------------------------------------------------------------------------
----
---- This file has been generated the 2020/03/16 - 11:19:27.
---- This file can be used with modelsim tools.
---- This file is not synthesizable and does not target any FPGAs.
---- DRM HDK VERSION 4.1.0.0.
---- DRM VERSION 4.1.0.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=128)
`protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`protect key_block
L+5c8xKbjiblp6p1goQ58UEQzmqrv7yH2Y/+xYypFn3ROjgzqPEfPDg0U0sEUXA25ELf+yHMJz/q
rPkRTZhGniuXVnEDfo0Rty/XV5S9UnrXVY+g1ZFEfhV/AW/4MS7JW+UznW6wATS2qdkmLUX8XEnh
g+xIdyPaS+/xQu2iEGg=

`protect encoding=(enctype="base64", line_length=76, bytes=839744)
`protect data_method="aes128-cbc"
`protect data_block
PyfIqqSHbY1Mavhyutm9yOALaWkzCIFHAvKNWJeF05EBRiY97J7s4SmlBldJzx3LhDO0axK/43TN
UTXysC9Gf9xd90lqFFTj2MzBXSutEnpdu9fg6zB2Li/hXkk99pknGy7iQTjXnGtCnlVi/MZVzxcw
iJb5RzaTYHAxDGw3ssXxFOdwiwHP7li9stFGpNInG/F8fSIWePWeKDdUPJhcD1nsoMtkHZaI93CG
plUoR9hzvhAguHNiEKczAOx3oTgEcc8b6aWpRrSVSbk8UjncQJc9DFZxAB67HDQboZiC3LFSrW9+
tylMsOUx6s0hyjA6Zr6Fpyrf1khOqFkGwpjA4EPtDh9jhZoaDfxznYuRKLC0QTtIbQD1nAoCvN+w
BRYHtQMEryHiuAYqXzzJ6qljxCidc8nbL2bw7DGbyu+ZhS4NAqbmmlmZpgi9LPX7bHGC3KqbIJ3/
0YNzI0kBdRt0p3uiOYp3gzIbnHwYTwziGR7IGS3RyclHxXrFhxuSNqnezSZrUvc/rekQpppL9sOh
IsJNb9/mu9OuB8vEfFrJ/oXdpj1bqSZtOVkjiGjYBCjeECWiyzVUgHSL/bB2wJdXmRrEJ11Pe33l
ZkJpqrDMwlNK4UgJwMddsOhefaxayuiysBjw6A4jP4PEyLbce1cjOuSUkR2g66dvGwgdL4F13Xfr
BfLMrW8qTUSmrDq1N4BxryPYXfMZFlE6YBGHYziKzKsqm01gVM1lIFook8Hon6W6R/bvcTQ8kOcL
knMF4oxwY6N1+tKz/utl91MMCQS0GhrO9012F/HZUVmIrV4wElWpla+deBw8QnxQXHB1VpHVtIsQ
OFbJLb2+a7qjxPgcR31fMePIYiGHU3w9M4Px1pPkHG6lGbjyGPUZae6EUuJ16TtFdro3D96C7Srw
CzvMNuQrqMOPMcvzGuH2R8gBxtLWU6Me7yg14ATd7HqeIIKndQ84+g72Nf8htNYsRPmU2bWfBZL8
T2Ldl+r6UpUoRWHgu/euH1sRmmQqT6kjIlTR+bhR5ausKrfMLY0E8pzj7JLQbCYWo83HBo9FSrRT
MEv2l+uSXdMdQtPCQSosNVVycgE4iVxVN9fUs8TmUeAlBqM3x4Vu1V75m4iT2gSCMGHcC/kFZTTV
r/OkQz9djKTlMoslRxYg4FkQ0rNLFLoi/pO86evfchZMptzwtgOxV9GHqBvpLUn8iNjH2ePSWUeA
rWuEuOScaqONxggekkd46lq/opTtrE5tInL37CLDp4NXWYr4aOLkE10g5aBl5xMlmI3OhTt6IZ0b
HxwGVkT5FbjkTXNG9Kfuu831ObX7ZyVv2s2Fx1jNYX9AhFWmhnzVDS2XTpWfC3SgQiSWTifpYNFZ
3+14GSaAzYHYra8GXuIupN4I6z+10uXZrVw5ctWj85KOxapnyyMWW56s+qfoo6TuO8/rxzv7xu7b
54tQHXbs9nEV/1ArwhJO/kLCsgnYh+S5GE/DDdZO+YJ3p3X1BDjGTgMKXGwcrdkLLWas6Ah4ZuRE
Ig6Vv9tr/F985MY3KMf1M/HAnKVxawwwDAkAP3FuMXqpOcXLz1Gca+k8ERtunQOsSBsdd9skqYJI
Yoz85sLE1/hAYOXWDHZTPIjzvICOVZMDmyDqfMc10SPaGjZHSd/Q7OfVhjpE93lFzwkVBDFQDLK+
3pbzPhEP0ZyvgU8FIwi4xd00Viplvbul4wBJ8ppyobzSPciCU+DDJn5IFTCFJ7UfXQUF3WN8XZqz
Vu5I7qEZr9QWFPWHU06NzkrWSxpJpTnME3CT7eUaCP59rFnU5os5I04u7yjumjFsjFFk1kZtvPeD
1cB0lhnXvdZuhnaXvoLqw+sfQqbpjjm40szOvd72uCa0Ae9A7tCXKFOxBbjKff2MMI3+80TUHpmy
ALhzB8EhjjJFjFI50XHj6E9OmOj7aEY21qQ1Ofj0kk0mN7glQoeUrHFPwerXTYPBulP6JmwXMPwx
llGSQo7mGi9JZPqOikVo3gcwR96hMFseMUCU8+aRVpUWsrbcC/0YWLCj4PxMsEQhhGJPmxSTTTUW
vkG5cwSZYGLrWmcSze/npby2Y+WY9pZCkkmnE9d7lgtRhMRbqk5y4g+gXT0QSjd7wjgSj4RkQqOL
Wta52fKGGrvIQLeq9msMlq8/J56NFGF2MIKvwdIxSZLkw5+oZJrI+vqcZMDDMYIUhoMeqvoLcjrm
QYWaf3wYhF6+9ChHURaOiNmHERz3j9pfIDJqmZxYJHUaBY6P76w+aR6xY9LQ5fyPjgKtcyaM5lt9
+5WWSJTHsFI8eVgInouTtkBM6/A8upK8vFB3PcEv/vXcBV17u8Q5TI35GBhqw6ZnNXxxmsTva9pk
2bM3ttVkCTfKFC+0Xt0bsNNv5AH8L+Mt6ymcP2lf18UD8VCicIK72MzE1s/buhDiF7o4Z4TmRzia
z60ikGLcprjJRuZe2KFfDIxkNqL9VC14HAqFOPUBaRHONOVhQ6o234DMqk0pTrOu+wC/oHXFPlxn
xfnWinC3YSR9ul2qYNNXNdcyVbuMW0aMpMoLVd80goj/t/jrfsAfefewJtINo/jO7PSdf2ye4oY5
XuVKR+dygSnBuWwBXv9JXb80ZlkwiIf7KDKwfZqrTkhbD9R7WnDHM5YxulGrYhIH+I9H3FSEFGSC
9VGkNsX4wnn7W7aksHjcgwlL62xnT+RIJpjH6RZmw5kCFDxhTzsJpM1MuH4aL52l+JmKkPwXoacz
2DPt70nDsr/SQcXQKqM1qgO4fCugr/M6dKNjGWBMDYm+Idi2D5Jn+tk/6h2uGeWtR+DEXYsiHRno
Aaw5odnxijbtoNWspa5HKJC+YYpJbpV9A0fWA37uwM2F5yIH80Yit8o4sQDA5ROQvIVQNSrgIShN
Re1zR2mfoR/VxUdCZWGDWgH2CskbIhracwlDbGPzlLjgx+ILjnPz65Hzk7d1aLIfz+LNmMe1FOoJ
/9if/AmRSKXm8mpGhsqjWA961gBo6lOlhLhpPiPq9L3+OywvALScYe0vvl+IqkfcyeVe8m6XizN/
roPTxBSt0Tth/3PV0jmhfLQ42K+KjvwvM2u8devB8mULwh3PyZ14u58cjqJdi86Zdpt18pS0MdFh
hxhMhGRNkDNTtRP+Oy9PAP5k/j6A+WLmaCRc9OznPh0ZRdQ+okE6Ji0nFmcaDPZPaVLH8PHuNCb9
u60CgOI99TRl4SWbWTAmm4RU2mb6kmwVO43qU7jiepkFkjMdxuigKgBvdmSRlcwpzkJOwQNFJ41T
dcezfeI25ONwXHOlJ7Pnk6746rjiIsL3/1GKnD1/7LwvvuJTmu8szbK1nIRMWH17GHQPXAd/5cUT
sOpznO0ZeQ3dwCeFTpPmGb/v91+kXZBHWvw9sxHmEYvIX0lSR0Ctuji8/chD9mj9Iyn4pN3zA0U0
9XIgPP814VsbKc0GyAscHDS/+7iwcMP6ZrT2BPcDr9VBhog8fu5nJE6dIW/ZHv2vKIr4Bft03GDt
xqR5cq92n7btiLHtr4zpjJDIJ/HzL9Jw7jaTeb/ELM15AVmbH6A0tLR7fppn3XZLkOLucQXE1b7x
YGKj2OqyCkNFzDGdoh+t5hgtdV51AjA44IXEHLjM/TymUjRmGvZVlUqa+E39y/ZpRmtxFA8YqLhv
OSUzS45xanwNN9OxsFkWBsRtrM98bkWQ0QTnkdqamkGBj/3H1VcLptUSxbwRAXssp4rWp1DO3qSq
OrT+i1cPvhXEv/K2X7BFfl4uTQJO5gTgyF/py02jJvvdYWafX88eI0h7+uhhQFrdhGyRia81xOlv
JzsMdFbwFvGxvT0KtTKp/xNVU089/lEoA3YXhSKNt6I9kzvxISYlHL3+ZLrJjsaCEFjQW+gtIAQF
dbDQCmvD2oVd+h3UKPeW0Q+lGBAj2xMkajDtDSvJJuNaeis8OdidYs0TBlf+QQVZlCoy1obAPMgC
qjraSjJVpgJ/mh/jb5iekUaaHhY0mQQafzRT8EUokaG/XyQcPwpaTJBXo57If3LZq8Wgp86G7xmO
zfxaXiW9frz9UM24ozINnAYiqFlNfUx0cPRijdFll4k/2mdTaiHGdTJkYOe2TbirrR3VabdhGMFJ
Ftal3eJ/xnHwqe2VnjHP3RgCh5jQ3+4j7sZ5MAaGGk3KpfN9eDaG160AK1rWJTtk63+GRzTqDyqi
Avt45/3Yi15j9ZfU4G4jpzX+KINBXXysIsHoPEnef1+jmH07cYn1bUI3wTk6nT1NCkUrIeT1OiDM
fNJaoKQ9eym9BrI8zUMjvvmC7X//zwftiq6dqdOIOEzPK1tPtLx7C4RYJU8lWF+yJuR/EJHwBC2p
VaoqtzAxxgNUBUOCL9paqd/msyJ2WxUDFfpnc6FDxywHYRyMyfyd1BPq/uaBo5pOKsEodsKfhHKK
0u5hog6LIk7lrzPvqg4TJoQzGq2f1n+ACGYamSkqNFVzU8oCp4Qw+Sh07Z7lBMSISOqoEh9enCoh
lG7bszXR17nQTnMDWVD+BmV2UBwb/patufzwg6PpIXpPUsfTjQiENRiCCHZC8HQJke/2wd2kMVXl
LvdpkEG2Sf7TJcqs1t99ZbTVj06fS4iYsHzWaYs7/kQljSzVzFCmb2um0b5ABcKnZtuM4dpqtcHo
HtPwmWEmCeZAyxRVP/8YRo/5c7qAEipDXTs1gqVXuIgfbl+8qX3CiAW9aJ5b1nUbldxv40I9UmrY
yFKUWtqUkBOKj9MxYQxUKAB5Ot1ALyEd4vBFyPfKDjB+QUycJ0ikVR+ZypxVhJTOn7QvL1lDDi3p
A3VBtxSexnjLGjwLXw9eDj8CXGX8thaX1Wwr161k1Wh3cl2Pg4Homi0ApOEPC3b5DySKtcavNM8/
lOiAajU0btdpE0YBAFF9cjgI1CO75TJ+5wY29OFJG4ZCfn80nO/clEFs8R3bPbe++ekJi0gsN8su
V3hSrr6rbEtpAyatoMLQ7gWBpBX9Lp2OO+s8O1O0SxoTSKtGN/VA1g1r+dK+GK7c+utksufZqa79
gVUKVM/pGKlJwYYoR5upjupFPaRjIDZCJiXiCWfCYZF/LqAwRPHArZsCviO5PcBivbqHeQU2sM0o
IN7xas/yoi1E6qheLJ+7t9lcRi6c9T0TIjyzKNyLDzN7YcSDPSchT/HUtRb7WrP38vd7yGOuKEDb
uYAaVwEWM1LdXs1LSQrPd9a7sBAsYOiK1bbRf+LsJgOj0JkY9XUH/fGK8en+snqlHZrjLBk7oN7S
AgoDHCK9nz0byMwW8OPz3iaAEm/nxCDug5Ifm4Lszd8myZTC1u0zpYgMur9JDVTrItt2iTBpnVUK
zev4Y8x18FmdzGLBFI1S44WTRYabIH1hjm4322eqt2ef7EjKIyKwoyGybtZ345z/uo5xMhAHzMiN
E4PMK5sfyEb/KQADT+yhPdNwGotoFEsrzOzrz8D+7bh6hY8J6CKSDZwImltYXBgKyJDwU5iIXrG+
ZvBrDRgAbwTK0myLAdcNjVjdjXTbopuUKByMl7j5daUff0DDbwrVux2UoL9nSZXTfrxsh+l2lfkr
6P0We3AzaIWVn+a7V8CrSfouHTHp93BGjDcYQkZ7OWoQVg8LKXo78AaJZ/3qA7Rcw7CbGgR6BR/I
NwmxP09yJKSZhLzZKiqJ2OBCty5QBHzeKD/i0H1a/OI0u55+JLw/qfdjy6PB/VEyzkevdm8TM127
A71a4z7PqGNpgs4ZHirC4ZX89mUcgeMM8psd5ngNcX/xRoHH7BIcW38EgQAER6ja8hSbdrFThWAh
lDDYAZ9NX4Uu9XLSLq2H5U/UOz2thKz0TLreJdlwZIu8Olf6Mr4HouavL19C1LxVIz/isavVnFH0
XCmWHFZpUL9iR5+B9DmnqYgEo66xU86FctDEdV8bMtHj9j2c7Tp3i1jCqWiZfYA1BFM+W3yPk6Gp
6w8ncWYWYvSAIQZVi818xemHRKMXEZ0lIZ+mTUfkG/MjXyecqucBemeiWTHfyFdiDsFn80FL5QQT
f5ZYyr4Bp1EsLZPgEyWcfluOt/FLWSLSIsPccRX5N9O9W0VCQ8FbPKC+Y9SICyfE63lt2MOnB1x1
VPeIPufP6X6VnSM3u3gkmNBdpCQ/a3NJqJgisWbD5/ZQ7PLBMr+Zh3F0xZjBNDhIVu6a3awmgJ3J
YycPB9VrCUqcWYZodMBAJnDkQpw/cJnTTk6sRcPv8CcOhcLRT73KvGPlnfOiLJjSW8ppqP60X/eA
VbxQLVW3RW27gTtXz+ZF4PRmxuxoE0oRvyPNu2wuEYO0DsX0mQhMYTllWs/7Ez1pZAhrim0XX0g9
anJGhWUp2+ZkyLWayPJL+38F4dh3jHzeH+s98+7/AqBBXLvHk0ZX/CjcRmcfsCEb1AIGgsqUfqVy
UQV/YJdo6ReqgNq8qCJjqDUXm+EzA3BoSA0CX9Xek4Lz2rWVgaXubS69Im/4qVjX/brIErHvek3N
hYc27Zb7nUKNObkFTau/Muw6FZXYf3sARfhMHdvx8ANWZi573ZYQOsxFzWk3Z1jeZHRdjp88VckC
Oz9Ry7TDtuzXcijF3UdbMpfV0OKY0oEdmRi0e82i1bpuIVW27+xlJQE6McNyB+/tvmm8xgp9UxGI
wB/Exx9cm+7+dm6PwMQJf5gMYtjCmcXJfeQ597BLe6TvTGcoqVHadDaP85XhmSTW0WMFg5y00b5k
rKWbs6S4eWAoXKt7YnOGjWOz8ziepEQ6EAMyoiBtRrAL8zLkoC5CHf1HEODOCv+AOm8BDWIF/wQh
z+zwETImVBtzfd5/N/ZGgg+2V1M38CgMTqCzLMO8bYErH7EwXMHmLawoPSk3dvyVWi7QFtl5TQ7z
SmOiim9eeHbqo2C2f8Wab5Nnu6XRa6yi6Zx+TR/ulI3BW4gbbmrldDowLpI41zeO1xqadSzzOezF
5foHt0GJ0mJpnlZSaMoJUTn/W0juvN3+MUlU0q9G0aTaLz5wu5Ym9JE3eleAcoITNA7vDQt2NIjP
kAu9h1/jYt25eRqFfuVitT6HnfJb/JBbu28/TGWjC6sNUfwMt+2hlqZbhDPsbPMCxc67vBk1yp7H
h3hwEcUHGGJfu4U3QPy9pNoGZlM9bUKkj1dSlfXf7nZByBkhhAcSijx02SgKuEE3V8wAUZRA+oDe
90VRGNVPGzdMttAfMXSMM5/er2iyOoY7Zvq8SAnP5GnEz3sbPo/X3hzcF/uI7pwXYZr/gcRJNIlt
HguuKeC9hMUzF4v5uA31a1KMMQBWSCqurVfBmG3p4Tu65kNH49A5EApB4h5SU+TGSLImWmYH6/DG
76lW07Bw/0z0HOUIwBC/vo+JzLwSfcfAd+XgOdpJrCXoiORnm3wgBT3MN/jTHCzGx7fmmN376HFA
v42y+vJANqp0AA+w7snYUw//dlfY/9vDK+mtGeV/REGRrW3iw70tW3/Tr+wczS77W5T5AVQG4z18
VX6yhEU+6sZ0MN0PdIqR8sxEq1UeTdnlFr7xIjzDE5mHj5hPpEtdhQM5csrHJlkDEUyqqjcfrbi+
jCfQE+QbUjZ7xrHr952pIl93kHW0tze5Pyfu5TEd0foWPjFLkcOrw4JeSCm26zVAhkmxWRAjn6Wg
vkbZk8s7+Efu6tV47IkXA2H6m99+WPibdWdWRycTBwQf8AqFMbVqMNl6My37E0cGUfUhiyS4Ve5i
CoUpRa7JcrcXtlETXdscOv+/RIVLwToZc/T96xjmFGFvSVrQM5dYt/dYRzm8jnVCue4T5jhz/UYK
s2fbxyTcH5AAZ42/WSOxKMJS1UoxDYeRwIiU0EeQuksr5/54d8nGPwM7NdlFoW/hITdtFkrKoxk6
dnyepgbty+YapGhI/F3E0kWCq71Itm6VqqsqqFA5Exx4zF4DZooNF5rAktR7IZszNF9j2zL/ld1N
HRueWFYxMN3H4mNc1zG8//51TXnOGwvsGx804cStGMlOcW1JmB1TglWx6v3aYxsv6kl/R8B3PxT5
e/am2iO8XY0DQwijbq2yiH5oqrZlOn6u859/+9sjExUv+Fwv5+7Niqe86X5Q242MG5GMElVoOX5n
vdq1YjKQpgTwDj43EaIdCpHwSWQ2eo82oQxTdt7Jk9Kt+aznUOutH+tCOTJV2zmlq5lJy+uc9uHb
vHj9lVYvuGXaL/zKFL21i0l2K9jlWdrc5KrNJs5puSbSH5ZebZDFVh/yBpBnr/WhwtUEoP4L9otZ
s10H6Z97FlQ5cdN5rSv84Zl4QtQ1JILpJcDWq3f0iInVoT0Hc87XRxsDp7jC/iNSA8850jngHI+R
jy3JWu9JdocPiXHvcNQTzikFI+lUoUOGyF7vZNP+yJ8NVZyZS9Y7uFFvgCNy7Ar+OSQnnIXPIQp2
MDbaZdAo/XcLluJXsJELOnIrMlI4JPOb8SMEkV/MISs8cHt10/ek+EmWE867wz8pdsw9gbzlZRg3
G524igCS4A2CpcKDpRaUDFkPAcwTgufhl3uzIy2BsbtDMKfPWMaD9SMNGu8yDpVE5g96ouc4GdpE
MpstmuaNGBqOrciXIWirxG1zITKJrOAnsypgZdIcjYU6aHHWUdyx+2FLEkBwx8SzccTKD7HN1CaR
isyKi16ewuUXOaXkfsJj8pV9xUTZnCuY/MYsp4tuNltTwG/q7JwGsc8RheUavwy9rWUBwVY60fDi
47/RDSqOK+OcRkko5Kal7VVeia93BqQFSKGACMjDc4BG3M9abHfweL/5FwHOHzH7kGMQOQfp+Lya
fBHBSGYHOiJ/bpQloLkZwv1Sw/LzWL37BXxa1p50Y06/uc5m/DZCaQvbugxPvsyf+QoAIlqREf4a
CbnUpZ3sc1i60uvtXlfoWEMBK0cvUEArGy/L3db6DocyiCEml8p4QK5iNcR9oB/UGyOS7ZE9OW3/
7IqmbREJNhzlQJZdMjq1p5trn2AWIg7GA9JCpFzi9tgOkbxdlBMYFbtcCcXmW+Y7c5SexAkBINDb
f6adeEwLaQ4rbETBVtUuxNqItpsucbpQM9KUxNiuiVYgIGUbH83jsIsJO0vX0KzugS+pIrbdTB+q
YYIZawh7jJ5UZ9ArmTfeO4ztGx31nZclYiIo2smE3mJbI8TJqCKsiYgKbWCDYWOdHtmuBjl+xiEh
CzWJ2gUlnVjTYCypjkQkP/TpLDM1y3J3+9DX3YDgB/gICAk5BB7VLyWKE1hXtHVdW6gP7lo+s/6S
Bf11/slvxgIaK6o6bRUgEDXOK5oAQvsxLB6bwiwcyl8DB+15Du6yA+hN7SIOdqOuKf+kLfsndaGN
pwDNgvBp27QXhDweWi+ugpm6f0wyyF7xali1krBZ+kJytFm/JsYmo4elwpG1MhkGOalC49iZITLv
x2EEVIGInDvcX+Aow74NMhu7pV+bpRvy4GXbK4PIF/ecyRfjE9K9l5FDEqrBvzJxemoKFgE2IqSW
kQUC+TKY4aM0DFm2Y2DjI3Q+y1oSxl2SnTpbF9ncWHYdWiHEZDk8h8NBvWLXsz1v/th1wDgijOQy
sRBGbDZk6t5qPY7rQCWFovUzZDM/4jKOXKeSYf7RkN8EwswdwUMi6LQPI61V28yupeTFpKz373d2
kMCRzqANDs3M5I/djTLgwaT+rvY5JguNhGotrPyztu1kxBm2dmbJjXvW+yKRytSFdiqDztRTS5Nr
ZKpdV2UhRehGbF1n4msKYC+XW8N7lMjtt9HINmV3T8Z+dOZ0D580iwj5U/R8KCuSHWJTHL/+lz/Y
WbjamD5w/ELIEFzJbZXgIIwOZIwgP5vopnQYu6nmhABH4u+E8PIHv7qR0HCmYiITy3CFfLSF+yzv
1CXnhirBPlAjvhpY9Y2WcXiY/wmvkKWRk2ssmSTdum96PrJhW++feJTdK2L2n6xqEqEv21ddnjpN
GwAQF/PafM6vu3GZ7JZhKjN4mnDRP2ptzIh+Vn4Ch08cd0ANVq8zy03ry1H/w4ZZemgj9yPNJdSf
yR6rkDWQJOFUjmCwvI921JRIdch4yybJZcqgVcRQODE010bYVOsJs5bFu9odF5NIq9nAIbFpH6Y3
5gbm6q19kR+00XgAloE9RcPEp2p9+7q9V4pL8kXkvjQdkUrXPFFdB4vtqjyPtzh0/peJqmHoG010
/AGLtHMmeh+qAPY3CDkuN3EBqWxoy/2MERRtRKAsLzT7XlYm1Q6XoKVCi7PoqWTzZUC8kRJMDXNt
ati/fMjrAA4ROLVgfTbCbYSvEmdf/QK6O9iL/Ld/wxN0CVhOAZTx/pLbpgGulBP2s0qA9C9s0W+4
PM32Qd4OtaxxxkQOJYKzvGOYcpbbg/aPrfG5XvGT0iKDpTXEDMNb3vv6z62cTmGEm9iXIleCWqHU
/IFcM8kLf5N3Tzqhn2c31lNzGoRc8ZZx0PVycFMxIY3VER/PWns6UOWiFfa3ZX6RDqqeGihPpSOF
41TQXD8aVDIMDtnsL9CkQjOa81Cm3MsSU37kcLPAmX6iv4f533ZLn0HB7GKcob0BqYJW9NWrHbY8
CKQbZ7iuxysSW4AAli2MERQDpugZiPsTUB/ZKUBs+64zpyN8jzZIWHinOnYy4KqH66NKcflBFtM5
MxsRRyETalnwOPxWJvzBIiw1f0eL/8KBKhi5G/HP8RFFHlW9S1e/luUrUqQT7eB3JR42zbCXToFS
IrqoYQMs0BkwQPiELy8cq5LDF2mizZXgiX2gcCUiLXDpiz+lSEICWSCVemsDwFX5fuqRPzKji74d
B4QoFOu22u2Q9OxZCoAAGNCvu39+rnAd61/MRTZzImi+H1tRIykcmqVgnWEkvjRyNsEj3JLiJFBY
NHK02Z6zd9Mn6ypVgZrrMcKnNO5StKuioDeKonpNfGp3icUZ4ZQb287WoR8bnuU6SKjlbNL0XW80
WxlElzLo0BT9M9fN+bK7ryoNU+krGMVDQHxTpSEFbmdFzAzPZkwsIcmkqaJJ5bXWv5HqiN16+2ue
kXR8muprMEF3GFkt+fBHenBL2/lnZFKIkLu8HPClmBFHUrA3Ip29oP8ilbDXixt9u3uEjx9O9jXs
HOoxaiMZWXLUNEhGqlBapmWQLfkYobS4kbBTdLfWgM8ybLSbiAjuY9X8B2uIkZsnob2+rLOLx1u4
zCRg5OjQjvfIksiGMo8kkar3HDtXrKrp9MBm/iMGJxTndB4bLhW/jj423AB/wv912wdg+Uqg5Xrg
1MkZDrpij6BVf6DvStAJXEkvOZofQcaQho/HYW8e5Om+hQir68Djc/y0Q4fkbnM+8JahRhqcmRHF
IsyRmQ09IKN2HR2lOV7KelAlKZ8FBaVXP2XziRs2h4jDrg1+4/8mvoA3opLs+PbiruWosgwS9OMI
t08VbXgU2inOnQoc2RtIqbtQhUUGxc5pxgR40iD9Iw7AQkvVnox0JhUbRnZccqNNibJODaEIu/Kf
dqUGBy1DWuklkwpGBzid7xNagsYBxRRnto9fChYwGyp9w/hAlf3dj955FyL9Xw/yMJYyr0KATCPV
Up1GlbDnOAck/hLoJbfGnMVump7tEoESvm0l8YtchbhfFN/3DQLWQ+D5HZfpxh1tSDqGJOhqUxs8
j/f+CRPpkA1MBh/loqJdIp53RQC8S4iA5Mxe9NpjSB14wbkPH9mmZhBQYJaa2imUuHv0fdMSvIsb
pYZMY+VRgETnxIGG0/olBEn4AsE82pthCj9dm3Tr+i9CMPtRX4gKZTFw9IB+yy0akEl2etNqdB/t
Hu2R42RHev2yb1Hn00hFFqTn7cLIDvjIXYSBgRIe7Y85mOS++Ud2SuYGTbYBFsEDvby7UGzqzImm
bkkftQSSApjhm/GXdxw7JJoo+1H7GkTl6vHgqXns206mvAaYdjwLs5C6wYsvH4j7KMTen5ypkmcm
PTtgiCr+9TqiA+FJI89vALgPk02MM+hGKexVVBCOjFZ72POjMsR2XWwyGSXhpsITx6Z6rKmX8Nnh
QAcircxSLLBbXM7OY+Es3r6suKGnRTJB/cGdUwWBQeEFSHTp/iRV96HOamxiKyPwYVBeU4xHCKRU
IAgbjJYmen7tfMbtim8JxaNWEdSmvjRR8B+eB4XqJfMIrHX9WpHxwItbt0jTC0YHJHNVEFbX+omD
GyfkofilbZje0a3qrR9w5HJFv1Rqf+7GeYBzn7E9SPpnQByYJaJjJWQO4Wq/9W/4XlObfMVryDFA
HIZC0P3Ygk5aZzMXT52TiCd2rvxXg5vpeqsZ+V6GkKj/vWzoixM9scYjNoQfvPoZ08usIOBHJdYb
BWxfyUWdErAcfj3Ybq2YPhgWfzWDtT1B1DDW02SFTJQL0GWNLberVhKzMaHjCQBnLp6KvmuHKa1N
UKD/L9HcSU7WbE5alm/jPWZF5YdWqbksreo8s9LStdPn12X8L021QK4qMZYsc5L18kyGZMbZog2U
qWZPnNmYLU1NyU4szLU8fCuCpG6VvKwOqLnd/jZ+KMpJI1pyE2qPcCCuUu7O+8NnwqX56ad2CqvD
Rs6jkMwcVyp8vWyPm1PJM0U2Q7AREUONxMCNSxNG4FUWRV1KR35gg5M+6kfJQ8js1hMW93MQKE1F
oPwMhbiROTPyF2sddD5/Q1RYS9s1ieYOlffU8ZbqdHRrJGOrpFDtoYpuK++rEYBQHJ45yd5FgA7Q
ImCCcvWK4DAwXx+r3pSs/XHwSK0gWXG5dX2NsB5l3hCQvTKlea4skoAz81WG64eiBeG6NobH9d75
ZRpn8iVQc3cRQTcCM62Ky0VCIM23ig3hfNa3LXHxBWwLFL0XKjopDR9pZeZZlrXrT6J1Tr8RubzU
0eIYyQ9yOF1xqHtsxh7RL3q8qc8xe+nNFSz6tnPClMGkmZGAGzewwCsYTF9SEtHmSZXECtsGX6L6
NFh8sQWMrr+2zdLY8Y1FWg4Nb5fmlfGmCVrF/mfkfB6icTkda+HScnDpYcmiQhKUJ2RXz/y5fkhA
EWr+57GURlB2Pb2C9LXlkFFVJ2l2QzmsOk/qox2QrBtxl0NVVqca5uiLkCfyBLslkaX+yhgNw4KK
9GHcnz8Ky6BBuVM1wHSsLHp5exVOuYZeivQs2WU1AYGkbT/RbILK6coi7+aabVL0vfWVjYK6Is09
/4K6wImMed22WgPx3VihxRvaGJUkZOz94veVQ4bSqX7pAyIdxgVBQlJR/qL9ZSv08HjvymsvXn+l
BURd1EFwvDBavdvp0dg2K+QS2I+Rl1NRPDh197UlAob73Eq1VwpaaZ2g0qVdUKJi+y9hYHUkQipy
GMS+AuJs1RQonx/FVq4+C9/V1Fj9mLvcx5LUeof/hrYkUqSzDkhsNjviHr1nwKf9lJZJSwYT0zEZ
sXZoGzA82+a5vQp6736xi27AmDmxlog1JAtxJ30SGxWTUrG+15aN+dKNThLaTf4gz0Q3Ngctbbyb
GfMW6utVkoXO4MrFFhIT2VrgmuvQ1JQmTthsH4Vj3AbF1Pn9TyX/hNeUmwyluKXxqjVWXr9jES0d
w2m6cG8r3nGCWEBuH13qoe7jRztK8iIvwheeWFJNFfsYnVowMYV9bqRrKl20gdYzugrKD7aHFcZR
nP4++MoXJ0hxSPI1sRYaD0U6X3dHp7Xbn4awAxqzZ6KuAbjDPgz1tUWwgW5wsPvUYLe0Tt2IwTRe
vrbaxJWV60NP3+9hbiht779gqz3zhrtZVrMZf7lHKqV7jauymCArwWf2ZblaNq9ERnUxHkL7I6gk
P8pxMWuV8mWANLL3mAqWXVSq4VleiVEPMUFk9Tl1yzmONf8T02SqHjf19GI2SLoGb9KKcFZu6usP
4M5ORW2k3CXFM4Dq+tCoZiEFZyXxjCRXfmXK6mLpJue1IIqDO4w2+KrBLQdAnVL6kq3Qqs+D4BU9
v1yc+hgeeyT/JXU/mVqlsGQ/lIMNBs0RKToSJWEyR/HHomkeyUC3iKOyq6ph1NnWQEV3EmymK1vX
9kck20dMhl7mbrDhNm4THF0FFZ1VROhCbQ/KpBv5eVbr1Xj76qd07+l185s9H49hlOuFezgGJQMB
JfpgcI/uVGY09Y2NNwALU8QmtJstvtFXhXpe1AVHI3kXTNH4KGpLzM+Brh5C00sJIjld9YhF8iiR
OrWwJv/oC58pyC1+r4HKNNuU7tP0ESXuaO8CLcdulf2nvuMwtKXjPVgu/cC6G25+7omo1+WyUXZ3
HKMpjY1KKEQRTTcaUwYhc+Ih7kVYx2GYjxqqCM6Lsn2BWmOdakfSVEcO6uKeRy1aJ2w95YbU/MZE
3o6CNzLA4R0gZjyrS0DGuESgntq359hkINzaLq2aTbcE74j01/lY0lcjHI9jbJP7N7sM5+5h8vqM
ARaRj5fSoOqmPG7LsLr9q6KFN+c6mskaR/9xbGz3NaIHreGavibFp9ImZsQDs6C68g86N3B6qfg6
XuIHX/G+dHlnypz/UVUzagGxvU3CoI0oNpq2FwMmouQWGQbvEYs7xS9nAcdvd/6sQqLr61qB191c
Dn5nu/NRsLcgi16y6nNE0DMEntcN8zcNf3fYVYPbzznP5XGjmpS7sqOhJNnCgFpAty6xSFTLIkj8
RuX8ljNMGj10O++ftwBZVeHyOh53soz8aWhO3xgBrHzs2cWJn/1AFjViGMW3ecB2N7Ty8BOwGie1
QCHrbUzpWPOyEjsPQisABl/W7XFOXAWbi9LOE6JqGw/WmA2tq3FtdDySyr2uoWwk1gTIq4rRJfVF
3r7YyGybkLgsUatdCEav95kkBACyh0cEqUH82BTyMLecL1CqIKoqYblVuoGe6g7ayZwp28ANaofQ
VIJZoMftwZkq4uEFMbF0GDeNFHeTixhKCa8X9hrKRvx5wUngpomHZMAJvXUqk+m8Bq426yBo+1QM
hd6+tmNxYKzYh3KWf+Zx+h7WJQHAfVRN4qRe/vyA+mt2/8FSVcYGAbVHkt8hQJD22D+WldfpV57d
HW3f0aOPz0EosFBkzI3BeBiG7Je3ji6GN0s+qwYEqKOuirebuSpa3/zVLlUaVCq4JJXJMq2PANIq
Mj1uIelMWzH1A8HsydYjdXQuvs38W3ftv4XpXaqDFSjVlusbjrlJQNRfA7yHr3I0aD/8DqqhNcgp
BcBXbaYjmwajCbLi924YXT1w9vB8bwa14jT83tu62QsYdNiNA5yv+F5fUTs7ZFyGNpIfkY19aLKJ
ihtkDQQAuzNx3SMKZhNvWjH5BjF+pVkXL2631yX4gdqqRDDZ1vD3OcuqAIa2C49aP53QoxpudHxw
bjar7uZmBcaDuliqgB3nnqLJzoo110/DnqEqKt473z2s30rsjZkhpZlIYqvhGqOda/BgTdfNEhE2
DfVgnx5/+QJZt7IHtuZWuFWWWQ62uzgZZVtxIPJvtPbyskb5ruacMzXLXKRAjoPRI+1gOr49mDS6
1nhssj47jCyeHxUopx3pFD2A3eGSPgfleFjwcflt6U8/4M5oH0dG4i2VY123KG61sJQ38j1mt/eX
tKwkCclkdfBB/N5N5iRTDBLU+MwcuOsAURUQqAJ7JW8iprtVrvj9K2WXEVc0KzEsPJvu4+HvL21v
jZT2ML4s99owpB/XlaFrUFauhUeWhQkq46Zxo42o7SHkVLbTpWevvGvwsIdeqWl/+vmD1SW8dZKR
qtSwcBDa3CyW4zlOcMtzniMsF2qm03YlFSPuty0rdBrKOR44CEAzbQoVFo16O9r1FAGIUHUhzcbK
lA7/2HvEEmESelMIe9V9pn1eIfUTJ0czpXFwp3VHQnJt+5CWlkb6B1UmmTVAfMuf5pcqQnjR5+XC
qP9QY8tbKvp8sqnQSd54thIIqYkzn5SgWtfi/O5q5IKhLqcPJ5X5te1rm6PJ92Nux3oqCtmyMaMX
/S/4VZOEvWsMP25B2d97IEw6m1cj1VAOCPnnTZxnXQ4Sg/JfH5Eia9ZFxtkg/ky+XLgVaQ69eCWJ
1KSGn9w/7ahAvjXeWxJn8yzlnRPJbmQWyEu1Q/8EqcmSD6KYLUicPswIpkBdIy+DnINgQqwoDeIk
sZIOX/gPWB8hXcAN9BuQPGnTZAU1sakuuSh9EKCk34jPnB++vwcbvGTCb475MaujYLTTgaVuqD/5
6+G4FKpU3nrqFbJ0BF+W/Phpu8e2LvK6ybIQMqnibDzwe1XUoxxq6uCjm2gNDHl3/+EAKNQgl0p+
iiAnN79ZgIO3HLsd0hpVokYlbfuvPPPOW2rh2E6BUbAxRI3+Qd2HuYMy57R0aGT4H0z0c4YIxUyu
NirZsIY4To0ydws0LuGyU3QrZpxtL0AScph9BaIlfU1eOz+XUKY2KjR5f2ZyuaXK/T8HNm90pz7H
79k39cKAwEEXnpiEeqdG3LhFJVeMN4sbXPFDXbjrQaxglSWTw+3wLKLhmCSIsWaV1uLpnGeoRR+D
uoWGBw4aS6xMtysKcshlvniZV0uJEYj6x/NsS6ZzxSQF0l5aNUvqfbVoXLKDs7pPxof1e9lXKXjl
8ZBe9SCq1TOr8+V0zHB5Z07xM2vhmWDZWSWUVwT1DiCW+iPVKq1aPBkCw25KvQxqFYV3M6Teun0X
rfz9puJ7K1gcj8+byeIG3maSKfJCQcakmxAYPxCqarxCm+aWSVagk5ToxmARbKvCbsnfeO+p8IuN
QUYOgvvl2z1sRaCFNC7fVz11QiE9oWVasndGirghhH9cBYgb/awztShb4qKKENblJnZB6H57zMgm
PxAYrb4802BmGL7ixUkygLAycXuE64uyf7Ad2RP2Kun5sodY5I6oFrhTBhvjGT/GobPDBITNnHS1
NCP7s0mxNb1O21RPsjwiRlO1swo5fQf47ufNYWCmzEm1lGnyRYniXsLHL+g2CVbDkgUAdHQRIth7
XtiryuaAcxysVrNGjOPritsgLWeOGE/Yb/BLF86kQtpfbLXF069T565BE925WKd5P0bcBqQe6m5B
ew+sC3/4HLKjT2/kYkaNXQ8J3v4I7KIkJuPr+0ebeS9xI3tiw13dFYibRiiYsalEnqZAu5dLbxfq
ZCki48ZuOQdvMzWPfzBY7jceRmpq6NKS+fpvVo+VOAahB5e30nWncQtlW1t336L+KwRXvCJaP3Bl
Pm8LogSd2oRZWET9g3uDH+MM+JrnPlkIAAAoaUpfvZXt3VJvLn6pSkwuU6atw6JCSEXP2nIxblKl
9TH0jHE6UP8sbtMC/2R84j4GUTbxkHysi6lY/fReB5KnKJcC2x7lWv44K9E9I2LcCSy1pZwCkF6W
XpNs7A4G96Q9ifG9vDfN6R31tWIOjsygemEekBbmvyM4EQfWjh6UBl+qLSp8js67/1W031RRLF2z
sfyRaUIlBX4sabUPlimziCIzaa/AvvP4OQcUPkI/1iHCIZzrs9ROgjMbx7omSRBPq2Krt5pm9GnZ
Nho3bQAngCd3RiFLX4bYmT+bkf7M54xqdq2HGbWRcNj/te/UWvBrQWnPi8SLazIb4TcYN2KFL/om
wZp3KXNhoe77pLXDIozNZMEMzxYM234nwlMxX+ywzriAtfr6K8xAjK+NR9gHjNHuwYUuSIeTu6ou
hC8zoEjLeB20UAjaz0klgOVwhUBRTwQcXFeQSzhO7nQrPE10u4JA+zqRavEU20cexlKvulpg0HuE
EdNuQF2V7HImcsCOVgK2H3kckW1ajbjxdtPlHc29UvSKOT7P9inuwVE25CsVtu/VyCZOu6692dvE
gZ3JxvW99F0CVIybin5zbjxsIfFzJrVPJI6OxB8CtnIxWSYKqmx2C8aXODcgrotFtrN1/8MAnjQt
hlHarNqe9Qp6OO7pwJ/2ITG8fyH2UVrVXwRPevSePgXpJPhM6qBxYve+cw2Db79OZQUe76uL2P8H
QGCgg5HH0QW+CxhRpoJeawF+P4/MHY25TiRzNk6iYHL8MT2v7W9DORXU5/Hj6XEl7isWgur9Ai66
+L44MGVPxcfwViqPRygZGECCfwfcA/se6tNPyoLM81yA42R48qPO7rw1ePaLyjsoGsmDbab0vd8f
e903CC9SO6KlQDfN3gKwYRo18DKxsf6olFpr2IUbVVwpKVLAjAWWDTYAlKmwBBwjJANNtjs5HIfU
EPHhLoqyQvb7rQYnWMXgvyTnkfCvqiPbJd6OPg7BVebvsDwe+ISTTI9Bd2UPbUb1MsQz29SR55a9
hvbolBTB6qlAlfZnuIbX8oHIbukOef5VmHiIGqi94PYeKgr4yYGFpYQjrbRo7HiJHvXtiUrS4/ZV
lbeAfn/M0eYvPFoGbL4QlDAe1zSCc5cDzpeXwHUhkyEcNoWSbYE+pNy6A+Uk7i6iVwnNJc/YRlSi
5EY3ptVPm0U4cO5vmDOXNHFEtXcAx7NtBpuGIzAQpBNMFU+EOA4geBtxGbVkEtVPHFdvV6KOLyOh
3PNCswqz/qB8ApFaSgKzSrNjoSKbGY3R2+Zvl0rwjUg0yNBhIHkJFvSGGxdOcQv2tsrr4z6tYnJN
ODBS21JdKjkVhVM6t65dmvV/Jt+qQZkZIHSp9684VdwrNA3lQ8qeD0mpNkpq9VhsiWSK26wSF74/
KR/r4FxdPfowhWFgVyWEZSs9H3+5IuPyRaxBNKgWx7CvOQhBmL4NLe+CbanO75urT8IvaiDRmTjS
MXW/RmhWs7jh+5fXLMd8z0psMzyqcPh9eLweFoy1DuHgHW3TrZPGvDr4Hfz23i2itsz3AM93OcqM
i6YEOTm250NAxmef5SzK9E3Wt0HoH0HwQblKazsuNB8OziybAOJQxfv/y8YSkMO5QLVmcnwvT5Td
nNcdIn8nuG2oJ+pTrGw2ei3owoO7mXM1ahiJ0Z8Fi9/Sjt4AltzCIoda7jhPxY0PSPnh8zC5YRIb
wZeAY2sg7+9i691gCCkoh4lxdpa5CAtxbXeayucKOZAgL7YMFAhvsfW1QL9YRMEzQKSpjOuw1zWE
I33idqLLt2VPqT86Vp3xwyHlPakbhrxy+TNBzMhyxaf+CaqaeEYGpUXGQ/1HEWf63myMHvkxXCUk
3ybMM069SMNt6PSaoWL0+PDJXktIvjopucUpJx2dDTqhOkfKfC1GGl7ZufwTOMmjicXrSRpSyrq/
6eiDrSj4rY4lO+S0B4erXfwHorsT+wlcO4vuGKJLNKq3CAQ35OWOGiZlPM+KZ7a2bo4QD5E7KB4V
DVV6zWArXA6URUy7kADGjtAWmUITjx/r1OFjgoCp1A23Rw7Iy0V6rjkcZ5Ar77EbgQZXT/TkJpod
j/zRaZBk8HcbKbT9IYNXU6XgPGD/nJSp7ygefeeospP4teTMA1xUXa5+k45m9uc6TCASHj4hKcrj
/mXk6Y8ZYb7PuvguJN0M5E2po35AEQOAS8p2IFr3eI2HfE6o/FKp/qIbRNGs5su+zIuR8TyRweVe
XPEccLTi54v3mLDreTrxDoby0gblsNQ1OdtU4tCqETHOEjmTptBNpL+kb4FoHb/0/klodNf4FEhl
nlJ30NBrdFCH+JJxrU7vOwVruy3dTmAIyyTQM7CGdSWi1Bhx6v4jdxSjj72Ii6CfHl7cKGpzHUSJ
VRKEesV+iSS0cJxV/dz8osmIW1TP2fq4k7c6J/a2dazx0Nkw80KCzHFEM+bGCPIbMjJxeM+9Cqp/
GVJgdkfTQUHg6uK5+8/uRqwiWR3QSjG6gOunY9yMlZC7P6957ynYap/cC/kCAmm82ko55lbmloKw
R6wOrd31yuO9Atxf2p5U6l5bnC3rxbyDkwdH7usRNv8OIv7I8C5GoqKX8CEp2PcftexwnMogW77R
bBoAsbeO21WQvSa8DbVFh0pw+zUpQTLB98mppXhpNhW6iISjmkO3NgvxbtN5SChL6rhiHiyvqQZS
IcuafDh5yJ+edtZzh0pBYeP69qcrqtFZGYu3e8KaSLeDvVwFBX+OHVKsqgDGJ3mtmwbbJfifyYmC
Bk1n/HTXPlb8ZASlradToRWsLnWYg6Q2hEPGmlYgEAmX3hiqZr4wnXNj41n4mskX4Ze0gFl5VmUv
zBBgAbbcycOguK9S50PxghtA7OZmia1RCwUphWu6GReOuiFK3Y5HM+NgKXSqtu3nv1ZxkRcshTNd
2lCLKEMB5dh9SshZigT/mlZlL05zSYtk6htF61alXmEsLSc6C61SfX8/IUKE+2uarJFOMtxC7Ove
G6pEVK+vjmMGSyfhQbg69UfzBRNvuNvHs7f5v4WcSanH2IWC+JS/WTQCi85YYBPdM3mXeS09f+GY
h43CtIvK4uljxyVFgL3KPg346BYgkFxdFMf+uomHqkc85bjFqVNxw8khmjN8qOcxFqXP5s8ymhSq
7LedQQCOD2GwOFuYgX0byIsJZvOBXiFMuPLa+J4e2jK9HaCNz6+8SLzJkoqHosbRnV5jfCqJ58b6
3VGHyvUrZFmkPbcdjve7vJU4CvMthxWsjrgg7mHRiW1DQ1298QD61PuVlSCLGgJwHpjv0jM8rDxH
Nj3nYc6wl/9n9CWspuA5e9Qzr6UjWSUuuYg21Aj7UKCf+NgZQzkcFmdPT2ynVvizCi4UCOgb+ndr
dAXCNosZUlA8oV1iyaYCtJ4mlh+Cq2Nn26w6ATWWLb8xMKHQSkRPFpq7PATEzczn+XhVtCeXU0Yx
9MaftN/PaxYvyv1nhZzs1YsiR9lG3yg7W+vmkd1t4BYTv0YrnhnDxQwvvlxoOREfOITDjeKFBlr8
GZhlJcxGT/DxTwjU9t9Da4inPoh4eJmwWh/i/O5SQQ6jEhpkYyXDznwPeF003H9EYOaAP9ReMhcy
rAVUrikUcm8oW+t3rrljMBT7Oo9WxgSDgVbcpJ/Ipts3TeG3imjm2+9CUyB/A2e/IkwDcVvXaS+p
q+wkefBSDneI4SwCzstY4u4xseEJZ//utgXxpsU5wbmOoxafOP+f6LoP27psJGmH56RuovC9XjWr
14A+F88LJUN7bhqMKqf/hPPD/8SsOComUCGMaCBeGI1t59DuKg6nLnmpFCrGCEU0SBd1Uj+i/CwY
KNTaU4neTi58HwVwZ6RhiwuUcc323CI8+S+KsC0k8WvugVR5YmEpT3iCGdqOf7FLqhwJzrSKnRhh
Awt5ZObGCkRrZ53qcqwhB8xNBZuPnX8liNAvdB0B24OqYbwwnrIoFnlvfcHjZelewOyip9LbRn6Z
KPX/wsrFxR6vJ/mpDABZtTVjVup6H3u7c5POPWbZ/gBwT7AAcSGtuuxjCPor4OcMhr8d/CVxGOD+
6+Q2+60DF7h0daIcKDQq8l9U/K27Jke2h1OTBdZg7Ng+A/BboLAkHc9c/JnlrUBZ8xHBNUslzX+D
qEIC3ZixVzZY4xj/tAhGBzs5eeXnZcq+XgVuQwLUQNuqhlRoFZHjqHEfIlc0kxkqjSlo/I7kLYox
IjNkHT6dhWOH/bHb/5YUbBD2lzp5tRaedv7+tXKfmwfWm32IB9Y1zyWyhRRfxUh7Jyk/SeizbXY3
+HVYqsy4Z5l+0nj1Z/XR/woDge58FZlaI8jEoIyHoEMUj3CwQexjw9JxsQhYR6R7T7g2Qhl+5JdW
oxtemtKOyvBK3OJYm8RpjgwhI8yIjFYKnzIoWzCye4hYRgXrOHkMHc8mtPqlBS+nHcWLBwxkntQV
Psvvf8RmW7NJ6aj2B314vWJfU497Wjj99I7Ul3XF4+l/5wSzy6ixiENHtIy/+jGXHBSdWx5l8bqt
+7kvunemOFMBnuAnjktp8w9j5g7IGxAPeVdAebEwDkpyYRRfB3e9UpsUJSmLR77pzmAQA6pWe6ju
6Koyg9ys7FpCG97ezW3M+FFmuFdjSIppbivz3UUylTFEq87Ipe8+f8ek2gF0OtaO2FhRdNTQ4xFS
e2jVTemtrsmHTSx3bH6mQdWxT9noZM9Oz/8gYqLBZPYdmOi90/0k2o10Pfl62+jG8/c0ioyhoxnE
6b+bkSi593wPE8ZYkFbqW7cSFz+T7C77M/V1pmokF7z3VIfNY4PQoZ9HhDwloRIWL4wnw+iawioD
7IIO8ss7OwPu2z8U6FHkXZHbgaGbhYwYBVpYMMAmZ9o0/9jHgDJGkwpjYEX77DwC/hVa/msEIyDN
FWq77D5eetaLzGX8TZ/r1Pp/LtKbR1aDX684xmI9FQalczxpBJ2EB4jtQZMRHHhAK17mPQ8GrMYq
uKHtxvRKq1jqtMwQIFrmCkpr5ED43iXOXU6cgoy+tlRI1+kwBxj3PFeC8bkdo9MKPaSyAGxFm10Q
GuSPwqmM821NMqfk8VHOeuOfOKdrQy4Jcl6HZeVC9OCFW0ZfbeowqiPkBTO20A1mTTDytAvH59fN
ipVl1UT+RRb+HaOgwGKdDtyfIz6FAZXAwvR98f0Tyk+I5RT7l/FoFnAOcJy3u15Lbu0X8x9TaN9C
Ygkkg5eCI0a/X6BFFADLgVDbRlbmGEJDb5UFwKnp2uOfl9EPnXbWk6+tRaLh+Bepc30NbpLiiv42
DJKCLLr9Hh721HXyc0N5rOpcBzodZb6CoIAzJM6SJKsG3DC1tJxjaAnrprShP+GLveI9nzMKZxQX
5Mp6KyJfMJlWtig+kbfQ7JOJj+emxt7xmlo/PARBNcTdebVCvoHDbrIR9re1x8Tlgy44ohrni6hj
0eVtRdAy6ZmmCUvO2UCJxQ5xJFFHt/L82Z+a13C83bS3aQ1FY/TpSwMMB0lS1wRiIz+ZxWA2BlP+
H+WhgyqxM1js99JdYbnkB/2ppap32DiUSr3sMeKhzWfnWGxVjLCMwy7m+GWZyENRxdIj2n9jvlJq
8smkTV7SdVIL3g6cEVSmmOLH932Y7DwxgBKGOD2c69gZy5111H/5rMTlXY8VnhsoITqTl6RDegb0
dT/vwET22Mx8/tukDgOAclQADh9NdJ0EZiXlSvZlRUQJ8KTJZkZU+iDivpdAeKxOrgZVQbQMAVC7
bpV4jNps+dJPcNUG46jKMRp8MACKdKDyASE9G1kgcH6GnpSs23P1ABS6ce+oqCCZbTzPfybNTpkK
/mLWC70vTSmqNo5Nz7l3gmE4n0BSj6IZTUODJlIwfhYA6JRzvyOvu7/n7avcWj0L6h9mM+NCTBkW
58+6gNkTcHtn6BrteJ/xtxjZn6YWuwdb6cEuq0/IXFjuDtCNYnfROdtc9RQyCF0J4GgfmrYwLJkr
UEEknlh183ffC7VJc6zzErYsGj94bXKQJUNyeVKRMf+bZPCXeElU+qqVtCavBlx9bpM6o0taMTHk
qI4uBqey0x5O0BsSDDLJlDTjc4gIClx00m5fqNft7ARIo0t16whxsWdmFjX01hAgcrTFM3cUokTX
/+ljV0vx4ayZiBN1Wh905rTGkEHhiBs62u/gJYqLTlSe9pAUW3T8l8HgWzAxgzGfCPykLJll8e4d
QDm/6+0TDQD1Igt0LgBzgc4I9VYyrm969yIA9mRO9hy52hOJH+Iydqh9VBFDEpazEgwJ45+Iabfy
7OJKmwuUxIWW7Dj51XGVAH3UTSVt3sQoNt0HgI7bwkFn1RR3t7Wx6uM+8B5TDBLPZANJL6eYqEoo
Jhp8caQXDwH/tXdc1Y7POUJFRVg8K5on/rKxz4XYOp4Nai/qz6caEYj3/EYiU3qijazkYZmRuKWb
LXHh0rULm9jGf3M0KbxJeNehS6bBufLVJlTSN5yiO/8VGyKJYTmlMS7N1LwIZxIs3Xq/XxAJHEmB
yjeI9A2RgDc2nEd0ZPPKRE4K8hKJXPfclg98Seoj78Wuiwpa5rpY62VYtJW2IchtmzXCdX1ftB5R
fUROVkSBdC98ZucEfkfeqiO2/1JxZL6SZq0vRb7/GDq0I5qGH7LgAcfGgdRsZR7VRcPcGJFvt9Ce
mVy7Bj8z9cJ4vCvFPMQp8LMx06QL+rcF5Si1eolYPuDxi7lHLa5RH/wH6Q0i4wBmIeJfBqXCnyOR
Ly2I4/Lb3JBs/dJSB2S1tSQdslsTOzn7hDfSZTUoqBsliyHSPeLwNwHhG3z2JppVQ5zsRGc3kKg1
rY8xhlayeZH6D6y9ObRHbEHp2tN95gsVdAClRFonf+83CviLSptbD5DCh/8znmuYuIfqVapRUH7p
cwqLuYR+DBwer5UWBmgIndf+MZFEULT3CgYhQ+rF4SwulklIotV9EvQ0jdXMlh+U6/o2zBzX9Vqu
qwtkMepveKr0M0ZqMoOBGCQB/taYnrhfVlDABtdffA//Scq0B2mObCjy67TjPd6m116wPljDg0FH
BgdRuhdDBWSDF5ETTM9mcG9RED1bYfWjGWXWK8et4dmA+0YPVotEbeloLTjKcXw7uHpS9JZL4iAa
nu4qb7thxhKCoqTMdTf1r+xiyYAbTJu/ieAdi+LSF1IOwq/0MkHuer3Gka8RvTGhLlQD59LcYEve
68tbMhnSyJihccw91SlvcX2AOKRYUSvF/UzzfMAmZGE/3ySDkehZuDe1YSvqo6Sv7fGuFreiHKgW
2VrXT1RgnI4Et5n3uG6yccErISeji1YgUJ0hvjIEtUctIyNurL7M4clWmghUqi2H+649d+FjKi5o
ITX8HekdyCZ0gh6VVxPJXzaOurs7L2mu59wE0hATo//6hvMwN16/tsQ5yFEheUhOWlb51lmCV2HN
CDFyiUWj04gxtAkQoop3lmh/hWjbHO7oh1L6zA647xTxcwx7se+8bPkPm25SLeqjP0w2OIJFC3e5
QfplKICfsO29irr/2ST8mM8DvfD4Nj6mEoESh8H4sNvBaGltyVhcpLMei97gqP8rHv3zz4qGszw3
0XjLmxjkC6X9V8zW6UJakDpeCY/6OA1QeR0HfKdrbN2QstXCxVPivAUuc7nXGMQVjgX+6Xp2Z5hz
AL03hE//cAUwX/I20yyWA2CseqbieTp0MP+5Y2Y7H/x9PoF/aqcWNEDSvtmt9PMcKFPtLLDV7ZpH
DDyyq+UE2tLSL5zAW8o0zzOBB+9LlTpdjLa+fvbZX/H5w1sGkbOupLtt6GUp99nBvntnpczNKBQ/
u+5IvQRvOh3L1dPH/n8VlFqMpFZqUuKliAJ/yKpk2JAXUb4Ds2xoqYYrFq0gyZi/fEWLa4lIO06b
B1izQIVsvM0hOkMokc/ft94Du+r1K9l1k1j2Vlhd27GFYdQYcCrrfeyf2qmy20f+0PrJANIUfBOO
ahkcCDw2r14zO5dD/9Mms5OkCmFYV9L8Nimy5r+kodXBqJo6TgQ839FM4no977M5S0IIu7wO1rUZ
pVJsFjWOQjve46m+x9EbxJUrVeBMRdjTMjLfMfL5+S//g0OT4Lc/Od3SazhkBb6Ow8oqtUjOlX9l
ozBwaABG76CRQU7zne83dN5MnOEl9wZAb5BavTR85g9x5/iNYWYVODCDcR9UO8HOpoajbSxdZKyN
GK13hTvfsMWrsYsWOOG7+p1438J6k7MyuAMBnHrQq9reS70TA+AsrDx0vsbTOsaHNAVoXw0W7sXv
FD5yuBtXr0kC3N74hzJQS8zOzSzqPHY8JNSsaPjc0zhea1JpYu7vACUyyOqTtS7fr2czi98rOUEv
PQDerE66ph7vfWKbOWKPlTTEoPs8xnPnMJ4wJQ5KQrTCxS72KJjdu5srNnDzws8J8bZUXTZV7g5z
96acwqstQe1hQSnwg9XF2pytYWN9wJbdaBuqqgogZ8h3Giwlb0n7lo01pGNzdk1Xd+FkbqTH9onL
gK+goNaV02HKxcxD4Rdvxs7ylJVqhCMXhxIQv5d+0jffeytHDH21NbeFN296AlfPo+z+C9jC+oDe
ClKXic8VBh+h1wWrtqKBjP+6rNEzlfeOGpivlWdB5rX/KXaI1KDYMKQ4n+BENgRIXd2F73Yhqd3N
S7S1JxNXXj7I/PwkMAotZ1FVjnzIrmZ0Te09gR9oEP1xHlD8cNkiYOYHWO9Eql2JkvkLZgGrR+/c
wnU1XV3WBJX/ooQyWKIjG490VObYwAjitRyT5VBgr4AtLayOyuisp4Kn9nfTO/lQjbFzM+4OJU8S
d/sRA0ZjaNlx2utXNOhKRPP5YsSGPQyrRdeMVkAcoYLtq9vb6JZLy+CKEhvtcTE25tEZ0d6lzAr2
Z3mPa2x5qxgNuTN6y8Xtg7PNbdNXvmkUy3o0aSV/H1WPOvIbWl4V+JGAwA65bbom3Ag/+hQ29z9e
1h6cnYwnzMwqqmzhTC40LAWAMx0Q33vc1tgAHGVlFBMPuql3RQq9NksFylZquvyE5Gz+Ge3XOQgb
MVFqQYQAItr+cQn2iFa7kdbYzt6MEG0lQUfTM/cGXVSXgpQXvLeXajbjLYImMH1fDFYUTwvPowX9
EvtFsPYek3EAca+s0LvOcGOwJ1j/MRzyOeNHh62JSUiNdxCxxDYTFQbnbecwHsEcEexHW9deuF81
pQDo1crcx3lkXJkth6QoVh543jBJUA/AiRn8r2HvfebfkBudfs3e4UT3Ff27nCsVKCTbrPDgnuOw
V1s7UYP52HzvD1Xy2/AiouEXZllBzWHprKhgnhIdkOnDJ3dq/lcWXCvIoBwbggt2eNSkt3ykH45y
fH2Lt7989pdqUiVsVAVwPCXeEjP0nc0xDjq6/Vpbd14atCkshPp5idhaAwxj50t0XbEaN7Cv+bA7
UDW86TfuZ02PEhfaMlJghHiByH6JTQLyrLx9lJvzK9CgXLiCfSMI6xYVquapA2n2aF2AoDAbk4rA
t18SQn8xYMyUtkXXnsP0ixvwY0XzlV1VtGlggWM5ombSeFLmVv7k42wlHjgsILXCgttN+zPCpenA
nWyPgr0PCbFMB3/G9VJXphPJDr+BjnlhJp0I1CtOpilRX1m7Mx27O/iAPYCsQiCqqVRZMGns5kus
tIudKwbnyzgApSrWWJdyhXSAKmA4yxrzr1dEG7r8NBZEjin94d4ntkXujFszs3i342MHWykZJLj8
brWjmdP9YslJjiX4/IJWygS1jivSAmEuIQzy0v3Bn26cXNRLO50pJF+VHOJ3Hggpje8DMXadf3O9
lfejA81lVgu7n3cnW29Fa/0NYEeVrM+TP5321ERVJgTF2FqJvqv+MF2KpReT5I/2uGpyHAzw5Gk4
tYuHmt1H1/dUGeLBYPfeelV3cr11LFd50FfStqddU+9ls6sewjmoJ4AOL4/1jvW/jJiUMrnTxyrY
Bf6PFTxX9h04VW4j+yw8ue9YgQLNi8Fzx6kpoup+kRQIb2UsKKUkFsRQ+VkwPfIndCPxopf+s5to
Cw1D+ubPOPWP0Yt1loM6L32U7MaO7mYGFL9N500fzbMiutCi0ukJPVflwOMhlJEAPNF49DXZGwl7
Tt2JOsN0P96u7nC8lC8SzEi+FDkVyMYSyaQVtpV9RJrGEjLtCoVuD8hfaVdERl754Xw5qvVsnMgJ
mTussRqbS98Rul1gjfGd856H+dBQTIWPpVPX1HMQ9VIPJgZOhvwRUymoOMMDNIYZk0SrdvWJQSFj
t/S3LFCUNaLp2vkPsMGHYbUerdmuwxq6CYbvoiFCJxuB3TcMRtDdz9IfZS56iyAveCRPEhVWXsYR
pZF2Jz/nuxvkiK9DF5GLjWcP9oppeFMY8m99crEzjVqRRnCzREK0y+874hwxia687Tl76a2Qv1zm
N2lEMLQhCxKFfoNBZQkC3CzoprKfGRAbVOAOw4tOuxtVkGqN6/Xx6LEIPKUfc8Ep4iP57Of3u15x
IZ+wuaOBSYKJ6KzhZcTdPDWlFKyTP2tPF3mZuz3rIwuzmW6zsv0whTForJX4OHj5pXWbIfmSvVR7
nAZJqmM4hS9dyDShCHmCFpR8Bd3iPXoChTwEfnIGGy5+/ita54yHJRp4xNctwJvMIJmDUvIfcq88
zj2klNN4q1a34EqlVfOELDOdzwaIhNfWADoF9Vw6xYRASqy71t8iHlbwsgMYTduOODVgtQP1u+h5
Kr/mXkYxjza+ATzDdNhcvcrfMU6LiAROu7M4tBWF9iTLOk4Mx362ilsi4eIx7DlrqAYa8nm81rLI
EozmIvIHSsUgiKCJeDA883h4nqr3ES14XfTtmNy3CENQfr4PMvWgIE/eYxWxHr58oquln/msQETa
dh3XaXXQRncpO8iOPpiMzY1Bz27bORcWyBBhT/PQ4otBD0Ly7Uje6gcJBVlqthZwxrmKG87Qocj9
NzYT4AbSzjqiSAqUhOub7ZgeTJbUtn9uDntLXfJrnI23vEuUM5ZD1iquZr5d4DbkEApdxtwDn2z7
p4MDAXvGZN0/tr8t2JI6m12UqFjL1NVzWeam8G1baH3XrHxVbmABc5VqtNzgxtzn3wnV+yJsiclj
BY8UIV8HPqWxWpejAv7BwZdSsoq0KNKh6Hwqh33FG1KIA0DGQ01VDne/kmHgDCrU+4upHLxUP+4e
0bm6irGilA4fBm50IPJOF5HEaZ/CHUi4mzLDhh4dJkDimpHjxLjiRLSxkpCdh354x0yAflHAtPu4
EZOpZdXGhQtox92X9FZpUx728AvzcK6uAugK4AxR3KT4CmvDLwCWx/2UXUengI7HVqrfFi4VOwoW
uXHNcZSu8qCOtXGf93FlVW0Mun41LpzIpKXEOeBEJ1tC5VTeymZOMjjxM3Z1t5EwY+MPKj7hbVSr
GDGqBdabtbE2jEpySAHa+3HzVjqzb/o8CUhBAZgZyXhlO3ZoEFzZM4d2Y8JyxH7x5rBA70tl5av7
rR/5Yh7LNLkVPSYHIDfV8m/nh/g07Mz3mnHZfG6qhyfmSsM4p5JVKvjZ/oA78Tn9kazmH7mEeoIP
SgbZdU5oULEzGRQ/LrTBly/rjOhVNbJOh7jxU7Wgjw9+ciPq7iGXgsf/aK5QXmVpWSl2b4xGbND2
1dSUXpJ3Q9wdF96AVKx8/0pMTWbzN7GFJ+TUyf1R9oXzHZW5pHnYCQSPlDHTW4qbZuJYvfsXR22f
IT9DdX5KnBlKAGojYWSIl48EmR7tGQH3KcqoOnFWfaKukd6jQy/I7EsTSOCHaXHOtd0TEi8CO57D
udIYKHH/qBXmoGglBt7iUgia/0QyBj/sI5/KjRG1DRypvbgSm8jvuBNGvTEUJ40DH2E5ZTq+qg+o
QwmI7aHFiLDc2TPcgVFYs46LPXn7HN7IRp/iT4Fe/tJa5SmGrHIZRS0v3oAsiqatMXOcgggB0rZo
1LJiII498NCBFO5+Rd162pYfVLo0DITbRIxxZmc66VD0E10jWWR2lVwKDAbec6agC617E1IMhaU7
EPNVKKZbL62PKgLaRgKnH/moPLmlz/eSHKuHVNhrKMporKV9mFfEFTsQkp2W6ekYPj7BKk004KwQ
Uw74LL4jQLf89eQzJyS3iM7CMFSgLcWbflsDeA1ikpjokhds6znjc2D+9WC4r7xltGcToP4JT/SL
VzOjrSg+pGFzGFHeE7frUCvGU785IIiZLo+q8sm1P/sScxdcQJvFdUPq1EOQEYL5hC7yKWe87JUg
yW3C2OBe+8KLl7Vs8NgEEIB6xRxn9qZLDe6Yjp3bM67ONymkPzLAYeMQdK0doxr2akr79zQZMqm3
/dsPme8JMPArrSF2mCLi5LVfCvaJ/sES0/9p7/EysZTpQsYM4iP99o78iLsAmwKN1cCyvrs+kXHn
KsjMFD5FD4fEZwxPhsE6dFn9qdF5GjHmbdYDG3ZPYeGgwqSeIzLA3G3ov/TOxlBT0RrPRfQwKiVY
Ky2ozqrEk3sqkwJriCSoiEs7OImMGCS9d5F9y8h+0x3UUXNa4WVFSQdwRvePpGVw3cpL8C+6s7nl
UXiagOwidDPuHldTInTySab57Sdpqz9wcOGgVL1gtHQWzydS+8O8K0UPS4RI0LSEXu4Py543n9jt
7ZhfcScko6Rqh9BENze/qLeaC/1kQiz1LFKG6DNjQYl5cjX/zYQGNSfUbCkolFG7AsqZ2tX4iOEt
F2ixkIAxnYROt6nCIEg2Wsx1iYClmAz9rVnS/CWnqyarGtL4R6sXaQz7BFQaeA0eOjiqBJniYMRn
xUzZ9QsQY7Rd1H4YPPRcc+OYd0k7+LHCXU+leIVjRaVf1bfQem+IIVCE90CKxDfqqoXf2yenlMxA
JUG+vKPOO+D1d0Jv4rKILs4GM7Iopr+w/SnERRuelFbY0Sg0Rj13xOCuIFLIf7pj88NNwoebtsAn
KkIJBvGa+KR9HmS1pZHPpWsy74n7R6rUYHjD7DZrvYtfsonAvz11StCrhEo8r4fSVpjpWDDYX/No
fSbbdVUglA7/jmt6JFH0Zr4Qbnd0zJJyVQMfp2F4EIXJKPst019A1GHXiIr2EwSBojVW6FcJc3LJ
l8Qb0kU/a3Ma86UcqBhuR9jVQWA2N5Mg2eOFlC7MWMfQkSFEZRZNgvOh2fcnWHNFHhi2K7f5uYd+
SDd0tYsBnz6slktYWZyZhWP7UJ7XJSRRou3HXTrweKNA19K8WpaLokxOrMun8c2sJs1R08PW7sgM
ZWWXOCLdtEFYIgOVhndBN5sNinw4meAttv+3vjjTs6aUcSmbQ6IWTFk0DCGkzVI5oRAY2YYk4SP+
Z1RpXxVSnwxsuQYroMJOs2IrcJCM3DSKJBPY7a3rJouIBCybX/XrjeRN+7cGMX2CdMIrhB9CHwL8
Yj0695IxUQchzFVIQPj+sb0ZhV3XH2Me/uHh0cf2KKdd1ocxZJUilVakDdvuQNuJ5uC0rMyGjGKb
oPVGnqZdlKRJ+B/Lm0mYvXzrIRy8LhTAeN5VxkunvAdEsbdWvYQDyuxF3O1FuzLjpSo87RrUNHc3
2REZ+4YYIC2L/qX0tJJXsSMrXiGY+Zux1RauXVitnAhG7FB2NPXPwLRxFB8RbtA15FtV1r/sS6/1
RHYFRjA2e3rdATWCxnkxJaF42v/C9xnU+WTsrk1uLUuYCpGqH1iVyp1fHY/ufNyt6+K3nrulSglL
gL7pA7d/R5KjXvmD/iMCI7cF7y+x2C3XcVyk5VCGzxRXuNqM/Kxri3W585X9IZMxzTP5H98solfO
0OvUnA96Q/mZhvvAPSOyu+tAOhRYRMFEoshOthBC5t39nu1PsItUolg9u7YQvnZHsoarzJLaXXpA
AG6d6UPLbZnyQV6JgXlMT9f8KsUi1Ma0G6p4qvt74J4Vv9rB9UeicpESD9jDQxNNjtPDjZFzMr7F
L2vKQfDa+tjXvCGTX4ehgJB3eY1V9KW0b4p+l0ZLmB1ZepIVoEYyaIqqqKC5yMyp228930Kxz6iY
PeLds23vHIppXJGoI0rhh9u5fztal5/DpWTWsP7OcZImL7LTbhIGlRLZ9xHEgkfAZVNY7NOYEggy
jhActCA2AL3ok1PfDpF0RBRDSidsQB00MyF7zjGzU3wtT+bjJml4B3zAumIQjpWLfIPdxbF7qxTj
aQ+GMt4OicDlzM7w85oKp+lAEu51ozvlQ9Xq2dBLEaIhlOZ5xvb00eVesla8MG7KwHkH+7QR9eC0
2FbjEwcA4ypcgIA2cVckcMqSuC5iz8vGQEciaDGQya6fSQf3uGVcCCTWsbnEuP17SzH9l3t4QR5j
slnSFbGZQePueHE8nXwLX7JYbjz59bg9IIGB7PiErzL0C2fiToDrbIZ+3fIaRz0Ee65wDsu5X15A
aAs9PY5DZTuUotgewm3Uv14yBeYNMCVg09xajHpMa3XiKCi8U4ZgolLBSkfdEuVMQnbUQlx370QT
t1SueDkP+zf4PhK02SDe+JWAcS2vcTc9wWt2QpCbfYC/xqI19wj4fIe9wgxLW118DJm6p20jJl8d
YAHu57/m4FJtjYQSHKnM0ewtzSjcPoH2o/XbKWl08eqA6wDDr8Ru5vUiw6sj49V9gAZlYlUKXc/h
m+JaSAklpC1w5q+05j1vfEhbSjHpaPukfJp2k7zamhis4jldFyP7nRE4xhD5gfra7y2xb0ktIuh/
ozthu+d6liGgNWSsgSDDUlhOHUURAiuup3ma2HsOdyRx6lVb7sTR8ElTdJoZfiNLQm8RDPnYpHqY
MVxYCc5W/dxrvVsrHCLcg8F2BEak1GPaJJKj/pSk6y3PAU2eZ6NMc/y6Q5qp8jE+dZQzkPBtEWJe
UbCq3WG4h/1grvxtyTtOzP9rvM0fpy93z6XEEi5eFSsHGwiHwEfIxXg8R9vZl9rzgItuozobhWGq
LmEB/8IiiS1Cop9gNsgQK0deVJ29Z0HtW4q3tRksVXYQYnYvTpFwg7p++h5+LCqNQZDbVqg0EWNW
xDrQFcqoWGi6kd1osAtUQRVMBZYjzAI+9Ku8HtSI8kRZX5zNohR7BpPczlvjJ9W3zISDapzU0iJI
qN2NtgrxMPBsL7HaZxVBZeVx57oB28XPi5yxzorWhylyweu33lBg7j1muQHHUHG3nJxhNdLrUD+u
nAZSw0JT+K8J1YDqdABVxjJNtzN/CzGPpfDiJR2pDA5k7EXT1E61hdNm820m2P6bZSBVtFL+Vq6S
Br9WDmBZPGsWCJQ/guB4uZKm7v85bFk2Us/S7a+2ZLhllCzJTpNJ56LThm5aetP1c3mXbPe906TO
IcNgOdOOjIMUTN+4T72smbftmIccI5E4MLOUxYwRqVlGrrBR78rRoQ3QyqvsQL/gvHieq3ikobUG
p8BbiqEya67qxe8R6U9iDFgtCjQIzMD+3gNEX+BaKiB+D7aspD/fa/qaCy056HriV4OsoXLctHyj
0PRH8Pk60mTsPUSDmOUWkj1MjPyRHUTfVGm1h5YCfE0/7m5+MW0Sx4dh2hFwqCosR7q7d1GfJ0Nq
nfGTMDrgmh24zwqDMHbpa+EZS5Vsxkghurh23TBpTUMvWs+e+XrurYnnkeDcyF1dKYigyjJng+FL
r9IdDznmW6DqjEnVWhEW5ywMqFOvVIkVgHq+TFegXx9cRnSWgf9wLGBtFJ+jJtfI0n+UIwsmN0cw
RhIZw8x0TZ36wVUVApyDMOOHhxtn0RD5XG5pSNOR2bQ/5a+vW1OnkI6Cnv82QAgjmSYkowWDV+Nn
sCYHk6gbhigBr9jXUcPbl+RrYDqW4MAoZx+dh24BD34dvB4rRjl85DVTBa/tvzMkFDZpsx5Ehvus
apm5jcV2WS9zXyKqmgQfFteLk+57e35I9bpYEMUV66QUtQtRlrdVmKAA1vbsK70obFWDBt1dVCSr
Uj0O0PzQecoq8HJBxfWjRviDhvlEbc05g7ZX8ZBmKgSS4Q1gwQBhHRptjB8g8jtZ2KAmVVH9Dny0
9cTstBACmDJveUi27XjntUnXsSl9Q88g23Sg703jw7M1IDE0qhUpmeJgXAj+kCDl387czCKK0L2h
GQMzm9eSSEujossC3Wy0xt1N8BqmdEtHshfPvsFMMtoi++ckQ+k2MxvnenGOhxxS7E5tgNX8pgUy
yjcNz6UlPxFBhbaG7vns1rwjLPce4FPfquV6IAhd4hwND62FSTUlwX6R+tOgCxrT6nPM4aFPiHBd
gOtbfkrcg2v12RLzPoB6d47oB5N2EVuAdwmOq5Vv2NKahKzhfIgEB9H4tFKjBlp2PpxO0leNvov2
kRPX+spwxK9JBIdMzC3Y1AglUJwSzxIP2p2nHWAS3PY9oqrwfEJ0inkpo0zS4Xa7nDMIxtBUuXTW
OdwIODbsp1Kip96tnt6Un+fCzEOj/YGm5eFd7yfZwCzbBl+LKhYA5eztBLyf5IxmazYhLJ1aQqNa
6dDI/WiuuUVNPcyNuRDOm0bkTX8eHkKsT5klakqLTQJ5APb5vJ2EuirFllTTRAUcBlnmvSvspSJN
NSxc62PBia17Ei0zXGghl0tdXPHOHvg95zdQZudThWl9eo4iwZ/9ZtDlB2u3yrgjpemR8Rca7qiY
zHBKM4SnQAuOXeKf7NAWBwZ4l1BQUypcSxQ8rwPFRbUhxX3OjYtDiGEtMW5g9DjPi7uK1KtucrXu
Pp6qZ6SZvNBbBaecg49xDvf0AKpwwhWtwclpmvf7Z0wy+wp8rdrVSXCXvYdTMqoMk3VKXMkEM8jo
uJq4ewRIEhVsU9IdG3gz5u70mclT6cxFI84o0kJbPTTEQhcV3PC0rFbpvctGpH/5CcmySNgamxGy
klfFD87kOWoIzQeYLrvfu3rPPD/lO3BacDzVC66gFseCn8ypIwF+Wz3OGIsCu/x7XXTfQdeZG+xo
pyaLvf5o0Xz0cjtWeR3Dx59tQhaBSJrvl32K8K+qIJ05WNHw3p/HDQ1lRhDbCgJzCcdTh6poGxaX
X58XrV0yBDgesir0wAuvVUmuSk6cxT7lLS3SfZB5VUqmcRfkrfhn5FowzmB6FV5/0KDhaYPTjQyy
xNXmEeAbTkWY8BSVWkadnXdIqXbCHWSkt77LUny6DaUebEZBqM7xb40YnRajZLNzx4zHHzAo/IdU
8MVu+diJcJL1W/S+Wx8sMpMGpK2bjnEeRXjkz4EPcxuRRhfzOkw1cBqcyPgzhpfPHZOwhdnH6xbS
QktDv6PlPNoaUTlU3sDAfq+ALeYNGli/Do6fX136Y+4m9RjroK2/aC1dsrWZNyV6ZOpRkyvZR4Ok
ulw01h0S3Tz3Tx2Jb70kxjk2A/DyT3ZRmMd36vJYf+SnZvEnSeUyxxe9d/V9lmx/qzUGUX/VBhLN
jlEk3qgKO/NDLucmknCDQMCD66rJtH6LBzfvxE4+W+9vkVCEi6yTvcdXv5bsNllnF2O4ni7k5dqz
XsDftgrkHL0krdLheZTI2vOPoW5rOo2cf4ti7uTCsEszYvKgFbfuAWRVQtf5u6UByMSylSAsj5hM
aYkPihK+dT/nlNUOiQbcSe4RyGdjBC/9zC+XB/DaSnVfI+EpS6y0EEbAqlgg4m3kJssEbvfMIB76
/1kHzXNPi2alCUwb34MhtqlJP97a+rICk0pGuVLpKx6/JXDJoaqD88mam6tCyo8UU8FfFcqB+IM6
xVXNqud4hA7uDs9cK47hBOl1aOpvswJVE8bUkVFJcREn30+Z5dI4gtr07Yu85DAN+YD9BjgmYBLp
M6Sdmvv7LAZaZ7t8j1nFxwZqSz4An7ahwPU/xBvd8NxEafHVkgCAbh+8tEidotu1/ndejeNbyhdh
CvvEyW/MxbWoZIFhBKv8wLNry34X2IgcbVNIC/QPgLJi7ly0jyOV/O0PCwM3nG7bgWCGuCNcuzD6
G2t4tDhujATg75zZ5T6IrzDHixfMXIcjZXetQCunwNXCoE0stm/Yuuplvsspae13DpiS4ZCQCrE3
+Zuj6zA7TdBuddG4v/AKTcy2VuDGEr1hL+TsAAsR45zuoNSZwD7FSj+MnSiIR0o3rjblcWb++SeY
f7d09ifX8PL9LA+TWbmG7FSfnIIuuTHux2poLyLSTq5rh9ph0KhWGN9mX5D1IdKjZTUql8T7VCAK
R2DoIXvMIUT2y0cMPxJB7BjdFKUFVunRgcGwhdDFbjGXgwkiIIM4a8d5/jF8BTBMqyqfInvTTn8P
lXtPJUUuHMqupGFbDar8JNtKgG+VwK+IE85ppIhBSYBtUERD8tM9MO29udA1rQrJ6EpIm6BeYq08
OEn3lTpbLalH1g4HvEbdvpliXAkc2Yv9rQ1DsZQxmcrAomhu2AVBx1EDv1N1jhUsMa+xZDown4EK
gTenAaOIQ4zgKQS0a8hbPF0Uatu/11lUgo7XgrVTRiWFr0zfJzY0y+tDV0YxrOcPfblPuCIkyguE
byUvm4bPDYh9fRFb+NxHGmeOdJ35QObaxSIKOhuHcipUvxuNetwkSTcKB9jMv2e073KnigePQoeu
suF2aySIuTWFYifecDEJz4NIHjMqAz1QqIAT6++B/cgXnbv6zEDjxVwGc/snr4fglyyoR2mqlivr
l0d1O9qKbffoo3LXiJ/GIfhbNfHbCupbZqpTUQijIgHvzDwAalfuJQF+UvhLFwqzu36Jo0hL5cMJ
UdYORK7GaynVVnKYSvMvrOh61XOy+7cQE9I4EBFRRCfaHeGNEOlZJk6OyajAROakEXlyeurvURxU
6PyFfovUSIKERtF1oE3SHmuOX4WgabTK3O+iMel7Gf+kIIEiUDJXdOv/go1+opmqOKtfpWgAKEMl
4/PhICOo0+aKv8XUunuyf7k4kb8FJ/2M0rSqohFxfIDp93dtTQ3WyzJwK6DgnTZe/buCjOkurrdS
AeJ/Jl6LSOimcU6f2nNmphknqrecg5MZSOem3jnb97yVerzKJoJhF7X8Xw12z1JRaXJUkoxN3JbN
YRkbYbr5FQn3okC5Xqy3Gl/rfNHuRtS4kSybEqYmHykJu6VQot4B8xnvDVhYzWzxFlXK31HVW3n4
NE+4elAyuMpqnRGM9Lk8Lw9tygXw/mETFOdHsAWmKBRj2IP8EX4E/2otJfudMqd5tgB8bi+xV2R9
KqvttKcRL1PkhT0P2CGD+TTmq4oMT+hfFHX4UP4/4wybj8KHQ9frrWhW8gyOkzU9DXRyzbhuQCHz
+fKZdJSv2AgdwMaBR2MVNefOI3zsKj5Hoeg3MUiHjoAuQY7B6VvJaVIvPJg1/D5MdomjHa6T0AM8
D0REQdhM7QGrNIbkFlSwuYB/jjbYPCjaZJDkJXAgu+ypJno6MYIvDqYnqKoFkIBMjweOc5uj1/XP
I5Ral7iPp4m7JehzA9uqe2k1hkw6dJSyhDK2DnW5BI28qkv0DEiCtMruJbQ2y/CxLks0acVIc55h
deY69YliHUxWCHJ6/XtRQ6A30D3bj0E2WUEjkXUce0JiOkZ1cNbprW13EukbqwQpzNPTj+WLq9UP
IIH+wdZGRM75wDVUK2KL3NBu/j/Ey6ICeldeQYkO87I9T6YPHFDeS+dXvd3iz0NtJeXwC2mV7H0q
h4jwralLyP1XBV570oMwohNxOIM2JXDORdptt6XzTJg8aF0vatIYdvo6jUFIwFu964u7ayg0HmmA
27PwsE88vIXLkm0zPAIaDNL/h7IIhfhz+kBXhkBtQrMbM3EC7IsdBLHjgfhI3d8scJ5pp3cx0zYD
W1GV0OtVCjCPEoHMRZspjFeAFv0WYEWMNxIJra6qlkg0WK77L14OjNU/I12gcdtEhbYHqAuCBrI+
xK1UvDob3dWWLBDd8w2TjSOOgh4aNlZrlVVmxk/BzCgrXOJwV4yG1fHNexMHdSkwJykSMuJx18lQ
OLSz5Rg9LNrZAp7QrWabo3Xcax0KUJFKjInIhUVr+NSzkwKww0DWQM0QVMrQp2FCYVV3BiwIgB0N
vWctQSmBvCsxXeIk2ZOhUlEmlm+ajKVjPSPNMAUj3sbwTUHzIQ0q2i41x+wLPbAp/5ALsf27+iTO
gZuMtB5vVEXbRiJav1ajO5VpfVI2WYFBlkyU+V+Wq/7uzexIvxlamvrjNd2GL/SI+H2mNxBE8zb2
Z0VRyzfPWnue2c7c66YJ1iJsDMd6jPaNQLn4Okir2LfC+WL0R5c3B2tUL8lEppyJPtxIGgCVETvh
zHcvneMiMKmw8pDYE79CJ0/YavvIe70bhWNFxTtCw2Lbj6ESCV+JFt56FJMkaGXpRgdozqcHhfFF
8eXBfKUExqjXvghiXpuwnLyGM11iSk8Hm07t/BLnSoEZTDnSe1Inv12PRbCzXyGwNc7bSyX95a0w
PWWfCMI/QMt2MyMdHTlUDiD6I+25UHaf+CUREzccIC5w8arB1nH0NCJEtXONw5t28YJedTPdrvrq
bzxVCVw0NWTJUlFDzgIgMbJuguz6jv0eFzmJJiDDuXNceaERVuN0fmHhuWHPEPmylFlm+nDRvia9
KkQ/HIoRHbAyYQkD0mPbWhX8bcayKp5H4yy3rAmjwMRR6QiAavmGKnR9+OQjH3hfd2WZLzYbOGCQ
A39XDmsZT8yPsbf2aD31tordZRIG3MXMLRpSUCXzuhdpWW7v01+qNay9SuBf0Ri7UvXLvb8NUXTn
WFOMbUqGQsYDIpoNYko722/gNltRbES652rQmlcfqXAqrxN2yKx40BO/3PvJ1M7sSiIwB2xj65H4
nxxZa1BXJCuu3UAF4WwiM44cmDUwQRgWJiNXUNRb5ghtHdg3BxxbRaG7bQCS8YRYaJQnldNSSdUW
V3tTrX1foVB+ZBryq+HWBSL3cQVSemMlQiICazJ/iy7e9zmX8VJZ82/lqLmYyLPrioMkCLaDmw+J
CPZqpLQBJAp0Bk88ZOWxPyLXtVJJda14PA237H7/PakTwBHr6ec1i7xPN2Vz8vRlVHI3w/l4PXhv
ajbYmnOuLq1O+/zXSBzBZZQTo+rxXReKEYSewpL1WkIyuJgNVujv15dFrF/fb3KTuPWzq+WLgC17
nTZo7Pu4KHzmc6jCFDfOV05f0QiPZBu/yxwEiR0F4GOAGuOFaDWjvMuBGyPC4brQ3vv3WxxeDNDb
CFUWbAbnDnA3FmF8cNAJ4zmcnGJemiz1xthpwCFutRzWThXTkTkhUwJC0FVa+nNumrXCZaR1g8i8
o7NhZ1PiVT2sMXh6eagB+RFuwSMYb+4fkST5i7/7lSYumgda87CozdUqP7qaItJw7M3EJPPTsXyu
HMzl8Jx7eswNjX8fSBb9kqo9S1A6MbTjhjW+7VHkjF0GbuaMQviCdj4RnGG5OhG/yydzBzoqbmtp
zkL2fAw0N1f9XIfDdqdqHVdlEfKeqr8wY5RYlrmIzzYabCVJW1CtKgnuP1T6KPkU/WmZsKowB40X
yfOrK64jkhVqEWLLBrcHkYpUbGvAVEPBuWmicuubcg9P1eYdGhTgQCFdxPA5GLwgCz9iiZejddmg
IFHruN86MCJNrYi2ygMAmLqavLDjpeFw4YfoPrIdAEX3UQn5QsvtxTtp9/3XdFEztkDYMzahtFmr
WGD5Htl7LqfGXItXx9YhvjKkTh2qvIZsoXmyPrWkLBWM/0h85yuFv1RLxLHVyUs0O6snQ3nDSBvj
mfte8AbqLFxVrIv75AYwLHEhlLAJSPh66+FhxbaXTsPh9usnEnnSa051EXZYHk4jhLrkyTPqOhxr
+6KifAX2pjmdV42FAUZRCzgN6cTT/dYfKrgwn3dz+iCyglZWO5XzGfPeTqMM54HbVrLquqPK0T67
oFebYYMC6Kk9B074epfTB3Osch4Ix4MAIMnHQ+yw2YQncuyOFdF5PxzjJ7VsSa2CW9x5Ipk8N+KG
NTNCz6kr4Cu3O/cUlaEVK3vdcbiI3yUIKqwDI1Zl++zRvF9+9rysyRY8Oiztcym7hs8rLBSi03zz
2MvkQEUiAsF26Mta6A627aJsgMAyv6vlu8/uVRuZOIce1bta875P79yYQzB1zRvvVg4XCx0boX0+
XyCWPJjrF6hZdn9MFhCbsn2iHy+k/q/YWnG5nhEgHR8OiCY2Lzn9qMdTNK74miuOi8I606m/g67g
JX9aBPQPetSmQ3mzGiw0L5yui+uUs9JLYXX5wOWeGeuTtQA/JTl0dZHLqvIvlzBB+lVJg5+Ddga4
iOgAeQdHzqVDP/xha/TsZKA2wnX/ym7b8pRojcuMaE2QaSj6iBCYQVAXZI7vN8CYH1umqqHvyjeg
zl0PdEX+ljH1Xth9pAIOXxe+OC3XX9kS/z4l1MU1x4wpn9uNAcAw7qD5RWdNTbbkvLzAkVU6mnRy
aVNvvg/z7kYQCKlHh5lni2itv8+g0SeC1HoIh0p91rRN+FYoTLI4TH1OmucWWkAMGuQIibbQZcF7
Jib22WgYWIek5zjQhFp8CZFChjeoKcsB/jC5aoA0d7K+gQF/p+xidEzpYm6zptq2htnu7xBk5JGK
akk7OTe954stMcuV1AtggYHZb+q2jyFYaZfIaMayL5m+Fr7CctmEduM45ovUvWeAuyBI6PSrMMNz
SKqjFOG3SUQJDZow19gh6HMaYoQRSLNzdfEohlPIaNiDhiFjaVhRAi29BHwy02U7L4T/t39CtsAl
VPUbIUjbQh4ON+8eXP5sJES4qZ+rpnO9SEq/nnOyvRkM8iQfHPau/I8U2IpgQtynlCUxrA9Lvdnn
g5NGbs+4Bkr2hWnYGgC9HyNpMgPFVR4NuDOgSrnPSHZKYWzQCvJrrAuTZIhwrIm0YB++vUpmS4cr
bWTC2vi3uZX6PEYQjA70Lw1iVAC2K1qskOc4dMaHdPL5P/0vBM4mtP4X1q9fx4KHz70FCOVm7l8q
9O2m2fuogj5G5IRZCZPXlCUMgyaEIuBJ1iY+JT+RGcpiVcp8NsPdmarlcRfAS9i5BN0E9PfGRzWr
SFq1px3vsj39/TOwiFLdOvPIQZws3d8EWRnbIH4zY+IlW8W9200R+oeuYxpF73RGSihWX9K9SjBo
+972lzJk1RHYeTEaASIBpvtOVekjd2db/DJxBh023RYrjvOEgAtaHrYw6yx6Pn9arH+UsHaL8E/R
cXYVQSpBUChk+ocJfzzntTzyuDmmBfnAU5h5F6ktC8U2hIJqQ5HWriBOBgwnRDXF9eZdmBoA4eOx
qFlTcZcFUbSRreew7182zQRtQ7YmHpjCXFEms8kXeOaF7oinBV3psZHcMHdZSgmJtxE+Q9e2uCwr
QeaIF1eaTfMqU2NWEtOkIPvP8w1xzgH7dt6580G11Fe1D0gtYwHgd5j8ZOaLjLKPGBW3lDKagY6+
ZMFJosl4A0RT2ML9PboDOeoGdAbPeOt8jG3NDGVnCnQWB5XNhjnzlAXUPzgYaBN4fKhgS1LvvuDU
f6Xtix/9zx7JHgUwi68FRrlmvMb1zr+eLVTLl5btf6ugmfjbzApsToMlN23EUnEwHvYClM61jd+W
8mQv3mcGI1RQcUdeVbcf2ngzeupSnNcCaYHXs4NP18x7aHgDdCzpjZvClbtTh+RAORS+wKYQ68bV
EDo57hYZkje0nuhe6spFJTAZM7NxmzYIVQ5g6el5I4SRr0ukxx2JtLPuXfPVvbfWsHV82P9odvpR
aQRZkPH+piicHoDW1y8H5/d1R4t5LaB2Jq+gytpssbVI3hCVkGsT7nh84W9RNV6A7AuY1NWqXoUa
DN+G4fP0lk1jM9nHeUyb7v7OLZba2XUIh6I88HJqhmM+ge0/PtVaabVIJ6DXm3hYd1+oEx2RXaVI
kgwuqauJhbwcjm0WW5eXUsImMX0iOV1BF4z5rmogI5+zIqnpPMJrRyE3/TArgx1XCm/eHfrdpAw+
PtMfNLavDj/AaYUt1S6N+xbKCXsv7Wl/aCdI3tkMyQ8IXguhrid/WdBr45YO/UUcdvhIxOIDsMup
ZtTi7ttIlslLuos/AfAXH3SoDS2rTnPyRF06cu5XwzHW0PoVWKPhUu4N+qXKtldhJMiY3dKCjlaU
Ea+fwtaE+Hd9mWxrEzHF7CtrryXBKV/M2kR34su52VRSZtT+1IhwVzTlKct75sAj9nRmBp09eH1o
Dkwf77CjN5w5A0iEB1A36tScIxBB/5ZbOw1u/6kRM+FYhZnCv8TAA2SdQWVyBIjTroLLVyBZBAr2
izn16g1tKFnNGsNXeAus7rf9grLfKQegxpUhLtRGE//VzTBkFwCN4m0Luw5EcjklqgcFcbM6cpgl
VQI2WT6o/YbrbB9o4dZqintU+UgGfrwElJM+10f2oVz5FqbXCKeYMRIQxeSGXaz4CbZEYUIJWTZY
4udZtYfAnCmpE4uFaiAumJ4RnCAn1eBWyAaZCdGv8DTrLlvM4QttvdfXLvzTyP1ozfmaimSoLuzt
fK/d/KfDP06cEhAVXT1nb+J0Nsc02iJL99t3zi4OYXPhCdNPfpvsLcLPCSm9eK3L34QdKG2rS+2m
evfk0wyK2DEnE1nngE52CkoNRfnEqE9s1b4cBpb2sjO7J4FGJ8NbVqangIRwY4w/fR+F3/0FaWV/
PWnClZV5Hg9GdmwZFdnCUD3H4Y0HGAiLUXmdgP8V3F/hSgVn4FlgiClND2phuS+gBRpd4lq4BULq
XKU/cSBMLecCwstuIeftJpk+8DFWpYz9GhieHbE2xj3D8iavFxnxbPJZoohCQ00tmBMXQgo3Iscv
9ti6F9sa4L1WyF08VL8PmiXa2628+QhTtlHmyomPbX3lITRQlZtZnrJ2Pbve8wZOxerGiid0DdMG
K1Gw/mLAxQ9MCdJBQNqSJu8IXHbbvjK33CUrPTqhvjIoZW1/pL50ZIWt2SGUK7aSfcwUiw+r7YBk
CwWp+bBE3SK6zWQ+HTNKnVlg8fgJ4PR+uBBpyCqAoQMNLewzxWlCTk236O8nX6UaE6Tx8KVmdtfN
JlG67nTmfFEwZm68oeWTopUQVmtc5TS1KOO/AgUr1n/XdIhjgMb5V0nGKd6Q8TLcFhze2vIpdw77
e6vCui6MYhZubQov5VZNtHVelUYPLZwQD9zkehVzr4Gr3Oc/gWlBHA0sp57yFEaEHhmeFvwvsifB
liL6ukuERWCRpyDwfjzJ3JQuElR7eUKUpZXfrbgCap14wPxZYNE2blsqXoIoG04/FygKVkaP+58j
cD4DdaJKSmNI6kOn7oZOWRjzMuXp0iC0QDr6I1vlQDATFhE8qgS65OVZmJObg+UMuNYjPkJm2AYI
j11WncU8gGkEgY+z6w+PXPKas06ZNYxyMYLDWZxH8tNiSLqROMkmcPxxtHxiphLoINFEx3yJEkXD
ACT7XGXiiDjfxA8UX2DTqCBYn6wZVFF2eJKOA6MD4T549kzG9hkU3Qx1MJbvtZOdMJCmrFEp/bMk
IWSHJk2Z9+U6qwnXoF4SxX0wgk8DsvkanpaB2SRflEkIdgkamY1Jn+XLuiireEyCYWiHoWrH0H2T
yMKUzpMFfRYw5DCnh1IDhyi0UDtSPMeA91IgxeRMDg0tGwScPmr2bm91w/b7YUXDYnml0XrGPr5A
gSQoD0GbjpgNA3HTfZTHzHVqV1k15Ni8LaCAxaBt6PwHxxE8/ReKnYs57Z2pjg72aI1UF03BpOL0
ZZBhEE3mPks1scaMgECVp0PZ0wTklNuYGkx1gHq4BnCPx/iZ56X28SHfuFjRO7mwI4pb8HQM6mqC
+bhXHLKSfwv+CQuHA3w09tZuUiUvIt/2mH6CsEiwiWgRqhU/oOXv9yd3HRcaIubUMV9dlRvVvaHH
N5JzmTq8xzh8MrBVdgX7nUqH3XnhThAd8doHtJtzIe/XZ86ci5WppTywKSYVCOiySAeKk/0svwah
VGe+cxxrIeMlCDoQoFCmA+wyCl/6b/nPWaZI2o4x0+7umZ1BzKD6im/QampgB2vpeLB/8ETEoeBh
YJVXBveXS9xdX2txEQpR+ZJajkTpGXETWqlEgETVaYC4aYIcJ05cCJaeYS+k2NK6edE7kH9QIJgQ
QlXORJD9pN0YTFJBUO4p3CCu+VQki5uu6gQlrd7l8HlwpMtHbQ6+xQlx/xftlYptD6B5uwm4qslw
ulJ8HRpRbiZfWdGoNECXvdEqralog3Y6k8aSanxQrpkMPSRcY45xQR7WFAh8QrdKJ/C3M5RZ5dJP
4pAOCVZ4jTXT2x0UssLD/csEa41efYkc2DFfk+Hw3Z9HFfYuEDS0LdFsNrGFi/RRBaZiH5HVX0t8
WiRJh9Wa9HMqprMOr2VpoR9wVqVdQExJRX9GAFESgz9huKhaGF7L5nHXH1mJFsZJftMB+t2tfNDG
or5ejqMCaR4ZEaM3GcDmNfdxxmJDEcaNoS9YDcOwJKpn19Qh0gWHS4GnMrstlv0cQGBjNRDCn9mK
tONhvTmzSKuQb+O4buvU6j7ku1FKyrntv6zf5Rwhlj5JQv5mPyGXQ2tpyWCqAIeSOeBY1Mla+MdY
R/scxVJQWrtjE1KOSHMoJ1JQtAhFgOGQCXWv7VUOn8rEjPAR6AS8j0RLi/0UvQ2/P8tGwiUhKi9J
2BBIwmKdHLVpNfF66TlLD+DHkjn/MF8qFEwqhL9vdfmPp7+Zd20ppuKSyIWKi8FAOGM+q5KN7W6W
Z1ffG6nOSCKB9JIPY+ONumEzT5mnQTGJirJVI4I1zidvs91OILnRbOvAAlbqMPK2yehmKq4xAYgj
J3jjRJi8y77S6d0bclYs/2OE1kT0/qPpBc8ryq24zbx1pm3CoEN9j13jXycI9tnVksSk0Ina1SJB
Z178+ScAzm1SYpzJjfjAFOxvfI2STtgBDF+T2GbaKukOpKMHntMMx0Xew3KLjWDVJz143fRYZnCJ
M+YG1NIZ8POB3C3bXtlaDNw7+usrkCoanRhvgryxzGnStcmvOkC7xvO/+tFYduxV9XFVR5kLG9N/
0CGhvcqyod94g8BgUtKbtO2QbHQ8v4EV8venMJwXNYQWIpV7cvoVTbLdC5vwGZMfwX+PCM/xn2kn
H5FWJVHMx2HvbmnlnfTMEsdLNdKqQk483eZN6GMHSIGM/sH//xDlYTkB13pbP5WyrqPEsj5N6EoW
n+9S73a8+qy7BvmUXWoSbOWCK1dNAiDm1Wto8wnqLarpoYcO23/XuiQmd8gQduHmRGPVEAOg+46W
KQvY+R/wWaJVJr7pcgSlDPvjF3/Rj8zK8vTBBx6NGavU6yqKmf5TfQAJTupbn1+PmC3FBuyLuMIM
RndnV4E+O+X5uBIY5Tf7YyqL9mzs2FNZmTMzWWp2CZIdYXXcJrlOPZ9Nntz8MKVOdp4a1YOkJCEw
RylKqqm4q6a0/muq2LJHY7gVM6E59zL4STXwF+9LJQ6Xf01haSiRlpz0Q8MH+3fdN59RmacCxrSl
CADQiosICHXtuj8olGJzie5TklUcnz7y441CMo1n1pTBpePZua1H9SxtCj8VbCaTTEQcvKdq7PUz
tFDIpc1GiQObdrB31GgRHvxiQ5mof754fVtNeJuyY4/O/LQi74gSm4nnH1JHkOeUw6SmXsqYBfOG
Jw55Qsgw9nWfr7vgiADg1dnSdjVx6c4iIqaM6bPivANA+VEVTFaB0xQhpMjKsDPnwJI2yML6wHzn
pgQy7OKLx9fTqdc7OkRWV88Gls5xidIftVFOwf574OwalWucgUYTF/bWYJ93guPpg51x27xAg4k/
n/sLMqBPNSbpAxFP/NBOAPJWPXdzkEUF7sdJdhaIl2GF+Cjy9WSGkqJCFqeBJ+2qfiBgJW+eWLvU
S83YedUZ8INS89KW22hHAx8ApU7ALOdjHQwSc4gbemgVygB4noeFmVHCDOG2dGvtp3ndxUv5BFS9
rXaDt+128FfyRYG/7s/nZdBw10KNCPsbzXyiEHU956xaWkWl1mP0V7mK34EeKq5ud6F/Rd+SJ2ja
9yAJ1u8i4xcc/BZeaD6Ci+6SrqdwMs7kD+UWX1nyD4ZY9ChCk1bdSv4nFMwAlr+OJ49Y54fMUrNa
N13uXtGDEp3ANNPj4hLfXq+oUsseFMH+7PJqd1yzYael7UshNie+89LVJIEoxf/ea+ad1ia/xhMn
TGz27p5+Uq4CSmZ/wqcERL9kRVlgHLX/AESxtTYxV+QAb0WBmTIs0HQewRPyYO9t/bL79dLJfxi3
qktHzhZV6QY283n72V9/Ey+SYS/q510iPmVo/Si9D9oF8PP/HXNxgSwxGbf7/90teIo8jNRxWcuy
2NhbhTpdXEcyMjKibhLMkrav+JoXDxw11CNiIEgdq83sstSG5TNvnqOC4EipOl9UbwGUP3leOWRu
yMqB+OTo/HICC9E1DkhhCr3F9xQsAoUup43hfE7L/z89hLsQol8uhWeojEw/Sc4XA6/o8TYiZ3s5
Bry1eVUDufzEqwohanzzcCxZZhwX1bjjomgz39y5FKQjGxtr70AInH8vde4meXVLZPjAVRQ/Z2lf
mUqUFYGtpsfqAerCGMmBpqqwDrm/2xi1iHNHz9rmS18Fu6BLJLGZWugPlp37f+ZyBLeRuMwDgKcB
bn0CcRHDFo5NnyJwZxTppSCNnOf7PBSFM7qRutLLUEd+StsfZvLKbvZAge4XIYztuHd6lNQ858CK
o5e9fRLU51P+zrHR1oSVg6CeM6wGClC+ghqbNkHtRznpuNkOUl1pHNqO0RJK/JOERSDCkFXFjSrZ
vjWBeZk3je7XlC1RmzKuQ0oFMYx2gvc3cE5HiLG4ajFRsgpQi8t75wa2BWjGaZYe6BHbj/mffnq8
kNrUtES/ZiYEODSrgHSVmngH0ClgSEixNxEuhjHC+gkdhqJNIRGw+v0MTH/d5x6/c5IW/t/80wiE
wCBnCdxqmbylYNFZs2y3dusquR0ouJMG8kxn10wCXuGzNmb3azcBUfsHMt0eGTdMqFw7kD4VtAvG
iPNqInDik+DZtEQ9SITpRPW5IkDKrBbSb99v9XoGGjppVrda1fKzDr/V/NNz/oz/OeZWHCfWxwad
ipYwUBPXjlxY3xLK+vzbB7RDQAgSC+8XBZVQ5yd1I5irgPjCj4RhbVpgU4t0BirLO4EyKpFsRm57
lklEfSwbx8NztS7S5JeuTSks2p5cowTxCYMZqJ7p59uGc4Akzqs/Jg/nMO0OUZBeAqnvPggG/mpy
gLlvwMLGo1ME2ROclX8Dlg5PCHbsvLfgrceW1CYBmSiHlJAJ7DHWNQhjEwzlughzh4RlETndZl32
Ru4Q8g0iVvjupvDzmO3Dyj2muPeuOBRevb7/iLIzYgmMdwx6Wrx0/U79i+VCOvRl9Tri69U1jhf9
KgbZkhZJoIlSx0aAL7o9OWy+VI4XZaIU32Keo0ommK1u3va61DYz/mJoHQMIXMyuC+FwRRDqtIo1
uSBzHoqy3TATh0OYpUrDXQ4a6xSlcJWrZctd34XXDyDg6u91zdPj4rr8UUjn6rC5amcnABykW+Ck
RZ7/Z6GLxzS7EGTgd6PulBy180tUp54L5IQADY5ZUrJvH3P6UePOgLZpupFaqgpw11ct20jF2CxA
W8b2uAjrIkG9lu8F9VzuqDL2fgTFC/2G/9gM7GcgaPQ21jqRglpkY8r7uirdIo7LGuHMFOpG/1wY
heknYObKUFTw5pM4UeCcJIaGA2FBaAbO2/iArmRZLJ5wz/dE+QwM60TZlOgWxXWGyLoKZ8jewPZH
EYOWss6PrwI63Cb7nHhHAIA0vubmwAR3TqwuX3lo/hCgOrhJGP7WYVTzKvw5Hw+/CTOg5HwNQaOm
ZKTufuMBJ2juhNU0mfT2vavJQ69kPwM8Ks5GoKhmv1jppxq13C3QbA+PNYkjvHD0RXGw9jMtZaUG
CaqVViNtWT0OKsA1b1u9DItZbmT184kqyXNV5Vlh0QaqneyI0b/f2ulIPnBGTa0WsHkRHhcLjKzt
z+gB3/+OgUPtR6Ml2iiOCOvxeggEU/e9NIy7hlvOLssEpoaVkYcRG4rTHA4Ettl0A373j2fRCvKM
6E2N+3/AYCpZoAT8wKxIwapifSsz00ukhlv16SSlMB1zWyaPa7ioGPWJcz0pF0f75GIMHsR/OV7k
IyfgMyN+5PKcUTu3QgPsBqddR1/Oy8U9wHoFkkOPz/4uKyQkucek2/jH+QWaam96VjAwL3ObtkEv
BMimpqAMRZtdWl0e2Q6nQDAtQntoZSpyk0MxEkryzwsvM7kvS07diFmX2kDK2XwIQlay8GA+F2g6
yC7mqBWlINTT8g39nVig1FkOnQE9zqrzZvAm6KHUTXjoUsx3MXPYoBRu9Xsh6mDdYzZvTRxNWaY6
j+M5K9YymsCUWw6UFT+iIZAYQjzf5R4YJXestebPA61aiqwpevEjHNSexVZOnRhUAX6tnpgBDnmP
yfsJLBoyFWvWc3p+nRo/BE4XYphLC6HF/m1uCNbmavAdYSb4ivz46GnWwkAKrxmv8d7KR0XGwOqa
jZC4MckKHQ9O2dreurlAvPVkdNgtn4kyopGy2FRFifs2TiPInwbz2/ShAQ7QriOZqY63Hq5lBvv/
onFtGUsSemEDlDm7cLVfulLOIickGJLGeXhu+1IxmJ/Rq8keQoO2Fk01P8ZjQDqIOlnYYv4zEBae
gotSfg4Lsrfq+fk/4iVbByasN4m6O/WnYf0KoZIt4sCN9i4VEAhJ3qRceFND31hy5O0CdgB2xyQI
8hYBs8nGIZKWKlhjdLGS0jeDS0pRdB5eeZvSIfuojX4/xyh1I3OV94bN744KK2gfLLWjZo73nZew
p2surhv1WLV1n3b7xnOWn8CvfpCLqrwuxBH+bDxuNeQPCumit93q25P3GhMgbQh79TwSp3AFOnFt
qBr9UzvsM6gGckhGN3jVyHb5E/M0Vhhzhg3bKKAgqtn2hUht6aNXPE5s6RgWpIcRnZ0RgxwSAuug
sV5MOEqBSFnnv9pAAiJWeWUVHr3OaykR4IIoB1A+dDHxIlUwXGTz73YpWxqqgvP63vq1XmW1/Dhm
rcPG7yD39VsJRxhHmPbgx4m/tHUTBsCi8wDJ3HqVWICKLqJKkE1P9aEPJ0qB7t0OH3lDT0r9tWDJ
fATa1HFKatwVxr9aDL7skTv77Z3cC0UrsSuukq9x8exsgxYCk7VI0IRdB4cVB5+kyEKAM6jKKyIp
2ml/lit5yGbenyqF1ptRuFcbjx6/tGI+w/95iy8MtkBbo6JqsuNNT6AE0zhwQED6PU1a8NrlaIAj
rwnbXMxD1jFr24RXNwACtpEtTF0w60jsezLVc9Giyy6XzY9OYy5A4YkQinN7ELXtCAeMOgCE/7mu
br/6VCsjLXUP1Q9Fi6EMmISR+kdiQjS0TaDswXy/9CX/WFUZGn7OvTIqJ8HVa28nuuJM6H4PMMEZ
MUctfQjhpFlic5+oOR+8XTw5wctf9lq7rKoThB6UpHOH11T06RoIZ6rRUaIFVNDqFgUr86+hsYQH
MB2JXN8Gx8IYFWbLO76kw6vezJtO+cxawYTkLGG82YV+PXxUcmNfOC3dh9fk7cX560MOfV56eX5V
rp75F2DCR2ypFsrxCgSWE8iUw7xkWPXzgWweCIfgUrzoPe2vFUNvVS9EQqChqY3IGzlBBFad41qB
LDXctJCkGLTjZDzb1VOeZxMZpjVVR7RysUp39HYeVngwkGHRerFRfGiUnh/nmKG67K88mUu4f6Lp
7s33IyQibJiKqn5+OYtfffICG7QyXtY7uvdH2+bQHz/012dgVFAhMlv2DbLUXRfo2rUS3IT0UFKq
zPCkYx4WnlYiPvGynmnSVPjoPE4r7nRd5YBUgNNZ+NYewpCXESuO7kIF3RQ++MchQ9W0kAGYmyih
NDKTrjkRccjoDocs+umkA0H+nNFtZ7HaiMqtNUdXeZvsXY6C8T9OFCeO6DAd05FFJ4uqzhPwkVAB
fM9rXLO6kS+Z/weS8oFZjxUZ2SmLEJ2HiDn9FsyxN+RG6n/QK22K+pOiyiJfdpkGRshjzynET4sP
j0cF2JYApSKBQhzH3EJgZns2Vg18uOEpxVSBbh7mVdsWGN4fnkpQxg3JLZtxkOt0LiSl7HMybjZ8
FGLheD+uxm8DSPXyDyeJGFVTUZcSpS3ptOM8ks0/8dG0d+CYoHo9xsb9DhUIxU8PBPZwJ4bFlch3
AOLJQLFSq0kWtGanU5vpG/gdb9jGNluhV92Ev4Yg6cTssAu6qgQa23ZjbXKJB3AT5tcALCOtEcDl
sNj7rO+pjH8I4Rkp7gELIWwdsiKb6eIJTkVYJktA4gCUmH8U/8JvsJNRLl2WXbOBmYTa+eUvovc1
YgtXEyP1/9d930YXY2uPDvnpCNbq21mq2fGRDeQYqc5mso/FppSFNZAnF/N5zo7RkfxHuPRZ35Gz
L1VaZRd+iICFHnvJz0mguNf1uRLNQbyazQv+gIvK9abdnTJUIfYYxDiyZSCr7lsWPYRDS+DOM4Lt
APbb/BnaBDB+jlytAYyL+dBx1NT5//NGIEDM5EGxk8c791bTEftoV7CW0knqYHxswbS5DSuFYTGA
HAhwbEMwl2ukT3lSUY+Dy2hTyMW/498I2Nq2NkCKhn2uNDnUtfWVy8mRE5FXEHzy7LKtMtiA3iXu
LKGrbOTVUaACgtJj6inLnWoKTziev1fZznaiOiZTJqcmi5CcM5GT2NyTyiF8AylshwQavRBHIWmR
qByFz4aIt9bkv5aligusdEWWvh7FjwoFn7JRSRKiuMaG7kx26rlO/MblI5IHB3rebz0orFi9tsmF
NZ0lI+EZA8XFgDr37vovin0GSfyWX6tD7rlTDbBHxG05DJ4IhwARO4A6a9wUoVr2hTkB51diR8Ix
Kl6djGjj+zEua2Ws1Ca8Ba12wVyNPRLrqESIaHB89TCmIhvgokJ0SGenG/YbOXCrVUH9Mu8Wr50J
MtfWNn4UEwqqWNeFVbMXjuJleSsNhSjhxTyaRrPtj9lecIrLm4OHKxP6adq5fh5NwxCaozhabN+C
YIDLKgjXkZWRQRO25XugfdqINfDIUgsTxRdoCbQePS4MkVk+JXm+WfFSoYBl+ejm8mK3UIAg+Gy7
GOuIz/G67w6KNrMgVfSGa0xBGL/uii1FX8HPe/X1FlWxhgU41wzaayzCQAFWl//x8sM8M9IzrsP/
1fRoezhcua4foaeekCloZCHfAGIB77vyipH0tW8lGEnKdHG63eLmIOFOFrZodyWCM5cP813258O/
1uu2KwYB4ZS3oT7+paCcZI03Z5s61H23jZDMz23RBuTCLQjvPWSCrFjp4hj1BMZUWn3QxMdPiTu6
waGAmPZ/iH1W9ha66CCSYlKiWzqbxT0mvgYC98LnxKP4UdqFzyr6jh8wzpY1UA32n1T5rO1tSTjz
6RbRDzBQt1UHhUP6rG/9zBcqDSXmr7U0ohQpAG2ac7RpT1E27KeV7wLUTCD8JUMdPe7Nlh+Lo0A3
+5rh3oYe06fKE/OawFrD+wVFss/CquE+a8Nw9OyAbxeEADKxpCpMwBBf4q5hGQ42SsAQUcvM0wap
pCzzPrfRSJAIyKxyR9T+Y/ICXl5Fg9F1eq0KdVMaFHnjavscRAKR1ZNpH2aMLFzlSYNZrNooPZuE
eF5chu0FSdo5eda6xIZJmXrD4Yy0DPxXYmMu3i3oRDIdMUCR1GCXm1GlWrZCgvZ/bmNYO01eWz2t
NNej3bJKiG/t/aMpqG0Jz08FUWGhwPtpPdxp7nQmIJH7iQWUOpqKzc4oBE8mmaN5j9I6uqvI5XSe
edSr0EqKB+DP52uNdHmJWqCRWlxnxpsLPk2wPHNU1t+fArmZXahMWQvYL0FPMfcKsD/GIZ1uYMBt
X9IIAkDnKacPDaMvBc03QkSJinF/sfoWmzm54W0gwUIUKPuwwUQ7pX/88XJVRGKMEQD5zxi8bmpR
fLEpt1TRts0CcIfomcaGF03hYhCrkPN8DuFQW3v0n3n0is86QOXSF+NR2vVLdtqJ3qbIfrQD/jKp
54B0ClY0oT6HN3XZSD5IOjnzK9D/EfKO2p04aSt0YjXd9YHcIqPfJczfmzDY/PVKuNEMdgj3o5bN
2FOLuPfaAzHvn3BryEfSdUkxRJGCZj5a840GNyLjdycrO1mPm4ekeOp1Z7nvXCCOax1rnZzhO1HZ
ohej8deStomhpKIF/B7NebmNk6AflURxJE4XA+oxLv8u7I3UosLaYamjp17dq+9royqZcy+/RUn5
CK6a+55BPzmTCq5lfkGjvogI4aAAUx8PQV1+YQ3e4cv7Z9AZGLwil8CrWqxl5LJQbjspIKje7a6+
vaVEWNbjehBEpxnlNjkbKdXy8whXl7ZupQWsLavcRvg9ygS4sR3+Ufkwf4ytOm7AAH7xTN6tH7//
szJuYg+vYD7GVVCAkWJXgI1IZEJBQ0826eQHaCEyh2fPTMZkxRdtOBVC7ZTzPOBnB95AIpDfgdDe
4L3qSzER4FIB1Av6Y/9UTBjnTKpik3DUh2TfQgbUAwZg/cM81IyG9ikYd0I0LsRA1E6IVhEjvYE9
VzdaCo9BAMhx9/QygXkkpSjBgtRaCzLRz5C2bsGNycDD2RUyyYPmxRlJ1zSd/wKW6NWOQlxiJB/W
EnDuCZTWTOQgIpzNOj3sdPvnq8DU+D6WSm9lVhph13AEnVX46aG/TLfBbaAC35cgVwpauvP6MQdV
/QC8oeo1PBuCtf3VuNPJGodERWKoLl4QJAU7HwR+IDOI8tF/fQdJVJ9RI7UTRpotLclFV5ORGSwU
gIZbTJ8mPjTKowyPapI3gVgOa3MpymqncQ4WCTp1LZOgtxQXajs14w0V0zDWguPWYZ8D0PE5UgO2
ddFcBo35esgK61Wi/wTevujxtDmR1Z1Px2jc8PKD4CH8fPRTN3N7G0QCrTfhGYsD719Wlci3cDeo
pA7V/xvj4fHe3sRBZf4cW2aJMnJW42vPlvow87vcpYQqVmCTWk7iK8syeuLyLYxB4/sKMbHwy8I4
Bejp1HgCVPAUmxBeBx4y5B5/ktYCftBSh80bodpzrRzzy+zPscP4zWlOq8QZ0lBGveE6kjC0nP6L
gZq1tt70dCV2IpwVb+Kp5uMqfaigN+2Yb7cBX5YOtgMUCxuJh39KLHJ4S3DlN4D459prgQ20cZI3
i1eu0EcVhxQIhZkwP3v08+Ev5uc/FQ/5D82A18+LXCn5+mqUonVh21gxly8fuUU75MrHdNx2JaYu
2xWQrsluZBMHI9CwE6VQsAhwYEQXzhNKxPXFpOKXfTez/VcdwbVgNQpoMx9j6Dx8iZZIFa0/3ciI
SlHzBWcxz0rmpwxZ0pdAU5qE0TY9vwJ/jVBNXJSH8KaWfh/GGpOxsyfK2vDhA31fqRM4VdODHm6K
vFOiOVLCFNeQtvoxOSUlKNA7WcoIKitAmd3ylmWNVNlZJ3XwnLhs4beqreEKSpJK2rrWE7TdjbwW
scpWb2WIHwRcUS0mcNjYsJsgVszhX62C8IMszDqdsChApqeSe4Q2atZPh+oZLWnH9m+l2dvnj7gN
VE0XQjyWEekq0mPbqYeRQa3EF8wu8jjYPc2N3OsQsS+vZpdWc5U4rjORDiAezWwQOsHYROVcQ2gv
YGec84VIyLHAfBlPWxcHNb6kvwZsnFjSLqvb6CGQw7feGdxLuxEja1XxdVW5qHbQmJHq3gqS8AeR
W83/Ku09O5JMwe+552fqor3B8BKcukT63ND+WlHVagcPPjozQb7g57Bgc2ewWxYj8I/ql6C15Nxp
L9vs3R9mudCn/M7fCIQLv0S6GLNNjhnZNrnVaMfRh6KH3oG16Ql8GJGE550yl6TBKeHnnbAFQM7l
FApVAarf5Z0QhibzN0xz1BEBLi925AGGaBF7w40/QN4MUGop8/ekn/VxbYdV2LHRZM08osA2LkDB
yggklcuWsFPP3ZrrNxIzKQIFnKz4SVGLZrdRAv3aFpvQ9TD+MbkGor4Wl9ffolYiDc7v9nO4v6D6
HRjXoqWFbCa+OVyUrXpdfM4NN4cDWzSytpmof2m7X4c2jJ1zfzipqXFH4fPtcPssy+ISMOp880Ki
bUD5FSofT0fR7b1qN5ouBkJjwttvkp6RGGNn+dt5OVhVCmhBKRg8EctLb0neziFB+DjuwjMAQXSQ
iufazdSwiEto1GWYBISWa99an6HtgL3WPOUZPMsoOwCGXc4ms2k7GasDXs7cBNo5b4+0Q3F6Dowu
2SCP6nin/CQTPayE9qPx/p2uCatf4IcfzWukd4eiL3Mx8oT9Bv37EUj5qZK9gIGH/0/yCQOcyLWu
E8nvpsc9DQbb8zJ1ULBDMzLliOsd4Na/T8FAMaR9VI1Wjg/8d0fm4kRlJuubakvmx7l7cRx3RpBp
Tj0i7affdPAux3h/ecJslM5QhpjmiUcTzwJLVMgaslr9VtMFuGv8ZzAJhucn6LksgIct61JZTgZO
7TxCcNToeCrgXIm69KOYLnt5lXfnWfceV4IS6+5bpShfTsDpJY7O9P4pxweAElAQY6nr557g+dOd
jqpBk/alTbPd+VlGyPNftvNxY3wWuJGTgPit530mdsb3vFZfEH5vuxVjph4SQ73pTbbhG1AoQzvj
35HHogi0uNwcgOn5/UeZr00M9NXKAFVYmlVQsuTGU0TgqtWtrCHy0OU6fyIZ9XWdhqTJyW096EJQ
4GulM8gC+HZyG4gaMUDjJR9oIXhnc7V7QCn0NovW1yyJl+rcSbEG+8eYGtdQ66mOD1T6xKo0Uc4/
j/XfdunRkBbSdGSJR6yvE1O+xFep/tuz1c3ceYkrmb2ThJx4aL7oTUGgzeNYZnWmy0IK7Ag9NmMK
gwx7IVrNrxCK7FbzYa0P8E4049AIVS7w/CFSB+RcbbpGAgFJYorKdxjF2g2rFrdC+zKDnnpJsRDF
ZsGIEJHeAESQBHgpMdD7CBHuYaJXroO4pNEvZjxXBdr0G3UJPsbvWmUACzEG1+nToEO45JarUMUM
RAgkgQkwRUFHTEThprn5MKCEM42EygyAsX4y1ntHz+v54ql2hEDokFHIFF4N0fLR04BCSsb7EiP/
fzNwE3ocGag0Z7Bu4H/xq3cGRe3CGTzx/lea+0+iBLpknosP7bMUSByGEEHMcO1vhZozN8lsRW/4
j/GIrlwHhvpXFPWp7Zj5HFf+QyysygNbuSBg6+hTdG0fMXjhomfwbwOjhmSls4/5R+L2sCi0qclM
wTltNOELEUapRAW1IHNB8OcrwLplUcJMQfuMuB8oGzXIAyz5NLr72CGnQpVQ44urvyGJyPBwVyLQ
kSoIyoC3R30xsn/tX5CffGrupcXXeiDj3EM47N4al3rxuj6aLQW+Nsz+bJvN68xNxkFvIlXpiQcH
IYK/FGAZjsUcW+aFPIpKd7Cmyte2L8v8THQYSQBKs8+EzIpn/4eTg1shhCumZ1DvguWvdPxWrp2o
0YfwjT+Sq038a6FcR+ncmCngRa1nCMVnIK9ubxuMY+557qfb/HgbvQB6fa+8L/DYvEwHi1qknZGy
4DQE030l95inSc4azXMJvKPPB/xnecgtVRZs/nlohpy/tW9lsRtubC6h2sY1qy+RjX9Fglfs5rny
OAAhrqVGvgAwvqJUQejlW5ROZ0WG3Ph3f+CtDfTn3gK+K6dCxitU4WEaP59efkR6MWa/TU1fKJ2x
e6pvmZMtiYd9KIBN9scbbtkyOiq8i3eI89S2/5ehdWOeBYhBSIJOgRGgdUi2nsdPq8/GLfrUKlAC
G+nfYgFwKs7lGHCL7tJ6jbb4mBUFJQcZ2KI6naM7aebIuHdw+uq/tj7iVBSRV8Sne8E5oAC39INY
mk6tjBIaBusmQvDfMxgNilMCZ9UPUqr/CBD2o3ULtOaMnU2aNPdHQayXPDKphJFzPyaAGkS5g2ip
KIJ9/wc9IRLXeSg8prY8lSBYyEmQpW7qvgwoaxVNBqbhwgX/1SXCjFzwx0YhMcBajjUs/pXKUEMf
4rIRszTwSsPxErkOUuV2rRyABw+246210e4ZitkLGolYxeHendua+3Co6cSCSE66jXtuoj4bh3CK
W59/aWVwdbibmxAjpn9ET2celgh8MJV/5igAQOnAtN3B1LHnBNsgUuBf3pqxJJAlGDuQFjZrrou8
OKGF8sILXL3+EF2MUboy2n0PiWf5467hNCbwfwMQMIqR2lMex2jiPYPl9qV+Ak222LQ5wO24msli
8ULCoAyfjMSZ8iMztoQJpLpLTG9baIrMFk1g3mY+Fc0B+EAXSFDozHD9dTeA9GfLW9dEJk9Y4m/G
8Xy1BtfPVYeru7D69tMtBprmKKNApphqKf0nLjyMz2V4QlptR0Yy2dHm3JqzO4a29mwtOtyo8c1P
nlBf6uWMkTzlCJuanT9pHOtEY5IVPuO+GG0rtixCyfvSfnjmQP+2EbnWZtao4RIrTrr6BJJCrXoQ
e4lwdBSohNnFo5dxgQ3SPaRk4yNjzg/TAF2RLhAvY84LNLmR7ZpbmJCGaleh9L8WkScoyMkjIT/D
5Ic70HZgDBIYayMtS4b1J7e+MfYpaeHw/5KsPXJ7gNkasLc4jqvsyoeHCUa564zMNBJKGZXJfzwD
+agsoPu+qNFwJtpnJqsKnQYRIVfA0vdm2JcWz34XPW/oTRE97qSGx11qts0pRamCHCn3EYBw4jBO
lHnrjr5rxZzddtK44uS6IwVj52+qbZPD5Izkc7/i8cBaoh73ddjejggcutCn7p3fiIiFgU5uSwIM
ofvhtQmur4XAGfqTUp3UsptlC+cKLWQml5yqGdwR76tb/Asv5mJ5/eqBzASTMLyMV6FqCiDSr9HV
d91ZFVH1SULq0Inkp6XMEjXl3TkZRiJnengBc5qwFpogxs0wLuqnOH4uuLD+39LFWwlmV0PipnMM
3KbCdZCsF1XoRUdZwvJPYlwfM8rBAM9LTmFzaRXkhlJQtVEhXg72uuMHXXnrV+vrtaZxrMrwc3Sk
l3OZDiv7bYm9FqX+KLjYr+SPb9zmh7FcIL6dmWDLL/gyBnTR/+GWhsNqTcUFNFw3jpkQ0LY+G4Ib
60xXdXKu5m7mFDFF7D3juD1QYhh1Q2lufwg+dm74Hft9r8ovVlO9CxOvQJ2l0iaHjtT62No75Nt7
/kecjovEi95iyqm5ILbMKt7UxRQ8DfN6U53JrfWCV80gjL4+gZX7SPRyYIQltzx0CmH978DfXyvH
yiXRz7/vYX4DZE0UOejuLdgU06GP8OcqrIIv/fgyYpyJFVBhZFo8zfLqTDPNsq4EiZqYML6noZbg
bCTdcbSXAWnk3IpYCNj6Urk7MWBRBCLJxVBjKEcLTuOO1yUZ3GxCRi7V09SIysfD7IHN540hDniO
8HtIddf82OugJAUolmq6Dfj7vxnDrT8amcL/MKSi1VbnnCP41+Ol1Yx4haT6WwFfz/vsSh8vXkrv
kgnmKKU9sXpYNvqPBbzTNnYLh1zpYHNgDby91PVQbPoL2cIVXpN+APQCVUC3z4qQdNic1l2Evcsj
B64Y0vnPMERmNvG705HbCt3HajoEqHPmoisYhQu2XA0Iis2pbf4QarW/+8BhMV5rZy0gzkiaWlIR
6wwXWdJSvPrqInzhLRs/YrCHnGyRzJzsV/PjNhJw7XMHP3zAKzf0XdxFWbt+PTB2jLSOEkl4OQVH
2zEpvwDy/l1+On64o8GzpE04WqC97G7zdV5Xu4FWuikZlyzaR07yqmwaMASp0V/n0zjVeUvHV4ei
nkndIW1QS7VBVYg+l/LgVRavnT4z0x/ZXOb8n2KsazKXl0ABM8zgIDBl+Cuhmw+ENGevd2g67do+
Qjb2rEfqSV7u23Ovy0/jnu3b2HwXpMGBS2DyRKnWRNc1XVxkPfb4Z/d1YF+vNt9rrjI+kMaM4kMi
Wf+iUpMAbMhY4DhBlx5+tOP8+RWZGzL4DBhX7BAz88EH70+LDjkK4N5PpUwaPj+T6bqYOCzWPLHD
0s1hTTKiXmk0R8lQyEm5TRummInKo9IQDkWrhoHl51+f/UmCjlKONpyuPS6s7QrNcVJ+ju/LcWVJ
kviiVATnccXB0NV6tPB2+Wrt8x4ww3u1NyS0z9gK+7IJ15VC5MdgQSnt2Nhq014r/xTn13WWWy1+
gEvVitgqHC2kFAfULCYiOo1fUvyvo0wU67n/wrEYxR3LFyvLHbK6HvEKc8wAG2qbxer6WHKhbHlk
j9sLZTIMPkjeGouhAeqqL8AAGOqgWue4h4w/2MjmGqEHWe+j+0s9y0Dkx7RVQoRuMLyX/ApdU7FZ
0Cb5zI6DD3BtQSWNIiCuYA+LN/WgdB12jEtpzlBmdLwtppi5ZIZscJ0oazlYqosIxAbNOzkftL7M
Y89z/U+j9I7/bwlTgAy2Rf3HMzQneNzyVWfiiDi1tQpCQi42L8DqXcoqwDLimw5CXwne1vPBIDxH
ZAYFE8g5JoQzEFwhAGY/67QCBDzlcAphu+4Ql6tmidbZ8+64Dtyc85ShZ+zQE541yZhJvgq3s7p3
ZiuaS4AZzslbmFV2+7X1/ba49L1NhK+imZmiVlLc8mbn4rLAxF9oR4ohyQ8s0gvzjfpgeVzozaqo
L0OiU+txRh4EIh6IgZCvLI6RdWkD7AW0p9IL/Gh5n4oznYVZInyaXh5DAEy/V4z4xrw6MpYNkHsr
urOjSPNDaKK49uOgigKohvL4vJ1HnZHtaB8hjaC6MvPzvQb+GgIOrkrGcsgqLZTdjjyvKQVMAzFa
9B+u/zCJLElXARfbk3W3IKeBsZbYV00DU1VropFxEHz/Ohrf0XoztOpTuQ17MeajuzmBAabK8Vrx
ipPH8oUbWjXuAxfN76wzrRYaiPk77lfLibZ1MMlNTO84VoNa2IoBmFUj0D4IOMV5bEHkf5I4Zgxo
2RiGKZ1X8frQKgv1wzvM4ONfAVFmamWbnG6BSope80QBhufVoWrBTORIo90uhIptV2lA4LFeU7/w
Hnz3F9OZbvzUIhwp2TiLYCV+f3N0iX+O/kAO2EhF2vKhGsKp5P6JizmGCIIymvUsMioFkIDUfaKT
jqV+RTWKJNjk6WSOv0u7jLh5xWP1YzzBHEASwDyGKKO6FT6m2oTjeWCJMuLGwXUmAk2sUE9IzrEF
SI5Ui158p9i3DE6g+2cySds9DaYYK/TyOzJHuoKLnAeaMGqgDtgvqonCiHnsFn5+5Zakj3zpXRt/
qWIUFI/9iQ+7ioFYGmUMCx2uvPhbWamc3wmtL+e3TwmPfqBtkxg3elpBrJNZ2Q0wlDErAJfexohd
FJ/TFg33AhNnZH690UFKpWMZJDQZGHouUS/rNfp0rPVpPjpl2XaC1M2BboA7J5/7uCvcRsw94fcT
bsYFdysU0K63pgBm4ZDvuhh3D/c5TqKVGZydOH2nGpNGfNx5dKX2nxC0MgFFDXBVafB+OXZqdWyf
xUZ2C95IbbfBSEIoHPPqnYzr1gP1zPPaNbB8n3VdFE7Jbo0WWIJRcTCSkGQjhNcEj2GH/5CKsowQ
VMyngQahx+OOeKo4wEuIWuNiWuT3WFQanDfON/ifd+HKkA9LULh70dfopZfw/EQGGInFQdALSHBR
yZ/QAumZ14UNFynlPB80sGiSABKj7+yl1WQlR0xogw9GON3pUY1BKTAGzrTGvrXRGZXuFHg8IHNc
WMSik5+z3oGVqyBdZtaE3iSt4/oMvgegxigxfQS35ijeUBC+3KgEHvA9K5fSe6FUoWd9gzSHpYbY
Q5wb2rEP24EajDWNrmVP7q40+KGVcBCow2fboLcqsOojZ2oKAKwDdsKcqkg6eJpJ9I7DXcncZ6JS
Y7GFmFywM3pD/W8EVuDvWdGEFu/3d9r96r0YUL/HUueuaRPOEcWiE6FDBQ3hwnZc+sSRcY/DuYat
xb2wjWxDOBixX29DIw5EMrl2JwJLmnb5BxGjeENiQ9S6xZpOcIoRBNhcBaO7w+1xtS7UMytS3haR
xYQr8YL3H5Tewl/FOvT+fAglU2safMu4MJPD4h8hj4vpynzoMQ9Vw2sxuGsmCuqkybMJ2TAIVqxQ
lurVE7QCYp3IoPqQGgzkkMR/SgXtx0icKvnoBC/6EsV//ddE/zyws+eODVBfZ/86TPj/AfxYgJO5
GgGgR7R+Nx2GYFi7YBplM1iK4tDgnxVj2O1URpLtW9+mb11U4MwhRev6KQaSIRRW9k6NSRq6xgec
J2qZyWx77yWlopE82CT+0bBD4kclO/sQq7U+ZRvtqIdRb8hLNNSdu+CFuB0mTVl/5xK4bjb+JvLx
5oWnwZxrVdHxih8TYgg2bEUnyC3lG8PhkmALHVjkFzxUqzObqLGQbD0r99zZUtZd+Ku5ROdgGcGU
T7aT2qi6AZ3x5oyhe1Co2DFYK0NVlrpkik2qXknC/rZ2i7s4wNCjdpKIjLrmKDwf5mEF0eXsMeLt
TKtsi2htdn3GaQJHZXA3L+LqdPCazndzUzmgIGQ2qEmXcdBOyAzQbyDzNw/aYIERbo2SF9aFpsM6
Lom8AaFazxTVwX50icMW/LNln+kvrR94COedKGf1H09tXQaNnDpWrFCITIVuf1ykZXaUM9uZgfNq
ysdti+l4bqNjvQWoBenD1Hm8Oq65NWKf6+tX3gClanjqAJKi8CKXmDaV+SLwJcND4UMW3H3rrin2
f1wbAKkxV1DNAJrILoMWb8tXvSi5w8cd834PjSHer4ywKEDIZyO8eWRD/QH7X+slM3bWULVBjvVH
63Ive5PSAhR4AL3Kj435vAFOrxWMXCPUv92chvvKru3zjm0PDCpIgmHnVVhEGh7AqPx5KxxOCigm
lY0v/+Fy6Zc0x2DapyBPIOl6YE66C0nT11j78XmS3v9LgmJCh9tf5iDLYjNN6pvTG8jwXDQBcx2g
2RYlMKeCgg5MTDUAQtRFZf5d0x0qC/6RkuL0xB59ZtMiKS3azcp6g3DlcNwJB++4AlND0SK9wqD3
P0V0HBU5fgMQSRKJhGvNmqKD7PJkfRyBzorhbZ7DMF9dWCpBNfgT2IVrQBU9H+7y67qdMMUBkqjR
tFryF+IBOz5T530DByxauOXUszH+/NJcoS16H/GxDVilUNeihRUkC6MwxmQF+fzhL4OfOX+hHAsq
ZU8dDcgYihR8StaU372MYWCLiaPBjgLZIOVpjxhdJGCDJenwLemYG2MaiCyLDsAAdC5rdsnAD/+c
IEoQLcj3u9QNDw1Nw+VTFtps1txbeC36XrrobHO1HhIVoGAa8o+ZqBZ1OYMvNTMp/AjH+tBaW/kS
wNuE973BeyBM3QfFubWm0wO3p2XkPplJMJTRh/Oq2b/1f6hRl5/NkIDaPreUWTH6EBCpVK06yj5K
7/HsDFjwSLUbpN5sRzTu8Cevc/AKr/yJMZDV4907CxfkKTc+rWM6VCzvWri/jnB8yjDFmoJ5bPGj
lUjlVz7nYxLBuc7RpU6CTZsLWkuUEt/IrWO5kyh/QILwBRgHel/JQdKPHDzbSZZeYSfZi+k3xZeP
ENozFBc0M80K+tXV76vL8teHD06Y46oNLLQJNQA51zM5Tz0jW/JtYvd4He9I3u/Gb+f1IPhaIBFO
CYG8ro6Wf+xYs6DvWLCUf5xRkUF6Q+iSodiJBZs4NDCjOBoLRMpN8Rm6oj37p5/UHcM29JjSMPwd
8ISMaYr/7Sz+AW1DWZOY4x8xMxb7mpdVqaJETBaLJCUihAv6cvEx4tYzt6TpskV/sSkRymhxeCEW
EPKqapxfGPwpvPIoHJJA6QhfmDBmYAGM9eVZbcFl7qF9eSrkpC8ddsw2Vmog1fhs0za2pYg6wIXq
9EarJfVCLjs/FJ/auxcLp9xj2MIk6fsyHEfIDOQIJ/8Wo5l/a31JVQ2eX9YGJ9fFnDyNkOYr2ire
T1xmiF0F1I32hV5B//f7qqEqa90R+jDJwY1FDuwWSbTtvA1ZM5i92nV6ttjU3eUnAvVF8xckg8XO
wXBSSPsFSwiizChshBBF9rD0SOtdTxbAZIpdtlyXheVNLAZDfn7sN2tDUr9CarGqHTCl6YEXwKqJ
WYj0zOf2kr6vG50q+qKrdmzSKMbB/7OXkKyPfBR2H+Id3K/EQAmZra/5cDikJJOaZ99vMhnny7/m
KasL9puc7RDQfgNdUYlrkqmjSlesJt9VsIPMWK8K9+to7Amrc8QMzVwmE/ibTHBr0VFI9HUGmLfh
y0Fa7aEdMKMwt28rQO7pM/SMJpkUCTON3sqZzVOaw3W/Ixr8i0KKdMriAgaSApZafRPnb6ORS6wR
BEda60VuqtRLwbhqt0zQlEJdQeFeJptA+Bl5bOnIq7taIFTzwB6qXnwBedMhb/bChv94suUoGoyZ
51LMXu4XEqhvUZXaby5tUHnao7vd4tDx/UoVwYujsww0OnVLWJeJK5GyATo8opOhNYct5U82zyAh
TpIqIqUGMuUFPWUPw1mnqoNBoVbbyTOYUNmKwYc/i+95Ygk+h2XhTLHbnni0+m2SFmWRKwJrbgRZ
iUwX+C2pV46L1Y1Vemh8Smylfo31HkD2l9mYEKauy7HihOdFupqQ6iNCMPv6K0pgtummd7gIz1tH
1bwTxmqbZbe8lMdZg9GdViJflRQmVVaNtB5+TtjOUrCEEvlgCJvzBims8YIZI3oOoIiOHA2+VW/A
+b+fBaA3qwEJtCRhAMhRhFdbEK6ROtfSGIFXbbCnzqEd1a/0CqkLnZk8pV20PLoAB/oVvxF1y95U
N62HS20Isisp+eRES3qYx7lKWx8G6IGTro2ZGtQ5hp7HYVpYCXB87bdhWr7qgHv/X0CI9OHXlrYi
lgUIL8GBjOzdnhMlF/ZeXVLo29816e5qv840l1y4IPAQQFxotH8VTWUKYDzmtgkMpvaoNOzoUQgO
6apVdS5mnECMe36na7mhn/nGEvdeN4dyy7hCPt1eKOUm3qT+yQWS0K4saHdJ9p3vHA9d2aPBMlc6
v7MIN2bQrxzwbhxNV5sypjTLI9NduGCQ03hVIaVcjdG3vztXIGmdNMFMC92IZ2W+HJCQJlVfko5v
Wt3TDAWTwIWXRxmYKWI8SMnjJdJJyJv+bcdrxWGZXlo8/aqIwRulIb3ObpJ2/JIAC9twhAtWPYgO
jRyuBMusWCfirJw1MJCEDSx7tsQRTGSmpdd5UJ2VQAVP8AQZAPlQkxTzlLWkeBi56Hmb6POjHasI
WiFfNWZI+QsKd2aTTQFiCbk6ZWocw6bmpff0ToJTOjI0kZqd+W7k2CucfQfcNf13nBbS4sd2wO8y
CsXypmNikwEYO2MuN0nU3u0UPLprLrUWwTS+gSd4ZPjrfoSgw18JVo1ROUfSZVg1KdCj00+vc9bx
QSkg6jNvcFC8wyngkD7CI8Bzm5tiSe2vR27kxVfVKQljp7RLfsHQcGrPLTIqF7FVVqM5Qc2kh8yd
gLoHuv8QSqwrjdS628JucQ9ScMbVb2ftUw94vM+8cnhIuc3FvedLwCMXsDpakSJEb7w6qyE4LZk4
ez4VT+nO5Fyd66u7LjIDFMS75r5v64DwgOdVagJ75+pTIDhkoKB57EVk75v98HtSB83RhYcDbpvk
H4feAMwwcI7roq3cIoPigty39HeY5QPt7rnPCf8aM/yCum2kfjs0BdIwiMLfiZa1tS52DU5apBub
tDH2SSur1sfK3wJBbore8KSSUdAtIoohaL5eOJghvD++Xxtu27IZJzrgF52aboI2WnLUvnQwnv0Y
zjrqcHAhR1/4nZsjLpxkZYFU6fct0i5LZTzyNmKX8eJ4Q0mhCBDhN702rSmGXatPIIrwDFa8n6g5
nuwdVk0DZPSHoRAjn45CTwG5p4OU+ZRmOQAku99MKje1KKFWQkt8v2UQGucl243GdcmxLD1Kza1Q
C3JwlYg5dR/BfBAx48sfSjznZFkdm4QnFCHbSCF+9NS9Hu05m7vmJL3BBezhktoDuzW2eUG7uOgz
fL9Rt02ctON0EEnuDTLMy30N60hMzeaw8gopwLvm6qfE1Q/2Rlc5KbbSoIk21x1lX9Q4V08dHhLa
jf6N6TSuUXwLNjitm4FsG0HbtR/LRyMtzYrqFrZYtx2EL3+PQki8g82QK44xVcjsItFG6XsOXNwF
mNNdh+ETyQtWXv0VgPup9a9CH1awwEdCqGmUA+nF5TQ7YhzjuD96ScyA3qRHgh+561RGYE9cbO/c
5DBy6RtQGB+uugFEqEUvjt+B6ixBhc2nAgSarS3NcBCK8JHRUZHOhFKwz/XAfAgfdd3Y20SSnymM
d54nDAgd4w++1NISGr01uaqs/PpmagABCW4dPTrRlYjLfG6BuCmW+ZamKADWZ1YfijDlpLlSiUtz
2XZ2ru5Xtm192f2T/zUNOsleWPMWDEcoFDm3DGFslQ3d9+/8EkdB9Uvr+GC75YUlPIqnpXiBZROq
oQ0FKZ5FH/nEIXMY0uVjOnHbOE9f3n8zdsZsQItEiAYRnYo6M3mdJoUQSeFQBHixHgNLAmknYCQ3
R++JdwuoFrer/vtSeu2FlgOAiBAV4BMGO8whk58HoA536MT64gb4SgK6zhHxIlUi5rcAQVA0rIpJ
v1bHjbItw9bYBQN1/07z0gM4j4/hb7pHrMMqz9RSlt209PbgGRDxzwMuzjlojHpXMfihMtcB1TVk
415pCOuKccowyvhuRW8GXgtYyPyS3OX+UtORCs17QVxQ6p2nr/OpU/Q6qhTgik90m7YFINY8P/aB
esCx531CIazhyuT51iSGzCsUfI9pzNmlWCalNr5dptMGp8X7JjQV6UyK+uq2Q1pJb50OTt8zeTK6
5295csy7sv+OR0aE5jyaoUB88FHrxzSckUpCsh1wEr4UPIVUuLvoY5xnIs9+e2+h//tTT8pTbu3M
xYKXesWyfHXpT1YncG8fBITT2Msrb2GqsakU1AoS5zpbW2wHYZfyjRvoEaX/1eKijiQsYWmlVbQp
9+/Fuml2iNRMkiE7Vk5K+wBvHNrvubcSJSMcEUTANsaglaOELF0zVOcbjccICEHwIW4lI0eq/GQF
FtEhF7AkBAcG85aH1yglIy42wm21lXmH6dxax/ywadwLMkt3GISF+nNH4mRiN2qqpJBISxpG4HFA
/uKMZwmrrVyGk3RvQYV7oTjUdrSFaUhHp/s1X18hd4XYOn9NieRrAZbbtm8Rxgz5v3cMzevW2oEN
S2sIoc+5ntPgX+snFpUFHRt9Y9SB3Ni95xsgtTeZ11+/lyNxiF/ZeGLkIj2mR7lANp6PO3rYhfTg
AWAlQs2B8vYvFpW3m58RB83gkQrBTrROS0t2vluiXv8Swmz1JpnVICEt71OKdX4gofSKqsHvlCOT
iVKsDAaFHLmlfqKX+ZOaE5r9jVlf9fWzXQAylojylrPRflfBX2wO6L38yjAQ1pL9D6ablrFbDlN3
C2JoMdzCB2tZ0aS99libQtuqnnA36Fz4JO3Ja41dwDvOq9fHEwDLcoknMz8qY8qqt7YASHxvGrvO
cfJ/So9+pV8gcIRTn+se2fnKS1d/1Xs2IYDyibfDYmya7gpKW4Nrz5jgQJKPuw9iyhEsfhTRtxAs
UItEK7dQqx3fl1447GP/uWz3JdwKza7dvZRepyEsN9ZCJsVlliX6lVvE3mMrq13YXaqmCJc2hIu9
dZnID5A5afceXGSTesiXl8t7ybC9r6ybMoCyJ6sWHZ/yfMLqGMbl8YFKMCekxRTPmUwelqu2zgoS
2L8/+hzszpm6KwhC5xZl+ellUwfxcwdobFz51JSkUiF6YxXDjGORSAWlsSFuvTzE5CD8NR9UJs1W
66P+SsdstOcTp2P321slua5xiULw3CFFxr0XjVrNnW7rEXcKkfqimN+XLWu/iNr6bYNW9kAPjkxN
v08TO2+xePjCC6SPVGV7pBKtH8FB7iQ0VCwP/b7fYMvEub3+8ZlZX0VmhRLNc8apgJL4M14fP2Kg
4drISC0VPXrxL6mFvoz390lys1HNwVB4yBO3LqTihy5OWqhTG1xQuIPtmy3IVzFRHrNB02514T26
4aMbnI9Q19eYUY5UY6bCvxdzIZVsXJmbrpgTb/9PSbLzvpEkEe8r4WqUR93mvzDa/OUz1fw2fP4J
wKYXZ5hfGHJKyDNOqF19O20EgFx2taK+rc13UpJT85JXykSJc/rwmxXZ2hCTQwu7G/et/nQvGXNK
ESXA5RNC2UnI7+Od0z5m0y1ap9g7CuB6/rI2in67fxDP/hBjVrJzAY/ywEbWO+3brK7BP5vo95eM
YRJHz3G0lrkxUNUTHPp8/yEPgiNcR3EY4HwTrvR0ek9FwC344+PNPlLE1wmKR7eVcna3/ir9xBa2
EthpY7FFrOZpOY1CsCuCkWa+IqPWduS8SSB5kZwWJQmvfxr/dn8h7/Pv03LsQWuwerTPoZ0xkeO9
xmVy3TwlZIdWMK+THBQn42MFV9DYdZ+n9J4J8V63zmYbV1ImCeEiPYODnhT7hYWFiPP96IMTGZs4
gl6elr05PDOY7CdsNVTVTb3Y6fAjtA2G33Q7jaQuAGnvGf/FWHTwQ5NN0HmaPM8bMCJdbuqunW7H
6TUfPfmG5TfnjKn1GUDByeF6KU+9O1MlnWRBT1YmFtYcpistKyTpfQ7ZL90f/8p1gLl7uzqA1E9q
E/twr3bdn7CTG13wC/on3LaBqjFzX48+GDDeowV/n5BbJ+SwvG36lgsLoiWYbY1CUymc3Q76CK4T
/cj7sbMavRcFuZuI9x6f78hzRCKmhpwK8i2qcnt+D5Mgz87uk0IWX/Xk1yUqlDJXR0mEiAVsPH2h
93Aw2E3XLwd43HPf+YPWDKdlRa+b3eNFeP8muL/rAh61uttwvNeQVmf+I8L7MsRGRGwN+yzNPERO
NQUNSv5utwuqNpYA/aNi0dWltTGlGeqVvpzFTNMADvSkAOM4pntQDtIuzZ7Mro/cHDyxhCN2gKUQ
b1vpCeF3568Bv5fzKiLza7FjM9sy/fL6cpJdgIehyk/qoEduio8hJ/vYuoO2/mc+juECUtkQWca/
X1GI7gJiAgDrA/vF+ZwlXVL1O5WKRNTAxR7AL9ywoignHOuRNA5ixLUpBULVE2pdPSoWvh8Z8Hot
zIBqnRNCZWa0nof1CIKxR3OW3EuYCowPeCPeKJUyBNBIZou2GFi+u9eQb2mdzbXEnpgy7I+eUVht
gOuhkdaBsKwJBYoc9MRXRrxW0XwyNs7obNOUCPI8wT6kOq3kZQugay04ANZMxKBNGLG8TYDxBhlj
dXUQkQWq8m7GIxUSkZWx3F68/j31KOcSGT1s79vccxgRKFr1sgYepQxYWzAdA4s1Ooca1TOPfvRz
rMoy1l82nNIYJsquWY/wibJZXWx1M6Z/0R9UUkZX/NZwkr7IGziyO3IoV2pVzaGPy9PuCWvhqg9H
fZ3zX1NBQeNvqR2ViDEOdXVS6PAJQRT28cTS2VbKKXl7ee0QXuiC8hSjAkGGdwGeemXv6aQ53JLw
btHDwT/owdrkveBzg78bPTn4EIQoA1i2KzJnEsmigZJDnrSjFKx312gtj7K5qGqUG9utkNPOdNRA
O5LaGFhSg2T55nsFpDWbUY4jEcjxR2Fmt8v5atUfB85M7K284Si+ynUQABUbztlurmvxB00RXKsH
dIUut5AnJUwSxWrBzuxPq8UImFqV78Cz2LL4x51FuVZ2QKuyKzG2PXOxHqR5E3U5jj85QrilfcIM
PVLehR+mxIfTsvhiCMNIcfc8MpSIuFG55r4TG14nSYGnQmGY3sfynInSxCTQco/ZEP3aIu4kQ0Jh
rhiBNTVL+8QsN6M0a0IZZm5iGguYeD2SPo44P6y84YfItwFdJdUdb4++v/cSEZWng6/vTKokcyZ1
VVH8QBeD5UWaV0goMCPeLkIOFc7Avnv0mWcAxMOdjz45xUlsVHlkR4jM2xt33ajts9AM3URMmZn0
7CmT62ixo1lQV20IbI7kNLG3Z81jeUowwGM8ta7qRV1vEK5HrZJnT0tKVbvh3Pva0nhQ427MQqXJ
Yd9rJaNERjYVf1mwLbBja5GMPYMBtZRCRjPzQUub5Kvs0cmcEire/t4blcfDwgujDLAwVHVB5ejN
W1RSbi7GQQVLLWtx/D7iBDxREMKrR9AUNve3edgn3a3PYNwUIHGddyRWmABNiMe1a8LGeonMRKQ3
wrg4ZmVM8HoAq83FxNx9rJVZAfaRcIlwBiCHFjQfZIlSMfzl5lEx5U9H1jBkEm2jMaJYS8m5cXi/
OvOvDse9bCZMEP+fVISHDUMCtwpH0QOsjoTLD7s2u8AfPGweLRCqtscd2kd9cDqWMho6q2iJoiWI
OT7LWEqwz9sGvYCbvx2fcETuc6WGJIDhJyY4AkLBSFUzM/asiXRCeU/+S6kqjdPLXBxocttzEhDA
6KBrDroLM1NvFbhthW1avQcJp9UxSvD47jBmwbuLe5hmqUwJ/IMJX7UAj27KFYRwTmrC1JGR3fZE
zrrahUf1bRiyj8whO8fJkg+Grdd1aNd01WJ/VcAKGUPtVZguIL3l9sh4tpOX1P6hfbKC3HhhatTz
m7nyajO1m4qnC/emWs5YMnPTwNtalF9LPmJwe4GTWlQb6vbU3M5y3THra+0leIlIeg6x9dhDxr5Q
Is4HUOOkd28GW0zU6T7ViurZKgMaVBBo4ltvPcQiVtSrojREXudk7rgKRvofCzvVYh9szS5nVihT
tZ71Ft0TBh7nnIWME2GmYXDiB2t8XavEggJCemeCO/K7epMRkr/CcrboBRJoWFgmREsbfUH6SCsn
dMXN8OHUAVfPC7BKDkSCmexhqkz+ZWDHMSWLp8xNl1pz82haAO7+cBEng7LeumtPRderBA9w697r
1snvPXAvc5KYQw4f3snRxLZV9fLv+4nuyJDLqQGTEpiq6Ekn0bV6oo0L38XYNiL4VZqp8h9GiiLM
/IIb17g2nZNPibMzP4JSrfwr28nXNKL5vqHcG1+Wsxsu7VFS7qUnFix+Xx6NrRZENqMNUlsdFsZw
5sz0IdiW10DstxfvK/eN3xKcMosYS1+oGp8+gNnqBkiiSR+U6UOuKqG5hfd9NYzouvH5Ed/0QZjC
0HbBqLE4+GR681sLJjDMI8rXujqiHeByElLQ+dtIp+YwaOpMZKR/zxr4YCq8m/dLfNOd3tB+CudJ
ndd8vnsaI3U2SnKOfYz2E/UmlWfDkljoPXLCrrgzKxQ/HW8+5s/QGxSVtnK6iJsjP76OOckzxoLF
XB7lu6JdOmM7hrcL0AoB19D4K5IoM4aVrYbwKAz1mW0TMN4SwBmyAymdyUF7ciNBOxV332z7SQXA
giD2s6zt2hyXu4Id/TQpiEibSzFcR3Tol8julbXUhx3ZTvi6rLF4znQjwzIgShC3fUawE9VM43j2
RbhHnoNh7xFqqPOV37dA2TofTK+fNKbmcca32D248dyyH8MS8+QpLH+OZodH56OZCyCYIRWOjPeW
EIoTBRhypstbc7eDNv2qm4oihAtvQzidsuPUw/FtZu3qKfVPjXBz3JembtnTImMBc/5DcUB/hOok
v0sjTHwYH7WNlpdCFHVKVaMyr76j+kM/1YICdKj0pYEdTGV6S1wMXzujSJpX+EIlJlR01D/6hvAn
v3T5Y06KjJ8Q7QUVieqZLZnTy4NsGTq1/GqBVJBRFAP79rGVuYJc+9iiVLcKLyYhU2xl/BUmQ8CF
XPHH2HWnb+NRDWDGb8jhkrXm0LjFFsJ+tT2pCvYywgairG+Y+yIbtBIjsB0OD5CPd1qJg8Ff5RGL
D5+jYE+e8ARylKojl1C9Cs2LCORNwlPrzXwAFo5z7Za4vm3wU7dmIMR28WGwU4c4xsFIBtGzhbDN
oLNvyKEeerEbWuh8QsWfa2A6wM0mD2zm+AhcEEBqhpf4lERs6gu6Amv46/9Q+I105OHnDuWlZxnH
t5NwQgJJjFHytik6nkz0PvlvaRgRu/d7XPUQO0fLJsBw2fVNYfgbZyCs8zPimqpu+0BKhM9KZx5V
C/PlUT040d1G5OR5zYHP/aLSfXOHCQ6guoHQkxofk7KxHlTGJi3o4uacf768BBU9y4OYW5p8Y/y2
nMpw1+SIfpmajTsf9/GPtg5fmQ5Rn5IKHbAMaH3KRWj3cCPERFvsbMXyjQ13h79jvxrKJsxQVaM0
EpHUXVbKF6N81y3ogOyo0RJlockLKa4mV9PRnq52NxXBWfdZKZmek7JwPN4BQYBd6hNmEyh/wc6L
l7ip4Tj+29+qh53Hrd4Db4WhrgUz5kSu+j9lqnxV8X8sAf9VbeA2s5rpNphxOag1e7ZBy31aeED0
MNlcidDxLlSY7TAZCsuvhJNJrmaSNqNy2gQ36yQ7DAa4OaK1JpgOHMvp4JH2fIM1eZqN/9tcGS0M
7PTkVa5ZE/oG/EB9Z0pYrU/FxkOqG/cCJOzWf7IbsVf7Jggc9og+7Euws3bSMFq8bfBcP7xt6I1Z
2f/MCr3gyfPAp4XvCZAI1EjePbICa3UxbumcrGY8sL8ymb4J4YYKb8YxSnFewDYIKtitgvboegJc
xWpclVzsdBKt+L6NdVLE5Uz4A8mJi6eCIBQVBiHOZxxbpQD/BFkFVweFDQ6zyvTi9GZxqZf1TMK4
GD0y9FWhnno+AlyM7tW3B6Mam3erijFGThcmcm3EC74RbcCYdXgZszY+uUOvqL7HCMJRfsgc+L06
mhVDpaaAGNSVlRWlb70kAzkeXZOhBMjYFTxHMkHA8B9eJTgJccIm2zwau/vtBOY0ReR9ZIB1RX0/
SkQaNb5wxn89o+n/VFbeN/blV8fK5aKfLvAiCemWgHCJg9fF5A1TmmyXWTPJH9T4c/c6tta9W+IM
7tDtv30aD2ii09NSE7r65j2hDPUssn4WTVkg1Q17ONqX0D94SIaDm/5TSZgL5786Cjwv4Qtq71wk
NByycctIwWapWmcnjj57gZzM8ZY4vzoBdnI+TL16aKTFvpnh9AlasLTiGTljrQN9CmxM59+2GxfF
JY0rMhwZPQbXZMxYU4CD0v3NhQeVRhOxyKovc4EXPK1mSmm+iFlAPRmkTFSoPvEi2UigQQwPnfPT
GliORl73jMsWOErs5HQl7IjtX3TdwVzZODN+LyQ6loZqgT13JY2EAytmUsZxmBD/rY/ptUELY3z4
qQza2LuTOhw6U5Mgn6zF29ZJ8v0d0N1Obx5f2dr4iQdI1xoOnC1RkJl4SD0IXjLs975auxNhumaa
rCY9/s1P/aCyy2fQ5sh1H5LCmfGCYEnml3h6rW9NOCiVXxDCQddXUdDWxphEfFi1EqLILWMwMeys
57duJrdF3W1yABeb/GJcUP+2bvIJUYekPfafB3qvcJRP9Z3rRMPzcYPC9Y0b3NqVEswCofPnL2oW
iW0uREkGr/BgMGxXA46dH1tg7MEs1p+FeH9waoDr+QojGMwt2AGhjF64LThVnoAMN8o4/Avmlw6K
dHMlTG/McBprufa0VlvBkHZNdg/6kRLt+ExnbfFH3MPqzy1TblrISKMUppfWSYTKzJCx3Knr4blF
EZI8xkkmEX2Vs9hchsbJB5WWziwHVtFUIdZHL0z6Vm/4qqB4wPp5lWJNYVv2thaVVYoaBZEOQ2c2
+G8EFjgofiZ81/F6lcC2V429iiA+a6219Htcap+eH9hhkHfU3N9uLdFACiLSpfmVuY1PmkGgsbcU
HlekapE7R1z+F5b+MFDzxPnuBfvLr2P99ko8Em1XY1Ts4L2TiDcUts4Uij6KztoOkFipXkx7TR3k
RHwsCQwWevWkM62FfUxLeFLQqXfjPHJoWn4Pt/rvFJP/DG+pRjOp76lwgKOwRHvcuoKvZeCGWr85
kXtLLgicE60pHNlUloqtnSHIIZh+6YoKhIANwbymS8ZdftvWXF2qQu/ze+vvBOgFpKbKZP8MJ89V
hdMd0jiOfUKLGfgeMXlsMh/h3TK82kl/xKMcOhwQ39Ygz32JaKL9CWGtwTLhTv+WfcMF0szvrEom
52R0qnDX+86Y5W3jNwoH+th8Y3yHl/yFiz/8X45dRo93Yg8JCm0QiV+td+C30BexjDa/RiRabDPA
bhAHmJSnMZXcRrwOSpsd5r510UY/4LgyXChkeawUcwA6YKVMVQA/r7gW0LQdG7Lx4mD9j5rU7n8u
YPB8LdqrZ+d3ifOyzL/IRiPjb+Z8FwMx/bDG9+UsHIewfF7vW9GmpvXon7OAg0ibuwU6mqf5USRK
CiNH1uuixeZVR04pT6kufXgvcAuAOxSj+2NcwZQRZe3ev7cDGcuphN66TDPt7jqTaW0fUtKE+m9a
C2voiiCE3FUJ68mpjnhrPxtvhHqzaxu9uL8ynAmKr4A710fiMFA1hSIYmaMqfJsUEy3yveYcjGqa
V23EJbGQG2sopuA7L4kbNuTF1Pmk5JC1fxJBO5ZLn8BImK0KtIyckutjAMmCI3qITlvAAIBranHV
zg56AIy12Pbk6cu7D/ktpVPGPwNJn1p+Q9Jxa6wQw2WT8vY0HgBHpIJnWdAF+xM1QZ8IBkswUAtX
TD7zSRxGmOEMmHtiLqjwdmFqKyJchqNfUGtqZJU/ZFKli6kJmmZ7o28r/WXNNdtmFMUreuxxTh0j
fsMH6rGPJl27UCuGN1+MOKSHrms33B1IQnRWa1AnNLAhgDGnyhMph67nYXjoZYAtEtL45zYSr9Sb
CzdPuC/zQgVOwiepwX1Wa6JyCEJ09fqwmnqi+WQgyBuBM5hPAxV3EFIK6Yr4bXNIkEbKI6MD74oh
v4sqt/o8m3bK1yV1ACSFiC2Sd963+HTyJeT3IIK0zFfCWKIbOIG7OVIES9SQkYPzixNLwcpgb+xx
57uEUuIQLDiVbhoifcXjYxWgJT/rzHjNR08dupFlsZCZQdgbAlcD3TH7WLUJlJL/jup9/3bBaN4z
Cqby5RDW+RF9dXlfQJET8WswdcG8CAfISHVkTCksb+oct/6HT3CSsG00uEMobIE4nTaFrmhzHE2t
2iu7M5S88KVzg9jtrA4oUeF7FOr58yXV2XXjezV8EK5PZy+nm8gIY5rXtXto3ICHOeQhFf1ErYna
OeO0LjWBTWHcspHr+L0aGF1DvVHtaGM7n8T4P/qfmrOK4NrqTJEq/OQRcg0kz0awN+lysaq3VuOb
ffpUiUO5NfAUylxqHN8E8rP7TAEd7P14R8rhNhqqqKHz5Ffe6VXU3pI7HKBF41RyBufU/28zY+EM
TyGCqEqP0At3dJ9+aayNzMirToReb0NbTx82vdcif59EDnTCsxd1Of4JoJtD3Zy5isDf+old3m8d
PQIMGcfScBVidMP9TMHqxViENTh/z8pxXuImoPkHdcExhLutMXiZQMO4YLpvf0n95VKXVAMrHWy7
Rfxav4yz0QYqmqJmmamD8ZtMAjD0doJ1BEN9ZZj3nyQ6pE3e25K9+p8O8ckLUTySPCBQaTfJp6vB
YEVylejQ6Giz+QDD0k5aJF+kW2d2FsXt4sbV+pxbBFEdNamG4xF8RBt9ysb9RaxgFuGWQ57C59xX
VWJdmUKtpaa9E6070rag1kXoKCLjXnTlLAeew28dsS3tTewAFjc/nX8AOmEnHJj2ULBsFMSxHVeO
FvB9P5y1JlDKu9KeDEb5PsPaOO4+KC04RljzXXLi+YNMNdGUjfUCZy1F6CJbKNXLA5ED+s90YKRU
0Otjy6F7vUXcKmhsB7i0qePnfJIOAfIK4gJ/juB7n3fyrZ+JMhcI8SWpt3J1J69iZOW9rKl5JxN2
ewKY1fWBHx+XVGkShBJ6DOvJubJ/R30SCEj9Xt1h2Dzf3bOhVyAJEVjS1VFA5uoBdb65yBhynLFC
7/2tJrYJdH3hlCSZ6tgDUVOjd4RPsB1y9NLBZ4r41uWdy8/t1lwaRBIwauazbzanBw9xCdpC+XLk
OC/hKuRnibRQmPY7hnOoz5788WYotQdyMcWnMajAQeJOCqjM+Zdi++odXbmNq3nC+BxZzgUpAhTk
6Jnp8AyJ41QkQzJtgfeCaJt0qVsKRGxkEBgjlecHIw3wl48ZZWZ0aoyvPWD8MfQ4y//mnx0yqXon
IRMRPvwH+kgNmZ5ZWB2ZSUzee5eiHKG767HL4ZK38E17GMMbMx7fMeCI8s7ZYhNDO5E3vplvhF/N
OkBCvNoUUuCLWAKfgNQXZAjf80BiaxfwB83aTKvo2UKUlra7rj5tG5uTOtW+NRWjuGPXoqtQ57iU
Cy9T4k8yx1a3VqGI8Dipvl962ilkWNhTzX0CxE7/EbcmJOs0T8g43Ev2Hk5ZpKw1HtkifuyQrVeZ
Sfjrp5qgT2IMq3PPjWRhX0zGQTrRWu1Y5wPzK84zilcWJ8fsjOMB0s3eWe/O41iFq1o76MpJ/dBJ
sfPs87CbbAzZgKbv5UCBtr4KvdXPQtdrxmCWnUeSu5/23tKa0/yj0SRABvg0QdJkqC0lFkyxk0BL
6S13NWOG6fQ+C9clVgtMbcLPF67B/8ZEz0r+JaCssv+Wk5klSCE/aNzEnvo78jENOSjgeMIKo/PM
PM3fwF/wbEqebqZ+7yjzkHrVbTBEeBT2/kP+Nyz4ZpHPUpQi8rONJNgn/+VvhTdDt05y8BS9jukT
EwBUJJDbCaSE/RT4NkyRuFVjSDtNPRPClhXDnfoIk5ymUJNUlhy8/dHLHkPHMx4M/gKr/CiH5gAF
6/CxqNyaqnqx4ezpsfg0BzHs8EH0aLO1xdev5JVdxH4DryF2pY/gWIwebtabq27VbmYe39mBFrEY
Rn7bqjqbsIPi0ODomTT+u43IdKsdhMBvsTWSl3kfj+pV5gLHgoEPoQGSnS9+4DOqKEV0BqHgWim/
40MqrH8w1W+gAs1R3StunLRZBT/RpfERzMpf75mgA7y8rLdiHBNGOjIH8lK5cjJfFI7jEIJIUtqH
JJE2qYKz0DrjUMM/GMl2tE0KcN227Qfv4jLvuCJjEW1ULRaMsFYfgGvfVdj2ZNCrLIrj2buX1WL8
M3y0u6BxNlzH9G7OO7By6WpTCA/u6hU2ZsjGMn9bEY4WvnU9sRtipoDTmvNuv3U2iCfDqwFnPxkV
q8F/OsAnME7cLZ5pTCR9eXFCTVjRRvM5+TcIIHbQ0r7rA45YpNuXzDomzmToECCXJrCfCzMfUsDR
j3QtETz9JgBqpmVd2Mmj9ccfWGxtzxbdbgTCQ6ubo6U0c3dh370lUl9VJ9/U1g4gxJd0bMLhvNON
xUzc9CzBMMdjTbp5RyxbUvDtiJrfcRv2MKNQB0uJ/LNQsVpRKIZu5iEPxney69kzPrdTeLNtbtp3
NDGruXN6wPNFOwDXiU0jHTe138mdNht8S/nJ/+kmMpGsUhWssyB3sno+vwW0soXaSyd08PEDy9OA
gGWLYlTqpXWymqMd0BtSSp89IsctKfSwa/03emTwG0b3nlxJRqOL7RJxiamuPfLs2ZkidQ3QMvJX
xGvCQtEp0cuXoBTlxGu8ulMzuX3hIIss6BzIpuTkWJoER+Viv1PJf77JCOnGnImAjdEY3IAAm/Jd
+Zx/CPzPNtGRHZirZsu5jHe13lQQcl1OyNp9X5Dc6t6Eg1sy5/1qXT+Cf/DSJ0ozyfml9PwvVMwl
slAPgSiROUNvaVtWAzNsDhMVsHfN+YGs4Zx/i7UxUP5EIqVwl+XeZpYwlFnNeROKKoqjacSEmp0Q
76puSn0Q4+6xsmJ1U5R2zFIeQLIfVULQOTzNshsTkEDm5rO/qOGm4IPNoh5Pyp9WdgxnWIdu1slT
WJ5XY7OUaDnIwKFPg3aaTf/mWQBvDvH0zgOLQZkaufHU3f9P1hsooxdkjRiYLmPt/895KU/C0xkK
HAq7bFxW0gnLIH3QWvn3uE3TNGKAL8DOzV0FtJfqHCQFZ9Q/U16mHyop9dsqAMGuPXrVLzkmEFmW
F/KBvlhNjy5SaPnUweY+kd/J/O5iDAZ7HS3u0ILDI66SUlyRNPUQME9wLQsh7CmCRQy68PL0tcfi
dH/3ycDN8zdDVSexeFRHspqDH43Z4/xhwdED091xKtDtFkhrigvIpyMvMHBywFbUkS/XkHx4DMGN
cxD3ZMmODkvpO1Eg1moF/jQfZ7XwaOqTwOSdOhjx/2jkL3tW5C4I91Fms/DhLkehu73Qh6lNNq+1
KSjDZyfLxbuMAL3LCn1IMLuRWVl+Gy11YyK+WG30Lo0VhnsEp2Oiu7gRgPv79rauzC+QRcWwL9nv
ifHZdEkLbw2FyAmfGecjDeAusHl4NznoefAMPMpMgMSM+RM+zKWuUkv8a97XKivM8FyP7Bco4dRP
/IVBBbN5JyyAm9+f14UFU76f9r6Gbv/aJv6wS1WBkrbjuL2qJJPitaC90yxH2VclCtZ06gyhq0tm
BZKc7k+s5fy5OzniZL6sQFjVCMFN9RZWPEVbi+4IG/MRZ3SOVeknA9upVdyC8QjSP+sXw0YuBpRm
OzPHWU7mwRR+qe5l/SqlLbqw07EMd1PK8v7erhLdLFg23mmIvLLPKpvChmRLc3uLCyzcsOuA9Kxj
ZorH/UXkyykOhSA4scfiSF/iCyol45pskirC5Vwa1qR/e/gqAw6rqfBSuKR3ZaWB1O3I3OwqPKjv
aWvy0QSqqIq24XzKyvBfvqKkeOdzHA5+cgMRhn9dgElLYcP+ukcAgjNUw7llGnenNtlJrwq4YmBX
7rwmHoz3Thf8H42io/F+bF+6dD+qHfiIOfzogq6z4enZzuDvl8bEnU7XRFNywoOHjtD1FxYYjCrB
um4eIALdeNvuU9wXG+Q2UNj/Lt4JfPw5tr1XY1NxPzt4dmKa4ftQ/eUGTTid7mGCGu2+Ihkp+mPo
kckloEQcQ06A5pIu4wlUzj6D1fEqDOKOXDdC1mWxzF2v66cPr+OPcN5VJHAnPnw5t2Fl6VJ2xlpa
MTpTk+koPbrAHglhCFWp6h2WvXq2A6uYB3y4HdMhGVEiAg4wRKTzMnMKncV/qAlPUatGE2d4bgvq
6plSKaGOTrwV/1Lez76cxx2NuBBJwJL6lnzPcOHmmBwEvNHflpv0zb43rPJOJi8mD1bNAW/hwa+e
QL7b5wNoJJ41tHB9ys095qTxWvqoCmUQRcRMuF6+Ln7oJ7XHGHvdzwv1cctoq3FsriYXOLMKyaQn
yEI0N0cEFdbQmPAZWWyHg8WwDd0VfZ9oYIXbMghmxZv7Ptm0wcaDaKLiyXiSGP45mf/5puzXpGP4
5trYGJrHcjOAqKlK1ppNJG2WSO0BvJfCX3NMZdxjrDDQ4i//iVChbLHNJJYIAKgfyml/fIkNWx/B
3kQFGr1GwRD6UmxmdDevE3OvCB16sSALvJUgcVog12LHUY8IfPwpo6Uu7inx0WP0ph1twJ+Z+7+6
YAZUY+Ii/1l5RMo+MXgAZwLjgTuSD5WE1oDNqqErIAbpgHkUtS2MizaJKF8NYjv1RraeIoFO8Mic
U7K8bJJwDA32Sr3IRB66RUuGiQ7EZpZ1IKZcIomUdR2H6z18LRfkU3amMMVA4tCNlt+4pZvaw6tM
IWKJ/Bkd4MId2MI0mMSTsdUkbglngRYb75MDF3EFejvGUuLu04mz+YMaxpXMmzYAAdGom4PBcWVT
LSq/0WdH90mqcW4JDBxPJBpBsFfR0Kr2nMIZ8iW/ruCFXl9665ms6HMm5u3Yt6KAu8rL5TnT/u7u
+LSM6UwNZU3ZU8NDozXV4fDqJ+I2v3Z4/eshhPaaDWWMks+8+SwXGCeCirVU11+JhKsPB51Whs8q
Q7gp/jEH/VzzrhttM0PNTslZDTfUnnPakx6ZVJnMspSe9nRbCijl09Yl9ASjG+DkdRuX4M1rDzvn
iiSM+LvDk0cxvOewPlSe514f0lipLe+4rLuxjLdXjPD20Z2IBp8uB6PLeK9PTOWj2tfFCr5k0AWA
yeyg5kH17WiCZYJbk7KHMJCrmYe6NMGvFQOUq7V0G0Eqi2TChC5omeZi2EFUEAXc1hu030++r+A+
rNoHawdBvbgiODDo/Ao8DqM/sEE/yacXXQp92ttehRA+UDWDN9Rg7TDeHciiZMcvZ5NXkfLeN/0B
cg9qZHqkdm9GhO1OIvJjcXpKi5O1mswefWG1ZsUSzkp7GOiSR+QxNUV7UIhDUkLu1AM/QKqfYMJr
GuxvrT06tnJXsZd6QkbKzoIselXrKKN5C5KyJu1IVcXy8XOJ7ZQbxFWIXX6WIav8AwVaukGtk8he
eHpkxTUTQyh1Bwhv6/AXTbpB94unGNiIceaOPivRBaJQ7ig7a+CtuFJGFwXRKV9Lf2cxOElgR6lC
kXsY70tXD6zF7I1nRLSsFQH0pcVP5eVStKV84Xi21GBYPBe9npxvk/TSUfclvmuXjYGgJkIv7CTN
iV5NP8ZnJmE5fVUL7vqKtvvRldLC7KsCcS8FAJY68CGUDh4/AiZJ6F55mWJYLbpWE/RfeQqAi/8J
pnzqVBMLuq6dNxOdKDLLM1vrJFzSlHjokFphFgzWowA7DtHmuROE8ih77Ow9qSxiPalXYmVlfWEK
9tWvxuPEtZVlTd8XdrNNQ6IGQsqDAG/BklTe0b9TeuFL2ftTUjCdThjSRHgRfpNW9+X21F72BNNX
jTR+vFw6M+cVnNJEIWJInVJWyhgySOAuyuyIyAiSh1/ffwOhwtF+CD7g5Xbkevsws1TlOdcMRnvG
aIOPFfyb+T4J+XWZt0edfPN5c+KtlpbDFduGr6l9irPFbhbd9m6OuGMGz+/Gz1R2kp9uUjbKO95F
4kg+2t/uQ5eea7yPFRPumNBMmbUEvJ2Xh7/KJYmT7dR/Bc1YhqKpEHKBnW/TqoxnAfJZ3qBYYWB6
zs3GeAryXBAm2sT6NF6H6HDH+ZmTnmeMbHSHx1FZsOBGicsT9IFfbnoUcQuOuZs04avIVlqhclda
1/eaAGVYF1XvsFIv0s6tSzmO5YNFY3BqbBESKVYyt/0euqOUgDZEDlkHbbKT/ZvfgijuEWeBPdaW
w7ZkAJLkpUorHJSMlqDWtImoJQ+vspTXHzvyPd34+gC0rklKAm6zUl+70JLgmZBJeONypzTv1Irx
UK4Qgr9ZF8uFEDBGSqTlDhtUzJlT25LAIDM71GQYVp2zraQFNqIYbTaVY5aauRNJEVasNKpvmvBq
f/H8mN4xEL4lvA69PKbXo9ubdvQpETh9MwpGXvTdEznLP7CwY8fVlKp7o97Cr0t2VkskkKWcQyMi
AB+liC82FWeWXeYgNgvihnQ3mzLjry3qU4SaHL6lm4Qcw7jYL/nM7Sp47mYemO9DXohCA5MzPPMH
zVmlewGIbUeCcsX8sKjdiLs9+RyRXObm3oz2rHLPaZPspke7IOAkf4tX7rpDnD2KmwUirD0wM5uO
FmiBuVzeNhVpQAWEmP4Qr4HKW9e/23x3M8K7U7U88Hgh1++p2pMmHa5hC7xXmLlSON3DINJL5cnb
z1OuEIsL1xXCIDuF6yHRBPPlEi5flthyp9eH8xGxjQ5+Vc7l/SBltgFIGJzGJOOz9PlqJt7o3hRQ
txa1PHzeATt2eFtCfILDNX4bn1Jfls3W9H2Q5jyYDy+OCyQ/3FbOVJ6gnThxtvJtWfSfX/ajhOT4
knvtbzOIZL7wn2FNPiKWUadDR6VF8gwqH9rXGvHKtitSO+sq0B7KYxPYVqTJHAD5qHSMgy7JE8mK
21K+wHtTMFYEJRp0zrAwCVgjym9CwhRpH1aDtdtihml1LTCgiJ+47GgCsABpSoEFoG5IsHrd5oaY
rezCFCzUP7kQfNM0BPPugfNS47mvWTCtXk4a9CF3XpXii/33mvoadAuiCVYZ4NGjVsfp0SIMvY6I
6MgOt7z3PmQ7wuIIEuNpYqoeE/1mEFNjZOkepo5Dvjl4SE/HmWXxteQXceLqWJmXHciyJXCNfeax
FqbUxvi2DwITzsz4VlEXV67XMUxA8P6qjnYLExQrrlMrhKraMevLmJruvqNgch4t+wmq34qZegJ4
TGVTfdWo2cpVnm2lKB8mRnJm6W4D+MCge8wfevGW/xF4CKhbD2yfKeiPXt47bSDOvKkhGWinbEQ+
VjNsujJV0uH1ygKElbQo1H5gnLhrOADi/wQt0Wm2TBXZB3gjmQW2ZCMJboyaOnCjjb13ahmLqgxv
EHHEBAWrpToIySv5WLR6gwkpd5QPX0KKX4lRqaUkV706CrGXJCBY62fJ7842JccEN/9cNGE+R5gu
e8ONzXxuCLWTf+ZenlE/4gGM5GNN3lk6KwkCnvnyL/zQAc135UCS+FpzlqgYlaEiOx/70PS8DLVG
NMRMxGV6uVtnQ0gKopuk/XPytvGOog2z15vcNOsIAVad1+Do4OkHtwRIPnJiGBGblDzfaolk6PVd
wDWjDEhcbveK0fnhZJ96jCxZ6V+MI8/RY7aSWxJwaHZnKm+L0ix9J8zMQ0iEeqCfC0Do4Ks1ytoL
Y/AAZrgnLrICEWyw4bpn0bP9mpe5RkKuI0qrBDnQU0X0URs8+ht3eIJ7Rcr1IRa8lCTCWMUm1CAS
yeF3cAu3kVLfVE8nqSQZoc8ph43SOebX7+pcbhw2/UyipOCDPnWQL1CSlzt0Ry3mtFmP4SCDSHXk
KlVolBUHw7vWhAancbOKTRaG0SkOHr4YYHUsivK3xA8RFPruuvnFEA77LdM+1eB9Si/dx3QxXMnM
fD9IfsJ0krIbH2960m2wW+U2qbL0PJVcmfVhrjxFr104KG7INr6jW/b3TtaG5lHfwFdFpGKj0JoN
vvu4lvQbEiDTTomY6yT15Mm3C3yxshU8LL+dt801uXVlpFQtG9nPy3mbhUZkcX0sximFojasVebN
M51aiUfeKF45CLKKP90uWUaNjtYW1LHBBzkAjvRogCz5VjIVSK1qh8++lG8HzGiHLoPxeHDj2wbk
m/LLoSFk16uWpvFmOuu4EN+c+kFh06TGm88J14OHaEzTmS8k9F8YtwdOCJIBUBd2koB8Hvzu+zQN
HBsvlx5cZgDCG6SmNG6Hc8XnPRQ0CIugiWV36fnO4q7XwQIs/3qB/qS4t/SzaNrbqz2dEJgS+OvU
q5pcx+UcES677cCD1DXrsBJ/nJpytH+4AM4UjrwcBepcbpubYzQVDVfHkuyvQoGlGdzool8ZL4Jk
EQd4X5ziz9wDFhXXhiEJPFa4/fFcd0dfLxzikIJ8Qg3GsE/XEI1UCbVO2AH3ibo2sM8hlFAjN+bn
W5/9/NI9gvu4MNvmBAINCo/rmKxMzmOfkXzFsgumTMXBBs07LpdXGQX3wiD8aM4izINE2OczEdOp
f7jgZcmkdIFr/KMLhkKnGjuYIRAlVuP8OLRSETniYDWdM73RJ8GuF2NpnjmU1Ue2VngnCcwfJVXi
csTpF+xFSTFToNqMyYxJb8huqBxhoeNI+tcjbrYEWSXfVz1jY1WRq2X0Ld8Blnivfqno4B9CLSOj
L86U+RyXWpFKEMU9ttGbkUQiKuJXB9ZKFN412XvkTa8buGEfINmWHbtGFn3/qwaGQL4UWTKATOuU
iTvsEtNta28vt1+KgzCGTbbZXytv0Vn8CvDxBcrzxfhAxLD7Toxf/NfCmsuo2zIDQ/ubz9wGa7Yn
IT+qohkqkpXECBAGJDTs+dw1DKUYyw7iuPZiLr8EunmCvAixKnUQiLn864nXnAH5iUu7utN60yF5
UM+pOcYII2a02POHk8C1AFSLD+PjYxjUAgJR3S09qhy4TzUcEqqgCrJZ2jGt8aazD51x2LV1XQFQ
5qpLItlaLZwMBr7cizv0ol3N1gq3E8YbjiFrv7eQcg3AVK98DMufwrkSX062DtE7MFhK3GYL7sdy
SC0YANu1ZZLFiXlkggBMxilXEbsTeWSH/db9hZofqlA326j1kpeHIm8sEi5apR4B1QPKpH+jai5a
YP1n3Xo3FPsgHhreEbesDtaRFCV6uKkl/knkxObM+a/CAt7mDZYTzThQupxPdj839eRTXSqyscEX
xi57TwytYrN4f8+igxrrWcg8ITmVi259lhR9PTAXt000oO/0PfoprBy3oD7CW4TLmDyAe22CVXol
S0fjP77cKnKNOLkUOI5RVq2NdJmGcefo+Kk6UR7xaQb/l32yKdO3GpFUm5P4iTvLSe30EDDJbwAe
TCXTK1UZRGZoXa7GuPGugIJI5Pae/c0ZbHFaFRNoAE1OQVVPP21cPDjKJ9A0v4DP0BQXop0TzkF4
m+narQjKuEbIo5Y0EavqPwCSg3fwOmweY1nrdySZkf5FeEHjSIK4mSRymjER0xfElu+yrGLxVO3Q
YTmXDeWUXsNORigz9Z/sJPhHERc7vRpYZnZU/jziElBakJA3NfceXIzmDOukCeb1mVkZnULWjb36
NLvpXpoyq+F9Rr6DBLg7tGwVYf7JMFtPGej9ZVh4GIPQg3rQ+FdT2RA8sKJ4jqC7beTynDliChsV
6ODfqfkLsqdpyANtzu7c89Ijh7mruE6wh2M/BVQiWAkiX9nw1CAwx3wJeWiyVHxu1EO1pk3lHXxt
QbNhrYdNaRu92ZTcb93Edpo3dp++vEgPq6RY6dzEJqhIr88I4yn2DeW/a5IDYd8OLQ/t21XvvYqj
QqiGVZuET1jMRHCDWsP6P7Xlwwa6W0HycDiFYJr746WXLyrkMtaAgy+UoQKFEPZxMdtFdPaOPdWG
EI2cygAg8QHeBCcJrPhpNbbRYALLWboEDu2C9p5n4g8KzdvHn2641IhqUizXgaMfDZDr/2a/c+uq
JXYpQpWQrxDN8mkI1qMIXuvFkLwoJ1EIdEDiDbwVQrjGA4rkR8bTxlwVuBoUia1Q1t5y/pkAudRU
9ZzS9P69cMns82hn97A3+CxXEJOFD0Tlp3+/q/hZIcrY+LAWU6odhOnfMHbllAzizW1ehFZbfbhL
FvGlgIXwiNaiW1d+8mx4gJY71pr15u2l6UTqijGpkr7Lmg43uSXd1pKUvOz404MCzGPalparytfy
kYcyI6XEUmqpeToeCJF16G6NYfKtOsvxtO+yToxJ8Ie1W60EnRT91qtempwcJ0aCFGLVA1X58S05
quRs+g2kMml28HhQnuavDyvH5bvMvIYAps88ka3jPKU4av5yOKY7RQrlapgW0j1MyRVti+oYQFpu
sK0HbKKelbfCtQZ83/ncgC/CSAhcG8IdscbII1xJDh0P2VyN2okhY5NuYnIcQ5ect/rTZYEqXP7J
jP5wf/Si3S9xn+V7WPoH/dxMPGuypHBW4j2YCmwR78gPVBYR57hgt7px+S8oi2H0Nn3JvFDsTMka
VkIlGd3PX5UR6xBa236/xeqwzhP8li50kBN2MbaOJcJ3dMQ6MSobieHcsYAriyNiLGlGmJrIEWtZ
p3UL0wLrEmUMIS02adAtPwDrQ7nPfjM4yt2pQ1/aEePjks3lCg3+pYl94F58zAluW2xgnZUBnAoS
V2ZluX7HurwIRmp0y/GM1REgoERV0ZHwBoEIxD6RxeU1IHb2Xf893umPa5MNE/Xp6d3zbqiCEFoQ
o6Av98tnUpUbEj+XPqMElIVqYBQE7YeXVv5sy15fDQMqwfzOkyqrpxZmBem19NbLkaX22R8Cv0OU
9atqRpJDEeps11KXyRApvYNoHb6ql3+ov0QC15YEsInbO4C50bm0pHV8hWRt5Cc965tSpeiDpPjL
woBUHKRsqQAqTcxO92O+to06/mSkxwEABjsbQEwBMcGwLbslgmjI//wq+1Yp0RZ3dbkiuXrfrkLp
zY73LuoGv704g8sAQUG1JzaiHLqxQGW5GI78czWNO0sglInWxHKPTfxowYjEYxeU8lbGMkRdHNYl
daqw9LRfQMuwFYZDasbYZpgB0l4CqbijVgC03jO3cUPjnKU1U8FoIZLXC3p2Rg8iDISt6v/o8hfi
p7lIPQ09gb34Htb+mI5MGCbT+6Wq+KJdWy+/qWFDWFmRaV9BqxNVvPxTnUwQUaHdL8UjudGtRNO8
hJR/ASAg7PunL7ZfD1fUMwcMQUIMkWOTxiRxE/eXUObWWIV9EHYGYoFlvvUzmnnfZydfN9GHyHJg
q50Q7tjzPXmGaJtc8UacMoZzT8DkXndtycs0iPBlWY4zH/d5P/aAn3RF7dD55KPLOuevWeiKZU6H
YTh7Ka/o1q0tvxXr8LSM2bT1dlYYlxf8C91CIrxSeH1JqrPXdJUOrXnyrceRLbHvATwgWynZYBrV
tF1wWeWTv+U42mmtQyHPHKFROpwFbW5UGpCBfX6Xeo0zFUV/q3Gp1Gx4ax3HhuDg26BJVQbClWby
EDKEteBSrkvJHV2YUQVZLDqzkLx3Als97PCnF0oDcZhmHJPHPYUuyD1oc14W5G4+QyOX9KIGHzDe
L+OiV/zUoqIgkQmG3o3eLmRUpgdomG1+bxQsldTzkMFI5qJu8CA9buInHpxX8MxI5+vRnpHWl4zp
2ZpZKD/pI73ppeN/ReK/J3hMQghP4nVw0301bWTHCo5kfor1M+hE65im4d4ofh+01pgoHCmXOoZW
Y8CXBwJCkrGeCUFS2fLlCj9/MExJQuuhLwBzL9svLjIr8TbFAA2W968R7z0HMWlLZdfzXVTz9iB0
wXTiXAwR8FsFKyEC622I/ERUTUh20t/BH8QiE4zvQOUMnz4a6my3duICzHMLAHjYtyQmcowjw8vB
0/BhyC8F58YeguuvBqTk4WYrPc3N8GFoBlFvXJPxL6Pfh5nuHec90iEBhZXzVzeSwtdXcqb+HtE1
VYJfrpBcsyQANAirhIUJW+X/DxP+AEG3J//VtB6nZ7NreJKtLAoH41I0Y7npQjaTW8D/GYqF6MBE
9HopBJpPIy1+E3c53772XTRFxIVY3Z60D5Ib6p0gsrSzqCPjT1V7nKy/9K9xx+pcuMM0lRI6sT00
QlPP93kCwjEGyC2nVVmUowAbAt8odN30n933pPqbMXxKN5aJwfssEiD6cKXqEDCEYH/73VBbj4jy
jJfre574OSThjwlANa6oHDLEc1J/SFzoxY29tJr5kItYqveBEx0AIQwtaH5U7L7Oc/i2oCbcTd0Z
eujBDXVvQ4EBWN8nmXo/kYjJvQKScSKgDvJK/OIV9c5L78+u4hvsDXMHiol96SDSz35uh19xIF1E
Dr49v6X53hYENiDUev6tbMVEonDMghdZ2l1e5sEeAeXnEEgxMGO+SVSy4E3clTYU2BXhW6bxpREe
nBTuTyPghPMyXpg6j4CIeifL9pjL7qL10jNqzTNC6+a0JoK7hdx7glTWukF51Gm8Him8S4AgtfD8
0Ays6XpDX94F1DfBXDQ5A31KGI+q+oE99ctvIDq9eGw2SwH9gCUIPNfwOHm3ZrAaVHGN3KwwfdBb
2bqqcKRpG19KMuvGurn79/QApIu5tGHbpjWhi4Gtg1PmLWXdbybP++HvWPrBnQlmueuWh2uGKQdW
D428+ZhGhjzKRAUF6wsJSIGwn6mH6Il9byJsO/TziK4Xs7SsMqiMzKGcTqNXUPsJbO7knot//YX1
GZtf2m8CqKTey99Nj15Td/ir1fHfXKSTWXUu2GB/B508n5EtbyDaR5vVty9giledw4+oa7fnE4dp
xBr20WDpbc4AyuzoNh6HRWAT8hdSg5acQTAU+VcqFzwiqxZUUIog2ycqnkZVhikJhf8NhDlts2r+
zKF6p/Gl5nkbAym6xWcfw6T/8YMgBnk9trgLmCuHoy8+YNxvqXchsTSoD/UksZjr8iyJdTF7BkFr
ZVaOW+xehLm2CF+sy7ubPHC+XwgfEgB01X641JZYyW/AWbWEeCTYhX8OCmQcrVySq5kK1F7MxPCe
dWZyJBOpSgnmgOVAN93WX1li4bjZMOYesTZVCZu2wcr4GZSYiyhvFdWuttWC11d78TX4vdjBj65m
dAIHdWdtg5LaQVIiHIJt6R8uJFo02sU1mRJVoSVkwHQ+gbY/5PxKegtJ5yIV2YK2JtB8TbmTjifY
T0sM/GGmA55HufXeqmAOnvtE/j2WhQpSik68GBbdf7+3DJFM9zwfd3QOJed+pAdtGSh/JB5M19dH
oMH4UaqkG/gi6yqYuQOXPnMzfwjCK4zIiXqxSPgAlmb7Q4c/StDlaKAYH/YBnXgMvXt9v4VkN71s
YbTnwL1NQk0rgg4OfQc1fUr2K2eXrNk3SJ2tspD/Q+RY8bzjSzOICvSbWaASfwHqFmnV23DwKiX5
fJF71Gz3jnEhKcu1uTrNGWWl+uJWStzMn1k8v2gqLWwktgXs8BV8RhEGOhme28peTtXvWtANBWGm
g5iq64eYt7qVK6AcrQN8bFC9+qy3zI//LvGBToDOk4/u5luoX7WiRn2qBp680ofHoJiKRdn6AzvJ
9bld1OWacEQzbIV4paFibs59wKDnAyhNV82tqRn6X0CkYRRRdfyJ+DpRrUH2BnjaYKER4FagS971
EdzKg75ljbz1Eg3QOJUiKDPDlk7iQcs2KLj5kvL21OVpicVC+Cwpuk6rWnmk+90GvbBAbt0nMABB
34SuyJSG6OlrHbZJMVc0bmg5j8JKSfHQenGOFZ6Du3lncAwJ82OPUCMfFi3F5oaCVbA96jL+DP39
Y+oGwymwOVpU6aIs/OCYV0OLzx41+3kfSc9v9/u5kJLeI86iqfoLYs67DCkii99y7cRxFA2Tx/m7
b1S1k0WMaEm3U/JGLDxGFkv3tyQKOIKubkaI8E7nBoBYN8TWDYcu8HCO9VeXWmeYGJksn9h8iLBs
gY41A+GxTPu/NzFxmgbzmldWiA/ftuCkKVSOSC+m83Jak5aGcfeo3ptVz077LFbHsrafG4P8MErG
cUr1biBSJi57bUWYoTJdF2XGVuM9NQs9NJdkQpW9lHa2f+Z2k3jUHDSOC2qKVWZJG0WhMwXQbEZ5
2O1T79V3SiqAdXOVcqE31zzOqCWcHLli8060w7t4eeHNUHx5olw1hFihgKcsZ0pnssZ99oOYuBTn
pWswVqqAN81K1WrDMZ+foh+gv0/2YTaMClJpg25h/1K01NXVxY9A/Nu2Yk7Zl7dAG78q62zc88cH
nIa3qFGj0JDCO+cLJbnb4m0QbF+NVcWkIXuF6mAk9Bt4c58GHJe9RfgNutOYJC3uPvuILzIwZ/Rj
2vtagxk/HB6dXr4q2jXeH1wOnBX1xUbT/kBpdAfYZdls3wn6wH1NXrtH3OI6HnCR5ZVvwp4ls1Pe
EnNQn65yySK255qZtRDDKwxWgNnqpJc2X7/eFi9wRpIEprLEHm4kHWhH8aqIxlvBNsNKdrht0q9Q
YIKKVHXGc9d7NmY13LkX5/bvI7p7JS1Ftmh43szXsNAVJCXNgBZPdofJdy4XXBvlqfYVN6MhxpoN
gCxsza8OQ60pjtZ9PFq47clcwM4PILlQ2/PIbYe/oMLS8fldsmMK1WKqdYU462MrY2udgnkYWOX7
TKjDlPLEQjN7Smw//n7uIZdSmkCirxB/5n4S0KSqyGuolQEu2oer0sBK9JJ3onBpvUazY8awVBr5
kmhAlM6soyNltODrbQRSrVQKDzraXnqymYN5kRwsxwHYnRVXcmfdzreKMopl8wp7EISRh/29z3UX
W1QYx9aHAQhcflvmNmuQnqbG3sMwRIGkJt+xKS93EU/E4P1hj4gSesOYTJ/0yqCWBWIer9QMHhSj
VCPOJoPtI7Bt9vRrO2nthu/SXsDI7xyU2tJLG20EfqN6OHISNeZ/QpTkxz4XCQM/epR9u3nF69LC
+H4lWnOZGVLmRCcHTeO52iCSGSQ8lpkW7GaMaFYdygEeEdoZeGFdOft8rfsczXNK6vkN891N4LvP
S3ySalfRjoddCstyVLavitrtIP87OzcbB8wXDyse5gJLUkbbLIsta3f6CzosajM19WWmocUm+GPA
o4u4zH6cjE0ZYUU70pbr6NP1dLB9AnPMA5tJqGojEZuHPKXarbTi5iGjgnQI4CGrsh+6t2bAdchI
avzNc8G5x2dYHTRPMeW5N1ETdcQ8suqpo87Y+rSZ4+w6oasPyIy05KwTJtaySL5mAo+lccdzLP1I
EljaNBM/cr06rr6T9FAY7C4rmtPSXnN7+tMIk8b8umVOW1aaqf75hBI4d5wHk68Hgmyb/n580ltd
d/ENw5cDlN6q8CxhbOkGFrTpY4p67qpfTcvfvbyVUZr0Hah43lFY3UWde+RQWhs72EDGh1KvDrhj
d297iOinl7L+qeoV0fZwUW4qSE51xH1q0gXGhzLF4zm+fvUtiADQh4XzAiTqgKoqdfReLHNsSAE1
SRUrAjeyDAj7W0kYSVH1RdRCS1D71Zh2zo6yHpIJIW3NKLthQGnwwoMpXcMvfZ57lnYjcNZrv53o
sUf51VSNraBRG8LnGpQj1odRM6c7xaMLljQuvGBnpSAEPjfJvA0+9uMk8VmKRVSUvVLLzSKFQi2u
zoDykLTRswjyG5QT+m1irUE6j5uzlK4hJ8XVzCnkMLHN/ggGFpk4ofvKjEOmcxYEH1K8u6q5fxek
GazMnoIiIzV3BTJnVcTiB7WvgUKuVluPaXa+N/EusJlmzuywiKoNME7BJ7rvowSl4XUVP3HPGMQN
YuvzpSOIz2GyQJZ3EXkl2n/rcKBB7UnIYU4aB2vj/hyTL6IECWeRvIOTMYjlE4+yU8Ys5ZLBYkCN
j9hQ5oNLDNVYqfkdLM6QgIq+Ihm5NGxzJeig98wxlLl8u34pYZsTDkM9P9TlrMhTp6iGdcnyImAt
OI2IwZcEJupvVIlVFifAftRgqy5BNC3vf2GWN1TAQzwYLXDjl+aDHS1eEcvMHmpOOOKyDh89Qn7h
O1AIs9WwEaCeViufHalEdREN73jGPxfOhbb9R2w70KJZEqVepv40/pTJ/gHko3CpQ+SifUDuyrKG
rqko/bvSqnC5+Mqg8SDZzXXNOX3v9lNr5Z4XgoW94mWcCJlHootvIsvl0dlyxXm5A4JjW+x2aPLR
cHk4cnpjAg5xOK6F4GUWlbIVMIU3VXatbciiurKErQJ30Lqt6oJd7Ir7nxRdQNO5pvsl9LGOVGW8
C0/KdP2sxoVwShyOVYUi20GBqK+TzSprUDBR34ZJTPSIVRWWv2Mj9B5Dss/gRJMxzzMzVYpP3Opa
A7gj8l5okZSYCFqLGRBX8X+qBvkTZ/mi8n4DD3im44HQfjAeRKrfCrFz10EqtKzPjcUdtenldKkU
CIC1i70FbIK6XLzt+qo01sHk2ydAWIDGeT+mwiG5NtuuqiEGhzW8G6tSdcTg4mTcIeCpm3de5xAh
uc3/WxA5HcjFWrpcEhnwokpdSRU0UuRYfQLtDRWQjZ1pd67bX0lgd7iKcu6G1ml6YKCaZ01fPTH9
Qzk6j0BCDFhxFNsj4YeZzP7Ev8NH9UPe89rc5gRiEPxEt798PCUpynu5kx4EoKPodz5sjIuLdwsD
3O3mepBGbxyUXowYzDyXz8fDFGGiRBZx5yRhtQFSkB0BBLHk36nrwDAYYKa3FntqdqgoTJNtmLr8
goZKszhawr4XjabCM2RGyvZ0tAZz7Z/CW7uufUv8CuCuU+NHmL6QXkwYhz2MZ7c0bP5TqPWtY+13
GlOxI6H0sPR7gE0XvRsex0TVs0lSF2CkXvAtQNrQ/wTelERdbiSI5ZwLe3U5Ui1xs9ESq13d1ypa
ejdlkfN60BgTVYOXJsPxsZKYgJXCCojQK1WTRIJfe1486IQMva0wJhssmWMsdndcDRLLB+2bvpjj
ShpjarMDBeC1GF9aBM4GTLMs4wdGKKSy2BTdJgVIQjP7NaFb1MgW2NuTxrEDMJwpIu8KrtpgDyd5
3ZAAS1kTJnZORpEQXP1WvGxZX3iPk8KGVBaQ/+CgOLwO0vQ4wZ4FAjCtTwYWXCZjMElLZ6FRLKnk
mGB/r8FmEh05oJ//iZVVXlG8cXcO1eJ+tIaRfk05dfF9pdlbG4Dg/HXfM0c2HKW2qB5jrfbyv9sa
Q1WHZONaena6FHL9Ns7kJyUa+856y35qJUqH5SQX1tH4e4ZxArkZXKU5VCyKhSsgWcVPmOwCNb5r
C3nMGMTTePQn+qXmuVlyCtFeNZlpKfXgA/nS6bJ3wjVK9koKnrmfIlRrFty9F99ib1b+2Y7VzwWX
j63ZM2dot24sPCgqswkDTDW2bewpzp2TJL9jJw0Qzb7+6b25HEV5l1oyZfhkN0NikVZJWSEy6U5a
OWgyIPTgJnZnlbD0AEvoykbp4I2lBYybYmWD4Gs6Byl8Qxcy1ofCSK3Wqfbn9u4+wU3r+Z0vrW/i
HSQhfbli9LJUbVYdMrhpAatiMSU3d2t4gBfNiKD3mZt6Q+GB529Eb4tVoGd9l7+jxX4QoumAsZo7
ZUW/V6NlR1i2yytoe70/TsbpS0tPDg0hNDNLYqgVzkO3UDUA1QgNoVXQPiyARXTOqDOc6yp2L15U
7yY1fWQKoxmbsABgT9OVQeWU+PZt7jHn4VnX1HtkeTs+nejb8eo8XcfRyvABZTUDxfxWRl1ojLw7
0b7c0KkvDUv0DRCWmz1u2M7BCCNdS3rB4awdE/UvNuKP7lt6ubCefZFhHp5NJBqbJMeHvgcpFTOE
knioE8Lwnz2s3XjwFNK7UeUFTLA1TTDaldKPLFEot/uSuLiAaGUHm0U1L0/0lc9rMtQCxcFsRdcj
I1MRskJMwWUe0F73SwtNoV3DqqFM96Ktmz7ZmiXjgzX1n8EIWa6ftDltLZyPAZLZjK+TmBjdhNGR
I1Ksvif4Gn2paVVmLK8RnpfC8LDLD1T9ixL9DSosyjgo+fosqvwi4m6HvnSsPShKVX8rFzCXO7R+
fuBdsP5jrGkOqs8Svs7680FSKlRXFHtXDdB+SF1oqo1rJrLMR3flxkxuLZFCo3uzR7ycyb2tGe5X
dqRr3iU/gRVxiLGBfJpi9N8oNxctcy0BENKQ11l6dJl3lpaBucuq+DrieRooU07wZ2hLSSQ84J9Z
WggqN5LtMF0G0buGIohI0JeXdCugPzYpPWpGeGf6mUO53VgVaeSv4psIJUafixlSvOhkVDy56tkW
wIBXo1FQufJur/A0F5jHyDWtAK8hUY7QVuhmU9zVpfAGDlmdpnOsYnpxfknJYwf5IuStqadp1gzq
Tux5LK+fM5GpKSdTNYyB23Ghp5l3tlKotrRQ27fzaXtmrWfh6gnzMcTgFW3yqrS6+Ae631E+Q4Al
Tvo59FiJGNcZf/MzKh5cEGNPqkbX6s5eUNvhIOAicA4w7NuR2sqiutfsm21R4js2dv2d4c85mm6X
VUj8m3zJacwkaA3lGuIcuyhhnHXqYlk7yF05IxPWgh1Ygl1CMrfwDrjM046l6fWDyw8xHXgTRx/k
yCx0fp2QH9sSrhkx3OtT5l086uItpRb+NK18xec9TfVmavYOrYorAlyI6Z3ZA55v8hkM/Muusyuc
JRb8rjQsaIpkid2a5uk5aVSzGoJOxnaMmRkYJSt+wBFMeNHeHrvG5OuGPicP3axZxGyIVVKjqNOD
Xy4lrnWjKPaWYIy5pDqCpGxmoEAGhIKvJysyTAMcjB6X2a5oD1iklBZ+DHIc5RKq0pxm+PaDcjRj
4J+xd7XbJk9/xrTQSzYaSbX8iZEHxBgeZ/nsoey+eM6u/T7vyP4alQ54B92EAakTd+G0GRGq4DVW
iuvJI8pDheceRkbY0UfzdyUbgsHcZY7QSPfnO5soDoZRFLBNxQR5LMX+R8B1P+Z44kszsqng3Bu2
ndBmguoAcZHTqMJdocXfPTb0SGHuAVRulMFn+dgHoGgePhFq6EvMkB9X9lggcZ7AfRNUb4Hf9o0V
IZaWiAXztO4fGLhfAGfBTSB3qykUAdCVXQSntUbXV+Xf/vhgguvxDZEwpLE3MX9kRpSPAEBz+ff+
ZRm63eMC1k2vrgKSzPKq4lCV8BfSebdd5UCGQhiuhm3W6C5Jkh++xaJGUmWoqTRzgIoO1kxqtKbx
Kzpx4ZmxFXdo78qKdVP1/VdRasQHnyT8VBGmXTT6VmH6IvkacPlls3JiQXiYLlYMrNjtICZP4vjr
WEevcngZTeWBR1NNr7vdRc4eNYp5yOpEMujduIxZmUF56ds62Zo5ZAXE9oQS9vrjRz1Lo4zjryKm
Ku0zuCID4mbk/GAiIhlxfAE7uZbFEf4AObhO5RDAultEIkH8LYVZw46V8m82Gy1z8NciNRqNdDqA
cMlo6iWkpMX5xQMGdeXKLLoqWO61dxCFgUu1xKONt8h2JpC2on7PWBo7kKmqYyXFo9qDnSlkLtpU
0UqoGNJsQCuQhSsqp/cwqORYNhrWxIuXEeMcEzkk1ehjX4vCy6Ok4rd+dI77iLKGjc3YU+VpwP/U
TmFxO/bwkJmWbUfoEmx17sASOqbSZ1E3im5j2meSYHYlHOJFtwTxDot/+JlORGRcClOE+y90D1sI
H947wHT7nsYmAtHFZ/bzOtQxDBRpSNqM8P8a7LSkhzIiqzW0vOOmnvYcDdKnesvOKxvyf2KUw3AX
WIjWkss/zE8HaFIPLA6J0tTHc/J+XNCDu4y9DLZEsqvumAv35HAE03Vfwi5wdOPJHGIAeieBAQTD
YRTfb9Wrpym9D6NyJOnnZ2nr1r1LH1801nNK0Fmzg8+OqFNIKEAGer58pkafwDXcvHX8JfHfq2+b
qlGl1an5QnDTAFyYAl9skq7keUC9GxGhk4wqQZEAMbiRz6Lyt6UwXeQyozsoTMOJDuBruXe2xz+U
uG0GqeI+G5x3iBBf3af8+QEQTUJxtbEwg2hPwuTsHF8+4UNR5/vqH3cYQ94OgQH+7SWW/rjPHSsD
k09gyT2OBn0cbWdYJgjQC22xvCXjqTvulmBH/wWG49jpnGgEvFZ4G1hwIXC2SLFHvKYrar7jnuI9
yl1Z53aVZ5xfaHY4EE6FSS6ePufMNgIHwSLoSMQOBGW/dp3wTkJqwN0o1d4YqYXbAH0Hzbmu5jx9
6BTw2dYbzwfuDDH0AE16dsDKE/o533X8WtCIep2kTyOMfj1qWA9LNndDtC17nUvGM8g4z2xrtUfr
amCxOB2Kgnjt7MKNvrkJmoWZljv9VyjdqZpZFiioziydfNbnpvO1g59l/7b7YkL2SChnSxbQMRzp
mq07XTErPW5gqW5KFgrt1+oZ/anQwpW6CFqchesCtfz59+TydS5rFnR+USaovBugmPZev8ioAate
dFAak5quSHGg4Zufv7PzxcNouRuwHq0NJIEzQV4IAHLH1H/sjSSLub6kubHf8BizbjcXEKIMuxbY
bI5HBDl0r9fL4O/wo2MzUR2AEkfpyR43OngPwliEhYo74k+lPJwzZFVsZJ0Z0vkh2nk9ZTob015Q
e2ktEhx/gw1IC9V2J6e0BhFZyIGpJu1L/pZS7JuwHpUcn5XTly6blc+5uu12C6rhb4kAd5ZbdtYR
bsk9WPmLsMyz2GFKqmrh67bOyQx2br51D8bn8WKVCOPJ/aO4f0+VJZHQrH7TjLi7S1BgmtWTlXnh
zMKCzBBR67ADyXKj5KiLKZPzJmgsdHlA6gIPzo/jD079/c04acyBT0sb6j8ulkI4JbU9UEoeT51M
+/K8AUFwgxjcioCJyvsslJl1ks+q3v6zGLr8++tElZ9wB05M3AvR+hp+diyZZ8L+qQuUE6sO/Zot
paZZRc0IvDZhUSQRVeOvKv23Z/7vRUzCXfS/Tsrzf+bOp3DSn19pRClz7SZliodfLJtWVqkBhPnt
UXeztEPc4jgh1WMcLfVcpv+tj6Y7HbZPNBWJg//Yx9e0r9yJeF3TQveRLI3Ym7QMHi/irNV9tHF1
ZY5ogN3bdmZJ3JhLulV6KupWdwtygKInQI7HjmSVmyrpInz4V4jWwSoTFKc+b41dvAZ7cjmI1JdP
NYyc3FxWDNBVw+IdIq2BURt4gcjQloXzg75g2mWhEqg1WNmHPSdKgeyOgKuMMaeRBW+iAp67reCS
o9bH9QIfffg283WdR5X8UUIztyy5GJ/rHFTfDpi5QFL6JiutGc4imncndkjZVGMWrv8U3wMnGDT/
wm3WmILnbI9GAyWqPd9Fzg1iueqRGtEQqjbfkJja+QznPU9Tg8ZYS7LsNFeWRzEZ9lvHk9FdWO0G
1u7S7SAALQ49mU0dZySX65VqrAwLxPMuQvP9R4XS5rhVhtC94KpYPRgxOoViafISzpFTOLLOlJ6U
gi5RhEeE+PotsZTSlF4ISnvWVgegDEDahWZ4a9Fsj5h+brSjBnyo9J7kkZceuTugBL3n90QyYmI9
h+VT3U7fIWpgaNccBB12nulcOr8gqbH0R7N6RYKmffP08VUoj8J0leCElb7u5QNJzxvF1F1HcigS
j9V4NrBm+6fyXIqSCRMKoTB7axaxzyD40tScjIMf4gCvSzsoiWxkYpfInp28epdyCTO3er7wEJp4
nD4b+VtRoFHB+dUg3SHKm3NGsY2NWyOLQtl6hemyZPvHICryO5GY2OCjOAAk7ViBcG0SW/K/2vLp
eFwAs3shExJtOVbxjW8qwgR2EIhU/Ro0WBmtW73ivQwXDJwXEUHEQA4OYDMOsU4yTxFqPXIb4BBr
ijZeGg+MzSF4LoD0YdWA49BguIecraI2jp6kkhopZ0EG6HQOmo5z3b7lO/x8UAbJquJesjxr4rua
NKAluOXjRXlYzT4BSWBJd5a/w+sPb1c8s7R7SmOf+JaqdLpxOjdHLXTFP6U0fZ+xcztu8bZJMOsD
TdgfwM8eFUpPSyaBI0tw+/k7PDmKa53O55NFZC7zpsucZ7dbdoYu4o1DSDNbQU/fbeTM0l3Lt6tW
gR2Ix13dfIhmwpWDzgjuM6vOYmu7XKyOKHKoJ+l6Mc/4aYQrDEUwzkbG7XY3W/kwWXxBwD3deRXQ
3wJ2FkCGoFbcRM0NO0e89XxSl/Dx2KIub6xF8cF8obfw2y7NsO7NFs5Fr2Gz13dwd6mFnCPIDPMd
EeGgoggGulbuN8cbg4L50fnAExYFHFG0oRAvuE+PBbxDztZVXLgFx+R5p3vdAkEKXw3OgXlVnYSG
YIwB3oNXLN3F6tuxH1V+fpa4XMOoOYfDapsFCMIvycEUrim/QeH255auyIaAbBImLJhGTqHC2icK
5OhiX+PGVPq7UMwlQl+eSeYIl/F1/AGWpccpG5QOG0kA5gQvdZXQ61lb26sQpIpL0ZjN+zmvXW7X
17ogjfTNcWmsKYXWPO6RX+RMQbmjhEVjLwBo8q+yJlm4VP4T8IhYywKyQJMmZUxYlq7kzIziH2hK
rWs6w0aYt0SHO7+qdX7OnPAh76DhmdwHP89Iw01a87mj7Lj2KjYHUJdl9gZx7sUg8TDh6AzHaC2x
Ukrwq8WHdwpSEqAJAPgHZEjZnYu6dB3xkXQUUGswoqCv7RFpi1ktFDg1vl0tGNb+h+KWLOJ1Nyb2
KvtK68mmG44C7/P/xhglJLprpLhh7ynorKpkHt3YY6wzrmRvhMv9I11V9cdrR0f+OaLNOUBhOrJw
QYeMBADQ1yjuoVqR3eK9GGSJijgofoj9h8bT0Bj9ZS7VSbeI1f/SKTd5thxGPcyIuXtvryosNxkf
yOI0GKDNA7RYYEJpAy/QSk0+aiB3F9KcOiPb5Qwu+/x3LzjJUMa3pO2/rTNFB5HuBQpFfVxT3XpP
MCFxHGZeaaCJQw4aIDICxt3TozyJaKqAf3tKCOOgboZ0z0AFWv/dAuuGi/hHR4JZefapfdz6DCCm
nnceFRc3NVbnhGpcwPjD4LRcfgg87ed47kkQ7q0P5sJ92MEEBkos3IWGCQpP8rxoV6yNQPrYaO79
QcgadV2CO2DIvXY0XlA+aDl+3TJ8rBMuUYjPrjViddqRHkWyuVwBcuHz7WlQ+r4rdcvw6kZWufQu
DZoUeB0Vx9asQcp21QnM6HOuuWhYpsnzVqFZq65aXcsCGU4mIpoJIKFKFRraLahXaXplpNoJjMq9
qW1RbjYQNL0dfnzeyyLPY5RHkB+P/EFyqGk47lLet/fWTW+NpPwcj4HnQVZ1wyn2+0JrZChfJxyu
CPgG7MsOXGzpwsD5xOE0Y5L5eHdXb4YCh3jFfy5l23ee4tyvwqMd5LwR6ADg/J6ukcZUMKjAhFXe
Ceb64YGNJ4AIXEhxe0EsPBrxR/9hd1aQkUUOUuZOR9RX9jTetH6BPxvXOqqH+EK3gw7L7BzDqHKo
uLmHEpZ7h8vddn+bjrA2IqEVc2sX5MTcZkXRSmCtGrCttYek3fn8lCqg0ucyV3ix6aIpjwJppzBS
xDQ7eDMook3Cr0FC+sY3thdvbHJN4MpfT9fQ4DqbOW5WRjtbl3CWcVMOwch/Dt0uSWxBIn2RFyQn
Rcy4/yxoK0GwLEzVpL/buoozS6sXQzslji2Ppvj/XY/Vwo4ag0HfPznQ29/f1qVedl96syO3lcx4
IN+NwQBR08hj3wm2f2KJNEaTEFQEJRATd+RWnkLK4zLmeF/caUSRh/uGFFQYLk3A5ct6fpkWwqKg
QEqUvwdb9IGwCwdV7KgObwOW+5uiMzxF2MZr7n3j55y/agNoADtIM8Qmfc3egZ2razK8Np3nLmNw
KzSJYH6Wu8LaQJzyS/CBXgM3Q6fWjlnPpTptKIL2XbPrxCAyEKD+JcTcIT43zIXFRq66fa3xumbK
mY8CN3WjR7EvEQZGz+mPrY6B9uoXNiXy5aJ2iSVn1LtBgSdQdD25huSsh8u3Mwy0umSEjW3wlOZW
ndkw1x6l5rI2aoFWfpuUsk1K9XNBak+LXXNa8t5d2VOCDX+0hwexhBgxcG/va2rofpAkry2jZ4qD
k2TISe1Ih6YtVWBENfnajrCoqPn8bIlme7i3jNyVWCDRnEziSmx4tyu8OnGH2N8jkPplWQ6SKQ2n
+nhFgIVjHHJuTPE9ZmHomEavSLiwOa60r8L15RbcWKD8QTZXTriGMzAm+EupcUzlfTit0ZoqrkfF
ID9fwo3Fy5Gao2UfbaABnOohFys+V6F4xfX+pW67fsYnLCPVCeD9IRDOVIs9CrLJe0S/2gWCvITP
7PHHEjOb5wE0ql0bJ/U/VqKY0drBm399zMCVLD8528us4uleQJUxgAu6Olajm6HkxG6w43oONYNP
25+75eFdknuflPLEoiZwpW1S49Ntd0mXFP2gQAx+RVN0E3V0BMRjUrbauA2m5eLxGNNSmU+gIKCa
GSNisRRsC3LIaEuGi5WrjdYB6Kk3bfanCBJORAFKFO8MD/6lpkr5iHwWBEizxMwpZMYIevkC+mMZ
Qz+MhYAbyz5ZklUgPHqkwAb+XJZgYA2P5417BS5jvuSXoX8S7Vo8rpaj+/56VPOgKvE2CX8cgXdm
4dffNTJqVFmjwvrvAzquDSyTuS1MzBaTcZnR34dzjh2Fg6nebw53Y7cwjrcnfpRLDPF0juplddzN
rGEZLRE23FDx0FNsmuPWoFvv6RCCgGdxKsyp3Q0KEJxCauZqpf+GXjueEPKKCxGSweb2tUgqBkVF
fNbfxLFGNy+ZMdA4tseOiRQnovS3u5CcUDDKAIs4JVvjC+5+L9W8UzzWfyXHgyRwLy7HbLVm76PS
FfwOailrnW0spsRcEeTsrrxwK35vqM8B9BIDt093CB09w662XXIk1WEIvnemrZKaw7/2/DIRxMlN
PYGS2Chkbh+njNB92dT45Dn57xIdEfJODkfBhp4jFc6AYN8ilsO5y/o1PEqnwOay+21BLimhYTgi
MMbLcKYZnBBzGePFERrS6inApOjsrsgHjpSV8LZrrJ6StcnTiuqBQMsMhdQzj31KjdFj4N8ZreKS
YtFYBNnT/yLu7yMZITgRWUF8ciO3ML0TDjSoVeq2O2h11I/C3TWDVmtEFyRKtK5CXFvDnbgv7zOS
HEP6wJZl6B3E+IpeGvZsYJtUYJd9bPIowqAzl54CYsQ/nQDgUcyE5fV9H+AIcBS0hav+dU9KVwxn
yMCTEtniJjLuKbR435qcb0AhBMFipJKHmO6u9+5LHGgvZYG168Pejcmu+N0NS+IHlziG1q+uEOYq
5RekcWsyXXzXSq8i73jCaILKC7aP6J+ArJzjBF9qXT8oVgeHlgjhKFRB8kETZnbrJ0oQJpxivcKc
vV2/n9jDxKMvEWRYDDG/JhBxTaA7ZO3xBd5Tb0BIO8/s/CQ7jTkM2OD0FZ5GzYpnV7liEU9ASG+2
T8Zb3aoWSH/cfzAdtap4sKpk+V75sdALA/1ZCgWEvdoEX4sSYrMkOldnXo/PU0dXp8eaJ+Qqghfr
zNuefCqu+CDtgzNZUyWlIRmoa+GIMFJFcOA+cNldXzR8cTCxi+5MdzbVMXMnxuXJWG4Q5Zqivokj
D/Ug9H2oxzneyJtZvlki0lN6JksSKUBFohH3roN/1uUU+3/SggNDzzd61fmKRIwuXj6VB9zNhrIt
VgYMwFC8BbQQvOBvR56wnBoV6U1A7VIDljJIddSTKjAvt8l+Jx8CHmU4F/Ai4vXCamPhDJaU07n5
CfcoIjbEkojZ69FD5pXp1nFcQm3BBZUNRU+nXmGkS4o/aiPDUnVFfUozBb8MgYMBfVvQH3vdvFRO
KluYnl7io/1sgieEfZtQSd0oH5HdWHvRafQWrvSuFnnBGYcBD/C73rs3ec4afS157PEAtrQ6qVkK
SwnlXOmctsUt7Ffr42LlEZAQ1PUx0NxdteOItMNvsKBIkkcoP5LaJcyPALex5x0lESqCwN3t98BM
/h3OVU1iG+kLZAZWmrkqXQ9MROtXscSWjd5K7lEavSehyWUHntb2n6yhZ0Vu0YuL698+wQgxorEF
yp/MrLC5r7R3qPGI9rqK8QKslw4vsvSdT6+3rnC/dS3W/q/e9TCsTP52KTMZxgCfCoFzx0oqX1/q
57ngMR9Eqd1M5PD4bs3e28/MYaw1HVX1Hke40DWYZ7vM1ak823wXydKhlEcfRg9+6oEpFFMsOJI2
dAGqnrhrWyvUGxNy3qCieYNKNbV9NshqkCCbbWubGtMhvnjG9DgQFIf3Sbh/lZ6XE2xYPL8K14/8
pCnGWkQR/+zn14BFTVxZPlSyYb+nfXm+wojFJFCzTfWbizZD+a1pJftXeCFSX+i7gp49EY6ctf8y
0MyOmkC+NT4lvnouDLGYxnEIpWIJckfnZ+LVZonPvfLRoOfpK3kCH2v9oR5vP7m/VPPhMlHM2R3N
zorty6gugbm8tkKBspokx4MmxU4ri9lmMak88GcbS13US1NEoL2XL7fMMoTlZJd7vN8lL9oz/JNh
MrGuFbQ73jywDMxaSqCJIl8F6MnBVRuow6xZZehv2Svzy7kiytBEWCbaf6btoaZ6Tn4L3pRHry/x
FI+JdvWddw3OFU4OdRuTjqZj9SBU2vPwWDG7YIOoOoWZGzmuJNFq8jvY5MlqM9457DB7Kyy4785Q
OnEb2a1fiOAbOUVUZRsuOH/ZUx4Hlpg0seJ2Qrrgj59lZbCBrv29pSnT3jHh+HGQq7ORJMPf+/JJ
sK7xHel+kXIS1FRtjOFH+/fYOO8nz6VESPc9y2rWRDe5kOsy5sXMRl6rgeTKmL7zMOQZrMnR1XRp
MgyZPSx+HtJ4ydNZyU17CapIFiLfOl1Fn0FZ8gE2W/8VxqPcAamlTadZzQm2rh0amS+aSj1fo46W
iSPNoLbgGiiLPHNO2c3eMSWNEmXIVNWZ7AfIZuS5FO+ZK2nMqcwxnXTLuKFf1r2T7xQ5u5AYNPBE
xNMCW7G3UcNNEPrn+RhtaJMUC7xatIyrqGEH/gMtWlnoS3Ev6FnmvATbWatLqK2vG/k7IGExQVtQ
3W0RZpEPi9iqlSM2GPqBK0bRV1KT26EuIId0LUTqiqamrjfMF5hiJk7cmS0gHc10wFjjPyEBaURR
ipZg6s3UdSeH2tjU6lK1Rajc+0TdhqcNJbMKc5f5YUkIcF0ubJprpKn0+n5NRBGDx0O/QUJgbl2P
8YLTiROaWLpFt2Nncw4+s0fazSdWPvH7YqNkwncPRSf3sAWfgql4MfSIe69lfvxzo1jrO/ReEzgj
JmOAFEhDv9+XW1kYvNX/bUc/4y6EkkX6z/EdMVCo9u7XKoLjqtakO2lFEsw/DPjdH8qkh5ffpzbz
StofVjW00wu7i4YE7WbeUCMfecKVjQdPQhhwuWWqbwJIpaGxANlW61wVpFUI3hIxxHmN2Rq0trIx
iysvH/sZOIeLmtE0f1PPD8ZgEqV0Ji1MEcqv6oojOzIk9CmMmCsJa0BMcBouciKZQqJasl5jG2/G
vCMq8aGJ/IT4i0JuJMVa+tBfBAvCzMy7y1waGw+MAhr5ykMk0deA+Oz2cT1YniJ9qUWrIzd3/51R
sk4+PXrnEAYx8LlvB5Lh5Ny+6blIYukVhNMT81Ko1iIjxJHKKRysXhNNsWadjaQtUxXzgTOB+ruT
c7on3d+KAv4sRHCg3oJHPoH6x/5gQ0qyZoL2QD7Na2CfrmVKexbh3cKrk6+x8aVDTdTzAy8RMb7u
eDDI9xsQ7qeqVP8ISbMu86EF//gLWpfT+CK+lCwGwTgXynXL04oMhksAfRrT0zU7F8GLqCsqYcj8
SSy7T5IV/sHCxqVmkPTd1gDR0EY6Tqsaz3WjiEg0ATGjrFed8HIAupBD+YBo20x++TK+xCWOEUAc
WnkGIx2J1HvAHoBO+7gH95lgliWzr+X0J0pWTQQyhQwCCCDA9zyxPPyvTGqLC0YoWunWYMt3s6rc
N8LsX/FSBIk+KtIufNRl1eZC++dnaNpxIuu5OLDUEsPXJyGrE0KIMIR/JyU0fh7i8uY0/5RrajmD
M1AVWvQXXF9MKbv1j3dqnrbf5GrzbFY0jgE2f8zG4LvgyX6FJGz04yKfpL8PfIpze/NLsV4hQYfZ
ABIYUgXAouit7bj/cOMIBLmGaglRCHZJUMfyYw0+uDNCC9/4fqXr3Y8EJdFNziJcN01civJSSgAn
sS31gMc2ElRL0okFK4m3QG/E0iONDcoIWwPlxm5JwlRLnrNs6eNTImJkMAxaWktvXXttTtNufRj1
UgAIbOT31Tu+vR9UUnWCvdCZ6SFgzqK6UCL7p7BYK9Nz5tHB268Teb6w2qRfmV+d+7YtwiWotteK
SzgMQY9jpR4B/HC5XRRALUX56FnXt+NP4qBw57cU27AwtveaC4DwOma5kyBGPh8GB2MEYNaxDjZy
f/hkAjtZqyDMl3rHE0LL0UTDuQg5Vj4U6CvoRsdZ7/4wEUKbfP4LhgxJS/84RIc+4xZ5C9LMmlRu
qimn5egdh7zgqY6UxaE0BdSn7HgKeBnxJKO+rLDokBhm+4tiv0RYfRiZ5W/oXrRMKol0W6I9Q7OU
xZg+64aCbwBOF8Rr7o4FUhrEuW2Nb1EHwCEKN6gBkXKcbwlcsvbrSp8d2p9XvCfpetNiEC/M4eTE
a7fdyaYmQ7BkHcRKICFMjAGUOY8behFnb3Fp0RWzS/eaoN6FVvZNmA225JeS0RjF6UVR4pqRklKo
4jKWPlyZfS810tiaGaVttL1GK7gblWtJJc2co++kxV8c0gtrqhNSHpQsxAN29jPtoxywOwpSJygp
8YEhKskTwZi/aExY2p9UC6/V8UCkGGnFPYkTb5HCrUGLWOjDqvKWB46lV/V2MaivLuGr7kKebjaD
grYq5Wm2TXb4qeLS6tz5USHg2ghdTVxJOAhzOq+9B98Sr8DW1CKaN1LbIvOA/WCMLGtzTOTjz12T
1vMMfmKbecpycUYaMSGUZ5Zo9TLpcXZl8pR1ddbnpCxlpmyQ243/HidA8uHskyqO48sB0ckLgbWF
4dWuzGE/eVdwTqmqn0mQA6k7Ez4eEIE90kaT/x4u+RLuiih2Q3wIhdbzToP0aGN7xp/5wR/aPYWb
UvokhCc4Sg8nfVqS9ImY6Zj/jkIeEM5NPYERm+jdob5InV7n9viB8pNUmlJvqcNT61Ag0BKsx0j+
SNXxJTtRLFvUpdznJYs6r4hBSGvaQX1kng3fI45mHnwQBRRMcj7smrsFOn6fLX3SC9iSUcI1DcGB
4h9VIi/5nF8oyVwQEuPH5yg/5Xc2yKK5WkP/gstatHcqBU4QuX8OuU5XAk2ywUdHW0mAEs/YrOV8
09cfk4zmVM7fCBsodlGgaW/q61p8YAoNfaFmyb2+6XVA3zqFgLMrc0uP+ehZZJUMIm+vaHqr27ZX
HyLGLrZz2pgimzTu2szJmxw7SsJZoMY2DO6QIZVFBUUQETnSxWl5o4j14MqFPRxh+U4Bj6mGbOdy
6zztebm6ofsi1fCGQCDFSDDz6sT1CYM72AYiZGjXtiRzfkEyyxXv+2tD6oW2ZVOvr4FEmWbDq6lG
/lb55CLZtbaSowGFXS3bDpH72IKGEEWvjFe6sr4K2k2yDqqfYaz3b6HjGZJWGOacfx4xdl8xE4IP
Nxd2sEsn19UCG1qj+xT1c+dEoOlgnsp8v9mW7Xoo4r6bSvEL2/6Ejv7EGs9p6267S1J2uu0VDXGh
8ZIW7U5cKeDFk3kIUwNVs7HZgf+8lzF2TUPejLnILGisRawTnW5Xwzm/rCENGwb3naMd4+XFwfS2
uvDbaPPePpYlDyCHWKd8NGSw5YeXzMpctQOtjIT15imV4RAZ4ErIVkf2DbqF6bfXKOMH5U4azEdD
sdv4vw+cNB4TEsONh27BH8/8vZt98uMxWk+d8sbdvNuJ+HIxTdkGllQzEdTRT840L/k5pW4W2U18
NBWRsrtz3+0E4cX7LjrqCGjaMcS7AyQorWjuLkfJkVqnUkRDvgifocMvPf6BMXuBtYdbkN+KzIlC
OgTncevmias15HZsv5RDPP7MyvuWPAlflFxO1OebTM7u/fqLdbkfJjT8seilmklmPGjv3TThNvqf
kj6oWQE8AQveNhLk0AyfqyULwd4ZQS8K2wxvYcerPJ8C0Bk8wMm9in9laUO5DQjpT2pqg0dytGb2
g56Qt320fPFhYuqkoQI4OEsSLRZveabnQ96EqSLUCjcNLmgpdGUvt1O+x73jv7GjgAnmEGEFDbH3
GrIEji2aRgVVFekGEf8Lz/sgH6iXHRq2w6ELOQ14AyevkmsDhyQp7DJB+3Rb0ztx4QhokO57cWWk
0VAgrK2WlZQveHwgXbuXOpZBSVHqYn4tb4I4H/3GzzVgH6LsZEZes5kpWtHyo8C2WWQQDsJOcNPG
KJGhgEgUEqQ8Ms7i8ScrnrhNSOtLo18DAcGEl2g+bP9UtlnPrEPTsJupFxgoCX+WbEWEPDVDMH51
nJxUtpUR6PFmcV9EKxEVRN31oDEv46WEWMI48vNdf+L1vtpielQkesE4zG1kPKeXbCMCAUoCfT0Z
F7tVQq6lgQTCXyk3SrgaAz6pzxzPEDeeex81QgexAbFKrW9DpKey12z+nPwUATGQy5A/Jg05jq4H
sxjF+XJufwOu6fvumoKApaqw4kNQ2ynPiWtIu+uAm+CXlpQ2G+m8CuI3ynEhtF7KadqsScntqkL2
btWsANWrE/csRalcxfQkG2eV8it0TysFPsa2FY5VKQE+0H1YZ6CYdiT3geqT67/7jQJT4y3DN92G
dHgwT2w37+gItLEEWCIDwiE/JyCH+w9YHRluOsdqdgSH0YB/wMhRr/MDv8B+C5roSHnhIlJK5LTT
pALmsSG39ni6WudNWwPZwDagoG3puJtI2FTJ83FzeF72HzWgpn6S7qxntOzi9IEfssLs/dovnS0w
Nx3qSbSzbHFyEnOGC+7tGLpDt+acqiLyEivchoqYMAbZpgEDG4YvUlcZBv7qckWVbZha4WQOvdSu
0yI1CEUUoYrzs/vPpKxsM9xNsn2FEAtzrBW1uF6/1OqtQpr76Z4BbTfyTAdZ1xYpLs1ySawc2dhr
es7IB8qPqjjh/KLDRtMWWHGNhnsS5Tn7I94XNBbx9QWLKjlfBOSnKpPeYJ0QYUOLGhuQyP2M8xyJ
eaIBxU5IYNhpwTro5qzuQFAGld/gSHEwj04B+pixxNfAbuXOo9Li5/NU5UI36WaNbM/ha0fk3XgC
65Tl09+OTaWdcW/cLUvgIPQsQCke3K3oEL9JN4L8gD7ySK7y/HtPaXRbFn5sGLSSKdXcgM+IWma0
RxWS7PqpbZClj9cw982W0mlN2XynIRAUw4ZUSFvjTmkYD7e//3mDFZgjqc2T2363yVo1G0cd5hzA
BofxpwY41bLSLGWe1EJBpDgAdvpOW0tTW5BKJRrJuReoX2I6ZT+E6bEKdeKvwJX67D5pB/fWj+0a
zNhU8cUOLrQUuPneAj9VGNkpZCq95ycMfYSOvtyX+JC0wB/K08gDFSeYNwSgmrMGcG0pKuKcIGix
e5vM6UGvvsMNCPNmhcahbARGcgrkTxuozNlbevtKFiROYrVV15SJAhF7UCIcKxEY2q7irdX85YaR
daivOO2c2BVacy76qKkwEDXCcaym4qpg+tfmiVs0MU+5x7728gYPEDlW7IFD/t6CS4w5OnAuuGM7
zLk/kqQ+j1v/hIHUaDJZdzJdsE2669Ah0V2aY6+HktPX5DEGtJT6KlU0PX+neqiPJuzOnDvKEVIj
nAS1IRqDHFrZigJ3gQnLOOgdyMmvstnIlegqI9CcyELGRTYOGO53t/VJIzMYc+Y8iwGnR86zOGyd
QXLvlxI5TiJpI5NwTvHPvKtYFL55g20USPz7+oeT60P+goxQZoJgtxpD0t/1SOMeRErcU0NmUgc9
/jH+p7gnSe1E6nv7l/cd3DKxYel8BVheXvLXH7qMbJJ33C72WssnGfjjibwyzZEcbulNgCBRLdCD
G6KAYmz/SnuIONoo01HSSImkZwRf/V7yXDgJH2FR/awQxuiYZk9xruFodCk1z1QHCgC+Owo4ND2A
nF8UVfnGZVEgK3bUooAfvFYEMfuBZwCHljvwz03Kr6vUUlPa/OWEfry4WFPa+TBl9tblPIFolZiT
f0fBXQ6G43Smtacn1F2oWVUugjJJBwH0nzYybjtG9BR0yq349t7PxQSVgoQPnDILeUvgsgmJSc2Y
Mv6H6Q1jXlPMQN9H1Zi9kTChSvI5sUle2UhT/70ISWLLpRTIQJJONEreIak4FWOIQqTa1WoVASaE
92ih1t/0AXsYPF7zauHk396ZRD4V0UOD8vYFUsmnR6koQEm9EqWjlUdGfxnLHWXIZkVN8I7iIKmR
X0aw0Ng24q2QPsTUfjM1Vb1jgWJw6I4mB8/r7+9LufRdbgaC1u3kt7/Cx79gw0t928zqfDLFHnpJ
RHMk+XpmUMFFwOOU2dQsyWYwzwNJsQZGyrHpgsmCcv7dJ9NTR/Onb8QNU0G/JR0aUk3OP4t60gI4
Y8c/lHobOXJzgJNLtVnUxQop6+YFMuuVWHsoratVGreBSlRLfjOnTwwbvkxw/O4FANRzErY6lb/L
AvNEbLXC91KakkdSO03uU+UVSp6iFNjueOa3K8pgmYY5/GBa2ewiqiKg2XcLQnBaYwZjY51qt9Le
8DNMj9MeoT9lL94ZAHugWEykWoMOjg8lQBO3MuDy8CwkzrgJ3c3NNG5te1c8+atK+0aUrW0EWevF
FwgF3t28UrlzUaXDX+ZKK5ljKcwU8QKXDMqQksJwm9aU9E9E2hDAjXkho7pvXgpGcLJowhX/8X/N
/vtsI9q7kR26efYjE14LOeS9D/ljPwc2/onVzG0mSIAgUdkSE2Ait/4NCd7miwsGRETi40LBKFij
gswqUhK7l+GBfqG/MNC7UU3j2vN6cAZGylrp2teB0+0OOA5GSZo/mi8yQ3Shh1cSCQ7gdrrzOqtO
RuHrX3X7HKKIz+CQn7heowUZwkp64vWzGuLJgNm0x+WniLgGfpWih207XihcNY+I82RrYI3Mwisi
z2y0AdgnG5tOqdJL60B/cus0E5ZlhtahRqyJ5QKC9TB0DVhE28AfcpfGimhOsumA7WPB4Tn7EIWk
mVPwLS9Xg9qpeMIGLFCQo2/buVmMFrrPvb48gkcOVT+tAdGfvY72z/LFc+nBuhueA61j/aypAlZ/
29zzKoAUz8RTafx2N1kSsI75hDKHK4PUydXzqYZGVHY1G2Ts9R9VpPv4WQd8Hx4lgOJxuHtSDsxQ
MngJsh+jH7H5mdwuSG2Uz32wTbeSdfyDDDMNkvrpt89xsBBwON0EsyWYArXx+lyKHX5cVHfjaTHT
UN/nABh5qc5bntXNjny5q13AlDGV65Z3Ncopd0LwXEMK5mwJ9gzm+sfpa7zfipHdoiPLHKVE5Xgr
uIWtCfYKyfDf0W2dE+j+Zpo7RSN22SqJBZoommyNtYUo3VeVRWKK62BCsDGQQsCQe2XXvrFwVmxs
42UIgIFCKmhYNJJjBKICNjFSaQhKB6zfuBvB9T4SPvMMUfbcP/TIO9itXCszhueyTnnj9Hvm68ec
SPTIVYN/bCx5dmPsg6qWuInuGEFpI0xsyEdMCFMQm54ExS7raRhl8Q1o8tmG3m1xmD0XqDjjkupB
wF+XsQjdZmP5ZszitKCPBsLcFnRfP6re+sVoAgY8Apahm0UEcuUBA+G0IPzGZNj062c4KPV9cfKf
qjQeNgy9DaKFtg2gu9Bkr+Zdz6ZbeZWknzmy4k0oBhPUdQSeQaX2QrbSMxegVcV75QkZJe7VJQlo
47bIDhgLHNgxEx+XFQaO4r2hksPZBF5MCWuLU66HMRRr+K1kNGAHXPBzWr5YnpjXAsllEMDnhhDy
PbNI2N4jude1/JXxfLVnEVbgnrwfVq/gOcazzNZltKh84XTy/zcwj0P7qSvxJO1Hl0YsqFobYLzO
YhmOqd+SbgOhoGwgBghK0Lzlm7EHdqEvtuq0Y833s9IiB21MXlriQlzItDPOo91Yvu4FFHTPbx3Z
izCQSoJbLdKwJekUGy6bI2jw1LQJqMhefzJ34wbwZFfUXbWYSqfxEvkBZnBmWyEA9fquqXim48JQ
M+b/DDlW4vPDhOjjYZPWRm77ttCGWNZd2Bhh9+Ky4Vmn7UuLONFE2pt5RbhFFcel2vdfLZHMvWbl
E8tTE9IZIyxXUuwzDtIIn0kOnfyFOGU5BJEoV++FofGRv3gjoTKswzseE7cvZjgbHGNKu8rvT4wQ
wpXTckqYg3zD5YQpLhRKFtfHWWzqSchpcsFlaT4qyWly25xIxuo9HQUdpdK1i9dqiQSP/OA5BE74
u8u1XChzxy3sb8ZXAUExeT8SO8k9aT1B4MaWSdsnM6j4Dzat8/OrjyAyylVek/4xQ/WPkVBFC2Pj
9NwNBX9WweybSyt311TxtQvlBOQpHteW1YTDSdySe1r7k9XKTsawodGScyOmIqidhRfisD5jFVu9
3Sw5dbRjWI+YHSYdSZgioqVNROMTuf9rfdsku9vPG+pLAAcHso7fPKgZh6482jL6RF71I9Hfgk80
JhvWEKI58NozEUlsqGdTdQT8EH23jQAvxMC4WesvArLgh5FjHZTk97HB31ISXEN+dn3nnP3JO7m5
3jnxc25T103kxWb9bDw05mBVB/KVlyhbBw7qR6RZgrBJrtcYuQI001azy2klsgT5RYf7tNgvV/vK
hySfFBLe0/SIL7dfoWXKz7aimi2GxyWD5j9902YqNf8cnthIA07m0PJoSkdb6bv4tYf5FAbJlGy1
rfWEnPv4Xz2rbD2gn/KzghOr+pL8DLBLYaAYOtvOwL5pJ/6JIUWzHLi4GeS3rdu7zou5pwRvzmZL
DLBm025og1Et0e/FjBvP4ww5WtuCzTIiKfRy1rIf9RgDCyENSUIMUI0JQDPvgGTIGsQzAOowzmUd
6bI6RDDIFmWaodrJn7CUff5HCiTHkxZXO/ec935PZBCliFIZ2PngOCUaOnV6AmKCMBF9vdUnNdJY
cBtYvPJrsFf5uMkEVK7qvoAXv/3SP0XKZdwGxx+Y3z3NTt71krmEMZMUR2QbMVOscwbB8FLqyhFf
4J98LzorcriLpDlVbHLNfUKkS0ZxDFD6COAuuwG9Hrwm63yCbCjYwufBnCnde7mduKX/gdiIQ8TN
o61t8GyIzil8ihIekHsw6AMgk3QjBB78jrWRilmfZT6LxRVSuI5Hthxz1NOMmnJfplGlI5+P3yBT
vqrl9PxmxPovrVKQBH0bJgViO5+e+QvjgWagF3le7xovkza9KfLS+lOI0WDwJU3FLhRe/lYWwPFh
Boj7bhenFZf6zyXmp5o68T8gtd4OFwDV60yG1VRsqyC7zqhWFNA0Abht69LmF+uFjnzzuKCfTJqc
qLXczd8ENf8GOwH9Tq4KJ59ROvoP4LW855QGsszvLVC6ogVgvP+BFJXAh8hf7ijX5SC+huk5B9VO
aI3NtPHZX9HW1u23rusWUHc8KScyf9ius5CAt01w+kbAyURiTaCn2aDUMgnSNlkNQ4xoYA+M68s3
d1M6XDwULC1tfN05+VwBbsuKen38KD2Pl68lnX+BoqxXiO47WCWnCaB6l7oxWlkxLFKBKwZ5Hho7
4ixJf5wwPZNowWjlbcbztKgRSwJM7hw+GR0i6Ez0GbI2Y0053aWQVrLH+56yV0PhJAOK1KpwF19F
Wa+NZJ1UoVFmG8DWeRZrjWmXh8IDvsJJ0pCKQJ6l6c8XkdiPP2hudCKK5kMpS5mkJx2BTFWjLMW8
Cv49Evcx2tS+GEcSMR9aKP0svdi9umdAurwAI6l6iWGKT61KbCMf9pCGzBxHLq2j5Y0c6KhrBo4J
X+DlNv+xcysumFDKHLmEt6MwXveI7RwIHRs2trCg90+1wdp3qEtLIPhIKNIqWlFMAAZd5vtSn9sO
2dyumQslsusGXTFjpyS0uBeM/PcZjF/fnRSpuzucyl9ToY/jgA/xY0Q+lRDVfvl5dZtISXh6hHy4
Nmvou6Rp1dr9CALyaxOUrSvunIF0w533sx4e1YAVRfk+HFPhfoJUc9euDSP2nSOr87VgXbOonkEx
v+BpfS3xEVsvo+tL9dpm3S2SLF0Leb1GZ5MoGzyGWInVS1MjPI22uNkCiKLyHWQLyZG0NO1RdqUa
bIA6IsyyZ7oC7ZemidWU3pPXVc+ZPGhzYa9znMTx6lousVvt5Yw0NKH086ORGf7wlE3z/OdIFIw/
7Z9/dFw9yjUC0jCWyG0fwoZPEENiPVOtG1uN4urtKQi0FoVtZys2UYemgrrwG0ayBJpJJhmsSlLq
VAUnU837vw0BH8aPR47BFjJpFr62gmwc4LQuK4wOimVPJFnk3UdTEzs8YL2zG8FLXBfq2SE411kW
09BKbybUp6s62kS0Xz2wDVHZNN85HUZrSTKbWIvqMoDaTbInvFsfsoBFDKXKop6YOOoitZ/T+50j
SZJxmY4xqEV/mQ5+Krtg6ofuwnE41af+6QMNW2yVsf21HH/GSeyjIcvI4+4NzZWsOXjTqq7j2CiT
o9rYnb+ZgiiBEXqCyHpqWaBphdR4Gw33oepi1dtQ202x7ZX7aTApcgau81HCWcNUPPldjFSuzTB1
ZcUI/gIAEGN/AuRt3xxAmrcoxIbpEQqEVNjwn+BzbtiaSTxDKhUnzE5EYduPpzyt3zc17FOHQfsd
rPnFDf+u0TPK8gOps2M2UbYwxPrPxJ4+SriSHsuD0plBjkuDFjXOhxPCfKxXMNrtZ+3HIj++0RC3
sR+jIjAnHtxvGqcOE2DeJ9/GOevNc96nAhUK2iIBKUYGde5NBycbICe9rUjUVrzhCr+/0EtveK/j
k03kWY8Oi3b1xMVd80MqWbPf7zWpeo9MGsd2B6EtxgTYk3YTxpK1q4+g+kVSQ6z0VHeZmZ4wjPiy
29c8QgnjzrXwCsbGmfz82pQrNoUnxUe9g9ZYBjQM5VklcAa8wg/BChkf3Ksy7osn7fLhKsM7ce7j
toBlkznALlLVvcqQ0hdDE2oV5oMuaWyRy2XETKg/sugagt7skLEzskJpVMTraI5SGSLNyTcUfx0U
YsHohWiLsxOjs8p6JnxjrN8Eje/8Lv4Tqg2sCVQR0JXqqCqpNSw9UsZxWhv0CkUSg6nyF/do60lR
e70LLjS8Pnk/eHXN3z228imyo/jjgFo/PAQewNDM1msf2PHz1+4/bIR7U2fuu05X30/4UpDZ/v2F
VxOTJugtWOYT8Rve0sQQjA86Mmr38wPbHOAl5LOmovOU3505ggrWB8aPyGZBatvJ06Zlv0bY4eMY
LDl2Gug1cBAUDvotwhWXJcuylm9rpcQjqbMTZ84R8CtKoNKoclvZMMz/8XC5wjP+ajTVxt3ZjGC6
Sp5tjO3M4GEy/y7uk9mattdqYkR+EyUwRzdBDwLNFk0PJiqCQmFYPKoQZLp3/ayQEyfzd0D8YZTB
dfEVSVzRGaMS9yEHocE/HJuuIF/mNIP6A3L8t4IfPySsJtgsHJQ1MxF4W3uUoWazmPcWFfvR1FLX
qeALPp2F1PmrPya7xYy0HeVFfB72q6affRBGoRUmXGvhIBjTRH+vYfmCriQXGvghMNWNUpmu5GR9
5EijleHcQNFjareJqxo1eEXEWYDOkww8SCkZcnUIo7s9Iu8iFerE2nEorz69zmOoitaFO0G6VuHM
HR7oXwyZT9ucAyE1gTj+JNh0/Xu/VpVd6D8uXjR90LU/2XyjyyFFurPfxufd/71FJ12ZVDnWeanw
OgkM8EDpBiQB336hrxXzBVycKAvjDoecBLycMDDuayX6uZPRn8P+BISBx6r5xTQ+RCzxnVJoLPIn
FsDaL4mDfsWK68MHGVM/ZYqyV+jszfLBewZD95Ob5ntlMCwjlT0aZLadBvm1DP1T+JX2QtK3QtGY
+11CpWgr6kYzgMi3HBLFM90eT0rx2qWRl9yS9r7CRw9v/gh7OAJM2QUGYjmkwn1ftVcX1sF88aMR
RAwgD67sdARpdx6wwXf3hvUhA0cdBGev6dD5F197bWwNNpul6ze6j1OodNDWpdm89KCk/Fop4Fgj
szCADNyGG0E73ZWr5j67MrjLuY+nTHn2nvGypL5jmCWzAG2PJH1DZHxqmKoftHPgP5ZwhVYOmbnS
pG8nOAy1lGVoWesVV+ST/CPS95ozl9+0SukcHDM+raxkzgnOuQHW7+zEr8QonKTxRNScE5td8Gvk
bVQeyx945PnPiddhgbBEDpuLhosD/TNsW88AZSyOfdy6cirmfA/0m/M0JvmDc1/5FI60CZOiatGj
sBzQilSCKqVdRfCqNb0c0T4OmwAots8Gybcr0zRiKtrrwiOaYtg+WVopQMUupsofp9MAjZotVsx0
O2N4ArHDcHxwGQisy8rvzJzpPlZb+oNbdGmuWHZfMLYIO0cz8qKAorVJc27gTq+f3ajOUvR1nij2
u9teVz8kdguCnBYBGZBtkEc1UT7zf2iSlKt3eut54TpG06pj2uYsQhdTjrglWAGdgfv1AYS0t7XB
KCdtwY1bRgx8bCnbNLqOkAaz6obFgbT4UDXJyfrslzdwa2upns+uvQjyLsUeF22/W4mbcbO1kG4d
Hk13qi7myMG0PVap3CIj8uLekgKy0blSnzAMhxr0JCvqFqpZUYhyVvd1JzZ0IrgdkLqBmyVNN94W
TydMZpL98LMJ1aTBRUeAekkuX6pt9P7Jj215cxrVaqUpedr+ULBXRe1HuWTEjRmraJnIhmrk9vgG
08r3NKwWu1fpnBMG7AH37+Y4tFhvTnWuVYxs1mvZIkz4yb2rQXeWKZcv009m4WQk6P7KeGs0XCjl
GPQ28Hay7E1qRe4A5EetDmTWafKLW+RfOdNPnn0Bab2D1/N7ljjG8+zDWJWVuVX/JP7yQ192r+en
VvBYFy2edpb9Mb4GuLTEUAk3gTu2Zg4CdwDddhIptghfars2U/5zzrH7DGj34Qt4+/V3uqBuS1E4
2DouEgcGgkx5woiRofc0D6bAY6n6cW31N925eazsgfS/MYRAE6KFCzDsVk3a43KX6V7uqQlaI+yY
tOIDEuh+jX6r/TEGR8iCJm1o/71xREGbgiBwkMifI+IR47iCw+eH+ondIuKrNArxZeU69kOiVpFM
NH6QbPf1CIBP8jDRAaYRARDlq6FnHamBjIpM5fF0PE4bpBBbPDGOgDo+0NevETotyOHN09Bg0Yog
BDyPCNaaI22ymh7D4nhKABoYC2IlyRQAoKxRDL+jQ9FcBaUPIdXl1BjBH6CFfIgn7fwzqQJVNCNQ
lQXmSgLKrGGn4gcM8PsGD3FvriTnB+dLBopASBhv3eLnyl8pSt6uTQ5xwQK/2ZGy6Wt4iCSMTwQA
GrasMhyjPggjkEIlXjrJu/cAbFxUt9YCrvp6JvSyWQkutNIkkymI/SClmCkB/8QEgASBfBwNrWRZ
TipjJJO9nu/upHH3HV8Rs7ODmgP85JFpGewBf1JzhKWCBsiJoY/Eq0fmVaT+2yTDfXNzkq+S53+r
g++BNg/spp9gS4pxn2c6xE8peesfibYYTYO1+Ory1Tjbmuw4gc8x+tHKsguJ2IfHMIJQh9bXs+A4
/RAMoTqhExyioYzN0n0tjGsNZZmOq62Son1X6OVB87CZjjgq/IRAeKsLOBAU1Vn2veNVHhAoWCl3
oUR77LklDRcOiiX/UuBy4tJdnU/5awWpcIONMYHgwTIIBJeSkUt56PfzswXmL/Q4GoEHbFEfMaAw
pd4wgJWgq8c2yTjxoVzViHdezXrHzk3LvB5UjYUBO+ozcn42BnUBtmTjcpRzBAiZSC3cp9wGGrJZ
KyQXKcssVBrPwbkiBkd35CQhcbUpX1eNFdRSb0g9IVF11GAL93r5ZeG8HFAcnTIUEwXkZ+/9586D
PzbYTXtqt7xDIbB5xK2pBDVYbUTxYYbUJjbXguLUdU9V1S3zrPkxJX6qokybFEfyQD3tL6PsHnBx
STMb46lyDV/t0EFEhGBMf9/PI5hdmEgzRcdXlR514YPKsy9MMqAQYslEqWzWibmqu0GuTAiHLs6z
ft7igOwx70EqkPn72m8Gmatxe0dFta+PH0YK1VPy1oQtWjIj32uo0aMkEsr9YUbe4876mynk9n5r
8J+SaW65QKaKsP6QDGdKwgh+io25gpWxrTv++5Y/4CPDY6rqh6HqSnt/ynUNZ5YC1QPnjH4L4AOt
S/FEeHc0RHY7Xc5/j4jRQ4V3z3OXSOh1Z3j6YlSyHb5y+rOTs5K48HXeEye30pjyPcjONqp9uoa5
E8LbLjWW8azeekItKl5InKq2sGQ8OHZ2qCOJ0Pj+V/doMmj6q3hHrd8d/nohx67c+J4D5wUgSWfD
bwicofFbNi57K3bU8Z/fu+U6IyhXdDdBLpF/Dpkpy1mS6skNm70YexFJjlMHv7JoMLvrhesRbww0
lCiuyLZvRhbyBHBEeW74hkIdxJ+2jUIHEKqgJ208yS1uCHwm9UV8Sg7beOcQAHgekC5XjbAVgGm7
XBI1am+HPhrapkuhnO7sHD2ZZKPm3gmZm294fMAuNh/mD6vGJIPGwywOhva+O9Ej6sxNldD/B9CL
nfdDWqQQQg6LrgrYgN4dwePI3KXjNC0ItHIQHzQPGe9HAs0qF/HtqhROGv8+/hPLgu46ojxGnHwy
8MuXd8Kk4vRJb4PzXms+dXHl1wbYzvVAZkVhkueDVYUer/lRQOZuvRqsCZtpSHLwBQguQyo4G9Wr
PnMorTh+IVONzw+vg6MB7qmxGfcnk/hEEBZd8CnUJtmoF+vh5IIw83ROPblXlptynl3VSkeDCgoA
e5LseIJoooNcbwlGP6ZzElbfYJkPO2eoKV6TGMgpt7hqV0Hl65kcCBeqXcimhbpe1PdUtgoaROok
DuVu51L84WMgyVV9aj96JRuouwNDChLYipV+VdeQibCZ9WBE4utHzjZIxSMuY9O0XtzzEskWqwcR
qNv756v7nfqQ0w4L0snJ9OkrQ3tyqI1cdwPHzyTHERhxgO6t0QkGOKwzryypuEOo7G2kkSoYo/gk
OQf5fOXpoZVSu51YNnA6WNfRb21ZnTlkMp9VkFf1hZRmCPoVO9mgR7HjX61V44OWR48zHhnitFX4
JgfHnGansF2d/Mfi+fgr34fE1V2W0zyvp8GK0tmGQSeajBSsXYM5OC42Ffsq2YDsW1ZBSHWl8BWe
4wEuBJGtoxgzFpsxsoCOhwag61WUa3k24Z7GPHnSKikxB77QXba6/+8tppZpBRWzRiLXlq22uxnc
03lTUCI8yWFZjWpb+oLTMP7LYOCAm0Ddqad3N5bocRFTCckSc1mnpyr8XVNKYMo4di4kX50VH8RT
+abPhOf3A8eTPDtHdmeBsLLSEW1X6gyWuT+ZXYMPFqNtKEA6cfZfD+qWUR+/pbP/U/o+5A7QztF0
RzcxLXV6I/UJhL3C9PRHpnLw8rN7QuHrfdCanTtqJZs+bISW0GOkA846+k+A3SLsziN19+w57hie
RC+6nTLdUDjTsLIMiagRHnUa3exEAis4dckj6dQJAMxuOjJ8Kv/bX9/p8BKTT60JBonONPGIFd4X
L/olFKrsXiUzn64QJuAjPQs7lC9dsPGP6ek3kLlKK0o3mX5DdeLy6zYOH7tsdebxF7WUWtd7Evsr
YtuuR/uBqmctDkrmC5yolB6DKyvPjRfMZviTn/EzCXSrwYdDFZnpuOMvSSFsEFG22toVkAqQBqcT
JZ6DSREhb1aUM8fBmbNTkhhMiNazZ+9m/mXrnvSYXGgaF6kOcetETtyy65rSEvL8oSOfbUJ7E9uH
+US459jp4QyK9C2nwXKwJfxg2yn3Zn0IRzNl8vuzRVd/sMT4xd0PMzOdD537c4WYP+Nb+ivOKueg
ddKlOVGRQl51qYXSshTVpiaoXA8YCusOEEUqankpeUd700XCqkKxKqTFuXU7rZQ9xREH8tAKguSd
pYVv2LzmN9ttGKXUr5GHKWFXxKCRvVklqb3iNFYn06mhql6UXV9Afu46X8Ubi2axt4+7qDpvchlN
0JsaeLwfJ1BpBBtfzq4wNory11smXxaYl6sTAGmywdHFk8gwEAMGY6hLkcqxE/Z6LBFArkqcUw27
meU/oH0sssuzHY2FmCs6Mj0FutH6B/YE6p6Bfp+X1DMVc1k3QmZ1mkJpZDixs6u4LxnDK2U1jRTs
cCY0bzyapFbeT875YJpe5uAnokCvkdE3xSjPd1ZfL0Ge9IO3iO1Om3Dh172ZNqjZfVk9RiSanKei
srIRI/OiCXSQ9YAEKajnLsZFuOiprPEfxkzfLPqBYjcEiQyMtBdR/A27gs2hXwkfem6/UV/YyLlA
PDVfeuJmgbDKyRHWfEYxL3iOz0YF69SW7/JalUvTm8XEYDW38oLbxpgfDj7Y52BU2b4lKSsnwoQT
SsoKSccbfSQHpJaI5uq1aoIiDLZIlla1H6ES58MG1rBSQMYOZj9XwytA9Wc8HJmX3PrCmQRwvFOG
3RDDz9LSc9vYXujyknsLtHXIkOsS5J35B2pDuA+U9vldotrSXsJex+gQ6n72XAR1VyMlfwnDAEUO
JxpTCB2cg5y00LlwwkAfPEr0AWGDk+MXrDyb7CiyatmQLTKfyeUCPC6axk3yB/GGWIMhDJweU/X8
TPKbWbBKbzu+DO+hGG1vKTUBNfWVCwfb3gNVAKbJrSo0OInj3jzLVky+dm/aHxl9Kf/EIADWlvmi
ay0gtx2fTFWTu3KDnBh/EMOJeEAt+DTwwMwSstnFCv17eccIkJlUnsL61ldLqT2KY7R1euoIcsht
KNJAB2cVTtMcYND6siALqN7V9JWor7J1N1nqpzJqI1hQ06VX8qs6htQ9l6uK7LTEJXGCoJjdCV7d
cX/GaMHol7UAY4ASgyl5/te/Ogfe52QRs33u0o+Y8LxlE/QXgOpdByx2/HPpbBz0/708SVv03sI5
XgvporPS0uzmJcJ1H+z2NtfgloiuSZ6adwdCcIIFszrypKvDvrHweIHp56SMts62ojSysHBtexZX
Xv/fSGjXA1KD3tnrNil+Fp/ZXwqYH1qcW+C0GV0WiWv83IZfZwjb8yF4IqNBqhWz+FyHGdGAf7+d
OHfeA3+qAZy9K30JU7nufHNqCTLDNKGmd+M0uGnpz3wWEqEq8MAXupE5jis0gSC21ilMu7CyilZP
1XsI8WgY8kpqWMxlFGP8GD0M5C1tUEazzKw0Kmur/v7YJTD1LcrK3uZTi9gkptyAuOqwdRfmhygZ
BBNkaNA7ucMwLEersQQIXPWFatBoto8cK1PN50OCOJHN15lFt8JFcudeOG8wtmW+QK7TUzmH/msB
xmfrESmTZ/YWBPVPkbwZwqsK5M+RtaPFhpF6uex1AlVWSGQyIo6GY86GqHMxLqTCC0H5Al4M8Dq/
UGsJYDBtES/k1vwI/Jpzt59c9e9WHplpVC1aZKK+s2du7zK1lQevLsJJUqEXmjR60m5eki3K0L3v
wyRrS6gxXzojpNuU+maQAZOOeZBAT+vspKTvbhvOXvs2TdQPE8MZf/Cg12XKDeGD8BFuQIzHf7zN
BCZMZ6d1eP4yjCQb6PKyWMyovRGXxn2nmn/RRvSDLk4WkXncnGdHbAd/S1vefgPSh0Scw18n/oaJ
2CX3KP5DiUS/Ne8Qy7A5+vP5AxAK/CXq7GrUDKrh8wwwPhIrrSsEx8ijghVPlPYpQuGedhWeXz/e
6UFZBetyGsukjG58POnX+69HpadobQ3SHnONfmvz6CPNSl+0zIEDQrudNmYw1L+NuvyemRpwulQo
Hxj7KCsCwfRuQMaKiSqyeCkaFRDesbQiwORIy7aFoQCfso4aRYlbkIozXBFp/zPLA4rBEYMa4X1V
0pG+Q4kpH9/ffYAj3In35VFHhjLninCdN1RFzC7TzMOmY5aMyYH/bM2vRBtA23+FcZnRRtlucnC7
C8ceRYo3vBrPXjbaks6av1SXyUXssrXltwwz3UHfhkhPpIyTczm9PzLjAHj8zUPa5AGB/W/F1Hap
V1arbQs5kUgIgCYaFDvgQkIj8SOTO+D0s0XlRzge8bHLLFn3eIjglnZ8V/Iz65mp2cF4K/m0bBQL
7LDR3rKzfb2ZWnlUZ/fEx6JfEKfbWHafJq10vYajy7ZKGv2lNTDC5OpunLsAScAS71BuVwuah4iY
Y77hwYlSm/UHQnjyVJmqDH9QVcpc0mqTs1qWenOa8x5I7iJFPZnZsFvO/xOV+gp/2wVWYQA7yPBu
K8Ztu+QQnXptGApFJWCiiaPi1bj+nzewivM7m4lblaTrGgj9yT/qtJX8wfWbvqfP4DY2U6yQDi1b
jBTmQNftfeLG8KwJHfNtniTPhUP4NVhaf5O+B16Zoffp1elJEv/MgjqZ5EvnRAX7hAZ4pPJo6Y0h
5HBdvCT5FpdviubkKrpwH8Lmtv8bznOkS/3UfQnsffXPvtGYdexU/i9BfJKUva8s2FT76VR7QZ4E
Ogg7wHS5LNCEtIP70EJ+s2tPawPiuTGzPFPv2JbsHoHl90HUoySEDUO8gFIKQUxFAAI+kp+qsVaW
drWwAjpbtNXNSgdZn5gcP+64S1ZjQUOyNQSidWc5uvpfJqnYVD5tKqVnoRAjiEPKLcZSbj98HAeL
WMeIoCiuZeJdXeppCLisvylnumEEDFX984hfTxke44ja0lPL7ZGyyUrlcX202+RoRUYU1ZTRa1iK
h3caEWoh46Xrpe5ZHw7RBzNRd8+2Wm47EwnGbx3PApa5ZsQr449BosPxUaDG1yBVN8zsyg2zEd7t
IFid/s4ux87tG90qH3x6/87E8qR6Yn5+cOe5KPGo6a2kdmPc5VLDinRqaR7y5GZQFQqRP8F5mGkt
eFRkmL0IghJK8P/SBiadQrGqm44JIM7LrOeG6d/KzaAqboC1rz9mWTkGOAnFlpV5MywgxYjjBEgG
UB8f1c9bhaXUP+voApxlkYvULooUvGnbkDC2cxnTXATHKfsJQrT2qRgN9mKNL+J2IjHw44YozvcQ
ApX3I91axCsM9x3VGkmCJes2I8I8Aet2T62KsvVHKkxGPATW4uGaXD8v8VVeYPb52sHH5Li1QhqK
05cnax1A5c5DiUpHni9PACt3/yG1SNWBdOE799agT4FexwzYhQW3TvDeWttYBU+2uDRl6/RZUhwW
yLOQXM/tWgvJgtnBTPZm6bQVfrViXnP4cbD/gUyMuaIeIDWVB2n9gR/7u/wD0EZMW/l8QTgy8Ueg
5Ok1mLrZECi5BqMyUF3HWFb5s5hFhD0zgbIpXKU/kqD+EXRHC9PQgebpn6IjL7kZVgHmO4spR6pG
2IpvznKM05gElkIsdrj3hZV/4X/eIJOMKFmeAag/kTMJBS5F85T4hQ6SUlK1bqjJNTN38SaFMPz/
jZMdjooFKyuUII7e4SGlkaptN3UTvrEnkRy1ViwmsZjG/Yo9xeBEW0jixwai0kHGHhJMCp/beSn6
XbxsyCdGLDi4uWzLNoVpUegrESNcy/EdYogRMhX118YhWsj1YOpRcXfFeSt6/ODkaN6PCGy9AUAl
3BM7ypx1t1XqmJlx5dai/P13s5Br2VLL1cne+HfnWZ8dCfquRNGlKjDgX8vt/qyPyctwk1VbsXLU
tdF8Of2iK2MNzyGMlEj89zLNn3TtY4aKScbz7PpLl0Z3/Sq3xAOBkTISazUUOmkdGG9cYqxvjGjh
z722o6QC/WsO26KMCMqTv/Af0iFEKkgJ8GLCpDX7/mels+uYadpgQw+qpOFz4A5OuYIgTmj/rAhq
TIh41Ld168ItnbXn5EIO/Kfc2w15FK2jmsPIKaPx87B8VUsgYQiOslgFY1gcrUKJNHAuHanzci+x
K4lF5Oi5liWH1WZrQUIgLXXbCADcN2wWLI+0St/WqlRcsw5eGU7ywiEKVTAIGg6AwA0nwRjP44vu
Y5o8jln/GEKusT3F19ylkp7ezXlRFW/j9sQKoWJB5C11dCtiBnQ4DP05LAtY7Frdb0ZYJxrGZ09V
P8JLhvmw+KEb56DtshlQFM4rOD8PFdWMpwCk2+a83toNG84AhR5w05hBY9eJS2gIqBy+JKMclaaH
ykVExdFJntB09udL8bm3EheKppgx+We4+rHmrqJ8IiboD41ZAmPxxL9dMIj9wKO2KaP6znQS6MZ4
9y6qri7LruCxMWUOai9IHvrlOHzZcPkuX6h5rF+/mBhnViAfCNt51x2RXTHsofD09buFzYtOzKO/
Yyg3VIwVSUa2aRdG0mbtzlmHcxcsPj0UVISnybF80y5K6xPjvnZaCui9tr7i2kwxWbSBIhgEa0rQ
1nT3dMU+yeShtxmF0HMM2tZfuW9J/WffEBzhdKJf9v8icD3Un+JjNSCoU6TTYoHI8AOPzd8DuJEc
qNlA1Sj+t5koUIw2Ilua9HF8rIH8zZyi9n4rjsEKVK+Gbt81Jmgo+ykdVJx+CNAGxOzyCMHDClPY
cdMkU4BSzPX8JrZ407F+hnpC2a/Jo0YjvMwra8GTgkHQnhO5zdH6VbeMTxTvpx9nzo1LcmknIf0L
i1Ud7FPwC66rYgZ2G3Xx/fiUEjrFuT20dM1FTgRPxYnmnJlCKF/pe24Jqj7cHG7A42mLSxy5dXhF
dr+UhJQxUX0OMyTc4U9ijljI41OgGzboxJg9x9v6TjhknN82odIE1oKqlwJpHSGGj/zUXdBZ6xqx
F5hx9ULsrG0/Keaa4FuFVnK25BdSZIWite9XpO+xu3ipPzfzs3tk+X/BK48RwW0S69CNP9jV95+P
y2dNv8ILNQeITM2yPpl3/y0HRmBuMx/AioBNYdDM7XFflgenHp3e36s3knedYKjDXF+1K0baf4RH
pesylIL9oAjqqeKYijRrlQNV9KRfpD07pretWYsIU9Ykl+9HRMSg0K2Lfa0U5/Qe6DVXPGk8jx1r
D2ofdVYrGiGxMZ8TsXo8jRQITsUK63zoFQQWNwANJDD4YJsK4QygwBlsYAVZllgXVhcmZe8d5Z0a
xfVZ63bOlTU6jUKjBDf4pBhiEyafqT6PFJumkMlftJSWunTegukLNhxhpJmGnR/iDXQzmTKaV8Q+
kHOeW3lnbKjwysoth6Xlpm/nZKkcEb5c6WIrHSznnFw8gJ0bXzzLJ+vPnRXxlGk2fJ/Q0NxGRZUp
kP2a2adZhXgAyeed8L3SHVqJsaZTlgUGHdaQCP2IPV7aCXCSnasddPWcHRzApOf+uaoM8ybJByRM
qGcqB//TsWmJaFfbcLJcRePv1Ps2jF4TCSm4g3XbvBzeoGcentLQZF3AoDYRCBrTmIRA7NywF2wb
6cCIGfLqz6yiJE40y5rnzIxFgJMCPbKsRCYyiwqN5tm9P4dbwFv8yOz/HI+9t/kRWgNHtwKD//dL
flFftwgMBSinZMx19Vk+XkFEc5orVwg/L1XnbdDQNw3mRBJC8dnPQO85CzXozSbX3lLl7Y/3ny16
flBUhKPnqS3nQhI4+VCCc9WUKgYlpjqCBF/axNpfm+JncJRVb4MqaCcEkfA54ZV4+Errqicbo9ku
bEM/AQiTpB5PVrFMG9zLH/rlqow1gsvtxgwQBnchM/R95IaRxUQoKPb2tfvbxpZ2sikzt3B73C6C
aWOR/8VHumFtKTu3qiC3k8QPYcSsy1zGZBh8Bpwg6dGeSQvtrgmJrKW6iXtVk6/WNjqj35Nj335N
Gii6fXaftnYPr91GQa8196liZfyS4u0UhzE1KPxW0O6YTQC9Yb4MmnE+/FPQS72+qBEyheeZF0TW
+ACuyTepsayjbjAbamX7/W7uwwEvp10FDNF9u+OCHjGQpaomIMi5Gh3GU1pIuFirWLvgDeTuC35R
UrX8BFK0Nwb68fOthKvHyujau+3nVjaBI7XdhYdlEdDBIfMTpi43QP4seqU7KNBlkNZoMvYHE7z9
qSBq/fOSUsoI6f3KsRxdUClclPNw6Jf8Vcld2WJPbY1SzUdErOWNYSx9au+oBXu+p7XsSKlXO+IP
/7FnITc6JWRAQrH/Vi2lU5LB+il8VDmsVHWZWHvnfnrrvnpW4/D04GkanZ4qmGSNTQybHVTpaaDs
E9JvTP2HtZEYPlajhQTffP1lLMfPtsi+q4Jv7g13wEcpwkL/rKkCZhOxoxhkLPJOVLQ6rtncRQm3
q4UqxM/IqSia8175xxHmGi23Qjt91nHzJAeWyp+IS2UkUnmpRPSpc5pPxzt5XwyzmubpZahJBgpx
g+vroQI4ntdTahjYt+p4qbD52Dtkb+4ELQiPExYcMb54szd7px984hmhcSBj83begDwwH/yjOuJa
EkqsqoKBDaHO8Kim+VqeyMskBsyfLL4Iz7vvD4LOaCnzSbAzhGWsV7LBiiGMp9CjN2J5W0ISqvBN
sYqSh1RN+/9S6TJ/UKzEXfL8X+nX4gHmkUU//qaQ07w3qza7Dwd3xlym9uvnqufFeJYNhyQz1e1G
ECugZYipjYOWygvMY3NF4Ttpvo2T5c8tfjDjMrx803gNyA9lTke9w8NNnnjhDxpRZ8GFMhD7dHxc
+okVdGsSuIGzs6erD5BrH4h8Fo3fHHhG2dopwYQtc6uDPurjbk1zTzLLcrJd4X3tZ8MWdbowqFz2
L1q51Mi3yf7D0mfRlvd6H/f4W5kfGrneAeEEY9DOf0nwVAmXAlbsyuDBlLwE9kYh0J7wwffRZeLt
iYpDJzzkA3Rr63BeSfwL2TBTgVrgwyQMmTWotgd/gBr/8pN4jCaTPuFdUGz/Mo4GEP9uEdv/uibl
dOewcumPMKyo7BEC6O2G/LTVpETOclBuwDQ1mfD72jvDCWD6eQ2xIB7rEcYuj3kLTlqpWJj2ntAq
Ba6KYPA2NDvIx3lpjtaI4Kr8RikaaRbOBZ7xTzxID437ve2XLhEYY3TI+nkTbn4jSsZC3beuCuU6
VPX8m76TYYM8YXG9ZiYMneLPnTxunOK9mO5M/IujVjsuIxIUtm6PzssA36yvQ11QB2Q/5WKizn3g
0NZiXUjFwsYvDuFnFpcxALFl1nHN2Q1I/DAw+vmiJmBddnH34VEdBwrP/fclDQik3yxlQEeOUsAU
h2lkSMKYMw+pBaWrAfRsIWqKc8ty7kX3cGTX2ufxKHj7pFvMLN3jfRVGUhYRpcVHp0CMwLkkusAe
Ap+qXdcEbxmDMCogvAiEIl6eMj/qEz+CgbE6RD8X9EjBexgEedTav/Jjlo/4VQgnhnYjq6wFgOYP
5u7JLRqOkh72UZ+AEv+RRalpwke8lwRxv2ESFfQ5aqKDvIUCxO1wCMfPVcxxt0i5vnZGGoa/a2MU
ZAXRx1qkWDiU8przbvra05vKbmjTryO49H5CvvFd6OOH5ezF5PUY4KwUW+xeg8Mn7qzK/6facXHz
VZcXbVDx75MygNl89n95SdLEZh3EIBhNcwlqbvQqUR5flPn/Ad98C/ZKnWYKfqb5OIXyh0uET+ZY
OES9ll6I2sQrjt7pmQWd/kxBUnrTrZcrZ76S32T5tRwCCm9L8WO3Ad3jMuzOYY6c5sxCm/lagXp/
s7g0B2L+aT0KR3UjYqRMTaZUSCgqLq2gfKCQGcwEeGHe4/hpQU3Dq5l5H/jijBKV47SXrtuNvyq7
f1yWxzjw/hAHdlhCc7TvtWty7C5x34uzHYXM4McyjkM6oLzA9/xqU1jhFSIgbt5mIfvR/APH8DCY
/YxFEhkjzW792O5g9IVbroKNEfa5XMTeQzp1tk0tee4Wl2CIXWDy6gP7iio+NZNyDVENsfWsoy63
SQy5eDa2c5/Q9XFarRqBP0VjI9/t9unZoogH97ctgJ1+15nKQbJlzUqe5S9p2ha91mSDE8rx1QAh
u2hRB8zZ1dRDIq9Xv7wG+/Daq7rpeQVQAutPOjkekfGj0siXjWG91ecSRnAmgcnrqtTaXflDkoWw
6fwzKv+7lEM+FMWsCuS089hUeTmjdJMi7176VXiEb2/YW9sXjoA+eiHmviu7iLvBQUGcL7sg4uBx
egrYzijPKMq8v8CosuVQqB7m6NgHTbxbxXRediq2fvO8Q2rMoO2Geb60/2OcjeFQuCslxnmvEyau
/AKLR6kFggHD/eNQeriAjskInXE2qslB7eNYtspR1ljDca2tCXciZGyHevbH+wV85duN5qjNLi3B
crW6QPS2fh0FUSvGz6xu2qgn07WRwca94V2cL/1lICEVhQRYZ0cSuQE/f6E0VWk4U5K2uJgNcWz5
NhSIzmv+KUKNKvuv9hERAWBq5sGXtXr5Ox8OXkSBdJVCNIKHHLOzaSTJRInA5n68B35pnqpKQiGR
6zXHi+w6x31pKP2OZfAy/wDa//kpPYqwro26NI6E97kCzP0ot0AUGoWvxfpuYTVc5ZksyI1ZP+Vz
0OKJ64QJRw+55fusmoY0lVLbNs+XPIha5TnrcETAm+pq9HwAqJyinX7YhsncnTXwg/ti4pbChkey
56zc7qjn3kFcQH2WhJyOi1rSVVaMQNXOxaIGyugjstNs5q7kF0S63t2WJTx7HFo8VYnOWN+3R8Pc
9sHZQ/n66tGr+Ax1dRPwf2HU0FY9ETImzZwmXT9/r9X4lfJPdwYOxo4Dr1dhoFEyBqfUG1dznvh2
iSf6s/Yiz+Sw6XZIKQevD933RKd2LuthK41ENumwIvS+tOTdrqU5ufqgOICXqm1hG9j++VBmDs/0
em476lAFjvQT5LuVYDNYlgozEatDLuMerCgn88mmUAohMaSeWcZ5V1qEnfYhuen05vGgiYZ94k5A
9rsomX4HhgMsAskhepVly1xi0icBB8HHT8gjQXcJ7fyACnqd+V3Pw0b74DMi6imW0Q8oWk+Gz3U5
9nK35b3luVhjvwbYCv1bIUxpJIEiHtq2A99TZMVrM5P50ghAZe9ero3dvtKfEyVLe5GrwuWkCtSW
9oAJfn+mOtPgPc4kgns+pQVHCA8SVkIUseWYCeyF6M+dLt+VBdR5G2aXree/ATUgzX9X9y/AkY7P
bLSCAa7Gvi4bnaExjimsquGvahqeDhvcRn7WCgIMm3qyr/W9DukefyFQj8YADv5kwEr+nsaYx1dz
XQqzxKWBvXSZwxV0AU5DADqGoLvSapDygHWYvH562/cfkCqtlztdBVTmMoYTufVp45XunYZFcn2N
ZaeQrIQqEva5X0AmsmvSYb8/DxwDgxRJq0gBrS04v+QsCVn3aL4fuGwxH+Q48ly77Z1/oIH2vd28
XArlVoX8xQNvM1McfeWuwA3Qr+IsrJkIJmdGTR440Sp5ylZ2oJSr+xrcBxtwTkuZld1PXENDjAPV
W/nxEXU5GC1y3hKnebWWc+OH3lKHm2iRtZas7+Nz6g1QT4m++F48VhUc4YPy/Jt/l9C634WnVs/O
S+1Gr4ca7o4yXRSbtAopJ4Ib3GhyaG8bkRjeGhmZ71Ns1TT3UGPt/la0EbkFWpKZ3vZ9dwow/M1d
H/5DoDtq0Tu0CUVoFjLiLPK2kTYTPieIN4h/0xqY6CdzGT/Za8/Im3+PCb/YOr0+Y7gjtXkPAqA+
9YRxbGS7lUCaKphuTgGLkHReyzXoeNuhY//vESRhN9vCog0x6rTxF9K00q35dknN+2vnttTx9yt/
EBROJLmMY/YcJi54HGEXnKtdqclrmTPmQl9HEajg6e2bx8iwPnoEva9wrPV1f2RvGnuTHLlTaETg
CkH7Z+NSwNWIqsuK8Uo2HpxLIgPL/QxDfcrRQya8MktFbp6U0Utr376BKk7N9FFJle8xZ1FaCrvP
sFaTKPekCKPPFLOvnvlJHUjr5vZ6jVjCyUwM6Li3ss/vq9HZsX+3cKtjxRzB2hjDKtNI4ryNPdB4
2AxqaZIynPzmz5Nb7Mq4Alpu0f8MuqTNyNV37XGRWlzQrvUOdkhxC1PN9Yn0SWEOJenyzwukAvNi
GKM4dmVW9W7+IvzwoulVeUGmXbM0WkAE0GgbyUCKsFqPKZtgMl+5UW1JAICUXyjXiULjcTO+zAII
rFr5RXTk71MjIYrATRRIq1DmCXxE7qkaW0QCPROARHZWN4TY2cvw/CDMjTVEdLQiuAquSk/n9BUp
denznYE5rRmik8kzcZem6DN0BzRrgxrls3U/hDkVNdjRR7BuOIHb8WpJ8y23IEpxWUu3cNkRAkPS
uvWoxiM8sfeBVIeeMbTQ1ds21oJx1z5HA1UwubUcyhyeJ5HQ2SJaqHkQ0W4+IHwTwAwkGzJF7vt3
mxkNF2Pe/nhK1M/zoeLUl4tNgDAw9FEyTlQzl3wfgsxYQ2lNPt9nlA2QgTUNoqZT2OuGclMYZPLg
eyT5aadO6RTDLn1RIl9hqKv4ZM/3XV/TUAXDjIHZSFLxSaIiq1f6gwxzyPgIWyH/wvIedIp4pcW5
FXP5vAqm9KrcbfoKfPiqSDE2GaPirNQt375QCHv5IDbPGKkiKV0NGyXBLcr5yNiP+QG/0uNmp2W4
dw4vqg5NodR1nVNtABgpJJVeHza7JyyQ4vEcMldaf26m8GxRtmCjeVbBs1fsQ0igAxWmw1NKqYWI
/Q+mn3dgiCwN+nL6NuYfC7dXMZFAo8ZVD7iLGb/SdmCpkMoeWo/d6iO5xv7VF/nA8sYc9xb0MlkO
MdeF21iP1rX3zekWkwVYv9J8VXqBzfMBSLYTO3RYUyWFFKmPPsr4LBSAQbIYO3fx81wbCuMgkMrm
aRFrm/wEM5sSLt9xzCJHBjGkUb3XTG+JQ8360RLo6hWk8jWc2rAxndd0ek495SCVE/MLf/IohIQj
tcTF4cVrf1yZE7ZyMUJ51748n5HkNbPyVm9t31t12Rg1X2kINisLVZoj6uq3JTwbjuQWJqtnZ9wu
QmG4DM1T1GbuvjdiMOLG2Sn07cAaOeapjPCa/KrBUjgbls5cIhUAaw8sGLjK0dqtlc0XZh8LzDzW
ASLDbzo7S0LNeD0n2ZGZ48t+Yq7CSBv3rG3AymlR19ncDDhFdeveUI3DMt9BETvQM4QJFxWSK/JP
NvcBI2L57C2yU8Fw4RFrf/BZdNsJ5euXnekxM/RB1YmfUwSMOOisFPMI2JsW4TWDQ6y03e9pEyeP
1lk45k3Z62kl2OfgeoDTVAlL4gbIEYeT786H79Y45H0J49CPrr4GgVKIjyRTHhPmyes7jB1+/49I
2JozOfvTjsrThqnvJO6pHL1VmenzPmuFy1Vv5zytasu+Vtg9FVpBMZ42w0faxOz7RJtDgUWpbXl5
CHdY+duGrdQPZqI8QvVj1DHeEG1/WkMR+9rXDb7vwpzw3GIYXYw8iEagtikao+CBM+yVKqB1YaSg
P18h5rTFxdpq49/0dfLAQIa/ox0jW3fLLyIyW4rvt8EorG1kFf3rkHlh8kQ7Mos7e9wBvq1QD43P
SHEYIgEwA3R87m9wgiqQa1y2G3KkxIHWcPdR/3rgCCQn3NHcm/oVraUxWXQ2OAVDykEHTktJ52Y2
FVAUY7YrPItCLEHBginzt9349jnejJAOqpaXEooL9+TsH6L9TaKgCpH5gZiksq2yfrc+xxjvfqfo
HOT0k7Zj+bGw7YisVKWx5yo4DnmkadHCD99c9x7vJFyfSBybAXb0WsJyM21+qPtkNUabvsgIv8KQ
0A91wC9872NH6B8mNQF3AhFJtABQDA+7qir1Oxrg8yozcppkiOQ7/3NznOOJkqpfXDHhgqYAMnLq
huAxqAGxyodLWckCKgcvrJdUI+dhMZkG4NriOPCd0aoCpBp/BobHjWyHYwC9TfY2j4Brukracrvm
rmC4GS93JMm2u5CZ0SmeDhBNFCDUi8X446aVIWLaiI85pjhrg9ayMLkSoBcLhZ59DL4T38AEgeAp
8+mZm7qFcC+5H+XjqOEjVFjXvYgVwRVgp1zZsNBZStPuZeTcYfYZ5dji8UYo+Mo03RjGhBZKUkZz
02jIk9Jzj25qxSAiQ1C77XG3WgyGyW1XuVdk06oXOnhqlrE2Azu6IPJe89zZ+tXkEAy53PVtu2Pc
HdXw4HCj4io2dvGg1cIT0fXoC3FGrDZ3SiHtR9en1TMcy47WUz9AfRtlvn1+67HGOAkw83yx5oGz
lB8vJL96BEB+afoazk7SiskbOkcYqzVydUKY/Ft7+AC0N0S/2Zsry2Sm0e6ZXQ1QcfAfbQ2dcS/G
ZSJGBfVLKbnvfp1Vyilq947J1EpZzuTiCff1wbGS9cwu/2EAgJEKtoLQnCwizfnYL+ft2E6cM5sH
W8C72JO94z807hB0T4sW0uLoM7twX/rhEarTf0UPtp2gqLhNZPNfpUTSr4JHSwRNRkIk3UgTiGgu
skEpkQeTouNPuTWN1P+uqexB6b048uhZeIuUIK2bYxEC7vKZX4K2ymu9bPEsc61QGcilfN9P9mXH
AfNh250Gyh2ctj6+gpHxFVJd7rErKGcvgl3+Cdc3cSAS0nC/h4ZZWWq2jstiAlhlVpsGl86drw5k
wp+6wV4q2GMgFXHVRPCHmdOM5vCDRQnKGqM2qw/k9HmEndRFitfjLoE49fSl+yaGJB7wDfkGkECj
zh5erq7SvuQD71MOy3v1bGvj75RVfZf4K20w1fYbCE7/GuQjtbMGszmSilrPQiIVHhtmutYtVzWh
9yluDwKSr7aTFMPeTOs6FCe+ZB/iSayZ8RMmwo0KyRvInjH+syjKv8EP7cwmX1gY/NyFwQZYjDQT
ZA9XKByJixYU0kyiVJOaIqSrAdlc8QS1VDMyeIH8WhSV1VTMNNRNPryVDXm8aLdnUEXcWGRRjSvO
EtBHFdxwLTdwRJgvArlUKJy7EDfpAPMFpY6g6WyNVbYvJkp6Id7TDN00Rg3XnHiS/IM3V2ORrYb2
spky0hZ9XCD1X9Q6b9zRfj2QjN/Vx2W7PHeOHGAeO8C2lCOqOQ0cygVQZ1c4D82FAO5DKHnRC4Kk
Zf7SMk+YMXillfnVFAMXLFeVRIz4LCiqf6yXhkNIeUDKf5tK1hfH9sjF3hVk8T0OmEooPsJeRyHQ
PmKt63AUBLItGoPNny91NfseCSLfUJkqgKDPP6rr7h7hiyekaa5GeR1V/b/Q3wvghTOT5I0rHVZ5
m5tcQYW6g6eInjqhUhXspcnO42gH6iiXkW92hoRFa2uhelmpm2kU61wL2vvk7gn9qv148AG8ICet
ax8QL3czuvGG0JoX2BiwPHUDuGrKj+0LDoig3xJmbLSBhbh0z/QarLy3o1PBwsFUp/RJ6Ug2eNwL
H5SfjkdG3yOaPpY1S0eOnToviUQmZrThtR0/MxH/Cb4s8fCETi+GHfz3bq8J7If8WoyI2VlIuCKZ
FBXdoQEG99evPc5HarMjlWLA38C/tvfe/gl+0vORYN5sSQ7sB4qKaxL18YzRD4LaqDCfvFso6//Q
1iGeM+kdWbqHZGe7La+PA1s/MCgofJwfZ1T9PKlr91LZ9l1pk5TyFdreSxwFiMDGqvu8PLZ8ooif
ZbxS2BIsRq/X7iciDkdspTt0luwrWpp+QNheOZW4px/suADXVXAmzR+iQzZcaVMuhlcFn3a/J9fV
mK/efp5K9ivHghtjwSDdjuaSigd+eTlrbmYoNDL+b1vEotU/+8uoMl36vZHvTZHRIr5qYW0Ejeux
wnOoOQwr2oa4SMwftAP8TX5Oo0obo5zlO21/krq5epMQYyQH30TwPQLw4KlqaqGpTGImvgVdLEcd
jqh0Fwc433DTtFG0hpUT+6zVenWQwK7uMlI8/pFlJgEdMuAUoQ0vs1nXQZF1O7Ifh08jaFL/tL5i
siI0k1srgabeFqMSeDUXYb9bJKKULVg5rxsJmzgEC/oYiNov0kkQWzKn/qQxczagG5gcjLQq063G
bDVTGTMSRgtj7MUcXgxBvuABHbDIPof0VrBTpGGOfLk7LqR7FjfB2IHICPMpCJxr3gZtC3c4F6Sv
ycqTCKL6z2PeP5Kyo7azfTjS597UDBevnPRRJFdZFLPopFMMf685CDzkMqkYDJ3MTY/d4EF7Yw4G
LxEEjmBgaSAEb03eDaG/DU2Vrup21+wrCn1RsEpR3bJwMod6lrNprViOXVgKo0AKhzOCQNYW8MdT
lO+110gua9becXItacrqxLOXdYzAbM9QgIrTUd6IzG5N9VQH+SdlZbZtGH4fvDQrghQaEJg5Lp7T
W16wIu84bASsUW4NXZ+qjWk1lJUuLw7i3DP3RTn3+vI+bmWrQ6kHPonzmttF1iCm7p4czCBSEg3x
1goXFu9IsvQcwzmSUHh4wot2kjy2LnK2L7JrAtgs3AKvtEMlGhZ791vccsEHHuvK3nFZNqORLVqL
rZTz2JJ0VPtj/dNkmt4CGol6fGXV1UjobpAfz87Z3/WnBDCzglZOsWbHI60RUe4ygG2yeYVzxdk4
wtdHAYJlrfrdPIB672hrXypfy2/DIJi+CyBLmGPZEl0pKIWFqYF9sgLISUdea7lXt8I9OpGxsF8z
ougJA96UPtd8FPOoF4U2l9GJx4JfON3RUXW7OL2vD1ucLUv0XvPctH7jkYojMiOyNgyZ6S4z7WsM
zNnh3WvNOMWOQmqY1JA+6DtOTQpwoApg0XSX8z0DXVM28sShj0iZlcfjW/th18ojlh1Y0feqDJ/X
Tb48fUbfSQ/lVQ5/kKZIN+jJaqq3pbomxtFVlk/x2QnQ1W19MJLzE9U198r5MNFUp18gO1H0Dh10
R06bPKX9OdobHfSj6jbJbgB5joTM9dg/K7V2aY26GyAMHlDVqJPyT3+q4n4NhtGK7s1F73BLBlIx
JY3IKmyuNwHHarF6aIcBz8j+l96+pIbCEbeMI53OunNU98+tOVfqm8ArtbqH9lRmpdNqmvRVqRZ2
F89zsC9bKzCp+Zn7opq7kIGrt/lF2/HtDtiEYlhVMC8qkXPCaHhnqN50P7SbqrKacnDijtOdEgFU
3Z3EduFWjSYWf/g8wDe+Z1gHkMBWMJGafvWrKjB5Wm46TgkcEQh9Q7GdTx5obq+ALlD3jTkden/w
AwjJpNRl05kCIQWmTYStP7SDiOWaGqTQV4Njp+cbWsMxVM1yUyfINuqNFZgpKD15z0vEOVAXI/qn
uVC9/3YZsyA7tGNGMyQUXlxhwZMaR1lWL5ULTqSAz9RwzbWXNgpYGH7WQ6cQMWus7ARTi4bCSnsD
SQIz9aHsfu44IP+SXweTFpxUd4t6hzhzV/mWkt6r+9a3ITLSwqUxc+dtYXZv6DnDPnYFvdYiV7If
bHLt4duB7M8B4h7Az0jtRDkH0IgXPX56LW+ihlUhH/hIjHw1EosM6JHFitn0PTVE4LL6sd9LtdrI
EodSa3IQsrdgXQ0kcUoIdTA9CBWNRCzZp0YnuaHNbWj1AARwJCLKOm41FEF1aTzblrAHRRUimmYt
z5+5sro/YXfStleUA2wCtIrh6ux+2+v+Add1Sv104nnmk5ekC+5NLMysmk4a1yO8AJPQYy06MkvR
KKZVoqG3uHzmdXbyvdyMt3FPC1NnSwqIVKBDcgK9dX2wgHpTNiUQrHxXMNilZ3c2NRKRPCXysWy7
L9MerJRfh3EhNsrLOeEA3xPi2l5txpsCA4MzDiXdrYYOPj9tRb2REfi75iCKOr2JHkLBvixfacUo
dZ4lCaf8vqcoC+SkqFknVDReikDWP1Ou0cOX0wSW+zVdzQHgYLRDN0Xn80UUb8pykdumDSUBUfBf
67+ewmbdXZ6e3hF5WJHVq6NPgeZxPM3z3T38nZ6ZLQik+7dDrGM7gJ7x1W6lH992j007s+OqbWma
1VewUA4y1GZGbZGDqzO9olxBt4MBCh6+3AIhfNw1rG7Ok+gyvvnWg2PCcjgTfDZBrnXAmrxdEhRh
3h9lA+QEzurzfLfNmqoTdyJYXPjXAo2DyZ17stcUxILNrXcKB5zVGcWTno0Hu0C12/GfgMtJ609+
okLOpITXt6s9Lpnu3X13NMUsSyZB8m1tgW/FSfVSpekYV9CzTNivkkGbNvYRk+N3fwk0MeXjnO5g
zd3Mj3aqoMl5/S/Q3FePSlfAfLGOiwEoJaY2PI9hWYok0aGF34vMZOem2tz+W5SSJ/SzJqTOHHjB
dJthXVj0gk/cI+k4MfyB4vqTasrly5x4uYHvgCAgGO7RvXbHPAchlgolA8kTkb7taNn19/IEyvJL
0CVblJgyZylxDTcbPptg1n5qXXyxGky4pO6nOyF7en4tjyZzBs5nVd66DtsgNIoUMdgXUMEGDOwg
FCr8l3ElL4jTIx+MDsvecoOcO5R0eqh7/V8deyZ9TzwkiqJeqt0f3pLiyj7Am9GIksEg/w4WanLf
55dvZrjMICleqBdKZnNzb3ZbfaB/QlWpR2cN7a2RtFhfeJiFxtKTGWVvTjCy6fP8+8DQJA7lTHfw
Z+FNDaVWSN5HbzUJO2jVhDGGZG6aCAZ79QVRrvByYxhLya9fzj8lI5iLTBNyQEjr6BnoqzkehFbF
8rcsY1JwTQZ96h6wcCRmxpMgj8BlEEUugKzEqAJ22KIGN+m5lFbVBnkgHjeuJL1+ArVg3wjSKdZH
CJ9mNwBwP19q9G+qNdKyePCDg/H5+C8Y0Y7Q31DYK4qDRNW5KGAfUzyCmauHbAZT8Yu1D8JMRFpz
5dvXhZvAwh2mpwXnQeOOpcUxdoZzC7vcAxI1/iRNv/3AWSwKi+Jx1XOpX89oqZv5CSlQk85R//Ve
YMxHjWDiqsmYzWfOoUcrNAzKlWd0bzmGdn/yaIQyHEfkH3hvq3TWXW3+Bl60Fpe0J/8KAu1dZKOv
vwbCb4NBZygQFVnnm32gIe6TF7oPAZZXp7oMkB+IGj4tfqlAWjSga9cCi5E1NMxHu8NWx52YzSLW
uDnzbWGxJQ+2eoXIQbwo77LTSnYkC5uCKW125F24KHJzpdd7RyeJmh1UANrY0lmK64hJIU1mn9zC
D7llsZGaoQzLN0XmJZrBnZkXeeJty41uaWKsT8aQz5MXgLzrzVdJeDES3xzIS7iXA/ntYsQWgxqw
SBGhtfSCf1TBgrLErSHSk5OzV21EEKyVe3xnMVWXz/Yjux0iHC0x0m6dH8GoggZ1eH1rNtkQ3ZP0
HIE+43b9AYGI/LaMqdfeuQ/W/zS8cibppEG4xSi0uZzMcPf9hbazi0GKU6tYPVM2J5/Pouoc0L8I
wPeaTPVPIi+/KMLR3aFzg5RKnAW0/crWws+mUEVg38u8azeROVKvsrUUw4/IHQNEcGOBtR5pJFa0
F9igCab1DGIj++ErAIsz4Q8DewpV2fv1pemKhrSSYvJBWVipLNptm+b+M9JeIRL3BrWEQvmhJcD3
v6pbnt9S0VLa17DE7CpZfc0EX/O7LCEtd7rYW+1l1lqrJ1ozyb4xgW9yEQDsJUv1zj2qZlks1Fm4
yoOeJikPNoZNYZs0ZkvmOKOOvo0WDk8jA8gTNfDF8ePXlL8bNoazfukec1efx07ry8w0bYSzZcnH
xln/bLmfspvZbnFf6DTEz5MShYdvYYda618VnSa6mLZ04kPzn7477NRkGQqFA6aPxEghAr7FXFwf
QUF5/pT2SEcdzMDl0htQETscegHdDhh3FfiqHF/oD7nu+7qXz9IGiDqQa45VkH17zYGQmnIKifiL
2pL7h/TOlTpMknlGFV2t2JHVcs99UaxNYyFoO5ZKoXyPVdGufa8Jpii/HWHSssddBO4HgMhnE4p3
m4F6XO37azB+NsParm939jNbqSCTTkqGpVS02QcwNbK4xQtLYTi+pUr7vudLvgP/29mIGuFyLhAX
keYgiXxeZ21LufU5BIkQZOULTKj/n+Yanc1CO7KEIR3nIOQPa5RSy/u3V7TbMOE1kFaDSSIRxAm2
nVGbXhSa63FaMsGCQy76b+3qOrn/ajEMwITuaLuwM7iljLz5Vr7PZkAT5kH37KDeWmzk/oVPL4RQ
Rus+TUactNdD8LQ0Su2XyelM4Ljo6AdC6Xzp+wTjXZqtmhmdtR9KpHJxqnXIZUz4rEjBJfgzcNTP
LsgYh+XbbQOUo492HDqk7OhZAZCbi5cKq5Fa6f+Cbvy3LNLrOnx0fRrUMb7ndj/T9VdPhchYK/Q9
UJVZgUbio27p9wOQvIq7OWplDlrSfxnJXDwtqak1LiS8ZbiqqG8HwYsEO/uQMp/A0tupqvgvJnol
UOwhpF0IWNX4jKVn51PS/wivJs5KCsgmrSCxsvs8rKSs0DnnaipxXI7FJh12G19Ob2+QPRxj6u20
Pi7AUOov2m9meANaC42kUyFxtm9BWqstp51ACd+2+Ruq+72Budp2Cb3iFF4dg/wcOljogyq4bBn1
V/RJN672wcZMUnWJxO0Lk1pirR9nN3y7uiFsUd8Q4/Urn9Pow2flLOrDQYpN7dnR2BFv3RWOWy7U
1g/TV96CkzAyiM+DEX2KDiO++ILWCDYFicqG2L5Sn+TmRnjI1TnEs4Erq6fS+/kBwVjwYT3c+xKM
cjTG9e9DL8ReSgbMcu0k+hLyhVvolWt0qqk5MASsVJ1gviOp34oaO3pk+i5rRvkvY4OWxcTvguAv
TzJ+nh74NBKTAwgVmdTGg1yOHW66YuxEdOTY6zXf56j3Lt2mnBcJsXuY4LdF24oCzCllACMghXCR
JrXcrMHffL5EHF6PFP5ZSWSBPZs8vX0sf9+eRvZf9ixnuBx951iduXnY2Jtiz04ySYyVNwQxuB+z
QWlWUf7zlfonIw6MA0m4sAhReFwYESsHwYPU4LHWHsjEOHnxqolFEgNso8a7cw1Hbfji7TLJqwCp
RE5/IbR++gUc1cYAg2og/G/8mj/jm4oleotLblWlDduCHCJj/yMLfRPE/BTiB3Em8qt+Mz2xgCVM
5i14D1u0MkmbDAyqLm7F0YkemJFJYg6kxMyG67r94D7maHrldThqDI1pX0p9B2oGe65qBmhTykUJ
VZwErCDblvk2yCkXwBV3omrKE90wv4sQViq4yYHogPm4rIImN28q4qaloNJ5lfIbDNaW70/oD/s/
vnC4kRSinzneohpIAz+mtDnAkWtBJCAAyV64VNbO67Oa2wuBrX+8vbyFNmv3M3CLC7zzFCp+f1zM
u+AJdCPnjiEWWJDiBX8VWUFIk1oyoQWW+yWlX4q/7ZcuB1GgdwbVEGntBoPJaBMTK/3Yo+j1jSWN
Wny106Qltgj1wPJs08cs1NL9JRWifssFG0Qfz9mIa7hh2t7NKX46y1eQIb8/SmMS3+12terlmyxs
KZxFGLtUF6hk/rOt2AHgHb0M36bF/8nPPj7c3PAxlpYb57s0jc3+mYzzoVy7q2ac834fKWqEKhhQ
1ve9bju1Mo96Lhbc5lFgXqJRqBgIKeY26Gyt2MIYy63znLfG0Rb+awFCERJxkVchiGkjAaAUg8j1
fm6GzGbBnFcDQFFq0hUZ5qjLKI6DI48CqnlkysazvjgV1mayEfGOc8zqaRa0G2UU4vCJF362jaxa
LDS8YwSWm7wxcjmYRNtzmfkd+GxzPWvSYi7ECM5CudkC3FvYl7nJXSdqlC5IRU4BGSF58llLaQPe
tJknOWiNFN4f+6rz9oEQco0pswjxVuTFVFx3dk+Vblbveo5+Vrx6FwgNxhtgy8FQO2holtefdoCT
EoulCJ51f+ekNTH1rmZKJzru3Os5EwL22isDnN4pssvBu+q5uQWTzrL2Wso08PqFXcYDsnpjVtYO
IvNKmicFXf5Ge6VpDuBoiUvci8sYxKfRlg20MplP5B9Tu+sHXxSZgihQBV9FjHCovmgEoX0QE3ac
mbeshdoEznjVlVgFALSIxKIzUVsFDkKViw82LpHtK+RywSmwHtNgEduBn0HvCeWdxa5Yg2+vAG4q
sOjvtV4uB9fyq1KbW2mUrXp0fM2aI0ZWYPoUoXIbl3WCSkVKq1k1wELz4TMuRs9dIhQ8e6IxkHJt
7iHfyoqvOFoR8u32NpLP1AzxoWvz5a0MyEIRJVPfv+rfvP6muANvhWqWN8gmmTHVTP00acECIGb/
97tAppmMiDU0AIVJ9hXaFsqzvNZ0apTcpX1j/NnLYYg3HUAquj05vMVep86jHQ9PAsF8sPGloOrD
puEYIu0uLoIIePJOpHeB3gv11Dy+QRLcWts5JwBhL6/fd9je68Vdqhl6qso2/2emPoCCRhEXsKPV
bkKBSU5dPLTU+vhE8DrPUzvtoJACKa6ugKGbB8FM64efJN9rFT3hQ0Z+GimX8NgUEfpuGXoa7aip
2//2Tv3K6mquYH3OihcvhHdQKV3KgHlv/EtoOjyvNnhuOWyEu+ofrxYsywviabu9dq0IEdunD9As
fNcHCYz3+ZsKAIJEhHF1haRZA0InCGQQED2Ki+fdBom2B6BA/yZgq37FxlSokyX7hkm02jvlp1xL
N0iCjnhJ0wE8MvfdDmaR7lH5j1hfdsK2+2k03/UlfGtU+cvVGxbUAbcDnscu0/ehgDGYFd5cj+Pz
S4HTLwhkwJ5vBW6iRCwWqp5TwBAD2RbHLEjwRqhEUPzPglRnfZaxcBGZDn4AQvfQ7gt38U6+5GO/
/1fXx8BerkDg02+7l/bAO4S20MYECG0Z4h8ew9/IxoixTDfvXuY4TFE2hECJuKglxqFAGnCZ5ppC
ym2nlVtY+Lq9zrvFe8bhIAhdbPunapAx28zFshtOET9xnoP8AKIzcA+9vyoG4wATEy201DmOdMDJ
ll4V5JDWgC+mIm2Eq3hGg2TJlV+lqR2d4V4vaqefMR6CUY10w+8f4uqSruSfr/m/GMrfZUjn1YCr
85scGw8RBTJmD2sXSabUYHbEeeF8Qz2hiQg5QsoUqjwUEJVTQMbC9wtVPd62ZC1vnk3RLqb8Y6ll
vuGJRyyFZVYdaUra/aJ1lsafeKULTyDFuRtfEI89ZRmWPvdAX5GA3ru1UAZj0McZa61T+nHqhpWd
9vlTitjGNQEu9067UxnMSsKzAG2ZHDzElHrem2Rjj1txuUXt4kbiWVLX6Laemc01vIivjBnYpZfT
VmjPucm802KWFNVJeUMUJEdpGmp7uQn5ZexDzao/+qk/8lsRNiLXxRLxWNkr1jPdGZkQd7y3k18G
s4YOrCntaVSBZhbL4WK/Dg8hly1ATwoCJeiDRW+6o6pkeVFg58Xtlf8j7j2wKhz0sZh352Yb2zWU
qhDWj1pewSPNU+DqYd0hH0w7WpSxZ7uFZ5Se79W5ljb4OGzt+mINZRqUK+QS+DwZU9Oicwsfq1zK
ApdD+OtZACigze/Yz0lEFZfv9PUkIJFTQws0r94Am1B0DIxxGqIuscHuMtqf+/S+KnJ1GUyTv+By
nZqf3mswRTLBJp9nUw0KlUWXvEiN8oeK2WXm+5lqkc6QirEWqRBk5usoMRv3yJdVbN706osrXUAQ
iCphWRUeFTZFwKiZeac1DNbd0h1Brr1AJgBta6x2ssz2oU9OWldHdIcQMcbzClS8TGuDItp3tKKp
XVV1PwbQ8MMlIfqUB8yx+OTKofR2NzpFzLpULaezxStW2xHFr47hBWZJYi2nzWlJ8PyDhTRdMV7u
S7XjaKcVwyGOM09pZbHYq7HspqbAxZIr1V4+qNkgDuht7FsgQWk7TqM59JEKT3U4PlmnDt5vHiT/
CNTeK+cJMXAoy6Ej4w68qQJCokw0TSMefbHGvsqZLul42/jEFOjPrx8Ghwwdm1TNGoDp8F19zEAp
ZFbdnheaa2lfA6e4hugAQ+EffuDzyPQ6wMWbtt4U+F5eRGt9tSQTtL5pm/ZmpVc9s8AWc/YqGF0K
b3LyQZTxz9gQsg0SsP6IEag40vQK/jz7e+bACH+eiO2MVMUrVWN4Zg+tP2eo581+HXVMFN+zEEwN
W1ZQfNlHWLQa6YxjYnqZX/r3M4DQeiQ8YkFkLpxXvNQt5dDD5tdu9w0+DklQLi85mTSgCycp6jgw
FVLKmvDWFoVLFngNr7JuAYUVJutkTfagmQ+54IGzP2rfFcih9pZbsUbGMGkCMrEs2DSjx93WWqk4
TSrvO00M1y4cuot83iDRo6wqBYiDc3JLghYCrwv5kx5R0B90CTPRWRlErGMvsi4eLnwiDL23NfDZ
qxbQGhqIqYjArD+S58Tg5chUC/E8IE4Pc/+BO/rFvFCTRCt6WVsb4WrzQSxMpgz6GyFNCihPvi7u
7f+y1V2xU32nEU0u82Swp7aG+jNn/9aHwD8bPw79rF0PonV0dnT4nvMaidgFb5xkp2lKd7HMTjkn
GnfvVbj4+L8nYm5qVxP8v+Z8WWzPY4sbNqJuZyC4b87t7CnnqKCV/e9kkqrSQtYYl0FU35/0lFTK
/uHsj+heE8ylJ+9geYVy6gw2ofv6lz9cf9uiy5q9icgtbefk+r+AgRuFn2NE6IDIAMxAN/QMeIT6
ra+wZ9jTZ0gBi3NM9dzDkd/bSIO2suTlAlCNrBGoHPhyDqKP/gqBx2xzVpYOWpl+orbMMGD1bHPt
fAOMKu5nGaava/1RkEzPZAjYuOnvXrGA1ruYJs717XZ/i67t51GRj1wh5P22yi6HVJEN5ZBqmgj3
/DgbMBgD6pEU8n9DLUcTZA7N0Q1oT3zC0229huMgCvirNN8OZCe0AOaXl+XC39HwV3Dny+vBSm/m
WV61fs595ijakr0xjvXvLL8IgcUuyNE8VqSfrfZJQWdx6hGJJ7saXKZBbIKkA+wGBEXDrzZgC5Mr
/P4X1A41AESXcvtlSkIsReACmSfTEt/PXbB2pdkOd790RibExBUnxQCTsxXyZm0zqDKxYh40PqGr
bbbIaxVrg6VgaAQ8rVT9JOdqV3lJ91SB2DuxX3hFSLorRNplK7Z5tVJmst2GEbqqryKjs5MCcAtd
d7AagFITS1lgNrh5aImC3mjOQmwwMa7VViqNMvgkVfKDQIBU/zTTvMW+EhaO82q3VyI9ks0Rcoq8
/dqsQvcvkHFeR2/RZlhCmfFc7uB9ejXCtDI0Zw3p3mMDOdlslXaiyhv4FOrXIS6fcjP3OIUmqW8N
Aa55CpeCqHQH9G9xoiHGuO+5N6SRzvqquNKcg33g/uCKguouu4KbuWKCL3VH/gGk7G+PX6Hmev/Y
LESBYuOvu7vpUSTJySA2f/WOcgM0+rnm5c87/ezn1Nrvk6Z2N4DxRyNDlhRXKF6rHxt1zboXJ6V4
ZFtFgrs+B2cUaf+FuZvSSaetO2gyd/++RhH9VnxMHLqtx24K6rGZukNDatNLQvBSU1Fo5lXq82EK
tjlNQKDITmtDQqS/plh+vz3QIoo3yF6wldUBvE13nNlcJFtzm/78QpQTibKAunLBj5RzMM5YWIU8
e26RnKdjY3UsxR2DfeuzpzKYvU8LA/OsdWH9vkr3sFzC6VktbjYlW1I9REYZ197lvfStHezAT3q5
U50YlhwWEXrQTf9G1WduQP0QkeP6BHiqs7EnYZgQ9a8y4KiF6Uiea4bD+MketjiEhR+AHZTTpGfu
UF8WVROWY4x4UUjVks4cR3HuNse9gvQa6Eli41WLaebniS3xyhrJ+dth1JsidIHQAeBLVPlLXaG9
ZhFojTwob7u5quToqRDtyQfeDq6usrF2iNXjLc45oTsieXiqK4wH1jZ3EA5HT3AbZdlTojrfW8cD
gWsGrEYIV/yGHKXli/tM3x69MPg+EyVRZxYtAq/Ca2LUeIiz2xsNcNwQTCNiqROQXVyOJ+GcZvoY
vu4Op1pxiYZOVnqAbEQZV+aR7EB5SbXt2lxRW0pNlffLqCS60kqsA7onRyXGKNm6UzaVvxMRYkft
Lmc6YIr2VHLIGIiiKEUa7j1zqWdq3kLNtf+IVwgnLXhPaY55/sE+g/2AyBh1X75JgurBvj69DC3q
EYzAEeZ/xtf6neCWydH3po4On/lg2B0Q+et4dyD+gjgR3tiDO5Ep2UVG4D9J3aepIq6RUErYVMjN
BwOi+j62Q2zxJPKGnaNOXVHdIyyS2Pe6BDnkn/7ut0niZqSuOGFtqUBxAYjN+qqtnsD6qKpqiK/J
pDreXqF3q5Ys9q6ePGNli+MBbNDHb1UcmEso5dWp3yCKde15WyuwpT24ufs4DpQcxGm9a2IpgaBs
fltrtUApYmsBWk1aMIUAF0mU3qi+JUA3zV9NiwTFYHum41jIFM08xwp2cKCUsgJY7s3sGbiUK7Hi
T47oCxxGuTw9QSTvJZrymHbamXnGLrHn/QtzBGiXhbrCcNUJ2wPlVGz80Ma3dwxAmBnPCZ94/efy
ZolKaAa2ZyDbYDVVETTHD9t2D9je2aJY7WsFoWuzX6dunTc5Ry5UIeeOBgxupPgsH+PPa+soh8Us
8FEdnWf+miWasi/wB806DZTfwe3SSi0wTKK2Z3F5G2XD8IjdyCtnJLy1HsPuB/9yyaS1SiacKCp/
PwOtrtNJ6xf0fdQwVgTaY0GV62+WAzolYz2hZJ9Zoh9kmVT1e2Ka/65PNkPmMQolJNqf6cnst3kt
zzC2/HXv6eXltebPqxH0mHs5RAVJtqWvWzTVXD2uVWH8JBDyTIgN+xHTtOUvGb5UsVCWVKruqBkl
tcPwq/kvR2NfFnFW+a1/cFjihcEFQ8L/VhWnAcb48k3lypW+0d0X5hGFURq55xbJeo4OaWKsGp7N
JQAD5EpEy120CLcafuOg5KLj6d9wzu2IvYvmf7oSZvN4zxcTvLrnDzzbqtmDoJNcvxxyBTZyPx8F
+LPk2C5jmVavH073dTahjCB3PSIDxTfiI+Z1ebXxYLDJjwDhcHjTCC5lh2ntm1wmSOS9br69D2fg
29zJZytDO+FvCDp91klju5tnjuOK30oMIT1Hfn7rHnw8V2rPiLdz/jmTNQaBPVGJSlzcrhxEW/o5
ur+OJVtTVkhIuyrCCwwS6vyaCnkLYIN/FdIp1EZXoWVW2poSYXL2WlV21ERttlEHqybOCmfT7y5K
qHDcSaudjqtQ6xuU8fiQWxP095RPWI2Qfhq7ED9ImhV+b0xuC8JKvClQuccx1OsrGXBw/E0x6wqb
N7Ypl1nB/vfQa9BKLhEZeIBpfZev4DGVN3/KdejH58gSqhopSEoQ9/Wc6OYf8FKfjpxfBgxB6mRl
vuL+qKpCQJSnosxhGMdate4GiHZF0EpLchNUWCrtJqAr2xa5jqdz0z3IjoXRFwBOHdeoCMW3S/VB
4TbnkmOKJZAcVHx0osMn5LZzrNJLaXvTl2oa03dLOANoHoxyLJghikRrJsb6omtTqV03IHPD2srp
LIH4U3fPhYdvsLuSxjf1LOCYAfhgwQJbYwDjqvNtgIrkaGC1YlQKpooPYylmMp+GZ3TwOfeUdvgU
5Q/I5cLXtq1fsZQBXLkVSYXbCZEA1Kg3071OA08Kg/ZDDr0IW7d3MIBth7YezCPWyHSmNjpNP+2T
rREPS4kCqVTPXXcsHZSYG/v7UUd2F75XVjpHWBCKZGXWY2r6TgesDDakm+JjBe75twtBKOEa4EkC
IgS/Lf/RUhO2/4SGq7c8cIkNH6UibaNTt8lXRlOnixsvv4B6O7ps9zoIyC2z8NEkfY9uCc9Fck9r
n3HZlb9lhh5fjCMFchTueA7F7avg3nVeepVS4w9Kq8bPYm81KmolSePTBTfrkj953EjR6grCEPO6
03ZNYKEYaVQ38LFpjfCSDfOwggCuiX2wJ9aLv7BAre2TR5sXAT4oYjNnIm80IW9Qo+ZsjGW1HkNH
miZ8NBiCI8nxcmTt1Ue2De4gAuyyEq9Leq9fnFaIGMJMA7ssDYuWo9FMP2B0kWEyV7xvKyAStwh2
A9vaRCBPy5U9+rXZdGOPB+1TfYaSeQ++iIxRn3BERYXh7cymRH4PNV7y/WfBUVlCeFGBSt+riTFL
Ae1101vGuX1y0QONjbMrP1u452HUTPaNK/u6zdHEaIefWVPUVwuRL5zI1wK/e4xywS/dkeT0L2dc
TsiHvLoE/YXSP284KTJ6psxRY4E56saUsAg06szZrFXGBAWiALtB4iw8TqUq50TyrYsY8jovTVjv
GvpRiglJ4sTbZ/I9cOGh/bYCi6vdOc39P3orHIZqnycbrPzrBWZYVewCYRJXBcu5xHqZ4woiYd/5
W8eLx8ooVJtisKX7Kr56R/oywOtWUaMkkVtKnvWFRBZM3R+M13v6W/9c7Ne9IFJr1/JpDSShfDct
701h4HPubTh3qxWIyTZQ9wbU2Pdj6F8p1gf53kIsbqc08M4YejpYBkjQYB86vwmDUbDLBjBf0afY
Aeu1t5yKzw40KuglQ+i4DmYFJd20jRyHva6edQym+ss0HnZ4sSZEdttVvEVOwBj5MOhW6n8GyhjE
vLHLqHsY95ZprdtLzZojzcD1vh82mlzIyFeUDwk3CWLG+IXm5VpOsNM6DYH1P9RerPUWJMx+/lXR
izGMxemF9/jtLpppLv6eVap8qzpFRvDPlPg2ssyF5HosqZepF/LxnBFt2v1GcBjM5KTmuC3i6C1Y
Qc6C6ykjulPMohIJd+cFFcLA0WufeQZtUtqU0Iff/EzFNZAOl50AZ8wnONF7sAYSQ32gQMpGcLwo
oVFEcoe5eXU//Eiznz1nx5+yxG2OGJCUO+IUKtB87m+Q0reJqUWRVAwLKilvYRkg+GSrfTcWI8Px
2sK4/rPr3huScqcReL5sjbErqJDCbDqH+JyZ40T0h3RP8wqTmHwlJ8S9XVyfX/Tth59KuA8p61K3
n32n3EZypTwbQs6lVMwJcqtrki3qXoLLfTQbspVUU7UiR6tfB4c6HE+d6XcdxcE8tSPkIJSp55KW
rNgExxcGfXfaxUioo9O7wc3kFPRwxChWzK8ndLpCaBd6eSKnxOgzbeMF09OTlEVcjLItBN7S7qmH
JsaB7VMbTxXE2KHCzeYb6eIwCODiueYeAcGePkTz+BrOKFbn3bBZSPQjaNkbR2E9UXbuIRW1UXDQ
xa9JJxtOwQ0TpMlIVeoqMyfSZC8BbqAUEMyxofNUJlGqL9A4IJ6fAB2BiV3vv4jX2iI88S53ph3b
esnTubvYE2rfH6Qhb0V2pnjS5yUIMVYyUUwSf4fwXNesF8jt1tQarBQ01cBKHBLYSlK1YfqL4XKH
wFonQdlwIeqkp7v+sRiPIPIA89HXJtthn/sb3csz4zUkSoxscObGtsaqk0QnrjNNPvfE5CIBvZuf
yGfPN5zbhlLcGlW2xO71eNDwf/mFDnMzLnZPFtlgVbhTAwR+D1rjmizSvp24/xll9Bf0QJBRzUDH
Svr5HGchOhyVUYfftUWJ+DQXM/RwymtWuBn1L9TNifJhOxboZ4K3f40Ut4eUs82uttDDxtek34ca
Q9ItrPxMOnt1W3oqamhBFTx+ce9i7ZYh5rcBmGFQuIdcygpMtBIk4VgqTfv7wfeUMGihgfDfVZsF
8ImojDVRw4OK8MWd4pyRGdD3COMjbNh4ouN96wwZumvnJgTvj+oJmOSzDNAnwya66EUtqD1/bqij
n4gO3nvN30YVsqPMF/ZyR7V0LdL0DYg+UZ3w2Umv1XXyn13xDKiDdWugs/H5Sd2TDeivDuC5ATa8
kjC111Bdn7Dwsg6bLjoIYaPOiGFOt8wgXNm3Ge+WUbfpFP19zgQfM80fDJFzK1tl69QAyvdQdDUw
zexdp33On5BEPzSHLy07/0gfO8tQ+EocS4XjrvDYFqWrikbWkKw8N5tFjD4skTAoAp926xPKWmzF
S71uU+i3futUokiwGg+5SsiGMbwTByra4jjcysENNgGH8oyvNpwmOJ6uEaV0cfx3+MxapVUn9vrg
Wc49MxxyNC/xwuWz5sguLq8RkWQX6EYTwOM/ad7ZjI+Lnq3BQ+GtftukOF+KYdirfGRGX+VSGxoB
CjOS8Jkvn+rCDbB0jPA8OEesFY8vWfWFtOdZLyU+M4fPlH1xbUFcaSbnHaLVCHQFgjo5w1I/eRkn
tgw9kDTAbaSnvlRPaAGHEa7y6X3oO36GwcoORQz706KxSQTyfpAchStc5G0cbJXf3sVRruDlTsbn
kXSJNjJWCniycYzvSD5chDNzqs8t1/iEMuzfFt6c9pHLgcYaqlbyi9BGzRODv66Zpw6ddSzFtiMN
KDmB8CI70Kj1wjUZNlCroG9Wd4Wf5EwpjY64LmkmPjnSy10AbHBP2y10YJgIQfkUOr1oxDE5kpG+
QTilVY8qI2EM3FRQ+FigRMtRN8mnCeIZiYErC9ueuSakwv6T1Cly06S2fFmSx+XSwR7CEI117Tin
Ce8NUF0BONiL/EWHI9EQ7Fj2Iidwk6EXE/wsyxJv61zrojWVTTh+frgkiFRu/ojArEAOLLfGAS/p
+hl3PMADTUwfMT2ly1byyxYI+pSKXz/oKlgbEEHt1Yh8uQpz82bjmzQN1FS1M8MKf9Bm4NrC9hi5
T1tOFAi0iIsyRWk6LRVl6tBDyBoPVKm1SH+VYxgbqXwjzK6XQAY9iqQNOHV1YEUqJWlQ/gpIfEIC
XiOmjR1A1Vaf1Tc4k4ItXsHwZdL6dU7FixDOUPAFNxNtIoF9cPqR/iqY4BdaUMAbxqDp+AImusPe
zvClpxlQ5PeuD1Myc7xm1m1moeupCjVdW+CEEXS/aQrLQc5s8uVx+YSsI/5DrMOc1zPUiYlxuJPm
jyXviM0pnuxmUoQ0qyUzrtNOdGAFYdiU/NL39GqmNtYo4bBMvaUrQIyMuYhXAFGocGyA/oCetO4s
EHf/BnAhiKBLVjuMvqOQgu8r50/Q5jXDhYiMIfKAHbwUXuwsi5N2ITVz0sgIcGSkbjwxzGNjG/Tw
TkikNavUGkP2gqKl2RY2sf+gqDpKPS3FZshTN4W8dKcmJdCyZ9D914Xf/5gdImK7B9tWx57LBHTg
4NFa1VzW5JS4BOGkcivYKv1fjkuo1nVdFli0Bmsqb4HNxezxPS2KNKp92XgdUsNqTyGTQF+GDgwB
uaueAXSw81fG0Od3fT4CqnCqKbUvvJwtYwao63q0SvEpmqaRkFi7pE4sfMwIBqXIU7QOe6PZuY1H
jJ1smQh1jzIbuzmDHVbFZiNnxx7hrgnkq2dDTcIE+OtgksKmeQE35oIFXE8gqmILhcc0RbO/hRNK
pZP1NZ+7P3jAPUnMerQv9u24lUsJjYPHxo0Fb5K42sdBJgGc5vqYuM0gkd19zr50ygFF9TmBqgoT
QFVHEtEJDxLVBXXsFK27pkFhDKcs68aiL+SfS02mp20FTZf1MCBp7v45cbnbcce5A8MG3ea4DBGm
3wx9q86YM9uNEi4/PFbfRe0dp3pJvxZAuBk+Nfu0EeXueXsjUgWWYoqYBfrMpPN9b5uJzJbJmuaR
Tisp7KkUxDfgWrs2ZeW/PVr4VsDyFO4lNgWyFdD/A3X3hVQzrOutLBW49YpahHkCCxk5UwJfX2lJ
JM7V1tfDaFOIGCl3XfiF6lci4zBE90DRnHeGVovF8RTT7DNwVrfc41ILUhblfgRvDGn0vAj8m2qZ
EFX0aF9x9Q9aA7VV8/qDODu4M+ae6RPLYtFtSMtUil4pi5oZCpp88xtB1O6d95ugkLc5fJCfxouZ
8Yqhy9waMiK2NVmetzYWTG93imPMKnaP0KtkRKJkhTOz5ZJyrxvlFOZO2mb9QJEh6AIvv5mW1dwd
0W7oKR+vGzhJ+J6f9rioaRjB0diUBgvVVzx6e0ay4lFd4oSfI4BYytOk0emR6KdclcpGSUTFzGQ8
o07MjF13pjO2Lf6k/iYA/w2bBWz6uQmBYcyuQ8UctbYDRWF04f8mK6gxJ6nbH3LNFLslz9EjyTDa
ms/9+WbPKYQt3tjVe3H8cdgdFtAB+wr0HoL4jxKbDap4zBw0BvdMhwImQGqrNEwWQd6bLm4roMcs
bP7n+6RZtK7XyhnYQNzqSrGbGfo1WST4SyZryY+mt1QjgGKVpNbxNowxEFxiEUda6uHhrhIJg5cJ
JFTVVWHiNE5O6Gun8Vw4BHhR21kuSAQ/ugjIqPPhWIHo518aNEHXTiRg5ZsZNfn8xIeEWJqCx7Lb
YayS48gWrqxyZF/h1M1qmc95z769qyH6e2PWZCq6/WpG8FAV2dpkWKn5RlpsuN9tUlyZReVjBWzI
PBpV/+p/oOzxbKMIEmvAOyDRqwpo3DOW3z9ljhnU+kQmUxgZDsz0II5ZLbED56wvMJpc0L1mpXmi
86OILwGlm232xEhhRppe2kwVcc+brURHAtcVctkv0zrKarA8pWNrQF9B/ZH41nCCHHq7t3jVtXfV
pgf4TP939NQzyFouAPGpDDRO1o13EqLr9XVRyApOi5vKWEiIcVrNOaHBJqUbJWFWdniUmABt1mZT
yjFfcQzpvd5yt9JVuWkfC3whnQg3umKNEXaGRsimziMglIhrqIyYp4JA5HN453aO5SHxuga56zQm
meQMCJlcbErii21Z8eYl+mc9R3KhUXtr9BnhWjGxhp60Jnjwi8rHjZBuM75fpQAScqLdQb9oq8wu
6/efOkd6x3/6Ua4+vfktxDsn1DBsFgpwdCosPJFOt4M5ojs1FdoaHhFkXUaYgeW3hXvZ9/URUxEI
mBO0lnzDP1BxbvEEXzzey7n32/Lw1gA6vxRJ1MQhuZY2wPreyJVfOlET3YPjeYqK740T0EroOswO
MvhxKNRtR5rphaMoBdRNCs37K8f2yUDs7mN06wiB0BxZHgf7d+JQsiN9qtFNVBtTO/uSa+QDbrTL
JmJL8hFiRYDWFGJeX6n8LuxrX9iSBLbIVzJLekPW4OTGo5Ik364DRcTNGv45QmZ+H9uoZigS5OHl
QBye2EVnA51cHeDdOIF1jzNyBQQffQpkvBYG3LgDJ++CzHBqIV8q198TKm8XpbqLS3UPUf4tVcKE
UnTK15jhJmaM8mqgtwOwc46bQW6V28kRaCXxR1798Gdzn134YDtdB4H/B+bdjyEp4PXnu6PjvReh
uZmO3z7XxyefqERq4L4triVaki/kuOsOVYeGhJBxHvztOGwy4D5sU8gv4A5n9YODDQhoi1p/6cUM
wf1m/V+L2eEWQzMiN91nzyqo1OXtm9k+v+IuBSAa2i41Q+KjC3FKdx7D2TRV0zpvKTWQrlEwzZYI
65Juq64BXNOegt4o1dWpaBiCIVPkHq4JByLKc6rPHmaQiO3I+SF+jpgcdUamkh/kJiPBT6yoI2UC
ThZyxed6VtFZN3RMwGGbC6y+XGWFp0aG8YcZn/Slp7Ov20hZ9wsrOF4B8X1XZ/L39pbp5pNykG+u
gc8ILabFE6HjnjM8rrk4k3nQjMXBqY9GJc0L1Abo5YzCGP5iG7WjqxMb/JeR3y5U8x799DHYsiYH
tBdcMSki4HhdpK42U6uOkyPVN2+6hBO2BlSPHN6sXxLiIXqqg9u6ZF+FvMZfEfi+7mzjn+2IAOr8
bBdRk7UGC4OJMx7aYfdkE5utWRcHlv4IPGx3rpPe4Ehk/D+7Tj6YXXTZOIkGr8XbaxQ30AO3c9KO
0Ic/h3pHDzhiK4whqsgeLN1JbCYP/qnvCDBeKpEcjJRjRx/vg9GQQEGPp2nuaFl6mC483eF4WCGV
aXj69WjWqnqD8B4TFFJ+UkFXuLD68pK84tD4QzE36jUgX74mbkdRp7joi6dCHTMuolqzdQ7hdVY0
BGmPtxpkDmqfOtQfSzd3avSJ8g72fizXweWrnczusxVcNN0Q0yQs+QfpJbGYmGYlSUd4RBWtas0H
tWQYKsWDgHQMCA0uFQld4jLmOdriQ/N5IGOB7bKgMxcHrA9hWcmWH6G8HjESvztOp4QPha0VUlgo
byVF2F/xLuvrxxYPj66goykCPlpjR07VfnLj/9nW8nk2ELFJuTN4d6tl5pe7jGQlmZEjtGSiq9qf
bzCJRjjNLasdfHPuLoNcZYvrXpjzWGCaUMQDl13lsrCSClLc4WrwYH0FK0Nx3lq1jLwpMLT5ns3V
g+vltQy03euscIsilKZbJlWrShYWrjU5nckusyEkYBkRDSRhSAANVV+9cgQj0Ae0tqOIq/wkqrqN
p/AeG74QjQi8D7jftvJWH3/ksBKfC6y+cvd6dp6yTr9CL2EuzBAlNJIkYQD04k1cHxiswrf1xaHH
1x+cfiYCLIHlzO3eMKXLKHBYKjdhULk+4NaNGo29Nsocq0OXIiRpUYpUn6iqD0r/wS6DznhZVRud
poDUVnh93gldHn9zijq8l7ieeRxseRXJEkSCIs7wf/E+x2h7wD2DKc00J4XZljdF+I83zKUqV09x
knqhDHSHqPN0jHUy1vp3bF/HHE+iJ0pVVnoZEmrCX7BfhfoGXnEHiJOi3DHnqaLSRK6Wjt3eCp0x
Dst6P+cuuOx022Jn4kg/3kLzrLhHNdVec2naqP2avGLMk6V7AomWchW9BSxmnYxUb+JVFxxb1VCz
Ik+RgGW73/s0/GtZ8CMxetlBSUw+b/5DW/DyWA2ytO6ioP5roZvqQ+M5nE6T+4ck/BkrwmiAot1A
5J2Ea0cmfnchC2+4hteYXS6lE5oYYKMigKvbZSwcQBsCyHZ+4hxvG3xpAgf7jOhQ9u2DTYRk1X04
2T0BVmTkib/Sef5frAnAiNkoZ4y0Km/0ojw/nqlAZ0g1XZYUG4IBD/QgpJWj1Bk5RofL+RVjDBLp
zWWLDETOahV57I+XU0ewGN8k8bW9ab4hwjTGXWZkVem1FZZpPIwp9pnr4bBn1VgH5s+wdU3Te4/8
S0vdi4UnEYC9LspMONRQK5nyPdsr310h5qN0Z3DV4dUUhGuGA3LXUKIEQDdqEp96VOiK32iksDde
+3NxsdJ7IZzsNK/ktjwdvS6iG7+BVPeIB6EgklcSvc49sXawKdTE8pFK6Wo1S2uy4IJGsYgof3Yk
pNDETzxEvY1A/GlwVX77bDSXIGkjxprlh5XQWrUc3DAL8Eom8ImjTbjcOCs0Hh36UfDCPZ10tacw
S00IOesRdNpY6GajdXdb+l3X+L4oq9Y7YADnJBhUw7No7XnrP65FqVMAV1tvxSK/VKspAinCAbHV
2midwsYDHtuEVWKMth0cslQFg3p0a12uUT5kVRB8np7wBXNNFbMunpJWE+CAKzw6NMm1bo1Xj6sF
9pEzxT4htr8+2uRAoAfngRnobFbcu54+Gj5+9jHyTYP3ANCv6P2V6EyM2ZU7rx1NDVxHWrbS7/Qg
wCjm+h/bVnf7xWl1uXARyjIF19TWS4inqwb/EfndcxkweVSr9fgsHY1WK7IpBcULKcEELO5JmBBC
BhcvmGdTloyvB8O8ddUlEMehi+gEZBdFF95ZkD/NsBbZsNEvNfs36VB8BbbGqjfN0q04enA58c1I
CysxtlBg24ZpnIhAWBMKvG3zG7VnuP00VK/8LTbnZX3EjsIv/RDjuj1ldVPNh3mrev+T8W0PiCNa
G6sdT8hGojwhxdcJYtpPnjd2MMXdstio8GUMP8ZtDtHmd2ezdir102vPZzOgiN1s9Xy/FukoZGo6
kuw/14/Hiv1ukq//L+XUg1QswPb4lGrO6WB+r4kpsltW1MKOInPWx4rOaXL95sf+rTdN+XnvRGXf
u4lqpmb2wkcFHPf+Dp7j+GZnNVyaWeemDGx5yUUTPN/6AykWZScRqJ0yMWwb3ls1Lac+Irw+cft3
xINn0Ua8KPF/PPrHc/Pmyo0jrGfqbnmq/ZN0pKKK0/VK18Y/TPmEPdzH4DCAJnYvilDqrSrJwA9H
V2dsLleYgsOFrXVRYCDpGPpjqQ6Misa7bQ9+hG/HDuprA7e6xrB8R8+/9tVam4LTc507SYVjB8F9
iOsmPA6Uedh7OuzEko3hc75a1ZF0+5wOLG+NDXrF7SNfFBKztzG7DozA512KSKyV8t5T01CgE8VT
rFuDRFQLY7VBfMrvSP37/dqk1pIXwYztUFpd4FOYdnseMlLtRAjjJYgN1GX1zXTMWUAUnOgr5uT+
vFFMzlAH/D94B5k7NoqE8zOWdMiQ7SS2OpdqlrJ8CslRN7maXBCRtRRccmGBmVcHsnWbGTLy3y8b
lnkFtf6S6GKd3t0t7u9GdqWvJoUMEgkKNc5/EnaImsSkaREI31Pb3GW9AspIHd+ArAdtp4O/Yr3F
7i3ec7O0o1KwGGqhXj5tNWaAx96UkqXtS/Y598KHI8Ry5pu7WJnjf/yq6fmxYcYCoHwqgx9Mp8bT
ixiE9yOI2QB/pgzKudSMGo9UPfoBV48otYmxQ3EiXWZelKZhL/SUgx88/Jn3dYWHOO54OwXe7qh0
nAmZgbMHRz9NU+oA698DKc/U5b1C4a1MqWJmRS0U2gQGLkP7w0AFjQ+KKJ2G8soL+Rchj7FhB8J+
ys4kLrNtbsT+RR9fcUOvx77KunkvAKrva97kt1LlgzjhdBStFHRph1vuhUp5c/veTFWyOwiz9YL5
1H2iVyzHIBJim13Vos9xzFI5zaEtGGQem49MBSeaXe0XuVq25Euuo0F11GKhWaezE4VEqcfvFqXb
j0/mwnrKJE2XhtWqr1cuF2PuxFyaseavKNTrmaiuSqqUWjbcFGHUmUnfuf4yh3S+U/Y43DI7X87U
+AQtbTXBtOpS2pqa4lcO3fNqFt8r6G0EMc8Zb2gBs7ZJT4cDFFNI268Za3Ab1OQKEtb2Mjjli2IH
hpxF04LeJ/7ACYpC9CUXPl1LZ1OmceG9gvsnHYTgSNrf9aAwxQeo9en7HZfblygV74rI4U/eYEq9
PQX4DEz6vnez8RVZsL5c/4Rocpajh+5zx6QfE2lZT66e/sM5XKH0j7PJ+G07KJbdWssZfArvfHOu
t21moIq4I5h/Er/s4h+BVS2WLizb0N0NZJamqJkIT9HdrSCukurA0Eia9hw9v2GCIOr5e9n3TISB
b8GheXjBMmgVvZWwH7n8JaPt4r2vQmVyvpm5DNYF9n/3HMHqbJ0kck0Cu66UwYcY6G5T4CnRolgV
2uAJ1w58Z0Lz40G1ofDkEX8ECafFsN+4RAayBDCj/zVH8Qm+kGIiR2yhVmAeL5Pkp4KvsTnLfJtN
YQjm4jfbR1Zo2Fq0YtlGGX3KsWuOXZqvDlqQX2sV26xyCGyXKfxBpcQgQmFIdMKSoqQNUK+DmK8I
PlySXHqoMBXS/nFjbD1kVISD2wd2sodbLCJ5b3zE2baDs+/qtDzmQqmcOWWIU+TYRRONsRqbBd2l
yDdalYQQDEGbO4Lzq/huBp57PykcN36+QWVf/SQBsaBYYISNfWb0lW/Ivva/ZeOsxpg3ryvRs2zQ
J/90MY4mHX5oZxVi1yJlDIRO8xnp6PAH5ukp6+ZbbHICQfB1gyrYykHqykgpSAVMK2Gwe+AKvrG2
DCEPJazLhQqI8dlCcEFGMRFKQNFDaKlqQc1X00SFbp+vvHv0pUUfJn5SfLVqVNaTScH5M7fPm3X9
fY2hxucBav2UJwOXiOX5KlGTMFOJ3+sBArFMMAH9uh9vBwGlgPZwWXq2QwA+dmLBR/ARZKWk6L2c
8l22Lf1/4+c16wIDMFZNtPO5E/ZikKfa/Jo9nP4KH3fQegwjCoUmCdpIEi4YW/uNTuiIWlO4aBNR
K7xoy4EjQiAmI6b8ZnAmGtK+J/0P+372JFmeCPqJvFLporjBJsaNDn9s6umPIzFi4vrkovQ4gGnf
DkKmIMaNMyb0qgb+Q2/NkHjyDcJ2wAHoAeGL3tBD6B9UYpwjQLsl27/+ez4o1CdHFpZ+Ls/dZa+C
UqFQ6fgcDp+jDQEJK/960UF99H6oqCj8qBsj1zdyPqxHUz3aOhSZNd8YXxP4suzbgFkwsHmlDUwH
66ALeu4MXzvuYGO5pIEtai5l08lLDLcReISII8pCEaSWGeczC3/36+NIk4UzgbysYYrYBN/CdIhe
qDQ74Z1bah/c/Pdw7yn82MlB1LMJCi9NkIfUIXm9uWq5GadK6n50k8/mocEUchR+pJ/O+2XXr/hT
VfKpOxVpL6n5kDWujVOLEqfypHAgnw4xObmqPrl2Zb+FGEtkF8eA/iyPU0GnaUJvHD5uqTNY2GF2
PU7gruMAhzU+6oYeeWP3yAi+KEjMRCtFiUg/F0jgg31oY5nLJURIQl8WHev8W8OzF6+4abX3oVTt
54gTw+mbeMHWoWxe0UHtoV83Bv9QWFzRYikaBWBAmiWzOUgSvME0E9YMu7QBFjiqx2FWWVHrhSp0
GEtTJ/+N/Zmu93awxIij2Qsjwwi7s/F8H5KpB7K/iaWaqV48fzYlw4U17hYOwSmo8y3wX86EmWP2
DUEjLCx+TN1D3eY58CIejAdljl/Zc6keX84PLjKR0aY2IjXWjkIeOnNBL6qyXzFUOwTYSk/qLhnd
oJqhpbrbxcZ92LRCxhpNZFKwAv+WmOAi1hwn1ETceJXpsNi5Qvm97Zco22z457p7nACkf/K1B7/+
VT2hDsIs0LJeIjd1sfdbPzMvjfK3CeyULYICpcZ0cHKcUruVhsUqBPn68SwISqbwBivI7GyM4yk+
aCnghuk7+blMk9KESkE76tTZEuDO/o1C4DTaaSOwvgxJYxpGjERr4Dsqajyl4XRhui7HNZ10oP9a
lsLxnbaJcsSDppNcURE/pbi3cJVnT8e0scdcxf84/KuTZFI6XXR/OZl/W70E3QcJDTQMuA6IH28G
CQA1P3U7lgwPPzgZh+E1Xl2yqxhTRutPCWD2nOhB7QbXlYaADAdIR+X/geiAPe+B53CbeHeO06/j
rz0bT1rcAOjvQvgFkLtnZDuy//gfWX3BDOm8v5wQPlXO/tJ52MQms3JIeomrPFM7pEv33HbeHjmZ
alJm7VfVeGL/iHI50bK5UHfw3BHar8pM66vj2yycSgMh5jH0P8Li/DiSebL70zkNsfeoYlKLjYz2
ibDudFU9QkL7LqG7OR3CItB3nSe2htbECOQuRLfCrC54dR6MLJv0SqMNkEC+MN1gvm0yXeJiSRED
tDltqq2iPDBfyn0t23rTUzj68/nTJOY7qRjG/zpvLX8JRs0tooszLbOGWuN3w3QUWe2o79N9441d
Bav+gguR9Nvcj7oMvoRLkkCzJHay15TKiA96vm9z3n8cEvpZOogOafuGNEYvgitKRmcfs3YRLmki
BSw4f3rQdatnA+HFpPNJQdiQwRG8p1L1ODnG0O4c1EViQFvNGbkG6HAT1IGMDddJ5Tsh5eM8jZDM
DetLcwwwX80rbxQ50JaIfW8YlM3pVD6oOdnv117p0WxKHknir4IHWJ06aQh6yj81ElDgzBo/VvHl
rRbXAoit7nPsNPZGMJ40sLJot/aoFu1JL9V9YxkNQRhJeDhiX3/JeHnDe+yC2n9DFmZe3VLBqUMI
k1/zGcCSfvwP1NYLRpAQZMMAwujO8tfySsZ7Ex4WnId7EaP27oD7t9qRymrTYPTP2rVUUGSPc/Lw
uMhSJ2lMlNi5Np2K0P8cAIBPrzrRwaRiECvRYo9fD9jIpn/ghBgdRUZ/QdAhrU5vCnrEHvAtjJpT
LDvAY4LENqfPQMKOzH0WZGcYDmh9nH7kELyErstld4QdCd/koN72JelT1AfY7BimDIXkL+3QBWco
yqbkjYmcj6zkKyqPoGs6IBTBPmHelxxqhZVMs0j3EX8czDiovyApK1UFWAyzOHV2FOoeccDT9mxH
4+x1KUf8cIALJabSm/n6uIKT4tzUDx7QGCeFz22Yyle4uz1EHPr8MZRxEX/tRXD6HPIe5LbPliXT
hsrdNmG4QO+NgUAWEHU4t/vRKOCDgr1jp0dVtsB4+InBzQ7hhRoxtFnuH32PVySz0+9aqsOsPe6c
M6ke0kBV6zUrkup+tA1KgQmoQWRWIVdi1My3xBnovexP5iELJlBQcTKOs4Tlr20vUEu/mruBHTSW
BDMR/ELAuggdKZUALMJXZzkilZD6LPVL+69L6Lih60ijnHMJDediX40S9WpeZCKNFCW47wlVefGR
XlF4igUOw3uxflBzjdRu/cxUJNPWzaZ63PxevtXGddl5WhrotIFlEQ31x4ELCP0p/V+75aZitQU6
pKVGkM4TvlwoJtk2e8A7nlJAVg0ebm1/vGoO2/+k44KfmBvs94O2fR5HJb5r7bTF2tto3ameh2vl
D+2DcazLzHJgr/IP5amBSSr3elSEiEem/wHw5oMO40sXMjtrPjiGyx9fwKtNZuDMjxJgdPqoWItI
9a6jrdSVKbdZr2MbzMra8ORMXJ6w46C85nEPgF7Qe9W7WH5pnbrgpfiIu3d7JdZ6CkS59ZRLHgzq
kQI3SO5v40QwaQaFDcQDZTXLUS7kp3+119+MPrsT7G5soK5Q//HVBLShl4NEAlY9mJrufgJ/P4Mu
9l2JSASfQiO/nOtyKaSoiioR2VL9Of5sPU1daj4rta7B2WYmYJy+Y6u4y0IbyHw45J0WRGkTQ5Eo
14pqn0khCZuitXx6JCB+0v4E2oFAv4d66e0mVbULX/mtCokr8wW97o9laHEWIgzNkCiNKxSTNm7S
UhniVCvTckBm2rwrAhmrOhot71kDrRWQWtcolDB6YEf1R8NenKqi7ALlMHH0lI1mm51mTqUUH0hk
oKrvnVRW5YfRYai5HWz+zHdTy5H2RzLe9TrPnjAcNuj59RwiC1nOmIpGvwgrjNTbc6bllUxRteF2
47ryTuxzsltm/WD7K1nSpmpeOG/HCsx9r/mcApUkprA3vx5HGLz47lHPElMKsGK6EP6SkAVEg6sc
j+ed9qswhbrQ+/eR/4BRf65vU6+sBzyG5TYQiwO0f36lkG5HuhMFbMzmJVt8qKB/sVbt4OBjS/qr
coa5iOfxnGdbU2Qs/xmV26ug6uXEPM9J0SG9AYwQ/mEzLfwQ0q378hU7MbzbEJKeb6Z8XtaCo5QU
dWcX5dySa/8qvl80bpWMZqv4ezpV00P/D7HXMCS9LHjesUy6aII1C/9j+Ok9s4YST/2/9s5MHnZY
tQr/vjp9V9XYoOuLnNywOmFjVwsfzynZwo4YgCez29yLNe/8BuHpMYIylViOyczUnbjZ86yMOEnd
iuVaUrbziGKu3b0DceJJULOyQoNIinbZr6tRtLceNu0Cj6n+YLrU2MerOVOnel1tP7rCqtpXf3+4
SvCtU7B6X0fpwrJqxTwuDZcjfQxtUmsi63y4WcXMi8nTGoM67vR4JCuSthW8qgXU2S0rzB2stjwh
CfgR4knC0KhbtN7ATXwq3MI6N////5Wbnh5ZJlPG5qomxI12cT9rkfEhkfDKrQf4Ie69xja4zF+o
W6deqaZaTuZn/ZElxdrf5GSFFgWJShC0jJuiqzLoi4UH+mtRDY2R1dRk/KJeShK/F/Cqhe19uTmJ
Nn1dig0v6SUW3c/KjP3eJX/QxTxWW/ETyzqxqITf99VbyMgsLMTfxPjVewMASk8DttwysvPgXWuN
6T1pbj2x3Ci0w3JRjZNkHclR63/2CNqFiT23u4pTxMNvb1V9MaMCiqMDzLcieAmWy7rvVsSGXaxr
1GOes3AOMJB8xB6kG3uglPbfFjgCn6D6uLwUbESNPhqobtcvMYpspm3j/8+WzSGRbg7DG63UnUCR
SaJqD8UGwQiEpzWHDE5ugwpzwAcHmAx+oGpGtcZrjjRc5kHDF74wSApgiD81CxDzEQgkgKbkHN2T
T0c0Tiaj0B5tYlIMKtlET4/02UB9HnvKGghOOew88XOuEwiqIaY4XKteyKM3lOy2DRW1Ri74hYz6
4FOxEHz6IebGQrghGn8UAjR3SQgBMEAXZI+EzcI6YQzQI1DCV1aK11fXLVnMKNBFP1K5ecRMJ8g9
uqOAfxfHDP7g3HumE0weal0HDX/Vq/lDFboRPM0bIpSXb7vdInPc1Z4Go8uPBJftf89MUN78jXJh
ZRZ39ptfeVCO4zqA8b8C3KkRwsFjLmZSgCU6XL7MYZBw4xy3C0ZZ/e0JKBvNMpR9fTw1z0a4EmTa
/CJy+nZ+OD6TmoUkd67mNX65NNeuiyT1jshBbql4rnVJR4JF51M0OUisjmQCloRruKQeBMc5QEys
zudzBaBpxVfjiPr7j9A8ro0+lw343vFYvlM1QtQFKxgqtAjAZe6PH+o2Ls0b6mIqWybzBxh68Xw8
YTpGTDEtCfhyYe9JYMjypMkOFpRE/iL/nzl/su280gSUA3HxgVjMBzX/d5HaEVj5K8jOaeRbL8RR
DjjOrggiOKxLREoJsPK6F0xQZqSvwwMCres8j3y0UP38tstPiHbGD2L208QUhYliO4Zu55L0/gBV
wCSNnUWVx1bLkOqjd38ZesNq3zD7G3hEaGvBQN025jGOemQ0f9+oTmWRzcbKrrkyny1JDN4HQwZb
BcjJhayY6oXI0yErj0NrxiQuS/Bdmq79HkpkEgOF3M+bdGzsoL/pD/Oba6PpFQVkduyi/DHdF4Iy
vBc6IOxXnonFVeGJ65jCTcPmtZeKwVlPPxUfUY1uUmWe21n6mzJhGJx/6AoPZcELoy2buGxtcyoT
Heb4aowWeCvXNuo7FMTNx3AP6vNjXOuDIpzgJKzQIHFcclCVUdLWYsZHxrpN5nQqp/5B3T5nOG3R
rGVQVsfJlRNq4nu5kzAJo/b64wnObBdddppB3cNmT78QdPGLeqg4c3WBXYxwRsI5uGACA42lbLsP
2gzxtkOfq48nZuJUSRcSTYtb5KvDhCSo6pA6d6Nu11nXhpt1ptIz7rJP8m/ypr2EVEF1qdnpUdX3
Y6QKqwMJWgOcDwAIaykHt7ttZ7gTNC9ORj+tHd5UEwX/DgcliVuy+lj906zZMVHKsuh7r8mM9Wj9
8dM8EsqB2J0utMKXS/4DN1eZXrlBDjysJ7+117IGFZIv21Fcq92lstvQXXeu5D6QfyaLQ8bG7AwN
SgtrlmhV0M48/0t1HIzeLTSwqltMH/xb7bFKkf9Y8WZ6dnimU2R421f0S8jUAEUxc0uKKadW6OXB
hCszTJMEEyY/y4inmtuENazVhYV5RaKUQzmVUChhoaDMqzx9lIzzMzCLIk2PO+TMrTAtkiJaJd7k
PZ0sm2UF68Zq+miN5g3MowOOmYVVmb+GLR6d2SmUCaVZ6zvjs7nrv8es9rrXFH0HKWRDLmVydzO+
qxkP8tsj92XZatbRYig3yVQKlpfJIoe5C2qIpdsjUqsrn8W3K7eU812gTJfHpSscgMsXi0409eaz
1TsFcRYXFRFIySlQebgwrskgR62V/WtH8bwup4joKy0p+ffY+8fhuJV5Ah3CQ5PXlgl8yNouve1n
aLsKZE/bkE4W+95qKR6LoNo+P7OzDuY9TyZrsRYODrYXNuyX3gAatx9Y2xUrzsEQENY3qfjcmY86
J/A+qssacbTb9QQkD2EwCAuExiyOS696HN7qrNN8Pbos3PnW8UHKb0LpJo6R1Zb8EqltE3HjmN18
wD3OPg7t+FoA9/utHP+Mqz1royDK0svP2J/LYCmqWxYDwWMfOdSsql0Zc7FMRFiTVINzG3xpi/tj
EqoJwNwOBJoukiO9yBWIQsR4+EMKPqtZttHLeXLWnHPyKoqLjORiTaYAO0dtpFSizKoJOk4DVutt
wf4qhLTAPWU0AM4Xtsz6LTHlyHSMTr4wWDIzJOT1EOtASl9A9c6lh7oFy2JCXJ9q2h3porvdokA0
UYCQqVWJ74fLdh7YzRxX5TASdzFYulIPamZHPVwwnLwCofxnnMqWw7JzncYlVsqO0QCkc1919JUy
nTCDHh531kWMWWME2pPJqDNMCCyi/26Z0dRBjio2o+vrTQc51PFQzjOnUCVswGQJh9alC7ZL4grk
wXm+C1B+uBIu+HiVUtjC3FtlxvQ3/gJ/nnaESOPNEOOC9oVkzkWyV3SF7LQeqUG3wfEheVT6TaZv
tE25MrizU6XElPAfDZtBKYWJ0bCGPlUZKRegpp00HbR1l4hxHyV/j81XxH17fkpaDV/zLXrO9JOo
bFTxnwlLd0VPo0eriJ9deYrIWHT4cnoNDaA1qLGBGpttNyVDE5QB5SABXEpsmEnVd+imcdU+xzbA
UPhzlnwSckhqEBNCWEF9ZbA2p+SdEOWau1Z2/2d3vh8iUIxo4ukOHfg6htjOuuY+TTr0DtYYVcwe
RoQLuEdvX/+WusU6iE8OKSvylrGHKkEdjBGte2D2xc3UZMyHX4d9UkynsTQyND7jyoJpomPhDlUy
4CpdlCAhfLaNF29fGEfJkMniZWVvT6cRCYd36cBNfvGiGQQWzSZ3MhGxzw4V04Xj+u3jV6YlApDr
atfsMpfTJacZrn5DEIGCP2vkQroxJqijqhfz1N2jJpZ4M/x9mzs/Ods2STD5qCutyK8aV8e56qku
6n0fDTw4NAYR4tdw9hVAZze/oZPkj04MvhLIhQ8s7BXk5KIrL0fYa2EGb9+qzGZn6KYyscktcM69
jTUABtXUpVflJvUMmHPFNvSp8UE3UHL2TfmjIs4AvPvA6CeFk7xamaYoR2muha4yrLwSRCLBZ0RT
HS2WgY4Ra7O82Zg7cBQ1gwEhMTItJjUm/JwhAl1SyPJAxiErLZwsp2ZAQWGlSdUvfX4xKtuE94t5
6BjYltIgzg5KDTAiKY/iNnPe6rHxlMmd6gwnZzzj8wAgE9jO95yDQFC896Kr8oto8N2S9Lz0Fp6C
2ujaJhtzanM0AmC6SV38fXCB6Qc2wu469PelxWn2aI2q45o86cfDed+aJt75IarZF/MUzcoTac6r
LGZ4zTRrcokd7RfoPXEbOI+h9RKz89GigNqNc8NwkkEXSgEQs9fGGHI5Ke8Jh+59DdiM8WDfbpOj
SlOtpd5u40K7ejFY7ds44dSSTjVPuhgEjnl1ou4G4aK008t8eqaXv6NhE+hv3ruBHVvO+ahhJrUi
hOGj8VHlBCv0WVb/2Rr/yczzKyJJrqL5lKOjdls9EcGFahG+faXm+Zf0ciHnqatkJ5PSkrOQoe5z
pM3l6k1f8pyJGJ5szzBUwU72c7om9ErePfI9o1E3c4pBnL98R8s8pZbD0VeldXSWriyQi9N0ybEO
grQ5iDRtddLber53ic/Zid1sTwhNyMw6si3P5gd3ABzoYEfaR3lY3aGvMIOEi3vsGmqTl9IupDW6
dqj7fm0fEEgHh4fPzDD8gTHiPu9S1mx3ZxCMqS5Ox51fn1bALlhkoeSUnpxBEIhjPjapsCbNLfB8
SfJoZFEE5rfJI+quTIcbgm04vETrX4prjofTmQqouSQgQ2IUKljH87aKJtORvA6MPbMPv/rfZ2o6
elcHYj3nI0mWDODiYiBPgemtAWWfIyhtZFjAKgTWNZnTA4GqN3JxVa8sAC2gfesJ3KX/QCc7lv3/
eoRM4D2I3rgyaGmriKdyN3fO+mrp/TIQs+h3b9P/5CaooZKK9QI6RPS19k/fpe44DGSLp609+C5G
c4wiP4/whfrEB1G2RF7afW9U26VFCopdQBl1LLM+f4h/XRLmHWlgQ5OAR+HkB+1HZFnEqkWR7eFt
Re1wh+0k8DWaEA5ketXtNslUgFNvKZ5eQBPzHFf4YWLRQcKtpagAK76TEjIKogys9POk0Bq7bR1c
VpM5+2N/Ugrm6cK1FMyrKTxN4gOOjm6YjX5Q7QHqFREogw03KRYcvQpNuZiv/Z2KHLGQ9oz4bmca
Va/ExL7XnS0oBcqXNx6KLbvsYSaT9Y+xFM/RT88gDxTKtrZGCHyamHgR+ZQcpq+uXx7ypjv9eDMY
kl32m7rtTj6CMqkJvLqf4IiGrG8o7n/V2QWnuapcE/UwRO8gJ/PGHs2QKqrsMGlD9r3a/s65QmeA
UMCfiQIwhXf4E+Sj6KMkYB7i0DUrzk6fF/sxzu+eLACmfCFUdQIg8PJ9i5ZstCyOiw00zw+AhfIp
1O2LkcS4QTgCMSJGZNQ2qyP8h0f1QLhgZbNj4E9UUBDIWMiY/YI3euQ08OVNFbZPKTS1hHFPXuAo
InMC1RXYsRWxj845DhBwKE7vOcfJd+1znGxgS3GYZNDPldYM5qJxbxtWyorGG+7n1bhuNHmFnznR
kItwFjLa38RoJEcCKS6n6HUa3DUoKgnO0KBrDCGuUvX0Cy7crbkxDjfF3jyte8m7GTtyKhUYtCvg
nKqaZIqtWzCly3SDoTDBoDHpQe8T9jvfBKSOO+EVW2ZS1Gc5RLRbct/MAhCwyhMMmSQsMytnGle/
uE9NSLFTZMJzoe2pOLBBtOHPANOpvLku8ZxwcfVQx8Bz3bQPcMwT1xWJs5uf0md2Ho934XxWmU1m
I4JJ5wlH8RODJCSpNRzTRQVk+wh8jOQVPgzYN9XvcFFjrmCH5rlfd3enopj1ri0kFEOxsTs0+bQj
xHHvGRytlnk6L4Wo806aMFH5YxROYWxXedlWTCx+auVEGeQ5bY16DKYnoYmfsPhX6xzeF2t4AuXG
YL6e64OovDLjGsoUfQtmpwSXLtU3WjrVaQ2B6OHnYM4LuShbjH3WKhaC5gn7nPBZC7EYFcEKqgWm
aT89nMTCOsl+BPFEcOr+q7tlB2+Z0H5Ifm/4gDMsA51x1yFP9bg8/vbT+9Y+Qe9RcMDUf+ERsRrL
NFaQ9ToyUvoI9tIEUdbyt70ie7zNoIvM5mBWOOJnqEJT7c8R+XOq4WZcVUjf02yShtLwsA9OxhiN
1wGXLD9nixbw4pVdJ/luCjY+XwYYwCFT1cVl3xcCp/5NlX7Rw8L0wTez3NTmbBlNDIoKcxt47V9J
uogqVERieE/AWFOCEGwql0cQGGGtZrmFkn55F0sG33PHhUN/woKfj+qndnP57ZBgXTnOv/pQBAcT
PxlsURNN7dNVxaXUE5UBIrOXzggLQWKmMJtG3k+CYAjL+RYJ7Kys5yMQ+KOEKOMaWRCnn3a3sqh6
HeUfitibBt4gyikq/OUtG1Axa87Vk0awKc3gqYqhqybnC8EO+asLX/ugsbv9bqOmiZ+/wZOqmSVM
tc1jlfcMDk30YRT1rUuFa/RI9iGqHGkUgLKEeM6Dg5q/GPdUHZ8Mbn9S0ZWo1coXxGBUGtF0r7yw
58pP3MjhAdC/rQpWEg3ORxK1r2NSo5+6tvh6ypS748mi8IyUag+TERUwVzNcYr5y6LfJbIKR7cCM
w96koAi4m1KTLsPU2FkW7NC4HB83uV90m0g0yqL7UMg4Hd+OVIMAWD9Y63BKrW6Zl6T0gDRkDE/K
8WgSKmbtttKyC3CMrw50G83QdqGVQKEEoc29a8RauWGc+0VpeBiCuyVU0jnF/WvvwOwPi3OZhr4l
aXKwRF/MRuP3g5Ux9Qj+KlhSZWtbwToxk/lqYpPCJbpkNMIGtf+wJLj08eyFMs++u0MV7lSdKZ1b
nudojwMDdWjVK161bAxXpA3IhOBS+OuelrcCYCuvJzIGz0j42r0lrsAAuG5qdhjH9kucB41djI/H
uRW9/2cwoio03hJkpL3n8y37ee5XZlxQykSeX1NR5V4UZYV6otEPJz0Mqj3UGzpj9PeLBwyjZsRv
iEgYA383ac/Dr0CFeEZ+BilRMitDM35iKqnYrj3QHuG8HmGfQT/7R5RMaFxmfv5+aPyg1ymsDRjG
Y7UJf7qaRXJoBS1qtGZavlMyjnmmZFchvDj5Zx8gKzsCKFLDE+uwY5w1mvq1M9RvJx+rY1XLFdGQ
Kng/a9Orp9+A9uotxOgS9z2jJqjxVb3I+KkCiNlzE1CyBMRN1EQFCQgTb61xz452EaQ9y4AtaWty
LpvQ2YKjHQUvPAiaf7Mf58jqTgQK0D58incmj25TDaXL/oGNqCgEysabyldRgZSEUQdB1OX+IO4i
KhiOZYAAzV7nnq/EM78P5IK5x08sR3/ocabyLOeQSoUK4KvZlkD0SKKiA2WAvTaft7VZ+e1E96bf
x9Ka70q8+WeHBHYbjO+WeD8QcZh6dk2Ifd88DA6IJOe81GUNDPgqjES9dlAF0uy/xDIxgF/Xp0cc
jVzZZdXRlkMRKasa3n+ky9364KFBzWr0qR3fix/G/Oh9h89G7aSG9/09NyOuK2cdGkqVsWkv35oZ
k7R9/mRpMmjQSXyHUL6FtpV7lO1BBXWRSxmIax85K3WE6BhfXjGxO2pQmRrvbldsG2gAYhdmnGFk
7kvnDTXVZrt+k6YySzOtOIw9NaY7qjWzAPv9UbOQRL92ef/pkMxTs59NVTP2oUW/XhjsUwnh6IuX
UKFXVGKSDVt2Xgv3S1o4+FVNE+hN7q8OjGsVq8VIThSgCFU9DSXaa8JGYb/53gJCXLXO6dtIqoua
hBFnF9TQ8VGmpdCpzI1d9GnMKKbjWf1/jt2E4bXCIcr1H22caUPVeg6R5URiAxNBr/khF5jS0DWW
fpZfEcjEKPaa/3rPPdvgmb3VvLjFmrlQa33JZZdnYUbCQCwVKAGvAHIJXA5FuZ9Ms7TcHqe1EJyS
syV7bSawfohn5jP5QNfVN6ldCVsJRaKdWjULvrig3I7nQ27w7r/khuroyeHkRT0rnufIpLfY4TqJ
f98Wl6q7Nn7MSOwIbTVuvDZzkg172J0OU2hlArVvjWoJVvolT+ph3fJzPhKHAtfWOxzs6EqimwaN
aUqRlVMdXGpEbQsfzrl1KA4KBMccs4bOrUTheAEAZhS9ZO8HwxVD98m067SU9/ms7yjPO264/oHQ
/S6viWp62UwdAC5AK6kLmrKd2fA7gBTEDS6vrlWfBaXsBz3DqFdi+nSd582CTBhQ9fw0hcnxbqtI
i1n9dBEVAj5mzyHj9xR8LV5qgg4DuT+5QRWAK1Z2gNjB6I2zh7fdyg+dsGk4JGGht4pY+Ox3rJYj
U7OYUUjF1dPaSLboqJCZ5HqBuCydvkYVEzXWNoPNzsERMVuLlApoMeU6D2qaM5A/ElEQGOPWkk8H
6j8LrMzSq3Uj8bukLsGxsXRUfY4hgUJy77damnZLBlEWXo/bBt6b3BWdCGEivCnr+jpbPo485t0P
YdCAHk69uIwm73Pti4+ZCCA5E9vPBUBwNwrQY9e9cJ+jY9xXGUb1NDU0Z+29dbI3cSuzsczgyk+2
h1Xi+GasFjiGpYCM1RjNW5PvGN57/wxrd89Kl9gicuM/NoNBp3s46t5PaOO4uUNbZgx0Z5KIWBX3
ApWm3GXpW1VT6116eErW7iIZIMTIFLR4Ed40EphtFoUM1QB+4xTG3V50Mla4kCAQiFFeYEv12V7v
gNgggQudMY92nms6D+mlswXG4qJLi1lZvRhKH+yzG4ifwErclbMimxqPh/oKv+oHPxBvzxSgVk1j
kgbTosMAvEktxyu6QhISuDp5Jlkn9ZafbuNUmXOEfWAUKqxvYcza4TsW4+yAqyIycFbU1VZT9ZQd
5zljWDvL7rB42UJqGwy0NcQaERt6vXDZoucDcO0HycWLgLfv+GZX7T+cylUu7ymo78ZwpLqNhlsa
Mm3qt9UOsJTVb7vMrT3V3lCzWeIz4ts1UzutBhJO1CGocVQ/0AQjJRRHl+lTWFCDb9KqbIij7RzY
kCqlQmBxjKDYP0yL21OhzgZbzX+5l2hUtJgSgkJCBfEd1TcC4N4ZAuB10akKieoLz+FeD9WfOLwK
IxVJt9wF3O4ARyKFx77N7q/aY4whtKiOTK5O+ZWbBO40lRqlQYscdCXuUUqG+srD+QR1uLgLDsya
P7nJ8yMbNhKw56jw7/OKtSvg/TpK27C1oOLpRKjhIvAODhK0JDvAs2YWf+f0R1TIKMFv7SNuKGQo
Dbgso4uj4VyBA9zM0h7JuWs+92mW30go3EV1FUMqTvqP+tCxuMHUwAN0jjiM1UY4DGHUH1r8g0lR
ONK6CpmhO2A6fvJS3rR3jecWfTIEDgO7cdNGwtjDOKQJgeb4hKfFL3wyh9StSYd9U6B+qYshPF54
txAEBhB5PM3dY7eIu4h3SAWUbkdGvReDJ1kHtUpRgy6gCLc1yuJrjwmyv1FRqK89PyT6+sBGWKBP
lrmTYOAFNz0hih8s1S1BFB1IkEZdrJEF4r1dVEt90m/4e8SJess8ZWt4bjJk62pW1f8Tsy7ZrBmF
oQOybHYr3lxR2ba8dCKvjjqElYM2AmfzWcKHipxJVWQWIZ9/NXWxYDReCA+kp0yIHhPWuCTOHs/g
IWcbYmzKlPhk2gsBFy9eNYvnSqiLGkbp0gJU2iPd1odZMxvq44vVLFUVZArk6XcdcWnRnRWKdHff
Sod4rXJHZEUIJ3HpwjePWJAeUCUaFDWu/Dngqu3CgRHamkdSOVrWK/zjuYQ7CtCYf9z8SoktNtoA
Vnt60y/LO7lPnlkkl3m5BxyB2NeZQakvxAHCj/9gYSj+Qei5fJ49pawz/5NQD0rN8CQHp6DliFQb
yK8qwz4VNxtCdu8A3cL8wOH4VsTDb4QzgOlFjpvi2QFa6gGmTjG7SWlKXRxrJxPL3y6yRjsDrFz9
te/mnRjPMkALwdxgDd3hNVP9apB/3jAgY4qNnDZmgvlDo7pnXN5wcOO+FnxCrtFgzNNQFodYzWK5
JJ39NxapDYN+YffAdnZloirradhfLGvcrqHNv32hgRtUWtvdloei6F4JH0lvXypbZ7VUCjph8RzG
a5nJt0GkkYde8mb1uKH/IEDQkFu+0yHewaUmYTH3cV0+hHsmvctSlvAlsqyQiuB0tiQqUG1FQuI5
Qj/tbBIrRqCtoV7R0lXvit2xu1jvXuaWRQlRAkB3Vif/bPa7ePAZFt8R+soS6dOklzKp66TOoKxE
fWjiHX+Nxiq3BTnLUygX7O33KebMVkSW+wEnY4PppZ4JBj0u+H8fnD+6bVOhyPhuRoM1pgfTM2dM
PHBVDOQJaAr9YcUhnj3cD8OclPMfAR7iw7TtTB+dIUSA7tPJhVFPTVC9L0UlGvi9W7b8/ETJGXYi
2KVRclG70bJXmTkHlWdkaRIMrCvGmi5jd9sSXAwpdyiM6fAYZ0Dc4coOw8v+7GvAhtEBCW8dzXgv
0/RDEzb6OPBWC6j6fMGGfph3YO8QeIuVcvzHEg26ask7A32EmRdjskNdWep+jS3YTjRBiidY9+PN
yAHHKjoekcXlt0lSdw3ki9a71oFuOFgnWbZM3N2qPFotR4qrEGBq1krh/tUmySSEqpPHkLmtNGPx
DmhzysFQiPEfiF07TjPdf0Z8hDCxR36Ss9Ue8i+6XeNXnxO6nvZZOmV9gZSJWtdrfl7qsegScVeh
GYDjhZK4ACbDzOApGgdNDPUMZwzii3r1+vFapfYZ1M8Rjfbx9XNhmT4XhmtaXoR/06x/+5tQHDrq
7bs+sYuJS8LKnL+B0wy2UrrBEl+b1XnByFuoIhucH+lph8pI6/QvDLRgq22R9fDtxyo/ymWgfxyJ
cbesTKV0JfVarsF6Oa0GPlN+i8KFOJ9s2HW19wId9iTuI1b0VK5cVYoDLsdtUpIt40jCm3jr985V
YiveeL7RFX2cmbMXwBVgDXisVW+8eybEwTIV91g8OtY7WLB1mL5IET3vXUxEJRizGI4x6ddP+ouP
I1p7KRbknuXZAR3VSS4wdMKMnz+3XpwOim8tMP6YxmN2cIP/ShJCeKqfTkUXNB24jwPyuinkI+QV
OcJLcw/M2Wfubq2nzVhslLjUDDMJ+BlisjRDtuaKStRMtIOS6tOE4GZog0CcsnhwdSV5ubhl+Ha0
A9yXE4de2P4ANkv4eTJXLEzJhmKwLvyyNNL/qTKNjteEg9lO98epO/BrmlVbhImMr6X9TKYlLgwE
sS7pDZdxuz4Vpr+bu9phv9P3y8URnMvd7tYr2yZY2EYS/dGs7V1twbOejEGzmKEuQfWPuxHuN01Y
+wSnJ34FiOkA4u/OUcRO++X2CqUBb+N+oWkyxUjwsU3z6fTeEoFnYvlxEGJDFXRkhWiHrp4aO5Q6
h5X+g2M9Gs8LE2gcineKuKJR5YknYmq/2BE4WqrMBUPEEIDdgfCk+dBD3ljlFUH6iDBC8mofb3Nd
+CJ5bVl0IJwBm+JYFGKmvxCyOtaZ2xl0j+EC3SyfXdQmwvoAwfKvyFh/WG5Pxm8RFNeexrt+64wG
O4J/UU16jOxh5NnTZwpU00rN+qHulA/vY5BdmyC2wTNTdCX7P7zgJyGRvcvvTUGrmeVyFlhxiZtl
ZpMuhHNybJzVomGjNZQCulLsK0F0hKVrrXt7FD0j7MOdoOCGcp83xy786vnL7l7/o+4mRl86wFN2
/rpR3IzZETTWoUJjdsvNbkPsKMCWVOoHBVUkDazmR8EeJnyQGlC1punEbmoiqHaWxzNGKuqeHbw/
oGTMU8p/jReSEzwxMtXu2Cw+dJciCq1tKw665jYu001POQXgeALDVoUSJsKeKFvkF/bdXwYUhOUt
WX4iNVHaJgLvQai6/SjHLD7lmvjqVncVzCFr+mnDq46B0r5TYbM+GOkOEWDbo9Me8pooszcJMLHs
jQddsuGHvhwP3uI0ZsjB1x8yMl/IRV7vJB7nNH95qsyi0EPHkE5NWe48ail8O5/bvgIR6Q5DIMmJ
BSmxIJpeydwo9FX2IGOJQ2HPJGlldz//Go1MaNOasAt8VVd4VLGwNzioRfFnIedlwaNKSfeFS7b8
3ESA+j6032ZJQ6NM2WTKwCgOeFLUFXZCLGLJl651tUbOeEib/teHb5v2+oejFWEvADZ1p5oh8P/S
Zv81M3Hq0jIHfhb3LtpFuEfzNZTzT3K6ttC+xA7W4iWNuIfbk7vM4byluWbxWuY+6k/CFGX6sV3S
6uX7crVo4VoCn9LlLVcPVoRbBCwkuL4wuUNMwK+Uf4jeHUBsb/rij7+Zot0v15IKtmZ151QtRps3
svmvepaG/rp2TQEEkKc59WhPW0p6yqefhY77fn9MJuKdwg5WHsZMmj7RQ+PKzMMsjKbTZuBERQSo
avvyce46qAW+j5FbN1Y+W6RxaiXZ5y1cAMbcUt0Azx+Kb81iFpI0oKJ0J0oRzShmtBhR831pKfwf
0GMD+nSO3WWuscld4wKT7OXthh2zHcUGBjmEZx0QNY4xB/AiSr/kKCqJlyic9JRY1AGhEMysEwkq
e9dMA9hA6c/uYpG2GjoJPXdqBa4NRxIC/Ur/yHDaUlwojHVCghoCXWt09h48eGifsOiqvOg9U8dD
VDoylAqOt7YiWQoHOmVc7DyuE9+r5byeNZuKgC4wIEZG+mKBigq5trx62NETTV5lU0EWKbtU0hiq
JsdqaWZ6t00UxhIJtrs7fWaFDu1SwNg4ke6w8QAsacYMJ9ZzsbEa/QtnVTL8JRNFK7vhM8GFfqt9
Sg8fxEKlSV1FdqVNqgoKWBd8/2TWGJypNjvhivKl42y22NG9wXnaHRqd04uyqp7jSRzK5/Z8t/iY
RXkAUhs5H+d2KLf9eDSSXbi9MqqL4BDenQijv7rTZspJjbQIaXhbjb9eKFtHiUbjWq+wJ4HBtpCP
CuxJSFspfc1K0j9YpC2VPx+5YZywmUcZGxth+cIB4ZwtjTtgY6cm/uaOiom5RvpCxDBIAQWRGiCj
nrrUGnbOSRRcHcaaGR8cAeiyD8i9jrsC2+Pw1r/qbd01ZR/umVbmWSv4ANetNs4qtkakG5/7yb6J
qM96hUFTDdzN28HWyxt0fW+Q/gVssvIvuKuHJlhK7tZ216XoY8hYow2lk7+2BcjuuzBPsbyRvlNU
UYz5XYBWwE9grbfTM+VFhPsx37og3kcOjDech921OMmyDmD1pFZG2Vff4I7dnd900JpI81D2ubE4
vWbL7VVrb9rber1Sl66zkqfsbg4/17BvM9InaS1vXEgf+vW59q01JQO1XIBCkIcacsgCfXuAexmJ
B+L9xvKhvJDdze6weTXAXhIqO6pfIJDXgKiV5gDVxxJkYq4z45B8ziidRdQgV9BV4+kBlQwAIudR
yt37rcIPqX7hqBYK4iR3kCiS861q9iJWNtC9vk8OrX5/YFu5vmYrELHnnVy58sPJetAxWwkhJSBU
QdN1b5fio8j8bxBKIM5VHmrlqY+EU53dv8HViPM0y8qdCxegIH5A5u8p/4IWrwG5fnWm06GfgpKN
9pZ7uAMD5XH8rOiDkEGIwlpppzW1FzMWV9+M4ABv71m82l723YR7iofKImJGBcab7QSHDVhR1xY4
iBFk1Y/1u1oa23VasuQIiuwBKUTtHJmbaqX6NH5A9qWCF/p5eRgzrrcGzEy2hMWITA+OqyP1Hb6L
hTvhW/A0Lct9tL88zZqGeQyzUgMTEECoCjAHZKkV5yMRZrHQnaKDoyNWNI+E6POYUVJsyHZVfrDl
5EB2B+wpDDlb3s1QjNsRpahctvS5i6++v2T6dGBzDRe7MmSxzWGCh0EffIFiVIk+QJpfasdFGFhw
tiFFt/+w/fU+iKBmVD8yEzydhRyq1qMM5M/IIK1C4wyI9PhOEPiGrOpxhSNI0bcETIw95Zb8LnDp
6CRAKCRySTetFGR81IYLoHpM+1Vh2aKxKjIt3NnazBMfe17R+a/dQkX7jqYiCWsOXjrYRFpDyNv/
kUvNKgXoBpDnpyXHsZ3zmLLBYveJTmMnPCXBSBJslpdXl9kvO5iSQFWyR5kmOf7erKCcFlRXM/FD
arCa+lkbr8DLHqWptSQCfElv8/R6yMe6HFHWBmVm5sYrRVjh8Otqf6hhku5P4lyaaJMYd2kv+Ybb
5XcBybbeDcEkEeVGhTh8E0uuDJy+P8aM5yQBn5WUc3TDXmwJNDhQpgI4cWEGbfJJkRtEp5PH4+hK
blOdy6zc41bnIm+fTuBlMHFyz4e3pSwUGDMILWfXkTNH1bpuhvd5hzpknVPeQ6buHMD5x32AXQIE
hVR/WHa523HACLonBSmyAzSNEWtrV66lvXHVUMeurmEWQ6PSUBKEPg+29JofPSv03jgb2jTnZ2UD
S35qW7gkffYFxgd9USUj4eThRrGtJS0WAuycs08n2bFIqunKUvF/1hMwg36avtUMtZWot5/7UHDt
PlherPNaPb8Wk85n8pY2pHU2M/rhnzT4WhRNMKMpMFCPcUiRLJ8SA5XHI9PHw/c+MvhKkNHhnopn
b2y1B/uCWGRR0lRaV6k/aMUhb/q9S51ia0UhdMP9+b56yje1iWAMwqjxeDbrnalW+Wm3GaNQ0MX9
MhH10tRv7Jh4mKtyoR2I40XXzXz3ceV+2+W0WkeOEYGYrjOfR0nKc93CYEQ9VsCOMdtKPAu8By0M
ppXjsOhIqeNTjZ06FZ1qL15muNfImrQoj2LMqxwnEOlN7Ric/GacOnfWMCFwkyckEdmNbHvBBgrI
Fn2TNj9qDpZ18VOewbzyYYOlbeTdFOozaJi3Lvg/lUX4XHyZdhfBumz6A/P+NIZJx1RP7H9WaXe5
OQL8M8FAQbIv/cqJsQAdBJy7Qms3jZRNV6t0AksDvVZZoxLGSvW39JSmupVyBq8EgyBAx3mf1mFL
pC5nkClAcSGuZBeXcOHAZWvVg0DW4LAtZG8eZO9fc+8/xr+L/mXQJNTRMT/cIUgD/azAfm/3poaw
lSi7/l6b7jJea5X8xgAPkdrQQGngLHS2DhMl4rtpX7Ckb8dUDR4Db6PieN270ecq5Q/7qAgDdBcN
pVS0LQQfQCNGD+9BC9cJ3NHlZY7o0Ndsak7CQzxBajs4Ggp1JJUj3zllnprSQ7XQz1+wNqQemtJF
seOLM7Uqd3RWPZ+3cjsrFXpjZY4S0c6QZdKe2ZnJnLg1WPtpBsaRIcwamU+g3kQOz63+nmMyr/vU
XGsC56MeQRbcZFrImJI2OSgtI8tdUjWMhykIwG1ceBLDjaAcSCyQGcjipdjWxnz27Q/Z77u5wXoZ
Ud2mFUSHAN+PQNL2tue7nL2o/twv4nZq1376sSirfzoc97F2Ek1clWRzNwGBcnhYqSfP+9xQHoay
bPsKZysUygBXSKClKz7z/HtJwP4hsL+YoC5ovoy8Ljtg34+6/kqFWYuO9FsIxVjAx85vZZ2A1iS3
hGj6RlZyiszL0zqdS5kmqGVl0sYYkvsgSjeC0Kemh9QaoHq+3yvSjBoA4pkq35bre7/+6LY2lDa1
o91xBry1HNzvPND0VSM4AYJf8JmjmrfwCUJ5/ALwsN4TkCG2eoZK798hK4oB4FlWfbi2+m4cFa4h
YHbYKaJIjXtHQithW58JiOhC8sHvkEpyb515wZzktCMY1gFkpbJ7UPIparAyGWsvJQY2hQeNTMxE
9IiiNHrsDCEVk1Bx6ApkqfRK796ZhFK3rmkLRD9EXtJ+WsMCofVgcPQT9PKbMfanmWvE55bnm7hd
hhYHuo4x0QSzOtkkgoF77j8XGw+fJ36Vx/+EL3Y0VWcYEozewF7ADGng0aespjVlkdych+mFvKyO
esJPukrOqinv3l3l6bXbsHGGJbTIhRbYWkg1fKbPUZvrjhftChTtcvpPhMA7YEb545fav12x0ldh
Me7qI/AzNDiim5+sVaFZAiTdSmIr5aFjiX4vEzNZ3+VAzjby3Efuk5qB54wm3Liz6yB0kVmV7e1M
9z+sp5e2DekPx0urgAiX1j/80SNpvibF1ziZY3LlCYBWCPLg2kupNc1Vsf3yv5IFvcJe/naNLeW5
wizCHrOP/fHzDY3YzWItuOJ+2Sh5Ko1wQO9HXMystQqvcXkhaITIrG9yvZ7s/D1+M82wg+AP3Oj1
7p8GiZki73O82xVSMGAa3CKKe24BaVSofiR5k9v/V638nu77hjfrftdnb7D93OvFl/cleUSxwbuC
O4XeDXaPjTSDYaSz6SEWCB1PLKeefsLbXSimY7qB66+hAqGr+FzMSmORpxgrO3ctJKJ7lnOUvOtj
o4YuzBJESTtZZuW8w3LYOi0B3GhRWDwUutgtvEXDX+3ruPUKlBh9c8S2HK/aQraTibTYf1kEgMVG
b808McvJXlpTxqEO9FTh5Swj6SJ061BU9EtuLLgvRN2LhAXiPvlOK0xfFO8SzE2aSaZlm+vll6u0
xhulnJ7kSpG4jqiKCeZaq5M+cveTDxvIRKo2YxeY8JwaAU/uwb0K5KO1yevxTPhbxcEOKsDAU2e3
gb52YS/pixg+AwVAOXxESQlxATooWaqYE5VAiLzfB+pdbz0IeNVvOj/2bFJDpjdidkrN5a/5iY5I
eiOoZkUo3a9ero3CQW0ipFlhG4MxoarU7ziQdezOqLsSWuNMQyIMVt7WLXQpUr7vYI1nasjdgCsL
WAnpQO2Shg7ECgqCNqZoJnYE2x5UW6s/AMFuoHktoiZxp99rP1AN6NkRgnEn0frNbzmj1wL7k6+H
55V9FXTX6asr2xKYybQDtuDGLKMDTGXHDFiNMvLeH2RNtsg7lzWSPvtS/iPxnEWAi12vaBDkv62X
klv1kW73f9USl2vpYJno3ekCNUKrpyWciJY1l/GMhOanj5ql1j5U8SXVjEXvbhE0SNiAhvu1L3k1
a7kzxvxTCOva+auQYcL9NQU4i5pOBe4Z7EU2o3uegFedHNf+Tsw/qQANHmhl581beaXP6SvlBpTn
CP4MN+od5Kso55iUpjKhKyGNHfJttpwzGrXrZoHw+OwTJOcNVCjy4RAEuiESLyFRqsHHVi6Zwe1Y
vklg0VTpbKjXDTmP+hAq4MQCIXOJDIe3Qx39X78MmpNYbxqWg7gMLIOVRyoQEFCp5398GN9Q9ImG
gnZ91Ycly53+ncdCx9drM1lrJeS9g55FRjgAlH3BIB4pKFmjrTPCUCu5Dq/sQVRDYwr+WxLiSfmA
YHQ9bAJ7tetIDqzquwGIliTRuxhhX+8eTA2mt8Gvqt0QYXFRBS/h5uUhQJM+JCIN5+xIRvaOigO3
HKZmzFr1sl7ahdW9PQ6IeuiWVbjPg9ADrkYQqQhIunOceol/c0YACH6hQYgoPNyyUZUoCAIHatss
YB0pkmIL+kwOtQOowUAnACcjHYOjrz11oCNhVVjvGycpZlb1M+R98yHBOMDaxvqWCnBET2snIY5t
1W0XeuEqPYOPZq+hiiA+dVW1hx51tEhMchYdP2RqAv59tk4gPf9VTLeBAbEM1mU+3Wu98HKuOkRv
db55U19nWma0RX96eo2nIVfcHK+OG0CRixYJB7WJ1qUNRc3Sq5xurcQv3kblJP4qq4W2oWCl6miM
E5k4DvKY3ex2ZAQOFANSCvLc8cmfffVtUcto5qEyPHflpHNwKWeWS3z8S8820UpQrNjtHCw1z1ed
u9/mhXrMh8hAizjj2wmdg1nzvEHiAUCNdI2kq0NOnTOBOR86UyGdfITMnVV34wDf/Mi8PvL8ZfSV
eZouu6HVGNp9qBWXOJRPEHlh/V/nCSordEgD4Jx/5xHM7Cnzek03AL8/Q1DAeapBOgVLAvhHxqyn
9lojQ51Q75fK274+CQRN2KI6BouZ863hSE4eK+YUjLK+4wPbggDrIBiUMYyKHoisw6tj9LPH9NKX
Ia8CSRIvri/CPHbIUHZBEhDMbaYOQ1sPAjiIJkFUmfn5eEy42XBwQn9AEMkXjHv0XBBkguJO8f/U
UYkVVpPgPtE9/DjkRrcAO9gp2lllRPRUDXqUEVQBF16A4gz20uALEdOmQ7oKHw0357fQJlvSDotN
i9s5rKiFMSvo/KtZnTA8ZGsgaeoBdtkY5Si4uHhXlkrsWwG2MSM5/gr5kIOOc9raDh7FgBLhuZk4
0Duww5/PEwrBZq8C+8hoNPNRP+Y1xXR9FOq9xcEkePKSuXJ4XqVtKaEIsWV1fliLoS1jW9uVjl6x
SBvbWuWPI5Lr1EoIuynDWV+hfEjJhcpyWK9Zwqvuurh0WkuCHd/+EkMjtakV5b4AUT/stmmrGydD
sHFqBl1b6JIBzLJBaL0vuhOD5zxItJPKvtzW9r83/ORdSkvrB94dz33z9oLdWd64w1M+xmosEpTR
L6DjHgoIXjshmynapSqEmmwMpJSV/m9vViJZ0ocHW7757A9DeSG9CccjxiCc1ipX+PJWdgYm4sq5
ASAZAWaBr2xWgJ4Dayfoe5CkkfHw40Slnw12iR0yq2c7lobo9rDJ8V26AFrh6EnqQusVMFeeC0lK
G2fNZlzbcL/rxs9ukPzS4gKOd/Aq0bKFrECOr89KMu8tfxl4A3qfun4sblwHLzwegSDUyVasSE1k
tWN9ga66IRZSv3YDgszJGwAY6VooQd0mgobMLAPias3o6wb49cZXZHrFxejOBZ/e8cF4L9Xb2iIu
kvbrjQDlpNenN8dcVCUwsta7/SO7C8qBFeEWJTVGjzNX1Ne0duxqyp5tmPc/8f9kT2mfJMTVF6ri
JzxLtVBiplMvRxgfVO3VDXxhLq8+ebWrFzFOVqwmNXzaeYlDO7RWaA72LTPe9a5AXkYa3nmlyS18
BXVIN5PUpFtqCHmb4S6pf+Ed6mqWC6HI9rPSV86M6cbOXQ5ZxKpdoB+VOEYp28ZKksQDNj0/ziJw
oumKJTQ6mNaoLq9koP5r4Gu+jN/UOq9y6pR1xSrYkTE58q7Y0xl/N872pxNzrfJt2P1HXtYzVVND
XdAOh6+pTyzHzJy2rcdOUdlqlPHJZP4RA4PXA1dBmXR1FAHq2fF44d5Y1BlIb+dE7OcgR4KEI8EI
bRltck8PLW95Uh95tZJ7xRqL+4toxgYNuQ7fNThQmbJkSThVJf+KM/oyFAcNTk+nYioLkCC8HoOK
n8qylyuU600kLz34zlRxHckOACFDYoJGmC62opa+dIPgXiQxYwpX94FN8e2aGzM28gjd9jp0FDyZ
mvYZSw4tI/MIcJpA4vN3GEc7aPIUYo8XKBIapWnP2k2iED8ENm2L6WajVmzhUyEUUglJfQvz6lHL
qzp0GGUk/XfPnUDRmEilvT9slWObQDWx1iCCqkt2o6h9hIvpqDo1fObU5v08nAUIAIT/inoVCzCM
L28Cqn+Sx2Z51HxxFDz9VjmmXyqouWMUJOoUAhK88nq+XegDF2XtNAC4+B1GhZstuXe/upZz3loT
H7B/LLn06pb029pTxCGdlIeY8FsYlHGOa3KYhGn+4fljMSp7A0ATaOQ6KfOT7O4GU5O+m9GzqGs7
NRKDrCJC/VOubYswwq34MJycR2j2lq+dwsToBJ32bVhdCpGbpH9KYO7LAB1S9Yc9Z/FxaHIEAa0f
iS74FLUTqKC9TLL1bS3gq+15OHiLv6gW+eFpqpWm6mrgSclIrRSP1lPn/Bb8ro8c9dOBvLu+MUPP
VViCLwjbUYu/6m525e/AykeATetyK7laoNdS2jH3GxI26lQAmo9C2bdhPDUNnuFWosEDdLI5I+1m
Q7cjyeIe07iqpDt9ytUI+4A7plHdZu6Z+NNhFfah2mpUUzML9GReJuEsQ7PsNxMWHV+a7bOxiQh6
68vrT/DpoJl8uOm0eWAPe8aC/ogAyjWgFhyn5Z3/Hi/ob36kcDAAilaras6fvuinezO+iOSbBc1I
BJN3/IgjRj67++qLDQO7tWrWO0snOWr75MW8dmaYem1q85zmhBlgICm8hX7280d4X6l2ghS16GmX
7Njb+B6lKUJLa6xKuP6okP0jyCqkUzyBY2EhoY9+jLeGh+xUSC1QYfzK1icbcoLmTLo54Q8zRh90
ILPHFJx7Kvl7CnYlD4OxdV6SVae2SWtVN0TzbAoyr5UPDW9Fl7rBgaMkUYeS0WJ5GFfnGNNWt19O
nKYbrgSSXZnK8I21hxOrHBlHgw+unCUoBGpjNiS2VY4OdyRs0hLJsR+ZCZoWNwrkPRm/baVGh/0T
8jVLyb4ILyoz8mImwfIsExlo3jeMqrjXYD3MtescvYM15inX5JQTTB6CtnxsI+S/GHgy1m12b0C8
lftRb9oep0Dvj2Y4G+fDDegWl42Zuli7CXSu8bJCjLXbfsqAVplWtTQ7yjIQmR0gYqlk8aF6mdC2
lUNQjnpVOzycgouczbRieRwqVJomwPTD0DtUGnpzz6yHDgHQZHXdM4hlRHyPtxm5EpM7DklBOOCm
WM+Qf+8C9o6Zs27Uqhoy7zCg8zaUcc3wjOD5TcwtwpKWEsNcUU9rAajeLulAon73fGm97EAzsanS
6xSNd89gXVt8z60hJAw1afGhHdPnvPrwnkKb86MFAuI3PAnlz3Z8XR/l51Nqb+U9xHlnuOKhoc/t
zhcdnsaIEZaBmDrUz9GCTm3f0e6rJ/zKWsSgO0398bPdGl83LrWauOGPnKCAazUQt9uEAuQli/Vj
bQuk6VysjUyOxwBkbmSEydKh9JRhQEaI4hvwWlQ+nJ3MAjJxtz2DpAgJI5kVuy7xrEC41Blg13Vy
JhI9GywV0mr9PAyqHzaDWEDEPMmBUvzVFnIzS4BcFHgkADcU+qAbgL8piYuxO8qAQAd3koSLgnBX
o4VI1ZKih+L8WzoL9Q/DcGEbGtDx9YVSYKhk/i7AlIVFoLAySAYSJNdVx90cuPw3svy/SNSudHZA
JkIQKrV/5rJi8NrFzTrgce24Q0Kp7AWiuRWebOM23UVaKZpWuxvAO+zNr5gbPOu8frZuOWWuYB7J
BMt5AEXXQxV/u5phO8sDt6EGm/mRon9Tyg1YGVjvMQ+lRWo8YvmWv5MEMmOidOzXaI3oLVDYB+HO
/UJqVEYLYGjzLkMMmL10Tl3kJ498DG8cekbVLFzIzYl8AbJy1SGUzpw7lOk2SPgcwRHaxpI4ff0M
7sN7xN8sevQ7PMDHzCQhPd4l634rGwiaPDNqFxKh3TlfMevxUiBslyo8LUw6ZSxABYiUEBF3FGoE
foAAooZFOJPMcDQ47QjxvEm0NCcUYv3IPyExPrKJzwtBZi2CF1gb1h4u1mbZ8C7lxW70qAJGi05F
NWrl3QUFxjxmcYsDPJqGlpvm6nJmBVGau3Rx/vRGQ8Z39ZSG/ZtpSB/31W/O02V1EKxE7RN2eenT
yznJctbmlYaZhRpaOHBjgXIKvmfHDw99eI2aZcQ//eModUNX08mWPgdnbjN7eNnWJA73/upTbvim
4k0rZnyyGfwDaMT5rw/f4nfPj9SrEoXbuhNOLymnufudncRFKSHv+p/cyec1rx5e1i2xJycPkd8Q
JxezqVvBkdzkfmvIapkqMCvnX6oeIdxIeyM2xuagI26bHj6HW2AJCmmqHOyqOfTJ/puGPkl9RDB2
sqSYbd3/J+lO/ju0NJ1i6htNYClNZw1Hl4ZMk1PMRNW3oVW9U9jQQeQBoyjY9lWf5xD11IdDbPhs
JhwoHtew357XtKhHYDguneqcL1vzI++kOB5bkL1+o9k20brw/m1XhSRPZDd733JhlKeLmXZQoReg
KZWI11RPGpaCMHEnJdVoF9+aJJ2adZA8xo8CyIIuGlJcszwr2gzXS1J5vRsb3ZXm2AOzlwJxMx8U
mIdnpzHV4TrgRIyeURYaD0wsU1juxyNbaizeEnY+pyRozJmjIwknbzUtHRDc65MfoPNvqOLLczYQ
RExiIHrrXNU/xl0rlK1nZ9dGaPxNJHfQyFqU3jUiN7r+TQW8PNZKtwaFDXHZCbNHSzXxZ1LYftt+
iPZyUwrf5iYdSLwyhMi+oEXdiqEgtfvSALfniMdl25rQ8buOnDQyi9PS8kX6otNM/Czrlo3DToAd
lLtSnqTPt4L7guteM4I5L1Q0Wf3U3791Tz3/mUPi168aIgLPviXdzO5CnoSnTj5v6mV4iErPbm6t
nGIPJcOtHV7Dc5RXvgL3EKyKGDX0vOqveaQ0gQ2nF5Q1yw7u0tm6jHBRt4rq8H7T/JeU4JlSL8PK
5sDzsL8dgY6uwTzVuJLW3p76PIz6J1eOeLao1nXtdEKyfpILjOx2KHi08Bnq+HlwCumU/npJICm6
21/Tt8MsCDFXDP9jnn4vbuPEhvTSci4Cas7nmYU9evytDG/Nc5qI1zPwQ7etn0l6TlQIx2h+o8E9
XdJA5/RNCZvia9QQk6Jrukryyenc+pZdI02xR0pitGVQCJ/EmJ7PAzVurMGp/Y+sN8lVFBV78A0M
uWx/9qC4RyUTNLo8RTU3hQA91NrnKy1WdQ7aHB6t33MQOEn0eyI/W4QIz7MBCBSE0eWYDRgkJzI5
Qc3mnIcr1XmtLZE8fMJgvhdUN6+6nF3Cd5FPJpyOgRCzKLm393pWlnvpxdR8QYunUzAl5Qrzsmgt
ulmPjjrGrMN8/Ga0ZbLSZxW7CjwOpB9B1mwY2Dsbi9zU3h0riw0vp910set5ETOSkah1wM5V6pxo
btcZMggtTp+0tTHmYu8FcEOO/yIElKkzcSUxMy5q3pDIzmtQuQRgUFPa8c2IxrEyL0iKIhAhM0qI
+dSx3sweFaLffe8h+mQKKBziaPzvryR1O95XQA5KVBsOC/l73/kffTpgTBoW5pkdzFULJCaoWTHU
8IxWw98qlWCWiDQl0Cjbp3dkiwMCC8IxFAMuvin51A6a//tMc5udIASGOAkPf7d0+a/Ldc7IN/SA
mUeFbzPUtqWf4o3XKfjRUcKN7moGs49CReC9awaUTV0UfNPvSQG0bprqnDqIssdWqlZs7QuVb+8j
2Ga7jA+1zU5mjRWRQzanKXCDBU3672F9WgggoKQZCA0eHJxBiqSpwcnCoJZgQAfmQe4kQm6bKCEB
FB1Pf80p3UOTGHUtewr4M7Fw7HhOgBMgzY0cJLLU7XgKA3H8kcKu90SwhcDPu1Woz6CdBzT4e0XN
PqZQspxkto4snmAa84bEEOi7F0OpTVsGrmfMwXaM9TY8T+KZEFRK+Wrawdrs4n3tYl6toH9x9YGi
GWdG5BcM2tI0cfWHIdaiRYnalTQXDT22PQ3hCAo6e1WLJeCJ4fJzs0CYM6y3/Iw1k9ZnR+BOb05t
B7HBLqhFdKqiIO7wEl8PCvqVgfwbKD6wzDbQ+uk6QIkKeZCVd3d26arTBqYEw52NRp7ib7h8mQqM
ZcYmZfx29cTqNqQ6bgod+S49apxo9SwfE9UB2i/ba2YQRrZ69VWMDE3v2m57kr69DcouSGM98knJ
LlkDJOwnHjP0BU8AptxQu0y1TvRU9TMTA8sssAbUi37pKJX/d6zuhmnkP9biT+mLe7B5lq8yssjF
l8MjAkozqOjdBj8cMLiBZxfYI/2WLbl8rYwC0HEaI/iLmO7ISnCNO/w9uVxTu0JiOCrBd+5shqDq
83OlAW3QUpYjrk4f1InCY9oUz6Okg1POqrGh54K7PJthJqVbt+XbpU3Ktq1GjaFZH1QVZ8X8sjGE
FLoAcy5oFZrqNayFB28ZHbjUPZti9xZRPvdqaD2vBBamw4adgE8oDwwFT860ERYRBIebNXOyLZtd
gZqIJWetufiM2hhjxP35EuOl1TQNpcgmP/mF6LnIHJOOpTbdPmCzmy78ZpnZ+IWWP8utG7peT74r
ECA0XiNs3w4K4GTbHrvVmjbPIDcMwoyEC0Kvmjl6Ih+Rl61wxAYn3M4ri1uunJ5G8+trmDIcyqeb
efKeASBjHO5ohPWZbqNpvGv585Wc3LpFeheSOc1yvkcyRWTJ+w2Goler2izaGUmdN0Hn4c8N02cC
eMJdhNa7R7IFq61keJDj6JNeNadoXY35Bc7agOtvzteWeIWzGxoU9nlfde5X8OJlKk/uTFpYMoQo
8c0Ay3kUdV520BKZxiN2d0xTmQ3eHLWSp2nqIS+3MOeiIXC3von26L8N6b/kYbGo0EVrjR7JeE/y
I6Pc3yjVjFDP7FX/34EtP63rAdYOwVFCGExZAjH1VhrYf5d12W00L3Qw40ND+6o6jHPMXFpfJLJx
Rx5TwOp3tXEQUxJfqzQVZyskxFxdXKNKsRbeiNZACDvtI9blTtdN8LwCeFq/MtmAV1s17FCS1cOj
R+SZORIEabCVb99ISt+VH8/U3Ww7+B7QLk9JrjyCS65+aOseWpvNt+An6TtgIljl161wuEUGxKSi
r8C11cLBZ4lgvSKavljNY4NqxeK418AMxPEUtr36xQ4hJEmi8r676WB0XKD48gRZeSyfyik617vb
sFm+lxTEK4twLCDSfFE4RlqyEGnhxnifP0Ob1vcrnpx+mnROSGB4e40EKhquJEkKykr3XAGoXDYc
KsTVaAPgKAVQVjujssNHmkCTdN7vbSSrVJZy5zt+MdkSJFF1KzflJ8sfvZQcs6L3cyIZiwaoU7Zg
yutSV69/A4vOOtLrbbv+klS4INHGZqwC+AjXoB8gLX/3GXkaeK8i5kAm511B5PRHGYAc2+gAUk6Z
nhJwrOP8K8WNJT6JklhI0Hq2qJatzoAUUBYY0CcbqkQ+v/a7si6A4oOTNFFlBWTkF74557kFGD7E
sAFYApsiC3b5+Dr3c8qvX36fmEFDRCKuViqt0g/NK8b+XbAa07HoK0P/8rIhp/gZxmmcxte87GC3
wIXhi8naBRuNAOODSi79CFEJNmZ0reAZ8+6I5WEKjuXByjIUUdayeq9/4Z/lb8/h1T8ZY9DcNHTB
Ja2i1psmkX40z/ZB/ip7deyrZVqS5fESxhcD+t6JsJEo+sMjtlzkgAT3oHDMX74SwCKV0Sff8r1u
oS7t6NpHBbV6muYC5Vu+g2PJsLRNN1+kJ1Ei4wrk7NY4mSIqzPWpITCe6ewbuWpAMKH/ysSR0FEZ
R5NGFhOAsiVXCkbl4VukK6d+jTK3UkD5NyapmEcmUS0EnJTcnugMN8PYndyI0KLeyFZm9sHizoBI
SxaCKxs09/hScqXf6l5nxMQDPjgrh0BQw+0gn5FYJJuyH0G4GdGXkIfMgzyUu5ER+zxB3rYFCDLH
4TmfRAigCpNUo5ki3z5PLV9mYSCCZLtNW6lxy9xsU4VPMn53juD8hs3ovaoL+0POZ5mvmvpMSam7
8PzIlIRtXqohhQCpNCPacmIRn6JecARixQXUXXtYj7xt90g9Aa71TKybCeYSxQm0Wk9Y8W8VAT3+
ep4YnO7DPnMaW9gC+WefHs66puFno2Lt9KOM14nEod8nCJlFSZoHC+bPAHcCd3ekQSZiIb6SmTUF
sgRVV0JVdMJlCVTgJMiF2npgeKFr758DNd1/WRVbnYQ9mPn7of+hswOp+2/Rr7eHMy/3uQOJ8mPf
jDESR/gjSH6Y/gQtA25JzjcS2qTxQayMvcogFABeB6veWtOh1Yg/JkoR+5hq20GfJDKXgGkvEnxl
7P21dxJxZYs7B+WwJRAipmySOSfljCnrxhSibYJl/ysNOBvz8fPlbEe1whV2Lf+7ye4feB1Logal
D27GOgF2O33ryFps692FvpbNLliwOMh5TS6vBxmdSSvYTDmWjTmj1k80EUPGn6YKkH++YUdtxKUA
IIYAmeLG3c1+jjgUarDFpyVEw827QWFwa8W83sswDcBwoEzi3aj4E3Wpp9Z/KaxPlQH/2OZ9HrYH
9PWGsNHM8tYP4gyi/05jyw6ZoZAe/n7qEDHGzi9+g3/M27TNZCj+ncDtqmHbu/LO2D/xZ+pjzc0r
5ZYM+z21X+aK8lAvnKDg23KzkXoGT7c9D07oW/hUv2kXsmd+e+aDaEU4FrkwIDTjsdFLMIki5jFx
QH4sRL4AmL+wVkTkQb5s3Y2wU9GWnzW9jL49z8ZX0ARwjGm6kQVI1zadw+px+xNy0CpAMou1kE1L
HSDsnzxZbg4+bMJtcSyueFTIQLQ1aGUH8DrPzztQ/8bDgbOMFGyCI6iFPCBVBlk/2i7hH2fkZ7Cg
RxDrYqxwglibZJ1gDuMBad4mxWT/CTTC7MXT4K5s9DqKWzsaHt3idP9KBqjTKtfoVNPW+2DlrMjL
u96L4k86InMVhl+1FHz8QqRMIkNG+k4DSmcNXiQazGoMyHpsJh87KNlKFjPZDrRNg7yEkC4c5aaB
wqPEgsn5Wp+j+I9JGFEAfYBcuKC14Xkr6WjxWWjir0HVMMjM3OflQCLDJ3NF6f3nrQpubMpumMxP
MqD7E1GYa/z0CcRxCNJjaU75EWraLUdYnHLU4avsSkTp9yBhqEnR5VErShvNzZdvTtquVEjF74PL
0eb8cKXSumJDXXCj8VWUn2SRiqpal0vUNzNLfc6OcmDSULAvqUSmtqfGC99MuRedrN+9JgvP96MT
Ynvtyo8cGjjzQ0TG3yScSu2cxA7RX3KJtjNy1OnnU6pmWlPGLyFj7A5swsxMmjlnulA7ufT8J1cX
svsW3fApnZBMBM3mHgG0zHnCcwBvwFr+rBFOTds09m1fWlb37NjDYZzEPm+rV70KNVhqn7+e6+aV
xocWDHX17a5rLohlkng1FRBd9wP6N3YbI3i49YBMF753AIuA6aBzFaEPAEUbekHcqsof64vec7/O
Fxel80KWCg+9d3OrPqIdaqbWrYfuZDKMFIzH5uJNKPT4BIwojSNYBaMHytJvmVbIA3eBv1yFJsah
Zk9NuFwc1N5p9Vg8JNOfD4Hppgap28Dj1MQSKEbm9GKNixaAC8KuLOx5q2q4auxpznzr124x4xqc
6EHq6FPcm694HHpWJcwwFnscHRPlh4DqMwgwt5BPPqZnRcy3NK0ezhHbxWcn6HR4EBfX058YH/88
YAx8W6ATbQIfAvRP2ViqFdzyvNPuHaaU3eFzwZhedRqBOaelEr/59cD/tloyFkI++PqmPxlZXuCR
8swv4UUfYOGnSzP4LXNBB6OMS4FpoA7urAnlQqspNNYxW8ULxrTHkYp9sQY5LSfOayfpS/D7iF0W
e9TNk3ejRi40m5Da7I9Kum5uGBnJ1+TqBX3MkipZn59zK/MYeh9y2TBIR1NetOI0WHG2mpzMYgTx
KSU/fBQdozLXOPvd8m3rFnPA+BSrYIaLc7KS9GAkHtWG5APFjy4Ee6CFz9l67tnb5XmQmjzwEUjM
WzENZH9aT8/A7be522HIGp6JytXwuu2tIAy/51hyQ999J09KQtnp0HCGNz3JOuAow9/4PpbrQ99D
02RSpGy6/xtjKOIlFT2V6JtPsK+HrzUu2eu9+lBLgHdYxewXlLvA8y6EilTYTFpMdhNJyXYfwvtA
Z8vKHd0dz4eJbylzqGamDpkaa4YbNbuInTncPFq0hcaQzWLKDI1ohFJdLwujoaVLsqTJDWavOUKM
wSDON3tmwia+uPcRKdSxIQ0kQBNQT0X83qEANzt4kmoXLEacm6zRp0cPmoJu6iOjw4Zb+KDQdWx0
pDaie3lQJG21r3dUldgfOzB/yie4AM9Gd0iS8CGnv9ZeBv8GztZc6hyRPjraLmqHxpGz/TGgOsI2
njsHlIRyzqW1SO2YS50NZuh1+Fo1CMG6G/aVIguiK0hIHun9kbEPXL6nINPfYvlTdl1iFGu1M2y0
U5ltAIA34fWXKACLqsRobv/JlO4HWDXVOE24JvtM8M6qsG0XC9+OvwbmqJMrThihudLAxWx8U6vh
LctXNne5p9oNSmLKK2dKKAhdBSlQ8V2qTUsfrAW5U1/IHQnkeYDzfUwfHlDMndQlijOoVX66FkQP
CdICwAdOizI72iijVDJG4ucAewihZ6d90HtTDN1cbFFAdhh4gGh1slV9lC4Qzl/pIVrY6Qqi1dUt
4hSAFsvjF0KE/LgZA+g9Q6qaURIrH/gBkWsSTffTqXBxi4cFLTmG2I0gDIQCqn8HOsfsLQb07kTG
qoGB8MfUOujborCtp82bXlC/r5im4wRSK4gMKfGLO7EpwkaKQJahQu1NGgekiRkHR6+5xE3J9WAm
PZebLUPJcHo7jmSoKVOhVXYWmo3I9UrdBEPQ9/S02ZlnGW3DrdDTE4aYa+ZTs09zfXKNxIDfUSqk
lqgFN5kaeX4Y/wGlXlmGpwQq9UTOFXSJVQ2R+1wmJDViqgu4nxIAPYeUBw5cUGZbMtMQ1PgzH83e
D/9LWu7d9R+wTx7vd2wRuWkXusFQ/tVKcWq/1EiFFTVdn828dzRQ54jM2uUGJlNb3PkGHaDm4lMu
K3lcOTqkWWf8wUBB7Gf6Nfs0PXEcwSkIWlyRqXLquQ4e/l560a56SYK1dl+fGjaH1KMR5YFpwesg
UR5bZp/vRdN5V/2fmxcJw8aXwSPrKppCF2YAq3BdCW9PyNtnZVjt8EElDb5jsCTg4hZJAYrPAs1k
iF+BX3pfmSH7DxBDcmraj8X5Dy2S7MvGzeh2pbUhE/G8FjqtL8fcc5FQIfTKgmDE1Lz1zxqgj6KQ
IuIlLpKuVObuHbfuX55+NLXAnwoUNZsKI0y8jN/EI+M4flz/i8lSmw+oU5qkol+FW2x2MMbi8z6D
NalSQBaU41UCaC5tRdit6lswDt/BfLIuc35eqXKoCFP5S7fO40/092eVRoVwplyJbEEszpdg0Wa8
3U7ETTDRWsmg7scVjDc1mUhXGiAHOp+2gBe2SyYF47M7sHo37hvlKLXbTaZk7joc9aBk7zl8uTrt
h9f0FZle1GAEWTR7GLfcFZagrB2IHgPvhFaelYoC+5tSpstys0h3QvpjMsuSHjJTKUgSdHC4Pw8q
8/IupgGQlPwaEYax+rBHX1K9aRIDrL+ytcH1sXNETqSQZyKmMGWSK/sQ4lBCoLnkTF/vRrc+J4OQ
vY7ik0v7BDCSoyGkXSeqzA/jAQgdIk+JShPgdC9cXCB3+g8A1MgMXGfU16i02IFfgavtnSnh9qfC
rxcTFXtis0vtuPQVRyf7Bahu6JViwp25hp7MM6ERq+sF/qrYrh9lTqQLwLANmNlrPUDvdFOPiKzR
a1L9dOWm+BoO5iQ04t+bPS1Y3lMKvL7LMvRceUHBaualAcPFhFqBJNS38N3rdvp9mOB64uJc2/DO
/9rRQvzH7We7/SC19FAa1UKWUD/AmD2Uzlpt403UXlWKg/f56QKOJJQuojXamg7JGjulOYF+SwZ/
xQu0Mv4C7KHwf2YFfMj2W1PvBjh7Cw5ZqKltgugfxAaErAagelJlvWLWrrjGCzWgbKKNBBm/ZNis
JZ+RsfuY9+Va/V9Gjo2I1UwHLzF8qgz0PuUsSKzyDL8f4BR8nkR5ZE4QJT/FxSjs+HtfxANVFXPF
XEbqFseB4mrdWfDi6xMNEZhcJ7f/SyzOm8bSWks1t2tiQXjZy5zFd9eXJIH1pCzfHGX4x070Dwpn
egndytHtaPDM6f6Re20GT/sCHgmKrxKCpEIlbG42Dyh+3a0R1CkcnaVdo7XRH1zOCNwG6RPUab1I
TW7/OtF5wTKMYE9xv2Apped+iziTqkglVVqSNjElrwpfD5r9uVlaIzZqJFEbLxruqLCW84fkMPaY
GTG0WSj3XnHLyACx0I5lu/s3scDwItyI3pfjemaYQmqbh54GsmJcqCtQVg59Q/JdhG/PpSDFjO8q
+J3rVYKWu4fUT5jTDwqqzKjzo+EC9unIz/cctYHCaKypDALAFnFHXUKDQSTKgaA9rbK02roUBpp1
wlg2xW1EkMCInKSk84D0ym55CiyfU/nuec/XbUZSooL17duNTlhNsA50EFEAt6YlSC2Pjq0Jm4ik
JLFnyzhiVWsh44eagg6Yc0uI4ayr3LKZ2kAIT25fBT71gndXSsVYj3RGk1yGw4SOR+E1uwVt+9Rd
wIz7DFQLxvyUq6hGZ7F0zhCODvTbxJ5DyKXXy0xXpbyfvH2/KFuqqRqS5Uk+QkkFcjCh85CIsgsC
vlj+iE3MlggHrOPFv3mmlo/FhD7Oi1LkglB2et7L7IafD2b+e8VbjQlKlrkCvvuwz82KdvoBMtJA
bIfvRI1h8c+MBd/K1o6+GepKy5j8Nqtepi0HhIw6B0ovZaeNu9v4JIudkyQHNXS6XIg557Zdb2s3
6RA5p41BopB71TanQjHJN0NISdvvr0a7HYfW/98IvLTLsrc29RBJuGlVhXIEzOvns8rVM1hYcJAV
MHmjjGMsaeuT9K3MxfbcUIjCcocvLKdgq1NjJpeX8uOC9ajB+O2lMyTEyJt4iDRrIcaC2fOYWz/A
k7GMMho4b+wP8fxhx7LMJqrW76Oe3KbrDp6URY1GL2NDw6Vru94FV4p243Fgq1DVEqlUmQzWwHHp
mJGBPgBz3qdszuTMqYxjBxfS5hyNqykvzwtKFnSnHaiGx70DrK7xDEnSTLYk+Wr7l+/93roTYkOx
Cu7m3kd7gnTfSlP2nhD8YovGKiImQcjUAthtB48dr6MvD4HxV01Fz4ZLr1rNsEl1g7igjgEl0LzM
g3vnNEzRIhE2AfnhqTZw9sl6bSOp2UX06BgU6huHKwzzrIcFloQFOt5MwHH+Xaa2e8QffbTrL+p5
q1rU5JUq5vVxCuXVlZVFG5IEbJPf6gsAR+QkZNtKQTorytEZah3gV1aKmnFida4rG1oFu1W1LVFH
ouNXdEGsDilijYYdBX/GF0fAbkLAoRgyRDWwtJcwcRM5YFLwwU6F6haH7YuF2z4qPfzBw/OmjAC9
Q68616fkJzRRNdmNloFZaDYpRVBXcqkmV3PlBLCMm22xvEj6baxA3BaOJJh+JzQPXTGrSkkz+gZh
RsNde1FCLgsVptxLfttlGaLFNB/PKTYz8Rhicts1+zcpuPSDEnFRLud3oT/5/TgoatePSOCPbANa
ewPfQNGYAuetoLb8vMKr3LNR0jcNQ3+8uPKFr7pN0/fHBvdP1NrxQ+en6eQHdcyiptAJPsqHRKou
FPTq2vNA0Z6Enw4Woyzexp6ixllrkPaol6QsGc/iM9zS4JW+QOooIpnUZwHSPo3Z/JpNsbLoKaR3
IWlPO3pP4yxkTvPHGzmewztWiIhvXGGri9J7TsMlmIHIDYxCaguAan5VZjjDs4TrzMf1A7yfXLJD
WqkeyBRxbAHnrLurooWjyAreN4Mn5kAMtF9SK2AgRE9EcUPNmK9mgPESFq4xTf0gPDL3OoKGhPfh
AOgrtKVKqoixrfd4/W99wHjjWGcWEFGJbNVUvjvBoWZu2GhGdanUDpmvhXdQPes6aBlMlJmmySHc
v+IkFMPk0v2sGjVh6nVNwd10IO16SoTMRPshc8PVFYSrAQGUTEHOlx3PaqrEavfCF62MzoJGI9+h
enGMUjYId1wsTZz+563iFRiZuwpmI9JOxaIJ3svSuCwnU5SH+BmpA34uty+jyiyOfRYZo6Iu1gsF
FAppa4X/k34SJ+EOshOvvMrGMj9c3uHuGIJtZoNS0q5LfandB1ykV8Zy2D2Yu/5sk5tUpKkymcON
jN0cudKHk7/U6DyHzRPnpW9Xw9on5cCOjs8n6FUkycwZW/7WUYzCsZQTXQeDC2D1BAmJdqCsi810
x57y/MHl/bUrHBqxP7o0g94LYx307O4cfRNETxYhNcKw1OslNAPjby/LfVISMKEtz0wFTShmD9OI
vIjuKWUrMEBMId8MCeBYJxsKM9SEn3uWtaRNCjIdf7e5U+JdqqZe40DBxadtBPRlCtZ2nGB0N8RL
k+2jZ0Yr7zsK2C0dH9Mc8SgIqGD3ohV9hOiTwDQXqdbQUKtLr3LS4xeleDcuRCs69UL7Xl0k0nJs
IcTxFN1jXDN+L/FnTdIHn4e0oEr4g7ihC+7ytnqSneqZQ6qqKZZAPQj//YWMFMEAZcnjDW4qHAa/
Smwb1WciGpP3PTkCEwmLCVTI1/R53aSZVagj7pSshuHBOaf8Ghs6qWAFY7k50X7I0kulwNz5Wboj
sY9jxTpbt90JTRB40Ycm8uYp8CpLi2Z4RfLNj4jWmhtbI7mLpsSFoN6ydv2/8K1EoxpiQeaBsSUe
PKS6OU2OeqJycPvTKgiLMUb6UQSeglIUfp1xhpluaAE6J9NoK3JNJ5D4wUQVZc7gE9cKThgtECiq
bvT7IuaLySkbZEAUd1j0U6RU3JiRjcyBhqhVZO2lc31/3hBoFMFoMaRwztQrYCehITsHwJnBP2kz
NZUdetDCDtP0v8a0XMmTyvy5aTXvtL7vUUyNQy9/PHYqT94mXSKijuiPiokYnshOpw6SASw88bqL
fH0Q4XbfP7Xh4s8kgB1W/XokjukLZChB9e+t+wavp0Dx9emCuMRixzWj0Mln+vqPE2uxB2i2nyWU
d10kM2gWRNvSe5+ILOIZXQSYWqWhitgWKeI1iMbCkAUw0ehQPcFkPMXLZnPVpl7AgPfMvQXF7kA2
NdmujtEkwIw+joaRJ6mp/vloTtIgllqfB/bf0mhhZRDcbb8VO/uDlU2bxmC6NHJfMO9NJeipOrc1
WwKMzngaYnBAmmzXCnLPsuFWkTzYR/2P027o6k+L71u6palRtntvZYUbIZA+RnpJa0hWY6T6mLjj
eC+ne4WaJSVz8UaN9AfYcz4MQ3F9h8S3kILGoXqkQPWoRLZ+LHOUbWxx3BJELQEVmJKbSjqZI2Y4
nugkTIsPzzTyiqr5mF1RiA8uA0r9nBsxE3k6ixezlmKoCCC9CbpibiQjcP+AfqCofqPXYNgK2bSa
zLdW1RqkLnaAwCqGmLKN4iu3Jmzw5heIitg3Pxq7mMVYgcHXhzzo7GsZKgYmmGL6/BFXz2cNffQg
+JqwtV4Mv9Gu/s/8rU1P4ZL7qgDuZfITtq8V1SvXUI76+QTEmQf2NqHpysK/dvtKTsgyf1uk+Amj
VXFzW+VnfNqeta6AvGBVBGqoj42zo/Wz3CRFSmKD69oBVIR00CPaY+ZDyVsJgcQfM9OeL5qvPheE
NM6s7T7TfGvAzwGBOk3/4FUfEcRZXNm8R1O/afI0K/GPa4LXKjFJcwkqwV1YxAml3BanTLTM7BKb
2r22XixPZyLgjgqy1bOZ/iFfkjdessMOCZxV2o+/nIRmtCDglesSBgtZfQWd7QAuAjFamvGFLIXb
yRw9z3AyaiaaZKL33xJaTx8sLyna9RfgRvU2BZHdyBslLdoWGG/La68jSNCbnnEVWKn3KR23fPt4
tfF++UraNF/kWX5vrrqP915lWNWQWKONIzxwZH0kfRH4r7XPpdYrI5zKEPm6mNTJdpvUyJuCh1GN
UI3+pvL9mVHG+Y+JjuN9+DUqurArmTkr5cm+3+38UgXFjHVsiMP4t90Mvq4rdW5/mhXlfQou+34C
fFV9xYM4KDFID+iwwIudAtz2YULzsbRbUfeQJF6EB18skFOUGG3oiXRl3kpKyBoSlqcP+GTKhHX5
Y6Al/jduedoSGxXL9xNaSZwffSGu9CbJ1ZjlaAofw7urR44cX5b6HsHqY6WkOIBRnmnyxFtgX1JI
SQWgLSIeMBAqCpJ3BuPIvFfd827U+TdwaWMBCOs0a3dc6jFUqEooYo2yJ0i6f/t3OCj9bjycQHS+
bSXLnBN8IuC3S+1bXdK7Vt0xKqeorckWVpJ1npVqp355ZHlUYnUp9IwHSaLJyMBvVfSPazNJkalE
Gf5QaBhwM7FWace9rn7YBPZNgBxBUfCDHXlr0Ndx3TiF/eU7kLpI72Sh4it8TnIJwP3QXHmpQWgP
w0DS07W+H3Q4wAPllGzGKPj1hkjbDtrxeW/B3gPRmBbHiXcXFiEYIHzu6Y9seA7YE++L4qNo3lx3
xj0Nxy6/ld6lsnmUexQ8NfFVvD+Er/baQHtlH/BMcCvv8uZkdeZZHbdpk0p+ce70WgAOVXmGhjJ7
BE/hYDNzpc4cNj++wj+l0ASrrH3TG+GB2DhwMeUvfee0kC2xDhs/T56IfqqhAerT5Vdm73/2BgwK
swXfok0U0CR67tnideCj9HA8iZC8YedBSi8IVl+gk6smJbV263TsTQhU9pUq6wJq2UPi+nnayJM2
zAzRmrf9lfeEj4g4w640bA67ArTq3SoouOrqMRlC5wlshkkyG8rdQcC06mn0wwtVKM5D+XuX4mNM
lvPze/ZZAdhzm+VVGmKRiu9hCd1IulLzrKTooJtWV/xkOauyQBDB7SpG9Fykh5azpIiKNzo6OZ8o
0xsWL/EUN8zcj5kr7AXP+22eWX+i4zcudrvzdNjQmbFkAd/G5ScYA1/MugGNLS0EZ/o99Jvfa2TU
UGEnj1elZHWB0hEihL34UEjweUfg8Wk2Y9Ruz71AD+3y65xznS+DqF3qKSPczJgmy4kMK0fYq0Tr
LhRbQuyJ8620VweFRgeCT7wqrgrB2tj7i8pq+FL0IjR3utumm7KyUuBX133JGhPqLPQCUaoMv6Mp
4Tg4usjx9gfkM/kDwASJO1adquKk143EaYFDwYRVaNfHt66y3zPBY2PrHtN4NwR+pNTWjwjluIGy
aPmh/scDZOf+pfwafuS5CH8kuhn2qgFFk+Q6LMakecjLN9ZKlcvqkjoDAAP1hclqaqImgIxQfqmK
WCcVG97Cm8Ugi2Q8VcpHgwiNCzH8DGKs85H9nw5ekRMPKYxvV9hQHDT725DZyVSGkOj8KqsNzTRz
yAOHZeLTgp53k7Z9xhXH1Cq1I4sM5L+XvR2XKNcxVp9Hi8BzRpIdL21eRSRzpN8wCp++YJ5p9bRt
ze685VtmDZmGy35FJIsheZ0bS1YRGayTebB/TrZE+C9OWQKXRbp4sEwtsKoxg8P0SNtPGWXqCqZM
HX5OadjBK9eWICnoymet3cXIJgLE7yTC4e7Em6VYnzya74UQYe4GgcceC+xhQ68jSOE7l6U84Z7P
qKbWnqpjs9pwYTlpE9mdAphR4cIi3LzpGjIaJrcHXSYrXoGDMkC79FgMnhr5Opm/P2RW5naKyj2W
CrZdW51TLW5xLuZ1IGX/c89eaRM1RL05k41iWUkWzNavUDAd217RUiqyDDh96UgfhFEZBMZ5J+Lg
LqRaf15e28sKT+buzxnneMuQltDEwJd2tgkOfWKJhJDyeXdWB0TtJzske88KUeEf7EeKh0y2aGaW
PIxyeLDUbBtR6oNufPIicZJhduY8R/I82DJRn94y/3CAc4RJ58xQ16OxQOv3iSHTmulR74nFkNk4
SWdBt53cw11i93S5A6OXrE3fxP7mkV8aA0WQdjPas01+xYEmrJz+M8ZlrB5KLR+FiBeY4CCeFEuS
JLS5xrvCkYgoaOm+LGj2m1CRq5p1iWbq4yv1RVNHsdmi6MxzTK7hG5js0OB2xMEg3/rhROZMAkji
Xu1FFUS90/yLNvMPx3sVM7idCJEGyTRqTzXpcbkDxMzGYIPvlDL3eZkQ3aMcB1jS9hIn1vxvUk3K
nLmftP/mdfc/MzrDPsNQ9UcU8ApHpGjeia2j3d20cEoGuLn39b23IKeCG1LLGcb9mq42gnFslgDy
dCUaUZnMX0YHBncgHNMnrob5zD8Dqk5nuNccVCqfv4rgdXWn6OCbxCm8PRxt1XTSBOEansvfIHib
9QQ7Z/QI05SLsz34ELRiL+mmFoXDks2rfVGXqeasPRQgvzEbk/0+jndEaam0IwIu6LzsLLI5nFrc
sVf9j9mtBwmeOZfIPvzWmkx2xP/S8iLd0LSoPBgjRMIZn0JYiJ/qu1jJhM5hLKoe2K7QW04r1GUB
WqJI5lAVC2dFvWdAplG5IWs1upYbG4R5PflAnKKGiF933Am9poSIMgTXG5zq59plJqwvhauAm6ys
7ONyhkqj6vcCIEebud6vWtmbGAjwHF8690yHnn4eRP0PRyf34GyCmJIeEeo4dhTq45VptPegyBUP
wnNk+Ur+T+hoDC9H2TW1IuMyif/VKRtYd2m/N9sdE6S76HoTaeMFkmo4VMuvKWgUIKvMxhNsK7fA
MEjkZQ8ynnQU0xDehpJTHpsudq3qJSCqnfTYbdx+ULGGTRSa6eEbEXHAhF9JshNRsZeBPJuSsB8b
Tm59UKTLg23sT0d9WRRRfKJ3wz/nBVU98by6aee9nmoW/I29vcxzfmDjLV4b8iL+Nfcvhd4EwdfB
2FXYO8eotg1GZk7NFTkxBPjzXzN/P7Tuettas/dy5kWiaKGZLvUL2/fInazFO52UEOCI2EoRUbPM
6e9mlPhRXHMJHxMj+sPbqunOCf48qPhMcHlSog46op7AySoeOwwwASgkxCYJm/pqLxZPWBLJUZ2X
xUbY5c5yUoIhfT8GZRGsYzPhXp0N6Q9kIUo15+WSvsgm9p34PlG/0l59OdO2nl63U7S8pDIRbSus
mKhMokvCCGff17TTQOAtoyZW/+wEkCycxGTvwibX38ITV+IDJ8Q1yWQ4x5jci3nYDwzT+/Bas57b
hOKdoDVQKPOqLKUUv+fpE0U9ecb7Hfns3rfW+GLl690pA1hQdH5/3+zhsvYP3Bge+I91IjBYpXpS
PHWQkgvZf2vrB0R309BxA6uPMVPfA2XOqpXIiFf1hYk252uqddasKdYmMv7zLvnfD3weh0Y4vlzc
5OWZptng027EQM6hhYNm50nEVfOxQa1R9GyHfITJgnr+RiB6qt3gudsUgHbVpxF3FPAV1osX3Qe0
RZgbWwltzyy0Wcu5pinQen4klbMxpvwYRPB4nQgI7lEcEMjAohx65sChsaddy5BNsH+qPp9Rujgj
DHwr7HTw07upahBKsdK+zsuxXbmkjUp81rLvJcp3bHFREZ+8kQlmNxjdD8EDCNdfHQTNAkjUkze8
QLmrg3fgKUAMo3d/KI7OPmq0xNbn491bnVy+G8AHZRv931PdFd2e0etYT791nWpomzL8c5fb10pV
ADuJRUTV2iBcyDAoV+2YHp4dh2lEmQeGIiv1zQj0KDtB8c14SmM/MubxUwvCh9CVZ+dgLL6D3iHG
424ZrpZBWNnTrWFH2+xcliwy4umCC+oD1FaPP3r97uWa1KmpIfJizuAHBTR7nT0gtSRE3aSZ/eB7
vfXvXcaAU7ErarnjfzcXXxL1TvUE/c6cTfJRWsJFAi3mse2omU4KfSPUX4Fo8r3D5NBRxGuEfqnQ
mq9arORaO/XITyLTJJlXw70M2kFXIER0mo1g8zGCybzFcYODqdHaRSnamjOaGqWoTw+X640viGv9
TJhi7ulpMwhReuIOVqpYMgZC+GlmUlolr9GqON83vsc6PFV0o1m5e66GL6lkt2HL3lwI3TyzQ/z8
s4uopqudw5VW0z4nLEcjcd+Ski2t6mr18lG1G7AFy2eInC6Bes6kXmH0tveXyjLYYHaMEAg1iA7Z
A1a9Pb1MUEymDPyx2g7ZH7YamPuSqXdA/68g4DOjeVG1sCMm5ifXTBGwWIvyuLltqC4BOdntkX3S
viZuMB92qOXB7b6bkp2hCuXR2S/QZ162ICHJj1zPuT7reQVBDYQQx8ABaaon7hkLaYy8UcNyiqYf
0j8wC9uXov4IDHDiVxtXrX+OWi7Ln+HKkqaRkZpX7CyT4dqBGY/YFd/oOUrzzQ7NsPVpQ+nAO+R2
EpNjS34fa+h/7+G8V0ITB8Db4mYPT23rv8MviiSoMhKmVDkYNSWwRx9/fUnXdlg6Bmjkz7lZdEcL
w5qikif2IOGgBshOJP6GwqzjJA85WpxpCp5bVThKrPBffEyQ5OGajnPgulXyveY50xuk2TEBHZD4
cckhRbG4Y1jboOEJy+fAzCMquyFIWRniArxfUSmrBe0OVZw4wJ1AnCPpbH5+tcCGgn92KFBlifkD
apPmfG0wXxCJ2xV1FpKWnnydmFZZksUBKCICOuXwe8cR4cK7CCNFL8CZ4+ul6XjkSF+6vztdAuPX
Vlo3zdm8ZzwmQdVzESqKYSd0jmFYt2KQLzLb/VbgTuZ1dVGCqO5JGmZwMuNlU4rXSMuN3wwojr89
v3AMXif48br/a4cXWnwBGYEPsDRHZltyHdF+jkX9pM3Dln2dEf5f6wobsUPD4aPMaPaAWFiiofoz
W3NAppxhXWgcXMC9CKf1wIhKHYEAEA5dppgftTMGggpTA5FZ+ASGTzAn6Kq/frz+0pNMfF4DkRCB
dh0Sx9BAzEQjGNu112NQD4S1rq7LDBAcfQOwAklP3v7MGkwKcUZhTDvovYKNR0+xMVjpVUiIvffp
HdkkW7CAGGnaWuvyorxFkGgc0B9P+N9rRXMcUK6JLEhBbeyfnaFkvtA4c0d3nA+2jVCG0bkzGW3r
u2DK9svgGJ59mdF203BCUtq8mD9IAyVUKZEQAmL37vMCzbd7RD5Dr85vokI+uq3wsuGGC1ATJTcN
WuCrtCfLiq+WSczu479DAUuJ7Qbmw2Bvlekf19f/TPNYHELmsKqErwvj5OZddJY7+saHhCf4oHEK
EDJZfykWiB+Bh4dIrOaQLiQA4E2l4qOFQjoB/yeSyQBJ6F5XWLn8/fbBXs/kgJv/knFg9oJmWyGT
qHbZK67crPlUx9+3KMGGPPYd8rFi/1Onz7CbCO62gA8wK5EF5U1tnHjzXqsdYs2mMnYu7UxUHDFB
kzhnHwj2giQmdrypSckASOKpGAgOSkkBUHOG3yvP6wvX7RS45YvI3sxuG0Ji/PK0jczgVjpj3Nx0
SRVicuU/O3O1atOfnzU2IAsw9cz8+N1x5QmrTaByE86MqS2QNErTDKm0IGRZVL9m85dBHVSofmU/
a69vlIpftIY4sEMsTzHHlAMcRf4o3ob+d7LFr8le+NK0gA92Ynt05GVHJ3dOjQMaIBBjncnP+bDw
YG3BqoO+4vdg/g9k+WX9JJlcKzWjkoSAz9Ir/dGRfUkYyjbzC9hIKatDnTZltAiERjcnhD6fKOjP
laAayI+jfio2UgnYcNv2QNKXFVe1aaGlUszs+56oG7TxjdhPf2Ui25xbu+2S2C9IcfefwTYmZoQE
k1U+y901L80vJ8/Pdc6OQJe4xhTBCaR2J1Q5lvQZoItrMi9Ju4g4qjxkFqSb5x1xZRxE6Yzsg4Cl
aZUMkJ3mvwWeVupijMCE/85oXcpNIpJ2x58u8+6tyI82Mv6gxGttwBePl/jDxjp+zHw7oVYjyTbw
ddo677N8sFY758v7DrTj8YVEGoalTNWLFtj8AbtcWNYw5QaEBqjcLrZUlaGPwUanIzzryzhNpx+j
FxWia3ZKSqeJfZaLWL+viI8KRcZlqkHdZNNbM5eA7VkzBFk8KBPig8udZFmJ3tK+mMCwWBofxy1W
XfzvapNuUHQuns1WdLMCpWYd9+0oF3qfrqDvTfAOEnouw9uds/d/6lm8x9n6ElUtFKq5w/aw0geJ
p6eC1xM2r9/eBHRjOe+l3jK/QLx/eAAE5TlytjgqurWyH3pMI2PygKhTwgVHEt73eUN8Iu5c/i8K
AnTq0/CDbrHwHI98zPyNqNUTQZ1YYBG7LV2FBmXtnJaW1muSps0vlwfDTX495f9Y5Dg1DIb+gQqp
AqMeyN9a3JsClIqS+eaC1lV9+fN1H0eSESaJZPnnFEF4XSbHmVd04KWxzX8cwLpx5VvL9JltTPLF
ThvK41ZL99CHIQzSwi2yBUUwVNLsqhwlhkLsfdlZrEVqXTPtJHZitn8bgJL2VtW7U5a+06/iTvFE
oVFlPlqbq5yWxJZ0EhlGtDl2JTf1HsTQsRubOzIgxpQ348JzQEz73MgXNYJvWj7tHLXZ4TQaManI
gG1jvqquhOvWb2dAyX1+s4G8Apgn8/NnrD+Ny/17p3JTPk0UYfpMSOm7RxN9EUcYEZCirdeFMeFu
CEwp9ALGYZSDKiSBr2ikhbiM/hc0h2KVBilefl/xyfvQ5O8jLve5TeOxpszVa8BI/tM2spmEnIpy
jyOyvYfSl9Hop2iOzWyuB4RVkcd2yM8HvMyvKgd8vCOAsLNzEKLt5PGIbt5udVnh86MzzhGprpqH
9JEPA4TMJnIFJwJa7ZdtxH0jNUqtmJYcqke7YTZrY2DumrW6zeAh0CdFCXA2lxwp8JqlJ/dk4FRX
88/O2UHhz1hDV+SppY+v7t4vg5W6d/MK+kzYedD0snNUO0yItVWWuoSkH13h86qy1IcWfQKQxgl7
C/eifeziQaidwVuVb1DruOA5epGWlggsuTExUi9r8SfzJt40IcQ2jRheBdu1AeeZY1WuCOdtSmZq
1P6sglhp5ldAps1ahG4ayZ4vbtBdIDk9dcehT9fFz86NKCysafph4R62G7q6SbzzI2Ojx+3V3In2
lIn4MEK8A+FzyGnH2mEKuArla3/pqa5ie+3MNxwkix9idpwbq7Aw78OhYltQfTYJVzyJuOWI0DtQ
umy3zOWyF9Xh1Lo+ZXd2u0tjTLBDDFG/qhfHyfYGPTbfz/Zz9w0A1zMSPoJOwhxW+eoW570+Wx96
heSHoF6J3K32reaUKLo2lOGDMxJByLr6//Cck9Mypaw4bCQ/xnl/nEZsgKkCs+6Unb1CQOpPNaHA
KoiS8v8sfxDwZyxoIW1u9EMQ9aSKvAWor+y1XwGOK4h6fkp5mtpKEOP+sgHoYjgu7XEidv4LKi7q
+zL5ACrsuirBHZKGyK9g+ZQoOATfhdi6X+dZeetl6hZodo6KhxBw8C/NMKKP/esURKAlS7U9AVxE
7ruS0ktfY7sJaZ28y9TUoO21XApCW/Yye8m6pw/71UCqLb3/wzosmPdVdAWNQjvJGC0EBsidiTDF
9p9SuVI19AKavGIRH3NlyxmlnUDV70ObDTQn5j7LezR+zJj1pbHEHkAzP7wBNNG0UmgDyvyVTvdR
CKw7Lz0QWgq7laVzTF8/1MQkb52WpGk51oB4s8NZiFUvD8QQHFrsDweYDQrRmByg/aWQRMNTmlew
NpRq8tUnUxQ/F1bo9Tet7Og9/IZ5uLCjs7lvoJbMxp/qXrNmP1OetJJ/YFCsqTy/YRfhnDYvFdRY
YfwyeuvAu8PQk8pEuTztcdwq6T6f4mSXyBTFVZpNdM0eb1zaybWC7DWKfwKR3B/HU0No7wO3m+aG
9yGL5DLdzVQwl6nXgxJBfh2eAduV5yoM56Pi/DejjjxFR5dR+uW9MQrPI/HuxMA0eFDTL3Z1A/Uw
9ThwZ28uHjmgTYJ+Zm7Yd2UL0rkw+C02XEyhJ1QUSlMaEwnih/rtInxl1ExoK8jtI/B4GkAUDWnH
+ZlxMWQi16qCZLTYa7Lt1nm8tNZ8i516YL3gXv/RhT8qJsemxqm7FjueT53pbo/LVHJVt0M57O+v
F4EL68EEfZhGVQz9D0lKJOKRvbjF9EIT5z54PSCRNmSJ18Nc/kzn6S8zsZ/+drM5o15gDqAZUBRQ
Wz/5gIUf+XL6/1EocA0tp6OIk0flpYpL5yFqEeFtmn5GJ9KirSl/gph9P4Knn19/UsnuyoA0sgeT
gXA1IzbaD7mz1RXFweOofyUI+UQm16AlHuLb31EGCXxNQ+OJLViPeJK7Hb796YNv7tcWGPLKiYYJ
ZryUrSjeQh+L8UWwDAMx+0zW7N2yVTLF7PQcyza6IVQyMMjmW8DAreduy8pAS6qhgAWMadztv1vh
Bz9AZhamN076kzWjSFwXq0w/kLxseQq1SEW39lTpb2/NTABToToaEXXkW1/cQABCgWZ/ZQamubD1
XeqUy8a/CIPJDTvewwBFshfZVXidKzxtIHXbkAL92Nd/Hi90YNihYZ2YMqNgU4ir6BNOIspkDmNM
GEDvhIMUKUpBXTGSw5DO6YzTNBahbAqNaH9OUTxwwBHgYNbJq80dKuP+x9t3fJXI0y6U3EO7BMvd
OJ13XUjSmzSHxl0vUlIQgK7JWu08CmCxoymjuXWK3Mv3zWqsibAdLQ29T3dkE+Q7Wk53AEblaU7y
dodONR8hP7b5upYz9799fylb1LgJQ8vFdWrVKsATL6c3hiC2WML0bkzJUMvhQBDFGO18qqhcKW7E
9aPpLPicP0SOvVAkESvW+mc2rmob/ybOGaSN75ZA6t9VqGad0urKwjrQwENI0eK46e5m4eZj5RS1
+KJS/X0ko8xYPXX9LPcFBuIsGQzucaU/N1agcd/eEjq/mV2U/f8fa+yHvy0fBAz+oRcbGK1K1/Za
9fC3hiEAsXS1QEotHpZjXbDkswTIHy0mJ8CcmJjpVTAV5bTZoLmh/VAblR4aEOwEdArf86pczKBz
+UpI9988wdAq+QumbbN25bgwpuNrToz1QHcaDXh4BEjELqX5OxwbranuiJqfhDXobQW+yWMa8aD1
ZHgaHRfm1McchrVuqxujdvhXfaF571LNj4muw4tEEIdi0U0sLrnuuJ1K6EAg9bLz3h1hzeMQufga
M0kYhyOvQyS9ZZ4DulkQ5aliaXwvxO2oSwU830U93QmcecmAgz9R9YzZRhLIMhH2W8997KE4Lqbc
LiMctbLII29sc5fqNY7ioIG9jUBit1BX0pppKy7A2fzE2uuiOG6A1BrUAS1CVbEjQ+7IyvCYBmrd
fS9gFidrqAAc4hya2I4sKofMFNw6m+HY7ROa+YcU6B5luxFNPvNl8JO1PfYnJcPS4Iqmf5598cEH
fg1qIzCHIba4hutCio0GPF8hwPvrfo9zi/s89BkM5rSaxWeBMWQhQXWCliSlJanF9wuh6iiCMXk0
f5G26zCNCiQiAthqdfteyqvQhmSfRa3GvbB2kU95gJbxfCqXfvJ6CcvUzVafzBkx2+xyc3ZOA4YZ
E/sF+Ky/N8tEdn82A49WorLWzk3MjieFLfpg+BiFEqWL9JGeqO7iz2dxusaa0rl8jEfyZaqNsy4A
OsVhnOeuJJgSPBMFiYHnL8xP0EsBljbxVVDeGZJAB/Eb/Jujl1OAkFa68DaYD9z0z7Px2p4mS2TQ
aPal2zTGPTNL6F4S/E2NS94+aly8sqHq9VVP29KxTusnAKbm89BXVZmkTR3zrqPX8I07i67+HKHe
nAuYyBX4z3kqoFhq72qwHWx3aQ0r3PbiG5uZPrkav8CkYlYARpQ1en32Ypu1nC5stsJgaJAUceXl
da/cr7oJ2bMnBWfMB8qEV09feFZklo3FnMe6I5Z/YQqdYOL5TKAodzJa1ICAD4+zrIW6RHeoWWyO
B13FTodg7swiQIVF9ShMdY6liDf2JPmB23gQOWYfDyIs5RLcxgnC7W3vfbnX7ioAby2FyovTR0nw
GNWpLAQwdJi/2vtS/oCh4CBH/5Kwmax0ODIe6E1UHB20Y8Z6cvrUss0M+yB22cb172i1RQwPhvmS
H0TJlqSH7DZVKW/sdAoCNnDbDg8Govjk+2s06jy4IG/ZV41yp0aKpWucZaN9ZbufA0oPoE1RbmB3
KRgDZK1XoxGyhaBsznNovkFklEK0ajc/XtcE5mpP7zpORXGPYT/kAt5tUtuqnZL1GdqPw8TG3FAS
R6omlOrTSJIuexoV/6O2c428wJBocO6b0XBSvkJCPia40iew3iC/Huc9toGhRAhrj/9le5nO+vWg
2XM0dEB7+wT/v5JqksNIBMwU5XyTb6lAFh+tA+JJZlV7zfg57OQJRNruU+XJxAEY+KYQGfkfREti
Xc3ToJKSr0a6RiuzxHlYcpA/nBzs+0FyISICiw6RJGL2f32y3TeH+VSg7vyhLuhulywvUIGoumAd
RcHvgYaGdyL7koJG1TjGH1hLvbQ1sgLedKMl5U9EoImLerPiCKlz1nI+Nt0yeK0uLKuzFLYNAHEq
M4Z625Cv1lz6NLejAJw5DW25Ju4kvxd9Bt4S9AAPa2/fu3eX74wV30tCQhvDhtMFsQVgNfULNYTM
U0a1hgV0dTNn7UySKDIUYeNsaS9eYm5bvWw126zEA/RPG/n+/XFPrOQJo71tAjNppoOruEkBaYHl
lEtdRERU6XtnA38EX9vt5WLJ9vER/29wyRbhhBT7174r5pMSsXFfvfCuhRB9VvQc2pJ5Mz6QxCQE
IhJntccupOFMjmM12/5xqTwY1RieTzZY3rT406A9IatFvdh2bHUMmWWl4w5LX+xFzdpJltt93QDQ
KxzBeDQXrNDrqmiH9gCvavXJcs/dxPGlBKtjj1CwEJdaWZD2WBKYVp6oArFm2ALHHGl75maUBMaY
PSjx1q25pey3dOElRoXEpDvzPfGZmTNMXRWRZcNl2tq3SoX9L6VNmBd4EnTTkcbvlGOCtQ4Y3cst
uz1lUNFqNWHoqn3wm+uw7fr6YmLHBKK2F+lhjROuCoqU/TrTaZBKWZ3xexy2Ca5ov9Kn1p0tHi0I
S4ZImHeOPuzQUIdW0l8OjEivaPbq4/31mnNH4kteC/VLPrbsSWwi/DLGS1En/g3iN9CAjDnJpXoN
3R8dGsFR9X2zOotphdwumzTf5+GyG3ajAeFUm+vObMA/XlG8++MdsJ36+LVZbqe5mSdFIrQiD6Yr
v+cdoyTpzIESrX5/l86U/07vOX8XQv/3XITYD9/declj0iXmqSbfLsmYOuQH+HhRR76h9GxUT5nG
sqzSZ32fTbN4cmCa3tZOil7zgkfouzkCuiDvxlUf/kSTCzJWeLVop00AHmkqHpgnqC67WiwIW/cK
yWM1Z+yJZTVqz0zLYPIFHwswWKPWZ2zledcRe0aK4YaOzEsxSJXy03gqAHWOp4x/TZhcOgnnM59Y
rgMU0OIddL1u3JiD/dn8CHk+0Mz5rMbrIumdYWQF3JUXcFa06cKxGpRVq3Wax6dsWgeU67Jp0g9I
sdWShbAd+2dQtWsycagTth0kvAcsEkjPiFvKaN5X2LvnluH5HhScGsMCIm3yrnl5ePQpN00Q1Mp9
zNASSsgKoMw2ZNka/S9QHqoLx86Mvyc21nkN6FuD1kSRzXFu5+0VeOzWTOs/tdCtUXT27TT121qk
MB6T6Og9QH990I0KJdEG1zrJ4KjzifBqwP13rt1o9ADqZVEOSrOu+CHZrIhXPhq2E4+KM2svGjEO
Q1g9BQTz/+ZCmQh3GyFNv+bhyH36i7AwtdKKzM6a/MlD/+f9UA+YPUylI8Dv0miIKq33se8gbs5+
Bz7pSx+jJjasROchwLkLNM/nSGVbqUjGtEae2mzUKdoLGVXaHv6/EHESdaHcq6uasPzifIFAhXpr
fKSr+6FwLigpOtDxJjKdXGMIQ6URIkrNfuaHEOsgR1bBWTSpdXeZwLefomLCO7NFBrFUsdaMm05l
0psxNPOf7QQ80WloCt8170fhe4mHLBFVxnpS9TA7tlN5iJaqY7wStgJ9F8T4wogl+W3yB5txCOvK
5MXnIddR1nJ49hP8pLpcpOBKuQQK8e2uoENyoiy2YSZo63ckUFacL3FDnqI/gsyw5AzNEVZazN3I
bVrCdFRnMXeCngKOuG95RZvl0TejuxXEcw0RTrJLSLWPifwyndaBDjuLgrhCOrUR7d3raELboXCH
8FlBmQqAodk55HxDm4JCMRYOzSQaltjLp2OTvIhwaOev4w+a1Kb4Vfsw67RMRm+iXcggI4HUYqRz
vGjZWjlQgUDt3S9zVlHEowImxyhUPD72wsNZNLVDmV5g0DIyolzeWJmaJWKpNkfP4mYUBN88CdP0
6lyzme4zORj9b1yIl8rY0p8SKD1/rILIpZweeoaxEpEKZfuUseL/kwe5oXX8ahdxYRa9htUi1dLh
yMiBg3fd7Z6cacPB+Qr8Rw9QRBj+tuDULN3RmfLw2aOTAizw37jrb3bFNcp7nIj1GabRCcZ5GFZ4
a7qBAtprbyw0nEQIIBuldhCUPOUeRWDfYjhI1xOqXA9B0C56wOMjgoZ59A7xW7ZShM6SRf+IMvKO
EivlIcwbPhSBJxNdlqmtCINyLi2hj1HOBkNsUXqtHPMwWk/UbFQBO+EjWWW28on8hCAmhTNYHnsl
Me4DwCjJXB1OmiScjFOcxE9n3jLETYElTqzoLonpz1Y0AsDF7/NT+S72d9Ym7cIN+jamfYw9WdgP
R+E25MxIsxRTM9uX8zBfF5UlUcbs4KKdJbv6PSKvizgStyfpaKTfOr4LNSQFjDsIMYUfiASAie5S
Fh/waxZouLGoM8QgWcjVp19IPIyXR5Lb2iakn8zcdB38wGYVsE2h5Pf/xZmddk2Y9gUziprpzAyd
1g2aAwSiGgLfe99626Bhi/u1piAwg5CJElMOat7Y8o+ydmoQ838sRFn70j7rss2tTRimNxaFC9RZ
SfbGj3g2AxWlYmUTZCdOuctP6+T7v8dR05kFiF6Po3Y5Kwsoyyu2+74184cjMbUWxxdmMux7IVY2
kLXsznI94d/tBmYmb416rf2B8AdLL+dHHVWTjwPGadjtkbo81NU/2u9XnbHapqH60IJsCC/ng/2H
oCW/3TYUC1uY/UscAUCNcw+JUFn2BIwogIc2XzFw2Pc0RloZBcTIryJuwIWDqgc3WXQZmtZmYIkp
PnfIlUHUt1VEja6RNobiBp63TUCzp77zXXONBizf6BbWieLjaLEcAgdr4Ids08wE4jDJpViPPnae
DOfZAa0DORfLjwTtukrr+SFVhcZxG8TP95pvba7l24MEUgErZQPebkvKisWe+OEq22Md8b6BySHM
jhQM8jtu9xPDxpqFHUXqO/b5DeLTfH33VYpky/B/vdc8pt+41XA2YhR75L/JpOQpHJUGcECnjf1a
K6MJ+wjRIgkObHee7NGi/fs9GXrg/wYT2t56inQpIMqLYz+BB/zt3y+oC37BBjT78MZUBvQZFOry
Gioq15yuidzcKEsnYrvOoiooAiJiuRaezwQ3i0aYnOYqLD+y0QnbqS0pUIfc3UsLVJC1YaUCDNQP
KxgDlu1c2wrWFXvaQz2EaDcwN3XN+1TbJUDDJOQ6HeRY2mvAER9p5lgDqIkFV46n2dl+FI9H9MAE
N28lhF3/AcYI3yrKHlsYlgtVR8PXjb6WFF8cXHvHsALN7PITyNBXz8JXuDwjUTh8B+uTVWL2rc72
zJ/cv2npFmhohVw/aWx6FQLMwZwRKC078LpnpKmszGjqgBHpAQNg+vq4gK+lSKKLKswL06az9Gl1
hJT2FQ/LC/69eg4GKb851AEok69mcbStTkQZi0a0uN7oCSK7NP4UqSGLSPqxka4Yo4TqzNH11e7c
ZtEbQ3JvbScMadUZHhPmEBcUbqBaXYk1ZuFkK35F8yXSjZoWJ+BP9jnz32BvD0RCBL2J/p9/Clu3
VKzL1dR117eF9T4cF+ESRXi0bwOOQ1WQaSHEQWzfs0Ly8NlA6p/CYDACqlh+vvI1Mbrv7686y8yJ
cGnPx0/dCe97Y2oeDGFqhB5NxIm5PJ8rMamThyhsld22xiVFBPUADo2OyVl5TacbWbfPEKymtFZL
ByKlIumNgdIqbMahbwBFIFy9Jz3cxjtAhUdq2HU89o/mfqs9UA0rGSPxhW5RwBLIqtY3WiQHYdTo
+e0HPDf9Mw5oDKYKkDkLNbHFJatJKaRstjPZYjV2DXfNj+aapr6+h0joftLYvRKPRMiWYGSAkbmn
3SamIPvy4qgtMVLZ4K011bHckH0zL9pIt56N/8ihPjJY6ltaqPy3jKkm8mk2qQ9Aq6LlRLLZ/c8c
0RZc3v2uOzifx/1FsKiyjApHHTIM2Te+YuMo4By94NKyq1vZPU9OFQHegKHB2Fn7tZooN1rDMJxJ
+Sws1EsDpYwzUfrb8cpE6BUyCuwuqpeSrGUFkoiApnPcZiykAQadvdJj3lpRSAo5/tVUCsOUlQdP
j/2txPSe3R9yFVyVtkYf70mizdQD4yQeVSBIgg0oLtmfa/pcsq1nE4jZt6m6dIoBC2HD9LKy8bqT
ID2MQmQvKkOf+hvEWnp1xHSnpnhFwyPGs1S9PSSs8riVUAqxlx4VB3POOxOzxA7ToCnSLk7S3UCV
msOXNVI06m7earJb1z4Hjh7g5L4zLabacD4CzUL5a8ci5rGcsBEi6pPNDOVGhm7FkiI3Vkh/e26a
t/ph0XGSABFrXohc8w+zuLvX11dujE7+BxSCGvpSIPeY5jObezQDKF96RMM19Ueyyke99irtc57k
sXAB3cU6TKIVGLAJ+6H37OflZvFPsqisXXeYtawNndm8631qgq/r/tGp4EJ3XwfP57m9WLyZ+App
Iya6X5ViX3PhxhddMU2hGsWWVoHZWXpHYyvpvEKLIm2WnUikakSnNdBa30nbAuZKP1ius3BY7K4H
CWPglG2s9Jwt3sDqFyqWRddUyJ7j+6u99JX/3aHJS+s8mrA7XR6n64IOhGRJ5AoMzaZkEifAoL/J
I5V0mmIEtNidPBJOKA9vzPnxu5/ekhy+dlkxZyz0ixOcVDkJn6ThFHgRdjwX53Rr3laMGvFtr9zr
BekfwP5QrsXLX3K+S6lmjnKZeoxylaqWLiGtw4nteGasedoJnSnRjvfoT/HIHAtPailojHC1/0H4
P+L9bUfE9CIvUfeYaIQlRjQ+ZTugKPwwWFxwYJVuEtWcF3AFcSFl0xHe2iJdrLOtucbUwTtjJ30+
0SdmMAnaJhRb2BFbB2EcUN9sY9BfuWxuzqpaBfesfrlImgb14OJVeVP1MUSvqguBso8a0QrJ+nJo
8TDJIc2eq6pLQc8tWQ+0lf8At0emFXMIFFcoTk5vmzuDc2QmpjzwDt6Lwd1HA6rRLUyEW6sHzMr2
D8JvuLAD9gOjz6ckldvhyaTqAlrDPftvmrfve3xjIAJKvAkMiKVvUKzFZ+4ZZTtXE9cTR8Hkv2vP
Bxr4mr21KfAMx8AgQIAYaVCxIaPppvvuvje3/9KAAFc5jFQ5q2RA8rSnvZLCCy6FKa/8IFCnzbh0
SoXgLwyG6EHuFuBOqKzW6Efph3bTheA6fiSqN7SLZ6AFJlJNd3nR80nUCRBouCA8868EYPfAWlpt
tqHop5RnljcuuYpEJ2Sbx/E4kf4gTrLVipMXGBCwd8vStA8gwJumlYKqVTRVwDWRPtKN3VV0zBfq
nlG7kIGQGpfcO0QLwMnK9tCfBPqak2YhFLe73MOOMBKjsznZmircYA8XCbDUXY5wT+BgcRqMQZrW
GDBxuzQi640kE4RCuxGdObj5P3HtflDR7MjB+lsk+JqqZYVhoUXaDjQsuUXV4oLyIj2cPj9ZB1VM
0DlmcDn3A62pL461tqjZrjVuSgQdexelUnkxu4zG0LlYgXQiZeFN71G9AXDZN7WZtEuRBbvnYqfv
NU3iXE4WJ/bsPe5IcHLPXpzcjpc86kLghXc9OfUqEoS7VPnuUTgHBeyDAxV/8X6a+Wh3CBcQTRqj
sla8sn8uzUOmvY/m7DVyF86LXdEnmXywpgOTypzTIRLJ3Q9aAmnfUSiiBdDhqzzYvVk6Gy2RmpJ9
RY038KQ5nQURQJk8qg9OZUYdTUi7rc+TPZDWDM6vKEMOiFcn0Z+U6seSg4AxpBKbhDqOOr/pOFhF
hEbDmpykRzgjTy+PjlL/DT0QuzS3uJAuOyRsyNLOvc88L7ndNyjlOwApGJdLlej5ZH5jvZ1nNfe7
fdeuG89aP6Jgr7yy0eP/Ie1Zxqj61fw43Wqehh1Mrky9k5bG4tq3xIFpvHS63vtRQqQXPvNN1LrB
9zPNzvqXD46YaBBnu5QlEcYyTBDlPD8QA68xJXbil4mUnCERUXGaCZjM88zpHHRCZXRTs63SDxG0
1wxZaHpXijjxCQJCGsiZRvVKc6hPrCOVobkXzegAN2qBWqr7KQq42m7vxarD5ihhv2yRFIGRTxsC
83J4rRi2/udgrJFCrsj7doggrhcg82IMHUPatXAfFA0fUhPDAtrUdBeF/qMi4q5d1XC5bMfq7SiT
T9nyX+VMwO/slkPpRgn3PshtKVCFYTdjBlM4MM0PXWGE0dVszGrGFNc3USXiiCwSS3uUr6q24rwu
ujGCCAxPcUP4hczIpg1JRNS7cXd7Fb27TSdyjECdA9b6aiEvxeeFB3Y1fyLgA0ry+3hcMwphYEzU
iIrSUzHijlXo2NVPW+U8x60hcg3cih6aGcMnCNStDsKDs5bFGVlqXT4zblHzufvLnJndcoqOv3BZ
HkNzquN7Yaseh4ngNHpublpQBshvWwXWCl5iZqG12LsLLR73d/gbNuJPxRBIRWBhrrjANU24/hcz
mzLawkICZokHPPAqCN0b3xZ1iL4r2jLpUpyUWMvaQGmqFia7WzTkAzgaFemd764KZK5c0U9YBR7B
QK9t4jwDdEsR1v9myghds0L84UwNTKdIDYQoNatVPeABPLDqYbOsWmCZXs0Kgw9U+saWdk1ljpiG
Avid6VNMAFLoVmL26F56ZWN5V6RXnW7i04RsdAJSAJTivKenp2YEADzKfWqD8j1imAQO0DcMdlAH
iIW+Bcv6poxOT0VC/xoSU+bsTZsSlBSzi/XykugSLKFVZWd90Lu0XgUJe8kTBUfRn8mu5xymdhP2
s2oI39gceZPnFjUzhNV9ZD29hEz+y+ZLjkdPBQ2jWctJ4gOcOAT4oyyx3gZX6n6MGg0s9LL5LJNF
3ypvc91Mlr40pivwGueRIdRrwq/3TIuIOSEcocyMpVFlwGkL5jHKJnmk7yD9rmDTNyXWxe80uTg2
e3Kc7nUXrGLrh0fiXSKjkLnPdGmnSpBToOIGLf1XW/4uyZ1pLT5Mi4QRlcG4BOJhFqTmcd907cjT
iObBjx0sgxGLYcEnrX9MNfDmIwwlnco93ReTD8aJVORU9hMEv9GC8pZfMaht2VtAVcge33kIqTaV
4ShtVSQRxW0a7rTERxCgBUtnDf3uLtbebubrlWUoypEfmlLxo4Nk0GsubPOrwznwTJ4smF2qoS+0
+2QeJLseqW7gtU6SCPX/KMhEZkhfn2jmH3+wseL4watafeydB39DbAP0rsa5p18ujm5FOw6MegnJ
LTyU1yGH00pg4rzuVmH+IAKrFTk5MvWdn3zBpACwPRA3MLdgVTmtbbY8F9mpa1E/rjRxBICPJdaO
aFiiSCPKEhuPgB8IimSFyGvu3E/Gc/Xi/5ZChAJ2bBUyVDAqn2bVcFoHTnKWQW+bscaWoRg/NKMn
VqXDfu2yCROBQb877+Y9jngFPr8lD1UzbJYfUK9C+x8OWzSOY+XM9I1isvGrYd/Mle6Gkkrwel9E
iSPWK4DBlXp9ZxZWsHIGI8X6+tkTw1LMKhtYU4aIZmGMl4HXr7Tq3a6jVi6OT4UY2/5n1DEu/Pj8
8YoUellii8OBBfN3lWV0gHbu1zl8+ov0Xay+5QQxMyXGXrFzhlVncqoPqHa7nzN8abE+ke1l8Soe
S2hUDbJ0xlRKYXbDBgXm8yuNZQKkQ6Sm8egh5gwzw2kpLEPD3EGYFXGeiGJzKWXqjiQZdSf1jo8k
ImGtkPEo7W2lwcOwk7SUQQErEpEoTQpb1ZgcAvnxwoz3npbbkwK5WC/X1NE8nSGmyXAi0rK3S6jZ
uF7Hj/sM2Nb66/N1d69L1k24TqhylMVG74jI4/TBu1XcHvFSRCtsujFCHAfx0zcAgThtXdgGh9p5
nNad9HLdmEJpQT/42Z0EYbv4/RnEt/zbGmzFJ5QUmgn7mrQbwQEdGhmQEBjeGu8N098235CyPfp2
6n5VmTMQsEPIMxFtSnPb8i7f/0SFwEazbxzx2uwax8khDB/NCC0WbmE5gIdgA/NUk5xTvdK5Nc/n
SxwMf65kKwl+6cJLgDskjiVAoNku4KT6zB6DZrGj3VVn7jkX4rw1BuMFxS8UY8koIo9qSlfQ2jpX
c6AXPA6owHpwRRX4Q9N2EsyrF4mR7joQH8qA/p/1LC0NV8AB/5yUnNpOYI48qLVJPF24gzhkYIFI
tQ5PPdg9p2hCilOFRrxL97+uh5u6gXu0sG+cx08G5/bKlwKaHPxB9jiZe2IoMmIXUqNytfbZV+Yc
J8O1k2W38g00l5kMc/k6d2qVqir4ZD3xd3twIH/IvTymhDTC23AfR7os6hVbdzikxYyhDogTnqa+
ro9iIVsk47ZlSHH1zEoAKUBGZFW6c6jVvrrJJE3j6aDWVEV1sl6sAAEMceYXDCT7RMZ8psgqIrs6
svtUK0pcP7P6JBNugXiNdGIcdWIpfiEIeXgaTi8vPAbDMnbhfAwKVBX0jfNOADTVNmXf0ZXtU8n+
rAzWaCKGw3hMQq1U5+MnDb4aoXnJ96x3QB8HEjhfoZ7wQphN9zZhWUfFU6ASk3/44rGnPOUZBEJw
2qQYMpIqP972Po/Y2k0q5oE7UnzUjAZR/X2Ukq2lHAp0WH8L00rE7Pj5jEkFONP3ieNgryMRxgbz
QnjBTQWLpVAjwk55bLpRGTWhRosPL3dQXVA5n51Jhy6RJBwrDzpS2Ixw+/JjgX4AvKglfxB/3+HL
eZmmwcPkMPOdLzAf4HGJBznkaJ5CdiXdbRn6pbE2EdDmZKJSroIktBjjzry9+Co4Knu4oLq5NylX
VDDFYKvx6P4WhMNICzrVi2POE86H8HocsciY4dHm3mqZo6OPHTTB0PXaHls4aar3UZexkqzYJ0SC
/KTxP+Uz8OK4ySxHOZtqg0ES+Y+XMgFF++Ou9E5En/o8O+Zz5CmspqzqTVt2v7mVTnzd2msngScz
uMa1h9Uhx+1Rka02wxqBSmzK9GbbwWARxTQTp7dD2jFuw6OmCFudvusoNbv/4M6VZ8ZvODVv/l3t
ejdJ3lNSyUy1LC87uOh+DLKNk9hUKh9Y4W1PuqtoEmuL9U6PeJfKx4Qjmh/MUXqPpggjNIrmKsht
yJtWTdm02KeKdktkrNsFQOs3rEBCZcGPz7b09ZK6lD47glfvLBftutROZpfpOUY3/K9iW2Ir4Xps
D+rNnMI546kW8UgoHzNkdE5bqNUAS6PhCepb9Rvis969Lus8Cf/OrWjELEUchQm4B0yLg/mDFKqX
hAKOATN+uXy71QzpAA5Xd03iANhx6hTHXIYQaffatvjwLJc0X3mZCQmt0caB66t+MsBSfXovNEgb
Ld6nd8gocgK0nQnSKTz/EvlSl8GpQAAmaS7JjFHvRUqWoAtFm8baB+2ECCLo1DYLxG7RJHscmc7C
A5pN9zSNRzFA4gKagLDdb5U8jaknQVb4/7JsC/h6lnagR59OyRJ68/yT3HxpgP4kpLqlngFb2V2V
u4/+fqx7Vd9EmVFdsVxgC2hmHBWbJZN5STwyIKrtUaoV8raaSZRxTywV5N8MXlpm52DIzcIaNQHG
orR/o1G7QYsWthUMypBYO601RS68Buqjroh527b1ZEcco3GdiHocM73PoxCSLYARsClaqOYp8TXf
c0w8iSdXx47LIDoAWm4ny/sk0wO5pMmjZmT/e+UAbA7mu5HGUyL3pwxUIODxnlLOW8ZDzRC6LJH5
did8FQboBRV7V5b9dzLDsFQ1L9689lYs1MO4Wza7koWqt1BVTe+2Mogiv797RubmDSq7yCJmgnA7
J1g5OAexw03tauOOBMaIJrF05EAjdhSs3Q5xGe4qwErSEbcgEVdA3EFl+0/7gmVUuUonFqITdxSl
Pb26fSyn6gwXlxfB/dASWLGtoxlKIo+5VnZ0umcXKPzJuFPHSNv/5OJRvmeMZVBh/2vMwnVQd4YL
qQp8G4Qtjvlw8OxsYEYU3Vw9YxNF3qNXSvZIgG7U683FL6YPi8+qG+68kQUDheyR8cHoE9x7/jo4
kxIMIVYcPy3bw3j0rArFRFt+AJQ1kouCi1zj8kX88i6S9LND4mG8SOmw2NHzoqwqzR/7WZ7vJ6op
LRkFt5XpccJDFQO6TqyyXhUA0J4nj0T9jmhqmW0jZysZWegayMSdG8AP0RfibqC5Pmhi76wJfgF1
PUXezxAdjoJfBrkVTaNXKxb+1BCsVCAZiFsR+3jJ1XxPbP7zuxP9AacJ/LH9EGElwj4EBA48UY+T
sszCBEInspG30LkVHZealoEYzamX23MGLLaaDyow8onyJIaZwUSAHW7I+jSFPr6LRaNSAhfww3zF
lSUijN67p/QnRk/9ZUQSY0aUgb2YORL66qrKVYKz7w+2Yq/WLGWq6DFcbvEAI1J/9cqyR8jqCZ7f
c3IT75xsKGPeCzYIUKy3U3Ee0w0knSVVy4vfYd7HZiFURcaxa3WcwB+r8fGZwES08yQ/8zh00sGX
ctVCvjBTHwZ+VlBXPSV2mmfqinC1M+Fy+HbVnum6Kn7qdZ6A5/lHZqB0UZ1O8kojkxH1tdjpUH62
qN6z6i133R44efcW/7B3+BQ35uIl+jvlOSftz/YNp3ZI2gr/vY65EMLWAL+jThEs78Fb40uPT6vz
gWLm+D4r7h+UBnncqWg0mEg564Ne4NAqQ8KBhAa3ksTuLDHCVzh3OlAbsr4YHY78YpN7xHu/hWAl
IUvE0ppq0i152Hg7vW+MGLCkRTKK2CE5YGUYEn7yG6R4olXbdCwGiiji7dguZwX8v1nc2cxbion7
OwBWsFNXq7SY24KZUjW7ig0bM4ddAwzx87RVFDbJ5fETs/Zer5ztuXFaGaI+4xDD/gQmtc4v11OV
UW9xek/QJWfzl5Y3sv6qXuWoPOiaUhcnhBz1xN4m0jHadCqRaHVRcHjSC1NMrYUBo+Am5QhQrLid
OROjce0UZQMO+JF3YeFeklLbjjQT+EwsH8Mgw+xAqG+WyAS2pD0LAL4/elxL4ysE44WZpLFmS/Of
NpwNBLjyQearW4AY2GJdw138Ti8Jv+N/oT0hZRaeGzykW6pp5GwBKpUXNUX+G//Wmh3Y45fkUaso
KHEKli0S1cBrmzpy0e0uf2TTMpTg8xu4GHeS3vIEV/JURqdBQZmbAIq/L4aJleRcj1MHu/VEjqwC
XrqxImbcp6qfNSHmmbfSzMGnM5wk/y/mO7bjgTxBPQSoMoDtVMTmTJKdEWfufZ3wWrl3z/mIPtwA
55znzZdrCCdmrv+OUgl/17T4HArsjesACxRtSqW3bpYuwRMkqYPAZSfum+HbdzLLe/vpUNG9CNti
PbVg7ozYNjiwboBFGArUTjxS5Xua6CCyRiePmSqqU7KQe1/J0BNGGIJvUHCXmWDGP4aEixCuu0SA
yQENzrwVZIzfewYHEOT18FzSHYkXQEatDpdY/SiqMtq8zwPlqHDju5Gz5FPN1Zd4P8s0Nu4hBbPo
4SR9skgFXnCnB/n4DjZvYfKdWFaqxD6ZVqWcOLUW0kA0I8SOEFXVNWzLZxpBBTBP7xiXJAYJKqSH
x9YJv0bKSOaWp40dEUffD11v1VIsT6ICJkpXAI2TCZFJ1G9/SJ1lX5stw2a8Q/nIujh6QqNFbmYi
bXGa8A+PbEke2OPkkz8uM9eXCW3Z6qIwEIErw11rYuwijw/0hYpNyvLeEwEtUEkH7BE66Jxv4BH2
t0xWttIg0EuxRaJPbpXcPZdUb4LHBwW0s1Ux7MEBRFWh5VIN2i7uufPRQznsPhlchoaP6zBIkrSA
z/zsKhe3f1AVdoHBFFrdFbs+M3fXn/nUInnZzETJkYYi1DL+VoGKyosOZH4FVHSzW1ZnKoCjVP/a
quKpWce5QJ4P7an1iLnjh0/PS8iEKMJ18OEuXX3bKYjk6qNWpkudwBQZ88VACG8qSP89DSIVt+ye
OVJTK+RrVe8PMCQITtEPRU6GFkDLXDWibBVLiRkp49JbuAoyBMTi7hPTxfnlR26j+bpu7llYwig2
bVuoYu0OnX9ulgbTDN/lTTIjz+NKYSf9VXCV4XibzgzSWOAwo+NrWHavnR/CNy/WinTbjLUVfDlk
cacKKl2r7d4N+Xyy7fd/289LA5HYwHpIcsCc+OTIMZ7GpGzGd5fkGN8R486+wdhpesA0ZsL/Wt5D
WpCd7Fj/gByTSXvRgwrk2sTBoUlSKly8YWRmI8+e3MLtUao1UTd0oiQx9GrwgKHFiWSsly76sojn
i7bF+FqF39tM053OHxEAH58VBZRzsAvafs71oTX7T+konV+JAwEnaV/7zevy4s+d5GceuHLTehGc
/93nGtdzcy+KueaCIapbd1P92CfcJnN3rldYBPrZ7R0CEHcoPKy7JKg6bkYNmwp2zT7IIxplxp9N
GDxWANWHFLDsdqD9kDQU8ZUU1WomGThxiC8qO8BXGhfIwFQ3fbXCuxrwiS4GZiXLfQzo0m+hB/b5
+EFrGfEU3GdJHM4yQCjMmb/K+XtcLtPGS+hlJhlRGV5XfBBgH15kn6K3aKDWSDrzlOg7VwhlVDqY
PR4GxLqL8+zJRyp19m/+7R/S1g7TbDAfSTwhom99WofaUoQquVGEVSoLcLh0YL2aUW2GG8pcOH4T
2myuqzBUBhwXxKUtQqd1oldJvcSW/xKLYXp2qGYffoY4gynej2b/G23ETuhePBRB1g/BjRBRzESX
bDT1mrsmtqvpkGgeEVTVB5+GiOkYTzBV+fkaOsScUC67yMA2A6NyyknuVMDrlDf/g+IMzh8Z4ED3
qV6Ilv57WfxjIRYXDyO5AXKQgzY1R3VFDLp25zijXPmYJdiFEYNEPZRlIliMLnnWmXhSs4VtJ6Sg
kq06HHVBl2PkxVfa/eRjDjYXFFk9jebPT8mBPwOV6+KXUoF+0zOrOTeYy/teg4e0OWKtjKosXnj4
xuV2cu7qOOgkZp11VAJgjktyfeKZqMkW6TlcHhsbyzlJf/Zrex/HI90M3/ZwNeAHjZ+8k10nmyec
iG83G5chf/VbpX6F7pUqmRJToAmqPV4kIgmjy6a6uSokB59DKWyyll0C9UDCSwdf37ivCJ7pr23a
9KkMt+rJ+XpYlgiTNuqmpvOGjecO10xExYc8C7Bra8HnLUB3xT1tLX1i1iZ2jgx2K07BI6E7DMpA
KyQ2pLBydBrV4OVD67lFO4lWIluAjzCvATu15QPGCxtGM6YQsYXoKC/4k9aYZ6t8oAjneiJp2dfH
PEUq56lMQN4bhzg/N8jnvfC5H0cL+7I7DwbjArZmLoRILZqScQyjJxNuxMcP7sWB1kpPopf5h6GT
glnfEUY/b3c72aFG/zKWDmZGdJpBbMFznYez5y9MyDQj167jyyNOxIVbUzpj17CREBZ8Q6Yx1ljs
bOhgR6MtSd3tJgQ2Ii/93yIM36m9jOggmnZBNOyFi9yq+L5rr1cZeRhxphbBT1yfcSB6vopuZSYX
dMnfX+AW4/uVHNtl38sNOc0armldB8E3DvcmPwwVR+94og5mVZmJXt3gMuKMFvWWEa3aXwzXOEI0
zXL6gpuiox+eJJ9wOzwvDVigdw03X2u7NVO4cXMtQEWTZwe7ZHu+HQYJqLKopO10rmiNp1qclWpC
hWL6eMIbNdHHyecxMjIvivSYDxI6qEYNVc5J0b5Sitih1Cft2LlO6NtqL4Xwz1XgkzfGvbiaKbJL
DchirIda6Oj44BbTZkwGhRRH2fSZrRnRzVaqhnzhBeFDydd70wTO8lDTEw8wJfDQPpvh2SSOGnU8
cHiHo33jwBulyCwbminwMfZ2WQckgut0QDgr6f+lBv2lIdUOD7EW6O+o969ubQ+to5/nbVKcNHbV
JDJ41XFUc2hk3qB/fQVo0Y9rvnQF/DopolqWDEvy1w53hz6Mh+ZyM7gW/qombcpQWY4sBER6V1yR
NE28GR7brlYFTYgC2coXA34Gr956TyVfa+VRzaqd6xtyYtgfZEx66IVw2z0rdYGreo5VKDn8pc38
PO60zoCGAlBeRntLa5wSjxak5oMzwH1PwOZHkhVsw01M5lHWzfi32VBlETokJiwXxcsdSXF7KWMG
j/OUqG+uObQ0ne+xFOseHazDBCv6jJ2cydWRIvuvA5Utu3uzGUXsA5ezoYxWjz6EirI6Orraynhz
nAYxdw3G4kXQSl5beyUvuNeTyCyFBg2Xgz2Ebe0tg9rcyLBq5WS/l9boHbe/6jDpVoZy2544RFlI
0IxCzvClDKfD0piXQT3wDeHfvqsF7Hq9m9C/QTgigM/6oXXQ2s4ghJPfjmmDFNyIlD840BE6NjxL
uPOLUC6UMc9JEWafS2QTXEvk5pdP+3K23BzMUWvuqKXbldueVhzrfRl8VxWuBJ2MEWvFmtTOJU5W
WBqfPNA2919NJpIZXN/5jYLtOeBrEG/iuVFuZhnJQmcg60jpD/opldZ0bQK6l7+UQUmaDkMDUKMw
0slM0VRi2/y+G7Cdv+5VYOjPSrBFmZH2z1w8mW6aiXHWsrpVbeEECCfK8DZJiwf4EN9svqBU3MIr
mNSVSnx4+MvnJFOaa9FIxgw/nTTE/sACx48tAcGMQil6+AqoBGATUsyzv/8Fim4kEn786VcEW/02
69tTzT/O8ZvCDAeEFeMytJozQBME84Ni87vOO1gDlw2jnpYS0EoEpVqZZT8CpLjSKOHKFITPKr7a
IDfAQnbgrAAZ3/CgXW0gHY0a34G/uJh+MHkHByPtnPuuWMwTZPtzq2AyMy2jT9rRAlBW1r6e9wKI
qKxzlvkw0o+USTa0dOveI01B0dBCH0fjZEbzGh0m1gey1aYhOvEwXRAGzcMKHWXA/dM9Dl8CXcHA
b6x4OIjKcM8IMdXHMNLu4iwXQ5b5gPIRg+lUlH2IGFlt9y4hO/5QzrMKTkdmV4V4Um2o/BLne/05
G901nc2EivSRuO6mJa5cjGuVkHdxr8I8g4/3aptNmmDZ5WOmWtso7TFFGdfVc7n6SPvWvUi0Xtqc
HqfDtPMk0rW4fNwdnctnjWG5dlYqnV0DcexRTe0uJU8MDCFkbLQKKiTxRouvb6joFFkgmzR8oJaB
50tuW0gXMve84479skk5d/WuIvnn+7XHpl8+GckMFz8OFtXiftmSNXvkCWXTl0uT4Sn9JQ/pwlxW
kggfzsuAgvYLCvRuDljwtX9mJ9rg3UbSDBZdtvAzyk4fugkI0r0XqItvfQtBrMq9K96MtF2tF7GW
SLTZy6RzMC1KGLqb5qjfBnU8X9RR8gOuU09OEt4Ftt2HhbrDy6IB8WofUHaZdmoERiucgEPdU27p
N3VErSY7tp5kS9ZJzIxPyDocsIupULtERsQe5+ydA3lsaSb5r/+jCUo/XHN4E+5u7JX7D8ueTS/S
J/IUzA9Q5k6777jCBmCyygwgs2FUdxYOUGhMfT31GlcfbxmgGGQHExLlkBrDKxF7HiTXR9shwuk5
jlq6BKkmkdBVYbYgS4iD5Vltm423AKEsCo7g06JHDtmDbeY74kDrTi5tmq1iwwFNk0fl9feHwBhz
Ged9q8WWg9ihg8+jYpgr54w+frrmnAZS1DGyGT3J6RIFUrd/9Hh6zrCpT8lHxYi6TRCdv/VS3OCL
JWV4qwnmG2rP5J8M+ZVswvRnIQ+xeqsyLS5yS1d+PpvO6JYMbiSbCSfBnkCJTLTadW+9Zd5/9doo
vjJdWXE/pBPr8asfLhAVJwAKvK5jRQVp+ndLsrh/QrLcd474B7Q+4C4yWXKE1XE+v9qQFhe07sRX
72UP7Nfya55DND3NnJ1xeJVAni6pdNSXrEIJeO+0EJc2ojrq7FhUBwqcNzY8wFmknSkW9TWZWx4m
sz/y6M9ov4dy9ttRwIizNEWQ2E4r0gcUT3JcqhwNPgkv2ul/UXsGogR/2/qKDJsPsFX7U/R5ChKI
MXWpOLDuyLrFNqnoLNxshnFfd3+p6L/XMv3EdJKtX3hzzdl/8jVo8tULMJwG3MsqLA1dSANEazsw
blnNT92Hvv9Kh+gICE7lpacKlNcnsbSW1yJ3hyt3GPhOFHcubjNdZZGFcNPI2nJy93dxTgIfj963
KUWt3vifZUJYQrRaCVE6qmJ1KvXlyHm/ILAduBxg6zwsnDgaBfNB4bQffr+FucdjlS/ls8MOngEv
mI6mUIk2sc/7vYN/RN/83oRalVHQDcC4AX1bTLAgPsXPeYaZBJ1qD0DAUerdiAq7flmX4J+Q5Hh3
yCjrJqrWeEwR9yibp0o/XkVHsqLvTdKL7IebWByiWtQbKsupDityH9mzQSREswcKRWBg3RDLI2FN
puc131lyplXyqVhWNAXtFDrlW/ImfxHEkDhdydvXGQ6Kr9aE7Rf6ayAyc9R/S0FnNlqv6WpXpkFq
9ooLAvnSOaKiEc5pZg1nz0yvml+xWinTAS5j4SEnjsTwKP+J9/3Xa3s3zrxYS3PrS5M3yhufAB3I
MywCd4CvXX2Ti4ZdgwLAklu2KSiWP5eJkPXWfhgyYoshv1hIPg9kZyWGu9zXE8JkSs2OR/0FVxxz
2iTGVAaS+lJKBVuCYvvbAKL1IVtHwJXi3PlS7nVOE0Gs+pMmp4OQeD5mhJoAqalRb9v6QnfiuZnf
l1VGS6bpeLoAnJAiRe36WBZL1auFFHlUJCpS4tAMqOyOTzl02RyoaXELTMkY58Cpq24u5xhGTk43
PWu2x5JeUtrsY6Z8OEHdxo/Eptwbb/XfqMLprz4hre+ruqjkxbIsJxtm+MqpEFVFxyki4kg4btV9
FOW+b0HR6QrDqLN2EK8oqU7XRrCCqMurMe8KuwKCKkfXKM5M8k/BpyttCnU5Do3tIdMC1ShkyNKz
JKkGH01fyLtoQYbr3e54HJAb94uRZXZEpmJXzO7SMsfLxs76KxElvk1QRh9faEi8BfKADguVc3bi
q7j4cBw/uLnMkhRXt6yU+aHItjzoc/rA5dbrW0GlCOkUFcCVUH17dJGe+BLMHwZcbLluLxlPU29D
HtiFAEo/BN4+X1Qj0fY4eIR3PsxypisrAM9G5Gp5kEMhgnLzSFGsZV47LxM0lE1LRfFXgYwDyd5y
NwOixsAZQDT1eTOC9Ent4Mi4B3OA45N5C3i4w7ddYWq76K6FxqjwRcEo0HZUGGJ4MODvh2ahs+UF
7PpCizw6vakxxM/Y6g+WGWncHY5/GBUKlE3S8fmnI5r8yi3QIKSXvZeFfwffa8AefacupzWS1D/K
uG+JrEw/LQFIosYJnoX4BqT+oSO3VQL2J2brdDmTKTPPJRN9U1aCGdNuaaH/kJsVMvWPlMfFd20q
IekEZGzKi4/O7fTzeVpCLFcHijIehtAlHwmHC84uskIP5sqxFUPI7F0nIZAfA6ZcK1LpELMadV0m
IQelma8FJ4jNnqR1W4py4LVVeTR+NnG1GCuXJRu2HXFljhyerrSTiN6liluSsgRxTyKRV8ba3EcG
cHf54KSQgH20Bbz8Vh1Otl24t8pCneKNlXCbz9VmTbjdH9O1rrHTpMDQSmJGBDRUD+EZjVypKOkR
piKo4Q6Oy1PWwQzKkWti0HKlzLgCZMSbOq1YRdoT8zJMTciU7pBCN5ejvOkujCuYagFUVOfDMIBr
WK2GR/TPKo5AsRkGml1GLHlajthVjR3XI1uDmlF7/IVCRWjbk2xFDWnHtMIHR1cGcOQVyQAd3ZmA
+dfkFMfxPDm/Ofu3Q1A0SZx/rjTEQw9hHck7F0TWr8S8uQaaljCD9fY/EIWflflzrDEPRvzJx0VR
2myYf50nyygAyfxc9C3GJfBKkLghA0eiAaHq0OfmYD53wu3cVZ/bkiQY9BTb7zICcDoHW124Ajb/
hM5fLet6BJbpD3PPEXaTc0X+Z8JWuYWSs2Rz73UB7tZtviC2U1X/N3KxY6C8wXLq8EhaRoMBmwf7
NgEQRYPZXhc5v7UUZdCNpik7DXOUOdjRW9h0f4h8tZrUihe7fAY7n8LSuoFij/jBaMGXslgX7+i8
kT9hOw9m/Qf7xNtubiIXufc0SMifN4PwHic/jCUZ/2s4h1uc7ObOBdM3AJhlDSHYIPo+sMO4IxtV
/8kYtnWhWHbf7gr0umcfHIphwcBz6CuXW8mxS94g02TSaaBtWpGuyE6OT1YIPbBxKFpCOATan/pg
DKlPB3PSqAj94NoxZZHHx25+UNZnQ7eiKNMOPi4lBw6Gc7vBmEfTTzIpQ2pRZ+9NojDyEKWUb8oI
VocZN5ECQhdSAdzJAHiYRBNny/68cqsZZmAjM5ALyAASbUX5QVOn+bIiJd8YbV66Xry43F4jMh69
xkPpJPYNzJ+k4A8gXVIoN0dQ/8eENSrpuRSEsOsdvkiFIfA4ZEzzgQkmWMQxkJGLt++sqyX+dGud
C4EARN9RStzrgMcgQXxaJo0BDNN+EoTOPBv0t6WJfrJSb6SKmZvMXcr9alt+Zn0JGXIzKatC6MUA
OrX6Vm6QxmgGs+N8ItGfo13QTItIZ4j88Mp/hRMCzVh3BKxK88STidMRvpFEN6Nbqd3IQXFRAz1c
txgqtzMsi1jzElhXVVAHHHmXQe3yw7lAPIwfYKP/PeCY5pocEsiLZ8MYa+kTVlOrF0rE3zz5UeXA
92ls/QsiVerCFrZ0AJiHZRaWSNYdMfFGpihK+ip2WbVggFETei5YJ5dUHeNIkAeqnsYn/55gEkUD
JLIo89JreTGq7uklyxsa4IxAq1glPJWr/kRVmB7pAqHBT9v7MhvQ40FUNFL/xOHb+mQxjjZko+ex
qjroWuK/6b/DfgCFLhuKB8yZCptciFee51ve65/AfmutumDHjmabJZ3wJxESaSbRCJKaRxB3NcbU
cGu04VRmEudyl7lsHFLO1JRJI3AQnUc6c/GHEz1zIqzJCrCm4yYpjK7Zn1ahwOIZLJv4bOFbonON
hKBkWN+ngL/pAnZLSjeZ5qB6J7RNUYoMyg5MggVvOUyco6m5ervSkRWEFQbmsWskozLbr7ydmW+J
da31kZNS0daoNen+INwIRVQ5E2V1v29WDqcIF4/QxhzPdGeVB6ZRpOSF2A57FMEB+60KLht0OoBa
wDYwXRkDIw9uFKMHQNJyQuJYAC+mRs2ed2jnzl1bblwP3JObHgep5s96DeEUk+5G55jmWXPY1hFr
hRZJYEH8Q+skAfHROqeRKbRueI8pW7dyY/3ebHLSrkExkp7rKCfeiQdIfOiTR+aqxITsK/yFNbEU
1N4YCL5rwZHCVjim399iYSZXwR2ApNcyzEShJLyU8foCv/k3JyhggKQK9Y7bcl1MPpjSDSS2tIUU
w/bAvbkWGwMTGg5cWfCzRmRSBc5ZR2x3eQfXvGA8iR3DQW0SoB/dAEGnEMGmHDHxwGO/040SpnRA
OajnQURk1CEOYiysuRuuqqGnfGQnDqdZKW63R+RiUqcjdCQaYC/IDtL7ya7hczYCcY1E6J6hVzKz
fj/O1hbiabM4Ei6gam1LXu69081tLdOxv5yPAbHbVURNSNjvLLpK95XyPwT5/pZLAWtJBQyZveq3
ijw/8syhcBeuxw+2MCYJiYf1uVcG3cXSGOeJkQwm2DcZEm3457pML/GFdijNMPwkKfSfxpScHOnd
cWm/Xtl4OCe6qERrCMw9gOelzPZGAQRYuKQ/WN2cPQ2VZ1ZAMTpELybXGObTK5pFGFAwzGv30PTD
wuYL3A9jy9weL65scctnUBbJWpM3Usm6fcN8+gmaU/i6nku/sCi0NNA51hDXgqysVM4U2aCUa1yC
tT+eMkzzlI4W1ta+xnyMkgSVZRacWiEQlF7jy5UNPk6kytHYGcmWUqlDHuGy08VLvbWfjZQAXiI2
6ceq+5IwJLNSmJshO6kjfvKEQBjZwOGUQP8cZLzHShFQ95Yyq2iiWGF8+V5D75qvwpMe0c2Mqwfw
cIlJ42iH7imlbqH4110porB4drTcVwfGk/x90HngJo2AIvRtA6XA1TOaTX1bAkSevvI3OCvhGi1w
tXfp+H44H6vvf3TX3zhECrrDa7tlQwwpkNHyeJ0HGgweFnzYBNrDowmWGhfXC4/BcydHsrJKvwJ+
pktPF0gIl2szC83DkWEJqOHLjR+tYtyEMIOqvHl0TcvdLQBy5NJklvula4PSPshKuPtalIU9yUaG
edqFiSvtUoft3prQRveo8YK9Q0d9FzS94YI3UEKDeTEiJW1je24blCP0y00/ljqNKwdmWjlPsOoa
4gO2Im3kiEHjc3zsXLMLGumRBjQI6s4TgegCtw5KswRzNyXD8vgWkuSUniIjPOk8BstfBWWanUyG
COVoi82lA2n9cVL3apZHOXkNZkFRISz1FGZvNriaS/jCSDVZB+oQXs1kQx+/GU6SpDsWYVbVmSI7
/U0S19aEBT1IGNTHYzO9Yd/9hW7ubu3Gbv4AVosvAYadsFwCZpygTXJkvi7f94JutlhrMlPAYx0D
QNKOolrhQ+j5l/FUj/CbK38vneCODhdEtxVs3Ce7Y2RgbslPTLgZD9YWqTur02P/nHthq+CXIb8B
rO7H4Alfq9B5s9YQHIAFVUlAbDHAGHW4U8Boc2o8VNYfNUOPe6/+ly6Ba7QxdtjgFVEFmdZrr3GQ
JJhMlb403BXVwpqXYhPBWxyB4s0cqVfqYoXwCjYOAfOMK5WBaJZ8qK7kfxknKyxKDMZssbZ5QtEy
wVswPrTUbti1vxThhCyyFyzggtFOVViiPykWudOrTN6EiteGb9YiKDBez9Oa8SEd7JZskNVNys4Z
3u4uF5wXijnQs97mUewH5INxr0UVMw7fUk3BVa2fDecsNXTSa36GJ9XjOWSJIdF+04oQjmMBvdB9
IX6nhwo8i5jh7krRWxHUsljUpx0TYKYrQsUVPdAogs0BgLkR55uT389BeuygOvXtQAf+cA6vRkgq
Lxwy/zTMcy18sYY44AFfRyPiN8SsuOueHcQTatp2gVGlrvnTYA4hNpRO+KMWdTQMTJhJQi7XQGk6
2nkR6JKNOUstkbEhnypFJvxO0fLzOZTXnyvffXceJApW2Nkl49shzd+//mMOVrkON7qjHRWY435z
8TdKcS4cmo+qwZwMwSTJppUBTzPw9eIaEqGANvcsBQxuDQ3ylRrULKYSkCMz78MdnkCoZ21buk/U
55BRoKdNBAkv7XiK40gt4Bu8iYUWLeVIeBqpnaRcmRvKy2uXuk+rLmC+gB1mqQkI188Pi6UVp60N
h+iM+PYP9STL85rxkOp+B0q6GqVznqYhJvvyOjb2tzYdjbF0QusmRLppbzy6Y/OE7adejPl/2dlH
b7KQGle4rGryNtQOAuphWjuGRX0kvvPKMmf56Zz0NUma3/L1bHLWRThwPJm7CcCNnKDxgEYrkg7E
GGur0aW1136nHhzapXFu5xpcdA8gByPule/2bzMspnyOCxo8+5QNQQ/anWJqm9moQKJ1Gfwo6d6Q
CJ5Fh0lbvHcR0qMnOoyF1e8V91mGdugesLVshwmVtrr25bq7uGg98ypqzgF3E3Qmb4UJFkHI4Oup
UgMGLQ3VZBlnlloHTidv/J5kku+bunz9JIIa8hiUmNUBEiH/f9JX6FfjRZJUqv/n/BHa/QcLVABV
jPBi5VE/gZPMQQa/FyXRXGHF8OWvR3Us5no+Zq4AqEjWdXCOELw7pzV2jToLi1DYjKK2KrcUBbWh
KsQUkX8s/RI0ERpsgkZ6N/56zwl3vm7gnhseeLRRbCQyaMym5G+HxPGQIVgVOPLXvUNyMETTYQ4D
Xt5C6JA5cRRq9K0HZ3wwRlKWtZ89Ztr9FifCZ7M+J6Ul3JnGR7RLiEoepskC/95vWYU17WbxzLA5
x1wO/eB6nUtDjxJen+YeZCNtPg1uVX/X1CrmfjC6SIybQC6trM1IDXfV6tBbdt+axaUqSnyFJXYu
/Auh9yrlCFzGU+3fQzlY/6vi5791CR98RCysYxE/YZfVIzcnPRWCn2vE6Wne7Ht+UnY7p29l56Av
eY9SWWOmG3BESrExgVUXpzb0mBuQTjZLJq/paWHD1FzDHfoA923MQUsuVWJJ74pvD09FCTuBQB9a
c+/EYpSFdxbfxWKrmj4xTjDEJAdOhls2C0arJAGK2I6MawsWBPw0ja3L0cA09noDRz24AG82otPJ
bZedz0KJGNirZaPXvNPJBdGSJUD8NW4ByKr+3XdgSHTsbKvVTpj+OhA5EC4KsEL3nueh0UZVpAn0
AyE6mTEPdwI02D/FjJ7TyEAqOsINd9iuGL63t1zc1vGRFTQ+4nYOavE2PG+zsfDTwqu1KTMigam9
jANALe37bdnoXiJHyN1/tnYnTts5iKbF+ij3fF2IgI9yu0JkKCROVgSf5wUp4WmUauz9lcq9AeK9
FJ5nP1Q6uSYd8S/m9UuET17dRX8u7uFjy5RQT4fUsTD2bSn+HzIZOxeYQlLGZLd6N//mTRRCvb0L
tIDGJzGV+MuRbI6dzFxLaSZzDSdft83IMsSs7ZHi4kVGgoQv+uoBW3hEGmkykGVpTCTnM6DsaLQ7
yJANnRnJRnyuLJPpeDQFMsDNAvRw+PGFje1qDK1BZKLX+XWjPEDLcNFq88eKRpj2tNucl0R8Yhws
LUc+R0iBbxxYcsmkEXdfL51Wph+6XcM6D9/9BxStDMbe5qtEKPzKWLDGX3r5LS95/z860QBU1IyQ
MVz170BokmvCG+5Zkfh97rc3NUOt63zaMKgU5+B2yUiTbXEtuHf2cQNL91IMnelZZyFFwwQoQw82
Q2i3FilQbvw6H2WKOwRSo9Ivn1prXXe8ukvdhxxf22dzkH5dMEwQOrqeku6jxoNoe4X1a2IO8ZFm
FYT3w6Eq4nAjddc3gyP8I7Go3Ensj1MLaIWsBSk3QM1biThqUxVPkTR6KzZDLTxGhVjYczsQnpDP
GlhpXdiKekWHWU1qYKxvyh4KCFd/MIh1/fwJ6LcWEZLDnEwpzKWMAzAOcP8O8Go8FHph1hisUuvK
wfTdWKDi6Q+RgJSaG4KSyFdmQEF2lqoTrZ58BCw8c1ltYFB7M4WRhrbHkclgmavOvn5ps1sqoqR6
wHP7oZ29akuT338vsYgjQu43dkRyuVUjKgxa0kTiptpG7Wip7KtIXOzT2hzMwQtZu07r4w/z8uGe
5bfHRjf+OID37OdVv7vixURQnjHhxoP1WPmD9l26hksGzeBEq8PGrT8df2RuYPWXlcjlnshxGqHy
uy9BidGTUP+Vo//OZA3pHcRiNs2QckzvDGPJnBW6lxVT+mqZ5x+3v4HzEildKZXQQW4wuNoGhmba
+XPQbEyBGN9vqvCjY3mTf406rUdYebvBLxEYxi13cgADfOI4si8oXIhirn6o7kc9Bl2Ap24Ny7SH
alq1Ad2Y4FNredinL+/WK4NLANNaJlqzqv/USQmaXQumoJRgYeA/33h7QGFWExH5qU7s1yo2plk9
9aTJLSsb9B7AdqzcJ5HQfdbFLwCr0jx/gCQ+6RFBC7Pw34CSRkwpKjAATInyyi8NCLW7vfHK+GwL
bxyGpNDZ/2+G/UkugD222klBrL5p8qAfpgOA0/0OHS8rtuwhrEm90xOkNAJoTUPwnpRxJqh6woLy
i4LpoYGoofRSHkmrBuuEnvVZXtcZ1kdNMaFKtIWF046vyEAbMqN6RlSGYEAnAR7fstUqr/l1+S2s
wInvFKaBcuvKBHXu+qGfjvKkbnffEB+czQLxMsMIWFLrEmPrvcDSI6EcKFELd5x1QBQkPJ42aqCc
QuLAQYbjn+hdPHWjsOCsdTXxvd5bnwvJ1iAZuzM/nqfBwhbACjMSmDRJKqZvrehLwrB5ubodEuUj
42V/ttLixVSESDX7fyuFm6TxA4b/4dcSrMwz0FJUbc+ap2NuBVRoYikT2HomIBgP5HOP8bVgAK4t
4N8xgSu6yPSzI67eD1g+4LnFL77viU2ke8IfFphLzZBEOk2dScNLh4F3/6r7UUCEklufzXEqwVyZ
TP0QeWB19OTzhHrIMKlCdXCOfMkxNFPyeEGO4saFFLsd7+KdUgs7Ofekle2uoOzZtfKp8KUAieP5
ciYynX4suMSC04dPJZaiEdBXpJEEET9P7D5pg7tYL6ZiOg5UmEuzjptlZJbN1O97AZxdgl52SSmc
bKXQj/OmyzC9e8NaBsFAQHo3ow5P3J+VZPPSQniNOYkbO0VaX8p3aySCJDh7XQA7YYWRkIzoWeUU
rgiFStLSZ06zGXDPGBDA76fZcnQuv+wmwAReHO5T0H7gGC4RB35O8nfWzLFLLLhQ/ldrVUvxnNli
rJu9aLQUw2rlmw3WWA1gSBNgiwErMSbmwAFSQ+gachY6BBjdnBkzYSrf2UgFi4j/Et1Kf7kFcg/s
SBtZaFJJOgk4Gkz6cB24pWC76zLjwL16pieq7LKwvyYvpLc+MBWJV9E+5WT47jlVnoeqNIPrXL9t
febA95a5NZxcrMuhYsYqyr/ADtX7A16eGmEA4ufkbFhkDL2RWHQOZfCG24M9tY2F+AttPzw/GS7v
4xkMd590u5238OCkaIX3v88+OXiYiIVSf32Cw3nOHMGu+sHvtS6Hqe7RE16LTIhWb5C4aaxmS/eE
TOWhQM2Sr3ze/AhQZ5TUFi8dO27M8gyCXPSV9Mzhb6gffFf29g0IqndAEs7rQtN8zs5h2Ee6unpW
CgKAQlHM126KBIig8XYww6jybWR4MDyKVWGFEdeJfdJp8MNQu/9AWQElVt7Pax7Ls9cqzMlPB2tw
A/jaAX9hUs2ACvzZuyrTpc6XC143kyqb/LzorinAej49T6fmKSrvoWmkg2hYCsIvYHkuByhtNgJW
3/P/mWA4QT4s1xcBN+NmBZZCV51CJiOuqC8AIV8XG7eWfM4WC/ZVszXu31leJVbGHto8XO8EepOw
HVcy23BM/83swf7emHP1ngzSWBCt9G5jnfik35wu8e/tXp6ugn81Fr5ohDDC4thyOAenFDDsK0Mg
bVcH+poKkOJyRxWarVjCXdDOfO4/H2/4UV+eOMk5jXh1bAzg5dINTDtaT7q3H/wTNeXZnk5ZMir8
QQo9+3cnmYwK5lYrV9YgFQrTmDVcG1dNFIil8zmQYFEYFpKCZybEFYQ4V8DP/PbEmYCTlM926tju
ElPhPr6iol0Kc9YEFDNKvRCfCyoDz63Wg+j2saw769NEQ1XF1RMdmS9WSFSPPp038Dt8P9Z4MtUt
n97xVPRB70SM5MslnG+d7xF3aWNa163q342ARdk5EyEyaJTZLndf/Hn7sgzOymvHBFiNyta9Px9e
ZvrHVG3Au0QliUVSVJl/ujGxf2H311WSk+ptyI9Iz3kUV7cXjGHEd/QgtQoPeN2VtTOZdNHvqNRl
A97Vw62JHbarAMoBE6xuMKLc5T05w0YVsbl0jaofm+ZFygRIreaYXh83tv1uv5AUNXHjuOqPkWtu
yisumzmEldUscNJqTj2kTombOs0zqdvRbMHHNnApCCnUDwgs9rKyLE5cBEw3eEVSp5D4uIyu3meQ
7JdK4KPsaGGW/pxPXe3VtqZDUWAusJ185UODzTWMZ/+If8cNjB7NOkkqIXaQrBhccN17rYh1OKg/
Ry73VYan/mvW9RdMKxs7enkmbrDqDbgRg+ayDXgkSdl6ZoM7jpYXfZSt8OEYJ3+r9UCGQ4GesUUt
K+VSDPutq71nvcvV/QiJKqf9rfxiC00+V2uOsb6udKXfk37DA5a+QVzsLKvsdN6aTucElZinc06m
Q2ivq+/fLHRiqRC7BW3M/VYUvNJvyGuy224jNVDIi+XEt6Y+MEebb3pQdTJ6ENDf3+OPijhWUfMc
TiDkWmnAXPegWXwgQU7Onz7V2TJr7fndNPgI+OQmexX12SzdTin7OvZLVE58+lQ26nDaA/e2St2P
DFrRUYeB9nqm7vG+ULh5iMGhI5IBjASolvwv8ls0PR6lONLhkEHemyEykzSk2mLdg5GJFyOIX7uX
7ruXtpuIY8lZRuJtMqmcoQWXAo7YzyqqmaxpZKB4BXmHEqir3XzKwhYJQUUzFP3w217l+JKU67+O
ccSJ5Pc3MOv86c+paQuTWN9/Yjp5RWZDlndKevZh6opRQ1VlK0XsyEwuRoZH4EeaXCj0peJDCPEH
cQRv5T8B2PVDOGd9iEcCFKzPmGfksrLJbaahoIjRk/dqpF9IeVfGy5N0nRaxlC4jlRgzXGQjCCsV
Qy0+iAErBRZ+/9egB5ftV4Mb7EcwZCDz0LgBTRpN//ZVbZxr44MlfKU5a+FPeQ9tVmCkLitPJBTw
okbOCuotAY7EVfdnlqSgSmLMDCw1dwPtbZmjZ5rU2NMfwKQdJlzW8vRxv0OsxPcSQSx2DohS9/+2
UWG19En70mz4CVMOIc1l8dXDB8LOTwCHJWfmtq2TOiuj4JnSlPdZK7nlFH0oiRwmm6SYiSk0tXzv
K7n6CbvmOlGjzeIqQpPUKdfSXybDVLBffZ5AQJxJsDFq0LBKzK6B33OXvnkIQPJM+uBuy98MyS1B
kWCdsBHgjKmy4/uQ4T/AZ/cwq/Xkp7IpQqJ7/iuGS50/tVJnwZdMH1zMseTgoOUe5gZ0qGipuY3Z
iT3ZUEYfrPYOljg/UmaxgOVqnY4rU6wXfzKy59le4sYAl4oeKL20ipeMjdUM6W/SDJKOhjmzAk7m
iPL+yp3ff96CMSBPhFzpLAmRI2I7lOZ2Vupz4EthzHV6GbHKSzl6u2KMte/aBskOKh57ZspEDpcl
HNVLhE9+mDtgK0qHuw1ANutpGkM5odSK1qzkD7r5LNP0bJ6i11IiGJbTqtsLe1ySTVIRdXk95QeO
3ZD3hVNJC2bgdieT4gRf7b31AUH1qaNTIUhaj7uxi8j3hzpIKhE3dx7F44p31b2m4rH4tw/ZwBL/
nrE0PdEC+F3DBJ1X5vP0p0BG33hNgUO0kslRelWKZX8pnZEnOp7J7nMF1CVt4VyZQDTXlSvtAVgl
EuXSVhdCp2z1VtJM/Z4mB1PzyHfopVlHcH6e+Izfx4L0WsoVqcVjfGS5lW/nDd40MMNraSYdHMlZ
ckJNwgdsGY6961r73epn9f1ndI5aUdCFpWYCpnv78MGmbj8cnGo8A90ZYX2h0co33JKCdD56FpBy
meks+Ehj0MwWqNMkZRlBJAnY8mvh1c8xTroQyKxtWK5wJ4TkbNXGEfzWqSB1MiHj1njzOPV9+eZU
jFM+QQ5/ZmylNqlqOnZnJ0Uz5wlmosN9wInY3nCzR6vDjGqi0JvTuqjM2B1Dml04UIwvb1ujiB47
iGpWpJb0f+PWEo9CqUPYhusNolXotuDlLFl/ZqBWIFaD1Py2WETTK3ESB3QidbE4dH+xXuza2vnx
YA7AsbuB69oSRSwv/WeKa9VcNZSNZvu+iiJ3iHGYRvcBE3ZJ8/jkptrtfIUcfqWtMAkHqVbHT+s3
1SthlpH+Nw3Si5QbWJzoHIW8/zF3/RH08b6sMroqzmmwgya67H/27CAmpcF9E2d2KZo1LvKK/VWa
3qcvxmI+6uKikT7ONvbRyARfJY3VNwzWXoR89AUjFTtFa1rcjCTdDGMdPLiaCKk/XzKyN0B7IXzf
cw/AglJ4w3faJ6phMCLW1P7Nc8WUODYeMQE/fwNLxftfWhv+wan5ooG1lqf+zMf7ONtSqMQALNNo
hrNrUIgtQOIedqtNFTXcV/WSkN0+NiKei826HHQ9N0sFZ2ifPT03WQuLO5lJJYq/mYotKryQocO3
lKmSdr72Y7/TGKdjFB1ur8ShhCoBt4igXoWjXWxzfriLXai24zDInIo/iThkoZZFUVN3dP139wUj
8zWRn6AEl1AdiffJ2aEOxPb+Y1PP29b9qTJ9lWfOvMFq1z5akJCVW5cLKgtGnMN6TeHPtt8/S0oW
OooyU34zLC1HZSXMwmiEyyMjtf2jYJxMywakcofTTFSurCMDC5HI8/WYeDU9ppqvCfKJdusvwixi
02eDuzZQKaGNizg/4HOwwHJm9762kAa0qFpqsLBMleGfh98Rhlt8JPsoy/1D7brH45511Bwhbva3
sJpF9ibW4+OMAOuv/QnMpb2nS77qOB9+VnyK3+ssq/sCLA3p+um98MIwwxw5Ckelj/oaqPVWIgim
LH0/3mOyLbnwDqzJQR4lj9d1BNL4Ib3vuuhJNqTBOPpe30bgxMwwi4lgJm146p7cUpmaVXGGS5yl
RT+ZWjrZlFnFtu4DilAIfr9ZnDGhvwfbAMdHH5+h9d8nqRoTsdxBZOgt8cO7+tpgTrO9DXq8P5eU
IZ3jBUHVCNJbjoX21NeibSlhTT9Ca7QJpBo72LvdiAt69nAYx7Bmjvs95RsTmPqXoRrFzsvIUzjy
nAAOFM2zOV9iqtObuCoj5M6BDEAtRYPFvPds3a2ex71YaIH/YTdT7+8TBnl99NU8eE3gIKj83Od1
fPt/Oyyg9j7LHqxq2nYIYCmUkM+oQKcW+T6ftO0kGh6/BI09HNzkmdbWPlrsCj1V46UgXyPsn9DZ
RHkAhZM351ukgtUzVw4+Gp5NV8gEESoqPVkBo5Mpdxa85D0F9tk1bFIIWB9IdP2aK9bxMxi4rPy9
uJAu2bOt9N+HkGsyuljAmqMilQqA1CbR7G5SPx+0YhTRfrK9aB3Fg6eBwF14eOxHlFfQEBP9C4fn
z6PV/8RlxblqxxsZrGlfstNSDEQdvMIxBrfB2jE6mrHP1R2tjHuKrrw79f304jU1PP7kRfHXCJZU
jb6EHmoYe/HqyL2yJhy+NITdXza7qykFH/IAg55P8cZdSvb2YYXhKYRucgCafx2FzVzelHACM2N7
6BhOQmSYIqXc6A80Ilv8oah/wmQ+aOLJIV2dX6svsFia1Q4pjTxl7q/3NOkTQf/JicvM9nhTZOVI
nc7E2CyjrCOrfLmb3KDHYlhKqUa2fkTsa6zgGNlz/atSXsPmbQ/jMKFtk2J7WWtGNeZbN3r2EN7w
bgcQHrqrDDu5BviwoYRtFj/ZNYZ6F3W/K1x1gjyrcwxwCyp/vZOWBjIzuSo1c60EgesW+I4jS55X
TO8rwvmp2MN8fmh1Fy7MQbqfZn1bydcgiCrbSU2MQrHtGKdzTSGB+PBuYJvRZPv3hTezf5YTPv1c
Kj3PjtomAwZHxQUbSnAoWJQFTcgbee9pBASpYif0JOmVN6Isy1OVo9AK8f10XoVNvxQfj4oh1Tn7
r0q29XIdtSkwv4u5dIMC/V+FNy7kG/2yTq6xtrXVWPf3UY6xrCibVIqoqJVM4eFVSMiXPydgCqbG
jvUqzjbhgz5E/cdAbms6Jsil+GmDttLwnF4abpUAYdRh8TBOD7OgpIglvGohB8Szpjw9V/odaLU4
yBNlOlqLhRmdzH0Umb0bI/Mxeie7iON9wv3VrO2RM1F+oUuAAysUUgZvPevDiaUQN39f3qUKyYrK
qI79PRmhFVAi8oQCo/qWfb0qz5ygpWqnmesm5uDbS6WRjV+ZwL9owCt5lELYwqu3DGLewRUPfmd2
hV1TYn2eyjzB4X90eY58T/+FY/FI5KCKCnWcFVIGdPA/NS5nE67ZEy7q6KWuyeTUIDDZk5autiyw
6bhp/SIIyv2OX3HWMSUzCaWCWa+zSOqMg8lvudOj/U5pOg50bqkGXiuzzU5vkG771uLOGIJ1Cwuf
O8KxgbUxwd6xWTQ2yhmWgJsJC0tMLmgRw/IPbcVXEC/ag3Qj7IJNQRVNFJueJgtqHxIOs8a89NQw
SW4NG5vu+3MRZH8y/8sOFaJ9v7O0MFEiQ9E5jIINTNNo8PEhBhtQGYtWmhLjCppVjlr3Z+DSu6m+
t8jHDWlAWEVohbn5Kfsxt6Wo/LCU8LPunMxhv2eGqznLDvY4fZcIRUQEmZ0LTBke18wpsFcOb5Mv
N82Vn8HFaDzp1QCMssIq+NnjbrvOs2QFdBLCuo2NG3Fazy5ptQbqBfEjB7GnDSHot8v6D6iV7DRO
wvutSaw2fBKLQ/o6ZasLBGRT7FTViZn7LAXrenFAkcluhPQuY32YytjT6bfCux/3UnxL2bc61HBC
reqqVcXIxS9kffndFkVvQ4Bn6ekzJhRGGeEGnQ5sdA16CDTv2IQSle6RQHKimWVExaTwZTnFpHdc
lvtdCgcg1i/hauSHuEgb+x+qlnLCPOY4RiRFJuK6hg8R7DEiGbC4MzZZRkxRciAuwZnyDX+qx6+U
/tWwxBJ48TAgjXu3XBg4KRHUG84dwbuSsz3aMbEqbBwjryRhDlMGwMZwDvsXxOIfp2vYVg8uZ3kz
D6bnH9hHufPY6oAJIq9ahnPIEZeEB3qMZ2l4hvdZipCX3xx+dNeJiCNutj2+E2vt6fP7PWn5gs0v
wCAWnXaCQlqT2HvwPfCdBKWyNjwlWfmBlGds1wWJFXVbvKjKTwC47f1/0tAgHr59GUnhwDaFvuRr
qxrz8qSR0kuj8YQmqNwR8WaQKHEV5wSOLyzayLpYHfl/CvT6gjGq7AqTEft97VgOLrKruus0zNg7
9psnCYrXBlZxsaeOLTbNTkFzj2PH9NyhJUIbFersYO6lmMfcCU4M4TfCFcUeRw61BFjTUH8OZ4vX
VTqu7jBBSeewyFtRQ8UAIlhKNvh6HEJ4GfdKw14mgTAE6rHlqeGvLr8wX4d6dPsJMeolspJzGtCV
sDGvfYoQ9AC0YM6urrf1CVaAFDQbZVmNel+fvcGLoWtUotIGZ12A+Mlgm0YGbuM5uPl1aN0cuG84
tIZKZ2b6RXst7RinvEfOF3uXbnT3EbDG011WHlXW/RyGPNZnTX004OqOfDYLwB9MKy5fDYRxk4Nn
+9C5CI5EKNRq/nNwaaOnHo6CUykidCzDsOT6XCqZ1ED7+XqOhrJ5peqHfHPne1CZu9hhmTpSFxNV
wv96UO7c/mBDGP9/0YivbPTh4b96bktum0fqu8/Uyw85CapO1bIG8szHAwaPsg3J28c92j8S89K8
wLCgWwcmclya0VbpYSZWx82NoOEgbnAl7ydzF8qcMo2K95luUxXksIEsoTx2y7LM1uuDgXgsmk1J
mrKkCwqU6Gve0kJwKxCHTjeDGJTJDQrNMqek8PzGIxk21uUacmm6j3jHs89w51KChlZFhRqAimUK
OBPOAKjqS8fJUtqeRiAkS4ITX6T/B+3Ez5/YsRqGngxN/IM1lllCb1aFHEuRCv03ZSUEjUCR68rE
OsgTaolpEFRqsaT+2R5kUhVkYG3cXShy1DjnsW2iob/6XqfQhA9H8sQK9deQwTUD5afFhVD4boW7
eNiIYou+QilvuQPeBz0cp4piNn4zrZqhz2MKHhAsziUhXV+yXZghd62zPNE4l7UyoXPSEssNSEgs
7IZ5M+ZOlEboVtRlIgvCkXGrhrDT//gHfIuVhSaDEKmdQ7lN3e7UumxSTg0JSVDgakm6gezqG2Ms
liNYSQsMP4Fux+RESOqz4hBZ0T61PCFbvpcerSMKAFhpiqiA3ZoPXtpelDRLpDfYrZsYosDV90io
5QgHVN9m/zuluE/VkrgWhqnKgGR9G3mDW0KlvrHMixRpwYgqfYwEJTF2sahF1XJ8O5MRYqS9VtO8
DKOIBY7fs4t2LYkMPGHL0mqdPuCPH2fsIjLv0b2p9vEJI8qKsHKkv8YPF+pdnou6p9+ItZ4uMHME
eVM6JVjabtXP2+SezpifIqjtY1Fo7kWdfGdmq2b9JKL+Y+o30CDzBR6Q1hc4A0M0gODGQ18Q1NEX
2ad5Yl0Tq+lCfZh58HrZf8g1ZkNbRI6twKNrTsc+wzYYIzaW0gVfQ0VvVhd1ZcgROyMQdKuJJJqj
B/ITtD2Ko7ILlrYdGAbthC4nvl+4EPplHvZmyXBnx8krxPPoLnnVah0TzeoJXmLfpNT8a90zamhK
fnrqXGmQGvpZMsZR5OfC8c3vpYcBtOnIOkmRcGgcRf1IvfI8eHOD7MMJd8w2ziCRv9Ekq7ACus7e
I3kGZWrgNvmYKdO36hFNbwY8T527sSFDdy7tnQNNBYp5lySMtA3Gg+bIgqG/2HjYJvemVZwOof2t
TFhBc5JwTByckydo0ac0DamuQ+fO/iz+CUwH066m1rKvQ5jhwLa8lUHtmkuZKPBoGLVOYvnOQ6u/
Rg+dGJ9Pe8Klq6uUr0UFJDpf0iCT1xAb23FiWGeUfGc6266hCTWdvHiUgA48a3zfyPrvQo0cYkKY
9R5RoyV3X1b/cozcSCCDoklJr1KDmS+/OYvGqhfK2/yY6KzSdpVyY3d9dX4JQjohdGAVXRPdp9A6
T5wcN7PD/S9cSTv8r224HaJBIQQrBwIfseFgMRf+aSkR07G7b0NK6kSlbKRoAwX7v0l43r7tw9ZU
Nxi9IsyRz4wyYN2kyqmcxl3Eriv1k893tfzMyo24R0DudqWI9SvCJbYVZMkKmOrjs11lIxXVjHm3
W4U6eb6BawwuGAClOlyrxI1B9CeJyD6sfCszpWSipoIwQo495gEbRrHlGeov/YTnC9q66StLZYlj
1/p7t23b2tBzLynz2wYV0nGylIJ3TFc+4kfYDQh2++/Ueah/swHu8q8REOjdbGrLsmgu9ny0sKX/
Mi4/dVv2M0FUZYEMztSgp39A01uanyklbPvbH8sgy3ySTlGZ6PulwcAx9+fBmH/feJrU3YRR2iQg
iy7fobGQfTfzSJnieEbq7QQL0oN0IwZbd8hUkSOObig5xKlcqaTXiabmQ7QUXEpJGtVCOSxpaFLh
RIUtxDRRJmCiO27OMPb2ihl5VLswWmUuBe3DcQWsu4ietF/HdZrYV9o4J8rBR0XRWi69zqobSEkD
LxhLDUpVxfgm3x3ydZeb8bkmmtwPkFzqJ02xK67rx11wfBAdtZAwbV/IdIWfnBMdMJARUH6gkthI
y/4Nijd0ksFP5HAkmqyRxZrYagoSgg4C2GIDHcitAWop+XEKWydr1bGRwyf4m0qezIoMFSgvNx4d
Xnzwoe5WFS00wgm0hz9KMKCE60AHtjbhFUK/1626jIUwwYTrWU2QoQqqnXF/FzzUKdt+DAU0Z10W
OhUZLhzERKeETVNnkqRpI/vrpj+yoUSNHk59aIflUrmCx3XxMsaRhY3pt0y+Gnel/KlW002Cd4xr
CJh+/JC8QsqVp72zb8zVzIU9zMOg5y8PmnEakAty3VYDCeKOq1iW0elQwQXUZpDObrCkahanOvL5
Y26Akwf4P41xiBMcUfzKtlRdUI6xxes7hR2tt3Ve7NQvxvdRezf73X5Cn2oTJjyR+HWdfxxL9MbV
RE1ZkAPXES53BSoWxGBMtCBlffAkeIOPTYimnD0UYh6Wg8ekHDynurG/eaLZOEAgujdGoAepatxb
dULDX4ZYNX8JQeA0FKayyIsjOVfT1VlG8IgaO/KRRRW7xLwYhtaWCTCq9ybPV+NtUwoovErr8Hmh
3cr79PgAwijiJrr++WTke2OAqkL780f7+ivu2cx1AFk/E8gFpCINOK8QeTpyzznorTiRknXD85/7
/4kK7oTJ6TdMZBrgl5B7csw/y3eDSEQYW36bvNE8wkJJ8Zv9jR/7SZjUhSwIVJfr3zxz1PJQXztV
UOp70cNCv5mCH1AbWrTu/dGKCBRGmGQpAE4H/uIKRqj9ek0G8Pzjf+iATfjVjOKvLYWqC3He+ta9
GSSd0PVxDdKfmjHzsPkYV2qBgA+w3y28723BY5xuaQhyDgBSkQ+2vZeZxEyfEAO11h6CyPKNog+G
nw0bQuvN7ijkhRzpMC70BMBMeTl7RalRhHgK/el3jLKoy8HQV/TkDdcJEXvQCk0yMr/Gwei4Kf7R
qXLebpC97bpOM+dWK8adEx6WSbyh7C+5QkTcFo809EyrziVv6ElHJb5lgXfKG4RCpZo46sCPVfJV
R3Nx/TqD3K4aSISfUxZaGGWMMONGCaQfzikHdnLgqDkmnBNbcGEu8nIAjtXTkxkbAkC1Da2kLhNT
9pZbKsQtnpJHyFnuqRMhzBShX1uhopHCz9To3R9S5bau0lR5p2J1e+gsApX1ArHrr7dnegFU+U5I
prqaCEDTEDpz4Nt/e9/iY/scS9wamPCd239XgkdmDqYruBjJSMF+uX8RcrYmuDu5YbYDjNl8Phcd
ErM1C8FzInmYd5nfcuS2j9IUHwX+kmyVZnD4lT48PMMPbKE84sRwdinX9OgRU4mrBc0cnk/5nsdj
az7slmFngmbEIc3wXMKW1Ca1kIa0a8jBN5ccNdlSvRcvy/ldppJeLRvr5O5jedKihsNBZnCYhpTU
u4suo5pmUrdsPVZNdwjk7Hz5fAidwJrB1SGh5/sLQYwxWfhIOLT/wp3rBKnicktFMBOe5SfyDHce
bhUKfqQyaIN/Z0nl2Eyih2DLkvHwlG6IoUAe3TJvqoJ+njOEvyEpu9VqTT92j4l+ODB/H5XJg7PV
1tye8iIBmgxctOhzpqRrx1i0VVtBtyE7KE4K835sA2TqKsIqhYbKUGndEfYvFjDah3MexkukkDUL
ZEXOjJsAfZ5rpxhJv+ddWgho1ogZn2TA7zkbP+In38U4nVmYBA9IkJQFF1eqAsTf/diJ5J8zlzoa
E60pMBoiTpYp6rf4rcUpD7UKTPI7I+jiM/0ZDX2Ie8YjZoFGaEseV82JU2cyTTOU4AN/3yEzgdFJ
8GG7yqjC2rtL00seeRZT034d98EBqfz+W4ffYaSvuYJ+sYXEXBIe7JKjeUm15aZ/qPlSV4i+UWM+
625JSJnKi63UGuVogCbhzApwYCUPJrTWIoFumJSrSyybwUdpZ5d/JgrV3RRGackE+NLDskfjJeMS
LDkMvPL+STIWNP1W5Hbp3BtSxECiPjgErYAgliYDs1BMV3LbgldTMyw7JQK43idAFi/aMw6Pk45D
uAGiwohCv4Rv7TpF8x6fxbSSUOIeaizzsJPMmSu1A9g1kH8gKfLTZnYXxH0wMZIEnMnWEdIKclIr
Rn9q+naJJPzrcyw8xNMFYsMoJQcwJ13XWTgR/hOx1yQo96itSdaqO/Iu6wDny0pU2V2Aw73cTAfL
gNhT4LOvhfl8do08pkA5aykt4SwLBdECgDek65f3Ta9UNwkESoc0oIO2qCLO5SokJ5Mf3+T8Gmss
UGhig18BUhH0Ob23HoFqNBb4GOjiKAgo6Yd4a3/Zj4FtXVpSWFYvqEiaJztvwkGGGLY8vVVUckBw
eS06WER7oNIhC/tp+pwh3KW1QjSe4j8vFEB7lP/+JwJXIqNPFlhs2zmdAAwhWutX7Ogpa2xKqgcZ
PAAl4AoA+aozMioiFcLG7RPH7CfCHaqdKDNTbJ7C+uPMbL0KOlAqPlqQv/bvbGIhKhPA+yg7Nkql
g8dORJqP/YAY6Hk9P7+vwx8oETEpEuUD4mrZSc8CIN1X9ZbLdTnAUMj1Cv++BWT/0EP8Ci9ss/Mn
a5KYzLZgp52mC8YY2pP6vetGYumjaBm4Jikw2uSG051vQo8C9wc+IxKWX0nn1y13x8l/GvSuGk93
qK3joERP6M/pcer/nO6HmL3gPmQ15CsciH4br2CWd9TRuMRU3y0TkMamqmNXt2cCks8PVjXN5ekz
ADXfZb21/M6xKbPRLgB12UmOaCGN0Mmm1Hg8/M229vT2iGVLF1Nu3s+J6EfMGy/VSu0UfDou0vOX
2DhsDlzDMvuSFL5Xu19OErAbxhzNQQW7jaCUl9Occ1L9IFdrG2eK5YkQfslodGGWoCnth244zpMU
0TpzzDTkuwTbvQppWWYynbHvQLtni6wRynfR2wvXDqTKz6k1tB5mCrk14YNQSz/lsYw13xVZOKiE
ca7B+xGZdD71S/hBU77OiGsLq16qNh83u5OkQ+WQngeCdzvlLFyTkuNPNSJAn7uP2E3O4itpBMvr
kdVSdAYNDx2CWjJd1Abih7RYlJ+FNOoJy47fTRNP1cnxFG54nqmgFVHkcA2uIrR6xaYqt0FDpKo/
CGz8gTUtElL1bkPGn49gPKxsj9NnBx6GMw4alNEbSvHxbFY4x0YYUI5yE9kGXlciukXos5V0TLO2
oXGF2TFkrCMddpFnoelio0ykdKejxIWxXNkqdEDl10QS0jT7N2EWLILsnDURsbL6Y05bzxf7UXjA
hsQmnkrhIcG0ngIyPMFvfpxldo2NUb8kWwStaep03EMNDwBY8JB1rtyp6QgmSzzuLmol0nT1pcIA
ZJ5bNQSxeVSXeHtSgjPG6l3wR86dqliDgAvqf6NqFxgQLIDvjZ+IP76uWrQEG3kVrEu+ibX0tuNI
VpHpc2Sju8V2mM2mfcdS6N7WIpjcLFEeKeR0PepB+QxLw4IesrV/7ixCYxFs2RQggjil7IAD0OyU
WcIhHJTezpjHP6ox0aZF6koevT5HhlUpXuiKn5CgFVehV1w4oqyNAkcrQb45WqhgcjhFMCUFJzh5
4HzniUlE+yJxaidbgSM0BJl3w2k+gxUg0Wv1hmFrxjgSzudwfis1+0gS7VTGsqfZcfOwLUrwplsF
4DyKmOtM8nnknq9PpqEEnId7wYtvOdOc0CSUcrYPSevWNF2ASAHKpTSS5ICToQe3Bct97UvwyOOd
yYqjzJa+/QWgGVdH1/X1QYbcM6k3sasWSKO8uXQpq3tprt224LHNGVq3WIPWbnzgOOzQU4cwAMlE
qWe5e7Cf1knJvHKLeg0H9HwjCZkYn6/HbenqO0itVxWrMm7Baz+vfT3jsR4/siiDXwanMb0ee4CY
U/RIhFh+kqFTM1fIVYE+v9W7WhGISUibZt2Ec7vSwTMmsKvsBqirI1fUxePrTccd6z/XonBB5Elh
2kP1xjYz1wUzocGbhFTAdw/AwdcItqjMeKQB7Ef8gJeoAbeSyNrCqQGdZjBUP7JjCHOQRqua0eoT
u0YdPKwB8oToxz11/QOJGVBxhkwGWeITTWfNhX/pVMybcMDrOYBGfsXMR9x93O+qARmTnEwNmxwx
0jaNtGGOoJCozkVWBTw8TJyXs5KesML9jNcgRGzRvM769wPssK9Oj6hovBi9gV9RlOp2sTN97ksq
4q/i5YGHiGnx2U+IBlmhpOUAYNavcF/CyNPqaO8cyNlP63wRcK1I9jsThOLGwWnSCvyqP7968w0e
/UqmL6kubTZpCnlNYX9mSnb9CtJ8LDTDmxrvBc9Abx8K3lGGlTlloVhsuudeTn9Kbj/DreE3U4w/
e/8FOvjw9valOz/vm4yyiTYrqB5jDvhadhRIRrc2G8/sy0RpTyxIIYetJNkYJsOEf1QTkHj3XLVY
Snb/epZv8HQwQxRW+a0VPCckwdPN2CH6cLVEKJiNM5CGpS5OLnkCEqqvpu6YxagVjc+cCNYoAkT5
9UXekm3fKHWlBS2iDNnBwqRXv0s38qt6Oe82QoReIhdrWN4vkCM5UZJRg2Ys6vRXQBCqOnEZEH2e
j1II46y+Qt9ny/HuxDnrzPOku3bD/bTimcH742TULxvBnGO7KB7x8UjoCBc23Y7+9cX8X7t0Ujtg
OzFQks/A/DwCbFiMY9+7/oUl5btELWqrz9HvLZ3e87w15jybgt6TlSxYawDnDRwgPQnCQC6hirgy
LNeazCdhQvbJDMFydTl2HlLvHY+xceWcZ8yVW5MEwcm/41O6aDheHohyedk56Fmafkiwz5StNI9e
B0fdOSiQaAfyc1244sAWtEJW4ErX2v+eIkTNV92q0eePQdpPLERyNbolzyuJ8uY4JkwUdHpXbytC
gZnwq/pWRg0OUlfRhIDdGcPFZVk1BmbnsF4DYmvGTZFMtrqLZB4Q+KfWE5FNZnBhVIUth+qkN34V
Zekx6w5WxHwxmU7Go1YuPbNaLpkCZNKsHO3pzdIBvwKR+W0WOIMXDQAiHueP8oPhtZtiMxRHzkNw
9O5x5dnuZVF+s9rxEoUDWyP+AaOha7O1wdzpTiJyOl0FS+M6sKTLTOApLtRLer+ReyP6WxifNN9W
TvyZU8kCgKePpxB+sSpfiV5hi1mU4hO+6JEok6baQSq+d4RbKHQz36guLSqWuPTnBf45YXS8rBjw
F6q0rsGWcb3ab03Qtq8k4j9lk/0QGH/j1SCsKGHw/Pg2kpc5t++iT2s6rgG21Ncc7UozpadbjOh7
L7RCWjngk5/4UGkGRTuXpiOvKGVRIYPErSmrKRPH7s9SDDxoSe19HOGV0QDUO6JLW5JRDnbrwR+i
I9HzlhGr7Ey3LFqXULE2vrOH91yQ3/9lnrrNVVf95WeRaVZHCXKa7v3ZBKylUvTb7pkCT/uczcnO
RTu/MEPTdqBrZyKZQf/wBao/2QNi95xmzWQWQ7+58kyDGRUIMP8R0EdKwWV3LUxwdRE5bCB/O7Zk
o3DniiKNf/LefWCg4WMXvBKk9tL49ZR/3EbO/e6AzXRLYBfVVJUcuikhrxOrMwCNW3D/xLObkFfW
ZzQ+VYj07E83qQ8v/oUzlX+oRmUrB7U3M4I9itIdNwA95+l7njjEGF7+jcj99JLxwjYhctkE6vXk
Zu3wzK9g55Tv24CHunbRne6OUFpVGn9y9wohTrZSI8M30JZ6PkBh/kEVdshzfCaLtmR1Tj2YDC54
7WtRbRrIGdlmAUR8AHuQ2Wmk8r5uB03Z93APpOxFmtcmlgTJvn+dmu26lPYCIJVd3Dx6HBCLoUmC
JFibk3SATcZnDmdefdJqvNPVD6MuAiGfNjgfzteelaQFJIbPBOThtDeDZ0RIrtFupDKpyiHfoL5R
r2yAr7oewWXzOtIYZYpAKMLLI195zDyNhk0Nwzgrtui2Zo+eHMTLnezECYKKXZAMhpcsEqs/yOo6
7jU3iJ3n0KE0oIWJA8pbT/cDI4T938nAsAR/2FT/M5UKzV/Izz9o1zZQEbv5pO+caJBxpXf6H6TB
s4rajidJDpQVskROjg9+Y/q0NSZZgcH4/gotEdeaipG683vAhZgMA5wFl+AvgizvK5dyOI9zd5rL
FtZ6uNr3WCOFeIDmCBVzbGecI7h/RYBA4XJcvePguBjgdu5Q/ALEQ/9EIa8tKrklEUsLkqeSsEax
6PFF8ptOAm52+JckZOnloWfa/cpne2rMBXmNgT0iQjkVH8xW8ABlCg9bWxdAHRnuz/h0ziJhuvr5
lG2/GEyj4mjj+q2AEFJbokZGRnSMb2aavtLLqN4cKaB7eXWvunjf3xFf6LR7VlfhZ7ejzrU3iUFx
J+L/BO9Z5RSr988TjDVD1lEhqli/Nuc3X0SAdd8EOHOtQMeHN/czViq8bwczFTcIzKPtKNaJUAK+
77anBgU24rZqMI4x44821f7nO/ql/5vipFJd1YHSGev/UaMwDwW1ztPj6eYYA0xIzMEVRWlXSa8D
UI06pdg4az6Au5M41kyuWn/2NAcZpiH+f9E8cLUYOU3whrxP/oGrHW20qm/A8ynhYncGgIB0x7Ks
R/QcXjCjA5wZSLbBN46039YSEn/iYG7w9DxJdXCC10xdeJ/Pl0GMC239R1z1nxbTWNXa9PQXJu9C
mlec6dDcyvFF3PzIy5UZW11npZCxtDFYDVUEt/G7/fDvRr4gn2vm/GBYmHVoDea1/Lrbx49EEjmJ
kyErsuK50FJIxqrzC2msDUY9uyFIjh4U/Am5x8KYdEj+QRPaZSlogVlFqFw65P2+v0qPkLqzEreO
hqFAV50HUxyninHNdWMPVAC9QyDvVTiy5zLIY7lWjcJFspuz1i+VDjSyoZ/h7cOLThN4RzYSEAsB
4GZc3/BnbGkFdGsa6l3yi9MudagAiJnflvku/1MoJr5tT/vkOOcBvi3elLm1FMSEkeCrYqcEFfFN
bnnKScoSQxfmg5diHLFj25Wof6zs7VNoU8iNUSm/EvEhe7v/+gQnrdBmLGxGt3R9rFv/6ppUPQuk
a6Y/Wr8IVM5RlTo2rTgescvyvPVJurIoerQRf3PdeoBNA+haNPwU6H4cOaoqjSPIAtTrMwnRz3rN
/jiTCGFwyLZa4M9YcQ9JETUNHaEND9p5s32vuhpQ2N1gnZd7K5wuDkMlBzhF0iXlOorgWvXVWMp4
oPZBX51q+rkRCVyU6i7Q82usxvh8oEqYBm7vUq2cJC5qKj/wsq4gcdP6b4QtKlMpUEDoDw/MWE4o
lI063XDYrWamtLUQgzkRC4sy4mot5gsfiio0GyFdhTwc4++VL5NairRVHdLrJYKOtqcSKVRsJBIJ
lJrLu4y3tUKO0ZFuZraD18Z6zloXeZXe0DosOF/knxl25BPQWal0V4LJZu929qO4aKrBJSbGH91c
+tSeC3qXwVMZmSXj71zRmu4ifUZcvEHtGeq/4yFA8w7eN9g1RJQYHiUQCHRUd4S9Z2ti85NXEJB+
j8Dhy0YCGjIWILCUoqn4pKvWSKwcQ4CPGGiuoQeleeZk1l4SNfdD8MFyUXF1j5B6qa2z/+3yF5+t
arLhYC6Tf4k48onBrvYvvco1ozLqm45P+rMatbsoihWcdiRPtbE1B8kxi8ARpx2flJ22HAmjhrf0
5TcqbPVs2rQ3tzgEJ0bgxLnS3YhSrr3a/F/CjqnjmD0rNUTdAGKVRXpdJ9+PeUZLaloTyVZWM6DO
otKchoeBTF1opXw8gsYqFC1mqEt9lV3FkUbbsabFETpFrffQJOp4ebD1+Y5Emhj/D8bYfSBPamUu
MjSqQCD9QjECEwLoeFtocnZeuK7/A0cVQrSl6LdEGB28qWyo1s2k4ad25VPgQqQOxKAHvt8ty/AV
GuwEJEpmh4d40SRcj/GqGZzYRCKg0+MuAth84k6fmOVxMzR9XRzBG9mWlIBsLYq9Q18jp7r6tjyB
pLqXE0KLnNfYP2IhTKx+EHUavdPGxB7mBs1rq961D8znGVfHJRNPvjOGwKzkfG28prWJFmSQTNGP
ou/3IBY2lMW3Cz/cmsR9EwsNMO4d89AB3/UXZhTfp1iB0RpM+fJ8fUvNywrTIMJ9TmSrfEzAsc4X
BElsTHJxVAoTKaiwjmXGLVq9qo6hH8nyYb4cdE5z72v0K8cFzVXEWXJGatvWUIK+MlrHvg86Mq7h
ou2OUjIzs2J94BRq7Rtfm41cro8yWMM2zyuVCL6onnylMA+/gGmG0CMGdDa13+Y2d9P3aY9V7mib
zFY2amvIN2vtEtJS1Cp0fEBDE8hkDvk1P9pqYBO3rGv9JdEDqtDU+hjngzoydR/wB6oKCmwRtfDY
N18yruHp72X1SM4j0LqXVcz/bZmc+L6+HrW3ifhPyktd2mZJOCl3eaYwykYPtxzusMor0Hufv6Pa
UjzyV18neIf7UDdnmP8v8iaFRrlWTGNAJ7c1yV3+m0fIR0lanCY9u8t+1RMT28bi+/Y/SFmQOotr
k+7WRRFsOf+Dlw0SjttlRPkNMcwx1VhfUrOrfrrfVAkT2Ii7Q4h0woHZnDJcYmGbkxQLYwSy5ua4
XU9UZDhW3MinKCIcfS0GhqAKjkXbHJuk6ha67//655UCXZMcw+PcHIIYPNmvynR0fetTT4c96Sve
QpqG2mrtI/QS1v4t1RU28pm9NuzVrvfFJW/azPj1AazgvemAyZhYiEEkmawadytrsZK33VE8RPf5
TuJNHZ19ulHF6za+sSN9037PrN0fHpPZ5aMzaN/1AyXANIZTum3wYV3YKy4MKaYBpYghyhUyIJzs
UkechA6yPM0G/OSTyDwyvv1N7giMPIL8fJPRY1B+X5pTYaqlZCJxKvNojuXw//pzaSp5t3D9U6nE
QBs3OqSHY9MIdj6zp+dV9dZ6VFPP3XVITAjpvz/tXm1DpmVYJQFmo+Xwz8jf+EU9Vgd2/Uq/09Wz
C2czeaX0iXKlSwsw9sJOtzPxsAk9ElCGi+Dohz8bNXV4LfrnV3J/tSkqhYSUD5TOVmC2m4+8Q1nY
w26dX8WJCWGxVC7EAomyiEFROAR94xWOMIU36A2l8m+wUlW+cIwz7RBPCxRzS1nXG8Vj26oPYXuB
UU6fT2kHLr5ogajmMcdpHFLW3fWF4ZtaCPkBRUQCVekQHLYFN9y06XaHbgyxPVXMA/PJBNASlbhL
YNR72zaRUJjm86aCF24Po1y1JczsrLTYNfL7iJOXlWl4sQikCXt+/CiMdQeM6mN94+q7imrj9d4d
sF74w3cfA/G/F/CPSuFCc9z39TMK732Lu5nYpGcwLlg7AWKz6gugKp3HKOEBl4hiwSYoBBoIFuGa
b/zgmSE7e0g+OqnfYQAR38hI+yM/nbrvef8Fzc4s3I6xPJiJB9dWsla+0Q9rN4cRXJn+zabICH1e
4QzkWOvLIJMUtKZJkSrcCbF6p5Te5RZxzvnbaum/dCJuF9XiPBLieKTj2SvZfGvPMV9z0kM/bBoB
CQS+3ITaVZb5iHKE4cy+31kaESMtSy3hJKf9JxbJuEj6p8QO+ebdXUdvo/+BRSUUKpRRcns1HoBd
3FcChTJcnLIzhypvbn7JL78JlQM1/arYorsSQyrO19OTg/3iUReW7EGsupdgqK7ZD5rLXy5/n3qa
1f/Ft14PCgoXNjXjSKpH27GLhCrhsAleB93PnguYxiqxsgJRM8Ty/0Mz+xiMwD/+quVnFo6fWZnV
xLolUvEy+Q+5Zr8l374Z5+nanyUEyu1r1j3XfHsgQdFfDs0U4dwtfEe+2A8ooDE50UM5uhIGoQzi
DYqWzspTZew6keFkfgA5c5slG3GuTa7gWGSvUfda1yIEIgyIEOhmjqilM45E20O6HkSFOK9yVXgP
kBtdCR4Sya3btb5hyvx5DQ6P9DWmGHq/aQ11VKVz0ofbaSn+rW2NUt9ZDU7VrmItWkYo7xIyccHG
PyjMwLVjKGj5tJq9x8ixaEVDEDUtotkS+472ybKWczjXTH3eRaREimZ7sxv3vrZo24+Hm5iQA+3O
psMPb2S89gSmupNCSHSi+J94CZddtJDf6VZyDxmQeMlosxELrswEs5GRo3JcXJNEceSO+yzay9m5
h9gA8oVsgo0Y6cPJL7ptsdfmA1+CTcVyoLLTD4je0VhfYU6fNwiuQIZnqDPdB981QFQDNdAipqHE
J1FAQj+heKK6W2t9NcclcIOemolfeCAGl/rIDwK5uN6MKdrop+kJzxj6/SfiKKUp8uFpKxlYU7OB
zUnBLCIxM39eXikr6Z/Y7/cnO57cAoJ1R7S/dGUcnmnJ3fUAe66JjrCg3JpUPAjdShgLej7GJN0g
bSdUImIeUQzxOvXGjg+tMGDqZAID+CuAYTJq2HdlckPexUPy9Upx8OpQn70A2++TIJgrdExrp+5C
BfpBFR4vfgymsy4rtPd677gy8h700oCpWmifd6lU4WvdGZmQrGeLBbF4qZKC6S9U8qsJmbPtIEn5
eYh+VsGh6XxAic1Q0wYIgWvimzBDGUDSGxoXKomHn+BstsV3qPHEoyJzFG7kI9a5YOpOe0bWw3eN
75X2IItngrPPyFfOk1Nu2htI9e4GF8cggn3Faa/rPEhBNDQR5EbW2guyuzdcXyyqJfADbvH1VhLP
rXPmfOYjHay8QUGNSSEkq+/nyD3kgiCIoiwKRQfjN9OcY9KR4Hsi4yX+dlUvEUSCx7y/jp7e9+bV
2kXyHJ6JdS5LXQB3ssGMLlCbPs6GDGqxdFGimQoSEYweE292Ua9Q6Yj1CE9kCn3IXJZo0uvrbgEf
3Hy40+7jag/W7SmOcrqhbuh6wFZwjvs9v25lERfuOAo4tAwhHLXqdIcl5dSSGuXsqgIOFVEokg4l
MCPPAflppL0lFtfOkE3fN7Y9lwa7ZmrYglNbUfK0VFUJark+yn7fdu6BJBE2/S5Xwe3Ko1nVpnwm
MPTppQ3IyJo2oCmUfhGRr4QNqeO5ZuZm0ZgNrUeK7BzyQ6RizjKvgwuUCoQ8352U5DM5B3RfqJwy
nEtyavTAGukcgt85qCJPpi6jhAQUSjit2OyQp+gFflImAqjIcDNLfDZncubIKti4wBA/xYE7u5hJ
q948zNohYcXg/zssa8uH8iR/5YMDviVQiE3VKbhb9d8lYYQJkF5c6gze3mE+sRnrd6YrJmoALdPu
gMkgcThrJ9j95i3zEUvOWeY/0HSJtlW7vzWpqfTtzIfH50h7lNEHeq1tNhYcUref0lKmuWps3VrA
v0eAecgFYL/u6mxYIFonPYY8w5KQSo6v5ox3fGQNTa77dypqG8Dsg/OD9Up109J2apuJ9crM95J7
YjZSfVVo3181/MulRXpTnnqZh7fhEh6Apj66gFKlzHcCFVQTi5WhFsQTEkhXipmuVGPPqxjrc0T+
Wws2fsF+BWiIiwfhJqvcP8943Ucr0M6abUWW8Y4kC3nQcmtnETSn806mTmE9ZahbUkC34O/nFq+i
wX6GCmMv40orFW6P8ycs8ylVrQJw1Kx2zhG9pVr7J5CfYxH9al6GwBp3HPHAmOCJRd59xl9ZhkJ+
mGDYmHE/q62RWWaF7P5U1oc86Zh9iZolD01lSJ4Sv8LGTv58L7hU8cQ3Boj5kJHkCKW6691ebxNk
dDcykTIic6fDYnKH0EQrwl8AhMR1SMR7NVu/LNUgJR5CqSDJtY1vTdiOYrlaYkSHFnMznRze4piy
Y7xiCk/Nrtjrgau3bVDlhj+Y2oS8vlLE2HOq2sWiGqwdk+2XnyJx4xPQqMQAEdSKeykSAe9dajc5
TFqG2K2cVnqJSxGPg+xDCHkUBGWw5BUIwfgqwTY6hvdLGVEPtZciydPwyvY4llJ4fEVRrcF17ZWt
yQXFeZNfFsllCY+8pe9JOYTA3qCfscg7uIpmDdtLxTtkSzf6IL5HFB6u2JQp4873d83LPWtKT6X+
1y8Fj3k/oPWXnzP2o7Ci09FtV5yTBGYO843igs57Z7P64e4n0glnzqodErAhv160svDuQ50xmZSD
YuFSoUVD35mN8SPtdGah3eIvpYhuhqGnAm1DW20iExCGtTfx2NOldztxa/7ErKeP9mzib1y3rxTD
G+iRCWj9uugcMDc2VhycOFsRfga6WQv06d8vJrLJTQ7S3jbxwVpufHX+Nv2Dh/agQnE5Zdne0pDQ
4xY/31IEvjgZL1mbNHuPPUVV8FVFeWphKw7xrseoJtev6F0CN20WxX2bhIk72gvXAnNnSm5yJQVJ
ghFX4ybH8F9a2YLhSSBf5QcMuO3DO1f29QanNbBgsaSWd/RvSUK0X9ZO3WPpSa23nPylAus7lWKZ
SPHPQlJHjTgf1V1zqzjwaqM6LFAFIXUxizRmR2irf0v6NHOt5brEZIccoWMUFNFQPtD1HTA9nQ2i
yk0iDfYdCj/3dxdnItqA2uRp9HEmW2m9j5A/OEocyY0vZSwNl8e4L23EYO1OX//TPEQSIZvw95Ud
aOm4RwVTQ9vcPOvxdrQCDNL+GqflGM7p3dmLAfBKzn6SyOgMEi3uza1j/gE+N91gEunnzJfRd2cA
BMv+3YbVooR8GeLZ+yqVqASeHPYAPnipSXDZ5NCV9/iHUUW/njE5OrI40oLvXvugyDU8HObPDTex
wcmAzK6tNetVDgPXRsVCHkTpJLHmQzI/U8k/qQuVe5wUKnuobXQgF/tC5Pe5aWl0Im53qmEukWj+
QI+DR8iw3AB/o4mlFuPlLIf2z3w/vS5VmTjZMDVGfoqp2Hfk2Xi3svSA2qzq/HD7puqjXk/0kGb6
nDqYgdByZyrvVxMd+dj+mqUmLGXtmuG/PfFYGS33WDbWD940TyR9m/pkn3JDbchceFNdwJyUBdTi
2ttU4jnFkMckAwnAdjVTeoIV8HnLShHZ4fjq2BxNUIcOa3OXEB+VQ6huF/681q+X0g9yGQ9qQFSV
5MN2rSu6jSn0UF/uKm6IMWkqVlLU3s2LRel9OQy0/mS7D2xkNSMdGzNbbOOT2b3umLskFy3m56w2
xP2fWyBZbeTW1NumQlS2a/wKccfLmRxX/HdL2dwGGSIgBafyTrcOi5HvLC/f87Jkz4ZRXmaQzel+
a9ZkiAJxo1wpyiQxgYFI+HhkZnDS26mSwss1TjuPlvmQxlGKR6124rxY6BW1YzOH/ieK+hok2C+A
kdyN41sTTQ5sxJdqyIBjmM41/vcvLsrk7xYETfjjhZc0/JCFWMr/72uxe0SGjYnrs1XdmIviKRsc
oVwPYtYsTnJaQO6OBGqmP4p6dwIqnpR2pxFKwrnQ9a+ICGOurUflcdPsl70Fstz540JeWse0iNdA
3rqCttKZn560qCLYFaxd8FmueWh4yMQAYaaabMwjS1hCw0pQhjCS7GqJPD+lm+TR2ahhB1yaTI8+
bIXLPw2TBwG+UPpCrnI09b6BCMo2Mi0FjJwZNFE41Qs9F+eDNDhDtbCzq7YjeZ/UAk7OWm69ao88
6MX39K6vAXFC/tVaaTN9p2EjTHejUM7RRHSInz7ScDNnBCDuJ4DNj9BgCgrvwNP5jFLCSREoag2M
VmZXqZZ996tiDTPbcCOs8pWwv+0/9q064do9raoHkJbh2cQ4Cb9QGtvuh2eAfHJyGvV0jk8ClU8y
6dykvVF5XRQorSSAxmUMk0Xgs/0Jd3B7X9GnX9dsWNtWO5TztFl8Yy4oshe4KSSX1VH7mMBJJvZw
34ugk88MlmUq/wpus7Ro7Vc1tBxJ2gAOUubOuczeja7C/QCjlln4H/zH3mOpVSgceRCgnk3ZwLsw
cxHPGhWdgQDFkgQ/Hj77DW4OMZlzAbBS3lVW9Teh4jqptKaR9yTcOLy+bi/tOl+HXAalTLl3DyHl
HUvecOtPgVC8NiCmZLqNp1TH/J6lc0l1dD93/plrpcOG20Gf3jcMDMRCzFjw9GX2JQUdeN0txNqR
BoWDppeiQzTEMZ/csJsiQRWggTvXA+cCTMIaHbOE4+wgP8dfrD9Nl0Or/NZB61SyyPXNpitTYKje
xOnb053MeBi+isiu7EiAuGQIqS0cG1wO4MScXzfFkL77bu0aRVK9z3mswHc+jPTgZvqJlFjz7bmZ
kuC82Xc0CIqvKna0voRzn8ZYk4tYPJleT5261PB87pRqQ6yUqEvwQrMiRMkNSI4bgzkz/7EFF+yn
lBXsAEEuXXZ2PW6htvzJMsqNcYEgp6QLf5w//onDkbdDw7By0tdmp89GhOf8UQBaUG2n0FDLI5Sl
FkemOmFo2ebQwmlr9A0owGodCbxmie9dp2wWWQXLkfw2fFTBdWp+OonpYWaO8Jefr7KtfDhPRZJ2
0ALHjP6ZBKqUYCoBwRBv4K2hJ3YI5FgFuy6tDFYEEBu8VkcFkSTqAwtbAdV/xh7ZI7S1+X0fsIBb
YmzEFwrleOV1lSuBcFTqrSFTxNUO6jYbV7BbOPBtFc1tiJWUlVQOGPfSCvSz4u7CIO+zJrUl/Y07
IPvKRpMMRif2LYVJl9ofwvP85iKwaoImURkZsD+VvOvUhOu/NxJaQY5Rj3ul6AZViKBlfDA2Vngf
x+j5/UWLpJTG7uAnfu3xEynmZfB3fYAfpWzgOpm2WSEYJ7Y3aT9Q7ssgkcB9Txpp+l9Mn1AGhF9X
Kou1pxKzGQCpMDk/viKAJgcf9FsCrMY7yrsB+5bkCx+M83j1DTu8pSzkKHmKJAAb6MnDdjlkICle
L/1OFUPo+UDW4wjXTOixssgJa+SSmZU4jPB3MXyNCMBDmNSYrL1m4bWFqQ/tDU13g7zO6TFezjlf
JzfV5pDLb+iQ0XW6v64th/OFAcLxcC1k2/J30keUeK+18D+TDoRxiyog3Xx5jvR2PcKfMhBrOfC7
+x4hHhtmtftN4qouafGvboIdQDDBz5lrwqLdinTxwZjqhBzpR8yErBiMeYnLNqjVj0cmoFmgDIcF
u7LvZLoVmZJw1OEdnoXYnaNEKO1pzH8v7X1AK2jwEFatx6vGqGVw29SzuEfRGnVMxd+OhUdXyh0z
MjlX1+nTYA42x/Tqd2E9Tm7Pz8TbPEeW6Jc+5vPrt7e103fnDnw6WKFQQbMCIXKHSUnhGakbdFuC
r+ElwZ3rfByhY7cUX2dWQEdrgixGpsrqGqRSG484bpDYnIWEqHKjqNPTrnvnHU/yywZWrUJ8XVIz
5KPP861dgl9N7hY+U2zcbYkng9NUlkhvmc0cvty43HNu15iNj4JsKo51//8HKq8kQgaLD4Leqqyl
/zkaKzmF9jxLPvRlergWQfZCFUMesPI43CGs6MX0dOxCuaVIZArs+ISwbdX6Hv4tPcx0l4yHeuN+
PYRlVmzkk6B0PNCSsSSkCKnHzTuBQVOAwu7PoltjOHtl0AJNEfEv5h1R+w005I20PhkYCp0smiVL
ca+EbbT9+SEfc6u9A+9oWtl5DfojQxQ0GdJ9al/bbE1bp5bolD73u+wPIbJNPLxzZBOMNra2DFGl
eoRWiKhkvkAsy8T/dOnAGgAjruf4MA+a2iUzPK6q8Eou5igdH+VXq1q4cr8wznifeCAlV0D1AKGy
lktymW34IoqcbWhKIM7HpGc51KN3uuR5apr/BR8Qm3cVOXH2PHRAlQ+9uhtpsh+zkvAZ/Dy1dpZ7
oaRG9hKGY5Lg+sGtoONDjx3A60EqvNdUPzmDzqS1HEA8hXsBXDPMvGUHi6r7SI5nrk4T32wwhZL5
67FusFcJzVmGu1ZEQ8SCMCQ1V78TGrd/mM/ZlUZM4HbAEyuJgKn7XYwBQ8ng8PsjRPJidd0zYv26
G6GwsOOSD6rKRBjcYEqRGgCC1SlJ5C6PN+/ZvdAR6heGQz2YvFael7bDB9NxGY4WSU4wt3srGe2q
E86EwO5GyLeFncG5eovcNEXR9R5o6WGJ3qXEV1Ok0XvptbNSpYX9A3iVeSUsUlDzQt5KRztfC3Jm
WggNpcLrcww6sV+S+zl7E2Y1wfCk9Uqf53SzAl+UV8GnCnQ0O3u0FoeW3DZ2XB987sfIIdF7Ed6Q
kTl/gC0tS1KILK7lC+ueDNj8FMREI3Qn14jLtsnG3RZewgO2ByANbrklWowHbjAYyoMxX4RjZ+Fp
q+6ROE7ZDgRiE2kTW8TW8TgPTlS6PMZR7/pn3zckhrh3rk1AggwPDbg6/WXcjYh9F3SYn/F3Ei1s
nbyuYOsgl3J7Helr7dsj1K9yqyaz43vp6NFj095GCu+BrxmK6WHAw5YjQaKW7iiVNOROLKpulfnD
cookRv1W/G1lgHL3y2xRWQ/KlpHqcVKdA5JpJkNZsW4W1eAVXAZ8bVfR1GwIjed9PlZyrejLSk6N
/cPJOr7OeeTXGjqeIvtmmRMVkovbjj9JjUoSQKi6neG2xGOieAxOv0o5Ft0i/8kfdjLnZ/0ShU2y
TTTQwwOVhMjypmTlCmFxhjwRkN/6yXXr+IftJbOH4pOsAXgfc0xuscMzPRPtmYA8CmwwIG/2vZHm
IJl+pAGkiRewB3Pj66S1QzoT1yJl6bgAW3X/X0SFuXqGj0wj08T1QR32M7vovANP3e2eCA2BQ1u4
awD1L6aYB3RDl8Su2vxm35GPZUHYoNRzGYw4o+qjMUbF31m+XsWzEMaEL+30ACS0LTSa5pjcp8pD
BN7F7QFbkGfQWXZKMlfdvroRiHSQ3Y3g9K4MVromCWt2lspPwjKUYi3AgQBNG6fF4C4g2jenGaRg
e6kC3HP4eT2n/hIDsE4TrvjihWWm0DyX56eE3zXuwSKVA6qNPxBqL9aPwyS7y5PetZtnAuUu9VXS
xTHJHEey29mnF8RQx2NQAWdqHm70rbcgO+otUyvCdtk1vwORcjoEpcoMDXtNhYYTiaSEr5or2hlq
VhalFadxtMf/fcKejIf+/a2rB4uGLMNZgi4nUZc5Ryh3UKyEPRzBOs771avbTPr4b86F14H8eGdp
6yNJVrNPP/IV4roQTP7Jzi6XvmJq84A0qHiWwlox9UCV65HA4XYV6U7r5qBdnzpBf93rMGJ8O47V
yJuYWcAdzS6P4sK5Viqjj2w+bIdTggcxpAUv2ZfTfASDFYgOxQ9Gjsiv+1fiLSJwBL9mNEqPB7vy
NZf7yxBeoubhD/rxHrWj/USCKPAvJs+cxfWkcEfNOMXFyT4kI1FQSCRdhL89XJMZ2Q75wvS9xdoq
IRQe1reUFsD54vYCf9oO0Z0TkWW3VB8EgOdTQO94n25CUZqRIvv1Df3ekcsJuGw1PVsSfx9kRD2n
eySQ1T7cJPkp0CgS1nWq7DVYW1zEdAuRirb64vd/fHonSEzYjAAYwawC3vnSpSeyMFnIpZSt4UL3
dWndQ0qrFqzarCyCpbrSONmIgnzed9E662aRF2j9Fbx1Q5GTh83jrdhDsdKu1CyvZPO7kNXlyvis
OomihPvHMuVcbhwWwiqP0Sye/AeasFPmHwtp9JB/kENdHEw8rQzLm3lEexi+xPPKuVmwN5EglBFN
eMyPV0X8YMyzB3O6GUrsxS5t2rze9ToSlUpSRLqxZm40pw5NhMZraakwgLEgM81RanhNwMTbQY3K
CcpeaDrbiipRCEGvJcf4MsXPSQbSYo9vbnEELYjrKpVazWRycZwdRDbXGdRwUbbsmCn3bpiHgLCi
m2m/QlkqOjutF3xf7t3MFBLaYb11k6bvojTl/DjlXWM/cZn0BlHCSdg5vN+voXhcY8ZmMj7BRvOc
ZfY+18Z/CTrkPYA+A+59NS3N5gQ0Bkaf2GexIbvtGTHpMri2PSppF8z9kFOIZO3If8h+USA1EkGl
HQOPOG+UCdRV6f6rYZuX0OgniuVB/d/4iLYjm3r+2avfYK3HUVEA7tPo/i8dixDjjjJdVjPtb03V
FX2qEIlSbHcFuH3aFpjnrqocl55UiAe0NM/Bll+a5g8VOkgYVjTNY1s0aoPHKh1bcBrw//FhIUFS
MSGDLHpq85JaZ7I56uttMf4ERHA8+7saV1nq76fV4I8/XPNRqth48Deiq5Ey9vaIvFwzRygzF1Fu
cShTPGHue0g44d1FrGlmw/a8T2qXQ79PoKTZRQC66lbMNW3PNgSRuuB7aHIlt+X/YRqDxOS4oeiI
zKW6AGhWvGABl8MnRHY5CI6zw4yifGtBWpJhIvPTEteXmkDgwyD/8EdCCtPSgF1dSqc0xuvsb70K
dpIX+Nuos0JpZ+hQqm6LUnZCqgjo94eCHO00usHqx5HcJEEQKknAIyY9L9prkskumFmhf4Je4Abu
Y5Is3yj9Ua7uwVZ836mTxbPBZFwN7FgRldoHX9dqEXpXi960JIGECbfRM9d0cjue8HZhyesUsCfP
pKAoxSiDgT+q5Smg61Zm8RztXbypHyqXL/mQgq/VbDs8UNdreFfDUATt0gQsS9pKpbxx+RiuyvPU
ToLceow9Tfx6WthqHZlVgi8vb1JK1JirbLGyQxAy8F8KxRzhqKuhbBNACE9MK6pK4ytFh/vgiRak
IhRin5hBLu5Q5Br46RYec3SnhtUnNg1mr6dT3blQ/BQytmoOjDUCgB1CRVpDOa3xidl6JLPlhn+w
ZKeRukC5J8sWngJHiH8mKisidhQV41SF5ahcH3q2VNXNoUMQ98IZTexWlC+1X8utemW44HI0nk7s
pHshxKdHLRCGK+rbrFjqT1GsTTB0E5ViApUwgzO9DcRWv9ZzbgKS8WokKuo6VP/8YL16zy6D3v6h
mF6d8mHNvPmqmyYnLgeF+vy7DLBDEvvBhBLmc823ku1FTBHD4/dqqyKRq4ueFomhQyg9SZXljpyB
gFMHnCbv9b8kUeMpd+tFjit0IBlXpd7YhFaB/5qcEGDxyMVpd+Iz9fRsqGh5xeYFgDixA4CqjHte
OXjftKeppRrXRP2pklmduE8y7Msnmta0oQD4nwl5QsonP4UFkOs37O8jUjt+2RuXmjcas2VIK7nn
puebP8itYCAMH4S1yBNI+dSUHFA4aA049QyDO46azoCA5/wfaE+oOk6fPSGIP6fQfzINTlmKdnON
REix73kqRogpF06SqM4R17dksj1vBxVIlmstinxNMRqrou6NXoQ/CfEiGRAF9BgrVtFOzGAPauaP
En9UCniI7HY9/qLNfZMjhl4gnW/r9iDqOl4qBaSMXW0t+GDDGVJjQLBcBvEvFsoHYVj/TvvKipbs
Tl0VXM4cgkSckF53DyG2TQ3GazzflzmotWR6x77H5Q22QD/jlXFp1pQe5E6U7OQblPAVTr0i6njF
fo2ZETHFxIPSFhcw/MocKLAmeh4TrqZow1LusBOqsYlq8LNUaYAC0Nu0210PE1m+hlGKvHDYCIrC
B5bFEsftzFkbEGAGzM4xS04UR5dGZ7kkaFRNKfD/nHiRKO/F6KGVY0W7TCzMBXLm82n0ixO3opCS
JlhwhWfuX8xHZZAUCBIJpL6lVrM3Brs8DKm+8RW135tVsEaq4Mxx+OmHboUdV3xz3QaSzMGE+3yp
YVKZ7GMm0BaIQ5BWizBjqT6RZg2sbRP1BDkin07JXVCZqYa+CL6Qg4vjTM6GSO8RiWvZQTfNnpJN
jYj5eDm17dLYbA35ZWDzEk8OKzkycD8+jSqsG6xycO1Ie8uXMgzIXr/ER63M6me7m5pmN07CVYCx
kwXxUwoZM/U6cMFo58wNypv/RBmv6xecLJ3yWXYuiOSMiXztaNXR5Bwp1jeKKeN9SVIPPDptO9nX
QHRT5Wt791PwMOnBZklWvb7Oxsmrit6gBC1JtDJrIZve5zeWYNRHwSQQUGOiiWiahcgCA5Cb9v/b
hNwM+QQq4FHOu6I8Itw8yHzTVmEeOj5N+uIdrrNsoWUUwJso+Y0l/tzu6tEv3XExbfQGNnC6ggCn
KWIr0yMn3QjkXZxLk81pZs4zK4KhiV42UFvTZLyL7RztkVELLfGSZ4l37P/XpQTlBOVYTjxE0HlF
/L/SgEe4KQZYMeDq42grjrMxWD6a8VjjOriHt0rK9H9UxsXjCS4tOef5NSGNczZfsesD3Os63iC6
U5IpXIJavGJq5bOEG/S46OcVQau9dVxGxL6o1JK176GV8DrRNnEgomfXoudqEXs3BhY/dLvkpv4W
JGb+LB3nxLU4FUJrOcPbCBXnxcXeFXXC9G2aw8gVoqwV7xY1/utgCWqAZd5L7YqWU+gYrnXdpG8P
W6xwiLY7Y8NUyT9uauMs4CZkW47/azRD+CPyKL566scM3X2P+BmRBO6RhMlkueMXxrotWBiQDZpF
kVOLkYT+Xv2tEbsxuB4XfrZS1LE1zdRq+HsPh4Fc4zxBP2+fw5PPDVYsA6sXP7bkjywq+8Y8lk9K
s5q1ZpSHABnnhroUve+brGV6DdAB8OZth4tXTafeymca5j45Fgyx592sVfPqu6SohWXbJSI/CtmT
KtC6sBckI5LGo/OC15K75uOM7m0l2TM3UZS93hUXFxPUYSyJAjoMevv5QXDWPK+oyIgjIznTZfoq
nwJvG0WU/k3ojRk5xa9yknyQVs3PJzEOGGtsHEhuY32Wrps6civ434VcjvWgU0MZtLX4roB2kIOQ
wrjg45eSlegoadFhBVDSKYKLAn9V1rByi26YBNGNeYUjsP7tgz3SUt3UQNWOjbFitltLVOdvx3vi
zyt0JXvJFTv6Sq5DgQj1vw5KGi1+zCvqxSgdRWPfwimaDLFrCaeoe2JTQlKwz+yT8wbDdXBtKqsK
5EkjWJlBEUlDgeBVWiwNkeiV0x/96I9/L5KcyuPzhp20dSR2s3bgQUhPZ0npK/SK7Bz5TSVX3dhT
y0bsplGn+vahKXKz+iD13UY5mqhgiyMpiu40CDkOlAzH9zZ34FQ+j+i4EnuoqEkbbivvb+SqG7j8
bzEs30Z3SN7M7nQE/IrcXa/0j0VY/M2lbY6GfR/z9AHhTBzJ1jZH6ymCLeUPy/bVxEp5otum2t7E
ES0bRVXYbcPT2FR2qUREiqtlpvIRq9KV+FewznX9bE7JdbV5IjaLHJUnHMrPtv11pyK8+PONQbAx
huGP1xok2E4NFWIdYUDKK9/8dDI8bh1AlqOpISkL3fiwNKjtO2naNWZRokcshwoEBzRSRNZaJnXF
rr9XVLK07Y/cMbAzIQPBHvDxl7QiYl2K7i4wK/be9h18Q18QAMwljEUPGNy0gLXhQrk/5kRfKY5u
Ss9fBGPznauRCb4x2XDYTLtdX/JVRhW+MQNT7XRrTJGVzD3QaBSr+Mbet/ObI6PoYPjw4n4oi4Li
yUzvDa4KivqL7eXyoHfwXDo2QBXzX+uAyalx6MeNMiaMyBIazRdUd3BM8ts5fce12N5wTKvFMv7R
Hoi3GQRSdz7ME7j+1mfuQwsgAkqgG9F9EmK29VaWVfhAFyy3VEO/0DjVqDRvpBuKnT98UGTcmtX9
N9z1AcbdaIYX5NRp5awk9KD6w6bwdY38L1Zrhx9V7GwgOEkh+OT+AQddEJY9VcDj2QRAOQyeHiA4
I9mJefIyrET/GjyfUFKnl7fPm19rY7rS+lx3YxVKSWjgrQogpElorRAbsuQNVQkANaxccYyRbeaC
OM5poAEBPfHShyczt5zOvQPStz+jJKnTUpcm8O4mCPh4lzptqe6cRpZB+CPWT4V8gnU1g9GFutsb
NR3Ooy3btyIpUosdrL9k43jUR93JjFIm94Bkj8o5HMfmTdv/qg3iWqWlXLW2GNDCYk2e4sBm2r5j
IDo2FsVjataiuT1Z3+ehzUqgQG3WfXq4CT/Hd+ICeqfHxUvm4OWlLGZaosdYvKGnDAwano36JYbF
fMlG1xju6YE0lgvfKd7e2W6wW4n6PaYKKPFrZHfavKUwFZWStEQ2gZek71NyPLG/kYyDFbVDA9RQ
uoQR0kO6ENP+d2jiOGILOyIfXEPBHdr66PyCN8aLt92giyO6Z6B5zfyvOGmSPl7tYm2ZwedAdrPD
AMHMNKc2y3AG3L6OoDRgoGz7qbSfw/OCg3gcYuL1DCj8HIYEdgfj2pueRchRw/RLz/qrV3dzfy/L
TgsAvNYgj8AFZk3g9xBw7N1fxRg8rxyQ7V2s+UfRZo1qTBETQSyfT0LLGGCFOLwoA9ea2MU82LTC
F62WvEll9HV4dJ/i2TW1UZGVzm4oN5Q+KflNUsr1l68tPVzNIVcx9R35ZRVqc/y5rlpQIYZ2sgRp
J/CuLIcfYUidZy4tp33bf5sbA4AAc5UhHq0hHYg7kJMzEk5n8qyK8rI9v/CWIeS5ipqxkj+B6doL
QNGWMdbuVIN6dp66WlbI+AxekJhWmbSJrhMXBYb+on4be0J+CYhzLlD1sibPRhVXFEvktH+Az9Jw
A6/EXl/WVVs4BCl2RKP3eTrYPE+pWBZEyfkd3ujXAq7296MyCEiljowGixRT6QLgZfcThVwEGqOG
x8m2GGg7N6+60Ka/XAkBXvNlk/aRRYilh/3w0geYCfaM9LRsCYbzzTl6M3MCERFnNaPQM+z2JE7B
WrTkFTmdIZeB3lrhgm9uIU2D4bgMwzMngnPpQf+mxAHafCC77OiuoN2Xvt2BSZnld7la3vms+SZM
rW/q9QfRE5/LORWcNiISmefBHJy1FcdRkzE2UlpehCoJmdqmI1a5ngw+tusbRbYaTRtb7L+lrVHW
bLPDQmFR9NkIwe4hqEnB7gsCfTf1PqzTW48CVkI8F12FaZH3coHXp9eoPNjM+yLcvyYsispQamMq
AX9pNFgF+xotC7JvacjN9G554F2Uw+lDQy+dpBqKHVYkQcMSmTGWp0PcN7Oa30fALc88VH1ndqmg
TYw0CsRW35Xj/ZDTExT/4aCRfXJeXdgDyeRoAzF0sRXOWAmPjWeWtXBpUmzsepzEufDh4XvyBh7l
p3UpFJtCRtr7IkYAJeAOggxWvqN0qvdu+htSdQsfcM9+DYCYFXyENuCNoa9YDlZYR9emtoOyPYiJ
auecmo9V50xYH8+fTURs1Cwudul5pH1oO4EML1M6vPZj9wxoUaIn75uEBYBgP9BlVxFa3Ao37q86
zHgmpEewR402u80b4l4ZtpuhrNK0Nfu0qVrP144o+lBxN/bXLxs02WTygzfxa/CiHIUgJ/yWtAE2
Wmp2Wd1i1FJXFTnyQcRwBWJIYCFKkXHMu0dCq584VWh9A0sPn5WPxVzsZQlCR9x7ThZlaVyFlTJ1
ut9sVaZuMKnzj++GlNOfQQn1GVPngs+N2Mfu21XqhbCiYKm5wpbK1b5sN6oD9o0rLJSjmPvtWI2z
Egu8JM/LbBt18bZC1QlLcVxekPmKvvTNMCPZKgNYiI8lNzmb9mjQk4ZLTMplF9qmlWDQDNseKv57
SotP0ikL5ktvlRGedb2zFB/4K6bjHeyhQUlWWqIwwWVvsaPEHNdTUeCXwbOPBE7eY+tugfgNw1i5
yr8hNCw0O3xQzSaskuP7DDXfQiP8wzIZfOGlNr1AIC4oTjDGjFqqdxbLN49kk9Mr6KpJD9J8aDYn
wNVgbIKnzBxnxi0uEQhivC9/FdFJNFh2mwvfXGvD88Yi1WkBfwKIpAcRm+HESip3Pie+1IsYNXtU
bfzJLni211VAPyU8K94cdveoJEaQpN7rtsNJrTKtAh1wGxT/mdXH3ms/25M1+zfwU4ZNb2/63Ubc
rCIOq9W45o2N/cDHzJVK4QTL00xM2M3VXi+ZLYsW/67rNlrnC8OQf44jlAyMiTPSYkjRHK6n/+I+
ozzErjgJOLdD8pSe0v/GNURY0Q/YdUvyvyu9asXejIWUUdMNHJW00MphDpHT1bXAr0NqbyrRb/HL
Al3r1cct99MO2QGc6lH1Xq+4S3ZEREoJ7Acepds9tKLwL9ktiz+OTD8X3VMkiYTI0SzovQM2yTPb
9Cyj2I1JDT3SQoaYatHXB5xHkprDhhScOwEG+cdTgqAeCUz7zc2/U+WBQ3vlozwwGsIdG8khW4x7
VdWZpoLzWGhZOq4xu5dUXlgq8zfB9rtJj+qcfP3Mnli0QzF0GiX/iA+XOi6RR5M5OJxor1CFaqC3
wXVh8vmjeOmPhFon2eMTa/AC6sgZzJKLPx9ozr/tO6UQpAXQudLE+47WJjrn4NxVxnrQp7PpbIuZ
UyvcQgPyr/SuDqdbniSVL94ZfHVNmaHm+KjBKY3XNicrPpQHvggj6Vpen6rt0WXL7UN9bjo2EZsB
5LIYoq0N88xDLSLyJGfazmRwizT5Nt6yer+ko9uhdqUY20n2YqBjurW+klnUBCPwP2n7LoDXVM16
c5ljCpKILW/8NEr2egskbzmYBIGkvgVcU1uovwmx8cWfRjVED04YGTfQhQYsb+Uk0fWjUEDIfdmK
DC5zY47+Jf90pHatio5pQpmzz8z8X0PGnEX8FBpMlwv7ZDeBRxxg/sdOvFvkGRvqs9nBNbsnbWRC
9Nwn6TJ1p7Pj/jMrchwxw9hZyT9cXkQdmd9AhPHM0NxvmLbYHBiqiIIrygC97EgEQjK4v6Ay13Qi
WBauRdiLpOtytPuDHvNVU7lV1fcJ5VS0HllXza0rX/WXFCVibdHru9GvBv282Z+nRaEJGnd1LW0e
qGmpPQZH7Dndtdde/WyxfQj1VMvO8gpz54nBpNNuy9piS3653h62xEBBHDr/haqSKCEyYw7QDVm/
Q0KvoVit18ewQrBnfBxIZCfdc0RS7hSijKoO0sqCkkGACWolhqz105eRazHfQ+MV6tjowSB+GSG7
922BAKc+y2TKXe1PcUx0fjAc5rQQgO2fqa2/wYVEwdTtfYA1AViXoRRssoI56auOysUSSJE1croz
ATKT2foy8O4fu8MLvd8hafXJ+e0OhZGfrb+7Va36EyrrkwanTapRcDCoIWci6ZQvSSGzK/Oaak18
7DmI5yHkhV7CmGcy9VP5421oWYw7vvTTm1SdXoyiBcJTSQrDODD66GzoqavkFs0uJ2n/tupLGZbW
QBYAOWrEKSSwcZcokw64DujW3WiAgSAX3fizHdcNxTG+WZxsFDsbYOu5oYb/N//o2pIZ9/30/jUK
4cC1lAA19anXAWTAQPMtBsQ04tNC+RPTWn9xd1fzrczSq/IKjuIJJ32cdUlFcnr+PTvxzzRh51Cw
WiL2h7w6MhNVfeggwfDo3kU5vR8S/lwQ1/4uRKO3Q0SYEJrJ6meli4pZ2WOiGl8dAKvilxWU05bs
IXF9fj+HJxK3/gV7K4Clwh7zcsoXu5eoKqk9mu7el/Q/9IXmY+IPXcedIUthPypHIlwhQrsKHCYy
eBqxrPeovHJz8iuxZ9DUF769qA5n/CAIn+ozokEoGgAk8tWHmnWkHRSr08f2XlXfAfIbfauCnitp
Dw14hYYmJKuOOa8Nlv1wW93hKEQlWwUQBgZXT/Nna1/aIOeeHIrooRT9nezyOjUnfQr/Zpyr8fVP
ff+Xx5tT5mYm74IDBomVMxQPpfal+jXyUJA4Raet1QhCF2oGDoE2vFRmOOir7TLn1bc66Ae+O6qI
Sue9BFEXQ6y7hy8QRy0RHFBwtNblJvPzZmq1dTWYFq+zh7ZfLslXJwyf/7s2/eOF5pEDM1PO0EVS
C9rhzCVJfaWKWdvnvTrXe57nJmMeaXIyvMb972zF5Ga1aQhkOXuzE4ka5niMR1mpEetztP5QKt0N
0ikvN6eUOU5RF2KD/pY5ZfTvyogPBc0Nqujr4aH1lkZYGSK6aoMkVZxzgAWFIMUAs2RlAE2nQn5e
iQ1q90vecbsrICB41omon+VdtzLv8m2Iq0Xx7AVIlffch/D9xWiVb21oB3hntZpvdz1QWhx4xLcC
NZFj4W5Dri5wz1L0p3wG+w7DkaG4XXWgy4yZUipNar4TRGBx7xqlfO6+NUTt7ZdHiF2rSpxWT/0Z
NQHiONpwFb/X7xH6PdCM+qIxVJZ2no2ysPTwrEOVBm0d/vE5DhQyqkgsZ87NbGlhYVlPkKRtXUar
iRxxvYykdcTGJwzxp0G52rfsbkVSn8EHTPi2h7BIe1IVSr4jXhE8E/A+M2yKjMhM7Ae/PmTJ6e12
M2s+h0qyNvI6pTTcdiy4/nonDeN92i1+KjA0OXtYVS0rVF8Op4VREzJ73SKYxYSCNsqmyoWYE/sl
Ck5CAqS05EcgRLDu/ibAcvTg623SZyAF092AJtQoLCDPHpiE+BRHjgu185FR0HUeZ/LqQOhjhSwU
SdoY/lfB5PYp+GKeN4Yd0a1bLpynagg67Oy20jzGM+hnwFMV4OrTYEhL1gjqinD7JNdz5AfvsjzZ
GNX6K+2xSkLSS8jIO1Y5dKezMLwuuG7JgUXTjIGNmZxQM/H8Zuehi6J+deH3MxhhgD3uGTmRGnwe
8bCY9oQsJRe5PBFqYUbkGEKqYidTHm4zCAhIefm98WJBE87M3jmA/x6o154452pqGyqiTn1eOSm8
gdpeqQu7ONyDrH0ZG3cSmNbnKmd7ycs9KZ4C+GD16MDwK5FvBpxJ7Kq7sA3asb1KXSxZNgFV/W5Q
sFKEfkMjDt7cksn9L36rOEgjdf+IVWOeYke61t3U8BAg9ckn5qMyEmyD8X+yEqjeRB/PqJg0Ocar
MeOqFqVU9VxVPd50ERKvFI7T+ZPPBYfBrmAO77SFlLBd9kfAhdcjrU79caRlBigxOO3ODsZbn7Tt
D3B6e76rhuG8kxbktGXCqZqmTyVOtOu83kfu9dKYi4HuJKwA5iIbUR8IsZylmUXrunJh8mH3DWW1
B0XBerIxf3C/HnAYwZSI5xui3M2HpWGdttU4Xo+n6jNzoKLvicDpgl5Qb4TOJv230EcdjyKWO6uA
feRfNZmA9F8Uo1S1eBsDRb8NSpEMSHI1S5zpdA8TfjJQELhOmNYqDc9PqJk3Vt3RYTxyjT9iYVjK
nTHcKpiU9/L0V+dvjeIYnoSrGG9KfjynF20eUk4tASlmAHlWPaCANmanOC38z1Y0AoI9PCpDLwaj
hEBNika6fYjYNBcoAB2+CwOZ3Hhop2SeoAfjo50WkAMRfsoQ0ML/vLNh2Y07Lhdmgh0ECTOiADrT
WfzUF6DdhC3PjfF1luBQeoI6PeGH1GuNonpNTxgaMJBEh2Mfx0ynwea4sNvF82rI3HICPj8Ko8Yk
SGwx+Ne85E1s0UFIavE95ffhxy5u8vrvqts7EbjgW+A67kdLBdYIRe5VDRpk5ZhzUMZ/3ahyd2Gc
eUFZyG9qnEhlFT0RWhOY6nWX8o/09Nf18mvXhIlQNtchSkw1iXDeCtmATg0kIJ68vg5jd5Tn74wN
s7dC1mpswypLK+dJMfSsn/3cPdp4tR30+BB02UI9EqCEVsJiM1YQWUqlNz8TBaWFT1b50W9JKwE/
sKmihcmmP2lt+QFjFEvhUZ5hCUwnOSc3BmPh/bSVciMpOZd4MU1QM6iRxjhem9XyTqCh+klIVzvc
95NX6TOmjTUwbzsnFJrMFGV/KSJ9fsAjuWMusZB1fde6p5tGRJfH/HVWb6IBJwHX7dcCL9ii6XcO
b35q2Eshs+4Id9850sHx7eMZdwP6DwCddttpzohoHTWXIRZRjlC8SRxoQ+q/so2krypQDayajdAR
YtdXOyhZ0nnzxhpaeBInJt1lJp/vtIeZl5IisjY4Zl6i/9M2T4FdXtnP6U7oUkbyJLqKsvO4iRiI
9J1B+ajPSgm1VYft8qcKYEiRde4V9gAnFOyEsQzIxYC/trydYky/xEdmEFlLsDvsdtxrjqrrQ8OQ
jtZEq+tWCHL2P38MBc4sAeFWUcwufqzBcQ11L7ScipNtY775MqVlQegBv2gJQ064aVYn+k2dk8ut
zc8yCnUXyRHvtnSsY8IkzormsXClnNEgchP1dFoZ1EEj5OElEa5AC/X1ZV+L24S8gr8TlYS7RcRj
d06L+Cz6fxwf7W1v3s4QFU2IFhKwVaprWBYB0MqkIJLgLtkwMqymyDld0vWpvCN9wrUkM00vy095
dps+YXhsl0mN/TSbo9+0tPFKjUf+J61O/2NADBmbc+NMqen/s1ZMUHE7K/R09QWWsz6gsuhebiV5
bd0cF7XWRXOdnzsvtvr5cjbNDYOlR5FywYuGU3GCI2OrY/FmPBN8fGk/azR/xVv0zBZtdHU4b5Sg
u6WqAZPjgOOaHE6gaEEUEp58UZ3ONPTZR0jBkmpbLhCsFBJMLuV50r0tdC2ZUf3BNSdj8ZDQfcIK
m95DQHkZcCLwiYrBaPVX+yycbdxB36BaTLN+stK1nOOYq3LX5DG8lOWEgqiU1Td6gjwv5dtKUdla
Vqalr6kCnXq5HaVpDQ4EnAzTBcE0OizhKepFQlb05O6E/yizwvnpOBQxcvd9+J2tan5POvhblMhx
7XwQcwzYVs/qJ7h9AdFAdrv6mw/5lvHrIO3FJZR2zv8wpnTcQnDVC/fKm6houYfctLn/ojafDcbK
yQxPDxPjFNqbaH46T/BtlXxFvC+KsFM5HrwLQuq8E/Q3M/LStDDA40PGYOyEIc9D1nod0+oRyLrN
h/9p8QwvjSnrJnPQyBtirKJVROJNtpX2kyiLdVir3qMSrjX89Li3PU5oogesh2mfMgXnjYmj22uh
ZAFV8VomG+kr/NBLQiIkxkVgqjIRAZb5hq3rpY9aMFK1fP/q5QOha9Hq9m6EyYmzEygBtvBFhOMV
xQLYxK1YI0+7vXmrRQblXU/bKWwNRCGhSy8GOVv+kBTPMtz6+2hU/HUJ3RpAV6B4L1qHSgYYtCLr
immIW5jvPLdUNxz8h19ZHpI39z7MbtRX1NKhqD0zBB6tfICBZIHZBVrNk+12QR61baJMhaI/YULG
iRmAdziSRRTmfG0L4/RWUM1n6ivpYFYAjgG1Y/JhX7Zphqqf9pEtyBomqoLQouDFfJJHUfEqknWa
8i7jtkFpVdG5CLqI7JgpIfqKEzvMHPCUyoniZ+XXBxfVLjHRxxduT7ewxEv+BU25/jE9oVzoDtJB
+oa6z/6uU1JKGUJjlMKq4gnXnBmZVvOGKGxYXY08+vkAR+o7sTt2+RQVeomfdhhTF+QYzMOZZRFM
JH7+TtYNjFOsuJB/UvvbXkSIsl9NQebtX83zU4tEQj1LyCyfAMsVELvt+3C+kQ+yqR7f0UZKaOgZ
HHAXmgNrgWfFuwdGqhZ0jfQGuqa92V/yYzThcqi7pnAIL9tkitr7qgXnyQRsX5i7Bn9CgTZ44+hK
bsDiTf0IrAPKkyisCXKpIs4dOvlFqkzRauGqA6xOZkxwzLzIf1L0WYW2EOPZdM4UYNdzgKP7Udc8
kHCQ05R5z0UFzHIXC7sXupOrPUGCU7WJNmHJCfc2nDTZLTw1zakEksAQZrmD6UvK4U5/sA4ldzyw
5etRQz5Pr6t7GouPT1LgJDjio2jjTfvVvZMV4RaVf3j8PwfNgzv/j2Osll0nC/I8TjRf3dKtuCN5
pMtRTS/wTusbKv0swxbjU55BGx/bq4RoTGhPb40yacWHnu2PpuRH+S+ra/HAbkI0Hcl+6NTEeSjL
16hr2zxDn7Gc71TD61YX+Qr9i+7GVL2foR5F68zqh34pF2HRZTX7BR5nd+CBagSgNiHoY2YOs4v7
sIsWXdrsiDjG0dlc7Jj6nR7/82o5N5UJy+ZA9M5mVO+FPtMbScZ76lreICbALa7gfD7nqgYv+Bos
We0FI9o0wjUj7MbTSiHb09TPf1TJ7aNzc3idU06fXYHGAjl3eqNfkplyqLXzvwaFFfDo195OCOIY
3nWwjB7Gke9qH8/Br7Up4F7VcYRbqkFPQcD6phMOxtrtaHwEJ8Bx5NCfPnW1X8oprJAbe3VjinDL
hxrluGmxEOrO/sY7Vtf33kShw/maNOAI+ROxRZv23KuaFwOwAIQIZ+BeINYdZ82lgBEgP1nmeNkX
ita0zmpCoZ4QVV1kmmSg7wpmlFlOv6ZwcWzUEvxH9MYksWH7Ap54UxjlOzJY/T6s2OWm7FMtNaJ2
Y0jL1Svv+wjsCj7VvWcKRfz3ezRdwbtYhHI5ql5NN5OyLaQGWea7bog139NSzeWxJKv6OIuvmKX1
9eTxWLtzrSMgsrYJour6/oblZvmXYYXFAot6oKnl5nFsikNlH9wEVCD97boehUjMpSLCQiHHDhyN
AMs2ahI1HV/Fxs7L8WXuYn61OZAVPeWeixDwYN3ClkNJnKnAtZzdeq9wQT8yI6MHcZaOikCSFFv3
Lsh9Tk7nkHAfL3EMNxGGnFvD+JZNTGy+2NArvs4Qb1avTTJ8wDfGLeJF5cxsP3Jzb3BCiD7f9uZv
zNS/CAJWQ7htbCxwWX1uU2+XwjDgaeV0YhZvZqdfxi+6Nhp7WcePSv0fstdYK6xkSfVdmKmPQDku
UZn3Gqk3YQR7ycbZqh9tlIMA9mrBXpxVJqAbub6I4leFAfn4ozErspJeiGo/C+rmm4POUgxV9Led
vUqqxdGzqwIGYvPNFatt1LVDYyHXInax8qS62cCjFeBaVU9b6prEObbvBcC91A95gIBgyZsSKUI7
EUj+BTMYKPxWRgnYYOPfRd6cwfCE1WGk3T3MqYutdBJrnsw00LRfIWRhLr7nqlayOYGal68hqQCZ
ykdjo/KlGtKQzKcFg3M2FHLWx63iIE5t62CpHmOgvj0/TGM6D0mr+EoF3BNcRrWBbLb5J0Wj/ZZ+
QwV6GuKoc+AYjy32plIogplvReRHcRwvdp5E1fTKcO5l8PnQfUEYe4I+n/mVQSc6SmtN9MSE2Mkz
22te/lUYiRpA4azxGwSV1fECSswdHuuroooa+iDf9T5PogQG7o9QJUxwHevvcCHHywOdO4e0WRxF
K7neO3xrl8cs9ohkIyvKDj93nriBZttDUppsHWVbhl5y85GFKAwgwIB6VwuVmWcyb7Vkb8dKf+t+
RrABzL1T2TlgTkyo4pyPmfNmSXUqOVqJB2B5D+MMS3Q1IeTkZIaXI5l78kCheBMc9lSikb+AUbMy
lpv75hOv6PXNeSIVk3OF+Kvs7bUYDsiurcbH3q+sj4XCadKPpJRF/FZ11wRjopLgpFNAc2zcW0zT
3KKMwjRc42N3nojWYMl/CRcYxsYSrT5cUeab0+fSco3oYEqDdgyB5eW8WKkH2u8/XhDk6QuTEmZ1
qsbq2nFuZJPRon5UnO2fD7CbttuA54yaYl8CxuJjU34nqC38sCX5AY8AucwP57L8hTLnkK3ju1lM
DH8gIuRDbOlFznXFSXSHJ3v3EpZuq2qig9ZclvKUgZ3R7B0ceCD+LR8P4ukMW/TkEThhhetExJTB
0dA+ZOXoRyBUlA+YDEshI4bd1ChkGq+y/X4t38jv5uavKegSmAP+PrFmLvygGJ9il723Xdjr8o+I
e2oSkx45alT1sLsZg2gEaetahp6KlwrdCZNCd8Fpw9MUAQYBv+t+N3qf5LsCsO6W0ZLlaBl0Wfvk
3krf+kwwo9Z2yGpIX0GpVlm2vb17rtLTIa0+Sqd0wz/0C3McXbQ+5j/AZViO/qi4EsdYbz/gwd6a
yxsB/61mx6+mRYMN+Ows3k6hi/qBQ4NrORDX9Cz0NESlpy3J4oCmrmm7O16RaVkY+6We8Otl2lQf
DP0efgUgE4coV8kn+hwdnBXJZgVRoE8WfwfS8+NpL+Sv1VnCjMfYhbPsfYLmFLWkWjwqyTCKL9RZ
sVYhRtuz1VSh7+9znA4/DIGxI+5UrDpb3lYRMP3WKBqGK4y5vMr+WRmz2PNSz52jUEEIDiD9V7WW
IBbZ8brm89kaNqfo3hxPCwkqWHMInhhNmPWwcFtQNzDeR5ZwDSmnm9ggTiLCK9nNVvDoaQpRgH/6
rhudoA1Idz8NTk6PnlpMTFOKyuOuSe9pbmAIXduEg4aoMtmkacCw04qIiUvot3YER053u3PP3S9b
sTFfS584G+aACHP++RpiUy07dGYL+ltA4vxGeGA3UMZL9fbFcv2UlryE5iYedYDiZDeqkSn8Sv62
VVsNRBBbYHCfSoaqAicI7XHxbehojbzVixSAcx3fkTkv2cdnrgN2r8D2teebNWdhpZ4np6+U84wU
UdHNt+6RZ2/XORrn29ljV7aDJIRbc8FUcbeqUsq9pjbyy3/7O/g2xbHrdUue5IHZ0WYaLbBokLh4
+XWRrswlUweZGNc7lDnzo2IdTWoIZTMxcDEPp7UXJUw6rYcrkEGgvsjfdfSQbG+8ahW62JxrWuE8
AeiRQJBwsllk91dlE3aKi8PO3Ep9ouBWvOltGMmQsJZMj7iPF9XTTJX+mTVAZfB20PfzBgB8QhaD
JcF5PKO9HDMglWyxlMW9UXF6BCnqzs4C0l9FWN98t3qhMM2BaGahqRmyGrP1pM9un1GX0xOiYXjy
Ciz06mJjAxlsWlzUDyyF0gaBHFAX+S+X2qCua8r47kustpoliN3CnrnW+pJW/8mRm5rP6DHp0Zr7
iCKTLFF9uSpos3LwUAXYrnHlN7c7lz0hlGCos3m2TNGirSCBhn/KQmlzYjENImrhXGNMhHktHu3z
iAFVfLg/Ij/ROyxbG3Xl0kP6aNHuGYAcCda/70rexrAbPmLpkddKo0jerrumq7tgBW0R8ClDcbEM
TtfgtV9aYS4gHevaZ8uwgtqXHP37/2dmOlvK9zHddJTxFvx+de05zb3TFbMQ7FYsa5Z0TcsTIsCO
ZUhnYHQuI30AtLDlB9BTY6x3cuhUT/zxmysvj9ouAw8OffzCZOAEqJyU07X8YbfcJyu7ZrzJ4l6n
m7hUlMhALjcDHermVWjfyc5lKFqUEZ89xHTn5u/DJ+pblB/fahoCBodCQctxH049y5kdeBFp/BN4
/JSSWIC6Ai5NnQCsvXqac0suLoSP/0wC/N8UXwYnIYH6WQFsPsOXkcS4Ja0Ka1aKJUm/Rr74ngRi
e4UajAatsnCeLM2HpjWC5474OYr7HIIFH/zVo0tki9vvO+Tn4UuHidAWXTAtYMnnZpPgbQlbzRsP
xgO2xSqSzs2I+KVH9VyuVdXPS97Yah5m5NPeoChOIQqRV1y4dwqhkRG7aRc6kLb2MIHWkjdl5Ohu
xfxlMM0tD0KN0YCEpuym8xftpaIuT8ODw7Vwr4Yq7Ng15UMobEpGkmbrm2fDdGWtQ39tK/HHtwbd
T7vWqyqd249KJa5FqwIYU3DWUsx6ya+wW2f7J9VII4ya94Du3uhOEE7fTnMrYboyNjWT/C1Mze27
DZDHRmCqyKQGB7DEe/Eh9kZNneUM4UaFLml56Zp0b88/VMd2SAe27ic2Lfy450hRMJ5Wm1OM0J84
Uc/7cxH7bXdCK20tu1xSC2bIR0JMbWimtO20aOFeZ31tr4mtrfizP1/35nJ9A7U1Vrt9XXRRyfkg
cqPITQf2XpDSXRcQEZJkxRrqm/Re+B3pYLScW0Eq5jTqDUq9rdawRQnVEdDWtJSv5IQQn+fGG3Z7
hCjQ0/lvCKdy0s2wAgsfGjXWZRxRIIwMc41dXj3/zF7M1tjVWuVYwE4Is2SV9a9JdAgk/gBIRqcV
JIgHsacMeCKAKLoaKBRwrh1E007EJ6juonKKYMbX/j+GRjMA+kC0XXe+djkN5rY1M3vsWOnltMXJ
rUA149et+PQmZJzvg4dgDazOYCFCDCHpDHKcJCmMc6bP56W+HLkd/OjdiiuE4T+hdca1TzmxIXej
ZoEl8rQcDkp/E9F47ONVvhk1xUIfRAIsR2aQ+Wcn2uSC5O2769cKGcAYaiZv+h7ZyG2KsOt+/Kbb
CC3+K77xf/mp2oL07U3POGumFiTYDi+ySDnYA39/kzq5FK4B+0o0WIjZ1Wg8cXix1gydP3s48T66
3Y2KwRMv60MBac+hWe6pKV7O0m/+RIl4jm7AJHZ/AJ41UVmd3TJj5Ft0JRUpTDcc7wkpeq57Ovox
e6TTzIZDhnNC2CoItQvkshLl2jB1ra/3rWnc7F9nmq7mHPLVzDe3z1eRBnlNAWywwjnm951FTYmZ
3sccwb10vI3c1IDd8ANsmXwKyiX8fk9WGZPAL7qhFx/OzFGXwIeubZ3DoiB0U/UPyn70+5VxzBVP
gXJMIZRDHzpg7QVpXX4d6i9Rykovs/bffSA8uaVh8kXSdU7y9Zk/nPg+ry6LhEVPXlsFSYRSTmp8
XoJ6PGgSQQdZ6Rn99IIzqxnko6ivSzo91jCezxvsgDEsn0aC+0yHbR7GszRFK+ABNezETkwNZ0in
cKsUNllqINNsmogQvK0LVujvgwqSrlStOHx8Jc0390X3lIW9syrjVsII+5g4z7kPYKDM5ie2oKKz
NvV4C9YrPSTkwEHM39rocLSAZAfkjZcUgKZqYhTgbgQS9XwKnpW/MKelwzj759N6oKKg5wvJaHoj
V9mQsOH+ju+E+7R2KdTgB2ovmtU+nfh75vwUNt+MAychg0D4WtbuoUh9M0D9vORsRkhomHhLQ6RT
sPf3dnNxHX+ttrhQknA+fmYsW3OGhwnbVvzjsLCBjWmOvBolYTC0+xLxrlm9hjz4Df39HUDl7eoO
H43CAZWnf2/YskVQHF7R34DfmEm9493MkKdwn5/MYMHjFCU5jeIV4I2aIg74DZgEFw0XrDcF1Ifd
4xrWHggyrv5JohfEz4Q4JeTZJ/QKMnNkurbBdgve6x/XX+jR3Gm1SqXuEi4pDiOsrHwQrs6yTKVi
xa2VoUe/k6CCAJjSRLnSsecSGhALNXv/gtQIGfTrwLT9rPk+cPjnRPZrm8UFn8n3p0wcBob8SbNV
blDIZ24PWxaE2hhA8PPnmAllXC1uVLiolkHJ936fPdOkn0Xr7z4iovAX/ZxNhoJETcsHxLHlroCj
6gV7v9D75bfiAqK6f6PB5oT5+4Dtw0uLDpCJkNy3GBegoAfEnPTVmETE/SBbswEqi0vqVDwmSl9C
F4ugaAAetGZmFhKnKffBiJ46H0CBW0OEr5Rxb5QoLGHeVEH4b71y+zfx3WMo+lJcu5YM4L+S1xEH
jw8YG+nKoucJIsXceliDo0vt7NsDgVTy2kS2O1VEtQ3CXtpAVle9RBFRKF5VjONoEGXgUXh5W9BL
Q7otcg2bAcDUQIGnsYwyfzocW65fDegcvpq6/QNgaKaKn0f5fKPvozCwI+UyvNES4N5DRzL4DuS/
uNNYqh0jOD9D09yM1NRdnNiBhil1a4LitMGKxi2kSacQ68Ra7A0rr2XZKy+5+zqx3Opa9U92Hcyc
3wCYlZf1N1/ql9427hZfg1GHmqyeDWPyCskgzAcLHFF/2h1gbjqVRxJjsKYSeNLdYaN8KNH6CCnl
OWv2zZvOCtn50iFFlzkUGxHowLzI2/+O0yDX+QbXdMGkxm4uGiXatjyEFOy8JuQxHClsW2eGe94i
ceKbpocc2gMEFnCq9WXcQjCvj9cql8+vW7MsAESyvGLBEfSPxKlnmkdwjM55f4qdy6a3Agl3AGBH
HHVaVtC9/yfkzD1GD+i66G3G971mVOu3TzJHvut+CrWL9cUxSsB+wAgcyJvaHaTQSss/9aAK/uWd
Mp8VwA1f//5YvW4xfp/hfwHMR68APcjMwegkGIZF2C579y5HOAjVdK/DF9vbVVKJB1RbsEBBCgSz
mM0B6xNJkbgOwqetgDqvk+urtvz3jkKSzXigsS16W5zxFgQyd4kG5TarM40qI7uOZEGNkvM76jO1
Rq+b0BmQb7RdIe+Lxmp/W/TSCTtCpWIgYrBNKexX7O5cTRbMeda6ogRbxl43+eZ3xuQn/C7IovdE
tT0IVQbPOd7S+F4wXtPMS5lr/BBfulWtf7gWKKVSyCzyziLZMhZIXspFd2uapRoJEOHerlzhpC7k
bu503iXQBO3vcr+mhHaPY5G44XFCm4ygTCYzq5dMTQ+uA85dWPK4uLp/HHE84tlrcTPxYIwH6DO6
N7KBKgBQDRsWHEAMWar7PSJv0USCWr2zmQzyiWMVEM/nW4ZfeQuq6dnsF83VRPKl4kQ/aXLLJOY+
E8jO1hul15pC8scXXtPbfhinHiM7r5Ez8KZF68dRcnyOlfd5AGoWl1Ayb6XSduk+iv9+ZUSzc5Hy
K7VyqoTcD/2hmPQFTcLxrAY0bpaCgzd69aUy6fh7OYoe0xfHr9s2P4feK/bHOpgOI7F1zDtjtbpQ
bPqlPJv/9IHD7Brdr0+FA5T6p89+cmBBGOoHwQXwbcHYWk9wY+DSXaSeUf5gcLSnz/p+KA91Rrdy
IZjGv5z2oC88JTYGMyMpjIchdwYJ57IH/GiOkUR29pMQWveehmotOAiO78Os7o6m30t/qQlEsjjC
bhFvqIpqjyffSvSko7R4kIZIcOYwFMPX7tdYn5TEtR5ErFKMkFFUMIlRUHkHxfywGY3O9ljfvUjK
AM/O6m9GUHoW1QFU+6G1RvWTDAbQ/d3/RJc7O796NhXB/0PNBt7umJqlvWZq8an1lmLM0OZngfz6
6tWm4zWo1PVZz3tgEBlA29ZBXhCI4zj8024HZhJfVGow0PLhKXgLLp/ZRRmdP/MwDVFMV3tsxOpx
V6DHRK2woclhqs/6cNy7EEjPFvZUSJLUEJYWyFy8W39aJ9yXNzvIiW3JEzfkuJ4DbsuEeWMKYdS3
5Px3ydHg+tHZjMHtwviOlygjWQkFrS1Eo9SvZtdrqEVAzRBQsSbY80SdT/j+Ie0k1x94cZ+4NpOY
3Eh5fnTfgVjFfuFiPjFFVJ6SMVn9rHWTwmecaFdNigLFtv7TCNAKsK+qhSG28Y3zX7fq3HMdlZfA
L9kaSm+eGqvtXKqHeFhL67QnlsiHh5Ib9UpeN8cM2/sUndzEKdWHWb50QaiHD25lagsB3XzO2U8X
5eXliHWLar7tIy2JaSAp9Xbarb3NIte0BivI7BdLGP3guHvtCI0yBl4CtRugt+WLH0c5vCwtr/B4
0J+cmNIKismvr6cPjKX9/PLcqevWPAnggmitOlBj+PEZbRzZ7+MMT01yE5EO5+DEg40VmRYmNqja
zmMICEGlhSgPA0A0VgfJME9O4hJ8DZlsYIO1vQNlZxQBbACaCKyJOKjkSy3g/QNq36CIflMoZkCM
8edFHNKdUsGe6rqOLFIqBBe2sV7LlW3iHzZsQacJ7o4o1vCSqEu/7jFw2OzVEPpSX9RosqibYnPl
/E/ADTt2lVZvb25cyhGMn3qvlUOWB69MPz50iUpWuYlGnUkJpPIhEv1bSMTWRILQuhH4uOy15R1i
RMnaqLXs07rFzJg+shDBVud2siHBKP/fIviz35cNd+yHwTml8JajUi9u4CJRMzmnxQMJ+Iv5kTVl
lmhn87N5Dk4bwCjb1jKPVnPoHBwVlkTfddfbC3uvtZXDvDkSDao9cWKjOs4+S+BILshD534qYQ0H
DsqB4NjQ337dmoy6a5DOFG4Z5w80o/9n3QQRfSg0LyB8o3NAX2hDaboKHNf5ITwlXgthA7I2MW1/
XOxYn1mcJK79IKIArbVZFWrHHC4ganDXoIhZ1FkK64ZbCqrKn/Ja50U+ZSLh1cZg0NRd8Ei2CVHc
GDyrgsN0hEsRCM8mQ378kt/k0XbxWZvnPyKX/HrLJLiErkoOMydI3YHi9dl3NwkDOogapdbdMFo6
Uphh0Hnr1N5qq+UHQxouHSZqJKoJRbsgCMI16i7I34BZjWIUcX46QmKtH7AAAOju5eecNqJ+2cna
CUjfN2mE27O+XpKKhCJWzOl35uhP6yiFsg35ML9Vd+LcaRlpYDmd7oHgwNan5uRtV9/BzglHyp/5
QzjqFLqnnt6lnaquGONsbxaRn2dJRbzAgB8ZWoCradcRjRbjc4FaSj7G17lJsbKLCE7x0Z6fslaB
aRLhaeuHbAzOdZ5pPc7sUHKeElM5mCf+eLvBaasPWIWw6Co1eob1LU2pi4EHnhrkg5lh2vckR17f
9g8vCLxzer/pdwGBS9szghsN4SLTTTSfB3McGcpqOUngDUKdwnmMOfj/80NcTx04d5Lcp6qjvlpN
6uVToE6a10oeMiWnh+eIFqJCGYgLxPA8gRgh7bT322FvYRqRLWQblFLWqLR3ZJGIEhHDKOSK22Yr
563GKa/qdEVLScLjZYfp2bms9I192jKV5KMcGx+EY/NfUbixzNrT9/DRC0qPLVcDdFylFS5h2Cga
B/MGRZ5iRJ+XJp/tq6rbdrSpVjQufjsu4kf2hKPSNlya1ENyv+lHOSUplW4+kN8iDbUC10jFn7Kg
qj4Yom3wTXGLeKDezoF38vnZz2iZc97EMI27Rs4zmCb1db7Y5bJU0gFPFCvmYZKog2+Uiqt5RD3q
JBUcgjQjmpvbkbv4S38zHMoEB0P9yPCuNialOayUoF4ursSEOnnboRCC75fV1yyTzDpwNf4NEdcD
RXeOFjkAZ20OqE3YiOxCH/s/KsksLBi+of631DaIe716WrM0tvjpHYd8/nAlvFCLKmVHGnXHxqym
KjB95hlgg2hBfsnCfXQN9mBPqxPGd/HR5f3MX0HkPSZEXwIa9R1vtZHRBsaYlX25tjZ2J/05Mi8E
aXF+5ZB7NrhU5emls4RKBSa2LUWPH3av2tDpcy3e3B23TR0zdy8NfGdqbVyIqw9ITNTKLNb0XVoO
IsHYA/MU33W/t3HyNL7KRrkVuSEklFubpa59pwB/UlFSyg/tSvcJ6ZONLAN16nRh2snQZ0R6Uu/v
RUsYKxzcFfeKU6jBoEcNfxLIrhJjbDJx5q1fzGAXnFLVr0axckGSkW7lclx4oGp81yHTR/ag+JDV
kr37dDdprYpXhU0qN2MCnxw+JO8j4aOkYtZMuilUrrdFzim4C9NsJw42CCaqgFbbcJ4YlqINfvNA
BfzyZvwqigfSP5OctqfpWPFKe+EqIBP+n1ZBiOkITungCD+gJc5sRXtsPizRVE//rAQLuN7IN72W
Ln0VDc43GfhUQIQudrpDkDXeBC8S9HKLUdoVmE9RK11gxMdikW0tOSUiih8bJZyLR0ZALaPrHtO9
5Tj88NR2DZl94nnxZAB4u9tXbhsiFcQYTuC33XdNphLJJvFLHuSwK57CKDnuqZmvHG+FwS/dduTe
N3fRqQogxptWzcRXXJUBNZEgbl4jpIrkhIYZihMmulibFO48uWDb9LsO/mqz1fcCTW21IhJaj0FJ
kBzFo3FqvAshdICy1gtrROLlvn5Z5nOJRWsI9YIF/pvh7vCfiA9ZHuvioM1VF4a57DTZmTzUNQND
QRpwykaGDSG4gy7XigkIydm5WtuGZvWXHuGLesAGxOy+wpFnv1g6+h46yPkaM9Qe+tCZjO7Xig7+
B8y65grxXivD/VnHpdnivaVM00VDZGZgVJfHEmFhPnFxmTO2ihXfVlNA5SFhfdpiyfM/NqZzuRsh
oyN/f6tnmCGekAzhZFnPANKeuYphyKu9nvT3DUeILOVApLmWhbXy5AgHBw2vanA1/ehf46mysgbe
rEbLx0titAhxWZc4WLGY+Edc/fK+6kYTRvAmkfiljB6Rq2lJP6do4HgoKU4S4iW1H87X3uH9MFwi
MuO5UxriCjzlFknb4Yvbuq4Std/50dLa5BTT1yMX+jo+SLK3VhD1LbDqXumNdmV1b4SWoVZ6/9ui
RaW8Och7LZVMJAaVgTNCcuGZCVv0zprcqeNPErkt89VTjjPRhu8zNbRFvTwVO4/jmzmWA5RzQAD1
Vdf6++BMGIZSUJjijGjMP3HsUAB6Klj58VzbbwzS7LJF3gAf3pkrcYYdT3hu1TyvEs5nYde5xgDb
Xvk5n99+qmKxDP20mxGcEI2jOE04SbqbqbaSQE/6ExFSiB9xl5TxtPtZaGSFGFa3fO9vOP83cgEN
kxsjkFKHOWnnRDuzLXrCBy2XT9gwtGe1FvHLbQ0P3Z7G3zR8pxNrzswyoDljvPMEjykusRPDmOsv
/MbtDLukPHY9hzR5Xja4z1LF2ZmlOKzU9V/S8Wq34JFojGYujplOOSP5G5gnpRYR7h3hR1z1In1B
VMOJo25SlSxOPBd/4Ha8DKnltehPiwFmfWLAaInjnoRL4ZAty8wz6KoMBazVR7ZDQzGhsTH+wZGp
9Z+PokdlsLwaZTdsV1ZusMbJ4Ow/qdEkWQ6xFKLMBk8SAfoWO+JDMUYIa/rciO15ooBCY2/otGOU
68fjiKcbTR/LMky1j1JqRqxoTW/z2yFtEv7X6TrcEoioecZh1VIWcL/TflPBRfi1ppptderRKh2T
AlqfUwXveuYLasUtgbohgMl/OA0hYBekEW++XNZNJRT92rG832/01UbaQZoVuFBhv5/LTcp0CEJA
YAlnT4KzeNiaRKK4toJOeBJHFKGAFVxsDlr6fQBGGmaU9RmPg9HbodBPAHL/jl9BmmC6ygGCcs2s
P9BLAjNuiRMa28RJzytzNnRdJ23apDl2ZmIu0j/poJ7XieuDXAxgJgaGGneiK/Gao73Fp0BWnyPM
ZYCwaKCIDr6XHFJDzP9jSMqjnsOVFjQqxfU6DpRGJy83BGHzHQGzib8odCriyFpPqf/0D9/l/7hs
xcLp7AuCDudT8Oy2wBg53qfqk8Cmu093y4K0hua9uCFh+744ozfgAld9GdmJ+rRRU+/9Url+9wIc
QmrlAgB5QYt64Ed2erVWes8pMJAcHTRWznoz1WFbcu4H/C6IUgUtYpOHzAkxnpWV6YE22kSLUlxt
+UV98UeYUOi0zmzA/PtpwLuE5EFXiB1F34iKVmhRXR323GAMMcxDUKFHKdEGnaxS/1cwMkv93DQP
K7xHpuThmzrQZBcNo3OFjHnrQHNai4e53YGfC3nl2YAQW9YLj1H/M5Upds5aOIFLBGtz0Rgy9+k0
T14aqCZv0bOaopn8hCHek0yLVLG5rmV6Egn630pnL8h6j2ET2BnEsT6pHlBg3bKwiS4ZoxfyMpwO
4OCeym5OBrEdh9GXx+HSKCKm/wJWk7VQbHrt0LfpcAX2vNajSniauE4nNmjliGr6DBqDpya1G8qf
+bktPbm9XRCtpOyxRX80WzWO/z6JJtOT+oEGymc83o97eLWKW8IInjSTcjKDMWEuEHw2GAB6w5x0
GYXnibnWh00d4zKhqLKouVBJI2biH7d9ofoT59tX8q31PVtps9Ww0DCrmAtTPhqKbtAvugT+2E9N
mHCsmweq4TO0gF8grsfqJlXpimlE+iSGMF+E5Ra5AX7yW970xky8iNSj2VXlScmP9gH3RK74kmNs
42SDRMxUuqey9JviTVecmgX81M5z6T71hSIi0KL4cQwV+pePx2N9jG+zVH7eteHN34JM21lX0YPH
cGoOGE+Lc51tc7rwmGad9Pwr10IwKKfwjB1HjvroFohKOZnqILqCvr/GivI5PMVIG6qT0+fZ8Zvl
N+l8vjuxxpb/ZQxAtVnTJ0/2gSNh/psWsF/Y1TtuFiN9WFcyaMAYpk0dirYD+7at6e7ylr1avOMW
I9IbGleLXm3bRLjpO6hde6tVeNAWDmQDAIzKnv/beT6lPcXVJb8HDauHEGaZ0EinDToCY8N1ozX/
lK32HBnV85IRo/xv/WnEmrJhMr0H+qEhwd7JtE4xeokPp7aMnPa1G75ySwZMZ/E9MNucUrm/g3Vi
ibQq6XsLNdCvA1P6fMRuc2fLFYez42E18H6JRdQhe2LoqSn9hvMxzzHmEBLhv1mo4oGdRnfJ6gg3
/tJ3aAb2K5OUnNmS36IsxxX7iyfWr96t451R72XvZEApKcLC64EdVGtl3EUsXdRHhO+oOf2a6ABq
qsIHEzS5Jue9vDzgMB14PwBqJY1qhiaBX57nwE36Aigic3/FEIRp4FaVCq0vk8iFOmNwM0HOBzxH
WzBngRRToiYFUv86dxRGWZXxU11aNqjKijSaBUWtOAgbSICMBB9w3yvwjXbbK+tv1eOhztKKHRta
3xS2TwZCTjp5DFcONLcMnC67EssHA1WDP2ZHoDKspypdhBXMtVWWhAQq4wOYPwp5euGwswfx1W8E
a2T57JKLQwZPMJ1hF0QGPH805KCVmRv312yZEoVv2H6Of35kf+ueuVEO9GSN6ItsOKTL1JyuEOVw
jJ5pv1xDUj1Ecq9wfqpC9SupTFu5+l1wgWuqtzvH93mPIbzh5ICIBc9rNu7FUA8Uj+ZPjjUKK+hR
7h7uPE7PE0p/Ujc5gxzSbb5nLlw3go+NGUOXeiXlMCqiBBL5fseo4kdYbqnBtGptT4+NxLt2TZee
7DPNavajdIMmQ7Dvp5l1SNO6cIARPttzMv7dlUSGDjnTs8Q80i7U4l++l+skFhm5V4VskSzzD5O8
GflWLmfczjxtJ1aIQNg/oDz4GfI6gpHXfZ0zmw74XGFiepJAk5TvHxFyuEDZ+W+UsA0yYbHV+3b4
raxezD2zXjAj+Sf9/AW4OI2Y841ZQjXIfy0WtZmrQpWN/j7EA94cTdejblZM6VF+55Ix9hk6gwaZ
fzcpWts6e/U5FT4+fdyv6bJqTe00NI/Nx9zCFdXakqFyGbxZZ+9mcTDjXuCjSXPeIESK6JEtAs03
Vd141Sgoah9TfSd6J83jb6R1U4A+iLQziL1hftSELzdcHr6oZGKaG/xXvv0dd8wjG62bvx4Qq9HU
v9X02jdE8/tTTBp89po8lTGHeFIPgJ6CtNletxQE107q9sRTDcEOSDBOp0D4L3v2DtYrnNuAEGx5
/J6Qm1izcJ+9tOuoUggGOlBpReJDCnImP+XyvWWhhbvhcdMaGYbrA4HbG6XFphMp5EHdU+MmAbCp
KwnlsH1ZQ7czjUjKdO8blVmlzVXtoBBW7Rg4qLQttXu8MpV1qptbBI9ZruTQu97Drr36WXRvXN/u
d1RmvUXy5qHg64B0vkReQKbUO+841rsPWlpVy4QuBgixNAgnK4HnFY4L/8wRTUaS/dn+OR4YKKcd
ZXe1xxGFt57hxL/VCMD3JiPY3fM01Ez2EeAkaFQvFtGd40AKoYUzapW4VB9kOsD5vTorxMdXEg4B
n/5FW8B15WVgQlUZA1BzoquzFLU1EGw8s9lPqDR+QDwyaN3FHp3SwqOCEXYSuuJ9+DihMMHx9ksD
vuwhnyFMob+s5nTM6EkJqtpmwCWfqDBa+ykbG4KBBx3Xa2t0X3m/mTrn+pUUEOGwJvMMX3bREf98
6zgVm4j+gkRgGzO8ldId/IA6N/NoHNCyy3CnLbsz4ID0Zp19ZXYLA+j0mSWqCMk92QBbXvSK3giw
nQmphWjD3yRKYvJtUMFh9RpmfqydIZx3FemrMoplNlK9PD68TuWrD7VGvEhnCtWUfQq0MSvspDU/
jfelqs6+S4Lle3a7kRk3Do5Z0zuYCAO+1EzH1d+dleTXPhe2l/ydkiJVe/oe7V4EHXQnONzNM/lr
u8QH9hstzfe/Wr/5ewINGOLWZRqTnJUmIr7hZEaBdoyrmXto2Q2Xx/0iCu6/cEb79FR49sI1qZR5
WXxdEnng9/fDkenw3k9z96pI6YTVZJiyoBqh7426w8Fkp91iXTUqY1xX/fE/RyH+tGue7NkhbLGr
pW3JAKWVg19SO+SdBJAmzUjEcJP4df/OCubspjSTJYq5ZvhwL4y8kz4f9ehAphluz+pHxkbp+bq7
wcgHhA+lA/GbMuCsJYVE4xw8uq1W0mzBMnfTP0PdppQIUl1YplQzBuvNRut5hcsES1VCG8w6TOze
pCRIPA1EWJFZL6Jn9Dpt12PSd/qOukkob5UVcW4TislBWVs9Aw1wkJ9C4eABOjlnZyRur2NQZ3Ed
0Qg+C088C26OUrYJpcVnirpKnUnwsxvHgILXaw/Ux+UkqVV4smrugqOL/wNN2/dd3oL2LUxs0mSL
CcXorCa1bNd2lGvR0zLRqfO1kFssnfHw8OZ4nPoWhf5xdTs/DwSa7dOqSn1S6nr9qVJuwi1Z3cjF
muq1MqyUeBhCwWQjeMulvzsnwmPwShoWtIYCDSvnrbGA1zmL27Q4MoLVPO9F6NGSvHRhQeF7+nvQ
9Yc5deanJHAu4Jua/sigO5cbP+XdIPVg2HnLmNC2XOV9CRq+83Iis9h9YRUm48qgAoO2j+/kiVHZ
RWBnQtkUE3HHTroAkg9je9jIQwC4LmCic8xzG9SmXHFjo9JQHaD4fuyV6T2bTozug36T+ilum+GP
cmbeRTw5MXmxcHTD8sTaJmndO/1HXP/qRf5F+J6XETSCK8Pbty9yC5E9arFqphXtmaiqhngFxQcU
64WbcI4TITA9PyyTGKLHD7rx83B9yPYfvEP2ZHI/P1E2RhhcUzQAp+h4VNSIe/z/Yl7nJimrA7gG
4348fJ1JGFKfwnJG2phzv7hy2oqd3wH8WpUNd6dkMSrstoUmV5l46qGNIoYRpAYcd/Mrj/RmXcZn
Z1UbVNwD9FlZwIOwWs52Dmfd8Gf8k3aauq4E2PDJZHYKj28/YZmJ67cWm4dPsHkdyyEibL1pRWHQ
THNxMBiifahj+WEXqk4Izk6vo/701N9Ajt0We3HuHmB33X0TiW0yndvAvbmyvUtUu7QV/JrLJVuv
GtEJu+yIFFVdhIX19voOip39d7zELiisuxhoyJQBNcPjJUfPL1JPSA9jerwoMDYPMV0xLKFS2jl+
aWiqaEVsbqogLRO1sHaK6qQnD+E8NfHyws3PmMCZd6h8ajXNHJa2xc2GY/L3hklKO+cDZXQgS0Mv
LhqKs2rWELRTsQr4+GCbUIlE4Elu1h2eCvv6Nwi+XpSjQsP7tJIXexZPOp/8UbLqFVtCLoclx8S7
hhypPuP3aiDRMOvHmxkwduzexn5+2S5h9vjhreR+P6sEfKfVhuuWm0I4M3wvm8fI9kbjD7WDkpoJ
wTW5nHDbHfL+d6o2hGiU5+4VT/fRrsRmsROdQ2nAhcamMrEF3JlCfeKyAO7spKTlaAxp40qRkF5Q
GgmBxrlyK29Cc/sUfg5Yb9YGLNF1O9K6f91iJwIaWMhV6s+jRpud5gPbUI/5a6Jb4hOlLNDieSrV
0Hfqa7utLjz/4JtjNRVakxqwHVbJ/wZereDAECUJHQTkNPTLW9g5ilTv1MDuLT0eYq8kDOJhYe0I
QOTfCwdZ23JYXKLdN2siMCzo6u2/ULAup1oZewBkb5T1/+wjrBL8Gy80gs06+oQQ2DCAUf/DN0P+
FUsEhoqQc7y0YUGrX/1E066V8ID+RqR7uKV/R8Le5A3EDQzJeFBG3KZ+utIWG4/mFn+Dtg/i1S60
KueCkcPBQDu6Fq3QoIhmjm1Z6gKEmtKsJB9jvW83XIodsPxYzEaDBFQwTwvvZTCY9aMZmOqvyAig
mX8YCAD/GTwCUNjs6Mhacb9PW3MUwhEVyES+EPwGgJEnHN6HHZgj9SBU34wwewviohtirgcF5OQR
H6MEzehdEuDvJP+m5Bmf1dNRA80+HFyImKVCZsYuc1bLnWCymyIPCaGf04zpIuu9d3LYz9FhKCsr
Gxz/RFi3QmrSIovxQ6DQDf3cACad8tgrMrW9FFYiPL0L1dx46VxCb5+UP9cto3X/Ukk/pNkBwPYu
8QURYJrPavMECeGF57PLWm9PG/fC7IwZWbgYN4skDor2QBv5RXprb8xp7ddsi1P2UnPuPBuDFnrs
HV/XtijlRUVSvxqTNER81mhOJFh1ykTwrj9FVumMQjqm7jDnCkUkDmiHE1fNynLvPQrsjDVyKasI
NAmDf6JjIfXPbkbrrS33tnIUU1NdwPO/KZO1uoqq9uS0TstaZ8RvKW1PR+RTyre5d+kC9JGFWeQx
Z4WW2KHwE955UOnSvyGISoVeeacVwMLVDPcY9ITF6a/DDdlu7y7AXLyeWwQ3nJwb+g0HPG6LCOfn
JK8hcGmOrzr36Xk+2Dekt8j3GlRT/iHdEpZ/UccJ/DkDSZJcktYUHS8d0H5M8rNiMpdha+ef8YE2
rxiagtavk/w3GUZjT1a3A63vRMc/npTijCY/XNip2hknkJX5HA8LBkvM5BwjttFXOKr2quAV8Dko
ysTT+KrOcSBj2BlZt6+VmfYY8iGfzFvz5XhM4dKg35bwpznHziYD4gcejC/jOx1UzSAwKQUMvcVB
hzFog82+nHGB2d5YQ9A+0vrbWiTyAp4slPflefRE163GRcGI+Oqo4+5H71NxxEtUVM3q6Jjbbz5r
pFLIdHVcD9fmGDxPsVYB9lHVDXyOx/H834gICtcBhR3s67TqjsfMO1EzsFpXbvDuWSrOgpycslJm
TDWd+OP5050wH2Xe1aM/YrSepulSmUL5EjM7HENIEunkh3xP/uCkMSWKukcamXP6NrGGhvBeak18
VKSi6AQ7CmEnOi5RP2E1Wb5Xd2HNDScXbH176uvwlVS5Tk3RMgRfcOPcoen0eEi+AVLfEKpzytOp
95dGqaGqFnb4eeMhBmATTWaLu3zfsftVQVgyfKFvdXePpjebAnTIpzUO3sASFB6mkazhhcECVnFk
H9Yoht833q96J+ErBJXVQyCrIVM8BSQTAH94wn8tVUCTHug63GBGUIkcExyQ4F/9eIaQwn7wmtz2
QNgT5bDJ+Igi62ZK56uju/j3/BQsUFA9sd2LZUuTk3G9BdonJBTyn2/uQyjpBlRHi6XD/pzgZdx4
oTzjxQvqHIZYQKwyBvQmFD2UBhsFhbTcMGMCm7lPCTZRVqOgV0qc9eZGuw0kXSAVmB4IZEaT5KPz
qKRLXEZXmjlHNDC5jAogEdtbKizNZtexAhZf/vVE1sGdz3Qbu2awkfESEWFlO9gd5tV25rQ13Y94
wlIK5gPlD9dz2Qd9ii4Ry+r3qjK7xZYAkHs7GuV7OztukYvgkC4raZ+cwP65XJn0F/6YmWTxqHRI
1+sctDd8YFYMm6JPf3KLnAJS2ctxRElMCYSHCezNSH+l8v8uMlYOGuf02hAw7YN3B24pqoP79PCg
+seKFFM8PJ/YXFUZIRDhN33xDh7CPFrN4YTuzjporFD3Aohjfrr0XZa6bG5Y+MV9Z4Mo7pBreQiK
kam7pFdTHWXFpl8NssohayduyjxlcWS8GfOCB6ocaNk3DAEjbCtuTyUbA0+SwL7/qVczIfiYBWxm
WrApY0OBT3GNeaRRJ3DVQM4alPfX9vh68IURzKy0SXYSxbN1COET7cd1eInVU/63e4BzoYdwT/9+
RgZ3cegISD0IRvoD77oJEO/M8s2ucsG4rciFNNujPStLwJKzpXJyqciUitfhH5fN4sDbMe86HOMg
p2eQyNvjdEeMV75nOPvMJ3GD2T0V1fxNHP3h7iyQWGNYgftXQYmKNFCZEx3FdgSlEizay7cPhrq4
ijpNwTwQY1ELgDIvXOWCbLgshDJ1U1frRT7FjUC3egpQOCS8N+LckcMOaz9v5eNGbz/QZ3ysWq+b
2Gnyv6WVBwM64m0YLS0ao090ZNwZ1MyipniJg5eUV1bCGj3Kr5+ns7r415kTTjLOHFhRDeJcWLwz
Scpst9iHzWj+GdBEV8Lg3JxyBqye98n3mpPMXrGqHTRDcnIYzB4AKuHgfs9BMOgTH7iiA8SDQ5Eb
PHZArMnUjo0woYxoN0i4Ddasg6QnKZgf2zLImC2Jv3wC0mtIYHEz6BNreGp6Svn/ZKEvTP3puHa7
g6ro8mGCWGvIR3nrhxJpL/+DubpXMt8vLlsviflqDjKsBp+a3ZTDbHT80u+KJKN6tclvLpgYvHeZ
wQdykbp0qEeioXAJTWOlYYqn4ztw614j4qCdjoI+hUxlJy3BYdnPzPYo0NsXN8RxwXkCmLOJFdjQ
TmfUnaPWTAeeBwT0iSQqU58BPH2ZT/0U9dRiexTpzWbQmDVV4IztdgYqOCpW6sZ81F+nv1qMIitG
opOFrO+hW6WnVdf2OB/SS04qnrFnW2NEtBfAF3SOw3TNXPbEWHc5BDgzIBbzr7q+L4GvaPNIBOfQ
iKTmiLzSD0ALen3GsVnJQQfoSlTo219xv1EQvuIninuhE1Sntycrn/TULdrICI8wFuHTwOOBTPa4
6J8yNWDQSrN2m0C4PEqPHL5FQOn1O9m17ZjsEiOLE5gEEe5liVGp+JQnVBi9ITTpK+eUSg4DoKL6
tMBCQZVsNrTO8ioPKjxFlbsfBqpeDk1b/n3l5lOPcR6TEzHzUpXtLvNBPemqcEJG5AZQ13u0YRVF
mVjXShBTqCmVRZhDUyMLOeFJxV68a+fLgaGPrikAxABosTGUCyuQ1tkNFnmjlrAKtXzvSdNewwmK
7lLCEK+gOHbvGX1U0OEWZfkjEHQcc8LZy3KTFvvg41i1h73otHHoKUbfr09BeVcoNAINT54JaBFu
GlKJD0i5pWvJSY3Af4CvK89/ytoqxvnwAFLjeodWk5KXD9HlIRHOuR+9UmKzvrfCHArgJwRLRCid
KsbpxHLNV/CdPodLcsnT28vBjejYTYdFpmfzYkl9FE62I+C78l7JlBxtPe+TbjHxl9pXmtGWK+sM
80tIQXwtmYH1E2ks6GpRZgwsd/Q5sY5uwcMS4V2SpwTtck21OqtYY2VITxVVf9rLzW2tIcMHgR4/
jVhu3xAEOWG8TSsb1fCjsE1C2KiVCJF6t2XPXqQg/jGBT12frP/zw+7y9IQ+/PLzGCDmD8UlVsq1
Tb+SDhPhYhaGlaEkOW/7U6nysABL722FaMhiDu7kqjC4bfC2mqXF+W/SmNfNT0FyhEsTATBF9IUX
6mQPfzeafrsPYqO9LU3q5QzgeJKeHPvFXZAeiOaYSzORnKmZEX1/SMwTA5A3GWQsELaquX2PazUQ
+GSQYcCAlMfeglqWnb5nmHVajrdxunXubuTD5ryww5gqXy1o4rlTPWBhgMsJ/i9ndOu0O1vIYmOS
oXJXPRLRk5mriblFno1cSFl4I1/6DK3YzkzZTt56OTCyt/t0pzRq8tvHg3vr/8CA5vzfvgOcPzEC
uyyM0t8qgdH8Jnn8olDa4g0hZOaDWnbQ7zlDtBqRXTAOQkCa4PvLsso72rubf3Xx1TG414xkmBni
IdnpZroL51AT2zrd57jC+TWK1VhRLRw7MjVwgCDcqWon1/5hCj5B7iQOSBrT1R1mFxa6ERODXgx5
pZd/adpgh1ZExVLk2Zjn4+hinCKdr9qxRTpPB1tIg1Opv6bEY75xY2HtSa9kIJfhzKoVlrRE23K8
z2rsBRDivS0bTB9d8ciNejCgtjDK6fvaarfgF6RsWO+y+1vhvzLwsqgqU1uaK9aYxCsXQKZokONq
Gy/bhJjJWN0nNSkNMvHMmgY3EA+7IDbMKVysJKOEQyvqjZIOBtz3UfU6oXwlWQ+jGvzWeEdR17wI
PvOgJ0e3ypdLc0+fi0quFlL8qXIG0J7Galv64ToQxlho7AFLioGG95ptS8fZqSWxNU1DDFQQylUd
qeuxgVO9TFnU4P7RZ2lUQ1JG3zATE/Y0fOu/4D/uoTV2jIEkwErrR48DMXf5q6itRgARqOQKPCO2
obSs6vClHqBgt8zsddipT9/7o/QMzJW9uYVtOVTFbp6Vah9AME7Dp0tNxPqxJY0Kw9IYoCHCmsQf
Pm3FWDWjamFuYarFWC/KSWf4R+Y4/n7m74oiKHcJ7mdU96sm3zVEDCpzmerszbpMPiDSbxGIXBno
OH4ElNkzQA8qrwjssDDcEmVlDDa8KrEoLxmVYwMZn3xHJYN/gtLZeSf9hX+71ChePKJd/13vf2q7
yJpdqPTkYsy1vsGQ/YC5Ss0WEjbc7HnhwvF8995Wz9dSqYb3ELoPvcOOhHIj5qa9NmaJm9kuk9Zf
kx43odsX2plugEQ40hAjV5VoCVPFbP8mpCN/8zekqnhbZNNVyQM0PLyr6RfCulr3Xe+2EBqsC8tB
0F2xwAr73htgN2aOGoN/vMfh/VX5eiZLa3WmQCkTafWMuLgql7DJ/5wK/eFpM5//bXgWHzVXUOiB
L1sn9LbXunbozoxgwaPnsRNmMLbJROHTnt/83NOz/mcyfe2cudtJsNtLn4x3Wd06ZXuua98Qq+HJ
/y5wHr0apYeKrNUfXCYd96mP1xmrjwUZJZ7s004LrJGGTAKdPG8CZ4ZrYKEOwUXokE0DynBq7GZV
mC/QeIb1Bphoqbo5txtk0DBiBsrO1KlbsNuEv6wlRfPxG1qNQIyG0zikDoOeQ43XzzQ2lxz/bdV9
lsyt4ouqxNh3flN+ME4p0cyyRTkSfVfpket4REJJpJ+VZmWy+UEnCyeTkPXTDYevZuq2NTWhqJ0T
ENQnww7giU4/EnSynoKrXdIJuVj5ZSl3mk0U2FCo3R22I7ANmsgH3Fw8q6nMWYUnczl57NKAxXSh
oF7a0/lz1jTZFd5B7MKmK30rfykicQrRrrKqYbt89MVupPbR95wNgcmWSNS+xuPk5WOZV+BNmhCB
+Rdf3sQQUjatvNL7ZGtlDXf52EA83BJgnh6VYDxSu5ns/x5iCRrGOJTIEV2Fe4I5kISCeAKOEbVW
bejnJvBc4hriNXzCS4zCobGoyIBArSgS1kf3dwT+jylvVXsBJbKhrUag86R2F5LoWFk2Sv0xS65s
XOGye3tT48rAEl2SWUEEaVmng9ca0twcIqT9NftEKXUPCDcpJXPQKQuxozGDZvJLmfgcwcSW9hqN
4+q/B+ary6flYKcJwC8G84zWF6lYzRwaysj8LQ+P7nIS12fpUJSXIpIvcVt0tMGgRtV3eAhB+aay
BnK1JNLCcdmu33L78ELA/Pq+TrTEKBGxF7xdBbgxYa5xinn+u0K0+f3+xjwkvTo5R1mmi+U7B+Ur
FY/OVdJpqvKA/sH+e+NWtm0J4EQWzWoutmKc3pWoKgr2DPNO+QGkbE/RxcPyuXGg77x0qQJRH9pn
WRmIxH+ct5Dw3RETngFksIrPjTyaWxVhvjHj97iOQzuJcDnUNnwqLuwPSCtdPeB5hiTzfPPG2dYN
MCTP+EFbhQCame2va4KKbQvOrZnFSi/IVbsxaI8yexNe6Z0jiIjhjKbzp7h+zU/ADCyk2lwSZSLR
Ev5HbZ3cyN/eZouaPOCwPLnf6BmXwSSG5w/cXsXWh54N1KSCQmtxQSeV6MD3+Jlappeg9fU9+OVr
0y06fl0SIiAuZh5SByNRfLa1jbKNyJ/6hee04ffIVXpDmPyPezylRtAuA+arHNyEJcQp74YfS1VE
/iZsfMsgIlW7Y8XrG75ZKqJBodLyd6EFaMrKz7zEYqClThMMEV02raq/mfm5zaZfRjuPSTpjmE5Q
flwwVacP6ICaQuA9BuIe3jcy9MR5tq/4tVf5zO6n0NFzv+w0IIDpU2CJsv5Em2f3Lcx7YZ/inumZ
Sy3s2Sda9YK4gmYElInaMeRh2ntXwKl9aApzKTP10nzbphyi5G8IC854S6AHWbEFEmqaoe0+6F7Z
D4Mr4cPcPaIQBUyubdIGh6Knsl8aIZIgVI2o2RTPTJKJA0N4W3DyUfgkFKAxs6vKlRszHeyBw999
AdtPs4cTswBvhumifFEGaXYpJX1So2f09Gia/kTfCakvZwXwi41/RjC1NkGCEt40I1KRPIX/wcHh
FfJbWCqHE/ZsE6BcZEFBjjNU1MsxtXhHBL6mCAUDeUztlUBLUdjQqOxE9EpSiO7PIJy5TRenHHwh
V5qwpJQh4INtNBPP1/CJrvQCZzAXd3SduQaB4D98HPpDPBFEq5U+SNbuhsjichyK0rvRXUX/Hyyw
tFawe7aV6iLKL/GqCx/m7h3hW7ptRROhzidKgGevJVZZmGMgB/buAsfmg7wvCgcQ+Isd3qJmVrX7
+GaMHb4tmxqUVc4PisQbkBVrwb6YXpLWFRjnzqi/MhlJd+3XvNZ1a0U9GhL2klxKH9XTzt5TlyV5
U7Whq+lzVjM4sPauiYznsLObyaE0ugLZ0ORTTLvR1qBBIfEVlYaxb4M8GU3u3yXj/oZq5JhJJk5K
Paz0J84nAnzBlj+0sy9Y4nWQSRYUlcmps3cAiOtgX3jIWSkUQgIaiHGWkeA+qWK+bwtJoiTir+AL
gvXjYqXI1fYH/hdxbHcQJQTiIWvO1DoIc9HQqM0T9RrMwi9ChVnL7nuq7ewD68u5BuoVCjBQnCNw
o+zvRiCtqNAeyFIFB9E7HVXygvTYApfM6OVHEIGZCuAaaW4pQPU2Q4MGnfCaGBsklBoj93mhmcKe
UQiL8eEE6EU+iCDQM9LHN6OEymVJ70nPQcuiDKYrEkPfT8gC92mfpxS7vcRq5YIlmLsuTgb9HAl5
8NSiDzQIk83vJzBHTgu2FgeOemHkVYP6e2H8ss9iHc3o9e/AUaHBLGpmX3rgE1zRgPfnf0vz6JnG
ZgHhbEceTde8o62C0V6V+8vV5zb5Xgl69Raixtzh/ml1Bj17ENB2jaCBf7OmBQ6oRuKWBgTheNPA
7dRehE07inHMeFkNmZLt/icWByLB1MO7bF175E5uJt51wgj3Hn7rdcOhK/Ge+s95v+O/x8oAAcuB
jEwZcI6nP9lFbv0k4uCBoSYJebd/kWpHNTyZe5fu4z2hjsloJsTPTmApDa73HSWbFjcYgPyh4DOy
LfSKi8Ftdrd5yh/HD3fryp8A/5uoRikLFmt+c/reQGfQBjQrmnYTHbuZ0P4NYW5ybRzBL0HX0jFP
BAkLmHFkvXu+GbD/VCHKSWAwmL9dWOGvviIiDasB30Q/UlxAKnOSyd2UIS4jueRZHeIJBJ6vs1jU
PGYqHh2wDXpjgZL/+x9bmOUbw6ARhdCvkc7BN/wzYto2R/gFQe6TD8alBqhOMucMJXhpjKuHRBY4
QVEFey24GVckAuwfudn2SEWSdCic01D2h4JY1jk8gLlNcNdjTxn4quRyBV6mNbRqLx2rNJ+WAYSu
65AugpDaN6le4YvnA4ROlI2QWChe7Ifl4tyVLVObRbNpcXTPT6lPCTkh0aL2CL64FLhY2dWCc/un
WHScGT0bTGOHveQ8ELSJjdxlJ6GxPCBNb7wuPsKYNDZp7irB2+boRhqL1U4wNV8M1BsStWPqPqrx
x/dEf8E29dwcEgchR94nDKqGFQeuoNoVoceeYvVh4+QCy1/ZsTaemrfifrqTSe0hIz/pjqeFzZVL
fTtzszLY9GlX+JjJgPp6SoqT3Np5AwJhu6lxt2Ls28EYlihHYDI7bqHi8ZEscLyJxLizhLDKsOpI
XYJSddKbdbxFJ6bqppKQIQSVSPFSWO1T1Q2oeSF5G+jsr9Upza+pdDiVgWZ2CRVXSuC0uFbhKBzP
PVGo3dF0v49cDo8/HzVaGZhA/pURsuy/AKnOy3XyLSQ9vy4h3ftakXhYyHATc2tE88fh5INks5UJ
HKvtnJEMFafZAeak299kF6e6CwF0lCq9XBm0t14/ppYOvvcflxYvKItwfXVuGoBYFi7biLT5QKcJ
OfCFzWTFvuDor6/P0/91lTeqkA19ZVOmB8e8/yPG9KkDIabmZjkh7IlaitHQu2K8/cPiM7wdR+tX
h0CH3GlOu1sBcpx3NIf5hDT60Y9JT+hXIAXBm/j5PqHaHrZIwF5e+HmlcZ12ehkfPvCOHtWMdaJo
JKT8W/Ol3aWTIX5vgIzCMAYUjiAKQLmjN1k3XFk6fCG8SJKIgnKbzwykIMWBJqGjRNLK8BkC3gnz
S1Dnu+oKO8krMWbF4L5yynw0+DCRBhpzpg93hv9fGlOs85oSxeNPqYrrqVqoBs/yGpkGVLO5euWv
9pgI5gz3qpWlwkGtpuey7waNQ1Fw3OjWn5t3eGjbNibZrQVfQys4IRDpEbAARIL9Tj0Ux28QiAdv
ZAyXJr6XagOolcbHQybPxENyPIRNZ21I2Pu/fxWTG2WLNMhoAVNcnahG30pPJF+1UbWdJCwgs3F6
Q510ZdagMBYghtBxpwIAp06ZgKQDHPigtONM+fdlvyKull5iJ5sl8jukuyWBsdW/nKl6wc8G1uQe
6g4wXqOH8s+9QwFytbUMvsE5PFMACqEEXEJ4CzM0h88qEh7127pCwpHrg7dAweFiDV+obmFk6dmU
PuuIi6CcrbsPR0LVWjZpcMRsPujX086cctL9S9euFHLkCSMwgDw4QuGk7rYOmrl1hqgbrq0ihu2l
d3lezeAdb1PgOaZ2W1vCk9DghpTimknZDMZDqRZ/6KVT/yGXIBKAdC3Pqt6rdqKLit1Kx3/TSlbs
24ArDaotlYmOrsZnDBSj6wByJcZ3GwPBY3/84EhkwLGpG/2//6P4FOYuV3NwQqxFLizH7CwB9ixA
IFh3Ofi4b3IZSK8zXboQAl/Jhr5HwV0DNg2X2ZhwOtUALmeyCWL75LF6CdrkoezcyDU/xbIImw2S
9Ikd9LbRzp8eRZCn+Bt3yoZmvgnF5pI08IZ7q7QPmGcMUuJZsDgXb9q+YNV8i6Xzf5/eEYGrI75r
j+5sn67NYjMDca1LuiE5vgnjdkH9DbnDjsm+7slvPz7CVMkVHLVKXASBthkx93GfhmNpQ9r5VZpL
bC4ie8NlW5JDqp6CmmvHBgIN+PMF7yEThGLY+tYQqfaFLY1/WBz809PKUhE07dA+WH+mECeUrhaA
HyOyCTgDoyba9nKgpoIvQm+YG8yY05MEu2wBp11ReACAWRK+lU96G424nxqnwN3BdRUYMIPeQVCl
w4FL5aiXshCiD2uaNPOWOJ6p83cd003Pzvd0dvjC0Q4JnIuIQUa9NtIrdis6mJ4PkMyCo3BhnTwA
9K1aWi185kNseMuT7mT1hUMZRhbY4LxlCKE/LH5KgMKCReLYrDWSeyA6wgo9tMcwYJVfN/GUrF0t
tPl0sAmnsrCAqBv1EB1rjbwN0aeo2iCzaucKEn2hKVuPF62m/8FyfYw+ivYjsdPXjbn+sAajTcBX
ZVeXkB87yVJXHoCPuDLaCTkrhldT5m8zGjWfN2L3kLtx7Kuy/Z/5CL2KmXEd8cwg2IGIU/uvUXie
G8g9yV5t5i+wRNrriurbwhsRwf96ywEUAHZaEbIdVKnDX+Epn0hxAoMi2xx3GGGxg5Q7F0mPQNDm
03IpRKE0sox2YW4H9LE5ijG0VYHdmEux/EHlXFPSplzSPfzn+/mj/i9UO7UYMzb5BMq3b6EwyZtl
vYaHoSWvYCikA6XegEdohsXmcpg3d3nU1y9+f0SdlUj81Pi9+7UOD1wGqKyXsFi0FduuZjv6Q7RV
7dq6FG/vRRgZcXq3yBABtdhlHMTLU9RrlCvz169t7yzZS1pCL2HMMET8lay1raUC0HGhQhbp/JOw
bfR6x9tnllOvQY0774G8KlHW3poWv1JgEh+NiuyFHEp1wa9mp0SVkw+fYJ9762/Mmn95Wk6WcIfS
kpUGpz805GfeLja44EcputcD53Tg5nUDGBN/7fY5Pu05NNc0mkCevXqliFde05L091c/ji4ev6TT
xihBpGpMyIRyi8OsH/SSm/2NZcVbDnTU6g3V1+5eWqgwrKz87EK0KDLOsZyKmDUYjh8pblqP03wG
7m6yFeVrioq/f1nY/aEj2Ci4j+qhtofFqbb5TdToNcalBRUsgqzyI2W4Exljh30lIVfbvpF5uzHL
UsObs1Hz6KNu/UAW9o7+EidvT17vJnaSnjZHyIIOi/uDTndS2ERVRAgcCks60ongI4JApjiagAzC
V5qF3A6JlCxeg2dpI1rwBdYTnA7CHw6gmi2WvcgCbfAgtYF3BdRlR/HCcaoj0ZgkogqNmQXOfeII
/EPttgDc3OCbnvHS7yDcpr7FrYeLWIKHp8KnZ6YRm8pWXMMiDGL0SSmTLWnBr1lFWkpmfuItpYEl
HYnLcaIX/+7o3kGjXNKP6mHYUJ4u7xm1ECHOsTTLxD4vXcGxeWSH4w+Mq4e9RAnr0OhBlLrRJLQz
dHjya8/GkuoC4uL865FP2WO7vWZ9BI/i6e6cUcWBwG6JOF+BKdZt1QugO+2o15sRd5yKlViVA9Nm
mRsqKr8GEyTOvy3VEnwg2ZPUi/jC8+mKYgnVl5YejStSBsQ/MiFzf3qlym6u69vHHI1ilY4PBlNn
dWZsn01l93KDG456AOqmxg+llM0q/Nov+IhPDSwnIlb4o7pNVFOXBLpCje6NCeW4xAjBRxBhyHFe
4WEVz3R/5XPJ9pSbi6BaZMXfiyvv/NOJuCMc5hWmTyeqZcQUU6fDtSddPvo5hs9vqNkfyJ0YLwe8
qOAZENC0KPmK254kjH/rkEo6TRGzpOFHCQvys/4GypP0sAhCUyi0HP3PupzjZcNgSVLN9WlO1QPA
LHY3iusCOk0ny6fmXBsktRe+SYta4jil1OuZzeByyufa9BLlRBD+Ke7/geDjs3Y4zECi5A9EJnSM
SoAPDMfP7jBiBPuWMH7rDFAEnqbLvj5pNrKzmRacyeuRpzQM5pQ1rQsv49lYdWgaNqYHqIzUzILA
XQ2iF515cl7JWp7eR5UJihItkq8TaigkWxaA0RceA0eBlQEoawaA9H7Arem22qSv00wWg3QeY7Y1
mA/MBRi57U4SqBx/AzGh0V8QYoVBxBozAZ4JWyx4jL1VDvWuaHD235zL3ThQV2r21aG37j1KO9EY
tTQM0hj+CsTeEb1MvZIhQanZakmol977G1wy8nh0LKFcB3ltj5PUwePpKRmzspiIF7wGccCM7P9B
44+ec0A8O5JVSV7RM2lMPObYhrHC2FmKQDUGLTsDcKHmqLExQfcq+b9nq0rHrm9cb9lqWF6PlEQK
avJtfvmeh3aUu5EeLebjF6W37tEHpaZLUb3itwLpyn7d2IvRJdvIN6YOADrMG83lD2J6xG/Mcqrm
s7nMAiNVxxXX4YNLqMZr2klg6CKMQa4XtJCewI2VNdBrTHmZwopPt/M4x41vkankcSYoQXvs4/MK
1RfG/f8fER9Ih59Yk015s/zu3AHA7EI9fnzGyQyDVtLVvNz/c/0YI61dmuhF/jY8Cq+ZYM3S7Dnh
2SgYqC9CEcbn24UszAks4xVaC1dh5wTmrqagwGYD11WYGDAYhBojuREISFGHX73Jsjrp4d++2bDX
kCJ5fYouwICX6wFveUlhwzN+HX3eXXFlpC4Pup0RXr6wv1Q1vGlQzDriOsBgb+5i55xGHpU6HkUO
ccsmV0c7ddnNbL7SBWGy1O06CzV1RoGGdzRcFoUrr4efPfSAiCDqRcPuH3eAoxsy5TFnBVc3b4Nk
skGwqfBHhf9hfCEHF9G6Ge9UnOeDplXql4/K26W7vkmy4Rpx8twlvupkwz0sbC81+umGMGAUekd3
SomwRVwp7b8fKAyJ3a/wJQKTNrXUk0hhwReXTQOS9Yk0cREduObnGGbiqkDneNhZXNlI5BHu6nM6
wQZQpyYnBuGjnFvetXQVxukSsXtVfK06TPiIZEWJUna/65ErquSLpuVx9JJ74NrOSGmHuhmUnRlz
enbkyyGQhQUgDcSwdKnEh9UBuw6pN4X6kHf9yY/D03ty944N6na0P9iQK976qKlyJ0PA7QHtO3KA
sPD80RsfSl/bMXO0FY9wtZYEtQEKONZ+sTut8sZ3NgNeSfttMKIlyRGSv1g5QV3CXB9y1LoA6zPD
+yr8qeBLPkySu9LuxaGlLPs7XyJBS1Aivb8uMW+6FgwxhgVw7oamCO/qBWlUm8Pu7Y8ApkmlFxpe
0bVv1tahhTBg10bIzb1hm+SXxMfkANZGDrHNedEe3WLt4qZNLpgZryrNc5fslvVE2j5BX8QOz5s0
r1G6ZNw9k6vd6524V2OEzYElqegwcCCqjEpJSiAguIkgRSCKpsT3/0WaKRIPHCQvcV++FfgBT9Jj
tbse/b3wrFDSQcca4ewz9o5mWg5vHsf+KjGeTk2yxdWWQcuaWaZ0xrgmOA/gbZxU/op96GjKD1SR
DwkOO4jGupebu27TlD43gzPBW6CpaWrloRcS8BRZldUYniqj6Gbvtjyl7JVNsjJE8NIg1WYhAts5
RfsfMSVekDG6JrKx9bGRnDVjfcAhoTKRKUjd1kDykcMzhb7uqhJ6PDFDnEvjU2VQmCxXd0pEqQEw
vN1NAJU4YiHjpcHOjkXjkhgZjaTexi2Cy5mfKrofw7PYP3MnuGC0UGHJU7wMR/24sFZMGH1BWfJ+
q/qRvImJMbha30/YGvh04Zc5y+mcsvjxmJjSQpocEvKAwGhDNR45raJfuZbxH9X5ETgvejlFwyEU
MbEsrH9OpXbDmrcUSzG4XCyv3uv0q6YoZy6bsTTXSGllPqFhxNYFYkRhZ4ooynht3PdH55PFNimF
5cVlYm8z3qoskjReCCyzDMk+BJBeKEvBDy/wSCozq9WXs6aZS29mmSgaM4VkRykv6/vVJSkuFetX
8BxNRv/761LBfln6TfRpaxXmrriJrzLpGURvbcTSdUcWj4xt6v6mGwC9FtD12DY1dHNCYEysGw5E
0Z2298qMQcYEmfEcNrs9bmfDynKwuvRp9cTA4/7bFMUEzbusP57DgtnddqWLQ9cOWGyJXCHq/jEI
rlyuuVzU4pwtkfirhiQ3nbfRKUpbyaWUXHRZmob/d0XBopl4bMVxo6AORlWj0Xy8Xe3YrLnCQ9Z3
1QWKxIhY6hsHzFs2HiKsG9DA/WFamk315ut5hbUNyl6W23Tk5PoNKia26bhXHwtqULG0NdgODell
tS0FklBpTqUqSLYUpypdLbd1WBwb6N2k2ho/hDf+sLEm4DbmrUYepaM2cptFU82sqZg4R6xXmNeZ
4EP8Hu5CQbSb4DD1UOLdHfpGoRScI0TOq0dbvTDXfXrVPT6Cc4y1PqjJrNRM14eqgepiiRGyCm4z
gca2zBLK6uNkEVyDjMVUg4fTHOutdDqkn+jBZLKp/YBgiWVRWav+9vw7q55k+P/NihCpaVp71DjR
gidwFDtmocPt5Mijol1tbMLWeeCW6vLIFapkDzKxrLlAogVckxySpj/OT6ZhOBsyO68gSyB29N8/
o1GC39k+EwMxttzT/0ONDi35aX5+2pAU1pK//qfTCNipy89RMy6dMR9y1rRgjvn7hbeuaGXxcQKE
Opaema4SCWBbRJGwI6GvBfNJQ3N9WrJ06EeMGhjdUOKtYgdpYz+VdlaTI6SHs8fBXxTu5wl6J1ey
JsZb/wwBS+GIphXts0XI/GbPAx5/xqbaf3d8aqMK5VkIFtkX5IEIme5CLpf7bDTYZNBqonOlEWZR
I7pnJgL2rCM9uUG7rovO2yltUNB5sytOLRBK2H/u2IHY1wlNreG7H7ZBBzyIXcuUURheqRjIIpy4
7vpdUVBwUmzdEHGFhBWyUSu51kMpmmTdgCXq7M+IG6qKpQbw3TQvuoiyDNF3OOM/FgUYatx6su8C
PuSdu564Y5Q8u7xlSi8uFCm9q95pat+laDGFMLman/y2GX7bng7zXVsEpNKTsDB4pmww/cZP7KlX
hDqkoRDcQ4wombvW4OU5jypAW+NpDTyYx+80sQLqYIPYQeqsGD1vVo88QS6VAubvubZf/Qsr3wlq
RjbBOA0RiaaXjvqjclkDJ+yqncUSCzDC1syit0IzdBWV3si4727AKw5qvjclr8rquCeWK/d7A8bN
y4w6Lev1nJR2mlF/pFI9C3Z/DFC3kSYjkDOltgSlI9DTupIC43Lby7OW3IKqOMV8S02vOL/asV2C
+oDRVF5xTzVKosy4FdtAlFdgIkUxh0Vnj8p0N1rLjdQN5qSf3g8sIHuNeNExpvVvS0rzbpXHO/OI
BRR4QaFQvZkZmWqiSpOURRhzVslhZKLOTB/woQaQRizC0AMmreBZSgQfV6py+78P6SEkoAbxfATQ
ynczqAeQ7++d2XSWWsdj4v7whqsreuLXZtsLEGbPGYpsvdUQFmuJM7K2cAmifH3tJSvIIegqsgBs
w7ElT7gKyTkHRRc/at5eyjXpICCgXHk9PoquIy+kS/hB7GjmcBwt8FbpLhW70ikdeC2UL9PW6IAT
yFG6wZMCqcc1nqIGWM8G4/Xyzmlux2kib6KaZn69wrcrTOUdmXLFfy0zjsgS/PwRV/GZ/a9jkztR
W/qxVXJCUqxIQ9YpmhCmgHJSWArRU8kDMLOuqH3Ui3kXW7mppOpcPk+gk+nYLS7beeDKQ6VQps5Y
ONMBJBp8R90BapRYXBYMGpqstGA8nrkjiiNP628uorTXr2R1Au5wM2++Zfewd0OLkyTsIuN5Ti5m
jZU6oRyeNsLyjnSpL/BOzgTgjXtn4OePcb8ybplJxysrenJkD684a3abJX3Xg0k7qGvpXh0JzEfu
1HkH+nAspNMjWqsTcnCYiXVMIZNdCAjSXfswTFBhkLkRP1XcEl2qMVuc7HLVN9REAq8WZoy+MUp2
l3Pf3j6EhrJy5RTvY4quVXPceO/nyBm2p6JuXnY0Tur0fCbQmjEVnTQZ7ykPnxhf6KfNNZ0oKyxA
BhJun4KJb0kegtHnYzxdg2C4l+JaJYkJZud4/U2ZUhN19vbnDnpqfuPKB1vk/4i/AEB2MLQY3Bww
eFD8Gzj8Bv4QGLL72rASK89M9qgip3VnUNwB6T+hfFfI6YoWh0QaWXYr/XKicrOEWAN6imjMNlpr
BLVJNnoFWkQYj1Nvb7Fi5/RAHGYjlsEMJaJoAV79IsVKWrkHyTwJvtP4wzaPrRkDzH6P+hiiJxIP
eZETeSZrbRAl+ttis+y9wP/U9cJZgTE2xKiO6I/0r6Vg7hhWTPPrmqk5jVr4R7gkYYBEi6kFf0qv
kNkcTXeqCuNg2WrSs2uf594M2Xy25oVWd4mEizN9PLTc6BdBZ6jDF8abaKV1XWRCJzj7+mCcmP4l
YGAym/TKAztD0WrTI7HnQ1/HxKMH3xYJ+oFXR1cjasa+u07LpEvrE6IkU4xVkWZHOmMFgp51M45v
wAs026SNoFx8+aG/AoWVs3Cweu+7wmUqLuecYRMgpszKeU/bc9YqRA9PbJfOI7IlIBTRzLZIgkrx
3wEd7R0NlqkKOW5QvR5dv2NyfZH8vIIMAr/SETgJ4cesJbAxtl7AhrBBKU8XKYz1VpHZ6gaEr6ew
lTfkAOYEkv/IN87gRax+zTV5AqaltbMh2GRO+KkkWM/BwYR8vJU0LCnJTlzw3CpxWj/xRsk318i8
XmInCV/WJbyULMYzRkSm0Oi7ozcgTP0zS6z9eu0GqkNTOcFCNvqnDddEkrFrv8lzK50IHnp/nopV
8S0S0Uk/D4u4O3VBe6QOyodsvjIFrXS8ZWJMrNnf3+YKpabBIoDHDBGuIw59QTVPcRdR+R2qhS8L
Ir8Mer7AXR5ZcSAPfEXf+GXBjg9VjHWfSnUQKIKqbgB1Pc+9ZESw2aHd1+78sPitju/XcEAF+EjM
ZAIqDpHHpIvtfuShQtEAo7AjHb9qQ349+jpSP5onmQ7v5shTCTO99BskIf3T09uY6RX/5Yk6N9uf
vbkkM2wvBtmds2e7frcoPAM1rEYFNaVYXijBpxYC16v9nmf38j14b2BS3C0SMQiAdbVIry+xZyEM
0YWbADixBY7m6hh67Vz6dUxEMUmoQawDcqDSwt0emq+q29saEhS3+4K9VL5RdJ0SdMHqKC1IJtFm
t3Kt9353mC4m5PxE2ndA4MEuH62F5rMSF3LINdc4i/A5vN8w/17p+wn96HCyLrF0+j/M0lz/OVlg
Pyd7j6FH7fYOmeEMaICciAiFeDaK8hXfRZc4RHwIZED+bs4RQsOPWzHpJ/VgK7zsupsjsy4NyVeD
NgyNfVB6x5pUOUxA159TMytjxM3jgLpfW7wa7d/Wex4T6+lOZoQWrstZqN6+/5E+NZYDyQMh8AQU
sal/Q72/3wOzjyOfqGl06THA75IJG8825bDt7paHm3H6zYr3uzTftTbcgcefAnvKhgs8aN94zAtP
WPReK4wllMD/q08ySujfEXvsS+5yF8QODu4oJCX5SqWbRoKEPYIK+2uKqqmH5zOQLXdqQLcmk433
J+KWQ5rX73KzXJ97g0At8NFhkryQXuGUqL9FM5BGuaVIHbNmyjS/h87ditECFkoBUeHL8AQKLHSY
I/s42qWGL/FSA/QEib+i+RUi7bchos/3VaCOx4YyjiAnpVExAdqFJzTr6sKkgVcSvMIeHGvfknn8
LqMB1+cLD+Pl4H0fGJIk2hjquzGl6jRnuI02Xw4VnXpBKhj4tSH5QIzjc6xmHFywUYMYTiIBKWdh
GiSw3NqLF0Y+mhXTv2+AIUVZx6WgKbWrwOMzSEDqPNqU5JDoo/py2YPJvbS85IsEWOtM3O6grHoJ
FQnxjIO56SbQZTz+5oQndQOa0gABKagTaJ6IPScHJyD72fybMGHaveiOxqbqdnPeLoRhSR5oVUw/
H2D4WBfuHl11jyNvEBKppzMFmxQOGg35M6XWWgUOiS1Y+fTMYmZWV1KdL5Wh0jpwv7a3IeihSqXu
HOdaaJksuZMTl4mlmUfbPkwnoanb5nbH8+54MHyZyGl7SqEZIWGRXAeT6cZOGOoKZaa6wYBGk0QE
JFdfOK/BagVoE6Xp9Qi+FR2lwPhxiIZhATE/a5o3N61Zv+0BfidTvWoEjuMagllgWAB/7ZYe6qFz
kj+tK3lBrq+ZgdU/hGRwsQUSMZLaqFXUAyT4a2vV1JfPOqsrfSyLJTCf2g7R6P9OJSYjp6hOvS/P
k6WSRJLOFaOAgcLVvgYKc+bD9hZLhiYDuATRHVJtbiA2LMCl7HP9NuoYRxuvBJGkW3m6oWiTYL69
bXbA2FI2qzXgP0PFOc6kLEYbbJl4IXiZFAPrIJSlAO/M/FDfrxJtzIOc/hCMZrkMA3zVNKWyGu2f
yjJrAUmlUlMeE/6w7vnnn4SsMYalhNaozeFlJqGMT6TgBlWHoS3M66BG9Vjw6kN7O3/V+4drRVq7
gLEXwcEYnj6WQD4YIxRnOw3AC33TwWRmMLVN5PUVrScngY5CYRmpAmVbRKchETBIt1ngO9q9MoKV
sMNmOfmZSKq5+5RPewDTbJtvZX2eApO/roskJv2RXQ6KeW5VrQ0ij9ZQHagmKntmOdlKbRtPtA49
89kWdCGQIG91vdfD22KYfu2I12VGaF1KSyN9tvTg+nfR5I5oco4Ib9XwXPKJpWVqAvLs1GeBPQqH
2KZik/dFSQccID04IpWmYSMkmtWlj/mf7HCyszMZsEHvnriuDpdG3tj1jAjjn+QD+RcE+Ckd+/8U
XFaMpXO+9CqPSVuTJpVMR6lntoLZyrLqhimEjEEmcP+8H5pX1BHcLIiJBdncZlGxd4KcXdZtax6p
gIzqGrCDQUhZh1g12L+tRwGKY/KDALaFaoJiCf6TlLDiQVwq5gIhLpZY1iwDg20qiuQApk8JVY6/
FKnIB1r23XsUeRU5m7tKLKyGOleB8o2YwZg2aGvVz6zPV9bly+HqrM1JSPT5WPiOCPQ0Ycgh5/9+
l8TAUbKYNPe7p/EtkVCcfXt0JnX7C2tLzfyFQB6HxxRtMSlFG77JORDvZzlENOC7xckWsx5KW96F
D61Kd+s+jfKsVSbHBbKRUH4WvNJrqjXuHPb0XybLBLu3bHLFsuI13LgKO9IqlL2HRyhXIpi1TRFH
MDr9GnQCiMAL3+Hd01h8CyVhlp6wK/jl28NvBiQ07yLMRy8FWq0VHbsPA+rowvDcSffaSldHMJ46
6CMR8/2AWyNJK2WnVt7t0HMeRCWwG1TXAMDQ9IS3q9Z/iPbQ79s1jrpDcNHMfU9Dyu+ovN/SMhGt
XDQzltQrzjTFRr1ZsrPwFQkTEOvjuRcYZKhUVg2qwBV29PDofdmwA6i8D/gayjPhmmi5eve42zzr
tI6UdLuQz003ioX/o2LW8oZZHOeIADT29UbEwGnrftwYP3DHo8CD5V9VRGDI1uy5bKHM6KkdVRzm
+4moX16uhlxaXLMTFAP8qDfoWCMP30fGpYkisiMF0A3etZ/6tyBqf9FgpVf6t3kC2maKSTC60Oxs
bYbtwSS/jaCTVHo58qF20NmTt8grErkIF3OchbPsFT7uBpMIhTyg8px4SpmCHe8CvZsj29/N9D+I
7/knD9rkHkG2rrNrWX56Q3KC8H7jwryqWZcMRu8uRaSz7VRKHu4DaM8mkf1iAhGxedfGN8ew9m3t
QfTfw3H8Gm5euV8/+fbn4P4UdkX1HJG1rVQlqorAwG/DUme0NGJ5cVAKi/u1Bc00/U6OptToZxtz
6EOQ/uW4UWlvWKoRTTkxachYzc5tej+nYo8fql0/Kx1MZvtvSdgyd++X8zqmXqwnrI6hb0sHy56h
Wfl2WmhPS8UN9WQDS/Wi1TYse6564Kvud8YDfsnOaZ55FHSU8mZ3glVbf0FxXkPhHZ1ScOmsBxQA
32D4Na96KFarnYRBLFjwrJA7Ar3LDFsDsM4HDNwPUllAstqmWc7rQ1i1i9+fZI4pxuMOSehG+Q+N
e6dh9EB1MRMIs/lW5fVprzGkk7R0J8qx/0L1ZFFipkOPHQNrQXOCMIk8wDrqLkjvCC40bX9WDL1Y
Z49wVGXkH6NqzB/XvbNK1Vh2Yi+Mo1t6DqHpRWsGKIsZ1+HNq0hNyvkDHCwEHudUDC/9JMQPVWKo
oi6FVI0AHsiZLQIJgMTbGZ/OgWgUmWV42WEgT8fI3mRfEBTkwq3+L3Pgy+Z2ti8HmIS4U3cxPtg8
cCcXuVG3lKBmuqpZjnmDgttl33ZkeuITEmvemWC9YenMCxbLfb+nO6YNum363Yg/jtlZypUo4djL
FGeY2w13Poii29PCh4Wa21AcY0ei9Y6MNAyVY3lKAEGQiYd742QyjWwTQ541Lm3VGx5VkTmHcy2G
rl/ZEcIgNCm2lttOR4C43BKG9j0mSh4b7NUOFxHB5k8zMytanjhlUIHbOtzwHWwcrpi7d9K8FIQU
itDP07LA8awhjQ1SEJPvjk5+XmTlgJAs0jvxWwEtrfbhc3joY5V81EzAT6qRFx9WDNNPjh4hq/oc
0tuJuToDjjdSyDfoy0qLBjj3EXeaDdy4/Ryzry77vaFa37p3N7VlcZz0SNiLPO58N6TI7K2WKjfv
7xVLptH56fUgXn8M2+O/BKafBAsgKP+w1emKFN3bbhBKq+V7tm2eYvtKoaFu1cZfnMVz+rfSq/wk
058kPiJufesAHe6xguVXMfvnuy93mc32XlPpiJ3S8R4fMW+prBk6bzPrcPsaNPdx6oAo4yVWdIGT
PMK8Pv263WsEF5O7VebQL+EQCX18wDZpN6p2Bxy4NWe2/v4+lHfCH4gUwnxlP0bC+RZ9JaeM0l+T
F6Q8QJHm51tLe6ib9ON9VMN+NKE++2rGZNuFNPi7LNPY6XM0q9GL/2x9ziyMUI3ubav7F7B3BXTN
wZ//iqwCO03td0qpJJ/sypx1+j9U1yaJKsM9kMoz1QKu8jJFVSp340hc/UtO8bkOXUBHWLE6lC9W
esuj2b1qMgkazqHMKzUncrCHikrJGju9snI3I4tQtArOfGxbSwuj+L2d+Jzg4ClDOxlthr9bYJtY
jQKNqwUbBXu7iMrqMdP5osMsm/rW24T3MDDoPWYEqu/LOmxj5ZBAMRgflMfV56Xl7wE/1Ywb7o1P
1rvpraIVyBO5fNYuBCW0bZHTkgUKhovjKFFqaP4gWsh3rwNMxlok8DM/qMJ28vKTQ+ZSCfJJvDtj
FFAOCH4HypW3xaXhcQ3fdN59mrJUidisauMmMq09EjKXBc7yFuSv8AF9n083PNyRGePB2KLhFnfC
m0Lp9jBkAosMpasAz0dC7HyPce8xer+rvJMCEze6RA/RUYTl2eFwbBDBsqHIW+JabjtNbeM9Q4Bi
y4kFh0hMR0S557ctkuoWz9dCZ3iH1lTJhvWfAIl8W4VrVssbxbYVbeEo0Zfmbm0aQSkYi+VQS5kJ
Lurarw0VGeqxvIZ3+XQfaLGOI8mYe/SgTGKIwIxOZxQBrJIYBWr7NKhqmKN42o25Td0eBwEtsUsn
OIcWAM2spqMJCds7iZCKdVK5geg5Xp0M4RrVO9yxCMEyRpiikW94ZqJtECnOYBUUvwupnOP75m+k
/6lfCrW9gt1Vsv0bXJ8TtP0zHWC3cKFguS/Apb3cuo4jUCJEvnfO5+F3syEbxPe7kcBIMvUtQ69o
UKFttWRbS8PubqqH5MKwh2MKHE5rixYzi+Hku6JXXsoEhyabpnN/4/MN7ZmqLWvkr532yCBaX1wh
pBFPVPHtGFf7ltl+ctb7QPzVgDtXE/yKLumj+WPDAUIBUPiFrI666IdVhz8CAiFRt0fmy2+au7Qf
j86r6oLAVYk7s+ZbqptEmZ89dE3ezkajBi3nanAWuKF+0aN+B/Wyb9uZgLmM3vFFSBOg9j8ZvaV8
JOEoKh0lBopvsTci9sa4Aal6NOnpFHz85AI1VelGg7hM6/5cDQD0uSPmX7Wg3oUb4WdZD1gOPMvF
vdYsZJjqjkbBtQs6OYK4kTckdXYbkUfZ2G7mr8a2OORzAdBHWffcM0r8fVdml4yBJLHATPjWYMAv
ktt+KA/wovxCqPsVa01CrWpbIaWk7La36vnLK2XD5rc1wSlsVITQ4V4x87d8IZeHlgHFO0HAnzeh
PVKiwLh+aWXYVI2fVPXj6v1w19nBwkujAoJ90gc54mkklILed3jlQZCdhoUgHYR6jVv+zNptFsYT
O6V20olOZto06DfO/N88+YsXiTJ6pEt5Vw6mxU7sqIBcyFRMTu+C8XjXmRbntHld4ZXtHBW6eEQS
iIsbu1DGVu8PQLQ6OHzHQZBwaKkqN6bDjIj2navXKeg/l3w1iaWQVxG7wdzdSmuU7uWHo/E8izpq
70FjKQs+nYHPQEMTGRZG4hM5ykIgtjQSG0YVcu8ao0KcFseSZHV9MYj0Lf5OvDosfqTqWWjMVm+H
71y3RG5lrXAM7bLuzlBFBWtBqdouAjXpNq8Fm9yMO57YhHN3gFdimHOF3rFrG/JKrAD3mgFwtH3X
m7k2dQD8gWx6VWYFf9qrp2DfJNMAR1durApUEsTTazV/tYzAKD2WGakU02t9q6MUk5316qvvD4uM
wrrb8oJLf4HO8j4KMqf4GHsdpl5zmMD04G7qUKei+PHQuSTMzGQ7Im9flfuc1WqPxsLP9ShlzopN
UNnwajd6HWpGrF8MKwIchg79+1ae2mxfS/BjX9LvzzL5/bCQ3AfHHrClzK76pRohdE1LagZy2J4l
kbbsvdG2HBvReClsIjtDz4CSg0UYhCYi9/Qd1cy/F2N/Yn5dyVoW5X21rzok2jZz5BYNwLK4RfCu
NZAlc3Ij/ehJ9MLjz+BoSaCqQyhRVijOch8IKFKCFQ5UDF8hpPz7Xi8GBuABAwa9ZLouN0s6xy3t
Zk10CudOuQCPygFQcPwESPy3fE24tOOuo5DBKHJoyrY67+xcfJE5P45aK6KNS3LXbNhLfruQIKN6
1XWbQQEUkDDvepevxHLwZUjWIaSo/5xMExJyjSh4KqEhj4/QGNjjxZoavyGf32LS+3ccsAT2OkPN
IyHqEj/FJ0sFVbc52kWC2GVPiHRCrxgWSGtDfKpwYJkjSDfBKLn8v+cSlh8IRFy6d9vga3/6eTlL
e2Wr+Iz5T3z/HhH3wrpyw01RC5vBQpIurhWINP+bTe8yl3HH7VB8ichwSOZpZYqeYwbm3fqBnfqA
VTbLv/cmjvb/ofi3wXufEWsqoVoJFtdx3PK70NgyajMsKTl/9OG2U0m53GpwtIK/4qL82L27GAx0
+csxgnpIYwxCv5YcXZVvLLa2S2P6yedmG8CmcoUAYa7w76HwuF6g+CPtkeR4AW5BFsYUkddZlm/T
NgxcchdzmVoCbBo0Q5TLivNEJ2yPRVKMS8argfHLiFpSBchSICHnliIEuIceN/2D5i3w6WJqjc7N
qqTEeP1iu14DihZ99ykTk1AZmQXLXQLU0WCyuEdYWj6EC88oxfYV8wD5cd9WtYxsA5f91S1pc2DN
SKeXk6Dlbpal8tpAsrAmbFrqRKyY4/iVVlpEf+uTa07NO0za3VrxiSy8t93sTfM8jS4RsW2uZ0IY
ZmwNudteIBFPn5lqCJLs/mbg5MZl+Zv5xBNgY0gXmtiLpLlJ7IITrWqAtmXAD2xVtFsdQcyEd0JH
adXs6BmWsbv7vs2Ze/T/7RV1ankzjaI9GmCdg/GxbcEG5mTnMzoxu145QfMRoxkp4eMTlvKaYqhj
UybsrnIj0aWihBOcpd8LPkiOz9qa5Os4xxGzBFLG1ZjiBYTZk3B8a/JFVfHluWfg5n7DhzMcXPoJ
z/NGWDDaz24QEuvAuHyVw57DaKVxkqUOkR3+3TybaU3IY/XzO23Xe8WC0Fq2gxdOlAtfU7QPONRK
sbePK4E2Q6SrU1f22YQ4Z+VV/DtqdbjRLTY7w83os9oG5hFucBRufzqXZKV/4W9NAoBqiQd1jnT8
ny81HuZfeQu+OIq4zm/7IWOOs3yKc+uQKCtRpZfd/11YxpxnveB65YomusLBbPQYI5mJpRN96Ql6
JNWZT7743RpbXS6o5m0fgHPZEg1H4I9VNxM2NRwsF9MC83hpKlnPko05kFqSdz/nsWRfLPiJ2yLj
t0/hKk+MckIO5pHeVDWTy/vgk9FnuWcKxeqagS5tme7NvbbUca9CRgmH7WXlxEWA5iCTzhvZEFdn
7lTcJPFCMC61BNm19cePE2JPR2hOHy9Qo8RbDwDMFaEUmA5Nd+HGHRwVoGjr0ZpGcmRkBUJCtWmu
pkZwp79QUtlR2Z7f0RNR4QsNN519AN8y0xeODyVCOKTIP5EcU45IFnVmoe820i7gjFYbu1AgshyT
z/4mZ2HOQdM4m5A3pYNe38tZaaYNmf2csaZzY4jHs+OLxlUHX+jgRbH1qXveTGpQHZq9OoeIT/Jg
MpbMVsO707CRJg3uYAZfrv0KXqpz4vSpl2lwJR8m8tAs7Gxc88hVUVXWJUgOAl6pcOcz4GlB4s0L
sI5KUuIl6NZO7ahm6wkJ2W3JvdWWsE/e9jM1EHr7ClWFO5PyUAqnSj1sl6WHJhVt3reIrfCBz3HE
zNT3m2Nkr/YxleV7lI4Lpv4RFSuPad5xrUzmDKt3KYSqDNuJdlsybmIJToa8r1ovB0LKNKGdNukk
llcP76jJu9X+DEZyzS3TKiKv7kb6ijtlB471uJNh6bZJihHUNO7ieM3Tt2gSlkrXu/vPH+RlJiSW
giYrOvrwg6nBMQndGCnIbjVtTXH7CNHNyppwH+ajObVNOPEp5ianhbcm0Oimh/CMBiytqr8S7Ezd
pzrxXgv5Xwo8IrBictXmHorWca9+/eee/wxX+SEIPLmI4JQoqDvkXjTUUTXzozZmEZBvyFSTpYq0
ChO4WKsihHA+m80ay4nrXOn8bY8mYfknI/sqRkggvJqhPzP3yPIi0kjk1/UcG9QhxXA0hgSWadpt
rgn8Ago0oUY/KXkc7jba0xA83mNHsQ2liO9nS4KHasujBoc9DE1sUDAys6iO2BDyJsP0qXt293WN
vBvUmMysmBvtqWQFLfRHglRz3ZYG0LHiUqRgnsISeuXiIsPVbFbr9Cagr1XmYIsPdHetALg/T3/6
qTxa43lx1PsqVAeRXxElVAYmRgAjWSm6prrDsvYohbTTjMBV6raS4CgBK+n5zfCi1NeQeNItrPXo
UzZmF1sBAxaLQzHAMScZA+8pSQRAZQX1WqfH8EOrPcNtuLScRp2CPA9VimqLa+k+Vg2azjPMoFMS
77D+4q7pKX9OV1lvC+vfNZEWDCmFh2e8WwbYGrwXxRkrTko1gGtiz6llh6yhg9qeDPV1Gnfvx/U+
NBJgQzfiSA0dPM6G4/CX57gdKY0ojH4nR4F6KoUp04rB9HQywtwFL06NtEzVIrSMS4xehJmPN2T7
ULdYihsXFQsvKEku0gmq17SLpnCkr0fY6mZUndphsci7KubH1eqLOR3fKAJDkXSCdmSP7kA5wBcm
Tc9SaospPou1WXq2HCca0twMVaRA7Jeek6QDUw5aRzZnrkpDID9o9XtL1wtfQWpZ6ug8qOAnoqRs
Aj9+MBAalDYUDDkZKTx5PyvrzxthiWAoDhw+m+YAV9MFGjKT7R00SgRpP+l5ujF5F6jTphRdKgXT
Q4aKYnpmfwbOXO9nHTwX4FQ5ovH98bDVdxyRNR/Duf72jjqDvrYNMFAeUbAse88enDe7siZcUVLo
e0oLZqhE1HrSGmB53du0HmiRdEJJS6WZhw/7cwb7yWMSJZn8G7FCOML8MWmzcDbo62WYj/7zbuQb
lYrRQvRLbtBmJHeJKAYr0JE0hC0CMKRHYFcHwQpCn81M4IqpiqesXn+Jd46UQND4Cdpa7H7cJ5H0
zwwHJC3BXxNcKVsykOApyt4ql4xUshYAoouhBy5fQnImuJGvCY4Eq+n3NEc3RVvQaNbbch3rxKPD
aDNa/Ew7EawglMciJxiRTyfBjKmcUgDijy1NgMvANFtFU7ON0e2Ltv1hVLaDPa2UzaiQgipuxA4f
4p98r4gbzcZGPsvccq4pL9ZAUdTQ0tOmHNJ32QAHmC8NmIMSvVb6Welxy6HbVOJaGRNbyD3eOnLJ
g6HkMuLwbiiChf5fevTghY41vYwwHoWLm/7DsyWGLL6BiYP66XXF4cwNYQcGxNjxcucWpZSz043o
P9C4h9OR63YqqHDDNdSYeZTEmDCdZPZ6ZSwyiFGjg04iwOtg07ZMvOE674NMSo66rMhBTgf0ZFDk
d4d2ILxRYDdrYmPbbzd2pPF5Hil2++Yu76JH8YSjtd4VGlYCQxPGxyaLM7HHNDC4ze8KKULR2TqW
dFBUjKlvTHMZbcxVg5D01PvTcewd/Cd0/b2l+RRgPftM6vEJfA8VJ4TvPXcDD91P5mIuIDJsc/qN
+dnwagqUcaSk7H9p6Sepo6BZIIpeGPwZv5IZXawSx1M3sjVpBmX+HT7rb3hjVQa1UHCjHvkdPAev
OcchHyI5FJEXmKBHWObdwb88Q1yB8UpFnovdMvXrESTnSUUyJMv1GlqY0W96i+YHrZo/BLQPBnfT
Fg1WTe/h2yW/ospzorumJjU7vUX3bg5KwlrEir8Q3gq9bg2KJkIXz3DX9ksYM2B94ppZYsDScLgF
RDsDgWfNhYA4DQ6NMsgY7GCHiEFAqLZ+CCslwXcGKPmJvCg/0mzqSjsbaALBG3jmRRdrfAlaVMAb
mt6KtN0gUIEop/pQlXjYLnC1y3Kjb6JbZc0A8FTc31vSDeaCq8SN4CAQkghW8pAyWvIpOloNfDg7
wI6NNWljKXMd/GPGJ4CMb0Db8rWVKqMbJjecomOrhRNnyM+1b0oQnIcysVeO1Ih1CX30EBvlO5sY
8ng0YkKHR09uPQ8oJJZWq6YXgXKT4CMMt0ZjZCZ5EuoT2ZJVkVK2z4hvrUnCwrIMf1ezAun9rpNv
AVYZvKLymPzcQ5BQvygYgcx56XhMSmN5oEW2wkEXe+TpGZqdwJJjcUH+tpAoAWAwDiV9y6ZqI+SJ
Ac1Qt9Nu0Cb0G9ZbOjqw7PlUEmYsUhAhrriJlxakC+RQH2MWL88S1OV3hGUY5SUqR7FTZzCy+YOC
AHyMWFcd937xEUVPSoWs10fkuuMXq/eaZkBD4K6ArUse6Zh6rngErI3H0Nwbs24mDtBNdKzubLjv
QDTjMESx7hBwd53tf+DEuA1S2BKGe6p7lH3ox+Em2V8CYo9V+t7Haqzz+s29Ql2X7qnkhB7EpRGi
2RRgrcvBVIFUhMMczGwS/PILhRqedmRO+WO1qf7qfXZK9WdxQK5Qbz88X7a9jjV4wq67PHSzrtRB
jkaUoqCFLweoTsLIXB1H6okDeOIbA7ZGWByX6P9T4jMeRBSulQFi/36yL2e8RTs7nJnAW78tocoK
GpOhkS95T04ST49hpjS7r5CuKnx747MiOoD2GFuXLIvr5r6CnWqm+yFxJCLBdZSxDtXzbvxYwoCU
GKP9spa33rnRftcC66DFzuOMlB0nrGqz/pWLWZlkIyv2OsshnIgBXRDATXQY9G+fi11HX9QtF76T
7U9X55CigsUuLP4+DfnI4Ymho23HZo4U8vrbkFyUAdYDX8Er1qfBRJAVcTYNqjLtGb8Y0lZai8e0
P0PPBF5Clvhka+aoWgCN+wohKyXifGzXXWwT+/yKfJQCVydPZxXWIi1eLRVJX9fVqa9mzHg/vpD2
QkVQiJ6yYgA5MZJt/ZxfEF0GBWMFspaKl/PQAhc/tFrlkiU2/s+zQzAa+jX4fKmglyI7m3ipz1N2
mhe4nroU80AbJqwg6woJBnHPjCO4AZ0PAUMeHmmCD0tj7AzJhn+AybQ4VLxuawiOZinq9KE/qgG8
vKu6z+HHU8j0v45JTNS1i/Dil9y0mNMCh0Y1EJTtgaF2hhBGr1uq2zwkpgc2+TLwg4wXOQw+P5IB
7HWGNIV1PBsNsHE74NjUDjKDeyxnokTKBOz4q7l4To+mJmBqzOl4HY87MTJhb+eypvQHjkMt+qoZ
bh4xUQKc8S5OcE2uv2vsCK1xWNerOyEpqvNvYHm244XXe8KjopLCNxAsUAhYzOZJNTeCjSi1aK5J
pJfMGbXY35SunxcxzSKmDPgW2qpZfq031Aa0Mq5MtifLA98ymyZQGeQXCpo4z5NG0vDC+h9K6be/
ZAVnRGisUHn+guAXw0qWjfftFPyChrUOssGMjMhgdxCqOGhcjIbKuVPRCQAzX3qZfB66uYGVX/mo
FuUcK0wWOGxULykNgG3jT/S64Fhz2TqQJ3UEPBmHEgAh1gHSCB7GkoILPq3xK8p4RjkW8LOso34l
hZpvR5EgmRL/IROdYvn+gNZ8OKWi5BuuRhVwPOwBmhrVPNcDZm9yzYhloj3fZKDPY6cuX0V161w3
smFQGlMfqIXxhgCKkG1UafGgABisHumGFawirttVJtnqwZh/6U3Re1Hcujq/DTQrLn/LHe0TwVno
HBAgNt9tR5mU95TmM0Lg+bmZyBAOe3v64SCrgLCy2YYwJt4B+gFFUdYiXCnzLJ8kVyHS0AVSj1h6
icZwTJkxs5f0vYY+gPvPTt3CefsEZb286BbVehnBSS6Vm0rNaroOjVuClGfd6/ueWKNabzsLgzvT
dNk6vpoAUiK64VJZnxEu87scf3/MSZtc8zXJJ+dn8bfWIwhavcRP65i6dHmlkLzLzre7XDS1glmJ
4BdRwdPWgQTuVlQvfRqqri3mfuAX0D/CpH9YZJ8GSN7w0p7ezxdgoeD+zFAtEA7qV5Vxz96wVtnW
DTxirimcWtuVo911v56USyBE5hFIY2fIemCFttAfFB2d0WQuyqgI0Od7X3ysYzGML+uYtByagWIX
0ZxFynFwCy6a3dqsJYNiAYPdiDrqR3hNA5t4lDnYlAOPB4RqdeUjUp0OgTwgmb9/bjlfk5mAclsH
napOwb5sEh8iwKDOqW7TfE2hhmol14D0bJCh4DEqWfFCtFSe+R4W/oeFHgstayadWSTmbqjXVwb2
gYW+dP5V8fYnQCPKq6ESMyuPPdKOLaJcQ8N/JG5ENLJN/IUU0AfqRFd33M564G7jVPvkE/VyLLMl
h2mtKTikScIagBnQgu22YIsTPrGFgTV+8i+qn9A0YQlVSLRHza3bspa8zsWHULYv2S23B/qLzFoU
Xgu2rJ5jlKoP+P4Ak/8HZTPu0Ur38pMYKZe7oF0fixhJ6nDhSNGO8a6APLGHoiWoJs2kqQoXMbVy
bxrRiWQxIsiJi0IDzSy4KPn1/72o2j7ZJnMnxPdQN9f9Th3cOZVbr9Cw/lzSk3mLDzKBMwWGy178
g7nM9PS0E66yKsfwB7qs52InK/kh5eZ9H8rzQZqW/DzemMoPR3VQVX4BzkSZpAQXdmU9nkOFjbeo
4GVkBp+6ETTafXObPSNpQU73h71OrUZ9NXigyA5Bsrwl2L91r0f4+F6I0ZHuZpIGBJ5H47mS0hU/
UFCFlgSjC3BK1PTwWzCZagnCK2x4wNGCCV0f5d1swEOJ0FF8DhrNKtlTaVu4klTh+5Grs4gj0VGv
7b8rfMJAlJTZ3Omdlf0z9GvowrJcK/idVbUrSKxUeyylFMPFOQjbp8IPNX/EQIuED+E5BUeZEChS
tSyZImciuLQ7+JTZu5GteNxN/XQcTF3P8cl47sJ3EKzfFIjGYvKwvwZMZy6jNsUv1Y4PyImCE/Oy
6eEVdxMhd6PVUlZb7qhg9XG5Z7hSXWY8E56962sl26UV3D5Q8qeOxvcSE1auhoT1s9N2AQId3PVG
t1c6WloBgp1//uJ7bUVC0866CxtDCS9GSzCoVwrbi0qCldsAR9OtnvFqx/zUYnnHiIgHObLL54Nr
vHbIDyPlRWDhC3D7jkzSnXgRI5zGIJd4pV1Hc6Q1BaPO0LKIEnS0F6I5NwT+QDDXx5fRq0HN3wiE
f5DL44LuzpFjGTakYw6UBaqA9HObxYs1376pjFmAQE+ui6ENOxPodqEWRbgwcIAhblfyhERhtYtr
iR/pXoeLTJwhiWqAROIKjEbtG4pXRzBNs6oDvkeomojxQsfPh5cTiAbYsutryVLKFsnxpengJYNg
KkhPWohTv3oG8atgY8NNEPTyyT2G+uagDClr2DwDFL8nd7xleUuA+hsqVgmJmTbZUb7SO5hwleRO
hFFQD882S8phIw7tCe0B4eP3rH6ysAOgI+yFZoH4csLqVRUBDZFIOtLcBHQsu6T+y3Bj22kii7Dq
Ydhwo2vmJSTbQElnm3CkbduFkv+i0YxXgSouxjHbPZKZPzvUvtWPDAmF5BhQhJegFHdqVMFeK078
pXRCG0FJRCgH8qU5hfNbpuMoTYW8/1OQC7s5qMgElqmN+jLDnYH5RNPQw/aJKhmKj2IzEAwQmqrz
wXm82D5j1ev7+sAIekf1oBG6EhqGZseTbRjUP9iaIkOMuFbRPIVVLL1xVZb5R5GHQK1tXFdAb6Tr
MvHhOHT4kquaADpWrf/TVVoppkrXQ0Gm+jfCWI2VZshzrHN58WfW4hSkjy7P/SzpAe5LUy8fqe9R
t7r0dem+5jdQW0XtPCL1IMS2FmckA/blT3qa1DhYMZR3aLxEROnYLeacQbmENXtN7ntHJ/uU6s/c
gavEdXSbVK/0Y5knglStyUx9gnc3OaFG2g3GKp15kvHddoNWBGTLZDKh/V1rc09DhMnA55rH/RhJ
KETRu655M08DIl4FErJxDHLyJ7y2UGilcdC6YKhCsdy/PzYOfBaesTpFCFbpzcpRPFmcqm40ns4z
LEFMAhDMlNvus1Udg6J4tCb6aee+64sfMKaIyabimSPJljcQw55T8+fLQioCWcVOYhQCYZ2T2Q3h
tugo10d2/ArBcg1HOatj2JMHPHNnV64w6+3SfIaKRqRVtilAXYWtMlIhN578VvdwPZr9hiVpiWUI
3b3CixFUQa0v5QtS+TLESzl2uVK95kyyqRyNZZjRp5MhayLUp2SzawceuJHu2exKEira1EIqwHqg
jFwHY59PUqjKNhYQsWfiCQnaXRSI+mSY0YUVfzzqM/4stu9s1xOe6SK11lLGcZxfPRmbT0KnyZ/E
DESW/WUMw+nw8B1cPKheYhMp+y1MNSD8NufFp3zQlFE5BI7ItLF1r3mUVPgL4+5+mWdnb/UZXgdF
yrjXFBJ2JhGDzepnjGBX9D5NvIoNvaXtnYR3/XQ7RpsZq9tYQsJJpIgDPfkYm0mfn4rgGrzCzhCg
Dwsitvu10F/ogbC6CCGnZr9vjrLEIdCfAJ7iLGxDRrsNeqz9VNO1ZtJ6jlip6iuL1YBkUUT7dRJ7
EL/yX1risHOdEr94ErEJV8BUiUdTTlI0gvOk6fEPgXDSuZCTC+GliIaEKBhCNrgRXrGobxmcU7CF
VsUzopiq1MLvV2L9/J4NwOZcbtyx9WHAiPlqzjU4XJhV9/f457wtX3l/KJEk/YPnQpg6H7QKPOOi
hR2YHqyM2q2W48vWvVSsWrq87NC3d1PvzN8qHMebupEyfm3ErdctKKNghs4ZsWqBELr29Bh0NlnK
nOMM6YvCPPIXa7/uGl1dTSVUjMcz34wmECwHh66vxAxZoUg4XL1f+TCDVp0u4Kjpv3ZDREaSELTG
O+AdS3/U+0OTWk6OhF2yCMzEffgCYAWBhmasY2EBeeVYH4AoGW1y3gLsk+nCFmO5fojLHvdcxa9G
OuVfll8GhiiiczynmNUHOk/NBK4UaISt+IMH6HkArnvOtjbRWtOhAO/77NXSLuy64dDQ6LQ+bQIO
KPCnZo7yeJRQoHwsmZW8bW0wh5RqBVtxVXBS9/bkoohXKOhUNamnVV84F5PeSjr7LcR3ifIeA2TB
FkABVtG07ax7VmJfr30SFnssckbmLuf/RuilIA4UhLoq/6BkNoBh4VoLsm3pGq0+21XIoH5bOj8s
nADX1F5XZpKliU8ZLv0gtqS7tT479hXfSmsjmNkRU3bTFBhz8MHSfPGzNWCWh6r0FfkgabgoQpkt
1fYtGZMFfA7ogIx105ZBRgb5CJ+qn3HxHBXNfiJ8E2judRMsRpXnzeNIRWM9gJp7WHPV9gguuepg
+NBbiSypK1UXtBOElCM2fB4X6ZW5yOyhh8TR71XHYupcbiCmqT7Ic7BmrMDjDOJddKcE/e7d/68W
E+knQrYZxEDZu2uV7JGwJasQmFV7ZIB8F8zPQUK5O7fgmPQaBn3nkwCJ2XLS5jJFhWcwIZ4p0hqX
Qr20wbhVHEUtkXE10H3NHoWpZ9UetO/dhhffy3BSXiDrqnxabmcbL17AfKHuCEhCqErmfn7crIAx
P/cvZhyZE+NTtUOmY3wMJwWCK9acyXVpeVQ7wVGP/mOYWbqsT52JlYTFpa31aXUPWfqFgtCWdE7b
aiVnw7ZRj/mIOczS0Dz8ZfWwXNQiUhG+TcC6iMISQjjxjnL9aXtfy4nxe677mkRVB2bZHYmkI79F
k/O3rW9LskEBxSNKsJomJDhNbBl8bNmZZdqd1UTl8dzTd1THfUzTupqgOJOWuBwPfHtr6hJX0T3g
K8oN9zwmFdXCJ/4nZSoTmCFNDNkfXaNwDiV98ix17Ha+c/ZQU0ZOjXX7ZkLROEMegwSyaGAABe+t
CVQMGnsFO1zKBuXUfPlYT5cJGmbFcUSWDkTFMYVKimAzQqc8RvoF8FG75CPmlKrNC5nU92tX+aP8
YWcS09QKO6+fZ+IhsTzh8ZTDAX1KcNYPZRvmKnJ8IDYCFuXTSMTVQ0NgB3BzV2ggEzKhq34DmaNu
jQXPQJXNSEOWFt3l9c6KpsquLfFVDNYVc45sj8ndIkw1DzZY9kX8+M+MEJmRIOGRF/CIOqrj68+/
MAhw+eLKRP1zS7iqPvIoFIj4YtxdH0+8rAVOEW3lxpsc/Wa2rrkJIdcu5p/1vZ12rGXA35I8Az9B
6UqfQ9DQ8xWWDFjIQ9iUxSnum0Vp9SLhB40NRmpjlcefqu0L3JuVX+pEZ1bWt/pBUH4eBkgeCIE9
tN4Xaxnrj0QTt4d9Fpt91cNrP2Mc5RV2UN2+p9K9pKhspNwvj1HyG4emIPJzv1v5IlU/knJX0HRO
KW6F7GH14u0cLm0BtqtHei8nEAy6B6jtS91ahM9C/+wMjTr8+JJz3EFxa28MhbNuIZ/pi9gQ+nPB
42cy5m2PTcQvniP/G3t0xC+u7beEk8b+mXNtwkWy7sYBJf+CcfApWdwM86vrNCx7jCwDEXXgRWo0
sybE6Sd/Pu6OiXM2qa4QZKdLnLET1zSjgfh6ggMDU6TFu1LX5h0JEnwehbfV4HC/z5X/Amp295Ss
BUK6kk5oAb1iSVT4ZmHb9djNkv9FAhEinl1UGsEg7xXo09HtE6Uwn5MLrbkNohFnDeiI3zNNff/3
vdZUfVPRWgn7Ov9iOEVQAyPvnAPnfUBU1fU31nf6regEEbAmXfoJ/1I1WcRl2lqoSF6xWRZS5k4D
ehCgTB5oyujzfEv0dp44uKm+cr3QOZgoXU9PJUEnoalENvW2hQhQbAb5Ax/ZCRJJR0s7hosSm79t
HcRPSvf5MCy/PJXo87r45UlHgdnK20w1xbBPXQYuY8ixtv10INi2AGuhq4EVUhGbsBpfedAkIt30
AdCeuNzMweA/V58sH0LL7YRqJS0GjdV99WRNOyNSsVwkMzsfgXemFs8L3THnIl5aYd3lQqt8vDFJ
GF3WPZmqDZUgagZllqJvlZx76iGGZfUdiImlIeMKKSLwuMFFUlcQeIbapmefxn5AXinq/ocgov4d
V+IKiyW/Nl/OTeFogKlHY6dr+IbzN4mODg9mz2Qp4pLIUOA19ni5CYIlSUlVkH1jOONwgYzMPGRT
WGN5+Gn7Z3djJCYTu/kIZ4jTQmY7n8xEIQkxiIxgQSyyeHeFiQbZwXP6EBaQc3DlV07Rd4PQmJ9i
XPtpD5oUWj6Qjb9bTvjVCTRWFVfd+gPNaE+w0EqO7aCbOWyULPfrZ2u/SK2wlneCxBX1Due34rl2
9wq94AY2mYi+hNPJoe6Z9W0fJ0wXC5w7VQBM7PaldXE6yh4B4fUVcr5KI41ICzEbQa9i7sYYHRNk
x7fm9M4pmAzu3I80t/0BeVHN6zeh7cmMYR+dEGZKAOhpxDgr+Ymy7RvsUedXoRHttMcyDIbTuSwP
QKxXv0qFVGI2Raf5y/6jHvLR2eVk5bxT706HvbFNeo4TIlo2sIcIhobHVEHK4yXn4d2kOU4KbED0
BIDJdhGCtKEAWNm/mo9NzRHvlHvOMcMejASOX2WJkgLHVsgjoMl9SflijOQsmP6NKW/KdE1UQQJ/
jq42idVgXAhYIgCA6rksTCGGYVnVIgeiMV/CFlOsQRtHuS14GJfo0A66QFQ3gKARKlMgtxHEoqdB
JE1KKCmCCRHQ9lCl9eSIed8b9iLJtIbgJVp9VfyWMohVO90nD/h2e1gH3b72+y3PSXzCvGncq04T
tMmBlAj80mioAbUFHgKP5oJHH5Bs9eKDm2ZHSY0QJCQ7LIqcoNm/29tzMnchk0fE2MVjTmYpXIBj
ByMgpONPGF3q74mnw1iQrqzDK1KUQeAwhOlBJeW+Y76mfiBtHU/HBm2riuVRyMfo2U5LQjvjv/RQ
BIjd4IXtyXRKdwaPTIBMm3WSPbP+wn11mWNWcj8LAkXVJ1mQ4OwN/IWae9/ByVNPynLwtVx+kQMv
DxPmtSnpz8NWyOU51LvRB5Fa5UOwQ3NZQFc1ic/jJYnd7g0dBq5AztdsO84znyc3qH3tkPnDR52+
SnsjbeVOW4NyITpA7nSB6xskWS4P+ZbHpPAnXZWqEkiV7fRPe5XktrW6khgpQXK6nnFdh1Khit2F
kyGVS8PdFu5c1AL0I5JaIf7joiVQARPIqkBsklkGeo6obx+ZoLoYJWVaffoeLEYxuAFaBvc4+3xm
Q5FgJCIgBdb3nTNmPA6+a0r5tfIgUi7tD4lJnEp2BI2rfut4pBX3BOqCaqzvZdUHNUdoX5P7C6NN
7FRQNQe/vM1h8pbtbZokztgV99rccUARl1+qxQzhrVE8S2AfQ6yRMxxcxUPeLEf/P1i8wsARd0eC
qH3ktMEDVuxKr0YElSL25LJ1IVQuvFx+Ki6oedQh4R2jF+7T82KjBhrlO8j2p+13rVuCnxMeDeWy
Xixz27I3i1xfQum0xugMBIHE6c3XU0gjMUnj7JKyJyLg+mO4WxFqphGspriNJzL8wp33wQeqh/dB
MdO8wO5LdShb0u/Y5l1RdegIoCOq7J5tpF6KdI/0LZcdWdIfWuy5o5KDIq6EuGjgMML7v3dQ8tlG
mvDpPTJa7gRQv61gePJsH9R3ACC/jJp+cIAL2UryjKzNVwpbFkxQEwoJJvGUy/dJtitptxlaf8z7
15FU62uYiVVYA9YG7qvXSt9omUQlAXXP3P1QIJIUKTcrwUm63Ihf1rP9sPDTmkbJlXx6NNSm+ZTr
DF0Vh4fy6h07DteTfgeppReNx4H2GCmubg2DJowHJdkAP6HXxBLjkP7ttLcRtujqLEaff48XxAup
R5H6TSEr+k+lT2foM+Htn64bP5X7qS9xjl2bl6FjsnbI/wB8/gKxe11oylJDGv+wiPZNXEmHbOAy
qZt2Z2B0kFCf8paFSjGFx/osgeJ6wc3GViTBNHgCPCddHRFHkKm5m8wyT5xk87ADaHHrbgxCpn/d
IM4k9yVJTsCKhsxYouveDcgKVWvds4zwuKuo1ck4aTKXQTdFNKPLEbHkiABrh8Olvn9t4IX9+s7c
ZnbHI/XVVW3HZ2fYxDhiyGX9G32zY2UBW2bw/0q22Ek4ewfH81mS0SEJakuiJwKX1L/TiVSGrWUo
QM8Woh7u/limAc2PJbaSYXzH+sDJ0UMo586baIC//3q7Dmi10o9yE1aTyQtb0o/AvDHUkMEfmh2V
D9s5EvAQhN0pLFQWshfCOrcMF4b2mtw9Yw0Mqk/1xKjeyR1C8f2uuShbgeLgcXMKGYxkm8ipahav
5PPOqEc8bRbY6E8CwOcoW8jjyEDBHo/C4as1nnOzyAgVvM6aq0LdOZbHSyhnVryfBXCGtF+C1VhM
XnlXT1GT2URp1Egwzuw8ZRbsgf/Ud5Fsy/5a7vEVGwHPjRDShEbLf5VD2oPgyUEhTAPUBCPGwVGU
Z6Ph9azGC428jqhpvHHgtcr1aACi2PktsOQpY2PcDeXC1NhnYOOgVIjKVaupYuo+XWuVZp9uSPEk
bN8zm3/+AyJq4m60rxlzMwYMCcjqzttJ7/j9KlNv/jxfrUzWUmiB8phfzcTfAl2Rq9+OeFNKXRg5
wFN6n1NisxJEw7hy6gIP5sTVVISncTHy2e771CaZBC28LEmYQOVzXyDoelMJ85pH+zI5fFiQ3/ur
11dCSK5GYMp159LBB3p95ihpDeqmvuH3bMxlWi5O9InxBfdwcWq8qwByeU3O36+i4pacN5Ir/WO+
XL8ajGRjNbBJUT96UUvUVZIcH5nfm5gBpMe7rSH/s3ihKF0m2wtA5qJjsqHoPK93FHeTQRJGpgGx
9hioHl4goptgGm3yaCtieLLgBS/CN3dFrTqH3TrzftbaZNuC2sD+56Qs96vhEiwTpoXeJZTjIwrJ
yd/l7/VHVRgETyuB5s79+Pg03AUu0pEzR4efJmafB5YOKeAbg9ONHRzCYoT5ORv6iKD3DKc7ZZjF
tnIxXthLF3Fl3/Ue7Sl0PNONe2XHQP5HW0KHa8LnaaqFv9cJYdHToytwn8tBqJqEbrDQniu4AcAz
ay6wTKvteikM+l2m575uM2kWVxFwZki/VIXPGp1AbP5jsF/o93OfFZGxvhXipdbce3bUh4vfnEQS
QVyZH9+dtIyBivqXreWHh6rlc/Y0ntxi3R3b0gE9N99YT0qCr+WtOXM6sEMbDZD022kCk5GM41Hn
S1qnEAyQcG2ZUwIKTXO+R7eyuquUSlxfDuscL4ikXerUg3GZsvWVROXzfTnGaJ0GjilEBGsdBSqL
mpzyJaZu2Eq7cm6HkAk4tncaoQ6gop/PBiOBbqCP+zhOy6VFG7VY1jRvmyOP5NII9nS5MtTuGocR
CaEaOLx/qL+vRpkUQT8iz0fYjg138dkfodCUe8nWlhGHfhnsW/ZLGysD4OytGY5ckplxtK+HvEb1
xJ3GWF9/yfHUCzDAhlbMO+/McUAet3ko+/FbvUd01LBfCebUyBlA8yoRML9KTLl+2WVamPCOH5T1
irVwPyIbVoWxj4tOu/hziVdG2r4hnVxey/oaZZPC7piYtw1fsgzxMBvlrmW7UATrFYEyIBAPwYQP
/gf9I5nEZKJGhoYqJZHV7YoaZuzySjWHeFwra9ij0d15Lhqm5Zt+jreRjYMND3CB59sMq3DLyO9Q
wLi6fX+vaIQN/rQmxjFOxfkZJKf2Q967pAw+j66WDIsPIrVeOovxUDFQ0UPJ4V+ApvaBgl46RiPS
ocZ972pjWhv2vCLlwDFj06NHdpGtHeJCme3SCuBP28zsdlFBFCQynLVfnYLW53XjdrfrHeGP3OPn
X0WVkMAqdKG+WbQ0OKy6eoRdKA9DITu0Bq/xKv2u81QfsLgF1Md+s9iMGlG1z/NOVQTcVa7PEviA
i/af3J+uJRF4kyA+CWh2y8ia7HBZcD7rdvu0BR5xRBv1z96/Ujl2A275TJEG/mF+iozg3lZv4Fs1
Ep/IHKAZGCiBHSzEWnXC6KWHJRSE6zEoTxntEOD5Dr4cvcbF0lCi8QKXu+Ndcw6icj+fooSB6stY
x3E1tW7yoNzXFiDCTB5Nh6/CJIxzOaNUCqH9F5bpc6IWeWa272pQEbWVcpkrRBt+xVv2xKhUrk1o
E9bPPeKdc4lTlTfbPA2U1kt0n3EhJOsn9BNh8d4wjX3NI3glSOWxUraJbJA25r/6knJ1Z3+6Whn3
bdZOgzalKJwQrhTrn/IBn1ri5L2OPRdJczACntywgdYKkuAe6o9/QyFI8hGrOnRPeyb6G0NhZ0wu
QjJh/6DHcwqanP9sEPBU3hbAakoUsIowVDHNxICnYL1PgcXoTF5wRlt3CTMelHNzP/CHpyDbE1sS
Zbj5Ku+i5bCSUAmpTZURT4BancY/MRptGT5oHzlLjHHKbFjedoLVmWwcpwIQjUZYv/yiMup4lfk6
96gQgNPWvA9Xw4z6ZS1LfiPipaSrBqR/QSTz6/VsCuueT7HrYGrejbwhz/dYUwCHwCV3unAK6T/r
K7f8r600hC/6teNIVfjcXdEguBS9OD4cpfcQyL0mKQ903z+r6QMqlO18uPXXwQOMe1zuMDJkgqmN
8QjNQs5cFWpTvKEgbgQsObYj0wlSpZcbVqHmSvbKWlf/OrdLc/ni4K5jsld342lhovRyvwDj5vio
lRI9RdNMaeQWy6LYXTx2Gq49iKkpl+JChg+msO1YdZ6rgarZInEeh29ITAUsk8dLl40ypYvim/HQ
tOsa4nms5bZUYCprCRtZaJatFkVMfA/7niasFQGKRXwVB1m/XiD4s+GBu1eDiqiqc3S3D+KqekrI
dbO9/oboENPmeDdaD4wTH9LZqKug0/Lhk4tVVMfMQwm41pQugsTQO/5OPATRU5OLNIJwhDMbkIx8
El4w4Fw46FNDXrX7lLCluK9djELeJJ6Ox9ACiL86gXR2io9kowx18ON4LVKxTBq/iWNAUKa0RDYA
+qJt6hdRRrjPNSwP5HycWBTptYWpNjKjrjjmTrxJoH3dbIgkNycDkhaXa5NHrpw7oaZh6SmRhYcW
YmanaGc61gDqfn1Z5SXTcxswHgb2KxfsemmX6c26bfwSj4B2ni7Mv2/i2/R/fMT6QFmWORdcxdtj
QIkId4ZLlS9IlqbEW55bsJpW2edY7kvvvrGqRZcVXdS8I43+sGcKKhDgbIYyURyFuWY6F4kaTHvm
L8F+Zw+akMpH6iCFx8OxEuwZgeYqDSZtkKSJpnyw6CclLvJJC97oNAo5UQCMm46aH3sRGmwiKEAo
B1mckxni72P+Eq2s1zqVHG+2MvTqvYlFii0ctsRF6iNriVUvzFKtrrqALSrlFz7F7Y5dFcskajvv
9I1m70L7dMb8UV9dWGQLjjJx9qX+lR55cLXhN1ciMQQhGrm/gjJtxerJCBvZ3/rQTKe48CrjdJFK
3kOFPTalzIBSvokQug0yOKpAcaHaw5x8pWErfj5LRwZCP+8zLmsIj6SwWGgCobVrh0fJAhFLmg/n
lczfopH0BgR3jo3FsxBhsnb7sHLmr192zmooKiQfsNH64XGKbxHDKKaAh5Gz6HiCOU/4Ko6LSSS+
WtAL6PJgHUSVEAQlbrVQXTvwYnY4Voc/m5RHtOV2LgSc+MygXvXMUTletXn/xP20eHv4miSPh4GH
TD1VvALDKcpx8V3MDMnjq1xScZkGWmjAsU5gu8aLYuwovFRlMc/cCguLtjTe5wycq+FgHot/p41E
14ZOFzov3KBCV+BFqC/YlWVX+LLZrpsgOPXJtgZI+liBUOYi3IFho3H8WBGv9D8S0sFizA5OO/Jk
b1bsKsyAcputwUeqAl6/d5jZPHBbwZUrgPnNfpkZsta7NAkX1WVbNkftTYOF/DZ5EYzFrt4GZBD3
MTwoLz2f9sIiOLqrsrtwasuN7gGnZ1/eMVYQCRMT4zuILjRUlqlgtMhPtuQ6AwIT7a/enOBsbCeV
FcieJTOplAGv24WLpPfNaDxD4eg83PeqxE28/gS7mSWzcx2N0N4dO5jd1juq3ptLPdr34FYYCR+W
cGgqOEwcO4aypvqPPGYfgYJ+lL4oM+uIrmocQYTMc0lfkwkV/Wn6RMVwBoJpF60TBSoPHs1Cn2S+
euGRUMR30dLgJjHs8UyQ99qf5i8kPFK0BBglHkff115dGnS3CpLvuukZxUdspiLZcsr9l9xm9iCH
Loab/XC978D8RgnmCvXK4twOduSKwuuZoF1J52+CaBzAxKE6dgIqD9nmzPzWZ4Gg2dXMIOsY2fzQ
I1XQE/j2vq5d1TSpap71uSGsDOQCUzg6EoOE9JtJulSgRViyIQqEVVAZIa2+7IRvFB30VewiQnH/
hXRIYynsAsV8iqopDsk2yQE+wf7sGqBLFwcEFINS1n1SVlnwHL0EDMFKCli6wAly5G7T4rfrvOi7
W3FAX7yZQmPZkCh/421a1aG9Amb1PN7vlS8pE2sFNp8LqUD0o9gdW0sEWAv+0M5cE60ldemEJIeX
D3tYeOfD6A4ImFxSrSTmdEfHjeYQfaB2nMEfIO/jwVEDpRvB+i8htinjS4zCt7ZvaErLvMsEWC9f
5S1cxj+npkzr6b7ma474kZEULH/NXGA0U8uMJboho6EYvxh7ffVZ/NQZvfnh9aR5B9kEWrdPW+G5
v5eusN4FlNfWU9TCCgvd34oT0Jv0V3TbGUcnU/4MJAi+L+5l/kknvjcS023Y43UwVc63hUrz1/Zd
jxP8rS4sEJ3e7VQYM5fKe1fD01j+IMKgM1wNGhZr0XDDgCXtRhbKkDQIgSjmhUf/1YbGRCYNUiUO
vtb7mlgNzbpljnH9EH3h5K6sMRTVClz3CR2zoHyUpLZlbL5b3iJaQserfBNCARz0DGKbGIqKyXYV
qSZQiG1D5GqZ5cHBStwe4/VvJJjohlfC20eLk2uz9LQQN0MKUJ5hBWyE06csxuecYQZh4cbxHob/
n0UauXXiSlbxhiRf1Jw91SVg1vhyvmO26kwDuCXvYWGdP0Q2+rPPY5cExsQLoeXK6JU9Ri+xKcsp
cXLCszjiLzVshtYBS3CTJpmn1KksJvQ+PA2ZPWAznZFsb1jYkSakOFiIFiAIESu3e1VX0jcie+0x
hEkXBHdFAR6/+zalPm6h8UBeTBN0PjH9W9/wAggsGEp9Lv7Oy0jll4bkOiXU5feVtNZGjZkGT1I8
vptNbc+UWdtBI4u6poWhE5gs6wUwnQDrgxQrm15wfdt5k7WbOW1yuim29JFlaAFEeeoawBuv6WkC
bv+EnSGm5YycUOMntp4CZ3sW0DRHAmvwFhJaaaHQv5uHnslJbcmu766Jzhv13hQkq6Ut0EwQzRKL
7TA46lkCWZ2VvzZgkXRXPpH1rgSM73EqholPqQ2bAUniAoRothDDSV4zf0eTiK+lyaPfC2coR2WW
oLH8q5B3KJDtXd3GSOhYuVxeA2QvNlUxEhGm0kKuFfTI4g7D7qrWOQFK8PgX4ggnxbUQn8JF/uy/
ZQpuUYGspQsrDvFNFgfmYrRgrfxwJJffn69sqbItSRGx7AEqc9/NgL1Tp+eW8TTZm1vksx6AWiKr
Vn3V5S+o5au+lSKN84k7QeBsg32RPbi8PPR7oPGCZFz+iV2dYovx1Q2GDBNihrRBxIQ3ojWzN8wx
oZLUAEoIV4GS7wNt1YLfRXQrSHcUzyH8POSWmmvumtXrwLVy9tNNM3LGmfPb5drDjFl9bXN7vKP5
ejZOBzSX8u7iWC6AeMx3aM/tdco3wJDY9VpcutZSn15WRcuu2igOWlCjLOpOeGBgxnGmYoDl5bsL
sVeaMNK42WHDyn9SVoFa78HttoqpT54OWeqbMgiG2Wr6JJwYDL1FuDasR20IASEGbUiTdNureGbL
5Wv7OxUu16DWevqUldvhrVtwYDJynSpWc8RNSApFlVLfqfCaJ3rtkc3XQ9PC6e0ywyNGCHa6natD
pJvMctEzRAFutdPXQ5TRpJ+A69QF4ZC6Vc/Fca7IwM0Um8qQ6MLxitV0oRVkgPlOoi844W+9sWaf
a1ffPpHYxbCjh+XoMCo8pxRBlCpSL3qjkGiuu70Sc2XZPZv4nbJa0cWBHM11kKOL9fk+CCG3jfxI
k6G5q0KJZ0yHBUWYBk+06gjJkstb0QluTw/IBxmle0RRE2USi0uweVUHY8C8V3PFf5CLJ+k1PYaR
Mz8tbUjTayG3o+LAe5Y2XlEP3IL/WABudungRHCFQhFjWoMfGOu2GqRqp7QPijNyFsJsGSAeD9Or
HWmhQbFfyBXBaNgWIsrh323u8E58fdpHPjAPE+NBpp+BLcIXNVRY0DUfkrkfQx5VDqrf75MD1/Cu
V2NeS0ODWYJ2lTDP/16KM+Ysn1GWof93/a9iM5AqLXtCSnbCbswnLuQ3YuKoMbyZRIBne5JIqLOm
T5mJzp9Sjrtab5aX7+BiYdOjBjlmIU6W69iixNmAmNpJExMNYbphBF/42121WTLazeuxT2k4rTgj
K8Adqu/YvtDvbXmW6jftqb1SFPTgP5H/W3K/pYgxsUNirLWRLs8xWUbRi5P5fsdgVhgriD9qwQrB
F+TQRwWloCmAbtW8wvTyzA8tsbwwmcJuhlK1FqxyWr86WnaeDDSX7xWv/sfduKS5HTe5xC6j+RwO
UjQKQJpnLNdjsvr3TtU85D1hhTYWnas9gUX0FBEXTc3xIHB4Vhe/YBUjR0w5U3makGNZTHQ17FIw
ZwU51m4zLYdtPIdK3MWpbzs1qPPEd3cBRdQsz1W+9Hg43uLtZv9EEEaUhE7Y/sbhBKpmvzcAsH2V
Iey6FuyjBbDFrozBNmGypPB9FnbdDEtJCzQ+YxUb6AeaOW0hk2u9KQpdaSUtPvquBTrPR5A+xwBx
MOsBs4aKku9pZz10v1LM/n+Miz1hMwSX/oG+HCZRs1IRrTBeYVfp3NpOnJJ3T8lv0fTfbjfY6EtG
0CmG2O4l5DG8liTl8mkWz6JjDTyr+rfS4xeNK7Aidpens71/pv2tLVScd1qWWnS75tpz6aCl4Wx8
U4czUH702Vh9Zjl3PPMrdStYd6RdFjf9vTnlnqSoBq3sfGHEXHQhcVO8/B5bZz7mhAUs7jlD3eIE
15fS+UV1QVgya9fTYWRlkfZU+Br3NxTw68thJKEb1oKYTq5PMd7yewY9CIwqwL8xu7RGsMfd1aA6
tGBubUSkB41rD3cOT3tb65cLR3JRbKcOKJgJceBq4rU18bUNdYhC+q3x/iVtX1UBCo3e0nMKvjKa
kB6tVl/c5Ksq//0HB7SKLOrek20KxOgoEpLlukn9OVRH1l+FhKd1FzO1tGxxyyrz6bbHwqmvhO0b
fjEiZPqx7cau5Ck9jO94/BdXH3ITQqmEOKsuiCiIhWJqOKC8c1S2SyQ8cnZd3AjifWxHGJnvqb0o
sNpbqQmsldaGGNBhdXilvq4gIFrQQ9Gu2nkcFlAeB2r0BrU30/Z7JuHdJIKccINHD1d6+vaakLVr
9S5qkANUFyyNAQZCF416wzfSkqusbIoYFBDwFYQ5jboLYOt2kJCDcT4fJnGitzSqGM/X8pARpjIL
kIZTcpTTR7m1Zdlo4isGeMJYDvwpkVSbfxIhBWddgwaKcUXaNZgKfrcFAJeHx0joLURUV24NaNAS
pJbBGsZNwoLYivRxA2Er8BCUpXDADvsH7y3xQVdAwV9AO4lXETyNkvaAMn2P0esJAHUfT2leCU+e
oK6J55aS35Z3kW94RZAXGIQwbFRoBm/02937ug16lKOA5D5IADda6q64/2Iowxqi4sPr4nALEJqg
wd8rv1MMe4IDHmfELXq/EoH/CRHVAlCLvNT7/FmEgzSA7CqVVFvyLQtuPwTCC4h/86EN0ps8WPS0
0Qqt3OE26GUeGKVXXm3oIQqDw5otqPk6hGqv5nGIMZVCVg4oEegEYj7NEUNSZmWPIA6z089nvwGE
GdGE2PC8TA+KCC+iEtx0UtjlGwJAT+3gglsSvYf+bWHDhm9wM3L4hcuoe3eVz07ugi/H+YExffSo
lbgCikpKphHm7VxjxekZjbId5BewxTZKDzp8nwu0HfQb8mbBnzpz8Qcp4X1eRzaWsc7+ftQnB5Vt
7mGSKmrCuE7RqGsmGxYLHEbOQrfTPIf758TR3GwR5s/uwI4t3XcR4yTocuOa1SpqXEnIHuiBboU3
p3NGCuWX+mK49lM9rqK2BRDJNiQJW4SjY98U+hwMPHVOL80sD+gXUgoYIlj8iHI+nWd0Tdyjgw1R
KOfO51MkCGIf+A9Hral46mPnaiI1YaFMg3JwkjkGzpYQQF/pfnNxGL/UYZmFoVB94RZ+iPLqAOFz
vG0hEmlHFD3l7Y4OrgHWOoxADq+ySpionPzsNNBHyBYoc/il2825WOJz/Hp6tLXoV13yfC7b705F
NdJ8t24XiJS5vY1tQ6MbTZHsMfT8TOZ94JNVPjfIYadHN6AkUjpxu4Fa+saZfvrryFWn409+aI9+
CWR90ZP9EjZhk6EYAJwZZRh1HHuVEeW9dEWpzWvSLV5cuFJHpmAvWTZXwSsEnmhl2sKM63pZphQw
3lbQTdHX9pdC0epa3yxKGz2+XuskFeAm3dmcL0VHGt0DFpMWH32qHC+8LN/NBVCEOLavc7D7+M5g
VzIaGBWqxZXS0VOwG3Vd5KkFRYOo40o70vUoTzE1S+oSu7ndgZyN30CKzqdRKtLZGpFiy4QjiOXh
7mrNUHuDIddz1FbIV4YwDyEVNP+khq84LS/pp2vZD44wtc0ovO7i+z4TX0eh0/f842K9+4mCMrT3
7lCMMUgqz81LsLwiIMxGj0zacBU3RGPq+pDeoEFAag9efXsLZ5wce37Z2n7q4HZLrnx1jksB/4/n
g8Dx5Jp9TDpnAw+bUj2eq6dDGCnZmVx0OvQJIqIafdAAKJ0hacsJZfux/P4shrH+JXmsYfI/nc4c
gOLeEGnnW6RbpEX16OBKBPBLiclYDgI5GaS7ERHMSXmTpPo8hEAfohhPiMaSuzkIRbKuGmbdW38v
NhFyW+2UlNeRz4/AgFQbqjOUBFLDQeWKTcoyZqP9jDQtFj+WwvpHgnHiGn5BzFVC49ZvSAW98poS
dLBT2JTirXbPiiji3zJqLHFPvpReD5oG56/+5h4Ztp24XKIqylLc+eUKwkZ4uwU64GkQ21cXWjwf
hgMoMwZFMDDsrAP6pDq1SdBnQlNL8xGFyFlDLKuIh2bTOibYcHHP4dZsEDNiyE0hRwKtlyI3jkS1
wvdtq1npJ5dyGq5J/SvaV6ujiysHR4yP7/CL4h36nOHfOTUT3WYVYaqBWaCWqPCtemZxw6d8cwvK
4Ka9/VJBMrDp6MdbnDhJQSRNBL+Uvph/OhJwuOgmAT1Sfi1pYk2P7c0ui8qyefkxz5DoabEWub71
Awwxc3mjurdN5Cq59hk7TCCl4u1qJBKH2dn1li6qeTbb91qXHE5RP4YP5yxCVITgDp8ZuDOlynQd
hGD4zqAOJkamHqOG/fFZvHZIGTodVbfIZBINsh2lB7L7rrDrjd56pQb0T3vL/GMnFMaLyU8cDOo5
Mvu41Jr1tp9RbZ1oWpJbU7pHp72q8xeDEEqWTWoepNxxIfu7X8THT4t2Mu1vJ5pwkDJ6VeEgHEJJ
0G0JApccsNTjqPSMPvRzEs0Dl+t7JzfmgrQxlES0iF0ifcVu0Cr5/kTmU99fZz2b7x2pax8Ioegn
nsc8nY/9niaoMDaDf+P1QoQOewOLD8TyBYVSAx+bGZpk2pcpHWxQpXgxqM+x+Ii62VlEsXPMcXCp
YzIC2XpTxzUzcY0v6NcHAhwb8Y+pRLZ3abwvdCzKhWHQ83jVnaI5Jgoj52EQss3KIJoQWghzxW3D
7DUVw0uG40/5Acp0M4SgbJ43M90tbgowjOb7wFsGpqTXc6sImTIJZSui9S05zUiAgLN+K701hKOj
4KalSsfTYn1PU6L1G1Q6hQdDgeiFVWr8mkE5/qjlU1yWW39R4voBEECM2sb0I9ddeGITVXGDLDNo
Wa78y9rQBV2OGfrGR38O7+TvmDRvNFbPQLVLuZ8T89COnHQKgiKKY0DLM4uR8ijh46FRGxAWi9nw
4gKL+6wmaeW4Igj4Zckk8pXvW6rlnYXV4zMGxANXP5zF9+pjzU9fonJzrf1AnUOAilGya32ih+Ns
xLKfUc3tMxe5JCV1y7LcsDLaKA5AXpoTu5tABFnWBni9g9aPsl2FLiXin7lu4mVYh0FcUsc3mqVv
Z9ivYfW2/3Po8ccpR8DzokZele/rHlgHTRTLCg8+hsU479p0oRN2AO/Cud9Tu4r+CmQW+Z42axY8
97OM7AOHD9HQsv6T7IH0aNtB/gHNw/OMyvTFerJ55+EPRPwCTBey9vQeZWT47BXb4OrhoGXut6Df
6wYQPuJwFIC0KpsKPP9iuL5MoPARv2AKnyVS3Ab3LOJEa8mI5mA8/YaWpYd5E8y9XAkUThq03aDA
nSn//V6dUdGr6UYo0mnnt6lF9AoNmFCTL8dwe4MN4hJ/PZKz5y1zfFMZA8k8BlJz18yLF5x7/+hi
kb+iejq8jITPop4bRktOUQG1LdbTlqGqxaPJjNn+4sZs+8+yDMPgw9Vx+Wz/6zqcLjq6d5RVN6kq
zFXL7Z9+i1kqeZvqTp6oaqNoNTvtlxbbJ/hwGPH1Iktav3QGqjVU/KG88x1d7JiARnOa5kGZDgGQ
GNUV0DITr6mK4tNX5Fczr9s4u8k9tsnjR7d5psZkKZkVw4n1x0iqFFN4AAQ8c8oY3dq1KGpax+pO
iYmKOOG1i7jd67tJk7UYUhsvVrcKCAPgM7VS2iWIZg/k7GQ6KiJpRjmvSn5Ms+8klNFY8gjYyBdi
5hds2rW4r4vvrhC+Ht3PkgqUWbTxv//Dwjd6mAlxYD0iqgbnzwBkUqTKEkD6oXtJYFRFWaMjwvgg
Dn1geUL3CvZcyRCJkqEMtOGUSxOWDznAcxb40xY6PNEnzd8gfqVwDfWfZAjEFkkWYbL9RMWWWlXy
n2kAEXyFuIF2eIjp2pzXNqT+jxhtRaHl7KE05amDYuvoaTLFTDdDKb4U6otHnkmMWMffeGTWcdLp
UuRWFKWpaKo8SstD0xurvK6LiNy11+aiaomD0pclFCvsRTR2AZJbdqgTC+22z0TfKURN+M0T7U+t
od7Pe/Zuq14GxSfitEKuF3+8/I/cZz0D2NO2+KHC9wXCu6/+6K6MMtvZg8JCE9p1WRyeAr/WuK+3
HkTg1Kn2WvOuQMpLH1YdMBt+16LjkaRTOjHV8XrSrZ8FrfSRtenByDPxR6R/MjS0xBLXb/yEACU7
5ZliMeppTj/RXFoU9a+Wc5oN8Z3grXuImMjlzwHefMr+vCM/PDm3qzL6MfceaATw4+tzIpqKoLID
maGYnM0bzD/fvM4Sm5WBZSfxRt9GqCKDMEXw2lAerQiRRYjsH+UW1bDPPzJkv6jIuf2QgIUNCK56
sI3SI+SmPPFjsxvnawOqRx635Gcg9bHizqZOr+Zc4G61yMFV3JoDtnOlZV0aRmmkFNCeV3QwDR3I
eRwJ391kO4qgn5T9CV28BygCEJPAAkdYbqHmL4I292xJStIHB42T+UP3Avn+XCpSCyoYRrEZASaw
R5lBUHy7aTniM7b2BtoIaaDGWS6Ot9mpazfG4AIuoKviHnUoCjl7FaQD2LtztEp8fdYbpfc+2AiV
Ks0ebyFEc5ZMtQjDHsyLvUg1f5kj6S6d093M3GvhINfC+0wfVq7SmetqgAWnIcgsISsgcpjKtXK6
ysP11ZatHdGsr4iZdYNU3hiHB3FQPKvtq7q8ziz9zdbqeTnLiw6r6Q84Gjey14lkfKPKG1KYDxcq
M6PqZfYmk1dlx+bdrE+h4VvcmFHh2TfPuoIGB4b6BfcVg1Rhs8BucNdHm1kDNLS02ZF4V0LnrClW
Kaia4+h+t1XNKqMFb+G9wpuYgOxag5SmIOH7jpCVPqFAzZtowr5/7VK6V6Y5g3tyqfRdCOw+wHAQ
MQN4/px6FH8RJbARsexiS/A516+7UUhjg7Rg6qh7eeSd5iwfYY+FQqyeTdkfnL2P7fo9Y2y37e5O
9nOe8GZTKAbbVD4/my/F7hnqlETZy5euQxLHoGe1T+zIYqFku7nZXktZq/IYYJ8uDXRxaiEfLYUt
nlj+u3rTu2SC1vPKhZjrzXa03ehQqPaEayAPYjSH2/pfghxzMnwC60CbFqT8/Dj6nUh7Ymho3rV3
YudLCHAIyeRcrfM+goPFn8uwNPUu6RwXUfrVyWC33dZFv5I96mB/wjnri5OW4yMs6g2bhyreIe+S
cfUPE6EdyrzmH1YeACUy8uEgDi1TRx/YvBIktgIxqyYRZsgg2bYoUj9Ejw7oxznp27thFIatO+IZ
Hj2qTdxL7XosFoPq2VFhOI6lLTBLMYQSKy3maJvgvIIxkYn/T0DUh1HO//2LC7+Qbz9sWA3/kxGe
P70oazBT0yCFkOz+vSVR0QzfJbiOWd2h+SvF+uu5sTjWrKb6NDMYV+loqgSe8Q2JnbAX7rwjOoNf
l4x+QfvxKxt6BQzUtnx2CLLDpFO2zMvL69WMjtbU7IZg9LXFBZfvmJKgjwevhy98xaGbxtQNHJ4N
bceBWnfZqAA+YIG8n/ir1kdVIl7tBFtWmMZzhVNXs9hkPS7QqlAbnH7tnw/mfnpjdAh3tiH5eCu+
fI5t0lCpRFkj8u8+VxNY2Ie/8uxwu3NwLwA4Tq+GoApeDQrgnM4Xwx40Kx1bGCUz/Mgn6yohewCD
V210ugoY7kfnkNao31eOK2ufLCLJcEdmLFtMxw+rRL62q0GxFXV75Mk9ws1Wil4ZTOA0dWmrgmGJ
QukPRYRiEAiHQafcmKcLYOB9LIS1m1lDt5JuhA7ZaFpXFl57l0RS+N7OtN9+2VI80cp6ByREsRes
VE9I0xyTvQ4xf0GX1mKkkC6z9Ufi73McDDIBWTlmexsP71r5rVzPysdH/ID1YiHJGEXUgkk1GEGr
a5UoBXWxQJCH1YlWGiL/pHjCcwHW+knb1CKF78Dwwjz9Acyk3TmaSsLdLZd8AJcw9dbriA8tUUIY
U/qkF5xEaRH4AaO9lY0/VB/0xDHJiK+IAH8jMpXcNIDcjoBSBtv+u+R4i61rdHE3kIYFLmAk2Ent
o1RPgz2shVI5bPPH1yYjwf6oxKwdOGntXTgSmTzTYVCppal7hK1WorrsYOfmKz3qFNsWu0f4GJHX
o/WCQf0GtTJrQ7s3jr1ocJNlyigbqutXcG+jvawRwuV+5YvIpm2eDbS9EkKVuEPAtsbCY8qGEn7m
qTQ9E1VmXB0cA6x0RBEI1Hy4G8rpyrgs2EX1GANB5ccNkP0qdS7O4DiwPqXslotAAL+Zg5bq2V8V
qlJRPr9DrBI3VU4eWNCtMzhbQkSMiw1thraeNAMnDl3tvkLQGay1/CAjUo8roCkwYVuYhj/XkTRv
Tjy6FhpzY/4XhHlKyiVPeWynVpR85uCNwYEgVf/Dcq8nJr8L7eWv/0BjFgdCylEHC1WEuWTVpJZb
nPL3jGhQvXjB2BtDSpJH/KVQ/Ce27PYaubqJhh25oseh1r4sYxMCkApb9G7pOqNBoHhsN1sOJykD
/VsQosU+qsGucQtI+i3aXjqeDECR7FiCrUOw2/aQgj72p2wMIrui6tpaViWjhdZsbsrF50SQrIPE
HBkbI7BmYteOtBeKtM1EP/xmhRnAdFfHI5Uu/KNEY8FrWd0RgRqkNCXKGJ3NDRged0u/a0KFKXIv
lVeDwoFa7w6P0feG4Vp0n89lyAqhfWrkOhTVI8hCNEpv0VimQaozeNsLABHx/qCOlsgLFgR30HIm
F3v5S1ug9oPG4BfFRyzhiNC3H1rKHDPdIKscIzJaBNf/nShVkgQ0Q6X/2ua0lcmAN2bOYVNywYp1
brWRJIcSRj92z5sImRx9ltVUTqv5V2MtcSmLWFRP1MTBxVLyG7q+WRc7vZgLLILL+Nkn/B+vCoHW
8ht8zX94wPtVViZIxVoFYEy6A9DKvp3wBO/6tCqROln/dlmpz5Jqebk0RzSNt3N/R+sK1ae1oHNQ
BBVIFKJQY9poOF+KvMJYN1WFbVrFFbmci4mbt4CwWTnyognLRqkymcdxEyT5BsN6lvTyVbuDWzao
RV8R4zzH6Qgd6PtoFkfJG7sJKbJ8o9vKUaoyq4pW2TKMq/du9bTXQiINFLvr02RYb3bddoEDAav2
I/u7LkqXSg1wuAkftOP7l3np2U5lF1j+geX6872bQi+M5l4SRXJ0dK/vk6C0N1WXVvGfk64wrPP9
NOcNzQMadq2ARj/3z3300s+GotpDSnJl+/YwGu35gZ2CV5wTJfdOtD24/yGXuY4Etr1L+cGf6TSj
ER8t6s3ZZ2EvVk+4ocEaCkg5dWqyuJFhM8zEiMD9NLyDHS69CPzdRidPkzGYk4tOgj15CJrOkI9B
X8w9w9fBRQZAROcDOeCu/m95WllqxkBRw8zQKPum5JfpTTIoM73GaLtAcbsXltHopBvPzEE8JgDL
1GG4vyf/RJRhx+Wd/js1KQUL9Gy0GZ/PVpDGKB+IMyeOSYBBGu8SVWGZbezE/Tg70kO1k+w7PBvg
f5Y/5dEYT5g6FWOihRzrwoKyFmL0AN9al6My4aiHg65QfqREXzBRjatjqaQTX5DowK9BEBqrqrz9
PnkuI/p7tSh4BqzO0/gBdXRxNbKxD+i7OR0TAAk2ATNp0tqrPj8toAsMTx4bOnfQgvZfDqA6AjTc
qpEsP0ir7Rs15azrg01zONjU70kB9Iv5Ir8nduu8mRyHtz5egKyKR50CGAu72Qw5q8z999QfF/ge
1uhObD8LcqASmlGThJdBEKqEUKzkPKxL5qFUSxCwvmXXA/s+B8z+CRqYi9ODc5ddM18iEl3tzOOG
65/4GnAOyMwdyGV0yQZPyvmNxO/J0EOwIunY/JPzDEFFB8UGpobQ/elFfqZHJgGNqH2Wa2T7YliT
Yb5Ta85J9K/MP06nVoxTNDIn63KzG2ooYkGQoSc6m2EzBvEqUdmhxoXRYjkei4BNr225X9W2cG/f
DTCcRqJfwq1CEzCkRRsoKCXDMnKlm4u5dbWgqoRtfUPHER1NchY/OrZFLibaVCeoaiwJrNewjrrU
kGNFoJlT7zfTORIiFRKGLqNsmfJpj8i8rWm65BZLJ1viBMtE0uNpvY/MeP1rOaJhhpTyMh7XKI4T
uKfUWQou7nMsFkvYaFkBl/nHGEXlefpigYxD1/Ug606a1KKDQT6kRiBx7AZzObfUs49fNBx6gp5p
tk679z6nl+FG3gTjQ4SGefRqYqKM5zIKr5s7ZzStCL2pp0tQD0GI+1TeDVz7nEOiI+OeE0ylnG8i
XmHU3mcsX9+pgtmh25sq2fQGHxyvJ0WmQVFGcPH7myCxgy1mPl9PfZzk03T0oJIQ3Jqo0rY2PSLd
BqFnRWar/yLkjOzcby7AXFk1ME7T04aKMpSl8lW9uzlAeyMvVy6cAVNpYxV2tROKZ8pG4fys5Hla
FRlH62VkswPdEKPGmuuchYZ393GOO2XenLN+MviTpghYPB6hjWHrCqDlsPnOAbqu7ScOQGtNf/G7
YWG9Jh5wNY8b81nGh8mAJG9UREzT2EwQlQjzju8pXCPi1QeuUeVV29hyIfvDM67/Y8pZBIZ8dxNj
OjTlYXDiBTDDSmsunLbkNMV6WFDtZcfKESU7kBji0Bbd2BI4QUhYcFZ/OfDWpgqlmxFKuCzyl3LT
RhbFH7H3KB193VZoURy6hFGBhZuCASWD27HBIAqkKkYqIvBuO7+QeSmeeEYrGYm+i90R9pFZBwLr
Bw2MQcgWfqr0Pq7ph5b29DCEWBlCDF0jtCmkipqr70+7d3ww9hPbps4SyEMy8mtY/krZBS1B6+I2
1c7F+KIX2Ht+T2YMxsDfVQMe9eio2MXDPDzl448VfoDPpTv+On/zvV5jGgN4S34xmTy+JXTevW6C
kGxJgQi7uBnmwQKAdpigsQmA/RZHHMybbhv9g06jZKnuJQDFAyF2FHxGKbxUnQxOCAAfP007ZRZt
Q2DC3bFY9JHr7mKybJYFh1dyn65GMXdVBDZjIBV1wTW8AOeFf7usXQ8dsElGKFlTylBcmreVPS0b
YrbazWxSY6j9+TC7Vnh16cspgkAZGkgGxmRfazxhaBJ+gT9U8Hq8q93rA++jCFBgcsFZ3NqOilok
/7aMswkR8krYt+44+0ZEsPjG0u+bekO8v+eJqzuI2UGSfND3O+mIhsMj3FcsdfkF58TZWjR6Ta2U
YMpFLyltQ5lOPGM5V+nHiO+PV756aKGsLF71QEr5XuParp+I0B6IAmvbGRRI6u+p3Am5FMrftIrI
zPRrZwkj3bdabGEdlJHilFJdMlMjKXBxZDjk8LdnwyrM6Y73nn/4ZPtQw9AAFY0kEGe1iRsg9UMs
4oDfSCv8madPe2s55SJlf7ZhXoMvJu2utoGIf/9dOxAoqv1ytd9d/Wp2TUh+vnyMj1Vbju0iW9gW
OnZEAbFsd/20JaE/SFWGZ2rJNqk7S7+Fh89Np5fO29CsqDbn4ZrpvsASsLCdkHSfjSNly4cJJEDe
w5UTLgDicqBOJPONCigqIu1p5Jc4PovdjHKp346fDiK32uMtkNrLF/B4nuNFVrc8LZRU4I+0eIcg
UuRjUaVIwbYQ5Z9uRoTUg1mI0sqkzPSuoPKVqn7t7/K7ciV2DGOQQzt3e5yuXIVAsYt737rG6S5v
OmYq9xg9FKkGeLUZj1xAARZgbQu31bgaqmsMUPYpuiIHBSu7niTUOhWjmoiFC9gmIiQId6KbnO6O
05vweMJ68VJgaQmdl38bUbYBKCsG5BgODKUPcFodJMQhejJNcOsyfe1l6jZ8wrbAaHbt7iXlZRme
0SzWJNVhr/LQEzwLpPzvdKFs1nMRdgk+toWixRwgdBwrNXXK9mRF19KXoaIGm9DltHjT0BUMcWSH
gWf6FmaIqtmtYPfmOqS3nGwowuH/Uz80B1+XDWnR8sdRaNc83cZlrI+h1rU8cvNx7jkvkoHwMT1h
m6oY67B8HWRxcNPOntTc5EHHTRfex13YClzgGzaswtKvHG2Dak7cyvm+Sj2qDsUKDRhuCNuqeH71
PZsUzpB/dXrfZlxCaF5D6m0rKpBfZ0Z2PqPWZlcE6sRTVQhjV8i4Flx+IEe62k0Ev5eAnyW8p61s
36X/+UCJaQ0xGdVbD4CNlsjpilt582FuYLlc5ts1x/yc/NFr27h67Worlx/RfmM5WXvklNPi5Lnn
0c15kiMQnfmZDDDonLOIZ8nO0wm5gr/Z6laXRpKApTiEAJ9FmR1qhqYuq0LTWiDBXSl3RqaJp7w2
25UAPzf5s/QVO5iPQxJehVuClPY8XpC2mvzd+r/ngNNwRnL/+0krHnkEZDPPuxs3SP15tJoYwlze
NNRqtBxjhvXI3HtFkjTUg4cM8iqlGky3A/FUQMvNUhByYaw4RJ7qErB0SUyFTjprfwF4Dv2Fspo+
rfNIykjGS+AYKUNDsnaY4kGJaGmcyjcDWeI3csIFBFRucYv36pp0w20W8eiulFUkMa9gAxvw/qvK
s9ldQM7mG50b2rPAIbw9BKo1I4iRGO7XE1OMpOsjpESUjgdD3IveyH7/2nTtXZ4FnLcjNOhMZoqt
ZARCaGAdPUqRxHoICFeTm7U1TMHbOUAV4VESZQits/hyFmgVKHUt2g1J97XRKN6+AaZ8V+/A78Aa
4ljgmNXAMY67dZ7dlaP4U+c8NiSSWm/l2YbHVVmaB//hL5UxPNJoCjRvIsJQ4i6lVveiDSfBJ+36
dUsMRrO/rQFzl9sq/roXlhnohfx1Pp4sm3xnHa7hRKGLExIi8br7qM5uetgknayuZNRUninWJyTV
o1DecGjebfaNsnHVStT8mhblT37g1Qn2N0u1S6Jb8/hvH09k0dxyi+rNwJ3sThV0vhYqCdMgjGQy
CuTsSx3BJ0EdVJNWrWr2lgg5sA6mevgbfheTqgSCTKhhO4lvhhub3KbZOR4MVwJF7TGh360c64PN
Ohjn81eqxcBAtbB3TzqtqKrvZxUFCmL0SJDZRCGSheOBwUFWYb3VW8kj2LsUGwk1jn4N/crFagcR
42pXaTpKM1VLbQMAbMAWbnffaY25Kc/uVufwg8BLUJ9JX50Mg3Mkz9QS0JE4SUGdf58YzlZswcmT
cMJQzZeclC7JEOychh4GE1HucLusYQw+NPF8ac2q6kgWH5AD4vrvh17YxdtHEsjYfjQTWW7dhUxy
WlmPNvItGohlbZSurx34m6dBK8oMACNATfYKIWl+kI4ve/v+umbOFCwKY+2vHaQ4wnh822ZBNMjE
cY5ZQsHGoO9tPx76CxAIa6vV2XnP0qwPPR9hqkafMZn+rYbAkdDlFcO3WQAGro3X6JOXluZPsCRY
++VDqXbKroD9CgdtQ9QeDV8mPeRSGiHQtPkkolK2nbOqevj37uGjQYqnIzCrJI+u3n92jY+pcgDU
nmDiiTKU645aDnaM+TxlACUfejKT9UPtpXwk/5KTARk5o5DFxHWIRzADn95sxoihLyxLGAUx79Kb
5yQpI+fuVbzzcXIknentAk78veuBwC51gXY5TDTzTMBoF4Cwi+D4YgM8EbPzlj2q6dVPI+/anYmW
PbFGtZIaalxoDKlnAMKtsb8bCt2asFzULEFySPn9wsSZjU+ej5CUVPfvBVWB0HED5jz1uBRBbo76
fYKqghWds5KUDeusWPiT4OfShYv2js/PB6HmOs4hksuUBvLnGDgutaOOIvkLCq6aKuVOAVwyDtYR
CvRlUTtEjOBwzfBOxlqppwBfUoJiBy7Ax2ubCTO9PhS8DrTUbLbQ8AsKoEZzmHgY8kwTEYnASKUB
6VU22H/09OhufIcJxKexKJKq3YIFSNnjoglP27EZ0GMuspdakVS8Bl27DdDlh/imR82QMsURFX+c
AQHr/swdjE8RPXO2oXKlQhT2Qt60DxO/7gCxPEhnxkmY3JpnwXZ4cyIe7neVq/kGnj4OmbEcufGt
FJPU0ihT8Krsda63oG/V3u4PAEDvxtnFFSH4SRCwgKlmdsnzIQdgobiOAvMG55ows94FEkLYE2tU
6UINh/BYM1wdM9Rj23KNRhpeUxgxKTDnuf4LGtms461iK/bUo94RukzMyLE8sbVtwiG2bCfh8aMJ
9vqdKrlKsCWo4sVbKnqVQ2FUzPqKVWP35cZ8lYzgLSZhRPbOeVGaiK4Ep/aemgTZPCfh2hZhw+Om
nZX0gnCVlxrLyAMYn6aiFM93QQz4Y7hu5nsYeaBcamplE78lHBqsX6kR2fTXtjL7u0kueqw60Jc5
xFA0McXdUo92LcA2ZCGwoaNbcRemnBNsHSGv/1v+ENo2x2JULKLIEUAR8qLz7V42w1/vAH70q6r7
VTRDNGBlFm1FMafSrDnMxH0jQ7BdKaMNmi3c5c/huXeKxIR+DJf8H0Glp6quBvSFk6UDlkXBmjd9
V6fpAI8bJAWmOs1Bn/dMFzRUyEU8EzpK74QTvgNdkvf5yVH+KzjDl0bpmnmWbpBlgDYxysdsqNKI
Hfj/mGFnzlSd9mkvG/XIdG1e1A/unth/aGSTze8HpVKwmCREo8ZKpkgZyIQyDvYP0VaWr1C4BB/n
8LAyYWIew4veU5zQLAdak34B/s2RVD/prHuXvYNTIuzVVOv0ATrWfOiLpedvyb/biylVgPi3Xjvy
xwPL0Dyzm8pIcWfrp5Ac85SocoeftMy2WH1KhsDiFddl3HdjCpC0CKG4wHEtLi1Yl4HL4McXymKQ
6N74zsUruSuycB1DFWIcIAN7qQzwn4/aZNUvUM3SgO6OcY+50RranP3axU67ySMyDU4E6dY7mD0D
/Rigy7lyfgEMZq3cnGmY/HdaqpYo9Tytpxye3tKF37mG2e91kwaogpsFs4qXaDINfTqtePp6be5L
KRKJutYNp01+EBcSZHJny6Moils4FtlXIHf3lSgOLWL5/8VXJ708zqEfde/XanJZfrr3VLUTDZ50
HIqQnnsy5le/s2MBUD8Y49PW578HVbN4h/WeJd8X3FtZuMBlA11itL9ZkP+d60zsp/ti2JFraVuA
wz/VlVAQRU3Nlg4klxY/BkMO8MnWSAef9qSFs4J3wSf+8p0i5LBUaPKo8Mqy86/jdRmzQgMpx8D5
YY8r5uM80j3I9/2BJ2qd1oMarKdScHgmfXpPVMm7OxkuCsjNF/hfAOrOmKk0F1AewoKP8Q0+HSTs
a3oMLJrPWxyTNFgPW3KoiTJ6czGI0f6WFaC8GE50RIYNU2RoQv6IJUntVOLDcr9da5qrTQ3UROAp
PrXxbwxduKgYwjesqH2M/vyffQaPC3SgPniucZ0kydBhlGtyVTvh3oJU9SRpSZeERaizm0z3nRcL
OKZVkXifQSzHPZUcZewUmStGz7i/k1vhTFeRshsXy4Qq0tT/iCgLtrRHRzzV0YcZt4G4mDYBJI/Z
BJ9/54+eXalVzvlIcH+RcaOje0/viaNNIbhpPGHOvk430Qc12vkMTQJVDd9SI6nlL5zU7+MMcxcG
mnUarNrvYy74wyYGyIBSeC5jp5osA0/A/0C5wjQ7QpLa2urYAjFwubO95w40c0qhiwERM3ne6om3
HYU0XMWFufzReP9xs7SxV7LRzfSLJsD6YypAcLaXWPQRhPAjsohkmOfM6z5JSy3RCL4vGsb7KtjQ
MEwE9dhk+BzMOlz3xfSfpeObqiiZWp1AATphfVmthz43rlwWesQw/HfG+JAKaO9LCi4dXfVqOFDh
vCUwGZXun7/I5wHiVCDCkMxlWIY/Ga19rlrFdUH522lazrN2EytPYUd0XliUUWEGE1+kTMyvDm5t
X7Oltzaopn8m1xBjdW8mit4dB3ZaTi1AyFpcUQMv3CTX7yLyf9K0JTrl6ziTX+WW/dkxbgep2+pl
3TTKarQ5itOhrOz2v9vTFmw6nPlyYgvDxt8Slhj7eyJeOJHyQNqBu6xOoOcM8Y7RmI6xKlJ0Sw6C
9UDQ/lNmBmH7Dm4k1iTs9PrZoFjCUhKtY0HXf4+afm9sh3roM1Lae0GPk4LRHXzW7maKBzrUjgjx
K/oW4wn2KmAFIWwYrV0u6/VADoamAPbm4p4hkQXVSIadasIiFlQtHSsPhqUZpVLzcsQ0GySNdiyv
lrRXJQDdmcixwtgFcDk7cfh4kSE5XSrXAiqNyRhRJC4MQn5cjnoel9lT4XsmB5rni0X58Kby/l/A
xxrU/Effpb+DsoTsD/Ku+E0dibZjwxzBq+juF2xBI6OIBBQsBe10CnvDgH4QEb53T/NE5kXQRLN2
EiQe0XAphAlZ0ypMsA3KvKcTeHk8JOUKHzLb8t8bz88ne6C6/T65ooR2IMqbBASJiVAQhZCF9WMY
OfHlbsSycAnFZwDTxY1PYOBTzCJow76J6VzpWRG1tPVxgFmYBCGvhqo/aWxhQfCAsKQstpNLDBAn
xmzqbN691itFvOg/AOiUhvFXjk8P2dx5MltULpd2MBE0UXrFYoQZVqniLJcH6+DSXOTOWsgnh7uf
tXv8qdBXA+x+L4Dw78Le8VEgb0cm+geu0F37Yyh8HGK8Vq4Z9PSmEILAPyF+QINj2rfpJp9Hamk/
w4nzC2A9I196QyxWN7Kc7gyAue+K4GjExwDbdgkQEmhRgqpvvY9UsEBlyIRIlJqlH7vb/qMoxD2q
rLIjExilQM1bS1A3k1Y1eA1mPpn+2uj3RufIY45dk54Xkz2busGRMMd3CpSD1EwKAx4iybtoYT5Q
7LaTS+X/z6QFSrFQxPWkfqtXFEwLpnVL8nqj3EaS/1O4Tv70/gJ4TK7nsYGNoA9qvovJuRGxsza1
j8QjfZ3p32QuKNk39bfSC+CXbYPoJqjAzZm5/ulemwl5LeW5B7xL+I6PovpQ+upgfbgUZ76hH0iJ
km0ZntEakPDrORb7iJUFcwVHSalm7Hz9JSkduC0NcBmkgZxSJF/qerx5m3FVewsUo9nNGOC9vrcb
LZ8r9X+m5v0vAsdeCkjFp9dZ/c+d0m53DGNbShJKwgxW/H2bHPq6g3B42noxZHCy5ofa8Z6ERYzE
UHkqvT0j4r320b8iZqnbtvQoL94M5cDgJtRzi4pkRdUS+KwssMB5ZBLce219f+NFjJa4znGgG4Jw
i/Pi4HYHS74jTyQCi4UoIm1BUSmDjAamrTfKXj4msSTSVFIhPJn1ITVdSrzguC1I2sUOtyKeMkn5
axK/ux7l+t5lj5enFsP1rkK2EC2lGTQNQJtWVy4SMheeeRCIWLC6cWufp729+MSd4cPossTM2Weu
tQD2hN7ky5jMPBKgfCPM0Lg5+QMeQCbQeQ4XhzmhxDZz/cdwmpLTZm0d2FsUnjnjOJnWdJ0CEqU1
fkVnHMwCpAViVDr+6gZvrLx3WKylZEvJnqk23MrJA6Fwqi0Cb3VuYW7NZDSbAvXzw3PurLkPqUdv
Rt0NUbhOZX2rXs+mX9l01OASh7iRPbwFyBpfrOiyMNgTVyIPDwlrZn1wnEnvCjna7vc4k7J29BZt
a4Z1z4uXxHSkt1+S4uz30z/ayRsjViC9gEaLRKhRtLPjYE+aR549Pqcw7s/YGrqm4IcOBHXF8TG2
mk4M4QOi9q+uiWtlU6giRSv6kIz/8JXRq76qAB/JAg7a55urkZo49avC93uvw3nRiTEWNjsH5zVh
r088uj4QUrv8ZHwa/ZvfYHp3e7ALStoV4DTqA1bVeaHuEbj9C4ZDKe8ZZHKzn2Yn/pR92u7NyskP
dZxyriSNCpFMLMTqmPn+sY9nQEw1szYT3ssk4W4fmtDh2WBAPjWlKMwqQNzZvIIjnAL1FmihZq2u
lRcGDJ+2jE/Q/yFNW2m4L9OHbGMe8Jv53+hylU2tM9tIdI7WcSVxAH3mkahIuQI7b3RYK2JgBotN
E64lcrbW65wQYpToxGo2XMGf2h2iqwXmXdtsGOi4nf9dNdwUrSeZOVqIf9RsyoS7TbBp8IFRP2QR
LbolQtBj7ob8bjVucFO7KNgAepdSUSaiMyuukzClemu4ua5bnJchOaJARvancsYWzqkFKK5LP2Of
GNAB7bOuqIfMpliWIfc65D3zXqLsj70TFqzQXlHL+gbz/Jl6aNpiVjDUzbwP82ZVnJFLGX3OA8SO
ayZuTcumfYIT//UN6BYJY7cL0Co92dMTYUtCMMkkoEDABmy7G8RFBpSYAw/qzzwWYs6EwgVu32bb
uf2ApmXD9K+wbg9XYA6m4/qdFj0CfyzTrGZ0nCQ0+qRWUJHzJZW4pfwrhViFfCFVxlnoyiVOfuqF
bph8mwmwLKYE3vQnPZywHA8SQexyH6b8/XqXhMQbdVuiBezeaeA1/It/uQByE2MPBD6BmKunIJpJ
Yxh1PM1TSRC3eEMOCL23SXb+ov4Iv1mTrZ2sgz7hLSBd+iCVKGODIIo3CqqXTPuwCiulROKD2i1O
XX6VTBPkFG5+OeHiJQ0JuJdQHU8+oVP6yiXUBrV5tWu/TMWLoh28e5b1k/USKGFs4MWhsE77gqEN
KvH6ugCpXWGGfuFbw6ylKnFkbKf6xCNbrLn+51gzgbaCtXbE47KjXPUoeDFZi5icc63cU19boZXY
uLtLYFCyZn4H0DiROtXiuYIEE9ofqtDScARc7u7mUkuicY2MXM3+/FKo1ut2Vsart11GHVE3MPnw
/k/iDS127u4EuBN0SniGHlOLGfwixbqtcSzJlY3AdCKrL3YFhfbh46TYGUvU88TlGySVazveMSyj
fMA9hp1Ku+XAilSdWNc1j2yvNtRvNZvBKdqfEIDR6wU+z0HR124qWK6FtSejeLQFVtpkgIXX5j8D
Bn3imVAlTDpwdtQlSJl/94DwBINC3VLaUgIlSoq9QTfhOnKT0J8fH9WLIjNP+15QxEcW6rFhTXDT
AqVrAyUqcqT9JexERqxz5PI4fnqPYXtg3n+qdBKdMKPUB39fzutYhOzzMQV3lxjtFoW5ZTm9MvLv
hkbSlPiL7skSvW/4v/F3zYC2soFJBct0F9pAt+TNDXUm4NzD37WU+N/FIIWWeqepquyYaLtOX+sm
PSqtfXLwSL1yA2pAl5nvtzyzub2zBhYVYw0GeTOIbCy5dOwX/HJkvHLa0D+O/JuAyFDpgXX8i5RH
f3crnpAJH4tWOMmj+Lrku61ZloMj+hjAeFeT13xEozo4g8/4vcbnQwerDSRWfQ/moGK2EtpUsUKr
A7BOJhA6ZVzv2F8LGdNTWoAbM6raloIXkwLrBUu7f0D1yE6EAwkCKMhLKW/UaBGieIA7I7TgYqVB
9MEJEijZ1CKXUzUOADBzX0FafAuZPD08F6iGOPGUbS1B/7ADZ3lCHXL2k5qdxMM02p7dYJB+7jcE
l8c+5QkZdgJC+DOQAM2MbuQg3rUhqZEB35BJOry0aaDRnhvoQJWhLm8aE/Idv89+pIETwP1jfsUM
Xjw8OYNE+8yt9u/+eWFDK3nJv61MVU6Dsot8UIYZpO7AAS3y6tkBJqKph/KfsB70HpqUzoI7JmDC
GCQNxUsMYxqUp/KiBk39RJ3Zt2YktdZT7ExWp6kBptYZwXwmncwl27G8wR+MGgf098aN+V9bYbrS
pQTm1qDdTVsbN/UfBiczv6Wz/ESoibj2Z4Guc1sb9rCZfyHUz03bOUzVEkB7qmcsYe755Q0Z1oX6
KgFo6L6x2CgHEstqLiqG5yDWK83gpziuMyQwIayU+wolrWfDWnYdnqbww1KFDPuNrSMTW+h+6E47
7nLO8KGPmXActm2mM268ayyc/F9EH6A4ZxjcHEXu/Yn7buylZ/uHcAZbHcgZhztalQOhYAHg8c9H
5tds8Bdi+8yx3YABWD1tW+lTejHO8Vyr1EwsFRtf5MG/5TOC2sM5q/AiPhjG6NcehONF4aGo7lr3
KzvTANk/BuEmXzVfrQCcM4JpFT3OkxMVAe3zbcVeFQbkhhgRfNeJrVt7JgwRh+LAuM+GFPHkphVy
RiNrEZ94HBsSgTRWpgZhEKR8RFQNKYUf32uBq2sNYVMPeimJ7ZilHCcaaO/4b9bGRAZv3mSVJkfi
0KVwquOG73sSY6E5jBMZdp8peR26VReAwbAXkDfT+tjgjQL5QlWy8XVJFjA32HZ/b56sSd8zTJD9
rZJxu2xs/0X/td8vts3m2iTl+r1PV/yrDxJhqHsQSfDYW9oOeVuAAPHEvJOvDlObXINbv7hKfyQu
tGKgwGxrieGct9U3lJrQ06cRaApkrgcrkmIP/6wBtY4QafJeXrYBujtwgYAXZsFvZaUbF8g7sad0
Mgv7HMYE0Rh00OyGDFD7Yb1rYgZrP+wRo3QSbv0cZNkptegzsGSNf7sgOvaWfn1Dr8vH3m05SzXJ
6/yu5dinEyLLevtkVQv5/GYsYT/6BEcMFu/55mKYfblvDI37IyOMUT42NelPJyZzQpdGM/4sC+io
FdiBABJdbSklAX16D+aIYVddsdqqmNcWhB18hmTQTHuIpJqClPYNnomJwIW7lSQ/eug/HsqFTeM8
R8KncmKwJKup7v4lU4+/U1PoIvni6glru7OgiCrxxxU5o33EdQAjARsO3wqZabyGw2VZOTl1Isru
qXcoiOIkjIvsiNbVn3WzZSi8ujyANjI/50hlc64e2bjHm2KXDyI8rPqidOvT6eTg5Cs34fSKk4hr
c6f3W11vSbQpnDe2ZMjkhZRT03irXC379aMXUY9mGrQNObrWTWKi4IwnqdnZrgmpJJCkg8uPuxBm
WK77jFF5DaJPs/6ETle1iUhdWrbtwJMEqXeUC4mQNOrAfNhEvXak+lZYGzGzPbcUr00pB9jor7Nm
grM4gDPoTLce/qKmlNCmz07XYuP10RqImBWroX7mv92Is9grqPNn0ACiol4IkjM8U3x7Vquu507M
A4VyfTWwBNU1H7LwhoqBL5COnFDPootZ+5UdTRK8499iJU0ZVW3rYiy5D5cQZe6E3VMhZM8gVhfx
c8E8UxyGPzFlcModVt6B3hkozT+eoBX9ZeorNIeMTAUnhxkMcOkndoLCvHiAJa4gs2Wr8tKeZoo7
RbJpLtcSRw41f53bUSjoCfhheTo4NwX2TL9e7wkUL+tQ1yCHNuZtwhrcq6Gjz5tvowIyjNMzFc2w
loCzoZEZCt/460AyIubQgKFqLCIe7grwaDM18AhXOK9IJT2DP/vbJh7R2wMFDdJf1ebWTwyAkIGk
wKUCuuSgrxo7yrbT2BhBJh0smq/KjFPXMklARXvRRhKN9k0ivH1dm4UyCNlIo5ag3o4eFXy0w2L7
5EfgRJOzv6PnAsqFUkEKCF4P9pOGgGewWzqJ9TTD9CQ0KaczUFphONuOfcQLa6sP1uB67NSag2B7
3l+QvbnMct9TBZK9Hf3pfX4EkZlOXcvUUMtnhpUc1Ft/36td4d/3W0tYHZ1tKHyThC+OzSL7tgSS
zUxRbNaN2f9tzo0tyn7xW2jAQqF7mEwe3GfG5R/j0Ag2hpDNM18u4Xei+izO+shaeyq+neXem7mX
TKuYluU7/eb28zEDec7UkMdRcsgLKR0xWhLC6KNgR9oHlYYlU+9iEdKeh2nGtyJ8JRXr/Y3knrFr
RGt0DrYykTvHeoOQaJgRqBz1kqtwFakoDDsHDeubAHwvU0yAIgGyn5KKPJExeDyRpB4mriZfBFsH
h9z9ajD5jtfvdi5zvvZqlePlgu6irU0c4T5SscoOTafmtUsX23E9Ln6Riubq96Pbt8CRHYGGiejt
OI/OsxBoxm+jAwZMCMVTvdc8+zZWT5SJeYnW5uYl0TiYDA4BgIWLEk5rLqhnVA9HGO7pTG6BxoJA
ShV81Pw1iOO8cFt8nW/iVViu/OeNUzk45aPCNdjTrGtdhL/yGTSxsWv0wNhb7NHXbaKm96X4XF7v
BxiEHYedJmWIYZ3Qf3eHc2GjHYhNxNkvWywvh4NAyhP7OZS2hJD91yh7s13bXkKT7YcH0UdwKwIH
KVO4KUxbldkPFE2ArAFF32BkAQxH/s9+YmM2kWTeNTmE22pv3X0bSyiFhqy/7fV8gJf/wLplwRJ+
PvCOGt92N2dHVu5lkIxqtxq2J4JB3BKQ6GTdRQVEbrLKwzFJCFM+ZF31h/j+fr9nVGDBo98egSCX
Jyxn070xOlVkptvRNruFXiGkLhnim+kk8W59zFb9c0jYpebu91MHADGwb9cWpNun69hGfNYvRnA4
keGs0FQGRUSd1ful48fis6gKbq0WWOGIenlP6Rq8v34TD8c7sBN9eNKUu/hReShnsjr37Czs/6nm
BcUEi+IQPty9cmF4Dd4ozlosC6rqGldFFjhSXrwE+fjT1ma2Y0C9iy54ukT4ZRXpeLMuLius4skv
hflRjrBLfLIyAoPo0JiL+oIz3q4dOKJX2r7CUL3DmuASLoAUxoMS8MLZ2MkcaFki5+XKAfnR3fY6
+7wsJcPmr9+9bKV2HUVW2/Hoe9+zPH0WwB+nT0TSsFb03PGb9TZYM8asxGG3aeus3D7JRXCd1mSu
/Nzb1v3/eW8FzK8fdpjkTH1SRZ2NZVEmRmEyUI5k/LDsGeSM5G+RFrsYL1mvCCk1WAKiyCeme9B8
k4TOIa/fJb5ySWsCVCU4YAEgPwcp80geglCGKZ7sIgKW4m1oqg48r7rE0ab125omd5ZrTIQFgRoo
UB0mafBKQ15Q+XbECZYq8NSj9902XI6zhwzqhrpCXW/4UDYsy7+93O/DHlfj+U/ECgjFHcBibU6Z
tkcBkmNrcK1uyHRO2nNLkGRHMKYbj56wotl49NOwWbjf6gqHxjU4GuRvSn3IJd+wH6ZQZwc6xVT/
7dvc8vfpD5PxVR1UMVqNzoAgVqkA8ZXjlFnY1QtyaEDD4vpq+dImRDG/xZZruUDJ0U+BBCMy0z7y
SI4kXuBWv5GsVlNo3s161MJF2N/Mnuz+WsKtMVnVN7DpmLEd/q2+aR0ZA/owwXAkSLqQ1xg5l4iI
C9mHD+OqsK0IErg1ZuR1zbKqNAnRpGv5UqmDrrCF91fe1BLAUuncf9Wz8JBZf7byMiq0ta2a1g7E
nyl5CP40tpl3oYozYHI/F1s7ZCJoW6iA3AqFBCjOZC+cCUKuLtiQ5U2vgWYuXHH8qqWxVNXhbuyB
UcjaPN9eTiFl9gmClWQ1HBPkUudjuI+eJWzCTENt1s4IBqr/EtK9o9+MDYgbPZhlgP4PkSK4YRGG
XApOqCPQPJC3dUKiQO8DWZ6+gWFU0Rut4P0ts+8H6GYL5USsswcVB174MzIwoGnMCgpgzT5dCrcA
5eRmnsDk3/OjOvvS/763Vrg1mbz2II44YBlVYjkAvWFZ8WO/AAv2LCLERCmKgb/NrQxNjxoaw+tu
PN3C441CiWDrKBPwmwoosnkDpFP0qAmm+kvd6AUvqKWzhBnFoqLKcqwHF/4Hj4TZzmX3Na1m+ol1
0e6zGlwkXu2p+nuajcZe5ReZ758N7uXILVC/wkGN7qXuwtr3AntOXHfNHh2HIuJlcLMO12DWJPaX
8CqwoAp0I+/R/t5nZAd4pnBGemD2ievcfb9TP/noqkAotdPOJpIsMkjbG12/R3DvULeemf4PbYdm
Fo3lYK5MZ+auAnjuxBtZfaHYMKAfsIQjMSc/mWUEZjjxUp5FE+zi+Jt7XIpQOwwZjvCRRiwHeFlm
cdbaaEGoy9+cR77j64QRPiv9of7KeNPbDrSyCZ/EOJGKUpbUk+FJ61ciXTF5ziS+Jxa7G7JHk0rf
/sEH8H+NZ5v5OZpldEngQZ9G6+PDe+bBD4u89M4tk3s9cwtyLBoTqIlV8xk7IjFDwJ345B5We2oO
FQN4ivBkIoXWZhvkgf/5slAAjTTzhc+mKvx95MQy7Lq7LLiyxzCjBB0oYS5edCITKJTTRHimVWGP
b6DvwrY6b++e8WqXjWcShIOZjlqUpyu7sBHqd4u+5/JkX9bw3LMwYjIJSy8f668w8eENaNqHaqJJ
YTonH4ows4Z3h63IKvy04YZ1bDM2Rwx2SC2ntkBYo+B+UxcXAURV9jMS2vBnNl+PuYff5Dzy9k0x
vZ7viehR8yMy1gzno+rCSY4c1RH8ioNqsxIws+mU2tBE8Km9A1wQxb2yFlUK91YuY5f2EATxSrEQ
Mq7rmY1Zd1uPmVQ1TuhC8CpBCyz0poCgBejrLjEG4JjvYPzE6fBM4dDvd/lDoQvLMBSkUZLHFzhx
sI+mJe1g2tr3YtFr4TD89qeYxEq8y7tp6q7uc8Z2APKKWcj8EoFX7Tew0UiMapbm3y8nWtwwll5I
pUgsPUKNLO6nHOxLl38P4CqIHZKLE/99jaLullBm9CjFDnFbrlYr+XUcrxaAYPAur/hFxLSjsdsr
dKZk9NfFv+CYlb9yJjdV5EUhG6lwrlYZSwN+H2s0wKtAFzP63M4J5JBXZh4kKW/T1ihL9UaG9NxQ
21oCRh103oMg67WqO98Jmdi2sN43/+Jb2PiBjUWIKmqA7aXE1OWikDs2JUbAWgFsgZ8seP96ru6f
blyytyIuRVghQxRXyghfdVU2LHPcmCXH5p5AUDsO3MC84bbdDDtf1Dc7ka9rPEqsAYdgEWBvr/y5
kBZZkaxNmEFC/E80V5Ei1eVVbvhnnFO+TUWTuXxFYkIWLRgEg/0r35JbysAPWshIZD5kwuthsDgM
QHjqt3U2PRTM6JcU61VJYVax3LdxpkqywDnM2Zj79DwfsxQEh7eWJEX8rffcjPDftCDxcHLXk1PE
jBTgUzlvIKLKIlp9uG8+G9Bsg9UR6PidAxpky58TwA+A1k9pTGkcHI542MQYT2/gHSUohY9Y9bnU
WeyBH+/sFbOEPJFqBGMI5jI4kLsQSZpYNjirwDTjEHu2N8L6vE5YYOfVQsj++zq9A1m3U12PHXQ2
sClV0G7P3TruOWpyax5n9BQJhxpvgj0X4EXitUN3uQ2hbmVxTGXQ26V/3B3A9bHc2Bzay/pyLAHQ
6zT6pwDE9CWLZ7PxvX3rYN8cUbY6EbOMd+Mc/aufoYVDbM/kX8jBqFPxKb0y/zqHT7dveJ4zI1/Z
qHK0ItyqmeJ3+IJl9CxmK2cpkG6BRIAHrm3tPNaj4QLNRLKYwjHv4PbIzKlN1NEmWbsdp1B9Ympz
Ke+OcZuHaMmUwz8XeBLSPfLK+KyWtPH9LQ5MGg+O8O6/RUjZI8Gy9IC/jI9kcWwGXYulUXvJQuY7
uPdy+QGg080IFF2YVHGaEUeSF0G564rA2xRZsRdwXtCbuOpSfhtXGq1Ktj/sj3MZycHCfPVVbuw5
Rsm86pX1voOOmet65XxsHnvTFs4OL0dfTEC9yjJatwXrykjo6slfMik264eH/BC1YLOIi1+HY8L4
ytn7H7QiFg+QymTE1SMDfYLBmiRioKRejR4pyARL1VLxu7Cwqfr8JBC26SYV46gEOoA1+uRyPPTv
1WzgDofGNGjuNrLwEQ6VMfBimIS/kMQ/w8AnJmNnMnBJ86m/67AK7lKa5+dcYQSV7/d3aMey7NvR
OsyWT4MFJV2YHRmufelD7PUKcyjAsNP2B58KD2KrzCRfsWGWweaAfKxrUU3boCnP3B7Gx3N7rCeb
pU4uqaJIGjrcu31gFvB/dYeoaHKEbEL8W3+KugpEC88SjdMfGvOiGlzX8boWsjdcTyijNWJXAhPT
aLECLRhUG7wFDiYAOP4gjIoECMnbX1nZ+leLPJ0JH8GdBFLg2gauLFsz3HH4t4vIvyYx1GqFRr6t
W71q0fNaQTuJfBza5bZZwgOhXYqO6H/Dz2iGZkDp5iasGt34andeBJPPOdoK9CNc8jTi88qN1anI
g1QctcvJMz5a1mx3SlkQ+SwZ5bfyfxa32ijWvigLHeornUYAgifmYVeqfZGZO6oeQQWpz9c1+9f8
puGFB3BHHplCKlOsJRiXHHhC7Y0gXIVyO+qs1rKnH1cnXqSbGBW7/YXsUjkdlAwOm4ePEuSsecMl
amENw6oDgS0sdjcs8savX3mx9ncMpX71vta4bA7UqAYiznksM1NjuossJJSAo1t1a+RHoyLSr69W
lfbSHTKVVvNVxxUMcovkNuXCSj0I1gXT08nLORBlu/oiKlGyrd9oSpHK8CafcgKp0BCelvuX8KkF
DKdssD9fpeBce4Xv6CgUPoT6Il4JYRwJ/n/0sp0iRRkmBgl1w2QcaRbJPTf15ASRZt4t7sMXnQXv
4t5cWLeZG1kGqX2YDw4Ow+f8elJZ7tPvWVYnw07OZmsr2YEd105TwZ/gvfDS2/E3I+MNPdSlF1e9
UVbOHm6Sq/a6ivA5RFwm0PtPzGV8rPQShLcRzKO7M6xLdO+9lX8z/wFKVdw6D0MZxzdNtkFpThrl
/rXU9eeP7W5KnzB0+/JOyzUomzm0w06smiHiCiKitxG7s9V6hlmvqvEewxuFbixUcf+wdA4DI6Dd
Ak3Hkh5XhlSl7OJv0G18AzB/ALm9Xa9Yc9Me5QjCpnr5n9GkkzUh2mhjXFZS8cyeQwCNVudOw8Kv
mnx+umvTjcyUWnI226qjInDEOoRWLEyIRDnz8u93FpkrcFG05TWffDx08upMIBG8aWj0NerRMmtQ
gEw9c4EW1g1OXrong1+JaOZ/PYJhyNvRZTKpLaUSGK+fPPqrsIhxT/2gqLlR4FYiZuiynkI1AGd2
FHULm4PiKsre0xBnB3Ke2FBfhoZiM/Bvn4+Yojs1GAdcSWBv+iVbdX0aNLeyLOWOSpTK9cvnvKWc
0vpshj+/LL1kqDhs4sXB/WtUyKQhFj/V2S2T+izRmTVLZ+SL5e6rjuJm566ZA2G4jYvelNmzA0zz
PYdllr/JOFggROmo3OXJPmiAuIoz52DEwX8O+/i0uKgxdFN73v2B+aGvikZQ2w2px+1RZsqOTIXU
+j+7cWJmDI3Rn1ut+e2oE0GRMX+po0vt4Ej9pm5ayGBwMHwIxUc9uYBg8/hQ2x0iokExr28VdOIq
zBE7sRUbG3fL8Xo2w0GWYhMjA+C8OLINbpdWNsUiSk/pHCJbbC3QbGH8EWtkBcwJmwGJNgvZIMRG
monWrAePSlI8KA496LfqM0SDvm66XgkfSsDEDlfYkLS6I6Mn+3lTr/IaG7M+eAOYLdXEZWsivpFp
X5B8QiTt1m0GlRdMHM/UXdjspQ43+dLKW1/aNFTFA4FTYMtXCPAclCOM2vPPOP/HqA/L0RpBibcV
D0FXiT4MPjcli5rsC9YWnJ3h55oVNrqE9Wfd3K7Ey6h3h1Leci29E1TUCSwt77WpzyZ5277o2vLf
Tv8gKn3lMLBgYUcKgxwRsWR9OZrsRFO4WQGFtly/vWHsJYUsvByDBcPrpR0cyjiSh0h7fsykWb93
b3JVIpGwhf4rmZdXyik3hFGltQ4xR599S9UjIot9/y67BAsZ//xZHI4FUZmGrQY42XTJj5R0tGXT
H0JnryeEkZDq2z5ZMjKqDNb2hJQ9oZKe5QYG77OaEjmWwTqQ7l0+cixTW8Yr8PfH4l/t93Qe+gNW
qkNQL+1IkSMx1I+R3XKFnJd98yJSWCkhsKUeBGv9KCw6pSUjARmE3ZezR/ZPpndVG381M0GotY8s
iZoxteLf1RC2VqxNhIA7W3iMqTC0t1nmikcMDplQPAJDqnnBZFBSIKJViZXCUSbv3OBAgZ7ajMhn
aJkML1CLOJiSeTBwWClf0h3k3CxULC5SD+XG8wglC97VQ/gxVVye8uDMQekrmoi2YBv1b0ZKENK8
ERhpOgtx/jG2aVysjHp1REUcU3jFBILWFJEJ7TiP/7MsX1Ko3ffmXdlJXabi7HBB2lnoPDLGyGxD
7dX4iSvK9ElTSPxuMkP0iCF942S8ubu62frszwiG3sFe3qZ6IyYpPG8X71f/w4NUVgcRSBwOIYvs
qeJ/QgMPvB3QlUJNh0jLzSwtDh1aa+LuBK79FIZRTRUhIIjb6inGEzGdMOnFGx3eRv+B3dnlHEdZ
Ni0kOrVAzmT7Tj+09hyL8s5eXd7/S6Fmu2k6595ITx9jYJ+a9xdjIK8g9FE6c9PITpa1Fpp3r8pa
qA+pRQVbr9yh0cwNVgr7bDN4t3wrFfcf2f+vxelnLL7EhV7/rd4ifqvrSBNPXHxd49U3wGsY/UpP
Bs4Yo0fCpT6YlG5cY6qdSplWwOJy5Sn/85jtZQMm01ISe61VAqlkmPlN4QdxRGD7tNUyiTAKVtXc
yzK+T1wfJMn/YRCefPvdVl8S3k/spghLGETVJxVkRX91tYaWrTUseMsEnp61zQ2QP75eknobYiLh
LN3Op6a5ajiZr2/pyOEbEUimaJoGBsnttqn2bffXQz0+4kNBgWXCB/t0+mtv4ZHE8OA6dP1r8nWg
lrMPSOVBixcwv8UtVmv8ULo+qsQMyWCUw+AX7MQYEyDEYembHihflj31tWMV+yfDPgzf2ErTKeG1
3Dc/RAPX1/F3VfMI1Rb6pAhmfpg7yHVj6jvuo7sFGx16Jx/9Iu6RoEm0PAviZOZIVUauxoFKfelt
5M+OOvcNEXdxuBRsQw8tVKh5CJnrjF/IMGfU/Vu4WF4LLz2F32q/obkFzQwdzT+6bFpoG4447Lbd
ZlmlEYqxEQgc1j7zplodHKZOgKzSt2x9AA1bvMF4FX2Is7ShRgOMJ9B37zvpCoLCa761eUlHLY0F
MF3ZD+XFSnzdDap/2XmW8STVbXUm3iKbXvT5gNRdogPtwEg2s6tSD0HMivBPIJTdPAV9VhgVBctM
hLkUVzzBw4qqPWpxEJfkhdymH9mzfrSSJKMOL+7wZeJ5ZvRZzXyTOfXQP2KcvqIPuWrt9vV2Pyzv
HlYYJZ0Efqc+NrPMV+Cd842B7lAXMHCkx8j61XIIwEPiWqXChXP5iDYaYgRPdx25uVJB0f/1h6SB
A0UbQLu0K4sdBNXvaPdT4y9ud5WM5hpConn/EZfjo8Hg8pSHHwd8Qsbd8AU/Slw29CiTJ6/18b0S
NYd9UlRamEZxddaGZQkvoivrWqHJdKCy03dNv+D0F3gDxyhtaBkqQUZlbd2WABQAy/uFZU2T6vIc
ZaKkKkRRHWXQzhIq9renUSayVVxmYuqbreistdIic0Vb/G9nS4suwFjcq8eXHAUscl+OPNcU6NAD
nqkoEoizrAjoKdHI0lw9RtJh8c4jrtdKkD/CdOUliPJ0Lo6Diq85vJjxUfLp7w07w5L88rAlzH5v
zxyB5pAv6TJ7WBZci0ftcfM3EfwnEHAeglYhuvNvN+rQgjvLzY6OjUiUgBTbvKLl1RiRetIcZgHC
TpDiUdM+3AYMSFjnRDCbpOqbYqGHjJWJO7m8nQfesaqKC9aXBuXlzPZBToxC9RY4P1Th4eqs4jFt
ggKGV9kj5LrEsQaWP3ZZCqB+tI0dllw/70cmaHQrGvkUo7s9jG3dDa1Um47TCcPKMw5W9ZFh8sIl
Vam+ho+nt2nC73peeBvsh2nq1KQh1FHgr7knREerugfd4huJyce0KtapaiYURGOLtqXcICy2IJdb
tI/40P0TIJKElfTAEUU47pyoZxp+O+/gnBXwq6ie5wD3bGFADJ9lvboC/6K9XZxXNXOuxI2aSpmj
kq8iWOdu0Po0fWPlss6jTvl3A2+63cGz7iMoDvwT6ul7mb1HHFahqCcn1zrwxhFjHC4BkWvpNU+N
eDjQVYceyLWTl9/sWXKoS1vg15OIoHkybSMaQDZTAmNTgdaZGx9D24qA6JGfBxiqYxHkjo0A7Ni/
WGaHfjUO53L6bqQioqUD/xjjdoU/cLlZAccC3cRdhXM9VbJRx7ADAkEjY1m0U3wPsXTlpl2L8OES
6W+8r7OGFumCwITqC1lI1nA9rM6nmwx+nslQMqRkXtYFP8lSHkiv13h08SXQosJ3HGzqNwVL1KIu
SzKSElhVRIyeV47dENTKbRi8KhKW6tswp96xm3DcDR8NQjdwWQQrlNyjJRYLbLg5m5QKMNU9dkoD
ohtVSB16MMPNCI7bAbvThga3wb0JaiiR5F4znll2/CyXjeTvwXqQ7IF0ec+1loHpfSjsMwNm2ZoA
2swFZpfGb3UX/bqPwrXRTagYKTCnr9KgPfPmYhohk8SBpEuLc97GGrmL0bMVv4p1PThQyrln11pk
uXbRSfaR5ixb/q2wX7wv/ihrUzVsAk3EmHa5cR7uFTFLzAOGp7PAeIKx8EnWbhWC3Vz3KHrb9T1T
ZquLJj2VY1jFx7Loo7jGoYUqkkxyBAoxYDARhNgqGJnr+e3sUSc2xYml9xpXDAtceTV/Msv+lTLf
HbeVhfT5M1kfiMa+6B29kGNdk/ALQ3DHMm71QHf01h6rl7K4i3SCy5K2Xb0AQyHkGUzbqtsKzJjI
umZGASL2+ev4123hsMbX50SuW7WMsdftRpbeGgI4zZp+nMip9O6qCtPp39aCA+SZLDy1ffCtczUs
pVMilZibxoZvsZMSdSGMBCl7RQNjiL8iE667H8bTAdcia+JEu8ppfYjlUXuun8x28YfAj4t8h6iH
gzXSpDTLWG5gSy7mhvURlBsTqvX5ZPurL/dTvo01V7kBqPqvQzYMNC+VqJ3ryisp27H4bFeuSVIC
yH2sO2quWr3leBHLtNmJSuq6tUUE87Uh2CT2rKMfDfFRKIy4DE9lFJFMwNK0w0dRMl9xf8ahUHZE
YqwSPMVNMPgRUo35j5DeSUJ9ccCyNmCngzvuTWn7QgYDKAuFQJuZWMP2P0L4XlChJ6JaFeuG1bzb
0kyh96W4ehwcMOS7tGDZAdy/oRxzMFudpk/ap9r0vWdqP3nvuv8RsvdbIkO+slC3Ts55Q8mneCvN
fJ/qgAmaKGCCWUasWWaylyi+I0/q/GcyP7LNdMSOlLeNf5Zcr+W0Qi/y6V4kpWazovgCnaNvE9Nm
n4L68fhMJGidPIEVEl+lMvp84V7PGF4PN2tUgyaDQqIdMVonfdcA/VKh1GbZuKJEXe8Y5xSEiVUT
GiuWy8tzyKB+R8Utp9bggh7vKTe9VbVIDJArrS4B65to3RG8Yuq9UlWJYQI9BzvpkM65COa+LoIx
6OWRCFyRMbEWj6jNz7TRFD1ZmuulNqXR9JhXnkjpUzsFZ8f3xQetERGn2fVKBeDo2o1cB4jz5/jX
s5E40mY7viL+CWmxPWctvVayOMg6ZTqFrXo+1x9obfEoelrRoIECsEZQYOUNOx0gzWNJA0sKgdJ7
pl38YZqbX7hIaQS/ZbDZqOYWQiFePGX/nkMzB7UL55h0pcoLDm6ppcGVr3HgNh1GrPG8k4ZZdIq+
84TlDqixJa4/AUHS198EU+Y94hcPobJDvALEHfGbEOLQDQ3RqJxlL1710yvJwDP/vVJs0ODaZhyR
R6NOzpryF9cILKEP5WRubbeRxY5/n3zIBWbT/812VDCbVxXHxCRRk9AnEQbrU/8vQJlwDR6M5N/w
aILReMm0fLiLvRWD+1Wb6Y8nelGBqHP7t4m4nTR8eRbW40wZghwSTpavn7PdZHsqEp9m6DICYbOM
M8FqicMN0ePYkgs8EfK5eKsPkxzAilZISk+lnBJhQGPdL56KGOWx8uN5e+v3WltGcB3AWtIVa8Yo
+zbPjZL2CaxI/FTyGqt1dRdOVUMj6dWuWkVSxsveu0XE6AE0CrX/+s8gj2WMmeY5pWrOnWXUa+Yd
xXLUpx1wwYoOcrWV/jAjwdX9kbVfeIAwRIoXulLBaqjkZdiXDSNS7CzAhB4VEY+QS97PqXT8RwLU
zxDtMhbESHEiel4ciyHZmA0qMqKcLQkuizzpwFiad0DSoNzrc1hK8bz8UWeOxRsu+EuXs8KQ7lkm
OrPrKWnni3TjuCmIncO2OnUDrSO2vySKo5GW/mvGMXwQUqysoW1gTwLCJsRgl72rI9FeqdvVQ+Ax
5O5dXJZBFNfMpsH9pd6PntApzdo01U+t+xOs8S8GMXIBHkSYIcGspMvcctMNWhbhRMKEuMCI5EFK
LeAEFE0RxvzATRC5VJUfWI0d1w3W6HlDupqwyTjuIXGGL2vDI46NzGBahq91aBxLinMAYSEc4kwg
AYG7rpc15aBuutM7GjK4a2XC05ni56n20oAP6mADwf0UUBuJIB18nzGWMN71cTyt5wNVuTStUFIp
UcIXB2CBcECF39uyNpIsnYXGCFVn7Ch/u+//AxHkpinsI9yLB7h5KSQMqyk0K3j+gmlUaylG+YiK
4HntyPQt3yl5vbl/yu2XGyJ9K+qPe4weoSEgj5TUVODak5ZbWvlU7tM2ug4kBryLIDdcUgcIWP2g
BVcKh2EvBGwFmOeYso5zjKaUruz1Lq4yywhWkacm0yUtAkLlFSqOLXhbtK4lPM9Kq5VDhIHCUgqr
EM8G5Re/eK5hc5RCezOjBie61ByeApvfSBWJ9+8ZVQ4aq296AeFzf8hlrsD7V2oDMvHCy374DPpq
NMa6HuSQJBofEKik+dq7y8QXcpczjdrLpxZM+piH1AQ6FTdLQpeeSi+iyKbrB48LAQU/F03dvrPd
1FEdvqrCw8m+4hzZuYT5heNcAq5JwYSahP5Ru4YvTjepRD8vC+zfvxR3vLwacgFCAqgEJcMDv/9n
9qy9pi/qSJkwj5/Fn7v1r8UxwU+mBNkjh1I4wiOkiHfCywhS8EyWxRalrkS9MSjS8yPz5ZGXgqCG
n6iAW6LPQGPV5v8RbGuATHP/uq+Kjk8nsskoTU8LdpC33NuxMLopkIwWlbQ0M4zIXUoBiP+WH98s
uN83kNjUAutmmgv0A2Vam/mYPnCsIJVsGJ9kDJX4m0qGga1rS5naXGcDlbpEM5SwdKEqpjgkrIsI
bQdrAMunANWKzx8egxDHXpZANEOuUBivnsBjqjcO7XgUCVzeQoUNNgOQnaIE0CRIB0ngUR416w81
jWPVSwACdQVg6s6xyUW7P5dwCFcfl3ydgM2Ncgz/Me8uNzcvatABJDTKvvKoqCw7FtNclUOEOEl1
L4hu3GFKHXfL9J6z1p1W8GNzEiYjbbbVODN21WXmSGLjx4u5+9gJmH3NunRqWrRQluetM07r8hm8
9KI4lp5pvQ0HR+m55lxkBC8HGhcCoOZKhPd/eptoIbn8zvwdBjJ2kLXUntVHjqr2PrjsDTOCYBUF
1deorZGT3UYg1WXQQmycfOSU5dQTlTRZOJX9rd8AYdugfiF1Ke99Xuki+3AWQRTs37TspxyvZA4g
x41gqTsgT+/RgqQqpqlwXMTR5+tI/6Xl6lHYJb0vjW61wCeNIGfzwqel1c8flRXrGWNB7+v6gtnR
AH7YJJGCzDKZ3IWg4fu/C6Hzz2jwwTh3DPTWfOqb9r7rmeua1a7E3GUI255jOcj4WfqRx89MZapL
jLqoTuvvx6JTYK2Mtwa3Uf+cjI0qxQL2nLQPoVzjnkbT/TUnxDgJ2SPDrS8RvYedQ2zlxnj6DKNN
Ws9DaxZyaVnc4QBT0PqS65nNJUhayOb2gW/ZYYamOHQP/JsTSmITX2U49r+tA+VfwO8W0VN3T3By
/MMA1pyzlXV7WaBM+s+HGqfU8YeyWo5AlWhTGEmj8IHUg/NCA9NSYJVpWtkueAuQNjMFqfqPfxjo
87RqGYj+l4Y3kM3Z0wzlXrnGMyajaRWFGU0w9Ew/i1lFOUDbgFeZ+t1z6dV4T5yM7ux0fe4TpJ7z
WKd/CCWUU0/UPucck1ZNniWZJlH0Q4NOogzjYVTuoXxZEP/nol4OR2hNKBLsM9oq0yF3GF+LkbDR
KagfpM6s1nZZsUfCg6+ClKOXlDqLvpM6hYW/mydRrkEyrjyxv2tyAz+Mp3tBb/umBppsp5qx/vrg
aB2p+oODxhBctTO6FZ9gJYn1tP6CjwoHufu/HB4+9AbCLLt/geAcqwOJrJClqyT4HctyEzn3v5YZ
zXZmgul4cO9LrUIrodCzN5C0rl6L/dh+aAeVJBs1hHy9n+mNuaoFtkBZ1Vc15sKGgkcCw/dvnIrm
OPfvNwGX9d+dKnlsMnyPqst1+dxe/GiFftP4FpUwyrASAjk2+hfKwPr8ymWyfWl3XEqosMKhhxOy
FhGPiOGJgmNHG046T8QtTnV/tUldB5bgGFmxt5UWBMGrC2CMm5PaCWPYUwyxhjy/ipcOBEclvuOS
X/tUkXvuGMJHe7QNwzDYvfAIoa/hLFDI0AL1LumIwqYipTpHV/kVUVCldQg/IyN3ZBtk9yegkP//
mTZxWXDPvopIM6NSC+/6k8T9nbEelZVH63KLmfUi7DTFuBFl6ilN/nju3h+11QwT+bxgd0oonFQt
dw9o5DsF9XXLcny2UW3lpPZqUAg6pfNU3HIsqdicg8u1ps06Yr3204bq/RAlauh50c1xS1wiO0zZ
o+WcScFWQzxv3LpGO6XTMmhMNqZq1b+VpzyQGsp2yq9myIBR3y84Yik9gvJ+Vf6tU6AVbrj3KiRQ
H6u9NE39MLWH74YBspmFQnFSXUT7mUbxLxlXTm9nxtpo+HauyAyzWdsQ+SpLHkio/Uq4Cy1ueh8G
lFHbM0EdAuVwuR6dlQ0Rl7KAlbHRWcPZuDfQH9RB6nRcMf0uK1eT1lXt2dorsvup3SyoGG0ZBa2o
pYpReyGvVqF1wpVTLnyDT2+0no/8XlJYX6taDoexavGx09xBedkkS6GxH0suoSV4q3YNIOM5NyH5
hhAPEM6sJ9tseH7aQueTEFm2ZkDBKjnaGHSaHe8QHBP0sN/jsknx8WYV8sgrOywtYhTeOIpR6bjq
4I6A8FUBEe7nmwVXGT3xb7Stoi7Zojc3emZlc3Ld+UnzLmCk6DJFTy9xo9h4gmQIa4x5938XpR1d
rlk2qAYcSnh0NhogMANrBb5aAfOIPyL4QDMAYwOYfmoJXmoAu40cXqVhU1Dv8jcvUI3ilf4Nwk0P
G7gOpb8MxsBmTzroPMcKx2OiOIIgi0BF9tee6Ezqfj1hs5V2S4Pqe2Mt0s14AodBBu7RTqaqNik6
xTF/S0cUmVYstiioZHhmK2P0S8OB8Gc/5VfDKnJQJ42b6/RTl4PbNFGmUh+X8wrG3FJvQqXP1oVo
Iv5HpXZp/lBoi5IFcqT5eBIAlCSkBwe6kyJp2RGBd4vsj72AQzFmVZV5L3gRXXVxkCNsLxJhlfNG
jk0Vyu4lWeAg49++QoeCqa3MtSwdHiHgB7mgyLc0277hY8ked2ZXgx2f/pv4yOSrxQZajMSA5Iky
R8am+AfoJ+EgN8R8qVFCbPBJfVW3lHmBKroZlFjOO7SdQCa1GbDsFD/LJkMElj+YlWXEpFbcT4IK
thgtcbieVWeajtknPXpQN78zMrhznBw62QAvkGmUzUrlixJVms7cbocN4PMxTTGWZFRAawtHc/S0
TKj5Gsq3MDl27HdFYC7v11Uc7L+2XH8CNE0PcNgBuW0aMRXFvMfbfTOs+xTcLG24AMiNMpWbBDuO
QHeY02732Eix6Z5oIIkdZ/QXZTZKL3uefn+m+lfhnFEEBN42gW6pou9RvKovPOuQxRsxRfe65gAp
eqrdnHQH2665ZcxSXtjNP0w44JAbLipxKEVJEw+9M6NUUUbWuN4w5VNXx7B0yLCIU3A2utn53YME
qKlRvJMQ3Y+/lSE6sscDrWvoDubtVadmxVSL6UyKHds3f7b2jIdn9g7sZP1PtaQIuPx1Yi7DdkQu
KJlDeMN4AJHjRT35IHy0lDhx7XtWtCDABa9XU/yhS1kEzI4xb/gDpat90Iam3FkNMalx9c/1FQqa
VJQiNf8SZo7V8BO9Q/8J3mf+YcYh3gJsC2MXDMXlAxW3m837dr4JLv6YEoy5ajJaq1/hqUes775+
FJb1e9QKiWgzebFrWXIwfGNe6L4ZMT1PlI8m6HOvKqOTUOjzkK2vPfMK2ewZ+sVvMX/jJjCgRjah
LL8tqjsOvzY4qI+y/DmBvE+dYpREaQu1eIIKog5VjLoN9ihfcta59hAIMFCpHn51maW6rOQMlTc7
/9K1Hl4cVfzABugaXhNB3wOFDu1qu8MoCixJgW74JI+zoMx6pr9Qo2uGlWHQTfmZAofcM+f9iK95
+j5QX2JEbMyr4nDaXvta6X3rAC6UH1Tn18Dnjtu04q1KqtORQ8r7IxROnIx7ipC0OB/2G9NAzWI8
xb2g5bGBZtINeeRrgbAAvUakFGzKQgzPa/ETj1wN/WvLabcXjeeOhuKQFKXD72pB6R1jpzvHlJVl
Rvm3Ac5mix4O9sbebfVuqXobgX4j/NJJyzdJf2ss04zj/CExnNHBoTLiPQdHAdngYU17kOUbTpOa
2x2g7v7sBZBYpYgduwsZRhx5J9QES9wpWGEVT4mHUk03LqDQGvJOIKeKN0pI3oKmTs+6DypMrdg/
KyxZN1GaTABplxuVU0pZPs0jB3V7BwSLDU5dOlQgQ2j4IQdgUcfoefvDeBv+AQ/EhIA7p5v9C7/e
nKnTuo9fdchdy+A1znMQbTSB/y5G7tzYBY/LfSWAwAdTlVZ3BehILoJLAJausGBg6Oto4k5CXxdi
0GGZw+Ffp08WwCle6T4R1SwjRazYae89KkRmtEwQBpCiOU3rjjMWH0IntVE3UqFSOaSN4d6I0ahE
Kb8neoIPGnr1Ao3BIkLHgfpvgALQ5JRz8YhaCdN2ZNPR08fvDbrlBiJj823d6CgSpZUQwIq9lZ+3
RnHm20l3kCOzIoG7IV3i8gzjxtCZmzcpKEMuVa2EFfdpBHyf219JGy3fNY6PT1tPmXPyz2WtkQ5l
FEkcU56HFi6qeblJltXDdXlCkkZo/YJ9DeVYUfGFH7yvSRGk3JgGPLCbX8WMZY4+jwEbaYHlDbcQ
3+R9bAw3PWtbxAgJsKruea8lAIWcGjOISp91nxrt2dM2wwFzo/9m+xssrB0x95EgNGn0brS9AB/Z
f6iuTI/WHi2T5SERVdATGxTh85P6zi2ry2qzKHlYA2cRYe9lQt00ctt7ZlW6g8zLsXuglrVBRHG9
+zuHziaaFnD4vu8KWcZdHX5aegWPhR6v1TOQr1DOrWjd0Y/bVQfEN/GcsnwWoHiO5l4HE28f56Rd
8adKkm6Et6jveolitTBTRwDxL4jVyUvyDRw/+E5ELKHh+V3kE2o+3tJQVmobhknNqLxSb+EXRvhK
NL9RBY+4PUr9nUBZ55lwDNyR4bYYDCdpgLp276nW9J0LQkulbzNX1qAoJZz8Qx7/qGnlF2gslekx
oEuaeQUrcy2Ks9pJwtnKTPClppS9PAa6r4kqwgQxUJUwaFpdNgFy0Q6qC2TTeMML1hNI10XhCHnQ
xTDZ9u1J4OgUJh96wEVoCoKsTE0RMVDNVdLJrCooPqxSUM2BMOtaiY/eEyBxQaNzQis3QvzZE6/6
Ajoc3eoYvbJRKPihzKDQpxCAGmluh5Aq94nFIQt71MKeHMuFzA3ehUS701gpiXnOYGSSIYxYueCS
GKm15xwKiGaI7pqV+HiOCvulF0xqTwkbnBIA9iW8kLRcVBOv+zXMo0S+A8b3e91px9Wz8UMI0Iss
emwl+ihbjCtqenwj2yRYMqOXJGjGXForyScyHJWJLZKYmPpYD7gMYe9qTVn96nXRjKShAna8raqt
O84TVO4rWpHI7gXdLmB/TOWcVAxra6SCHeiMKl/bPIh9+77dghV3MGhRws04/8QZl+tP2Yc1ft7d
S6zRmWwR/ziAb/A817wZzx0ikahGWmvjJVuXPczFRLoHAtfxXhWhBm2ev3LT/879gzUf7ybWnbny
0wKlDP+DwWNTcEVErxfNxJ0E9Qyl6i59M6PD6bMlf345VC7nDs0dXcEi4YUXNirdwB9PL7iO/EEW
bBPyyofXb5URJDHHsiG9fuJuwRkbXkfhe5Gtw+2hLSQr9cP7HhqK8nmGVxflBrDSABXTSnlex2Ep
DLA+bvxM6my/+Rr4hGs9ybdzHzL789U1q2UbBjB/RnE7kQk2zDBA0EaF4pAzrRMr/R1BRQ9iuNzj
X+GdFLuRr3qLPEC+HQKb5fODNaWLIczfCSjknA/qmqwLkhuYRjUSNGfn593jCeMwpxfSRGQsmHin
Sbk9ov2VvijYrJNb90sIGyOtuvX2VYZtrLwRzlKf2Pwy9EPUEOOf6qZeLnHTvQHAg8oM7uN4OU30
i43cjlF9njj3ngHcffC+DMISIwSNGdEArNvrX6kDNNAkRDUoho4+k8X7ffykgnswErxjWNnfGmW4
82ZdRJutwy2kT12MxtH5dv4ko1iVW9X6vfuGjSRYqV9v3HQyDJEWNdl1dWWoT2r9g55eT8/Xil61
5x8suF8kgu1FmUp6xq9hV8bF0I54q/NIJcVCj7tFZxlAflruI7caTea7Gzes0x5NVgUHEv0DFrCG
D8JvU2xkmxdpL69tODFNq05p+TXJ+OPABWpdpHQMkHQtIjoDreVYZcedTUkVKImX6cF7VqxUiaHD
SWzNh49ecd43vsnUI7plYx5hZcOaSpdmLgUeCf/EAgKgZdwyv6+igCBQsyjOaKrnMsA2gvf7FUEF
XBmi+Akbtesy9GUhV5epFt4Wb/aBi/QEcenO1h60TgvyKM1EjEmHvxx22esysk155dnFpNhARMEU
zsojClxkmpFPq4nlH9POJExcPHsvMGjy6V3ES9tT9WkUVmFdANFRz/DJzpyijR5ff4nUVIh9d+ga
WwG17hcoYSvOcypnGIdLGvzhdP1NImH+Qp5jGS7qI8kX6Rxwsf18Y+9IEmeAMUiODeP8yPz5RA/a
ewkyXkHdTlpcojcC4YjFLs08YxQF6HRx6G/qnffKDjMnO4jsgwvDTze9lQevCDu44XcoXG0nmFeO
Jmb1DUYy1+jpYJ+6MWB4Km5oLbYz/wXlGAdUqobKqZrCHWtR/JfB4sU2fQacZze/Fv++N3aq77GG
xn8MBQt9ppGEQpowCOZ0a60SYqpUjwqdd561/4GDLhVLePvX7I4UpjvkAekVZQXx60HOyrKmFbzQ
QV4Vp29dAu4d+NGXBwmj7NPjssKPnemmhYss29hh4+NsVpvlO5Sbxw8B1Ns2MSFPhgIrBKkRofXq
e+h2nfbR2X5cuaMMKS2w5rl6xPB4NrEyaPPJC84M1VKcbYvp3orSjkE+ZY8E/h7I3nCue6voxFOG
6mY0DBTwGfX+Yx77HKoPDK3Dlw5g5YoND2ExRpt0mcnRqhca0Gx6Qvqexv9d08+/zDMv6VGL3URA
XwukMjpzI5xr79vINMtzfWEYFo21wsXaaEl5eDNm39GEu5YJCyjZL2E6OO9LOzQAKbY03xJ6oJnD
vvY/biU/vau76ITtKarXJi+DxKqZ8j3VOQ497OvJye6Yr65DwOKc0idZEA3NJioyvPUOJ4Z6SsOk
NufD8rwye5ZujGljpRhWLyqVX29m3jzQvnXSShuS75bqMvfSE9wTj8lYyIcOXT84p9LejbDjbBIU
lpt0e0Nc80TF+wsRzk0WtW2y9rz2Y+d1Uv6E+H5V7PDxP/M4ahkBYqWS55dHD4GQCtvaMu5/ufCR
vjzBnuOgZQpmkPhZFpRcvfJKGB+V12EvSyo5GnA4DqaRyFeo7uQu3PxDf6gcjDPXTKCoCBcbgaCZ
nh0m6TxYXCMJwN+PzOPw6FZoi9AWZEQlJ9UbSkHHQNIG+uAuf4rrNPfhGLzcY+yHIUG82r5IbCgF
7e6mOAy7FRn4olOfivR06rEo88Og8H+/ly9kyJAlJCul85eAjc+bTGdrRMPgV0qcavkOpAwzSJ7+
XS8y5E79qplF2Q6mS9T6TdNtm1g6PXbEI5Kfv9QJfpv97MytakBtGCjQIlFgPSRnH/UtwU8mX6sO
XYbkBj/spSwaSgF4sUKeku5CdAUN3M86Q0/mSW7kgAJTDBybNzSzyApRleWnRka/etKeBFJJryhB
Y+skmaR2drxTQ1jCIkYn9rf07W0OMujCWa44PQG6k19Wc/a4mEM5/uSLOOQLvuKU8XYINepVrg8S
4a2dC3eK3ckyWZi5ICs8tqs42v2MXuY86hvGODNPZQY4dTHDWFxoueMEkhxhAFT8RpKJMngVjXbU
ADgiVU82B+zGUCEsA6BRw4jfAzLVNBBYM2LVySqRi68CbLQPcBeoFMuIDTymklup+jJtG61AL07S
glWMzo16fr932qHcJm4nVp8R2w5DDre+7mLNq6kiXMk82g5SqI04EsN+HgJuVLi8cEL8m+4HoiOc
HRiOb1KsKJ+QdklUbOihkB5R9AHa34xUemsDTM8NrwZExrHD5r6UbDJC6B8umNI0M81StNkqlwSK
nZkAQn30CqyQb+jfbdqx8IOL3tzaqLkrS9qyY47q2J2ffz+Xca5WoffB6TBaLTRrueie83fGMdya
XPqZignIX62+AAJO/D/fWbPyqi8YMqq9p3obWvC7HK3PCQXkC6joyYwbKxjiJw75/fY2sqzmX0Tf
8Imdl4yIB5uDuI/RK0kNCc2oe8yVm4m/BPfsE0i5cFCFVpF0YYEp/IhjPCvg5uYYQnhKVWk8j7mo
b0TY/4sAQcSESkYIJWjBvBVe9aHEaUU2xkjg6N8QCH+fEK3fUjEyC/Fwa+kRK6fSa9N6CyNvYS8r
CRVg6TKjEowF/qRzDA0Ca7enQU9kAGNLvLXBpspA9m1l+ZOZz0xOIzzqcPXWS8xgcxVsvL1MJJM3
ZaIbQrO+PaMilEtufvWJq1HWqqQwbik1mYgv+vrlB586j8qkYC7xTOGVRvaF3wQCUxQSazUDrMPp
nBiwJmPiJ0jt2NrZ3ZGm8VVdtcDap94dh4OxkVdZobtkKk0evPqCSRptUfHfMSGX/ExNkMH7WFJ7
4nkH9Du0C7xV9qcl7apVDajFKdMVKZOo77Tw8HWfJHSCNb99GKLqwZZ6eIrHuF2ewVXB9wMT9Egt
Yi1g8V6R+VdbXZPmWDrjK4sw+7tLM8m0ltlSluHkhDLMwIQbew5GgnT3vMlY1UQH9n+Npdq3wnNg
bo8toPLBrZdG3QutYXXRyGZGv6dpwBUoKF0eZM7OXw7/aFUQcHOEQC9si2niKNIMr7iAJNiYbkzj
xOLAguZ7boTwOmxsixs+p0HHBp/L9TyhKEitH0s/N6wB3NvlJylyx2oQK7/vnzBeLZhgE5CyjexB
xFkXHoWwAgwJTB/mLyndPeIGRqlgyrtX1wT8ZxPqv9fsqbum9R2oqcALz04MgxYlkqp/bMIKvehS
hKExxH17x8Ibe1dhUnY3trYqraKnk75Uwnlwqcuuv02qcC8aquvXKEhPN0IIiojauW5Z3Zmh41sv
UHEjgu//4aScQ49Jt9Ja+3TPUt/BWFK7ogAVWXN64NQpAZrz6YXFGFpd/m/gYjtJYug2qtiDT/Fx
Z5tfsM620AO4l08JDOZpNXbFLG8/dwNvg67ZCCGf10bpLoQNUl9lPLarR42EE03pesyZEKQz5ci/
gzDVsfxIbvYaL7VQ3U7f4iP8Q4MIPxsA9a3CiGh4SMUr4PVHo73RIdMxYIvCKXAIwn8mUmS91E7B
h1kK9rhEL07PNN5VKnQsk4CueNZhJ4jbOcgJ3npCqwueX3r7y+nEIa8eXaeXEaqfyUjt9sc629A9
hTknMjCskmOTzNU+AKkGRRHesNMcZtVHcX3beG71JIKCtbYSvZmrcLrl7uozU7t5sA9HTL8Ppjc2
yqBRwWtWjG6ijAdiL2OhIZ5N5v3k4GCZBXzxcXqpTg/9/fQOhz2YC+XdBOOg8p7cC1ojbS6TYin5
4rJPWcfahNPDDBxUV+1+X2+IAIgpgAaUotYuz1Sqvn8BncrkF5asGjgeaguhJSeY4TeOV+AOWTzI
RwrCJB4E6QCRBp2Qs3xexBZcebG9wlkG0DDeKVHkgtbfbWW9AURmZ+x7SPXHO0NE8N/FBWu4xbrE
I1/tEbS9iur0DTP77OjY6bOpz2P9Ct8ZNgF5HUyOBCXl6qIttlKHS0GhX8dbWaRWazVVoCZxBwNC
zYo0HI0Rne7Io16rjv5Aozyv82pP7OOH38JWvjL0ldU/vNkaQHhxHyCWz1HCN7MJh0844iBIpvHO
ZtH5FewI5RT1mMrpJoXAzlCT1t6+T0tZW/gL5rEyMWGc6Cyr1zzaRAMTu3ApCYuNDo65F5eo23BA
ry/TY1gh1MHI7A89p7UApep7ma6/F+V1lPZwsH+dj7+0Hrb8e/MVgt76cCOY21RVMIBCYCO3njif
CHOJ3o62sXwylpFJhbxYC5/CWnG0Tw1TS+E1ZeebVJHS2ycQWmLiyXagcsjVsP/Mc5ZJpMxh18np
F9pvaLq8LOEtCu6Jl3rMCsFOA9mfWIBariMHI+95/KxxLZeOdE+qC6YzmTCm+M8GXV0dDSih2Bkf
20P8bUjUiXyJSywauN5t/qJ/Tf38NtsYG6Snwd6fL0xdTeYRnpS83oXwi4o5LzpbdJ+b2ObK9g3+
fWTAXOB9an9znvSfOkmrWRQIhGGkKhQNvuQZIG2HwyTsgZa4EJdZbD6ZUiooXm0ozduAYjgG2DPd
0kalIt70csohOneRj2yFiadn2C6QfY9yQDDB5ntG/iXtV/Cb4/T12wAaSmS7VTGnukOIKr7WZiiY
83tD8dI+eS+oTXRuBdH7nYSXHuwGnYok484tX+3RcddT72c3TXZ4jgbGy12ZKQNHiVpeXASAYlv8
L30FR7Ej9LEOkwIdrCHKYUtmOxtpUZcRXVjn9mnjdM6ORNha+9pMt4ZO1kdtGeYDChtohrAAcxaJ
FlLs6sI/p3VlbWdxzfqL4UoFtYnYnoVc0PvzPwjXFkC3UKEvkBLq7JZsIYNxGr9WCXAh6Enj7sMi
GX6aMiPY/OEFw4Ny5SDPTFgzyecHyIW7pCPBE2CdoVXH0lZm14oFRVbH+jySRjZAzhnJr1Ag59JM
mgsjBrvGCXJviLZg1CRdM5sgHESH/ZrM6Bw0RbaNSdGtFq2I1v6Y9yPafqq9uCiFSZ5WbEZPrAB7
HylvgFVmI6xR2LRaiFJm1PLx+83mr7mGt7d5DXB9dCPS2an6slkpzt5ZmULtMKxDairUfaKeJGt9
FnoOGWtAF9wREYyqyhoW1JsxziIJnaoUic8v4i/mm8/4H5jlqtYZn1Ph0NDBjv09CSBld5/aNQdG
9VrGoQFtwTqeamX8zxtrT0B+V+2OqlIVbMVn5odmrpimDhrxuOr/0rjUG2t9nBm7+3N9ZP+rk5Qa
RUMBujyNeOza5Prk0g2SFYytWjZFt0qgsN3mUvhhuTfVGvfIknJDrs1yXlrVMjoezoVLbjHZbNCS
LBzyXogWQpaMrfUG4GrJ434IXi2CXUJmvGI7ZgRRkDp+YoBLCQ30RlLz4DTByYb9gBCSrlKLnAbE
9sUa3f2wfN5PqdirurL9+RL3hFDOfoqTmyLCTQnzVtsKOraSVcdNFq7WdsDcskz5uloW60AQT3Ot
4h6yuvMt0AjlvkW3yXh5omPl0QQ305IG8bx+aUT5eUQEvqL+VeDSdH/xxdCj/FaSupLBqzNQFfNZ
+exra9hhiE6Clbs44EuW5QLrs2lGIsEQ3AsG98AFGnftTSoxK6IUDQ2vMCB1lEY6YRvfFx2AlLs/
EsweAjHON35PypTNZeryLFXZVGJU2+kUGVQNX3FFZgg6hSfvWxIc+14CkwqX4zXMr5rMoUeea7ft
pOvvoo6tX0EycxkiCtAtXAJr8U3/c4Ox7XgXgXdavgya7JjlUUX1UaWYMHgqqq59v02jMeYreCYc
mt85bX3xvmHdTpUmRtIRK/SA+kwsiLLTCORMLLUH06IJ6SEdgks10lyEuwjnGKC717pinr4/56Dp
y49GQRTfyNTHfJb1+tZVKPJ2hzxbfRmg4E415eCPW5uz0dQQ4jPC1HpNvI7wAL4EFevo3VgjFZr3
iv8Og+UJV9/bZZHBu7TTxEMHR1Zn/ltqD0AF887DZef12URXaMZ5dXfv4RQqP+QJdCrLI7ZBcFdP
J2sswxjuMvVfMWa/89Zwb7cpKwGKrYCUgaicBwioXpWS97rg//DsLDkQx+hanWJHiTHU5YZwqO1/
5j20IXOf4jeaGLRYJsvTDLM9KBLwFA7nUtkGNkRLWZmAZbE36MFGtlrTOgJZS98hNxb7gk0vM562
QSzp6NFxuH7TpXEQ+OF/g9yQzyukW1Hop2JTdpkVyDKFncU1YnUPvxdabekBivUHSYVfjDMqyoD7
WvbBrKaPBl9Md3jSPZyt1abrvspVLit/IgXSBdd6mc26qiZQ6z0DMc+YXS/KjWZ1m2VvseqKTzDK
5A+JQg8W9p1+vYcrhcJH+WP1n6UH0ErXDVQqmyrywRhbXFJZw66WhvWYEZMt2c7nKNvsyd1uWPhi
yorCiHs3hjbXc/I+7ZGqmQmVN1Lh6AbZ9kicB0E3ye+DXXKrYML7pcnWdOFoYZSwfuXnWN34tEZQ
Iq1GCG62MB4DZR2an1CdwVYVA+XVJVRRHPquFC2EfSRoWBKOMCgeUvhHV6ADV2Qdhq94VUtkfnBE
YcQ9llFsByAegoMgYPFGX59qx8oM43ufzBlXy5s93k58smb2NaGEq3BPa4/GX5pZqFbugXl6j/29
NK5LOd+oMxXUTLpPipKWD+wC7rDJNMhgJL03NGfWlyFod0jLjVZkMg8AbKEzyRlVMD3Ov8bR6JyE
IQ3Og2qS3A2HXH9tZqqB+HxnsXqE4lXcs0EUsoJV+0MNRCVB8piqvQwnyKCMsfK7GcGIbs3NS8qo
2o1SD6d7/6oVIgJESe7s2HamMvf3HvjhYdvQcgZdikFPgZaiUfyPWn7dGgTMGgrLJRuXP819BrZF
Bv2+vlWGtR7mX6essRj0YtwUaM9huabeqewmPRsaFMaKWtHhZg9ETtBWDFZBbRJHNi93gqnjzIGR
eA+hXDPyoW/Xv+oij8jI9kkhAZ2t/7waFk8TfaavOrCZD4N4/icc07jD+M7yacvxeKZn4tDAqoJu
tO7LFePprXZhfwUqbCOz46D60VL9s0zQpvQF2DsUhQDEoK71mNFtcBW3DoQnAtfLqqIn41xckFn8
4lLY3g9ILO75IaEQKUzTnayeKLADlyV193/BR8IFpMXYEJ6BjzhcQ7vIYmedEGI3w9bBkOqlHjHg
yKj+rQaTWBIwdn4LOZyUd9kKqS1fJew24n/8QVr/nhcjWpZFUnEQbXPPvjB+qo1P0rAew3KYIi60
dUeq2hriGM3J5c9eSuDa1TWRZltoaeXyLsHQtgIOb8mREjdTTCIjxLfnSc6Dm6p8snIkax/FnA6I
cVS2XDdBt24/DgnV16mCTXONBr8mNka0rBuvlgD0V+TN8TWK+6Ab77njlpcb03eHyp8wwZeDErXP
Q4LAAOxaaqaGAGos0m2yQ22nNRfTdgm/sH6ASKORsC93UktuVsur4mUvDPclem6Ll4f9+7dk3M42
SzgerGoqWY/zmnVNq9ss1smfNMXuJ/FG6iy8vn5L2e29SOV4TLkPag0vhWe32ftBfqWj6Uvogbi3
/Y9QYZAwFHgRc2iBKYNTNzoVMytJcoHNpeaWX9tFiSNP6sywet/4wxbP6M7vTIBJTyCXzuYnHTg9
lGa2Yg5hzs2FJo2SrdED4DaYBsLeTKqe6+qodW9pcyBaPDuhIQyM2klxZce5Ewwt3uzJm4D2OY2J
ccN3pYysc7pUbge6E0ce87WIwxNeYL1fTS+IttTqN1r8c2HVeboRKyk3S07cXIH6VdA1biu3P9Mg
QtsvshidK+xtiQfwzuV0HWkXjbiHHOMJERnXBXAcgx3/6ngy/3ltCadRnm1nDzrM7EhHW6ELxE7b
9kTsKZ/3y+2Bg0BHGFEm9xKHDRavF+vjaJ/PZDEQI9tdRqjpaewO0FzUXkvR3CaVaLEGvvhfoi8z
PJX5UVVn2eipWZKe41QrATID+homQDRDEqfa3CC1xfGw6sOiCDJJ40541o8bpJBLBT/MaiioCQJT
uNv6E/1S5kDLCm+nODW8KEPtA9PWj1mZuv2CuXEzikxx/RjvVUy1Jrz+adiNiGwL7xGQsQ1gpjan
mzrXDLTT0VLOOQYAXpG6I8g4URA6ojZ7k1OR9sWoQLJTp9rbZOcPzafSPS/eeihiPc0M5w9fA3vV
cky0bJcUzWEPcXKekvgdovN5O9D3+7bSZ6dbgJ4ALoeIVUHSA6NAchzxq5v04AfeU2Nuld21Y9hx
Xt5ld7bbAaXFI30Zjglmo7KdG01xxNLdSjnFO+kBEwA46yM81RAIVOi2t5WrwxIrjdns7gK1NXMw
B/KEZnly3twFTzT8Fu4Jtqls4dz+zqo1AL/YP297Kx75Jbqi7GHhczy/oqAPlvuVAsL7cAEMCVMS
Vg73IDCcmsmlFXA+bblAjI0RR5YjlQ5fCJbZuHMxBEw9UduxKIQxem+d7sF92Sy9C4v9CTs6L5WI
WiToTsngZ9O1XokVDNPHEfCXvu0xtHNmicCS9+aGiX60VNsbbtgGgWKB3WIdXApfk6Q1fof8x8fM
9+hed3smaKQjB34g6nhzvA5/iKJGho2yBlTYgAyyxcUM69Cyl/cC4qDXzgUsbGrHXLl3Kjcg0+5q
vmladY7o730gC55tmOZ9VvIQLPXT8ttiwL57/1FrF1Hbea/L0d68DmYxq/KK0FC39yNSxG0joRBo
zDxzk2onA3lX4+7oSdYNznLcw+MvBEGr3ikIHfZRSUWI9Pt0EnG6cPYquMfdp4wkl3DvbVOu1Gm2
y0llujDtUejeQ0oyB0XiNO6Y/jqdev78aSyfgsarSKHbvmn7dGfK/PFhIl+djpAqrOkJgKTT2UfQ
XEDBUS0RqcHoac2lAyEbyGAQFCd5EgsZhiGVWIQ7Ku64gUsnDb1/7+VCBECY3qN/+a3b1QXD8TRn
YXaV9q3OoR2OcZZ1xUgUv4GsdqXlLAxhUxcVuTTNVK5b66reTpnIxFuYTeAKVNJWvUeDKEEk04J9
NT4xaa6f+nR0L3/vCwio6X1FwqwyPztliYW21xQtcqifKyoB0llgYHHEs757PIOqyfTfcP66QT3Z
FTsokKL7+QgNbmz2P0HS1dhlCOOz8kvUx81Vz/DYMDEqaIydI+gHPJ0LWd+bsDRi1aJl0gVub2kC
3/1nuUyYzCQcd6h7iWpXJluxE09IEpbMUUM/+9fhTWrlriR4nPolHBFaqm5PlVrOAPJO4E13+gUi
j4uJ8AYo0QgrdKVME2leBE+FbFcUn4K1lgCUb9JmNLp4zAfo60E3hZ36KC3SRFuhd0SbzEEQ8hA+
VmKBkq8PecjeO5mmuAqR2ZFULNDu52b3g8h6Q/RQOr7q/Ge2ddIBsMcPlLNSPEgqRDOy50UB9XfY
5z2RzYnmxJM2B1f4W8qOLpRR3BgR/eLdpZ5pKxwkwis6zvbgpg4UJdj7bf95PWZAV1iKj3E7RL46
ympN/HnfpYELyu83Vmqa4pBVcGGctaB+8Xyy3ucki1OzZWTSpF/vOWZtppULTX4wgNamx55a6+7f
rzr3ca+YsSAUrJu+o3qzzNufEAXt4UFrqt+T0zG7RqFE8kXPCIGM+cetDxQ/pgDIvjijn1vgpMvf
z3tr63Qvz22ndWEpB8zmoXuVKshW0En36SSWfEsCRcPggan/bD807LL5X+rjQTVDsqmHjOoLDyJD
sMZyUWnFvxrCaykyP0VTYjAM0IR+O6aD30PgVeZ8CNwfOFQdeGEdaZntQdbjtiNIo0JRoiZuaFC8
IrI0XGCGBeOtyMqEozws8TI8H9G+U8/NS6QQU33Eg+UsPBbNyzWhNAUwfYl2xIvTvp9/x9ochis9
PlDo2ze3FHlTWGj9gOw3dAxMPhDyUWDsN+T+qmT0J2dVYfLcyPqoOjGXPFJ69qS76KD/pcK7FGmh
pBqKo617D1vWu42pAHKh95J/DsCqpdH8/bAVderxoiv8YK/Q2I5jvx6hUz69NPpWI0hvmEEMe25m
QT0tzFPAZGy4Y3T7K0ZNPC20MzWAZ0Qg25JlW7ouGLHq0xO8vAFN+lZ4em6sWO+bjWv1NsBcMuAC
tJxj0S3C5nbrDWuC1NEBiZXs293if/LpJbUnQkZd7IDDgwishHAzAaTfTwZ94w2G6J1RXK47geuZ
2GzfVPADUCavnxKxc2jbhYJVlm+6eYOazatSzODOqn7CBNvtW9oFA41MyjQis4i2RTnY/o6I8tOm
KW1HfOfpjF0TjWME9Vf8ekpJ8y2uoRdtyGg3+96Eg1vmF7HfQ6lApCrZ/zxSphFcs9srUrk6mlzQ
2QSOh69TduCX/hGK8kV/gzQmGKZyuQ0pDuiltqClg/D67rIAzg4rlUf2JyvE8OzaKtmItYXEeh96
+aL+J7PTnBYDbmNy2BekJhoyTbyHSFBw1JGTOCcrbtOaxssQN3Rpeie/gEw5lX9PmdCrpKEx4bSH
a/buLCNXaipe/9t1gvpp7zrBH6DjMvnWTTmfCt39nNfUVacp4FdKOagexZF3VH+3ihtyu2kcFoVz
E3y1GoPU2Lc3v7LvNbm5CuoQppPUbpb3VANNU3BufpY+MzCv5KUKvHB9GNTCBn1Nhv8STR++QHFO
p2VnBglP2UpbH2Dnq2kZK0Y02VFiQ2Crlg9gqxVIf+NofKZK6RB53oB5UpL/eZtv1hQNwRn0Zk/y
1J2sMQq2YNCIHfHXCX5HEsl/GtqKgQafbpgHcThOswCyqe9D7czXTJfB6u2h9pHAbZGCh528X4jH
VVKNHZwHRQqjqvOfEZN+bg/vuSMFmwcQ7MKw2AcpgY9kW4nPM5hLekg21p+820pDjdv6zfnJmGwH
x8ylQJII0l+fLRTK6s3130ZxO44XJ2tDkOcpeyS5B6nCWNfOF+W2FbzcPAeJXUUPr5XYdZtYcnwF
lOGXTo5+5+1IYBZHLOrweJ/SRODtVKaDxdJhqy/1OtgQsWndK8lUN0rpR6DtZpws+msbxFf77vGk
Wt1mxYlU1t681KMWp0g+JfyGZZqcq6ZIrDFRhvM1MjkrIAMGKZFjV6L4aEVru1/rRpk7yFQEK/3d
6ffDpF09Q57cYuI1NhvwkTvhsORKiLY00MILWST8WvS7ayaI0MW+m+nOBdM5RbZBzPR9MoSA9gzl
D4GBJB/tB6sgYB13NPK45NZlynITtxg+23dPagpsMmiY7jXW7cCvLPOdZpyjvbQmzPHaYwCaOCnf
Dtn93RaKWVyqTNFtEhhbIeY0BW028EMA1eAgqkpuk2xqhVXZX8Eia3Tk+n/XDI+6ZI1lCUC4B8vS
cP45GEaoXH9piVoA5u/x4rFvxobD4OM2X0TY6idAVQ8oJEjMluOISiuh/APxYOcP2ZCNfGgpkE9T
iHeokSGazprAc6/cX3I28eWtyxXCGPdHHNvCqjlEAEla91klgXDZQkdI7XxOqGhitdgiLQHa6YYA
hwmilaVAcISR8Zm4q202JGUpo1W80mlnUOdeQncz0f87BTWAFgLgwDyINsPuaS1o2qNlVjAgpX+f
z5XfhncNa2WbheixYhvEnsoe6AEkbtD7yoYa8lKPIu81SchuKrgDPHzTqltJrJD+z5rwEU7UvzMW
IHAjvDubi0Tb+QTeurFMI79DiR0gazgRo+ApxkWiXZmAKUEmHd8JfUutqO2PqFcjhUitObJZjmcr
ldCY4wKyvGEYT1/kSWqJs9O+Tz2i5ViZNAuzv3Nv2+4OPiCJmKAlbNeok8Llzftlc2/ootnZn/fA
kvN8rOHQLmHKMTtnac1JmtbBjePQnod75lEsci2RiY2PeaQUPvbKtrTd7tqzoneLEjM1KgR1OujM
MhNUaZ1awVUwpoxpEJTLUoAAP2R1yrXP4Nc9DtK+6WC9OefNxkSitFdSvJ8jyzgHwpZNGf5TPvJJ
fAOSIjN26P1GxYmnycm7ErJNoOFnoZ0cXeeNv0iIryrouL+MFMEIccPtl8CTQNbmw2wJS1+z9SgD
wFZfLuNENwUcm2yiklgkBi3QVzEK0oueHyGA3//PzZzaittmvGBklYC6j34O1uNY1J4avXkY+eGM
Lgqs3liYo8Ul+mAPl0c1yA3KeEkGsRWJuNAuJsDB1wsy/X0O4znHfJ7Bb6/3Ys4hgwqeGij3ETvy
IBKDbyddpLq/oXVW448Z7csp4DwoU/jvTYuQ8B85tA6jq6lqSmiKC4zVVHmdi0dHKJuS2R7h/G5R
WSpwB9l3blikT+gYAanVNZDwgVAvQaT840iyKu6vfg8gcUEtiz0twVQjhOy2Qtg+jQNEN9Tc4mCX
7aoU++ccQJinIZBPdSFlzWCMKYBC3lfqG0WAxJ7XgVy2cwMtmBI2BHXLHbw9S+ImcNF3bDux4l8E
49RBa1o5bsNz0Np+P/yHDHteY2nV4ndEt6Q96Qkv/J/0IeaQs2g4Otb+qA/kSEgj4osKWq78XOSx
ZwdwbtgmcyMqAY42AIpS6bYSwWSPzR3ko6kuYwAitKpZWiZGdRg0HCLHX08bZNB+ClGKwLIJiAmG
OWJOmWj2l1b+t8EljYnqChmlbSbZBfmM4UwqAhO7bLAEMYjQAJM4xqP4gU4QFd5FTPNI2SMjv98R
8p4Mal5ALQlLHs59i1cQqEVtJmY3SSqQDFclemAlU4joc3p4a6T9dmrZ+G9vBmCnWXTmOCQKv0IQ
qVkWPBJD8+vZ88Nu4/198je2Q587TjO8JUjs/bTeENdm07Z7Wkav61yhW2PALmsT1U2gx8UmOk50
zuFHIjkmHiIH8JxWe6WMLxD2R+n5tugZhHggtHTpzpD/jKp9OiM60cQJbmUlbNZPxQDDFAA/i4mu
7FJfxwTDRITabdu5etDWl58QiIkzxz98Uwf7nf+q/c1ENNPNN48YQ1f5EXnSrZ3QveJHMBFvUmZn
cel8WYmOUUDJN+NjK4W3Dkqws6lwdteI+NSuEE7+7WPtQGiz1U534f3RX7ahzHQxaoY9Usdwn/La
2FTP3EeoSjGmrItadnf8gMmjqTAvjMVaBrXAQcaLaOiBol5Odm/y9KqFfyltZv/wrVpb6jTY2XUp
PPOiUitJ631xGC5n+zq1YySSIbUKyF4TKq/z5QgwxfbJERELIMrPeUgEPhPBlBMdeHimOowPIqx3
3bKEh2Ae+4YShVhjNDkDys2yT1lHHC4dc9fYAb8BhdaYjVJyZkvny5tbkM+X0Oac5l92iJ6RNbGE
H4RxmTn9/GoR7feHCd14V/TPNYljLrQmcSfGr7KXmSSkLeR0CBt0em6b3OJpNv3wW6Em+1Lur3St
njXgOwmWxl/q4oUq+QQzx6lagBJXtlN6KCMgHyjswxGC6ZsdblL7W10AGflpJR8S/6UEcLz/mNYf
qHtzb0Vj6cuhbX15I8JDvtdtCblPpwVHyuYyZTQBnTrW4ZVRy2PL5XwvyQCKLRtPoLMibOhlxHTH
hzywbI/sL3snZlSCSObh/XL9iyQ5BKtRbm1KmQnHNdakODwPjvnbWRH8rE+heIizToUUDGi+TPmV
kr6UzZqcTifbbL9aQFybqOFfYMsJye9LsbYWA21UvOcLNkeermN5zpipMAQ2+HOm0bBcntdJqYvo
6RRTiqlZAOyrVP4zRCqTLwwBecficvlwVV6lg+v3idgpFWfEJfgGxuC26CTXVoq9ddM52/l2mYuU
4smwwqTCtY0rdSJBwrMs7O85kpeIK6+BYTvMtG+4UG87ZTqpSbJvX9LlVxbJiAJ44VqZQZIdaogj
gSdxdZGxQMjBaBGFfQPzehA8yeoD7PRiBaZ2P74tt9EAESlklCO9kkzydQZ6bKCfb6P4CpOXT0S/
GFEI6jbAdb7DY8IXRftrVqybhr6n3pvuSfDojgMSLsuKpWpLLExTd3/JmyMEVzsdmFv07ymwxeK8
wQJKeyoFdizc01RUtEb5VAfApyjZVgETqzEJ46yKQeRfWvZmZZ0Mdh4QYA9BWPEpLwm49D9I1I78
dZnS4jpnUo9gl+4Dl9gG3EjFlOI6eDP7qGzz9J8viQpH4VBMYJZGb3aY6SV+R5f5SwiNDZjdAoTP
QUVvopsgiQIWd28Y8XSpZy5Euk0sgFVRPAc1miKHLa54gEan5P75Z5oD2RD7g/zQXoyLRWAkJ+0P
MWMIsfBTYw5FGZNsERyibiSpHbtxHiA6XLNKcQ+gXqNJaZ/NAmzEBWjPe+okk3PDoAVxKVXDSRWk
aG2ToxbUWhvWaZgexALcMiL/xfqp/qgVAdIJ2IXzeE02nN9601IKXrIEf7VjWre3YgXRgLYdUw5Q
7TLx9GvKEW54EfNtdC+/TEfW43o//J20Z5XPCZqmEWRjeuggzXRTs74FxVc6xTSatFoigM60tkoW
ByqwMXz3lMuxnIsogf2Z+NGfV36r63aV4aennAJGBNSabNrsWfxPY7eH1NGI89Z6LNLxOLqJeSiU
CbysT87immyeORh4K3HVjgQyg4ua3aySn6hqhIHORFTOFhxQO8zVaannq9uEiD58FNLsnHk547Bp
dfqUTPd0HrqHsbG42ualQAe6BYR+hE5TJun9ZAcbv03AlZjQZ7WN+WcK78dXDfFPoZb3BlUPVeJH
jemu4B3LJSr59EfiH6YiriTcVWlkULNFlXd0yGzQ08BuyvDIALYRpwWJAAlMLhZMdaJKMVamXqiP
Blu4erGkteCkWBfF8Bco1ReInlOyigamPKJngpHnByiZcD6LoSZOi3kB2SUVI17mi5outGLFR37F
6qsi7gsmIFlA1+zPtEF73Q2wlB1O2Dk5C40JN4zKInPz+msXWMW9pkCDpcn7czoUDFzs1zyhmtD0
nILlCprxfk0Sa0EQzpQofBEHFM21OJbVIDE3G6UQC/ChSwgysTGANM8+HQqn5+rPzIZ+JGgNNk/A
gl7Xq8t4XB2ozg/VDmAg0YPdufsZsWCKSoxY3skmD7IsqwbGVUJPt4AtV3YkUCkcEl9hejDFi2KT
oIQjGT6yTCxMlTueEWqyj4g3dSIfxou4JBkM4jO0A8OMYGbOTCJB7FooGWVc1XtRdXngrorbF/49
7sHpNd6Glt7YFj9eiwtkRVIqPtXg59hNgfrThzkYQRQBc96/d2GVvctZwJZiBRo4ua9B4qFvTUcZ
lTy3IJhYemAVSYvQDgUjoeZWiG2cgkVIwLSqOpJOUqqXNR054/nMR33uQHrCh8h+G0CyvSc75M0a
NF8boVA94LriFqna4xxyJ/K5i1x6yltbgXwE1CDYuAVETTF+CEjEDmjGUMp3//FlfWaTgJiDMc7z
5D0iSaQJvGm9IjpdUfAUP6dlwuXwpR1JvbC3vp5Uw73AmZ9s0iZ8kCzqzJzs4+6toukfnBDnKKlS
2/0YAWPXlh09xt1447TJfENhkeVu2rlHbkCP8fXkul/wNRyT61tdvZHVrr8xvbuI5k6e5pdvy8uz
wGlmvjYXvTITsmER7SS/yYxmk1CvvrgWlxgF72QeC0MlF+g52jXzwSNk0izcRQr+eul9sNHL4LsE
rD0VjhLo6nNIxsIhnczgkF1DWFmY8OufGA1B0YFjpLi5s3UCpQOSRCau/YSdczfY/5i5rZI6STw4
sO23qwlypdZufJ8w8p/6gz5j53X4XZBJGSHq+0cu8GD4MAtDOwrLdj/nxPG9DWluwCaS7hs4xPzi
Q/PGXhD3FhpBG3MtBGBwGo3hliGCic9jRkVWO7OSf6hej/bsltD7MIJAEFmbk49AkYjWs+9CLIn1
AlCiZjimkfPQYE0MUq8UChEp2BmCvzz+03dco2wQLdJ2TVrz9y6UK6nkrZg2zOw4M65KLobeZ4MN
CRhHQjmgMN0uotGRx43Q2i2XGtotf3Wq4NNJm855/SH/wu84icE9s+SqzrHpt3c8Yto3gF52QVYC
G+xCafzyXeZLm7e1xQctrs+t7uaiQLXUY8iFLNyjJzuMcnW/hbJ6MIddlMjgn5KS/eM4G0maqL80
8iK9ha/tC6zn/1nWjzrj3PSETMGREKCJ6Fx8zkFbZ0JzAgu4C3YHm3Qeycx3pHGnfIJMeTYJWyKe
DLiPYWxgo2o2XqzsG1h1BKUmhvwWeruRs8nzgUAGxYVu0fyfBWxNt5F4PV1ZxnqTncM0vov1tL3w
YbpbtDcSS3EkMBy6v+dPBfXzraacJ0vc5eEgQ7cLmAPaAmWDEmlgJNwNmOuJJ08X1xBU3VGBu3yr
BkhLfcZzgq5SjJv9AKhX4H67EFRRlSUMQhGoDbN6dF//gtiFaV4mV+RfDmSjvmSufNmezrFLM1tY
GuABd+t7Hl60PqhxDPEdeamf+Fsxlxl3NXEQZr8HIsmZexXp/XLbMEzIY8Z3XuwbLzHboOEpOP90
/socwWuMpFGVYj0adVVE7ywnHKFTiFH3/6HXZo3ih1HPYjjolPKnFrrJKI6rZNtzs3eX8vqVXgCQ
tERczjnRx9G+EjksD5LjKg7x0JKCnIR+m9fAEBKtDN8zBlBttacHpmnBJlb2+FZR5wtbRRMZg7xG
qpi6zLfz3xgTYhhPTy8vmPYAeeCaMhUGh0EXIm8aj7Cd8bdCQJbsiccDSmgyhV8bvNDiYsVn0io9
GNBfdU8GLQRRU34XJTkgFYzShS28rYkBKtgZR7+qRn/Q4DWJ8ybLotbu1QbkpvEMpz6/Ps0v3u2x
fecj2diiFRvKOp2wxtJQk5DI9V+5Cq+Vgyhy5s8flP+v5w2MurgAU1r9AEyLPNhWAQUK9Ppx5Xfc
W/ZydcSeMl6rQLVTgfX3F+FgRCxaRmKpVBUFfGLUsBwHETw3SVqIGVG7mw3+0mXSucTl7ZimY/qO
EpLs5z8v59U9QxPj9jlLotobcJ5wUPz7Ztbn0JvWHpEjWZqCXKLYGtyiferwGqmbdJpJzVIvrOGv
n30e+6uWdlChYk0YMGBtb6+0xLf2sQ1CdPZn917pgaAu6KE8hagDYUQZtL5mN/P2sr9N3Uqwf4FO
gX2eTfsBzngUwhLLcM4ZLV2STOLkif6EKEGcuIBgKlvyacKzEx22rp95pWbYf4IZQ/UpEi9v5vMy
6zVmP7egQmEd5Zyev3I2NzOLVhISI8VM7aDzQA3CoOo5PdnUphabK6Qzt3qWEywlQMAA57/rWhCs
ymcSWzA8HbEYLXlcQC3ep/meNmofzpe+9VyKAmywuPObw/5FMjZXvhohIiAaD7zK2A/ZCxe6iwF7
NPE/kqPkcYaP+E1LOHL+QkmY3kx20JS6k36WSWq1ctDeDVzIzlN1do/XKYeryjJmCN9CZx1sFKP7
WF6olOlACYvIR31FsVapIl0VncOLFTbkVi6SejPznTKF4plnHpK9yVgxCoV6nE7rSgl9jRQb44XO
Y26uI92KmmyLY/l68zpvTci9VXjzfWsaN9OMZeNcmyNEJReUA/nCsykzlSyH4h+cXqgJ4vFj17HQ
EOCAg69hRxGhdKr2h1ZOrV1kBevZkMJmwsdc4moJESDfKi32bC7+PuwoWK9Cc6cLRpLIrg0Lzcj1
GhvkbR5dB2kHmKyye0z6AwCUfpPTsbDNen37y9JsDrzDhLX5/XxjNeoVZbG5L+8vZINZ/J9OEBWo
TzybbAKKZhHkTmfj7K4iNGhjPkcfUS100l5LIQr+4Ecrjshnd+yZJRJPq6+K/vu1eTrepXKqlnxS
zghthEGOwfNv1Sugi2fpXvwCfhWMSw1ixX6F1+h493kZwQ17JgJaK0HoH+U2xoDdbiZmIoJ6LAQx
5T+wyxFLs8iyX3AFB+dR9kpX2t9t0nrfHJSKIkoHL1m7S1cUscK7W0lW49TtmwolCy6XrAMsIePi
mZDjPJuLj5lHEsT/IqhicQ+D5jn6jrwFSeNftVuP663jtgEpqO9s1WIPa4jkXbbpPFwOAr8QdFz3
BaJbaUjuZVTBsN89Mqw9WeoHSo1qA9FEr6HnbDiZZ+TY0SAlbHi0usvsvDvDrdimLye8RKu14KmF
lnnT5XK8IxDTU3jgYzj2YD8tmOjpzGauyxqv3blv0c5RuzDv0xXnPyy9j/HwUlWuBt6GaBdcIJpu
XkJyN5SD3WK/vvzSBULKhaysKfnfp/qyF9KZrGTFxnOzivCYvDdz1qhkv4WmDq3LFWct+inSbHwF
zRH8kjATrH+Ri/bYVkNlurnLT052QHWJCbpZKdg+Yl9h1PgN/gWXZGujUKziwoyMu5FVCIgdUIcJ
KaKo3VwOc423jSvrSWTMPT6hCnhzgEpYe+jlEhz4HRoIkQDgEsg69bYRMTGEyfv8FVoz0+lbiy2J
spyT1X3inKrpZw4xt+OWrtS3IpxhdqwwePMh0cuBFT5wMN6FJ0DX6e10/WPuBO5pqdJc0wQjYmg3
bD2P9pgvJIAz+NbEoTCMpYDx/jWWDkQYDPH/Nev6a6R+2HHcaM1nI9F66xkdW/y7sJKOqUGvtCkQ
CD+NX8zvf3qJHvErc0fUJbB5RAuEfjV49tOxEBMWGrS+tT1BBbGhMjj2BE20GcMs7SlpjMZQ5ipW
8jk7mCJ/tOMcq8KB1jWbOfOtvb37qmrfZSJw6WGsde5wG+SGPVKuPK42fHVbRagAG3b+ynwQMux0
Nyk1SdPl1gakMy5hkgcMKrvuHJEB7sE3Ob1n4eZE0j17Qq/UlcchNFZxqFNh1UBowqRk8iBhmgvh
2cpwfErFP4M2NulmRGAexIV237UtsPeYilZdeaR4nnmC7eThF6uk/eSRzQV0bLQKGSoQ3FEGEOhJ
Fn561AVaY5+/MyqK2Y9AGsfEAle123/Ky/eywt/z+2NuLcCEyZujOi5B9AgEwrfLZMe/Ms9Umc/8
oFTE3ODgxlGf9RbdQJ3WFKGxVJP8L+Sf6qHEuw3jbLbFl4ZtDqOqrfmcI5NKoJKpDTl077NkmvM3
SfYWQeZ1gFeJP5SEuLE6cl1sd8iEfsctJAJKGil2hX2UmIuTgTORCrdUpDyfB6fdrfpGQngdmK2R
ahqDsi3QD+uEa4swS0Os8JRjAlxJqDMNjTwNKd8PfmQDPxhWsuIIbgeAaB4lWYeHOXPhdj3/9M46
DHi3HY/lDmd3WM4TmCKUGB4pXlHuh0WmoLqfU2ZqweYBmvppcCwUrEKosXd20VAjHzNQbPvsEH6D
E66HP0H9JAxhO0z8Gy6U7BWXHQbQwXYgOTmoJiKmBVSf2M1stImrlfdh+EY7x8FuARtxjU72m89/
5pwUFHaxH1ieeBcx0CAa8lb0WQd9xWcUGZLx9qIJnX2V+7CTIZbGecqC7jd0fV6XNGXEvx8HBcMW
9+HYE/MSRxmdTM5qQBBW0D2llFZhuFq+J9TqEh5XvM5ZHDn+QqwS6P2kDFRgH4sERs0gBfC4LgGw
um+wkKb2U/2J+oegwtL5Yrp+E5E94QR3J82/hts1waIkUBMHo0WwY629eihImx66JVNH9Kd0wP7l
h5bozORmvMnNiHsdXKjy3A/y80dHsTIqorNSQJrqPAvt9JnQGxpkxYgi+3OOBTJub4KIp8rEIMXQ
N51ahbXMSaoWHhZl+blqvE5vwZPdhGeqLAOfLZSp/Li1JZ3VJthlaOziFQBu9OYSxRELxrPhD102
qTa2/tMaTogdCILXJhIycVl3vqixCtfDGeSGWB6Av8xj0HMEckKpa3NASlI77ib0Usua+fcz81/K
k1aTyUysuKtdul3igJYwYTUhh9cmRHi1XQeXKoygPfUK9geXXpWXy4Lq5RPXC7vPHxNv+PcmwUyt
oJD/HquVZY+abcSNL1yasNejevbMagr2qDsFy7LUsQ8Ytnf1rwKMmQzM7WCkOsAq6b30pwhwrmo4
NIK+wBJAVyFU1133hWBE7MKf6M89lYntT+f0Aq4rbTI5Xm+MqmWv5s8tQ5orY2m8aEVRwCnG9hM7
atDGWQK15FLC8iiJNuw1QoXAsqvU9X/qYFepLd9e97LLyiZ9sKXbwX5viXY979GpTHBSdKFgzjaT
VIsoqWxgcg8gq+WFF8MNQw0GhRFaqxgLhqUHr1Frj1lHFP8oNQh26ZX5H4/EEFIJFMcuyUcSElYE
wWTO5aocWxFIRW6gnTddAdoNq5BnlaPZ1N7x50AqPgzyD4i17e7oW/Ha+hMA2d2cIBct0y+cfCe5
OBckEA55fd8cXpbe7nGhTvGb/wHZlkCnmwsswjvOGyA6BLiHtmMRLd1/HDSns4ZH85RPPbdXx5n4
AmsTBM974jjC+Qz6q0yxPW1o7kBul9wumm3hKThLcVgK+LtKN5yDXJYNGUYfOsQHckPFlld1J4ZX
nANUKRu65WKxGVrauKnIP0+IDnezjEOsvCLpVo/6B6MmUCedproU6oyWYvHqSodDAghupvRfy8/X
HpJpbqcBCzfuNcZcEsf6RAPzby/QHkcjdh1BT2CQtptR9/JPYRlOe7uUUaNACJFfvCfVUNINJzb6
8tKgx7Vg6NSu9yjbEglkUbsR1IpzWMB72XlAtnWSXBIaDhtzTRq5sLHB2D+KfsXATf6WaHr6Ud8q
QO7dK271Wd5J9CqmpIlN5AyhHYomaMxp+1pHe0FaqIDB0DsMtYJS/Hh4qh/pbClO2yJB15RLC9ng
VaOpIv0U7Qc3vsXmWvfGNEhGV/ToYNFEoo5m70+yMX8ORu8yuqgioX5SpBdgfk80yH/s0gE6Z3V9
n6pizSKVqLcTJ+x+WDwz+51Cglzh7DhGXLL9MBtyFnKE1E60w7DwFESXo5Frvz/uqCHIZ73AV0pw
QjAE6oEWgwc8r9I8vNDkklJqauCpIpH8XjRDTj3dr+5pdsg6/vQlrsB6swx9wi6SJD/3OsB9T4Xp
baJVnM5iL6ijY0db4q5ESK5rD0z2z0t7AFejzW4Kb+Mcdg9lMqaD02IS10XNW2g5Q5p4KBi/tgA+
oebdmqZghG2H4RoWxQzQGj5qM41Er1E0pKhlIgNwplT+QO0x6fx433EWNcU5vcl68mplTyWH4A6f
R+nuuv0f+5dYWmPKjraZIIq3dqExokiffqTmjUScqBsK210xBykk1HKQ+W2Tzl1EGXl6ipdCP5Mx
xsN5/H94pTaKLfTh5oRerYSAfrBQ2oYqDtPqifKqCrIlzKpOb+IZvE4dGnk93vJNFOBeaZp28WQM
fsuo6A8gXGIXfu0pV57WrTNpsHPhCKhc27eqS1vneUzDVSBDPO7ixmNboeJ/ldnBJfmKDodFRahP
4gMVBa4FZIYjtW6v4h7635jggJREivT/uDSUJBcS55U/d33bk15Ih/FCth+GdG0jHAvyeK0wlMyK
y80OZNQoDRbCh9hX6i9zgi5LUL2HAtBU0hXP6lBw+Ovtzo4PIbe23lQS5S2tVliCFj45s7iYTNBF
WjxN1ojbohmO2oYLWLoPDMyonc1VSZux5nby2oZSdFQnrrh7/czlNI+WqPD8387o0/OIQuGNTOJV
fmEXBSw9Z2XGVB62aJRqI1JsZ8qVEIEw/XogGCn6GFAw38DtFxje7X3CgSMqNg39sXqpGCwV1ixm
4iKzBkUxjt6lQknz9X3+mQY66T3q+rpkeuU7AYuJaupTGrqLLUihaUsNfWoaF1BIHN57/M89GEt9
7uc/Jf2XL2XsLyk9MQ0u0/WluHGjQM28ZAH/+Zbdy0oq9tbLizs9OD3jwYfDjcu/VQi0DpNUMRYR
4UdIjrNgvhXL2Dh4VAuYoYVcu3YzeQdnjML+KheZWwgYN9lIwguQ3k01/SuDUa2/yC1P5nLYgoaF
eesZMLRSxCTpiD4Djd2je/qZ6Ch37BznpVpPGjWW/tIxAPnyZhFdHuZqRey81UW3D5eXmuI8/AAM
xv1RuN7ZGrBMhdF8WLvZkMZh3StMyXTpWg/c2SiMgdThxCvSkenRtkEVyGpoKZwsXCH9v9zwPsFc
jwD2SK+0Kn5dxXPNdn3b2t/1A6e/qFht2W8NjLA2UBHWkbyBJw53c7r8xrWD7KW54BS49GPm44mA
lmdGwiDVZ4E/onExa5vVEScu8J/8LJb/z1krF9rQn105h398Jz9p+JochptasZQZZNCYW9DeFWAQ
J+VuACAs8gmqpAfhUTsSUG0MumkGm3j7XIGwboSP1SvsjEDRTkpmN8T7SwrHoQPVLrCjJIg5ENEi
Drrz6zCZ/0gDRfBTpw2+coX8oXIyw5MV0SfvDQvrcPfHhokve8Gah1K/XkdZv6tK8GhH+JrYbvKz
CEFQsnP1+fo06RwGXZVKdVj/mkjAjaGg9EXJR/RUGYzXHUA1zegnbOJgC/QMRsodVR4cgzw7zyvd
lqkdsCfZ+dcxJddmvNQ6+dqBejUweP6pZQjS2A1fPnb8L+X+P/ZXUrIQxfasDNoreCxAydFjFIQn
eIpJTw8Z1D38sXp5APi3Bxij1eBe6PqFJNl49hiZZcbjq5TX7kYsZRmc+KcJ7h9xEsUGcIn332bh
KRUkSak/YvU3lmwu2HxmWeyC4JsVR4rrgfD6p5JPRBl8WrlN837NI/LnFyxz2EaATa8bMNG9IWSS
DySPFplXURKiVJeK7QA30mQ2XOutfGHzkhIdVGhdKSp/xKDh/YWyjapA+O24wxr1dItuKRiXWWaP
zZ2kA8pe22ophyhfyCDJjgrywY6Leug1BHB2d1gU2Rm7klzaxvyZ7FPoM/WPMm3jjqHNa0F0LZ9u
vZWK4Keg5VGKYxIIXLpMu7j7ZFC2S9M9CGjmdPpoeV6GVWEDwaLLtleqFEw512S1kMUMR5sw6Amx
vR4WvEUYeBQ0/Rbwo4C1AbFtdrWndX2Nb33veOyxMrcX8L/1Sd9sEwzBGaKV6XQrJkA7oc2YREBt
Y4zMVtn/4Lsf/2GzomesVZ9Os5gzykPQG9TS/fTVS8WLtAEKFkuPZb8/+j+gzRzaHBi2dd5CL6Q6
ZkEEOfjyEUaflb1owaMYeyQhldDje5LIC9UTeGWtQ55nqqEYsIES9Z5Wb/Pe0YBN1NKxuMNq7acW
Eh9boUSZFYyhe+5Wm9gYYs19UzACW8fblR/BhV/kUg6SwDlSANs5xmFROfnXxUxpQSrLdqrDm6mc
DFdvsoJirGZhPAzD9nX3dO6L1zSgyXcDHBpjxWSZJO/lVaA95ua18IHSQTrjNvHxYAOSroGss8MB
H747IboGTn80Ug1sbg++xG5c8D+W02IasdwF+nRBswwDhXgbwlgh0iqsE6MWOckOZDssYDspK4xd
6x9m8gGnpGLyr59m1Q1J7FxE2PnlYDU+excu40RKeo41YxYs/Wq1GCxFJ+YV00yJxKnspuokoCvn
r1K/d3zjPqd0Jgn32ZzPN7KQ1Dt/9A4UFdhObEY68tpxu6znDgS5itMYfhV56XVSpJNeEcPJHTvn
F69ngzbx8+dFD1jBjjoSryGbiPwfI4PXDcn3T/S3/Rs0lAak2H1rotB08mD3oCgOZob3MkjK3uUz
OLNGxT8Xmw9TvC8TWWgTlnyM69xW9BbUdHT/5i+hghlHbhiFxzGYQrF+yWM436ablipGOVoFJiKW
FBNfOrI01jkTAStWWUHjQp/TDfFVbI+nl6105/Yxk191gN87xSWLdT4RKL7hnx5qL0VxEPB7yVcQ
Cu2K3ScL9AvV8K2YLT5DRj25PS3i9aTcHFU35R5D/euGOcY0WnON5JBbjuz5Do9aUcjQBAfjRzRQ
Kh9Bwk2qML+M+fzBYUtwIcU5fh6ZxbVOP1xPcldlcMVBOKjsRtnNf2lNmzeqp7EiH6slf07zECM5
Ih2HNP2n2or8KrNOL/I6UrjvMyforDJyQT8nZKJERunr12XMHlp2U+QKlrdQAVwz2U+wpnrMkDsA
R9+92O6UkACpJU4kTYZCKyJGV/w/krZptmtZdd6Ik+m0kauhS64WsRCnxNknPLo3whnN7QHECiYR
CoybD0z7pTb5Vh4N+svZGpRMa39FlgyM/V3/Wks85Aikc/u/7zKNPYS7CmBOGZIe8m7iXxVDOkBz
vlsOy37zoeB/+s91EKAO4Qnvr7f1ikTC2XgGBrRjV8FQQ/qpP7ns5csxWVg5zpKM6UAtZM3aO7z4
WzqiRmnEgfWi/v1g73xvsyThD2sutoRP3lso/6UrVdNqP6M9V0FW6ELkBOsNRrXfKdvv/YMsJTOu
OSKYk5gUciSzQqlWH/2W8FT73ZBOXRzb1njebYBcv9dQ7rlac0h/R1qtdW4Cmq2y136uguCgjveB
7kX8a39SvR4uZvjumsXFJJrqcVD+V9yIbZbKQ6G/eV19c1Aj+06lMj5vmy0HvKLGqUONFl7TwZRm
5la7vIJjBL5Y8o1IBtv6MAoBrU55ticfn/LZrd8sQ18Znda9PAEUTrzT0XnrusYbegW2PwK41Q6+
69O2vGBgsUj2s3Wp9u5rU0XNY1Kr9hN6zioj4nssIiPnzjs+vwbFgzRKMTW8ghFrdarTnxasdVxz
ijcF0OVLW8wTxtA9W/zhKnFcV+xN7bz0/lLmwoluNTA2Ye1QWn/hrhyngsJaZVSRV87tdQ/sRZ+f
FvNIVL/MJ3rqSbMUvPuCgYyQNsfYrcCex6MT8PUlVkAmDTO1N4odSwWJZLxUGvV5cpewR0vXP3xA
Mj3Qswke7nG4VbgWhQBaV+6DQQalSgjiKd7zmV23wgyUoBcjjyw9p5/JYJNtGOkCVtcFDsxJB/xc
cBzx8J7fMspxvF1bH6yyu++/eYBHspXUgg3GgWSHoXyYc8KIERpmPFAtyN9T67KaoM1lBP7CE/XC
Swc34TFQf+KeCD32RalUKqPU4OY+4Ya4PqiiD/edXDuC2OqfQC264mGwPDhTB5s3Zn8Z3a5KRWJZ
OyQOeQTHKnLKgRFIDnKI2R9KWluorYrsu8h974JQmF4Drj/UxXlPi/byPUzq1jYNQ7oiPLoDhgfz
HNwet2eGyMT2MecMBXi6KdkJkEIwd4qc8ZJzCmYOIjtBscHu+bj63anM7GfWfn1omzYeWC1bSbLI
Nz0okc9qxVv+SpPLDTOgfDF7cCmoMI8RNtDAfxBuy6f6KOHpHcW5mXxNzaWIQb1OLvw49z+0oH5f
LnEkzgBKEUlPNgSTmbPuYnNzqDbqNKL11Sa5uOC3wk/rUZSCB941ye7j2fp5wBzCXeMWylFkWYKD
oTWjSt51ryR3WXzGQUPPxuYliFZsVbD9KMx02Vb7cQyzWd3nKFJeX6UsFcbTI6cC7SFSCvdUlOBU
mfJ5B/9uTFvXlbeCHiE1WuroGJfavMK2KCF3IsS66z9tr9NTzQHfA2kOexH6hlb21m8r+el1dXJ7
QzBJW/HilJ8/9scad3Xza2nGFvV+v8oTZIBDyE5D2/dMor+HtLZ/Gr1HQRAjJ2aCdTp1UxW7zY+W
mSrNJ5cSFtnGYVYgb58hAjwhTXZE7KRlyVoEaLJVLnR17G8x+KCAZEed58d6pKaDGLpPHjj4mCeB
49o9OhhnaUwqCmHqs3KF1bCGMk8a+N1NL/ZXxgAxTPX7BD+v0mLVW8y9MS1ICC3I9a97l0JFkTuN
X4Cce4gKxY2mY1+AoWd+z1jZdEx9gKq2Le2SXGQj2fFknLiVm3W+EcmDR6I1hsM5ro57B54emyKh
p3ZT09Xz+d/yOQK/DZqnZ3TgwBl/RAChGeTw+0g+NxsNcONyZ28j7654PoFE/YGfpFvaZjqHcbUa
RWWChpKa8mywaeWg82279SCeYpOIS3aNye43l3nR6xr3G3a9goy8zdXbfgRUOtdtVHzvxLaR2+NG
WsZL0AaAmMvF2I5srUw78L0hce4qmKOq6be8eApTGbY5NDikOGL3HM1vtKkDZZAjuhWiVnH8xbwU
P7tssa6f25mz+B5LoEYKFjTxFYefqqR967DBn6LzfTixrudTZmP3/VqCm5siliDM+HcA9Uynb3vj
AROlDTNI41nhpl7cD4s5r2TsTsONjL8Sbl2S3AsT0CLiX/FTvrjh37/ahyYt2WvIKr4vqXG3Nwpu
RuPlr8iSwuIjSPxEvsfhV7hI/iKkb2dJo+Wa5fghoJDOM3bfr0E667zNgHrm83xoFR4OPn+mLnH5
yCan4Q6kWQgb2LYd4a2EXuOYmwGZA3hLb8kYnabaQ0ynYQ4kJSY6281UioT/12vbvZbhr3kioVQp
w1f+ytsP/3AKjFnWbits+R1EntfUQ/HfW48qH+CkUaEdJ0HHDER4dJjwSqHt934t9t/RqmI9dRQa
stls14wZFgCP+MhkEnVXU9ic+ePvHDwvK5seHFrB6/HOnHmCp4CwIZojLHovyiLkaxZXwVdN9oLm
qg6JzjTFkyeOJyc3IIGbU/u9hfzI21yTMq527pic+lFf5J/A6Aa+h/DWbd5IU7nzDcDpPDsxclZI
KsUjtG4ayKP0CBnRIKLJOWFCrreuvIFCyF5QsO51ieaQW2mCHMfHLyI3sEiLoGlvoOrLv8hH+7fp
mIM28iTgfxNQ7Rqf29pgD2OxWIHv8vPch0R6khow8Swh4IW3PTSH9DQttlVrUKPxAw4s6jX/bb2U
Jpw7Lt2KRuWebCfwTPIiZXhuMEcSXrq4RCX/qpKzN6hPkNJ/2aVzAgQf2BUTcfas1s33pyoVuqcK
9tR5CBbM/ANzVrmu8o+0zRdOeMwvGqQRT0HwUyqT+CnFEh6/dycTfV0oR9jiEdk65f3o6ula8YQd
KMWkXTfFM53IewlxoST4bj1UlfE9BEUkDyhZhQjnqPATHv+4/TL9DyAD7FAK8ithgiUxOHeui1dh
mTY7GBx4qFOPmhfsLT/+H3v92Wf44tOR52AJS4AUrnrFtm3F8yTtRX9HcYl/2AUYvyiBD9b8rlYr
YwXbPtmUl4nML873+/6fnsNYjE7S+UPepMqNQXTcSj0d3FrHSk+Y8wHyacmoGBCkFF0fYtUgXcFE
Q1JycRvuF+lzNDylemjXjxQPiIEIyWqRPSgxRwri1v348lW6PBqTzzm5x4xEM3jKpWN1EAgELhuf
NxdTW+4cBadTbg59fhYRaLwZWUlkJrhhuRinYubERVM4m1l7/HKduB/43slQibitoBiiGhiMBqqn
Y6i8CmSQS+lNi3HVLXbM7H5FChttLviuWWAZHT21n/zoQCt0e7thCS2wwYvwB6MjHwOnlkeFv5xG
1qMwf09lLMbeFLHUbJztYW12z7U6ohWnn2BYB7i8mbSHUbcg+4GjGRbvKYYQGK8PNIUUgbATCDXJ
l7O40HjDf4JxF1kfDySoVIYSOYALuZb6yYR2axL5VUzR7Tpgtfr8/TUFTEme7RKfb3TGXECSwJ2T
rdE5lJWzXuprfssIOQUvDH8w9uSG2F/eQoXwogeUBWXJ/W6Gt4bY4GAPk4kgCceeUf/Wn/j5ilgd
b0z7/3i1gAZkE0QzvuXlj2GbA1S/uHr4pLCutkStB06iSRXB7718Jezfn4RcBwzcQ0+9mOTeuRCg
6gnFLZvDh7jHaXPhTyp34DlGbv+lohPto7rqytqp2YCylhKUxCMO/S5d4zDwr11n5WXXVipVBvDI
/+3j333F61gfwiKnDwirJqe0i8Znzc1Q2c76fGSmAS2F/3g5S5kAOOnRjy0hRSQigAiTwPdv2pcj
Y/Mb6nEDx/Ffx3Sxojl8HeNSCZ5u+hrnIB43kQYxIG9CMBdao3bSxmBNhed3ALYYH7AoEQjMLyoj
R+56aRPAEuJjYGmydvVWv18lJkti1ae5Xjq9VD7pLZbajywqZ/+nQ85crtWA9zeZ66urkSa3PJ7w
cOIqtB5lad9Fd4RqtYH6VaQjcvWHDntvpr3ODGDxdchjz4zFud/vcHgkU2sJysgRTUQ+/nlGzWqN
o4Ca8QHEE9jRAMU/Y/hoLgSZwj6YLUHb7f2hcrLItmjaXII+b21PKAs2NOuTy3/SMtU4mR7mhazs
vKBeEzHmUZFffEisjLgMeVcIcLpGbWyhrGoHxbJOKkd2dQq1W2kXNy2nbpm88YLAU2JwkNueH+S8
rCVC6OxeuzYIWEjZ1yGL/b/aRM8Su7fbeKfAQEfO7jfRzfTHEnHmsAiC4VfgYnU6uIasGtB8i0qk
lWAGds58V4qfY9XbaVxPSyT7pySz/oy79K32S+HZV9aap5/7jqppDSzS2UxJPwk9aJTPldx6/HOC
vi1zkdgbnP7afu/NaTRTOuSCnE7PRjl7Rx5puXTY3hVkMaXFjUw2nm74CWcytwC5J2SoZEHXMeSi
sSOhT/swKjB6tibYsWBCIORgvLyMTxo16sXn9asykl/NeudINdmTNtXeqrJuP0tpuG1+EfH3bHOn
jpIbtwMxzL9VSPpVoS2286xjzvB1eOUZ4RMK3x6A/vQtw/gzySmRPqnHweSa+Z/T2hgZw07wedrN
BewtdaMVj/+wYJ24GVVw+Gfs3CZj2rbfXf2y79kU68dlYGFkxbjWF48aBjhJu43YA9jKSy5MZ8HX
6fS71iUKh51Jd8h4w6z8E1CTWtDsffR4HggoaVq2UZtJSIP0d2+mX6xrrjl9C8UZTDlG0X7GgPw+
d+sI7nb6H5LULmHT/pR+Z7EXLgjY6jQ6W4iADtPWxXCW3J0CnnB7PZc7vFrJpWidBI7C/NwrUOa8
0l4LoHIltm2c+SfCA5noqK0rl9yPJ3vkkrL17drts/ekRnAvu9EfVSBSSPvsOChPBqQSA1Zcqab+
cRrbqZe+HDNmhzPuVL/NtgARepMOjJI34wuTVs8dcIZFThRL4MOAorMV3bPWkpbhIbQYPkvaBe+g
UnfbgQhNGrQaH3MsfOL6gWdFfT29jVZzAEHHk0RHiGUCZKjcl0K7byPnxAme6Pv2QslDfaYfScZR
fs+0aEXa7GSoF51ELeuXOnejzu6LcZ3WUAoQ4c1sPNDtMLgcLIqgEwBW47aJZpTJ3z0SWT5D8Pbr
7Lqt/dts4scIw+ZaPIIuRPJJKZyiVvd/RYbBjhbvoYu7j9BVFCBugnuu26IVdDE5aAo2NEXUM6Ez
Xhg5eWhU0lbkSsWNP/55VJL0TiEUpDU0OoW0UhfYRIs9BymJxgEibYqf6DeFu33m8pZdF3QXBlbT
ow1Hc53Xz3Zs/9E7yMexNXp+6o81ZOrIsyRbicojYXwZTVp3FAbt1bO3X9VDrcFyWJjYodPeOekc
mmJL6xNUt68FRNVag4xHMr2bZcO/+rJFqtP5B+GxwsA53gLsnogHPMKfH4GgIdwmfYCwPaliRH9l
ix5c1S3iJvYwR7qayOF3gdDZbWVEimD9Yc3vDpP/E2hYF9bvBvGL+RBoLUldL+m4n5YKgnd+tapw
YFQB4XcMevru73uuLbb/VYNfo9MJjVek1ESU9PiucmOsZjc/lneaQ5bQwB0dm9so1BrxSJCjj+Em
k2GyHyBWQH+/L1xDhIgLI1+kY3+0+doowDBDzWshot4H5JdMElzZtAYrm+WYPL5sYds4JLGRMZe+
AzqCpcGuhwyYSPJbIToT2l1rKdTPLUwfKGfS8oz7TXBpvkatqJ2LtIEKt0eRVBbnYb5Oi/O6nGv0
JWaOHsH1WXSZ1qc7Z/xqrnwjMUbxxuGMPHdJfmW/Jl9YuFae9ab6Fs+Kk8CONadiXXcPJUo2n48f
TKns+smzQo5GPLacyQ3WJ9xCGQG5vKZZgo7ddcNopI/j4cf5+GtbARJRbMFCuKvKSHblaX4EiY0i
MmfIbslV8RwYV4hH9LCy/YnW44/tjpc6p9Wfgh9dvghAEsBP+XKRwOLePUh/bUSJ+fXqmsh3Cood
caOXOCs96TI+wQpOrH8+3CfuyrpMLkY10JSddnCTAtJ0ybZJhEDbkMjUEJPj57rYa6YpfFhr8f4S
7wZ/kADugFnWt/im9NTLVCQJeqpu6M4Ypw/3z4RVEHfZUImveAeSwbWoMn7WGHg9xKEoZbJoL7n3
j0/AcL7Og8pIxd7DoYcd3hSrO69xJx0M4SGTq6JsEkQg8CSIHoXVvjK7I5OXEnxMDDQwc7h+0pHp
8NPy3gADqITN5pnVeUovLNh4oCpk4Efn2FXZCNRd9GuH3rZKOtR/JU48bkMWHMRc+N2okaQn/BbX
EOX519umZnrgT3EO/5fni6b65eWUui1Bq3o25effb7BWZT1daydhcqvPp3Rh6QFy1PZBq1guZ5Rk
7AoeKrP2X49CUo0xCt0tacJQuwA5dkYioLKCVxKUd9jDcWGn+1eybQYV+8aNGstXO23sEulfTq4f
T5F/5Zq/KC6mEHtsNPnrLM2tKgVbT76YgtwBXh9X/wVWydxkbYLWVelPyuUsxfzbFrnwWr4rqCE/
vDwiVcz4TPX4QCbQLv6FuF6ir/FYHItaUNnZqThp+gbfThJm/IFaW18VwYbguMr6ks9GArEcYgy/
y356ziaVlnbFTw6WKOdqpDXgqVjwh3Cict/HEGmd5Z/XPYh4flkBnjOgR2H1jDpsVhD3mwkdU6CC
k5EDAvmw2aAHik3onK+6XVaJp+TBQkthE1kkx/5DoP7mqnOGKuuBZwnmLZVIwdwwjsg1e79zScUO
H8zYN8W07WMJnCB1+NXxsYpjOdPqTtaoQ+yI3zDQgrYE0ED0TUFUv59zBg0dul7tk8Azvx2qmavv
pbNyFCXC2bCLXgEqDVnRFcYeSvuhGqP+35ZbNwAT9redxSC3qgHAFpBgXf0DZjpk1uLWye/S2gBx
0wWN+j+81GdHuJ+59sbBNW2zo9HJwtuxFd8Ev0uzTmPX+poRaR2wXmiq0Fm1BN+exB5DM6Wo9AlY
PMlN15bG1z998fkKWC50FmB71e646iBgX1rtnZTeHmcvuTa/2CfGlQEYiFgq6CeJ2vKc+MsgPhCU
muodxonhdD7IC5KoakIfdesTxUoCrKNaZueT0rWSY7R/0p/9EKUmIsmXlX4AVIsVeXAsVuDETVXG
adKMG/C1PVxUtRllP6Y1TdjSH55WQH7JcFFDds+SmPbt43Fq7AXSwlrd9SP6f+CMydZDjOXcUb8e
/6zFsyav93hyVP/mK/lj5tIlFBcMAxdZXYceL2l2gLAWQH3Bc54lhC3pFCe1rCx9LLkiTGPwpRwN
Vkw9JJg2onrBrH5AkX9RurdmYSa2qmg/WEipA7mcdQcOYsQrh72U6xPCxylx+gUCObkgq34IJBsT
L6l9S0Vq5fhNTi1YlRYnjV+6c4IRgr0gef0dkrvYdjEGwj3OunBsHgQhbkot28ZduMR8zvVdP7xN
fnoDcGP+4DaADM4yE6B0PRanfBCIYvjWDmLkCVZNNeM9Wpd7Dw0ZFG5f9RMfbyrwzMhR1GVrN2cg
B3Ii1oaNJ9h3Rdzt7suHasuJqyHv5tnYd7Vj6uheHmtFK22vhVlF1ozlvka9+mWCwoonxHjf8xlJ
/rdb8DacyNKlfzeuU6MtHi8ioMBLSPokpS79eoZdq35zRW9tUjGkMyYpXNEonYSwtUg+jbvvDpGz
NdWeXPsakUdYy1Fl4ayjZPZRgVwGZ+59yVaf1kW7BYKFFrwWaQ4g9Z11pyKIz9iChghoQWn+ozGH
C20sXH7uW7lNm5T7p70Wf2bZfcAQKFdAVYzphdwcguRklRyq93v3JaUL2x7NsR4CfInUn62dj2fB
1zEW86UiLqJRyTpNGueUL+Hj85Clq9HQlSfB1VuhgrMClguuGxAAHU0ffz/GNCjnTKPgTKInvjIR
z7U151hcBz5KwsRarThqvBbA0jJVv17VyDmS11lXuEQ9dMbSiUaRLBM1gB72d3v4PbSD5cxSAnny
5dg80qWuORwYp5Ha2zSqYi41MNcXphLDOYAG43QfG53bQV4zTumirho5kaJvHN7TOTyapkAv4z4d
piP9YdqqUmviiE/dS0rvVJZCo1tq9ZxB8T0PzLj0fipcnG9bp6oe7ySt7XMml68tSg1EQk50Do6O
Bm44SeQTBFBg7pXrXnyvno9inb0vLX8v6fjNHWzG6xWv+nu0HrSxvIKQw8OY1NgOF1np7U2pwPDe
2UxaRDePn36FjnZ2t9vn6qTUQGg/Mh1cqzZ4/eWOVe4MlSiJ7IYmi9CXDoU34akAlr9xxHZ/B9AN
qENNqltmxawWyYjcX29MqV3ihbyNa/1CyDj0mL1v02doYlv46TFStGLCDRcIG07CtmybcLNaSMKK
c/SYoLxnzWYatG7rYtT1ww/phmcBzc7c16p3nQHhyyr6LljzJ/A7ywrJnifIe366zyXb6dwyo/bR
49FRBakM2mDNkPiEvzguszpck+vOJ1YyEuQ3Xie6wBAkJUdZ4MlrAtmE400FdelCaZEz9One9/Ee
mnHWTluVsKacC85SMHeYvb0L8nAlZo3kqPoaTRQwAprxYSXJjGR5NwVWJqr7HoDFOj8vHqSLlv3q
Q2TSsbx0iE31n0VlLouZ6mpqNjCWhwLVfMrgxzEWnS/unhCGhifKAc110fH3tnMk7HltEJNu/LxX
2HZrZtdGW5OOKdo5CTCBcAY70RY9Zk/8K6Lb4B0EVYZzboYFEAPtWTv4a3sI6FRu6i258T8sHnTa
RJ6kL4gzl+TYC0Nf4TyhhssQ2DHMzzRD5mmcjG2iQHwjlkc+jtVcJNzDTkSDEhGpwnvVJmA5Z6LK
bwwaz+FZNSt1J5YyuCndwhUyzfA2Ir+sdU/nQB3o1Zm+NZibNsvIp5G9fjew0bcoJjdQVPYGJDHJ
TT3rZRqSYjIP2TSkqF3Wyk4Q2K5Mdl6BjSCCJTFxmFSX+1UE4F1ZIasoEV/Pkj0SW3POVcgPeUT3
V277U0vo4ZxeNJ96q0VbcPf+qTOs1EAWlJf+ZaIhSNmLul5arpMUGbnKsyNz/wRPVl05y1IJcZdX
ox69DZemzinkYd4ds/srg5yRRgshZdhZBVQiujxEwk40BMeqXRUrQt8iLNbn7ZP1thtsMS6B7FpH
pM7M8f/vs/yX1vW5fNYXcxTMjiOFRmNPI4U+KyNqeO0uAHbzjwx6uunLE4j25IeEerXVeg6d3bJy
oN0SL/W1V3YSlM4ho8CW0dn3rvuLSF1Ye6YnpLEUMtLrD6sxBbDX/E1oiw2R/PPz+khKsRvllGCa
jEOXQTqrvIBc7J4f+neRX6UV5gFz74bPR5c037EQiFyVRaXyjToDYK+wEnWRbJT0sMYcCydhaQHb
9wVUbzZd8/WZztC+rh8exHxJchqNiRbVNgEOAcpBdRJsI32XQjlLAmOKgIdqbaDWoz+H0n2HvXKD
Jo0cmQK06LFcG4ZTmOsSH1OkQQjk8eTqeQxLyvoJSPLvklt+2w6HcRe7wiHIE2j2jtBnxjw7b7B+
TGf9Pb7PVv5QQqbC8moHb7IRNjHXmYJ/YRyW7lvYDPRzms+Zgnv95Ei7S+BkwoUy+ltfJYS4mzQ9
NDmnkk1Jw/WtCS7V2Xu7JYVd8ic7g2ke/rUOsKUcp9t67et3iEku4UBIH6WkCIB6tUBcJNdoMEhY
Nu0Hs9jBQa408DpF5s8w7wtQKLA2slzPvTKScv2qTrC5sVzbwG/8CHqLyqk2jpKp2bEuu8hyR2dg
pHC7UCrRedkNqYES6glY4XM00Gjyh5FvyDY4/zphsJvmwpU6NbXjkHhTR+m3rAShZ+hK2Ch0SkB+
69W9rgdHAJQjqvEiFHO8+XZHTpHBk2TuKJo8MyJufshJbgzqN3iE9luLdIvDMzOn+X667q7O/I1K
ixTI1OFLYXo1OOnCibjEVw15erqLw5OndQ2bZ8cMjgDJFFlv0pOtEUW5jhxO5542CrCMSgkDFJVB
thg7THGvvEkJZAifLglNsH2F+w/zeaWUF5VqdkqI/60LiKg9g/yhlQhQYP3G+qLfG2iV0GpRRx7T
Ah4UCqVBy1hpN4kgtMJ6rZ4/3PW/EVJU4mWFe52erZQUGt1ygjt26SENQNGCrWfHJuGseRcbqnYd
bpwqj87PWoHpO/lqeXkiJ2hG++GbghmO5R3WJdDf1aDpZa7vwAHd2/J6i95K8A4q8gCV7/iusl3N
tsUPpbMFkpvw6jzU518oUzxrKK9yeLnntcMeq6sPLdsFsyFhpeJSJWbcdpkn24Kt6tAbbeHN3tiW
eZL9iF8IWCBow/TAWFyq8Q5JsQ3AR/Kmzw+W80hBAsoDEuoTyOIg9NTRsDv4IX4bpQqAp08d4EDR
6ydoCLaeTo/wjgk1ps7idTJaZPVJDYAPCgBh++1dGgR5jdbL3AewZS4KJ2COo7JD+n5vhkKdQ8Ok
Q2KoWrLZYd+tw6i0CDgH7O5PoIfAg/BgBTET5dt/OYJYqxB1lIuAMLn7QYnJKIcx6Ib382FjgJIp
Lqx8QF58x82Mw0qZch4o86CVwBtDVCB7WA1djKK0O6UAJO5YwQzkkx1s4EfT6H2faU/yb2puQh4H
C7g0L+xJJsLcJ19EnMnArtcrVCK9jeX+smHaWRqXxccITBA+azuq0BbaqVIziiUq5YgjhtIvTiH3
AzWzH2T6bn4OFYOlyMmsMdm1MgRJW9k16U1D1S+HDaGPnyGB/R+ZCruswuUqzdMzSO4sTUIsu8+g
lZ35H7I5CRKuCTYtAz3kpcVgM27qtTuF+PLOhh809Cx/mWyNcr7SadjAJ3ifyIuG/0Tp2JkB08V4
QKw9hO4DSa9gaxmweWhtffnfUOxuXmWeZIQlY0ZKLEL0fLohkQ2YomxhID1DerOiO3afLv1v/wI+
ecHynbGvz37dW9CfAxIg6dL6VBJOUJO7qQJb+zmhkZWcnSFftCKPX/xnthoIoiWioZuDP1VXlmEG
Df4JDoeuNM9d2Kwe2Xn2NQusp3djWFwAHZayXW9tlCEStsvtLwjHdh76MmaYAU1VJke4lXU+nn+b
uk2keyL+zMU87o2gpw8cLAyCh2HStnk/+7VaCgcUABpDFaP0Jxfw9HVmN2F2Fgx1e4Ja6kh3DO3n
snIN2SLRwKOK5I3+pAbi6h0I+dbzOmYLJelN/cTnwCn6rW3aWxkeGfhZW05jZW3Tlw2yCT1LPw/g
ZjWtCQftCCn1UXgSosNdHYbcAX4M9QQD9+8EoLrkJFMTIaCRajVPAMXHZRI+BnkLjq6ZCTDwvmRC
9brn7WZYdXkoO0Vb37UvK1hBaVqFO0Mi4r/JAex/Nw7tRwroN8GwN6cbMaLxPlq0dbTNPKOQ3PXJ
A3mUhgDSr67UZSUe11X+Erx/fljvHvFS0c/6JyyYkmEVXa7rx7K9nokRx1jNUZfhITYoyV6Bmqj7
WG4NVLwmmfS6ZVFTc4JrCuj8SG742BEeOhB5sv0Vx1VpzgYXCI/6GtUgJdp4Gk1rCc0lrcV4aLQe
g5V+yENLhFME/QjHyOBf3tmT//TfbQVoH/h1yhuTMklESdAFC0jJlptmZtyEbKHdN/6sxpwuJMjs
NxMalBwwh3QUZ5uo66avLG+HMCpRcLENW8MbYxWMRGe63mIqPXq+CWgAbeD9Rgd/a3NV+51/FPgB
mzr7auhzF5VmPjf4l2hdgXAcspQSLKPsq+cjRuwwiebfMa/D/VL8LL1Mbu69UpPaQe4/qz2EyEpx
AgP3cL0PTs95wDyKUoqVk5LZMgty7qrnEacT3VrvGb6cSZqM85EXZ5x8e/6o0A8bwKPbVjtMDkYD
vAKoUhFaHSXwJlleoGg2qP+f4LOHuKl8HiiBbMpKfQunf/CYG0qw8YjPpTNqjYSLc3ZbIy5HgULG
Hjw2/ruvqZC5mjbDCh2fQIV9QFY+ZWcsT6G1Fm+B0QfJUNhE/tmiMfX50+wOqUVZTXvQy0ZWMl4t
vRHxiAwEQ/+oFlq2bLMpktMZB2mwZ+9BUK1OnWQPiXeEg0vvBze1B6wa3WFOXz67yYq0LmsPcJCI
/sciNENNQxpqlmdxJQc0OUtkJfmTBe7Pod5sNZaDY7GMcGB2a2Yty6ZjfBYBLEzPE0fnNHTYGqgG
GQAJTdziGbLugltt6tciREuGBRUQ1H09sfOJwRM93NIEsBdUqdtixE5ucTAiL0mBvnvbypNhJ/gA
Aa3302z5eEtmKl6XkWNq1/jEx8pGXxdAPoA1roJSR20ePrP+GmuazcndHAaMYkM+YcedYjCAEOkq
Q9XydVw38A2n+z+AsnmVJ/TWRpNPXvPsef5yq8suDYIAY+2AnwJXBVOnFxulNNHCXkAaCNmigmYk
oujx2FP+A2EumWzWmlbCiKolgz70QbLNJdHJzv4g0v6sm4KLaPIztR3N8XuTzVlmJ+wKMCy7v8Fc
UcBkheXTLVTk9MZYSKQVzivPzEQLHNC72jnJRHYBoNg4z48Ca2Tpv8OBNvSw3PBsJd9koWfKc9kj
a/L8axQAFqSIMZb4/sw25CgHIlkJpgYCAPeZthT6rRMYFhrZu7axa3JhGW9yUmDoBDUmXtOSlsmC
GK4UImovs0SHQoexBCMLtaXl7KDpKO3U6VCLwWwkM9GNFSvNUvmfzu6xQafLOpuFWfhouTkH/zMV
r5P6zxGnbQY4K7y91omR3Imts1ftL4lxAG5cTVsG9x5Gi//MUVnM+w6kX5K4hp5x3lbw8uoMLZUc
hiT4R5T+K77T8+HVXQpbBYqSOFJkgUUdGvJPcL382YQLoW5hS/cgGzgXJZjH3hgyI+JcubOeDu+H
U8dy9xrSIFpXAdzFlcxluPK6tPUZsMzb8nYBgY4bR2beD0C0lSEGDnCwlNr00IOAr4zu7hkmPoA8
3TZobKaFZbg4CuJPiOzFewTaUZpfb2wXd/Thi25ZOSKaYwm2brio2Dfa9ImxvEN37F/twcI/cXW0
nXxbJ1c0VTyW1sU71HpUZIH5wHD00cp7UcTn71ys46XHyYPHQ2d61WhjDIEsphSeyYdtnrxXiUvJ
z74o0juzDtdglzrrEQSmLQkpmYopSC874SAvpnqulQztVLyUB3PXSwVCBrfYI0bEuD5hJB7ukKJo
Omn34vmc+jk6gENjmogvE6hR1c0XOyU1CUITp+pt7ksB7zFmpMbWIR6CiEIG0BOU/Cc5aPHlIDxs
Yx7JOIsHwtX5mQ077jtdlQJASGif3rxs4vX4Z64dKm9vVUDkXy7IrQp2wtIh1+IXRizbjp+m0KZS
BYikxHYtzFNq+8dpLJ1lmxLug3UD1VHjR4FdWGgqK+S8dpaL1pAq9NEjBIdHY8k09pRb84Nib8ay
2iZcMbadU7nD+Wu+jXokjzhgDspQO1alo99z4OEUICA1b25TPJuYlbIVINsnO0dxTCH8jDxh9jbq
wUZXJB7nQRi8x1FALwjwPrd8oK13FkqDFoD8Q33cL/XlEeE1HDy7hwxfmGUCGuA8cMcdknKYA7s4
5ODYE3Q1a5e6VTambdKVWci2aTQIDGHuVhlmafNAJzoMy9OnI0qKJBFNkFTUcntql6RxV2AuELf4
oQpErQg0SDUrlk/2G65q32RKMpGtTDpfY/6I8G1oxpRfJDSXA7856zhUF5DvrATZnhesasfHGtUs
4AKVeIaOAAIhTzkB187o5ASw2KylkTOSXQcPGYvnu/ni0osfM4hznTA+vpqi9TmYnU8qRgb70yfV
ouAPZenCfcPGDP+duKq4DvUH+SOOOR8ll7Hz5I37R0aS7MO0rrF9DhAmLcVVwrATvJX07wxrEqVP
o9f0bTGo3IsiIY+c1ARVb3wfQmVlpJMx3OR+2PSz59/XNYgHTtJ86b4jnwcWGQTEhrFStL4HuKrt
VNjAZ5iTzxkMmmRuZPhdtnWf1BBCwy/wf4ughJqV/feZ3FAJnW/XXqtTPSLw3zyWRguJl30wD5Ky
OkIB5kELMEJhBtKlD9w5abkp4O0swLjatYguIa2e+5ldHLgeP9AJm5iPZVFXbyTkrlUTKJYu8fdv
5QI+sdxP5aghM7Pn8p4YHjy58fE9daCmur1SRQQQ1bULFslXjRK0tR/SKmwIKtbC79IDYJ1Ts5+p
Yy9d6XjC8VrY1hCuyte2+3oIx8zgK4mxQN+5dH1f8Nv1TXLJjSe4NrUIZQcj5+XyAqsVCKSjVADC
K/P+LLJU9Fwz+m61H4nUFqfS90d9uuT5/Fu2gPcvRik/LuH/+wM4XD+kq/zSBlCrFlf3WhiBBu61
4Z/OA/FBBWyeS0jgGYqaDc+4uR7OSuqkZ4CxGhvaAeDpxqiG4vPjPFiMrvrLSDYGVULtRuUxzN0L
blbFI2D14ZjJC0d/aY38qfU2JJS6oQxvH1RjMhOCkGU7rYim/aTZA0JL8H//AkgCTjQ3y87T2lP2
O6Zr2QzcdQjwdSb1sr4IvRlds/vnew3fKPlQ9yXc9WelN8hE5Naj5/pHND4oH+mdS5iWbe+c+Wl6
4SWRj55w8lbjqDQDSRnw89LTYfs4Y2D0G2s+xK4J4ffF/PtWzHwzsYqKKRHBu78DQj1KPwyT0flA
/bYFyYxb8NhjGloZpcUtiYENHc8IV5Ee/zHvkMXaZ5ZDfyQSe+V2b7ElbTJASEDYkV1uvUaVR7xR
UmK+dnnNCMDo6++VLah2BWw1Pzb+q/GEslj+P/RAovi5z3T6Lza3D91gbuCkRyUpmj+cYVIYWkkV
YxprNqGUVD426keiF+lHU7/36wLS5jQbPPRZr9xHuKyaM1CZuu6d2qVgKiujcxIkd6zzdrmbtTw3
0iYPlcE7fqZTqZtkPRR2hGbFTcJNTEf+OwXpDPYfWTWVhEs90aIe94vmXFhgE7ot2+Nz+tdAZ1P7
YPrp89uh1/3C98O2LJ4U9FEV/aPqkeq1tkWc4VdGC0pnLzKNo//oIP2oK65hAmR/rSJsHBX/W5o1
zD2J+f8iqLbWcbqnWGgyWh6R9uBiMPB6QQbIYcXJslDXBFhDzbsAmHUbKlPTuNMVZLTn8w1UIE3X
Rpk/WMUCiHe0JWeByIGvVjrqGheB0aaDvvY0H5SlTU5iXdFqWvfhOJwiIv+osUvsSH+ajOw7LO1z
yyCT6CTcvUo8igMaLtHSGJXMz/I1EyiHMQbORIfKCYoyXVa9+KcfvLobmK/VW6yw4KFgm3ATjv5S
p7QPUUPaBeaVXv5vBsW9QSed9caDt0N1/bnkcrKr+JJxYzWRyuceTMddUGBM2fUqES34G02xs4dD
+U+F8JfS2f5bWSr0b+56qSl8HWAYt3FiW/vHEPLtSvhWegr8/mMSghLQZwe60ibkrCmCqrbo7x1V
fhnn/V3un7PRa+LjyWSf3fgE8AxyaaNG5MQZfdHw/bbn0h8v05bkZsMfd3s83gH8JRVt2mGE1vTX
Y88elp7BwxQ8HQ8Lyn7pbwsyEwcSiu1JtxAHHARN8mXfViHjEIPZ95VbO8wvUavGglCUmil0XOSf
9U/3EvWetYaH6OxsALaGzrzWxw/KNy8qBeLaAlAPLWk4QF6bkQM++xhvC8/jWGi1gX9+1Kw4pnUT
NmufIzpZLueGWTvVuC6yLV/OO8jJDoTjFOIw1jTBxPAFqF9o5auf+vNPBSBNHmywYX+cqx51ga8J
2Djjblk2ATRXADZeCeT65nkrXNjeqIC7TAkXY86eFZNOj/di72rhtC0vwKnILEk05eY+yOjnTAps
gDezgJP3YUZUDZ8Lwb3RT79h4z+vxDwkjtQkEnglsE+4zYbgVOil+6bnbHgQyyBL6EI6eITIhSdm
/cRkJDfSseSwWWlz2I55Wo8QRfgllva2sy89sVsu4JnSastkNFPxQYGDqZEMAI3RykNsYZWHwbrI
lNxCVNUBFcOxfphrBkNKrglYE2mjHvK1PWEpuMTw59/UXRgQ33fwVq0bKzoE3xmApZNsU+HNlThj
whqm3WDi+Cnr4aYGSi/FGn0JmUvS3k2lv63cJd/ITHb8YzbULXkN4dp0V1JrV8opCBkn3Jl/iIv1
Tl5M246wz8yIMvpis3d1rz5sWxEEPwxyf8qzDTY8eRzH45KuiC0LOaO0qWfwVcPvoRHB1IzVibNI
M37WZF9t961qaxJovvEWpC5JBvNSszgtyW67qGRFXIP0bWLo9Ymit0RyNtTnY3W8YWieAO99vssM
eK3K8exsdzshwSAdoEgxz3FPycOt6z75mfceSjKtraKcudy8V/rMsHg7J1dKD//HJ1RKEaYlCuC9
73NEkTNNlpnQck46nIsSbk1Pne+RzeYhiKliKHQZwgOXrvSqSIGvedYD0/WkinN8j6Uf5/MT1Rx0
5LM448UutFwIyKycMLc07cZQbEH2idr+fPy/QBg5gJRWxp8zA/3lCOvwIHCLfYyTVmozzFQ/PzaC
qJOhN5oTUNd8/2JNsPrV2wPSEd0dogoLxkhvBeJKCuDm4JM81LDgf2Q1vSSKcUgKAs2jF+RT885q
NgEphwQYm5c+SSi/GXEk/TtZVAJdDcZpj9zPVpQx+lTySEcWGCtPIYMh0JhQrI72WjlmKql9eilZ
ruQiPioJW1xuCy0cK5lH8dWMJ5DXEixyUIgJs2go/HLqSNuZBdpKL1/J0N4HqQGfbzHcJIj/4l9r
BaODOE+2AIF53ugexEBstrrc1KwUZgIbf2XQap/+8YJoqmXTlygdoTUCla3Y6Za5B/eipFIaCklV
w3q5sxjtjaWoxSz5sxCQ7GKd7SDV2/1FwhJsvvT+TgmC0vVkMcLCbXiFjv9jw/9s9jhlSAw6EKxj
QnpqXdKRo+iwGLm7tdYPP97hqaYSWgiEmNSyX5VkIXg8J7bp0sW+RTPmSBcyDncfMu3uXJ/sYH/A
gQTwpPJpHnKhibeD45Wh2wuDT7dXQah/v9B0bKCzC4+Vm8GzMXYu13LSJ81mn3Lrtwz+9tzFcgNs
FbwI1xccDEiuXKa8bWEGC9r4rFx9711ej4k2mU2pW/5qUzHDEtIy2uMWTp6ze3AZKZROKzEnZIY3
47+XejiaWL3+KQFcUCm8cEukv3i/GgPhTTQ+DlaRHFuXm3B7uaEbyE47PzPVrtG1wwc0jdFslhjo
hzK/mrcgnczNxos/jn63ZllHwzTJqTYL9FZ4o2k/pw+wEZps/XUzN6RCPZNYNerhwZGGu8jfKbh4
5pbCSGkWpxZwBmOkwsS3oOrMsz5byZa3pGys0Zgmn/lBcxtU0RsfqZCsT/MDffEngmkIOyGCT63K
TzDgncw03oexNtbnBZ84c78to0fLat88EsTDsFI2N5FOGCtvhZz1gn9Cn7etTeZGCWmkwR+nzVW7
9n3Sd4AIRpnDU1UiGvJ5VJlkxz7pfvGaT4ICKukvIoDeG1S1WgTukZrOF0kfTEGwrTy1aHBhuXce
DkpoyDHTQ9uOs8inqq9iEmwR9xrQMyQdiqSCKOKvG0MopcL2cxLHO/zJs1eGVdodO5P8NmxpfX1n
F/bbSpb4D7L1BkJ50XZsd1vgUZSJBaU7J6dNHwYZAaCHdIDgjhUBe8RvlUbKRvJC5Uvh1gYglHxo
LuZ+2w3XOBgck5LvZ6sE2FO2DYWA3G4oMV4PhiI7V34ZmLEhmkPtYsjWb/LABFF6P8och7eaLs1P
rRdi2OdBXxiy9Ps/d+Rt3scfOoDiMaTonO6HjLFMAMBMY2pehSkLtWfWsa0s5Nf0qvaPGVeF/oFV
dtf31rmRLT057u+bX7SgbhCf3R8Ufk3rKnvnIOwYIRRkiIzGTQh0MsPNxh+6b4kCbLDesF7HVosE
O8Z3ZzoBShTzN25YClMYnqzGEoq7vuClpr2MmOafTZi992388ETff1thaaj61giqpDIDFvtFK5W5
H4iMXK6dS2IF/JWX6i/8A6VAbmXBtuxi4XiBvORskWjvp4EylqS/Nh3OppmK2gNQFeu4JuD/PgKP
ylFDWucRsOHZT83bCRx1icAzZ1WXp+ANpON/Z7k/EKj3m7kfryZK/9KRy/RbVTyEQJdVenwVcc6T
5jAKXwWlJPEoLwa+kfSk84+b19xRbU+fYgbxE2LxyDU08+xk5AuO9rt+YfbGB5oIgGquQa3OxVra
sd+71X+47c+QGiS+31oB1meNwJr4AI8qEDg6/AFiFz/aSmoWyQUcWjgxvtJqHvpPZjaLGnjxB7kY
eBaXd55w1pSuP8jgM15e7EAAQvxrltmKgYuvq56KSms43jmePgO4rjwutCdlRqqPtEKZfilZ9KzY
/OnpJ2uYnqpBY4801FYMG4XSqKJuQEqyCOjFNMPNDIhPBjregX1+bOtUXL8VyooHXnmSC2cHX/XE
UrUwOmkBxOvIEhL+FTNdU8flvEUjed9ZmnkX23qie8kkSjIA8IhM7yIetLZv3edaL4u2LHUpgxF8
gL3Kdacr3lBFbDjBux7ZR5yd5p1Ot5bjjYXWV/iss/086AwjVfO1BEQxP/9WWlCj4Ak+A0pmuQeQ
dxoxqXa8QafovaW6MTAa9oUgWncz723Rot+4hHMbVuC17SqW7JJZjV1ImlDTDzmzN9gkmEDu7Dh8
/y3ctgHj7+H0QvPMt8kdKQApI/koylu6RWP6a8+HybUbQaSr2U4dd3RglkGKSaprZKz/ETvUIL+u
2rmNnZn0Cf9og3+ZlHVB6L4n0UPUL7w7rFP+xC2NOA2H8hbBGnQLuBfDEQVtqTKaS8Hb+4gQHSDz
oL5c6hW0YozbVKEMA5UIOESeNoQO9UxcMY9w3lWND1jB9LLjKk/fgiKH3YW8parUaN50IZzCuk0a
V9Rx5WzXH2aHdgYsfDtMRMvvDpr0qfrJzDXm9iNOtfuJJb6f3F5bl3RGq1tH4I5Glr1/LqoMuCow
S+Q00CdS60cd4W5YetwwmGh71ZiLj7jw98215BXwUWExrn4zttoVQMphnRnIiLNjlUiaycJMSJ63
7ghloPZlpADSnGHMvItlhJ3BCRGcK92q4o0eo7KagMihi6f1qr8mHwIs2oONN3Td72xeibIZ5gZq
BIQrDgMjypb50zet5wNx/nSdAJqSHfSK7Ewuy1iNpKHxliOfm1fwG3EiL2fSmcTslX5oH0MQIj0c
j3QUpY/eSJMjaFL9hGSsRZE78ZMR8cZNy1yjiPjms2c00l2fevY8tvCBNNwFWhJVcz46K6RfcEoG
yCxUt9FNJXXQws26MfJHNy84IHuDfsrmqTH0/fl6lLNJcKAkTp8N2ti9dfeESsFDTSX9bMSLndQD
+dO4TFFsaSm/3vZqulrWyPkI8bY/5n3olGHKuV+AXM981leSz/iyCW97cEzvSlLf/2nmgI7Adark
cRoQ6voLvScVmoRdjQWRvGqw5ke1RODyiIBa7CU5OsymYzOSKmecSKffxGLfzZb7vD93vwaroQY1
B8DHIz26MDw33gbyn9us+fF2rMMyS36ZgSxYwGOCglQ1h5mwzkFRcIbZkP5HRRuGdGRjDOGqzeNx
NQbGQo0FRZQDUJULbhibNn2SBxS1aXIkmMeLQIqUa6EsAS3AA/vmvmMi86fv7fIltNQDh9RrZFc7
dwqpWD+RHAESOYk4eiC4j0swCjQvFLqYks4Ch+VfgcfigS/006m85Rtx+fBQI/A1dGTvMeYORw4M
hLLBGCpX3G/CpV/lphEc27/sXT5glBEOkyyONL5ECV5TAPs+1oHkgL+0wmxfoZd2VQwuMcynOAa1
no8WqqGBAwubctR6J2nMVwcxw3k2VvPTTzgGwiX5kistC+/OJUZkc8mB5pWNVnVUpAmuE+p6WBZw
pPKa09l11YcYV/vAtzhIMv42FZI/fnLgC0l2fKT8aA3WUPCxgLPu/Rjdkt9CEF3TMTFgVNV/DQCe
CTcvPSc9hKSz1O3QsKlEcxDnuSu2JfOiu+JHybi5pwrFQjJjw6VEwatn+pO3uPKH3sVWWgBqFl+z
Gz2PQLZc4eySNsAcfTq+I9j6GaCO5Vk3lAYDfCMV2OfxctjR8cqYi8igpFXY+YIaLGkik5x4EQxe
IxnoExWLAxzCmbetX9JxsOEEdLaIFyOgVCdxySSfKji0/Lkl9PI4VP/+Y5BLLuye7deHbKZRJTkN
q58iuTb6zwDlFDJl0y0fah7AVf/rNW92Grgnzt6Ddp3IloCV2aLTHuAYUZheFN2y0nNP7a8wWuzV
YHDKcRUblxTaqG+S1PAbNGnvsp5drVRkMnDmMe+PTSezcQJsakzMmkhCH9T/6Tj4Fa2CmXXfn2xx
Y48WYompSeIfrJsH8TIG8PMbkghLpFJ76uFjPzX0lVYtrw4Sa2QFScUJu1nq0Jv4OF+4Q4p/W+bY
Od+CluheRv+1Qj4GNKhbf3FkFrw+BAS0GmSRT8IQhFZ7MzbAGTPg1EH0YqtCKVdu719hVgYQdU3G
goop2ClG9JJQ5+UBDSBetjtPSDJe6dJY1KZWzQ475gQksKFK1JgHB7/f0yOO0vtQBIWNp21RLVGV
G9wNxvlwmHxymEzCXOVJk8x6mFGX/HgPBvzrWb7R6k0SsAPJB9aaJAG+oSNpvQoF84IOI0daO0VT
AcJjk7VigrHPS/Qz8I1EN0U3nXJOtF87o/C/Kzr3SskJYryaLGS7jhi2L7Z/HcOx+bBjOo21CvT7
xHw6jnhMkwm5s54FQwp2hcQWfrYTyVWXRY1WVy9GyABympiOnMQJXpde9X9nFLUISyUmRqt/w0vD
Cec/DZ2ZzIxpnNwhhO4IknNjy6uV2KV4ng722EmivPtDpkzXt1kQh+56iOeAyiULsMtZXCuWVXkd
gVB4iwJ6ZDYIY4eCK6wBztEDpY/qpCZvQz7eMr2VpNMVNHWoP/mKpNIqCYeAuIxcECZnjRvCV8yc
hdWyNsotbiHimTGmaUXpwr+BMCyEK3Tj5dpODdAiKnzddIH863Ph1UIgCx1Y/bxVgzHouKxnYS2Z
hPR9z96ddDve7iFnn2Ww061rN0oM6uEKyNN6EWGZjwnbsoyIBVxwr+wTb/X3NuNXbm9OdKgKISEa
fZiCG2qp3HpaBjEOCRqQhkROLXE7dFk+T7SJd2yMRylxSw5+30JxJasCuAg3G55/nw9iXAhTLSd4
0plK9UEIY+xcVVfkrmVdVdyArwvmj4pzsfISlbFfqTnWcfarE377Secb0Os0UC1AhAU9dVZ81hS8
fXPG17ECPxGTtBQIVxcZO1ysXvHR+rpQzxPHQ72jBekvpsZNBTyZL25aeWFdAkk6/RZi2RjQG87g
+fDKsxYAdnaTCtsNnhpxSgEhNgitEQDt1wXy21kjnVzS4IJ8k0Df392CSX8TxcVjUHKLboZwtbDF
x7iwD5IP/vum6O30xY01vaXYdtjQ+UvKlIsENhfKFvVFcXAqc+EsvqYNpNa0eyrvBsYrTYqvQPka
LRvi17nW3jvFce8RQ7vbFrEDWpv/NwI9UlUES79ELVtJ2ew4qDjrV5xxDrzM3zrgoXuHuQzWd8w7
0dR4NQ1OVkKXiha38PLOVLrg7ToOI0plbgpo66EwXpY7XhxhvcWJuSQJLjcCsn+/CU1xMn3RMcas
zU4traL8+Ca3ooWE7K2FNsoehb2LOMRpHSrAgEbG/eosUWFK0o2PF8wSGnHwpmjULKFEnQGla/cY
rYKsGFZCaaPAWk9CNvUA43X9FZ25ye8mXC4P/lMPS4DQ02wMUwgS2dbPbKy/vRypjo6CxYe68+6m
DSbVruln3ja3VagsqnMQivNr4LPRjw4kCisgEA+3TjPBl/XPRdMQtMhigBj0ZN1I5o9p36vVMq01
UlLq9m3qC602UQ284Q4RUmYnYlI+3kE/1JEsxjWDdpqlqmaxmPKVdGopPAtJDV+LCEIcuu7c5ma2
Kg4Ni1VNWNQwZVPOVPS/1MBPTpTMZeWv7EDiNQP5AHgeZtvqTdDQScwr2CZZTOKwri8udd2Q1ZKE
5N5JGAa+3fCPnWo9IebE+RVgfnDPB2rhwYrJu47/bPd5A/TPI5tPSG6ybeFyFXbSxp6Pad/liO6R
h48sSWjaIpkUKfnwl/uaukA8X7Y2/NH+yTzbFne+v5b9/q6qmVK7vVWx4i2MZ+2BtKwXuN2baQYM
s1ZKCDXwNgyLkz1eGvIjxz4B/Yf2nh5iWz/6iJSwN9sbexcj0fXkSS649FdRA4B10xExzVk9eIDi
oarX/RW4p2teL0lyuvq4uLJoYxYXwoIzpjWK2V2zlPkOT8z+tOkSK1oEOjRBVLuQQS2aXcYQrO1W
Xc3lanPfcmGKV7JpXHHMGcTNs4zOA/bixFPUCNUT1f2ftGcfi9tAaVxndaplG0lMWdXz13Unpf1A
meOZZGJIahhtJqZE1CrGq1azub/4SbgAC2ziHJqOqxzuviiJeQ+UMFuENMMyQy/uCTDD/D9GmOTU
r0LqqNjMHnbdLZrk2Az4MmZDH/GsDrSrYUYVf55R1anRY6Ypyrxm7J4y8tSmlo4gnyj3R/6Hb6M1
Ulc/60W4yGlInBFX+4fDkfWzg3chHRVcRElUcj+UDhCHtwaB5V8Kh8pxb18Z5PLcQeT9RsZFpqqW
Otg5PxyCB+jhkVlN/pppcDdep+uNHlTgmAi54sodNtufpbutCplJu0ThzG6xkY7mBrHroCVo76Pz
foDoeOC/PgLe6eCSYaBdFxg9OXrVdcYsUVW//O/TQtCO0VlDeretwpSifzqNql1Kg3iheW6VTmBJ
sbUhfa4XIhtxk6peaunpFRM/oHwXLuVftGwsrJvfIsRJfk5th5BCC52Fu+OkCf94WJvM6rwcf0Zr
/JtgEcUrauyQlF4D1KuepSWNK/mNGGLvrgnez+QyTT/BTCmWGbLZsOct+5q6ugIP45XylOO9jwtk
uyKYAJWtSipeTygHPn5JdlmQNRCbuG4nm0i0OefHtzKwqKpwlOGe+lxQyd7rIHuMtAkdZYQ1B26N
6KywPh+UEgmKib6JIijRtI4YsrNmtJUK3fdPuE95CP3fKn/aHXK1/TqwYYVrNGdBzrq0hkCt5UVu
fKQMx3oK7EXp2ao+pOzjeXK0GNrKcJ+QPuZj/EArG2zopziwmj243jst3AsOJO9THkukz2HrvSwf
pKgLFEN4bBE3DD/VnW021SX2Il9IwYYotAsBvicw0AoEmgNF4VHDO7aic5UxeYa3YP80uG1KsTvC
ZpzySZ0Xd30rF1bl1c1obMLqsWspDmuj9cm72JOMNUL7leJubNckLUx//vmd4DKocNPCuLPPfuJh
rLBSqYv49npSzq2ZIcx6EoiFlBnX2q3ffnYgnI40LUgVe9A9R4CzIwiwrTY1OSYCCgLIh1w+dgZp
lGz5QOp+2OFIyB8k8dt/n9MbYR3M4pBFVtDnxwik+L1Fc7G4UxNuqHi9NuZ6LbULEFy0cHFa1Zyx
QPDV8EAGEDsytah76OeBTdfmflgAYtAzP8rLf1htdcjxXhbTqHAVr+35eNQP+nN6O8KVOAh8oHmv
/c9TfGF5BErdEwqwcDqUMFrMuKwCITpP0OPt6OBf/p0T1bUohbIPzvoEjkP20R5tQaCOiF2/x9PP
rJRml28RAhdDbFH+TmtW1RwlLUAjEtJPn1zMMCMGkg7bcGEY/sjq6D7XtzuzN6TD/Yn7TQE6jVYt
pju6NAnAkZYWprce9OeVWTWpA3XbBCzp0eAkHTJTkLnNDxYLWlWtc+znrvZT5jGM/tMWWYPw2nm/
Sit3NxGJCEcHDEyscq/ZgpF9ZC17tR73GqcKKeItYNfJdrH59s6nVxzuUTfVrTbCUm6EvBS2Qpf/
qmtkNkvFrTuVq9++Vde9ZweBCXM0YTk7w/sn0+ypRbIA79xNINTEheLIlbzunWFogtjtIUziiRcu
siFw+bQDS2ibhltOBDaHsTDYx41LESszy3Kqo7A+tImWf+4/hMJGkvTHMsRLINuwnOgwzEiy9Qyx
pMdqmRgHQz6thlg4knwp/uxCCXBd6lB7UglgBkdQR7EQecNY3itnnPni27cz8N4FIglCuDe9+Wj2
Kekr9Y6bdRpR4K1vlXiKCiJFso5jaYZMxFeJFG/zq7EcD35qucFG2MyUE7Iyaskp1gE/jqslpnXk
Fb/ffHMqXAjb7rtOJ2zDJmZrbrmFFQwI3W08ADuJ+ytlST0VohJ6siL2XhecXsMKTNd8JivSgRrq
KqxJps7SypoUCFJ/fONCRS/7SpnRnZ4tdLOnG+qKt8bwNKJiQFBP4i8fm0QWqsY6Rk25bRxXvCKN
BhKsWCuqDHmkp3oftZeS0NSqJrhD6O7HEmGNofDBBjFovJPWNfLn8dhlshsrek+t9BG/dwrMVH+E
dc9M6KndXirW24QaijkiGjV5HPZG4iC4LPKZnOQguOjGLxh5RJJAyEO5c+t8E8kBUkACjcQrPHXE
EZVLwcOvnkmKVyyOGb4LO1Z02JJ7/aM0QT98wYMzZk/20roC/v+JXd7M7mnFTbu0jS+ob/95+7ne
lprRPsTLJqR3EbzF7aLmSXW9ymqsPnwZlyK6Yw2hkKt/RBoW3V/wloDnvwzMlJU/kTHi/L3ZSuWy
dsd+1sdIfhxBI1XPirIrTX709v1mP+MkuU7pAOem66C4cmIV08YGXIp8iC7pRCm/jgfa0KTTgSGY
MG/A4muijkt92RsqNcnmy9pvyglsx9XB6Wk8gMtjgmQEYeAnYYRe4UGMcW6GkTi2phoU+WhLtqRG
kImYfjAiop95Wk3q4bEZkdgp7QgtJpPAyRmqbACg/gp1kYFaj6yc6piRzYRrQGoNwVjHS564G8BG
SPR6PSmrS2bNJm1eHCweA5e+wmtN2+UItCbTV/WUmCr8w1A3bUD58mBbWSY+ba0A+5n7uVbLMSTk
r0RzGlWrBKfU8AiRiXAhXnij6cV2sSYOjSdia/jVI9zAKufneSuhOiVZyefLvge2lDM67nrnd+VS
W+NsT7HRW52ClioOPFROjrhDSFtX12zVEJyj0/io0qrVmseQ915lpmuYrL/mvp/4aBQ1PMt38V/M
y4kWXv6FrV9Ta94k1ihfz9z1d8L24lOZaDfihztLYNZhnj9wR4qrvg9ur4cviB67M5IKIz+pGvi5
yWcZtOcAdDAD5LHxuV68oEO3ZF0cGlD5KREohhexZTTi4Pk8wLND/jNwWEUVvvMwv/dOCsFA94es
k0DwoTNStF3nnQmVr3ywKIAxV/s5xKf20SOYLvzmiUBvVrX167Lq6NTyn+5x2dgOfB/AkDvbgcgM
3TPvXMsSVJaPCVRvXTD/PYdzylJMA3BDCfgFaVJ2xxcH64rdmTgOCTDiHUj/VF0dMmFOUuLnuclJ
vcuZslJeZJQJ2tMAolExS2Y99vMk2a/c0k+XslafZwlbzF4+sxvXVNrR8Ez3OlEzWDXrGJIv2L3l
SuMHMhMZLRj2FQHfDvRCW842cQlu1ESOslJOCA9Hrxg08NHykmV+6vngtx+KrW/6GN1qDbhOBvnd
TQCzmxtOPUYHRwWjJPL2scdu4m80JqDb6OchE98CBPaiE6siDc4kUuzFtOXbnsve2+dZ8J1pAZQp
Ije91pKMH8e82RPeRC5IAljNWICwK7z3hVSRCIDeQYrpy6isNWtcrEu2aQvBkpAC4HohiMa9G5Mm
pO/go+y9WsOdwZydYoVwONcCIs+WI6vihULHYQTxvRmf176VSzZFyNsXOzmv9KjXTJR59oGE9S+U
sqYSCA0RHyDFPikU9rHLjsRhySb6H1pLVK2i3TyjRSe0lAoLu27ZkH7tnRNUiHaNNZtk198M1Qri
3JP8E5BksGkuMvEThlFpOmfuPMwzsLEWGOhEml//r6LnIobymYu1T0LlyYpQ879coJIiHK4I4wCW
qXcVyEED2F3hQq0Mxsd1onL9mLHJmN14TTnmvGPKg8Ogg4k0Y4EvXenO5bmiIPd8KDJypD2EpRFb
Vz18J/YctyUX4X4+znGPX7Qg/8qonf6hG2NQJ0qlQGh93Mf/yIlSptohZRW7MY2bf4xeRQL+ms3w
h92F5vDN7bpS0/dO7Wq2cPmi0JnZQRerSjv8IiAEDzy83PweEGVCyZOB71FNIKkSmWLu5gNxH0Ey
MUAKjDiHdgg+7cWnE+Qa9ePXnsXXtLCeT4y6bimGSRo10wH4HiYJxH8S9O5IUNp3niRhPf9mxsfI
i6J/x4xR3HD8lSfD2o5J7EIcVAQxsZYhIdg2s88UfVndIuoHgmOOBJBPn7FncXfmAriz1SW3NsAA
XBpKXQID1tiejCdzzo23x2Tf/TyxVm7Fnpw0ToYEzgodQmo8e+vKWxAvzxWQLmrlVlZzvQ6IHxBv
g+wP5HbwY6HKYgMbcMTHyANK7sYgKyTLNmjc6JiztwvrYzGIoTwC5YBTofx9WLpubI1nHQoLd7Yu
wIxpYUZDcC3csnCtoj0TWh5pp6AIEIvhZvJCwNdeO5gFRctvRK4zwTDRdXsdbKcPfDYYRgtoE/HG
3fjsMbyRTIUv/h4wQ9C1gu3k5y+7aYxsLL9NlifkqRQJ9RcogPXfcHyYBhHMTuegQBn94SYOErJV
MTDiGesY85/sbsfcr2HZDk6Ppq9InSWkl8p4QZFnl73tFaFZRo7Y+5GOm0hsVvJUoAIUd7ZLvWgo
XRyJOfN01RG3t8x10c9rbrlgkJVoHcwp9Pv1CFnyyu+dVf3DSmxhUu41GBnGEKhk7LnIJ0Y58lTd
beJDmnhMAXv+kJAgkKc7NuQPeo5FK0FNZHuYX2BtEXS2+FkFfPuQi46z5AOKrGy19rQ8We+T0HOt
8v2ogzGYmzqPQEkyPMw4MB4PM3TPLYFQyKJBvIO/iWTv1HE4CJgmoa/uI8g4vdjjMGjSAvPaKwci
qn5MXShBr1upy0v+UPOkZ47rdXZzUa9b9+uVmitQDm6w3mx1BVg/J5poZB5t46jM7hxHeT5oBdAQ
LAdxcLjoQ4VergZ9A0EeYGN8eMz0BJrYOPTYzsU3K7EJo3c4JwwIZicHNQKYq4dBRGu1/wm+cGHA
IS9e+cI3pXCxuBDFAbIqgGLWpe30acnyxza88z2GSTDLYQ32GrZFC+tvJ8RxGvc6iF9JTOHzYla7
xmEbPnR/QxsKguMoUkKD8MO5djoSO6TWBO7xSUvlUDpMSS3WUrkcUGXF1Rkp0KfSMNZ6cvAc+hq+
k1R9WeDmfP7HLuDJRZuZD2Wf0gAlClheHL4i7zdBI/upfQWF8XrBs7FnEAbzODVBlb7GKIp3Q47J
SWrsqrTqOH7OlshltQ2y5cGIf9ZIO6KyLFJ4o6U3aLY/2ZABzBk+WBLE1h25PlhW1pXHFzDEEMbn
naBBxwcXV/s5Kv5qbVq+9gpEwAaffmd1ngdjF1q/ka9JyBUvPY0AEyZkxHB6lw5m0NTkDBAVGAhh
aEp+mOt7kOZy5rVHAFC7ehNHpftbj0OBB0teS7K/LNYlN4GGed08SeOhvWDQnRglXK67Ih90N68P
9+LPNVc03Zyltq8iIg7et4Immi0uQQddwihacF4S9F6+sqrncHUk4oSpeebxI7qjtTrvKyC5Nb6j
SoI09Z5ainreR64UGzaW5DVyfJeUMhvGthh3ydXTEvv7wAGFAgLXeRw5+T4vpuRjkjk/Cg/4T5b3
SfJRRkoq/qtaUEGGHMrULb11exVqBeEpL7yrTr90Ul1619hnumU8EYdSOdSS6ZpaXku9mmJdBh5Z
uNFPK58c4qaeCL2RK4GO7W5pMAXgPoFQd2z1vZ5WTWllF0+eK2t+b35sBC7MKGqC8F9LI+CuOHXb
xonpeFw10eZ5BwBcPes51GHlPa2pOEnKTQHUpv+nvrKoE9qRy40VHcdzI/5fslXt1XJGRhVSHhE+
8mnkxMS2N+k28p4JmyuR1xIKAl/mWIxclFjnoAk2dweeHqINAwdHvhDzqZezK8p7mt+G6oa+ag+t
yM7CXdf+x8BL99YnF8Gg53dtjxiSlBHst6wsjhf33Ej+buXMosVSdxrU2W/xZHPmbQPPTXgGfugp
Og1CesY/w0IdxWye92/Q1aOED9eG3jRU2zx/0WN7Oefo2kyEQgFL8Wj7flowWCbzit/oeBiIMHRM
m/dIq+YJx1VyZOoqaJaWjieBtOg0Aq1tsUDVHk2eL8Udb0lqDMIx16apal0kTyBnAonShO9WahFk
7GODZO4tYS3GPh9QDGu90/kMq3sVVMvXCCrfBXw4JzHaWp4LYh+nLRrCPpSq5t3Iz4MOVROudHuL
4DsjYN4DKIifiMUgqLSmuOxW1iMKzxBqlYJWOhK1XuqXVxmud2KKJZAjNG3D1r4cs6M6MwEEttxe
/rP6fCP1Ojs9CYNgmvRWEEJno0NH3E+6KnfdQoG2Ti9kNPUrGruGoElO5BtKmlEmMrpSLQYjfnj6
Rp9tKqh8GUbKxfjvq2dq4mfOjtcMxusQWVBXo+sqHlMYOs9d8DaQVhD/S+au6L9EvidLSMhdKpa5
pElVrKqkmFXMd8l64SqmV5UFRUGTKmXQgmKbzb8JCQ3i/O62DmldYlun1gSj3n3gpA6KMetwrkAo
X995uL7KI4Bf/HgbV+wQGGg4XSI3G4wWnmOnr5x9mSyVaTsOi8LjOOUIiiNYxs2fTES992qD89vI
7XbhvTcu4b2YV9t2PqVZrqnz+d5gIUpIAKo0wz9Og+o256SISLaxI+ffQS/JxulWV8BRS2BWMcdL
3CFAtY5FW1bktuuJfS5pCNNzQR3GIGZLNGGVA2C9WzprMwJN/tQvWNwWk0wZpYVX2CPLa458avic
K6DlBmHNwhH/M/343ig4sNtXNvB6xXhclHQZWWaTLxLUssnRyAKxT6JHYy34ZBqv/LzRgJG1PfU3
IB/kRH7Alo10e8x9s7timT50qqlT+rRbPaMgl/BDvu+rJqmlf8wc2WDdrtMb+OXJh3775tBbdmIU
LfwjcB/XlrtMOLioSRVmTWU15el6m0VW2yuSFm5U6rUFgmKcenh/Gt7JZe/Wums0sa5RsA8A933g
dbUuRsE6U3acWKGLuWFv/T6jUMsh6D3B/zez5cv7l2k690Sr77idqA72hxxldcLmI/SvqYvFwp3U
g0aqSj0D6gUTBL5ImwBpILuMiIVeiVCsGeKUTHK0d/BJf+jOFBQ2MxyFzdIIbTavcT6d9ctdUOIN
ILdF0vvtTLapxquNpC5qem8WhT/2OKMS5l+UAko0BLQ46O0tIuvdE6q96F5WrH7jkZnvH1TEYTgT
iTII5ESYHhO6yN0pta5z5Q03HP2TsVHidzdvYEJiwfmtWKSHlXJFrrPDC1IzbYaaDmtU5MjZIm74
fuI4nHlTaN9mbK8kMQH1bJIOw7BzgzJKUbCANQidGqugklGAZS8nNwHSAI3BW9bZAZpoZwXnKA9c
3Iu4BJMcJIKuOlP9ongYmeU5l74SbXSff+T0DSJAHlc88URuBHgGh6fsU2D+mY2pd5MtvbYXPxRz
Zt86hcTZSgDCjroP1nXdN8oBWK2H6l1SU3WRLrYYZCaUI0PGO3U4OsiLVn4HmQsheZI4hGkiZdcd
vnSVStgv55ch8ewsC/OZok4z5JGubDguqgCSWX/uioIcgZONkkcZFiYPx7bGCFU9+6ahsLhmrugY
IST6mU/yIWP9VTfSpbQICTDHbkQET8vGil9cVIt5ohEX6VuFuRk5vds1La13YaRxcp1faHVFWEqu
qnal4Jc4IwQv7DP6fdW4vSgxrqN2Yy/nTAgrGRYIUsq6gInLnnfbz9CP2Gbg/WbfzffO8WU8ZwDr
ZqQczQrUVPYbC5gGc/wu4Lg5BmI/kXj9YKVquYACdSxNPNIQdInwlMdh+uESUYnRG90JvdNsmkJY
ezn2xfUxLp9+UBVETzTJ0l73zJmmBKS1EhGgsp+H1Q2tdsiBFUzZ2AOFKr7kDdV5eTwvA6llDeHc
6i8kHWE6cF5isGNwe1HStx3ID0l25nC6Q3f0dKAHgD695dMuCIbRlAtsngTsG1qdRfndMAWsWroB
eRoXOmr3E/fd2Cc4N2zpjsD5+cw8gzqny//pFMjJDsQdOVhlTCR4hlkUL2gIAfAFk70QIzaD4MsI
x8bOVu4gAjE63c+ENyInOeJNk16H6Pfw0Nmy+7QqIINw0MzWZjV6ill6eGUrBSv7nlnSl/38TtCG
Ewqqk1KmryvMfhbS2FTVArtnOzLu0O+z/KTF3t388dDnYZykiDQWCRDBe6Z0Yp/oVcIWLnhDbgh9
mirw5+uKH9RwFoI2IhUXr41LTYxsQUMnsqf5lUF3SPQQ83F8N2zZCe/VAdBfAV4seqSfPsoNqod6
Xu8WX/8fGZ05YHOE2E8EHIrmnS4+jAw5yO8gpv25YfwQxGhgSmWizrsju4e0Rp1ctNJM+BWdH98q
9db6qPUG+g6y29NJXCDnew16gkBl1g6X8Bt6fiNZ7nXXk0aKVZJgUwaGK5Ir6gKLdPiwrwv5gy3N
p9pVoMQ8ZKejYIN8qOLElfSByGenyfeB5t1e0KgIJgXVcsM/qVSEiNOsPX5UZRtfvQD2MsOQMN85
bKa9Wi/cFC+8cnlWhLIbIpMqv2LY2T5qviuxeqOQEE2JYM7B3PaNWYrlPFZZPu8edLFgr9t4a+0+
4Y4s6V8/Dk1GxWibTFV6XJFi9IdJyV16vhbS+LZ6DskhWR9h0oUUJCROtW4IAmam06YmSShIYce2
3Qi6SkGBVeqvyO/p1PLlWlD0BXSVq4rywbIBqi1VzZYANaDGuxTH/cDbzE2zXT8OzFwzEQlIVnwn
tDfYAquSYvT6p7EVCtNpCFqrQz6A//neFcvDJF6EEkglWEPvUXvjZnI4Ovivfvb788y57wItQzZS
U+tYzMRXf/oroubsLpdzCeRwJJwC2kyv2J9QdNYCuAggBecTLU1gMT4gP2kSsECgjLQBDQyXIEoG
/fWbpoM6nWkh/VdJseb0Sjn4J4WWJ/EBUYCPf5qq9gkFobmIF83eLR7SPP1Q/mZxZGSlP/27nneN
msjl4zU2Q4aslKacYFsyw8MGEHj9QWLmPEF+WFavRFWwEWgcauTDi+BpmWR3IZIccn37Ox0yJ5YA
8hwsVHL5+PE7sUYqrUlkZAo7OWXUVBV/UOTXBjDSXd3FyNTaHyjYBg6KlaIb+qV004s3F8XBDjpd
x+PVwOMtAUdmOv9c1pdgc8l94FDoheigikvGeuuAgCfnnMSte8xOSjM5P9OkHe6xt7YNzZwAu71v
fSq02PgDKJZ8nfxb00695a6W3nBAvyxp19zZU3faLHlAPLYOaCW+SiXtEDIFJmWRURcPB/6pcM63
/js4EfMj0H/6f+FAlFJEVoPxNwcZMVKXozU5Sm+QPRGz7D681wFzwVQzcCMVro2YRA5FFBzjqey3
32pv3x1Y0Chi3+FYZN05wJXkYgkOuD+mxDy0LMOptGomiXEquWM9bb/+nMyvcY9ZJE/p6BdB5VUq
y8XeJdFED5bpg06NEgWRzzZj11X99Et81IGympmz2YUdfQ6fw4kXQFTqIjLsHnyhSiuKWm5WAJRE
gYRzpZHFftcyiHJ1vlU/J1rkLJcK667oGMYNJ8jf2fR6vK5H4trVauVRCMGS1yoHXTwj5Oe4/Sy3
nbimShdtWJD8D5JTXYMsqPg1BhM7aWQqG9x2qaKluuo5+FHU8SQz9RJoNBgx+jG7XfNfdHdLjiYr
AH09uPoow6CyYMdbQxkGOV0NCWo0TwNRoSHVZv/DNuZV9ck5NBnvfAQZFAu8fg+HdA1XU73+VK7J
l2SkJls7+IXDtnTKcKVBJ7yP1o31AaJHj9AZk8b4gnrgc+cHOHZ5ypejXp4nMCcEfUjYUt9W5GHt
ThtDhfPxkEMrBP8kNIVMI4gCinkKgz8nUBaQdgbIE/FUHLpCY6Rz8RfzPeIMX30w3E2QjfJbDZw1
+xOPnKX4j6BzirnZNkc4/q+GFw0ADz3MDyQYzAUCAIww/wEngh7rq75z5+7kojubxl5ybgrR483w
aRIqT2isi1zS74HT1ymPBKFCTErMgse+lvHZTAj99vNRWIhG0Uo5tEAezRAkq/P5Nu6N9jG59o14
pvFxE4dxRqPotN0zxO7g95tvIMJ5AeQbQaka5ZdTwFr/96LoRZtBAaP9ulCVX1jt6ckCtd4ScLbp
kycwshtTa6y72twEyXssuML9htMrLxvEyH6Nt+aiYihDR/RT5TP/KSaAzTu18cJVBgp3JV7Yrsl+
Bo0kZNyTTNIbn/j3+JWYDET6EOMhJN5YxQuJf+ZUw3FW5pRZvU0YOe2Cqdf/JIVKew4vuSSxCMtM
SnHj/7MGohmEX6EuMMqKMWH9iI39PdSrE94PDCp1lU2nZYnsYxiMi1XKCBgu4FKlcvxbzEUWDJ37
3bwr3ww5Z94SoVwyLRL3GhGDWDQzkKBv6pEMCQUQ0J8ygcCQF1zCskIO/sSoXaN7w0badIbKsuTP
WOivWNdtF2kCO+kwx2UGmmCz07dJoRgqEb59KdOp8UOSKr1Elo4ORiqgJbp8wARglSBptx7WWWmb
kWPZxl4uEwA9ZqMGHnfGbvrqfP/slXTZJVSMiLO5pz3dVg9fno//+G56AUls3Qp3f0sllaSDlucR
LhVu9jKClyZVRBPNjfMeATm6Pj7AmRpSXLde05pKO4nLT/A/G7EjcXu/03tFNBHWxte3bBY87ipg
Tz3SkT6qY/CcDAVIZ72+Xqm/8Dv7nO88Kz/exQbKv7T0V/BNUhEsRVnaWjzeHuD/gAJaFDyv8eze
h6NWY0+047wmhKiSPkswnCvS91TqAHc3l02lF/VMsawAue5KRaBscA3V5wpowAGfdMkhgai7eIO8
xMEAq6FSLNX3dBwNFYWgm7byMyACRX7lTSrzHVVzmzNYLo5Pv9Q3O7Hw60awhXI2DyP8hAfHWOEY
oxj15Rx40Xk4dR3CuKodlFOvq/AnOWVh5lKEtXV0iFBmuXFg34Zcebf9uGfHVFF3ubUHSCyFCnht
1YhqKGqZm6vBXyo7vSjXijl5UfhugZtqZPFKR15VNlo48BmE+MWjF7CfjXzl3Nt4rGpy5xnnv2/H
lfduhFrL53ueO8ZiIMHnkG41eG3naqS6sksAl8NSdH02go/vfaIYRzdyw4M+JOLqB5+F65ivYqwc
KaYFL0A8IYx22vSnIet0OB1bCCQ+vdW0/y6OQH2c5aMN9K0rMwC149KmfPhINmrN0bS6ZV4KhLq5
fS7BK53yim50szxV0XpJ208iemqX4jZeAxM1U/xEgr8cwHpBgMufmtFfVcBWpqua6kRxAxmZ9QJT
NQGBbcEM5PBV/KlFAKKg85w+1t4Iv0lLx/0468K/10ARsdOnVHdGFEj1B/uCt79Z+bKGblWPiWHJ
P3QrPG0ioYtB4NNM6h4Ki2FGnfj+tjiNrwWGHTyYEneKGCOCTkk4IiXHwXbTmi/Gayp1W/Qz+cEP
7lFV3yoO9LLLA3iv6lw0SGv1k6PguB4JqqkThzHahjuOodOvoxhzEl43XdoYrAPqEA3reQmBIm8p
ODRPdixsQ1zhFyGKiYP/KGSpIjL4I2vEkk3vA5pV40oN81w85cNc4blCsA3Uml/wIXMTSXJigaNr
G/mjLW1RKU1sSSNa7YyhgVydS1nfDxiImGI1G0HFkU/VJm8IWieq0qUN+U9EkKNoEu/GhBBg8orh
s98/d6okPV6HjN0DcdSf1XO7cGTspqd/IDwKU6/Ap95bZ5yVvcY+dfD7VpoxRCY5I/bLXjlp/A2e
gpo05HqPy+kN2VjOZJCgiXQctbIBo2G5lYz0B25uKG9Yv00KtlDUH3DxdHbCyLTe1Ys7nsjk3uz0
0QtW/aqewa4Aim44VMX+YNV0+E6ijg8F3H/eyje8454o9BgOOTlNvOdZeNVlwibmtFF+uZrb7/G1
pl9hAOhAJ/S7KJoXb3wHTiucNq2NFbejT968qJBWlTt5KU3vvmsEozeY8iyKqIwgJLyxAotQXvnI
EiGOjEDgILaOUk8s2SLkdCWJs0yZtJJEnFnEAs3txqkwZT+LSu8RVLtKaDv571HkMuTcXB+zn6yC
MYu1aPYDHAnEdNXfQTjAiKuGNwyOHhwLnI3HQnlkeymTgi3QqjqlGnkzpifMkpfN5VOsw8mzpUi7
M8K3NiKSV30SiD4XjQTh0boAAi2WErOjOP1Ng52bg/VqdUrIvCjIy3QIP4uRO7W76WHMxaeL8Kfu
s4ywLpwfVXqtcZf5rQ9Tpj67u87ERtVItU1arg6Ow0RhVtdZ1tEzHsCa/PBGFNND+07fgwoMGW8v
ku+226NgeA+7CTf1tmifZA7YDG9uqF4mMfdsAv8gI5wfPobxe74c/qDi1o98Dvx5N+TKZtU5/6IJ
hImrGnO+I9SU3wxE8C44rkpsGIpOaQOpgR2qqxEl5JrqHQqJ4FndibGUS1LKlL4hMI1XzaosXoz8
0zxqq82VuD0E5aXM4s9/MQHde+r0ClGpPxhRSOg0SS+AD4RFjfC0OD2tt8O8yPkH+AWQ1tWVxhM5
/f4L6/6RKVXCTDlMkDhxgr3XVrDpo5KXVFSWaWyiP2TquYpDpx+3QmYhMiu2w7Q7HoiqKkuxKQFR
QzuWF6dafZ9Rjl+cxkcPG+aH6HsMGl5xyLl5T5gEeRB/OoeByX5Gd6vSFpxciUWEn/3mvKaiJetZ
qUwY9t+D5t1Ew3U904OMXNgYga61iKOyDNdqH5SX3W/usJ9PnFopDG6h71BbBVubTkWTYWMl6PlA
MgHSO6rOAs3yFcXtxz2rqaBhkWV5Ss549kSWU+VE2wR8gXojk0mVzKuCOHvnXPtpm0dl225FivWi
RubCWECU3idBt6m3siQWnGQ0h6gx98pVYVRY14sQ0F5PRf3TzMWXIqUkNMEd507Rf7/DfitgjNnj
oAtYYwuBTrZY4NBT3h3oYCdd4UHOtKEA63Z4CnhldLLqeIOZlxymZQx2BQLGWkHgoc5Q+NyTPFOD
4qw7xa1MJgUJj5Glb8MBJa3rBpib6tsjtSg4dMh5IazymgLXbUMYDUXF5hkzA1+/mq8zNrg7Yx1v
8x/XKByafbz0zyb1e0Ygq6oAM7CAgiX6Y23nosfgzh4iKld424/Tw/2v0MHghDnXI49P4VWkXhFA
RxYOj42uY2KRfM9T3z3yikQssewe8mmz5aT0KBAcejKWJBF5bOgKJ2vPI/EE8m7AxCYvMObAHnEm
uzK7HT0UWmY8zh5vCXgTwUl0cNsf89r2iyE1aAa4KWjhgMvXE/clhPhspFFjn4Yxjp/o4SdMTKS1
KfVRu0/VmG79FObo1dBRAihVAzSYQPMZMpu/0FwgYbWhy5hprypjcn61Ata4vtVBMy4+owWiW+jS
fhs7iBgnTGCEAczSrkC0c3msBxTejqPqAI9AZpx38a/eHiFbHzGg4LXZt7TCdDmAqYhJmu7GIjXM
tnNsriK1nMJVSAA9i+urCSd2popm5OEKhsAUZTB9BnphXFmQzzvbIrhQrTgRym1xt7oA4RkvHnXc
oB57zkzCpWRzS/Y1gm+dRERTfU+NOEjBn/FEjkCdrqTGy3V/D9PtpMCcxL/0YeglH6rSdmaBb39l
pMIM5FF3li7uanXEZgqQGpO8efGFTaaB7wFZJBG6XX68Zp9JbisTesBT7/dhbBe8gAHfya9mJ7Z6
rdLyr5NC8K/ja9EEEGWhRwnc+8CmMO0l1f6PeoOuCb7PyVxa+G73lE25Pvt31tBvGWwigYSC/e4B
kljQ7qOTDEIL9IIUE5CCwyK9GQS9pVE7065O/5IYlE2mjeAo1Kf2sQVuDT8i5mMKBiXbczWwzpHh
dJ7nX3//CZEcWFXbNTUeqKGC/yzHNUECE7JBpwgC0KFBZCJzflUggDuEuXW131CRlzkTO3GKABOW
TkWnuoVZsA6zqkEcszw7jaUYtZVCGFbIWblj+WaI9hOZJx2noVxfzbxQyp8KTjgLGQBWLF6hGNGO
bcaD6FlCscWsIef9u2SuFyKizt3OR6jIEHKR8/5Id3G3HEZxvItENI+f8GGj430WkKX/axbpshNN
tdfh3D0PDG/DWjBcZcDK7XrCa0ZM5lhHv7YA73PsZMF7K7qzdEzpFWiMtDYkBek2wEBE3K8W7C3H
wcfpPzgNWhyRZZdRfZ/LnXCuiOuPpwGLjmLV0wb1mQIDJJ3HW87jL8S8PIm+jKW7LK8QfDy+l3+G
GvmOxYNZLGOw6T/NgS8hOTeDF8/FvLJfxc9PYxv1SM01w4BV0595IgH5s85x0bfnRpPD8WWXvozw
X5faT+1lJj6LoP7v6M0JLImddbj0LVj3Nd1mGdKtF0JuooiIyumehvp4lfUmaGlOctIF2cAd/E4E
pHN43b79/Kp/RYBR4lSejSMbWngR2IXI2RimPOVe0mA7QdfK3t3UmT8cw/EniXrE6ylIKsczSiiC
sQ2p5+/B0ILY39sCS8FpoaeD79qlqcO8D6ptjBqhabrlovYnuy71b0EVQ6uHDiWPTvXdjSTBRpP3
PrV2reIWt9WR/QRnScHZriFEjEn02+xBlElD/Vdz/IXX67akZoM/xQRd1wSKDiFmkKbp/prlSINy
0lXbXO/r4WkKaXmjHFv6O/HwP35ly2fWGzi0AaRVtpFYwONzM5Qq/KSawGKg1YCHBRg+uZeDpLso
v84P7q0tMlx7yYtEX1jQN0o9adyF0IvBz3f850t2gnMkJfzePN1R+8QKwry+Uz6OBwW+cDBRHViO
gHkfs50FXdjV+cm4CHMcZo0cHqGi7BCG//3kUHemJKq+xXkQJ9JFFzh8ECx6JQ5QCdpcgenfqP3X
PmqfPhUW2AYUTzqtTvgbpEXHl5bWsD/W9ctQQxo1P0hCJjjGelQQ7pWRZNmSXMK+ef+61At+wWgv
oAcHzOO5921AJMUw7nt298rNvXVEC67eWPx/IXLoAOeiUV9x/ilEnZ0XSnFRZaeOhmkGwy/Vse1w
4wVNaGRgVI6aazoY6csPDvsynO/FxCldPl76pIGcGFA/WgUjqHtBzQwvFfAA7McKEwpffWVGWR3/
pBR9mHVOISQsOyrkpK7COTzv98JA7ir/Db4eyFHN4CIFXMVzIoemJWil9GSvynh0tB0Upb2nct6N
o6pFJ709feKi+3eX7M1vZBVvw1aeKWRiW+YPPIEJWSqg2qBVbQ5X4CNFSjXQW5JDjtLJuHU9yZIB
V/FWt84O3o1Ry1RtTGRyTdYt3l7g+0HKnbmZqQdldoBrXiSxn1srOM6NHh1xFbi1w2aDsbF4wKJg
s8Tmeg9Sl9Eeysc2CrJmFOZKYqvitEMV6fyhEvTUG4z2L6vidDSHzBKBu5Fr/jXS2JrntO8+i8v9
sxAt0qJReIq0xWfiDXztYaozod0W5li9Hkw0yP4u4FQm25qDSZppnWYE+jgFPYTKrCDwgZyZzgfE
GnNVD80fOQERR08inH13+Jt9u0cICgDpiLmjBNegJ4i6NrmS0jCpN3A7n8bqQQc1EMnd6yzB0oni
yItChvD7B8t4vqiY8GgiYBgLlQ2f8Mmguhp5+HB3w3B/m8zz83ZImvu/cw7QQVtwEIqteZXiG75e
3N/Ymz5PquSHG8ubqrc4OO3wdn2p/Lc5ndZoGzjeFw26+oinGfNAxg50eR3QmXdTxsepfkSf8hTy
yqtvpbEuDpRFBypcZ3iYuVAV+b+o9Y6k7ALLlsF1ZJjYkzgkpm7WYocdIWeD1jG/z8P8u5V5Xy6p
UlV40dLsg3xYah8rIzE6UPv9Z6isq7Af5qW1Qfb/l20dUINrhMkudkC6hIu4hl1Isei4iFKyiRU0
ZYLegPYVGqcrAiNBzUo5Wy2YtwFoP/zMs3Wp7nKIjsDHXzRNBnK+QFQvy8N/sDlYYTAw3z7Ry+my
8g0pvNRL6mdv1uRdyBoQKpfWQn3ZQOGr3FJEG7pHhumkHc61rac1XKc29WMsCn2lceXRGyfYJiPa
OKGYLbu/lndc5d5lA56YvmUi14sgPWAWTLuRvxdOrN6cwiT/SIaTVAvxRVCDn+viv39e83FYWIbP
vsaCmLgcqiKp7WF4PTYmC7ByvbNmi/N8KVRn7cAxXyla3Mzcb1XEIBuVzcQM8W3cVsdBT05uEgG4
h9S+pUySvrQs5WGRC7G1SB0FBVFcw8CKpUjAXvQXT1sxR5fUixUAqLxjOQkWgd6o7GK1QrbVZF8J
10sWnnYWPeMr5pQpE0/GqOVj6J6yBDrFbThcReGx2TK14MvRjlw1htcMz87havlRRfBH2fKV1GYK
qTPbHxiiVoVdEhnf0jLKX2ttgpKwMJXAde61OOjObwAVUa+bMusVY/pDWSeAn0qcyeUOCkPMt0Au
exSj4rphTf+YDS5xMhT0rESRjzBcGFbnqQQQxqzZVWu1/qdENYE5dZ8mipTdXucwUixJCFBheM9o
hUy+xHz0GttNIoQeEulArdLk4fS5wFob4EMIcB6mcutY3k1AesCSkZ2MKnWkHURtSogHNN1Aceji
dvZwLgZVnzjnhvYa6YBRctQnwqdoqP9CdomXZg6GDMRe6xBsYy+WSo3/CY3UjdQHIiyXp9EZ3phT
cJEJdvoZxjhr9qnY9jP5x1GpnDrSqy34BufsHG6x8zWMeyr8JwA/9E46bokAzzlNHUXeaGgVBfrb
+xTuytqzu0vGRBm1LGCrihlk0P5o/v+oPF4YSFykVPUfb8ltwJZWXo2tJ+ysHAx7Ld/R9B4Hk0x2
rWGWsfSojwJrYvEeTzkL+2IPWFc++PoqthqzKibgZyTRFym3m2EMjpHYktk6AezOp1x4/XH46KHi
BpmBw0v9Ehcz6DpfpicayZbudV9JUwX4lblcc4dhSoolCvqN+4c4bXEHgNO3PHU9sC70VcSbnthz
k1y7suxrR5QmVtfZnlyDsDVTw7PQZ8INdy7wBteDdWK+tCOY2Tfz/AzNb9tWYWCdmZSuFQXxSGyM
TL50LMsX+FRZg1FXPF+KNvWR10plw8P5jhgrERG8e6P8Q9XhDTSzHAlUnWO31+QPn/6FDs/m0HMA
dC01dGrjufJt+OYGJU4HjdS0mFPeBC6igHP1nL7exdYxLHnekpZtj/i+CaiuEt1VRE7ItNHiqJrA
B5LeZtu0nX2BmrlY2bHRPlQalzeuqw25atLmHok0/mpW3jnGWtvOsVy/5P4ql5Ns9quSk2Granq3
pkzvill+/7RbGEiNTGzgrdWM7wwtxhV5a1PuFQZRYMdlRrWAPd4HTC829GMFBs3D2HRSQFNzuoEj
UgrCvVHfb8MGzQr/Vb8eTo6K6hB94uJhhCVQ0o/nkylG97SK7kP3aDDZX7PmXNkOR9X9FvruOH3G
+cooEuO7Om/79+5dNkgSUa+1foTApntzFAqAVZwNv5JBxRQ5JjyKG3qKdZ6TmrQGJdjs0FlVWJgk
R294EQlbtVlHvqYBNf5wM4fUFTTtlz8c63uT6uyDnWkFZCDiledWtHoBDmKalEM8/5FDNpRTOTpm
BJeZHqNnh8cdq1Arw0rXQkyd+TOyRm7c3YHVG8KWj5IrNlaEiQ3YH0T5El8eH62B3F9MZpMpjhM9
JAAWLEXs8xGrCZgppYFHfFaWlI6S+Ha8KDIbPy8Nn/KMew6zOKk1PG1k+eKYuKHwJAzSEjIXeYfL
5D0dfamdD0j7TnjBe09wsIpVjBZGbkI5oBMfbhJywdy39cgh74KdKcN6D+97oMBGgeMa4XePN+TK
fMLXwhfXhGVZMCzqYZI/lAFo3xm9UJ+0mAFRE5/IBB7x+XAKX6ThBz1vGEii+IUpL8HETAqGWp3q
nbY9zvWYsIvU6Z0Fp2M+hX6He8AmOsjY6A+5lgTEu+4WBh3nKaCbTkIGu4jvYlAmEA9EoLw8VjZp
NFOl6vy8pVRlDi7Ygt47ugKQwB5YoyPv/XocCXWW84Xw58oZN4F5n3glu7G3r/jw+uvN5+YcSbJa
Pyj2yKAuk2enaBCc93ItkH8MSizodFI6xpgL8WgF6KOtzFnX09/Ea8Is3zZCrAE/NL6Vox8L+unE
evJeROLJFkVg/KIidn9+sScwvfYYRKv4pHeXVdVRYt4cmULWQGyTyClENPkHp9b5g0CKzQl/2t9u
YywFVwQOJHeIg2SmHaoeYCbw66zB694augpv/0TqLngEJaxETMoQFan+A3BN+moFlg7B39XDun91
/wCDw5S4bRA1Qp7WqZcHs+vLEt9eYZF3xoHvWzfp2a+9+/rxhd04QWvd5t8J4FPPmnHROjxhpW3d
Hy3P3AgUtVuKnKguMD7Zsvj+ujjrENuCsaBPLav5cJSuKvtj78XS1CXd1EiB/vy5sOqA8lge5gP4
3pvbZLX6DT08ECxu7mhNKLUYRS2jsayCzZa5mmzLHsocKFVWOchs7vUOgSzskmN69eFx0HABIsvi
iZMBxbGPpv5PCbrZJG2G4qCRDrSgiKZMHixxPvRYOMsPApnW8Jqi7N7MlOuKwkdXW6bEQz66wIkL
4K8WVAeTIj5SuC4fhUY/bLKXwDPEODdbyQB50+j7mdNCUUg5tY/bcSmAQyRCGtz3ngHuPDviUcC/
RIt5r1kOQl8byCQ5qfv+FSX6V4BjrHJFub0BZEz+JjFqV9s+XXOySV3dkbNR+7BaLGiI63+s+CMI
V22kc/X7DcrjBqe0LXE/f7Grquk1r40Mhks2v7HhQmB/ojIz6mzg/u1XcqHF8feFFrCNz6rVnvOo
Xcdu315sz4Fg+U/cVdfarYDYfGEnyAK+nSX/tbzMozGX9+3wOZpdh+PMXOScWHZ5RWoUA5UQgRUp
D/53HtQ2PnVnquzSTRlSNtDt9EplplP/TG5m/tjZPR1FAPSza9wEBZLqBfMWm0HD3x3A7yzuRmxd
mv3hWH1LMLOz5PzbBUSfHjJnL84V95qk2DKJwFGr722yYYdgIreDXUDB1sUAvSJM3QGY0pPa5PVz
XhZDpMTq5Ax2a+aiTKKq9nGvKfXWo3fNBVlWifLUQ4N5NL0EzOq6JQpEjtlUTzmhbzX0q/nG69tF
kdSIU7ura+ZFwE5t94r1KfovZWbM/RJM3n+f3N8RngZxokHCzT7lqrYuHbiqLmHfBOtiqlh/7nQW
E7RvbTFmilv7jCAYK9tMGeDKjTr1/pYL++x9XoSHQV0E0iH8Zrkaqq3409V0seJ+ISCGBgbA3njs
jZx5kuI03jUR3KKvTDm6/dw9hupJZPixaUycCweDdc22evJ5xJJXfuXK2HMDd+VOOoe+W+cSbhH8
rCBuGsrtg377jtDpFz2ZwxMgILuQCvUfQp+HrZfu8DnvRekdVSJyTDQXUwjKnn1Rv63mRvtUxOkT
ht/iG7CkbvfF+72kp97498/0X4R+CEgkW5kM8e6xuPsHiKUik/ntWYaAbFP9boDXnLMXdzMu7199
4WhW46kddhn0ZV0IfgPKcirAp3Lp7t0ngEVd5QpiBqu2NHkYJWo1PMlMQwcDa7zQz2WNLcmZzq6L
hmjALA3IKt3L+beoF5x8CAA4zqsAoUx4bm8j/6zdz0GTOFBVWLm2/ep2Cu7nr1/v+T8CbNcAFJz/
jdhOrmi4gg0SrBDNMUBKOcVc2TyO0rOWsLsU2x4irY8+T/C2fJovA8/MxGBts4COTRUtJKA+ji0Q
r6X09bk5hPx8I7n0IeMA0Q1FiNnEg8DkNJvuKgPJ8wupoNEtt7WgPl2iL2igXz7bN6mShhUlfPiN
Cgtns/KzUrYo6FkRDGHUlAD1LE737o5yruLXyhq0IEdnM04m0ikB0VVJBDq+/XtRojU2f1mLbtSk
kpNA2IG+EFKeX2vWp7yfnKGXiCVJQC0HbSw0n4KRke5e9PbGkSuR+7K2VX6Ot04Q0quy7FHlAsOk
FYq2tjIPiz/aRkJa6HVnN9zzKUsoq1224ni7OZmb1BkKjlkoUWiZUZ5qYMZAN7y0tBEq8tt6DfaE
lfpgpkoHYpfm0S2a3Wc901dyME+RjInbGiSelSNSejnUoF0GRT3bATLQzgNYP9jdtJGElUXbD0o3
/ORortmWYigXE6yskMixXPwMjfSdVVIOctCc59Tx6oyfyfogKBwCtEylUqaUESAZ9cgKnqyL34Pf
oZTsyLBN3mAyyKmTgV7Poz9bMvut4qhhUZ1/Lw63Q801WIGiyUfXrvOuiNdJyWCd1NQbhSbSo2Ni
BMVB9g/UJ1oZ3asx0+h6RNNTTJ17RP7FIOT5n7ZCCOx13X5woSJdkg7lIXrDa0EEreIkp75lzX+1
t7D/09alIGchwlODURg4n133KXslNfNEwa49fEReqWzgtWB0wWKr9LNZb8TfhY5KYZsRGeGrPhYB
qUfpNVlGx17LHKpEPlzxrk9okZ7sTn4agzPiCvwKPlPM33emHfasDnxd8vUYxcbxIUw/6Hqwx5Vd
Qn9SXmJUvYoVIBIole2X9W7SsOBHWpwUGM4x1isgGWaCBSD8q57s46DRfVBlSy5j4ER68FLW4sPj
QRoDGqDPlJ7sHYm6JS8lPES9SNv+rpqkSvBxgBETcxwLQicYKi4YLA6DaVjJfpLqq8aLm6xKVNpK
OAqenVMVtUXFfaa6mzC9IhOy9fPkky+dEOsd21sbt6L9qAt1+M8+yRZQ2ZEd0uwMVeMsZ8apT7b8
KDkOSyFGeFWQF73wv2zRb6tb+QM9s7jszGlo7MUUf/AHz7MUhgasRfIW7FtFto+WfjMt16VlnFH8
5QimiCmpS6j4XjgeGLsh4ii0qVj+nTmT8aZNNpYz1GHW6Rq3D6VctTV1DQFua9Hu5N/MUZXeHAB9
G9UorNAPor4r3iFiMH3Xvj+BIE4ElI7B5SUdFpUENKg8WL77WHygXpXiVoXACB4txXXxwxj13aA+
8IEDY/Ofo+qwzGKNhBa95EdyioYQ2REYKt32VI5AaV3qcXuNw1GZn80OcDPbUROw0vIqr8Tv8dRb
XonlE/gfnaJ2g0x+4LfdltvWPrxTOCUuwHtMkzBxu2ztNbi1DqcVva2LpR1juhnZjmCJKjEhgCBm
7GqS/RKQOhBbCEst8tm6NwGuyligL6xdVPU4kfFZxvWC66zE6vzUm/BdI7TEhRO9WzChmmXm1wXq
DbWR9xqc3BbCw0DmOswrlsnEscEYODsJh3OSXNBDd4KNO0aZoYL2r9Mhcf2G7jtxJxJ8nLz3xfD2
kTz531KDskT8EmQfaHVSUPE5SOrtDturJlQ5fsGuEmAvk6iH3Qbu3PivQYZIm8NPSouYiERzkzSf
esJcPJPmvoJEL2fkc5CLNFZT0h+PqGns7t4j3c+YjfnPnJNXFLS1uEWuHVDRtTCK5z69BI4BPSLr
HJkD1m5oPUyOaoZPjGyaLRnT728gmLlvC2SYFCJh4tJ6ADzdfcZfq5KhFFgwbZRp5D8bk9cIG0x2
+dNodweFPY5aW4IBDpOlmzE9plpmI7WnW9wad2iSvuLXsTvaTi/MvtZ1blwLmfOJOawTP4tgZfpY
j8J4iARZVYhJ4240qbTJ+M+gF5bZKYXsUPUcim+KeTaG0ShB7TSNclDZUwSB/z7vBPE4/Jt8lBLH
X4gRZEABzR+S9ry9/NrftvMxoeIu5GPC43WlWvDIhgHJQKE4+M9LZOSFNy0w575y4P9u/3ozUtg4
7UKx1ysZX87T9ktd9csMxZzAjI/bBwWk6E2iqR5EtYIL+St+uDNk0B2sn+822eDPgb2QODaFRwl+
sWjrkRWZW2/qYy8EHwiz3S9eKxPNJuvNP6qldGbD14Pt0Y/3RdQlRIkWNdB7k+6mVxHmrLCdBhT+
W6bwFzkCouB6ZNqyvOT1H/njFSgSq5SVivYjvZGgsBQvzESHTN+DJDv2es+UiRgJoDK0bhOLFl65
cRGpAqEiPwXxrhmlfTyMEmKg2s/GFhHOSl3LyxN/0s3N8kPDtJbSfZtzPUVEzYRJqvXspYQiJEFT
9axQhYH4LZRjBgkVV1mtZCDgz0hytpCabkePSoX6DcvkKZjNwudMkZwWQNUl7gZm43JkjHivyrXr
ME8A/h3vO6KOXcWMDfcUmho4unSLRGexUXNezNuftwYzfORY8vgsjg3AO6ZfHbrjB5IhBa4jZ+bK
nBcbA2mnq1khukrc69dQ2exCWYEvV8WNIZSB+2U2rwgr/PVaSuAjUAurc/UKNUKxwJl7sVgOqe9u
y6AkLdNfPu0lfzeSVs0YXXElDKTcFDDu92RILwRwHt3Umpk1oEWM+l/zuhHotrYHSZmFiX3m19CP
GoPbCnjIE75z1TJSVh79ikj8mHEshdzrCkeWHqqy1h8TIsvLlc0qw+KxQMDKGigri29JiIw5fOKL
NceQm6jgk6jNlwXo/ClvaDiDh4nXQJY3u1UnKJ7oc4/1uI0UYe7fEixeEWTQBGjQPCyXhMbkg7e5
VGEHaqXyph/2wYsnU574CZLbRy2vUU6pMJ88spRs2PJSXsfP5weof7BzpxlpUCQuPbFBZ5cqdWZp
eC0KhAqgLh/SrAhwmy79vu+89FMS2bn39TCSv46jlz2Tn7lNy5lNTGyY3Wp8DH0sMfciXZmV33jI
EgL3IdRt6Mmy1dLVZ5lUg52qWgykpb4jwV8+BRwmgWTdu8jqwaXwudHRZcIX4Ly0KRyTUKZXiBzV
cY5heKeIxLa7NPBJ6h6hTYZx6aXDRivnsmHQf7KNPimc6PfpfZafw+Npo+7ADIyf0t635rs2LEpE
EVThnHWZzmUiGWJX1MPQOr2YK5r4q32kdI9ZsQD7nn0FXlhZcHpaUIuLZYE/ieA3qTEqi9o9tMsj
qJw9W81c/lHnxd9+npX0SUlqn4eX9gsASuan9+qrzp5v/dXJq09gJGDphEbSMEehht3Wu9Er1rNm
WQeJAJQwpSO/WuJtpQU2Em+J71mCLRqoUlvWnYytp1tp3p+kAk3jU+QnLlrWJr673eo3G/qkCJvY
U4bcEt9sl8x6bXvPrxA+9zr+T8G7ZtEF0skCbYz986FHR/B8rn+Y4ApAXEdkpvUL2RIyzNkpYATh
+P4OfQ8OnaumUoPDEWKmuPpuz7CnLHg4+u0mT3OpSLeCshmx7qcs5UU0V3jvJBZLvH4kCjOZceHg
n1hq0I+PlpAeUSclYBU0V6jU97LzgpfopyQivs9MHLWsHf3pK73scyW4STwKih3jwPhpkzEvrsnC
f0J3W7PO6KZEw9e5uk6Z3YpO6oFGb4VAMXQJdnzMdmeG40fArYD4zNxMc1E6S9DbPs3fm9vjcyUc
oSGEJXUDB/mDqRWwrYQLTEaR2yxQkBFd0m7vTaF+ZBmSIV+Kxn0hOc0xjGmJ94xL7aPR9ABLVQ11
DCuwixBMQqy6eE5i95a7i0yEeKyItQob4O88LJMkWZsxHNKZem/uyLlyLMKPzOq2SrwJJXUGV9W0
2EMZ2NBaObjskgkSpoATTx+FjudvlZK/poSds6siScwq5292wwX0GhFQh+k01LAVSI6zJW3V307A
6ezy0DWWRkSlAIKTmwbhN9BJ6G1HI9e3xm1+jrkdszUOCE5BcTXo5ezBVtF/1Swu3ovEW+6HMQMe
BNTOZZoe0D/59fWvukh67eeAMTkTws+MKizT3ApKLBQoTVAoOyW1x88JE22mSxgvzfAh2Ff0WWrM
A31YCozOc25Al12A3Ot5YPH5vApiWi6Vcwkg7LaHPPmIB5WbPZYK5u86RFPmVoOp1JFEqMvRdalZ
Je10HPcgHgl8grVGvnfoTvte9v2gloqem/NOgO38GIpuaK1vsVyWwWWz59j7LZikBGq1RuMxia6y
rw6T+aG0yqtWEZE55BA+BsG36+qOZy3Jf7by361/bmdm5LtYt58360VSnh4JfL62maSk/+avD05d
ZVHRv26rWynqmfXcvowyO9W5H1x6roPNw1DXSvY9PoK0QqJKqZfTalicbJ4iDeqXCo8JgcvIJn4a
znWttxI02p0cnYGAYCsahiYfSV4F7qdLTYO9kWz47dUadIoh1r9za8tK6W7GiyZ+1s/DoUtcvrna
qzx9JoXok+zciRYRcgIph+Qt5BEXdjKYFj5npuQ8FZ8TASLy1tovrT4rg2IN0OCc76bRd9h0xVUM
ddjxPFFn2UcNCQcsagPbMjnjoGzLz7+7tKbHmFiEBCNlX51sN68J28h1NJB7LYoZbnlW8oyVYnX9
Um9WGTTsW5bgIJ88rAhly/+jkkAwfxZWdr8cRF2BmSDOxJFCARHpsspuby2v814wtEAXKKunsVkg
SHmbtOs5WbOtHNIQgd9oKuDWIatHw6cpi+FXdVFmbB/CIvsvbYid3bwb9tovRnrKLKhhbpp4TBb6
kRg5XatjneOvy7WqXZqJZmdFQkM2zXpuaHnmlxvrjbx8DPghSyUtM7DOZL2/XXvs5AlJD/qTDWHA
Q6N0BfUX8AmpMYUr5VJapqNd4ukbAf9jD5bD/b0gAuvFrh5FpypIagaLDCbTBhqX9K4luMdQwB3H
cPo5li8/ljdEq2bF6/lHPnCzRFDm72U0kKEB9CsBWa8rwH8piRKK9+PJ6scaZYbLliJTUAgj3PDr
3gPFkXFEYdI+wpl/fw4ncCg5yfdbWrkb9hDC2UHr+BEIBfvxbSQumYhAsnlJskCKqLkEsRsNLKMw
nQcTAZAYSe8SmvFQhV3N/LJXBbPy8tB6n2mdnNhkBTPaHHmch40NevVwv1Hm8+a+zLJnzkDxG7ZH
6Llnfe/EK5kpfz53cX39Gk0e5e8ggMBlqCq0IsmAEZzpU5vPW6LoZ+Jzt2QWBcPm4AXMa5rnPO/C
C1z55HqjcMM4urjhcI0BhjXlia6y+rKXLg+3a5/YNyZz+hiWbL2Z9Lx8bVkxJrjetcEToXWreQfS
z3iKAEQEJSYyRyyLecOLjC4ZmylWUtA2HV0HY+eTCfYHNO1a+LsObSxXWgmWqMwqF6vIaIbGyhTP
sjAc8fiCGe2Idnqj10fhKocNjyMLyoLnaOOUqNEiDXQBMqBf/xisG+KyNmGqDp9H+IfUG6ujJfM6
NB4HgrQpdZ32wwu1TlMN6b3I6HWal2kOz/QX7cGdBrXXeP2MbRIyPLAseuUFhwojFBDIkaI80yEM
ZX1zUNpU6gDYI0Xm34orVdVuw16lAZ2Cz7vU92l+iWvP9D/wWmUkg1QNOa11pcrBi2BpixUDok65
ity+jZHHbXf3MbYYNGNSLuidIW5kAul7k6vVxVgKQNVNK9VrqN6o35Cw2BABIXraOrziounbaENf
bSaAOvkK7k26aJpPzW/hFLtVAPwipCdxF0w3JZIN8VkXdoRq1C4yxbgL0y4T2+R70yOxec3qkD4P
Hzo6fZWZketP8V5D3GCikQI6TtijqUR+Ziqdmyn3PEDPKnl9PnItCjx/vTbcM4re/qF9VdgLzCNY
ODNZMXCqEO64YOgGBjGheUrlJyFqzfpPxYvDnqqy0DX5pbw1uypEWpK94q8HUuNtda5d7eQLgBYx
4C+j4dg6x/KBbm8t59ewwJ1OQOzsxUwl6GXt754KBgYvEttlCsmSVKZ2Mf7TmC1kVMxGcHo63ePu
qux6nZWHBO45YirF8/Y4Uyuvll6T7SbYajttswk5SHDX712U0jeknIzrgWrf9ego1MLeHIqUvK9V
0DHRGcqXomB5eZCswIprqg8tNff8lcqMBr+VROa9JW6AWJTD13uaRaFB2SEIkknkss+kbsdsr74a
dKJHpm4h7Ukld6cUepQibVLyjzY03K0do1g8hEgcdrC9bw0hgB5ZYLT/63rMQiEya9FlVNGv51M8
Gz1SDUhINhgmyfoBkFtFoJoxzad1/ijRmOjwl3LuE3xevGPFe2YfiyE6DJZOoKR76SW24FCLKaBB
EsscOPoPEE7J9siNERmhj7/TgxAlKfLWgUl3XjvN1cAcp6/ShwEREMnJ0C6rAX9AQ2basjizZv4x
p2xxCuvDflVXjTLxP6lZjJnzPp/Vux7lzGNI7chR24XkCdhWXk+Xnw6EXvpa4b3LGvDu43LxfHPL
02kkvjt+fsOdFkitdA7xhf0znIKrHoWZ4rvNprBjgmo/nshzUwMRWJEbTfrcokf+ztUCL7+1Odys
iVe9w1TWs2v5ShvLodywPwyzBJlqkzPW1WPiP2uTMuSlxrrE8BrfvvXksdHL1JBQQOKFV+s6L8cG
pkr3DVXyfp1l0IJMlAEo1i+bN9ne3ujETsV0BoHBiSyVwDx2QYQ70aboto6FksNZ8/pjiWW9lY6t
PnFv7lNh2vim8vrV7QQVD6KlO9+NbdzOgUZgLEIg/Dvo5Nf5lfCV/YzAIPBHrT8fnoEyfRYBwnXm
B8yECic+jFIDScv4FkuDFNaADyecEU0O2UkNrkyN8byIJHscgbza3mw7AzepBmzhRjNniSuUVvYK
BSHa/qiS4hK6EJKqHCgXQd63rMyfOlJxQr6iQZByT46Le1YHUSb0Ft8TTuCYEXC6Z8hqSj6xslUj
O55SBk3Q9KCTGuzmkeuBrzXOoP10zYXWPz94qhXJ4Yg097z6SU5UWWPxXR4mxs3cnQ452+7SKWCX
97tI8+gjYiM6wf40X7FRrQBmxWwmgueORFfAu7aZnDwQWAfdwBYRPrDKTk4/VYnYjLF18/7UO0jb
VNDK8HCKBge8aerGz+LaLoVWgcPjg2zkyM1W2fLkJikxlLyBE6t4hLiGUqwpMwHFdAHj8Wgqtyua
PL1fmy7kwxD+MGYnxc9PPtHyieYSfbQZPoKciX4IHVdpUhQ+UipKJEeQmuoeIVV0w58P2jesUNds
+kPDzwOLcoiJVn1nc/zvFA6bL5qoB6NaNht0QnXyEHj4CkckGXr+sDYPhMcqtCxNamtPu55SelBC
sE/g6SqztIDXlJlaH2BhCf455b+4AczS8MJngScAKR0Lxs71Gin49jQ5vNLQ5FAGrW5mZhFjowSV
1FnW2/9SdREAWb8ML78A1AmVhvuEJ3JdzhlY5AjyLRn46huH9901B9jk6PjjYsKvY+PrivlEQCvm
S3a8QedosX30m/nSg/Jfjkbxnla4kleMcvPcOjNoLT0yIAOiyGb6L5ysFuASDrVAGwVO1vHxWUjK
1/NTjp/BpwwAk3UmhASi9cnuuS785AyMgpiwJNKUSDA9WA2ihF4Ukvv604CQiEAwLgr/D5JBgkBI
iRtWOvrRvARg4elakBoA/hHSXUJfG/AKggsZj5vB5qdYUUqz9loEZvLl7HCXoQAQrOp+gXxaOKm7
99hxFgfl9CsIS6s3bBVsWJYVUOpdLK4NqwZaUrHfec4akmWEMzSnU54q0E2hmDXb6uZ7nalD3j3i
BTsDidLx4gFNhSRC/AqaYMuwzby4r4aC1ncw6iCFzA9MT4nIGYdlv2IWza7BmfVRsKXei0E0O33r
S5wV8A+pEtsHJjEo7Esbu3w+F/lj8Na4iq7hrDzQpp75q0+U7XgAJcpYbta+RAwQ+i11FCtyksyl
KCptuny5bU3jY4yAm1R5HI9ZCT/T3VJjMwbxGp/SawE+SWpJmLpjoVseZxf8PcMycyykqlhFU08F
vUqvHnSXLP77G0xqxLl6++/2P86GV3BKGqvC61LCjjCoZoEJcgCdKG3RIeVmz4NUOWFfMOoLNw75
Lm07XM8xtCT7jbiF58LrHlMMg1BGyYQkdYBUM8m5T3A9maCbTK7WyAoyknlzXakVRBR+KIMn4hrU
xfMj4irxhCv4RVx8SISkVUajx8djR+EyhvUQEm02qnuaYh4uUIEqmSMYo2VYI49I0r0bOEZRlei1
w6R/B5GNW5TypjfaCfhhW9NHIhAe/3zpO4cLctN+Kg00g4Q24vOKz4guuEb0q1o2IAQRfy8dEPrx
uEKsrcMeMNUn2F8AyKQVQw8dw1cgneW92rFpFB0dCyN5qpg4hBJN+OhfXSKacgcImojrlYEgWsAX
uh2dkFC/7tAmnVVf/qE6+1GkIPe73MjBAvfW7UgNELNnRbK0iY+bCHWQdIh1beMXq+EVssDgMEdB
x3g1w3mM5ZInnzpZ034VeWWdntYgrCT/IvHDpiOH0zeKB/x7mosvlN3OeLDpRlUhhm6b0FTrVBtA
DDmMFzKQIoD9cPruLp+CxoAFtBBMpRsoLz/3XLpd7Gz8g0UTCfZviynhKCG9hCf7O8F2PjJx+YbI
fFdD/6k9ZGypxwzowNi0yS7R8EmwcpuOYhaM72RsRzrxYeCVc6ZkMuLolherKLvJXnhbt39E50cT
fkYoDBnaGGAFL5faXg6Y707xBiTv0q/8qJWYx64PACQulqZ4/ic2SlQOhaHfU3GJQrR+gHV+8ve3
/QRaV+WEBRzOxbVUImm4XxFKthebIarvkWmjxin3RDMQ2KsiVSX3ewwoQ2ADGIMun/puD06Ggvum
B6factWRkLztMoj4wPSb6ZFTOsVJ9ZiyHAN5Vs6YfvCtq5/G8TcO6lK5xJWx5NzwEgBLwgXIa8H0
1enBDxwWLOUyRuzrezEc5SaXov4xm/5IwFh87qU2dH+Osis1V3e/L0Esptig/NjzJGi8alV7XXiM
AuJd3a/70RhyyiHYnaODLyvF5ZLtSZIBJEY59R/+ULsWKN/Cq/NxeJCQVaJk5R45hp5i6+GzEwM9
SqXZ58l++3zEvZuEAJTg64lbd0DumNQDMV5fIY4BTa2NiBbFXkp1CLYcuemIZ8CaChSoQ4y8A0Kk
ZrGQn+Z+1ToTm6fKwxbXVY07bUzPtie4S5xXeiEXngNe5mwx6v1PRiEXwERvazpE2s3wN9WSV+aY
3A5QVq4aT33ljWc+iE9D6Ny98oC8Uux0q5+ltY1rPzlPEeBfls6+cFME8Zws2yCnO81gWj6c29E5
k3uXBc4aonbE0c6cPF53Pnsb7gpXWog1mVvnvi/kgh/hwcOPHceuhWlGrE9k+CSOqauQmRlYlzqu
lp183sBbGi6FoirGVGt/MOUiOpYd6FibabWpCiSXcokE1Z93XnDTTW+LtqWS3iDa6h1xceWwj4tn
m4vwoOOglzQUYnbmdVrYBGM9lxxbCfOzs0J4WWLtnDkfEoeuHgK6GyI1L5Bo4S0X6wvt0X1np+kO
MpnHfJf/Nu1s3gwlfcI/m4DsvGK6vSyKgYpMHgSbH7DHfpbbHsgWqesIyCH44++R0rKdsLwlQFzV
Owy50pDgML7dT62FZAx0/Y9HCru9KssZXAIDwqItV1fX25Cv5VtOiK05W9OR7G334R+laJqOi0f9
mPiKXG/LDUdcyNUxlZiwMCzX9n4o68Wy0hf8RDmZKJYj7Eof5cEDLawMw0/DxbCTP90SuzlnEFEk
vycRGASkUJlOMYw4N4U8a3uN4q1tvOfRVza/sIp2OjsPUFYbd9jqSRwaTLYxIO7i5hntKBpPXVwQ
tEqAYUs4m4q6bmCI6qm7ahu4C6jp3nzqx3+4bKjkQ4KlxgjpsH6eqLkSN/ezrCTmZyvJCBiqlX21
39cS0LCGpivDZJljtqoOKst2qe4lOcO3qo+Ve5sg3G2pcICRYPuYqD2NZLKVsKo3C2YM1KdsC/8n
bbsrrgS2hxYCt7tVQRdRDE26N3s6gX58gMMh5xPts/FATLag9HsrcI+4o54MI4nNZaGAHh2VBY17
/W+69j4BOP5dXE9z+gHTO5sRjhubY505Pmpb6vmPs//zlQ1kmaXqrGWVDyXfbM/3ZE+90HGLqQVM
IRkYqgetdGp72v0xmgOX7HA5u23a/zW0Bn8pacP2lCD4ILjKzCpU+T7+Ms6KwQ6aLUTzR4Db3mT0
nYx6GCgvZi7zsBYChETk6MT/gWkWo8v3dtuj21jwUhVsRy4kgxuXOkMNJsOqdqB4yT3wWthJUnUs
eFXqtqIDjjKL7kvgYkZbZ5DuROH/+HhYkoXFiyNADSBUkOpKdxc1OyD+6RZtGslBShhLezj8xJYU
ruCx/oOUFe1YQvnJrr/duA7qb6N0ECBPgwu1SXb6Ou9hR3oyEowOEh0Qg43eiIELUqtlyzNw5gV9
V5bKLWEOFaF2pYNwvS+UdEBHR/KE62Ul5jDoZMgxbZzAq0zzzBTfPR5WgxYqJsZ7k4nFrdvvCzF/
97T6ybOnGFRXRbSJhnHJ5PvenrE1GY2FVVbm+WQpQLpUlY+nARO9jfajHVk2U9lDB6zlyT8Om6ho
69yIkwiw8JCLF344O77ORTPjj+98vxP1D5H8lZGdto1lVlRdR9NzPg/SjWR55cVup+xsU9Ws7gXo
a5UiMWDS50B6N8HM1x+h94GOvM+R6q2adk5xnNXMbTEzr0gSpmGRbeDXAE72F2UG7PF977GCMpSa
fR0E2pEP7WZPSQzmHgvktMI2EPRfTt5kWmWFWyDkYZKirVIVlnjgg3vDGAGEQmev7m2J6pMoDEQD
G/bgLCYRsZ8agc821MdLDdN8RgQ6AINOtBf2TWPip+U4t2atzPSlfQpqApwCWVYIrYFfbpNY1WRz
b7nbFiUOGgEQJsHVPmTU0h0wkyVf53WyJJvewMGL5CoupdcU10sOZIPoGUsqDjZ2ib2XvJzE+1Xg
MHkX5Lg2yzTjk5cMdO5K5zqYtjpch9S9KKFLl0EfzUFh3VeB2qwiTwosVTyAUcBTjvMzG7W2N+pP
/oHRMXW5UTgh/uMB0NRTdr6eQGx2GjbBLyUiyj/Szfm2/6SkNSGR0PQ146GVOja7KTnioQNIW2Ny
Fes4by6IYttKwg0NauySTnVSayVboZQa+XGfwOj6SpvPL2RhfjUZqtn9AjI+oHIkuH0kIvZnH4eO
sXCp0KyEP9yycBAHgM1nWwXvSiGjRVP3y/fjHDEcUqKRJlw7w8KcNumki10deBLJZbIvz9/rNww5
j+C0xB1WOsBF039Qvnh1iHLg+O7GB0ObWJ3bEBoO0v1T53ULt0u8I8ZCTTyPJRhfzD61++N+yywN
6n2QOWhilW71uAQPiBNI0j5hSsioCmvAByDxtiYvIEFxIgBTWFpRZurzaInWBmdA+/VFdf9Yzdbt
2AXzIf5HKnjjJzaQg/7tKAHIyJzWF53xXaqLciwLosfCOaColX1LjAxKPCfLOZLwimpEFcz3wb5X
K/St3EWJ9rjmn6tUZj88vpmSP5/pNwRXxkop+5w/M4cUrwV5f+Gkvuq8KDVVY4IxSTSKVgrHy6pK
Yo7CV1pv4B3hGyh4/54hCh8pEdzL6tOvWHWjzdhLm0PN3OEAMbvL8Ti6FCJVpojbSx8tRortWd15
Efl/muDpCv35P2bTmWcpdwJyfZsJpSlrYE4ClQcfCu5u+KnA7pW2XKSTMTgNHfU0erYdENqoFZqp
Prqrv0kJ7XQcCaSUwM+Rwkq6xcLjBR8bZ//YKxrKa9Lofztth7vxT2CghqFme7Fbk7hgseMI5EId
QhlpPKxp1DJD/sGqbZMb4Q/EaAsZ/XLj4q6itZv6oPbxeBTuhOrAoADeUhZzW+DIbuFapw/H3nUc
gIgbSFZSERPPltuwetUhfguMr8PZnZowlJXYTXl8IwWjagLkFGj1rQnWh1ptfHkuRj4Q5mT1dK4m
hVtmWMnWoLFTAdx+y3+6S1xfhN05HG52Y34psXH3/6eoAmb18cR3h8cyA9DC071ARmbvqqS/uqfO
HDPR80InzQm3p/AVgolUuOV86800KRDDKL4TiYa2bpM/NcFdV7DMvCBKT2iuOZ036M51OkNHrMxi
rA6fLmQyLAtzbYDnEz/WvmcdASUG2Az0zkNGCY4GiLuj5WZUHYxmvfQ070dFMGmb5VVFb45Sr1o2
473tTresQD5nUgRIXHrY5M0oWSudgTTE/8lgERahmd5QZpVVTAS1Cui2/gpVuoN5cM6I2ahTWlak
RP4JlFPndINSDgfI8hjr6dLSSQwO4lsKAr8beag688gkdxZwelKRQCz35/NW/Ycbr+VkWHjSH0vh
0vAeD1S+WkUBxRO3NnDlEsucxRxUgY9qZnccZKPowv19kfS0Ncrbo1CIRsruOxzm15Md6CgpZSC5
9SYj9KE5IBGnTL1x4ZC7fJDXJAKT+yx1T9/ukt6BoSl5qooZ5cdy+uiEIkFw3O2pRwfBVR8JpGYX
aUHr7CiHaPZv4Ajge96onXl2HrJv44uXjJruWKWgXzVzJ7NQsyhGYNvu6cgjBW2lel78wLOfxtJJ
gGReIkgaHz0S1GFr5x5X/c24Yezqsdg4FtH1/96mngS5COEGbPONYE/PBKjUx3lEA5yWjfvWaGfj
27Fu1vZME+JnLHrnvPsJI/T6gNXKYHZWqiElKIRH1/cndoBVhoqGe2yQOOUR7aTFcpnhGcKbTiip
7oDzekE4TZ02ubOJvvkJuv46i96eyGOI+t7e8ww67jFqMoQr+SJHsapQRgzLg66Wmj9uYK0Eiafx
l4SrdKBOB4fQCypPmxIQriS/iDALt9B/qToSba0bS6RDOXVhpTBVsIQkwJ0cKgbWPqfa8CSDRI7c
Pga5rfKdMkhoi3g7dZtDBM9BU5WprylN6ffE4sQpuLen1q78MfoUFyMijqjgqL3vpKXXtdPn9h51
2ktwxVmiLZ30AEEszXk2ucFhjtossQPrwRtsCGr4tqXrPyGfSXNBfNl3jkYbIgOHs6FL7u7NEq4Y
aquRr9saMvMQUSywVDAHsFqfjmJGsZRCw/zcT3QCpblfB413rH4E3k8yLkcUzoMnLLClNuVpXBil
TO6Y5dCqfPVQHxVbnqv7HwMW4BLnZEfm+WMIOyNd8Z30SxZjotCAuC6idbW8sRWBzlZsmfkkfFac
xQpGZwM0d76TGQia4hBa12Km7WE5O+B4hI55d0pQGW+MC8gDUSLDZRvyCak3Hnyifqy7yCLsDpNR
CIGoJ1cOdtFUH5tWDq8zKh5PSBagDwGr8gde6AI3mT966vMKNMRs/xGJRK3tfM+UNB6dj1imY/E+
1LwFNNiXZsEwr1hFzxcZBdDJkT57QvLy739oY0q5fNGTyXgx4EZHFyORY+P7a2xEQi2wHw/47r4E
ot0n7bes7Ad8bumN7UNXRX9elxak7wKUxyESsp3eI4vP3VYZ//TEL8KGCi0IiyvSfLvb5mwlITdg
XJTIfkq36WLjImjcapJOTKEXq81vKARTzvLM5GaR3MTomePFaMaUaXOYag4IR0AI/OJO9GtEvGLZ
0pgGGxsHCb3WsvrPCKy7aJ4pQ6u0oLFl+L/GrwTTrmtX5zCzKq/HiibxRsLM7jem8BNDAaBVmgIW
R9uENsqs2OeUFGW05OkpbYUevsOfCp1GR6nVnD3rB4KGvMmIAp11v/tC5LXv2LiIjLlULWDRObfk
3l1KEgVgDGlFHeX3bsWTAd9FQTKU1UAktjz5YYkurF6jGLfcb0LzBTUY33i38reUAdt9Yvoo9p7G
16jjZJFyAcijU4H/+4CFdhBhakpHqVkWF7DJB5AuVhoffpiX5UwVV4u71S6rCHCY1SY51zL6BUUE
W+apPnifCfj+woCrTENNBDIF3UBHe5nAU4i0hxAjAsG7REJuOnpu0TPmnJPhDPdR3r6dkEjoeOg5
bEt3F7rWnRFO8WmK4oCayDmyZe4D3REEQMDdCeGCCRlpYe6CRUtd9ZN/OtKsGQHwDdVJ+gknNCTj
NSN5hiqxKwEG29ahlTHJT04frSyOn5ECVXuaDHtvn+OguMEWwJ+b+p6RxZogHSwnMFwfos/Xq8kT
kY/rNWX4CXrW4cUROqxRHcIgkdWP03BRIkZ031s3LUFsP7kSrlPj7fwYKfVNlBONLNG0lP/rI7fq
nzEi3NmBvICzxvmjpzYUSwjvqQFyX/HsSRJOJkXFYOwJ1P2cxiEBa5kuWPzcxKkVq6k3+GZke7F+
a8G/AtQn5aBMLQvuYXyr0guBe96t9OG65rhjoYKDj3PDwz0n/ao8risj5u1e9aTPx90c7H9IdFac
YfgQojfJUWnObYIHNmShe9ZKkUsa8PL+AFP8UP1JU94HC2WMnpcDhDDiqkJhrpsoS9SF62nUY4rE
ZOe9/y1uBVhgj0+BFdjPZXMIo+jWr5TPjEiT0TAV9xg00dzFtiYStstGeknNE5Sxd0vlj3R5Lsmj
tO1on129jRuMN1xx2JSZ+Ij6jlKll8yJjlvVc5QESO7nkzEJBIoC6w2EmCDG0L9muONNW7sH0bHi
xg2vodI+zLTquydQMOLuSURRBqyD5w95L6zuK8I67fXMWIUdeG8eKkGYeBS9TxR5WEEVJmLTsO9P
wKVQ4RXuvdsWjFBMmEEo+78JQdL9SfZROuwJgujM2mhRbOcIyo9PTddDXmKMVWQSGWuo/52cTXny
XakkoJqj8WnM5qmaL1jF004M9ssjYv4mxkswAG+6bdw4i0yn41y52zy5AqAMKTy37yslD55svBm9
5cA8e0UiujYjAfjYCgeVMpeXbhF0vdRtuPxqhlcYdGYSFcFUvocftYmQ9ANI6+I6ue2bI54QNYU/
WG7g4lsXhU4OLgciPLuW15jPL318a71iwyx0psBg4vcW+8pTs96IUcFY73v65dJ7iXjdKo16la6s
HA6LpstMUk3ADJG4mqdNdhUDjyre1JBuP8/AqBla+WR4wQS1fl5dHD7Ot19ICAeTCL0YKxZLLZnU
BtVVDzlOkgaIsAjJfJvaPV8+8F3Z7P1aXA4B4RqbHYsF187nPEKcQEk3Eb+qvqp2fdjTA01J159i
4ITb21wgX4NIhetp0+xuLQ21vVjxU2WSB8asG4SnAYjEsSCThq7ENVfj4H6jQxlp72GVyy1hjwZx
/cSE65cER6yG8zNZXFAunB9LuuJJWONrN5Ges/e9SyzBCRy4+YxhfuRj90Lm/yVZFDZPew7Sy2YL
mFaJEQXWTvUvN7pD0E7ePTN6jjp88bAzEbQUab33SnwZWIIwiarzWltLtpmCCgRKHLbcNa7g5KgX
ZDNo4gfnU6YqToGA4BLUUDo2fdDX5McXKBDFx/MPZFMCX2ojP2VNTacV0zXlkIhaokPBGINx6G8f
I2UAIIp+qCmIeEBlhyDiftaRwhoTzkeAlvhWMVqeDkIxYgjKM1tUJFfTCKAqBejmnb/82Jb3jwDN
MvuTQXsaMrxx7NKndTJlmx19+9BNDzyCSLmrMLt5rIJWeSpGWOBhJzghSA95yQLNqj5sL7R4BzM3
POdocAQHq/8GvREFatEOcbWYgd3+XQ8Q+ESGlWC9OINvpa30zIk2oxuWRk4uN0utQde2F7C0FV/W
qTgUp2bWybqersOGDkOnro7yqO2SLlJx8T4KhjwgfX8JMFXsnZUwSV6rzW7/r2bo/IHJBKfF6Xch
QOtZwLTIR5L0k5TpLNV45JldJrSz5dcjuAaF8em6TcQOBtTBGc/jAV5QLo9ka8Aop33O9KKe1Yto
8YV0wCMJQqeL7nhbUSi54iHYPivFDsfyBNIFVNPxxcnsOwSd15HzT5dLRsor1NHhMc/guNPpkHcw
CPsBJleeegA9M3LxzhAK0XfF731/vpScjk5kkFwm9TKc0D6Ll+dp2cgeVzNsxEOjSzakkLsKwbDX
Vhs4BLtmhsfDNpwqdnI6inQ+V4QCPR7uS9564r2SuAwxXWFpfpDZTxV8rxfZbOUltmcQDh/jXp/b
tZBFqqbctSm3I2MHsrnHXyZ+dKplkfZBnv26PxAVYSl3FkBfqk8Ld+EQlbi3I47ICbqOKHZ2WQpN
oZRW8PRErCFu5Z8XICt0tkTsDppbTLiYEOZw5+4KxSbDttyWwPz0Bcc4TCvjSwdrwBcgur6yJkzQ
YAPDg5TMGuL/n9JOAZM+IlKIpHeSDqP9jTQQH+z8H9Ky4T3guYytaZja4cSFz3faQBZlChr3sjsE
opfNxRz6fraNOWZZq2wXZcNlbNG1uweW1h+eN7WiCszzbMl3LXLGPZnhzixHyH8BxolPyl3pYTsh
s4OTiOGkt+ExUl+2ejpk7gir0o6S9SYtM3KzGnyxT8csb6KOBtt7dvLakVkYcbUS33f3IpnNgNGT
pL1cIOdDDoFNZgKbtRxO4DccxsQaStFIWY1n1hOEr3we/gJBSgRa1OeFigIGGS1ReOzMuCQqIK4A
gwKIjQw4hPPjwpX5xu1DkxRqj5gf9d8lGc5pnure7t55f4XJqHu78le7V26H/6SUIUdK5kEZFwEK
9FGM9sI6wdMmig53ENsB67hDclvIF/2L0QsO6VxX6venZRZjcVFvEi+iJxFkO0XN3jlMSfVTpWKC
YbCZwcYYkbu+9juYHtqDTu8jOA628vc4p4jHLcX4iq/Y6Qo+l4dAg546lfjjvuuSRCOFvfKgjBbk
m8absHo6pfju0mdVQzshNRaUXu9eGt67C4nc4aHVdvk6DunBzwZHNIUwh8yoyMXKkk99Ch3faKEl
en+Tl/5Gjs5bT/ZYiYvHU/B1lohM9H6jF/UP8Nc7XUI5Jc3DmI9qWn6N9H/e0ZF17mEjmyBMr//V
2Fgb5uyBrmF6QdwciHFqaCxv3IOjPimewjsj/omNGVa2rqq5gk1SsjpKunLCgRdWt0gBPvC/EE4J
gvG+j3D986gJv6Rpp6/DEnJZSLoj8rbg2ZLZwil/MxeDz0EvlF5nleU7UtDNlE8PSROMrABGCBdq
z9is+rUa/Ey8kRV5NQK4KZQdmoyMMau379hN1QY+sIH/05YGVjjZR8otC3z5nRMMBzQYFH8fCA9u
H8hSC+/Yxe2geSoZmkYcZscFTep/btkmfbATxPIDAVlv5Q3S1su9akNCi9lSYRmqG+pZv5e2YjD/
OAKptTYmkrfkwxN888ijgZQWgCcRwmrz5M5V2SSnbhLMqjkOFyetzv647Wo//kSEG/wUrrZUEIH4
LeeuAhZeGMZjib7MZzhgeCaf91vxbcgTScu1IbjUBBjsyr/KaY8/UhhpA1fVbwjRVOF+gLsWg+qz
umKW+gJoSYteAgBdu3IIv+mm6emaTOMKcY4A5q6kCf2pC5zuZfIgzN7qDPa5KIFplCLMWKY91fqz
BEQPVYGrYZ9Q5Yyh3yjN1Jubz4eMJZRl0t5PTxbsFKZ5tHZL+z29S2on6Fp3QdT5Md9fdDgfxiSu
f0Bi/kZFaSVEtNp30uWTZjHoUyzzKbY30QilI6zS5OINgDYA0YmGrNRO4eclIgGU663IKWcKiRmK
3IZV/OMiDqWAwRMK4dItL1DahIED/94vmatJWHwewUXg1gGwGu5saUOeUIucjIuDJiuxnyYtVokY
H7pyVaEq41GrVD+QsL2NxrGikYcdjnftMDp+10BW7JUoiRfZTuXeBR79h73yJh37xPr1e7HJvNAN
vr2sCJsvH3yiXtxVuyEJeW6++BPd+5Ul04x1W7S+0hnVjAlfqalJdOUHR7qQdn2NqTpCyV1MYSAX
VbCqwNGL3wxpfMmQjx2k1EsNBcHaXw4eunv0rrlTxEAlVnb9xzRIZeZrx1m5VHghrV2nwOx9aZFi
d0x/5wxS6f83A9TMsnLs2eeBrT/GpMqyqlmxLL0vejLV5wVIwJA4w9U4dAtGr1tCiwxm6I9V0NrK
9fxHKiEQAJoz0X5Tn6kZH5psWb1g+BzWSOvRU2rp2bvyST9ye0GAGvdj4Jsjvge/Yy8b2MOWeAKB
rvtPUdLE8zXtL4e546jQW2oXVyS+4AfoyOfBErpNr5LoK4Baiw0mtAE4PCEBDPY0tb474E6Lg3ra
rJNaVL/+DH9w14Snx/0SvwdRIcH/MX2pZXbgHzaEkcYUuJvtzWt1ZfnWtMSMEE2v/7lrGBbQ5sh5
6j05SK6AHGMAxRc7hEGIvOyN9dgvcpvQpJsu3lc7/4YSkDq+FJcFDLgYbzy6D1Ey9wMIlsBiwdRF
weZAN2XlwGWjOS1Cri3O9FfYikO239wlhivkXGkycnRIzIEruDdJdxbVpA+2re/ZLzYjlrjdwlQv
hTO9nPlZY13Cvmt1THY8kqbam2xVo1nVXJJiHpXoTUFqMgyMV6Lqc4G3W0XMRsq7DTOvxr+ne8IB
uavgQO9V2B56EP/XrADf9O5JLnSm1yhGBKj+e1pNHOrVYYSm6oAAIZWZfD+/HrhRwpex5GvWU53L
uJhfeHkA6AM3yg2fbDE4Zj/fzZDCtJZUHVroVe1iExz3LHPoTS2P9LImK4Vsp6PLe9lwo9O1mSGY
mDvHZafzlwELibg+jfG3JRiyagNNsBlBdKHsLsX+IRcRsrr5qV9xVAQTGhYlLqwBHnbNsnh8sS/1
sLUxw0dyZALm/++ExZQ8Z97qzh4HHOEEJMH4//ouWZGN6x3eARBFtmTToOjQiWzFm3uGh/TBbAVh
RbCdmYh2BYVFoyS74S58Xk/uYu0A3v4h+y8IhRFHJ/mV4dQCWcu5MzkUFqaBnjOBU7YsPzZWz/cm
/OiA3NhMfY2Z2HmZgdTka2ZbKVQea7ysksw8IFTu9Iz7B8xHvkq3SMB1vUIIRRhil/GLkZcm2acB
n39IpTCFHvVJx7Sjzs9dSXTXn/WJIkD4quBbnYwXYkKjeIguaQ8vSozEsYGv5GMCOaqOwsGldmoB
l5J1uffjSIi7Z8XozFaV1SeDtwJa9fRX5R1XvgenZTVY62BlPWRrbdAg1vb49HySiJt1PFVx+WMH
CFVyg97RpAdo/K0BEXK0gjSAMpau5y5aEMXIybSz69ssvSvcla7qKVEYvrGTK62RZI3++RsOlvKG
376W+xtbwsmvd8zC+8dpyWbZ3RUShPQS9TrfCiaVkoZJ7MQ2Q22bHjmFZO92nE2xn0qLA4CHLDDg
EqC3xtY6fiVKF6nuP2DTqGX4+mQv6KZAL/xeZhBQLCKM/DBzxycK+rlxyNBTcMB7qgsPgw32a283
qw5PAGG2wPz6AY7ywXX8LcXtOI+NnThTcLLNUrOzajbGxfBVHaT/fJNaZj4c28umGJvJSe6+KZvU
KqmxG6yqkW05ic+FQnBYB22ZHRqpFa8K/4YRnxmc/LxA7mujCzDZpDoxTg+d0I7qFIEfYOUF0BnL
434neXEuZjQW6TwBM9rdNBnI63qG1mH8ZcL8215WHtGyAqPw4h4p8spZ5fB70g5uBClFaUA8xZdT
Lfd1r/OFhpiYi8UXdeTsNW3N+tMTV6iQFCDQ9StTLFwIG7nAIhnaPAg9bDle+223WJaonLz1uPrZ
83qqaK+SjxlpNld3T737+m0EmtIZvd3cP+VCh8WPozOWkwVi/dUlZnRsXWkRY0MdJsQnZ9tZDjRX
AMi8v5EI3ZliWBVP5ZikJji/Ida4Z9S2Kle1RgXctvwwVFNAYspPSIY92Pzg8wyCu/cX1+oObvFl
tJN8V5T2vISKYu9QnnXjiOT7OteEplaB6vtqj7sVb6Ho0U6oy+J+O01bs48xuhoYr66MsOJnOvJu
x+r14kxeFC+Si1RI54IG/dei0mVmP4H4Dw6hk4RTy9zXMGvs+lpLGSU30hNq/Adxi+Hf47ihu8vK
FHGIR9vlaBtEL1+ZPZSm1bI3ZSwleXy7Zg647Tu77wFldSELlrR0vqURMFSw5I6vVD+Hty5gikNa
u037rtranlw6waK4MOf4OrsjlaPFAd4z7sQ9E3mFCQAyr5y39Zclvtw26Yw6MpmZiKPpEQxWGWNd
OHLZJ1oKwqZv/GSHPQzxzlSP+hHAscUWgyKnmK+jy53Ow9BrmhOLZdI5g6hoGReZvx61gB9K0gyS
jvhsbXwjhg3r5E/xetExPRacqdwajVBm6QAusndk1P5rjJeqCLuGewnsE0lTCiQIrXuJ3oNjAyJ4
787d3pLEbnlWaN2CYsh1AylT2ACtw0Afkdi/YWEqTEzJuS5vTxVufYggkw+vRGREBdS4BIEGgGrp
HrsviIm/MRpJNP3IEsH+i+83onrkmKhBxR82wnTZ9Hhv7cn6Ox9h3k+wLNL4hbZNILoTiqH6FAVm
0/lizAh3+3saMiXAecc5w4dW6BBd86DpwqihzvubgdcCMtZtiQbcdb6PcxI9M0hSs6daHu1Fa9i6
kMLy0OAnOEy3IYpkd0LRIBsjjwxdVsUmHI5vvgnjdJ+pfYSrPVETm07Xgy6zUdyUruxz8S3Cuwiq
UB8Ot4lqKns9ZRgcpOu4vMLut5awpZupKkl3TZUXhS9KtSbKrqchIMxgvmcBFvhDi4ZE5VJDNwCT
A429Q5PoVXgzl3lg/aaxjZArWpWqMrK0xiallW92kcFsIlirWhF7EC7v/3vuV9iTdnhA4wwz7+/i
d2mwxEoeNLvLhvp39uGNZD8eRugNImhantM6awnuG1RmMxCRbGnp4wkv/GQmdW6pZPKj26VP4K+u
vUi9HbEPdu+DfozMx8IVUUFWkvlk/dTsh4cYYdDyML7sfvoAcm9dZhdoVGq/Kvs5srq8xeh4q/3h
yCvfUz63/I8MqVbfxSYrtj8i8ZdQCuZ3bZy5W6Z8+bEFArbuwvx1HwGkHQzvGsZwyZMOjlve+HrD
tTQsdWEMvLOBBWjHdU1KHjn3g31X2NSgJ0DWVc6Wm2ZLdh32INuKFmnuOk2ApHsFuUBOgNQoB17/
AlIhce3+XJnTqnWwlI5I0uNCe1sDzJEhRTUD2lIAUsBmJQrDlDFUK2eGebUOc/G2eCTNWlUh9jQd
vTg40j/CecjlC9p9WDHpJAUqSEb37MS/WJ6qU2549a39irDJbALECDlWGJFIvvKjPJ69itZbKlYq
GPdk+1t2CXkmxKflHH3/vSIGdpLWTH6nq8boeZQH/JQcMTGc/KNsBOTrGytNP9RsXN5bCevfbPbv
cT+E986BCv46/ziZ+kkPvxAek5Svfosv87Z8EbNVj3PcrNH5Z0czUYoYpv8q+ouCHJKo36tkIrr/
zAv1wz3ELT/Aa5sJ2F1xXkyMYQTNl/LeT7vjX8pT2QhNC2/1h1nRbQy4XTKy8rM7aQIpRT/SXBBG
8ek/aXl+AQ+dlUpf6WKOBiwuNCS1jWvvB5CdH49CdIlN4pAJItrwDhu/XsSeQ63u0mHNRtzNrdVy
MyCRFgrpehi2yIC7kiEZkRw9yIOzkqYKEjrnOsN9fnckWq+6GQaKyJXmjb+X0Gaixi2kD4VqiW7V
MOzygCB61AuUlngp2oevDeA/RpPTuH9Cuo8CRM/baxbMSnNyckg3VaJp+5I1Jwsgcm4T7ln/ghgG
leB2dBS/xDEkeQA+OblPIOFTI9A85z/Itn4NNaHkV0Ax7OZ1G4bcTTRgngN6IKAq+6eYaausm2Kp
wXskaCfHmugdXD2TMBRIh7q3KgBAQMrrGZhSgkqeehw0kAESqEXu5ULXJrDR/p+zD85BFkO+QgeE
9YJrn79Z8qbChbLYu5c+bS4HPtfZkjAQVedNyK3o3MFDMAUX207XMMoqoSbihjutWBgT5Vr9v/Zf
sruVCYIoPzWM9EaBZQELryqlDIhF+qB6H7IZm+LDxRYESdwWNyZ6hF2nMEfBFvqgWIwJCvVeSKat
UspoBKTcPfWQix5BPr/EJkukvFXTG3J49nET7uMTa9vxaDRRgrJZnCH63o4eWlmZFzHy5YccFFIb
VbAGFggIci+ZCa4uYdM+NnuOehzv8mbdZo03hVd8dk1h5vgu1MukB4WpJFJ1eM8nxDGQE3Bn890A
HddhSVskReupJeWdyJd6M+RhbwKS59kxUhMXoajWxQRimonIId2Daa+fp3iQE0Mhv0LFtv5UyaiY
fEPO6h7Akq285PB9Da5FpkHjrnK+RNHUFABGg7MSCPA1KILg8thVBZW9CTP7RXIGKETrpSzk8DDE
FfeBoAvfaeJ1Bb/xF3m51U80K49a/MG1ZFkHI9np4HqY8uXFq7mkCeHX0CcTVhguSeG5+S2MyZEd
Be21p7FaeLDdMumQgtA2z6GLb+IORpivHKZEafCnOGneEC5WWqUZzDyoEa4oN0hBtq1NZ/iI0mRl
j8fPSWKOfVXJRkqV+Ay4ZK6ykou93dPIxwbOGrFpjmZkcCTHZ3JTn0+9VtCSXhcD/Vcx+ENDjXZJ
H+s65pUKgxXNSSk6qEDT2CO4XmwFdg95Xt3VcYYPpYkoX7P8B0KjX3bICirH0ZJfK072Ae8iCUqN
LSiOY/JXT/pH6h809yN18bvsrELhYTlVNAfyE/mQzgg6ipgc8AdMstL01Y8mmzqZRToMjLi4v3YD
TOwo/F3OWN/qLp3B+kFf6gLHR4qk58y+VRBs3Q2RHj95Hogh0xl0hHmYi9pEh0rfb2p9wgBK6hGy
hYNAEsTabwAsD6Dv+rAasDva+pff4QZy1EFi3VJ3PmhQr1nHHgqOgxfwRe7PjmYZpl4xEBRuDEmi
e96wPugtZEogWR71oGVUuvtLt2vRjUfAXPARRYPYP5tmX/LRn+xE3+NN5gionunFJXFvBup51pqy
hWjq08cl/Y8vJMlraLkPyp6qf+UkgykvJ1tntFTIcmQIvYrG2G+o/mh3rW3gfIgaYS2F9cAIKH/F
zC34kibA2kRz0u57X3Y7egfZlQMbM4U6n0E9AqbGaFSoPdgWh00jg/HnA2FHeI0YTJAZ3KjBcjET
qrWyoD+y72ispX/IiU48FLh0MX7cfLC/vpQFJKTCjvKWT1zxl1o2lOZBjW4wFQvtKRNtNuJyi+1P
ROp+WKCbHaSWpRw0bUErNVuXFNLwhCXx6Cbyo7/3IUane9y+co0lrl39l5dqCJfj0SD0HvYliBtF
i6s44Apnxn+hytoH/z3tR23eMBlpH149D3uhkiBUM2XNiZ5Ep9XIp45XaoxZTVG0OqVVlLkl6OV6
FMtia0E4Ug0MivaFxNy5VBRUMb6gQOL9I4avBZqgE94hND1vm3jA/fmzhpwhVRGBS1TDAf15I2vI
rQbvtXKv6Hq8NYwJNm/biDXrqinvIqW6WWl2wwETGLPVE/35LZek9ET8UiQRwcJzuIwnhNdiuI+2
cfkiHT8RXzirPgshc5Iw5x1ofYjlGa9DFuxJxTqAT1yoxymNkMkTwRT5lCrP8xcj6oTbv+/bx3Jv
/mMUjyNeANWFeToh4/bpSYC8XPsvx9SKObjEamE6xUmC5mvmsyHoDTOYgJs7hDbbHXAAXARD+1AN
aqLJqmNY1oOdM5NgaA2pVm5f666Yy2c49ttFaw4eL30Tz7x3W+bDp0HgUe0OXUdVNBoxeu8SsvPV
PA6NkLwF92bOATrb7GbZy+U45JdhFhGrfRZdqI/xah5ndrVV7RcePsA/vMjCnihnIxXRrfWNtDel
53LknqobQAFIdoUDy16OFJy8gwX9+8+qY2AlvsxWiRwdi/KHALRDtqR3C0CQvfJjiZ9ceR21c19y
Rj60UaU5O3eB2UO5mTSmyxWjnUax8wr/k+eAspOUaaofJPjAn26LF9pztkp3roCfnwleEIoaob63
xV58TWcUjzoKC/BKoKlYCo1F/r0/Kx1HEE0a+1/8Le5l86EAEuNZVxsdtThykWx+QKotJ7HJh+Ta
SyuL6vr4UwNhMU9MoDfqwE5eZD1ixoc6O1BODRIF7V0gMnY9WCJxHhFZ3dfDg6dvLldgCXltIQbg
iaK8Evl/9e5AbcMUt5nmFqz3HiNd0YEOKE8ZvXFox1iw2Qv0QRE2OfQWouTy0GuoX8GMYPVSmrvh
NbfhA8mU7m7Gew0R03MZJM7ctsHf411D3lXPZgIYC2r1LhoXupK2nVhom4q0AKRchwO2TWlLoDOk
ZUKgsapIhTamP3qW3rE9A+i42u5U80/ULt68bHjquyAuo5nCCK7c3Fx7RGuC87Kb+jEho/Qua0oZ
uHra7G1Nta9I1kcASAvQ6bH1ZLoo29qv9hFJjAuM5aTDbMAF3vKJS0h9QATv/oj4fmnticRvTFl8
bg4Tya1XHTxm16HYXtbY6A7iTn96BFdZ+9sSz9pPJ4brd0bga+RyjuKZmht3ARM2babGzwMJ+k9Q
Br36H7D8D4/JozhG0p3y5LXRDniZq/PwozpBsOQu8uPi8A5U7bWF7rBWGrpnRYpFKZAjtLZLCijL
QknJQyrDTfAsl4fVhvBxHh4i2d5qXvtg4Q1/dSq658RNwkBz+5uJCDTuCyunHl6ZhfNQVQ1sHUwf
/0GXw6LMkUQXVbGTRCcl6IFfr4JtCZS4Eed6XedN09wI3J6QoUpgd8oiA9tNgsWwb+Wk3lh7oeH3
y/mGX1hYervTXJGKQMZR/p4P3/cczZ/Bgdo474q2BKccuX4lz9QhWeDfJsWYsHsZX/iTPLrXl6dg
33Xnn2KuGRsKpLXQRW4ny80/ViX/2OYEelUzqHp3ZT6SIDom4VgCg5GKmIMZGum1NwTtewBc37sK
va1/aVQFMJiBXDSuQLq3yIxAMG9JueYtrkSplqlV4Q96REkcxWcbBBy2GW7O1lV9be5wfhZvIIbx
7tsk0w3LBdr5z1APZeQfNkFgkDiPdE+SOtw9EFPC39PKcNSy28S+afmM63txmI/e8T9rIGwSWDSQ
gADQYR0q5Ibunr1UwudlWl3s+MZkxT4F4tzxktlNeqX+uTIRZmctzTLHM/l74BKWLBlQAmxf3wyn
GTR+rTREa4+ahVJ9CW5Cg6UqfE/ZTFFriMP/btnbClrrKX9SL5OTXAARgeXPL133vT0frjiq1sNI
7S0vnTFptSxvAO/z/Qt2rtwFd/S12tiqNaSLQFQL71KzZZrHExmbTxJp06F3H1OssXtGkzHojDc4
FW6ZHqaHqkv8UwlbLWI4d37m5j+TJOgHtu2SpGG336k8ogOTH5v4mkZxe44fNVmVXAOuMFGlgAHd
ZfSQCxHZsqUJuQF7Yc95fogIKWeRlVK2rbK8hKCpRIoR4YEFWfJYpcAwswUMbYQxOZIUowEmGm6J
Jq8e4rEcIHSSxwtvzwUhVXQZ2KoYUWYy24bhhAVji2/nqtBhvJbPWT258g/T1Gm6ISEDrpc98/H6
mT/RAqQL0yyuxLB5+vehRHVrmumoCq57pJaa2Xtbp2W35JG3kqAEN1aou/KB40yW4j+C89KiRwob
Ovzh08rSQZv2KijAqJpDpDvrEcMWLVR1YNy1b0foz51I5noAYHlaPws2t/UzTk8Vzgj+gn7Feggq
FD+XdFvcKq37XdY6e0kzSuq4VlVk5A0KSBUReJQxQYJO4xV2glHA67aCI3w7teO0NMbuTwmPPrEc
oTuK/Up4Y1ImEhiZy6PoVU0fOYHSHZ3JCd7G0cNXZf2p0VF2+sxEWTdpmsZMAPuBAFWXpRzPQrno
7w4o4FYtVmQkB751L8iLHd1klj2uUzQA7r7iLieENa3NPEQAvmO/ZxnZlu1QGbW2ZyvydE2ji9m2
bdlCSB4PGFkC/abg4awRrTN2i+8TsqP25DjL/j+Aet0o4aB5gFrtHtzlIwALykttbMg0v/F667kC
SgyNjsgXdluFiVO2dOqtdx1Fwq3L1DPao/hd30yAIEZOgF1VHvuvqrQmuaOaOOx/ujffKv9C5bI5
5qlqPUp5UjDKM2ARkyhF5EDzmfsurvnnkPTDiBiS0OiuTuQGvSkrUaxPTfZW3GlufA+xrqqnBRcA
WXIB45XnEF9XH9OTWzraLFAVP4wki8IA7GdxTGvBuBrDF+ewX7fnIovJXyaG+CGo98/BxN58a+C6
iMhqv5TpZdUNsCj2oqxFh1xOxclXYhx+Ok/kyl2p8qP67p1wYjIdLV3TLgdHsuEdDqZkyf4WPINh
B5VMAbm7VZj5WozSdvN96bfFxsivX6wny4QNZF5KvnrPuRfgOZVrHSsuhm1eFsgzcj+2MT0coTY4
S2MAx1J0TFr9fGFUQ/bDzaDRk/GMNSalBZqnb9TOgc1NSqIHGy6tPGL+Ui5BZDmDgT6N5tf1bt2w
Q+5Fwr+asiCM2WVzeJReDKPpFjP0z+JizefVS//IdD/XF2Vq7UHdRT1U9XPqEQwiApkxXsduRkwN
Rto1XbTP4vIxxbrKnMCdrgaUYrCrPrt4X9QzP4vq/4yqb7AoX4XoHYfKSeAZVlJX9YnFfJc9d8+Z
egQEmwyqOH7pf3XH65jw3Y0D5sdb8EZLW3xKOT1J2D8C0lLN0g1W628DDJq4plORTetAgr+WZwbi
q2aeT5UwePriKaW42yqXxAvDYqDyiYWoYau/DuVsRRN4uBnhUbjpMw5CXjZzWDE0S4X/qpGzbvH+
mWbzhLw7J+Dg+BqKlzg+NwZ4H200Wffv778ExU8cGQIRl1IdcRgIu6J7JhiN783WNWEiCH3QRCUm
z5qeqZ6ByHIqhXvImMBhCE6UcgpgEoJJ8DiyKjFR/q4gO0WZIgJwLkXOIpx8Iv+dKuImE2UJrNnC
tiZpUY2cAmkjlBXY8j2HqskL0wmjDnnN6c6XKhymw03BTQWWkQhShJ3kV+fID/lZsigsM7BU5y1R
KoZzq98yoxacpTO2CLoQyVU6OjyzzB0KSN/fgsEWI2GWwU0MSSqCok4HDsQDj90/8I83VY8HVmfu
mE7PT8r7HKSu+1cBpDkxj1NFOqHjJZqo4W5B5bJErvGC5aCJoGcbM3UQ6CEQXB4WhWZq1yFCzBnb
GNnkvv71LwiVAi+knREx6Sfv4TPP9uyNTyJzogS+FQcXXta4tZbr03WoXPdgzg/PJ5eOEtB+rJqg
vhqTyJ29eeUnv9+ugs6yzMml0sfI3aK9kgEPJqoY1sMeD1jVjIv0EviM5OpzDKDhHUTXH3W0px7N
T9nINC8FBV/R1LHXSCeFgj9tkh915zlNBsQHa2JQFLhFKC3xfWMqkEK1rZLrD6xADKCD0l8uGL9E
Jfnfs2xAtcfFm5HAk/8lYgohLYPyHf6uUTkpQ1/fV+pOuFt4HbCppslWF//zG//avLThDi0Qj0tY
zhMKMKSi+Gl9Z4jqzHdudrYUGPF790zYQSAsoAhpBwBZs2t2qPT6eY636IPQ5SSjnrZUpSSpq2YU
XP51hCIGewBrJ6LFUkQKOQd2zuAsW4yVd8ErnPQPHPlagZKQ/+6xDkcZP6FkJu+ii9L/nRoKo87J
BS9YIixXLNBnmIl2mlI5e+PAIUxMGbo7SZJhh3g2v6EnSJGFLzhhlO5ZS1hHU5Dvp0uhIBulBLwB
qgobeTZGuxdp8fWXq9isOOP9snOYkIWjZUhEiX863bNIVhOZLhURQNHpAJXvi7gHZBftcYNRnBAO
u7tyJaHhqcCArQCav63OPVibjiZdY7P6uvcVvKBYDGJ38w2UmheR4h0pMd3KHLONbOELJu0C0N+e
f8DWLpBQIwPp4DCi5Nt3GUH2kPVOoEWhDIYyE6Fg1tae6eie5B6MjzO6sR0TG2/tPAB1GGY/7v5d
3AuQHVZ6sdjAuSOFzb83iBvH5Ds/h50i1AuZFEPHFLvZHh64NxRcnWPH5hW2zZ8Mjnu+1sVzAD5S
7Wi6uMF874pT5uQTtsVaRYzFV7M7uePYT2of4/NlY2SlG81mv0Q86iOjxX6/URScOBvKgs6IIPGz
12ArCWyCYiqsxEyIWYOBO7WyWxuis8HhxlBThR4UhL8m/C6GGTt0XvnPnbYXa11Ci9c+QA2NA2Th
NwVALFaQm7JPuX0uU4IXCKFyVObqL4ClLrqFBJIlLDjlMVhcrXum8BPOgbnFkyVCEtWgGYt6z5vK
E6VgTSs7xNwKPibAgnYJtis4DjuLmaftRsPkaC+3UCVCiz4jHk/hlVzThUZajs/gH5tHLbBQ4CsN
6kQjMj/sX/h6xFT5KNpPPt5sV7U3aoPX0+/FugqC1aThRC+3bu3z6QeMEQCdzrYm2kzH8lYKYC7N
cNm3sakjZMQB/WEYbNPbHLZnWL7OShumm8uz5R9gEUv/sIsydDRuBPfCQoOa5SoJDOl55PycVM6k
YBloqdwAP+hOV9H/IGwTuZukch+fzpnwcfBcWY5353yrQ4ekhtefu9LSp7TlS4Pd3EE/vzpvnn6s
dpK0nd7xvJ3Nc7xd/t+kUI5fiqAN0+hOFrVmDJQm3Ky/LRxaB2hd0/X4V6EFHY76YOBm8Pg502z0
d83mZzQ7LSt5c1Ixx8IB5CxDRZDOzwlkbP2rHoEm8m6fyAZ8mDvwaniYZYVR1o97Z9yOlAOM3r7N
tlAprK1dpDWaHaax7QTmGjgyjbwEfhvgAoD1SW72CNSI50XGTgPcM1RfecMnqJ2VLOiyONWK/SWJ
15eGZ0iiZZlncp6nKMr0eXtioc+Armhfbe/D+ASioenEnbu8CsC6t6NmK8h63IuibZKJqo1qPkY1
mXNFiY5fTSKBHemcQhnTt0PgeUKRiai9NzL94GIqNwQOv/tcNOaLGYWi0gujka0VgOzQSQEBxW0J
J0G6w5DnFdvIq8TmaIf8Ik5oMBYEGW0sG5ZMTIg74DxUzOrD8rvs0Oex1Id2lLJpbJmC+9wUTekn
XUz8j6cCVf8XzW5q6Hf/n/K6KXyYkSOZpd+ZawSz4rL4zFtdkI5cA2SVbMQWPIWnhONHenbTQa8J
HJXH0BBJ+24ShlPgqvvSCF/6wXoOnNxbv3NgppteuSbp8rwn1DcwlgxlnByBxLqK8j5GFkTp5W8I
M+1iTCHJ/vktWbDSjc5eYzYdNIKetvX1MhHBmYa2mJVFOgF+yOwrpqiN+dLgc8FVQY4vSbgildhR
hZcF8pvG2cIuwpZsu+4/S+CE3zPG3PKTjOWvCESmOHnKeBTmxJlyTUfbuFMFo3h0mq7OKgFPLjN7
sckVoLoK54J2JLN1qugimQkKsO9uuW+WZ6wlBH1ePuF//HbP3fI0GT31YNRf2TSGfdMRXZiZXSez
0+GWvO94x1Owxl2UzAy1S1XF5nijIIjxaR8nodhUrpzBXNCMmHp6VMNauuS7KYYeePnik6D4FyKR
ARloScutaJx/jtjIhW6oDHBDI0FQBP5YKusfLsfZZ3KHpdudkoOJQ4P3eAwx6R7Gdr+b2Z+Kcfbe
8tFbDE4ZwdkoseQiAAasrtYKze/6cbHvQySkrRMf1pIj5zg8XQ2mZldtoa7pXbYzoeQukN4tN8p5
0fGbwOyEFXM3mHD4jcVSizkAhaVdSd1FC2QrWPTxf47hfUvkJ0u1HlMHh+E4pajgwstfbccbRpM4
xwtoul3jnuwv3xAIKqxtInCKV3jfrZTdUF33TsGUp5gsA1stAfTQnmF2aHqiGo1ntfsbqpX0jH8I
vbMlKA1CX/GUgG5ZfbfsMh2RSZCIjpidDlp+xw4Y45Q2up0Kd9u1xZmFx5Qby2Imt5ALeBMu73/a
aoG2e9elblX03eBkOmtktLlOZM1JPvWa6P1pX6xlciuckr93gJ5VUdI/uvlxtzFsVz/n3s0yCq4s
vtzilHqol4RhJfLo8e48c0yYIgKFoH2MXltlx73pCHquaLx/f+6lZigjnaE0fj4lg/w3zJXzx6kX
Ruo2biolYn96z/uXzLU7pe8sKzXQKwPK6e7QVKpD2UlL0CrKj2AFibXCKiQcrLzL9kjTuzcaQsQj
UfXk2aMHoXIPECV8reoU25TP1jyZlSvtUIDZNIVd3NkRtrwnWG3qWk/OuFpVsJ7RW0eHUH+oZ1Ab
zbZutaEuBGssiV8VidKmrE9M7WQxA6XkxH85lQu2MRIeOKxn7sCkmPQ3bCrmIwpBL0o0X1sYuP3Q
rrorK7OF4h6YXi6hmNO3cr6hpNK+7HbIOI95RjnsWBbmVPPfGme8kDAAwaqOhogiEfbgXh+qlrOu
AlaUuxHHwmqwybiSK/ef+AqPHPM1hYDwuePyfjWy2xCrwebasF4YnR8a3c2uqLMmxjBJI4JAaMiu
RhMgqCWnfltRyxw0mTQKOwdSF8CdrBvTVER+lug8xJysOkTbmMvWdRYxZoKwxO6NZ5Dpmcw6gmGu
CsPfSwxyhdJ5DkHMHZzN4rf7Uy5/nblh+CEJQwO0UYaOsKoivCPv/e3vpoxHBn9Eg/yBXE78lgDL
viZ5a5UI5loB6zvuDS3+j0/cpWVGE43qRjIgsvIgJ25jWFOFqWN8hNTSS2HtUepHQryeI4bOVnnH
XCCrHOBY2ojghBLjHHS7oXgJqmjeSWCvKI1fSIM4xABDXBBPvaGvkTMhpS8demDIROZRYKGGZ1oe
SXSDTEX6hI4uq5KyF4lrsY6PPs7OM0atscZCv14tsg7d7qysl0NXCsFUM067Lg2eX5Vu7eXqtXJA
S5crGguzRJ2biWoXZPQZz86VmgcgxtP4wbDvFIobod7EFHtwDKlNNv3wb3L4pNgT83lqd1LUIwIw
Di7gWs6kQa3biAaMCMh9ZjjvMAWxKaSg0BxZviaOf/SI3vEF42IkbCzvps9XJrnhKrYIIuxFYbDK
4awNMg90OvJSaUuCTK06tIsIeU3H3bWVTtY9tahNA65h1cCeAWJjoNoyY2vPcBgptBVs7ffjsxjX
UrsDut/Oc3pt0fx+WxibJ4PfbfPVWBsAcLKIw7jXa7xfB2Qn3lGpkDQpVTKrzAfFmzdFXvF+Gibc
2UuncRnUDkpBE7yecPU1dlcEG+761z6E0bK+OAjxhSEcbTB4kUd5Oy3y1Eanrx6/RNqd8AnElPIN
ncB+xefLPJMSfX6xccr7Fdmc9KaJe0jssVmYcV9aAYn2wdXMpRhl0s9tav5R9z3lOSex40Kv3snn
2BRYRHJYwDB2NaMrwhIzMRjl75Z2taaJDVlR9KbVe+XUwBcgWZPEwQmlvzJzUg30pG/O0jZvtRit
h4xlhCn3hzQZQqDJT50jH1iCrLeM0WBQptWqn0qftzWViFu86+lVQzKYH0XJb/gO9R5QyUUvghzq
E4gEZ+NvjwAkPXLR1cBEzYRwHemS9+y9xd1c7E5JH+8+zw9LAGepTynrH+/55yOdAiKZINTDnLqm
SF717sy4hq/NtPbmhR6StHdYGzzyvWgKfpgzphr0U98N3Dpz+LPYIJILzGNcgqjeKPViVktJSb7Q
wcGueuWLmiEbG3HgvpjplDrwO+UL8hZ3ZCnxQ9iJW7jMx7ggDjnucojo9cQrnL3H/Vy45ZJOS5q6
nEPGpD3PJ+xtsVRDx5zR7YUUnjtY513tgESv+BB5ha+6ivs3HB4W07BA+hX37DWfgAK1UvETop3W
mYaQHlya/yRIm1+1Fw39FeNEixOTYU4FoeG9o+WeWco88AE8+jbgjoWeob5lohXzoZWU1J6+z/8W
U+j2iYNyQfRtjET65r8h94LBP2q8702J167DGiTg10S4Gfgrd/PQCRKdVDq0uCjSSKu6tvr8B1z+
M/g6dxoiB+bX/Oi1ai7Sf0zXTdhDZzalsTfiboOv8bgc4mruE6rN3Cs9CL1rnKVaj7PZ/Jb4eWLp
RJN2DF4GMxYCJPDfVZlCYUFnvupDHASC5IASLpUOL8Qm247RDbB30Kxynv8gj3sskyij25bVy+by
T2jSSUcW2+WQt0IY05CC9s5nO0wfOljjmlHQIh9sISIytbjnKIScLdPoPXn9EtldlDnKWHzItlT+
91IcHKGjJhtCrFTLaxX/gtv6ObL2PrY3lQXE7BmUeWE152DBJ6xTxslQtWtjJhpmtzRHd7TFOyNr
M7hQwfklX982B63oPo+2+LhDe0MyjynfzbITzreTSj/LDPgqks4Y3eG2R9Ix+lOKkZXA/nixAkVa
rh6d1qtP9deM4Mnny4soxubMfUdKTRpinWJo2u/5CnKM0lmKnpZTPKX+wNkcFEDfnqWXLno/q5EK
62CVad2GtvLErfjAQsAKXsG8iXNuHb0tcMoc12vfphe7BHJ2iREa8Trx312wC1eoE7XL+2XlIQoT
BQtkUTZpXkydVjRtmez4uB8hZXCc8Y/APTgHBCjcq7rnn8cPl4wDGINObQErmm2RU/gWZbzJo75o
dfAk3N4p2UlEqFYbh74r9oo4HW8hzg5jfi+YmBeT8XsFi4uIAekOYP3CnO6gCS6e8x8/wlDcjzb+
jKu1hgp0KQWL/DVXYyx/cJyYFUVdR8k2SVJYAakHOK3gZhDiB8Mdy8AdQShOxfWWBxHMxoDW0ESa
W2FJGK1q0PEdhc6wAyrltBZYb3KL58T5FrS8TdqMHU7oP/vh1kzPhn2wZuLKDoAZseTv7RrBgpBH
vT4Trgp7GzpFe/ecNs/jbu82NZernqsMbyXAqvSvL8RxKPtSCORIfDXeZ83+I5an7GLngQ9P+czi
F98yxr0Gzhz3zjD3pgguzr3+1BuTigXepMo1ZkDLtR9AsFWPt5hwxhXYYZVy+rQvGSZw2AKxLedm
6uxsgUPxQ6d3eQoSS+goelipuLagOzKoLpH4y4qQcnNNO86OzRPf/PzKiojCPJHgvxA/L35TAJ+J
RICLSbkCxzguBeEGafb5dMCMogI3sRNH5nnoxR126PG1yTx0XMwnYK5xBS6ls85kNJlICiIeVIFv
5notdV0Y7f1lBJVc5dMDPai58rCE8qtwaB4p2F/ZFeaF10w6Y9UbISVvYGQobBvOCK2Q6Jozgq8T
HTdkKFFfnsP82iTQmQMQoyN+xYV4guteD0ceUDr12VrEehaqEQyHsR0r0Pd+sDno6WZunAMdl7I5
U1rMNhQCG4GNPAKXfAgEu/vMFB/vStA+CH4uUnMnzFIAVWh7kTLLAKVBc8ih/FMDsYBiVzdohftb
G4BLeTQmeBqTZnLd6vgU/MKNzn90/hPaVps2aQ++6lRjoEw0Tjx2sQVFGv6QXE2v2pZJgZUOoKyu
rR5zoQHB3WzmF0KBRQMxUNKzPhjY5wyLhkK6Mdv6AZGe7JAJEr+4I0h+VG+yLEljeoJN/DNWUPMr
xarM/JdtrCLKEh5NOJgGKY3mwQoLF5vvPrTcQJCKABSRYDCOoJk+TUP5/WVo9/QeejmfpRHfPcGE
Ow4w8W9U639JvXWvUkuSIbUbu0MYLEwmJgitsDPidhtPuPaeGA8fnyYZq7P8Ijw89xXFijgN5puG
1P+DuDMAU+bUN9RSoL8VeoNZkWzPbxDZN2z2jkSu+t9nPIhA0keHyTNiCSF3wqH6H5Bd82x12Bjd
8ItM7zLcZBPx2VhLXLMu7Vxiz1BvEe+pCKAXGrGS7n8mMANiFj2hkQW/9ZZYgIIEtFHqmCvnF2MG
KUe2bt9VpCAAmPeURn24KbmLfDeUV2Clyoesk5D8NNy9LmRJp9mhSe8fAHGmf54/EDRgNVJHm/jB
jpakkOwBDiAC9Lo4B6OPKYZr3w7B2lem8dag3WSRVJfsILxvWexw7Rvi4grMOnYdp8Przx0MVfWf
fttIFuov4igbcqWBzABNCOIL6yGaWA7Qy8YJxdmS0/mE5iQ4MlfU3xucxgKhwZMKpgANXc+DmvmE
LFWwS2IkuwB9bOdgxSZfDSobuFqcBqWYL+BgeHEs9M74vcUyamTexHHFpMtTQfTejssy415yEK6Y
qkFPmpvgMWzW29WpRNnTJbYiYFfLxkaRr8Ahxu3HbVLTGEd4Wy86zFJXdGKEFUKI6Vb7XqyvNAff
wvWZcMGheNYHhI+XXEQbrBRRm6clvq3jbl5JzfL1eY6I9X/R5uXx+nudV84nnJLhqkvlEVNiLCZe
qytubCWNzkiJNv3yLjHJob6PyJHi1Qomr13YvBrlUUGdjvR5lm5U/nUcOjB9acHRdTx1j1pkxoeE
posXT6k11kpOXPDYGAFMUUbYfIp8p8zg11RzTlqe+T8CuFg6/cdfEAXpQ6edwNjHg3yuYjnhI9mH
5ObQljAKgAFInxaKqPtFnFFTrcGSZ1MIBDXDxRL6qicPEYew6GhPDZdpp01F8/GAq4zgbos7Pbts
1X85UYamu3/vRi73QZthMTanNoliL84wMJFykyBGoYR7GyqvcS0JhHtzd5TWXNzuKfjsFkgc4/lc
y5zUFFDfRa3L2u2DN4O1NWh3Oxl/En+wapnvZBzIhFmR6J8kZw3MQWBJdcE+phihB1dF/05RfghC
ntxoPp8sRMPInKXMZYaHOeXvoHD45wRM5UpZEEXl4W983EmbL/QZ0mLAYzCHolO5YhzwoLHi79YX
oytGtuLyMihH7YAla2MIxiN2FjlGreyMv+cu6dKqe8WrzMJIA1wOZkKtAs6+O8fnYWVa8hsd9IDL
Ls8yygo/k7dHoTrX/u9OBdYlahBWf3cPt8Qh2GvnVQk1PyaT8YI0QdXCIBc5803TKcwuHQWd1ded
/l+RYJaEPLwsdAQDWFdTIkTe7lx5+58yc4X9zgjU0GZEd41xHvPVjHbaDdded2ycGoUowlXndLNu
wIgW6ypRLEjGA72HVudNSilMeA22Piz/2gljZ85yAat1/PwRT7gh6ECXMouRGRuZKKC8RdCACIdx
RsXz/+LmeR1ozudAwZw0BKNB9X6GcnrGfru9IvED5N/xQu7umB8oTPkIIcxjW1W5xZ9nNg9bfIi9
Pf4EfA99mjqZ+CgCsrzlVOqt2ZzQNOPAm1gB6zMyH3ghPsM15TqUwtQvgGzZzUJK5JEwVMDPL3uQ
jiUeqJkZ962aneA1RlzHN3X04Yg88l8f7uTGdBF/UJHJxFH+qnfY6nuffqsfSOqp3r2Edu4ZTcEV
CgrMBSJUbBl3ir21aH7ndylyvxnrLDSKN3lDJw+dbyVnRQzw0HDIGa/s6AaWRpH4KJyNYU6EPIML
rvkDspUGqaFpyadItGLaZvJBYdpaNQMwZbD8+lVuZ1fA9UFQhe79e1k3dea5IDJWWMi/3JiT10Yp
9pq6uhvP8fq5Gzqeg0iJCRq5C154IfhSk0/GDidw7usUuraoDHGepsXyJTDSmBM0k8kLhZUrGSyl
vMs41urfFhZHe5S6sRMMeg9kCcsyR27a5Ibijjx5jfoMVCOTf/HlJWPKrXFcwUMj/kjZClWuhK4z
57toOlj67GfYaHLzHu+gg2Z2NG3WpIUnbQTCeo5W45OprSVTo9aqEH256FOGf/z9HsoP2Ms7AeqQ
JUwtibpvnfGq4SfRlEWVTsJdRAA6qU7yNIKHYP0ZOizGEGMBiJANZ4tpJFEQ7U89tTP4xzHR5hI2
2nu2JS/BE+YQREKTQqxKA4d8BFVrYj6NSsOGEFLrB9izelV33kewPvjcfCVWfJ3BREWCvX705OGy
PM2v1EaCrUPre6ONcSHzcOyPF/BnwdpGllyXB1K9s9btaOhIiHZU9yBc1XsAuAz/zHfQQ4AURV7z
HnEIrbOdhuTWBNY/b35rKRltYfuBbb2g6SRmabNYRreseISEdlX0337yoNwXrlvecN1tZVqYlI/o
87U2SKQpVU56KYTLXASWBojHe2r8t8oTjRrhmlcORWHadplmiorfX3dHWc0cl6RqWCYn6OdrE2Sh
QE3Sei+u39Ym96auRp9+mV4gizFMdUxKXiUOm0KK9Pwn+5tIIgtUa6YKt72i/qOqB8e/UZdrar/1
Zj4kzBvRtynnf2TC0s1TyJe7OPCvzZ6Mc7RRl3TXj6J3lNGQJIck10KiOlta2a7UlZy41/4f3qGz
ox9V8T7j+XxrMMXG+5M07/GnIsH5lPXHQBOmfl9yTYa4lMSybnhlU0l+c2pIPXFFjm0pOtNUwrdU
qGjtSEtlzwquwwRWyD5/0ntdSLjeQwU6Sfc6S6lbZy1ryNLpG0Aw7+1vJUgNpAlynP2ld8eozNbf
ybKCmPqwpHwYIgE9rqH09Zr72jzlYxoWttQytei4Jg0CkamLlCAW8dpK3Osxu8FYPsv/Gp6MfYcG
Gk+6sCH/TADmrBQXrTBNNi6tUkhRHKVCzwppkIH1SmlzA+Mt8oXSIzTdRSRWYY2h3PgH9oBqtYt5
GllT6MT9fynhijAXjbNXk3TqM63t83Z47h+YwpNv4q3FFthrJWqNtw8B+WlxhjFRpAjA2mjrcgaQ
0Txg1OAvICA/0hehEvjyrmq/7gjl9UbTLeK4nkgi1CInpU1x2cqNpnpw4yaAlD0j4UmDSo9Aml+p
a1Vs5bHgdCxgvNPjOnqJEdkX01j8zvzEOOzK/KvN+eYRymAvD+0j/1ReJmjjMsxTIwz6OH6R6UDd
r2cUS5u6m+JwdDnlDnOq5VHO67EQug1P3G7d6qQYzMFgIoEUcjdGeuqYuOYbjfeXgSA7R4RQtEaI
gXHW/Htg9XrWNjKUedFt+csspq0we+pmp8vyPNrB6C0vm9UJlhsU9+LtJ+7gNIWJn0U0tbbG6zwb
KL34Emh9EtkyyTOj3iFh0zA9FV3jh5iL16PhsVB3FF4PPzq3khg2rDrGgcBPWYHRvGLqqnIuF6v5
xVX1LO9bbvwVvOzHstm2m5Ib4haSWuISXd7TMpFZbtWRACSkNjK6IRlsPvFVUPuHWqwX58aPyYJC
bsEplGkSdVrPavzglY0c9kTwkm09Az3Lzoht0TTXeL7qlIT+VjwH9/DsrBtg6YakG1YkpFb2qhfa
6OLfZmsTgbB8tRStfAN+f/PzuOnMZFFd7W6sQepdCUeXPdwWBj83/79lewUkbpeVDywwOBmNITkA
LKn/0fIaN+eqwDPSqO2yBA5nwAdMNNYVlnqXAfoY5d9MJKU0Fu1mveIOoimJQveBDexhiYRZ9CEo
GAI1yFNH89l3pel26DU6EW2HaVaSklByKel+/Rsv+guvi5dIJPqsym7hZp7drgFBK+2NPXdtjkSJ
cEt5NeCJoKpAWv41eOBVhMkOKCjTxJuvyq7SgExoFrHus5niGUgzvElSS899+Cbejr6qIfd/XltO
/wZxWQJWIXa52+sRQmnIGF2z3j8uR7yBuKgK+NWlQEo2E1ztlvX4/o+LrLtjaqDVO0P6JKWLVSTG
CVDJ8jZZZdXo1SFVuq/QMBj9bx2229+g4+r/32t1fCxjZ9OFR9djrzdbu/WX1yIZ5BowcYc8Cojy
cUmT6qpcowkoudafU5d4dY67/aWGekCNMLlmSCt+XeC3o0p6QK1DxUGyVC+bq4oL+riK70hJSdHN
mK5gq2SjX3FKGQWlU6hZ+tLbOM5ZVjQX6NsWdhVH1Nu17ACi5ewEmkRsIVCbPkQB2nbqzZw30AXe
C/yxenlArwOpkAhFO0aGvAVXcsszd4Z/TGbthcBoPxHFXTMtfnwL1N5mXiwDKWvEhGE4XtKOLXOt
fa/jg9XKHgYzq4R/A3MitVcZbEJUU+ZkdMtqhM6SwW6mFvi1MH0FvkyCXmd5ctf4V145pcJkaY08
mDC53xRruo2GRjlbmpVI8f5TyM4KutqXyrzL4/tp1I4pcloqp9VuDEOQ1hl28P/911OOCql7LIxF
/m8Cb6U8IzGZcrVJQLT3PMOFqrMic+JaKKgFZypD5DzaNmE57hjw7h4YuFArbTNdqGihVOkGUhxn
SEftrFH3kq+VB+IfDobMU7pm0uZZ4I0M8XEfErlJgoMKZHr97UZcWWpiwHGt9QJ8v0H2zAlBLKV8
BPxZ8mibdxFKHhOyTJ6D66Qs8xF6TICPXHj2LacBiLnK1c+CgYmAfzcwOgoliExUgAKOPHkAvgPN
mJn3aAZ0Be+Yq6i6UqHE8omWirxSVwp0zygEKkk4TFTIRzGL/l9jIhdsLrhJt3JxnmFUY5sqFUCP
zU72g4tENrpK34jiOsbvl+LEdBETGtAcCbX6Kkr58V2IeFGHCChXQdcJ5Cc4W2YDXqQ2n65nwb6J
DWjiST7dlC8HWRNvPwnPlkf2LCJR+7gXsFRQ6ncXbq4tGRdn+CJM94CX9tMrJHnoQuSvtXHHqwkr
i0OBTxgjJ1e2jNdZm0DJsSoAYeUit8aqe0SLIBDE4ncOX9btntXvkWG4qTNmOX5fLEklcp7d46e1
7iFCFxmm1y07iSbyZ2ODjbkYs/RhghFuyEdRlt0tk/tGr3qe+PDmAob3NhLU+VGMDmYhHUXLn8og
vbbzH0t7s4uPG9mwn0oqAGiKjCnQ8x/FYnznlYup8Agyb5CSYh5CmDusCEt2q+4QCy/cVHA5ErmM
rCK04seZZp5l0I2IcI3z1574XC2TktSOQVRaQpPVSxgSp1QaWBf8q27DyxiLJm9R0yt4wT0gyQ+n
TwNY/hriIUotHxn5dErc4JjwS6zrnBp4ukwyqGlbkNyWvTtcfZU3HKWFBBQuer5u0TGwrceSFBli
uwR3YbAxNHIgsup57XZ/LaTM+rKh/q4O54iPWO0BFQIG9vSHLRvpAcDcd8tUQ6IydCRUQcyR5WKr
hrNqILYxhsI35umtQza5JUmxfmo0JRgiBBSgEYOnwiyvAb6YwcmvRORTkGcjJofpe1NS9/nT8DGv
FkkBLlxsaKDzQc1jO4PaC9PTGeU6pMsWdrQi/R/Bc98T2YIDUFgHPiqJn/ZDHcsNKTAsIsaj7olY
xwmGCLy9YadqoB3mOc9xPxIrsv6iNofCF8HM43slCz7lCRGW34grBON1GD7rRyg/WvdNjtQ+WbFL
nekZ0Hs0oG8/WJNiGiHI6m/ydmWFJAN0Krq4XAKmgG60mX6bkGtUN5ZRkOKrxfTEGwPuWKsgPZf5
6iAp4DZ2Rtsjx2HkoUhqH1/7WjjCqmXa2c8MZVExi4G/O4Ox2Aai6VMFTHRlK1MET5Ia0uLgyNvH
F7N1OFT/Elu/XIOcbbXPXy3r4wMMfWPqTu90Wq/mwv4wFFsPJt1fYzP/TYKeuiMSpaZQUegPx0Oa
sXyFAJYZ3NX2IqRjyXqWIW8c10D6p3w2EU2FMCm8WxYNi3NaV4M1YUiSDk/DRbNtMbuv2wqKUh/b
LnpX2kJkK8Kbj4OahVSgsiij/nhttgGtFJLObMsIE7mLeXgtU7rAM4kkaIIiNrWanIYSFBw5wjZO
4YzkifXQgpHptp5tSIYBoOVj9/wJrd1PCRw3avsezWO+iRbrljzjOCB4G1II/Wa/SiPqcjM6dUB7
at9HcP5Y6FuMyqZ3Kz900wxLpKhV/SuE3zlzgaNaS998dF5Qhoe7MfMZ8XVt5X3Nx8rDfduSmC3J
hLGN1AMFu4HAH3Nsk85Z5k56feKAx8V3hVJejVaSvO+G21SlPT9gyK/2cRFFXGffqLv/eI4KGZa9
j4EljNOO0L4jx+0gJvzwHGzJQsaz52a5GHYRNaOZgUmNbSkHj1pAsy6Lw2B3LXXW56FJLvyZOibx
LiaRWtbLfc8tRnjqbiiJ2P9fF0a2lss98G9fAlokifl6ZojEbMLhCAcletj4nypchcDO0q3IldNw
vPSgLG51UYvlrcC0vCyk4u6L4Vzf6BsB1Y6EZWarno9RMOdX1FLuvZsWu0icPeksKgPd2HpbEfhw
QKzoUNv6DLIcdgAJ6ZhS07kcv24Hq/3IP9HEesi2n47ziZ6cGiQUYzKdJpqalAJwPVOxx8xhA/zX
hQRDEIJ/kMy2gM+0QZWObuqzsrC/nD1JuMSNEPi2qxyH4UhNKo4cMKqEA+JFj2NKHynSMUgGWFVg
vhX+gXmzIAr4cgt9nxZ3lkYGAKZQtvPXtbIMyvmAF1crgMF59Lh5drAw7ilq0Hm07SK5q5lYza2s
m4F/l4FnEmsWqIu5fLjKDA/GklV1qCYxJNDCJRhbADyVYseDw9yvGKVYOtZAu6StAvUPGgScPuO2
4rKChlGsQ+as9DdpDvvtCZjeMA3so98y68EpjoFmusJsmdhyYILdqJpKy3SH+k4qr6bZf5fRytpy
Rm6+QCKW4OWhUfolKVTU4jmswxDnPcff8xiYRu00JJGZGjYe2XsBdyKQMfnejRgmMLdClugmRi6o
SxELQdlgjkkT/lAk5n+aFfKcIw9LlkodeM8q04Af7UpFOG1YJqQyb++FJ7dstEnUhTMiEkMAn+dE
3DiDjbTcqbKCzzAQGtbwyNab0BrTiO9SfAwopaRXXyuoAVMa+0s5F+dcC+CX6uomPdSr+xqv7TtZ
2rwJ+J91eD8yT13B44rhHHhG5Z/5S4Xn3cwwZxSkh5QkzCEvBjWwvsdjzZ9WiJceiJtf2E2ZK2P2
loyDbOaxVmjGnh4lbYtbGsUt8p3GrwChcyopbLgRouA3waL4UOix2U4pLr0JjKkpqjrwC36RJWNh
HWUq7vbXRczmnUxMoj+tSwyeyj+i3q/btOL8LZ33JhCRb6MmadxASYcB4Bo4PoDj7YOS7HauRjlM
SiydVPYr5WsNXJbiOeTZve9K6LEesJDlxDfvMwh6LrRnI7IuPEg58E/oCXQzX3F63QTzHPaSs1Jj
L2N4axvF3D2TJHBEGgy9QzoqXyO+054/yZzsSDAD0PJ60Ybvtx3cNtbbwTYOtkuLYlPXd2rQwUQi
e1tEwBH0xnZBC5MTek7M1Nzol/YkOpBRosAaj0eRuzCq2ZhBlN3/VPeZfGN3SmCxAGlRDs06hQ4U
ofwoyQX2Brtz6nQLcQR5H5TPcjIhPa2KTmK0H3tI+VAiG0wSEKVM1iBCqqJ0JocWMlVsnNKNlcLi
Ao6/bEUvB+BX5zm0wQipTG3Sy3NZ+5vpMy25vZ5GU4494ObPm81yamKH74Kl4psakCBGGXP1AU5N
4xC9u/yjspOewW+YbmNFox6S53xJM9vm1fFw9lyyPi1Jcw6lmPn6gF9rvoJVkIDWIGYGzn182l4K
C0e2Tw/8Lph2n/4UnpzQvjpgP9bQhGjI0VGBvuVYp+BvwNySL85YFAR34zt3fcjMt/3gyaTIh/6C
X1O1TTaZhKubujb39yp+tYPl8p7iZkT8nVAW4pXIToxGeG79VbINV4WFgavaL6V5rHRsCh5bmqSM
swbrHr/U6CIzlMKFqtp5nxsgsG0O8ZWjug87s7EaqC09UdereLrZF7E4BPHUONU4VYA1MMvihjlP
57UAzp1pfFIODK88wTri2IJKLo7t9mBYiqtV+xR66ZjH0Pa/UFWsNieQr3Mox20W9g6kxAUST9vg
oAopC2rEvUGLHSIx72ywg8fLMEj7kfR5om5xFm439w7ypUPxOoJMdIbSBEppQCr5Hs6sh657qH1e
KM/twapbrEH/36kKYuNw6eMMLwNufLu4T889lTm6cmpJGVSZ5uKItJc32ZUrWtJovR3qG1uCyQVJ
le0Q+xmnUTfN3TuiLZsxD36MbCn/ew3MVI8lj/Dr+PzWY3P6K6Uz6lJ+A4F+eFfXzQzP8zylrrRw
tC7jvjqmM53WEUGgSyqvrGjBUwQgmgPZAHyMTBsMjbKVDsiiVZXT/tARu8JD/gT2+iLGGmPyLVTZ
tIy00mikLVDDkbCetG7nSvlia7wttV3rLlGyxuQN0795E7UmcjiNgN/t/A/UZOYqjf//AJinhDG8
vvRTpAmgNpkV2gn8yOJ+nfqOIh8exXhSVW3OwGgYUbu3lAVlKYTD1D0KmwoNboczB1/jLqMveTLU
pXv6Hnu2wV3T/1kX/yakkYts9FOlUxDG9Rx4jrEp3NuZWj5LhwYzEGa5eLGYhyY4/8uLQm35tPoh
LdPXC+lxMukto7kop8Dw3Sktgf58YgpFcq9FPn9LkyExSAnrUOXYYQhdWtoP8GeySpL6NtjDimfc
vyrKChbF9RGneALEi9aWwLUbft4SVFC4ERP7vg2EcCT0/LqPWCswFr8Nk4rd8xvjGVOtrslxG/oN
DM4ssSBnqjYUviSk5x2POv0wlyLXdLlbCQpKrBoqO2CWy4NcG+KH9KHWIfMP1T9HeMqeYL62cJ//
j+droEi0kF44ldnsxcgPaDf56GHyZHGNQwHos7TT6qS7IYENiTkdFpgYvceyk/Nuse7sA1UfMFP0
+kiZSbpne9fiJeFuPPeDpbsxZyU8FiCJQjq0O01RLsZohLU22pfguP4dU0nvYFQaQunUhj85cEYX
eEf6Tz4PpZo13v1yQTcUThYnOObUwBUgYVlkxmWLgdUFtDBMb3o3BD9gK7GFuDB3wKr0I6j8/5yG
UBOQCivkgBXu0wGc2Q8QWPFRTKUiWaUWJpKyZJwbVUg1Mw/5TPozH8CTi+JYzUkxogIlCS4GoNau
lSuk9SrwNkskkY9o9GhmE2ab68n+1/TMg8CaIvsfpy6n76M1vc+F3eq0N2bN9OK9Eb6jHuAyyNoj
yBX2xJBVEEDL3sWNAc5+vxCVuT6Fe9zGaFB+D8p45uXa7vB2l68PDy4O9m3w4d9c+LFr0vBH6Yxf
39mv2nuTtdD+wVF/2PYDr2CaRMSgB9PHSxWydFhKYuzEvYGUQfeDhXbiJVd0AcYW/vwrfTthY9Da
6mc+HPNYx+xHx67JaUND/VUJyrlvnvBqqE2TRDE89YoRmgdMVeiQl+salLAe7DluosuxBZ/XPyBz
nxj8HM3Ic20RvjYcSfekwEm8Ct3dLMbGVLlzhHSZbYpJWzRsnwcqzUJ8/kbrQcyrFziv7Eh1AJPT
XGO9KJ+Hp034nQO26hfD/48Gr9paWOpYmKVlCqGMyL9PcYKhKASNUs8+aFw/wRzQY29ZwDEvksby
w+AipIJjjfqpsnVcxo7h9/QGq11/AjA1M3akTfngY/5Bd2iJ5QjGGnzJ4wSHapUEZ5x9oBESCBdh
iSyiRyk+3SakVPOjk6Zw7sRbEJU2ibd1oyCFcZm589lNZJQTZI+/ZnZACrvoXXFVznPngD5o8mTO
RExmi9J4LvDGChauXeuWND8+0U+SVuRlxTtKPTy+aalt91MUp3yalzHgjg2/yC50X5oftObSKSCa
Oyo8VB8cUq6NwRvvXamg0JgiW6AObQ4GVNq022wnGjUq1PeKXuYJHYnsq/oFStqrEAArAyWz7YOZ
lRLSTNIYHCN7Pctg7FDP9CDBzjVlaCmzOgN/I5VU0dQD4gHs5JF7YijqciLE2PHwS0Hcf3YVKnj6
/gQxjoC2wwVUdv1lUSN2Z0juGhZIDZ5LE0x9JZClhG8EjZ6VkQdAR0LEJGLuUz1zhXzqWYUwbdHY
nURUVxCFXmcWcP7ieJ8FKVCmTvFWC/n27Q6z45CTUgPcAO2cdfIOXdWbn7HmHFTyfsHUdNWaLJ+8
a89MynfnYOwE8oU7Ny8zcylF7TQfjLOwZaSGYml6pzOgv+h1o8j9M2DYIh0QqeNhHAfOSYwvFcwe
k4SXy+7OZmOoQg/9vLgoRxjJt8z63hJ8ZDyOFXXIggulxdu/YG3ZArqnzEWQQCWclIMRMULk8mVy
eSQQ+rLAXeflTJ5gVobH32x1F8AMEzvSCR6citB70NQ8dNOeZ+6x5DXjMVCZdOsdmbocgsZenMnA
SOqHcgPvVTZdh9u73Pgjs/ZFYHZKgwNpxvCPMrjmIj8MRvGj+QzYPZNRGdcrc5oOnyDYqCWh0ouJ
2Tqb6/QjB1KgLAEHxqbBD3pD/K4ojaPLSUaoAgTr8mriGg6DvhTH7g/TWC+eF81MwM9EPNWzMxEI
lTHWsh2EG75WernK+JN3kzAR6gmMR9LE1aioQHD7t7nyGci4G+KHix6WLvzOKv+pRSeB3av8jH1U
tC43qvVu5O//YLvONNVWa3LE1c2sR1YGfDiYUsykBQSxZ0F5nH1cqiBANFGMfIh0CWIvzd1aRSDR
8j32C+rZY3cdl/6yqXrdra774a8gr2ENlWCIUABRuHvuX0r191DIExD5ulHNhZreezgBEin8N/q/
5mNUcKZUDuBNOWKqUJPmLGWaxZPr+ac1T3FpY4eGKWQWMxCb+IF8HacgC+FyCmw85Brq7hkns8jy
jBSZlKBqJUhNT18+KroNq2re4epoE5gO8g6mIi4Qe6W1+effNUtklxUEPkQWkiiQUhNQ2sBJmWcU
VMtyqlqROr74eWIOrnbUR8ycnCnb/2tGqj9vIdV+TwDmlcb+jUKGKi5nV0hJEGWM6V3aeJBT2nJr
NrBPYfbqHDdhqYtrou12kor+myPq2kE5vF/uBBiafSJ4CLwGa/HDqpyqHzwdcj3uko3lC+R6M7Tk
1PD6ciOTD6GtgbvrAPhPkqK7vSg0SbOyLdSzhKmrdDfLf1Lntgk/DaLA6qjtP+6aDU5IdY2qdAN4
Zdk1kT34ZZ6R5W91oBYbDmdPDcUkmrcUyfxRRyUIbjmt8vH+fgsf+coOu4rVLxmW+G+I5Vwkm8Em
c9+XHqdIPOb/V1hZpOym/lAg1arCorC4qLpQN8qHXE1NQdi+f8R5HeHoUm07KLPsGzoCDXPIKPJ/
3R9C8YQNIaGKZQUj3/Iq4gY2Guc+mqWFVf63YFHkgU5MMsHzxvYNq6jXxEk4y9OuCrlJe5oPG4ew
aUdGokc9LBZM7ByZZx8m6TqJNCBujBkhU+9STpIwwncYTpm79RNKy5nVavzM29gpUW+5l8ctB2G5
SjqKTOmkC4eR3yk08V9uhf+N9JaH755naaNESrR81NIJi4ypJldSii5eRkeKhEz7rxJ0aNVbISeH
HBkYIQqOwDPKebSx65GHNpvf26PfIjy7V2yuCNZeNilg+3nCCKEjJWIudK87JVGQEVhQ5j4bDzNI
+/mMukXvwd5q2tFannPMMG5El2zA/KfZH/uTIGK2fi12TGNs3Lt9IZQ344Zi8tv4nUumbMqrTOcY
TeUJId+lHLQQIH71qQwhplBCSjAzpiqjfJX0/bqPrX+p4BVoJf2tcpQiC046cDp3TK8Y0tqu23QW
OdzKKyHSLQ2JJkuB/7usykIyu2PNKDjlS/1moHd5SiTOou8etemhhPHPaEmFSrdYaJo+lr1HQ2Kd
bo3FdB7/QKXMRJIcj6DRnvkQMBjYvaD88Nj1efUbo9zX7dYTwuLhe+b5LFA4vUA7wA0IKmAAzYXs
mNfvIzd/sA+49qq169IK8Ms89ACf4bl1D3dbZAvhn6L/cBWMCrjUFMzoBJV6m+6W4iOpd3aQQgfk
cj+rumrzW2uxlmMUGdNHlH4UPpblX33/ZGFy/b0CG2aLrbJJMqFxt8ofsxQu8/4wAElclHmCEY0j
9NIMu+6m0OEKwuBaP/znRiFB+Lfm8gBSoT2GavLEM0Ki2o6qfuR+KM/t80CxzD/PpTnKDIKL54/k
t2l1Jd+tMQeTZfiU4xcUeDSvw/92GPTVUpwCtlYFMPlaXYyrdg7Qm1ahpzVSF5Ir8oTceWdp5qDW
3m81WOISU9IyzVA6SYDWkGmXBoVzxW5WHoxrWQKWY4cckeeaygKFOPtCtgMei4bbwzBl1H/mSFpL
HfxU+fC2DjFfU6mwrt3v6JCVJK91ua3Sy8bfvkk9CKvDswE1DB7EQe5yaxIAHdqrzlFuwdo5xEAi
/RGx3Dv0kPeP2ZdBdJjptr6Z38Twof+Vzuogr01jceF1V0Emvx+nho+zkei5oSRaGUi98HOlwguS
pTi+8VowLCxPlngRWe+I9xMLHtf2ECE/Lw5qVIMvq46PBodubFyuRH+LgYV/fJSfhoUv6fr+IAQd
ble0eScShFkLg2KyQ2logYVFctGaM80FPB8wJ7vzqIU06xQdO43p2mOhxiSlDa5TS3Tc+6VVahjk
XA6VgZ4kR+v5abn1P3XBbQFZ0myhW0nfFp8yUpojFmeWHWrvuSbVe2L59o/mFk8wBUDTXr3bgeRT
7N1JSk9m2u3F/GZUXndkhMlXcbHtJilwKoga4h1T+QoMG6sYZVrLJg6KkSQ8ngzNQ6csJzOSLxiT
OwQjlBty3AWsy00MIXICf0boNBKo1DCNVYvscPXyiVvgBQqugvgnv4bcNM9E0gfQKxVI87xkP61e
NcEpTljcdE/1zhlgXxm2iMf7Ikc1SBKH4mRsIaV3h1+99JBWkGskrXvuFwZ99T7nWs9ZD8F9cMjn
9nNZazPFfcloJW4tmDNIFcMgGy8En6BNrFvnpZm5S+JkyQRES1myd7cF6UstcIy+WUMEoCAgzG1P
ODEYpPZqwkQKtAhWWYIXxDqcXRk4V2SAr9w4WKpmcDziVYrNcPUu/j+PAe2hOFpWqBRaGTTqB5JQ
EnD58AyRCg44wwpb06fqWRr7WxZ1yZKuzSFj6tb2OYUHucWXIWdK0gd9pDR2kVNjjtc0hf97hiD1
ms5HBTAyP2lBQ3A7hY7zg5BVrOWmAETXWIqLPKGfc0c4fAwW/4C1WgoxrSaRyabXB1O56KA2jB/W
Dpc5shCgvnERgtKb0sQQ/CL8aK5gFZCfinkjhmyUe2bFHYHAt9GRD+Yau789SE3gvgoLvJ0/Zjrs
1clJv/A1nQjJrayxxZLyHndJXpTmYImfjZMtfActkIOauMrV24n3VAuzY5U7O7DNHYHBx7I4YMna
aDq/2T/R+/nzGFa4VK/wyPEv1DtnZOLh/RX3MUqnqb2aQq6iWORvGaPFKh9C3WaY5fm1ZK0Gydu3
5u4A6GSAtWgxIcstNyXRCUKwvdP2tkO/3yWTlS35SqEP0ZXL/whzPbUWYEUK65/BYGTh+gTZOanY
09d5qwduN4l5NZ/NEdSN+XXtFW043IGNN1TXsHOoRo/QnwEHvKhaxmKkkURTggjtEBI/lv9mfPg7
rNiLcA2Btf2yHjhRBAbUOYhKIdjUlgVK+SxnGOqXfA5i2QVUNVucP6jHITt40jTxHEAFf3KwPmD9
75WfinWNV704D+gJ6He8wwvkrDWb+MJGMV7m103/5DYz9iDQR20oDHdBOcfTpOVzSd4sFgsLTp/S
XmRO1ZrUEwOlnpwW2LFSBhrjPapfZtGTbOEtkWwt+32VIdBKH4qRcRvl+Xj9a/SleYgcDIATAxTy
HTMoT5TTUp+k4zmyUVtu7Is9MRecZ8fh93/qmQFhZSdoFXSOJqB4jwpozz9nv80MkIJtQzsLvAFU
2N93LYnW/TmJBMi1pSGE0uTzwLtc4iC2JKAxQEuD0eiWQ8CyEd2Mb8hrl46DYq4teHGWoWSe3Blq
Ljls/o9xATq7TLMcUP2yRvXAvW7PXyzE0ouRJUssM+NH0RWpJ7VXAbFF2J2d7XBYDHJ5RYK81ATx
EkogcGhBxiDoq+CNUDd5IyClCayo0pQXhMZO7Xcnst5jEbNXeCVKWHQ/jjKGz1J4xD1pCE662aSg
VFjZXiK19AaoR8DDE+MVKh5ID17Hs1ffYIUYu8A92oD+QW3fUqMLTJKAw84qqcliy4vvpGonXgDy
ERwQOK5IbKMRuYdAlYW8Luovo+MKMW73hYwMPWh3ZY/W5tgSx7RiQxV65OO+5o5l8ztDbfEFycW6
nV0N3vztgLxvmkvHsESFSfF1bdf8zLHwJrvkoNkFRassmo7dC8AFwMP4s1Z4CBuwL6sT58OdY7s+
sfKOrl/GT60AU4pyepODDPKt0v/MvWGQnCvunM+fD0qJtHzTRMIsjHZ+GZjbJpeO4nV6Z9gBVVnR
oCMox/HFe9YnropKgb8hIav2jkZ/R0xuZYtLKLCza74srqdWvKS2BdnNslYhwf9UGvsBwHP2O7N+
m+z9NwJ54Yh9MW0UcZgUwWXynfJWv1O60nwdyZp/tz+juLbsBPQNK3ek0Gxp87DAW84WhnARr8LA
fH2pQHmeQUFB4whk8BE5Lqx0Py+MSBqMX1oHivo2O2Hfqt/IFQGilu9pIvt07tZOwU8MBAtX/gO9
lJlPOuj3gqnFcLwfrJWc/wVdFiulOPcTHZpuIsfRO+NFDbNlVxz7jpvIo1poXhwzmkTEwqC+Oylg
LXFHJYLgbGqQICzdZHq/LgVqVg06XfWq2aJopETU1WQ6tjSgjOFdnm9kWlPrqQJkYuYVlodVa21v
wRrKgyIM2R5xTtH7BQ1T4FU6z7YhRQ+/quk7Feq7T5QOVP9zetzncw6pvgpO4pmbM8NZJX+zkE5l
gRP+sG7lD9Xxcq4LwBGWywIxttzQNefo2B1C27AEU630pue+swSe91rlW4vHgaGoxfQVDCy2UUM5
FLs5QTr7xOWLwcilLE9p0MiupttIqnMacAUjlZc9+uMBudSLhj8t2l5O4kRVojv6sHKz84qJHyjG
ezpxdK0jVx+lActlOyqhnFWCXxuJR768LSXOueKtIQzw+jZk5tyAMFmPsSc+xpDg5c8wHf3iMlNG
fDCKmul87XV0Cn+n9BgXUPQUL4+pa3EqCIqXGjvyf+UtlopelkBUPRGVeiqnIcWMId69KroZ8Mrr
U3wt1b0n46l9jMDDMer6ErBPstt53TbLNDbyfzG/XX9gnGKZqSPq6AoxPVLO4WJpicSzl+p9ZBct
DdBiqXR56u+llvrdIu9MTxmfWOp7gISINRFw/AGqc/kCT2VGnJ4Wv0T1G4d+msU1Fx03D/53vdNZ
ezpGf5kBUVoWfKUZ3LZ/Pajrq9PruzOz5gMeZhhoQMbyd3LSOZB72f1TK5Y2n8LpJkAuziacWjEz
KjlOTdfR5HA4Q2MZ4ir0ZEWlMhq6zdCxLsrncmKVRX9itpofq71LX3g1hRoo7DoHsDv+P6BNaT/A
NWrlzqyJh8WAkl6MO56ZBXj6k8uwsvZerlizOsbJ3P6syTiYXA6FCaLrfKxCwHu6fAL+U6qMO+8N
oXH1v2ShI8rDXhmJpjmyL8f1KXllZVSwytB463vRBfubaFJkdLesnLfIBNfgfCX6PbiPJuAB9vXv
EMqWDTs/vUyWeUvjMPvaSMtC//4oXxqpX/53ZM6TviqiUtuHBHs2EOL8QnXvynCQ9ea/tO3uWMUi
1fS4gtLEkcyOggLZvUqB/iS5IV6Pq0Xr3UT755vnQFCcUcbAVcJs5vjlRJwuj+8RKvswJOPbDVLo
mM5XKPdkrPuEq5c0t1l6q0WqFiA5bRnYkF5vyva9VYYuEOky19o6k7ifIku03xeOy8aZpDc8oXyD
eYAK6hmc2pU+6FybI4puf2/nkEPJinM96jrQlHZfFvmdb5f1ZW6k5Z6YNW3L5CcV8pQa1TOBDEYn
m++EDosTXmjY1OAbzIXfuxHnLiJrBblxQyMV5dnbdF3cXpji3oDdMG2KCEoiUed/blwy8WSde8Fl
yJrWt9REkW8s6M7QmKUuwF44X2yi/fFaMnm1rHLwN+zim2t9Y3a0yHIviKT92cez6E4BMsYg5+5j
WNQRfegD+Kv3CkkWzepWfZ1kcq9SC01IbZ4seV0Aa6j4L2ZYgodMa+l9FNmNP+Kvg5IMwRLnzcST
VtkYTm4+Kq21JoyvYioAt0B/Tq2RARAgz2zQNF34wn+MP2Vn4SRJFPwoQeaOUEt6SNVuAO98Qrct
AJItikqdZymU70O9SKZAl0H9kcQIk699DErY0pzWaXUSXSjPbJwKahq9p6wVvuWCQ9DvZQirah1S
8QGck18FUtHJufSr4OyTfygFvTCoXpd9oVuoMMvk54goXu/NYNVv2rDTKwq6u7K+v4qfsUM6ZJ6k
/vPTLBI2mdMuq1DzwYPcD4uQ2RqaCthz9dHn58JmNw/qb5EW0yZMA71gpCWgvROuqju+aSh3MY9G
pTSa0NaVazOCdT+GoKYt6bPL7LlMDnI/EnKqSaeNAkZ3MNuWg0DZRYZp9DC1Cq0Uf532Mqy+/v/M
XArfqkSIYbAr/dn4H9h2TQBNv/3gdaSJHIrUqjUgxg9gC9FDlHlyPXH0EW/TZ2MxhlPLcGMylGWV
epgphdzs8Sy4VmCHGugkn50zaTxJP3ceOXlt38kG7tbjpUEZ4x89IJ6OdHEjOHzrH0Gs8LMgdGJU
Nas8azMd2ZOCYqjPX0aFqCRtEaAD4H4WfpQiVdjuT89czmQdEYzwBicuPFQzz1FzcdGaC+lOhwiS
pFCUaojWt4yfuYRqh10w/PDqiMLE/NLRP0aCZ5rVqZbuuhJA2ZfbhfB6Np2aSbrpjTFv03aOzpj7
O/PYecX787ZF0irpBrjcc8gZuXUhao3eKH8/ayzgfArSikONhtg+0bhlTcC5/tarG5ib+E/JGrGb
zsu1hiQWMgorAqszGyeTfppUz51YbhAZ4j37sK36BfWLxguliPH4j38b3XESlL9D0YsFl44CNuch
FutvwbSlj6YDAmAVQJ2roQFu7IoXPVO+kwiwecyI9csiFfoKSGspk5UHeHisr9a54o4D3r3qXwMG
kg5x7Z6HWPe00byqgZudtfSfzByFYjkI61QQMuulDSGFKOA8DdqjnzCJ36yERQF+7L4LV1pnQlLO
sNmaGtnjN4/WtWUCnJVpBxAKqbjiEyroTGGekdD2y7G9EE6eZr34x0LfqAYBzeTIJx6CnGh4y5UO
93HgesNlrvhr962tf4V6AipqHDFcftBYD4qtCYBRWEl3Qh14b+BubWar1stnUIJVG0RBX8H5p9qL
BDhUlfbLwACGgQuB4F5HGVpsUlSvYsIMpCQF2CzENbsL2g0vFh/TZS24u+xukGMYU6yOHdN6vu8W
sS9mjKn1Vs1mo8HWZU4PQgD/E8sGWr99I6p+VthQVNOuMgm8DewND6mQs72lBaBbYHR7rWvX0tnz
tc90/0MLpVlfFk+G6213eRt1zz1GHj8GHpA346a1IJLVD249fJO7gsn/2t4LlMbzBZ9m3uOzHzlq
79GEBHXbaSoxofytyueZliOLDYQbdvkB2sGuXrDXtCxb9l3bql26ECakGnqQQNIAx67ZF890MBKf
TbI1ZG+mtQwg8j9VQt0nqUWUgbjIs4RnOMqlQfaz6aNAuObu5DCAmD0z2YFUsCDegE5MdsDcc49o
khO9y1apUCCgqW6IEmBynmFKpWM34SnTAf+Np58cZPHGnSLp8t/Fpsyuu6rV6dF8ONGp+lOVBTtm
zAerAPEDQqsyuup1FP8UTOQMvm0NynhAUz//rsXZ12uT96KZGhCZGDom8V8X7Ph+A2LkAD+Kd4TE
pj8fk1t8oop4v1FEeENsl9S/EbdqKB3aibK49mFeMiv5YZfreT+SI3KNkqBOT+WxxUpUUOARxKcm
vWOaYDO4usfjLXIF3QU/bi8SLbrFjMVQFWhTB4JVEjWJcevhXIdf0d68U/OPyXtVWLld67rRJ6GB
gGSBv4fkPjzBHhLJAKVF7RNj9EmjEVHdU94OfkXGGzItHkhCMLqRno8apjDaBNh2QkY66nA0hwOe
4ubUqbSuoDLighebi93DTkmhFB5eKXtzc8d9q/kNDE2pt6fosKOxWSfTAFfvSoGcTDwiO6Zh2ERJ
WFMWjo8PrGg52GpIp4VCwni5WXYAefNrSA9vLVo4hxhOhdHDoiAuV3RWZA4VG+B2meoZdiL8XEvT
Zxx/67sTcyL8yfaGK7KwV8p4VbTSf1WefifZl5YwH5fdfaml+X3eVL7EsM4SvxBTHGrsM5w8fo/z
fTxO/G/3EqY1GatQnRWXrL4ieAUtPW8hKontWh6kPEOFHK1UWpL4mSPwg+0hFX2Hy1ed0e9Iqu1I
H3WYJQMJKoi5qRvSA1EWFRk3IBxS9goHlEz5fNOnTam32JzyAXPB8DbRdh2045t5rSO+fi0i0+v3
0qbIgIX8HRmA2wyE7jaou73f7slaRpcqqezWXcu5XCmrV7HeXEgYjGsJPdEIC1nOLko131F7O39Q
omzPmlePKk6HKWfecZXk9QzT/xbX53gFwLnTPrOhBgmGABBF/uBXN24d4/tvLXzytmecjetZwR8J
gwnLQOdDwpxVtmBoiq0wyG4Vgzj9NlrsY0GpTCw8b1raXBhi6HkOWdEWyn1x31XOaXt3e1OdhhH6
nGkPlgd5Y+WZFCMaprjz0Dz/6ZMqsRr9rENS6ERuzG5l8Z+hN2qFmg+9O7dhJX3QzUTTkqpud0ND
0DyPHVoJ1qJwxH9ap0yNw3Vz5zwAgU3cshw/jW7PWn26R5wv8To2+9Ve5n1+zK8D8XUbF8oGN3PZ
FS8DmHLvX5wUhOTLg82z0iP/Q/WQ+uS0b5t6glN5pJSaHsj9n6pg9uCJJd8wM2VVWyBD0m5nkKN0
P9S9h5gGg1RzXTFX23jSxLHGfyp3veBE4XxPuEZ0LqoYo5sg9nvNsho/kewDonlp3OLJLjHpLRJN
rE16NQOy9W3Zv0vAfd4pJ2pFoBA68b7aURR/3yl6y+IJXLu6cg6oQpZu+CCuOH22ktyYR9814IDg
S3d2pnyoj9Btp9AIwl/5MzMtKD/jaFg1tPAUKP6f5reAYrN9x9eYWswcPd9jhHdSYrHQR/U0nZVq
Vz7M7HjpnbasBYD4vPnST6L20pv8Lm4MEsbcv1LGbPiGu7zV0WdsPq2Fyf6umEscTjl6gU12Ip3b
WMrLShTE2FXWZDeqCpZXBwA857zKkLJfPwncV2eXx1SRg7fySFvH7zNT7CotTarsp1b9sQv16YUh
FM78dbHbWQ9whnVuH/NyXnOJdIt76Omtnt/CBFsHjKcYNo2vB8gfU0bO94DqLwVb6rLIwE2Gyuns
SIitYrcY5FVfn3A/qES0XxuKVYanTyZLj0AcD7oknPhTariLlRC2zWE6o6HBvLNNjMMTKSpUBl86
I2AXdbwFA98u1TSd+xQ1XLo77H7pwdLSckkU8lDPFG7dF/Z/dkjyPxQVvBQSZi8K28uOQdDq1VIt
XuPp9yOOxBcNLDcrhWOSNUeQYOfIFTPsUF9Wma2SD+PQ4YjUFhaONm3R1p+bprhD4jBUPhFB6aq1
gGmSzyhMLxQCOizfWvDglaBOWXeC+ugVzjdn5BYu+65DCKktT3FwN2e34/z5bHH1uKhxgiIpr/5y
ViwpfuRafbNBkfQcesher5QrtDqnbafEXChymJpmQngVKrkUqVCEnCwK40cYCvTfe9o+WTpZLUrF
oh+v/yUJ2OLTWFruioQfkeNmrycfQ6nqXN//+Y5Dj4P/0CUJXkJhwnRAB7qXkH5+400kGSvWzARx
hBDXjhwNdiIBqOfAxTh7W0RFHQSLTmLYBprF/Jym68WqK2eVUSZlz8AkWVqlrGPGZiQYrSumfBdv
+wlZnnbyswB2AbATmsBH1GST7xeqrO6pXghQJAhYJNREZFzEi8TeRGnwYFmyH6mFVngK+17OV9kv
iUNrd6ItunXe9v05j4HOT6UcbadG0q05Vc4VXCxxSo9jTSaDaoC7IZhqxfb4Rf4uByQPKy6czkcI
JX8nHtSh1dPXjSBtsqHXCE4W889w4bkYZccwMQUAGrjW+r42pA/3BJPmrP/NXwtlo1n/SlQSpVw2
qFOZvmYBbFidpYr04qAVpu9xaFcZ1ZxiFsv4Hq57ExK5nbVII47B/3+hhWKobPlKCkgP7nLKKmyw
6x6Aw+oITSsT9Y3CKJNcFZ1izWgcl7ZIv3Q1EBavnw2Ng1Fxznt0OdR9iOoj4q/Ez7yxh7zsr7CV
wWehU0YRtpsV4OaG0H0MEjTFL/zGVpob1hKQ7QP1KirHz+zwV6hbKJN9IOrQf/uAVrjIxKTcqoDn
4IqZnoS4c+PASc2yehH03kMahYT3TtBlZuyV53JW3krFRO+8DIfTNggTJfUgYKWb1IFJu/US7IEy
wCj/oV7I5v4vkBnxgo4tCp8Qy7I86JJt8NGy4OgLOe820cOQeWj981ArcHzATGgNIzqOKuDXzmcx
6PlUoBNH5qzJqnhcl4kCPxHYp06w/LLBYdpRQERhBQxmES5CJpz7pZjyOPB7DhvfA1Rkah26GaVn
N7Hdkz//XNxT5WCL1hlhXzUOKe7jbN9hPJvulaP/AchAqcmJzWOMekS1WcyET2njzdUnQMosX1YX
nw6kigA7Wa+30HlOfcmKVpceuYSv8TB2F69K++6lA53HPWL+xGA+aKJdhMRCNki2UgaA1Nh5Oj0H
uh8g48XQThGrATLl062+V4a/5JTEcDxaFn8KEQfGfuw/1WUrB3hn3K9ndlLRhFUtK2f/E1GgtADl
6qzdS8SR33HvMa368Ahb1PUH9FA4pyaDVnXXp6rbz8O5CNVPPOAdkWZUduR7ltwUKdsPc/9il7HD
m4RUciL5iZxutAWoFCpRsMpo9Ww3h6LDQa3qlrzfbWAYiLXXTWRxbF6gmVoBM29VirzvfgYb60PC
8Hstjf15bzgubAF0KjIbAozdBuC4R9AN/uRR2t3YIMmINaCFB51ivZiBq8JKeo/nIyCgFB8i4YR4
slVuHMr4pESNTef5PM8lDpBZstDbm5ub/tYvRg3vuzUhPLO0aLmTwzRsyWe0PMBJ1v7A3HNO9YF6
Hgu2rzm7PvCEwBi6d6kJ/RH34mYQqaumVJR7e42eYIeDA044OwNKTIBsjgvyfsw6JH8JWkL6SJzu
UpJe5nByeyoj6QHcrcwmd2LiL5tK4IgC5eEQtNTpWVjckRkhWYxhQDyJZsHvJhCPUjLFfyco+Qfm
FI8bCGyAgo8IOGZppKWeqFNp0GY/oyDzEBTVZ73MlFZIKHGoghYQatEdOcZjDsIz62Mv3Jdc6O9E
essV5DMB0F+PaiweC9vuqc80+jT4gxV7C5UOiuIpIHY+hX552HmSLaD70e2PPRyWCvDSh73htnEU
iV5hcCHeOVOijysdmzngcLH2LZb/58jGG1t5ADO4mcxWgU54I6UfE2FIpbiQGhqCFR/RzYmoOdaf
JKfN/gZWTIUG/E/LqVdF0yraVl4FxBfnUOeEORwOCGhwpGwutPwaDYNF9hOxh/vSD5vyNUofFv+T
LPqs59o0T9+4xqlo/e45hiigdRo2EgJMQ0ftUqr0ZyFCfhsqJb8lHn/+YLZ2h5+LQ17VsWVj46MI
8KI6DQjzK4QEafd/+9pE/UVYeYQTI+z4JtguBTdAiX++r/BmDGlOPJPGMpunfOmgF1mwHQCJGC9S
r+oJCpG6fVW7hJvECOYa0H6CmLp29b39bMwJG5dNbGomRrT2Ha1mu72uE6xVYHXcHWCvw+HCleRn
bxdmdqS0ncklHm2yHQczFXnPfeQp4KU3i5YQgLHAkwxXf2m34r/jximTFy1Jf8s/l9gBFGVYNg4I
SjN2rRYgqh5l2yR7yDQI8sNYuEp+YTp+l+POt6cdkRdsJ8/CeZWPoKYml1e1h93VhpAHlpBgbvCx
UZlnlImJoP12eOYGjeUXg320XBeEO2jkNawk7+FXWLn+Ipk1mLYHKqNVTAG6nRsJWOR4kBqkjSPG
e1BOCiPSkpW+IVIYKBlbo4WbSULHSeC4UXX/ADyjJ3T6LExTk0beTgRHNJuSdzbOGritpllDhiLi
oWesiZ33PE7C7E5fKieT/X53xWH8RWjjI73KWmGbNbmQ+0urECcwgfan1ylHIbG8ZzSsh+oxvDsg
fl7UCMHUlLCFWltzbxfrweUlLHlQrn6PDsDv8omNGDzEa4ktJaZ5GTOy0UIziO2IcklAYiEJSj+f
VLV3JWvSlQI42/O5b//JoYhoN7E5CfrFTH0rvJFRwAqZKEMHmSOMQRpd/GvWwVypP92/lN6UiqkG
Eb8bfbhpy5Hq8tJlsA4R+qj3K/YhT4g7BSJkRM05+Qzg16YsNj53pM0ibliAXV9jR8IqJr5udWge
jqtWJMfF999lo35cRJ190AXjqqG/PeN7a7IsMzEeeY2hTD0IjgK2toZs4IH8sWzc3PYvNbpf7nyy
fQ1W+Yg76y8k1zB9kwdeLcvCrX+qzoNtYKtEWW9nFUqiiFZqLKMBxcI66I5R9vf8NUmX2wYLBnLS
8q3xQT278jwSjrU0y7429rxkVLtO7AG5OeZ05dyer2MPWUQVEQhW9Sjx1VOs5nfdLqIAbBK+FYCM
QbnPgMLLldagay0MeelD1Yyt7/+f9T4W/ZLs2hamYNjB6eafSLaeG5p+rQ8oTjSbifjVTGcVnHZ6
/IXN0s5gAIOnY3W3YIZSezIN6Fl1FryP5hOQhQ0wLOxkjjEy8BQ4vn5Y0wCVKvSQzplHy/8utMs9
JckVM6iaJ2mq2fG/eveTD10ykbL+15nN4m/DyMS65V6/BUb2fPtv8HpetJ/fdoVxub+yuVfazG/p
7sRDQvs7R6nuw9Pt6ZayRktBoMa7IZ1yyjN2PnsFhjRs2xch09Hl0+HLC/9cno6kmmUICuKFVfLE
uvpwNX74x2b/MB0OosyAFFF90Ta5++1nhtUhsZgUxdP0yuwIJ2RPG1b/zD1NR0rsNChkeT7tA7Rd
3YRg+QlaFuKEi5sI6EnzADw++oBwqb7j9M2CUPboCPgcmbvCW0ZmJqpESVbo6c30Z6Ieis1/9TkL
XQnZxLKcIGifFrcwAk5KcoJ+ic9uoiPNuvZNqOmqu6ZA0JaH6iFhzUR/GkY/sZmEyi7YhQgpih6G
qdQn3O3hyrXSeAvao8DoTwgbB85/2T3NDkVC+TBUpodRqe75ZklJJasZbE+VqFcJuSkifus8Ua9Q
pUgXTu+Dpn7i6HchdVKjOWtlFcUQYpfIaYiUPgIOW3ZqcOAVM5PxbSXwNCr7kIkNtvuWvA5qdXT4
rcqd61eZrfnyldNr6zMaXvjwl7P/RYR8LMMkoufrBbykI9E8fa9NG8r1gP+yoNlLf74IZdukiPzR
B5SryZI1nec80p69qrfL4gNwp3Zj9OyFTi0UzwyelwSjLjRq9RwF9PPb5AXtJtk+a4qbY6UZFN6N
8Trh1pHUcUyp0RkxEA9d6qiJsbDOb5zXwKnHp0cq5KSGExUCkFnvWQ/YSIj73z4YWYD4wWOprF2q
yyqY36RVX3v+G/Wxzb0jeRxd6FZuGWCeKHzaq9WzXY+z9RuA9CBYQbhgf7w4YzelRbnwte3c0DKs
FtyP6rbW9o0F0Famzj0Qh6DekH2efR0H9zUzFefPrHm/9e90urFKwITGiqgiA+2e2d3aC+oDt8yf
ElC3qCzDuHe7eWRGJI42MMeAx0wnnr/C9w6Ct4funqDbsX8gigdV9HhLguyqKPHjJkNS7dDM1h1n
2gOdLQWJZAjhO9osMns1iqPTQM2Vmkh4LbiN805LOMV2RBo/QfCwnho3w+kqLWzDlYcPYhafGne/
np0yiymAU9/iYzQzTUC5kvLdDUknuO0MTQ5FOaxwHQHi5ImYa0LR8Zm30Vp0ruircF8oy+L4+bUt
lw38JeFG4XUId+1084P0KDR8kV7LkfjfguOaNbgrW1V8/O+QoicV4JxX/d+WR1qSg2yFDzplvmFa
aEfjH1p8fJYsP4eZveVUGep6YVUBP00g5xmH60L57izvDwupm5SOo0rh6jPGo1SoqLBQ3Aera8yL
YlNRYOrtgZxMaQtmYr0UrN7XsDddIxtLRiQQb94TAMFvls9e11jKjad5VG0cm7ftzexB+F3+pKTf
tI27tToM3hwC/FF8FpqfNNn+Z/+tEhmxxF4sttXsWLMfdRvzz6YhYn7LR8jEt1KL1KYDSCS0pHSJ
/iwS4vE3P4lkb/Sz/aQrMJLfuVa8LCmL4u7oYzUgfKki6c4tzpnNI4w+xZF5Z52uXzjcEtXcbeYS
vJkQGi5TNXoDvHXoGedHpEUrRXxuxcYMRVfIB3aoOBYuiTwFJ78DXID67mefQJmgfvNWVuysqduw
h5oIzWSSpXQTSRXOLtPIU0ZjxKzzVdqEsgcqfmbv9MAab9g1MyNpUM1EltyW18IrHrcToZK83WRk
Q7KSgNms/Au9qd5vq+KSpG+TgkSH6Q0YW8VFZPVRai3+0vSv30hDMUdNU6gMc8JftV5Cs7rgR+Tt
G8x6rGlsQdjXFZuuRlkoR48cLfk/yG5TROjfKhXwPsUVYDUrrOld51y3rXaC9RJ/cD9L996HGifG
r7SzsHXepUDKr8/iMHyZy3stgYaNEEv7fIlr1XH2cY6mr6rRrY413Mu2bl6wzlzd70XQAvrVj5Sm
YIAnRi06q6MRodYuP3ni6iuqjnmPWKhpmkNqjG9verrzf41POR/qWLLkutWxKz+C9vpZDHYCAXFt
O5ED6QeE/A0QSKWnRhNd4liuNj2UepMzE4WHQXKlxf55Zc11yBIKqLaWIBrK++94Lj4cxT1hAW+/
vW14z9BD7LDMaNQWNDOb/nvtR9bKYRFM+k00bbIH3uKfUkPC1gW1+iueaHDp8P8LOBpWT4yjBZhZ
u8GC5T1gaYfvTgp5izAFVHdy6/xc0TXJOvF0HTDlC9NTlAB5tKlmu8yy2OioiNcmfcwIsGhyC/Qt
dRMH4wLZeKksN2lTg6bVAh+H5Yi3Mbg16JOjvERKQa03YS3lYHyOXfikWq9nXEHP/B5rwVDgLeqd
oosk1lG20YNdlDICiUS4PmegnXLT3awnkJY+3Y5/sWfZVccr0orPJ2fngFlsq5Wj2ohGotQFjvIS
4YUQ5ZwdNRO5K8AxkZmVB2GB2ebVlaHcWyAD61LiG8cbGCUtLYG3HICik9LljLpffunDlhmgWtrb
+qpoIZBrahzWjWtPyffuuMZ64KQI0b1LigmFV8NtVCgYX1CXe39vFPc7vMReIvg72DNu0MlASyz1
w/z/d4F9tGUX5WpAWstaba4XLMmCrYb1Ooc3ewHy6HXzDHa34yt+zY9m+oibWFVhJlmBM2+6UfQe
V9oIlglvm9sLaWZrCHNKFNzCgTU0+2fmqseloZ/5dXPl/kOkqFJRJYGMU+WCvOC3KtnYx+rkEMuH
Yz5UltanPLnuNaXfC01cmmAxRsZNXAFKVgFbLe26RTkIxNEO0yd8V9Y8V9EcqEheYbMsG12vyc/X
BS1CMqud0RZqKlhFOmCFb9Pr0dS6HZHyPBYwFBAxY+k2SnYMlMaS5kxPvOtUv7xZ0n5qpJ/7FdKr
oYSrvB5CSlF1fuysFuPykSFcTjgUPUkZbR6+uZFh6yzT0IyXuA8kpmC0NjcGBBRtBKRQzflqFsIz
LqtLQT368N4FdabFf6W3/ymPxIcFhOOQ4YRP10sxTD09T+mSCNtc1z4W01CmM71/U4kQO9LFtHQO
ibXHct2I6JHjGjU0IQCOzNfOEZfcEcWa2iwDRE3te+rooIbV2zO/hSnZHMKTFskChKUMFjfT8z71
guxsAbG9RfYP2sNI3DBow0ZoCAf853Yjq+89fhQNVvx2tyKFwyvNgFvP08NyXdjCFW6dqEACliMP
I7Qrn+DYvUg+PtOHLpqLDqHj0Jff8wMAAhYzI9C+1uibvf8L1l6qM2fJOS1BFzqiVl3jzc1Hna4y
f6IoLx2VA0hYdzvPWVY/yTgRbuD7IEQKrQGUckaT0oewxXxN56Fw2+Pw1+V/Yw/BcufyuKmSmxM0
k9M8sSjQCWI4JJEH4fgKfLiU6ndG7J+V7jGsigfQv8u032mK2mfx3HpcxzMrZpI+H5P9jC0g8xep
K1Stm7+eZLVhroHCTP0WgMLyYI3HA6UJo+X8jJfqEM6teyK5MiJgPFMjctAnU7rbWjymmafVZWW8
blgQ2jEymskmSYKD6uYGem5jR6tUryVlXHTlIaoNtTADD/99N7erT0sIC8nCKAKBlg5Pdo2UDOSB
tg0jPEZId7I1RDZWRLEOnfRn0WKIc/3tDHTiZ3jXdHkpmWk4T2EVC6HpvTdmHNhUTfA3QTxx6dzJ
L4Kig5rU3jXGzpzfd5dP/wLTpdeeQ49CURoTgtYjNaNAvrsU8iOZ1I64Y9KMdbNenElKUHSI0XFx
9Gtzx3ip43th8pbaGModh5k/pA8B9DzulqtFP8kqKnrOynXziM8gtEZP1vgsHA1DY0yRJkYcDFhC
82LWYZ8BgFA8jOvJ5lh+UjJ2lxoQm75p5iVlU39zIdPRNENzPPaFv10iW28ApNYkNJ2EBJjPWsDz
kXwqu7ScMZITG1Wvd9IjtHxkeX7GRYbNxzqaatJmrgtDwzPgKE46izEmZAK/y/CyKFWxjNxJDlFj
DjFDp9/pw85WOBQvDghaliqCv3geDqPw7hw/WszYIAHMYF7UrBh2lGmvKwjwWPpNazsNvx+/UNaq
rMtJXCVvCX2sPtY+2hHUD2hrAaDcBJFo7dSemoW5VaQuU8tr3ua/JoH2x7yxrYkpzeDWYBaTjBKQ
XUkuUiFZ4IyhYAk8mVyH96zKxor1ulKgwl90d9B19o+y8IJjOVeG51vIOX9vRXZzSODces/jky11
y7zyHNL0q5TQ29OaFLOOC7He3kSonaly4mp2nNrT0D5wVdfc4Sah6MERkhN75HTaKMbW12qSRj9n
AQ5+CilBTp5aOeVySyxr/58d2rmmXDtqQ2JY51F8ZUXsX2Xc5GUMaRxXXJ1kfaPxWjz1A7c9apmJ
kM6HCXD5CMZmafLSmZ8xa0kjNH7kan0IJIZYsYsaEPGgyRkwe6Ma4wZoPxUoVeNtjiwtb7HGxuXq
4e4SrFohbbED3/ujX4vMJDEdMBhaSfsSVmJArhV9q83/y49qtCIjHTUsc7QMsOVtnsx+Adx7PYcI
TWSR59PMiw0MT/C/vSvVkgCOGS4HY+VNA37hsglgLL0AETd+HhB6m7Q7+H2VArfwKYO0m96N49f9
soBTzcI/8+iZARqNwwio8mTLaCocyP4fGTSUOZhfVIBgg42lB9tdM9CL3DBVDZfSm9MrfhwNdynm
T+D6j/dYrU5+3RuGDCXib1zNrsk+sDPtQoAERlOF8QJ9S9Dsqn4pxuOepR7+ysOTPMtHzdU/qFQh
iBVtbcAshuqpMFyemR/NX0afD9HuDbrAIqKkdWr6ZHaFSS20a7ZKx/IEC+TXZH+XSOYHFjSI9QnV
fZKqvikNAzkxPQka3u8PFZuzUBl8MHK3Hb8kf/fxUqyS3mSYPBcsKOkKty/v0YViTDBTr1jrSyFP
hSOV2vD/5QqIWrChJ7NkVcpcQPLROfzPnxwot88+Hpf+r8Dr6u8UB9f5msAnrsL9YzxOCFZsksAF
Iiaui1z3vQGezXlHb3cYVy7ofDqcz12sixz3Ts+L6XQW56cSBpG4l78UAi1fSkikUDrVQNFS8803
lHqEjc9QdyFn55A4z0W9t0BiacwwHtB4140SU3g7bYcH/A7MK02DcHkcAAkpDD0yBIYm0csTK50J
WcidJ5ddH9mMZeOXFaj9yz7CLCXTbdZtzV4Uq+NkXtZiYiGWy4zknzIFXL9XGrU6XFR9LzEYvuqH
9kAnhQfz8W2tPgCVUvVFdGjg2FFyaEEfz9uKznb+S9zh+N/BFUHA1LYPKqSeS4SDfVlW0jx/2qAJ
FwYN7gd15I9jlcOdNMQ2RxBKPOJ17f0xQzp8UyGIc/oSoDiM1s4g9NFyxUxDeETrhVKwzOUmrlTj
JKpfQcIT4yLxRtPQMeOA2ptcphfbqmzNut5jNELar1H0Eljwzw3PznI07Ls0tKs2UIkW1zL3r6z2
gg9Al4tRbAlBKdkLZcrbAJUTW+feE6QJaPcQBFBWMaO2dg73hd3B5/lPXTfxyaFm4Q5sVQA2zgVO
TVJWcosKs5GGTFvjac3VYefvpb89S9n7bY2lBF419EB/DIN3NjXhc3gvmLiY0syjeb+Ent3zsABr
PP/wC7fTCloIl5U4oGVYX20OMWzMFdJnFrPy1jZy1HUt6Op8Vs3DQWb9aHPPJws95MQ6ySp63o2l
8E3WQoZwxBUyzz80BuNIvTa19Aw7IFR0xEluyE1dnohiftzb0J/JHq7tLYR/B+Oz3yRlEtzgD1YD
jbhho0GpeVqNmgyiQFZcf66wsSKzmEtHoHvLDEY64Vqo5GXQ56dJUc6HpYXicOcWTb4gLrr6Wkg2
jej5MaOYOL1HQyfsCAoCwv38nyK92eVTR79Ld2mHIv9cchNjA2rYtaEGjacdhVAhOQQJ7DpatvzB
7PndmYT6SE0rtE1hqzWncLinxf6IAEVOxE3PAFdOPr0eqcT2MHMqyMqqVcmzENyQW3G8/6qTcFJl
b606jyBZbpmnjpFpbcJO1tQ+Njv0OJGNZpwXIe/SP/8YVOz7Ho00Q2U+DM6NHgjOdwWZ+ibfd+iR
JcEslst848Bl5Y0K6O2EX2SPBgZk5IokePqiXmgiYuXCQII5/VPD+0TwwKaMQB2jTAjSHBE+gid+
kYDviGR5CEcxWCb3tcAEJmvozHEVADe0w8m7pUW6DUqmvhDO7w4urYz4Nvi4oIBywTTnEKfi7xmn
KrfODKRfU2JglSAQv4zlAkahwtIi2/NMcntOwOwwFhUQdNjJTjhjuzATMuiZMrhla2YXq4JG/Fkf
efQlcJHa/O2N2bLgG0geNypYgTTqIaMPFdOqdSdOzwqTpaEiuFvb95O53ftY8td/ci0b/7umucRp
gTw8nltbcw00pNlm4Q5+cmZ1n8/03r5HYGk0BzohJUSQlt/e8czuxM6oUzLDVCyazwVSBNF3hZ1n
wU9pC8M9WCdy2/B8g3VLoqcl9S/EWlfuqOFNzlR5bZCkgBMwzGyj1zslxgB8Nr+Z+AP4pkI98Hw6
gDqiTVa1xq1DwX1BrxUM0UodtAQX+JH2+5MVqLQ67v4h/bwfy3iPe0l4nshfs5IN985i9mecMpX8
xOldxanyriCno0WLUiu4qR8OaTmazv5dulXA0oNYMrsuEMJ3FDW/tmT1QT7E3lkLy2wu7SEcRiLd
LahmLU0mjn2O3ApH3mDQMbWZwLvC/reIdH4nSbnJ+XEDC8AS6NcA2rCJgdhky8bPqXxhsqbSB85+
GN786G3uI1lc5TZRfmzEm3vkuIQxynpwxkWnpVX7xjRbR7wTZW8kTAkjbdPrFJoUyOGjF2f5GpPF
nQTfUZUAP2gSCb5UISB9VVJ5S30d+hAsWZ+6EFsFOAYkY3Uv5OAPjcRGWihoWFrz16SvgoX0NXRM
QCEB/tdvfmWVhBBhqEowqxV6ELd1J1RKMp+2RhUCnZifX+XAie2Nv2QAJpOreOM46iliufUKx72Z
/cZZb0Wt1+Ky6Mrsi2LaJ3xDChxXc4XGCDX33hJQSwE8vV8LVDNJ9sAGOTkwQAziT5RmngsKbCcL
D3ppGGpI/oE2Vz0IHDKrQV9Q12vb6OS3m2UZrFnoj+pOi5xLB+EFNo8mRnX3VZBaYLQuLi/nVc5J
88QJ1tbS/tKJF9DbIWGvQMpgyzpDnutvIHghUslJZbhKD0HHsz93+OOzpzdAvG7pnfkj3oYB05H8
kSWWSNOdUG28a9msF4V+UhPHdtOlpqWI3GtzZcZgcPBmvrUj6l1cM+Eoq5fDXe9dy7PXjFWABamw
Zs7P8WOEBw/FXmmfgieL9SEfO449NzDDHveE4UVIu5EFMiqUhBGXf2H7vrPxZB56PZs1fXnrCGix
mACcFkuqHCfpcec+OVf9iNdujYrV2AcUpSHGp2WBfImNI/WWpyjbkdZwaeQPoDV3pcKaGJdFzz14
ftU/9AQFlEm+hX83s5ZqY/mmNdEeIgyAmg3Qir2P2bi0qOIBLeCZQ6sM+RYI8YKF/BYXquW7OdzZ
OEtZ3azT/sJGaoX78zErtLutuR4S5S9ou/MNnf+RawMWqKaJxQuSN1bdiXy6qnVEgxm96mvzTGT9
agZfKxfkwMnJLqCjE8k1c8ytWgzlkGSHw80kqWwuCYMC88lhIaL1u+ey8v1P5s5//mlvnNocTyLD
+UKCstlqB6aJVYd3a48cZ6w/YPJvWZM8wzA4NYh90TXxO9LmYQ4Ciog9mVA1QPzyEujWxMuwB3Od
sJJPRbLjdFsligdpmz6JxCJ+/Xrb0XMAqu6qFqA1v3iGYwKtCXam3m+K7nFsdtD3lBnVJLmSO3dV
1gMJXtYKmkppZH3hJGxs+W63Q0CrUAByb9Cd3N0Hzwg2jbjT7e2Z+i0P93uRdsiF1IFugoqQpTUM
8IPAmHLg/TMsHTu9RVDEQUwXcJcsKUpA7Ueiz8bnjsdg4gz2KMBJZyJu7IbdeOCZERa9AFX9vv7G
Lq4jnH7KZHW2SIRSTNOWw2obKfLoFX/ZNViDDMeHH0TD0IZpUm5QLapicpeOeAknu524eyY+gqrs
wSzpXG3Soigi1Zjyet4oCepC2WANOSIQvKoZdyBEmZHMdpwW5dbqk+SePYLYsqzYT/cjcF0mfsGF
g5TYWyF32wRw5fOOScv3OYqJp2s1VOPll1zt6/AXutVqoJ3dTC1zg2NvbadtNKEA+/g0o2YxMzCt
DXFWFt+gx73gY5GB9pC2V8gDSFta9xz8OWw2kUs+N+AGaHq5VcXlEP5hia+cbttBYql4I1TIRF2U
QJT02PoZi2Yp5mXjG/jXNJRXgrDvRrrUdkdQm4tlBryh5YNtKm2dKpVf+ics48vD4MjvD2d2KB78
BEQRtqfBpn9uk7TV2L0tX9/2SvgrHOQEXfIfA/ZwuGcCizR+wBK4Dg3CpTRUDHBpbIdNCsHHE5GC
u0oAX6Z5g57O2lEWrAuGs2Oo1CB+j0G9XicEUOYwB4PCOc8jEI8TqD5R50X/rJ++n4Df5Itki4JW
Y1Iu97mxyeeaMabQODGAU1SuDCwGEn4AH/0Sx3RjR3ihunnt4FC91StUfAsZE9WgryzvlLFlrLwA
um8ka7BmtSrYW4NYLu3l2SD5bRN8vCleDJ2ua2YumPL7Ev74tKWoaaQ+pL4j9KunVd7CzqV13YUH
nbnuGJF6Lg5q3VAsg3Pqngkd23utUYdce/XbthfXCZVfPVX4E0dx/k6ib3xLpamfof1BkXju4Hrv
ij/SUuAajoaH69h9prq2R2w9M8cmfRcz16FKigNVpS9e9f9iSa02qebWtDn0v+f4Q8QzLJUbeZRH
xl0cPBC8DfB7S331KkxTAWX3JIJNPFGppwffmcxhGZWdTdamhKoQ8iz1soADxYF02BJxkx6uAbK5
cNoITI1S9+1qN794lg7vWNFjGzHcXXnCea71s/a+zaWSI3RSwVtfNqCPQMjzY+BFCdLOFnNG189Z
Aprkh587fnhTNBkiFCckkKDMnIlJN1n15RQBxlFQ5c5iYPQJ1EZbpmQ32H1Md7/ZR9aEwEvzR89V
7yh9GsHIpB1Pc0f5MGpkINkaP6wns9y4nffsyPHtZOQV70QGKntY/wehoXUPTZk+ygiRg+tUUXXk
qJYg8mIGRBlayvRoMpbF7durCkfAjsmFaT1JG8ug5r2dMzdQ6okFNZxWbp3NYlyaaQ8cZJ8lQ/EH
lQcR4VeWqRBTUd3dXqmmUmxCO9krh/aSBM99EZ2mMgJxKwI8seNO45+R5ZmwvPSpczaJZ5CH8vLb
EsqXY82ShC1Rnjnwtylr/EfPDKdD+v9ZgpxyUHvOjoYNv1TkHVjpQs9xsnPbN4DXzKyGyBmvuUjX
PCmjYOc77T1fBv9wam6E7JFfuKRpfgRtr42vV4VDH3kGDLnBL6E2ta07+HEqxnzamHzqXxIfn39a
iGvKNOsAZhcnW137z1wnnc4Lyp3MMMPQ98mQQB+oFAnk5om88irifbqhLHyugTe9q/kD+iTOnKyL
0M5RN6lxtqqJ4tKLZGfZ5EBuh7txXBDvpV8FvNiiZQbn0HVXmxSks67XOmjfyJNF/0cpv//Y91jb
06Un++6Je1HfJb9w5HbjQBJVEmkrqtaHm62ps5AwEcpShv8X9GbgxylAZMVt2jpatNW0DwVzMpZ5
MAGZFzMWlnr/jF8PzJlgMoEvFcQ3rOlFgn0okJceKwiVYRs4QJx4N/DV0PAdc5hLd+7P6MYtsEim
c4xTSkWKOCLlIS3lKVDkG27/ETeNthWwA+OsgRilj4TBENf0bUXFpmksY3E7aTmy8vzYeY+cMTru
VPgE3EJ+XjKzfMAPTYABhgkl0Nn99dwJAfDLUfEt17cTX+Oji5EWfCvALPONv0qoIYTsz/sq2DRN
ma+53kTgoteE0KtHkLrUAU+GefTMkqAf8XsaM408QfZ4CNeC0bKIOeah1BLV8S7kKlkUVIquS3NW
u0h8P2tT481Re/GnmatqhypELaV01vJuN+pT31khw9hwTxoxn19FY52Zp/lzYl5X160hdfylPCBY
SU79OqkbJ18plNLTFASNWQlrvQI+FE8gmkP91qkyy5GgSqls7I4lDIceO1uJiYKa3C2HBImOYISQ
s3khueURMpbqn+r2zz2ZT4ZSpjWErInI4EvMs8HcMEUbtqlEVOz1zbktJEs83S3U9pO31A3fbqDk
NTu7pSEhDHyUunQWXpWGia4rAE4+FH0ka/teoDJ2jDW39Cm9g920Q6+SBA6wtK7sIbGlJfsmGTGm
51gPfhfi5L4IlRRm730hRTKBHwD8mvopXZlb+WEPM3wNE2LJyNpZDsm+RSgzdPWWSlDGbVxmjRfZ
3kJv+IKsdaSBpBXQZPef0Ay3mSWynNCukk+gAprorElS9Gvr/VBO41vywkPacfXYrFKZboyF1yYu
X1kw1X+PzvFUEReawCAgYwbV1tKa1j0+FC9UxWyqFU0ZGlMaL6X9lV8O5hCK0MN8xaVX0ky+W5dN
L1IpIhHDZNjjMMaEkvr4R57Na1KwovfdXyg5hCCoWzoQqRKbdAeopCcfImRTe9iDaEi1EYubraV5
BQS8v70q6wS2M5Qx8fw/Zw98PBtkdkTu2RGaHjxToAH2iT1Q1hpGbHT1kKYQxiOpOSP6U/LVJNGL
VKumUvBeiSCNr4WI8ruDOC8YZcf9UJEYk1TQ6WhHlEHR5LFHAZmI5T6H8+YJLJBLT45dyEn1xB8s
iagnA9eB9bRFTQM4NKQHcuyndFzsEPhYMa6vMxMEE/HVrOdnyft19v6T+feRq6FYq8Rhdoqr11oP
12WEoJYZwmck9eZh78bzW4pqdP0j6U4bx0iSeEyHrfPeifGuyYg9kI+9wT6xk5DDw1lj5WW31uyO
IeduEKA1ocEGwvxtiAkB9NUrMGgirDMSfLmL6qiqBLDdOrzZrQC8m2fuT2U/GYGvmoxYZUBOO1/2
nGj8BYb0c6wp5z44Y/RKf8C+QMlB9Tk5oCzG/EkbAwyR1HoWA1wU5vioGWIvQm6GhP81szFycdOy
zrLN/XrarmcVWYz0YFD0FQu7XTtMigMD2yeIa4c4u/qr4BODiHfSObrH6SCMY6o2oxlMG1tD32Ut
qtBwvRnxFr4gjQRMVh4zkTcMGJrPBx7FBE2lYu/mlon9MOvuv99yrUioLObc6QZTwrHdiT6JUs/r
jXiyDlJUoB7yTVaHMtJAYK5TBDcVCIfOeputZJAV5PBmAWR7kpKS0XZnB3IHvo2SUjDKL7+sHgxn
h9WSxatsdsmqqRa/mABxyIX0yo+NLllYBCEGMfkCgKQZihIxwe67i2nOQGDlfDxVuwOig6pshf0m
5LVM84LNn/c7deS3ZAc4FfagktjJHL8rVybtIOQX9Yo6nDx1xRzHoBEmh6Jdd0kM7LtsN7LJLn2s
9FA5ZYCzSaMYKOe+qXj734nPktNTfCOza6AJ5BShf57HSo9jADtztoCbBM0PZNRbkoFg3DC+bhMM
HEMQafXcOsM3PW3Hq4TszNlwgJTklRMtU70jXmCQevuUF8Ptbi2xrwYTibl282bnWpFLkJ69gwcK
Re7PQYyEPU4vdv3ja3msLe4LygBwBUd+kl41r+0jwkPUGNcbA/PWDSum2si+at0aq2bLFFAYHP9/
O/O7WfzI/EDQev3H6fSRRp85UGpo7hlLzniah2IlgRPINGLIcGY/WuJTPhvbPE+FJzF8s1skZ7F4
AaVdWSbFhdp5dODwxTP4Zr0GEQdmYjXwKL/ktlRuPCJNxTcWByTcCwzxj5GEldFML7wloEjhNWSY
UlCx8gdHi6Xt+KMxMhj31fP3q/kMx0wvTdJXYO7+scS6ZZdyQnAAULIiT7KDryYWrRTQyNn57W7f
XaJt1OaD3wYSiEErqHy5V1HkeVnlVI67T+yFV7IP7RF7dJSCc9SMVSQ16OxweU/5QtzxwimEN5Vn
bQP81zMuAtZmgG2TGsXHYHqglc0Gag9K0csZ2A5d4gpbyiAusTll2/JUETexWOM2wVOmnaza0pnZ
stghzXIxYgkDTiUWvBzFiRKxVRqjnUDm7mBMbPclBYNfENgxiJzrSRhhPzOQNO7IiX0WBrhkMBIH
AAJDgFqbKnbQVi9ovaaRAjd6XkDAJeawvQVc5xFdk8nZ8+MeWT3zm4kYPluLHjSErmCZDK7lJMms
TBwTLzaVQQYq/d/IOvCZNy0AEfqAx+EwphSEdHE/dHEaUw52hggM1X22G7ahQQQhscJ5C7nGEGYq
YT8dmNGi0hSjiat2S8q/enCeDk8gpBmBr9vwqAOwagSOVgGYnZ06cil3vswEuvSoXb5pPFmzzYcK
Ow32kP6TItW4k8nqa2ZL91nBBjctdL+uPhJAHQIna8Kgai/fi3SYt74gEqL82OBB92SLI2yQuIqa
mFQw6ErA5aQws/60l4zPdwMBgV7MwLoNRTGvXSnRT3Rm+oAEP7QsNfxlgQW39YQBPue6d5EhmGO8
3x7IlIIj2ux44eu3ShE3hADPZPiszTyVBAAFQ+rgpoGf9arE6Xviqd8HRzbG+q+ooJa61mc8psf1
hjSwEdOdF/jWl8Ei6Xazt8ZEQsi9lulVoeX3dGDpimb0a3FbgxA7eysFKOzy9Gq9TymvfD8ZxZ06
QQGw3A3R/PjYJQW3aCFhEBL+se2QA7L9fRvNVDxfLs2j/jF9dHaaCb0G2eBk3eqJRWu8j8vIs176
qGWPn8/geKvQbsYTtj6/Itn+0fxZV9UmaLNkoN15ADWvbqcpVKMHCbXFF+p59G0wHGg0kjPHRujF
ewDVMpEWnj/RYh0me3JcLqp3p306LTbxlYnM2HHPr1Ap7jsGgMBYUyL0AOiTu8s1MxsD54VL1Rtx
Fq9X6Dfsz5FXmeVngZAhff7SXpD1y+mvJN43LLT+Yt8vy58oDXTZ0BQxP8uh9JlrZ7Wg3+lZYu8T
1TLCzDa3PBOxVl6J2eHz/kaC0B/utflKIHJuW62/+ugtkkwRRcDl8kQme9ptsdL/KDXht4OTJamO
o8TkQP/8hGVvrDs/J80AfZ7N++NwQOgU7q+vo43CviaVsnAROfy1Gg3rn4XZSLdT6/OMY5NEUvoC
Xss2+1ePbKNmWwf8AxvbJBqtwjxIwjwl9ii6zEQuJWJZpVEAazUDo6y5tnq3VIYGf00OhIVDpxoW
rRltlRqZvwUPPxfZ5JdvEXPhMFZjE/wUbXYj4cpJKgPsaKqkW/+ChCMUtBYYDFLXyeOIWHkD0rCZ
VUzoHBPd5ctoVwNsL62Ukn7EkmibFACcP2r/jEXW6TjldhlgpCGETqbahJAXEuNJLncZgwnyUY1O
e8k+xWASySi0diLDIm0MAEPONJoYPkT6OVK81kPk7vzoQwZYGYGue8urGLyUCpmTZKJ9dWXxmCSb
6IK1nM++oyfYN03SRpbOuNNTmYArS4749P4tWEo54qMi8Px7lV0I318oHaaHs97bQRWOrr3EF/db
hcQjnH6EPCbyIMPuEbkbxpt68n2O4Qjl4OKLKwEZF5F4tcsWWzZY7h6UbnUclxPz9x42/yiQ6iB/
oqEjUXWzGcs80ehIAjLCg919b7AM8zXKQzpc0GLilLzZ/FktZEN2gokW7FVCaurKhKvmcjpOr1YD
YhjbpO8PXfxSt6Arx6H1yCjbdgXU3DAvOIRd9tEYGXJDxUIqMiBjEDoK0lb6N5/BT7wHW1FFwQv/
XPeaTe1LQgYi7O16vRlXKGdqPJeDC+3Y9VbUB1jrDuJI2GrwKwRgZEhr2MUprzcrxdvTDmNn7XA5
ir1IVyfyQN+WrAGYuYbDKhBsXvuVTsdXrGMz+ysV9xn4r98EXEUdPtMpdT6S7LO13j4gJtGej+9w
RRGhkfnvoeFlRSu6fDnn5yoGn6YTNB+51bAYmMyxysVuVi0YldXad0JHzlixEDfGm4ycFmbi+WVa
x3Zm3lyrU1Z4dFWoEvv4a4zOcYDFaNkmHse2+/AMJ7Bf/kk7j8Los3c2lKL4EnhIwzOFYMkV0g/j
4nCq3In4XORge2q5kdlS7LrrQIA8UP4up2s7H7Yr5ACDtzdJYC4jXBrkUuPJ32hbKcfJxQG8fpf+
zqbb5YeputzeOmkIqahQk2T2keL+sg8FMsPf/N9hxvbDgygCIqjSd1LAHxv/qsDWFRjpFfcUTC4i
qSnVT9lTW9yZhR7lFqeY014uQKJVonDqlzn2umwHr/uqMyFpkWSiwfKWdT5CsVuLSp6iTlk+zByX
GhnKCmz2D7a7oYdNXQRiBxj0W3ULVSifbyKu07RGcCkoLH8KwDKGVWYvO5GsPAAkCxq1lXKmwQvP
law1gI4QLoiRPzxepaNLmlr0HH0nLYIONB381vavfkhwIXUfICuRpF8U/Tfrw6HMXrwNdgpk7EJn
if2gOce2hZcEeTMg74B5QiCy0k8UQ1Uohi87kr20LEVcfMkQOxG+lo0D3v9MCD35yfyD6xaYh4n0
TIiNCRUZRuYmoheECa+8Z7E58ZQ6B3z83gEXgHMEnqJMCmd6TlrhPJUcuUOC9+HanFwun4g8gUKr
yyFS5wW1p7LWjlxP1Ztv/uHRByF6PwY+QsRdVFQA9vYtJOiRqq9UAM+SpcL+CKSrgV/KjmwH+hIH
6dkGTEbM6rnD0CUiHMGJtadLcSlt9WVP0yrRulPXNWbB6f18jnPp+3/hlWD6cp9Aitk4QEoJRJ1Y
6r+VDNoiorrAasW5fknDXznQBpkTbs6lmB5T7mY7yj9TbpZq8A5pXS78MYHEO5UEJjLhwKjDtT1T
SbScr8cXtQ9NWZGHSM3tHG5Y3A7YXyqKl6F74DOiDlNFwz5w/bP1PY1y1wovxQhDi0k5blVWmnxa
cyplyuMLbFUv81bAHb4owntyH4tMPI+HTLdFXfsKsHxGfV6gkcaitcQSJwtnc+vwDgathHqw8kzw
Gz1hlnTdCq7jJHOxxaH1e/C1+yh8TrnwDCdX9FNn88frKAxCR+FXjSyt96f6XO85U1VAwYDf0C7u
NGSk3a0W+iTGo0TqgnJU6kldqvu3SwRM56x9noy+xD3lFz5u79H9fJ83aTTchXffP097cJdEF67U
D+361YkGyQbzrNyHMmP3Lj+QQNuJGzVY/q/yXu0KXaJUgjtZUQbUA3UrgQVOUXZ+WmNn3YoQPoP/
mmgecwzVw1RdRsKiVUQDF++YvdOhjHBcVrbqwLI4EHfeCP516yIP/gIc3FOZGI/nr2Nrg0gyfOnF
8lnW1iGTeuDctLBDBJRhu15wDRbaYqVzzC2asp3upFIHkS6qrkmQocOWZ9ke4GQsvWgzrOzq6VsK
71DprntZYK2mHgS4iBldhrJ3T5lvcZVmnL9lobhVUezxI50IUyM9ce1ZtryAoCgBiaPyk8rnYUsr
7SCvRhiEQ/kt6vsLpzB2drywKMuMOAEs9yhsxAOxuPsRMPF4t2IO6k9n+Kk578GCecya5qrxdvub
Pc9GoUwBNq6Ejhs/E9NExSRtMKbLF5up9KcR0MsCO/+vNdtUe0ZN4zqglhUXxrERsFKAnSJLSIDC
/7DmLvVxLCbJPh/Igu7w/50uAVlB4FDjtUhDnEhdMLY3xn0GNi1FyCo9QzViA+iwbZmzrapCM+I7
eN8YsJgF1/icldI9lTbCBatuaJ9P20TStEuTjT7hxcmXUdvQDdNGRqAE1s0VxQNacXWD+wDkIR1p
X2+xVUbo4ZES97ojLEUcY6AqJP2K2p0xpyhOQoBWzOnxXYchq3IOLHCZUCyqiwSRtMzo9f6QwBic
+Bfa3A7mP3uKwJcdt2Rnu6S3yb/FnP0nUBgW9hk1KWjgBFHJ8mnyQNmwHldHxgIyjhI+LsjYejl1
AARVDUTFwHyzN+X5CEBHlD/zXfoaUPg3lcMyK54RyfKASC9hmKx3tdJbFcZsI3EQL2ivOxiZnspZ
30i4io93fKrcEqf9wanJtCgTmFagQwgndX7suTlyR3MZ4Rd858Af6NBCyRQIJrCOy1IIKwu4P/F2
0GAYfAjH65pyF4FBLotYoRyL37kzxyDuLbk61x2ml5jonD0ZeCKOzJP7pbtiN30uSJIHeIroOhNl
kNK82botNT7Rzd/69wnWGtEpKVlFEmgBFCczKbV6e5oazhixTpIR4JtmSW3S5XhGh+w52SVP+l1O
CT5M7HWshD0Wv02Cc+iYBwFSM2Zq2P811IJ/5P6DGSDFzpwmYnDWwy+JUPLGYI4NZ6eSkRV7tOhi
lhnwFPTiCcuq7oyKM45P1BF7AARYRMarKApxw5limdmiyhAm/449BMEOK3nSRnRaNqQ0xBYLG6cF
124ueFqH5wTeRCDR/926fftfmdR+YTRjuFC8flLfeBK12gSv/6uLG8FxEySZaq4/hVbmf5L2hyN1
xDuEPhy4iMe/hdznhp9WXGGlx9h8mvD5z5KVuBnDlTBgJCeWFbvUcluf+6Q+HOHMOlyWkdV79sTv
PUA3WH1hD6rMRK5HzyB1BZkd5pTSQoc7MgHDD7Bd1QNWOki9HvJmFVPjQv+Su6c26Zi+S7RFTlTj
GDaP1cGvMcmwckulqMSzonfFocRAF7FPL6yBGka/PHE3UIXsh1+jNkO1UXCMI+Z4siW29Dzp9+Ao
NphDvRRugiKmVzX9sLDPX6PY6wbtxdZxZP5yS1IAwp2PckfVpy6n0vfsvOorKUjB+l/pQhdhkXnT
QG1VzRURfgKkK3TinhI0wDyBlpcWCCBQNur155LAfvDR2I0Z2Pf+FK0PogrfsGSiYetUpTDhSoHk
F+CdwcxqnO+fa1g0pH8LT29OWL53XjuFoeDeNQuVmxjOjiSqbrr7Iq90tgW1UoILzP8ejmGdnfJb
qJc2Bsd0Y2cA2of11PtFEA7BuVe/9QoA3OoFgmwvJL/qtz1qWAFj3LL5pyik06jrhaKGRsmfrC34
v1FDXZnPvK3YkQMoG9MXehneaWdNuQ8M2aLvHxmYh3fhVPCLmOJ+NNytKhN/GVzSkRExkg1d6M29
8SlHIWNCUdy3SQ2Jx+JSdoDqMg+t/K4JdfXytk9kEKFfq9csWwckiW2UOOxTYjq1PQnNTNbv7Z78
HE9XIXSYx7ytcpmqjyii/VAsKT2l+tri0gC1junJ9g27kP6lK5mL1M0Qc0V+9ZJQZwsZPRvSiYJq
XiiK2/m/eMhkCgiw7AB7Jlj5AbGzBefrbKM4ZwQkdvAKEsDfbeTKiF+p9aTaY8sM4M9g8xsrPOGW
+F+GFYGfjlGls6Kt2ROmrGZh4NFm+ovelaUuQWMVr9Bga6S0QzBnhp1t6bVhMgedlDGmis2ufWCN
W7rGb2C+u9OUxlieK7HCb/bG2SMcJkZxV98dzkzOzEdN3xt2ZzZSA5oEg8R7sO9q5EfrPM5D5NU0
pj8nO77ya80a/3xRqTshwyLHgpqb3aaCUfk7hvYdQBGBaayz9Ht7TMS+0VUiajkIdMvxGHDDZ520
ce6d0iwCvA87xc0OY3yNZb8u8A0U5hvQngRImJeca2G5fL6pAxqxnHOVJJe9KG8odIrVoMnh0ppe
VplsbK+5DVm1eKp8jTGQkKfj15xi4EnbNhmaF7zu7dO3Avd8Ub4MjNpP1u3WpGKvnpVDs288/qvv
cmxq0RL9cEYXyimFS/d1QB6d2xDBmlXbOdxfFO02iWQi/pDFIGoeNSfIaotHKoxEfLMZi3PasfUu
STIt4ZIZXFwQaadOh8RDwtfQ0QT5oTTVMarJrJdpZZK37KR+y0C0hobpJxdN0eJZAz7ZARSf4py6
2fCwOmWNlnzTAI2iLV+yfn/z8E0VromLNBNkt7gU1FA6aaU2eYWW59fLCW6r5PiVvmalhKqcsm+H
i/GU0fF2Q8eyZ6pMMfTgo18q5y2SlR8T92vafjposq5s8GAjWBfoiJX1R0akV3jD/eMydbdOT120
7n0Y/PyprwtJqaL3YpfZ1a8s/8onST9qYaPouU3ZpYKTGvhfjMam56ZVkUkX/Fdtk+E4DP9ezBXa
YVgCNitWaLyYXiIKbyF99mEHgv5vQPNmUR34sZRCKCHi1hqRdYG6hibhXptlddGSQIx3Rh22xvos
NXKatNotKSiZ8/F7CnRgXVo1hv7T4osK/TI8uckQJ4XVwl7mnfzSiLj1tW4Ba/6bBWkLHIu3v7eL
LyBz5JvSAW6Oqs5+S1ColnJjAfRmywmEA92Ak21pD0fzcbJ9YbIiQxoC8Z/LH/YPcWgmWpzLRVQi
A/+bpDeeL4K0fhub0iZSW9EFKbH4qzWoquXwg/nS0qIxfbHKSSv9XTq1PaDSfioIcWDGtsnTLhTE
J9pSHOKUKLB4i9OzAj7DUr9omqRHtJn8FUT9uIH4Ua2TpildRSVE2Mg/pdvNWrb4CKZTa9i9lRtW
8/01Xe6MjmtVwr2TMTAaN6rFu4bNxyw1HRgRCnc7JTOO4u9In9DOanpIVIadChZDlRb3jCgOk9My
cfOsTyXKcG+Z+zSpC0fvsy+HqpzgbMlhJJ8ZH36x7KiAlqXpChe4bJXV2Rdl2gO63Mi/AGqrXBv4
gSFFIRjwe/nHyC4c25AlsrcJP21wPXOx3KvKcITPm61YRnNbjKRYPKCRLbhxSuuouGorqwP6Iopi
Rye8mfCq3fVsQQht+m1j4UdDO+cIl5PALWbCxUjQ5kApBld+EQVZeLkTnHvCCQ2G99z4qWYpyFVS
JAzdG57iwq4QZOVRxbQfF5/zfG81jaCDexLJpYle1nsRWeZ7s8ZArAmXmSx3kTIIWwQ/kf+KzeHj
Wr36Y1X+QMozpEhdJKu7kGCw9p0Wjte5rVtuJLqKmbkjJ6pO5GBh+bMIoBmRnxzwGfPBJ5YwX9HW
PfuXEaH6XV4WASP4jtKSXQ7KRV5neVB07lAj/qeT6ph3WHSLowyJFXkiQ76cxMdZ52gv3ED0b13/
o8XEzvE5nxdVoPRlJWjTWbcjKyJnE10rW18qlatsYGkR8aE/0CmbobKfsIU6t8wmsj3bV6J/Ma5X
Rb/ahG848AjUz72nFGGygFQYu0CyG6Ju/PMpwXAMShtXbRdAn/BU3XUgjpVb1FFfYgoE2lGk0gyF
bRX1z5eddqQESv8Q7KoLA82AymTm9NG9pnpczq4vJQPJC3ljwfkkg31GQUYqEMri7qChDMJttPng
uoScEpT7LmlQzOHEdsjJeMprldZuZx1FFWOoPIszl5nZNJIvibGwM7G8iP0FGBIcnKhndpsnMSAE
mnYvJ8i563xuiIziqb3Q187EhxE5LD2T6mdG49mZ6iSSz9+f+M+YMbN4PNGcl7yg8l8ECxc/STA0
4CWKP+434EuPzTjousUSilZj/W17Xvuhlke+jIBdLSHL99RwbLzfzu3t7bT3LTRIuOY7TWY7dU2h
g7de3lcL72V7873j5W9e0eHo8rO0sgFqutsdb74YDYe8GED1kCs6wZAP7Q7qEXJhnpObTFtdIr3+
xWCjOtJZA2h6s2qNTweK//EDPBmjbWIKqGB/8CRpWaprWQxb6Y4RgyXJ8oChr5A9HjJrxKGuY3xB
TONxexPyo2wXYw+dbSfuLPN3bah0vF/6tO1kUAN4A9JcxBLp60cct7Io6+8PcYqnh14U6Ne1OnQf
HY2WRrYh5I+s/xCKW/FR2X8OXZG8CvdhrSfdd1vX1u7RHohqAuddlsE6qyT+Dd840TWTZxmiKeQe
rag9pc+TNuGwbz5sF4I5d8rQbFyun8RbdHLYkgfMopQQHk5ktJ+NlKF0qArNOE59Jzdx6xlIoEyF
kxACGNIAvvaOrCj8zhik+KA7XKoPNNPM2vAerbLHuSYhRf+5ZVb3YJbXtQtYbfcnCevsoPXOzjW+
40+2xUIoBKCnMlMrjwiPCi2jX/H6hfyQxYIw3Phqxaz5h/efyMMzNOdzQdqi5OSfQyxNteeLnDkh
QKjPQqseGC9eN1ML6v/w5zznz7lYIc7aFIXzx/hirSWwcOM0x1ye2/8d9GRHNGsUMhV/p4wlOXr5
EXiWqrjN2OVSnSXDyBQJnvdyUhVfV743cB2/cRXV09Miu4D6I877b+4w3hkYP2eV9THNWqHfo9/1
HdnfuxV66FIYZfv0ImJ041b9UZJKuaIUQUmCnb0CsmxXU8X+sDCCpBBbOwMZU58ZkrODqHu7GBKH
LKpfdXLakv4WlFUWRRPmhdqW04jGjwpdFYZdmy9lZK3zE8b+G1FVNGSVGLntmJ747p+z4uhxVxYl
H99G8ROGYVMW65uaPhDdtJPoPRVr+PqBX9j2xqScu5kbuYqrxXNzDsep1rtpJVhoP6KyNhVwR8yb
sqzPADHdgCa3oYkxRZbcj/Mm24QflGSuCjz3tXHgq3oLQwhZaJzxs1hWEBsrAl7dlbbfF2QL7GUl
VXuHQ25xqXA911uWuK7DcHFmtQAKhSXYdS/Edk8hAFCxKsoHCTNocMoRu3DjRDMw28SpB2iBJhQG
YPiPc3bPuhGPHzDCsLuPLCXpF900EvO7YTk6KXuL1mMNWRGrSDuXncCp28W5jWOKI3BkM48Pt6tQ
3blkSSR6C5mUwTlDz/vD6S8y/EK2FGraRb3cwxEyqEqdlarOjJlZsG0+eAZgRjnghq4uXCIrNHD6
sP8bA9ulwYX/I1ncdTQ6jP2EB7bmqcXuK/9WHbsygXaK5WgMXzYJdboUAya1U5ebd1oceJRJ/Pp0
++KCwh4cct+xn6ci0AaW/3QN0YZYicuwA1RK07QKoc27JqGEm2Ds2Ox8E6JksOa5kgSlEOKIgqG5
QmM+d/1iqt8Smpsi5eFT2syijhBQGxTvLSzqtfXrsdO4LYJ1rQoqRU0t4yM5mIdReAfK4EcMbR6D
XIwgL+DwM2QPJF1wAV/VfkAmLG5tgRJDyIdJ3TC424tnjXJ4JmUQLczD4EyeEKtWbU7hxrFVJ/Vk
wTXy0VNbX1tlf4wU8T8/d8xOiJQHrwCwB6Q2OqCucyCbp8CUxfTfHaLNk/h7NHDYc/Bb3lcKnnkN
lD8ZIXNf6EBa8nkmSs2OI1FvRfp6tWN37sVbGqhCKgiNsyRCse9TT7Q1v16g9TCd9y/mQxlBNOLe
rxEcl7Q+iKGRP+LIXOgdgvboEofvMWjbvhRlkrfm4BBWSjNabSAV+1zTAcmYQaiBWhoIMwNJRmKj
p28v74pjQI5bmyLo2xVYJWdlbbEA6GxD94YxHBBR8Me5SaqzWLRPtXp3E08xAYYKp3rCWZQvCqKb
wQt3C7XgzWPlXilyT/AzOAAQR2Ln/dXsryu1ziM19apmuwu4O7OTXjBZtK0XtKfQKGI57lLk2Pic
IhN4T4JaRydigRJ+AxsxzVbddx0q0Pto3saOecm1AZu8o6nPUCA/qau/KgS8Vyl3ACnBExWBA7CK
DGVWyVJnwBsFKj2b/wC0AHZluCDadz3fAxwiPLZs6EmZanssXaZLsRiQLWKRjx7XbGPT6mmGgZz4
gMGlA+aMsSsyjiMvpUNZdKYox1iBuCxoC81F/l/R91bZKc2G5ZIJNh2pE059d1mhEuBRjSF4xoQU
vMzqpyMqbCD3AoCYNWMizbCl1DOCl1yk6IvJR0P9N5VB8cv/By6NbqxPT9+dQ+AtQuULc0tlheBj
WCblHozUtOsNBv0m6zaMlUurr8VYPMwiNfUMYMC1baJXKzOOQJM36LF1VmbGgxj0aYTsY7ZAPire
XufuRFIROI/xn/K5SZmwnLDm9I8VVDoRD+7/ZGFYkZ3iC0T5iVOi6zJoOrgQXKwEAnw6MZ+BzZ1X
xJ8p1pIhrEtn4hmPH9DjC0Nhs1U4iSjMDvfhqJMmgK2HkEHUpJ6tT0zzzp/Ah8vFL5vl6t7ewfCA
WkROHN5k888kRzcaiQysFg264aN9n+6YMf2a05W4FRgJykpvnsZQTP8iLV124oMNCgGsHiBSEBEx
9NlxsATDGoBfBDgoCrEIzay13jIpDmY7oY3hWNBCGZwPFb3T+ldR9EjOhaJVsZKCLvVb4j/XDbg1
Y51A4pn2A0ZGclzUQHGtU8Wd+mBcsdKdTnJF6Mux8RD6VPcNt34+T+QXjjjlYtLVHAhNfgRmrQ1o
9pK+I5SorcAZN03Rg51lXr5OndRl1KCSiit96xgLFWnBnfI47NDYDpJKMB8Lp9QfqLS9zYYHq9uW
3E5G65Yu3jhFr8kMb1upC1P7CXIdD+t9v7gVh3rAhBhZf92qH25jXtOGoEielmulvxByCrWC8T4W
bZ3doNeWo/vbcULwfdBH+5mrxnQfz8BQb653HABKpZKyNeC9IKoFyj0oNiGflgKLDcIqkAOV3EYG
LKXOYBd5q1SqC4LmQxapQyDpny2/dpJGzsa9GPzOrZmDADfqy4DDOeZ0uDuMEGMI2IUP0CTUV70B
EAketL+PTVO35N3Xbm9KAeI4hqJDaZu2rOHM2KAV4yxN0FrP3/038kpYPxUMOMgZRrI96RPH4gzf
Vf1+kgqoEhmGaLjP2QWz54JaqAU0pvOsQpU2G5oz/PtR+hExEB20A+t2pQjfOuxIFZsRj25O4O3C
prAeRT5CYvzsFNRjqYSUF97mfB0jxU9H7+AGwOFTyCjTMd2IWLsuyNP83mWafi2ky8mCG+9k4PDK
SAC3oHlDcxeYWLjwfKuXIWvzmxQQB1pENvveOG0RptMtVwsr66DlZASnnTpS69SdunO3yMwzeYxE
x1aslv80TqssAla60Z1+mjJoQbTpeATmKzT7t24Qq8PV61gq+pW/pRMJU6LoQXdr6jgQ+LZ5Vf+D
Odof4wV+jp4MXcidIP1T8H+L8c2eAMy44CCMAYoLMRY3GT6Oh+9of/mSf/VGrW2TGjntBr/8cTPI
7oCTzYn/LAXNvcc84qgqGZ4Aaus9gPJiaS/RM6+K/r6smNqMfC7s5X4EhDKc+rouBXQefQdG9WQe
1LPkwPE9nWCSvgPsl82yiHP/+vf14Hey/UB/D4W7IE06kMbKnsYKiVcGIuPApdVXZRL/NEwLcU+4
lADol33bQjqSGATfneqQ3poLJTaA5yyj4S6iFHdnmVF4UehG/VqNOSpNNzByGBfxqX5hscqTIApX
cabTI25gZhcsu5EHZttfGul0P3hBNQGD5HryixOMr6pwFqqnSKQbyc7pe+c7UctNZzMdpJU/tnrs
3jwZ8al4TmikoJ+aCR60w2CqjUdiFWbi/J1sJz8/aO9RxpasSaon9UEcXXImRKse76QuNfvDR1QF
pzmbjZ9jNCkUrn8/sC0kQYd8ztT01QJDXB1Vm0hLrs4HtkItN8G/XTcABbrwRkMZbpJTNIUvMf2s
YiC8r1Ri6KyRA96Rr+vB6CiEyE1mXufmiL0Im9xES9bGcF0x7e8G5VgJx9oPUrVOfBs5vlWai7sJ
xZB6GJBdfJfk/sd7/Oius/d2CUllFPP1dLIcTTumbwyL5n9XsKx1ogjXsMF3PN1mRufJIuTZ5ctF
FoWtaOrXknrk1jON9smMx8f2z1eZITb7DLbB9ye1PrlfC8rirzgIdf2XKPEbQImrWfgfwz7ZX9HQ
7lzQvLysboyl9MyJQaQLWn3GVKj0zIbyyXEOetR7NLvdw4Xw/UZmfKd8Ehk5F6Jnn4vj2+VZPwZB
G0gWGlMZHq3jpgxxMnTX18CSwCmNOasDklj225Ocu2I9FipCdYTBY6LjgrvzRPhKJ+NIwLwUy6eL
0Ln8CaFY2EgHgbvegD1/Rl0XbDlWB72tmR92lKipdLhCO+bGnKRs5mGHg2EeQv97mD6VIEeHwKQv
+j20kyXvC7nkWMxDxa1CcLgTSriQu1sVVaBQwqR/zilQK36FA8yagWjHpCP1mzEVupV8d7RFjtZP
fdcsVj6de/OUFnYsb75tQes6oc8MnpDRe2pp3vDnA6EkZZf72770XFlxQenIpsGNKJEoCs6sWrCc
mbYBDjZo1bQXiOGZEvSivJy2yNMhXCEeSdEH/HEiMtfiqoULvEU2M/g6g0ozx7zTYr9oOe+5BViR
NJQGNDUCDp++c1yQMO7v1r+hwxAei7gW0jRxL/WRkZ5xHeZoHwaMnA2dijmMN549V3ii3blaQhsW
qmmABFT8iBCnCLyW7Yy0cB8KpEjmAakvoXr/oITqypCi2DTOPbXtC8t9ucR9S/C3Nzrconmm+UaQ
idPXh0qvWNwqyZxfTp7/nTuzG0C/6W9NhBDNKn6q+uzn+D6EpVjvPca6W0yTed47LzaeExBBZIKL
NiyVC7DJKwWjPx3G0DqW2+y/0vJ0OY+qyKGWKYur/LTjlZJUkXgbU/yFyDqLNihCm85miQSaTvGn
nN90tGOudgae6xLzBzjyQVNxXUmcP/NsA1QwPvw9Nliv+KNOWK9qv2ZrtdFzZCuGZMNTB66ETqBn
QPF0TI87b1WSKtkJSuGhk1iF/tqlsPk96Dt2a4yN93qoaU1sELzlS13gpE7vNP+FyFQrvPM6igSW
Ua1zTANx6TaKV1Obq6QHAEEyrm9zo2kZPzzVQMqZUzCeIxrHtHv9H3+t5xKmKkfQtdzrY3YqLLZd
F8aoVE47yPhcqzOm2DvG8ksnU7CvKJ6Zq41/v0HSYk/fMNWvR5moQwHvEusK9Lut/xS9GEzzKo4K
10tZjy3g2vuIWCz/M/yBkASSEbFPGE5VXrcwG4hSWwf5c3Oz3fq2shJSAlDF/ou7JnjLx1QRuBZu
ee2RtnNEsV6+8nEzrqyCOAWFdGSJrlJleNilMAs2gjb9jrfrR6QQJA8kwI/Oeji8BtjxCeX3RFO0
CsppCHMQ4YonfH7SvV+zdo0jZcwy6pmnmQ0JsSW/tbBNCEdCUB4lMJeqO+HI7BOd4TUrZGeXqt85
aJOAXcYFsbqbXiuMAbfk8OzkeDWdKkgtkpggYXx5AJUexKqij5oHb9Lo4A2iCQBF5kWzr5GJBWyO
WypFFXhkqGmNr2cWgjKSbjkuD+Yd+YAfAmwAC176mulhxphHRfYK6+JGBYVS1RCw6Kg/xxE+B+ht
VxBExEGVb2GOg6wyj/mgwAHbka567y65QvtA5QIhp4E9yr/bpecfhzxPxFItDOCwm93AN+nJrhE+
JPV47iwD/yoYJ12gCpEK5MkogoRbRYvaLQLrxYFlLg3i+Mzie76rr8P9LBsmg5In1TeVbXB9vM7d
TuAD6sflefrCIPQvSd/nQrV/JdKqE8aElTxInr0Vscf4aT/FAoV6RdzI4GrLbhlM7VddBR36ichx
LxUUmyT2ORWhSHOa6U+wvFUWPXtGJlF6GmwRkwBLczPesaM6FBq5zJSN+1IDrrgVSqB2EVQkuAW7
fd9xYYUoBu/jkdxDqi5+ddDanSakZHovl0ndwaQrsgyJiM5grjqSERbzFDCls4GHydKWcrSIzIbi
Um5Nmf34edRwJ8xh161DoEfkT3s9G0lurgA7k/8Z0bgDiWQm4GzJZ8fBxPcAeuuaNdJ1N6sBvvY9
glja+2ap9ll2cxEf5dxN2uD5Uc8GNSXpoiOVCTWfGhDUBkLKMJ98yr0wDAiP+nPvq1zxCchVc5w5
eTkOTnYjlSMrtMjvaqb9tUPcztxpb+m2nEYKcnpl5MuMMhldNYIlO37TWk6HtJ4k8InMMMuqxVok
DyNOzYDlry6PcBqL1Lif4MnJd7eDjcLzUNcQmLMrbWBMLI0tD/2yLejrSVWm9e0i4orDasIWUb/H
2NS2Ksy/sgYysuM1KWuP3LJBdMf95jLOwjfFeU8xhVurIjHaTjDgAwN7l8EZn83r0jVa3qV2pR5A
6BptqfENXgsNV4IdVs4NV2tQa3kE4YF22FvTHqc0DEx2lJqP++OxaMVhzKgkXYSpPzd+LGrkYIZZ
jPIqglTKOoI82IHqyIeiBeXrciGYP3kc3zlwcAh6lxnFSk3Uh3t4JcInCZ4JovJnSrqgN8yDS2U+
dxyQzdBrBYVtG5F+pY0vgIbQ8CcJaIZrkMH+zayL2DrXXi1jiFgTplLiV/2Zoi6afUpd7nSHlKOS
xHSNm+hCUtZJ7wa7BVDpTQQ+HyRJkwYnw99Y9IK4bOXg5/M0ZmxN7pu/m6kvZcSZRBvwAsRytZDT
i0rXeELilusmLaiyFqAVJLBzyHEfE1xBhYaTkoovBv9piUj6kN4/4sYJ7cM+F7ZE7ZhxIj8XkFK0
idKVDDnGL0WzBEYpKJWiJOd1JDXDMYFqrSSAOFenEwRa9t97GtzZpu4CgEEvbq/cObIrR30O25TC
on5JALMjpk/XdhxBnlY4Y/PL+2udp/UT6+2GRLhvosY8SSNefSFx59PTN7JcpSqUHawL8gGKxucW
hEdIMYeZrpeFPlJSyUQvARUnSR+keGeqUI2wCSqLLfr87KRChFED+WlPZ0msGaG5R1wEOLVRaImc
lhgVnC7Skg8f+4ZSE/rdu0FbAFtuSGEWbaxnN6POyxeSJjVyaf5lkketHYxMd+BJsS6p6Beht7FS
yBh0faH3vv041ozT8dbszcPindYI5JMILAuZrxWMCn/RMABDIP9Rg7BjeSiQlN4kXdCyFuqhw0s/
EvWnysghJ/Kq5cKlH+pgCJCqZ+RYmE12Ql/vyPH397QcNEBFzLJue+yfbU3eM77UXWfe/HtChS/g
aPq1PO4Db2V7HAGpXljOlgqYVYlKWJWV86m4dFAOX/d/NAeIvJsV8jrDIhycNrlvZSS/05VM9qNk
aJ0RTuL+eEAVDjzRFwShls9JmAn0s4UcaxbOwyN2NQu3iPUJ40/A8fKoqvBocnN9laORhfnL+Ngd
09lh52B7iDuc5+UTnJjayw3IygAujNt85G17zCgvB7Jv5S8uw4wzBWP5oJeTP92SkyWrLxpk/WyN
/kr7rNWZApq0qkbjh35x38NdqQqD1r1DR5ZFUgCcNQaHeULayq0EU2OFtTiuogG4jZj3MgLkEFc+
8KmeHEB0KgpXUuE57AfatxPnOauVAOH70Ro+jOON/wFGZge21YOQ7wgfXzylLk+sZfkgSiQ5ap2M
oHr8yGgl/qT7cSQL6/mw+B82V+gvbON0b+5FlwCSGc89gAIzEavjOlPzV5pJsy4NlRRNevX7mQv9
ZlpPbRi6lNh7xTRLuaCw5zGwT0q5bNj1rIw2DKUuEaGSJ/TaZU/YkmbCMNFSsLFooKmCu+A+/WZS
ypb9bpgR5u3ztbSEZX0vVTkDgcK+k4eKwcI3EDmQFuM06EYQhQldXIT2+4T3osnqogjjlmSW/sb1
5GJCCWjV1AnU8tc9VQc2InG2uUku/GNN58VBYDgMN2Qf7R52i3hjsCR8Gz+kFIxUv7jyUnct00xZ
RBXarYoozzyvHrr1QGZPeJjggqrssdTDSVXGidkwBkRnWT1CJd5NANW/vrujBLN+e+9N9z7fpHtm
1tf+ith5LIDKfAJtbFOkytQmIUFiJD2R1p95agK0VHB2a/8JPQ7to0KzUL/NCbUeHdFga+ylqaGg
U3q9l8sdeTuvnLA0tQc7ocgK8KCfA4LHGawBE5A6GbdD9P01krYYTlsSKlckroweHoO8I2X7ADlX
KCvXEqITSrmxDvVh1pvK96D4+hKQWFOvTNKDwiMrm/wNyYPmslz4F+004Uy5kDoZrEWpSxBZvhdd
TNX7pl2K5B8rGt0vPZYtbX37rQidUCP/pBW0WGQjRjyZ6wjNYOy6rkLZz2jJlAhZZnbKIbd2d7zR
tespgju1Kmk6VHbbHTW93wgsw0bBA+4zJk+gGNWJeF81MufJtQbYBhLztljFSrNSyGJTsKSk9iaK
W9ztXshdiw+GUqNebhtLoSDpYKRCcNyfxnJW1n8i/h1ZhyRRDpy8tjEW0pHUAuWznyhd6DZ1MSHr
C7aRI0elrxBR+EXKBcebdXdj2rVUKat/oBdH7rton0D/7saeSy4Ev7HyFuE9bnxywYB4Y8vJSlDb
ttXbgmgt+fb71Jb2LKpAPyl9TZ1KM6svFo/i3byVZlNcN8EDbr7SDARlrwOzo9dDmbCFMCr/Lcmm
brVgMBMBzqiivh/6YJVBZGWs2TSu0/E6o2fPpChUmjSNcql7fi+GGQ2L1gJ0hFl2pyzaE4skYeLB
/1yMw3IUJyZEh5vx6Y3SgLeLskJ/ZEpuTt5Zl2rLJSruTThEEVxlmxNvqi4E7qW65mXvS4Pps4kt
7iKOvrv6YYDg4u8yrYSUP0W6sg7ntR+DkWLaGgPYEs+/WLvy9VfXt2LsfjVeqXDZvy2/HGi3RANb
k8WmL0PnI/C0EukbJMX2d31UJtuKwYz0fW6qPEt6owQG4b3qOn7tTLAonTK9lzphI/Z8YmdnOHwg
VSoWGeeOIbJUi8WMNQPeCoCV/sAQfxbE6NVQV5kAFEuERB/VhPQp8QlrFbCaBRMKFlabJmLfAf7/
lrvAwuINcZoHrZT+DNv8YoOOGHNB21SZQ6RSIiaJNY7SRz3ZH4ShO5XZxQSudqIHouumhxrBWuNo
YlCe0yRcodzAW9UTIcykqPSDZjMHc4DD+i6vYCyHfkoeJYQT0c1+bE6jlIFDOBF415JhaI0SFABI
6IoEhtkw04Hz6HM2p10bBfa5kU+KE/26EUPOzLm5YIpuAW3VbhpM+koZhIyO4qv0jUnG2EImFJxK
6dFm22KmQiEzLaRYJPTO/Ea7+9RoECxP8rk9tYG+h5NkofgiEIeHFIrYegJe7qMDKVoS80E93YCz
9j4KK5tESqsPspBHOasUhyjOgeEtvWrLDcE/KVpekmOnObxIqSLV0oFe+DqZS/TWTrakOVoXbFBu
7kfA6XhnfFTM7nQGDBjm9lJ1ZABURINYoPy03yjGBly2aeJp1ejeCr6jIZd6T3RGFsjOxBblTWtj
76GHu971qNqv08s6/PJ5tSgnz0DGyjKJv2JmLyaOIGsPz/O7hWyXu1ax0Wgm5AAEFny5ISKri21G
JIqha3Oq1VwWhs3snDFRyygIYrR9dKmPOFfuzxSkwKhrIjk6PIz8JAHLaYz7Ru5rVlryOyDJaSpY
ZVu7GGOpnw46J3yw7L0i4PUXoDCPNNXcLvKCGqJjPM3QtotwCuGDilXYKbm/6swjbB7oYamA+46s
dAPWuNf3GgEIeLawo7mRFlq1yp2KspAFCACQKicnxRV8dwnNsn9W4WTc0oRxYS/TB1QF20L8pJMV
Ck2tm2a9SA1MRRJGBYMfhv38+C08ipaiXvOQWyikrdCw3XeaZQluXz/fRy28r7UhMIEQ8iAw7ALS
fzzxNEDZ3kMPPfmN0lrYanx0s+bsOek901mS/RW3avwf07FEFE3m5r0ofmdKKAfmhcU/qY8xb++u
W5wjgDmghlP23kERJrM0ZfzHQqirU1ppn7aZOKEVoKHD0ohovXAQ8V+4v8Eb57rNSwe35WOO1YCr
OVPShOT53XlStD+rdho96J8vNlc3/y85csRlf/FOD0D+yNEBD+PU7b82BoSqpKFCid3yLYCd0tHZ
DdJ3W1YUaVB6Ckf2XhjdQigmA2u3Uw41RWxXKIjVPM6kGXqKMATlY5LY4WvM9vnpNCX0rmNRTMoP
AEwZwC3CaauyCxrkTrxX5zwwUMMqVkNl7sfT1cAQH++JS6jvDnNuO2FB6Heph+OoF6cGV6Ym1S2t
VH0nIL27yNXy3O9vwpj2WF7dq/WuflzLNRc55cG2W2eviK0jl60xkBWGOt7nuYyJ1qXjw+5WptNv
cDjxlGIpNjkfXaDeakrgt1hpubXsOCFJVmcKO1He6M4xRIzZA5KYd9TwPyoFYbP1kji34jw04AgW
9ywxjnVnNW7XcxEyc1Qh0stTuAARtTcAwTnCRILntE/jLbcB92CL0/syzKCjK7MaNLgMOLKi6Hck
qmYHc69lNtwyI59XEiV0k3NHeutt4tDXkBSJb7saguDMfQkhsfZWJifxZkTLnSmC5+eaaVqgDoPm
ZuM4pqCbATGAmg49dYU6exxB3Q4yEAgKVbuang6Cxn51rZiRMaV5bwc06l9qqz4TDpxBTVUB0KeV
PI13t+AGBmBMOAuq6ysufmsOf07lK28Ekfk4vVumCt8HvqGJYn+JpPcxzqxVz0hCuC7OKUnq9Doa
qe+2bzOuLFSEW4SN5KInLkeNKimDN3GDHw+pQ5HSe00WgrVn06GtemAE0uxON6hAUNsr3DzHxll0
dllX7Acw1KkZ4VqPTpRU8ZgYNSbTGW2DD4oOvPhKEKYjA/G3RNrBnxyFQUzaZ98dY1bpJRmD+cTW
+bAC3xu2qeKg79ukWLk+UzLD16EWtqwzWF/CBMri3EKQmr85xv7Zw4i+L74h5b2ma8pbVZ4BFqUN
a+y+x1sTs2I2mzP5VLPWyYiy0xQBef840KPXgY6GuhQt+EnQ33/YKoY98M/qPoTHM+1vvdfZLrOn
9pSykjQdqBT4oL79ZLUxUZg3WoiMZCvKTtLCsaMM76x2ooCCPB6QBCBu3gYF2oIu9A8ZY60Pg7wr
wmnA1fz6aNhySPg3SjIP4MgFDAc17uDSjsz3MESL1b+gFhSu/IrxxYKtgaTdt4g/NvbwujcVfgU7
ouWN3oBti/bCpgOCji8fM3lulYSAQF81j+2YPzlzCoylVKYdNEAxOdCmrPaQox92A6DxPGsJK0W5
ojk67V0Y3m1chZ2MT1k/6sqM2QZALsV2m/sqSmc9Y28txc1+0ORWAd99ouEPMPirYQCBLOckY/Vs
IBBA4wwoE95ULTxgijJMtAZ09jyhm4AH6at/+1FsgpFDPSWbWV9eo8wzDB+ZcOGzgWUBOfgv6gHs
aVK4IYzfpoF+F4uYH3B0PFWrofcYwWwKCGEMCvIsfGT2GKqK0cfNIKEw90tJYVQa0BTKRt5665t+
lWmUCrtfnWKRTMe2c5eIXTR0UtJ52BIYdYj/hSwiW8wct7x5mPwKYHARduSvMv8fm3RhhNHnP0EP
M43hafqTw3YD1fDqONJ2CSuidI9hevvfVNU0TCjVQQzHWSpSPp+SnkF9zy9pOha/ygAb6k6J4mxP
jCLlUw7AGBTSZXPlqtAJ+JXmSPmFs19CBTseKwiN5+hdImsxAbUou9HD3B1pnLTwD3YMifCfnwIN
OH71jFbqHv08svYPvDetEVDwXZk/0hIrrQFOUHCksKfq28uLfH7QvwodgDQdlQTQvL3IVfjx/dCT
g9oAZQt/G4tVFZpXY+1pE11Mq+tcJ9Ig5VYde8flO3vqPiE05GCIONcWTo5O7nyI1HdVaBnA5CSF
Fo5ELHBgkwjj5SECmab2aMy7DZaJ03TH79iiVRNpQW+Eff6GAw/Qip5A/VgQeUR06kXMTreJ27qB
gdUYnqP877DY/STui/NHY9rE2ebj7Rsj+S8MilRK3HssT2lUgLI1zob59z0wbfdgXmBN+0A02pDC
o5hHWByq/SxWaA87G382HGwJ/y2w90gc+kh8EangAlkkynP+GcRABh/awJI3c84lrLIeqFZkLMeB
1AyEjiB367GwgX8zpS7zvkc+UG9nSlgQBeb558+QnsasNv9qrL9yH1PpF/uL3vPFvrTLBVKEMF2F
EjdgIRXw4ojTdDYWQErRVlrbRqZXFbGkXbtaLAg0mYUncn0H0mrieZPy3z7/4pB+NkdXSrqq69Wq
jD5xn9m6R7A5IdX7J/RrZYXV/elcvaxBQM6Z2836B63hcW4GpPYZytfU52G45jko8/hi/zL/e0G5
P46Z3k3sVy7W1gIZ+FCUlL2CdFfgiKN4mKOc/vkRFYmWSxjgegqMn6mAjBuOVz8gCqptSVtq0I9P
tB7Fq7/qwv2u5qHSnSdU4sbx5ptYbmWcpSVnrQAahy4ZGvhwIiPZiDPTd4+fDBQuCt3tz89wX33n
FXB25nlCGkG54Lf5y2IG3A3VLVfIOVycR3TXJOBXIEcWsusPopzl5t6nXu17IfqtMltnD4dBYiv/
U9s608+NUXg2J94d3M4lPX73ANL235Fp5h7nnW9ZaHsQD2k85+C1rbH5QclqFZavDHFXhRjOFAgq
HC+NN2BfVyPOtnJucwdly0VytMZAyfIBOHxfLZMaPnpLg7/NksD33OVuLiAryU6xdwlDTXpb367A
fvwyRZxmJpI3enwH298+yB+4+hRMlyxqTcGPNzB1UpgYWL5U/u7jVubz7kHp9q/7ntgjoUOg60jT
kksLSICAV/tbwX2tlr0FiTbvLd5km128YfjCWnbwTeNl+REBOQYI495a2WyiwpESoB8FuPrTKwj+
YDICGUCN6LjCidd1wx/xCmYPUbMSlmQFQijkCcVyAg2qWpJX4XHhskgoaZquekTcCvPmpHG9x/ZU
Fwm1yxmg2nlPqMTQztF+prDw4mXql+09i/KJxCzrkTaOPO/96bQx9DsSRHA5uzBepEDOvu+10hMh
Y0cWIAaBYVcOicdEtMRq2y/iNYQc2nHhQ6XnBiasb59xnfhJ2lYk41VKud6wYTjKxvDhAUJXaCn+
StOw65Rspsj4EtaqQfR1OGpIceK/NiuykxCY2k8NEpjaitCoyfbLakaA8EuFVIWSVDLBvfFrpFy0
nlXli0fbk9YMgUK42UEwUFbMfDIF//MdJrTm/r36Xlk27WQ2oEGnBhZSyGFNDJmZBnUBZ37c0/2D
KG12adIi0+jSEiLoxGFSFPp+y38PEu1KmcTE8qVri+dfIOwePqbyF8M9CLdwBXdpq0/3X2Qh0VSt
z8R8FtxCYxb8eRvPKpKnOd3b15TpBSRj++ZMYb0PGvaJvWrphqEZmbPVYbF0AWV9NApQnfn/orJ2
QtAiZC82/BTDZT36RM/f37/Vj8h3oFFCgIQWvyl271OeNewzLJl5fe9MMYHHB8WvTx1uriu+SWjy
06a8vVHkMqa9KhjryLSiVNo+Fwp3iD5c0khN++z1chj9PheZ42sNbtsqlFE+A+SEGrS6OLVPEQUA
WivUqMxs+DAmErucPOG79VvkdqY48L0qGtM0TBEa4L+3bMRSs9iWx+Oy42Syt1HSrbhMKUn8E8QB
OToGYnok8ZMvi3I2SjE4TAX0T00hQcrfSuExPjnepx9p/JD+RHOOvnInGQFxvfSGfcVfAEbDU3PS
hUYpFihoGf4IvKTwCxmqHa7u94pC6xe/k0GGwjJBqKAg0bavO3BYq1xe9SxzU26A/R53p78bQidD
UkgcghglVWlf6MjqDQ/iLJhHnwtYjdnzF1NcagahHZE5AU1bwxGF4OeQ2tvMhp36xNSjMp7qyRA6
pNqNCpHK5c0hTntjVQBZJRi1AhZxcsq0FvucydzV+o9/VccLoyIiZkuYmTsnw8Q/wlHPbZeednHS
9znbM43upgEhC1zsJq34K2fvsI4eEYRe0unxsj2gysERo0dCvqhtF54MkY61f6V97skcBzG1JW9r
iQ7PEY0TYOPiGUYIS2Q9UogyALAoB3OO+CDEfF2hrVo3dlVUlZLyPSYzXpcnC8omcjFJC3aWY4uT
qG8TeQagknk0AVe9/hvrR9z8OBROO1FcT5KkCTSBkpmDws7N+fWndrYiS/9b5wOoYsHVTVmEupmb
tMqpVwCRze+aGKOtBBfdC/OBWai3qtBivBa1uoKfzLJp/M+YNoDDqthNjZVhuZpjSTqOLt6/gKhm
ve1CagGfRAHO/Mf1WrUGpz1jHAF/To3+3Mzfn3eQa2GODbiwxpk5MpJRVeSv1tb+lE1nrxidwWsc
yzYGXf8OLqr2jgJgnwQbmldF4lZsz3rw/idvISmCAxoBXuzGL4kCnPaAn1HP1dJKQ1Dth3yB3m1v
KWalhBhXhsHQuncyJVQ2F4pilamda/Q6eZ2DOhC9KBgYP5trxBLZRW9HlGnZSvQDeMMABIQl8YMv
1j1NrJtp8qmc5Jiz6CgcfupFHzQM/jJFirGDN1s4EI6zhAkJdFz+DH9TRadEuVgoF9eMX0st7ylP
wQ58wYJ867yjeTr23EJBmprDD55chHUqopCZyBH14UK7fSHN3DtGAbyvTRq1RYGcWRMfwl+n9Cyv
w8Pmkx5tHKZWksoIDZBbBTZUq3483wR3iyn2Fwae0Hw0najoaxz/klyzvqFlY464qctskd22EQcW
EjpfEYgNwulXxiRgt1ePNfFsPYuNlCJYwgHmk9kzDf4sedcmaKB6zLlg0LYAzVx8qEkxGY5h+nTs
O0KO9RFHbZ2Eim1qAs+CWl365rJcEij+mUAytWgsPstn/ogon50ZshjblWMm5VFZli/5+KakKzr1
qNNNuUtt3/OLbTtTiNAlv6vxFZtGDSgIxTSlHUGilMwABPq+rsD5s+2FVaOdnduXEBzBBktwnpPJ
rOPceHc4sHO8RvQ/6NzEeoBpF630O7RCyFI3tVySalJwl33AB6eTlC+LHQrZMeWsG0qYcTod/dIv
nTTzg3ZE48eXG8r0EvYPq33HVGIVgc664Q+f8pVMYXii+/w6/ireiZ5i3VMZA7x/jVQAu7iMb0Z6
TRBNDRPfsVG2wJh5KPinWVgEs4tMAf8rLber5wlvcW6pevvt2cAQV+2+gTQ3BzVwdxL0nqazAfio
hgWuymfTUT+7ZJyii8vvl1s9Iyv78acpcz5O2xPWoiwTfvkJdO+x7jA/zmgDrpl4iKMRgJnnetnT
D02PhzEkgIp09XRUUSAAHYy028QsfLR0ShyWbKVMOolYKCwiDTpwmoExz32BPwy0/Bm8TbUtv3Ck
mEPeNTFMJ1ghRAQfoy4wB0wJOX3ItADmL0j6RTRvr4Bvkj6UcHlpPIBxCkI6hsT26V1PwIJ5lK2N
JfO6DTAXLpigt8ZDd8Ak0Tmx3Wx7RVHAdMWrYcM4kcThQEQfLv/lTb3uFfTN+RiD6uSHNovSVPmG
ZG/hQPZIZYrt3jwt58AqYf73M0siRr3uchuMIK2wYsh4rLwV4IateCniPpnwCLm1dWVDwDfrmzN8
maPsVsC8JVWp+d9cWyGMnQFMxArW92UW4VYO5mcGeq01Ky8mSb7yGCDk+LABPMRXSpGq9aS6l1D5
YDOTwKY3jeVadwzSn/fF88orXY38lrKGETK8hmypzEKp8LT19cac93JKcRIPfAlDW4mx6cjHg41P
pgF/NWqfrWSoES2zRskBYDR+PMONC6R6EJ2plTq4wYnXHOqfLIu+s0YpJ6B5XT3dxr8kb4eRmp5J
Lc2cV/aDyvLrfDlKhCv3fa0DV2e9q7T7BT5MH2N186q9k16JcsdEFmMkMPaCHf/sHahCRvNTiT2z
5zYcMiQjT/KfNx5aL1yCRYIe+k6UHgKwEO8DWrCnOjlgTmivUM83EicQXQzUsd29YtEFVFBYB9/3
Iv6K0Cow1lu9BW2jARaiI6WR1jIckZUX4f5XFLD3/N0Ey+QaeBJgRyfKX2LGsnilGSXnZ08aVLBD
C7GCWv/0pAKG73EFmVyuVIQH5WUIy1RRJYRH/tA3HqB8YsPeLjb8GjInTic4fmfhry8/37aHxqXT
4W5wAhdLXZ6n41veVu9j4ZU6NwqgvgikHEVn17eLFsFD9wpQ//2xTKB1LH4gKSmGPKbaqCYsv1mW
NmRb6Lm3smg1z5WLNfyzwa/e5XgoucAYRlr+v8mLmCs/ww3gLfmS8IqV+D6mSf73BehsjllWoBon
bqgOkVcrLZyFAnB5GzSc0xqt++sV6IDzLd13HI6z4mKBa81jIesLCK6P4gsjgGidghjsdmmrsVMB
ikXAUKc2nnTWOmercaJBIQj7pwgSyxlw3tp8V5xKg50XZtdDQcC48sYQhkLpc2ZIbE3GzOCZED+Y
RKUfHhzW1W6ZU1EE9jbEqAyxCSzZkZdJlpX5MgkySsPtOFlTcZDUmpzSrVp9ehJ5zN1k9ds0HQHL
TC51vL20Qq8k/+HH20vtwj3pM9UInq805/azcXSzOHw2GQQVYujZ6WqdiZh6pOBJrFA/0aRQtXGB
Xo5/ZCnpt9fCh+rcFK0QqYqpiiPzZxXRvrhEp0uawxaxXTTTA3+axF3Sq1hIvzpClBBUpjpxqlL4
bq73RO3nSkm9AksNyYZPpPDEeK2S3GrMKOfS461zHVNQLwFExiI6kRYHZFQjEFDq8fkteI0PJqqM
39L2ibbIby0V4Yle/scpDM1BIWIfAevC4B4pLOE/I5Vrnu/juCpMdr3AZEC+177Iu7+BXJg74s1Q
Q1m2iVr0tbr+UQhEOjCWammWuSIcYtDrfOhG8olhFehqVCFnGyniX7N6zm/s/OI3ryeX3amczvIT
HfTRL6rQWOdqLtf8wATTTIcRrOQAmwoKMi/pmOmItXiGlQbc4Xl+blF+ptKK+ck/4t9g7lz6oWa1
5m9ojDSEO7N2TZXgune8/OJNtTwv631yYc0Q1lwWXl+wyy/Hd1JjdDe+oZFthbO6gN8l79XiM5kt
0uM/rUGaVxaq8nADjDSoE8Q5DdxOgz/P/lNOdWW2d4aM3ZlBVABei9oRKdWDZAkKxkFfrJzK4Gbl
zRwvV8JqXn37HOij1ZLYXLys33NIpDwaIANCUd2rmGbLj1iXgXBhE8OmW6oHhQk9YTDYTvEDn50H
AJ7wRoVGe83h2/bst2bMQsofHU+tHfWtIORRIsvgeddMW+MkIc1o+J5K3/xHnKlCf1ilHC6Z7UT6
KrUde4TnsIabvgLzxTE3U+s/GGjCsIrumgsbj845mEHNm6F3dt2zQVrEiVyRcUSDxmJtLgHN1kjx
SPCHcbPurh+g70M8/SunsijsKRx2b1TIpRG33fX/MWxKckOC3GxmMQn9suROnkPNMuYjVTVjtHLE
V6XIdN593HJlAtbZ5MqHq1ngvx4sudxA2zPZN4uDs2LScGlV0wQW/TW36tMlvYaBlaFTVtYdO1a2
MchldiaAILks2ya1AhPk4HSLwmsiSmFyzIozJMHCNsQiitGIu0m80xGo6We0KDIZQYDZrJsdGrZ6
qMzlp/f9wr+5247dwjfufEMS3l0I2sWZJnNpyIEWxk+Lrlw2wluBIBzlGHshuZeUpfNYpWCpPz2A
HdSXSZP2OGiAmrkEc2hKZhBOEDvX1h3I/5HKG1AZrJEatd+DMnpPzJDa8vw5vmjeQqu6wFo+sv6R
os8gpzTW9sddxrqNjms/qPudQ+u+nbxrMaifvCU+RZUqCW28GTbbV8d3VMPG3VBojSO0L2W8qIg5
5F6WjXutND/hjV0w4EnbMoUyqL/y601M7dX9woVf8iZj7PJ/CmRi4juX/XY6QFiNJkW2imG4MSMn
OQhjN4XKZE8xz1iqzyUv7UAztCkoea8x+xb+FKAt3mSk1nSCwrP/gZKmeSRUgqmySlHo6wTm5czN
WqTpdyMrMqhKjRA59QYGdI5dkTi8gGtEngCk8UShxX4WNf8w4q2r0u8NcpV8ZVeMDOTiy7U7aufa
Pzk7xkbTm/XJeIzs7ErFSHdC2d1C6c7bB7sucdhOxkLvjdQMVFQ3tneFjsLqNybU4ui4HDgclIuZ
H1OdM8wfuG3rwYGRxcsCjiDkrVlw4SYGpK3WGXwzq890pMUNp1clRQMXBVeHv2AewsQ5xKwopctJ
LMhUkQL0y92KtDR3JY0TDdzbIKauM7wFiozfm7Jf2MTE6Ue1zLQxsuCA6Grm1Jfu7YP8zzZBEhHv
0iIlEZ1q0/7a9TyJGvE4qdaAc5SFbsVnCdX8Jhj7yROVqZqoKitkYE+nae46HTLp5+8F94sMiWUZ
a1/cxbnF+0wkgj1J2KQ3QoL9FW9S5uo1xOzrsHwMjz3WkzRcrM5IBI/E/IZ/8f6fXtl68H7O3eaU
XXMaZ5gYdbUNbfrSNA0S6GMM3APyDYzlHbpkyxZfsdSr8xDVJy0ZUkqe1c48JMlwpTtZYIOhDiv/
NBCXp7mqAzoGlWKZqkMbIxMekz/68LdhrCrmEm1E8I0Xz1zIZujV/sT/AWIKF8s12a+YkKpljFFK
zcFxDAhOrLnFN5JwvUbaYNHw+m6N7lyPRT9LsbWT9ghLFeDhQHAlWOuREIjGHrk//dtCP7jXza1s
7RmCAs5CmtKRud3G66q/CfFr2lU2poP8N3lPmBSHCDuXCfanmVF2gxBPrxkFSoumn0eAiRL99wj6
/PiRsBWiU8bfXLZ4hNp6TZJUPi8Fv2tz2gXbaKL/5ITZdHqzldEj0EU2Z+XBdntmbj50Mx+6lb8+
R2yci53pwWi2wfdl2e/hkgU75szVqpXQKb/Bw61ngATep8PQt+iK09/xnzdyP3J5B6j6OnkIpMY+
6KsY2jfYU9juVv+tIM92MvlORsayzC2+lqjWEczVKYYIN1JlIlzo6+GW3s8AtPCrQZYQL3D9hj1j
BZcQiR0erLcOQvoL9Ul9dlqGf7ypxKSjZS5Js64LbVsYhIyb1Vdkl/Dw11hVr6zoSZN5HvsU/h2c
kf4Oof0B77edq5zKKbWYmZJfRH+P/emzM0cCD4wzRjUDtKLv5Wyx+lGGjmRodxKn4lEqKkadGxWH
Mvowif+dyL58UTKXaBF92eSX0ANPkd8DAj2i2ksm8QdKLnKDnAFPE2VrPShkPMoynXCnp7YiYqSf
z3BI4fFU0IQZ+6FHHif4PtXiygLxZIrLFgcoDqOicqP2zsGoF2o8shFUkQ5SjGyzCygocpXxDG63
TVvrv6ZOjdLLjFqA6QkXH72rgsO5PDBvwlyJZsgcMzwo7s6FoC/l8aRfIrzNVEWX8vH0EX1cbJiu
F/ABpyy53GWYLPN8e2gP1mpVsjz4WBBCUz8ugrCcztNH69FxTeux9slFgV9eHkiR/5mfXoRXQgfw
vWpeEl2zMx6WSXVI2qMNHW5Gxrlga5GASNFO/bwapppC3nqP+CjcRpa+0Hm/xno7dGtwhwQU4cGT
WtfoQVFEjth+wV/ZruE108Zz21gR4jGZPt2+PKO1EnbumeFU5rVm6+iansHxJDyxYMFq7PGU301S
G34glMlQphtMEUWQkJiU1x0BiI9mw/mNepgrafNDsqxvSHT1CNe9SQFJ+Y2E86qVJXQrG+1qYrhU
FpJfPbB9p1ZOUyVOw9r3RPzWWmNgOqJQ4yZnjRHf6WL2QS2NWTmvqhj08VWhQCCVgnpzDlFv8d25
LSmkyvc8m7sSZcoXmpBa7PO6ZQpAh9C/w/R621hVZ4unX//jt+MzOt7c8iFh47SQEOf1nzNPQAXy
wQXJp3l0MypyUREMupMEs2FB6iGaY3MrzFiIiA3O2YfWMTRJ17waSx+d+nqaQ8Bh6yUioUa3EiWY
AaQdKPgsOcGbbWY4facf3bJeqKWlPA2VTl6kYNQiMkMPbpt6dSzq/buH1dZ5JZLe/6cZshbxob+P
K4bOsy41xirTM/GhEhlAxewIjUG5m8O3FKmYOuwjtLYbmerTXZKZg89QB3ILAnCGo7KtTPX2LaJa
T56xhFAZYmdj9IEEw6XnF7X5FwW9P7n9Kmuf3RmT6chwnHYbDGkUHz+Ti881o+uUgvueYaegCmqH
KGTxEndJzYJCvb+AjbSxZXZXk+BujAMuCkjfh19cGkVBJGTAf8S77lfz4sEd2p27qbuxBAvALbmh
aInBYqolBcVegVNx7muSI/WMWI9+C5hjAykas6FALYGsRokQCmaIuj3E0wpsTu2cUbJycK6UYfjB
H/NasioqsSqJlp67q/hiq6qb4x/2ZPAY/rZaXQxtKrXyk2MvzHuGWMfigU48/BXnRWSZw2+Nw+IA
DNRarYPeCEuOTr2+Xzs1PWwi4dWgYble09YSgcK4Mny/vTSV2MqZ998DtY7VnsCbcBTvL11sBwWT
reCe+AKWSLt2szf5hpkHIWkx9yhsYqnb09bnstLTYgWUtfLaD7KRrAP+VK7jFrfdYidifv7aOtlf
AobaVj3345VuS7OxukI7w+aO92TCh59QDzWCKkUapkqJTDshOJKFJwjLdJmBPDkc9hnG/87L1Zxq
xXToJRNKg2vtG0ZyzqcFQJQWGuefxZsN6HF6rFvfw5sn1DYsenqKehF4uaA4wud9jzYIjgmcOGX7
Sf8cl+C+V9igZBBDm95af+kdBsNQxYoWAUGkXS9k4BlK6JeaEUvqwxC2kj4jEpw/3hRN9g9jHsr+
v1MF8ChYNfKd+mWVVTkSe+rbkMxz0zyiTtamxq5ryKoxiqm1Os1YtK10tzjTfYQus7d2iWkOrwA/
es0vMGoGBLY/dFdfrhebeySOnfIY4h25sdWD/2ZYJoZiR9DUWuf0S+o4bzafwAsMZ66wKnswABqD
MXxMcwSJ1vBwHAmHYyXQiEbcICpDpzq1det7gWTw/e86OEJ/b6hDkfuiON2zXdCoyXY6gURX4mSM
jb4orPIk2OV3Qz/d/Mgd6FcALatmPLvnRW77JBTPNTyJJtoGmo/os0a5AEWQ642RBhGufi+y3p7Z
TXx02cQ91KD6CTK4EAo4La/BRtcSrIlpl3hC/eBpCDwSFN9sNN3AL+eQIwQAuJoBTdnLVd8phfSX
PATIX71evjT73VsrqBSIJk5fYlL28va4c3o0q6P76/cBz5Z9RKypg7IfPOEcJ4QrYhari8uUtekN
pvjwTHSY/c2wmzHk5Bv1xnTMlb/bIfDuKQNAtQVhCwF9yUIfKAx7Od7YbmyxvPqxmbx9lyVDW3eu
F+xsNLHDPIJE5q6hye4BThhvcsCBltd3oDR1OPO034JnCCMzE19jHoYVtC9KfW0WKgXb7sN+yrTT
Ffm39PbQrb8KQ8U6p5vNupsiQmTGW8zHr+G73bZ5AKfOLNaPR0Ham9AszKQlZryFXK4rq1q0P8cd
mdYquazSm9n74lWVA0SffX7uC+1BgdyFyE/yBfLHLIrTF8FbsfmjLmcGKXCNWeU/LDN85Whtylk6
N/kQ6mSwNxcYlX8p5kIPind7I/lyZf0+mpqQmtnHPnpR63CdV3aUYPBUtQHVHAXCIj+xNIdqmYDO
lA5cn180jILK8BH8wjZTe69LdGkA76R5KOPxII6YiHO6tMa6SLH5KWzIe7PmOIaeNqDYXCwTM0MS
fMEDWX7djxtnA32vKlTVKFXqcUyl1I7/gskP5GeEga25gGDDzK4533bmqQc005YTnsDE+eD/fG4C
oqEboNL3pLg65MV0OL6CUlj0M14/zaAaiZGhRK+LRdrdCcVT5yDQ8GOivg5S/iKE6PLezwa0pmv0
DB1S4wfI0hhhJAvvXkw5WzB1br676Yif0i0CyxzQ3AccVtGlhe/TbsNm8T9s9VTU07COmHglsaeE
pBy1ScMiurmKadU6YIJnJ4ItO38vqhpVaIn8/qHWslHYxn9hCJ6Em8TYPw0jlCLuj3lYJuXC5GJH
G7IhMzRcmjd+OKGzIZ7e76VH8LyiscVqAdYI6a6frUPg2ZFWuXbk/nNOIzu2hqcf5rgVXxE6pyNG
pY0bghpCmF5mJx5E7cIxXxQgWrBie2am2F8gpt5QhjS6jt9Q+CaCta1lieJ/3vPa2olB1b0VPRJD
u5iIvx1f6/V1m+iJ1uKXs1vr4A9J9aiZaoNrYJ/Dtx4wzAEDFfIIqQihEt5xCHlzpSivms2r8CAN
00aKnIhljmIKwJwC686blaJLY3J5w1OopXTI0y+S5cELv070eGiHa70FzG9Ylb1cfinrLwuDnAAh
CdLlWtKcF/pOZZfWRo3u2P6pjPLg0F2L6O/jlGf+/SOBOeI0hIp4GEm2sST0yf3Xd0v3FaiGmx2c
HOtbGM2sDebp2gwdmdz6gBYjU1J9bh901G4HKEWOFFDDzJ9qjuYiUx3v1hbNnALwUy7FrCD9JWxE
dsg+yWQYTvsR8rnTqC4L/2tixZ/Acu2VceWwHb55qskPCmhuEnYxxbaf/PcaJrSmfhjDeM+lvH3T
EYmEN1pHscwmT6eNR/y167HpiD5iNCnBaH8GGAimRqGJbAR7m0Dp5i961pnpRDm+rITtSuhj2628
1IqmzWNvJCCMaw9b6PheEKhDQEIEQkQmkls9NGfWIXhR+v1c5BRr/ItJIw51ky1XGtP604qdAvvu
qko/yMD/aVIL9b3CSJdOacvp6JkALpEbdRa3cKX88g/bJ+V0K4btAP1RcK/RbTLS8kK3X1I7f6uJ
9fh1MdYCmWFH1NqOBlCqnm6sd5JmQuAnb2j8c1N3odGPmFPOiHIcrjO6Ij//jUaO3iuE4Gm9nMwp
J4G+uH+JGEXJC/yIo4huOKYYXhrwnML0TvURv7CBzl9y1BjgeF1DwhlvUIIQaIMWr/0prn/q0wol
a2LjW33N7UnbL7KmcqXHKccTT+t+geUEGwE+WfPG8uq2i3DEpwNlTG922a9prxZIOsd6c+g4svqd
uoS8vnOFizjzvvx/ENdtQ0JqcNKY8IgQr+OzPKWz760UA/n25FtqJQYHPriMg5ge63gXEoHEAp1O
LbXmnyVt2XTnYu9W0lNRT9l2GGtH8bvzAfKCi6Q9DnyD/P2NIni0SfKQ/2PJm8YyfCfNcG65Xwd0
TgKiWLBBNsrG/1dAn2rc1GmORbjXN8VecUu1iLH2iEjNz3xR5Ti319zYvAOhLwTi2BiEz+lDt42S
6vPjDaKc4fphUXcpQfYjMZbnEFYwgwetvxKBYOF50Qumdv0S1Kd6FYsFr/e/f6eCCqB5ka8f8dPk
Vn3AJyjp8mYzLEov129j1dBNLm3FlcfEEULPCw6bKoewnZ18eHk0vm8ts7P28jVu+Y8KxRZajNM7
CRUQAjOm179wRQhvi+ByC4UTlrvWtW1pLFrDsV+BGudkbbWYIvGohbz5f74t45qA/cobt2h8Va84
tvo2TaUTru91KAi46AfCvM0JpBp0C2yKBjmsEbREuEuULdOAwjgPB0vCR154kvjdm5ADHAt9XL5t
WZm4pECxwtDmEgVAtiXRm/ImRM/mWnFH/UQyvO/IT/PqCwsmpmv2jn/Znktn59o62HFIO6ebjd3O
4m94uEjmYsZldWbyY6Eg/tdM816KqRpOSNp+EJxvebfLH+VtOJVPKDqFLPXFEYXm3kuM5BAqEShp
sO1dOluFMzOhWdF+shMK7mjwLMRZOJRY9QfpjG0adwaKTVJarjbF4zzLfxryPE8x79w8Odg8EgpM
FUiF38n4to9TcCjOUb4sKAYOWw6kwFk+JTjk5n1JxLti2HIQmptBrC1D/asVWh3tSSGO3i6WxAsT
f37FBF56t00imSRaq2WT56/C/9gkS8v66kcWC2sG+d0S/1bsp68RLtTPR3RIVp7EU3p/2ORL0ZWW
DbOiDhWesTf5eeISar0cPXxliZLFnd8ym/+3v3AK4nKVttNGMSkthvqhvjbbggKOUeevda1W91R5
soHjcQkwQBuHZ9221L224mT+8qi/KsmhtUUBu8RWx/8/1WEwYkHxtur0jHePZrRFHKXaw73Uxgd2
jOQAbf9niDYn7ku7NTARAH4ZYy1Fi4QhJtzFfBZKRTFufeJgRDtqVTt9aUZyoecjsW4Cy6CqF+Qm
L10HZrvbimjSMzQ4OTiQC6SIo68k49OO11I5SOdck6qraK62BYD8Xqdbj4fB2wuOEhm36HrGrlUe
Kcqhw43j3Gf2L6Xhxj0Q8MMgfW3KQmcjox/NR0YQM7F9G6nG1MxygmE+0PFNOAwVQNXJ8xgvHk3e
Px1Zd/UCHgiCXxCCPaD2j0ucFZ6SgylwPbvYv69E7Iu043rExaPuOfodk8/4kpbqPvxNG/LVv0MG
WEE6UNOoosKpENytj67r78bfdJ3ogefPAV0EcqyArztBelIOKx4xruYhgjQzO8BPLpO//XMXi8cj
XkBY5ilG/CY1j0aruARLjkjY07RqupBDiLiUtzwSuu1WuVMAbTV+X+JEwvRp1W2iRp2dTsygzB8L
34nh6KqcKpFQAPE9xZMvQNqp53/NgxToHT5UqbkqlUAaiuZdwn9H9WkOsuOSPopJn52Ly6KLEuow
PRlhvweBm6hI1Gpt0D6Ycsb1vXeCYvY25p3kYu/pSLLzcDCsVrIOW5mYcrYGAYaD+vfHzgC4anB3
xErcLEl5HlO83W7MisQT0GETS8RXbJQK8hMqeKqnj23oSuH+PwSkkpuSm1Ne3H3jrrMpz9Wq9g8z
O8iGyxSbpFQSL+qU5hVhQAgITSLSlp3eHZkkyg84wwTdQQqXmX21AzFVfy2L8OVdKjpF/lLSMsAQ
Q3OSyas0EvJ3Q2vqQAb6JwIK2GqUzo6rR2HO+V4hmLFcEubaPccRX4zS+njSUdcBtf6asEU8ER40
hGoBjaTVb2bHDEfMkB4zZBgQmNTA6yZ1KAcEbehB3CqVTF0gXU10U6ytJ+U5y8QbEovBcBx1RDdA
nDNLyRawpzhZzgpMgLFYgNkds+9GGeuEH7tVt+UDjfc0YSBxniSx6cgX16d7WPcZfvmy7xGiHykY
7heNEXMmJeCA4+zj40yjNmV4twqv5NtrHpUv/pHtH5d1XhNoEeuH193lBCg1WfdYnS1ntpsCftKl
Iq6qi1Q1nLmJ35t2BPwia9VujxwiXckalru7hnHM33lzObObbB2rtAqaq5HWgCJ2o8h4tJxXesWo
7yizpx18w5PWlP4SbchD1ev18CRfUwWmLZc4nkeWM0w0znEgZexdQXrhoNaFXJpHrKR3rcAXp2MT
1Cp4cdxC6WwJ7xq1A7ICUykjNmnBjpX1wOoS+d8Cods5keuRJvXbIEcqSflNsESB9FR29VWaYw3T
6Rumeh/TAaYYX3+wgUyirJLup+uK8iA8uBp44oHpx5bdVDVdIVs+/DyoNV0lrjsoLqDa4eVB69MN
9uVobXv1KP2wV59NBhAy4vbBYg07i2fQDEPJYPQOlYgoywfoEHdfF0Hpo6LKsLrIuKmbfeZQSzpa
2bUZWwyXZwl6hQQGu22iTBOPdWBVu37h8kW/YkaeGHvzxPmoUs9HH7a00DPGrtQer70bZWT2OoJ8
jngxF1sHNdEBTEHEWjmesRjqP5y9f3alTcO+mUOuvXMvgMTCM6/scvBHypAMGGzeGc80YYcm5WAH
WpZvKqvRCuXSMcXdmt66lY2PFMlOC5ZY6bEG9QN61cCOF2AUiADgsN5NdWiRLs1UNZ7pJNxtHzau
XSgYwsNfxQVqHEWdRE4Z+Z2N3hpY/Nw8QDp9fYbpxbMamHzdM9uXCiCmpcgcweJ4BZb5k077kq1n
jZeDFP95h+g9xUcCsFqYmZbSvmvqohypQOt+1RW3SoEAqcFhoie7+6XlstljaSsiGIL1vCnFFRrk
htPc6ewAJpc7j9gVerGY+3EYnfdg/I5gk6snaM1/B3MO+mqena5V3G3LCP9RBclrBuiTAlxqbOOE
HBAJLx7rF4cK9CXrS80rKmGXuXr0KfObh2fQbUv6FtT6smhIq8QYGs565+DRUfmxqd78vBDMoPME
MZzdxsrQCZApLgg2jqyXaYxpb2Ktmh3fXhFguZYYIXYSvRQOvDRWXKkLlzbE0ojo4IFzb1AyBm0F
cY6fikHZNyr3o8howep394TZAyOkbrRFw43iSVKe7tix5yUliFmIJX9xuh8+pAiE29X1NXWXs3A5
bIdMNAJzicwf3u0tR4WhMDKe79JEMniAclkpmv0y0AkypwBym+DFFbbegd656v1gkUZ38ZK/Qhtq
MfvJrd6JyF/h36bwaAE/yFi/ltbySOPvC6foR8TbMCjikisp6KCDE5K7A/XEHZU8LzJ6aQMmHGjJ
R4yyvTgcZ+97CGeqddds6gStA35a18WEjrW3q9jqtBvs7/ujoAO98t9ZIchUu5NmjPTTpydnAoQR
Bdxg4xtpnXuPMuDduHPfMupQatuusHGQQ1ULa6AZUqwd+P2REQytRZp8oMrSntxfbfSAPyVZw0bx
W4eiozj18RsdXBASWkKaeMbmsqSstF9Jy7aU+/T+bbfNdc4E1iPgoQntxmWTK4DhznL3jOuyHfC0
NcJJOi2TOvjZaXHTZk7OxoicNuaPXGQyIUj5SQZQAAWWjanz3R3E0vxSaFcVUrsdz4yugsJ9t7ua
ltbhE4KnDZhF5MnKIJ/+PelySQbzcyqhe8za8JRFfa61cPVn3aIguCt0sOzAAeslWhk4+PoSIo/D
mKvZNkBJz7AQxisINYAvilX2gaw16uNw3tWxPaNWv1ZIzT5Ly+j524zrFRs88JycXWpiMyd6jvGR
XAwH3IZsYAc+MluiwcFAT0YCzD+MzIxq0+vMZez51rT9Nagcp+YIOAnNsfrtYVkNaY3tZlG+rXW0
l05dFRDPx1knEQTMe9wMIM23Rg2+fctxQYjuqrikmqRnf59erHnU6okOUCSaua3d7QHG87Q70WeY
ZJvsGw1p5d2tMga2KYSDJbnkcIxyU8VhRdC3Fp7ziLlRWho6gAddaGJDAEkC0NuhqRQND7JWcLMM
1s/VCE4nNrfLgslWiYTpKKKKQ0c794o6VKaDY+DJsBt5OBsuD7Ro/66fwRHvBIPaPjq/dulIZLhC
4Ay5kwz+nLzjfiTnuInfb3+whM2vpvsCCWasAGmvJxUa9ARNw9qKyrQ2UQr929i8A6j4Z0Gm0nLF
gEo6FiEqx0a2RFL5VgUVH1/+eSvHKGMPKC1tJbcGx/qPpTDc9/BOMv4vUCkDkqvZXyxFWh31PLCE
LVshRrdElpGXVcn39GJk6iFhmEfEtTyWlx6pTQAgjRm54ltc1eQyfA906NjtG3LZsfXYKdZKwuQm
Zo0/bQRr7yS+idS/FxKpD8CAT82T8hlJknv172QJkVCT6ZvCJYnBoBn/V4r58vRrl/lGg8+EmA0w
pQXoK5LMKKVPADZuMjb5LlUu8lFxwleFBvlWrq7oryYiGoxNGjp64LGjkNKs++aKs0bwBAAJR26K
awKcrx99CsXV7ciEsLKDGYrggzZccKKYJINGNwtE0bZsqN6JZL4k5nrGZL8yt9AhL8Y4iFHteJoJ
UmCtoB0R2Wxju0ZTqA9gNn7nVSDswjQ6Zy3QwYyMhwEhNNGBNTI1BnSb8YYevsdpFXwXbeJqk0Yy
43Do7bm7wy4w/RI9sV9MJzUft1ehVLObuJmEQ7SBG9XGrXqf6sZMBt00fpzWBs0dqF4wojOTeWJo
0qMHiJMO0RYSsGeM6V/sOQMswmOcfbX0b78NVhYW+KwImqPqIcCqSJc3nqSHFR0FZYh9iRktldW+
JthdQat2SWOExY3aLTm207FDYE0LrguClbiT2kIK/pabDNuYpsP/GY06ORo/goqfWt+uHlqCBIBG
VbK7zK2fVk9yA9uqzNt7rEo7iErHY+XUcRiaYpckRyGHybedyrV5sl1AVpHXypL/J32gabutiJ2x
QBUrN9rmuBNM4zk/DzspBlScnWRaaZ5D3lGcG6hGIDfZCGto2RuzmfzZKMqRIM5wxqAeP36zZgW0
u4YNKaLdmR8iyDzwQ98PIy7zk1WIkyr66FrZbxS0v9KnXg54U9yQIC9DnyRTGOQg22M0wKHwq/Hm
GnS8MxMWVP2KYa3tfrMzGkzIzm2n3P8Kn+s4tPPu5p+EMKj6rtx6eOybpA1tH9iV5WIv7EC02KZE
xL3cNHY97DXxMSZMEnE2cPq4ZPsEpLy9B1Sj+sxCl2vTgmctvZJp7YPj2uYMc19oJzy+GY5Rd3CC
/dDXCckOJ0Jm04OHZsIRROC4Bq48geFJ83nCEo44WPtQx6SOIXyh3kFDTcDT0LLFxZ9A6QiuERMh
eWrQPNo/FvYkbi6YXB0CjpI7F0JF4vSX3BdZSg8qV55XNOuL0sXRvfGKKXxsaDbqWWxPzzGdpNos
NK9tQLJ7T7o9BJuOKPZnIZHIJUrNCTN6rv3i+I4mhcsFf9O9qMgWMrCXc1PcBBD3/bb7Rt6uE3oj
bGUBbZYRm0dRVyneTjVwoxDLSaNWlBXA/kFbkKdcbFQRQTacCkuTdmr9scDW2MkKXieRCdwzIdZL
hbSygYTweylyohqvR+GKwNX6QW/gU3kle1NwiXsgStqQ22BqjAWLzANhNCCW5s9abZv3xaSu7m4s
4xTGHURaGwiqJ4ld+36P+6RaJKdvPYl+Tv6qvKftzrnCabG23uDN0GrT3qutTvrOECovW2SRjmxs
e21S4NXyMmfqHotpvbt5Pe+QgWb9+nkiRqcOVuyqz4hFUJS9HGzXML9BaFELG4iPYfufoYqgyf/6
ckZ2rXkcWCPWhz4DDorOwE2K6vrwnmhbDtnUw9xZm+39UqiSf2ROr8KyyvJcI74SEHQH5iP+EbA+
EjaUx2EFQV+eBm4PgB8QA+tQfsIP83bl5Xgt07fT2yIbeLd3N2s3SVe1VXipE2rqzpulSzCTesyw
ZR3JX/aYUw9y75nGPSCWdSicGDI/gmWsgKe2eD/6xmjrOfp0Uc9xlcfNreKofJozwhv+JzmvV3XK
2VjlQ3gLZRUSkvcpZExzRXcPcpx6t9iVMZfQnVIYzQdP6T22+KIya/xhFuaw0iuhvcSUvoyokQPW
tzBOqeIXZrE4xx5OE/RbtKVuif4atjIhL7SuE5GSwhQUFRs0j7nOxKgfFBkuX+1TFugcXcosoVop
Y0lzsH1EXrDZl7uKCQgZheubfyC+wf9ApB9ayLp6I4TXKhAP8MM1XgfTyxJLYR29TTjJrCsFYlt9
2w6gBy5R1Nji8mJ6QaLyaNlN3hfgXQvQ+bzUX5pYWeZZeJ2u9+BfIlUnRpOwZA541MpYtzrW/OHV
BZa4dMWtVDomEgO0KAesrV0xVtOkgP7Solk5OBaP+d6idXQlAlIk5hDztIMLhqEKt9gWId4zvFdH
yn73iRRm1P1n/ACwB9sWCMme/1kYg6muCKH/GLuXrjqkCFQ8d0QzZWb02Cu+KnwBkJE3IgR2Reaq
xxwcHGJKGDesMlykokNOXcisCpCbpQLadlQo/0lSAz2zo6vte9I4FXuQadp8joAdCgGtMVRk4026
rZW0Yyah9ieCODKQYalKme0pgLiHQxDxlJtFVlt9DarYUF9aK4NUu1kBEWuQWZ1du5ypnnPN3q78
37MX0ijhZqn/89emlb+h9WkadErdzyX3QWTFsCv3RbGEgpbqCejay125KuOgQn+LxwUAPjTROlhd
54yolh8mhZQrUesFHJ3dITEOKgvyQdjY+CoRPg6xKRdOC/EeoUkjNSnSfu4OvXVoHuJxhxYJmpbj
AZi2PjIpCDw2yCXebLK4UV2HGov+7RbTySsvsp5X+5mmCGwLEVMJw4Ga9kCbN/6KID7AwNDVZIOx
fRyWc9olqYDqyPK8yMQTq26sxpAA4K758jKZPT78aSUJRQjiBh93hHwX2qZMH1B0gqgVDplUxtI+
CtLj3Xgg6pp/UkW7k8tijLRR8NYOiNgPWMCDgm8SXsHX44IInUAMKnk82//fnPRos9C58/6oyl6u
RC8GxIqrU0dtc/E4kz0RJ1/OXAbkxqwO+iGkLUkZGODv5RAvHFlzt/ybsA7NnT0dwXsCqK87FmvV
IKyEvSPyLC5Fd6GmNSUAXWLCXQBA5PV0k/Z0BKbffwxkHQhUgZQA8FqzPEkZ9qBBfW3Cy3N/2H1v
96eq7J+94qoS29JMr6kZLE3oHOtQhrKSuGWrO1enXh8+kmSB2zbm3w2j/zd1k3XniEtT2PXnH2EJ
00fSU4EZMpkGceJYh0AjvkYFGF85Vs70w9seQsSl0i3XkBDGVo+E0spVvkTgHSf0KHnxkVSFHpAE
2SBA2srMZeJfIMPRaf1nszAYOKQZ3mXe0c2s1RGPoh8XwAq4HDDvQJDtsVP5KKXcC+TDGGufUUMH
VjaSp5XYdo3XNITbrC7Fd/dI11bjqJNsx7NVa2LsUz5XdShcgLIDC8s15gbqCEu626+/CP+HZm1q
ASxa6kAfS66Wy0ZyieYgcbTMHxc0vIFex9khL1XripOZor2K9GCQuuKNCxAKSUciFMfDf9XW3Rkv
Etx3XOeJ9GjQ3dfMlY6Jkah5I1f3uatBopF8M9MhyHJqk6c/QmYfgHsaA/kF8UUsFUXFivqXvvAw
vIfugnwhtp5i2PS2cufuzbseK/xfERH3cFUccS7dmcbxNu/jKEH42zXqxfXyl8fXxahgDt5iUrHM
3PLApGkVPMB+2ByxQg/zmOt3oBNzhXsh4l/7+7TmXWE0hMbqK8cyOEPep0oUPvXhSkJjA785vOk/
W5b7DEJekEP8IiIyRRwDtMM119C3BEuMRDFTtFusYsouYDfY2MePs9+g2cqAKLRkaCUck/tvGx3g
hPlJqLgWC3/dKafMCQn/3+/TnsR5k+z1T5u9CXcadlfFy+5N2gr6Q3SE0dV1F34cCI8Bv2WlxEb7
VEeNiPMFk4d2ZJfKw1Bfs6veWiWazMv9YRk7Bf0pjkbonOE8vPswdNQhn1lp0AeWqHRWdo8skYkZ
/H2iSyRaLa6QVzR5kNuBvsjbZEesaoLzJ1QyXvGOPjhzeFcD9QiChOUdnOScdLURNi40cbdPvcr/
dcuT2da1d218/TksOHq4gkgOYOCFA7/j69nc9Hr6zJKUAKB9dQ+aZ7W0bJKMIYPX5q5jd9Eg4D6D
F9BNj2qoed3WnjsgM1YA4VaLD72SlAjlYUTUk9JmXl2T90Rib74KJrExUxrpPnak8s2NlQ5y90R2
xBaDXBUMv5Pcsm+rS+ULvFSgodyXfBaKecorxVX9LYgyuhOvEIBA2baQeuKNodoiONZvh/4fjKoO
dunMclnYsg410rWnUYhHCyPOaWtEVsrOeaO/w+x7TI/lx4ytVXNkbbuxK9a3D/Y6jnLVhtHiz9iE
Y/gRMg6YyShR7S+PilM+sNDJGLFAPWJfrroOALSPV9c/blW4Riiq/becxkpw7sIwYVBlGCNh43c2
B/unz5fSuK1Xnd8cDh6cb2X9VwO4ie3qpThkSk4DPE8SqVhCcd1QBmgSz1twXOCd+fRJUviiMWwd
sp0bvbiihtjAtyzZn++B39G8gVwc3AbRNI3SblZWnK+32+cKiVdbbYGMmdUwKVM3xl+ocCVzjUmY
wC8M38yohHw9POlZXSvSzXKeJEWvYyoimiYeH+5v9sO/EVTNspLWd4rH6JnWqioR6r4gn+9/6EgO
vCbu+bgkC8Ec67DREJhr/Dds5AtDyJXTtMsIApudUYaK6zdn90Gt7a8azqIEt048fH1i5wHyn62i
HL0H5jTk3Ras8RPh/MEsrJ30n9HzDKIw95HaASMqQtz15abTCybicSDADa/4oi1w4Ug1oUa4fPl/
WOF5QcGezaoZaFsO4YdlnAxVqMvxOFdJaVDq8THUjYtE3CMqZcfCQZq8UbOnEgjj1aiGeGzkRWKR
pOR9F3JkJCfplBcZQ5xeRq/RJZ6It0gT7vwk1yX+CfdmYfgurq6+NoALzQ9o6dj7/8tEbKjfeRRE
2jnqO1v1JDnizDnJondckuE2+LWiTdeoD8GGj8x0iiATs/YueZfbj5eF25M4Ig+TZrdNS/YdTu41
pM0d2ocn3THnnKfMKkzrednAUSysZ0Ov9x7stlDEghrbC81Eidjw+XpUd3kmIA8CYnXABlef1vej
HK994c/szFIfob3VKQF9yF612Bhfz7m60CCLQBkJEqjyMiO86q8fSUEVi5MNQMOGLYAD84/bOKMl
cqi6uTvFEglcsY4Gi5KtleCcDqyKDYyD7FA+BTpe+jhG9N2TVZBcb5pVYXlJodfx/JcHer1THqQy
Kikat49P/e3mdPA6duZTfBmxA2tXvgPszhthzlENn8hBc+ZZ2FFqEZ/c5nIysCSc2NfH5I3OUaAV
MGubQ+WS5O1EWnEUmG+Fm8QSmOhwunpsZ/I3jAFiqzY4qNk2NDzsH1iVjLpg2dD2dC1uCHTrMFTE
AjFEo330qelpRzW2U14gATqD3CKnfjjNQLq/r/26uY1YqbdtNcMK0TDRPM/Iua06cWxb6mAK6DSn
phGZWGaRQyxfL7ZsxPp6+7ATa0SDBKYh1EUJfCuVLqMY09NF6cPbc3WoqdVOowVHWCG4YxsDtxqa
8TBiV5oxsvN/xeFXEGn+/YuypOrvIn+yf5PmsJf+Twt/wFJpwko91MgpEvNc3UKFvgIJsTfZQGc3
TOBn5T4a0AuxzLZotkQJSoKanxIurUceWFvb3udaIP2tPf5uvMimzJwXOaa9Fhz9OfLBuD7acMH1
+RZXTEm8VFDOPMluL6bW1XL4G9zU1w4XyhphPlK6agU5859Mm6mltjnHJ01Ja5hKHMYFxlFCsgyA
5oOgWb5o6q6epeg2f7qzjM0DKX3PKq1WJx3ir5hDOAhLq6YsqzUrG+OHKVEMzC0qZIk9EmwHfyD0
pjiOvjeGoW66TzxJqdNwG4+b1LtyskqeTFtDxhUBZ+MQKPWWfKvL0CFMpZUC2mbM6uOV+edAAY1c
PMBBkvDIEKTcEwzE11Nt94r4Gq+UPx5YI1dQhMj353fJSmN/o344sabxfEhK2omX+GAQ4OgCkPku
94YtMOhO777VwOU0fnOsIyKIuVtaJhmEnDS/mndoWJIcOMioOoonWhmysvciiBDUQQ2y80rODWvp
+T1skB7wbWeI1K3pMHT1mnZdfvZQ8XwhOFMtmvLzvgzrJZrK+Ik92IO+AQYd6qqzphRLpZDrUBP8
x19VO2mtatJYZZ67j0VDf2F4QkHPWgXrBofirQDEVLg3N8J45OIt23AUit4+6F18FfGYUtqhgWtG
6ucNVyonKtaoBKQcf5HnxxqeWBeUf3H2x5gNcNtN3O/hfRS6fKDVqhge02sg7QjMYh6lK4QjGQAv
O4w5V82Wb8SSPAnunYTnTY8cJmF8j2OzKsGjNZBy4SCLiYIOCMcAo7FO3O8qnulIiLjdnKSr7zvJ
V+R9QG/AGnzGvR68fYQPnot00XlO8KgZUbCGXCIScIpj9qh9KWiVzi2i+yZBppzEgy0hXfef9Qsr
q6ASTBim6KC7DFkd/XlIxP2poOtKw4S512Ga08xlIh3DfigGO0bV9Om/VvRUC+GilGHfgORp0dST
s2cK62A8WNr+/k8Dn8wdz69bggqqJtr6+yi+EMBUi9dfOvjYhh4maKZ5xwPY5QVA954Ib6G3/P+P
l6OD+rOeYRPm3ZgLe2Fn3TZnYOD1BERfJerqus2m1NcS51bninnuSOEd1O5Dy8T2GOp/2IirpN97
X1hGqN8XldQhbASEQseqRwkyusRrAMycxL6uf6x5kPpIcDDuQ/Yoe3CQNva28yAYhte0/7wSDsYt
81n4nF5fD7ppz/or3X1OAP8nQ1uEi+ybWv0NYT2gbzXR3JC+I8SBsATFut6HR3X78acURhGiIVRh
XJRtcW2bo5lPwbsffI/rhE1TPRj7bmO4pOg3An3srjRWDgSR0DdolUuKlSdNDg7Yubx3QrF9zSa1
7n7jvyuv0w2+3pfJRnwXzGXsja3FEOkBgHHZxBH+jbcq8yHmaoZVLMwv5ekQtQbSX33az2ubwG5+
RhpgnX66s+Phnn8A0OSXg+WaG1AIv5ExKA7C5XqHWJDj5mPs3catwNLxCnqusB+5uEd50HQEgfcZ
C5ybbI35BzLxr/kkTLFa2l/r0F+xi8FLDle+dAFlKF6Pq0dB9dY5n0bvWmVJLv+MX66S2DCpD4PG
AFvGY76yZQFqbkNhLuE8tgGs3IlkLXr8AbneNDCHNmVvhAGL5PlIav37RQWx9nyX/kforlsH81n7
HDuxbG/rQPzchBeJtDc+zMzEgCi+GQjKgqiQkociLlrSTBtgwoDJ8i36ye4koZOcbbDuVaVXhfYr
8s0RhoJgZgdFb/kFLC8mBIrYEzYmoHjh0EmqFwUWf8mxD2yoFwA1tJl2KzNM+c5o3nHgl8cfU9an
jfPRvegfVJBaZtKjJxUecjanZVHXQW7l1v1RYZBnOFDJ9xX+9jbSRizzcbZzKGaB8QoYAFdEinQh
eXhIzO+sQRwfyx6AINfZXqu0uzUXuC3p9QKH+QDE1023Z7nrT6ho8LM7rK/sy2JjLoWyZckFcvGS
vqk9ybTM9DgnoQ54/K5o3L8AmGen7H0YZygHw4hllmKF82lbPBpydWEe5WBLgcQ+f78Vrx8H+axN
W1bS4PHFtDKvwHwZmM3hCKnneiWSMp7Sqi3EuRIVoE80kyOQwg/v5Vc1soC7pj+e1qDdQ9qvsYH+
7bwTx0iwjyVK0jwL9HAG7Y3Wr6v2taaIA1K2PrOjMYCOFLsxGzc1n46BPv5e9cnAHzuHopS6/VPI
jD7oHIAAPqyi2vjUcc9cRaWZvafBKXtgj0p/dj1qii/PK93zfi3rB8el7K/nRb5/Yda75RoearaC
vpRgCmBOey0m6O7ZPLZAV6Ut6j/vAnq4p+b+iG+0zU6JbeI7+KdZJowrILKv+WhcgmMkBkX9ku45
oNz+Ho/9Kros4PzQm15VWNlK2HvTdLRh7bccioFWaH8dk+68fCPz3xQGGxjHWj8X5N0RKaAtC3UD
7QrxlzKWqt/05VAeeLaKSp9jbjT2zPPWeuq2kg+B5Ee+4yoeQ+NWmGkU5h8+9Q58gPqI/+L1fu/I
hinajBJu09PvNeofABThyNt8tScte/G1G42upcRzgRuovX3fXXl4QhcXwTxrismwtfQ6sx+nIhzX
jtudG8KSo62YiGnxsn/v/69GGF801spghy0Umoi2a+o8eAu++rUHNy5RIAE+owBRVQRkA/mJ2WG5
GbJJQKrdKPOIxLMt/gxXQl2CDsD2jCZ9Owgarnayo7x8UtXdgFNrPLl4KFUKy+LUuzYQaaBYrvs4
0IjA59y8/84n05vkJLsl7NFvghlhDIyX+/U0DownnvkXDAlJ7iNLxGlA61DvvojnpuGuY8oozLVG
wAxtTrUa8ixJbEoMh/fpKlCqz8BY+z2QQTJBIDUWxp0m/uSl93+ehY2CC7MX8bcf90p7bP8NVkIG
B5+cYmrIwACscAx8daYnqt7yy0tD5B/iFIMOo1DppuFx7Db0TiG164ta+MzAbcAw+4AmVoloUjTE
Y9q7SlBrN00xuQcPaxvSFB30srb9tOA9ElBIvVQ/fZUco2W3CAQarrV33+U9JRnBmdGpBFtkbb2j
aDaomaxZ8+lyGkF0uwke5yKOzDmScFX/zRkyj4qk6kres0nAC5NKjuJv2kRWhcr1Yd3nrdf8VyMJ
7iStXuIqm5p02BFZdu6j94eH6AEB/5WXsYGS0HG+A0B69en32Kpe3v2NcdowdiJUbaX5UOOOO5fD
70AaYQbV3FI5cYJyRIOhUs8G1vdWyx4ffQdrXXlsDiB/7SCZvSW1oiqh7z/osw5emeLo7gHyXVsM
66AkGIorsgnls2GojcSG3+NLKSd9IijUHkzY+eOIqI5XH27ec2RV0SjZjVyoPyXob4pWM+64wuwE
6k5dn62srHRjw4pcbr/JrJMQmDKTBHYRHotj0gBqeuhOpNRvvqDfFzUMVUR0kV1p/OqcBp5yg87o
Ib25kYb0EuhQvj6GIjnb7IciBiD3qiXYxsDssmF1E5umDWh7p+9K6SlSTRLguVwBENVE0mYcgSj/
x5JyMc59kSsGMBSIQtOic/vL4Ak5nteNq9ZI/KtELzYSnYQfNFeXYPnBnjYT5MgqW4U4uuMhQUB9
r9M7+r8IaTMwwO0npMWT0e3G98r0RE7lYK58MtJTIgt9Q4dBg/ob50GTDtlWsl1vKUNVEaKVmuaX
QQTDwaq7XXuR0g8YzGdzmx0hmj/l7IAspqF/oSjNAYo5MyoAELo1jAqJdl4rhkfyQQZ+Izlb8yBp
b/O4XzVSbSx/8QV23GqeKDnpmSGPjekgIJXRrxPgU9f5JSzl66zKsOhj/AvMLMikHao1d2xl/aVS
m1xOe8cEMkoXfE3W9fBSVE0lOPwdeeQeacnIT7KOn7iUS2Xqs+mY+hbjSGgO3fWW3Fc/9HCpJPA9
MYBU/EYGkT9T0Mzo2S1TU47Eh/+Nzoe8vQoshrsU7IaszwsM+GJxmhleCnawtlGJVIOt7lLR3pP3
bbtu0QbyxfKjPs42XTgFca583dB77y9fXnS9CxCn4a4qWrf91ETBweJDekX4WTBLlY1LxVpKcvx/
YjDLgxfU6cHcSa+skmN6Qa9ibtl5Tv+kNwkhDM3HQSorFeEcoCwZnYvXk4LFqmnORpwOXyaQbFmL
vJq04b4lBTl84t60Jm3r52d9EGjU9jv+E7KTLFIIx6qRc8x/FcZOMswGKWIGDAArBWmIfyTnFuPh
TIbhFu9aws+r+SL6+28c2jQmY+vX5DbDzyFOy4ETamK9yiywRGprshI+bDA4Sr/l+1Jg+OGldN6I
lXh4p0iB8VU+wqySwwcFgKC3N37pmqMBZvdcU73YD5cphF8QkhAcUSOq+RbHNbOLwFMKhwS7onTv
gf0t1UcU7YjVntXSlCtwZLBDJ25PCZHvkclvWqFrVwSFlw7mZBAQIxDCAJeyulEsXABSBjj8aIgl
2fljtiEMOfdGTD2G0DtHe1zLBRHTUu0R3zZ0ZhT4fCC+yMUuueOfrefuDTBxlkFhXx45MdzW1gX4
dFUCqC/vm4t2tK+zwCj8U6FitVOS8Dog3NYeX833C4neQVlDQX8pYgd+Rboxh9mV9E6fM317zXI+
zVaEaR2iFikBQKaTL2CWAPu7CsImx8kIwHY5fejF4A/cfGuOdOJZwoadawwnLGztBh4nRfmcgOXy
GQsdZvpG/LVbviDGB8HUm42vyD3eEftqAMTCA1WCQ/xV/UntXjleXjzk7BdwKYB6ne+PGrJbtpeO
kjAvjfxRyVhMWda/Ein0VN8vVfuXhm/zhE/ICFk9XYRMGAf8IZ4xTUVpJpBWcShXT4SZaoVIHGPL
K6Pl1F2YgRlf8s+83csUm8HyDkQ5GeJ+EpboYp5NpRFglnCf+TVKVX2XoxXeSHF1dTDrXjlukss+
WWveSDBbASzqHxWoXi4lq9nVnIRrevWkiVcUkJuNzkGGK9XsfDRzUrVvMROsPqURtb7v26EKh5iB
kDO0W4EXeL1wODkdtT8hgtAOsWpH2kmeZSdpXc00Mc+sJvCRaWldRgVsYJ0exNEC1Um80FOj0Jwm
LlXo6uF55UlYpsoPlfmQcx+eqivFP187k3wbI9zW0JlvOA/lfEYYun7dLiGVQquS0kYCjPE2XAPr
sKhEt4D2aQuWDhuaHkxuG7HyBff+vpLrRcUVqz7J8v0a+v7mk3mGLTnVZUkjrJr3L5j4RcTsTva8
qzCN2bhANU3DeOky/o4EA65+e4prf7xfh73IXR08gJzeQbInu7u5SJLgbmX650/gWfibKhIGo9ix
4Pel9AoU/jrrG+Eie98stiAh5OvVYpeGOzqFMQ4/E6jpjulE7edT3xvuUDGcz9OwZulLqL0N+BnG
JuR+WQUf+JX1m6Tqws09Y5lvyQrXKZejcBiAHI2oGciLZe45zbvgP1nOdheHLn76FskSGnmWyDTZ
RX2IPWx+UNKWN5YUigG5kYSwPSv9ffhOm8P70TNCVsiaTs1GyLK9aEQc5J0Fr2Zj8K4KxazzYSky
vUPbX4cTUlhEhTRG5dgS75xJbV+ysgks51W/74oFKi5L1CO3iXX/2BI+u/ZY88ycNOrpGWdrgjAQ
FhSwy/TV4vlfwpMdvlqtXtetIBLme8DiYlaCbrA+zsa+voqexbwZO2jJpc1I++Gd3FfE30HlS/Bs
f3pjNCzPyOfkf68faBYP0u1HQVcjw05607F2+PvIMmJAY4OPYyOfdtkm4fNmDTJmIJRrmXzWdmV4
jXNXn2ELgUE7mepN4ZesxkEhXRQCWzAUlhyW0IjvrZsZU2P6blQSr/c+N1jB4zHg9CXggm0iKFkM
RdhrtOsMagrwdO7U3JAJMMTkEowhUrLugXX9tZ3jd+d9wRq2Lw+CLeBZe1g42WvL/O/WbSe58n94
vfDU3UcsD2oqXh0YRzQGGZMQ8GN/Q/2K2UVjihSLd57bqmHgU4Y0eaCwzsqa0N5+ryKXXYSGmCgL
ZO4dvCSkoL/Nu2vgrfHD6acQwdRDMP3qnGYizccucEkFDoC8cf6CKU3AyoWbH/r9zaKJrLWJgdDr
Fe1uf4eplMAoXRZujssEWwezol6IO1x0ZOhbmbghQNdOIerPsnagty6hNG+dAS+GhxyT0th+GZdl
W7DC2na3qYkKiYA5CbzmC4IvXOUA9ydDIzKjmkVDdZFMN9iXG9irSuK+eoI+mL9RYUhTJ7aPFq1G
3eDYHqSpti9hEt7xaITgWje0XjdL6KNeH7LoKphwDUbf2ylkKLLjnYdUoI4VuW7RRZyT/EvA0aJK
t8wyh8GIO3/SSQtuZpyZHVxvKb2gty8vak5h4rf/8D46R8xURPbMUyQIxarLYInLvzAfsPOCBoIg
qrbFAql9iyj6PCohlh8QFydejlZnuriCZLWkjsfYHuvja2KyaNxrIXQEtA+80VzDuMXt2J57wjIn
5BejTj5jQLaQRjVOULBzT5QUNcx1GF4h6fAqvjxbwUn3IQ+RpiIyHK8+3BwRcuipAmnrShZs9IRf
9d5FykHFnnPiBagxZujcbHVfjvyEHS7+Ao2qoXg9Pxi9lYtP56kxCBHuXNF4WmH/kuro/xj8Pn3h
eNaCHwdL6xdAPjCzOBYYzzQAtbX069loZ9ZstNFXQ9Glhwe4P2CwLdKJqMjrLqXFEWkZSNZAQeSY
c+RelElwcg89JXywpRvTa/RzVgV+YfNalxcOdoQd/RGQtPH+Dui2y67Z9cLo/Zt6qrqloTV8E/WV
wh4ZW8EAIoPTE96sRw+BjVpRiON6Bs3bvkNQ+FEGV+RdiyhledFAIU12PTgWZlQmPWLGqXZFqZUB
fGCWhT1Rr4Ws0ccqwLIOw+FrQjH3Kr9lbDY6l19xfdQipzG/XHfkwBAJ4OkV1oOsUkWJ5zDyi4BT
s/bQz0eZFJ4OL3gsuFhP0nP2bCZYiTO9aAoYPNMoMt66bTqW/PT1n8so4/myG14uVhjkXgtSPmHF
SSaNruWcCbLX3KwaP29db9M6CA7g+9Y0IMzOFRJxSYciuD4Y5eqpgEc/YDP3H2Z0A/2MQYz04+sO
3iIZIJ+jnwFqGknzc6GU8jeWVaTuVaj7iISXYTwraeWdhHw9ORJ4Dn29NE+XekX0rQKgmiZn1k62
cxQfyU1fj1AQwcgiOHHW9q2SevQKNCGcjYNJT8Z3C3m9o8lXPpgqmraXqwQz6ZmTHGslqQqrxlAC
fF/vln4/Lz5XwZfBnv2eurnOWyH22KLjXd1m8B23nZjHuDvnx+Qk01IPztBW6yzO2po2V6urcF/8
K92CyxMth99Kv6BUEU644W7FaH9AdwXhR+smgbHwC0bPj/7vP2RKluy+eXsxEixqQIckB8+0GrSY
2H4JIKuUVAQYOZwnSX5A/ESiY1ZrRtNG4OJ53HYhPy4OpXvXN0rbcxY1ldcNCk9QurqiwB3RsQNI
oZQcLRSewHoDkp3EJj5UKVsnV+icMxZOdlth84i/XIn7AG7j5qKbNC3XCZU85XV3O+glQPuIpbHy
XkT1a38WiKSNHCKpBqVvwaE95496Sx3UHe00BYjp3YSOX/kxIzidu3zoJ/HdDuv5qtXXE3UK0pEV
ziqzmXNGfCdBoBcEJbIY7iqFTeHASX/mW9QwATqvSw2z9SaHP4gWdbfHzzKBRoDouifS4UOIVR0R
h+pKUk3rNwskWb4g/IjUaGM8QIKrVDmX/yMbSQKFfAWucNjdHKREfhXfUuLg9da0WGFQfbdULH52
QlfMdwIbzy5wu5syfa0SZ8bKPQ1fRd5HrAQgWyxx4p9Nc5FWPmz9Jh/E8yYoNW4fn0UyTefDWLeO
Hn1syrejSun/MnzDKmQbOtXd5LyhsxTE5a4nUxhpGLXfgQst6kk0WTq/LXnqvp+TtHvcMoJkHVm5
655SsFBE2chNDJXtHiseJBYN3ipgtpuahmo0Z/zqEaQI5SipvmshW9OWXvjzcTvWF8FbU3Ur76jv
tRzpNe5kOnAaDDW+4v35vdAb3vSdAtPvcY1KxQYu2dc0EUSGBXn1jHI1ZjnEYpiPaRTpwtaiydS3
gNUVwIo2j1xoUFlTmgexE1a+C2wY80xifRMlYGc8slEk7O8fcqt2jCzAacYsipQnDWMJWX1YbxnE
lOmSMPG6HtRECpLufc53gqRgov07P1N92UlAN3KBFOL9nghjhdlTVAKHWKk9dvo/BJo6wEVXsHGu
4WmNQmrBBd9W3f/dmbiStDnSqjodcRGaaxKxv0giC7Cen+noYDzmQIcks76pfPgRMafy/KcS9jw9
7P3loe1uyivIeFOom/V1CeITEPOBOBIQVJ772J8mO87rBokKZIAjU8jiDOOz6FQ/vBqFumP3KVaZ
7a5wzvdJ1pO1O5qmP/VQAr6Wi2Y+b/+/72U5VQ4RffP+ekm14CLQjfsjT2GGLbTXntSYrjK9oKLk
C4zw/JMymX04bh53fcCpJtGUL2yUm1AGzbRxlKLj2ffRxJnkMEu8/tU4IqY+totY7F5uYn3I+1cw
q3wBHqRzjSAbeHnRO2TwwVT+xF6TrhAr/SGhJAzxhnmqeB4nyOzs72sODudvbb2jCF6/q69w4xix
p5E+v6Kp9B+G5TT+RkM/oD54UuhcKOlrTHmUiM3KY+IhQj+i4HeUCfbWqWSNhh3MbrnC3kJj02G0
veLv4OUQ2MsiwLUY4FJMGNYUoSO+XhxkM4YLbv5RB8LPQ/q9nOx7sGkzmTJCjWgYxHbpXONY6c7p
dWsMB0xMzEZNd7cQcOtSisKdfrmQp8uLL36Ix8IWZox6gkgHJ+Hv5PU17wZJfZklG9N60DbCSO60
h8uCZkW13WwRrNUuVqRZ41Lvrdsze10ucmZZ5mp6Pk5Bx75Cxt56RSIbz9eblgsc2l9yv1T/j7uy
dknEQruiLg/2bPxQuy4CkdmqWZgj8gXL6clAZk7GiaHHZkEqweMLAK0LWtjsWAbnc6YCTAArOYR/
BhyAOp7cySqYzMXObwlq5hDgONVcPdE0u5/uOqS8VKg+nn5Ev8+p8X0A3x7FSllW8+rwdgs8BT2X
nCabXasow5St0iGKRamglr0RaV++h0bX85HApK1/b6GGj06WIHlW2DeN38vEFPl+QpBHV5LONpVb
hOingtdLtUuG3gKhV/Lvqas6aPYFnkFOlTR0Po5gK+mnKxVxfZ2EioobKtU+nnavq/oU7ubmB//F
y9YrU3SkkQ/8HYhRw5PgTOngi5l6eauvAgTM9XqW6PVT0GHJtG7MGVpCh3fdkmKsuIpLdrT9T5wC
zkECXxSK2+UBGcPk4MHMRZzvdwDLMTW/kir71w8477J1iqgtfNOImvhoGLk+0t7MdU1fhlCFKWnJ
3lTNZQGoBa+gNi5DM2Hz3GlbTtpxba90L7IYUjpk8QEoeFnDNqYnhlFPiD4UdDSyKT2luKyEPzb7
nb0xNxUKBXt86NxlF+kT5ORwfppaE/9J45HIzgCvgDyNGbukQ8fqU06lTKGQjYe+hApRJ6km5GOn
ifeeC/0gO+DccIJHhBJYezZCQUhjjyrMdDZfiDXwb/vt9HEK+qxZmDq2bEvCNNlBi0qbKOqBYD3A
yXYqN+/Ooa9Xdghta/jHhvmqZDL0Gmqb1TtAOExm2G4ZBPJjyXiBmypF1PWcENVJ33hF9VodtVt5
T3q9lZIalfQ9iGrdxli0Env4nFNRgdC2+pU+JaFX8HNWgp7dsJUvaFnEmy+OMJS09qgcahurXvKE
ltaH4o0JJn2Wb5RoDmJOwcqiJyt4G29x21ykGfRT+C8qK4z2rZeO5R429at0+uYEHBOIvR8611iU
QGAKYSJU4Kwe90Kff65w+zuui5GnWi6PuOre2nEaQdnmsTOHvVFYAtaWoAKqROzuW/D8+Ada7pT6
0wGrqcW4FEAZKH2FoeNzw6eCByJRtJBl3uMXktKWWBrIr5p1zxuASHrB13LWK4NbjP5gSiJUF5Bs
4eKpbCcJhSOaxvGGCa4Bp6vIyLSTzqMWjly1vdQhEjw0f7QzmsTQMfPEh3N7Jo1HSsJh4YqkoZ1Y
xdt5sGgCOG+aoVzgs4WDF3plSGCxDGYZc2sTw69onxmhOD/+Oc9f7sIWt6d1PClYTUtYcryEtOGg
sAvQmtYDj31XTb91b4HkRVwXk+J/QvMoOLaPS/TO5kY1psZDIC0HBHboIhUpttM2JHJnQgpvmw7n
weLBrmmGdFH71+17gZs4Z9o8olBUB0W10jz+MLZMy6e742dHgXj7hkXkWMoyPuR6DrWLUDwHOFm7
HFmkCMu2PEVzyD3+ABFOeWzetRbLKFJAEfyatc3QmN6uOuvmNwkWmrXnESphn3BtHiQfB4ut/1nY
TzuJFBiJmzsDhK5dERUhLu2o4tGVcURiVrzMFenxhsSnMJpm1lGQRPUUgEXpSqp+zv3cYjmnBPqL
YnePoRB/l5nkd3pOrAAMCggWQ/Ah9SqCjjwBGCgzlUDMTD59iMEPEmOOzUyV5NA5EZTQtm8LJce/
8bazypSC0eNQUCEBGCjgmgstYTSuXIwQ40SAeGBFj77nkNrkIXMukdK3g8GgK61One/qlzPtqRDy
AuMtugr2X/ErEayhn3/y9SUgWZTmaUzBDI/kVAjUMvn2s784+BCKg9gp6MtM+M7j9C2QTQBf/4En
G0bURoFCkJLYiR5OrCKl9NNXqL4/SG9Ku2yBTDCzWg9ezx1T7CxP9VuaVH8zSTa+ltivDkAvPqHX
87W3xKn455eHz83rzW5oQ4ZVsUHiLPZ6hPj/uG+C9qkKn1T/1P7biQRhNrO83jg+hUpS96QJWG5z
JhGDeupmXPl5735vaSJZhbMpd1DEDlxCRYdw2nL13Zo6oofKB3MQHXmuyM6ig7kStvrJ1PtADm+b
c7jq2L7bhBUhBkGXq5Zln9N8RuR1vv1NoAGhp5LI/hOulO2HEbNqBcn2XDs3t77kxinH07b/yLqq
exb9wKz6XkRtTksYVwdhS+zaj/FNquh4JxLQhl2SrlSvMs+NQhot7rThj3/XMN8NLv3CwvKMIC3Y
HRPif1LG05duOF0KmVyIHePCaNa7KEPFcjuQ0xf9dXZ16vw/kUi22LWljHzbYBM333ziS8B8pp7Q
AJftU2tAouhS3/3hLw+3j7VvSdR2jrl42xOoooGJcMNz+W4wx+xS/q6TOQ+lm9ffNuADiPX+7w4T
qEPzQ4dG/rK8f3KtaeL1Xx4l8kOdrXHhV3ty4VxgpMvIbZj53Ik4Td7PYhJczGGmYu1m3MAHxh1g
+cSKWhF5D7ypet7G3/JoynI1NfFQ2fBhxMYp8x1f+wDyH7FIv+CMO1F5g+uuhJUUqdpI+WRvlZF5
TJUYWDA+fOhGwNZwxHX01mHXqzmFVcvNBE6zbTNfXCxalodRKIiez/1qMR0RLtB0OEXXRzN4w4ye
Bsh+Ye8zd5GXpH0DhIF0blQCk30uExxXX5+30xCMlggLALfCo1X12FkxJlnZLJRCOx4OJLn1hfhl
r55TnfsJbLYoIOJkgMd/+h4joocqASs79vwGQhp9iHnvjI1+ZVBSxvjKW4K3afj0GuuVStb/6++2
2qrUEWna3SOtvzOf/MewxDy8rA7ZAz4VA1nJR5cRSTJcsaFf/5SPYdHNSyaVStdDLVnWBloXNbzH
gzgtmPnhpLnx7ZwnW8rsOuJ+T5BQ5m1svlxyb9bbVQDzandsj/TQZf/xIAWeRMh9L1qXXFlkMUUZ
MMZhwuCGUS2AC9jzY5YI4M9UAzL1bALfZpwPnHYvTxOQ3cjHl4mSsIw3g1AuNrAc98OAuUTxbB4n
sYX3eBLC18yDVOPfmYfxC1ryS9Qr/HwKdoTw65jNdLB3NpVL02hNG/zAoDru4WwkcPQn5RfjkB1n
nBQTD8b4AQN+ef8bLkAPxk53Ue/trpGDN8iFTa5I6n999lCyypvHHMnTgp9x7ni9aEKNAdVpVRbQ
cL/ODdHD76W8vUaYHBjGJ/NAxm2L8cJuhU8p1JRLxLNREnrByXDls5fiWc5f2YgETSNT9gkKivrk
FEvTN3iRv2ZhLikbupOO1q1dZR+jZ5ZnC8i4qfpd9qu6+kYcGfzczxUEU0y44P3Ec3kEZMWNNGsN
9xI1p3Zihl5E6ZkrGVvyaLiu9mvF3La/tcFIkBie871Iv95R6rXVnGPbNj+LB92OdKjEIvNq9oQy
elaleJhdZgEEI4CNjxxvIoie2TI6UwPxOYPpi7jebLMa9a4I8PWPEi6xLlgUSgNJWkKaZZGquNjO
jgGF5sHEjUVqqRwV+rW0KcqenTIvAUj6/gwqb7iUi463WWPxJX4MA/ntymifvjnVMnzzAXtkyr5U
cVRHMWn6jrf/qLQYAKAhMq7BYBYLfKFYmQP9zkBd5vpb1c7VCgjtoUGbL1ONcLxRThPLz1LiHRRH
BlniaYxdrm9H1sQOKVCd+dvxhhSNncXu+DQUpjnwckEVCRIBg2Ebb3OYLgJc+3HgVymhnwmqq2Vw
s8KzJDcGQH2TwGxrJI5HzxjMR1/sByMqmUkaHVysc/FSCnayA7vHxsddaDInbhZyuws68x+4nPOr
H15XPLz+VK3ePEWld8YtlSwZxG7xaujfEx+Kzc46DfkJ55LsxptlPY7+mrSs6MYvaQzTySZIBGbr
pYVUfd5LiGKEv6/IfkEJ01gZq3OcBLY/DTSUpHV0pQWKGUwvbJqbFgG6vXWY3QiTqYCtdQQFlkOR
Xiz7EoQTZICBRGmCcgOOdY51GsVxYIMZ2GuQKLJqIILkuRSzS6BzUzj/jhqJ/epoQo1iGYA5bzmr
cs1Wvfe40DrndGZn7JRmFnNelxfEkKaVEsmQBTwhwMo9qyzzEvHwFXWaQkZhVjngQXI5wCGfdbHJ
V+VXoQB8NXIBfUy5JntNlPqN4n7mGEOsEYGV7wdZ6FARUEsKYStmgsUhZIS9K4byKpS3tGGj84Pd
nvOAs2e8RnhCXtZLDiQBRyrGqC3jnBMlzDglpgTti3x452A/UY2TPIAoDD4mjgpY/perTHYznDKB
QjWmDx7c0sQgNSdGpT/gHQP8Q9bygbdHOFGjZ47Jf7qEA5IaMGa6bEWyc2j6Br39sFEie0BNdPmd
9hqa34yteddceGcIdcYtUN3iP952Tu9lnXSSTMX2gWt45lyf93DumakwmvmjKxUaUgmCQLYLa6Th
L51GzCZd+KqyJrLRdm+syBdblBqKqTue2AWDxuSDJOXrVZzBN4R8hiB5bN/PEvm1k+FR6bRruber
uBGfCpoXB6XS9fY1r8yd+xVVzEWuHFw1W4Rg3Dl2mJzWeT0JVLSoJyNLQHy07hBbGW7o0iA9NZPO
eATg91e6kSzjzo+sNSODGcN56teX/X2MazPN/BWICHzd2cOE1v63PIe3Fsfq0UE8P3oTQxDVnxRS
ZJZG3SLirCqLrzXwzmgzZcEzA7GsDrWEBfjGuyp6+kMFZnmLygdahLrrxflPrlB/xDIQm1kf2SS2
RspvdiREJDzVn3eaSxQxOaHl1xhDsQKx8Le1UolT+S8gR00Sj8e2hsCatpwTrIuOXC/rRTepgM09
0UMFOuSwCJTVo8RbfahZtGDRpGKoF9xYH+NDoKLZ/Xr2Pz4Qpqbc/gtY2HxeIUvM2RJJd+lqKG+b
Hil5T8zsfsatAQEehkOMPkJX/o38+mJ1iSuZxB48XykT3VJfpL3HnPYsEYm82s2SHmxSgn3b0ll3
Dz5I7gRCbIlsMmFrnVKBPpv26+lTufYLVbV8Z9TIKNKmMYp3kjNWnDMtTfzhK1cRMuauTYzPHp+y
64vYrPQiX+CD4JAHI8C+exsa/E0noVJ9Wo13gzmyqvpldYdjGFJIp0QvfL9FZBKfW2TKtuI1j+Ek
OAsS4er2DQ3A3aRfLj7De4k8AG0CM2ojp6H67cu3pbEWzfPzbzfDM/46oyBIgbR3GZNA345E8Lg9
CDMFjO5dT2hFjaqzCaQiEERnqydCanDl0Hov1KWvJvaTXLrI23yNxw1wpk8gzA+/RlRWLjw/v/Wc
DoGLPQsjBxmJrTUc1/LbuiyrCLDn2WaNpdGGjiLsGJS6reGzSNJEftH1W3G/3SCEzJbcWTWb6PLj
FI0jQ7Scrg4UOwEx4A1Y76fhNeCHEsANC2e+44Wi6q7S5bUS2IgK5UdTyr2OdxYPWZgmVAqPIOHC
Ft0FY/F/0jAXPnZZWKEGyYjvRJV569yz1QDNOb5dW5rBU82IQAjam37yTRJvvDZYFXjEqcZ7BIBN
4DFUAu4u0SnvBs8NRF4xQ93Ymj4iB0+hD+J0fE+bK76poQFglMMIyGJ7P68uPjaIh35T6kJrUi35
+8GrErxa6TQPC/POAsJlSzbs7sedbmh0K5SKWxRO9dSs+dRnSR0oUNEo4SlixzTpnMrJ3gSvCJSQ
Ae7DRJ8NvLbzWRYyizd6rXzA023vDkbDeQYpSlAMs8FXxhkBGgXGHbCA6uiYUtV0XEhaSKeHE7jq
pewUK4wtWGQ66sLC8Y9ZD2VMxJ9u2Z8au1dyLIhtbaBuxO/o+zDzCrvX8NHWvex1LYUV/sX2QaPd
/Ki8xe6JQoMunhr/CUIER8XCCFJ5dv1VACA/FDg0r7B+6FMcunS2b8OggLk/XDaFaz3sBuBVXQe9
rzl1GgHvshGcfsJ9sZXkRNjFmgszqo8aiWOEH33k+NkwdKu2fuNLQr6+WSSWo9b4tCdCfdS44mLv
O6VB0+mPE8VQiQAxdlxZQ5Gizy5s4lC39hWkHOYMDk9lxAqaodAuzyDi9/WLqJxWsxwPfy72jF3H
Th0bsybFc1y3Hj1gTS889eHLcJTmO+EOq+eK3sqjnUgzMcRNFm4GEUsHEd39PHsoPNQE7ytJANtu
CQMsJwvAHHlgp9MQdObO9hW4Df3+IOMZ7Eom5o/dh4Y5wLqNjxD6zvwafwPDY+2Z7PGqczPSKihT
lncdZ08aJQDsyjhq5I1Utc8B5aN4VNctQD7NtvUknkBdiTyBfxjfZhcMNyzWV3ZS7822es7MHGch
uWXBsomM28NPZank83KY7D42W6i17zSxLLiMQ8IzKH+cqVavhknXgXTn1YLhaYKyg61iMm9n42/Q
/EJLq78KxsUaOgcjRfZGFMq+KGDS+5IwcRAvE0lrQto4cCi55uhGQ6w8NjWKkDRmPc0a2DNXT230
DE8+8bTsH6mtArPnAUXTTO3T3pR/a1GMSs0cqh4QpQzPpwV6emR0lA0Y5APkYeBUsfN+eTCWMvIk
G5NTSxsagoO8up8h2wP24CU/qEujBZFc3ZghTE4fusdZhhmFihTmjTHWioIDzKJK5TON3rP5E7L/
Nv6ekdDNQdNuVN2w9mp3k8mTmN/ASjIIjUYnwsM2AJIvHcLABD6lcSRihS7SPxvzb8aciK/dG4IZ
ZOTWVO4NHZKKk0WTvaeVn8w+yscvg332xHXN/nEqauebxMJLs39kQDmnMCp3lq/jT/EnPrFdb0u1
iPaFNdLFYshh71Uh/SO4E07Uo0Gft6LXZs47yjwa8VqG2Ba3wPu6fI0EQOv+P/K2yuEJRgDBNIzh
iAQB2+rAhEapcqUsuw4YagC5B43qoBNIyGOgiT/+21Y5X+zRp3O5IPNcNnJsKUTgO+TvYo+XlNKM
1oQNGj9tOHGkywMKuuIdR+vPYABuh3UQEt2dMO6VgrS5nPUTfuS3SCHO5yRLlMWKlML6E5annE8I
rifoTr594YeWuw1SvolqqThTF59O+o3McMDH4XnsdyO+Kv+4n3H7iZB9U6jEApNV6HsSfel0O9mo
fUAw47XoNXhzMjLioxDrTtzjHZ26WeLqZpGhgpeohF47WEfVXHez9tNqR3O3U6HNIflyQhhT7ALE
cXHt2FT2mNE0Hznc/NKquJrhUqHciT/RBdCHRYZYP6Y6niUtC2gbhIj1lkA5EpJ1ctdJ/pCOzo18
s9B/kDjILZ8i8N1b2erI5xISE3pD9y5n/V812p4sYSa2HRjg1rCTj5YIGs012AatCPAb2ynw3LA/
zfQAAi7JFUscBvF4mU0wmuGl/5WncOoc39ejoXzLGWkYTCGr9TxaYqbD7nybRUh/UlYUVPKWCRCG
y6cJ6nfZBsH/uSKL533HQss8XtuH4YUs8/un1ihvdzBO7D5nKuZIpXklBnptUgULBzhWsu8VxXFW
s/EQBSoWEEpNhw5YK86Pr9dE70dLN5xXhbXOPY4qrnnJRFgS4W/sSkFyB59WDkV7FeOXWH6yZeW2
0G9Ul35KnmvBHsBNR8r0U8TIUT6YqikUYtDKAz7VZjvQxuCy5YF9sArFa1PfWm1/WLLI9GKoXuRl
3ahYfuBYqtfwrbiYpApgUzTXgOHyOTm9Ui+meVCm/K0jVMWBVrZUqBUct8NRbZxgOZW/qfdWZDWB
3NWWFlbxLM6bLVFLpVGREHJxVyPi3o2kWzpOZMRXy4apDlmQ82VVCa1IczVNHfNeWVSIiFyEfE7h
npaJ95bZYtCYfRjCnKNabF1BWPvXleq4/T9ikbJOO17lhDdZFjVqB966E76yhXv9tS5lrecFH+CC
fSs2JYU4fV27lBYQzMfKPXn27GaYinO6Mx5HV2kZJBHamM50IQLixSxDJNQzqPMxKyaQXgQwGmf1
wvyYk2ywsHeDlpqqrlpyDQcnrGFyxbph8ahEjb3xoPh5Qm1l6Fq72ZpBPMpGA0kxNKaqN7+dljm+
7whYR/Los4eHMsxy0/E7bsWMIa+GBE4+XbWYzdd7b+w+LUGFCS4F6w/rkjLpMhXKk815OBDcue2Y
FRJmiZY3+vavS+CyHoo4uHfr304hZW+57XF50t8PPVPE4yXc/nmqDKhL0AIN6jlQh0M8V4TSbPuZ
7N/xGhcBzuGbs/Vy0cK99bBFs36MNU3GhKmaIddXRGIbJ1y460fAgMlcvpzp+aWJU96/f7rocKjk
DQwg22fTCdarad/2SI9h0yLzl2yGGRBXZLYVpQ+3GXO93jiwqrt77u3EKDfcSkZjqcqX5nrRwTmh
tMYaHo5Yku/8vLvMc63IYEUKZ/lVEoptGgK11351pzOxghdUXaD4KyEa2kbEL+XQGMtwdAXp76hL
F+IZrsJv0wiEUKVud/431cS+s1bj7Ag7Pb6mMfciPcUfwfuGjtZnge1mvXv+wSf+2FcsYdFnC0wk
0Ec5RMqEB3sBjexjINPCXIo7k0qNEMQRW1J6nphYMREYOaEpUtHMjbx5xVWAFti5A4HM9TYxmhf9
rRq1FZsztsLrv9MZSWnqL7VF1ZhvYbwNcLJJB3mKGpQ26hFdXRYwbMyDWwN8JK10yi9UbVxvE8FR
04pEr7kYNXWsCozu1YLGdvX6fNdgHuO1l1iQGhZtDScVKe9XbnLs/d7i3HGHgkDefpQyxQw4rZ66
orX3SwjFnj9CeRlUrpIsl0KYiSIPqPBbtEWzk38p+oaLlsLLzJDX2s1TGIzU/Sacb8WDTCGimZS6
gtC2TYzjKDPYlUtEfetfk7iO1lAj6fkkXkXm/uT3qQw/QRm8fD4vHT1yrwm/wvjRGWc50cGktleA
KG/ohGsfVW/wd320SUsHlaxMRCmFk0Ea/mbFegq6wLIVHUgQQuoS+iEWgPhxV0siCnRxVOG5ZFnw
NBIgvzBO3wgmKOkpgHdLSuQnEnOl1LuL7AFTHoQJZCZ81FXXzGvtlozLPLxBymYaSEyBV4zqiaLS
eK3JxSlt3PtVHiuM8yBgRtCHOk3awiwsQjB20cdJYLlCGYt+AByijmJoFgJvu9uUiMEzxQkb5HyR
LNNblUrePz1s57mDS9tafw8ekPfJozO4TfiiIErOTJFv70mld8MqVA/tzP6gRnHzTnVQJdz3rvFZ
wpePDim1+JIBxujLTWmn/sw7wfODMmFnreDyWvmf6Gbi0+NEpL+wzEF7bwop8SNWSvQGMJ0Bx+Ub
Rzc4PJavcA/n6VmrK/xDRbNMShrSXCedqm5qLdtWCXlJSBo3CqropPUnhSWEvb6jAdZUOUUaPMXh
WFUQjWE1KKr7JnNfBYJwYuBstO27S7fhWybKQUDkBt+f2oAwXazI1Vi4CYKpzNoeiIGeqerehUKO
mP3gg3kT6Ok2HHa5woFN9jcelxBQLVbJqYJgQFzhEMo8GuvUMDaPKNcGIQIKpmoXwJ1cvUD3eeX2
qkeDipfIJUQSKpNxVZiKc5Kw5sUNt3jJZritGkEPVUPxkWTGN/rvkx9sKcNet5pSUDIH0jIS7cYO
v2y9cVRtbCl4yJfJUEIKBB8pmlF4dzX1oRYdc8qrc9rXiSqhyMesvRtoNtUCUU5bMm/xQE5KWQQ/
4/yHk+6+COZyLPC8nOfZLl0rxr9ktglWNd3GOBKrEITkIZj2ytT9vUmFMjK9yDRcthldScPVGDyj
t3TFLD0y7yUmDM00HhmUzK13N+NfOoTiqQIr37WAh0uWrdD6LDOMQX7cNbVl1lmOT3Hqz6RHtvTs
5aVKKJEYP8LOCCmcC6g6oywtMGsoJ3NZxHOiVx7b+5g1DMViTvDDnnHCdiRik8dshWMomqLlkZod
HkGCINmVfd/FA1XlpNDFdwg8z7uBVx6zCEPdx2e47ckgkeJALGuGDIx4TaKCOYYmKyZIPN7So2Ep
dkpPCoxZR+aRowoxAmPiQ3WL0L8HOJkkkUQ+5pUERVyLakhUfycFAiI0oyQUk54sw4plCZ3A0Usb
7mieAz6su8fdnoxrXiDyR5Y9/OAwO5Q+auG0rIw7zhzFPwNGCYMXJVj0ec4hTPOPLtOSrDMKfWSJ
VAuOoOrev3hq55iUtxzcHgkKdsow9ERpHHisjHygsgWKyW14hjuXQyx+fCuorzVIR2Q259ShmVtG
3uk4kebJ6UBj2JeUPiR4Q31EXl9VioC9RnnNrYaSS13Tz4BL3xscqHjYSeAP3gd6RYVxomH8E0uK
2VE6Wo1RKJD0/4WzusA57mfi0Wnkm8kzcjGVCDavlGISH04OFPyRnmJ6N6xWKwE9suNbUWHOshcr
+9r0ngA4UXKBjELOBXEruyLoe9JDnEBDMrMG0Ho73QMtbdvg2uUyax82KguPwMM8PGiS6afKASOw
kGIVgWNuCF60NR88E1FJWJZFyuoTPOZkMr29WNGexF+zebPDo7kwI25hYTIRpE1qqxGeK7ssmGSF
DMO58RfkDUv9t+X6ltzVZis1gjhsGrbR8A7fzXgiDswZBdibVdKJXBmihRqmy8iNRviVLFsYH7lA
aJFFlwyP2FXcC6JetaTeo8NC6I21SW+nC1kqwkYU2E/xGQNEsojPw3cclE+UPq2gA4FOMsLKmSCs
dkXxJECoyXRa9TZZ8TOzhYb/B6ztNCp3zqs9WFNNCeBl+DvE6NT5+FZgIDxkThqi/fN+iz04XBe8
8kMvsvUCbf1ApUQU+7A/yG93PQG6jKf2emRwqDWRKZWtq+hfSQuCy0G1W/9rDC2gQwGRLkSUkcBV
kbcFeK3ssstwXAAT0rSESwEcgfE8xYXeO8IOxIpx593yqnOVev+VecFaRiQBdKaYBIv/Ydb+0Wi4
cVAgwEzgsHytdvZkvhQHoUXVubgC+NgaWsQn3P6YJ+hwwaxNDqbMJuPFGyhp2GNnUplokkSvCUdp
aR0qu2fKhCgpxBboVZNIEsy17hdZdKdIiJ9OfzF4AN0/Yh/KiowhNy3mc3vLcfGMPjXcL8ph5mET
NQ0korZiUvpOsskjDjYp201HExW0ksO1lyUdv6QAIKFbXPeC78WF4DfMYJkyz/gG6+ypFKJtVjr1
q8vp1+QWmWq3/J4ZM0elKLrKv/RwiBHrzddf+r0iyERQT1vqIRed9KHaHPWbW6FhbC/5PixLN8a0
Zq/ljUUtKtAf2PhgqwLawfXcnuf7F+cFUDeifNUs8tnpwOw4U9UxcOsEUkIqp9lwCf68fBvRI7x9
DTFGtMY6vo4+qERnjXkJtdq8GOZqKQ6i79Tj00/V1J82h69FuM5pC+jIe8G/H25OYAAOrJEcgFSu
8GNtAAL2r7BpFPDQ/fS8vF0mYXct47quszkSqnYJ+A6Re2o7Vjw3s04j0XgnqG63Ic/NjTXMXDAe
MgsB/YnbfhResVDNsBhfMrLFQzdRRYkOl7jvHxFKHSazQ9ldXEYD0u3vTr2mp6aJtqToBYuBfuqs
Shdnx+2Zr/v0L1U3VousXvU1RIg4Kaj8duhhv2P2uA+kNmKDLv3apmsRM7qnW3mAkoKnkShm32kY
kp1gziCk3gSE05O/UuarPHXp23z8Y1pV3FRAl8OZn0hgxgiqZqpkOtyZRCi58DLw76dSe7un+upw
hF+txeDpv6BdFiIi9MUHhmPAY2fhh1qEjGyMhb0JUcN3i293TGMY5BqpmVJ0WOYRSN7o76BG2R6v
xsLjuxGyLppprg19mh1euviLNFXpCneUlM5bdMrJFxh01GB0m0hASKmlF7rooY8DbHqzt6AaW9AW
2gvBCJ1LUUNaUmgQQQdp2iSBXHrglADkI3ZTLCWOhwbRogaIQ7K9VpMoo3zCrCrBhMEPoK2HDzAF
GVbZCh3hm1C5OQQn7CQMK3uGiM5g+Krge4ZMyG9cFUeHK5yAWy99yvST9YTFUhkFO4IrR8LGC5hW
pIiNuS8rSNS9jF3+wuxkdB8afi9gK50lRG187kJUZoGSu2Pwpi2yG2ziAs3vsJOvIjTryEhKi1Nj
gUWJwte6HnosQFFkLMTXYd+mQBStoz53LOVc9A/QO2ThiIh0H45jU8iL+QZXr+E+4OKoD9jiAmCe
QMlU+eSqWBR0ZekkvD3ieTf2v0vhnCMBL7xo98Q/pS6LxgsVJ6WcVT9DCRszrhnBACI8845dCnjm
MaD4Rkp/YMs9mHWN4FxX7cPO1GVenbdPprHIH3+pN/YWfdxRgMR+sOcrz9oIjbOtPbkEtRJh0wvg
R4kbsIJ3X+vj63vYe3g8e76he/uz9ZPHjTI/3vqFym9J3FRIKmEIrBGh+B90OGjWeAkTY+241NB1
lWat866LCGelZVjlUklUKyLfzHThpj4RNxzkWS1uBDXipT349TpuURmd56b0M1MNt2q6SCjQOyi+
AMYaH+IZC0uphErsEem4miqxa3KKQX9chdcTHVenDnp4I+sf08plABntlWhDEDDk48smqVeA5yGY
oLRUsk5aYlO5N2HH2rSns3hVcwcwU6C1uoJwcWJiktqT66sl48XcD8VZJmD5sYRNjFZFrIm7kKU2
ZPAiPRbmt7zwTJHr93gc3Uegp9IeMIIbDRMBj0isow24zlH2fayFX/I1IBigoYltXUmT5rCqiaTL
dzGrIxxX6RrNMuoZexX9H4Y1oDOc1ZSrs2oSyO8jVmIe7UiLA0EqD01G/Ffd9F7T3+7zulGWM2Hd
W4nV0NZ+khKWFrLa3sYOU2XiUvzekgQ5qa70eireg4v/cA9ZdXHRn/4EZNVhoZXvy2Z1Mu8aV7mn
EG/JWW+f3CMgB4mzqdtHHMIUOlDeNBHaqCTFMBex9tvKGDksKrfB+HYZmnhWVJtmzJL21yK5G7wJ
Qa+t3p8KiYDdlfIOPOxY9Srz+LNO4Ts5VYEvwIcW1IDG0rwZI5zTy569oZnfVc0w6HwBY1AxHsaU
ZbHrhGPRsTJ3ke0SPTnlTg99HSafTeOMnRO6/GKox4eXcXpiwkE18PviKn4JS8ng3KQfYILoz7qO
Pyhqrq3pOzRgx52PFEtZPgypmmadEIWKLE9E5fHYra2/2Ae+lN/1ZNpmDvuECN8h+au2dYvN77JW
SILl6flKhL8FaCFqlCkE+3hQMsehjyzSicEDcF1XtbOAxxmryYkUmHZYS8fOz2nQIMtlT7G5UDsU
4+lg93+VhU0vyNrUEo8BIQlogUw3oa2Gaa4C4HhlFKOVM3i8ONBaQhEFqMWLdKpcaP5d5A/siLkZ
o/NLWe9K0OpVGJXwpoBq7m7tHpY/BLWHIv7MJ/Q3n2HI+qXZX72zSk2w1YonA+2+ypePi/ex0mJ1
s7R7x83/EbHrkChPQIKIf72OT806uDP3p5Jl2o2zDczSHUStQgUvkTbneUXKuPf6xKI41Rvluq1O
2MbgT5a9BACtT+sv3tPBKoQDB4vOoq6RJyCGIOMiBQzgNSVzlnH1fo1BUKUwLTrCZr/3vJTbFs20
e22ukRS4mgDu1ey2EtmmWFvGCaToZnSEKGs+XM19bZljwhHnHRcEp28z1xpEHh2GaMJIuUtdturd
EBfDaUiv6M6v+Q2QMhGnREhI0uPjGvyzNof1iQGBe8lcJGJccUuZ6l/vagb89MQ1jG3Lp6pkvVx0
WgFn0WegHxYvXlHBrHeDQ9fUX7DJcVWTAQzCdcHhrwXmL2WPDeTH9sbf+Ic+7bKr412pCureoJXC
lUpGYXiVO7OHvhSHs8Igmb+SDNMsmFkAfi6ntvuKWYFc9l/YP53anCzP9rQ93mKo4J0QuYffoQ9D
bKj7TSGmYd7CU04euvLOLhGIDd1+7eVRdgsrL3RWVG1GMPIqS8Ftd7AxNtvSS9UyzMcwoYjQMzhj
dWafJogbzQ7TEuRIelw4Bjx+Xym+L338+84DAYFc883bVLiYfwEwRpKgTEH7UrFX3fgOBYM7HNq+
u4REzOw6DSOxkj8wjvXonsL3JxrFkOdU2tywQT85J1hqiFlVP8xYaL6zLzzdVrpwnvQAL6dGvuR6
g+5MEVP5BapccYFrHDhsfMNjpv24mVW5I31FzszDs5MCweZrNVrzlpHsCjl0rdkoH0emiGwrHAKs
aBJGv+bHfbr8p8hQujlbDO6K6SKBaSZ5bhwTKAMl9Onq1LQ6ddCg/af7dXHaay8H3pJ+hdOZDbZ5
OIE4I4EwYv52t/I7Qj8Zo/LBUiz3GLl+mrxIy5TUJCPrKB+xhtd6KkQI3ZujlIQ8jU130pn11kEn
ulgA3pyqOeCqurE0McLCW53JoLqZrIgR904cZwjcusU3pQIsZCO7AzwJkRb8WZiATJzRVpSmCA+8
mFrfZQWUuD+CC+kMbNlX0sLwoVdNGPAvPWzK5hnk72hjdWx4YOpqwvvK2ryzT6RmkksXSXV14WYF
JHTqp/iJvewTx+xI62pC85kxnx42N0hZPhj3Zj+kxzvUGBqwsbVTj4lreFotUQLsSNn4Lyajj3Uk
Bwr6tY//MOsToMMY16uAjG/WP9nRYS9zbHXiOxJ85li+ZISPWGUQiufOhrC/56Of3TLH2epiLRKk
6isl0w5rdtDl6uuHzi8j4Pxsbuw+2xCwkswyyoTTfSLJz0Iul/FpJwcrxb52vOB/CfvMD16iJmKZ
//vBdsBZNGLGfh94594YYsvjQILF2OYn/Pd7tVtFUn+jsiWHvlebWOAI6m8ArlcJCvStfzpl8J/h
qaPbIaOjTEiJFyC3s4qb90KPNsAh37TNYMhsHgtAVpIwMaLFH3QAtXLfnBpMgg77rvQ0a8Mfsk86
m8Pi9Z7xMkjsuBmfl3TnIvbOGWVxYBCct+wuo//MXgdIrx8LM+GC5LnrT7AZfjVNmHP+wBF3l3mG
aXTe1Vy6f8YKf7POm1kFPeDFz2+pTyWXow48l8Q3+Usey20559ObQVaKLI0mSzqTxi5lwSpv1nXQ
B6alYxbRooIT2I0WX28TSVwBlOaYwrTQImW07EIEt6gXc1/pB2FGrfMxy8eyk0JjzFNr4jP4aYUH
CNizMxmbrxWu1O4CD9yXz2MjJH+AfqI+6/R6iQIz9PgbCzaM4ILT4RaTavsJ6ZhcPSXXo5SkW20H
5q9QoemziGCFfumHHFGLOxU9tJM9vThpXdtYQ5tgDsPqz3VfUU5eIbkjtTvwFHpN+NzNXgQK9bCC
RP6yUInQTiG9RNTi2A3un4PjlHsAhHZdcwOzC3xHhEBATbHP9MIY4QMr4V+g+gy4OUgvGEF2Hz+l
rzcvNI6OIsa4OpCS7eXDScWFUQRxy3t6JwcM+3HrbGSsa9V4b6Tw2E4NOJGb2jL389wfqJoSj0j7
im2n9Nbw9IvMq+PaizsgTrclIqhd6l5+GHWE628Qb5g+34T9qiBdIdzpkT6gg17vO6VuL9RLMd80
VN7zLYgArvoqkAkGa/a8Brtlx5t0JMmzIMqr/D+9+TZKtEFYU8oj6sH3QBAJy6wy7OutXJsBFSBH
UbldkbhQOZj9Xqd/oimMMr6/k0JdOiuEKgBGg6rmLy4Caf7e2PhCEjuOk8T0nPAjwjkU1jsId8Vd
1lNVL4lZYex11nHZMOQFlxKzVE47lHYj0nNGsrPrKG8eKgjXlKD2jhA5IKeQPl1INUNHppmTfQaW
uJG35gOguYJxGRZ59hWih7NhltAk7stoNumm77tRnmVnZT63Xf8yd/XCpzrxtYJnhJo3nsUYOCE9
T1Jh6uYqURgNxzC3Jhy6vfHXuxLL2vjGOAkgpahmryifV1h/aoE3d6ecBuDOBNx4v8r7AORyscFO
ga9gIZAKyX2mXfB+ZmdVchXiMhGBccTIWxpgb71uKPjBCO9wPGFOryINfwl2gVRqraZPRr4is830
rQNoG6Qre00DohNEVLlvfr3/fDnpWjkUIgI4IeuRCHjaHcImEZJwU5nTREOB0xa/LWjLvTgy0wLm
yjlhYd3Xs1ENXwJFM42Gv3BAJaNj9BPTLPxUHPWPCdZTRvDe11i0At/73RZxt+p6s2aEsxhxG3U6
JyM0+AdCw18+t9/zkT/0757QMdFHfRYq8ut6SxY9IYGU6HHftiYcxQlOZseu2p9HYgCLvW2RZkBM
ZhHatL9nJVDALancMqBnLUn+dF6dZnYayU3DZjMAgeJuYmm3GjW8e5GhNJWVurRzkcEn+O9IMol/
QXdq8gYRoGLuxq+YdDr6bQ6s9lNdToS8ghT8aLHuvG6AvFzwk0fkCSZLJfqkTc71Xsqbf2cnmPnX
FYGKpt70XU5C8IFkHDyJAObEiN+WrYr25d80TWivyP6D30hY0uns/KBucEaY6zxQkwtvMi41sVkf
FzAReSWtk0iGMRKSlZG9ZHObm9pnEj/qMDU/C8X40kE9Jx3B4/bn3zaWc39Tfv3GeFugGqUJI4j/
Xz0rxLUPVOQKlmIUgUeX7nKDQavz8PvhmPCJo9wifRDwwMD8hdU4b0QvP5Z9v7/9jVucIdd5xPTM
z3dcBqCVdhi3KcbK63u5jHvKhQuvRmK433skezC9rbDfyqptviF1N5rC3KJmW49LFm72hWBbV0l9
QHm0ehfCit89bhSuWev29jaCGrfr+Cr1nElwgHLoQ9w5Yy887uW32nYvT9tn9r4550YhrVl86Cns
Vgi+I3o2eE2d6M70sGxN49L5JZzpIPm4NAiijqPbMX3TWSJI0wSYcTksmtAeIp7Y+UWF9a2GgEO6
rFkGsaokOhKIcfEjpyKexoHVNu8hOETmi8p7DWy0dTr4JGaNKsEu2SZuUnwp9KKWUf+U7LaeVpaI
oFUJQPEPu4frL9UWvqfudJnQTm22qm/QKQaRgSGxJWkdvBUwMBN36jw/2vxjs2p+pK+31mn9WlCH
MviRE0slslxJz6KiigPyAzJmwlugkiEibZipXTHFAeMKeRHXQRs5r2V+ozIoSpvEVoMt74+IHWBW
U0M+3MRRuisGF/ElPHLz6kh5lzEq6JpcYTt+h65XjmbXNpZok+vkHO5ZTVfI1T3myO0cxIcHT2uE
fCGZpdiTKzzh4e13oE50OahN+dqMQefgxb7yrCkIXHP24bkz67hXjOaY0iM7V+JlQritGekhvBOm
7QsFk6O9FL/RbhtgWu0WXSA0cDqzA+Pjc622tpFBgv13h3hjNRxP8PcX9b63NqH79jMbPZQWmH7G
OZ/5JbS7zKCvNidSpSQ4LQhe4FKzqrq83uF1P+WO9oAgZklLt9x1H1FskXN74g6GeiRsNXeM8nFe
xwu+X2KqEOCYYvUNizxIWsy3EdqeOmO3VEBOtjX/g9NLUhx6rxF8/pAiBQZ/eJn4v4+1vc65Br11
5/BbCOvb9EsVQldetc8KjwooPRNZ+gDGHcffR2LUWEr9zWRvPJEP9zzdYZOCeUO8ZZADy+YKz8+y
TOx2ymQGm/h/kSNDpga1Wi2CZTp0X0lTp1Gcnq5GCEQjCWnAooGMZC19SMWdSKHlb511DMXxvyQZ
pYTJZuU5/EGxvhqk1eoDVGv+Du41xPp3eqTZUOoBb9f0Dy+O4bCLGsiFMnW5BPnALDvNINNkRuYs
vJ/8b2PR1yLlldLQTmJ+h+KQ7z6mhvWI2LadndnDJSMGCLI7iPljJvXVQndHfejOfMSYk8iNAbRt
1DmajHUanGfQAt62D7Mi02FDn2bVWA4iyPCSKT9WCJtjNt+72HI8UZ3mKoeNXKIyeLF4qSIdGsv9
xIWsO3MVX4ojt+GXkgNr/GCevPgE0zgLdip4AVpZw/sIgtRjEMnqr8aJh6KHOK1CdGyjmsnsSlgi
kWEw7l97kjZJcpH/mRmjzVNOG6CZcSR+wKXvIyC6YRYwxGzjY351BlC3pHK8JY2RAvqdJDbOZGc/
OpKp/z0F+5q+6GSdKoXfPchbeXH+cGBEAklrCat9TduyXWrICwEEtzFV/0GZT1hVYMadvnlSl/g+
oteATCWPcRefJjYMGtLnt8hwuSLJ4y7k93BgePrs4I+DkixxZLUE4EiKl4K/pl8Z6lRboek+hJO/
85+wzCWelHqpFmAHxAlTqZKipQAqnJxNLKVrmmXhwRAEhJZYNUfp8FXYEraBVZSepvAh7JyRmuEx
jsthzqjgaqz/qV6XlMfewXYRgV4Y8QoJiF1W43HQWfNrK3TWv1AuvuN6uXpCSsRkESQtqyGQTmlM
AR+KsYIvk+RiCrLayAyWHvNsBEty7dsPfxH0AaBlI3mpFE6k5DmG/040kXXejDJ7u/OmgijJUgUP
XApzHR7yDQJSH3SYD9V/LBdDKv6k4JOoK0QYyHgkdk21ub8gdSUJ1nb1xQ864rByNu52ePNoJFn6
YtOoO6I42oVsZKpzpzU07mRXhcY7TVb3e43lHWfObsyn6l79G9LIqtFeNQr0D6sXNmucGPpA7eoe
a4kJHAQJDGZeCX4olLx5AwBLy3pKmgMFF9ECZ3ok44HB/BBjWTNx4z2Jw00VOd/mFqyqPyy5sbIm
BVZKAZv3mFu7IsrMMnGst5mlOcXMh9ug7iEiqMNmy4wCn1P0bhXexMZd1TuPl5auOCvyWv3WbkgZ
ph+p0xgHkmkmxM5KbtFnIpbm2QsawEI0khelRCFlYrLFmy1bOQOLDpIaypgHVR1Gyd71E+HLXKaq
R7cGKysg0Pjtid8b6bwMMSphajtqFyuRYhuQikn2Z2z9DSZBu/TQJr5Gz+r8tOHvvq/SIZSz+lGW
UR1YPR/wiNkSZ38051IqD18gtLAlQ7mmvt3d2orphaTAaoYelu81A8PIMQz5nhYrhOipFO13VcyS
JNV3FXtuc1Z/Bd3V6M4wNUbF0bWLRMwuJXc5v2CdFgpz4r7kIVDPDfjFAgCFl7Km0JiojBwIOCeN
0lBlTDqXaANKnPQFxryvtyO3N/d7GuPnYLFW7G/pULZp6eZuZ87liQJOSppApigV+TkmW3QlDh4a
VIxL51AP4niMY7WN7SacSzOG4oFciB+vSfGjU81HFCALCTU9SWlm9/U9A2pS2MzanyDsU9JB3TCg
c6iqPKRTwO/qrcPBt8EXnJVt940QMVfWT5EGyBBEsPcNNmkYapikXqAuCI9jJJBIiSNDnpDkBtS9
QSBOVU2/XvTrePELaqg9XRYqpMfHCMXDZseV1KWRItk+G5eEaz0HCcjkXEkpLCge30tKaKG7eXlE
4Tjszxc7Zu92MYBQMEEj//QOSUlLddSfeQBEPa/c+TMD2CwlWY9h1uEzIHOS/bgwyt3QXatceFmP
TRGEfAnNeO2uXf5WYxkSe8XJPSGEfwAYNy1wJBVZa86xhTE+gAmQQ0kuwT5ysdnzsH87WyyzqaRv
DxiEKW+090RDEF+RM4l7c1krzJ1C4qBvFfrVJslCksNvimODoX/o3ZGF7T+jr7Ql2ZGl2lgcoMWg
AvHjQClLl6hvdIgDm9o0qeB69+flEfdef2HW52IrCI4+G0WHgu45ltE+qXN4SEfz7Ez7wzzJ0KT9
+/IYJJY+M4QO5md8Sjr5kezqP/USBs/qWGobwkTFqsTrBMXpX4IOeOm7OEYyW9OIC064oxmKM4KF
Gz5ABC+ddFwKUBWgOQY2aF99K/cDkmIuCZVDVujN3hjTh4lqMrC5sRWUjPDXwB43sCbLy6Kk4TrQ
PCiJtZHTyuFDBn8wcK04+jWJfU5PuXpHxiryCHnvhvN006X32E1FYU+t7pnPQ4jNXXBkdsqJa+Ep
76DoCfYc6+RKklh7xNSp04qB397aQRiSC4D0FbQzHwelNczVvr7UYQ6X7NXm+nYgiq8EpG1tBMEe
UuOZ3QzfhCoXfKVvPH0iUsQiBSwQsQJIfB9cSo5g7JvxiqmBKjhEFKUuzDWn/5Zrr0wGDJro8hEJ
XxLwBYmjOzwnQmEPOwW+U4aL2LXk6DbD5YnEVWf4XZN5zfsZJZI/abeIHjNci+xl3+enlg1DroG8
DHrrV23dxiEQsOkJcUnANTOz5dcVWX8Jm3q7mbAQuRczOChMyGjLDGdsv7UxIVpHnLubkQ8JRAx8
pB+i02adgtrgT7TYoIG8AxJLxFh+QcWCw+sTmIGN5YQQcH3j1wZKnizRza5jlXkaounxgwiM1ghy
7xffr5h4J8D9c/L5woOOg9qQm8zDv00ZK6wdNKfFKlmTSO7Sz65jJ0sYs/SHuv2ZSfaKbL9luixL
FpM64rVeU6p8oIi/Zf0M1tM1Ut9L81vSpgklgF7MX2N1wrWQ/TghW/KRjx1pxI+EpGlBWQKeWxjq
oxbGKQkOBKd4EretX5ugPBkEhmgRFGuscQ0XLhlvQurXi80b9t+OpmYmnwj0+9PGPWwA+/A73csb
rOyytXrpEhByS2lBIOE52mNb+NgmQo+A0Xr85IweqVdH+UWFOS2fbUWmDD1qjD8rpJ2RXbmY9tHe
ZSCkPF1M5h26YdpF6nQ0OVJ2q5RRlZzLukNbsz2ZuKk23N9/mYCIxJ8km1bFHu/X7XIlhBHYE+28
ItPnXn4MgkXLfQjtyC26RjDPG7vgRvC3bYuaUEyGJOEfOADHmyKN6dEYZxSGJ6MnSw1pQ9AkQ3/B
9+Re2KCGOggBguG9bmLHBCneDVPTa4+x7/06HMNkB7SKp+xca1ualy3gS1wDu4yxZtF76G4Q8AVX
ekhXGc4zLzUJbBBtO0ehW1FxO+f7Z6LTE2KPQXUnAwViStNtI2mBh/Z/BO85ouKJA7B8JNFNnjba
Iwr4aE7YJx4VDYlfH5WBPEQ2dH8iZGHYB1vokvKDhjZwLYxCWJ0D5BrbNHx/eT3noz1TI8ml1YOu
sPOON91sHaH1MJcjQvMsarEiMWy23dPVxbd6Qe0goiQ24ZxzM/B2JqFG5n8RLqk/XwXZT1Fo8J+9
v0/NPOIXOwF1BPFIi3oHoBMlHJsbfl0rbUuzTLtXurr4RVTqlS9EY+Pjoxb3KNPAjdRoIpslqj8y
0Zi+uvsVS368VH71zv3t7hm8vz+0lJSAVXcg/gITlKcmhHYXLEpAm+xHOmowC6FrJrMMjTcjsnrj
2MDxS+ABQX1Pj5FiV2vcPPqen5oig4SyG/WYqn8iY1ji68fmBNPS9Dtr8VBYB16Hi5sdKfJkhGTW
z/9cipTJpqsVJzyGyzhmM5Axiia6UkqNbuhiCOseCZXucsdXoDygYirwyHgsLd0PfNKThKi7VN11
kQDsp+Y4tpwzL673p6XAwdBaI07ajzzGCnZe9fCa1y0mf3XSVko5NQwr+qO6dYEtS4uuHlVcf2Vi
EOC78BZUptFwq1N8MkBrqlkX7erzNqJ8HN9q6K0UCmm40noKbnw600X0LR4yZ2pkgi7X6CeQE0LR
hfrAbhAxAwIc/JsiHVIoedNrvB6f5LoPUS/iT4pUSkPY26A2qMr5Ax2kizdwcMYECBBhXIgOpmcT
OYszCxnrJ1+HXDUFJZF+AWVBl849Iys1exIgF7wxwf7A73tzkhtwWBi61udgV+ko8TAJvH65+OwL
XPzEoytZXPXIkgdC0SxghhLNFf4ALzZ+TvtIjnSPYB3Kg1I7N3rdpnwokJhTwig1A1u83Za47LND
ZPmJMBkoUXjIctaix6C04/Gw4rKkROE3oJ2To8GXSMPREA2qIvdJaJDB0YwKqPYJv4AjtkT7ea8b
k1Ufsl3kXq05CKm7Q1q7rtHzo0qz+ligGXQE6PikelYQ4NUGnvUN/NP6ww+X6kaDNmYo3JC8jWMd
CZ+JO0vERPqgze02pUEPE4MXpZ3kg6uzs5QBuhfwAckY8fyDnkCGh5qHb34P1zzLBQ6hvaPq39Ke
4YchrzJcyH5B6dwNo+IxEutLlC/1npkwxpiN45iN5fLSe4IcUE/ml8/W+fLVofE585sAKoE8vpY6
uNpLLzCQvFNqw0hf+wxIP+Z3tTGgOIm/bXOmY0ccloxHN8UddhxRc6vnaWGNO72ulfNyij6+VmR2
lnuzC7Nb5TEgLeHXeqBp4nfexnw3/SeUTIeDrXGAyZFilfQYecCWu9eeh1hWuWqzuwFWGeHuxbfC
5M5gv6CrkhJ+OVkLmZbd/yMoGg+izRgf80mWm4coPxNBj746CpyN6zAXBUTAPNbaSYeszZ0Wp03y
IoRkWuK+5tpC4HKrkX4SasLiDNYPu/uOJ4knh5qHD1aY9KTGI2+0ENIv1U8rKjOUEH9dxBh1pUGT
SGGdiL4yzUnd6L7dE17jj5dOiPiVbDbwEbDp2qi4ST3u+EKDzfgXNeULZivi2QMQSy4Stx2rLvYi
bI/wDG9zgfqjMc/mWGT3wa4csgm6qtRFNoq2h3JGHgzie9TBkeMgoVrr/JALvttUbSDiHM/Rewkp
25pRe8Mbfld7ebcMAPYTNEPv9lYqCpG+lS0OXzG+5cM5UgtCS6WCNe4Um9LC/ns0q9Ovn/yhJdw/
yLBKEQdMdcWUsO0iqnZALRmiJDlRtCVVJruuGO4wt2yJUisvNWfG96RkNvpxeFOPbXK8gGJ9GJ2N
/7y1fnAxQ9zES2UZ9PUvJ6nex3ckXNeJgqUBibtsvprpgOoHGo6lB/lA+/DcHirPIHv1VCGNj72x
TBcsL7hhQ/3TNJayIQBycVIaH0msKjropq+6JYuJ+BavCxSP/7GrUCVQKucrup8daP0hFfiU/WFz
+SXeXXCmlF0k+E4faR0P+41qQgDQZL4MeyQnlzK1dXW1mCimKtyDu3Z9dn4d+nZ1u2lqc4uOZX0I
UDUWSuKN8b5qtaeE9niyYh4l6g5noePWMp04VI/B1PE5yGpU3+Zpw8Tyw19ZpyVtb3JZrPYTeeCE
f9rl+n8Uv9xnZxwANhbJqC6/sXS7XMWaO2jNi5dWuAdyF+eE7XixRUa61I72gjDx83Mw1umyADvO
//Xkk341jJUeVsIVQvcwVPJNHIyAedPkY/ZLUdG3RoTSl6G+kvHUaBVuf2Qw4B92FDLuW104oEvn
Lvy5niirgvmYxfzs6NMfm9QxVAN6hVkMTRuudRUcJti3/sxswyy/so/KautzTIyTcjyc0LIbNNMM
Dm1ARWvR1Mxfy8CzYmNC5mb+7gG1MDEO14LfLUQAQ/x7ULpSLMpNKLT5itnW8KQ2EfBRBVPFR3Xu
6kITyHCAPXmnALIESnycxIkKYTjIXeiQfjAlJmgds/myXUsC6jCjrr22Uv2TgSxYxilMiK1YxHWK
RMEsortuTpYf/Mo9OJAyWivoMuwS9kLWnvAdCSMdjS04HfGIH1oBJ1avAfNQzh7YYfWmkBa09zeA
4mmlEfFMoURuLl5MPf4LRIqmXvbEewqYYGI4dVDBQNoq9LILMdRpiPi4pRcgwIzUTfI0pszLLIq9
Custu794q/jrCr9bDkiYEZJZH/49xyAyLgqKZOGproocYy/d622AwV91djI86PN0LIYnpgKRrCyR
EsI8I/7f1llHKhzAyKbEAIlb81BKhtGglnGt3jyG7bzQflkiD4eianATw8S04jUOZmgucnmzi4PS
zYQwsaikaz+7JSnYQy/9q01rbCYePuZznB/0PMvWxDfAhRdS2ujAo9OJuBqExUfug40nPff+FzOE
7LOh5qdAhKt17lSOlllz9vTbBctFD4qxZ7gZ+AeATIz/NozpVYuDo+YSeAH3+zeE2LjT809CkZDa
PyUfDbERDDOQ89G6kbmp45rT2Kut4EJhecB6fzf3DqTAFfUHwzYGPIILcoFw2+W/uqttOEH6Gtt+
uNBmlv6i9HRPjX7P9+kLZi4kIfy740Z4yZZhQsIeY5LtT002iuzAHOXTAfKCvNBG2FDPihoc9quM
SsFOBilT9lZs8Kl6/j+a5D7cPbZOvj3N9veEkp+Uhwogt2mVJqBe638wglcObgnoGXqvEpKDXadB
bCFTvwto+aI6bo9s8bRXj6dbPGVbWD+XW3A0qwoFs9SHZ9K2oKYPyC+ode1Jtfx6+yvs3w4LC+7Z
f8pU37ijITu4HL0Lugk7IUobnAMd/bxMfp/gkKWKzIBxi0IwtbIei0c5Azdc9J50EPmqcx1mzYng
/QddOE81wdeWOePdoFWbKmz5Foi0uMYtS6hivmc8gatCW4R/S6kyw/LKQOW6kGj9cm1Rr50vNZSp
foGmtihVvvsFDODAhYAbXQBalNt7a7ajsCAeiqozGpq3Ut4vrN4lfo2koOmPlR3dlPuoDdd8ymEv
6uxRoT7NN1vb+12fZHTu19jVx+VWfn2xx3bY0UWrKADeUVdwo4XTOoMZd3oW4GmVAscXgo24wIu3
MfKeawQJ+hIDZYRd/YSIqW4qpRtikqQXGStKqXxwp5av2/nGZfte+A90mU/LPDrCd5D0Nwq7VMPf
UYnKmNZqgDMdgEEHgw0JrRRo3fsATAoiVfzbH596/UpQUBfjWHrZlEQC6Fdp/eSAmIi+JKWPA7En
HQ85ALyGHE5eWKkJreeaJN9eQqGpE7ONpOAWLBPqteEb8oQjlvtk4/3NY4HUY4B/XIaFQrnmzZHY
9kQMwjDlatUs/gNj8/u0Nckrz8HSn0JIRpyWTw9dGkUc+Ad0cv9oRxbJF8rttTp/UWib7/KrE/bB
0bUKeNPEWMR2WY15l0E3SYt1qT+bKrDBA/u2IA39Dul8ecCc6w7/y8J4u7SHFoBvfgTOrQ0BlCoK
3mJQMe+ov9IeZKRftTWLWOv6uMvUfz7z4aULYNYPpST3q68QR6igba2zBEoI9Ak/Pgo56+5xPTk1
vwjMAFxb03DWSF/5aqQMNtRB18d4BFg092qdqqlgveByf72TXBVUYrxkyP21KocUBkwcB9tHy0On
u3OrNAtUqdEPP9n/5iEwKtu4b6YljtAXRcbNZdWFAsINdUxgS5YC69QdekQ1nhlK/z6JHNI8PSig
Gdj1K0DlFaP35j2J1TNMWHgMz+HuBAV9xdoQgGjf4MgfVnHyEIi28vY9JgJEw3bbV2he1ycQjKoA
Icu1iPUYUn30HJqWd3Ffb+PVPZctAp4FchKYCMW7b1bNxonZuYTNIbPVn2CwNVzS0qAmnw4Irh2K
3iheBLory3zeIZPLxngTp2Pz2b5AupOJMSB0AnhE8eJ3rRbZnQhTuCVzR/7OJLDLPLSPOF+MdpTY
w/HOplbuNxw8xfMrb7wHyugXu6oM3FfTo1U3JYvyjhx7ZnU1wyx3Hz/TYSfh4fQPhgHeMQfkt0Cx
ngY+OZMPeuuuh44mtlwdWhkxfO+7jHGMevYLNa/80owRRiEms5NzyQlIM/L3dEuxi63mPdKVxi5h
uHUAVm4ngW9LQsAyNL5tWLEY4CxX/WT5CROVIG180eVDndp4WjyMYSzufdsCPP+m7RrEMMOKnSnl
WbmpIGYdHD3uYMS3kuy70G/7IIz/TDkKQTlS7HWxDDxjI8d3w0FdctipmSvtKe2vwc4T4oppuqp8
vuI+d8+Pb2rK7o12VrIMELtlk4WrmHvOkKFswqfY5t/O1E9xvs4efhoTOGs2RagLWspP3r53HxNT
9dzEOrjGFdUc6iIpGrHVb81mShODDCbKp4WPCXscM2PHzbou4Le3LKxG3Y1cYIXLMhswRtufCHik
Ahj3NfDLimExGdDAWWvHeaWZescv+brnDwfd9TeYDLRFt4GWzyQr5fmlyTsNguPx8x86SW0JRv6i
s/Vqelm2wbHMyohSfjsFqi9Z3oRrBqIrs2tVZltCbDHeP3GvVZrxiZoLeGMKV+K/0vGnjjhljWqJ
cqc9ai8HywF/v5bVk+2CeydpMIJY5lOLXYRGwCYMAQzziM3A+KeV1FI9txRmqbyb7WJjuT24woSg
y93+BvY7bln9ZT2tVOIXpRCjXJdwzRgmYzsrzSvhkOCTsHht4YbHrvDl7cUGnuPgQdhXc5oFbIYA
KP1WZNytfeECTZjk/By8w7gaH8uA+qIc/YqzFUBGBFYbY53a5Q5lo1bdgW2mMQjScoQNPTYpXIx0
+3CBbTdI+WQ6HC03d2aXI89Rnf6WyJcWMbdDtRZJszmihsXbAKifyTNDb/OfDJHbd1FNtLVr/dDD
1XXHo3LlXKBLc5NOHMKcmop+If4RK0eyTmvcEVCeylY8XTXt5TB0D1gJBWQ5RXjzNJeqFnl4Cq9v
sWndpzIWhEmrrIrijrN+UuEbXLh1Q2UzBWThp+MHkzqsgs2WkZImnn5UbVnjcUcd6x1BWhbbdOeb
PHQ2TSqHX5SavpcgZ95rU3/P1+EeBfxeifmehj/m3Ha/rGxVEskte6qes6uh0MM7HCWmkwodYr1Q
AiQc8Qcv0gzD0ZmlhcU0fCd8jzSv5KhaqCPrjWHz7Dtd+Vmy2myDRNGEq97Hpgg7ZwXUpoNhJReZ
NdqEMBNNSf/5eCYbyqM0LJsQsovoW6+O3si1VA1OWl9vGo99svDscwg70eBRtUl7SY56TrMpd2cl
FILvCUsDJFtQPxsrE6Sdl1uCLyX1/YUb3UWPv0HoRVNYKYOdPDz1NY1qZ9DXVCAyKTest7hx4e2k
WGF2MLsclB4aFInPflkQOiO6e5iykUkuJffujt459kXH8bO4MC5I5AZ7p86IJuxzwg/AGANqQdw+
O9bKWlv1I+mv5FGSAZrEuerocMterP85ChU2x/AYupDhzMTplD+JQMCbWK+jgAD8ZzwXuahB6ML5
8RsCLxTX+SScUDRP+KCrBnL4dZSu2in0bGH1tL/Npga9LPSPolbwg6J/3Agzf2WNNnjjXSvz/iqa
HGxAEF4SpLLBSXPmjDC8tKUqPMuN49TGTXIN6Ghq0kCDH3KfGfFK+yCAkuvk4AYHCv9LrVhEmDFs
aPk1O/kuftSFdNl/Rfi8ja/lTh5LuKYHxlkFWfH75hOA+cQZcaqDKtTqLHJHsWqdsa8gjwJwWZKR
bCnx3b6sJfF17rH7Du8+8o0OrCLqbxbdKKRT1pALxFICq8rXr9AExXKh+Gx4ll5e3qKiQYyvBYfI
03iMMkRnbZ4VFKxUBuPsrz+isTRBKAEmTvNpexEFYTbuaLIxKwnuy9HXRVrvHvarX7Fvbn2VGlKr
Lk5aezLMQC/oR32Eb5Aq5T204Q/6b9i5fFy/11zeKSHsKznx3dI9ctxC+Lwi/0o/rE0UXmvBxvFO
rKUdrcgUOAMVyzTh7q5D9Ii9441ltnG5i9ioyjzq0dw7vk+BJyk4vkZVOJGbf5LJgPBhTH3WUn9J
nY+6JYJRfdUn2B2VQhg09cpIGh8gZ5fs5ltTzcBv0Vj3PvfXAyVGPqmnylWtoMsCDnTyMes5aGSg
V88+rcDRqhTVP+U8mgDS7suQsywStUxWgjJhKheUi+58ITe0GvkAHfIPDDlAh4AuwunclydRxrau
kICwz/sW3RiTetch+FXPgARXOude1A/+9UqiI9H0FqOVQgIyiGw0ojNxXxLKFNhpJaPBKQqSNcJS
aOjWyartgBbPb9HYbiDK4ZbuB7d4Y/vxTNS9ehI2vW4YKOzN/8oEE2ZLld909s+r02SxempkQBJ1
UHPm/kvldaNLxuegUqB0rt15OqU8Dvh57Fz41ga26mfLzv6cNjEvHGUd08w7n6iKF2KIvHGfx4wv
d4VxpFtggB7Mlax1a1qaLRmyHz4GJqRawdkumAgY0/tC6vrRgvfhEnMYBfeIO6B3SrRUwUVAHqNe
nipzBD0j18q2ABPkY26x8GlqdE6u3L8coBseTNfhrfkPVWtaOGt20QabLZjCHUapzLvAZi78KBfB
0bpsi8Lmiq/Jn6Xn7oh67XhLCuJRlqA9VK9WKR9y87Ve+BxaAY69asHpal7g7iDEdkYO5hMmTPoW
tS22btv3/oY8brHdStZzhxmsG/Nqtn60OARpM9kt62TEqWhogJBjmND0bvwQpJ8j65OhaQFggIKg
Rg0J0NSJ1VwMRiEaMZDEHXXRv32pYyq6KXM2TCyuWR99BbvCxHIuc3cxZpwMvsGEW03gjld63O3O
P9URyZm8Oy+JTkdzuh0jSN3FNPO5JmCPy9YGhy6SeSlDXrOQduIPt9pM1w2HNmlXzqwFl5+SuhyX
FGyJ+l5gUvqTxEfQ1UypBmTjPn/q7gKk4xYINGFuaUNzrXH17PlcDhqD8IA5iuXFPxhszmsum0Yn
DgdzjZ8J10lEKNdtsghwDmUA2fzMt9iCvOTzNhc4q6m6vxKllsmL7SDsgMqDCUiC9NQ+Gn69QxZs
EpRbtW9oWHbaqrZsfHRsSFjxa6CT5gmeVCEJnukkhbTC3MEDdyTK39iIxoC9k0uRPPM58+R79tA9
JiZWl+QNA/e/QpuDWAEhr37wK+zh/mrNqHu3uDUtfUgtiGG7iQqZLar72f8ZDdHDv98HqQv2HQi/
oZtSgU7GR1Z8Fb4FbwOTNssxdDbDOEHttGIP6OHhGB9Mjrok0/xg3oXg7AxuCE+FMTLvi+lXLsjo
dBDeoqAnt9rlT3X6j4a5p3hXn0QZPx/tOHxletYS85ccx/oaYu6+Rb3BzjJFO1SiAi3p/LCzw+dB
ku7BO6Eyqmg5XacqU+4IJxtMiR4BExGEnBVJw5KQQ682nxaNy3F7EBQ5XLiB9S46fH7NeWHmKGoN
N1rMBEYlZb/64cXIHh/JVWBgzcON0HCdnCVGAK6GQTETL8tTZbcoGTqtBb4bnKrRQezW/VRIeU2n
8xbV/W8yqZCLsV3xRuWCj5UzpK2phkYqXZly7giaw/Z9wYItuERsSSSUe8z98rgH9SVGtvKrXnkQ
gcQ+97j9dCdLJJyoy8bPPDf0QKGJyFI1v9COHab+ER2tSj3T8mBjZ8UhDM4H6/fzvJaqhMk2JAHZ
gs9+r+/z12zzBaYqU895ovfa5QjqglyWylhMdbldBaLRphd3sX7+dkhM5QrmkVV2zgHRIHWUnNs2
fq9aTcMM6wVCuFfX8NTDD5IFeIFBEbqwIblfK2oW1/XFx03NOdR7N1lqrtFHQJ0OQBCgABY/PZ0T
zefq/wJR9VyBeTSdjcEGei4SjEUQ/86QRRidsL2x2vYPOk7eYEps9C00k4U5+lQTeKdcGBZno6bC
LwdNHiuvDxxN1n6IGo4lYIvv2s5fSQnqxhgdT+pMpjMHhJT+vvH5guBzFDdiDf117q0UezReNP/E
2jNXfavmnaKf4mFSVXiyJDtfxeBvuJ12zVY2xkoNcVT7LJ/TpqcR3vMQk5sOYwggNnLu42Drclu9
jT9M7IOJeV3j0Ca/wlPOYR6EDlxxeQTanThpRWa6NuK8wVraSsrDNFpwlzag6dJbuc4lL7IK3MWD
9ST4WRPFFS8Ui9DFlvSvsKSUI82qdjbwKLqRMgg5zbyKJX8Y0giwdnq+jCkIknuYb4cZlRoPg/qd
iK7QpIvWYCtCW28DimIFQr6Z8liyH86wFRyygGA0qJFrCX3ZsYI8jS9lMPMqBzckF5Z+EvVGDnJe
3sNr1N96v++BcFAr2VgW79Z9j1z7a9PbF1HeOmQdfmJWjbZ74RhxQs3g5txx0t1NIXFkkgH+Kc2Z
IYueCQd3CJ3qe+iZo0xbhlrrTvekqEvtyxPfEfP//Budo2jjEUzWudLvH/9+qltYdibSlEoml5dO
3XS01wbfkBODwce2QHqcwR7ZzmPwB/YicJPt5FO5C8iTiikXs45mTF0YnfNRMDsyqhkc7PgMps4h
D9NJEROnmB/69ipIIhUBudOrs1P9H/gnP1mNgj4x6sp9FYzyLryToRtqazlIau12VgU+jWK4AWn/
TSBYVKL5LbCmL7vAFPffS4D2oB3xLQ7oUx+l2MDWz7w6q1zNKqj5l1kRFXO0RVlT0aMSkWsros0Y
sGy2umusctYfe9FDpGCqu4KWzOvcGhGSaIDaZayWESmd6aC6KOi4809BqPFcclV+7rQmSIgNQM+h
DAZH79jPQ41rV/Jv5k9eYJplM2QGEv0c6tPMJxZxfjzGd+zcUAb6j7SphPf6ptWJAwbM1xXNr98o
4gN/MCetvudvK24Lu9KZDRTQH5KluUtZzAX7o9fpdIRrtiFMxlkhnEcjmczyrmB8R54zMPCy0w2c
uCeyHDIr0/+iKDKi3XGISjsFn3ejcQ5AkCxLtP8VaVFhFhyDGkijgfUtjClfWiZlxng4l7TqOqQc
0djc95bajkKCs49kAn3mqs9CMDK2o1SnXOxyPFwshsqZysJTyld3EIkcunqzEOwrqkgKd5g6igp3
hlITBzVWkesQoi1fksIvIpFdKgjQ5SA13wdysOA1TDZk1QALlVvb8HAiqjv3WfpoNshFaQRcyqVP
xW8IMeislYXMLANzLrtKQDzAdGYOC6cSWE9CS3Bln2qeMC8+UUIwFWOey8rV5rfiGKRefLSGqekb
AwwD9BuoXNDHrQosdJAlFRMPljnl3CUtp9A80U1873qNTi3ZSwjneRTcGWplf0OAqhMExQ4EEOT9
lZVFaGrXZyja84VnNY2rpVYV03pmTZtotSaeiDcNatRHLyFn38SYGhVm0bmpqURWZp6Sn6zuNEHa
JvMxygORs21z+K7IZ15WdR+sQy2N9WEdmoa80FpunFfbAFSTIGL28YZUBapOQ1ise3MFezbV2dDA
xIr1mICt9OsceogsRsBCZSEe6U7WuOdp46ocgWQctSCaSATCaj56Pz0St0rYqC0D2Ke7oHO4mwYm
1RFp5Ud/cp2Jv89Y2r/DvaJxZ6w36wq7+fiqPIS6o6WonyNRtAu8lT//buEHzugtdQ1KABSIq9/B
GRkPRclgHattP4gxIRhVH9DcVxwVka/PlpMcs9QqarWF8baigSoZsQkryRJ0FnfoFnzrQA55GubX
xOq+qrrHuHAcN45ol+izyWVPfvMQSpMdnTbMW4bBuAjORGmaZafQ9tt6E4MXVKgeQhxg49S6uIDS
yF7bpG30/gWjKFL6pZw7tsMqRyGziG20NotyiOi8CyBE9FO5AdX2z2D3Kvvrg6OOK19lG3eK/V1l
NiPL/C9sSZBy1Q2ZUUXhm94fJMfvMBXPTBPISnVuamrkZLGSiXTdDpdUFb9sF9ejs8z1Q0F76KdI
bqJ7EbfsQCHoa/IRY+yjAp5ajI6oR6AVCBsRfykjUT6LzYv9NkjId2MJCeR6XyjOHI+afgX0L/JU
iRV+CGHNKfv8IeteC0sg4ODy1Ptc9TfFEDR0MrzJpvlkYgbROd5a2bAk5KzOwRDtbGNkm6OVgk1N
qzUvxgXWvHwuc6NWs/ljfHe7sEzIVTx5e+FwQO3miTSMaxPmWo0/DkBnF3YtnKDQC/AGGFyEe8aW
XocxWPVaEfJHgLEkPrwEwc1pjXPsNZiisjCDAx2/Xd6S96O+LduUXO8xjnfWrVA0BSqwtbwoJfLD
+42IZO8DToG8yGsavAKnA8fIo4VdlStBer9tIvH+8jM7/RVDAi44ewkPJoLiyK9PDUXwWBd5Cjh7
fCVxTZwKvkGrWSGuShc5xYYg+yROAUJ/UEKFjLGMJe4LPNE6xim/fEK+jtQ01S2tgwEKg31CH+EC
EHFnWfsneqIj5WLJPLG6COuUHqkbTY069rGLt2iAtQDpcTZf8tlO0jKWvkvgCQ0ytYb1TSjsW0cv
MuPsxEEQm1CYycdhXpUz9dhEIGNKi9bI+ofHL3Lyh/eFqCOFD4znnmyvVHlLokysnqMU35W5ay55
xem4jSA2f7PJGgctbGZOszmVbGu77boyjTYw/Nhs6OFeNSIu/xnoXATmxms9IdAytvIAv56quiDJ
zC8r0xwmxfsqFneEzFMxSs+rJ37kMm/l8Pwi50siwvtPDH/oIDPPcJ4aVCnPJWfgH+O92R+P2snp
bSOBTAYE3TezhtIRcXmCFbTg3uzKCSW1blQK514WcDb9B/zswtx28GvVROWt1m5W5qn+6s8C2XOE
gy1Nk6VU8+aCZavBfu0LciAU8cPlqvQmFx7T3t94m0TOx/h4EhI1uLWZB+se37WBzQHBmmi1oeSW
Hd0dCzb/lCYMM5IL4uN/RxIL+6e2zUjF1nlmbZyFiXUuF0E6z+4KZ7c2YNyoBTcqInOo9wsticsz
0hW4hUNJ2oO0T9QEKd2kBvUZ9pOE7siVj9DSs1KTWNTZeWHME+NGheVRtoSpsYRqba+g9sPZVfxg
d6Qs32tZ57Q8sIc2bUETyVB36PIUvrFVhSxcGGMYSf407NTyTrZv1gTGyDn9ybPSqYV9F13UkTrA
O3nQ/tjD5xHk/Gx7WQ/GwEg4hV+mbBbkjoWugiOHni8vXGE28Z69dWgdnAyYY2ZkqYVaLu+d7ZNe
6qy2Hq/hkgCoWNeVg8w8aaW2+FbNwAHiKm3DanhgdTZyhSKkjuTgjIAkFesFTErS/lK6EUSjANbs
UsOb7XEQ+l7McNqgt5QK+dPKJJFDbsI9AVtiIbXLGSKxEm1munD79DneAbvsa1hqp4V4ucFMhuyL
OXJFhcF2vGKDy/no1VPrS0cLjvnBL9FLQbzC/6FWTQvKEBgAfsJmG//X3nk8tAZ+ah/JBqfFHP0M
bYMCPRlpsOWR6RKsHm+7Kl+HJPgDfMpqFlASlGOtsOB0dECv9C3f72maXXQ57RZgOxBSBt8iVsif
Bm3xqh259o7FVLlB4/sNFnNFZmSph97X7ax6FL42bdu2N7zSOGhJMBEeyRILcic5QPMuI7zYfaZF
j7vRmfl6/6ijDyVl69kqWJhjh4bBx2Z7zssMV1NBaJId80Mp4/dF5MYR1bHcdU95gDz7Edx2NAIP
w1zzIuvtzp183ZIEvIjknGjgiidqJLpYJtNp2DvKddH78psPKMQT4ruFyla1eGUHTOlpczpJAlcF
rXuHyKyMIt8k1ae4xHDs7WiqMD3PZdkq/0mIvFAD0CynYRSU9tr9fHzw9zt+BrndOYFb/eaI4+rp
c0T44NgA3b4bKebBP4gLFiV7WhYhp2SJ1J5Bj+q8mHCA7ecXxYUwopsDDvktUFDVnHaBONSXVluC
27lqCGIfPK+2vOU+cLJYcDHSMAhqWqm9A9ht/5FY4XLjKHDtWSu2862+uDcN+PSu0UsEBVmkcUBN
W3qAAibNDy+G4OB2YbSatVccX+GVUlzKWk37f78hajGPA0+VYikffzah42Sb4pAk59FU9WnG/hSg
Oq/4etbFEt5VJQ2h8ZDN/WY4YtVAPnd6CYIxPMv1XCTiNECIBoQ8QxxgHtZviQLOzQGTg+CFUuBD
JLtGdNnqaiB26h+2IIzfkYkUr2/VeUK0hzW0krr6oTgdL9JUxW/I5nqJpWbEf57CXx/FtJhpfmJu
Mzo+ag5o/VjdBrG3LlqfTXsVfLqRt2w9koKUL7aZup1xCvRuDWUqKN0olcTjQeYh3L+aBTghakN1
qvfFW95RyuKjpV1vshrUnRqFoRucfwroIKvK5B1ehOqJC0CbF552jSofnmWbEnbI/VjTno61Ucsa
njghZ8616rHBBiLyV2Mc+IKfdDUh/TxGBdHT8sRRRkp1Aw0UQOvW6QlxbtCjQFrx9rA/jLWI2jIf
FO3jOVz2wRncjrAfh1ujfqIDKP4/fHxvVV9Q3wDc5j3zhnZTrjz9rbt0kell+0b6pBMQkXqvEvHy
vt3PIMcj7vggHOQMH4NJhmecHHhQuyn4mEZlIYdM2UiFjImBPzbPjZ/yLjRTOTI/H2Ep05Hai8k2
GIs0CkmERDH6FdkPZdYnZ9rnf18R+dBP8Od5a4457ZUbHkY7MjeCnMAVZqPSgVGmT30nIx1AzuU4
g6LfosD/ZIqHo9jJEZgC0NYEf7WnPVkxXoAlDYXtNfGE1xivnIktFzpmOn9e0bu/udUZUI+c2ARR
zxPMItxnQj2fVVmNDgfkUwrYNS4idcwMZLZjH7+WiTnv4I/R+z0S9a4zY2EiQdT7OwnybDmnsn60
7vq9HM3cIC8D3NUrZcswPGY2CtLHgyRfIWgAhg9Dugd1+HtvCn4IrdzBdtPNYJgKc51i0m6lXywq
mTu0N3fhQcV63X/jurp4YEW1E025EFFhQzbL3SyDkA7nBSBeLYAD1h4zWkjUpHfC/Pwi03ElNPjO
1cmJ9ZLXcP15q+eKqGPb7dqHDc9BEFeeEky3vqYiCdAYR62KIZK++/TWTUn0eBSUOJX7EDllJyPl
7W4mhl2S+yHCo+5I9agE/maoBNPhKOLD+HbvmTVjvU17VQY55lsdEfhsUBlZoIoKq0PKfSznQ2rX
6QzvTdYO6VNT77xMp7lAaoDsYtNybGJ1MuFg7iJ4V/qnuSrDu9SGVFRRps+yLc53BcAYmF6cc5F3
cRQVMDeiuTK8flt1eNZol63W85zTdzd88P3ji1XH0SK5gTTWUBxKmeG4QkTWbvTtyCMd0nZrGk56
/gWF6JFBdBQ3HHFkdxfMvs6d6oAf+OkBdyXbkG6gmmEmxx43iBXHhgIaFDNwRxU5b4Amb7I8pfOi
C648YhqqDpCdWzojzgE3Oxce8ACj1q4GpyjWdYVdqhOX+pZH+RoUL7jIg5vL9k9O7MGUtYvtUmWk
oFcxhDV434e3gwV4SWcZYtIPS0jhcHp7aWCTG6krbcZ+FSSxIGvkvd5eh+mMZU55FDob4n5aUXHy
QS/w1HbKyqxIuNPe+S39bjrc8lght6S9YsSh4Jpea1cTRKvsuQfqIyG9DRglKLriZKvPg76/OzTI
/U9TM5XG4YuW65LVkgo5FsJ2DqSyFqUzPeko0PKjYnm6OYICaTUeY2N/8diLATSGjL4mTN5POv3F
tG010bGGPL21jlkbEmEvsGPConwUt0Ggf2fNf6kYDkvoGPJhBwp4wOMHz2iKr89Da/UdgQzaL6Ou
LbZVf4GJEA1rWNX1y79J5vHy/Wh/f5mLypkgTCLH5IJZRYgYus/0YtsDEEsluODG61k6+9EMzCRD
pItAujtVf5jPpLLGtKQTfAtC28Kzz9KWbLDTK/PeDNm3gXwxEL8EYuGi9ND9Qgpefxm0lTxGzpIJ
GxC6w/7rdvaj9SUy41/DXAHEd3WrEfRI2S+slwkI+q0gAQEm4VCi6SMjdZk9Givc0UeLQJEHcjDU
U2EcUMeGQMTa3oSptZtt4ExBTxLPZ6mUXPXTifJQMjlxijrYSXg2xew+Fc5Zp9McuUB9e17gIYa2
dEiRSk4hNDY1ecLjy95scpkT8tIbwIgT7Dww5lcTeU9SqPl7qHFz9M7qih7BkbzXw4rLFHLujfDr
He+Yf9JL2899VLdL1pSz8Rc5cw02WY1lOVWYgSzOi+uZeu7zrHPidMgySYWyQJ9V1aSq1Pcq+V6H
TcR5IrBJo1l9KVpzj38h9jIRivA72mKhI6j4hWAzIRx8cKj5CwV0XG2lfbCzn0HPPTolC5WLHrcY
lgtU3rUvM7oqLr2rcrlXyFFLTgoUQ/57PRs9cFkF8i8RO8hjZElqiEDZzF8YClbWNBkGBcECS9zn
VnmWD5JM5dKXf81MnisxjvwrtA0y9qScLIZkv22OgLGB1JB3HquzhKUhoMJFUasvGGSafAG8hhj4
D1pjeevWzTD8wYeaLFNxbOfm+FLcWbifqQldFkP39QSCTbHdUkOHD2+kzqU7/grielXgdE/rgJqi
kDNNEllJJo+t1zHNMXuGVWSF47AFrVJfn8Fz2tacIVp0KxUXb/6tJxL0liizfiqL6NhcBlma0rvZ
ZduxWupsRYIHljnsB3yK9z0OVP499HJSco8G3BdfyaDGuBtTtC026r+dAhj2ao9cUyzXM6ZeY++9
jeZUU/+92yXz+7GogtSuoKYyhhrOsttefUFaM1otlHyeAck9lyskQwlNjAkeScz+OtWBTcMaLQQc
Sfv1tOKtUhmwx2VodamqO2Z/gzSdzg7yYgtNBrUFvdXOKkyZFylEWOuDQVIzjqUvjg9b7BFeBUJa
4tXzHudZp7edEaLf8cI/d1GnzKRWnivpaHHwRdpF1uTQ3uGTtwkX0Di+nSA5e10+G9cYKzpspsz4
cVWL0uq4W9ixLMV41ixwYdLHDdwffLginmHEXzm3X3W9Kb7pDJESVMw5zS5KqKmW9e9xI9z8XfvA
nMMTSEx+o5s0e9dTJfrfIjVOWjDWezwjvJFLz7YypMYVAAK5ruUf+yiBUXSlypk8yn9NLcWbN4F1
7O+5l2hm+ZHo4UFE7VPUFMyDf12kqi4qXs27/VlPKcWa0qZwu/1Cvm+9gc/EB3brLb9mlPOErKcu
ugKSBpZCbA0HKBQIWCKb9Ssu68aCtrG9xJ5vlD1VplZPMkCzfQk5UpjaOh6PApTaZN7fGjtbQIVn
Q/MxW+rPg8CRYVzeE+/FQbgqVVlAbilKshGghPaXtTLvrkT2OGAgsCkCYDSdl5HGVhOf0MzXtieJ
+XiXRy6r/0ZbVq5Fifa3E3Pvl44wz7f+BxFdm37Bf6bRBfg+RUrqe16HOeELSQ32l4IODTfPlVQC
iqKznfwuhPC0+iwD7R1x/MazwVz/BCc+2ZJ31+feVNZLGYK8Uv7NZPdNlJHT+cwkniB2PztSTRsi
LB9Fw9oXwAWliZJhnJc+zhlX9t6EoqMB+f4kxBJgYUugQkSX5LTghrQBJdOf5ZIkl+goLYFLx7sW
efgKxYclOSfm/gtg4vvPXWad7FEHAu4yaCLNk/hT+lYX/WccQ5uhFW4/dc40KF9sEunVioO4tkwp
zENoIzy56AEBspGj3RIiI0nqOJd/hm+6GEXO+uH5VVLU4xHwYSubxj2oJ3DSVzGGnPjc1j0T6eCm
dO5F+ahZvEoKVXLV78/WqkLJtlGeFsFuAGObCfxhrw9gYDOWShHZLFYymjW7pKkK3KqNIUQYkhB5
Lp3YtOwoKgjJmQ6td9tsx6WFi7k8G1vCyvgva+NtEC3K+4vX3LS6Yc3JgacGUK1arM5AbbbXw833
GXpVzAUi+PqlzpmmC7jigqObfHu1qx55qggshMYsPatTJqp8zVEi1OPvDp223YZrAM6ieRV2GiiC
2lqICpDh0LNYS0C4QVK3QQLhfpWKnMEeOdksyhjZY+j3zfGkiCVxG4MtaaTlWhOuCqzTgKFQNVob
whzz2dHHspE0I8T4C+HAOyDvXWxDBYUklsYIbO8a5mCekAWiHhJWvtCeuRECtvreLAcEbJ6U/MRX
p7LHKz/UtKjxfT9pqmxMs5iHkkhHRG4dPNB3aSjWwR8DtXoSLw/omWnGQVPbJcX3oOoVb08rltYc
NU9EfT3W7xnv2zpfDVlQlLRVEJ2qfJYP6K9Zg6Y0DHipWYTAMVyHFlc0/weEPCfmHiH0rfDsMffY
5sbrKK2ui+PF5eWJSflQPyxV6PBJAR+0FPPXJjMt77vL159dItiJdYfhBgrd62H1T0PIN4WaiDbm
ZWE207hS8vZ/Q74ETPLTdSm0lWjTGGXJ0GIDGk0/PwIifWQSRC2rxMmF28SH0+3EZgG0Jx0f9B95
wgCODitLlr64iFQL1GAst5H5E4CkWmpMvXbZf4suWifKJFYXL1mvdDBamfXLKWSQFmboyR4i70x1
vraH5LGPgEf7ZNXAvROG1qwAvjDXD1qI0qA9He1p+K2E50GDWgI4Df450D1VoxLpASFb0EPm2Tut
Me9K1P9OMGF5PjH8ZqCVtbXnws79HdMP1BFBe5XW+VVVbwCPRbhq33bBKrXcDLtfl9PRRTXbsVs9
ei6vxb/Vo0ei+ZeKmiQIIwswyUyusVQDi9FgtdsVaC/4u5/ELb8ISyphrYF+UgNdqPKqIADzXlU4
T0Uyn5LSqJvH2trzpB5PyYzFAWxKSRgDTZk+AAXYY92P//vp8grYvkkIc8IG9N03U/jSyDfefo3k
Of6t6yLXlmnEjFf/tAvplj59YN+ZbkE7IAjTwwibDEX+CG3fYYrxekmoAmNn4iO02+Ezdfiag7SK
pzAK+acMdAksWntmU/QCcJ7jbuDE0hLXfs9rrN+a4nwwjZ8TZGLhQ9qPAV3B5nkE1vrazEcT7LeH
PgjyQy037Qz2ZBnA1G344mSXGhUef/X4Ga75CD6b2EawPrksK8OT2RCIL5BavhnkmgO0DTqiPV6/
Ea4+xM9Lw8k8hqG+CpSESJaaRJrDgbDFcekqsfdaeI0KEa6/2LIOh8YTqkVH9SL3pb6jgxH4nGLK
iTIbvXYhJiY77slu3e+cyJwJMlG66jqOkkX00WQ84AdBQ2Y4RvcXBnkUnL5XVGEkPcW+Zz8FJKUE
LL8dbtgwmR/h6zyfnsirL2vsDyjCOfy6qUnMWi93VPQGLhI34ljSKR83CxToWw+OqZEfAqvkBqVs
GFd4L9rhcDWhgFsbSU0MKhw1rlBcIhQveoOjsYSgAH1i2fqHnX0LePNeeStsntQ942YstFU0CaSh
fEV7NduyKR1wJXTKnOYtw5eRDHFg2NmCEMmL9ezKIRqaSA7K7+eNvXFRMgvc19tZw8Z0IHx+SFBS
rbThYbEfz7aF9gtsEZIssMzMHBf1NKE0zjIIN16IuMLkrboqGquHjuer8v3tuOfvO3ppF4mc7388
7DDndA44PKvefPImyDlx8JQSwJfP5IoCEdxE937FnMqjcTFlZ4za9l5H5WK6K0MLNuZvy6ck0vry
UikmVgdWicTmMT8ZjtIcZnpBIFaQzb+RZ2MN1QKzPSIW/Zzrce26WpCtl7KVi0Nw4+msLQtw6IUO
stnM/fnEDVWuf+QtbxXYyMLPwAv1UvaB+M9DXDsCUCauDDe2mC8JvWcK9g/pgGq8zLewMvRx9b0K
I5sonwtsWRIhYvQruiq9wl6v6oyr9h/R8Z2Y2jNJkUgiHPn6/FlyNQG0dpRDRABaNOtWMcAYpyUm
F1k8LOM6HpcE+kbWdHYRtJ4A7qoNTPuY4XxKVGff9uswU1WkIXLyTL+QqO9JWLvScN2HVx8nOMyS
QWFIlQoKPZS4O898D1Jh7y81N1+fPoOE6sbzUHxQX6YFtikVtDI+J00P04D0EF7FYWGpuMPSV17f
nY0ImSBp8qqir50f7YvgrtTGu90pe30n6ra4KN59ujb5TQwmqZwemUDyxksDkhUuDw0RU8zK7Z7w
EwjKsB5YjmrhdsipAZvZcxxAQsAXwvQm4A2XoMCLuCIJ/9vY4P7mepdZNfHaKGFW1nJ+bbSn5+Ru
qjwRUnEon7+pt5vLU3/vAxsfMrccN0dPSbibziVcrcvHZ/3GAdgyM8XoB5lol08/685X6cQw3IPe
5EFQPSElDgvQLHabv5To3r7Kn+k9towR1HoamHeksCd1uOaACgA1n+oqTe8J9t0qQW+dhLLWYQNB
xSyr9ylsYIiHC1g+kf/N2A1MxmozOaN0SJBGeWMGUGXq+X3vtWU/kV+SUlx7xuDVi3l4Qbl3Zcvq
iPHV8gIgcVJsz/q/ZiaY4JQ/3ODqDtuEk0PNI1ehYaQJqVwyakn3ZulG8YhpLAegMiuJEXgOI5bo
wcKHZgY/fj0SHLS+n1//sDFf+pTiHxg2c6vl0kyKkyN9BIXlxHBzJf3fCBxxZYHyR7DOJuEjoedT
jlzp7KCvfpziPMWW1Mjsz/ok4fIJ61/DRqAuFyPOoBNdzoNvZysOZOHlGXDRkahEe4wrmc+pmwna
Wtizhhb/ZGiUrsuqcT/LCggceJBsXC5GxfRsWtIXPGEtnb+Z/My757SZrKsiqW0Qy/xpKaN4wAbK
G7YlbwYzaywo7aGvLNlPFn17DRQPl1Q+3H4Bm5OxrvDIdJRE87wG8qAMC/JZR7LrS/UcyAt8hNF9
5LctJxW9h3syUDkTBoz7rSXRCLgb4srBt/40rpm7hTxbWXtOx04Nrp99qEaIWR/K0fgEw9MmJwF6
4nr1JpS0nghJ56K+J3fPsiKWZ7UgnqNh18mwvKiRa2I57J+N0jGVrxhHg9+pIH8vqpsmxQaWxvSh
ScLIn93NrjcQi1RcNrWNJkLniFZUiql21vZ4OyMyMVM5Z8YpjRm0V3u04CEI5uUAdF8Ru6u3y6vW
R3mAizk8xEpfKcUK+klXjRPWIIoLDhwaqee33y/d43XWTTTRoh28U5u+b8+LkQGYJ6YHCwiDmjPm
NbSepgCCHORgqbDllyYGbU+UYPHp/hGmIo7/gQXPkTZXSPUeJSE2E1Nz+gjye3+PPFaszIos7E3q
F7awZGP7AXll5JJxI0U0wkkXh+4vv4XsMofjClbpEY+56A5aivucOc11FqWPrFVWk7q+FTdUvzey
k9eV+qquN+VwyI7UGVtWKsLyj1U8gNzpV9o9yi+dAdXANB8xCN1Mi1BOGXW0Woy38NEfrC2HlEzj
0HN51FoQhmeFhFNZVOKytLCoy0oeOAavYFNQn0aoUfyw0irgui6G6JONVM+vgOBwHXu9NydVEJBJ
TMzG2En/HWeEtMwu12tW5d2ZrtIU3ckqvvchGa1ouQYvbRcUvXiE7KKVEpil01dzvmctM7XBWq/S
HmExywvzCEerst0814jMlHJ7C1es8xwVSSNhVVpaAyuKvCKjHzl5xG1xyNqyZoIOPAIz2uNsQofO
iLVO3Djv5ActTWXTxaImsXaq7BxAr3p0CVUAo9SeeoxVt+7mEZ/RE89EasLFFkFBbdsWDozjGcku
UvOfhuGqgNYHQtjeAwDVLUssD2oipaNIl4y3J0xn/OFxZZo3dItPdLcgH439ZEBrPXciMNuhHCEO
lN/7lLjCm4hSmzrym8w+7N7ALDP13pR3Qckbx6jsXAQEnrkHoEoW4LMUXNLjVjgm3pTxpbkbnnii
MhlqpXB37PW8HuSokixQ2VG94cIunWtaJurfTMHpvhHzxmONJ15sSca0hsBnrt0CmogLarrz/Xin
UuqPvLk4+3itO9nUMVx3WKwgG2fWnuqdfMJND0yvdUwGPgKMNHPLylSu9/mWoM7Yl7/CyOgv4FO6
X6hLDKcAv/X2mvT9CLrtKh7T4KBqbfL1/p723KWUxqX38qytKK+guUIBytJBQWKdDVgoNBa/cLw+
pDiPencp5rfL81WjNEN0nIpGtfPWexHFyv3x3Pz5bZQNLzZmVOkfFJOq2ysJkbYzEf3og77evHEz
5Ze6KHUuTYCiE5K54xHHEQI4BK0CkqyTe02G3dRYdCtb5/cpskkvr/JNFiHbF8e2YcoxLivx3KgQ
vY3Ill+LDv7PuIJuDtKJQRxBDJ8tMq7d4AHDKla22tmRBN76npblk/FvzosSLqTd1sreMqm1G775
ZnJuEBS4FeUDx29birsJGtlMV05mE1B4JsfTDomOfBw3fxGKad0nCLYSd+i20u5uvNmNT4P1tuz5
excHkzHoygv+F6Gbk+MpCRek0Y1u9oLHpjGNtdxt6MnPs+xIn/saTGcHLngpIMXkldXAc/ouRe26
RVaAJxsS2POD9NBwl1mjOt7Zt1y4MskcgDHxvYA39dTB3HvEf6VW14s+yUAtLqaei4gWoCWAeBrC
O/2tZ3OhUEwwqZIocsrUofKF/AyR1KVfR4fGusjPodhrGW2Zt+OMK5GLQGGp21Y9vv31Trpgsyq4
bYE2Sz1tMrwKLOq/6F3Zbho4CbTi7ck8Ll/tdtKbRmI62aUqjA3qWDd58g0EYWpvT/z98LpansV0
SVydapPSTewtsSuBgry5t2uMMKgTF3fE3xoOQkhIzYWLtnu6mJsia81aq59t9K0/GvBIhvgOkoYo
pW9ZJN6AxyFTUlvUCGErDKDzrOAgO+SuYewNXX9ZSag2h8RB70D+jRUY/Pk6iUNXTYWI0v7IGCGd
1cTk0ecItCcYKCzJ9/RUUbLwNjj84udLbi35g1zl4S/1ZzNQX6abNpp4CEvFvZbnXD0MO/DCo76a
3tQFDPhktJd9qvVntBlsofZNKiqbWtvKC+3tTj4qiQu/y3whbmD0KWrx+XrzNo6fbWimDzO5TTCE
LwvhhD3v9Kasq73WwWqiLJSvbRmlZATL7+Pv/8IYa6WIpQxYBZ/4ACLj1POp1lFk+tMvINNnV9t4
9WhtqKgnxomUKzEqZQ/J6ZuUrpiaYRtGvZ3jMTJOG1hsg/YmVCyjR/427WpD7/eOFs/dMJAcXjBf
NNB/KjqPFabqiTn6kMPrpszsRlMHYq/LNikqi0zJfNJTHu+spW5xXaq6RTLemkMiarikK/DfVAI/
SjDQ+P5o6azy638DnQ8XaPwTEuBWnP7pBCeclKVOrcskrEawbMvRbS5gQ8jVm2Pd6sslOm9iXd0p
lU2UTv80IqUxV4x1RKUUoJOXujvCxIvfquw4v38sb2Tre8vjKE3nnE2Rn0MmY71D5LdnqTPJMfdg
zzlT0Z8Yy44JbxX+a3RoShAgnhiMPLEBnaSKXBAFNHa3ePc/G6OPYMYlmB4zIfulkcytDxS5c32w
dT9usbf7PecdRyGlyKd7MwfGcpJkg9stU8G6wawOq58FD9HzJFnVtOvuO1tvnF42xWa19cirZjut
rNm8472Y70ZNqfzdvK+1ETdLb873+7UakqZXnPXYmQitfjLXvWLUZTN+1EjXJpGoDit6Zr7SPdoQ
F2qlawJrti2fhGR9kC+PcsGYtpalRPW31sxCM2a04q+mPmeqdKXvIrtPGvgA0y2/kHXtZ1C+GEaT
I3qel4beGOKvFrnc/+qQfqVs2K70ft0t3qE7GTuRh6BHw9/MJ6Aiay5fzG6TEz3iQGTBda+pINky
lhuYxiu2752MnND9GFFY3dEFXxmcYyllcPL4i9ORHEktzykj7iDr9qlbWjqgpJ/3XFAHaN/VqE6H
2fvQ7+41mf72wX7zPyhIDKrFRp7XMku06+UtEniFGHZbS+OhULujnKhzTWSzkm6jGgWnSPtSW9J/
W5Sl3KbJsJ1Q44An8i5oxOsEq0SAoTyc85MAeo7OU9JxDRs3m6r2vZHc8PuWVZkYrNu0efa2CyUw
sEraUsx9cyQg6rVWZzrDMsuRqF8NxctGylkVu7wr3loJ5qrROWJOVYs76k/hl14gaYh3g1a45GT8
/W+6g/q6Vdpe6hOIcdszPaXFpP4fDd2p4MCnAxX5MUUllJ3IMymjlUK/62FaSK752w0knXnqNfW+
r8mnUINOq0rXAt2esdkw4TI1TFoV/bkM5OnyBJY5ZUkCiLQDbZj1rWf+BEoVrGQD1G+mHQRTzOHT
yUTIFoiCtKdH8gR+MIdN6OXB6XzkEZqlJd8liBMxg2+B3yP09SOuKxtgz1RVHxZyT5TGEHHtaPwr
poNFyXT1msPf0prgK6nzrZPFn/PB3r5q+43E/KsdhFKGXC8VlwEMX1aSmrN4yDp0DBEVbUx6ECrK
6Qh0qgKc1tkkUAuGzV3jslF7G1G86QjNUIULO8lrlfql+m4WaX82xqlhfDgQTNuB9ywZOa+JsTA+
Y9YygfyWPFhtAB0/MFI2GRWQfsATAKebJFzXS58cU3p8NREvJfDY1RqMXeeZkJjR5OQmsbUVpAyg
NeDD+YNgyaPmpL7e/FB7X++nLVIgb564j8UVi/IRVABOU55s3ozf3b3j3sx8D8aMdxSp5TwF66DV
8FyP1o1wImc3VRp5FI1dcMNNbwoIKchQ+wv2LFp6rxu8vZ+lFXpS5oUE/lMQYo9qoUXbEPT0sxx6
RmC68UgFGAhiPKgUp5wbZJXhk27omEV1LdfK0mGUkiyYDDVXg2tXyk1PX9l4+o1uzhx+8IXQuJI5
Dej0CMdpdbOK5DshOn574OPswV4hbd+mdzBbyuI3RF7FtrjNmWSEYDbYRMMzrnYcYTcqZk0Xvfrm
PvVzntgaOpWCpAGomxt3G7jDKFmqKbGooaqLjMITmYdjNMjlvr2IZkZqth6czeJiSFpj7ouqk5nm
LQ5PorBMMtgUf/pOJZp3QnFrAHCB7+ulEvJUw+HMphwMm/QHHjCU0gMY1zZThwEbPFSOmAuRf2OR
Man+vHJxVpPJrIrGU6kte4H4B1iGfNRcoarZdciChEIngDLyFy7DX5VU6tkmX0FUvtQJEn+b/2JP
+AUEpupE8LhxpATscSPW1c6M/ZmSkUdsQLro9AHmSR5eG/FBybTZNnGU6KDOGQmry5LltlvniCIs
nwwISyEBqe1KOvD4GUdm+ZVNG7BgE5MdGmVT8sKy8vEUxK7XseC6XI3Iv+rnoPn4Ucsdrnp64Eb6
5fXrzEgMqPeZrjSjJsNjCjl4Jzi3NaEurHbJa4EF2e0eVIjZjjOYNm8QXKoCXx7d7jFn9eHbN+S+
Z6iRamgQ2kb7mOwPT7mDgr6EBTPt5vx8n1WnG5sVUtiLaIbwi+mGTQAIlJ32TJWcuHRJT0Dl535M
/9z+zoBpBHHU3wEMWMjSa2eNZAbcgN6+GIAP6JL4NuhM1ltszVuxluT1ZzSq4wH9JnUBwoZCXaVG
UzNQWkzEMfCol0yKMraxMxzaIKvZRojTKuLJvN9zFTa4i0LeFcMt+D2DpCkPO0+TIGEMETiUAptr
EeC3m2EzGRyXgGdux+VZNyg0iNDhfHIE46gMV75LQOHktS4d2Ezn4Qp1BN3E1lPzKBdX2S33ujGX
YRCSCkmNM8vqybvjWCnnvhAeIS60SRpfzFQdrzOoJ5BEJJ8JpeHvvuvmkF0Q8hewO9mLSKtFrOFk
pRqF7lL/vkOlMeEtU8+91cepIqGzSsIrqVf2Vm/epZadjMdwmF+WDpz9rqb9k5FQff8ywmsvqnHn
TCp+ZAug0SJoYUs8c0J6R60SwbuBc3Dac7FLdhLFfTMabImDlJlxYd2BKkYtlcaDIxS3bB6RSr4C
xbi7RaIsGa++IGVR3RUAEM7jFmzfiIgRofic93vv9X3K14r9Q0UxARoG0aWj58psHz96YKt45DdC
Lzo6xL+A8qts/I9z3DQoqYCEJM5oVDQmneSSPkYjB+PpwmCkMdR3XBzXBPmf9I9/iZu8mFlFARqG
xbsXBGJqHsXjAfoJYWnG+fqLetwPqJXXyQASq+3Y3E3kHr/nLwBV6dJ0WRWYiG4P3XsJ5wq/J/yJ
ZVHVgz/0iFrg79SGUMaPwbwjqioMR+qwpO7mySyOSxbW3Tf0MwL7W3uIIGtLtrshi2JRBDZm24wY
Pr29bA+xUuUEQTP8TNHN3aqecgPL96hUV3W5FSJt7IMa8ffw+M8oumG0D7RiobFHqcdllDAZ8XVl
inoo5/+qTr3jvveUSFAeKeI3k5e9aGsQf1fL+j0WDE7mrVhb0Jr8sZ6eTLhZUCgoHj/ybbX3RS6v
PDaNcwftkHfTnc7NWUARZQkhRnOMOflhJH2hC16P2XsigVAMlLoviOpMkusR8ytaxw8lGidvsy4U
lNqcy6YkFsDvsRYbhgKUiUOJ6UMKsY9wCRlYWdIaEAAOdKlu/mZv7XZnTmtP1ltGuk1F2yjr18MM
dKqPSACXyqVbrdtKhI76hyOl3LoxFmiixX/6+6E7UukdOa2FtcgE8SIj7knWY/nL0usN1NQ181ME
E5AJx+2VKMN4qFb8O8fyjM/0WtqZBMh67ji6/VJfQziTYdrghLwcOu0NkAf7vgBcBkgjk9KIfWTh
o4+nIqiBMvkR8ACTzbR2kNyH6oQNbsH4G4zE7OVvNupVfsucpSS2ql/DjcSUn1J2bUQePEWM+ty1
zsHMUaIWsCgOqlTRsABIg6pZvy0UuG6QuWzZgG7qr8IADvp8QntGTuC2qo2x+6TQVKSfVicOpwos
c/jHKQGz0n3bg9DSn7ekQHDP2kiMBTbXmEKlWsJznJlv+o/ZTobKpAiz7dg2+4XY4R0Vo9iyUaYZ
FsZkechvRbTPlKpbBGtZ03eQXKbSQ8H1QS/hcAltrQUf4VNgInPybIPgtMI8SmND+mZFdGusjIE5
XQCACaAnqsPBita4u57Dt2YwH5peR7afKyHELFXYbq8km8+c87AtzS+WJhJh2Ui5W33mm/NOuv1M
YH9kQrj9PGGDYC81o3YV1Yu8QtIj3f8BGX4m5LaEWIbWBIAofzMHe2V+GJCoMp7VlIQWufsMN2ps
cA4lkMhDd5lA2WzpBYEj7Bc3iyVkLEyuh6WRFxDo3i2RYCZKm7Wy/D1SRVPgYoYDIwTgd331QPBo
q8rs7SeQGtx5gsaptzhTa5SpWL7IwzJAWzA9LRO3fpGq/BnhJR5wih6YhWuHPS0kDJgu/vzPw2Se
q4p3OCqRftfVVvxZ0d+krzV8ZHyjdZHC5inQH3sCxM+DFXaRT2aczrpJ1qyZuhBC7cJD+EdgG9EM
U+zF3Uar0n0lWU7JiIgCqBxwX9inNqn+XYoefkx0ClbXlyR1xz3NHCQVXDfQaErEA9F2RCddcuKV
qCc1ntdOIpPv7BVXTZ7p0dzL2XcQWZycehOOpqtXvtrK7Q+j5yZ9IR876wdHowiBjh+VLMndhLkA
qGgtJv3prrG9nJe3n9a0tVDC+CQqod1+U3bsdlT/ox9KYrxoOaXhwwRNsymy7/kz/UmcLnALM9TJ
DS8ItUn48bXzH87zMcHF/8WoBp6/mv0rgD1KavolxV/U8uIzZHeZdKD1dnQ+xoy+zCdRIEWPJ/QM
MsR0FDks7q1xhb/Fa2tfFSMeIOqlQGFE4lzCYCBMnw/N1JiOL5UCvYPHiWuY4KBZvqotDjUEsN5r
4y7eTJtClAZuKY7Ag1pJb1B5O69g39/YwoadjSW5tXgE6f7g4ORvrH9zhAucsUmcoSHqjUZG6oO1
C/bnuU8V3Dv5SbDvr6L8MsUuSGh9QJEspY8JhkPf22OcQQwREa+yx/zDRwRCy6uY16ajCNfdREJY
+ccjA486o3qpuDhintr2cOVHtcxtuas8gvOa5aEEsaPvxurk6SGtGFVQeYZ8Pbpt3AZ65qQGg6A/
cOIwG/Hrr2bZicA6Kl5DcHCkbeEwZhPlzBZeUK6ZX0gPCftPAELUH+mUAWpQWdfJetQGNkmFUkv3
vDLke7oD3Ss1N1VtJ+clZX1mMGEPYVLuMDcu1InZMv77Mwx5i532AgcJQn1lfZeO3rPIGsjdlNGk
Zyw7v72RTJ6btcNr9BnG24czjO6vd4TH9kzjU79HTybCqFndOVYp3dZhjn6eQF295RKxSnLG6WUw
EedDIa2cZbE2R7aRecEbExgFyoToFNyLuBQEoR3RweqX1dduJ/QZ2GYbpGCiMUyTHH5M0FRR7nqr
eS4g0qqt4APGbrcxK2KCg86TK6j3praxz3npRVkrCU/92OVA6URs4DHnk/ApjDoA+3RWzVKD6O1+
8ZShDlzoiTfAZ6wsEbfDEMoxXMprZSfb6MvjhFn4eWHnzI0xt14NpoKXsfjsjSWLaDj/vZkSAZMT
zx3NnB8k/Wq6CNeMecFVUF45IVhIwo+pbuvryf6jUfB7R6dotK0EEwA0pU99lTYnFOBTVd+kDywX
VtthxSwgOMW+jJIQ746AeJ4pf9qzS+Ot1Tw3bTywPUw8U0v5Uv8Wpd3cR/gC1noU0Cyi2ugdyDLv
/6ZiY1mXQdGs+JvbyLMyzz4zags/Y9CuLD+GKWN4Lu8ArfsQDaDEVTGb1vQ1e9IHquIQZcXUtenS
ZypZSfRgtxrPN7uy2sAla/IEWdYDd7zrKe38Ba6v6X6wMsH36xrVk4p4o5KnGdkOULYz9DuAtQIa
YQ9KGE60R3BosYU14VMtze+eVaV6+9k33fd5AhxNumXlK78Qmqvkf7LjJFcXepi//9Tmdzhqqb5g
TxAntyxtFTNwZoCGxTdF4YTiNslOM3SoW+uQVNwljcScqE4+OvHqzdYkDx2IFaqqEIGKxOM14BFb
0f54KoSQnIB4bEINvVYqENSYyAgLUJBpeKKV6uJCge30vgc/pdJC5JDB8jjKnNHqq8H8Udr+RXV+
AdeMVo6ihxJRKiKs95KgnPHknaoPUmSGRI3yrEICdowtrhLWmeNbtkySUz26cSyuiMVhYZBfHjPR
5hvY8GdQKY+uvs/gXLQRyGPogUhZ5MTdnJoWK8q/tTQcCfrSbQ8hQICxsDrAkcxb7z6fueGH2Pei
kYUPbjBAiCQ2JP804+dsvXM5D0/lvmpR8QdtGn/2SqS39S/ReFFDTx2NB/HUulwzkLh9TBhwZvFr
pCN+z7qF3nO5qzx2zeKpoFZ6VUqcHpxqRWns/y3IIILA+PTq7yerVU4K3bFpndJKQg/wAI4ZIUPS
zLZ9DGLzTCeFMeEgXn9gZSIXET5VbCla6778wyHyD1CRvfp+IOE0Xc4SgQSUBx6yPf1Aj5l5Vs7Q
81FQ9MNRevqG1Z6nxR+h193yrgQ7EvW0Rehom+gZS/ZU4pzXWB848l5nIq75JQt86qX8Hk8H1Rnr
RNo4ptf6d1zUS+Hs2dUiwKcIQB6z6YLkLeu/w8QJjbm/vRF/qinfAawdvdP+60oFyXqMYwfVKwUh
kdWLY0WPKYXyc3icn+ZIfOpm5qfY5JTu2FEmWyj9NzCNE/RSb1Si+KIrg2MQHNBndb92lYmtDF0P
av+mr5LRHscSRqLMyc9rPvGRjo1yUzzJChZmRm8hddHSYQghUfsc4ruQ4+iAXjYKmXsdXDMAWhuy
eMm7gV5qRJYN7w4S3NHEQbWOVvkVeCB+/NFg+lZD3h1W36sbARBCOJP3SbyW+TO5p6i9YmjgYK8H
XV5V85gtmOkJiobHdV4e9hHK61oK8jnOfbCyS/4U9NUr2DU3aWHVohy3JYFwnHrk0LEP0T1pB3hg
95kfOFIgih5OPrcMsVxb9OkqquqQR/5ME6rbVtFAgh4mZQA6ytP8kTaWDZazbyJP2YvVEReBa81I
wZgPCFCY0X7Qi+8TfE5fucyjAfEqYP98ETn7UcynhdmhI0JsFWsiTW+BtY9+jshZ+du9xfRUlDXZ
L0IkaBp8Zl0p5PULernlGBYvlp6euZibQJ8RdmIIzhRmO8LbyR/14iNvdDViqn9q3rSLEmCP0Sid
vXmXAHmgtBnXSGVq2oEda697Bvxe1xs2S/ucZ9qX2YIQRouuLzFkIrf+GLZGlMEnGOLL+l3UBQX5
hB354WpInYUsabiXiR0ZU4uqd0L84ylmoHVTtGRODsnuuxIBTrlmRVXPzJyMGjdbWEc4QjjoamrD
lLQTDlmdvOyJ3kua5QC5EOulZX/FufVXSIjUwgfVubMf2Ek9QFWsC6fjXjeIdpWB5+8FzJ9ijDXX
g6IAqTMWBpHCSdN/77N7/tSBnvRRxWxXJj51Z3qRQiDteJyahneR90568NEnA4/OWlA4ueCquaRD
yFvXtEaMXthHhzPKAFtSZ8y0Q0Vwxs/2/zSsnyEE5FcHxDsTj1GU6cwVPI+xEpDZPbldxgjEGvQI
Bbjh7NyZI9ARj+fAso/NvRRvTCSKRsRLzaWTE2/s9tZaqdZgeDnbJYd/deSQgISBGeOeSp8AZwrV
qtgiDClnNjY5sXfpZ9C7L6Svkq9PXw4Q/AwSuaJfbevc2Kq4FYJ0d+es6Crl2YhVY5yo4S+EFlHI
r2GQEtJExJf5BNMwM02ZHIWJ8E5tgkQ/2wbsONphfH6adfjJd/UQgCt0d3QLmeg18vMu+4CeNSM3
e0aYPzYP4oaJ17OAuFb2nJmmKF3BUHhhoxcrJaQVu5xNVfOhmkwfBKwTkPwmZP6ruYcZU8VK19uG
0GrWSqI0gTUgD7y40HoohqPVc9w0DiVlrfePmSsy5MHYyMQWXyWgxkm9jnvBqfd5eAk5e+xei/xe
DGuUWRpNr00FPKQPOnnuQp1vKmFkRQrz0WOo+vZHDNopulnFHK0eH/Vxzp7bv/cUON1Br2tSc2Vo
01YTQwDLCjss9y6eKd+8R0cbQSEtzOl18LPDbkrXriEtvPxPUUgygEg9S89xETYozpEKCIwihTvE
TVPBk5e6zB/+0+BHc7TD2Fbev11WM1Iv6p0gafME9mgcwreLzU7G4YaMCg7yR5H+pypZ37qs6oBn
EXatRrt9l0S84Aa4dhwrItUiF5WljvwuCJgy96JffSd31M/PnwrYJDq+rinAaCZ7PyR5I11mG6sN
BTzv6kDiJ6DdcQGeFSowC5LBgSbjxieS/GZJbiO4wRVoQua2eH+4bX5EzxiA8sZ4CjEOb/mbWHPx
Tj1W2Qwa5Y8TjyVPopF2U+iuqKb5K5d9+MphyeAo5SyJCPxLVRsQIaVagUY8SNR/JCZIY3ImcYxT
cXLW8Knu8BYU44OI7fVxhBhEUN5RXPG58QxWiH2oOihx+MI9Mve7N8Bo52H0/Dp60x5qzmAJcm4k
EBswbkHVTzOTeVbQtcluxnr70trg2DWK2UmHKLwoDmk2BpIxxEtA0ecCRm2xKcCmW70kaRcCcyq6
bpRZQ6LcHNzslJ0w4H+Gp7ZFx29SHciKXL+asHC/Jj1Em4MPIGDvhLX8f7owRpJgqSX8KtJEPfAS
IZydwpxa6lWkgZZSlMcq/MoM+b5dMEt+N9EnIHxOwvXvz3frXWw5dJQ20CiOxxZLVaqGugnMevF4
SIR8vbfvaJCSKbkQO0FTDbrsSM9RsNZiJPkS3ctegGQOoRIFHv1pSFYILa/O8VjPa1ZeISm8SSu6
8ozMBWyFqiAox8n+dG++C4QZfnTqso84T1bCiZsFXYdRDelOL42+RMLPNsyK+tJkuzo2AQuGwLM8
eHItucBlDOT8uCLXU5VxIk0OPqvDYj4yGQjkCZn4yMyA0Hw3m+UkxOUvZRyU/ixONx9t1q/KLrXO
8d6ZyDtn5f6lb8PSQ/zgC5n5oUEtzbbjMQp+Bc1EGeNTyYjh41lMysQy9Bd8nEr6K5+PQ0ocFRJ0
VroASGbQAo9T9unpWswI5LqqudtKW04cQgog6zuvV5ITUTmR86mRYttKnagGGVdckSIgNBgERmWJ
WzfYfeP4iW2/pMPffOfXUy70DRlO8rSfuPvGqI7mrZLXK20K/6KdTMaU3Q1hSBYRnesuu7UeLiap
DBKle1Pjb5bZ9HkwW38QG9YNdCV5cTBah+DnBDkChAHrSyLKKq79i8pnmYwneGy4k+oNyNNgDi/c
t0FoPTreAHz3gxMmoj2C3M0YBQh0C2/K3hUXMu5qnrCjl/G/KP+TYin0PYU0Nbv9HvmQ33Tygt+e
6EWjl54KsvdaqhEeEgKcOIaxEPdVfFHvfIpyPbPGRIDF/jhDVMCYyWJnq7WntPsYd+cTI0GuDwAJ
p94XbguXOsXa0DX5MxQ1V+wJKMGl9Qx5rUQ7y+LC7SPZL56W+2MyjYBr0JYWD6hStaC9A82nXBFb
RHnkHuM2rdZOfP5mEbR1wnyqervH1mIQho819fUFrz4oXkYVN3BXs5c1LlVJLsKAl+yNcvR7EcWj
QSCZZqm/vgHHZGwfodDhc7eDQPrzqHJ4nE874NsxD4+RiP/oLBNpxFyBkJq6IAtIUbZh01klUs1D
mRu7+LeGTV5bWovf5cdn5FObEQX/Daw2FDTGSpMkShfHFNQC/cCL3VKg5OKjLEWYUwX3rnBEDqKP
H6vua7TC+HLtKd+ri6W0iHidfM3H7VqdtXuc6HHEQsoDNeO6jz89bs50Avsv04W3i2LO+TUcyLZM
uxUQzBVAw3yehhelJXxL9wLepx+iGfbvApIxt5IZhf9DSRGEqhYut5IG32FJOtM5bG64zpzhfDEt
HgMXO/iDW3rxPY1XrliNBinGUIrMYXsMyl7ev6uirgpaKncNDOFabX7yMO9fLIQttaTKz7yuIqrW
QnjOVS7zwI4zGsXRr0oLyyMht31/fZ/LhuUt0dodskpK/s5l0pvScZ9oFaRMLEO04Bwg9rAiLBAU
jqWAvJ9PUTGekxtq9nWk6+PypWqX/GoLMk4GyXV863c05ZhZthGKxXXh92jWSqm2TcnrqQbBNyKX
W4NOhmWC05QzHyBK74wdChKQLLd7ne7rvmOV8zCMw/m5aa2YcCKilv7NR82qRBvOsfcviDUM68wo
IkHviXyHNseqOCYk+EC2OrcR0pl3ij78fWBWh12wW4135ivt6A6nUltSV7Gzdep6cVbJ51jHUZeK
Tz1MXAD/CVVI34LP1uoR9tXGODrBsb2nfZkKducWNn3aitEXLgoIDaE5KpuVM27sNEs9msJ3PGji
qtPWIVUhLH+5Lc0bSB7t810REbVtGc667R3eSbx/10/JAD03iiH37f88K+3RsQkd6Kbx3lZfZYY2
Z5oXkm82L9JpZ2t0EBcfyEiwKlVUCIUeSAzdWbLWkXQvug8u/iakblWrl2YzycYDHI5cxvmLIPoZ
esFZITF0Gozd8I+pbVDZBwOcbhCfq/7ooYsB6pGAQKBem2h8OaSglTs7waIUwdIbMM2GjDU5rSml
ze8QqHgqrahp7LNrVSih7hG4UG4IFUr4bNzUJCVLIIznfL+D4ls0MClrJEl/7mnYB23IbBuCoCx7
NUfgOWM6KIqn8THuf5OG6TqqMichf86QHlyoq89zp2DPXMqpxMEXJB+vbHN5UZeIjxuvvI6Xon6a
JseFII36xga1Nku//Ls0uTwiozoZfP1x7ExW1Sy8mneEmfB1SKMBZN7GzLlcHGeB1dBH9KJpSnJy
0Ar67dYYYhvo2MvRi+1zAoJoA0e4CUttCTVdvNb2V7miyy4TdQRcPuczf9oaqFqBLtFvMctEoEGR
3JcTXBvEmV3Zlp8RuR8IU47dr3CXEauUAZ9RkU4h+LxPqieG6Aw/1IRNWWBJcsE7B6Y0E054OWvw
743Gu13vMTto2PSsQOjyhfMcOmltxXr0NlLpTsEK3rO0kk+9zKKDlx+tPjWO1yUWC0Tvx+q4C0SS
1zUYFVJA1kDHE8gF4TGjoNAbIwTmz9ln977ntQe9JRsxNQa0wn1t89/k5plKCnetIihLDaqgFaY1
QFNsPeMPlk/txWTrLnME/uvcWAYRVeDT9T13MgySdk+ZvWoAVkk/AYP614lUg6MyZO/TBONTjCT5
Uh7iu/srkgXH6Bwkz4fTvfAY0SXdn3t4W1bo98qZPIBwHUTEkN62dBu88DrW0ZvOtWikqIUMga1S
uUQuk2e0SNRAcC0JJAHuxxpQhhb3tBd56tUSQDjd4Eww4lmFU7rdsDb0iXxN7SoGdyPvnetw+UV3
awV42Nu7gQ2DsRiBjchiy0tAK/p0MzBveHvbdYfzwT/pjT2cLgiiuq/okk6Ra774/3GnQWm1sHzK
3PMcuo4DC4gMm/F9ORqWclDJMa5oy1r5bYcSUg/iWohLQxQ3AWw3EVyZqCkmyuvndUyNMVoKD+IR
NPS+dbDyVXzILdBp6goPpnBATzr/zz9oklSNVc0cSnpicZ1Ob0FJq05hsfhVw0bPLnC1wVi5oaEl
d//YUgo0VMY+jZ9ZMogMfCVpBh3FdMtggrzUrQTdgZ3yQur39KojzPoBhhepjijGLbl4pq19iFZq
dV/RybMDmBu38dCCP0f/w52ohoA50gNlzUuIZn3HvTgxsvROQpvu7byzdbfZ/++aOTwB2BdX+TeV
UgsapiAdUz69i4m+VLVMQWzvSeh9EaRBpcDYCHNdJ/N0BkrIvsnuzwwfGj4xKg3AKosCv+RyObcA
WkajLbEQEd45/9cveg9I1EVl8H0MJxgUGIonlf2A2ekRdXU2BtWE9mecvYwRieZVtmw8gbpqQvFi
v18c3w3Vugr8LpJmAjLYd0YDwbR6xmWT9LohIPzevaYXNRJ73hSgAelPzptea2ZAqQhEUdHwKa6v
/cq2j24vyI60riNlRZTQg8ZdiZljrTzawGtfi+tv69i26WFXaSQxa8jsF5Te8cApYD+v/+vAmrVD
VAF++yMNUO1fKWOwyG/WKR5+n6yOHM91sdG3qURevpWERpad7fCw10abUNmPIS/upAzR3+knunR5
5pG2KKEvM/iuyL5HIC32mnGCoDJqIhmKJCHMswFysuV+X7eBN7/ob20cu+iuYJENoRDeykpKAiXX
IB24BkWCgoMtgRxpE8HOkqMijLFSlUHXQNMpDNl9kYqQTaTaH5uDRKhAe7QBDWGKwA2VQB4Ox67o
QS8fnapP50AgEZ/76hfUFFSdVWonjUDjEIgnenCWpXADOLUMHq5EYcX2RS3uXZwRy48Ky5OOb9bQ
mssGpEhCLuV9R8b40m0iCoTojlfPCJwUYc8zQA0kP43IjIOj756ikGtDdaDeeDZTOaFB7zt0332E
ep5MSztgZ3JfRmoJV9v8sirl5sXmAG6JtFbSWU23rbUke27Stghm1mW9ftvTJYnrhDyQMTbwrgzy
X0KIlA908lUzP9F3WAE+Hlk9pIjKM+0QIJ551r2bFmPvskD5VcKDF0P99KxORv0jxMkmkZPLAJuX
MY6u3tmXbIGE1V/mJajd+M5OlmBZhcdQEwUk2OHtpRkzRiSJcP49cEYtz6ZJVFhP+zgrKi/63b36
FwiqdbFVGn3LoGLuL1HOaUv4Ls1PVXnCTxO0G9T8nQQk20CN/9m9aSeKBFpoZcrjmz8DZIhGumfS
j1cJio5hFECGoUC0FHGW1G/rpC2TWUZCae7kDM2icDTYV1o5ltZLd2roxFcDrYoWB3a4b+1yjD9s
y7gpGRVL4wo4k5E5Hn+/7wSecLmlXV6ad1Ko67w1eL7zQZxQjWHv4hH8KaL0TkKjiFNTU7+d3gK4
st++Zp3j9J0wvGtpQocMuxZGR8ZLadvn9QXBZropsNB9UtS5W2XZ75fSoVWqthuZcWR+2ia7eV91
DDa2l/IFXDjUMaEqzLWmHHKT8wfIs0ypEiddnr3I8OU+k6aUstg40GRArNuteXHu0GxwtPkN6T4h
90utwcXDxnhnf0Cw4v1GfRka3zN/yHZTYVf9QbaO8BLlo7ZtdJMynutIx+FIwMmAkUiGphWxb+0F
mFWtdUiZkjQeCYXzi9zlMFiCn3jX6G/d2FvYs5uLfzIqvPJ5fy7n33hEmf5xO7YzYi37behbVyC8
4vwaa5ZuCdVD+UhntQ6Y0C1hFXYakXrMXy5FbkmL0s9agiuWic2v1cXDVr2rGFsDtITF8RyfoYX8
FwqQrYdCD1X04cTt1yx5si2Sebt0mjEtXU5fGl6+z42hBhAdSS7Wi+Lf0KzwOJXM4ey8PHG/Rr9k
kU1HE3CTawyDaR2uINsHxB6YzpKt2pmepOHYmEMTjGWAb7qoJCbYDYErKHMCa5ELRXbOU4syy2ZY
XXoGubbIaEulAwDJ25SiejFzC5qXxSvLkHtwMi9CTdFANPr8LcMVzlOx5DUEDg4i8y6y4e5Pa8U2
OpUQmxrMBuuIeQNLnVF22zlWC5T7fqgID6k79BsLDOz6xnONPukLOoNZ9BF2AKqmnzgrImF5WdQ5
r+ImDntluTWpU1RNW4MS+wci9wwD448G5sOH42PFbcejxUTcBBV0zmEu+KGEoLGW6WIwr6ORveuF
boOEudzLLHj7qzh1aqyOOITbe9fxYnyGNT/My3XKN/U+Qwx/l5YTLhPHLGf+bXDMQqRgY41MyBro
4Y9Wl7Xs675lOeL7P1lOFkW5ZcC9/Gps6T+qUZCkZMc1RmbR2dK2t0knHvNySoAqEJefdfw1M1gF
9ubLGLUFIyQIqyCnriG+v/mG/6oOtP1FVLRqMWu1Ti57UGcOChWqk9CQILLOSoMN1cHcPxcl7uEB
0MIRYuCu2SL5i9PxWyqr/k6CVf+iF0s3RB1OG6WAlF2j90ro7SIw+yevUXMdhiFCRlXDbJOfySdn
OX+0lpb7RF8HKkdauTmM2TPGcThA4UZm/OIHxRX2SDT2n04Jv9St86ALrFzJqAfq0LyGqKKC1vS3
74rqlAIuMYxDk1ZZY3HJAuLGTxZsnFWfGLEDK+EJYNWmBd3NlMoZ7HEAYEibFUUhHNN+Zm/cB3rt
PkwLy3ZQtzIW34EADl0VHE+knkI2EHo09/5ByuRrfpYgz91ZJopy7nyLWwOpVnc/aiqovov6phuY
oN8ENYjdFymp6uWb81MBhdIQaXuGAIg2uwSSnjogGKRn2mLxxtxKpeL7M8XZUvg7iCnf30pWHkGg
uYrdbZeSnHkU+bv/aSwVzUJGMQIWjLqoa5qgUvZUz3n2dCY2TJX6Ibm9laW3xoZLWnjl+VG2tSdj
gF/rDlx+s36drT+gq9K5Bn9LnYOCLN10AeDPAhR2FiYfLeb0AllHbB+U5LuBTlMA6EGR2ch7F1Xc
3SBNO/5A5DPGFD4AXpUa6NyWvNBLf0bmlKKro6crIQut1Nr0xWzkPr0vDnvGZ5Yvo0xFBSO0YSHR
0d134k8u47tWkfPh75J81q3Ndu5oQNIa2WK3De48Ocout2SXiz1uAfHDZ6MiN5yZjo60sK8h2e8M
e98NRfLo5315pH0LsHC9KNM9bpycAKz73uAKU2ZdsY+a/WFYsjDt5PPHoHieA7TEUZta0qkEFDha
Ld3Slt8G8NNwjmgLwJdz4WyPJoP0zpLW9ji5dJtiCMP24vmUUa/8qkhu0AoQ4cPoJRO41f1Z3qlX
bkyxjnkItglWOHmRWccfwBIqg6Pmg+OSO7ot/eo37Fywnn9aFZIbgbRc2HkB1+i+aZzCwkbQ8MA0
tV4fj8v5yV0m5WmpEVDmNUHdjO3ndj4REows4fG5gt3NqBk03GK1VdqLtXQCk2+m2MIqPjMvQCt9
Vd3LW2CfrdD0IdKmRJcN5ozJnEEiZtJ9vDQ8AERiaJxK8aebZkn99dT3ceZytOEJ4Q7f4VrCBj54
N0jvb7IdHnXqZDMZ/6fY8+ZZbscalZIjHHdnaWNuMUdmfJ3t8FpIjoj4K82/EDTVXTOcp7AqjZyI
rkGenRKOb6+SrlHQAz3R4QyZICv00OtmI1lP16ZCZfFiLx0JCxnW9ZnYysshZma7a+RZnnJCIwAR
Nr6LsLepnpDQEiXrnCDlhIbJ36jIN3R0viYMcXoxtvxUb1eHMOvDRmQzq+Qz/1i8B+LZG5fb7RyL
olFh0DCJHQrc6xYZSr4haZGhXluZiQ9s0YwtexEdk4MeGeuw48hEWoGPJXMb9tt42seFPp1p+1sO
nEeGkMMt+BxwL4RiD9SbLC7PtmclEOM5bAEYJNUdS+GwumGl3c96h22mdfRQk4b8HjMyxnXQCvLo
D2/1+v4yqFT9J1enekgcPXCfyHmIHiVGCcBxdEc5sTyxDKbyv3l0BoXb0mn/dbkIy+35JT2mkUZ/
1CX7OwqCk6z+AGHTZUhV2Ryu+9xGeepKipkXDobf1FreZ3dM4whi9aDTvgF2owRTH1cFZnnQvTea
n0WUFx9SD3eA5n+NVGWjfJMCyMEQpwqzPHZ+49LBs6jjDSD9LsM/AOkJPKvbJkvV3asnTwtt5T2O
Nk22LpJ0sI9Wy32P+VyzZcGvjOdU6NiKMB4XUIPWEx1gRd1Q3/KdmVAyWfv6iiBm3IpCJ4GM2UQS
4H2V111fIaRixkCaEuC426Tb8NJsJdwBbjuM1t6g3C+gkA8i/IPYjGH+780ximCEo2nL78Kp52M5
u+459KgcWHtJ9JbImgD0d49/hLSU8mUWe11DoFlpwQkzTuXwh553Lci8nTI+KSvGDdTgpmoqGtIq
AIfXqV0eqVLdcHcVflZt07ZPeUgcLATrKFqRCJHqOhzE0Hocxaql7YCPKehAM1WgP14HmK4JJotI
pVuICE5+27OrzKVTWuPnfN1thEGk479AS8mDIb7Iewj+TEu0WcwtosS441YeN44M95eIr0gDpvbY
mub4n7C29L6wDIKGqDTaKPkDkqbXzmO7O55G8rfErsMcM0X7rBPVszdnsZO47wB3wmM/ORke9ATo
5ZxMGajBaQF0csn7Ljzg7QE5uqu/hcdr4PBpBibwQWHuhnhhrJjCrNP97+jWElz+RXOpAr+qU+es
5qOO2C0qd0Gj94+90DRMk+Z0UxF3PykS3BULvlkPsjZg4jAK45I35FkP4i79n2fkq3ykLJgspwYf
XWoVi3PDx2lZ+A+DUCDwlraRkhQmoOYlI1BwF4zPepvDKMDFXfLLNvF2zwohnphhlJ8oqAIYmPLl
0O3E34MgSpLQfwI0szpK76OmfSIg3UkAh90qym+U2FRhG6t3+Td70VmRhutQgIkORbp36YPgLia+
AZYE8SSuti5cWXhYveZyBNk/RfpTgYqglPQr+VkKjtJk1sbifiElH1drqOnNMS9YMXToOcgqSaDL
G5+izfdltkQJ8iH0f0Pye/sNb5pTMXPSLsGZSbb0peM/2QPp3jUiHTtwdWmJkAC0Ftyv3lfMN8Zy
69ciS6fPt4O0OfBY40W3zffJA9/2qgZwJ7dXE6cgE8ySl388rc3C2APc1Np3A7NOp9QjMd/I7jpQ
K22Q/bsASb+RznfqHk1ClcYGcMcqwYGUOH19FbAGXq1htfOrDNv/QJ+IAQx7WqQwkUxJxTEMOZBO
VjBjuU8FaVKmtLLqBYtgfBbQFnU4Qdf7Jdpow10SxD6cCdje7g0z8liagx0Yj3UW/DC+nWVoRybB
L6v8wV4HaCVnEhJavHVF1/4JlQKdnhk6Zjnoq5ywtyo4Tkl6ChKPQNVxvBeqKaki9c5g4zNyxlLr
Te3Ko8Yglw5USm639R93ktNFA6N9OoB8m8RcJr6ridGWXBZYBQLwEYLSv2zVqbl4ElgI+u0NI7Id
szP2fWqTFm06hAaB494I+OgW1Nd3/YhZ1nFK0B/QlRVzfgXBepGFeclGELckQZo70XUeaumKfjjy
NJGrFjBqY+rH2CB2BCQOuzytnaw7UuaenAY8xignz5/wczqzBVpKfBRqWVqko2husIB7wG7IAb2I
jmYQKWg+H9XMZgDKaiOXZ/RLgoqW/IVd1X6Sa5NkNKKILztpo5+kXsaT26kfuU9e2UhVSYiWm20I
1Scu+gfMFSL/VnqmUT9sYOF8PMCbYnbD0fMx1Y6u5U48tB0k1GhIStZnzRhZuTtHg84Fve6O2KDA
3yvtbLT0QFFbTNcoRA73fLdXSf+DGkVrdsEOPbrOckW2RVkT/za/Z3MRRFqD4ZqcihFfJ2XwoI0Z
YC3APOuko7+SV8WcJRI+G5m+Tij6cVWTSfkN4rKQwsvfy3G6PKHTfpDxZT4KdNnuDHbtnhSplvVB
JBthXrT9Ih8mE9rcBGn6SkIo8JVRVo23iunioRKLI0jo1gLKzqGQjnBVstbw31JdnWHF2Aa52Lrs
5FCIGLbPTzNMzxtCQs36FSbIJ8NLHa48uARzlpPOVVKOIr0BizMxHX5W0ci+zYysXtXhG8mizPOh
XX9a7qiK27FxnrYrU8SljpmnJk+ajI5ZNUwhlxLjUCH56XKeGkRGaF8XXQfjvHp1XZoISyJ72EKz
qFoutVwMmSrCNoWBmqeEM+OzwI/dx5PjCmgj90lSAwbOYSD9d9+z3Ko674X1e2eFjU5vNQfJFHa8
YVrIfpghfr5jTH399YpQYyi7zu/orSxwhvhN+jidV+Zqc6QLU/1gqKHVgBrfnDRuJgglDneTXMWQ
0lghn8ZZWsg4VuuMla/57pCTls9CGz5RbOVhlwe7LHWr1rNV4V/dGcFn8QQW9N/2uZrX22cwgFFM
SzC2qNHuxRMBX9LgudigiiZZctBSdPxWLOuBBylEFSgaNbt8ENg43UFyX+4KNpKe8yxKU+sKVlmI
HrWYIiCW2PC8HjypiKV0SkPnpw+xaF9pHb0UkN2HlR5zc1E52iGTeCTY9vAe4nfiO6opkqz0Ko6V
quavXz2R9R/lMAuk/DPKftLK7kTt/CZ2/MqzJumwH+WFW4U0GdeDVc9SBjkljWDnzX+H7bnG8Y4q
z92W+qXkCG+CV5lu5dOqsghmY6EHFvtse6239Ct8+/ge/gHGOkXKoDuL2D7Iu1xpgQ5sY0Ww7YyO
s3Z4CWYk45wRrAFJ0gFUbVlPEWwO0EWuOPFjqJJPcaqXCz39Rb3J8ipldQ68SpIHSk/5NRLGwbE8
ADvD9EUnfbReKxmiQVkxlUHLjxgp1n8RotPhLYSB1uGu0th4/4HaGUXR0rG7YyCrbG45f/jpcrLC
CaSUqRxFOwcTdfKzag0XfYAyVtyGBQrE2iknyBDSZwXzY8eT8Dps20LoVEJGebkMny0bMDoXLXwx
pVFQw8o3VKCgRmsqh9+ITgfHZ40F3uSN0q966LHDmvTpK1n7kfW5uhHzT8kqGEWQlpjeZngcqqhQ
0trVRUHjYYz2hBz0ithA+mqBalkpEWWeMRa0EpI/zX/g8PK1gZIDvIVzVPTcz2YYiKE3oFsCaSRw
DN+zBwHJknRhSyoQqOePxV1mymsOk0XJlCIqbnWuAv4a5aeS2UfbdHsP18Dbn+FQkCLstY1DdNaX
SOX6fQoSgEKVgN90do2wDyxbGDSlow2SzmcrYS1srax3mchj9zT4ouXhPkD65S2TSHLkhII8wC7i
20htsJTM0zM0F1zrLIv8pCL3TGRpDM2xqkrNEPWnEolpOcOCXfqh+067a2XdHmmArPPR/Shnvlb4
bbePM6/fAo7FPgZ+MGbhfGH1+D0jVMsgdai23TmXOrCxT/52/PEL2egMmmw4m92FRx4/LSSa2ULZ
aVnazVUCoeNinCzGzL6LnyYeKGVOqNoRyJj5gm3KnhiMrPW1C8sp6O/rXi8VQZ7s5VCXGm6mWdE/
uBySM4oLAX6nQnQ2VxRLFopDgjAlvp6uBMgwkDp1jetqd801nNwS+WMZN01YCwckT9O5RLtvlEvx
S1uUkINgIYt6BhTpXLacBLp6AaKoy6jmfVrm6mOu1sZT61gUpt6/QkZctlj3kMPGJClNXRGmwsPZ
b/yRzHO/C3DTPMFMPu6yqW2imGT3IZYxnjr2lQCZwU19uWFGg77SQ2UF1ETSoO8GbLxHYashdQZu
aoRfvt/CFlnLSe4K084A5YLtOYkNa6nqX+gs5Jv46g0cDhG6tizAmaEDJRUN+OE5S7ZP0ceKwtar
f5QOjy9Cha5ZvSc9kdpJfT07NvjoAimovCvNsBU1/UeUCkV95Ype9qz6Hk89BAvQ3wR3vp/H5+MX
s4H9xQW33JzqHuMDH7nXoIoD+RRcb/plXjpORV2FgVbNfUMY0SFCEUFFW74bWPeUDpt5rP1jylO8
HM0b/V3hlPyOVfeQz1nlCLqFB1B9nk9jmaVWrsqPo8PfeoX9TfY8Z0d3qMqTp6VjEVFoHsESl3Ky
6NMBCCdRpnDh02Gb8Z5RpkUkU5rjuY4sHL4NU0l7lNC0pGrbJbIa+USwd8H6qZ3mgXwtsP4umJP6
r0qXbsZjUVI6CBJzLpf6dJ6SGJ45rHpWspkdzjSJlVPbWJlTD1wyFoHX3hvga2MitFYs6/NVLl3U
oFB4wIWDJHWAp83vba1KwzmUyGbBFefVAiPsd+BYp6dWlpWqRXila2qnSK2eQmp6dnMPVvRFhfda
lNkNHKvC3WKNYQUWenptDfIcrcsT0ybOt9nbxAX+KZ4pCIkUY3xvZzwOD/wkyjb2AlHwk4Kai160
ZYE+4G2OPFG6YOoFVg/10YHDN0qQOzgj1NgIBfl6kfnXZuwyxljm1f+364vBlGsulrnpuE/vdiDs
lDnYXHQR85LTPp3MaFH0Wpdn9hnk/nUhUbmN1FJKDDDngy641qOH5wGM02F0WaaMtZBL8xAasqST
lijn/qocG54pDQP02syVg2bI9Kc6vcy2Zz4YxjcMZGhrko81RiVnnkiTlf5Ak1E5HJLihJtrwfWZ
kIaqiwpNVCiii5YxhBWn/K2c/shzEe2MXuaAB19yeXevYECq/LQjfsKDVM2qV5eEIQPLkcyTFEkW
AMSkNoH2OJfqxk2T23vmmZSrIrF8RGWaes/gUM4ZBKXMK2DsDpnoWKIRrmzxqQ6aYE9T4Xr6iaI2
JNkAvgxrS0+BN1gozVSggtVfLig63UTUe3tD0u9ikgOhw5Xp2njtA0hG2Is5uwAFVbmiJE6LbB1J
Pwc4CTMGyFcDViHmH3KYfmMQ5zQI/A2qk9b7mA+zntPoMaUFxl98G5qGv39FcvKwYISx5WTwhJ9E
DFfJZZhQPPJO5FM587njXwrktVxQNlypTIhWAeWCE7ybuwxHzhpn0ZUk26K1j4W50QzQOYa1rAmK
q33cadhvEQ+7TVD8y6jqki/7e/DSZpDiY/RkrFHjR1Vm0RboscYNnk1g4gXaeFovga91V8Dvklur
bV0QrxaPDBgpNjKDjm2Ac08U9X2XhF+DAjM7fKscqGaVN1B/Aw5GkC4PKpH4/Hgd4U6ikxdN0+Kb
tfoONfFtN+GDBDUz4bk3EZdolebMxhrclG+h6PoqGWdaJcKW/TKDyRluPxCavUzvFzEA4hWqkzWx
/WRi3PYcFNT4NXRNyH0CrjThA9l+sFpl904zfZSnR2n19ugDKe9RlUGjkwW0hfuGJU+SJ4cF+ZSU
scRak9dg1aeT55FV3e6O7mwtwja9XZV+XwoSLERrLJvKL8WoIOs/KfXwFD0AizFQffHOZqWcr59h
GVKyrdtbUYQKgdT/CzSt6xjGZaFDTYYt9tohBHmcNNMWtQm3/QivsiOHh9A+dG6fExzjgWDWeTfE
uXmQqjhXOGyutkaHfxtgp4qSziIK9ICqmM6we57cCVoBC/OM8pKjR9/0/qWdPDnQqSla9cwAoCvt
5Zlm2ChYuLDNA5mVZ96aaPM5DkMEr4AS/tp5z6peAz+C4ZP7f5QNGYCyPibV9IajvkPghfrKMmFl
zdNnuvgqKo6hvdpu6mmRjypOYiTOndHSj4p7FRhp+AqXYUNRN9DqJ+MJa+sopQeFFhOQtInghmLE
LRuY1ScxFcvOAzOHObIYVPFjC0nh9rr8lgqxSxyn7/HZtYnz36dv9+Sw5LAkw6SIY3AyBB8wE70E
31E+VS/qCqNOXuFhH2zXx287Hbqfsu3g4CU/Ub07cDfO3Am45tYI85s5OFyFM9fO/wCDPcd1ioW2
R1kT05SiFKUvcx82fX7HtkclOaOC5VwxG2p1kgQ39DaJvZ9TZ0FY5/W1zxrER6w9YEfPdCZjALmb
SIIxw/f2p8lPLz2c3zkJCIIdxM2C8eFTzadqXl6EWPAj5lFpTGM68Y95mktO86qZwkUMDGC6mko0
3ko1hCVjM4vK+nawJ2APN4AkfFn8E6pP8B/PeI7zJNj7o75j1PahEMrpffDngIFUcPfMdWUf82X2
0nPsw7E/FxSwUxFNLn6x8uJcYuicIJjh6vCb/jNyruAQE4QSn2cTAjkxZHCKu3EKq0HfJhqrPHPq
dsM4iK/cVNwDqnZsR0tittCoFc3RDMmR8yWLX3sMuNoJAyLwoBzoT1hwgQ64WkolHfVZ8C2dzzar
aJM5t9npX4Z2KN6R0YRFtXV260RjhmqWbLn2a8ipRS96MndL7IygvfyVB12OByEU/lUQzCYKkBKm
EYCoTrNuTlj9za79LJD0LVSKgAw4YpJLdc7vL3XVIeABjGRyEnXmfYSUFthgIRtvI4d/BJbJsRFr
gwgg/FPa3QQuhOpDP3/ZTW8/An0okJRfVZ2Vi4CZc+HQDdibueycZh2kTU4RT7cQohbo9shyE6Zv
U2wIsL8LX6xkHur2rBRdFwAYdmUDShuwSLHgo6HWL65pAYJVQGIfLct4SILPtO0ydSd+38o6uQus
UiFNgJMFkMeOq64hLe3TBkgqwynC5hxzZWlAvCt7MybW1SHa3Eltv4kSIpe22UnrhtiTQ1WWEoPl
hIYI8erT3fhzLxD0ip3bPquuCtUACeqpjkzncr6ovFAKsnq7kpd1wysMUxwUtoEtersWhmkE8urE
FurUOUulB97dlV1e3CY/xQbicWT8E4M3VplQw4l501a32BkE1zDffO/Wndaka5DXQQ5DcJvPH7lP
6Ikkqy3eF/yMIHDa6IemRgFD49OFxVrdZ7P0jTyDsJyCAkypUCOZ+an2zq9kfzz65MOzBOUQI4lk
BgqFKcDofMaLsaic+tqmahYRJl5Vv/pTQhQekNeECbehaLzCBKamti9mVc5/SPx/oK6ft/Dw/l6u
Ag9Pg9JZlqLi9GdINYg7gNhZZlStpChQGDfgfe9oX7wIwjkB1E2wpnAizRIYfsLHhlzJqKPLyF9/
J3kpzzeGJ+yrfOIcqKtySDyl78JfSoEJPHDlgdEQe5WUSvceQkiX5lhAZjvXH0bUdbqsrWKsUdgI
Xr7gmwaxr1PSKiPmLjlGpYRqrX1v8rDGj3bLry9VkuQSEEpK3yQ8JYbpzn8dYj5U/ljaQIWoYv4D
dt1jPi5kaCTOvTwuZrPmnhwAeTjEuXIUEnPshn/BJGEagN6vn1QI/zoBG1fJS/Odyq1neSBmwaEG
3liNC11J1YPOcBcZjbvsPiyQGsySodqKMMmTupp2IhbfvHSbg3arKsnfzeJ/ciLastnm+uA/Te3+
8iFkMrconvrfw2nURL0fwRZi+p488DVL3H+CpJx6DpXXDg0IsXRuXetJFNMtgIw1pbQ0RbdkU/06
JaOgRDUCcgkHkgkAYGxI/0Ty8ZwvA62aY4Nd+opzLt5G6o0vbcHHq9JsV4QoX6ihZ+xIw8HINXrb
IHxpgs1NUwmFVzBBxCBAhvgjCklGtd9b7E3nsxpP1r6VGv6AGaTa3S0h3vh5pSTyr/QTEHcotMx0
7m75RyaDHGA1ZMjKpCtWzPTPGy9RTW7reYtEkbQeXeO5hnJtA4tGz7ZrSX5CrjINTshNrg5lGzbq
398O1uqEN2/BxXTxehtryHMbnoBdam5YH8KjWtyw5RcgROZRc4eP3G5UOpYViy4YMLiQPiPuTuL0
+tn7HzouL51eHrEKgMcvGrY/9k+BoLR6je8FKmzYYEtsqUXsqOpNLVTUi7IVlmD1WH4Whi+CRLzm
CYYkTa43s90B+QY+YmgICbWPneHqkIFNMOUsVKcOg2ZSfhL9M5mrEptHmvkXmosYcsmP0lBURa9G
aINZLfZEQyBDK/uGLeDtxV4flXGnqN4nnqy1Z6MSv/OQf3qbNRo7luBLMzQky5F/ZQsIxy0czvvR
NwHUUjNchPt5GI0n2b80GSeW8MbEvXBlJB5FnJwP2nHhtDMgmOfcSl9RV0f1tjfRF+PlG9LUPBOm
dkuqiWorCeNkwcY8cDfhpla9BfqZZ0/3Kmts2P3zwDOOiKA/C3U1ESMAQVjrmH7boNK0lONn6I30
W9wgqhFM/iEBNUxlKic3QsN4hVe925OZGuTEBs5Z3eoNSeu+2UijZZ1PE69UTMjDE5ToXx948Dv6
UHxpvhaen7R/kXT7282aAVVckT+i4CpyBkLiGe2E1jb5JDdYsWOiVGLyFMJlQHsNxTBMnEqmDdqS
0ufxIcbkkTjmNb1zAzNvO/R0AjX09Rb+KDe70riu9EAGz2Mi9k0Ef/jOSB4eRkRvNqttaB01h1NG
mCo2TEug7AwcvwAqU9YCEGHQgQkDSR8mYQw66i72eiNEV1fUcpIVDIvbAUa0g/naoel/sB7/xOEG
aa5y/tgUPX1QOMUnyw7HBVvmQlcnHww7d60Qrvo9pAAHmDoPuhmES1zK9vPFXGHHm3OsCEiw/kSO
09FL4dnqO2ngWNJNx6Cspgsw/Mg76vKOMWiXpkHjJNc5EIISU9ebgOVo1cWKy5RRpT27QDvCG+Ck
XZ+BR5ye3bcsNvCNZ/niO8OUeV+XMuqAbrb3pKosRUDAudCysRJvFVHC+LfOg5Cfji4CIiRh562M
YTAXLhCAI27oG0gsqwew5taDsgiAkt0Xd7ZmAGaP+HH/pQt+N3j3NyaZ5HUfVnzG4TPfIS9L4itj
DfOHh1ScsqRWEhrNhFVL485ujGvougoHoEsJl6LBzd3IVcpzb10o0wY1rnbOrTwV8uBMVRUUgsdW
WSELySw+MZOtiCgost/61eB5FfQ0O75FIodItlavfv7kZ9SNSuCC6IyWZlbcCyPwXFweI6CYXtH7
/f4eTJp+0t+3ISkekE0ZGU38eO+plF23jM9qXuroSFk7B3tYGYCcQRX6Zvsf2bN00hqRq2zgerzB
YF2xlmxSHRuc8LBhBQecmVPVz5hgYqtrTi6R20uoS5l+5Is+qlmYdQrbcslacXcxn9Mt8NSZL7PM
z+pPT45mGB0lT2DJJY2V06Vd7bgbikhS1CgUKy0aDvCsf0uqO3jUL9bpIGNXC8PUBPjqkSNTcnf9
eQGgzAJDCPMM1JGguefb4XMOtsDOG1QVTTTUrZOI0p0+fo0v0Lpoe6jUAKS8UErvtvJ3Pv6ith0z
1GfH16Civd6LIAZj7CgtXcFdBOjaIA2SEEZj3mN9qkXfS7ahXTUSawU5aNy01blrgjHxlQFlfNv2
wUHFlDaWDjoWlQxHQr/N1ElIk1NrCbUkkrY0UWWwoCliHdiwy7FvQDmtJMBWsPlNBByLve88VrIp
J/5zFGOL4OSrCL+MveNTB0/ZxflopeudCDJukyOq71diHMrKTFNSPdWkYL/DZlh6q62NMyzKvfq+
8DiMRnxw0iEqDNcGmkuDUy5C74IyOhbCFvykDIEy9zzbLJGhF1UOSHSRmdRHiyx/jyT3guJ7DvYl
+Sewuu8vjk7fqca3i3UqosXh8AXf5blCHqj0acBlFbnguc3nXSZM7OUAtfaHtZjKneJKe9EZ3JEd
iX5SvHFzcOGU9mLpErATyLX5H3OeV7TAbJKe+4YNsq+AR2CQZAiziJZC+P0kzXroGETrWSvhcDOT
rbZMnhMiIXignXeaYBCdO3cWtZfcMx7AcCuPyQt7sHpMSDArhOW4YW8++e4DyuT8Qj62W0SItMT8
hRYtM/eNvKxPGvUD0LR6qHicL8KXvNhWcMG1D0ei/GkB22QL+YjGI0sA4a5Ogg64q9ivl/EMo5NG
U9cf9zdQXcfgKJobN2vlVPRJLWVPj3bgdYXePscLkJTKuvjuXzq8iKcGyb6M/Qf/aeP80Jhxit5x
R0LMaz2w/JxAoogGjXXL04AVEjVWJXPdQ6Lg2Oakt9Jlj2TuZQL+vbteoxkmVOu0+u2Ku/yBOy+2
doUzTHtnYqAZVXKSQrdj416jr+i0acQ/nGcrntgsgW+y7vbOtayQ4BUOhNPU+VttPdCgao3OYcB6
PnYQW228+pmjs+MXx4Rd4ZkZqQr+YN1hsbK5ycGww4aQDMWho9efK4CA8MBlHv7lMWN7lsxD1LhT
phYE1ACv8rn3aAtad+7DwGqvdPqyzwar46YkEg7wgicDlgBoA168c/YNaNHQSQa9di6liNPUOAin
a0nFzQrdB9xcNNGHcZ6Y7SwCn8GAVLzqvc6KNl7rIQPV3RFvreNhFa6AV9ii96eKBL1ChPGb8U8T
8HNnp3BJ6L4zWq/W/OfTIsmVSDBU6mEaIHFFkVFt9qxMnaRj2tZhxtYHvQ4VSn4TMxyH7SRTpDN8
rroeZZjupH38Thuphkbe0uYSWFbpllylb/qJZolPIhNIVuif4do+JRM1hAt4xTku2EUv/27NbA4U
/pV4t99w/Yij9cVrX+s0AkQbvv5PYd8/jWP2ZJ+As1cXcu+zufF6TTRvbiiAGqlkiktWzGRpPJwh
KQ+jXadOQFmXQAjimreW4athqXGNf6ksBOl7Ysj36FHtqyWUKLOxRCE8TCjsVGmEXEi5jRuf18XA
+mQy9HtvFfRKbacEja+iRXRWNMvSFZ0N7MqkGoQ4dxRzeCRj1I7x/NQHNH7Qwx6/U6isNDKXHgOd
cwBoOv2I5Te8M0ahCYOqNX87qkzb2eJ0rox+9n6MwqjDzqr8qt9y+E+BiEHw7ROXwbJKR+swgldx
3FgePU1/JDXJqTnItTRIjADPg+NljSUeQv6q4nK7aIL/IvSGXq12vjJy7PXNdZNTzDlRBLd2Jvmd
4DATKsG+tGj1XmC4BUlM+z816ujtuDFNY8vBELM2SSFnFdjTka/3XolqcDtTInYO+qIZGHTyGJEF
PbNjBqsg8KSRqLpB34EWT2c66thyB7ZO8ZzVQ+U/82cMi2QgvqznSA0Tu8ymkm+uFMlH5cyIGQgK
SAm06XhdKJmCb4rtG6PEZe1jfcsNC9EU908QP8lChmI/hoWj9hKL+dHQyWXPPxsj7q63FNI1a7CV
HaAvPTfCCCGZJqz7xwwFNjiLyZ5wTOSIXGC1o38chon4rC5DZLwhOEvdhPyoD3xAf+2TSsa8krnH
mSu8BXJasw1KTkLFGiTyzHuMrudQQpGi58Bo4PN1svD3BGy8MqEZfJOIxpNsVkfnDeShD+X24Y5F
sBk3msPfRveWlgSIa+N3ixV2dBUDKBM2amMhNWfKvyyaTgC1NiilVgA7bGqQ7WkYbusznvdgfdtX
RJiYdRMyMmY40V4BO9PNIVG1ML9G6SaYEgqwH1HoX/ByNg8fe9KTP1RnGlG/b1pKU1OWd2d1ZdvV
TroE9sHXdHEhGbCMc4CzwQ0c+o3ZYH8JHtWSQlE+2GCOmUUgTfPfCWqIABLUE8LAuff89bb/EbA1
ZVxHSA3gOxjGSWT+TO+7eCxixUe2EJNHkdEU9Iv4OImi51GAwaw6HTHv3/lIUt+Gy71N8N5/OFBl
tQrUCu3ghAPQv5m0a9UC1u6KXRJCfGDK70FP8EaYOoI9aIR6hSsjtCd8dcuAF3svWKzf/O6Aq8c0
YZlYdR8c2KPPSRyTiKszX1yPaBjXlcbO0ArS8YARX13H9M8tikWDa0zASap47RB/dvaoC+08IgO+
k/x6JVohxyGE2T2A5B5wULhRXPnc5hEh3eec5a8W2Lk4VPN1Fl0PfFcyBs3nblxuDXyHFV3njQPV
n8wtZkyCxtKeBO8mIUq/u5WzY/8lUNIK9Y1sGmONG8Qeo+W2x3MNuu+gD5yq1u8rjzVV4gGXsflq
pF+KDcTZYjktPFBN2MMqngrUeUfc8xA8tsppY1H9E67Bj4ZlXggGLb1VABIrRVctWrlrsSTEareJ
kSaruT1GqjESWSFK3TqFGRGWX1uz1icci9Jc8OPOhSIOE2ZyionPnet0J7hbKZVPfO1r43baH94z
53orXe1E71rohGJkb0oPN5bMUHE/NskdlKuGXOj3TaTVItoFqg9Akap4sAJpO85skpvcDYgoYKDV
ZvQpIKDhkxVmxsycNB5FSLvcjIYAWMn0//soV4Wvb3+zXGPMYS+4fHW1cFMizPX0z2kwVdGUVjYj
6SrezFlWLscRAQkVA6PDvJvCfRnqsSqp12i0ewWWQTzKA9IXS0J8OAlSx+ktSde1zF5ObODtHHaM
SMx21Tq01Zg+IGDn/eTNuuIlkJY0gtBLdIUybCCmP/VO6Zh7dAXh/sQpNOxbXV5XNLQu8dzYHrti
XsHnFDG3sUm/EjD1qSeaaWOs0/LscraCSAYxQcWO7iphxJCJuwW35Zz++xOZvVtmcKa25ZeZMRMD
20Sf61R5F9KrvB6INdfrn+zaQkOcok77axbIVD4OFOFi8AslS6YVIpmzU85auieiNzZhP6Rq1J/h
mF1R6hmvXmZGjzs1/PiO7T9Ty2Co5R5JddXKhCRGHnSaKhJ3YbYAUHMULiBzVvEyKjeDdhOecahm
fc3+VfHvCJA1eYbeOCXgHETMfASFrf/lPWFExze547luN/kD6iXpyt9cR0XCoquhMzBH6ed/tTgf
UPnYlMy0ZvM9AZogoaqtr2YGWsAEJzzWyYevS2t2X7NsvYSVS1FgQMHvfydE2flkici2wyZoS4nr
JS6/+jAMgDMJuNI9gemlJG9gDStV+Zn7961huWlXsEHQ3TRCC3itAslgYwkrRRIbm9HTohb/Ifk9
qCUqPLQ3y+COWtRjI/2aE8w4C9cTmu65j2SRovR4aDpavA5/LUDF34BCDH7tYniugbpdpalUG1Gq
PmMqE62460qvz+PiYxakhnvjuWUNSAfcK3529CdbeJQ8SHUf/EDoLVbkMsYwpYjwE+EZcbOzts9r
oImf7Xo0ivxD/ipLcCtsIHtW4sV/4ahZA8PYIbLPTudMb6+XDjR2jyOSmLoNUGAuUtqMqLYSziY9
F65luKtKh6lrg2ZznVptw4fpNrLtjs3UIHZUJ1pJCxfN3kJibJSogwa3y+/Xp2ePmogjT9wpHmrb
7aCahme5OVSOmxbo6VUlqTMaVgiu77UFGsnDFfQ3sne8K/g6j5phb3cf4kqdymt5iUwf9xvoiZRF
G/kMFMAQD+lbErewSQc0Zl2DD8iR9qbOiqQqh5rhWqo147fCnbIuW65bIXSTIEnPZfowDIPjUPAe
nojlW+IqDW1cPORpT+xhB5N/Hx8owNMUA0maS1ItraB+sKH2TW1uF/ZMHnhj5e6PZHIFcLwYai4D
Av5rfO7aQSA40TmiU4VYUxi30OQTnoZw7VPPr2qWtqe62CIlyQU7bAgvFrWk/IXuIm/7nz2yUmzu
SrhUQ1yEEWDEOdE0AT1UTgvf43LveZEw+vMwN0hwoGBJKWo8ud/XTqU68PBvf1ndKb+9MwcYm2/n
pWiZ2L0vIXxlTVKWLSQ1VWUnJyCmJpvDfEOX5GtJYVOGgSlnDFVtCVA6Rtf9XSwxGpKm3Y/+bdAO
dLuNA+IDcM5ilOG8pfMj7Zr7GefphCS6tZVU4g5kA6L1JRbOUvL3+wwQRtOct2onbcBujC19T09/
aPFfWOuZ+77M8XD8xiaAj9SqkxS/HMW+VNbRmz2D+tAOL3y+rznZ/sH6EAp+9DVR0a1jkJ4cjPrC
SclJ5sVpeqjjHDgswLfsgg7tReoL4ebBnEs2A7j7kygVVBBm+UH+1aOtesABHQ4sEYEu1R+Iy5Vb
CozJ6kE/YHhKTRlqP5MgodExAQS3XFJg6qg20D8/mOZoLn030TsrMYDA1QP7zY6olSLMTMWNR3To
W7V7nJXVaJC0dE1bUTCqwJQ1dfLP9fs3vl+m1J2BQX6GtqQBGSTsm4b+H3hreWsh3tDNQtocMNEa
k0rvNqw56wKUk2+/wyYCpIkxlfLQIoW8ddG0MtZCo+edaWWOg5bHl7aB6VgafzyKIvrBLFh9EK26
0a04fQUL53A7/KS5S9LUbZXkmPi2/fKZ/gRH3OUh8EZNky0on5+mTkO6Kc4hMm9G8afeW79vzSOU
hD5k8NgtYeus7DAABOq5EpnW4u6YNJR8ccat9wWj7ZLgb7AGqpp4tSalYDjaNZ9QWUvLApKPboVt
xf1fKT7o02nhP32L68Pj1spe+mwomzD5Zg+68TdBKUHVp3y/JZF++u5A7WYaY1k2ddduCvA6W3TK
RXdAtnhW7TWHhsqcnhJlRO13v7M6fLpcTpNTtXBEt4+m5h0XShThQpe/HWULKgk2f+Ip04TzND5a
dZQedQynSiz7tVvBp0bvNHFQVyi4oGYSeggzJSR/FVfdoCs+m4TngftzJ+MsRd2Oij3pEcJeslzE
v36PD38jAobniY2Gm334CFFYQvvbZ8vojwu5nUfZd8xpfE6vmQnuCyIlbbDyY35FwTTZxugBwnRi
CdtdistyEFAsDq1BGAQFxLtxeraGo3q+imTqGMsmPiCr/sidPQ0MtYrGPPl50hHEHW8SSo0P35b8
Q6FFw0kpT1H9NUdmx4jkpv8hKivYsGBl/77tjIjj9XwzFTxdEmZqRo7fLxsKw4tynWxBl84bd0wy
ehhWE4LUpaIud4x3nc0shKzQQUuMDqyEqkratkN3TCCpOlCW9Xn/RxqNZqbmTgKpSFbdw0eJo1C0
U/jFCaqeP85RX9n6QpNTdtQhZv5Kp7HfaxpbH+0Ym5TmPfn03+MwOdN4DFNPJHYEX5GgpTvyWtJB
gJZVy6qJIW4UeKYaaV+9FMB4gG3H70dHoNilqZaMxOnk2cc/dVpS61c6PLNAREmZalRmyNgtxBYM
ngEbYAqHxDs1tg4h3JqU+KtbK9UxgYOXNw4wklw5h4PlrUwDjGkFmHrEu60QdNx3LUxzxF69hgl5
bkiEJnEpe43TlMaeLunBAIJtZYKye9oKr2WCyFUK3IX9xRAyNCsIuIrhxetXenbn1yubmeBoWkkz
xu330UjTtpRCn9qsO9T9EEVraDNU5mNF9lXmDU4YrcQItqVdsKds4QENCgelXcCSsvKEEoxKGIhT
L8Q1cxqFeQPTPrOfnQtoTxeOQXx69XjsYvMwoSJ9vu1LtRYaf9K5KDhAO86QZ9L3oSUHuwHV2v9k
053YfHhodZzm8iWbGtTTztf1inJ0HdnPTbsvyq3KpJhp1w/V7JAnCFx8CtyCamBoiiFHPJ1HJLS1
4ctF0yDh3l7rDh/r07eGVKdY4ijvyQ4ExsM/Wfer7CmYIBQFq0+GVySsIoavnV1kYkiRf3/vLTy/
F05Iqc69d5YtQ/vw7gDxHFRYI/T97LJQxlIDmRA2yq8cTwE8KnQYaEJoNk3GAZAVLBRFdLNwAlhI
BG2OZcZHndy12Z5vwuRxYNoe7JzeBpAM0UFmTABdC5TrpB+O+B5lgUWLHP1JYN6HtN9vWaHpf1JM
EWwwbdQEFn/Zny5zmhBIGDWS5hX0ooSAzo1oz5BtAcJ3OLjEh26TUi1XJwfPgigHERs+NQ00+CQr
osSl8DeONU5CWPOYttNeTtMh2RuWmOCHD6izVV9RV854riur8yk4l9rypZHJpCpVqdg8Pg+DNUs/
qPA9OmCh7rJnkJNX4eT5vvZphFziPhZlAbv0yGDuRJBoTLGkQjz38w0LeNnfl01tEX2H6b439o/H
kkxBDv1JSW3ldaHZ/Zg5hFQmofRDjFw5/UXSseBZz+qPi8erxtvhqvevnZNlQLJJjGCNGruUPBHi
cOUXIv69CiCKQxqGEKi3Oh+ssIzp1gkIqlawb6s3WkviKlXKpkaErif1Z6WNXEAmncSNea6VTEta
TVRY/6vXrMmkeVg4npWP95dOPxmCSstcT2++qxz3i6XIyXkamITGNyrJumb9fUhpyyuK6pZBx3Mc
nBsJzvox9+zS6DKkifymWEIk4T0B63CIX7HTWGffAJ61aKPzRbWMKHuO6ICau7/R5iJafkijq2vt
d6wEKZP9cmrhmcxlNtgxm0vnrPEDKGoYlRppUD5tRZqpfy0TaL3UuFw8nbMWQ+VgGHdNwDKePu/S
0cNb3Oh81cgfC3p4NMJrD0HLpJg+LnH6vZ0yTIujY4vMtEVAsR6eZ9daGyMha0K7GTmRnxz37yjs
7DvmathU8886GZ8fejbFZTCvpfXBW/NvIDO4mlaGDaUbpDf/vB3LxNcNPJKswULdvjQgymRRxz/v
Y4f9w8fQfPAay78ICsWZB0BoNLpwnIXoBG746eMD8MRQ45TLmxdvgisLRbmB25QdMmbLqJkL2J/T
1ym7WWFnhXP2QS/OnOJ0w8nDvLqjYIxTnEfLz4o+dsAc97tUa8TJfCTBdIcvaaQMNsnBTX8bcPrl
oR/8KLKAVJJmkEDU57yTfPmW/AIqwC5FXYV0vandKulrxbNvYK/1CCaxufucPSEQFArM8/oGzcvu
TAI8QHbnRBarYGPl76JaNaqC7LUwJlRuJJaA+DqsLdYCTPRATgMrsFmJ9VQ57efk0LXD+gvXdkYx
G/EUVBgHxgXOc4Tgo3fYOi8orWxDZRoSojY+tYP9JjN7T4HNp/SkhZ4xBGhu/pviMTI4mSgsP27H
vi1vtLZmBCJ38TuBnQjbpe6sviF8IN6BsH01iW+fsi0tzEVzr9swtlesA9YhvNVE9SjAxnh6DvVe
TQMToWrm4A4STgSxdJ5pk5VoRifOpIJmkWsY0lcgL4LnAzRTFQO6kYz2MVEOhD7iFS9u4sWdp6lI
MBfFWcV7A2kz0qLq0ec76KUUXEoU/yhnvt47FUrGEUPxiIiMH1t6a4kTShuciC2r6mAtd2OCk2M2
71/Zwo92jm5X8uuD/AxyWN4hujzuYUSBUBocCDIRSjjW6HqEHspubAxIWT5PndSVHRDDQUNEdb/Z
IbSId+L9avmXN/maUq733XEbPytQCQSkpPVpNh6uoPFqQqY+PvLD6Uj3uNZmV8kIxv/LiBxinQf0
WRthMePdRBmBUI/Y45zhVA15D0DlqFUGIwGZ67W70UJD2jPynuwoqwaZ6f3PuGpCOHzm1Li0SBux
U/bg03d2icayKKEqWffaB3n5PrEpkDljh/yqlJlaPYawPCWP3NHCxqaRdPD6/Molt+3ylKpZdxZF
XO1C6FGm9zrJyXy4Y5n1n0XM/woZ43uYGzTVNs2XOoDRPKY818O8SiOLQhedXMylFO5QYPtNb22c
khPctGubFg0Y/pMkbDZeIIT+a/tFEagaptubHcbzoGWU8dlOVZaUANc60BDjoj18UJdQPwMtkvlF
g2ozF9RSv7PSQTz0O/MHx6UETCm9+bmX6zQjT7+B+rncV9UqmDGofNCxFLOVfDgNuIpIVGixXUzz
RY7cLuYM3tEDtWuILF2cKDGbDW6IxcKm++tOuXaHnyPk/bXK0SueIfgrEM1xHe2KH3tE/B/LCNET
gLps8xC1cK0glwtJ+uzE3bTlFmc1gWrDlbPznGGQ64OjnlMPWuh6qBcUA139d3Yh2AE0sgIu10hd
V3tsPrllpqbhDbyIUCrAbr/9CzIjerVhtoIxd7TIipRGZgpCGdra13SBAnL81lBKlryzMGVQ7KKa
xNp1p0cyQz4KJ+kqEYRHniIo7sqMfSwUckmDHscwcE51GBz0h6mS/x63mgMAVH1BqheVjjx2CYDR
nIVy/9DHdSByRC+oRDdAbR/X+LDdX+bycwKdwLCllwlDiaLjR8yZoGhU4QnFxqyjeweTulk3EW/Q
cQCz0RvVqI5WMANRrDYjWQ1Sat2NGYTaersWa+XN6Wsf+iSIJuV1rs4cs0Sv4W+YhLaEHNRf9k+7
FTpzC+Xa8oPV4eECxEXARiFE4GpY99zYyZcPVnflhoJ9l0txVitKEc/SSylFfOqpdD38B96+Mmdu
QWBJCpTryj9sMxJa4dll9iOImvfnJK2T82KJEaqNlYuTRcPGSd50og/LiEhuFzFzVDGSS18U4dpz
BplzsV9RkOLIx1WMU0O6HVYtKZQfg6sYHeMO2lv7j2i0o/VOOKO11H7+kJnVjns6gNty7oQdMQeh
I4IPkXkjsOwOMcUncVBVTce3GapFko4uKkLzSpwAckjR0V13SpMB0RYbTgHDVaBTXMzrmqAAsFIs
f+GgTI3kZGrLZbCVpeFP8sfhmN7qNQ7rHcfjdsESyP0PwR7nrndXOAzMV2/mnxp3QJXcKrcXAOml
u+IlyO96Usw1T+ShtrhoqSmqaW59G+NGJF2gPV3TN4YpD1vJzpje5PAiceVeErkTnl41S+lH7HIO
NWsXweq7bhOmskGz8Lac9RTC8e0TBaNjfYS1EV9dSbsPFXXuWRW3XCIVPd1VKuL/ruj2LXcr0AEz
MSQMRm7iIlQwNIl0Dzz0EeW3vM0cQvvfC43gOMIMGcS+Uctxgp9U+5TR5R+8thi0LrqGtNieUcqR
TJOykfzFG9iBLTvrK10QCtMIY1ZoUqaAH2xap+DpVJjFu+rFZJ16w8+Q0OmQjy1dwNUfSUzW3hwF
Dy37ZOwTjlBt3bgfSzJJKurn8zw+Ue9YrqH1OxGYsUXzpYGgvvqI46Q1/14e5hd1l9sOe9X/u57X
pmq/18QERSFoKNZNQhbl8m2HJM+DScpYLdrWg6Y7268nC8P1D82TXI3LgldZ3kkQZlMR2vImKJ9W
i4GQhiIaE1Tjh2vdSODPi5mE8FCYpnzeTJxQCYpcjgbCYzDB5OoTkrBX2sJzjpBKlhqUaHCRLnk/
u4sX401/E35kcoGtPWlZaHt2P0V5xkxWy+BWGTxBgdaC4/6dF2IOY3P3KhafhYyt3ve3A9OWwY8p
bw8ogbzAJt/KyNMjt6sZClZX6bAwAq6HhHC9E6Wz+ZOWheGE+nnvkTq7nOuR5dky5k/uF3NqlcNj
AGdRO01DY2QH39YzICilVYBJ06AgrQJ/lTGQsbKukYKeD9zkTovB4lFy7A/uSzZx8zGrD81GOqz4
U/ALiIO2JCIftRwapt9D2TrEt9yiV8XrcpV45pnetgVLSH1EvinmvbnrJm2nbM5l9bDstnG58Bt2
YU90YmoYRhfGZ2kj09D26/2bSq+3euIQ3a4TYHTBPz1BmBRysE9t8TUiccQX8ZU3VSb1kCVsKm8w
BgX3vYk2VcpG++2Oz6IaB22h2qMwZ3YRtUisO/P0mpSx1jlGr6Ux/nJP25H102XH8Ff2rRHAXXWx
4QncQyHqQ5B/kvg7XvcgQ9dCjJ0DqV+rBxhV9YhhN2mdwlY7xS9wlo6fA7iaC2Sp4rsqO/S+1dRG
8meqMlrXpZa6di7mbsuKvwh1JQv0XgHM/wMzaDt+nKloLrO40WgbHZhp2BR84lL0oBB3+fDSM02f
pnjk7KrQMf3k88yalgROyaqg3L2E77nxvIOSbLS+OwWt6uc5Uy4V9fA3qQzSYxBtmu8uunnci6CI
um4CCRmsfUFaM38C2/7x4AJEbJ/giyjIfYRoEYdbM6gwCQqXFLy/xUOYP8xPDfsd9VtZBtxcOx4/
6tRHlvrgwtn1FmAwX225NtLfpGhD/jYzuZy72GBedlRTB9tzoDLDPVeHvoNES6OOBD5lhZnFffRd
cOeZufP4ykZty12oGwGpYeI6DiEoGWP1M0rwSSL99fbQfI4RkUEPKtSvRNKVJB5LJlzFaMQciGvH
IJuZhEeLbfcZx2v5IVdR9sxGKRtoE2KpIfEdjuCIwmbDMgpsRqdUmzLzCMWouT3lrQ1UVoqx6XiX
zDcDMRdspPDEACbZnezt3UeAbZm9esZLuW9FNzwmmNnqbAA/t+TLSD8vVVWxnDRu6hO0wrCfeMDX
W4hiVNhl1fn4H+LjUsVh/HExcsMBaekyvUTOctdynt8JqR/yXT4azyZbry9UyI/CdXymHnB5zgh6
c9CzZ1lqQyowcwuCOjXfnFeh/8Vinpln0zRvZleHh5egvLbgE1STTspuNJkWJpVMZNf8WjH3+WrA
O1gtBL994+m1SMAw2x08EEiE9SsGzHspU5i99vofYq3s8VUGsBKTCDHARRMJE5uR3hysi9BDTkz6
qNuWe0phaASHLBUK0VqP3x90xt9YDu1+AMRYfsW+8WdDdKT9fWyjSBfHiagyr8CZV988E9wG9ex1
yPF1+3qpj59zdtkQarvQT5FWvuwkRiKSioN3+FhfxlaZI/SOFkv5kL08v/rw9fVoz6IvSxCBsQme
snjBodcBPudR3QMS8LG8Lz/4nqeDdgOjJpEUPmS8yzBEmYHKPoGxSjOk2e7DQoCByBlIESzcSu2Z
kj7qqFWvhVc064TqazYTkwXm8wgpU9rVuH64DMkf8vNzl5q5I4cbbeuTYvFcxqzR/q7P3HjA1hpq
cqaedGMiP56sKKDgIy4xQodqDfXwbd5PKEdMpksLGX/1kCJr5BdoaGIje6FOwyn4WM1pEfCgQGky
+NFVsmvSABQTtyfSgX33IgmVHg3gRFfB46qmZgOPD4Vf9xLh62avcpLBW6W5PgCiWZ55sTHRLf0D
niyNmrVOchkO775Khp4dWCXagkM67zLj8vbp/ZebsKOkoChegG/g/IdshcQuwGDecb1ZAUbO1ZFq
TXxvyoo264Kn7P3WtEHeGhv/iTFZD3gC4U2PNonf5i8yyevE2IsNCcaUYBBvuJ+ruklpeeXmACYZ
/YKSBAxlJJcMTONLwfasLdyNQBCgf+Z/mB16EaVu2+kYsrsJ8y36D181bmM/GTKAhZfOtJI58Pde
oGtLzpQYfj7davHFCIVFEwP2ceeEbUjbVnCQdh0PQjLSWY7fX60IyazTTtgl0sZI25s8ek1wRVyS
BaoidLzv5LeGc7/yK9kdmx0+5kbAhPgB7mgHaVYVRQ0JCYWrSP6CTXpLRqadz/WoBkLJHHRBYXbV
JEkhtjYTT2K0yy0hzJJM1JoVv3Q1PC+Ep1KsCCfX3J4Q/+NxC9cqjSDYBRID/0TMiUmZbgIYhCpp
w3GPB/O316XFh4YlJVVhrJ5OUW6E0k7RXKi9qvKodm6gfzPwFWKFinES72KFjd0XERAn/hLMttZL
ViIfmHmDScGXgv3kUAXzJaNzJo29/q8P9oyjtmZfOntAfcc59+1lo0ERa7/9DTiT7hJlzNl04DTV
9LB4oDr5qoX7nl8cJaw4dkr6PiJfPOdS34juriau2gqMZlVMTYodVbh3UUepQ8CJqwpM4Ir8FTX5
muFBQFkAmgLVT/zmOANF3vGKr9WE09xRtP+18LCwYvNrxg1YBQrX9p2gZ99P8WVwfSXHhFeUQldU
7x4COWVDMiB9vpxVyPFPBGqc09RFYHH6CcXR8RCcvXiMWYtwZ6KctHym6nPtOiK/Ab9zHZshj6gs
dxU9AoDB3As/CfUuKIjENBI56LCbmxDEsvix1qB9mVHB3bJXUIM4mFzeCmWLe3fXo+hPOiTsmDk6
FCTu2o9OjEDf2R2xN9Y7i+boU/ZZXJfS4PwjqMqZ/Aki5ilKU/0ULH0Ezv0DAlXbpXbxIAySeV9G
+8Xlq4qVa5cquIM84wURNpOTSYJKNqO67N/+bcoklDyili2WLP4rdb3uBMVi8iWOOnPdpFB2sZyL
sJ0CMCwcrHKFaq4aAdoRx5lmUnhsAeGDaYo1s8Oq9JpFenFxWGteQR6GqkPod/d0RCE8nK+mHYZ3
yK/TXwOFsGfFgAGX9JnL0F/TvKjpFzRBWTyzOXWVaP66+F5WAFyCFnExHxAVcCCSsqakcAm72Nsc
FC/dMXMxFgBYjt8nU4NXwMIl2blF5AhY2DIqxtBixCg00fwIIDCiF2S5OWYplHrZwiU/P0i1KYb0
rJESvA55eEJGAzK+lEt1u2NzJIm9hQlglxvUP26BL4QBK/DFEE1YrSduSfHdcxOiobM0p4+LdrlR
yrzcTBzZOPyj9/nMt3+xe+xyG4gGcGLYqStGf79KltPU/6NGE9aJwG6TRifqz3WLHlp4KONKcch2
lf+O8FpkwScO3g5LxZuOEWKPp9qEsQKhCGyfB8iDPOr0sCu7sakaG085LGdUlcwxNrOYiNTVfTwg
rJysSt6reAVfyf9jPe6PrcAyQ0eA+6/R55RIzrhxYYojlq9k6pMuiiFxgdO9p2s7vxmwPyDHoatA
nDALWb4DDLrKvXfdkOt+55hPtdrmd/wPaH98W1Ug/e9bGCMPfRtQTistDGNnB8BzrxQyv1+2ta3w
fL13K8gahXD9/X0fYrDEZpBTuM4rW7GUQdbuS7GKoGYaKD/AXFVBBto8L6a8Dajq5Y+QLy2TWcxg
hirP71IgSEgyOXVuClwt3xn+wBCB9I5H0fngVOGCrS6tRNfZXyhIlCdyyu/6TxM1QOcKUobYXnOS
7YTSzfz369xid+Q5uzUN3c1DtVlmPK1u82X7Aqc9acFyQQEUhlykj6J8PyHr5cJXn++BimWcnTZS
xrZ8ey7tRetSuUvL7GjdX93HKeRnPh9jy9WcAwQO7BHtVpTSo3UGzz8Pw/pvcxBLyJVuY90W5UVl
NzjJVOO3QX1ffSnZxM9MSjYyek2FTIKfVJuB7FmBPiI7LfFu3FCOwg2SPe5++CdnIbeAaTsn3oFl
DAl7KBfVikv/uxHOdz5dGS71XX4JuUWtSxWLj8nb3llpw5IYmP24vi6BBwEE8+c4Df9WGihQdYzE
w00qagN4zBuDmjnwR1WMZqGojr+HrB1S/s4E2YYQorktbn+4Ymi+4eBbXsQAvUKO0C19Nw9Xfw7s
9AcFC9s5dUWb+wjApfVy8dBOBahcDmtY5QxH4PWHqZa30AXuXzwPvcrOFCLqqP9xIay34W2bmkFm
gg3kYJZz2hZDCZQ0r8dPB0BQrWcVOcmyy+bWdHw7AuRDzpdGUDb6t4XhOEWqgYxJrMjZkIHqBg7v
ia3k5K4Y8LF3DdimyYPTvBKWm/0TGRiGWkkOkTJHt/mvgUNMMuzVHmGMCAkf+g1c/b26W+ti5epu
X1YCpFn7+GRJzNtJhUF+I8wkl9aS/7A4q2r3ms9cXHjr8il78TQnjzbXx0sEodVGMsXvWVQOgk+h
sc66k3OuQM6qaQpp+gWDHmp+DjL37Ayu3WKbtOeWjmODGeZlQLqayk0kb4W/ro5gFMn8hUiYS1Mj
CbdEnTHe1fNpVYlebw26tqLylVFpF2uOUFbXC0+jOCJaVzgOhjyed35zz+OEimclZuT4NrXNc6MD
SSXWEUKfKrYNEg4nNS+aWhbphIcF3jG7m4DHV+I2G21hHXmZOAHlVPzE4/RP6f+SEiH5wSSr5iSV
LiW4cUT68Vw+9YbwjvY4y1wP0BaQR3twIKI/gWCtZcIbxhMYqWOA9L9eRRCtHVuAc7V04qj2tIuw
zPUd3u14jr7KPSr3YZnzb/ms6p2XshujtF3Vfms5GGsJo178UUn2jzKkKEN1qOiSvJcutUjJAQU/
nhK42sU2vj02M5OwOeUMOsFktGm+T7/u8SJZf2QxLL61dgCOEjaM6yjRsADDc8emLPF+5NU4gisY
+/3ETwRDKy7dB91xpa9tCeTNEmQXJcPcaYi0dCE9OqooDvqDG0/Kf5+5PZEvuBGai2ctMV7TrpZ6
fj7/32zxHOj1CrF3iWOx+09lSW4Wt1E47EWGZt/NPLS9OoWgAvHn2AKA+MfTQRc7OPZLlKnuDSmP
JBFjANdMyc9zkhUb0qThE6pOA/FiNfxZg1K9mf9NFyIFcdiKNZouFq1usCjlBdOrY0z4pvCrYIhl
vJ4bvwNtiDIUbdumDFOYx3mxaBjzxycHJP9Zr9tGuNsX2hx9CteXnhPmsmeATXllFJm3oi+Kggfz
sA96vMTYRc7VcK+2XsaAq6bF/R2mfjRII1j1NgSbngEIP6Uk1QzOvjUBCNvDqOUqSIRecgbcth23
i10qjODvHuzL1F+edFfdJytftni7t69zrKPbIQdmfy9XJVL+Y45o8jO1o5yg0EQ8m11FoxwStCQX
TR/OZoB6Hx5+JCW4fz9fy1xeXtUtmzRMDzTtlbCoSnDAf1u5fCG7SfzKbUVoOio7WaMKCJUuB9qK
yIGO42N0lpuVfo1uUPd2vBgyK3hXVbvUb4Ey0XA6j2wJdA+dns6uumYsseu0E1KTmBjKyZ/s8fz7
nOLY1pW037YFAfFE4HunicLh1PaKilxlrLsaTkj0W7SnWW93xeaRuAsqeM7e0UD86EOkrSHOEvpK
2gt/IwSzXGyQgYKfUM9FAxRHoOgicWfIFiPbLXhVeGpwVPXtXlHFh+H9AjnzyQ2ryW7qXaH9v3nJ
ew81/ft1E6AL6hvvX94DIdqb/B0R0W1DpMCDeBLfpFde2z9AVfTEGiNTzm6imyBt3dG1Wqr8d0cC
hSI/9cYqPSgk+XLAIEnayndO0ZoXVntcTAYszz+xIkf+ksOYT86Jt/xwRVpwi/Jg7Rnf556Jc7Td
Vcqr/2I6YD936NojpO/lqLoaLdobcEHKMFW2gPbmLIX51uAyw9UOu9Yqn72lWOedt5UIThE6YvIH
jPeLK60ooGYEEeP2LTwIveVMp3BlnJxlrnVIBQuWCGnGS8admGl7xBvv7CYwQ6nvktK1nqHJJTUe
CramJo17WQ1AnHbMKzTqP9sBk7CS/aiVRUIbuyJrveez3Fdr19pLkasVPrFrAIldmC3AcZgYTfzL
Z6FRFm8PelpCQks4orFNlzqvqLuY/U7E6CP5j9SBALwKn7r0GsOv3dsaT2/AONP1parYq6eJBGvz
vcy/jd7OnwqgWr0n10DRVmhXE9Zkt1BV1jGFqvPDyGc+IddqtvYiS1hmw1jw7FEzJRfj/f5Jj5ey
zILrOpXOwbZ0AIzYkPFexXKjoP5y/KoDvGKs20KU3kt4/4yExuaUl/HoUvwQSWv9WWpHHa3KShI4
q3oxY7ahbWVj9go4B3gz2k8itsFWzLecigX3oSrlxjC6dkEmU1YmBafbzv3whCLCLZ2b5Q1NfjQw
3/9Fs5md+eK8Cp9f8ZVGzsp/TR4gf0k7x1k7vzTifiYaQaQoQHKdPUwMkdm+FtqdYsjUVjTWg0v8
v+iKFmsG2fma44Fp9R/Cmq/hjdGojGfiewbvGLJ9eGFsD90I+eSwndVUM8LQnL8w0FBUhOe6jioF
uegtokXjUIi+NO9chjd4ase7sBpO5/cH9cvVufXOgpK6pjFeCZ8YYFBDLa5y93+A9TpKdTFmSL2W
zXXzwtivWek2aGyQodcjt7SrTXXlqU5W1VEMG1uKJ+7PFUo0IFpDsc5v2cJ4B3PgZoileTX4QXl7
O3E9daVyhJ/AQmqvY77Tshq9tRDx28VkD1gyVIwAeQo8W8cugMKYS4Qtni0ZUkWUHwNBdZ55q+CT
mf1ZYNLVwbGs6KcWh/wsruVtkG66KyH3jgletY0oLGL+xxgpG9Aq48nRHRZfLGTX5XQfm16VSieu
AupGo+B9/GkxlPl8Esz1LLgP06flD5bGxQqY9E4W/ERgSRpWu6DXtZRSdgPrgdgRGWIFqQmUuWeC
cVKjaP3tdug++3ar1Sjritp9KhtCKfYwYUFzJEdMuxR8nbKgD6XCAv30BO/ZhHH+TMBm6OUlkTfu
OswuM21Fkw+WZIO1g20/yb4ZbV6mGxy3lUyD88gLGZHwUEd2snr0ZF5f8RYd7QmyHWdtBsYT0Acg
kV8V+v/cysR21XLnJK9Ct1VOXXddwHeogaMXABE6FB0QjWqKhfhkZUiynzrToGYlwqFGb6BgPGRM
EQX5RjWK+PC9lHgUG9lyv3eOvvKvEW8RbUX7UjYt1XJt5RBvIqYE6gWysqBT/DSiHWYE9pIgNXMf
K5AMh3ArDXbRhILk+PNMaW3c3OA776VVpb10BsWfjsmiha9JbSyPbs7x9m4AOYEK5vKjZoCono13
kMzDOG2of0l55QKudjQ5r8q5bmQB8Q7LSnls9z9EMTyIr7o9EKO9SN2t8SpgyU3w7t7dfhFOrHwx
i1SQPGM7NUf7/w8jaQTEMeWOZu5R8FIScebT63X0XxI++HsUvE48dewm/z+v8ZTFJObMIJaBHB+G
hUMqISGh5fkveSyeGGpUsVIl/IsRmQ8FFVtQJ1GC80V/Jk7Lmax3jf0UNsirWFt3NGVIMvLM5xyO
Exv1slbxLkav/guhdwYT8zOSFmfPCigr5t5zbyVF6vZvlWYNiM6USEtYETuOmRJDa3ZZvWwZnFjX
OH+XhRD6eL+MX8GMAiDSIVZ34G0vWQPrI63rx7cHDOYLsbfgjaID1NzxO798loNZKH1pj0y25PDA
F3+1e7zwnDaecIYgV1dQLFb1NZfNZcT3rorZWhug5oRFfST98eyck5Wy7yYwAGVwSPmieJ6MNkxf
tIKii5bqk7pTOzfrBKtHqDcFDFEpz3lM9xbehO9dBSsQ5HXqIcKwQOUv/CcGkEjassJCUjtJholJ
eSXOoq6ci62wTCXwWAITyqE2SMOZs6UkEBXL2wQegg7bOkKzw5ABlsPVnCCZZXpD502390hELgQz
h1m1jH1x5x+rPC2Er+y4IYFHO+9s4+9EgiHWLanaOT93G9sKCxjMOrsOE4kM+4Te+mQuy5drzIbr
A/7H3Y0Q9YIKzhntIugqG68RD7OLYoGzBXFrmQ6JSMs251iAeM6Tq1OxUWn5dfS3KrYIfY7KYnQc
lcc1QIeuqHcjxgqRV+V/hajhCwOXx1UZ2uEK98YsNVg/TfCG75aQJqHZS9FQIrzn6Kq7Kw2Y9X59
zfyh4ktK6gHZUL/g7ekxVxQlKDoYFN/SinvPCMWS9B3SbgxXPMMHfl5A6t2U4Ex7MIs99DosP4wl
hKNgwI8FO3oIHR30wcsxpYfclbQSoWGp2GyHG8hmbKkvyj2b+L3PPbyQqgTxV4HSgiWJvbv5Cxhc
ackaTgcIhyB/BpdOmmQ5aUqxRMOuzZ3yW3+MvwBlG4QPzVvph0H1kVhzc5XG2DEPbR72upDZDIzW
Ip0nvaqI5gZyNTghBVF10cbr1fol8J1FA1Fd7vdZR6KnuH/FUkUxfcm4D0wuq4qnoEnFheUf/o6D
f/9iuGaJuO/nAHhPE6o1ivcoIj6XXih8VmPduZDTOlOdZkDfa0z9Qo0CYxUuPmdqPpgNfktgzCQr
hN1GqMsI4I2aJ3AUeJUdwv8zKUL6WudnHMYhJ/RoTBc+H9wz1ZsjWsXypoZ/TXVCB19s4RlE6Yjc
aEs5VsxBNlM8NsaRMtBeXb9Il3LXBE/xgSZImyPw6xos691PbEz6pP0WGP6IwzkiG2NwVwt/FXPm
d1NBBFInQm9N6ThkVy1FJRZTCK7G1X44PHo9EWkNvpZNsnzlI0WQa8HjZ4d3LzgHRAI/SsXYgDas
LhYhOyQNKMXp9SmUOdSw3aP4zXY7Tx0vH/K6xd1GJfiZiI09JiZQ7fwX/K8vPf/+53D8wYata+pJ
zGZFybuALOe1lY+Y2HiF5UO+SqlJpIzCem5OPHkX30rXg+sse7aQaYb9rFusiZnY6kupqtVMPPk2
KJDudPDH+inHkljExVR6b8u52xGaQeNgbYCa61gBKo2s0lgj72gyXVesfbMCZ3V6/2meGbAGvEGd
OcIivaPc+Z/67nEpu9p3SX+xL8MhoRb9Aj7cRMftgi34/7JEYzyIjEqc258d6zulS3EY5LNlVxTT
mfeSmPCh7nyQQlVly5pj/U/+oYOBhTD3iJz7efw6/5YMqnyyAC4jj7x4uepj90jIhUfwhvlkWzKx
V3UG3NX/0aWjSD/pSyDDfyYgO/zESzciSj0ww3LSX6P4oIyNN89RAlSRwHP6B+3s6iZOUwW3I5Tv
1joFzEJmcHfpa9TQ2fYekoIszWKw0tNFTTqZqNmgjaNsiVx4N//wlMG9/Jp5TQqgQW8H+WX49tIh
XaswdNOoqkqUjQUfE7Z/eIinp5XMrqtopwLRfJR5+eJnHx5reZTBsBWItJgVoYkb8lbFzkVpBrud
mhs2F3T5OJiM2PqHsc2JanOZ4V7a/Vjyw9Rc2CMyy+lZaFsFy5mT/oWyzEaempe2wrsEgs6dK/y5
pj0xvF5aQiVpp30yZ3ryYmvBgr7aeIGUR0mwt1Drw1COTJvkHr5qRwEqndi46vl7Usyh5+qPhtFl
YiBmQZUR0vTte4ls/5/PxLq1gapFTxLXHric0HAFOkwFHkDK3RhEnqlJCVBavxVkVvGnZjbeSMHc
4ZZQmL4yivOA+ttGhJIkpn4Ror0iKl7xakOJ06HkgruUvmkp/XwIMw97tope+PFrLB7HfHsyrYLb
OFbtnoUqGbecRNWyLueC40mgbcX80NCxYbsfaXxXh1UOWyB7Qxs4y6qPmiCIYxB6B8Pgg1V3jH8I
xNu9fIukUuG4ypY7GirciJK21WcCsWxb4f4P9/n6iBKsangmtQLTGWCqKnb/il8o+uqzp3J3OmIH
o1E9tF0VGSOD9yWAKGXXTxZK+p3BPRKeChAQJS60KMb7DWVF9alxQE6kgiaPnFb0HoPQEvdt7vLH
mMPcoiAUdSL5iyZc66Fo0gdj9NqfFEg5MHW0zz37oHPYc8niKRTXu8knfHs7uj/QqjJo9gd5cvNI
TLLyaiLkmcvDpuUyMAwmvqTS0fh6muGPXCAv/B8tx4MrJeHKpQWN4yOHGnlUlD4M0XT9GTLPa5kI
4gaM+VQJKGHs+49PC5BgnWN66J0/UpsivyPm/cwy4IJfIJqC1++kUHuPSGCFANiNB8f2URe94CQt
Ey+TZDuTSy4Ndx7VRKBL1O7iixUqS/jh4J/6rdcRNgReRyQ463puC1HpMH9d0zHBrjqGPS8Q4/kA
5PRBCJWrE6ma37TFiUlmBaDKqrYJSmEd64mWWFAWs8SfD4hZ28i1JH+wquE8SfMgJ875r2MHM7SH
FrVCCOyLl/PvGtG9A4RGZMXV1SNxyjsbTyhn2HGtwnm54gWBRNZm+nY8Hh8JKJnQE4MpMYcZp2/r
zn9KBE/3zuNv5JJP485i38RKv6E1a8T9/I7m8vP97dU7S++msEdVpSQGjWL1OVgmGITYRY6vrT9T
0g6FWCG3ZYWFNWaTTZpcmyq0nZc1vPACN8NA+EYRDq87kMSBBf2v8JFhbnGNFIuYiG9zDGLBizpA
4HDYHWBCXVyEQ7g6cG+nM/tA2QyCiz6asS2TyZRFo7WrVHKk30MgEUpKFf5safz3bEHUyJcCQjN8
AFOYnkao6jB2dmjaWYxlHeMO0BXq3r9Qq8CTPRM7/iwSOWzKE15rYSj7oRcurJu6pvUKpcJNVQ+L
fMWOaxiPGMQ1DXIgiaETSCvglX8xu5ByA528mdRIxdaYcCYhh4v5LMDD11/NPWaTy/onZkZqeBUR
3len88VBjguNpr0apAd57iLsmQjrolTzWWkqWi+rGyST7DEbXC4RzIbf4tyybk4zfo8qxanuIvIm
QmQKW3VQ8xRRDWmcoJ75tKiILrjlu7g8beYp6FNCppuQBhFvvEcsliap3WarePLl5YB6vcGVUwYt
2ZlhtCC+SINX3dx3rQlKyRDIHkxM13v/ADk+50LJLeMdsmmqLy1fXHR9JrFE3l/kKqEuh8u8ODzL
ZBdbQhjukLXPgAdy3rE1VDl2TU7OQQieOie6uFbmglk1dIRxp01/ODb9cd4vQPd5ag3EsykxI6uO
jpjuilTy9b94j8VHz38a2NFta09x8wCr4NGJeHuapADwG4uTQHQ5K8Vd/Q0iciuFlO6VO+qAUrH3
SaaiAINOnohmYu/DSNVT4RT9Nl3yHrFMCS34+DC9HeCqD0GBqjgsxWjUwcgEU0M0HkRTJ9ByR3Kl
CWFCMnZzFi1B3eZoq0YNJp/jhzAUw+TTWrKGhif7HUCwuS+Syss//Y0flHzeBgVXliPr56l5oHEQ
Icyl5L2ofNwOq1DaJAb/UnH9t9Z3/hl98/YN3qjP741oxskI7AgND6lRdLYO9g5Yt3U/B9hZOpa1
7IOrBBvb06ZfvhPEd4Wbtv2Mzhx598xeX93WoNRereG8E7/WjF6F5JlH8f9Xq5U/sLvUWUOy1/5n
A+HkBJ/rDD/LkIs5MUx0bfvH14MoLeiBLwRkn8QWL6I/pZIbEV61derW/epfbDx2lmn2JqbhDwNZ
7UxezKPrey/shZkb1EdwJYIxdUkpfpKsDw4vMPUlS8IbUgO7wzaiAukRnK8QgoebZjIIWMI3DiNW
i7r5JowKIcEPG6YhOTwZc2Lf0RDBkDErc5zwlIUFg3kWCjXmb9TmBED0bchaAS/kFaTicAhOjYJR
TZofc0evzHwQWBmp6PwOGR15r/4rZeHYOBe/4kryGwpbztI8eMhjaRMjiKBIczKGiwkuXUWb7LSP
WskhJcTSurjpnxNH2dODCKt8NtCD8ybJr3+DNFMh9ls4d1XSByofM/+f0+yRgxp8VdWg/SnuV9Xb
Ik0KYi/IowONGLocsZPOZcILCR40ujQnabZo2CMtfJozbwcEZsisltYRMRez9M2eciwPnJdHLzoC
jA6Bhs2GMsRdEOqqnARzg1CeQxp6WMAMca7NW7K29tCvwYvTtl80zKyKkYquaxmuNv3wj6/d7DaN
cXYcpg8MyKeDImoQjVJ35vdH0HCbrc7EF8Zkoy0EMQTPi3yISs80ZuTWQUXFyfPAXvAsj02/HQir
agLELQLBthHlXMRMiEUIxhCjZy34PDtcpIbLkUoDfiSR+or/zWHq71Zz3hc0VUS5ov04Vn9ky68O
TBtu9f3U6s2ZR4VSYpO6c1m2fuGc+5mJfd9YjQhKzk+v3A29acWVyTk5qBg1MhCh1iNsnT3QMZTk
YdJypeaEmmZLNumN0kKn5WnLRbT9+Cdretdh5aKoC5mP7g6wk6S3FJCFmPZDMfFt9b0jcQ3VbAGu
FYZKM4AJ58+efsY2VBZRBWBh+aQMAnUCBQa9gbI9rErpWEpRPAR5KWFCnAD7er1OKKGi7xtqC8aa
zuZ1mQMFZhVBphnz5gyOcLt3kpnAUP0TJgs0V+wqekcELv+jyV27GXOUmgfho/kVsyG544SWuuBA
LZ261OGYKLzZv4/6xcFZQuh0LKC88bUQXt440BsJ0x0RKpI0Fk0zAD2WoRgTGcQneT+uqLcl+kIL
TM9SyGijDsgxfsjcyypM+VRjNNEXznXMaRvm0O2Ko4eaot9JrYjZ1FAU7iIk1a8G2gnBKLnUwr8B
PObTcvr1jhnoC2Na6bAXXLLHgLx0sVkf8CEa0EXtSq8cvPu5gQWcxe0S7rLAquiP/fltxUuJ2SK1
abg3bfd7GoDAIl/qJXXpOjgvagYWFI0oPIUTxb7m1dGEFiuC3NXb42CcS0CZ/b4EP98HlNT7Vogg
vBko2S/UmGwp6Kb/ngkAFdvaqbC/qu3xaRnhi3P4b0v6xR5FoKaJhJmKN9WcPBQg6dstxmZgYPWc
thiXxq869wVEi4ncqT0HT2NDE5NXI76jfnplYi4rFxWhNgtrzuvIVknpiAvafgtPgYrrUh6hb45T
IIMod7JAOgnrHWN2MiW+LPaS1CJOL4sY3gZykkzxi/3fbEBEwEs7GWgWG2w7RVhwcv7KcE0C/7QQ
2x80W5Q14gfiIQl/SrMjb3xCXr3tW6FRKMJ3AETlnshhbmdYUtYT+s+tZ1Di0Fa5tgKaDlu1VZmU
vBumJHe9eVwka+VhIUFlHJPPgXJ8D+fsuZJZNIplZbI12Crxs6v7mq7Fmci0ZFUJ9RIWx5v7tD2E
Mb/KshujWcPc8Yrd31CFPia0RxHGOpXws02ypqHBydEaa3voFHd8PqUUhCnZziPOxqTmx76M7+Qz
Ot7maCaFI4AVu8lKjUcQQyaft6ulgtIP2eBV70qsPr4/J/ZoofsuTjeMOEZgpvbfKOrHf8lxpbfg
x9XLeMlvLl39vAq16kuBwSJ1kkbU7VHj/Pj6KYOkbHsbaev4RGHD5tnsIhIDiFx+fSHC/eRi9hQj
7uP2hEtdekHn9CuN7oHIerzzZM8zEcHra8DarPmbZHP3D6GvqxyePJpD8j6Y4zHM2hdaYKgjqzZV
ZGItBbandCEtlSFQcfxjpLUKlL7i2HZRyjuKoykfXypyqUlytR5IXm+WTgb1vrG/FBhjd/ceTRaw
SMho2rDMPWsLxmgh4SNJebjtwgp27qRSaejh3Nc8AUAQxb5ko+qbfqhNcLSsFMDPIu5FShF5Wk1U
KmfrvrVPAGKF9+bUFQE+GllkVJqO+vxRjDfEpJTQLGnwSnzlCC/qQuVJLS/BtkT42cCfbpjC5H9m
oXdIZKzJ9ab5VtHL4IATE7mSMYkZOT04JPNd3sW/zAAwJpFy+8To8PEhVyP/K4Zh+fW15QgR3M0m
0AV0hu3typ8v/3l/dash0q2dXZmle6H3vPWTDsr2Z+B4nqFzKwLLOo62YwR75D1JEQg1GAqQcSw4
mUHlpKzxCy61f0rTX/cFDvXk8GxLVQsd8aYb6KFaifzHvba0GnjhxmjM5SZftQOu40uGLi45224w
TdSSX9jqzL7Ic84OqGex5w2/eO9m/rfjWZ5QUlYMP5y6z1da2rrGXZea+dPEj4aa6w9jmGynKVBA
6JnJQ0IeaR2Or4LkwUDZyZsKTmsDTU6tcD1VGl0FE2u8ekNMWk5KB2wzxQ5JdjXIptoNyzhnx2gs
70xuhpzIjEDyZoz1CoJ9RvKjvT8M1dRqBsp02ngGHlaxf+NNS05xEbLBL3osADQ2QLTwbnmMi3F9
92/kB0fcJgb9oXZlFwODVRC4YCSg287fmq4tUl01g9L/seJdR7qpb4iVUHMfyTK/99/uCOKtHORe
DnLRlG/327o5rou/Im3HTmHybdgVbcklY8PoRLSDEmP2Vrz3mfEP0WCuDf3sBdodpI/MZLDW3HM9
HXja1B70e7HUSR4N8FFXDY9QjvA8f6tiGFjT2078UEe/ABn4+xf/ychexjEUsNQLsw3iH2nfQK7w
Wu0IzpdvwgTH16pn0XYvx7NR5rl948wBqnLJNZlFzXxibZl9pv5rY/qG6zWuO1zABOJ1Cr8cEyYx
4IvekYr4YN9TW45Vs8s5+JpfuY3U3eJ9QDIwYP/h01oAtWf5Jcm51ami7oDbcr6illNRKbSlN14q
MIx3oKhPz5Y1REAu1e8s8YK/aFJWtKkpcCEfWzd7Il3Hf2pq6sFwjsmOc/Z8VZZGxyAoCiAlBpeW
cneobPZD3DozrUsmcKkAFuQjhnJPVu+jTaEIbasM1i2ehuaNfGVkL+OD9zrs4RikUvmuEC5F5Elp
rx/FXVnKPEwk/IDSdLmYXaIuLcLywW7U3pCFpSK42A2TtKjoP0rvozLcYAdxI8noNINJCu4fIe0U
6sMwyJPRf+IgO8eXUx7CYlFVFiOw0nOqNEKl2D9DrSZv8Ou/bgUDIiIV0tp+GtHqQqvmV6X9TUEA
82DEHWXuG8jHH/7goTIczlfjxh6OGu+R1H66i/aU0lWMuR6O9vAjTsey7tNgIUkuNo5ZTPKAixTK
H0WryKQ8FC+QQu9puxvJzZpddqaYQ1vyXqEA08QKIK4ypKllEl12IdS3t+jQzJY/XT31Fqnv3lr+
cddtydEvcox33kNWPRs0McCe1/j0ieP5IQgOKOfq3KWDdvQqAJsLUUNFGfaAteIuSJb7kZOOZqNF
rL/5dRo63ZGQ0Yks/c7Exnvuhsg3O0GsELHmYgbrFpIHLMEiXnh9FKIW7/FtceKgJrY+R72tabU6
ZHrUB/ki3VucpdFdZzkCWTXcGlPx+DReOhLSbmSX6pEq7r0e1d9uW1NbZC6MiNxg9WbiOJrQU74Y
RwJnNOM+LL2SroOWCg/ThUO+uOT2FPXyPlNfcSyX98rpC1JAsJEJoDl6ZL3Dp0I3e6UTDENlKEnH
8KV89AxserlmE0ejbx28BA41lV2vk0gE0qFFJciil/fv6LQaMiLTkdeB2oqrjZko91hlQDYZmMsB
Ti23RYeDB6TYmMiV/7U75OHcCX0lMFPX1qC+MxQQVpIXiuSuXt0W120c1+HJYZkiNMPXPCU9ygsc
EgxEDZaeVKuuzP0VL6LgTmol6ueZIHjEHC93T9R4lbUL5lklfwVcWgUQL7JqacH8Y0B/YPWOE97v
iq/N8KcunrMtr8J2E6SKRRs4C6289kYB4YgJ8HJ5UiVAf4I4fsXRA10N2xIs6kpW4RJI+Tx+6B6I
YlmrwLS9B57lBRXZT61hTOIZTxz5gvKDy3aFZFSI4GEsWzHKj0d02bBvBEur+Ao8e+dvYgWoDxc+
117kLst1BCmXMg7xHLeMof2iYl2iu6e+JZlgCNsG5uqvcLGEs4owVVJOuOTYq9jerSqANxTe/m7T
K+g25q2jSvEnabehnu3KUbuympO4t4dHrlG62bKIZrA2PO7vWbhkb/LiZ8TrXNZWN4hrdq9q7VCb
0QpY+sfU8skIvUFg0kdPvQcVxoKlyt61zjWndNw11hfseyaWSgubgTQD7h/lq3zw8q1XQY+qRzpI
ni/8KodOcR11xae2AL82su/kJvcJLd6ouewcwPVGT8b676z0IgTEIuDsgO+kPxqOIQy0wcQX5Zys
sPw0r2DOW3rF8zwqrYSzhXF/IvD7LqJcmiwsxEmAuJfQgDHLohc87euL3nyz/uYoL+4DYlNdn1Ki
7/WgF2zPfxNESSKypsPnMzQ6r91Nttn0Vywk9eiU0yXxf3KAfAOFoVSBf0zkV/uH0AOmnkSSJe6N
c1Rc3uPjcbsazWThTs6CapwRCmZoSf/6obBndt+hM2P2Om7V6a6hrT6QCsccy0yvHpkDaR3paQtK
mnqFLxXP3JxVoJnKRD+mQDTx81h2kS9U0TBfMxMqVJ5yjgasnNhdlce3S2oWbJc5m9LPDmFbeGl1
4J1SUvqgbWQElsVjIZPkP/PfwJGMRdSfmiYkk6Icw1Hf+nALiy0RNgBRaoEe4NpBtKSBj8QlBFaO
w0d7t4teY2mcUZWnv801U+inQX2FQJ0eCkSCRwq9x8kZvVOdnRdQe/6xBiEKv7LcyL/PFbKq1kTm
2WLZ61GuftJcqscT97P2zaY+zQsoKsLjra8WSomOKxKp8//UhI7UtIPHc1vKeOjQb3PepLilv1Kx
gfKzxwDbtzSMEZw/PJ3tC03qADqew1I8Ro57RU8+lnH2drGWW9NYL0wl4ZOoI2lFDrqLCUbXwPaf
G/P8MTm69ZA5bPy6d2iqiHsawABESv5xjHXDSokG5mx6bOYdYlKfCkvWvqucUmEVVV4TJYICqr0R
SQ3+N8ZfBZi0V+cMKfW0gN4A4QRKzXcODpqKYSiwr4+QtdCFqCwSzve/m+XsRghM0qhJyI2l2rtZ
2baiBdUmzOYK8/fB+gvN0+HwkmWp6h+wqslGhIa6bpHgqKeMM0IizmR4eUvhx73kIXBlqPvYPvk5
6Zmq/mkiHqaYpez+Vfneak3a8rJhIStaZ1jKc8teZOaleKUDidoSmGJnE2CTfdDa+y8wZlivJgpN
+m7aGL5yxYUL9Z1AQeSyViTZZrWZ2sC8dw/xd9lllN1R7QCtyjjode/EV9LZ5lvjDke9EEZ0kzhU
FtlFQDvNGLT2rPg+SYKp3si88iRtfrKUplve4TPgZ5nQnDd2RYB+e8eFOtmlEWKwAAUkgoeNjUJn
0JM8Aw9zSIdAz4T4Bz0wtEDVTO2ghou1S2D3czyiuZ7ntD5mg41YD80MUOxcfv0xqIMBYHhMCB77
0LBSM96RTVVTCIxpHCDS5XDMcSrmDuF7RbKQDu7fhr3q1k2PkA72/gaLx1NQ3XLaYFOzewRoSJk+
MOBzwuVzg/wr8bS8mVRQvOUPfSccNmjDzoaNyq0QAptxGDpPqqbntUvynj5FiVvp1hQLm+FcFqgy
JWb1afp90jid4Zxgt/zX+TNtBwETk3MHd/hIhtRjc6DtGTmYfcUB/CeU6oz5HAP36PeqAYOgHwkg
vqtEnq2Ur4G9CK+Or+J9rwY3wNOM2VM5TbQ2AY3PaulWPIbgSRs/ZIQSAJfUn2onit8R5sxk09EK
KxTg13OlDpkJnsZA5xK+a1feVhYb99438QWoKFhgQ7b9NZQ2M6I+wifRaltVJj0cO9eiV1yCId9f
0qzzn93oXuFYPurhll+MZQapIMgoQ1mHuYJAiN8UPgicZDjaVsrv1sVO+PChxghCLo/53Lq18gUy
2f8XPzIEcndlrEhBCRb584+hcXtBHLCioxEeD60C2c3QPp6veo9lNFDxrG+wVRIUA32Re5RtxA0P
J6DHm9kGEARdCCwZl9y6V54Eo+oZztqd0D5ckZYP2ZGBJiejY8cvGU+Luni5mi/CWsG5KjSuCKRJ
w5CloNVPB7tX+lcIQl0v6qvjVEc9+aiH1uZBr8lNjh+0wJzbcn8RUXKkg+rbt/uj84n3QS1dvfdk
V40CvrU+Lx7j9b+yP0ffDUeS6PpcEa9ekug2YzgqPiE89rqeMqaAVZsMsWZzuaQpVETiLKivJ54x
ihICD6UZfYBX3hGQtcS8dYHN8sSKUK3+9rHVLYXHHMwTAUbXuTjAoiQVV4Z6j5T4ARQWInY6fnV1
NRIF+bfZu8xM7PUbHTcf90yeEcWGeptEBJt+I3F7Ypia5vUMgj1qePeiPfARK7SbxbxV7VMpqM4P
EGgF7Wxc6FFw0toJzlwYHMTsedpz+gfo2CXrBXM8B4GlY9DaDOr3VZU8HE/mt7NPLAVKeWwxcVp3
46h4Gc3avoOoM7NZKwAD7MggQvu1jL5Xh/gAqXtWZx/GKmfbg9zlUFvT9jw8L914JUQGUIr+bfB+
RKSZN3H8/kmv5z7azrw1eODnVUialbEqeeVj0Tws1SNS0IIt1Bl/ODIXGkMQ7GLWh6MD6rxbFpYq
cpQ3TJ3dLtdHd4klep2730yurSt5pl94gYYlZbuPW2FT+DTRscS4nn9RXKX/IFD0dzBZcaPWDKny
j+YDL1sIlhu1dXhgoiZ1xVpmToaHYjgYHGi2e0lmNZvjgSenoGj2eM6VhYpH2H3xCqrodz58Ugz/
ZVUR3sgTYx80nACpbT9IQ81bMM8hjSP/7/lGuEpkpwjmrxCGuk8vCAkfcxo1Ol1bLZEdYYBbKTUh
Wg9kqlkyPt6VOR4gBd53Ggd6tKK87oyjj9cmX9x68S90Uku2IennDJqhUhE+gkPF48Clo/Ch6ytg
zu49mEptD8im2zeMBxAYUCQvvH//BNE2wvgilAjewr9AzB9JIXMMOylfBXt1//3CcoE4LlkNxWMe
kfZHjUn33t+kzVapw/UflhV9ATYpxNnyj724SLO9J/qh6tQhP+Xx6zPZJAB+qyZwRo7rVl9LU1gO
xwUXfGN0keMhoowwCOT/7Ya3F7e2KJnNWTB/K7RveAY3ijQaolsW3C2Ts9pG/WHMCEnGhw+zPLY7
jqLXGzES0THC4w5ScNvgPSK+hedgymvJxYHfIN+Qf1To+XxSm8m6F7KtJhlvxJoxCQzlPUjc2Xw+
hbe/2azyRzmtgsmAoFsTuD7iHjhuXI8RjJhDu3O+pstEZq0jXfybP7ID2ZMaBDvRWl9zZ/MI5YEd
1FL+09Ou0hWsdDHxymzYxIt8QXAsBIWLkcxvCJuuj6I8/uS9I3LgR2GLg+i5gmgBdBamxrGjKbsx
yJyCAtV/T2MXplG7mEWrtefPOQ513a8cH1si8wpvY1W2tZukwqG9zYIZCf64yRaT3cIaCTOjcbKU
ekrabLnidZls2yzqQmjLisd4E5ygJqGKvjfx8UmNt8YAJnTSvRWBt8KxL9h1ttsKuoB87Arl1Crr
2JC6lh1wY482pl33vzFAKgP87HFEG4zCLSA314i3ynHIrxWSrzsT3d17jj0fqFE0YFx9Ps8/AkFR
9WgLzKLhaDAeWE8rqvl7lxCYxTw9K/1jWv2BHRSYk//te9Zn652jwDqX8lbF0+Yh64UUSX5V3qac
3+3CHu/4M62kYNRs68GNRBSkc07r4yicOApIajB3AxiyBoXtaX18RylokL1tbIDtocfuKwAIWBqM
BtcN18Fgy+BIAzFjcl5QvRIDXkLto53iR16tkG1xrDOpE2KtXPuRiTkHsJtd/wCPPPqLufYJhJ9R
ELIVP8toj31vmxpr0PMKNE/sxySvF3TIX1gt4gmkEEUGQU5eSmxeN6uDsQnksPLE9bDiVonU6Bfd
Mxq96G08NocdfrIjLihw+1xPEWq7qCsmjBYWBODiTCbMpN5HwRyl9PXOFJ+oF5Tr7k9MEAAZGXyp
7yzBw9wNkLH3gwpeLzwi3w/9Z3MhFpSANyBLLo3dHl8OuWcchi65Uamn7UOl39giHwxReaaq3kHs
GyTm1gX+uAr1gad7+pnD7bK7HzpFFsVctW9y+wiPjtXFKAR3hRLCf+8CMBxz520CY65m+2NfWmWZ
RimMSACGqL+UBvRnNfFe9pk9QvKCG/TxDSEq4ye9BEFP6k0u0J2slfq1iaAOpWJg5AfKVAwS+ydb
qBKQd1Axha+XGuqXNzE3zOIe6cvtIDSORZHsw4xd/3uMFn+NTVGwUWRgq/CuigdG0CXQGxI5VVul
LcKWkGoHOGDOE917mu3rgH0cNb3nLUb6ZmyL2CZBq7WYOdmtQRklAx8RMYlqzXJLb1NcR3oC4kth
+u8uNEr9QemvHn/fqlv+T3f7SrWqrJ5eflRcPwCSIb+DZbN03V8WlINg2k3oX7zqoAySodQgXzYh
ywr0dSWo9lfLN7qfKqlIjJji9B0jf60e2JhcjWwIGhbULdDaI3xNQlpHqsvKgQmK62lHoNPDMopd
O8CUHuoDZ+g91DX4c3L75/bh0iGOV14EPcXGUm4RNufmZ6ajfrmDzVoEO4SHppx8L9lIn5/UhDTj
6XaTk3yHsneREgHTl7Zmod/4Zfn0E49bRJQ4qzdr1Tjb/Sq3cZNiaLYelX6bCNQuAjxDb+Q73dPa
Lv5PPxw9HPl9HJO/T0M5fnhy/jS7YPTXKdmdCgxgd/WiFzVKqYo8Cv4jvYkWltE7E2j4pMUUJJ1K
aZtc/C0yLnIaiRmWgQfGUcdY7DWb52YkfZJiLIPEjwETTu9UTeHg61XpP5ycuzcMAaSr8yaiN3BI
p6IC3oXNV8DY9tH58CZLQW5mtF3mKI3pgf/itGSj78gygF7nrfjaI9Ym0VGGoMpFdKkSHVpXTOZ/
6aF5uiOlQZeF+CR/6kWceGjxZutL5rNO2ErVi8yhj0vJEf4XACjxUIGQNZcgiiRsP4YenYu7WZZ1
KO22CnlzGFYvrfaUXHlq7470BhAXRGexqSpHmGBHA117CcSHCxIY1FWjDuhzjpm0eS5UvU9D8G3E
NfJ6BzzG4tjz4sxBkvzx6p1uWwVTFHAjDFYi0K23+RsdK9Tquy/cQu6VR91nOMJjKgx8oYutvVtL
cYXDaEkJ8UcypG+48nW6KYDnNwyNYZsM2xWlXnDwCAAwhpY+SY7A4UoIeK+p/9Yuh73Oi8Y9EtuF
B6zVuRbR162/do1KOu7AMugpBWvJsyZnTiaTsB1c/cqWO81O5X2LyEovF9IkTqhvHmWnPVKPKxg8
1h94kd+gTGMD38odCecV+mA0cRaTsuHGjEDgiQV2DK3EYzga8QbL6l/o4jRv3ydtamkCi6OffkTN
VVLPhdwr7xg4wbAa5N/MgmYK+6YzNMR2hlafAjTCk0jmCpxeVJyhybMt4B8V52v1degVaACjE3JL
fH4iD8tlc2wX6UiNQIW05Rw2UJZ6J5gr0/btCieP+cMAy0cW23u4v5KrYn2Dtt/9EuVJFSuhumKq
buRnNI9hfohMjn9K/oGYnPUzxxLXUzHqcCXhxcHXN3/Fd3IMB0nBynuwFRbJUU2UHMQpFCV9uT3N
3b+9i4C+5IyXadl8T0KuO6/UmN7uz2Spxks8h86qxdCzb35ekDkN1uo+K4riB45FOvpKGHkPgKAm
17+ZLV5k1PAfT6eOZ/gqB/g+2qCQdT8uPLnXC73uxMugUYX+o8IQNeTibHyS0zR3Co8hsJkuG9wa
bNye/R+7gRC64Z9DW9Ww/1tVGQkpQkSB5Qnu/hIfNy9rJ7lz5jivnYzm4zG6FudvX4x+KXvSJ/p7
eNqUmzlKOcO8MV6fcdtOfC22T+VL594AQ5GPrf0j5lr6MWCXgiKwW1GoA0PgabzPl0iuZBlQ2EwX
jLgB/pA1w3WOwywLDrTrHOi1Np++NhJ9uOeOhOeE2GMyqJIozFyGc29HCl8cyd+Cm0Jallu/KOFx
wPyxIFsewdu0iDlWSV0pg65hgmQxn8VbSUA6k6heVSmoDKsjrAcx7fMu/roeOPDf+dNYtHmmhuh8
OzsNuqoj0nszvydzaA2q5OxqpGXc0UO4AYl7nzp/Nbd8g7Y7ZMr9wOVAPiXA47OMoeW2SERov8NK
fa4zvlG7APwsTiecc2WEuZnTv3hKbraWMaV1xbC5O85FdVxuxCvF5AKEjno3aenXeQzeP/I05dAB
9YVynh94pMV/KCY+iMYPxqFXfzRY2zx2vRVeDPG46IYRaxpPtdAVykgHk8xfFea78k4qgkj/1lnA
8IO7El0AjNoAbJHtxGsW9tGTJP2LKPdKfhrQNFUMBdZfR6+9qTRdjrRVFJC+9g4ETenw+4RMfDQL
AezcvSq1cOXHw1+VKyg7gvRDLn4oCEe501WhmWVTnZeHHcBR/w7k3iw2tmR62cHrmhCcQGXygo0W
F0hMfncajVkBI6lU/i9ihCrpwqmbLf+en+4OPIJhiBivDAdYG3PRA6KOHps3oWHddodblQzUqAG2
QyZxBADrsZp23/CI1tw57hnC60muY0sVAeS6/+ojHm0JCRN+mBSXkJRKmeEnEKdSbPsAf+ZCOcsV
xab1AkcmDmdiOsST2MlUTyGj6FOaY+wN49Pvou+ddoVZn9bT2p9ExWAHAh6XUdvOC7mqXle/9gf3
86/549QU2rtWl18YIZ4QYFGo93qUrvp/zFBuJXrxMxsiihvuH3cjZI6X9642aTV++KWQpSbrfiTm
6gMpB5m9a5RzZKngsVNrQUmNSltIPgre7XPLLv+80UkS+Iywf2HwhcROkXB3L2s3jCGyXvgd6iH0
oOKCF5TeAQXkXHwY4gSMCabXSpehNvU3i4iKN+Rdb3lZvxNbK81J3VuobqHo+LilN1lLlTC0QjD6
y2oL+dmrYlbtTOV01yxWpmZP9e3TkucmDLI8VNWTghVXemjJ/UR7LmtpC3Ey2oqpgjvCIR0pKtB0
H+VeF1GB0tLNgdTkULDqb7XGLqnH3XPb5IhAer1lA3Wy6Iauo4pQbzRwEgtktePqRSuIUotKeARA
HD8waGkM/VRdm91dM0gObXYpEZXjuPaxJUkieNKceAJK9PpEcWrRaul4USD4PLdhd2wNVMPs0/KY
OXtV1DtARCthtPmKCLt+ls0+GkUnEl4Z776lLDID6Mr11uAhTx7j0n9ZkKr0eplNdzx6GdAiHZss
WuPKwhRn2kkIlj/SOllPeL0ylft+cgHiL7YnP6AW18iNgJQaG0E9G91w2q7iGJYBiD+tRnc5VooY
hK7MntvheUxzCS1DtlFwG/pVNNCm2qvNj3bZM88wQiE7HSlvkFm8ZlZrAeXimzUN2scf3ycM79Ay
BfW3EPjGcDmKCvZuUQbYALd7Jktq+FFEDEZVeVGqso6latZIcXWAnlqHk2NJJrovlMFmorYhbgPB
HBQ17JuNXqWXB0Sv3VP982pm75eR2jPB1EKk/8fle/K0/F+2EuAP5g8VIRAeNtI9seLyIsW/yBV0
mHZA7mU8CJtu1zMchHFfH6jlLmvv59lUid71v+XDXYs7RISBjC31SPxv9d8mp8i5jmZtUbZRi9hz
ZPJS4eBqx0mF9bg6KO3+6akkJDm1c9FeRtZhhLbtGKberWHy0Wi+VLXahjSqQWrNzAkoz+Hm/lMo
Ld3Tw7z3T6/StwEPuVRTfY/xNFLSRGQ7tYI0/hEUCJValpfGsfGhxZm0rbw6Cg6WxV57dLPTa/hs
dyCJ2bR48McwDUTt1nYXfkAGE4Mckf/RppGQkPnLLgDReFY5xLIjXHiyuBd1fmdmvVKiANMhUJnk
s87CMXQ/ji1XiCztLUD5M+Zz9+hhdnR04xykwsbUXkEdvOMkwFDNfT8ysoVni2/6MzHQAlZQ6geh
v5w1f8qPTPo4WjaZAYOOnb3LBPUSEyG7HfgrH4wI2V1N0WmOIbM9KQAc0vXlq8qq3aFKo2/nkLil
1eyWgqzpMw+9EfPiLERmDCr3OtX3huvt+I9L6RpRXxL57wUEB/6iLx0IKEWeRz0cD/zBFlYZQMwj
1ogz2Ofx65+/CA/LoNdeiajBfkncRytkqmEOVAYp0wsz4eUYZvmJnACiA9zehVpBuXWnpoUrA/A2
505Eu/3L4oeMGbntJKaQFHJoWA/XdJLVZ9Qba63PnAkcbIqJxcZ8oGFz77U6kbh6FrIe8mtVknZ0
P+W5mTq60vYiG4VHC0ZXRTWu3DKmSthEgt3Mj25twGQXwCqbMP6AjiPefJryu/UGqrrB+X1xXKT+
PiD5jeArTnTYoWFJS95G0iLox967PXIjUhY9wLWWXT27QAw5wj3jCvH81aEXapPfJcr0xNsK6lBd
Yk29sxkhYQBx8ALRbPIxIdnWtx3H6VwFgpWuNG4AcCjEKaqA4pXDiWPGnnIJySNzg8CuoNShwLx3
IXqk1fRzqefjiNXzqGDMjWGXPIUM/C84dXfsal0xOofFdDmg6JCG9QanJraPewuaBIXGbt8PSsha
OHmqFklvO5xSMsYFXFkg6snoDXuktsnSd4guAzX4jr5zoTNX5p5Nt67q8IXO2uYhsOiYmGjO+BEB
lblnIQnhdVcLusMJoGhBI6c2qm9S9+/OG3BX7CY5jm1NJOhNMjpF0hbd3+uOO15RajfCXA8WraLN
Blx2xfjApu03asiANBACit1E0wQeIEDSKZ7DOo7lk60clsRy30bqm2DdJdJBAwktVvE3Oi3cjVzE
Tetaorp8Wj9o+vxd/DreHjry3VL086aJ3N9Pg6kUo2Bzu6Pn333bw+yYKx1/D2QWTC9oXkt/0CRw
dulJCtPgOOw7UlFK8JdU6uEXGZWOheV2vBT16Vd4gLEIRz3ge60kNrEDleZC91ILV1Vbq39MTjjS
RRVVpSB+vx6FpLcrqPHX+EgfY2Z3EgiFcJNWgqBeKL5RAjC+pxuMyNAYGnCZtSRPb7BU1YC+uHGd
2x1/Kqyd7SNoDe1XtlIdBOAj/BF1UB0t3HE8YDyrH1h1NI8jwJcxx9mx7Du7HsM+0YWKTlX6ZeB8
9gBrFsNTmzK42rhHLGLNx8aeaWLs+DtdlL9pRToSXZl23FbjtwDucEu+0QnU9mL+LHbSHEcHd0yB
JTOCDe528eIoE2cBQvVJU4DSorwHqxjI34vpGRjqdxF9zp1l4WRIBIsR/IzTn/0CmwqOmFuzlz4b
6GonTljvRv3+gQyt7ZJMtp+tde87YmFC6aZqLS4vIOfjNZFl2N//f0/MV5fjx3faxqdHfaqKB394
9KqOTFTj+JK9pObukYie4uia1BKg4EEt/8dPn1ziAxrHvB4nY3M1H5rRcXYpkITgAuKKoZNjBR6g
kjvNJhKE1eBLWs8wTdO0SJdLZ3icVi/khiR9tC9cGBaChcalT/m2GiNTwKRKI+neFse48926Ze7m
FUVv+DuaLnxPwqFsaiLji74gk0pxDhpS6BfDvcXGc4IaJ95CnNPvWrIixZmFmzLemx4nObN11mGg
Xy7dh48PADTkD1VrBBZn/Wb38gx+odoakpgwFKokO+8Ni/tE74dUfEWuoCl09sLVl9/mtFFlP1GH
IeD/2nRaOosAYd3+jllYvGzWxm0DF9CVDjfT/8aLD0Ox7x+8BQOwL00IdcTTMmVQ1mOOwY8rk+tr
i8E4ubIyfRUee+PImK65KExZPf6ZpPYGzzs7Rfb6F/bYcVsCCyY73IdYdzUCV/SYm44HDc1WrR4b
3z+WqKjqEJtJoMZoDuPqdL2I0xCAxaHcqbFiOuQKQHlxc2jKGq0T+9hnR12Go9Om9SvEgT1CpqoQ
Xk8ziwrniDmUYVCUNDx0rfobPTV9d+vKobKKt+FNX40nc8n3nLY/+z6M6v8LVU3qdGeVz/Vi813g
9BjoOOl3RXXgFuBH7aUXWrytsHM63KGdr6v0orbNg/xKIMA4WO70f/CaEtQIh5FxgrITg+NmPbyW
sOPtKfAKrxb6jLLyHMdd9l9ggIZAaNpK4DcVblWnCEuMim5dM0TNMMEqTD5IzvQbMJbA6nc3zIiY
0xyzl1GLqBCgLYkFImKMmDh7YYaNvOixm7Gh7PfCtbiFBm0t8uoqH5o5aVYF7Bewt+w5c/NMaBlH
rYAvqZY8hzlauUpWVX079+J0U5pHJhZoP6T+I2Zkqm2ehbnywUlDulD77AP8s7AlCkIMYJjddr1N
5lHDTL4pmbeKqFW2zJjQgVOhHn2i9E1B2kpsQN5H7uqcMOAOZ6X/sxmphxmsLEqHULZ4G1AuSNYD
clGbfVVyPFVwi8DKN29sx/Rm58MYN7U0+sAeakEtxk2IMX8syFI27LB0VRQjzaQ1oaalo8SGXhso
vCnYF5nEzDj8LaScdZM4RRTtRFEGSbYHzOpCHxcIAhBYCbsSgBkjqDuMJw0NjQ/JjEX/dpOWJzxV
jnYd+1BaK1f7WwhAhwhZ4mhjgazxlJmQfd5hIyLkB45WrHUKfWluviA/XRxFdJpBnTbYkD18K/kj
8jmjPYI5jmIKhKucoC0cnLK65R+BobOJSKoisCozW0NKI1fRQadqohIcpcfBUMooU7Eah9wIGU6w
JVuAGtNwYgl/vw3lwvWBA/vTKnWro6eCWUc8YnyZpEbh6QdJDxQF19gD1mwd6QVCUqgfKgrj9A8N
0NsD+S27f8FrMagIpcFRKafPNXbey8aVzABS6+A6KNQCKnacadU0V/RgXQj0jO15E4vL/irfIvA3
oCuNCx/PLoOfelf9dYT6ujxYbfrkWWjbd6JNYuPWdppLS9ENpWDpo+ppWCUppXiEdK97Hez3uVxj
cVgeEQqE0s6wDgg+Wp/TzNZqAqglp9v7EoCGe1ljCXWXYoZtLXcvMTu1uj6p1nxiUO/Bfz3QbSyO
qCYTqbzL2O1h82PRbemj0HSBvCkHTcvzn/YQCent71MHvbc5nxQnAGKHu2yvG4hM5HKesQwSE3Ml
FL4mqP0yiBoRRCgZlX28+n5+07FAVgzSlBSdmx3b/WHupX75gcaVExXMrJLYp5Sh6B1nRjyP+/gO
u7vTGlv1Zw7NbkU6hd4qPJO+AvtDrbNmADRW+9scOr/QpXRQw3sfIGLJQE95F+bto0yO2vh5AxeM
UBhA8Vw6A1Mgw6S/EzQCc2Vtu36nO1tpjgrG2TNm6+EjOix+6SFcmvvKaHqnP5T8lCMpYILlenl1
VAkEtKJHuR9uhwJ2obWx895DWzsYQbhMT/Ci6T0g/SRynFpQlSv+hoJJbn8UNnMs4C9Jwu/nMglP
lhdJwrosjt+zWCaydI4gxtZQp2G+F0QQMjQK41pSmxFsRQJEwtuIIsd3QylBv8FMkTJykpeREklf
5MDapPMDmgBqohnv/JgqviGW/c0H8ApD0UFYBfll59SIUn7Jk1eGCRLP0T7vK0aUd12qrtc+0AU5
FLsUO6PIgALNQeUhwuUCQb17JRJoFX3L3UKzXTLcCXp7DzzPSG3at4qTHwHS76sSdAmXXAfNR1OD
FIU9tiURPf+v03FsResxXjOVPEa4pIqYdBzTAZykmwlY2Rn0XUzi+XcQiMGD3mr0gT7my2Ks8SEX
I16sFqU9fHF+88FhqpJE3f0AFhYB+NGor9MxR55QDu4k/L/VCd0hd60tgtEtuwJbEPWqLBuAsGY9
U4mFOApiMOh4ypeehACKA4a4V3KDn8F8Kdao+duLfrlyrMdEmLQii/42qmGaxE/LxGJPaJEHnq0a
HlwSvLVAzDz2LC0aSukOC69FU4vu3LEo7hyYpxlCl8uSZrOrcKieJ5Bk+Vavz4FATXXT0t5Z7ifT
M8y2+3VEhMIsoUlmIgYY6FRPeknmj8+BGc48r1+F0+fnEWROt72De0a39o1xvf/3WU0UIFunzJZy
pcqGSmWT7BUsaZZlxq40KbT77+gqBu7ib9D9rOF1FNfmHEi0IvFbBLUHhVUdd8lHwam6skKv+tAQ
qd9tFTme41Fz8rqNpg2Enx+TD8fvSrb8+G1DKCJIoQKXSV8atNiXW3I+Hi5lVgrEYe9Bjd8YJPaq
uz83hy3zZ6mLcAwdUKEwXBBuQS73ukR+7eiFTcDoPgvCEjDJDtwWSMoXJmOdl8auELzvpecWB+Ho
IPtaKnE8XRnmpvH+ovL3NWbzsDFKskBz4hONTd0137At7jBCMhXI4OsO0UGIQvVHtZTwFy5H+EXH
1nD+izPcT/le5NlmtwqFIuuPuWZ8Ltalof4UWhCG58mi7jb5Qzw7OYbLfo9UFcjJc6jp5GWNQzFI
s8A8nZo4uLoJKBQ3xVWF3K01HCnRwgOyNm94OfmDT8vW0X7ubty2baGflGz+ARm4T7+zHHNzSC9p
zha2o8yrKWFcTRbtKZIvUmC3itsjA1KDIFJBVY6sM5aMtkbFJrS1R0TnPmWaENuwy+ol8Padf20S
tLlamxbXQRbOLCJ/v3Qi0LuSWyM+Gu5cwGmTYIonvuhf227d49FbBsC+BjwovO67EtpL5v1vlaLR
05muTynWwL+dleIJpghXC22TCX7ApV0O+13lUoAscUhM1msNcrI4fXJO3ZA42iIwChIOHZIYrWHN
KTKpH8FVsM7sQDM6SrdHWjT55bzsdi9qjGGtC6Gu+k7kK4Hbnw+yRrKlqkQoOPrLuhlvwVkQ8Aq3
I1JaGpVKjc9Q75s9tD54OHhd3AyvsyjNmyrZqe3VQyGE4++cRFqEemN4JXI3HERBz3FlPlHq8+Ss
uiLLTYPmtEV1qj3FhvED7s2FcUoZHF/22Ysb9XGC4wmxUcjaf4gBD5gKqik7Z06efzOlJezuQyVS
9XakSr4yf0ARCtXnmDvNJaHauM/8B1fak4ZZBYmtGjrj73G+5V7V2JZ1DbjwDbcJSIAEx71UECjV
qB6pvqFBYqDI7K4UGq45jTXiM8uyD/P2lGfM4nDcaAcOru8Sy8qDUol5GTrbrFOgYjQM2v28rMx/
MoxQrj3YBQrkMyI2amrpU496g2+Weckg9OIq0M6vpEg3cEJzJ3Fh031y1hNcY3MR0aOs7qSfVkcI
lPhr/HsmdkC4+y1Q78HUn3VY/3zZXHdGD3LmQprwzYjA2R1vQws084wrwOHrT3OAS8RFLALo6jRv
ZTsGOtItvD+MQ/Ip8DbUVyRz/9TQAmuIafUDv6BcJ4cKf+NAXZ24D33WXhXPUUEoOd4SfhuxkvCe
LFnaP8cul+IZDGP6ZdHyZwkdiebHrx81VjcL24CLG+qn4UkbdRyw6nYhPyyfzSgXPwalzp/VfBh7
w6wg0KDp0R30MJ3DbJedEsM4ReG2kdvmhuETr+yP+mY0rymXpHvQhHdTMloytLGiyvCmL1O4S+IG
eV6TkI0xtEsDhREFFjS1PtGeCy6TVrUGSLMrZtL/rvwcywxVJC/i2vrD8rGOqtYvt9c7Z2Rs/cgw
j8Hg9qp3HG4CyD7kIFbn83yJ08O+exLs5OM0dD/LWGCN6TR7EIOte9A9zykdxsEVBH0+OlunSxjE
BmsT3hikcNeGMH8lQ5+Br7GP0FQ3OZ1FYkbeLry9LgbICAFxBStdAHtEQQ6ErBElpuyD6a76eZ82
VhNcZ7mWWTSc5mgFmDc07dS7smCQfkPW2UDhY4FTfzzM0yVVajGwUCaMdfUG3nm4Xr7l7qq5Pum+
PpjlbplOv16iSnZmnn7pdlavz2SJ6S17ZgIebXgUMDD8y/mgHxmvpJPPtwkjSHhRZFjjpe4g6K4u
KZNaIVJqQx9riem2p2XFGWorG34mLHhi5P+3z7l2LgclVLqBIPJsTMs/K/GfkCHPbOjUVVqlIZsI
7zkY1NTN6RO76/LWPcGEX3zw5V8JVNnI+/mM6ZFKyQ2w/K2MEJ96fUZqFV11siCieT/MXVSMTMG3
uw/rq4Cq7S0XzKrRN1Gzc88NhnI/fRx8X5d1HPT8npgWODI40S2l/jLZpf9Y4pAzcw+fWuV7viAz
XSr5qMXIAYxvqaFwe7rK26fYqyApizfVH2dfcUhTXeWvMz8OnJ+3ohMFKPzzT4PT7UAajfIoZb6v
mOkfvSAvNMt3x8GKgz3Me2FQSOAiDFZMN8qHBggIFQ6f7bJZ5Y6MUoy/nCDSzJNRugQXztB2LTzF
Pzenzu4uXEf7zIpscHWWWtz38JwLb0eYEQEmK1S0tiVCcg5juLMFnyt0G6nvCIBczGJQcFZ+CLLm
SPpO0WOCmo0fhsqVvy/VeiNGcHqGkMCNjEMxTQLrP+DQSomGzevSUk+96vIn1mUL2tlJhqUAniAY
2HmxaPKo3FPYy0LtOXkUhrL2pt83h4k17mz/iFI2qJy0Xa+opnwNbqQGVAbQlDtd7auMknCybDQn
FPgS2Kml5w7h/9B0QQM1eNhC/K9T3zgLv+yscxNa2vNzr3oyZ2FYBa+AbgLxkOJQAA9lOLeCiVd5
uQy1oA+DEpjHXzfUuyX27M/4R6fGz4HXH8pEEXeyq2U+Ape4pcNmWo6KEKiC2QANvLrirNU1dKIm
ubD2Sp4w3CxOgVPXuKJ2oq0HB3O2Vs3d+bKVWGrYTe25JeG1/epbUuO6T8n9+llgUX8FcxphxfzD
5BnaU5/PmPxHFHDEzlI9awP8msDzLgQy2UOBWpxkebwZVDjSHRhkjFqH7csc6/MnCycDq18JU/5Y
QvSNW1jC4HN5qyPijYOGmJbgokX1I6wPTL4/dmLDWSvTqvKBngD1x3tghGbDkccOMt3kLJXI36ce
+2lXbkP5mZLSvvqQ8kRpILtW7IYfpReNMOWSZk5bdz6NpHH18ZOIVSD8hKQ7y3dxQBuiJ1Qnq/m6
Nrqyjkyh8D7PgRdPcxghJCVHMxVymkTXeL8yvsnb6XFMGhz/11sVjSdoUit7tZUfQet+1xOrJLEi
NqdCmxWFk1FiWs25Zo8R4rBtU7MHzBJ2OeeHXLwWUzbb1t0WfuMDgUJa7VOzc3PdoV+2xOIezmD4
W2OZABX2KKJ0sYUzPWR0NGnR7JserCh9Zcmz7vVaH3YSdPdeXY2p+NuwSBLMS6gwf3NNUSWmozKz
C7jgSWrp2wG0QUNImJhPsIYuR+1qzhnUkqxsYBYxrDOL4yeo/5cAG3/MjhCf+/IPbNLRsEX0q3ux
mM/fdXeS8TmUf/ftDgmqZ357qH37BaxWfANdnG7QlCrtF9tD2RyXbencl/oLH+7rVxsxt3wSP9lW
rtXr3KKj4+UEpPL4/nXhUj1ln5xC/s0Uo1iKvPa+wJgtk0FVahIHJ+i2fDafNCPEvt/QZ3LuaVqF
/72DD9/Qd2v7IPP9YxYu4ITlGZcZYPFDo2KlO8OfJkJPSyKWTryhDyY3D73SKyCOzFdfXsi6+MS/
s8VU1AD1tPaOVkoGXxHnhdFq+FPG3Fe9NFbhAX5mCz+rsyGZ/UBaJkMgKWS04kICQXD6Mpnq2XdG
jb0gg/apPKlGdbeKlrQYR3+KLccoFrzZiu/o8DuVUGxhJ0YQXp5VorB+BT4MGnDmikx68XuK6dsp
E6UE/t5BQofomHrN6q4fmq/FjV5EXyKVrbTC5+IwPyUthrrkI/BSLEDEsN1MxBwj9M0R4vC7fxle
b+dsjlbxAO5CLOiC3eX4LLmYLywjAL4QwW1IEbxU38UwvKh5oO2fDL+4+DUddMS4CuutwktJ7ft7
bwPiKs7j1WZcgm+W3CEL6ec6HbNis6hrDSnEZBe9EDnZy0F8RNTfJddZtIe6EjdZBveGjOKLiPwH
rM1TWboKlP962a/MHZXfZ6M11cJKBnraDNCKoECwbg+QdWjcmRI2NOWJLDNaWOMrkB8Wn90Qvfmf
9gfF2u+v834zLwjnHHne67Ap6fFqCQSYcorIDC8rKJagLrm+xGCA9Ghbg2sxUvoBsoKFbLK0KsOZ
Zvy96luophBbF0fEz4pL/X7KEZABx1lk3FLFu0TZlUmqRRtJBBVzwqeuPsOztVVaAHHEZrK0pLRD
npMVJKIYJsmzNKv9IJ+H18hw8Lnb4x8j+WDYF9oPoTI9FgzmB1Sv856sHOhg6+j17XJ7GhfjUr2M
hjmv50Sj/J5T7g1nl3AlJ50A3vUZJhSI1jie0rWMgBs4vQugG2b0B0nen9jZuBdvgMIqyiFm2k2x
n4c4N9Qzb55Ytk8SPvvqCK52N8JJq9Lh8EIu/zq8uw3ja/Jmv5ssR6k/bKfFpiPsot+rlrBknQGA
C6mWxm+b2dDwTudAT8XGfYtIQBLwxePsnw04iK9BZROAWMCMqwOzH8caxpyQB3FhKXzaM74gH/v6
JIgnsEkXFfmbrkKHerFlHU7dXWYD9IrVzhAF2NK5E8sj+xsHlsOGNc7bruGK8e4Txdx/lSXtNO1G
eHbm4DvNR3FLmiDtb3dIk4MEms4qWCK0wsL14LDn5mXupkwgrlVHOi4bVpWe1ufszlRgSWUeVbeg
j6Xd7pf8RHwy13KTWisttpBLksiHTQKURgJwdnSUSanV17pog8wSjV5xNSCNvF/8mOFXdEdH6soA
jz7Cro0jPeM2D1wjoARqyERjhHAS/foRwoIjME5BFVFzPgm2z/y78UXR/FtKZvrrjqS2eM+72pcP
aq5XZ5LHFcsi3OL9iWXNC3+o2k70FOZ5byA6sn4Neg3YLOcwJDEORVDiun4jbHmCKfrSF2X4DaWC
UoPpYCMhwytp5mpRCTEA1JU+Gcqv+YDlMzPNjcbRpdWccoIpSFpTM9l6DNu1jHBJwAB+QbuRQTMP
PeSpHwptv4TJw/HeluDiVNUR0M5kOj0pTyyX+2CatrhPJxZegOuCpcxTINjDbNf9hhptS059BkqI
6LW6gaL8F4Ct5tz5awMwnd1a+2vkKcgrxattNCGXyTkZXOZscgA7sFeNgUmWjASDQBBkXc3hrpRF
ouLMDXl00wDob2AUG5PqYiQ3AdP0knynY2BaTrjlXoHKHU/rpKb/N8DcMDClLBzZixCu+p2P9/l/
YjVGrmx93Fyp/gZhlMZhvDGsr1x0lAz6cWBpHwnY1b39Jdxp+aan29Xt/ueLRt4D40+piOL2Gnjv
5E9SL+yybeSIyO6rMMJ+b/h0GFe9at8FIsGfBpLHaVRJYMHJZIhwtULxiKSV+W+02rrvq3sqyAPl
EO5sz5r0akShg1D5dY3qwc+IW3lcmIA6eoDh/tLXLxon7olZy4l/XVVUZ+Ddn33iL14ucE6bUAd9
Rdn2Su6e/POTYsdubv1ngLS1vrHtooslC/Kh0vlGB6e3tAH1DOdSHzkzf4hsTQaH2WVKA4OXRhP+
ygEgzK/SpK9kQtD550+qKtKvMNxQ9T42zM3KbyEpjvgosjnaRem7kBi9ztB2DXGLem8ZRcD8UHos
WxdGXg9PFewFm3KiGylUUyXVtJWKNSF0SOgLPEQs6Wqv8O3fgZ7xFZczs8vZ4grXpuxwLr6y/C5L
nPuCZx+auGPUTL8VEIFFswhP+8AI9ZfyjIdZc9oI3xfDaZVh9HSOTg2t86lWD956WNGWMaBW/7cU
1i/wsyvGQYh8Lx3Hl5hHLsZGsQXCbiOXB4y11dY+3LO7GaqTkU2CxSZY7Gms2qSz449NYF3SrOdL
Le91WYhq/bXdScHZrLkVlW1VCz2BNuTvZNxitIt60RBNfuyI7P3Ut477XsJXOEx8YM5/J5b2O/qQ
WJRFaf0in2YthNn1ZNCBMGXa0tZ6VuzMa7J9JXmsiwxbezNuKtYRbW7deS5mfEfcXJs/sYRg7K4R
y7jZbBDN/a0n89+I5mES+JMlteibWDbvcE0b7+mWDKGvxUXm0K1retQs1JBM8tu10kJwhe3BNZPV
3jO2dsRUXTxPgFOM3dy9TGFtWZdKrrXX0/Hu0BMiCXRnDMrt2sMCPrOyvbErXVR+t9xiM8YMqvjq
Ya5GRsasLSeF0kAZMkwaz43f0vxA/j2MH12OVWFtuHgTl5iVWq179m7EmJiVBTjAmg0ULf3FX4mi
+JhAVSy/LZ1svAVFA2denBSO3KhoCgMbcigd5c0uFqX633UoljZ7az7ZXqfW9t0RsFChFKPBcDRl
eu/W6DrArRHzK28BpIgWeoy/jp8GmXi8+g7Teg6VE2jiWCjkCAOd/7laiF9FkJCAy2alPAPaQRIc
5zzah5l/KeZt7P+v6J2wShXxF0NBaSRDXhMo9lT5hfLZlh5p6wIeSSztlfcdB8att2A4FnBG9nYb
ZvcsH55oKXArOBHDPRG2O/BexO6BXxrC5wR6sv5J8n1b/z69ta6DWCjBGkAxo41SlmliN437VYRy
WiN72wA9WWBSZpGo1blHfXkuo/kCaIiz7Rw0CSc1MtS4qIUhhCJ0Kml2fwOz492OSKYvJ1R8BvK6
U6h7pkW+W4dh8dVODelv34fv+7HkyE8pGovZrN4qyYO0Yut99SSjTCVvyGPBg+rXa/oHFZ1lNZGy
l2UfwVJt/1bhPmqPz/qj/72rM8xDEnAGP4Lruk5Z7aKBQbm4DTo+TD+mwJQZPASB2HzahCGK9UDR
q6NOKzqNhTa5cddU78vMFZfbgR2mekt9jSZOPmbSipdxhvKqGlptCHmtPpPDu2sq4hTxxnHfofnX
+sUYCY9Snre5M42Ab8tjdqI8VzrSDchWUbvZJh+VkjsittEcXN/0chgh86EeIKbyNVZLYZlPYPVi
qfm7Hj1wsGBSRO636Uhp7kyoc4ioDjpGqlC41lfvQiwXy2Irnmdqel3Ak/2krbi0ulp54SR9akew
7CU5MnPq0DRvebGy4TBOZ8Z9rrXcuJvuN6N3JEnOvmZqrI7Ze4PI47gqDhyTcJZVZdLoblG65VO5
O8f0pQ6kZqSNvc+GUWm/9VbJGeoE3SgpXiw4z0530vF+mV0RsFkCVG0yH++AO7H1eFqqQiO22ScQ
nREy/E/rp5KRinLVuRN9dClpeAINANxfi4d8l4gkdHAZP/7pBKDLErBag0moPAwM9Nnu831be2Iq
NIRxsuigWK9CN++DbCJJyfm2Y5iVHTBmrgg+P2idD7hpsQeo26dSPGm20KnPwdhxzKu8W1BaA3d0
dWBo1NLqUTqaaU0rHp3/VoMDg6rKl1FRmnSLRB8z58gJl0j+J0bnsszeF3GlGXJhPFWSgAy4Tv+j
AeCzNz/5XJTWhZ3rPTsXy1UuQhxxDteXqEv9IZ9QxHmvdN57tj6W19kbBXdBob2k1O991nGpwzaK
I7jVN8D4TMv4IA4IzmzLdI/puQcGLmpvnZyiieGErx74mc8La+mbOZuQ+Xd+uOgeFgY2mGaU/rw9
FUU42SryB+zzHDdm3vj6FRIOtEfrRoPRQiUENGIn77eV+hw8J0zzeri4m5pacgpql6gzdhMaTmay
uoSNufExmLqf/2DXPF9b+Ecf1/ev1/SAZItUYbSAuvCAx2AcekBJKxLT+M07pbyHnHuLnigTjJdg
QZti+GztskX1wcbIKdu/knPJnzqPjpumvbqY2FiOzYpkZX3b7mhr6+7RzD0wJGHwKBTcqptfYW3O
WKPwK0/N7h0rdU7UcfaXYe//UM/JvwTFilHIRKCIktXLMVjutGoJ3ihm9CNi7ksNSbyNsJ8OlKUn
mdAuj96jEpTWAhCWBaVHmc2TgFqMazgnLvX6Kt4ZDDj1eHYyd9DXXgFAUhSyH5H4PByCgFVraMgI
RU8TpeYoBdxtG/BEbg+PM3BtRcVgu4hTLjXY//RcEdAQQF0yBK8sqOrmZixT94QDX8K/mcQ2Yhd8
01LUOzkQo0770/Vbgw5MYMrFoxJ4n2IjiHECEOHXcjqy+UZR3Imbhl/PnZnfKdUQbaz0VrADgybp
mhGz2CASIYXeZG0CIEynMv7LBL9+fH6GjB/nL3H44l1PDgO5w/nWCq3Gej2GxeKfnfMxUdcoSi+T
RIZe7j+FQW26yoDZQMj3D8ibQnSIKa/qNq2+oDZlOB2MhjP4BQt/atcXthdaE7jycrJS4y/EO8tE
eonNcbPlobCOMoNZLjDWMol7VWKvm+5Am8AGKHPcBvpM1jKrVc3/NqOiX0pWnW1VI1xqHlGSQNCL
unBk9J/GZ2S6ATsv2Euw2cwJpJZ1HZp0ysZpuRid9sZnKPw/gZ5mBuUtk2l+q118UFQU6g/87DqL
iMqGU8DMLAFkygt2uh7Wr6uJb5J7rP4s8uSXBkscNBPU5BV3bHbx4t21weEr+YVTn7GJ/lt0nvwm
VbsdSRLmJzIXlqYRv4gxzYZDrH9YNjaqp0JrDN9we1wD4GJR8MAFKDRgmdRgrkCQ8YLGun7EP8mu
lvR58pbt4Rpb4h/QPLqdaEnNHUrEfunqRFrITm+gKtYNixSefKZTZUwzZvtUriyIJgeGQqCBiIZb
ID9TGqBNK385MrDuo8PeZY19bbcS3KBD6beJD+HWsGqWm7FBVYTr+ao9v8Pp+nE8IIfiEYS7RfiN
mBiWK8+AyUIec4ogtu9cevQZ42ZJNFnNDSzjpDQRPnQFJ4sUNB1egvChu9+B5+BnDqnn6+fdEG6r
X9WklDY7zkLFSQplOrRK6FGNRlIsxytVUnV9Lk29DntdtEZ3VhhcNHAkVpTo7P/Zd9xMee4DMzKJ
cVq8PzYJcFKmWQoTDdLPgQNWC4rrdvQJpGD60rcXKOMY4IG1QhFNuOCp5CknPM5JBUAByKuhv7kA
W7LD1nzR1tfptpogmxKSrCk93fgrKXSI2YEGC3mT8Ha7EaiqZb9TduYq0+T7JFPMn9qBJMC50fdW
c5E2bj+thb1adgb+1iLEV8GFG0Qlo3DDTTMI7mNJsvuWgFLfjX/3LWt8gUDiuJMKRS7K0gFQANdq
4JqRxgVWAAPdbZRbUW9ieJPyy/T1pan5FQD+bLbXR83BH05x9nwRc4gj62m2iPM8oINCFC+5FoE9
aJmQxAqCcweIrpA8DuL2AabqjaJEpnIDcVoOBVXTXQsKnhSjTVyWC76EDCQzQbI4mpDkkrxvO515
J0le017sr+FvyIz5muHGuUmDfrXQGE+Y6pefuCf8eBiJLVbKKVr0rM7Pl+pHaQmvqhraQCzgDENe
9VUJF0nS9AML7F7H2Kw3P6mLWmvJrJ57TNNVtudtMtAOX9YiocI8K/e9VLO4XaGOC806Hepk6QmU
KBO6swnUUPJVmmnLF0nc6tzu3kSKmehw2eldhkkGAReS097DckpKiYOh/D8ZikWNUdh9lOWTp9NX
1IqVFlWMJJ9TLmm+QP6vIjzguuXFD7m5T5sBzYTwkVFwtqM2jOOHNtxEbZUuOEfVh3B7AhipNgme
xk3cMU/rA6lFvhqIca3XabLMApN1Rcbdlk5xxXRXq6ld+kl48t+UzJmQjmGXQaVQHDH6qxu/VGQY
XpB2wxvMWUefCmY8ejIJOSzAUInY5Q2cfjAE4UQuDT99CylPB+3B7WuWcSpn+Jhu8Le75Pp5ebSh
Vu3f+D3OlSIZdeTRAbzxly7UcOr4YMh0Hb5v4KJGXH78+VOnoezezEzzO4kxpi620UUo9wKd6KFB
HjJY7qh467r6H6G1YtQ9ON70OST0v1wDAFSNRh0g1Tv0o6pojowrwgLCetZ7D76PgdRgQsVXC/Ls
U0z+muL1TaeO1UrgnV5cBWofLLR+Qmuf4zUbvuc6oTksrrVRdKKuTIqohuSUwOTA2LMp/luF3b5/
+Qe4GzwpWKLTFrcSf1jemTUXD62PZNMXTJ2zoQmaONzALpH2xjJV5DhZjE5BHcrtY/mP1k5IJNwQ
K/hwoEhRFlF8TdLbZlSTV9YRdXtOmrUEjR9e12isor4PyiyyHvsD6kgEwuRxPtGs2CIFv4Zek3xx
5O8A2h9NEnQs21iRjlB+DI5roXKMtzVQuatGxDJA8Z3IIYPjjcvZhoH/ED3XkHOlM0vXE14qABap
qWvhB/4IiM8wR0IsbCEh9l0XRiwk3IHPsp17emoWclmBtPXnT9DgItSY2dnqjICrMudb2PhRgUqP
dLWoGH2OUzwPV35pWkmjhGR07UgeyUSKRbZB2xEldCCtjlpR9VYqwG2n3X/bi6S/LaOoolJuNZEU
1oCUzo7xEcqr3Xb8FVzVni3afYM9Tg370ol+mwXVR6U8QNOhh1f8Le06f3CNGxagflFDPCG6X5En
4I6u93KrNm2BHtXznaKkMTjHXiDP7vBTWwa0zIKau5ZMoJphDeuUl2tyPstvblZvJTEskMSLk903
fPdhAb8dvJqDEocUjsJmX8soZm3NY2LASa9wQSvmzwCIB1fj6itKcbGqKUyGaZxaVESeXYzGLmjW
S1QzFq8UHlcaqGOJTUpIgcJebVmnatmL7iPLWLXGTghsLBBjTqjbK5OVOVxpYJmYhPNvMFbsfDpr
P3qQ3/UgPN2QQDGs7pPXvmXuBDYnYcf1uuFmGqTWdd59kgDz99eJX4WBvm7PCecz0Z6q/tqqX8z+
6e+60yUpj7TgEiHnx79s+CgBXIRP+Kp67SoOxjIv/eZcxXH4at3zf1UXJY9r6zhUVijqI77xSPuI
6ys+V78P7KhUCB4r8U17DsDKnegaOwFRcn0yQYtN4y9vqXsZXcF8YMoq70BUdzai+5VA51jsw1Yl
DPxzGLStx1OFAvd+cbSMmz7iFCM6JdCEO1lSBHMlrEArxNMGnNSpLBWhx9zBJEd892vIC2nX0K/y
0eJeEInk6XYfFe29g2QBNNN9+SCEesQOA4OyWokK4YHPOJ4yr+tGTlHcVzTtnizwCr1HpRlEwZ17
cqfkDMpI6E4JveYl8rcHxvn9gbY29F6laLnhE1NEBb0PQgTP/sYmEktXi4E8A4BgKNdHgVuDR7oa
v2Kw4jTjTA9YZ2lwK1iymNc6/rKU9M7HQRS4d5pgjFx59QbM7oejObra1tBW3QgOKCL667lterVY
aASEC1YinRMMO4uAaBrLk9ebfvotUA6p05mir8VGgXvx40t0+jh9xSo1ayU5U2FHy40s819fOX1V
vH86j26xiIj8vop0F+CRh2CpVrHddnUVCfeGmUXpudxFQeNefJOZeMftxbEh65KZAu63YjVbNZQ9
cl+wPnNLWrhbYy2ptPzC0aWp+P7rimSHDwVuSWrnF0X5mX7GadgtFOtBQn4bBNxwlb13l/DBcrvW
yw38F9Cb07VN5Ayoehy7SsJBbNNGkNzL2LYAtbuW3MM9c68I9eiuQ+/wx0VIkIx07J78HRrdFAkY
U1OWbqhewFgnmRBTp7BC7dzj7yjcFOzuOqR4Sa+qy8wheeEdJ483f/Hg4lB+SKsgHw/BXPXqwrsf
DdhSdBtbG75GGt9vDI+p4nJHVvnPule+ZSyk4Ieae31dYZSjIX4dx8ZPdPLjiTL1A3sc9ZsspJt+
qHe73Mb1AR/Z/mx3IJ3hX+uL5GCgdNpRGy32V1zHDg3fR8DJcUyGrCpTBx0SAz++HRSCz/3dNxuw
HdO/2nYsKRbCSKBpjRPsrGFoYkaDeaE6dP+OM/xvVybmUrdSwJoxEQWz+ZaIP6w8Tn/03ayNoHf8
dVTv7SdcR90LIAT2lf8bkxbE4nH1bUDeNRz3pYYL1xuELa/wUvRO9RwxAqTpyJJWC7kMEyDsDKMJ
lyH6U0He6QFP+cyWyeEgs3AKgvs3VdDVwQGZsuyLpaOz7ZAQ6mdSk/BPuCgZyu+YxwWfzE7GPUaj
EGHPAjU3juZoNAuPDSak10l6B9TpCYy8lRZtoyd2Vo1mSZHF7ZgJcfnbY8uxhST6T8jvDEfWXnG7
UXuEAC0ZACBG9yVjJiPJgJ9edm9hDflTPPYn/NWm1uEVGk/5kDhgGib2QVl0JzOn5R/ioy8Sde7E
NQeMLV3uDJ18aAjZY9hHOqUi8rkFctvFp7c7RUYT+kuYiHLMy0T8sZ1f5E4ZelPNXf4osKITMILM
6PTBsrxjmyYFqE0RwZUJSxwCXnHhvNFLndT6bBCFEtj/uumCQSmZlazx7y2emTnyRvSAGl+oh9Pw
w+TSiIXA5UtjThZHqTpV9IaKWM1OAfbt9t01iIHiEASB971QFg/RfnZPkJUY7KVFgM/0gjiLwN/d
gpubnjJBikmd11a1LeLBHzfP2WqqdWxUlAR1EJ2aHx5C+DikaY/W8gIu8IseUbHOmOagcagoX/3F
ZhLrfZwUfjiI94ACpppYO1o7P8HODrSKEvyezLGsX1L9s0jKC488YLXtKci+5NBm+w5ahlQdTD68
mNIzNEEM+yOFOE8flfuWbTRTzJaJ72aCOOqbyDPEyDaf2GHdXnUKX/l/y4Gx3u8b3dQoMUasdS4i
mO3DDu+Z96ntVu2M6BdD+oCmZi4sFKqVpUkQTb8AQs5uDo1rFbrmDnrmYXdxgK73dO9P8M4vrlbi
f1MjXun5jzBUXH0a1jGY2ybh1RysgLL8fIcxyU2e7s1MwFMnwuLibTarbWV3ju5RYKcb+7cBDXis
L/IyEUH3Io6d8kWS+0b9wjhWa3ZM1g9AqhyvYUrOEnLUnuH6RQVcRrGJpwEpyt+HhsCU/QQJfknH
XULREze4WARccresNJOhmz+/VdFbViJ/bHM4jffTqti/xtu82WqajYDOf8omtOpdC8Em8Vfl8xe8
jL3/PuWMGIa+byGTxTsvFkSl710ejuAMLT2EGB2/HlrWo+dWJr/Y2Tkz0TB43BT+wVnPRjh0djwZ
ZUrzLn9eetoc4tG19PENPemzx0bxSLw393vmmaBOd6WNDpeyY6XSBUO/3HT6XcwUvwOTWHELJ6Io
KB6Y+qbHLuVhTy+xbQilUX0SSfqc/s8CzWX7c46eD5biYCW2qgR50/sWZk8WyIqwgwtPCmDv2h6Z
m+fLlgzvNscUrdgdPL3xtOSvdsxzbJmNADFCja9f6zMQhPXi0lxvYjICQyFoLQUuZlB63RMjwmFU
ragpcHHz8gqwVAis+mNw6ruOS+SF5PpXJhCS/Fb/fTCcbxyj8MveIpM0DixDO2etso6aNBYF7zTh
YrmpuRIubFXOl3xBslqK/iVhVqObKDAoXPHouKQ0mghu6uzu+vT33XI7PJuwX73YlEA/dbwqaL3I
SqJABzfIFi7WSPP+om4t/0sbwQsAhfCVAl+m5M9jDzHKXymZCLXL/m8XUiNKC5Us1Jk5UucHObGl
M3qh114AyBZq0SFNfidIbrckGJnRNOKH/kJUtaiPm18WI83WlS86rmpQjoNVIsE0tbdxzJt17nGj
70S5MlBRF0+IOmrevdtVFUgX5jyzbSF955MpOUDeU6KBHH8qH7q+XabX7vM89yziKbwr6IMIGU6X
45dzulL03HkFOoPCdqPRwdw/qqj3q42jDfHa559GF+y5MyGpK9jsBUjsiwE2cnGqOxKCtT8CNeiN
fAKutLMlo45TVQg/fSff4dfdTsvZzrqP1nyWtxG1NUYeZpdPlSidvxnUISJBNn2JGkj0plZbPHhu
VRfVHpWFEeCK5F7+vHtqxMBkNcyBM+NQQ2sAXKrmzCYp8m+Qla5B0nSJ+jYzcJV6wU+gpTwdBaxQ
cgGV9gIqykBEVH6+ioLMaTdYK/GBxR0QJAhDy4crc8anA5OsOe5xBi7wjLGYkvdWG29TrIJRP64t
Y7yggTT3UZaN+l/9wj8hbAnXJHZSEd2DWkk/eOaknDgG22utualpk8txe8K8dcpybndPYsdoxOvf
HvX7fb0QX+kUmFJJO243a1HxX7T6rwXe/64GpkE1OTOqBeGgswOIK6/n8ohSuw1KS+jDROVwsu8w
VAI6cD7KYGgUPK6pihizu90WzPj/NIGOdXWZDGAu2JQ/xEPZPa84Y8+auFjcFg7oX3JVjQRk5mnt
5PkH+u56WMOkIlpYg+xHjn/rt7LuA5cLicppYtmubqA/HYC4iNMkQqEX+jOQBREpwLbKF2qWhoHb
qYYY3UC+l3/ZBGQ98ka/RCebGjm42CCce2iLYybR/CQKYYWv74VDXX/HP80GrBW63kuObZHNZp24
yZFZsc1OOHrrLPg0TaD6RkZByfCQ7Mb06OOGuklHoUj5kACiF/nGwb1Xh0aKdeRlWrn7De44UxVK
zt4CMR35rZxFY1YeFMLPLmCxGDHSVZEquhkReZkabG55+mMFlKkREx2b7xbKFgBORim7L1z74J8D
87reC9KBiZLBZkNDchTfZS3018mTTyJG1r3xXcKcsTbxcWos6i1JvnHaa+u6wAxox+Dii4Txgjca
pFOW/R37jRobFWGnGHQeGHsH1S+XNn2VKRd/Fv9SppkXV215/pB+HDfOQpX/qcVc9Vy+gkjS5/5S
q1xzh7xlOP3Y3z5ID54RSlP3+PhWpaLFRyahv/NaDnbN8ToUNy9G/3Y8BehRRfQ9MMX6EjbIYFHR
ko/sbXwXb7W5ox62pfB20ZshlAaRTwbJFhL1nranh+NPjSBmkA28BBPmD7Wny8fmYtQ/Ybq2W4MM
o8usKRSxu0lD8miZpEaILxj286FjukJj4SXIDBsYiCn2kXZcXUU0kdJOULol0VXn8PlkqpIXurTF
smXK9nH8y2paL6z6jpapB0MOCBOLDRsN1j/cP/23jAZAwamzh9h1ekTffuxpoRD2dpSHSeo18UYX
nvVQOMV4bf+xfhBC25vSyUTZGeEmpyMR1W34mvt0vbwE9xmwJFXfMxGHqKxG+ifyi3Ld19VLqfdx
qpx7dC4POiBQdy+G+Kv7bbmeAQvI9zUEyeAVNfKfRuMJqSgs8+QC8fMyYJeKSDe+OCdA+CXBbYRZ
tMc3+ViL3Bf8LQMq4gnJ0kx9CLo2+6Px4WtdBER83iaV24Mi7jj8FysjCfz8tFV4Akp/J40CpEYE
u6Nwp/AY76P6wk9vJeoSunNo/+W8s+Tmc6FWvPi93L30UmpCVespYnFHwHd96zdmKFPp7nVKzYcs
HBYWgnX/bbQ8l3QhJc4JEVaZydYNHi5lCZTjy3bDiuoz4P3yQ1AkoA3h/FMRylSCmRYDLelLwtnN
bZakqiTQGEhFCi9abh4xI2PB3tx6EOzPVA/HG7TAjvqTD8JcPz7+JHTU6trRWqtt6zz9+eyQ9R7r
b8d3jugN5SCVL82aH+Gli5s4VTI7W+AZqhIiTpUAC3FSS4/DmhVryHPs3A1thTCSrXc1j7fv8Nir
5LJDxeEWvp/hmwuUijifcsmf7XDnWTcK/gcn8RqwJu7D0xuK4amztCGE43IqQkQgkgEya6eoTdJg
3aX+CCkr174O9qc1eppoqEps9KAhRnFwypUiv0E/oEVglwCimtQTRuA0iHZjvH9Z9lIqJcnBxvOf
KGT+YvJZwLJqM1IKEBHt4xIFoN8rxbbxLviLVFwFRTR/AhUyXR6ySDYMPwhrMRHFLnPB0HzdzoBQ
tEoidv/89FhWdGMklTgl6Cj8YXFBDT1eT4ZYHhJPhwFSaw6PP5HS8rMsup27kooDhiEt0ffn4lDZ
WZjq26JzjakC2aHTHDFgN7rpvoDNClrby7/4sQBAkGtx4K6rbJfCMaQBU0z2fMQUsAGU9VvmVPnK
TlvOtmdUM72OX7bfAVKJ/KmC3kd39Gjm5rm/tNuI5xcZqru4wluxrJs2nQOA+M7fGi3mDNiz47sU
5li2kO6rlqh1/7jTKZI1lHYAxAIRhBBB0TG1IHq2N0wQWsBU/lqx7qxqL1gYcf9WM59pnMUcCDcN
8+6f4En8EyJO9RarTAMxjiGJukPjB2QQQlZebbW/dXcg3BKjJIIdz6ndxonBmVT9IbVsPNeZbb86
glPZT4fAaFVO7twA71/4LjwLR/XaGvfXou0GaWtQ1q8NyVLm3qgNkDqBuCpuhqXV8l4l2Pn+mhC+
dmGnZEOoZgoj1eIPBxcID2bSNebT6Qm9CTk5R2hZyvvv+Tfdk53ElXJDIPh4/d4JlMFvElEqfzDx
N2HWoZYwqyAIqHoU5uux86h7CYoVoayW7Ms8RXzgketuH8/Jm0eM/FAeshS1rreQ/fduODeuUUf/
YNe/EzbJJWkJcaQs6ch2i1wpEEzmQeKjwRjbiuztZBCcll6T+2HvHu5fg7Eaas8nnYb02A9YqC5W
5qczfuQlnp0fK103Eg3nJES3df0s3zrA0SJbzoq+DG/YE+S7GIozeMGGzhSNhtOUh6Nih5I/cPQN
LO6xJGD2e2IyMceo8awkdKJTt+b2KQ3x68GdXZRf8cjA3o2WoZkSsK/irDzsTPyNwfjzjVRdcDrf
Tb7W2yZpEFuDD7LVoIfntJ5QdwdeXj12OBsa6NK1GMRl5UkSeH6JIbeBFaaEflE/JRvI/XZU18KU
fCheUQ8lAXRy20L9hgeHzq3fPpoYQCdYfg9JyvP1nFbNMF5EPgrERiSCZ++JHVLvGPjWlTx1nvWL
zPBMoXFSkM14KPx4r/+K+KJh4i+9Un+Vu/nJXPg01t5H5zxKVyixpMuJie1zE/lUg63dV4QmZKwA
gcSiEINBunKWX2+N4r9YBarpgFXM4f73eQtDAUlfHIowUMqJGYa53PHBhFYysTE3GxQO1ZkGvJx/
RWypHLxY4ubJrCjsfHr9X2omIDcoLql+Hz+Q2fnlflmOkol2Eo6/GeAoa30wLzl+pkoA5MOnmmYk
A6tEv9IANdvdD1S6VbXSXfgAyW3Ew+0bw2aENfpoLApk+D9DH6MAUADhgKjiDuBdC/cqgQCr6CCD
iY9AMd8WQf2p1evGifFk+KCSOWgA8cTz0TsHENrdIet20JFhlDDUwEGHKwiI57cdkC2mC/7r/4Ns
BHVbbIfFZUQU1TBPy051uCsCTaLXSfQsMCtaGMTVghpA6XlGYmMXKgF98PDFkisBTsFxM6JX8H/I
0AiQ+eb2U+APfJCFh6I3+2uYUrk2Dv/LDyh5R1xw0eYUgBpXNukz9xjD/TqEDGQjCZWHREFi+bqm
FoDwrwcLFEbboHWvnxYXGuvKgHbIl80mBkA0mplfUSMyLIGAm6EQXmI3nms/oHSR2Ov+BR2CLhXI
jDDVk419YIQBZskWZwfoseAQK4jhGrCtgr9qHX28FujPAahExcerTUAwZUYIU0AM8nj4nkgA3/Fv
shK8a0aPGobZgcDFQZgG6AN/GCezSy6yukJKQXGJRZtG4x1fDjZ3UgtMoxS/gDbFTxgdag7ZjXvI
k+DqYOqOqDp+CFkLrNEMNaWvm4YB5X30kjzzbtW3CqWp1rkixTQtkV4zv5KF4wdkvf+XbePAaYwb
wcN1egT211ksnSha7EVeeGoeQQqTB/6kle4OXis4leEkTxZZwkIFOW+ErKp/os0xG21KtGP5Qnis
u1rhhbzWNqQkJmSbtzTPZBjqXbZr1neL6n9SyhFJbBf9pnaU0l/l6s3Idxjm6sfACHIb6elesfaB
dNpmjXK3sYgPboVFA2fcg8lmbL7Z1QIxA/eWyNCXPKBoSjotaefvx8s1C2ztf/K3SKegmETXt9v3
GlxhRX6Gld0xxNcOZ7sLJcUrJQCxAxW9tA3REq93lET0JF4/co1TNAvAS9ZvLJ7F2Z0FsJn8/ZZt
7TZnqoO6y7iZ09AbtCV28H6koG79u7UsgQiAvvtko0fKwO40HxbHYlm2A0TjHLkxWrxM/IJAtFru
LaCdTcmBKK/O8YpoA/dgUyzY3LPovG+YgvnA3TPwQvzw6Hh8W7AECfWvUH8DGhkP48ivJf2x5DAa
ZcwNSbGuWjHi1gmbn/U0RwpGxZ9As4ApRrphxJKTkksMcRvDkG9cN0bhSmL1JujTE6rhXtS+HekK
84tWyi135ZGkSnLLbhAkp0TkGSSLdfDW/r23C0l1klKtDaxe1Mw3r11jnJTOJQ+XAWcek8+Vel+X
ZJhEqeMTfY4V8Oa3114izAt+LRzF2dKFZReij5OBBwI999OnAYISc2RVwEWu0caKup7hmSAIEKrZ
oQU/UqZy50EAUV+GVIrJM/rB+HSPerGYdUltmapnU+ko5rzhLG6mLshmW4enk1IyTM4q8BD7xHoj
lbQYZAsWfZLBRi/E4fVM+jbDI7sDlsjhXtD8WEQi4CIn1bzo68RbcPZe2JjWEfQggMEfSX2Fs5ln
XHaPvkK8Ypje8vpPG54scIoAtp416qy8rCcqYgWagz9MOK1GIL4uInyBXDMtfLQ1Giy6LVaQkYVZ
oDOh3g0fnWBxjrSoVJfvpNZszUoK49pDNZFsHrRGBtu6NdpgSzc0kKrwLVDNmMAJHCNvCnVk59U9
ZM7GPMb6hIjsTbs18C40aWoYCvvudrIkT7dqMG4DOFV+xsnSd15DCwJleHWW5ZXmxpewZI6BTLXR
1ZiMUVwYIAxOfxQ27gD5qu32o2IVLIN2+S+sH0I+BTCYFiDhyY26wrYgvlBFHwqqFw9Q5D007Rsp
0dSZLeA7mjpID/YLKG0HKvG2sXIPmUuJjcdXSvAm/Mxn3g4+xnrhGHmerbfSUrBA1TyOwGIZyOZ9
yiAa+ysulqSlL8l9BY0ntAd2TiHXc7oHM7GJBEa+le51xIGjtdqQWuqiEdGbZkGKo/GrO5osXT1R
S0bIGM33sKCldAg+duH+NWgMcO2Fgpk3SgBZ2fIJQ183Roao/OAhNFHMz+HNeCSjusV0EA/KzAnP
xFSK9Fl/War/HObY0JFFQ/9K6n8NlOuWmfLV5pLEzsTm0DndRjLd3AUkYKWr0Zf2Z+/wlcoZVkmB
ItKFRG+g/NBwQfCvI+QkBQuF+lUiW2qmcFak2rKrRHWQqeo/SQ5ScYau+DRGoiGxRadXu9M5hQ9V
vkoeTG+zRvHwoVdFYJla14g0PQuAz/w2dk1YtmDYyd+e7nD/cCyMwK1ICbD4pZRAlrRg8e8YwYcY
1xmpCgEvQv/O2O+lVaCLE9U9reenz9lPF47tsnrMVhMYjdVO1GKIzpromF1FBKQns4Gq3RwBygl0
6WQkUFUtWug8SkDrQt6+rNTMBIcdRTppqsP0QMxYwgjWAXvGIz9W9JJSy9PIo+UsLd4/pjV8dZuR
4MOMc9capGSX3MvQda5BdBQER+2DfMU1bjISwB+xChZb+BlJk/BPLs4qzcze+FMyBLkAECCKFNXd
PNa5LGNpUgQFoLD9oABtg1xp5T/ehLAhoUXKJS7jY3yIrF95k9XRVAA4K57sTNvC97HlDldZ0NmV
XmwhBwiF0LnThflLDAuaATzIBbvXB5XWHU+Hg720o2rn1XQKLbpBkrlrxz46yztqh+rBz8hDLs6d
QvT0Qrqas7kho3extaGJ5z+xRmF4XOgQK2p4Naq1lM3eAYjVxS80o0ud5rDJjgCfzk8dWwl/F+HB
AdFjczgQv6B5JU8y1ATLe3RBdkqR5s6EfOFaYayL1LOWhZH4jplx4vzbAND+EUCww2w8Pl/IGMkd
pRjzdhJszmmtaRqOSLya31ajrpA0lrKkv/76WEVHLloLXVlmRPN9P8mqfuJz13xrTkAMX6stGAxh
7qwQpV3DV79kQJpnP4F0+ho81KfoYMxjz5m6ajOBmyCvDu8vH/ZN/LHclWuNjb0IP5CdkktXseZB
5S7mJWKH0pB2RD2SNvZ3s5j1u2Z1lIy40PvMNJg0O23vB8HnVBJdXg0n+8nWsQYrCKs+ZFrVTtu7
D2fcuiWqm/MyHVdENmFvCWPFBwW/d8MpUYOkAZ9fBvvxVjDDtuP+wOr+1c/F/ovZX81vK3++9S7j
dAwYHmN9FWj2HwRac8sWSnQCH1lSWRS+uoFFhcr/5lRV34TWf3WJEOKcWN5u8KyYXGFx7b/rbfZc
cr0ujt/dR6lUFG52cyE0esKxvnqD7JK79ega276uQGEMx+QWJzHL4ofP+S6ybhXworlxKO5OVS1r
z/dFEg63bAv+yFiQF7N+Wp/TWB4YMrUGH6eWzCN6XP6pgVewBH0j2xaf2ejvFOoJzicKc2UFDwCC
sEnzZ7wIUZmlnH9bhhcFAVzmJ1iNv2OTBY+Y4NEgOBcNRuRLjWGN/IyamNRG4g/WA6wAbNrE/vbb
Nyr8C3zagHwEKuFiL1QUTr0cAumFmcEh5dH03zjISUElyp60zsN4KnZ1vRDfEqi093iZVq6RW7lo
zbGHnf066CVVF9iHHbIXVFLl+g22IaeNJqRQKQcYsyjNPEWJuDWt7k3+qOVq3PFly8nSA5Lh70Kk
SlWuJQASjP+ouq/AQ3hFQ6+F3b8mxUyoUjG+h7v9fhPibsx6q+fiN1APSRJLxEyVw4/9ggKUS8VB
jVX+eXTLyMYHGQJ2+XXrAaKFqjmVsgVP4lVv1x3WY/xmnSG+A/EK7SjZ0UX6QFyfonSzOcSe1ceT
vL2ufL02WU5ujn5vzPRVQjo7Erq1r0iTt4zHJhl6AHRJT3xSzFD6VGo73Vr1k55Pb/UqLO4hbvef
33+XYOodFDIU4zsSgL8XCYflxCkmdu/v8Zl/v/ICl0PCmlI2SFA8adnL4fVx3Q+OIjDq7SSVN8a4
H1pKvB3RgOIDlTpwh3OW+cd+foBE4iGdFf2NFBp3W72FnJTuH0ewycq5CUe3cIu0Ml3MxeC1WDDs
SHohrL/Ro74VwCa225WxMfEb6/Wkdc4zko07wA1nVt/i/OKq+LyvOpGAdvWVgZcRGQtJwrFxMEa3
m/bgNrq6Kld7H9RzhpUM9HHuKaaq8Ktf2pbzJr6Yl+Qzz1t61gpCFYHRE5T1bc+ZP59VVV5RlZnz
Xd+PLAaYuxBZqKrqgvQ1xu+b8bNAFJkVvEqfpACHFBejwFJAAHwTXyRk6Zn21AOKTPSR0xmCmlr2
9mW3qXnRpS0lXBUHal7D3kQyquHK0eGaqX3fWRvhDjAjxoBT6tMk8l/lTx6T8kNe6zMUjNCGho3W
8zd4WerK4qgVTxLYvl34pHPwBmNQDp229/bRJ1vzcHJaJyjt9O234tWR2kOetuw66RxwZI1nQHC/
wQ2BKCkLPFlmAT4IISUd620EUpVyDFGuMKJTYfF3kGAL6xIVugNSUe8yTSgUvZ5IhkbZqBhQNvv5
5wFurkX3Wod85/XgU2HlTtyw/B9VYvlt3fjMRjCV4UfjceIKU6l49+cH6Q2T4WZVbdV1N1UFiaSR
GY1Sgy32QpBav29fjUqoWeT6Ixa5OqS9105K8YM4GiNO2w/+ClMvFoWn/6bs/QyQKYKqQxAa77LV
BATqwCf0e6ADC8/SzwvQkoaA22OIH8mOpin3v2TGgIZBlIdYmBrGPofxY0wJgf8w40+Sc0UZryu7
hSYOMUptgjZQq6Wz/PrPeqsjiIBA6FeuXtnz8b9gex4DZfm2QApa6QPNm5sesfmkGMTso1peQVti
hcVA0YduY+ia6669QQ86lT6vMwO8a+Iy9vGRSz4xdMZziE8rOn2aU7bYko2Cgys/oN97aZyj4fE2
vZjgmf84Wc1+WoKdw2WneIdF/KpJiH8yFK4AptkBYTJA7jWOV8WGV/Jcnjou2blhA5a6dd8Lzzh+
LgsqIIpMuGEy/iZnZfU18Z3/gFo3t7nCAIMiplyd2KQKDZyHJdKtR52Q3lo9lA2B5pVAwVEFrGyu
l/3vzi+WNib9M6uO/PvQNn5/h19N28CSe9RsZpzZBtEEg24NGnWOILBdpmf/x5cgdqLLQ03gtEtt
Q6j3C4wA+PZEa0UXzivMrGg28kZmFyfLX4Z5Ke0BVF0D2cBSi7g1i7ei1GVr46lFoILewA0WYnBO
sVQdIUk0CIKqDqvG5FnUkgqjAXsOOuxi/D9tnbVbW6WfxZ6mlF3v79j5vHzqV4pCjcKMPVgzDCGH
DTy9Fhy6mq60uOpLDj4WvzbRbtYFuyfhpTc+6+4K2sc7YwEA5mjkU3PF5YumpSMzK3RtYe/EHIWs
P64HLfnD0DSv5+leyb0LH4vJHquJqQ+6qzSOJmHlI+TlXopTdpDz4u9Us1Rpsx90wuHwaJAHKwH/
/Pb2s3BNhJamaCk7gd+uy50crrASEHlLVqtp/5jpGI9N5KIBXCklgLG9oRWEy1S3P+cFY1PIxksZ
8+v4SXuSLvkQqkpgdhsVMbf77kEoYoxW/i+PdxFRBpLzKkYbk3/NvvpJVU7x8XLknohzX4BiTFmS
EzsS+ZcP88w4gepApwauvxg+9yM2aDDHcGLGF3Yo3FiiRh6TIuYbOCbk4U7tFFPlzPIaT9Y1aPP2
+KoNDO/CKJeM4ba5MaJA2FboxgUV+UsG/fcuzHEKSFAG7iNdqBgsNalkRO/HtU4yLnl3H1bYiaJe
Rz6HY3mZ6T+TD6BBmbuJZ7CJDpE9v3UbfTRgC/S5PzNlQwTjtzdIyQkVhQyBkiZ2cchndfjCttOL
veG0bAJs+c8x/HZMOXxN7WR7Jr3OPAJFMthhpxt4AWBsuD1iKNUjFRVW+JKDYQR91zqOZYaioVeu
mb2XVA1UPNDuhhp80Mklg7x0SyMI+bfIjRjBQnJlAF86wr/DuiM0/9LRk7lRBwm420lhpGh8Ql40
W4VwN2Mdt4CPZmCy77Wt8pq+w3aoOqkxRQmW5Q1CLP429A7/74oxnDEoca5DdlPL2I2WZfjLldIV
N34jslyNOrh0QkLuhwEdgJxpvGvoz4z+39NoJjaIzRrWIob2PmOtLFAhTaEPS/Wz14mKRmX7Ai9p
eWVgVjXIlqdfH9MFPqCBy6NKao8kellahDGNNNp97kCSmg1fwZ+fU7mnSDPogqACSJq9B77WnOx7
EJpUEXJG7is8s9puTt4+jH2bd+Czp3AlLGxeJEZO0KH58x1DlV3X6kkUZUYIQuewJx/ttJ0wkjYA
JFcVLcrJ7l128utRpGctkSx1aZU/6XOuCO2ZOCPCzvFtJcVLCMOkd7+ljfBzB4XyhI70VMzakfJe
Hd8vNvNeWAQwr/GYovQCBUzk6359XD4Re2gMQxeEA/1WFJ2jcucLCX2Zw57puSaRr388XynWvZe5
Awq8TckNDFF9eBeXmIqIcUOu4CqU+erKQ8lyxj/7klTypfk2gxb6JE5NfMgt4MIBtbljmTcSlAiK
47O1k0ywbbdPaHcGdNYcwo/+/1I4OBpvmJm9it0VNQS6BOKpl7JcnDkNsWC+oCY8I9LWzfzh3Rfs
uBpcONvRb8J1KHFTcBQOOxDm+zN0J3RxMaEyPL/HDyGUUuxXQ3Y2unMDDaMybtaISy4FBCOanZJU
/L4h1r5slAXQDoaGRMwx4lNTgjfjTsqunfCRKp6SWUJ7wyuXaA2Lyskb0SFCLqwPRhO7Ya1EZrsg
LqzKRCWSdc0Z7hdEUtzvHV4MUcBKsPKuMom8F1RB3kTE1tz8x9lja8Pp1qA8cL1lVxHfM1B4bM3q
+tb0a4CzbGk2gxocD+Wzong8XsvUkdGWlYEpKx5UqJ2ckcFPwc6jNmRSLJIOeWQf4h2pI1gMz+gO
0SNQ/d/ChDAicovKjBJFMiDGDi7nUaRUUuvCM3j96clNmNd1R4xRT/6D6BBBTLgkWw/luSHeK5LT
n9jKuWnxpLPpfQgUtOrgwh1WphgcqlJFLY14fX8VC9+X7tZlB8nwEDuC6ZVgi0J2pD07XxWMegY5
NV/trppc30XtmcdbiJbS7wYPTEPrRU8bL/lgyTdPppUDpezJ+aFN4BjiVx/9Fq2CkSrYH1XOMUny
TDIRdnLj2g63dujJUHw1VmH1e5IRTSCwSMHVezd+z2/sUA/vpmVVRsyT2znq0f4p62WaZP2cbFnf
ACq7MrOhnUH8JSXrBx3zwyKf5/THbHLiOk+DVg7Hqa9TzbA31vSjdh8jMcTapFvOSGOHSKfsut5c
Sa/xReTo02pwlCKiZbtmXxt+u+eU4q2yzI8E1ONXln1Nw4zn0Uo1E59ahljF3rzmadHHZWcJURXv
3PPg0Nq/IYWjHRv3w6vVV4m0YmF1CDIiu3iM2yxC/6dozt/X4g9EU0ANv8LSvNOLsGCNzmAjCTaQ
7fpotFyuAtk+7gMvdMFhSVE81ha2O2/8TR83XX1G6Bf9c739neWWSk6amhQSGQ57gz2pNUi9XaN+
HYqhV6sAFftSLc9KzZgjgONtfcOTKXq95WHxcKo6/J6H7dc+J3sH1JPLcs4QAbg21VBGx7vL0LBQ
g4ErSP2hY9zpMGdCDeND7zC4ZOXZmqVk66IbNpFk377vMSwlfFkHl22rAT0P5lBmHTjgwuLiH3a7
B7RH8quitHV7CwICjZMfO5TjPla1nxr0F4V4j9TLjjwKjlMy8lw10GWyFmAeSPzDc9r0+fCZr4Q0
vW6qBWLU+zXvGdK+Y4GdiOgKki5Am3kUrsLRjbX8y6lPS9P5rwS7mWjjSNFKlbfBjOPbL1Guqp9q
ayjEjFNoQaN/k9q6hbyH9bs7eVOWP7N1gtvpc1EuLeEWv9OtcPcelVuh1/oicn0uEp+rvZtcOqzd
dbKG8u3UhkfYKsd9Ny+3vj3pOSSl0TO+9o9zccCvT0rU3xfRn/d1g91XX+XBnfImsPlvYn6Ypk1q
0V5ce3k+z7q9558P/b6SxVEIVAuwuP4cx13vhzaNTJdW+5jrNdAti5HyzfUKc2WttS/bQ3sLAwZO
X8kvRIu9pyZ/5573AJkq2FrO0A76yba2FIA/MapHXO7VnlcpnwakfOxF1NrqY70I5b0jcHWq6P+T
8h89jq9mqa3iIRfQ5mYMZlyChN9ki7aS/QTbfQlRU8LQ1zty/CDgo8+PNoWyDKO6Sjprm83Bg0XE
bNs//KXM0SFlRLGo6QDCOO2uwcOmZrzC6VPben98kzDAKupOZTs0yUyZIPEXSlH4P31RBcHah0/X
c7HpXAvaOEMpIxec8wi4ufTWKyDOSLiR0kVvFI7/iSteLJAZUOwTzj+VsTJbatxcAfPlvxINrdzW
Ul2KkJ8xPd14+PCEi129gMKUUoa/bdN+/tKS+fyphHOU+rHwLNypdmL5HqCY+oUrK2TNBpcaWijM
AnJJhi1eJPGFBFcCdo9pDKUBDW5lC4S9h45zUnn6Kyt/2n4N7FryrpNDZ/RP7OQGc8aqhOmGZDU/
lqbvklBJcBCgcCf6rEgtIQw37TNiI4VQ5rOQzUDOO5rieZxw5vgzotKN31NBtbC0AUagB32UmOhH
xz9yLebAdBo8AR4HxUUvO0uNhCL4+CIVvuiP2/tSRVy8CNcghnhsWA1wp8DjUL5/+hIgoXpN/iyj
KJnGSMoNOQd/iU7rUSe4Q5wg9L/1RFX1f5FoE4obGai2R30unqh+6hNm+O8WZ+ePkrZ18H7/STns
hcG3NOngnJVvhBkh2JQVu1OlUs9GFJ6d8Od37bKFjvlpl5h0esgM1EPxTFg5zWBjcbjGpH5o/Vzy
b8FUbYPGBWztNhiCre4s2xWcCqxLY1iAq/SsStYaRtVZpWfBYv8TWR7peuE4hC8DUF9JtGE4J72o
Y8XbQbqe2rU5HexbtG5Nj22Yc4mJ0cLQU+Snx5RhOPovBymlU1EHgOzomJN4qGG+BVoAct1WK3Pe
Axeq+Mlwv5Pf3IC9Iwt+q+nsPzDYcpNpJ169yqmwJXlIrvpL9tdyqjx4Zn5mFC8z0j/NiNJ1B6YO
F6YroZJ6MpyksTZwuteg9I5GfliK04BD2oQiTEaUWfZuK/d7AFPv4sDgraV9FLdLYZg6cbZ/3pPj
lUlYTMDnpUK6TMTSpGiNGNq6mw4zO17p0SGEGyscvsTYxHJhMbVx2IzJDYk/Cbd5sXqq8/FPsDaP
LdD1ROu9KTDIFyvVAmgFdzVwh3LjJRHNmoxynTVGZdeQmevRZ6FrRX4lDNCqF5EIjDucVY46h8q6
7EVx4WRtWdaOzDNkJdnyAXuOlwkUoPqQqYG5hVuVIQis+wcX5jVG1YPmK9BOPc01wyoGtu09cjWn
UYetwY2qN6BPsjWRHdbuflQ/bbe0zP2neg8zYIdGzLGU57zmztOG3yUrNfmN7V3JOytUQHu30oU5
Pc9vT6PvrPRWr6HcdsZ3CY5V9ltWKFnVXKULXuHxzNFhbmnBfN0ZTSbDlpkm1hq9NCe0oHp3PX5I
WTVRFrP2exw7+9oeKXcec1KNWRLNch44eLGW0C0vFTlxhZSFLF3kpSXACLfPvXBneogLDJrNoB+P
mtChFbtf+lNg53Ny9PcQDSiyGIlp9cMTrRvxcDZ9SfI/MJrKPFFolx6nGCx/7Wr/OLpvtmhJ8zOX
lXc9msbsACXy2uUEEVX1NBo/IVI00x7huq6Y/J2HfokEqNgeBk16cNPLjlQxKatd6PPmrvLkUltE
HyjKZbuVzAPur9WDiARHj1QWfobOCuGJ5Osi2zMUHRuRfmrD/+Isd9L/mLFJ0IjJzrrGGBhMxovr
2cgFxTAhNK8WjL+Pdy08sWfZ+OUh++3YEdbfe4Oi7A8VjB4ZL8Zlt/v6XTBQ5blz32Fa9v2WUKOR
W3tK9zoL3/E/JtP19hH9jWYItxIjejNBZ/f5FEQw8JTaIOiGgKkXaa7eXW/g7WDD2UVj5S/qnz+0
AX2NmiucjotgU6kEPTIWW3DvAntKzxffllTu7PQlOS/bZ4eVRcDT1TKsxZ822lv3854b6ZHefJZC
tcDJOr2tt6qxOdxGka+KQhltrJ0lwC01HxvqPI8z9LxewDGj/A9cG8fi2hUx0lrdhtQRh5kxheFN
FWb5gCaZCBTWzLuaTw746Kir4qoROYpwFcetkb7nfjSABdGv9sf5ugS4e1514Dn57pQKvvIoASU2
e8aCfWszBagYkix+xhvL6MmlZEVAFe0z+U+oyh90vIid1ZUwpH5ZqFrMcXDBHO2GRmbAZBuTycUE
gf9Gva93hH293HLwvAepZEBlaavp5Jvh520+TJJaOM7kvOp4B5vUvOm/MnVT9WBHutgHwLK2lRMI
q2O8ltQBsVz1ZC45JN5rkc8+1Xb0+2ecoTlPgYVuM2/Fea5io9fQ/ohnSgYD9yKRa8GwkKOD+YV4
WU2QjLERfz+lYQ9oaa576t61O+/bkuDsD+T5qUVBPBxSQdg3BXcxiLmk2lZ+oTsPQii07QWkBeN5
KUyMCN1PZAVWzZW8mWypWYnnswWzDolVFgVP5yvhFGxBMRBqAo/9DwC/cHYH1pxIGWEAh+0Wcmuu
bHNBO+G9tqMeD773AMLJb0vnwOb/HZ1vukiq+HphMl9msRsWFrYPSqrjoEMLPU33aA1MQuRPk6dD
4nzsTxz4J6ZqLxX9rkOxk46VB2jxt0L+5H1/hPWsM18Tt6MBslyUARWa+tRDJVDkP380wW4TTUYm
uqtOXHU/5jwS4lMJ6DcwBjtPy42eQvWJ86N/Id9Hy4xF1TuPicYlh2fQXCxn9PmSSk2K4XqCzGzQ
YojRC4wthxkkw8sdxIv9Wtu5c+W5Tx8/d6gWpQ3VLxUS4NfVKSWx4tYOS07kTBXsZUVd6ShhlL2V
MFHWjnLjxI2jiJKsJ74eT6c8NGbrr+JcwHrNegHJLxwmSzjOo4SZIv+vA7kF2g5WVJ8E5IKLOZ7R
GguFq83DkUVs+1oz9905lCOQNr4Oi0KwNB2EYn/gbXlnKK1XavnRiNUYWKhCCQi5JKaokPQ+rN4o
Oad+BcHShsmuwQjxOWB/Hw0nPPPMMvo78xUXjHQKNmXK8H6Ns0dlB2NvBdGyDIuwN8tTJVvVtXQY
gYjpDVBVLh2/iJf8MvyKehSn49MaiQB6zmmtWUh7xzNgU2w5Ib2hnPuw4F1L0DnN7lxH8fvr+2MR
/sfnwrnTiv8myJuK+RpGnCXMRu5hz9pdx31+38TQ987Lz0mvi7PApqwVwByYxy3xwUKpp85aVHM4
LUplMWCQQMzWsqukjKr3neijxgSdjXkthImpiK/9rX5o5EnTuwQQX9EH+9nW2qyFpNJ+ysT+fsJr
ohFf6ad5w7MHro+tLuMGgi9ok8AyT+GkS7l1tPISG9EKOu459CVpBhTI7O97/5CvR1AlPYIuWVtL
nNLzcQSPfVsOZUgpuLHnrIb1vnd2CZRa9PAWsqFDGGUKUmyd1qSTiR8iZJ2BT68GDxc+yc258NE3
Eg1BtOpzwDLIIh2ut1jZZS+A1TIrzum7KWso11u+FQ/Du7LIDniqPYm66Y6hHC8plGKYzFhilLPG
RzTLqDT4I2BQXNTC5ea+tPrhDGMM3RIoT0aJd7p5dSAcGlAj9pQcbujKo0R0TU3TH+QU7mFCi+1z
h+ZmHzuzvBb/HcHNx87WQzTGwpvYz6z4ETB11NAMd/T3U3RI4/TcyDwNUyPo0tH5+6J8AEXdkrIe
1cASsihLOqKqsjOMjZ0DFXw0rLJTmVtfHK/5eW1ZWVF6EaYO5J+xtJEBXUpv2PQYSn3fTipPvNJu
5jnd2sT9gBiuXPer9cZJGybKqSsKn+w5aLp4ZoWfVzh1m2+mhJyVmZ0Xd9LVpt73j7g6npOZzgkS
USnNXKjtF6ogPQHxOh8TmZZaBh3qEBFp30cMUg6gWKhMMbWOZ7Evf7dVJrCVN07WQR0JE/Mqzuy5
vln+wamhmXzqli3U9McmBO+mO/xVvLK1n0nqfKhSX4qQ43YbwQTZcEXAe2iAOiLrAEB9B9WfaZ2h
YodseVI79FkocAH2KBtrt8x9tdlKvmwupkKmzZs2Hzz9c3QujHDgcd+fJj6zF6zF9OSc1zC2CBDN
5V/pg9Xo0aj2LIiLxFVJLl8NFKWV+HibwF/Zxjgmt5HcFcbemf2QfQaKDbcVjxSPaTDUVjP4aph6
+0G21h1E1fpgh3YCprKsEWW/QghOOQ1mbpEI5PXTA0gl5GilWV2+0O2utHQEC6d/ABbwHBuczBey
NwEEZGKdGqMHdafNwkxSpM/vO07U4+jlzrKxh5VSHEx4A184dUQzpspsfuHivLgkWTb3DvSzXKEv
O6tO1nlwWUbKpS9XkUQK2hbEteJRNEJZosj5K3EXirJhexfeKNN9ma8sKqGBZvmDSuh43F2Pj4y/
bcsNRj4OL5/h5+SQOdqMm1W9YBLBe53h3AsruCCuzYeL1x5f39iiovzuhNQ6h+Jcp+Wa4/X/UvSI
Z9ru/o1MMgX5p54rgOnJlzkWNgLuww2amr9Gz8sLgsqKOZ7qPyrRFm7YmEM69nlkgo6Kamp1GNER
hLlyA0NFbXEIYNdPp2AkZZRe58nCdJtx38deeWG/j3kXjQMst4icL+HyfdDvJRn9NbHkYwZpPQ4o
PjrTamNKMq+jzhD9pl9c8MvpteceE1iJyYRv/K7sqceJ5O6J0m75IHgrwnBwl35R1khG23C90F89
4Q3PE3auw0T8ikKWA0H1Ae9ggvLKQDilGgG7xfp3lol4BVFZhNhaVjSdVhwwOfKq3UZbhTCGfymG
81ttxsSUPVzw2QRlza0gagbKKjP/nKB0JqObfPIeYVNDn4npfFglj+wqScufd8k1iWJTG3BWxjUb
RJ3yunZaiJOR7cZewqnP11iVnETA9fskAhV0Rt2U0FWBdGGRtb5cOTo17rZQun1yKLhaHpC1vKtT
2Ky08Ga/TWICy1PAEJl3Hnp2ZPxMQ7WBmuf9fwv5Kl8shAJuuT4epx17SMF1c1gA3LBPdfK8pdpO
Nff1p5/+q005HTYxVOoLxWGR5+Sax+TTb4TsFGICBv4d6Yv8kWusTDi3LbkuHu8lXIUChU1NKwl3
S98FVRUgS1Ex2ZyElm9ZNX9WDIrTBAFlCuknnC9jG1j5Dumz42tuJPnBPpiOCEyXE7SktD0tXzKk
VEHoysVvw/Q/7J0HyRrQH6xlRsExGwSjoh0uC0nxGUzpdfh14IJ6Lq/SsvHtCh6gJyynA0onHJrh
l46egv2sI3cvWlTKpdK0HZz7aJP9SPVtDPj0vJcXQ40p6LHp3r6mT8YT0Bxoh6k+8Zpjf/CMi+Oq
3FHiWEw8O3RCMIC2PvugflVS1txMGpIeLgyhh5jg1sYodLlh4P1V5Q9p4n7U+txVXSIzv+Gmy9I4
PT4Ko1IVk1vPCjrbyxlZ3RestjdH1XzignaanAT0XbHTvodH6umtd0eTPPHKPab965VRSfNokAVM
d+9mmeVCx8Ltd5AfrfwxiJlTpR0zX0UFpIKBQGqXBePrav4ghZUosOCjtq3xM30eDR/zhOmZ29mm
CH1dTgg9D9m4q3a98KLid/m1Crlm+EZgqdA9gNaKbe0gEUShWHfdTAKUkJeETHzpFIGXS8ZLyfFX
UDRnhELSa5LYF1FU+kS6wAiiYr8iIYi96Zl+8rxu2vQ2z0WtdTLuuTdgjUfWXFMrvd0qHUEA0uer
XpMhgZWHgRR7jFMSc0HWCNKSxk8sFFmKT6f9KuJNi0VvNpl2rcx65aiP9HlCnlk2MWHnuqCa2kVH
EMASmH/pcblp5psfjU29YwIqxstx3/WvIswnvvL10iOuVr7Y8P+RFS9S/7pfMB51TViMepn+QO/b
ItvMnVOcAPvx52SAnBmJfEiOXi/t+4BjThrlpZd+2+RtwbJnWHOsjObX2qvGKcE1bKVQuokIG4kV
6SQ/90m8xrIPKLGUac/wRDYXVFXK9kcmY/IPJAQdGhOkUdwiQziyaQm2hPRMThIjpU81mnIaydjs
dZf5pa7deoXYZ0+bV11LOZ439V5MnjQWUn6XRubpWHpoN9l3O7Ak6P0nlknDHI9tZC8JpXDe9oGh
2AvL0NCyJrz+aAjsTFHG0SM0tVK0sYjcNpvdJEJEA2QIZsmUtlIVlV+7IJ8F+Vl8bAYnOQWyMkQn
huErt0wUIJQVKlHb3ocHuWMkEYdpYQxtwyYQO8231g+9HMDvyKVjo3o4eY5OHcDWnNah1FS4+2JE
pRONxUwqJSVgeN/hYflbdgdMa4/m6EdJ4ku1Zo6eL2GtU4bKsjM+UOiAxZm4CyfmpGQ5GONhFxyt
GFUOhd73rt3ri04+GvfkjAXkn0SkCJyvy3OWcAsEnBB2M/UtBEJaWYa49jESqG+aADOFhQOv0iNK
ilYUSZs7m+8G5V+OZDTFuGpsLkxTbNHiKfcn0Xr5mc/PbGUR8Vs0irdBthAhvQjVx/mCTViAt3Lw
Dwia1gqBDEBjeVoXeEdZ8TS0Brjaq9lt49U5lTVRvcvrcEkqtSMHgizv+ERCa/l1rig8DxtzNl+t
p0Iw+9eRaEyu84YspVTQC6jLEO9orvauEIhLLILrcEKzAgF3CWtz9zPvPhoVhDVC2fDl6vCLCGYM
3clsEqNK0Iabtx23EAL1MtfeQOI+imdgA+ojPVSzh0s765l8u+wkDe2+Gj0IeIV72i8WAL0kt/3x
+OSDE8X+0LV9cHtTqq3FZ+/NkfFWiok4K7ily+CT1hsmiLO1O0q3v1fJoJdLP5UvWsUzzeGLzFah
po1k0TLeOskoUvJhjZsFRnYN/oHdZQyMjtLc+3ygjsov+csIXkBPkrbodkibyF3nn6ByxAiDF1nX
wtfXKJoW5gZZRy28M8aGgjHgXIPZU/+mo+rMB/Z42Pz+f9Lpphgf/XXPjHQyPSxDmI3By9ujNoxD
ZV4JvGWe0wJbqsVHBRWaIygHFdNtmEFFnqg4aDnDQ8H23u0/HVJAT7zQI/KQKeSxLEq4snF9js7n
KIkHLjEjnvExHKtzJ8KXO8/nnISyAtBLpmq01ZrEyzH98jeSnLPwh1mk2s29RmYmcptIF6FLSuDy
LK2p8iHeikgPRmeDr8ryZ6L884r32RjZpEGjP1BzoXN8lfWeyIzohzHQ8wMKwzv8tGbpNFQjJDeJ
P+w2NB407e/Ae4kppdmXftzcl6i2GYhR14GsvjZHq1cwbRrjhgMDIse+wRMbwhV75FL3cMqAgdRT
MdkcuoMVm79reVBJuXkgRN1L9qNp1PjIJL9MCvLdK3/BP4rrc3Sa8eBhiAYXRk35pDkog0NFOe58
y7xpPTdvHzuaR2t5bior3wAMpLnoX0VixNZEGKIn5vRF0KILJo9T9DtycDCFTAmhBGLMQLpy+iuK
FeyVZYkyqMPTBUnoaPiG39wG7XGBuqaPCLR/i5iCk68BL0Vkhcu5mAqojU86Y3Gx2tOtp5CnkMtz
yv5kBlISCcJcTofPdrRvNGHjltY/eu3fvAO2zIl7AnAzBFSbQeHbFUf/9wJNkZyhtrB7awLRpLMl
kryegqhV0s3TPTDqaHA0TKTQxCXlsyfSKJW+CRxPUjD9ZB3ncLS+w6r17F+oucbrcDnCI2UKqz2z
K96e3jLWEuVb9TbakdITeW6w4fCn+8+8misthnmLHaVofpqARrAmucOGSYozyOi76xRfcl6hmd1R
3xSEcL/AYPOH/Rb4AEhS/7ekZ5QOCiykKxFgUWSNCXOnbR0SaCWSMA22zitMcR+nLINpCgvpa/Os
tulbu0wWdMkX6OFUUOvW3kKhAf2ajGiiQrtlAgPhNueUNF9RtEcVAe7nJWlNc14XWvsaTOBoS9wG
eW5402KqjUMXoX9JPzIaq1T0bELdVs/pJuhUrxfdV8rzI4awdqY4e1jnHkl+B7K0kX+wf4cGrvfP
WfgoL9BE/sHaByt4o08QLDBQ40FdwQI9PPXQdOypfVkiBI4gxaRxLwOb2sKigJNQtQPpnzEx5Rnr
YNJtr5SGaKrkOfjgpYT83jrCuR5Fy67kjdSMg+EmQkOncJaVjKvKDp4KcG3AAvICwKeUbcKBo8O2
ylTaIGFJ4W3pnFuRKl0lGnk274DMriSZEnntNSORgOkF16hg51taWZnCwra5oQHFGBGJU8MRAksj
wi+oech7VNtMqRS9P3+SEnpTZGFSESPcfBvJWgBSnPMgij/0olRzybooTzISdzI4diGL04fl/BTT
4caCEYBgHfsxg+6b8T7l1XFlec5iGR+ILK24KavO2/bIIlRYXwu46Fx13ZQDPmGuRf5zH0IERt9x
HBxrh2V15z5WR1+ka07t6sRLNURoZQ7BP9fDICmSDUYGvhSwiFxr8l7+Nn9dLwTYvuvNY+MFhm7N
HgWNaK8skU5Ii8GFJkD/sNCh/NBmRsKX866OGb8YMZss7zyELfRBidQgWNnGb2gPTJNDOStp4Ost
NkaA39EFYepR/B51WRkHxoV3EKbQd3Kz39YhekD++XlYs/yxFN5quwqmjPHR5rTpYN1QomttX5sI
LgBhGYBh+ctuw5KJf5Xr4gZnT6FrYK3ruKnA4SSBTqhNEyODPWZDsNTEWHBufsjW6rMiLSQDSZ8w
y1FQsRnAHAbo3QjptzlwyqFT0u53F7cOJkRMmU6AyBGdtW6ojIEIeM7eI8Kf11/wS9TWFFz66p1f
KZqS+5yVjV8K1E6Q2E0P3narE+5Pf31tPy2K/WI/PqnfoHc3LbJMB7sz77Myc3z8USz1diRE+hWQ
ZoqJMOA2ivTkZm2G/tUqRFbMo5fTy5BBaJ2tdW+M5JTXBx7vV26jpDWqee4NMWhs0CDJvzErz4V/
5Y6askhoT04uKHFapb47OE+UnKfhZDunenU/fiGU2F9vqnJiU9jpIFYEMHQTPPTjANhAfTjq4VAl
H9RmcEfPzRsTKBKbWJ5UiaZaOVjDbm7Zj0pzcAL31axrFD1U6T9odu8zyeLuoqP75ZP4JN56OFRh
sW2JtsEiUGxsfm6a34oF2WUWHn9BQchp2Z2FNs9zj1XtjiDod0xJg4zdaXGsFdPazKEjYW+JBtyT
ATgpMGcFUvAXu3KjVB725q1UKnDU3N7vC5g0u3B5B+DwamQYylUia5OfqK/66PyD0etKniAhgLH+
3T3E0xSnDGXUt1qtctI5LuaOP8fHazyma6Hbc9AuSw6mqrcjtdm/GUvllCy2x1llqLKmc/juso7y
U7blQIYgPrX0pr7MiAjjUPmuO+m1a9ksuy6Fwp7KEycamcw/OFBJZAoZt+xuG6SfxIKwR0mFOPa4
dbt/DhaicVsOhOLa2Nst22YWK6VxBjfjYV2dtraEg8Gky2cp+BaiGjzmgYb6GozwTXEyJCEVjnmG
atctgQ5WA4CmeIj2nFPU/bH4lPVhAMmswA/LbOToWcZssAN3mSFz9Juv2ffLxpBqksYLEfyXeP0h
4NydbQRwlrD6Z0C+7FJr90a1AS2prVt/NCJdVp6yxMXxRyMWC0O55FkkYCcAWvbJ60++qrVK/gig
+0lea4e6Q6Aokp4SPs13C+KvtKnIAETArDzkCoNmTrlSPVJPXn3STdGefQp+MBUlv/9zm1ADO3vW
njpicuI/DcTNrH/t8hj7BczsNiyHdHLEjlZcPkuUx7g+RxjHDbmmqV2YdrtaSL6xWdO+Addh9SZo
ZiuYG93a59m7MbPJ0ZkRP5DbemuB6b+/UdeYzXg38fDYQKLWZPutgYCCtY+M2g6A0M/qH10W9As2
Z/DaBZG7z8IgbWY80dUHw82HF49xQO3PM8akFRLLpNDTfXnDUJn+jd2uSf+DXTFyulQDclKGPGgl
8+3cN9sl8jYhEY7CQ/MehWj6oyRCcSVdPxR7R0giGiaJat8R1cTGktE3mAULSfcY/8iy6lS+KdMN
qrsEOsY6fc6/AxTlnxwuIwRfZsKIOYKkZrLuCPe7Z3IRshGgJWPTmBNc0bQFqKKBHx6BXQ5T7//w
srb8W08a+9tY+IrVG7XsWLECEKR/3OYrYyEn+x9lGJjLJsMmBBgHrRDjGhq51Ikw724bt8nnqei3
4kqSW/RIkPhBhGhxY2PFkv7R23Guf15H0FxkfPH1/r6s5sqwuiP4HqDY73yXoOshbRMi8fbWSlST
hIBFx4N0Y6vPx5/SEJCHeeAmTWDTX187cUnIXrR2f1+hHrd4qv2bwRsMNmNw/exj/ZGTAwK49xJ4
5OHJ0VQ+C8QGllDRsPdbe/8NNpqH/yuUN1I7rI12ETXhH3pAPWshdDX4jU+ucglODlsSmtURTE+s
69Un0STDl+IvkkwQTXpG0ZbxyqEyQJl36cYppLT2oRJ7RCY6Pcmx2Zuf/vp2C52Ykf99BMMCRPnJ
8crDfunDGAMCvOf9JqHFvg4y0NqetlLd0TdA+8qDtX/HvW8VArPnbNHJQueWTUXChxUKYcrIHlT9
0tj4AGnNRq4c53zXCZ189nCNsVkEiNz6rTIbmpVT/E4BpF9FhBnsqKVxFweTZVzDhPOwWRhToYlG
3B42CVA5vffJeRsp9ru3Mj1CYVDUuvFObuilgxBWKfEfPKsn69TBvQI/yqMQWvNSI8Spsby+1N0I
k5C2Dh80MuE85fabk63+ZKYF+aTNNYc+pNJVg0WZeg3zQTdfH6Su1hHrAmF+BlkqUNMBb+YzgPX6
SV4kgomjyEeUP3Ho+PeB9AtXFZESKRrdWY2+ZkwJbXkVcfRwOPMYHD+Z0u17lUkJttiL9A6plwFr
H//XhSK7zDbiv5ZhhBcbl10Q8y6tN5dLJ0oorZ4dYWfmjLebRusf2nobjNFh8R9opIhCs6wQlsNs
6hE4wZRhIC/n28IaD/08S8aoV+xa6prhspXv19BpZ+Dy+FWS9nWCVS42d2qjzWt5SE612dJJ5H/j
59fmhDRr4j80SMI21rNsY71GufAno8x0kOW6DLqURrQv04heOBG/RnMzhorpgH0w6ciPx5VNhJN5
f8aOoa1jS8HP/aMFY5dWi01R8Lga5bKwLRG6UD+xQp6EfEYX0Bc0U3qOSQIGwLP1hVKp3xXm5fbf
EHfa0l/Wjt/Tc7A7QF7iIyCs81TDvfZ5vPYe5xuVYBbILjo6eJnK92jvUOpOLtiD1DK1K2d/JBzG
RUw8pQM2Mnl0Yj2BBawprZXs5qow3I7wm+dUQo3oEJYEcrHeobWM5qFnAxQP9huizDO8g/PFX9cc
+n85+7xLWAF9g93oIs+pHtxbzOqf21jKA11SyUGpznrLdl6RO3RaPzJdE4phVYEvVO/KNvwRA/Hl
U/XP/jrRv7v2zQJrbohX9VEDBmLo6HHBOZPniOrsjD6mNhE7WXJhyi2C2o2GOgd/54+TRDBuEYrH
tr4Vz0gre/43nUlLxtqk1CjSvtNsqyyFyMpqP+5SLUNLNYfLHZ194QYdGu2CnHvcbZL826U2rAql
hmJPMGtL3EdNnvA3UhpbTVoWjWZ3qou8Ion26A6otIBZlc3Mt041PDdSXRGZ3AnCOgUgEXYF3tNf
BZiUAEDi1lOTqxONtoilyRfqQvShRTgMPZGAQXCOQQh1H7cF2xuwyuwKwsjEmYjCd09XQU2y3GJW
pibePcU+iOg8hiM1tE40wiCvDVSeX94w6U+xXtqal4paIEYklXKXR8mKhFb4bfeRRuRvilISGOtL
gUhQNmTsibjNxdRG8JTZ5Ct4+gJ2uCHZxeDmUg79T6seTrqFzWjWTkhKyhvvLkRZkC7N0769cvmV
Oc7zGLuWLt+/ekFZkl3wuKOpKKUxdlzjyv210YMvKV1Cq4rfxuqbdDj/ovdX7qfPlxwDHTrDKlLs
540WcWXE/+Geh/dPVwaPZVhbcYo+ftgk+hj3XeWYqiL/ObBaPWrdD95EKPsQ9RW5jZsEhDirwBem
8kasDhCQwdC30LtAmzJvu9VIy9/Go5ix7MWODjL35RtQAK9LmuNBzTc42rmnEyiXAbQeR3CfGXyS
aR90emsuTgr82bU8zMNKGoevkTLqRnwhxxYUOXHKNJhr7A+6L5SvGd55kt9e4NcBg9o3ud9iuDI4
WRJssa2tTSXWFvPwYWctH3gOoZi1lMq1QhNEJt967W7O4encYuGUTjf6tPzh5uKVIAEKqkzcF73R
XuKcfSxlZMB8pFMjRjFVo5xiIfc07TJCZUwoWGrmjMNz/bnbQM3xHqJ6xIzlW3d34UqPlupCewb3
tDcIBvwDAQ+QjhOvbnk2qepabu0paSlB6A36uXAHSpQx62kjCHs4/7p9z4CrQvowJXXqOq1no4LI
Leym3/Ad39cpYEAPmcBDyBNV2ylxFuCEMtBIrDbd9trmAm8Cd1Yd65dZJdj+pJrg+inyMxiO/nqd
hGeZh1FcxzyFnNJ1uFhB1H5jNvES5ptafc/K7ItaIHjG2Q3Hw2Sfs9tdc1aTo8wqj7p5qi0ooAu8
dE37+v41wjH7a+UDA/IsgTsgWPMulpuSwsBqA3ra+iQ1IsM4c1Pj2b3wD/0ieoi+8dPEVs2Mhy+a
Onkb/G8snD4qIQhR6Ri/gDxb55nS44KdIUHRuPpV+hjaAd9XjeOgfcfnktxyiGsOtxD06yLNj3uN
BDwhKws851LqfzZTs7rnPHFFCpqvogySKQRoYhc/6G9zWEeAQBw9zgxtOTRQ3z9yW4b/WzqP/HCe
YezOjFu4ozRvoURmAPWu8JrhDSy0VrKK01DxZ5fERuQ3jV5EMPzQmZWYry5BgW+9U/ydg6j9kaLT
r3ysSlvJVUF5L7I4vq6ZsXSXNnqkWvlIeH4/1/dZl7yXXUPLqsgSt+Y+fEp9EuHa9SQUcaCRIEOi
5yrABksjUi1aORq8TdP6c5DVHlWkpYskuAiQfJgpfyJ7KsR/UEKae4KuwRPBFuZRKUOLaTTroLW7
Frha4RBCyYe8Yc8PDZVsUQSlUNKHoQEUrLkkn7++jM8c71luZt95vElRh1ToXt9vR8dStKy/i5uc
O1P84ZIa4bEXmDFxMlsEOyAdxMj8p55kVJBYJIIHoKDlS8o7c/Yp1EEhj10p0VycZAQi91YN2geH
opB/6Y/LyPf8ooZ+OU7FeISIGeQwogxp9sr97v1nirmMWF2sWA4sxi+zLeGPplnfl2rBXy4D9DPr
zy4qgDbI1hRq3oAoROqPZu2IEVBPys7JM75DXcVqhAHX+uiGFAj46bgX5MUa90pcY9SDmNlDJfdD
09QqW83zsY6CciTw/Ip/VwA1S0xpNIXXw+/J0zNJafuorJSbcSP7wI7kVSRPZHr1mhP5lxYRIYJf
k9ZCUFZqd0Xk1BwiY9HllV3S42D62eCmnvW1d27nRZI7Ls7NEEfJxi4DeeUg17/0J7G14htsXHtu
GDBt7ykujxTxQ8cXGLfz1Oi9vVo1jad4tmqyppbqh770aBjavZv1ZbZpym6z57AUCsC4kYAeITeu
//3rGOW+NCG9fY1gzTta6MAz/Ye1uLR3M3V+zrbggX88lC0eCaKT9t0PhehcrDbpoF6+11hFWYef
h3+Ka+iJkeRGXHkUwvBMevsytw3y6RpmsBaKfNVuUtqWE7w4BIfwa16757kR6W+Cu9RRE677N1qd
KIEMqn3Ebw9OdRMPSE7Dc6zJG+mRPYAfyEt2QC6SiFGaL/m08jKou4wgh7wavYyEclIip86Uz/jv
wSzqdGxPmzIee5wbIvoMhEuM798CbUiHD4/HAgXwXbOt6KdAoEWMYng/jls0kC698nZz2GmiEEOt
QKnkQtX667+FbBPkmy+YQjKFacpZdY9qQ50iz8xiz7qyL0Hk7kDZp9nZ0PAzvsh4KwYOWHauPksX
68euoi6onPtjnyUV4zwvOSkA3yLLenX40CLhIn6KqeLCMqzGeE1DXnzNFuHeO+0VC1TscWJD5ROH
SImfmymf7o40dwSl5NllL4ssVFxYkcKAv5ahLqxTAA6GcIqn6wSnzm5qIAK+QHA5FDRRZOpaQ8qn
7d2ZGEjZrDSTBgZDMehpZLL9FRa9GnRjYBkWY7YPY2GV2oCbKnPbs/2I/U7VDcNEF+Thn+4cuNAG
CpdzhOqWxqbhaRxM4jQX5tz2jJSOUFRPJtsXnWjrlVG4pcpkILcrzLX09oqGI6fEQc46GxW3pmvT
FMz1BkWtPHuuvpW89Z0EvsjR60F0fzRvz+zEwoURgYNLV0o5KJb6DGfbtiHZKTR63TxvIymUGHyJ
xLK/42b6RUkQUQ0nlAdrZROxmXH00bGWb0OQz97gs45kheRuici2Q0/Q4BUYw1T8VLDFUv3wfH6X
rCPAToCDMDEfnpGPbln4ikGs6bkTYjbAP6mO/jhJ/RfYTA8hyEQtkEs5V6ctU75QQd0H5JG+vfZD
pjkFfV1WpnOTen4SYGQiymuD1gUckwmSBOyXU99DqJDY22Z4H5/NBXJMyCekZHJYQNOkQhCDtYV+
vRdr8354sTNNZ6TFg1rvpSDiAz6aWECta9vRCMEPDib0tLEzg7ATFZfPQ/on7nY+fF9KpC4V3lbH
1vdS5rOJMNHZYC+npqu3Hwx/Qjm9H+fIn4LtcBdKAogtr5qnos+KoDqbFB8nOR/e8485J0PSXDpI
vrsI75ZXu8yQaZvwiMIDj383smehsFEvoScjmH9b2l054Qf6e2F61/widALS+712KBt5is9KiP1C
mBsdloCtu5QHedBzw1xYYxTd/figTlY1SSzrVgmYQKYW1cWmFlcG7JFSu4YRSkxNpcOiYsZYCydR
t3FE099nKKZqiOCBoZAuAwgTiJNhJDFnpB0G+lbkroQLwCwpQH6TTcDzZm6dH/y9A7g1Ql3Tte78
lgocH957OqCTX2O14eceefWBzHA2QXW5jpYNOzwqO4I0aKfapw///AAr2KJNu0Z98jOytkgOUKi6
pvGguZcbi1ogRDnH+2jVs8OjknKYJMh6tNknZQ/vO1MTiTXAs7Updmkj5jWQHtUZ1P5vshyKyYT9
uwA+TswchLP9LIsRnNI+PmiBlSJkKBkb0UgHzxVD7ixaMb4mHdq94J0AptClTjzf7XEaw6JfWoWt
XPFlAWMyGEeqLnlKrnhlD2lwVWwVtSiOXikDvmps7LN3dxW5IpWfNUonsbL8J5jgUDJsj4SGQkW1
SNbuQXBY8mLqaSDVehlHtSM1V9lhNLrFQsgwXaF26i7+Oe7daVGSE+32VJU5KlybwfvqMMX50VAp
yIQBvCth90yvk8tMZ0v1/ub2KqX7A1VQzMU+Hsbl476ck8qdSIgCsUwmRG/IuTy83fx1UEw0RXU1
Ja4GD4JpF0IupMrkMLz9nyjXlv532Gje7+06ISpkss9IU4/Ld6JeOfI1zStdHAnJKh4FQSONJpxz
Bee7lf7q3ym6p+6Yhta7QkJl0PqGS6xzkzzkkVL6yAKlhbmMPiVk4tK7ztugxpdkJyt9ataksq3X
0fKThic2zEu1hZz3d1JvI/Dx8XGEvf9NVm8q9cAyxKE8d+FwVyxro7BmQD6xp4iJCdbOvmYkEHjU
+TDQPDFO1mulxrAI5EhehLgMFlNYu3zwnWHPSOxtzN2pJNcDYc7KaBWXuys3fAB6SNheWOghJL8G
4w4ZB3EtXJvPCediaLsZ3uySDniXs4yjiRsFWpUCWXpZCI0gow0CfQTkAaX1FMG8Wl7kBTQZz7Oo
obPHOewDA52v1Twr8ymhXWqzpnNguUGqqsTroTdjEI2gcEqnXMBr0kbAxqVnWYr0HTHqinmQiBuD
09+Q0P0eJn9LkgAw3UvdgwKA3VFVLmKfbVywfWQ60Zx61T9no/7cAbJpLei+L3+qw0OAhvhbbhs2
Y6NKoEmkN8rENW3xoGr2Xmp5VfWrGGTg4d5g9QlRHVziDO00nyielklUlv/IKAllIjLvqyLCHx31
0q10A1Ye64ULo7YbaCI4w7kA2p4EDYg1ChJ2oZPnuhf08ddq1ppFQad7FHNF06jDa/cNfhat4crm
Mlwim3Ondpm6epug1WBSzMvYxYhi+CFNk7YoNPUW09amLeDSncHssdv/5zxDT/tOXpQa8tjIKJMH
GCVbBF1HfzTHPfVTXjPBZ3o78tMrBr1pAxwwfuN4STtkkar9InCpz8GMKlopa37W+WUYOBgT9vZ9
+TAFzaYJtIn6PCMppdhu+0cb15fl1FeWqWvJ8kVeeWNI/1IBnBdVMXVtRj7tIco7QxMHBsebcfGA
JtVpriihddG54EKB6uLxySWER5sm+ft997LTiwkBa3gypCJNlxdZWbBoUSdoSEQoqlKMqNjhQ3P7
WdrfGLjOA+68zPBHCKNWiiKWiDdj/sMdTP1a2ol1fhOB8rD1lLHxnSWUx5tGnKMxC2NVjWH+l/Un
XP4zYeftEy8YzpOOiK/o6e87LQEog6qQZ6k2wJuLZYhYd4dL9nNNvvrWXiRj9s+dVwZk3t/LHPpg
iKCCyNSkGdiyrikdJ4yOkSSaYoVhTo/tMZ8RHbX8C9nigB906TFuzrbT6CeSZyOJ6DnUfuCE2czv
be/mUUWXwlhlSA8t0FiyYZG9k+V7vl1VwWK2e5bcDkyPYDIc+jeabN9dZ8c/kvrmKTr68qm05Nxl
FjkwieXmf/yOfspKTQO0Zzs1xMejiEHqBoHtX+0kDCj7N2oRmwvxVk2bx2sDyOii/bGjQVF1R4Gx
ANaFnTyo9SmzxKAamzGLl4kJFaWAnSZ0+sTFUiO+uIgFTpQR2KXPveRhCPkP61ZFXD1O/GwJYmde
+n5y2KmLNAjITyiK4LUlGjbFgSP4K7rJ5L66XFAHLPkpp0ezW1GFoKHccGh6KC3JSH66kFDiHExI
sS/HlNsflW+VINSM+ueb24fD3Ej3MPmxgsN7CVpYSRKXstgT4XUTOUDG0X1Zawx9bUiX362XdQGF
8vhw/i50vaItUJhD3rU6Owj38ulbAgdv1AEsGWL984HTSATZkFlqG9vMFiO9pQhOQMNdmeY5B/T5
mzzqczsbmr5lhWF7NyfYziCdJ8nFEvQNos2snfjFfX8s81num7zuFpDF05c9aCo81OepMC6U2+bF
E4VlaQuoeFnFjko0iPBks8mNrgiNzlMJ/xlGEn2IazHi62RNyqWCL9SsjLSn3MaYS1VFVdhuBZ07
HWGxp/toD+QUWrIjUBAg/fNvbJTZpGRcLEkXdYEeOwIvbgqkT9gUc244153JJdZOkyP8rtBDGBEX
j3p4+QuCHRZwcV/Nt+bMNKcJFYr3c6wlhwyoEVzVUvDq6bphS+ul3P+o57P63DXf9nliQiusiqs/
A7obTenyABVwnbK9s1iT6tBkPFLJw2q6AwHCd2ht9tCdIsWu2NzepDtduFoCRf3exYSGwzRLvddZ
sqxk9AbeC7rd/Q4qwKo3Baf4o07ACq4p+Um7S1QUNlRYzWw1JSUfgB+dpcNRPHCmR/cNV580Y/3o
C3Lk/BDXyy2vnFLFj9zZ9/u5TXbeEEFM12oWFAJFre3DYt7+9Q1jKRawAyGETThCqGlq/7xBZR2w
u+2nU9SNJMaqLDjf0ieRGWstCgfsUWbStoTUuLIjVR705DoMjsiKeFJZFILwzDOvgEPUnA53f1Vd
UiMWuwxCI/HBlQVXRYarH4M0T9R/f/IQ+NSA4zbPF/kwXE4qedzKOIQPSgCjGUUC1Hh+21/VAXvy
bo4sXZL/1JOkI8N/gkWLrJ2O6P1v4EY3HckTV+xMtOOOdCMeza1LHYX9iXXEcyEkIOAIvZuYj/JT
FWfYAuBb5iv4jrlA9yXCYE1/aAsUuzzZOUh/UEFRlPvJvP5Nl1vQE5lR5ja6AwgzObzHJyrZFEuQ
msjEONJnJ6AcTeLCbaN9GRbZw4WtPS/Rk2kuv6eTJIrA/zv9MI0rBCpZcnpVilqkbzlltDlImjFE
M66UGanX6gM/9RH5D0+XR+p8ElfACRXg6wpnWg/ROBA8ObxM2WlKe1JDA3hrxnW38kIHBRyIWNk+
0ysW5rN2iVTM7Ekx17ep2Nw+SmPP7iap7T2vpmtcYwmkTPKnmx00op8H2p2pRuSeM4xPFqCSuBEG
Fcn14sFR2H1Afo2rvHG8/D18f0kD2KSSaxGgT71TZjhBaDEcVUs2t8osK6RLDm+WS0IHn8XKwgXh
00dGm8Ec7v13UxQr3Q9R16Tfw8yiLEGNr4KPmw5DnAI7n7OFpRTFKUS58CTwalxyMRrgAnEUiDSw
xfevqggUD0po4/p5qXKNwV73j3VhZsS3uZytQOB3l01masf8F9wBUQ9sedSUYMCB2wdHviTyoR+4
urrGGaggbt/SCsfaUCB2psFtpu8yYCS/AF+p+X4vPYt/EpjVA9jkaTUUkzG6l9HSgc1ItRGYE3jx
SrIm+92OTHXrZ4paX7R0DT1+7Kw1HrBzwhwvExZUqwwCMZmqKYuDQwm28xtV4gfLQDcA5XOEDNDA
iuWryjSrgGncQMvQ/p970WmSoUJp0NIHdV7eKD1PW2YUqoNC8MbeADLSUt3EjsI2TfXsl5iNvF+W
C7jhszKIW0JMkjL6VNC7yeGkm/gtjuNcPsUDmy9fjvIh26IcVOm9wrjY3bHC40vL/vv6+Jpssdoy
NA8FnEk1Kh3POinRqkBK6sfLc2v7SEvZN2r4oFI9HJ4V6KGwm0XlF08EAWGQB/ctQhRZBDZrRhuH
bd4qfTEwvS55C3xQn0i5l3xCmOl0HZ7CU9sYQZgTLwyVlOl77vgL9yPDGO7jiK3pmBeFH0I80EkV
tY967Ayx/xnuL5rHai+SUmzp/Bat7u/sEjryMHslw+7wSOpB+57zqZVLlt6HSrQx7iQLakW9jqcz
YkrHe9tz7S4YGa2sdezrykN4SiE+mToWKpH6MsxxAxESOwCMISMx5tbzf3SKTXyYNfI0zOV0pKrH
n1CVZWa+6X/NE+OwtKcn10TshAbNCynngVTHk2oe18A9Xw8u07puLBV2tqmpBxbdHCi8VYnHshgO
IPjzWy+FkmnLR7F+3aH4DRtJM+z1GezF2/CcZpnDlMEMMHkotzD0q+2hn7sTRhzrCb2Cxjwufxq/
qMPS7AUgos7bse9aadd+bAptZ7aWSMU8zomF15Tv+YPjNTJZehwDIvkqWFgPMuV6zyv5kt/K0p2D
Ofviuztl+PZeadaYQz/BRYB5fpkW6kfSanVCJc+2gZ4PwXF49zv9Cp8O8RQPTJAJMKEKTb+p4pAj
v+nf2RoPwca3tqzRfgCuu4vFzkRq+a6wyUWwXNT7TklGY7oRjT68pgGR+9rjv6izHdwpG5SP8aKS
TNWE7ULnvdMWFaNeQe3+FxwejA2OmM4oigr0y1ppOxUTdAhDItsk6OlTDcNI2Jr5zLLIMdRjYwvk
Kk+JXZxl70g82srAv+mVGw47+OcKxKHH9a8ki2ivRdG0QVcfqpm4mZ7XXTqNNE7ro+cb7EYBweKS
x1vKKLjItrpyUGaVDhg7XNoUB/rsg7iCSoJ0+/MyZVxM3ICKwAu/bWacr6ZTd4z8Ds6g1VhPPZql
y8n3o/KE8PHnFN0hloDHl4mMy3smA3B5U0cg4DL9f7k1VaGqlNfS1dl3eJWez6g2VzP+pUyo2obW
hesR/tGyAq1xuhtlWdGxVWQmuQbpUWFBPvTwK4rImID0L/sKFW55OneH4ezjh2nknNftIV0Bzj5X
EJ/lgC1ZiVyoD5WHbEPypZ/8nuUXI6HNwBGitczVhh4c9H7ZeaSvVj3YeZTIMROsqmEi3Nc2Ly/7
omDQWcgLN+5+Nrd9z8Ep1sWA1DGP+vLabauxUQoWj2q7ssLU8z8yf4iEoJ8cHnnV4dGVoZbYf/Dr
2/jHUleVCqcjg/h5/qmWfmNDPZKNLUwcZVLusBJXm7Wr0Ff/Ych8x9Pxzw+GnkJ4utkq0vS+b6I8
nN/9EAYy4SFaCoytx5tztoVwpBf93G4IomQlny1PqakcZSRQFdrI+TnVhW1p/Pyojf6nEW3wi/68
GlmsYg4f/+lUIIJduyNOdxoJ2FqqNwNtaZcbAWxUbjMP0ve4+gbpbTYu244ZNwOLmymmJL4IUFXS
ZTeTWZQYyASF1R2v58j7k6RAcM5egmxfO6WiNHv1eH1XFInByL/ySXPYMfrtbw63B378EZPCWwP4
R0tvY91nHRzCmgdiiNOidcr1u/0lNhSG4KF7cytScRkYWAYFowwDVN7pk0X0wQEjkUhhvG8CyMm0
9uvBgDwwCkARwdcwjy5OwE6xWEy+uD0O5puYrmrGVomXaBnwwI7hzkykZT1/mOlMcWlos95g8tHj
4M61cIJ6qcup5qGzcFTpRSKrE6uhbhhQ1fyQNGWRgzgtSt1IzjaMtHrbgY/TCoh5S/6/2NbeDvY6
S9ftZupJ0bVbRsanzaJqxOn2u52OX6yw+B65Mfe5e7/+/votsqS76fHKOH8Pe9iLomJinxkA0AXq
5GP6f0qMMB7Nwyt4a6bNdboGtKccF5Sz0w/3qZSVS9f1Zo1+y2IbrsCPPiUDBRoKF9aH65/27UWI
PySMKSHC9CUpJ1R3WUUFdohJVCXskcioIFb05gZKnOGv0QFJxuXLYewB+13yD5tIOD2k+/Xtt9ld
6zrlEL7p1KYqi/VO3DLkpDVLRhgQAN1O7MbAqcouXq0cQa5m9pTwAk/3Kzfvw9rSRo03Rjky+Azp
9nj/YevAgW6pCRroRh1gz/0Lh7LM2k4pC/RTUmIMJcYPAROzKa+ZE6Y+xrt3sYWnGr4emfmUKXxe
eE04WRfojTGasoH1ngFBwkuegZ/XxNU46ssv7+Zb2q925W7/+8HlGmyPVvePQTC+ZSbKYXgW6X94
FfuOwJ5McZYjadLRTGE0wCOvxvexHwGuh905dMKfGl36eNy0h+sYc91vcH1T8Srn4MSn3+ii36EF
0O5mFDjCexFfHc8BgQJHMarv2ra/Jj+DdoVJaVFEj9TljCfLjWdMES8gpL/CYkEyOWAtMEiGbn5t
9UcT+1ZfNY/AJvpnj19expuI9S6UcAYttRagAdOJ5e+eJRVwukSTypSuo7t7MFC6xR9bjOfj86OX
aZUivJkFo5wxspjwqmNYVSlwiqs+n/aPVTV23sh3jxaQ/9r6PEskk1bWhi3wpcBHdh3yGUNiBgJU
9BfyjmUTxTWAb+zlQ6EdJoPWWWxK+uAArMW6P2gTu5fYKOe2g8YJUpyw8+Z0jyGF20a8Wj07ZP8E
FkMie/EjG8giNzLfqJILc0aQPohbd9cFi4ynSvB8nYdqIgTQCmyWSAmONWMXGXcWSy2xLyFbyZnM
wk21GDmse96FtTeoN6QkTHmOlvt0lVu7pnDv08XUnLuPyy7IHFIl2hoi5AAC3lWwxSNG1lmDDayN
hHffBDQOQmXSmJKsagTMoEqcV700PvcOWrCY9NdykwNCnc+/07CqypEsUmx9moSJg+8Moe4T7Lzd
GvZWQ/F2zFxBHUJw+FCKNr4dQy4nk/WSszqQySmaUEXK4cbnmrVW5QYy6Q6gvMSCiik4A7FLOpsk
TeQXIrOLQyL734x2/eOV9lyUTSyQ7jDIdKkT0db3E+e7G0FW0P4eff01zB8EHSuSZKmo3/MJ9Tt/
aqOI/suqDUFdWurXf4toHPqg2IsE7Zpf0/sQ6tuoNduZU8L++5RHc1ivEThIO0P2zVNqA3w+dymW
C5cRvbQ6tPoSkVMT/LAvT6M+F7xqiR5NavoS2rwSuITynugppCzjhoNhVdC6+rve12ZhhdnBPRjp
jKjFziw/Vij8+n/NLXOQL8djsv+cNKCqkDr/R48cixKQ1sVf+a8Lr/4KwRjGjx+N+HZJcxOKppXO
qjEtW4R1ZGrcLY7oGrbnlTf0PEI3ITqCZq9diM+OLrByYbsuYhExsf5KjbvmJ1JFmeZbIYD7FcyH
v88JQHYZogXmRMbv6Pbv03dvDMsJVJh8Z9WNsWQbtHuISAfkrm5IHWHPty4rRZul8ToYFQD29jX+
jUGX8wCD9bH6HH/aheN8WGhHTGah/wXXzagFzCNuAGiY46XwNVRVrgFF2ACIMZCuxiN34QgJFgso
aroZcq/pM+seA9UWxSu5B2TTcVLbeewMWgZHfCRSYEgZJEScuylOPOECwbMbG15XmcbsJAFE3RTa
d/HlfMdhm0XfiST1Uq4UZj28h5HMxaLDwVBr43ORKnnphwLWCKK6X742uue2HhmV/C6v+9mYruK4
qwlqdhAJQDYvWr1xSBxzWA9NXy5Pnlrp4kLoy1P8Oct2FrpqPJvcQN3aeB1J4Ka1JzWBAWr+JJ3e
HeptWl/+cC7y5du+mzLhqcUFUTPcHDZr7+F7BLWjES2FkD5M6WFdAJfWMdmnT1Trw2syZHR8O8M1
RbzYA1D6Kjs/jJz89FFRGgwbdXcvgzrgbgrid6z/A6iBW6E2X3lUpbcTSP/dqzAcN/r6z5+XQrKE
+WkOYvJSNahhniXwYK6IBk+UAgbPQul8xVWbjdd0PWZBiYqwykYsukruwFu7i8b7nH1NP1+QomZE
w3K6MsH6KTdsdOTVfsUEbMug5yWes3wwKen/g40KkK9sXKtQqqabxGsWURA54ebzr21Pt9NkXzVN
nLJGeFsjcZE8zVGkmXOL/wkg1awDQrG3cQZgsEZlP8y44XoI+sJNEKYDKgE7OFA9Q5BfxEbdPckz
fa3tSy6Pth+IKNkvqAYlA0Qf4oT1AiXcrtHBd1rIjFsrXNAEfs8KbvyiWrPCrniUGVnMx09QiZF1
jTuSCUUWb7en4eVkJkgz5fWHczULYeDQ2E9SrzLgFgGaYgB4MPtczcdzNPltduqb1tlkYdlGR5Zo
DJ7oSk0wFiX7pGL6F6BQJ7DgibxNswalH5LO/RPJbNoLYnoCgE5/7muqN4Zne6ReZMKybR5rsNfm
igEkX3KJAlRHhjRg7EXrlHpaVCE2JQRFZCj3pwRfvVH22K+GLfzBgZcFcvbgb2yT6GdXECQVCDqp
zrBazvKF61PDJ2ehU8wxNKHuGLtvjrLT4/QxGz4tkOxOfsK6gGpX8YGa4ISEy3wWUlVhoYK92B3b
K+0DXyyfp/R5cdtBgLxveod+17ip8y5Otw6dOExh7xTlzvGXFU+0I1giVEOJKxYqvEyo+sdhJwGu
g16tCadKE2KlUMZQhue5Lxl2cg3RQEG30CVNYQHNBdBDGRoaRWDUBj3P4Sl11IYUFlzNEmdPtGeg
hspL+adl5nt+qHyrD+jza8Z886meXj6GGMyqiCT6hsaGgpA05hSelwxJdh9ScuQlHs8BDo8XRHNQ
KV4XuvdjPURQwsVmY8QBFix6VoB7mPurkIQiDitfvLKGcBY+r2jIVPZpWydn7NCjUoG5u07Ib1/0
PllNrRqIH1s6bXVG69CV+VE7fskHP66i1RgWTgrQDNJbTw2KlY5GhCg6YaeS20hgm/C5B10PFG06
4+YPNcxVfvr3FlNr8y+wce5Q7GNOWKHCTa2J+KsLpvQbsY3B5CVGdpf7536RBv7rhtOZCcCAfpdp
+uGabxtcHbhckVfqCh2RuEEnYmp7ZCT9YYKGiX5j+8z/z5L5YsprFl9BxWmfPDZZe0r3mLWdx80y
/n6KJKx49mCwdcHzk1KU3J4embTuAvWSCiQ6jBxLwfMVHY3VJA0EMrXCrOal8uKAiuP+V2HE83dM
QxGpgAucAsl+UXFPwGTOORKwjJHvVI5LzfoHvJvEMw8MA1rQ2kgdMh9IK7FuYu9jvsGguJ5d/lA1
jiFzxGWX4j7QqR0P3cqzVubDpoAD/U5azElZSkotIGbOmraGQU1EMiOsJSbiDIFF2ahokSYPcYlG
KeJJWVt7mdksL7wFBrGtm1tHY3VvbDJAMz0JsRHESea5bkd1ddR1fLbHLmMCmNq7bbkduSsSElSp
VEUgE1sTqbrdM6t/HAbxrfVOLShmHNPjwhaX895opRlCc0LJbVa6bSweC9J6yHvG5sGzt7jbhup9
C45t1Xr2FDj3deYbg7+262g1vaQ6HGXZPC78Ed0YTaGRcsBmEZuiyadaH+lcbhHf/9c57R45KlpL
BK9F/9qfEei96rYO4/aqG9pZwYLxLxONLsqDYfbhfy17EDa/763qCgJh3dZvh8c3XmGZA0yA+DYT
9DtyBPFDTWvcNBJUumpzNN32UCYFnjdEgNvde7VKOpSV5sjU6YTSQfRgUVhhWPi2ye2NhuK4q97H
ZRX6dv86wy9CJC6lcK5Myn8NrXDX2sadjWgdN/lcmUCsyuPmtsaEjm0cIiob/PfszlnjBlzkeDNS
y5ti8Uqkdg6ZCj/AUJ4g5YtaUx/mPEK61B0bYeF+DI/osaKiDiGLTYcBf9jZL2tQuLDsuQl5pWau
11XrSc6E+NSiC5P2GTqmS9bNQCvQllgjSeGLRXdjmoRhbHk65NbyJVk260lg9u+ZJq6q98a+Glej
R91k2YDqG/7zNCZ1nM7DmbRwANrzA9CY98KVc+aFQVlKFwKP0EUKkE231gTJcfKJvyaUTRC0oO7F
h0IZDHND344V2dJdRpyloKdnaV5QmRdbqzC5phV6cpnxCTERrswBE+AoTOfcS/Zp9k4hkYIWD3bO
0vCMc+ujSZMyjAyujbH9uWFMlAAFVb2aTd124nqtxf5G+zhN4/oOs+kRJv9S/WObTPR/0Rf6iy1i
Q2u2vv9HcCZDAB5WhSiT7Jg+duzuhRftNm8Fi6WB6Ov/JVLYziacZvfX0iKZJIP29Mca7xGaEUUo
rkeYlyxe7mGf4O55CC9fcemiATMj6hb24aYUuLtDDTlHXD4QohIDdrdJiW9h/KC4kHFAL9ce89pJ
iu1OMOSbu0e/2GxHEySsEtn8/LBXySvtCxDkICHKr/gpTbLTFZ56X1wJQmjQHcJpump05SGxBID0
BVpJLWFQOL7+oR3mYtY63696pI+cCvDEiQsM/RQNHvuBgjvN6EG8BQuX39PuubciHOY4o6yAehg1
dX79r69Wa7NR7EOjoDqp8AejbsDhr60Ba0xBc6uwGAB+uPhjUfr/ihcoS9dasvFjAmR74VvgYogg
pP8oceReLARyfEtY10coEsdq6BZEyKGo/GGOwlzaXAOFntj1QgFKvjC/FL36R//sDcrzDYOedx3S
JL8c0yYngPIiefWCBH4lqEz6zzMs6h8F0aui4eyfodMCS+lH0pSjrC8lQ4v4VYRy4gCc8EMbjBnE
c9zij4GXFXvGQBudsLdR9ArxftnAnvMzSoyKtWsAUO2Sra/qyzMgLXBhF22qwZnWwsnZBoVdkuVK
bZdRLmO/RpPH+P2IN7fTq2gKJyWOJUQ5j1iwRcq1WyzMg0YBX52+q3CWkHPFu2QfveguFsL708mX
8zG8AtH+8jUAPwHgHKgbEJHVIQo+C5ZfZd6bY0CMgJUlA9oxOGcBjHqP2xfZRv+oijfPtvdTFkiG
ErR1t5nGb5vyE+VfqLWpvljwVMQlx7Z13B+NvVeGoanU4Zd1aaHmNleF69pvX2dng5a4hLDukwtH
9fVjWB1pz8Ksm0MPGItgaNkVgOqz5QsgZEqp3o5XjOOtoiqOtrFDnmVM0+Aka2x3YspYGNyYqxCp
3G67Ix2NNdh0WUabAhmz6Z3wVIKG7aSeYkmkN3/DrR52oHCbfw25vLGYG5fTOD90+vb9DMmgxg/W
ASEXPhv8t94uA7PC1CD94YpwIixPSeHKsPI+8WiH38J7+LpTVgqccCBAm7CiEMZykLJr6Rl0u7v5
Ruxd7+UFEn11IyyzpMnV/h756N7tCVOokisXAignD2avo2v7e0riWLGzlu+MbiRUiz3ALUxYSXZ0
bCp7MAlAT2/Op8ainx8tAN2sVP5cI9o16EFYAeif3QcWw9La4w6Ew6w4CLfRt5GSnICMTWUL1gBe
RmzFu2Wj69WeMTrvsusffJo4FUFYpiSbKnHq3NbLyiFdkM3XClvSUTqOJ/Bi4J9Xt1b8/I3rnt/e
XZhmnIOSzoxc2J/RXXc4dV4wrd0uCU0j10zszwn4zKqt7+oBG5L7WJto+nug3tnTpOTBFcs6tj24
pd5LgkGvbvRGzYIA9jEI2X98UHZLZsHqRUL4lz3KNUAc0uEh84VkHoRw3CMbLACG0QTxWVZAmN9N
+PHRcanJSHA+qX4vHQRUYY3U1PJWqXYn2BFRHeOdt1bERaaqKAfvej006mWIC2jrwbTs5DoiBIUD
jBkpZtgyYdr7QTuPbO0PcBQ6/deOA1G3F7Eust0YH78X1H5ZOHJwL1Ftjrl/O7VrIYXPgetk8YMg
gm73H4+gVb5mO1g10V0pATrOiod5E/N0wU42b+P8jMQtLDXF1kfrY0nol/a0L5KLvR5Iw6pBruls
9eP9kpffzLzgiVHCZWNpz/5hxXuvzHNhSTwMCroA0+L1HyutaGcmSAwhKsz3+btl8DPJfeRXAQdC
QMoEodloYv2cRDD6CAWGTIHM8gxavYXSyLWE8q6JO3n/WHaocGdC7ovk7APa2o8Tl5LMhgLWYucB
WkrYAIp3FN5Iv0Qnvlz69Q+V0CaoBEp5DPy7s3SnPNbrpmfGCuAUCnwnXVwnqc1MI3gdgOlKRszL
75a9yQ+y8vzKIqNfn0rLcQSqccqT5Fq2mUNGBwPbd/9ETYzbXGczQ4AmdTW5Q3uPXbN6HWpgumrX
6cuiWvuNKfJ69AN9mNt0s9v4J54OwEvuHtFQz07JSlzPK0GPv/rnaKdIf+PcAy11uHOgOGJDFbxP
UPbRcf2cuqiXVr/Y5st7fCYRGB58SbQO2ieUkzJFdVa87KwGjuvvflsqc3jNDe+r20MXiUYx1RnN
7DuXV2l4gfq3vMo3yc0p9htYLd6VeexQ6/7JVoPHPa44Ywj6MhUPpmeXqP2KYKM8Zz1uPAfzOS9u
PCSHGAb6EAecqvAKqmVF7EG2f1EB6ep8oyiVc59h2u57Lkl8Zg4L6UCrr6ffS0OxqybF5yHPzJBB
6wJcr+uggOG2VF43ST/+tXFCwIqVAg7ZvaXXgmgh3yFiDJom+nI7koNQzWQjCECd8FpO9+qC9xli
WFUCqK+Pdj0Qj1idy8jJtMDZbgACqv2shalCZczuMxHwLb77/9/24z9+0FviQ7+kcG/uBsaLKnfW
QpnqJ+HY0aSXS6AxxOMoccXgbckT76WpUsMKJ3Xzt3u1w94KMfStt+f2Xt4DkfzsfaAVcHSbSJrf
DsgYjWMkzDHgGqJRYBaEbEmOpXw9oVzl+eMVMgHiu7bALlpWXD5Uce/gIf29LI18S9/h3kC+E0+d
E5e9c9OyQh8FLHfWJHM3yNTECfFVLR4ksaY6GMD0nyt6vNYFjGnerYLcWvwUP6jI8XW7ThFasYFh
UlnLOTY+5DAZ8lDZRSyvkQPBuvM/3XY5MUkoCub4oftNBFiMGIZpvu0B+r6ENdaF7/CfZilNoUxC
prk9g0F9l0AMIjiu0F8kRn9sfSE7mzFo7uQl9RkfDerOJhjNHAa8rb8XbTyBgTJFxxRAmdyANpqI
vI+Soydz9PRwFmct02t8b3ThlmEJrHeXma8Q5RLQwUn/W4lrjBtujW6qNdXhgg2C9OiJin7F6sTZ
s04L/mxx02P6VXgYjyVw3jclxbmXpJdZeeXCBuagQ0zN9FT0OD/rYkAHEFbwYMifNDAO287f3+Yh
z5GVy8Cc3P2PFodZK2smDvsV1uFDbheYt4Pw6/DoFx1wxLOqdNA3pP1BLosqy6qoCh/osERldYZ6
xQTJpNl1eo1Ih75kBKV18UWyF5UbED43DwHUc8n+8gfErDdy+5Hz8mY1MKW3MFyyh55UZE3em09y
kkuZDbMQjzJ3mpZ2SlfkETroqnt8jWkMXYkBU3IuNGcJmzYQT8H7i22iw/jg3MDtn8hMOiJJ5mGI
Q+US5yFhOEHp80hEtmCxICoFY61mRNBjsanCmYMqbEAnMjGx0BH3kDQo5rJZbLyHElq9NBV7Qfov
Q/RJmLs2NnVyMgbgqgIUz1TaFx/KKY0BfsfdsRbB8PyqRoJVUD6BitqDTeNgXRyKhhdh4la2VLAA
W0DFZ9s27VhKP4AQxTFwvKgzsa63X0eAia3imHHKx6PD/Fc9U2VZg6YZURAK+g5flFRNkTPkaIXW
5F5hUMab1XsxqB/7Jw//Mi5vpY9iVrs/X81oy1Rij2KBb/C496hUp/FXrO/wtItsPHrl88taHD1i
7qPloGVDmWsLqpJliUQRGLmfzlPNeTFIR8j8/N9Xp49McrtRfPfWOd74xdHrFnqP95DxSEr26uat
mK2pdJGCJHOe+Oy+jmABpRDf20qrGDg8ELpSZ9eesrSkJXpNCfsiHt5z7liWiYh/tv2tooqgUfFn
TzP9pYEG50hYSmw9bjJNp1CqJ9NLrUl9HgP8tK5NBJdFX7wZcv6pHUwAkjaA+rXtoEX0R+JP/v0F
c+UtW+LhqDxomwlkiK3kIQXyboSgDCg+al6lVtOq4EfZ+zsSekBXUnk1R2ZEZCORyCcl9vNoZ0IR
Fcyy2FdOgiN8EXw1xg8Xa8T8NiIWqp6iUKEzEek7N+oIXXF49s4FE7YRzouiiQRsSIpxoa/o1M8F
P5rc7nbmn+YsYuQFQOt8+md4/AUWNREuzgX7Ba8kmzuJG2STOYn+RoGleSbTurHnbz3y+/RlyaYy
doTXkvOK2/yx4aBd/UnFEJtsc4bO8o8mtRz3HNvjghWclEbUdUERfRcY5KCYNtKaugTv44vnAKow
MyanWWqKdkluUGV+UFtV5mL/ojMi+TBlxmGYJm9ux/0+MZQ7/lBENxWsoKxM2irYRgzXlHvJaYsV
/8L5FeRQzT0PwRj3mcLrR5azQPLjKKfqSpq5rez9EP1dYF2JEhWM/DN4pD8lyaRveXmXDngCvY93
/Gv+f2ZlUGYCyux138qUfbYS2re6eS9cGuNHRpP7VcT3wJuHxUugT4shnnZjDee0ej39jIYJvpoT
YrlX4MQspE3JG9G2xcF6YI7KEuPz9OhvG1CSNNkwLW6BhiUF32t3nqxKFS4XX4ptpFF/xAcJg3/o
7Wi9fXDJejeSjBKaYTT22I0x5mN6tD/pAx8nU1iyKz0BWme2dvi0+Z8ZqVhlBE71l6BA0K13/Pdx
q9/8BCJe7azp7SHINwg54IppND6tetNDdi3q2wGs6kXzCztpl2IN4ilxSWdEiGNqWHofRDCY9HPU
+Q1JmMdwNRY032KAuY9l4sCDG7WB4cULV2eXQ44muFZsoODHl1oCTfbn9u+yMS2QXBASq1OfjhaO
IYzhoIu1BcltrSdk5BV+h6fLV2P8inZAFBDx5RAVpx9m87ZqQ0jK7PwXa+NvP7+sImMlk6bxJbpy
RRkjR0L0qZ/O7BKil6vqms6sjNBbCl71YL86BanrykHZTww4jOMLj3d7LIvWSTbrVgIbAnPKvDC4
9cLNspczKgHfoQ+ExmGrW7suJ55TVs+CcqWaNDoL6wdWL3kng/aPIFdQCo5CAShzKADSirYc4FwA
YnzyoTi8joX8Vtq9MGnhSvMhuzoryZENKqBli7GeJW+WmleX8qJqs/aEqMxpOXnMEWfsqRf/Lqil
023FQTB9lEaw5O9pn52qFv8NyK+cQhQygZ3zm+pRHyb/LBd9X5eJQiYLmo58zWDcahYFZbHsKoDl
V/6+EJAW6OETxUz2V+LvPnWiWRAhqaDtJuWltbUk6WBlMFKUOtqsqr0h0SD5sGVSKzUL9d0VNfDE
urNNaNklfu4SfOgXzSjYAWISrlOZwpETtnGdCOY343HjXECx4upAxH6P+IAp48a8Uh+y6stzQELk
+APNo1/txvSZF9PxdYPu55ir9gMTo60cywgvAj0/lM7CFuvUdGGjJzYCHEnjCfhUHMVYw8XBYzZA
6XITzSnsCW0/xMUN1f/0NCMw9z9bHUvD5dt1l2R+AXdd2TvnZeUAOfR+wt3PzprGCda/ZZzXmGgT
JbejJ9PsY4LvxhnfQ1x6As1tdZzutjMfSTdjhQD8pOgRoLCInqSDNcHw8+tU+0viHBvmMHhD6SCk
WRywpgNy6nrRDtjaFXh28lFLEf2ZZs1hGMHSkBFcVtAzVP0/oONHSqPGi7q2MlCgSPCBqSdR2XGy
fBLtLJEi9k/QU1fqvpsx5S/1RLmMHchLGNSQ/wqFm7SBf700u2jO9/zx44BTMriyGTX2yrOREDzj
3zisTMXm2k86fEitkW4WqKe+Q2zHtFgfcZ6baILt2/InfEGkhad0b3OkzwJbptvuPmY+O28ZKp6W
KEU2pfRptrCkJNpkHL9GChooaGg63CrHR70vC1KYR+ggyS97ucrCJJBTfa3rGw9yvy0S5Hh4p/cN
d6oSs73flZH9j8Ns6PdYcMD82eFNy8WLvKkYgloZtkB6l6E+lQb1Hp7AJqxYx3g3aDgnQsY0tWqa
R7u0z/dMy0mxvvvHm3DribZkh/dA+98Pn6WknAKvXbxRuSvJgbSeq3JCWWHhRYFCttuOYEzmAehS
AsXDMi/BsCILA8MYaMIK9uuOTEze6vfdZALpW2utEui8Vn3+zocawxVEChbnHYMcsAT3BX+kojIc
+jvPr/bTVFFJYCrKe7b1PQfTc4qUZAhqDRnqi7mNaJX41FJ6tN3zG3BnLA6eSJsIn9goZ95jMStQ
qyhJgzxJJytkr3U/yV7t4PpybUqyA7YmQbaTQPlXEjI4hG73vn0NA4CyBjKX8J6yjvjkUpDFWjOD
jKk3mmgztx7ID86kbj1sVKIIcVssq1KM9JtTfu/VlZFHHnusYcITuhx/t5/iY03Dcw2hc4anlzbW
qwppLyzQG/jxqFfGrCTRZWBuzsivqbucbO/gmZMfMruLXm5eTQ5Kecnvo8GNXSYv43CldNL38oTa
2fQVGIDBh9ja1KqTPG5Awl2aPKC7zYRg8iiIp+S3sut/M0kG7vwX6RC4K8YRSJfKrNNQlHs2mfb2
HF2IBSgyfKVhCh+tD5vKNULT7XSfo/Y4j/SSEkyAlV0wmAYaPhKFCRRFMp93unEl0K+k09HAqSQ1
oug+KKlJskugk0AacSGNcBMDWNAVWW/G/22EO2GgwajfpL8tozj/xiaA16oVURQBsnLGU2bbzIPk
uL8mNxmejdBNux9OkbupdCqiD7HCOBUmBj1yZJnbHV1XeR9fRsx68FRn+pXh/sjvJyjRvZopkT5s
hN/ocjJEedi+7jSV8PM2XQFdYjPiWMV+id0pgvjyhbfb+t3R+uPujsozEwSK5QDKKDORW+FDso3W
JCFtfJiy9a6/HpUAuZu7U4TynGgtrD39zXMybaeLFTfvgeFHivrsH6Q77mt1rchCf/kwaJGd5sBc
LRe0VCbCeHmaSDUVkFSPY+SxPT+p2r/FfUNfp9JWjtCG6r9KCyYVCQQ6EjaZqDJlb4SawEcimCcr
zEkdTwOaX92cxQtRjHK1+fPqxRrmt3lPIgb/eMyhw5tgZnzVRi9JFZM6BtNjqhzTZW/c4m/OoZqh
Q0zFlTgWCM7gvHUCoiJo43vHhdK4RXGjKwB0lOBsrL4TtWJycx/S/VaGfyRgW8nfKHB0OJNhbhTY
94mmUQsdbjVmU7J4KwUMSoOVQwc5o8qELwF/lKBbcljE1O7LlW8ycWGVXvKt3qs7Y1aNrxUxC0K3
Psjygq7yHgl316R69mZ4md+q32Zg6gC5/VogFUQMIRtyna/XFsFS7cAWz9lhJSPIliE0EuwNOy4C
QF/Rt0ytfAIzfyGbPU7d0Gm4CHbIO+KXPqvpo0LAstp/c8A3xDTOsnB8c5QzG46KBT4xJMNd0sA8
qVGSqGWVneWJeaZbTWPl1Zzsjq0I8Ke0caXUjwiVeHkwmP5Rj7vGEISYougtRAYh+WHDZozr1EVB
eRzsM1waq0iz/gxW7CRcMD5UDbl2ETzvqO12bE3WqK5z5vzfSjSEbyzku5iEfIWfOo+Ht47UWgjB
7wQop4ACx2jR2pmow6QF6buvs+riOSCXsjyDOytURJEf06xa5q4QpKcXgS9e9FJu30U++l4uT+9F
Gw+PWN4saSNF8qeGYyfTa5UbBVMgnt2RU56y1K5PSvmh/MqOpvRVM+b9c7rv/NWfs634Ot/qHJOY
W+k3vJQpQyXwp0ZQKDKKjWs+s+DDVVRiLvMbfTGzjjVg6XuLXe3/sk5RHvaxo6g0Z/F9zG+Gmt+P
p0RAR40TzzKnUcDdTOtc5rzTLOhB/8wTBr0D4sE5/hEV9obdmr7iYIxeR237gY1T0H5l7Q4fVs+C
bbFp4/7YqnbsYaS4iUJnidfuMeQC2pR7npnVp+hH3wYChIwcg6/KEpjF0TfkoUALCTxXXYWYM84w
7SowGeuM2rHxJxQIScu+nXJRb45/sjg9G1Z++LlKjqwzEt54s6aVGZYf3sTZRZocTef6SRE2gUEN
uwVCFcravKA8PmeHweI4m5SeXquxZy1D9gW8lWPe5JANY4NW0v2zupEkRNKmMcht6V78ybBoH5FM
1+Hi3o8m3RixBJoIuXUjq3u1q6Eb2OyUWc3AZK5Zi/cpOeSF+2trV2/5BRgCS6oKFQ932q5B579a
BZ0GvojuZ3y7M9WyW0OakL+72dXn+LR9PnEtnieaiUqr/AFoOAZ/LKkVITqNmA0/L+phicuI4Q78
+nrgKvIrEgMTLE09MT0K5eudy+naxnIM1cB6FezshIedZiRqDla9m6+YzbqecVVfSlpwPP96TyNy
AYwmb0kfnf1Gg6eIG+Ydi71OwWw2LzoucU0wuMzngIs0lpwt6z0GbWMxYXW2GceSGYBRpAMGR6JJ
G+aCt+AjkjC5cjVERCZJSnmhZr9P9FmGlJHo3/b8qUijnqEjfHBb6YC1QlCq2XuAZ4YjSugitFAP
EhTOGRjj2H7AyYxZEqQAnBMB0Z7lewhYuprp1THyVzs/VqUcArE1GCMfRXT1+g3phAX1EuLWZ+aP
3QC++uQy+6+i/ftKG0PDleU4rL0ihE5Pbkxijq8258ShDqo6PESpZDi9skggTjQMwkYsghE8mHBp
OklSf1eLAb7fRXPrEohReP+G2rAv1/2P8vBvDEXizCHFYCc3pRa/lemU3hgVXCe5QkuQWMaFjjDf
KcWNlQ55eSVsn/ro2rOP+AvYFn7rpvIRkZJjw0drZ1qvYw0VuGHr9ngUXcXriajo+T+BZ5O4alec
2ylzTFaWZL8lLDYF/lnBgLxITY1+THeKux+wPnJ7/TysWgZCOO4dZV30xQkCTR8gAkl0aBZ6nQFz
iN0Ux9kQkyEZ7hg/6/fq5yqmSD5h/dx3lv/ItCdrdKObCs8HODFAKUKdrfRN5rO7P7EKqIfLsUqM
vjNU2UXMw7uEHMNC+USuarzziEzZrrwAZO5F9wwZpupI08lsnUvsz/rJTPurV9cIVb6704QOYzvV
UhCIZm4yuXtSJM6Z4jgIw73MO0GX4drOr81kPINN9MnT5Rjw/Cu0eO4mHINCv/kRvoBpqUEcwRob
tRoB2APP203LnoxLf50uRTiP5JpVMmvn+XVLtsLRkMBH51azF97kfhu2gssnG+he3y0mVHOguo+9
VbIzuq5D7iurSDSIziNXwatuPh3r3Fz+SURl993j/vazVoJUMjhobj3OJ8ZOPc7Nd6I72OrJOg3+
b5ayWRZfkp35W9CkIt8cNQUNJDHgrDEVe+4tEHTFPgyEWWIDzSEMKlfnZFAK8su0NEbBF4+AdJnw
lh+J603mYV5RQ4WL92Hig0xA+axQ/UG8LETcX+YMZV+o1posL77K3cxHtlIxEGZ98lnERBeGwvd6
0S1Sj9gbRQ01NokvMwmE1eOo4LwNadts5tqxlsS8xzdYaYxpdtYjh0iHe0MhJPP6fo3ErQ0V2Sj1
ZonsZR7YDpKGrg+KANtFzapv1vKa5jPd0AhAQKTJFsJBTW5jYQcDlE1csBQmfr5JJaYA56Et1TjD
Uca2K4+ZZJhPhJsRqfTLtXW37h2mPfR1CpeZgMR7s282azh5A1droZuooSuN3n5IJiNIsmNKJuxL
KOx7mD2oGXKbtEfxyLJKcC6EpCGF31xB9XFSBgDYK/8GZvYQDIitTMuqewATixB5STXxR02/X3cw
4EfBpmtsZYLv9plBkLe+1Lc0j1F7dKSLZ+ncjRSk7tR8aWrdBRcaI68pKM4e1gyi3bAPLUZIi+Un
clD7cibSJyxeTFIiV6dC+xWA7NWsSMWx9tlzXt6LaiKHXHYY1p1a+0ZSDzAnM4xUfOE0K/yq0L2Q
qDObEpnk5sJ87b3pTR1qQ1O7yi34ETzP30b/PM6Y6T7zpFS0jYQTUFu1B1IZa/2XPsWNptWJHGRY
ipYVmBFzL59Zd5MLvtq1RXs2kgY7B9tpXAe8iFkJAgidDBNEuGBFaNTmwh24axa9SHeggujd00Ux
de8ovWLK6vMfKdg0eV4AjHEJ0wBbFIjhVJglE4jIJPdy4wlcaopqGefWCYhPfm9Pjt8VcdBpZAVc
Aw4gDK9+2IKXzyckkb1DypnOiRf4EyRlh9M472SejFqBKv5/QhZw0NseVPoghef1qQQk94TqGf62
aol1/GJn06SqmYz3y18fW4dwFLqikb0A8rRV2kkxaKLAMpmZ9uqcYMf97SLOtlAJx9lH+/ZFNC6J
SPkO+ss10fiOLUvoWkryS6Qv5vaxF6YxcXmlLysxzEFGZ6zmngAk3ZkS5934fwZWmZciJotdyo9q
+sZTyNpMV+kA8d3t2TGcQTN/KbEp3xeuhxFu6jQg3dH9/Rb2LAHsdI0wR2HMlGkgapNXeJpvYYue
YvFrFK01YpSKvQyTASZlfmzTJoKfGBPApZRMTH1pgHaC91bCPMo9KZlfgFigbIhbaS48WJPyIdwf
QgZ9ZNxS/QLrwv9uVnOc6oHpT2ZDavVb0c+7c902X6DZWbN1lepe3E4H20CTgjsnLkaAd/YjXg5o
xVi7/TzAXcuHQ6e6B6N1kBQMGdVOJBlkSu/QUpxutG1YmWS4tZeaokwFEMt301/Cf+ijCOiU/XGq
rAL8tTgp3XKPlx0hzfNnOsYahYLZSG3OpjHX4Usn7PshAHsYXV2uIrZOzoxTaEe1hb7HviyaXZ0M
AviteXfWCJltCxoWBKPnEgAxf6aOyHxP7RIG89hPT5aypOplpiNaKODuYbfz5S0F4oJ7Icr6Us40
N7zTSD1w2uuEah+7BW56SdwlMVv0kcrn3sSIpQxaKvA+r4dNsHe6w9v5sMNjObY3RXVP67cXBn0u
URAEEtWtAlF5vgRVCp7P/iCSBSbHaGB+4DAofg6eCj4q0AK4CUClsMcPGhyWE/D4sA3o4oNeImBi
InFEnfsS0IddVBeslQCtIvRYWd88tN63ZSGrOnm2N1Ngs78hPNXqAs8N3BPQH1NCE7F8/GPFi99V
R4t7bpSrL5kxQequL9FREHIgW2RVjR0lfgcbwAHxXscrZp2GYiKMoxJE4BvJCWlU3kGTiLgA3dsk
CQ/BRAGEMFW7H0wT1Kjc7bzN9dmr3fjE3wIG+jUr4JV6nlpb/4lHpTxXBy3zavyCNUm7Hk3pBIlX
3Gi4/qeL0rj6Xt9WA9pAipXNoSXpMQnU5PDv0CNOBnnOop3nxQjv8QUfaVTSxxJDexjWE5Zz3Kfh
vaZoH8Va5VG7CzU0d5BnUW1nX9RymChu0DGNn4dweccFqZy7G/pQJnIXQlqkKwb+hjH04Hce/lO4
3Lj1NhT249wG4Nh4TlBNi9AlCUBQXLdljr2aLr8qFivRE09/wWyVS/zbZui8yJzZaeqnV1rHMfEK
e8oZqpNfM7c8L6d9sVPRjKPdszadcOh07LErWpPxemziVNB8AV0dkHwN3jTDZmSMSTnK41c8vecp
kGTAi78YxJK2jdbP1HKZO6nVBiUEPokJ6yGczvaiINiraib5EXZo1NvWUf0uuw7dkKhHMyvyVT+U
XdZ6vuUlYt6pEzTYaGT8yNF+8HOnGPs3td948ZVCb49pU4R7Pezzt0EG8zVyQbdo4EaVhl4y2PnG
I4P65S7j1gtJzeNiZuBXdMkI2Vq8IwmrHy4+qn5qHbR68VgJGhtpcTNMYaAyUO6cLdEWo9l86mcY
JZQwn9TpcYRb+ZRYaAacuxFfDAnMtmxJlJTuxiglchQ7km4nW3dYBUv207Azk9wr798Rar7s1ku4
MeeQ9scro7At9h6FLwcdlhcXsF/F5GsLNP/AxB9taoyBgVKu8aNdfXhQrbgaFcrRdoj5MXvWGfZ5
rx41tw/FgSZB9P416UZjpDovOqcDVoc3yC/yzwUa2PoqP6ZUxE8ltYnpuH0+rmEH0pNxDeQaS572
en3ieN+Y7JxAKqkV6ZitvToe7If6OsPIuLJZ0FiIXEYPcpdg37YCY8UM4+T2AGpRlvBd14BMDhWs
h6VPBmDbFuGbq4izZmk7gYw/BwhEcYh5MHN1u5imLaVGI3ReGKNeCEa3i5br0ajW3qEqhjvFOamz
jU2Gx9LIM4NPVSJCmj8Y8Yd4JEXsJHIsS9VTEpTL5fSEOQpDQqXpwnhw6AFDymlCwynWxlNgzmGr
rT0yHOCpwxLvTUhCm3yAO/kDo2MvvO2qDV6uTsz6OrgDry510H7scMCglOAifbVQo0sYPOhe0QgR
BdQEtUKS4Z/w8ewvV2353TEedr6pTq9tNAbAV6lkCCP9jZzG3MXbDblNmOh+WM4NotVbI0iwM9R1
3kWeiQhwXZS9ErbVNtsGyERJ/u/vbnYRectOyzCTV/PHycEH00C3QHixJHZ4RILJah2hJG/8iOJM
v9ftZabCfAT2PmfDOyAK5YohuPUjI0WV1FqLxd2Nmq4PshiC6xUAq90rtwFMiXh36jxJpV9HXQ3M
JaQdAPQGokclsJ+716nEh4PcfXzrTDMshVfXXGo8/wCuHv/pJk0FKEn0kvbxIIgkGqRkNaQiS8+E
xQ07fYqkLRFnDahdJzZ3MVYI7gwxvlzey4jOS0+Y3xBwQ78f4csQnSdJs6keL5SEeK/CmCmbQkK5
Qrxt6FXEG1oypszK5KmAKgTk9InjGSReabVC2GKFJ7p/CmcdkodUrb7l0cUPbA27D6h0mCZ4FCrc
0hwwDq+FL0nf5UYdXR4fqWYGIoG1J9SmKlqSsq2v/6xlfEVzqz6pcQ4WprkasQeGt9+FRmQW6DtY
6OTPvDjXbZcUWO/vMY+1ZJ5UcfWgbd4aWlkeUkhtUSMz/eTFgNDb9RpcdqPT2ITMnQA+13W5+R4h
J+oHRVRAS92+5+YpARV95vwApCJ/kcxMI+1/MBHa1tihMfYbssTW2X+BULHlYLzIKmvGFZeOyEei
9dDqkdu+lBxEVQCQXXLp/slte0a9CpJu0WCbN6AdEZVW2Tjl4nCHV8EN9EQyHsW7Ni/T7sLWLxOo
5dzIsCl9SRqWf/InmKznEwbZhY8ncep3iXUDSpuxRZQlMU+etJ+EGLH6WfvV5KrKG6v+OnyDKXoa
v+hgCUkdnvHKTYd9UYyANNizjRqgO1Mxkw1DIZVaThos1dZ+tdxqRfc3MfCyfHyh3S9NpWLljFft
5Gz9jcNfQdceGPs3YPvQdHGFK+yg/IIdtnlU/RAaQiRytno9nqrFaYZ2GPtkiC0Oj6vK/CffsPHn
sDeO5Har2SvJevPkKL2ZDurWLjXMIvZYzKbbvFWyMxf5QaN5UsrUqBHrsx9kY3CRjXZX0TxP6UPM
zM7yPGmcfTcuBo8h4SxoUxJ2OaayR/SnFKVboDLGbnc1lUwl0egb/hjfImajNqrcleuFxfI+77RD
HTDsIWSAw2U1KJCHVv+VZIvd46iGiZm54V8MIz0s3Mg0xegjJvbQUhA2Y3g7lFNmL+L1axmj+iJj
CAuODfw66C6/DhA2qLi1O45CM84/rAIsnMRgy25w2r5aU2VJCQKdArEFUcFXXgzGaWlj4kYZ33V9
60htfTR3zVvqi8j7PUiWvZ2v/3kC+n0OV5nEicmfAG72tk6U6Smx+JWRr83MjPnC4+TW37kKgRC2
hJs3l8+4MUpc24Pu20WSH8fLg6D9AgpvN8ASMIekzmHc0jDTWf/ZQ5DxucOyFMdM0jldTFxqGOdY
wgVV7p/O55BHvzKOqkcM0AS2uZBRVluKRw0RXBcVXBo5CiEkRUa123W/Bh8cgV8qjX93BNnKFjEB
oFOEkkAOXPpax+zgWdWwE2AprZ+ZD8FZxjs7L3mVxzhcWNaXe7vtfdRvfS3qNY2Kf37aA3ZCJbKM
anbuUxTL1RQnPHSdnPfSO5HXsoFaxJ248YJnHWjsNxZxrvRD7+BX9NLrngoRgS/UG5eFsvvRWELu
IHKe3k6QnBnLdkpilOUq82mbTGHZPiUz+Kj9iSwDNkSmSWJYcb2yVWhBP8Tu6q8zQa5LX4UgnhuS
0kaptsHYWDDTfKlzZqlaNRCu8oRBcxFFLezF+vS/LtHb17zQbaG1d+G70vJ6y9gm69KzjN0vOXGB
sgF1/OX+1MKw/Ji5sRbz9kXj90QK2YuGUW2DAQwmOpbhPgLCDD0YfzQyaLAhpxw1zP3AfFxFiARc
DApPqKyRmK/gJgJ2aPFJxxYyF2YMbu90l9f11VYf7Y2JJ/0OU3vjRd91d1o9LXuR49xbkkA/4Rqr
ykoBQ9zk8JNwB0OFHeNIkj4LxS/oD1wKT8Pw9ZLMA5SwEgmQnbRp2Rj236MttKWWayDy5Z0nl7+S
I156kP+nDQ2UagbBDajkHpv0gRqhhTrDKSXeoCeMlO+250wAgErTiqbjgrGPQYZryJoTTB31hAEP
KPspw694EfOJ9Acey0dxK9LOM4eZRvV09OKggf+7z438w6IECcxJsjqO8Qc0SsVYTdpRSc0yyZby
6+f41b+7Qe2wvuVKgwQqYbb4eJYzgi+OTRCjsRUCdxhxhi3MwG/5LJ04J9993GYNdFZRMW9J0Cvi
ZAPGbRpZGzzeZrTTpf0WGUoqbRaSzm8cidd0X+n21i/GoqM/SncQbtx2evdhF77I1sqTXC0Yujws
YNNTf+Kx59csdy6C5gUtXLwU2LPzsvdsBk+rPwpDQkF5Yh5GwYRBMpVR2fu9SvtLwde15NjRh+va
Vl7bF/ybnu6vmRcWDqNlJnSb6Fy3NjTwoRD+LB00SwinqFkSU3D8OxfdcRDLUme8K13LX4SGoxJV
92CNVfw+MmSOOGWFJNwUeP/ubBkF3KcyoyaZKQmbmoia5xdXLyBG8Tusr1xMau/Hjo5weIBCKMrx
+yMt8oy7fh5yCwRpNF6jjregO8adQYZl+yoeBT0Lc2b9BmQoQv06DCk44md2BZPCTm2gMCnhLAbI
0P3nnCT1I53BJqYLrkWniZiKBSk9L1KmeDCxdQIGAgRXuKCFJRflwDx1FTBA0ve9EtVUkxPAig8M
8gcqT50h86wP9QTqcUauED8AGgWv7oTH79SEqFWv3AOeyAEM6EV5Ka3fUYYC2D14HtlzKzkKPquJ
mZwwyUm1O8/IR7yXT4qDoDi4letIF1PXkJcpY5mKKI0HYITMUnWEz4jSRsdHBa3IEtIf2A9hu7IU
YNABiNtPN0xmEDZFfwBWUU2Kv5+e+9TkHbGG23WWpzAsAMKeRtlC1XONT45ft/umFTYbosXCXziv
pTIiERMYBhqGWbEHceqVJdizwzY141Xtl8bWRj4PoUQj0S1l/yat8s0AWwUYvsK3Q0WKZ60IRm2w
cWYB87by1qSnstnWbDIqPSOokwGFMG3ufBkJ/MuJLb9SOgrnuPgZT0qHsjCTfgzEMUiOWMqkOiaa
t061YK5GjgiXxXYWNvBGdD4BjS6dhr6NLH1s44gCZQjCgpLomGZaIGlC0Wa7BeEPKkfo9ONCB/vp
vS3beVYkGhJw5aA+A/o1zLQDX9AliHnlLJkUEYoeMVip2X8qRhbmRhpLFSyHZRidTMDnVRdkUybu
AQI6vxRROJ7WEvnbhSu6Cs86DOETuMVCHlzVBgXFXCJBGzIX0OApRT0845GwrznsxcpH0fPxseW5
oOQr4cTGMVCIOQo3mTlbbiDgFuVr2GPj7WCiXk4jZnRN8MeX6Gf8OCgpcnFu5FGIKiHdxoZ5zILb
tJiohP+/3tHsTFdGvky1Lc7G5O3pgz7V0CRon3mLwLuW5MTMDd3TPlnLEM+ndLr+1UugIFj+s0WH
GtMwpfUH0Gr2LBZhLhqrH4QpaZyrlue0w/emA3g9aXuT5gLW64yV0s+Qo/s1hXM9VnJZpJWJhff8
t2VVknUp4hjxXmQKlZFeyLpOgQDoNDqkqPD1TcgpLwIC/kdR834bcCqH0IVjCZDU9K/4yniqNJnA
QF/xg6udZpa872yFECylYUlkaHwzmQUJBD0Bx7kdNfxBjqXSQz5gwsYMCBN9v++46DnuG5w72KC6
qGmMn2sDWfwrgu5MzT1zu8trVHHHcT/CN7L4Kdbgio8TVkNSHAyWXMJIFi133t4yewKscI2PaUPV
mS5mP8xMDCiQaIeGXWuXsu6PIvAOub/T1eBxeL/8AjhfsOZzt0m/Ngt+UQwgo3/Z3J04xili0QvI
wPh4htNzCh5Pg9nf85xGmiCG50RCPd6Bfd1fbP9UtdoU0uWNNIdbXenVstxishs3I6L68ifKPsQV
K8xa4dCkHLpyeaUg1t0FQeukRTSfCr97q4gCmxL9i3tRdEHskzYSpMtUFBl3ECT8ujDn5tIGkWlI
NBmrNpNppVyKUD56dxEyLLbOuiLkasMvPInBGyN+dqPD8d74d7+Smu9kTxpoFiqHsfcB2uE87bx/
tJwhgU1JXvMzRXE++2CeUJFxm1bVcSec4lhqOB99C9kfi8nBfQYRaMYfIHkHxVkDl+bMPDbgc85f
VuavxtKwmXXTPb9XCqNSMCtJyuGBR4+cJKVAd+Lf1acSh/9o5Lvx8F4OliYh1qAthi24CSIJTzkk
hFDQ09YSUMmckkW5GCMgfsQC+oGLaBpNlhbYAdmbZm+Jn7K+3BY694s5IG3KG4G+VOv8sb8jYQUq
KimEIQphK6a9HzIF0yG1z0QxWNDHrBYKppe0j5LoH+uEP016ArFCY9co8mDCXzWxRc1rmFt/HX7U
Lp5y4NQSH88fJ/NmGUqhK2fOHxXYx/aboya+oJW6ft81+w6reFGqWtVsu/GoQTnKm/LvN0EjEB/C
mYX66AVTnpl9y5kb5i3NwvSllo+JMtt04AgNaHZck1E5+YlejnVYj4NSQIv14YmQrJNkdSKLtEyy
eROfDNFOFIh4OcCRvSUmrZ15R2ScVQ2Mk4mvhpInbAK6YEJsaanhXg9d2l+V6CQ8LSHJhAroWB+L
O+FMiI7rk0EUCFfJwtLKF7mY/zBG7FSq33WFpDNwd4RB9ZGsL2+VxKua0CYUJTGskP/twFQW9ks2
Q5oIm0G0Atse6k2jKJ7LxPiMpfue60nokOeNzSMcMYSyvDAEua3dATwk+NrZ+kfGAMikBW+oGZRM
WbJ9reX/0XWflwG8krf8vlFknzjwHrvAZQishOiObvRoG4VqpnEkC9I4rO6NjVEEdEFojuNmKA8R
ZeLShl4WEBx9Gv0cQ6L/jAr7Ml8Uq/TFdrl+oyJVjKcRtabaCQLFRFDl19iZTZq8R/h9ckkzTczB
+bsm0VJbC/N+tj/uhG9l5MFwUmn7HAA3eqeBInoQY33L5sNUg5Hl2bYmr3smRr8OaKcJwbQk8wBl
1+iuHcwv/a3wrEMlDi4GVSUw6fCSbwPzTemTkPmrnzpCJL8wOZvJ2/SuOctm4NpI9sSMVXggW4aU
z9T3wEbYVf/4QPnYCIkyf6FehH4XOU1wBg56LJXY2mEgYDzmcknt38LsfHy57gWGsxPRylecd7pt
z2/euvr4FjePFLYXL4Ty7Wzu+urXLJSIcYSieSDYoLNgbz38DTuY54JcqvDjNBPKIGU3dHsmxdug
FCrzSGpvnga2iuggLovJURVdSVP4cnNHVsuq9qLnbo1Q4u16zNmBQoOAWGmDCyxUvSvjZi/IGfSY
rnAKlPGXCoCM+u8nDSXttWnRlarJOIW7Lxv4Z1HTQeIvDXashcB9HdU8skLTIixoHCqJaWlv3HbJ
7k1h5C8I9pA7+RqbGrI4dgazOu1ZIV6pgbw+XrAvPnl6cAQzRf/It9k91OjwOPiO9s40dvAZKZyc
QKbjsTMmKq0d/ne92HonXzGDYAopD5/6wuVPKr8rEjcwjHMhErivZFsf+GkNzdk1kMtKEb5407lY
fYLrwa09wnbl6r8VzEgNllrPRSvLgrEPxlP4099jtllu4EWymSklRswkoj5rRg+kU2A0wjZzRGwa
ogyNxuEbWpRr9auGno7lVi0GrEKmEcGyEWKVJi3bgPwNPCwXRONbAyQoV0HUYLsdPt3deGwGe3x4
1QGsg3nMP+jOys61f8gxHJ6Lou9dCdNFJPsw9TfGt2Z2dnJer28UPNh2FFy+m8C9zeQjbhZwjlBn
LqSQdIqxYp52BKnzXTmlOwBvqI4OK3sbbWPXT1YCuGi0C/44yPKY4je960XVemroLvsDoio3U7CI
HaVQiEQggQh5nCC3VtIBRle6hu/2KSOBkVFKlLRXTyVwsYjeQJBOS3RnMgjl4bBSR7ckMupT5Pxe
shNhKp/nzabj/XoCVi4pC34CICEMZ0NZ602X0jA1Qn9gyLsVXUvcV7xydPwtubzSleHdLTLaL6BI
5DBSa+Mq/J4oDa6Uji/M2S/oMxlGqxdZo5vpL2mCDRcaZNzesLUiLm9jV6aMPu3jnmazE1lSjgs+
U6pLb40WL4vY1M58yqdht7HvTvYlWctrLyUHrEZZSfXA9g+MmbcC6DFeM+TfSbQwVc9tl18/5rfD
pBCvrkS5m/CnDhnB0qYDzZofhjMP2b3b5DdPAazsqpcYYiUEDFh/j0VvxZPflfRUt0kavxAWeiv2
DoHtG5gc3jJaISOs6PsyDlEyS3fn+pjZDvVYmGtGkgq45ErDSy2STpXMTbn99Sg3GJ9lNrPQxg+w
pDHYy194KqnlLbxNMZz9uUYH5KbcypcWCcP/LLbSXS5qGcuPcbbgFkLdT8PYCureOYThqBTaeDKw
k1TLVyDwU/77CUpKu9JQktIOEU5UbnkatyCjhYLZ+AOGAZggWtq0FTH0SkRAkS5TEwMABT1TLHjq
bNzECnVaD3Fi8nfIwwiDvYGyASPSfgho1ZOgwtz61Soa6GyPMphLGib9t8a/YaM7u530pbLSiFPu
iE0MXpbLC5ttUSE08G6MW4fX0RYYsycNoCl4rdPTZGGkQCxr8OeMtWbfAKHASBwxuaXKeZbAp5hL
ec2vCWyWaCPjrljXDgnRpE27z1GirUhFBSGl1+Cz/c1/KuZNNawP1CslV+aRDgK/5lTcXI4xvu6J
E7mQdbZgHndGhSJwvr2WY6Lq7Urdg25l/Nc2fGnHnpSWTQgszgT7s1goe7oMXPyCE1TcEGQyMKqS
nwj3g6vrcCYomswm6CuRpMxn4z9spbRGxqpEf/dY7QgvkvpCmx8puaiXXx19vhpOoORD00ySmbiB
DKMx3CEAMbd8mBu2aOF6DKsDK1Du1exAv2KW0SkcV5RRaJJhgFuHzQ3kldHB7XaaJ7dHQScERxlW
UF8WUPS9QLDwlMbWp22n97krRvkqZT0bw8xpCKAaCyHeFtoG9fwNbTZBpQlPnvM/2hYlLwQ2fj/r
jP7Hc2wt/xH4z33VNiheqgGi/ZAtw3rFbV3Hsz762rpnR4bMQ13YT/OK6kNNyM8pyNDCUzlO/taU
xq10NpuEV9hs/bGMeUtWx9l4I9th7QN1XjXePrBFI8F2P/xrYbegoYydpVD7r3AnEi++lU783ltq
VUHRbbJknkFCjlNdfpSrdvckR9vRe9Ko6HVCfHkigHUp5kt0lMAsZzwZ0n/l3NH9l4o8U3gFypM/
jtMqbWgBEdweSz+Z2/pun8+yPXBW8mwpShZUYkGgywPlBwlwSOcaQXyT+bJrrqwXrvJpHrQhzhiW
IHlsB7AyAhFMVZGpjqeKOc18fvlk9GR6waU//8e6CbbvuVB+pFybXwWOZ8iC7ph/8sKrhtosf6Ku
U9xke7FU8bi/7fi2dPrLySl9vBD/DVah9ejm32tF5Tl3iZ3eQR9w1Pv3sESVN9g44Pb9pu26HLWf
IiYNTqJOphB5oyXBI/cThok95LV1HKqLiseZSFl/atoX43Q0wU2ZMjMv3IIByWYMPBe1qJethCTj
k6DolZaaaN6Es5S7D2DX050mq5FmykyDOxgIftTwiczTUYkfIRWG4weHXc+TsSNK9waP1U3qx5Ta
+7QnYIhIK0NBvebB3z2wo7PGpAlazC2Toyf+6IzrATpZtoy/oX/ugmUSzKjV5vF3okJYVKtqLa8K
OvHKFI4cukPtRFJ66YOb7vrHnMVPw4wMte908zP3YEp0RR3ZXk+WMXg1BkF5A+Wwa8Kl9Z6FeqFj
ljz/rndVDW4OBHxI6pD0+4342dXplOJfG0ceCRX9hw3gteNlLn889OyI8SnLTkehuTGQUx9oaAlA
ZoqhErkv8oIJerXbPA+dydEjgI8Ldsb0KjWpmQwNS1uviwDkn7laYVzQl66bfVRxrbWCpp6rOs+J
OWjvfqoHSKWYiCBDE1Htoc15b/WiMAKNFege9Rj5NeOABH89ijSjPkN3CZQ1VcUPkRgLIOWJHED7
iCpnfvwY8gunbkhk12JuO2RE7+a1dZqePjkJfaNw+qa5gL9+Vrs2xPh4e32s15QDgc5/mL0dXGrD
cd7SsUVm1+0W8sAxTJ/G4gxZFb3J359NT1dNYRcSQ+tXyd1+v64qfC1/eNqfqzB2K+yie9hvMSsP
syph2rEy0TCi1WUxGHbsFEmPaBQig4W5gJqG25Q49PfghOEg91sm4KF2X3Z1rcaqwok1hU6dPP9O
R3byZIYjY9StUxLNIxOlzBbEEXUoJcX7LXufG2VDvYmwFoVKJB0tXgTFQ+QCH3nS46aLh7lMNGar
92xgdIFoIsIpUBDK4bHml3edeTWFmsx1jjBQ/3eovGcQX9nuOiEdz5ljAkKOoV9fiBv/qU1oAnxp
4dNaPEYtXN799HCvhVkp/StOo2mI2RHQh1SY3a9z73DyodsbwSrjON4Cwd6yIgu2RGp1GJsSbPyf
nI+Sz8FlPGhu29LveaWh3C0k4IbXm4M/zCZz/iYsGxMb3YjRKepEKlqbs93rKbfJEfeMsHMf82B7
GYkZGex2DXv66CVYsdI1cXquYl6sbmcqQUstLgPHSJ9ejIfTcf6HT7KNLEY2JNwcrCshLdn61F73
SlMNZKNQKhvAJhcFx+lU/0KupzmCwrLWqdupVLnJoBmG8KOzCgI/680Fo3XDRT+aSYiKpiXEqU/l
rPOYQPeQ4dqTC1VXebqCf4hvtcGhJnzDnzL2POqSg3NesKE1wQSnhg36tJcjbgOosjG9+jzoI9Oe
K/aFnRvpGBAPX4dIrAZv2BUKfMmaQMVAmcArIXDzvgp0ALt2kkrlIFaOc2sdNyvYjHJq9J8Sx8gF
En3uVvTRQ+L5WgFKDuRKGD16Qf3eFSuhTsjklG3ukOlwaL35gGmgu/su+rvRcWtOA3h1guVY7gce
GjPpPVvyMYuMDsL4nDFPYolE1DXV4W6K8uT8Z20HUPT9gZP6b3yKDg+iJtl8d/XRefHFOYimYCbc
kWWHNzfqEQOpYeoYF5fLEkPyoBhVuJko455wWUAgoexA96tMl69qWKztAjpMOVscbWveZ3qKImhH
FGeOUyf+YK+VIIBeWrASqCgDOukyZxaPGYeoCkGsHxTj/bO7kHib7RG04s0c5rbVlrOGlCjzBNBE
X0Vjf24TWb9tZt4rr0PkqbARYcZE5YQ+PRTj9usTfOKzRywp8eyqepzE2W2150ud1Tg7A8mqwUPm
1MPEe9XKQJeExr2zjaWaEfHOBiyUZicq0WMZCn/NAy1BkFTzwx2CDENncgxqrLxGbV9mxzoCP+KZ
o2r9yUwh2SoQOACFVcUELNZ+ysBCS+tVU2LNsM0ZKgkpzOQcx2ZlhKs27J65n2u0KZK1Id2Zhxhu
F87GNTWztXSsMyiYFFM/m9eR2aRLnHFh0v5wbIjkE3hYBsFEHwzKakow0Ma0IYKhiyUewgKA6KUz
N1tZeDEUrwDwtQGzhezDWXWc6c9RcH6xKizJHgEzbxQ4idqMLNvkvS++tcMn25JGKGxjCG6CdDlZ
+HHh92B3+cgJmEpFFg1pLQndwBPL9Qj4WAfNo1gYivpjjg4n0fgr5woCs5JHt/xFuWthXjTA2Gma
e7AjZDvtf8gGZxsVUBrFUE4467ODqSWWzqc0PcYgfN4dMW2AsxbeYCxIi91K9RhLYF09ZRjBCcjy
+mqWk9V1NfovbFZBpzzF56aBXuOUMKL+Tyynk0Ee5S1RX5TupM4PjBq5iLEC6/UdFbspoig4O8Jw
x2iKRhQ9yjHb2F6svdk4NbpN4YdAA23g2d4klpMdvv39y+qIQ89T92xMmy9EhztPqi8kU30QeD2W
pXVPT5+zm65+wKdWrL76kraPnbeZj49Ep2DgZo3uAeG4jmUlq+EB3PVxyRTexSug4rOUeSamZp8n
o7dk/gPbB+CkGRVkfbUlOgLRf4oq5mqyEelIIL7BgnOAuxmw47GImMypUKx1DaQtAs+1uG+y++pB
QN++n/RZxj+jC+Fi/ovR5JBb9tHcV1jEPEiX7cokr0g3xe8ZtgbQIZYHhZ7ifEai8iMTx6tk/KE2
JdZWIPcgvl8zdJXW6L5H/Al+iA7TsXpDufC4uLjJgja1Qc3FRkyLHihdPGW0qjb+XOZoE8ZVA+C5
YwXgBLVEkDbaioJFUCHgo/n4NelFG7SHRzbjNuPLwS9/ijNSgNTz80eKAwWfo58muCS9KMBrDTs2
oJ5Yz2TisWNZ20NuqL+sxYmHu2eoVbaN9/IQSWzINZbvL4wFnGQQvR2u/CWfLZ7qbVLcF9zJJjQA
29yINKyaPZs3p5UktW5+6+SQe6sb/Xu5uDJHDFN2GVku5aElRZv59QT3t+kK9QLVgSpfTT6XS2Ml
+a9lhl5Eg7sDmwyEHRIXO0Cl5rANODNMf30fRGMoQ402KQN+pK0xbvqxuT10q5UhhL0sOTzyqbCX
XAPQLmvRMgSLZkD5nHxFIp+uoewGB5TiBTajoe2HSLNAn0/s5uLQWQTCPtXKYTf1uo650NW8rmbV
3rFIUMZEmX2DctD3M8aq20uu8OxgLEPS2bHk0nlalNfyf6hPGz834waG7KybzjgHMMgpmiBXUFrK
X49grPJkcKWuJtibkUucNI8FoUcVSiUYdN8Qtt8A7t8+FYS7FGRAQm03u+Ggpd2PhxqV1nRJzV61
YlxXwKLchDkt+IVnYokTDfG7Fj5MW9HAFAhO9PEctJNe/0vVpMcZN/qIQv4o0vOAu0oX17ii6RXo
vTzI45nJaZms4d9VkuoAEM14FcKrR1hDzkLzmI9jP55EQn2mSQ/F+vBMB+IXOXYZiFu3CAqAIvVp
bCvSPncze7DdgoDoflLe2zu77ZcUdBDXWm4pDh+8YgYq1puExwu216FEZYtIHJPppkDf7iV5ZqOM
Xv1SQ2Py4BEraVAviuEVZeMM8xzgA1KWO2shmKjUXXIgCr6W+1i5NI4DbfShRhmeSkO5oqu0ZTo4
U6hFLm8Dy6smWFYcETbntdDYVyJqq/ISO3DtZ2rQl/bPEcvCYirx/l/fFmyk2MLmmAfkMCJvz27g
zikQuCKt4okvNtYSWj1C2ufLptJyoZMI9w1u+8gSJoqTN8G5uETY0m2vBDF+vlAGiMHU2NKVrAe7
0uT2mkBBtY4oBbljmZAO4rn/DlIZs9qiBTYL17qQyckFCa/mCuvQjfknbGT89L31LylMXjfpmnoB
L0H+UxEW5LWHLQ4jR/SG2XvwrCe7H4o2UOnkh2kYJL12NqH0xkbodN+BNU4iIDn1PJd9Ldp2ycRB
BPvzQVIUWSlqouwMAIpoTLnpOtdmEC2l+8eGLWK73HNQOcK2+kUq7RBNk1tnFmgbQ7JZGzFdHTuq
mdYlgNt+BdsfBE/kWdWOdGZzlwm+DK8qS5gMpi8tuyDQIms3M2/ObWVjW7T9hjRInOk+NU5jhO3y
kFplukxQldirgF793qx6bS3oZXXkEvk+J7C8XeUQjZo0uRmj3ZVpHdZewXwuMsthF/jhqA7+a3Lk
nzV1qrM0LsRs0Gte8ebr0HojLTMWXJ73SixGnMdrlBE8Bkq8thEX+fD1yXhyyowo5lLfLtCW72KP
wsrBIokXmun/MUPRruksjcX09uw9u8esFTNZS91qkrVhFshMJht99GqTBdK9X0nRcEHQLviBxtaO
eJKKKPmgDRDTJ81MkpE3UBJtiSXr1nZ0fotmpjFEUAWVA/znMZG4lyKd6YZz/lLR/pmLqE+TyuFN
yYhyPDUXcfN8qCpklA41s6tN3Af33WjLFXTBlPbZ9AGiWcwsZoTuoS35mvOUUNlScQrDgO38QpPA
leIUqUvuqJObgws/YtfbZt561qC/YOXJy600FKBXGhvpfy82UCdV8SRrh02Ex9bK8JnqJAjGAt5u
SudrbYjbft6JUaDZwyIT+Le59ccyf8gOsTfPCA9MhgaD5MRhbMso2NrUMVSIOeJDNz7O4UlI+igL
30yFggnubVwPCtL9PVCIfBrIevYkmnWs2l0dXNyvW4hz9x6Mjd2lgmaLFmEN771x0TkLLJOPJjmy
zd4Gxrz34JpAyCu0ql4tw7qTnxucBwRX/4h9bB+hR/zQtznniOhgeniMkyyLxOKWArqDS/NsGReV
MdoYhfZrOJSepJ1y3BWxsZqypiLBUBhJ0z8R/EamLLnP87oLUj8dzTswag3bhDOHOo7RJOBf2z5k
wpEt9bqfimGEZocieKyMbQwfeceD3VAEQV0tJ00tVREfE2YW/CwGij+pdn7hQEO6GdOe/UPYluU6
33xcjufGpeZFAOgDvhzkHpVdBRIEKc46+VVu9F859b2jel2KJvU3MgVJSWAw9iRg9+NHx21Lzdwt
uOtEwBiNthdmKdZTCoCvC26GI/YuEtJXIR8ZFvxruIWmWTVH8BkcwVrESoaZlSwqtli+Zx6igyoC
jlktqSANvp795jgom1g/x0UddoovOaNOSHIX32GxO7P/1E6Czcr/SsvMCNcM3pQ2v6hkmVgHXi0H
25NfCJy2aaC8NLS0R3vyfwLnWgmtiWhtxfPXk7PbXC7tga2KMPuDr5gT0fgT6JjiYH1weqkDxKWr
Rnc7D/2OBcF7nTTkazNLtczuD+s9ymtLH0IGL2irQZXQMs22MsXEZYA4BXugiGvKbKyorkdOph9F
ErDnPWZhY8RfHKUp4bSPIv6PbtXt4LT2+EK1xsNHFl5MYlro4E8KJMZ/oDVQBc4kr6zRO7ymLPRv
YZipIjuY9u6oGAW2M3qHsMDtJfkzZhL3YAsriqfnSnbtU0Wi00xq0ZRiOL3WFqsvVm0RBdv2AIXl
SiEiFYh6vS66qFamwBrjNtfCII6BOUTFOcz/X5OxkfhsKCAs4jDmNncmzCBEaIyfGVjN9cWbHleA
2AeG+okGqjLAvWkSvoAtKabG0cvBoc4wM24X8r3ajFctU8Q/hp6+KdSBH1EFQaLx4EHAGSPt7bnb
LGfgbMGLxa7RWIcanGC8nHgGCmjhfz7tU2vK1CUNTIcCzK+lBgmaOJbM26OfwWcxuwPlylZ8kpUx
/lU/GgEbJ0FrGNKRdZE6Gs1MealYPgCXtR0S/Z7a/HM/4yfmeuamaV+4QxSdS8rNfhCsv0m0gRhZ
jqDYeVJcOjERk6TnL1ufO2PT+yQv7pj1zUlfAyWKPFIEyuZm68ERqn8F+s7a76T8rGj7T2tDcghT
OPf0jiifNhwXhFOVsRPNih9jdoYTuszJSsVLQtyLSFHetB565GC7Lg56bS7yfmzSvRv29VRQqeCP
R8tcQvmzwr+7m++ZMoj8apT7lQE4ICmZmJyBZvA4xYDAKQO0GzbGKNr7wMNfludRckBzOc+Y7oen
SPih8vEpBZXmfMtXXeP5npeEi+NcHmbh/EjKNxqB7JlX8a4sJsgxBtF1pEMLs/ZbW7qbzTyCU46C
c0qRMOLsOo+ii9Kyqp9/JuLJp//SVgtFkhBvfLilACSFbL3i1ZyhGXvErsuJewrSiNA+87zIuZyY
tPHQW3NSITuaMWGO2sDftSwBjr34QMYdmE+o7jf53p/EDVMUTBOhbEdCDaKiQyryEtnaXgd8r2eE
qGA00lLaOFh6N4hsKfjQZA67pFylBaKVgSlcioMzIqFag5hvsMwnHn/UkexRRVVlD8vnr1eha69c
w9ZQaZXgTh/gyxORuVIlJF3R7CAn+qFkkMiZJN5s9WIxzXqfYsYmcGE+yNsI7p/OAlg8ZyU8bb42
YfM9ycEqPsnElj/39xu5ztQvUMnLS6fGZmRUpfcfKjsFZ3J3cXw/Cap/T1K9Lmdngz5vLj96gYIO
5iYcg4Ss7WR1YiBQsttxSHxHzp/j5s/7kMp/s2eYJVAoTWH0dyh9FmTmy0r9ewAw+kaUgp17lr97
RxS9OrVsI/B7tcYXl1L6LePZ7tBpSuhMgyfU3Auw2KeuVVha8+kS3vMB76Vvulkt7jfCxBBT9v91
gCDFsAsSaIbLIjg702Z8XkXSWyhTu6pbth5Dbu8PjQRoic+kNonC66jduIc2NPu2SCH6n/cxXGST
k4ylfe6bRUWTDlDDkYfYAPeRBXz50ixz92CTtMvcMzTX3GuQozC78bx+adOR1ROwJYHHYAIYL1B1
ANVuKEOfVU/H039JTimaCAgvTSqucbfJrfhf7RkBpJHa9vFRqF/d8DXn9DpidIfdnNhOPp0dwnbY
dhlHRWawIq/+H3DX/T/G1V9rpvC+0Csu8260GNooRd5ST4UT+O2vbxsD4m8FESaPrTbQpNyMTAJQ
um3oIQaUtqbJ90worzsweVHvlMUiN3E0IgzwWwa3Ht6HmKg4JS0tRqyQgR4NMjRlvz3BePGWzpH9
UEwHpfP0TJ7G3j5fbhPapnSOih27Thl46YWHW0rOzfPsJLNh4/1tv3qQtBF8LfbigPca9WmB5Q8R
1yqrshgAbmFV4xGnzN2cRR6GNWkfhPMQxVLpXLJQ21FJLnLtBy/ScZJ0iqlN4IJS/wDeSWKTv6RY
j7aZ8JYPKANoAuLpX8AnqKv/BLmA3LpvEup1xki960OUWLZ4wbxb3o6HE6aw30HmEMImewbfulYu
/57vkSJZuUHiDHrswt6gVGR2QlVNIxX757++iS9ux7/CaieBNJUrQRA1W6V9dsfggduxEoeHvK01
wARLROliYdJtEcr8qOk1I/3puqX4axySzjWQs1MvUVvBuuEAozWuZiFBV74+cDYdoEXWqln3O+G2
mSTBLe/Tna75j5xL5zrfGxTYeeWrOVo6SZGnTdXHDQt4QrMA3gkg/qSjixlFnxoR8gyow/raFt+m
w2FPuTYGE/l3slkywXgpJL7onRsHAZDh5CKbV4ajPkjZzzjYJZS/uZuIlXvtORSocsPmtnVM8Obh
Saj7NlMKpe3rnoSMe/A0djHr10L1HCSk+59uC3eojvaX7qTcP9gDGOqxbrFo3Wj8h0Ti5CnG5wtW
FiGOyUipn/XNQMF0v7LEqccymd1ouksFSubh4lhnT0fYmCvnzz55dctTROcqGhF3ZjUgbhMEgYxM
23NjXLlTw6nPnaK8iBCrNYsV7FaILeH8nKQNG+dXCEnEIAwSq5BJHLYnxuZA6QtV7MrnQFSNxgvt
j4Gsj/AJXni/4VxyRuINB5sKdXIirQC55hxqxxyJPaMclXAJs4dPl1CFla1VUGGsYiO0U2u7+228
pOYkhWndeDcOBmnVSLDGMT1vg+GehoY88xtrQsajro2iKJqfp7VyY+aoFW2Ak7ceIFmfmaLQ/+EL
5IHVYv5cwRLAyumuEnSTg3mn7jC4b8c+j3NPyChqkUOTMuRSho8Z9ckPvmo/ds0AlIS+aQ6S5bpd
xko777bHpWicUIo5TsfG8NlWUgwBKfYBxF5cqCZrKUUfbjon1F+Ctgn+/kASyW52aCHOI4orA7fP
J6Pd2U4bT7nDnqKzCsuQYetsqpdZav+yTzruwdx3uhHyv2Scn/5RJRp26nSQD7/BMUHLv0IQBH9+
bc3HD9dk8UwhcUXIYcm6hQ9ilT4GYv1Cvn7hL3zhg8u0vik20qwpKk1XyQMwfcdyhsbldbLvByKK
BzMBAgbutLMR/es72QJR0N47bht3NmnRIfzqt3JnjMpwYVwzoreBMJ8YZXuJvLwzuOG/lC+3rath
Dm8m+QdViRegBB+8uNJQ/Hvsx2B6Gaio7kqfhpOow2T3agJui/ACvaLmcoMFOjPlzgaEDxTD6hOw
OjlP8J6SYhBgaWXMf13L1w6CkPlqFzCIlG48nzpMyTlW7Hi7QzD5xpBBuuO0vVscRm7Y0ZvPGIrK
5oL0Iz53chmqFE+0eHu/G7L8bkzyOjQqEw/VOY+izTWWZDd2B78FklLYo7+753ORhdP3LNk5Z782
chrnhJ7BOkHh1sBAMtq/5X79fyEMsnfY+QRpjj/9hdNXHUwBJYvZxv+dMuNkIfyvJxfX205YzPN/
GAYmW2+1fRpHnigkcQgKJyQJ63kiS7hwFn1uhhNsEEbouPDbYOux4Dyt0XTHc3SI0kbNDnujVOE+
4PZbyM5gVJMmlQCgky40XKPg/9NmAgii4I3TZDcrAoEYW+1e6lCRmX00pIVE5YC10c7+vI6aZIOt
9CAIhEe9cZEHq69MMdu2TkpXpnRya4YJDffmX1NZhwe7nTKappVS2xOrw0g94uvLUtI3K2YJ4f8X
ALnXuYiOdO3Etw4G0tahnjAactqlJcwTJSP0Is/qrDYQqkh8auc3I4lre5s9Ok/JpHHPzd1pGM1X
b5lkZJOXN5eTLnqUJDDKZxgfLgo0jpdhIdY7i1hyTd+MLaDaOz57HUFP82NeMsxFYPtcA4ci61cN
XRKcKQM2Eias3LXnnqHeRmvxBEVnGlZzzl6MkbHf78P7puY4oN/wKobVFbZmEpGH/znn8irtukpD
8K2RJHe2O5aQpof4EyHTHRURdHQ6Wbki/JyoI8LlfiQMY/v9IZXYLX6edME1RlPbQTQ2ilY6bhrY
X3rAbP5U294I/goN8a5abGcrHYcSdUyDS9Pf92neLHloqsCY7rnha5XT4LkkMRwztBy9tD0nKAKO
F3MLVcbuGqGT6kC/4b+1JXpRFf7iIz9NtRE0pq+auT+Lbw3C0kIWS+v9AtTaua9/In49bX/kPrDX
bGT65PpYMyUrdmorFhmeKe7CEvUeLikyeAs1q4eEpjs13T28UDC7YBRLqZlXUhpy1Kkye5TdAygw
rV3yK3AF6BFr/RgHgeCIfcvpfcxMGnQgRkYlssDNkjAtAjXPyzwQdEZR6oOyxwhlZwc3C1/zH4C1
Vfrh4e6/LFgcyk8VxbnUb4rV6Xr9FyeRMUcwqLryf/wMz/kTejrw6B/mL5nfmHMWM6VTlCfb0ASJ
d017rb7JPXieIUqVYR+P3z/GgIAY/UZVaJQDXQ+LciiNqEnl82yBYQUbhP6iWMltM7RScSYzLyph
d3VDUnnZBL+8Ay3HZkzT8/jCs8HoMiflnKjXYK0QqUMX4+jCgQp6ZB3Jn/dF0dbrwtngTUdF040R
jIpdoqpbAUanPdmRRcWenvDsfMIDeNGPk/diTJLFnUfJc9ok+2yvq163JonZIWqDyZbIEDFrZ8HB
CtQOPCwiC7pL1fOIS/HhDLvxdNpvDIfF8f0P5mY39/GQxVpFP5W19wh4DlcqcToJCodSbuqNYxr4
pTfOgGzn1NHqKD9YV9J3yjyzrNSCQeU03PLrKNjw2kwM6zayjAudAyv8lo4mZ/tY1p1CvVaRB/qH
1umrIabDt10Jfx9hurb4av6tIu2qzLUweAPNlhVrbXDwiwOr1JEvTiPiXsJTFYYka/DmhLv0caeN
fM8RpjfWeaYVPQlhWh4v1sF+qJX3tulSQh8Ezh6zYFEG/FEJJknWArbI+31k9eTkQNVMuwENl977
BHMBC+uOdXtJ2qPsZEMxhjn+IqpWCN+42FDar+IvK8YYAPgzW13x62MXC0FY3L1djUDTdSwxnZqN
QFPkm5z7O7BHepHh8lUoynd+7n5jqzZmFjC4cHPDO2My6IiyDwKor5qklGmL82TcTZssnsaeLgiW
ZyiNaR8y6+XiAFmWsqXhfhNYyoyceLMHDFZTajUyEPPMIB+nkRIoV55AQ9A2PPMPbVbZyNF9GNJe
KXA7I0LvxgpSFtNkf/yA5Or7zGYTDWr5QSPjPDhMmuj3HIVhZOVHV0LkhSJmKoeiQbD+YQ8uzgw0
y//KUBGe1r/5AVjxQzYI6KjM8edlDBKtiVi6gVy8ve8M4a4+9sEvNpvjsVRfp7h3GaSyqLwC8yUV
X9V+SxXEUo3WL3r+4pjyAsB/XRW4Qsq0cU5e0WxaVochTKJjoz9AmKF4mG44vogFqogGL9XIq3oK
eINbwAXROrYreoVLKhISn/FjomFOPf+caVlgpeo1+npo6lwCR5VUWG7WcTSN+E4nwsufcUShwPmZ
0SfVyKiXD01rj+XrC/FNJ5wfl1D2yQ+jGFh0wokdq0qQGxlUwNarEQON8YiD3OuGmPnweBZIPlI8
s6FxMbT1rXo6hZTP6qXVDll/9WJZekA2lHHtU6QfLiC2qCoD0tAiqv4BtYv7/kDu9hB0dyllTxSC
Lq4kxcJkcoAeNg6Lfhp9n1nJYW+3aD3LSeDEXKk9l2qBCcg3JhyKEAdOYXlj16stxeNBE4zPgXvP
steEXi7kuOFwNsE6cw5QkvPjpHQRfRCBzPyNmyRVQda9iFS5+QZDK3FcluYZYB5n5AWx0Xp76aXv
g/eTEiQhNu+NOWx+ChwW7lpoBUvz70XIh1F2J1O+oR72468GYD85zVZgyXHgBxy+lg73cUtfywJm
SureOoB7JR4uxYftkSyk+v+n65QnXAekPcgxBeRhOGU/XFVCRKrysS9ULOS1+vPb+YoGKaYq8AbW
G93wztgzrP7QIxhFSiNF3unsUVn1/LSur3Jpvs+EllF99tjFP2x1s0J/OFGzDR417jjWUemryH6j
RU3H34UE3CtGnEOjXFGA5ZhQRtGNxIws40KcWQ+nIDHXlHYnBlmFSkfKwU3/smHKvuybDe+u0kuZ
jReowUJHuE37sBDpQwwQjvKNqoVRfICgcQtKK/eUeHAmyTM7pPVGfRVwxiYdQvy2YRDSVBN1+XEj
T/Di75SYWr3M9WzbMPFtyyLQ5nVMLEfI/BovfOcKz3KD4nByli6gaPXfb1uElnP7MKv5yYyAganE
dI2qu8nhNNuNOBmxft6AgZZBRmkeG0/eeVIHtf9owf/jBxgnXYJyvc6yz/1N4qIg3690r2jDiW1x
49pHbkndT1VvZ6Tzd60NUwFEAZgGsbG6sz6aL3FhcNU9zyve2s3YjLXTYlls9nKDQnRfIDhSfLBI
cHKBFgQ2MoHlNLMadzlgMF75RUUiW3m6XhI5cBzI9wPcfekF6bggPNS6eTpKSyssQ4jWsE6It/DD
aXqoi4LFUEt9wfE2Zk7wz3luMvIqj2hjCWd4XuMNn9+YgwN7mkd8cGZ5hdfaUcGHgSiPEYPSssR4
Fu8emkCQsbuQB0uj5O2QpUCFT/G5YrVT1fFFUHPuRukrY8L/+RiR8mTii4AzvaCzAhER/vJ9pT99
f+5BF9D2Lri9lljxnkgide0EvHvYJKqF909RFpkX58+8YkqpQ0IBb/3k2zcHzDCS4aHfMJe5ityX
HIglw2c0vSmhXaya6/jXVtgnvxh53o1zddbPoxbHt5DFjfsXJ3QCeI/F9GoaIaubyh5PcTnsqZ66
6HKmQm6NtZVrNH01rZrZuBdkWm1vIKpvhhx2pH7se4LFKuxUp8AFd2L2p/xwugZ4SM37kErGTP3F
kqsmaapcEB3QiMoo1e8hVnSb6QXzPQhvTCVAqdIZNv3nwodJZwPQM3PFMVrw8XtyANW2X1jvNAga
fYs0kud0sygtGqS7MTOUc6/SPlnLpxBELIA7VUfvmmDibGG2WO4OHJKVjac4fMS90kh391O+EJHX
7Tk279wvnLE1+CPMgvKsrN3dUuaWV0UhyAVEc4AzltlZaj6CVrRS/cQZpw+tHHVqPAu+ctus0jeq
8rkKkallaTEcLl751/enB/5tAic9cIHYa9iecWm3c4yE+uCdLWMvPtkqQmGVE1PMVIjNVAt0xyVd
VaGCVKH2VOWcAfExOA4sK/F2ZFTSOSVHqCl1tQAGKK/tU83KWuhFNTYzNXLoFuiD8V4iTBU7axDV
+lFNhbx1ketp88173ChlQ94hZ89EM09oIOtNxm05gyc3pcwd8IfaKrnakT2X8nZjFeNyRCQd91+O
Pprti9Y921MaCfsG2Xm+8dy+IoTuLoCVhWKePwYzyf/6temLQMFhg+ZWVxjIX9MAK/p/T9j8kW38
4UajRtCdbV5qcsbuDw23+nYn8EYP2gAes3EL7ynsn5bN9nOo0HEoyfzxO76dUw3xRQQDypQ+3APd
qVyWC9Mi4Yu8p6Py22yQaF6hQUtshDiYJAxtr3K8olQ/SLIiVYBRDBeIW8HwTXDx86ICfgB120qO
ou1mTdxfemFT8s14ENAs3lJRlwRztC3YEjma638xvMu3lCVPpAUFeBKbJBsfG0iNlTRc+13mbvU1
LOB1GUqwsvfsVykd3dfwC3myAcRFO6A13lDukdJY9xvemmhrnFKRKWgsDxfJBnDXRXB1S79ChCIn
pcNQtDLdYs+HxmYpFZVitojkpWBv/rVl15bu4VZnm3Pd/RDqcNnjLRnu1Zw0ZSn570707/JkyHpp
4W+qlXIKiSV8Qm6pNweIEG24j3RdkktnGGj2qw98klE+oe/SOCFtMosPbmuuHVw4n5eZN9muoFxN
kvelsSxYYPFekA2Ifp83pjGGQdrZ4faT5tpLGk20uu1YT5FbAMacGg5QaF5DCqkN1RAL7yqPkBpD
HzjMu0kJ90rBQyoJq+Av6NJlBX5ViW6iFDJdJSkO0wZloOc+HKIG1uPtYXr6LIALNy/w4RQNMHHF
N4PhJpkqIHOwz+9LyQh1n5VBBr6hXbQpp8DQsbLgZfhHBJG6VTfIFUOy5mqSj3I/X413xg03FEtK
J+VfKEbFQnWhB/nejOs+7+lD3x5LMGnz/VqkzPy9PPk4PLZswqj6ThgQ0VkoQGNyLaCFPVFG5pR6
POUbnPIIoe+SKsrA7yCJjS6vp3MVAgrv8QTVrC7nOFq7PRGPgJFI0E71Wc2Rj1B8v+BtprUvIZnr
6cOKed//vu/pL4TquMrAYmZD4HRF7rnldA5/sq91Y6RveYiQJrGikXw6Q9vD8S7tH8G37x7HQysS
q/DSv7rJKVg8Mzx7aQ4ad1kpY5tCqMqWely/Fjgd6sY5FfNBLbw0PIE8Bclq0EBQPCFjxdUkkWmZ
3OMIjKCovpxXaiplsO7RDtGLGxF1FNRtrorHQyfFeIQa4Oo7KkzbpbOblPMqD9nqk36ElwsaawO6
UsU/bO8ffucMMBGwNY0nu2nyXB8BfysoS05Cvtm+LEfHWdlYmZOfVikfUip9rY4LUzsSI7hTPF+E
bdoJaOBjSF/5lqz1X3IgTmKL8poQOSFsIiQQDe+lV1RL9+Ta5mTDgsUjKGXQQAmwqFMOhpUD7F0b
TDQgYK8HieFsxUm0c4bcCHrM8YB3K80Tk27mj0/vkSLKXJpoxKpWN+xl57TmBlYELN+vvMc5umqQ
KyXTHKEteW85wrE7FsCgA+BAYf5xD5sRqyMKA0b3tF//pTx6yLocWZEcq4OYhXqZis5+8+RbCqNh
eI1lihhnLcm0FYBR1Q9jwJaXr6P1PK+w40mFuKWg/Dh9HGj1uKc4mCje5UuqCdbu2dgSCpduJ61c
Wou41y2bd65lSRhw/RiyB4/xGZ6n1bmOe2tEjotNCTTJ5oYdimNdn1dzQtEgAjOpfxkqBn8/Ffdk
xhqAQUVwflF5mis7dT6Ru9U5eQzEF624Kugkp6FfgyPu0TKE3E3UPvejDoGbfF/ofBKJMD+czwZE
8LZuM2X2XhportrqTL+09v3VD4izJrlhyNcNrvJiaceekLbMDU1Ho+sfql3TExZflKiLQ/PeEj0w
FvdegK+abvdwfUF2HMQaf+CvnTWRtF5A2SArA1YnT6dOQonYZG+ZMUfNi4hYr36xIK1NB4tlJv8t
lSe7BgTLowrdon4NDalvrguxEAqHt6mNlfY9XkCkjk4W8jfv/wKHOoqse4EsGcnm9erUGezc8W1t
ncvZ1xZmO9CXdVz/9K0MMtdOxPib1DsKulnhD/zFJAPY0zKFqE1qseoGzQvEcwOc+ZqAo4/ApGYN
XOXpCa/V4V/yjsvpitYHbKO65ou0t71aUA2iCr2tDwcuQ0mXotCJOlYDFQpU6TnONYu683863mYu
lQM9pi1nqxHz4mGb39MAzYFYSHrfiyeroHVKhrAkBMI+h89UVEzj+k0qFgWueAcQGcoKF4iHY8n7
vI4AzyGEdS/Vgh6MkhOG75eWl5IAI1B8Q7VZnbOTUpabFVT3TKTPUncS7DdqnVxPHPqJexRZFWrP
1rM/nyARwaR0HUlzUMhsdtFlxvdlc3H1lwvZuZ2l/Nf0vok32OoJpLKNoRgxXiTQ0l71MzPSE2JJ
ythSCyNe1bDRd0WdqkrmXavRYH+K4akOIji5DTI4Oxw9oo5xXDkMITH0BG4cduapd8EPlJjOyvgE
XdSjQ2j13WMQIV1VP+tSAUyBfkKpkM4VUmB8Hi0XS3E9OifxkqoAHmHoHb4Ksobc2t6EKVeikM6Q
2zr7BwlzymUOqvtf4vrDeWh8z4SXYKviLGwNX5vNAz8NTIaHEL4azGwk5Q0intGeTZG0DY8ZjsQA
8wY4FzbYRh54And7mVrLAo5gmpWSocLSULra/DI746rLbYN2OvnO90d8bYQFMZRb9KcqISo3S1su
s3gYM+igfowJy8Zfl05VPx9b+ZvJhkRijqfpmqcpgWS/YjDfP+YSA72jyneMH1pXbBlA49wtrK/f
OCBMd36HUgr7MxNF1VoAFmmTWD+J3SlVwGPzt8NAHNUkFr+jtGRD4A5HH2CKnDG0V0GofFw6W5zs
VKPoDkBpXXvLp/APW0xp6xP4OIKc7FOzSWVxTw0cTb+VR7uZMMdWtL92QCCB62lgtkBG6/I2d8HC
AUYvYPA24HkiTmTVU8bFrssmkbochEHZXClRqoB2a9/NnSUWltmGttAR6BY0LBA/kT9uAfYGkr28
0TnoRHrZxGAfl721zAJNWl/WZvakF8cnvGdt9j3nDLa8MKWM/FhUEzt+YjOhf/yodFryMZx8y1ek
VCexnF0ze6kOFA/wgGlUiVWt/FuPMX3jBTekn+snjVIhUPCbbeyGwb7rQy+ERFCnu8h/zc/v8Tur
3au8msKboX2pmfpkfW4eu5CqU0X45c5o6Ga/J10elccKBBkzS8GsZogiosvqgNUQTz/EzDaZQNJK
WX+2VvgWDd5FKNdurNpnJUgikENyCbECJJdkJDV3MKRcg1RStX/Zjm3k55rizYAc4GR1q+WEyCly
bPrYaMcPieNdVJHHpj67CiyB7bJVAmuafzh6b9r3TJLz5sEtWQyjjwlI4gEobqVVYCXiqPb4v+v+
qeQF2wXz1QI4JtOXz6CtZAnjL2WLbf8xd4C5WexynbOQw04T4+R4cBAqJ3AudefNiNwqDUZCpxgz
zMcuwknIYM1eCZwKsTwE+CYtFuPJYHfAkpcq4/WESnjZFWS4OY2PcGZKj4AalDVWBScCNziKBBsv
jq3WZdl4wOtuOb/dLlkW2ehyZeLmqKJRYoiiFFyJGQeweE+QUFqZtjSVcb3QG6VHrVAxOjQeFwgK
lmG4ONlChhbxLzo2IPLF4KKWTFbWGKUr7bDutKhD6JExSs7Sown7QmIe8HMh8yNt/W6lezrXp1iV
t0a9IC9eYxuYhcu1YFV7z/oVlJb8hBghOziyGG8D7CtbA84qwGH/8NULsPm+rb1Buz8THaND0Dph
x/twVjO7+j+oOFY6A74vhPu5C8Px4opQHhJKomiK2nvOhzwRrH5WxT1jBe3dARmx14ytYLfxf/cE
doso+EybEUpl4ygS21+gRu9+Prbn2Cpc4K3lCg7LanP48It0GWZnGmtKKBz3KEiwgHWstw8gY/qd
h6Vy/f/V+L8MyH8ZYCUPCYx1hWMtlsQRHcgb5AD6qQYiJCqj5u3ZCi1EweO6NlBMDRKF2X/eNu3J
XTcNpMiXEo4PeaxG0x80ByvyQ8OMb2Uf9KRXDU2hv4BMFv5+9jfbJgzFZBGOYG8yLi1LE22mYHQf
keNH2pWQ3VWAR8NSLmsQsYrdq87iD+3qthVZVkssdM+nJQc6hKBdsYtsa6hweA9m7MY2j0vBiX0V
l8Z9k7yH6nJPTDpS/G1pEQ1/ARSji/R6IfApUqAzsPOHzFwgm7m4orqkuuAGvi7i/yExkGhmmxNr
Z3R1noTkTMg/Mz2OuVzBPXT2yrM3ulN9tD1U3ysiFC8hSJhl60rIFQMS74Jzag7SvytFAfNS7jLn
oCecT7e421rgL2v5E5K9PRIYlgC1x2eY+RIiJ7vp4Efv5nxpJTLAqhOHCOLOUWttVZqyUYijDytI
1I5Bh8CsZ4bOxiA4ye6G3LYFlqBhVY6DEB3i/q8BLaMjx+2XGhYUhaOi5sq8zANs5EMFT5AoE6Ho
+1tskPx0iCBj/51ZJsfKmQw6sEYc9343w8nrobcwVzFWYV4kCSk0CpdQBMbXvrZbAV9bhcw5la7n
4oikSD31cxJpQx7L+hW8loQPS65TtUhNYwqwSPpdUwY6++8hx6fNAgACa2l+zYVPJJ7OB6Aq3aH9
uoQbPaVgfzzYOp8Fw0UB2W70gaQk0P31qOFgUCO39rV2kReYZZs3nGk8i0mseyTuBr0sHQ7bEyln
ujnjqiI9RPEOTvcDqlaOp2FiCcSnhW3XSkGZ9Rodj48pWsHjDIgeQv/stNRNTxY1vsX+1CfAW7Rw
xt7ynypHtaB/RTKiOVv+RgXLvD6UYHtxwL3BmuPJAQSkMY8ZJaw6TOLZtYx9rAEETZd+tCxxRCB4
cH6Qgk4FWfinx46lfyUejz4oeery4FsyTM7ER2x8TnNZNbID4GuNrSvTJMQ+JBmMJyTmtPM02JB/
t1KDXqgh7LT2fYGftr40RWR4FE0+M9nJFCqqIOZRBTQgHFQA9pl+GNeTRB40sBFyg1r+CgDJHPlM
frReiOmJmjgsp9blQxsgyHsxpJjvkVqd7HmkjEB0p9tk6XCskbIyM8QlWmNkKjdESMDd/4SvwpwH
hXXwXiHiwliGcSDTRGcphX09mFJMMRvyphM9+lkBP+YgO4fMpy2gC7yKbNS70Ew6P9OWqUY3B3/M
pOyVbXX9BDjZZNWn36TQo7shG0W/4648Gwgu77fi2z70RBDv7yTPPatz5JfuSiqUR/S2adseROez
wMw1ym4CzKGbGwfjeoXP99fV8dpR1F8/kbLDDlYGxvj+9L+twWxb0xwlrqcydexg4TlDxdLMnrp/
AlOqk0qFEDMH57u6pdtQLYphw059bNeIzaALlzz0RpYftvpfO5zaDvlu4MzqhenjtCyS0A9bJyX4
5n8b/puEh1nKUZWydRPp8Rs7vYgApFFfcp209Nvi40A0NLnkpjbFji5js8fP3Y304jWE+MQnRhSN
Jn0c4fTPbvNhAzDhlK5jmZuBO8QVcY0AAckp7hbP0Tz1t7hdfIFDNfGGS2lyNeeYC3ttZbxGk5Jz
BKYNgHd115UDcuG5n0rEho9ecgGKWorz+UDl9AkDzTMdQxHnQem3L4BtDq/jf5IyL9tjFx2Jnk4p
f1y0Jt7Y4slmXWlSX90x02aoZWqT1KtyrVHVHpnwck12faZ5Kihz9XQyw+G1catcGIQ3y/APJ4PT
KpX1ipsf/vus8ROnT2HJLxTFWCPO1wfbxBEOvWb2Ucl1vDhIm1wJid8n17ZroBBdl4PHp85RmFn/
ELViKVBz7GIbf7pVSQ5u/s62BySpb/FDWPCkazFO8b9AeBiypz4b6UuxII9aUBVH5uAxcMwfOsMi
k+n+7QQYjO0sQ7tAF/kPgkR9npRmNjQhj2gG7hcgLhOug+XusptPGO20nWae9j7+KKWG3lV2mz8f
dRwxhFDvLiqtV+MLhBZasCG+jwIgLNkthCdhEMTXxicqwzUdloGaFhNDvxDY+QFzSHy4udAWUd2v
m3YVsrQ1ipbGdmOV4iw5ghIZFOPL+kzjAQsh7tRxHqiuRfjgdXhTFonmy6pHwvG1FvENJHZr0/52
HG06oX9RTKW2A2vK163K0o9ABf8kWNIb6GvjkJB0fhbBOojUxv87XP2G4drgV6EPncXxuRJ3LDEU
ZB0I1S7V8W5usL6FqHptND5xqB87at0u4kyf/KsFm22IbSwHetPQlEjydvS7onFQFN/m/VcCaqpY
npmVfFU1KNx5pJMoE9HPSXlm2FIPGq9ve0bqQo1FMuoY6vp8N2bw0vJljK5EEwRAITk8XiB6EMdR
EBceAcPSy9TvpJ8ASCoFl8ZN95EhwhFW5fnfbenlh8I7hzm90V4q3CoJKAr8CGuGo499bUeWqke6
3SfB4gB9GLQJN05yC/OcbnsxUg4fSJEU966305km2PpxICek4RBPKwpZp6+0MASb/ZzjPQv4WA18
maCl+uEb6ix7Swd9sdDHzpE4yhhpdywwJGQu6VgryArr0umlNtGaW4pk/PgxpvcMioiQme3SxSaO
XVHKILAe835Orxufi09a1RTWvG51GuilTpxz748GHjp+fCVqnIHI2ZMgwB3J9/qgXGVuxtUIJkEr
QGRj9E3PnHgPQSv497kDOCdJofObIYiX7hF96OIsqALXOp8VnWhWO8NLhMSa5opXWlhHo6TQfu6c
lSLB7C6J12MqCoSSTLJoPHx1h39rWcpnebz4YYbG4jD9od7zG9C7gPK3Q1Svz/DIRdx7G4OIJ8gV
pNCbhmTGxxTotAo3wqmq49Z1QY6Eozz21f8yt3pdj3beTFoZdsSAPMFdKJ706si1EMRblu+5qtVg
MjIPjxGLClLj4uYV1a3vJ6ov6BZdxUmCVMakOJq+hY/l5KSIvGfU2UM9Y9SdFo+PcPDqE5oZrMon
/9vFIQslUVa7BpUUt09E4521XwaR5BMA7zpDQ7Y/FlmIuK+pQe86LiGmrYyF1TZxeniAffvw0TCq
++WURRuz3qRBlH7X2kNlE1yBsZx1jshXwv4+ehNRFFO81DEZqL8+Dq8rMbLBxL+Tn9sjP6fjXSIv
0D8yLFwUoOSi9IUrqkXGmU7S9tr2f/Wln0ftjqcu9cNJx80lCr39G6/psHXi7YJEMj7u+bFLA3TC
BSxIEMi/NCWGVUqjSVl71gPO+QxCRP8M3I1bMpxyMrdzOmqZrxqSb1sHLgAtt1POpuhyxFCoyuYw
GJ2GHSH3FlgCrxz1EhZwTevnKapWzj40o86dWpgVTsSRmNgVulHnVN96g1eXl2GTTGO8CLDAFEtk
i6UxJKI+fl/hZW1nrWa7e8OT+4WXRF/u5113aW/X+tAdtNG5OCYui6TGMEAL6E0lJiUFnm5dL9gd
wVZvE9MOPsAlk9zW6ureCmC5cXjuAH4Qq2fpO7se0HMhPYjzkkkD5tSzU/SPpn8LsGZ6bD3AUGnH
OKr9/j/FszOhrjvXEokffUhQRT32Nhak+YNemzJZif7KBwUiEunIMpuyxRnDq3oKWMDXAk/jaq1h
lr/vhOU+/F3gH79evYjbbi9bgU9M/XEdncnIugsJheGiRBF7J8PKkvLPHyPoXT22WgPbLiPIYG/X
TA5Fhm5YS0zLEK7+/riA3rnJPc/3Il6KaSOk5RcDNkY6urp6HFfz5t9H7XJ9Heg3RZ3PeBq7WTfU
R5YxVXj8h6d5LTybCUCX6XR5gAbwV632eZUfrevbZRpFA2AyAVxockHM8Nx37Rj1ekYIB5U84Tof
9+E2RNPcON3qtbS7yC/wFzasY5YC5TDY6vKscbPkPDFfKW5+20kf4wBS5wl1SnGYufWbgBgcw2aF
8hvPdkSNUcgfhoDbqsbDXG3YdkSdvCuYNzBMRljyOdvpUArV/rJwsZYepl19arLHLzBG5+eGco8w
GA2vayU3GjvvZhoo5pZTVPXGD0lqrt/bzrLfTsgavfAEjziepZPnzrCzb+uMXN2KuRwBVw15cIA0
nOw7VAYdCPru/2Nsze30Q5/3MXv5dQ85y5Qkh7QHfTyzEzJoMn/f75F0Rki/+tPqr9D6U1j4Odoh
DtIvj9cpqsTStXbAR1Nz+OJR6trN58za2jkf4PBuM2sGp4awUxCZMk4d94vv27TqAX2QyvdVh2Ow
682UJeg8nJexdpIOwd0DoW2p35MlbX+lIbaznZYypL0Cw5C9dXCUrkyFqcR6fdcqK5/2bsGOp0HA
0SWjOhK37t8UCm+C02L8pBPZiVCP0/98bRSPrgIUE93MxsdTSratUYbxj3lwIurcsFoMV8vuW1nF
vlp1iKwRwiKAWtbZ9owjLvRiyFX0PuzbCHfq27FsEOGdytbldzPWcZ6aKO1LBXzYxDOt0u6dtsUi
IhxKdaZfQzU4vPP2GAzj/Kh2UbFK2+u2XhONDQnb7v1AGmYxkJW26pzAjtp6QomsLm9I60dniF+p
IskBnpQO5yR5KMaJoBpIoXs00wPqkt7mtU4j63669F/uf9TonEEWANCBk8gLMFScAWw2xaInaQKQ
qKCjAz2qgq0FR6brHn6B0sd+9CEP0Z6E4qEQsVx2Osu/KcHZ2skCOb3cRKbwNq+MS1EA4diotUj8
9KiRYtj3eAR5DuCRKpcMHLjJZtXKUXrMesqFWG4PNzPtgOfq7oOCSKv3SKrMpUodgfcz23nYgDsm
S3S4dXxD/Tl4RoJhHoEsy38D+VQ6nQnLaSFczJvRye3Kj6FYouPri0iw6IM25oq6lGQSpUMmxRlx
BAOH1En/3FRogEu0ykcYLFGPz49hjDEtmpammYx5jfLvKzXNEK1CM43lFUAssH562uV6w88rQ6QI
uyTxuhLsZR4z3qOt9HdrqWpNzdcotXQpXWBxR21dcVTwNpk8qeN6Y+NuJ8dFUOf/CUtfJ5AALPzG
oG0izEog5Q54U78a+6vmVEfR74x0EYo6fmBWnuhuZcHWGslZcG3PG1CLtZJ7r0HAdYQ0MNiiEUrD
mLBFqYhyLzQuca8eK0SLycu1SAk0RNUsdySs06mUMVJEBtmV2fT7OYxmpOIZCBb+xjJKtyxOhmjR
LouIDz4OO0yxiRyMkT1rrZptKMt+xBKzXZki3f+tz9P6X46CLMDgL6CVED5hA7h3hFa3gl7LMLEl
hjwXHMxeD6hhWHIbTeSUI6QkHMHSHaZU+i0nrMlKjiyKbU3r/6FX8nBoYDC4MO9zzmhPhYR9pVhc
XDd7XtUG3zchA3R4CNuuPju5ptzj5iFCAp0QgF9tGjS0/Gbij1iRIvueTFWrz7gbi+HNY/3zDOzw
CqdhhH8qLT2RdvytJYVooUrV/nU4kXmElxcQToPO0eKfrC80vqufKwWHRthUDfr/mhm328vG5uvO
mdpW6C+FpHWkOSY+Ft2i28h19F7fhqv5lfQZcDUa987WfHD6wYdqBqQx/VSyRZgLqi734mfcG7ry
9mnioL2g/Zc4GHsCoevIgo3GQdHTmlobmdsDik9qLyjK+X6wTUJrHpR/Fb0Wn2+RN6Ra82DRCt12
vgE99yZUgZz0VA+R0n41ySdeUhYQkWyPHPrGBHqrLMlNfwBmTFuNKlXQX4/MJLqr0B4aN6IxEeyH
0atkXV7qz9T5ijS+IoCURXbrtM2BKGZx3zech6SqTufrUYFCTlmLBK4Dr5mlCiNPXnXTPoEL53uw
tJ+T+x/83SRqdkwAQ6URZEJEutIe5u01p9FzpGE49HO8nIv9U8Dxw2o17ZHQ/86ObsKy5M3QS4ZB
gRVlZ3lT114Q47Hb8CVx9zsFa9RmWGEvxISgkxker/NjMjEi/52+w8CIc5glFQ2mzdsK+WT1kLtS
uEzo0aO/JiIpb9T1C4SSNbOz2eejmCzWmZGRPHFppdsyk3HdR3nOD1YfJvLQUOpkQQ3iCRuW3mdl
kkY5RCXufD02ECqD4qwmn1eDC1fSL9/OSzcGqFeLUmzYjyM5hJYFqH6/z4LSa1RzlsW9Ezr1Zpjg
hxmgNkzst7DQaXJQiSdMkRUvSy2OJ2Z0nbnPDOGpge8K5apNcuVwShSPNbTFdyOF/W0/5Igz21Tm
YevUncO1WqyRXjhkgrVG+C4qCyuawqMzzBS8T10g4URKpFnB17sp324Hy+uiSyido610nuKfOC3v
sK88OEC8Oa9ASSQ8jm+ad/JXSkYNE7YkUOzwnuuYYPrSmUtXW3A/XOg0EVf0wAS1v93pkljWbjt5
mO1PK0CkC3z4OnUqOcgdbKOUdYB1cBFJ+3/g7ztENtU+0jLgeA1zB6YfwqVhqTkTQ1RE4Rm/qnv0
eo+69906qnak3dW9aH+ujAzMSeBPi27Akv/xr4bgTIw/BlFd9dyLQHQuaFBra3+cBSJkYTRMVBiZ
OwD2fGhjT+KlZajjz/XXz9AVsuxeMo821klNn4sUx4nQTzMBNCGuXIilfR4x/r/Bzp8Xk08ZtzwJ
vQW1M/VgBgydrN8JILvWIrkcSbVZHO43X9qY/KTMHzCBuvh3jhD3+H7WMb55sHHKg2dd2b4AP20k
5hRlvlU4IQeJMeH6y8xVAXjmBFbvThAXJSyRiYuoNqs3o7hmn1FvTCmHrYrtChEkNP5AaYrcI1Rz
VF8FUGJEfLs/7lCioTlC+f/jwGTYX8adcR+/1IfrNTtid6tbtp5wD0dZKtDTfgOo/eA2+N76rAVc
MjkIy17qCWFcxkQA4VvtPPMCF9KtAM72OeGGhlM+6W3/4IoSJdB5JWSB0taY7d7uyTtehkaetmC+
SiNG2bYFNaG8MhPB5JXOHAJy2DgdFw7Tpp1gHJY+69r3SviTQzKNz19uVfl0P+zpF7aujapGoTay
nFbPUFGbSfTDO3cjHu3AdJvqz34JA+OARWw8YCT6NYXhL+cSYdj9sZhogeOSWzu9RtYnv9oin7TL
9+Dai8p4Pe6gTcxb1FrRs27gqf5kSi8c9tjpUtesLScsFEhdvGonTd1bUSj4IrQykQ5CaJKpMIwz
ETstpAS8MaROEBUCS+W6Dpx35m2YCrqZ3Vvf42q54Lv5NDKzqQ/UCwehQmTws/4ZnHyv+1mfDY6S
4OHs6vbhtNvV0+U3a9bCOpxZg5k2wS9pc5vvz0DiDGVo0NGy8ZmSvZKz4D6is40+DgCHkI5ZmCFy
en8XCjOGetH+Qz7FIXixisndiq5jhbxgrRDoJaOcXhctzE9aX4EbxALQRGoHG0+KMrlS1DZrg/Sn
wVcZMmo5O3VnXILIOdareAQ99HmbVLTDPShwGMHPKHj4ngsE2etbB1FQy+9RtRQuXeSLzLitnnhl
FyEbxAL8of531jWKwn3U0l3oCTyYTMjjUGkbn2ipUtxCCnPGD24qLdYofFNcmJflFy4uezzaAHQs
tVdoASv+BddqEa5WG9fN4AFP3Gg0Zqr2VJ0fRMXSleDN3tYGqVUEIp7eGqFdaoNuWamtrc76shUb
L2rMxnXQyCEQJoBvFJ46vN5k13gUzrYiESB8EpSyoNKKlDCawcia2EejR3HKVZovDPW68RC7mvyc
/O9Mi5cQs/6EVQigRHvHwxhmj/FsMf+YnsYQNNdYidzIOrUdawLpgWaXf1hHG79bkdjEBPABuwVn
elLdlygryzEGA6KKjsMfmJgqp3XeIlgeRPg4QyZauyPOEFbSiPFg8D/sgqTAkl5hsW7tsMRYKx8p
9WpnOLHCtXNOn0ogO98MT96Qaiw19Eff71QGoxsXF/qtjD15kIpYx4vhZqfA3T7/uGHktwP6j0Ba
W87eeXWqOM1x69LTPmbumCbrC975bQZfJ6VTweouitW0sPf6qD1xA5Vk1l2C1zdTbTFzQYqWAE2y
zYI80ekRtF8ApTV6oWYxZ2MYlsiU5F5b9RMEIgXQ2O2M02+FADnDOsbn0QLpwG9YNG3pB5k8aYSi
XnKoUfkyDjgV1RDcIT2+kNIBH7Cohgn7sGQ/Gx6UyvnVX1CWtWC4WBbRRZY1/wvZaW88+qxZo60i
6qvYXsL7VjCW6PBAwJWfFNYtaQIx6gBE94X2UJSO1YkNVrBpKFlfnJokMKiXS2ZfnoEZN30exujd
1UHETu2l+H1zDtUSaQc0dPfnrvbrOyawJjNFC0sF5qY6jr2znZsSh2VX3ERjG3WMoy2lTn0eYB9G
/be73ArMufv8xpFOz2ODQCOrDVNF+AafN/Rc/N0BbXL2rMSwVNgId4Po5s6R1TovTmlZu2lP+4dr
ykOJAyHqUa9ac4RuJn7c14Cb9GYfUMBImkvI8e01Olazlp8Oc4eVlSzpXOVFRgqfYLLmLltLw+Z5
EFRbuB07hVZvaCzfppmSo1Djinf+U8px5E6FrHCA1sgyx2aRjKNVBimbR0354O3VtjiLU+IBf2uT
vL8o4snKOsByeoRLuQDrQ5QqwTqXwWcEzhQd8watrs79pL7ACtOiiA6DhUZ/4kObULCdGdOdPvI2
/iGBCq20tJNAs2h4jBkIxVQHg0ZqbRaVreJAn9krg8zjsxygioaY1/Rmp8C8T51YZYz2k0n6z7eJ
gjBHHCPqjsQrT0vnAQzkOOGrxOkZg++8cVPcbexQQGI9W99Mj2RLjqTnZD4rdTGwMHhfibNqWEmt
JH8eD9GCBlvQFv/ph7TT8gJMuLBmjx0kzF3svd/qkmlP4Kc6PVaSSBjBpiAtlH52CVMyDxNKqyF2
24FeRGo6VK2+fT6axE1Ql5G94GEK8VUH/H5B/iW+oIt+sOiloQCJPbuxRpM09QeOLJH2PSx1fPF7
6UJMBbW932dHBEWDr50HR14Eu6o+REL2fs90VFXOeBc8M2RIMjAEdTdkV07vGetXK6MAC5mfSWAI
6xQDTWiFfvh7U1Mprx0tWtNSbktjLMq+MlAnD3al+XS18pZFcXnoiB+EP2UbhfGUumHN+Ln71gCq
77dFWViYPutDLspoafH21vTR5cr8pAv+P5m51WFfo1/uY1ke6xer3ZN5kw/IlLcctFrLCtr8Sg3o
uXOaPb2zgaV9Aj0I9NMTscdIrynIUvzTJ8INmOxjyfL0xvbK7TnJj9TgkELRvKnWKLJei8YN5kyV
h3L3zYcTbaAxoQtLfv/+ETCT1g9PhZhSZFcWl4behuHyE6VwMeo5Gv/w7Zjr9qt7aSBfyWJojnBY
NtcqGmSOethCwxFqWrmcW8ip/sBojxR6QihsmhPRewOFXseHtlcFEbBXRXr4fynzUGaoBGUK6tDJ
aUEnM+D52JeGCRT1R5nAUbFVzJ0YSzMusbAXnlSbjrocj+3eOaudTdNFX79Ngkxm2KcZqotywUbP
U8rHqxb1lilwXVgNfRgsFBK/YQ5UIWuwxoSVD1Ju+Nl0+zQwI1w8+YFOyH4W9ZTCTlPV+z+et8fb
OE6YwO0o8lRUZKTX/4HMAi74OwWqzmxG3dUcygZ25K5G+Cc8awwfvUStOLeGW6VY4unvEgc/Zgty
BPhwt7aRp4CXSGMQFSFoc+xBHN8zVzmUQI9y2VLNtUOx5SguzLo7iFyogXZqFCeDsfoboU9jc7FS
NXlKHqH5pAAZlQ07oddAo2FBKYqU2N4eJv9nmt0lxNwN4SYGGfKHaGaoREVWfMgPXwCc7FYVD1uc
dgcM5fqwSrJyhYaYRoQEnHZbPo81Kf4HpPoUpxs2ObiJlssZjtcJowxx3REJD1+A6wo1AlrZWQli
M12WmjdWcAVh3nWY4jCt0pPfFHWAKMbS40SsFIRG2snryDcPQRWEBSilb1bgiwTgaELP62cBsJI4
EHlukZRQfU1ogJyAme8PJdfTORV2/tUjo4Ols3NJ74tuhmktnVPYE5lRkhmkGz6bGuunY79Vf2Mo
gwAc+Do4k9DJqKoUCv1CUdNC0huJVGgLi5r4MgkZV6l4hbszEEM94XrGlLyPQsoZ5wEaRgk7fGTS
tfg4nICbCdzRwRSI1YzKbZQDtJzk2UUxlMH8ckgXwRKCXHhlkDbf3UeRx52EAJUI11GX2XipXkgD
RVJhqxSjuwYFr6xemjUJj2Ut0ePTXouEv0bEiIlz3nbs/eq+/6fjWZqbbHbW3YbFe55G8chRCFDu
ykImQRzMsxk8409Gz6T/ATxrBjstrJBXEPi10mYl9+yFSZkk9dbiWM46coElgNMNRvOCzwWo7GAD
VHqpXmPCmSChq6JVPJOmX8IODbCuU+9v53rpbLiwEHfEqF7oFqjQvk9dZG/6Z/QSdf6Ctal3PbV8
PJFQf9v8/nI72mZG+hQHv4agg8ITfRm+KMlZn6y0GP2alsi+Fc52d+GZAbn4z/kiy5Nb9krxbPS1
n/UHUo1FsxHlxguZwaAmaudhlVd7B84TaM+P689TvGJWlhyzGN8eIgf9/Idz5BsvtfgMgBHvM3qF
/WOiZ6H1mxpqDXRZeAPrsqCdV3HctiDkiABqPF4b+QV0SAK/m6cWwNDw33CH2T/ryyb+m/W+zzQB
jKrO4C/NdwBB++G3bKuCYhTj2crNZwhd71j48uosRKWQPPmZfaG2bjGupM8iyXy/l8x3XauvFxAk
io3NW5nNQMt2UA6Jb4yd3AIoRcNhx3gvZSi/QADk+EtoekO5P9buowKBiggn7C8FPsCR69LzQgAH
X6nCEnH7KZW3Fqjbh2RJm61yCeO/fYnsmXrmYS3ozQYFkJ2NQ3em+K/ZW14klj09+1SIy4993JPr
AHEO4+4vhNx1e7oEKusKWywXz3rGcDAh6rnm0+okf1MypsshBDGGL/QxzALK5+qie2nS7q29WKZn
q2m5bXiAT7jsf+hRqtERlJRVgAXYeSrOKR8vfmSQ8kZIT/HEesg86tvxp0UML75br+SC5k5eQyq6
7HHcifrOY8zHrtzBC9NJL9TESgh/QDJlF9/pVdKboV060wVBrZxaQrxXlU/hZW6Sf0zTWsLV/wpG
yZzV2wKMPUCrcgMjt4ifsMFXSB+O9I6nWPeCh+pNzUfU9Wcfh0Uq8DQUjYnHfY2OgydPdSziyCW9
ojungsjUV/ku8qQhwFLhqL0JuV7bWctkW1lgjkIOudWWd+0o56heWoCrmG5UFuU6gwSNYBn+fNyy
EaFwycXyhf2XqKno+cpqotxJ0o3gO4c+2VyBYFR7ZvpZcYZZr75ATRnx6lDqyQDcpHSdkRZJoeMR
NE+olSTGtx/IDMpA7ZofRzi2MJGheCTpnx852uaWvU2MzIk4pkzcs5uRKAvAc6JLQARmRY0HtFwM
iraIIYUv56YRJ9p56/UIskF7P131sIotvhVle9j0krSlIHQ7+lOAcCfnbcCAuF6PjXpiFjxS1I9p
jk5yAi4rprCNhcs9mx/4hy0hMi954keoNTRJicFxiFQ32PPgBQ/2L6k7H83aSvxViyVLcy93lE3w
V/CzqfzfmHNFyhbYwjk3PDmxJvEhdMOTeOl3USoqrsZLiE/gVTYsBJfTYYNGHVi5CBdBKS38GBT1
/W8i4nm96WYYaXCJWYdbLpmoheszMU2+9UGgyHCZmzEkSRgC5rCaplIXDey3kZ6I1OPqayLa7hnR
Gx4LqDeb2wrG9Pj0XFI0sib/dQ7VOlPTIQBPmMYukfsL4lv90RmwSNGHhs2hK9TZ+xspDW0tSksW
QhniuCKigE+WQpTeDLOLLQr49xtXj/baWbycOpl6ngr2kSM5n/wY7cYJasegs+ld9LU1AoRdHq2E
8j0uRoBrYzLAiEE6XOPq2YM4yLgHhfBZwVJWsYnived+mx+GOj2/yhG98vFHCphj8I2Z1TzRwtfR
t1WOTWXjXM+TsmHra/qQjWQPXxvGqEDdtDFLv2hPl6hmZL/sPfY689PMkZFhZCrFsWMZbd8SRNrk
9Vzc+ou45oq6VEuflMFyAvLBjV9z8aoeulccdN5BJCFxIMuOjppDA0kO4nve1coc4tlyHy+NzJvq
vFvq5MMDP6VWJbhst239ta8+nFnk68VSatz14TqfK2SvHzKfpGPLuwuYgInzV6vqpDuUPqrGqB/e
z1W9YlqBHOOrPiPXpQrm2HJWayayQSHm2wQSMM6hHw+cNLypj6qkBCxVmg5Wu4SlFbmd02k6Usta
6wYTmtUzCUVLrzTm+hY2htRHaUzezDEMWa+0jM5rbX8LwfAFoYlt8zQu2sFMuON5WbhaPIKPDPQe
f6KvRNsykgUiystYTHWoxHTfJ7P8h0Kt2xy2BJKQkFPq6YlvdZr52QhsyZXslOgPDAXhTfJxJXl2
M35fMw/6I2nSgo+zViBmQ+J/w8jy1Ursdq+sOpnq9v1AUJxk14Z1+f4a5aRMUvkKi9oMgAmJ/9cl
xaLocP2Obi+RRrNGnfUH6nKnkdvihbcc5WW9a6j9rE63J7vHyaPqupbJ5jhiVoEoorQLOk3Z/nLG
9VznFvkXYPp1IQYmRdhcriRlFNetKH+mtkrq2QO6g0eUA+vsHWvKMTxPyh4PzY1iDX3r8DW1Ezn+
CafyKC2l5IwyC5/nbiYx0WSYgxjZIqJK72l5EWG4MUHsk871kbu8mYQE7MEYCplz1luGzBXtxyXC
PzdgbxUUb5d5y2iMGRYCqFm+NRBV+B6RqcM2S2N+qg8tn83v3ISDFEqYvRL0rI3/3fVF8VdVDwHj
04pOT3NGFFGwc6qcwpmwdQsYkHjLRrkK0cQoFPMMpyVFuFG1Uj0w+yOHw/u3Nt4tc8yib6zc/ZX8
ZcbmdSkBAlVMAuwzr0f1G9pycoMDLMH6BI1KHNsr3XIdcfTwx+G7dLLrb8EMERVCXMMY/JhagPbO
8JTzS2MGK6fIQI9mVZkFdlG+fxqWDVIPANveWeFmP/e7oEimBSiydPmx5mfSQfoi+W7x+r81sn/I
zEwYImF29DocGKl8++XAOmFSRkyAWghXvnaal/DY5WRz+BHvp3wUuB8R7L47PEkQbcFw8IlcxZDl
m2SPngau5UAVk2yqe5PjWIjtGZe7ruJzpMx49tIoNN4hdNH7XXi4Y5nfu42OnNj1PqKKkIkH+Sni
9wFbF8qTLVDlEvFGoVY/QMk2fLwgn2B8kfyFy8+VJTrNuMdXOr+/sVvWKRxjDUv0QgH7Q8iIfNWE
mXjnosze9PA7YMEpduqISXqvaycOugcwgmQd+vRUR0QF3gk6INPGFYGvCBdO1BGVPKnU8friugKT
Beof22Fb127m16P4PUU2NK1Wv4z0AfhRLiNqzaUdWoNYaj6aOoFFRKh4NwNa+Fo8uCLZgX8lAzk1
A4QhrKI9uwQos8zh0wTf4SI4zvIyBH1wptnjWVsMXaWcr8MWXlPhGuk/MvbqiQPOwbXLemkSEuTt
109Wrzfcfd+6DsydBmcjmiZvkTwf4dcAsBLjzBGfR7YdsMnU5uSVBCp3iEw0RhdmGPWTvXWB0WDS
q2ssCZq6KIKNeRKMtPSEYP++hic8ceO7IawPvwQFXDNQV/d+YxWPF3+dhFu9mCSzpmUXuyCKhXrW
EXYurKiOpuiVlirp7Iqi8/o9e8quy/cqhNRqNbU8gA0DOogZ2Dy6Yoo5xL5eKUPlhQ+A1TZhkNbS
yOxhC82ooZ6spZIxexch8R49wRSihAqFAKaf+VYbOqPggPIkxBfMo+aNSVo0w0CJlgMe11TjMCRS
KUQE42h7QAlP9ja7PyW13CrS6uh4SP9JPuQAJwbz4lhV020I1z0o+Sv69FhV+zgkq1nOqPdjBL/E
8Vw4yXilnHqE87voRiNxjozmwgXGHtgQrhnC0GvRUXNLL6HGUn23sBbTtKIm69sXofucmqVGP7WE
AW46karV1YO1NfRm6sq530PciRW/NGKWPstCynK9KFOg0SG5XryJK1oN7BeY6VxdZblAYBpc+45S
JTiiTA0AkMQbeMsHZg1AoUDBavTTGza5MbXfJLB2gD3CzyXHeIDlhcl+BqH2J4ikXSrB009lNQ9w
sS99/mcf5ENXFCEW8h0O7kqekaRiwwgAPMWNUNT0Bj06/mEgubArcEDFa89hflKaYco6HSpRpGq7
wCtPji/5XluLD+HHhYHNZ5theajoYg2Vt60Ax1pZ22U89WJUWU3Z0NHptyNZyCtG2Cj/rmr7wXrG
Iq4xh86BoqsSGGFc1pHrZ5JR8A+BJcPF8IFjDgIUXZwjY1qXy/FoibtY5Grf27LlDt645vghIxW6
/ZZKn0OtwWXIJbP07z4hvOalN4X1OXzxwfSMicJpgnsiEVti6bbDKuDzQtLJgHuQZ5qTktrLhyv2
ZhQ9FgMxVQb50V24qvQu8frLVH6Orl0uPSBUaUUi0vvAVDpl90tZL3gaJMVz0uUYGcWNRxcNwBHK
nVFazVoefFoU70M48qeN5ICUNrNLNj5zL+zjbacqI0Gp/PRnbqVpQmsloeIMu4riiNpNUsoOtRWH
qnR87NYXx9WkDL8dg+YfESCv13NHD6V6R64UIl01zHrHvbpOuHTptFvwykUG9m9u2ha2IeSFIVhz
e6rMeg9RFhsLPdXB4/aozIE1R8XD7kLSiEzr771ET8YNe0fmGzilZbJtmi0bB6Mglujs2WRyQt9C
gi/V1JtsBndGwzXwCGnftFzeulSEP6Ju0wedDmwZ9FP7Y6jay/Nu0/bil9VBQNU6WVn9QKJPu59M
CJknq1vIuyk/RbWjUY3kG8VhDGbb0WmClQlyBjcwgwlXTqjDmff9DUbocSMd4QAKxxQdwEFrrDwr
Ar0Y5kIU1a1gCiU5KUzW7JrPFnfOYx6mGg3veGYAdF8FXjlTWNuFbbPpHeRI7C+LCOo1dutqy/MJ
YacQ3H2nw2WA4WfyHrYu6ooM9onn39dIoeEERKq0OZjBO0Lsb+g5QWJx4t4A+tzG4/+I113nNOD2
HShvuwVJgw5fYuSrdB+AAVvBx3anllJ7q/6+IEvyzqJp4UfoV32L1BatEYdjQEGNv/llpg4OaJlM
9nabE4eppOqAjjH58krY1g/KCSuJEGYpoQ2csd0lLrd/2qjZxbdDxWSpJrQ29hFGgabiw3pRT6zl
WhahCg/ZkO1MyOp9n0RVzaHNzXo95CRPbMwZnkg42LPdk+c4dTe60NHjUQKTpd0GsyiRajG8LKPv
TdgGj5jXWlEFqmK7ESCtPvmQubOPw1UHeS87QXIqUG6gJwq3AI8xH4+XOTZ3bDGOT6thQWWiGrqy
/jtgIOd4JvsDe+rkGpLkE2CXLp7BiPNpoaOS82nokqa/YS8qvudhexpfZKzeRSSjlB/WXFp0WM1n
HY4w8xhMkBTlNC2RK499N02zmljSJx3WrLASXKuFdNKzfhiyI67b69NNoCYxNMUA5GSt/pwszg/x
P0DAvhAReQpqepXscf2ZpHfBp8B6iInZhrrwIX4+9LvX+aqrr5tJeJF5JxIdItcOPcKFo3egKP44
f/T+XHy07nTsF7j7t5kVjrQVVMU5CYZZqcARAL+aPXlVDCZXHGUF3r11A8KY9mh0mSX8TsGcrd8a
MlgdlLg16COgFbsCgtJSjDsKE6tTCtGFxaz9EdZinBH3ZD3Wy5hG9+rf90MjQXHImAUMh4FZVhkM
aAdzXbtwgock5FstdDRIGPkH48HFEwrl7KNSWsiDWs18Ys0AMt+1TcIjeM+zZkKJEttsnkCHB7dz
cEJCD/Z95KQANoDCLVzCiXMpDGSOMVzQTAqunrWTbFyUGRgJcbUdxDVfpme/4xFct2NVlMiF/POq
QIbKUNxFBnPF5UYveFM69pcI3aWw7F9W8wKjtyaiC9zW09MsHFydL6cDqfYin/nEMSVtKdeTif9z
g5XW8MKLG5ljJMBSbUJujxVBTK90xJiXfHNjDAOo7NZ/Ux4M+gj46D9byMHhNlhotFkYprIBCLZ3
+7GKAvvpNE17CwYLblc0FBgg30a0strjSFmwQwk1sDkEb+tOl28uluyVes1IcxRCe1CTS+eJfDwq
3v66ayVegFf87GmjCydXIK6cUB1DSYcsoXW30DXCr0bmt+u/uJJOeE8PnwKr1Q/OfxrlkVCOkWtR
viZroOvM9WsMq3Owai3M3FSE5kYoRhMmLp1EtrR9zLjQwjR6kcBQlbO47eJv2VOLMqAfRyaiYXTb
Eo7v433JZ8cLrTyNPrwvHyo1GpohU1nxTftaMQWQe5ZQbhAlTd02/bHrbOtJi4bgHsVZnHDNgpNV
rvscvxaImB37mmSLNBo2AfbFiLoKodoLovnHkRC4IkHexaaL/p9xxDGsF4dI5VmtqupZN4kQcuRK
qSpaEmpfOOBAbq/7kfJAOD2WF0rEHVgIftYXQn5UtSTdWqQUba7CDUrHZk+qe/UMOnRdJqOcm8iw
7MudmMqalxRbJ4qiJ9rHCdqWXDoJmIGz/IexKOVBuvNeP18kEQOLJxcy8ZBgY/W5oT8oe2JjixJH
GHGULD/YRI4wp1IHx1f/oj/YHoBjsDZgLiyGklHMcOMu8N6T1/UBwgSrOKQBndHeqHUq70Ae0gHf
SnzNkvG6zRsRTy2QTX9AGmGv3feqghU3IEszNArBgRrTPWodex8VRcTe2Vt4v/tVn946j59AF0ht
b24qrYTbKjnAEesVUyRDe524pwieTh1I6b3r9dltgrYS7EI+RKxpBOIh+YjpHl1tDjuVb5Irjc5d
DrtujyxzJOXS5Mm9Z65NDSJNIYIAE6eSs4OxmEsegxi7JQI65UcW96BAXh70cJxKfY6A9p8Ryrt5
Y8pdsJaoNXRfJAvTl3xOZPAj6km721BDVBiNczB1aHO+ov7VkuDcRIPbNr4ED5eDz5y+eqVVjXcX
5Ks34wpyGYOJKjPNJlm8rCvIX9hrZcODxj+KxDeKDpkR+KlcrFcqjYPzPFFXzZbLSXZR8dYQMvYe
9OIBCwZ591Ak5D5XGKt2RMHiis0KBbCyZ/L2ESQtmc/MJcGIKZ42nFEnKERNADOfAhNPLFykhfy/
LBLoD40ytLDnDkTqkqOI1Bk8viZ9s/mQ4acP7lyu1LTxe5dsrJUEuxwLwNI4/QfiVI1m5AG/OZnp
NGn6KqIbG9Qvj3D+F79miWwZQNCATyUJfCwPT8vu70PVVcE6VlODUOB7zCH1YdlKb5PmXudZEv8a
MpvRbgAsrqbjmyFRbuAaaN4Ij/lnGhHfqzKbVZCY5XgKnj85L4k7X1xlUGjCd+mSa/T7mAaioD1g
QO6L+JJrv6JJ+B3x/kPF3jeB9STiQns2NRSQlzEZbb8jxbDFQkAe5WdQOr/pI0rx/bfU/yG2FZOB
jx6Xw7bz6e1LxRb2oHkFJiJftU5LBQYyi4ZTXjW5gK/Vg3tkh78ebnPQFziu3epRhmnqqaXlsG28
lmOmXdmolfuWYy18D1lokkeRAEEyIiw3S7Yf046X1IEsrJF4bImt4IYhGOPQObW17H9v3/0mbrWJ
UaA9/owWqfEfM1qwyh/FXj4gOsdc02HRXoQFbhjV4QW5DNx0VyvUDCfeCzb4xKCNG72xwfUb0b0r
ZDOoWzpLfXgaxlX5Zq/v++CsVfZZiqBG+wBfp1Q2L3hvNGukYip0Wg9iuPxpo/8P+lSuSfOc/edV
AgjZB+nYjJWwE8xxcBk0zcVnrPnfeBBbAhAlWZIeahqfe2XCmjjiduBquOBaoH7C7z2Oq7N0uWBr
vp0p4OxdLqVIU6W8V3mEyXN8bEcwLIOmZAWkmUOcr8UtjkWUn0VsU8oejg8LE/SrbIluEOl4r8yn
8lcSNVTo7zsa/3MZQrvrdkWcdIYTzcLrjIGeEZ4HYNjui1HWnW1bgAYcI1iYB+7Spv2+5RZAMh7U
JOZQVDe5eF9lG3SgQk3UuwoGbz3RmBZIhJA3v7qoTfHSUXp90JRtDuAb9WBQ/7/24ODNuyaVVgJc
DQ1Qtf/8aj9bQC8im2QW5Z4ZLRQYOMr9aE8zm44aiPA+54woIB163huBcRCTcfLqE/hGjMhd2W0G
eXCtk9Ma4uVLKQVwu+wU07uycU45Bzk2d/1GLJsnXa5E2xRHg7bVz5FeVZjqA4pvAi8j9FeTATbJ
QgB+99Fhe4Y5N+7lo+fzWmv0msycmolikaIwU6ra2A6i8UjYcRvClU14g1rMTRMSLID25bIdGTlC
yERg7eWdaij6Im8PhpU/Grjd3A6yOh6oOyUd2YfJoUr7YWtQj242Hdlsd0Wy5tlRnGgwHQFZ4hEA
8yNwqm14y3smEFtXF+raAC5sb3kiL4kT9CMWr8VcS8leh3Jyoy6mq5zFYmuj77EXVU3TMnobekr2
Wf7UzTbF7/5tQjDcIej0emULtYZe97zjRXPIV3/o4nXAndZEIJSJ2LjOKwlTs2kbsN97ieumZCgY
JsQlSu3WOSXGTBC6WAp3E2kkQRFfQmZTjynXWiRBAPEq5iOOHA33yNHTmXHz8BfV+NZHlJqLTfQY
0t+nP4bqxIqo4u6ciFNuk2sBoljYIkXV/m46k6X45JdhF4YA2LibOUxaVZ6HgvZnEFSS3GfpuB7S
cU9YOGHigJyRm3a5YxzsyEBMVCoPu/qllrcvHMhAHXusnzsazxfKBRVI5fWJXz0LsaD8UkbIpoZd
RnL/43q92Y+sFLVY9b9BCmfrqHUsUxfyaSd1mIsXTuj+xsoWuazwHRWAKtVqVUg7DJID7UAHUoI6
s1XtWKkwHO6Bkc5ZmZS2PtpF7Jakd6ePUgHpUbhF7U14ACHW1KrBsVGg/mjksvMQClA6imAjjDAJ
6+MKr2L3iDWzl/pIMS+WvYa0D6/z97QC/DyVoFugin96U5X9QiDVLR9Jmig6kdHFSOEF1BIMQGtl
G54eYoh0Fpb63FQehcFgVHye4GJjb6MGUeXqiWaYcLalztAnpswE5LWeQNVDTL79ywi0zIizNeqr
lu656toNIps3k6c8Q1pfPUl89E+pencarVTxTiSU/qVBR6n10REbzhXocBzYArwoI4P7ncWtUL4/
ticsVXCQi5oR7mOs53ohJZPjHmwKvQoClU4IIflcV0vofharV8ZYS1lqoN25v7J/IrmW4svxUigP
F9D8qcS4XpLln8ETX3GM1DBW0N8baEqzt2coVJ1WnJdAFYIaa8+4tsABy27/i8G/OyeR2Y3jQDQ/
hXeVVJtDvK8sNAaS1b2jQXCibuCh2UKaizBKtjIjK7E2ssh5W5Qw70/QskqaygpX5W4OKHftBSyC
2/w1HhFDSwHe6pF3mOefugDq4kLTu/r+qv+W96Flg/oxi9qtw+o1755nmVxGD1SiTugqetwIETtZ
3XPUxIOWqy0nZbywuyqyt2rXHGJI9eR+zhnArb+Mj2S2lEbFqnRihhL0yzSgZ+hHl/wBFOJYmf3g
bFmScte4kcg31iugXWROic6/jkHppBT0y7QGU+B0U2YXvaxqg0ZqCA7Dk4ITkaUmKAGPcKEb4ldc
0oI+lbRZz9ciNJSEMiuy3UGImdsN/wmdchYt7DZzRkN60UEAGOt8FaELwa+VYJfeDGOI8MtJVUbm
MoREh0JNw4H3XWgfD6cpOADAncydzCkyTJ0Zy5e64rWMqKJhhAc08lhDDi052sNxaIYmuDfRU4NJ
dgeslqmn1famqdrGFte6OBU9haG2T2yEoyS18bOWm2HbmlS/UGRwxMb84NHFKayaNcrHuDOwRDLp
BkGcrnM8ypp46iff1Uga8oS4/pZ28+rs8ZVTjkqm2l5GR64vUFAuD4Pt56OQ5DGRTuDfBoJj7AfF
eS26FSQhQ0igKqBY3sPEssshaY4qrnMtQhuhblT3H7nXhYJo1+T43/waic6oV9yD4Jk+3N0AlG8U
YUmqyYnbfO9zU8aCEw2pYDaUPpaGm8NMzCp96qfFuv5vnk6OoMTdu14bd1nC4Mj6UDekvpsyI8Ne
VHVlCI+EfykZf++90HhfiWFaalvXpJcGpJEzLKj1fC4jH7NmQven8QKiOwdVddvkc7K5Vx6U5CFe
JOlKfXg/Ixfi7yvRo4zKTy7tpgfn1ZijgtS5vI/i0uZ8c92nDKEnRTNgIUxlMXPxdyem0aGEdDTV
mFMDF7Jq5OUPcGRnnMvQuX1t8Ya5IHkLgyjrc6EigvBpwE8Ui9v1mEV4JgPg88+gM8biQcGqNrCW
P3qoPSJPv5nzFN4mHfHc8E3gcqaLag8Ujc6KA4FkDiLs9zmJ0GKD9+S6sMjMVE8hbmC71sdoWtX8
fb/kfh5LpEx7dNn4j3vr6Xz7oB8k+wZSvaPmGr0vsziOxP5IPL66XUOl7b4+j9Tc1o1PKWIqCicH
5WaELJmvJk/MZubkj44hke9W3MM7UUZsOVn4YfBgBkVSvZo9Mwp+J019lO+taioAmeMFNxwG5ep9
Ccmz4ntECySbf2QAgdUPHKCAz2mp5DJJaCI4Yqo3LJMunP/y3TpHjbOdfFLNIn+SVjuW3BAVT+rk
nxZNyzZESlnM7quqzYI3T5e+evqVqs+gJ+M8fwvlMCjRoUCDXCUo3kLADBgX6XsyqHonHgHvDcpI
bUZ2WO6flOzloMI+uCtesdl1wu6K7FBJeK4I6Vo7As46Q/wuTKbv+oElsuRCncZD/vDsrZ1A0LTz
y7CAxqIba4lSCIz2ZUH2j1WrBmg4jHf1OKNBwouB6Ox+H4pQFinQzlftPltIqmKVrmfll5xmpFtV
57fGJBnVN7QsjNQFkLOre41BeavDUHJXejZ24U0CZZ1S1agRWBHWok8zecawvpD0iM/udwkZY9aK
CFp0a3BtQUy86h5F2XE/gnSqaJ/E3QDUKq/bQs9xaTqyQQ3mxASGro3ijngO+NXURcNZzS4qgBf2
W9xKuOn/cEZVzLAHL/ss8JfnxUoK4sjoJmbZjmA6yicHQhJr1JAFiCoSXW1aPPU7CHZm3vB1DaP7
kAfUDTUNGKFbTsfT/QDUbk44+VswHa35Kd/NS87PVNNShxhRoFXbB9nDTjAL9eUe0GL+/qJnebZe
ZBu7/UiGk/j/O84L2lg6g+5YECV9pTO05RBT6VxDjIRgqtxZ2+uMZBjxVGFqfWQiDvySEqAgborf
RcPMOz41Q8McRlaQANl4qnV2r6rWsrcgvvKq3PA2k2jf8VrHrIkWF7RdMb6xom+pGShaSvMn5ByH
nfXSbNBer64J3ydkectaV+8AYW8HTZutkPX5LTQS2QKfQyB3xsXuDiDqYsZ3Ri3b15X1714HC+Q3
QR9Q8I5laCJORMFvNVHeFTLpiXQFuj9NhDjSiZUqxWmjfFHse0RiXFpm1ZjHgfUN535Yc291tceq
C26EgF1LTnM+lHV7eO6OuMMhJhH5q6s0Se1LualKbHXsp4nuicaYqFNRuhhRdwnU3PGBqG9E8/gk
r1vxPFx+fGCHkfyLqZXvKMRV+seN8zwkbExIcPTUxbEC8ZiMPam3Qc5xIAh+Oj3WvGbtJHp/zK7g
HM+QnHqblJS+KRMzMEQYfccQxfnuWfP5WvjhgRGzm6XkFtwEjEaIj/YRQDRUiwmb625ax5gEHERr
6NucvUhIx9p/XthKp9yPLnGEVLlyxl+gjQlS8DRt3xdISDaZNbMsqhmIZJFGHMD6V86sEBl75iUa
ZprCUMTJbUASNDxZEFbL/ijBwgpw0nOwwX6N2RyO8b1hBdOaGKU1maMp2lbaF2AweK1FmCX2oVmZ
10nSPpc/WeYvG41b6F1vpedQn8AAN5CtpxvO/cz6gSuZWAjc/XGNsFF0lRIxwWzgnAjHRdooKbDp
mLrnLrLLxhVavoLct5YvgfrE5ZN+OEN9iL2pyVXSwE8WQwOGkqq4gqQJZO3QhHgxQWPGX3Jx13Qd
R7inXgyNIUBtDl1O2yBt8fOMxIZmUfo08mPxICgR9qR1xwci3IzUbtOZXVtBw7/eBUU6LbFhgB8z
/fiDQDgwCRZ9uGTNFCw4EoXSx5SHpsnFCx21Ozydd2w1QROSPtI/usBwzKL6wo1fSkwDDU4ByZA+
QmXKznRc4iHsLFTxlTfjxn/WgAe0wDRJUUXQo2C0CpJtlmagqwMaqrBvCtkJs18UMFLJNC3g2ZN3
eVviijPe7z6CPrUPUlVRw4Tj34veGaAX9s0B4GRhNyqYGcLJkvrt8nY+Fh/qtdnkiyfyvcyZ6DbM
Lcy8LJroVpxFoWJFMzsk5GYqaII/SGXfltSaAjaJquwd7piQcFh7S+UcmoXb3jSFuD1aUFeV8/0L
xKIJ+zKYkMcK53mfjqfBYeUvod336J86HgA3Bcfr++gBMLgWfmK0C+cTDjWX7R2MZt9Xmsmf8Nwb
TtVo6cVuQ7MBjbLp2JuscK7nPhcFbADjGq6WaMxQbC2MBJE7gwwW1qGxR3Vt15Wx8dThYkLi6dJ5
Qe5hChI6iuyr8ym5aHICZgsb6oQ5YL4LkgQ3tK7q+N2ug8y1RugQo1pkohilXORIMzxLE+NtxT98
udx5MXCBZkqDxUlQOrTOdo85bCl8ScS45OqnlDj6H3Ya49P1TFiJrls/pTQupmwXiaJYCXKiD27o
5Vw6yfww67jMVqmkGJrw7hCj7pShb4Vnnl0gkz2eNrgJvVUtqNRYpCzAmt15v/r9KHC2RKxwOfAQ
K/dTrqn/ZTKf0O5HsPLwZ4q1fFnD44TOQ9zgLRuOBNrm9bnHGnos+qKl9BE1Y6AQUrWY6kPO5EYx
gZlrFI60DeqAWg7WAa5Eynj7+iVJ9HBDTSCNZUalYYSu4kHq6JJV810ulnRSQVJ7LsL0KQjCEbkl
3oltSS9+KKZo752ej4VoP8/XgieqpxwHYB7TGKj8xEzgohZGl5U6EM+wNgmQUUUgWLLbFQYor6a0
36trivGZt22vB4hKU0FlO/Ddm+/xqBsmA/cVNBoiOJyE5618MWNTZLxJpnRInZcZzUIipeGJHdHG
gPoO3bn0zyHAfak+6B5cNv2lflusKXUtC3iRBkdSPQ7LONIcTCLZepVjsjZ6ymrykQRzrVxXXkMS
5PWBl5hUwnry0An0xZWhpoXW01ja8cRl9zWFNydmtli8LuYlhkuEgGvGD6g8BKLw21K1CEK8c8Di
ao9hkv6tX4KS+B36iTQ4IsZfS/mkDCcKM2WOplVFbZK/cSZ78LZMyRMyOHGbF0+tdOdWXljPoqBB
bTCLG2VZot37Xw5GgjunjXzjjZ+y1C8FMrZsBwRdCVXXau+dVsInZLy0lCt+G7jUe8EXJ8QMZupC
x6kRBZf/DJvlFg5lxJycaNkafxKXnIwOl2xPjCcZkCQiAO1EZTk2YcgR2+IpLZUF2tMu2U0Imtlc
35bOYljMlbB1lr7pt6ytzG3hxjHvL7mPgf+AOJ6sSLFUQzM9tedi719W6NH7C0ixMbe2slw3LxZL
s0NE+4rKxbOSdLa4JczZvAfqVzPrvLtcUgKZJkdfuPGt1km9vSqIblqGIePfmvTqkWz4OKibK+AQ
1LDjxwEzn+x/PipSmJ2bW0Pf745UnVgqKClWDtp9WRdnAW6N1EZPWU5PnxzQXY0dXbv63XOVOcUc
9RtDQD11kY/78G5C6WGeA1hoiMdE0WiT94xSC+NGk+qMt/+VdmCELKzd1ViPa4GXa8piVOP4bOYU
ZMwVIKs83KM8ShQuvDRzA2ZqVIeXMp+YBbh9BsAVc+X3K6GXgjlwKVHOWZtmM2BpUqGsGIoMrfr3
8NZ2uncCY+9YnTYJf2YEUnJlwT/n7rEId0380Jistij3XcmymoXzNTvsJzjt+y2QcXdns+bTyxR8
3j7ZbWc2WvZ9KrY+XxsYj+uaJoq2hfdfQf5P13Wv+mnPuGZkfL76/lHBg5Y0TE71c31EwYQGlBwf
zr3OIiZQ0A64mP+TqKG6PZUovXL1+Z8Xnufbpx06/Tv2YPkFYknbNvKMUy6uC5Kx8Blzed4EE3Ow
Tsnmek+7g9dMS6xCgZUol92wc1QD9WaEGuBHoedm6IP+iZH50y/UG2w68/zBG75YIMGTk7QtF4F7
aXekzzAxo06NGx/UxZjOkijegX4hRPLFkfS7nuMRfbm4Ec8ncBJ2/duN8HA8cfADLk4jBycRWs8m
pCqQIVSDYMuACDSFk3yNOakMn5OGwWR91Ad01JuYJJuDA0tFbkMkNVqD+p1RXoagdvYMqG3tOQiP
KnAWvDPldsicPVOGSnAFmn7rk9kiEOzBb5o9JWIpAQVzZ9yr66XGqKFGqeMWPQJV5eKy2CzGuxrs
9Kv7l3B2USLH3s7WECGLKI3/6VXdxfer22g22ZrRsJfXj0S3UZ68P/aaNQSeZGTGb1Sm9NHEK/DO
UQxv7Kby+7j44bUlCnNt0qhkj2zLBOePEt+eRtmXZ9xVIVgB4+EDhYCfN6ezaXn+BHrsI9acEzqE
sVynhtjG/lgdZe+wvAxp3fNPXZk8N30qv6c5aGJTt9pNDT36iHvAuKF9n8wZcBJJdaL0mbsf/B4j
zPQJMAJKgJC/GF2k3K9eiYgyOs/Nxz0IfF2OxAfPkpFtjji/RuRs+NTforMH2+Ny/ulLVIiTzmW3
+3MQgFL8IoQA6Y7SZZ0NYT/AxyHTVqxIeYpW8A3ZkBnU8/m2mqVkTCI8qpszdGYKYjhx6pBbbxt2
aJDsO+0lDVFadptH2wSmKghJgPlFftXWOkuy5Ex31R+xoIhdR1P6TAo9k+cIFpr0CGFWD+Y/sxvA
ky8wBldP0ZDw7LIgUvrvjNOz+qpKa86JA7p5kqaaOzop1uy/DVZDZGEJq5RpYxWlH8NNpGyxHELy
TcVZ0uh5AplE4wc6gFVwiyHzrrJQ9gBVFZQHVtXA5HYAYvrdoIzlHoEa0AZtSW6k9wcWDWhPUdvX
IXQ+LOXiDLQWScU7sHAeDb9cAAjGBoezVmMCk+QGw3x8u0wOB4Y/e7rw1PVkzSyKLPU6nMnwc2rA
MPabEq13LgZMsBsHMTGUji7YBzuSv3xOGgnCgJfzDq1lwZrrEUr3glpOOfFp2Nz2i7l3gpWXZLev
urxfmryQC4SxAgyC8SuvVgJ7U3Kchg8vBCrluYujSmX0/FqZLx9Q5b3XWlORtQmie6LCgmvZID8m
0KxXfEUvv/y67WDnDLapRotE0YI9CXFZI4FRSTCYon2APC2PZCnxlOT7e4Tsha35Pe0DHK/T8Btf
akST5vU+pUCP1qMKLN1Y6T5s4iPgYZw6fhrJL2cX1aP5pR+DmntCpdzb3MKbJ8pnxrEKbOB98e9g
T5kk7IqxNHRJy+WvnzzkgbQw0W0VfmJyP9wA6end//SBLhoyEEWLLmov0CCuzhP41utokZ73KPDv
86eylULhfTby76+Iy+jO+x0xfkz/TDuETtmW6QLfnAYeLgfpdT4/tD8KD8wAQba0IFGemQLhI5Ul
P0d3UA5tPWYxSg3+SftqhGq2oVSCqDK03tvwqF34aPY13RoIjUlAWp8QHkp/vr0Bs06RHGMFv/rl
Sc6YthxG/Ow+zixCrMPIMLtLtChFpQ2hA76pwEgG9oIfqpn6QYPfkeuAbl/4LgLL3GHl9/JSXdiu
4PGX9l+csz0ylVFhsh4k2ThA6ZigD1LTcUd+5h6Tg0HqIGwR5LAHuOICIAWFkb/LAnRtyFJzL+J3
zokUJJd3hThYe+DvT0tZjMmxnoxlrv1/T4f7gUyUfCqzBfAKMl6DIKDKBkQB81mwDpNMSJFY7hct
BfafnDpLn97UzcqrR42dIHm6+eo4pRsFtaYQ3C9MiXovdgCocUClmGDwL2QePC6FqmnDxARCqGMS
14vGtjc1HVnio7MA8NHxRWNlDu3faSmn43AupE/TOJBcUojByTGngmlkGOmjFPebI0Xzoj6N1Xkb
Faw9tZsYdNVXFTMM6ctkZ5B8p+V4Oe+cJnQKkJGs26NO3N0lcefYIFhMzCeLXCWZ64VAtgubbO22
uFis673oSO+876Ju8wpKzRZ3qhBA0P2tTasg9FSQBlriuomNMUJk0XxV6rkNJzL4R/ZOTmT3hCWP
0imGFNlv1ff+QvWpd00MKSMxNm1jwqV43ixWiujS4Ld7zlP+XRgxwr5r2wdfijJWNE9hVDIVlpo8
6OqLlOn2XFPPYPt3linBzpNKtVcp1k6fQWOHS236Stgtqb/KxXH8XteNfJTu/MZZN7FhZD561Lo3
0027R/rtWs4Gktz/bSvAE6b5hXwdMky+r2zx916MoqNFDDh2+yATuUIxNRJrMgaWc91RjQZGM0A9
hLXUZWAySETEjgZdjbLF0SKM3AO9fwn9J+WGGeYNTMBRfxLBQkSMuKBnYmU4P+ofsjLCKBxy56wC
EwTkF5i/rwpKi4vDBypT3iMiSQ/GT3tHpGNJsI6KTI0TrJrm4uChOz5VCgz/8apwM4B5voygj+Jm
PLZz9nKCcjZjqpWwSC+iMOpSCXc7yu7xhCTY2+1wjX7VVQ5tN8rsg6WkDs9LALwodZhPOmP+w89r
g1Kof+fR/EXhauLVsfMPdNl6DlVns0n3YpFrkQNePsRS593kCLAIDGliGE6yPwAq3NA0IVQ++yjb
CfaegnoNn+vWa3fpJRLjm8wVdSOhzM5T89ZGymBjF4SM8KEaolxJHzzxxjq3fp4QDznuLgh0VWKn
aeCuxlWQkabF97ASB1Mxl4yDiCdyxvy+0fSganZLfDyd3buOn4CpXGg0Wg/X0E816TinozNuY4iZ
3R1j7LmMq6UsE+7+e8cdScYgY6A69uk2IX0vlFYgpCLlmsBG6+S2WSiHGMjCmHwyMrxs/8k/HNve
3KEBvHYzf5pb/Yq0aK4imjMJu92gP3galcASevJY7Qp9iEd8DqPr1RP3FHVjZ2FzmIL9OXh/GRRY
nj6jVB2Utcl3b/JISlmedXhJSN6vNcIM6KB3WGz3qoL6sfv8VEoCZdRE9AdSap1fkiaOBqtmrEWf
Q0/hJ/1FvIu7sKO/IYD9aTMdvY94XH/PpJhrmccmMJ5bsj5Jy69P4iUyo1v8qmtIMONiHpndS/Yn
RILc8w0yQXNdEdFw5s2CNLvUkl4DLEk18Hku6l8Y5pbzBLwE3AK0gzxcUnw3AxpwmMpGZo7g7GGR
TCCAEuk8/N87ct3vHi8hmrGpW4ARwa1ueV4mNF0nGhR9Jo2e2OAgo0R8xCuuHa5Y7egsaEuYZL6T
oIwqkIbPMrfcIky6tJEjUXLG/aG2juvI4uCmXBKJG4WblOgz+j7PffxhtCrmi/l0/zzbfc/m0p1F
31zmOWxgfuzauFvMmAXgUtn6eYj82uErRmP5exkRCRJmcWGjDdP2CcmjKKdbQiJ/8tk5IEDh9qXV
Ty0eHcgzExBHfTtQiMztU8IR7oYrQPocHAc93msAhQr8OBUR5vMxpEH11nUgPAz/pBX1lZHTtKPg
ozt8XMGu9UEMW5BlmAiIoA8jJ9uWUe63TRgQg1DZbyeMljUCYa5X2efUHFAwlIicNV3zOpRe4hvE
JG2Ew4A4bmM3MPPzbi9dbdUQ5GIdF3LrjiZ/sK1W9QDVQtkSx1N18x9HHCu2qq4m4NJyx3SviXQL
euVm3vgyXuPrnIVSb4yENhQ6SpebgBTl/XnK1FTiaKsFk1zjiwUsgF+exjAKvNtL6PJPJ5lX3yQg
a1Zeb6eg03z9QuP/2L6G9hi2pSwYhsDxdzKiLelzbkVgv7MJuwR0MHiLe/dEXnB63+i6nWB/0OO+
idpprFUY/eF9BJtlH2hD9ccrpBNL/RRF1zM7Ck+6YiqkX+JTKTlriW50/0N1hwNDNIyEU3d/oi0a
pkgVRLnKoZiDmt5GXWSVvtY+4HadhZOPyBf0QwW5sM5aLiB5TuELS6QnGqUG6GTSlVPlkPPIzqII
50Q4KX/HzL54Ri3IhDCbDDjqEyC1ZCi/WjjJdUioS9qsLAsLYMgB+6ys4oTB/guMY0tycOv0enld
5IvHIX3cQfxyZsoWTLUTj6/SLAEb/IIcBvqn7bgarCiGxoraxUV+kNgOel5+Pe3SbHTTE8O6kewt
H94foDmamZ9eBk41oz1qXsZYYhx/KxZqhakbyrpCTA2+MjtFjyOdpM/h5or88/RkUWY2MDYHhZgq
OqvumMvZUiKgdhQC3t3tKtCA+YMSTZyMxqQRprPTnOMyZQMGoNFxTXl03xBI9PFRltCNH/0aUbEK
cB1+6/vbYx9B4KnI3NAPBFs4iDokmRgESQLdgK4M90J3Gek7sdZT7nqFJz+TV5WRgqSKqwHP9Hr7
tmI8HZKF2OnfIh7Fy8H6rUmjJM6fbKF2ULU/sgdpl0BEP4ONz/O5FJfOkduZl8fx2Qsi4CYAENjP
gsGmnxDher7vfOSovEPtkmJzqPKf9f4vr09ZE0+ACxlWm3aJ23jVp9jU9VV2WCACdcPBqI9UKeq+
V3tvr0215JCbE4iMQXaLaQew3kN1WfTpaI6GfRsSzEvWkr/IBDu2KYzZ4kp2U5a5TUkQerhaDjPv
F3kbg9y46XWJj4NwfhaLgyo9PFiRU16f54se2EHP0SxtNitsGsp6tqcQ/y+kNPXtIfGj/FhvWrsP
xVCJeBR9a/NOiTb2hRSYgmwrNfR0UUS3mbpyWrtFXT8ixudLRdPcfDGcNZ8NO3/13XSXeY2nOOhB
a8PgSLr69431YtcyCmKlfO3PA/8++HgCZcoFSKxFx5/nHErXQK7NUkFh4yWyaKdTQtvXbTaTPbz7
b8UkJIx9Puz6FAa4n4yhcTAulsjgAHXLbmZ8ptwr/qo5AI49bnAvpxf87M1LcjVB6js3jU0H/jZu
f+H4hntux8Zciuyg398cuzph64tGdu+Am2YysYQ5skB5AeuqucOet1mfJo9MVO8FXWnQfjRzj8R6
nOhZqoKZKjVj1KA0duYnmi81bjkqsV5p/8y//oatJ5C+DZSJDcXdylypzlYSLW5eFIixkVIZTY4C
vJ6W5HhTSgGGnGEriGLIueDDETFHjVGHbcUT3R6Ctvqw0oBmakhLwklPNXhyHRNxjQmaXibVG2gY
tqSqkFirNxPIQ5A+KY9diiukvyjWkgAMbJyfPZRXPyNaVACeAAHs+OtmbkPCNGwKFh8+cugbVs+9
8u3WamrTVclURPiM1jBizV4wj68pT7aJMTv9dnz/bGiNBj7UCE3JqZwqYwpRhIFb1Jj0bWf8xltY
i7gV0WgCDmmi7Sbhwa/y92WZcWuTCmgImD7SRqnJusPtnG1sVYC2J1Bm7cs3T/sL2vo2xy8jodvf
cIEKoN8Qov7HoCijj4FDvXqM1tmO5YRjusxHGhKavszqHXVQzf9N0bH/socfnjZwmYK03YFcpoYd
eiHkKxeRjBwfmzeu5tYGsKxlUvEGHueuCR+EC8/kMcRQaxff8Fc706MIVscZ8G2sP4d5a0lICYC3
X6BgIJU4kQ22saN1Nh80Yg1MumxHF1vGulrquUl1RZnVfmQgDc9M4wUbQioTKAb8EkKVNtiRkaTF
hoIzs+kTcjkz49XL5N2aKQ5OzMqNKjZcO79LvH908VAGlpkAgEIWi2uXwOLLICVYja+yKWKYaEM4
kM5HmHn3eyKMfv4mPSHeeKjjhttjUki2w/iuThQLAC5k9O03d3q058nONdEqjiHA9RZIzM1x3Rqn
Mj9yPsNYf9CRTzO0/dDY+Ge/31qfGWO3rYoxkbMgw00ZuwsMwMLV9t6q9rg9iSj66lK2F0uwu4/G
nEOudLPPInLbU8c4nzZVhtnMJwuG11Emc2T2cXlkaiVp/FPAAWzrOuAzEmP3lKw54YlZ7pORLS9R
XQhWEFIqJ5gL4DtaW2A/fEemUmXsWhYGkaB9epgpJ6gmkaN3pRiPvvIym1v3PDEIYnBFteu5qo3Q
EBV3nhxKo9TUOSmWVy1qfEcjgL25KF7falEhDdRft3pe8tXZ52ld4mP5WNsQEz2j6PO+NhOAw2U+
5LYjk1bYFN36EGQ5bJUJ02tkSnfXXt7nEidah3kk9eRGnkgDBcvFmIpogmCs8jBj9RzUi/UF3ytW
HDHBuX756zf++teOV19bp7wy57vCc95XOM/70+QNOnoWupeYWC7ONunq7eD7DPyJCj+PsRJpQAZo
lP63Vn+yjmJemiq5FrNFjHsZhPFIbgeh40K9IN4iUh5kYNsyyvXdxsLyN4O9+3ApnEWy69uEIIRq
q7gqfCVvWEFsh9yQQdmBZft1D+wn5XxRDUPO2U8m8m7XXkUqUIllJdEvRH4pi8PGpYdDTEDiXvqq
uQi8w/rck2LisgWQNXdf/50KYttt7pqGNNlruNtWqmFwrUmLyKFmos0rQe94WjjqJBuBUlshHagL
KUzJBPANQuvYPq4yNV7v8wDHfHNyMbHSF7RvdfJLhfSE9zeO+itB+NyaFGgzPnWzAa0rpHw/7+Yq
y3olkkXdIcoAwBbAbeP8ghxjtEFVBwfUcV2+2FTcuzZf7iDaqizdAGfrMWdjJm2+mEUG/nlOxCq5
rgk0DH+bX1YzF5ziBbvF/jp2ZMIfGxwNzfNfyRXwuwPHiZD+3KkG0g/1gcc9mfeSRmSgz59w1eSK
XQSTbmvFY5NSiJdcv1Y/APim5AUdnn0yq/AKGEnHzELCN5SjM9/e+lao3v6jRDF+P1473dnd/rag
UzXZfsRdXOQ3X312Ut0Tk5B/0Mg3g95uF4g7RXfmyfQzx3xOvkFkCjj+BWXlcBf6GRUu5CCWDiVg
FhunodMj9kAdwU27kRxd3LvxuAOTJ53k3YnQvlax7OazP0l9VidadqxZgONsVFTJIcwUXSdSB7vh
E0Xy6jmCI/hIyIIeySqnRMBeAQL0/rNQecGdIdsfWn/SjXru/VI3FuNIl8ZO7XpLQpzUxUwW27nM
0jdPLybyFGduxF8bhkW1I1WHlJ7RBbJ9rcyBpoKw31sc1nA/EdZeEJR9v2ffLTVXaCDojtVU64le
A58B5wcl24u2oqa+3NlZBaLQiZfhDpZGzwGAciLXUGkRv5YVTPmhYC1Tv5Ghcjzyl8UAPo0r2n3S
D7mS7r45rhNtDxyVRH+N3BJhQoDPIT+9Xjwn8E6lllkFzwpxH7YWrWNHwqMAnuFAoC34qlSos9JC
2gIVO3UHfUqJvhTkl2U0sPvXnBV1MX1+0Vu//LWN/Ke0HEh9M/YRzZp8TGS427jof5eJ3oMu/9FY
gmHVXT81Dye+43UsWriVOYa7W1q8iW4M8gQl1auvbm9LdCdx5uYARqZ9wCsqINfW0cew0JQVtzAq
1dMPNeoSQTL8ObqNEtqIRmQNnKJ2tD0dUvP1Z1KhuETfWWUj2vr8Adp2iMsTXGxUgLS1dCrJeTuf
v1ruq9bJq3m2hanbtaeMEGrMH8bGZXEGVra8EFtpOcPW/l9qSqPJFaC7UQk94hR1aaabvbt8Hzvf
3cRPqgS+C4arKwpudQrnUJ4zR8C45VbYS7IoevopqVsmN5o96uhbg5RybWHXZljWTCSwaiyfpP/o
daYuxqbs7clVWuFtrlbmbkN2AubctDwvs4lNWE48ZtxfhZFGpfSayYBIvEvmVnhRBl2W2FU2itqL
q7ieaf89D5a98+sL1j8hyUTBoJSq97pTvmBSvl3LH20j5wQCCqnq3KIFrFIKphEoYei/Dyl8qGN4
1UEjxwm8iwnJmv4jnltmkmX5QA7P3OySM4/9AV49Ea1tfmWnWmrigTnxV5WFmdxt7pujA1ijvuDL
XLRHZlErkeBMDdRnEzC7SJk0MMvt/wqYzfgKLGvukB6DkVP4XMdJGsX5GebXOA2TcE6qrjafH029
H8gEl0qx99Rl6QiF+K8aHlvt1N8daztIuu+ldpeXUtW5Yuo+FFIYzfgzHk3RPpE14dJeJ/9aeDev
muerM4UWwmVLVYqC12kGBWtV44KlDSn4gn+xYEhIbj5ccnffGQMD8qLaJYLzHMhlXSU4EztBahM3
Ef/ZoZufv6VdAW3iycFB8bPMaCigQu/aSBDvPj2kZTkHvJRbAou6FCL4yyIDuP/VPN9Juklg4X7i
BhmPTg5ONK65xl2KYtSgGtdyhkngqRXl1pAHlNIjV8cdTpei761MN0kwMugyUO6w/MtZMUHxP/Ng
VJBQankNM/T3kNr2G0B8zWcmN0X3N7p6xc6kYlsZyc8fwQNAjIVoafLibmCd9K4+bmhY+Ew6/FsC
8KIc9+8q9Je1mFunW9gW63WuPyXfgzFzI31yaN58th49bzBLS3Tu1Vly7OppwV2s21M0XBT9DYul
sq9FBTTC4GW5IgY0Kf0WaVJTRMaQYUFtfdQzV5FQZbl8lQdUmwQ7+PKIzvZOdm5856jd061yqjym
t1zvpg0/uht0swSEkKcXxP4kdthmHQsS4v8cH0gP6O26bk/UIlFFuEseyzGS+SGCgF9ZFhrAz8Wb
ZgnPN+Gy4K9MLEkVJXTMc84n/U5TKxnxFfOkxp1hkE2ouW8r/IZmJnxIudh0d2RolsmDJHa27QlI
9ZatcE+0QfJHwAsxT8e0kB5cbzBnInkJyjryY+IblFQQizxutydPKVwpyWCOqD9rOnLNBiGIyiLI
4OA5jaY2ddLNrz5LOsxUrY71+jrDSW8I8p29wm02Ea/95xGaxAiD1m1HhUABzBJptohw9nD73AIs
VYydzgMpiPZ5IIF0C9oxyqswkRPDH989L9CHvuPExCplB3d3iLVkvBqiQvijVvXiZIDUb0r96WLk
vLnLH7ES9ejFLntKBc1F0zviVlc26DUKxH16my2TKVoccxGU76MT0sAkVMCXsqTAxP3VrkcMBmO/
F9AFRV36xK7qwdbHYsHetpfOEy+KGyuWiXbLqJ+aRaVIfLQYXoH38vD9izbi4F6GdWdExg+Qw8p7
nnA4nWHFIcr2vF/xCH+bGkahPaYE0G7PZWBaLNjt0yP2JEDsUwVnBfgr2l9iP+uaSizxKQb/NZri
dyz/DArmrcJ8lDLIiEvwwi0ehp+FrE/GXlUYv0LQmEFXBRRE/NNzKx/jInQU/+ltyeVHx6YWiA98
NRkm+7PikO1+xbYzlQ4kEnD1+ml1QmPT5XREdsUtffpJhAnt21rLh98xtC+HrTKErGSnAr4QR/kL
mgBj7RbMzMXE1gWBkcbR6J0O7nmKHyV/TVIQIAO1gaChU7aJammXTQppaxfBD8uCPCPacgs1Meqx
o8Yk3OKQNM39D7L/UF9OQf+EEbD/uuRr5GVMmkoHEtE2blz7YDpBYKF48Hs/zHYBhQiTiam0+NhJ
3S0Q9d0My74RrpCVcuOtiAPS2d69GIrDyj4FYSC2+aH+x5xTTMdLArlOfLYenWYJvJJjWyqXGs4w
3+m4os/YtUO4gmFjWyr/QwlxwcUwBJZvXPYkXjiyTwpJDKQuClEjW2jfPyNo+D0vQLXztOPulFBv
/uujtyZnHGFVNIIKhGIKBhA70gOq/XXwRyVG5VtkJVPiwi23NQKVpxL+kHTz3HoCcay22cl4rh1L
GsOQqc+0qq6j64jB9eLsHB01FA3CvsN8k7+dU2XbtMPXVIEzppVUgNnnQ4TTICXqIQ7OUGwFepAP
3J4jmIRap0qNEo74uCwIhSmMDVxxMTovYrvwiIys7VVyj5rpjpZnetUm0SQLrHt0/5ZJORkt4jAb
46mD3cX5HCV+WtuoOVUIM27uX7kK5rrhyLQRkTei2izYbmS7ZGpwv+c8A2tAxArPNNDKwQPjl4fG
/qHaU3UtVG0A+zjRmR/z8RWGCQvRhv2Jx9gK4M12KFUgxSZ8YW1evBvx8x5dlI9/sHzVy6xnZYmT
98Z9dnVXAWs3YW2KioXkeDN90nMbfZ4cdLsR9eirzR9D1u2h7Rh0I+Kj5aHqL3hFHz3wslILPf4R
CYpraNFouDRGTEgB0c70eUNt1D5j0LBLZqGhcEWEGZAzrdPHszvHqopD6e++mfmzNCSLJE2YEVyw
Mxr0F4Mtrx6lnSvIPWFJ6kz1IPfotMT+nIVIWE1ZQqaVcoqMscPayDuKI1HwtYecbNpi5SjPSDlO
pfFJb78pbB5ZPQrhcpeGDnGLiXcJPFgIkV/Ob4DAoyMpy2dACSLnAoFZNBV+0YqbQgYeawk33JL5
iL7LUV1HBVSzxF0b0QhC1/ZKnvudFBfwhMICrcgr0QAb+gwQzIlHA1YKARS/M/hPpBkAh3n9rxBp
vONoIKPme4vLhKQySQ2IyRV1hCrJrrRO2kSZnM8WWW6NfCU7RNc8FS00QTnJ5PfV6vAiezmzZchD
LYs3mN5KL37EjSHIdfaNiBwRR31/v4fI7fS5mZyLibBBikYD2I3FjxbsCgRB7y6PU4c5B9OZay3U
apMSgY/nf2bVTbJ4ZzDfxkNE+xgeNtoHWX0aj3n4j9plL9S9wFn0vmpyh+GFW+5p1BBSHgEgHRIO
HAH9tVoimGvbp9WdPKvRKTpdqoLB/cbn6XlqbCi3J/7wPQ6RO1aEtgiNW/wAdXATT4xwQp+SMHh4
1VfzSoRYi2khQNr6Dib2rmfQbeUFU81Facu1U1fqpjb1iUp7XBtQ5Uh6FdHfDHK2IZ2rnq1pxJ16
X3hZwb0bmtiiGRGdLRNYaWJMAYBxJ21xJb8/dquAGk51S5lcVxXwc+ZqfVhHbMNJSqkBepU9FDa1
5H7bu+ZUCg6e7Q0NmS1eIiH1f8hcO5DBthirgpX+tA3TIYxJCjMVWulftQHgFXqqZomRXseYn9hL
apBVVyK5gzLu1z/5fEDFSMETZ80xhWcvqOSSPK6iodKjomIx1/Q2nFvezyuPX/R2cL8G9ACAfXZp
qJAFnFA/G5TMCoCNyVgi12fwMlKRaksBPmdHkcPs2ZHqHIPJ9Aa167senWLTZapw/iMzrrXHwuuI
WP1bq5rJr18r+nD9lHxTPKujEAQXpSaw6M2wCnxH427eGjOZpSHEOGHcldV1W/udCG8a8XrlMZLI
Y3EjulHYjryumE1XavCwt573s8hYixvWYIFLWuo09UFsZgxDAi/8sLCSkFObnjeW9z0OHEuysrzE
YZ9bfC861jYtcK3x2QbGjhwqBB3v6pxpott+pYuGHNzjf+3G2rJ3R5tve5tJ5oYU8cK284o4mpff
v1qwPAN6w+MStREtdfa5z6uSgJfPS41ZiI6XN/6z9jHBy0M68bK2zhBtsWAYqEXpubrFA7xbsDeS
vGfyagWm2xlXfB3WNDPrOBpkIsGFXTs5MbixtBMmtcQZ16hl4nKP27uNe7RTMPtMQuY4OHn1npvc
/2gM7pJlGGAUsIfoRoHt2ApX7odQa0wDUrl/7P7B8RBHr/uJby2FS69AtvvybFbexIo+S37va1GT
XCNs4gERRM/kQ6WVa0CSv5QM1SsVf9jYGzyucE0BXNmiL4CLxeEC0OEEbYwmOtcfH2eQuB4VEu9/
oDPVE2L3ws/xZAYZUypar0y5vvzSNJNJz6ITm+HE2VMEG1uMLomfCUL1Dw4TEJQk0WJ1fG/lZ7I1
DdXEynllinPzmzXepXMvDyiPo0Ni6UcJAOW1RrvzzPAUccuVeMrjdgocBZJXQnXf8rr8zR9k7JUX
k4v2adFcvdM5PtOnQiKfLMj86DX6nYw0JNXclMvEw7MJmKS5EimyqFOLT/vDUCsNLegxDiW8656G
rHPc7cMaMQR0dtkJNgwrx63IIO/S7xNCe6+LqBg0G1FsSBRSJQh1GB/CRsw45XYjqlzPj1HjT27l
tP/Qabo7duHsUacUPURgqqNQDkC6Uv5o8cjhPrblsREDGx/Qh/4DvJe8pMisOm8fsIkGWJ3uWzEO
ioSvQ0isf/bXCzPMLDqLK16Ru0ApxUSq3AGfXFBhJFYbtZ+6FVKLdvOy05N5jHPIeywAf3qNESJ/
StpxRgd7ZaJvUPPAR4q9c2YipUiUcyFYa7MYFgSxtDzdqvBugDBCLkfH8lyc+vGP4nqKAlKPL5Hn
TFwbs5Ek7mUCx281AGvJNPzT38xFT/mkqik3sk9wbYL24glchS6/cBf8RhsBci/GsR7orw6SD7TO
vTyzgPgsC55OKV9TYTv3qVsoBXAIPj1gNcSFacuK/O8zRqK2UFygl74JQQXm43u36F2RA+WqRw5z
8b4oeLtpKxTCp6o5X100WgaiGrHdbWPF8Sc2lt9B4Z2fJlr8DkrrF1FjgMg8hnVzyuR4TLr/NKX+
CRSj474QzU3ju71hccUEneNUxeU7o5Ub6TWMaROuYE3Wyc5E8TvaLpnkZEeeIJW90FaZ/hkpFe9A
9/CoMik7JSn+uoeY75PDrycC/H+s80xYYJiNi1misSs4NNUTtqLzzYJ/Sh61iH1HHWlHqf2PcTNU
gO/ndM3Guqri51qDFYJvUIMYPXYjKtrXUN7i7J0GuwjorBNAm9xQnaRLiuLmXuWii/Jmx0Th/QVT
GjPZJgUq7cjysjmD3Bt6084Ww1Q88Y6mdDCpO8tWW0lmerl2Lh4eAzFKuBOR0lyzH7HzYbgjzYnP
aleH28EEQCXwcEJWlSvkEkFK10WhhxLFy6E8R8SSeuhgIPayUQqTiy7GDVLC+LVoTzJpJ/vwjT62
vVawp0p0lcBN8GngGNTeuen68b3tU5F2gqCjZDj9EHnFJOS2fapwh5yDe/PPY/VqQAGvcQ3K18/D
oI3ksj+wCF7nQfNyJG9LHqJE8NdKKc6UqUDezzSqBCIQH+/pDFUBioOtWYDJ6GEIwwBZsBJ3hJ3S
dneFjFeoAhhLsdE9P07KRgWm3ND+NVhWBqwuOjHLqkb+9OmWYJ6I7eGAlXy7BrSgQw1w4I//WxQf
WF441w148bkzXXjoS39ug1ZmCVrYlJ6p82P9dadhapoeFXn1bQhSe3BWb9VLDHE5vI6BY/GUla/h
LLP4jYyGig2UOHSGXYWzaaXvchVcPCVQwz8h0NVETNBWqk8twKw91pbuNkQ/bO4hLr6P6TnjzWVa
UZkbsdvH5gKChb/1E1VmbYTuZtGVurC5RyttQ5YwLy2by5ImBqNqLuD/RyfA5rjMYmUL5cE9BWgu
uMmNsW1Rq81HjpGxvcet8BhXdGeg3iQaUz/HnHQ8pZXWnH0xoyMrZXl3iVdlyvhMcPfPfH2O7RVu
X0sS353rKHhyDhcWdFF9TIp0XzDy3uf1G4+ZKSXIf1itJoTEFzC0Uv26xXbNT8Sm+/LivZObxjum
fiUK/7opXS7NDRpXdsCvFPdyqcDlTRaVzls+j2lbf/Y2T2BzQfasWmrwq7qe6tgbXOYUSZEhyaR+
uVdQqSlmxxmQ1X8fpYRTrIDeiEbtvuJJReODZXELuJPj0tUk2gVfqEKglk03+MLCge9qqvgQvTPG
xEuTBtc7dC5Qam4qY9jDk9ER8lcDw+TbsfIN3BtsBm7WhZfrqOIEo63IhEe69U73yCnFhvppsZBG
G+bBwf2ujYkcWzrOv7mqsNBYlA+ApZoTJMV2qXIY1Qe35FcrWJm1S4i5iJ4Wp1CsukExtSlGfXDD
9WRqDpXRRC0EkjaC0yNE8xr4lapTfAZcrGZJ9gLtbzy+1FbZzwKQZYZx3laWznt/tbYSAKRmcUVi
5M7jQTVq9TMep0N/IDBifbUPkuxYZQDs6i6o4iYZXi5ua1CPgN6e8mVMwCheOA36a1NOyEL69NGt
9uXzal+gj7zMnJ9OcPDQV/VoNfi0/YZ4bgOTsbvUUUyLuIl2QimWfHjnOx4EGuUe3GoYlIoOiVDU
5dfWNKnHt8wmx6QPPWC+Ouw+oaDy1+KtJ/9Y9IbbHCI2om2fl3QEYDbPV+YDIduoMCGwk5Yluw58
/X6TZWk5QCXB5HIBQPV80C3bhrXIlVfYsGnG82cwYqHpBnumUGP2w2sP6yZc1ZpP0ABpNIG92TCf
rm0/SHeIsQpmTaIyg2HL5OLx12p5Ne1ouu6aMuW9PLxYkPp6UFrL26hZuvP1kQubdaHdK+ZMMG2t
uUG7U3dzLhJ/Rzf3JK82spd6cEzb9wMCz20rPDEhSwNphVST4g44bU03WU5LJxoGq9yLtbfkfav8
nghobelMKuGHgOElg/mlB83LfngDPnZy5IOKmH+J/I9fbppOpswVt2t0Itu0bXbYpdqqiFeuw6ro
Yw/U553WhgAkjguUAzxGMQBUlp3Xbq7cvkwdN2b4Vd9nTE2VLCqSnd7KBeW+0mjEWmbU6rriDNc0
ablrbeHxBM40fFR/MaRGPGJdp3PHYi1CWEbisY8BvkVH0SiDZxlmSrz8bPPHfcGWrrhTMosSaDjE
XdcxKPhjGl1wdXdJhp1+t6XFGhadfxUuuv6oCigGadRnD1SxWvjPj82eR/0lr6d94SmcWCU2Q+wk
Zb8bMzN6SL9/kQCpIs/aJn1zVDEKevB3yvajgFHYpKOaYXXsDVUHfs9ayPshw7K9MRG0by9CZjnK
lFaYnJv4cUFDAuDNXXNnGN3d5Nc/vV+8lxWYjLgLLqdqDcO5xds1/tj4KTO++Dtrgdgq8+Ia07jx
H1Z4rn5GAFIYztLRJmJQRNqmP7pOxtCOJpVTx1xe7VYa8t7nKQ02zg/mbjc1W5jyl8BUfuAirX2X
4J//7tBHU6BXhWCDJhsg3NTYo9Z+eI0f4e9fIWZaR5mqm/RtREr542Zq0EIQJa7RfzVpTZRG6Q6Z
NAeSUqK7zdoVy0viaIWReZz4NO6v90J9CJsEANrsBA7wzJu0G98IgMZDqv9cluvgO4xtJCPHGqbc
OYfB+pjdk0SExpn9jlhcD/Ep6E/ZPY2DQEJgUBHG28JVFQjlGWmHkP2Tqb07QERPlLpXAT2ZNDGX
7ZIhX+8YtX5Q8GIB4+rmD6pDbXPy0MBOEr10zkvvs6IoAtfNjvULtXbLfEPRngLWdSuJHnshhPas
HO7jPIxGNsI5Uw3Eu0qlSANNsYgJCxsTOw29d/OUhqWyHKPOqz1ZXi7LWXCM0CbwJ9nC1T9Y9wyr
ym17MVTp3jn1KyGKtZFOtHe/jX9gk/3B4StndEspGb5qFKh0RwKW5Wiy/QE0mEBSXXfTpoh5teyj
pM9FtN2G5INkzM2qJoo/9OD2coQOtIYPyZSyiejGdInz+oG188uA+csfvyKG+Vh05OIdD/G1VFHi
RxPC4WkF5FeMwjIs71zxQX90xNbSlR+8dLDeogZDyRmkqS+uqwFZQr4pYVFFmLcRtNtyn95Eq3f+
hcislrVdqb8kxvUqKfqVvLEuFGsg7nboHrRDN6dC+jiqIt/swtoabHtetoEIFxt0rR0H9CWKbkEB
jruQc7InYvoIzorPHgjpsWdhsUQqNtEOfoAnq0RVYpdSvnqPB2hpI5l1nLQXo8Bt6r8rXEIYYdmu
YuP9NwipL9+Qvbct7br+8o5LEhznvh1zczoCNtzHOptEUU+EUaqrVszOnrwTqPeBu/+SCQ3dXHSr
Ec1qDkNAJg6BopjcX4sYnwODey/gdkCsmE+o5U3oWxRtYZd5kky3ksw13y9fzx3XocGzvjXtbhBu
+Rjuop5zw6rCLpi43U7xMVFAPpdCIvnuPH/blYgyGbTmMKC/HJHjQE0CixnIz9WjVPzxQtvfWZdR
hfTlVyFtIp3UT3NqoBvvt4wfH4tqikZQNvaPLKUMVGHlSp4kqVnRAOiq4D0u+Q72muYfYdovIz8E
i4SsoYR48GafbxePxnOT794kVop5OQ37uyeZwRxSZozeg7GduFVsI2uI9J/x8zhdQQXRB98OxPQV
nsooVL+mISJeznULIiP2YbeuUnvvxmi4puDg2KMa1NLakFh+1WNTTIcObFZKOD2SP4FouKnltW1S
tEAoD6Z2SKJdi/PKlHYohGlt/K/cgFRlImQ7y5rOkPxdw72PtBWLtZ7QFeJDk3fvHYvWgqCkrdE3
2exBUpkNAxJpYddxsbKxo+D7d84l9X5zYmshhvgmAS15O+BqO1OENg86kv6CF0m3Zp5fAcr6Bjwk
aB5aDv71yPKbJIzlF8dkfIXmD1R/htKwT/21IU7DCuuViDE8tJ9vXF8t3T4NsEQ87mLJWcX+QFFa
lwuUVrQzBZWcbrCZkcriRKP3aJFQmHzv42Sos/yIsLSespcXXPrd+8Ep0s04CvglRxqvPzEqvJm6
RjLC0MJvEbUReVYgX2tcabBAMJWrqbAMqZQbVT/s776DFIxFcM07s8j2haPzKCJkUnfFn1VM2Z7u
16d+OvUKjbDiefo7nYCykzG8iRfl5mAfjsM1X8M50R1L4UfQiJTVoH7aIXo46u84XUIRD+W6dP2Y
lnNc6L6WeAugW+FIpqwINjxVI0zsDQzp0M0oGkJtmCX/z13i5ZyA7FYOxF2HckTIceOQEyrb+jk0
DxQMxXL1bgud64kjaJ3vPcq6Yz9YDUTlhsLFfVAJhSqbF7pmSDoXHSft5qMyCZwRC/S5E8oZIF8R
Ja+icuRd9nA5i1o8JGQqV8j/cdGZwUFfY/mUGk+lMD+dxNrrrfT2RbqjFGm7SXJpE+sNazAJI4t/
iWgupV2PGvWogL7xMJYoqS2RSuaanwzPBoDNrZ090lb1CMjaK7JtfWLHjGCxUmlIFvDb9i92/Ba/
Cnr+/+YVp7djT0JuotjIcaFOJNis9jAbK7+seXEA7DC81hht5EUXrRxKW4Rt3MYYh+X8bSKlCKZp
Oc3AVpFNqd256E48eOy4qzJprl8yDJlQSf/x+3cjAkv1CJ/1s9x0XlS27xyC+z/UsTRx4OwYIOBS
uPNTdL2Z8ainy7pGee2qNZ2/px5Q/DYd3rGOsa0eFNMlz2z+YzNeHDul2HjK6J3oZssnFp8eRATo
rqS/aJUMphPLXV4F1xqTK++/KetODnRrN4FZ56j7EmmO+QkD7gH4vePnVML6V0cdvZ7YxH5mxazu
im9B8QuJM8MTCx7zw6Z+SrnJ1SPk4gMKI9z37RiMrK1TpI0pkrw3snCfFTrtGz32LSnBDUUuzZSb
ibbaW6led4TyF62LqcF5qHGCeNnbTKU8Ffb6xZw+qv8yNjFyCUFaRsrj5+pQnA7LKJ6oAyLhH8wk
uQ9PvXOr6RUFqW05uQOpOp5XrbGlEZ8scqFMyX1ybuF6JfAUkubcGfIl3xz9xZe94yt5AiUNi9iV
VIG+iK8a7usL8Hki2uAuI2nXPtAEmLz2WlYlhX97UZRFGfroM2gA6aXMLyzoLZyVWnaX6JtBpf9g
pWz6tKGQaX4bEXDXiQ/bL5SFp5bSfByMaE/70sPrDjFMsRzfIYJX8K/0GaHtYBLfsihSr6kYtUJh
ABFHlKocJZzbRbmRoXLIeNdHhwqmNTQAoJlsZUBb0C4ynOfoVpPatUsaYgg7Ei2JC+bWiB/oQAdR
GBJgIehHkhL0SoovdAA+th7uFAwCjmtcDDD3FyJyS/woL+3k4+ERFRoT4+BCPqq62ioGPY4VFh5q
1msC1vKJpgcA7h6soZSamvsiiBDOARQYrhL3rJ//7Ig922X3+b6fLS5WqfQlBYvJ1pIa2f3iTk6R
7zabXWDcnxJYlXTq1B016YpB2zGzE9b+Lw+g7KE2HViYUSjPbVF5SWUzStOyDhnVSunsZqMda3P4
8QRWS1fpGo4w/snsrQF5f0MZmQ/6LrFquXhZkCKdthoG4pgfHT01YHpDhc3brmKe5AwmjSzilE3z
HnkdsISj5qkJL3lzRbpqU3k3XPBIWL/tyRYlQfj4po5se15VOUDzX2NiEoT85qwDnvEEITYPQeab
Bvg+VW3ubqdG9qT+9LsIksF5iKqFl4+02e3lYSI9yFZWDftaKSMFUGBaPeyUpZPneAwR/sBfvaMD
Uz0M3P+QrXU4bbyO6g7Vi+s/1GwGXilkw2ZBMQSEwxsyP5k0zvjbkjVbaM96knea1wvcqC3Uvtp2
Bi0/KKkE/J3fbnzacljnGJ/wck4cgjGgl0t+PKGWCmao08zsjbr8urlen+Go/10aqnOoL2mJXCjZ
FnLXe8JfuykdfXc0D3y2sZQaO+52MUomqREgp/skLMAvaOEsoaRSsZGl0gnLcFzn0jBsnlCb2z9r
X3lMx3B2fC5q/pYDZsVcCpjqku/sNRAPQE5J61+9asNpRKrU1Aw9ocwDDw85Oi/Qhk523kukB/qp
bBhc4S60cRxS6MV5kYO2E5FDaNW0ZDKdDbO4NJFeabu7uxZfItkrqrXeYDn8tSgL497oyKYwWblm
pmfkbj7he4A4ozQNFxkoEB5mupFpSzrC6ljkc3zHYXnUlNb5WERgHco2yZApgSt+5ohZwoWpKG1Q
lGiVUaUqWUYACDoPUyvvF0/Up8FKKDVa9PQp3Zjwk2Ft7+6imAoCO5TvorXhRgmsAekooDmeBBm8
aC94WQfzOx+roRdlrFEFyXSRXIjIhI//7s++kHCYYauHKbE0GQHsxVEpGXlZQZ8vknTt4e/dRg09
gNl1Qmlkk9JWomgmE184qmU/mb9/B2CUw+QC9rKh2/ZTxN6FcpiLRuy/qa5eb95kXP/0ngagEQw9
s2j71w+uaQEUbFzMwXzSGtCCiz5h3jCo11d1vZYptKiQSt5gKxIYBmsSbs6J76t8tIyRJ8QTNqq5
VoGIK6hVMjC/w48hPuY0+zkgOXmx+hadqYB+xT9hYcbU3BZfVcVnDuS1ibWFbfc6O2nDYqdfVq0I
RC1W0PjpCm713RDQ0f3/btDQachcl0vkWIavQd+3MriVvyhQwiKv58k22+aDysbR9L6yghQgeyxy
Trp4SYDhgyKdhMXlyQiWgJE4w0Os8qBC8CYOb1H53jyWhu2k0/x2bRPXVcZLJ3cfjGK72wH4aJtE
KLP3d+Oc5Krphpz7wd1FuWJiPv7BwJkCu9UVItcIwfhBEwgEUquSAZ5oZhcmKvT+GyRvJnHI9XPX
gvLj6X46JXWruKfv8X61L78s7qmEAcG2ffGFPorZGRER9le8PzhNucBWBWjW3CziDTjXjmLT7cJt
b5P6EPkuG9DbcZ2Zuq9lRMTDRTSiu9UW+b5jJRIXCi48dVP6UYng3CDp3xQfd2r5d3BBzJYxCa0G
w+Tj05BS1PLvWV9q2CpPh1jcWd8hXMb012NoEYjdKDX+0sbxSSJL4Dw944Y/9hAxJNpNKmDplIa5
NZP0lV0J/npa1TNG8XyFmGSGp+RAxUSnNTd505Au4rBhaAP2ezxSPogP3z0CZvu0KSpsE14bVsVt
jr9wKpuLYvSl4Rf08inqfuG/UpA5N/6T5l4G6Hz5TlCLgbpHhPW3VmfWXdUHN/gw/Kgw8K3a6t08
zq6pyO1yT7UIECEDUooE1fb4EFuqtniZq2TL1sWpm0mN3K9vOVS0wfrsqM9sSK1VbfrCs1vQWQwk
iPiwkAPb38X36enr6RZ9V2KmxK7+T2E6qsmfVgvP7jgXsLbOglE306WceFHTuPUnPtJrXnKs3aSj
jEoLIW25YaehmEUbH8LniJr2HJAnzqIxVbq9YKdO7ryEOCkqqZNG4tryfJvxLxGJpLxHQp/tzh8d
4m2WSc2mHGDzs1k5S6lDdkgOiJYpzwRbshaxWhh295Q0/b0vwzu0HKhs7Og+pr2G+JphEJ7x/iXz
nj0ODjaITnUugCwZg+KkKoauZjNMM/qyEwgLYvx1/YcMaDNH8zZYKzUQITGe2NqshlZAVZrCtReV
Ov2GzO2AulwpqHUmPujQLOlpQqlvHi11NukPkcuL9NEgGHDqvTGl+WgDHZRiaJR8gXQRV/xwnk3m
y6zMfpKmePJtTrX9RQKuScB3HVaIWUs9KpaPmOeTL+dC0KMkzMt/+Nw/ATc6l9nIUqs9R5dKx1dh
exzlDBMUVgusUJd8vjv4zMz8KSRbj7UN/TgDQLK506btfKYJlGHAJBdQEw3/we7IWJBFL8fPJFt8
5R5ti3GiN/H+uy1A0MbIXvIoU5Tx14VyKQ0aAzhNYC/dTSB2AEG6A7s2405XwjIXC/XJpxgo8IHY
VJRtwwA3D+dECFy3q0c4FeDiIHDAj1Sn8UhbJBDf0k6fiBfwCQsmG1gJsSByyzA7S0suukb0HxAK
XOAfhMpmrIJ+1FSCZ5GQnTaOrggtiUO5gnT6DxWLyyoj6yLBsS1VYL+tMDE2VCx/ByudBCk9aeDT
6e4olLo75d61yz7Yt2atYKADzfhI56H+y9QMiXe+fQq+Ss2ey80EO2D+fH77Qx4I9m6/cFM22Q/P
tcjG/V8/5J616tajdpwna+TxNmqyOqxb+jmJQgICQu/Ob9bhRRTJiUOjqei5MZS6rtdiMWrvocyS
6TwP4qfarH7oioUQ7v4zcnrLFrwgEVX5iT57rdvn06WyvCMri2GTJRZjCj2s1k3O4m6FH/FsNBvs
/uAYz16fgA5m+4KQEO+GPYPzTdj+KzJRLL9d1Ip53Bq5EJNEgM3g8vOd3Lmaz5AUgsc+3Ahm9igl
wkF0wHnch6FrkMoX3B3DSac7QB9+0KpzY9lEdy2YztYUjKBCC/Kq9DcfaCUTWQcbDsc6/6dZ1qTe
qmXsLrWiZaogjmnM45kFT5u7khoKMOChAV+wJB7E8hp+HmjtvmWyyBFELFCPFR8xsFFMEu+hluUt
pr++FyEY9F8tU23O4wgwKkPIgTmr831iV5xSum8hFD1Uwu1O+/XEGrrnjMAUROy1QjFiCmGZlHcO
XHnQYFFFLEZ8YcL+S2R2tzOqi06DykoV5eikSkhftd9o+sofVTdQFFRMeQBgHfyfoJE2IfUcT/QK
DAgMV0XUYdXCClM1uK4T7T9MebMCY9fCU5wgT+Kr68GQmn88BjujThdgnI1FSDtnBd2N4RcIU8oL
1ZPh/VATZqXwV6pP5HsKramLdobxTjtP82rKnH1dAWPZK6wfbL4u8H37evtdajc3DPSR9tQfBSke
X4olOdwzEazth82I5nLulC3/Y6KC8kvQ9DW1cAnRe6aLM7c9vI4Es6/CH5eKltH8atSiE0eHgDCZ
T+QtOAw2a4DAc9KPmfllmkMz06yhVWjKqZhupJ7LMNq07jJVbK497OaRovSW4S0+EwzCIBxZUmBJ
12S3d1e13GwTJiEV5hO9R+311f1SFmGgIbtMawRsgT9A9q3pxHWHwvcMEf3AzYHbWODYXX6oOJ18
5U6Wn4P45dL0GAVA6Y55hiMpV7wwnX5vPvXtcI8++UaGeYubc55eEN0V9B7fO+vGF34R3jeZPmHX
4PuJAVF81brzEFaJVWeJh4hwrMYJCuhD84ADVBQ7MGQL+EAjT/6YKEDBQb0rkAORURdmrs4uD7SA
74zFIUYJuxbQv4nVkEIdE5FmOa2dkG3FPPjkzb1vBGjr98WqIDkyOiFEk4Y3TRcHPf/5eFU3eTEE
qkwtr7rbXcYIjfzKmyrXlvzy4cMfWut/6oCR2ku9Q6cX0QGUOPYu2QTZ5YvmLL0b7mVoxkzo48Ic
tFKyctl3DVE8hdlBhXO452JQ7rdke0ssjIiV6oF4wsqtJAEdHNb8JAVCgzJMHCKjyFAJpo/kO7u8
5xhk2XIRco6l26C79en17BDhLNRlAw9agI1Fx1fLU1qHslLobQ76CGtmZdNLUV6/KsOHG83TCPHQ
hQkW733bC0Z6anhJZY3mngKLQdCEwJBm78mcUffeeFWCW6sNGHTqcnehG07hFYVW86VEe9Hb9lHD
RyF+6O4fGqbcLj8vt9jPzXdxS82PKttsdPIwwlKX/PHmJeAttbx8HUtegc2+124xd/OBtzJDQeDU
xHBbNFy9QjAaLyukgKYLdZ+YRU1okE5Cwz2yV260OFmGI9P1sCRjeSY820msFwNDqiM+h4XFiW2N
/IYygPEtGIEvdygMR+MwxOIOJeevLGotDhkAcv+LfR18OfCD53m1924zRAf1X/lEwqvvhNctZ4m1
0t2DLcxweC1w8VmzLz69ebEickaCxGDNkGPfZSXHX0/EwBCEDFTw06m81NMnrMqzJ0vlpOvDYu+P
uu/HbBqwAsyws93Ppd0/8p3rpZ3F2YL7Foh5DdfVOtnRw68J9cAKM0NhQZaUGeBmJ85nxnXqynvc
gXVE9x9Ry2ZHwdErlAkiyrRF29V6xo5xbTBjLLTn6bxdZbj0CPLgAXw+v1aW4BsTA+yy/N/g82ul
Y3y1o8euHozu5GuGiAkgpQMK9gpElBuJ39OEg+bssLAV0JwTLcGMWAKdPhPyS+NLjDz7FBnfnrxV
WvzLQGPQQ6zwApCWa/DPfVPFJfJxZLoUCH4oSmNYWUFNfsT+OWsokF1vYEV1XLb4w+VhjNNoz1E2
AwmVmN/XzOgl6y3o61gbMUt4KAF3k+UMkzQwEyTVjLtMeZHPFbIvyQ53HcGR0WRhtcwz0MXD7LoA
f5Txjlct568e3wD9JFkTFFq9Xwtox8yYgLaFID4pzSLsQASxKtMB9V5o8iuK90H16UkEC6VSXD92
MxPR0lXl/i2YyVO+/P6gNPTiwD43EWQThuLt8/Gp6tq+we3GpRflOCXTSz6I02ge2klZPtIemaD5
b5IBgNprchoVWcRgKpoKmNfo7pmW/jqxamDQNsztZ6zqb+97flU2+dlM2jhVXNjvTlkW84OLKp92
VVIMvLfG3QmwQTQoga/1DbOyANr843OibpZhc0G1OCVTZTl52aLMyRSBGeqyO6+ceLFAP4nKhfGm
iPyCgEEXpWgLmEx3MHi87Avq4uLkT6sFaJZwOSBoHP9Bpui6g81IUBQq0mZoHN+xxRmEcQYVaaOx
ItnMpk8txi7v8uIKV+w73GYtGPQ6O6eNj+4FZGCUb9PRf+R9aay7ZlUX9XuBFUPk0OiooXLTC5Xl
6Ya619g+P0slKg/o728vRCpIGU5dbAtweiMlhOGP/Swx/2OqRAvGKKn/yDHOVtiUv+XfM7AiMy9O
bJLvWULRRex4Afg/RER19CU5KKd3QNf3oJUHuhpTH3ohT7Ka1PHzxM1UO1XX/jf+9s7G/0HF8cgz
VVwpNHqSuvp8Wh0wAyLmCWTgHdKYhZmuLvy8sYVvj8RtmoIemr+lza/Zlm/ej/XiE2tCnIa7FWz3
lyi7Xk0GhESsOjaCGyFyZntRe5WuWvR1VBzIXeSrAeujf820TKSqy09/JBKsvouacDKqt8Ea6cOG
TDPxb9v2vpqwjVepNc539UXGrwW+XsA7kSguYIRhPEMnzWIeicvp5JLldJP+Q7LjREUSCpOUH6oV
HtxkvoNDxKSrouoUcz3FXZ8MHPh5WOiSf6SvTXay4Q5hiED1GC+u8YsQ7uTCFlis9gV3nlHLcJDe
PthH+Y3wn1y3BqVnEu5tNiQ19LNOd5jxORWjuhzf3WeDinNiUarPuq0sOJliGftvrndwZLLLAPoN
nfTgi8Bvdrx5/i3LxYaMV6nO5I+ssPb+HsZZuvlBOsRUo3X8offJtfv/ebxSpjOOSJ8Tu537cC1i
WMz2yaWv1YYd/LLVd43PVwE32f1PFoATt5eIsiGEL6op6FNPRpsDUf+1nfl4onA4fc/zYhyzsSy4
nfINwT584U0YoA2jbkJvvnCq88utHRmXcJiTMJBRW3tmncD+bgWf6FO/e/amtX8YGWZoEIosHus7
gQ+6uDm8P/EOCY0dukRk39O1qZWjIuZn+AJGsYADpjQCsGe2Df2yP+pVEtbG+6oyaQ9y8tHbqB+F
eSw0d19zqn7tJXpdPaxcYwLb4yzdTkRVt7f5V5Cgl5CFNslsz2RwmorlIA53ks2CI2Q3CxZSGym7
SaV+uyNBN+SdSR05ozqG2m9f/SucBug2dZOfcjnlS6911kYmBchzozpHetEmmR1upb4mnk6culOd
0xP6Z7iBgpitBx8z1/EhYFWlhyacQQQ5zmabW8PNItRQ1Qz8t5uNH847QVKMs+YtbJ7btQH8oIqp
PowqT++P9lxHspXECH4V+xlZxJBK2a4jE0h+ulZFnCQQHShSVF9Dw6eSKgmzu9eKFMkU38ifWmti
MQLuUCnlK75ES/C3X8x0VxrRLFKzpDUGkwxPUH2N07P4KU5mPWhKJE66ItaJoLTbb1tblt3H/taH
Nk2P+KlX3hthgp/x4ijcHxnVfjgz3yyK1DdPuBUN/tbLfgeDVIZMZWgj/ZLcmtMqdf3vSJ26Qv1U
oPTat5xB6PGKBtUlLm7JAlF2scjd+rrN+sfFcDsM+aPRtq/tW0bVZR8id30jkNYLD7SrBleWdOU2
K9t0aDzSrceS2kKFE0A6TZdHzQgciG+jzdDX1yogb5h8p+gvoyRg0G81Cx+R5iMh270/n08V5Xps
B1cnAofcA6Wpxf7xhW+sPadKHzUgxAyfbHkXC/mTKg28+kFkDWImKlmMIO2c7Foq/GHlVEzhItuz
YUncHvQNWGB9Glx1U4VjtrSuHhlGu0uMNsN9D9TmsAK2n1C2Bz7znRCxVrmQjzeB/+II6cN+UFIS
TxPhZhiDEoohhZTqW8Lt+hPq3EvlhvzUAulgQ6WnkTre8byzQ7yRrnjpzWFduxCQDl1hbhkm8YRg
hQsWoeatNf3tG58qwm9PHD1ip6G4wkInRB54tLfh++7G4SxQ+sL+n6BXdZet3hIDbEqmmr3lbytA
75nIU1DeeKr1mZpzXE2Ps3ICPDZSfZLxljmZb1TTCWHjTJc1s8UOqbkAQVK6h0fu1EEZxMggkmAN
X1KMloN3nsQsg/dZVfXIeP5z3zTJcCHA4bbABCm+ryod0WypDLbye4RR7S1sQKfQ4zmQk2vqZ9du
vqX3+N9hXF8buhEPEPFyJwYWDeE7YWnvj2LkElXdyAGfa00PC3A+7TQbOiFM5I8imVQUKmcmr1fr
bjrMsDLKd55wG82s0krC70h+aGr/8/1qNoBPmfdw7pZqVUhMMWRpYhASMp+KCAZuKAebGAHgR6GA
zGXYwexqScqC8QH50BBdFkxp3ho9LpdBLHYwdcQUXgR4+IXCA/hJrT2+T6TPzFTqUrINpqvFpp5C
EOUaIXnuOpjGTa2ljUJCEAIZ/a2YNGoP+UeK4cA1m7Jy3IoHvbjIXboZgOE7iXAqzfVNggSld/Kt
G3oTTEzSnpat0xdqYNuh3Fp8AJ18GMw9jG1v5PmzJN1J5+DbhtWTdUQmI3uRaKTSd1x+dHAIrLU2
WQwieG/nrAZe7VoJTmyeIzVwcVc5k971ZQnxZIuGx8Na0E+bSDy9ffldOZwZRNy5TNAy1lBxkNc0
cBWAH0XlV9I0XD1Pr6RiW6Go/E/YmtJ7cBx+jrYU/9dMabph+9Unjl71YOahlKTESEb/PLW2RorZ
5DSG4EPr5PHUgAXc0B/PtuPOPgbJzCo4kr1CHtJyex1xhJbayEzb+uIGAcdPDT6PV0w9EFzJ5jaA
EhjeA/S62UZJRr4d5ijoCeN0Hwv+82Le3LeQcwUweQ4vj7IkbgDvuscpOjsiX9mWrBtjlGJNvCTR
vEI7mva2/PHTWGVeGX5ds9KNRevninaxAKjHaqUGs2VuqRCUaJSmefXMiIYMeYnnKH0EhQfvLGbd
0HubvHMdGivopfHgyzN37F6EWFOJI3O00DunZ6ijc/FFaPzUKodOIkKBxdm5ZGYaEBIysZYUgHk0
88ZWTSYX7ZOcHBE1QYA35gHNV/FZScvmkSBL7OTrDhtYB9/MsKKAjXYsGJDTVdkr9n+oD3Q7pmPL
xfwxhAlvH+Ktk/PHKhD6/rWt04luhw5FB3C0ZwnVAxSM5c6gfnEAQHoXlkU943vzsEpBT8I/JDj8
E8IxU4G13WK3pf1uJZveeBQkYzRxrT30sBOMnMzRvydiU9OIqtN7G3cjQ/0TOJ6hY/vqd/NjBZ+n
IRcuPrSssp7NSUj45GTZh1KGkT4ubgl1Uf+3Juk0/xzp5YrAgbYkY0BuVwCMRaaJS/iHvE6/CiIu
mY3Tr01DXt/YUxvUhXBk2KM0Kf4qTgeoHB9PMueZSfD1dDSnj7K3WXoBDtvYZEZiwhiYE7eJHXMs
Z62KWXW0+W5A4zNw0CVdVxLwDBgQ4WufaZ37ecIxvNZh4t5FVkhm2pLvsjeL8rkAi5OURqx5pqal
Ebh2ZrYNd5FMnTsp2lwgRYHp9nDrwbjA3dF4rbXUkPHqjZpfqEjkeSRrZBGpshRVXysEx8YoytYJ
fIq2UspFgApx6HK7P7z0bUx84dPIifRtRhHykT4T1EomUfCIJPIoLGYRJIi5P7DY1DmjGdXuHHTT
N5x+uLZ+x2rB84SUam+yqZYu2lkQslVIQwo8Vs0p485gLk4xNwhmbQSJi3lEpVHdSGGjXp4r4NeE
+eoTtWcDnhoN7ZoowX0eAr8a4qhNVP06FUmbm0iMLzbVRCxiVtWiId6ghpJjDg4W7t2YMXH69cxi
5e2zCc9ZT3IeGXjl23IAjLiQhgrweNOq0QBdo5GFmf80JQij/zV/F/6c7MZR4xQAi3oUj8bPQEvv
CEBPNZ0pDW3ZhoOWwCMu1ZeCSSAxO7sc9ldd/qSHjYLAJvzaIfxyvcsk3OkLag+09b22mxp6WF5o
OSb8Lgzj9hQXP1DIk1M+Yzs4UbXw5G6yT+wllGXOqIIBFUBr1mP/P2sqpDONyklByCigkIv2e5Mh
i+OI9tOsLdM+y4TavuNw+3gOC5yPq8BzxXQ3YCnM64au9GfrB1KFDJQ14TC0AZFKd1EkuYueYACH
EhNcrnVBaixnAoi7+QKNhUdcSqjGemsKKL/d8SnSg/GKpHfBXAdRASA1adusv3vqxlaMXKytW7Bi
rFpuRbkAyx5SlkgC7flf5bIyhd9cWDeDCrp1vCi3D8aXEXsEbw7a8+fW91gTVQGT47HbZupDI1oH
ViiXQf3gcdvMyUBdhVcKDOhBzDBrSWGpqtYtyyNfimjSdfsAPGb8bwAzZliFmLqpyzRlkhgm6VyP
Byu+AIpOMGN8lKu7i+VmNy3qm59ihrHHlEMP/qzeoKD6AXoYVCZSY8/D22HSk6PN+PVEAO0BLadB
P0pkU4ct3SdwibD9o7HZX9W3Tvv7B19Dk3caOoKBo2LYRvWGfQGerxJxKhBL1/aHxjST2eGecHSY
tAliGVdNg2hUm2NoidR+xdJd2zn2iD3prQDIJ/0HZE5LoVswsgcVEMqfrij820+aGjNWIw6bV4aI
MfRgMevbu6LGpNBNkIBJS6TI4VYxh16UMK2s7MWe4TALtTtRO02J7FvuqVncf8zbLUt97X/dyAn7
XxUQWFMahZj5Cukw0rzDtvUPtqNCpMYc4aJyaaV0GHsDdzCMx+2rv5AfOGs54k1+B9UnwATON70F
koNPtcvgwmxVPOTRBzBAs0MsMOCfnK5mlGRgJLW3KTYA3diNO7sGhHcTQGSslfPbDNViHxfsKEm1
zJFho8XGRZ8m93Vxvjdg118bJP2QJlF2FL6KyPPIEoN9i/Cli9KR4I4ui8WtcO3Vr22DHt0XM1uQ
AtoEi3SpkQ9yp9FpruuG1us6DBDbcTd3EYxTfsbJt0726ZidaFuHr4Qjm28V8vZ+VglwwDtPQuZc
gxoUuuaQndkSOfasJE/YRoCjJLxi5N3bWC9W6jp6uPKtpFtMdeDClBgmTpiiuGHdudLeBBTKpGDz
09qehCYxg3Dgq9yyFeuIiyswcZbaY+41Kxph5tfimnzp6cLSEvG4FpdIeVbZp2fEfBLkUB77kZWx
fj/jBjEF7hSWDMzLWEMR6VtyAKaETXkz1CiOhSWvvvkJDJcTRgKgFuFIUgK2wsoEifdSi2JkLUv2
igdt4HBzYOgcjFL9w1ZsEJqAmJhWFvTf6ogISyOv8wnoZlNx83E8uWMW2O4mNuMqFY2n0gieXVup
m3qmC7IRQVv/y9N0tJmkRyAqABFQTkInbZ4kSBbyYNhneCK7OEZY2q5gY2TjsUy0W+SxWFMJZG7Z
tvIQywgoVMXRZMLOZ7sRQqRjjfFn8UktpPzgfLB8QoiCj6x1VfrvtKzhnMLsIjfbpvnIS6R+WIST
A5kYtotC3ReNSdp/C7CEJQ6S0FHdlbd4Rz26dOHISSmFwhFg+53eu8Z6jV2QL1zNraQw2OC2vBsa
quVdOL1fR9bDKabf9uI5Le2XCWNaD9slTUl4QUnRrkgKpJqisdvBVTd3dCQz3dYpeFpD6d4DS8z2
WbvoXoVGEO1PQN3xaw3boAkoMb0Uasu7vLQZHHUgmwmSlWIW61F2BbMWJBp/STPZnOqDgemVPV0C
3g7LbFUfZOSbB71ri6/31nk7D/YxVp1iX9Fv81BIWovmejvplEepCs8ycPMqM3VqPtWu9Hl8ZfVE
eSwB17fb04NdUojG3EwKERKXETppikyonSwqV3sxPfLKL5gCS1gjsMZW76h8kpCH4vF0ydWmqF/H
yZuMMLqLmPWW/3/Uxxa9S4QnZXvkPMcIdHS652bjUM/Awdpt8aC6XgXYk+sYKckWoWPHyqZrfKbU
++nET57u5LZG1LUCI6AUsftd0dKkyYbpQqJ8SHw18aokDoOnNhehVrEJp6qyfZP8ELZLtbcU3W+Z
KUQUrLzbGFPaoy6gXo9ZRPB4yHX5py/ywOhW3c+I3+u1RwN+HoVKte0aNQT0ZAlS08xiH0c1hOCG
ZsaId6ub+HKpOr6oxP5brm8PLFEZntYbfQWrtRf4fkxXiQThKcbrc7biPnKNZqaYylCQMMsy66fN
pkpIL9lS+Etl2Ty5b3mmMcX/L9RaU5osDaHgKMOFm9cVTmv6/ehSGr3TBcSCFDyGxFDGRTtwDp+n
iUeL8mh3c0pAP/pwma/GDj7wR6ZM2xCHlaFxo39awsS7UnA0rX+syCStUNadnCzF/8QUoW+BOx3x
1dI6IG1BMegxNpN0b0sdWF19Bb1C8ExnBhPWyvpWohbLRq7nYaTgTHhZExklofZMWRy6olBjaQK3
ga9oJbzJjaL2uahmjtqxq6bSTfYthZH6px0ZwophJpo9XhSpocnlou+U8cRZdILxYHiEr1AxfUBL
q/LJBZ94Dyh4HB99i7nEq5kX55QuocelJUdhJUYIBgssYUSp4kH/rCU7+lNkR83V0S9zH6cMPuNu
WegHCKF9srSn2X1elZlrK5uBLvZJx/jLS8Ac7wDoF6DVepCpbrcnVq8T5F2u+Q1r9K5CNkYZpNUL
LLTFwJd9OHqftzh6aWeiIYTH4pD/D5DbI5JMwNgsfZQrgsx68WMVPL2LI7HMOtvRzLO9rs7WFgaT
onksI/qmoow8sqShrhg+dFciQpp8sS/f1rLiwm30mfbUd04Sg8besGHglehwf/SlrivPn9Lydvio
isN9mV4t1tanElSBAHI+RKzFKnwsmMVD+vLoi2AbR9qwM9HK9ViutxpN4DoXTA/8FucaiJhQRfjT
pwOWTEGRp8UQN0Gad0yd2sGAUh06f4etWnM+VKFEQPCgfiN2m59NPPtryjkZ0lvk2XJm6hcoChE9
bmkqEiK5neXZkOVpb1FzZRjcinAswxPnBoPEOVKQ9ILhi7t0ulNTwFleG/CzL//VhVTflSZEvvMm
wx0/kkG/L24bqt2CwVQY3EWU3CZL6lFa8pSClzV3CMrroxQg4TkcvcpmZwLLx3tegpnCSP5yTyjc
EOEAsJ85V0HNXNqoYuu2qPBqOXGE70EJ6Qf5KaIdX46UfZmheMVYZP6FF3QMsImF9QI+hmArEQAg
Zj8cTPfzuRsi1hvZCb3j7f8Vr1tBRbjmlAmPDV+bwNWDNv47k00y7ILeAHx3H+yZM9d/oQ0ASNgR
osjM2NouckQ2xNryo8TFOrVz32BMIDEDkKog6Ehv7bCHb/+07DpvRhDZrPvjC96LR2ywlRK3wfrq
TcP59J4PzKiJaq24j21R8JfXWQZHzuVbldlLySKggZCFA8N1eI0M3YN3kzGzrteiZntkdFUDHhbA
x3kif4oVgwFD9Gz7EbhM0R0o9PaveP7Z6T0zXwi+AX+/yteY6hovkh3hatY+0YlV0fU7+Fexp1ew
D65dVBsWystoshySjs/MIkow03MIvPFNRSFV9tjcgsHhJit/v35fCGd4J5pH5c51UdQl0W50XFfl
3QNUFh3ILiVPv89wf8s1HMfPXVXFZ9LONiNJg5/fxag2kVoD2R4Bxtn1urYlwLo1V98rUuAsI346
00IX3atJHoIV2oo37AGa4h3SMvGNou/lm/5mP8B/NEM9rhTxyIcn0JqbUcLk+SRUwnmiaV8VMze7
c9f8xTVodKiwcRBSzECndhq3A34zxPQzLDIreaT0NIWtfpf/ykBFKxqN4Co9Bqx85WDarJ3l6epZ
/hxvpg7TfC39Lny22KoHr5c/sqmuAoloCpnthTxPAiGoFqReZQFm68SxO0GJRPx1/DGHDDcPASbg
rkm8k2frVAo16vEOlAUpwbdm+S0j0+P47qK4xtQOdEo6DC4ZgpeCam2rMKvVzGBwQWmt3+f8PRZN
CtGMnf6khCy7HeqXUmWPHSJmS028StIlyF5gjzxj/e8SPaa+hQbh5TiMriSH1FWf1NYttdEgX7WK
xLCb5BCNCE2jlptZe39n96Iux8CAJjuQleNIpyTKU8h8Qyubo43bJTiwH9bWMPUWLmoG5pCoU6NX
hAV3vj+zD+4TF7kSG24GqY4s4Gp8GuvqY14T4Zd+sU88MI3Ff1t9mN5Oz9RL4O7oh7qDcSLGCHpQ
6VgMUfuHWPinXwC3RjvMPxAMi7oFNx5KuKGtD2mIHNvnZ63ZpIlLNJ2zSTtVJUv5oWqNhL8HCdzA
JVC61rL6ln0rjRnPPsZzdm4SVXObzN0Ym1nx9FQ+wnWZ50qfnJAOpdJ/3myEMgtXtNpf9vzd6NZE
IJg6TNZbAt44scHvaNKX2PowJhcJVAdTjg8nVNafZTluXPOaDeyl6hITZwO1KXoMaQTFp7plLzSq
NDaB7XXys/Qss/1GkIW8uKJ//6NOgebqFvI/dtcpP1CJ8ow7fVcyoRUXwB62i5+bEnuUjuuz0Asc
cmecTTtECp+LNpchqn8fa6inCQvz4alNg1fJU3HcFTM0XiWsS1xT77AL6SIVXFsMlCGco1iZ+zLl
mBSwhXTIB0TegEoHJJg9DH+brQdnFRRu30dvRtUqnuJDhsrpS2XKkjTU/oer5QvYr3UWh/BYHFVG
SrIGp4LhKR6ffbpqIPxTsMpiJJgSGHtWrxUyaeXT1sbl6lqFtL9zBQasyagCk8lu1dMyXXB13duh
aD8EaguGmQ5YpVb6RKVcR0z2e7I7fwLmGwFlywZQvZIXGwJlTy1QmXhQqQbgyUH5jta0TWGsu+EM
AdxBjz66J1xvyaqZLLjNukkIiSnw/NRsFCveJf38qQiUHOWJ1AjK4q1FxguYuy/U+erZZozXjAJT
71ce9ZLtU4xLo5p6U9ySBsGFjecPcM03qEP0Gkh3K0tINsu6ar7U1m64rOZphajYSUbenKAYiXFB
i+Jvcxq2J53O0pZOAJDYFipRqGBiKHmhJF+sJyMi5zDcBYW9iMxWZ7CGhgoANEaxXR0cc+PWL4pT
hXUyAAEnuPFmML20cvradDj8B6ouIoahiJ433vqP1mt9hG3TeyAgwToYT4arAlNXL7lx19COi/AI
gXhOFEZ54Adw9GjhqUDcfXuO66paSN6w+4TIS0qCrlMaPJKkTqRxHMgdkzKS1M+d/Hm2biwfpSgh
Usf2gcml42Ml84xV37oTRN29/u0bhCsCHsRotJcX/XBSoWS1GEIDhttYktDSXTui0Som1muoIgAO
LZYMmSIrDhQZYCLIuIYtZarrebC6d/4Be60uMkuM9C08PQoN1JdgEAzakRmjlntNXV8yDiloKCBf
xkLUY1R9LL30O7OH/VHxvB+ZSmW426WyOlDnfwV8BJfGMMSAl9RO/dzXhKEQ1qFGMp/Gs0awCMON
uyV0PG147pxTBpCikvFARJTVVGAxugd+EaUG8F4av3ekk74p4NoR5ENOH7nicfgGivr8qt6l6bxE
cwggOVv5n5FaBR8pyv0qhx5W8hP1VavTXOEnHCPJjAge0HzYLwv3ha8JH30FwtM1UZXrB5rJfaGb
pFlIlH0xVxci2V3TtwIzyWWfXyv8hMwevO0DF/Z/sgsn72/jMnx93e86QvY+fWlBsk0LxbonBuLX
ah6EoEKx0XGk3T0xzpy57zBST80bnI2K9+Y/48+dtv2WAQmBX/RqfwVGOltMQpDO16+y2xiykAMd
NHizRwDa/VDIn71QxBreW2itKGdpQyQ+YCXgMGZasK9pajC+gtNTiSqCEBx4Sd2BJ1r8wn/ArsPF
Y/iVlrdPqCI5Z9UXkVGoeznBfvurHDcTzuriKmDVb5TJtkS6gws+RloPpaT5zQGpzzQfIzMK+Ubf
vwcWz85pVTPOP9tCbJZ/3cwzapbUfX4FfWLZh2EAYVCquyogXYC2mg2S2tt4QhkSjk0IYhaePhTb
j6U5xJLFRWV88DzeGgvz1WRhDiyVNz8Mq3BTAubDBRq4sa2sRq7UAvV8VZI2Rjeg8ARljkzKdqWU
wv4NXDMr5dApu8VY86BBQ/ukU48Mt1wFNfflH/ldHWiU0vipBRJ8xz+dvyiSMS3tRyzCsCdSeli1
wByObMSX46AaFl9vK/g+b8+FJQQMPk0UmreYhSaEvDOBIbrbKX7L/SGDLmkgpehNtDSrEsw3myFD
XMYJ+Xt1aTeJ/XFuhMwd4FpYcOmp5Y6AaNGvht3ZFYD/RirlGr1zPqoWmjtIp+V1oASga9ziG47F
NT96o5NFY2z64JQb+V7w0nYAq226PIDneHUvhQPbyUOSSAS+8z4b+Xpf54UWBAZEBWI/ArJWhSdn
efgGMAYF+YWeaD5i09tWHA327ikg9KOAz/MxWAmpXz5Sgf8ckUz15EEcr+HSjlWCSmNAag+VIVNQ
KaR54a+sv9pHDK54g8haFlN8PJSVrh0pcJOE7UPGZZM7OkpJylSWkIUVz9gcn2CthWzBLT2BCwba
RI18Gzg1ZZWS2jfU9F2qp2l8rfFv5bLTncBSgIROf7JaASFsI8olCxujG7L5xSJLhtWgSXb8XOjd
3BD0IfGhcz0OQ+udyMTd26YXKjtrhmyHRX+9DjgqSiT1cuq9+eBuON8kFiDc3Uv95sghcQsHyBwd
MINam3YMvfVBiciDzOKEIIx0q63rXoCw2SD69D+B3BwxNnNPDE6EHaHHO5C90svadVA6eRcfSQL+
j/u4OTHJ45ZWAjSUGwDakKtUJF1dCje2eT4M+raRBOzYRgdrL18h1vMjGreF3vEkm3g6P3RF2WTG
k6tpv9f+7G5PKxPV/N7RKjAuiwk+L4sz7eN4RsE6xDFuoxANsjRIMDBYb/zMMoQgkWUbCiwfQnxB
U453HUjIopF/etm5cibI6p1ZfZ+C1ZXWqg6Eui1Ttl5QZASKwYRqME1Jq9FIq4CTKSG8yaXoZjfw
/2OOVYzcTSldzhkGcdxQ8ffb7OLnTyn6AWYLmiFtcJSp7zviJTV1JfWEDV984R1Azd3U+Z1+o/Yl
E07bNAZpb1FZ5n2Sbio+9AiC/yMphg9E4MozMEkz15LAEO4xMKC/IEv/Xz17J1GZ0JTO6kGxxR3Y
MfA5+EIejBfxJ7P94clMy+nyjiKtTsRfN3HkYOHjPI0WgIjwiMae6Gitfw5ElIPnKQRmI2+NXwSp
iuRWSDZdxRTdX2tFgeFoczfgXnZTNqDqEFc5E4+j8+96XGNiV5lUuP4JiqfGE4l2Y4PJpy3KgbaH
SWp8Nsf4dpX8E8GLU9rQxCwEvsNF9jsTjxJcr9pzmSbsoSwKI5Nw6YxiPYRh8cP2SNrkN+02DxDT
vKS+3HQUEudktH+jgO3qiXw5+KpsHP57YskSiPrUNclJ1cDkfg07wRL2bAKqSkx8nrGF67CQsbn8
90hQXyu33rsqDd/vCuruRhLT+uo2OfSq+LlQw/6cdG+MAfLS+km0EpkfcsegzNM6VvxSnV9yHbhl
H/5o77LgQkPjYNrek6yQa+q+FSMzTQXBETAYNe6tYXe9i1JBuRqtB+n2lN0yGWnhVHBDsCvyOUqT
k7lTK1QnGBlnL2myEvczvTsdLIFkyLEh1FeN2XxRQceVuykZ4j3v5nqINqd1lMmljlUYYTewEr2o
e4Jvy0yizTG+WtXl+PRUF44rj8iUqoe0Z+fA1F/Y9yAkzsngOLqYzwD3aS8cf4QTC1wgAhz60LxR
JFG+1eI15Yy2HmGIpB6lR8JEQcrfijBy+hH5QnQ/iW4ODJxNk1OKhXpoJZGfopTkA95jt+fTdaCG
AsdeI3dJlAX4w9Ew66T/xS84Aj5/Ctu3VsOjiHUCZbNnyVgkaUmt7GndNinmj5FAF5fFbW5d8zoK
DyLoz0lHLTVeH94B6B63aeyxdGOUEjk9yrQa7kwI90RuQPeUFlJ1Ma8eN5Y8ncYGXi9uMHtjefxC
YmlRrqCF2D35ctpHLQg8VYxA2mfXJw81o/40DZhnCrXg+n+Rw1EZgcJL8+cWGSA6n2LmUMDo7MbD
pj62TuFUIqIKyrz77w5vZzD69opmb8Ek2uTwdfVrN+Z9MFi7+r17PQyP+7XPBuIbtt0ZLiQEM7Ua
Xl99HCNN8HQnkLS0xL3xBdG7d3nzWtMWG8OC5lCe234QsvS8ceqCpeWzcW4nI0G1WUkpNZhwQBs2
LgwoOri/76saoRm30VUe9Wd2OlM/NhUKbLnjzARJmb0mMLTubWQGw0w1+ehocgMRUJH/jeuWcNq2
SGE02hQZDDalXgar6FVrINrWCnDZjvYGRbaAHPdHS9tAAg9wU0gxLjblZJ5MCGeDJljOYjl2pJ4U
dLHqnfqmgaxAw+6bbTrKAqvxDW5RaXt44ITyDt9YkoRS8QdVnY7xk9wBwy1DnkO/cjg3pJjSmPvH
tuV/Dt5BpDIiZLKT1gW4y3g7fTM3YnPG1bNaSPOUWHdrAOgJpqBkIa91XLsJG7Sf/fiR4Kv9CsHo
YUdUj1vTK4aUQycZQK1/1sIpmqa6eX5v7xIwqSs1C+LH9c4dQjrazvytz3d0/bKlPmULLsO+0beq
JcfZ52ojGaVGhkmd8qmsGHx5f0mVyTWDkzZt9jDeNXro1hqym3Vbur3vp6peHy6hBT3SML1Xahw1
z+3AGEv3jF6lV2rq+KqXO8vHG6Fnkqk2nfluUeUEOls5gA11hq5SsvFrAruvkMo9DrU8PqshffKZ
Oi5OSjPed41MZIJN8d/WM7BUyssYR625XvOVqN3OsMYgdz93lPuEzqvwmA9Ex2ydFQFksHNgJFA1
0frFXs6ig6Mq2pr0ulk6lF69+J9zzPH9IQAxL/V8wl17rRYMCUN9BvvnmHQEL9pmQrTt4+w1GyuM
OeIXFXQehPgee5dZluzGGHjtnv9+3iEWWhr3POKZhaaTTEN8q3AG/yJwNQeIs7d12JXbTznVJrn4
grjcFFXBkNK12SAy7EoIJ9LXl+31NfuaSNHc0C77ypOM2UPuN76ySzoUGky0rp/X3RLGVIFrihgF
sy26VGFdIqv2QYlpkCfl/FuzPKQWOAvqU10hI6Os6/dmzVaFHoTmGYH2hhqNAR4ljuvS9j6/EOzX
ognVrk2NVqS7rS7KsmLh8UX5THYK3tVxi0OmbC3ixpJwwYu35cv5J+3zySPV3KupCdT856levcge
dXf64CVoWaKasZ/rSp6n3++gu/WtbTe0Jrd7jsF12rotTQPqaEEDmrie2XsEkNVu9ThO7LkwemuB
NzywX25qpkE0m0HdXZcc8EixUXRBg8Rtf6Fo7y16PBxcci1HJkZzO8TGXKKOp2ec+XMk3+aNBXKQ
hzMwyOXsfRdHcu0OpXZaWO+PobXLvoeDjtiwGigX4BKZAsmJvncVkAFIKIHo1wTRKTz73v7yTkMx
wn/VfmEfiFQbBx+ZeUHT7n2c1v/Zf6CyUuxXt1UkgdaARmk0QkljEU1U/8xSsk+FUwsj2c28f6DH
G8Rkayz36EXR/AKcbeYKCg5slc34Lr8VJpPLeNx2jUTLEXjMqV8Za2OfWRc+E7CBKE1Ay6IRg/td
QcL9VwIy3z1I7v/mlX+Gq3nik6MWno1oQveyWY2EUy/0C2pzZW2Hpry7lGV23fIKEFrogy5N9GxR
Jy/fA7HMXZ+sDSBljoRplBIUG4DcJAPxjuVhat74j/Z9G37B/gvDSJCSWFl/FP90Le+9BkZqlj9S
OC70Lv/EK7P5KTfFxSfRp/4RkVth5x882jKq5Yl/Krzasss3pNNuxYcBo1f0HcWVbFnJHz948195
4g/iqWFtvbeVP38RwN68YkYCG3zuNnMljN7+MTIZl6rHVzwFf5mMP1r0odx7jSiECykVXatMA/4v
pb1LWZlrLwKdgUIsVvS7iW/SAdMCMVCzNcW/IUFJCCwOcYoX1xFi1gRmV4xxiuvFzTHcRk+LXSdl
ewJJf1li5svKsnPBDjvO+VrbhrcAWiNDV7xtDS0dmakpXfaeIS3nTeYupe7Cmzd9t0XuyuL89SVV
gJx5CydG6igQlZBeTsNuXOwDzXRASwmh3H+ysv0LYUiK392+e9nR1ttbZi9MJJB55xGWWiBybQC2
IyoHu7wFCSGALq7W1o33sxJpsR2tMSMyf9p9FNezL9dNFSRmVhKJXKNiQlBejyCgvvch/PiejPiL
mmFRQ7v0hgHDoUybM2S0jIGUOXKMEEqVrk8fBTvtwGBK2EjtViNU27P0tVk1euE4ImPJ/zWaTzO1
6CQN6WmMnVK0SfoknlcitXlF76pPzAim+3alqMS4V/zvgs/ez4odluekfPhiQQnpi0etEAuo6+GO
e5Cv4UF27cfiTPxFb/zVTWqJpczPnxhsthb8xaEUCZSyLJVUSb8awewm/DXUSWEaPvuQDAJVG2Cc
ySuy6Rn1k3V6ryWM6sCYBy4IdeIFGJ82V4xPOS6AeU9QOoh+gch+XqnezV2mrfLcUFeb1MSAKv4o
PKSYCPrtaDguntrcM2cevdTqB0ftYEz24IfYwn1qvArSdu1UeGAhCrnck27yiEQ30p5fwDIvRf67
4CEdJHPOfs7dLptvQ60R7KSkOenYC7CsMWdQu4btwR22Yd8ccdcWGe+mZRkA5OtOe7VuAtqqPgCe
p5zAIHxPoG9+IZ0DdcWWj2NTb3CEgm5ufRJsHTk4v648ob2C7/mxRf3vbBlIB1VM6d6OVFoXCsX8
SRf133lIvwvijyb+reegexudLgssFfD8tGRYDeOPDzBMMv2x+34nT8ORmxjaeB4UZP4RzRFVCpCA
9y8wEu/iG5gz9/k6kZc2iA/70prUPdr1Czmh650eJeTQ2esMBnNSi6B9c67Zqj7ef55pHl7XJ1Yu
HoUEC5/d0ejrl7GKPc8PY6TfdYIiu14f4D1j04aFmGLXzSR04nY3HftLV7tqrUIDiZ2WND9zYkuv
7XrHXhsdCGtv3/sK5Ep4ej1E0BPQW6V76uv+WqxfkaSR6XcETeTknLRU6Deq79dyuG8VSxgOq5qg
XY3oa5KaOARD2NgdclXp9BBI7mcaimDtNntp4N+fLpqOAqzNY0ehgdsm0H7C5C0mnqN3YVQJl92c
PZD79TbwG9In1COf/JWX4tZA59jrFteTlHGR3F9YH9Ni161zfLpfBviuHHUau7TGvOunQwgrf9j1
CtY4ZJNAdv+Wqt2X60E2bWiT9wDgFQ8Odw2sScMoVSyck7syYlbdNTqOx3eDkLhIUmw+zD8ZA2Z0
DHz72UKK+plw2SDOFEls5qcWt6Sw1ROVqYgoxnTxqIOT/6cFRJQgxbWHv6Mi1ojQufy13qestXoa
mcq0vX8mWTMmt6ujO0CX2nk9Ep51Cj4J0XQUArZkkvLYukLwddghrxHUKhOYgWIftztaophBSnyY
XEjTK6oaElnwLDPV6ofy77kvXfCkAYpdpDD+wjcVdO9j8zoXfAHek2ugNCKvHmlFAMpCOvSqTTWy
/cll/iyKKuSXyLa8oXUAjXGWrP+c+lrT7AX+iuu8AAOBJNaF9dGiXF56wk3UjMAX5DPV7mlefKRt
TFYuC/lxgl8/UUIyOdLHvYAp0jVERfw3caCm6AieD6hMaH7LAl2n0qeL6OwtZox2iSwG6lZD6kZj
apklcLyjcE7Z/oW5k3MLmR8TdlBtouOTEokeSxGITAhY2UzFp2jeiQQu8fZ+Lz2rnaL6KZWie7KH
oA5JfyRaqsLHcVfA25O+/zBVHOIZs1BMCQ/Zg8b4APllv+9LtwVqlEOQD2fKuQG1E4MkUq/cSz4K
zPmuQwqgHzfFnP2nBuLpnz3m++lvwk759kVBEKx9AbyuAdjls13h8jxU3gjjKKHJU93+KbvW5DQN
MAWtfVJNmtSQjW7umq6as2ylcOWW+kNstQitT2xbOZ2OLreNCgCyjIPHyX+ds1qviYVUQOZXutqM
0T6oL06hJOZ2kndlMYG0mhh09VfA/Ok4OKyap8AAe1yXXMuh07X3bPdCUgUYHqpO6MxDK5q78p1L
7E622ifXy7LQg3px1fRu0ioz3GFDpYPkLxk1pMDXiR0o6nh9g8kTwMccXuR9bKMdvfJj1+TkbrTy
JfuhilNo6zyBdWjdWBYb0tzKavTYhB5POj4uKNAVrXKSpTQa87C9DP6LfGw9nteb8QASPVcj6f52
9fTguoWfvVbGnJBTqpYFoL0ZMNVszaUANH6nVXvkrv16qL0FTCcPHMVonge7hqRaPmq1jSpemsxq
FjuHbTSdH3M5OpaBvoL9xey3oE2C1fhPGlxoMLO0KFTbiDfMNXblTF1I1t8iQfQVIlycYPDlWw0s
cwGzazFm9BxR4otkirwWmMlC6yj7UrrxVLS0j1jx9nM1RFGW/QFnN5rPfhaM1aKgzKoBvNPSLCsA
1FQdcoXfxXx6gguTuqB1iJ+XeReLx+W05vq8h4ghaARBKV3JsS37SVRcxn7nSR4E0KhnWZXxUv8K
992oeHjJN5sgLB43PR5Dvvi8lQHSrHwqUgpGsQtBhXrtlIaf3XwG6QVJ1oxbJ0EE2TU0e1Toisdq
hlgUSx89rrZP4DVX22WkzWrkQDQY/g/hDBosOHFkPPW/5ECzmXCt8FYA0ngfrek8TcJEaApIXZVe
YE8rlRrnlHHTnmHbOFpNkzCcd9NdwTqmCdVPcF+sIPC7BCGyCNcxIh32YDOAiEtCQrIG8P1ORJrh
p8T0WQTM69qvwlYIvUSAgHKTFshdgjE+UUi+1TOEFhJAEJCjq4q4Y8+rO7tBzQ0I4oD46Q9o51nV
xVt2OHzBQ/6YHdT4KBobfzK+IP7PRmH/Mnj8vlFF5lCRsGUVO7GyYjaCS+i/yYRGhPO7NVIeEM0p
bTa3LYtEJcQGkcpWzoq5dhxlhIJEvrmOBPpxvrCtr9RuNP//ew74tl9rdbsFjc4VYVEZMj14vY0N
zljCjjDhA6jDWWk9CRDXO5PQ4SgoQmXI0IJdgiIwO6QcLkxLY6CYdZJEKiP55exGXkrrdRXo25YH
/gJhb0L38NkCssFkndqEkw2Jwi33Y141lTMK49553KEXvnD637BoJRH+GXF2tDT2abtYnDGVjDvF
1TWEN6HupevshpCTcrH+4N+OUalCJ08kF/sPEGNkQnpsf6o41UM7ok7Pg6ndQ/FwtP1dLw1VDcQR
hLXmQtbxol3vtAXLOgg7BNIUMAb0Ya4nwEUP9n/GlGrG/5MSLTrK4HJHs+reVHE2EQ3GREqsTsBk
YjBdAfMQM7S2M6c9oGxazVpF55K4ILCErHIZzVJoSkLiyDi3Y+hNNPTwCrN5JusIBUOmN1QQxnIU
TdHS1cgxb6DhPNpSWPeAGKgYe/JTmUCsvqh4y1B5XnrBnSZ0JAnfm+aI/mtkgH0AMg1xPW9H9aLQ
adgCBUOMrcLY1nfQrXwGkLMs14vlaCc68/+408WKfNtV3b2/0Z7MYqIhM5WqsjIarbWBGDYafVUq
eCTjMgN9e7RV7+Fwwp3O3cRkixCc93kYvt9rbk0JExnaFQWrcwhzEF+zn8+hGgg/U2brJWMPNYuj
EosA9dnsiW6yE3tRtj6MPbzzS67etDsIEwEX2jdyyRvzPXaEhBO6yUiAY8tE5BpjVm14D2sID3Nd
GaGJ9stN75o4HsW9ePOFTQBf/p1qtbKOeSYTj8IkPP6I9wt+gTyb+gwlf2Me+1wbAgAeJsFsgnJb
k4AQPDs3yZiKuIT32W4ynrqlkg7c+83VssHJCm8zxSUwwoWDv6A8StlT98HJw6syN/q3w6m4uYBB
VurCppS/ZvRRXmip76qlYGcLt2QsBK6fh3m7e6eLNMc4T42luhJu2oy8i7CD1jYfGyRtcySG/b56
LE2wWk7Jt8UGnZI0Srq0xR7DEWA16qumLJfB04OuqSnfPUxZgd/ki2ARoYZLYQm/VlcAy5sjqLm7
ivjEC06mD2xXklbTfteU2YQyHm4NRl0ebe0yG4OxSPdRhUvcnzR1xI12Ulx9q8oLcPBkeQLroBis
4BmRssAsD87UyWlomjAr9u8HkKeS2tRdqm0KyQ0SfstLFjquy8QGZht4DPZr1pQUJ9qCeHwSkuSC
ayXp3Bnorm46OOHJK4KPPPGtHY29H3hp57bb/TqRywB9YPV8h2HGMOZRCsYvbxg32RrKFTJx0MdY
tjXYg/fmaQO5lEvZ8Z9GKwB9bYPNQzlm2ujUGoIVqgyrGf0j00U01jKeD3wEsOnCUPZHMg3A/6om
VYPJXk17f07myRSbNCanJy3ExMADp1/I+5NPCF8HX8Tl/vDmd+W4RXZWBsq5o8re1Dq8P9/gNZ7A
pmeGH4ZvC6w05/FfVGdNp0RmKrmXRmSy4UP5b0xdeDorIB9ytHRiy/U7I5VHVVSUImvjmsNGVYKA
zH2wq9Pk5hWMT4i0zo/ks6JNVObg6M/8GigTYfgZ+eEhapb0E6L2YmXURhFpCBZzrhfzkTcUe3HU
Bag+VeD7t5MM0iZ/6lSaPEmaXB9XW4qnHY7TfW76dVDVbVlZye6w3Ojo53yJlPL0d1XCNoVrgabj
n+SevRg5yNmyW8ohxtoL5sv9ofoqQezbHwhz6ywHxU78vqac9sG381p2Ab3BBkb6WMMxLbVjuYsX
dwUaPTTaUdo30iUVSTk1stMjcEu3gDFlRr7qVdAjzJtihMFz1oxqYodfp9hP7x1b7MTgCQ/HX9V9
Z3PXU03M4/41TIlqMzWqDL7MwyoKGtiwCpnNB5K0zmV+NoJhH1zE2hnmA7zSlw/RhS2h069N0pRn
PsYK8lrRAsLHVo8FuAR72/OlWBewALkR8dIbNvOzEwaJdTy/D6evRASOa+ebjopGxVT53cd+Gq+6
SyYTq0kAcptbuKopIRMYLLJ5aikUgsxPvVTTZgEv60DLjvmnoFwb0r5tYg4mhUoBiHzFeTkzbaXE
epSdcDOHnn2sgW1zLhO/kM1K5ArSH5psyndLjw+XDJPwDbOtHQvnqBKCCfU+zdtHglvErjmF5Mao
Ag7JzriLA1vZuKHtfTuMAOeUZ3Pus2M3Yl7+lng9ccM8A2IorkCk6fG6gB01E8cECUkaOnRVZ7+d
olufLq+LCDT6bSwNffKHyNwqHHeKGwu9LHhTVISDOxTzabhXtNGlMNHZ0MneCkPOI7WQzp4eI3Y+
F6EZeH2JoTwsvHbzAC1AhAJVoZT0GkZJKCruncPZ4mK4Cm20PFOElfP0V5HZvoDg+lFrZ+CY19Ul
7nYQKoTLZOz/dJZtPh6mI0/G2d8gABxqBqQvgwDkRZJdcqFOMQb2kc0FyQ+Xef+pWbvfM07tQAx3
3fBe8nlw3GfrasFazbALz0FJFripj3aHE2kBhNuT1xE/InyWcuc40epHR7b/AMyw3xzbnoksksLi
sAeiwfFaGUk17IpWmRkq9uOKGG8LUr7xtDR9VAgiMoRO7XNYEdhX8QxzN/obJMTkgvN/9mKr6IOY
avZBkEOfYPmCoFW3h0tUScRTx1sBUNcLHOezt6vhR1/QtJTSd65MHfoh7NrWFfaWKGjy+92MIBtF
921MF0MUWswgV+lAsQSkur0kwVTaCafYOXYXkn5RiKpd7L3/okyoU1CJNoa4JT1RPdPPgLZYiFId
iCO8mqvNSi1ZFt6Eu7zRXYU8YiOnjS/VCFzdN6gfKJT6HvkwmE3xFaZLiVi4Zam82Gf7iEDtUaKL
taFV/lDe+vU34aeuIgrtm0B3qFnlLq53eKzrfQivU846n5e7TjgFl9iYec26tqD+Z3j5Pvk7uwnN
+4RMIZf75J+obTv2O4/z63bdzWcpY6ue65y5Ja7LlH0pBQAogRRoKuz5QS7VI+oAwAPWbBBMaeYm
j8HgP7L1tUXOaklv5ew+D/BjZOPLWpZy7c6Ag2IVLIW7FSYgdXE8kW1xCqYadFO6Ek5p5FU0ZaO3
Iqls14IUnMSZ49VOvmhJ5UaffY//Ue9YvjnBfktn/k7RQi/pFc7IgSnucqc341FdnTDFzWgZMjMr
K8oB23vrhAn4XNnz51HO03MTpjmL+U34ngoUIh+REnem7kXE5GLnRItXHnzxVLJtW7yFZutgsemG
Bc8aXq+qUsbcJDQ3+GacSPhnpREWrqCy8kxQTjkXPL+70dKyF+EDVAN2/BkME3PkVGfZcsJdzpSM
RIFnuCikRIds5NkkgazanWZJChFDkzJPwdb+i5JPY/m8VnZ6tFb8S96mgf9pe5sODFM7ybrwgONW
A0/h8PZULW8cbWIcrF8akHiHsXiCMPKEIzBQ1JCeAMRBWASH/LKyNoHjtGBK3UTEwd1Xituey1pf
ToJDV4D6bYqLuESSPXiTVYmzMewKIKHbxwLN7prAytjoE5+PNAkCBRZsyUivnROERcH9i5giBszk
zvoV9ob9F27ez77dreqh3kgwUZ3mjOdZqTvLMwxSd1/E6pICMZJjUZtha6MV9aqe5BL/Dpn1DHkN
5Y6fnss4VkvrhCfRL+SEmggxen0ZBdDC1y0b5ojT0AB7XJVMDIBpGeSVzT3A9I6YXNteMlxywHd/
gE8ij+MV2PNZuK4i54otz/wTdXhR/8Mppq95siojivZYe6VQ7KlPnCXxtP7+oCEDqd5JgvLIKQqh
oLGLfrOwPh+DDDkEcJhj1qkLoU787R/B2W20VKaSl3cszL9IVKDX893YsXQr+XwgME1Y1GerkaQh
Kdh5fVA+YUwhOi1/7nEbaGui9LPLP/KrSA1PL55tOrHnI32Q9txGn5xtO63fIsgrzhK4EG7/3Wo6
9A3mIQu/5QFjAFyMwVT1VE08BewaVUo8FFjIE+Mkjk1yybYoO1EBE6Y84b5JcFDgMSHqoBGsv2ZL
Z/tt+ceJ8Oe0UXza41XGQiFcOXWtR3dMgZcCjjQFW5Fr6g35/3djLbod65jIsmw+yYfDnQuddFyv
6JZXxvA8z7WZ4dz5NciTwUbqXPWyaN1ka2mueTCmO4fcm0YlCTbtQxC3b2OHtUnmWPKzdw7d8bBI
POO5eUKF64cpvanWssD1l8JSjRHoP+RYojjrxg9v1i85kRfm9lPZdXOwYaxcV9G37r4pTLlzNXw1
Ue/cEq4gWWAp8FeOKi8d9SYh6sD+hvDZ0MfAp+8gUpzjqHIxG3+GV2rVJrgAys5A77l3Q135rodc
pL7muFLeJsWf+bj+YD6dlSgcBLjtGWeqcwc1F7Gw1jv7tNAWB1/StSMnAGHzWwnnTQt0tppaJI/c
4qkGL2G6v9woTzjWI7daNDou9veBjZrqf0bn4bJz06Gf5sBtgMaKNNcBtbdpcRfxsyWZ5uBvSlHs
9ELZBTa4JpeQgK9k20bTzg1xg1ZqomYhLy3bFwa38ZxQ3tjwYQeTAFew5QHpf4g3kcbQtYcqTufp
3oJscbJFwalDOMR5qhV9Vds1kEKdm7OvfY/69Wp/iaLL7PmThKWKmQVhFtO9bUhKx6qrRpLpyIFQ
vzD+bi80TjN2LeisHhuteOaAa6KDqKkcFzTBTmpQuUGXC2wn/sNQBgulN8BcoqKiycJNDOm90H69
XGRJ6l4kw3ce+64bulvC4p03WE6z172RzYf08wwjASQJyT+qBCN8sx9RN7jAygjdDZqshPqA1mAj
5KGxM83YJ/J9QIO/X+xyOwXTTpkXUAth4e0wiW8IbRzDdALBkzQQNAg1MvXyFwUlWbRiwNwSulfV
UbVZaUxzUeQ6lLowoiQpjBtmfAWaTuD2LLN4Nvqb/8efH8xTspEN2vzHRhoU+eWM4aZb6+kmRAQw
7+Lh4v3R8zY8xzqfMkiGi//SyC8PFjXBEyy5k9W83dDk59OtKjgtIuSKKbPIIPDZa4xIKbfCd01E
xR6kospfN3tXtuNM/k/ognKb83AwvBz+olQTny1URurW+7J9l8VpfEgDwhbbMNFMXCY/exZdP/vE
CtqTqIGoQzJ8Nb94FkParDlSVZkV8jq9Ao4OC+3RhIqTP3j/RVTn2Dyoi0/3QO0jyIjNe3MCJZJK
r0vRWXU5iulUWb8p7jLJndcamsytBqMHXsQLUFrIy13I2WJwh1Mo7sBSdYMvxl57NHfVfyzC9cUf
Y0pzcr+MnRW3r9s1T0FFlHSX/yIv7UDRYISD+uAFsM3WnOx1SfBC3tfoqKnJs7oOYLKMQj9arksl
8anxL/Zz9iWZ9dtWYkDFeBc5NnYxPQ11AyFM9se+SKS+pMdDNGS6HjtJLkVrzOoJQ+W9oJ+8WS9A
wOsk9slEGAsYWhQYcJWdq6nLJDVafmRzJq+OU8AVPPQo6zDEKcW7NqlBK2Qn3+KCos+cuuOGmA9r
oZWJ/bX+stso3S2YHNBc5Untj3i5PHdNKS86zc6Gc+8j9Fq26bVe8YEjBkr/eCCmekAbd+jQ5D/9
Cnr/fdXnRCXCVZUCPdLSFSv6n2s+k1Z8fGcSooVXXzPmA3Chb3k5qIWhn1tVnyvRxr0w5p4zo/54
43zB3fdK/gubIjtXr+xORKott2QOyBvBdEm1urpGNsJQwCAez2wp++zCbKFlIr31Owb8pqCRL0c8
TdJ/rb3aFyrgtk0xG7ZSxsI4ee8OXfPZH+gOZG4EkOh1sg7y8RfAWdBDyAPjRwPsPxXLm4zgyHGz
T5A7OPu6akyfjFxdWsPIadfRoiDkh7bInCi/dV8q/muN7GwgzrhnmVsZiM2vWGZmg3VKxpxG/BfN
sCxvMRlL5viUW6Y0RT5QvxKKE/+CspR+p7gIm+0xaTrpDzmwIcERjzzOt48CWbmP63g/vj1+7ofp
3RCgxgxSyRfOZWMzWKZ8RyYRlSVNRxex4frB+gjXadBEkzjs/C8Yrf72CZT3CFyyQaWTn9+0KC0H
Giw/aXWbuuRrm36X+NHJXpE/IZfsq6gtx/T3Da1vNC3xZhSQMP6yqgiaQ4sP6IRdNdLsaHRAjxKN
JRnnCfF3MQqEYUUd6hcHaItVxfUYvPhUtE0ZR88nimGRyfaDWi5nEFJ4w1wi+Lj+psRyvAKUWdXe
btpHDsDvDQQ+PKNe5QIWwYZFSiaTCOiHVblvM6DGfJ/WGqtZkT6dLq8iqcsgPb4d2G9KbwUYZtup
J/fRv14xDXEclQQ3d4GwKgaxiQaevJOh8VVh9TSK3vJOsEPcYqBjwtcSm7/9iBIOBskZa3CPBXCt
1Efjnyq5yli6GrSu4Wk8bM/QKW7/59wcvqzOtWghOTi/Z2MM5m9WNkyR/fiLPRikBGEuNBcvXxLZ
7vY6cDcdkHYmEkNEOWBRvJNyFAgLcXlwahPMjZLmsASfAWCZBAkwUccrul3UPNBC3fM6lnl3ZSsm
0T4Ucri8U2vh3wx0cnu4vXKUHRwKfMaq1Bl6397qvJNP2CmwDrN9ghZ6xw3KtWRQBhm39SY1ZJ3z
dSNebz4oplfrbpzDgjL0On4y1131lkcpzA308JP7UNWgfNeJ1/JaMC8eZwkdxB6mwHmMy8QZbueH
960BB7Rw2nbb/AoPDMp7Wtv33/e2/eke3UV5+myaUmEVgq2zjbR8xl2pGi4kAiIKXyIhlHcyOTcw
LlD7zwy9X7wH9tVWFy0AF7JQjzvtTW/sgO12kgfkAW2CPrFW+VVZI5vQDYIhn/aX4N3cnHoVEnnf
Uxb0VhoMx5FMNBS8WnvL0fy/w0v68r3EP+jNExlb8ZWvqzgzPA9u27PUM2SvnbHhhnky04xHS1aC
kPDoDdtNyO5x9IqttM2eSf5oFNhKBw7UJfYC/uIkYfQbPjjpRQbwuJfCoUu4bP9zEZym6LEBI7KT
mKADSqSGXeERFnDSKprmWb8BngGmEVik8MMpt7dDny+SUTxWxfCWvWvzHBOczVGI91g0bxzg/yKz
pXmfoOG3WeS/jBvd44NRbcink5ammWWbJXq0SFHOFtJfpyyDZfWP8FyTOTDkP4jH/r59YmJQH6KS
r/QgdSXEnqg3Wzl2oaJYI/28DCH5o1wUOh2kVORTiXSsoI1uk3HlBbIoPTpvrizobu2afTIYMwsw
moTeEBMZIeT8qRj1W6v+Yya9XMWa6/FT7SF8iZ6PuVCDAgGRDRdvkyKr7HvYOfgVmURE6bFiY9VJ
Wzma4th8aogG0nCYi+Ig69lQTPrH700p8q4yYJ0zTj5daTZhFAynYpTuaH31CJ2Iv8+4miMg4xvS
9NckwKtTT3W/10wKh9hLbfqJUkyjRsqMvI2YIBKfDeacmLy37A//gZywwFa/saNWoB9KwE3yw7+M
1OWqzMR0IPMBNAOxHKBOM0dDlJGP5Bpb3LP1qxVaK5E7yHyKI9N2p0xGdQm64m3f+/rEpqzOyR9w
JAvoIV3r1YySwOxNrNh4xp+yEhK63cWgyQnYlI6VAuJn2wAvowqW/cE0NjHQQp9lqYMSOh8jpuF+
DIizDWCwukl9X2o8VhBodc9EVKzW9+8GR/50UwibRHk6P5nOss7tkc4soQ35/JAhEUdGa4AkXEWW
OSmDUAwhT16Iu2rhLRxJicjEpl6DdlQO8/fQJ23uEe0ci/dvEv1wqDQ2AZT6v8ys6xXnjOKcVUSW
7/sToPbdD7FpL48A327lpm9203Pj+u/isnaFarMcdpbFOjuPxBnyQtO1TDfdsZi/LGC0Y1z9LoUU
JQ2L1sZwvZ9+vDDPo1PSAu2SfhO2Hb60v9nVAWPhYhOQMq47CJbgSfTu+UN5g7zPsPdeDLbYpnf5
JmTr3IxgHyH5GypTdo9IcILpVGNnXqVxhCxXsduxQPHc9RTGhGdcehqEVizzR6a0gWrvBDkJ32SF
yIxGgj06gStq8RQzGggkwfk07bEW4D97hs/d45XsOjCbKQzjbyh5o474+0VQ0gGsTzw9Y8607d3a
IBlhNXdWgyVQjLCgQhty4OfOAnyD4mf2KnTpPwezLEPKxF8Lh5AT3h02WZhS8OmghmrF3RJPdLvL
RGrdQUX7k4/VcMzMJ/1rlqlUx+E72TkRt8hboegIy8WRPcpEjz4jRxWzFUNbXLulBc/QSiAC4qBi
ixCCqNRaMMRo2cG35fUidn4I9QUVJV1SdpXLQcASSW3elxKqEJBox2L3GP6vKZwI4ftD9joiEL7C
vPnLPbG4wwKsVxH0lM/bfpCv2duN7GAfdVCOhS4wMp7Ntrq1myarEb1wXwP7JjZ6nsyF4XSG/4BI
d4XdqLmyHxHeX9/B4jyEgVd9G2n1l3AcLoKAt8Q4z+tgbZt2EgqJg01f4/tBfKiKeaPiGDJ2Z/aX
8QXOmlRvl6blYbA/Cgh48rhlphqNcgMapoXoAXlR0zZRlHr5WHl7Vv9n+SlCe/RkC3AnEP4pepfZ
8clCJmd//ttWTDCfFpyRjBaRaO77PoQvnyYklg7luBB9f82FIwJeNSJtouuI0MJEjmhsKB4/qBMJ
xEM6F65/FEnliJWllvbrEnhTz1wGSb0Fbge1mZ0xw89/gpzgP9+iyiwDEtN6dwkmCNyh30WnnEpn
HsRvr9BVQdZRhqq0ZN2osUBPqKKN8Evr3YIcgw+KihcyBHhYsluOdNKa5GN66BhnA4sxaRHq6cRX
NUtpQD/4yovr431dwsvthNMLOoUsk7574xSUUyBVtOpbG4b1POwbTe0BCXANgIwjGJo2pvzcQaeN
ntfq1GV4AmdwZ0eQ+VDTjJ2WemjXYRpQld0Cf1hk5oFrYPSGihWVXBxQ4zuV97w6W4qCYSAb2mGH
HNCYs0hDNXPM7wIy6bMaKc8RlS/4m3KCzjk3LjbweJerIZfaCel9b2eEb+vIkliAfpXj37F8fAQ1
zKjCyfEJve86pTbRM+PyvxaquKRBFYXEHb2rX9LKtLM5JHfjkZAXxiGZ2PeHsHVkCYJFCS2ovRUp
0Zn7/1ir/B7oYjj8RrwK/sODG2pbIxBl0G2AOibAjIQfKYMzo8p5N3R3vwoZXk3TTAtKJeYJE+oI
3bg+guE+YxzXHB+GsXWQQUbeY2W+yhTAwfRXGgg4r5whhlMmx9tFBv4KARh4Lbg1YLN65lLfCFNW
h6lj8TVCblDTdJHmJYL4bPkqHLCmKUedUnsWbh+lCQAsrRxBhvRIrGj3GHJ0E4uLjdAd5geVFnzS
FAmDbKWS6cejOJGlftVqHO1Fz2K5DPvPgykAMMyVSoLKdlVUjWaA7Nu8wN8LZI0O9M0gvrKyaLIF
r4JgIR5sQuiK6WX5bcUZjAllJLsBK5Aa+a6Uvhu3HK5PY3ZH2sn1TR8LZZr2gO2zZ2kaNBEgrxca
AmehgzTn5Z0iqgA5o0Q1I3l76djR7VWW3Vn+gxiT8+IY7oph7K9yELctN8CdlSNWgnWiG7YkGbEy
ag1kmcNvZNDsQCx0/rOQ17vybChYlXUAtTD5df8HjJJ2c9UYrBqKPJl4TtqKnVCsB1nAdq+H9CcI
xrUi0eIVAL52XZuo4zwrB7FUaTEZJnCkXmhAevVimiW9jxEg15Wl1zxDs1mCrwH+jN3FeeQqKjrT
3rJ+KvBUARz3lkM7J3QXksS8fIGPWKCJNBhNs38p/xFaQD5cpno2jtHPY31pl0c79D2gxBG8T8PO
aNjsjOhgDA7dQ4Uh5A8jw16rQkMnLjVDPTUuUDG8tR0qTxbbDtFhx774tjcbSCcxrd4H4j1qVsuI
9jk+CxVg9MOqlMqS0TfGZnG+pP4otW45kj2oVepvbLsQhO+c74tFoycOrBRSeWnKSMWsVdGaR7jU
tzTuol0hnnFjtKigMBW2KF3f+fxkjo5fBAIWemJkyEmLB0hip/bTRopuU43IrgiieL1QIGB0WTRg
Uz2HAAti+qetZlcYde2mW3MYet1wGW56mRn1bh87dsNkpDcc5Hi6wgf/Zo5BdrwCUERuBaWnheN7
Qs++V9HgasDbajGruZgRQ68WByct3FdLIOy65MdLF+H4/sJDftagwnN0pMykG/8hxxMQsL2N88qQ
3EKeXMoJB+jF7He1rcICokMbMkLAax7549SK4x4MJdXurQtEMhxsqJFIz6Rq5CgTbU45SkhEayQb
n06SvhBc7ofLXfnGes5mgOiMEJxJOzt9vFp4cm/D0E6zwuQFhwXweCKDKsgJOJCXKjYPDINxcu9q
3PGYJFlmqv6oKT1499VFwcprCbj1SyYRVc+Slf+k4Bl2g3AV7e8xQw5BTDSdHafKGB3dySXescgC
va3lKjDSc9euyd4RqmfsMhUNbMndW+DhPoJndtMJkcZStX1g7Xk2Sf4wui3gjiOl6sZ1cV6KW93G
cWIoF/b0pBnP8QO7u6HuAV32E+EOYROSayuP7NoR7WJJ2ze2NBXwv5xH1kPfFWGidQw1bDOfkQON
7XCVyb5H6TWiRRYwYtF5qVvpH1y2VKFKwfHZ+KGo3NGxKemIhilog3vhClrOKZnwKGVY26TPNZL2
nmHaH/2vmmNlGigotKa22Nm+HgBct0bHiSwB20066nV0IRg0bFBti3MfU75EDzlA5Nv+bwpeWpJn
E5CtireEYG/3jcOBkvDSa0aFWOBlDInvaYb5Xui7JC71JgqOLpYxeZJxe2h51BZqAWIKc/fayZd9
N60mNikbxVevJdMugPzbtWIJCrgsuC61dZzQButxsPmM6/SafdM+LIdjpl2Ld8gP5HBo+WC3frQi
1wVoL41bjSoz2U96LDzf3Y8ccA7SNkLtVtLnIshaURG1gMmkAM1eIFMQkOiTh8hNK2p08kXrL/ma
aVvTIO9IHVIzzHlD0aGloVc84hwVzxzKBSQqFHYJRbdXgySsGvSkzTYsH69EMrVWar5R2lMwss0C
1C29bBrHzuUfWUAzsk+MaxsBESbIOrOklMQn5g4ih/Ca/0P25dZ5Vdri/mhQALeijBmH0YECsfPx
4bT2O+H0sY7Z2cxGQ6bMZ6MOZbNRP6imCihtV5JoK6+y0QsGZo/bwTR47vVB8COObvCZpaafGlaQ
B85rKYdGo/x5LOoWlhM9+65UPTzXmvuqnFsbNv94uYV+neJJDrstLV6JpmCNXuaCI4L3XDZCjFE9
IrKkjiF6w9oMqSHthfC3MgXKnElna+dbZXUdz0U84eg8V1TEPLd8eC39JM+SI/DSey5zstv1wOWO
4gG6d+ydHi+0UAysWCSQPMkIN9mRrXT+jX8YzzOYVzPwSyd7GdZu41QIj+lv2hUDzRoyomwWHNQr
LLBdXUMb0VtS8pNN09s1aYxuGdx7nWS3NDqf2DAEQnOIVWVpGx1I9jdXOIF7YFNcpLqsDFO2SfSh
XRbOD3PzeesejOa2v+cSFNHsY1DkSVrQtvLzIqAVlfm7ag/n8gOrEpgBdDCjY7PNQ/xXgJNsPcfI
z+5QWuLz9rIVWB5oBOAa8KZIalTArMwkMehlHgSNuaDuIQYfBlWMhnR83axJly7vU89V7XK6UBIW
v8zq87ibHD5tlOzA1gT2ZQaE5nzjGdJ4UWomSin47tfNBHR11yrq7cGtcm52DzMxkrXVk3ucl2AC
s9pwYQnMvMV5TONmqlzgFncgjQ/Yml5ZYr7eQSUU63tI56b6mafZirhSXSIrtp3lvDj7ylMMB9s5
5DcIGdD04FXVlTuurzwwEyTCRx2wUEVslG2Y+GgnO8lyti1+C3lo4z1HYkkCJwTf8HWxDpX0Or0u
Usu+YZYxuz72nfIKOXSrX9Ltcy0dhOe5f0yRQNfLI083Tog+Ev3+1vA75HXVqreZvP8uGUjRacPX
UaU9H72DLEbLFHCVwT6akoBZhoyUcReXgJs8H2VmDAHcaH5KY2HrBm3vLxrajb+KyQqsHsE1Ugkb
3nbb0eBRXb2FyiJKCPdOOZQ9irlxpG66qVolFIX5myuzqphf/3YSOmxtBy6DjUYcZPN+CgHIam1+
RfVK/L0mZH7u8WWDJ255zJqaGTMJo387imG0+iGgwuNwenjZhMVKcWahRpxhUCzo7esZckXT0ceN
iXoY5B3DUeuK1dnAVlN+zLUr9e7cwfGLlrSLoJCyvFMy4Yw04iwaie6INm7nSWJp6l8rW6l3XJ9w
/AfLwBo1vhKKs/Q9Xwmh9+1t9YUlHQaOJPDkIpH43JYOz+yyQB2RW9DsG3cuG+mn+Vj9WVMGboNM
vRY8lkQgRqUZmtrIb5Rgu9uj6BdUXQ6mtSO1CAkL41TSpB384Z9vDOX5mn1E3sM7w49H9s+1Lqkh
6ZWoRikrOeS3yHUj1FJ/DRm5iT7eDV0vwfwlsO27Gc57gDJX4cy6PVxO/++sl5VZcsgwDBXxLbln
JK5YKqYIKZW4yBqg/10f4pECj9wE8p90j5zQ1fqvu50Xq9rkh8cn1tHwUaiBKZqjudZ092RPb0QF
4RNqNXnv7TY2Ta0gyZO6tsRmK/lURQwDpjjt7tzjk/iBOsky/6RtLi3P/7htADOZldAG0VkS5doW
Bl48c7ukQkvXGzUOqzbhUxZcViA6BB8AQnEWYt2DJoHTtsSMyVEhascr3ES1Ons8jAFiBUiozkKZ
rTPioWzvF4yIG/26WDxWgfQFQXu2rr0uIVPDa3ZwxHA+voew5PvCmsAhoyRLL9C42ESEDYR0aBPP
HCyZKpErzZXz8k+hqQO4bH6zCtL3KGrbJMsPUaL7QulWW4a3tsL5sztS8S5NLWusTgJnfcsX9UFf
yLzGgSshEjSRVCwFT+4n+ANauDcEEMY83LNwSTmHQyuktLUX/7lQDseP7oWysvawJf72B7rAP+B2
GlEDfZghmBo2WEy9bv9bBPRg0E+MKcVds6Px4SqZkmdzfCjhyrNWWuC5Vu2GupQb7FA2x5zu8l7O
rVJyQl5Q5n943gWm2AS0CgwTKQXGDKQUWccyGVs0B0w8tdMjRcnDc2N/PoqkcDCCxChg42Ce73XG
JCqG9zVjwxG6SGPx+bvdefVY3RcYK2dtQhMNMNJER6p0RImpxIflsZfmy+gcv9Eez2bD+GxBAeT7
JmqTI15sha5PXARLQFx8nObBnbnloIgluvuzztxtywMGPcc+5TTjPB4u0qGdSSKYvMxhhGmsgz0l
6vGM1Z6PMEznKgATJxoIIR9tSPQje4If8L5SVaHAuXkzBvrW8f5TkjqSXz2c4MJDqe7JAhlBkkzo
s5VGbs6bDOoIpjpFpSQ2h50rC/tC0wS659olfy5CD5hYFl5HW4bC0gLiA2Cc/zatCnFQ8iK2VtWB
S+bNU7ngJW6Qtcp8QNz5FKb6OQKPpj0CulmykTxrJ1J9q6iguMBmjK97+5mTEbzVTAFLb+pa6ZV5
fxaL6mORjC+8p6RS4TJ909aLqAlPZ/QDM0HZfuPfwzILuwjfe06W40tppICyl/4qbCrbT6qBUEQ7
iwFvT0DBNF2VG5bEhNPq20VtdaG1JAhxWTCGG3qgl35welLF+NO6qu1zrouFU3j2u1kcLCCHCywD
6chzzkSvoBt1UX0OSR1/pg8szg7KFkuvp7sqUA3JzvepJYs/+O9f1RcLvgluTZS/ufxhu5kIykeX
5B4Crr+QUIgtPs4DxFnI7azN8LsfVaXGOlcEqXJH3XGrl2/YajrtrP4tBVvFJI2NkeIkKv4vVmCW
hvqNi6sZ5PefBWQIerK551H56Xp33D2qvtwH1ZEZWd8/8vSEhJxHtICrsljj4OmdnytABo3zXHaJ
QmNAfidNvZCCj0WQ2asBb2VZo6QK307eYHLx0IzobngxdDi7V+qA+CWAxcWvELDOsABZW4qk6pbz
4GyJXNOXsgLryfxe4VyimVHK8uORrq4Ds9tOgxVhnSJmsYfGqFdbKBFEM1vyk6xYscXUU4Nj+lF9
AcYGGhDw+bm7XFXH0tVZ6A73S5PqFSE6/IwtDs5+SijUtJPlZMdSgZ1nEv0ONuMQsMppHdw2uG1k
EU38Ri3Wlpt8pDeoZRsIWhVtHD57DqvykZvSA7ufR9cnKaz9fhlpL9nbTPpR57j207ccTGYdZXSk
Kq95msYBDO9XGDgIwwjzvDa2nYQwXcx2mDXgSCq6SXM7ToIcBYSBSG6X0+KxcBnzKxivadV6UzeK
LagNxsIU6wdF4YzZQIbATkSe/h+DtRG/r4umEf1cI3lS4gmPzgQL+qCvIm+sQV8lNN4zDG4ibOBp
dV+1ri9jzRqJj6I7DeBDcw762KCnGNA8oHhSipfZVaPZmWS5zqAAhOndQyYz6ZBpVAsU2rf9Xai/
vG7p8k6dpWh7ROh0Z5wvKEeeAaAL3BgU8Him9pccf+FtgGkBulvAHm7PrpuellGCa55pVKjDbzHn
VSjoV2rEaMIjroiAFfttk9rc7BV5XO9aPGTQNESIGRi3zmBoZ4WaV+HXp3ef+grQeiZ9UfErLezR
cZJWxrMt1en+WLig5GGX+henPtd+dYNqZPIVMmP237LrgcXN27UCDbuF8VU8uRW+GhcSWSGXNJEx
NLw3GGqO2PYUq4mZpCd/uTQ2nCjKvwKKugwQm4brSZVwgTIualcHI0yXIjxff8TD/Q+QE2p5hum2
WVXvrZ00r+51H4ANL31X3EG20DHrkIB3IDH6iGGn1QN1Od5nVdxnwqHuBs6KBL9p3cMtfk3gEDdY
d2C2IHZEhusRrAumpw3Of9t7q7qJkqrM2jPY9ZF4bFJRVO2gVTEN39Ad0C2okQ/uF9r5GUsq8xVz
6YouuTO+/O1LenULdz9E39d61nLhzP1PQk5MQYOzzCYxglz4wkkzpD2wJXXp8eODGiiLj7qeWFh8
jwRBYKbD9avuR+UNnTQvK6oKEClugC+MYksmtnly7d0qX5lYe6RUllx3inKWbgCBnoaXExnvkh5M
wkWEmxRzhucR2dTZoxrptXA0+86nzafymdh90OlEdM6j2qCMT2veVeW+VH50xcP6oN5lpUXdh2iz
hgQZioH5T9N0YacPkCZVrE09COec0va4B5h53I2t4WfO3B+X9LdZFi/YUg/27y8RDo1F2fx/t9oD
CcIKQk8ygWJukUd2hq03XOYxaCztokzkOYT8kcbW0aIlA3H/c++DGogZSdAO3mFZK0uOvl6Hox80
aQbj5aVWSpsZdRhgeKaIGlB1ap69/0svRkY4lpsrCYHGW0t0a/IccGYxbAjQDRvdUOYJHyBAasXw
HaZ1ZjV7m4GEHh/V1l/OyEvfMVT8MZVAvhB/7hP+jXg/VASZ/22+gLH7EzwRzx7rUnqy+18YJRCJ
9ZhwHQYWHnLc09ONg5QXx1i/3n1IhSMsG81ycCcT9fobXkYxrPsVdmHNCDosmkuRHkY8SPNxzAT+
C9tUoURXAcfebLGnyfM3ncKGY5dLtYpKrpvRNGXcRa4QxQUBz5v676vpTA4Dh3l0wD5iIZ48tupQ
bWalpSKG9wo6yfTDisbzSHfFPk1z1PornPKR5mpefsq/416qb/p42E7BLCDQIKmeYo9DgEsZ2I1V
5Ek+6BFJlnFqR8s7dSgH0cS9upq6LUUb/JNhHoYhOSjhWX/C9XzJWvXyIElsTBFNW+JFf4SA2RPd
x8ekU5Bfy/LK5RCUDgtDfvkraRGIEKhrU2BI/BW4p4+ZM16W3QgdzReSZcdj+GX6JBSLa2QDgD6q
hepWjnBL6wBn5yDfn/dhJQFNvIJqHqJ2sFwfsVMVduodUSS1ux9WGyvXxiNhG2OK5exUzco6Q0+P
QBPE7aV9UWB02CFO0AyvrXWMaEPWMBF0HwAC5Jse95yVbKAdpBt8mTpImBuvU6r4b3cLMInkZ6xo
/d/z2XPTZ8W/fVb4Cde02SF0QxukXjuWCu9sE8q9Civ1nAAB4+ECYQxMM4r1Ni27dlzAQUsfoM7k
EBmf8UFsuNqr2+jhSP8Alj8NWxQ7bZ9Am6vnAT73cAxm4K3X1iUR3ILxL4uvSMxO6kVlvpdkDt/b
v4Zyp25oFSuIbr1TVjCD1z6yWH0Zf4o6Hwv5kRfxMr6IrvEJE0vn/i0oloBXj56xxm2LFbXktND8
/7wMlRHP+7PnoRtkk9NVIYVFwpTvEUK7PejRZEzdDtwT9zhFCr1dTXmKbfrmdqwSNGviHE6FnH4R
JrhuhY0KVYmFYQcViZMWqFRkn37hfG8m3LpBm28+9r3midlIzkBLnUpQQ77H09DdQtpVgJQ3ceiv
CvlLnv+AKUIqRNJDk9fLaBPgBW3u49UEEaBfokOggPhxRbtxcfPv4lUgLS99c1LZYoUyMM21yEKK
1ulZ2g/gO4oqa/vEETXTcoBy2UwsLRyOakqBtW3QtnI1bWY9juZL/kfsfROcvOpr0CxKRzS4UPUD
WqT7+smP5NOmQKJPPOwr3H6Fi7unxgXXdAOGqCf014M8d6FGSH+7dfjFiJ4d9KtpB+2b73W73twc
CM6Ar2D+P5SkSPrBxJc2wa0o1pwJkF5Sna9ro9ZC/DsEqK5XcJlqbUkk6TAyDyYjOQ+DAo2e/gHx
BKLW7ioPBcIQ3JMtauFhnWbNplUuZzdXQOIw/PG0e8CtFZ1TXH88AuKcbDC8buUHVjnCIEjcyqMw
Wbu18Ur42suPYHzVrTBEh4p+Q3Vbt/CDVefk6XmXztKkZsprL9jrvCGPZHllyYKB+3HnY8z4ZUrY
rCfQ00EN9QMRvu3iPbv1RYGQTA9YIKQduhTqus+wy3BP2alqoetIt/3iCGGbD0KHOtJMKeMuaXAi
zoJZBdzLEUNO/1ACwUdT3MktKdDdb1bKUT9dtl/jwIIbsyoletnx9K92Dx8FvsHpctQ1/NILId3T
2ys8oEb6WZqm9yZyr0D0b+Xyj5If3+eeC0cOG8ldReWJCoypBc/uVjymjtVV+B+cMTUc6THV6JyG
CB7kyY9cmsn1cwQeQK1V8JBwRXNJ47di2TUKH+etUrTak4iBWZVDK8OXluO22ALv/r1A93+dWgdm
uKwsz9p0aGTG/AXxlBdFHMwZ+gI/zE+VNtScOAYNaX6OBhZ4DOu6siWIaq+FDclgwWe2MJ+FSyA3
LHHIKvdJdKgt8kYtYDS/lkvRrU1TZLK+nWVm+qPC3YweEUOf3G4ws/YY7hHRIoRllQCEtlduQAHF
HTDQqni2MSxrCEPmEtNVX5K6SCHrQkSHkGx9K/6yDn/mw7Mj8i35WTUwQ5CVIG5c4aIb7mB1uZgh
paVZjE7xClBrXuD8FdM0BZiDNbp8yLBwuNKFvhX9NRAwBWeqa50EVcTULeEAyxNnKZCw+eJZrewj
V107IMq+hs1JFjZX8Dc1lWVaVIuXn7hZi+GcVK++gd2lvc6y5c0GRpo9Ec/AgtoNAY9bmIQuZRw/
NpBlIytBJm6u5RdC0GUIkraSzsHKBpCsORMyV7nN+l4W29cR5LusiS/G/MisqQlTKoJiRVKxEvHY
s5MaKOOqHryHeNeQwU10ToTxSQ+I0DbihqSQ1lhnQGPegtZi+7K2SFErE+TRPMHM/rOXJ3tAVRPY
HydkaWF2EbT093Ek7QyEsDhpqLyqPFRPbd2aoiry35QGtRnRoK6j27f4NsUq9Z2cWWQpQz/t+Ynn
K2sjH+esjadWOx/TkqDzpJ5RQgiF8G29kh7dx3bA32XHBBLfZpVg98lhSZ7gPyeBWMqi7RgHL9wq
0/cf7iXlCpB+GdUa5LZiEPAkcHhH7GzlDKBzRSoeq2w8vzZ7IYYH5tOz7xRYjHpPICTxMSMx9K8n
mMckXM1/iSpG5vm/Vnj8sRcsBjMnZ2HCUm7parVl3DJsN5Hzdt/asl7kb+2Oo6w5fITQUaMdsjWH
Kh4kxnZHKWCe3sUDHlG+iyb2fwPclt3tyCk1Kg4EKschhKLKL5o5HPTnL7gv9QkEOt9JcYn5A4su
75+w1gIJqkA1REZdAKL4dwwuHNWTb4r53v1wf25SB4C3Vok2fq0rEoKnMRIGu+/ekkfy8iCTBOtI
RCVSCb037VUqfcEN6/qtYoQJDloKKff0mkr09NeKhgqtg42sCsilqMXU2kdCyJsMT5/gfcFa7kx0
2HhNOkmenlw03MzuYQ6I2XU+r0vZFlTaUvdXeByRcHRB5nJe0NINrXUZdcUTW7aejGA2LWGfJS70
xTXOdvqHR+3tDl1nxMKkpi/q7bKMpr/Fo4KUKjbVtSLUd/uVPeeVx6dA30q7G8Ld/NNq+6fr/Wd3
TRTHRIDB/F6VP9rKaFWTuH//hSkFxN/fYXq4Blsssfylil94ysbm7MHy6xjavSwuE/g3aNTgARi2
d7XTv2ewMqmlgJeiOkLTmZ/1JeKVk8BF+t7qOz4VNRxwhXUHc6EoUgTXnO6CEiWB3C3cChUaPxdM
/1D/dgAc4QDCjJsChhAdNCeX+6bo5pX4P794s6GOQ09cnwBSCY+GjlGj5tpNDFh7REy477gJmKBh
LxM8tspmLg2pXkFYEhzv/XjNc0h38slQRKv42REkpIMd9UX3Lgv9UAYsoZWTyHTmpqKcrI/3dbDz
mF3KFblgP0r6XZafDGruJ8oroqV+1VwkNmj5xcGiy9k+OziDuLos/Bux56g69+ZraYlzBvOuVpvG
aM2HbVqNfwIz0O/lafRU+9lzkuzIScQoP02sDz/41/a0YBzHZHjTtdPjvL+QKR51Tp9dbgCkIqyA
YnBnXOWX5U94o4dyIiWaz54gedV5tnysHi3cOBZRK+pMafRLvh5Nk65+DHm5f7C2kfIai+ltvqn5
MgFKuugnNoq36lzXpuLtb8LyCah39aAgh9W8OFE0jLSOH6ANRip1m5mIgDbP2x//IoqC4nnk5AvG
Dx3pZnGmmVZRELyTxw/5c4zY5nyCefBenMcaG1Yr4FYOsz91GfcuM6R78B+DvD8qRvmWKEJGZaOV
YjylQioyM/k2NbLlXpk6gj73NZUC43qmoNYJ0gzInQNuep8/iP5a92etXg/WYHmPDvz07yKCFKtG
QwC41dP0cZj3Bmzv1hbgJHDbZTGuW3xn/ft7n7PFiqu6r4/phvLqKHpFIeeXKok4CF8vR3awBFxd
pGxGCKCjVETWrnR6JHDMEDuIl1s6ahgcHO2ecB6bwMcXfMqnzMtLokIEiJqkxSkE7CPMRbKKHeAh
BHA4Ira67/EpSLO2d0c8BrTv9JmSqF5w6Ie2FRZpiGpM/ymEFuE2IMCF6nvXFqKnma7vN7fKumJu
ULhGnNyj55YHu3pJXsIBThgdTo/Y4v5XbDHDQOViBwyUJqT+aUYzMXab7OIqaqWOYOFoT01FJ6sg
Icr7AnAOyFmlTk8JPoShlYM87mOGs7j/9Bf5f/d58RIglgIvrB+eJS+XMZr8KKE6a039SYwkLS5z
sBZVHC7C7hNGc3U7aGKjdQoGWTJu1tWpeeI0gw/j7IRV+Cvj8bnNLUZl9vvKC5LMNe56s9nfg47M
QGIBeSmMOcUQdHDzH6UBb1Fs1Tb96ElJ+zB5jGrAS+/WNqp9TS9tMqVY8HdPeyguGd61e4BG2lpG
tKIbi4kQNkbkjOxe7xCf5jEEVoU1GB/PNEFKV2EheaVmIouPS8zUTq4eXtz+RSjyKlcNMq1xLekt
FLj78uQqxwHv0uEzamPmobHKRtPyTw3hx+7skHGcmrKW1tbegc5e7IohtKp47+2HXcP2I8RoawnG
ErXqb3ToFQXN7BNI9SUA+qPYsmfP464jf041iJSlGmfmel5Z7v01k1NvRqaB8piGuL/m3KTqfnig
pvFoB8qW96pEXOcFJsWjNzynlWip1LmRm4CRQIqIx120jSKwPfWhe22xBZeickxPWS+D7+rZau7p
s7DVgvkAPwlvoWSbESeZ0Zdy5FV+naDYk+JqlUm73WbnzYgnyElZdWW3JXfrtE/6aadnBMiLOzHu
Ltm3qgkdktLB9oO3SU0MfyYnI4CLMQI/WB0ZWqpJ1C6K22hmLLLmRQwauR+xCR+5fQX7+FdXVRgK
/VI50TM4qXArXwdRlj2Z9J+sFhvrVBdI4wnGqk8Rq2Pw+tlrNZLQL/hpSlmkYbuj++pShB7HF6p4
H+M3TZNC+quK1u4W3o3y6JlZdkMbmapriM/qORBt/eA2AXFNtQ8T1ltUahKK+b8qmq7kStObOoUi
7F00FwaxiXMmjz9Ws6Zndbo5YJD0GjN7/wZ+1bSJd9tPqBD9EfTt0l2+/KAb28SK6PkuXbEZ3W2R
DAY5+NHx1CA2HSrNKSFncyn11j7wvl+HcyztBrofFQnFBe8R+mFcLOvKn47rYUZUovfWPv7jMLeI
NqOtzX//32C3BxlWmrKj4WRymEwSpJ3M3z+NmGH4042sTkquz0SE1ViotPBfhsx84qCyqZVQGAjg
o68YrMhSPMBMZb0cz0Biyy3Gg1RQEm4X+nihjYGpjMzifku9q6WWRWncDhkvI2NtUnXS6gLXbAqW
9w8CLinKMJCzG4qIMaVu5YCIkOGDiXK0w+2s0DMxAqUGNeER1/nkarVynMcLyFHn6IiICAWZiW/r
O5m60e6cvfx5aawMSf3DdD6zD37hMvP3sj3y70MO7ug0yuW8LBr1yTdTmB1XAdlXkLi9XiS254RI
zFW/WiPUvjPkKQHmXaz2JcXTXiHVz1luE0nre/TrG5zNJT55mCGTH63xWDAchcpP6+IkmjquPcnv
bm/RK/TCoCNvccCwf64ec0lZL8c3z/bqWmIBl71bqUebXmEmgh1SS9RBYqgx6yporSqAIOuhUepL
+CwqSChTkdngXYRt0PJoGMQcluXfA4rQI2cG6bhqY6n2SYTqI6M2jlpmSvwQzgkdup0dKwAneSyS
IQF2pSM/nDfbeVAZk76t6Fo6XAOjhXB9YPK+xo06kEuXoMoE9Zs7+j7IO9y5Hw5mFKNm3i0hwC5U
ebDVgPZ5JxhlsOeDHDTztBpkb6AnuLm8bZvfTytJUiakP12JwdIkEBtnnNiRqZgeZYf52jYwCobG
rsYGKkbOLjyZRYNieeYNSmIlTXL7OtgW1MQ7fJM7Iy/V5ZCn+C5U8qbI+4GCPLMYxsELsgK1pig9
9CLtFNL4Mizy1wi0BN9+4I8L/8E90zZjUfdHst2k/5kBUVnN78GdbHuEc2bHqMbzWkTmU29WiAt5
3/1cNa/jBlQaQOmtC7/IAw3LfYtv/x+Nm6VovTmivr/osicJCzo0+4vTwEkGUtz8QK9HPlaH6y+F
Zoa6KNSQUqXs/pJOYZ5SBPpygzdfMy+gwoqLNLzE1QwxVOeQoPQREwCw0+LmuJUYmkczTzKDB74Q
XR6QV45p6jd3nvjRi/gnc1WVWj2b5G5jkSrjvc/IbfmiKpRWOkNLsScwpJP44Fnh2oYfktKYlg9H
FC1Xl2lE8MCtFp5XPDEhB1gy728Y4PUBpXo4eD7zMTLYBuXDrjBL4XTcB/ssdN055Vs04uAx1INP
Sld+Dd/j29XhQ4VOkZjwK79s87WPxZ307v6cMi24T2oaR05tlWipSq/yquGE2zx0BSvvgB+pSLvD
Abuca5EXW5OiNogKBa7xKdESAdNpPTUksTa9kOdiUWq2TxozoVkw1i4qXJcNctQRkPehHra8jnmW
aXSXDvrISURjzdralg9k/0xO4W1gR/CkorlEhX0CYRxJzSiR4h/vGYIGmGZQsh8CuGzN8gECaR3d
kuHkLU+FMgu4bMz5D6JF8t+ufRGEEiOQ7yfzvM0HAT2abMUs/SbxLVniWBzXVV3fkbnsZkg0PGtZ
aDaCGDWlxAL56HC+tbrsIMJ2NbNo0ckYdt2quN6dsuY//VslWUZxHNDsaCL0gu81EEU9/Ul5PwZG
Obi5vfq5UHH1ylPg2UfhZ4svW3f847Nu/ZttMd1PnGO5T0yzhYoOUTBcNiAKmGVQAcNOV+5DnGio
M0lgdywbKCX8n0Kb5p5FDWET/JHNN1BtoMj+UcSTo2NExccvz98ViYs/kWmZapXwjLjWOVCDTtVO
5GokZZCD9AHnmqTyWi866WfgQ3Jr7c14sGvfma9cn6sMekcG5b+jri1+DROpS9yShuQ5nvvc+Ju4
nyD4JuE5UeaGie2ogk2bU/CirYs5eOlXPbg03+MpD7g49KYfVRR+0uzDcfRfAMt7kKopnpGJnFGL
cYWMUy/yIKjaBMC5k6VQk+K0COiaLZANufHfs/GDynmwHwIZ0F8a/8WWoXdKFUfS6ryprBG8LcbC
mDQmqJLTjip4tSc00yGzB1qwc7/I0YdPtxGjwWl7RJI9bL2kM0sQNHBTnd6ZwwjvuTb1x5ie4l3o
pDCRP9NShpZ5DEcK/+E2fMqpVN7ncI48uJRF1EBe0nPjLdzs82s13OpQ7GdfMYLVqhPIe3GCKoiL
ZEeNmYCONNfNu5AsRCtEAAHDZVnvYF/6ot60qntspxK9v4fryhpjtiEPwSg5H8+j1gmkmCh2Sdv1
kw8TrePEIwjItYW0qpA09kLfFKnXj3/cRa0yUaioTN+soGYmVC+D1Z3tbeP/90gJDmrO9PXsERKq
e/CsG49GcU9GCOv0ULpOtR5EixTp93ri83rZzcczw4h98XWFIyP/O4qd0hR1E06puxSTyxJ6P2i/
PMo74oWQctm8CekwnL2tHmbNgRzaUhO70psTU9c7lyxpL5zR5AHwJRaCX0v76GAwWLKMBWSj2bVx
SUzsfDQV5Q3fqPk/yoBy9t2bYwDSOouCRGKLaPJtQTwkIplRbVIuun/RvwVVUlFe6tSSgO2et0x0
PZ1Mek4xkY5Ne8B/rprUNYHz17KdBGb48Noh8e+ngL+iS9hXzk0lgst8t4Kg1yQ72QBD6eh0MVX3
WdhHpXA5t105cECJ9YPRJ2k5tTEhaSIcl91NfS+K0i/4z8EkNidA8ZQrKNrxG9EsQWiaUGyCXpOz
Caz15elJ+zKAMcQKd7yjCP1R8yNpc+v3E1SuU+kZ1C7KbWzqxla1yx9ddKpvJQVkwII8ToomQ2wB
msh6P2xQI89Ml2eZJUb2NEEcxFBE202zxZNfWYgUtADSpgKMNlrM66AxCVhsAXs4U8NbpMNrMlQx
wCQP6sGwrsxe1w3KfDJ50SG0W0bwBh+q7jd24h0zOZhkFsXaHBxM+HA9IrJr2p5f4fNv1tRRy6i3
tyjWmYv/6byQtUoL9WT9PMRXC82tLid2uq7erGYVCftHXA+AmFcS3Et1y5FuhuxqSmlKhIkqkpju
INw8mwXcAHDoApya4Er9SqKWwcKT1bFcw0sBwbAfNcpO32nYKUl6H2s3QlKN+Xi6cUXMoJxtkBSk
e9s563f0iA7anQN3SsEHe2oAGxfOoIS2BYrpBPoa4BBiBMsD2YmJRh/ynrea79PPpdN8fgaDaswj
fZqOQdm+3T5l87x768nqFEeb3uRsTv4ZDEWUSjMp+ti+XaPMS15IdSpcIBw7YmvFRMwNGjSEWuQr
3Jod9sKhLEpHhiDSDX4542lghfD7dWQDFQmfA6NpLsRVf2TDBa+6MUt/zNFJS3lY5fTyxKjV1vVX
B0RGgfumarE3RJy/9N6FSFoC+J28W/pm/eJN1+uxWqNFAbsBPGXNmfpVOdB7+pdNi2J4EiEURglc
DGQjR7q0zLIl4htRk264x3oblVhMftzVWqr9BbvTcoJ5whPsAJC8ybdH7Gf8cz7KWgk1Hc9jAALf
DVJb+MEUlD9RsBdX24vx3AB7ZDiIC5uceVHTN94V+tGL3te1atxDMJ2WsT/0MkMdb2XfNPoLPDsG
5x0w4os1ptKa9k0R2Mr9roXLtVUAdlzL37yP7HIRBAnmKgW4D8vjItvkn3XvfOMIpqGBMkUFW1G2
5elxi5pu7gGHXr1TKm3ZXeryDi3l9SKdAy3liu1cvf3WeICiJjrGnGPlO3PFEBciSpF2bnd+m9bK
pxP2itFkG46J7NozeuFxC3W8s8aH8jFF0Hs4KjdUEyTv/mFnl8X8BvTCcdZFXP0jUHauL1rDpFKr
6P5daLx1pJK3ac8tiHfXIL/aRCQq+l7Np0J1N+qKsT8hiQoL2cHUFVZLqNNZhxTpzvt1x8jTwY+0
nba1N6Mi/mhpLAt7/OfizAQn+EVkZQ2q2wEvBZSAIcQPIg2HLCvfYPhdE83cTiTJ2evfGNYn6pgY
Nnfo3XGgEwymO3j/fVQEtmFsHkdi1mPcq/vBtYK7et7D92iltnvPq6IvlkvA5meXv6H74rdkKddv
5ycWEoVsK1SRvHiB/le8kdgShBKlVW7bjBzwtdspn51JL27d6PexOzrBRGwfn2DwzwckzDflJ/6t
xVyWHkaVJ1UyBB2HFX5jYg5vYdkikMXHijt4YL4ddAtcxZhJ/mHF8YOnnJurl1sNdyAet9zNr8j/
6Wc+RH/ulR7kB/4tRkU+f74XI8cYv1oYqTxqjlpL80eheO7vEybCUQcxJlvJ0WE84qXt6zokTjoM
rQ3b0r2eP9O/m9sHt/3S1XO9lk0BQ92LoE9SKKmkZwzhUbOzkPpPxzNI0XXPc+ohZ+DHGFaUIHta
5PtKhLVSUUmkR1e1oF/Bvlkg7Rhvwe9lghc+uqnEsqowz3e08VyI3PlSzT/eWulj7V8Ehci744g2
Vd6OshZIbSP6B1TMke5lWRd5AIZrVyR7M6QX+qJiIoKVQQwXinn2C92mnhQPe5wAWRHmDmSBhiUT
kQkokIhtgsSvl35PTc2Be6bmN8VIwbhj4oy8CLMFtglGgqlSR8ywxJlvSuWH4Q66gx4VZfMjDARp
nd9f6BwJth9rqkiYKL5uTJUcLCvrCSdmrZBO8ckWG+g4ISOUko/iL694T3n2sLEI0czjQ/GTZ4WP
7ywQQJRgkLKe5nEudhipcssSMueCped/w1mkifdCHbFZPqCjtbwbi8jHiQJ8khV3iooKCqjIIhjd
/uYF9xP/Gpx1KUew2L8dqhLXNcj/tQAPZZjn5aTRn2AiqTJDaAniRqpwgynfOt7yThRs9JlCcEBn
oLmOqgh+BsbNepLvtgNPsFHJ/5fmSy3CvaFLfmP1Gy8mYvQb97MGPX5bdq9AtgyRynfdERKkOpqX
kyBPlNzJDQroRNFvm9OEzrAPkQiD1QJ/3+4zyRLKH8uiFGkdznYtsR85hdko9+ltvylpmZM6hKnp
XjMr22T/FYm6yVRWu6oh3awzU8zU6PAwl8cW0EPnpQ24jC3IqvsggbvOGhA27CgrH1aEFYs32hH5
fnYmpVA0K2tn7gFyns8g0PJuX90Jk6nmd59umWl24iHaeVic+0Jm4ljpZse7wGR6ytDOxmg3wxbV
2R1TpSkZeuC35eReWmuFjj6znTxhxlDwJ7Le/QWgLGBIrmayggKEKm4k2XDGqUFGcWPYWf/Dpz/N
XG0p+mekLQcfqMphKW1DwBJoY5xviNFDmVpY0tQ/Mjgr3l+t7cqTiJCctoEHc8Bl/a+iDFpbsTHx
q0gpslwbHOvFr+h2TLye8egNM1t+VqG4Kj4aVSGcqUQzkef72Lbw8H2GWMG7MLhtbHr2m4imS6Nf
ZKTlujt69eiBOi9XO8Ev3nw9s52R9tw7dMPp7RQfqfqqt8OPH/5goBjZO7P/calUYzzo8+QSKAMa
ckcE7uuFVAhp6xWLSM4TJ5TVqDHZebAevmywchna4/FmpDTQ5M2Xb+tOl5XxwXU40/o0bKkIvc4T
w3xftASdYR4R8xg9gce1mn2tjDOJ/tBh4Zv2uJe2nweLECzbWlBNORLxiBl6UlhV4BUpXcDSmbaQ
FHLekfgkl8N3B3AHBf38LiXl3r78kK1vVM/ec3TKTAuIoTuQc8rcWUCgiDrNVvTBwKaTem98RHMl
OQS4FTgQzmwIkF1DvqEst5HyR7i/nNbwZSOZXEsbSoCClDy1Il+7Nh8bi4rfJrR2BrOLTO6oeWFb
ivv2iMm+aJZKdOGsluVf0VQFM9Sh4FDTe1P2MSsHLHRcr49z8G3YNoUhr1/gzSrFHpG/Gp+HAYoH
dFrlcw1bPygsiY7AoIcF0K6hJwYCDUFUNzLXW0IODskLdi8q7vv0lF39Fo/kT0eqWod4GrDmhzkU
XEbqjGqM4MK1kHhITLSsApJetNW/o3UuiQUZ87huTdWt0/6zM74H4kIoNnGp6gNFCUF8melQ68j4
LfdNjADbQiEsDylR0d10Poh05O1EsYjTdhoYk9sUYkEt8XBkX6MIEzdnOvbi97v4fl/vkhZZIcjR
K16JYu/STsWzzuH8eUDzm4Ipa/DqniKQlsWgTXO8zCpuKEj3Bn23pZM3gBIPxF30eoKSXuC81hbM
drMSTO/wj2ikCMoiS1mVJs1hAfAKCq2OzuVKvd7djXOHeS7dWaFsiMtmUzcO61oWowH0XvdovCFZ
gkGEK0Y93pPppTlWcBIA4COX/DLn5picknplImOwW3fG9DxioIUCLFiBYVa0mMAoJUOtIr37rbpe
sA+RJNvU7Qqj14J3y8fc9pB9kxZy72Min5zEf0/xA1CTsblSx5CkxPgb4pKw9+d/d22L4DeLNGyW
8QEX6jIUeIXvqyY4aalj0/Parj2ziSyMAowvYtkDWcQfmdJzz3WwSm8jwxONJEtC6hmOd3Q7R3xJ
J/tfqlMVchHiRB3ZA1q5W9ktFVWDB3LwL6mKUQ+wPpIPvxrgOyR1TCLHcAefhrqa+zAkf7x0cnkB
z2/JZIGCmnfTSW7wsAtgahTN4tjyZrlpdUbHRHssBqQ/bzyYr5pACTGzXOoanCMGwrU+8f6DkGOi
ZXZeHiJBJTOVcUKucizzlza4GlCX0bpLp2KeHdG2MlCRIT14H+r/pZX6nYLKjtGI1eQQSFIeYFFm
ydpyKCJbZ2G1aOebBP8ibm8T2y+MGc4bua4rWTw5aqHspIejt0bf2Tpo3wWmyisqP8+XlV7KSSGQ
1TeKWMSPPzBQNSxrpyTvoEqLwU4t+v2Q2/S44yJjA1PnXAvOMCb9lNnVRB5DsyB8oCEknf38uvHw
XYXNuBNFY/clsoxtToKiK6Mn3VuYwgdi9KSwonkNZJXWdA+/JfAmpz6zYDwY5du7YYnqCBdm1dqo
RoX/b7rlG7dTDsI+/Jor+5zY49xe+HtNMxfP7jQFa0Ig6/bD+wYczdaih5K2xa1N+YekNB5cvj42
l9NH+Pquw6YeXOXKNBGW13qPSYeBsPZTxPP07kFvTQi7CNDYshZ/2+ycBeGE7+ZdmBQN6RRc1FBH
qnhGqjkxhJCtAGURCJ3C5gccFMUp0TJWhVgu3go9eLn892XOlqIos++iEAxcYZe15rlSMsJmS5PH
ms2Biuj1lKO7uU8VGPrYsiZgzXZHo6BTcyNBduz6leqQHKQxcA/D6fNNDwf+2R0soZARtJ4WZkvx
NbVhHuza1UnvxzercbLyvViASDB0cLC75kmFsJHzPfMPqFRk6AXzuJpYAQRm0/3VJshwK1RZwNfz
lxTyW664wv9441Ye3/YWKcFPgLtD7GrUU+Up02miAsS/8ZLF4KHKA8BpHh1Ki1ySRN0nanLLsDR6
GchRlXhuxCqBnIoWJYcdu9KJtkCaASXycl3Atc2sz09o48DBWh1i9Ail0ukg+So2NkUTPl2A0McK
/HpDMvvNRfZnomNUMluBGnpkTBZXVVaQ5feziQlrJjCQj9omDZajOcnJpZn7FgYHRIviAi9JRIUE
VrXMZudV49aHyfl9oaWGycDI+hmKMrJON3HPKt/LxPNRkByuObjFSKfQFzPJj/cbkXdmFVdRqlwS
RG4Se/a240myjntfkuy/3zoFUP4NdgY+oC5TCNnVZ6aLuwsm9M1UW74lbgP00IoDfVY/fh40VJ0R
GMY0JPxwkdplPpp3GuX7jOx0zx1JaIgCXP0ob5p99SEeCrmOGauTGd7ZxNd44zfKloGEk/0NcExp
wd0EnwuU8/sqksUiU3QITQ6VKuDCpCuOjIoVsoEOo/oNvimJG9G6gdYXCFI32Prq0z5zPB7UbwON
Y6MIy0jIdLaqwGQncjdw5FElEHrSS4ma+Y3jansfxxa6wCw4wgIWZ/6fofK0EDwh2WnzrpeKblII
BcUYz2o/eC2YvZmEt5NYd+KFheHM0Y081ZXr4gI6SgFgzzYOb5hoQsIEbPdrvqIFaoFEi9+oF2gH
NGg3VC1kzytCvkeiX1Sfdc2x4vu/Pw3Y61d2N5cRkNOTNhyZaNhidPyZP87ZnQ5ZRB1XtUS4OqcW
60I9oNcx9PcCldLOlKaB4YRKcuLGUqe6dzNAIKwaMl4tXWiETYM3hg0INsrHQwBOUGPen+S3jix4
2214mcJWWxiQY9pToyFxXvqRQETrM9rxyAbbpZ0wAF1jH6ZoCFkweKTNAjCAJyrULAIKSnU75jJl
2LNOQbq2k1rPTau37K7ac91h4eWM3OmX9JWb74BqWh2ofy1VWWe9qTMGWZLFB1bTC8tH9XpupMKg
bcAb3cyWFSMMGhzrb8YyTjo1aGD+9euqbGjHyjt5IGh+yRscyJsSep3NvUPGo0Ff13LGMUKzGqgO
/ijZZbFLMG05SVoC22AJRsWllrPilv2rMwYhXbZKmJNInOUR1zz/fr0o35f2HiiplWf/dqqoPXTf
D/yM4uvoryQsoof854bQda+MiYqRjiJR0Qtb16XVPDtO9aj89hWrs/voLlgFVn3aoxsXgkMSHjMS
d5sSbwjll3AhH585G5cTSbViZx30yg8zjyhdBc/8GUbd0S5ZOvMt2K6S24teN71859OM83T3x163
6SplBXVkLog3z9zGQg5lLkIiLAwCPq/1Y64ze3SuLR8yDFqAztGWQ+3jVkF0DB5YgzONgnBXX5Qq
4Qhj6Xyph6WM7VrYk/tNSip5OLjUOg5O6YNSBOcVznSAGXOE/dCp+321TAz+nCw1xtApFPANAQbJ
12asqQfnb9ZnGS2CtmAlBeZvnA5x5gIaDmxrq7lGVcSGwnw+hQIfU0QE89ZFNXX1YJhFuXGdnM/R
KMPujn7F8ARyG7/skVEPM3R6YCnM+iiLiBf07IBaE4fnzhJF3PkRkBr1V+3jzYV4/Hz+zyC/Vxth
Q1d+WJkX4LUhlVrAW3tnS4je+K5HFghZ9BJgH/TcRhtiLFDcaSLxhU1qBz88pT+ArMXyoW2ifZJC
caJaDTe++wcXHW0Fx/9PcrColi6zGrzzZ7H8s/qqVaLIi+2uj8OAIQX5Bk6qqNOTEduFCOfGX1kz
N/L5nFP8IR3+W/zu/BuyjLvSghdZ0I5HSiNhAzUxY9ODDZegBYHeMqBvlMBa32noegXIcEVxMl48
yW/5KVYB+3A1+0IBoCUuOLrHovJIF9vcg4yeLccqqzGWRi/3bHe5K+gkM1aNwTKv3Rzs4HLsX79Z
sMeeBeJxzF75cJc1BwW67H8X+eSiUEvBnbElUhelHgbgx5U9wurQRrJ6S6tpkIPfBZXCA4c9sKa3
VzHWeUr/YDRMEG6Zz+z4mH71VmZ8jDtgkp6roAuvjAixud2sUgqYbTL7Y17zVtheNO7OlGgNgd42
exqrHULQBR/KV44+ofyZeCANvw8EtTgg25dYS2lWNMIZnInNBiR8gBZEbnqw0Njl3PQ0MOob6UCx
+1jQ2qQEIEtXntgW9hKfgLZUnBexQ0ll3p7RHzFfB5UcmNsSrMgaX83aZewcJXbtRQPenX2vPafq
ReLDLL8kZ5kg4qGdfBEVJ57vuPatLG8r5G/8s1B3AwDOPE6VZBk/sy+R/s4EEtOXsda9MktBn2j9
Rl6dMjperk+54AKh8FKY60hlCjL6hFrQywxKP5qecgRIRNhC6XmtDaad749hLxNb9qJXVvmpQWVH
ZE9c7i+eCdmohrhjMbzUGgoWtmJU56reLoE7oKuA/xEKVdMcU+tfC/a5IhMOPsYlZW27M6t74aw5
wxCtdYvOs57UhIDBTbgT+ZJ+OGzBYS3Pj4VcgSSf1OFt6eWi8AnNCDiidhNUeiDdsG+5CljCRykS
v0yI2aX67zQwVFaofxHfdFq66glQSKnR40nfelBnhogJ9ryfkE1uXf8b7HuQodKu5Ptf8MrCYshW
1ZB64ItWcD/zj888ccJQmsRt6B160PqmnoX7CYLWvhcAxR62OM1f3523qhMFJxtjID3zInW81jTe
wl4EEmeJKawE5U4382koNztK24hHBIAG4JfR3iSe9MtCCh58rFMoWS3XGxz7kNdpZprFPQDF2Hsw
eR9PH3mnNsioGidr6ncIqWcVT5K6oGapJpNAWPXv0PQmlcEHH+lnZnNEg/br0xAmAgP3gWe5mLxU
hq/vM1+KZs9KFYFkRPWTCZf/IHHDs6RZDWLZP2pOnhvPOVf+TKabTmY0ZIulpiVwgBkpRuLSmDLV
Y/9ms2hAnIpmxXanzU4wneFpyfwez2dsuPG+nj+9kBr+CkbkFT5dqtufgKvUdxeFnnC+y1e7qjSN
0+nlC3es+YQ7SFlAvJZExatOrq26fu/j/H6Jugx/YikyVK4S+/DkiFNETAs0HxLbc+xSB4mteIoG
hmfoRZvxG01wHipSesW2JwYSe7ittR1GQKmUKFWmB8PM1iakv6/TfLLcFmkRV5gISDDsjp1Dclm+
GC7hg5TUQS/5JsyFy1PV9I9Cc+ae5kXZ0IzAaOCTjDalGJ0SS0GF3Sk47Uw4hu0LMPg0Fx9JsYjM
sKoq96/1YlUGFqRv1QnP0ZBmrT1wYSesM1r1h0FaA1MOtW2duOblrz97mBLj0429OVUSGfd6agWB
xvobdY6djl7Bq8Xm3Jho3HfPkyKK6hXPmI1e8MBqV+T0f/hg5E5nro7h1NL5GR9CTJaA9AvwEEDD
rRan6+AdgvzMsoqxsGG8hVNtR4wb8NqFwPyGcnINmms6D0ZEfe0joq/V431QXHhz9lkyG8KU+lLZ
41boiuF0Q5cX55nuMZAC2aJ4xhJ+yp4Ar2AUKp7uOgDTnZv0A4Q7TBlIZw3aF0dYhp5MGyje9EVc
0yyggyFGHP8wsJUx54J5lk3F6qYqOTQCIbi4oIYalv/JldDUjOueFSDRGElOfHWQjARNRujLb+Tq
FFmwB6ajGLxF3wWbQoDXu/+xKYW8O6r7bV6CqjmOpTR98/FPNECp7AY9bd8lyodRo7GxHjB37goq
maoh9IgVRs1ita7dvujjaAlw56GtP3R8pT4ubjAfy1Vb4l2XyUMZKQpi+F0dmxpi5pREBbtTCdcX
eA7yyolMGOx/5F26ZJDpfud1XtGI2+hGu4KhHPzbCpYLIhR9x/ivjO2+QcB19JYeTg8xSaGweOWA
cMfRUGBAXji+uOPUM44YZbvnFZJzZU9xy9yyzBHCRH/heYhZH2hXP87Zxk7BfPtnY6oeZgGA7f0z
6qkg32lat0TSqpqwKE+xK58icp2Q/8brUiQjbrhJ1fIG26O60oEFkZPFCSAhOY5zUybLaG6FSSnN
VfsWzWlPJnW/0HqIfMzFpB4Q2lLPuoyxKybAs1OJnymm7/BFRk6V8OFuyfmgetzoClHfg3r68Byu
+4SyxAPoN+tuyjvzepsCC/BIcT9Egam2rsJ6IzlTAgozIGflch/jWoapqrbbEHZMEORhiwDI5IP5
veb5OxmBB7O17dZEMSv7Ucx1RwYoGAZOCWedT3Df6IsgngAZebAT10HMnk7hfRcmDBFMsbX+1J+6
VtJtXydJwsTG6Y8wnVnZEeolPXkvOW9wzBP0KyET6sQpGSBj9jz5p/mk6AAQynB72gKIJFW7r2yy
yJa4zCV6lcWGCF94dWOq8KUou00wykojLfdZEXHh6LMW+PO/Wy9DbNc6JJ8HcscrC++kzS3+TQi7
DhFOFreTmqTosU9J+rGC8vXNIzJ0b/5oaea4tzj4mJ2MRft59En8LkkfqyHWrHabDWI0op0cPg1t
xAee/muDGqR8KNjUFpa/Y0sY8Kqocg7IJKcMbXza1Ha0ZeMKMrep6W7UGIizf0lpsEL2w1A2KPNJ
/QHodod7iXY5z0AI5vmJeo75ZruJLVkPVo0gc7JCidC3k/Ayu+6OzJ+L4DMvg5EIOsoKhrE2Mo86
ifi1Y4P93X4JfbWFnEtOLYCt2XLg1h85Wrh2raDmjmZNUzmM4HXC66ZIBaXClIlvKPZM/Lq3EteC
MKmTBpEd8FLpB5RiS1dzzikTl/xgR5kT9Bt/Ng3WbUWrjyYWCfcZ9+kP+8PuRK5seOYyiyQItfIr
/7X/7QFEZcZfMMalKuwvMFPMSf/YIbtzwSiJdUQWUAkLsOVybkiZH+e817f9l2P4s+cIoDjhYhq+
K70pAeVgnAoaYEXNZMeaLQ5MnHU1WQMjE8H2FSMXrl/xj1xUMfImaI4FZzOH/LFgTtt23Q8lwWdB
FtmcM6w8IuCBe3/Xijd5Fol6prSHcFeKH1VI75V/J4X/AqiKf+m/rOm8I6A/EjzUye9oP0R4rCmu
ttFVhjBg2z6198psvMPd96z0/cFImV/zEYMPOzToL7ZUKQbFbZ1cYofzRVRgAisAaB4dU0dQ3u7t
fwH20XJ6zzu16ISGTqbLCw8/pnpdfe1U9ixk3pZ82a5R51YUOH/48e1ThYsbr9b1RSdDjdB1NCVI
bcHJ0dsmyquQQFkiJ/iGr1ny1/VH0lw+qdZnQLT5xUgqQ+UDKIevOONSK32ifLyi1iaWp+6insv3
tcXbjCGMr77/+CXK4mUe3X9jQDSv1VHhizZ+CfGnWpywPW6X7Vmr4EYd7d12cxz4fpv4fWsrPlNW
JkYMyV/dPdkOdP3Gv+Odz9OGw6qoUgOq2+tO/xJf6qKmYf1+DIlgIot6QqvlxSPUTAwLKTR/hx7C
HQSMdKpMUqAGXY492tNvjUFF7aPbdCWUWQ74e6b6DE42fPe4mLULm9yu37obtae/VXaI0/nDDXlO
k6353VwYn+6cdGQun6cQGMeDbIrZHwShM34k8SUmSEA3VCRiopixIsCX7enA43qr//7Dn+p85Ve2
kg1sguKXN2ryF4vBrd+6AGTpvc4jLOCpny0Xa1JWQkkb2zp4n9I4kFQNtgnaYrfvdtyfmiT8secO
NU1R4E2ahckXSL1E2XzEyrs9vXCzxkLkTk2/kxEirbQztbm450FtJHjlLe2PPX+7nNvhdtFGMkr5
SukhSd74nlaqBWmJYSGVmiMJHUK90Gm1uC7EVrjtMvmFODb80cvt7r9XJCvBNxw1lFkC13IlqNMg
FKxnWVoT/9besVLxFzhNdaqHNNSOT75r9x83U7mU4PCbBBXW+JCey+0ziC14ZecygqoM2YD4JQ0A
TUf88vbT1Xwfg4I9uo3TVYnGwNgUvoWnTNhYIwT6hALti3QmOvvZY5x38U//cOpy5jvi5HYLJs7X
IKCmVQXTRw0VYtF30v+jLkIgDyu8pSPaUICIQRJwjkTxj4AEsELbzR4RqJ7lDGoHprL8AxYOlWS/
DI/47wJAyN9M0AYiuxaky8Bc9+mCtTOv4/fJdrAAqnZPYTsShSzxrCytOUlBF218V9FbIjtm9e+O
+ETmbzzpJ72M/DQed/n+3wrQXWCeByiQADHvEJSWkuoBA8QnNHS5b0hUen9UIWEnHFnl7tqKUx/g
wIcbLXGN6BKHkQy/UDjXAuRdLdxMu4Bx+V0miTZeCAXyUR1RqYNE/zolyxTCwaYEcF1bhjv1x4QW
lLYFRN+ZN4D9B6i79483YwwDGLlAGlJmqSxOP9jaPuyxZU3aunpcvZk9f81oK/BQnEl78n8WmXOr
f7b+jISWsifQJIOStc+6RG0SY23ikSnc75xbzKpuhql0hwqt34REKA2qLNDBnz1/jV5IYlcKCGU0
BI1FOpvXcFD73qX36homa9Dhm6C06agGACqxepAd0x9+B7OTFt5xP/JaaKIF1L4Fn4uzC8Xah2kS
p2jkqKkgY93iRZ1EVxul7nyp2ixaM1joThylZGaIxXYuw+X3dyenUa4VrMvqyW3YFhxoo6dQHOSm
di70abipejI75A2EnO2b/WoamFzeAUSpaDIpmgaGBtGS6skhzUfYOfb4v7ovSLsVsMof3NKlwljL
4RoVBgH2R4OMOShJ604wAm3VGEvCQ0PRDzEFQEo6bOVjFknkOxflbzdg/Cs1wRPtvrDiuqiOrb+t
QdEy+o9KmjxTsm7ZK7ScPtrUAvQjtcTstqbn7RGf2UGH84oTd3CzWQuX5DVRR9D4pCXMitJLzOWF
1ycan4nF4fur50DEVMSangYd//H5mtZojSHB/CjWVZFQUG0gRr6ikdcIHfkO3P1Q0mT/uzhZFIeu
I0fvDveghKDoqUR78X4b8bkvLlhN9mGOs5DVYvSE/RztTLzxJcMZokQ7UHDLU52+svOLxW5QuhxY
oCwPLTcLPOQMrr+e5/g5jD7CqVM18QxOuea/oF4sUEukcsrGPm+qsHmxSj9myGKpZ4YmzAcNKi/o
/x8+Jg+ZqT9tvVNQz2WdGk6Xxns0+i7SOT0OCPnB2BT+F7pzxR0aQHn3Sz32NuTfvROGch/iFYOm
eRIzoeaR0EYeIQuDDQ/luhsbMF7XQ4+uaarFaduV8j5tfJCaXwcVin/KjeRwHC+aw2N35NFjlGoz
+6s6XlaJSwnZ069kPMQR3j9t34OqYYqggBevEGwaH/DSl1TaP3iw59N/PvUaoVrX58b+soFWlCQj
Aw5xvSnbbGDEL9r/lb3mWchEsLekIqnid06k6HyxlqtmhW96xwQp/ly7oSZUdWmmMo/DSzTR0OM+
wHVMwoXhDSCDCZLGjnnof+tRR/atPqIGrOFYtTqL0IAdKcXcIpPC0dL6qnqBRlizxj6NRoGQlTi8
qNmBozVWJZNIenuy02nmudLeoYzr981b14RS8L/H/THoqTmwyuyr9vTwNhnOh0U1t0OEUQf2PA80
ZFzSQXN06VAB9flBX9UYzbAq06+bRR+RxN9iKNUL3Sjtu3yo38LPS0ZlCyNHq3xxwNpmXL0ySYPS
iJOAjGDax7UbZXBf8ab7qhLWP9LwwXoJrrlN3JnVUm8PiZ3r52Xw80Y5KFUxVajT5bq7pUpvNzjP
cnBVlVm8idYJLRjY4GPIt8dOx6ZrXQrnL9QVKKNN1z8uGbiS8+7rQlCB1AtFAPFhKejtTDoHyRSP
bELOU/UFhS52xfP8prq58zBifQrG4rvZyU3HdL3R1oQQ8X+l4yBSV1yE1wEqK41/1Bdd6Y6TFI05
Trop3Z7fZelrgCu/E+eR2cvVNdGlSwhIYYVbrhfronVdHtesL1I9nKXGTcU2QybIYiAJsGJFxR3d
WqVcE2wcfoTzPkPCJy0vX2a47wTZZzLjh2Y6QjAb/XwuzSdjm+1shHEMh1T7tRSZxMGyQi5PTAxP
e1d1QXTTbGg2sOPGUVpuQYcHYTL8/LJjU0apkN/km+KfndEhXdzaFehPnorEtOJMMzyIa0VuMQKp
ZX0alrI//4x0pcN7e25HkSm34w+PyRLqJ/CnBWirYIh2bDKiEC7xaqZY8C8Jtyw8GzI4pJU6Yixv
eYcynvYynJLnHRRbTkNXc/Az9xNt+1DvAoKbt1hNKcBOZQm4stz5IZ+v+tnUG6fDFparnkRwHqai
41+olxp1K6KEoUNocg7lgC5E1YBfjJ8ZTEkwXOWfO/4KZo/np0Pu/qasToKU3ZFDrWmnTK0kNCBB
7zAsSYjLfzKictvRLu1yWooLvSJZzLIG2PP85MFi3MEN0y6uEKgD8xDrcq5j1ruB2wpyX8L8Hsv2
DPxeJJn/nJ8A0pJ4albeD+dD4+xmXwAP++2CeFV4v53kXv00NrBuT9q1QJuLOT3AAKciHtCvTQrj
JpGPLW2XcweXsnAW/dxclFQzUcUis1L/Fj07s4p3q1Eew8tuCtMmnW4Rjh4OODTlyikFuOUp/tmU
nRMc+n3o89DsK3N4QjxWzBGN2eiGHjqJqejgmb4AOUEcIWXtMy+scR6hHffR6PL79K+KQktLfESt
KoYJetD+Hz7Ljw5H7HHUg89c+t7zaYZHUDdHifCUwaYxad5gfH8a9RWLW0anFkAMSl6JMKYkt1+K
frdPBO5L8NbGAEBneuK1joHYb66NQ/OWd4Qcc2llgpnUS9UgvEz/3nEz7HM0yDqrKtICl1OHca3S
g7v+76pmLMKshwgCx3hAU4RtdoEssXXqQaBc44e8v0x68d7dkCA8/kJf8Epqme8q7tr9EzirxIUT
HkBaRBHV0JajSIfAwtzYbnEkNbi945Bh7TjiA0afl56OJPYtyT+CmgMZSH2p+03zmCC4tymxdE8g
aFNULYtEz62YK5MjvRei7W0VpYNLZdWosFySR7BvoMYrwnsAJT9REMa21fMhoIJko4ws7iLNh4Hz
ZECytWZ1Dnkg3n1t05GIbPZcfFHlH9ArCDvq8qU7yh/wU5PSd8c8LLkBojbfqAx96Urb6zAUvWZh
fi2CLQ4qzPwdlxeSxc8UgAjck6+jlLqaZFJmrt/6iV+ZFEys1ET+ckL7pyk6L7F6gc59w4C01ffY
SnzSMQZ0TNtJoJi9XQhN0qGVkkH41MjrypG4X2KRPefX1O/mdkChDJSVq/qG5eZE/R+LByvunaO+
GdGcekPw45odESTJPV/pVIznXKd8f4s9QKmZ4c2ag8b6TvM2LaG49NWs65rQG3FQQj8Imwobsl2c
BRP9MkycbTRawix9766rkN8Q96ijA1lN7evu/vpvdTW/rh+CcQcOvFjMmVL7TQ9wv50srPpIopx6
JwaqbVaicegJEjoPkEe4AgEbysfowXk5XWQrRnR90Yg+8Nqu72l+AGxjSkBiDQFPI9KlkSoL3vk8
O0QPn3Uf0uAuVx5c8tj5tUiCWYQ6OyjmdTxcIAtpFswsHToxUOwXqcZuPPkhUKQZvsrJXWaNpZkb
7Jkad/MgBZYfYAQlIowBsu9hcbPvjbhOYH4SD4lCbDHPAPw9D73lxa43Ytld658gY9TNZr6sFvrF
o4xV2pnjE08AfRs9Bo0SN29NqYOr1zu9psjdoykuHZdqFDkf13j7910shvNylQMwfBIjTTp3QeKm
NLuBZnj3enhaFkrffKHQFa+9bsoYl7e4gipzqXnZvfsigvqUy1cxzdIdA6EzxPfplUCq04t2bsZn
7pzPzol9g95PgnX0CVujzlZ7qbkgyHJ4zzTH9WFV966DG5McDkp5qRu5sPqkKsPd9qFq+eOw8oKf
FTZHOdEuIRhF86Guq0wLIFMbkdVehchr3j2a30pE806qWEXcV23AajV96ASZNv4+CDTxZYWSlCNT
yT3PykSAFl2PRnzD6LTt17Y7MNnm7gj7Oopfc3hAkxK2umLg+yN0j3R/q/NwHS8eoMETm791Us3b
SuDkPxLIuS2U4U9e7530ABXsEhdvZY6Z2aQw0SfuhM/6HU9THFwwf2q2ECBCr0pSbbnt4vbd3waJ
1zFKVBPLn9vQMnlNbhEffPgmx3akh8+YRg2ghT5bKzz8qGnu2BxMpmPLclvm58luTvt929lbXC49
kd8oKSJh7PpJStN9c19jQh4FXhMBaNrKMdn3wFW6BrnWzakvOPKpuLrBkqVrnPrSP4iKBYj3KQlG
OXUj4iOudLuwUwoAvgQJdzPrNbIpV3RL6bZiriuaFuF0cebUFJ3NGM5LGmsjrtrqL4OLAArPnlei
CI13ydbHq0fw2i6wBDyeIcCVFn08zSxnlokAEHYdDOgDb2Godj/6XosQxYhOM8nePcKmv6qARsuL
9GJUyYxHXbIQQ2B9rTG1+VW9MhKPYiQxd+W07H4xRIDIRrNJ0Mag0hnWwX3+4Q3qIC8mQ7gLSK9W
m4KUFvwJkpkTf+gW92YKbtqs4WvRFsUq/KtvEVzJkxofn5frMIBVU96+OC7H8mrUffyol2wA+bfu
31mS1Sp8VDBo4NxEVcPWxPi/dVzvBnpWkpXutzQTjbdU/RCB1afLpJtXBstTsktUA6NFpoHxzE4I
KJqMKZObtJhlTcyFAUteo6Oxih6qrXwZBbr5q7ZdYQ/nmXzsyxJYnOtP0rguNqN7P+/RKiC3QPyP
qcuZ0xHLlzT+bGkbzGTGzU5WrQxO0dbhiCtYcdkHAliEqBRC21MitYrdUfbhjerN2TJ/1vvqqlS3
ORA4WxTow2dbcePu7v5r62mv4awJJOHoE9Vr9kwLG61GgtuTvIBSjq2PFEX71YUvZQiBeQrY9npW
/AVSrUBtqMV3oR0kqPOUpf1boJMrIWFwecfrLqcrIfqr/jD7HAWQZJc12qWZGb9iCm8/iNs/Du5n
vuBL4TuV5wKqo8eJ1Vl99ElAMG0VHKftnFDY01p5gJyw/23Kvo6EHo6xf/1yamf4xlF9tXsVNJ7C
d2KFwDn0XsxQdqU6mMlm9T1LFrTZ4sWbzLbFLFZ1LuiXIxxmtSTdDegH8G/0hWKuouHyOrwzWwUC
0xNnQvhIEZ1yaXGICNHKpLAEkNS1ZnSNCl6+N174nSbb94Mu6fKzh6ZlSQbzzNDil73hsAcBJaog
Nyq3rBp+5igceZjfn0Tc60h/V9SI7S6dkKGLRg3P3/Rik/7gbZBTyJY5Bvl32e+bch4q5SRRuMk4
1DQBSwPnDSUp5LtX8Cv1j8cS8TRFyrJPGm4mxMb3hFnLgDEKu1Hx71qQiAITx/Xs1oHw+1YhtdSb
ShuSEt5kmtJSvPpSiI/WYEcXX7G3GR8E8P0/rYRkbdXeUVaHrigkQUIyFeyoqLc3HajOI2FZ8dMf
IXhzJGglDZaqb2FtUDlbTsjKScC6z7Sq6m5j91CX5fxQT4or3uLeEJycU9Xrjk0jI0iebeKxqYdd
l45JaJCjsGKprSZ8sn7mWmSvRqXr3J+qPxWvLVNxkCiwclCZzuJDpzXL10LkrQagT0NrcywYDUY+
oZkG3iMrMiok3QA3BaOSHPn+PK6b9qXtbPI3W/blwXFG51IcXhjzHfP/K5KrCQgoLsuKPotHcZ0M
6mi1MfQIYFVz3gEV7PgIYhKpW34db0TUUWFaremDISowvZYpKKiQqdAh3V58UrWlcSValLQLY+O6
5UJ1MaPhlkAkEDQktcko8hifyd1PHBueYZ8Ulzz6QLF9jRLqW9LeYwM6FenkDbIC3TFc7FHm/SR4
ChLvCKKb+4TD7e3fXHAn6ljQu4mp1b7wXc+VICtd8ZEnm1CtwviZIWGtVw1D02UnL7n5xLhqCSL2
tER9c66m/n3Zhx1Ffk8MF/hg1Qw5bl7aT/MxN99JTV59+YMyY6PWgxpDafYDVdz+HOCiZf7yhmZ4
zHjM7L/DTlO94030MKsfnVh4VxyY7FJvJ2F3KlD5A8eW+t783fk3tcclMXokdW12DGnPmoubtIx7
kiD20TSdDbXXmsUjcFwRPbYDvC2RHuh+QNSATubpn8V0tGzYtHDsfpNNqOqwWg9K5NQN9hH65mG1
1GfPsM6AOVvdzl6FpoU5C0PL/C39tZuDtje1fCQIDstt5wvbuSm+mTxyDwhp9EgJixhnJU9GL6tr
GgiveKHxgaiXqkHir1UswiLG/EoI4lOD9tRcaue9Yj0i2bYY0A49ToG2YQnTOZNUxUEhwfpAYZZD
MVcikFKXttoukqfAotgfObM0cp+moDNeQfvIDaJlp616FRuI9Hu12X1i2MnZCE7zujN9lagtcQdj
kmNOqMBbKHt6kKlyegbvt5ggtD8xHgTqmmo0LXRE5lAoxRI5QB5ye1pHTeyPl9aqCv+0nab0lNDb
uQbvmsAY8TBwbhX0vEe3gRCq0ZME1NXqOZDnQTRKCtif1UdtFPzRT0GB/tuHXQiHaSa8zdyPIXHp
ToWkxuusKuYd3zzuG7frLFuFO+fd27rpn3Q6dZtW/DfVRp5eupjzMYCQYHmev0IsUBily82HCGpy
SEHHK5TdtWcLl5HZEvTPqAIY2eH+xxsxiqXf81kaVmAZEednU/wFd94GQLICMYUYiNPzAzr1+1O9
xHIEwPDVvkKjauFhWKoBWpe3Vy91urab8h3kAD+zAi0Y9BdElje+DobTOpnMOtyEE+/wvM15Do3N
5Slyqrlmx3Czvc0FcWkgmLj0z076GWZZ6Jt3zPOrVyGyNN6yfT0B7p2o/Ga1YGvoBvqbJ0PFeZ0m
6HBLJpL3VCK1c1ib5OhQeOWcyQrE4mLnbG7pAVAPPBifTNWf2JzIlvxPH6Ni49tJeUUVpX5nogM6
11SK/6NLcekKFEuViqRxF9v70wDtaJshNGE5yMWbacr1rapdUw0cvYuF1HpsRS/7PnT9k6i2FELr
bbE+XojxyR56nzWzojy+EorTmB8ntGPRIU7G3yVFekwHO0e7/VyIjcg9mMMB5shF8EZwYDfTB7y9
4ktuHAKQzLmh4gj5Gdil8zINMG/iwAHCuiIeV6s0j3+ZpzWxnSFO7rjj/Ar7RiWqxLkm/HjJsc3s
Kfp6g2+nJyp/Ry403PlayyAB+wg6BS0KYWfoFm1LrjjdCpqWZO/lFXOZCNXzfxfPxvWyCYzeYMZx
SWY90Gu56qp0Rpl5P6ik+l3wEWaImJ64tbNj8LqSNwhPCs6f0w0GLSIAFynvbVuvt91V8ytJJuK+
ZVNvGxk7582eJ1csqSg8zHgNdvqQQMYehMhzTEZLwyX/ZAiUlLZabcowJtKvCBp7RwAXy5Yjfcd2
xyg7W1yV/eVGPATP/vJXrDDtZxP7utlGhPue6aD2o2RhOZ/+69wZjYNJcXME6yFQWuqPGcm+0/o6
Kd6UNOEK0+S+2dWSmLwtOSZljq28hx0d51zEjDGknI97E+1ywhoxxRN+lIxPPFzQYTS4jgMiyGkt
uJVeWlZn6OQJSHj0ZukdQSlbWtP85Nm/IsdNdwgBzSgtBBq2hgUKsbbniKgc+m+/49g/2TRZqYoX
VVhTJEFi424BYWAwlA/LWQFVMWflYY+nDcM5K4WQngofcb1vd9wtSwZyuk3/wiwiiPfXUyL+9eco
zZwv2+XtEL+SJBCLKCbnGzZXtgFn1t1IK8nftGQETqf60kYf8HVXe70glXhCzRH8KSgqTAmg3njC
RnL6vE6nek1Ut4fIkUluRWWmWwfI6fL1KokTXtpy7XqywV10pNlju6PSbSsLrTpsdHUfNybZB7i/
EC66UtZK7NAFR53LdXJV+yLWKG9yDyjT6NB/2e1aC/MCqThyp2H4nbqugvWoKNtb/stiZJzM0VCd
VO25NJfGXWQ+MMYkIioWtIihpLmCJG261Qob1LAepzle03YcWkfxbzmNA8tiNAdolP4LZLMieveS
LByfJAjnOt+PMiIAx6DPbhYL6T+4jv/x4E44h0JrLsFoTymmiWHequkSV3fsoaTSUT4rftXx4Z3q
SJIgkLnF+I1sMgYtARYFzhoYPFPWBAOsVD18nSy7zPa1Ug/nJyWdhBhIwwmEIknE7Bobfsb/qxhS
QfRuTBT2g0YZY6MI6kqcTo0ICw95t4qklWPK+81GDyzhdg/DOIMHc0uKvjQoPrsB111WzJC2qjuJ
iRxgJ4tfEw1lKUTqUdRcBPBc5HEzFXI5lvzhKrk27PDIh7DaE583CftYQ4cKGAPOAYHb8kjQyXVy
TV4vPKQF7tBCetOYUye2RfZcmvv26f+RuSLh4CAInRF81HvCkr4hAsHhw31KTM7MwW9gUaTd0frA
52FXPqoBDcpWRodqdpaDx2BvgacPOoc0Uoi/uo0h6DJM8b/UmzFYTKpRitzaRDy+YGJRHVJp72Hc
xgNSwFUr1wjfEomK+XyOB19MMeDEm0zJJtK1TjT63EWUScgz7JJ/hq+ACqNzt1SkOrq7HqlZvHPq
YyMsehAKrgeCcLprDKiG9zUJD7WVoNRjaxxVPQKpWzc1Km2x4ahkB4lTn0IrFoJSi0zsJkhAioYm
RYSgezTre2jBkcK04zxTvmfvaVEy9WkNMB9FkqohNfJNv6aYynio5Th8MB3wHbDFD6eJvDHNyZUT
2omNteXkeqNwPGX30XeihfYKXAWAAQkHClaE9YRvnm2tE/jJgTKP2CN9OX2swhOtzlKSmS4BfeDT
7dX/y5KhQTmpmH1qLnUe/7A2B69Cc2z3c8QiVfV9XMylC5Lja4tfmG6VTpB4tG1ad3MMVE2q/A9Z
wXXx+7VVg/AORz/XdLlGEImo0crRHPzTACbZW2vE+IDqBxS/u3SQ/N4ZGKEBK/mVvFT2EED3viKN
tnSnThOlVcI3ghZmqPFrnKtuWWy6zD7PWxcxDDR3p1ZzXp3Uhhv8xvweaUgHTFGWmTve7oExbIIT
UujevUJqKydg1RR1RCO6v2UEPINuVlIXAR3UdlS9YghAhH7X7wkVZ+UsSOF7QN9+4hXlo7wGuJS2
SU8U3qFYJB58srVQIzhr/O0lh6/0sW5Pqq1J9EVgk9rosQUHWpb8J4+ooGLX29fK+UhqIeYU9RFY
DAGEL5yr5eJOOBgFJnDYUNv3jb4bLhpxKedRF5+6nmBQbh8R92bEUnTAI0r+t0KULqXX+5txeNzE
TuNltWmzkHvCS8B5aUMvtEly7qmlrAuOAkxl9ywmsCn43tQl6MsIGG3LzSlsQ4HIKkXwgijuTfTo
783q/AwBu7+eTRbnZe8F+DFVxFiF64emvWdz8JuBGgdTPdo2W7Nf6fYiXXGiK9Lw/5hq1gJ9cQDd
b7oKIUesNYQPE1u/3lZGPukqL4fSnyzI0PUDkezwrjg+6MHIdLDlVDNhQVx2rBwWAME1m+pP5Er4
poy+r5vo8N31Dui7ouqUlmE0cC9QctVSYHT+6NwszPTCQHpUCIzkdQZ66J/R885+Xs4Wj6o7Zes3
fV3fYcxBZmEpIIRuqoGDHf6/S+E2iprLwEmCPjoAaK4Uq+WnNcKBVpAgZsSci1dX0Js9ZvGGm8YH
wM2dzcmWehnjdWx4jjGQrjDvoPRR6A5wLPeICU6vGs77wQ7HKi0GkoWymwVF+nxVGnWfkrHz5kZD
W9apVZz1U3cAy09E6Vtazdvy2YQHZEpyzIDmGuHbr/a7hN0GgvHX/w1NfqbX2FTbPsWk6A2oPRQn
XYGAyjfFPyuMP1NXSuycmHMAAyaBtS/f4d42hlyeI2fIOzIeMTuIOLsy98GzaOxLF+wSR2BWTBaS
HCCRIByIZ+pVtAKSkOrgw916/MQVwpESsOG9QH6Gupt7MY1tmWp3+YEw611sgvo70LFn3QR3PRpW
r3ulztU5JDc87PQUDBtulRn8NDoVN3WYMTZZEvFf54rJyNJswGL8g+NGVvhDE4SwJp8G61OSWsoJ
lf56IJmwKFok+Zfw/u3+qclyhM/9lVZL7zn7UdvKMpCW7GaUHsEG/2KIDRj9+hn6/JqjTi1tVLt4
LrxNRSx3OS/WGFKzX+t/hTHf1OSLYwu/KUywnOH1PILZLds2vc+SOd7bNqEM/ABW5S6AlFjkI926
mo6FrfoWYmBoKLqrektZqowRPxU3trh4nKGlT8moTxGY2tKxgO+h1lv2CW6UjJ0lwNJock1Pbkda
IyEViv6b04O/PxfNVaiIOddNPeT5S8TqTB0HDaLcMx6oIEmb1tRJcebgK7YiDsgYIvjx1zvFnP67
ESHx9M1Vzv8kCq/hxbzUUp93Pg6OMbZhxP5kdB171UKiDRleFd7sJfZqIJkggMiXpODXuaTZfWaD
RLG700cVIIcIfuU2kip6ngX9Mq++wiFwATM368Qw9zW1YiZv2c6dWIn6qABu8aA/eQkAVEBn0Zp0
vIPJw3RjH6A6ZWcrCWkt6osqTpZlzC2QkA1p+pUP/LLTMVWxARhketel3wj5gzd4HsxpJdQ5/cdL
y75IXpcOBDibnVn+wTzzMtR3zwkXvN7lFagDbr1rghmmlGxZeOYJjNz4UwMV6K/Tjt1IFxQ70xrm
JVGxWUgD1nx8j7bYxhfE1OK1lsBuLHyHxjdqKIyy0xmUY2JvGRWniZE4fbXisSiWN77yMOQla4Qr
J5GRPm55wkzZz4d+awGuYuyoesnEe7tHojEIflQLdfsE5ljWV6PPkso2layOhKHMmQOYnpCzbz9/
CVEs4CbvWeSRyXaF68vOTS6QW0H8+Hpdfs2nBjUmJdeIfolPnzbdzapPGic/gPDV6unwIbW8U7IF
mAeticOOfjcMty6IsXEf2ITpyWcjc44T/kYPziXHZwZefoCe8cknBubm8HRC5ONo9D4IOVZmg+ck
pp3RQm/KUVfZDq8SLZEXrSXyLF1GrkkHfBpGWp6bkqwsUvX4vRNKVMlJm+c5yhe9j7jXK8kxHyOw
CFnP4TPoMtDS8Y4IB1qrfzVizd/IERiGLckE9eGPYNCEpr86X7wzs1ciUIMgWgAsHAvLK3ggMxZ3
k8ZM2k8djsLWvDUSaSCFXKE5N7Z87+/YnZQrLag/lB7/ax+ut43GhxeRJwEJEsu9LD0mGnvMnrKy
FiHtjoX/s7v9oodjepSLgW63URmlOl8EKMzi4lypBt04MpTdtI+zYZ6SrEi6nRMTEOyZgVrzqd/M
tE3+Bb69l2Jad33VLJZdw78cMfSdEyLE2JQsLFgKlHXBOSYMK8Y1wdYQ76CQbxX4ripuRGrCT5tY
mJisaDfcQygZj661y94JAc+wAyC3Novn8z57qu4wXXWWZ6bQy4SZ1G6bUhD2C25C0he48Ppv0BQH
m4qkI7LOxvGLmFYFso2u68Ag5AuOt8YNMZ7/+nwdZPjZIjRS5kH6O9MazwV+Yue83bMwePujp+06
8Xh7fs8zQKKPsKdw8b0/1Sbil0ExKhSZh3RItlQKSb1AEd5Y81SdETdatJJ+9rIjSOKFxzqe3leH
Wk/p2s8uftmuvCyw/xlcNoGKFhFf2DQaLPwwNYSxmaJTloIwwLhO8oY9b/8M7hsLi3RcgSeCE/Wk
dSwda6ddNt4cMLR2cok3lJzS91umzTWpQqhLIj6854QIyfjI9aYEXMAAAWpBZc+kALna1X3VWWcQ
rQQBmhxzaqESgDTjEKJqHhxeW5TKOQSCzqNYlFS9Mknztt0O+zDG4CCnxv0Bub2QkZ3hKxyzRlZp
h3CKMnub9Zu8AN/KRvt6fnW1iocGnvxtUYbf9aOonhv18mg6NXW/VXiWseYWp88B63S68+i1ajmw
ylZ+7iofcw3GN5Fa30OHT/S4h7wEz2s1z/UF95TUnhajIeSyGGS1YgaYy3u5PBIgM34RuFAsW0fS
50QED5R1JvBsDRApfEE3/rIvCp/v50LPpbuvb90IDzHmSfMABK3ncoUZ/ESGoHz9ecEU/ybLEBPu
IpoXBfWOHu+9BU+eMt6IWPfFyTohbEfGWc11q5ILmCakvS19Yp5bKbaag63E8O+PhlQ3EohcPfvJ
hmnwXsh2oIkXddfOL1lKCqG+f65M/u1iLpNfRWjxfph1Qvi64xiq/shPVqWTtOGCVB7ovw5FZ4oa
5OlFmu1a50OPeqBa0C09H6a4n0LBHC3BGRRE8TZY4XxCOHFwpCBz6eqnXILBroeHCixnSS/AKWCV
vDFdlMrgcS92z6zIV/dXehRdmmst23OrgNfhw+SIaYi3Ts2m7FewZs0oLa3MAniuajkCme83Bvsq
zVMmeNCEmwYFN19c9r6iv2nlTc3vQh16CrTljlwCOcHXm676WrGFNzmP0qJS5IvAl99oSTxg4Uyi
7RSnA0jD7rBXRBLRQdnGCkLAYk3HyW7wCsCn2IOft6t61sw29zba82dP8NRIGMxCW+NA8uNl1Rg6
K5y3UcImoUrsSZRHd88EzgKmoB5sPJ1fYXkVjaRYFObtbY6+lkQu9kZqF0jGGwBce+7AIk7wBpmD
RSHskVeFKbDbeUEmMT+S3oBqZTNpwS7elrgvfml02TlR7FB9OjomIY5rr/WvVkXe/+RCg8OzB4SC
cmghs4jS62f5nBnVhpjP0OntDrnH4R+6CHmNn3ZCKxbDrOS8JkGbSd9LcH86OW2UE0Ckt1AFU3Z2
A8BwjWf+QgY5MtM5voGg5DnLx/NESiaewIW/SI4V8v5lKl9RgZgRYy3OOGwtwRjrPgrEGRkzpJGe
LMK5rGY2KB0yITO1FSTTjCEIEfPimQco733s6aBtaaszUSrJOaiITRdYCXzBfITrs2gAcRkBOxyU
JFBON6FgBSDdqAtP2og7BUytV3YXEW2ICrYdh744yHx5ueq763tCEXhG0hUIsjHdEoAZCu+T3eRZ
rrgUyPxkUpTNVkXNEMJ2laHvhQuq3kaIwVMOq0DGnqsZIPLElwRiIYItsROVgt4xTP40FqHseRQR
4wjDCKKfV4XvUBFXgbwlfP7pmpvHRbqgMomsKpZtujuuHMZMZrm6g/XpXrGwtuqHTe2fe+YRnTEZ
gf38fA0hHalbobeDTR9voyudjPJPJDz7e/FxW/jzlGYvsv1kMGuFbKi2nbiIzIknXDHt++xZgto4
8MtPjHMwAP5jn7Wr+CzFWZluIKiyGpWeuG7bwG3mF6S6Ul7H4xo/wfNv+/55q8fy7+NfT9j8mzba
Shd7haQNYb41dRrq/Sxa6TJ3myPMCjH7Lec04gS9diTmkk7s5k5IZrh8LV/Cd8yBQSoIYgOl0fAx
goF5fXfu1fm8WGsBgN9BR14jnCpHJ4HYsVmNs9codfECSx1vuKGeBB49y30lAPJovHSVZXgOTtB8
pMzGmMYpwhFC1rdep2q0bDm3tosA8sqIf4MsMRZ4cC737+bDZMBPMeit0g41BJFZ0u65Z6omfXRt
qg4DivcPEaYiChh2UlZ+raMs85iNL/z+LUNppJSfRRwd7Y66LWjh6oaCuAIFuL5RyO/wDfE/f/ne
bzErBYKoRCYwLXRwxW5SA+tKkcOmZsqERAiuqwIiqPO80bTqnwGmfV2XXIzcXCeTqcpXmH08Fyvu
vngB87QCVPRsyAzS81DbUCf079kUy+MR8wwZ56E2AKfV6Bzo9+r8B8+BrMj4JYLPh9Wwi9CX5cD3
/GkmOPLnY1L4YwdSDrx6TjtiFaPSAhBMBeSKXNNex4SThehXOJOBb1Y5EBsDwDSLcEmCmtXbG24S
eIGXUI4LIFyR0US1ced3uGApwNxHtpLnOdjN4tuIB/hyE7doUmycKAK7EKZuXSMnnSyYKoSqWHZG
ZtaOucQBIeBIf1XL+gy/KIiKQrvLsdlXUHCsT2rI6HSBTJpVXNX/24ojtD5CTfoAsEZnmyH5Kg4z
GJ97cQJnhuBRN1+KDhaO/Qn+YI1JTGfJK4yEMNt8Ht4xEa+VZNZQjCdBbgsEbeFNqsvRzEbPKl/j
gh2yxmvG1ycEvBEwPtu3OfTs153geLiyCwUfLogIakJV4GsNHDfeMIDbEzMxSsnsc6D2EC5ayI/r
/W9uJcGEVRLXl6GiiZe9GbuykeI5GlOSjDgcXhGb7R3aZgl5rZP6p02KGbEMEP4MvZuiObevQ9kl
DQMTlj9HpLPuoQdmEV7BGtpuIn0Z17PsaxXjOv8Lqul2vImP3v7lae/yRpzrm+ya9x7pz2Cr9pF2
45ntF0HQ4sUzpxjvuE33bpDNcfBiPZYLDbX2RaChHLCzh2cYQ9EUgBOwvMVhJTIKa5o0LlUtFEfQ
OhJqX3IT5toyk9sHPUE6I58bqX8/XfIvYVkldpBU1POSjSvDcyBzqbs4zh2pE0uf1oxwBctnwHkS
3OuJyPhNORAP9MlgCv4GP0LPFxj2brK4/FRLtVVloaI7YHhUPqA67NzdRKxPJ1/tsgyCMJEk73Hn
K5hbS5l9Z1hA1H+XtpxVL8+LSrgxlPbt4siO05ghDLC0NELHMn4Y7mka1A0RB/ENKDiRmto2q8kM
ci5bnux25a5WyD7VwikR5/3B+xOj8PLkWJvD5buVBT12eoTOb5QT1giAoueaMItAmkkQnJKLtCsT
gzXO2JhBEMFUirEvXL3p4tMITJGq5wYDTmSae8ZFzhXndMVCCfl7NTXU7QEqXd8Ki9sIB5zJonJV
g+G9/Gp6xOTVitpIwN/wIlsrAOeL+ceoazlGAHweHixC0x4AoBScdcEXKTh29uvVmzYEeI35Re8g
aC8JZ94BYqXBmXXih02dSNfHXv9SGJOA3STagAuARUT5apUDJKG4uJz8vpnUuQyNnQcj3iEpVwth
taJNv4rjLdVgXQM/yebqYYECGQupN6HlreVG7YAE1y6cHEkBwzZUjes5y/cRm6CAqXUhnH6FNAMy
EDoP6AEWjnb//gtk5FO5PfppvX2/A2/zFehHNruSxi3JjqdCXIlzsaQs3nIy3QMvwo8eyMtntj2g
P7tqpQxIVW0ka1wGkgvxgyPd4NSqrGhQs9Um9bjWlleb7IGyA6Hz1CdiTTvp9iSK/VwNEsLUHr3C
QFnsT/pAu4ewO7ekjdVQv2e8EhLqNytY5T0eRm0I8uzW6nsiSatFRSpmQEjthDnfbNYgZD+NVHWQ
qoXeuqwRmyLJAxHOM4+cMG/bTINwbOYLJZWdpTp500EfNGHZNcOkzDu3zwmGT/FkNt88czWtk5nS
lXWifn6b3W82/T8Fd8Sm1lpKF9e0SrCyEmgOYITKfCniv1BwzfATK7e6TUWr08svvcta0o1K1jgU
3S+vXFNpdt1kk6deYWzz4eOiwtwa3JdDvzjMqwO1NYNDx24JOA/vZ9ecr9ghr1rgr86p1swUf6Am
J4vZ0MOyT9ZfneiDv7VD/M524iIjf9Z5yaGiq/FfFyTHyf8pO+xcAObQN80Lx4dv3A2wzWFVtBEk
LgAETXcFvsKPxJgLjpRAELx94mKjDO6PlZOpU8aN/k36Rd8gFiKZL0o7EhfNKJovuUuYXd5FHTZT
a0+mGh2BHA6x+pT4pe9fvwGQMV7iqlpEFJ/bg9Xn+6OamPlvL20Svq1E5exKoin/5Kf/eiHveVeF
NGc1fdu+Wy0514NwChnNmFjR1ahEPli9hg0i8VVlYpHLfWfSXV1A3stXqX5W10udFtKH3sehAadX
/u2DMa5CrHJRTI467CZEwjwf7lfPLJlpbelItUVfTCnN3+Vh2xQHzvOV68ANsrcMu09aYPt0jRTK
2r1fG1+zyVlsHhKWhzCYPzRhCVnSmxRb3+4TQ+bWKSHqfX2IpVmz9H7O3DBq+g5wfWEAiXvHX0Tv
8S6QJyUogKGUbOs7W6mtbCOzGIBcR/WXtDkQnEGjSQb9LutbWI7cvoeGR1TKiLnMadNKO/HnGzJF
K4X4nY1irU+VL6wR2mk4NfHLCH/tl76haS5EoneRlIFnzUbMaZnD9SiNKxbzAtRZcWiBC7EraR2N
N6sJLWVa0OrM61Q0+w3s9CxVr+4r5F5zPhzfKxVS1ABp2J0r53XZM2EnlekDERE8ylNgPqrZ9lMP
x0eC/FFWDfsdpfBmwtIpd8MOfQ6NSNBgZLhss7sd7FXjj7Igd5gLRG+ctRvskP190j0SdPUM0vjt
k3orJrnaMGyFt9ETQ4yUykfEyyjhq04PqwI2VWd9W2f+ElTj2+l+WwNjn2SA4Lgeamhz3tVhcDCG
jspVyr5L4l73yz6iSr2qyrNLbuDZ7xcngK2+bRQlG3Ek6E96Cazj7Q1kl68DwxU2yqj7HKmaSvwj
Imnn1FtTnoh4lWFCWq0Uf8PN+bbN6pf1ho0mU2Ow7/c21cM0jAtdbrIkow19P3RuI77ddM+zGFeT
w01aH2qgCOy2b5KDJAfC4KAtBPfjs7uZfdLZkj0fjaEdsnv+3D/fNG4PhZl4cVohAweNSTuYe6pm
QQeI7r1zG3jMUyL6iMBx0xfG/8hltYcPq15+1FrxoDQwqaoAZDWLLNtGPIlTXCbCkcYaAwaYoOnS
eOtJZHIJ4z4BnsrFQuVa6vvlqsU0ZaZ6a7GmeMZ91486GOCrLg2RGPyiOTsTrjmuT5LUws1JadT+
pzw9xfdNMCxTVPruxoyX3B8OUYQVVwKpLey3PXDYuH6JI3KhC2fuGdi1tdk04vMDYyUanb6eDUU5
YJiMkB+RgjklaFUI6sz7bvVPoO0WQ/s1ybU6AlwyRjZ4ZbCm7LKzyMqBE7gGKUeupm4DwkSu9tvu
BTawekxcVy/hQBzmX7lIN1ZMW7PQZ6Lo48eDpR1xZE5QY1sZCFEZmnxtwrvRWO02fxA7HADKKEjM
uzoUwFX0LQtC29jF7Vg/vPagRAiM8qF3qNn2Ezgdc+ThX0spETkwwqVpvUbylfRH89pYpJakiSOO
KE5EmC3CWQUnzDSJgef7s+aE/hesFy1JX4Bb5Hmmi+aeWYJzv+T0vUOHKJs93J+lEFzzOjhj9m2B
IOW0UTa6ifgrKxPGgDv919+EVwZZ2w3fE+Gv4CnBla/EnQQHWbtWGzwzCtiYlNRvQ1VVuf3e0ZVg
4pwl64+C/0jLgIsSh771zemR1dC7Bfc5yJConz3QvfNBdSTun/uvVeQ/Ye+XltyDTQsK2UJb1sNK
kCGQsAiP514ugc1I6JZF1ul/Ci19fTTHR/S483qKLOwlGLusquwfUsDf4DscWeClOAzVNSft6UXX
7xfeQ5VCOQETOH+2b9/Cwe895PQ0jfMiKLXjWNuGuO+bYM0gkLHuDgPJkoPVs0ZWMzHO/GXfgdC7
nUs2k6qjIK8Sho94k4byOZie+rHGLKPSmNzLQ3ZbVpSYEqBJ2b3o7uP7uUx7h8pujzKijCxHsf2u
ltt3dCvHU/zZJhogO7x7ty5uJ5STNZ7wvbVI5U2oQ9fBH/lm7iWPGhejsUGzG1EnD0nTyCx8/8YP
PeKygap66rboGVDnlQ9aM3UoHP0eGXLPbMtT0IGQyRnK0t1RasMEwHVA/8Lh+q20h8GJ+e+wpIgT
0e8CZdCfN3YJAKBjaY6Hx8eAOTYdIx0eXx7ESQaqNMqvKwS1p5/tmGHysZPLQ5fDHSUVIR7Tq8v1
CM2zudAue65K36zoz07+DaoUlEOShJCCIrTV+kH4Eo2U5yD8Q6pQhuxF0CGsacDgF/j1qX6jssm8
UGO2thPzF4ytzoM3Os0GGG9vteHioggFv+UgFMzoRWcmoBBCIk9rC7HBnJikkVJWxmV0yQR2rx0B
2ibGIz7sU6gnwcv7rnp/mC66DMdJKkt1ERNuyNpWdaSEyl2mHfjgi+5Iw+IO8wKaKXuIGdGipKfT
M6ZJeo4G7HC71lYO/OFaeiS6TUio0iK843DBz3yDhx22Mqmc2aCj1uMyZgcwrFpsP3upd0WlNgOA
bl+Vlzh5vYUoq3X56EZ5AwMDjFe0WDz02x2WocpGi/H5Zh/YLrt1R4sTptTOnzhsY5MM4HCFTKHf
9sCIqbHj7405MZHUnnqzb1O/PurXJmzcz41HoAR8pEN+4AFNiIFD7DDjhCzQbJ/kGHQ3GdDVymDJ
zGTMYT44xzKHKunGde1kYWAbq9PlDfEM1WH6op+Zjo6AUPx+FhK2ADciSBNJRPQ3Wt4T1CLv7Mt2
sF8bIXERhNze6/lX2aomEbZocMz5bhOMX2Moi0nO8mUZzm+tFAch3ylQu4s450nPtNHZt09hBFG8
/NAJZyGGT+msdY9ZalCRogXqDyP+kPyANTaEgdDsqY19kU8O+JV+ijbL6YPSrCrijMU8s12xkQSl
CK/0Pk7MJRDO0XVDVW4tcBqdtreHiHMZ7EXw18jP1zxq9Da2ZaL9cgonYR70Wx/2OkLPAFu7p3uu
wR7V53Tga96tiqVTWAa1M8tqv/Mtl4ocNFWivmVu7TRIdaAeACG6iX9xX7TBfSKCTON3HH3JfDIh
XuV02xYQAsriGKwpZrc6o9XKhK1SsFo5wYLTiJ4SoMihpjJBP+CGbiLlr9QOT+scb6Ztm0DyhWBX
5hbH+jUGjZ6xK9gyQt6dz+Rg8NexOE/UkAs0uJySCmwuuiQ97dM9ZzRjiqh7XcCzdVCYiD3T+vJi
1r9FhOI7byN6BfR1+G9Oz+L1H6PLO9W1hjGJ66ZboxnFu9Xsfp2E+LQJHyx9wIIBBKL52R4vw3qM
vRse7piCrvgFAhulEDk1I0MvOTBAw1ZPkXvqUFTuiylCOvyURbHZIYBtc9XVGMtUDITNZ0shgAOB
YWKaFXJhfyqcKi3SSi2gZYo9UvwP5za1p4M68cTb1TMTeUAJuHjT4G2I5/0lIKKqhxzYbrS6XJz/
Gd4+c7XKOjV/kDwxfk17Aa5XuyxslHRZsz+uIoe6YPVj22L+Dvk94bkaTSFXSeweSXh07w+Amyw2
vEvhGF88UnAytQgPnY+uaCnff6V92eNjRShYUYK16AUROe+6X3PFw09cunXUn9dy6XIjkJpQVBug
N0YQckINqgK0FMRH/LQmE4fIEw8i9p9e9jM2yIPHgfZfydoTdQLrytAu2L6TWORzugnCYJkWx7NE
cilhsqcNXtgDktnwh1pYq+LJ49UTGvoNMzszqm/bWEgmgwKl4qFYkbUHnDOFc7JaBHoUIDrLufsD
mpmO65U2Yd20Rp/6FJYT3tq864xMWa6gTPVnKpqKmWENZCluMqjklvKy4Xe9CYR1zU3Qnod1AR4U
gfGtL1d/ebIYci+Ka2TUrMZNh4dxLFJc0T2z+Su2RpNBh1a//W1lkNiJ0Z9l/FOwg1cc/VyXg1VU
UliPR/RvQjQfYgZsUgxUJHCC1JVkOnqQvRZwMLNjd+XOM1wcfgKeEFOLlWfqJbrS1olapSJjd8fm
gO99Yy4ZW8+DNQ7bnaO3L175WWn102P9gpyYiO6rvXH0UqotTbYHDdUOj6EVVLnrv98AK/NfReVu
YM7wWi6PAWMQ4TPIVaUXnSmc7O6z5MSKnYJmqHBCVoSVISxvIAmAFJv+FcOfnk7LWgMK3GA/EE05
VmlyToUJscl0ptcUU8ZP8W6MZjc7/1I/hHmqsAg9VLTBAUn3uEQxHhDomb+USEUIGIzqTONDXwTv
7Yq43tnIXtCw2DNkmeVy8gU3ai7vB8CMur+SCkq4/wmds1vLmww6dfpsWQKJkNIcTsPKWZVZYGBe
npIwws2TH1TTqRtHX9ENE8CmuBC0wfaaQsLVJeXeEsfVAzSLJ3P4eyKVhuTo7BDziIarJH5VokVC
CTYGKpepJAb7RlKQcmZtf7IrsmZwguDXfseIPqEV0c3CoUC6uzw3RMjT5hDHfuIuhB4EgUZW7ray
uYCaX29Iq+Ta4+lXuxZmfqfZF00TnfDOdPB2xNaXRNQTxxk1FhdNuIjOX6tHHGLvlpnIA1lEP7qM
4bg518yYlENP32pLpN6Qp8F0bCq2I9cKfT+C7J3z6ovxxL6VyZE8RKOWOPuU7yEM+xeiCUzmFcbb
Fhy+n3zy0z2OKkCqKBUpbbbvHao+DtdD23UK1N+NZgFWNucPFxsucbdilOuQ9G96LAoXEkASbjET
/xTcwHxG8j+GL/jPxRrvj5ydZZF2vxDFuCxvCOdTc/IWiqdISuF/cUa+1SbeJKNMxqo4cAth+OkW
IYV2YK/P5hRTdeSLmYl+rf6lSMAnY5gd/MJKzsYbHBSvzsVdCuWiRB3zxiuvpky5WgjLORooB1Nl
ETcoMukoyLBoxdHPrXrqYMw9gEviLD+pWqlE8RxWhzY/OhBwxJIaixXVVy9SheYQgeG4ogHzcP8k
j8/PXzFLTxT7+CK/y1fgenOb3dWA4EtEm2Df9/DJrut38FTPTrxG0cMlRv16vcMILPQYiyM2q+8Z
gMdH5L/vEVrto3Aytel/HpQJbQcwJmX7tkcGoNYCXSdHJF4ZZy+whgPUCjVS7JFmXYKdqeZUSgrC
xaDxeCevTqBGrpq28Pfnuz+fjJF6q8wH1lvq95OGsHMlrLyArVXg+FEdqwUW4PcTr1CVfWKoLQqP
htOoHPgC4MZwQoacrI9uYPa7WV/VsW+fXkWdzppc1t6ANqN3qXEioh0fvVNMF60xgx/HO23CM3yR
biUIB++5nnLVt1ylV9ZTEV6Yr9mGpFvSn07tByQnVxMkOBZsMazKANhzGHEyxbR4o3gGDGo48NNf
7zw337koMGvJnyM/DYrK5G2yWp/pxLQAC9H0FcYDHSmn1Kh2bKjTml/aqmMJERYleNj86WF1ymj6
TMKKpLuTn7h/394b2/6kho3RF/HvHk5bYQ0/YGb0LI2EEJCo5WYITOudf12yPDPnsWIQF3Qv8qCt
Qtne1uWBB5ob4DGNEoOLOPjG7cOm6wS7kqJWkfD2FBPJq8a3Gsp9SOIsUt+qVS1Hy1C+Pyva+2R8
c/aI/P9mapjCyE5rhqP6cQWHsINJ1DUDWSYPljpGq9Y0/caULmUI4sip0cg7cHXOSwp/3/lmGEpI
N3+SfQxr2CHkVFiOgZc0X9TprPR+kIsbDZPFRQOgZ1yOfOo39CAOHxMO1gQFhurXnvioqN7VDRuJ
ps2bwOLSnmTn/2n0QbKNQTueFAHndJHPdraz1Po6fZxjsHHmjlk4crjWZ2mXM42CARqk55VQT8Yb
wHD/q9x6zxuFyJg31kq30NE0xbPnt/YIprbUmhjxuNKPoehszF9CwvGKJ9Gq2Rz1ybRsJHLjFrg0
S17Q8azNfX/VE6SmiQGibGj71gq1up0+Gl06OfUZJqdTifHjI+HVaz6fSA3HfgTmuHOWH8hUhOqn
Sjm+GcycJcaS+8btnIN5aTIpW29Ps/TJLWHHmCO8CiOW67Th8BliO/M2R3kdOak+TK33x8P0KOPy
LqeOnI2Zn9fbWGXTr1hWWWT/Copxpl06IRYReS3RTb+dqWAniMkgOvvdQXGs58/9BpC8j8/uo96W
zCR+0C77Mn8+f/oNjQFeVJOxuWWJe8g/7k/IoqOLQALKmbmyS2TELhdel5noWpCDc35Kl3NDQZFn
7diHHPsGWLHvuU743SzVh9fq/x9Bxh1AHtQz5IngFQX4/q340VgQmUL1iLGw9nN40r9kxrto8UJK
1eUKAZBHoOA8k8OREPfKNYhtmqHyGvp4nOu7Vjp+231m47MHgZkMte9EMwpcSSfeKaCBl2YvHp0h
Cb19LvcREQdb+6FI3HkjooDX43V7SC9ULN3z8XulGerRlw1ygdfU4qtPXQqru1Hl2XsP4Cn0OGic
Uauk7Loim3EQrgT758YcxXd+gYzxAU2EfzKzo8IH23T/ejvLzff5TWWer5RgbNMvGSrWfR8d/GDA
DNj6jUXHlC4ULFy6rcE4HP4n7CS7lJvQbYLtTTLgivFvyvc3Yy1VcP67eqQgBQ6VKvp61u015Gnu
NlmFm0eobe96ZAVebQpW9SDyt+/lubhnHWYrtkxzBfHYXJQj+DtzQWT+uMqHrE1awh9fHyhMm6Ti
MpA/rncjJbJ09WzFlnhI/xKvsVwTSnvZjuSs7xFH5zQPLP5NYOjBGwLfRK6Q4ogfdZEuCqof8Uql
ne44dOfKZU7Y0lFCWojEl3XTTTnYnS7L+CNCtinGbhM4NGXMybd3RA0EMjui7Rm2712fRMlM+x9a
1rVhcVmAIsMxdneeJjIydyOOB5WgKuf2nF/IvqFcScxXhJEskTfIghMraJf+i0xTaCjUK62opCJb
KcmBpknzZ1hZoA+N+ws5jq/keG02cVL5os95gFHYbxnecaoaYh7cmH3wZ82GfauGO8tqJMuDiPIm
/a7RdNhS2BgA+QbKBL//krnIKID9eYqURRoxqaJqDJQA0Uv0iyueIGDvdFrHMl9Bfes3shaKim4q
Kj0MKlPQzG/i5jktzkLEoACvdZ1H/IpQ/7O07lU+5S6/TIXLc/lJGfzJmO9d0Nv93gewyngSfb7q
M8Xa10dib2LuHr+8R55LdeNitS7x0AvCiLAVR7MbpoX0D6452ucSA3fz29Y4PUZgTAyYW5Z7Cyop
RB3w00p7/S9Jbc3Km7XraEoLV7eKF+XM1UixeA/bq5e5xp/KSB+u8lORHDY20ERl72O4eWNCi7rF
lg7+8rASmpXs/0aTfCr8PmDN9XkuZe+JWNMsr3VvqA1eBUpFmLDDSdjtpVjo4O05AI4HQznkk9V3
YJwWCKwLMHWKS8EWhZ5mATBAbnR0u76lhJzhaXMxCQgv5Tkx7mOsG5PTnA4Zg9zVedOQ92L+wywK
P8Lo05xtR0Rm5P2pigfmSn3fMALi4RRUArsS4cnGoBCNAa72tQNaglEiqHZCatiPn2Yq4EFon+eG
VmEg1aHM9kPy6g73qfceYSwodtRbh1JQ59scSEgwP9ovg71++Flj44C6EYI1ipRUciD3p4ChHjv3
kamFIcfCx99aOJlAaKotj6KbMFtA5kkWTy/IbY0W9XnKhIsXub9dtINJAG2jlUAu/AD5632DHzmA
qXgHgLIjieoz7cfaDr1FTpK1AmqlWr1MMUy6OGgpx2hTd1McEidJkS62dJ0H7vwxA9GgNtz61+ZX
lO3Y2RKrq71YmRytfsFNANR7F/M5qszJPzxVguHwx6V/Eckf26za1c8Ph7wewc6ucpMMmMPKr/oI
2f3x+VP5v6Kyyi3Rs5xb2fzqnQ94xhM+Uu5svH5oRLhJezja/2+QPjIpyo9FZPkdtPE6maqYURfi
umRH9eSfYWzOYRlNfmoQ2gh6NYDTZVAkVTcA9priVyhOJXx/VSYSMXGVBCXdZmqSGilKD9NVYErD
azLkp9/n+dt8uYbavMvHzOT7EYQSM8OyjdaI657lUPbLdOVYl7MdBNKsLkZDs5lIbocHZbmuu3c5
iTg/mV6HTLmyz0SpJZmW54Y0Hw6xwE5uSNM/z53eP2Z/Fqy51mGxfQ62o1EqaLCxkRTnBmGtY+4x
i4xSCbAFOgfNjNgNUCoHBVL1bXd2fy2CBUj4lro9CaVgRuGUmy0jZNT3DvPBtmeZCfcH/KdvkkvS
Lb+Gh8m2zpcPs3tUVxR7yUSZVUr7PFwlMMSmUEVgbhgeDTKnHXlcui+CvwaOyjoPJHVKHzTnYk6y
lWhNAc8KzDJ/1As/1KmtaLW3KZbu9vUUCjzxXrplEq8q8OA7M4Zhea9+7aPNlGy9kIjWPP+/n4hy
ieayy2jZ5tXma88avl/sNG/hjSC/dxhrl5NVYVG/mLMPMY9Pz4Dp3RTTFv04Mpli8rHFxVBDMPfa
uNqcGkw/IIh+kZvQ7WBh3Oddd2B6PYEVIF3WvVb3gR3uR2elbvSPU0bFX2AZhywXGgAXkObdpEYD
3DOUj+YqNMr+q2BmY6R7eHJ5sieihSBw6KrBy3aa8pdAvUwICLEiQpgZw/vCiHJpBcsr8AK6AzoB
RUSm4+BMlmk0IfEFHrRb/u+58pTDrnVb1HMgJX3pCnYduSEnBfP8f68XmVqyNo5Fki71e92OHpxY
tqUDfLZov2bQAOnI2I17Ll7jGluIlu/x/BDn0W5L+epF1iDeneumEBgkho0rINdJD7RA2NtdoRTu
Bp644BSydKZ5OUdweiB41nx04Orch+nC3eFY3FO/GSF1zzWYw5qTlmNcuLLTAQr1tyS6CKgyIUWR
zm4eflcAPZEoGKvsUsQdb37RdH2Cx8y9gLHcf1BIpIdtAB0+Pn+e2oMCqxCCn03+l+fwji4JplfJ
q5mbL3zwo9mLj8+iBd3KXbkxNhTewz5/PUan6VHa7zURKcRp/oZvG0RWKzVlHimpWGIWZNno/4Ha
G0M2iA9arjlcDSI0Q8dtJxNXf4XFlxqBbj8oMjUJ9EF3O67BsXo9yrPRgvFtyFA5Ed+69738sRzD
mkBdUM8UTMa7yLPSviT+xCUuZQ8yVxDk4tcPdSQjacshnBgV2/tdKM0n09ThantspjkoPQky5Suo
oa7Gir16jebOQUA+e2ZAqungpiYVRpSSJNpxueeC1WP44+oGv0kyc5qcVNaRGN4B1oFXAzKPqxl9
TsV1FDFkBZJjSNA0kdMhBW7AnipHRbLzdts3ivzfv4GHsgUmQYN2IHpyznvAtoHSPsJtqCTkAwp3
OlO1fEYNYx2i51BnOwfyzXW1pKi4Ayv6rhFz/4LOKsWAWVy5MjorKF6fRHGKMDwnx/0gBq+CjAFV
MzT8av5OZLnWpi8jPw2E2BuSkBvHPR2vpM3qxE7B9N2YNJnEpPjL0zgbbBl9o1ryNfUWS9Cntu3k
vP4Ew0rBDkG+nCZklcW2K1UJdZHXxpMnNgUhpK1LIoKcr7PRRpb9Epgqpo0PIE2pC5Qu7BmvyaiY
TqAtA9rTHdOWHrjFHxkFrL3e+Rd6qSJC+mA5RP1iPbRp9zQdE+JLeDjHpyrpiqRoqXqTuViPtSh1
CwVosh2lIr79oCZt4YBu/TWetsArKdYKQSguVNaRHXt39Qma/VNl95yTEJfVgcgd5dezCPhPU4uL
gz/42T0Afpf6d2t1UrIDEAVg4uGtWm/5AQg2s4dE3Lg7qip86ttaTGhx/FCSjyywPsQj2OFSLHF9
qtolxpi4fyNJJXHMQmRx8GFiZ3O827/sDDSE8HlET52qgnl1eRVml7H9H7UzGWwpDMRYYRGrHu2g
JOBmwFcLgkN3C5CXxRCV1FUPO1ZHQN65yBGQ5M6W6Otq4obePQKlIZraQmu/K110CNgmZ9Tb9iSk
uRJVca98zQRan8nLcM9PLf8Hr7CV6ttCF1McrnTKGXEPxpzbkKZnAJML8LtK1JI+vCVAwCE4oQ7R
xrxPLTRCSx1PNMUD/SCzhkPmlF43Gi5CgnCn+w1ko3SeoukQqr06cfn7jZw/Ii7y7vFWf1SBFlSA
t3QHk8XCc5TgADDhpuTW/5D4m/hEEwEJolmptgM3METU0azLaYMNZTVkGTQWnVLKDSRoTx+TYwJ0
e2pe+dmdvbhSNPx4xQGar6DeQ7G1LXvWox/N6px/m4WFLsP+sPpTSdifFLLdE/kK7Tko1fD8bS0R
M7n2DzTzFbVt0j1s3S91L2M7ZCxKxFKCN67eU19wpqN76xRHVcPh/atMFcXX2IBb+SanpLhV5/4P
4wmKRVLnkjJZtDdSlUp+P3N1yhEx1lxTy3xqbplw+6is1XVF103I2hkzsMDFmtbWzcm3JfPhrv8d
4lrgHXsseO0E9Tz9VwO7YtoTLDzDRK7mFIIyOcs1Y2Fw/Xg53ZaVSOLYqULTz2r2Xpgg7QkKVEBr
jGPPffWcpFggtTCsk6W0a/D8eZPSFAnB50TsnigkWdn1B8klXPGYQ8nVR6UDpP6tsOfzRbTr8uK3
VvRI90gYmdJcgzfqWdZ7XpPU2G4ziBejAttc8tJxFRgMLh/WyhHwEZVLfh0cVNOMm+NDlSnUtIHJ
ANq0PDMZeiGEd6Ily0WoWpWJqluC3Xg0yW+PlokgQNu7nJLsLAdEIs+UbvYMw7zFuBs0LeqwDdYh
qnmQAtDCwkkv0OeT8HahJ0UAtKtIATZkYdRmk3u7fbYy1C9PcHAh3SaRDATxRkknE9rUcWSMDYrW
LfD0Yuvh+0hf7aI1h2W3YA2sRxBeWD5pqAlyAkmyatGdzWZEbpu0ux/JiTsA3vEvlKV/oNJOAkgF
zGMfdzCQZpKthz6UCdTrsbU1GsApPjx7efb0PanfeGtqv3RDbdnuqZZOZyhRhXZzXQS/HcfDFMvA
NhX64gCF4vYwKt11S9AhrHvS9ErE8TwqQOvTdLlmlS4qtKb4e/f7rpxdA/k1I6VBsko2S+csSaas
JBg+VWoEypYuctvNIcpzQmNVMmjeMKX4qd/yjTGEVKEHKPifKHU/tViEu52AYoHaJn7yu6wbdf73
rJZuChrH7O+JZ8nMgTtpUeThxok9qk25jv7MkbzV+uVi5Sw52X8Ev8xhYuFaZXFX4QXLm+RW9acH
8sU9JE9dka5LlXQz9cy3UcCMPkDPGpj2mBGQSn+cT/cqDxcMUilfZ1BaN/M7Y/B5WzyqG+jaEfUS
wyMjzFX2kK2KMrxSAXtnI8iwUlo74V00tIu5PeMTDduztHSH8t3Mn7fQaKZpAt4bigjDDnbeVrOl
uumHdK1ifiga9VvO9+0DYFva0m45LMs5GH81XBksqxvu+u99SyAUMc+GjuBPLBjKqOW0hhp0ww+o
eJ3G5g7eJZPgMtfq5hlet+CtJ0NGdNN/lWydu8TUtdFlquKE59Jr85/TodDQ0Z5AO+yXpD7UrbVo
ITsjW98GV0nwalf/JJt/+KoXhv9o7/1lAlMjyMN58hvcRxs4eloZV9iHbZuQzftHIy5o37Ss3dpl
ZKYu34bBFy749KpzKwkVZHVRwVyxbrF7vN4FH7ZnBWQeqKbpstbmUGP/Pzhvmp2TQou+JLolLQv6
15JHZhqc7UbRmBZxdVKhU8olBsa8fcNwv0FBGmBp7O6Vc5DgRORg5yunQqmqb5f1bkykHUlF+QKS
P9hZEoabjTJixwNzMrm+I5gyOol8GAUF4kO+1dvEnFvsTDkNjWy/ViJwH9hkF0UytBkqaJBzwH8Q
pj7jcgTYsjc3xYlqtqv3fPfKAr6/SiYw3Q1mzZTqwLVOMUnrf6eHGrGG81vNmkAUfVG0U25T3iMS
xbeWVbA7335ZGNSW5sfWct+qOsdQJmNnLzsAN/DsvD6E9MUouiG4X3X5S+7WKCsr6Pz+SvoPp1ye
8efnH5fq/9zgf48l49p1JAjjq8ocshtATCbVQ0GOd1VCSW00cxWbZc8F2tBEJhnUBE/hDVgvRDwZ
/ySZLPjA0aO5rrqb3+R/gVHMvw6MnD6A0FWwC46nWz86PSfxj3RL/StXJJVBTU+XQV1j0CkT9puc
VJ0BbI39aUalY5mYDvAScxSMLwgZOWEtc++mTRTF+gMoIkr/TgULkfBHUN9/wNg4uZhvvgnoHbu0
Zzvj+b41vekTUOf1+Ykdulk/WvwJZTbqUeXE4vE7YmkevLUQD9lTt8YpqM8az9w2SToin+6ledxs
3p20fsdRINn5FLTtj2yDh7mruXYuZNli6aKjVYDc58YX/lySE8II9N2SQKIIQk8FatJffZuWB3zi
UzPyAEeq8WxD51o9fiGNM1rkvEqtAgQn3i/FCBAPzX0FGrB05idt9XH1Ov7wLWEHfour6ofHF3cO
CJq07obyKgfgHdg890iX6L63BRmBah3SX/4IP0k7RWLowN2wmYTNiCjjN5cCHHcgOUtVbx7H7UcI
CWeBlxRSoXmOWQOHPTQHnAh6fyG+E7j7LtP6xSs60p2cyKYsbBhDQBKyQQOSEPRFLOV2ZELQOL3b
ZTIKnBSXgrZ0By+moRsoTPHe4p6l/4VcHJ6fnwv53unEJ6VfoASh3oB1c1xBtjRRRSqmK2obd3Cv
Y+TNMT66nF1czVJ/3Y0uoLXIx3K+wsHveISYVtakBHe5JU22IinhmeJqkA3hGpbB8Ed4OigOcqtc
j/5MOkG5jgsGLJ4yJW7XmkFNIioPX2XPOop0GX9q5LR3CtuB7I+J2YdcCpbcvuQ1gmCNoKkWBzTV
ZCP9c4TYKKt9h2apUhInT1d496FFJg272EaWIjezc2HAJLHa/Dqdad+o5pr+XaA67fgKeiCFjaMg
TysZrnrmu8j0dRXrjUQq/JdpVF2wE35hKtgNHtOg14GWRYYYqAoCBna/vFoGNOaJgG5kzUUNdd9N
PNfD+JcsiwgSo/T8HxKTp/jU2qz+J5dRwnsgPYnKQVLZHS9bmTXEiwzPwIofLgv2c6YazIBYUJWI
7SxzJA0FGfrAEJkQG4mTpL0EIQB806Q+W39+ip60v7dsoIj9MwieK+8SG6J568uDsjbbSFm/2kdv
hUBM6GQAadvrSNGSAAXOQhR9jGfntCLQjeOAvbcE72ioDvRqikPe02rMfap2MHiWDG3HgWV6iAfC
M50nG6X2eNM2Y/7cPTr0PEtP1RK4XnWf1afRn4w3xS/SzWKqn32dzwSyjXaY6Cj7HsiCHWfWufhb
tUyw3ONnb1CaVfwjHr0X9oA+b+NWnfaj9d4Hx8l0zjxjnv+oQHII0OBdlxcG/NBPY+h6fNYjB/9u
SyBCzUD5nZSP3BI1JnJs97l/J7GBn1mnLXERr3r04U97Ynz4KnyZ7J859HIb+HxsHnY7gUnNpkhW
lKl3Ub8CR+DcYkle/DgBXE6Aq7WYSe8gvP9ekPJLg86jUam9oVhta0Nm5rWMgpoAZesfZKEbX3jf
YGGFEj8VL4RLbJVFIe3y0tTu2lpOZ4qnLWgza0+/h4zDBQ2bSK22lOFUPXHC33g7U8vnn/M1Fu5m
fn5pDhnK1OCnBIr1K2mvc462SQxCYFKRKb0l6IQzkqt+Ja1xw5XRkSDv/g/4L7GwfrhuZCECoqYM
Tw7SZEJRjUQHBdkDoE7KSbB8jWEkD4YCO5ZJn2xyK+YVfOV5ns3D4bRexrSYHm3iyoh2TpiqSrdh
Y7Vnhc41fI84qZ3BH6+n7Pc62Udt4nl2lj9V+y7QQbbm4eTqzgTKWY9CLEs/LHZ2j05LOMnb8ZN9
i5zsM66zHNek77Fi3D6JPxr9v4gET+ivfixdQJ75MuS79Z9UxsFNCmYTM9qahqbet906JcuRZYV/
rbdIbfmkig+Al73S9LNM/2TyqZ3CbWlAJx/EQvVrEKBHjEnVVlgUPpCLNcG2EDDhN2WpJ1PTShkI
9/l2fj8QXZ1mqEfTrV9R+5Vhp7Dg7xkYTmWHTpOTSERF+syiYLBEY5Mv/t4yLSrWwlXJ6H9Ktva4
C4pcu7xP0OyLhuE/ZT9ow4HjFBVHXXjY1iNXjNw8Sn1mutSr4YvnZ/DYtYSZ45RlPws22WeYoQwg
hSBNTwXKY8FgbW1IyOgzK90K6X+wLZyzeanM4sv3PqF0xZuzzxI/DFv7f6WYbCkBej1/5nDroRkB
xPohP5ZZbaY6U90Bx3zFRQHMXOjffWKfcEbWoqJsBjTgcuZGyttiniZcHx4c98whFuB+pY+SHFsm
nua+1juyxS/tqm2amvMrpmWKBzizByzMnJyKyU9KNxyeCCssT5pu+OeYOA+tTn2AA8q1xj44LvNc
jWxboWlsNkvtJFm277o6PrcwIl8UvnQesn2Up36xCfi06563CAgbdkF6Pfe8VOvRYD6vpok+E5lM
FsUWFTXJVh5n6xpDl/zH47Naad04TAsSx/hdi4VK2NlLa1EmjOg2HCfmf3cnYTK2agS01M+UMumo
IKoRaMq0kU8ufWaLB9nLpVwfyJWY+ckcCoVylGR3VoVPmemImZlpJurVnayks5Mn4yfKSGMgxuLo
L0DIV6ZE3sUiIhMfXiG4gSpggDfJKpc6SQ5GYzhQMk01RUk7y763qoJvn3TXjo8kPJDLcG49puf4
5ZH8GNFQgUFjIrHrkV2EBEhqz24aHYMh+ylkWnj6fPLLd7TBu9PzNhGIEmjO5aBOitSyo24r3hCW
dJDUI2hiV8JcHyhjuV4aLReC8inFJdhCmZR5YNXPftZkNOf+pnJoKIPcLrXttohFR1qpXXqXOx1q
CkYEkerQxTAGz1v4V6N/AsNk9jpce3WF01UeNRJzL0tuR0ltzm3Fm2Jnr+1Gu2zscg92lBdBLA5i
tYeQk5rWZMuCFtBbViZe9xhsFNF4JFH3ybFDKZLX8ZN1Li/ftpjnNyC4HJ65xCuAioLqi9hjPwua
8J/u4wnYx9kP0h1z4hn3r8YxdLGvNeMDc0jgrdOCR4fSOQX4zUlPEADs/Ca5aOsQ+JHlIPj8mJdg
AT4UGphnuPoCaMzA73WNVGiiFRfqOFJnm1edAbyUBYVG0XIMPyTOEI7wL0VbvXXvHU8Ix0hfboku
oP0ip/FLMc2K0kgaFXfFgkVLm0DUPNnyRtDMWB2QWma+f/zj5b97OkVU3Gkb0VbXVXa/tWv2qeUB
iSHDdR/WucjyAy5tqeJOLLPAZ2FRfAPo4lTrS+dUsLSu5QS+KHoLcCqjGV3voaSqDTuQYOEf69qm
DzGzIwXUCDexQcPGaddt98xCqOutCZr2Lz32nWLGL2LNk3ibqlYbwA4YEVRDfp4I1CtttXYGT3xo
fQ5L1StYmTnUy8PaVNNv6N40sQH+Xwzs5SaS1nGIXkmCI9DhYojn0SHoFkyNAsxSHyKidb0jBFEu
5sPCpJ7qZDWLuHmfizO4uR8Vm5+3Wy6nDfKCVN9rul5kXf2obZxopEP0CR41NLr9Ea/Ck8NLV/q5
zDOPf5aMIK0FkvWp8PwhKxPRaNHhFXcnwAu8xN2jwxrtLFNizCj4KAth8xoIJWr2ByAHjlhxVc50
pSOdPRRi+VzZfKJ6qF8z/tlG8AOzEQG1QWuLP7mhh0nvxLC1SgOx59cRSVMRxPg2qY08hzCKmGWD
hkN1NQcw2r1cu63karFNRshFsuB8bpz8jN2JthxVUMOIdUN8n/+8AIiBQIN0Mek5aQsD/DCt43tX
DZOYUPxb0ayBEudig1MWX5M605WkINMbo6TywsvaWAigPOr58uCfl2FP6Y0R2Q6gCxtPd0a3vvh2
fesarFq54JHLUBzaMoLOajM0luYvFzZSlUlXn8lQubnU7SU5eQCCWwbw2wiMJPV//35YM7OjFYdy
5l7S/tj1/Kr7Woyv2nESOWDX6iw9HFbkzSULX79lk2KfOgqVnKRZcCa659VM7Y+wt/6Ae22Xm+ad
r+giiHfxbdazw/PEsnTlox3nAsik2EA0Pt6eRUgjK66Bto/QYBc2VmV2F/5btk8tY226XSo2Zl/Q
aEN2h6z/5GkfyYZowVEN3OaeOIwOGscQtiFdYPpXNWfDNOndUpwsFGvdASTEb25GWgMmxzoMy5QK
fDVBnZhWkucDDpu0BQhJAM4t8L8RU/6g/SpsJkSOomKVIJEhXIKv83xh7UBHUyxJPaoksedRbJGm
FEMw5JXu9JrPkYrprpQdYqgXR+/fply4+Sf+Bj+LhThUMiJQY8YOC2BFdxlxLagnH3dz71s1frO9
KUDaKk3RnAGlgPAIFn7twuVS1anAfEzJRhaPvV7CqkhwgBOBCuezxSrBaUSeTa00dYfHp0NKC4NB
3T/WpOmrxAHEjsmtihAu7XDLVkfJnTK9GNA70wU+m1kATFoFhlSSoCwa4wk9PWSheg+EJEbTiIYC
jlGi+O6dWN+hMD/VKg6oDx4OIIamOT/lwzmj2kiba3cYptjn4Y0OZlY2gBPVBbBvfG9j4UZoWfMG
AJfxdqEoX73pFwzar/EtGs5cjWoe22Qw5ocPUSiNFBsqJKi0mYaMsyImfV49IQHopQ6IsaIOe6HL
fLJxyX6PDN63o4nThga7i2ZgkInjrWVjbTzeHtMvp0FohvgvtrVKwVAHa+rj4QWc8AOF0w8RkkCq
21NnQEtwEsIvbcH/k7Feg9QB8BQCalrvTu7trGgxanBxlHOmid3U1T1LOxyJrNdolPfJuNBWjL0U
XaP14FJYDbtK2Br+y/rYPcva6M88YDK0mDLh4ma19AXqx6zIvGBrOSYB0/03gx0AadcoLwE2eOP4
0XJq4CatCSGm+DhQYBJZasp74VJIETuNkvJtbqzKlqSZ7fJw1k27U+87maE+bppbvZSqYsYN3HUk
CNKkQdAy3Um6QD+GohJDtr+52ZUOJ2vFxnrHzl7UL94wBKcoe01L0aflaWsFvkLVptw5MmV0szFG
Lqopu0n6rJyh7ExxjA4JsOAVPK1zw1jGTNpx8CkYnqVHNJ3mIhlrfvoSQ89bm3IJPKFWTBMehuOY
3K56fv9CWosiKdq8CWkkj6/5zNeBjl/YVkVjeS3ESGQ3BdODMc3oBjiv5XMUkp37gxvHwWhGfu51
Imynes+tiR8Cgm4BCbzpwJCSVLr9zVbbywHTGsAJImXKTKiZRbbQKKWqMRmU2kMfGN+e2PVT/suU
OKAHz/gAY9p473ZfMGnCG1akAhFIWV3BgmIb1qh6ZcAmjPSobE7x550fX5PfZCFImUdKS0wIJT3p
CvKrUdzXL/P4WAvw/pbttsJqJODHIQu1dOHIrnwcDTricjLQm4TL/asNVMe4cgCR3my8s7mu4/k3
74R63PD+RIOjmukNNgckfnHX8p7I8xL8QOiCdcBqrA+vA7F2WBh4KrHL6t/ZMm/aXqaJtPHneQrf
pEL6kTwEv0rU8jzeITpqN0enQ238vqOZ+P9gz6daDUPkNuwXiCJm1yJymb+kybxg7imX6gCjvWQQ
30uPEReWVm7dsJXmvPHhUIt8XqW0EMu7h7yltSQWB5CoQuXQjhISXKTG5cCioWjS8oLzB14aPqVH
Df+c+yc8w+IttEbijUU2fa21/hp3AuF9wWccd5ClLoJxd1X6ZyaPHnO3jzWTcAPEWQH39k51gXjg
HR8HRpSJetkh9n70eLpPy/3HW4K/tbGUoeT3Ur/UiZImg2bmOnZbftP74NScwvw8j4RAwrXJQTSA
g0dH+7MEHUqzVBbRK+IG+cB6YweK4S4LG8QvCcOqWT8kJpx10l4UZrqSLlH6nytD4HJt6WHKBA2Q
uqaJeuj9DgnKSYwHAO4DvLE3zOYmSFuIgR+YXiGm3CY36Ez4zPWaGeADqBp0b6AZuMq7I+ZppoJc
k7h2l7wXzUUl+lf+0pr02eQuC9FWJ6kmbbEp8JRM0/1I7ugiiNl1I6EcGP8OC8vOoVi+P4MvVgcd
Qm/FceIwBhtVF/+A/TNcicYvfONmnbQg6sWVhhRTJO3oVCsJos0PD1guBzKfEKS4nhQJ0nGnM4Yf
D5HQ/5k/sTBbUgdmP0HsL59U4IcDpw9GHY3+oPgN1qXrr0DLav8yHlpaRYEVqjPdKXUn2dzRdn19
Dhoqvt+xyxTNhPTqq61zFypC+pYVCN7+OYAxPzZt6jhGNnZOZ/anHS3yGox55iHTQU8G2p2bEyXM
GdUinsEyAwhiFfk5r4QTwEDRh/q5on3FBh1pEf14EaI/13Y1IjCsRRqKu5CSvwtcOid6mS2Zh4pa
hZHuTREqCMdno+0u59/Y5sUAZmV4C9Jo5A8nPzNxdOXL3HGMiFtWbEq9qHqcjsHw1BtoDWhlRrLF
gmIMci/65NzEG45WbfZYZ3BP1C/vs4xLymFlblfb5z7s6y3KbtR17VNdc2j8ka5w8zVSNwaBjyuw
r90RWe4RBJhPrVDGeEHsrw6oOo/xRPgbaezYPUc0VdeT80LQJwyhnIlGaOoJhnxVvZC7R8lwmtOa
6z4PdA6f6dWm+fmzShED61lUv2+vfi3sQdVKvFB7UDC/fGCHadGb07BVl5kyqsR8Jad+WFlKFloY
bMiUhey9Q4W5sO2QdYfS/iRD006BgHXlxoynzuYwo0tGe7vYtx4ifVpt/Sff2gIkrz5nt+phSvl6
mLVItIEjjyUqiA200ZYI51VBQqvXQbSDaFZ+exxX+DN5/VuRZ60XmZyxGjbQkOOvD3UkaAc7z1sb
J67+GZVcqVcZSxe8elcUcmzhUc0y0KOyTLuYMxelFa/awgeGa9opl8we7iIZDEhFpsKPQtW/a4g1
PJyAgKcGH/Gh1jiwMf3f9iru7E6fgcTeupeLmqrr9EneSOuLVch8RZ90YmoJ2cjmgZi2PbfXY+kk
WBXrY+1PF1QOkXcoIAqH8PbN+RIoYarLATJ6951rCUl0/F8WGZEM2KfKQKMkSDG7voEf8cpoWlJ3
YS417uTc8BWy+XyitjtRRToK7C3+eUZCLNign8vyZl63hSRjX/PZwYojELW0EaMn2WvzFzMsFZOv
K3lbelWVya1r4+1xGG4Pccp4O0E6pNs56oc8YasLkYZo3IgfMdiSB5vSnQ+gSLzXqRGJHdxJ8FCY
YBmTKvkL52rZ1u4HvZ0ZQNnBKTY1nO9Ul2CzftyctBhT6N82Si4pNAT1/BVgMudXuCkWYfVhZ6LG
cnb/xh0XozBwy8YGmYV+tv3g+pcE92zAQ544W6a5Ifq6RHwe6IO9xM1EyCaR5urUKIqWlfpARhrz
pfkeT+IcG50QHeamkI0+XhbczwI+PLD0QqonTzvp/Q09OvVGKtFPzoo9wqkJGrsTZmp4s5ifj6MD
qaDZVrEXNY/2TNBQSq5ha8eiGGvvG5Mua8D+tc8myjEjGjxcaVxMU/NqnQJlH1U4SEu1qDN8YLpB
56JgtVVh7VEhzZ1PJrnLPvJCWz3UH7aMB00Obtb5DAz5m+cQgUPYjKDThhTLiN/wPPbDsUU3jxH9
c+Pj/32o1JbGO2a2MrllDaaBzDtho1ae5drgqOT3qMZT8WhTOA9GOnsFAf5tuAo7uTkemT4esKfw
oJPCZy4A/Wurj5MUVebY4fSUBttIbS/HY+lGH475noJgKT2S5DO7PEcVzmGPJ0DEHETVYdc26/oy
tXDuod8mMpM5MlInqtor/3Yi88tZCL2lilNzzQWaul8gLnulrRsxsa93wqEHGpnW8m9TnMExXXuk
qD/Dp+iNmSvBLh9H4451vUtk2A3KIhV/nXEHfUuK/HceYgAKMcbS6L4Zwjnf8j5db5LsM/vizGcK
x+aRG74bBU82DxRZ7EGyh8WZvujrmQakQeNldinPxdp9czAaPZjFPHn3lbw9sw4+qfnPtwy2VaFz
NO3as946v7DVcL2LijqkrfBWf3H7RqoUnxpotUP5+qatG1d4dvwerCxiziGS1jZkhj3xkYVRclc7
HPAZK2jJEjCnvRDOYR1WBFqXiQZhzVNy0YwXBrmvRYktBi3cjXzPF3mDFQ9YlPr3SVSlLOeBYbid
1Skj7lOHUMuOZzaTWn2hubqW9ve5H143pCLiIBofOI4fBvLgPmNs1D9tiG2RctLuYKybA0xPMtKg
I/455Dp6uGDH9PgtgeDqCS2qHRyAgUIThNDct4jPWP5Kq+c7uZf9GGsmFTZ1E95ipxMCe16FxipE
xZOyIrneMir8IcPkubyaYQWfE3HU3uHKQCE11Z8zKC5DnUaR7VdLnGhajESCgBPHO20puFt3l060
fLfjZc8IDpUwtZnnm5IwB/Fk7e60SlQd8KJpa2ScQEmcapOsT995XONY34rjJaRPuSREmPmT9djD
SZP4f8k1y61muJWUgYtTapIjl0y/O1OcZLHBv1DcEuXPvn5lVxqN3MG+tXQzyYw4zlWC5mlxMe5A
uXsL87f79jIXFImoRLd/fpHcHdnPAAQz5CRE1xGnI7e5Kre0YKoTCa2YDGapuNz76T4xOpgHK3ff
E7Y3eY6+dN4+ZEW9P3grvKPULZ/Req28e/TKNISH8eN4U4vytalra5GJPJV2UHDUjtiU+LpYO77c
Y+THo2Wpg18D5t90MYKhLeG7PBkZAC9dVEiodzHOO17wccgN/jCPtb1T2XwWVba7H+CGMo2TUzfQ
kXACJF3KoYMQqQaM4Q6csifOHbHVWy6FG2Wht6mY5UtgJjnd249BjrWw103UHlEiZL59sWkBVZsi
aTQdhQWyc2m0Qh92duNeB4R1HTmuxKmZ0Py/rprmmkUQEZCgw8aEmPjgqdZ+ALLTPOlurnbxrPd0
dCcPqBZq2e8o1wUr0RDrmEDAn0s/gdpkcTq2yhXz80MzdmADdb4/9YYFbSvPGmj9uY7l1F1JMBDj
3S47kyPWAePEYzdozWxfspBh4oBH2OQbE6pSNnuUUrGXrDz2QOOulZv99LAzc8pnmsF35Zx57v2D
J2OcwnkLKrEZ5i3w+PLpAu0KHhRdkgXAKPDgq840cPJ/au+t4tkCFNs8xHpikqN428ivyNgr/elL
oKb8x+q4cdp8l0oBrix25TMP5JGhGhXnMXdLk6Ay/UddRclaQ0cpxxriuGPvAirRftnSKM1SKdf8
Y/mtzhpnLZiaRGdiIRmzNc9HURF0wdxISQWkJK+xBWoX1cDFM/LPmHY1qMkNaJEaCwso8cT1uWK1
VUQynV9G9M/UWLZeMpSg3RKbpKXdqyKXW1Oif/RkRrx6GaSMIc0K91aZP26lVHILg9z5vmtlaszF
N6nO/rmpxjNDBk8aXrf+2tVx6QZV7itRd/ozs3BXe8Rp9n7EoSrgWfhrqpEBEFSqFv9PJVGU+j0v
jScbb8n/3XSIMmhX1zzVduAqL+EfIyXW46sC2QA8p1UohB1JNf4k2P5bt/5Ps1ar6ikFtFvTGXCA
vCQV76T0jG3MlY73F4RQ3Rz7/xa0tSEGYdbacKza9B+8CQHBVkzzjqPPJhFrUDyFTTgLb4W+uXKC
u5iIFtlUQLiZ4PMZ4XAB5oY1I47a2FaRpSdd/PvVmnUFLw8JoN5kYGxiF99w/p/Db6R3Td1f9WGO
rPcpw25R89hk4PQp+r/pLrtMWsC/F9jZw0cxXCnXczz01LhoRN1df+ls0/2V0dEKGGPr856qTeuX
Z0i10G1DSABXAWezWODiuSWLEINU2jaDuXWIgdGvZFQ/2Z95TnFUjOqt204loGT+8Fx+SCdqJ/wy
ON8i4bfUFz0vS8+xsUK6LLEyAk2p59kQ18jRUoUvzM8gYCCgPjrmZrmrZfKKR5wCtO+yWa8W/QJU
X3omIjCbbGf3zF29BwQHXkbYqhg38sWvxS8W3qS4zb0RPswMF311iYbF7WdCmadyHypfOMq4Nzdq
TjtWrGPJUjly2cN3GB5nM3OHOxO8HpSpHQdKtTEnY94SYRnqGajrvw9HKQd0MltM6Li/3HAVvcK0
S+in8X1p/g9ongxhsQEDLKpIsIpkvPhMDLW+9oa1vGfSFt3ZlxixFjpLSOqG9aKRSCXOkh7lRMJ2
qm4qGVyrJC3gsZoCo4djp9N5TzHv5jDvlkKJHJZnqrkWBwhawU9/i+/mIntZLPEeeN8bewGDa1Xk
7AeE7KFcTXdXS+ZwxyOK+RIQJqI473kqV7p6wE3Rm6YpUOQCpEfFUC6KzwoFCBcGm8OMLWW31UEP
73vR4shrkH61uwSLTooGlUGx0rbOjWNKxmKVHU60odMi38EyjMeZkuSiAwkzKxP/Ft8axezarkaA
dzfd5EgFMfXMHXyBeitLYNjcEeGo6Y0LesNAraNTqsiTbdESMImUvRYIeE4ywlu9lP6kQaT9ktzL
HO2jXs6sOlE7coecKbsQTC0lVBhegemFAs0NRErJh7X2RVLjmqBj00Z2GiHDlX84gjZCOy22b5MK
acCv1lYbusR/om1iOby035Zym24gteiMYujvnEGUszUtAzQ9Wds4rwBFUuSb1ADkF0FuZgRGgcQr
AXU5dCPQMJt/EXyJSDPISrWupsVZ5Z/pP6o+eONxccgneisMf4BLWgVxUH3HJsPIyewz5GWYQI2I
hmdAT3yMzuYS5yI8uxQRvHFvfnhyu8A9rYCkdl46ocTD2lX1MK4HtAjZEZF+hSP0J80w3SpmdpBo
rCto/gmMCJEa/FUKa4M2RH+JahmKlcw21WmFcuwfSzLDLRlvO16dD0mZXknIT4b50IVMfc8kYljA
EVTiZKcwLSF/Mg1MOEMPV4murI2Wrh8XskGHrN9UgNFevFjdE6QxjxH9W7Os0nYgDqTpLRF/E42s
cmWceVioIdrkqbHW4xDFQW1b57ISdhbLerg3Yj+ebD+53u0JuHvcwQClZyJoUCSqhyEsYJsufpPv
pTTBVTU1ubJahnpHQ4KKrTdqmmv7/HjxFHxxaZpr6p4nMVDhPxJRBtLbhHcWZ9eKYR19gZDUePvR
HtkyW8eDtEhcHJQnYTgnZclZrrD51lloJQkjRVSR82xTA/02vG/OqyN1giIFGlf+wEWkHVUhCiH2
1Rkcm3VuJVJX+GWENYw6ok3xFrHtmKbNPXsQ2W2OBxcWEhG1RKmGHRSe735A7dpQYssK9+3Hg4l3
qHjjZAdMhb0o0kIUzWJQftnIymVB8en4iKIqbokWRBMOAuzTlCkloJ6AnnkBoTgkS5UuUYzNfmyj
EiEkCaVqgev9E7tHIiFpYFxjGFPJ8BVSrKYFV8UxWzFCS1tCqHIEnCi9rMhgEqzkjypsfTKgw77L
+UYwLBvI6fxDBdBQOp4fN50alJ1kahtCzyF+L8GTPCe4/Tl1G58ZS1xpX+izR40+FKPDQ/spJRHe
tse3u4mC3Mf5cxU/G+tBeawm8Sp8cIOd6yMU9FhRfu+F/SGKIIVQXLlo6MXPOxoKMRi+h39gxup7
eHN1F5tMraUxUSmTZNixKgQ0nC5uYVdhT8/wghHVXI9cehl0yM2KwDZpA3ZJ7vFrCb6i62iwwA4u
GZP0OUEKI0X6RqZTF0qCZVJyuwQ+jA9O/R8B1ZFEVW9JT+FufcAZZb6Ou7HbMYS+4WacMU350MRp
lrRwYhU19Ki76JwhBSng7lHuzz5eEOg41rSVQ6q6JpXd3/HaZgAb/mXyqrBX1v6a7TINz7hW94/g
VdK+NSZDbq7RK4mJXDvGA4v+9v/UEgHMO7WYqEZE9Gs8iDhnU1yUUSieAk0XdVdkf3hAW7WOMXKb
kJEKbQDUokh6mXwVSsxDD0U0gVzJTyS5pmUbPBcvny3ZBi5CXkX3hW6zw9Jjh+0U/OHBg3z0SD+B
fJr4KQ0WaQjpHyM9CbIDRGGHv5KPQjCnS3Hz92IHcJBwp6zAAK8anrORXSh0mICqZ6pTlpw57UT/
C0hOK8KD/XK/N+PUHocutCJC0vBdX+Wnc5E7mavmisVVR8C/f7yLTy5d8RNMAg3K6qv71u6XN//i
QXQWqlyL2hv6u5sqOTAAshwk3lCaw18zv2vPnGZO48mf9jWl+l1Vl3+tYSOYVSrPRzS9RYNc56eU
sGe23r5J0GI4aMn+yhk325O7jbfrPTIhZ57bl7OKV81/TBegvQYoiX0bt4tjX4BkD4Bn3Jbd83FM
o1Z+tHOnoS6wdTCrtAqGJcNQUOjLNNFvfhl++dYpAOW3k2pdxMHiZ6r3aRC21L0j2ld6IgDzUSPv
MNq30npxDqutu/6WFwzElDzfhoMHN9ptndDD1uh7YymY0IEGnd6YQTpQcamEMyj0fnFSPPO5qxES
ByA0sTSsA4IgHVatN0yg+PwDvhxqapG5Vmh0u30PLUvdWhaSjoTMOwfDZNgojs3bgxj3QItFUqtK
q4fg54k6f6aaqMuUJx+irPc8dJYWK7eFSA4uY3yWABy71CBLBQqo8n/BfksYCniOcrt8bb1gmey3
rB1kKBF7uJQApQ86RMmW0v3zPpgKZTdhVMO4J1akZ4TzNgGlDK1DumiYqHaj1wD4ColU9Hwqkrmj
/e4USTaPd1rR1nfEAo5DbpZE1igbgoWaFeqyWAVDGIH7uQ+ri+dQD6LSf/JObKmb5T2QBJTF4nzt
jn0UhiUTHMP/YcN9Vds3ZkJqncynzhr7yk1f6kf0peltJyiHcKayp9DYR7uIq3q3f53UDeu0ryIR
pRJRm/BZgjBvopV6+s1WceAUlw2LHar3JqSXU8y6tlY0XvOF026unpYSDc1icmnrKrSiQKtrcxg1
wrcMka4YPx3/ViqZHk01Ifw/GAoYJUaymTv2vYhqzAxHrG2YLlbeE2B7Tx4MzcPaWv+XuSodklAu
2ukEkjzfhCM/3EUDcabbvx56sgc4kQ/o/XwgnnE4xQfyeGjwBO3J5okS51JfJ+KDFYRVu50dQ3QJ
/B74vFCutPKwtAcyZgl+b0rfOvNxxLEJ9NJHe3h33oeJXgdyLhbyMa4jlyQGNtE4+880JlDIC1ol
FePbVq4gAd/aL7H4Y4CJuAJp91FFA6U2C9wp2TigkOottDdvLIzxXcb86es+/0w/hMZOzpYoHHc+
aGDDAC4gnNCwRAhjAuKgWOgRj3oKSw+XJvhZQf2xxQA8aZy01WdpGrBC3h/pKhB1zg2LaVYjTkxQ
sRPXdDqMQ4fMsQ7TSqfwMAT0++Ov00JWRh5Oa1LX36blXDxA+PeEY3WdIKQgl5fgBrUTXenTKZaB
HgWKJ+Py+UXRWQH84yD8MlHMe9GZtSozVWg0iUQ/Xlg/Jm+LyASwkabd2oWqTmNEte18h/Q6qjyJ
7qMjJ5tvjYyZHhtAFh2x0bq+5N6cFViwi68LPicK1WvYAXFAREMRvaxIZibsbXxxh1tY7V5aE3Wk
ZB72jyOKpH7ghHFDNFReINXtGLAFZSZYiRlr9ysuj9twBpr6LMmEzATWzYSS1mPeMN15p4x1tsAb
qml+jMuszG1eQzD4Pk87g/GkV9Yd2C2b1+ZLokcT+5+2OjNHALSqtOXsTKzzBt8nkhvou/bpxACL
+jggdM/bfprqBwnMvvVrRI5qDP7MU/Z8qA2Uk5B14yZvxtqbxJA5chW84S7S78csCjvgrk1pztYy
PANT+gmNX//mnxhLJ+u2Sq4PS8BkdpO49dDqAOGTuK3agrwtWZWu4kNwrpbJDabDXBFyxXVlcX86
xCuHvWntU0QUqsjUp2KGx5Q9+r7BalZ9cNz7a0uvXPe7XgbO8g7pT9HYzU6LmkypKDORcfYnwFfJ
z5y5WZydTTeEjobB4fchMhC1wzfKT7lfMVSV15yxPrC7x5pC42f/l8wH/c9Q6IUq0XsCml3w5pzV
1iZNDmKKOywAobMIg9W12rbX4jWZKU86FLASXz//kzjh8yZrTHU/wmFgxEAnc0/MPy/o3stxcq2n
4tANcf19iHoFDB/gxjLISGCgrdvX2aPsdlPB5EpqxrR7Bf2H3nZEPoLsIOatnVn9CJfMyifNAcTb
FFF49PCYKNvFNb1L+bgYwSLxRRsxwgF3azdO2+hE7ihSKbWS+AMHgjlK7SX8f2lFAIZWJObxzuxA
IH6FnKziOh0WO+qhPmbIZzZ0ZKnNYJ04QCBXKyoqhaK1+WyKtV7Ot/qaKFmYOsqB9YFQfoNNYs27
QaxCG3ip7Oe0ooXOF7U1vFsVKQ/RrUAFPP3gjyMLlmWXTbup0NMi9zbE0JAQ1z/HxeYXfE1TgqLd
lvP4L+KH+PJuhazwTRBiCRIjd9OuKAa4yYwhuQ+C17xeAtXQUnfIoZcmWp1fdyad9TWia7kvKgJ9
JuakOpVaYrhHaeyZ5AulS7lqZ7mXGGqsXTaAXfZ09yHduAv19nljf76Rpoxvy3IlSy8sr0LxfaaZ
YKiONLTprZqyscd9wzMBjiVM8sPtz9jOGIDR1JBUqt43UcBEvdHZGboed7ukSGJujHjKJPUVZ3/U
TaMiGPclasE6al6ZSBQpXd0AKt+YAZHmZQzp7C9JwwHJLLZgbYObwNdeJgt7Z4f7Gm9YUhXRf1rM
Za3Xc15iJtlyExuuzGZ6lf5jcy1a1A9DluRjoVGflNxYKCQx/uhQ3KX3NUREAz5fw4ug5fSAzauR
Lk1H84ODmGqm2ALBN3wB2Ju4sVJ8RQdXQVSOOhG7LeXaVEKlsqfL6fvxnNc94quOkCJ2TI9oPSr5
mGo4D5Fd7ygP8aUNuIICwCgcq5Qit5dyD1GomDiBpfzJzgSOk4SUEXWU7U2dtXBO9K443cO1ZKOV
RTrxT4bpuaNIgPqgCapf3UrTwsG5OClSglsu0SAUhEgqoXhee3K55L+LxSjMbFxdF52G0go2fBBv
SlGOT67vGUfo3Ma/gfQSANqp3UNZrwMxP4QrorCpr5sNxOzyTG89Bmipg0kCafavP67OB0EfVhUz
Fg/AvmzsJayKb+BPbygqHT8jyWLW2DjNMSlJUTurW11bjdWqfr+dzlAFrgmlB00euY5hDDg+Uo3e
sBG9KtM/2e3QaFFNq1HcDO8xcodHHjobvZS6bM/lsQ+zQRvZWagI3qjRcEpeQWXxREKPlf3hwMPa
u1JibXb70WXOcXZEaqQsQzUHcSatFbZO0yU24A7IMeCA4Fy2mIhqzOfn5OPtaQkjp/ugfWz/X1bJ
832gW70jLsHdnplGdnCmWaCtA7D2v1gVmlIYo/IjUixQn1UtMNANAOo02gPYMolPqjxHhhnYdYNt
VVpqZGxRPYiVV++kwIIHLohydNtGt70WLVJRLEDb2+Vd2og1+cFWNJDhneReIaZv84TLLs5Ce53/
qmxjs0H3kVgXOPjGziT95VycjN2wjTV+X8dU56ylD2NYZu3yPpZmtG9sjGutiTTRNAU526d00KAr
2fR3Tawgw9GiEkQWAWRIeIPq1sg40YLflPlRO7J+/X21FZNlEq4nzZx5MVCOuVCFbhHN6ajLlZzB
aso8MMF7cKf5R5rsdqfT6OUXXjoLh+oDa8DMARQbkbITkTP+WdE1csbwMtDNAQEHbnF1fNjZbPZo
5YdgY7P6iovIz3Lkm5JztCjDpkSrF74mcu/aA8zJmgBq78iLwrTb6vL7+wB35dy8uIEMS7R2maMD
VWuAqAAXcDoisIR+bswYiWqYjIF6u+JOxdJxgVwiFIrzrFubuS+m143Kph5wogms7EPwbSCLnP0l
vv3q/6P0rulgQ5a17uRhedAXY7psmJ0G8MzfyNHImxoeQ83NjTJHv1VUjfBNJEdx0A8ZgRsjfbju
Xx6J3FSZ96lJjuPSJREf8iTSeCLdgn8JBrjriQqgZpXEJ3BmjnYG8WrNU/YhXqSHSrcd9ZJsf1VD
8Vj4k7GlfIgbOO7ULtctaer94QLAPOzilSO0Mwj4cBRN8+9irS90ndLPLOX1m+wp3MEByFFM/iHl
XBtQM1RCRJ0tzS9SMDsTR6wiY/Ld2IvQoJhN8JX6cYNMm5QkcYlcw7o+zqyPR41snH0rQ/RJ9QK/
ZWrqaMtPVu1Rk2MscTY37BMbqSFBbTtKfAmbYxu0Wh2XW0mOOTedaKAVd6PvtQ1UBfCH/fKK0e50
o3FkYZB4On/A1s9ywzK6EXaP2Kluta5Umwk++SjARwCfYKHAOhvlJXT1tgCQZ0YurEp3L2+8/Ftk
wIAy6o9NHgzYXnh6HLsUHERgU2SLcr6gks5m3adipLBP79QIuFgOhP3dLJk5LNBWqYED8lycANAz
Fe6c5cdVlaZdUtSkOEyaRRhnOZeb+ernsJRFexf8zHGkrq4zcoomz4vxmJp0eLecalD369Oz/9Nl
Q3+yQnEQpPXWmee0PVQkBm3bfNH6vuSponKtvlxKzOHvqElDArfJlj8aDdWn9qw3HC3zste+MlCo
mmnTL20Qo1NZYRzocSsNVI3qhDMTzOO03xR21mFXwHg9Zc2XmpDuOhyV0Yy48UvdUB5MExhIwTE9
6nopfKBJ651ici7ky8ffEVgmnxXx9H8QDjIJDu/j9pFeolBfscLxMSd0FR3lYXUysfkEpoS9HuXp
EW387LfxQbaX8eW10a0le6mvOESIZrgGkoqObQ+IhrwAJ1CcF0vso+3F/BjgdE3flxBqgxw6fvgI
/tPTCV1hJXIZm/9d/L+YJt/jRBMqpKMFrRT0BpwIQRPV6QZz661/aYlDJ1yIHLu8E29D3XxWNevQ
4C96n2Ilk9C9wN5VuElAJDlVLrtlghI/NMp03bxtIWOX3uSpE5ShsHJROdr8aGdyE9OYhJHQJZBs
/Bz8lxpHwPrTVUttB3Trcq+8hqN0oBBMLkIR++69zSZmVOVsGtIg+7MthpkIa9VSDYuaSveQVL77
Deo8vBYxwDooaxmQzSa5FNcChoAu1SIB+revnfuWt1RhDNkFl05kCPZ3uG+vcBuPm8EV21sj44im
+WcnKJujj6CHXmnPQmh2d2wz84E2J3cE93dDEvUj86ki+4DX6QjHF9dGQ+dzyKugfuH9svA2zP80
fRgUo/XD24l8uq16vmQiAAQ7EpBYwqzivZoAgicYV9czR9WfPSbs2vZTTc4QmG7cZ58xQkeAVIu8
65/eQmhBzjqoP7eNZdbPH29HpMy49g6+0JTPyPMF1WoSpqvzh+xaVL1V3ja6YYl7Glyn+fYTa3wm
ztxvHtpDQoqa275GIK/wtpUk9H02xMskWHb++6Zz3ITrcxl5HWz+iY2H/wb0TMiUBVXiTy+ZvMsX
Ys8TkBYDAAgMqAGibesF5y+/2HzriIcy8sC3/glhYjXXC2uFLDRmqVBUXTCGu4UpbACdBQ7f29/G
LVTrdjN3sc7xgOul7y7HeoGq908jUD+7z4kLUp2PJWZWPcv4HhLs/GBcoOmvDBwYZOcQsb9EMQJm
oz8XeMWcPBTSAuJyVkUkChKwOirXa8mA7dPtNZVYv6ige85E3RuOVJuekW8fpXjeBhUQRZ/NVweL
NP+gJU5jTwzV8OlbOJF7DK3g5LJ+1e7jyEqooK65YQFeiwMkHy3R2CFmOJkbxH0stif0RIh4AdCR
lIC4AswrgHKoWhjAqKtUqT0q3/S+VMNOPlOqfIsLAYcLsStUY1xujo5eLdSaWRfb8ABpb+4df5ml
8KQ1g39rLftC4J52eqL5hq+aj1oj4+CW7kZEoFNpv8gTHm9/XTgaAH0aVYBjo3y6PczVFjybpEK3
m1ralJiagUan71XaVh6PhDXiVJ1unG3bqn8p0H37EIMz+rfOLKsrS3RYX8/2AfnTlcWb07EKMeDi
Pvm/NbJPi33xL22WP6K60FqtRsuw9BHoZyYg2Av29iVx64NuqAG6WH3UeysRfaY9yRsscsWxRDmK
o20YHhr1hIxAG1SoBP/YzZyCZmJXTO+SAmciVYFn5xXHMCoQ7KjmGMnYHQxipbZ+E/rDLBHDWVPe
8AT5blEtEkoUVidmNvhuuWDqT/RoKrHGVA3yzXgMNxG/EYHFQQOOewrjby9wSwVzC9N2+fyq54cx
aLvlb3zAUGAELvveeLPKsVVf4d1zvKgPybfU6yapbVSd9J8FYlqtYy+y8RpxkJe1KdP9KqphwBo0
bKrsV2tGWZrfvRjnJ92bC3J442H5SzQU21M/opExJXMwz+Ne1Se7zxl+uZwRTDD+NtdUlOgpV5Uf
UNdcpy1mlfchW8PxgKFD2ZKT6OG2ezZd8PedjpjKW4TeNcPMcDeKIZuLn598NxfZfHx+3P5TmNkp
IGoBFywiKxoTYoZWsDOLmhguQzJmPsTmBwZRV49yAH594XnD/BBDkG3qREOc9e1C5auVUJ4zszSI
1rx2LfPlLdjSIUGKqjKkRZD2rzqiMAJIn4JRu6iSyj3qakqyFF1cK5SMekS9bhdkwVPDa9wrhkyW
p02E2JynuubTzG5eFnnZszPndyibY6gejkEbmpUKP9h4404xYz0CZLHY7ooVKD23v2QW0YzoXw8U
GH+WFYfIBM7sBewRDHbQT6tDVR4Uk6OyFMIdGNodImC0u99GTsPDlsrGk27frzeXDn6dmJ/4FgmH
/8/jhTvNCUgzn7qTrxS32BBT3TaJ7t9Kb+cOtcLl1SfpThqyu1ajO23TitjMQZ4ZCHKQIBChHQ12
iPEEhMrb3oSXO085hjRL3gQVlWoX9OYcYhmI2eRcq9kIqAdkAEkdVoCxB+Y0sHqbyKFdqpKL/x2N
C92Sz5m2r74qSGlfnUrEwkaLUDGl5McqzOd85l/WAT4hKjMAI3gOC8rwy2YiykqpA0ATf0GX9HqH
4v3hf/wL6qAtEw5WjM+cKyBaeFS4EmbwrAScaaMk5MbYiWwUX5ABcusT3O7rDkn0of2fvW4jDI4m
3DLpIn6h82z7t3YmgM4No8RAKwI9WvrwIfQ+cfHyLNnAU1EROWOynuAy5VEMG2OszPkoj3I7dSeB
rI0BcSA2DDsEmiHUekGu+0LgZPKB/R6LMYZRmTH26/w7iOoZgboHPd4GjA+R/LxSH/0V01yyflGQ
+2AK1DOCtZVXEoNhbKlO8oQhhLuMd4X2gNDtncb8ve9IGlNW/XUh/h1hg8NfdLaJr/7yeoHzIl7q
ciKUxGh3rod8HiPrlVzR+8ktzK4pq7BVcRi2FYcVdQXp8eGLcahi4kxIMY35YOSN8yogvY7SCMg2
5F4LZeGMadFh1jbVgMroWngQVZFtQPJLkYPZs/zDWGSAdXQ9Tt6aAWKu5x3UwDYOg9gvrtbCKP5R
5KyYaU6V4svOrcea/rb2/9ksTeOwLz6gwsbZPDXqVMeScNPW2AC59Qz/sdDl10amqzWfaQza6GM8
vocVS2GubiyIfIS+2hDFEhTWCno1M13u5T4RuRZ/bdyYT/ZSbyG1dr7hqodQhdYKEb/9LMvkjMMx
yxQF6yNQGMn0/ICl3aIvTOzUFJFVKnYOmbfCiu7mYE/NXhQLzZ/Zf1zIXlkk2cbSGcCSz7IcoDL2
HOExLTe6Cuix9he25hO+q2XOf9UbkPyUSJJ2nVSUpYvrMMgkQXalRVM7pKeMM3V9IJlXEzPRYeen
KhtmIX3ooi/y8+H7R1HqW5zVAXvi7amqEh7X026KA6h7HWpLjoTK/6cHPjofw/Y7MajHrKD0rSAX
JuT79TAlE5Pb5jXLNZBm3zgvjU4eBAevHY4hNHWwOlEDzh3+WX2N8gk1JeTIAISaCA8JteOgY1pC
CI3Kx4cWT3gP2UIryjo31XF+qCTpLGnH9rsoaniVtNsD3iszsBDERJA77oFh5y2/4EQexALi5sMt
EfgsN3fW85UCjuaOIzNW0hBZGU2O1MoYQNasOOcPCheFZAEWpaS8wz53xXs8NqmKxkajHsOhZYcQ
Mwqk2aAOk7F33ICa8iv210rHiGFg3h8j9Jh5UGvVU5ncxoe+Ff7ugAucrbrnGOx5+5tAAdymXTic
tm8Fm1KysoXAH9W6ZTsiHOSUDRMUgIfYm7g6CozMbgrGt8XnaMC4CKi0x0sKWftRLBXDnk2qd8hH
dtfDo25EM6NyXF1V1EhmYBXe4gqElgxeLLONLprA645HPLtBCLgLJ6uJBpBT/gDw8/X1gRCb0iZ/
sp3zNTUiNAaEeYFl6EeQCEU0E4R09FnDKI0VJI0y0Ddh0YsjpEVR9hrPcvsne6H9hii2ZLf5SFha
DwaLylvE/nyPaUVsJfSd+qOHfrvy7AVvSjOw6x6vRdr/u8xTY406EdOYcq/RjCHqwVlB2xOLiam2
PqbAZEz4cBpTse3DQ8OGtpeLHS857npGqfZBc8E+vb0quTCiucvpfBt7vrJkM3TnypVRl7w46BAk
oVezVsxiaG8cL+SkHW5y6Bc2v2BV70XX+rlmUYngG04rng0Yr6Kq9J7TnP+oTJjSM8CZIWHN40RC
qkL/K/jzN9AqeyvCcdcMj5BM6ZomfdPkoVNHrCssf2UXiF3gkO+AR2qyQK2RXgKrk1Y2wugG6PQu
ry9KwSC/YwC46BmOKjy5/Ibyr+ZAcq+8ABIWcpOc+Ue1+BAlilTBc4GedsxDSDImw5y6UPoJ/LpV
+ZJP5x6OJvtpRJ+lt0VutN++NcGnBrWE+nw4aHfBUuRJeYQ3iJSmiv8NjkaSuhzDWp9s0UNcfleP
DyAl5Fi9S2zaBJnR7jZFzVyridr1RopWQavPntbXuTQFHnWKWe9e9zDFAHeV3e2KBbUKBmukvoaG
RPQ0+4DIeHZt+Dxr2ysKypGdLej+75fR0+r3X/Nad4notb/Epg2pi3le2OB33HDltEhdi9+ddYjh
wEIIDskDr9gOHg2aWMBhyTkY7q9z3J0tCvVW3liReHYE8IXkNuiiObit1TEELo0w1ybtI1kMBzDh
HFlWgaHaqEJO3D0WP15+tAa9m9tIaxxMtWkIpGrG3Hnd8AOBd3ZbkyUhwadHIhzWarySvbQBkY0+
Mwz6t53Iddz4F9MOdAbDetp95vQQN4jOujdEOqunmgb6ap5L7j4Hm2g4hfxrSfZxO1YhX7o91BTr
KosyUkUEnqx0v+6w5MbDf2uZkdp57TLKYP76ZMxZ01jUyg7YUm2IrnAPLfXJS/tlYX2DB4Io8rvO
M9fRyc+inD+Rw2kGXDsK5syC+LJXk/QziBVXoscmFtwuBISvu/DYdU6vJX4EARJdXtpFFhk2uSGp
RRD/B6m3dopHgYuzknMncvotHj8pHzrDl4gwNrNQddutEn/OtdD58jTatsUDMnNBd0fQL+jpbWaL
VLQendRKw7fvsxVmZ0ceXpeQBpxI10iJPrKWgWERbgI7m0wfgvEljmAiy5Tu5fheoECXAM1hXAbf
A8zHUUMLkPuF/ezWIrWyG/UbgTvDGGrp+mMKLEzG3/7HcdC3nfSFOgl+7CotFfC/6kpJ76FruGT3
bh+9xWjLFg1RS68TsNkWSiAzGGpTa+gu4P3PA5MtGKgtH+LdWyPJAidi3qTktfCYg6GYYtp1++vC
yrEELuQ/VHh9hVeAxTwb2GMMqi8QS3TRkzLKPadW3cQtcCHhEPMtZ6/S5AZP2g1AySASZeSFM65d
b8GwKp5OidQZ1oBi1V4MSEh18bC7ynJFPySwJsaieV+8JAXr+cjvRBsS6Vw59sFEU6VUx/OIR8I4
bNuRxfWnxvFpf4Q3OzN2t9D6ONLFHmve5piKAMitckHeXOgYb+dmpIccgS3iERmphRjXZZRR6rLP
j++mfMHmUK0e5Po4gOdSc9/ZdSmKmmafl08+NPgs3M3pj+yTs6s+tX9ijMl7ldBv7Ct5Iz0qgGeW
Tldfu98IrSxK4QoUZYrLbzYuP3Ku/edoImTOSzN6pSHj8oGu3/dAqaI46QmRgf+ezb3xfRaa+T0L
08Q2vbwoauPQ6QMrp9iV1BzxZ793YqqbFpFkE8aDTYtp0FW2gvav5/PgHqPenGQqmHA6Y925rFrU
iY35V9WMCsVXjRNt68RKsLiKFBazt0TQcYSlgC0gk1y7AYTzxROlPgMxZ7QnNM53q/iytwG/u1M/
ApfY3ziSluU1FDc/Jarqnh11UwOSKCANz14eya6hEfnQHmKYRFaoJiLpT8IZsAx/n8+wNibqPfZK
lkjUCicftNXgWgU8didPbeL2uA1whXA4Q6cPR4z32VVMwI+FCHBjVAXyVctbJ9uXAtkoqS5BrfG0
SHsenYu1lKahNuPn1ut+oYJzYsVYQ+A04wk7jpc5LrCieE9G5tiZHPqqm1CIz9Y+VjXIJe2MMwOF
Pog3RVxpdlsOdz/P8RVoPZbXIsGgD0soIwIpG895UiUUrvQ5vpmr8gtjhMaHC3Q9YlYUlc52OnAt
QTCJYEdWz6lWdyYRICA1w8TvUbdTtQIRvJhWIBT7LFoy0MslWES4FKGEpnefNtduxrkLXlC3dGBV
u++7gii9cLOEkcMHGfcDJwIx6dD1t5uyilkHheknid4JdYxVt2GWipWppaF0GTPzCTDUHQ6DvQXh
tdvnVuIumRospc6EWyvadw2cIhUoFAeUqL9oL/1b42Y6szjF4TrAjHLsXDVvgzwaoDRzh0U0euu+
+kBJ+1mor5P7yl5dsUNLGsUsvfugfEZmYeyBLgii5+626S7CSmPK2MKFe+oeq2219EV+wq6OXeOo
t6HkKwdNPaiScL6wowETBpCnvcpgUllFsFxDXkgUjFCTuNA0U2ZwGfVHSQXX4jP7KLv+MWR7YGmf
RSHNuq988T/EmLZ0Y7WWsAO1vlE+wmwi1j0pKO4m/fA2kque7bsDrZeKpDLHrzvTgk5+g4zYIgrN
PZ0kqxUtB2lKrwNBHjtWqIvOgznESn0mccphKm64lhDmdcTze6dAjPjk8Y506UmR3WnIfE2PvYQH
zO40MErO9KYPEqUgwdavbTm1l2nb5XJ73FGNNl1LQgqXDUbFQWF+kDUQYZW5AZM5uWTQPa55UadG
ng28Mnzys1z0XAhdUS1obEPMUbcqLe5EeHv87/Pq+NRH5bvhg0VytdTqxNSxZP6o54kc5YAD3A3l
PU0wPPhq+Zlz1x2s9a1fLyqHVHCNuW+I51e8hbKnzS4J6kmgK95johQrSDNCGb8zA8A9jitW7+0X
PkNssXZGHySmiUvkXBxgoqi5+Snk9PIRcqvlZJs/d0ipS7sN1buk76ow2APk51uT9xSjwukErAIt
RPoiB8ZRB/J1tM3drVglgL2hawfnB5R0kvswlN6HOAzjFKHdz3ld5LPyg+TIP3DbozAqqn+7ywM9
Gh0RXa7QOVbzCDHXhavL2Sx2HHNgbIyD9w0l9ssbDDwskIEjbbAOWbeSORKbwZKtc+Rpa9kLe5fg
4gHzTI1mfdm/HmexRkKB1vNXqGmWe3rSisSIz0uiAPH3ge9/IG1Tey0JFYW9UpZCIHYnP0Qi3IVA
G1QX7E+mb/OakIJUDvuT4qg6mL3MWVmiELgbgEFSgkc4MP2DVixkzD6372oXwJcvJBUkxbl5rZTx
9JBW/EZ/QWSy+uCaQWBRg4YNYvVFsXhImL+Il8HMA+a6xqqBbCv9fXf5rOuY02klIuuckPSFqsdM
mfzeTuQSOc+SOkcX32zfpxl7LTvEuxr8KqlEwIy2IMaBSSFLHUzdK1NcNiwpOsU2mGUGFN8yeEmU
H9CtPYZToyu0cyTPzRVVN02u5DECuS9/2N2U1vTRIsqyem8WdYzEwjNhP5CM1PhKJGwmRBGHhyMI
sEKlcQCtjVlsXk5STC27po+IYnkmHOgUyzQoUa0Y6V++1Qfr8OTpQuB8pp+/c0Ke+5Ony7WPAj8i
UpzqGEGfTP8Fn6GAE4tVjsHbj5lYqG4Z/pLzFLeubvTILTllEfDK3jIa3Jgbef3NGom/iIL7z2CW
3/LzRD5wzSSEEXoOakY8w8DM8EmYFejljgzV+V1riCeJKmuZ4jTJb9pYYo4NEztLd4ZszeBiPP0S
rQFHCFY03Z4/cwo+j17uYuALL2NDgklffE1zztp8xEJz8Baaf3hJ4CXzn2PIoC9dlY55pYtFU5wf
jYNvEvsSB/jXYZOX1heJyYEQXpPXI+vBwYrOEpnSzgdlJYWBl4Ol0oQPI6Uqy+bj1Q/YHV+EDIJ5
mYPLAXYB36WthPUoDButPClvKlGICzh3t3ifzJkLNHWekQld8142fBn8jTXBnitR6I3idXRC3oic
9Wu8TdHmFUU7iK2d/p2FuU+LBrXrvDMeKH1XnvRLqu3/4zqWoEcmYml7r89JxrQG9TZM9P1pdNbt
D1B4pAbHVXdA8jhb/qOFWI6QJoIZUgHJnSoqHr0xGhTGvo9KunhsZysyG9cprT820g+Bs+i8SWLl
wQJHNH8794jstKxLpf7GBcZlW4ogqrRIaV6WeaCalTb/L8egTCqd9v4gmwrOw6Rz1FWYHoNlU7SI
/9vNpX2golr0z0SUjU7IzNjwbcwlpOUB3TRlT1/qQb1D258l2oYIc5IrXlq2z+YpaBx3PISol2Ev
zpepbC1Vq6pzE5Na0S326w2KO8ozF2QpqirCDYsHeR0/UZxfrT6Z5LDAhjNWk4OMcz6yg3P3e8wL
1Na5Qqdy7XOPDdENix9mgQ/QII8ISuwqr3h4jNew4MmoyaSPLPI/N/V/VQ8rcb61mu6fOpfXy8z6
eBQcuBw+DBO4oMk+BL+WnwEGvouDVzcN2uX8qQ9G5ptVbL9pUKXoj0YgkXXa2z8whtrIXwdOdcyG
Fs8x7z1yLLek4qDFz3axBbqfMspDlIQOuZ0sZlNO4D+hXmfQSzKUkZWneEtYfVvIUT1jHCYKqAX6
ftXfJV5itVUqPrvyO4rWV+SuVaiGY8L7ODl0FjIkosnrKkLX0pgNGCTEXWnd5ZjrOqk7RVejSOAL
ArYBmPQm6DGPYCy6sCOChjf1Djwy9Vb+9o7cOwmUHhvHk/gY2kUL/EoIcMCurVAJ7xywkG2wxypw
6DHkLPsVTqOfqb0ARcoadpsPDygwvdGzJeN37Vsd3Ub1QbOY2YPw4XiwCYK0avix12orhnjpnLnp
sL5BGHInI1fg5Fi3WDsYadf0aHOhbcav+1TVfJdWOSzeISikC8jQQTDr4wJdh6KmJVFRgEEzuMNg
6hu9MxRMPUDh1EZS5tf51kuUpMfqPiBlLQe7WNwqkS9XX83o15dvJcmF8Fyrc579FDYn4Yq9l1Oh
vw7sYEROdugVtiHW1b1/RnoJl7JSyW9HH26x7qDt/wdxOpFVbmIcRbdUV5mHB5M7BKNeOOU74iZ5
5LaM+onGBARnVahhrOzoU+l/aoZGqc1Rh9fl8pBh6QP2E4Tv68p7gKtNqVKypTQd/sEfXcMLpjz5
MT7mFT+lAJvMidIB+bDNJP5RJNIM9iFns6VQUfU5H2Pgbpj+YPmCLmA+EWugUS2CnX2nrtke4382
bExjUl3LnhwMM4ukLgGuuvoLDdBekRU5SmgjRCR+/LUTtEcHAOaL1GicU+j5tAnUoqHvVeFYn7Ye
l8yGzaXPFvfo8LfR6Wt9awQeKMQlu+GMT49RwZKDjWzZ56xSl9/6PaDhAEAW53r4KhiF3ul/Khf2
9v4Gf2GRR9p0is+wTcJefAjn5seVhke7i+j3Z9NRJQ2X7Z5dZeFYDpUy9FdsH3GubiKNqulSr7Y4
ijEFj3sZ1jLVX2sPHLAXzK0hDjvXu4xTHsDCHnjTIP4+5glwM4Rpm99Wo5TX20ZTEjazslBnk26p
2AceNYtXQhVpLM1ikUEWCjcRFAI8EuQsFrjfc3NAQCuJmsNSFQd2hKaIkVYV3v9BRTyVSoQs0Pzc
UaJjO4hJA00nw93SUfDvK9qFHBjfeZA43IYaRwLqni4xo4Vt7/KUrNLZiXTi3jFP/hzFXocRvEGD
1UZfaFyMtvfexCojiqHUgkYCjJiIoXhhm7j4jSL0rJh0rzOCBc8aA/3CksjXV6QE27+diUjrRq3U
OvLrzdMA/eKv3r1Gm71AzmyH8gWTqDQ//gQv05p78HCE91ah1fuKJSDsAXHMbeUkdYLVclRtaZ4O
VlFLSDt51JuHyThl7A9mWRndAsgffeqA7vpW+ayXNlKLmXubEfLFKuuT8+4D76aQ1zQ/i0yef10c
Wb0RQYBQTLuucPCNtqrssTmIpoBozRqtoILhLgIA55Z0hSddSJnI8S1GLrH7WDYboYaKyhPawTtI
POz15ja2fRyEAqqZbxpP1f6MJEbqBEKrxO9W/0CytoSDRr3Q4bHu1vwgmv4XQ3s7r7znKZReymdX
r/JSO2/1lZLca2I+VoWBB6MwlIU7Z+UCPYdsLW0RhmHEBZwF1Yf8z716NMwH8L8B2fFSG/1mVHEZ
AUrjdyTKIhXcsuk0HZzOBXkkAhW4tSCarTDwTt9kEyr1qJOUZMAMU3coMAUXIXP+7pM0763anyIN
i8NYpLuhK5oKfRstnvwR6CgYhvIm/rfd3YEyFSAyZ8E7mnqlbA4NxrtFaGheDTURkvHV/TWPFif6
PeM7JkCiy+ZrOLoapSaK5GLK40Fff1yM7ZEu4SNOlbaTKaQL4btYk/RhOqRKkglJzj6uW2IrnRYP
GY6lf3HkD5Y4C8Xjufvvl2i9UiUHYJm2UeG0Ww17zk1rPHIYMoqiLpy0BQDUO/XAy5o3arhSUen0
GdYT9pxGibTLr86QY6oSkN3ca7prZnnQalL7cyLxNkyQaH45f8rOUf7EeDGXTSwEyT9cynUBA2C+
SWzEDkZUNzmhP/NTmlh7reH7Ka0UYKTkt3me5h83DhI09YY7iJmMhXSKbhXdo4XxFS4No1OXdZKn
mkUfQoO7U8DGVHzxKJ0776ffgxboOlStP7RCb9sjQIad7iqqfO8W1HI95KrpnXRfkweVD3a6LXal
xH4AccHvHuoZrH2C3Og1zUJAOVEtuExVWmewO8GCtKCbb56Q+QZt7aOp0ltXf8dLHhfVDPfU6kHb
atP6jpsdFdtFXWTxNvrOsebdG6sVH71EjLlgDpO20AzUYDiMcEOGuPQjsZnHw8yBNzX+zszT9+O+
F+6IMf1MWPDVVOhu8oxqdBswmtPouRrswXOhHIL3bzPlg91YjxdOPS0l7whZUOur+BOArd25F4AK
ocdFnXvWlxmZQA8naLv6WMEfprpCjy4HsOsTsV1HkaO6mIIiEwK+1FynoJoTGqFWIYi9Ou3iCLnW
N5f0qqpHopmqnT/6oPUpN3uElZHWFuC4zrHX7di7mjJof1yIrIKZXtz9gu54WBeCoxOEOsbxIT36
fZ8tNe4pYz5A912j9mu6sQBfU+W/YmU4lwesYTqiBbtzWgRxWrjOW/1Odzfh7IPCBt37kX3Ii9iv
U3qKDSlKER0Fy6OjewAlsnGj4+o6Dqv7rmuCBaF2fCGg7CzPLqz6oc39qmjQumClR/fQztz92tu+
8Yy/SoQwqJ6H2hGaUythtnJHTw24wXNM10VRlsstxHOlXClUquKAiulTtNWhE2tZPkJIY/EY2/K2
uBAcSHP8xUdiFBVIYi56EtXMwSzP3QTdFOvgsw8uE2Tl4RsRFmuFBBAmcfjJNr0yPaMVsvM3hHfR
H909qSmyAMzk2GY83Dzqv2+qJagESBHEM1h+1kGZFQDJlPbop7Vzs3CAeV/IWOsgquiuPxwfqJ9F
X3Ih2qkvaKy8aw6G6Fa7Md9o0XDsr7AzozlsA8iaHlgcu/CawNF9BwuSQBh1BbWX9iRbb7TvCAcc
asrldLe139U28iH8OaR3T9gVR7jU6jauI5Huaj10+HZ4gapHteLPIQh2FZzVY9YOoC11hViZXCsF
ujv46QF24C+WhlZz4vivGuv+1/Nq/0AIlVyR5Y0JfAPUoPJB25xzshowljvNPGGkmOhS+f+jdi1P
yR9JxhvsyEhwr05SjrmAUP1UmBPOE5UEVdN4T+z3MmUu03ez2yEsOdB8rUISLiPCGrRqFSp2bB5P
8jLNCsoei7+5llvkn2X/nS7t3A/i9x0OSsZ9kTVSfOznlsJBH4XRG+VnMx1vpGUprdo+OTqj4Cg2
jBsUWlZmNeSym8CGp9QbLRkWKARupVw5Mt1IJjuUyJ7TQJ0RRIGpo2Sbw+46DmzPW7p53/7CwIUS
I045RrNMVwk6bXPcpRIydxk3Xt+6ibNGShKnQo+hiMIjBBJoduduPPTGnsaCfpzB8ZK3wxHbbs6Z
mFduC/ZyurJUzAn2dY+BlISTKCnqVmcpEyRSUIrZtilb4iMHxyDBhJ7S6cDehnEnWad+/fZYZAJ+
YSsXww+orU1udqCadc7NZSkKO//I4eYBiGN9aGVWFa5waV9h7JWIBIPPiDieIXqUE8mtOfltgzkG
eeZwtioQV5bIMgVK3D0EjAa6fzuF8BwBMIstFXJyJzY8vNcxwfpn73bHcB2T2GB91h0jboWes3rJ
OEaXAu1pU6RPbZz85Zcj31q+3OecgKVWLcAVd0hX97ltDlKTKk7Ehxb/2vB2Slj2w1A63CO+qn2G
BruxWs1ahXH5SdOdC0IluzdbDoEzmh+OF5pqmZleYJmX1VyPvaphCl19t1GTchstAqsC7gCONa18
Tbnuu5Bcz8zB/tBHFjTIUx34EQjwNbY4xj2KsF08wDEQ3ZS0/mWXevW8u7npiAate+obVtY1qyFx
YBY9yniNMA8qyIc5IetgO2bvxDJH+X0ve/+5rSHHOr0O/p8SpPkgvwP71P8qMXSaM3NISZooq8t5
82Q8ggXd6cMgYlGC0wscligEF2t7i8Soii5f3UW+diRG3G1DmbcH6dCSpSYFhYxzwTt0RWLswOO6
rO29/zfukjE66Bv8xD6UOjNps6YvkMuYQqHz4AsTzZ8fJ2E5qiajXc71MT1Hu7RbYvv/bDL6bTqM
aMUCmCCRez2++/NFFVaNoQyRS2fXJtJGBA60xH1yHo9xQgnanRwNQvcEs/fvROcM9re2xCDb4GZu
T42JJlwtNOL085kBQW6E8xEHZvkiPAZLwakL6Uzc/EKr06GuYaa0BPNn5jbFcmIXbouQ6MBA2fA+
iwtB8Zg1lrZ47gqrvzqG0WbyPO2C4oxUsUzonb9mJMGzYBNBbI2ZaZys9oiJpfHsMZyfHhhFbEd/
wg9zmRBKXr7nFwkk5wK027axYOFtj5lpDRL0DLjSTYBBPwfE9ARWdG7887W07p2kCh5RaKM4vCj+
VlAI+oPV1d5hwoUX55pqd3TfFvuwl74LwOll1kVClDEzcEkZ8u/AU3SgOlIE8OtTt2KEdqWI52Ij
0sn5SE36fCz+GYCDmHPRaCgJcp3RcW0uLfLd7Pl4qteiqtlPJyJXdvg6l934oG0Oc2K5EmrHXjOX
ccHjuOdQLhkqp6qcErGPJs4OCSU8YP728TlvoTu7eK+YhjGl+BxOhFTWAsM5B/TlJTu9yzd3Ag8r
OGx2Gl4dJ2YdX+h6M+jsQRt6s8dsXiduNRSbDat16kVCX7Phl3d9YG0R3n1cpAuZOCR44eQqETm5
5YLBoV4VbwL1RPorb4Yzs83Ev+xKd8AH12SJvF1J/1LCvP83t6lUXQe681Xmr0dItR/bJb6j0lOv
hDKw+bsih2YUyiF0AzTzRBfzL0SIl383EFJ9qFCE/dGpBYDrL4NhXYye3ns2z7cqu/fkXdquBrWu
kUK93hoXeVnUC3P3IPVU2SSmF+apNGJf0AFocgzL3/N1ablLUKKBFy3FqqiBAJRBJn3zRpuzjPoV
SVigvpPe4oE7aiJDZayHQHoE+7PUVgk6Gg5ooEBjmeh6AhUSMY1G80rV9Fau5zt40J8ZWFC2UZJj
1h/s2QFp+kEU5rrFZKXpnwenM3IQ+4MB6kM7CwItECB2GeyrDaPwKh5hWcUihXhvZufepBucQT36
sGxp+yyfI8mVYPCuURn3c3SWT/OdZMOka/fuo6hK8ZWpqqFfNi3jSrD5TIS5vOA4pv6d75c0bdNt
hXeZL7Pczgir3bSRFDyY4H7FJZTokHPnDo7Sup4ge6xhSU4OCJsHijz6o02vxexBHGcX2kWt3KSI
bn3i/TfPQDaFSwQx5Gtc3sSf6UpqnMZd+7ju6lD/7wizr0+ZiG65Ul/v6aIF8WpEq/yVYkx1O2ZK
UPo29v2FpwLx9Mzupw6Z07h0Y4ixKYPAPDn1CNLFSiqLZ3Dm7CXHudAlMW3Sy4axsM9kTkxU8hbc
fFKmgMNKPeqtBexKbNO97dm95Ru/v3/pYv1qMZlWOR5lraGGs7EgS/o407Lu1Y0ZkdwNwrO+c3xl
ShD8kpuvTXeXc/fDJzPoB5bv5Z7shw3Ymf8a9MVulVaDL8PwxdX9dZ60rq4Aju8tHH8kgHR7gaAL
bHY4xhk3PKhWddwa/2amWV0pZE5odc2D+EnY4IC/SkQBOgHFRnKfkTa7WAztHoNjU9UBQMyFMM34
k/Wumjg1djCUbm3h8nz0TctG9RGquGqJzNnSCtG/i/69BlnyGoUVoGOavSVa25WnOtZ6i7aC0pyB
vC5ZYEQCzUCiuQe1p2UrfqC/QOieysOqTYN5y4dP6FTSbsbo7qFrfYHNBeVLWJgqcs10uXQOcazT
72sx/4RC4KDzC9pZ+mxSImkAAYEuB9Fp9qeKeY7fUHnSAuteJwYqpfqSqPeCV1+cR7/XU4mVf6B7
0uaRZgsSyxmWi3yvjFwjtk7MiWUeg2RZKZPi4q/KxrTd8vtKPvPedFuCGYK1UIo1mrAHxLeLHXJ/
TQMWNLpN3ZzpMqVnUycQ27xCLoDJllyJrUXU24lddzsmMqSSIF8TpKgsNOkjy18n8ipCQeFTU/aJ
+pIX+KH8YjcIvfZccjCA6djMNeNsMfSwlfZ/KobE5+gUyHhSoccKGaQTTYuvn5TqjlpIo3WnWO93
9Tzhmu1rN06LaZ0ytYhkv3l7KfDZnLXfR2Kn7mTD6EIOk3wTwlRrh9Hxp0bv3YNrU9Jo1pv2g0ZL
gp5VREWpv01gz074NmQv9z1G860yq8sSiMAZDmw4FYWAfwCCZJee5yQaSwFWvbaEV9rlYP1k2Mfa
qbFF2tJiCufdpk+4TBnOh/kNmtP+lcd4ziNeRXsemQqq8nbH/cY7248yYcjO6JAiOtGw8WeaWHSI
uLfa7I2q2OhULr7nwXikmbGHoTe9Hk7gBT5UHWuWGnqSwOGmPvbtmtdZoOoRYuAvrOpeCPkb/Lhe
OPJwv88BZWgZsRbYk0tiHJLk7t2qj1z4X/sutO+l2jIsJzi+37mn5lfYtsG2gDfmQh0EKrduJXZk
j1n0I5J1uSoAUqMW9QOvqHnCKYatQQHSbyrp9DG4YAHxQXtwNgw8a2my2yyq83ktZvWfCByiUPui
yGfL3QjVlcRHljd8E5UGoWSqjiuq8rVWtGIcT+qneTESPzXf7QiCetdK0r6bJnpGX45Z092sB8wP
KkkV7gPzTM2S5gqqjwX+ChZHcotTcsuF7t7F3flMaUI+o7WcZHcvw+BMkqU0ZK/e1i97tOt10XVY
VIw5RTOhYbJC1IJDZIp5B3E6HJeBHXOnRQ4YSjSItwfh/R9p2115Kvj2hT/KGEpM2CLhYPlfMb6g
pbURtRvpiaQJqTR6yTfOqNzz3S2oNFiIrsTJbthHANYBsfBovVb9Pnxu86aqleUhd1zZipbfQ6y0
HA2aVGVwMIBvdB4Ll3Y6Iy5heySgRIgWOQgo0YUY5mBLaoml2AsYqLsI27SbAkYT+6s7znuk1Kvx
vm2EeIip1WycwIOY/uWpex7WzZpBBIMl2DjPsnmUh79XmGRPP2Rn+NjVQ7n99yZc62C8EHimojM+
3fe5OAE8vkB8o144H0Ql7TxI37y3gGTM48AyI5RRWyaJQFDHRD+oSy7ngGWkyZFfsUqM8JfSn20S
CrTaQRIm/YNyOsf5HWna+ooogLnIjac/cuVy0gZgZoKOyeWPcOxws5P+nKhFQopSge7/jbxIU0CT
VpwZkcelZluGusHu7sQrrxQvlTpbDPy/813w9UnuZsGB/tjwvU52hwTggOXVINqU/iISsLshhXz7
Oqs5bjAM1q1CB0frNSVLqVznJlDeZT1JfMRCK0Z26X2vNpIVtWyE5ioXwHda6ouDxlM97L6SvL3Z
69ID5stmF5t4VdZbiFcMJUwq5Jne0+j9dW/dK8/s10C090HQ4r7ZtC4nkIuK6Lr3TTfGV3eevXe/
q/aPQrsP3ajeuuPEweX8xRyIGHuIMhh97CKifWj5psXUvzQtAUyJEi+yqrCqcAauVpJ29HZ2HT+t
RJvVyTpKlkR3nBufBzQv//+NfYEQ8FOcUh/UR+TGiVp7CyOQSG0uwcL6/ZoOh8e11Ed7I66KfwwG
2AfJSg4LgTeFe2PdcirvFUvtPzThL8XckboBV6c4u2vTNIpr/Q815shVLprQE2/Epdg8TTYMYj/b
WOD8qz8VjaDkPRTZlMj5ioRU6jJouVd6OYsi5m6Pf8ezDcKgHLE0ucFEf0C8JmEeeCNFX1HBUV1o
thhO9rY7ZHDgEgrSGHxYPWHeKj8RDv96QbhAsnyoOMXglTQvVCKKOfGiJZCkIcDGMSa+K2kEekce
MiReFaelPRIWvJMce26ItyxkoeQydh2I4VNPAb3Fbkg0aA0CPsIPqshx8W0Pyk7ra577yvoiBWa3
jk2TiVv7B9f26YDbZXVvXTkgjAlRnstFUYgL7jKtCpc1UpaXlchyDcQxOo1sYtpUd8FR9pTQ6+GM
iavZyiNcCHesIWvbZH/IEv/VPvz+tJBMF13bh8QApU1nsiqRY1tz7iBGJcCIG4daxe8d78Labsja
GybD0hKlVWKtbRyV07uRf8k96dzgoxfTd15zhmhU+37a89xuBovOqnik5DgZvaA1cOlDSzA/2kat
Idvp3VVXhh79Ot9K6pcwaxMalXypYiWXH1vZWyHvKlbbM/ELqHqGEIWSzyWeC63nxhJXea5jni/8
6y3yLWm1Z36broJxuWnHa1ia6WhivwfcuhfQztKliuyR1MemE5j8HojHOuvKqpdQt4GbAoVPRqFi
AGnPcvPDOaMSuvbuhOf+1CPz/JGf7YHPbnvKzyL0DLzsskQFs4PTnUfb++UjerjYDv7FnO9Tj0/a
P5Pe5hO2oo3EjxjTu2b1cg5eVQw7A48UxtURVpgyIgB78cvx9g4rJriKM+I9bMhIZ151Au1JhWC7
hzC5NR9zmV6OLb+kv4BQNJ5gmUjE3OykO1RbEEl5CNT9vpmruSrryq6owWvBdj8jhgckputi/qmE
xlNPb0IiN49naeLxQBLuR+iRr9Sbt1myR+4o6CiCsLQ6LINUaKQ82knB0JGn2LLEjShf/w0BlZLT
sD5d9v/EXKyzJ398Y8tBsE/hs7YhMu5VKfBTUaK2XkbFupyf9Xspdmglh+mCBGryK06WGNXIebV/
pwntBKZ6FNe3YPrRHov8DjRd4yilqxfPqFQx/rn5x8yZoGwxsKhdaBVTHLWJj/sy8+w6QPmVK8Yv
5ikuHvDbxRXN+Y4QgCUpagKzrmaPQL+KidoQBdND1MKEkqId7kw36CoeTmFUbWjDbV7WGy2psGOw
VBvnzpttU9SzGO1+qsY/Py1VRWq1PTf4XFXbmO9YtIgHP5RgDBqSMg4qTV6inPxKUulvE7KB/e2L
ZZb3+DRV67LtYBnk7M1fpJ29HkiE21B6cxvfAoeoMCHmS3QoLYc4fpYgDKogRpuM9IJrOOyLX+mh
0xcrt/OFzXg1rV20heXH40VFZEocC4eiQvI5IuRkvrD1nBJOqWDjQ/s/AveSKUIgCcoVavGuILs2
MQPa4WWILgFGzSLy5HWzB9iBgFhYQryyx6J5MhH9FE3nqLnyWUzFIW6T8p1GEqmU4jsOSIPbHfmB
UbjxaWrDNr3heJMW+qQMVsFT5Yhp1WskeCH79kma31o8kmnClepHlakvdnm/r7n4IYJc33cnTuwU
ckDa2zWGhH3RP61n3sWkTZTo8fNuQNvkpO8wNCXRGD3j9OIaX2mGUsPUoVTIBIvgvmuoXxs7fZKQ
C2+Eg73em6J9GFDa0h9tG88E0rns1/43qdC0QuLjXtOhW0H8JdfRKZ/qooSAQYl8zq4or+urmHp1
gqTuqN2xhauQ/JInCY4dDiYcx9Fa8jy2xCD7Dl6hjvJh+gFGCpsylJpWFkFSKUnK4OMrh5n393wE
eF/NLDYmw1TSet+ECaJq1OKsSyZhSJOyS30n2GFp0C3y9DXyai9ZtoFLg098Gg6kPtM5b8wzcy3p
/08saC6KQZH5n+rz4enDhDQ5ijxeV4Qvbu5ZEdhiOLEffIev4MBMDfZ9H5n63SZ6FA8cjTKJunU9
Ukwi/v4GdBKtYlmQON3Ba5+XsM0KeZdjyS+2bLBqjQkj+3F0U5WPjiEkM7a+F5qDGK0yiV/pvrpU
RP66WAeEP4R0DvULbuvM6KctoEiz9ccPKudgzuWLPpW9OX44ZBNx46ihjgKFfYPUn6iD1XvwICS4
XUVtDF8kzOE8VdfAafpUa1UHKheDVVIEGZfv7ofUtWhWT0ZVD+U4fUXkYQNDNg97IZSyzZ1iS6wZ
QWFrxBDmXsbwFlfYK1e5Lu8X80t+03nQmqLNkt9Ge00izleFulmLH1i1oVQLkfMEaafobGvH2wLy
VBWP6Kxj3wkvgHd2mEhn9nLEGul/HZb6zzUprclSqDih0ZtQ8llvsOLmk5s4dy5sRbgSKnLNRSYa
ZXZT1lQsO71JH7DNNhkC40t5OP0+5LWoJkXJjVeTrkGK+/hgGDIMtaZ5XvixuEApXwT04fMarzEM
JA+N6c5/jw9droP33lTfO4fBcMtrnzzRbq0LWEX1api3BtHclg+mnxnwsdB2h5djJn+pUBGS6VST
muaJQDjVlV1LCbN0//1TxYocrQCNxr30iH8PIhVg/c5OLcaCveDTjqfho5YigFFt/PF1lrHrHKg/
qgJRSMwStQ25eGN5spYhSL6Xa3P1vZSepsEo8KZQZ4aKOkR0sK+GFR6rldqb1gnFVF7gtqFJaYyC
I29GIxt9uswaEL/lK5B8vJeoy3UszgQ1/Q7ruLsMs5e6WHfIDGbnKYeTZAmAjgXpJA9U1a89ZbMe
FJAtGWBV5wukrQuQ7AzDfakHVcjrAl2SbTW9oewphpv5zET48O6ZTu8dxsr0xMw6tSERtnCX02BM
XeKrzB7XujIdSKhPSvcP8PTqtXRz+VvTTvtqmB/AW1qx08wm8l3RNRTCgiyhE8ZSSuRPjexTijLP
JTpuFPj0Ud+mCXEVayG+wLUkFyHe0D6Upkcv11GYEufjE0fRPoFMkwhlH8twGKCf4e4kBcIabgGu
MceUORMBbjNpoACJtuSBMfjCDNzTHiWIeewnXDRp+DzuaT5J/WXYTLoQp/zzTSkDCZ9lczQPr5k5
2NUv+5+09JU+0108qELdo9KX+VeIJ1HfE5LT/J+G7Uoj+Tl2vtL4dm9oJY6xpk6lkbXG6CASoINI
yuQ0zov13cPTJ4ZXLi+CVgW6nlOTXZz1nERGXqzkAHBkeOGir/2Juv/NCJR0ueNmOac5lqWb8Lwn
tgzl6qOiOqKE546ZSuB4pKjvNOmcjJFJ+ewomxinuwVuWdK3pLHthsMh1gh96MvPzBjqFtb7OJc8
YO9okTTWwHRgW2TURUDSJzvXbVvp2fa5mQcYbkvczNA5wKkPP2l9EYqb2qBUWlT/LR2XU2zDGidV
enUKmBYkTYkKKGGjInIIYSASvy1ebgjj6ibtIidHuie0gIgYstZ0pybuFwKIF0rKLkhKHr3fJE3Y
l3u//R1qnhj7eHOn9Jv4UVBRAkzt/YBr5HPrq31BgS/Iv1UGieCIfxZfttRF5UFLEFYa5PWzyvk3
mpAFi8DbbIxL8SkOMHASA7L0K/yilcAC4UxzvFg5rzfewWdFt93Mf0qJ8CKvGm/CTfaGrGTUgesw
UwzJDe7fiOGP6SkQDe0YHDki/FfX3b0Fl3Cw7R3pwPpvXmZgBYoAJNhHpB+QRQCyawJa1zA3FlSA
xHIfZ0M5YiTZlB9Uial1wLJOhT5wuY5Y9cKg5T/O/6KaLW9UWQR1FdzpIBQDJjlrtOmNh8CvSrcU
NqcUdq24J3skg4VmWIKaZjQzwVTgw49zBUBZ8UoB8Be9ry0RHb6E1KDUrIiwli38jC1S03mE8b8a
NS5KP7lz/DHdsGfkSigjLlcrwCmUTV4YIZLHfRhQENWG/+/41ZodW+gFFAKf+qLbdf0BKQ/fOtZW
GI87Za9a/3Zs7VD121qkG2oMjQ1QqO0xedGAtXqw/u4wlu4Bw/ZAi1TEHHqxs6JpjAMUMuc7qvus
3gKDXSY6b1PNO2o1WbakIJeEbN/MBhRxsOOauq/RjcbrBisNaXolCGTW6CUttS7K8sGd4yQjnXJD
dnGg15nh4kuyzt3X//3WAFkmB8rZ91fH8sYAzEh65QpxQFPRY6OOK9xsnjLORl9rc04HhHC6Z2GA
kutx4Xo7zegGmS9b5td202Tr9CT4BytlxV2QC0XFANxbxHrAhTl7KDmALwkcpWpW3MiuYyxwieW/
wn5tSZHVADNKB9PpzEVIKQRkGT5Wr9kSeqqJniynPWT+J4mCmkSC5+yykzWGmnqOPJLkAQd5O/1x
xyRnuh3L/CU/8RiDJakpGZOcc5I5SqlNTUwhounQJclP8tBqq3pU3B9S2jJgPFvrA+43Iy+yn7Dc
CNMjNIvX+FpQzds4C2RokIqY5vhUmTDbqiqXfZJPV5yoZmBH03Tt1GRBMqufWPjmuVmCmNhp2VdW
jLtUpbu9Tjyh5G8AO3W0dvvjUcYNYuEH48lr1ShkExDmmlvNzwDT50zcYWDDjYHjtXrdKayK1nza
lIWtA+FcEuS5aRmtfPaoMKcKvZCGRlOUNr/EFTTzw1197hvSekq3w3IcR92zUE5qkaVIbFKihvsU
DULwC0EvJR8Du/QufMnKJgrrXFw19J91A5EJpsen/iBwFBXy+PY/zjom7grWNVAjaI+cGqOW5N32
us+nAwV20dxcW8WDLpTRNZmPydcgveh/TQothOgw1tdRLL7/TjtqX/1A1n/PaM7SDzjfvYx5Cp8S
CugnSMYhXeG1rp4yz1uRp4PAqHFQG2Jaqf42qRp2HDVonaSG1Fc6rZUX1O9gTnXWQ2Gl4Y8Ksp8V
dWMswcvBjKuzM/7zfDu25rlf4AMTeF7jvs3f8OG56tRC+qAtWeZrVvzN12nk7mGYwwkO5l5ONdre
uh/8emkLDzo+lx2REkQv9EE8tqdSM1ZUHcqMLJb/Jh0EgdNBqT/aRNXzccsOmhpxdgDRGeYsYs45
Mm7cZi7FoDzN6vZOKBefiC3AX5XY4Qh2xYuquLfsGVDfyc/8MjpTDNIVt38iuN8oWGki3kZaidO5
xEHf1f+uRlRAPG2lmRj/7DGvf4z/MZN80yBJVbTBRrOTasj/F4L08KlFus+VJz9z56378/CAqyJR
XcZoq+HPDKgto9VPhd5j2eErVl86yh9OFF9SKAa4Hp/gTkgP7Slaq7xFNslkCNwDxVpML3W2nSec
IkAQP5shWFsP/3IG81NrhMxQgn6LXE1DlcnLgpKrLKwe+Qfa4YWyVcjaB8WY0l1IQmHxHcvS5BCK
/4L/dNF1i5IAxLNDtqdHXL7UnMOq/Y2YxkXa3LlC6jyIJyc/ytU8kK5GcfqxpoDHOA30o9dHfOf3
DwV0NBVANskhAz31a8s4C0zP0etQvQ+hopujH+Cer7KV/hPzyojCMX7abR9j96uOtIPfbNCEZaGn
/n2rXIQDXOD5YLHuh5X39bPyH6KA7W1Zd1SHHAwwuAkFWiiqNtdHhfkSZlSLNYXTbDcdujARLyhs
ICzH+k3N1HeCD84Ht9MjVW2DjJpGypP9L9zqNCtqgf7aO7sUfva4hmD1IKoyrbDiUGFDnoyMk23d
mOh1epOtRVngRQh1LoQQJrJvonQ3jZxxfPvsSROnNX6oLzlBd4o3m2QbA3X8E5ssEYnSVXN4FodX
u4w/3uAFinz2RwSqwCBm4g5lNQLs2pXMcAa0d+AsTEhitQtPREOXKcfo5frmTTz3q2ZBO6T0HjXZ
scPhZ/FJET7U81rXmKIp0EB+xX6S0hY3fQLA6jCTf4NuLty1d/tPCsLwcwtpGxgV7C93cLku1ghs
xgQwIwS4dBUUkergfBG6llxSGFE70R6rpJk6iL3pvyAp9sRxGy9GEKva6FTIUXTQ113G7BwlQ37G
7wvCR3k3rpRx+yFXEGR1aURSo0HCD2DP61WvK367QsHXHB0s6Q5cexWggVFr+/xruClUGI+cjfBX
/OTDGJ1HXLLPQK/QqvHdiGLxaJ/BZamPJp7UBWLug3zcLEd9CVPT61AIV+XIxMlgucskIYX0o5gH
LE8qGbxxg0Ba1zv9TJZ1vKP693mSFLG6kPjBjDByhs0q/eXA8bUnRsGD3sXaiS5NYtWGb1xQ/6Zi
02ia03NNIgVKisxx+QT2jDkhGLQHzAdCkNP1F3Ig1iXknAsofqNQLji3YI51bO35kvIIdlChdCG3
EG0R92DPYf8dKrbTYd5GrpWZqUTMcTptDNsDJBueSSMUYUr9qNrjABIJztHXRS7OXL6LsZXgh2UQ
9k8/IpxounCO9sMtGAQ19Tp5bmXg+DFagmvVjS7abdDr0pgPtb3Spx7dGmdjt1zfwwKAXDE4RN+r
hkBRrmbzOuI0pqkLNaPW/bJv5vmSUXqho+8QruF5IC9nNOPY9wr9W5+xU8dXXI1RAQm4M0ss3t5G
CyeKfv7a4T/brsYmgG8ogwrZC/rfPEisbGCHC0Cg2DQ9jt8JjCkXtJOlk0QGlEt7+xQcWwTpqOR4
mAk1XW94ou7nS6jzuSpMC+iHr8ezCEb1qwU/5YRWiVcQ0i2LDdYWxacW+4i3wR5G5RZ/ZikZ58mS
4YYP/EGIA3qi+Oh8F6EZDNzch/xIX1hj88KQIcrcEX11h2TkR6MI5IIPv/WeL/XcmLtNfIJkOwKT
ke0tJv5GPePgwYvg8kEjabGYWcfPVy4wA0sRZWAFbrXIcSxhhkG8WcigIFN1qqq6wZ4oYEu9T43x
U4e5LY0EBGofIWMWjzWr6UoaJ94t9oZTfZWaSCr4qRKaAwj67/JUkM+cS0gnG8UuaceKt++W0ogK
04XgHM7b2YezgK7L0uxyg/tJ9Uve0jiPDwF95LKsom6Ds6reWF08aw1vAwx4QHB1CPiVf++Cwsza
c9DZt0dIcaUeVKpru0wOgYtVgnwMjmPOu8Ht8w+GZjxuswHRbMv97HxCaVS+CJrQaI0hL+G0c3/d
Hb/lo9vVTHofrUKNXIMWNXcFG8RUSzEKxhmSHtl1ShuAs1L7mFaYPVJ+VjQudzHiy33VHHXZpQnG
rQMmw07STFhdAHHD07ZY3bTdmXXtHgkU9d4h3aSytMmMJba6oQg1cUWq7o9yvogTqx+eUGli4tSN
RUbYTjcLHSfIjOKPgS7QC2zYzbyausCnvI1bJTz5W1YdR5Df3N+Tw4zggF/ZcIkMdRWafjUSpWOW
VvcJLHPewq0aSrz61Mxuxkrgs9yjSfgwQJRPd2GkKF1RvP2qfT1htz37OjU6IaYPvZ0M5v7qaU6l
K/E1nY+c+F5J3lUQ/3Jr3363eWtKMqu+6zUYVhJQHXwX/UIowM9MdZldPvcOhvUNJ9nkJ5d0kXXM
xTtuSUgVCv3v8LIL4ca5f1D3JkCVEuaVXHSJHHdaEMN0YO5zF/0ISYoEANPlBT0atFzPtEmUI3rH
kHWbaEu0+h2mwQ6PCu48RhoT0rww8th+VbiCv1COF6biBnST5dtFexza6a+BaNrAB9wRWDrLD5cQ
yw6bn9X8YUIFV5IF9qFEvh21MY4pvZ0Vu3r4eHBS2aLrELOAVdFQbpvP0nJt2qORU5g/LhEENKbK
OaIy+/ygYl0H8w4RXCUnk/oyBXfYfo6msMDTFK68sNSoLVtIY3AVZvvHWsCDaCmCvhqSrjMhYi3U
xZd1Dckuf3/1OcL2/RknMLRLgC927LaBYIEVNYGMrtlXS3gp0Fpc5S5Pm5b3Q3dPEG3VpkY8eIwZ
uk4TH4NrzRl64sCtg/NvuV/FYtJfz0tLJuNd+Yd6XjmJDEO6TEOwsXS4EWkjf125hBkFxRMHn6x0
/cdmBCuTsz0jZfhR+8YDHOVKrM0Emc6bSDqc7JxCPGA3JHHKPSgoHzvrxDReeoAn7lS6Q3zsNw4+
gpmGrl2IqepyXpIidK+Drs/e3RLynsA5qYCfivmEW4IDB/ASNAw3w8eg5GC9OoRPvhi03Wx7sz33
EBoLo/zlRJF17eX4P4lc9sMMkTkk0HR5lNcp9UgsI7ScIG8AKUMO9eF90DG/fwUj0WrfQbE2Tt7G
O1a8//40o0PbLYdjVE/NLV6D8Zi1774kTRLO/z5RPkKgF60dlCT8rCRzbepm0+mN7ekDkdNDSQxd
W0U/4sRmArAVbe9cKXAnz/12nNbqYmHWg5izAfoxNsq86W4bxT4MqypUO2b/mrK+8F3ndenZqQ4e
K/uXzHc2BJSjjGHFCgw7taCcs0hTKLRgPeVfdacqnGs75sx6OxC7ZNbeMdoiuPKhg+zGopZ5lNOO
obmjr7TyZZPbP5mdG7/ieVIJPcrosSXQ5He7BKUxOL4xQEjA/29rIxvdpUP8I20bP7CRVWdDco6Q
JN1OZxKvY/gLPawNFaVPQgTAjVEDsi/w1eDOOsrDXPpqu4/+vIIhw4iHhL6awrcUe4ZP3OVC4K0e
QG3cY+13nskA08LqrXWjyMoIgPeqXtxkbNVqnA9bszwLPnlmPfBcUcPrmy1n0BVsp8MlQkoeHjJN
A7oImOEwVfr0QZ4sv7816KkXyU3Wv5IexbMVxovruA1cAiXoPZ8fq46j7XP+Kyh1UhGSoCxycMUV
ZjhPnrgz4wp+9j86Wsg7/HRPnIAA0YiU7DvbRssXnvtjt3Ryxtx4vg74lY2PYpY9/Ha3Td7Ud0qe
Y4M739TA7WY7pJJZKe6LqSAIUzFHo6EQ0SQhY/MtQjm4KcqUdE0SxFDjcjd4T95FPYAttItC7jqe
6LRF1BtFrQ7YGSGMPVAiEVxsNLcrs/+eIT6rmf9YFv5X7XLP0nMlq2iZ5/XpdfjCQSmde8vnkP9v
qQU2KDkRPqzvwvWtNHcgTmaPLcNUgYpJSMZT1nsLLwXnlClH5irtN3CARWGOYO+72StrYe/Tx5vS
A9vkhCMMn+pmmq05CbGgfZV3J+4rNeKEQQAERZVEDMb5cAsGSrN6tPdrCEC5zTVJaSH14hl3OkG9
glx5Xa77qxF7exH9pVTfc6S0L0Dl9JiY04Ewlzk0JnpRZnBTDpRnKZQIBPjqkId0fIegxh4VpZHW
DnbSARBy9Rgosh1frFQ3+ryTsRxFwf6W8d58B5UH2e0C1ubbzZvvxdJ5Q8k+WPzEaapUbnl8diT5
/oSOA2ZEyucUWFmeH/RM+YZu1Sb+SZMZjfT4XlF3mzEX15nqv9osfyrzXx1z2A1iqH2QXBlGovxM
Iafs/CVdFR26voa+vBNItyZOvUlmU2fG2JL0ysLXmiNS9jX1H9a9o27KhG63ciCdq5US42WTQzQx
ZKs7f7iX59eeE7hYeEuRjo4pfYLg7hVJx14htVxCdG2hFoA8WY9Fsg+wKfhq8TK6gMlg01mmWs9J
ieIOXWwktj48lYLwZd0L41JfDw/FOuu/fYHtTWNL2mdjN2L1Rio5seyBoL7bfTlBZQUTIbGlo/V8
14R3aa9yjMTf5h2krNTqnDP4PYtt36kTTyVYG4Tg7x4akNnk9GQRuKZWT2kezNTvYbmbcB31z5mv
ykb/4hq0q0GBZ0J1UbPw5CXt83HOUhMOu2l1/VcZJIMY6O2QFh1wPwyU45gTluDo3vy7P7v/nslJ
uUQuj2OMOo2ZmzrKbSJ5mL2K5spjEp9ls85i7wAG+N8K2C7YcDeNRoOQTKI/8sfYrOAugJMAJTTA
oANgdnqh9oJ1ihU3cZQdZVrQECYte0UsmT7WHj/HandJBAc6FmPKX/SMgtq4MEfUvmMx6SNUuJOl
lR0MRvwHV0gCJfzmdpBi6jK4+lijP8S+R86vlbS0c0d3ayr8aKRnMZ27CUrI3/ymwTafNSom+NHy
JMsbQ6bsFo2WP9JY8/J9pXCnGzSKftngTIEbQ2Wbb2n2WZOw9QI+tYU0GtmjtcIc1Ppxf08Oa870
eEE7SxbIqFy9kc+L40XdGC907jzg6MugNqARSu4QsPqQ7sH3V1P9meJfZu2GexnGW9moLzpn0L3G
xGbrssJpoWstXul3nlNmFhiFG0E9ngu3ENjhOjP4YNuCo8sPtzJ2gLzX8ZBii0QxRjO6DyhBlolC
ac26H5hp7epJj2nziAR/8nChkFxoLG5uhAmezfyA/0d8VIy2Hl/BWJMLLPecAngN84w07w5AdIZy
dFeM+xLDz52VHq4brSpfqq09O/DYU7mB0rILNO/veCJbwjVcMm3Gf5MSGGbz+f7/knRulza08rFi
L+bNeCBzEPZJFpFGGZF8b9KhSK5aCUPXXBBhOG4vpozqvV/ApWcqmwU+pl/4rJGWJqO4yewZ70xE
u4c40RbDPvIPkwrdgHJGFcv0iVqNlNr9PayuKqasfFGOcBladXBLqQXv9rrmDGnIRXMTiM6Iscap
ZDGkLp0wAKW/3dyHyX2Q82nbFrgnYZLdBaZiEDv2xyld8gqVP7sjAbJ4eY7Ntw4Ek4pQknf6RO9Z
9U2MXmgVb7ZFhIW8t8nVmdlUm7pUjaUswdID9a3GeKUBi6ikrrdq8RU5NHvjDhUDZgTYpu6Wx5KC
+IGEfWIYXl82n/FIXckG88QA1kKQn9j0GmIqJPCJi09t5SJK1eJ65lghfiAe5gL0zGZ3UGS7bH+1
nyz/LaUEYhSX100ymsq+5PJSd/wOIrlXazMTnwVMFIPS9LsWEWS4UHT0n68ZLAoNTfzuQUN/1Y+x
QlIKywoY9Q0G8nZbkn8sDWpK3Brg9w9tMQs7Gq20cpFtepG3QGeMImglXf223xFk8SwL9MR5J1j2
bj9OeGHx+friyvxap/ZXsYWdTzBNi9u4Crk50in4N9DRxOK3q6pIdalPZEmzHEHfy/kVV2SHrPYA
dTRF1swNs1YoFhn8SOD0KRJ8OqvJXHqwBRnP9r3OVtgkWTQ5MejxHvd5R4gaHmqAEPAloKmDPfMq
J0H1hKy6H+0lsH/YXQAqHbv7kbFqg161ntwWb+TzmIdqFViux4mW8Ve42lQIrBCcqqrBW7KO1gzV
dpX+fO+/rbEQrSsmahe003mqyeaoB/YD8x2OXWxqBnMj6nTAGe1GqJBOsKbV4tZ3U/3ZkWbPa7Z/
sWMsRzM/vZyMjskhGOkMcmav3ARWQlHZxNMVE3jXJnRETPuN8pehTWdoZdiGkYjN0MXjikvr+I/w
MGYGwxJpgTQYbmGoLRFBe8zJWA5fF1s+xgn0ritsbhNalihm326Xzv+BvjJCPudvEA7qv2koktNj
sGtY51AO/sbLvJra5ygdpTcHVMytIZFeeOnRm2m27LOGkEEcsxCN8urYt7V4KwcS3DmCt0TlQsZl
vykYODd9SPfe4LCPezPYq7tkmex4+zOtnNCkl+eWT+UQifmfdsZMX7PnIEe+xfv6PiUQAvjqF+pg
iF8rbtcZOPCgLfq+tyPxD+crQL+bUIl3o1iLT0m005qurQOiZLlqm8vEsARPrtLqnLiKzYqBSXzf
vI98D+pHrzjJjwk5wlmjD6u5TIqEkpu96XQ7oh1zU45Jz5AP/x7hxevxt+ISQNTlHa8x3nd0em4R
ZvTg1UM03jK3/vlMMZLG3Xrb4rqhXQliH8Z/xKGDnSjYh7ZeQlHG5RwFubFjBA0IveDwQ+oEe52L
bwWeI024GSdAOHDoO9earXhQTH8lz7dURnFUNSJ0GoQ/GiGwsi941FNNp5f3ZfEKTHmSx6og9kV0
PbkMazn+XfRXuSEDdEgkhudWgeuBQ3GuRFI1mOvClChUXt/iN4MCwa6pDxkHPv7spMqa2LdfOEBU
FZ0aYscasjiuSE8Q/W995UtMgs092Qla7Z0JtTV7dstHIBxPVRjiMEabe9QxWnNFfwZM/9vs3WC+
YBo4+NAN4mj12yCr2Xna2Mt5xmOWzfQ7soTBYncETKHcNeH+TQXWgCyPijj5/dcvcBbKgt5nT9fi
2w092hLx+R2rXrccwXKBbV5QuqS6tIgx3XrSMqsjVXqk/Onk/A5w9Ha1IIMhb9GYmxitgwuLcmHi
L6VZQQq9G2f6tjBD5N00CrjGT8AL/0e5lvl89IqgiHMr+Tsqi3fASFL155BEooLTaI2L9YQKb9+Y
LTjmrQhhptFgMrynxC4SEZ5KIGCmoBE/n7LSQTd7t1vLGdUgPL+DGjuJnxAk9cj6kpGkMZU7HYwH
e/LZNtM+LZAvOZBi3Pnl8Vijp8H3Qi4bOi4G/124q1BgxsvczNY8HCC2Is5kVu/YUc1DOus6l38/
eCXO22Kb7VoDgqO5eBSVc9an5Si7bPEnGU/AFTSsJq6P4vGhyWTktm/UDa1EC0PBkZRcYpVeEi2I
jHNnWI1XGrv08kZgXisVyoX1gdosFrR/DjT9WcVlTC0bRygwi43x/RpVx9dzWI1Xk24MooPQf4GY
SCmKlycRcIYjdjqMWVzD7isDLVSdkyL5kQ9YzhgSBR6H0FvHicT1ZHl84JXIvlUV9Sv4hS66J8lC
D+O8yljzHlZYcULi4UWSZEE8oaD6SwZvLtiA2vZ80I5r9ji0kszAN0dJFJoTfBwZxrzCSX9P1iAe
jsi1oHoVa3jaAx5HR0lwN57IqrP3zNd38kSoLd4XiqIQClk+AIgaN4krptfjVnZWgKRkn7GBX+nz
i5vDJcTSqq/6B4vNTxJ4gX3dicJH5H4jr0ar0fMHy5kNGWW3MRO+bP2zVATGr5Q6f7OtWLd/4shP
ywFXOE83fI1A6V9Wgkkexf2BWBwSKDAfaP2Z2pQVx2aQ/kWWj4Q8AiuwT419FyBekl/EFqfhdsAD
5OlVellEtd+SBTAnUre5iafLdnphQ/byEWFffOTrhanX/TgxmfN2iJhh15cm5krX0uTkslr/grMe
5BBvu6NAOmu2Vu+wvPF5quHWcQpkerDsRGwt0AyDhUR3Zg5e4x8s9S5reFWPJbFLaoBQraaEXj1g
Imat1B0hF4orJ7kFx8IlVrNfexUkcyiwuHwltC44ougkJSC5CzOq6WAHv6oIcxHWCnkSRsBcHQlP
U8R9cwH+7+0VGux/UyW5BdGYoQjcaOY9GgufAulbMBsYhciiL7wn4eBazGWE9u+RI51z60h08gFa
J7ZpocBGsCVVxpSYwmE5O7spF7VjQYjQc6+1m5wGy3S1LMsC2sM0/GvWC0ZcHyMsTg70lfmsRqiJ
70Q9EHqXdM/zFKBXdNGuIVqTPCOpSF5+v9NYi46tQieZYXCeAQZYWgt/7f/wIOJMwU6v5Vn88xEt
nCXCZ0Bppq/RhfsCDmjTAtzBtLjIHzCYdXFJndZYa9Z7AqhZtvDTDFBO/6Hf0UDufiatxd59DuC/
4CKef4NXjWhuTFQiQAk1GZ+gnDtG+QTibgPVinDQVO4qdphodgk2cSU0gxnLQ7tzmGLrEXYuVXc5
2EGOI+LumSWl1eLrmPHS0U0J1gGGbRU8Z8PtXV/CskIS0qam3KogOmVBQqTO5Q38quRjmu1Hw4n1
qFNODNOr6uOMaCr22BvD0UkZ70qPEa/gxfZiZZXbmkSD+lWgMfPsqGZBJHk4ky1IKjZmmgQsODDC
yjJGWeQdm/nCnqlQy4qCTNbxQBc9x8FWY9Ei6/ghiUlQMcwpF1G3SysTynKhNqG8jCktynvFIhLf
descNAKb9Hj2RwKIw/7Eebj4FEZTLzm8SrM7Ly2v6lVQNmlj2yRJfXcmzpjNzCy98NL76zRys2IG
y17HsO8B4lU968KcAuI8/RTwa/I6elAUSx7tsjzTFgJQ4+f3pkwYDBlBfErltBdFtU2K9FGgWURe
cJie3MsjJOO4PVQJEvK691TtY4noRqG4eyHPVdIRgX6QQBn1Y/L+SPtkFvOuenc1x5Cl9FSTCPd5
cchfV+ujon+QguSigHcoZs3zz1F5HeIOFtgaKNiJUWm6HeTcWCWc7h1qfa+gpRq+R6oV61yk5LM4
wFjIINxXWbSXPlIM8Kvc5hY83GCAC/FW1p4MQV1gS1OTjLEWIuGYbr8yQTXASfIY5H6R+weiIHjG
jw0xciAyxr2gU8AjPkEqfkPGL0m8LJY48OOkxDMckV4tvzM/MDV/0FwbvhJatxwl3hF3eGhBL9Ho
Uxu/souCx4b5XwQSZtQnPaT6Wj6H8bcarGrmuQBLXlz7kfQ8cbW0pP0OJppxcFMpK0DcWHVhXutR
cfCojCX6KH9lofk+JUdD8YCnb2KBlBEaaYVfiqUaQy2EETjCvtAIWW3dslvZEgAhv/KvVf00GGsJ
8vwB0EXUhHURbWZhg8yCr28QFmg9Sa5hKJ+MVLVCAY+oFC66XmCg4dO5RdoqzlqbKoy1p6zuwbVD
MP0j5tELUg4mItdEKmlJUVEbiMszWo0QZqd8ubt/ZKSctNbGxPvzINyh0Y3HH8MaWbxzDaHMGqz/
1zhv0pdA3AuqiJOp/lsUD6X4CQbJaBlHLwidYO8QfHK8iFWYeLxF2vUGH4Ose8M2+eJr6Uj+RrAm
xPsMooRcOTT3moEhWNybzKnXntjS9IAit7Ervm/YU8rRIhLrYyPnPWfF/UzcAuJArlnb090pdM9X
x4NKPE56aHrbWXJ31/1hqvt+QYTeNMi4G5ANxB6ogWtYHllo3mAAjOXkG+ihYceZmrq4g5aFDnty
J5PGwKExcR7V0/PsuFxo899GAV8x6UlgmhyGT+ugq3yJemMI6qrISSx79rcy+3tj+FLlSweNGYTu
B0LoH2YjcerqpWu5EtMNOhjKtM5/4Wl3BHTQGfDaTDvE05iWVS2QzvHGrk0B15nSZUIDwNn5Uw/1
8DpPsWD7E5I3A8TilWwCoMiUHV7ddFB22eIEouuvBfxcJOwfryfdEy4OyKuCrnaqZWmrfwNKa3iI
v5Rh2ueiSYZeKK89N+Q37KeiRq1UiJWNjaU8Tqi1FJ4VrbcbdFYkLByy4d26aB9UomxmON2GZ0Nn
SZAgMzyMQL9sBezMARqjbZfzuwr1hUoYuQmbymatYvooyDAPcHf5WrIHzk6Q6EEl6iV5FaDAGQT9
1dTqYdmfj3SpEC5gNxeRBVldZihqWTki72Baied79YUUI6ga9OJrCBDck02UvTLarbNX7BtNvEc+
d3+j08VfzoIYKZ0s2rhneq0zf29cCaJ7066ODOZa9jVzDMKYwT6RUsuirXBR4Q/aRLeoNmKnNax7
7+Yiu834uxp18BjiMVfA7CHeW2FFbEbzvw6kDU5XVg4uLyw2YOyNsD/mTeG9y3kuYwlBw0s8fnfX
Q/mB9B9ssBgOs+DmABqE/pcIXXgy65OwPQ8r1kdhDFVU5jTODbPOTVxyx7oKHdL/s5f0+sGefyA8
uLTTAZcsjJHG9T3P9p9rWpuRvqX7dcm7sumxpnGOZP6/p28GMPFV+87iitqcHsxPql4bd2ZQp38N
V2/y+GyXLC7Ui6bBG1HfOH/laj0G6DazNNSQt6Pya5hr9waTy0IwhwobRqSbxKFSFwC56wt5PPX7
AHlwrwX9LhiVWIMm4/19tSIvbx3M9Zk62Jzg28MUdG4GRPr7H0VzQyUysVx86nWWqe309ZrYQBJm
0FSjxERT4ghdWfB/7etkeZz+UN/XPc3B8uZLH1xFxzBxSGCNk5FqXWSmHh1kxVSKm01Ub3/n0BG6
uiOw4h/x0JiXeSraM9VKga3pfH932KlnGKs4nawaRK5pZjrGDBjJaR5u2surwvZEDNvJ62Nhc/hz
dw+mEWF6LYh5bImOsZIJcKqu0b3ZAYUpBdSVKyxdA5NeOmEryVyyR3FHCzV0CjMZM2ULTINZl3sN
F03yV1FLPRRljQyNRtKU4mJTqN4K1ODpH+ikLCyx12zIoLZr5OANDq/lWRzpBCgQhU8QovfkeCeO
B30OcMw6RmCeFlYn6BQPgLRhB4mLKHzDHY4b6laxjirHj34GZBK8rlQB+0+BQa/hWAEx5EpUfu58
AL56zrXQX6lXEMKtncVkUf4ac3XQiHf/9xmTNzZw900Z3og0+n12xeqak8npm1rwEzXGa2c3uRuG
52+PXMcTpkTq12X85wRlacC3pwg1RysUL2uDad0UrJ2jVUMHy+wFEPzwSLqT2iPBgPq3RYLrONpJ
z5YZrUbKpRasHVnKbmCH7HPLLsOsNpHOKj7PNCkqfKsUBKvkCLNXHZg2dO3kjBt1cwWTYVna+kiI
0LUDcO/YUJvp1Vbwb0wM4kXrN+tzbR6GJFqCieMIjFew7bdrXn2UXX99Bsv2EdK8xmcpJqAFf9ag
9P1aCfbuouVO99bhLuCwUe9k+vPk4bV7c7kedgjs3TcUC1tyy0KNF9IiLefmAq4z9hzCd3c5hr/c
8orS6Dv/pyqH/mR13LW5Eniaf6CCzvIo2A0LYkhbS7XqqkA6h1mao9F4WDUIh2puotHxrpC/bjBF
jJGwvMnP+mtYW7ddc3O9OL2LkSgpTIev5+Kp6HIB5H31/UK4e5FZSlkiTpBI/eQYKCSVHCO8gx2n
PZTj5GZohb/bJ57q4juAm5b9i+Updy5PcMD7nfLwt39ZXuMGoPO9W993XpsvM3uw6Kkqtrs0GN0R
e1P3OleGjjWJjuzV3I6nunEshlcX0h+EzmHTsKJaAxqCfwXnAWgw64M5bUjXaTnLsAsrMYkZibIt
arsulAeZxD5FZxv8G4+pb0lz/0A3utHCZNBlDSjT3a9sQxey3j+4LBpUqxaGQKjK5s9w1usaWKDw
fbNhh3CPMp58VrWueJeQ5/4e2jmiOWbdbudMZBKHD0PmBpo6mRYmoYgWp3EaiIzO5PNd//TtDy//
lhVkBfOUih6vvo5w+QAU+vDMv8PpcNooUsSWp0RY6ZZIpnQLra8UxwWPfhViMgUVEDUVtJKMWs2Y
2QDHmkPxZdUVyv8He3o5cpaBaCQkf7tuLEJX/Pn74glJbBzXqsGUyJLaQMPwW3hm9b+5KlPkeadA
fIHHAyvja/MsHlIdSGLCN8imIUVRUjXbNfLPdUDF4ALAg1DQUXXEt+K4p/kqilEYlWEOOASplLx4
1OC2KuyZ+7aUD3/Z40AGcd5K+yPtvRC7bIZ0Ea1riMHaniMalGbJoiwo/b3fv/7zIb3UPUm4G0GV
ir9ueyyvJlvldlg+0TUDFkkMhRMXXN3q39A+HlM/9HsMOpZxy8J2r6rLydVyedPsjgT6smSDeDQ0
WNRpg1kOM+UDlfA1/5m3zFmleBtYv9SoPwOunf5CB8WubnuWWw0wvf3AdnOjXj3nMMFJ9RYRzY+F
PX9YvtzusgT/aVJUV1Duk+NnaeUQCM2uWgpUt+P7140sCMAeDob64tIfitcUEMAi2RB9DZF01U2s
sJ1T70HV/zZmNz4YAZGhWxMKbV0K1mXjBA+zxQv0hNQKGXIWYan4L3ABvbCt4NcsUqdXFov+cE1X
QTIkDld8BLtZAVa6iP58PyN5Bff1mLc2BHk5m/mFCVAyj5Kbfk5dfcgT6oyIZ0Qe/Xv8g9AHS2Ys
rhN4fHkGiYmMPzQ/2UuRT9xtZKAbnGcIEU2mXJHi6B42iMU7C1QBM0TrUlCBQfA32olrh5VsXNsS
b4b/57+kqofMqgWFWP1lqdq+GWX+1cYwV3n3ummgY7bZwwORqMkaqOpa+7ZgUBb0rmsDcJdFXuVc
7S44CZqI8CXEcsP9QOORtr/A3jtKpsDzSpd0yoIf+o9nJBo1+9fwkpTHIeUmkrlgv3YLPFmiMfuY
+oxkCUSr/QrUJr61LjVNTt9eYt9UVi9mw1pL9PNici7IVXLp7l+2Mum95ug0WKZAgQqUuDYb9tKH
T+p4xNDKVYjVcIe7CP6L8STHHXkQTfKWF983J9+PRGEssHDQ70Re22NVXpIhDdo7U8CnMwuy4tt9
VAdAQyDJdmhqaOV/Rexp2xLP3DlFdVsezjJiqZ1KHpTE2HC8uzVqpSg19g0ne+luXT9RBpzcw9d0
wUGFpGR4UKxTlpm6ugQKyv8ZWgvHMhmRNvWG3wnPrbhhIEQlIFgPxmoKPojwwwYHgUd7CIAfAm0K
c3N0eoa++k2qU3WccOQbmN+EveWozR4MG9/J83rN+MJRLJMNm6C6a1zLQO82DuKp9vLUG2wZ9fVw
lTOoTKYckRuaZwMDE2RLZrr5/LZ0e2RGf+Vg18R3w99tPBPnniYOeKVOkTn2rP/3VtOTkEArmlYK
4GLrrAGja189muOgT3VGbYK+J40ErT7Mklk2gc1OgW5DKiZX1yY75yx7+1imLdJGCbZr3t82mXkd
ZnhvhInohWrYVkVvqjtN0LSoqAjfZKxRfU4bkFubzu5ORL5Pwi9BPFL3gDeT1JRwBTZvcRDkV8Gb
9H+3LdUK9dtFVO/02RMCT72e37guYGnZm60npj2ytTHpml/4KcW3qBNOPQYGcaNmj9UOFSDZ/UsB
xKcy9ARQuRjPNEOuGGMR6XFOngub+M6I/HLOWL8remgAu4a/gtnY1qjfSEtDvAlHDW8HJ9tv9f9N
K4QAhHOBPmpuO2rjp6DMB3ilD40KI1cJ7GEWVL99LrU05ZZSKgbHZe8O8UU+1nQQgeny0btord4e
RVxJS5hOGACmdk7ielb/PnMVGq2v2Ksg7vdtDUVggF3fKX0X5OmiCSJfFIGUPLlFS+AAZ3E7Y+w1
PTjibz9WLMCRj02XUWQs+NRFUv7xXNeHwQjLKBFI321Q8DzvS3PsWDQZeqp4/yv3NnGJgYcUuvWV
Vxlzc8gG+wE6ZeCXvxtOdzmqxIU3092szt0c6n06vZ4tAbv8nouStXWkS3TGZlfH4wQlm1rBnCga
x9R13NScqsNNZGWz6zzPRKt7/8b4Z6WgYCafzMX0zLppGWssJIPXGXLaMKmi9klsmbpJ7NdxRgy5
1geKr9tXixTXdPL2WEQwx3g7F4CIWjLOeB57Viu9e0ZHrTY5MhwDyrUCM8TKFjNX9y+NXyMJsX6z
p6Di4jPIauSnGtNIch4W0iC5MnXPXT7vkxV4GpDYJ9+YIF3nwkA6usEU8rnuW0Ned6Hjz1oWrSbq
Eyb+CFrFZtLvxfEqIfT2uCu1hBPA7jDZO+GHXduRmi46S4YTZvFuyb+056J1Ezvo2zLhHTE442pe
1NZpCiSGZa//Rf0JF6N/O9/dFhm+mciVqNDdxTYA4keJCI0a8HrToOs9vviojEKadqH8IiNQHuu1
/oYyLsK6D/JztNX/YxChTXiy8DEyx2En5HurbuvIe+R33vERPF5yvxYgBMx8zsn6X6YTnYlRjxpB
0cqKo/sKWw4D0rL5uYK2CV8zpd97/WyYyp2KQm/Dtl/YmQHh2kP0ofN5tjWh9d7MNJp6gHWP3vKE
+nZ1QlKir2xwiRDBF3kWdYbCUufPvEPP8sFwvRapRpXgvPqSEFOGFoJWlkEk8JKcOMPFcdY553zw
oMU8aAgKidI3QAZaC/1qFHuor8OacE3qLzinqyoQu68J6bw+nalaQveIl9O08vcQnPTto2KGJoHw
O5WpHhut8XYJ5uAiZb65CYD9XIauseBa2xl3R+MoUqieBOZH4AX1+mJ1tgKWcrL9GSi/+3UC249o
Yj76ZzqPMv3wcoxZfpT86nQG/6JqxNcBYMbFDVhyHhtPySZLtINl90mU5irtNbNzGJ5F03RN6HSo
HkQ20/4E3PMQi2QPWYvgqgyU9uwuwrcKtZbeDdjgBmRG/FVAmtNMfl4JRClquql6pgBXeMwuAxmV
DLapBHzMVyUeReLpQyJpkajj7L/5ZMbKMD3PrdQUsxoIGnE1MuJC6tEslcCxxueEwDG7v6HOYB21
yts2W2SGTQ4XYBqSVJKSaxtTDp/D6pk0mJ0pLlfw3z2utAsA10JfbS1mdFCTBkmjU4YiiLC+UM9w
MYRm0tt7AzKjxZGGIST9c7RpnRjOd8iVxkSndCHSqDlmrlvzRZY3ecdQfZffsYwQPqnlWrJ8R87/
Iq6svTfWUQe4yaxT7sygJCvnQlyKhxeBGfKhhJP+lwExOQ12SpI3r4yrK7Y+NZaY0n9YCTntV2cO
6zFdn4NVkhbpL7aJQere323q3vimpHIUdmPmzJU/bvmUHpXtAEfylGPL7/5z7R3jdd7URjD5NcJz
NrKDz68l1pEdiyIj4YUYTdd5nzJMhneYcQTKlACxqbUZSQs6y/LwkcN9OvQ6tfZtKBiUzo+6Vy5T
YP8YAjC8rm6CC7BMxMmc2ZH5E9SpzqKIFz/APoI9Z65LWeERt83p+fJqItj+tmZ6nL93hCu2UAMV
wF1rvJi6vLfpc9j0QTo8RzH7bML7sYhHqJzCc+uAIOSLphULC6qUuOc2nUKSY9c8htT9U/ws6uM3
1iW0Dn1cXT0hXqwUhamrcrCgxCWoF7ExkTqCZIicbGp8dwrxa9r++9djFVf/Wr8O/EwvknmS3S0W
tUXlrZn6rYKEBq6t2BBBz2WfHeTBAEDNF9rHLdobgkIBJVCQ21Ku7vwH/8QPELvJeviLrckk3tx3
/YMWjLrwlz+k/W8JBe/rH/LXZro1pQLZb9Pwq0qZppBYuu6ECjbD3HQAclwb5jv26ea7CqpMEu4e
TahbfPO0Jk4VyMg9BcQ1Y6oeFDzDklFjh7lyLKNu8JIYUqcFBCMNtBJfemtNa+o3dgSWegtwOpWz
00CXf0z6VJ1P5rTpNUnBMgCBFj3hLn/RZClKRa1AsyYnNZ4+csDsRYRsvX0S+SUCkWKpUVsSLAKY
9q2Fvcp365CS8qdcLNyJsnR79TO6M7UIoIDSdFz3aULAyE9U7rGdIZa1Ea/3GyUGyUnUEcD2qknF
X/vdWzqoGYwZ8HJm0k+cE8FnVco1CHCyW+N9Mh/Kjq+6WexjB6IZ4WF+Chcc0aXOxKKYi/JuX69H
NWuuuhL5I7Lrv3r38iH2BTd1yHh19fGekYU2oNtQ8S2LoQBIUnhNz6rRvH0aJUV2Vt8m+NG5349p
iFiD7/Kec/ymsxSJqAYmWIR63YtzQ8uCDdEt+4nTqq3NwojUWGKEgJB19qqYKglX8d66ciAYgKCt
u7sCLmXU9Ls4fVAnEw2WlF2VPeXRDqL1zxbZSUlw0D7sPq5WK+Tk/aUVTHwBJoeeBq4fX58fx4AG
vinUplxTh1MHW0UjPwabfaqZ7Zocir7mqO3syrb7CPEctkLnuOtg8W7H2B01UDTAyFySBL8NNC2V
jcitOfKOwDQveTsVMmuxCMLhvRou2WToQe2/VQggnjZuFeL7cGtRbHhloujAKTS+H0PGQUV1DjkI
3AU8bQa7ijf+UvkvSbqwexnby40klRxMEaIniODXO41Lr1LFYcwD2mV37aXLyIABWDT0ba6FCsky
SCjoM7xd6PjNpSMdkkL6jZcdNHBwtb5xFCKboVZin3h5PiynERBadtaXasN4pX2qJu1Z1XiteJQ0
5Sm0TU9KzGvT6zj+lZfzm1JnL6f0FGgSUQGN9NpkX8MZG0M7sRxKghivuH/+7ntpFImK8md7fDjR
SK8k2stzllC/yXMIJ8gdBLHVXlvtn3M8f0nCLbpoWZbGnZSo6LHBvTZUbyKJ0Qr50RCpfom1VfOn
9dbNpWYlC8vhmJgF8T5skSyBE+6q7+6WzTQ3cn1dA3Pfx087KJvwjEz+2Hl2kg1J+hYVyIkTsAYf
tvQmylJBXwf1gxLceLie8uy/drlyBz9NnJIGnc6+6el6fcv2+Ap1xQLoaQmRK/bcGlHlmU7RYmzE
kadlGPm0+gmfQfCZiUsaLUFCI4L1dRS3Rx5ZQDHpYs3xtB0ZuRt3G8GwgAQjFaUr3p9k2cX4LSJB
LLWQ8kI/fOYMLFnfVYMysraXTkTP87HLiD/85QlCi7Qh6sFmqrcD/JbPGD8ozI73vLBebsiuyq9E
vhblfGAvLWfkfWZpMHGiuqtNLCjK8CqCqlEN6VAqvLf5DYYesmkf0Gf3kfKum8fBPj/2OW0ZOgvp
y8wwIEyMeJBt8yYosYyH+eNJTsy2mn+kQIiKPcIwqcPi5J4pr+m7Sg4jJwL9mjhJPdMl9pAZJi/C
PMDtmtAos2jAzUlbYqAHyqTTJ8KeZH1djP9hgTxBxmYKONz82Kg6vpxcXeUPpJ5MWLdm6A4pvZ/T
RVvecINXLRHowKfkEc4/uZmP9DnagLUIVcbb1X3fLgupSxDhGKHJLEpNHQZ20Ca8ykL6zotiTu71
N5vvmqtxVwZsKuTQQoIwsu7+xqWDwjRtbT6MrNa2qWt6aE17mEbtu/BqhrQXzD0VIh+5xhEIcJ7M
IzcbIzq+UoVNQ/WsYPDwLCazaSjzcgkX4Lf7d6PrDow+Sz9+6wxKqMhykMTLHFL2zzXPImvZI7dH
drVCxp04x9KnFVFkKTmK3qcI5BBcOd8dkqxBFA2jRojZCbE4ggfrHbe0zi+Twc2ot0htnf1DiZ1p
BEb8SB4kKyarbXp6N/D0SbOL44AjqYx2meaDn/VWlSlBed27qhDQDaq1+p3IMYTMvckaDJK2pxx6
tYw3k81vmMCYfAG3Nm9D/NeawofihzV+6yYVt7ZWstLvKbnEfbjAGHQLeYMtbNrtgDxSzCtz30G1
mg8S5fctTjMhdXYv/8Slj/q4xNWfn3MfjfGlPxeFkoBwGc4LWAh8S2Sn/IOQf8PMbS9AnMdV3tAW
YyxKGTym2ucmAgH18s5BlgcWLTxdMik1rMQWhv2q6Djt+d5qBDVgHWSqhhy9bllqWmAQlqUyDWz7
O0J7R4YbtvOCSfZVdsc7b5LhuZdLCW9NgDEzigC0Nzzyn8mmg+PaaWN3Ltwu6QCHcVLD6KrvZ7V2
CEfxBIUWVuVKMxwQjACcT4JNfnfiK1f1Ay7gXfcGCOduc3ukuGRH+SofZPtUXhNbbsTe4b1BP3sO
J5AzdMP4jVhShyZUMXfmMYEEkzhr/EdTGzK2Ke35NkbIBMeoNwORdWddv93ul7xwqNJ4CntnaigN
It/Xe91axDZAruXnAA5VtMwWXLzU7OSy69HRWX7tQQpkg02rBZIV9EdkagNdEhbyrkZ69Y7BcW4Z
4rwkEVnrR4l2CeJrpBqOc0+BiFDgQMLk+vgwIQZoZslzWcYn2QLBrUdStjuRxs3tujA+LKJw4jTQ
NQQ1j0Pi+NydGcaRkYuFyoLSVzi9JdCpBjeEAVG92oAdkyXl3qMREODFINJjkiZ5CLkNvLgv/SMs
qIq2Y3re+IIA7aHQgRqukRZjDdVLNTNTxvDghJUWipOEQ43qjhsyIzLBy4mxXaZoQGFdURjMsx9a
9IRGvCefDBgtueKSQ3PxA2uETxDs0pLTxunKCsiqIAFzDajX1vePOvQihnSsMjWhb+QcoZesufQN
WzJAn4Zl/g2Lae7IuQTbmElTQkigv6Y52MRQqMMnvwnif2IWLIW2KFVqYkhJo0/iTZweYjcAXVl9
0QHgfXe+A8iWxlo3LEePKPorn1nJvNLe2PG6duWKlUYUPY5K5k/MTo1xik0dptWSIVhq+x5uFb52
43YtO+TxjtscW2kNuOOj09BQP8vrRfwNGtIbS26dr4VQ7xo4DSUAsXuwqHEdg9g1flYzSDmEHOL7
TN5qgdG0k2xo5wmStVLWGyZKAEpTx4gdJtRw1qBE5tnlLImtkqem+QHTIMFh9ZctjZO1WeEcj/wN
VA9KT/P+mZim+ZLvdgkrbOzYCBW1n2vRhwOkzCzWX2wzRd/MDYA+Q/pd0Av61MLfM+wOLAZPYoUk
cN/t6F0E11vWDPBUomCYnJYIuf639Li24qdHeneNXsAvgUOxkmbZlpsP698KkCL+7wps+48S9maM
Z1t/TJRRV6K9xjmNmVOoHRXbH3WyE2p5qUvlOpqwHrUuuaBqmk/oUh3fNYSryxxF5UkG5wg8ieMp
0mYm4P1oRJJOwkFZVFAySwYMqX0SCAhTm1oJu7PZwOKamoGz0Z0HKQmXZaBUhj+AuDrwmnylrVvt
Gm5AMKzobMKP27v3KmD6EyyLIpq8WemZHDE6A4HwdFd/WVFuum8X5pgNAsLpcrV6S86sqGXNyflg
a4ZD6VRQ2k/A4sCJtB5obrgUvZbOIh2NDWf89YQue+vK1eQN8CE53ybM809CdHzjm4Z9tx1x0itv
Bhs3seKOTjeQnSYnuBayZq/4bXd1Qt97tIN0JZpB5jZ6zLZ46uq+8RjmMee1fHzhxFg54J5b0BHU
9DOplC0xM9NptHAvcJWs8o0pCO76SVf2wNeCDJApLwn+mZy1+jUmG3C9OMv7lZWyW4u0+76bMZLa
IaWqhU+nMZD86a7FGZZl5djcICVn3T46hAxaE1uNke79Un1y0WSJBq53nXfYJ+mn3ZoCGTPGypl5
D0f01Y/CGi/7fdFUe9IdGZnBXTwee8qFusl+PoDxq8pC6cEb9P6DleiDmlbXBcqNFp0LuoEgGQ7R
UJj2jtpCAWAXacsjbGMePO0nRad561cVPrk/JhzddwXJUKtPEw+LA5fyPqHvF+fJ9cJVsSeoSYTY
j1Gm7ctZeHXPqfehdw+nginAEc5o0vVModqS+bblhDQC6Lxr11FEHxY2J3llDps7Huz4srXvKFqx
/msdwziyxaX3VxgtNBS6HPh2DZF2s/POOzkiIctsmunBSSCKxSv/HonsV9xPFzF0F8pyG8nYMHfu
4spZaZqGNgyRtWE8xGVwWmbgZT7lc4S2yxiA+QulYlpklEzWvw97W4bf43CO/0c6LWhK3V4eUixl
hdSi1MpHlURlUgNrraEFPzrNQ5PFNNGJv0kwu1eypCmO4TBSGTqKmf1hB4brxZohSPwOm6WaBZFZ
9d3Yx9PexXxfWD/ixi2114Dg0WD4hcpSIlSkR8NzH0FNrTkqbbySAji0XsW2lV7g4VuDfEnyibv/
ZmSiFwUad5uTBgEKIXo2vBMWY2kMO8o/IqONKVA8GslKJn4USyAj0S+sTgZGgWMHOW7eeUbUNooJ
q8T892xjoioqqPju/8D/s7iWDdygS/pNk6l3slA5m+HfLMTEqWCUoJSShvXbRoBRMhjKr0fXCu3c
nDk2xUo2jUDnHJgl0UURR3HwHN/ZSXCkgBng9vIVDR45F8cp4obMUCdUKQ4OzGZzUxF53UKiT8r+
57dqPutFLIMsMyY5YPP00EQJf6Q20hJGUzxBtK0JkKx/RAwqzC8/lNplf++wUSoA/dba3Cu08EUF
RCWmFZmYQD2xsECuoFF9yQKQOi63bR3/e3a9mAhvOpnEEQpSgsDYHvudTRvIFrvOn6OFgkJpNh9u
zDX65xjHy3YOmpNeGX9MtZ5E1SjRfKL+zQXQciEXGVCKLQkgv6ZeBNSOaDLupHLdqyWX9fx9FOQM
RykzAdVusJ5jm9PoYnT01X886jpyvbsetcePu6If70qcb7gftSSqEKSpBPSmxYPAeKIKIxGtulvz
ecJwrCbzfNXMgGuaqrND/j1Y8ID4UHFmZhE4wrYtXhFnd2CYXTSSSJvNhb8Ym3/R+XoaxjUVT3hh
+5L4anGnD9fWGNuVB/pm6VKDKd262GVgJeKdHFf5bEK3ioxtpyMzRg4glWQoK1UCDYslZPMOQzV/
GrwFRPaWfswmvg/zDet/uVa8uJtLyJk5lnLL8u/0OnLFIqFmGbhwmg7NF5QFlShvP9Lu5jwOokxr
69Iq3QkT0Y2QyPyh8vKbrEmAk9ECjAJl2FlOslDyb3h6O94pqBywbnZexyiGXPDZAPdW3BKhiRRM
1qDMtq3RC1fqu7n0yVzHcj4rqRYW4h+egujax9yOLvhE0MY9347qqXhHCBt6cE3BHBEReuyHsy2b
ZtkJj5fl7Ceh2cQKQ6Q0HwpKcWivgN+3u5H6nXsL0geTOASjLj+8nEbyckuxGi/js8VrkhhPQfsY
cXAzE3kReVfgWSZbDJJ0vEEaPJP3GzubDVy0inRZp3UJI6Ne6usPYRC3wu/PXhuSZLh4KcBj9UqG
klTNc4eLILSSOXmcqKB5gdKAmVcKOIGQgB8fNYvaTPXOrzhQfVuMFxAQ5p3yWDbQOVgDsSFGSP8o
t0POKEHsVGzCroZ+z4MttW7dx4f5+EzEZuXCC/3StlKdZIeEGptlhUCqsLPt9WV/p6FyNTFy3wSE
4bBPDeSKyI3cmM2QR0KXhoZ8/hyxbApB1Eae61hKfsLLBRnBir4WziIsHrYRdopjAyvU+qWKE9gJ
Ni1ifysES1KEF6XHjbqnVJ6NEwUOKz360j/2iMTSJoBxKQVvqjJ5iVacWIwWrCf78snjYioEfUzI
aCR6dhUhSi5ESHsIi+AfzVQu3X67GqnoFXysbhq6fBVj3JZlprXs3gWatiEV5qIvMFodZLnWrkyl
2OjhqXK8GOjwFFV6ApQjtOVSrBUMVBCLdDsI7/Y2OhjtyThun0aoXcv4NZSYU2uXaIp/LyB20XqD
barWRoqCMXHC8C2nl9ceRlM6X1M8yunrybHez7D5qQ6hac5ST4J18DjKHq8/6EY8YzixID5uPu7h
aMFV29OFTYmnd6I87Vq5A0xuCWKe89Bfro3h/3ox4tz9yWuppgKr5gdPrv8shNMLWxKS2QolecPG
oe1fuownE+L0KWQ8Pg1R984exjFb9FXuCiFZCoUrAc1wuWVid/RyEatZx5NFjDmkpbrcuEqWlEP7
pmRqw0cRXGHGf3d0CB61OIi0U8KhvOh/qplchqsZkQiE3NFtau6XHmjP5KNU5ZGd1pfMpT32jv2H
uz3TyiI0yvAbg5kXWTsHejvo2aGj6UkgFp4vGMywiRqoZBEE8dwZxKHRZKnNwSbqo/Cx85pBC8N6
yYjKbq+wIkFIl+zQ0HYipnVunxPSyCLyw3b0fJw/k2KtAk1KlyQtBur2htq0nIkYVBu5IDp6mCPl
6hFeXfSf2nBiszDowK1Zm+6evTdTC1FaomlBHvgHUMYMAcSRsNuPaOMtrXWAizZ42W/fdwWaTy6X
Cnr7W6sJ+qyM3fXM2j5Ty3kpDy16MBlGHrsG6s66lcmsmumBsMgGsSnNevWs0dY5BeTcLdmTkQT/
wDf7z2X3yOJuiv4Kn+qB86O3YMZ41d77921Ki8Gdrli0jZR7Y2SQOEj6QWqMD1SZyODA/9e1u0kJ
lXzSYzU6HYAV3r0SnO/qlYGMcz9OUtGhOP0ONTPAJjqWaJc9dvaf5lq79wqXOx5EU4iRpoG4jmGI
w+tQl0yr/w7SR6CvtzAXDKg2TheS0lZuKU2WdoHrnDazji2J1RNxFZtcS2mADCLk+q2dvyC4qys/
oMQk5KPASmubDZpiYwjSjlEko9dBMdNwF0FjdQwvacGdnOJG9PLZrNkOJsFzeGUKUZVjwZqwj7U9
LfJ3ynDUcvUSLpPz+eXn0lTr06ogFbeo/oiGvkF956ws/KWtH9NUNThRuXVmUYsHTT4zpXKX1s0v
sP5Zoj5PlvAACye72OSpgLWWin+cSvdacTySSHSTh175By5kH2wLnHg1GypjHgRJw5B7HnOPJbda
5pDPmkV91DyHLsHLGq6IcezGMPT7uKCMvg3Kmuc0DH6H7kMTPt649slZO4IHe09qsLT1u1ttkN38
2X4Id5IMO5sUS6MiG22PnfBR2dl5RPJypo+xKvqiRiCNBRj/L5udXVS6/n0U7hoyLdR7plb7jVr/
BW7V77/I8O7MFuiSV6v622uGuoDbl+HapPTCTH4MUEHzBh7nw/Ba2TQnL1kJUq8SSYzF94gu07sv
oI5cKkyuWUH/vYPSmr5nYtW6PbodumMwg+J9WrpWs7vFArdGx52JO9RwsN6xJ4D4n7DKDjTK/xH7
ZLEXwoUeak1CMXXzMXv8XbmKiSgGCZi62/gvc5clAvuyVEcMa1qvQ0FHtknXrBnMM2eDDCRN3fzS
C3eIlnXMiMukAABczJA2iwgISljyhUIh/mgo3nQjguQ8FQgidtsiJuzRf3aLf+Vfj6Ia/KGsAyNu
D5vVMUBbJaOe0RbdY5mXtWwOfKwI8Dd1LopmnEIQ4lgpafpzfxL2jtStxZZ7wvMzETyGfYxKaS9U
9Itbb6xwCn2ovTJb+K8rersADLkMAoh/0FrmZ6g9bSaAcwtzX4lWgCqRZYeboa73S0oH5DZ9x1Q1
68D0isK3kMZPMIrllPHyRVa2KxOWy+dEG5rcM9EHcT5mJume8KTUTyN3BNdXPxQTW5K/J7uoQ5YX
F/+JVR6Z1Rc+NYDkt4eZsBJJA9EP+VbdDrDnarS/obd0KeoYX/xhdwjE9ntVmbCO4CQAf6QNUjOi
Ect5RJm94lbHwlOUXZJVs5FwRY9iH/irTQdoXXJuSlw5T7lC90y/rPPrTy0YgshBqNGX0CXvsLKh
uEsDwr7qTP3AcmIIYJu7zNP0EVrOs6G5ikfYQKD2sJ9daNm26bFdlYKnyfHCTZCV5/sUEziWxZCj
wX+1LS+mfBqjNe5Z+XUUUQmPL5T4O/8GOga8BJh5bldfOqGqMLQchOCiZC/LAlRJleoWEEmZbrws
bYyGim5hucJTKVisjhs60ob+ddGVOZsULCC1JDtOB11A9oJ9EdiwO36o+YGzJ3pLLA/WjviYiqSr
vTRLNB92jIk9dqpVzDjxD/cnuWMIX8KraCM2XLytxgjWW6UCGrPPdaivu6md/ltQYZqao1Hc7Ipr
W19nH2h1VNkYNudhpkueUHHkhgwOay56U2DfKDpivldhVeEiIXg2SuGWAXVSbMXSfpE1ewMElGTr
dSOPTcvZzCuGxcO25/QBwISSZHJbJ9gBLfy5SwPq5w4UNJYpFGJJZPtgAJUMEv/hoz6gimStGOTG
64D1xtUCqfu5tth6NVN1fLEW0si4kcKFbestN1Hl+iIvxXCIPPfPg107vDKKKk0IhuHHDh1/PEXb
pc9N/Txict1eiMhN1hcyo/yC/0l79V/+MIdCK0qv91p5MrD6IWubHCBqz+kIHXAvbAcxUkJ60Nqd
RLlwhv/OpyyQaRpHfk/kV3Ed/2yHcQ5bnJPlY3ZZzhB5MyXN9wQ/ECr1Wr2jtv/1NvdTcXRFghgx
61ke09sUqW+/oWT/VuDeFad1qLWG8sqv9Xahhq2gWDq6tbzB5gzy9GZq1URw6zzeDvdOCR52VMUy
+ckLktiA3w50otsDDpOw0RT9KWl1LGNWxZ3I/4h134EcFvYYrKGVnK2/72wP5x32vj7ALd7FpU+7
Fl7wXnBfdAYHjg23h7eZcaEVD4Mla24ERaL+NpQ62NAzSvxV1C5HSSQtZ6OP7YS6iFSXF6JTlZsD
mMyTpyPEaxDOUvCGw9MXkZSIVcT1GO4d5yJ1uON38DBvrelNCDU4dLmL4dWo29KZ2XwwruxP9spu
LPD8j/0e9GTyUIeE787GJx7ZGxra6YuGpSIs8FmUjAuAAQah10Hplu/qVXKT+wgoCB9zZB9x/qyw
bNvgukl4eJkBVRZtxb8sAouMbNdp61kJaE4ZBcpkK5E9j+jtvsQF6xHD2MCCaM5zjdY2JjfxHHpP
kjZ34slFDx3p7zdFOh9vRtX1AxlnVRJzqb9EIa8p3WhcY3Xkwm0wJCHAsAxndcimDyc06wLPijSq
S18n+hxUxG2mg1ZwDVXtLydt8Kao2lpRdO5zoOIpgVxEOrW+MVqCcHhvWWCyn7kjnCvOIR9D/vK1
8dHEgQLvsTeAvWzvkDx2QC3oEPNoV3lr/tLKD29oGA2mmDgD4JyN+Sf8y5ed5mX9IB3ji7eIk5lo
68lFujk0RJ+32uuZKBTMnipoFl9H1+P7n/pWmWVy78B23UhZdYG5O4M2+h1oMzJnWJZZMXgW/7Fp
sUh8ebQ9O4lTmC/QvBJ0ab6vwe35yVnGmv0NIJPsVk5nYf1iTIB+k5iZwLKrb/4T9cAW2WHCYe2m
yDOa4T4nXc+mdoEX1IPrLxeehvZ7VeYwktBh8QL98Mc5MMTRBYDuJoEIS8wbEdd6zIbH8duVjTcn
Zy1n1RWEPRhwjAAL2gex3uMfLmJTJAWwHHobtiLmUS7jD3ki1599gSJ3XTJVo1lq0bZTL3x5xNrw
eJV+D9TmxsAN7W0B8XrFkVKO37vR1lzAyU+bm6JjLW8NI3SEwrkjTNOts1PKDNCsxKWPhVByyfVI
TRs1y2nequSTsJjP7U3hQBt198sYPr7MxR3rBtuKaGNxioAgruWzNQS+uOtSm7BMHTR4m+k7Q013
yj7H/x+ARUwrY/J2QOIu824vozgfoggfM+c9iwJV9nVVqn6q6sZAv55SX/Cv/9TrRjYs6hC3zScl
VHv2jEek8IAnEAW7XzLIwTa5ZZzza5WuNLf3181pCaB5+MHlmCbHXTM14gsjyM3/7HlkoJYo++rd
2uJ2MO8bKUClCIKr1GtA5DDBLSAWBrbr3UhvqBo1TVKh4FVe4zr9Kt0OB4X8ComhX3mDF8ZI/Ov+
98P8I+d+0nagcUP8/xvzqb1sdZ1F8cYPDuy9sYj2Z+ZzrHQdzEgSBSGyq8QKttj47cTC1HrGnR2D
9etpRYETbyrAJ1cLU2gB2Zu457kx1NnPTG8ESrAreRnUdJ9E1TfgAcID9vvfejfeZKUE0htKJlk3
8P8vapMN0IvW0yrtyhsnnFrdTImocRT9k/RhFAhbrMmvcF6dF8QisSXPGKFmDIs+epNTu7OtIhBw
uR7c+ZngqTFA/RWoarIf9p5cI6H0oj39HJSc198q+/kqGBQDGpCz2mg56sXFx6jcYc/9jXbCYdyy
yuJI2b9N4l9pRSPtRMzbiN+W9zApoK5f0HMavsyadtgDVpK0K2g1G+kaLW77ERBJ6FKIWvffgQvQ
u88bFzRNfjEmHL7LsBEXSDpDhJfNXQ9+pxhICAt/eIsXSAz5Sc3IT0cOT5wrsdBbpKJYl7+JD5ul
Mwd/uwMdbbZNdWgxeCG+fARfbb0ZTk6Ib/RgybxTe3vTlABEjZ38xaozJNSCF0DdLPhjn3dKVPLg
mKy4WOcnO5HEhlHWW1ngubVNx8G7ghO/TynEFfMffBBpD7sfs7O+qUEIIfHpK6e7X11mXmpLS8cT
GOLPjO7L5b649EaeOw4v7HP7H8gruCdj9EwXiDomt+DojyMATEw4YefTRjD2r/PnO+VbHy0s3XPl
n4aHf8DedkiakYLv0xum9EWyu+tOh0E6w1jfq/khSQWRcrztGX/QgjEh1nr5XJ1xGm1uHOzLfbhu
FkwlrNRwi0u/q1Qv0iB7nqZPTEPyzjnqqkc0PslMyM0UnwtvQ4msOlyS+K7ff7vNlyiyQ1uY5Kgj
FdX2uCTGVYrQKRvZHWeVJ4UCesM5tIfRNpOVYNQNSBAqgCcArl58PX7B1IpGR0VWTZVISn4OzY9v
X8x9eKSU7KzDh5Zk5r1U/bC7f8B8mDwYuCu1sCb0fuSw/oUMAeCTZ0Ib6HPbQrJNx618CTnQZJlS
RXtLmbZXYxqWL5W+WHV7ojjM9176l7wMNQwOOtCaXkUgsEGakZG/zJj6tsHrjxyNXJHEx53QBSIH
rPF/ahv//pjhyiPcR7goJ0in/hM/2AUruyyl+o3p+ku4HmuPesZjIqdu/NjXBTZqTV+52yVLdgR3
JrN9/rPi2aXyHg93Quo3A9bMF+LGW6YWv9SVkQ3LTmvk0lmNQruMGsx9YpKGDZGyRgZQ4eVS13IR
Ch2JtpNRWkMTN5AE00xB0vcLbu5e8rF6i47sMuMRyJW0DazF+3qtybU8S+SJhmAoDuUMxjJyNg7I
JkMSlld3DMX4Qzs6K6B4kYeQkhVEav1CIPi9jwXN/M8NfhF1T2+rTDcg7gVXFcm7qQkTff5TpC67
P+eVCr3gGAOphyyBGYz/sBDaHU1Aobzl4toekG4IJ3npxYUmSgYOskiPC3Yfb2LShbQHwQ1EP4Ju
bTqBa8nTqr5BMPA46/A8bDJ9X4dTKp4pxBcKhU27mmEdUFumUszeB7w4R39Ee33l99g2L2qYZojP
JkAh57wtfhGr/3hZTYiFN62cp76Khs/yXh+Ih3qhAhb1xyez9uUudofwKxdzGYNytQUMYbZjXdJy
HZbwmngbaok+QA3eY52wjsPjWxKDkfags8sn476bHVTCXv257jOBFnz5UXbXgdCcLK+F13n4daZR
KgcjGmXhhiO8qVstOIVCTstwxUUB4mT6EGARpzGSYvOfkSGS5VGoWJkq/iKdQ5P8gmJ/xVkA9CsN
bH7SdTNaKKluc3Lnbevqy6JIF91ctgIZaKJ5viYKwFrLPBXjH+H0R/Z5+zX5it0CDChIx4jBf5cs
1pdMSgSOF7gXeR8UgWxyTRNX8QNxQ3IxWOm7BJT7Q074dbKQNJSkJyyGqFqJAQfHsLITXV+yaZBT
rkhZnz2tFa/AHgFZkf3cM8f4HJSA6IdOtocMAiOaminT2ix/HPHRoG4S3N8C2zsFk2VQV6nmQvbP
1l4rD/SiaITlCu5LQzyc2NbQmfXkjPxyxjaMtMS4LL6dV378Rk6y3uoZ7X9N+Hs6u8OpW2ojLOKx
ePQ1U2qzvYOgB1wYMR5EcmqJ4Zxvj9GjE5IC0Yz+osWsTB69JiQpv6uAVEw/fhku/vUQnliOop8y
pivT2tGP7YmsPXelGmMamizu0wRwkfmRnHuN7kUTRaNC9aWwYif5AjpWC2bxvEwPyar/W93PYfPc
O5f2T23guBI8wDSEkHBQSzks4gVOULypFnDCnana6ZQTV/Ey4GDo/kggx2b3Srvx+ei/dph0U7WM
ulUVK8Z44F59A3U9mXd3ZoptOBMtr1r02pynveQOg0jdFGivRzuEb2jxy4yn1PAarcTxFTw/V0ah
jzuGByDXQGrBI/iHoRUmwBcMfWoE50+UKEqvi1VG3auEFjCpYDs4uaR3lLzVmCcFWGptjPmcXPLp
cz2r8rdBgMmHX07Fs2Mpe8M3oEHwbnZiTTzt63jbpPysV72kl2R0pILsD/xFbkEYnREhC31ioKc6
VHx+eRtsr5qTFR6dtrJMR30avG0XnqMCnMGogoCJAV0WuWFhr1BDf4XyiTM0dph5df3hTp8p14Da
B7C+8zyqksq8WptWoc1kh43pvOajOqzPz7hwaWXQ49+/tR/2ynRUxOFTZ//uJyV4JIBGKEOrNQHS
dSollbSqzEq3R+AZyLAiseSNuy345Glw1cAuEUDSC34zIn7hLyLnHg79Tc79laeKA1f5z8wvvvM7
dINxUBiU/LfCZXN3byLhQO/l789A9vle7Jhl5FZBMRsvFAZU9a2VlhsBh7QyHjNcxTd96l3J5214
SlMBIhLIMwm0KkUSc5cL0H5Z0hlTInfB8ei/0t9NC2pueD2tgYkjx+3vZGaPHt8sFAEkTiSMOx17
GZYrwRvvAqPh1nrvtyuuYGnFlYti6kKlNDcKuGIrEg8wQ4jUhEvcQkW8LDl09xnSxkAdo5sI1ro7
YimzVbxcDz8XZePA495dCW6+xbRYohjkQfwQWoTh4IW2Iwsq9puyehBlN8X4yqZEUrlIEjMm7KbR
6jWy9Yy83NH1eIA6xJlfuIfOFuNosRfJyhNefKYqCbXP36AfK+LWeyqBw/q7pY8bj2G6UuDdC+if
Wnf6FyeEDfd9b3sNihyPLIUpMDvqAl3dsogP+fuV0CYB7qhV5M/OlmG6FMqFpmz/i7V1mcXaD5JW
HOwsQnd9WnwPWMdUuHTIk74WByexQauE1W6xL2rB0S+JEy1BS1CFR/5Gt7gL5rDtSEdRME8ICJSq
Zr2hNzqA79shShTQpRns4s00httrgSF2eccrGRq8o2YuNkeiY3ODQXTIJ2aIwjRAjMo/8/tz/Bv9
QT/aw+/Cl6GuKCvkJm8xqQk5g56AEam0jfkUrTCqSZaiNrNhhPDYay9zhaRlIzQYhiUhRo6BVDdh
DPz+bRWVFZBqWJMxQ3KdGJexpjSr8vsj1anRh2E7JFYBvgSjw3X+i998+PqcPXcGBB2K9JBzxPH+
3/u3jdXs5JgYPl/WZv65y1XLxu32HEzQWb4w4ZkOuRMbIm9p9exQ/8XM1aZMncUy004U9GMBJQRS
Iyq2HYh/b0EY/sWnoewnB9f+sdll9k7GgPdqhwDPQ+6c9LMQzdXbEwh1sa296/wBvvaTXLl2adMS
TF6zrlKb6GigAItlJ5V8WKAjKGY5x54gvVxLqpA4lQYlioZW3o4WPI7Usn9kfqz2lJeSasxewNIu
EBfoMlveYhOhNRvulxlz2vuogAljpv8oBKD+iVZwerSLj8+/TYI/PUN3LlKNz3BHHPfHZjLL2zU5
rP/JlGhTXpMF7qg0Iy2lOdM+NVvv6w8VNPH4dzJTXOFjxfP5dAwOzKdAxTSXNevIp0hX2IXBrtM3
GSyt7dG7PasfUWBgVWmnQGY/DJWgrjK1LZ8OUFp5tjC5QXP8FlDAlJYeu0Ob0Wox4qMQue/6Hy0J
73k5y6dD3p8CsqvompB39dGNgzafXJSYMudYTavk/HgB1KJ5szxOO5RLMmghLag0/j5lBuuFrwuu
qQX0zU+2UUQEbp6Xv1uZsEP8u55dwEK4L2lGLWLMK5tCnXchyVPk2EJUAz///gZoQhOh++Os8AcS
GTUfngw2yDxU24oEcrh82I9DowrM6mJM6SldqWhd4nBQlf9xjxEjKzYkn3rmnYXb4bfCtNnaG3YU
NYwESYD+s+qJt691jmqKV62fTVNA21Hsnmgq/2gzNySghW/pUH1Uujf7+oHXabhafDWISkSc/Vvz
QcQiH5bRuSNjb+/aefXvhvDSe0mmyRbXK1vwMF7EjWIC7vEZavc4JF5zblnuBBriGty6IWmcBGYs
36cpEe76CFbZS88v1PtQwWV55r444MoL2UZyEaoCuEXT6fN78g23Rn7y2wptagWObFJrEJBMrxFM
ZI8Q07pbP2771jrXjC/F+UiO8NsU1+jreSV7UkO2t1dm4dJzDIzNzr7cJjyKQVKc8ch6YhuacEnk
gwO0CDU1vyu3tJPA31FO2hgbMZjIwG5e6MAUjF23ne6eRtoCes7JGYrs/L9rEVjuTu1Eqe8XNAiP
1B2ODXd3oZB8z0NjJJkfjqSdN/60z+/5K2v5ad71vPTxDOzPiv8zYk5tAWSrXzSfvlFRqfsI5Ac8
4zMLpsfKqq7/PhxD+azozfGUGkCBGVy4DDgrivEjToKDpISzGUusuM7cpF8tXGjc+584C62b7ZKm
JhzanH3pBCd5P9Y/mUcbOOL+MlenQUuvH79JxN0KgO0TA6BS7lCZb5PNh3PTwZLAXClk8baY+w1b
E5KjjzGXFOXnbjFN870MdP84Ykq56NDsvjDpUysZz1XRawxByBpDmRHbhtWEnCixcoUka17rU9Sw
31dckImGfz/ACE0VoEGYc+JMGMjhRzIHnm20hLUsXBd0CPKrcM2YqYJEP9PwWkNVI6RCUq8gVd4v
N9jH1I0UGdfhn5JGEE3a3tHQM3OKtm48AEcUvzJF+3c4gmxMhZL9VKryt/UjZpYX8RoYLGvNIfge
36dE47RT0WAQ9eYTUovAZ2JPoPFS+LYKJPXuSFO/ktNbBqqiFXQgwKdP2lT2I8kK9hzSqtW60902
WfFPiOsrgvZrbjhZ9Hebw8ONW8yckwJTCjXe887TDqbUAfqGqJyF8sHhQ2TyNXf/cX6ApIKYakSt
j6d4UjqcF7GWo3uF5dkZ1CjlkXhmf9OOrEM8P8qTr51GCn4zKBbbNtjI8YnOJ3mxmWoTPMhLrb8X
tFMLKUBqFxbtsOfok+DFsXxqY/MCMKtjaA37z2R6oXp6huuE8zahmVdptpiC3kmEEPvmzb/mteZU
uyk6MneIn+4lUzZcPUhA+AAFrNUSlIoCFPzRJJlcxdMuvPAXSDDHvp6w+pzbvguuEx1ZagKQHBlv
XQdV2umA+I2H8KPYVpFCGTPGsDhhdZRc0cqkM8onlz79tS8RayA1On6Lop8KGRaHIyVuieHEdmEW
N/iBTULvEJ70VTBCtYvF5S+8ylZ1/XsS2x2T0iLbqygxWMwsRSKQ8YCdYZO3E9x6YxebkoF9hvJH
TZqXAk7qzVUL59VqD8U5GyFwyrX0xILrZm+MJ4fHd0y+ShIJQYbEGzPd0s1NKimlq92I2RZMEf3z
sFZwgWnS3oMvgOmJ/em3g90oWCqrQYGoUDlbACQGo7Ayfw59EQUz38zskryUFhhZa0Bj0/KhgBTJ
smgpUvHAcV7WrygNMGH6qOcvF5g5isGX+SpvCULU4hkFqKhTRaH7Vi/kJ91+MU2oU9uSxiotoOHu
ldBuCuo41yQJSQRK57hhU3PWU+4jNizzo+nLaWh6ZFN8B5hVdQNBbR8i3fDdZteP+OnzDEwWoalJ
PjlczXRo/R6TgSsl5wkmF/gPt+2nfKg9+CDLZo/oJvUek+V9OSRs23argw5suupSsEc9MPTnMzH0
lhoa/zDrcVNCT23NDbQB7a/tJUAz9TKUOt62rbXZMIm3rBjLLqPHX7lgcc6HNFcXcxHcj+qjvYSr
AyPRkavqIVmZcfzoDVGrZg6wpx3D1+uTIegsDdJXm4qKG8Vw8ihAhd9LxdDszvkEkPcSc8VgyGcz
uLXN9HsACTzFfSFg9pxyWlvumo5nBQAMM5CjkMnA170FPW2T7LhQ4sjGvIrJP4D+kIorfkuGBx3O
ZGr7dea7HAKfQlWDrpg5XI55jMmRF8MvXAqZBfL3RmDjYaKl0hwlssoXIOnQMotD37lkMjcYbOKe
A3h3ptWrmHxfnEijIiUkWiwBCIpdYjEyWS+o8nr2haM/q68Smz7KeYxEg2fCHNL2WHwfaPR53/cn
WTXW60Xv0LaPNJI5oqknGGvU/83kgxVyU81Rxb1MX4XKhCfhmZUoaO1kBBkFvGNjE1uUZzZeVAml
hjVQBxyIa4NyJu/xJDHx5XcmZTilDg3IB7Qc2DOfUUJVR4yt5pHi8zm4F/Cmu8x7qUjiLN07DmQM
OXg/XcxaI2A98ukX+b+HP1KMQPremPqmNohg/3qxwsaP3C+Zik34bzkkKKb/5C0td1MxFCylJ05R
ZrmwSi93jew7CbKwgLrImAjtr7LV1Qe5irkIj7PUPTZPQN3tTzMnEdDzh1dwlFg1Ny1RwPr7zGVo
j9xy8SmsrFs1cmtnPKq88OdyrQxXfTDXgO2L6bt2v4k5D8A83a4DGWTOf022W/yDgeXQH1IienFI
s3eKqLhjOSvc6hOmCU4qWLXJiGzx2CgVV7RbPVdapUlRjuRP2IvmI5YPDWn4Y/LgbChnX6f1XFUw
61efhoCJwyA6XVIt8rBQVM0HcET44df3utu8YZu/sSjm/7kE3HdpDSsamgZRr504KhumUnyT1OPT
tuWZ/w+rsnKeqiDy1wm6JYr7Q3+uU6bVxUk0XidBZD0KUtm3pETtogpO0/SjRKbs1do5vAlVa3t6
JvPrGCgoPclUdC1sTlYDyZyRLXCglmj+fhwIVw7II0ec76Mx7IzJhOLd49FFh7I7bqYtzXW0iB4r
GhHQjEBBH03vqlRp5izdr4dsvGlPvVZheOFNwwsj6CQNjKDIj0f1HT/a+jTJzU+7MoG6XO95iTZ/
pN5C/qzbW2/h1fb+jxLtdV7WDWC+cmVcszu0Ld+7JZcHFij2mxA5tt8/3W67EGMolnL1QlRMw8fG
N5d0sFt2RFW/bVu3nOAftElGUposm/KX9raMxIjPF58StTmBVlTMr6IEzTlGdQ0cJtLb49EcifiF
Uc+3QQmPHx3cKi4awPHErzu4RhIvQ3f8ouYyxKD0rutDl7/c2wpJ04odSI9hxWYopg3JV071rbVo
qjtwtDFRrHwW7OzfTyNDA6GfaNkpdhrmM4Zs3rVxQagPdcEH3OuL4BpA+FGk77P6VW4iW6bVeOaq
tqLRj//3tZU9bp94Z5swkzif6VXJRvqJ0mnfeHbBR55Ls2K0Zi6eyLmNtjlN2wnaiWc47lTI5oBA
z95iQenWaDSZS/BQDpywAbXot4dfuogzHk8Wv2ejKO+oOsizQaT+feH8iSR3rcF+buFMJ/cEx0GI
jS9Yy69ks2An2S6+bLjQBUX7HSwbBcdmW/5L8R+nxg5IibtPM5/TBF+TgVbppp+WbqJNL8Z3g0RS
Pqzr41xxXAwusr/aaTimRNvQTaG/TEJDV+QI+WkHmhs9YwKjGFY/StFhv062+tPKZQ5ZGDD7Cskl
Svp2Kw+EWNGP15Rx3UgUvS0Ih6RucQjXdmyPkBAML7tBPO551DEpHUb5Zvn7PxFfPpKG5FpZsPYU
EQ6ddSvpf4ck3cduTSl/IFcOEVKW0CYK0PJTxLt9buM275bTqb3gRKGTHNkPdsnbHlJcOMMlGbzr
DxA0QT7Cc8h5STX9EbKhwlqeaP0m7O2J4iS01RzqYhLBXjm9V3S10yyK43bodjN8cnpSVgfpUDDU
CGeGP5EBWDrPiSyS3i5dGwAs6Euie/m1HYYq3g13ESYCl3suPGHdHe5w6ytlxMxntDJcdjl/OaC5
mFfiYNagwegesRWu20zCSUfkN5TFTi66Ufy2nNd+Lq7j+f/kNM6/S9qBfmlH6w8HH3lrNSrSdwyY
gaMQwOoLDetqg+K7+flYMH3DiQ5yEfq6990Ty7TJ59P34sTy39bYRVjH8kjwhYQsh+bT/99Gsqjd
YTT6VbGzXpvK2YwnVbtroMuzh8GjbmDDr2268vQNivMRh3kRj5CpRitK7Ofr4hLCFRxl+ARY3rKU
cqYC+8PwqzT7c0qmcgLr4SElYq5wt9fiGzZQTUN6c+GtkFb/3Xj9ItYILC+bWJC54uHnuJzZ/mkf
FHjCo1gbE9vEOX04vzYVMeo0AxB63w9sBqZxDd+wgd8yyH57UnxWR+qshm60HmAVvK6X8iyOYaBw
yzmOLlQLY0iQvXvxU/TjF+fqDOQDYueVJwl2m5lOzS7/8cumO14YnRU6QBDdm86aMrZ52v9Z27HI
wpqI/jJ0PREo2WZboWyKY09vSKCfaLx7Uzk86fLR7OL/MNVP3V/SzX9xWtOSDsj38ZTSJHgQldQh
K0KPwp+jYeDbe4S/JlicidZdKq01ZtrhcPl9iDEY3V6R8mTnz0Y6ToUkk6eTukNmgXtmiw2bED/F
w3DtR2yzUk3LJPnCu6J8SPI//8aKN9gCkIG3piPecnmVfbPsZPJWwaV1UjJ5fI8I7Pbwj0iW9sHk
Nk+EhOuPBKafTam46ZvI8Jq2bCSbgMG6vTzNALORZ2qTy/n4FHSVagMxE1PVMKSBGwt4SP3Bw7Rk
6F6qO38O26prvVCSSwGTtlSC3VXnIHRXkE+gN2DnYRoYm5LnM3H6xSFdbSKpFd8gtImo1/F0wX8A
hW7xU9J/+5A4xDAxqS+Z2rg6WgA5NAQV0tTT8anhkmmvSgl5PkEXc1XCdaUcIl8kWVwMuOs7caHC
kcUtU6TqRTBO4/Cez3JPAME5YOFsFCWDV4YpM0ylkm4SYzgH7X5blpBJa4xQseg3hGhIvmJ9cl0S
DO2igdGEIvGiLxo7Vy6T+QNFoSBX6/K4wY9ng15p04fnGg3o4dmI9/tcP2Lqzs+HWDlkK2/GPQvA
nMuMNW+55I58SFfrycvB32sQ1uW6lch+uW8WiRnAUU3nXzP1C1WakBWl08d72XoTBbrJCqBCDrVQ
RgATITpx+/ENPVHKF9bzBzKZcnZnc+0MOvYUWQh0yFQqR+KmBStKhoBJdDCMB/NAQlx26eY+UYxS
3zuJEOio8a0FUd3SGzouCYdD1G/nFiX/hGPHuqVJyGC1hFOK6MghD50nJMCrNlxtz8LHRgs1LX6n
f+P12kJnG00VwBGR0s1bYV/3TSGOd2mbviecfNhyiM353Thjwhy3aUGx5vsPjUoYVEQkofFyO7yS
yHBqoNGFMBv190+1Uy/rEqVNQTnnaQ/lXq+XzOkl4SEN+4A7YMjwfK0kAL4ZIbbDYloN+T/JbO9f
09qVfcs2lSzzREEn0fRm7Prx4qzNAWoR4V8LJIxHP1AvlLXIUxVkFYjBqaZxImPnNRJynb9uM9To
gvg/ldb9AfNcsx6sPYygMSzT+gWXj8lPQ6Rp1fPkalkzKha3j62AnlXWLp/ocxrSlx8E4CJzOQV8
QH8p68rLD63pT0up0pM4PGNXydoN9omKS6EPqFRCUOz/3mpP4GSRmwULorcjDR5IMirMXi0vBXWV
fCpkK3uF2BYuNLhyZYaCaHN6j417buyNdXhtrP/1CuP8gGLfXNAVRViVIbxOrDJrSFsj5/n8PlcS
UhETbopNir+oNhoHvDgNT2mZQKpbQ7bZpwaqnD/W/rifk1ZHIQ+rmqQRW7q0qFhiWOtlIf9oeT+r
Fm6CS7bgDGqHFAJpHU/0aIEGyPFO9yQhaVL4h29FsIGMQdKTrdeSreTLuLa1dDB2VEuAw9MttGu3
IwnM8CaeSvriuLjr7HySDDmDdxLKDs5/erbBjkRB4LJKu+mbZNhJ0GZnpoTnK3TcDNLLfHeLjsyZ
8odhXGBYTPCqEelczRP5xLj/cigHM+MCihUdUj4JY2EiTBuLU4ABKJKKJzCSBHIeWx7Oo393m9+T
ZhTt7ZitFs05Ea2mIEQ+zILod8Wga7NOM3xozCxY/6Qv+4AiyDI5vMNsGiKkxpdqg9NrD8T0wHlw
u0hnWITk3KGHRMg2Dg/Ye9btxPLp0gI0Bqug2EEdOGvQkdFcAHzk/eG/on2Kc+nuW5ZFde45CEKu
62KTHU980rjsL61tXdKxVXjxdAzVWT3/vPF+VS/0E44nlHXlm2K5O2jb4kyZe6PqO6e8PHObwlMH
IUwStOY2zumyIdhOc1923/Pgmp/2V4X0iOxCmbi+HaUPA7VvOj7sF+BqnwH++uTbJiDK7lyV/8bn
Z3oIyv9bMigMBx3DfZfbGNBWEC1g29GflfdbNg+YTu+IcQu7aXbQoY4EwBf4E89PF+R08ACRBTKg
L61QxmsKwhk5T8tFBvy/KiYdfA1zHivb8u38UZmIIHG4dIzE1S1KOvl2+mnE5OO6a4smb1w5Svcr
SVkVT9bCEm8GlqQYgao2WRpd8UdbrXVwGfWs1znqg4XL2i66xRLNzoKBUWO/remhQPoM+qaoWqlU
B3rqJepWyV2zQhzmdlqy5TXM6Gd3Sh199dJmwpbCffSxUgS8INVm6pti4TYXzjfGApsgErFpuNbr
jh26nER8LR/PDaPlACCg9yx594z0uCNZrT96uJD/c9SH+O/bENUds9iov4S51/hmj/8uU77h0DUZ
yL1tpaHoeBaY9eseE1t0LbVV7z79mtRMzqPyfaTvmBuc7rSVZYZn94wyx4ibCFpXJr8dHA1i2UKJ
aaLyVsxjzU1DgM5gTPojuCQHM8VU7owVpqCMEOmxvi/hI4ZeUXV7zVNp2EaBTqt7GnzYEciwNrZc
T/a3TvUTsrhGp6ML+1Y+wR4X4+eM/hCnd2YDcC+bL67DuhJxdWOW+4bFjwUifdOWKgH7z1ecdEwW
WOK6ohppAhdq8xS6VdvZQFlb6MYCb1px/nR/9/i5x/mzgAbFVdoQHz81YOrMsFrst22KujSVsMZ6
hD1cSmx147RAIgYlEPBmAHrxMzINdi+wrMs199Ibr1yb6s2UXUFzRkYeSBfyEmmrSDAO27um9wT1
GZWiTJAnGwQyzaYyodUUGGI/NAH7Wam7Y41VeTHRXNmcs1Pfj1+0O3M4lGOnRzMmPDGh3nlX8EpC
ijD4rUgdrmc+MN9nV7KZy9Wd8KpjOQ2NAZAKEXvJuwp0sP2yk8EXJgjk8q6mmqxRk/VftrDRZEy3
igtboM5ruiFelVA6LdtR/3k6CD+ody/72xFPwtEF05NF2HIpLLOs+rLPm78i3SKyiLu1qi3fKCH5
+fsOLYCD0C+Of1BgM6eZ4NGJF8HRCegeH5NwS/QgMxQWKnr8V29/ngihEmyZcSdq+U9aaI1X+LSg
e69KstmmR9kuB9abun5iIXAbvA3y9XlHtmocJ3w0gOBfimgChi17Z7kShsnQRUnSjQQzLz7sq+zj
po2ZemsIFvuc1p6iRIqQPI3/iYhj7zqg7kgMBV89NbcMhChHbvPv+LPmHKISbSWCVxR9l/zG3zpQ
TJmVWxXPFnV/8CxNDNiEACabikMVO74YhQCRzXOJgbKMuJyK5P5J/Ywu7/2dQiu8O/PaofztYMpi
sXHkY02+gUwgrP49YVzgC+Ee0aFc5ZB7zXQAHjP+LRuEEsBBy8fPG6BsY6mHgBG6z0JGfTi3Ig3F
SyOOH0zi6qZoVv5Pd4iSdvohhlxVVYqPFatOb0uCTPAiniI2SbuG1CZjXt2XU4JDUlO3xRrmvM1i
zhTlLSmLK74HS1rfK+0J9vViFXd9JFOahw88o6VGGmBTgjg+FVBZr1TJDq3IEkA0osWo6Ne5DKBa
upWrU+6Sqio0YxulvcEAaPHIK+S5hW+ecIhTCOx9/dsdBb2SmRUTrhE1B7KmpRWqPympRfAnnzkP
Xj2BfIUzxDdRi3zoekzcEoQfv6R2uVg8bInjKgJ5ElHjGdQEQWbQvc12qmfbXL3/Yin3ENxcUWt7
01M3VEj8Tca2O9h4Oy3zW8V+uphjYzoa7ls4TiDrY8fFNYzBZXbUcWBN8d7WZWtmgYecfHic9j+a
24LT1rsNJKXqCRBCVHqbyAjlNrmHJZdirVWCz3UkKCjh2S1qeDwl1ck5405/WeSUqmD2UUz42/Mx
mM4AIBt9zEUuUXp2k5ZayeUNl32mEgwzSAnVvw//aXg1qLTQx2MIaCe/mNTNfQr7w0ehieHN9kUx
hbY60Zj9Mvbm/c8IBEh7ElSeKP+wCmzzR1eSO7vz3DZefUBuqdBuKvp3x1bR8OP08WsPmMrYdbRb
JbZmURyqBGTVIjqK4OpgEA0S4FWOYLV69YggwPO5gGjDklzpKu4syZTthOtO0RQnpB+drMpDTFVS
1JFRcWoROjYCRMWdZoISc9u3epVoujGRVocKJCii04qF8ttEKM0SY1nfIeAd7V18zMhkcQ+qo34q
0zeL4h4F8uefQ+BYNKbYhh4T29y/Dcmz30Gmp+xnPGGqcUQwvTUkPhn/nltuwO8z09plIRQenFvN
4LyXXiMWHTBee1SS+yDOkzefXBPOxXpsgPglQ8eC8maO+HgonyHb+5ksbIyTdgS7G1aje4Z+z0oq
yyqf5wAsHN+jO2AOYM6HjZUgbWZ253C/KSf5jjCKMNNG0fxwWnCTCS/zzAl1i0C9d22dRp4G4VPf
S8Bop1qqG8yRMwvffsmk9U25jG+y9IVbkLVbDHFNAuV5Jpz2BpfrxcWV8VESyK0I3lMMGYM3hb2k
SgtQOyBRfvdUItkPquF9bAmEXSC3KgWkINGat38C4vywJ2ksmEQp0DU5rtoPhOVaAKxmWZNkbhHA
9vto8VJc4Mo3Z/NzrmZ044sVvz7VXglN88aw0k4KWKtksALLvd8UUhnXjxB0RuPmobXtTYy/R3FA
BrCE650OYQZUgDfWDHt20dkZcxkm6hPO9EdeANfOykT2EkNS4l66/iu0f37L0aif90pfxMUroBEX
92MVhcAUaZKQfY1r3eIRPOVsNAsDw/mq9F9QoeVo7a1nkQ3dM/yWSV4gV1qpkx+3xR6lPNGGUA6G
K6Ln1KGjKvNcw9JdaXS10rqAQUlgUJ/f1O9b1odW/Kmn3Zi0qrzcIYDXlGCkpCb/ZYAB4Jlh0Z1B
KGsjTt1dN1ZN42EGGvlVATNyYCYlubV8ZQojuqWF5vS9p3whFmpMrz1x3DMDPIg5YXnDjVPxW85M
V6qow+mwoOBLQ3M9AtidcpAOQSiCVnwEKLOJ+pilrXRrYq/9fioYTRLrwf5q97NVbAqm0Ugr/pvG
h4MoaWHnXXxa0bIy+EJDzw84UwKZx284ACqH53enyWWqHw00cmJdB6lrmbisFxholu7m4BjB3PZW
b1Q0uD/hrgFi2o4ixHArk2XZ5MEimP2iAvpUQC2p6b/4TmZXYGs+A3+yHzu6rPomLlmYqu7dCd73
qVzJHyaBPJW9q5t6OOBx37ZMIM8RH6Wfw0eDrqlUEHl4Nej53EObMKiYFhZ8UwaXeFekSRMTu8sO
zLjnzvOr8evilNdsyX57G6v5ikJsy/rAP06GIxLEfPz5Sj1k2qn3DxHFqqiAnCA9i2QuIi+i677j
BCaTOiN8obz5xDcZJth+dkE5AKRsfj39J2+lmDQ18xgoBrQ6sfKmdDieIAlE1pJmd32DN7qNJ5v2
AWii4qNTjSKeFbA0azCGRWJSZzPuE1Pl0KXsf6PaRYFuN196pu5NB/heo8GR1R5ThHR0WDjmSOu7
Yx2fn6B4CmQKqRlvbcijsGs/J+vH4WIwlD5g1NzFnrTgA25dQfmOvuJBokDrpLg6+X1/5x+hEFBB
umLNU6E76YHmZxmTjYr75Ob+bYeNEcgJ2ytv5TQKu5JD1C6rfx/CCW1FOtecP/jtKbgDSEDH/afR
aZGVKE+EoRyugUpxz4Ln05+kBhemdb1qTgDQaby7Ntb4wzvJQbl8Nb3n1jpkeUuuQRFnCyRy3jFX
1itL9s7T735N4ahPvEQTF6A0fqfxRdNTB1RBT8zQb51fGURoPXqswNJ1+FIf+cE5bJUlbBmX8yQa
fYyZlzvUgfiyV6bN89N4b5GlA9/DT4iWGu+odxeoqGKQ3JQDW4hLaXGveCIMUuwoaQu5YlYnMUhi
vBAfrBUFwEe5YbCfk7zRJprPYkrubijdn+2NHfc5fSP+H3+4BbdCFcl7DSalVkqgu3quNyQLnPju
XDrWG3AhMo0QWM4C+S36w2kwYCwR0QTl1jnlnxJxgMhdCOHIEoK5wI/t4FquhJ+ve/MzjmK2C3yO
RKEbHE7syKsOyQXI5MrTB87cIl0jWm7KYlf2RUIK8zI4RxX4l5nKqjMt56OGv3EBr6CaZqK61fZk
ldwUt/9uU+K+cteWMtBu5MhSbejLUOxjBBQEtV/RVCRLWr6PIiJAi+6QXGm5I62E5wu1Ex+qdWkx
AmKOS86crTimrsZB0XtqUd58fq/2ajLUtlh87GsujFEhkV0G+PGNED1f7arvtyGfleNmirjoIb5w
F5PSS20JLZ4OW3J+JCqW22agLqB6QKYzoRhr6y2w8w5AeRc6ah0ODh4ge5EOLrqe5LmozPRwGXWG
ku4u/FnWO1eqHw1QvjSWMIWrxexLDUl0JXDIDBgBRoU/vmyU0aJbZvXqweVOUPtA/kY9MnVzN1Kw
D02NT8JPh8KIbHbvJL/qTMg68mQr8AU+4aJTKq9u6wHv1/UGBi0JvM+cGeK56a38K2W13Sxe2IdG
veW+2ejsl0Xceu8UWKW5xhjhRyvkJcpZlyi4iyNYlaPkgMTW1AO4yLUr850gh2cmXa09DQq/RuLw
52KiC7KatqpwnTWBqtxv8OtUrghJ7UU5uKOOPrp4+wzBiZQ0v6ECgYe6dkqpgh4XqLTzzzohqZ6C
X3giON/yKa4K33s9p+/fHh21XgElIKND9yuS7QzSIU6PnHqBs7eFsScVsUrH41d+ATj78V76IF+R
1lSekvliX7Eeq/+1R4RXFaOm6YI/p6KZ3unJIMrg22TaruxeMeuOQa1LI9BKGGGao+HJL5ShEZia
qF3IMtRG662MWz0lrPLX5YMDPwLX4ArV0T+VxasAfXXSeJr2o4rTNszdJpeOHuBRxTAq7eWylVCd
/YgM7A9yBFWNwR2eQNrx/Pol8JzqsnVJGXXqDNjf7e+2TueSYde7j87f64NmiX6KcY89mpJSTviE
FdkEjEoyOd0wIbARKKOWW+rCL4fhRUL8YcSMMN205xIhuouPz8hTCl5U1HMpx1w8Im8EOLRV7O4X
54yuAO6ulR4Rz9QGMbPQtCf5QrezxjpqoGwsPzZvVBHVAP0WHZodu17/WTdkTHad5HmZsOay/WIU
GhtqGLvlKyZQTTiZoDlIN0GS2Vy1rZ7nVsuSlOfMKka1xIxCVC0qaQWs7tn3By8opSPjMAtYDWe/
1n38YjsetkcokIN0dc5GwxEDnvpjD8BpE5i0xeuK5cXnxwK/Ofn3/MHpCx77GZW+mazelVOAb2gg
sIgRUZhkMykDUXLL8hLunayrxmaloaJHX3ySRM4zjU/JfY9UJX9IhdYC4iqO1PMaCb1Rdy3YbGrz
YrKPBMgqjMGgBtsENZ+JAi4wo083GkY/k7RvzfII9pxK/qmcblnbkA91Ti7U5wh/+QEE5TmKPFry
/Gz1NfD/qiT7+eKlpwG8lzpKsaC2PA7L8Rqym8y+T5RNduM0kYX+wCT1L4q1h3INZrmpY7ruMWGE
Yx9c5b5QvwE0OBnwdLDDlVc0AjY1WJ8dc2ISCNFjWr5TL8ePfXdSc6xonHHC9sQb0Hm1PQKRtcww
XlQM/9+LV+fzm51O1O+aXUyFtOCuU3v5JmwHN9lYa/VOHC/EgMICDdTAvOB+Zf5ft4+It70+nIhY
Phrdu4gBL3IYcYyCqQ99DT92LO9PzkCzu5xZ9kX8xrSQQJp45Czp4hVr1fWhQN4vhwh5L/VtZ4Fo
h5RhVKM8bffLX1PTMf8A0fcphwXBwDI9kuQfg9+qurpEWZRAbsD6Rjh9nFF2FzfgpAJYGmcpA2hB
Gwvc+gkEveSEYnEJTo9350yOxAu16ugzhK8sy0nz2mSGwY7+7MqxdJDkVveVhCoBiBtOikim97X+
7a/LrVRrY+EU1+nizBR0qxs5I2cAy1z1JIAaTZ+wcVmwH0UVGa4L8AEmHswCEzmY6xsuRkQBTfkL
Q3D8J36OXmzPjJUkumtz/42kjBvvdMM9wobBkmCY6zfwdNx+ksx5Q2vAakL3mJPPeoYJ8Xxwjl8w
sIgK+j+KM3mOAV4VMUBNohghiL2XCkjWy7rE1LqYq7ryR6hW/npzmYVvmSp372a3jkvoo4hSPmUX
netG7veKSfnCOoIwcYWD5RQtExe/ngSvKtXhDPjquv+d0UjDIWEkxC0s4+ACUMbtJiEk2R+D4W/o
UFNXjUBLCO272vRrdDn6ZHGERUWzdb/07c/AllvDRAKwQmofGRAwH+3VmOT4aWDbA3i/uVCJc5dI
I5KFGEG4pWxDPWExLU+IivNY/O8kOuSD5VBeNIYfOwqbmGapLVHINTA/o92vXDLO6UjYEKgoztVk
hVdXWB6dAeWCSWQJ0dCXbk7ORKtXOcjzuqMbobI0CmPp10Afmzl3s+Nn24p7gqOMwOb4MA1Hm4y3
FaY6wIhcTqf9eMvHsnlXOyUla7g2cyaXYLv/Hpojt3yhF9T5ZtXNMpWZ9USXILKeT1cMexfM56gW
hILxIkoZsrLYTX9Bn2TcmpPHROyl7DbiXXqXq4nGDWHwbyDjV2AvOfu9UfrDESS/EvOPW+0w0zi2
uNhnYfG1bQsiDKKqkZgEpLaLzj/bDZ881+Fy9r7nmAtHEPRzFAZLPMkGnvzPzwoKaQB36Fx5O1Ey
6S+72ZaOt8Bqd+zA2nFmu9YrWVcY7EmkNfh4GWan+cxF5U/3BpaiNbdpMDv/EmANodEsQolDxSwJ
3cHMdBLxuah9/eBSjnBQ/kdcVSXEJuG3ZdjSiIQsg+yNtkbg0PXmCuK/iNGcxQZ7krCgcF6tRqKe
VGYij1Cjc3c3klPzCmPWXfEJwl9rMAw4PariDVwxMtAZT/eaHMYx+jT2+UNUNlB3uvZEvHSke0fL
szW9bNXlli7/cxgeHraSzsMNBwVj2HjIguzhAW2KMc6J+DrO4Rmb4pcIf2JFFPIwfOrU7EKuCz+L
+ufvOm7JJNd5qNrvEVCro2ARmcHOhaSUUtQpYhi4DCip0crd1bgrO2pXcUYPbk7VT3gaHoa4nlYP
bBzVuTjqDzvfBuIEwL3YsUgM3BjC58aZBStK0aUvck6ygutJx3tgl9D4xnIuIuWiqi+HMQtvckfS
lRMsAlUEguWLSCuZYJFe4KdohKaADy6oI7YfX6Wyy/M4lxFM8G/3K+VkJ0VNvdO0AFbxpSgZfbPn
GgFRMCbjkELEzRWuZkXyf57+fVj3MnaJ5Yhienzd9kZ1xhiO0wcVST/JU6x7VWbhuJ4Ds+P8Lg9V
m/LhP1KiXD1gf6Y1tsP/aMDQEHudwIivw4jZM9fvt/kQ8hJRHmwXbiTkqUbSCmrquJ7nGxQG4AOE
S4d7Q1YkbdHwa/bjys2O7kd+eZprUUsaVjGZwPqQhwiVvKRq91zJNMchxq9mJBOh2Lx3cDDj6qCT
8N0Eren6ULxSUC04G6LIOv1adUHsBc4QIavWcqb3k7QSEIlMa5q1dr8OdiHUT9NERRZrOPC9bWR4
hK3cXpHzoll9oMKjg6jWA9wPhdJVg1q1M4CXKvR/nKnu9IomIphnLSF9Rn6HSRJoqyXyAsQe+oab
nieeEPL1XH4zLw66h6nYrmA2wYGwjFv7FQE9bfOGWQwjkgTAXqyEZ3imaEUGoOMNCzAtCuHmfDS8
T140ZyygpxE9IKNDm+Fvy6iNRA50yG761WUFrhCJwOTo99P/LNiYFHUqwKpr0TI36x1Zq3mJRecU
7FFVbIO/upPDVEC8HLpSL9PvkITznpnO+BA5GEE/Cfsbm+QNI4EAn/7KFpP/ChLU2likj+mmsBLo
BMcgoaBR4ZPfBAjQalnhCpfZBDttGirez5wWKlbx0jqD25HH3pyeaYCFGmEVvwc4jZa2np9DrXUT
gsNjevfkDj4KPGis6gUYY3Eq8uYkYascJa6ZeIC652tPePmx96cWcyhi/whnwMiywzGLSp4zMtru
kmOSeHDqfXEmfezLa2aaV6bz6FakEEHhYdn2EdH8sQkhKZexqTbOGx91rw3DLiNixBH07Kf25Z03
3mUhc7gNTrNrdsqrBQRfsiKPtShzQhueAVL8IgqjZ+gu/HOGIzktjqPD/hVP/gq0yDubQR9DyV7b
VABQlcqQP4fCc/EYs2LvMMDqL2ImhL1VU/5dgm+ULjjVjgylXX4qh2t2wKFTI99Blu7OxoxzxGI7
HiCuZA/NscMErWPof84Fr5y+OuU+C5zsChNFlOFQS5plk5k8ZmaYoS1ro0QKE0PHmhKfGf6tV+SN
aQIwE/bkB9D8tieGRz3GjKXtWg9dVfXA7g6HGZHq34XjWSdXkE4Hwa1i4Zrbn9w6MbIP+CIZuRRD
KPSiNofY4xtn/mkzf+YLsXQoP/YIjKsWnJsdTKkS1VOsygzS08yu+OT/8kVFfwAJEdwa6WVFRksn
pKlRyLM4/SHgX6uRL4Qi2aC5zvvsqdLDPK1Qm9WM95KJ3v/c+pf0lKbguvPuFE5ZTVcr8s/UINy8
kBYdm+AMPgssgLB51aYeDlsaEJK2Gi4a0AQjgibNVyhoaYoMFDhm8IF0q9kQF1k6uKEEgc6+mHdI
X/z5kaYEhOQFqvJeGOURFf9K8GUouvQ+W2/O46bDetgeepwCLLQolULNTHI49qdoVqLTJC3RrjQM
i3ZXVEvhspfRb62TPMhqXbxvQNppKAOIerQ461vNqHfSi/TyI4zI01Sn2FOtdl86hEczX0AmzksI
S7g06qvUIc3aBdYwopHZ0GF00YYfQR/70qwlzGJ8TaSN+rAyhx1grmknXvCR4YHpRCSfcxuzkoU5
oosYoDJxgqPo47cpzqAAgG7NBrrzEm9ASnUvEpDUJd4IYVCiaV+sSYgyXYDJvnZbZt04ql57/KGj
m/LxQAR3QYrc2Wn3/oyNCchiMNnNHxApkwwHV/2e3Zrg0n0fS/jNinwKjBQf65lsgpiO6fcIJZEg
fohVNEholEQ2kSEg9fOobt4GRXkMiR4Dddxekih3gDfTgxhUhd4CZ78ZOcHGjNJpIJyn9hzmLB4Z
o2CR2uZYBJFQWkkwFoO4qpA+NziV6xmSujzZwIW2/0BsS/5lKWyPakgFWAq64w7BhzG00FKw1KnI
cyfVdLJepmPwf2K92pwEr23lLTyfbJFRju4J+ccRbi/NKW5EMTXJN9PjAMRoLrsWXtax4izC3k7z
500kN1E1IfCS7cWNlIdOz+KQhExRRME94z7fcGScG1ktyyKbxk5o+FQZ0Qk1UqJwsRDS7QXMAUFR
J5puLvGdx6XAfFSl+PVgc7qzdkCI/w3TbLoBZXzpTIxVi1lcH99BYYUetTQrfrZzwrBS8EFpJGCn
2b8Lr9dEPZmqswUvUe8NInsDaViNHjdfuWqrlMsmDtCFiqSXxh6uoCepfx5orhBVPTg6FkLN7ur0
zcuh6FdaAMo6qsLSP8GAUcBNvZOErV0+ddAyPRv+OfSd6ABUtOyJjbqG5qxmumGFsiderdne+Tuj
Mym5moVLWbEhMzfZIhKA9wqn50M9q5ZWKOkkCxZvUSYeG4LfcvRQP985MENYC/zVXsLru6jja5b6
U2Z8io0YMym/3swfut3cgNUVBL4TSNmAQyBlLBr+E6ssm7mA9AUKo92+OyXvlTocfg5HJrklK0FS
9UutbTRHnpIRpIfUbS/54rDfNhKi9/d4JZV3Qvqdm523jYW4Cur7e5LGYP3/sC6oa4vDcAVsqg4q
pSPYJ8UGw6M9ny/TiGq6UF3IdaM0BuX4MqibPU+4nkZs5/YmrO0jOcoNNaBhxYQOqjKNIA0Ee1ZN
QBAjzi2z0sTV/tROzZHTSmgMkYlXAg6he57ZU9IlKERCH1TJrlq3KQxRoTu3Zskl4M0hMM06kGcS
3jJLGvCciUb7ZkwEexaar1qrWj/S64Mf2OSD/u13jlfsasB99n/5Lx94RcP0MykHpc2UaKgmu6wJ
oYzO3GbNvtINPPjssig1AeD5eZC89L2hwnwfdRH4RsNZkvxeoxcaC2TVtd47InHpGnqvX6t1LbDt
zReLE2qvVTw0zmags7u7dQ43U7R/GMhpBK5oTI1jLBTXkn92gnx8Gf0irplrMc4AOjJ4fg5UQR6g
FfKtUJ4pICKkdkuXdqPOmheBrGFMEfX/lKoOkUDt5mBis4mygCB6gY/tYkjE4yhcGNO2UEQI3aWK
dchw97Vd6ata+PJrI8HQORqObwofWlDt6Pjfkydx4ojHUoVi/ZX6uwlbcP1nj1AAoaxw+XSMq+fS
2JfafAFJ9Hn3nqQ0PV/I+egpaToyPYgB0BFeDaExYQgnCoNeJ5oRvYYz44nOM696OiVS8ZMY41bm
aTgtYQWjip4yVgYPOg9dJwE9lSDztFZIbSgeB35xWIsDs/XW0PM2k3BB79K4WmaP0irhvZ2WuNh4
SiAXw3trDl+2DvMAIqmxaLQunDB3YiH5CLdm5PFIauc94AG0ZJoruNnZr1xDMvXnPrNGyZ55oXDk
E/HNDp9veUagXKuOGErsyZG4WG+5qjbo7r6sN6gbfdEAbJrobgDZ7wLU/6P6RZU/QVZCodU68qHm
prxvLZPE1L/apyhPM9A4mxyCVwLwFQTXTghZ/SJGof75n39AhFkTOk+Dm+bnfbflFdnZHpjSKHLn
d54BVe1xWHtSLiPPX4iWNG9XmDN+pygL1nyw3q5KPwgHQLMCVq1L1jWzviE4dPzVAzVDf5uWcG58
Pg/k4f7dlKhVf6Lo1qLIbxEs5PdfrNyTXMgsEXAy236zU2MxRYZiQqjoyKwr8SFWjj23Vl0a5WB0
BwjUIGLX7MwJtdOD4Kd+LWz9KfLQq6GElNRTY5XNF3lptCCV4QRiKS3dbpBTM2XCiuc5IC5TXofk
SmQzxGr33tmIk1PNfD6DbmkxL/Z7SCQvRraI6BsY5X808peLHXwHHGrgI3vTS6J2RZnIVwxzDzFu
4d3jU5hDzolQTBMPnUrYnGHT/3Owko/wWU6AgiR1bVQEFSlffeBPme+q71F/VTjWAaO0eDSKz9ZZ
IneNjS37ceAPJPl2xuU3GPYdIhc2QzCHLpxGE0S1b7D/qRqdo5um2ckzdxDA3ni3XC9I8kvoHuAa
4nDHdd4LGEFSEMwTFjVWz9q+teMRyQ4JOLrn9ZoCU/6i7OkkJdAKIoPYmsirGmmHv54i66TD1BDz
4hAg/EJYci5hbB6b/k8R8Ce1HXQhFFYVjsnSmhfECEFkAQ2QRPrSwiUETfDAK9aHC+Ncm1JuY851
0BJLDcgaBKhoGA93aOaIulnSspuxt9USoydw4EjlgvLkxmjlh2WmfWKComorY32yboP7gUBe5P/6
twgxvfmVHJbD9xC4GTMO2+kaTG3Z1EWeO0xUkMFz/72pgcZbvwMfJrrn4d1JPtxil8IBN1t/30/H
MaMncpcWUl5KvvdmiSdHQ7VJjMSIaLx6F8aMH73zSahYjY5zA2X3OWPiGNs8ORyU1Wx+97nmaavH
qwXu0AejAksv5r1w54iVZLlnza/0GxjRoV7HHW+azn5WqJ8AKz46NJNl7S3v8oU5Z+JRCDtlAfRX
GV8+KQ85MLcHc7zcdwCe9iAJ2R7mWTvRrAoYyMZ9JAdtvVU7Cm+i+uavN2IPEFhxau92WOgtPfwk
wRSctdUIau3le3oaOA2vxgaL118qlzjZbff5U7waCqWP5/jiQagt10sfquRHzGiLDuujDKith9XY
Lsp6pEtGCr0RwdL0UlOSqFv/slOR7WYKC3TyibMnEg2LRf4m+ZGTwnxTWrpl+fOjeIekTaCOjlJK
VPM8iqn4mcRXRXfiDttoEZhXhCJdxAWq7VqrgMfwnSjs6LyuUox5Uolu/KRuf8y9jANwgXFVWV61
Y2mMgWu1eeWRoMuEot2wer3yCeaWo6jOagFMNzyiS2KpWTlQBrXys4OgiIka6M/alWMNxRyoD0Mb
FM5Hxid2UuQkSv3XZ/aPa102/+mDLUn5fJuIUinOuq7FtCS2LMVA+pGzszmSnOEq0hUZSc3htVX2
JozYf5oMUTqvT/zXs/tptWGWLziiEhanjxDiCgkSxy5UQszQj5QwLCaqTujupi7W97yR5hGEE5nN
fysKQAAxaC89FsRHE/x/n1cVPzs3Txv+dY+NilAWvX8DQfJea9Pf7t5kUBfwA3wRIrb8cT7td9xv
Ivt9K/0UPg6Cw5fmvG9EFigz4bnGPRSsCI2WP1FBk/82VN9QDgMqgZrfbHJbIyYd6lMW7n430GZW
ZGuFLkE6UtqLMk1sLm2VhC8lDF86s5aUhfyzBrXappXnHspvvDUpzDU/OAH0QpVGr3huQVossRTP
uv8mUfE8KgvPULOuNRl/ncyTEYRN6UNc+AYlypA5BxMrn1YmalcmMvmsG7Coa2fBPtUGUXkoRvOj
BEc0WWskMAkLE5YjHF8PWmBYz3o7SH3PsbQ8X8YFRV28DR3i7g3EieSNaCVX+nfqV9V2PPrfcihX
DBDy009MsP9ntWR8GZcnN+EYk6PVS4J2dOFeFCqyb8qFQ6OeHNXSzk5tikhm4UPkfdUzeOrTbqs0
XIGV6DqlnO3BRyWZFIl08KpR8v7qcVSfwKFJ+U+WY+YYMyZaN57KePz5PBzSUiy4C5p5/AXLHfmk
SwVK7KQc9FQ6VjT+dkS4dVNbvjDsKaHomCa53E5sf9F0hngu1fkfBXGg1UuFouCYOFiWGuySHQTS
HW2dxf5ray4FzcNgHA8crLxmxHOT6QukdJNEYE6YcEkUK8FD8v/zY+d0YUJ1wu365zGXYuFnykoA
m69HyX41JaDBaWfrqqEje+SsVGImBkTs0zpppQJMLW2CG4qT1zGoCAS8Y6o4iBOnTz4crqiPjVtc
6IJS7NVbd7IePRUNvatsh+F1+03DsAF7APEg3XgLcNb1WCSeR8rjuHFmlCExkHcWgLe/wyKOxBWm
O/70uTw1eHNNlNRRMOTx84g+2pnYxtwT5QMXthxf9CUTW/nCevaoxMKhewvZwK5LllHc9UL4oC+N
As0sJJTS2S7MUhPU8ua6pzGe1HmS9NQTogynh6Fhx7oTSY997aUC0OrLfdT4dww3SWbPWR4YIgE3
gzOGsypfzZ/YAr1o32ssyU5cefeCsT/LtHP8cEkizNZalgpSr6tyDT1/BQLAjtul0BKlucHMQ9J3
Na9t2KSrNmNtaPIgsj3cky094t7Po0LyQSIpOY9c4xmnnHTHGGJ07uUqmwcG/XsBQ5HW1pcISR6l
kVWp2xx//7djSsuPasvUe+UthJyzfaaljELQNv2eUevuH0V1TEfBnEMSWEjCQda7vXBCN36DXGMi
NNxx2y1EZWc+bWorPBEEsDJoVsAWxJuqK/GRsJBfG0bol2QPwgcj3UUDUI+y0ChMNPKImWXmcvux
IOYIpaS0rBjvxlD6yLQwJKoqjVygOhNG8o8Z3Ql/Agk0eSLWyxjj1mjQL9RZJr75VVE+x6P96AxO
BPmQzSfnjTHpGrWexv22sWYNhEPynF++T0XbpM2PVet2+6XJw22Cl3I4svRacNXILqFMf3OdFPgO
p+l7w6XwSO1G0enf/PCsWtHb8GDDWWJLFmsEAWtCXk7kzpdqIBjSoZS1TmbkN20vBjPhNtpy7F7O
8xAVZ9hLr6IS62RKowATfXi7cKRi7w/9dftBhnOKV4+aePsY12IKY3Bhyanabj1fGXZs8l/74m9v
d/wR/CooTi70drvR1PyzdbFy8rvyaXGtwxroQzz48J50KJ8LllEn4dRfmSh0r8xv4TLNe9eiwqCx
tpSC5p2qLXj0VjxY2fRekHT3QiNxuI5rHZ9Ye2XL9NEOFCu9cD/cldTy2skHwa9iIlm1VzyVJIpt
jsKfIr+HEvkVEvPoSxk8zMOiDNruMpc6yufiShdDiQJfcDPRL1xegedfImKYCXdJAyN6VpHJWmb/
u3JSdZc9NjsZe+bmidhQe0VcZvpqkGB4b/ebFtIcTMyE9Sb8CY4+RUTq6aUhSa+nwkD/ynykIX55
msSavCqANgqy/qXFOjdLAjt8A4SCb/sw2IvSbYw+unIjWS+AEQhq/Ynn/QAvPTWJniSMyiNsOm+7
E08KVZG2XXOCTUurU9FAg9D2bjs0o6KYMKA8ZBIJRhBvJk7AcL84HHPyUqC+58z8aio60PKwZnZN
5iF9bIxPUSuZu0hNJ5g/coWuemgIbZz/yJ+ljFMttyFjeb/5IQrWsdAl4SalxiLy6KGABiXhoxFZ
N3o0KqxDPqngxAMRKVdOP0LXf5waE/m8XyMDpS2qtVC7wUhv+p7uQxzkR0HrRrvgQm7P0+p3kCGP
dPPlg9g+7hIpfWaQ6/Th8uExMebOeEt+uqy6xhaWkdR0MKJy8yNj7WJnZpEUR9Zp6RWgDjR4M0KB
8iPYffMmvjt/iccCOS6bNn2Uit0OliJEywJQz9SRVTWqADiDG70eAWXvmIvV5ewvoQ8bPn2RSR4t
umV7SlXadPiXX2gF/XiVNhEIJtAuPcIbj8H6+wJ7/JsqDfHu5kH7A4clyLtVkQmZ7sxRpsK77m0A
x/4YJSB+2/X2KN8scGtYbrVhxASl/IreqoY0oM5RxaMAHm6Tv52cVRWoGq1K7rnNItaIOKkJUJdn
75rWrk3yu6WM8zfrswMZ4hjHEGHIJy6unVa/pJXDrX+nAyUxkgPK3umLZAdrfnwy9NfNI+fVXsA8
TLT1DRxQ/+RPQ8QmWU2nqv88yJjUfJbPkXjCE4LNiMbl1NSRR5Ae0Da4YMoWWAg7N2nSRSO9VSau
iZJbJgNvN46K6bt4AimS7pQfbkkHz8hzVuxwI7eBnWuaoQmzNAaZNDFm8jkoOnfvdCTyT50IATgm
829000UB8/pXh0+C/8TCkNDPgg4ITXV7vfBW1wLZZ+IdWli67CD0EgRZ2LPHIQUWc0TsJy1H8CFC
qd2Gq76ZgfT6z2OOkgF3QCID/iXLgW+EatruhyGdualrXjrs1sjAs3reY35vJddnUiCkTjGDVE13
FIIjBGxbVDJlBNnntaJ8ij4nGDtbFAavTeuz3RTolN/TUph3KM/GMye8Ckj81XbzcvCriOUYExjC
vp5E9pksuFXjOuZ1J75fuDrTAaQCAathnECTG+6Gh21MQdtpIeRrre91JOH7hl4G+9T0YXlu2uxd
h92RtVi/q7zqb9Mrx0rr4WexuX4Uaim655XBPW5qAGpmrgolfoKqKu1geK+VaFifAT5s+AivN/Q6
aw/Gr1faQi/UUVu+sautzpJhXMm88Xb2rDG/gxP4u6+26elPKpCFXsK++UC5tqVbaHWNWRGybFaM
+GSWtGmm2MO7ZdSpxdQ2Pc3RTZCTKkAhJrwRQktjZKLYysn6xx5K+8hdpnS8/LLXwawUx0jG/Vrp
xa71INaIAkBoXPtyuxnUAVxPB4rncxrQXmfiragzlQMPQFMw3XAHl2LmpFy01ClhAnVzuEqu7AxU
OMjPE/Ao9vuGTy5GYKWU0TmbKvZlTY8rSzpSYkmmYBs/EDcawIHeaMSsrqfnOZvyFf1Y/0bPMrll
ho53ylRU6rZwZB9dltDGEeWlr48fx4s8fD1XESqBFr4MGxZuv7vvk/1LvwqEa3cOtCwK3kNkv5F/
egYAG2YWEtDxTHqLhaMMcBZI4PMZwkivQLaOGPi/F7NQpiM0E2crX3fnFz2VN86/8/vXHkzu9nvj
PkRdfiWvZ5XnM28Ks6+MZYj9j7cvuwelagFLd8u/CvCUI8O3CbyGoCHA/IK2KVVre9ET7RugaPHw
K1D9XHl2grq+0Ml1Z2322aSZvj3NbIvrZLzpPbhX4YGPtvoR45/1MBn0NBIKnMBMtWJEc+inqZzJ
wNsqYzIHr3pkg9nh4f6Z0j8IMNKj4/KG6ssMMdNQ+GSQPKo9VdQADEiFSLe2cVvi8dFn1hIbY6et
Zs0s71Qu5ex1NIXKGBxm2JsI5K+uEQiianjcS8qCvOen5gHh0g6ksMFAFQKM/xkhZ05KeTi1K/pn
yU3QP7UqhsP3mpJ132sTHFv9oaBRa7Ui3zzBn05fnc7PZRRxaopqvBpyxm5r/UQ8oracmjvaADAJ
kbRrgBil7kGiimEqHETN0XApCfq4HnGwhPMYvqAx9uqKoe+D39Xkm4leGAk1DEyQwUgU5whx5TG9
U4AU53+YUNl67W9qTdwEc9CNHndS4jFFOMFyEYJHxCig7PeBhHlNiuXBpm8z6NDnN40gRRd5ZsIv
fIAauT01nnvaJHSqwBRcZIBQzCYsKKdruE49ZsaQclN7DFzwN6/NMTDGdCn2b+KLZ/7R9EYEFkAg
4JXlhnBhqixZ36odh/ni1GUtXQmztmpsrI5pUx7O19Zm+m008alrOhghPfbZDf965Oc8LG8fHWsL
KeOkVHpaRX/nTK7RqWLu67AwM68ZejS27uzt5xxSRvqXN2N6BJ+DQLJPYQvo2S3JNAOkjySND95+
ic1xnLtaq++1CEqUwWZp/JZGcujtZovVYFpSXYGhlrrvM5Vd5VVS6tjwHtjI+exGLN8sdB1q4LbR
UFvDQ3PgXGAVUxC9UXGEXsZurW7hezMQO+jaKu0HwxSmZeT+yHfmm6k96LP/igv4U290tnD04vYr
Y4t2wJwtxgIFb1hi0ac9T8tw6fvw5Uls8RSpRO/uxUXQWJtlQFtw7e++ueUpWEh5C8DHQV/QyWEY
A6iD0RV9ZUzLr+GZo9lYK9BHNo3tfwtZ0aCGqCqjO1RmPpolnTdvoFS5ih9udbASwwoxZ5lrZqQB
VJFGvNF1UpEbpVtL+Z8LYDKz/yMNyfkHaUvF1htT15xkKajqCMAPoprnE1Q4+piBPqRTHiwhU2wZ
1cmr4kdIRybL56wsXza5SCP7lul4NMKYqFmb0o0ZjrUmAios6PKqTXS03N6lJWeiL6QsWdsyfAsH
+JDR69drDKkoMB4cbF/qFXB1kMlBblkDR1FwjUC5jIOzokL849W0S3GPhTaYraWRJJC0d8pL6QKD
FsCPxTfhcZFvR47e/ijmbunMFxI8vyJkYfyyOLEhv2E2bVxumO9RbyLk01q5dnMBNXKdFs5XFV39
oWFVSnt6PktgKFzqSWd7HQLbX9NWEvxS5Rw9x5M3gWiaZxaHYWRGOgYz9ya9YifAGUEMGqCen99y
gtJ1uWoC8Zhr1eWv8kDQ8WvUWWv1unyHn8POpfK9KibkhzgRKm4S8gZ3RNfULU0yFcrKkb/B+lMF
Eco6NvEMGRLH5hWae7pUotZIbopsiNL7KAFN5yb9tTxF4LONj8a8LI0+k6KvXoyWiNywr83PL9dq
mr7P1ZLhVvYcDCX3xVu2dQ3CFWX9TuYFVe18UQHFBQ7i8/0ZQgPwdRbldfLiv6058dlPHaMnstsM
AloUPkg+QoyjIIz1m4wL4wI7sy8f/BoVtcOudrgJUMDZyoQgz0PyfgySvYN0fAtvZ0VLQjancx+j
7FW+SAvXu7OUfYA0uARYqZkv4LQxGk2QplvBHJMKdG1mZZW94Fxj+iPlFXqcxjQXXePKvQnGWMkh
ziA+h7IvAU0wuU2L2o8SFyZRavugKsX+gyp3vo9e06cGBva1X2eQ/u6Wl7+DWzhmh6OvKM8dH4pZ
fMoD7wp9OznXtobACOWulMaGhGTI56sMKwCiwYXQp6No6T8nh/dFsD0sa9cOTGraVZ16GoOTaO6v
MkcATFp2Vte3lhw7b1sWHURVbjE1BGKhuaiufs5hhSP2DvHgLFWTXI2WpNY1Lbh+i9zMYAoVERn0
FsR89+ZMy5HBIqJwFaenNrdBeYsVQntR+It7LKigC/GOT/wmxCg4yY0Mxb7OKSuiUv5vtKPrKLzk
d6fWnNjZcc9t5f6gW/zvcNlAZyOKoLwgX3HsBMsyEta3KVAciunR0VREAMmgdk4vAx7mrbuEwOwF
lBeoFXU4QW3kYxMk9RK4ZjMg+DeRhjB3a5lKxHh4yF+fFLMBkP/aabKTD8wwB4MQesD2pn4mu1Xt
QZFMhtaSXsvIRkbGQmfep+nn0ocFYEgXpynpCzmtUWdIb4J/FMC3J7Ph9WfGBkDemx1Qw7/yr75D
SmEauD3Cidl2/KvlDfG90hunkdzixGsE5mPUDH+5PK2WO6gquORqcQCugG/xr/9tzocRUOY+eeRG
tK/kdK5aMKtqsrNfQgm2E5pDxUj1loLDsujjitD0QEvxOti1SuI4C9CtzMEJZ/pdoshR9HRhpJvI
0jILxaYam1ePDQhhMKUZfusZBa1cGHNGZ3ZxjYfrbp0mIbUmZ3LpNgE5t5fQHOteLzWL++f1jyfa
vvB7gWRlGAysYFE8D+O2sPnLZFgX3HQbWaNp/VEw3cSw9lWm+zhlYB5g+FVuE+rDOMTeGMefEmmb
rSAi15m5vJzUUmNVruG5hzBZrX3Mm7GakeFg+ZpmUEHAmLZOvxDyeALOxgns3iCAmVmSDLx5loUz
XxogS0D2vnX/oDP5mizpIVw7EThy9fjVyhgg+UDv6SWDMqOF0luvbELQRfRXvz4VFXT+YFZ6LUig
gwSL68AcD/H/SQsncX8C4Yn6PZ3KdFOGvL35Yl71uSGvtA80p4rr4815Nwpc2cPam4zBS6ZbgzUI
HYj56w2f3Po9pVuQ8KjLuYYf2fmaXX35M/jkH9FbJqXey/jUw/d73Fvje7q/VWr9VdrOOzQ8+Yhv
GT18Ej/63P0ymbhVMFf5vLYRdzjgneQZd+EKI8OsTg3RDFWo/g/OND+XRhisBbvfaFXWxyBVPA3s
Mbj7E8ZZmE3Vr9ouPtwWtLqniFP4K/FkDBknPfA6oZPosl1d5j6YE7/I7xO7IXqZfkykoKJG2wHW
7Wa9F/+O2325qMx/RZiSU7osTTLVXJRjxH+gQKU6wDiCB/OY4EHAFs8AnHbNPRS4X12T/KrAOfZY
0hBBJCiYTqo/5X6KSPigXctIUN3lWrZYrWYmwc6RstRCqwmdMWMUYP4lnSi5UbTXZ9KXwl4nWLj8
3Au01eUpXWaOuWp+TgPgP7a27uIW7Twz5hrxbE3Vd87uvaqyrDTpaD/O03Q6DeDz/ioOoweI/ZYf
sUTSUjPfm/75zGXvz668Ixfdt5qxMB8zmUwBaekbuiWjph1xitRzeOf26TgVDDT3RRtX8bD/imAS
lKQ2glBLsZzIwwQ+77tG0UZGwzqSwpBxOjPN320dJPbel6BFY5tCgHozhcjJ8vb/bmKCikYvqLnm
CjUShOesWVq8wXkOJDsHScsOWgDGB0kBgyiQqX4GlesNMmNVAYPooRSm9sHKBCeeu2jKXuo/g5pg
k46osmIlpkzvtaoGnikAuK7I+049Jc2ElhtaM8X0ZqQ1x7fbRjqmBJFAcFZWnG77yCnybuOQP70D
pf14jmcl5VvEYXEOH3d839rrCqRslMr7zcMpXtABN6tLaMSUumKvBkxwO8NpyrtWULOe8BjUWyYF
CnH+9qEj1wHlbmONipvU23EyT0Onld4wMfeYq3H+m70cBjRGi+J7g4j+M5nNAbbSplTTf5Ktap4e
mOJdpmUteff30x3vTn3sm45UX1dcQWjR+c3NK/3AFHyq6gn/ycg9ETfyMCfyZrnU3hFZJFvTO5zg
OwfMaIBNYo/ON5njV2LGmnKiKETT4YUih6LRjOq1mgJDBCA4MwR6stBHobwTt5tCxy6ql2SBPMey
dXhLmFJTcwxhCTa/6DKOuBvpNM7iiIFyQ8Xn0dJ+9wEGmWenSYE9QJvxAsa6rLFxFE9yt1pmjT1p
2Y9SMgvdipl25ccCrJdEjXinXV2fsgeYC/uYkUnY/N8Evuhqkk415cMpAzJrerayMUgt5VsXLDrD
t66Zjc9NR3RGMqzHu/i+eQ81ca0/rVA2x3kCZVOC0quOZd24T/h9KcP/c5tk1nOm3cwYaWmyeFHF
nPD6qk6b2QRo65dlZ95vihBp6Y27brZDWiSGbWg2nWrvohV4HQ+Ju6K74WPKcbPMZXZSMJUaLMHd
QtEydg7QcLc/jCSCgTnYH9NSh7Vx833GEi0akJPKYXsPXcrmUaid4Z8EBHL4HlrTepZb+lBl2okF
VkS7G2FIm+fp02hOIeOmkKHK+VW0tB/wkzbUciXUvGUU6L45r3h2GnL7m+9iw8lFz3/eorulhrc9
/zygjM1x1beRtltWbWOl+AJ+vZiZ6H3kMSooulv5lwke49NwCrK6/+Rx56n1BDonnqEXvGf57xnD
Ju2GvWuCb2ERz/CMpTPsupHGYqg+8cixQcsX9kMI5w/dLCq9KvD9h2N86qhk2FXmNqbAa1CeX024
rnpi8DcV9/wmNHUBdL/Qcv9O0POxM4K2FTkTD7WBCir4XU+wT0zfb9hZtYkPnpbeLgTMYal5FVpZ
F50OUeEbyfRw0Td4NN4cSDAiOw1hiMsuLwNUkUkFnqlyA/whAmyuvaP3UQ7Ips+vl4ZCM7WcfMnO
wqTcWGz3DdwkZFd0MzlUEWuMWnW8ByQ9ibHgOnIfVLoVgLVOuuskRtUQDaWg1ZRaRwL0b/5wn9R1
FDKc5I+bCj7gBbDRtVan+tmNAZO9e/Xa/iCVWy/TYn3QWWHnS7Y/TSYThzniroa7dpHX4XJzIKm+
L/i6zV0ztp7iRhVofjN7LkN3wFmyMbBDWZuyu+fW8sfnfBI/KbVxLbOH1JubEA4diJVJ8aQ/6KbQ
+G0TkE2Xf0QVq8HPJHmPbIBysq485DKYK4zLFkRhSpY9rgpEJb6CfrLPPm9Yyd7j8Ek37TCN52IB
kBkof4Zh/RQGUPYTrl18SqfA9DOYAI0PujcLNSdGOfFWR1TzhklLrIR47KGQ9hrrSvDifzPKG0I3
K52kdjrLY+B8aIJQmmqvQ+pHsIkAa8r/Nx760xhECsC5/yG2UlIG5BVpdm0V7cYp8yMStAZtujpj
JHHck7KP3SDI4+rebA/FOclaEG7OYJ7F9hA8590jx7tUukf2p/XoucK9mlriAtl4bNPy45SfzNnY
G514RlRfQsJTle5cw1qFEWZCfOw7zIiRs4D9a6ZEFEMwlMPHdhpw/7LaFn2uWFpBCSuvBs4juMfT
2bYbste3vIVmEr5MrwHYrBs6qaNSDGd0sM7jzXedyfwjqr//YVj1d06bJOTmARWjAOD+vaTLBpGQ
8gHrT22CCWMrmEX59ZO6xiEyLsrylr19hJZnT7t9rehkGssTYmh789mgKf0k+8Y50PFRevKwO9jT
Yzxg8aBlXGmCk23/ja/iwoAw+hMoqJ65EUTn/gd4c5nxy3hDyj0nxukqvBp6m4vXX+vvl16A0rnf
4RoM2XFW3uu3Zgsl/AYclodBVoVtWk3jTpNaKjmCzghH/7BbowX/RL96tmc+D4R2BPGfh6HZx1YA
qQaMI3LZwlxHLY/0Uq/s42K/1Az6+RBFaC9pC21nP0WD0khJS+hjSfPoqtcrKj8WjbnRjsSU6Tl9
1WC7/a6ksz7Q7lCmg5c26gN09zPgtmjgBcynBkHj7NTTuRlvAt8YLdjJD8ME/MSLRitUZ5CMvvxm
X6yy/T7gX+Xn10CksD98/4rg8otk35WAhlCyXNbPhrZpYjh8XUrWGTTrVVq8fX4yWUK1vFtiLlx9
bmaXMGB7nh53U2EcwhsSDtVkU2RkMedRgVe5v1mGVFuUjNfmdwxAF6Yl/XaNoDUsTjnTWk6XJVJ4
VJrzlL3hkEokUrWVcJgcXLeVYvpzgbL3V2jTi7YJ+OY3JbVwXGedmrJosWQ8Zz+K6XpBG+hCrrxW
Jqmnxy0YWFTHS9VdfHsOJ4CuOS4e1dAR0biDefAOgIgau+S9ua1pc0AIeEohmqUmI6XkC9eTlFGF
4zLbYTRkqk7PbOjqoxtOQi8VIPCBGNN0BKvEe73DkMP67YyfyTD4Aum+uS1F9yO5AWQuNqRU8pQP
EDLytQQiYdJboOf8fj0k+VS/QdUKn8iP6mwQmLlT5fxjyPRqMdLI4HwXx3cgjCQi8NJ4oi3qk9X2
Lg/8rOE84ANCGyDbvtB5hSJiAZIQYk1LOrpG+Noj4AmNppLjrHuIQJEDa3hh38AioLT2k4+YjsjZ
7bmCU4K1Izay0ABKReTzi5IRjRn02/sLwrZ7Tns7/EaO0JaIzTtbhk/sZmZIP9GHY59WPY1rJUzc
eKRfpl8vEl1abNccsWQqRkU3gWVVQQ/iFgAUbYaPgUHZVP468hg6iepGsaEXrTxnKF0N5GJT822v
6drgm9LAyF6zgWXw7pFoepGLmwttVLN1Q1yP7eL5lkGkNHvwx/BMDm2gr6g99O96BBLaVWaSbQW/
Kpgkr1AtT55PHr3hPj/PnXkff9HrFM1LiNp0RaQCvyQbQhqcpRG4TFBmXnB0C7Tmvc/pJMwRKttd
3ocZQbePhdUNv48x/kTDHR052O7W/Rcb3qdrcHOnyhLUQFZu/pcMc2YL7jqcMFOhudEO3iKFd5GA
cgw9gjl7ybKNbuIHU4XfiLU/7IaBEDZY2+cy9lS2zuN4nW2Ae+dDjUH/xhgHcKn+Vr9dHpQPlkO2
x2M771zyJJofB9oGgcaM8jc6f0TED0jSwIlT9dCwFjeHY75rvFs8W21o+yfFSG7O7HQIjguPzyu7
hnPzb6snGzNuNjwROZ3bbEiEgmsa9j9YdAz7dUHonrPZ/Gq8LEGi9y8AtfPujFKchkBqMQsNUUal
D1f/+sRtmMM9ZPmKt8mWA2F3X+YMxZhTEfP4+GFwXcR3BXTQZpSEaM0/1+Y/+dtbJaJNtNTrkFtu
SNhuWcJ7uG8nFthxmn4FEUDwgT4Qx3raWSJS1918caR/AXZnSORSfji4nTNyxC0LqBI+E3tB4Bi2
UiZ3PJM05T3gTO06rXOtuBSExB/Ksmk74l/CvTLw90FEELM9bgXjs6BDy5z54/C9tzaU7xZInjjZ
QajZP8OcKcjimuuvevFn9gwMH0+r0vb0mNH+pZJYJTbp6RluqJ63tHUabfng95EgKy0SsKVNAHm2
DGxWRLACdaJNXHdt4cXYYxH7MhmPlaCKKAnC7KGYQESYvLVnqMkZhK2SrSmBrtqxmFXJD3ntNWlw
d9JCshxEpkd46REEC0zyjDEp9XOecCHS3NPczTPe0aBGjpFegyt555O1t3itPnRTN3a7jhe65BGC
WpsyEv3CqV6alP9JK0eF8R2voQfIoysz1ExdZRWDloXyAwQkeMKTHnR+m+Td4aM5IIJ3xLP9qVdg
Nwjr0fjk5OARM+zBj0bsVgminv94DaKZJQkHACM+mwbYgWwEZlwDRLvSQQMXhBkTLawh8IlMCQai
WyZLZLKMIOFiFG3GtGMZb4tFKP/WcUnZu9U5BVz+ayBTM+x+E8i1fjYHbkmSmLdWpjJyfXa0nyKz
1RZHNHe3fL97foF5sxCFcuccOe2us3Yf+sAGR/jNu7uj8eyDE3pOj9DsJ+CaMgsj8dJb5QMFDrIW
07ug0bRbeC+S2IzoekxqroCAwP0w/r4Dcle9uPN+f9CC6WxkeW+hsNUk8JGMZZCswzWyZjZKzDfz
VxfCwxPIlFSWB7kvgzMzQUqQ5evM61QbTSkSPyVK8ZamrjIISES41nxnc1mIlRT6sZ3CTN2/jO4i
s5nX02cy4A88OENKsyNcOMSM58YlQjJ+p7FM69epOUFlnc12ylvIuvPijs1rw7ggBnokvS+O+0Hd
L2GOBDZdz1Gvo0CEe/wTJ14MZOxC3SkX9S8BXmq+7rO24a8q5my1pFe3D/R8mttCRNXnTioxuxNY
bIeZoTBT83SItyW5EqrfhZ43tCfnjF8b2eqvbkmOd2SAib+SPyN5b0uYOC3bY+xLL+KAmLWBrLbU
OOaIA/N8e11Oz6+jkjgmFcOC+J1Q2+ZPI0sPvptEgrQ/vsWsySY+jEsSI3nk9JLbWLuhmEte9Lff
j5Oaw24kRHEkmZ48MRE1rHCY+k7h+PxnMXdj9oHfY8e1xJ0luC/8nfTU9QoEGc1M+srTJkWR3uYr
FaBtXiJFRA4nB247kbst6KSfv5Vj4czNv40YaRnE4PwHoarxNUSQcfyZTXxJe1H3uPXFupBJL9/X
nC+3y+qimn1Ly+y2HAH+881C+yJTJpio8AC+XXICvZigqcpylIYEkfzrjwW9fRMkFUZCCndKx7HT
qGrmVWZpSbMsVG6bDoEev/XON5aodWFQD9VBw5esHKJDKCT24QE2sHdXcwp5roOg/oVF4sGucH1a
HPuPQ1EIRPTRMDtD9MHpZc/soreqQ3rHGkvep8lhyrytXMWBrhDik3kxdUvzFzxh6LS9v6xRj9+4
GG0R2yIjK2+bAeicybcdIFpwYgl2EISDHlAnuq3+T3QynMZQnP6snHU8kEzAnI9oVhdyGQqOV5ph
TWxkqAgOD9oCCMdDUKewryJNlJxxjbVt7isNjNYoppjAq/iDNs2J86x0psYORo5qwkWQmGfNxFvP
+2EbhDKuS/DhfbihN4QJsIliCS43MSqhNqtGHEYzYBAcoIWoi6IyGEXTyHXVcFMtG9SVHnKNigyc
xtDpOSqXqHmsc7mwI7dNVy16/E9MpbVusE2RwjiI44/btbWQADRAyafmeliY9AK3x7Px7TBFdKZk
ksWRYdn4CZpschbkxpYuqFnHHpGFhZSbGv5wF/prRclZ3pkxKMcRuT14nNgNkqIrLlYZmuN4GdCX
Yxh22u0bvTrUN/Ip1qp3/l3be6nIAeByYNMtP/ZSiSp1SP57KXHpZ+dKx9EXdGvYuswwSaKFsIUP
iGwn+DR+j1wSY21IYmqsUm8/rph0TlGGzI5xSLjScLEa9bzEiq8bICQ0fuDpVcK6y9ZE6yLln2It
gLCsDYT6Nbeq0PSneois2Zm7CHWnRRw8n36tQyYR3xMC86w6QQBhyjiysrGjE1a8bH7TrVirAI01
2122CnDpmDmGcdQqxQOhcrzwKDVKfYP5gJyjOGulf2N3OPlftwMqWbzmAS6nNrWogr4ZZG6TtSgg
0vptyo3cKPjJO56KV0d9P0ky5H5Apbx9Kz+TAHkQc5w3RHRHev57E2QK6wj99dd3USwBEXT+aUqb
tV+DKBs3wngTkFOTBcnhcrjIbzqVUm7fDlPosQiIUt0pK9EbZ3/CxwGt9GZll0W/PbZp/uR9R7iu
oZJJwIcrUjI1Hu1snexqY+9aUoKsHPcpRCBQ5BkNERzE5Ilt+jzfT5lvwczNJwSlX8rsyYC64D9V
BMLWNfVesE+klHKkrbcGYwkLT//xq0OLVt2n3qZeeo9WptS7AwptWflnT5TokjdMU+iiuGLdvi3g
UPfCLV4KRZFVL7CEa1/5U4ieTpppRf6IhysGUM8A8Kr3Q7YWyIE2DIzcUv2DUUqTmd0ORrj1pGNJ
9eERxD5LTpMk+JJBkwwv1rBM+uyYkv2YspzT9zogM1AWUdFzOVecKleXoPiLgOmWs67wowPL5JNT
b04ARXJN4bWMKZdtAtejTA7NKSCUg1l62cQd7/weIBwGhn5EwJCqZCRBpEtOwpKoBmMqkS+6OqjB
jP3F/s3lduQgrrK1lC/XSmFDYGuuEGqDgAlmqJgP7JoDSn7+KpZmRoTjEgMoFGDYEBq/eBk/JMMj
84bcjVJrrHEUCG/sG7af5RzpaaEA37GrfY2RjoUsH1xK0p4/cxQzj+73oLb/45n1r/e970SN0SiZ
1j/wCYBIKdZja2ZA39WKQnggpOYPAh3N8G0FsGTU3sLLMbOnSalUo0GgEDU2hPjZu4QyIpsh/SH2
7WOw/Onnp1gSX5OSpccCinDPdvE9ynRZ5eW82dRYotUVUSDN+9mbNujCjauzZIeZ0jH5OxT40dCZ
w9hyVKdZy6DYl1HFTNTh6EFwUWg+w8x8DzfyX0/65U5kRiGlv+9vPA7MFNpN3uwhJxjqn773ch8V
u+10Hqf/JuxfzL+wUZGhBvsyS2V//8hXTvmDAfT5Uffe7aDWRhd6gUKAcgW9YM9bEzD3liB1cGC6
gJvCw6snz8RCjseFf0jAhbRShXObLZlqPAyVKphrB0VPzvXE6EHQ5FiFeMtt1ziWd9er/BSkMNF/
lBbxD95sl5GT5rRbURGujnhEDYfIBaiRUOr/IRtx8GEdWWxb4wdDqJJx7lHuoJko96rj50TAZ+VS
DIDMM+dfmSHSThg7PkHawg5kZmxojBYmWvyFjHPqDVvpHEFiNfRma0wM/JVcpL76k2Ljgdl1V1BZ
zmYlqk9g9t70xyLd+Eqn5yzjzDQKeF4fBPlhhwB9XR4Eij35OPnG+vybdBaUQryIbvJgf09Mz87s
NjYi1UJPKedaIUmob5+7DZ0ICK5aSt9S7GJ9PyvaXiKoWMgW/J7LAGz9V9TeUJcelwxybz5pDhpK
GES+uOUKP+0zI4Hv0vpi5yamJKdSm7Wv+yFV20MeogUSm3R1XsGmDaNrqkZzIh3Ehc5HjrPXkG4k
FqJY1RA2yV0X5dCb+cPk2rWLTdzzQpF/tL0qXLWT6Ty3RRJ24WFyInJfdkaWLva5by1BVrmKJCIA
8i6kMQvIkhGMuIQtei39TcKt4P5l5w9Y0Z+6+eG+n1u9T0TM/OXeJpffhErCrc/5Q3QLJUqFWFtH
BhzrpOIPtydGQjSExQnwtsacyJAXCyj7EVzMXagKlNkJxuAdjffPeCq3BNbN8Hn8ahINLgXwrk3f
Oh2LcBVYN2S/9oD4W8oO2WGPRQQVY9uIIL4YLHtO+tvLELX5tjMfeMAMXH2dIhaWFPE1zlkQ945o
2sJ+RLv8iMjH5i7Zo/4HYrL6jZEODa4no6lPFofeeFp6OfbtQrRPXDaUKo0ZyhzrKq47+VUvRWy/
nCZM7V5XI70fqETQAjnbaRolQ5nH3WZSNf2bW6Zw9wOygjx9WM30yIA5hBQRLOIWCec7H5+WHHF9
apHm1Kw2fFOgE/nGv2Uhszi+ziri6nHUT50BqMAZU/2eDUbf/qh4/VbubSftUwwwm8u1rPd+q1fF
4ysdKeToqMdSrobjzMhKVLOG3DmYu6Tn/ACHrczKvlOwynnztChqjgXl+xtMs2QwQYrkwnV/p/mh
XXZgCXo5dZ0Y3qWb/AP+g+isNIBRSyEzVJX6f0rYWv96x5XoFF5l9d7hmzqwayWVQzUBgWmCP3lf
m2gU9C5vFEpsr9ILL5dIi/gKpgjOAG2ziaV1L31mwnmt77xKzpgwotbYRsTXi9IHfma3+tsCHCQu
QBniqnLVvc18bQ7vwzlRFrEhFr8DItWc51GmKIJz3CGF2ClKo4wIrRCh+V9WTl/fhvSh8gqPY2bF
7yrzibyeOGr166KHXlmdHnce4RWB9+bIQsKEY1jZUUPoDVM2wQqz4j68GjR5/RnOsrulg6ElPk/J
RJfq23OZxcafp0k+b6hzDPyhbld85rSKv+GkDne3u3gh08guAcjzJhBomCeJE0Fxxf6W0UfDJkSn
Cb1zSK4zgT1Px23uHbFfumH9K9x26m9S6TZvnO1U+X2aIu48nFbJBXHkK1UFse/iprLj/dXCUV4P
N6VItDvfXuuB6tqSE4ZFjq+stNant0ytjPsRZcgqSYDhfuCLV0tDlBYAskcZRzhWMskQ9C4XT9Ff
vlP3o4gGzDS1xuBvQUYIkT6y2l3SJmyTISVyR530slf5pFYy61d7238PzMBl7H3TKVOW/rHvofA5
cROrRXvFZYpDQOvybmDmiUgQg+sa3i9X0pyccYi3lwK/12mIuzN90n9UsPY6gMqWKCLdoUIktctc
RMJMXExI4DG8CHt4v0pPh/cMtimpkrSCIffPSfqcH36+EHBtsjVEsklxFeD97VkQjKpw/bodawPZ
FlIFQovL9JpczJ+lYR2g+inTso73hvth6CZ0/DaYz+dQ+DJgYW8evL8MdwTuAtHDG5sF46fubnYs
vaWgU5iTzS6bZt5kyTcmQ/bqmNKSzYhXLs9PuaSrRqN4mzTJABpDBx3uSvWarbezxLG76a7EdKqp
2qJbiRW1Xt3P8FLJqu7TQr4WnSXOyc2D5belbK7l46sMRiz9PUOf6vhmYkgnRrsWltar7j+kZJLL
2eJB12chu3BLpzPv1VfEW2uszRWEHjTTEJOTVxLtPv0rG6E2hv4ClqwKqdc4vprhKG7lBm25Z75U
Uj0/mQYFFbSmUkk8re3rkrTukC5e5MfbQovHTmUyoSnLd4y+aoTXl1kp+/AgsqgaSgzA6CCv52Ty
SEbPW8PnExrXRbXN05eMV4cbMY4f3EWjlDmrMIc4YdTH8RhmV6MNXsY6OXQRZRqig5D2OiohsgiN
CgaZu6jVOc/8LZPiRdtLmII0HeaNa4QIP+/m6tExQJaLgL2+UBIcF/YLN/gS8fiI6Zy4V1o9VFLB
hwy953bKDXsGUMaqfZVHIHA6fB/UbGJ36ycprkYPGzguDZJUvfL5y/8BskFScaR7xcgmCDFUTtzU
HDovSm8S6kCFEdZcRPdv/aBwrJ1bycn+B3tt5yMykWfBLfUaKRSwNu2x/LHnqrujN3xq9uyh5Ju3
42c7BXS0zytRBWAHg0+bYkTb0U7i69bE4qOZxdxdjYZmLiyBwcbwAVB2XxEeqWt+SQYNUc92YFWd
XZ4R9kLlXgCzFWBftEE78ajhdoCBG9W1cRrUniK02DdbUGuWmzr9sF+DreS5uC20SX2EfBmq50t2
VEG7cttzS9Kmx+QCcxoEVMkY+xIGMGWF3Q+ARJwreNi2kKLX+Wa6kFHLEedFgZwoyJI36MWyqSA6
WarxIg4p6v3XSdVdNARDELGO5LY8Jm3pOBjKHu12AFgBS3SCPbILx73XFQXGCqpIvNAQhXSkeQje
FuQJFG5BCCVIBGh+tn4/BF1tjpK9XCAb1cMs3waYspJZ+RSu8diQL7tpH+ZudNJQCNdJ6tKLIDU2
uqK36oTkhBQHZWaFPonRvZHfcYtETkxLYA8ZTgWc4x/IKazRPh1HjZNP7V0O2ahA1cXr9ATSZwMZ
goVwRFwUaGLneTKzYOEhhQXEIQZmzuFvAdBann9Nz42GVJ+KB+L4vNYrgQMmCppGOA0NvAErGkYg
aBOb3vAKPf3ay/HpaSd/M5J5hnUHbTWAmhYCa5PsH31NhvFu/8fx0RcVcKkSmUVAvAwJZgVXYnlb
a0xM4zbLbUZdhsjDAk1khU2uUHIphCRfPQ0vTLEIaWvxMFa2TL1z8QklgGUAXSnHONNag+e9bSSE
OQ15ecbqnpXql8Q3w4bHBpDAZ3uXaAApo8KfRZggb9JLZWprDB+yCF3zwYV7o4k4CjMArNR8YKHO
SHw5l2puhxJJ/hcwJjL3jwfwO0m/YzQZABBwHfIjtjF8U543cOBDcwAN/W8ue0N42uWXBnvR+BbX
Jt53/GFRc7916L1T1hbgBwaXQtOQLIGGJT0JtB8pIKW/bZUoKN/T4/SRYZNONY8TXu0JI7S0p0Ol
fRvDquL3qlYmmeX8SZjtPNpaXwVDEzIadxXJpot1BGchqQOx0xnmPvkO9XxRAahWzRh6EiiKq8vl
mEfLRVEd8FGGUgcbxeEQog3uS0vIXyForgCIlDeA/QAn24uY+sHXh/Atit8UUhk94ugxbVN59D8v
STYJBORm7u5Kb+yjsWvjur26sEF8z4Dk8tBXtSq7627Kafl2o2UayCn4knSTn1ZwEbGSnigFNPRa
PU0Slai2Hk4htH/x9kHMZpJVhVo2AaXDFwkZeit6wfKyvNdPzpyGPTaZos0M2Sg1GEgtG1BFtM4+
M9PGuUDV0dlIFgmHBMYimKIX9xbbyTfOgVGhk0fHyJ8+0QfXjLNv6gvY9jckUv7hVc0iGdcmzTGT
5RAc57DwlGWefZGHnW7yQEBAO1veNDfUem+YHotpA0zJzh3HSWIT/rgt0EQf7rnNHL/GRBZ/+N3I
oVZTPo1zZqoIO/B5toRAEZFQuNQG4lzc/UH/mjoXOwichrABku6V2pP0JlYMYPGW02cn018UCg2H
whd6L2/I6aaT5lY7HoiIjfNxCXQqZ7g60LbHS+62ApO9SKV7WiGFTUzsoQ4qeWbQAGAqGPOGk7FW
wykTNI7lrfAvQmDjCqO9f3ADjv1B4Jdg7lzv8TunAQH9K0vH9ScsCX5MEJVJG5K4ytcOQcgyA0uY
NdT7uqe/D30tWmNyRzyXykDMxC+0vkgrO+TtQWhZX5ZMGZtMuwShIBaAbtFVDS/b+LC7uneyB3Xo
845wvaGyrO/NKv4TWe6FRoI9rTjS84JMxrtniv4vV7N0I+AhCbZXdbvyJKTHGd8Rzqro9+luPzmQ
/nGAajNAhE6kavloVdw4/LV9gJkTbaWGi3AaoswTkJ074hoxqR6cmrDvZhCPF4WzoNv6eUBl8pzx
DQceE1DgyvYneqvO5nS3AHHvKcc3qyWzoYuUFj1lBSZg5ZNMG7qOBwffenDyYqbWOT3RTkrW6E9H
YF25logflyGoySzrcPUmxz9X7o/xx7FMIdhXdNmezwYdoBHlq0TGLRtF44MgQobm41KVKndkG7zo
IeOnSXWivGe/uNVv+T1BDuFjDjbagCVGpTtJ65H9Q023U2kCb3IJoiPSMPgGJBmQ/X2gWnvePLTd
SVv5GDQRVy39QRmMufTr3oWl1FKEEJzdN1LRLB8skHBoZDL5NFAWKsPg/KN39EEexCJljwq4i7/v
/YUL7JFzNBhEv/kCSFUAZK4qZFDi4CD1qJUv7LXlBHU9YLE4jl3hX/MZGz8LBZxuKYl791ZmpeZR
atGef2aLJYW/qiNrVyC/9Z+JVI+GAQQMriVcWMHRLh5e1xDAil7Uj2XUmjzZYSsJ5Qyuad42dXMt
RtnvBEWtcDMjfQMDXQIquCTU602t3JD8nt8xLIakENdYKIOSYTPMLdzf1L+j2d4/4QwyP7rKOasm
Y7QiYiMw8RFyaJtVxMcY3VxvuzmXTtLqkeQwgGqW4u1MEhAtmcCIuWMyhwtanPjKHXLDDLJF6Mmz
QedOg0oBDbxS0Chde4TRcNExfFIvfdnVrCeUfmkSQ7BTd3UgIxr2Sn7AKHWaXtTZEv87e/mzFq06
H6yQA5Ja/QyqA+rvXigi77V8hVO466iqd929beG0yxeNGSdjBjy8S7uIN+R+MldyFpL5ypjTfPub
T6H2oIQ3iqb4h/I9CmAZZDV/xwTtA78YZ3gV8YAXyGO0950zxHaaQdVW/WhiFqmy8nNzzsZ4lHWb
/DjkA5KYql7FMYbZoedJeJZTf3TR4MxKdksekOdYHq9rPajz1apIb6Fr1kaKaaZknozSz4MIPr0u
HhiB38nMZR5kjuChfxRCMt/ARfe5YpxAsUOx+MzOt8l5slQbXvL/GEgiXKfGMMktEhdH3Rh76U8y
GWLqf+0SAX1C3VYQWW8eZGfluc3Qgx91JH2LHcdiE1GjetfurRqZyIcjiR4UrAhoIqjZ6j7JCGka
YnPTNMA3lu8YOCgWp4TDjumNZy5T4gXc55M7trawPNINCsCSzOqJR0cBwGdLk6ngjLo1SapWKLR9
amVAYbl8c+i7wyhdTQu4CKlPL19Rrp7Pb9MtYuZVCcEIyN+UaBKpk1EOyYQXrAFzGX0G+KivkYI0
rwogJMGN/M/w40O1aRv1Q3wIEZfDwO5xHifJVjLIhP/A3ZhTKaAkwO1jmgxU/2kAnqzSzae6NxP+
hw0zXj9EZzqHtZxI3d1FvWbKYs6p9Qpp6Nql9wayUEl1wm1EUdK84rw59tqkY8C8vXuZJjcDaVwf
Dbi1zxUt6PAxviWXioDTGp4zntS52bq07ITLysj07tSOcy/Y73bxyrBPxNwlpV8bUXikIysOLDTp
w4DqFiY3wgWV9+Z8xH7MZPbn/vRVf18CyZbVDfybTVMHuIFqilS6aD/fFXWm7ae5Wic4VTydvcjp
rHlCQARBNIZDIDz/nb71i/lRv/fZNFwEumSaJ0d/qENK9sFu3ENKIpIOto9Wcq9gR6k0r378jNHo
gVMbjRyxMWIok8f2ctz0jjIfRKUtTmaZNn5z1HJEmKDCW77nfJgZOpQnhbBhejvz08UqgUZAg4VM
7yGrWrYJ+HlUrtBZeZTWZM2kT+qUwB/m5qg6ZBBWPPZ/u0WDNXQS/6JXVDsnn1plILc9ze/X5RXT
OvyrFMaizFBogAM0GjxQy7Oe3UfN9HEA/PtZQaNkjT1hwa1Bi1KDMdnOCh1iQsFnyKtaLaCRvJbH
gYVMc6L4/RFmLSJWU/LTGnyBuj3uxNn0RSGspwneZ+7edeXhNolVC2mmDG9WpzgnH2Z87bsxURkx
CxIaWtpe3/4tr61LGU2TcLLafZetlb7sVIwoEC502pqFl18v026bIrnzbp1M/R3u51xxJDeCpf+V
V0/WwyPYBUBqRZLBh0Qu4x4YEpGBKJlXXMFjuAkHF3S4cYyaJjUtaspR38X5YAhlAdfIWzqw67Fr
3WBWlv2y9Uoe3of0xGZhNdZr1l1mDNZ9kninD5zcPzMbUEM8yKUz8tSGWFr9CcHhew7r0y59mZ4u
sEgLVfgbqJNuaj89Q39DnvEw1loSKH+iFtHPpbzWY9aLyQqjdnCbZTRj7wxe7E6q30WNvVEgaYjY
GtNdHzYwlo3E1us5ZQub2NUO9CTt4kBkuHY936SFLKkH10hNIzaXIZokxsVJgmk04M35a+j3oKLp
cb6uR8lnjBppVSlCCE8g/NqHeGFefFUudtjv8ns9yiJjvL0fRuWos1LkRgUB6f99JhvpTYzKg9p5
bbatMbJKUeHguqHVrgwFOZV2jdaXwfVNCJg7bFMkwfXchnGWpLpR7pjY/jjvRCIts/A/fz9Vii6v
hXaqxqsEX66lNy0A1NSSJdp7Nr1C9Ftr7nkY+pQ2Og5pIZAJe13LT+OgzXlV0mhTo5vR/rAzcrGV
FjUz/Bp2DABAPuT2fIfEbV8oBW2sHoDb6ppCI2toQber6StFuQHIly0M+QliL2ChZ5SULbX2OBsN
fVQXoop+ztXXcQ/+juBvP7j5FKsGvhqBgNPatlWcd5fgsc0+48BIta8SGbCBtdQuBiV4nq16bS33
SorxcHHpO/9E34RbSJiMc6e7jqyKWRUfJax/ODQKVRPVbDQwpRQ4zd+/YcFpRwlRqNfbJSSCrTFF
6iHuXoeJTW95UhNgWiVRgII/ZFJYv9suPJ2C4mQr4UH2htvpc6vp0it/++0yTsVAbg1whaasCqHn
a0uMN0wemjItIEsVjrWwESmd+ul41QapJyAJ/4pRlmuXNTO2tfy2P5UXzG/i7NGfSBiI3ey33aU6
Q1BhSQuwfDTnYehzf79jdVg0/sc5SbpTb+DNGWqHGtscoSvH+tty7O4QYPfydeoqyvnBe6KOjhnE
D9Yrdxs/BptxdTX2Zp1/NHTU9XvUghjx5ju0o59gKYY0gKcQD95gPB5FvS5YcEXVcRcHJJ9LmJTE
yp7xjuCg1xXkXREcICpsvMGZS3Fm9h7bFspkGmd5W46Kx4OocUUSilnVA/i01eaVarvgW5BBSVp/
+KvHNBdRqX3XnjoDFl5GydTKZKPoxGDvqQ1iqvRllLe87HeoLgWiTgdDBvGOGmZz1dr+MAIwevOe
EcUQd2cvuTzUvS1tEAI0kghD15CSENccQHNOJ39sCeYElkMEgSw6nQlXvAZ1L+VqjzRV9cfccyDf
9cyH1nF9cDzuQhcM5/Taj7gHr5vpMcsjW8z+q/xvKHafe6cwOg7tyoFouYnXUxY/r77k7xvVjqWl
5DdMwLFZMI2Ag2F5XmiIylgd5kTmNapw0ddfoQUbeSee0nOVYORlOr80fi1sGZ8nFzeP5r7StvJZ
DE6lNf9F4rCYjTQdfKFOJ+5Zq9Xut1V6XCcicBIUT19EWuf94yY8escOPa2H76ncHU7E8LgJY1l2
Ay4cwClo586eaDCzVs8aurYUBDjFhpGJpAHkDqLBN4TI7Ods5l16uDM5QMZTWvw98Mx92pdzgeWe
4CGpm+Cxn8neas4pxZ8WApQIZGC5gZ+/cw87CImV6Qj7wn/RtZx59FeM7wu8WAdl/nZTP0PXBvnf
zhcbjt1ng6zn5o58Y1+7G5RYBwj7AjVgwDjBaDNf7MLLwX5dkTzjhz4he7gCk+a8KPw/9lhVpgrX
Y+8k8CCN5PkCqgkeM0thoyP+8TI/KzlxW/4OA8YPRbP4Xr98mXq8GuDd53obUxqxsTt2zbskWIso
TE3nZIzCDJPaBmh5y9lhSngMdsgWJzALcRiYhGIZ46FgnJxXZtOI0tMKWoJ/RoUvqIEKZV66sWre
xleiLkF1+5HrU8Qa8Q02oyn6c3O2uVeRJuvIvPblHYFYCoMpmLPDEpa7urlWJk2lIOYU2FZ4BXDw
cUwnS1ZJ/acOR+a4oNQEYCKA/NzTinFLS1A8M9l+/E2VjhJkHIpw19m64R1agFHqnde1t4Mn3DXn
A5LtvU0ciQT9v7EU+Ds4aN5fd1vg3ZgJIfXihpIm8jkXgN5ouo/04Sj71zW1kMBXRGpawj/pCDCo
VmDV8PR6ihXcyep5Qu5BrrxoNiMkWKsDGvFsWgsuSp8SxawibPsAIi4O1fuu3qzahmtAZK4QaJOC
tGiUO5E26+CSNQ7TMquSLlJ8EuB1FgmZ1nT84dc1XtFu5XFGgTYSVdaywWyQy1o4N9rYOHHrkRrP
YvaDIAjOERAbfJpSoXbhg8c4HeWe6FVccDYlm855Wje5Xv9TxA3q9D38Blx3DuOwLFIt0slnmCrM
YVjxY8fQeBeOTHUtzGhPiZr9aiEgiWRYYVkZc0yeFv/05NgYCjrj+T9SBgBC+S9lQOziM9j8g770
h0/R9Q3FJqGn25IWg1b0edoS28Fao/GUEcuPWqse28qJQecC0OVuTi7RuE4Dj+vjR48HpglcEOap
bDORysNrTY7BPOM+6i69H+zjvcdVJpQXySA7I6wu/3pAFl/bRI5PO1BUsbfZHvaWQ62pgjwJr8Bc
UogO9HLRt9QZWjSq53RSgr9MG1ms+OO1OUlftqBOquQBHKFxFfsCnD31dq7KWhggIxTDb1g1YNk8
pXybwX/6bdOfsNmoqSg+IpQMYb0rGbaoqD0zdT64lCvxN+xmZN70B01nK9QuapIsRhIVs+h+D93k
ifv34Ic6yrbqIiXy08TkizgRi1JNTg/QOK5HgrzOBh28+HOlklGU0sH3ro/2bRiIviUXeXHbeynu
sTa0BnDdKczWvsKq6Tgr+X288C6v77OQ2+7o9rNcHxyNy0mG95Mon0ypMzPVt1dMWuOmNJmbozZ0
lZqxtwNYKF8qVGK2PXlOaHid/n4z6opf7wvXOyg2hgy3sq5+XgIOIK5JwEa883tZgQB0Oim9szLo
lyOS+QEXRcAetQudZpMyLPnFZoxmfMwh03QTbZOkwGih3MCTcIzS747Cpb6yMMVtgvI8cTpozgrv
yK4V44Z02QGQWY8H+gzk83b+zfZyjJ4fzVK0/QRRzWlOXpEe7pyqwmxxNjAWvMghQOidGKIMwOjf
yrfiE4vtOCN4P3P0A4OCVtSHJWcPdFS8atNHoJJV8qPouiW0VqMQHmiANcK2d+dcVzfA3TBkkJnF
DgAasb7jHHtZ2RHCV0SQ8SoyhYTiInd2UA47cPabDAasliDHrG3d9gBY5pVEGk6OJr4i4Rg6PBAv
Ncf20V8TCTsge7qM8uVYreeq9HyTGywa6tVqRcJilVro+kYvRetyKIufY565c5oC3uJ2EM+4Zg6k
PKI3myTO/SiKBBfl44GUba79vkHbz+gGrrizIQQ6yt3gPHxS0olovc+KfeADu4Ob6ENPHrxfQqTb
iQ4iRjt/KaGZlr05MY1I+DfVvJcmWSEoUR9zpzun5CbpAVepqn8C590nEQ9ljrCXwm3oyUeCXdbH
EMZHSuNrRZ2wijb9Dhly+gXOD6HBMffLnxElhBIDAwUwli9eIzKIjui5erd3hDNU+79Fr4vJjIq/
tW5b662dyvVCou+F6EYpA8mzdulGRegDi5h066zFt6vwDNF77oNjn4Mvs0Q70LbXJgVc2dFWmCdx
dA//KHg9DmwMfe9OS/cMRrljTqXgbUHsbICdcTh0EHpdLHUFQUIgkfDulqCeN3uxX3ja4ao6m2TJ
rnb16IddXKwTzw/StTEZtyg+yX6TQc+YW75mlJ8o54juL7/yYUFNia1+1gTcsDlVtiWHNSLR3yYx
Ls/8x4P4HJSA+2jTDM3bFUb3sBA6S95TKq2RFQRsr7y0HnfRTSo3WhQcRQpsGhPeyw6VklsDumI+
a4oMsHlMszVN7h2Z17cQfx/6WKe/1LYIuikyryiTNj1wuLFWxAnRMf9omRWNEKNYDe7gWxGIVJke
8AC5xRyS85gU5hYVhuKhcOB6KAmBINzuPG6h55lwDp0rUwyzEiLf6V//1hSvDN0ZlEh3L9UhW4L7
B/dNhUNVLGSQdJmJRVxfARTs/dABcqXcyFezUOuA8w58N6Os5b/X8mwEF3c0dDLs/f/f8RBFx57d
NVekCR8pqdjS2k7FSD1jS7Q7F5NbW7FphCiUP5a2Jlh3XfXlAQO53omoN2DAWfaT+zGTp+zKUho1
sLlEqw3sKhQDCHwxWzlNNyaEfmkMaozafK9N1dHb1cU9bDvmi2dmKIf8a+o2McisbNyF2lcOxwJS
XlB7J5KOBo6d9edcr//kf/AyqPnQHace5BVSJhYq4R4LxxWe0DkJ60KJcpgfdp40wEs5U+vNI+bE
jo9I25DafvdIOy6zA6xNAYhaiVeWP4KfJKzBnr9RlbIVYMhfpyMJD05WWaQ57q+AigDlEvtmlw58
XPOdjFC+P/0k2JkmYKRaVgM1yNB+6uAob6i1RkjJWoIdVKPFHbWD4ZSGkpq4Ll6P/0P5G3jtKMYL
JTvdtkRibPEiqtjy4d2Z2X0wvecGSWervtoBw/SQ6dU3iWqBdNU6iqsoV92Vxe0T8ReZn5YyGKnT
nFBG5mIR9VAg83owkMt4UzlQqXwT6rCa7fxsNnG2X3XRMW2GrCeLoZEdR7VtFE4alquT7g2vr0TQ
H+g5sOKBzd8nkfZsARmKMZ3FPPDxawJaZNh+3u60IqXmgzNghqR+ZQsfUJbmHfknJ3K39iZeSupZ
PazLU7o6l7wVeqL4Mtt33agiHhFPjfL5j3qYtfoQmXo3QNaw00jMuYIb8FnnJonREn4KkSaikaGF
IYeoxri7SkUzsrS8fRL2hPKHZ556jL7S9LWVTuo3988y733kkeoRU0LkS44D9TbhpHXqvbPKqQ4g
WNky5XTqQF7VbVlTEfuAkA49TwQSanOfYXAl2OiZoaUdWLWudxaPudgKGiAaKAR6QL8IiDpQcCTA
A4eb1+TjouY7nzpfgFFm0g3Dyxon+8khvHMLrPTTuL3lR65r1by/cZlRGutkP72yZA0WnOGBhIrh
t0WKgnlDJjW/OncmLb5VMtjSeyZbTkpd7Gabu8GadOHmS4INkyEmPLBB+SLoFRmDhwPGYQTkG/0j
/nT79Kn2bZGv6kNtaILJwdAtzH1yvz2DEm5hOE+doPUuJuOBuiOviFtWsdegdV1rGyNZyyt/sUyh
57XSpTy1irCSv0KA60bZtrpfWXmNN9RRfLYGu2W0tGlTi9fahOxVCPqu2vtQQ8tB1ufBQIKW5hhr
lN5/5IG1Mg55snORp33qxpTTRzkMLlH0eTjSoCthwI1VhCgNgqRUbyOZpRI987aElh821YhDOkKR
V5abp4tLnduM5/xbyQ9DcGWRQ4svGuAFG9x9NaOXdOuGl8k/KgwIjkojsW7dGrZGZlhG1fMD/2Mn
4sgiJY9WrXymhKPsQv2WSZF1jvoyLqC/AJJlQkaq2JZTPaXqJnYRv9ytUvUxYnnadxpJHf5Z9jlG
//Lu1PeE1gFFoHNcm/oN9p1ONVvZVhlWhmG+3LlJxB6hyPe+qgZc54/Ytpcb7DFe8GeSPh6wtSfG
GAwvlB/P4DZUdn+mlTRP7B7uhSLVkJrS5pQetq85ETYLfLCnNl6tsbr6GEGPFKx6LDU4bbEie1W6
aLJmCXxQ3oq5hTYdxvZcvQZUMgrYFE3ULanzJdhCVZ10lxAaIpru8sq7vtV5Dq+iQDKZmXAbLokI
eMylsZcQbj/vO1puD8YqHPH4PGM7rhtCXZ19t2PR0a4F9Xt5KGziHbS6YSTQ4o65jNZDTci5fOrY
E72fhsWWiTnzdgCCQxkO0bBgVqBazNm6bbmsQ4Xhb2QdYHvz9QmDqQAxA8wW9uwmoX2S09TseI10
rvMTwNLWx4MGTJJfMy7FC0AdHlT7uoxRueqGVgz2SiCmz2lLq0p+weuVOmO30nzJ6TE+B4ugPNdd
MjUxkMNAZHwuPrfURsXaaWQecwKeHfNiWfHH8/n9wHENg17CldmjjvT2f9DmJaJJF+xSTYY8u6I0
35MGOLt8svN+8JeURUFgQ3C9+Dr9rJSvL2vcZ/cehV4fyh1x4DmbZbjab7IucsbmAtCsIY+EARIh
vYCQymzMxzic6cXPs+rq3K57mR3cNeCrGu8+Bb7HYHurSjTFN4XLEgJrdq0ixRaTjKvBSLNAidGW
br4dW0MeLhu5vJS2qTICa/JuHA99tyElJcY5pzjU7z/mw20Zvo8ZJyvh4G+LLlnL+jzSqoU6EQaV
3YjyrSSIOWX3pzcaRjZpYcJaGdNmnkndyqk5tg8QOOM2GYN7SUQw1QIT0Z3tHMmWdv33gv0bHVsr
yi3t9bSmVG7PyRSmfsQtQXbIjGtV/dQn4xAJuKXxxzrkRcym2dtWkvXAgUHyaDe+dTKy/vv0SDWj
Y98TYZgA016lq+F2xAX0oepFXEpPOrtdMwk2+fU4OwiZzkltooHPgyGmLVHxx021pFF+gK+ELkyZ
cfK8Hq9gBCVrlURiJfOev2UJTswFna8C6xpUAotc8T15ajUqQ7RylwYBuoiSWExEgWePBZgwETd5
JTUAsnipMnDOmLsE2keHijl4TKZbEKzi+r3057bGIxZsbwHdt9M6pWiTZkAS6FpCNoP2gTe0BseK
TfHMSMdNcIez3yRsYkesd6MLBs+8jPF/kAOysfHhUVwTi334TPlFy0+6eLYcx80YpZXnXUuk7FLs
sng3oD+4Z1MSe7KqIute5HYci34CLtWUKCROPMtLi7Plv+ibXHPltilghmrv5QrkPOe+fIGKfh07
q5qdoZbZFBm/CJ0X1ZvwSaJwbYTz9da6mqz6C0MHFddXVC6LbpdaExVVEeceqKSEUVKeIyTzmfAV
JUbU+nT8iJkojp0VR8GKMd/rIrRQ5Cqhl+YyBlAR6T/QrxorgGezZEW8FxFLB5qHohMNsiUoJzxz
jqyLwiKNKnMXQgqBKNnrXHM7LUtMxm5pJGceworvkr8TQqA6tb+Ev5utg5nQDWRVbShQXXsTzaUU
gQUyN/4oW+irgb6YJ7Zhg+kjTMrk3i41qZ3HAIyVluAnulXbUOgEnFJkqKZf1RCD7+W14hsrMkLi
Zd/O1gvUmCDPHJbLv4og6x+KaIhP4Ql2GXa5WcFARCeZHQ1VedobS7tcy6oFNK9dcy5cwd3qs2lb
TUVSFoPmRym0SBe3eIw1CCs/Kqqt1DI4yg0bRX8924TWVEQZSSTKsSOkGk9QAito3rdJA5VR2Zap
ysJoruQGDniS8elFuXBi7uAQ2DAjjE/o6cMABI7txMlbugz7w34necfahzCmx8vlMM+AU/Pk9Yuh
SwrL/SMa9W0MPkNTwOz4+t9VIizrwP9cI2CCihhgDOlHUjdXjkYUQQLJk3dHVUEVV4hGN3qfGcjG
tH/pojQKIcWDmpMIY2t8DohJmzV+nBY2AGjH8dMpHUHyVLNA1YTt5ZEXfyzf8AwVAtgxelwZxeSU
q4kei5vvAwI2ciD5T/c/HETSR8DjuPfLZvSK6491n1Rq8B32u6eBWeGcupi6BNgCTxF4Ui9iHDGZ
jIQ8ksjef+aPkHmE9iyJQglglhyBuaCl3FXMp8xW9k2CaWWOU+aX/D8QydjqRR9SKgrrf3+ZDln+
uuwroBG7qwjcy/aungKGzeeWxpLHfaBpkZIHZRHxFpGxgBjp9MiXUU/d6T1zX9gETDSY4DiN+AOE
c8qjIFsHACxAP4cH28F2jXsmlINZ0yN8LVidiAEg/ptqKMN+kxdHapnIao9ZLTOpSmv0nRrQKOft
yueSZJ/NcrxHU6vEsT43+s6x/2xyjsG6Ot+9Kgu26s76RGd1Csr5dSYPdBSNXrFd3DmZWNw0vIVN
bKmJb03ER0bvXZTbLyKKMbzFdCwM8KvTWexwPLKthGH0qvT6EE9f3zNKcEBbiUNvjX9M4+aHaZ2b
mX6aVn1fSbaV1zQqd3Zi9ms46XobwQoR+7SQLYuM7obEAvP7qhR0FyJzzEIaBAK4KgoNifU4h4Xe
Vi7gvTu792jUWf+7iRfDZRjJBsv4SIl2fSIvKu61Ds8eGiit73I92xXGRQ57O74QoMkeIJc3qmAk
YYjUCYuJYX/K75yJjuGsXSebYFLD+kYK2W+gpgYkPp51cpnFGjkc6RST6ZVW6ukrF3A75X07WVij
k9UvGrLjPPpyxtORA2gA0cusPPAq/G0j+L1AkYe47n/c/DP6ycVXILS/V/z462IekH3adSTBZZUJ
Ocuoh02qJGBVaIvDs2fjJA144VoIotkLh/mEjtd1J/zidgsPV3kwnMkQGrHt2OqFfjR8rgZcztiL
UgoQRgIWeBKQVInpZi+5peR4shYy0O4sdIRUHGKmPVbgw0UYMAQiFPl9DUGVYZMPbKKKrgVlsi0M
ipB4cQNOIXtLvgqUnhtR/pIYMDnTtPK+2HVOdMdFbGqRnZIvHLd1MRUiOXDLZ0dXQfeBAv4iWfgT
uKi7YNiVManaFQShFsY5sYNfhmXDHtJ2Vs5mI98LoL4QeuEv4vNigT9uPb+TQw7KPzCu7NnTPyQ7
VnF6J0m4g69dsA7skgtFo1TZc7XgTw0uEAa7GDsY8njdSagVDrR3GvaNKQ5KgIZJURMHf71Vh9dn
gbGGlrlus3i4IzV5A0X1cMBpkMYRM1JuX1j9hZCFyT5uAxSJIvQeXAQcXhdJsGAN69F087uiP21L
GD5v4NQBPpWfj9EUfM7AaYsQpjkDRNoP8vgMjfxV+80OdnPXPELK5WSWuRL7/BapGgyPGL4OGMdu
+KS1n2UUxAJlcHF44sl1l8xCpLqIo3mGOvz2simQFbqCSeXIYApIEYUE+LB16gMwN4P7zwHCFW2X
PpD1jsCOOOkg2vFPxT4FQFm/PCZSo+RRbUR22mh0/7MemYpzRfKgLauRMxvoLF+LQ4n/M8xnkUAq
nyFT4dQ590YxkDtVsQkwNOtvtZbzmXQU7G8xbNK2CidwljPadqdCNpw2Kl0LIZDyjWEKL371xaGK
9kxpweYGdneP5v41Jp8HzteasnfWqzw+5gMmgNBZLnjDohuGeSOQTJheoLLvXlNOIyWiqBm8bEIN
Xx1GYJ2eEwcGfvMr5hRS6+eMDateWLgeGH88tv3IF0Suqb7BSZPfoo3ggyRpwX7Xk/CHFCqQ83S5
nd+3+KxV64idvcjbJImvs3+7lqm+X0V23jX62iwcxTblKL0bPeEoyyqQ+ayNc254TNanbiV6nJiZ
vMO6d3/4m8w1NXRKB5OML60U4j4YyVRheBkBU6UagC82Gvz+QSodbRKWwE538OfRD8Xw0CAM7f9y
NoxglAENefievHMnkyWq6/7p9D5e3Y+sdYxZ5aBkktkQYbsL9Xov756IU5nhjM6EOn7tiR58vl7C
jh+RWev3QNJotFjK26SqYB36UXkOknNqYLuL928r8zh54GiTFkGGLOLBJLEIFkJjdkpf/u98BBOn
6QP0zBD0GIorJwOZXSnaI7f4DkF5aL3EXsOgA4CejpcN9BHN8F1z9Z+Cs3JfNaYugD8wrnUA+rhL
oDAjctXNYRVcJQXVfrjdzKl6bsCXBts/F9uaDjJh52kOq5d4Vxf8rL/Wyy+rJ4JB1NRVhS1XzNdk
EDli3amPaTdBZYWf3ItOTZZawbOUn/9x5eU5Wwri7Pos51tF15OC7FnMhL/rbjRQJnwBfGqp1Tqh
myFxyiJf2Qwtw3IhYQnn9Ymm+48WSybahJXwRMH1bLkrl+Mv8curlZgOJMMbVzV7eosGhdTXCFQ5
LkWdozhLYPYyBHCNWRVd9knL4w872CEVHlEmS2yBFg84qgJIFb7ZHSxNbX1/JZ3C3GIwiF3DlP2N
pD+oU/HXXdna4nZKtqieZp/HBq+OkkkgmxgtRAC64mZ5Dy4h+5ukLONa4Lev+xmod+5x+J0Qm94q
rrRvsPlVf36sE/9tNwCL2X0vfqz3DR4ThT1LCQ75CqN0sccLAaFQP8ARltLZDeoPQLsxLnnDPRYI
Ei7EFCAt21dNoNaBhPvrUBFOJjaJ4BZ2e+k+ZudJ2Sxr8gYQ87s9469CEUObHkWB9I3t/Gup/frE
KB4FwABPyYfKAcdxoeHNhJYZa/3rK/QmuX/uk3vlTPaX04ht+0CZg8bK3pobzLDclMYg5dbXHuV3
mi4FjfUo1OucP/lPULDWSiJrZ83Sx5GH7ox54Lk2+rzJQFb744xaQrgyT2zxzLesY8psF9dXge94
cFpJcu6YsWA1UOxUMVunQ48PLkoctaaz9R4fx3UagOw3LeNAtLEosLpMlxXw8LqwzG4JrdHsdlu4
EXQfMYFrInFg5xg1YKHzp8s5i2JCYrPqgCCEKXe77O7GKYw9s22zP0sZrddd5cTKEziQxwshassO
AGT4oh9UOXE2RCwzxHmo+967LNnUZIR691zV/bQeFEpyEwxwCchcisXL7WqXQbqghny9UyKwCDBI
v6kdSz+LFxAzbbfCI9iARN+xR/YSyalNYsuIO+Wtcv53crp0uekwaxjvMjWdVBzIripoRf41SYWH
Hph6n8NKtSLxvJc0xP5n7xhtkE3z1pLlynJVTjC+HnyLnDq3leG/KQigTAE3WJA7TmlyxMYicwcl
/ujdAZpE8LdQEGdxJAoD3XE1yZw3ZyhaKIe5DjEmJ2T6ubPioaKFmf3fOFofXZRDWfRgqm7lef+m
0wT+xM8jqTuhXKZhDvJl4wOePWP9ulah5F4ZPwuTf6k/pKrNTQOtmekZgrSwLI+86/CDnpktd4ew
dpggdxkemB0qSLL+vQW+tf79bSxuAqwYe6EXyiG86lfPgws+HlSgblq4ORTr5yK4KNvpGIAfxKZV
RlNG8P3Nitnh8uuJj+ChM2z5ooB8L2d7micNoC+ptQy0gXtviL8csxBvW/xOfgLnkvwnxrz8okMv
ni90G0U7eW0rk0qGgcS4pu1efveluTak7LfzVPHRYXAsAsFttu536BvLA5M7mnul4i2+Z5ULSBPc
uxzOWSXcD9ACX9MxmlC7vOYQsyibaq0nfbyw8t6ff/BCnvw3l8Apb5eMRxiA1ctejdH56wunjj0z
lKzeh9UXq9WlvR7GzjClF2m/0oXwnUvFNNhn8wDcezmDPhTZxv9nJuapK7uY78gSlhBL6ME0L8Vb
kTLnUdRgdludS0mLgMRu3XaFnw/gua0dLaxo3DKuDs2ppuan6Rz35D3xWlAfIp+1WARd2ok+zx7+
IKPdleunw8IghJwFTXoEIZMv9RcfOiceW/f5dqftdkW0LLPW9TlwfJNFJlHWR6SQ0VBYXvv8GDxg
3f7PehVrBDES77hpd3LNBuceYILmaFJQBB5SVCsaKZAZpY8o2QIjMtB/XhaQr1EpIM4Ns9gTDupW
RPjYsxLsXT6QvTObL7X2fXbji8jORa9XUihByhhuQOWHzzmFoggviHhWjPnyq6RJMTfuM7rGl0lF
/fQhzzQWwqh4kCjXWhDDMVVPsV2rQPRHr75/cuvjLBDbiZ4liMtirwDz3h2AY3AXGQp2FMJWRzJA
ncq/Xj+JIYdVGYOmkOvQmThqjuKG36PWpndDjw58RqyVriIsf3Lq9k46Uz1e7Qi0Jd4sXOYbKW2B
n7J7fVyIbkx+tQWt05HhdHAJTEsB7r8ZRH3AxHAIBGYZg5n7roPUn29dciVUw82obvWw+ZaBHpuq
jXWo3maq0a1dSLwDrp97i/kgkvfWjDoPVKbzLpvuvUdDc2uwRLLkY6kyIhmJiISbF7ihbOGCwRuG
w5Koxk9tVQtQ0ooFJZ7veLlwT5PGNqST3FReFjUFdxU+PVNESk2Uc35SP51iTHehT4zoVeMzxeht
5NPd6WkL/Ax90nULNAPJYNJmYymGD6oLWZptCOm5I+HMdRy0iOXlOI8cG4wRxQnrLWIRHdO72g5K
F/Ig2xsI/LSp4TuNLobPU61tJxelQIHTVw4N4isob0dDzhCzG/9Ws6kheeUHNGVGRE1mBp7qqCX9
tko98eDRcgPzWjmEsDgVQC4pqTJSSB3lagNpOweYi5FFbfrw+vAe8pjLyzmAxB1X8jxBTjeGz9nL
ZCRdRmHAEzKk1OpOXJTVrVZsryxsyWGyZ51AtCIgML3BqfYTGUFun6iLkUUM8XThNopUeFf1B4Zf
jXQYepw79kCqqeQ6mcUsj0X+sQ35X9E3VkbQW/2AcPA3fxLzMhdjsVjMPZVNHysaEfJzc5//Jjd/
MEEAbGBsWE7k15Ta55PJ2S1NQ0IQHpzNujt8byZsct7+hDxUI+V+mf3LfiUvK5h6BqhZCIAiIa5m
pdwDm38uuFdvbzKS4A/hIrvcGgx8ye7J+rN6pAajHGTIM2UKPLEsoHNYEdfK5iJyNwTlcT4yNIe0
5W/x655Eby+k9mL7AZINjJNVEk0i7VI5bSsK/2haHQlIV1nBT6lXs+hqCc6h+2LQHFR20YrnRiCF
JhyRRvFHn74CoGG88KgjjU78lGIF9JKNoh8qWy/PvS4Wl4BfpJZ9dawHPQ16BbjSfzcElwUa3pc8
9B3VZ74Y6PwFyLQ8pT99jb3DwsAA4pqXVRpVlWd4TPe7TqC+7NKBmzNjVPBivtekiN1a+gEqAShS
MiQRFeDJEMcJD7DMzQxQLNtJl6iCO/9cHuqxkkqSEeCDs8OgvgrblusDpWvzP1WnGQKEmDzXcMs+
E4fR7KmeA9PWp/xA0u7r3AL8IGGHc5Q3/6t9Fbpp3YsXGx749pPkGZNEmnhKeXOkfqkp4BFHpa5h
GnrWRa6QbtXlAXZQCvSze6+F71aIpyYokRUKzH3UrygBpbhXquW0EqHuy7dL4hgq3JvmaZHoNjq6
ScvdG363i25g7XleRSFUwgEkgcbPhsLJfbFPmPkiNj76rKTkx0OL1Rj3rPWFLi/SLlrPdT4Xrff2
74jjYGlK5rXB/eiPKXt+sDUWEQrFlzwBA8+Y1eXJ4jFlyeZH8Ln5oI/bP/deElcpSAH5HgFJGDPu
uk7QeLjsCDJmBZjitwqXGj3T/FD+tpXC5H6zcCC75esoEkKoXI1NngOP3qgOXhlKoR34AnurD4nw
4DYFcnKGMbGhMdq2xcIiFM7x6twcwjjOrkkXu/356QbWJMFZYP1KnT/nPdQYWRhh59yZyvau+7RQ
4laUGVFRl+E013OKAp/EhbsfcQkyZ8or1kmWn5aaGr8FDhEle6fHzcQ9qgg5ViWJg4el0z6MNPMZ
3+DimHEwRYRhmwahG1ByGd6k3qr18bxOaJgkkEdVc1/qT9m6QXlEpjUnvBMCOn9CdbPw8A0FM/Im
kyFIA12H6hOo04bBtioNVeBlt0uopmnvpDLaicGQlpL4p9IAFpSh2zebOEQDtlxM0AJwBNvSZBY7
kfi3oPUQe8Tm2V6nboRsdHqk+q/gXS8m7EiovanjfyemduE+90jGozgEmbrWjUG5c4bxwjf/EBnQ
YuXtS1RdYkQ3vTDncmHwjatFkgRgoTkak26gpCkxDh51I80wQ0HNA49F97hBiGcNKwfn4rhSSIwV
APci6Y0drwSveLM+I2hu/x3KOK7wnuN/QKvU3dOgs/LupoQgbdWY7bIAb1mmYXSfYyl70QS5gnUK
mRoueAn8fgZ5RZJ02vB3PPnSo3/MqGSHGNpeLVkulY/rTQFeQzC8r3XRGff4+DFmAj1/0nTTHadj
LPFLe/mdcmWpfR+pKObt4jaRei3mz5kc3kB4+67hQTd3H654vAIdDmbvDceMjw8M0T0W8ixnmbky
SYbU6y5h+H8acx158ic7ODnZsOFNTkwreVfkMbFzCj/Zp9QTZwD7e06RcEAcima503z5I26w0KVO
WTuiABPCjrwtC7bmvm4HvwdRRjlPRlkvZqEE2uAHCjhFPHvYBvOnjCbd0sfSW5W8JOLUrhJxgH0D
wjN4LFrd0cyx+g7UNyhajN/VjAnEM1LuKuAaceB0skIDGmlzYejD4oiBadxFmU39V6kOqXL+9rri
P0IpKN45AORxbwPiUC+Gy8tXUl4o8WGd5BbfwJDw8b7ZWse6lHDNWxOdbOWL060DH0I1CjZ6wPpE
luBtZ5cCiaqBZHPtZKG70z+a0xh/DvpATgpQ9TGHuGWewUJY+i4uD9dxMRpgscte3XTb3xI2H/iq
9RXpeX+gs3sd/lgJEgv9HOyuSaei67sSnaslRNA1WI4sx5qYPv3gKtCs8i50t+2lhv6FDANqduQY
iOEkX8AbHpId5DQukIII9qnbmRj/3qZG59nlKX4nqBGDrhtWqbrLb8mmDXlA+rMKKzzfpqorn8rs
g7CqiOpWhlcn5tDPGdrxBSBPz84y0PTiflkmpixMTTykNTgB3fyF9w74sjMlmQF/3RP1GDvTTah1
1D26/LUmoV6xRS3N62HyioDrG8AcR5B0xOYBOe3fPkqfeyO+vaeumG9BGbV5ThmJoEgJ6cFTfx/j
czAowMGO3ugBQRiDJ9ITwWq/GkN4tiOOqq5e82/82exM4UVioLl/UECsdTF+ZUOyRMWERu9tN2l4
93Ro617vqdoIZD4IxL72YS4EKnwmrsTW0+EBaTs6BfFLDXuusE8Xlt35QkhefaQdwde4/w23KDwu
ftSAiLMs8TewShmslswpHF4U9RYEMxr9b/dz/DH3VT6iwalFHOYjzv+ULmrLXueq717kuKMwc31d
MvgOKd9mxAjkmxjKa6/sT/zCeNc53XL6Qht/DiFgzASyzf4TbqmJHTss4HNRvp/7m5dxD3F6miNY
qnLmbtxp2DQgR4yOq8Gw+Eix080bKprIeSham8CP9BjeLzbrjDON8GnSea1CgG9QFpRLBFncFv3F
LFWkFIL7HcI2V9GYxLj/gnOGPMKfRuRJtVaY+JSXoEvFJnr24SjMZE+rK0PaqAsvLOBY6Id5g3xe
TrmmFCralyD1PbWbcv7r2k5t1bhDlJjyhGBTBthu69ONhx/GCTG7aHNUzK9PxAkvgWU5Pzp2pVYT
0hwGcW7wCfMlqa2vOQzeqVCLhoq7jJNmcAGEu5v2m8gw4VDMGY0+xSYDpFmqGYWpTxEvY72UQob+
tdCIF1h/nLuFW+8iA8XERwelbPlNFq4g9SR+kz3XxXDfWMr+wqSCu3Ig+jOCjE7Xipenu8KAzwDi
9/JlxpdxJoz1+OP2fLZgb98mXYi9vRoDR+xoOKBX+DELUo6TuvwCuiZSvfWiLhSixKogFhzXSlf0
jm3VHCGrvL4TDT2Ekk1Y0WMoYMqevEI80+BqdjCpokWiX2Cx1NAg5EeldI7WbtkhbAqhk4VA9pV6
utXLW+6CEW4yDX1BFyYpnCFyL2YlDBrc2BZc24l2Kli0nhEMlmA+BcVcKY1k3IMulEyGgUxMjHvt
aUW4+6eZZtJZ+OkJrvvzA/9JLysPy6yoErpMav0N9I0Yri6t1zKtXwKqrDyzzxITG0Miqrdkq5XH
7aJ9gnHMQ4YinuH2lliwwwdFKJRWEeh+lCzUn8eXTyydG8+ICVwPU/s6OQZPBa5rAYoSpWSKog01
JT+rDEegEYaLD1meEDLLxNI74ejLd4LnLIHKMzu7bF+kbakZ5ycNctJOyokPQHYw48wihSgtyqKq
1Ln6iwZHWNrdlnYyNn1aRSdvjwNydF4cx8ekaRGg2YRKrZi4IHwTuNyTArJIj50HzrbiLYexGyoI
Ss1rP5bBkLo/oAQ4Xzu0mRpYfyJ58h3U1KZNcJToKROrcP2CLjWLhc84zYUYZDyqWIxNsk+JYsLK
h2IucjZv+XyeiHCRgz6uGRtw+cOIKm0xyT0KdRMDgExrgLLtKXfFQqBBdvMfy+3wHtEETiOkqrzV
Y7veTqhO45ygx4uBgB3CTC3CDVgmOZRxrfOcC2Ua1x07tHPmsZCUgW4AN6G2JsGHsHiS7tu0O2KU
3NUNoipdYWFSWspOPOhEaKu6RrZXGJXtORfg89ZUK0MzVhzno3YaYn1FqEEjgcoBzWl8OCiPqP31
ZQgIDdEcmFDvJZF4nLIpVPTxjYmIA+/HTA4bclTKH945zeOQ0nLwQq4g8Ui6rdpABpcAWzQn+Rbn
22xK0ComMk1LAhonPTMl3aRnMvawQ/mBOHIz3f2EQF1Am8UvWtYr2ylp9fSkYaAqNT5ySFdq4n9q
7plpjAYlLIJ+g9I7IVLTeald8vCdROBEPmECn+v6/5BeejoCHzmy7c985JZgrjlq4EUEKA+nyjCi
qkarC6LQR1lxvjh04F2yuDSqveYwzmwQf4qdCvxhbS+SwgTy2uAXwUxtpmJYekzgD1zz/2tp0vIS
U7poEF9A5I5mKJdhIxrMn7H+SgX1DmsPMiImoaF6mJvORnyQc0uyDQmpxJLdsZxBvAUEa+Y6ZbP7
7qI9T4F8lN1byQzt7Q7CzhA49HFOPQx0TCYxas5GACTkvphXILGyP7miWg4cW/q4CWEAykPxqGcY
yR9SPIPaa9qRGPuxdfppfMH74VPZxub3BctagFtRcJUfEzt5a6e+Z3/XWtWc/hl7HASFxU/CGtKv
bdGo89vPVKIqpAA6MJRdMiBlrOWEZuHPT0TBE13DvwhWLpXU1LFGsaRqjcILYc66AAcCpaWb9f4f
FMg4fk9dV3oVOgcdS6zvnjC2pePcCF9482i65bKihJfe1PI5Gy4vajhPgwD09aUC3G+yrEx7LDvN
aKb/4JOrETjvdEcdQHFZzFWX1MwVg+YLub8InNUZq6F33B/vFdd2SjQtBvpP/hfFc4Vr5H8WWuil
3b+QXuPok5O4olQXvtmVQ7Ph37qVZJQx1XLSSoxz4UVpcklymkYLhtWnlGDs+zXkg54H36OOiIdo
3uGeurpuX6xskpLZNOqQRjOz8Gkqow/YzwI+3/HfD2oQimmFy8Oom+0fkXx/bpD7nMQNJ1ypn2zE
efdyVcTEQWh/dmWByr587/+62hWGkTEc1LHem0XsF8kg6Pkr8REj0KLuEljVJjDclDUhKM7u6eNZ
vKE75hWUth80e3AU03xIkoGuA8TKIzwhZTZmDgtXUIVMpTVx+Q9dRv8yMkJ29fEo4K5PEF7diWX6
EWuxaie/t2fZRpzJcypdElfqXvmfRiJpl1nwq9qTX/UTrt6NWT1Ff0mCIBXNYTWqcL1GvyCCOGT9
uMkJiN2wji2ECC1tXTx9KqNlUH9UonzDN7u02/jGpoD8CwHrMJLqMfaTlX6xEVpYc9b+sjVKiEYU
+YVeWZ0p+tkhXW/0A6IyBysdcx0XU9S1OWWin4Zrd4WISr8liiyinBP7JXMVkAM2TRMLOAF0vbTk
iMd/XiZJMjJFor1UsgheaMijcdelFYicDKqG4YCk2K8rAPFQ0/A2PuiFOViNDWrZ28SJ7AGrRmK3
Rg8FFZfDxkTYr24dS+8ojGEyubF68GdWpfFtuCRQqPyNVtkn0XdPz/bVEb5hRPTUYWujRoe1IrR0
AHyjKywRNkLMxxKd9ExB+XKfgvHH4/d6w4DzrAMGjlLI+MuYUsFFV+H3VuA0CrFyGn/6LCaCCEam
eKEBJ/bHdBdfIbmfclaPBoY0rNQByE0SQ0o8PfYABBw372IVR/Q4qQTYwPt9PKJVedBlBIGrAV4M
HohGc4J90wwF3zR319hwpl5my5C5aI328olgPRU/iYhktUEuILpMqptATis6A1V2OohXMPK8K2q/
091kmdLnNPVTgPvTlTsQ+mWDszAKuFbXOwwl8eIWloisxPnNcxqBD/j9WK8J1AFuOHyTL47DXWWO
VOuucUin9JtB2BlBBrbrPknU+iAbgvOkSiChpJh3GMOaJDLfSQQGtC7JJlbgzA9na+JMitjkKrsv
GbNZeL+lq2jCnyaMH3NQY4/XwsY+UufS8EPE4Lx/Bps4On6wrVTcLZTso5wDDvS8NAuTd7MjhIja
Iv4Qfj9TCezn4wXe3kw1tI2TIdn8w5o4KkKnzyUhErn+Th7Ow8Z6pgdd/uWldT/MRvSoRHbGrpIU
Os5HM0CcaBlFqFBPLCD1HhVYKpzh1JYvMVjA38Tmybq4V79JX6LJsKvwBhLSeAvmErX0RATSQUXL
p4Ac0H1YdkcpIrNxzDEtVa930WVBaCd/9Qa0abcLCQw5t977lDuCfw41r8h9HuS+hjA4B9Osar52
R1eI5aDIKHJfjVmoDq8Xjx8Uixvhi7+odfWOfkEN6l9g/MSItPACsmwmK97F7Q0Btyy3nRUWND9Z
WkaQIbztdCGFri0x9KzIc+fJRej2hm/54beXXfXrXO2TL5uRaGTFRI3maPJHnjQemqyYm10N9dNL
QgmPESIIWvnF40WWSWFvZk6O3OryuDFvpAn1IXwGVWD9wohF2bhFMYeyRLCI7IpSd6YWNnUYcGyv
ZLcjw5megivtYNb7rQ/Fgyvc2wcwlgnlHOdMTFAzZRKhD2nHZP2IY4WPZSHMgr5X8ouY9upYsa6T
2Kp9sVxLA8OVLvUhB/3VLTiW5UA7u2oQYHrpkfkT3HQos3Z/CFTN3qzAGIxIvK3OrmngttdZHCya
JoOv9zgVgjs59lUPRKqgaqi15Q9hL5LW+4hDn16Spuw5z5M28Wc22zBjwlWaO20AxqpzGdhaYdyn
SQGRHSK2ZHs4aNIWBEwbomY67mmtO1xwATvtszAjmCvVS7FQ/wIUbPSGU5kbvUCO2L1QGC3j8BPL
vCf5rTYG84Ln3SUXKyeQu+RQj6LDSUfTjv4bI/iUW7T30Fv65+UL2aDdMLv4jslQo3/3YRh8aSLt
lrERcZYKgNaIUhQHQXNNbdZUZ3E5tPflIpehQKRzV05bc5AVn0tb/elDLcaZgRpZv7mOAFtGodnQ
xY+pnosRXjO1xcc/ngBl8U+yB86ywxhZobyonCZv5AqEcWaa0ia0GNSYqbMlHXRgu934Phdknpjr
PyocV3bw0tP+BOKdD2/ip/Keoii6zE0Vm/J0tH8y5EmSLjPfmIn3oJyRcaxLbvb1z3shd4Dk1yyV
LkJTGdOxayZVJqOVYLlTwEnTc8B/K1MNyCC/rPkdhprjJcX7E4xDIfQ488nQlgdzeZRFn89lem1Y
ZFiW9WGskWKEAxgJFklnjn4sjExcvlPoEQdzIgzoQ7eeHHu0bYbdmFtpRxf6zRksDUmaQZhJh1Vp
5nbhwPjgJzK+0HTlkCiFtja/6p4UsCe6AfWnv+rNuCBeRHNtPYpi9tQtCEu8TBBy48Gpg/N0XY9A
8DSIKKZfeBUfpaTARFG866NoUNwITY3D8T5c7aPbxIbyT6JDKv1UnH9hGeoQZ2FtpudX93sj3Clr
wBaeBU9OQuAq5+7TmOrTrBLsZ9qx8d9R6o8hJvAcDEIezKIhBrF/xcce1MFyUh2qYSoKJvOv3Fur
oJ/ZNRIwFDgfXWxS0vUakS5FNQXu0f8yOS4Uw7+RQZ7NM0D/85vXrx8LfIfv5jHJ5FtM37OgaurZ
IpRhuJvhlL41mDVVst19dddbwFyb2kwsNFBFafaUzGhwBDs7uWTOeGXZEy3WamKz1nppILmJ29xF
XCAb+JcbB2xAJ0BVtc+tXLE6dKj8HWchdBSBSTBmkSP7CW2fu13CRwfEvjr0J0pc2oogH0c1A9PS
A3uq/xXn2ks1/TBgZ7eUdcr24M3pQd/8P67lHt6iDNbPffWq2TXjimqmGBQlyB8zs0OciHxZn/0z
Kb2SfkA12YB8VcC1DzXyCe4ZH171OLVWCCKbRRbxg7PqGz8qItD71D6HsZHFpSTOsyZmEM5YTELt
lWAPD9Uu+0wPg4IkThySelyLC4Lsb6s2WTNlAGu4ANoBfhplOQEp+1+wjTDMh6Xa9Q3omBBk5cPW
ukZnI7Dc2BfFdhm/yMiw6thlnXLqo6wF3joxuA3pxuRhPYpyazdfT53rldcEg7C/kIk6Qmha2nFI
JiwyLxUt6qDQLlTQdyvckACTD/bD0f4mz1z+fJsOmsll6YdK5SKk+BPC6a1P3h3wh6+R5BgnGJfL
37I5jNLfNL6KxBqkKd0Yh/Hz17t4YVEyVSQc9a5wFsmrImCdM4A35itxu3a5dafiiLa3epEbl4ND
jg+Vc/67Fdjew2CxkmoOUBgpI6vGvhLibVc3V9sJPAq1ID7h4m8Ne1FsYlBh9tuhgo2/WAFo5VP4
q+qEiuWxUlv70WwVlQ9yJs4m23ovBFwpmkMt/rmLMuXpd5MbW41aXL7AvTy4pcVwxXZGCpqupiJW
rWLqwouvjzcL9QsXEDWqUPP06hxv5pqPIM4v4BNgaU4Q4kVRu8RMFHllJ1JOgsB25w+k0KidApMM
O/PwEFfskV5rzaHpNtRP0fdUHszaxZr/c2y8A7b3HeshvwNZB37TMVTWdy0L5CqaHHQrT/wljFZE
3XOGkRa94FZW1YDuGBfjsREUL5lG+e0dJnbDhdAnstS/sFTNZYjG720EjRvTXOAK0uupJ7uJKwGZ
VS/A0r5pclTx2M2DUEdLRHLxOoHZG5Em054A1o0pgTIoG231Axb77Oifvswkxem5zu1BHllsA/sO
3Lj6vIv5eLgDAF+bPIyX71RGbqKfdu5JCRfDXV+YyimS+xPo6OWZGmInkBn++8rPPcBiEZvtqFdO
MwMYFUrRRA+3J9X6q1frNw2oxj+bWuNBYmk4wkflCPri+wDyEB2HpWkqXuUOgv+maKzMyDZ63SEX
YRenpfwI0QPiRF2PFMcZYcJwkx7YzG9xtYaEdTGgwkEyqJh8hA3+Jgfba/Ezs12VpWAvhVPfpDJP
3sWaITR7U8BB1av2K1v34qC6BJpWKz5gj3y24LFEesKVWX5qWVzVcYnZ0dQ6EfCc3MSve7JOGEOj
nwCw2pglIb+s2x2eoL3UQtcV/N2j0azPsj+JQxGbQp3viRmsrBl7OCxFQt/jeRsLToPf1lpKI+mg
8E6o02HJDRQnHFIJb8oH4t9pD8u6GT/VdwN12WqNfmzg4XumUk7jTg15R2H0EaoEsQRtxTLD41so
OizCdY+LDPeffDzGzLemfxDii+B3YN7gLzSLQmhubVvk/EzkgbXZtDHf9AcuJcU/dNyK9DckT5tK
gwrIvd7DiMERDAgJfFwS19+eA0f3mqyAXJLKBQ/stDETqcozpH0A7/z7ic1l3PKsDzjMYDaEAHQy
hJunTnhv2XO61OEnnoixFmYOq396O7NRh0xlKiCXISTs+/wZG4zFyFFnDSaZX/zGx0yx2x50Zrt5
XVtbAISJkqc6Tw6pxoYGCEOWRR4CZp2bPvPELxVf02ioo0X91Uw/DNpUpP70ZIVddmpJZ/0t8Ivx
ErhvRhct4QobpkS6J9jEEjnPpmF3KzRYGSRbYw1LmyNcdHgvRBX/ckXZD99xcWcVYPo4Eq03wK2Z
Jl6c1xEooxU8wIltXjCjy1JD3R7QZ7KyJmorJOFHbGgOjIGyHU4dkPsH+/hTEO9zuW8ltOZdAkqD
bwveZSyrwmIDpNsyRoPa3Bj6ltfJvRBq239bo/4c9LbLRPu6huTUU0STNhwU9tXCqU5L52XGwdrX
sH65uT/QOFj2dmv37vRjdhF0j+KNk4STOoGptZg0aioUNuBHF3kutjkI4hX0lgVaNTHF/8VYkIU0
uv2rjrdWBKxZGxU+bBzgE1+vMYwD+P13s+fx3FwdLUpei9+3sDjcu9yHdxpM5gxRUABqyeoiCDzU
gTCtEuz9t4+1aMO96TzexJptCU/nwoaNYd6QOjZC5m1kt9P1Tk9XJW50/rlNv3qWKCZ1YKziRm/p
O9/W8ICrbuvxfXv2qurBU0gWQp+g4G1LJcnB88UWLeD6W1ALNdK/jWGFlqf8AmeDnVA0IQisWLSe
WBHdHIREPBqHI1SQ05LMVz7l1o9kzaiX9f/uF3QhuLdbWfaQ+YecTKrrc2Qqkv928HCdE3gF8eHB
lo0vuRLMSl/oHoIutmARG0YtVKbp4va4VbD4O0612/atIclJiNZRE33yffBZJV+Q78+xghQumWxh
V1XIL1+7YdAibbStV1vA4IT6O+B6z5h6Quu8vQO9bZKVBvYWN9lNacB4G7cbZSrYdSP5vyz8LyVJ
SFay10z51KqeeuSu1y4x7ZRX0Jdl+8P0ZUMVT535RDcM/z+NOyWsAC8EFzhihhyW47kIAruCCbgh
DZhfB/4vABioxgFKS8lUC2dvu4E47L+Mbbz+JRCRbGdQLrdXAHgF/CaR4AI07OW+0tz5fASH1DBf
skvyn+FXpz9JLig6QsOQthuZSJmu/iDvbqPkDE+ra1MlCSyTwVRQDJ/5KGjllqqdt/e9+XBpaZiF
VgDWfR7AqjdqbBfo1ukK6lw13kO9vZ2ENa9xxqjEchYGDr17kAuzkeCttWrh/SeM/jyHT7XpXl5Z
f+j78WA4S6QYuENKsap0QMYzzFiA0Jm2/Bqy9LnB8kz0UvOzZpEN9jY9w4T3WXJ0JJBBtlK8BWCD
Hz9hdxY7vj2wX+dyP2qVj180uKLNVkQihMSNw7TcsNu7o8/To7S6XCZUz6I6P/JsdcRs3Eahw4+V
XMPtfLl6OY4LXtIxde35ms1VEoy4BWChTELKUQcomhYtX3T5J+l4kvPAGtXKY9BPkvD3CPge0RBL
/UCs8HhgsnEQPXyDAS1X3G+FifeCRkgelZ3w7BuTkaExJLyT8ORBJLhIq7RBPfSwI3D5DaPLBNFz
+qzhTut+jomUSd/39QW8t6P84dgDPdYV/IT6glJ+ARp+0JlGdgzHzYZlT3nTtsy+cYZAPVYzJhBl
F0dDzcicdHO7n8sqWTP31UWm+YNBcbZRwU+jR0yjtUkm5urq3PCiADDFImCfvj4Qh7RNAa3noCmq
4QdvgLP8uw96sXVQyNvUH3p6U0QPS5f+flUYJ96EcYVV79Vyl62sRfNZWNHjzs0BjMezOnqJ+6nZ
rZy3lYAP0Ap0BqPCaw1GTv5CgWuof9txc3x9TpYB1EbG58LloIotnuBLX+pZ8aJ6TAGlFBGrHMup
dBqVy0st8UR5md/dp2Bn25W87m+BT+pHxsggKbGiDUeL7ue0Cu+dg6Unn11puCi9/WA/bifcOM9V
FaWUgKj0cJVQDw51HoM+xEGNl1aXJRMDV7wasgex2eTUw7Z9LSdnUUXsdEOpq7GTenEBR2PS/Gpv
3yAYkbYjsa6Ts3K2bVlCDXQrTUh8SzeITbA0bCoxBnHWXhOpjzWfeW3h/fHLrnES2Wyhs3VhQWTA
hxt4dMz40oopd7fQLL+UAgpMKiYSgZJA6riX6SrCSO0Kigo9iFaS+iGAQVofH+ikIcJClR71c6Ss
O0XeqPdh1zYY+nP6+Z/yvyOgHzyoyl9IjabDFPqOtFEECNb4LANu/mMKmeKg5+k3FgvuSxzhikQx
D7R9S0kKBkjWUEZA/ts5EESe35SU/pIZkLz4i0Kt6RQOQ3gWrb7QgD+NdtVAvwqW391GdI8bcBAD
vOckfuN5pAGDimMkxxYd/mdb6rhvwbLbWOFjkMoeShnK6gIuadjlTCXzfrDZPMghJOCujRgdC7Nf
FMtKrI61OFjhvTfQ8UO0788KalR2PQ5y9WBqK49C6syHmJ/PSGKNvjdRuzs4j0czaji1cmbsiBJ6
TiNQB4uIEzx+dHMx6inEEZBYnzIZXwO4biN0IB47Hjye6bfpHPLqhMyvf02x4nR2hsJXBnHlbH+g
Eg0kd/Qns9jcB33zOQCRd02N02yGTNDZgNlxG8zstLV6wxg+oZy/rhhg7q/KR5MQgNIdkl9uvsrS
LIVQ9Yth2JIKZNjqJUh35vmM2YrRViReS6K3kagXOcO/NPbG05GOOEahmeSOhICZlkjVgD8f2hPm
J70kYk1hVIf/wOcxZDO1T/X2gbythWPoIzUjL523B2rW/o49ryW/8gbjQEPsMe7u8MeP5tTUcg0i
nab3Ah1zl7M09z26eE0GIw1XHSjb2xqcLZlDTASK/4P9/wTJ0R0BQsgFaUaymlzHUbT0uSAFXLiL
MyfTC1amadT+ByPc41FcygAQExTIbanVUl9wFevqEfBRTjw4UVh8HhfexoWL96dcaG7EPcvAwyKt
2LTGKKGUT5vpa1ybB2aoTKu3lgonmmjmNqMn8o4wH2DPT75Pri/Qu8frdBXok0Mer8UfNQ7nTii/
k52M4mXAyWBE1wRYv61ZvXnvCEPKstJb66pQ9i0/nmXQyz9bBnehvERiPqXWWVnBQd3sZkCFaudo
ITtcAvoDMrW1FroqVOn3+wxr5dQLyPEUf0fJEdJREoO7hfJ5PB9rmEKajJhPMbgvc+x6zYDLl1Oz
od6mY+sFMiIpxtUJkCD7rRZdantzsk6KmcyqGsMbXiCTnc7XblRxkqfw21L3uwsQmSQNEPhIC8fs
e9zJe+EP0HZxXvRTioJEuhvtILu5n06eFIdoXWaCLT66Q2UrSxb3HqBf0wUhLrhTZGAcYTPkTrLv
9NFgA9zvgKQpXnYcvvaCILwuByk9OJlOq2MxOM85vIW8L+qs8m5TryVnaQqYvAcaJ2TgWks6aRLz
/tT2fVKCYJlvPzp2Lt3nNysrtFOMVjaH3n6IsPp9xJP8/CG82gJUENcZes6NkAgyi+UN3UCPpNkd
hpevtUaoWUGzzYegl9r6vKfC0B426lTnbHUDUXtEI+u7hxQDgeakftMW+RwfOZgj/vv7gtOKOVpI
fCf/++Qeccul9igF1VDQyE21i3hvuHEqXbAPgq8WxuEqwwA56RYS8HyGt4YDmUPbRKZcBO0S7jY9
eMIxgG7E8WzDMrstZ+cpnwTF3Ww8xXviMSKMGfdP/c4YwUvKmv7VSAi/OJGC18rNZrCH7zkHHy42
X1k0tqlzPuCdm3qmq6ClkArDEvV+r852iK93kPJa1I7IVKznZY9w/BcrIEEKDJ94e2GQ+/o6bkja
b1YRNegMtbymJZovfm+KW/tvQm4U+ayIjgz3SGeXje46jaVbLoug9l99jAYoIwu6ScascGtoSe4H
IQLd5DGnc7eQWRC/QhQhpf/nt0tVA5OEnm7FSDqFmTBknQm/emXf7P69ibFiB+VtO2Bb/2YeawUI
4XY2XJbLCj1YvvHXhhS6iz3qe+UMIAEQ5ir+x6qSxDWtkP17wFDbVxHvZxTrdSjchMmKdVDCDScc
uiekY3OcFW/HuxNoYBcTSWh+SvkhJImTA8QMP+sjtu/Cz89mrHFGWz1xcshM0cIqL1WY3GPv+g98
bgcFufQUdOinxkeEFTEupphjj5kJDwU7n/7RbxgNV1fz8oTF7/r+iy9Np2cwtv8fsTy7iGxkaJwe
NaSUJuen2BNsidJQQgJNbveq1WSRdv8PIVCZyScY77Sd8n4yw85/Svooj7tikwqCVMSiNVNvRsJT
LQBUzdfqSRD+sHzeeu4d7qvlDWEZkDVO/WbiYZl8QlLEcQeju35Abx+yS2dYNSHWtGYTkA0jTDLv
k4tqG5O1u4PAGuhL7y+kmka9FnbwicQHw/IIoPvGvqTsIkXafSqxaNsTWZi6SD3KsGsRz+P4bQNX
BfyFk8C239Arf4tfyUPzXjcPkCIpUDOCc32L7CVrQhDV4glRMuh/LLXTOvuTdbhmxUY04w2oZHVz
b4vr7eCJAJz81jm34qBm67XsBOi8NOjJX5CAHomEgu+NzgIJxEtHgZirdhpMAKugiOz4T+j5YrF+
CwR8Ppko/Omeyc+w+fxj7ytSznvyu89U70qb5EL1R9xtKxZm+O687GVe6YKIp0iJh9hR3waGG15b
VAv+Pvaw+Okop08Wdz2QMYsPBT9gVKTdgM/lzhMU8d61bFlKxRyWlsv0ZTtMRYUN52Z33AGFzR04
6IaR1wRQe0yeL9YJOzhSbqJ6nbvRM0YdzvUGbjv4NVmu8l/qKOJPIrJJwC84IRWB/c1Zuy6jsUTs
ZOQeyBloeYVU6Oy59wqKXEbb7Z907WDIkhF5jDcDrt7w0fqzirXDNOw7uxy8YqIC1XhiPLE8oUvh
uEf2VI+IsddpxM2UnJi9HY58vtXXLT7KQNiBuq0MslQF9P6WZ/z/pS1ah3IoYHWUSOwTNtUHjSbk
Ty0bpoSRzeYTzQeMTCe3QH0QiJR0IweQjuCPRXyh0TBtFulinmTuZNu3TV5wjdwMlHu//mDRDLjR
Wdrao08POpyVUrgF6W1utaGeP9mN/wZbJjoIlkQxgdRGxzPKyFPsDAxifzadgoOe0dqtbqmY0/+c
kHLIiXZeSkIc6CWhyO41fhF5jps9bCDopbHLvraw1lNw7TXXPaGpL/X3T8oKFT1fSDzS9OP6umjr
2pAIvUrdfuC1vcH73JsJDgzM8OVh9lNJ1RCllTQuAL5iRPnE8E6e5X4BMHTIGsDc0rIk+A6a44Jc
U3fLaqCR6rLtn0n7MQrx7ggLa41k5GtI6T14avV4r6V8HlevXnp/Y8nACPr9DcJq8FC58fBBrIq6
vRLYfuvzDZK6nB0aOtMXHhQup5pqFAjOEX4xAZAzA9ULAY8SXOrROMW+6E4DOX3vlGz4HZP6GEP2
ViMPQQOYyA9FCRqzxhtAiVndurMxW+aeKSTrhoSXBPmuorSBqb3ncAt86MO0yRR/AWTlZpgT6GHq
o10VEXAq4bsAGhZdFkM9DonA36yK4BcmSo+AIl9a85YBIuvTSKbfuF3fUqIuB5NPlrvvZssxoDNB
/gVem3PJHI6nYKQWzcpfxEn+yYC3LbNmCeb96Zz7W2cD6NdPcI/qVxmAfsJ8WRCg+3Pv/x3z8aBq
tY9rtiIowTVjeKJY4vCIO6kiahDUjRMK0GODcEJw5kszBkduR2VUT4qyT/wAXgboEdS2G61qFKHF
FEfeq+x1pyVCxuycpxY5gfeH46HFWNeFkofu6jkqhDF+lykJPORZ0NWltkrpGlyiEs5jSu0TDQwT
Ljq3ekftF/wfFJ9vDchNFxgduLXF81EdPLmq1hREqBRy2/ENVnGRvhMa/Zs5ynyuUfRvFny18I3C
XgNYa8P7Nq40LmRwzHKzWVffoE7kaPTCQbTl54LsJmlbKWZnA/BiHZ+0NGAK3R+H7xh0ZuSSF0VS
afC+2fvIdZiy+wbW436uKSGku3wYS89IjIsWh2K64K3p8htOpsH1Y7akutQY+VlB0oAbSkOd2whD
0JyVg+vZh/YUv7ZdJEEltOb0N6CiCNtG2eFgQU5VCklE+L5D7wHc5OVOB6sWk01uJ/+885iPzFHJ
0tTUzZ1twVlTB5p9dVJu/7d7y2gmZE2J/D1i4BaI4vKxC4xM/ETpjIp8aAFDAq1S5kqB+mI7nfx6
N5Y9uuo9dOz6GTsCyLMz+G3GdBR8thI5Sy4UKfO67LSZjKBBYzoNykgioKVTK1Qnbzqmmzav9mo8
gCwZnLb8V24MQ1gnuY2NOfyxhPh7O5QoXaG7BSqIrhusiq2NZNDAc2uR8z8J9Hns5mZu2AfyZNDH
1vPR5L4GHxrasmJ7DsYqIeVMDGv6EdHreO8VLpFK4nKSae4EEUUxs3P7mOr420/xPoXbggvpTPTr
mruvYcwSLgDXACzgBI+t2u0Kns8eKDiXVEXIAFVIXKZiXgtW3hJOSHh37FLkvQ64638oeVxJdbBi
pcWHcF34L0P1KSvh0O2dviUqNyzKS2rf/GF+oWdXZT7tLWwBIdII9I5KWlgyV66HTSQl7oeCX1He
rChXRMLoG+xs8XU4xUlR+s7LGq2RMckLuQBJowMW5o5oHcpJnEb9Jqd5Puqf6P1+k1GdeeHsWevO
k9oJK3jch62nG9s2zJlBPZvt2zPWg+02oHm7gif+GEZb4Jc+kSvFT6LR0rv9UlsbusgshIoJtZzi
TklzzvjmPWNWhS6t6UQiPDJAFc4E1pSc1X8cHT4Wr4Pg81X+qx6DhZ/LrqTju+bptoPV94xZz6cL
8LrjWFHSvQZhCg0/UpWYU1rvFclnXgPO2camehGE99MUN+ivnIXGKLGGvzwI2Woq5VcAoo+bcQ9j
By7JwquLPBwqOaX9BfeTo86E6tL7fVIUIbQJwFmSSl+oK+Tl0/QxQIH686GC6RK0qN+yo6f03aAf
UxsFpApH72cpDYOKfQPng6vgf8/BR5MyUsheWbnRaSLHzyJbeVsNEmR+dXfroV6yn1YwkpyuYtFb
sR+stxXLQifG6K08VsDH9x+glZ8XNkWgKQDR7uYs4S8zMepWmYdUl2/VaGWJVJOvW8PUFbnlOTPy
U6BNTSNbLCwG8CKCKV971pyZT8pGkg0+slzDLiF2wnHXwuT2QfzIViFO5F2Djq0Bw0OlVh1wxMny
n74JJfd8HPMhiBCHkyw3CtFG8DRV7q9tq70S2fCaTVTPGfQcO18Luk0GXgN2BmTolkO3njByJotW
VJhKJbzNmvOlulSbdLlSXrXqQOD5TPnCX4H0wHnlZZw3in7w+hMk1mRgpDzR78Ul15QCKbE+csZ7
cFpip/f3e8whFaDzIS/JvJPzAhuGqUKgKi2JJtfNnRLivzxIpVrCzuodcRtZmeRnV4xNZ0gOskMG
VkVafWGo7snGQe9DynE7qBvDGjwfNbqh5AbxoSsU9npx3/kJ/yKBlX56J95vkK1+qUt7UUMq0RfR
RG4f6NVsRgkVsq5CMrkvsEy+ejM3IFmZlEii0NzCqgqWXjKXbLLdVZ4z5hfIeRlBLCovn0oexW8M
xQ9SjmpRDifCzNkTm1MVdSrf0E5sXIylz/xBOs+W0uHnHHI4zItES0LkODCkjf3msZ26vLm5S5uU
KVQrTytQtZPac1qcqVoqiP1qSfc1VJOiUfbxADappo6U099JDlI1t7XC8KWi3lGrHCN6XVcygLU7
DoSISu+6QcnOwdJ+FIslBMGFNuTZzNqhaeaJOxsgnsKX9OrNtyeh5RDn3DcA3qTXZ8XQ47DkkPHe
79O0oQkmb5OyUqh1Zk9crHwDHq5uIe2eLuEzS8ejWc4jfqe83+gD/5t7P6eTrnr2nt6XtIdHP5P/
OVWswPxHZXTCWY1+8pKwZNvq87ppsotgqoqrFl5FSBEGii8U2jWo4v6w4yW3TuKCtD7GXE9t7enn
Ky/oC2HG/1HTGfVUnN4PE67w/FDikNB02yCctzAXtIFucsg47JjealV5LpnJyL81rLaRdnHQwTs0
CeAOX/HYHca6NsAPDJ3baI5t8hMXBIvvf3dz9JkTuqMnmhn3npmp/b1BJoV4l4EOXECsHUiVSUdW
MBPKTF4RMRzAgzaBQdSzz0H/2pUxwS1Xkl+1BEBwdTCuU82Ch2Dqz3GkkcRaox76ApbWwmYQPWMX
11Se0pTPNZ4CO9jNGO882zjf5+ZGkW+2kflKtP50V/TPqp3eUA+Ovxn9pqm+oUumI2pxLx2wZxnj
6Sr2gUs08lxaHWhxzUQRqC84FSFKvBX1bSXY8of7tiyYMmXr9lCeGpxhQDC/uP4S3s4nVHyQiNuN
HfNDe9xQYdUeTxFm2eK97EWsAl5usvVtgqSuZRhZ2NHX9ck0vKP1RVitST4yJqRcBRnzmS1FgKQK
EuTQd5mvuYC904Dfdxfh8iqv1hW+6JgtKHyP8rJgR66jvLHFPqx4Oswu7xWdpnOdcrlLc60irBml
mrncDzu3zNmq7L98X93rSwAd/N1qftCCTLaBAhIhPPXFjYWDQnNpXpcOxF8xzo7K3mkn500v69pw
Za8MbZjwjuw3uXn7ORVkFjcC6qD1he7k+btf3Bc6FZaq4eFBPr/dbG365fo1O/Uuw9ns4M13BpSn
ZdpLNXqqUjAXWAszXs6cwoC1KjHo6vweekqwXFzkE61QgwotoLn8eZtl7tb3Jl2S7l7DdQNZkhL4
eLfxNpJQF09mFuTPER0C/0nsJMCEnsbb15XELtcxjEB7fyovjr22DqcYI3pB5SpD8VqHt4yTO1V5
zTilpGQXZiAirP0ntKKqAY3iEc8iQbZst5XjmeHGYbOVyC0E45QTUcCwEtHmdJuLT09pIRyIGqEW
Q/fXqGz7pGWorXY5AFaGkrqnq67PXNKKoY4c5eQ1z0Fpi4Rl/k+2SxVXLrsnFT6pBzLiykp/noiQ
+UU5WqB+I2VSldn+xrc7L9YBlcpoONTt9NXFRLdDr27NJoEy8rZJWQZcgulXWme2+I7stVUNtmXU
uYLLqk97fQlrV0xep/T/hB6WDffKdNfm8KNvusvs24iXCCTNYIMwK+8pmc1zs2Znlw58ll5gMhJZ
W0uq1YyE74i+BDWzghEckSynU45sJgVynuSnJlFPHZ/dI3Yp0yRw9le5Mm3atOVmg6H2X1QTUB8m
5d8zyNDsQ0/meYYPIKDBCU3FzJcaPaeUofGAJsSyEAvCQviBuuAxiZyodFa7L57/hc5cah5fh0on
J8Pu4hBnR/RXeky/IfWiyTFrRlIHZ9Niuj1ztAg58U9V4CXb1UcBap41P5rCN0zbcuIK5v5QSDnv
Fq2lDxjcaOenIyCCPwq6Zrbs52N/Zx1Sz0Dhfg4gFrkzywYYDfwGDhgfHY2SZDT0UHMJjc1ULNv/
BwxnmBsZiYysdq6Y6DfeEgO9s/3Ck+nnkpA9WI5wSURKa2Fli/Go+kBY4geuE1qO5Qq3PfiRblXZ
S/eQHGpiVA7vY5kaxprp7d1vR9y+/LWnvdzsYebB65/V+6haB7wgx5ickfzrf4O5ouYrMOwUNrgk
Y4vdHA4lv5s0Vpx1wk2gIDyyIrdmT/wDshcuKlSNqUzsRQpDpcsU7DzA5/GGJV83JvMQJtjyg98p
R2OWpY9wfDohlNm9hklMaEtSATwQy2bExmo8Tz1Ptgj4QlVLOsTQJW0NS8t88nJ/GdkiXoLJo8cW
YpuY0pCdQiQL1D5sfNflVt7Z7ovtPkuhOt/jcK31i6gN62IJKs8hX1ODKXp03V8MSiIoOxRltYdN
3qC5TbASPKsv49doNE7LIukesZMyHkHaJid+alx6RoamlaP0IoO+VOw2kOWZZvHQaAssZUq/DOuT
UmEApYbVCnidupzPSX3UwWXLrPhbWqOOJ6sz995kCM8cFU+lHEMPuHKW7aRJQO/yxPQOTM8sgVwO
4PWzdGZfCWQk3tkISjQD/MP3BjR8esreLhYdzRIT8PG7Jew/T6jBqoLcOUg62Mxs88vwOBj2NShX
BVizoCtZ5nEU4MPqeCBcBY0YATqyLVdS3tzYdhLA50rVkowsPvbqjJ4u/KbQgfndcMe2kNs+xnNX
wxuCBBUCYPhBonx+/+hneWwz0ClfI7k27ToRccOQ9KC/QzwU6gG5sh/N+mlmj7eAXVL7HZAxZmx6
Zqd3WZtqbEzvbLIm4wjM0Liame4OfKbvAKnYRBNnVnnMnBaOU5AnQYWVSz2PEnHryb09+ghXn/tm
fBjwbeqL4jh1bOk7/zWlGv4D6Eew/LU3UYvLPwg0g2yANkN0itPVSkmDQfdM6lXjVbg81q0WGv8g
qhm1vm5hpmK+GQWeydG1q7lCbmu+gCglUVy4dg7AQk8iKiRBeKmZe3dRMHyi1tHtgdKxcMK2rcn2
lXLbd4VZ3U22zUda+983q3GzbJZA+DgxZtYcL/pS7K18bXRTjCWi1Jvp4mysCp82UFx68LZxUM9Z
D2Skt+xr9TD6gkOOpS+Hg/sWfV267SSY9U4f+viuSzomLkV1YV3LGGLscLNf7KiDKBrnGMmK0PSI
rPZc/LAfJC0zYpEQEAdTzLBmolIqbf6Vgyh+p6+luIwvFsbIEudloCoEt1w0uAE/yCAdbsqOZFlo
yJjBOvZZkplqSYKmMiWdkW8+VuRtoCxj1ImsRwxt20HM7xieu+FpVmV0vSRpX3MPaPk8/J6wiQUm
Q6NDTgj/NNxEm+l+G1ay/pmJsiPxIqCGevdrPT8R42cj8eEWhdu3S2AU7UkGZaOOzG4DZHHQXkjZ
0FSi5lEBbdG9yr1xjreGCJNX41TZZpPTmKvy2lqRqj062iRjpdPBlwdKMUrEDsBa5HTE0U0T5nuT
xfXufFPsjBVbU/jKY0brTh7oF+sv741PhmalLPqYbxp5zQweVWkD4hO1iWE8TIndvlE/WYs1UMqo
bRMeObhv7epFU37UZYATy46u4+mN8lMQCO/PwHxA6f3TbOMw9yVMkQpfneRyWRPMcQ9aablULTRI
GEt4aNyMqy/DpUSf7l0TByZlCbUQxyYO25Fysfg/r2eFcvOAbWVnsbAIsgO7HrI9ESQkEIgT5+pb
DvHV/g/ejWfaxqslHXnSlY93cr7wLu0bZV3V7lIzk1bjAM2c0R1TiqpX2zePstFZoaAlLdkztls+
akKkOXXuyQ4bxTf4sotM8tjwIJh686NgHw45q2dDYhu7ge7mVL0c/cZx3mdxWracQ5IDsIGQLrcu
kJsUuQNXRA3HA4erhd0SF8TyOcqFC95wayVcLjSSN8W6B1vjXjEO/rA4hA0cS7T2eE4VGtofL07n
HsyxGeHmkqTVeVM805wgHz3ZWwI+/f02INsyEfa0ULBeqNQWBGifgJfB6HgwOlUP6vzvrORcGxy5
4XicLxA5J6fPWvRmdL4d5901X2JKP+afswDeB9gKneZ6r3zd2r3oLzeNdYhU+E1D9HZgMJM4p8iW
DEzKbZp/yKoltquUlRya+HTt51fHQwa1azv8vvBt6HJlU4AMioYrMyHwuGrQ+QOhmIG4wBpDawl+
T5wpuZEDEHsqWxlsuzHEez1BAuQYSZaMMWqPOnRFZ6VLLsIUYdlaj59BL5RBk/AD1rp2GdgV3s2v
A4zG+GSXmPDAiJ97LdQQkJ4lvOfpWBQeGwrudgr3WM4pQFaGw8FzMYFJS2rIsLb3zumdCxO6UrAe
Zpe1ywNC2lsgydJzNeli8/KTpoFZJANeSpxLcchJxFC0U4hWwRdMRpYJ59lQ0GN3TRgajcjuMVs3
tHDgHNZqiDaU+y4uVLGqHpgGV4GFcvPaw7YcOQy5ZxkXbOqpypUwQUrGS/6b/syTzfFHcgQi/vKB
cyLWaaFJNZynR+dst+L3mubHkffyQNvgjeGrQShoL8HQA9s4032V4Mdrsdf1gHHscf092WMYN8Z1
HjUNzrIvteWLf0J/k7MnP623UI6EY79HaATXQwMjiQYSaorEm0QN9sXmbwckW03exRQb7wTuBFu9
wzpgdxBgpdkVQBkPDOOLAMKSpyJOymM0tcPjG8C6LR+VOv3iux2Ly8TibOXqb2/NTOj1+pNezW68
zXF3TTa7NhmY+GhnBtHjjTYFwofbwP/OuRtsSV9c5LqXPFYMbedLdMhmxhOdJlPkr5slUHOIOd9T
Z0dlkK6uxmvsYv3o1u1kOOqpF4d8cD24BJ5dzn3Kfhq+5hUEhpRRKcxtH/7uabcQ4dGmL4DyyTxT
SquOYEQK9yNezA3YaWXSVFm9IL1csKBb0pBuKylIrKyYTvbnHRmDWVuVMml/jlcikVRMrHJUkKO6
kkFG3XmOAuLLVwnYlb3BC8eEcS7GS0WaKNhwm9RcORtUL6kYwyQdM4e2S7WibCSIYImFxKg9LqYX
n9SsPB7lWWIUgvcHmo/irgTtHRrTzkk+jjH4Gf/vVyxvq7f5C+6Jmant/vl7kgCPYrBJnqhoHLDe
eaxovK/DHLJj+i8TuL86UZsHNSdkLuUwhDVL6qq0xpwqKKZ+R0FzEnShVQrTG+aJ6qtUTOHVgHnN
r9wZkdHB8QawWHRCVWrPkIIUn05CSbZUw0rQOWoofNdNJDJqaMTQMv+FgecpzLkgJMYUSlI2KW7/
8vC0pi7l1FM3HOfkTo5cgA1K1926xWFql7fH7Kjn/by+GXr+SphMsliiYVVPzoHNOR0EfHDQl+XD
f/v727dNnhsetnzHPliMF7MDDPOFniqsb/dEKW3dCpu4iEPrBL+MQHs3Z7md/d/wN7gIbwYvhOVA
ZUICyvkypsv+WPkUiSgkrN6XigVJ7LAqWtYOYkj8o6qrVVedUIDIh3DT2VVHnXSSNTJIbsW93Box
rqazsaz/qZ7L+VSm3idji+HklHxheTL3Me2nn7yfPdP/PoPdy9UGh+bexcLRlc3dDgXUWWjKmnlm
ok6IzAyDvvyxteF4MZ+IRKHv84eS9oY7BxqluteXOyfeuXCjhUB+h0H+r/PetCW/Spo9dKxYL0OW
T5Lvps5l8wCanRuvTdca1GdLKCw+xKQ1/rbt+qojutLHjJoUmTpgC3839lpqVmxLBcqT1v/Msh2U
n73h7pDEPXRSqXV9uM6dYFtvNhI/2Ig6RKc3IxIr0bq2AydtT1+pZ/+syBrDE6ZP8aCRXZSxLDbL
yaGC3KrkJ4DC9Su97v0ZkxUQlwB3qa5yNNLpba6huLjlF0zhqGCSPj/RA0GigOoSHsU3g//F8WgZ
8m5716PBy74O3q1Hzs+cmZazvq1D8mRvO0KcOsJbsjBMqxXxgZeqMyHZkRPtdxQfYOidyc9ZGnyO
VZgKf8Ki2DoocUuwXFakRsvYIVnIn0n6yTJJspT8BxD2/qT9ye/iJ4s7ECuU0W+VPwbQdaJftIBO
2CPT2ul2SWGg8MjID2s7lZa0u/3PXsrI4HBEyLKQ1yOYbeLVg2ToNBaWiGHr1XhdMs8F7B2tY1es
tfxGoxHOIFx8e7o0r3JC/Thu4oMxE7FF8KjVdrMz5CdJdc7vinaYsQEwgfiu2MwBOY+ydwy3Jspn
uJTMMqvndX5PWKM2MIaPUahg+hy6iaSRdejkbyS2lF0FTBMm9TMp7ZLoU6jpqugeTl5BxMVs0kmD
0kY5E2BKaN15KuEdbarsKR+tLuW1YcP/MzgdENthQkEtK7MNXE1SRR8HMVwLjUz3Lue4uAd2mP13
k5xAryWJVCgWPRKE1OcyJHPp1RC0rccpb1aXImsBQluxGL2Rs3RNGn3tIkt54amIuT+l453OJyzH
k6D80+ajpIwVtl4ub6zG3AcgkYTe1UC2VV1cm0oyhsF4i/sbicOKxIRAhL840ero2eEU0DKPyCSQ
7Tj85xJHHqtVk7E9WbwnkAYOPnMXRa3CHgyg6xXqy6BG2iR/XvcoQvRWi6OkkEE5MLC03VwJ/xbf
z7P7AnFpFDPo+cY+dcshFK56Um1hja44k6HZmGEIQP2M5wC1o/bZgYXXC2YClA7wZE/c+Sj0lVaH
Jb7KY3DzTjGTW1cmn8D5RZvQreOiq1XA7cG+tENe+MXqdIPMgaG0tWgwJcyRy0Jl8P25yGya4jri
sSqNZ1ukx4VtIl1q3wmxQlEpN4NvEtYF3m+843wDDznVnQqxvBbOWN5ylzA5OZFufDJVdFq5pPqS
XIB6jLmbYR0GDYjLMT7T+9vcb6wSRU2Y8auq+JMEPUadPUruX7HOt+kTjhv/ZWMRJ6rZlLiUGgHQ
cn9M2qO5BCgW0SB8e6PZeLvrIxGmaBP9FOOnpoiEyzNSsjWc09nFXETd/1tp7sosoGLSg6T1Xq7Z
BOtFmMXuY7qWjsTCd4xd8xI1ho3DPP1MOyf5f5dC5a7wbX7691bZ5aTC/p/ejiOM3FRWdyXwJKvB
KEWhq+3N48li6QbK0E50cVBK8t0NN7n9cRJqnPR/WcPFuLurUYTnmGagxkJHuNNucyUtauGO28UY
NkZ1dxAhuLFoSf2DLPjwTwr1UOkMb7aebMiqM9Z8IB5ecZICX7+R/qmslGw7qSn3rzO8H/IPh3bS
R2uG9VYbic841h5RrnjXOEv4c0/aTJWkqtqLjOVR4kQPGnFd/nLRi6NtK4c3UW3iyvyiPjjzKD4O
8mfLCJJJ16xNkfIXgagCn5kQMVoWYQqBpz4ZG8HD1R4vVfIGaprVQb45qmHhfmD7UDKkrPhH3kpn
J9N7k40Y+G0SeRyBwrjoRhpTfZsetZFEiGMAt7fIU9cz7kdVGKa+tlaWMZIDuMPn0+5oJnz1OKIL
rmrA6wzcYWITOwwrKCbpzIAgooJSSk0LGO1cCvUEA+pcsKDoKZYjSHoT3odKkZrjuGZ7VekQUsVg
eNxmt6gia29P0xqIMmgBwIRznMvX1HCbS5zlHhFkC5L8mqta8z1U3nHyeNqBuiAFup9j68Xp9FCj
xGvZEqtCgPSK1tF+INbt/+iumkPm6LhNExo5/JQaNUFBXOCcuBOJIOtfmKKZI0jioFy/UIuEBnIj
qsmi/4IKj0Ewd/BNKII6DIbgEwMkn1lRjEKT+sMH2kiwiHbzGBmxHQXAa+AElko6/jjevnTXxvnW
GYYdRH4FV+g4p/OT98lhUPll8dcXCfOdGOf8JZkoiNIc+GyiZ34m77CO2yS/JLSuDODX/MxcWknw
208fm3QKT8j/v5V4wGcgXG24QEeUcgWM+q+/yzC8+snTpxa0sttyzt1ZwoVM3g62GUDBo1oSR2zR
p+M4ki/IDavryetYlaocymTwCpCY7vIsGgNUD+qnnPItQq7ZOSSA+9J55RTd3wiEPmkauvvPJ203
g1GJKLe8XbWuKNzTMmOKwKEH/bToHasVVxs1ON/zstTA7tfhgZ7I99mQYnx42Pf4pcZ67UsNVmCz
U3dT2EfkkDsTJVaot3o0f4CHOeT858BETd1xit6gaYGrvL/pzXPz/D2A0c60swWd1JHnKj7fxFo4
fxUC2nnwQnxFl3uxOMvH+TiCfj/Bwzwpps6svu6UXEcPZMwK8rDgjW68EIADDbFAs6VFlq4Tmy5y
/auavDSStmW5Frd77BLCSuO612DwDtOpyW4UP/VJAU+M+veq8Tfdob1Z7tLc+0emMzrtKXQk2hta
jLr5B/53YH4tb0JoPCtjkEv6LIouPSyQSqUrk2dP6+Snc/6e20L/e+nZIoyqOeMrAEDGVOxmNP5y
W68DAvP5+sBQHwAOJP8ti6M5VrB6/ccxtlLY+TY7IAQo5dkb+T+FE8rU4pV5tL0lWFVDlrB0csa9
R2mV9zWwc/tB1ycUmhFyMPe+VHceIs25vymZyYVf+gavaViexHZeE8r8mLBP5pZfi+2kBb5XiRES
B9kq14q3S4DyRlNzhxSPSRK5ezl2ahlsRitZE8O8OmGQJkgWndrekkeIGbHbMPeNQ0K0toi8kY72
aQ4NF0D0eQ5PoK1niuJ6skEFIo/Mbu4lA/Tvt+nxv2Kvvqiw6sbxnmFqnu78VJ/cnqCu2EdgPH8B
XgchGEI56ityPaeOjQSh59grKzWkdarWm3PcGw2/a1YMdQ/ND72PZyhI+2quOXQdbApr4+8bkCUD
xIgPMQKzZoSdXzeOFcK+v7nhien4ayHxnw75E0+oA2I9hLjFCRj3aPb34v8SJta1VoT9uNbdFaJP
XQlSxmZurxE+MQhD3+DN5B89dEASeXdukKOJ9J1iHF0+e1NcoJAgyxl2THm9zOkD5ZUAC6cYjMDm
PWwiV3hf/uL4kxOFroHhftPvN26d/Po3Aa5PwKJTdBPaZwjicaz8FEVJALnDolz/Wi9vTsfcNJs2
fn/RQkxFe47EncZnwxRYUt1CTE9XsoLY1C5Sj/mYuxBvApRUEYSjjgA+NPvGhYZgIO729ElGuTgf
1DN4D27MCKc0/7JRmvhI/uI3ULGpIq1RDwgPwi9X1fUfFjOD3aGRjz2aBSlJz1HWcYbVrpUy4uUb
GmclIwU5GlQ2A3Nl4F1CyZgYbe0tXg/IY3mOllGnehsjsPdajN0iCUYepp6VVmlRm64IyME9rmuW
0uCm+tn7lQ+znmVEftWaHT+O7Ew5tKf/7EbOgyz2P8/JrfKQBfUKsBVyyNHCl64Dtz8LAKfmZbdm
uwWWnZkwFQExgudWzDKr5GL+6FZkNacsupgHUVwhtP1Dt9tBeBAj12gij9SoqwIplm2z9nYS++aM
56lPhdMVkGd5xoh8hCZTIiyZAjGYX/YqRZdXdxjbMEW6WLmdhs+G0VU46GLzFDxyE1nh1adSAx44
DJK5MLPDLk23EbGcmS0eikQQ+WuMpFbeNfiPzAv3D6M10oSD3GSJBce04A10FfdnfvA0q53wzmyy
PI7TgmvIJG/enY9o0zRVT7fsyWdukrB72560kN3pLRO+RlqPokChHN3Hdr2DSfR6+dOYk97MtbzU
mh1ngvYheN96jdi0/VwlVtc95wKnWaJG4iFRmL0hB7/HJmpk8CVjd57DKoLDo3thPRL2NWxzCtHv
Wc1zO2CyktVtZTCz8ZAs9GFbz7i+D9XALij8FYPSCTxGq+Eysdyq8TfWUy8QQyG4sDYAMX+aYJuG
SirLtW9cpIEm9UiKvGU3GBQv9outEYbJ7GAsD6He+cUeYW9DDUkCyKo0y6L1tzRK6Go3pJnopb6/
uz49WdlSnUtrpkHE5A3yw2SNGs4x9LliQtl8AzIYY55dyf5FmenTNo6jCiVATYwd2CgNHZQAw2aq
v11qGCjRyK/mKxVBJyCamVUkb4B4TsHNDmpOnv5Lii8Nty9JtifiISIJ/xflT5/FHkSpH13O+zag
M/sg27JR0kmy6IriS1CHsYEChPpkNOqsGsO853Ps+U2A/nBmxeum7xYa8YhdS805SrRiy7h0V1eH
inPk+UgvomouhBipXiRAJn4qahLX1BBv2pJNWDuGoD4+bOm4oKUKW+Rc9fZVhgZWelSFQSVI8R8x
NVVovDVfy7NJiMAZS3woSbuTc5puhzOxlvUCFmj73t60FYT1oHXAgh1cm6vwbcVgYOR6eEghGwPe
VqzfqWeyz2FaeQ/TJdH/ErWWqD3pv9FV2rsv1oUDxZHAssg6hP1BemeygjUBHOA99OC2VS0Rxtpe
YHVBdrdFDhcyO1Xwj7Valq6XoPGMZgZ2PHLf1qOaltB60hOzN0s6Yx8HbdJXGiyh0Zz7RWAoMgVS
XTnCDH2XmvXRqr9dz3oHXLVo/D7moXGC1FUO3IldYBj4h+tFpI5kRICjxpQyoQQBqHGcCsifCr6u
e59lkL8W3ka2jqE2VxwuJSTJ16ahDX5DlojjhhBwnfw67I8e6805+ZRX5HI3Evpik5b32y61vhYR
f4qsiOFQZdPK77HJAEzUUYMYgCK4/PR+ltHesx0WGC2YpxTphA0yyJmcHIYnERPsCmyd9Lg6sd0C
S+Z2NroZEEDPVaYSRXQcS1cgTzwDYgkJp5uh0xwLdK+SaaZUxTa0LNAl9ld+ziab4wSczAc4Y7NN
+zNLR4YwRHJRn123lPiqcdV65mzE+4hJr9dJzoJutns86RmEWiuSnDovrFg25anBSRvujfriaunJ
Nmv5YHN9ZNhnG6McLDYQJW5gvVi1cMeRsh5FNSINXjaijUlOZcPaipgx2PhEKKvyjSu6kQbF2NYO
mPoaFYeuI6xs9cp8/Y3BFt58zQGJs+3JskXg87V+Ym+8QmE4UmL7+XZAurXD+z73275KGXcphlBi
cGmTwfHecQDY8REhk6AohgXlhB4ytfCbYbgbNJe5lbCLiCpiYR21UicAVe/RvC867Yzm88dGc/CE
fePMzf5+NFlzLgTXgna7RwMAiri5ZQ+ZIh4NTpyUOVJcWi0QatWtiXsC2BigjNkTO3PIgAbDkgrY
3eyeQTOFr3V0snkgotGWkWB2Bf/YGv90nYMJMEpD3N3XAMAcZkiP4kLCOSf+RMQTtanRhp7SJp+E
mNBV6jobzp5zDCcef2rmPMk4CmyFosdDXuTyZS71RDSHhIzdX3lRVtvXzEi1NF85ZGLfi7PjNKQ4
1kzqIuy/AUOqkV3lh2o90JGZKi494Y86HMAF/QPmFUQJ4btNvKSAfoEPHmYZi84PJaIBfXXnYDI/
Pq01cjJVBd5QnAkGRec8CGkEoQRgDnfFWKCI8rLJaglaA/RL4mRiR/rXVqWVPXOXW2BAxa1CYjqr
sw7rRMVflHSoNokDPqjxeCWBt0HUl4aOaXVrge2IWlJE94VFcqfjC9k3u7a2iqMzieLPa4kY5P3m
iDsyWRBVxrPPXvKCOpQqdIB6S/IoOzb+G615xW2eRserQD4alheFZ+ocqfjeacrAIVylNMhG/Arj
YsUqGrzFaxp28yjVWQwb4uXUJWVZRy/feg0kR/kLrW2lryCoP7BTIKGAsiBRXN027hcuA1ob9yw3
k5L+dFk9OPHj+mCNOscwYHoWNB2f5yjEv/+EZjZzq1qmu5Y709p3zLVsnafQ3lzGjd4wDvqRjnok
BqfHbqciR1wb0N8gMObExKvJWmIiuuAZv2plzTGbipRe67Dc65wKiAw33fpugGKp0kpPDcduC3cD
kHHkx50/gmsZyXC89eREYrWOucHbs2Yf7SLpwJde3jOebVGOmb708A47p7CrQxHgth1DpMQm7sB6
6EEbTkyAmDdaWCXi0WLXUmq18UjKsVLSBywy2gpbaDU2PH3QFj2gMvODkFwT04B5xrvNz0GQADAp
LpbBys4vjtCWXYWP3LTiazaQJF6P9N+z1w/uQAJLqePw06WMX0yTyeN1/8IuFgnrsfXolGUZPsOw
TGi36WReJ4wB24HzHkK7DGDng9RmFg3OQI2fgOI2hPsxWkJzSOEp2yyNeQ4fai+M7Qq4OMBpjaDO
xBier8CtpbA1rThw2QRT7MysXiVi2h2L1wVLISi6J8Gd/hXlA5BwmiYx4ImFJ8bDgMhlGZnZfYrz
Bh4TpgK4LyUt1HRChAJ/5PT/a5uFXiqVoMrzbDZzESFltImTM+3NyzJAy1nJO9MRs2lYs3eD9wng
+6ZiaQYWjEiyI+I2kCvDjbW9pdqY97w4r0TAmELStIQeorIHO+trrSybzO2jpcrrLKaIjuIYdiRT
en5MUBjYDuIAU3o/p8rNjXQofmF1QIz4Saj1NEySr6aFxTdZwLAmq68LaluzxSfYmeHv5+HE+mA6
DWN+at1Vj1us+6+Z94myofWrrBQ3Z2ChDHC4RHbn2Z/5kDQPJ+MXpdv9/BIzi9QhcoWT4+xK9e2k
F1KS/g5iWsj8a+wRrg+OPLrSsJIVgIk384pEQypVpl5OE4V/Sz0RVAbtatNO6Q2TBpixk0EqaaoH
Vm1R0BHjtRPRRgKweg1Bf47hWHC9E57k1FufAo+BDcjbR5khThRwW7/WGNYdiwan4je0m7AbT7/d
bEJahgz5YzbGSMRcqITLUHo1crNmFNeCsQFyEcNgn9NJrrjLPSpPcTvfmv5d1NM+uc8GqQ7ilPLa
g4hdi0IEFPbDz4MlE9n8nFO+iJLu6pTc68Lhld2nNS+wCO6Msr6tUfsXIzuSJub5J6lZzNnYDu7j
tWB0KqgPyKPmgiir4acqmvaJNe56/hQoYqUGlPmIpKgTiGrUFMDo9w84TgAxyK8AOqhbuC2icFNT
QGeMtv3zeD1JOHz/h3jG9pGowfJ1226Ty7jstiVge0hGemshSSKZsK1EhO1rrjd5G/0UoyYAwvJ/
mT0vARXVdgWxXtr/ZDeL++/zqG6ISbpSoTBPI/837p/234gtNwYxcgpWZEpRffx64GSljsVRpu9X
0wxIBKe0KoG+B2+jSDfmTstQzylIhP0R7+q/BfrtYOhXPk7rllhMhzzECs9VL6vk9FHqm1j0o8AJ
of2Jog448KmYcCQpyuuqJVyA9hWXwdJGvwrmBmxCkjRUfjcHuN2pAI2/KT27EnwAkQQaM0s8CmYz
cS1loYwXa4n2XvNR1tw/DquWPv9fRCzvUs+XBLjfjprb1eHn5tXo+RsQx5Z/pZIvNI7ukcYcuaAU
734ywTvVt4850fTqyENfpfoGPlQaXdq5lmvtHxIhEVreIPVK+6Yz2SPmRQeadvX6WSkI6wRmloYQ
Tb537pfPqiP179f6Ke6MH+0nIWERRfi0hsjTWSsIuzl5SJwPR3jCqFGtNAqvCmm6hGEQ/R5edYmN
jZSWAyKgavEAXhG+y4qJNFfTFyTx60DYm+EAILC7TeIoI9iL+MkxcH5cXXRg6aCf2ulI5vtLvoq8
ll/ZXWOSXS2xzX+OfHLoHpaLVQ2ILtXhMsw/YMUVAbjEcEbigBisXfVRXiqIwjFqgrxYRiy6Pl9Q
R4oP/C8H9Yq8NyOMN9LDEVgJGYbOq7w/vzDZJGRcjTz/DPDdH83P2Boy3BJZNErrsIM5MF8cd7EC
Lj1zUQQN+Qt0wD6ULQaiChSRKgkhfXkQaHelk6gZLro/gBFONPJ2vcfgqrjTeBPO05JwGR0aKm7m
dNwyuTPmlnNowt4eCX52f8mdEBT8T84Rm6kVpHO4JntpIRFIGUDJUpy1n/KXTDIux8SuHzfdRjXi
rfX5ZyYbrQQjzhsl6AOcaW3ExCBfmegmhNVXq7TFsdNew5Ins5w/z22KcCYxkbYP6al6XptjowKA
WGIZ85HAw+2G4sJMEkZgSNjaXEbbfYlQFO54uqLW8up9uMD0XCOuWL99Cpqhvd0sQTKF+5K0I71S
OJLvpFjUT1MXXLRA61rHNnhUcNLRafCGc5lTEP4RSrBGsUXPOUkvu1ZLtyRDznkmWC+gP341PV4d
dcx5AfFtrfQB5TCAER4WQ2tQbfZhcLfLWaBHc6oskbfoBdnvrvOFazXlSSV42A8QCaM/u5w8S7kw
TaNHvoaKH5M5c0o881uDWnJ2gJgZL/rOjuikZSMftm4ULQAO8uAkgS0rNfaHywoomEOW7DNpOjA5
eh4yVHCe95sIOY9xFteRxoL/2hgpbCd+B6Jh9JlkOEGlr2ItbHdKURm9CNyYOL0WW8iUbrDRNm9h
XvVSOxrAfd71jCTaA6y/AU+IzWymiaSdcxIMLdrOysapNx28LOs5JfQ6hBUb22zeguo7SYCZ3ske
MntV1XR4kJjIdbEUzeZ3m+RTM7CKT/RFR0ElsvKv2WUTbiOn8cBO9AOYzUlbMOXvxLpuZdVrFgSQ
wYPa/sWo4OvqqXHWq0MkmImx/Dy6W8dqwFmdQ0LGyofDf5i76nd87VocGqbMORQ675hrBZLmn4oP
NenDjghIz3np07oiLfT4Q+4/1xIE4CffLHNiYZup1fy2T+mozsV5XuNgo1CfpHeGVGDmFShCr/tZ
J7Qq11BIv8OraWOG2oI5rr5PvFQ8dESqf3EnMmz201eYEqgyDB8vxdMvPQ1Ag+j8cYOXt/wFR71D
HdVYPgCyyr5bYhtN6Lm+pJCNKvoQTUdGwcSzooMV2NywCPZqiCzBFlFd56glpWPJWTlAJc0RkPP/
wEmV8CeKTnhp3+JKquSiSz8Q7w44B8wp+Yy0MJccVRjDLu+YBV8XLIXeQrr7SP2Xju61ryyr9c06
gBU1zlbhTW0BXvTaFwLIanRLKeb2gsjI7njMt9qPazw8YgmDVxZHU7HywqJJLZBSkCQHfw5iu465
VAmJOe2oKeqXMKb2jl7nsA4F4rBvHWlaQWeZ25Fb+8WJ81WZcuM5jbNR0i7sdD2GvOsTjpv3lUl9
jq6BzaPIN+/38tc7mzUwfJrTsR3riGidjQq61jslnSAVa5yu34LCsAxREoEW4A5t9w1CkN0bOxBD
X2c549DgLfxr9GHj/efFXZLdMqL4glHhFy1XkgRtC5Z0MCulgr3OxsnwP2wibXJ3jpNGLPLG9Y8Y
mocawhqCKpQJf5Coeh/oHTAthsooth/ArJa8Ln2s25TOoDVekr+QXvtRKN4Y9ICUFb5qsrQaR7da
GTKz+d0Yvwh+MM+iRhaSN9rF60LFHn6qEDNfqc8vIsmni0M1e/YP6j/IafZbMfpc1IGXsHTs+475
dbYiFIU2IYyrr1Z4mdP9rl7ljexfk9yh3GrvdmRuPhpaZG9yx5qyhI8m3Ny2+1wBxw99MS6zzS7O
zLGkXtbiu0xKvjbhltTRyEJ9GsoGdvz5y5NivF+2+U4E0hjKdXr0vkF//4XuaMOARIcun2rclt97
C3hWuj/Qslt27LvykY4h1jwMxNJKDNA9RuqCRPpFnIZzjFoWOBFNWRd7wUecN9vxECM9/Pv6Pnr+
ZyTDkrUkOvFSSxq6jNF1FmCI4CxO6JIymmw6T70v3FcstiitfQh2Gdjjf68Imoq65dhoJBs7Cx+/
pfVizBWV0hsGU3DLjJTanvWYSDsDem6Gn8Mh2LyBt2dQabDLecsb3AlUmYVZ5VRWgqaROlqc2jU5
cqUOiF03p+by/34Z7A9tyvo83KexHkTsvN9L0g16rpRRD6Gd4vvWi+Vq9nbrA+YiwqqqHvCvc8PR
G42H+yQHlFO3MZj+gsbgvNZO1+obYH15yQ6pgdaktTsmi7qiQja9Gg0cUo6Xq4bjtDvB7/mvCwE6
hcLQ8DsQLi0dVMVEFvIIo80g8mkC7PiUECwbAYC8O/96Ag+GpwCoAdz7BGkgZURMp3f6vwcbYYdQ
AIvSsHJqHa7CrV8qdF4kWwixUN0s4MFsv8wNLV0ol21gjYNPLqth1OujXwKq7lS9bfG214r5kYMr
sh2YqgGrKhNFE34q4o2OZOJnzYVCQqou4AQhcKJJoQzemoEkInJ4kqTSSEEjEioqhS+rc3nUlrQg
LcYqnocwWQNkSncXnu+r0k5X27YQ2mSAdZ1k6ThMimAV4dC0qmEX+uyAFkpbv8GeWKunNNR3YfJB
CKaTvdrayIYw3BVSYJzUDt35fEQGh9P6mY8fz1X4QvADg/XcGvUFw6dL7uVYmoRLnwf727+mn0O9
SPBZsQbQnezI9dUi5G6BPLrU/JuoOQaRLgCbkpj+M0re/fbf0o3K3T/2Sf9Wz/mylN0HrBsHfoNQ
9ejgCPYiGmpcMjVD1pRmRc8HQ1Hwy0AnRCDQYt1gebURCfArkw3IvYQOV/vSDuttyqwN2BXzPmUY
ymzUyhgba6zYIVXYjxKQ9MU3/WoESvn+9U5y12I/mhUZ45Lti4ecHSWd7k4MSrUuJsieWgOLY4Id
RmY5QmWo+j3Fkm7fw0KyAWGqZPf11DKpASqqM4OILM74YjoJJtls2x4h5iUboczyRq0u74kciCBE
4lhZRoxQu01scctaWjglFTLDEhwJ5M/YfIQWVflN5rDIZdU1MSnvihrwe73teFz+HfHJOsrUYanU
kCzGhntmlyD6uT7C0ItvBF5YUQCWlehBk/VyIy5I3QAaWMuUdZzQHBICHTLUIkUQgL60sodyGKpV
U3grDD145cF0a5b43MB4xiNtKPuJOthcLTyQEPz33Lkjc3yDvG/7RxCnO8MdijBpA0/yT9eKRcVt
sgAv5eaOXBxwJxODwDws/DX2oUCMyaCvNf3IqQjapo1WvEIorSZ/Mq1H60KmUudRj7RTiZ0RqLnS
EmJfPk/NH9I77yrV11u/29GkpXVDzW5kKEHBnePsBthE/ziWUfzfW3gkN7Rsu+caC5PE2AfnnGHd
09f7IzBTT82BDro/p9T9VR8YeFYB/eLs3Q1dORYSeT5pktVrG6hQbLGlQSzOFmX4VLms42js/8nj
8GulGqJZjoxtuN8cRckmoAi4bQLtITopERjk1u+x3akQziGBPtE/rtju8qyypeYvKvRl2u0b2vR8
LM5Q0VdaSRcXv9H2hhkHtAdtR+l9CrrUIA8rdcDIonFB5TV/TbqcxtVJuVt+taHsPbTHAYvLCqGM
K6IESvM7uFuvHF0L4nnU+DJeiP3Fu1LqXzU0nGDFoWGUN0Fyx2xHoq8c1l7QnZeEwUh7mHPYK9HG
8SfT35L/ePI+8OlDbrnB0hBQE1WYa8/hLZxBEziv94pnGsWUTLhB+RJX/XtljWpHzx/QsV6SH7Vn
jID2MVjBWMI1Cn9UJrpxl07wLRWe5MV2t0tbkNthYUv+//VAYI7MdifWp4YQaqO5Z4hnMnfbcxn0
d2aC8xXLxL4PW3hs9ACIuh+9lTfnwQ2BJYJoYeGaRGipFzPZh5id/5nsC5vcfj9ihgxCZ0KKtNwq
mff1ozyCUKL1GJy+Xk9IsZruAHfBWXwMjTgjSnYoZJP8AS0nnkR5h4URqG6uvmEP2mVBJ2vFsmxq
2gMUenHrBxalMRcXAsGBkYf/4jEG5KPZgk2pOP/OCD3I9hwqmJydosmYjYRGxZApzVQle3DWuO9e
hkWfVWAldTGDaNlkxk+1q0M6HHtR2RGQ6JlZ2NzE3c0KxiJB60/7FADy2ddFNqnYe7sZX+hfufPm
b3P02z011TcSEF0+fZ0lFD5vmzU1k0JoWwjNr2eoZZuO5rO8B4LYX8NekqAVgp2aniOLbNv6sMK5
3x2uE4ombJPpWJ/6QjTZ5ywuF4Y/vYlbpnKNhc8jbYCzlfKpoZaPWST/x0Juv2Tk2RMeXUt4hOQB
WzA5YRd4vGeF46RFl7wrhZqGtEaBf3twQfMaJmMa9JGqt098Sre5pjUgJ/bRbBdlc/SGWJKwX8RF
DnFsg5s3eOKQ5vbSZJy66paimeQAa/30bvP6m2q56KzFHp9ryvsZ15SQ+OK7+b+/ToP6kSGQBZWX
v4CuyDKo5shq+FgZ1md70L3lyI4e4fD/7pbIL28cr1w/N9d5zKDHKhaA/i7hGzbrHNEIU/51tQlj
RFO7i6fmOq+QFQRY865imNk97aCoWU0zb9yzlee9yVNGriklV76cQPAj8vv0BqrHe5dXXl92c9vb
HqfJkM/vces0FZ8+igIcvc6OKOIq7Glv1RRxd+SQmlnM2ZQgGtvj8iedm0pHTtSE13xkUrFSoYGN
qjztPV8BgFqbLY/Ra/ZGJc7BbaFsZ2KtYau8dWNNLDNHrIFk/QWnNhi66n5jNnP3bZX9D/4Uun3d
pDjSYQogdH8FCMDLh2xbtqOkG8s6glZP6yxSSaD4PenxqcmVjJHoEsrzaV7WBBY97Hwd7uSWGjIj
2kKugcRtIc3+uoid/LLFEnTrSCQWN/ywwka6YFbL0hrv+NEE69GjALrM4Tq0JdY2pv2eP1XLB6Z/
7ZpQ8oP3y5nuzMtZuSeR3B4SPsMVLSzhCcdfOfRQc8yWx3GbXadeE0oEcmpshVdsFqaWR0TolCDv
2j+m3f8GHQ5jsbLVFOH0gG6ht/xpRnlHceZ0VeT8ViCjyrRviuLZjPLyTOcbww5kAu63LP/ZbfMk
G8GADVbjdcU7414NTfgOHAGbUhKcUR00KIG+GoU50AMsRIv8aJNcuEVrma2fixzoUfAvkOtcu45B
A/LT9EcXj/Q9JMycPXmvk7pX7lD468yWznY1wZFou6OAtSnPtpfrH08S7Gv28npUYiGRyFTyWAHb
3WnXama+DLaqvMT01iHD3mnfgGeabYgpwFFCvVaZsXIjmrh7CyTVmIRimcqOOwnid4oGSjDwiwPQ
/Cx8Aex3tiXctl6ppziI2EbrcIr5CxbD3mmko9OAM/Psjk+O21httcDm/ks8H7TAXCHqfg5NEsTx
owXPKxejPF5pWCrWkrH2UbLkgn9+TUr0To4Qm6Up0nq3tp5NjRyaVo3l5cf6OtpJ6eLVWPiDfJlK
ipBxQuxx0nzxjHRZ2UA5aXlVWcGwimOvHeJXKm2JD3ZDLE6VNC3146qF4FqhvNgXiAdUnPKSRA0d
6lcmvUCxcyNlo6+tSdw9bUFrPASSHu7SMZhZoxizZO8u7C/5RhSnWzgJQEIRN/pJgXjdE9F2MOsq
PXJ36yWSdA0Wbdx3BPJ1yJYPUnPRVtBjVJ0s3013+BZt53z/BuZtmbd559v+LVMEg3uPGJCh4SLl
PsLrpXeRAwYWpw9P59w0/fKozpjejVmbcFfD4vUnzBFmKggJD0g5FGDiqCxg5rGBd0ML0wSy1e90
S/VVSDNcXB99973e9ZzUqRmUAUSeQT21W3CpKJMLVIO+rw4uOGlMXn0WWrA/LxncPXPIXKND2FvW
QBN8hks06gOT9N4kep1N+ODSD5GBu7kg2HXfmsN4eCKu44gYF2aIrsegl5LnwbHMJ1vHncaTOmuR
RK2xHVpYq2TMWPL/Rs9dv2dzJS/G8xIf5682rFolgbJ1jgsVZfVLFdC0W/iHptabl4L23ILww1Q3
TM24pmWmHLtIknEiO4QOMaLBhZdH7UxmUhzWP7bsFWQmMibZ1Fc4b7FcuUzqiM1B/bPnTrelSJ8D
1llnBq/LmBG3ljazftogkt0b3nyQzppk/vIxGIOVTR+KFRjzE1gT3oQnNJ/Auqkr7mSwz8+akU3l
S5mnT9wT91qXCcZgP1fS3CN9cvCMMDBZ+mNGbYHiSgrWa25ad6/bE7ihniEqtQkn2V6Rbwc5JeX0
IoAXMyfFV58D3f/jlT2TUpZitzZljXA1TDFCERC6X8FOLQRoS5x9Icpt5CgYmc6M7EsTTo9fhIbo
LMVH4ZOAUazdhtojxWPDFH2TosqY8WabdWwQU0lp1xR7aWOzDhT2YmDsv2Srbjdo7K5oPjW51BsV
ZAlPxTTMyW4LVxytm1743zNs6t1uFtB5t51jvhWdK8+SxHCP79CS2Go1P6xWMffPATfCChIfAjQ0
LfAWsPpQby8GkquNNV9cJNVUgkyGcrzn5kI8fyDi3WBnaIxDS+kXy2XKeKkFGcciL8w6JjPvCFXy
t6hjbKvplVX7fyUToTtotSY5oDfiR1hAkA+4S4H6/7Cso5hxf6THhMQfGmSnqbPKvJKNPmMarlZT
RsF9w+yhUYGVI2Jemthx0qci4gzP82vHDynN19rPfVM0FMWJ31PuHQL86jp+U+qXittZCa7vNrKd
/jzZnWAcE3tRw+fV1S1FQxMo+4swtXAp8h8+8IAQNFMJU+eVEV6cwQ0idx9j37YpmnA7Uaa4uQSn
Pu2sqpY71sit07SKOqYfM1e9A3dvxKOsHyJTYSti48tZcJr2y9uxyRl4qg3e/osQslcpoBPjfWlB
J3SupiPmxUVClt/Ljx6o9r8KmsMlzVXfb55SRGluiPd+m9jGk93GojW654gXYtyjDOw7Ue4KVkhl
nXppXYbaTyFS3l/mTn2D/bhlZmel0cT8dI62l7oG8dKEtnu/tAr3DOZymg14E16JfzXw6cQVkO+p
0hol2DFY5OrNRTGvSrXSRRLWCffXbKF0ODOWUUAxAM0aQ3T1dJvoYYtumadPMctg16rfY+ll5Sqk
lF7YyK9lb2VAyzeyexBmHAyGkFbXrOJzQAtbecjltywjEAbMzJakjQ7UvfezVNi2aSCuSAlojJ5c
HCYK/jiiIx7/zk5MCHP4PUZslV0c0EBE3BOS7r1lWOu9QD4rAcQ7QDZrn7au7mvxquBu9g2RrSEB
pwnB3oXVqU23mZHzW7kKSms+wteax3bUNAUCBuY8ZHWEdGwe0ap5uc0QrbTR2SyISp3XYiPo8Ilc
9p/RaFShO9H1BM0MYoelRiSGZQFxqyv92XZvgLAKuDkwnqqcufyA1Yu7PwpFWXNbfo6FHbyV8DtE
We3FLc65q8Q7YSuuoQ4DnKGdyUWyQQqnbvZQB/16dde6cSF8b89Lm0i1YDy4HJzAQQB+ahqIjW1S
OmabmGppU7OgsvTXOsaLS0cf8BwruTPq3jqV58vx3I4I6+B9EAyhFHT3an3Dyx8MVZ8Y6WLA+lD6
TBiuJBfObECVgeUJC87Utc0sazHuP8OvGMj9+GgTACpSxOlW4sZGNukLsvDVJOtPhY6xxaLgeJ5V
LNdgDmEQwNvvFCMZ9H7QxFl3SDaaYX1iDyDFqPGRww0+gdMsHJAAuq+f7X3WA0FNoMqceSCj2KAO
S0AyTbLRcHxutAIsQDFA5W7v3r571GbEOwnwYPB1qF8xAKOW7QQ1+If7ZLMA56Z5zbS/EysDhk8N
GzcMNeLMK1VDHraIjopQiiKWnvlSUaJS0pWOYGZxnpyz7FUtWIx1CgLSh/XeuICIjfcTLMG4X8jN
J0pf5wlaBqxxTjWGa41lq1K4XyPGoUk9BSyhBadksPvPUwic9eqEv2fAyg9RY0Gu5ZL6J8FLpe9p
/HV6vnQ0BKQd5v0jwE6c1g11/1BIrAkjXBoYERO4UA8NqBeAMxM93fU7urMggAS21AG8EM4+edW2
pRt1rKSPn5+3I3aPC0yVCqnyUMFQ1brrWAtnA6bnYAgeIjs+pxa4p3YOxvnfMN1god1kWURvwefW
2cXrzKAKRiVdiWAE65VIw2lS4DqqhCtYrP9U9mBBA3j4RiL2ic9J6pKKSocI8j4GbNK7EkI17pYK
hV28TFn3+6NyMgRWdv42zzSiFymW0K2u5Iys44vTHLOEZgy5Os1yPIoc8VYJhmtOtXLDG5yfG7dr
qGuCpepXJ5ejIB4NrEP4iWpCaxi/vaxMKi4ZFnx04ezlRaEll2dwxcsikBQr+aWS96cSB/rftCdh
Xcej1m4DYsDUO41BtGv3v932wuZ6CdenZkE2nwMO94+AR3nBl+1V1exVoEQGqYa3e8ycBWmvOmcN
UBbH20Y1GgsB6VhlAbQ0D9Qkag2gkRfF3/ZmYSiF4Nw2Taco5qfbip+nwZfOYw6Az2HFczXPMqOe
UiaRm1xhzrHMNqYtGmsrmHb6i+vII8SnCFU5Kyk9BL/k//lOESJbL000XFhw0PeLOlPxYuvD4mpE
di8hIqRcfL4MD75+v8rthGqrkNRGohGZAWRHBE1rq2AOz1+NQ3MKOVPmpFkdx30PSFwH1uazHuof
vv1emb6CNVZoetKEcj6WX6q7lUCMiK9mrIF4GceXUErOZZqL5iHvtECQgyhSK5y32N74GUI9CO5H
ZMqFSFw4maNhMbqPo9C5LPuEZS873PGtBkdT6tAoAq/npDJmmFIVbCvuBDgSqKBqLOOh5uwHBfHN
gWx352mpXQpMJnu9iAzfhlBA9fdHnQQ3kkzElXHlADIsbVZ+B1qH8BTPGZ91rX1FXasFzeCu+9+7
dFtNm3w+yALcXgSoRXt2VGxDJI63itzEoRGfolpxBEApsVfdDsBxOk1KqytYcDgACE+19FTdAfd4
wWRB5YRlHeM1tZgPPux9m3CXWJPsxQCdfhLJfp8h9TzwP/YqVdRVQikGmGniQMqOyPwr3cCmiFPD
1uQlm20juni5Dtppqbi7B8AmzXpb3VtKAZTD+oNvJL3rAOViiJp071CKlQn/3MEfwTdLrMusY5FW
HdiqHX/M/YRQB2ZrtbLaLDuD0yZktSPEE8pp33c/T76053R5HumU/fCtzkRwAc7WPzAEw5DZONVH
ejPnxyt7X9nDOTSs4Fv/IYKIxyeGSJgnnNnPzu21v/nyqi8ekzxF1riZymOqEtwwUGdiUmiiDErQ
g8Bcrxrp/jBSceZEZNKMaGlP3swSNRv1WtcwsE3riQhOB62tUBh6x0WxyPgDvy7QsCurB7in7HWT
jK2qah3+sp5sdXkaomdaHgM2h6CCLUJYwe/J/yLWeCUEpgjtglV/FqdzAha+Gwk+89WWki/HiYrn
OEs6eaeIY4o5J3u4ml6w5ue28iGGXBsceXYnAWFTAxLYskehNsj4W49nVhnyKPYc0D2mQO2VEq11
U9ynyQyaufeA4l1vwWqcPqIIkzLEW8KrYXvUDx2xnv8IJxf/y4GFmdQ6B9b3dc6atsxvImD9NP0g
yzq+FeQ0S4xlQHVCjVL10c/vSWJjdoFgCYvyXSj9bf5mCm8wEozTVKlUiP/0FMszPVk13B9lajob
peQ8FASJXGd5nJ8/3TIBcor6ZAdCxOn61EgjLtbzg/m3vzP2RepYRni9ZyhgQWumvQXHSfvI1cfG
l8hS2wykp3JzB6iA2Mln6/1Ic46B60lFhVujYeWhdmLLoMT0NGt2unCzrvaYApFyV1vZ+hQcPQW1
sZ9cqX2gEY1+9PV8Dx2rRw1KQUmBVcHmBlAbBmHxqXFX52WkBSOwCC/pb2y3sxcgAtykeZKJcObV
kZFVoBRkvCIWCIpu0vxK0ZzMZLN72ypaA7DTvyakyXyAaFx8FDvoMAwYNChPLcHbBYORbbOSDmOO
asbJoq6d7TwYpoNQCeurYvYXxtEWHBuXKlD0crelT/s0wGQBjpdPSELpW+fucj0xCcALBxSxhTsc
2y2EVPFdch87LuxULrFNfVBNdnwQYvYFECJ5srAvHf817/TF+JnUKoYfb023cQjFNFryoUvRqJfl
+AKxBMBPMOGSmY9ek4n093GQsnrnqAcM72VCQp+qlM2A2vIq4+SWTK7lBW7wkvQ2HZ4ETb00RR8B
Pfs4Gaq/qqYFNLX+mbLUT+g3YVzt7wE1EreH3swpF5XnvyrtuThu87qmrhoN/j+2eoHkk7Z9w0YL
rklEXaYWNn5oCglDFN5xlUgn9axzkmMO/OMlXgrUId3w5ruQQeBV96lC1P3VYYcZrn2HTvtp8FIT
F989YMV5M3dXBNSUwn/0AvDgoB9oZCD5+W8Ww/Jny0vzYlG6ENWR+T5eXeNO5ZXvBW1YUP2tI8kM
F5ogTi4bSRd0RYz85HLXPTL0K4NFe8ghpQ0Zdh9DbQG7lmokk4esbME6Qdu4mdcP/tYAf32O3+el
oEzOLchlITcd9Zs9fSjzzomVSoMWAS2jIhn12jWdl5Gv+bCCoIFoXeXqNIPENI7bNn9H7PvRBukY
6fxtffFK3Pg77rxqik684ei3czYdTEfj1bhNZ3+eOIVEHSWaNpkjtAmZgLdeZxonAhHbwbNg+6EW
Xt6f97xzscQjDEufQmqLqjeUFPrRP6WnQj3n8+hNMHqC9nKKVRVCQGzRw7B3KKmM0P35Gy7NvqoJ
j6sMgW/6Cb1i5a71AjgK2t9Tx1giUWz8MbhqM/fyZt0fFfZTWAQwebowh4+NpawiJ8jZGqpbV+47
jUDcr7acmPPTSWVTmWgJsFdRoCpWcepIxBwInwGHv66d4WcVqEHgQosPofxETKYhKt+uzcnPDZqd
qMOKpvpdoIYwQhABu5I5XpkGmF5DO3RMb8M48kuDtayYRkKmf7kjEJbNpJGtq2Pr5gHx4TtXZr6z
sagN+Oc4mcIlMvlKT18BtcRxRNhCYzmcQZ4x0zH9//WxXRu97LOryOo2Dmg984RCenn43+heYk0H
b0uLOtiJ5EIKl34w18OPh+AaxakAQOROX7zfMaZ96hx0nrViH6kDBXasFFfWvf9WUvygQ5CHGBOV
hoCl0BpmfyVpX2JCYLQ7qfZbaxBKIXmRe1pfwPXC8srFjN6mYnqDsYFQ96clGNVSZDYM1QOOYsXW
iUfYa3MqNvrLHXADOhzjXrFCo1rHXIpRO9Zav0uMyPWSKQv+gL30DwwK0qjNgKULOk4ArSl0uci7
OP+/AbXK4nRoiQMcC1FWErPCeV1YzyhaWo4KVAXs3IJeWCwlC0n4nF9KuSa598wSG28eMffN3xsD
5Ti2FcZX6oLBRIcgw9fRGezeD02/CueVSPytZJwpgOdbLek8v9cU8lnkZmL0wIwjdchnux3pk+lN
K0EIi1CnnIgrc3nZcwCEuLkNvzei+mckrEnyGk8MJ0iJa8ZGN5L2gjBsUjzs+9H78yHtLduETCEz
YKtEHgo3RFCsaqiqF3LlyJwN60PbnojqZ6ZqQiSoBFF6PdnAOAKqPdmrJwqyFuCYTfT9GmO7uyCc
1JzEysstVjWAvCClPBeWMrsJV2UbRm4HGZtgqXwPe6pHe7YxD451A5PB7/T3zOldhHxVzTEAmwcd
Da18/hRixy1JyZuzP0byox16znZm25dKCKYFwjeu+H3hpPpv6wlSAsE+fCTpQxH4JYEmKbzz/toz
1OEB3EQNDuP0h+Wq/4zZpbfJAXX8wxNCoxg1//F+wXssFlvMjcnIsRD5uWyemOtmz68gIivtaEAI
vORp371hh4RS44N7Yis/+GQueFZVxJCsZmTdrTucDFiDNh/bT8ozvsr4WnBDHEX0ma/TSmNHUPxv
bi4q77DF2TTMOEH9KisSuaAbZmzOcjLdz0Tbuy1RuDpJIq+RHN9nhbU12namNM6iN3uA4a9OAZxf
it6xRCcHOhsY3do1dkhhUju8m4UCW4t9BnClsb2GRB6a3IRh3Tj1cfLpQF68PHmkeqHI+wal149F
giTlJgEVCYfxGFuhEh4fJuc33yKfLavuISCFMNu/UqfZlxM/zmZwa6GEMcdRyMCgCDF6yx+1xX1P
KX28Fzu4UGEwzN8pptB2hLWVnteoHOFoqVaMb7CRbAUFrUobGuv0oilES7JYuA2AS2milBgovqdo
HjwXJgdyI3GFiERDPbhd5peB3lXN+06ypZTx4IIpcxt00A3lokcFpnusW9pmG0rP1cnmuv1cidIM
osdXqh6Cwx124NM7wiVQteGN0dwNyjVibuwoANachy98bGi6x+lyqJphtOPn3PTr+wQfeXjm4e0v
qlyy62P0/nKxapLw/cUJ77R3cENHnoxIMS54qf73j05wYKAu3kLOrVPiSd/+6V5Q6Z+k73xRkrIO
0UAkrNld7JfP8z/IC5m88vEPGsz42aNNiISSbNgyjV1MtfcVSp1KinKEIclY2TrXbTZEIMQVqoUO
d+/10gyo77491Lr0lNg0XfGLf2OF68D4nQ8fYvfq6UajD6142RjvgDz0jw95QsgB28MbWZGlqvtt
dTMZzdJrjXbrpvAfgrkzFvuXMR9qSqqwM/WITFX+9ZyOh76g6Dx6BNuE2z5SIdPmldq6dlEFqW40
GXEpqdjquMIA5ytiWt78MY2JPLyiR5M45rTYW8gF7iVDhqH3RUrME6ho0vCSrliv5VYByUBv4YP7
llkpUVytiRMNr7/wA4GQgjnM/BeWfAux+uEvxBfSklr/EbDZjtm7QH+mZj8xJlJQDAMPVc9PhOC1
j5zMa7aiT9+28BeHkQHeNnJ7iJZvmrgP3AENlUGylxxamhHWaz9txg91hTSENvVeo05Ez5BeSbLW
sRTFXj2s/BBz8LYCG+Nky+Rj3L2S86aM3FFeuAuQ85mX/ogxaF3qzKFFOmOIYo1Iu7CIrSsDB/Rr
JIujLNmVkRgMVEEqW+hRlEFnTIckcdXoxKJAnm98oYSowSwOUc8mRsb/a/zWmRT/DomHW6P4iXw5
IHyn+IEgyJfVkCjvG2p31zwDi4yVgmJpfMJ3XS+L+IkpC8tELeeDnhQiRBg42vQk/osVDU+oVE8U
+Yp8I668d3yKBieWqfl00QTfkYFKRDIPTc9alLPB2dcCpSf8F0Zb0+tmZfNDkvozRUDtNKIKLBkr
uEhttIHgW8bdt15Hls7TqW9FIOc680VATzAFOTe7uA8KripNLeD+FdjfePBcg1xijCIhGFWCv6NH
998UzD5XuyLDxrFy8owmT4woAyHyxFb8gOMwW4NWW5IdnY56RAFR0B6DDmHTJge2/HFl/A2iK8wR
Aw4mkOAg1URDZkY1MopAh1CMCu/wa1saLkGomBWjb68emE3cX87wqD6qKkRltBhm5N8zfhiwoZOR
oTPKVYnhcwcGv2nWq/ihK+ypLSfm9qNjfVHAKu1sAGsG3ETS7pNhR4fFgIY0nFzDMUUd1gE6iACh
duKrXQuUwPLdWBgKWyH5lbH6uqCjcciyZqz4WNxBMuIP7rVfBOb3XcuamK/3wcicWfZcrst29Uwb
Zf4j185A8HAF7x3S3Rxt5fsARIe4EDYXZoOzk+/NcHCe5RCzNf+kIS5E+WAVkdl1Du5q2ahmqpAm
zNbwtjvoHK9ylNdw3dTMh/Pt+WGOBxBLYP5RsePJSM6tBbGqqc+yiRKUt22ZeJ28Iu3ViN2SGdXQ
zGlubF2wAXv4RH+wgNqr6gL4y8V1p48IYe8l/J+eIimyPlbqtMKVRE/byCjZDMq/xXwDYkDsECS5
ftgb6lYI2Yr/zRiIkM+zy8iohxUiOeSCRzswLUo4XuIiV+ZLd1y3P1MOEyFvc/0KmxsrZB4CUTb2
z9MjsIc1wu5o0FQhYgK9zz5IlcXo8aukVjiDiv5cN1vIfcUXfhk+twHrF8iyvPEldjuuBWbWbHHk
flGQyCd0UrxiG7IBnnN7o83vtb9yKpnMm+QLcrjzOWw/Nd754O2IVLsoxWML9pO7G6PV5rTAeaWP
VTaRuNrDnYS+/MYcGcY03MPP+FuusqPio5Zx5JE6qXbUf5AsebwIFH0W9LFGAHe/FEhXXknI4tv1
k2+5sJvjKBfRds9RRpkzL9mLJLJRfBxXoaFQgGNdheo8oBw1wDdOgqXQJWZeroW4rZ1IGr89Oupr
q4kbeNO+EV40plG2wcT6QWOzxLtmpBpDAWrVdlnoILoVvCFp6aPSjRrAgRU51/Tib0oIKIaIQOo2
x0AyW5SADZnXZ3Jh0xP8i+32QjttKYdm0o7zl4hT9YuqORTmF4cqFpVj8KFxlGrb8ALO9zThKW53
Q6HMmsK1vHwy10AAKEz27hP8wYP2YtVZKKRmJgVwVCHspK/XI+47YS7Mkg16u9og9UwIjFgwuRRt
Faq4McGqn00hsyotBGiAjZth7jN5r9Bz42dWdDUTFJ/NDzmLs9XzOaWiPyssPvL4um4YDAPV4EpB
MUOXO8RIq53hNOOZ76BQlLBvWmdPOJMnSxcrdi+aOW5HJy4yr+e6LdRocPmDqYul380UKtiJmzgh
vbDLirWwGxMd+BD1KQvRfkv1n+91QXxILZR1QPZ36jBcevhjH7NlqFscOMfG/jqug7KVFKN8AQMa
DzCpJk3nwjs0GlVqLeWDFqqLuF9xGcQz8L6vXYt84wjlarLD2EgV2GiOkCxk836QOdnZf140KPkX
qNcYvXO6kHVib92s/dL38axT+uI48v4Vpu6533gFShYa17OyvsgbiLFkf5HtK2IioC1fdqHWFS86
cdvdt7+Bd+/Vsz7QmxOvZjGS4rnasQltuVRtI6WV10oowo7ZcPa27fpjih2X7WUm45+APrE7AEoB
qwDwMqXTcb1PjGc8mC1L0STGFnZuy9fTnUMVH5FhZbDsf2hIAyakvFAvxlLkAWu559Msq7O/0Jag
VXW6S0wQe5q//HrfOx0y95KlMaxnsduRszJMT+0LlCLtYLUkxATGECEUIm54tW4stNMbDAND1sFW
IPDCPgQJKAB/LSNf/SF8N1FWUB04LpvdDo6jroBHMN4BjmX5PE2NSISA+q+yWY/jTvD2swX5EPEm
N+B71RCc0hFfoKxswouTMbyd0eQinx/Lo3QCgmOuMcBIYzajSJSGJRQRymtOrC1w6KwA11mE+y4G
7XvtJzKx7gqXqDjwOlHoVWDZPBe6ViDDLyz5HRRlvIcuRbV13gNF4ST7koM0Al+Jn6IPjcLwU/fb
XzdClVkgu+XQbZhPxS+rqObPXR6dEAzO0KmAbsd5y1PyUuMhJ0mqVaqqqP0fNYSs8ErexBdP9lKb
+5EZw8GvZnq+m6UdLiGTDn5D67WTghN21lqUqCjtVvs5C3QCmltmSiu+FZODOzjQoQrb9jXMGAy4
35f0iE16sOUJIpvuJ0DQR1vpBtXk5Ay/DntEhvzSqignyAQssd9czg9zySQQeH8pjcqnc0IoiEy6
LgZhS1LnzYGScH9NHBQ8+xZuqfu+Z1rn8LCh+zA2K7qDw4/TlRYWo5vRQ3alIi0NebvcAV1/Oje4
UXQcxBkkvLmbjCaOxtDuG9Zd5X3bVHRSRtB7pF3zuPZSFIbNor95O/q9LG7oQsIq6lmGYmQTZk6f
rqUPFueAFrMMUQJMaE8Y0jEyA7HJuE5Wj+QtK5/r5fhYwX13mLEmaqApW8qc7zrpwya4DRhRd0Qz
HtgQW1QInF4eOmRVKc5yiBHcIKuMjWm0FJVmxVSWCmjhGAl/S/eF7WDWBhqSGIHcdCPP1yqK561s
CHuyKGmG2jYe/GEJTE+8Lj90UmvS9p6LkEYLiM/98iStMI8kIXGjl9peYmQPXjL8Se1q/A9dZZPx
tV4i9t1mKtpEU5FNb7MsIfa9MeolBs8J8N0Xy4mq+DanYkKC7E69dVvDHfl3W+nyHyXTcyywqksi
0AyrHo/67flPZIZOa85l10RBuZag6MXSAaEMpYrUoA1OpUG0ue9MODpX5kGgYOuR1W2j0rgImdn8
1jI8mTN0HGTqVUwA/2FKVtt64+bsFpL6Pu4doWcS/fyKtqpIM2o3kXWxExwZKFiUcPPkdZgI0ST/
1/HUNg9Ck9mIeeafx1KbYHG2pEjG+jXtSizJuHM1s5tV0aHgj9ZBZi9qa7WlV06M6Oak8bI5Uwdb
BLBcCX8IrRYrbBZ6dimR3JbqDTbokTCX4VbHaMeo8eAIce3I6XF+cZhmEapAqBOWT0GmixAyEJr+
NQpx/kkqYLf59inJfhrQFxEqr8Uk1wQ1GmiheDn6FUahRx8LAEMLg51oVPlegwPnk1tD7MhpDZ+e
AQo5gUQ2xY0I71wsDRera1WC8VYThEi7POczv6B8r37DMU+3tDiclh4RYISVO0xJlQ0SF7sjyyH0
m14yBR1aGpERcWGIpPuXhUYcjv91ZcXhODzIkkDcq6DQbGUOnWG6sBr4xdopByMoKDdyW227omT+
ady+QyeO26RWWZSv9QH1B9DVTcX3qDestf7DdVgg051UgzlQuljeic3JtxRNZE70YLAZpOlXN0ig
+QOQQxfX1kBwus7DXOZx1qLAdbB66r4TQghEuciInbqVk6m5cQydV7DgKzZ+n16XE1SF4EJe2yLO
gFoKMKttFVx7r/w+JYlM5hgzsdQF6SRCMzNxFtq3X0McQjNZUBF3ODP+nlNz6PlGgn7wDZb4//jt
29+kioWCcyQjO4xCl5udJRSkXdW9Eghd0X1bsJtcK3Wuokp18cf/CusQ30Fcnr0SbuwnoykYv8Ek
uTmZrRHZJzgv1szrNAZRLJ37TF6fwx+ZYPm7k0TrKigjBVx3TrcE+0xjujd7FhRqbpKp7PL7Kame
X3UrDjsyRN+6xB/GahS/0hiSfue4BKkEzcA16bs1jRcmaXJCL0TMb+9z2T1qpMatacoY1112lb5B
TLHU4Mm9dqSGHmWZ2EAJMVI3YjiBehRUAtXrMDi7ugRlRSiETzj8mXRLHiVUAOALSLJK28oVBKRG
/FgcNsa9KSPj4YEPKjO1RuCj4JJNKCZElGONSW/7aRKQDvewdzEuAqKs1EcFxXXJ9LOY8A8/Qqdd
f79+7kW4L592Ixix6ey2Yt8+2pJev0m0wqbq2XswkMnmyYr2fBUdLlJ6O5MrQyejKBZFCJ5rIGtP
3SjKBBp1ThB0h7t7ASmRiDYwukzgNHmw4PvLD3kWKtEreKLBygc3M5/WP2j6t/rSP3mSqpZ/UAmv
/il6N+eVVrsthL49M5d9Tc2Kaf4xAFPOjWJf9VzcojrRPU/BBD/HgY8Zv6CBofJ9AJxRCTKYvPPx
eC0mKVOCXYKyR/uXe7jJp6rLM1eZPSna3SoxnzQ5/Yl9bEJ/hKZ/2kSzLo6axEbaE2WSvBmjFYQf
czHLChGIEebJGVQoiMr1Jl43IOojeEqU0yf6lIrZbxZTiZUNUBKQZVezpH+Om54M5PNJulJka30r
nvEFoyTNkkfS0aF7dTJOLBncm4AY5eKo+lpUCuS+TPeclGZSLQ0APx6tSE/ypgPyzfMP/ay6PYFx
nzYoFm5JEVpj49ZVvlFa0b8F9sTfI1UKUjgwALFuPbJ2LnkiNzMlIpc+Nbzr3CRGoKDHwlgwGLuX
QO4am6K56jDgRFKXQyq6Aq2e5PSr8VaxIHGIrN/XJuQMhcjfvK0CLepr/srsspHAdAPMc6TOjXLY
73vSi43TDSXZiVwVBzmaPBpYCRu0sMu71OSNAqdB3rXBCOEvCZW3Uih0Z/BekgujS4SvTDfaVCvG
QnXm0X8EPlDlOSZKw5yfWwdd/DGhxIpMvymn9mVS+0bNDjhyOl6UJt86JD+/jhsOvw62jYd1GYSN
nUasxphzZKGI6640sMzLenNJt+L6Mztod8hfO/omdGRM2iemIY8JUXn3kclRoqAnCSre16gtte1u
v7W0a1sacFTv73ZRp5o+8wciiykJE5jA9IBlvcn+TOTc3SJuTNA93VhNViTRbnc/j00vO2o18nNJ
Fqf54EdoppiZzuWCfVJFaC7t7Adue9zS6kRhgEXglAsen8/1sS/NlC9um3X88XIUeFHRLvf47FY8
yjS+n5rShJmZoyr4MU6LpMhhczDVNMQhaT5sfjoY5wmTzveqCkR4lnYb8tT62NvTzY/UP/adILwn
fP9WI86vdrHAfgO28wjNg214LaYCS8Qvwky5z/6jWs2jh2KINoSBuhU32FN6gwOqWhdGT838l1oz
owfCA/fcoVFfdoMAsHmcWLxSZeCcWHwEqP/MZpZ67aiJcs3C8tv0nTMCEnLN2ZkUQ/2KYygbqnuq
X763CFO18smjSZZBWamv/clkZkUU8HBspKWUEWkjeL0PCGCJKf/m+k1kcVCquIQ3t5ehxBMhhGkB
5nfuw9OSh4Qed+2WndTGmqDJSWyQ79TmziM3xh18XJ3FD2ZOSGg5oEnO/rWDCHSpUbPDVx4Fvws1
BfYejKe/3LjE3hs9CLe9uuGmcLKalO+5q4HoG02M4TJwZ3kCZtHVKnCVrG/m//08x94AiWEjeGOa
oQoQeMLoh223HTT06uXFro1PoGRrbPolpkFFzDNtLLKkgFer29lNY1YhnIgbKliHK94EFUImsqVJ
Jmz53ggTH5O+Ntv0uBz2J5mDmgEOgM3XLdCwbUv4fpbCMHDeCePBRwd/LBs1DxPumMc6lJ+u1s6O
kXgNE4sjcvlKyqHsaTcZqMn4Z1WS+dEah09Wypn2VXNC/HajG+6Oohz/1rkPjfiwpo1Y590bXFLJ
lZFcHY566aVyw7rSYs2zW0vxPhUw/OmF5PuZHmdb79gOzN5Tx4E3nRvSI+At67mUxTZaa3MknD9q
mgTvNJ+q+aHNaejEKec/hX/UNJrV2kRlEHIGl3j7maOo4lv8ljl1a0famsImkaOlLuv/jY4/Uezo
lUU47yh0KuKl/6NqgQAiY2JGd/feuY3/MZpMmq34EPObHZVhcmsOEtXUIvHEOx+Lr3ZodR5LLMc2
A/xQCMIZaC49etZJVgFi5UJ+nCzLRAeJ3AU97tuWG/nKUiAKtQexrIhBMTrp3Be93Wg4MOWVsras
HBx6m9nlDq6dxhQ4yEmgWuDtEO3toPi9RtpFOQ/mY1+hn8EMxTeulPgnsjh9Ac+23JenxTgz8+OD
/I4k4iSqU3/nKhw91uD5yXSsUj5FCwX5QPDsp39uogVwG0EGw0sITKWmyihBBhPJchR5hcJz0lMl
kmg7PN0uMjpgYtIMv+yomaujOOi0+de9hAQIHiLEtScYwNG06YLK/Zip8g5Mk6KMFf3gB+AynHxX
tfX2OJmxwn34nfvPOoI8EvVCj6yY6mAtZDZfbQlgqGeuB/VZM+rqMEQwMeDM1ztUWDpf+I0qaggQ
dPpKB+HtLKr43SPyWOv2MgXQ2T46O5gRaY5OcpDW1kWi0innKU0mTpEG1am6VBBpaLm8JWtHbFtN
pjKiD0FyPrZXvVu9QbR1UUxoJ+S2CT/an67Ie8ROEsubsspLc9d+wSgxze3mH/egQcqItU/3JOgS
Gwj7WgkiL1RaSW55oFBUznsdQ4i+VsqFXOkTK7yg93+QISuofwrRKdglDVTRI/m98Byn9KveDmLQ
B5wCvyxBz5PT2jMQ3vgxK7rkAP1kx7h+YxNdKCJA4+ttnvWLngdraLxhu7qW/DRDFi6adh74FRpB
jSPn6S/wmvklMciBvtevbAt66QfO+ltaoYDW00cexGnx22rr7Uv0BDIjXCk646NTlHY6wtjCSQVk
d85puCOCDk002TGfjIj5j9GFLsLhcqLICA4k1aJfblZ+2TkHN0bSVyHhsaa6vec0I2NX1ri2Hm5M
GF+pAZ+293FBDT/2jVuTH4PDzsZgIVRetXinMZFJ+Y+uqnyHX50YdtmPlLEDZjBM68eqSRCUoshg
hed4R2K/ZS9mv3m7Pd0lnuwHCVADlX8Ljl2dXkg5Ys2bDRLa5x2qe3LRRr/u865lF8rg6LzH+cnz
JF9o2E6E2KHNrf2/+rzBrtypAqkz4scdInZSWXZbU/t+MO5DMgXBwPsFh6nvk2KYGz+DqIP27AC4
BsH8Jg0OCXYXYayepFIbh8d3LRldn0Nr5X9BbVcT7dq4UrCL5dSxmOCoFeE7HVKTI9eguRMUY/QO
c9wBQkKQruk7udE3qCrAnN++RtxtE7stpMwyMB8gZOR16QAV0mWaA+TQmG3XDhPYtFXal03gCoaC
I5Mjkam8Zo8VHTp7xvDTFhKwPmBcPEd8PKkPVh0Wk+etBVhwYYSbQP8cEqMGsFlBmATLvUMGIl6d
msaG7Futs7v9R82IkFUKO60isW5mRVMdrU2uDgd/6zRd8l8rvqPfGVY80Qx/W69GVYQnIlKMkgSZ
oI/taspyJ87yhELplcnbf6bXFAgcxM8PEdVsD0XovIRyWRywVj1l1C/oTIiY6d7QotiBzqH34nc7
NfydtoxwrAbj3ZRjmOxSjolYiJ5KH42l1Hn9xe60AKAbujj1720GPXLnXYJdDU/d6EdfqMllZyxw
q0NDNgg2PWgmqqC5noNjIAXzGaR9YLd709KWjpayDqqQ/k9T2tAw6cmKnD/HAgOdsRTGGCJmIsrj
/BKh6HkF8ha2CF3eR2XPwRqn2gsQRIbUyq8PMmoL87NCoBPNO5JZ2w/BVoTwjFpafWrtv9e4+GMa
kaQmTZTuVyt1ZzinWb8d54/EV3a9SMz/uOFejjKQ81io8c1TsxnaMxO0bigdaRAi7mXjS6M6AXD7
AP719FGFMk7MeazUepb+I4I1QHcIFLHJXZb74e1FeYvXuO2ucWxVIWtTbyzlWALG2R8pNMkBV2ey
fi1nL6cRe6cSk6MdQpaT+Anp8XCQvcFq6Kskj4sR1WCvT1hcGQHd1vZ0qrGQX2XFPlm9udhEu83h
qPBOx84pXeCbDcJGh6cLT61VuP2zrUZjzBsrSH7+/+Ed6XUYZslb/te+wDm3bC1WKpRz9awDDjog
CeOg/52l6cjvahn4wz9kGx5pWqWajH68FPpuceALkJM0W6hkseZYl1Jxhx332wpE6gK2KLzaCxwC
K77uBFYrqzXHJljwbbJAcUnYaMOfbi+k8J6RM5/fmapjHoa0XtiMQh5k6BswjI61QXkJXXxaXnaM
lo6EEl0HRuybTw1j2WcB3fSFGaH0301okd+XU12WkXFS5R7PWdHy8EOIfkflhs/f+g8LtuBLt6HS
hr0Vqbh1JN02TvD88GoFd0t7e4PS9rO1CrzV4ZoZFVBAQpX+mPPv+IMEwx5RMIix0/04CeS05bQa
CCU65Ak3yy65WCe6lk1kUNLqXMjy8TjgOA2K3dKcTlZJHy7ifyXAHi6GuyEa1nuJ7YBKqEc1BRIG
uPwzY4ruKUt9rCBtTMqSddLNMZvXbL1bEzOQe+qjZlzRnB94YUoSkv0+onKBGHdAqxRs6MGvd+d0
58HWnkDeJsRYjPmOYFTPPdgsNp5n/wUeOb27NRHLggszV+NTSFXwwUK0F4qTMMAkAwgR1h0hjdwD
r8Rnxrn6pZnnuexlzrv8T1V0uipUsSS2kOi1TOR5vLeE/IvbeamAxFxdloqEX8Bv9vVsNJyrMsJy
qH4jVf7UkfmINvw24S5jaKPMezH0ZEsuhZfAIAxznuDwnYOkWO74LZ3dXPzl+ynbzh8jT0qL5B6e
X4ZVthRz8SeNZWxGQkXDB7RIzvfEpUF2xdMTpWwMlIvD6J2LjRvtICuZI8Gw4u2I8SBVUOcMreib
qC2azOgvnyH0idyYLxV3yGT2ZX+gIXA/icwrUVb9xRJ8vlW+cbvgBcz7WYD90AG/kEUnGpk0KyXj
vs7FhbyE/qbJFCjuCSWPx6ntfyBXgcZGYCd4PddV3G864d25/SZViHLiSZ8dHfh6RQE5h2l1p9lH
+emWStiNxKm/7i7R50oJbdCWlTvf9+vfb3nIJ5Rud66LnVpP7dJFMT44tp2IVYQHD5K0VMjvUcYn
hz7p5KwLojS9SDF8W6xMo25QFCHGSrAkwHh8RSFRQ86f7T9sGUHNhZYxZgOA4jKk+t2k7zi0Fkax
XI803QVmgMsAjSB9YeF01pR3vFnKQJhz8OYKdWWki8+LcMakUarZJF/duGBxQM/i3Ag2RDUNe4H4
rni8r+hPB1sp0djhZrIV9iqs3uyaZvHZWyUOxieB5QDfjKN1DLHKpaIR8MHYyRGtZiftiM8Ay1rC
Xc/hdpDzWHE76bpk0Z777GpFS1V8KvG19/iJZo7Mhgz18QtPGsWMScYZTV5wgFdt4M6kcDWqUaX3
XlTqlhKuV5yjHvsUj+GR3jPHRkmNT2BOQ8+ZnmoIY/3uIGr1NF3yLpiUDOyXHErrXC0LbI0KWNnG
kMMxABNXqM5bFPqCOz6a5JN0rH2YJiULTpvHtOZ0lWzfJGK/p+aY8fbRfag68MfRrlfoqqDJ3jDz
/zh9UbrJ9h5lzmqAR4x5Uyx2P+gN7O0wv/dyb456NcE0hqUXf8vugXZCIezlDsIQXOzuWRhmWTYR
pNJgcxLYFz0F2ji/FayNI6BtyIN3To2eLhFyHbnq0QllwgIAzDp4B9ZLIYsu3as4ZJ2PRI+CzCfg
9jEE0Ad4Jt9inaJ/DYPZg0ZC4f6Ajl4QuOLWV9RD/7TzoTlNv1ym77ab0MZL5Ncd/4Yv6Q/Afdd4
iKYh0Rgo87hmU5nq5KWt1ng/HAhqovKfbe2sasBIph7j/zR1NEcxNUkacCcMFPoa3fQ7/eZ7kUxP
dfIc5RAIESvAqxF/uACgJhH5DEHeK1ZLUUYlsbC+nzAnoU+vhH4PXI/wifk1PUVV0d5KOr1STa1G
JCFl+bxilC5LRua9KSMWzOiVD4VgEEtXj3cnoQ1DXehXB2o21ObXhheNUg+0ZusxV4VFmBWqt2uD
KrxEmWwp17sc8lZXN8tLi3YSPxOqwiYgWlIj5RXmK9XY5ufbsvK9Mh7miznKsuAK2d39DPH9i6Lg
ZytngE1xo6RoaLi3TaIl6U+BAJfXwV6dtUvmlDjxBVPt4JJkQPxyRFz3wQcJ8xRkFDJmxFeE7+8Q
OA0yhfQ3KV76s1RJv9GY+G5LnfOCGsWlsW71n48G46Pp526GjR4oz3/wdDE3ZlU6lFSavCOSPOpc
NaDboqfjrmWbNAIaie4gJvW8uXvh9Bj1qJouOvWjM/1IQUY7wHxdHDzqGifbY7C5s5PRavzjV1Cb
pa1TBIUYbCk3T5BDoSZezLVqyGDVbgsdgYkodGCPNvRa/97OtRG6I9f9XIZ41ln3/722FKCJTfCN
fXh6tMwzXF4/AIaH4qVrtjZQxGI58SJDmrVbnFAHG+xmJYkKLNZWCclKbZoHYEDJdXxj+Y6KmMI0
4o955hue6VfUZLtCqtka8f+yxDDw31eycnH7hOwi94LTlgBeTKGNTOXPEVTX0ycbxq19HhQmbK/n
nocL4a9bF/2yGgYbOM6TmQxb/fbXM4m9AucS/JxBf372cXVtxzrYbniZwthPbIz270RSjZ5ufUfo
NXKYHO+ghODXD6bumq4j/cJokoupy5NolFyMvmMIKDuawavIZk7hEjbDkLRjFKjcj2AvEL635n1B
d4MwmHPdo/1i9clrsjMZC20RK8Q/A4egV16SvZW8s2eeAPnsqNghYzt3u8ET+VfDehpHIRAQni8S
pG4Zt9T7K2q0PEBVs8vH4G2oHED/bf3+b94ojPmjjpUbHTDCoZkSwWzqa3EW4e38vKkh1qkrDs4o
sRrwKG1guiXDU1tpSY8x38etEd6hRrmMlC2qCp8o09e2Eu5SBQ5Tr7J5pXTUdkkvOWEngZWjNvE4
T/0FwyMfAKsYevHJhyyRfvLgdyiG6Z8c8mAcU6UobFck9lJ8dVAErkBr9M1My+9Wmq+tUIjXDToX
JG5r8JyPBFZ7/FfqGW0CKaDnFKni3b66S/+154VhwykvE7956JoRuf325mhtkKxPx6H8PFgkgevt
2zcL+zmL2ePIB/2bEP+TMleEzOqOiYV7E/jwIUH+UepAeE4d+kNkj8qrTNdLyTmE5VtQ0tDSQEgx
K2Mv/Y7R9JQh7eQDSVy2NZHBekF0Z1C/7wwgQtn8nfvy2SKhIyNWz5EJUa/QC8QDZa8eakOH+rXZ
gnNA0Se87WLkbSDmwr1DO1bFHWpI4pjVMOD3CrNn+TOobPtSz3GooccDwQBZTDwEVyOK3yVax+Td
+7UoMs6zKn8dNd7aQj6QbxFxRGSQPYSIEAQsuYb11w5KcQbNcDwBv+oMvlgCaJJtowmWr1Oz4OvF
mAhtsgDb9rmUsGcl0tPMIEL3OrNJVnUwG1mU+3AO9efBZ+DqxY6ynNoIrtK/6GonBEOGCS2f5gyU
ha16bXl6Nqt95dvg9trvb21RoMK3enB8ZLwGLNG4tjUV3hh7r5lkG6YwwMoqHkXnk3xDMbUIjm4M
YHm/RMw1nrdQtfgyg2qmR+0kbdNCSecm0qrRMgN8sxtC5wqNzsZgdBPc+R1QT0Tb+ALUC8gozgCV
YnkQC8tAiW2I30Ev7ObifxZCBRK6iEzzocuZCk40dg74qDsvXHZhm5YOPduqPS7Zbetfat2ZIG7a
xzkHjSGd1WFplHjgQ+hSpxGTZSU4mzeVkXVgps6c+ce5Eb2IjlHU1wINvCEqHRMAzUGFeQxHysBX
tSL4OAavCqRhNAPfqsRnO6YidGFCokVGxq73XkASm6sxviBVtPHRLfOKFSRJsiyTA1/b9l+JcwIh
LdHYv/qDxsqd/AH8m2wneER2xFPbB61lgtkBE9znc9w3K4plBMH8926YT48rhXUZ6lHCP2BXHxZ2
6kkXWq2bFGxoDauUzEZLsus5WUMziOBz6Pn9vpiCaikIalSeodhVAwlzPzKR5IV//++x5uflkxfG
CSqSh6WpZ/nBBmMInhibvamv7MztFzzK1GxNc72KqBMxclWShiEfpjFzHXY5OJBLqqbuSS3baPqo
ZKWaE21l8vy5BdC9oTxhMlzcmnCjGblKWMXdtfr0Rg9w8pNJ2aDXOU3mOwRlVeJoLdbh06y3D8Td
Og+t0bfdAqd9K30OrLiPh4BL2RTlmYiIY7cCs9MH/E0+le8xC+zp4SbAO/DFBpqAqwWWYCpfU0qq
WZfOoT0VnID9kMmQAekqYTKTh6XPR3f+CaIbJGt5ReGbGExxFe/roRHv5a1thoT/YqdBKKPP73Se
djMJwuhTCdDZsQFu3NBmnkkhF5iuEHSzIhWUkK1AfDTXKxkOTJdlrg17kc7wGVkoeMh7PvBD47Bb
PEvBuUDrCRbHvFj8pTFgUMmIBUmpWkCivG0OoSGWT3yFk5XWbV2ZMnDFaLiE2nw9+uXMMZb4EWPy
gxtwL+hJnx1/5Q3JwRSuqxAiVLa4ORhnEx1KImUrJ3eDoZ4trc4kYyhUNVeayzlZRTYW1glPB1TU
afbk1HpktceEmuKVZTemuX/Gw/AB5Tq9KuqmUmasVAlXjqIfZSYtlB065cvwrOO1JFZHmvUSDrGZ
Yc4a5enPIc9ZchvjB6Ot2ZbijLwuIXZ4hTnHkpySSjvl16XCds16nwuMrwXnI7knVKZIYVmzpSQ3
cTTm0CxLoASL9ZE9rMzd4+bAP1eeDbs5E0k5lpinUuWN8NIYUZJh//kI+AkzjWKuCeB6GgYLQk4e
K8qo8rGKFwDa63eUKhfr6x4OHTJzZhcooq122INvjabZfPy/UPayn679b/UkqHkuIlU7ki1k6bYU
GeUOx+dvD5yFNx0wi6a/C+bXVyuF1qA3rZ28laGqf6fon0KN3Gh47nsifzGJ01/HcXeXYtDEBjRu
9U9IDUo95hDv+muI5nXj1nIPtIjC9B+jE4dBBckUsQ/fPNCKwAHcZKabddaHOC+tGfE0HkjyT75i
saJXOqwzVw8Whbpsrvmiqy4ou/8+PC/25OJ5lfoSsi/NZUu4uIG1iI12HgnhKqp3WyrJWaKK7Qct
PUiZuOhPGnGgUm5YpYPecdLlUawvrB3517ZMlRp5iJpxP4luFZF6zEkVGP5spF9QtmdMmHsT3sXB
/7dzQlEWZbTqQ8dWYIpSroAaCuaxEaSGsNISdn+SbNGYk+CpXUHIkJvd9W7SkT+RHSmos4V6Pvzr
Ud67RxlP6+gYKs7yplkuE6F17dY2bf5wfSm3TGUHmoRQSisFrWrT/W/UW2zKyJFZtxSmtu0sb1zz
eMYvS81lYqJwpc6i+he49YyGx95c614jFb5DD7SILup34M/xmB6Rxvkz1tyJN8xZCHeCk/9adXZ8
GWpbwOxiTx+wG6UL/g8w+MX14LtZxRWxeUg3k9CD3/5ndbTo2LQaJ0NmVLM1BRJUQPiWw8BdOZ84
O66ATFwHUK1hIFJXiq3sS0xiOPlT4sv2UvJ0A/CWffQeJ9V5BaaqkCodtGU8EK5FNsR2Vgu3yiky
U6zu77zx7wBhmmRDPZKxFbIdMVctzWVf8K3Eu8KBCTsHXtDR8GEEJMge8JXLOaCHGZlxuQHCTXE1
oCcw0P2GUl/24viJjrXuHmamlyUui20lq5RSIF88Ow/Zq/6L6Qp5rh9djUB8w9qScRk4Is/hfBaF
PBUy+XG90AdFZWmwg6Upil1rHsquFPadj/h96xGBMMIh7zF3OLAbuR30R0yfGJiDbQ20AJaHBqTl
FU/T2U7PxDP0ZXDaxiqmMB/K3cPZPO/IrV+y9K5doNISaiUJMbJIfCJo1Lhsn8VGRNCrIPzqUlxD
N32TqHLeF4IgXACS6C3m7AVWxw5OkeL7rt/TJOPS9lErX5qNAp7aPc6pEpoEL+4ImO3vkVYwwmf3
NKOmIgQqsuKR4OADA5mRyWwHq95JWiQvOOGpqLUQcPgqBPgrFbXb29hyE0lNYRlqUEWA28jDNZlp
VOfZvEuTMRPWzsN/GqsjbQK0IVeaZNMV7NGbAscyneTuBVunOkxxZk7nGN0X/ICH3nY+k5NzPzkM
DNdj4HpSmBkDGmjxSGqOnDHZniOsQKI19iwcsB31bkKVQNSenrWKTvg9L8HDA2OxU7o0swYSZBLn
shU9QTYYuFQx0g3n6WN8W0frslNjpATUM7RDmwGQXLxH0WKOlnK6SyKLJOL9D5fLP/SGozlMWvCf
JsG/8KsM2RgRGe0vVlM9RWoFDnl3rNkXFN9QhhlJOGDwOoJgCXgAQj37ov6OTtk/gJUxPQxFBWWL
Czfl33y9sutn4BcSyY/FuX/kaQjHocXCv5KZ80gg1i/h65lvFrzPyDD6PhpPAsOFWUnvcwWRDRxe
IQUZ1HhhRPi8bz/7IelUy+NhmxBTNzoUe/oPlHQuJln4Wi5noPgCEiJaIsQ4/J2w3Gmszt4uzePy
6gCg96JH45U66yUmrZecctLGLmQZ37EqmDo67j1cevhvRc0/PLh09C9V/OX1LztAddIakpb8hOYA
Wojd03GTJWvnOZ1A7CK9oeGg5acwn0ns5Ykpvrwqe0dj7w4C8y8si6DKIVcvSrBJZN8wQj60Frez
81j5/6j7lXSldHogxbdyRqiRaIw2rL/HGqMcte9uvNsNrPf33qh17viQyKiDzy6qXU4Z3ytgtPPy
NvKIYqD/RyWftYGzq72m1qQe2t/Vdbtd+bpkYXBrjEpPcvsyDs+twsl9PsV8EdwIKv6Ek+0yDIFj
KvZN0i4wmxAqTHKDXTZwDWVk3uoTzZjoCdaGDsJbNFufB2rsCsgWlXqzA41n3JM844vWJN95lB+F
1A0qeoeWNTT+Ow0cmBbTB+ELsGPmz80jSX8AzuReeim7C9qj+fvJoXsfWTy0j1mrlLsVnncp/c8M
0Nb32YIrAl5StJE1BS13kfMQOj4Y0kmLQ0eeIxlouDbscXRXZnJ3Wg0fqU5TF1m0t2qqXbyDTaF8
luuUw850b5vCunTxt1+tUSsd5UqgXRmPl7v2nmKL1Pj3IIhqxLipVFaZ6pewz+Klwxb2miH2S9N+
wAoB7HKYMHaUXJkoDcOcamD9XAkw7T9dKfqn5xwgZfZ4eovDe/filiZIW9rHe7i2GBMOxg8ls2m8
I15Hi/HCquYbpzZAiLGlRhMFlJOGIz71Ak11Vp9XoXKchmm67znlIwDhaAxy6XOuO/wlDi0cxID0
1l9YHZfnxcp9eUW4FBUPi1ZpvFEumFIJasD+PAL/zX7g2sgcZ5dt3Mah0jtt2sRMNUxwOR2lCwjN
p592vuAkjrU0PgQN7SDrbEGs1V8Xxa8ApJL0S/6GBKxA8+yIOnAcLyZN7orlatmL8f4SjI8HtKG4
pwmYNnI2Ma9BtpH5dsnCqfCsZoXIgLy/MS9XxcTadxbd0WQKXSIH46mObxZBFVRMqXJCt+HGDVSK
TJ7baQPmfKPk0QGLJ84GS57sXhiT9GgMZeYUnGicQ8Ue76PU7Y/oue8GgHIf4nCk7fsmoZd1/d14
z/VKmA0/UiYl98Z69rmEobJSC6Ujk+f9vytjqanRPEmlXuS8vq8T9OGXHUHLvOuWGRn75IsfOmEG
oBHYbbpPWGdCXuoA/oG6dCbGCWsw80BqRxHW8xKPot9dWoY087ee5UqxxabTA1uSYzKpOI9hP6GV
JEiLo0LpRq/PslK2O/uIgXqqpyt+1oNTsiEh6PoqupEDwDpEiZj3sVHN46p/qdIG7UL6nTVaWzcV
yDhcwh1bWPXfc7nF/9i1v6OGhcdrmkwNhaxSZTsFnAT5wHoA6/kpdvOm3GROibggo8A99bTH+d0I
UbSVhyoEKW/Sh51hKU2pnSZ9MoBG72PxZ6/A+jQvauiZFgOXujAAsiFkIHMRt0LPefqOo71UAx6A
eZ9+ScctTCtYpT+KebmzVH2OtKScN/arQF0GkCdQPjs4XlFq3NjlL38l/whX1CTkWHeLFeyZObjA
V+1OXBYI4KCLtfF/MrVp0aGRUqwNGpJs+R4efZaSCzJ684Uqw8c5/BD41mxQVI8Hu7TnnXvitOQM
RPqnseOWLDIuE8GFSK0wRZ6bdgsUhuOiZMicz+UHVld6fIXXib2A4G4+joTPQTM4HctpHNx6dPkv
dQ67iADi46LUZNE9JaqhRCnf+VW9VrNiImpsFZRaet0Yne94/N5dZWaMgw6XLOKZh6GvYmsYvGTu
ZzzcxXFKIk07kEK1C3dbuBUQdkb4Sjb2hOy7Rtrb0b+IEaz3aynecLnwfpd5PKvr/FX28L5RFqww
jt4yrxamdXNEvl0I8+V1mZfupmaaWfG8UAEKYbK4UMjutjrDfWBk7KHZu+qMx903PgkZa1fYazfm
1nYdkAstpgPVTwIwTn8z9bGtsSkdKDNV73J4fcVGiTvn0VX7sew9FnlpPvegs9wUY6o2/WIqQFld
rK+p8Z26ZZvK2/Kqr/diat8RMSDTxDc0etnpZ8gIOWp7lnCBa6PkfjBgBxEXQ0UWpx++wYeEJnUf
4WxL/RKGIgf8P8MDfx8qBjjklf4+GY+s4EwT6ul6RELVcVrrGMXXiMXehvvVGIF+jIdIaTjz0DpL
1FWsBRAI5W9GInln4U4GzsgaKCy1VxS+cknMSmagVo4YXrl4Lx3LcPxwg0STZgh4TQ9ihQe8KDYF
GZ0a6AsS/0hZM+aWHAqAUYmnlXYA4uEnBw8atJQV/d6N4ZbnYUQN+AsBtbJw+CauqMtS1KBBCtkZ
S0+SWsptXBmri1nwy6xotQT2CoTkKzSEaHZOZAxPcY7gaYHWgU+6O78jQ+Gjh3eST4ljU76Ll5UH
GWsnL0a+vpt4HZ9lhjkdoBQKNhF55HdzjLXjlSgDoK6vkv0sAAImtat/wcMaDqFT2rlceRse2LJ0
Vk7VaRprw2I1djBMk3wYvbfIi3X6y53+ffeAos8+CB6nbi3T84pAXN2V7sMbsjkqy68ilvyNr1GL
lGslI0avoEJIo4S8EbHZCaUzDuiwf0DZXZXHv/GSvZL5Oml5lgdy610OwG3esZ3IyjlVjK6+rksV
KJGXhJPbaYyY/1WYmwi/hYngMqyrcAACIlhgAjx0q0HmJ3TZ22Plaanj1O+DzIknp1L4oPUqehdy
TkiYpuFfAOyl5J2cRM7OLz2muH4cfxwNORpo8Jd314S1lJ2XGWJEvEv9GV4KSylQvGPOdnSb48L9
nnwPo75WGD2xDwHxnqLthA62ULNS1+UI0HsxhnFfnZcnfNQiyq15RaOpkr1KP15je6/eHowIqbt/
CVarsWuiw+IEwdbShlTdXw7/sbwEQAXq00wgbkdHA3javTMmCd2SZ04z+UFdWoMj9UL9tBehiqvV
VrDZSNxrZzFW59oVw8Vk046zE98I7moVhZKPuQi/xeZgnxCrTelToPzq0vr4Tr22UoY1Sc/iXSq8
gJ4GW2eJkmoXOaMVwcmE+QhKPwMpVWKyq6ScfDjzOm0jMcBOvQp1vnhgpe4eKKuBc3y8ix7CcdG2
nsGhG2YW9mMxjLaiJ6Y4EiKCuGyzJI1q6JhVNIpLBoobFxy2ZERiSFHMHGCuKX5szvkv+RluvyUd
gxbyvEGp3xWr2ZWYNyYia8M/OYm+LNBCfe4B2FULC29mTNAn0HTMxWuucAPgqai0fm7c+bIZv8z5
KdIjN7hyM5yuQCfrlLnODFwbH0QwHZteWAvMMpT5pROeMfG4y4q/GPocZsK0XoCRZnWt+G6Zc2qT
tmZVcvzFezNL1c2fK+qTLX/0JJSAdE58LvBYiur8Bx7HnUs3jeKX2xA2O1+N6LEqZJDSBUcLNjUB
I9Cy3J6qUC0MP67t0UtWoVOq0SqlOssq55qaiOtiH46fZamZC92IdtnHyTfnobPDhBD+dBTsFvw4
HvPMP4bGKVLXdNBAzDBS10UY2D4cK/k/PQQ2YTaJ1vHsMh9wFT/iZpLiNnDaRaYguvAxfazuejPu
NMVT2AyY6rnF1APQLMOA3gwhcxwPgVOrLoAXn5NJ5MDWw+O/8MCjplGpwqYD5fWcOasYARjCev+W
ECK//4HwAe3sEyqoipunXKfjDvXXO5k7MmzqRb4/Eaf2pdB2GaSwflumNjPs+DSdEwwWRFvjs8AX
VUmCHOO992UnCoOnCFleLYjw/8pWRhtGUsNbri9IW1IiLy+VHjgBi7HhBakSFj6vtlvoEmVaRAFl
4IAQuqqi6YPzBpfzy4A9Rf3aUYlEE/lp/B2iFloBbsjeBWS2TXP/vlj0AwyMAnDzsjZ38Eci3QwP
uhDpWTqWh2wJzQeJmjDpCeKZBK2dp1+Jsl5PzDTeMUV4FI9DMt//0/Sg6gWOCuLOdvydYWTb3mYK
IXJSbDOuH8iSg7lVfFrQxTz4fOxEyCP3wuR527/nYvKltbuXIwI3j68N7AqsjwX1M4R4xwww86hI
yuZkLjUINNlbxbALoQlzpcKM7osPpB91vGzSzpCtdaBSnR6DdMMcPJDXG0XC7pQEXRQokeYvy7n5
9UUDY//oyN6n7w+FzC1MHf02Ib23xx2KAcdRGGlEg5JJTGe5YymWxOlqom6wMHcMePAFJk9jiBAb
/2CzjRucs8vZFkzay03ZQjqfhiSDK7luQlLa1J/CTH6e5nxalq54JDRs1m1Kg9fRPV2fQD9C9cg5
t1rbUnCovEK1XENujm+INrcMs22fq8z4mM0N6M00eftlf449NXBYg5RBB8nEZiKFpkD5mHaNs1sq
CmhYeTYQAl4PA5uNjCHYgd0IOXiTC52TZv/gOPY64OP5g+OeWaNlhaCPpHBVG7VykEVv46wU3G2m
89efxxpDQRG5kwKRttUCHFCJv/pZ/2emN52AnGehWIpTsJxQ1cxn5mG8Nlcx1/sIiC/aSoAcXfTh
wGSeEt0Pgn3a/6mhp4gQjUar7WzCP2kfcPMEdRbxkQusoyYAYYU3FOfJuB08ZtCrJ+MH2sVP/wkz
yPv65/ZKFBNoLETPpBbRGU7rOIBTKS6NDMsPKLarFzDhXRL15t8dJ6p7OQTz9vLYFttjQJIAP/F8
8hyNfORcab0gHU4BVJ+S+z/fnuBFcRaxrtafBRrLomGW7QbTUKuH9NHQacpxZrKNAh6YkTN6R0/q
vpQvbZlL3H4L04JWckQQAdSIMnH3EWP99l3w+apeZ6hN4FvkNINBK3/7XtKLp6cemX44QszzAjZr
MnHutWGePwvg3cBTcsRckbI6rjG0nybfC32kRWdguyd4+D2dmCOdJJiNOnIdvtKssnztpeApP6Uo
Km3sYlG511KQXBySzQH9x03ZMxMMt3UmqLXVRx72rhcL5GfiydxIjYmvfAFCa6SjspVWQeCse+IW
e8otM+5nsJVDEaLKn99KbWhcv4eQxBA9L5Un5Gl+aNQIcsGM8QC0tV5KiJ8o1oCsp1qGGhRNKp3Q
P2pdYY/HZp1qjZPeIlGFHGiuonz1IGeSRSjdmTBw/w8JPwlLV9ma5Ux7DyMudilb9pdkFE+pwfY2
lhLKfki1beIkzKFgHoIeSs0VlbLpwwdbK90xVqY7QVVEDDY7y/Pd9IUOGkdxdepAxevWOEpsTKrA
3LMtIBytUqqKZivIImmoS8SIelunvkTWXf441Khd4dgIqempiy/T3dz+FKy9WPLVNuZUySn4E5GS
PxD7um9FR7Qn5EQpce7pkuhHRX0w7dUiaYpRxwbC/0S8ssg3KWM+QZhcPErGOYthIckP5ZnsEG57
i1QGxX+h0Hqh6W74nFlguzHxlbMZbK3tT7iAK/7LJhO3i0pZeVyfR11vj+tUgo2WCGOfNcT2veO7
vE3Wf1N/knfgWD9J5z+V632BqB/IhGpMj4ukk86Bpgp2zQNEbfjsqYkZp5gFkGiZqvRsV0L9BNSx
P2Rz4g25LGQodFyVd9kluYz9D9b6pDUvIwPW6mvTbR7d905AZur1XDYuB00cgZ/211KhfVpAqTpP
RvJ6DpylBH2UnAUsQr65wYbmBtbTreUOTgzF+TF9B7Sh2E9KagDMDFg9wpkzsMQPOM8Exk6egJu+
XJPfVweZ/9ZLsdb8FgtfBiwxUHYtV+5Iv975WbTxrh7VALT/7n8+3QanzV9Mf6Lvnc48QkdN8hb0
MV+LviIJT5ytiLA5bobQFndJMj+psxnhZq78F9vy1XY4ApDaqr8uzmAPTfjGAWyOWgMYiwpBuY+p
Nc6dxWMEwxTlcsY8ytoZ9HSCgbR4cUUZtbcXjTNO3Ws1BpPYHQiZ84NWoQivmXyxAxVc0jej3BTK
AdPUqvWi5pSc1CnJI8KWb/E7mwyNAtPyZdAc/AmvBmJFj45D/tkSk8bK1DDopnkbxWpeOCAyGCNn
uWRcqrvxuhsWhdf0m453iJzHWsYSr+t0hqrzHrv4yfpUiTYPPdUixjNuH6ALeXcZgGH+AG96SeUs
r8sclw0y4lNo896ffKRW9+UDcfMpYwNq/cvySU52VXzKcASUpPsZAFewaMlCVj2XEVVJSjrH0n+A
JxGR5Yha8GWQp7lmHOoFMwBVNtsY0E8vN/ZISRswCAdJEALvkGH3vOfKsIpIxpvuE3QNdTcRFROE
WdQ2n5awSi3fNnwMj0v1+H6k7OgfAaCvpY+Tl8fZfqcdfj2a2xDtTPi2W1RaTdGrPjT5yVRuZcCN
xyKFJ9gtR47ieO8mlCm0a9tPtIRMplcul4ud2U4MBS4ABo2NpsANob64YQi5ClwNEhKC2jZNe3AI
3aE/SKrAmagLB65Hw135b1mtWE/eOXW4XBOVhbyc9mbyy/gJdH2V9wBN6jeF5aO668ziO7YcgkWR
w1la09U8M2Q+SOY69rOILRogiHzxzQBLoCfRoWpoNolAEzmtMMSSpqwfAIHUfRmxi43YOt9WzmDA
eioAuM4QZ/HP1JoemdY3CtxAFU588fNG7mFSiUyzMI+Lx3+cU2nxAoGcCmKH+juMJTMCn9H7mDIS
3wfc086iV9k1mCEXCh4xLfQgehkn8L+NyLjwgySwUWVDpPi/QoPdiLU6UGZsWQwoJHgf8FzNhtj2
+5i1TLPxQ8X4d25mVhdEuh6/rh7OxbF4TKpZvOApt3Xd4YFeWvgF/xQysraz5kd8v3hqG4720jR4
gBDTQj/8Pq4OVkGK9FUk9htkNenham5Xq+CcV8k1B+erKzO5fATE2a5RniSYSHGOwtXD6hLaK6Kv
JzvmongS39kVa8S2+tgo6A2oQBwsSLA6vqCPD+jVLT/doLjSDhENltS6qVLhjFgeK7s4yiYiIn/j
u/RhnQn4fWVdK3sBLhveMUivviQzz/xQ0Fa2pNEr6OnkBpO3YdrjmIinFcGAGLT43x0tDp34Y20O
LpOBLKyFlI+7TPaCZbpxjWcGTR66rG/kTKy+AwODf+GAfiUt+7EWXo1cZiJlzYUaN7cP7MnuhL/1
eaJKEed2HtkMSJRKc4NIkkVpZ+3GKBq+sMAGKzbUoIywQVXGU2EeNIb3ObMOZCMzpt2sRd7JYH9I
0MjuKXPC80Uzo4BD5lMvR275wXLNsilwKdd1cBA6CxZ/eDVhWC8kiabRhinzAy2zYjl5XdJEOG29
w0Q1tlefxF7OO6hZSknUa7QixzBVbQBcl1famK+r5YwU+3aSc9wSe1ikFTx1iNYKkdgf8Q1vkFFF
U2iGh4+LyAUDu9jURwAlEKPysU383q6iJ/XzAMfzl9ezSZCeGCgLWuN2x4cR5qHGIcrsE83tZOYW
o2DVN0zxPqUreiV3RPIcgm9lhQPFynoejntqQFJK+Y7vPI1cwtqVRawKiJ7f6y7+OzB3CG5acPvm
FOP3uKlJNoQJ2LbId5jawU7gupvAOadQAp1MaIgyBr3AiHcQ0XtqSBG3Fu/gSA2GJaq4+3GMCzeW
WXLJdYbeoYFhIzxevUXpnKTzMlumtsQOoU+w2fHG4u3z1OwOuWKxN49D7byMDaLBS6gPBYUcWtBX
NcdkV6bjuj+BzB0vp/CTe8O8yB4M7KrWIBZNR8YPJ4M0OqJTLCZIHoew6fZbHavNG9R7n7Hlxv+H
7smV3A12JO3c4tupo8jb0mL6RaRxBEzFA8REShkVYfHm1GX3NKX3wWuir2zR8ZgPvO/rMaZOaiK7
XnHeI82/gIgs+x2L8Q4zMS6i4g+v3NFIiFEnIViJXsbxZh2ugHJsbh8jv0/68y6vaCgGZUjzlSrk
Unhf8DR3tj/ITQvENmzXPEbzaQjg9CG1Ekx4XhP22YBW4Dz3Ugj9yX9P1DkL3NFIaj41B3lRDe5R
TkWNq8IIlqiEjRffveVMBc+S49Werp0pNQOx/O580AEkag4IMi5llTWHHjafScdT1DcPMngcoLSJ
odzfIjofSVDwuTmtSzUd4pGxK4PccOtiG8VxT8wrIv+PBo80aDUEogkTDUkB5EC8xKLMPiUUlywj
ACJeKafBPGa3MqX+Gz2xe+60cKM5p9RfmXW6S5C65hT1CRFKlffykSpSze2/6ivJbk5HcEQn4B6k
wpLOBublb+eABZDF6Pfujbfee6fbih3/zEui5A9gKllKFJFEn7n6t41sPnxlS0Na5Ip2Nc1dsXcl
i+Ke3xFppr/YTrLlt+m8jO5blRc+/XfP6gA2qBwgGaIxBJbOUa4X3elufcBVOtmrTzdXmdeGQXlb
oT6P7oPvTDkF1MYX1qS3azotHSk5vjEXUsKFaL0gxitM1l+Adjw4QY6wse/ctg+oPh4aJ8zBMIKy
mnR7zY3PLdSaU6stCtGfrZnT67yqUmA//xafVJ2JLZHAlloeUTTsuIaPI6kzY1ZUu6ivp5ngAo8S
OM9+eK6PAlnb7Mvz/RWEDT9VynzdyPl08QvYGddvZbhuP+ymqAEyXuX5LTCLEekzoqa4o0qDpo/e
H9sTNELtmM8uqEVkXzfBYLLsMMRxW0Jy8gxZq08M3C2Fa24jMleJ7TOudrL6Zd3BKYWsx9UELz8u
innuWlCk7OON7aClzMvxXmoEoMhm3NFsLsMEVlQWgzA1QT27youVQFMWuRY9HCeS7a/n1C/7VjPW
QzB5xoaM5eVdrBjmcQxONZuTQmww4ZMhUwQeoWWyz9iV9HcEcwwPnMnf4n92N3GjCKsKfnzFLhLj
3wErsTI/7UE2Aeu9ERJxJTebdSjf2389qJQ+49ijNJR3N2/Urknlzwxw1FpUlfCTy4wS7RJRVwlO
v+ehTqKpEsWp0rvF1KlkqxS3vHNHI+38NOsKnNEcyH0CgCdJx0cChqeiVFYYWjDakvM/Gf6wX7PH
xRP6OdAMz6jHNLxSNvGB8ZjplMyCSRmtvVZaKRHowH9t6XfwSXsj0XpffPrt53lnhqQMrIPcQf0x
+z71GKpOH3Qicxo1xzWCFu0CVY3dkmfP/Nql3eLyRCPOFJyDwpdgW95MfPB+/EctYauFegmpxMx8
RYV32a6mYXlNW7JiNW3SeiKs453vVRoza5tv8EmxKDQfGmjVAtVtLQ2wZTn0vzmt2MdvqbY14/pi
i4LjCtTbbHU90+VFg8AmG/J6r3WjClAdCaU9eDVD/++0MG8UNr39PY/CRiD8LhBnt9bJSldwYuH0
zt2g10MyqSlkOVPFZ9O3x2BNcj8EICyCAJgGDwvjGzGWOZPZoRgMXuD2zZaq7flc61haqClNxBFf
IS+wNAWe48nbNZxhpUO3/Bh141XGIN6cn847mcEv50tl2MzHruwh0FGGuUDeJgWXjU2PWhimaJEP
ld6FxVQzW6dI5unJHbI+xqeJwKkAZ7pr+OFoy/vHUQ1I1mj7Elo7vBGcjWDhSEka1xstcVUwYPXH
BGCRvZdLhVS0p+Mpq6ojnmIDOPqQ4SlyCVxNeAjv8ORMCUMs4CIfsOIrmRC3UNnL+YVlIOXRAXAx
lW6hl5jPQ2QD2dhzFd+lAktPz5qUATq4qMTpxj29HcMuuP7Ff9CTXwceR9EvF4ZL5F8K0178grZM
B/xkqBOqAPjjdQ5WhizXZca2wfXynKBBZXe58pQ4qBCwpTrlJcTBAN3MOtof4VCD6zgdXNPIpSnR
aQilcI+crIgTiDXUoeUWhVfROnbFI6cNhBRZlWCOX9o2cX8KDre6cJ9eNJHms/bqkmGO/hTMSC3O
uwakJgRyfKPUujL/5BN06q33kT0WyXM4kcw405ogsQ/mnBPRai/DXtRTQAg+cveoxC8bQv0aRwdw
+2o6nOJHXaHMPFIF+KNHDDGKofZI3SKEOXLjMnbCpEPklFB5aa/TlGVGiMaIsf29IFy81LJw7Ny5
Kl5pQ88Kfscle/McNygYlSFyX8nZVtpa4yTsU++Ewr4X2XP+fRzuD4dT9wLUuxiFo6TsO7GD38VZ
/Wcc45CI8aQjMwmuerg8veqcx7ctwGVeHylBT44S3Bjoy7bC7IDJbzd/KBNr8sZrcHONjM9/vJQ1
b/wAWcf1PInAY/xBO4Pv5DxFEkZ/bxN6b1AEt/0uhzfeJVmIX0Spu3V/99qiZ2iDc4ijDxSo2PVi
Q9QaDx0kvPVbWdOuraK9CCnSnvT9Rv326Jk0P+QwpcYzYATkeew3dN3DdPb2ERXabDPNQaw07umt
G4CYGxP7tPuFAcr0D3jbYkomEh8iMypEnw6XOhr+Cg//Gxq9eSRsSVbmkrPVX9Lg9VEL7pycyHl1
PEGMdYLJ8JVyDQ6VQfCoxSJIESbHr7oxRjTEkbnfOsS0mbEuAPofTPCbquIJu02V7+Q6rC6i3RbS
/k7qExHo9+gVqtfFjOJcJqAv9rpH7bJvkQU/Qo7aJJkI7DSjQ4YB1suySilAzDRryvo0AAd4da02
y/QOShEaIXQHSkzKXi27cxcvWkNwKaqOwKECjvrtMVv8Bf0MxQjeBVfhYgKOdtuNbQqLmdoZzLmX
HARb+GeHUoUCEnVyn6+Z9i1uPtDphuT3MJB91ioNj0+VQxb1WsPay/pjfbmq4seBPDtjpJ0zqQ8d
ivv74uVxB0vnz0JoGt+G9hzxnDxjVORUXDHJfqqWCr4vsSGGhtObAs/pSLer9x4IVxR7R4qHGMq8
DoLLUbNzunC2Tj0k+HnULcpl27xHxJqcUBolE49rq7dejoDrIad+2CuyyTOyi4jCv2+PYLD+zhP+
59VYvzFH4ZvWL7JP9Zn3I9e9UdMLH8sLapOHYAy9H6Rgp97mqm1Lfp7ml98CvvcqEEB8XJPzCckQ
HxM32CNifk0PuThzErdi8OXhcFUQwaXQoX+TrTgSfVuueCJG7UqerhwWyN0d6dx1I08EfB06Knn8
m/xcgTLuHOxrXDTfYsOrOdBfFAT5wQJDGdjnW2G4xctB7dOYxYb2c/Qsnp+zXD45yvzMU5ob0na2
QLbOib0xpr39D2sbnNZQTkCz5ytBpoi4S/Ulaei7Zyeff2y16eGSQsYwQFD4v/7Su/lKCqND/HUX
E7eRi1tIZf0jk1cau+TJOZgGnxCOwEGYQexWoB+ADu4iGhtip0/kCOMo0RHAEGy0QrlKxhiDXOoD
BsPNs8iyjjTKyfpdfqeMBaBb5/LPHQs7Aazm00V9AyWV1/qhA8xAQRraH3zkG/J2HpRH/24d5W9a
IPAXiGmYocETvEPqDWc2VjHxh0MZ0dRHJvgzgT5DBZGjxrap4uJxPFsBsA+Dy+7emPcZhvCnA+67
57F6YcgPooMPAe7hAdT6NSrQSsgJYRUSMWvY5mE8kG4LjAK5fca/SbQHJRTHeggyKGzQ9rzzvcxn
gSAbXAMJ75z0EyMhH2j6agSY8B/wzUBKYrim7jpKOVPEg7Y40VyCBsrPc5/FXx4X6o7IH+kLun4Z
3v2oySASQtrdTZDXif12XcEdhqvfAWQjZDhlvJ/zfEp1w09BN7FytnFCc9Id7xLHC/y/IvWMSiXI
0117w2vDfMoSFndWzV/x6JsRF9TU4Rzfva1eM7KmXJiTDcPrzkOOix4uLqtF7XHXr1i6K/+DALFu
qNN+uHxt6v+CFnNEhH5eAEi+IEGMad0qFP3o+UtXIaJdHMjct8TzhS0jI+0FmO3XezNwtTbv84BV
x1JnygHqR66opb6cs6baOYMZIvzwSWYDEn/gafBegxnQ4ssiG9AgRUxJNfNJWz6+PBhCNO85aq+2
JjR5RTtVFvXFka7SRN9TKMSwKuv763Mlp7lbHd36/T9hP7yZq/ffZGIfzVcZmgE5bXpeWT9G49Zu
Sstaz8hyPCamAIR1y+cKIntEMnEfm49fT0EisI9Sp8YTuC2RhuXXC1koB5+KIbKsE34TLjcAMok3
zAMhOWaRm/AIQK38afyWelPZy8CAYjcBCFzL3aNIr9TUxT0tW03zUuC9efMbbwi0VhqjUUWfvB0z
NLKYFTwvocKzfht81+ZXSkcuZcuPfzQlPhbAJ9/hQshJ0tUctnDlKzr4cHK7kBgrXpRYtW/CSro3
I5zpIS4sQAlKJTjBMJWgOyFNYr1XIgSxczi1QgHaJNozXkMxZBWzI845apIM0hx5Ly+zyZNxIgfv
AkQaosOAnJ2+7uuhfgF5AFkkucoNWSRg7qX5sdrtLbZXFpp5Z4YhDX4DVcnfRL+8PBBhA3eUEsLW
OchXrfyxolVGXKPNWpPCeDAtNLNck2euZcpCPMKlJOfjR8vCw0x7rFE/XJeu27Vc9oyJgpxC58xk
BUZC++jFLfrWs9gR6atOgJb072g7VJyloPsNIdFc14VS6JG0rByA249EkXwA+BgPiN4fxsY1XPt2
NDvHOI2lDsBARZq8is4E7IrLjWSG3jOi+nTkzZmmv5V9zNhsBXGlMVX+1QUBzViwacZOE/a6K1Dt
5lp9RKpr2YnvHKQixYN9qqDI4302inyRUsmt/szffIxYPwMDiVRA0XTrUgdhtUTMT9nRNw+FsAfq
+B0NvxJ/P/T/3fY56CRt3QrbsLxrbaJQDaXiuqjrkMY7npWtcmgQhAMYVcthqxm5r2OZq+kZq/aO
8j+b3x4Hn9VS3aw6ROWBoNkn8JHjiJGRTk0kpOi4qTXqUFQf3lvGkkP9H7XnKzM7fNTLD5hrXrcd
veis0a/aYgMU4MlKUPumVsv5+aNkjGoT4+Gh40PJ0UG9Wc+6o7ZNScIFen94hAryAc+ChHr4KOaU
w6QMyjtx8I3v6VttCLA9zHG4RzWOVhT9poY0egu5ArHxCcQKJtqSqC3nbSHDnG46vO5EaH/uxUtn
i5vskuvnojuaWx7BQvhWdI0I6667+mzhMwnULZZ2ngo4JVUXXpIyMjH9TrqcohQY3hT+ZUrY4oVi
VKurjsGPGXG3lQ1SloAcmBIxGVCvPFgC3UkVREKyji0rRY6dxhcel6jhDg52PFHlqOjAXfEnrpNw
/z/PAHP22EhVad5PyLKFxoLxxQU5FEcF5asRotoTxV7sj1gL74jwa9nbtMjYKfI4Kl9Qu9thel4B
AU8FzrsoAglokt8KT8S66TLbU2Tozkh646k+qkAEaQ/7mA6it7S+OcTwhPgzY1PqfEjLkaFbunfO
I/NRJI/XC9sESkD7qauqYiakJkcdGSBGuH1B7irc8yYfWRlG0VpAKjjozAKRhZAmXiXbEXmKfSkv
dyq9d0GBWhW2dR0XmPUFfi+AZGPo9R+9IujHpgfymaOjV8Fvu134r9nwrUDDvwt8nYmPFDa2fYIX
fTIsxQ8rfI5HHzQa63M4eLmnVrceHLXQzmxsKwrnymQ8E5JsGy8g2WpHoAxt7Bzt803V/7k1ie43
f68rCyYIBPOv4dVIGVoJPY8VX599RKKwJKVyeGbuWkyXgg3v4PxSJpzRF2QG/HKECEndOhiix8js
pyjQrGiVbaUpYLk3dbpOBsyXmSOyYFMOd0jatca8DzTdOtWxJL7ToQVGRMX+rbXnTP2L45UeeP0S
8DR+n8j7pDgZ4StMJh+KSo3w/ZWq+2wdLCCqMAsLpEWu3AknciCGi2oTrczPikaNbhahm0i9I6bD
eq6MOiBYaVpT+NH7e9JlP9L8uvKTqQEIc8Zh+9ay0D3hsW926W3rZtIOzMK0775TgOaMWd9Z3PTs
GWmBvA9UfOQm9GDzfuHFP5VTw1YhfwBYqQbcPt3csrC2G7azFR5OFsRiip87hHsqTuYO7PIulYlF
tVuxpkU30N31CVNYZdg/YiCG+jHfPGaKcUVGHhzaZEt8IKxjwebksLSVf3H36ShGrwYPLH4jr8F6
PYkZ8fw8f3/8wtHD0bxhAkbWG6/xFQBAutSdhzE7fXu+e+uHYGeFSnc/rXiFm9lZapw9GcDbAmvf
ckPvpz8oUBf0xZnpIrcCOHty9IlRocLIQpB2QsUfvI3FaV6tLoLAiu7RzV5DdoJwk4eThRphsGix
q4Go6X9zqHlFWI/KpUbrGJyGztQBNUtnsYVsHQNpCziTe/WSLRKBmvHLMnFpAi+slvs7uxAZnsPU
T86W2667EouXGgoWSkQY9vC2PKogkYzQa5gA7j5RBXaD05u9+YZYAOLsLeRBqoR4iO7wbRCqwXsz
VxTATwJuUuvw/GFFXP2vnEUh0kvyfaw6ZFcIXF/Go0n/UBFGA8Z5fLkowmMItbbJyiPofm+8T6eJ
oSOqscfQMu5IYZSrHRAl7RrCsbtZ9KCPu3yFK1rpLPunqodSg9ULT/Mt9XOTB8BZKjyz3oG9j6B3
YjnyRxh3vUIyZv9KG0SSCv6VQxkgAp5TiNck4AbQX5pvTTGH7rFnqwWxLDKpEyigpoMaRNO4W0BG
pz+GXSZPwlJ0o0MJJ4WyHmg7WlATXdwPlQ4Yw8sTcg9IkWFFw5vatuw4fxzjU251lqzfH9zh8ocl
69Ah4roN4RDqJftVVIviLbW2ZWmF10rGfOz2L0OXV7fBBEkDzx4nAbEbhhAhg64h+Y+htOY956zN
d0sq8y0VMBDTQM1HZe1T87hb7a7lHacMXhNBWuATBO0lS7ehOr3tg9Pmr5Cm6dNLH8abJj1e5wRE
IAyJEaEfUx047wxUr23mSqsbiFKhClMNDtOaxYZs97r3Dg9SoAdArYKxXInIakrwA31d7IsTj33r
pYiz5aL4IM7PruOzEzkSa/XB7+51SOqr33XAfiDk0xdJhuiwhZxF1+daHVe94sH6NajpwsQk4LIs
/lkWAaYpBi3JFXE6yzd93B3sXvOCUxUh8RXdSkYKG8c3doiy9QOKm+VXgMVTTg+KJ3+tE4cF4Qzt
67zeCmhVRrLUzXZBA7cLg0A81FV3szkO/FWQVwmxUQCmJedo1kVDUJPvkcTmlqGNjMt52TjcaU24
RXX/C+RITBpGsLBaB9LW+dvXE00OiKqkvZgt4Rgm40qc7IfuSZ8k4xiuDJm+0JQ5UzvxHQOxzgv3
j+zuQEm5dXGTWiCfeWPlGBEUHxdYrgmClRAanxkV2xVWK2UDu0OG0jHd8/uR8TO9FNBeUGcVQFf6
7rNRjwLJleB4T0QUbtKWHkjjXfRPFxCLLrnwgS0qGo4VgYoa4Cf0clXNzZDpvxkAjR71IMSi1/rS
ABoYqE4dby/yHZStJJoa+h8LVdU6MTXEj/T2ETd6stElwDd3RIAOWUpuR8TTxo2RdDogymfkqjDl
9eHZMG1AF9PtyfSPEQce9QIbIAr9cc6Af8w9dgugS8qXhQdy15/6ozh7nRsACWLnRE1I3ErtCzxI
iXawjHbVLV9gfVfBtYZcZ3jR1F19wXfnH2/BzlFxEB9bQgvYdxbwy6E4JXsA6slKLsV+01RHCwmF
XSPZmSS5xZogmAPdTguXOQbzlFfpeaaXQzS8YBODD0H8GfBZIiw5ufy5vdH0NObI1r8eAs5u2qC+
u7TkDqijSchpIjBIALdfss7Bi68KZyALxpAktXFrycMVCNd0TilP9w86hpDrS1hafEAxF9IY9WGb
nJjJ9mBZsOt/ZfRlCPMsoohZ88gdEbb+V4gZYNmeuuIaKNoka+99t6D6r4Q83StKX1B7NbryUvGr
avyy/z6T8utl47maXJiauNnoyXWlMSl1XtFRAMxlmzOutH/w0/+DKS8EGcVM+T6LK9WWpSRyYqFE
IVFyOGYdlb/FDOenanrBJq2FAO8to0qDBMKSxtrQRzRLNNabAPWyhvI4BQ03NzfcbvoVXQ/7JzTd
eIjl6Mdk83clWiDLBa+Ay0qg2bKfOL66r3m8z7Bt+XNXnEWC3uyQhdvoVLR9/qd5FSrqApa9E709
3QIDX30XwQmgF1YMrropGhYBTQpeWVY8NSiwkMrl3P6W7fzBRDubEw/kforqoJu4+itRl8lcsSET
PGfMDssHHshuhYTL+kKn7qSka08AZh4d7Alt94QQZNU0PW3c8HUnrJXKoDDbGFPBi3iKlXmDcNhb
rO/9QAQ+i3mQ1bYyMql3UV1XZ6JxskFhJN/rzNYJONg6NwEUvf0qeshj0yVqG4gCOYiE1gzpuV06
TVmazig+8VAzZYU34i06GwB1DKZ+ntJS/hSDO1bx6JgGdotQdU5Z1V+gbmqako94YoU7s0nk1e3v
1MmvDu48Y/1zDr6TWtsQYI1yDj3DTSy5TkcUPB5becjxr3sGhOxfSvQEp+4Avh92sMJGyiuylUUl
egLglshjAEcyZdDsbLqA/i9Lhwmd023Pb1qh93U5tbyoRDdbm8d+Rgky1tA/bYCRGN9t95lI/ki1
kaUW/sXabfJrhh++gJ7uYeco5Y7J+dDOlsekuZwPWZbtZpPmjC9JBy7jSkU9w5ITmr49mR5hW9Rw
D/3I2F7UCqz7aHQKZsU97M2IU6j9cM0QXeXmTzatDspTkClakd2OR4gmp1YC0Wbcx8JmkHj+7z6K
3Rax5uYrDx86s42xpVOzcGnqK+nHfThIdIMNHoZYYHLa3RrNw+Z/y+miNQYcbYpLPOm2e4G6A/DH
5CAz1uUwMgc228uYFYH9sD4hkAtqyLDdMJHkzvZYYP7wMx3pBwNfPCrzw5i+n4esWWEuNkbIS7j/
jjAYealovjT0zyHbBbqBmC46SqxmuOr1dFBkrPmk3606rwONRs0L5cnE+0VmhUAAXwxG9LaKk4Ac
+GcyIZchAKmQaIAY2JZ5on4k/HYuMDBx572JyjttTTNDiZdY46EuJYTT2jhgK8/x4pgbx0ffEID7
EPdq/wI591aBQ5SCDUUjHaeNXv6DXfc3RD/uDYS2IhtJ8xyOau20j1M6SVy1aCWi9uoQrV5ol68Z
IiaZKko18Y21Ld52eulVoeqpZOTDo21nojpt3NNmk92oYCBmQeGUWHZhtjE1MQTkOxkiMSrrrbrB
88YTVfJr9FCMOvDNrCE/oUyFXxL2ISmzE0Z4v+Jh1sGNH4p6a+RDVl38xSvYgiyNlXH7vPUv6jYY
1lLnUrcQAr7rRnkszEv0ExAjKjwFfxig+jUMFzm4hrKJAt1S4bBJv+BQh4b+B7Ay3OK3RoeNb5w8
/FBLOPxDSRujOAgEaQRbWmnREU5GLo+Theb1pvim49i+OoAyG5UYAzpsvu+AdLcq1Z2zm9a46Gfe
U1hAKEb/FE0fI6AGmKp+4V95pcnUvbZK+ZPpcjJGMAr82tpnSpQKsPtK/WPAlFC2geEIlaic/pNt
f5RFESquBI+czOs1jkpPVWtx3B6YfH7BRhX8diuYoK6R2kqojq2Wru3faHtQ78iC6zoTyvzuQL3q
7cqPBahdWCbXBY2FFqdXtUMQ9+UDldBG0qhhJyMw/AK2xmiSCE3Of9g9dUetKeokU81eZn0RATxB
SKj9Cukc3cLT0W+JgNyhoOrI50BziNXw+3Iq4+km74vmhECMvZF9VcJOUNwgIWFNJLc8/JuMeYab
l406ioVCso5hvojcqkreHjkE1jl1Q1perHEugEts644sXs6po//6AepymGibP+jTnBOecOcBTgh9
vQ5GhXwDzdNHx50S3QUM1HVJx3AOkV/BD8JpgzsfbzUUCzMy7uoWYjlJnaX8VNCrraV49CL1dNu8
SCzOIr+UcHITUyIf1rjLLJeLsgZRU70l8BUAHxqVYY00ZLR9X57hBDCIsWdSRQ2W96dwcLseVikT
3h3ksq08OM00iaONDLIH7eB3Hy3uUqysR4pvVvqL24JqqWbGIE7j8lcpLUS27dt+k1nZu9rYb9Yj
lqNk3qhVd2EzIW3uxyVxnqS6dMvFia8DQDtIUSw40Xc+ZYHLDmuA18IAXM61NIWWxwVP+e0bz7MR
ztGneq3guHjzPtJJ4/QO7nwMEzpBJdgJ6fCis7fXZPq2j9uIbP/CjDWvO1ZiysQiCg+/auNDZNO1
bRwegj10Cfag2/d2ARt7gMFie1C17RmI4iGusY5dUhVoJ3rXNJh8jMXqs8s7pQAj7oYnymUElO2m
V9INoA896exeLW8vFgsSRPempTyHkVQ2S2QrNBBQw7LHPQ+lpgyBr6yhGno7rTYZI/ESqWksteVy
XjQ3onX6ZC+qMAI4FqMe608xns7wYMNEFWaftlypUK4wGEueYV53xrFZks5v2NvpfmIysYYbnLav
D8/HM3R5E1I2rHkNGgYNxSgELLH5NW1t7N+kRqfGPU68reS4Ly3iDMzwHZTV47nftk8h/2dKVLv7
ux25Fc0fiBvfgxMj7yeSrezAyC8Jl8hE1qN58VXSdeut4yODyISDmPs2haz6/lpEyTp9jnHw2iP0
kQuh5p7e5qU52KTZZ/y8pD+Boy+269TRsZYT60EIs4H0pmniekAC/g4KAJxEwXn/lvi4UIfWxHeU
tI0joDDIO9DEaeEOb7iW9pRnNOWw0CWXqmhnRzInjODVVI4/zfKUrbOsyuvHuItmXwfwVnPc46uE
Kelx3naRFzbS2K8r10RNzc4Rhmjc94QTIVNOkIKC4zEP+gh8w/UcsA+tPwKliiFQjIf9Hvb3a0Kw
V5IGZ4DQ/BNnQfcM6o5+h9w3Rzse2U6MMveRkMVvCGYYvmTyfBZVVvz1CT1zGmpwVkCwzIrkYg25
/Y5d8OwJel5PSEePcoo++CTgj7t5oJVCWDiILUoRJ67VEmJMAjXmQwXFzcJHjN2XJiJOd2KBiLuq
Rjvk43DvJfzjRhBznwXFt2mrZnkOBWcE9B0XSFBC78LbrfgP7fir7u4py4hPSLJU63khZ6scecNr
iMVLUMAwBvLDqLlRzaReo+KYU/NVW9qa22CKmvvSTGqZf/O3JDzYjkQPLgbT/79rP/gtNolZaw4q
ZCQ6TOSsIr2BHPk6O4qEtt2SKRxngnpyloiIJ1qQCMEbDIj7MwvZ9sx142SBve7qxMuIK1d32D3/
ecxyG5xqS8Ngfm+dWayJwqULNi9J2E4zPZP9oeG0u/xRT+Hg9gHaTc1V8F8NKJRRSrZ3+b8Wnwzb
FaZv4wlOZBZFW5sLZv5V3njsegyvu5DYYXBzmd9ZGeuVOYBxEB24szqzjynxRdeNRFLNVn7MB1uW
wW2Pd/yRnXdEpEL7pXnOxCUCXWc1Mg8M7agUFDoNkJyB6+QdVwtyRcGAoj0yODTMxcotOY72XHkJ
TDys2wY8TKmy3VxXaveuKyVKylFQcMRN1YK6l3eYItJD6hTMH4Ue+GEIsaVaFF6ByUGCpQSirXir
RswwxJ6Gz3v3veNsbRxEbOEOTSUOns+gR+Jkj3EmXuX6yGEJl2pNOJnwI4bZJGJ6cY/K3qfrEccV
r8W0AC/dkzpfiq/GUbV4vhDVQrJpNnpbr8MwNP9UHIRCPwsZS0/Nn+Q5UCAHU8wY61vY4mYyPQlL
FPTzAap2aM8Ez8qsr0eqKMSjgeHkfrxWjcoRTjQ3mYi+GmNLDkFP6/E3ssAs2gGmGW/PW8pHJAnp
F1Lg2NYTQqVVnKsvxF716FDXXz9d2wrtn8yCK4wI27gDQxON5VsR2GC1rm8R1AuOj9h4OA6zCiUZ
1Ytw/g3+SMgX30jdmnBffpFhWeEAV0Z3gEwN/19LV8aYkEyuVjj16r3/qFdkPMunEJXdccOC4mnd
UbxyEw/DUg6BjE3c0v5ZufGZ+W+t+zOJ7tDh9ri2ks5Pnzx+0iU8ifnLfVMjS4P9YqQiodYePe9J
fbaIdQEazKXFAIPEEtYDPhFXJ5QBTYKZOCxkqfnNt8ABvEn52xQphCDPDLiKnTAHYFIioJN4EmuB
38XJwYzOyltcPXMJRsluoj9RKFbuQJf5DZmzxJTSznqLbyPuSeFWTawxyS24weGsdsytSfzOCWPC
sHyrDoAlYyAhhxCEVSLOVnySthcr6HQZKMabWDVa+0hmsEPcJ9qUIF2q85xcs3rrvBMAitXAuwv9
U7rCyXT4fWgYxWIiUSjz19tm2gowaz/64ze/E/Rcq4eAT5vWKaXB3kxXt/850Yz34j5PUcXBf1Um
A19O+Zs7ZmWntiqBtuQD1Ysqko88FReycWT1/6gOCLfgOm2lGaR6JLQmo1+4mNblpbsYvnBEwuo2
P/rxVI8Dzd9j8VWdfGtGvfLqOarKHNu8TTg0Es1WNw5JtTIeWChB6UVlC6Mjp/u5D8C1jcrCmgc5
WJkYhfyiL/RTmgT0thXULoDIIq1wm2GisZDlE/Es0Py/2g0T5JjnRPkBWaKjAArS8CyGjBfvkS6x
B7buqxN06Hxz6+CtY99H2W5VGNCKFCEGDcbVqJ3orjK5LETNay7Chmu9+TzUy3Fp9IQYrFy0Cig7
c438X/7f8walCQqYXj9JXoidj6wQ+iD4V5Pgl8bvnN3g6QS9haVG2/PGmKhBZUWwFCgawUymnUC3
gl/4VLCE0iwbIgoXRXuoCvvp8GuK5njPmn1SdUXGfEDB9b2BcVJQ3yXRnM+S8Ieq/9V6dTt9Z4a7
WmRzUheQV70Urv8Eu6ul48vbQSJSJobzF/vXA1UpxIR58vwsHUP7MdtzGoPsll8vyVdnMwSWMVbT
uanV5WjHMqEHYu991Jvhio9ygK+M2laNvdBCIgt3B4yAo7w2Gz8mCh85TssGdBbHy8mDoPNMBd+e
PiTlGDP5VUKEf5ht0KvZWTygHEgMoOuLUEY2c5K6B/lbLADSOIQoKeDN5Gi8bEuYNE7jZeSVzqVZ
/8CHVJtJgd5Twx1oE9HbmLE/qXQDTMGotxJ5Uodl/B9zFpcn9z3TUJzvWaCX+zc2ZExa2sC8ORvA
w5g50+LdFOF7aU4e0faPHOxE5fKFstFVpSowZj4LVmGd+UDNREeNo4Tt5ONnQMNj32oGRWFIlr+3
m94khc9b4zBn4wEyoa2CuLgW1IhuQ8gXPPpofvusy6mezG7AMC4o830pxfsKYGP41oWn4FdXIg6i
MqLrI+OUkCeYn7mymjgiDkrIy5+OUFlanPJUffGEVd0LA2GS6IhPR1yp/zVNPlqp7l2rnBx67wuR
lM5l9FFPE9wYo07uqOVnvuf6irTPlJpWGS65jTNeriEgR4wjruiNadHPgyEkad7XPvMwfQkKtr74
bVJpj7lc1nKm1vcZrMJeLcBlIgSBwWCh1pByq/PpzRHIpkYYiQF+fxfN1wEowaagAZnDIPCupLlV
DAX44TVaJlvHD8IIMCGs8sTbTjys0ff54hjbFUgiFd/6c76KG9UvFhFpKGrvb0YG7pG+tC49kKhE
/3lU65A1eI48TcUubnasDWlSPH4QcjQQF1JKvSGHljoa0v0ktJepRu3lYsHulbTOEVUmHMjDXjmM
QglbuLZR3cPmAMXQVvGHDGZngl7xzeby37KHfOJDrMs3Ktd9j6dFZG4HE1bC/ikbap6MCewuvi6k
vRGdLPgOtWYdl6uutWqHw1z6qIt/zTA8XW9hbRmBNYN0rXoMvx3JxDVmNBSIbGzfPjZvTV/1tbjr
ellY1HrVobeugnGWQtZcHqMukjnTPdscOri7MEPtwJYoULkXHIM/kWofwLlUNDOKfKfQXEj4EE0w
HMjaxEMv+l1N2CGBWbKHTCRsMamnQ3JeqwC+cOG70AryyfDxFeDQwbEUTVVZIP++WaN4BBV3yDhq
Sera5b8LlafEanyAGHb8wChuluIOyx03Kt8nzFK8+GMpePE3NgAHUUa2QWomtEn7bINib+gwB0XX
tJ4gZel0qm47sBdQVD1eGgh0xuK7eVoXG3sKhuhj6nbZCsWjIk6BZ/AFxhSP/stA6bTEbXJquEtM
hChGjjk0n00BvbtZOv6j97IUl8N+g4pUZ6AAyjauuSiM5NLOeceBVS6ORGJ/qGPDXO4MJUkqDWB8
q/o6Utk8HPKq02xjAHNbmZ1czhocEg9VX8KTCHiyLmUjR8u6pnrYM1MxLrdsCXvrS1Hy8WkrUi2S
0XAYe/QOUWPjPbrhZPobmVNboJv8RT2qGg4I06hTmdYUHJkHVh+snXhrHz+VzWs3y58yaRPvy8DU
FvUlg+yZpx5dx3BB8MnMmypNjO0aRZUBusd/xO2pST5oBSZg1kdByW+hqq9IPh2otk0oFzNE2eZE
i+kNC31iAJ5wZ22qHR09wSJvu4x+rcI8uUYo3uEE/KrG+jO3D9g0DuUcNm2L4V0L1Dod+Oi9w4gu
UJoFIiLMhu9T5k1+JRSHEOOYIz1IfMELY/AijlwYhRjffpPtCqrbAYVZDmbNGtnUFFyON7nzUvwH
sXx4z4wp9cFWYcGF5Y/ssqJg1ZK4p9d5SUUimkK8w9Ssq6FHjptFQeWlWKwvuuoWuCmJjXmufbWj
LV0+4fXzy3MJK+Rj+vzHoEwlGxhJT3tYLSSf1iv+Mm7Cldek1RJBjCOXrMUqU4dUMrFS0WUJ6dtg
QLtN561UO4GxJr5bQFxBUR1Zu5Rpw3Lqm7sjxMKHwBuIMBroaxRmvH+MBBt3I2aTVL6bgW82sjzt
ZzubjeFafSfgfMtOgAWnAFriFT9gEfUgijmviyFAWAPzX1qcolMka/d7C0fModLI5YJb0yWroT4H
GlxjPPDU4FuJpRyUNf8vPRn339hYcpMJlyAf5Xtw2tg7bPaHwpNtLH2Jp2n9DmOEahlKmRviTGjL
ElSKwcVc4ATdvikcLMrB2i409D3U6LkNVwfbjAq74JBiSkl0y3OMNtvlKY9NOdWr2hjh+5TWq+5b
fAlJ2p4uCCBbAYGfX1nR03jCTR3MWhQzHf9LdVIO35jWN8AdWUpUzfe4+SB0rN5c4bAeHZEKDD6+
+zoJpQP5jw/XKotHyEb18lIZMhDExhALvFk6o2DqBwkbr7YLG9HmegjED7Db/6OsyqcQ4GU+sauG
GKLvkvErDDGYh38X82irJnzn+gszbAUUUV+N7hHtPnUe3DdGrpHM5x6p3mJmLrjfTYcuvlEvkCUh
5otWigkpSLlJF2LToatwwFBbtaQaZr3PpBL2ALJ98He2OqDd9R7XEVWITQdUvjRwtjzmuAULGLv2
vS3JYb0VW70rQbtCf4R3KrpeUcRxiBhCv//ZxlP9wsfBtoVFRymLmG1PR3roqK84oaHa/MSKYq+N
YDDzDyDg9dCTswCgTYFmZi6ezECrU1zf6PMzmAulupzqgE1cXDlJXNccZb8zDORjlaIC54D8YU2H
FGLydCRKnvXV7dpOu1/W8y2XT8pR9Rowld4aQ5MsONLhNepDbDdTw4nl4z9CulxUO7ZifPLa1Zgi
QebG1sFzaZO+6/wSLiJxFLkJNZk8oNnZ8QwwnhjLRHaDYFi9YLnH3TAPhaDCah+8IFZvqtNnTRRk
FbZt2FCpWnebAxqNfypWISEkq6IMzCRfQLu+U4jcKZNIUdzJ0FY1EdPrNjbAjsU1XQhDJ7/VqA8n
2++VXhRvRYUq77MfQA2+nGSjKjGgH0GU+tSf3w6tEtUY3mU3Q8o6s6OY2u+oDPoDR33npV+p06Re
dgjA5Kmce9nIffSipiHAcdOD//V/+5NtfyPrJallzJb9p16up+fIFXyZTIYXzRO7MJ32EO/EmmhY
E1dLkSg/6e4PCbK2vXjY2yCKW+RKSFAEJMJOw3eKmk0Eba9iTbTY40a/q+SnyF3noMwGvM3RPt+K
S5HKxsByXyiIP0VLqPlvIcrvvzmpVIGiAn/Tn0IQZ/tXXKeNnd2S9webwk8038nVfwbFF0LRmCGG
f7Zkix+TXLaYC34yTYAWkFMjlDuBCAqEZaKt4aOrSndYj9m1UYEhsh6rlKIZGgBrC8zBywmUyhV+
X/zOiYoAvzvAnd3tVH+hsrqJxqsBusjDdeJMaJQjsf+Me48HG1PdtfJwkTg3oVN/T8t2uLrSs2ZT
+xc+tSivYUnhctuZ4SWuig2KaoVkkZmJJ0Zc7+b0DU3LP6evxY8bB/KwQ+Xpr+YZgJo9zEHsSpxf
ZioOh8gq/MePbgRQzdYjziHHq+cXL1m6Vj8AaxotUnPxaV0/vIPixx4x5fi4ClQ3G3tHVOVPn5Hz
3DrKonyLMVZzzsrKpSUpevAHfiipSXOM2k0SNShYLBF4WaNjB/mpGy029fFHrABy6zJNDIFxU0oY
ZNvALLgDx2e0x6ocOWnE1lkBYwvPIKDpsSQmkoeUhAUi320x7+xgx7pvB6xopuEp3OwsWNcRUtRz
5zBax4R0ABiV53kwjukoOGHOk3jTmni8LpSYAv1gqE9qEKaBEg6ht9IBanFMMwMT9hLzBegEiyhg
1Ua1l74NgawmaTiKh/5EowHlfGS8Xt9JL8b7xQvXdwhqQdxBYCWpyQDqK2nWTDA4KrV31GfDzl31
FYJEx5VxSNnNFztml80Pf8KsCsBGAWET4K+7aUl1z9XYpnTvIUJwgKLblnkQh65ONzpJB2SJdg6d
ufR722OnVo0k8c6XDkeX0DPbzSWONFPnKYN0jwYTitYwHLlf3AguvGUGdiOgtQY9ds9Z5P7+9YKQ
YpSp3xpL+pzrx+iBanEP3Nl+xjdzv0vUjSY1WADDEnXSgcb3tqZu3qa0HISsKWvoXCxA91s12XCF
/gVCH2u0JwRlCLNUgh3ogBhPnilqkl5UEsEvf02NYOdZF9jU8wZeZXmkTmq2NeptVpX2sZSp8QMG
trxhk1KLfi0jjCM684DL2Eih4jbb/WPxPg0p6dhBKVR5qoEHX+2Zp1bpzPIxoFLbeYaPUiyWRmlw
iRvKF6O+b4HFg8O0A4Paz10RetMMb+QgX3dVLzgWyV0nAiAdW1sdB8W+eieBqpw4PWjB7ZjuchxT
DFmG3+6+8TM8KcgnOHbO0CWTWYjCxoihv6CZQ0p+ZvWpB5kA1ufcxpEr43jdhvLz3cixTm8LKYlS
FV06hbyUDQqz2k9KASaSxFDS+W2aG6P5r3G+usOCFTg/2CN/b1OY9qKm6E4ZY/sw9+kzHNQk275L
DWL0FmaMxPnInJDcct2oWzDgS/K8e+tsL7uW5X8pKsL8mVS5V+bqY9X4Ck+GqIACAa6q4974LLKW
UaOxtJlGzAN/YZE7JKxKgqpia8ezctidwRd4+hYRi2p8fjo8NkVIyXU1jEdf7iD5vAlHZd6E1DOk
jicflfW/q3Cc1yylO/S7bOG3tAXahjOMnP2jR2C5LLSJlSQdqEW9NIvtKSWKxPlDZRXkV5EoFYt4
/+S+9oEYJ4+xipzM+Cu6O3TLE46bz/d6Y4WRW3dTKM75m6ArTZwBOMJk0IyQRyYdOLchV4M/p+ml
R/jFHtcYpdgLI+TEYKzHTQ6k7cHhx1atLfalElUq2E83J0rz/bb9/DhLklTsQRm+vWRXoRDB5zqL
zy8zR3HR2OhoDF2pCbbt/JZLqexJos7qHGfJgqOqe5O2AyULbZtlFO/AvrYpv1iq0GZgtfyUyE5o
1CxQgjZyN8G8pY3ePcCXNrFUtpv5kama/LQUoGDt2a/fH/4elFSOkB5muVaXv1hAy1HE9GtpM0Je
FITFGJw7/EzKH5DhpGSnAIy3EO1ga2tmfvEpIX78DiaOS/xjJpygYsdSvGOTLQRBrpXSrq981gPq
Lex7wpk5rJB64YciaZ5gybeg3lNOSWmU5QEecFiHuQWNDjFsSkOHZMImmBveXlHwQpsJanQQnbBT
ZwajWK2jxsq1CiX8WWhBz/x4PnIuj0Jc1EW8hncD95VIuBqO0p7Vuiy1fHmp+ZTHyP5cRxQ5SfDD
4vVsd3ejP2yhAuXfKpDmvZG8kTQwqgLa74Qp3IZEwaAwH3gT9LQk2xkstqFlc8yDmMJrouMAmTjB
/WzLN4Es/+Fk5a375FGxYZUkhSNpCd1wZHpy4xEFywhqz/Pksoc44f8lhNRlbfdLmxUkMNruy55S
6/8tWwBiPYubsEoBHcgfEl2NWISV1iaVdtV8mm1/vUrDQrqccllVSDoDK/SzD84EV47IHic2LRF8
SqIR5fa+ttSjmlXJuxVU4RrQYZTJAU628wS4VxGwHC76vYUB1AFkr/VPmz3ljr8WIkksUQDBZJY5
uxBzjtX+cOAEdJQ94uV1YV2JM2NFWgSC71kW+pYVsK6EuUzLRfVA+WsuUXYLVUGLJNsp8QxiKdYs
uKObp+OEVlZr+eTeCjGgFbfcWSI/NP+RhT9UAhsfnUGnWw46iJXsJ4o/9PORFoKU6xPFPZ8tT/Lc
qHixiyZ9NNX4YHd59gZS+2MOgdno1YVP0FgzeJ3jvmTAFZ8SOZFuSPWa4DDVy4VjI9YLfCH9J1rM
UmK7QQbkjBAnLV721KTGJZhsy1wdEMY7RHdDUOOpQhU4DcPrKSFSAOXp42Oaj+9e8NL24874Kzju
Co6/jPR+wnUtpmqHyZ9hF7TD4pak0tTRfNdkEnhy05L4a6ywrM5vrj215eNb5nQhP92p4ohaANUz
uMM7790dV1C2zZvcsmvgWKtit/G+hJeI2mvzxtkYzlaKJNgOuRb4DGeLdTxBoWH5dgWDGRUdHQ6d
uF+1bJfvwUlyn7xW0rViJc6O4agAsXcYsJaRL/8XPkXNMIfkVT6bSI08PZHn0d39D/pwNBZfXTHM
X70zCIfdQybeYISIM6Y8SBZQOfbAImVj10TTditmGkIrmMvdsIWwDOYikYDFzklMp2qfJ7CLmxdM
F9AteVl7AaoiuQSR71xWs4O/POGMxF3GyCL9ErSBTQblrRgzDTuvgusH6JLgaqLrwwbv9UNG+qze
ldoqXHazrFsN0xY9TN38Rfw8UfZHfjB5ciD0UWiqbtNxXQ9icTqijmAVXoOKpeZDkDseFRXznztZ
lgYMVdxEdiOwWM9WP9HcOREomg4daa9ihXneqy/V/N3z1ucX9wstxpNyItrAN2pBxrrI3K4LYGmH
VhrvpLuQANlHR/KuKbzugwpsyQc8xtQ7w37cBWI3LebP+41D6T/IHNoPf5sOVSIX0RYZINAPYCGH
0OckWBkxv1Fo+NCnb/Pnn4zMio0hJVPHzDVnF7EOTj4Bh1pGasHOR8+o77pqbwzpZgeBZIjMaKJj
UqgoHhE+DL05HPwbOR0GNJk1S/qzN5UnGeXO4gD6FS6RyEcbjuLAXUcbxGs6iK4pCRXGmh5/m8Ew
befh7g9GwByCH+b1yVR4Yltw7qE3mCPsfIOtKWwMcxCmMnqJKqnA6Dt8hyoCAPeZPh/L1iq+Sqp4
g/A49Y9TroY+P/j09i6Yy/KO6LslP/IKHhpz06AHuuZdKdwtDbWkulhA5Lk/OXTj0UnbEfSaH0ZU
RsjGrY/toN2J2oolPcELtf9TNjbAcnopHKxcD72ObLsn6LJkeXyjG4UUtooedNqqMsPV8RgOtvIP
woDIKFPlmFLfQ1jjCUI0Uvs3oSFi1aOrMFYffTR5VPmftvdurFzGq6Y6yi2vGtGNt1vHguoNU9zx
bb2Oo5i+bhsnVKz2u/dXGEkWOBL/9d+P8osYCEySH8NeeWWzqmRzVkTzbxRoD6GStbWJT7FPOQPF
m9bcumxnZhBgySBgfq5utP9azEWBZ/+lzfY6FX4mxxLPt0nP/giTOhgX8+7l/mrN/9CMZqpYnZcx
y2hEKkY4dknBIt7oHIAbPtK52DB3Yd1qIaesTF5P0ucLh3eoFlQ3Q722IOPoltJe2xft/nmwoVw3
LEkDK/ZJ7BLtD1B3owzMERLu9ztpOlnCGjIa0Z23I+IiTw0Q7V8KkW92Cbxq8B2FDAI/D3VbGueD
pzOWlSg6tGHyOterZl3y5KY/XODcqP+dXkOEcMT2irTU/gJoAliy5DKCZa8V4IGOCJEhqFdySLIN
0zqzVNm5ldyZPoHogsjwgNCV2XtLLGbOJ0WZXpImZmyclHosNxjc0dscC9lhl5lDY4VDM/0BifpB
SAg+3fUC7bf8BQeJ2Q0YilpDBsoiMTGbjsAVqcj2tPBY2QBbbAMWO1nNi23cpAFvS8sU0wNfiWm/
V0bk3fay4x2hcNtu7hHh8t9Uvmk3F9lfCIY0oltFVlCTjgmJLjDMZvzD//8yClCgRiBXyYbpSoXq
/FZVzgbF+O6KzqL8m4wBlDfNtcllshftZhkv0F+Bo5fMjGRoNgA4ZrpWsfwafJcBtCgpVMASJwEO
u0XtZpPCnfLUGnA3beoIwn0SF6w6z1rNhpxfWBlzPMUvOjVdzAP0l4iBZDLO5OYfquGAvIx9nopg
pBL2cnn0m3BI5c7xIhMCaozjnmCAvKe/foqjYA0YswsR9HrsbIf9cV/DhAbqqlei6VOIzdJdWAe2
+RDAI8BpJPU+W0kMDIhf2eLlGqpBjPJA0c8Qd1REJlTa/2mB7IWyrWRgNK+PFwv4pBXyGRjwtfp/
KzksvpIjQyo9wIWpmMeaveNxaiTHi9O1m/tFdylLKEJAw4LS4Qesce86T0ixNIuSrt4ndHXRXELv
fKtgt/coomKTgEY4GPC9hqSqHMYNjMygJ2Rj734gTEzwaqAPUyXoiM3cvGuqDhs67dN/fWqc/S8t
eSZ89ZUr6oVCMOyn5kWYJukfvLpSOJoCGTl5yXR436OQQmXi4Y+QIkGdBPmuJn2PH0ljriRJVFUx
Vc0HjSddCJ2uH0b04yRGBGoBMrCs6HhAER8gJJ3iHwds8PPjde7gL7mushbpOr5RiCJC1bCQtjNg
Q7kDYK6/Hn17ZNAUjUsnaiDhvfHdSBO5xi55wULpK9b9HN6B0is8adnIS0KvLhQVsr4KqxqhXD53
1osv292PH7fZsp34nPs6dExZjK/RqNv0QJw83DZuhW37OHumaLCKefGlT9hrEGzTgQoA/saKbBsv
XCzlenMfnbrLen9k+u7xgPMO+muewm9LHLcDSgxju0tDr84U5i8qhNsDLlcEqWITSXmqGLZcfLRU
HhGP/ThDXWMxHR9vCV8KFo45sSHa5AehlFsqoh6xVzawpY/El6wMz3mA90lUkbMHJNN5WvFm1nY/
d9lnampXLMU1LdKfq6HPwWMtf6/5/24YTaFlZIXteR0MUn/JH++b+W0KwjnE3C3t8OJFDiTV3A/y
yL7Hg5jMvusugSwiqMKuxm071ZC9bxiohQQiT0KLNDY1v/cZHILTogk6+8Pxx2/kXwfUB2y02Xr2
Xe+xJzLMuUVdbLMF3ppt6nGPqKuQZQ2B/MvSD/z/mMreKpq34BFULQ+Tpy2nY2NFl2bHnJ56YE3/
isZPjkVuN1sd73k3MW4wVA4NCU01GkyjgreflqCZYAF2BTW7pKJmQlMo5PfEPgqVhDMNREt3i8y9
ebVfbXycZS5rCLIWmOW4oXZAnhgO1WyoveGpqKMvqmJRwIiua8QoB5SQ2vVvzPPwAGPYlVthjTke
C0y37/67ZuF9Sy3KiTl726cYBvUbZgvoLgOPeveltDkLuOjV8ZF1dDQ6y1yVR7t8K2TTYCxHUtPg
U25Tg5Ottlzq+7kLdAyOA3TzWvM8XnXC7bkOB+Cl4sjqqrqWxBM83UYF2QwuL1kDYVki0AatcofQ
Bt+lH5tOLuzmVnN8Z9INNVrZ3EBt8/ql7WJ4t7YQxLPpoV/JPtzpGlDufDN9goX2BuzsiEaDaxHy
lx8JAvmrCbqooW45fzA+lr/0lNWFNPrxSNVRBXYMobF80BLrZ4zEAAwCNNYm7iSLIsBwrw4O0RVY
CLmvtU4tD15Ck/AcyWyjn7g/RPwQTpEepFeJ6T5S69b1wES1UCRqyF1rddBgLhXrKRNKD1tkknn+
1RxrX5GNz/xsiLORtElimTprdY1gNYLZEWdUVF97eVPewQ09cHxuPbqMOKz+WJgcWD1/Rr4ZrCgd
qSzjc8xuzMIKdaoj5RcaRfKe5UJOdiy2wh5HqLdGquUXrrXd6dfD4rv160GR6DMkG2hX+8O8DFTs
uuGKnVYGroUscSHcVF/VA3IS0PdeD3q5OTadJDkWhV9UsLZl5ZVPkeZR6JoMP2hU8o1kzzMryCTq
WBJkwoGbddxN5Z5GUjKbtu8W5F/tlq2ziWqOK29VEukOY5LmpbTjEkUZKsZMUP/GXyWgBKCOgRFi
qCy2hmA2DO+fBT0keo5vMc3fSVEUqqsgTOkeKOAVigwk6J8gicb5Gf23n5w+zg3vI6bQDdtSGTWG
UFrqN52dV2aZfqUDb/Gi2hpBHc8ZX0lIpDlXtuowzpAsarwuqv8Kks1t7FfIhVnsFarAeCuW3qpi
DGFuwraUsRRno91CTU9wbHrMs9TGZS6wbkHZwe68MY8EJRiDwB2Aa8Qs2qnUg6HhftWAbZPf+r61
xdCZ/i2iuBGdfbniua+8qlnYE63yn/s9RDqN48VBthu9byEPOo0SxbddmEq4pkcRFZaGEh02eqmA
a4eGONqPbYL5fpZ8uMd5dsp16FBJihXy2pvR/GZgFt4DBIsNZcbWQJX65OslC47aESf8qUz+cjIi
yEQbfPsjqQKLdSLaC5wz7JjLjkVn9rx19/13Ng0++2tT9/Os9NF8Z9zsuc1qmBQGz5/VnqJ1N8Lh
EvOwxczQ5OYZi4xlH/g79n5MioFk3JkU7me3yyWde/t6bvDFHfsLKCvoSnSvuu7taAcvDcOf7mZx
MM2NfP/j8UHyN1jL6qljclxzw11c8cUvQnKVGS4lXCgKnDWiE5jfc/WWqo/eUYg9mT8JTMvghy0l
apIJNkvb/M/QG2fkpivEkWmWcIhxdqP5N8V3Ert3Xtekvm4cBy25NDlWHT3DyKHPcUnW2lpGHiFw
eGcA5a1hBxfOJxuWZ9Thlly8olzxAD6EOxCS9tdZI2xN7jcwVQqwUX5yk1S8PXMObJcKC3Zmjxv0
ItFdks4UxpdAJ7NmSJvy9U2gS+uBCh4Pw0FY0oWRl8XbCGa08i2UUklx14ZlLaCqAYFBUft9PGxX
7gxFQmzue66AyQK1qVRXxsSAUEUVgsN+/yntX15atku+ofDlZwpMqjymAihSP+p5N5C5bZTHa2wS
vG5zWbSW3fH9GKTG9dwnGUAakjf7sDXSxfthHWkC7JMa4TA7P51Yx/T3/wwhTJv9fQBm/BNAn67Y
Ml7KC5nS+yeK6sZNFJ6ktJaAyXJK5FCti2yvGqErV3KCTsUTCb3wGQqKPZVRhshGLE02OLSE87c4
mPz8Y7lzp13pWKeFg6C/0brB1Kzi52yQ3yr6OuayL4liCGsXkqvmkTQTErsGD+lR2JYU6cP63t1T
IYue9/meAKo6i1kIQbBJPtQJj72TuOZcxyuCVDO6FikbnDzuBuVqdRRRpoQb3weoXQg1iiCkovYp
cUlBdG5ajr1s5yU6ilzWkH/l7ncRnKxNPvEV7YlA+jRQ9Rwp/jw6+P7WMX5j+7oUwnvNTh11Nkd5
LOoaaq77mH1YLbezg6oLeL20Dgt92dXwyBtq/NjOqBXPAbD5hfzTAsyWb4wdmrGundqIgyexTKgT
w4krDRbkAwWphf70p0E2VVmqJhs6pzQ9MD11xmcZeRdS+Td4SJVJvXDaOiEy7iPcg6PSEWDeQ0AT
sczT2t9xhaMoh4e9H8L7rY194WNVWXXHE6bogpxfpvOte203B0rqOvq80KX0FECeytKAsJ+NARqe
ohuYK3oBkxlPqfLZdExrgqdcDWTyMurmF+ETbxRqbaULQLtTP1Ir0Q/7hoQi/lYh9Mqm5BDWeLRu
qe/TdqSZb2DAzJXJ+IfDGOZFkQKR2qGCB2t58XdI2Py1fZl6KVBSUs/dc2300ToqOLeXRzSOcCqe
GA6Vb6m+M/33qbeHdfYFmvqGTKPFDjdKGFX/SI7+wPjls06JStHUXqRKnuSuxE1GlARi6lVY9nIt
ri9WCiVbKrC4BPli+qBacfm1oJCDtTLeYj6YWVy4x3+qwM1wB5LB3Ss/3CMXQXyn8E2YlXeFqVP5
Psov3ThA+ifbV/7o34zFPBgPlyLjb6y+mAgK/evF7C26Ouf36dOpIaByeW4IlWJNnh//du88Ta8k
TQSyX+mbJEGGtsLHsc3Q+EuyAm/a6v1JUMv7ny99k7TioEdiquZyVh3p8ECIZT2O4eE4qzBEMQoH
9zC81VziLJJMPWkSGJXXSp0dEWB8w8OlapcFr7RtrT9X3cmJ59eTBH83VytaERiNP8lXe6rCKfvp
kophTRZzWlKmH5fbyxaH+RGOZ+vFK1AmV6pViGpKLfPOnwNxdrxzdEcPDZ4Wi+BPNJtCo0RyMJ+F
6OrXLVmGD8RHpLU6DSJw918KAz9zk163JLOb/6GWZpaRLVgDdLFID75N33uhKy+v0E3F2ax94WO1
eRXtw6IYcXoAzBauzX56+Jd0QDT58pGK5UlFTc8uD/qiYTTXMB7zq3dXSXMmO11Wox562qQWMdnb
kjIxsLw1G0cgkBQB7wPk9+oYeKQF8xLitKtXtpusdIbIJQdjvo8Rlu4mRY5s3Hx0QeBxoDW1X+b+
znQPmMQ4p2sW/COiH9cb6aJ4ihiUiEuzFy1bRr/vQYT64b5HlMrolUlTq0sPXISkWfIo/7gSMcD+
qLSMY65ZN/Anwii3rvpFd6ZfKDchYbi1VVTxLVGVkdR28jojVVpKH0HfkECq8ZpZdnP44Z2qg/3F
FJT/mb+eP/UpCC+7DHFI9/jCG7uJDFOKe/ahCspuS2F3xin13fmqCkpT8ubGIphp/eZhdi1Cjqzv
/yq57gchLaG5q0puT15lEb3TYXdsuXeuKBmWWC+EqxXDzNYgYcxOh/caD4/DPjDoF2ztqY2o+Szb
Xrk1BsaX1MpkIs7QUm1sLkcm7RjCwxCQv30/minCzPU6d/6g/cNVxFqb4bqd/LApdc9sV0NZ3o0v
MoQdTk+Ojfkn0MGvD+GxtlAe3mPNgVYmCAJ+3LA6ORszfwWhGjmRLBwlHW/T+tDPk54j8GrSrtIZ
mWjNZKxPb8S1LxvutqgK4k4EXh0QaQyBFmZpjqT5uQSbeyBjp/ZkWmewG+4awnunqfsmKWEQt/tw
NJ/pr0FfM8IIPfOqk/J4kWAopwwZEZU5U1jYt8xfU6X61POX3rzg+JutJ/GE+3jD2f8UpCkGiVnK
Uh9LCcN+jMwMXnhx5ki78oD80KlunWs1bfmE12ns3GwTlj55JLU0/uAZNu9t3Lm4DmMDFoiv8SCi
Dpn1FDQr5O8N/XMXuHFEPMuuAx8eBEvkPJ60sAtuOOV+q6kPYLztUVwcI4+uGGBz214XzNHVVZm3
NFbQeC/C1tsWckK3ogAYVLDW7G7PfM8de3xjQEKLM5tJlx/nTJALPJz2Z2Njt/EOEXOyXDb0Iqg1
6Xwk3Kpc2iwhFHmcOXJvFqGAdq+bfRMDeEo/gDkMdC7jK9XH3qm36x4t+Dvw05xufEncU96ki7zQ
LQcapQlrdCTxBmOUeyZDEliY2/HShA4cMNGd3UV5wg92up8O0s0BMMRG6TTv68HX0gy1/jBN2Yhw
qEznsenkFGWmzXw/8O7xWtwNdF4ygZHtdwycUqQQgHt76C/qH9QCiomZubKw/y4qH2Csvv6HQP3w
dlJYVHyLRqHbabZgXmWN1ta1YI6aZ3C6pdnsqFVA3gaKlprR6lcaIu9jRfHZwpi/VxYGY0er8vYf
fGb4t1TUA965EWxlZ2BKwh+5LsUgNtgiAa8ntcd+Np5gkunNZVltbvyD+aRYRtzMQR5lCOUK5K14
z+rjDgB7fUbdy+p2JQmeChumNE70JEnFrsyd9k+CXxkLyw+qA65WmoFZB01d56QyvX4Kfv++wHc1
Zs2Qh8Qzr3oCsezVTfHmJZ+F8b/T76GQ59JIJEexZod59bp+GUHr0vgqIihH/ZJNIYY8iPYjKi9+
KHnbqQwOk2GG9ndWjLESvMm28gMUURNdelYaZwh7tGRgGg24Fznwi1QC+2BxF5bM++bhHnt5CBLb
B1vUFcCd8kezxHwG5JLDnBjP/k//O6eoA+fuROO7bP4zMFjE1MPPnOzxAa2A0d+s/fMNzDttkxmO
BHh64BdPLrCIRFCo1V314yTaOqLIGuRLO+s/h44RWooPeH/vnKotlWGyulQO+FK7ESp6iW1mUpap
g6eNcEEcmjA2MYlcL38DUv0xFsE5fSKaSh2A2RQz+N6OERnIMveGc5r7NWbwn9p2ipeFUiZIxQtB
DmZom2FLQwIMwOxxmLLRSckgsiGSdNqsQKFAZe4oTeJBkG+AJpe9HYYJFNCNyK49dJo3l0XNPsBt
pZ3DJusPjf/Fk6nlqU19z+MwppP1+sKuz1MKAt2p44O5PqCwH76ljS1AbDlszvjg/o1iI1H+3qAB
rmkxYHd0Tmt8nK81ZUXdxSKVD7/LEnFVQER0Mf7/dfrP5jhXrHugg+B4h4v0GYDvWKuLevlPVF0X
jfcN0h+Oph1DvbAtEtIhKCIVYZ5Xp7JGzlEAV2x31KNfBZMLkxNopJa9b1kaRdMQzLA3wS1hBVbt
yR4cqTEJuckbDzxv8VIGKYvd6oPLDRyWKKNImpc1y3sZjuO9xkKoIUt2LOxERQr869GIFrWr3B7G
eEQGVawKaqmSKiXj9zL+SnuA8L8pjYl8MCw/StEwGSIZZA9VCtT5Y7psEAicV49INsc1Y3U+eC3A
0tyVTLRZ6GH2folI0yq+EcijaLHg0eOgfzJlS5Y+TpSGSlGRhyzWK0EbM8xY+Bw+d8ZLMt0NQ/h3
7nCTPPnsI6i+yfIcXhZbpZqdM6GT3lp7xt2ogWBkuLWbte4MzBN566SbLWBny/bZQwkSPZVJfXnK
AovzzyqUw7omN1m4iVBWV1pqoCImarqvC7GHQUXvD5b+gRe5mMeogExgceu4JJ0MF+6dVpwouGJ5
xQcz72uYiFfCwXcAJVcG7KTcNsrjGBjXGLSPoGe6APJKaGVUe1iifN9EAWns54Ws6AniygTkpakC
naBlJyqevSElTLTEKM9UESUu5EVIxnySvfgbiaqqFduAoiakNjS07nr5jyJlqo/vcm/QQQ/1cH+J
HrJbMf/dUeSc0qdicgPCrHaGvYCzK7dGhYY3Wy/NDHA68kZ4ij1S9ioTZLjfzjLdTIZyaEromFdj
TXPLatazvQti8jyMTjTn9GV5zszXZ1KDsKP1AGlSg4xNxXP+b5PsRfywJcAY9zwt3oU/rv1P8kgu
yvh9sKNwshac0fsBBiuMoXNAGJ4Hb7tVgfwzCix5e6hfvfldxMdC3ba/d+vJOvwWHlBl1NGF5QfQ
+PPV6trzJzcqMeBwU7IxDFzSjsbLetHUNG6RXrsSHyuaN3vPbRQTPfXKNtX72flib9lbLmauuZkw
LRvUFeRtMPsOPHMJ2nby0tH2gLaOk/lcciEUITWcMqSSMbqyNk8d0UQGI47JSe2Loeo9M6eAjwGD
Ftlrg+kloTp/08AmV8xaFNhJP/fEbgQBrfN4FM4j0iflzjDFQH1vpRqwOw3Rl5UZel5+H/XFeolt
jaNUncx3hGWRyRz64NcAsc2PD8NCBnoNEEN8esQn9icQ4NLLUp3qjBSveua4B7z2wwgEZ2ncpq43
+4yROLZL0/i+SrTW6fWjTfwvBNt4gwSGPfSunB3pNnbFRRMI0l7Kx1nNMnhYzccfiHknqi06EVqZ
6bGBjCt4fvvJDrleN0BdrfPMKAKsOIajO5dTGIfJxWzl13zzN/ci+funjYyol31y7pFd/W6gIv1p
4CuFCE61GPYqzgm2dGp8A8MK6aiMmoP+mHNudIN5pyotvlC0yOmzNn+zCwnaOjCI4jwx4Zq4r3+/
aFxbubMJUcauTY/O4hhlJZemlEInyZct0cW29ag3T448bgL82fE+dKFLv2kcan173u+sLlQ8gruY
qiuW5KuLdIQq1UzRTuXny2GG0GVF8kdjQCvMs8wLXOZIQ+w0N/9p+tJAWrjnrzHwIUkTBeqEATT+
2PMcaumBbg6arpEhUwOybg5Vf11gq2qf03JYCpiDbnM45oIA5DJgP4WVHxmL4XEhEfKIGNQMsW1K
6KwmYY/TTuDgDQVnsDIQS0WUskRGgpsYcLcF0ixZjQzBXoGlmpiiPltRwyPNXW8ZqQEA8IDuEDJ2
aIGRraHAA6I5HKPTYeI0Hry5IuJHSFbvfd0y56yLl+x1qP6sTA+ymmZdvgvlH+B+U29RMZTmDQFv
03JdlcmRdX9U088k1tTHd2UfUiDzP6PBqvET/B2GxX9UKyEs26JQfeyssUld/0YFyeOe/0D/hgKg
8bQoE3XDjxWvnFt4YSt4IJZbrJaC5nBBz/Eq9VXip9fd3jjrgiKhg0fqJSGn6XQVP8wPhdPCOdFq
V15vE2xwHYZHXkp6cwsYuEhxEEq/XDbjOsoqc0+JZ+cLnlbHeorGk0QGR+9IOucGrb7R4iSIhJaK
3M9VtORgTa1K+hwCURiGYXfwmbWRNtaFZ/i/qJCnQKP4bzHlYyC6NWTDjJZuaZXBqtm2K+JLxbzN
o+ifPFTuAm15UHPmiqeAXTQgXBn3SKJTkuRP4HTDU4g0ExQ4ewMhYyYFi3KYpu0aq/RHCwx7eHHk
rSp4Lx3jSMdeh6kHdo4PILHXsPZX0fkCPOe7Kfd/k/7RCT3Xfv84RlqAWqnIeejOq9NFJpXrPEAu
yePFJdQQsgkxuT+B1Hurr1znR3AN+dSqPvWINeFWDOX43ZB3CpUQEBm368DmFZMBTcPPMmXjrHqb
ZGXeINLU34PZUKzaKykeMrmrEAQ8f1zObo9pLFuwTIL7zVVNGwiL6qcrKZ+jQrwIM+CNpiEYvrT/
sQ1pcQLPXOyKgkbo8BwBMZeCXevnuy4MrOSSlWkV0Jyc7LoqDu6MgxXz/3S4eliRYjavVHuQuOw9
bceu8rWYX6wGDdgf0NObmtuYH/paDb28l4IJsK3VvaB1dOdCVD0bCR07auEdiwy4eZ3X8WxtwKXs
0/2zKYKIEnq8eZSVfwpapN+tS4B7Qy1DOdfkPwRFTKOfLXj7Y/SNGWS21uWeqdR/nSSVHEq2bH6S
mzZPb2j0Kfgiyt9Vt/R7I+CSYo4QIr4UKVlOHaoDjK+4uRXKuAz0RtuGCGB9UwtaWTFZ0M7XNOFJ
cOWVbaupda6DmvFtdTegRr+OtZDIu0yqL8xGz1FHEOiWYcPxgeI/5EoClcPPdcn5/D5GYYvlshCk
mDdSE6kzqP/3eYB4WdYuhLMl55SJp6L6EI8J9mSraezrpe7risKyAi9PJwpjIUwJ7DBVJjADBeIr
siHNvh9izJHlvRB37+m+eWPlc7qmFNmwYHXdRFflCohYfGNR4Dlf7vxTdDUlQciX+7KxRABUKX38
5zREunwXxNkLuGwyrZrzuAJbP8C0/1tAla0LNHKke0wzkXVxa/USAzkR/yEFYQHwT0ki6p9p+UjI
5un/eG7jwGS2BlslPA1eMTuE64K4q6LAmgkCGGBdkZkQjeI6nF46sFleNrf0zIpHu/+pkJbc9xy2
ozinavwH1jd1aiRtQyNmAc1KJnnEVqfQ2Xrn2JYZOda1wjfSrkZatWINohvogB3VevT53SKRkpc7
FZsNWi+GDAmRp+O83/InG30OvG/DcQLucBgotK7pdLV2tP1wqLTkAZIEEjWAxPSW8VRJotFPCtMg
/N1sRglq0MWhTWkQEm/SkE3t/LHPvI7TrLAfVFqF2ylf6hEe6/Gm1V2/i9T/sSwcaB6MgWuIfC26
XFUSRoopsYyXUFw141ytGt0cU5VMYga8pK/xf5KmHbM4b5Ba3PUGQ1wF0AtPbOjy9jtkzWPqrZr3
wjC2uixmTydcUXWi4J0mhhIBsOQ4S2EnerRmpsDxK8PDoCLEhkl9dMVbEcxRoDh/CZA6e4iZig7u
RF9/E66N7bqEkCwPU57WK1W1v0OQWCoQcr/GX5/Q1X6g0Wt8kYmkCEmFolA7TFjSNtQOG1LJdcFT
kOhsuHCWqtg5GVT9c4cpYxabcSPsOJlst5wEiUsyJSK2fgRBfxzDEFj02GUCJ9ALuKtlRG7Skywv
aO6j8FCK/BgSaxeZYS9fF2NX9w7YUx7bU1OX5zp4mh4LRG2qzvVzSG4vT+YTP7u/hxBYFiPINeFm
pVXB7scF8qae9aCSWAf5I81VmWwdZLuLUEf8ZIZoBBE/l899HyZd2lJti7chZI/E3T3iNdfDJJB5
pAz0+6i00Jz5F6g5lBa+iiQbTemzUFBxYjAgYio9biPamMYkc5SySuK0xu1QLFr/NNgkgCOn1TJK
2b9yTH6B8zYNc3MpghCd0gDh8nmRVvhhG1jlNBkhuvnlGKsl+0QIIPamDZ7RkYtkrDu2JouwN0ax
QEAyiW+xkm8jMZ2Q+6Q1sLGkZTf7wELFOyQ9YHuAnzepVtX5vct0iKEj+STG4jN6JnUgrXDU2LWH
S7ZvEKAHe6uQfaFkzI+TCJjoIJ4L5TCmVm5iIPSU2yQvc9kuEpVJCw/w4M7ONFl/oHE8JRh9SJOw
ajrSGZOnREUuIwKCi4GF3JNaBfMxgzDOfvBUorc6kfaKY6JPdY/Svp/wLuNhvT5RUSzik807YYdt
CaIIYfC9wxzHuC5mjG02mDvpb6lalnXIiziOVXJ0TNTfnWj+8WPBoILGf7ahMd41vAXbfhNLazTT
S8lIDqgzJGM1Jw9GNHxTVL5w5jsB9Tj4Uoo8KNz9mw+zhkCwmTDElVSsop2gVPTl1agGhGOK571t
6Iv5v4XLPTEN24g+zNwfJ3dB4FjPjrHcDJARkRISMi0aj4/WUVUwt/I58VQ0Rzw/RBMZimBpC7xo
r7ozzvXhmTH1l2grKigBQOGSkDsBCo5x+1Ve3EsSHHj1TUvo55v15WbqfHYSJIREwcOOkGDFJPYL
R1gSCAXFz5SU/F7h+oQTXiHLMRPmzBe4UA9reRjPCtvgm3DCcstYZ2aB/bGb28q8F2Zo37fRRN+8
65Tnlr/bM51PwhK0vtnT5r3lS10COkcxXkHeMa8nHS9aktL8QZ3CA0cRWXY5edVOdFKJkHrd2HTq
w2WzeBypKNuZEMFMAnnMrLGDJy3prlVaaMtEeYU0zKIqEN4Rh+lCD4XIepZSo5OOOzTuZWD3rTum
ng10HstruoWtkI0qQJbLmMCbz0lgnzboiPJl7vzhsfDzsaUwCuqxeQVfK1M2hCppWWAh3q7ZarMM
EzaEA4N1M3oGGuKLmDUoZhh4hHNnwLtIIn18EM7tO+VY8Ni58TRmvZKM6HN+jFXlObhCT0ZRxkEd
rPdNyUHxXr6omlN7lbVHBaVexdybhglPj/zIiC36OYi8Vo4ZdAPjqU/WkNB/RK4vvS4g9Tj1PACM
6knIdUSK7Gvy3hHM3X8m4bjRY3QdlPKIiipniMK5aYLwZ9zxpWhaFpNFuhq0T1+GvXDiM+kZR6vf
1P2/vh82yZgih3qzezfg1vQE4y0RH+leF/Uc5Q/uQuHFCPuHzDIDP8+bOBER+V6Lwy+WxIAMUC5H
zQRwmnjCA3RaVqsPK3d+abQ8yl2tPlTcbnHo7hSOg25ktMRwOnIOueoDE6kIShIV3Wdi9ZMCmYpA
CGf7JlHe4MLuC0FH2f7cq3Vjp9DliOHM25d3H8YbjHPe28ox8KYFxG+57s0OosJsSqKcQ2GL6wUA
nWrM36My3y1rioE5FiXnOou4mUcmD84Vr4uf7OiymZCGPVicOGntt2nVroSztMt++uk2OCc2/982
FnMLAJSsBII3VUjgtpVR3pxYa3n29iNWxFTi6xvDF7LCWDEF7qMunWfyD/LamUFpkT3Y0ymnEELq
KUsG9ubRhwomlq9Q70CT7f9Zrax3C/a7M/31YUNzq4+OrkwYHEMbVN6I+3TjOIClp3WTLS3l9Lnx
eSGnLYsWvgIzW6PGeBVT50EYtwts7dNNhDTQKX8bHEEHU6O7bzrglXHFW2f+eXn1vVWHu46cjOAH
Nunk5iFHtN4KxTgRgsSLSMcw4edJex1LebTHzcgdnjclll1wIeafYcjzXWmuEbSbeqnk0BLdSOR/
KA9AGpSfxSXQCaH8D4wLOH+CCGpnjBh+uRQpMLz1IaD0AaRV4NUxyAFree7Ic9Vkzllp6If+Eyi1
y82f7wEuJqICiaW3iqT/YFzwS4PSn5UoUd3ODh4spJ88Z5GFKSeZgoZUhxCkFHWsGszy/0MtdEVH
gBYRYCwrcmFbICCMUd4FN1fXX18P8Q130Q7Hd3QALWGIuklvjL7o4VQDzkpLNVl9ALR9HPRric4P
pqh4TVAgTKOLMBipZRGa/oQTn1SRaxiLpxXMJRa5nkmkBIY+mVKgmwVkPJ+I+wU9c8GR2Rf19A3L
jKt6ah4t18xH1wewNtnAkaermu+8UmCGU3v7SCKqnDCZTe+HNWWRnhE7kO3gn+PeRQN3dUdCl1G4
7U72whM6DdxSOWqd9wpjtU2iX8ybHHo0ZYCyuHIFv+2TnC1/+GsHW9TGGLAJlW42a8OUAzrvDX9z
hDNLY/GXiA4ia50p914622OplgkIcf5fybdvLqS26m9L6nnHKPr3c+NWourAJUUv0KXp0iCNUuEZ
K1Eo7/PvnVCwriRqvFot53VWYQSEB6VajyLCv45jXlRFQ+2qUjOp18fxWhovlOGzopozHKC0BiIt
3sa3g4QQXbt+h20G2qU/iRFIlpb7IoLxAk2zcOPCsm1qkOsZstJGebu9AI3QrnRndHGGk4jhpr7t
d8l+nKzL/eZ7g1JCwqqncBSXfZN5wQoP57bAsqkF/1dFern3ujGNfXGgXrAyvOmrbRJnzIQGtou4
PkAqgjFqYrgtH8PDVhx6Ajw2EY36ALkiblkvxnENDEsEZS3F1yuCuQQ4ZQ8unfV9olxwVnUiWBAH
4cmjFP6D2QbqMXwUa0VN+Gs1UA3XNnyz0kezpDpwfLMgNWaKZ3IGWYZl36dDCgl/fAbqmccAW4o1
AS0kOtJDxxLJJGgIrHYf5hd72Zok1ze89B2MY8oipo2ijcImU7sUfQDkt+3S9Dac95OEvQ97E5Pm
9q8x3VHks9/M4Lw0EXAdNc/ZXNXLjYmhJGtSVZPci3YMYK70HJH5kV0ryr87HEI7nUtV7tctaT2n
8kF3Mv7J0460S3qEDH35GKdyF0GPjNb2cSkZswWl9KOutGvL0z3NxrJv/+TdJ4DJ0Quy1wgTpMpW
rDAZhzwvlTeSMk0/A7H4+GxKNXtFK/IM/MSrHcKcAx6FEMZRrdvKnkcrrvXjN+hmdUC00s1+otNk
YKhZ9Ktg1trgxyUkmLoJ+L+726oB1qOUQ1VVLWqbwoC9NNAmjbPFqVx/t55bdbq1zXbJ4tEY8mNX
evwo/lEahLVKm4yLz1+p6/JvlaVF60qZep4H/sZfFOAZUIEtkgl1Ut69itp9Soo7ou5QuAHOSGlk
82q8ixW/MRyhbQeZpKRTHqGdTbiDfQ+cWwzC7AmmwI38rnjqUqGHHS6aqQtazmblBqHxQE+8u11Q
7PEbsebHhar2cjMxDBq6c38EMqfWeYUryKRKFfnIfoN5UJgumjk9/RH55BguuZfK1st+EqOeFaoo
n2sMuqqwLZrQgV8khhODa+yX8fNYorGwf9yaxTgt3wpFvGBoLANtNtzp1RB/LdIP90QWr9V8QBVe
mPIT8E709mG36e0qqx1TaIwR8R4xsrgPTDBLdUBgMXL00UPVwVdAsubhTRjyZnEdxIF4uySTLM8i
4tUN11cqrlIyf6fyM+f7Ipp/vay6XsvzwvcXDtw9ZPRkrhlcTp+fwHW8wm8YV7frfapJ68rcqt0W
d8UVKBNVT8U6UQXiVjpOYFnrW4pDd3cGVe/HChuAdo1oeauIO1uKLpq4oGyh8Mz0TPlmFRvug4Eo
lfWXaSFzUXJ/wPylU3Urlg+L2jcb1Hp2jFo4JEP9eq/2aFJsNCk1cWxKpSkOWiijR5SFz3RjVJOI
bbbhnfIzkZtARVyXI92bOkisXPVomNOz/kqF2HRB7utbRWG8ISqQmWAmaB1xzMCn+azvd5QwY2D8
AdZRheWAwR2o51iXPL4xWpmZ+mICcTRFAqPJSsOnvHkc8UXezI/rFui9Zo+kXRlKag2yRpXumFsB
SSjS55ZVOrHSbEgW5ciExdeQgl5oW0nsJjV7hSIAQoFdA+xL0+38Rg3qtWf8spriEkoyqg4zXdIX
90/yt+mlBA17KpCVGPkD/7YqofR3U/VvUXIQWWWwzUcBreJb/5q1xLzkQq0Oaf0I7/uD89ScOqKo
AWobnXigZkcXTj7I0Hf9qUHeUBjFlUf/u8kl+vC7rD1rpndktai6aMbSWFufrrbepjoau6JAKVsI
oy0aWNACnpJ9bgui7Cxk5rQKNQoy59gRxfMyLzANVY+azTa85Wi+Qe5Wy1UA+kVry3T5jdpnQLAW
MPNMhKeNScpwWGmxiAabOeGHQrsWdhrWRvTozryPEqYjIQx2XsV9CXTi0QkFHLA4730tRmt8mVWS
YkunEE4hfl3kIJmvcoGzo+Y+xodY6cZizZwWyCyhOcgRImGuMVsmUZEMUtIntxWV6i5LyDLmb5FU
y1yJ4ysqCSF3G/5P0/q6xoHkF8Yb4kE7Mqe83fkvhesTEoOEfX9WtB7mYlzoZyepmqJQxm/MmREl
B4SKZYYclWeNjVitSqC2FaFaG6ZkznMtVSBrEK/KFjkpmetZG8vrLafJUFc/UQaNKASSRz/G8KBj
59rKN1+6mxbA1oxcym4vqLYHeBvRU18IMlNGIfWn2OUo9HmaTTCB1sPJVjH42YerhRiKadL8itPB
okkG6KaQ2BwnlkOo/dZrne75LllG+ggPjP7BAlCd+pzmjRoUfSVlCKDpNyPq0T38ptuFLKjP4bGs
4X3bcFtFGJZweyh7SZNM+r50vPj5ePSmINPRvAYATDluhqt4X4diBGDIffFMQgPcGN1o5SdxRvSP
Z9+ZDU7gAnnUgtJsS3dDaPYKqTdq0FLASYGGV7r0i8WnQR+97YJY2sxhmwnVoW/gKc+rwBC9lZNP
6wqRMBi2MTVxbYWiESYxELrLgW73pYfqHINQiwtIoXlYHy55xyg0kFn5NJj0bzbQ/cjqk4uaAOaL
X71QZq0aC8764T0GHTd0h9yINhee8IruXWXr/+rr1H0bWWwdS8EQtlJvLKqBj9Zl1Lw5oe607x+U
kOxj9xiXZ8TtDdpDm83QIKPwH/FcHuqVuTznkPiDiW3P/i0k5F2H1162cfxz2M5+K39qeSux997+
hU+UqHiKQrrPv2skHXhZoZEsNoh8XXbzzUe87Q4edTE4JUsmZnkru290fsxen9OGMLARVkUMNjql
jB1bDHkAM9CEABV0+LhlOk7b71o7aYpZwBwbwyytxooeL3NZhecfi02buUUs94KW+cUah7yi/nAf
rWDtplx4JUa0kmHkXozjMC5Nac9vqLreVn7JepNGhpX2HnmcJFCUFa67TJgY4kXSQyG77LkOUQ7l
xVYy6FpbKvJcKlLBbmczjnwP+kDRkfwfei61YJAIW2ySEpdXwQGD9bsitpgBpp8YB0b97/dqXQfc
In1hnwHQziEv5+Lor8Ok5vG/JO5aZzxetWLiUkHyWBMCa+QIDD/YtFFVn+LteaEOgaQJrMJAolq8
uBbteU521H5jgdqkFblr6fZx79rRR4t1ZaSt3nYXqc2iUWMhEWoJCMpwXmwXbK7g7FnyVv0Hsk1x
W9OZftnHrXa5pmRqZZHRkNR8af5t5mLfK4bSVu0WLp6FfBjyAE6KZjFrw5i1SLRWmziiSuhA9kv6
OSgdry+OGHKeOzUi6fNxSLY3oxh9LG9lxx9tIVgTyW2omuqGAtgarmafx4J5QFeTd2JDINrTeAXA
FcMqjIF3kdvCjvwx2A9ZCUcSr5IoWH1ZyueyLHlrQufbTGenXsUJvv5WctxyZPrgZBSdGIcaiVIX
Nt9oUcMPaVd0CpYK7Q6irFYIvWyZ2KVDn00luuHAlOroWpf0k5IcnHJQ9eE8O5suHAJuLU1qMoLu
VYONbzhq0tefvJDnKJDlk0EB/G9E6bxdeXZ1hozPgKvc48nA9qi9iezCKwFheWGkgDrizAN/83ll
hK+nanPqn5eGUNMDuXXuQNpw2mAuy6RP66tIyZqa0747CmOQhUEZkOh7mvQpL7f6Zup6SavrrPf1
TTh13gKbUGcnUSbDO/jj1siRJSYJ5zbqaQqvZHkSLPO/oCtqoOnlhjlYm8+PT64BV9SBOLbcDed1
ZCnyNIZF4QdC6wu+I2oYLKwjj+VKMbIvniRPuO4TjOQJ1NQXk//0KpAjk6yG/QIFzsyzNRVCxJK0
A+ycyIeg4F/weIcNSDhwyqHv7doZf4EZWJ39UnSvRicY8WL84+D+bJf3qnRjYAfgAfxgDywCNLpe
bGpCFQutkelCsLZ/uKOHiLwwPR3yGLWb2Ts+AKVkIkxczndfJujughhRWKZZ0bScWzqTRzahr3lP
lu1WRbC7UkvLjw5az1ExTl398GoTt7R2nI4azQ1tMtefkHPxaGxSYTVc2qnZDgBZkOC60+b/T9pa
O9BNnmo6HRB6CUEl0QOhu1Y+Iu6ffoaOdFSayH9E7GMv+/uHb9rDP4vUoznfLbBQ2x5FKmF7KA9L
ZP8wLAG+sGI+vsipyefC0/WqdAhUyD7hluo/jRlqQXFSE4rE9GKakJcdhT8inpsu93Ewe4BmmIJP
hfLNE2EEWN0UWprccVg1IjVZwX0j8uPRQaJzjwxF92xZVEtMf1eZ/MbJhu+oL7khKmus7VGRICJs
3VjKeSYfGtgBjGxIcNbBr1+8kX4nstPVk1qF+KoOxl2tdKMcZud7X+DcePL9qyWe8C8MdYTCVudp
4sJa7BZybt5imL1+iD2vn7KZxlot5998UfezWpIWkY/VyCa1VuIjys74Vh0SgXeOf9Qym2D+uQqm
B+H3mwXNmE2IWOUP6HZUneKfcKTY580vx/Fq6gvq6fLJB1fL96FH3hAaOptilCx2Y0KQjt1xqJ7n
mdkGWnJr7hLcJTUxXFCrvF4uI8i+Da0SKl10K3BUvHDoBgdENm+cM3wagq1YdfQHV7pfQ7awn9Qe
mWVSJVWuAVLY/v5seG5xKMNJ63t7pA/o7Y42UVfmvG6eoQtKX4bHUOTYbysK6JmDITl7ZTG3cn+g
ASUOF6OK37OQ0xqBh7vMx4tV/PGiKkgUjfDRp2ij6Czs1UfxL2qZI/rvKbNpxXYQ2Jmx2cAfq8yl
EFJB4CQvyrlZxpMXg7W7bQ7QlNxj2eEcw+T+FYsNnlyN8JT2Dn9Re2o9FuO2hdZiuAIGNj9OqjtN
pOFcunDDyjXsfns4vNYACRcnoBMj+nBG1wltV7d9riFIptK9nMbUCIeLDfxZ9Ls9JL0ZeIpnCpFr
iSQNZfOAA41cjvLKLmAyL7RMYGLXV/SkDYLW9AQfUE9J2qcW1L0GSjZEo0tg09g9mAVApILIrhFa
dChgpY8BuQbGS0lVleuAA2vTk/qKaiMTce22C1QAZ/ikHUuyHn+0NXT+eMi5nb7Uv0Ov98uu9tV6
GP8W43SaHfM9nGcUWdgWEy0E55KiH7q1V/wwDIIBrKfzhLWAiHtsKv8aZfHQsPNq7humF5DcVePs
hjHeqrRB95nOpJftH4vMEy1lWwtrhCvLOirxZ61XgxKX0wFJo6LbJekHgWmxYu+wwcFmIDagpRPZ
fFxBcffo6mxtgw87cEayX7L7I9nuGsk0bvyHLqcEBXKG47zZw1vpOxe/urNwaMVHZn4UzLZKV57m
Ir3hROjodplzKxvuRVj4SvVXwnGBdGZO1sp1e4ToBuDaZmLWJ6HSvqKHPyHXNnQeBE8B2xnWIhkc
WrVUzd8jWMECsJkpS6gDM1Yyiz6fHg8fytnC0UUY8iTagWlsCd5wbOa477JfGrEk5N8KVysmU4VJ
nGaAK2qTj3D+FojSEJacWyObuvlYkwe4D9OxSVSMtuTloaWX1hiXl89IGxhFvszB9coiXrjggoqi
Hz00MGmjneT21+J9soVJ2sL2TnJQ4iPM6W2r7MXUnyAAKXt4UCL5fBNhjGo7y+gtqdnS3+S0cMyu
/YrwaURlrUWYxpdjJRiYz2OQqDmcTn3AAISM9naBy5Ti/nPGdkNN3pOQk+TTs0uOs8HH3KqYMHUe
i9BSOY6HPqQbZO4/nSb4wACa1zbUQvvDg9HfBTKGNhI83xa0q9febdsxr1VW8tbOurtXvUQ/Jv/E
wyoeiRam9M3nb/9Bb4/nOSLvVbn5ajFko8Jj4V92KkgVpKO+OxU620LbxVIcbu/ZM3HQVru7qjn6
jPvMZG4mTmWf0WZvvn3uhXZv4fcC8n1Ci1wSkVxUx+Xuzl9CO9ahOfzSGkZpTY1QsCwvjv0UtTnh
nXEtFla+JSQkZo6ZoeRS0fYF803GLClDa3yhI03HSwnY+l3g+aFqa9as2SEBjtLOWtG3lYtECCiy
jcrLVtDc8Yj+Dzd5FhiIrLXwn3kFIEcALn6MjF/8JUzTi2taIjHlB+5hwxCZrFAdog9zhHr1r4gZ
FKOzfTMS/Urftm7d2EWHoC0QHY6CcWoUgH8CtSXlVXGc12H9YAkoeryDLkGRSXunpF5KTap54/V2
Tsd33IoVW4Rn9HBRsggjoU+AspXhFyGlkYxhd9oACzws3WSmYse9/cd12o2YsDlFfBSSyWUtGWMV
RwFESq31pzK8aErmqYnzNhnpyAvKrFA+DbDt25rsDLU4ew7wuZE+GDdDWaCsJgASolqbOzyz3KXq
9FvaodIGRQAAjXPRmBWGCvGtEpU/gcAfFkq0WygFmbA7wlMP26gV5YQ7KkUzJCD8mwBEUKrICXzW
UDM80B2tcqLa41qZ5ZVqBB5A5k2S1fGZUJv0+5Y+iIdaY3zSn8BtHjzvNCUr8NH2xJRHXic/S9SQ
bmEhJhuFpiT9NlxN2rrx45eWVq72F7fzCmuFk9TI81M29SOmF1RfPR6eGPOEq2Uiul7c9WIsw8+l
pvd0i9sZUmv8nm35u/nSv+jMh9mSQkLsYua7zrzyjf/UpxPCHqn36HhB5nqw5HXyEbS+lZbUAyzZ
IiKJYGYF9N+F0NM9fVTFbuNRn8mfvP4rtkLPanR8Ag0fcUpP4ec/dtRUhD6YXyMa1IuPuk42eOom
zRahCROkVDbwWkmLbO1dG2LxWdn/NG8gUr9XYv1s4VikVQ0iz3HSilKhIW8MX5EhtYFPFH/p5+lp
7uJe/uUf75bkOylBl4fULbXBlJ5x1f6kWY2KPaN3mBjAqjlsFDJlaqKdDoshJipzc4+qcNm0Pha1
xIr5rEdnwbHoLtRcfne+Dry1KP3sNv44bHZn+vMhw+oJqO+5F4lqMjpr9T5y/fkVA4/66wQqxabO
fhjVZ7gGgEAec6R698MfVWnYMPTNoOmy+Hm1ryXF1SVc0qDVbfkW+8gjY4OmxnRX+jt72ecpdSvn
ejxnEKdXPQ0lUrdZZdaNS25EgoOoHUNubtgTSoFq2N8Db1wJqZG4q3gE+1dKcl2yQJbUCovE7h1I
YMgQG6kJ86qtNskFKUENnu50+d15bQzg+xNG8DjSFRc9pQDcyVYbmE1Q4UCNXcAGaJQ5PilEEVoN
zDe2MqA6OxLDeQ2Mhz/PQeqknGckOfETiJVdQv6LKejRUIno8VsrlLOo/aX57MyHQl6iwyp+F7pm
7YN1OnAxk6bBOS2+HRbu+hIbhn/ONj+MfVksHH5yBSy/+VBffrR6e+yQPFdV863XiXaQ9w59DPDG
BInrF6QxxcoB2HW/xkuZExnm/XoGlgCv709sLLz2+q83KYRSgJLg/vDhHj5lX5q0o3+u7aTbodK7
ImDTYzaaQVbQXguWqWzsCIxwLTH45TMrRu9LkE8Rg6aHZfmP/QOg4e2pBfL58LHASAFNrPiE/lU7
YYvzl+kx1InKPAnUG+7WlwMjrwULs0f0svQWkuLQ6EJ9rE5G/9In6qnH0N8+HTZDuExUH0py4E9D
JT79OSOQZoihpCaZNK0PDSrRyTBO7MzCSnpTVjcjHMDIsUAa//tgQiHew1VeX4Iggv+WZ87KCJgT
VigMEhrzuFU9BUh4GpoSsCsPqbfvh8Oq7B3sq4CSny5ceKtMtfJpTEJn2kiUp7R7HMqjz6YyKctZ
o02UrRUNMJ4qc+nngb61V5D93WrhbvvFEKLeAhi3kSoGF1En6Isp85EyQT8zUffMC8rego+3QQkX
QhKSctIpNAJ2ERsYu1UGd/WVVPFJz/u8ACsNKddlouAP02R2T7bBX9rh3LmohC/pZbvukSERBPVc
Vt9Avl6wOGgOiFjLmYj1P48rF4p+s1OCW+/+s99VrQy/6BK9KJFyqpzR/cVIqK+00+2BJJYmKfCB
F3s0bBxLTatWbYwDq0K/EEQnguErw8WD/1V89MSYw/7ldSENS9/+GmWKNFqKm9BED7JCWfTWge54
kBnmOagKqNIR/KpBp5MHqAQuPKsyGU7xccG56nSpLQ/qqnwM0nsxGhEdQOXtzA1qv73S7lOyOFjk
GIP3+icN/gEv1yzqV8Sbc5B2xv4ZHSujjiYRiFN1kWnEWqvmzEKns5bN1QHa9s305N0P/oPBvh5E
bMP1UhqJexoORvI5KQhWPgkVpeFTSMf8b40tX8VXGMRpi8qi4X8UTOkmyxrqTRlwBavZBX83gM2C
paoxWjMv3d9MKaz9R6mOn1yQKQBo1O4JT31uV2gncfpBMmjHLxcws9p9uoxqqErp+ts04G2ho0u5
AuqzQqn2cx19phBkO/4BePGzR5V6YIaElb5Gl9T+chGAzCK/TeoTUp+jScb4oF/VHsJBKTK4pinM
lsw2SV+KCfgLGbpqZ3UO7Lli89edXsCuLR5lSuUUXVCDl28G5D3GdVxhjBNZq83K4O7U2tsd7TuC
SRsrPBUx1UFo0Bp/uZRfoQnDTLCw7OudntipFHI+yaARI37cYaIEF4C3j/iffvBT3mmH/GqRl+je
imn8n2GRL5rUIS4SyHPDEZU+ep5lQVOJF7r7Na6iKzX4ubFIXJf1HWbV2UebGmgXLkN90nVYXzIj
w0BfsnyC4bzNjIOMmXAicFlyMquRfMxZMbm+kT0cgyO4RE6csvDNE4AWTUmtPaCVSX4NxSlplRPK
oGEUK1Q+/4nqMmKesRZsQ8dqBB4tR0XRF8Ogl6hhF4XNzlBrPEKbyDjJReS63xWaOs6ANvLGK3mj
6n17E2re7xRE9Rh0vUhymKA3r8yEfPBw8ItC7/Z/9srArWnAnmq4W0pRgybbcMh0WDVuk+oabtrH
Bgwng7E2smVZS9UYwmp11mDenTqQjrLumjx4TTPBhlCkLvEISN/z0wBimGwCYjtQztXa218iW/2A
nxmNJQUZTgaaP6sd8sFlS0BclvlkQobBcMzrfVaC/O/Dhdp1M76BWJWzz9yFAQLOwDrukgFx03XL
gPio+gSeUOaiBmzTDglyuzA5cwi6vaVg5YG8TlCb3WEd7hKFxPst3H2HHsgv9/5boVDf9RUYWYBP
c7SFhjxLas6HrBG+GXsv6NVWwIQNgU7Hi0MBgCJMeytEcNRfFkwmo/FMNefIgqFqbTKJNJgarUAl
zLljVZDO2usmKhWRx4W4xNyUNIPnGcI3dj4EuMpCtTG7TpSx9gkzzh4bjN2pkytRQyo4PwZ3cPu7
76k6t06adGv521dKqx+p5No+4ABtOhLFh/RvNBOr3G7MWKGwM9eVkPO3viR8l72r2/tMPFgh2i90
a9ZGcFpxM/iNy3hMyVFSEoGsxoGnAcU/B149Py+9bLuAdh1j5L2Q66TPhqcHJ3VkeclJWHbE/wEv
0f//JDdoYA2Cihkqxmxx+X7iZCraUZjnxHF/3oxKWB/3zdaWxXdy7AoWT5qXpHJzrUFTiipRKalY
1kdNdYYmGHm4Z5RX+8kwimE2n7tzeKjmAc6wUAdIfdy18jrIIpWoAq3shthMmU9J4LLTZ44Y4+28
bMM5rb0xafIibrYQBZjIuOmJ40OIM20qXZlQslXZZbBAJ532G3XZq9hBn7bgODuwMInVv+2Bje71
wi2zimMdkGYyo4ag/qTj6hRfvOX+AabINDUpd3V6GiCVUYTX8xhLf05fUESYVaYuTw4xOViTfUIy
9Fx3WopXmpYHP1lAe/PbbS24dHAudDZHZHoW5beCnsqpATChwh22Cq2CSNHgbSZHBj6EHH9id/Pp
hYeHDVKU2SqR32ixqqXu+soS/Vi+Tj/JO+68PNUA2MM0qWAtsvIZWrXzSiJmysBcvXNGqEuOuUku
+70EeUwLAylG/K+NTzE0D8pJWoiZyhY/XX8Bia0QtvNRMDMKKi3RX7ge/jiGZGDzFVIFnbmZyc5I
dTl7Egmga2yLHOVuOpexiyFR1vZRViQ8FW8auPlGnTkFrPNCV06PVrl16LaAz7AH4XoXji6ELDQb
FkOmhdf1RKZ2kWce9jQVv4U8YWvRwPU5pqV6gZeOEYki/sXTRO6LuJIWzeUwYCF6gdFFXK63mNLU
DJTpK4SFVDkEaZAMCDzwWRUisiqLavzCelB2KP7qGV6wL4ImxlGJniVpE2x+gq69BBl71GBz9kZB
4mMQYZsuhycrp/QTA83sqndfj5aB0X1tsXnZlgaBvZey2BRgwOCA63T/EkImyo5qVqxrGaWuk3XA
07fHd8mvUhYRP+Hbj5rG7lUwIpRb7fT1hUvnAP4bYLEurGrD7jBJ452gp2rWUFlzB8ltnqBLT4jM
/nxntRqakCzd81UND80XQvwiN6v74aEUP2/FJCld/+lw0PLq4t81g6DdI6lSUkoK5Q2drwspr4oH
DsfLWt1yKxQzp58Vjq5VhslcnRTH7r3RdLyueA+Pk9eSsITIHVtmC5uHzlx3vv4zzKjwLiQiEp5f
YvJkyGVLj5k7VRvYYLwG5JwtDMFSKMCWFoT2x8fGcLmTiKq0HmyXwMsJ435dPPmuVrjaomqnGuBs
3uyYi3CODUdD8BmTPk3wSVQahTfEVIsSVIPMLI3cBkiTkOzNApI5lOkiFnXfV3ZmlYg+5Khyd133
I9n7P1vBUj8KKyYsiKFsGjXS1ayLNQW+JhRdDkx2TKCTSoGFJlb4xGqgiOkXFYpGpxxQXrvwDpiJ
BAloSIP7gf24wSYUOM84q+SRNQR2kMSKfu4L1fusvwnEDzZDLBfIqEu/YkiCrqRcUrVnbpP7PtQv
i59ECJlITh4pr0/XDccMFt7g3Zw+BEnAzcb7lR8kidOx9MIK+VOT+u4JATacJCkUtlEXZQj2DrLq
rIHUpQtOeCDdfm/dCGQuM6IcocKKO8CliWrvOr766f0P9Fp0qHP67pP5HgNcKOkxAY83cEKEMy0G
LYauTAMRfRqOW34xjPgFsxo34lEEzkY2CMfnpUJ3Xrl5BNLIbhV8JFna7+lJrptoxnQVDR9IXTlQ
iQKur30ckI3+bwCO5/cwjU762Sykd63Ae3iiSCQGtX6Q/DFctU2tlRYTaIKM711Bm2rSsUZWzfKU
YY5j76XZjhUjjaB6wKGocPxFTnRFonVUIc6n7ZC5sZfylOp1LOb15gUy+qYfYErK8oy3i/xhNF/h
mBP3FM6TlLxxc1qbCI2bXefgqZQU9Y7y2xsJo/9BCosXbbCk1RV8IulvJOlM+KRrvfZm4KAbyj7M
uOPpH+RPv6WwIKCZGZCmGtJWpfixAGvY95dyzx+Ixkk1FUbqnlqAQIP/HyqDh4C+dj7G77+5OGaf
Er2M/QMgHStiGflpBokCd/BdRnURCeGUeN9KWcSuq/UJT8YyBzC13Z/mXTdekrEBKyMeCsZp6Cf0
zGDUXoGJ0FN4wG9diPPFmvCA3EZHGY40Qy+I+Ql7MzxasRe+RefDmu0F+WbuMZuPAR4pFLIBGQPI
hO4jOLlXXqc5O1DxgK0A4kWjoO8qeCJVisZdZnwvM+CNhEQeGZt2ybHlthuRYbLOhA9HDCCyfR2y
p0DA70BivCN36ilDj7EekibI+sL/O1bC7trJ9cwlJLxl7JyD0XRFwrShz7Jr/wQSdl4N+y4geiLh
mUZtk8pqaI9v7D0Et7nuKWqI+9n/5ekO0pboC2UGooWavhrSdPieZSDSeEEBjdWT9s9POYlAh7aN
qP76FKOmAcCMeaanf2HmSucm+UHREP/TSEnvMDNdt2SxeYhlDw5eUAZJmO4/RHlIOC//gTehahbf
OXI0XfkNCuSHuujTYB2oxBEUz6yHZ5JVmLv0DgmfvWfdg8/S4wRr22km3frlmKxrUAliHzBL122a
z/k2ImK8ynKqlt90Ktl7v3UtstDvc6tnhD0/Z4me1ouTrY6ThSADBogjmG/sAoUFCvtdEjVpYbhm
rPq1XEGPiHVx1bbDSRw1p0X8QOawU+bzaRYhw9MYuTNnP6USUrIcsS+/lGbLa6Tix8vaS/ieu2/Z
mJqhx3KlefPHZJbouSE3co54q6ehpg/HNJICWbr6VNAU9+Fzip2WQdLy7fJM1HPSkMRtL+0NxzPC
wSb+5sYWJ/sWG6JK5KK4curRj3cK2AYaWPXqVvzn3f/xlC/3xBnjeq/kVbi9VYRFejEQt4CBYRdr
a0huCJMbXlqWe4KQApM9G0SjIpmKzVtPC2F3+cLKbX7NwB+MpDxH2l5IGML76jtp9Yd3+k06wUy3
NMgmqGTZMN8h9LXOXcl7gKRJtSU4/JKSZVuIViSl+RmBVYMDMzAn5guAQVa0e8gjb9Gf7DXJe/+Z
+tf9OfX11BYGZH74/gJOU/HkfSZXBu10nAVxQmBg3hAf8OnE8guef5kkITRdYFX/uBJb31INZCzn
pTCJEYmkb84TOim/tBT4+pYhuBsysCrqaSHJqNtlEK6pUYLPDVjzbDLnQnT2b1tav9qE7ND/nWGZ
S7bQlZePwt/v/Y5JIzyDz2ZZ0KW0wDjpNMlCSPb1FqhWpNk/hAG9WD0PoO+lL+RfXB5/XUxVYIzT
OM8LPTTbAIWs7dbyGMYWNI5G8PZhONWupySUDWDK9WUgHo2J8i9ReMHC9GdmDAxgeFpkYb+9QB9n
s9oGQ1ZnsHPrUmdUs6aQVi3QT2ILhr+vS9WxiZbOXspqqEPqWiAVlUwixCiEoHwkG6wL/6DTLwsY
U+5EdkNwYhoRSXdDx0SIOohfcR/mqydEaxHq4KdXGcpv/LFx4hcSt1cV6nrkGGR94ZtLldL6Z4Qi
BUTbxBA1wNsyX0kHrnN21Z5iRu/0LbGUuOYUN5lMKFTqKRwMeRBAeRmuAHZHNQiHg6V/Mb/6ZPky
SHLxY6wD6V5cNK9UEEqBZ5YOEpBPQr/dvbFK3p42YmMyrdoipgWO2rhFNxUbqlWwl9614HYRXdjn
hXe2rYAHOI9i5Rx0EFJDxzUdqOz2Xeo2rYXJoQdPVEOyH/7yXPk5LmO1lSP7fECummcHLUsCH9nu
yM0F23wPv/c45RaWfHjeEF4qGljdnkE3qCVJMzeyqR7+uup0iuYzqWdT7orrC+5YyUM/NdSNFH6O
Wr0/SlCwoNArvvalkjn5vTvEpgA8fSz/SC3EbDSvojrauyrTUeXnLBnh51D5lpXdwC12uCIdymyo
rfGgY5W6MDG3DbM+V67IU7XKW5e4F4A8jNfJGfHTw/0/46clZ/yAtoLbqSNbimdjCcjgwTcXfKC9
/JLDJ35ZZX0g1eMgJbu2CGoyIYSLxbgbt7He00FspKWrgsvaGTyYaVhZK+57W93hBMdsqDPz290o
CjGuZBPDQHsE1+/qW+UcPi9jT84boBgRwEmEaz/4HMe15VzgJG6MklgNoE4h5Fub6cC5ppU+URsv
d2GD62PXggyVFlvhcAf3WbVp87n6ZEhCav8fvCK7tqg+A0+2xK6fOuQ/NRAKK+MZNa5WPg8k78an
HqxI2cpKadZEr6fwit+dwEuPfqfxK36ekftQUVtTE8sl5zRxAfqk6paREiPJIPPTOZ4iPRfUzKPK
dJh7zzS6NYOO4IZyTxP5Eq4QGLSf1/KOmxE0iiP0/k15uTPZ01+weHnNEqqyjjh69vktpYCjvqgR
Hg/r5ZtGiGZPJKqJ1MVfbuY0qZUxTZNlkdG5R/bBm0JbJptbTSnCfROl+trfBjtJru4DAVdqkdwd
/aT/gu2CSzmMVk6KxyqEhGLM417PvARn5GgO+4ezXGE37v60/isj9y1PlxjvtCQmuVHTo/Lji581
5SU+/SVcaqWAR7vCfOwxDH53tm60O9WThJJB9nXKwVL0qs23/I8LK4Kiup8URx9FvvUpQw0lTPlS
Bu+Md1iwBkp8idW6LBBKqMjxwDN4NuWKJ/kWvuNfvvWVTxLL/7IFkZhRbNxdDZSBl65qaLDJjnR9
SfCJzr/j5sqhAMKRlMHDQBcIlC0DpGbF6Plca5Je1ecufXykg5PsWQXSAbm775jySYWfYn3/nfBZ
DoPFnzJW1ql2jZVGgmohUWc+W3/hRfTFCC0fSm12g04cDk9zkovzH3Pkb/oX7ev9ouw6gdAmUB+5
U10zaFh/gX3PgB+AkegrEE8ToNtmhLCbCTa9oQdMjUFQ+7f5LvRpLDM83t9W0hBDCyy9KYh7VT4Y
2pVT8st0cFpQFuFFwOPxlldH3R448MD9/R/S4jBGDSYL/5YvPQ1W1S+HhaSu6FVXPkaRacrfVCy9
/FGJhOsfjYSWTLB9HXIQZUOl/xn6oargu0ZQWaVx3dN0FByQUsJcaLfg0faGz18l9RXMLIemh78J
NtDWVmA4vXqS25J9Ih19GMrB8QriAFuiULtRX3KCjGvo+tj/PM/lTTnxFWqLrz8hDfZ3J+7PBH9V
EfJtzb/y1yUoiH14LIXuNsivWVvjDQUBsI3YDT58UCGb8Df9gkKhj4Mbdc2CvzRhikEbRrugy+B+
NUDhtanlB2GixxDQw2Iy5nRFHYrSADy0BfrAoLvEEFlUmrtomdwv9r+eqhOfzVdP0oHnWvNAFUZo
rneg9I7PbLIjElKtHDB3TpRnFSLLPsoluiAmltRldZSHBTNicR5x6ATZU9sO2rdrrSy5KJC8pmSg
p8RSUwd4nQnT8MjiOelR6tyD61sUMe7P2Tg5rM3WTTs8YYhw75oFmddwNWbHMGOTdI7PThbrNlsG
d54SKp9c1eCJkZU0Iv2EqpgH1cUhZo/Zi0hU197w3RIl2Q091GpWBNOdpc8FzPHI7ytceXTtXfSt
25NWpVbN01Siv2g3t4uG4TQGi6uAYA/Wt8yo1A9tJhqWnrw9PSPuD33aaL/aIosTvi3YQkASlbqc
lxbTu+WAem6D+ONarToPcrhyY6YL2tdomUafqhfLL4OA1etPSvdgaRDAzbOXWsuXlUfeYkT6PLhL
GVed2CNxkv/woV5Ov9qMRJHo5+CCOvhHqLjiyBnkjvTOBEk3UmKz8gFz2DPZcUop2dRGop0JnQO+
hacykB5pPEstzW4FN0qGqzO8DqzUtxvxr0VJzHUko9hsWYVw5PTLrJCOoQDgIU5oLFCwiTKmcKdc
7bYwwg2+3fr7WYJEmA8e4/IpZ/QFCpQWvwgf4ZOg2PhbiocbOoY71fockyd+1pCvavKeHEVnWynq
w3I++NGotXKfRmzjGbl7q5Hx5l+HEQ9AdChlmgtkkhvDrlDLxmRH+7NzJvyKZsTqsnoXDflgMnoH
wG+xLPtYEBGne1bqhJg7Wr46Gpg+287nGcdlKjtebSeLie9PZhvEHbpt8A7eGxCxZlC2cZ67vMx6
iHgdWLhdd+QpBeIeF4/fSqNn/TOpqKAxH8lbtlz5mGgrIDsu9HhvI+zA3PTIWKZcGHL5I/k6TW3V
/xQC3mi29JksPfIJQqlM29a6giAdmzZUNpITnFaNyqsyWHcaoD/qDbSbh9xBu7RX20B+sUXfIEUb
uK1eMGceAj+uNxkaSQrwcvKV64x2IcYadXb9brJG78/rN4Ihgs/685+D61L1sM7G9TV76TQBqr90
gKYQFJ5G4PqKSsG4SgZscYW9JKmdeFlDRylJd394SytlQoW7tLfARq7aXgm3ZDLJEs6b3vVM9PCj
RtY2b/f06hqq3lhVhZt+bKbm4z/bEYGLP/dhDy5o1gISMd0NAKnY0wgCsvTdIEQHREnffSO1wXpL
wJ2TmUx/5bgr3xnPDhPQMUAB4lVHS5d7OObSAmgi9nJf6+QvizyMEF+bq+gEvTyJaI6q+gTaQuY9
uEKg8JG5AWGBc/5qNK7WQcAQjR9Sr3sTdRDrkJFK0B7Gi5GEuc98EB5yPvzRlYS/3zciu31DYY5m
rlw/PjauynPavasoSj/lO6aHwqqwZPHwW/G1ZcmPeyJEzYhkVX/fKncXWn8FC36QiCmHfWTXHjuO
tmzSdbU04V/Ly4MWwtzY494ws9HWxs5n0z3cyPcO4uiC0QmW5/O5ScEzL1xpKFWRY99lPSqmxjyB
OH6VVz1PuQu2TTXwDE/mx3GuvToOKcDEVh2CGnc6JqPGal7KQcnf/+U3IsetoV1pl9EQ24WkM/9d
6isXoCubO5Uz2U0M1R+sNgpUcErQ15dAO6F2UkEsh3NBGM79LOzLB344bJnyRD3tMbPZtUirrSys
ZY8xsZiWgLqGzCY2OqjG9iJlWjTWBVbcN9aoGhlw/g9UQiuVJhLwYumuAWqClR1TKYsffUo5RFGR
0BZr8HAL0oYJWvONF7qbyCENRLsKqjrY29MJUbxdKDvyPlXpn5LK6jXavPg6mCsG7jXLZMx5rMW0
qsEarC705VykGLDRaiLcxqIt+NLJ0/Pg6Q8FQ9rJmGFiuQ5CmPluhXFBC0y1+32Wrqxu3b7iJ5We
5Y3oY7cSkm6RsFwcPFQKZA6HwKbeZhm+ElLamv4NJhDk/IhZXdYhjrHK9Ju1lhwCyp49GdOdCvNd
8FeNM/l8Uy7wq0FtP83/t0ckH5UZArbF+aVgJ1e5luJNszJC9T3fekstf4TXxJ7m70UTxSkKgU/P
JW08+zDNmHQOt7GOhTD/Za8FY38sNxANehnYs4JjO4cTkid3Ebh3vx6r85ZdLZVw1k/tTGW3E0D7
NBfFwJQY+Ajvme0qO9giI9wfu+r6EPHW+if5OsStAJneCR+BrSMFi+rkKfQ9FCOJpsfR/zV7SAP8
2hXonYBK8OG+iGUl9vfQdDrj5Ya/kN8vpJFsWcn2OiX7+fCCiksObKbtaUtxw6DjPcwYvPkVmOSe
ToyPjPHljhm2T3noI/3adYog8djCEaEZpu+92vjDKflpog8FkIWk7qM9CWvytAaS52dzxiB1EoqL
yxuNHNcKUbIPpKnsqrTzsmaR+z+MIb/1QgddiRwr3eaGXrRzM+CLTR00mKOiJ/ais7sL9K//7t4U
jyojR1tb//zWD0lFtSyXK0iIBSM9Z8zkPxTX4f7kyLq6hNUonXG7F5ybt9Ro6397233wACrMyHLj
u9J2KEZF9cSCFADPwFx8OCiHP6M4hKqOAfcRHvYynzuLA4GVYJnQGYRb8kMs5mw5/XlwF5CWEP5a
+MqMjI9dlh3HZBHaRbNoZEEbSmG81kNjBrgC4JLlSyJnVUtnCni6NJ8qGCju/CxN4pqcPOgEOzPc
CP9Oms+8FGjksyqC6NghgXQ13PdOlzAlbJonHED7zNpOcrHEYpkGNYDGF37E+il+ix2lWcMWe8NJ
bgGA7PyidGIf7+MPe84IKx7NPstzB7vycPOBezJvpnyBRwDGCNyfCfiS6ZFpVLnELfYEFXjzPpmq
xeT7qim7gjLcXrCGTfqTfyfzEnSyNREjv9WHhqYlh5UWFc9x2nkILnxyoBacBPVDD2IOWQi/Ei+8
OSlTFCfkzSHLMDgzYTVGp5msaNPTz8Z0yrkggzmGC67R63LVSxMJWeOPZdh2gRLul0cVJ4qHBIrp
frhpIjwnkS79Iso8adDF39js2GePwFG1692VAdqZBmIsXgfiUpxd0KCbxJu/v857n2JFexOOuHGg
jV4ClRyCKu/kR7HWNDdZM+NxeYiNUZ2RB26D1lhdlQs/qpbz5Yk7NBgnF3/iYyW6QYvbGBfetY01
aLVT0tje7zpZIbZLAHIKXhz9QO2xkljyCs1eJnh5Nwxs+Hd8IDW6d/m9nw+ZA8q/qka9IQxwhEE0
vqmw7zARLXSfaJoJ+309J7uj+n6hMkE0ZihH85+KY0fOYz++rqlM7HL22AfjGKQ0xcpkepfp5nnE
ZDAjwsSBm8gKWnctOqOytIwRgfp7bf/Jr1WO3KU4zRmM9ZE3jVDWljL6VIv32rTxajtMQqZjxRnM
UoZfs3IsqsDNNGHiPjZCopuh2f85zEbdH5GAiHP17RifZ2cSE5Ol+flowsLiKRbcDAuBUGn6bPHF
5rTmhq9ZWP+RZGhTSrtU2ibVrnVSKNE0G2uinqiu8KOLguYRuY31DjCg3HRZg7K1WY3ggiwaZbY4
yxgwFoN1DDFvOp2j/0rStdSgSp9sD6jHdEbEYuFPbn34mzduawnVXpRIKlWCofq8eZ0SjnIg4gYY
diFpxGuQb/zqQGxF8rIpFTtPzSPPmQU52nWpUUcMCTaQzRF004Z4i/SS1Krvkje5WQALdEWu14OJ
lUwi9PlJeBGp+TTgpMd9VcVB46Rt5PoUi28Q94Z128hmjklCMryZyUkf/x6B1VT6B88tl0Xi5+p2
HT7zL+jFog3mnfhPbQFVJQ0FpoxNQc20aWKYPVLIoxUYJmDjVzeaQH18C5I2p1lxBtG0BXBcwdG3
4JYcW+A/AWvdrmpuUHdbryJ8rGYdpxTax1cPr425qV2VvCwycUu5LLlUC7hr/oQvEcSHwsxQ4QKF
jOkUFTuN0VbLqflW1fMH2YdRxWHo2VHckW2v1aNnZqukOHdwQxnvC9o8hXrBl0gscubQ9eKIBKWQ
5OvUf8+UWBubuCM0bvbSkSUOzLE85KWdf4JX5IneVaII/elW923VDfqgP4rPqp8tQI/Wrb4Yi/0k
3bb92mCBto+b93iIYq67kQ0N8ysb5tf5SIotWMYrmEeSTR6rtncf5kwc9lsNLIkZYu3HO+lGRS8S
ipiw6tyj0Dc0324c8SAXKM4QvbcJdGelcoI8ClUC6UgNQx9WQTQUKMsW11mPUgdUc+kvvw9/0JUx
6J77N8NjfGNclDh67LB/bQtR1OViDft0Cl0cSdIw9yiVp0qSkovFgUpHLFNrNXtAvcdolDGotM3j
2Fj1WIgRqYzJVQ9Jsnhaa+khmOU7Km5O6lwMFqP4447z0Xqnv42wPTKtS3tSttjEyeps/HVcd4Dp
uX7oakmKFD6eDs5bBVSI4pYE4L6JWwZit01qXHxU5wf2k73ccHGLxcGOVKN4dXwB7QQckwkfIgxD
dx1MSnBfgTsxvTODx5V0R6ZyzypDyCTZLqNLmkYWgm32u/W7m6z3Lc2KoVJrpdDR9+jDpW7BUeKI
nYqU8kH0hl8YU648UpsCmO8ZlkLwQFak2ZaEew7PB28TGzgKSRWwRzC68FWinSnDEav2jg4xBdnJ
GJu+gwpPGIQyFBVIbox41rzSR56Y4mxtRhTTwUtrN0mYgcHhp74sGXcyBBF7GOOkZ+RevghaaCXo
cJYahPold+90XrsXcxedbRHe2J9lcOqgkYLNI7gXj6FzRxiDYpumgn1MGxFV/vhMHC0vFC+XLwTW
+wQrUcMuFtewxYw6oGp33xBEP6/H1F6kRoBPNXIidLMGby/cPu9I/iTEsc97o5nMiXxjpw0qqTVe
AEx4OhpweU/tGtB4RqcrLHjkPMq1T+fOENa+EvM3p3TfjBvlue77yVe/jHrPnsFWJogihB2v0N0k
NInYC2Px0TUJLOwjRGRmq9nVE+rqUXat23iP583vgQe6dd5+Nox3/zByHUaR7x4EuTBx5HO5HjC8
YaEGRyIseuGqOQnvkUyKiWCEzjVsgCQr6sWj5ue5QqQn2bQTScuBVsPpOT60gjrkP3sWeq/EnLGW
okmgrkRBf38mSaGZwcsbahKVqdvR92y5FO01GyLGudu3OqLGN+FhAsiBda/3t5ihIWHtbMQKtSjq
DWqAUi96pgRgL5A/zuRPcypLaSBobZjCxrhqRwYQ8t2iw3FvbpNAB7OC9lOBaMODZB5YYeuWNL+T
CrDh8pxUCKXOLjTAVTfRE+h0wJy1qYQkToPAmPrhsGOxRYUQKXL0Zl5RW/xHSQ1nDjWfJSNe/GHT
BteFuaw4c8L47KzLcPeBnNKgeogHPxC3EzZ7w2RCLclNGWrSmO9lT7RrYpR8TLu8qR6Xrkozl1NM
9Q1iXekwXs3Dj3NYIJWy484etTos3hdM5Z8QSXnxT1g4L+mrXDNH8yqLz7lz/i4fBtITfVyP2fVt
kKeqfSiNGbuaUjIUO50pWrw/TON1hiHSRFMuhH0PAmiX/mhG/CvlnObZvxUEAxZoDNaxWf53oCtm
LMaA8X+08gfpLkSXSxIBpGk8ocJei0ZmFo3pm7kyo1VewPDfhAohcqAfBZoJlefVsa8UKgZDmgZL
s5Dzh5aCAdVcb7jfWuozc923WaXZiz/g/2faWonayzWkODXBHdjycnJzBkgf66dgFGQHjS/2uFK1
onN9ltctz+kqRE4pUgFAG0D1Mo06tvuieVq1HKX2rvrxRuWHSGU6rw/DUwUPU+coUu7zer7U5UM4
8+J6oLNFsSRp0SC/MG3SVpjqPLXJzXFW0MfLPYo1z/oASrjBElQ3QU4dVZerXKGyRGpjVUUcaXGo
uoyTKekE4PcgUARKs2iDgKDrylxjr24lZSC/MLPgR/nUjD/prOm1A4lQgCcwuwG5x4Xx23MFSMdh
i/bPI2uJUb4yMbPvP+aFxFoYITpEvNJvIOop8M0qbPsYfsftLYc3/9dTC+S/4MNkMkICtXBA+s9W
HQ6ltJ47pHuL6BN5ltjX7tkh5KYybGbz5vyfmsDRoAIz9wBwX80+FJleXRuuuQjPmZKSpTeUtQbd
GCX+iXgG4jPdpBHJOWZHHckqgl3Nh0LdjdI8bh0XSkso58idelcw/3khCPWm2cQtdrIGQOLaVj/m
PsMW+fovnc0udnrT4tqQjh/rMK7SQm4XF/MMjg12Nir+qj8afEpn6Sk5JGcC8kjt7Z5qlEjR+wBF
2PyinE054343aYqB21YBAJpHKvM6nJEx1C2/RloOdFoNbNUfjhgG1zSES3YkZZ7SEsE/z10UGlPx
0c4VlIXMYqzFbOisjKDAPrDBBGXyAH6hxzPgL8/YiwJFaj5gKJlwK+0WMM+ZvlzbanVmhios2OMU
K1GQdDhtqWzYuO/fNW3MAZ5gtUTlWCFAVRQRB/4mzCsJ1JkFh+s5rRmDN/s4PmnLWCy3azJ16ubE
i4WR0bYPCYeTkruTGgU5RCe8yKu3CfR0j8vl6FiVNSaSOu0dWaQ9wwsOgSBMa0S6gUJQyhJe0Dn5
FXwWSj/VjBnfndL7KNVXssqseSLnG50okXRII1ZYmTnn7hVUbTtro/TpAOuKliX3NhR9wy+swlMo
p4i0MUCYnr0RqHz8FwxIsd8O13657j0Ae0u3kSLaWoW2SkO4/tgXU764CTXy/hShyme32+cvWUyE
UToRQwyfDXTnjAAAucLeQ6z/9/H+JbUDVhMyA6VTcGujivbj0SVunZ6k2bMrREMmUMBfUn0OtnhM
edGK1CU9+gUzko/FTB0TjGa1aFHY0cKkbBfEylAtCF5J580/e+46X1AkdsnfvPn7yUEOTOWlmMKD
1SszWlW73UDS77S6+6CpwXGi/LMYls3OGL5ycxf81dZjG8mvbsrTa8m88FSZmHdvTXTmo2Vlqt/I
Tt5FLNgfHtAzHKnZUx5MUB6yAXWtXa9PjclBT4OA/EWGlWBsj63rUCOGQXMCB6tI3uCGtts+KTIW
+CCFsnS4+XNiz21L18SkBTky+59KjDZ12IGdY9REtd+xLK4UpFMd9LrbOctFU8jipM04C7B++yzi
ipTFUoX6AG6y25btSNhjvd2E7SSPbvONNGZZ/gaQHwExJwmcqV5dJ7mKLNpX8yR+6rkKO5Z7PNYw
qbzUpe1Az2BVPWFxQfWQ58WvxZEHxhhGNs+sZMGheuaxqar9LmSH1WvzviIipHSaQcy7QFrxTk71
mMFD8VJzhmQI95uzIQvXhkqM37kepJ9wZFXNWDZaumTKJvPCtlZ5qowHDZiu2HzhHDhu+ClZPv6V
2/znzf5jE3B0Ip/4JTFi08Jks4niqBfqv9OXg5R+0x5TdWbFLblgQ0s1PzWVyPSngE2VbVOUfJfv
W2ZoDUOigdNqVgHxAy6IZu8txkIlkEAsPiEc1luV6zDej21pI2+g8OVoaFqvJfVOda8NpV9njZoS
DDQ5bujLszZfECUNu1PG//CvxlrzZNe3wlJJHdTyCyMYFLuQDfj1GC6xuhvo4iFiFtDry+54s2rE
RyWQ5Ew8mbpkx8DYIvqBXexHr7zUzKk76EorW6Vf3HsRGEojTQCxRdYVUEY7EvOqaGrjV4i3SMH3
ccp+X+QTyj1whtTy1zptZszmZx3N20lJ9FYU0e2LwCBoKQgOgaKA+QAmCF3c8iZt+rZtA6PttxUh
rkygSOrPEBgb1z0PPDvz6wuvG+qmDmymU70apCZ7P1vUqovlkWxxs7i9Lb/fapHGS7cfowlk4uGX
455nlbNQpz5YdlHb4efa0U//bnK92kU4GJh4gnRpQBOsTvm8tWQYsImWdzck1KC39qwY/1D76hwG
9CnOvf38OFcQ2GKNTOLDPbc8vpCgzSEfURKit2Xi5oyfRpJ3r+e/I0wfOg7Gl7O8FcLkqNpEH054
zgewsk2bWRfRMV+PSu9XS9oaHlwU4B395A+/KLW754jM8ts0q4dD9A1Bd9R2pQNVXsOybaid12lO
xv8Y/zjJpCBWVZsYzJhIF8DIvdzMQQSbO4dtkxKfE/cK4k+x94OgjGM2YXjpEgzXMflJ0uauHW91
dz5dZskHlgTy65gxlM64YZ8HK8SRyKEg5DJt3hoX/Q1FgsGVqrYeQ2cGhRFESXnLRRMEtUmjxE/D
Wgl6jQfvCu6J86FHz71M0cpRB6CCknkerQdrfU2z7nxqeo7CCMVLykqcMMBJ9na+uLG3oePCWY0F
kv9WFt5rGW0RqlNc+MrOXvQXbyJQ5CvBSZbqEnIz6loOdwE8UrAWziQAYvihH6drloXdSd0TlYDB
5iOr9C4+F7O7w/911U7tg3njy/59RV9vEXGP2YCE1b3T73HhSMYGTWKP3/YkAvq1hPFm0w72eJP0
72ErYnfrz2GR+I44qL7I45eQPIkBeQQMfGTKfbD3/ZSYYJ9RRwebE5jbYMX1cdAp0DhTqJ/5NmRr
Ljr7vrazS66bYBFtlqEzL/uI5yYmrO6mgXacFKBnG9ikw/pCefk/UtiBNalPehE+7JFGWCJR0zKa
pi3L4qpy91QsT/eliz8BMHjX11m+2m76OJHRnlivcD60/+11tUwuCJBwnW/37GvyPlwxvBUXg5nh
3k2PQbpYFTd8dovciC8Cwb0wJqCRWb0A9aXgc53oM5K00cnjBtNZovEpAT0OPKlkxQtC0rHniQvk
fmA01WzFn7u0FwTtUIkEmKHC8BTZ05QZNGjWfEJ0ELHs3FvM8AY+GPdZWKDGHWA12OOT/1SGfyP7
LAc0Y+jRtRP3yQWQD9h8DRy0NTnzj5d8wwXjINuxY2AX6p4f4f8oivw0SDXHALAD7ZTm/NdR7M9+
vFig53oTp+bvrmNQR5tWI3jBU2rlGK3J0I6XxgWM7726X/QALEzVfTaFKY7BzJawYcY448YV2oJX
MR0UelrCe5E04yIL8Uf5ZUbqcD8mTeElY6aUoDpB5G9w7ZMdMUbQ06zLP96DQKwipLFtD4OypEBq
hi2EqJfKazNZj5wANc1xd6iIzmV3lb9F/t4upQDD7ONEnhtahUAIzv+xLWB+74fbtMYkfarn+CAZ
cjCghXJ0A8qOCxBRcG9qx68LddoIpk25Zc2PU4nGCv7OzHTfYRsRS/d9SAF8ydxS4P0jPM7tqJT2
XRn84e1g/xdQq/qZ2nTc1oGOPQdjl58FzrZfaDeTMLtUW1Z+LTl5IWo1JeP9dqJcztFPea3D5h8z
+4jkdy/xkRSTdpBjTjpbp2k3yO0aNiIDY1QWVjz9+ohxINJYDucR+NSkrwpxnDmL6eeC/jBrMwi9
UGJ2y7mJXGGP2nrT2ObYyYIOJIKq5LP05nIihs/mYs88DQro2OJYCKsdGahvn28FCnYrBjPxPYEN
YhGBprKknne+lgy9Zc+DT0uysoUesEsuI75WtG4XdM+TTgKyeo1366fkKp5w1MLkK9eM98bsMkXD
tG61OeolIyefli/0mj/XITwouqOTCyBEMdolr/kxNj+tpTffjvGbhJmNyKRYBrUTmqAJMZAQKTeu
E/GhQEZFXHyjSvciX71r+HV0mH6edhH/W0GacbL8ZHMKp7fNirMjgM0rSxQIzMqVWIKUKD3kVfrq
cBf/57qNI/H/fnIulqUWosNrbn1EZWw6BaiUmHix7Wd9MYT29L9soj8no7X0a2KP7YAnGUNJXVZB
a0nOX45mwdD8J/7Z/DztuvI4vYFmjoWT0a35Z3S1HInm3VLo94YkvlUb2jK0Nf0clWCa5mTNLM8v
P7KPHeJJeQmDJvrKCyF/furk4p7zT4LDqy99NnuX3jgMiI7U9yGDAJDQ8kq4wBXwi3YKQ1VsXVXX
SWoITgEMOZpb+jyuIkyxu7cV5v2fKJw8fCIR+4/pUfXh9tKz78KhMFafCS/zzNZtzsnGLO3Oue9E
oh0JkmXrWK56qUcyETFmZoeELKvsH+hFOaJ6jpw3M94uC4fU41vU1/VWW2Hj6OpKUR/lIAubUTsv
vmm3u5Qar69WPncNDJr/MiJ/4WDXJrNcOIlYjDtlfykBxlaNi8Qxs6yubiGtwdstUxGcZLk0cabQ
XhDG0MV/Y11I8bT72Qs1QH9KAUzPBRYSmkiuA1jlMoUZCB8MhSrPGuNm4MFUwwhzwprAX8MVAh35
ImMsAhwHHffd+NmSyg1zWjJzXcUm2ab34UJg7aiLOW9YewxWufZs9jDucM9YBVtc3s6BRyc+YKyV
q3t51Qiln3IRQr8nXQET2v12Ti2a+9TFVuQhoLxcdjHykcqZOXs62j23L7dwa21/QE83yPgYae/a
jmfBi+ZOoxsPUKsTgHV+uStBG4OJwJBb1MtAOMhIzRWrl9qvwrpoIFsOkXWXdM3SePosMhidaxFz
XRESYTAzrC+s5tB/9T+CLvJM1TTuHkg4NN0Zo33NCyXt6qB50OEtfT1/W18eWMq0hcqzBG9j4W52
VITIGVOXntR+6c/Kg1fE6XXm7NEpv7E8BFnGknSCTrOUvA8wDrv9fmaf6s7V598aa+q1+arp7RsR
nw3iC3UocU+qSnO67bW3iy3SgqB86ELjzI3jnFss2oBSTz86VQ7tWcjAO6ex1m5pVjGyxwsv9PaN
f1kpFHxZh02ieK8BUFmvXTafThQTcKSdUE4wANZTuw3Onmz8q+BkN73Xpgvlt6YTEC6CP32LUTbC
U8gqRFqVhleyPtQXjWmg+DeCQCM9FafkZ+A0hrJ9dQzilVgoCtSizBOTkvtODF5eVNSUHd3pYN0y
psw2BnU4lSE1wgWW7dm5l2HYP/kKeyIVrjWDnfL/Ju/7jRYgtjneazqnHkBCNspnahAlT93RsGBI
Ze/WIMqWFLI4CeyUU4YY4q5LhwcCFwY+qRcao7HAf3tsj2coiSna7DmpIE1a2LUylW19snrPQdzY
5pvRmD3Wo6UsAHCoYjmd6KHtZjlyIYzOuSJJK4Fry+iJtJji2aqtb/3N/+H460g8BNCfR96l+J3J
O8hB9jed+OCJOSjp3cg1F2qoW+XtuWv0g6ZCUy3Pbsp3BUs0Ic9MF910Sr4H3e/e+q5+JnfbwJkP
qOGkLzxam0J1B5R2DBJd6UnM0yPa44ZbG3aS7EAUDDQ4zkoTmU6OqrB2aWR75pXrlj1hwD5u4LTm
goRwAxfxFxwtI/PxqqZ9Pl+RWI33QtxQk2gTSGv9ZUcSOiVjS0EFW2VV5UXLg+cm4s3nmyg1JGag
SZIIDTYGBnlSyVT9S+WufP8f16bHcFT2E98X0KJI2Tf782Etr7LSMz09RJ8em7h1n/mNPai6kDHV
WkCuo9/EZV4S07nv/lVOrX5UCiL7YIBZhxxZeNlN/6zel+cGbRd0gXvtpItkfdxQdv7bD9xsMG1H
lmp1iwoOgnv+0vbQOozlra3RFu9ZBextq9Ktsx4GOHt58xU/8d9ebNxnvbdPCubbJl5QyMmvyggO
FllySzVjZ542qAL5xKeW8aObGfp+T67RUnfUf///XOTKseb1eiZdiFeVTE5+y7YPolB2expa4bV9
djDePlhF93ppMNA28YJNyeRhNcpZNldzGHmy1VdQu9iDwnE8j29A84wTRD7iyLLFf7P4ewaRlN20
2vA1Ao3da1p1xPZXvak4NDYt2SMiO5Cxc3n4tGkwZSfxwVUnFP7yDrgvHuqDf2zCYiTXfD6fLezG
zSk7kFffkDvo7sy0oK7FC8wX3Ga9XBSAg2GNL297+dMZgSfIjhoW0KbaD0Js5oElYavLn0RF3sU8
tBnOY0CNW+YWTqGNgxNCbiYixwloVThRukwtP01LFBvxunkbjRH2I55edbKaF72vXbO4hI7Q7Bno
/PYtc7U0nM4Dbk8rtjpGRTpjV6TFq9yO7ECFbPOdvhBH3NmQpkeFbti98GVU1oAWX1hkbOjuSol1
6KNVkiPaa0KHVPOQqA0SzOqCvyN3Sm3nLfmHsAMlvVaICzXp1HieTEyZJAfOG8WriilHvC8ZCJdZ
gTcVzZvGWgiBUS6bu9NJOwdqZbYSPd37xTJXQtS24UCtYDX3L9/2tdLxyF8ZZanEhRBygnN9wdEf
S/8u3roE2sC5MM5oHKea92hZtx0DtJMpuywbdRlwF5ycUih082KE8XcCT1GoAriV0zq5e0numasX
y5B2QBPvnqzgo0sb2EmbTNENuAEikBM+8KQQx/bFsXQI/Vd4RA79QnDU0LDILq+PDa5O2tR9StAw
CTjN2igajL+wJ5aF6pi984ozbUqpSBtjtuD/TMxa/jTPtsiHcwvyXV3NgFWkm0eLO/+ZecHZnb5K
WWwe6Ig+W9nzqc0xOZrbZMRmz56KInQu8ZUxsrWcnh4pY/HB4IVnJS4Z/spC9kUaiSscCL/QBT+o
pIeUQNtyC5uacsEVaR3b6Z95CbrYdNgx7pbhBDrzy+2/yMs/N568bYbuaWN1rZaHSxCrgEyFL20g
xblyxlX3/ppVbhW932IRNWHpCZwbv4AxfjGk8ZrCS2De2YblHvknxMbFRZizrxraaNpOATGoHcOg
/eDrU9ahD1bdqN3S6eXkUWwAR8utmg7mtVlGeDqMfWv2Q+Mjr+21m8UsSYr9cwOe4w2kjzk2JgAg
Lfj7rqz9ved3gs7pnV1cT/RYeKwifyIf7eUH+ApXB2QA9S+d8HVt3AcYY/h5m5ikyHllc1cyJV4N
9VlVwU+ZsfolzEoeOZBorqKzY9mpJANBVwsEyjksEMmmJ2BRxusCLqdhKo8rjyWGg0GDfM7CDwDI
7rdg8kPJamkDl/S8vTf9uwcHQOWdh01UCw3ITW5wr7OcJq+xCWWnVvZtoODBqXC11iBIAy9rzahN
o133JtM7fP9sWRCHXi/k+2DPtMAlM11f8srlfAyaqrqbFt42dpuTNkA0YQYLSsgGUdzWjQDzCI3a
+qX/vsPQ5z1jndgw3rZ9eg32KOVl7lBcQakfQmWktNAp6aIju2ZOnuFEpK9NuBnobmXEcmG32buJ
vVfOXF3qy796Uz/ed1PmOXuYrkYLMBYMi+QjLXjwj1nZrZoYzTETt+l5QMd1bHt3TTRn5/VXtuxP
y+ISJ8tIgxD6Nx/g2bNKqFPoKsKm+TUOGhpWO0a9JYrDzplKlrFu7Mys8z6iuXakOHH0idJHfbiS
b1LBa8zg9mbSsHU2qCPRrgaFqJpVQGjxiMoKSbFPkjTflk6JGP6e2xC2SrBvCG5NoiVJ5zfQ7VeK
ffy5YF0HsUmio5h6YaIcg6jxRJAHTe/QqoOBgA2Qi0mEYpw6W2qvEnzAjPImeKhQ10S0LTf4AC4F
zkuR2Ww4kUp4CoMnQRAeu6fc0rRMisILF3jkYzAME1v5H5peP+9GND6yLH0dl4Ma2Ht19pDTbA1j
bsQ6w4VQiwECAGPy39pnjgvE9rONhTtqJju5mv833vQd0mjZzjRsXLqKRS9UbDAVc3fcH0eZTS44
yDMNvS4fOzxFidTZpiof3c/0YURh6t2vuMqmyjXxN3jjl5thUzF/QzqIMJCS2MOLxQaan1+xVxU0
au8p9sbPeED9lbhb9H6TT0G+zoC1SxfBd8evPQNp6VZe9qveOp9vLbMEQswSzEPrLNtVys5lxenk
WznDlRUhBnfG6+fGzn0tzt24VXsVN4M8yVfl43uL3zF/W5rL7irug6TCgAu3eb0re3m5T7fZEccv
1Mmqat15hEiLvoYsF+zuldK+QS5vxqRiNXplXf3hqKMUd1NaagJ4zBv2S4clGqzMPXz7JqOrFtGP
SB3LPJv6ewhx4bpjHQiIkWKEFb6Wv7PTdF8yEjBOpDViprjdPBrLlbNc5a7J3ZHG+Pfc+jWn5hIY
tVqXG06D7CVZ6Afx8hMQ0EjLKslwdQ3S4UDRESi1GfsFIunhmImnY636kKPMAqtJeTT+nSLTdIa9
jGzo1sQ4CiMWKCQv1Fu1GJQlqHAe6P4kMJhhzKXWl/U9Ut303YMUOi2T8xoSdJV7OdV5EEMmllxv
/xl1wtIecA9g4wOYWgpNsW8gv+MZ2t1o34d0pPP7BCMCkB+jRJ7aVvoCNLdSrwAEKCxa3YkASMZx
dFlH1Bksj2Du1BGRSm7f/5HDiphfIZ7q8dsL0JihxHhsZKhszhxndQHZhJbFlsbL49eovFL9LWib
2gMNRELbWDemuLsojT7VZGqhvK/BNyd9NrBKzHMFNTWigIcRQn7Odq9N7YidrY4s0mP1as42LwXM
M7r5G7fDtOA2FAlifDJyLpaRexjooTZx2VXTYg/k9pio0QCh3xwI4JwPQduWDK2fOXdg6LaSEF/R
c1SkKPR+YyWgsrwrP9JAv7Cok9bQf4JeQPwgUQfJQhi4OZhNSiYOThezf5iGHBXP2jKhoD7uu277
mOj64bp7I5k9okDEc4W1o1rrPSQY0+g+6TCoTIKENK74ruwMIUYYZqK/xPlyg6cQEwBvuWCEXiTk
w802GKFihXRoFvrWQhXIgWdusMDme1yjqZRtE0oP3WuWHeKBGxxpTtSF3Y1TEhcS5bboYCbaLlNc
G7J6YtMzFe3ABgh7qitCFTLPVZa8+rCaWTDEjOa4mp9Mxn7S2RJcbG7eU45/V/uP9ZZmFTyT0wva
0HqOjbOyLsxUDAsiS2MmfTHd7y6o/UmRIREhu0vK7LTsSiidx3P1AsbO5dxjrb6hu+ue8bGf/Uo6
sw2uWh19ScY6LHTXY3dnyO9kUthLAvIri4nw9BPEjVy1xxwdHFarR2WfOaAKvg2t0MZIJT7tqk1F
EjGH1hynVx5VPWuO9wRoUykwbCecKph92JATYJ1p5zksmM6qz55jtkJ4hvJj0fck/s2HP5kVm209
Kxm1569uVpaI81leJ8Y5rG/g8CYrx6TQZ7On3JQ4H2zpNgpaLk+mj6hQCAaJuQU2sxzg/6jJZ569
Y75Zk6a3q78kx6+Y5Dam3xG6PmHLVImIcVODy4NZxNZOHdNnb6GZNsm7JzI/3mo/43nIiLAw+RVM
HOGV7qCLmEvZ+PfcKV/wBo9J/wiouRSKhfiZO7bBAvDuJ5VaIzcQtp2CjAeIBw2YY4nfPmGp2zUY
Z4ddyVy9wBZDNETu7RZU7qm6jH/d3MKNw4NLUcnFmkXIi88nxakxeSStoImZcKXNbPM//9Aeo5ZB
fonjtbm3EwUZM5m8pCxveTvc/+fM8E94EEXd5xfUJlmestiv7PTLtRValoES4ExeXW5HZJa2YeBI
Dx0Pd7volPoARUTyEyxN4sm/o930qNc0GoBPWXbnCPCLOMTbgqIKvy0RgJVMu9E7pY0heRtcKwF4
daf4SPQJSwoohtz7CCGoKGxncvmaufGHLw+thvbqWWC9r0fGttuGadZ+vL4KqJ7XUTBb+IqlY6Mw
+R7NUhcg4v7KIeZ07hQ3thlqjq/CregJJ5VsT0l5kMfdE0OICWiQSB37FUIs0vVIeth/56UznkhF
HW1OciMc/d2L+50EJvLlmR5ZmbzZDmo9NLlGb4YLPwx+ndqAexfQzefF/imaEPpuxCnhg6DMJg6x
jSTeo7MbB3n6j4oLsf9Ior0f0JEHLI5f//ECfkmGuuVymcS9N6WZ0HvKvsTescT/AFcb/b52yS4w
fNZb89XoVdFyq/vVqVAFfTuXXzBlnZ/ZZT8CrlKaPiabKXmxOK/tyKE3KXP0e/vOTgmQh2w+xnRY
0UelhwE5RSLmSZeYmGcHZnO5riCJhSrQ5QjHBN4+MMHookDUfRih8RdGIzwNbUHP1i1UFuhG9VK2
vD6iOLxEFNE1ehsuwgBpFpKkQ0dFCfyU2QpNayurT2jwkFLkCvSxdTJ15JqnEdnuoU0baryvpZ0Q
0c1gIRd/TBXXB5a1aTeQf+3h234j5Bvj4Urg2JUlZQRnhSh6wB9cnHakShBAIoRvhPf0F4eN5xSf
vfpN5ky6NSuiSuF6ilaLBghjnc76PTkFvvO6eFdRhwCQtJcIu5dWtHuPb+OQXuqNmo2Mv+ngMDea
nwoKWRlPeQh9BQ+vSrxfuJXjNECpso/ee3pqk1rSpxJrV6bdhow+2ZU9WSXEt9EUVtjb1LjZA6LW
pXlM1Pcj/cLQXiHpUBpxraSykpyG8M/zKV4LUfBgpTwhWlIhOZfXs6Lo20gGt8BGWY2wUpnyhilv
vhudtI9G7IgAxGG1EVd3epuzVKjsiHysuQc0rJh4XUtmIsr1vutk/8slKioLcmqDJYKKEg4QjiS8
WJkT5tK/Ce0H6XbZX/btoQVfkk0yv5emFJrf81vtv1Ae61y9dcq+f/VFqeTRyGss3HYSSPuWWsZb
PTHfy1XzG7rCvnbm7pHGc9bnhqOHuA5rVk0QNI7bpi+b/vpqbaJqVM7bh42HqQ61eFAiB0eaY0vE
afeWk5Z/AvqcuXS+ke19k4kKvkXBfyR86k21x42ixEUN0L3eX72g0lUQKKXMpm5oRHUSj2Q4EGX5
oV1hKBJYmTJOTo0LPUvHPEO1xj+HH27wgDufXZiovSf5fu5ARiQ1QMCdRPuSQaFt6DH8vo/Kytni
VqZMU2eFr9uaIODWRrxiNm/pb3yJB0V2urZoHtouAYOMKYar46QtHQ/auRgjxWxcE0WcpioL8k3q
dhXpv5+b6/8TYSMPw69XvtekfKvFOH5Nk0YzTf/BaPhNe0hzaE8YqJ7sTvrYFyMijTptu8D/lSPn
hJBp7tz7mlUSckKsJiZtp5FMGyTpZdCWG5wa4Zqoo2/1Wl+4SvsRP1VtnQTUTuhgwmSZWhPQU02y
J0Y1l1ipsbvGPxY2a5jzQxc5EUu9cgBfsbgfly4OQtqQmMiVcVG28WcM4IX3pOhDdB+D7XBX0omH
x/P1D60Dwa9mGFa6sKvr6IZ6gAzcKZdnDOAFHf4if+n3oZeZykon5qe4Ks2KhS3AahbDyqp+vX9w
HhXXVXABx5mrKgxAYSE8BM5fX3cYKqnEimSzTBqu4MkiMvEx7+3IAMil3zoenPN+81KIDo3gxG9r
qN7qsir2jai4FpjuUo8tw2Jb2lPH46zbTQ+fjfJCR00tZ/aRVKHqViym9Q/wmfHIOHS6QQ70tV7s
YeTpCrI1Tu5L9nssQDdel7llEcpRahxRKyxmaCb5WLKXMSzfJswlZncVNk/m41UxTmPJDcc3Bob5
ceheCOD/mQOwakSJ6hTmC10L1P64sbeEMQu4ze6N95S0qmhKe3HqvFmedlkTRAwwEOIYQnfadUVH
QKTuVQrMADayJgKMetNITPEVCUMzvl7rFUbVTVc0CzH5MJB5YJrlolS/DABOPl7Ja2YG1XB9OPMQ
ppxwwXtDaR7FbhmNwz+sBqwplfcsu+nymQpmensPd47mbiAhKRkZ5oYn+CxxvCs9F67Kg4TdDLSh
3gzSnTRE/W8rIzVI/2iZaKF4DAPRBhlkUqA12ZZgls/o6O/PBvHHkKijNKpUur86WJppa1AmpMTD
dn8nbPxOx9kGEHUMTxQ/vlwjp3/f2gFt8EuG6ROrfDlFWnFna154FuNraHF5dw/jr+n10JnCmzef
GeM4FQxqdEBcJykokBz88TcMtZSY2iTT1VT2hYA+pDnAfZZ7uc78ed489KpWYOF0o98wrl7YnssC
kdjTURa2ZR+bXVb/5IgA2Z+HNwDK8CZDnRhFOGFAFO9zmqdj/9Ki7lUDpe6nR0Cu2p8BnQlq0gEo
kMIDwZcWwhb6OE6m6d13w1poTJw0Xqoo8dLOWFGPNCb4AnqUCTq5x+si1dYsn2BI8mRuLvFoCAXj
EhOm3gHmg3qg5dshg5iRKmP27n+YeJq93LYpbLDisVC8lTXdZWBsvYbSyKGVsHpy+GdFiiOueLdM
bnQfsDGIkqzP9r/vq1vB7yFKohz4KjFTiWR0+Y6eRv/vWXpwLNjgTJzp1xQ15d/ID5hw47QG32KF
8xGDtMXnK6u+XOWeCV4tWaAGqGA0xSqS5UHMnADTw898Hku/eSCseZwW69fwscjWvzqD60Xr+s5F
NOa5dBlId0bqKr6uWdbI1GpN+M67yWaZlcdUd/2KtzVJh94tUY3r2Ohq95N7BendluUQnFSDnkL1
/Wv8Wt2FT/hJ6svRlj7RLJjylmPH/uSZhnlN2r0SP85uZ74w4oOCbMKXrC5Xn503jNaFHyDvfYnG
J2ZRmZbgDjKhZGXlXB1jdq43ZtJHrVl0RXd3FN6dSajc7NOv2GAMlZjdfTpNk2NkO1B6ooPnP32I
HbdYhq6k+fknbkeFxcy9uJ8Rpvv9s3yVTckKcGUpzVJSsWbb5ULfJhsnB4xMZ0EyKMev3g50kl5S
AsQSkOX7NhWfee2xvoJ7ViktRmhZKsCyrcLdnfgM/HHFgvU+z0kykQWir/WS53ha1q02FOVEAJO4
WH/uBjlVI2nHMKUVusMicnrDIG8Targs9cwCBFzIwEJNO+917u7wA8Kv81VzkwYuM7cr65jlnT5r
hv78moACW4VH/LWDQjHjAC0M+mJC3LwCe7SJWdLjarzwclH3dVgEVqptIAoEwEMhVNhohap1F07+
jnwiQlmb0EOLuQfMDChoO+ne51/QixlqYlgHG2/DYpxMeAUhTMW4mB+ZQZWTiRqcLM7OEIg9Z8Oc
O9z9I9vpivHqAR8AZhrheaufXY+81PRbXsSTiE05mJGfeE6nxc2llstlGjKD8F7zYQxHzZ8s1cbq
OeImHQCzCKBsl+GQbi7gvk3DfwGFHe/7k2f002jef7PPeVtlR0SXrXkozr21SbMPIVDjmDcYODhK
NoYIFKcz7jqJYCyWMCfwut+7H7qNxLY6yrft/KdxgyN+UJHyTgzWqKQ3sajunAvEYJX6JB1DiWI8
wsaTbGdGI6jDJIV/irGVznN9ERtlfm+hfxwLBHpZM5a3LkFWF258PgQb9Pgf/N1/t9+7gSGP460q
E3Fw9R/E7hIqgFssb76nP/W3dFprORJOUDmWyC4uFibaExPH8jY0i3VUjr5v5Ig2EYfRaySLZ8G1
FG47AdX8pGC+6lohl7zh682Kbow4vWpW4XkAGSrvy9C+SbJJ8LFroGgfw57ueK34cKR6DO7UIdOl
wjOre6gZxpLXg1JGuUHmrHYeQMQO6x6vBRDgP6WArYwZrC2pYkkpOQy3maib1JudYazPVHz0uw7I
ygH8yeqpphfZP4uyhJwsOtRHJIBFBerHuYxS0rq4x31AXANaVSXrxwLlnu2CBKAGcvcXxrFygF7C
yjCCmeL8RX1R6rUXb+7KDWO60AcOQUl0FLGpgSvCPZqkX0l3wJxoKAWtCAkcjbte59usEfdrTUDt
676qqZRneaG62jy4GF2fdCBKjqb1Bnotd2+mMo7jpUeUHry6M75/VjR294sG0pdItz0VAl/bH76y
RMVyCf1skh0b8LLNkx2wa6Ekwat5986iDRmHcfU0XJsimnJmcFYWIIvWOBkD/aaSOuNItwlZkuhF
nta9UFO0pwhq3cdgSmzXtxn6e9TgElpJ36sG7AHKsFTFQScoEnolxCGV7r9DMTLDrxyIX//bfNFt
qyHkjf4jCu78n0fuXdYh+J+VIllwLFAdkdFLbT3rVNaV3r3pupuqGdn0eAoyfy0Pg2AKFD9AZ3d/
RqbavaHUarWoX2GwioVVAeHIYfDr6aHh3ZcztS6uUvZjp3ivYuaRFk/zI0fSMH8VdQ97HfAElkx+
oxTEZBxKVcnDBlPwHFuhJhkXsWq8xkBymhr8FDdV7bgffQdGYjx+3tkNeEQ0P0Be1Z6k0xN/y9Ay
uSJa1MB9dv6xstyMYqEPtXPnxZv0cS8XavHE+QItw1J4Bi15ovtpfxik6x0LTx7rIdcThNA+xmhx
oR36tvPBtY5wVWoWSZh32NDDRuI4XD4zs/IOjgfX7j0toRQSJmtWhnBkPzX0zK/pCKXEOMFRpeYO
+AcL13cQ4PkdGGBCgZhA85wIaE/wi4S8FmulT6xcyZAp9YCHE9aT/6gCvc7mdkb8sgkyp4175u9s
pKpGhsVRPFw99IwdfBXtlrUo2gwXurU75wWSvaRm19+ms6uRsYYgnm3yCGivrLFgx75bcYMVtCXh
fx6nIOLwUMsHJ72dpvA1or18zro4hNZbkzg1pLsM7u4TKCFJL8HECP7rD3DGLU4J+QztijceDR9R
1MA676gEIN3FOH+1xkjfK0Gn+LhhzBjEYKnpv5sG1xb2r9bFOZev/vNzWkUjlzv/qrAdnsXfxQLH
kTXARzh5+3Ird+9YsBLqiSpLYcsbkBmMX/chpgD3Q2zuQf2UgrpyW71nn8018BLh1jbYXVQ9gBPq
s3MBM4tXigc5MOJMUlCgptYTX09oTv2yPVdQ3+ChWLtIwwcuMVxl2u7MQwgiLMUXphQyhp5nBchb
NsAdjXSE0zHtC+cxGTKVT7OfT/Sxsta3GhI+2YajvVFcAu1GRdhgSnuxisjXxMgq/H+rd6Jrb3zF
ixgdmD0jkF3FmoLa7vrJJfEp/61Pl3/OPu5p6Diy0b5nB6Jr7bWGEEf1Gmjg0FmkcAVlhIDFAMze
/rE+h40PXsC0pAG3CRmBaLu/88wACz+ext/hqAulOLMDQ1NHGs8vDxD1yMH7eIgFoR77NNnos3fu
0B50ZSgDrFDP6Yz0m67Lo0x407PpEofHaf+mU6qoavWJH4QEwzjDXysmORhlZIvWdZlg8W1W7Jnc
UCoAbUBqmkRom6mAqk6ZjJyRVB6NUc5wND6ZxizZNB2WmhWnTHntkPf45QA4/XASLVgAzmP/3WIF
KpHj+amLvZm115+lpBZ2UYkjtcYr9cZApe9Lj7ZpmhUHOgpqdPsNQk1ShFVLSG1OD9SFLuiVBONw
oD2tE59J8habSBrnhnln90wavVKPDl/1vzIlmzjbcPC/F29bfKtfpSZj2aZHG20QyGMUWnq4Jt4m
zXZMgCweNH6NJ5VdrzGYSvRHcQXurRpI0306/k2GlX7FvpIRi30RDssWPru/6+q/3MQUSQ2nirb6
UHo9T/mYaCO179mQuvkM+tMX/7NUI7eEvWFhv9ok6U9I713xDyLbzvRekXGJqrO1JFtrl6AiDqPx
3b58hsvyfJrek6iJLuzEER5J5HrZNaU3K/jhU3e/L+LKTcop8ptalg0/okxs9cT8tM++aEA8d3jP
g/rIedweEwk199Pf6TU+qN1A/Q9W8WiyQHznmURM9+gekllzEwgAV4IoeW6x5Ei/KL/mi+kma0mU
eYyrqnGCmy2NjAUcRr5u7BBSj1IGi3TqYbPlRTGLijWuLHtnPKkqwIo23dgWOzrvMIZY5PUiVOon
031hR5xhkbSO0GRBSVofQv1QjycMWpuz2UDxxWUi366kElFgUUA+/OHcyl9NYbtWXOHHvIKAMDJB
7XJPzr67rNf8e3llart3vTayo7FfGpRxAe3BIwcfa1djMAr9cCcs/UJrCFvspqgOoMPvCa9xeSm/
4/jKNrZL3fanxylS5pl7w6QkR3/mGTq+Cja4i/CPvDilhUtS3ZvjCNOMnS7Gf1lcNTXYOAkSS6BT
/fYHasSi1G691jbKbbXV9mQzrcy0eAsAiSINZrGxf7VMZPNiSfE6t402owjF7B7nxdF6Bgbo+gRU
HYGyioGsMUT6ivXDZTQNgRdXzz7B3orI/vAOvfQ8j/tZBh9CcEdrmbW7K/W7CvbHiSf7N5OfHEIa
cNfPN3pinFaj2zCm1eXtVw9op5ByrnMVmwjj3pCqqsByj5REE7mHN6tIkCSWOYWHaKlHzbpyLZko
i9cNgrMennQDgakJDLizY2TgIjiWrZ8s9v5Adhc5DetaF9sfm8fSW3UTZTf4YyeMiYonPdFiETUG
Prw8FThD/Th8ygWKoyskXnMe9uPOHYq4Nx9aW4tuBOV650tG1gr5oj+kXfqGWoNb/Yo2mo6sfzrR
Sjeeg0DOQVTBHuLtqsuzkx5mT49g5OhjmYcGaQYGLik0OJVFFHe5HccxUErh3nxLLqqRhJ4a/tZk
rEjbsfnTvEzAEXdu4VsEm47KOBGjEV452vAGkHcbP1P59J/lYwHaXDkpHjUIjl1357k0oLsuqKis
412gbJuzNr9tA9is5MZTTYo3pqjIM7lhMW6gnwnEq0WorhM3p558sob/ZMQ1WaniRHH1XOY9twG1
eN1wVSPvpngvetc7Y6CzW7OO46HNViF2e+UWeh9NsockT651ueV0dh77AVjjHXBwQ3rxcR7yIAHs
UEpXWmmymEN+pjOo/E8OKQQnNRuCGvqfcFdqqA4k80ignCcFbZZFQXxkLS58rol4Da0b+UexrIaU
5fyq7l+O2XddORKoUlGcG6eu43oNXkJxnclwpgGvZDlOJO6lXG37Uo8l+wDAx6XuOr4washZfG/y
ZdG6iO541kVJp3XE9N5C9D5ikdv+KB19+o/BAklvbHQecYAyuz1azCd1IZUeSQUFqNQ8AA63Q+WQ
Vi8HIITY4eE42zw/Onbq2p9KdgZNAsn8OkcmL7cU4enUI8/s/04ABYHFHbWiXOuhAf0fNnqxPYZ4
EWhZk643rOhGWvS+umP1ZIPGkOsJ88SuqS17gua49FuOlUFuQSDOmoOJCvxYN2M6Ljtph21DHOqK
+IUFXIOHhwYGCH5o+L+d2xW2RUUoDtvdx8ydH+e07EDOVGbknGhcTqItN+gui0TNW6xHU6MnaWZW
+SF31dgedrReZaAoH4JDCQG9aBLm8hMbUDhkj3GtnkJUbmkl8v26XSlycy/Ro7i4/GDckAqUzHKq
s2l6bSjUnHFL+S2izUAiDumyH2LD4SkvR7F/6QnxUOilqnG51gm38CkxtlSMJhHVHXCUvnYEufzG
zs3WTGrSC7jc1eXVpHnTJwmjaReIuSaOQdkUP7yu+TJGIMSEO9PWITksA7UIEl/EHhEKHTBSly0B
MYgsMLbGT3nadcZy7mYKvoLqtsLUAuP11d8iBi/FavPrEPt25R1p+xfRZrboKP5bSLGstw15snhM
x3lmwoDiIN1iKTvdImHK9g+McJLam4jyffOrGkgaqJH/knkmcPsjrtu+U2OmPtKIYXfjkbs5olz/
UsxWVMHt5/EWB3kqK/02PUB6KWkG68kNvL6iVAUNI493PRME8b4P4sex7ddMfCkIVayItqxKAmVP
m9TZDIqOwQ7UvHlB60KHz5siqu0U44MyfaOtVXYhOvfnaohuhYAcc85vBtfhLUuUBBBQ7PBhzGhR
xUJj4Wi0D9UHTvhz4iCHvgIbKmIJCA6OeuLDFSv4mqAJma/I/v3ckIYdpsNxe9Q42Q7x6mZ7bJzB
cRa7lAg+PalfVm6zPMx+60uV1u5KP3zidRA1pxD1r+Mk3I62GcuGaRAhkD5Cvab6e/nKxAFMlPAB
o46DATGvn2Iq75+rpswv9Q94JmjyTYW4HKhlA4cBwady2bI4dM2AR4MdgEW+9mAGPLJCdAIx+qpq
1kR8UdPh3jKvZG9QYFZhrtZPVPTFNWxptcMkF40T6PVUpOUdUNEiEJh8E8UZ+OYDnGnR0bmM4mma
EFK4KzenDi84I3Q4+c74ShuV1nvt5K5hNndMUmhN5LQTLOX9TZH+f92LHw39SxTojnWHTYCRWyVM
vEVbVk4ROrTN2jPifZU8i7JWkwbz3OlOvpKAC7GvVEZKI+OJKCxoKUzOF9E2RXC/Scxzxi9RfTmm
H0EmWqWMANDUwCbraDIwXHSsy6VhP2oqBRl99PyPeX3Iuo0oNMkxwWlhmdprrziSCBwZ29IkEiC7
csQ1bwQLEkGnrUoj+/Gk/x/jTPmseTVZSK/l8eciUpbY1iseBNW4V/8puoisbvMEeakc1Fm2XPYr
+X6XPBkZd9CM4TtQMhKqDaFixwT7mPADqva7QlQlw/OayDEr43IqklqWVMgcC20nNKzrvxKfFnk+
/gs8fIzmL1Z/OC3R4xf0fykaA09hfxhmDXz1ZqMtntKEwQ+7m7kPNhqKfqGUbc8yvAQfU51jtnio
4fnU68yFNLZAo/mxE1WJ3UWw/UstwGcFAxiORy+1E/UBf4iokLHUQIEg/Zkk6BjiGj6kD4aKjymi
y+bnfMLlEjagng322ZrEZUdxv0AmyGnQOofd5uiMwtcb9CqpWtRmwmt0kOAbzel0EFpcaTXh7gQp
FpjRIa/Hia/PxlAqzB5aEvlOrr95Zd5Vss/y9XegMbuP4oOgsyHXC1sBuxEqc54RzKF4tmispar3
YHuet0iWD9zv/B/r4G4X0F0xnMaaH10QXU+2+ASEA+eyPieNrAyGMFvgnWLe+R+6kaT0hwHHWVKX
9jTinukkFt1QiRCo+kJA/DaO3Xuoe3ZtVxv2EUa4uq91Q12vUB7FwTWhmyE0duhkoWt2++ZppzGq
g0j34qjhyBYwnDHyAeuL50nrJHztYGU5uI/UMAKGazzLnSFauvaMeD1xG2YIQJS766xuY/cTIkc6
ThIW3lDX0Lt7fOtsL2nU0QP3P0DsXVSEdk2roqKoee6SRs7TaiHN8D6b72SwR7hFcv3uFUHavgJp
uLCtfoqo4RN96kIY44NAhp9MKKSIjjM4gKjq2veqUT+oLFJxSO+jD3i3t/Pnm6NgSefagSKT/+Y9
ukWv5Oj4LVdTTekI2MGygdfJ6Xqunj7Ht9yz8Zjl+5ZEBTqmKa7XDVSzicQIdnc4I7eNp3ABQj9w
+B2ltXIOpeEf070s4JK6EGz6Ah7vkAQOdhHB98kli1VC9UMjIXDD5un0fFZx4/puFk23Nv4uTRtX
P3euQtbCcFL/psRTPuAP2PCCFXP4ZarQA56Rgk/JLvt0i9G1iqIz5goZ2IkWUf9tR+mkFHCBXNim
kzDO82AAEqgGDIsFBDGtUqlC8NgEDRy8ImNxWXun0f517FHSQaHVA5QR5hKe1oel6RhsMkQEy23M
JAw/quex9NaJ8of9udCkMVWG9rM30OL16mEpkNxacFmKl1lrnhacls8C1WERsa7GqZ48Hwq3JiL/
UM+yHSzRzubaMqzPj1GOQDgz59gejA0KnqwqfMouihoapB+7fXACIu4jl3H1uDj/wP0cXd9ogTSM
LZV1PW18iygMQByib6AYLG8iuXXn7Jnp0/eiLb70TDZb5/8sj5ymwMm2EZBqwHeeEjNTQlorSghU
H90UuT1EVRztCqTuv2HlhPAgCfL7aTopPngixWJ/OOrZUZ33mGjQyoH+rI7kb+g/wDrx0eTrtHjG
o7oHDBB9eyzS5sza3KNHOYnA9rjpvC9PfDYEkyPDVuU6RmIh3lYjRB6PT3arNYQjwzG1qG1G9JHh
zxbPIgKFjwvweqVGTZfTjr+iVOwmgTxlHvbjRazxo4DIm25sUD7jPF2A+3hYloaNW59ppK+UX85O
Iw07TSjGKUAIvQcp2jqvBQzof9oHzMwC2LGVwvnc0i1PCXdtfl38wN+QifYZQAvBBA2ZCaDN2Z+M
woXNQU1WdTwlHkWN4LAWZ3hVmE7oJOAyoUYb2SzDhLYWqJRoUsvsbN648cIroc1aX9ZdRxWfN2cH
cv8vzobSfelZMfH+qrrlxqKuzagda+7ta56td95wZLI8bjnHEzgriAf3aNvYYUzo0iBz/c5Qn63f
l2wVGoSzQd7q+9U15m4EGazH9JxZB4RvsglMy+udxc/l5gjaF7q/vaAQT/gitFHisvEHHmWdRZM2
DlJheDP2dkBmLEBWPfrvk+Z8gDHvePrDttFeN9wdSq0ZVuEk7taaCkwUzFyxAyI+YYPu1OriCUdP
c1t3OfwG6L1iFfelebZTi1SSXxyE49LBDu5iDzEFKym52uGrjMCeMJMbB/K/iUISzN8jVIgBIQ3o
GXbXb0XE4/gu67SO/Ti70EUyb0HvNt/hcE7yhR357huJ+pqtP+UvzBcauUOScYIheXdYcIOsQyaV
ucVfZrHmjEBdLcgHy9BN5RD1vor9PLCF1qxwPAtV1YsprS4krL0aXsvi4qjekx+QuDtLkSn8Mj4M
jV2yyVL1/8zonp1LddB4VqoFDtjWQ40cnhmOwW9uLHrbt1O6MUEy+ptXI+4fwb0iyMuz4a13R4Nt
KwWnubnuzlcb62OqC4kBTZIXIx25MR01uhgBTD3my8IN8TrTtIx1Z9XFZOLt4d3pjg/hZigS5PbK
IDdlD+qZgpu+n9yfHJGt7YUwnq9Zmz544iqewtUTpzVJHJjFvkmjyB+kjoCbdQGMOod/u7o4vPDQ
AEPF2NjvlRx5xl9oweCmwLpmCO+mNnlCNdYgA0hYbI78AplL1a+Apk+jMkzlplne+Wwor5y6CQeP
Wbp2SbDEQE4r8Qt7/+Dh6nu9B1CdU+wiVzSlRPiPz7gRmNoXc+gF+s3ez53b45e9i4UxFKmvK04v
kUUV8adyBsxQxE63RoURprqj2SV8hDQt9UZNE5X0Yzis068VQxZkY64/wSW6aC63tLEb62RKoucM
YLyHVYuIIQRra2+928vOtu7iGxXXhpS5taz9QK4kSNCyJ+NZOe87GFtGmqt/ckwSupLaYzBgj46h
HAra0fKV8qHQz5zjBWr+USaOhoGabaqs9Jng6TMDeE0ldCaqEdMHn2qMzvnp7z0NLA23ars3/svB
7geOnDB1jt1p6PllfaGs72mO58kXSgXHkh0RQxd+EyRdzjExkFl3K3Xm24I8k37Iujk/qCf6uw8T
QjONYU2Oud2gZbFrELPL8/9l5660U/lszYMRExjbWsBrnG8E1y/w7FkZBQXwzXnokoSRh417PX/T
ebmScM880FqJLXdgbdGNHuF7ryGVdLnBrmRZ9W7pxVscvzAJy4aaXNKVClzVq9J0Ci7B/WP5PJCy
P91rTFxJH2kSQVptZvn76rIy49AN04fW90fZbLLu3M6vtCiezL7AlOavLqzosqvf5GJjSzCmsEmk
iCEi4nS/yuo6cvjg95BaZKZTxaBJiGSe5+yD+IT6FCJjHc9o+zLVQBqnHsSSPbJxp3fqzqYRggZA
Hepm2iRonPfTL0czXveG2yvzfujiFEKQRHeN5CFn0x4D1nHIt8dXZfBjdPJntTA6qsc8N5bhr7nk
rHlIYADGLBJQnSYYt7jbDH48+ntJoACPWgLCBnbpfk7tIBRON0ydQX/eh8M4hO0IBr2W4CVgSpL2
Ula51TRxgjlIcfyeosGQXxbzI9WNlvt3+H5g1aReZH19CZicH5f6xAzXzNX3XhcNPc69z6UrY90T
Gp1hSkB9zPrZGeVOaQmE70rNZ0MexSL6/xaRkhnKuAwTbusANTuuK6jYFEiJVknBMX28qDwIEllf
93S58mA0BbIjFJVo1fauIjYuF5cCEdQW9ZwjlU7z4N5TGdWp1SNEYVNsGNwatgGeKRufRO66r4iP
I2KJ3IdLIDyZFiS9nBCQR8L8UiW+I2U7HjcQg0DWw0Ecpb5S/q9YVUkk8qo6w+zLxn9JjPmJNqAn
0Drk3BohxjPFUYhRr4790zKtFcwqcXMHWoVvNeYq4cBLu5gTPrj3LapW4yiUSIw8NVP+0B1KeoNZ
x1r7XhM3ZZedX6EFLscdH+bMMQEIyT1UaBwStS4nVYPY0iDK9fD6xjWPHd2faFW4hL4/T3I9tUip
1oCFhR7Qkg6+XnWCEY+H5UcblxHMal2QFR7fwfTfaCqapuYAitxH/5shAzR9XEC+och40mZc4SGZ
WlowXc5GN8KCDkDwkOnMlRyocH/3BeJ4VZ4ylu40swItIFpX/rxuGIWDpaOO5RgdrM0YP2q3rfFM
vozTwUGGi1Gc+pH0jvVOpQmUbfgkIrAy+NqODgaVR7ZU/zfofSLkOnKndZKu2a0gDpTCCH+leb/i
N0je6irxiIm56/L1wzXitGL/97+8P5apw9HbD83Le86epTCvrmKRex347ecxaZajrxlui5G7ybVl
uHQjuuEZWOH0GAHtUrDFideQbE0puYlfRhuzcXi4H/EEsZ+m9rx9OU/7vyAQvoN17ETdCGkv0OoG
x0Cv9hTrn+Bk9zoI376oKHr3eTFMPFzm0buEmLsFuU/wHwnAiaty+S4SJeS5ZjDm8++t33ohcf7l
yXzDSRhuWJLINUiV/trT93f8/ANS5mZ7c9tmIs3ETR7Ve+0URzaKSflwmytDFPqxLLshwj85vXXN
6BV/tKFceiWsDFvuAqk6rJxnNYoymk70qvzYcFPctch8zGZHIy5pcUhXLVuyBSgkgREVnmI9oJsH
ngUj2sfXYP00Muj4h2DY2vYCmHYUrktsV0qhpVU7udrarLLteG6JQfg7x4nsvPel5VneQNDXIbo0
8F/fRFzmTXwelkZSwsPI6E+p7/RQ1zy0qxM+edTGsGSx8sJmbZvKy8S02c5a/g53TqrI3eAqNj4l
LqR47XC161L+NotOyL67kkpFCqCSSltlL8W2tEd1m+U2zPut6gTOojI5hPcL8lSV2uQpQ2806hto
tAsnsoCek67fWxNjsoRwOIWUBwTI0pV1FfEymURkx41+c1RbNOwuyPWhKAbovOD4UaNQmEBkweQm
vZR10jsS20bCMweEVrASN4hhsmImOube+X8Rj0xVsXH+074C8StJ1mzNgILF8V/gFvhUWxYE7myX
HM1g2J7xDQpeW0mgnPpfVkiV/RhlcA5MIXiDK+8/U/0LQMiRZq4RHxbvFjocOySD4t2Lfw4tnIR2
bykRq1z6p8qwRY84JWkRqP/uIQ2qtuFXQZma48aRS7zoNltd5TX44QG5oB+Iw9u75yhIoQul2Lf0
qFYSqj+G8y1hU9Xch/n77kSANnyZcM2E97HWwG/N4HcpBCLz35Tg7t4lIndB7m40Wga0bomznSgY
U8rIssEcSHiQLXgdGQ1cQPIAEtLjwa1t+PCeFGEX90iOcg7qzjeUx06OVZJVbxZsYaTs3kQkzxoA
AyG6e8fOcXMsqzJhInSzHSkemvTF70HyQhh3+GsbnCDWS5aMmmJPqyhcqRJubp0fqWF8FxpmuNKw
N7mvIWi3feMs4D4X0Zrpmp8RJkyczXmrGPBouP8OB2v/Z+eUoUgxBE2Don5zeWQxOo9UtQCa9z2+
xgWvi9nul65ZPWIQN/9QiQSPPRFIqzPaiAhvLj4lkbbpMUH7oxSIB6AuzACtCJVTqEdvHv4KrAPo
KSAewWLvufddTm7Qf9kNvuU5hvpDAQRUj5XZYLX22hZkY9/UrS3XUkzEeP0+RHxBopogIl6Impm/
OzlRfY+LnYSz7qZlJEteyw5aJ29i+CyzUXnHaGqd0CW4jYkUfrFZEjDTl/Cg/Kilywhdbg5CprR7
K3sqiPab5h8qzexuVLXN0VsZM/PtlHbzULb7OFJVPZSdfbFWR+za2hphbyadB1druU4RB6QwXhYN
pg2ek/vHgCqms5168OUB7eb/Wnk5t9nHbx1/b+BBqmSc0XDle4sxruNUHcFeB8WhS5El4+ftmXVF
JeqeDFimFxDep413eSOX5HxSosqOfiQW8TUGCaUidT3jlgYezeju7fKUOjmJdiLc2VpZgeZlY5zC
7Q8L1+JbrPfJqg6ee83LwzM/1bmgD7Z2XSjFpWN123nhC80XFiWRUYIoVMXysXcgG+VJEtAoNc0S
CpCCTk8KJdNq2xzZn6Cp4r5PAx6zztHUfjdlh6ogGZH12UgqBVbauWWsHtpTCbZbfC8m2YJaU1g6
AM24JND8b4anyY2zZXLBOEk+3HcSJKXKtxl7UJimyMttibi1lb3eKfC02t0vB8ifnH3BlxVpOtp7
DUmQVP46u3OsFeVFuLyRryaDU2jGcSWOEFOxSBZBcY7ebaurN0EvmQAHc6D92sYgKlKrXfH2VglD
zw67amo9tHARqYqYrZeSqxFE4/Nkj7bSarhu0LTEw5e/AfTzgyghTMSgN8SXkZpB7jmcqe485kGJ
wS143vSdeNBrM7NrchxX1UdVoIW2MxQFlr1jHJELYPp7eILXa7btnCuJn/zWRHuMIf0bnKeRmeSF
lkD9y5HxOh4T3Ys0pfTzH8DVy2cVu/1oecQb1Ierz+kGxyPedvT8UXExRE/iM+wajo1ETJ5qdls7
H0zCj18DuJOGgY6eWgh4c6uamHyh9v2TKd4fZjAR7ALUQpQPVzlo1lDP4OP+BE5a6VWDMyNyNdaT
e2tWIW3JqfXV55hpYGvNAZHV9PY3eqbAR0OZPhbcIQxUvGtd985ViOqEK/SQRFjKwdwsk4l8XgI5
YGK+GMfzF30AQX9LA0JNmuTuWBtcutTnqgn54ul7eRsXvwaXjjoX5adRH0v25tygQmmWjHCozYfz
EqNGbgTO4F2T7DJbxQAyeQarxaa8TvoiZ1EIuhEuS15zSzegsNGr0Xn8ke/dj7NJrWOCFAmJRhoR
CUF/lyz9SgtBZudUYAGiYtQMWLNRgXQNZCc5bPsIIIqQm8cQmGvRjQeo0xOzvO6tB81MzTp0ToYs
edH19wOUOt+/aNvuSs+Rq3rT5MyYFGIs+ogMPI/SnWWN4JDj15BYxYnRvS6xZWYSXfirwxmSqvMg
XIdQRIHrGnH4ehl7ZfD4Zk/l2+QIgcq+RADnIrtBcsZP1a+3tqd2y7n9KhAP74VDhcLx1lVlXngy
XjLK3y8Y899roVCKyLvle+YWHIEpzxo4IZqpRKInh+Ukdg4BF8FFuYsbhEozcuHoRC2EpgfYR2S/
4S+XK6/m+Fi40sH4I5AymX4INEiBdko4V5kqphEpqjEuOzm8HaI4xKyuoWgSVRm5LfHdaaOY73Si
8g3mk7Ey6VWjkV5ADG29ca4BJGShBTi95nTzLiTJBjS6lBCc659HW7ZSAlsh0iQHRtcJE3/f/5xr
9wfJs7rVNyV0IuA7yR96NMGNupYkRSQI+jod+c3klYYs0On9emSG2lVkE/xqw/Wv0tH3KrTVeh7D
UyzcHV5Nl8JSIkf3KVO25FHc0BWLJWhFIVZvTNJyIL7lI6iquqyllT3l7nmE5DVHQaWQ39di7iJN
/FFXne19BwqV6n5J120lirEY4achjiZgNW8qJkql1sKrSm0dlE5N6tDbrFeaPBSru5SEb7uGGW4t
Hx2/4BPfAhegCfYlDYnJk4a1XR9kjB4DnB4ppGkL188CSsAjgKyJXz0XbQMmz5TQYb9VNTcdxUrj
yNFr0vTECQjUCBTklyJw6uqlahLHkinFvntjNlUXPeQNH/WprgWn98MrC/AfMXiXEI+q02tLZ2Ta
7FWHfLJ36KSKEYvCDoZKrJbJ8ckIaJgTsIyKkrsMXXmeYkOt1sJ4++7cO+njImtMq7my1zWBDbNW
ethJ4Q0JbhlpQG20FW6po18agKr0brp02zpn+ZoZZJ/kzq0lriokGc5HKUvgBr1A0MYlURzlw7lH
KQGrl5o9QkAdwumSStqhg0wguGhsUbCtXJnfPWsqy+kg8EM1OUH/u0QWJwrw1jpR/ezOCRPlyaq7
B1YBLJch3IKQ4fOK+LibxlCXEzk5c+hBLyFr0T/EgNMMZ5EjlClHuYgJ7SxVbS8bEYRvF+ILcIcO
8P1cs8VrO78pNwj/qzE2xdP/+WXAGHZBtZj875GC8jetByvh0cF/VXr/tMY2d+Un9tDiDIrsDXGK
vY+qV36kSpY5HBol4JBFIX0CgaY7MlGwSAKtbuxIMa9MMjLgy5qwtcAVQJC+zu/dr1+ZwIhoQwqC
l4nY9EIuaBV7KhNajVtsEWA8qof4b9yIZLcm/XRNAn/7/LfFR4PuCLe8MNWLW370ARhAffrcJhsE
Ep5oxvoyJxwh1jGMuBkAS0iY2Kd+DE8V7cBJ0py9OqkQZf0X/8pgcZzvOjLFtvIBYoFJMxlTBKD9
viUqPWzBeXVBUJhqmDSVgF9hputkXCDlVQY80/tbLcFIrbg8o7F2g7/1vVHy/5PiiSJ5CAgg8/eu
ZOqRrfpjchHltk9QCtKOVkXwl/euTJhjNOmTHNEqpdsHr58apZICJWTqD1mcl9pIWtpCEEB7oF3B
wjJzr6taP+puZGR1GcYTes41TDBIhv395NQ/K8TFJkD7E3WcT9qwOtLNtlcyLx9CB2JrCmAtoevv
sZh6QIEJR0fH4pK5mlt03yurZ3kOgwlQNUwlgEqx0EJEJLIQK2RTHS4OlNZwswsoQ6iZjmdCgO1j
ei91Hu1lcTkbSr4nWM/gshul1N6UQLfpXF6tBDgzcfrRM3GXjHQH1Tjd9p1CGCapkO4InO6+XnNt
cuj/Y8ee0/uzlKfkSDlGdovwzKb18agFcPRUixWK4qA9ON0wBX5Oz0WiZAdS9V8q6vTOzd9wQ6Jy
umgpWydaNUZi/j571M06criqGATDE5KMdyDGsaggXOQihAhkiwJDjL98Xh2KpIAyaRxoLJ5saq02
2W8MXRTxmI6an1yXk5KI5iRVAoZmvUZpeuqhmPK1YNV9WkTtKkuPF0dvYinyGIJ4lsmu6Dgr7U4O
eidhKkyZOeCKnWSpKYBMTAsIHMP7nKmUGRjF5OaaFHUnAwllbQWc7UuJ+fPuvH8uOTvaOEj2xfF8
QYpwMrEPVqAOXAECqBPkZPsG2iaYfJ7g0X4TKpC6IolOSiN4PI8jBj346aEEy/cdjA8cCBw+tyS3
3cjGQKa/TSIeeS6N4ijv0v+YRR5j/yHR5bIZNrMPfmLaDY1x1mVbbuqeQowWzUcjI/74UMKT8yvZ
4cvJ8aqgQ883n1NVDrfhC5ueJGGM+uYv4oslRjemCNYhPxmRB0J7aSw62W2p0uZzDTQy4HSMArYa
nPGpjCDaXVBpO2y6NhNKgbcx5DtXfyoq1FXqvTfG31lD4oiESGhuEAYfeReTYzRp1pYKhka0i067
HQVoL5apacDkyUB1r8eZj3NePdNanSfyPuUW5+ZJbdAuqBQ7mXep9oCIQq6fobWKF8gPHbTrFA12
MIGW6u3IApPjou3MdbAqiTLWD2q5Uou/wEsNwZDJs7I4/auGbvO3nSd9NPY9Fm8psv/kNnlQUuGL
Q5dVWDRKA4O5FZZukK9Ld+XlwF0abj84yR1xWYTQ7+tcxurYo1uInYsiP06zpniWf2wyBUiutxWE
qTNd/ZZ36/JAVLfq34PV75ijMZd84rjT6ujKp8dGlV2mSJAGoer0I4F790L0Jhsl91O0Zt5+Lrjv
pJlUqIeWEl2G6HryVbKXLNCdJEYey16QWFOpGz/wB53UhAbp7aDwjZhZxIEeJrrwfqev1L08YsqP
Xgw66T76EVTz+5XBxidZJuQt5wobIW0SZWjb59tYd7NuMFXlk+PmHXHJRqEBgV+c5XrUtG8pjQFz
NkhRRxqeupCWRkTs09uK2eooKtLVQSIv2IiW7Sh6TrTqJIuHH85SYeyu20NtFG1Y0eqAIvQElxFF
P/cNCoZLoHyVNjBm8M1H5NHlLRc8TiQbeY0SJnbK8X3rd25d8COUY8Bl9Zh7BEjcTokfdo3osh6g
/1WVvA3EKXbuULEhCFZsL7zg8fj98tCE2zGA+z9vH3J5C9Pxo8Gub3gSPMYE8kQ0qIn40hSInf69
IheI1bHztqXAhlTJDlN5Og5xbt5yYPihDs9vcbZEv0YqaI9vWPHXu/yUjBy6N7X40/zSdtzGbzfM
+niVBJ5GzpBO2FEqTquwVwqAe6Irqn51QdXypn4AsENLvSBzt4ENBAOPx3uO8a4SV1HluhubdX39
KI6H1Et87dTZ97R+KzBwzlizEuiuyfSZxm5YKsuQ1zc4zHMLwcK4M7yBu2RDAMGaK+ARDrImllb7
Qeaj55EmURbXP4LvppGe8VHHFRDs55gF8cNdlBPWLlkDhqPNPpwfuZWx8bZq7dfezLzYpTOxlY3m
mYsPXzdL+Hn4+D+ZajaH445nYN8+g0lTWF+twY4W5eZ2qpQ6NfbaruFcZnLIMcYT2gJZWRODcpRX
TgT9MAfUdri7YMQO6ZUXsSES/6eMVW+YHK6aBASlWW84iSntNFKM2SfuIOtFAC4Juu00VnSHoNxB
kFW/xSPooVLxuCu+dE65k3IO3DE/wsn4SijlqI9C9lJLxqDosGHY6utI/RQWI/K9L+RNFmPZXfCa
eMqkYThfdvbxB7JVz5BvBqJ3nyXY9z2S23DKTmA2jfXUzq144d/AStHJ57tDHt8eqiSiSaZ08gZg
QNjzyi3Tm9McMhl+GJs8BbTwgVB2SYUNB6yz4eMG5H4ulEkOcoGnUbubdN8rWBtm3Sz9SfRmDGK6
yyHq415orParNk44JKv4cz0iZTmm/qij0F2O3HK6CuWgMW4mYBWTh8KY3ZVC9o1cJ5uFyDUuS0Eb
y1xnT4ZizMGcgkV+xg5rCiPPJpJ88O2T5aLq2LIH8eYJL0Z2lp/YESk7+w2L5pOyTJhXXn2HaLBX
bs0XDicqJ2E+nyCqsCqasesBA7CXKmwySqXb48eMs9Xr0Yb/X4Tf7n78bM2JUZOUkZgwzEXWSiXb
J9sQzpPTUDz/HoUMSfOJzsvmVja4z5CR8THETYHnNefAaaiAMvlv2D5TvB/XTB/8V0rIxMyu7J5J
OIrEnYoktyVZeTHC/vZdAcP1npqJlwTt3egeRUUPeZoza+3AHpNiJUPAcY5ZwpXVVfHDcMp7qPmd
ZH938CgnqZ5jpzCXZAndJpNyU1HgXP2gPLd6wQieHtaxvqAOMeNrGdPdw6y7fx+6GSYvoOmSicWK
zbc7B2pXCQgSh80saS/QMc7rfKZWAs9+svX9FoAd4xg9vo/ZiQN98ZeRIuF3jqTcR1NAq6CBmXVx
obsoucS1jTQkxzFjB3SNE35yUvPUtTB31aVXHdsTc560toAaTFJr4vPqbJWSgGVkMbzrcRtrBweZ
9A+WGGpn+my8DIL9n12ljZyYGh/nWnEvdlL+4CJz4YMEmzJLGx9p1jz5GqF6JySfzb+PIGviK4c3
W4wIH/zoN0LG9gIWt12FomwKN9tZRoXrB2AutbRbcIbp0GBA72VgzuO0ht38hSV7IiXW8H46zP2D
xIMjs/bTQRCQu49iA8KqARklDuXKYpu3oRLsPlLdH18QieKPInR7qyulxJQlFTeOy0dlmAOk8yWt
pMOi5wydwLkmMqyQUwPMugauQYHu2E6BdjJA5954yKu7SLfibSl7NDrV058MveAK0C4pb81tTZ8O
kxYK0rSIeNxBi1ksFasFExe+f80o3QS6e1psPqXvH2zUhvDEDi+mt/GbjbQ1kuinvlP9UsucNnu6
qOB9HxOXxorsIUfmniuz+m7JNCAIK4glKT/jFj+cwG3d+jpVAVY74q+uKxzIDJIzNFYP6lk2vaEv
0ujVSW2FfrZyADJtrU1zJHK02u/tjShF96WaBK2/IZymfy0UesGthp7PUWzF5sA02oy6iHnPMGL1
jos/IUgcU1W9orRTN0YyVL9LrCQE15Qk+A9C++y9UPTWs+3oa776JRBK6ceDEka4SiEJJCfeOdmk
NgAdtBua+WsOCCYr4hmCqVb/xtj/HscmNwNRnf/U5Ur0O18vowNHP335AfOt5anzmHeR0QZLNuAz
AmpxaFOikJC+Tqi2CoLcOsHQW6nTsNPHcq5uqMCsnNDlDBlwSBdkWfPAgS5X6luJeRMCQT9Hlkpz
J+dJqJzJfolEZiEPUHq0HpZ+7KJyC1YA4KbwMyR2uHUD/xwMowBN4KUGpGgTar3pUuGCkMz/3kJG
0y7XC4Np4xKvfYcGF+O/Ir4gZavTjCWsCxx1B60ZBHNfAVHXlZwJcrdonXE1PXI7UK4PSriHC4f9
y4qGUI6ho1e6rRwmon2YaZiW2sBU/611qCai9DoSQa9VTD8bko4k3UChZqouT39vDRvyztP9OShs
qa3tWSnsVt+yM5LEYDcHXvewB/d4pbloW4vM7uzVevImkzwFOEpvY7FsAF/JaI9JPqMjKH0Xp5t/
sGKe8iHQlMxHP8C/qVhF1084GyE/mXe0bhDcPZm3BUcqnSjhNf+TlK0+EE+Puj6TaPhoLrW3CjDO
DpRQd0FrOz45t3P1hNyhFMr1tR5TG7E3uaYq5A98sP5o5s/tDeeyhNxUVhok7JNyP0oKsQg+lrvr
oDCBd1jdb7W6twdoji+xjMMVPPuGOaOQJ+TON7WULecPCmNwfPtHXFkTEv7cijrJacZwNeIpVM6p
27/1BgxXykO44+7lvI9iWFscgKaSJbwo0YCFD3BFFxIzXv3jfNwSHHNqT8bGBkJJXzMny0nIV+75
OoDf7lsLEuxWTfIHj4ffdBv82fpS+LvfDEWHMP3G+wWFHVOD4OlHiOxJcUZLogCD59d7wB6rhJ0H
r2eoz7aFYeLzalAePX0fGrBz5VLTkuiEWz/KaffnhmobZ9aYftWdK7ZOs3pHhakeCM7NJJJ+sag2
g9oIwMxGOhZWV3XvA9E3H+eB/vuxx/6OMk7kpv8X9/c78ztabOwdOHyg/TesKerzb7Das/uKL/el
sUwaIPLXmdWhZ69psZXlTHUVumME0/cRL5GQZBifa0x00RQw/chVjo88AC/bB2Wv3l0dJo6+6gnG
7WAV4aZB2QXYetLvAF7y6mR0/2m3QY2Xd/PQyhkUwvYjx9L8fa2NCmExT6v7kGFeIyqqMDfHZ8OZ
GhKqIWGLGJo2bIB1Qahe2HMAWPbrka5naiTwEfkdyn5F5IUa/RxebTBnhT2+MDwT+XY4nHjzEbkR
bp08dlFQAAks9pwEZBq2GBzQJKJYKUkIcjsUs55Tw6BcTfEsiUR2lfIhUu+Oizi6ZmevCvZxFh7M
R6CE29slfQ2a4YCJ02DpeXjs2gzTL/RjBmjb8Wf7VTpfxzt0u7rLJDXGEmTRGiyfzFELzJwdpQCv
llFgbbq91Dlf8f3dAyegMYWoOLBOHou0MdhIQMzPPf9a0h2ieloZ1GWu0NzrzW/ShopjxSbSl8Dz
bgdeKm0mmv1OvDfGBhTiHeP2MV6pTF8I9O+xnk56+GpSuLYw2yOvXmHjQZezWAUik8+iKjIXC945
UF1H3930V0s9ENKmos9jPUlEssY0xOqfAAw545KeHTORkvW4EucEpN2uCCis897ncwZmEVwGPaur
gysMOyFG2VEUNLGjLJ8Vs9vKCZAlJziXkQL1bFcTpymjyU9q+9G0WPitrz2iV6IYgZqpyY/XgQBi
ofAruiR+w6gS2X1okAc8R6fRyT8McF/vS7feq4LqT8R5Eg++zuALVILYIyVu5W2Y3KDokH41aopX
eh9EkbEHnsZ0a+Nn+aG2MEr8BI1ikL00ctsKM1WBkV/g/ABVfhlpO4rgV8h4rBIrgz+0bRM4EMqj
u7Bu9sXZyu1jFc0iMhf9hFIJYDlrJasmCWgRa0paslFuoqzO5FifSz+1agtPI4Iy17Cx+IDEp5cK
IKKSSL44j5MIH8W6CO5jjr0cqjInFI76FHUFNrtprbit+GFr76j67lN++Oe5AkTt1Q27wXeZC60a
4DtBxotbAjsmV6bRkqsDdMlg8lpeptuXUtZE1+Kd/srRciBvyE1x9CSXs9wCswC+ulmRkZrsJoBE
h00+PUZFd8s9ONha2ZKpZDi3roeKV4GV3yF9iijmWRV2lcXWYZ8dX5lesjnpbEyPuGpNaOGDO9tg
I9Kw2udyTnNwn94qEDdp+YQOo0RCdlxTR8+L+7x/+FeM0g+Ym6GnudQmzVWd5GZ/RL9aCiWOXnw0
mME1TArw+o91D1piRh2vHJjatvZzwSG+QwxDKktGfFUNtt6U15vZhIn+V3h3ZNxTXIq4YoH1+6ZL
Gy2nn42i+rg4JyQFpL502H0M5BUpV8BiqFmojKENvFJrfuBTpWkYAjNryG3zmWppXjGaanKdCkvm
xv8jG0l0FGiBZRymfEC6EV2g3KoSntBiFvbEZfy/TkqYUcttKBbJE0KG3rnQJ2l42n9hFn3Grd/N
iGnPQq64C6GPVAxeIhEGFvWIDDyh9VT8kED45GM9kwQRLYbOLvhjaJKcqGeI9alLie/Y9VeT8btA
EiBpX8jFtQFdwwCfzkBR1OalJjSIHJwPoecl27BRpOWDbSjJTxtgEAjRpCAE9PA5Thv+mQ2vO77b
kyLvqafW/vwul5txV70ZXSKQa2IT5N7kqD6oKYgUleMLgnhVa4SAvoUYHT4MgyaYaNzapVV5n7RM
gG94eE7lbGJ7eD3sJMuZ7SJS0avsj0/EzbnUbjhAHCHgxd9uELMPVU1GJNGHJnqWjgms8fg4NaOO
18DSnaQF6YY0fLJjmlMQv6GyuLeafJyO7/QHrFE+t8QhqgLwVDR7I6q9N7DITpWGR+DLbeGC+EYi
KUoYQYgKc+apEINDj8RvDC3P9/WAW93+u+SHGdmoeMmH+52Pb5608Vhqk5ULO7H+1pxbyM7So8LU
ILcBR9ulbZmTGFBuv+0vJJ8Ib5MPISXGCOEMUFBO7JPMq4fPeB8848ALLrl6gcvrGJSvpnJOL7Wg
xF7HX61XM0gG0dqgBno0W5F+jfjgk27m19+Dzcw7WLzKKGisdRaVcQ9O0W7nxxW0maWN6OfWJFaJ
kT1CrWceMg+ecg2aYWYdWWgzMh+wZ82d+syVyNY/WjMkw1zfksHRf0uuMwURFZ8ySZJ8u2OtMJJS
94dZForKgDbX9qymqyllLIcBn4wLFAXgNVt/P/H7lE6FweQQG1APSxNiYLC0WsMahZ4NGOnEoqMs
YQjs6PFOqZfY8NTXm1jopXXIDQs++b8TBiu3iVgiFBrU/BJMsLSqK8MYr+OLVPhbBfJnNioMbFCU
8r7m/Smjpl0ktmWAE14SKU4LTxGBeDhY1C+LFZSk7wP44/hrxDbEdIEKi1pZrijPIxXwQBgRiAft
USd0dc04W2HeQTWmMKIbAfYpbD96pibLSWm7E6FsrpKGyWK2utKXzn0LG6Kz3Nln7Zpk+w5fg9sW
0EiEwlrh0izuYkJNGfAvJM/acKDVhUNAIbRJjTGxab0RmPyWTfjVDutNhpENXDjUJaWeKpEu2lt6
yXirJsOMgtsJ2T3RCgCXZeBr7TGCP7zLlZQv/35Hfk7St3L8Gelx2cyonFyA976vgtJkyLN6FTUc
l5y0ohQPRDzo0eB/U4BFygEGh4r0C+g7BtV/ggojoBRBuptpRX0cdGV6nmg7icIH9+i115/4utXP
q9lrwBDXhMRsiMVcQCushbwQC3fcyzFot+CF9K+vQiM+wWS7kDgx+cjZ5dm8cMIAxUBhhkEGlkUB
tNNCdDFBVAuCYb8ZbiR19N20SQcaW4tpwcYOHyHwajp0hcqz1Y/x79ElOiaoX//sPvigCzalg6Ta
PDvFC1i3i8fQGfhUb7sXCwyJuIdJK+92+eC07fwfW0kfQTeN/MVl6OLcP3NsPfKbX/Vh0+fa0HsZ
TqK16no4rluW7+ubPtDIYKdCi+SvGrg5QYLyzFl4xRuhIXc+pXRK+z8tD8c/124Qfj2os61XVwKv
ES/x1gN7B3Bi/fzqxqBhwX/ol3XTibp0h+wPBbkBjdRN3UudOY/eicWNZlizbHy0N8674a38JJln
5BmNFJScC5KWL2+9PIztChK1w5hy6jwj7Xm8axd25tLl118XOjFvQZz8+WV40nvYfGPqEU8gf1gV
/++MTSGt6gmjqGaRaabTeIATE8bAvYnNGS7NVnl+oifryuzs413BWiXPB6JvSiqsYAcTtoj0a6Sk
RuWVsBAi+qp88bS/RAyCSmk2laoHcF7Q+VCdZ4b2d3Ge/K2Be78A1X6bEmMstqxDoT6rNXEmc7Y7
55ATgXivLktAE9xu5uaDKjN12cnQOMf2LD+0TqCWvCvcPOsMoCminEwyOTf4MutKLEc9R0uoiDoR
yyjfTwhixP/rN2JtfW4aGy6gVFlazLqV45gTLqdWeSzMx8fu7Xz4q+4ad4s7lzRqByrTaSaTzWck
PPGZigGA7HfE9zW2RI08v7R6VFKJL7Py0/Nv0IvyA2sHWXxOoueY2shh9rcx4sKsieidgBaCxsrF
tz9WpnY/OBuQ3KVC5YQEa+nsk7krFqWrRjg69kfiTvZG0IF5HAlrGc9Fr6GCjZNt5PmtcAWul6LV
2lxN4v3HzLHJHLRkTAhFexGOWaLoaYp5cUNZsb7m73Wj0hNWxi5PnQ/g2k8+E0iyBd50XWMa9ShI
UrvyKc3P6SbQuf/Qp0HnLsAslJXlSDNipldC1XQFKULWH5mrJSb437nM9fDXEc9HoJ37sHHVOsSy
auab1rvgSgiPAD8kwIhHSGJvMKZyHRmMQUmhR+hfsbR7Y/mjExq4BUqvXFXkLtyFnXZzdR4tyOaM
8u720l4nKiwzvTtHlr/qdoqGpj7/huyB41WV1R/7a4bE8E1q54X0cC1OWBxMZM2jKz04uBjHLoE/
Xje2nKbwXVFgitHmGHb+bO+A8AVmfClsaSmqfftc2igfuSCSeK1e9tPk+p+Qw3as6+zYnpQT10vF
Ncy1wfTpGeH2wMIMVxSoeEn7I3n9rK6PI+8WXsK3rSuW+JR9h9L/6mlEx44cb/Z6YLcI8AMS/Hc/
/KRm1TmuCnX9Y9anJYlCGbCe1xI9DLOpp19ddK/xGBmRGOZuKSkCS+ZEt9I1de7sxoRdXWxrhgDR
ZapDogQNIY2e8kW78F94jg6Gai461jVJcbAoE8aNVSv8/w+QESvaU4OzJbBo/l6+mGWgN4Dun8Wj
BjyQmzxVFY0y1Fh0whFvviKMorGaDu28bcB2lKusW3/9gYthz4BUliL6cU8Ui7+Yz6EcoGJE26/5
sz5AaRFgVZtqVpx/9JufHtJS7+Ve9IJi2TkqOCLr6amau2TWvKe1QEjP1G3FjbYDsITIs6tDhgW0
vV90cMLg0z4KcQ9x/dUgZk9P1owOKGHvyUMxEDBSWpc1inHN2wPVtQyfAnogLebJjiEXrONeaIHo
7KYjJCmn/VNCahhFsdSp/WVuL9DezEWCm9k8+IqxVwIPwSL6rEUBHeCupcvzVp8ydvtOstowKF2U
htdPmU2N3YfK2qmgIdCbonpgJ+5W14L70baXpvGlx77x6SfhwOjVBx+sH4dZUWk7cYxJwoeGU8im
WESXvccZzZ0NiyGesSI7poy7OHeWD+6LZqhYDINJxoYZL0pU1bG4Kcta8uPlDSIae9TUVUNCoYhI
jUFBb6UKOsR8tkG6D5tKaOD83Sn0AWDNa7Cso4Ki9+BHqYeZnMD2KJ1Q8uTQro6GkxQ9cM22vKCq
03TEwtBhVRinOYWJDeUrjRXe1SWfvSL2wivXQTX2sgUHUmb7IHwq2Udl+X4EGq1j1kJcTXASz33r
QpMGYUkuKbm4ycn61XtnpwH90kD1aEXW8qeLWxM++Poq+y0zLX97aqHoZ8r464xwkPQ6kD1zJ4jJ
StDmEB3+mWlS27DdgMfqd7ZWWkPMM0MrLuCxVQc+adeVcLCkyrnhz4Z9+W061ebBQC6PjII+LMLy
pqT7U3+mEdFOsyBTVg1/d0dj60KZih0vw4TAdljdu3p+GhzTKpb6k4FDRJGBqZOrBRAzSpYjF437
relYgkBXGbCq9Z+gy0lDKazbVfcC8JHQG3rsLnvRxGYv10GISlg0I4AcDpQSkYNsaHp8n2CeFqzd
POX98XY9z2d/RJ0lF60zVjw1MwlcW50xVKw9j5YxhQjLxdgr1puPVZOQ3Htk6gNBIhCf9Zmp4uAD
Ga92PJch0wr6ktjkUtfIcSFPWsQ5vnGMHj1Sk4zTRw0KgKdPkOpCznQGpA+gLJxGZqOhKcN4n0OA
j4QQKuz+nQiUgujupH+fSxqV6uUzGAmH0yU6n/o9d13hsFkpQcBAncaAEwGltfC/zdT8cHX3lWEv
F42JGoVTMM7SFF4vDHUSVS5NM3LPF3INjJW1yFgVr1hea6SVSkrSqNkcGYSVg+rB4JnHoyrczJxr
a0hSiToK2ZhOMhIsU8apZ5ah2vTbRPfz5We4DwQkcedmTcKL5zivyAal8/4lgn/kok8RM7/KNyPs
2MrLPmr2NuTdPta87nw391RzXWlKdLSqXw4vUFXdrLk6GoDXXJ33TQqZ79gA/GHZNUaafUfRiqOt
dyGDCguWstIIz9UXa8juodeHz5lnzmqwtHetdix1uhsSfhZQTiQ94eT+jcJ2HMNkCihNzONSY/Gn
zkn7qK2kd7UktuqqImzJqhXLLuf53eYx3SV2OXPtaLRRiYuhU+iKnKdzED8FQ5Df5t2VQNSb/xcS
EwtjKkiuee/9K9Tp2rJ49q7k8pf2XnmZzwvEO3ba29/ZWGscGlHNwCzugOqnJ8znNmqoe/nNjizF
uWJJn5eq/mvK21RsxpMbzgnwQBX6ONAuTKtYw1+XCSOf9i2vsuRKrh4k5R0fTSWzYNNYHp/QLnat
oDo49TJ51uP0vpzB8eXP3VXJXiiVwFKgNFTKUvQUaEqilrDVegfTzDgnWofvIzVZ6SIqWU62ecu9
B/1CP6/pOqQn9O33KoqB+ymj1Xbl9CQj87rRfe//8JEzpdoquPbdlKD1jXltxDlUO4Lq2U1jS1rq
e4SJRLrhsGpdie3H0tJPGcsI/e9P0p3clJaCQapPCZKraPVUhXCZ6DLabLQ18vq3k5VoEMqy1Xag
csD8O5jZ9yAv7jvDHXx7twwvcWTbnRooTD5Q5NE1nnRCLBMcAL0RqZLoIiWzUO3GYb2TPjlGv6UL
Ws/ocBVWiJ3CyT3cON6rj05lmdyQzwuNqWkYyUhDLGqLt3GBO1/se/h7vOfQV6uWXoBwZiw8eQFK
3Y6hb0bevfVEBcj17bRekdMDXt1IC+o6deW64aRf0hHwErrl6qsh2YwFhkqdvx3UJfzuaG1z6vRM
xHab17E73oKhRD2rEMmODgWjwMPSjq1LZxy4ixtyCvOzOmn7rUknseFwH5jU4J45LJJfyMQbauYH
/MqXuLsgJ9GZMi/eZzyYImdCaXi6Rr0S9dpZQuCZbgvj9QEeAOV3UkX+Wv0sDLY/UFCBLFWSx/Wr
LggeA5AfOwuLc7LvVFTM0BoC5++Sdga49EJ6nbW4ymg5AypsHnUZzrHjQwidpW+mzhy+Qn9Vt68e
6ms1bkTw+YQg3p1rIq0AD/F4KBkmsqvC3usDlzdw/2nCUNJoNnPrwwsxZPr05Qel80HDdCs7ltad
0kNVLYrOlyhdDXum3zFtT47UC8hkbbGgQcx4Uca1fuxxLn4PfDQGjJZyqHdhhyEYYS/7OKOD6jJ0
7YbY6wX9os3chNKWJngDmktv84BDn++nQLxibM+AdpxDoet9ThhN1LuitoALnQiJEUcuCijy2KiN
LMKTEk0q7FmQscFHkBd7MsLl86vj6ycrF9j4AhlbipkZ/ZIQ1vdMTYKzfkc4Dg7F7MaOVoWkId23
2aBH2V7SmQJWnMz2dODFlDnWowcyGgA6LtmW8TrZODov7zlZQayie9ghMN8SUcPqfqpAJZWQmnPF
/qJCiez4DT7YJnprrlqGAbDX77AzDapxLaYZxY2+VL3hYzrVvKbFqoF06z4J1YUN+nkdiP0EKWfa
MbhxjBMRu3SZkVuzsnkf1C4iqvwSQjCjFmDgFrcPwwShvJ1TLmFeTYrcTEmsJEFmHX70H9QUht4q
NZ5+JMLGXlLCdpzm3Idwh+OPBdtkPoO7zRGQcW8aeTJxU4vi2r9kfse7P6yhvywqjpaR8P2ZAJCF
T9TvEIp4tisLLbRoECFp17iWc5q8kFx6MjJXrcsWzWxYOGw5jAjMhQ0fNHzUEIBz9vfLsac4Ba7G
yPeJgeHOTGVfobfMADVH8K65KFVkYJ0xNvREIxjQ1CPBQFo1oXHAineott42rIZiu4JnBNSXw0Up
ngfyDQneNUf26JRRcrLAg08+rs2MxOoy4QfKlslMxqbsy61rgGVIGnW0axfDDKz9ZssQ5yhfzuKK
qn2Gwb3FwSH7EYwUMZooqh9VH02B8FA8b5mY1LzYzAL8SRdkl2pIToB/s4As6VR7ctY5o4VdY0HC
JeEid6e0gHVsaLNJEfrNvZL1sBgXiHT1zfii54uxi7uSFM0S8jCHJ6kBQ82dVBrBwD47OBBY6uGS
ArsMN5r4AwNKhvKV9lkXo5kpulU8bWFG/qur1DtGdmlvQZKcSOaWs+y2ZSj8ZXWd423j0jGQbwgm
L0IhjD44mofpA7sCDvr7hsWOlrMfWLSyG5iNhJzCTdEj2MYeGwIQh+AGSYFkV9Ggdr4xnbo23VAo
7zZ9/06XH2p9+VwDC5Hwb2FF891HgMftmdg4vjCfIcgrgzosaZ4QDuKiJUQ16Ocaq/epnVeQIk6o
3uhnXIteWllajKT+AYjdXU1DT0j1snEkH0u1O8bC+oDGZHkcGV/L/VUuNkV8qLy7eGRZRrItLOf5
xqi2v8D4cw5CE9QaqLRiMSVy6ZZTqDgYWdOfFijdD3APOSCb20mU5mZ1iSMaJVVjjHykhYqZ50ri
HAxhtMBpq+NixIibZObF10A155KCvsjq45OlOJkG8YcDBj3n2Tv2ZbJzSvdqsCGWKV/0zfcExMaC
ESd8p8fVl02Rl4BZzXecM0sqFrDp/lzi8njzkE80LnUP8Y3rw52QiOlOOL4WJzj8Zx6w9VbOKT5U
qc0smnSseF5p799P42LFTLZYYapk7PdH3BLPw/rfkDM34lix+NZH2QMjRTFSH6RfjUqt4KGrZoRi
EWitszCzl1eK2mB+bluLamiOFCqWdETNpF/PHwFq4Ilj6bDciKPJYfllxdBs2ggn2MjbB/uVypoo
CLdowTBf3cGNCMhTqEaJWFjS3YwhNPB90Ly/5kk+LY90tcG3+EROaMftqDf5ZZIN6LI0rfKeM7Zw
ddYk9avN1thY4coIXEtumELxzijChFfUvUwL9Gi6wUsLjrXudQUNM4Z9mxGLnXrxnZ2G3XjtJ3Wo
HdK6mIN7APB6/BbGBaKkqA6WfJHbCD8yfZ6idL/Gy8+yzvVwbpa1SkecpGc23Opu5opqvEkei8se
MdwK9wKQ0muRKwbsB8xVMtPMRZa4E04e+9YK9DP/LLM5j3gHVjtenPbprr7b8E4cro0460Ltet2K
WqwE4A+gswAwOuHzLHh5A+goO6iKBFkQARvNgkU6h5rHnwkpFO4cY3vhGhaJHU84LIA63YUPi63z
rdZwnlHyhuWZf9REhrMckZbIyiv/9gjMXtURteevJBZbr2VMMSBZYCHde8e9g8u1LqafkB8noMu5
u4Pyka32ZKMrmbY3n5ptamyBz9wN6J7CeOhj5U2CMEPeLwGbJhq95u9HrPXjYS/JjcUxNeuSm0OO
MxVw8wyq4ChaiuCzgV6FhCRAR0Wz3Eve6w1OfFyrdbrL3SitRYamGkcJoOVMh6wmXDQxdRVhyeJ7
8Op7gFyABgAcafNd24awSvXSViOKiXwtDLkRgmxuQKE4wyXipV8ZLWyngVbGN2RTNyifWAAUqnl6
Ki7z7MKTf99wGcxS4RGAfH2+BY715vWxix8Hzo8jpWjoPOGouuzltPx9BkgYefqDg1USoIcWMRoH
Au/ydTTvvrxwXY825sombxnCQfOKHjc9rGfbLNfJEtA0KmYzagphKuxPcuM/DtT2gTl32OzzdqZE
tCHmxTN++8/8AeRH6xJHEP0H0oGbMrvInhhBiefyAhQK6XdxaBASAZCW68DIxOfMTsU5GXG5kiMX
JPmIwpw+X6+kqMDXj8w5T/rsIYnefea0WStwHQ26dyXDHz6VeOl413aZT7aA5QDkPLlBDv4MZ0d8
NLfrARVLWl+mCZ9QnWuP492e2MqRlcT7Mkajbsy8o+L3dKhFJcgFsyNesyGqR44n4J66YgCyn5B5
3VlpZrTpHVuXAGCOubvG3JiDdcHcY8i7R5+vxYBINKLyH/bqiJXbSbYE3L0wWaH1ktn5XwCX9GOQ
6LXx5GX8ZCpzOqbO41FfhwK2vvyIL38Xidn0qJEjD5o2wif7rpRU90jdopBVh/ENpLHA3R9YCbcR
+JU0IEXUD/N+LvqiHe+nIz59xQaTwGU2ydfXVkdmWD/54qrzPHx0k3IitLdqaek68wWpqdfdoPab
7GdwUWbZ/ctMTUYSML23lFxkLgPVMWlygkOAe/pO5L6zH3BgyNfz2aOI2Li0hqPnzEkdS0M8t5lw
XJs+EWzLFG47v5Imk/v2yucs3jzs3yX0xUf1iN0yYNjE1w4YlfS86O9ZNuyY4ihMiTKEZYm1IHZe
fdlyStgZmWfIjV2Y0u3e+FJ+1XjXvPsr3z7gGpQ5LvGGJyLZpM1TJIsZ/abcd2p6wdHmnNTGt+XA
LYOufFOu3wbkqq2G6PMPa9GlDSRLbMHxiEb2ZmFX285MjuIFsxHwnjdbcZoPvy1YmnGtAKdH01sJ
2V4dbbqYfezTuW5rAaXCZlPV/FMcHA+iHgSBWqMBlflO9Xqc5rqFEV+ZlQ6Ug8DvLp656uprhGE2
8rhJB0rljcLUfHHOA8OIqqrQaef43aRV92ozbAi0+easTh1Y/LJ70JRk//egTfkuKd3k89tIq/eP
QfMln4l9mPnYiO2zPmyqV+7poiENLfrVZnbn/7pqW8w7Wyt/cdobJ7eRaSYoxaAOCUX8TI7M7YW6
rNYHTfh1678W1YA96dRb1wARZE199/cBdIXQWqreaJyYEkskYEwqzgAJFjg2KBTUFoZ77Mno3HXL
5sZBWHYnosMzVQIi8JzOuUc7zCHvJYopT+0IHBi/eNHt+IeQTEX41b1klY55ivOd5uKiawPeg3o5
rjWLJ6PHiRODvwJ14vdOMKlwnOccBLiu3XgpAtXLR1/31AxTn3JMU7+UcU2kktG/ja9Q8Npoug16
8qdYNrqWAsYxcU92wMX+9mWq67Qk+TwJQ99xJIY6r2takqI9VJLzVEN7dlDQt+hZJG1TZJmiK6nW
7cRQ3r26sklX+yVY5XEF6cDca2l0XxiKAod9K3rTfL/ogMA3h5spWtq70YH/5ozA+03rl4WgbdBp
geTtGk8BdZFF+JrIJNpGFRfhWd6RpO2ts+q2MJ6hRgD20DS7s7BA1DWZlmLiEOSoc1d/lA9vJWv5
MiVucIEDMmleb9FH+PVY0iGQswszCiuBaFd27yXhRNDJZkrHx7L4xqo9r4x+TBHjIVUXF5jfGuei
OAnQysKC6bpc+9oTyzX8W+9DGnjqCOrafWiSJrOOZudFtDN4VKVcjiXqk7ft1mH5b1L7HPrHIpq2
zOei+SR7/XZzbFeVu8yg78l0X7vr/KJ4EaWrrhKk6W6+JbLkZxOSD2oIJ4Pf8cve7IK3UWw9VSai
6/XKGtjoJdcgznX7TrB5mxWex7TeLqmT5gWispVa6dCTWL4aWzA5zEXDvrHzFK9XT2ASTr6rTu8x
RLXPF8HjX/wlZLfyGDXzozfMqeUFQrKpACWnH8RB2O8vZKT269WTHW3EIjCCOAml0B+LLDwcmK8d
gGO3FokdhfSfWPeZASavBiKjKMz/HmnpHzbQwB1GPezaaM+ZnLxdnxd6/iPKhIz13bTHChbhJYBD
/d8uqvqzxT2x4Oidg1Gb/ZL11OT4IVPttPM+JaiHS0lRrdKIPKn7DrYl/Ma8ku5L2PB0dLLfh/jZ
5uL118OGBIrFQD6k1JbKh5y9zOq3Rl8NDw76rYfQIMKOonMrO6mtj5Ht0YvJsNXj9GeWzdoKSUYa
HIK++BE9wBi/TDWIH+mG2E8bEa51MRVK0j3IN/AIWkpz2siZ+MKB3V/K1w2zIiwttE7xIVucNntj
E/yPkCtDskwRkqfJj0DIxId3r19NZgdrtJQAhc4nuYpdQHaFd07umQmxI7scf8X0Fx8Yc41rXzjD
Obg6xjR3po/Ml+uRI0IvkVT8679KXlr8/eINF6w1wl+baMYjLSf9uadRyMQoQNBW/ZQNZaFJgRr2
W/GviYcmrKt1e+oCwu4h4xV+QotwRjY9hVrHdSRatN3Lp5dvKGZeVVSjqLtpXSYQlSsRRsV399sv
sXtEsq3neSD+W+V2fQIkGuKFHJTPx3FSmppRVHkHHfH+QKFdswz1+GR9ZdE32R5jrhxLY4ocBYpr
BwCm1my95JcAyQ1hCipv5wc58NG5+kwclZVCRBLv9BMpPF99vxOIgiBJEkhbkW/88CvJjDXA1gR8
OfRiT7xStpHBvAbDFetapadSQPxXbrfZ+h737OfBEJCj4v7P61oGB0jCK5VZ0ufXxMycyxA6ZG7s
UT/Ql+e7RcU+FeWMyEbN+u1ywngSo8KtYGsC5pvFizPW7fDIa8a7bc3YVolzSl3WiGuaoRM12TI5
+jLurrVJo2AKP/WvLZ+CRL6EiG6foSNOwZiArqyoRk4kCEZ4l1wMI/HCFF21WCmRpz0g8bnpmdkH
k8XhY6qs7tELf15GaRcWMbFN9cUvWNAI1whZbmBgve5ZkdnKjn4ulPLPwLNWNp27idjYq11Zji6p
lr0qvzAP0JV+QwDz/yVu0y15WhVwqtl05SCML+wIidH/QOqIND+PT2km1uOyKo8Etby9TLgALWBe
bv71Igo1Dqbzcn4eVp8t3JCpDIEetqBWUh/h5GbBllmw27BfsOUtR9feIKs+8egrOtbKu/bQSNIl
Srqxx66iKldxMw41L/YhTKaz4YsCpeUnzDvZ3hd89/n9uwQkydsVMZ9200FrO1AjQD49zHZRoKYB
ieVlghpMueiw/D5v/4hPjLm2t8GXAGbSfABaRjE30MciaaN/heyiezjnLFoSQi8jqcYc3qNUkAK3
c9bB0UeOV4ZPTqDlYVBmE15LrjcCDkcMxWyMQ0eygTtkWBWmUeznluqkLySNKcoQ0SPpal+ooWGP
2f5PJfgZWj8TixV5pPlJT1h1NUWdV/NkV/oij7dGKGV0TzwqnLv0djvJZh4R3Vr4D74DEPHCQ+A8
WXRFgsktFhFiRtluzYLOyW8aptogj6ay3GU9BwmrDvf7rei+5uccIhlhIMduMJq2xHlkgT+/vEZs
zcd2LA7aBz9vXKdmOWXoLhzT8OXnPJgkOqqfwU4inbIyxPKCmJEJnehTKFtUC0qkkArC/abGZ87b
pW6yCm9DdKp6Vuz4znJkRIp900PDZbKk4ACqe0QR2DTapSTxjw1j0TEemWocIyIbM0P8psZKqmlG
L5ZMIanPe278ftgEDetn3npfuHoh3CAWVIOdvKS4TW+D/d4Bez25MBvJhj2noVqVnLbr6+Kn1kB/
U2XH+42R16vGChXWU9FP99na/xacqXBCfdGqJNaiyUlgZKoDiFq93YZCkGApMZrnWbza3J3D7Kzb
0XVA5DdzZgduYqqqV2A9alAJCumPEJSDbZBRdRSgg6L1leCBMxrmOyu3wK5U9bYpQtv4ZkqH7fil
5kZgFXTkk5xL4Omgb7n7GicKLgHkM0sn6Xj6gfeTTaZ45hHL3Em1W0nZR8gVirGxd+zfUTZDRaaX
tip77tnd47ns/DYzpoDOOdWYzgZZ/PVDNk6EuRkJBT5EJlSwUbSBrAQ3XGF+D8VRqUDJLO3floQr
ta0JjgAKy7HAIJ8481+V5I0b6o8iXB119FMdyz+NArREPMyIP7x3rRHvXbD/e+qo6WYlZ+mVgHVm
1didSO0ep/IS3Kgox/LqCZRT+yHgxGZq48Dlgz9dJr8vmNuRegaY9JQztYIBoDMrdSVbAMslZVTe
GZRWgFhziyz1FqxFnLzsLeYP1eq9NvW2FQd0XYioNi5unkQeMMfDVA/ht+C4m7PZtYThzMVtfF9i
L7/j879Dtx9ZQm7g3Q5NuGubqzK2HBBk6ivIkvHwzjyaW7pXUcstkpmXwv6P/yTPOWrNY30PqPCk
fR+g1E2CKyqqjDBr7ctNHRRrOEFYuJ4RfhppDVD7NtKueuW3MQ1j4XRvex0l8zCrc6deKha+wQ4i
IUdE+IYBOlduexb7ckVRLOY5kJvIDEcTC2wDnomDGU0o+zN/aV2LVcjFOoOTJNxPnfAa4rswICfG
FKAlqryOyGkApqooZ1M3lsYggMZaXh/+I/0Fk+zsevseE7ftvxagrnZESJCJ2EbaSANvu60X1ZJD
uN1XsmfykIMNxHl6xMACHjIahlwCAQdOMRp/AnHGxHMAFrHGklF1rICgtDWCU360dxHx3n7js+Kb
wWR2nWw1DErOCf35gdo6rg+uvq/vf1GH9r9QQWxfc1m3OXaW86ZpEuB3+utQ6wtGjyXxw4rOGwm3
5ZfnhyPxeZLR25fsh+8c+0kXYSkOitWyMLca22FMksrUFfF1OSlLsDn2rJqSSvh2di7gM5tzVGF5
dbE6CMbz7ytEWKKDTXf/JU3A9kM4kPVLu6NZZOhUVntgow6TPYLZs57V+ZB15T+d2h5o/4DBiZBP
WaakoPDpSsQlbaymbzrmATNf9h5GjUfQVxXaSxzsz6cR4BCl/jvrwQm9tNd+ZMHThJZ3mAAjyevO
iIowIG2WpeeDUyScOcjA8BJduuDdirMy1RV2KyBmkmtwV53KpIxFuO2rbR/kTvhN4lD5lYlkQpdW
APh5U/KM3YF6mtqpF9ihSeivegFHnDiQc22h2CKR88PTb7oPtophSX5qHxEp+Wlli9GXVsk6bfP4
UGePcvOHdP4371ofsHYM01ooaOJ1oa8FrPfSlhshrZch2U8Pc1HUTPOwcBIS6TOwD1VChLvLM+Q7
+nm/AL/NFUNX78Q1hsq1iCAfnLBufXbYqXvTk2rPg35hPKjJJ6N1R/dm28x4vfQcwG0o63NscSiA
zlrWtF7NOxNN+kEc/Uqcsf5Bj4j7KYodl6ScAlIrbaV63zOCQt7hsFMx3Um9ENfHRUoNw1KGEosa
CGgXWWfVN7h25b/10xKiInzmxsy0RLbeD4nbGPDYsbWwvnR77M3EULrtSBgV1KAG03LBK4i7CVdu
g1x71sP+S6L3ENt9HD8zPthC8jxLrwW+869azVJw99ehh9UTTwOkPe9ANJY2QR19tU9a8/1T5pgf
qZ0t+CejjltQzw7tQ8kUGG2vbB6s0hTRNuPOXoEM5ZyN3m5cSXjrI2DQLffJats3uH8/CZBbJOF7
+VSlosbaNa/8gIWjNh00dJzpiJjTFnWNX7UxMZSVl85cTpK/xWWwuT1nwfJVBlYgwBe9bQJcsqO0
ZLko8HHTBOihfyXEBbBKS7EhhOPX3/sXIQbvBv51Z6fkWuV9bJUNKEgEsEZwp6z0FsDAcyu/1oi+
oDLV0A9qs3tYNBvTYwN5eB+7NZL+D1tBUWqAMrzVvfCNxHqzsKVzsf6tvMux+CtaDZszayIgEMvZ
lFhwBopx47ZbNVtcM77teDYn4jwMNtCjQs3q/CrU2tckqAO2kmE5lfILxrX7qa41T2k2415SXfhl
J77+CIT8wpTczw3ANfoqyGsT9A0GKesE9Iz5kfFsPtZd8tC5YKLORVzIDKrgd7WPM3OReUV1WwLc
di+XRSBtJEWKG1bsXkL86IFURBaUDQlQPDHAjdhMQV+INq9Z1Qut+7jO3TAAbqkIwPcisW5EA+Se
gRRsMWBVD2wSxfpJLy3+kLfiOXCZsm763jmjEASW7cPIEtAUjqpqIZcLkSPneYzE8TX6BVS/t/qk
c8/g0p/dxGk65MHqF+CO0halGxSQWplG4ez0gp3t7maImZKpyNoOgLY8zPP+VNmfIwnJCqMaG6Ze
sVyt/CuPELsro75SPa3WMHLWt+Dpqf7uJPXcFtTUEu4IM6X80hwmlYjAIELUFbW4eLh2NqS0DhfR
guFFrXxY8iXlbTWQctx2QZp533moJ+NLr7LUVKMF+/pc3UebkxWMJaB0nT/IcLi1bo1iUDYxJ6pA
OsdKzRrJ6j99PzIn1iMqujRdUx29/627Mv7BloCv/uUUJaHP2ZduBG2KcpGBo2M6L+AEwuRRD9zM
JLd+4cn8VH8JZnkbAmKasEs6w6JQTziZOfghv52rL222G2m0y0MNAHZvh37wGDrnOmrrsGH+RMv6
w1WCOuZqmS8p2S9twoOelb50XwpY7KeR+HyXT5lWihwn1mPCDa6X4f84njUy0tBe/a1gqmGDphwU
l/60mbNPqvwMjCnWB6QHKmNdCj5JwtRwXJ9CMgMrIXu1MbhVB6gp4vnEmxfgWqPBzgbaiaxTP87Q
lma0co4VgKxPxbyMAfhO6Xfp1f9pOFR2g6vSmAWJWtqf/A3DfEifuSxL0U/oEGbSOeLA1P2KYcsV
qcnOs3YBHDOG9HWTgTuu61kfZaW01gWGVZ6el51AgCp7/ywWKm0ie9PMcuer4HZNyobczfpfDwNT
bciN9sRfEQ1PqVZ7DTxwX2LT2mSmu+fJIFWuWET27aGNiayBAy4rfKbnnwJe1lPMx3RcsY/o6Qxr
D8aiT6PlR36H0BJPWuPfFoF0afpvs+WeY6at13ZNHLw7p3kARlKzjbrpmVPqut9VMdm8VIlWASjc
1SlhfeNclaNjI+ijvmcwIDVCW84Mc8dBVzM/jLXeKCYHNQhpbK4NFdxN7RF5hvJjapuOwodVlCUf
Jgh1BFibjiZgQZFA5TbhJaHcjXGTm8hsl6HFvyoublU69pXOQ3MKSkFi48Uayk9Kr+BwM04ul6jL
rCTxAkZJ2jWCfvHRmpldc74ozx0CScVVJGRUXZZLa7+zh6QdLGnnyKc08mC9uJA5axkmMSZRpql6
UG/r91osa1AQvacKei6dfwzLZoZxEw1ahpyiuhwmSiAH8FxVHxcrEbMyNX+GK2CiSamOj5nC8Puz
R8PeUjFlahzohzfaEQam2BXEx+A4cgYqZqiCMF4HqYIPWUYn8xl93dixnay/p4dmTnc5f/ROOOfF
rhz7zZbkH6D4Du30/t//NPMAZNXqXkhDgCuFBaQDL3cImo4SwdaL7s65DLxBonuB9Ue2bOdc+Wa9
RZt9cShVIhbwiMpIR2NaXLvYAslflyDQ2zxytqOuQg7neW73QCTc62vOL7kz0waS4Y3wOg/W+Cao
yXNuR7mQNVdGxq/vvPN4KjbTtQ5y2cxzM9eHF2RDqqUrIaNesWYKMTg2yb2DUvEo8ut1nKaO+Vxo
UI59qkQ9+SNSEy5b0jRoFAbwYE6kBbOUwt4n/HyV6gH5sPSKzGwJQvwsaBu9xWXbdZn44OLOgquh
IhsbtH/DH8j11wAz8eunIZSuiy/eS/IHqHJHbumm7jOHUpHKTHzjjyJxUlxbN0wLkO904z7SmJWh
A8d9Fb6WWVhA15gAuGz74WALS7wHdUiXtwQzq4iiVjyfgSThDMvR/neJI1iqD/Qmdv8+if+xpv0Y
tQE+M8Si/ks8Rj0Uuude2MhWgKO78j8mN4k28BnSEEJkPUQ15OBMBX6Jr4IcjlpsMDE1HZix3hVQ
RFT+fBLRr/nvWUBgQpPY6kQQsRja3ytUENqcqQ5+qjxEYdV8jl2wqypQFB78A3XyFbMRmAt9pl+8
ufyYDyLpLPHHAXGYbJIFUDKeggiwTDbTk8tJWt2/5NKfixjCTtWY8kTHjBQoI8xVyU5tiSUtoXsB
hHwR7ky2Q1p6sAadat6h+7kSFIZZNN4p08RBgpV8lWUpyoOzKo3yqkT30xkZ3rkhTgdIMweliHIs
BbL/dwO/g4qIxM1wle3GdZzGuFdNm1f/716RLRC68vRLjwMoO5mDeHiXYlbakYpiUVIdGrEzGwus
t1EFzeGDh7in+Y0O1hCKeufrxshC11WUXGnC/JvOw8d7MGSfIAq1CUCbIHNaph2hqMKBaSlgZoz+
pd0Ytn8TMBTxmC+RFBqP4BPzCSxjoqE1+Mw+D0SRpttx4wiwO6YsNYZneaXnpUdFZUZkpbEHKChh
g+8c/GHid9Cg7+mb35qqTGUW6vxIxYQLMo2cMmIqHQvWOMUzr/Or1w7WzrZlHCMpWL1LGFj19WHo
mywOArojz2Ux1ZVq4Z39nlXCav1nmsFupEDY7fKQvCD9kRfvdkRDesdxUihfu2eUItUJpZOT3Rhz
y+HdLNHIvMjxmV5fG8SGqFBWqXHWZtC/MdEiMd+zhhcb0DU/ANT2wESxnXn2GErEjIzdh591znxy
IxhDBCqRmtxB81Udie5mP83CFQq0kXiJCidzCINSXIyCLQO/3K6LL8MItF/j/r5t+lUMrZwHwKUY
WaD0Q2Bjh7HQN5aNMJu26BLR20kwrQwZ6ksmPBRTYhol5zRI474e4JKtrv7QoEc1yG9xC1OSAWwn
GOW/YdLyWTXAyGWO9jfCGGf7SRw4GeuKyY5xkHUCKhqp98CjaLA2QVNDI4n3bWkNIUT3Y3r9Rz4R
gieIGgRgfDxp+CXOKEZ4sr42yFtWPWDg3Y3vPlx+yIqcx+TS/0WD7aI0c+rQ1DgMmpBQ9mBWefT5
ZkRoAHjVtVJfuNLSLautzOw6A1MGEcwWVbWado5EbMYOCPe+Ehdz1b3lyhuMU8828+peuuTYkmMN
B6a2XIPu0Whu7E7if63m/MxYLA68a1V7LQMgo0FEaf0kjxU50u7QSHgR317xZIdSbVjwUZ96xg4t
ncpm7NxhFgdru5ca/Fhbc3wk3DeYjSbyprZCDVmbV8eL5qYHM3TwM5kwp2HwPYjbV8bd/Hq4hgeE
5oFZzj1RAMNn+U7g7btQc9lXu20pGaFu7qPrsowy+BfGjlmNn4wLb/CyZ4hoDkk7FDwkWIEquDSY
9sU35DwyE5aTrObcbKsqkOTUejUeqypm3kXgBmpoGemyEaMSKVPEK1QRkxSaVrGfPuza5Iw/wRmi
HuYehIYzFdxxyzBYwVHFlQPm+R/H+rqQRI1EaQg6hRY8KbQ3bG8zNyu3qxDQ4S0FceYUdI0QpQW3
yFBZk+Kth9lLRAqWQTwsvInT6JqUYgsgE1HIvDKt35R74k21oUm4V3M9EhfhhcVV+a6CpdDVvc/v
wqZpbAd6CX3waK09YsYvGQKh6sc2Ta+oe3estBvmTjqF4/3Tmt7H7VwONhIalB1dHe6TBOwfve/4
5gryKUSjCIVegajJqPOJ8cBD+03LrqQKiXJqXlfc3FKGvuJZCrrpBZrWZZhBb6O07zw9/+oHo1yq
LM9BZiLLlcS43FZqKP5W61omRN0/qNz2Pk5NoIWQKSy8WJiCYzXBQVOgcG76CrW71emPP2/mXXnD
K9IaKlh5d5UOSS+cjdVdbzzLi0TyhGGk5xh7u7RQOFCardrASaHU7te2w3ZKvDdigtRQJmMGWVHF
B/HpKLiVNxExRZ64CmexH8GDQtfELmCdkdzIXOPEWW8AJpYQ1VEliUVjJHTxSgmY8eWxYclUiBqW
wNx8jkwiGpdMuRR0GGSwJ01JR5kIzx1IJm4fcm6uvv0ByHJCDiK1npD1OA707pEZr/4BnFtYcO27
vpEr8gEFdDs1iKHGXTVUkGZP1vKICRNGZVa6bJ6AISsnoguTPU011uGLZ+9fbIGuWsQyy1tZabi6
kzeVS9D/SjaziLD8Oi6nisMhylv6dFv0earzmRaSN5rbQQQZPGBtKmTHE3QsKSXRlnaqIrDYg5L3
SDuItz+j2Zd/gsYzxTzWPiidhjisA/RbBz32RYXkleXbVz+vP9eUKdHTLSTzbGooZGcuJRfmZBsQ
b27rPEZUJiYAUE+5DoOUAYjdou8qehZEHOvxExtbQH2LrcSNQOYSM2QG28VP5Z5jj4qWRKcbWuDv
m/RRUftqDaCadLsGh+1fylkVDYcExq4AdxMFEfNTj1N003ZiPHSqO3LcRlmyiZN905ewnbPVgkeF
M9g2oZAEUUycG+8fQxILZFihwLzCfF/YfSVC/E9WKsbLPiEsX1QYpGek7WCKaqwUwVaewuVT4Z/j
lU2oLG3kMoIAn2brB2MULTO1yo8yqx9lKEeNkbWgzNVch+HSWcnyeBE6tG4UbpeMysIph83mMhmt
qmkRyS6/xCiYVCOIYgil9hGxck3jDchoMtBzp1SI4yKwhtgoiRuXYH8AcikxOJEnCbQqGJav/EkV
/qT6T4f9qPpRJeoJpIZ6yL0Z9VCtM/dvR6LwkRL/4ijltRmQTsr0awkxKhodoDNQr9pDTanH0lVC
Kor17wC5bqoopENLWedHqmiJFb8M3jegip50SK8R8zlfMmg9Z6tkRCxcylrzbX1zaULLSzcSLyOr
/nUbFCJwv1CCOcat5yIfpZjwkJ8=

`protect end_protected

