------------------------------------------------------------------------
----
---- This file has been generated the 2020/03/16 - 11:19:27.
---- This file can be used with xilinx_sim tools.
---- This file is not synthesizable and does not target any FPGAs.
---- DRM HDK VERSION 4.1.0.0.
---- DRM VERSION 4.1.0.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinx_2016_05", key_method="rsa"
`protect key_block
NM3ChAZ5CBZFY41YzqEOycN1uwx/zUoNu7BOxx41RlqwVZa7zAvW/Ao9VOk21gDdfHLnG5Bx9GiC
OQXH1u6rhVpMzc+sFcFZN00s6JcPKpINZb5AUZlA47fVYBr+WR1APCC9FDL3st5RDeFkDITar8pB
4iRyypxZOZCDNhsA2wh4o4M6C1qMy4Wi7fX6Y5Wmb/50AZaOwT0rCwFOLRTHWCJpeSIqFyWFPd7i
vBzjOvb2GIWUgLhZjxElqPv81tqMclickXIvl/dgJy5tmcdAZBgRs45Q7PmFS22GahkCHjuCzJNl
BJ+gLUjIX4wRORy6klbc4eIJhuqcSebug3aY9A==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
YXzK52VaemZz0/IWhvz0+N6d0oId/7s42AMrs+0UBiFC1E2Bmt8AcJ6Pp99zpaZba3oQwTEUHmQY
6Z2Ctcsr6+yjw3RviG0OQY8I+U0HEp/EzWOR7Z863jXHNnBRLm63KEv2pBbAvyKOoYpAS/6UThQx
BpM6Ku+M2MKQL80FL+SDExNWC7AvosBVxJc0GoL16VrtIhWIyif/IJY3DPj5vmXSrkcFh2J4IKic
riAp7cVOdhtODbPQXuRAat81I8Pc1w2JSOG+Hdv5oYG+s/wqtl5pX2+/zYYAkz9UGnBalegM1Trf
DMwmDbpekBguagH2rWEXQGkKBW6/n4mjpVPG6Q==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2019_02", key_method="rsa"
`protect key_block
fnVWVwpB3IWiyzbNUE1lpc3bIuS0IEluQYsqIe553CACyCGunAGc+QWfLQw8LhIBxzNEUgbFmMrZ
S4Mm3cXVCBbcfpGwx6LJsGVmR046cbE88X87g/bbOTGEvf2EuijHotYLTZmZG/sZFq1CsVLp3KLw
/KI2f+30r4J9yZ1qRRp1oC+9Gf4ikL0Y4rsEGfHCCtO/VYP3dQFv3EhcXDhM6JHeD33yenrglvxa
yhwbZO1kHBM0rjoPe25lUoL1iLvDWOcvJBSEYKgkjFuYmSZ0vfTjpnjt1QhvpEzeq0KoZqOFefL9
EXySUt7US8gGDTDOJnUKN2whjaForhjhiKI/Kg==

`protect encoding=(enctype="base64", line_length=76, bytes=839744)
`protect data_method="aes128-cbc"
`protect data_block
t6J03XhftFN0AEj4um+ECA1JHfOdbZkhb+jrSBUl6Q9KBywAjckx/PWZAY3y5ocm3dYEymb1cnKw
AkBtMtJVxDJvvOzQueIexVIYxT1ytKZvp+TRlndZEP2YX/Zb91+v0I5bUDrxsjxjtkx1RaiPCOwF
3CmIFL+wd5AfVQKZMudWG/+ys0eZzpqdWvYsUwlXmmcJTS21JZ99kZ8pbbHIBjnk6wau/Vm1fpyM
maPJa3QYMbkCaRVWkqI8/+ghDeLL5ed5fOt0zbrfiGY4lVfFhLOWptvb1iWOoiF1ubJhKxZqmlgB
PoTGSdWhih5KvnNmbr7Mo5zhzGzHgm/z3cgJWNVH2J/ETANELorXjYrrMUgxU/2p26yVpFulijAb
lgYA/wZZMucc7QcN2A+bvWVO9LaMNCJn4sQk4RR2hDwMvhdruL7fhJmXfUlEjRynKvhGeLYtA62R
zfz3HVuk+/eSY8cB2PocexBEIFZGuP06tHzahu0MvAWzT1QxglrgdJjKzTNtVlKF9NBRD2PfVPTZ
lodO8WZ3NLaIxo6nrfRQ6e1I6rVHdBiehWlNdYX2ZsuVj1IprcpBx+0ieMnomrN5231KfA8qx5La
QKHhMDIaaLwBl3vwcmmgOdzrG3OTNQuKIX9zhwM6dyY/EBWLng694iCsbDNORy8N/SK5ST5RKxrQ
dmjob6dbYjk333nYnJLtXxYvspms3eDZHFQ6SrHFhSkmLNn7Z4H0o9PFElx2oQkJFddVBcUwe3zC
p1EbLNTpvTUQQkD75tmO74+POmEJRqOedxdq/SuZ6FQOVb5Pt1gWCVLpyO0z1mPfgJ/UsZPdLvhf
yacTRMXLI5eiiIszbtZXV5S7DCc4cD4iornQqvYOqIvA8fppslpl2o3KUQBI0rzKoB4JwFj2PwEI
lZ1tHSZicfNU+AAJ0wUQ2IWWILWW4ai2iSoDi8HsKN6JsyXpiSeYvscPAjneEte6S7OdAuX6l04/
R/+aGYdhMMfV1MfgQBbYeUQHhFe5s8OLdJP7U0eztJoowwclU+3MUN4WQUt8BeQ2IzxoUJhJQMbF
T+WxShSbDVpZO+sYALzVmb7Adh68PPmrHCnuGjc1mTfeVo9XDeEOIIYFt3/F8VVMDpAcxp855n1U
ukuKbhv2o+ZmJG6ZycGAHiNjv+ZMB+j7DBk9bJ531EztbUJSHs8rYgaI+6s3KU+6wUr1S1jB+ZFa
VQ7P1noIhSGxFCKhDIxOLRuV6paHYUbvztsg2p0qhdXSBXXSCT5UrD975tfEKBf1EnQIH6lUp68i
ybLSih3Hjd4sRJ8nW02yuB5CBWs/FfAEQ4NRs84VECANbZKCqmLNHyujZH04o3mmC+w6IkufjO9S
rfzU2ekPHrwaVh1V8NJSdSoQVbJNktsdqmLtEJCYEGkZdCpAwYjAJpzJJGjcMa6LfGVytJbf6G85
5uA+p5nD+Tgcs1IbfhBddjG7RDJZYlCRpV43SrWIdHQcFE3/GzjquS5RyWwER4YoH1ZZbWZzMv+g
oy2jD+nvLIzNgw6s4jUAppSaJkurLVXKkwLl70YIGOmnaKroqMKK63vwiaByyDHX11HJbpysb68M
+25+sK6W8mykgVOJVyxj+gX3QEWtCzWoQkwsDJ1Dd6GuFBRVvOx59AiyjqDSALmcojYcr7c9mFcM
9QivWuo3KagZWuss9uDyNH5aXHzvbxu086NKEyd0Ju4sgU7It12BXFcL2Ku/rYOcMEScgKS1CxSh
hSX+kK21dFiN4wSF13QkhfBYJagJ52UUdOweTGS21SZK4BO/kcgZ+7Gk81x2yBu210ec3Lnfc5Yi
Mu/yUbsI4wr80bEUY1+gMDZPDrn9IOhzV+RpWSUYFgnAUJr7e3s/N+R/e06DsCeyW0bDfx7A1rj1
+HC/DBC4+C0jT9FRRqjf+OcW+y8rvwucMLMF8X3YucrIqoi9LIvbxw+Bm1zKMca8RATzmggDAdK7
b0Pal15YhGZx0aVcKLFwr7JwzJzNrAKaWezihChLGUIuu62bnFE8IqOhZLEwgj07G7m5aCPZOb3Z
rnPPGC+XzkGn5SddETZ6zyR67FpRnUohvDlorJ0xX0ATTfHlMiqEijlMX62LoyFXoF57Nu9C7WHk
idGmok0SsguJwqJfrLPHfbFTEZxJVXVOX3Lb3aFbp9US24ouQ10bCS+eZ6R6drnFU9TXSLkeFCGX
7UmSZ+aSZ6ll55uOftROKpWcnF7NgZSYol0YL34VmFKWv29U2byiRqGqRapu9F/GZYz9ujr29aQ0
iPQjtsBgQy9q/8jZpDFdeSIi+Gw/+xIZ13qEOa0XXphffJnv0yogL+ISBXunXVtHeWbmPjBdFKgm
mpc74+fD06lAdTYW5kdTyipXkmf4GDImkDI2VJqPxwia68KeuXOMNpHmHAWZgnJW6XhMaMPSXHC1
5BlHhwhsIyXri1YrCq1aO6v8psLYnXz4ZWBnd3d0abYxiuiIDaqtjFjx+GRbkLgqRfO73K4UA3EU
Cr1ahPCItDm0izrSJgjcsmaYSs2Jecgzp0+1OWXlJHTJqc3oQt2OoiLuxU9TFrVRvmZBru1umWsF
BVoyANpeViJodXec4zStQftHPtFkux27EZQ8QZaRySaAhUf4KVQjW6B4XFUADRGsB/7jTO1PY+sK
idq6HQinO9y5MIQKeZSjnyAZBdwJxnHTlU/IDd5CpGRVRlSG1LPnFIVClxYRf0dfz3QHbl5uDtp2
u6Gtpe/2pJH42MUCVYXrrNHOBe2dSEBsE1G0GMnDDD8abK8BZfcjrT3NNMDgkoCshriG8MDA4uaZ
KpdZHZ86q2JMcqTO3Z0FAUFo2agoWsfkSQcr+NjtmQe3RMPJxfyPrnd1Zf+Vec0cC5HKKUm4u/ga
szo9p/hMeVTQ74idSh8j3NsGB7yQXtJyxiWZbQJevwOl5BnIVkQSpH1biAGN1fhLAKhn5sB1sl6I
CjXj0MzKLRVd3g3CwTGoHVBbdEXJR4oP/Rgr5yJDdAmWUMWPGTqn+QIwTgDP6HuKq2YNji64TaYg
nOaC0uJ1px6a0FV/ZzNuUPk611jBkDtqpmTdGUAnLR9RLt9sO56EYpYtapo5I2cLYwL33wxXoLO5
8ixsz1l+ZGqEqeVIsb8OUHF5HWeuufNXnKViQq6ZJu+CCr7dQP9Zp+fOA3CY8Xdi+2UefBEHupSI
3nziE436TR7ryU7XcPUPlMsaScT3zPC7766QT0GcfebOPF3wAd8MrocYOIwCyKfjlnWD1Pf0z86p
8L88T/MQdK4SfTPeNRYSFNbfHkXD+l3CbGUPu+yi8t1IcyUkx/uh1wJ3PTq4vRm5ZJYCOodMiw4g
eh9c4wBo0z0MQiDuWKmjxZQjtanvuoGJmB1sWoAXpY0XJkPFTMmP8HNLUr3qzfNakmWeULnoAjfS
ZGVgZH9KAxMP0Dk7nc9h29ohq1Js1LSjDiHrkE8L+DD0ni2tPnge6GnSCOkT3kXIK2JC66zB2AN8
4Gxhj8RNtufrrdhwBBpC9updgY+OQDM2ABi58hjLLtqMKSYlAhKjZfLpECSHS+aGZ4+AQ/3JmcOU
9JdII6cY2YlqhZC5yh2Di4cZY6Nlh5ZcojCE7CMmayIv43zo1N2Q7Y122EuG0OtVgaOYX80FdluX
SulEwwtKenERl7pI/qq/asL7FeoL6PpL9xSdOjBVYUE7wxt9o5szonR25HalsacgcdrBqzmaa3/M
Frz7DZX/wDhtEcoKWUU7DBLhtpF7P9LS9VNtM2nC6fASC2keRHPhwqlCFmRJM47ZNOcxC6pIWt2q
PThqra+oKGMsi99fPcvuRSXQEqdKII3SLhLJQ1J9JPEd5CMs5/ApoNecNLFhXQv8lVKhKeglo8pV
/V36ORsSkBZ1VkcLdz7xS5vmMKU/7y2eKRrca9yFvwqF1IiY8FIjNh9/TV5weF2HJYaL7JxIYwJo
i/VFqJ2Tmljhh3khoZG8GOihoi3gv8ZmrdrDva9AFhoAd1D4A3bu0A3G5DDAeZ37gPo15oFXexFZ
4BOEcq4dcSeDOsVund+9nbHKWuHIzM718ka5XvzD7qoKyRz3dzlw+C4QOvI3guc2C/cfPbDIqiQg
CgaY3VqhQL7tQa+v0D/6c8hsji8SFg8JRF6svOZ/Im17C6IpBNxuh+mTbjUGFDo2zX4NJO7ky48D
TBr5V6NNxGpYbJiVw5BaHUFPoqUvWwiiXBsAZ61YrleArWjbdJD7TUUMnzQ2IXdPJm2jCp0VneUQ
7dHgWU5DFjuhYTqIGAk9/Tr+RX9lJenGVYIZRN/Sa+Zj00Lkp+KULxorC6zR5dkBu5i/KuAFIY8I
EHhyng9y5EZdCVzMG21KbTYep+mKkk7DRSip6d8NfTPtsvfirl+/f1mXeiy1puKrNvo28q5YjsAl
W4SRIjSYnalBkYHaT/9jcMIK8bqpRhB8Q+r+UtMHi92LIqa3LNzXu6azeo0nA14ROYNQm3pOwa5j
NAYcuiMIKka1S7VUVz0qWOBcbbChXuW8sHWUukXg6PEh1Y+09PoSEdjeoaqoGqXIw+3Z6ktiAWaZ
foVsr2EYEw/qR30W+qcUWS/95g8zA99TfuehlVC+AlZTfw5GfwHqNm7YUt1xaVUQIfi2EMq0P4B3
QvR2+KEIt6qK7jUmp3lDiWPczOl8UDP8Hu+ugCIZPtjOrrM/HwLFcfjXn5fmEQzd0fJze9Jft8gX
RiQxocUck+Y90MwZoHOONLu7KMswRdcqY4mthZSNMO8IHq+n9y6wb1plmk44cgH7do7jfiQde8S/
U5XjrmkF2x+/tojMPkU0T2oo8TYrHBW2I1dwmChrjsD/6MwMMufH4/42D9PrhWFglMvv27GgTJqd
9zdhiJWOcF8sFL4bQDT8xvj+KU28BZ9UpbaOX6l9/UFj0exXJx8WOkWC17lVim9VHtl2ZgZoOM/1
Qwmi15L+3iDipKB5tbu2BvxvRRm+28HDEhP9R7km5zUUAJU6EtehA22V7prN8WIQnj9zCBnVOLzX
djlNWerREPtsxZcTCxMgJFvsKLn2S0YYnolFugZrEs/CqU/r5S5o7pKpGRRVco3DAFQATeq3PtGY
FtD1C2ueRkLE0xjeGImokLYSDN0SPlRsx3rD6FZK2EFjeUyi1HzPfIcc5fPcT/tN+M4/afWxSkB8
mN3JD+86NfszWjVlArRrpctoUg0aJbP/Y/XWXgneVofGhG1EsEFEAF4GhHVMdX5Srj2br3Y/aUe9
ouOpv3RToUux74x97Lk6G827BHwP3v0gWNLAKnrnfY8GVlhSK0SKHxBXuYoq79ZEhLFxDxrwNVAR
/z+KktzGEF6O6VxRHlHVNPYGLD9UQGJKMKzG/mZDOqSjrCEbrWfaB7df/M2M7V68cz7LSpguVYOl
K7/NxE0YpYJoyclLDXQhNpIjMt8e8QsBVN3o9ni4n1eSHLaPMylb4J2wTgj4pLt3laai7k15yx1n
tsWWNC6MUpx7zNRqcAWg5kKaQofQ6SyuvCdO/nQQVn7JdueVSyroVEwCwbJVCgBOVZ+5rfgFm4F5
MyB9uQmmiKRiZuMMK9WIyWTGdgiMWHv9Bp5U9to1RhgfSRXHGMreCNTFSm+LwVKMeeNdWxdQQjv3
Giek58SAtO5M3dwLwOx66ZMXV5CWYzrvCE+zh8HgcOIAC52WRE32F2wyqAH5bxyxSs1ZlN8tiofN
vb0thBMAH+lvhsbeVAQo5by1z4iPSfxmG4Hza2f3Q/boqsdcdDfX6MZWXbSU7JGsiDlRJcUMsO9y
d60QGc3Ja6gQju6a0L7yiQLTouTtZj9vAFNJF+iDT/bun5/HTX+rlNOk0giwfRs0oZ4ekuX0V5y9
yMe/WzkZiIrGZqU+l0i4qVgsqaK+tLTkEkniVk43UXaQLHQg2DSWHNQP5BQXC45G5WIVlLStf/Ep
ZS/RBaIVMu1vvpa0kYrdjfiHzJ0SuGUnibXydFzWwS0N49qm2PUsu75GC0fi4iAnAcB4AIGmh16I
6GpiePD7FuUdCECXzQtQSnFqY22HAMuglWexP4D7cNCaOcVoShxte5lmGhThNKy/NhkAorUIGQzX
i7cwJ1yMmFWSJd+DFFpabSCdbvcYRFtO9snXMrSJirc//HKWSgCd5ro5eA8nraJx51yv9b1Cr1Rk
ii9YlQbjXSk4Q64WEbu6UxpnfQsVtJP1Hfmf0dbsT+H7f/L/l+nl2Vu5JvIzKlmdULeHallB2dEW
Nekn00pg+RXC27Pxno1i0JN/6va0Rl2h6+kE/iCpIEA7MmIxUpUfmQhXd+/Mc568XwrvGP19foey
mQxWsYTRj13GcTYTTcB2E7JzW4WLIZzjmiu2HZ/UuB9x99KztG9LHu/+emc35LEwq5b3uXZ6LQf8
44NSqfApabv8mHDx/k0kMbdNaZQ77lr5AcQXtHStfOg+dBZVYwwyKy1DQ9oZiqhk8vBz7t6xyfnc
Lpfw/a43C0POoeke0rfItVB79/tzEnK7qcUAxyZr01jkSL4lPWSDOKABCfuJb3cuMoFjmneW3RNh
Hp3C3GtEjFEkAsMk4T2ocXmw8O/YZXI2aBU8JEJjUTbtuSrGBw8NLhiSn1DheFwuRxrYEi/KAz16
OzcYr5wzs1w4ugCKfZdWwYuEuswTDQsXmTwopsg/Q4cDgnmZy+uexNakNyB4XZ6p0nra0JpeEfSL
fUm7qkiHBOY01JfCayFiBYhuJpsEVbCAtVuFG0rM8p8wlc+3ctT7RGwT/IAxE1O2reLre3D63XQW
UU2xoETOtcphP8UKDuOWLQ5bfTI7w25biouPgNnDeJnheN4X3q8k57QhUAgSbDMVklOjanBhVr3d
546LwhNtayDcL4ZABOdsUMRwAqljBEl/nksmn3fNRZqwPIJkkuZAWUwFZ1rrSrA1PTWOfYK06EoK
gYuqLHy9g/gAJ0KeJ7h4OGi6xDrc/dfiI8/LP/5wh0N7Ox6mebm96TaXnt2DdHePhV5q1acm6yWj
HeJ721RZ6i6CKli9D5sVPa83mAgE3FyIS8n6N+/6LQIi73jrTEKTmJGx3ftJNddu/SdIdJ4S43ik
sCUYb9Rj03G4XyA67Xboy6qycw88GVUjUhzPjPoVfQoauchvX8NuJcro97aUGuG+R52nt3S+Vz/K
zsO2fUYp3OmqOu3zBkK5/bx7O4CHpQejb9XxK2Oa9C0JfLKNcNU0cOcDRIOhmYeBxscGi5fcfrbY
9mpWZi6oUG8beIm7jcHiivE9aLlHu0lV9zXUymwyAIWVKMI+82Jfpu5TVSV786RYppX7IaQBGucH
8+n9vGvytmY2F5JmZj4efpc0DwUdggZK3CzLdqA+xJyRvvhbpCfdmIyf8KvIfWDLLxAQaUk3z0kr
eaBouYEs1QpWhWNk32mxqj81dNvUoMaevbd9XIAW1OZnLvzNUXtbCuv1mZO23qqCHLOd5+q2Xlx0
oUugBrjpTdwgFvKKJPZ6EzPZwGOFXQ6WmGfSgdvdA7OWbroz9EzV5H8azH4/6ng4wk7a2Lx9htdz
9SqW/DgeswTDqd0Owpw6tY1FXvB1qxO4oqRD2Q/ZYpmuiYhvjNMm1IpHbro5XmAHNS7kL3wvPK91
LagYZvB4TOiHl40kqqH7OyqjEsC2t4ZgAvm/s9+Ap0yAUGsYjnAn7cww+lLr2yAxREoiZbqmCZ7E
yT/N2J52QiZAO1SBZGiJzKzk784lLYZfBNRofVw3hhpdbUM4pH6THuzx1NgYVnPsf0R9cSKb0vZw
J34cvK5Q++V9ZmIoIFcFqvjgnj6N+QJ+8XwS1wIDeAX41khr1Uld4UzSIkVL0VBYEWATrL4rRExT
boDv5amDWNM/2TutjUCPJATTQ7P9CIr0wgZUovjGs7quz2AOi9AZr1270LwpynK9btirZxvpFynP
YlqVW0PQKJ0T+JVuYBh3z4DN/YuS6Weyq7E1b0gboF92qskXxd3alTsq86f4GjnT36SUuR/4CppG
SXhLi1NR5JR73wJCkqvZNHMPfAHlSFN2IHHttt2DUIxb8GiqtGUgxbHF4gwtHrjI/90mx63xEhFp
+Zj+EJ7ta5Q8rA8aA3sUQEGU3Y1Yigd2eU5Egd9lLVjx+MQ1Gy3dzLTEOFu6Kdl3tvnHwrGP8ze1
VhnA1D2AsMicuIvnnfdsKm1MlFu4BwnQ8/pc6GWU4M4nEInuTuhBR4JERManoDusbib6gruwPxBq
jZ6hX+URSI8Cl1rHczBgcjwkagcOev4y3lqEk7ts6au6nUjiPVYHXzYe3mHMbl1qbip0KFmYSEHs
I1ttDC5B/GOA2mYqK3ZYyZFxeGTCFQ7U3oG0Ne7ecMtGg16loczYlErrLVhzAXhXt9OQbeJ7BqGn
QmpWcJDZXKbln45zq+X/9Td/rG0j++lrv4hL9Tl7lYUWKFfLTTBENs+IEy0kZmk3HmLnp8jMuGNL
0eJYr9JN2InZpm+2/zizJEg/AMnIjtX6dkRWvM+py9xwEoFbYG7ggZRhIzDAMLBYks/oxZ7OnfOz
YF2cXKgYVMpGaxGacDLWciYhdcuXp5xMWkkhWGxvRB8G94vHjrGsNSEseDd6o4Sy4Y6t7GtHa07m
NZAdYmf1yifGSENmJpMVyq8+bl7ZGiQ7Vu+wjZKu1D5E5O5FSb5ll/BdOzo0DUGQEYYr87htaNhh
/4RkWspYW7+KIFMkuqiA2NdWjwGPF+vIAYK39kb5aNEqk5k4pdgBU4JLZsxxGwTValZBqB5en8fZ
4SqOniIo27VuWUkBSodDwW34tkr+eQbBeBqUoSfbxuUPmBBO8X5bfnIShr0hDkCFKtjcF8FbTJbZ
B+8W2USLoH2RsXLSp3x9vnOi7JZ7ixdg+NnK/ImU96wmC4988Lr0Ao58f3Nmmz06vBok/+ikTh//
fF/clBjJQCFFT/yntI/NGQ2Dai5RZj2ybt05ggCEqZXtT8iuvq30q1SBvcmAnyxJOVEiSao8WYbt
1TtrOm8BEKMVP1M/nDiWBQppJ/sHfVDH45x+2ybtCQ0twQIoKd5RsFLtFNuit8931RzCWuaRyFIW
hTPzFpzVo+sqe/s0pKIqHRir0xR3DkDU58/K1Vb9i9FghItKLlo/H4HgUvtGHReeECfoOP3DhNba
Y5x8jarizKKx6c2U1CLT6oW+ov0UF3DbpbOVQ/q3D/TozkbQqmT+LNxsCZAgHCk+EpbJguIKskGI
lOxj+fCC6Gx4sh3pQqULVblmiUDSyDxzodcF1jlozUoka4G2Dg8SNm3NrM+xwjQY1uJfrpYJpI00
/qvH0jZCOQ8B5+dUnBrC+08a1OZlX0tKTDQQM2QgQh4SpMiPiqaRkFwdH2dTd2xuamX4I75f3Isu
5g9Kj/0TQCfz+gZoTs/r1xj4q9+Kp3OfVoHBdzWgnDThCXd9Qg+Q5S4RoGInls72CsmMKNIx+arn
XfUaFudQV+raW7xpo7vxuLn51Pt/c0bOgCuwLf8MLYitifPg+PHCQ75JBYN3TXrDv7IXh1LLG2e4
cUdMCo0alyonOG0Q05PdXbMHU0P+xxtPGI1wLUBtSEVn+HhJxlyrc8dYxB1w83jTTGe5QUrev1lB
rv0HOtk4ZWIm8Luh2K6W5vYfCWZjSYkp9ZbktGx/6Fp8pk9rsGWE+5xgYC5nM/8CCt4f9dEzKJMM
C8dYJmfPXky0Vjn9NAlo0+lKfm+CSpCvdHta9Sba5506Z2Xs5UJfdy74iKgCuWowLhO6LE1SXvpf
vqQ/kZKv0luXPl7GTq2rZ/39R//G3gfkVm8/4IzFOJH3AinC/sThpUWsKbVPbQwStwkcRss/Wv+G
y+zIR9hRV+sTpLTjY9s449c/r4gqH5MF2rxHx70HEFAEX8XSYl2T7ObGIbCYrgl8WVUhk9w6bidP
ROWgVqPC7Wgji3XgtJuOz0oYBY77jAqw79fftKpre9V2AfKMWIWKOrzDJsDkfgGGOWk7S40emAno
r3VjZB/q8FpugGIRYod3T+GcF9JHJMhe3prMe7JxSAdIQUTyATFDLu0UgmqlmMpkHcRmcOjsmpFu
N3T+AepH0gQHHVGKXcB3pDs04O5yOVZPqIxFWTzuD8Wx2M6/YmxLzGFonBJC6LUl7BSbGGQj6LJ/
IXsvMqIqrxo8LIJUuH3U/T4bRvfAu24MCXbWK0G6hInkgMNvfe8Oid0zOx+Dv/Z8ASGBXwubmB1w
n7+qUPQx0InVKOCGJZ7/Irg7j1U/ZrlPA2tYLAXn3NjoX559HzHAcbmNehzmk7qofDjo6Gi2WRLi
BOIqbu2dddpXySuAJAWsM7W82VOSrmidesf85Dgr+ef0fo5o9D1swg6I1NhoKFJR7dB2gYCbfDvU
Dpp/R/PD5eBqAAK+jqqu6yM9YRXhIiIPBTaEehVSUzrXhweabBKxA/nwmivnSk6JcOmzluU2lVrB
+XYK+dIvH7uV9IC0hPmo+9ydco5Ssyp3oe9WkMdbeyvpyBz9W3J888zpLFzt8MYFpt/I+zLNjGpf
9Z2jwVzBIV4mvuqmKD21KE9pb1j50WkEgrdaEDpaVOUm+7TwNo7gg7telz20sgkGLh+YC63vIzLm
AdEvul7W79dJaou/G0pcpNSaow4FG+7zjYJWxTxyIY0KgAS+ClyR9vy4qVt2g6NDB2LmYaOjkknc
KXcHR7eJHra9U9gV5yVe9wQ8wOfjnVQ3t6PTiUi5xH8YcI/ZTET4RwkZhFVDD0TW8sm3hBjzKxco
dvaTpn5M6j/fLnh+EUD3AdGi7DwNqmJfJ2ENs40WAcTMLxU4kfdg3s3UJmd/CCLXRb/8a+nNd023
Zjclmt9SKLlf9TI5Ga6ajgmWvaMN7hqxmAvrBb1zoMf9hTqThdn3n0dH5nmtl72W58Pxy8CkR2/g
zNtmjO3x5H4A9VOgyFhvy+XbL2n4ogYN72BCuYLAr21p7ClHtIfNbT8q1wXCZFklrMOqDU3zObsu
t4taF6FHEi2/7w2j03I7+n8nKEGFucuh8jaErGlzwOfS+W0Zu+KI/iZY9BZd93zDh7CJAHaR7yRb
be6SV1VoyyyhSWKH7lET/5zp4PFGnnNEKuR2pX6qL29XBjXHPZ89iyFbcwAsUMVjLz8yTHoC7Zt7
B9e1cpFjn5jaJ8oudnwAS0f2ay8u8c0zYGN5SQ+lkrSZ7wKGSGE4BcR3r+UOjQFfyEWgjDAcQCjo
IpCsEXmBMP+XJ2cxBJ+uP3PsHZQpCPhe5CQzN4nI2Ma5gs3jBMMsbyv/71P2TA1fcAh8GkfZ+eVI
IF5tzMwDHO3pLtM9UqUjFYxm8oZavz2h3OfZOQ0EZ+4gj6JiUuCG2Zoh4fpn6q6ykMVkV6KtSVTH
cC2PXwNnFn2owtIC/A8raKVio5Xh9dI8s6trH+lL7x18qTlcMTwT10s7RHYerAIiAqFjMFpWYq/S
aFahl/5LCCuELsnZsKuJ+4lWQHE7yyAKg241vcleUiCNayttG3LEKyOLZXgRvwV9CKMPGbvP9whn
U7/15Um+M13ppStn28fahKCcbFThlw1PzPKs8FldiDcFKLBfoJgSKdmDGQJ8s8l0/ZXvwNSQWqrD
kjhxs9q8WRhpArWHr5WmRkIJdrrknpGZ9OLau2M1PVrJxeSxvIPw/H0XY+RlPxNuUc4ljNNRqRYp
WKgljLlF8aYArDuFqplgyreaZbn44Bu1Jf/L0//ue8lucCS/cmw6wwUi89hn66FCKCBNVTYrmbi4
WWQB46/KylIh5FIxaEfcJ1MHGqvbtma0vZ27xuORVs8o3CbGvTdnWCYgvU3VBkxKFCxQD5LgY/SC
OoXjvSXle0UAbkJw4WliYiHF8Gwr9k4rUHp5Dk4YsJl3+AxlCpWp3o3u0p/eZlVHhbkrhCuBSvUk
4H9h5FneIYpnL9I+LQhwekmoI00vvvqlMdGSM0Zvfw1xQIhUSNJJI+fHdkzJ/BOA+6Q8yDCcmRFL
13wFxtx/L6X5QZWF5dcG6t6zmpVri9/+wx7QhTUmm04m7HAM9t4jgrP8l+mZGX2+jvu+CqkXofDo
IZzN/1yGLahOGtjmUuKrl0+gM/AlAyGFh/REDxfp65FfI6u7R4nOkggKIy2saj2ETdlHqOd8VKmA
z1kp43qZAY2a5TfdBPeaJkatE0t0LvIJUaspX4q2pDPgJBKuqAsEiG4a8BJ/5Kl/dXPw+1L81ko6
JyxKN5RvXslla3J9rRt4Cw3X98v1SMUKgNARg24XqdNhxHolxkjx9x+e/ZfDG7VIRb7vuGId/3i8
+2jvbIhuXAjgKk2ZZLSOJuHMbsRs1EXsVqoNSj1xn3Hiiic0WZtEfUYMuRU+p5EMo13HRSDa+5y5
72Bw+KV4RcgMlD8YIiotEp2tr2V37xjrG+ETwRFkFs/F/V5jK+5k5sSW5cTFGsg8a/h3nTmSrzv/
6ic8OpsI2UsjvhdSeLMOOkEylntOo5x9YU/SlLHMFYn7xdccdoMGjG5+Hu/o5Hd1rEXVBNAGsEQo
iTu4OY9Xr7oIrEQ+TlAxFMmkMErm/UY+uVatTGG3+HDhUNkfZI4CnpnMg0hHSE93mkf99lpqt6g5
6hkK0y+AYdTjQQ19rJCsp4Yx0azAC6MwuATwICFLeUfEr5iS3/kW8hjpuhwjkEgn782kgMFNvrrw
Tqw4ysTPx8dd09RU/QoxAArpmgxK0sPYqx/rJZRO7l3L+3S0u7uWxMI02OcQWqPv/av/l66VW9JP
Vq3+bNczPJ9lhkgKKfcw9xZxqbR4p2yaTg5Ht0px+5uSmS0ATuoq95YQgrJXq0OizGyo8v6aAHmw
7oM9IlFfcHdnbittSBshhQxycH+xr04X8je3RdVVzpRmrZq7DTEGQJb5HPic4bvZWfAeSBZdVoNH
Fy7DTYrYMp5xmW/+AGfESwXYj05x3d56s+qh/ODgu3TvmOB2+EBzfvdjP6nncs3Jaw7YzhNKS+US
YOc/aRn6fy4K7fwvKpgrwRLndH2AfLngDFz3HBxBB/QEDjjcoRNLUNn+ROlCNifhcXkW5v55ymzv
NEefxyRHnOeK46pYHOm7rWcFVRJEm71NopzdGNw1H/XS7vR+V4Ung927yRK0cA4en6GXDORyNrfM
F0lUssRfPLIwYELCRlC6ZKAROZq5KYKWEFP59YjmHeDv1ODl3DucR/mj0UeLAdLdyp7t6EEXtaif
6mssIIZNKF6kzkJXvsP8T+Ir+1aR0kkZgvc6Upkyo6/OD1gSDFc3FwQipAEo2cCO701rcuA6LXA4
mFLkse8inMJEqiQ2UtbdAJOZIc2LHKvxWGYhiuewCntOZoz/jWbPtpE2d/7Mfydw+EBDmR2Q+CNq
kFko7els+/igVx8P6/CDlTA6eFHjo2r9kePls44j62J+91VZslOZlfdrmi8KX541M9VsuvCa/Dhz
+rEYvqBb6CvwKPthKuuf90FlLhZGLoLaaGcJhrh2pXVRGxaqaON9Ji0Qwg4woJiKv7AO/88CAP2A
1lPKSSs6SQJyePCWGzWvmdN9VZATA681hhbCcO7R2r10cj/dXT5nChrDTQuYC/uB75wRp+2uXyP1
/WfIrJv4uCMMuasSl5vtqhkLvJg8VtzVR/qr7sWS/xO8iBimcfbZwNS1LWK2jZ6jLO0fUfGFewwn
nsFp7kv+5uJEt6drGinAPeoxv7IgUJCKI0Crq4m7c6ysAcCfhzw8NnVTJEsf9GcX76VzHqz3OrsI
MaBBsexXHYh/Ov5L/5CLROyZ8Rdb6y8XIMB23QmhA/Ie2Uky7eKQ7uwHb+VC37h7oqEMZJci9w0R
RZ4HSIl+FnZtV1rVNt8Ogl4ZaDUuouDw2B5+0Likay3pPLU1zvsQhynQFLZVuwoZoDnifjctF50g
yfH1Fq7P9hZ5d+QJY6qna9/2h3qhdPu0OO3ypow9oWyGIMsdYR0hS2WCedXhr+jGQ/a7av01OfMy
9WyEaqQg+xjbuPtfssEG8bK39T9choMO3oE9GgaSrsEOskjhHJdGntivDSar1XUfUuHNqn5GaYzE
vM3llgLnCX1ZPtArbUTdd3/jQ5f8BcxEFiQhzDEY9T1JkFsYB0G0xLZwn69GeXcvjg55wIkNaONX
eXEfaGgfNQce8AiaYZoH5HzBE73Lsd6k4fMDwHBd62Wm9PqG/daYwRv7IvBnGSyJdh0M4nlk7ple
HLSGrsJoEHsnMLeg/IK11BGSQQQ7v90J9aXXSF39u+UdbKzBFtwEAlePvtZMWSNZOUYr9DvAxs3C
f3XOX+bCZ7RDq5WwVCGm25b2sP1TSHM4QFdXIUHmIjP9vRbXkX8f8dn80hXDk+oz8ypg2TXR2u6q
/sO1E1znrRYrispUtyAduuzr6zPoMccGRhWc4SqDEq8gxqGjMMiWy1Jomp1BZd1WayiBvGUZC/Nz
/tgkHz3+Nm0F+4sZ5waT2YD0meH2IWXjFBaAe/Om2caq5sLNy/V+TnMaZ6tFJjguUuSK+UNy5A4r
jeDgi5KqNvw0y4OaWH36rrBdNlX2Uxh+Z/2D0P3TEsAWNPQdElKXGJ1GtbZOSPXvLEFgTpzWdpoy
2H62Jf99kkj6ZRMd69Ho1xUen1Vx5W3y4+7GC+3M1nCtCmLSxWQxDLdhgdJQM+Y+rWHC19Mdaive
qFD87+6QDWgrI7srmvHwZJT6pPUy5TEDHVQh66+Zye/1hiVi6ccdFjR3ECCInXmwrl/27MyHPKcP
N5dklkExmas+yHoMBxj4dE6NhHNDf/+Ftu4o3ZY5hEP6OGIJS89nWBhswAnoBOCcboFLMGFG6DPo
VenqkMI7+2K28ETSukKbNSHe1O4nE+Fb2sBdKQoiRkl9sgsBuOB5p11v3zH45+PnTSQoGQ/+ECr5
tSdw0v0NAgpFuWtxDo+L4UD2mNt+YUjtMhxFfkqSITC5eOF/Nj2OFkYxOEdVy8YkJifb+UGd+O56
ysOrwyUO5iDfhHyhwXsXRDSPR+i5KcpSt0GYISrciaaD35fKbDd1KwJZ1QKO75kvNsd+PwFpcNz6
rSU4SI9Jblv9CM9sEmqt6bMW9pKmTsTLeI76GGkaGGcH9Q95X6i6/lkWYXSUW1+WM9LHlPfGOyPh
+mOMNwXDi6xMKrFaRp0dw4GiWCR0zDqdv+hkwlayTeUdhmOD61dZVrVs9uhgjQYNRHa/l6dKLqMI
TBhJwZ3fy17MPSHrUx4B2Wss0D6tPcquWDooIbGMYeqyI0tfaOfxvFPshBprxZE2P2lHQSA5rWM2
s9vVeoImJL2xpLS3LLxb9nmMtfNhwT1yeXEHg0EYhUArSXR87XH+8pu3V2qUHreYo7xUQJaB2OIg
qiwxOeTm9pXKcKjJTlw8hS3te5AUniojZg9WCTs+9YCMAIKnKEi3GqL1Bhxe20SIEkoBbQekTabH
huG1acQi0AZTZChVaSk0zZJcZF+a3M3NFnuzLekkHMbtWJfJxrTv6IW6GYVSaTZchQi4kFv68ilA
PduXm5nacGd5yj2knOV5W0IsU/s+g2Wg2CwHdE4tW4jpQdbTKdGeZqRlp2AkQHI3rv8HSel1RwV2
qq7AMA7dBpMcFpOhZEz6imZ3aHt7U1grBX0SAo2sVVQlxRMiG/o8i1hqs+3c3jiUaKlgBk6WjNrc
ol8VZgDpfIDJLme3AnRdRRINVOQsWT3pPWAAJpcLmMX5LHrhP0JRMgsInbZhhPl6Pu/fuudVol6T
hZSJF/nGaotRSRtkTmMAmtKtKbvfQFT5Wx2QWKWksn3ovp+w17H8gaTG6wt43+W/0TOX4zNyB5es
S74jhhSCBQjshzdTX3+n/xd7N32rGLEh/+sQDN2fFzloJrJ/AH4LllqhBcSGry4uH8opKl6iecRD
7lBwIJLAkCJRDAAWygvq21hba5g5DATVSkGZGDu4I7GJAfEF3Z5fp29oVdAeDideL1r6Hb8Oljrj
Ozg8+VVl3FkwMHRSuAsBK1n+dqa2v619HLFDLs1zbRi3vAzPBUywiwcEiVem8XFnNpBBEddHTW36
ZcKim/sSNLbO+GGyDBh9jkXoF5z01H+tF914lbSlI06Sp0oRKJzcLkGBfNB7YARobQF7o8ZnPPok
3jyHQMZgtZQYWY41PUwPOGd3Loz5mLCihzXDtHARvMdwDGVvfpBufkXEczH4+m0kCRtemWz1ed+A
zbrL8cWpUag3A2Ur9xeZmpYVSSE1cKyoE/1q0L4VCHvqqYooP6BtClb+THkKNqyTu1c8BUuGBAMU
CEoGM39BpUQEsEG6fjVmWQcLaA0wfFydSTWOXIH6gVJbomRniA7WWJmVoNZ/AS3sVHDdcXRtihPy
fPmX45LlMB2P+MYkh5YcB3WzU5qsNv63s/COHS6LJ8F8sxJhytD96hxhFdI1raYO+suPdrh7Nqe1
rkXBjcXjFGnsYZ3BkKbe/MUjsSQEkoqJwD4qBWZtndr+K0vjfEi5EdYdYB7Chm5iDchZp1IOedM0
+BuJg6KDBoxn+6Qn+neuGk+pKYQIpefbeVh/QIXUaDbX9aad7nCyYCnsVJRywn0F4kLaE8cabUOU
YFxsCvLuEwyH64Q06mk98HU5lStXTZpDS5h3d8mz7gy3pTiU8TN6N5FFaNBVfztFW+xXZRqNdyyu
8SgfKeLKl0JYsk/zlCjbnUQR2yP8Z2KNegrEYwIxp4uVcsA9eclYY8m+Et+Jo8g7OWF4jUag14cZ
XcccGP1aRvvtE2JP8+OAj7nY6BsvyRfeOvCFbt/tmr/Zn4TMaU8VznGMZ/1n/Lh4GQQAtJ4PF+/C
rogvYsqO0d5dRwxxdebQ6z8BJfXeLJKfnwJr1lRmZWo0AW5GpSQm6CgwQnUwf4ESSTGnh5I0Ar9N
NZEYgdP8OP0em4iyMP5goyiNBS3t/Jgsd1zgztqh+N9d58myKgPMffUVEca41IXircnp5eBd/w9h
ncfqjH5WZg/YFYLYLalhqquJIMdTTvIJ5F4uNnqUSq13sA+14ms92vxYy7nmNSUmIaua9L7Gya5l
kwfAGbqEzZM0M8I144gFHNrzeTyrV+EgWhMsxl57JhH6BdB36RMuIT//L3CFtcfw+bKO7yyizuYr
OOC6FVdTol9wLiVL1xGAVY7QIyxtx18SOZE41JdgGTpT4AWbnm3KLxtrmQODrPF1+oHCz82hBgKK
XI69qqiV5AlehUPdrYxtRbCniItBeS9yZyxD0d8uHF3n0NJgLdfaHd3PDcN25R7Jwo6q9DBKOg9o
v3zAZZwva+pXLudW9lipTXE2C5U1YCAfhoL2q1l3PIIkm6GWhVwqxot9eFE0tEjwy0Da25/obTxV
TLv/vU1lIvWaRRwHxar4u251Nn7uS/PJ8PyPuI3GcaaYC1W5EH/nT94YaY7hV8ng52pOoFMA706Z
IO6x0Vd3m84LKkKm4O0AVeEAyT4/JvzjyOMe2cN68iemCHGB0FMdFoDE289fP2TzaCNvBwGlryxv
o58JQtyQ4phxJW7NlqKZ1TSdOWU13M4PzZI1hxxQHppkwztl2LuX1Pi5ju9DWCX+tDZ1eihmUC5+
6HEuF+TvyhXdF82oeWRH0dC67NM4OxG4yRaYvJ05QTNTBUfdoJyx11Zva8UCYNlSGivqdZRxot8s
rfZlMuPKrstJhb2F2V0GXBM4asdrYdudfzkhx4iSNdnKhR7irYoh/92+jIkQc97EpdUypORnLCtP
r11Ifsm46/M1mUhZWx92I9Cjx/sicubIHSJ7x631cPCwFRxKzDw6NHSOJuydX58myNeYOM0WnMD/
EvIEHcNvS49k/LpnHXcD1QnCVYosg28lkz8aregb9j11ixV9t+1p4WJY5BolS4JlMKWpyblZ+83c
feQNtBq0uVQs9OmuRFfIvD7IfRTGzQFXNmrn8TjYJfzZo91mWAKWcyv5KxnAcQpAsiFRi5q2r4RL
HZ2VoA5XX5vR8gtaCs6kMTIDWvcPTjE+/7dmyLv3Sh/xJyGjvB9w58r+wrQbNsII+hOvuPoPPS7s
ZCv/dbTYGyx8KT+9RgqfNJHtKOw9PtoHBoaCRmgFJg2c0Bych+oB2+A6fBilh+N0VKwJPeSiQhTb
Pw8Wmjcx9w/tybm7YafL/iaN0E3smvY47+9GSvi5u8bIwilpQhS85C5h732oA/oc6TQzHM7dg2TZ
jPsCL1+Kfrx5fqK/a1DgDLVKJtBaodwNP9iVcWdb+ZgIVfhdpJcb46x2y08LIi34Cwk9ykheNT//
IX8/LUNELzZL/fuWVcM+jmZEniu9S40yBe2UelLGx/Xg84HOmiFjC/yO/mpDe2DbKG2QRrKl/Pg+
h30Nr8KzA8rUTRdbTAO9qnDrEhZKVZY0MlLPtsNwMV/WQr6gvZAVT19q5mk/7xLsOya4XUDgNLzk
AIEPpnRhAOyl6M4ZKc5Xx2tx90sbOoj3/rAYoaH4IATryBjGdLOlNWwcnQNqQOVLZhdheuLnNmJg
gY6vC7B3GJrEGX1gH4xNozMWq/v/2bKqvjbl4OOJYbEQZGBxTuPQgS0LSmiv6SzBBj7iEZbM0R3n
umUVQ775H1BvJas09ptiZLwQsWTxNqwnuh882JyUfnnMSnNbHPElstkRCg+OiCMQJD69Ibc+rVve
nKR0GsiUiieWavn/8It3atrqSVC0nC5qVHI8TrQbpw4h8MdwVBSpSIY5CXReRBvgbpWLZBi+S+oI
FQUgWshXDTpEsdV/ICJ0NWh3GNLzLdZqiemPy/JhaF9yPv0CR3yz8RLt7jse11419JqB7s9unjWO
bJExVItdw59cE37eYTfdpgt+DqXq2cHikaIIqtVA0bxE8ksDAMqPQfwpG6Eznraf1X5K32GkzL84
4lS2r63A5T9IFc7RpziFgdDWjm17VBVf6nc0AGVvMvEAFjCKO8CMzIP8vZ8P2qrSgBTEJfiEjB/C
KLguPxJyoq5oUm2Y98j3jRA1Ki1LL8aD7uOTmkTGtsKVS2/LASrjW8M3uawUr8Id2ntcBvo2jQ5R
XmOHuio2PSJwrVjOE/V/WGTuLDxaz6GDnyCYMEUpG886SqGIUJO4uh1KnAY1vsRJ9FzSsi0NgYye
uysJgqGy0qTP7ngdIc6m6B34Ntd42aIu4CMAjZoBvBoBaSbKoC6m5yDUSwDWC14sv/zOX+QB2wDb
3nxSnHmdDyIlaXYMoKGoiKcUlXnSXzu9C0894bie8W1iX4AHdUz3Avkf8yKCPv426beHvBw9wtjW
HIAQh9TgNqGNj+7hBznXa+D0HUYd22JpkX3nwAiOTa9B1TVy7ZdMy8NQ9i3juKQ3CKQl+6s+dEh0
kX2X3904w4rMsLrnH4UKQXx111WXiSx5eozvqeiIW2sbmeLrN1YaU18IHxoqUR1aQJbRNS/qjdJc
Vj0R3er5i3/6WS2RBai522pOsDrWgFAXBWVTSgd+3pH0zvFj2UNt48v3nqOOr3TUcI/RlxRKDHba
bHsWrFGh8ee4zc6WNG+EdGfpZ279OdtkmlCmkUR7aOCr7/+/wemdiZrVl//dVljswJU92jb20E9X
Pa59+MS80o6KETl6U2+XfYPSSAh8jWCH5WUZuqwf3fAfaJco7H22oLal3ofBUQx+0HpJVEXd2iPZ
U/tHKW7DgnB9ZbEE/C2Z3Ke6StSgirXmv4NBZkjP8KgdEXR5EBoejdUjU3lyEZbR7aCHMijala0x
0ryuY2119Pit26vt8Gpm7RWsdsbV10seLYEsbjKOxQ0z0bPMhWZDz9KSH054Ba2p3claKyp2OnW2
27trr6Rd/Scv+Irx/1edfTsMUYSGk3gyQCKUClbTfDuOwOS2GgP5ICO+kFjVqui0P62kk5UhT7eP
PkxllfucKy34xrAdgohuOZ8Cl4a6TVhWRvoOKDPsotB1ebaJ1OL4d1IGqRh81meTZgT/RL39/6Tv
IVMPQULe1dqMsE6ouIT1cQ96uNULXs2pQJkZqYKEZMPOXefWpVVDpZjm8YnP/sv+Gdf/cmlgt4Kj
HNTuIDEYLQYsD++r4k+Uu1cTvvar90gZgFvk6i6Iag1ASRyNZz0idQVonugxN4+Mthez69pf04V8
OAwHyCybSf5AQQ1MA+nxR9tvIGWCoUiNJMSem2F3MPivpHe+GhmwH6Ph+L+PRGArO8ri3W/cz3bC
xmDQmY5YcV9B0dYuMHJN7Es9wxtLx0fILwSG8L2GzGEjH/PicijGodxwBoZDAXw2/oXcqI9AJQ2j
x5XTjsvDq9yX5IqqWloaf/Hmz8aRZDyZfzgBPrm/4WaKbwbcYl+fIyEhXsSyJLsiz9VSKWA3ZIzY
AywZVZBlcER/ifELNxKdt72GSmQeD0hknSvDR2p9PcTPrY8FFEPL/elOP4TYQRYUvwEdEKiWDdQm
oj3DmdXvFlMR0XE88dCdTRUdnLthRHVo+GDved5JpeZZur8AClhXGI4LpJCZZLg6xW4bJuay78Y0
R32VTaMVJENrswYyTQ7NS6BDzqkAjBajDcPKXONX1AVA9aqQnzqogNURn81xLY0m177sdmUr9xPo
ajTgDLce5xIufMA0LIHU/AMIzX/jCEGDEjrC//7zCUymMQu6RsnINGv23Gp8m0u9g7KatgjLS6fz
ztiohM1iWXMD+dVgmGsvTSvppstXSZ8vMNCVALt6idzfx+UW6Xv08Zk/hEESznZbxEBk5wmM0efG
kGbfvXPRTsjRIQDzJrAa5eFhXu0B8IYSVEgUCNy9UHrBAYI0QE2mqO0+YVmy6ffN7m8UI2Qldu5Q
z1Mk7EYoA91/Eg46rgpnSxZFcJ0nqaZjgzgey/5dxRd/JAGlIdL2HACy9dhG5b+yl3MWUzPeG27y
ncfP8c2L6d9snp34Z1POUR95zdCBrUDC3gWw3aoBEEDw7RuTsJkV8w5F7QaafpG4SYeMBQcLsX7B
TRysRCoCHOZJj/8Hgco0F97ulVFZ+JMn1PqdTu2eVfR5zIIT8+I9MaIOfZGv5ZhxWv6bdgSEYLCH
g7+d1Sl/uyNh6aNSteHlce60i7E/xE1wkx93bi0wRYVibrk1cVHmK+TNNzEs1vTJLPhpqOd8rV5E
VCbkmLffV0SErHGKRIWStlyZRrft447BMl4MajFslT9DWxW9WoofOmt5ZCdi5d7Ws/NFKucBmBED
a2wbi4gxLv+TTqzrwCyOsFqYVyXY7F4iYFsV2jltef24b+zMZTmREPRmPqpZTBAOdI58PPf9JhTn
BjCXNE8FUJ1By7XhcdEFeBS7PXpVrDKlpr8pu7Lr/SJAzko7d0cxCaztsDPbnxpH4CCNu55wcxem
2z5BLRNr3jTCtBl3c++T7uRC2NQ18+isqGw5ti2jPmoaHM3Euy3Nb3Cc8GbZIBbgkutgJ2MzifVo
m4LsfU7UbdJuZhbV2J9TeFaoddz8PLViyIFztnXgvGju5KjZAlzGJxzySvERFple5yDh6qxG0dN3
ULqg18eTSbD4E0FyeBft9W3nbri/b9ofh5zPZj0Mh84dLVZh4PyOwsRWVGosdjnCgTX2k+n6dvKR
swoDbxoiiId2cTq4Mw4qNePwOaIHDvt8myf4gae+g/Tea6jMWwJE+3m5WGHxsgTaRGnbTmx5h81x
0EYbcQ8J3kqr/z8RfsvlyRDezM6qCIpgcwthsU6AfJOwpHWAOIiP7I89nez6IxEOtNPIac8bg2Vx
cLm3YNn+5Xe07t3YlYnKlGivm+Fn7YYqU6En2mSCdXdiCgrhT3CSvhVEReX/63m/Iyg5+ugt4zVF
MRZ4ub/uHfmGe3YY8XGPdYVwttQtw/ccUrMlXJhIDVX1EoWYF6Ivuq7hM9XFevjyTyXt7WU3HAO1
M03fY00FR1v1tdHIQv0+jWJZVAaY/OO+svgO8934S+HEJEU5jJBN7A+RMVMkW/yIfnM0JooPPDon
sGzedVKAQl4h9xUYYRgXKpFlfc9A205wL0+bysDWHJ7Ino9L1Vvjh72oLV//2m8Lzcu2Ims22Q1V
ZTXbHGqSBRRe4ifdJ2YzwrUy3cAsT3T1mqEgfOhR0tU8mYt8hjca8HH1mdmMtSSJF7CTaoZeP2ik
r+crZzZLjD2Gd04vHGNJ6JcIVhjVNo0T9wXdg9raNb5uF62lVWk/fW+dmCbBEV6zL2SY5NX892DV
MGKkMsBCg87/1VjcAr1aLItip+svxtfUU9A1nibbB0nEJ408+QeObKVnzJpPrwz9y6Bm3bnO7eOH
cf0VNorLK74UBOE2+y2qfrH84AUvE3lNz1iwNyc976cLCuDcestmZfyr8XW7hAaPV7AGVfLe6YYf
bU5rMn8psPjb3XsJRWjXdtLrqAqXu66qysP9rmvL0dgAoP0v3dfRssXzYuDpYuzFfytUw8VmgBiU
UkSU2TUT9rz1471rWwEwfuYmshzo4S6176SLJSZlXgd3hFU5rBZSblOYRDeghuGFhqY/NRi0iqAL
8RsyXXj3ZFBCAkgtUdqypaWo+YCdkzzYj3xaAcMSKurwAIB7h/p89DQsYdWwfZ/wrE7h5qice3pG
1zLxRIDEytQToY6SRgIts3CuuvA8xLyLP7lQvdu46+VXAuf9iGTg5oTlJp29P5LmokF3AXv41Tr5
zCObMfOzf2/h/glqVuWeyH0m/eczyLuPczJyl+wOyIxkjB7JTjDkZ53ASb1k19BuchOqZXc8J41V
xdBhj96yRDzd6H5dcG9+4pjCHFxndcrLPLur+FwwhrD53cGZeLpwtFVV1+X8aKDqPeLJukpDaUQt
Z1Q13WU5TPW9gO/PSaCNq88BJwEq0g/PlItKiVEtiLt9hntaLCQQP6XNWCx/r0FH14Hp88LZM0Mm
+sOKt+pGo0IxTxgXHx9G6bgx2RYmlkCMFEFOFknqACAXYM3Z/r87lBpNxfZRvTW/myROQnpOtnN7
hPIG2Xg67dybYvH+i/9OB/cVxt+S6uAltcqTE1bUAgVaGPNGTOVFbq5ZxlCBcf4o/Jk1TG1yxQos
xeYumJP7ZpN2HoLPN8kvoP//s52PXiZw9+WBpUOC8nfcaZa9hEvz7zW2eckEO6Ik+ibZuRPYsxIM
cNd5nfZSBd24L1dpg9MM1MQ4hs3RkSTTB+MMdSpfW/G0cMjB/mwTZWcmvPfvZdcjxAiA8nqaB+nq
t1OmsN1BoUAgWak3k5QqBPoEswQXolJzaH60dWer98s8AFjRqrsADYOCbMk+aJpIK0b9uhnUhCiH
2PxbTNEbivoJ5EEroBfann6jSgV5gsd4L+FjiKV4Bu3mCPxjrEcniVW9VNlnqRiIRRy33PelwROY
gO6mAfLSsSMuNO4VtREp5aew4ce6L3P8Tm6za5Z3Q2aoPYoj5TYk9NqGtSo4RxlAuNNlNtTKXgek
+PCbulwGy6B43izGfX6DcfsvJVUeiXilNoIl7SFd9sAuyRMqMq22TNwLu3nYDh2OKvoWhGp+aG9B
kvtOa6ISHXksvgD54ennVSVSRLKuF+NNj/su/6oUjYjTTLMpgW/5mThklFmQTRy0zMWjbYrE+0mZ
mRGEgYMUfYVlngp7dQOo7kWBf0OYv6oqZfNx/dstRHb+nT/WFVOC7WufLGkFB0uaHXFXPMuvnyoU
zi1/FKn4aVwm6yyR0DgTm0HDiVlRuVnbEh2rYKccjkXS5Bz4Lc4ZvfS0EgjKDKF1dxhpRr5xMPkp
TwDreI+H+rcz35GWVJFbvfuhX0HbJfuHqv9wpcm4QXZpbZLxgw+ecIL0GR1mJ5HnZxKYXt/ELnot
B+vALE15mSDJ5YCP6tfC0/49Qn2Z+j9hA948TUJRnRCqj5bhHv8CNyrXSe4CYZc0USkL9D7N2n6C
uKWL+s5uds/hd+TmWoRgCYQg6StmqqIvDYAZDVajn1J63zEyb4M3dMbBpxT5WCV/pkP/mgOVtWD7
pDp06Qe/LmDBz6VtMELzcBv/o1fca3divJ78uxD/9PyVz7uSkA0vIBCePRO8fwfBoTiYwy4mL4Hw
cJzNT51SbCPvhHdBBGVvnEdCtGs2DaChXozUNq7+jil8dHelJgSs7XS4Ou6eGik03uTIcdHh0EYT
rh3ngJ0ZUHac4cIYsvOq8JkWS0zZnn56KDdbOD+crrcv/KTjPqHu8Rgc1ekUkONAR0ffhjhNXkHo
2RgMnuG3ehr7NRsoC1A4LVNVicbFl+eI+feR9mlfmBmvlcA312ZDaz1zU3/P6fsGch9WE0ySRGDy
CQ2zmZVbVv53zRF2PZawRaOc3RDPMcV6H3cCLFTlQ4LLSJ9vr+M9w4NQXfvLH+ZiWGfcdhZd1CL8
0pIWreHb9HyDnrPiek2vdzz4f1rtKTvS4MnJqI5DU5uuTShKYITx7mdPDW98OlN4vz20sHrCY9JP
k/T/xxAVG8jNKWNFiwpzi3I3+a4JCbMvcOqGKXy/jrJCUMN1tHSI/CjIux8KdXYgSTCKO73728b1
byus67rSMFiRDh2hF+A47EnjJzfZtpY71boV+7grcwINWOyH21UW7Qv7lGilvaIIEHBZt2YItxgj
XqevOQMMj02pRhW5l1Oe8SUrJdBU1vju0hVwKMKjjLoa+WHQQfvGcJPlxjL18Yl4fzeH3fyDtB2g
fl3o5c0h+agpyTYzD/pH5je4ejAkPCyHBpP7qDLNFs38vUPqOM4wgSatpjRHjvXyN5aK0zADexiF
djjKR/SczKGXpSV5+JathtEX6kVOCFQ5IP9S6k3YGbvggvc9If7fMEy5l7j7q+DVzBWK9zmEjUKH
Yx/nCcIG/LOYWv/ifg6qp+Y8uFKRYwm7MHdAIRtPX4qXAZ/zAlc2ybao81/oiJOaGLVCfEOp6G4E
qvjnyKikxv6NxU2e+gFtKX2j+o+9gRQfUOZtIZ4ypQB7IfyBwHfLV1BJ1DfUzLrLnYKdDiGXpYTM
ylJqyldw8jqef5dAx1Vs1Hy4jSJ1ZAfpOz3EbWCqboOuN/SXLuVRFak0ZNmnY6HeRGHfqaJiPSWi
QdQnfz7PLsb0pNPoFNBlvF6SZAbwDd0ZN/jrbs56pzF8HUDb7R8my7X5o9GRO0V4Co86rGjKOvwr
mp6CLfJUYGBtXD9sfOm0cIpG2WenW5a+NgpswVW3pl/HmP850oCzkoJbQRpPn1H0AN+lpQhbVhkl
vAgleFcKHlpebwDfDfD6HpF/Z4J4pQxdS3l28CHmwwXNpAF3uiSdlj/mZOsLL6JKAL4QJ6ixhNp0
yTjazX8s4H8javLoxRgDp6yB6ZGeGMv1kg6/Nqx74hy9wi+d/Mq7RyIu/ZxC3+2/Ori7xCo6eaUf
6mZDRcV8JAygSMg77Pc3S5pvzhmaDwTNW//nFeNDWELgs9qHhnbpZYhtgYPckzkZkHjeanqiSaHj
H/rWAPbT8JMA1Bw8/aOVCA42hmv/AqRIdOymh/GsSJKmsqLg7747aFI7aQNlF3k87/032FfdPBZC
vIxs00NYLI+OVmnOGHiSQlnN/A10Zv35dnaVaGZoiXIMg94TjG8XeP/5yXS+z+M10JZZB2PFjoRo
AZjhMHeSqEnJZznxnuMCWOL1ynlDdjflftpFMpjNfAVATa1AjCl3NR3WYZmLasdDMTeWAgUzX9nP
S8uE+aYX5nxyPlnCrNOxSBKKpXu02zHKku9AtirTc3WCEmmT5teZwA0LeEuU0McXVo0RvjJN1LEC
mgU8zna9SjOkja10jZJc9dLetLS48/tW6D1iIsSEVnwRnA8tGGcn/1ZVSlk1y7dai+QovgE0N4Ap
uJqYUzqi1tVpzgay8740EL+3U9RexAmYod/wzl4bCVUmc4p/NFGFODhPiloExELKpRgGJW69jC6k
uQLXCHkcvl6TSlOi+M5t4sgQQcuXH6u6NiVQZqxr09k/4ws9SOwgH4hcvS0aDSP2vuS9PFNwdDKV
m7IIek3S7miewMwZIoXfLa/0/UDyEFB1v9KkSraV8zhr3FQMMuGA60wUveHzsaiFvzbpXo05T5tI
JhaTVQoVPVV9Tncpx+lj6xsEiKIaSR2RXumBMk6apDwHExG5hfw/RGO9VBruK0SuHVhpNc4RWUn+
x5bMB6PJPF+Wn+F7CCb+ws6Gqtt8jOhj4/GH8Vv2sY44omzXX3oXJMdmkNTsDhF4LOClhB/ZPGvr
BWHYhD5Q9pjsTYcdyXZR1CvLPkx0FvCz1BaZfjU0I1No9s1P0EXuqXCcvsRUJGIi7wFEwJN7BSgD
CjHcMZQ1O/BtobjQP1Gi0lhLEqa7j4Nb8iISPzhYcvgc9vvjjaC0zXIlTNJBUmfxtfBEpdN0pVRk
3p3OpNa0zDp8iCarW9EnG3nBByL1t1IYbh174MRNCD5/aTXFNeCv7YOOUjtGpdJK7VGbVjwv6dpN
7FLuWKpVxcrQu84WUsvuQAqnjDqB6VNz9RAIcctzErf7pzByzVEL7E8ADoqda0FzD5VFmOvUHS1d
t1qg7DyOBqpP+PDqYqw1wA6weUmvBPBd2/6sR4AtE4il+GhK60tUHPF2oQwUDPIqTxnu4vBmo7ZK
HDXKIochR0OfmUQz67Q14uAsyBvrK1EX9pwc1wmNntYLSP8Jk01uIUaRg8TdwS1UbL9Yl20GmNMe
Yn0kxv9D7X8gr2wc+zPBnTIjNc9Lnq7leW95m1Y/yTS0j4rchf2javv8H/jv45utjOXgO5kS/2qk
IgBVCV8pM/ifqMNXV6V+d/VAPDYRoWEZAmlfEyN/iS9hRmEXaeDwrYFSX/I8n2mUIFdAdb2nPbgZ
Zhi5zlmo8r6OcCYsMFhFaGQyTecErYTT1Hmo7Es5uhyzjCWeJJuXeRAraHZzcwwjFALdDsFsVwq8
iBpv+En1bkf/n9SJtWGWUohVCLmbZ4nvRe1bsZTumN/nvACeXcnLMc3wHoj5k4bHGtCSIl499hNT
dzjH+mvsoYMFjD4MeMfvp+zcebHMQ0tOvCv1uCaC5ic8H3iFKTNvc6QNaIe4kHq8wXcMqkxkms3B
X7KHFegX/SeIx6csrA6bRA1cO14NeGwWnl/JRsTtAqgZf85pO8q5qVKiHKJquBx6A6gVALsfUYAD
0cJIjAxgHPfJhZBOn+U8u6EwuHH8PnKFb89Wtly+PmwVjSdb+968Qs7Q1p2hg5VDiYT0j+TNk+2G
rvGJj/R4VOBuny9inNcTtdqQ7fd6Lu4aqAV83v3DmwITCQCwVugtR9DYLsRkPOaZm4bU68B3kHdy
UhodyZQqJR3CpFTgR9yVfYQ90gHBkWsV9iEmStiRldxBenCEhSXhmXST/VC9JU/1G0MGKBOcdtSO
0yK145WEPJaH1eSWCxTfWNw5Gyou71UV264pgOqk72wO5z+VEv2sZ4z9fPfDZvc/P2YsgONocUaA
mZDUQBQS7+GnagA4+U5m2dX8DteDHFNxMOKhl7ehNvPNb/muferJ1Rd5CckhJcKzbivVa/GtadAp
GlaRH2ye2y/bUc0kMIZ4MyV4ZIO0C+o9tF7jfjRKv/66AC+kMbZ2gLjdVNwKgihlvkZcn/AXNLFJ
GAGJmnozi1Ly66BrOMg0MNW1i9XrAm5/WUtlh+JpqBZspkCDqqOyhiiNYNn1LBc0mMmXg6TSy0Lt
egA/tbyDR0W7LdTe6hscWwtl2NR6lvdVKM/Qv9YDicW9GKFhJnfd5YOZ4D9w7g24mh4QQNozRb1A
krkxVtOBBYBueSoEkDPp66lspDoG4XRML6/W1gZE4510cPpXYxCmMMD0l+1vrCGERkML4r8wMgv4
l+8j9ob1Qp1y4eetrVB9xSQTzs/7BW/0HVd2uLoOEYyTHUh4Za53Kov955aLNJV65f5bFlXh+FLt
0ZQv2SbQh0XsanwVOEwTK+vDWeAJE7R7gAfY575fsdcv0wMnPR5AFRgNSfbZJAZxhpf0IGjgy8Np
3qxgnQng8XCwjRe5K2gXFKPWqfM2naOSywyWRu/4qDDXLPBAwcpYtXqiIN8Q0G1ayD0+Ko/p+JP1
yvDHjKlpXUjVcr99ydbPg/VgFfP197AKvtaRT2eo/7KQYRvfCn8nYLK/dsmn29e+UNWaf08V72wn
LV4E3MXDWlkpKTZpgOddYLc9PVYRle+wfC+kcOD/m+qBtUsxYLvOegoi/oeyVYNeTyRvCANVrxOM
IkLqL3cQFaamSsIPmdvqL5wFXJ3suWtg0QP9iNHAYxcyObFXSEI7Il/OBe2uTQqqkQhv3IdpecI1
MqMclcMHgvzoWr14Xhk5bT+MzFl9vc0idO/lkbSH+R+X//cRLUUPN5JXBhCM0lNdCpXr2SeniRBZ
0Aypjl3bGRNcgUD7GGMJz439TIe95KMHgbllujpEweZ1Za6/oLJKWnvF2SZ8xBfL3DZ1dwRrl/Vi
cgE9+/iuoFyQMqSUSYUumInCbzj5e/ggel7oR+fh9SQzVlECHCNa/mZ30YGU/S4rbblNcQwUp+XH
Un9sEz2ivBttkOOc8jQiRPDE3x8qfyuJlfTcaKlPUvJJbfF3MZx8Eb8nJFe6e6Pr0ljwSWQPcRn5
T8hgr/VG1tOcZ9Zy0nohLtgBa1wlaw87HGwN8meD+ZBz4Cq1Yfc8lkbbjhbVfvPai3cxvkKp83ci
BGbyJMjtMEOXo4sB4g06/DOcup3/Imyn56uXt3iFxfZyZBhDb9D8MhvDKAT9hIc4aLV3eAtq/EXD
o/94Dx+nz4uNite7RvvdDy/Fl1Xv4kNKZkCK9c9oy65bGNhlbQIaA3kYeiIx3ORkIsbxV6B5zUND
j8kQ7yprrtUIRerB7NecpgFTTC/I1jvDEWBkVkbJ7jXBUUsWemBY+1EH+1YeKFivCz84HXAckIVq
DTO9GPZSdFsOZjA3hPNjSV6QCD1t8e8xZyg4XfuWRU1J27cQncbElpmX+f12RsvbsRRN1a45+wCA
r7C1zvVP0a4m1AEXalwGra9SoFvHz2CND4H/sd4DAOZ9K92xaIvQ40aPB8SFxz73cFx4oIxXlAgq
eCb+POjF7BpRdx7ie21UDYRHqUR92yxEWBwQtLKcl0xJwrIrvISbiTKa6n6NIHjl6HkgMxAzDRS+
mee1XC9Rbx54HIfVV6d7w0FeXDckSIo5uSYPqia5UiGNivbTaMkd6UEyyu4GjVkVubDqDShhRTy0
0P3vgQNsm5C+XDxNtFYCpHhgi3J1/8Le3vJukf3Pnrf1t28WFTD1boyneW/2tMA909LWyTzwKCPw
iKTNweO7GsRJLdDU5v+GQGJLJmnS0fJMmKoxLYJf9XzJ367qrSw1GNxdb1nYtX0UjfMVU78FtEoZ
Zxsh3T5pAz3H+QdZv0e13Y0DtLWyX4UPpIpFs4WSgjL79gxyc6fa6oEsxk0xhZbtoRvCOlGxtSoO
BHcHWBZXnOfLJ4sJ3iy+jrZZxJn4dcliLyBpzo4+6QbjKulrscLx7REFke+QQBkOjqmWXKtnXp/E
8GYYZPPsDZkR0w0zNhWDNbVE6fFtu25mlm7nhavUjsPSQWhHYKoFWJ71c9vWXHDFcaD11Fgir2J3
iA2X8ZsUvCv1Y+foO+ia8961sQuj24LvoskZpxhLOJ0jAosdEtamMDnO7ZTV7uNPhgJfBpqdUHCy
hJbomSbkRD2xtb0ekxcbkTrvsCIdIJ6Ot0oQ4pBslSYcnkB++6Byx6m6q0lfYNTMfe0GjfwFhIBB
VNuXLIQRkKBpjZZQ8hLT4yJan4YAckRnw48VFs2sgVQM/i8omgENu8JOUsgeSPnslUIQCZCB4wZP
5z2BsM9u84jtkZdl3P2GDiEonN1jIAyKqggW8CAH4yXmuX7+9Y67qPQ6qNDnXtCgDxnR0xHvdT8t
nApcf/vHBnMToYmXl+d/8LoyR5EPqJQs2Sonr5wMY2UUn8tkeXg4OrIp/sLEKH3Lh2NT+rnOSza4
0/9qcnLMj89Rnx3STkJLBZMZ3PuqFlcu/ZDHtoLWpmuWJdXOATArxooyZvkNs2u/T04dKrKI5v3V
QpqQS1q7q46vVMVBvakgZ1tkZAywKOwCRMuTU++eCViHNBfHdN6JdVB0R/F7AoUwJ3pjsiOdLc6c
Z2k778Vb8X2nUH0YcswpgVwmJqsxmQ2pjvIKsb7seLskUX1r+zptA1hcUX+xEQhvZ2AuUpBdZbUh
fVeeP8vHyi+G2HX8LIi/cfhIvwef93RrUaNkyCYQyXwXw/KAGrLgHhkRD+HWLiwhKnZfmbMTOs5b
T3XvgARdD7FJwybeE4miVE5yR60E5b7Vd0M54C2oWa8DRKuVU8shNfbvalI4C1II5WREh+xkIQ7v
2w4qfXOCjsnoi6VIeXpTL9I7ob/tPVf+OhJ9NTlBhwHliDpYO2ZekKiaoPME+ipJaYB3NYO7NnV7
skz38/4wZ8RrWUKjDAmoizzfb1kTUEMmj2jOgwV9VWaGHad4xNue74v8HtZknXGJsDqtpJFZdDAp
W1w+1KJWqBFR6TCL/YJNUDAvHkfIN61v9n0RFx81eHPRkObuYPWfHAu3+Tei5c3WhQfC/ks5YSg/
cJZQ4ql+cMc6j2x3w0g2yuP4OV+3KdMNwcnGeTMaJAsA8Zqgog3yNlL0wVBlAZB72lVF+JkjgJ9o
vRx+ZlcxZOXAeB1vpqfdZpGgQb21qAy19hj0CG0dNMIy8iJ4p7o8e5GgtQErbkB7Z6L/H+xTYeQJ
/zs+valkX/G/o+CVKvC0aFqPAu1J/n+TmHQ8yTRtADJUuiaSSoUAi9HDdX6s/A48r/nX+uznHubP
JgMaT9xeeoDq7o5ubRxBAQGq9aBGzGGNzC8BnrTkRQ6dmB6E0g3LRi0ElK7G1EEsG/ffeHSHqrSH
9V4WZAlOsmGT+SaYKz2UC5Jfp0X0uFNOzTOSCxnOYEbb0uwvNsRa0dKbh9lU9HjdNa8ywY9hw3jB
usCqjEePFq5XCZUJEq7i/4NRjB8fk5HckApxzf+glmwCPhzWEOdk6B6TC/rF96kyo3YVteOpu/KX
K/wjcvbavPhKLyf5qsjvCwQWVF82xLBtmCI80/TdbZS/Fq/Uq6idlhQ3j3uhTMK+kG74I72POGyY
SevM4hz4PSeiKH0+JbqYiTM/Q8pZfx38lKtNuDC11Ckl8+CW54A9RQWd5qmbS96xR78gAKYNk7xQ
gX+AG9oKNtWNLKWsxuXQAQ1zWEMdstpOTWoae5veK23m+P6qd3RiyrPoEtuGK0smwQ9Xo/g51yqL
J6UsSgYM6V3NEhmmKbW4cMKGpnOcLutZOmzIAbAJCFtjDjsQI9Q5oJVTkRYNiWO9Be2ho/l+UWUE
juCxkRoV2FW7MjogjukJx/7RXSmlkT0ZDNiRtfyNtf4lqA2bhUcGZ8vtnlQx5qnPMgjHGd7ejlON
B3MlXDnTYN1Ke2kPe1klyZvWcWASiqq9y8KW+g+ayrSUJmgXpSoR4VKgVPGdFXHANo5vj2Tre3zL
ihvLmokTDMyC+1R83eQkEBrfsXIcyJRUF4BC/KLHI280+wyklsyr8uv8Y1YkKh/h45QD1soDv/G+
1XuG2jQ0MVwg8ZRZUHW1s3WMm8I1BFzsNQ3gXD3ZkuLwC31VIqBkynIN8MzLH3ifFymxw9fgGBZS
X8wxUI78Yc2vPKPORlv2x/nTD8Ygj6uEmKy3Y+65+pMcvLQ+W31owa7NmYtAQE3opkdG/VGUnY6J
2FI1alLDMAoN8n3WdpIpBAAcylziV1AOp94B7nDjfpzXMP6mlKLfg83FoxOjFFywcsG2m2ytkWZI
r8iN+KsB0qQxGWzV1fS6cXHO/cIwkW4q5YAbhPHRUgNZJYj6lkDiFgQvzL2BxAkZTEeCyS5sIOuL
gRpD1eHEvsbZS2xjbwiUYE3mX3B/9TwHsWp7dpCqGk2vXy8/BF1OMSxhqsLGF/EzLejhRPqnz6G4
/Cur70WjGK/bRvnUF9IMPtlrEYXLBSWP6kTDJJmliYL4Qua2dEf0i/xdfwTSsO1dAD+sELaa7vj/
1N4XG6KmgZDIz7dylDbA4wP0sqnBFiYHcLiRl/4y8fHyRKHQ+rcxYMzTQ7hctX56aws3J1sMPpKQ
UsfxNepoEwMwGmpgiQFH9YThMlb1e45Ez3/Imv3SuFlrpsy+xB9EBABkEFYJI3XyCe06QNJ4Zn6q
MwTfo2733yh3TvTDId/TJZashGTUxJRI5vJCup6j25Hm16OvbTajiUbaMg1rEC+aXUPLHxAln1e4
kTHa4dnkBMyaO8NMysn9XYn8XRXZZgJxgHy3Xf1Oge1GjxhqKnintBBDEylfuWYLQtnZzdtpA9U4
EbomDwgJ3cBT6h7dQIFspK6VZgWFpZMODQxaebRgPcYOWiBaJInxQAX8lCrW5Sg/bZCRx0UQirL9
0M/aJeyz5t3xrKRTp+lO722cZeAj/5S9YzwUGjVDKkvnWWiEYu13L78jun9V766kwDZLHph8CS14
CdcHVKjbCJIjyA9sWZ5DuyqO5ldMctsE6bfLEK7Az6dsFUVniN8XS1Hnt+Fp51z5VwIkRRH1GXvT
ovW8A7ibmMzdnm580KZxR8CeCWMmBGr74imBOq5wn2E0DupOP8iMGJ6vS51sPJeyUFhSRhnJMiUE
rJvdRR6+iIfgy7kDcNOofu2JJm3QREUqTyyVHRPudhJ0TMs6NgMwKXb7QqMPFNmiCPDfV05Mstgy
nouM0KS+C94SNv5Ie+A8Waxf92DRHMbFBqc5kUsnB9VC1UsmSLJo2NOYNM0DtmelXrmlDahf+QAy
c+Ckh23JiI051OeHoQLyO9iRcBHZ1VcaaWKlqKGG0Fxl9jZ4y0qPdQUpSuXHhi7hQKyfaSyEfbPz
yiOIKi9NJUGMfW7wUqX8KhfKhEeLtMRtUK1CcK9jvioDRxj7pqbSMQ2/RJrxKJo0eWF8lQFMe3Zo
S67GlWYEd67oo2Fb5oODDXEM/bk74l2HuLQqcTy+fxEjphBrAgVgM7Euig8xHObvED9rbB1gE+Wq
L6nqHLSxKCrEjI7VqDrMGSI8oDOgjIyZUypxvBbPr/QzTqeiUXxnjy4pHUJ/t1x46vezIWqKrsFI
7N3yz6wG48sZtC2VH0bk+fs6JB6nguCj1SZU8tw8TKkZCKiaPkr517IDSRc51CsmnxlZ4Vh4miob
MpaIIpfs+RdoFsWH3G+8RPTGtBISp/9u8R560D9ZNFN4EmmiA7NkR/BZpwpAdgJ4U9g1GtyRlbvl
nfGPrQGChfmu8rXgWlHrBrbQ8xHVaiVVCGecl9Wx0ubNF42G7SKrwjWhydNJPUE0XWtE1/6bN/R3
6ltBa8c2LYylHw8+FPCl3DHd79VWVYpZFSbnps9KKf8SdVNzBKAojRBaSgcdAJJ2qlM2ecdCswH6
uuL+hRX6l/mb5/sBX9qeHbhU4vtX2uccmamRqgATCD43vOjSyOgVXiMNc11RZrg+dnsw48WW+IzE
hULuRERUsxX8LYygGyZLFUD/e9gEe8H0Zkk4zfbia3UxMKMGawVBVpAjoRvf5kQLm1mb0sKTaTwr
N37Z4WPJ1VQTXSf8KSBxTlmMS5BEBfMZwUjdz7NzflmEDnBRPnTBdWXLR3SdMpnank4qsQC9Hpwt
glFmTokZQ0V1btyahpXb93vSJRbIhMwxv41b1M2R7sp5Kv1pOai1eIufc3WdPgxyrFfs/gtM7MNE
zoxxcSbIjdr3iTAImHQ1vGDhTfVZpU3S1s0dpXYf5X4pBuH+m/Pk5IsscqAJoVLH4LSVApo1Oobi
gEW9GG6uv++1Q9w7JhzjLXAJ8nkFxXmfnx3S+yk3bFOeXgeFxQJqpFM41liFpW2RSmGIkUJsH0QT
+dgUzlGEstuP8UUYhxQdNnbbr0SQkFXHwJtJVMlqpzJRu7kWfvno9Z6NFImlYNbN7h8KYECXyue+
D6RderEuo3ANCR3UGQQMFRqZ0f7HIIQGFOUKYB/snj7tuQ2Jw1ry/rf48f0YYr804JKY2YgWy7Hg
PWx+lha39BXnQ7DxkHvMMIWobXihtZ6FAfOSbsL22nVMF2c/gUIhy0hxVULWRQo1L7h1mWUfEHxO
IJVovXy0eWf+gf1L5F7QO0VcRev8vpnuGuCSeNWF0YvmdylsgsmPOWZLcwXFnpyrO5DgrP0jJ0Jj
Dmv0Jhog8DSBzQdMKSipQJ8mX5RrNjqKNjZTD6Qo5MLCirrLUymCTMHhFfpoySGLfXKXxrb2MkEU
rEEi6SuUGriCDvJYgw2LkXF8SwtC08iXWdh2jO8jg3foSG2pKAe8nbMxoLmZ11bdLOBwXzd1eiL4
d3zxns/V9iX0JsAuZp3qN3IGyQ0awS8TYAVatDgugSTxnta5OjNHM23sd1jXu0Fe0NqZwa0BPfWi
dkb4bDulOIF7Nj3OHNCQbYygBi7GwtV2V/8zCTPBS1tqlZsCf2ryj7Bf2iLuX+khucnVM9AqOsdz
rYTGBGhozYkV5bsBitJqyibLk68ibwaGBqKYj87HyTIfQacXBsoMesVsFX/ID4Pd99V3DK1459In
wshjb9N3WJF7/qNLjfdrnq4FGDbtzngLhWiNe5wAbAW6JJurtyO8f1jmXlUsDEryG3Ah3dPQqsFT
rXQtLaRDRmZIRXoRYoOHOj2vE+63mPB8/3XievAu6qYp4LgBKo8JITcHsO6n/YnVjfbfYvRH89qv
BSYhL7wdm5rLdqJZtVu3CGbqdjT1cCBSsDuDpkLECM7JSzFQiTiR5ksO8wiMkrRPCjD2bCtTWT3F
2Lnncd4CPiqy/c7JFe8UQWxVuiG3d1YQtVP7xsh7FpnLnu860HKJM7izNvodRwliRUAIdZedoq/a
GY07rqXdn9OKP3o+H9RTowrYxXv6dUbNU1/jU5nHvTX7/EUHV/CXVXrkzOFSjvzBEFYEEZ2QohLO
p/VQcWyoftOIkHZuWeYDKDSO/qiIrI0gSj5x3B6wVYztTeTtmJpsNbAwSHW2bAX7T2ZXLFtFB+dv
JB6j8aNanITYV94PLsWiPJFoLcfMPzi2ogo2xsSeC3a7r9A0MpoJlr91FPdcMC3ex8UgO9dVjRgL
iOT/OGeXBcclnsbjPm5fZUQVdtnis8eaLhXOHRqmKRwBhrv2QBgw7joOlFIstPU+CtRAinQKzHvO
81gg9Hax4lYHxW/tyjFDbvDmxY+Gv2YyIJSC+kUuuPawBssXZzqS3UaKAIA7xmFJfUgk7LFBMTPU
v4FD6QRN/d2xGyBUCJ/f3+WLzejfQz/1cOLkG34TQKAWjljVY/kmskIyKl4ejIanfjFKC0HBYaVw
ql1IB4YgIus2f3LIuT+SvPCiAUGMKhv1EgjnqkaJjmyimGdqB6JMN+nO2yR9ECMePxTYFD1bLjqg
XrkKW1dGyQ/7ySepaUVsocuS9ScqLOxj87pYqKj/2NgbFHuhWtDMVA2HpnqkZZ1VmPzxf6ha7IVL
tAjKay8AA0uD3qPnUvFAyI1Xw3alLT4+I5IlbaQz70I7W9kCRRIalzuWeFWDzrzKJ43SlaSO+gho
D5Ew+6bWphuSPyqdB2Q+7qmZ0G9E3MWYHq5c+fUljnVDhNEPqiRLhy1rLmtFcxQXaHOuTmD7saKH
mkuFfIhQD3coZLddLSBwd/jpT7zXyQLm5rvQB+TJ9C2a6HNzcktIXrOUIyoAPXd04CtDfs9l6OPc
+ps8HvUFS4zMeEfvycpeujOUQf1F7ba7rAxDvxG4lkBpgiF1DJltXluAf8ViXwWkciDKzrdJKsrc
TVnx4gNsbGrloz6JpgKsiBiMfJM4l7wpM0IYXp2IWySvdC9KSxp4Dd/P/mEDZmz9DxPC3UAcURJg
Q2dKE9N6T/otA93+jMyOlp/4DlOOsMFrBw5dug01tvW2vOHf3MnK4tk142cLzjlk8NkTya3ZqH+A
KMb5idxD5HHxv2r6InHeYfo2CFxBQ8Rm0JpLSoHwwhfgDnrtxb+8l/NjN6C8aVdFAyw8qiCO0Hru
qFRrdZrATxFcB1AighcUHfzi/jmGzz9nWEPAlxof9ZwUcUBCMV3hgFVzw2a2rYJ6hfTRSeYbjphO
GIktai8ab1yPkVKN1xC5xKOP9/8mUcao6VoYt+8WpHb5l/8fJPwEE/SbuqV+KvIBYOyMKN50/cNr
VA24V81bCnOh9N2y17hzYT+t+v5eyCN7wseKbjvKzEF/gkNmSJVYWyzUHKC+CeaaoBI+FikKQpfj
xNT3dNYDIqFBvJwuaOZGIA8fEj9aOILdWUkSVkt8PU8Ak+e4DAe5IC2StrKExwmQ7+09AColXACg
1skXKjjUFGrPleMdTRYLCrQlXjT7O5r43VXgoGpL+9PaBo6YRKEsoG6Oz7jnemVAHD2vU21wLVuN
Y+fIiJ3uXhN+hrf9RDIhDvbfWE8mGiOfPwN+8mLNVAc8K/DP3fqeXyt5EpqhUS3Ca8EF0Ze//Zy9
8Uz+KXrTSATBkSrZ7U8rd6NInTRDrD2dmAukjOxH9dIS5ZOqmZ1YKBCDmnEhU83vM3F34F3w4rXB
GFzwqwJNGuibgXWX4SSgT82J9EbkjKjuw7f6npIvydBzMYH+kpygkYrX9qClD8vNhKSDVdHFFgXN
9xtd5PligwkfiFGxKh5UIbTfwG33ju4wqo1WluZhmIbM+Z7SsIje6Kh9GyA3Yf9CO60wWMIJNnms
uHFdmtAs8xiQCgHjxTS2ORgExbOrLzThEzwnnvlNXfY4wmRMyVWGSN9Knfgdm57BecLLiSIbfkal
WGLoxduy7W8Gv0MLyargh/ZeZzKPedDBZuCuVteNJBG6N1oGBqq/nlhIj/bu5z0w7zzx7xlQwgSD
dEXWNH2aDxN+CejzNDOc8MfpVSJou+QQ583prVIyjDLA676+seq43/5D5gS4nrQ9j/9KFlTSypH5
ITPRui2qu6Kzv6U07bieUU6nMEDwubhHbeUGI4XlirjBxIYkVqDWzUKHkBNxG37OD+vgDOaMezsD
eXmknd/cmZ+41moYVwjMhse5HNdMUj8RWEX9tpbTCpErvc9lxsfdFjuyEf2rM7vy6zyKnt0F055D
N9b+JNoRQUppyC+Q8djt5pvMHry7CLN63tcgMINhERaP87CtgwKYke2hsZNb4kCKajxGmcz3Bdp4
4cCQG/EZ6yDtuoG8ggzm2mS2Rm7+MCiz2aU5fS2pjksGZFUbb2+lWuoo9AyzX/ibD04cuqotivYm
f5ffvj0bzITZlKW5MR+lhKmaUGIc4+d/esDnCv4yAlHpM+AhscMqQzR/iLybHeoOKzq6nLFfEONc
g9Hvq113ZRl4Fhr6BBNewzuqIJtKR5/V0Qd8G+I1J4q+dXKycwqqOJra+3yrKwy8SnhIBwaOlANZ
WDNih2t0ImYZ+ebTrJCrdogF9EKQu8MRlH8a9tX5hsXGgopQNHQycVGBo4mVzkPAheCjVbIZ7maz
dcKsTRp/xB+v2f+wQ7wD8GgCmVS8G6LiiJ7OCsTEJlCP3VR6tcPMVJA9n1fAXgugpwoQ7GUN+Yuj
Be5QCGc7Ar85mvY/YU9bT6M20l6MHJ75HjjrNxPSogsjXy/2M+ocjODIVshbmY6uuCbjddSnWTn5
ObE9KI60NJFPoiGmrXKRMFXvhNm9dPxYHRmyc5lpBmpD1Dr5hw6omdE507xeNUp+MBot0xIs7cfr
JW+LIJeHas9PKnVbtKsbQkSxX9pwlkeKEBKli7JoWVA1pFoPaXCcyq665Yowry+Nf4X7+GDMVqEB
MdaX+lHrM0GLv/xZEYVIt3pGVNfzLBiqtV2gxR2l1oBQP2a+yaZ/OH5ScNP8cDqhA76dG7N0S2zs
qGbQRNGbZj59VU8S/cDCEWFluasi+6g3DhWl7/yB0ZAq2t9pYZ7/TAiMwl78k8P/3b2oj0xy2WAL
cfYpgL3R8//Jtd3tJlxNgKrp8HzUiLQPyuVTeMPFuLD15yHM7H8JCw4hK5EbjgJeLnjrieWbku6q
fl1U0QWxLuvdjAIt4Pk2QsIS5SW9K6ECofBCT7k5PThIcXpfxXCfWS2ssYzKUNiynlPAjANbE5bd
lfVP1R7Ba88SnlnmqtO1z/qmgzqm3L3oKwLFyi3/BGlZPbXRIC+auPFdvJOsjfNA3UfdTLzRFwvZ
H0zfxpEOL35ms8neAp7oB/6U+hl1uRUSIEHTNFACCOAdJXRbtGQzV0mqPM/MCpPv+GYr7MA2hLrC
lOyt5CEfeQ4y0beceP9CH4TuozIyCg5TjkVKboKCcKAsof9H6cb9YD1aCmCCd93nk8PPa/1UKEuM
P9BwgMwgvQYI5gnQ4Qh2ytu2UICpHjs3fx5umJmf3KZ+3kF2NyLSGaxM/kF9qQosegi1czOUwodH
EA9YyVp+xAS6p2sHThLmggRGv9YZMyr2PgOpcfF9pgnDtiYouVWvM4BwQxF+QFOpg7XdBYOjQCtf
SD+I7n+4gJIlJeS9iJxcB1KHh0DSXtl9hwRyU4D76NU0J4ReenF5y3/love2RvsVi2MjOYnr9lZx
NmpSEw17il5o1MJ3roKP47seQQ/xGArrqN/7tLKF6+9MWbcviCMmM2Br+5K4ZQfUWzzCrdDXB4hM
u3SqVLefqKgfswd3FilifZoClU5IwX5tpUquIVPVikgwQWf4TugygXt+vFppjEctzIyTuc5zV4uD
cQ4HZGtK3AjAyjyYOzQylNdOh+EUm0FwT4z9ngb0QMDTlHBk5o7tdO9AK9RrIKBy3EgsgPC1e8xJ
j5QG6iJkycoOrT4up0kr4PHG2C42pumU8kkQ+luhFP/nwQoUS+5jwehtjTsel0sjyIdNFGj/h5FU
vUmqE1KfmFVEnHjIUVWcjlZeWnwXIUj8ko4BnBJ9cwK4+Gu5PYP4brrg18asQXOxPuQKECd7+kbG
USCB6aanSkTiVQ6S8QJyhCFklOR2jK3ysn0L0VkG7QQzqV6SCI2w6a8PX2zIo0LSTjQQ8HDK0oVg
VFZcKbBIkhn0fSrx7Zrp6DIUED+cHER9PBKkbN8t5ANFx0mO65M7LDBrb7khF+deLMspXF7An3Re
FmKpTrZkfJ3juIUnMM8+L+bqq97M6SAPLaGZ2lrqK1czExgTD9Z8fXtysSGmXAyumdxF8vRhlYaV
CLLrgGyM61aR6m+/6SbatJ+DRItMVZJfqnHup/cS5bRwRW6NTspj6PHGcqpZrU+UmZYY9i3c2xgD
tYzX86VWgHQTVmIhV0hlWvY7NC4yXpaO1rVpCP2hNbYOz7XEqSvh9SRWlOHAJCNQO2kdGicLw1vv
EOPHNFVrWsP/dXlwy00I6eZNZ3B3hm7PUndtUCt1/pWuDs+HByX/xb2C11Q9QKz/XguPIMCyenji
EqKjSQd/8yiM1SziGRp21B8c0MQweLSk9ubNnmlf5783HoVhr632WMNVaON1Uedye6Pki1Lfs/oF
BHVs19iMcNjYOSCEt8HatDnph3PpzNCxGB9CKBWJfPGt6xqttXN0W4fA9zAuJD50uPjBhsu6baEc
SpwJuX4vTCrndHqPm3N8GRSpq6usZKxo0fe+XKciIyEi7xha4uCfU82aDl2kXcWQf48F41WXD/Lo
hjiW/uk46jsf/mkEGGvjYBhypU/5+Nv/v6Wg6+jLTlLXLwANYcUmcfSiDNmPJnHQFkox64GhyzT7
xjC3otFN6M4OuhClmYaoOexKp71UQ8bzrFNI6uLYo6ClxsS2L3xgitHs30G4etNdbeyLAUsqti06
SnNZ3ThWP8cf5/XEwHnPebdXGtNlKyWTc8zWLnD+k2nH9J64R7WknIRVnugEqbnoPfRK3m1qIxjI
GvD29gqnBUaVKJzy31RY8fEZn+SiTMxYmMsE6szUeUJWUhBQ9EXPaJRuDblEwvyGx8ftud/zBcHs
xxd2SE3hOe6pts66u2/J0UEo65ldRuFKl2EJdcbXjVNQ1Tjaxsc5HOrgA66X9ObG1PV3uz4pdP19
Kuqh+oicvlmmE6UTXuE3ImH5vZ8Ga3XSJl8GEYaOW0kjyJ+IsQD6a1v3E4hV2MfmFN81FfSuCHda
uI9cnPSYda5ziQrlfFAhJYRHQX6PU7836ezzF9V7/R7umTgjp+gHwUpN7afMory3i5BT5sYddwQA
r9bdax+9fqdn5ZrWgfYxcb7IbfT75IJ+2VUbJgm8YJwr5QjX2cgcLBNmswlGYC2eJ29p/msRKy/q
JRZcWHAtir6EyVrPU2Za3HRcyksrxBdPYzPFGTwPV98v89vZPiU+FxEMGY94b529lyJ5dBamKE2I
wQxGwwxDRSO1OFNbeuCNr9HAySB0Jdpr1jQGRVu3emGm6CUYupyOsE7Ybr1cWbzQZz5pAImN9A4U
cTKvWBd1459/g//YqH3/3vidaxnnmwiNNjyGqHeseg8vOij5HWItHjdikiw3bDyxHZ7SCoW09aea
A7IlsQWmm3BkJQdOOQ8h+UxlVW4HB3twMaPbeZieZPTr1Hxr2cmSQ8d4x5Nz29jCX8NYdq18I/J6
7sMNS14MBIU+lEOY8OhfBqs+AnWXj43jNzRgHLabb/cXGvrjKjfrFBTIg+Vp8shruVtw5J8eSAQp
n7GJ3htVWpKCdK071xPLIP7KQCF7rjCXUtBbN4yJwdbNNuW9sBW/Jc2LdxlGxeRDyu+MaX4Ao6SH
kzEZVK5vGI+vTjtWqFX9J2+D2JnYx52dHph4LMRgOBGWl3Eh4rIf5ASz6D/seLnO+E5dvVqUZQy/
/SZ1RCuv4LIq1oukHEsiyrF82CBKEd+Cec5V1qQNv1xaIM7M3XDeINhx6XeVCjWWp72cVFmTzi7M
Ei4YsggP7MbBNl/jBGqWOo1+6i01Ti94fpaNXAiKKFlQKlo0NhA1N7ogT7JF0guUXlRmtMuUwCww
fzKbVxTBxSur15jc61dcGN7HF13xw/HkF+zM4TGYUv4sPEu3YYr1vRKuqdd2KQg4vJmW/+gaeKPt
6QvqUSiBJ9d6MDt5SvJvXKfgU7/dk7sHBPklFuDxBFgW6dlJGr66D7TvfdSraRn8rqynX0oCj0C4
A06ytwjGXqS4PZZ4rtXjn23XR7WrOkY3I7JMfx9MOhffqiTrrq+X8EkHq3FtnZ56S6aLGA6g+ADK
eHfcqvAW+gXq3UnBzWZGYuJXdd7YvFUG4Z7DHXGwzwO3uK9qnNmiGQ3+jZ0ENUAN3RDysAqFRLI+
ge4NeUdi5njas091DejIm34qyn4kMsjA4Im1TprvihQE7kbQfmKb4gJlshgOl8AMnUcSC7t4v5JD
bPskWq94J4XpRX4gqu5SC+4JsTXOlLH1OgzjkW4opvxbnpkOjq255cIDRXiGDIQVjjKvK7flKWhD
7Vt2iJbE8MFDj99869FhrEPy6G5JY/jkEbaH9X3PFIzBxPu72nQ5CoicgXxeoBh3vn8gBf9sYg0h
J4KzOhziorNqQCR650zaUpcXouQtBGZ+tbWM04c0dzySTKFNMZMUz84b7lP1KY0pN+LSENdZTfdz
zPqmtyyLI4HvKnW5Ls5SMAs8vWftwn7bO6WsIDmNB3od3JPRhUahchu6DPACVamMW/Ij6kH21uBH
dpSJpg3dnY3ta7NOxoHotJPt29mHU17sCKeAWYEFOyAxUWsBg/3/ihgkG0oSG5rqcrPdd4k9dYjQ
c04gAe99QK8H0CgA+NPeC8PfrIKdPyefKPEcR4iYGHTwjhS56n74Oqs/SwC8yUAXc1lp1Fs0Pq31
xYKt9Hx1cbCiqpvAvmvb47W6HYkRbhOxC0E42xw7IQLMnvVziJ/TMQJSaeWd4dDzyEuer1qsx6A5
bPL7kv6ZUXyZY6WG1TiOC3D8AK/zUrGNQMTX7qqXdH5At7PuPfEzY4LZrfOiJBZ9sAan455+xJRp
n8woEPDTYmIYtIrCjxdQncTW9INULiyB20J0HlSylUYXfpujC6kcpABp4ZbZJjfNNwGB+PBgG6z2
uECISK8IkxnDWun72V6DBWp963U35mkFucUqUO0ppEYh+YFIEhdpa8wb94cP2NxntFIyTDhfl+Gn
NLiZNAmnC2J14Z1mX74nr0OKWm2r2rkAQN+4t25DBmKAcg6PIIAO7aj+HENaBPjH8TcLqNUpPIaM
YaBVmzDqbnKuLS1g08mZkX8gPSSogkQovDwNgGj7J8Uf4KpaEI6NYXyGwMYmSwRroTBRvApEqKw8
Iaepi6EUdLjZWCHlS4pl0/kehx1hprdagtLzdDvLhUnkC9P3h54At6jGlxF66jq9BRpjvbEOedWj
iCWrBuaqWHgcov03sjqb6BSHSriDdywZKT9ziR6g7BU/Srf7fMRnK1rV8R5faPNNOH4DuUK+5J/c
208k1Xga9tvNSWG0VNIDjZDYOz+Hy7oZlDIab8KmsxApOwei5k0n9Ooto3wh4V/GqK/Qz9efIdv2
lyIRT4cSqYZXfB45G7W5FiO0ls0LdvFTaDxp7JIQL2uEDBnZP0XWVNi3em8byu7+FwgJZw0gx8SO
DZNR1FEysaUGg4AFUrYgTxYuRrvLvPCb28hH3Lcq1/YGuNV8gQIoTYx8AwFiE1C6iD6SB/uMITEb
tYeKpuJpDZlxGYZl1gbMwbvfuZPlMUhTK4HPhBAzf5U5PfSVEh3Yymh+rug3MNJVRNy5GygJ46mY
iMFpfVrId7r00vgqjW50Ai75L2848boU9wGvbY+1aq5WzVT1M1CvOZfu+MizEyOrheeEbkydFdET
SjRBMCbscQouDaCzC0EvfTXUDzOH69JdiFekskwgNZMOMeuMlTzBVtOgcuWUr8lukKbc4shv8R+P
WSst8uBWE9aMigiFfGKm6ee8ds3U+8GFk1LwIYr1So1rQesnNM3nCU8vTkMOGg+ZyDJt6MrSPI97
5BBCF2VKE0wVEMqRa1543aQVpYIRZGpnF1+kru4QGWru0q5wTu+0gmYrOIkyre4TN9Xg2LMuACVB
tw3U4EOr+TF5pSeu9C+J4EQI5eWAVaEyQ5Hrmy1MqlzYdCYZwPEOd6UyN9ynl+7Z/PYCk9qT+smr
Fv1jPxD+RC030cmlmGikYHqUukcriuVnuACywo0DDF0D5TY7OqdLiqV9X7MFWfdO1u5YBN9OvSgD
BbNS2mdq8rRuehHkYcClt5hZIbHOleZtfs90zKGfSxOl9rSSxbqw8bdstpX9vIK9SANkNVTOd/T2
DpPd4tcWlZQbWdED6UwHqjlcwMFz2itTePNtDu1R0JWY5NGXy+jy92WvXXzir+qoNMT9YoaLvgOq
G8oJIzkie0gpSoBQ3gfXLc12bpIHCPTEsGOYAozHd+HPe2swB1nuTBunCitif9VGVMQM3crGX6hS
g2/Gfp9s1IeZZQ+TCgpLkLRE1F+OHinFuqQQWQqTUZiwRuXqV4KMPokcbXo7C6FYj2nP+74gGngI
3hoSYXDof2jwS93FSz7sIxV/gDwMC4uIaDgiu+kbOqkMCVvMKeXX5Es69P6THebqoNXbWQOHgw64
Dk1/DJoVxT26pkxze3bxt2bv4VPJtbotmZveXDNWAnneh+2KGyvXMFlpCtfTsaA/wjKlBzciWiWf
GaIscvqvTU/84AIYvZmukLJWHyLUdhYsubleHzAJCjd2QiOnaXkvC/SbPwjXmYMoQFo9Y8TbJD0D
E0LlkLfNwqvFCq9rI4hfGHevmxf4sk7VrIgVQzrGIFxE2zpM0EaJIDM2278Dgsv9lsgAF6WQbqqF
9SK/L+CKOIKfaU+gDkxeBasea2gXchdSxGJVq5PB8MsGeIJzYLr87IBnqnA59UObq/m6wTqSL0XY
BHg/dNLnKlojm9UGmHPlmSQW3UkRBIhgwAiPGHHHvQAMowNojqEeUENexWgTdv4mO0nvIf8BEAY2
HCExyqRFlDntKTXN7ICYUhuZKvb4buBbubGmIQfk9YJ+Q8TqA35z2b6FCJHN18WMyaB9etkasOmm
S7/tGgIESwIocfM6Ho7SFIGAydtAH46IeAadHlvKWim/i2bvqrzp4HSzKx1ceEXf/odh/87GE56E
1ZzkhK4r2yxn3Iqmf9L1E5LGnd4zVfEOkSJzwYljRptnGZxa7cxUJTWYFxX+B5zA5Pvlx2uc43+L
I7uwrUkB5LqWUOxa89dZWALbY1E/N4z/YCdt3rQ61KRP9BF4qIhQR5m1shfuMn3pzBA7PEJn0mgt
0ZLGc5dEYYaxU70YHAUr8YwDiQE1HqLkcxiS1ionbCC9DBPRhjhreUDq7LBtpP1YAbhvEuf95BTg
H/sN0TvnjndRNLSyF3X/2xHDjPuKkD84c0qo8OYA5GCpyS+6hmsvHGvMniNzS0kRFsOygnL5wA0/
tRyWqyFJC8pptIDUhMCmzF53TOlthGH6lMEcEfvm0Wsdm/DiZl5Vh/qG37rLBiuW1YrOalOoIUKb
pQztakACzVkZaeWCSCiqMn3wBCgMJWHcSgIcQpw6XjTIBo+WMXDhg7LMjZXH2OuYekPots1MiVyz
VxyAuBMGS1b011dhLpVpE/DdsJPbOQGeStyl7kbUAipKATr76Ms7QnNsQ28vEFVkNHlYd6rLN7QI
qfYg7IfGEeVKb2Z7F7TEGD4Ll8pRmOlUIZUNSFzod8iWiCC57xYXywoFWlD0fQVxeVOGu0EMRZu9
vxL7QsnZHdPFPdy2AL5Z+BEuHw3MXYpgLTPpGHowkTfQyhXwIIfoQ51lmh26CYpUZJ0zoEZ9zWWQ
Yiu+ScYBm7Uhg960JpvzEgqhgd9O1YSgMo4e2vJgCX+bSc4lWR7l3R2szou6ETc/wcFfjABOLncx
kQomixQOK2AylIpRSfk8teNNjPp/XNHbogHhsS4cqsAhlPAMPIc8XokZU9VYigqGQl3s4z5yj3Hb
Rubi0robBU6X186sEZotpBmETzOXfgZzHtlgPPmMRkqi4BfdtbaLwlX4N+RZbQUWrdhTrEstZSct
oU/ggilACuhmWLqgeGBCpD2CEyA5cRcQV7QRJ+pdJIbw6hTgDXTpbQZCdPfbKAydmjBETxdh+3B8
YAja1fLcRfWdnpCvqAITVlbj4CdNY8/az2mdYxtXBg58MIxsVivYRd6hJ/aPR0R8k2P5S6cBpHJ2
LCdL3fWEGd42+ymutkq/ISz6uB5Hy/vQgDIKTypOQZz7VVV4Z745R1iJ+vC5ty5rASaFtjbpnoR3
JBrMZyQOzzv3kJCWhe6L2F4YIkrIaVTqbIwZn/OFxcz63aPwk+780icXKUT64AUQEOzHsOVKTgly
sro0fdiByBegBH19RlefOQJOJCIFTXdNMYbCuW5yYWfwJeI6aETPaSPgdVmVGh/DiC9PuR2f/jI5
Xeu/PbUgklhmENZCvKi6239ZqheYNRwz8TlV2Iy+O+vQkFYmObabrGdFEfn0ylYE7i6+SBV5bckJ
2LcV5CkMAQ/cnYNNlw8J6cQUjha49lALpGfabWf6zXZ1VA5eftVjjEIFYQAzcoDLz2lZZ2YhinL5
g8ihk+kkzXz3u4jD4N2vLmhWzNnpxQ1tC5nc1b7A5hwBb2Tc6hAVKW50ZL7ZUZPyvajdEsRPEyhK
qWYxXE8RdScs8Bgn3Hr/+lbDNQ+8rDiqbP3clpKlGZ6ypF8Fepk4uxNfyQT3zZKVxpH29OdchMtJ
r4S/cxGxMeuXEbVoqDcxJbMdwnHI9L0hpL/maLQSiKI7cvKY1l/S+5zc6fxrRTVy6qCykdf8DL4R
KW/31t42PFUUkURab/BzAv1OV1sUVj7uspBOVuAszkx4mkZjMU6Bu2EbOHeoGgr6GtXeLSu5lcZb
+4c7k3oXt9rc+bkwLw5DiQVtN9+sBbuumI1L/Hsb8IqIRCAMsg5GsJhTnTTiLVlZzoKVJDu+xbST
VO5ZA9ojrKSy+vj9WymdMM/LQsZH+7UspUOxb4SFRA+E/P0UYONZMZb5Jf5SjfxT+uwW79p8cxRw
f7nNrJkPefSj8OLX4r+ad9shfkLdFxI5mkzzaML0SeRNUNXN8aKO6C3xJsREClHxR1y9Ikk9THNm
H85sM04JxKvHsAqOOAFZd7layfAi1npXJduSuKIUWzxz/rtwgmjHZ7QoYctJRgprbajVzR/UVnyG
9zJ6nP5X5SyCHtCNfuqaEG6kthcSm4NX2re3KclsldI9/VpmzqhFCGJgdGhgogQ3cBKYMDDDx0AL
qrYNMAT0i1QoAWlXTNNHy/aqRaX40DD6FeVhXXe6e0vr50K7EELd5vt+k7/Tfbcm9nTfCiU276Ix
w5l4SstrHjgnvFD8NJQ7DslIEaO1oD3F/YYE9a8chY/bwYh7g6dalqV+bdZfOqn00OXdaOyGiD2L
9sggd/VdhrPl5rWr23kHFhQ37d4f0yBqHz5qhCrAIhdZz6blqUJOvQ31Yhi4IVOEYHBojKUA/tgW
UWoyeDPaZ+s4l46ulZ3bVxs2e2VB5SVT0XVG2lRqwZnDu4gp2RcW+y6mJRn7FCJofH39dPmL3vXz
BDviFqMlWgn0nBNfIebbajklmCliiYoFfdtMCJr99GcErMahvJLnBI/rJLV63AHt+3XzkdJRoVVi
jzWm9l61pyeTZwMb4m7cnSsyASAQ68rFHTiIdmn1FO4xxTRzstCjFtgkEVQxaEU5jKALlAL1dr41
p3Wn53KI51WmSbNCspwFph9sRzi+qagCtJqzFnN+qOJSbcbosAebDou1Qi2GRTW3YWtDg/6HdtDG
7jz2Ob1oXIDsfNofmleLP0TjuYrrYytBXbVAC05CDycezKMroGp4zTht+Aft8YO6fF17KRCrXHr9
gAfWm7cznXiN2YowGB84hNZ9LECKYILEfT6kZICiOLucgL0AzKhXquYlcq08vQv1gUZx+OJmLJ5v
dP1zoIrsn/l1dzTRlmknBkETVynxjUVO2c1Aq9up9BMUc9GDRPNdK7UoE8QkLUL7PV30IL4ZLBH0
MRDQ/wBVPwijYgVYwzZLugrnJHibJieRanOBqLIzpzpg+5Rd1kSt3/VfMqpbjaoYPW+Ivwr1AcH9
8NkKFSoSByOGmj5tFno9N/xoIA/RvA0ToWDG0UIjcQ6tu23gruacwMlfUHKBDYbzr9u8/01Qi1yg
xpbXlf/8G07qMR4DehpeitiprESPB+61CV3tA2RiUP2MPYtZ1kvAaV1UFEKTaFe+3UeeLBki15S9
LPxpdUnVReTcDzwvo6g/e31ydn8zJW+TKDcAOJXpzzfWcecqQc4RksKYW9hNwOJiDTimcWjih6GS
YSOBxOM2JYvfPbJFrBfwudaymvJrMByn9xUu4K+Srev17Pp1+UOm1+oE9+Jo4u9lRPBzXCm/1hT8
HABvNy8nvJNlsyOK6MUeTCg/wIrZ1L0F0xtE0Rub5HSOhw71NtszpjgEFNbqV+wreKYI17OZcUR6
u3vxPpKxEBizXHv7/A1AWYZE6k9JWbZ3KdIXT31BQ/ph4/Xas/6RKUe7Q773JhUPMPlYhoYuAY7G
YUCRVMUk4mQ6NszmYaNMCWcaqbQx9MMiP0HTbLgPtdAJiMGmFZ02KaTLODYa+Tv3J4o6BvJkhlE2
FyRiJEWJcPHAq2O7q5IJzPtsXEtMNciTaDqfs3bF+e74TiLhjDJQeC8+JbsTV8WrqaJJ1ARc400e
1QrmayhdfeZg5BLrUOOQ9wShwlgtEJlpLjOOILbIKVKcLI+oJ0oPxO0lcmjlIMgNpyGeIWa5bKi6
Ac91hSEhW9jx47R1nIKgq33iMWUGLVpbmULV8Hf/R53KMH0EpAm8+Xr2ljdeO04042GjyX/IhuTb
DyeIcjSFLQ9C1MGg2rxyGGouy5ggCnhEmNsaXj5IJJAD1qN88OqXZWhoNK0vvQqBw555rIGbqWZJ
WfF/aT/FhwsK9lnA5Id4m+CtliVTJCMuGZ1gEH7L1H1jU+7+yI4H4xRRhK90GN4DxOovbClz4Qlh
nAqIZScE5Vbli0/Wr9557618SqR8s7uyBrOdudLt5WsZqbOJpzGO9wQYqjNGw6uHgSr3EWpotDcQ
6iZ1ghLgthIf2umBB3+QyjVKLqIpQGLl3w9f49z3hgMnVGWJo8GcFFoZWTHFmzWh1hhojQNpfIR/
wP5QuIaxC6nXRHVF6Gv9NePUBR3Jrj378eY8wLkJM5RKKHpJCtWI8RuqhTGmtGbWR9UaBf/rz95F
Hi++kCjJVSy21n66TjySQQWyyXaOx0HBFXSXatzt6kIzCDS4WhpFqPWxbwTtUr2m9ehVd1xbQaWi
ifsM2XJnk7YGRi2at4p+d3Kds8iGj86aawvf77+le1rZ6/ie/JJeBIoU6EnBDmZ2wcEd93kc3YIj
ws1csFyu1ZJCr46M8PtYW6HE3+KnQdkxhSEsKYZKaWzoyDK5v69S3yqvuzosFaqbjwugTHn8o0Vj
GCyjb/1jBClafsn1TGfxTNzsb4Tn0qe63A1sJa2bEPzwUYX5R2KlQMPIdb3zLg/pNHTkpysBR0FO
nbSxQGq1sDcQ0bmeJenSjlCUCa/8/fdTm6zxG0XORe/j6aY92Bp7vzNxEkNOwbUuHCVFzKevAs6I
X9dj1s9SXQi07M4MojmLEyZ0uJsaL/F8c9iLi+ChJZZkqA+l2z0oNPTaz1fgCJT98Ox5NYPSqAT6
i2Z0sKgVmxpeZ8cPVYWTTJ32XfvNvWFSX6KjSLj79kU7ozR8NJIAmKdMAy/sOuzljfl8yvLOe+eT
dcQk5+PgSeln4RRbeC7C8vpy0jHFIm75g97cVL8cNlADMq2cMEy6Dedzwu4IRuUwY+0qEUemZEhg
uPDjzJW3vUjbnzTsWfYLQXH2h39Stq/6OcxGz6/yG11jcKu9dod4o8c1F+4PxaLgqNE8wz1nUGFL
Eeerm6gweFhm8FP0kysVeMiHDTaaH4RrhmHunlFl2TBHVWJzedjKU8nZ/67Xcsvd+KZYtvLqDvlW
HL0zEUCC9FjuIm7RVO/Kq47lT7Mkg9CM7+BdNEH+MzfHBrEXmMZWq/3RobAgkAfRtd1L6KU0kFGR
lckB3nDB1HDQ24mO2HowjAD2ZpMrCAES2oryg2Owt2Nkz+CFgVyHTQm+QOyOo2se2T4e3hkAyQLI
lr8UlHisBOR3s0V4PWk7g6Yas2TJ3pIQo+9hzXwAEKcUhFIZjLrpZM0dLb8PwGyG+yU134VvlAG9
sgf+yUNLaJpk8fAYarWXA2TMCrs9CdEas12Aa5LF7Ey7JUyyrO12cE/Rf3T0ipy0YLGTEjZHw7o3
02U/+1ZwlRfriWzr9U8lQ/gCc+7+cObeEFjGl7owz2y8I2jQgd4H9WfGghB4JX9pEzmK/OR/rKyK
iZPgLNsmmCi6pXkbLwBCTxKptqf7onknBdnkhonFLALEHLLyYCPN8hDKnss1c8aN4R43A8jWIoFz
M6tfUMTtxz1ficm2wl1bD3POk5fA5m7q+AyWlkPEV1VUL3ZKTOCXKjcm5+N/39JiMHm3l7w7yP+a
k9IE0QVm5tY+YvgbxX8YFXOHxe39lDMwUR7PesqRY8TNdRieeLiHCUQKIv0WbWY47IPyoVi7zi42
Ylmhl1tWDDDMP6FZq02J9yU6IVOSDIbGrT4JecDrnlCnqnH4v5aZpKN0aXCF86CKlz8wwfEbC/ig
1NUr5SHOYf1mRTZszgGhfpS5W9ho2dEP12wLwJ2Nk5bXY8LFLkp6ziLM6Z+2gKnY1P2YRn3LY781
szNAe4JFZmyFvcWWyfymgnx4qR5OktQQMh0xXyqSMwpPm/5mOMdf+VWIiWdz2YKO/QacSDS5VZgt
bbTl8qEl5BZNuWbRQU4LVg1YqTBR8tgjOnvSeYV1ET3eq6um+NxUmkop5cwiQ2T/YXzYa+uvcim5
ugPVF+Wq2ouK+JF83CSQZ+qzUq+8sxLQeJfP6cflwjSlbZ137MYUc/yPfOv56pRXTC/hj9o75xBp
DALjW6zsJ61CjiqttJ2T6SVIT8f8fFPiB1pBnX9ofzJ6CF8ZiXA8vzruJb/M4XzXV5HI2nmHRbFh
Zpgmkbiwlhtg0G3xvLmexSy10Dh3zCPqmQiJCVw6wIU3NKD2OBRvNWYsQulOcvjvmJN37oYelIoS
4PE6WP22TZ7axg4r96RCQ0d+maRl3QUk4e6HuF/gvBQeFqRGhg63HbHRvKx1LZqR3mk4ypCYB9tU
A6Wg6+2cz77/YJnuo4d0NQJ76VaQ9qef5CLrE2lXcogPbAWuCzj0BJOhVMG9YlzJi4u8fYR1ksES
0CVWicKfOoK6PdyUOTxtSuvHfd1P1RJG7WGJh7jkd+6/4NmWvvdIdmr1GCnLY1dSkxbzQ0WcTULR
TCwPgiPMnJIVWUdofPxaXxQlwZM52nqi1HyAvGRcc3RZI/ilkY4e5Rh007vTimxCiNS1Rxxt5hAS
ahhOMVxhkik1GTzMTmukOxTElNsdFaTH9pZ6g/V+NxzLfGGyGTMQOHZu0dHNKfAflt4qPPLhrMJ7
jqHHXn/ugHr+1p9OqDTRvnKloCGpJsb6RiyWpEZ120ECqKWjwAK5b32BJ6wwCV/s8AiJUk8T7Kp1
rOdhePRAyl5mXNMQeZ18xdpXAWS3Wd4a3nWvsFwEVWg+NpSdjhAPElQUTEii2STteViFM/DSfb0T
3KMZ0s1hAjiWhFFdyD+sZYGWPGCddisuG7PEgvO6MfXIb7HkJUjorwQZyRAn1Tskec+nfyHlujFK
/9PAkcZ53FJolrCE4C6b7lyE4RU0mJxYxI4DQHsGV6g7ivmsN82FgSxh52w0EuU+osS2Y15R3iCQ
mqYATKm3UoiuFb4Xmb6VI1NvrvHZe07KdvLMmsSeX/YdDMJI/CM9z3Y8gmvP4JqjAhJjx4Kyh0K/
S+miW724ebA0GbqL1zoGWY3FpOD/6/J0/ZC/nZMXYojg0rpK/uCHM522TAlMeHj6nq/leUca9exM
Ofx5PRtEVbxVBDBKy/PFbZlVrDtB4jGMeWZNIz1O6++7Y62VXg98UNJ4se3zaVDqiNnwHc9rf+a0
NhP8AoTF9bxZFsqhx/B07T1nv6FUGMrrXHq8eVxm58zgJzLLMT4PR9CQ10X+Ps0Z3oT/hgGywCoj
s0GyltY27nxaUt9VgkMCnUbn1U/cvM2XtFIyLn/o3f28e8SwA0ZI7Z1oisLZFz+6biISoo1X20NY
aMcaXRCZv51C7D30YaQ+Oujcbjp6RUqGAfmsidqhIhsk4BfXm1tVe4x4O+NkxUvruBm+Rg2ck4bE
SRUYRD8oOS9rrPObdh2dyqu5dnHMUYVzsTDUWZtMBDQHQW9ibhvwJ0v+QQXAw8MXnz1b/23+Aevh
4paBEJ0M+dJExm8YwUJhe9Q0DiZgycQRGLzf9deEXrP+fQ33/12dsOxAPMtuWAwwLWvkwblszF2v
Q5FtZAv7ChlvfkQKYjtX0TpJwBu/vVlEi58KB/at8dG1LsXt/S7Q6rz8/TSstK/W4whp72njUB/f
q5r/lsflplIIL/yfCqDzzxeIuCDv9mgUiWnXETKYWzTyOR+ENZCX113XcE3OITNDQStQCgJFl967
GiUSi1eyGQj8dwCt7Zbl6HpG4bqje4Hdyc8FwxOSgDecAUB24twRZ33wdwfg/fL6mK3MOV/HIKDW
4X9MY12eQarssKUy4Uw4q3WFnpNCKNhw8F8nOm5SQHdT3A0z4dLnjv7dQ8YpNDbl8k9QUwxOQOj5
H8T/YMzY7VcEmk7os+rkYkxAkrm3+GTO2Ll8jjvzI2k5iKD+777GSDuftoDYb6haKcsS/lZHOIqb
68phpiuixeHEik7y3zc5sT9dpEv64cwgTDZ68fXXrjw3GdSxf+dqQ7rh0H3GN20F+gEC/uRpiF0o
m+eGG/ZBOpDt7zLCJrta/dRXQTZkS9l92EuoA5dPJshWTRYv+sHL/TN67Kr+j5+asSivw1eNovL+
F1v+f5/UZK/RQkX6EYHbfIBDkZ/ahhN/e69KD2WD2GXMlSlZAZIoy8xlGsKEvLyXcCykmykCo3CG
ekU0i6DWeOQqgFVYt//y2lhEuyu0ZYRPo6nLIbA0ZHMDVHR5yzQ7kmkCIm0s7o4+l1sjXg03IvD3
9PCiIKkvXRvBM0TpjuQ8HbTn1fPugyLOP9HE2OTz43I8sM3NLxJ+ZIUKRfVtQzp+lxJu5sSamj0V
1MeKmgPMH/RUun6LM6SVD2oSP2xu4DMefRJV739GOfpIClNcUsMMGkEP8n/FaIlUq2r1b7K5CH5O
Vq14S/W4KUfV8o85g4b947pHr6tEZfbtA8A3Ty6iSU8y2MmhphtKftW8S/Va9+b3tRX3X79AuISX
UgUt6fhhaIxH67JcHs0GV+Qo6TEg3VXTZE8o8XhXdomXctBQCwwvADqQqcr8RcelVBvJjtc7DzfD
zyuEXV6qsbaE0JibSFDB9ZfOeJ//7dv66bRg8DqFv/PgIpgsO8+YU0QJRsFI7275242y3hziJNKY
lz5EOO6n4KRMNk/zNJSHB5jVT7I5jJqCjiC88VXIcwc/hevKmz4IkLZgJzZXkmbI/cIWMT+07OgT
gAii1Bw2RO2EzDrk0Rv/W0qdLNh1sOOQYBL+rzzfPZOBVQyRDuT6TfcrXVCiqIMfGA0DHUQ2+SIJ
MzthSWexQXR/XMHlLI2pyluBjU8sr245vPwyEN3n4BmV44Etkph4lp5o5AVBS9plOCXIPyT9/DyU
5b3+Z8q3DM3U0WR/sTq2AbvubkQhyLpBJiB70EjrHYPZ77FDi0BoMJBpcWaBIniF+OJISnerUqFX
UfQs3KiUaTx5oj1VJAXdjYmR27CWvWEHyRjZj5xPXlisOxTv9x2d7l/RFkHpeW53xMkQOui5g8dF
tmWE2F61ijkxzP9LMSIrMocG3hOUHL5oY3p4ZxP8Z0XGPLc9LUhyIj41tGj+PDRlkRq3qxZxXfUx
L4XlIllvUNtcveTLK5HBOQ6mhMVI1MJW8sLLo1ZwzNCWEhtiuE2PyZqW0OSl2qVBb/s7M1nWCVNN
tu+UqDLt9194DS3LzZSrMdKvHAUq+HdKiNHOuEnICJzRseduemfy2+nQqqMZo9OjGNOJLcLNUaKy
DaQf8pFJqYSmzMvB5HHInWOv0oF92liMiZ+O0FPgLcacyXZwUA9XbskltwyvLKVaM1cEigDG3rae
CR4bBr8iovQZ/aI07notRARyaZXgu+nw3QAYhhNSZeE6cHMB5fVBvpmBevjPKkcDyjShZFv/IqBs
CgVdV1oBTkmBQ4aHtXfUWVZ4jvOUBioa1H1swZkT5Fs9cg+BQabfcegMCe8Pxyf1P4zUmIhEh5aE
ObsWjXjf7WSTfTtbAgnAA4hkuqH9bEE8BkDGcHsQdFKZpPF/cs/d1rmdlGgTU4Cs4XCWun0x6dM4
PiPnXwX3vtc7KNbgoWgfiWi0dJhwZxsJl7BA8WIgtF8NGJHQ+dc1oMr+pckSfa1aOtxfcGbMJo/F
QK2ndFu9GEvkyXzDxm7HkC9rg9Kf/PhOMS+leGGaM37SPwFzrzETU0AqL7IriRO7bJwwv22ZaEN+
+MTcAdpUIKReDmwPinSipm0kCPlRmLN5OsB+9Rqd0aMS+ziE/A8SslXLFKWXwiqxwsONNhWmVy4T
YgLSyQ40aFFpzpVDvkF0YcyJcHkxYiaTSGQlFpLPaTB67wSfun1uOVh/bS5iGJJBlZuHzWZGTh0A
V26OlxfX6lJAwftNMNI83LokeAKNNYxbWux6ksB148J4TmiuwnaIW2kWFC8S1Hf2nqdOb7OeNdTk
rboVugwMz/UU1PzZZBr49xeqSKYm16FGjJIKYmA+dYQhWxTB0vVHJ0dMNJhkPopC6gnWXl9PpY2/
Ta+bmZM0x5W0peAjfALuWfGvmOyC5tEMwPR37QFlLyjB4lgMS35MH/fh47jR5F7UTPjZUWWeID4t
Y0VEsWjjJQaN886R0FtPj1R4pyFFEFX9IvFKLsQDTMmjZqklU2b2ktA5ckHsIPDBNzgf16N8xmql
VQjGyLhNZWD9pD963Mu64oKbUnBPYJrhRiC6i2O3g8gt3KNDRsQvV6ur7OGbh9UpRKFueHS+xug1
3udSSZGSz+/s2kxoX54lcFbBO8xrL4NgEqje4iFZ2wLeZiPi0h29dNaAFRfY2JvM02nwuLSHTYUV
42JgHNh8/Qy+s1T82kO7fsCWrbb6f1xZuh37nruvK0qo+W+5oYY1BI8VL4rXe9IxyKIt45x6oCla
IYkj94Hv2N9FjHqiMiOBMq6M0LciTSVbld1NSypySh6EXH1V1hctvzsI8t42WkdBHGR0qkMubR90
+GX8hcA/wFcVlZE5A4o4HdQ/SgPo+Nn+5T19My68nwz99C3GJKtWK8M1qe+l/7yHghTnlqyR7kA3
zC99GC49NsTBfTxYBQblIYrTZGUiXMbm0jeouuwLOqVBC0kIJj1mHS0hIODcAqFZHYNUxBCOlaR8
Eh+texGYtlNjwEp0U8CwOtvuxUicAf7R6DjtZV6CkGrTlX1oziR4XEqf75HziQ7jCBxB/9OZWqx5
EuSzgcQ9aYauWYVDarxbHD3eKWzYVF/PuIc5Jgk3BRrjHN3Wr2VsPyb5PqjYbLPl/lZV7ZdA/PmA
A3Hl31jFxb1qobo2Li+tZjP5G3e+4zNk3LmeMEZNn2Wof+qgW7RlI0664OqW1mjXP1Ah/jdSgHnn
f2x8Dwfb3IqZ7LrH5/DdMbhrAU48XDD/IROjsva9b/2DnMNLSlRRQZ/qX1mPTI2hY7+f4U8RTNsg
z+jySFKfEOQksAAXecvxXDoVV4i1ckbni6EE4cpXGaERJHZ2/K8+GPLvjV6L7aAN/Ekyt8TMevOW
3S7JnLjoxgL3/8vIrhcJ0ZntfJ/AlMWOklDIp3j01pkYdP+MfTl09oz+rXggqJb8bWdgmcSgTZc9
4sTgC2rRn6qe4phwUzYDV2FgSWGCMUWhAYjvL4BRhefK8Rwb0uaDljc9DVrFmbxI7ceHJfD5E8SE
ZkINeFwwda35nf3VlxYqm4skGoT3oGrh71CtE6CoZuIFK9SXIT68gUThvxh+0FSIFPjvx8ZCT/LG
CH0FpN46MPPKRkTrGNA1uyl7q3MJqDwThbAMDK1kL4XID1IgGBOCWjj2y+Ko/FLTOPYKAb982NoW
r6k1h1OplqkmaDXsoLTHCQjhKS2hJ3PAUKif18gZdV5UpcBA1hPRTpvGKYe6V4hwhvgyjAL32Lae
pcB+QGZhkXO7qjx7jF61fTLsQs1SNNUTOUvgvFdS62z7Ui7EEop0tKgRn0F1xwMu3+xGHMxo2Y2Z
lHMOSF9aq0ifbeS2dpb4uLDOx7N+EsnBZmY3X4bvtCzeaLAI/bAPiMVsodlxIOm45JHP+08vd2z8
O1whL3meKQvQ+4LWfTVVmwm5SMS0t3/4Lql2WJFyG3o3aUK6GOiyI7o/2+XFYxwDYL/e2ZaaXoZ9
21kJYbTtwM0dXQ3T2yfVFAsnv0GyBmfOAkmbSFzgZKW0yM4r5L3y2c8vhyNAeQ0m9bkLz+duQjdK
mn9m+nihKFd+0dU5SCfq+6oiKcRDWgTGJ5pUW0FWDk2SJXN4dP/15gqKHHN+Dyyi/G6+XG8Pcoe9
+OCper+tYasLBYQEn2hLeavQMnd8z9bo4RcKG12CF/X5AViC0JT42h0q0uqmuzb2kcbunEsBi3aA
Y+KUfTy6Evae/mZQW4arMkKrUJeKBygOMai0+RxJtkXlLUYGWlon7MJoAhnvrjdr03iGiCviYnK8
asyr9B7UIRPHhf0vQQkpeFIbcuq+MPbChgA3XXp/fsBkzyCI3Z6lghDCCKKu2iUagJtOKsf+fbJu
5Yts6lPkznkvBjAX2r6tZra538t+XiDcwSuEQxsm9CEpaZemw9aq8zjcaAHrAACl72ys449SGuXS
dcsY2qWCHNoS6A5RMG1b2vMbd3W7na91KNvNZ5ozfFACvUAPtT2zSgJaN2MUg5mzycrxQJHI26Lf
5xaTpBnqp3X6PSOm6HvYVkABOPQrYU8SmWR5lyyUm6pC1DbwRHxaXadOt+QGr+jOJCieth+m9dng
B7m04E9YY3kFmGesR/S9Ea4LbAw8/RW/QhCX8NJVzXKGt8avxWtfaaP8brxkg8fsDA4atzY7pgA+
rYplWFb0XN+GMdKyaU8QulTztuozlJ6J/9Q21xAdo6CNeb3oxILIHbpM/rpqSQy3v1AdPCYlcCb3
TBKLUSpjumypcRJPXcJPtj0eG0v85+WWlExBplols8CvOkFOmy3bWCI2Dkh1iax1jWCsZZC3/PWk
yijF5QqetK5R4FXkpSxkDWTlaqBY3xxGxYUxGidh5UUqlOTKmhRW9jTPKlxZuvWxfXdbe7I0kC4W
hIKPW0zdu7DQnRFJOvprlduF2Gjn/378KpINOt9/hyaTj0oTxhEtxqmqnOy5ZbR8Qdhw5ixbDJT1
fC28vLlBCL7OIhbfsedg9tV0ONShTDPeztuoCamwKAgDMdqfjKzgRVTghb1uZCmTFQxkMQGvFFad
QXHS6wtvgfSlng2ZH8WlrgoO3xs8G3S4ED6Vh5gukhrR/VYvu9ZunTDUpvwa+gFMABftM9jYF7Rn
7xvXaVq24VC5BN+EFZhMwYGq7/sPe3KVfYCcydbfPLKjt0205IjsOnpSMG9a0A3v44M/JfmWenkG
Uo+Kt3q8WxoUcluhs6pP32fd96Z3bASpPaoxZKqx2P2fu0Rx66qE3OvjyNlAlMtFL+2SM4+7iAor
wkrcEM0cfMwmWFrabdWrTYEnupnOal0BnF4eLTHk2MM8n+xld4EzBQiL4XEODLkbIPGQk3TRw2uO
kYkjdRmPoVs2qCdyxl/t5pzd21dqKollzVYQUWLMAq7pREK0vWY+gmoXT3twOu5e3tvjZvgVLo0w
gRMr3kaI9hXef2no5eSQHD3jUd3OR8zUg4qy80IOscNtHZhjFt4G0N9vz0IEcOfnAJRGVS4zofec
1YAFOmwgPbWB3YAdvyN/zcBD0td8ydQD9y+ppqrg4gWVBXe6EgRX03USKp/RqucFhY7ulXArFEXQ
HTr5O2UYULNJJ+hboknFAuyI9hnUr/UNF+zyYZ1psng3C5z3HvaDsgnYET/U3Zv9bQpDG0ad8UDV
2nP1r72S3CzE8k+tyJVenrT+SqOE88Xg1gORdNpLGfxlLyq4qP+cr0tHLM6ocL8MSnMm7qY4dxNx
9k4YWO/OUL05kCz1VjgIaAJtMfh1MKVVaVMEh233AvbGFHE5TCsxFT+O8ao1UxJAjun6M+muZXua
TOPFWYdStd751m/AyG8XQy4HJy6Zun2CW+nwPlfHIGkULwfAPxSjekn6GtS3PSO68lwKFvXOTQpt
qKtU+GyW3IvJrReccbxBu9W3TwX6JkCACZQW09jb018ehcGW333y5p/eH56OlaaaZLbeABsoZSZG
yWYdafQ6t7XKuq3dohobLbvN9jametXq6AzsgfQU0Jc3IsxAtRVyJIlr9TGGhAvLubYzBHV+72S4
sGghVrCYadMihAWllUaCEljqMTFkgMhNcYVavEtauNk1q7qmgFO10mKlIsjEeCk0M111krUUgui4
PvmPFXJuNZz+Emz3wE6M+CiwnroFp3KeAtS6bGFmQKFPhHCQmOuCf+VIneGaLlRL5KMFYQ0Zr0ZN
r90GKY7UD/rlLnV9R8fuzQp/bNxKiVQhH8GjA7qt355dAOx9epDKN5g9kA9Ja0KmnMPWinGC+fIG
/nJ6MjX3DHi0YJQOxV/Gmq5BPuX28goaXiUvJoZcED5sBRR66PVCmhRGmP6fF63tMd34k08/VbS7
RHV0nMGTgTrCQCU15I3tlAnxpO5Ov1cRZM1CUQGaSKvlN73a2RdOvMBlTuoLFdrIjYhAyV+tbYU7
7Y4qOiChlOUEn2YI3k4keL5S4a9U7tAQCUMNYq5obprIRFGs8ERQNryMnhsknvivQ5CsgMlscsfL
JmmAGHJecdldAlvKywOOndwRo5TfGZ9pBrGEvj3R2jFcVktHzVc0R3eUNk4TIOgYZtTafF37cjkH
H8tWc8+byngIzLTuw7soOJMuXJmqo4ikFDTAn6d3s8x+bD8XvyqqsEMPIaTvaX2lPndnHP5jgG2b
BY65W8lk3TAl7Pt4Y3FTSjM/NPlyyMJGmc1fBdAmn3lsCJ4/RuBmAwR7vOQejF5BNSNyBtsMGD9N
JbUczsDiLsZcoHH+MRiEia3PrACPTZUSnbLCt69/dmPLynsEo0X1OnlBWvif89cqDUBI2VyflQrL
YHF6ldyYzghr0ji21LsE+Cf4DLhlvHNS3uVGT6VfvVXQnHCdxSTV1X59mrWKxuy/szULQumYnOkq
7wXPIpbXv+LRFyo+OarcXyg5/SR52W0FsEylu7yKm0gLyw0XFYjnfr1uaHrugu14Vf4YsJ2JAmxg
TN+Cs45WsmCUkPtK/AXqVd4WpokagUYfirL9kASwUukBNnbwRpGyIQdcJv5nYKc2rUSvCNZyS+/u
qxd2MoXtV0VxYhGn7GKHJoJ1bUkP2A6bRgxs+10mFhXWgok7wVtLhPG5JZOW3arOrLRGF2yM30eR
h6EDtx1njn7BJKnmrltUYxDN9Su34YAxu+15UStmUfVdRpxplcqz5r2lsBGu0Yi+g/vot09Sh8NI
tLfdpOTIgL9qx7V0DqBempxnBTuRLfqa5Yx6u0gUPRUKxrLZo20Kw+lN+WkTvEDjojU/LliEI2UQ
9RDvVkS4yyOjlAw3YSSjNyy2TUjJ41ByzhSEnQ9TuTclohTXqsU0EoXCbsTCxkWxlt2rB+zLL5df
NrSmV03AZGSKkO1JATPP9PrVRkYw/JmpBEfWv0momuwvY/La3iKx84ThMFq/9RF+vLYxOHA+81Lg
UFd4CgwiSMpp3z8ae1mAISGBJ2ENd3LbcMzm4/dB4zeXD/cG5iUCOuBq9nYo8lKLy3J7p4qcmy60
uCVrOUMTA8FbHwGRdnyy68R2SLtzHI80AXqpjC3ZuBcRkMrFsqmKeUg04nGWypI0RWIZ+bBqxDj7
NEeUQKD+Q3DtZDH3K4aCaNov/h2HZngPvOvkfH02a/qq8XMxRZwCS6S5dUOsHmioQNaNZBlfRD5y
3xCk6QBHBZ7sCMz0zoazrTjfdicBzCPAKPbjS3dHJx6Vi0uHuezDezDbHb/vC9QAj4HdanA3RdtY
hhT+OBKwLIikKsRUtxQB5fHct5WxEAPmogt2fTZsOHAxZlBhVNTKGLBFkHm1zkixnxHhTqd9mSZK
hUtNWJJfGLSDNge0Yg5coqp+lBzoxvjjwyJwiHq729f/wDbB6gwtOUmzAa6i3YEXFejgpa+B5epE
qiw0uhs84Pa7JxCc1C/KxUEHrDC6wNm2C9hqcC4nmNEWPyOMm3guzUOmfKS2oRRg8H3k32ahNIhQ
WXgPsseFLUIwl9MPHkaO2qUy64ZeZ+E2i2061c15kFLEm5PbnbLeByPNwfOrwNZatze92hjNvTVR
mwd0aVBVbKjU9juMIkkwJbZ3htkSf+djxxy5Qm5nz5nSRKvocUho/Cp/eqV3Rhqcw9XQsiGq+lHL
UBg8TZZwcrfxcMcIA+4DKx8IQjaMOW8RWNUAgd47XIZUMYC6MmZW1B4a5om6wy3uCoflJ3jASHeq
vMSUxvGH6ixV2YtAy+SgX/ZxtypWJCg8IhPTge08IVo6j2BtBbQbRQefhwhZAwvTCcn+tB89PLcR
b1xi15KuZ/8omU8nWn3hHChpC0BO8yjMUZX4qhFyFaqYw30jfSrRy7uhHDft7CP6rCIUpliecr2o
df5qXJz1lrEd5eFNlZEeWtMSRm+vKk8o3EQWkm0OPIeoVLGH7ZhO65L9gltxVSHCgcNGxzQcJE/r
MsUZxj3D2/bq2fcO20PZ+0zbKpllRL4xEydRFnEuffFwI/V6YB3LSEKTkwVUVgk6jHH4R4vDi4kX
74/xrGrr3xeBg1aLZqSzCRPfmDetyCX5NDUPa4Yfo+AC1L1VOnMBtzbJLW93k19tKF3iFH3mhR+q
d1o7K8RbYyEkgz7o7tSRtf4i9oGRk4/N43A2ApkBqbj45r0nnqTxsFjIbOuL1O0qOzxE9qMcYvmt
CTx6GTDKWaICczRzQeLYZ5p6fVAJL8is8qhn9ylXe/Io8udh9kk7g23KEDw8q1YGtf17nliEA+/+
OdLmFob2iwCH+WSVauvYx27RL9Jo2YdpYrdwHPW8cTtlnd8a6bRQ1ZDRAxi/RzjgfIyV1yLXTy3W
5dGijoSa94ehEUsuHbOXV+szWqu36SYUMk/8I+VNhSrtF0xKqHjy831y62FsgrWxye8R4LL/qWwQ
1qE9LlQ5YcxSOm7MSeD8dqjQ149ijS7o+stXpJ9LBbU0Rk9419pBQCImiZOmeHMBktxdsAQIgTzb
+lRxtFcWvXle6ib621Scf2GR6SKkiJoN5OuUCiadgIRvLf6yJ7sy1up5gLToLPZ19hHEia9OUVEG
b5x/W6q/iqADcPCrNCMYn3qXHDFGAXS0JOtLTUfZkHxeLqVotgHMCdWUas7bcPq/j68UPbRyZ4+C
ZSxCB3zWKp6nsZrugiBX4y2iIlY9wTk0aj/2vtaTbnyeaH8pRRPz9vK9Ph0x+qS0CooXeDm6mUZI
jdAFj9Ia7rhw8gBnz+ZBBtES/RTOqRmwuVIgPD7OpPhRXlqkmSVwHeXbVk/vDWzrrWT2kyRbtfy1
s+jIoTLkaQepcDYWc5Wtzh+gSAq8/ydIL9Ait2kFskYKwi8Vl2Q8Ai5mxhWwRut9vxL0IeV02gWL
PBi6YqDuNSyrajrk7rq2bAYfjHjM+7GLhVi0rqsfAf4rAIUvzWpyz4FCs8bJRRcXnDfdUa4G2d0O
SnqJme6JXKDNzWJPEsHrkAWFDX6/K26WLApJkqVs4wbpMDr685bz+oMGwyg3jfwoFkyfDRnyt+0R
pEgsbYme9l9AOKjupk6dAW+TnL6kCXKgRxZIwJ8tCPyD720o2Shq7AzZLWCsNXLxkiY2GwXrCGzg
wj1Omts7+LJVbvQUZAV5F72sWvg/TS95fzNQ676sD6aZ8MMbBBEBBbMtDN65vz+0c3/9LAy33/Wl
nh0IQHbqDfuffWsVOzCsZ0gBGCFiF4F7CTw6bb1ZYF/BTXSOdK0a2mEw6s301tiYYgmIoooK/LDZ
HvJ4YwxNV2wEhUDjYsBeZl+v8sLAV7cPQEXU2rbibDfqevtpmiYaAg13K8pHR59hx/1Ep/nSeT34
eW565mrXQFYiONcGYE6/d/V4PiiqL05CMf7fw449MrJd9LHp7H3xfCHjZfTciZRoTlWUnOo0jHhP
Loej7kuuTiViA1+hnl8vL54vBJ2ntU2aWnfRLa/4UhcZ9dtOx79HEDiQd13SCYURkzMRUjh2DOGj
b6XRK+ITwvd1zuVKnVN4XrFZDqLYRMjZHR/9IRsy9ewnTE4cFZ6uaON/nmp67M9RNTHvi9Hn14li
g5kVQLo398sBI+MaieO1TA+Cg2rD8cbGqr6qrTiIdJVc9/pgyf6DB0hTSASPS4j9Tb/9yvVoZv2y
rG1i8VPKiFr35Sf1wRCRh5vuN+M2GeM+v38jYD/CeIzEEcCI+iejIkFvY37rmezed4k2a9eUjf/l
5gUqgbt3A+fQ9hq0Hth29nlJ+G16jlbLHSh6/Zn3p5LEI8s7+ro3jMNQvc/BRAwEVvXdBEvkrzVx
sfCWE/vFjnwR/8ME+Su0f+tVUCzqEoSzERdFxXDH6oVOBppg/+4BoDbf8giwqObHTmzIzJY4hJUS
bLiicxpIg+in2yrTTBoTcf9xdv4tDwg4bf8kjbtEDoD4d8aNK0eQsOR8NQcqzhky23V70Af3BFzs
uWRDGX4c2SSpPZNEXRjFDZLrEWQBbdCSLMABcBz1cOTGfj2HhWHvhrGzyusPn0Fb7BuFQMtu3nWU
YsI5jBkw3CDrr7azlIjDj0kKWvvVjUFgL7eZtthFR01hSOfTVQ79thCS6m7zLFw0Vz3muS6r/mgc
HiRN643hWVxcWaq6dOupjgOPiZxFT91bnMINStypgYrf7Wg/2pm7U6TcVoINQoSucyHuFZzAjd6J
hrctiw0WOb/kZXI3r84rB6Lhk38NyJhwAbJhfOpd7Spjx+/LBB3j+DHZv+4bwS+Lwrg8rutMwUoC
gLt6H0AI/Bl5q216Za7aVdT/4bf/KpCWoAHtAIDept3vhHIRZ3yJyzBHM8+VvQey3W9Qbeu4PBb9
JraIzG10CtVs4romBBBvkrdwAJMRgTvv4YEVhM3mbrp+067u0lxx3OfJy9DUsefIZHwPj/xqK22x
G2t5IwuomSwNsKLLya+ETvVULm1LJqrGWE3beDdIvWwPUCzg0OnByj+4uysMYIvdYLvL7zpqfI9K
t3rmNZZ2IMv/508GId4nrJ1cX6VUFKnu+2PhyehN3jrQ1whIDPTz8gTsTc6tJpQ1ksKKEuqH1qBN
sEI3OTRyXwGJSMLldMW01t63x/uTRlhhn2gwHRr/rU6MYl9NO2VHRUl399xah52kMZLYQPZTzs7g
S1M2291OytYBAOPcvX2I0Gloy2ewbu6ouKD9HcfdQGd7ZFEiO4Lex7UMbBAAtLzToYTUUdIbAP3p
HdHuPkDJklaYY03EuV1RJL7yczTAZyaqPMMo8r/fF/QMhiKiopNNh1LMsgReD3amOv7L7RvfOXos
WvUw3O5Nvj2DYVgfmK4WPz49J1hQhGlmW2TRx6mWXC9tUH41vUlBn0NSl/xXbjSh6fdpAJdOkN3U
VTVg7sASF+I+3sOnA3RSGON6QqwVBMYlWdVwtM1isKGkINXns6Bud2RfdVk4CQYmV06PrZu0m11x
Z9/Liqp+2hDFOIihl+7oFN/2TW5FXwRVrVKIx1LcUfCFDSGXChdp+kWjFxuNP42WLyPoZXmXtkYU
WwhpW8mhCisy7LHdAtbe9Vc7XAxEXxkaaYC0dD1OzzkSoz03ZB0kei10V6G6faR4MmFmaoJ6meRs
wadth1+19jgIcD3bYjpoTRAMMOoFzbzyS9+uzWqFL69N+x5SkQatwXeGBGtg0gj7CeaToYlmT8R/
1yOKQ1nT6PkoNpCtUEd321iPv1JP1UC5cFRrlgI5oWbqns1ZW0J5T77v/wqcj5BbbY1gbDAWmNKU
2Y3OLnA1Iro/icEkn4i8zQngAFBLJ6en7u64rUZe97NbDgMLJhW5r0AB4wX80lAWosMSHLum+PWM
Kz2lOIPIRFv3Zt5485ZAuDkmMaBpdS+TbdKExabxkfepJe6AS+jkjChZiYZtyCmumwnSGjalwnKO
+DheJEeKHAVwNU1gpiseSnR9dGDCO4Gju1z/Hopw5AWududdD4AzGTaWU2z3kMK8kpzt2yzZZ1un
MzYDiSb7WRxcxWK0t7T56XvMPzM+tBQNe4P8uZ1aSP/dHQhMzgsBmjUHDojY1Y8XLIBcnjGo+thP
E1vri2BpVQA5yHOGWOAqhAM6S/ambOn9gXqOmQBcMWSJyRE24WzZKXyaQ0egpuwVBlrdpNan/ABA
ZINsenenAE3qkauldm4bBVFrYnsP4J9X/PDGb2pTBMoXpb9JXd3LmxNPU57Rgj/+atI/EuV2UBC1
0ee6eRXkscI4wFztk7LWkGGXxFqSpe4vsiRpbvvQOQxXhjiKXUl2ib+SsbHTrSlP0gEy1Y0eIEvl
tQ5N2Fk6OCYfCzZFTp2qQfgZ2DFsIw0PaIjWObsw6GsRckGa3MMuZG5IHHNcyNbAt+xGnXe36lkV
okMmuZzyuutwLm39KghKdJZSD24dHW3RnB8pyvWdUVtdNJmXFQDqtWmR8f2ee11Qe5wlYQi889pI
Fajot8+wFEbM7eb28BkmFyo4wywFizq++Fz7I9h+obZvE49roDmbFDLEDa3Eg4XsYjJO3zr/muzp
nbmHsV7Vk+h7gaK6br4GUZmqQ2qZrzNZvqhyfHmoVC134KHiudymNCUvIrrDRt+BdZYgXxglzucp
mTayIriwxuA8qVwKKlNFKOD5ux7gve3DOD374HJDT8BogijIdy6KGmkfmKGznpbB8ohCH2/KyQ52
C/bWy1Zg7I4/aLeC1KDIG7JegNy5c2p1ZNQ5qgqlIozjJC0Kjb5DYz6vp57QnIHZyEZ/aT9IXdsV
DHUbHW5nwoa+L//BcmW0FkXlohfZJY+TywKyYaNfJeCDsK/L8b2cbPhKIvdom43ZMo7eyjt7NsbV
VvXymd2LK6LoOF9oZ/ZcJEJRoB8rJadWYWKMYvdAopgJHHhua7Iy83WbLu1n57zsUaT7EXHU64Oz
eONO414MlHm5WN3Kc0x5kGf5MJXJo+b5q0iCYN8FvazeyQvirz6NkiWsmFwzCF5EFBZVOJ08uwDE
tqpYwH9gvvua8ZBonVo+VcSOwPZpuyGn1G+P8ZMZ29aytiZZ4JzNfTeQg5NbSbVeQVe5i7KSqw5F
AqlOKy67Tl7xUAD0p5FHSppuRSChaM5KhSzwXi5VtWcEtz1eBv+5ZmVA6e/F+kt0cJ1p0YEbIJxp
hSagq1A4FIu1FgzjhPiKS03Bv3owpERK+ktMAQW1trqlKtt+mJLOvjBS1gRtC+jORu7KI1Fu+oQl
liCfX+jdsGwAdaIX9GXcrGulftkyRxqr4gfYcbyEBI4hFuYgGukW1vcsEeqbaEkEMuraGDixYgfO
GpNL8xr0hbd53PEhxH6VoEGaz80tbNivkT0jacoteIJXkyN/rIEm7BtHWij7K6Bjml+aygOpePlB
hakTroaXoOqHHg65ppAwV86O9WBmQcBXC//6WI99uH5GnWLNxVfHB7SLAgedAjkbAQiyv8H17JmG
dZYJIu5UzjImieFEMKW9OYWLZ0zvAmq8SciDT675I/D50kA7224L+Yg1vUhMuMnwazMYkUbseFyO
/isxBLAD2CX9vukSmAJG+c8VEz0CKS2KWh/WvXBzjeUl1ZIwy1eRpkTnsKXabrszYRgWs8Iganpl
u4Acv1WRglLjafmwkhCAs9Zl5LSboN+rx/dmqlw5ctq/tUZQmnEvR1VozkHf8slglgxeiXDvvLVP
gVrrXqSONotDB+4nKE42HDLP36nNXA9VRoooXc7LkOetRgJ2TxjspBqQ32oQxzwkvDbDnB9yOW7x
549LxzorP/S9RhpZLXIZ2CEeLooARU0pjZmQlqbhf3FRRvpX/Ibe4ISj2dDdipUdkzK+S+YMsilc
x7ODG9CQKwjx86i1tQcdsvLuof65RxbFdRSYwD+3UPY/bows/mI6/0ITwIM+8MlfQRe6yI/0sQdG
HJoGeQHkRbB11ihQCSFedN9aq9yyi1QxuEWk5OW34uvpzHSiWV3JYjgleI8arKNB6SpbCHqoZuxg
j5AQToWxd/86+8woBEEyXbemCg+6ASiEo3ZfdCbQR94rmhxJcpsQcxP1KW7to253Y23USaehuhb8
Jz4bHau19s/0SXPaTeNO3u/70o2/NSszwVoVhsE0KkU9DA6vGI9siV8ZSKV9h6mvvCc9ZWN5wi53
yl2NWqz6A3svV7wGGXJSLRHj/jg5I5zjuhA5pqrowu6Pqk2yksrc17SpGGuXJp0gBBdNeXh36eRA
wsF227TeqFZlH9Lavu8tO3X/QdxIN+35wUp/0oCeB6/lE4bJxwtmNixV/lbTGYrBigqZD3v0wLMF
wR2u+VWeqXJejDRz0uPQsqclX7ymde7rd9zgkqsvlNcjssqJJtni/o+c/PwPjjhZbEMwZy6i3HKc
3j3DyCqBA6R26VlObrlmALhkCHbTrZmXxGzKL9v0JYGYLLn1eMeNEmgiPRx9dDlCz3imK99YBuTF
ByQw5U3s/JY9tAQ8GuUFJmX1gQ/pOD5+Lr0cXPGQybo6xVEPvI5rn8xiOqvCkjCWOPDQpycvpdny
MjuWTLsV6CECt6G8fIogJEcYm8cfZvkBG38ItDvj2v7kJAtsEWgbxzcml/LkRO6AjrtFJvIZ/M3i
lLSoP/jv+XNPdkgyftUfDIyUgYVewnbqsQFa570QyxV6grP9V5puJuSb6kJtV0VeLc85xeCrKQ1y
m0TcdvJNKYhAI8TOfXUyozRg5Wjva0SqrJkFKA9fVwyqNJTrVS+qOtrO80pydsWhIQlILs0g0Tkr
qCvbySeT9gbociKcTDNGzbWNU+EOrveZd2EXEEhJ2sJlEX0ldxdFISK+XsMqObE19d5jc6JCOLOb
yGi/IxcZmlzN8oDz1tYyVQjCRjtO+3y/efCAher2rz4xgLBY7vMxFdWQJxQEjkXcdOgweB1e5l3M
64N3Pg+QBi+N0nMiWa7RAjXVzo5vRcov9rRl5vq9WamonHxGPncbMQuBX5e5YwwX/Y8PBt/PVNRZ
quHyK4PGz7dyrO3NoZHnNj652LvVwlsCuIAsxQB5pJb2ipe0L7OotsdYGoTe6ao99KlqnWrw/byT
P8dJy6m1DUJzQ3J5wAy2FQo0NE6AIVI7DeZ6awdq8cBbCRSAfiSJZd2zJMuPCT2qZIZ/f7xngCUk
d0Wc9vBHWjztJTT+EfYlQdwNk2L4uTmrnvd0qciahsTBHaNjAeD8HEOCkh7nSr3ASDxJYqx24COZ
oMHBMvGO+uSEvSESLI+XJfzONk76QG4uO9JdvKdMTmNRraU77o5Ydy3d0MCxF3K6an0FF4BAJcHX
4gK9aee8DfqarAQCw4+F4XMSMR/EQyiLDUZpI7glVv8aeDVT/v+7ofaJFr2XOobjmhC8SMiiRkrh
ueJdbY5khrjM45XR8ZgymTs8DfMF+oa6PKz1gqroHCcqk0nQIwLbOYGzjVnDzIgA8O4GlJX0SQO4
CtHnjv72hOvnqB7UpafHEmDdLC10nzG7CqLTyt3yC/Y2xj0JRCVVmIz8cKLaXk1YEbV+ZC4tMyjW
WyXK+MDs78e6pZySHLtoPMc4DczVXcB0hEpDFMEkslJbQkTY8Lfq1OfIxW9+mNAjWpTDvtCZjyuW
noocl39dqSxe1JRZkByMQMERLWFgVCr7I4CqYxfXrgUYS3BcCKoOFuMvVsmsRDyiuDq2RamaEguq
M8n6T7Zodlpv27c/JjVnBTGg/zgvtyL2VJvyk/vWDI0e4J58G7fd+2SO6Cuozn3kGZFde/0XbejJ
CHNtmRWz8q7n4m10EssGF3Ar9IcWA07PTceqcs5ZkXIVFKQ1T8hXvXroTdGLQSI7KckWPf2yvINI
MmNyE3LrInU+yB8EgijTOwU9UgsNO5Nh0XR4wzs6vIZM4D2gsHLONUHnpe7yD5iK9ADiyaGqwl8A
Nfo8xDzdk+CBEFrdfF4kWCIHcxA0wrHNaEKvUqsqXjuXPaTVqL+bdxVzfzkV6sYwgTJRBEDXTE7l
4gT+3P5ff6J72i+2MFNF/mZF0/12Mqzh9EDTX3nw65bq03RYXKgl5Yj5CBOTJECL4yTzh5PQKOlx
2rOXRm6uQLBSTGFJVTaMtskLmtIESA9XVlsLJ3LAvmboPYWTwL/HNOCxmdPq+LnEWztmtIZ0RXxV
CHJShdt1TtyxxzAMuzhM4HehkKQSBBL2Zsiz7ytg7LoTWpFKY96MBAIT8AuzbInUIEdvFgFXV2K4
ug00ZyvX0b7v/d1fYs4O9sKKswZg7GHY3QGBxp1sxaf+hlno8jolZ/D9UDU7vfwI2I+j8C2ydeWQ
32Y5WgbZmow3BgtvF3JJxj2uxMO+5kCuaumiDXz5KMsH6tcikYsZQCieYR64uYN0K4wHnkwwe2Jn
X56MxNcQAch8Afdm5DBY1FEZGqhVH3GfMbonloo2khcT3IY4fd/EYdcNPcUWExd8wrUBWJCyFjUe
BkZLRpRepUIjpIVQaiReix6X8uwc4Fv8tjkqgE4kRgIs9DtDIBFLMsBCmXPJNS6au91t66YeRony
2qLOnglnTLqTNe0Yp5kC7eSO7Mjcop+5IjbnTbkRzdzdCu1Z+6LkzDaF++BipVeN/UxbZqjCPt1S
YPqhuqaYg3Dw290VhZcI7FoyqF8qz/R8HPml14LdWmXOWjL1PZt0RSV+sNFkLpruIeC96sornS49
oGWukVYLLzS3QvrOpmiwsOAel839ivjIZVtlMY6K/M6AhF7eKqLs/cozg92ByGBIQxm3xvps99RE
vTnpIbY43VmDRU7CsnqklC+r5GriT3WY4kEt+x4EEgSaKx2JhPC4FDi3l/4OFN0yaaLJJOM8tz6p
NsM6qDrqVFEP+10FJq8zs2f/QZs0eSy+kxIxCuxgSLHhAzP77qgn9T/JsLkiEhUkMtNo5PNvvWN7
cPSd/ZB1Mt6hwxIt3cyIeT6xdDl8RUh5VfBisSyJflCoZOs3cTUFA/0L/8ji/3qD0pPHLwrEKSEC
wd2zuOO314qFiiA3SM0bvh5VKvq7se5q12H1O3JFlj4Ja9codmzvlLBCjWtj2kzPYr2f5VwoPCrK
AG9XLpeVaTwkCxyvoFUDPDZ3+e9p00n4uBpbF7RMmKvQ60ml1KN04ldfc6QwIDvPIGJqL8k9E5lw
xRLBVSC+2YO9rLkdBxtAfCKQb5PFJzP2J0ySIE98S6DlX1MsBmM6r+OFTX/z2X/o/YrTt5hFJYbg
6hcV+87xnPhMbEUzwUmcPqnCJKsLcPyMfuZRLg+GoFhu5yHEs/sB6G/WtVTQ6yzmvBL0oJY44i6g
69YZv+/UdxQRJlITb2EKUkWS+Wa96tY8bYxmxrPR8DpM0yCTeiM9fbddMTyOS5StQ2dRbokMHF4U
J/OQygvHYTcPcfsSwdVVaDeenLGV1j0uM1ySEyBisA9WEocoRA3/ATZtp5/SzbHdD7U2/a5+rBSW
Is0kumTfvfoECE7+KtSghOyFYNFrpVTPAtuAKjbZSl/p393MfF+qVK0Vg4pPb7vLLRBDfmaI757R
RfQIVUeaGInkjKCnUWb+1rJnFDWVM8jbYmi26xQ6COg8R6PnovrkaMyJgEHiUNhNwxmvPbiG+GYn
5982uP4/lHxKNhJC6wy2B9Wg9PUvv6IidH7az22eXhCf8TT0uUL5J0/SISBFWkiSMyBe7SUaL08P
3at20RIORB8q9rrX81BWCTBb4jIfMQ1Mw1/Z5Nm8Q3n3kQf10bL9sIL23yOrCn8m1mT/mpFT0Jhs
Lq0Y9etEqAbZQUJXVEMYPYIxfdABc0QtbfhB0ETMKVc46MjV9EJeqKYSkpjUaBgYoBD98/qIIUll
KOUeIPwjt/D9yuVfvhX/1MRsjfg1xw1haNOJ7IZzjgUmbroXrE2/QUnOQz3UpNeleSZaJDlXLZzO
HpelwDftf/8CQXxtvh/BEIievKxd/y7OtE6ihbqUOi0fvw+zupLI6Pq55zz/aF7dytayLQN36DNO
JG0agm4oPtD7ILvCX48VygXWLkv+B1JWkPo0NV/+3o4Nr+aOCJjR7bJ9Gxg5QY26PxXWhSj40Ekm
NTOy69YiZIHFIdVezePziEx022wLbCQihUuN/KdOcbJYGGoiEDsJtnrkpGvf4UsW01WAZ07Vv3p0
/qxc1bF57386VHVA52Ae+Oed6C1KyYz9Xynny02B+VP3NXTBUTvOMVcmhSyTW2feDNSjcc7K45My
bOWARgEYR4+rwnHLkSNWNxtm9ia9dbteTZCp4dAy+sM6i0BgxnB6tVTa8MacctcacG9F41bHixqe
sbwA/WfxQYo3v5oFpGHSFNcCEdR49ss/EDF3Q/jBGtaL/wBN0O9zAN5GPSSFTACaVDCzlarV2B5l
R/n1o+KNjcliR44GzTgJysETROb617JcVyAM79gi2YnffpP9g/lT8ze2sarcbfnFHWcAjCMvBLNR
XhcaOT3hK4YfkEYREjPYl/cOOSMLwA4FCyUP3D34/8HpzcQzaHbGajTDnXfB2XjuLB2gtr2tua/8
aJbYIr32XGE8YcI+7GYwsKy5BzqG+xyh9PbQywHA2r1hgC2JUvUIPwtHjpF+IJrMr03Ns/Jc0CnO
rcoXejoBlwlzBnGi6rghBGpMU+GWV5/Y76cinrAwKG4ZpfaMuW/qbwzSWgjdjQNJ8To6Kl5FDB84
WytZqQKNzFcxdWSDwTHGEm70fS8Ne8qy77uFWizSKfhy7LBVqi9YRnkrJ3Y5pKzJtw1mIwBFh0vi
Ad/rrKLTBYqBxLVXtpv3D7YexLgQ3OEtQb/DwPIjFqONbtf8wtGdfg75Zq8LUj2RhyaH8BryFYmb
qkBU4p2cAwAtj4hjnUgQ5pIGE7K9cD+6h7wE4fFpbjClUdm4UsKGOSYr4zPZQHJDrPWfe0eAUYTm
X9WfpSVSQeZ+d7ncgHb4mrIEJ6mAjpN8IdkW5ZlJdrSYiAhZF904NOwzc7tWN1dqDzmPRztKYSLS
X9vEaUeFs6ktoaLjgJsQjWl5pz71hv2paN5W3VXhMbzT2A1PGBWCih7xo3GCs022HzgRrhBzrdrp
b4RRkZBvefQjXqYFbRxSU3TO79+lTfyEYabl3SUPZXE/44J4htqtJQgbZOkaLGsyYDp4lfXAYAl6
PeHobTdsywEM4xpie63rWrg3VuedE3hFB/rlWn3ptUWkKX4i5BJdbdvGcrFyw/Sc8zpDY6uHusVR
6YvHNQhqIW1eBlOoLruUSSzGv90nvm0Dj8n7A01Plmo9zVFV8gTQf4DcG/CIfGhm/wjHpdxS4jrs
AnKqmn9cFrVgL4bGFY+2buewKpprEQYYtMgT2XpBptfFX3NNWSYn04c6vYrf4lONZ1E4VcyklLpf
JsUvNh6GTQi7B31VVjMt998T/2BqTnCz6pV8mrWF2LmbdvpbahIbS5rXi9/t15SwAhd0tAwjHrsL
jQvrkQ9Bs/pJOTPj2nz1CguXsvs8/bXQkCusmgHJgrWHj2GIxydMyQSdcBnM1cbme+bzvyy549AZ
46IhuAiorpCWM5ikjXQeSlvq66eTtRxjoNXxd7fanhtsn0Z7VP7miS+5rBCP5bvxbAT/JTF3vJCG
awSoiIwyMfNyYn9ad1EsdReVcsYLf3ZG9ehza2Sbc+Qn+j7TQKpn74OO6sB8/sgYZgS+vWWaTdhq
4QNIraTZKgkUwr7qYWZsXK9kMcNO5Yr5EgLZED3+G7qxJbJsDzWg69ivvV85jFXbSJXcUsNVXxz0
7hLOS4mFGAba5/NonrTONF4B9fL7khKO30ssPEKZES1GqyWZ4dx8kOk6u+8BH5+0TTm+1lQ8mLLU
J8KwCWBhS+myReeEzoYjI//JCrrV9rK5mLNOVeKCHtjAr4GB7u/QaERv/72ecxUm/qk6naxeJrUD
rRjProzX5cWato+kyzvA3TaKTeQs3E8lpKWgrdGOOPsOVgaueyaF2Y7xurvEUj1NCvSbxvE6LtYR
yv0CkvDLWLyFpgQ3+W6bpNMp4IxnJjHSNENuz1SLz/NKp0ebuUx7sl2eXfAYEbk0WiLj6Zcf0HC5
9MbYYkBEuadIuBAOWWA+nkl60CyM945M1Zx0U29FvambCwlQoqBCmodsJThg6agBH5SMlWdk9GXV
klrYQmmyYpP17YW9y8HXd+2TfJluM/YyBVEEMNwKkgHu5vgfBfl1aXRMaW11f20So/wQIRamtcXB
iSCwZTeUrYjibFNuPuGcavaCk4UoVkwbMB7CDVkEvYz9x7PclXqupe/egvxYoL0Oz+xxsAJ9otB2
pH5GbsUWt34bCdl1TJS2R4oaIcWTmzKNCNLZYNLKqdDP3Y2J/bhrmTuYDOit1eL+1GPkyhFQ5Ikp
mJdhtqr5tGDn2SuGmiSJN9ySzW3CK/VLACZgTJScmwBcFKbdIQBEBh6Ed7aPMGmXnI0Iy7RIkQ/r
2FR7xvE8XnQ62Vi6nHtYH8fG1mWaO1EDW5p5wz/1yK1vKylzj5t+Zi27Z+FLl5lmR4S3Y5jyNZQm
rLjw5LS3yH2iMIgxlJBSSGFCAWBuFK4q3pipF2rVxIDvfN4MGAdygo6W5x8iz/I7zs7mc5xOQ94q
5NVd1F38vy00OHHFyftjsHhFjEHhr53oKVwcwJUBVQyzOPv7kmTOrex1MwtYc1aChBY934LcwtC8
SqgoGvpOAWC2coXBnY+UQNUI8Ee/zAVjHUxuR0/qoXGB11G0peBDehVvT7DJRuLSf3z+QpKTzvID
xGnwR5rLCRdpc0hry81Xv6gDaT11pdh2zDWBwPtalBxfAhZJJqxwuoB0HbGQ3hltpTIORzfIfrpN
7CsUpmweTEMcRcTzRLtnwLYjzssbPG4cS0l0WtdpK7i28pz2J2o4JH9W4jIKLxV8ZL15JrWwoieq
12Slqe1WPwl/2klQAaTsBBYX0eH6nrPzs2wps/3t3jv6eCPmCfS+UpdjYvGaHBfy+7HBI9GGwI5P
CoIDIaR48tQXL18nH5pGwVR5NUAhuO7Jj3vrEa9UTw921TRRXDSnmAScdfl9BKv1c8tZDzQUticu
icMoKO5ibH2Y5xRBETQCiTrs2xqJkQstwXFh8vbS0X4ceq2kXiiJtwHmjZvI407HELWV+JPXchTh
mHw2lo2PvhptnoWVNc4Nz/bjmwPZkuKk/HmjNIjFFmCmC2MdBZ7kJt60nvsXpYWehxW668qqRDk9
iLR0zkVmgn/SQHOSYQu2oE+zs9Nd8ZYMhZ+KpJhTA5wZ46ZGUrOELqNyeKEptlrZwhNYyuIMT6bQ
is+bRK1E5jCpuirur/8X4xU8O9yvtmeiOc5hQoO5NITyAiBAvCWmqH3CUfLjcpgCTLBRF/z7Lxi/
joxOYvJP6BXqE2mPxP20qJfN2PkaAaLtKre+26rschI+KSE0YWKX8UEaWqtTB5KlTSSWYg/z9LPi
gYzNdSGtxnkk4EQhCjwOw2sDDLF0UWytN7Ty8uf+mq6EsVYBRj4X/Gs3xSwQHAF/c0cRFGIKOMH/
Wb0X4bjRPya7JBBuGZARBMWcV8yZbgEfnKWp/yJZW8pFvAi0+7lgPtXVaBI4Pc95sxXqHVL9OmNQ
aCCH60/H+kI3LmktKWlYvaKSutJItGApO+TkKKmzbUy39X4szBXmoLjIHqSd4Z5JGaZ3goIDzvXq
R9ofzWC/WMUUbQ1uBhREJTZeW7JBQaZQc6RexGd+bvLrvbFFORyd4LynwXI0JWs++KOU0vRoye8A
golulnZpUFe7GDuBK4jiOnJ8Gq4oPVSx1I2DOL5XCtcyKSHCA4zSpTckVeW5lcelIlscFv6bW2I8
sF7+hKyEHD/OLd2zK/oIZ6q1vt7JY5G5WTSGEt6NM1VuLyT3HAkxJ1J9kx1AyBaIxrPR06j9ljvW
/9rctKkHSegr8Qwexu1lfvU01hJvaRnrUKFqWwcDQFEXfEbqmO08ippW1f3TP9OpghdY88vL5qfF
UZkcaWm9fZPTdBlVh6vSCZTdebr70SZ71swUSgjQ4F9gLYoujnzvUewDZ38NQ1ZM33UmSCP2PEtZ
CHIufzNuov+YC7DC6TL6+7KJxmlBHMHNlBaC5kBvR9ahbbhrt50o6ez+rwO1S4XCPsrZVTlYhj6g
RqxZghWulue3UwmGFK8JaL3WfdJ+tH8BBBL4fi8Qad9nMmsye5fnp6Yc8sHXN235SJ2PI3CNLtIg
z2FT4EgAUoHHyKcdyq+LVmxZbWppqBOsWXEAn557SHCK+ZGrK9iQqumXGOzrlDL8sjojCctXKibZ
GyDoNl+0j28PyF5Ze84dzDH7LCDNID4TgcbseKG3JrvGDW573SHF2Iu9S6uVcWyESyVZPDyMzaga
3yg+7DreruhufPxca5zu193MaXGS7P93IakOT0yuFs3mslusamyRjYnJOhZYhpfGy0AFwn9+Ibxo
Qk47ZIm/vMVgMqaVyvjm9m1sLHtOMtLuSBYK1niH1TMP0jUb6NseIrxW06byCUGjlSHNb253eTf6
oD2HSGVY6oSZXJYgbRtDRHSY50PrbgwwfXXBojzyGTh8wm5cnmUNARVjrv3EuLi1AKroeg2ShOKg
t0TOmmhyzhKknAXuWmUb1GQ1ZCmctJN2M2SqSTDeBZUKRnQ61zTvJ1SMPm/vjfx815GskmKMd+Pl
1gnVQWG2Hq13YHvadWw7y71hMEpK6PlrCxevCWd5wh4WaD0A0Wl0Ld+n/U5iHCWi1/+MXxuLyMzN
wjtc2g09N9wIoYh/nTLIpkEn/8KR9SAvJToKFLGwyxC4sZpD5lc6CHVCSaSr6dGSBALp6QHrStuL
JpAyObAdOJiQK3ymhMybX5q4PmL+rcTxuOQiEBI82Q2t6Ynm5Z6ZmNv153eDShhsDWuUN8+rQNBq
wToQ8D4fz4mQ9PkqQGQtdHfjEyV2vKxA/E8xQ8nlq1ke1rmpK8lUy4Oo6HWMJ+xtvKNdI7YO9ovl
ZYF26KR94SmeaAOIXpAomXIFb2ffVSzO7nVmE2qXMiswTX347fYdfRcULnget1Qr23WONOn2TIxs
8RcmR3wqNLYJLSRhVmy6YJOFhiQg64MoN2MOUl7uLr5F4a6fAbHFHaDbnTJxxjxo8wYL/G4UnFx4
ax8vYcFBmBbhLYDK30rVcM23ZGfZqFcK+hqpdG7a/FdOhmQbpuDWadnGqqEbgt6cnBrNXuYRHPm1
jWyP9ChYRLV9YMt9rrMsnJ6Y2GlqqGWb0+SZyCHIdia02quf3dzEZLcc8v204fMKn9POG+ELEVqK
CpD12S4MqalHU0PG6z6fWoxr6osoqqpq0orpDB6I+pcirjVB5rcYKm/bxgC3uPrJhcWhtJQO3oPf
xMocOcnKrUfEP90bw/bfTRe0e4sVjANMieQuhF/KIAIX4AtoXqqWZTUHG4IMfIIu4tfp+6dIhQcb
FJFyCocLPdACnGKK1/LLA6xBVhKu9KifwSfbwdNoyE8JaUXNVZ24e22S3VynJTM8jkR+7n0uJhh3
vGyuTd10ER32HxfXXxhWpM95THzFc6OMA1ExzNOBObPuNQg2ucr576tiJTXbCKxl/OHMPjURHhK1
jkvU6X5/Ebza1zGHroHiBrhKNGEuQaOVOpmyMt8eUYfT/f7Z5x2Mb/kUjQ3U6hQayUxBR+W1s/7p
p2GF/ycQG/oaQG0QK5FjUR3DW2ZdNCoVkyZvmgLXhCd6/f8ZMBwjqNFiwep6dukc3u+Pz8oHaBkA
cKAo8jXQzNNsC8QVc/GrW8TmTMssq38u0ardQFSgeHMpeUFwIyTgYBSwVOKPyAXF0JzKyFctxP4O
LgwpXhzSJh1EYRGP8tLxlAdVr5XwekOHfQXqN4GdXEF9J+yUdUhcx83OTUqFnwvRUX1Oj2Dd9fis
Jokc+XW8ZX3r4Eufd/C8pJ1E4QzGTnA9GgKaqJejM/Djer+bPV1eBOWUxh0TXLuN7Zfmaip/7ajq
0DIq6q1BhKYvThy4u23GIF3r+vNnrI/agcNFoamBlrEiyM6lg06TA8rZuCAD9tUgaOIx/9eP8btE
qOmNU/iwF2tzrg49z6tKL3NLffby1lx3nWoY9oDdsiavu0vhgSD8R/xbN7+Fukf2CMaZzoadmU52
Ci9cb4JaEU3KM6Wx0SXceCMYRtznP+j1AJJHwts3G8Ue1A/0viS5H/axjOlkJPUGkgqj46QavnBy
OEUVPz4QIrbc2wtFz42FwvT7WP+XXplU3I6iMVyfDjIT+DD5ZmxP35ymhUXMSzz3X+6cf36Ixsve
jTcvDlnKavgOpYl5GmGeY4JVnkbs6zRaFnc/OojqEVzsXQurK5yQMkdFrFkvLbeT2+n409kQPvIA
uems5NdTFWFgrGP1vPYjptOpvwfINaTt31nuSin6scJt4b0dL5iaH/k+Rs6+VUSZCm9BLjjoDUtE
rVywlZOPxIGUktQDyNNW3ppXyqeFaoI4z8gdf0949hq7kDRIrlssNS3U5vTYhN+oRTSxEP3tqie4
Ae/5wpGXV5Ysbq6/t3xt26LrEeGA4DlaQD8Vd0YnIZOfjsjooMdmA+O4oBWY+assk27BrImMfaIJ
SpZ9bzbmWZUpIVs5rwDCDQnTqLxnPM279oDXTs9O4b51iTEJIssltqXtTbWo9X82XvE5UVCjQMsZ
lQjOzurkgaYXFEv0N1YfUAYw1YK4ch7P+HZ3u394Gx7isYK/ehPxnfthLADu6P6aIQ4QIts6dQTm
hfyipjuTuwD5+ug6hFfgaY+XIexJfuhviEYdSNY0jAfdo/h1cn5+dFiTBide0TQhwnVHe/RnM86D
mBFWoruSz9PjXf5ASYl2fPmRF6nzGy3L3K44id9zesnTVsc19/xkejOVdufltAI6pjvQrh006E8s
G0GiGGZVlEXuloI8gp97Ysb/Koj+IUhay1rX18zhKX7C0nP1tPjpws/JWVcd64JiAv1IpONocZjG
IgwKA3bYVHhBQdOQQkMLp0ynppkWLZFn7j3Myefb5U/DIUOqMyl7GQZ8IQqGNMRrUquuvxLI0A6r
8+CTdm60edOvITsngUD4LO4SkqrCtYYHBUiIObZaxbbIUANGOIqTLqYmgGH+yTYr3lIU/Ab9GbLZ
A6zuXnEoo1BBZ76+bUGkP2/8CpYLA586+cArpA1yiomgdjfWNn0CxnaFFGMAlBUQ5ZeEPY7UP171
xDlykZZjsgTjYjNa4vM4KXt3lzk9VdVPrmTteAzqmwPUaPMGVJXwfTWsrF1LmF2WqvlVV3x93QtX
kA4/rHmtYW8B7KLyoRnuJ4MOGIVNgSMs5FG3KA4a5rUpdyvPt74qbB1nsGI6o9b6GdBxiWGjPDGO
EWqL2wspT3sn+NoOXHIHiPoaYXdwC8Dlu4pQaRCPlWdleqxr1NYPBuzL23zqSBw5SEAAJcjTFJli
BLEBmmac1Ldw3dLvmdj8jC4RLCbtnx3ItuFsiachTLByiy74bmTKcsEdxcBoZ7KqZ0eeF3uwZ9DK
qewKzHzU31A6a6SlCL194bf61CEmnspANYSFu6gyNWFQy/JU6IBLlK/H2pBuJLP263UpccppmuQO
FxSwCUmmyvkchLlZ4cqKQ+t6rd/iMCysqVX/tEDsk9usRd7ayhpoSsCUykWL4s75gmM7leDSu0Ge
Gz6COAWHO4Kto6zI4mAa4MKk41TSbxInUPQwAmhsP98q0JjCdMAKVmmhCUKv4ErV4k4OMTtwQCIT
rmhGIxTEXGJ1BP7AO0nxYVNMLU7AH7VE3x5gUgNHmw6Q0x6epe0ycKFYygmo1tNDIAe6+5F8Thsr
O+fqrAJKuBrborqdDyHY5cTImuyumzpNcROOZcUF+vygPnZwWJ180kZQRAQWBNT6+MRXTaF/XJFS
yULemo9eQqz+Om/L+6P8jpZsj4l2txSH1Svma63lyqGbAHXbqiMPHz5/zeskuzoGgxwJDS9zT2P9
Ise6vwcjpDiG0wQHxTBIZZFXqW8pSGc/TW7QZmO7uWbsRjIiYqpzrI1FZ0AOslThqi/VoJMpAcTZ
CB7txZbUj3k7A/IMchAqGbiwblrLlcQ6iZA+vYrc1t+757snWjgdhJ5Zvedc7cwHcyzCj8jd8d9O
+EZ0JXprAwClF6oOkXHPX/uAOCrkdu8MRWbbm0UAoU3SoVYvj1RGK0m4RvWhbno4+wng837iHHbh
npgPJ16w3iv7TY9BGi3r5EV9Tpp4N2Rh7vZCCHYsB+Zgq6znbspBtuz00qlz/vau9iVlHoC60iqk
EBllqrwpA0qmw+sPylnxKINzDBJQi7ymoxVWtjurs1Ho2YspGq/lugfFKgbpoJ4zZXCVOWqjlto9
g9tUEesk4I09Tdo21W9kL5ldS7Gfw9yb3l0DPnqbrR0jk1FyncGyyBBlVwl70HWdLNMRgEit02Ht
aAIMGhRZ7P4QPdVuqMJhWGa7CZZYAaPlo3TGNdDuc2Vq+UW7S+lg2zvoEtm5Avi6eWgax5vbRMJs
OE3zjp8m5JI3PLATLWbAONXn2MDnem6kOX95IQVFJ4jje70TJE+/5OOF6I1IerbrUzmWaDWwRmbw
zUkVO0hlX5vhyDL2gexa8bLRQBZoirHKcUU/5IK2sJAkKte7r9JkVBL7C9HiekTmkvOsPinCY+Dr
KBSFtrTuroRNfh1/6/MTa6qfF82T/+UTHGDR2x5h7JxzTYCmzs8OfpsRj7TRaDSjKfJxhO2xHexw
K4E81yx1qfTmj2wNB70hEHH3N16k3WTg2vY96G6cy25ehhaTjJTtprI13D6IHbEfMs/0B/Uh/2lr
XHW2gS/VQhtqrKruhHZhZL0E5MdjNZFH8y25G/KnrRKIhvGDd+whuS26pDqh0XC1veFxQXIyFtbo
kPseWy2WXWAcjbT45IyMUuNYTrlE55QTvI1mqeHmJYJ/mxUIopZ5QvigT+FRbvn0dYscSTRVnrVp
kYAAm4d3/s9RH1UXUjc8L2qbIp9+Xha0Da712vbm/4cM+KhoAPVzzuGXjO8RnLxvUbUzXZGy/pgd
blV1IgVDUDBywqlwcD0wB63kIa+Gm0bykuEGrFIRtrDHTPuGvKU0BscHjSV9G/knV51e6gA4kMfA
dUFhMqlaP/LmrJsoY3Oc5cdVg5m94y9ZNxzyuHsi2TGC5gDNgEdvjcjxlzhKKVqO4wo49EOtEVYR
THGS0ljHKxpt0N35KSUtKSW58wHkIwYv80GVHjwU/4z2AwmZmBEJ+ePDFfq0wFMMahpyxdE7saSn
YnCOICpQggOnndFv5r2e09jC24JphICZDQGGO7CRKziuMGP7vb8tmkqzIcinT2jqsbJssFnEPtM4
D1I3OY3bCzkqTRdBd18TlU7xYgzwTRYWFFDCYHPzXZW2WBwfMIfeIXIBUQH5xdnjSkLl/YbRyO+Q
5TcizlcDcGeDJGnIBuU9RCPrSvN5gYbwZYLX0FrG/v/ePIKvBmKneFt/zKtRRebUKi3hxvVICJDz
A6ndIbdcIsXqaQkS6iIR3poBZwehtYZFOarlbM8qspXQPUeVEelqXllHjKAUIdWiFfi9ww46KwW1
oOvIh24DioZitT2nkN4yR9y1ZPB4b0Q3jDm1UGCCclUCxVPxO+PjPm7tsg1El1iIgErcUhLqY4w9
kpcM2ug8bxC6SblFFT3KIOUTquW7ccVjWeDm6/AgjZ7E3ox5aLDodylteuJuAfFYPu5/vOuuEtBn
EI7fegSKRjzAXZyxN6npfv7zN1UgE1NDxZF3YbgkzzB3y8UivKEhQukTUcbvpFCEMjO9rTbCCrtb
N3Fhx5T0iXAToSf71RItUEuo/DkR5WlR91l2Fw98RubgRjjR+WULeshREHsQV6dMdMcAjP2gvqFa
tQ7tyaendXLhb8Ni0nuHENgHaH0R9LBKqqmxXP7nEggsq4qP5YS8VfDJyQy0itMFJm5cqUK5GuFE
3DjWj7LeiXlU9PrMB7/VM289Dcn/W4aelhujicgOp4Tv0FFjs5tuQ+maXI0Ot9YXoAxvxh+8O59a
1J6koDZ9FrNzgEMDRofurQ4LSL1NhwkP/h7M2bnipPFYYlGNnccnR3bVMfBqOuEK/keN+aCqy91X
E1imBl5QBHT45zI3pDlOh0oFTLYG9dQgKNIjeK9I5JJXvlR04VFD83rdLYnAV9TxnPP846Fzn1zt
4VzyKSaIRrGZMN+Oo4o+dE196iYH+yR0a32Rz6ymQ2lHFj4lKNVVVXIfN7R6wGce8dhvngmltSQG
Ra2x+ceZuGVcT/C9AV2Fz0LSnP2QvJ1TuCgKVacPJDBZO1toYOko7C698wZtfWKtYStzo4RyNXOB
N5euBjfm8RxY4n29EuDEhrrQ4kG/g3BWNRpnNTSKD9c8BqNsxBTfQMvGjEv6c6ScdKLmadh74gXy
5lmwYMCxZQeYc+5ajmT6Z3mzxnWMxlP7/6K/3tlfTrE/fzCb9RJ5NuYgCGTLeOn8qyKW8E5oI65n
GCd0HR7nV3DvZHdo0QmOSPn+LZAXC5y0vgGkWs8ye6ivmNxDBv2ZdjgMQ8W6N+eev4qXKlClDOGK
xgZuQMjGPUYY/Y/u1ZHa48ivYPi/MqMNAcUv5gvFV1fz7mWGzpLxa33Ymd+Tg/HfqmhHLC12KukT
30CLXTNh5/GaZMiU//riNRfv6KWsiv2ME4S9PfDPTWAKuDskkXUmd9TKtejDf+u5kXq/4r5+x2af
c/ni1vAh6U7JBn+62x5pVdvK9PX3XEbnxY4uuVXTW0rueosAv0MyEKEWnU5pAuMJ6lBUTNVtNkPF
4hUlIrWb2BxkcTeq0kLXDRx6X4m7k6IY6PEIg2An8yJRGHzWfEBFZQmZhhJSr/RvFEcRW3QD8rfw
Mut4LU8KYcWrA5fseXfTWDNqc7IYqHrsQlTKnBPVeyj4IRbjWeZhS7D3H4fuzWLNF8btkJvW0IXD
9VkcBdRF0uBvyBOAmbMmdibz9uCJTMVLeeQsaxjv0O9DbBNLT4pTF4xYvAsFdwjE6C3V7PhQ4aLX
OSjhKr/EPbiLRkRNJRCBUcxsATi5fdFlnv5Rjn7V1rLIrYbdm7DhEx/MkjAr0v/rpkphv+iiXOtB
AjXn5b2nWNtmTZAJP9NbRGe/RGHdgt16vX31qryHTfxqbRRhbE0zD9neI8Idl9p9V0enhV79i/rf
h+aHttXaf+XTvQeO2cC7RoHQxBYNh2cJRb0EKmoA7mIdmASZ2N6vicojMZ01tVJkG3HXnWSzvAYA
1Ca04Sbrj2eigGUNQ6f5/G35NCkjwiYGxbGc4Zhkr79AArGI1uY/fjR1N/sSzVczcB2yxfF82TV0
LU5SSl+pGbKzR6Zy7wfEuz/h1JjBHxp5daYXdw+GChzI6Bo5wdfFGrLzx+d6LxkDxsIoBKfyT6sm
QC/GYHEIVK7GkNvGArRLkxEQbSDq+X744xtLz37VMOSSWvyyxTZHcL/ACQSPjuHTLM+hVCZRS7Da
IKNZD6GOCn/3cbn9juNNw1WT6G28blrCJtL9Oe3W14C/8hAq82Ggyn7bv6h0d3MbqIBq9hfJupo0
Cr9l0/9HhfH8fK0wAznPUPjYiVCll6YwdYociSuxHyaLltXImX3kIi9ORnyP0yPkuBpm00iiHK+X
xV7Dw3I4gj5may60xnRk4VEBKKjjohzUHXOzSFpopKRo/xOOg4C7MYf+M9KWjzYM8iuAWEufd6R9
tQyxsv/4CuvdP1KrlJ/wrVIyNX5pbjh7yZF5sWiOw1z9LePgEIWo81XW2fZ+yaIQvqYYpZl1VOCZ
PI3AWtsLL8KlCq8zPw9QV8H4huU2D0F62ewzIAWIchaKthhpAx27ipe5qhBwTCUzPPBp4DQh0hOi
OunvF7o6lqyl+mx4MzrJljeNYAoh8cQCbjGCYtn9S9lSdICrPzplQmk/irImLlTzJpw6X8jFFcJ5
dQx9D9rjvKfcbHdP88+2Dc7f2uwSSXVFhhqSgx1I1ueI9ijWKWg7Eyk5seAP6i2nQE5lpuvvEmi2
FvCzhGNno2OW9tegoDDrejJZiuofQ8KGD6enqrVK/wZn84c4qOnvUsbowvDe7ts4URgXzIQymX5D
w1c43v4mGxnKGoJMthJCf4GFwF8cfqBSxS5WsRpTvVyFueyGHqnRwZTuqGbK7h5Egx+chhqOOewa
4GHsJj038Vi2EykpbyillhggP/DDAI7Ho0O+b+L8KMR8TLvw+COPgoNjCWwbZyY4djmUiSQShX4o
+u4GXkRr+75a5IlXtBRSq5ekXrHFpmxBc5EiQIt65NH7KjojdBsEoEtQNU34n8XxhfZDOVyYBj3p
+BvMES+kxqQimsN3xpP1ywiqyjpKZGEPX46ZWqtpNHH3ywIMZ0vjRxdJZ8XwUz5WMVCU2K6rl8GS
hapju07GrzzBlGcIUr7ldntKMxnxjyXBSmzIV7JlJkLiDaP3uAM0DKVmxZR4olN9OJiMy64QEIiy
oLgRDHibxjHhMJd6fuhl/MqkSl/sanSxhq4Z4OxTGn+Ir6gw0DmY7++effemw16VFfiQVcH1Qt6E
oMF5ZQZRVZgyuRFEqCtcE36X85crHE7hQ0Hw47FklVoKhXLIETcDwhn0v7E1FmebzXUANstbESBd
PmfyipiRu5IR9scwrKNvVR7r1IR45f4hrbaCEAh73fWe+dRhVZA4m91QygnpuANQ688A6pHf+XsZ
1aWqqG2gWzBcIK3O7msBLmCFrc4z7lm7CxK1ileBH1b0Hl0qtR9Hi9OJMeBvTSsnXQjfn1fN+hNu
9+kef2bRtjXQJzRsEKqiO8S9tnbmPix13EE9QNG+ASc1x0/tziHOwwg2EcL+IGlsvjmmHC/011Lz
rI0iRw4uD+J1jtlKy7b/x9Rm8wF8dltMDNp6gQLeI4YgclsS2VbjhKOQeJQu7sEqCTjPQzTqyGVo
puXv9veCJi71SrVIBoTPRYGqS/BLeMeiJ+cvMd8L+aOVufG85jGDJnd2Hjx0BZ+VAYsfeUv0T6kc
2rWRPg40GQYasT4JagyzQsdooF/CkLswF1NMgQMfNdE5aPvLk1tJ/eXG25id0Q3kQG8enSfflGUq
9L02Ndy0wC7v5ji31Hk01OL9UIc//Dulv+phl0sxHeMT9fR1R/0LZ5wFq2qPRd7FNoeTlY/SZMXs
DWX8V8rvGnD6glMQmHX2RqlR5VTdx+jARHiMP8C+l/Vpgtc8cCzhyvFOaW8JP1n53VI78QM/vDWs
6Hiu0mARMYvdUbo/IoPZASis/nd5Z9vmnKUyuSXKwry4K8UW6GaSwsVc9tVI8uQuQv2aykYj0Vy6
D47u3gnTgTwKXnLfnBdjDqfSVFKJoY5+QnFlHByVE+gUEwU/u7AZ6584ly92S5x0/sxVPWSjrW4S
9EbS7hKwld+VdL3MIMLT1gaG6JF/NoahaddXFGth556Wc7RnIyEm9Rl3tFUzgmxybLA4uBJqXiTw
Du/zumLBztM7MaqumbXuuKYb02xTWTpZy5n19KRrhyos4S2R223nYLHGXo5ROe1Z/cvmUG5tN4WX
0oEzvAMMbPrzWIk8BSj8Bms61sUv9IVgJYVqr5l3OECSp3cVWrutT6wfKTxrd5wlzCyR8AFzOkFx
6GvA+TsCc/6Zy6loiTWbpFiOXRnXumYt6Fec6D0DC1vmoaLc28gQ2iNXQedcPKRoNXrNm85cbJp5
Vb1IIg0OoPLqfZlw/NvgpNazVDwt8PNa5nEQkDYkkkI5lGr35SxLEBFph5OhmGNM5m3mh+i9UP0y
AW/yJUU+eIRLGaYTTDL2o0kH29h6pMHhX/vKFwPVD61l51eQ7ENHmZnAQoVLHwxsyxJKxtom3Ov/
R49xf9QCzlLu09i2QPbsond15ovc6fzwA0Of/sXpDqnYRW+YSQkjTSp+wy7Hl/DWnS2E1Kuh8XjM
nCoBheh2H2ar6cD9lY4G6+Olp6XeOXPvlebcXmDAelEpSv4YOQAzw0hxHmsoEQW4hYesvK9y5QIg
aEdBPJRH/xl3MQu2VIMeU+VESIEp95S8s5bQq+YYxTbc2UHU3zLMWlehWuhK4r+O6jVY4tOqLqNj
NZ0nBZrncmNGHRgA9L8KaF9RZw1Vl1SDD1wafdFbxxUKuwsreYXn0G/ei/Mfvpq5w9qoxPW7q39t
EVtLVKfjT0G1UoJbCeIA5sMD5FHQ9/oUNrLRDfdxoAqiYDP8x6gb/V252akNFOpVD4mB4UnHV3Tr
ZVBAzUYeK+ibFf6yN+OJUR0AGEzhJXH2D7ilrYR8IoenU7nHbqXZSGAOLl6OQG9keZu9dkVfiMKH
WA7SRyDwUigP04/MMAchlqSpPswDM+9qm+m5ClNYMnRdAOh8jaJdERicmrL8dHasDw8LWlBdaZS8
0DNZSt/5+x2I7uEQv3BgLSFJ+TAoFpA+PQEJESZl3XF5DNCu4ysq4QOpJF0IchEDTy8WNOetiQC3
mQxo31ZaXpmNf7c2ec8KxoADpIodgzMf8UVT16wlICS47y2Sc14Crpp6qeIIYx8AYa3XPTdmWvxp
0PtpZfOdPCzymUOu1cwduDYbkPaFT640mbRtmSIaVDvlXOwLMmSNz7xEka4SYtPp/XstYGb5FMco
sIKh7qIIXRHD3xzVieERCdcfSsOG4sH9TjQoSmacszy/kWx2BRNbORZnL9jOiw9Wl0yYSSLvZh+i
y9sIM6D3enCVXHcrqgW6c0oyAUvItNcsCUeDf0tYyCmdL0zRUq3I6vDvUg8ylQdBZB+Hefa1VyAw
UdS2avfYKkKmffWNVhfgB4S6DCtM6x3W9MGqvCoVe51DhRvVe0zAeLPt0BDpW2z+fzPy24wAx5Ws
rGToArbFU32h/elwl20eDz4pKRQ3TAOeNJFzXuLMT+POeBHpB91Ek8U2xIAQv5YiZyyoBR8dopo7
BXT8My/C7dyAJ5UnFuJ+haDyeNwFQo1BIEfhEuzlRb0Olqa/exf74jBw486GtwEbLTPLqsmtghRM
wCeQt8Qsmsf5aVlAdWHM2Wnhb+e4MWQQ7dmE9xhV/rtmJkAK+rE2YiIC7fzul2fskAotQFgntY5j
gjEIIT0HU5ZKthzjObCezsWYZazDGN9TiqQ9gxQ3L5hCIvcZQg4/qKzCflXeTzty8d6RWL42UlY0
WX6WzZH9mlfW+ofHEZdVYQUg7dHlVoB8qiqbVGUJ29JZyIBXeYANHE6goOp8eG5kl0umEN9V64sz
WJ8FiAU3Rj1fNM4X1+hSrX5aZLoLCY9+JOt0EG4K+zV81lnu/qma/1E3CDpMYkXhP1kZfG/BOXjH
aGYolBdNKBD5orqEP7PCw/Z1U26UjpfgLReNFn9Em3RoDL7ONWe3WPhg0xaMWuDO3dHm/YEllR9D
4XPmh5m2xjLV0ntywgM+va1t196xdrbjDMcjkgMzcb2WCeiOc1OMuC1CsRPhL96p1YEEsBF6sVYJ
9B8RwBt4TcqFGxDJov/AXP2eBMLWdp9gGdYiASC+komX3P7eeBGwyL4B+6VBAheqQvUkBssbRkvo
pY9PdZK/4iSd2XLALMN+u1B0Jjgnt7Iawt4YtmuWU6F3uQOL/5ASIjH6HkNp3wPv1OcYbg3sulOf
tYS9daM5jxFvmzvscQuMoyr22vTNWifD/pssYPkgCTb/2SmlCw/DmYGvEgyVyGZs1lJYPUtAFUQc
3l1UIlfuWSdmPtKa/8uBHRNSD1Bg9dj4gZQBOyDJbcAqdp9EYxzZvOeZRAl5uQLLbwS1TawDv2fH
RE2ylWWSiRnfvTsICVgfWPa20QcDplnfETzc8q3W9a3OxSHnlAJZ1wfHZGokh+12MYl2hLy3OB4H
bqZ3PRbLLDdeVIalaphhCKtrWjQHRBOQ4tfkt23vD3CfFfgvugXsiyEj7LF3o5J4X7OJvOWBrM8M
Tv2cMD8OCHmwN2liJrtpUx/cISgWDAdXu2mmP1M1TIX8HMb8tZEd7sWtWcZUI4I1iKumLlyJaxay
ttnEj20luY7i8X/iphU2aJR2RQAdCSazZKoNShyJyQjTihaKkgy20m6pIy0QBN7/7wgb2Q+b7Rh2
HMyagP8+iw1HN1+sk0OnqfgMSOcEohXUhGoljQT2stZ6E2ZGqKiwE49YBJGuqlaGZUXTsGWS/CXy
bLtfjI+449IPSuSEV2ezj4u0XOqtwG2n54ba8byvnpDxnBmpJnQO9xS4dYl1oZpz+YaZwd1wiIOA
KXn+iIU0gh8xLI9M7J3SEmuapOslBxTy9o10YM0/f8ksqwQb98yA4hGSwP5EOQ9QhlC5XwwNbuYr
po47LiZ61z8Y+2kwvAIu0zQf7Z6srOxNmZzYPzwqp1Qf4o8XCiiTs5qLD6oz8fm7vxr8l2GIlhYm
4PTDSKgwEjOOsgrZrzVLEqm1Jsab2EQJUEYg7gQlYh9nqaSPIK4BR94lkmzVZ9A35az3vyB1bDgK
wgzV9aYAXcAQhS6OwXTmd3bZum3CSd5/0b+otxvssTy5wS2zKgnluDaf41lmgW5TW0tG0poKB2oJ
hmcaNtwpjs1zRGo33Bn+e8b9Lbm7cq8HGiwjd9SLy2fhl5yPx1k5fIatwU0DNy5wrcKOFnj3XzIA
DHiDLbd29z+XHkyU0ArmuaebuQuga0h9dBIL7Xkg3IZd94JnvYOUomZt8lDXw0HOdcqlE3ao2n3d
7Eroo3PIGvviWZHKZaZWQQgYXNJY+PTVLMN2AQ8Ds+C8AYsOjs5sh/TXeqhLCR2F32Y0E1bQKAmH
bXL9BUiHZ7KH8HBnz2YGCEQe3XVelMPi641YP33fhAB7CGhs9EnOLTe7A2T1A0FyLC8yVnHGK24W
Lggjqy7KUkzPeTS92pD377+T//ncRrSa6Y08tqPP/7HZozyrtTyzLE5U1IdfPKSxOG8OVgbu8ShX
me3vvOlg8NTXCLNUPBcs1qjjVCEraeJPii1/Vj3u4fBZh84hLsM5NitiuhHMYwLBMQA+FizNJHH8
/WNlxg/4X79VLq8zOeE/myPZFb/FpNwHWdefRq+3AfX6Z9wpuMt7dzqg2sq7QdMaV2ue5Y1Cdh6b
JwPiuiZFSLRnNWpGUEXITCsvZx6t3OxSyNzS7JKAfUaZwS9E2e+5o1/ynt1qxZb+RpCxPqHXP3YL
dPpm0IQjfBOuQxU0PViu+ffT1FqLB5b/93JWOM3lIJ0wMHTzXVz/JyG1TUGX4G99Dyv/xZI0h/MO
weH5hGOlXKWSHA22q0wtg+wmYrD5ZdG4xqppNH7kCTaDCUi8r2dQwQWJQ8Rk/4rrXqTAadtz3Fdv
zFupdxxL1eA1tMqQOs6r9eOtZMUS7aJ438IVMlQbChM4BT/cEQ+zwxGC/2TjnD5KP2LTS7ZC+WF0
pjcnaYdKeT2/Zs/Qr+rOlsGvCmALg20yEVOCTnZB9uBxeoU8ntMCZhBXWMVHKz7FPCTsgmMy5Uj1
g6XAoTOjbdEcayWzTp4XWU13lGLh7/ojmlQ1yQEyNw/793vd7/JjaGN1DhCZgRfw2laL9kOal6Kd
k4XOfIX0xGnr7xWGHZPmYOZkaurB7uiwqqCHSYl6RRy6+M6Qs3UGIa6TPn3wG0Cnf/Nu5rtDoTIY
UzQnvVcBoTEedA27yKycEyWbizg0bS22M7vlWL9R8fVjVUNazX3xi+WaDfa+Ckzt1RFqEoWya78p
QYKs34RHXELF59v2PMQ0l9A8jvcOUSmx6fp9G9S8KzCWhawXmxSl29xEm2Cs92bjnUqMeXzeqR8Z
+JxIPi3bJIICttdzHb54xhquAVALwaUC7YqQcN1uXxZmJjRgfNJxAf+lA/0wjBpPR0uJaTQthjI5
YkR74vTlc5nVvsxyfaxl95Ut7ku4RilMCWImdN5vOtKCXAdpa5UAY+fYCALJbDdmsbgGxSXB0qmo
+YZb6Dpja2ezmXbw61fH5AZxf9xLLooByI5WGMeIGEjNilKNxq6VzLzEtjIrebv/dCtz9YGMa3pM
vVF6UjWnIcXLly8qG3XIFFdInrXSVJOZjED5zP4anLnVjmAfElPUXl8ePh8C9nPi5dPS6GwIQISl
QAmTVoAYol6kbJLbtaRggLgsh2S7BJktNZoXt331Lk2xDW4QOL7Sh+AqP1hNf8jVWv3eP+b1RXY5
RMaK1/dIsQronnZwo8yAbIFyD+7WYrGGDRX+pnBYMrpWZKUijSzkOfmMrCTdkF0Oqz1+4lM2g4ov
NWVmimE+eDPj6TYdqdqzoFKicrNcgKXfEVhP1PWgb6FdjLY1uOf+HlnMQp6ELhanTPBIvaYofZe/
IEDZNaWi9Hx23v5KtC6I4H/KO8LyY8fGwCHsaSpoCOWn42A7teyPdJMY0dRHLDAP88zG8OO/MdVf
QpAav4BQ5KM6LY80wk2Zlw4iEqQOMFjwQueACe1C2eoRCXPXnqi2kSyFo3eT95FfjxtBK2ba9fM6
xHzOmkJxFrfgpw4vtWK60XRxuV1TRF7+dDQoIx5DfqzF2GY5RW5SHRVzsKRWXzcOF5GmBbbnqOZM
VPPY26og9cCEjhQugvHEync5GdS15W5bXGMyzZjJistu1NWgkITUCvb/MAqNKsJ+MIQihiWdakKM
isRUlapbIW+m3E+k4UJrM+YhFLz2BJXy2HUBmHSzDrRD+ZYt4IChQc/0d8ms62YSv9dNv2HFEMoU
2Amm4ka6oBnIAgyvaMQ+sY7TIinHrcIZvZ8NUISdirSTYiMD6gvMmKAcBYBHZoplWzkY9Sl6k/jM
v065AZHmZnp4+i1yyS8mkoEBzZgS/t1nruDmYNeKDwV7YYDAJQQfsu/JlPdU5z9q3qSWCmK/9LyJ
sypBZrEC6mlOFuuKtqXywf+YYli7OyI9RKmNTr7sH/J9zdO1KeF51jTXMImqxxxIhN0n4Md74/sx
bn0/F3ERDI58rC+wXcXH/C5Ieio2zXCWpg9SzN8pxSLHjUDGb1jB7N7vWP6jiScEDSZUbIdtC7pc
SGgbiF4Pt6j4n3MlNfDqCU4xodCM8ek9Eavek2MS+uC6x8DeivbDjkyyOj0FOSmBypM070nczWMb
8UHHDScmFOVfFR4QUIdwaggeCdPz9Mx8pAfsc5oBpzsuM6vSrI+RuU7tAP5VDIgs7ty4YuqzscgN
TP57CngbQjDJukeAsQr1VHzEc4lcZPpyGWX4fr3y5FZ6qsZ1cP2bR5Vbn4GdiiPS6aBlWAapGGkZ
onSeqOGF/HKVMhmGPoJW3Vv2rDE6yePrNOkZtEOir7PXlrqI9VtMyE5/GxegZVXgDaJC5NSFHcYx
6m9pg17L0Z7nAPZ7XKeK13Rnf5xBNpVq96TxHTgdFK8IxQYt5DGX8WXxLuddqdWyl1zzpJd4WQzx
JTQVA6ty+lrJYBSX85idDgXhB1uLADQly9S3RBwrgtm/IdV7CcylxFnTC4x4ldFv/OnDYsMulmm1
6p+LfGBMzvS3NtAJM9g8GIS3CQdzLateOhHo0GY6RT4u2jpsnXhGsKcN1XFOEkYXUFr8YNNrT1Ey
mSLDT3Q2W2JuM2fMlsw2TLmWFy8P1yrdfRt6sOJzIBM2S8pViQEGkCjvmGkqpNs0ZlNM686FVqHJ
p4hGsTC5QRoywRfAQpmk4G+j+tkCaabVe59NRGpN6N14txv/0fOdkclylVp44nCXWtHkesvfCvDE
lyko7SVyVglRgOHxZ7nF0DMyWQuRhoyiShomioPLNgzrzmh5a8M0dC9AJ9LYsWP+lGkvE0vrZhIo
AnvKKevRM7xFvL+wdJ7LoJJqQl/xbzOHskf9RcOqQLiFgJ5N3X9yv+P48AMKplSuoDgcRSKqS2lp
vluQcAqdpctblfER2YbUwRiCwgEkjs5lmX3AgqsVTaOKxeNfN/a5yQuBXZeWt29qMrOSjFIlJTme
Y0Rle/7NoLFb/ryjzGwzIO+9oILBbjQkmbsINFIscSGP4PHL5C5e8wdnjK5KnC/l+yHO3KJyj8qK
h9RJ25qYBZoH/5QTVVYi2Nrv8w92iDuYaUlt2ClpSBihuqZ0wY75/FUvwaaEqR9o01B/bbSkF7Fw
pzQLXjFP9wpfoXWfRO76yV2WKTWb/ddLcmR0riRisRit85PLxYv+U7tKKi1Gqq3r3sGsyABK+it9
16YVmj0Gai2zk7GdQJu3lGohBcHJtSpp5zbBArhJvJozjaO7P29dkwlnnivKOYoTvnSuSJxHTX8C
aZ6OfTuFle1z5BsXlywubMqLBTBEQCIIFmBEjXUNVSFNjnugr/THMvMjzAQWmmI9VUd6dGCVYeue
NirI+lDrw5OYoyNyJGueLZGXpu6pzdVvihxQF94hluBJxUVg54U7p2Yuvtzk5qor4rsKIkvufmfT
ZaTMyYfBk3GvlQwjvRfVt2H7ONJpyeFmY6hVr5p/scsugvVvgf6R+IYWuixeOUVlqTDO3LHVRLqk
iAh06nmvmyeeu5+fAtQmth2Bi/mQOpmdjKL8qnrcME6Wax2C9SshmtCm4WICYON8U3Hza/gOiC4s
ioQPT87XJUvfZGD7+otBvDV0bCR+LmUlQ5xm9HZD76Pjd7zBd0Z2vc2rni0NLgseVnhFnTAX6pzX
mmf0nm6Ky9dwzRUSAHdCAxfAiBdXmCmKhsaRBFg1bxrr8EeJ3OpaooNp9n5L31js5tDEHFsaIy6D
bHTaRE3EtJDgC7LjTFx4HR0WlPRyZw9XA6p+N5D5gyBH/HFQrZbkbmpNLj9Oj6F0pJtHChGUl0Lt
8HoggYLOGtiLyCJiP30WdrOfAMMNn0Ciz8Nlkj7VlcOSEU04pgvGlrqv0q8i2fGWqIP3tatRoH+6
IO4b0AepB+GzuhroKY4VKAvMZ/N6qt72SB2b0V28nnIXmabc5LiAp8OwbZHjkE23CvJtX3iLR2da
fDTVBAAKK1hQQum/CQC1Fe9uPutlMSsav6B4v9Cj17D42ExztHxPXPduyyPC7VByrn2ALb6PHxdp
Re3qYu7BB1HaqhXBYOOisiw48/J+r6qyiUT48sp8FYktdM0cGxy30m9l96J8e17LHdAxTkrzufcp
cselwQj88I57Xs4Wursyc3iOiucKWMUzABm7AwkYHdCMhzTfIhrXCZd4pEp+nIBYY1EJKYSpw280
qgSxhpj65+y8rnuSxBzM5dU5Ff1E9ZXkjMUgswKvLlgxFup2j7jcLTU1vrP0H19aqTlVxT8frU6d
wzyrRqYNpRU2eU75fBeDi6uPJSziv8Maw1/Ah+RwA+pyYwBUqyt0eVeicVWzwR/SD78qCOwsEi73
PtweT3jxRBSEYPTzMWCkKb0af0ze111icy5Zf4g7ucuxT0BpaanEB5CGulnwiaMN9IhnQRemIST1
UGUp+EbqskzFBQUZ+ewqu2GL7jqZtYgqiGF4gddiBobaJJtqu+sTmL+52Rk4+yRsvJo/D2Y7nN9r
xVlEo9GaLcQC8XoMBSbEhzjaIpxD+VcI2xpaXfx/wCMXWQHHkZCcFdqp3SL8bESbrhibZU/iHZZu
/hejUzRN3Q7ZRGhK1GjIqIM3JN8hH0Tns5HFu4SEtMdKiOD8htcRTFXMyE5u+bpu4lLQNYV+vdQe
AftSWXzYNHXds1hMHgwZcYzLdvN7mnLt/Ucd84t1pjYOpzf9Xia4bAd2an5YhXdAFHjItFJJIOyq
37bOJUYyErXEkYnEOy5qvy9SZ7MHv2vywfrn2nRAIXv4NZTMK14L1EbFkTZSyWVyAWjGKZoRRjcU
P+82oXkFjAhifm2Pa4sCmNaJ7SZFSgVVpC00pUYInicLn/VpFvl2ZO/sjgkBdFbVd9Si14kff3l0
4mdfc41hoK1TN7ppKa+3R/TzhIewrqaR3W4+caCFRRDlfUM6y09RWKoZTC68dMd1b6XMi6xKpOam
qNhYA6tmFsdvqSp8xTnpNT5BQ1PIBg+XGLsOwopUz926lZW7qAeQ5krcfPBUP5lm7btzJA3fFCx7
JlM78EQx73BNNKF7qf/oBYoqbbUBaLtrR0TXMLTql1QMP0d9w3+agG8qfCSzdlaxYbGy/9WFz2XV
/zT0YcykDjxzqGCY2oamhJZnrr0E1AuKFSqRaT4LiGJOK90uby1KGrZ2ikSpJrbP5etVr4t2CifR
XhEsHn0CkmMAMHzV9Jegs5U+qQfuSwNRiWrb9h2T4WhYbo24u2Hfnn9RT4c20roULEd+u3iXob/2
ixjCx+uLZGkjHVzn4hZBybc9/6J1oIbitO9JtZHYEw1dXPBl6PkD2vHQA2xJfWbOEK7VwkPBUdPn
Z8NqRnIIijZaV9G+Ee6NsDLMP0H+FqbET+kdF7yi2eXyZRSwOyAaeENFxDBwdVvGgWnr1KkbNRDn
roQjgIGiHk+alDaQzoUW13wNvrncWQK2B3Lgny1w46OPCpqg1M+zpGq/3p2FBf1EOTJSIrSIJmA1
sl3l8b/ffg6ZJB/hC6j8ALzKYMPSDcpU/XuN1OLmF+slradvnjLbdj9wMSIwUly3q4RL2EBgSkf2
MqHe8KyH+q+MszJ4vFraEJ35hfy2TtmnGRmT6/Qd7z0BFgyjXUslglJ9a1pbD15ELycOq4CVokzB
8PU3S8uNCA5h5JVVahBsoWBtlmD0XKWNnezA+XpE+Mcuef+0eBCGkqJSHKArrzZSSGdYyVxuOKMv
cfB0SjjiG3XFBKrdjEU5n9ixFI3T5rvTpbaepAcRlvtk4RYDz9NlXiCv1ClF3QtkK3Ulx/zhbcic
CHwdF/cCH7hZu+rc2g7FpyXx7n9U1YQ6pxf12POoQBH7eTBz8OGJCd7DwQeQb+leijg0LlAtMfzV
tz03pHBjSE8ChfKd3g+PqBJy7OK0dWvsW6VtpPlrpUQp8KSjvLNui3zWEQsOO4qvPI3W+7a+W31q
hfoVt91ZddKV7DCOMM9NMf/6kdX2UQJn9/yAURkAYLtiS4AWgd0L9lTR5XmYeqegpmcb3Wn2JxF2
uE/257gUnofAiTGcrXBTJluT+gN2Wt/DcKsnF9a5SWNYATRdupm0MpJpNimyNIOtW5OtnccJmpE3
QIWadOKPK1d3CsFtAk9DtZFzlVxttyy71vlvjkmHqoR4pRJR1gjU1xiFXgwJD/RyJIqxpxHSS5uX
jWXRueWynCQD7HYY3CQPS6+hFXNrZINlaCpXMkMMGpfdJvxz5Xxk9jlqU5jpRCbSo7I9XJHVgY0b
3tRPjoTSUtbAzIOv6MfMRz3KX5irgHyv40B5ROygF34y6f6tRK3YpwGEAMCJHAJBfCG26UgT7dwz
CbUBDkRThUL5ohD65Ztr7mgJx+TJg7XEVI7oWyU105ALBXjVhIsL+0r+dkrZWkIKA6Bw2xdj4bc8
/Km7PN1vwZPL9SYM9a4lfMhwZ3THZIL4lULMo8pLCmYTN/Z/LxzhvKELpil0KdNawaX+OFzJcEbC
AfEqvpMWvAc789GyuAvGuZdkmAiNN72ahoyUZyk8TyRyOuYPAQ0JqPwXZs4JuUjoni5eF3ZD97fx
22DA/d8/4ousvKTBHrNHOq4fngZqHNB5ITDz4IdUeXVW2mxFUNhXa1EJKUaClo7mRfNYzX5BsC0n
zp+vb7CbYsi8UJM+1FcexH2n5XVvol+3sWSvUTemtM2lzgqJ0Wn7Iv/7mqYpIB3BMki38933bjyx
OZktsgAj7J2QHs4ELsX9pHo5bQV7ZpTWZYA8ZlJB5K8Zs8Aypln5UlkIuytxN8SkYVSHQkcXJrzA
nXHtFkXvn6utrzXSumACB+Jgha88pJI56+j5/JnCdSqCEwBrzHj4q9bzdZm56S6p7h0bvFzqCc/H
vtctqoT4FmEtYexRSCeFnasVYe1vJfIdZmuXSN5pDRZOho8gO7fsITZFZ7aU2O7+qeXqbW20jaFm
FDh+fptfkgw4KLNGXFEGUsTnPhhD6IbQjqplKTqmTPRF16K+gMArfY+gXFZpx/C8h4ysenFH1cQ/
EPPcR80ZDij64QxhoqOjCemV3m88WBdFCyxN5XLcjEhrRr1WrG3lk6TF7rtNuuxAUUKv1722U1iJ
7+slC/d/lcNT1IMsNzFxLToz8a8JlzXf1zoMh72Ie5x2HggT2v2CiKCn1alzNac8qmU7Jx71P2j8
ZEfl6mI2iWMXdE5SckWTwxKyOvRxg8tU3eZeBJDe80GtwAwW7dgDsE+rGvehhmMMwCDPZzNTR1iG
QBoh6qDLijJtnx9PtXB1gzsDen9jZsOoyV9ESBcVZnVXWVJWSAl7LE/T7gn9OrX+PtMwBY5uoSqn
zizHAXFrN0WFPuz8C3QqDNsphGQIfcwKQ6GknmvOvwxoeE1vYHyqkECTMcvgIOkDD5CyYrhmJ/s0
83X0K/GrqdkVVp3l1b9woutxF/IPAf8Gjlt/YwgPjJahXgrCXRk5vXVm2A2Pf60okQM3GeRQnyZx
gAPNSXi7SSKCBgAxPrmZSrOv1ttk6A2CcYJ8JhaYAukk7ttGYsyio6c3DOGCucKtlSqLnbqvvGpf
bcD+JuGYBpDlkNH4fqEkXrsBNO8p4HtJpoDFJbD3Z787xBhxy8o3ZccmeRlr2dtuFEPeXstjTL+l
VscNexJIpKb1jkgEepRxtwEDrKISDeu400kNu+YOug2pXPVcSYlUHowJ4aTARl82NdVbDhw/MXhl
HpWockfNKKr1wzh+a9+FTvfCblTzuC6cOeye3HF5qsxv/G0fVisCjpbVnyefmyDhq9TzDjzEK/cE
pMeodHJ+Gr5ZUeaBpK8N9e4uGHbHTQ/RBSir+Vpp4ww8k/xyQV9XRCEeqeanS2q3aPV7E9mhJy5R
nfj4PGRRTrelC6IJWyvxzrZtIXlaSrTWIs+KM/375Cj6MaqOWTxvFtg1ITYfi2nX20RJLF3MwJvl
S84jbtcXGUMK9Uj/IYn8HmGZ11dgjam9WxZQ3A3WsVMIRUvibbhma5fRxiPsT92W//1R2vvpm9Py
PRoFVqxtIgBbPFDB0/ss/RNuqBtvnkuURR9rwwapFqPkxJEPClahjBlZ/cSfpYGqFXoecWS2Kjbe
G3uV4qsR5KdfQcymnp73BhposFZ3KoE95v+clDMOdRFsi3tgEvdNGufciAKRAjnP4FN1P1PptSRJ
pYBsCKwjZs4xiYlDLk7bs4BQHEPzFfchMvsq7T66rVG5ImCoFHOiTFW3gnnZGfsFCfC4eyEpXM/c
Bwb5d+/doOqxr+jSNYtBdPadSy1XJBXiM1ymXaZZ5yZNfFwX2VMkKSSfWUCduZmefKUtkFqTgUMz
DGY1nWskERQx1Y1NGF5zOL12fbagcjbJqgAxQk7N6VcYZOakh1chGVhuFsZOk/SqHQ/Y4+D6dBVd
fr4kA5C5hRwk9XMnHrQBFBaAECmYLcERYEthbnlSq1nPgr4bATG/i2QutOFD5p1cESVWlM2Eu0Ee
kq/WlAFvP3n2mEuWGQ37QzsGQ0cS+dX7Avesn0XLuEXk/Hn6qOYK0/WiwBJ+humgdSblICAEw7A0
n45mpJEaVhxOGIRflW2dWARV2OBMuVB1Cd+UoD2ASBUjvO/euafkzfKZ1oFtMlMzGCfNC/xSuLvq
ZseRw49K0AvW2WiQNo2ruQ+hD4I7pCmIquHKIZ7AtN7SfkyCliN5GAtSfcb8n6HDWX9UObhOmLuq
gO0lFXRxpeorDlCSQobVnM4CtYYRJ2HeP+6ubSLN123IZlef+bW8xyTNg1S5IDhTHJktxMZYQgt4
zdbyzIgaYYxK7pYXB+eWXHtIgmN+BWIKP9OttXACXM4qY1JUvQ5VXuMGM9uQF7e3ne0ZtsdsjG/d
WnLHJNF4BgpQ6dA+sd4ef7cFNlx+OsF9Au93TUh77jx6tb71O+ZFApxRCccWC5CeBO/4UcO669ej
xYTOhb/qfdqxrHrXPr8gCyBghTqOI1vDZoQHpwB51RFdIDET5zS4+AcKJsC95PurROz7ZH+OU9vE
9XXaEPCOD4PxEv2spvWImhreyEc65N8IID2RueRaGdf/k4ZkEw5OB4vwspCLrQMwhurwh/eu9G4i
DigBxC1kdmVZwM5B4OtSRF3dKtQge6TTsbltcvDrrRrY2fOfkDicM0tygfy9HhwFY70vBPlYmdXl
wwxjePas7fqmQlGrmt5YA5dX0Ac/QnFcYro0GDm4IDsNOuKX/JkVp60ok2IheQ3I/o095sFzLfqv
lXUfigqA5tzt5kbX4PGI7/TdO8bxaYdBjAtqjbgldelJA80MEZEGpEtlUTk7hh3JgdojqzXj+oyI
FJwxjb2amoAxF4eAcqMtI7lT7PgCbDXvc2SSVgIOszHQajRgluCwygIETvVyFnuJOIkTCLOlokxG
0dqaeRCCo30g7AvibrV5MN3a+Fa0FRTT+wZt/5yecvHYOOmNWhn0/xI1LNT90P44EazcGMCZ1GX9
H75+gcA3K8iq9u2jhtmVPQxajemMfRtZ8cY9G0mnrSkoUCf5v9LdRIW3NS4SG/rpqdRZAQQN+X+y
ePJJMiDEN/K7R7NPw3T6UsqSFDMdGdZIo5GShLjlCY6mTI/JA3Z81dioZnP66mpDm95BRWk5KEtK
iukifJeMN6iRxxK/6ENaAnhPrS0brGnN/CSPAhl8s3oMmShfbHHwa306FYgtkRdDmwSPUl2Nt/Di
/BYhkAJGKUrGulH06ekL/n89pmzBE7IRK4IF+gq2W3ADNhW8nhdtqQFINgyvGJv+tXVKi4oD/Oeo
Jee9n6e9y2poaz1X0Yy5ejdNZfwnVQ0UcjrQh0NiBk9ZdeU2zIHEf6maKDD2WvoQeEx2fQCarYLQ
fEPgs01C/BtmvfEIxeGDjbshp3OjaHybO58MKFZQu+o+43z6zaqrSbEVIu6OrtttZ5/V6sYMR5BE
6LTBUJ2ibWRXqS/ghb7LKGJI4M5Hd6+3ZaAbu6EZCn484Jt7bemBeTX+BJsCAsmkIl0p4qMP/+O8
3LuKIJUUeYmEidKDr6Xlw9zcUvYainIGnAfvMsU3Sjij1v7sEg2jUsClCU8ZVyUxbNr4DOCAfFRx
IrrbcZTzxlxnAVvFjxc34BjqhbFSVIpog75vlFgF0P/9fTMpceU7aiIH9U4z+ZuE33AkKsoUtNz+
Ieq35lc4Zw6zGSA/S9hZSDUlKhlhQMttaE3TGOLLQ24kZz6h6o3my2RSo2dYQ8kmIdhPs5r1WBH+
eFrmK58ymmco1rgdRRcIV1OAyPGeDMQIIVMI2sug0zimaEWwfdAvtWTpQbi7/MKQQxkut1n8GSjd
4gL3RTZc17UKFmw/IzWFzs3PQWOluOJFK0uE0CtlWNeZ1xB0r+EOYPIK2eD7pt1x/4SsYx+AEKbW
Kq75Y+Dbb07wU1zlIcyMWzWl66t25YynNTqVRHUX1yjqm2/1wXQXnQEboxY2FPeLzhJaZBdy61Mh
2TL0hTFFRBilzBqtbjkpwMQPuQAKZsZbUUAkcqbHrdTmJWNceGS05f18e7T6Fkojk0T2nfsEqT4m
SBEsU28J4Nlf0Uc5w/fexfZWXvWho1I9isXcOeTig5bJMgXnJuTVGodhN0srxHsC/V432TmcosXe
XgNk8T02LTh6HGbFkQPi/M9IK5B3IBavUavafw7v8vH5E034j7m11Aul3PEkb/htR/bvmxmje9zJ
D2cslKnNb6LcEsmprZhXLZsvrAFy70GrLWYNdAjUdaOmK0V/MGQHQtpjEwiiSlS09Qu6rFAsnE4E
HUyX7HS9fzrPihuiP56qgA23EGGgbSwMl2Ay0nBPcWojjST14gsxaLSRNR0H6poYz1xWzpkM7U1y
FYfCRs1tZk8TErj4tzdd1KSGSg2XPhiVO+Plh8ul9v38wJW4HVU0NNcArOIv6uJNumKB/+yy3rEe
TuU4CldaV7/OY1rbfBAyxdbRBsvJuX+HCOVwLm9gqXpSOVmdRaU2DRcjJNqNlUIrVTzCJ41by/3f
tA+xCi2hMsCak1vPLUulh8KjJ8k1mFehMUjTJzPkNh/qsy1rtY4gPInArZkbrVYzE6zxAyAwJS5H
VFWLYr5fgloCgsIUXCTxS6wLVlQHPEcVrpJfnMWz+KKTFb9dsem7CmA/+QuQjx7ihTt8570/1yvH
zBpckooIB0UkHrmulGUxxTSzEpuC/NAwQUkb+P4Y69ybmf9r24t97nz4wiPgMaI0+2VPjn3KUDBH
UGfUZiFNJgzxCttfvsZQR+QcFv+6dsGXWihlE2UuBgk6UwpRg/K3j4J1Bfmv5ixvD1o92A+/2s+f
/XMPlm/jrXXrlX3r70a3FslA39Ol/2VuI9J+ks+C0V9KrHmPDo5Ut8iHrFnh5A87ynJzrgB9zzI6
1QZV2auFyXSH6n27IgL/lA0pfxyOCusr4yV+6SgzlIqRE2eS0uZAo3343fymUxtKywnWCD2Zhw7T
qcHcfwtc4XHYmlEEK4ym6b7slUJaVJT3Wdg++CAd/QAj9iz91tN6EMEpQnErvdy3McA9FqxuW9mE
PlVD5u1qmNSQ7lajL/OCNYYtxokHsrXACnH5mPnceQ88w8seSOr17xYTW7QZI7kEpmfQsJWPn775
MYBlX3cQUU4eWSZsfNl9G99M/kpT2z3XaE4da0YX9PS/MMbPbRGLJoaGTVSfJiQE/L+EYFi3bFTR
tsDUKM59nKGeEgO9xKNLYNqfG8QHdOd8MYWBqzWiJG4hGGqWlEH700zqfRDQXooTE+omR6qNaLS3
xTJgoVHaTWZluB+7nH0IDvcW7zQ2By9/uhagZcNxsLBcx7hukdpUsL97aE6xCx2Wk/gUKMKRrKEb
DCi9qL8o1zcMe7s2HRyDBkDzwP2evQxpgAE2Q0GVNly1TWTCeVsbTm0jftiApBODPh/FLRznd2Um
4yiovbSEXdZkMn3wg2jhj1JyhNKTkweqh0MxG03uLcnlxT63zx+WzQVW2s3mcIO6U/2dRH9YniS0
RLZRZoyNrkgQSmoRvszt2x+bsYc0SFAMLasdk16Yb9bkj7mz2DxByc2lMD+che3bHje8tu/GVqDa
LUwRODiMbutEYL3sndTu0AyLsX/lvgIiQhjEkEzZ+Xvyg/3b/Y38jkFuf94Xl5fN1+ym1dyPjyCj
vxKF2/rJrgCQ60Cw7fXGFF1kcUNkEPCvFb3da0XyUZ/JzAcUD7HJRXcw+emhigpeS1CkajFJugFZ
2HlE2SqDTKKGAk+qMZRrcfsO8ivX8KcOH7m/WVoGeaQBFjZvn20s1jwqptFWObXXf8munpF2WERy
kkOwS7sFM2s7w9+zmwz2Isu/XJix3bFuWywR+ELfOy20kcjaF+l10PwgtBnpooFmjG6zwjvwXYDp
59MVgcHbjeDGvImgw3CIWf23Of1w9VgwLbkQO/mpAGBOhcv8zSy/G/EgZ4hZKfNqGUsaaODq6Oeo
6x0Ix3ur2lnqidFcv+XkLsLR+1BdTHFabJaB6MMR2NOSYg1P61pXeu2biokdIq1VsER3JqEABZWi
OkPWuZyLX6yx0FxpTTRxv2XQOVe/nz3nowUWaiKW1M85hnZqseke8m9cxE6oWUz3J09j0pUEJuXN
AdUPiewiRV6MoNT1c+sm5QTIDCZfrtGoJHDFh8XsY34aGta+6hOQE3f7M28ZD5QqQnRBr+XAzDjj
7/y5rgzJm3K5FydbMJLqOmkGe4B9WYS9oc7EX03mqxAYz6H9Fts+oALbcUvVy9rrmfRZuqQKPZZg
oRkBtOEqLr2nEXolwS64NX6TbHDAsJAhBUcofdBjv5zoiN9jIzDq7mRaD/LJv+pP5zGNB8o/9j9a
Ag9lSLqx8XBzzIB9ffgYws2gZ5MMjXDaYf9EKipp2nw10jCyttrYCM1DoNMEecv0uJPpvvV2e1d4
dD3SCCKk4lU+9f2KgzBUoy3jtpfcbDZxB3VQTvc4MLjqkKqOHLZ6I1IlABVsftKBH0tMVYfRrifI
cDHXKAneOMJPpcZDifE0PwSTStPnkSCgXyvRwxY0+R7jsC6PM26N2RvwlX7Zwd8kP1H0zklX+wbF
5h83zwQKoqo++I102jqy/syWEm4ZjnJmlscVDozoZQyiNDMHPAA4I4DpMliA1CFHYP5RBZxjOTxY
J7Up5aLepfRNonl8jQdGZghJ5JvvLdLUGLenjuuFNSgN1xpp89VA0pRUHbq3DTAztWeQpN1H+/kp
rNMgG1SxH41IZEN75M1G/4wc0M77Etf/8Lsb6nKzsP3XSKO9rb21y25EX1aLlkq1zflv7qvVsJTO
lLJC46V0AjR0PylkLy57SZBt9/x9Addk1ByJ6MBjx7xaJ9dGjqJvDMQWhiEC7Yagi3KA8zG1OAVy
cSob8/XoGvUMhthB4RR6FqYGEb7GjmERjdbg8ggLH8TQK156xtA2Gmdh2VJjkcbMVGS36HOBPvii
N2C3mGOpqDOPd1k8XzMVT2r675oEe0F8yhjeGvzT0PTIJPU7oL25uuiCQcBANOxocR3cltlWK+33
ZxteaHHZWm0NidX9dTURJpklVokdllTkV5nB9Htx9/hCH0y4m7ulGqhbqs2r/OrihTqPkKykQZPG
VDbzt5W9ESV9wBaLimiRpbimm+21u37ta89QjRI1CzM/8DNFzRFwbmNFZqT8oOCmRCFcHItObq6X
sB8yC/fANnKFrfiBU+TLt6s+TJwu3bLbtB9CxacIt0sfVfGRBXBvnxhRAbhCDEW4xlw9mqnQMtHI
CGY+n9mWqdNfExkVbeIgjueQTnxu4gUSJVEzT8tv1FGLHP9xQu7U81PHIhrfpybgQgmP3fabK8ie
V5DPd6g8cvGCRHFYkfAQW7VtM8bYIizT5SVsdXqORhfPhxh+tmsJnC45jOgjiTen60hadyao7/Mu
PY9fQrlXhG8UDsv46TWkzHMf+lq/aF1vxl14Pvp35D0Lq5NglPitXdiN3R77yx+YNdHmfeiVJ4yW
drKc+F/4G4msLOihK64Lb1dfux9ldhUzSoA7puogwGP7yoH3q/61r9lAaL2LVg6MqBQTezXdgyAF
i89u9BjIuVDYnDW35kcTXf9wYIfLCOs9eYWh3L8fjQmMbQerQ2zyldHe6EI2XrPUdweS7Ya2AkAC
7PR9DxGcXLywAW7eMaFntMt9TG9ewFLfqNlswO89Lyd9Wv+/i/ui/zmlp3TQTeuUxS3Bie801Rs3
MQYghNdPm1VxzV6Scv/6ZO+f3VIIkW7eZXxPNWv6RPxI8vDMJGXHB4sm+JL7k+EfQA+ASfKRRBfT
xoej5v8yYG7XK8PhT1pIBk/H0haIdQkLiqWhdACKBwToKoNDe30ms5ZgMDYdEwtsexvX1ATVnB3H
QadOIItVQks6szVPzvJU8jeLS2UTvw+8JDzRlb4e/vOEuSXxFOP7aR7sJXB8CY/eM3nEZV3Bsuy3
nyH1k+5TUlW92+KptUjeuf70PjvqqcL9rZSqznTDHyP54LS3tzH0yhxbSfMYvhw87OZDu4gkj9Ia
EpVXk+uFNzku8Rn+RRkiDX9TmuC+A2oR1uuBae8uT1+J55XkeMx5ZWW0Y/mNc81X1qE7NRUfnV9u
1Qvp9sWaOaLSv/l2l/qc8LPfjoEVAi62jkt3t4VFwxEq1tA6WJw0lF6oK0u6zfKYhqx6XOtkoNja
p57liUUpaGMc8QIY3Od2gyj6Vl57qzTakfHP03Dsx4wCyCX/hB8qCGuV105aoFphLZzOwOihpgb7
bPpC7jmaW8GnZAOlSoFu9TpPcGopTGX3QKu5YaD9rvYvbmFGtlXfN7FaNMD79c3Ls3r8CCyTycae
RZPsnkNTOuvYw8QK7Sjy6e/wic2tSpsTd3SANnrqgmrH+5zbX3NOWijbGCvKj9eFDQyS2gPjjS5w
m99w0tSZ5MRRfVwJNNHosgunt7kdoapIaS0m5fBtgSPOfhs/hsjaGbUpVnv1ylD4ogrU22i7ZTUh
s7AwEQnMGWvlRJ8ro/3s66mgpPS0yMfkkka65HRFrJ8bys7EOzwUQAY9HOTPZFiZCQA+C55Z0XSE
L8vg5G3lwlXdjOTTW/csqdy64Go3Kz4HJpSwzFoaAqt26HIu0dQ54pbaw9Q+lvyYpYSoMQ0DOqCc
oolOAQq/VWK12Kptk0py6VLYs+A2vsp0g1gruFGZJFZseR2xpNLkiGZ2oVscrIkrYxdZ8Uzid3V8
tLMadTgbm2c1XYpnnK2ehoXXa3AQjomko061qK/bqoiSc9AqjvSfoSPUEOV5Sjdtyd/cvbuqAsie
dY99XSIxNltTzfIDHt8vf0eb36kbLOdxLc2ugKHEZ5tCJc7Ql1aUNjEdlKzH3O468CKX9H2KieKG
Du7e+XPnE2O0kjPHIQ2+i+H6miUa/JWub567ImLctFnx/nb9l72GAZBPbiX1DMj5R2XBagfP1gTa
nEYmtxsc47Xzs1aCj9AvTt/e/htKt7EsJ4gG+xmyjK7g0D4FfPBrcbY7jqhx3UN2DA0Gh5UtKgL9
/uZe4jDZXuA5GHGhLXH0snXbSFRb4hUb0keuhXEjQLsrLHQCKg3dSEAT9QLXXi1QXjIwMDNxXBuD
CbttwTGaEwep7RKBBbpOD9S/zgDJ7JB42I8koEDRFhfOv0w5ZqfNEb/ea3NsR70KJ2VUbvgdQNnf
0/sEkjf19sWJs8/XkPnazgcMmiIcolgEAMd+puCq8AeZLslbjY1bjE3k8Di1CN4eiTQRV2UTMSgm
WrIzXAXKWSqaPNaWjb5USgkVealTJOhC/wuervjNczfAxVAFb9ckWHZRYmxM+IwCoxbx5MBIH+HS
J3/WjY+4NQpk9f42Kl0CVBLV4BJQB8Iz3DwA/3SxD22IxPF16VuHb0YJawObWQvpP/lvVHhxBgY5
lAQ1KcFjZqJGTJWvNMXhtlNMYjD5HmBp3XD2l42Hao/1bUCiLFfl39QoFidCtzv2169YzirXtXhV
OKFgQO+FmWKHbQioVqaHDp7U1keLqFDBsdnQjk8dN4DGm2zva7idHSTDY9aQGeBCKK8GEXEIQ15i
z1tGAX5Zc+md6R0eDrhHdR5p0VOrtRoD0cefSE49KK7PVHEvkZL7EOs8we56ab2b9VeVZ+1dnpX1
DNjAsumpqs/tU0u2V/0fGyFJmSQnkA/HBYaC7PQjPpVXZE9zl2+OhowuEYnZRXCNjq0jbKmRaRbP
bmtveIY+vhiTqZEXh1K5rVn9uTKZpr8TCM8juCz0l2gfZOy982uTX6N5QqnJST5t9fQgvtNBbOSQ
ofOZiwR9VhFk+Al8ghaLaZ032rj2hkQVB9yRJ2O4uBJy5aYecrHei+QDYeUCK5mSkYXTVL/PCGrf
NRxLs0nSLVyYQJ6IgbrOZseXy5PQmo5HRpzfUXWwq76Rg+diSh/bXdQZrpFWOd6IuUd4wS09aORs
HcuJuzk3q5CqBmolT0HesVlN4GJ4aNM89JBsr0Lg9pOr9Aa4KM3whtfX1p4kNWnKM0dGsA80AOXQ
45fOAnGpPAyL0yTFXf/QejGgJIkPWOEQMHaaR8WGeF6QYZ9jEEKZ46LPSP73+xjrnZXraUKOegNc
fnIr1FEter5TQIbUUNOCqDpoqKnF06KV12uWLnsGSHSg24XOoEXzKzS/adOZnvqOQYs3QE6nJdLb
kL7OkKNexrAyLSGZGxl/RDBO5amkuaUc+20gad+grTAjPbYJNXFt+pIwFOd8Gm+kh/jnIdRIjCKW
HeFP2weWr70eZFky236j4XA1sq5+Y8t2uUFwdUqgtojT97ppHlDuwtnU6vwz0RtgEevzPgGdis5C
OXSQ4X+conAmLecO6iby1cmDmNr2IME0lt1x5Vi8GIHYQJHs9qEQxDbEywzLythPrqfpgqYLLF1t
uTGUD3uMkPrIYZXZNs8G/GQ5PRELc2TV2uSupZtZRMDMxXd81/OU25D06LcLYmRwc2Z2hd+Mcixs
/bhYDkq7hT6o2dl3sGUdJoeBmxFk+EBakJhJlm7WvM1tRoOsWP4dzZSjVkm1UiDyPK33sLispvER
akmmkDDuzoRP7xmEUILfitM2BirTzcnsXAG+kjrer+AJ12dBeG6ArnvfTfQma069OhUf9bUCvKrK
z3n0LZ4SNhLw+doo4HjlGQdH5kUvUVe/kyAsB85oj2o4Z8gnbOhjMAp5lJLNl+VRfPWuzjwzNxAr
VUgTzcO8/LTpuoSdb0U1RPABVdXPI+QPo5DWKkS365dbAVfp30u59fm6QJu17GaZHgunOuph9JFY
pDdlKxpvmyz+K9JK00nGL9yX6ukZIYTAxM/xbhpEl0UfvipSnnVqoPzUpT7p1AZwAEo/My7Jg/82
Glwi9mvQj8M+0Cevy5PiJSYi6/LBmJjnSGILnpjfS/EKYIB0fH3swOrYIoiqKHTx9jzriYKVo1pf
NUuC+1Yct3dUtqWCPUnniuDK3zasHXHjw7a2av/0IXHJeWGusYZ6/NBSYfmczPrleBD/Bk5zQavG
vyKcuUFM5jhNpOmuZ+X8DCCs9pkylzdXQUvkSsYpsOf3WAxet7qcP5ZeDt02VHifCxmC+usRfbKf
GAq30KhPW5NbaLIE/4CIkQwGBp2vViPQCgyT8PApAjxV8IcE/cy8vP8oH9O5jpSX4yhEOaqT78K7
h2+9rOcwDPNF+tb5sHdJw3/ztfaGvBjmIzzkP/Mm0gVLmYCyTO955Fa/iq6i6wItpdJyYuXCOqTD
ED+oXxPp/NxrQGwFetogcOwt9zQFz3s7VdzSGU6woO7Dt//wsEYJ9omEb5tyPKplSfSk+lo2yxUD
MS55a3OU5xWD+VWQhIMwLrA7D7PrIEH47KE29lt3Tng6IEcm8dxZkDUK7+biO0bNz2HHOO8BDuPE
pgrPDRiW3besYbJQq1V8yrBPyCefyoYUuDv7M3cPw1mnZPac8DqMxEDMtw1xzOkzyvWPPqu88OM7
AF+DYC5eweEVIrHxswXVtjtyZq29oym7FDtwcXj8tjmCIYUqssJK7DbtEerSdl5Q65bTRP81veTu
eZ8QF2pTpvlCdrxu4tAXQP3b9JaneEH1uRzXD7UQEuPeRrxu0vgAoUCjApDbm/wzDDuLVyQriufW
leoem+4odmtfSZrHrhKCOdJ/1Lud0AwiyQCbrQ4Har3bV3DRq4QnE7JDgBWxCTaG5SXJUgcFODMC
GojPjtfYdlLJvJu88CsdqTNxvBJlDGAIMLHub7PyLRf6oCitQ+T9uiu1IPjg+edOhJlMHqp+XZ1Z
qqfIW+xIeos97VbShEMjD4UtCrFsLUNhPUz/zx+Znbdfse88WqUrF+sTmJbgY2vLdNSkr0k0gcKH
YUZKLVtLuOXJRbm8wt7otH4ieuXD8jLSLX88Z++2xmU0i+ZkCdhW08jxTluc+h1Mjx0RwSzjUY28
KyqHfpy0bWcYUCI00NwEwRoAJAVNPiZC55PHgtJ+jVFB19xB05Xiwz870G1R7ZgLhgFJ7Y/A+ubw
/cpXxBA1D+8OEGLrsUBYPhK/5CD4ogzDoQPIZp1k8IcWboN+b2vVknleV55XiYQ+cbfojxHcqtai
la5uj6P14jsUUhXgJOJONthhprgCHnKuRR+RlGJW0qkuzoOUiJVZw5yBaL3G3Ltw9SCl1DwikuzS
kKu6gD1iHLv1+sW2fNl2IXr7zR/GTg2To5zZ5Ntzz3NB9kB1fRb6JgykGFllwspFpMLI3smoPuS4
BuVWxELdsDVkWIjrK3LPWXC3058Cx5C3LJ1IpoBtoG0mETBOkLcyVyzl6QCB3mLLBBwG/MJoFrkG
jjzX9vsSR/Q+GeYmmFscMQhIW7iZuoanwrioc9TLhRgLnjL73/IKvpKr6abxxrknS8TnTrWXptpy
WygU+P4gAX1lhW/ozCTQF7IeM9IC6z4sTJHGQ+jbUzlGP8mUW9kyAcyPIiuqrVqY/m8/RRvksM0W
EZX0mQ/bLTbQnIEeodTxkAVirjU+fgZ0SehSpxaQOETlF3lUbwQKEHCVxyGZorZnkUF7Mv2MyJ93
PXtJod5pkvqdtCCMrpI79rU02aqzrA5DHYfa5g1eF2i5am6QgboOtnp6ldFXqRtwn1fCGVPRpkHD
+Y6eZmh3VY2Ou7YA5ERwos2f8ylMJ9HYdPSgW1sH+SSkNqPW/r9b60p+HiBrbwBJKOg+rZ25a1wP
y3bEGYgh8fMsVtzzYvCJDqQU+aIb+IbVgoeFs2fFgFotXio+r/jawmO8MCTyqWdOz3Tj0GDBuGDM
+5WIaWStVtJJnJ5rjN8HWDykHW8tcmHTJEH7weX3S5cPXG1Iu1rVwUXEObQJ0p1KHMKp9k0Dox/t
KuH8FQSzuLFVTFbMD5DG5yAKsj/OWuVx9Qkrtzr/kF3ptCV3KZIAiRnsUm6yIe+y/zNSPc+tu5Al
gD6ZpNf2wCnHDlEabhWIiDCELOX72wtUMgwjoo+45FK9Ak9WgtOTrDe6eYWBVagLcXAtqGdSYyMO
uRh8X6Rfk5gIuvmiq13H7gOZrWMAS+ozYB6Ze/in34lEj/qN8LXtdPth0kkL2rqolZ7S4UzIMisq
z2VOB1GPnU7TXxBJD4bh+mAgzTvvYhTqlTOHfkGptbdf65S+6LmZwXUH1DEX4faQ1WWDI8nwNPt/
IMYrt+3Kku3vCtKEz5pTFiFGfLrNFFjBGYfc77kdXAjSc+/aauQyo84XguZVcQsszJcuP4KRcosp
cxYR7cHSc1W6VeNemNsWZDrz7Hw54fL5ol8cYOaNBYdBjsJWlELX4s0NlkEjk1siA0eyvNif4Lrf
Wr1Mo9aqM4+OPP3iwlM1iizvzxJE0ELWxyrGuDgELPvlsK458YRu8uuzct1OWcKhCITo0ckfLWZ5
p2DGleKLTZ9/uZEQUkIDOfuLOY/5LRoRR6ODVYcmPCroO6xjtgVhXaj4XrNCUyXZClwMbGIm/XRF
wpMnf1/20BGuxEdXsuJJfCuC1z4Q4tMpkfP9ZhSfUj2IPpoxPsyjHGN76IVeOiiY9Gq3VLyYXtmn
xMW5rBZKjIKseX/UjOoY8Qtu3uEOkoDkyKBCZabT3iFy9MsqSUY1UtlUB0L9Mt7oa6rEP2qPap1F
tTqATdoFAey6iSTtrR+qD4LMT2hqnlIlTFSuGh6DHqLa64iBFV1LZQm7OOjP9PH8+F0MPQGHHmqF
+SPJCq8le5iIZBl5CJeC2gxPP9K02u2/45oC/61oRl0Tp2ALmU9gAIqz3R6vh3uR+FodEiGOOTZu
qDPxN4WR4Cmq6tLsZVKXeRrrVmMgC6VZas9sQTaPoyay+O5gMIEm3oTlFR6tNSGRyMo7xOqDEfQ3
rVirWqkeLHeCTVNlkiKO3VY8nh43FXASScWQKRv6kmPLLNUf1YjS386wtp0uDiDDmUZ4tMy/54Zp
+9tGF3//x+yDnvLcWR37yD6kNqqKXbEFdGISX3i5vp13iZpQG+vvbhPmfGkDbacHl3mW8Igw5Xvl
Ei7PswgijQpuFjJxgwlSGJHJOBueVOHroH6zFwKnafsiWS9z3pyMdFxIMIQ03HktjjtHM5tUdZN4
QhMgLB+Q+oBjLPsTOJdqoDMM2ClxTXyXytZNnJ+VXgFtnSClybfV5V2VZtKk2TZc3nky94DfYwem
MW1zrirONlMD5FKGmKDCXHotL2LwUcxF/AwpGrU/dP7sBFyW8a2MI/cVdow0JqNkdpLr5tEJuE+I
TNvI3WZMzDNpgl90eNHCGVu4tDruye0PcJRo7O3/JBD0H9nK2oUzRP6cWAJ9bESA/c6ip64KZaNc
aoam+c3OIKeKkZlcThrAnFebWPCBb4DBiZTXhXa/Os7QS67lJBF100teM4xCJVrc/t9uVi7gGvN0
QZkxyhe06rzZbnB0L4Kzb9YmQrox25K0TGgz7WTUNBTeizNZl0n73pW3ZZfT0QaattPPDUFH9qWi
HOmxkkD2ek0MZ17+Oz/FSpHVXzdn3IfB3eZ2NV9ZeLa2iRvrfqrjEGH6ngfe3pY5wHAqQabfUR4m
zwYCfYx63ebCnW5hRANmvYbmNUteJi1fmdd9pqfwf/hBx+wKGue5MqUCABSxDG4PUlifWcvj58RB
+aQALOnTg5z5h63nYgqKyde3DYW0vgAB73JdGdhzmGLHb6j1OlYl2X8hT3bXa8WrQmBSwIctm/qV
g/SeV4ShQ4ykdPJtbxZm/8ZVm1YDDrDAITMj18ix+aYLs3XUe8e37eA405valvF+ic4H0YQvrbUK
OvBV9WfCDigupRgrxreePG3ebwovBgy4vXLRcfg8oIQCPVm/yEE+YhFi3P5wtDUJhGfbJH2ox//k
Tk1xn9/navaPPVtAFJ8soW99jhvC/yj0Vqry7beIrKrwWRjma6wmXe21C/d5uD9XTVZGUJ4onrMR
+4cCwjTxj8XM04sAw/TyxxQrdmHb+Li32fwyIOFNKrKIVEm8UUTZyvFjeWJtMER0lw0yCqN01V7P
2ua8fflgNUEC4NSGnlXO35gCtkYhcap5hfIWrvIaAaUCjIU7k/Wf/Oraxr/4z11cRxtz1r8wCgky
sXr5utYYSu9Ax0uMImQrw4H2tO0MluFo5GGrXADtVjjUcc0n7Fdw9zjE4xe94rymfU/D8UZ2uMnh
QCAkSbZpknPhoNQxa5OFs856ALkNmPNdBOooziGoaYtLZivPvgI32f3oux2XcqVXCxv3OAFDo47Y
jxAzZisDhAHmNY+yyUcN+ppOrkqkg+iZ+oULG+istGXVAPlGLmQKV+oPF7RFBoLJUWsWC/NyfOfV
GP6eROjj48M3vY8UIrtyEIytaEsTPRCDzt9ttPbJG3X7Yr/NQ0icyAvLQ7Qf3pLgFU24rNQbYM6t
G1Bzi3coSlytHIfFJYg23pPXd1rvMsVNk/VA8CZWSn0ZUXi46OMiLjsC19bHchjoV5IHk39fG08w
frZluuqHvSoQzkRvIjPL5Sk9BeeY216pgkp16M60Pg39M/Yv8OfeDAOqHVLF5U2p0ImxglqDQ98e
9/kMYbkpPY3baL+Wdc1J1QqWMmSlImrIpSAfRWbTRtRsurBZSkONfpjTewSwpoAuhqZa1VMozfKk
p5NFd1O6B3yi0V/kT7oQhMmNdtCSwbz3836z60F3GmGkiLWdrM0N+YPUZz3JiN4HQZ8nL87mVRZF
KhKzLg01vi6EYCk5KqU7KqfE0MrojlJNDeV2DnIyzFqBGXtLTYetDcZbTOn57+dA36E/UU70EBLB
pnDfYGZXSBeXfX1wVDzbX1BA3Qw4EDKoI4h/7HH8t2TaHfD1AXvuz0XPh8z0evLAmQ1iLLiGj5Eg
uTieB9P9QRXCllu3qUhIc4tLOsBFPXN0DeLPAVT9HVFFqkYNQUBRqi2MjwYCYXV2+Bz0C/Nayq1b
KGlPd3MU+YEp9qnNlcNASd5Hx37Sre1P4+eCguLzaPdTWAZj9xlNeW9GdhmopJ2eem0FPAUBG0yu
hzq12rolbfBn1jnEAuF2WMVpEQNg9Go0rspv+vCwqzqGR+v4EMxIqjtUCEcweXARqKPMLXhH0bjh
ZyG3RytLGB79XQUoDC+xdZWjBc0wEe/SawNjREvzxFBCTF18CbUir/r+o1x2QWDsfZ2dHCSj72jC
4j2pnHNNKvyu6YkA/BhT8ZuOwmRRH6CEEO6Tk1xTas+XZhhRUUT0pxzcN9YabUUyWkxKEMYGn7KJ
I8JQLcbQBEC7T8hMYF+JyOSCdviJBSmMOrJgFdYxHvEUDyq0ponQgFOacRYn2SZ6Ja09Nw/+LHmc
FEyF00ZVayvDJXslDtlR5Gu5izR3ITw2Cz0l0hZUQhlYRQU1UeIKBlLHNy0LPzFdIFS5snDasusJ
JwBp7PNnmmvdd64dWTNRpKIJt5S4vtvHWTZ5tpucEuszkHjoG8Jl9ICNeLeGD3lKax7Vo27Kkd6p
MPwApyuMw6wAfxtOnB0qyAPdgrt6nt6qU6W0LvZ7mtTc1oxLLWxEZh/FTXzxnoMwK/3t8IoVUwYC
PuX6Yzp3rlv9YKP9S45OV+f4ckoSRjrCvae2n0PFEbLuctEuQNqx2bUIhgvMoHc8pQ6WBEyUNu+K
0PdrYdmn+Bnp6s114h8lfGiksB1/po9HyJhmhwZGaJMMjEeLa/nUq/j7kjE+jMwpPaw8c+OUHNWV
5tduhBvqD3ca3WwTXnaSGQ7SPeWJeoSXEJREZXmvscZDmyBsIyP8TheLu3Aqv+jP6FU0aWDSC1n9
h9FtbOrIxJ1D8zJ/ewP5of0qYcOBE40jG3W9hTxhj3L/unfboP/YzYcJfb2vpA5qr9ZdqczgTxAC
8ha6Q1Xd6tUEFNK1pavOIcMQg9hPOW+spdSUYhg4c6Skey7RqN9w2FDitsxJCyIaF0OUKQ9TAPyE
NvfNbeFWWo9wgFn8Jo2riZLxZTY9w44O8ilPMPsni4kK6WZhKLBkY2qf7fkFeJ4kZLVUC9PWbatB
ej+urn6mkmKQwaOvk/HVYs2CQFmJNcCV3bK9AZH5COBXasl9qOYKiF86hZR/KhnE0fKd2NIr2mkv
lJOIDO+JCz8H4uwN9iZf3I/wI0ef3Sw+WIhEU2bXvM54cbN+cHu0AYO99u5KsjcIA7Q1/Ks6XvVv
B9ytBwmlNivFtCErryAwitaWdjOr3wq9Vc9Yv0t/Cm3KPWxXqaBSmM/EIRQcxZoUM/XaTg1q4sC5
TO5D3OA6QSshR4tES5PZzZQh1MXYQ6Fl5IgE8f5vrghbAid39nGrgMhPNK4nNeb75WWazJx23VJV
geGpLmSHk+V/GmAs/OuBw6dL6Ysawd3AEJJhSQwUE/WHDaTecbr2kAqbZ27RtcabNUUr+cJXvwhN
Ozfm6a/coCL9fqi2VyQj664YM8sT0DhRjbJ/XbELALC4Y/B5rTcHSD7k48/zaxmRXO3hzFo97hut
8bRf7SZng5Iapz55424W9qqi5H9z1lE15O8A7pPyx/M4VJ2dMquKPGFUH+KkHsREsW/6wby9dcNn
hKk2+8x2aAsYSehYq6kV2USoC/gVWaidw7MyeSnbeIqY6Sur/t7hknyv4l/rXWnGxeEHGtk1WKId
6D1miNNPR0V9aHN0yqLL9MEmnK4xw8qrGxa2uD3hbz1ISXtATpoJO61Ah6tdlX9EbdjXXOGQORi0
l96mCZiH62Z9brm6YtKfQznzXWXYn2o50BQ+WP0ciTq7jTtPqhL6QSuHUnjmbYRzctSZqWyT43X/
lvOooZRbgNFUTGWia5ZnNWoVDY0dU3kbJJ0p0Y9e9D1u3Hc57K7WvzoCAZdZVIMgeKH8CkIPqEYK
4IxYmxnDpXPrGExW7nQs/lMCWezQxAPVKHHpgdQl9AZ8PhR65B8f5SGhlUNlVSdkLG9yQEPV7nsT
/W1OBc0RVBzbmVyvW8Nhn5QpLjuvHGEja2PpJ6R/ynZ9seSR0b+eUDhgUGXbyq6vdV0tVasdwgPs
Bzx45XgAuRd34rNxSWZWInZOWnAVbDJe2uzqWKEjeSQ2De4OpQ4nXGnL5F6iMDkOWDbf2opBlvJn
oJ/HZSkXxVCb9rKgCsGtr2tEaRxfids6RZAkMPBaLzPXwJOe1+ZlUnejQQQ5j2YL3DBVf3btlC18
n8p3Qpf4N0adg+/E2uf9Vnm7ZHCVlkY+YjI4OrBZVRS0zLMI2ZdEMzBdam3Qs9o6n8xUfRA7C0dR
q0Knb72plxKphfWooxhs4x3QBgY1NCTtk79gYYibWYluISpONemrEPRJTf2xIg9/GkVTb/6KnIlU
fXFweFJrqlAt9rJzRrU+ugs9jPmRWyyfiQIMg7cLh/W8fDufoHsNEKQCoEhRuQzMLsojqLyy5WeU
/hc8xZVp3TQPE65IgpEOnQf6wHODagJ2AKNUxrf5InrB9tnl46GRlq7D20drrnBWJtbNwDeZt7jE
IADyXHjXXYmrF5B63K5TdeVFJ3SDl0DDvj7Oyj4tXquz0KMg5+tSJTWceSIsh8jfsrfDOBTt7JUQ
/2rU2JmYWAZxlUjs8OTijjopUhhRe7hUTDG8aJ8THJBpARUUq64BSuGG1HONoENpIiUk8js203ml
lqMCNcTX+jcEaopD/Xcev2bsZlRhaIeSPobwT2S/Sl6rvGlbMt6Z+zFOgPrWLV1sGeUbDC+jsSOQ
QA+Ogw7l4xJBs/hIOF0MdIDq3Ht64IBb9Ifls5M2kCWI3d3bIww0g7xoqeI4eXVL/3v+3quz3Mwf
Pvx0/16/8rQH3RDqR31Eg4EcF5N3imaH883jgWuLEMIRFMjm0v/vTgf4VFgpDHHh591AEP6fEa0n
AbzTMVFYNbFO9cBPKT5zHGiXJZk/1vraPewy1/0kHfnGHvTYDs1wMRoqlwQrPgVPfO+OKkQ4+dkB
te0PmnktJd0eIsvOaAyQUfBrJRvoYgC2qXmMMGzSXKLRo/IUt1QBwZSrkz7drAhsuYdd9PJXnHVT
XgpWMgnaXx2LwaoZFjwe7gQdZ/Cgx9HGyEkIGbFV/AnhDiRj9qCnOHoFVk1DNsZyvGqr7CbIOxsn
utiR2pG8KOrSYlA6ACrgofDhABXd8PLNwVyGP1hjj8riWWVjwQ5f5qYpwpgzujzVE+WNSOmmyPGS
XL24Ktz8ly+lt+9XfkYheemhdhXtrv3mRP9H408gXsmxyWQ27fis/LhWBpM/CoKkEVCwJG8ZNUsj
JQvS3PdZ849A3Iqy+azf2vlx9aB/6AZol0GfGHUGs51SFBQBzIqPtJz1CIjJeOfZ2oq1aJ2rm+db
UquzLTYiCqNwsfKZ2M2O+ZlDrAemU7jnmgDl9+qZcNUK0VO79X2pJU9tpuz0VFrjj94lBdjzh5VG
JxiUFyVk2MLlwu0WwRbjrtJYwDaj10LBRrXXllo748PI1F3bA2LvHaVZ57cfFMBzreOD+jU10X7g
WFvUISQ7rAojEJT849xotilPYUAnmYR8/djAfZ8ecMkvt1H/8Es+Xj4nMdoxANtWbiXah5PoVVSi
h/0ecRLCavpQ7vbhuMvu/ahhEug++7gtRyAB8u9aFuRfEBmM0/hvvi7vv6+9TzWwKHBv2ksGdZTI
F/zmqMvIRHzxLvOaG5hZUJJDoyjmASW8RCB1PkWFVyJ2HsnkV03iKelSDi6qlxWNq0VjDn8ujHHt
qHbyaYSuadRAj6Ii9WnLFPtS5BWsDned2UYigB06phcLK5iB4C+l2KbU6VJFm+0dkQTi++OE+EeJ
tBpEZuT5nqm++mtWTxnFjgyVkNoNQqlfhUG2Pz6zv3kKwHF0RZPEmqw8u6iFwj4tE58JuS+1P27q
ebg/ZQ7UYmP13Dz/q05WPKmX07R/FyrBVDH8XnohbDqHqr9lp6SB8GDZqPK22Ltnuy5lu8BRtivF
6Uk167/m7veoHqHQvwDccuRlOGQ60BsvMkiC5ltIv8HGUNNjemIHynoa5KFC5B/vjDCfjiy1W3Fg
wgSlgkzHt3IIEBgQa4NzDO7wcg2J/rliWZLr4vSkq8k12s3W+mvPWul5hOi2D1gjZZTR2scMfn/7
levG09rZMvqplchjmcNvD761H3Ti85UmiA1ez+kHZx3EsaoBe9gnty2gfgSi269O+pkkZ6fIDRLF
v7LlVyNJ8SJiaDtEVvUOh66SBgnkgPXh9v9WQctHjLSLL+r0l7Ghg9dZFkuc0P+5PZKiyCyL+xs3
vWgMn1PR/e4F3PoY1oPOKQ5Gaf9+hepJEL5bQkl/3k+x18VM5JFJGiEAVtD+arWTkyPO+LGFpUmF
xEMH3dgFFHNvIgRNLiIWPOTYNwBdrtw+QXbC/WkZtdRfYZYvt6K6EuBlF4bQQ6etd623F7HrP0Bm
Qs/2pLwrL0iWRf9fQqBY4CWrTSRQJT3fwdsUrDTli0jQSh6Xl2uDVr2YmWCpTbfy9sL2c8zU30+c
pdInTlEpK9CrZoYuSWegEt4fQo5NtNOMUbemHbXvUa9mwVRn++KZr1D9/05LRwvgYEdcp1n8W3/q
fnzmJ3AanToADFlaiiOT3LMcBLW+DLndD+1H6bpcqZak5/QBtkjLv/roGVSJI42/pS3kkGN5LZAO
7ZIw4zfsfSgNXg8gRDx2q19pPT1XHF/u4kBqqAFXtNnEAJCjhcA2kXpJVP8fWklwATA7pMdMIx8W
2FddwvWVWTfn/ve6SZ384lTsm6s9Jyk3260fNbrEzmIBFcQOcAAVyMyXLfADEkazFMhUdezp1AaJ
7QCBzMeqFEarMHaHyBoItPVhp0+S9gZuvSUxJqtOki84qdSFMtxTxLphJ4rKcLmY7c8L/vLsxEmr
0jiG/hnMnY9+KGeOccNyePiOaIUnZhr/HLz3PO2mxHO9h+06rzOmkpkucUkMSZ7fNjtXNKqWH4QZ
v9vKqI5/X8hVqIECuU/VVgw4zSvB/kwFmsPlWKYLRtshcaBnWbE3v4AAwou+dAXRTNTaysVkkUdV
GeP6r3dSwAwmklnJlK46nixOq8gyFxiEebZ2KS4GiKoZMnvak3xW+Q5Pywf/qbVZ0dGfovG7YB32
0nJDse66hBwGv1l5k371XgDw7N7V8G3blh16s7KqW1cvWhtC9yZVJAZmXQUbrQaIL2gMsssB9UYc
sthW8zgomn6Bde5wON2hrPotQsJHocWdl9I8CZgqu50Cmmg6a8bhdulScGtbNkgL56cR9o0WWvx+
Pqrw/9OMTe2n1+F3Q+9Sgm73lPSj4T+LKcMns9LgvYHRAWydu4Rh/BxMi40AYttZw6cETkYt4gE/
ZLmIXC/WcqiKrJ7qOxnIJe45qUSV6J4o5d1acGCHYJlqhFRseAunJh5+Baa9OfAqMaKgJCeSnUUO
unYJHkma+xCuSlwOD3UiO9KyxmUAlSmzWOGRnUhZgCl1mq39PwS51BDhwBbj4cBKcq1zgosZl4tm
Mo4k0tFxF/PJWwZvWT0FiKRIqSPEHr600Pxghcuqu2RwBRIUwf6Ed8r0yizw8k7kiE/P/lLWbq/N
Jxw2d+ytxn/GfbcWryyrIC7qE7CsJ1e8escrGdYUSuzqoEvtKYSp+bt+svxOA6J6eDlf3PG9X0Cq
+uZEJKVabD6iyT7XWL9QFbxM+YbeUBNod9rx0Xo2AYuCxYXDamRxJf0vK4kB5i7vI7+6U3jATAiy
DyhYnEc0kX3gwN7HGTdGQ3dFVQNK7mCscbXnBybTr0nx2YxzjjFqvtXEOzjrbYPUV2te61Pf5LBx
SCtWK+hHztmfpeHR43pyWm9FG3z0gYaokO7O0YhXJj6NqVMspMKLm8oGM0MwlnNjNm+SJO12dwQV
Xr65tNIgP4ghIzcES4zrpFjjwI1TMz59KjvShQ9pHnDeSHEt8DUPgJW3XZfaZ3TLYZhBIgu5sYQy
oiUsTgQQMrYRa9iX8K9IMh5i6OWmDFayQc3afTJLt4o1Qbss9teYRA3ldEksAvwOjGdrVX8NbGQt
oOLYqw2Aegqt/7sxqv9ichCgAZbKkkFOao9KfFou2Hr+HztLpF/6O4dmtK+3dGEtLhujpmpw5svc
Iyl5ipq1GF4D1hVIpouqDDsl2+LeHX81aRrD5inDjwg56sKbFPsBMMW3Yf0ubFTc2sMckv+qF8qp
L03tRXmNu6ygsfoX4zx4NswRUN3tZqtmaZP7wCJOEPArAt11KMkSwU05FseeY6UVARrLKO2GNLFf
6veeKkt7Dj8EwlpYe/zcn7FwMkxbPl+KWncskT6n/XioM8xFvaOdlvaSeB5fFWn21EwbdI/Mjg69
IqjSyMv7qAwrYq+/nKS6372BEn9a3mCi9vO5vZIE7koWLP+qksPiWdpbxAgF78Ca07QMp+odcQ+5
jibbe0JdCt4TIzGAwdwZBn9QgMKUTWaWGay/o9fEbksIglV+y6ja+Zcx5gQ4I6KuK1KraYhwuac4
8tnZ258oK8rGATMlcp67seZMBZsngOhvfdHCR00Hfm1rJ7P/rNGK6NGiglln5VZPwBIS7X7g8Kwe
wbhKwUpORe0FYsa3gs4hFtlavRVErhPW2lppoEmyWx03qDKcAJu/troGLgtEmoUKGi12A5MHmVhk
wPx+LZ94PXw2LvBvbtnTru9MGXq1LF79/ewRaXTVHquMFpVl9MFOifcR7BTQGso2+UrTDoavBY3v
HsaEeXNIYTvre9KN7a3vTfW6NjbrbZwh3EJ2uqdtbF40td5aUbR26C7nnchjUcRGuGelb5R5HsZY
PeGI28+g6lJiT037ezbMekWpPLKt4Lqa9ITXic2HW/uDRCq2m9D8UIR7PAWkLhczVE0HyTRj0Sgq
UlcWisGOYR6o48l/lUak+GVEgMadaxmwE61bMbXHwLMqGtcsdW/ekXjftEyeJUYdxEqfYugEBxaB
Bblw8Xrkg+kLK+QouDrjQ9INWiAObCpLmacMzVhQ7pzBU3eLyKvjeJOX68AREGOUF30HOSDlF+Cw
FRge4F667YiC0y1gAgM4/Pyr1Jc2UG8i3r6J17Eo7P9YcHNTiR3HlBJyV7wvwwWF68Oc7old1fAL
/mVHLHLQF5avb1IvUXmrvuUmEGg1kCp7VaLImi2p085iNlU0oEfZdTDiwSXNk9LrxcggEY518lwj
9p3yKzlZaU3jY7RLyerGBEZpj7bqp8vGfQHYjgIlqcOCX8tP+WZHwhJP1+GK0NLqoAYSJI4zNbeq
NJfD2Va6pDBG1RH1doCLt6rwY7ZOQbnM4I+E0i5rN6mLq4VowTECUdX2kPJ3QQfIGDeBs2fKA/mT
UCW0FBNBWZ8posCKPztXNLcpIyricGTnQVq/JuRnCuUXrLRNUZsYjzkrLl8uFF/XH4Bini3efviC
hdUNTwxvl3sxav8yKHQZ7Md273wzQrnzBf7eDiaK4b166HLxSyMiWUCu+3xRofuwf2E8rfW41eBF
yRPN9M/tNTeQ3h7zdig2tI2RqE/dn5Ee0nVpftkj/082iMN+YNcSKbksr/IcmMwmoT+7h/8ii1Lf
KhyrgtNhlDSRHlBo/9whpwaX2vRROJ7dGJ81eSsGWiAGZE8jsDeUaP7dn0yQKhYbEd+UIDBgUqaN
KyNXeI9Mk0c2qsTNiqVAfHQcX1cAIR0vuSAbqjBlFCaxUF+LfJXFlIoEMB/0r6NLznfUJLE7wNvi
T1PFWFRVVtSOf4bBKVygb4w3p3prSpgnZ5lY/9CnVPguOJ8XCtJYZxrr5aotGddtAZV1zcw1cX66
YO1x2g1PyZfaILcyPyboRc95yrZofJfEHr702l/rkj/w8ReztgvRoPu5gzUAGDJD7XmpQXH2Sont
GS6BSSWTjsgZhjjqbKvXnGYE+24xiNuY828+uM1LCQ2WGkAVGoi8oo0p9O/l8pYRsTPMisWDBZQc
5blfKBdDec9IVCs9eoi0ZqaSpzJMz60TNrCLuyNxi6Hn3Q6ywBqcflCcYNRaLUHJHLSVjCn6CxBM
lYcVGvjs81QA7sgReipjl8EEHcLftKpwMmUYhV1KLj3I1xs6cP9P7hUGuj45G+bWAFDhfXSQdIPR
UblvAQdZelQ1u9Nm1VDibMSCaCpcI4pHifPxS0MnrTOgqJVn3gulaY09S3squmViEyU470sBDK1A
JnYJuhMcZPJmMv4zzVw99LegEZz1+oAooK7NID94Fi19oMeebYvTOL4EWGBk61NKRadeKtQDvxbD
Ifg+sSUQQZYsTaRAPgU3zT9Qspxo4TPGv4eS0Hp4G0m1gGaxbso3ZGneneK+OYmk40k/wNMbyN+a
KF372ezj8jhDiFNWMw7+8ghTvg6aNbnOCIU5Irw5Y1zxSivzUc7Fdm0ENzPB+s7MwjRZ04Mxk7Tq
McALcw/UpZs6LXZfzvWR32YnXXbuw8Kc7oXqGqfVVoleCiS7Dwd7rv69EmH3SdiXKBfEinzfEy0c
hi2tUvlBS5q2eIclpmy/HUwTmuz2G1K0wwKT2/stAc/TKQRbE+CgHRnzP5PVnGd5kQPVu3wkH3xC
IXUuY36ifOUIw2VcJAsSVY3Qs3OtdZ8TUEqCueCdBBTRsuARHWEzLNoaPHSo75cIq4YmwTKEoJGs
F6/2iNoGwIreryzExS6ZDl9yKpNm3FoTWjWrisuYZQtOxJAbhOV7+YpLyb+htdTr3r+mhpPjBlxn
0tElgN8ce8MV1nLcUpQr73+2ybmWj6GmizF4XF4BQtHs/6KnSQOf1wqq0nlLPVrHu1AnwE/+IPvJ
02F/hUJlr5wT9sKao9klxbeS2WrYwucnMUqp1bu27xUUbP8FkJlkpAwl0e7HBARNu9smPiyp2dLt
tutC8wqt4FgPaHCqIgiiPEM7DRi5QjviKZAFJfNb3/xOZKPCdpPqDC5EpgCnnIK0qz+NXpMvl3th
pFEc93oqsFUMAot33hvGdoaqSEfCTJ6OYJTTnro2ZZ6J6dxb7O3791KXJ7m9PHKghKfZ9XmSa2tN
Oi63JqPvAvA8DGUn+vux1xtap60yfIinSJvETnH2VPWnfsI2DykoHbCUATszqc858TakAeFiRr+a
PuOgx8H16UgRZgmnE5D0mRDyhYVS6XV6sHBAqFCd6NrPt6iCXSgK6y34sNib8Tp3ESed1j7sEDp0
vuGY1myHDPJbcZMZ7F5v+g1LDZUbGjGCzoMWn0NhhOJZC41ACLzBmR4HvsguJXfR4J0klr/C2YFR
+rltr0b+HaK2WVPRRbY2oGkIauH0DTBQgUxDpza2lC+iOOHCzFCab4ZKZUYn96IuDmn5nnlSMwwx
iQS0LN6AgtqfUG7K5E0fFaMSNHKMCW1rFmJYPhGLzPaga4Ymi4TQFdL5IjZXtUdDyfgKs43ck4nk
yKiZKawPoMoZeUmOAExkKJWxh7XhcID2IFKZAHlhL0cv2oWSWVa99AKe0qOEY/6JEwPpvw5q9DZW
x3IGdhUEVsjjZmaIvQ7xeLgcH0g/DwQ6ll2hTWaRpJ0TA5bq/mKs+8NwdpLy3b/AOCA/tSD04WhT
8txw6kqRrRFohi8ENBRfz3pDEUkL//10G/6vJXIN5j5R21AiEEGwDrTq8p7C7H3rJUnBNW4vzPfp
FeR6GD6tx6TMcYYLLMPKPBxzXlKC2fKUncK55CcwZVtf5+G1MRDP1um8neqBhW9of9oSSiAL+2BH
9U1FCM20wS68Xd2S648s5OQR8EGl8AM6Oz5BgLNerebYoeKE81fTkn1pcxSyzVVbb54y3hC9wHIr
6Bmr0JKz0qi644aBDNvjSo+vzLYNScpblApivPpxYZqbMP1OiPxk/od7fVYkkmcqCT/utR8Kntog
hJJ013vQgOsz7drD7WggMwNANr9cTOJNUkWWp+CRageZjI1Mx5B5sn0YjpxUfjF+TucEqMTdevEU
qmt51iZRxAqlXYKIxAw25AAe6+szd9vN3XESP80DjLOCN+O0iEh9nSM/i5tg7lLA7v09QB9mGz2q
peI5Tc7AZvYYUGI1/m11dnzU4x4UWxBuJm2vNqkKcOo0Bb4gd/MWR7bjPFttCQ3/sPkhm7hwIvTE
J0wt17aVJcSLmTW80/Xz+vrI6McX4C0a5qru4dFMB8p7cZ1MwlVWJ2gNAj5QutXR0chZIJ2y/Pfh
4sjvUOXX3WsTZkLu9xKcQvOhQxZu6SeEog2XE7SMWa9Gzbf+KRIgKrDuz/YQ/0S/xrctufQMPfSh
pOiJ40+saIwpuKFF9M17r3Niv/lpqTwYWpGM5xIRttngT0PfgF4XJeK2dYhOdDbF0zNCWOvxR+ta
4I65jsbp8Sg6q4IrX+6//novt2yFRdYC0KcxgPSOJa//p2jUqt7CZjw1qmwoK/T2cb4qrHPILV8j
pfEnOjrS1IhxqE7kir4jy8D6U2epItQP1LKcFCaBtNGEQ2eBbjKlSGqjhTOjhgU9vOQZxAhK7hu9
ZUOFHLcIP+HxCMH6jAgm9QCjHSRyEbLczJ8ZGOVIxmxgtOa65jSPd4GNOuIvAQMdCG4BawMf0s2z
Ff9/Dy+WCY2EaxadxT3Tg7mnMmMuIc0B9Nn2/ioxPzduxDykeUgNLBAr9ASMyOD0fBAOlI5zbQ9h
ytJB4LXvukshGzEB8Q5kHjeJpwxCjTUpEol6FiAaLZRcZrok2AZe0+7+BjTC2HL+ZO3257AyAz+R
O7/8IFShqkh2tD9ViHZVDPp1LqmDRwC1UpVPWxI0HNbVkBwqyGTc+B0S6DMCyhOeKBldxbtKTtR8
Bn7+I9kjKjC9Vu21xz0d/ajLjRm9LdYsk8QC+pndTilZ+zNVL2rliNZ1PM9cU81YbJalbK4j+8ih
BBo6hLmU3cY2vZBU/CYFc2YtUYFKZTUB6AHJBW6HpSwerAZUJ8VJrYMCDPtVfaH6X5dBHbxHMkPv
PrKfInb7TNRpd6hNS1gnEv7reeUzUy0Qvv0NlmqI/zuLISD3sJCWFAuLKHt0JeInFE9On44v41/3
ZjDwlM4NQf0vX2Du59MMUj7hrIQoRYZC8KpiPIZpsUzQJmJXSNr3M5Mm6llf/Zh+t22q1Q1VuiOK
pTeeAAQ0zVZSfXv+sKED6NI63BmF46cX+3RceaNW+dOhJaGhPeyUTSPQ1r626TdWujb468m6pFlu
YqKMFfkffdIa2yJZEgSrr7HZ1klky9mHhwkJE6S8J9aElkRCa1UOOSLZ7vUY5k/uZcOMcG9qALqn
bFKApvjCsgQDG7WjrwAablCkGLWaTYgcqNLHgI6no71j4IiwR0uRh85k+tGVSnRIzA2QAb3T8Xze
/8rmjqzGkSosmHp+Z3JpOh+dqpcfJj55zzNHwLU1XCEmokGY2OGbhKQ/7vyAWpFnMzu00yp5d/nU
xYVXwvq3KA80DlZaSf1eGxeyfp2igyHnlRal6NL3vQZc4H1/EDmValhGsl39JBOvh/iU3B6adcoh
b6eh7M+f5IxGXDqxgKCe0nKVtzD1QTyLs9fdidjUmPahox81iKKJwNjkT5X6L7+aL1OlWcNovRpV
PK1HJwK+gqA4UPrcnVBIMJb4m6adiGS55Pvd6uv09zml11fx2Uk7pQHK+Z6AXbznjQK5o1NCjgJO
8dllfO9sOIBxfTCy7Bhyzr2KHdcFqLEaRKd6x071qSiMZ0As4KJ4YpzLnt8YPHzDu1WRJrpu7GTL
Wre2UOBMXwuRpgMZbxWzAeJEHrxXGnrbUDnZUtXkcHI7jRBmMdejzk06DSxNoADW+S75CrIE/evl
DWMjGP3wkNbMTUSS0Wj0HLpdUAAw4RWLudLh7Gpf0atFROZPzN+3z1pog7LdNqkfBxFOtZEZYQIm
pJnOxzk+V4ld2CnkbBwNUX8sX/49eEVeHZoHFAy0Dut4QW1zLBbqdk3xYsbLHURHlQPEYgctJ5jb
uvEBx6jwxjALrCoZQWSC7FxZhbx8er+vCasEMry7uoQLz08UNOq5BYpQ/EdJw/7+rQfT3bfxBWhZ
t8SIQsiOkIZqRUx7NZseNGUdQVl8zia6Fk5uvUPTcTVuoHDDlEJtA8bdJMYq2LzSKRdNbL9YOaz0
5T2/ygHf9hatN3mbdPoudXX7G8/nV8ru6g6PHZ8FcCZKoJZYppPh5a6/iecfjuVX6v22NPWrltQE
INgOx72TZwE0BA1znLRz4IkjiZ713AudEoxdKmKjNdACuuO9Xo0NrrgDKrRlo/cMbFv0wrKxBgKc
/jpCGm2dC4kaavslAh+BYvv0B3YUx3a1IXBfXlBPPWhPh/6r2PLTbA88jELfX3BSdp3d3LGhsPSu
Rrh2tODLUeXy3FDteSBg49SKQmsr57fgLd1nX6gXubh6T3JYP4uYDjw7wj3oKb35YelOl/JNsErl
Wwyc8rnwqC1efdJjCse1yw/Jw9zJFnIlYsH2+dMF2PpxbjWE0wlSwdPjRnN9DgOnQrrlLW6YVfPH
yeelwJOD6TVkXvPk4SDoz2zSf/PCwjvtcYu67LsTS5jpM7GfWeIw94PW7VNhsObAj5V+knlqBZiR
2cKZ+oXEwbgEwaUogSYitNkws1JwLtiPjKhztK4qrAWhzt0yy75RvlV1U/A0trHQtqSlctJ5PQGN
5RXroXyIbka9fyCZOEv+uz2PAJANqIFzZ/BGGd5+uq8CRgFmVmPVqaI6jWZx6GRePk9M9MfS3EHi
zCFJT21Palb4OvminAwf3NFL5AuQhJqiGEaGujlLjd8I9JIWHqstjBGAb0RmwcGybQlBCuDSEr6e
8xeaR9enchdp7OOsg1O7hxSr94d4qHY58U9p4OCPKM4SArcxE2tIVFhi2n7YhRZTQMjSYj6agclX
ZcjwvcQWAsY8RBYC0UROPnVtMtcaw147RqCi8G10HZHtKPsUBHe/O1SdVuGuRETdiUI66Y8iUUGU
VvM12BDjSY1KO2A8CFG2eDl0RhzaKMNPCaEDIBR4BSpxTlpLc5PfexULS2LyNDYjB1mLKNbcgITY
fz/gCGqu07l9Uef7lKgVvzEHy98ue1BeHL4IKPL+BL7/9iCjC8wvS+7N/FG2lLZOzMr1sH262Eqn
oqU8sE7seg+/G9pur904XNQzjc1lvbShc41KV/gcAjvsvWBS8KZjKJ8R0RK3gbQ9rf1qAiny0Vhp
a0JOK69/KqT4jBzSwoa/TwZlHQLyG+UZmMbgROgiw0RSgfpFxgFlBWTi6tfd/cPKWTIvoVFx5cNR
XIMUc2+MyMNkOsT9If7iEf14GUYvGRflheTRQ3YzqbiAC+Ik+WjaRI5g0yGm54NJkud/bhE6mzjg
gCmgO8azHkI0S7kid7sj+RIXJjYscVmHINXQTKRgd/lTHCx7jbb0GIrjFFjuhZwRNwbWGJPFhfBi
Qmik560rYM8OQVpVDWwVfuz6nX9YKkVdnccnDY1I6ooW5iuRGjuBPpr/JUDDJCIrFQf4wYqi02DU
2TaPDaCVEqLD7GCQ1Qnd7K0f5opeIUUa1mG2QSHMtOLfGu8id8/kVYShA1XDt1Dnf0MVPdH62Cxf
2eD3dDTpSCZu8Yhmx6nqIjOh7Ya4ae4fQxVw70uhh6bnRYci/Ry9SnjBanEMzlqQRFDBWdLjsBgI
MC68WDNQDcq2KcFpErJD3OeXegXl5Syf4vcBngIuZHXGnfYxPMFFjtf8q7sGIUNE4NMqoLbQ1+nF
TrG7UVNguDPogwbBe5J0x4nyPOEGpx7DajQQOz0ATbJd9tM4YjwvMVklfg5EEqlf+RNnVXhY5VBd
ZQKcfu8twGyn6UwgLVv33KwD73hGuYeTCXaDtEBduFC3yEJTSEet41ldtAVxyEOYgFzcKMAvPK+X
qbcMlo/xidlNIVsE28phWEqOZDDu4oyHoYMKViTfGn9in2GU8PT0WvGVQWWcJ2o2gMuXENTGXWRJ
g7flumw/Qoj2YRGObJMilONd8eWDdFlPCG1V42kk3DUbCO486GsF2VdzxANAtoCRGeeT0Y1rnM/7
R/8tkg5HlKhOwlxRSjlerBqXlbicOrlBwxJbeLMtISmlFjXpF+1B48V5O7PBZtrY7HyF5Zhd6VeI
2YV+DMmncZ4R/Rfdoys7ONPedS3Eb52mlSc6TyfxBslQNiYhEBa3eWc7XWPTizi0HAWMkYPItngo
Tv80TzLdPgkHUFLveqfqcPHD5Hdb78fiCVyiliLYSTPCYQEtWdqHarYyotD71kS21/QJREN4eW85
VWEUdgq0h29hUaCxZhdQCn3z8StMdnz7h5bUvybrX5Np0Tbj9x1+7kXQHwhzboTt+Sh0qleoGjcL
7u5hFR6zP7YN52ND2gQZ+G1YZnPnW5YcG4ZVKamjfAqJpf14Hr7mXgR9cXuxctz0osFWDfgkZTrm
QIlrFZT0NxFy8V3SEb3x5O8w+sgKHl+BLRyMQfvnqeIv5k1uPnToss7lq3v0+vNkzp+URcqD4DIn
+5IC4yeJgFda8cJY2nO1Ffoynk/lIr8V98dJ1n6y0F0oIVbYqKMPSZVFEoxiq9q1mDGDd8GnQowe
DoGxBTj6r/M/zJYU6yz9X5sIhaSJtEsz9jX2qfmS2XIRsLPKWqLgvEfgAqwzWXTjJNqFfz8cq/lb
LAdJzlMe4xcdbgB+lFWimIkxop4Vnc2V7dfzMQr/JPAys6i2duaPyKZCdyXy0yiQF8+rjOG6SpkV
ruG1F0N0NGWmcU69XCvUGPeFcTSoFi82xFFYt+P0VQv0aO7LzxKNi78AbuQPv7FISBtXFVAD2fE7
vecOv6oaLmJ73V2taEnpNIJzDxW3FgpeFNiZhwuWvHoOW0xfgQx9Kdic93eQ57SPDFRFm58Entjj
Ul2ny7DRQmDZONTCwSyt6wSISggoWIfotnl8jsyOw6gQobUYB6MrxaW0/jgH9vvsvqE/yu6sIHLX
qAQHbBbK9VJeNnrbvqvp8Xp0I5jt923Q67XysG0Op9NkqjMvcv0ZPJL0vW0j6TlVzu5/WLDHCRYS
o8eZkiloyyGJG6EkgoTlE9PYD0AE3CQ+N7Q8K22YfIRop2ijueTfkA8RQRCHeobq2z82G1ZYnI+q
ddupWd7PxFi4Elg++iZ/0hfrSwhzEcLYo3IRY48Q75Nroh0yCaT0GNH/NNBnSxuYvc+pa3g5LXZh
Nn309iSUcwgI69Pm1/wEs2LTEOPVDYgiN/rRptq45CK4lLawXvonpu+atL3d77a+8+I7q02EKNg7
u3I8+DZAHJkizQ1WbcL2N1bNU/AvXeoXYO0kBH2PGdJU3SUBF9Fawi77FMbnEGO5Qfb1UXaPTjvv
AC5GkRR2hFJUnOlMSzpRdQp7Jzac2pVyzd0DUcIgCVIzrK1X9C7434KeJ7Lbev0q4gwfKq6arpy+
L86aaFmvaLIVY6fmJtdqk317Y9Fsv3ONagkUEROTGFvpoEbztFbLFfRFEyx5BM4Ntj7kZUEGnfd2
fcL8S9agHQVbvVvalpRb6e8HFtCkH8jHNZmhlS5cEVMy7973+4vbnP4qVrRwfvmn3Kuis1RGUI1W
f1A/KOPschb/9OvMaxrPfNOV2w2wdmL+xjV/ghH74X+hnaPQEWKUh6ylSuagkYbRk0ctnqZsm4GA
LKXiV+Ys2HTwP89pJGQjffMNpuyH7a+B7LtKqSZs1veae0VXdPuRALcO9gGekEmtWh7YHK5aJuOj
ujTLZD56qb/6icMaz7ThED8lhjWfKeL1xwBpvOSOPdSMiUaBSBUodIEM6Igu6uJoG0VKdkRVyM8q
5A3IE/qEVkLucudhfAWDT4NMSv6aENG4zrHBOZ2+CbdhsvlIAanObaEot6mBy3nttLCoIFkB+bBK
M67PfNUBDJkhe8VgZD9OqUJIgB8DB/eKPknNQ8kwO/s8Eaon+Srh1SJjDPqh46Qb/lTxpNN7zZx2
a7k3SOdsypBCGX1FE9lRymsmJmbNkGWHyG+nIg9ZBZOpFw+aTP83dCcBCuIh4lGJi/jlpj3rt3ZR
NpgPaXMLCZ0Q4sk7MOtgoWpsz2fqIJ1zj5tQJ8F23eCmaFL6vuJrfaUE4p4JsaEinfWhEyHcPXvU
eKzxWG16Ir+Xl400W3JPsOI4M/lyGI4lMfF9bCczdkJZqXOq4OXOoGS0ztpQ+c5Qva9mp02vDXib
yOJ1LcmTB9yfzNDKS+SyP6bdcXosgRXQQUivGW9wIHV0LZFJ1r+YBEiQHg32QDHXRZBxW5aQ230s
DY4EBTPcptcvY7gilGVBGrB7dXIH1G8uDE+3R6bitq29rGT4nfBfuThjLqw+YMLshEjpxXldWJeA
Jh8LHs62emGiRd1Sf2Zi4XvGJvuv1pGiaksFV4Lg6TF/9+iqetptk3/zqDmnp2+PQL6EWLeMK4+D
sljl/p/uvS3JuuyIGmNXEo6pfLomK+Nkmy+7gMn0GQU96a+JQo3Fen9G2hVGLigoZTmNvBtSn4Bi
PKVzYguASLo8HWRUblsfRywEqG5WPN6hzX2vWHkw7/I601cS9aOT9Km/qpH2+hy1q/kDEmVUAxzs
JG6y/5Ua/oyTTdrZA2Ku+jjW4Ralf4zzVHbmf8PoF55AAU2Bh7ZLAp9l5me8eA9gampNJWvDpFNj
WWmXnyQ1trNjZ72TS/HSc97qhmn4z1VWg0MzMx0hXKoZkmqD3mvgUzg526F/FgGMDoFXOsG9fRi7
RZ8kIEsmFXOI07XOVk4S+5Al3vApt2JvcCOzv6a5UAhy5Qyb4H6T3EFbhZlQi7g4DOZ6IJM/J1nL
ez9DmTQA4zw5Zb/+78mkeTH4NaSJ9ixUbqGigRL058A+hc6dFifz4y7wKrU9DXGeu/QAzaZ1QM/p
36lZi4WhKLE7P3MwEtZ2QVXSEJ+iKx28qTArrIB6G0Xxske/wa07+sZ0uzyIeOxSCW3EO+WH3Y3U
d2SRdo6CHm8CBLmY2hFnU+NHsEsNgj2zgGbeF2XVsjCALNSMDncfBX/RsOQh8q/xDfs/gDQtunQP
371lgDP6gqdRimG0zuNupALteeAxcXcC14dqrTHvFqUQOG4+ELelKQrZVym84jbUZ66R/9bQHMso
0HtjrCid/Tk5xUQI+NoR5aw4qW13hcObjGiRG0nzN1T4P1fcuLcme+4nybStvZYDSfdlpV++dhaP
/ZC8nblHlKr3gx1Bi9fmi7cqtgVhyoiRqLMLgrBDQb8MznOE8iZuW4t17lFJwcKaaAJAn6YPkCbd
+Xqn7ZC4+KtHfJR7eP3XS+rBqtShcrsrjsltBRsbZ2vUBulF8cZaybHOmn7pr2G4S8JD49CvtwQB
sFWMkajcAiR29HSiQmumlNS9qYI6femoww6V8Ry6hTH+MWM80XskWVUd4/PEA8pnH+nTbpaVSrsb
knI962nbm8WznMgEu8lDkpWb4xIzxm8HN553oo/yWKtqLQwY+ErQ37VrXlMEgF/VKQA6OcqGDnms
edhJcBGj55ugSFFjy0tVmMevb4xdbvpS9RFH7wd40A9ifJmGmi/d0BEVnMIOAPTNkpm1idTGt4sF
Mq5wMCtvvbAUWi+2oT+3+2qoIN9Gal401LxUmhJkUOUMgQoQMKQtiRYV1D7Jj75pSMPr56a1S3Fz
Uu+cKXLDdYb3w6EERwwADCi2KSTXOOiuwpcf+Jh1vp0iHWgfc2EcyopkjIKvR8edH1Mp/ksGaWQX
KO2BpEhUGkGl/Y9//IpB3trGh8CvNgMZ3O9MfdDMPxKHi7Qqf89mo1/CS34apjUKeAt0dRmI+H2+
AzuKQMVJA7DLfCF5Tu6z7NyDC5b+qqMFbxychvHNYxPFYKdrnCum+8lNUXPhdsYUPrRwXX9O6LOA
+sJVGynicduUE4wWFm1x2bwPMC9hM8FKiKk+aEfAGIK/TEB10esdydsZ8bpm7iH317m1VtekiXbB
cdVk1WP3NIZiUBnO5jyXkuzCi1O7QaOpMFXUOaEza1oa1IIHEbSEoVQwtqJwcZzbVlAAPQUG7mA2
g4zcCDq8VcUaDWY8jlHsOzrFEC2KoVTIOBGycXJ2XcBOzyyN+9Ro4X0/RUhzYoFRU6OQsJI6B2CN
t3qopPEEAs2jpWnTh9/AliXXzKTTkhs3ECYjWP29uQpeguAF+mkGLESdH9xRdXbmf2DZu/1g+ySW
/4zuItdRBi3+8UP0fmHpl9760dV/nyX9oJwmL68z3yjBfylEr3ua7FeTp2W5nAmuFpTFJf7heNgN
0vrIodXT6MlgiiMTLW6V6hJAN9xlfWzpAqqWLs87F23tSjUrAv/0nDOsjPYGtNBPCivrSRWvfQjS
ECHl7y+9rE8G/TCq5snfzVC2LYbPbWcx1mBcg6a9K8kNYC8cqR+gfSp+OiKGlRiqm/gn40VBLhvg
f5ViX0L7lixQGr3XV/99rQtXNkN00r5oJQNMrdSiOutqXDH6P1/i60Mj3TJluCJPp2LjhrSjZwJo
9wzZKBGu5txmJ2tNke7PC7zNWU7VK5P6kaooj+B4XWGd0oZv+VK4VNEOBKPFv/QQNUWlSudESDVb
re1g/LjeegIdZBq1+Ot5Q4ll1LEL0pvCUmC50OcClSgUYWGmsWMqOSrfnEhN7MS+qhBiAyEiM60e
46WrjrKyEC1lIBm0OH3T1k9sVG8hSRAZ4wyTHq6lpf0alTBgZCN29cdzvi6ul5rfSVbWugryofIf
865RDNhxSmLmlXQY3Hi80fxDAGYnlfYM0A5tWXpeTypHusMdB/GhxdIGCwldO8O6jsMRgIj3nwIg
sVvFPT+0+b5bHya+2inGM9ulJf+m5AcjFxkAlx1bhDssTa0Nz1iv6PBZLcACmKnjb9zhjGL0T3j8
eFbBfhOOeyDzd2oSAPbEzIL8M3QhD391mMVmSjbqAB1xPwaxO0+uTQavh5sLXn0Nc7wABIKJzqYG
HKgpZzcs+Z0JcBgyd6G/rxWpXpmp9I4qm0LjaIUrhg0SifyD1ZB13cciLLwijc5jekdfDO9hh//Y
PNDBm7L0ufQuDXnTHUzJmQUt89CAeyYMMnokOsg/lULMu4yV51mE47o+8aU1JsmdT18jDveFXdlr
2g2oTNYFAINMHQQuB/CFcIbm36yZsnz6HONiPuG3cOWrvyP4gWCkk/xUDt22wQXYsoyXC1ThBmyx
7tlDxMPdYnNay2S8/TFMl4QNKF41OHtjWFSlHv0GGATgY1sIHQYJcNxnbPFZJssuCLOs8JVlHwrA
DQhIynp3VUbitgkvngnN0pJbQDKAf2kv19XfQvuGQ6hP4IXmsFQPmWRe8DfARGfLNYjXK5hSgZEQ
THoMVwfTzPfZ3+dR2YDi7NTo3tIqN/ddw2IL1hDD9ErREs01AodxWAWZ5j070srq9lVWZc/8hZsX
hZYHhvg3b37/LYDcvZK1Qf4CWiHmF1GPIV8V8qVMQjB2niaViE5lwBkeN8Jvb+PXQeolXw1IbXYh
CpSV79Vy98p+3uq0fU6aJSvgL8Untlqr6a3FOP9f7NUxyjamnQSeDe9gtYltX5deRN/QWJ8sz4cP
YD2M8aJF6xRnhwtv8Q6e4bJHfFx6Qi4AWk9lZbIzGI3nsxcx/2fzjeINCazS8PDSnTpKOCdFCRqG
83GRNHfDtEl3kxTjZ/lQUToiiG7jn1HfrtoyymRmXQAgSNX64UkmL+OoSiDubTnbr25AAGwEUbem
jMubpxFHeDtTgkznxkYFbuURQj/5WD6A1xrXjXAX9Ie2gcyshJwG0i8zcqAFj5Zzk0yuibyjNKVH
7URrN/IFja8rOLbBxP/GN0ilcXhcQOdOc4+DZ2W3g2kgnwRyBCjbDbr6pQ9f8TaB/AVcP+K3oEnA
RZSp4WR20JMEnOzaTnvawIchSVThURRazeJ03EjwAKsntDZIxkwpBrICI2b4xsn0adgJeY6iS4jD
GvqTgDsjB4uZY4OBzv5U0b8lVvBv4Gn0uWr0gZyTOwRtMkXxHaxvyInbFrUTTcnsIMAA1o6GrrFc
ZlyexFFBGeitSN/NEgcFnQty6eu54fsK10MaM5jwfUeGSbTwt0IhW1Zj6U9DC+8UWIPAoeyuEQCs
MyZBfc6845WqKeZC5lrpJdxosSihHifguBE33AzvqIE1892ts80uiRGZNtaROocINfM0Qf1HfxP9
oZeL1IMli6LLnCu3ON4eN2CF78TFgQiklb487HrY1Zggymd2snwXYLNv6nqBh7O+smqNozCDNlT8
Grjv0/D85OuLAz4Nw4Vf+vorZbgW7073wkMkcyLVRJ4w4SlLyzQiSZBW1c2BbApgCA0GF8UyZFSh
UNkbsUTvSNBiJtBCPULs+vUTFqprkVd9ZcOt0QoiRyIQ7va8ClwjFc5Z6t2Qf/yetrUp7RwJ7t12
tQFw4DUlqcWjTft6oxGPK/HWlAWQEoF/hEj8YG+FvFyiP8g4g7rWoSYfkS3qr0+x3Gmd87Xb7n8G
IZjKE0YuAT+o8mskV1iErBslhrABl1yky/I0eMfKAi4qztTKBKriigDnocYkczI+TaJtE3vFMZAZ
2pka6pe0WVfhM63N78Vy4eGx8BbJsHsCFp+CtVIYJRpWEyAHLi8aA2FXdLgLdu4kV7A1Z9oK8Ixk
26xKNAz0iyZTTVOpSetEi3Gp2pSVWDbx2LlLS9b4Gf1SduhDAgT/WTRI6VJFJTCR/fK+4RGiYEKQ
0yC09n2+1giaezzYTtj/kc6hNmrcwQoMU1zAaL2YP7FkWZfvYVhBe3SJXNNd5oTefdlG0kIXUEj2
+51SaDKXqtH0iF5A7GaPc7+baZOzPep63NElJ1V4k3TUoLflVgch1+iusbORg4JwIBHizRnjVlG0
dokkwwKekfCT4AqVBETo6nukw32Ri+Dm4IJndrgmqLsXgSoGjW+XD94sywWzKLZNp9svfmSKHcZA
Njq0tDhglQjR85RzmfvSZJIleeZRNclHq/pm/NTEv9JExhfhXiifQ74ieaYml/+saemdH+o1/YUV
TC3By98FqMaWcjsvwqAwbvCU116+n0EzfNNEBpWhANugt8FtS84TBvo9oesL90el5nqxfAGIAuVP
wA0GG57Fu9k+m1MpAoskSWD551yDOKWyJuggBSzSSsCAGME1RUeFvTOAJGYtKiVaznwiM+ctit7D
FXG/06rbLgtb10DaHR2AzvahBairmEsmam45kQMFn8/JriH5MlSwa3Hs3BKw5Xei7EtFG3Bkix0H
W3BHbuZrKr/hbLwI6GifJeRH7EQbq4lrho3onFSztsqq1G73Co5YSWnW4XYbyP2EvBsg2azixbt8
Y/ybh/+BL63+ODEx3tnc1IsIAK8mgNawoiUtcCvPwA7ujXsr/taoGxuSs9Nu7YlrkKrKtOIoiFpr
90Uct230BUp2z0Jj9KskDpSx+DGcHfxXpE6FWR5EcGh+WAG04ykKi9pBfS4ysKx2NxJYdQWKaObU
sr3+VbWTv9hr3qptQo2yehwiwFrDNCAax+YRjZIgWS3v9biq5FBKJIIZ09BrjGmeBOwMLvmu1Ahm
Gdd0kgs4HFbciMn9eoYdZrh74gl0nH6QdQDa3NATZFf67hhwtjZ4W3bLcV0AX3ul9QZE1mGrZfhi
pnJHgbMY5s3S8Gqjkpx/9tAOTGooZXB3mIqugPCVxwaIAplvQhBrICyA8tOLqbGqoNwTNUEmuTA7
+9k5Ju1mDHf1Yg/wTvAt5BUj7LjD1G9l36b93NlV2Gqc35FR1/tUBpfy1s1T2v+cGwbIHIJVbwAC
B6URva2ouZjjjR6sqUL/OUhB2NA8bOzHlb3gjAgsEA9gPjfwAtqulNEWy+ahAZnb4fOTGUYKPIvb
UOPy+YeCwdyk4dFEpdN4UYrSx2H1pxzBFl8VdyzVxcOrG5n0fNwDtQRYaIKn9T5V/5uhbHje0blu
YHeTcAvmFigNv5HkN1EtUdYigntA5fYCiocxEClJ8P4R8o355dWCI+Muftfbd+A1TKm8qRNFAogg
OtPa5fupPkkXQTlvWnyqOAZMHvBleVoZFIaIVfxvgoi4W8zg+E0CNBFPTM+6ePUCRFpATFnJ9aoC
4n9j66bmkGN7C8TRTG7+yHBGdyW5hzj6MZs0VnizFFWiX3L7BNLm2zZZsf2peNWA4IBOrSwdBSoK
hMFUcJZTVh8AbiRfA+0PCH/6FBUVYde5eI0Fc6/UcFWyvzlVMPEs8hiJcr02NBEHIcYnYvAwnQJl
bMjHIVy08mALUvTjRc6m9d88t2aVxID6MW7O9SCfIi1Nz0TxJhYJnCYhHML4a7NGhAGxC5WvFFo3
q5hwF/7QAe1aVPawQ2coHognpDblO8IjIFXqIeeJ0U8OIkQnqw+mcerqRfU6koaYIGiRJS3GV8sq
dE3WXkxcoafKAZQjXRDGWIj2XlI/JUHPqvyij8E2o3HNFtMCaNrpEVoIbA4xSxMLH3a3Fv9Z7dPp
3DhPEy/npOloDXpiA+bvmKWIya/4JVFwzjFSrYZiEj+R/SHKOmXL/AN0bGzoskqqVTK2Ys897BQY
dT+14n2DmmRyE3+eHy/bh0yITY4LeTWMOiOM0hpi3pBBG23g24L8kx01S+uXb2fmJ8hoNcRD3q4j
Oyq5PVh7Ms6APsQ2UmUQh0eAPfnln1Faieh2HlLHUz4fjLhp6zi6t43xiy8kb/VgbzAT01A7rfpb
5XnNMXimK76S5UFeRvBGctBJ2KU4rx5RNBSVdXH1yE+yw/LUFdHqcPBLzfeZgvUAwuTTeZtOptSz
LRI42bRnvKxV+xYS1hMRyu8TA0KMBA4aCzSMR3ojYPF9fiDShDsO+EaekmvRIeuHBx1Beoz5Qe4+
ae+VTUFpBxD6LuzT6AnSCqKjBKPrThXcsIXD4Y5i8+8ttSz/sVXVa/lfmXin7iQ5PF/xcICQ6x+W
UBfN6oRxzcgYRz5tRpiXBo586cKOHb5jGjadssbYtG2AATJYB3aax9cK264QFdQLEavQSmkHzZe/
/H1HCQ8fS665OGgotNfw4RMqeJUAPofkpW7w3C3+QorUftokQLI9rxji0IMFz8G4nbCtP2ikahRD
nXH8IG/Ij4ZMWU0tP5JyTnsv7c5MiGMie2RrEWoXbMGfkUuAGtb0i5R8eqwzGx7X86q9RHlQadIf
HF47hIiNh+RTQAeYoDGc6uLVuWWu/JaWQbjcIwy2SlyQOLrTeEsitrA874cYjoDJiWhIJ8tBocSO
aMeyKOlyVP7X4KrO58OZec3T3QuPijpWzTmSGuYuLPjmK23Ua5knokqmi/EhSh4eT7nWuUwQzOYm
zw2b8iAeq0DzvqzhG0CuhKZPb1ZXbey5k5etTNOpEB0v+YJqWi3LfaQKLPF16rZcYRcWCd04Ytiy
9iPmz3d00PSJm0dm1mUjmVNbTN6pC/RScoMHKJ5XDrexmJyl9S+KmAgFwi87ZCBILbtbJK0ZxfPl
TJV3lh0uR7V+8G/lTjxu4OBPUd0W10M0YMqg29k3Y4YLR32H9EhQQDUP8ZuFM2Md2Nll73yWarbU
C5GPlQZWdNgYXf1/69S8e/jcLgke2CxZJZf799rdgrEJTFpZ0g/tgoBHpFrS9OCUdKAWbsA42HmE
WpxcFI6aQ5y33PFED57VvVdn+CL40EiFyxySEu1Vbn8hmHdF9vGKRhUCXl757HQziq5h4z8JuTkq
3wbm2kpXTKZGkW+7qfZRg5wxyU9Yc3zhIlvWyJzrNU+vCo25U1mge3fOFid+Gx6MVNNhvXh/B8xq
lVKQ8uyatX/L5EXHjL/eUYmEYHqrTk0Cn8T5JJAC9SjcB3PwwebTIqL+Qa7YTCkfdgdKGskyw6fz
W5sLjg+iYAtb3Lm64jU/dZyrCowdGDUGSmpe0j9TX8GBHPjzXUfyocAA8r6LqQBFnWf2RTcUNG1X
j4BCTbBQbwZzP/gSL/MzHoz8o1HwjE6VSQ6e2OBIohVcP0vNKlJHF6aOGd7Kq4rN9o/a7wYvawi/
K9W8aEPmcllud53zG0y0AUijVNNN1MV8LOiL/tRYM0MnNQvVmZdb5TVe8kzbylKxfPKUk0Zt80ZN
d1PPg6MSKUAULjgWIGHA1uoHOJ14jTk99HsOxwnDfnwlWi2Ak+5ORqS6MIeEqpgqI8S7lxQLukiS
5UzX5ttUPgacAoOeOJfZLxYmbvn2K3Y4CrVLPeg9nJElggEiuL6GMfSAtgU8UzSc0UHp/9k6ecdb
i2XJ1kXDf011miUdKwhM2/T1WpTXc+hwL/ndd3Jxx1HoZnMVYNOuWwW9gkkdzbde2PceLeRIDurn
pAvPh6rBo3V/09bnJEaf+sepvc6xY1hJMfpJVWo/X00mZM687bbrAPapvnmjt/OzL139zJNi7yX2
R7dOrLChGqWDpxN7NiR/Ylm+S+QXl1Po4dtfJSDBsPD5/AgKBW3LYJoj1bR4xQzsuwwGFm3RJ2GA
xlYQMsvMS9qIR8A/rz/t1GNiZ4U97gklnDGq3FosfWQIeavqVNAbvxVC0dq0zlh1o/K2WnvRgmCL
Xc8OiRo/ZmZaVh0Tp3naJeBV2AUGMtctKQl9v0gref+ghps+ngvSZIhQnpkTQN2P86lCcQMo80j3
v7ukljXL3AbRUcdfQHvTJ9BpEWZkUuPAsbYfjrzzu+Mm4d8pgWGdHRhkrUn+0Vza8dqaIx6QlFPM
atfEGqgCu3uaXFoTOyLWcJLkm7oi6yrjgLz9nUNafJcTgWINZK9XM4zMygi0GPywiclKIG5NBWjh
jIYVujx/WLKm5GtnLLJN0IK5A6eu5/zBHXGignxlQj7qO8GkinT89D3INdwsxR2eZ+PdzDQetvt7
wKjAm0cE+2n4y18SCpwdoAQCTSyoxh66Oz/tloBagUa8fyNzFf5J1lwaMORJ/RlOJrZvYS0Z/s6n
rByrgDJn/sHarxgHO2QQ7j/YlzEk+wcGASqhT5NCkDAZRYuTJSYAl8PhAATamu1vIani9RorhOMt
EH7V5iCiYFNQhQjvbV5dceMpiKXchvdY+wTb6Nt5bUk4KV/Qm1cl/vVG+Soyco37Bj1Cb7RI4a2n
vAB9jU0WSC49/ErwaJDGIaJ943QE0FQzgQ/F3v0NZfVZwazI8gO+Kqf3frqHR8zNbGu+HYnCngMd
e/qXF0O7m6Zwjnw90gcIiiYpodwvXJ3MMF0ODV8NBEva9CPmXuYCY3Fc8tStxBGVvjMNhBjlDORC
ePA/eAScViQyoZPQf8bNHaPu76FwjZoyBkcOxdePalpkOeLoJMoLQDw8Oa2Pq1LF61GyzT9oRVV+
N3SvG3OqYS/7+3c20X/cHMvqDVVDmU6HEjzHj5S9QjBD3oGZV6xYu1yHm8OuWnONm8+qkDLQQAdu
EYdzkB6zd7v9ej4aKErP2cPkG6ANQy7x5aE9DMHsTmryZL81Ew6lWnHC34I41ZrEBIQb/LTWv4+c
jCD/JO/TN3YpJGq9pbeY00XU7L5NPkcExnit0iwT0ZRYWCdCVa40e3vKTPw2pBmcKowAjQuJcuM1
e3XUGTqOycoiDPjO5gAEWPhWXwGrfuj5jfwJBSBx7MmzFIWBa1iyT0xsrAhi90kIkod2ChcQJXOv
xf7dZb3x97N68ZQZ2mM9LQqcdBfKp2dYURx73/lY87ySXxN19TmqJSLZD2bt4D5RJLA3uJ+baYJ6
2Yixsj1usvu0LKGiCr1Y9tOne/Z5X/NpnuPIJ97mFdQxHX4OGjSvYdswcznHb0vtriyCrg5GDrZB
A7hoh5gDCXPBXksmIr7KGhc5R7Yf1Wpfm9QP1qpmAqa8V/FwP02euv0r6EPL4uOxwcuXG20u7NWJ
ateCzz52gPpv6utCKamNWTTpFHY6FMD6MRBsINCWDKhKtjfHKy3oJ1by227P2m2eMSNnIpYcmDll
Nlw/u3fGQK1/Pr1ZvmgHmnOayBVzzVZXsrqrcoyUhvxd6Tq6ulXvR8S26qsu5POhlqA1p1vQfHWC
Rswb1QQ6Opr93I8JwvAF4I7vYvvZBEKIgV8B+TUjWhqYX+Si82FvwYtlcO3xUppXJrWBMrlIzyJY
L4FDsQycuazHLid+GGr52IhU1zY2+a4CMENxRBt8MpPr8V/ipObhn4ZOKw5LI/ZX3WGTvHyxl00g
ukBbJCZ+6oVWidQeezIp8fJqP2T3tEzu7zDHolEZuc8f/1It5Dk1W8KuxF816PiMB11bdja42Tk0
4X0w+1yscV+Nu6bpB21Putha5iu+AUJHiBpFO3y64awTGB2DdqOSYEa4iXwEbWS+vcdQnHl87mvp
kzTIHusONXTw965DGuNB8cNDlJGgsTeDPR3X5dr/vT1uhkhInWrefLe4rwAJe+6suw7MN6gfc0ig
xOlIou0BAio4jmplUABuaX3mQWHR2n+jg5skGJy/2uyChm/jS8lyXAbZkNvj7brzFK2np0dYpm5+
fTdL83g54ACDmXjhibMmN7++aZ31oQ/hx1P+RTIaJp7FydKjZl5oTcmBdwPj6sZBEY4V0YGNODeI
ONBLxQJ7ahyO0MK8obATV90Y5+dLaStZIht7WAht6nKEPbaw2C+Ft4j5dtSQUtn6KVmvf2rKj7+6
iXqI3RH4B9pWqguwBAq0R9CI8DzQTGeKujoAiT/Im9DB6gIZzHSQh2eaDEI4WLuPmB5Cy7jE6P9U
BEm1RuLyFuX5XJdv9DZ+J2KtwV6/BTo1eVQ8ZblF/RPybNTPCjI5LysjPXIZc/W0um/HSmLDtGbF
Ddrlh6zfFPIg5adlJ7EF26E28wSO2FvvIGvIGo3Omokz6AHcsPwRSWxcpZ25NA/ACj1MncMWBQ5T
Tt8GTRoboX1ced0IJGNX1rEGt7eSqk512LntDNrwXst9LxtRPd9x9MZN4EyDKB9KmaEvjTjwjUGv
AufnwuxsidLlrRgW+VaP4Z60zxaJamhQKt7Y+lxd6CAt+pLqjVqQN0wuNagDpECZb0dO8SoGcKUY
eHZt6k+ieo92kywG4RWYCpbS4nnBLHgOy8HGjXMbQF/PLCwmQFWdz+sxH3HLW//+tAQiuuNA7iwQ
pTAb9JoG0Cl9P4XenSBhcSp6Wq+aqG/gju247/IZgkb/Z3XDv29BToJLAVDJxUVcbhU/SdArWSaQ
xZ/uMpHiRAavolB03m3N/KXbaMAzm+kub5Pa9jYTQJPI0DwN2rSgAhKVIlBkJg+iD56iV7/bGNy7
cCqsJwG/AougHoMK8mN3u1UJdkPhi0o1VoRW7EC80dTb8CMuioXERXXMXFo6VEt0adf2U2b4rNp1
yi1zzoGstU878SiAMM42v4X25fPaJHUP8FAmQGOwDbW3/6q2vFvEeEY0vqsdUNCBSz2mw7YfwI7G
O0aLnMzqOL81viI03nTLDnpxExNNdaOuBcJdOGS/U0T+g2cVFuJLzgP2iX/fSUmXQEXVAmimfpxf
SLrCSiTRJusEqOzxhF9DDh4kwG9IuIe3/15sHuZIhoRDZTXWM4Z+bgI53l+eD3e3UPh9gSbkGnFJ
blttLZSKY6APYjK+3Wdbxsld74iUKCQloXRJnQnyGvwvL5Jyb4x08KVQjioYxcyGpWdqBVZjJfLP
hUmGYwPFq32cDHonHs1YBbVY3CXJw7h17oLu1aqoZ7N+pMJsLRy/U2+6PxlT2Khk1ahR0ypaXkAj
t8AUplmwJS+3b12RlwxATjRsKNfpeFBEbc3wFTi5cqC9ENNQak39QFFi96S3Nnr2v6VUOu8nZl8L
bpXQjUUFcg77xRbkv3WcgH/mWOcNSIb2VdMzUHU+HgmN+N+hGEcxr/W0EjMeTuP85wppH9JhcrL3
Dfzj8OQwGK2HufmMA2/mEIUG7XZMygFjzt/sD+6VVQitmBNnSwfIK+aWSMDm2OY8jOHXOBwHii7K
EC5a8Ok0+jipMCrAygBwOnTtG8sbE0w+ovKTAO6+waD/OGci6AzdCW7r17NZ9ssu0wHM4TAv8ftv
RmHk7jqjKw0ebX2880x0Ao+bgDUw9vzXVcfuJsAXZPpJaUKCCdo70oH4mA5Kl/yzYGbLp6z8KQRH
E8F4vPxHh5rIQtBXfItD7yqfsNyJcB9XcgUfK5GPMHk3GHc87BBleRoz4VGi7/IqYCR2Na5s89SN
z/3L4btqiXMG83MTuF9qaaS0y7ALbzDD+F5fA53wVVlTCVNORPpujZK7R++WFlIHO/8E8LEQvd9C
VlkiupX0fa433+J/WP2C290la1/CJ/91pPhi0xgGN9DYyAd4LdA3qWXnjzmSWzPZJ2WMpQkSy2Bh
cpAlHU6uM8M7tHk+qwYB6Y2xNLfT+C63E3H3WVkIuYP8q20hi3ohEPdEAiqYyYS7Iog6UPmDgh1p
M0DQ6/EGLMCLfHS0hLwyi44RroT+gEZDas8KY8esjGDofXqcyAg4LmSmEX94nqS1CCWY/BX1Ge/V
6qHbWABwRcBoIYOmdg2LG4lOjuTWn8Kkiaqf4Uh1oMmw8yR7KzEv6AyhOUDG9KbB20uh42zRq7sY
zk8vTLf4X9vn8QI31Mbodl+ppfqlVjJtQe3/D/70PJPehHRCH20OjK/i7jjQ+ZPfPrOud3gmbFXp
1Djxm8D+MkFNarLSwRo6DHWCYbqpsTVlqSIQpwbf36Pjdw0YYaz1Az3ibxz/oK1ZZLpIadWptMEU
WQotm4L6o96ATcAsBRj+WgdrMervUt2yl+t3t4eBBgzbH/CCBTwrRN0h/PGbx39Uvtx2uRZspYZR
jAkXzH/Q4rtVJ7T/434tRNxZgffbodiRT4MMc4AF5iUjvb4idC7em3tTNAYlbpxMa/h2dpalm+2R
NhpbzAb2LKw7HHVkCRE9eJlg7y4sFkmrXZjSSZRPibD0r9zlBKHf5HQ8ZNCJmIZBuKGAMGzDAXk5
UX4ezVWh6eYlTZLtYbgeNZ8HmCyPU3YpevkBOqzHm8SORpwjAnUTh/k9TMD7kaXVOUt4CmTgXfbC
vlLYo4/cB/IID5HdF1Bo/4TfEXykO9bGgHq/zoQ9KGTUYesBMStoL00NsY7oP9SLAzm1VtRRN81u
aN+T511WSdy3UXDf9XxN/3NO4ZP/bcZSQk29zI6G+Q+Q8hV6Ndm3D006lmbHvNw7IqXDVCINOzK3
d5vXrxzquGE9997XahnVOML1372zq4oFIuxhTedwpoyV9NNSF5kAnA8e4VRJ1ywysxyHvigI0k+u
wgcpZW6KaLcz2APkc37yrwF+F4g3nAv6bZxPs7VMVhCMcdzbFgjU6c2lfk+/aSbOT1ZvsJ9vFx/p
i/FbegvPC6SvwgZWYvPEDg7uyhGYjJqJVVNzBe586l0bk8w0CB1B71x+LM8XDEYGAw8vM/vyDb9z
PmkYD2Vc/jACGBLEOIuCCzij5H/tEsrvjDvMYMxz0J/QJAn3mAObGpyOWFurdB2L5sLULwTgrqPf
FWEgbJ18aeIqJBc4MNMDUkqbqnzPvQIy2ftTk0N9rahLxyLApHVX7SSZNjDAjUbRwFrmPE+syIpV
/wlY0qb+AqS5IqyRwfRONaRJ3OJe9HwLwuc0w7kibLB7Omf/5VyL7uTw7qh+7kvbQ85pcc//7srn
ynxk19HUBxGjCSs+QHJnxY/9aKE+sf3Vwv9TScYwH0pt8SbEG0kd7vO4jf1uc0nAGWBy7ym5rj7u
u0ueoTlXKszfKtvtBJBnlUOaPoC824lE8ct3GnFFCA5dvzm7XEPC8WT5uUM7N122VD5875hpJk3L
ixLYU1UDKsG1LGreT/NlMV1QJp0U9+r++0KSJVk6uiWlrma0D27S9/3+hsI/1iOz1ylUz/ugswby
SdUymI2X54mq8/o4Ar8BPXyJkVT2x6IL9U345NVFCZvDKq6HZMT0DgK1nT/tCaHMBZdPubioCmIs
0vGZJonVX74UZ63NWPip7TVYzmpQgH/jjMlfuUJ4uePJlE1Y7juT/pF2Vh+4uc2hQ+YJNFYbZbHN
FVssZtERONaqUOGCKaq4IejCMFBdOk+4f77QkwYi0Ky8fQFagAs+YFC7k+bSsDWoqC5LQPM7+hTv
3rcHhqI/V6E21Yuc5meIJmnvmfarwf+RAyqVCJgZUauOd9rD5Z10rk4K4MmymqprI/Vx5drLFzjQ
pHZUnzCuW21aoFTUkyMmjuRjnkYfYNqF/mSiLXs3zJU7bYnEgkDU/PdcOdchEepZxmUyZg/qw9U3
JSJ/EUNOKaIxM1oCaoMc0iRYhHIuYE04zG77BLcZyaMtSxkYWI9u5MfoOdqAzDKK+t+Hu98uJAGM
gmn8ZU21lEwL7IpBWu8MljcxDKIgDHToX5ZCIlmO/gGLoKc8jO7BqukoE5vDckfvvwFqUuQansP8
8KHs2CNwNNipSOsqk4cNG8bNpIf8KPQN8wflvT5ZUFoBh/S2IjQyiZuX3HFYsIl21W5wdI0rgkuD
R6R5byYMz8R3lpbT1pJBd51RFlS28ErgDRyNyzsmUdYR+BQwBZBMNlqM1tpBeeMEQDnNZcTLSluO
uZq/XMFpdEm7O0VDRhmTNHTc7BakbzF2deAAGbFakVPapEHFRanyADg7MxoNdfZFdiyiCt+qJ5uQ
+gdnGqyHWVbq56+67hlVpRKsYnBW+3dLj9MFGcHBk2sRzOSJ3K2sRr6gjc283j00wjBOyhyba/sS
lm1/dkWqLFoM4tE0/QofjgqJBTXFqPYx1L4I8JaIon45xKvH/WtcMJV8OAOhdQ7vCOV98Mj7LzcU
agLbADO14jgVvujMd0txhHvY2WzdhGWQz+4eJOwt8uRUQOHpACoJTkOW/zYpF4+F0b5uoi6cLTNm
ClpHN+JS1FNaG6OmXDtiuaF0Rb0kjImD1U0GQXm5gPSQ6d4KCCjV6QrHl9l2cx5SR/JcbnsLDoH7
s0rYKJzdEXh0S/7yiK7WVWK03s8AmpLbJt2V6B41vQmLO2hV5OT2ejBHxllNvreD+0fMM7MKfNy9
r8y660mHAwFsLw+S/4t6i2JRvIGKSQcrLMXaJSGmNS2eZXuKt7bilQpblgkUapBtNWC9GuhS+NC+
6CY/AdMvzqT8ugUxsE8CYuUmDZts6KBi8AU+jkVbb9moW7BWTNyCmzSGNt77osOdbLjY7O3bwQ/f
FSGFJ/NGXBsuwHuTSoCUbt843RfS6Ij4xGf2Q7ZYbvXIzN1uS4/YP0SEbsoQV2WAoMo66UcI4IzJ
UKHro/wTJkyixdcgWLPRFbB+hmzDOAyP4P4gzDtQSx13SmcrYl6mcs3xfOfraB6trh3n9vQczd0D
s/aM0Ktus766gF19/w8nU8OTulI46gfJZrh86BbqjcdI7agL3ig6bw2SqFVgsmmH/wKmbUxtfh4P
vm9KpUL/ltVaJ6ZHrWDL0Gmfy0HDZxoX3pr2ExknZ/6ahZ73OeD6jh9jgw659su3i8FQpPRE0R1V
rPtGCW7hkeIRGkV/DCafyNkDcY5VGNgXDJ56bJt4HfIopwvdxcU9yC3zbQzabvu3vtM5qxd7jGvE
V2aEGbAgRiBZ/rsYm1FIJj2epMt452og3DxSI51dz/35O5iIJNahz/sSusxyfvXX37BIFT8jA3Nb
f4wWYnuHxKmZhoU/3FEZMyUw3NOXnFXCtP9wCXyd6nQ0eXReV1hsXyYJcH35Xc7MY6eUKRsNNQd+
FRRweVb3ekYK6wkG2rHANs2e9KOb9XmCFpDu+Nky9oH5SE14pt+FmxY8Fi0wYbI5AS4Jp7foEiWh
UtK0sd/LCfXybsL7bcij8DRY9ylWVxoC65oYJTmtyvsN/9GAX/sNFREWL2ybf52LKIJOGnUTOEmD
PSlDZr9/lVrJI+4Q8qVyc42VsDTnGNF7XoJfdMvPk75FldhPEsL41nMitp2s/31/3eDM+htKc2Q9
75EQ3/u0r7eE7zPy0fZ9vHmLNC4OCOjD5ksKaqts2Qn0CQA3Vd7wFTFBd1UzLW6kEF6aw6anFDLw
oUUH8mH7i7MN4asOGSix8PvheuEpqeyQdoFCg50YyV+RMVVEOoWCOoxZTscvLe7WBINnMFMmIcJt
dY4Okvr8LBdLincu4QX4AkfgfUvfDFUP2TzBq26AiZcxBUmok0Pe/0iCdADKP6U6X0Kq2bNoUB3F
C3J3p0XMt5YG8jy+Chi3mXh4stkgTWbVSiX1elPR9s+OpjPhhoNmdokivJECKiPU9zZOH+w6dHl/
fNN6OMdxW1u9ssQby5ziLbOpnfd0qs1Ivd/KNs4rdzLx0dT9OTnAStyXjNf5suIearKgFT9icyaz
2rkW6yEtCKqsJLGL0wAfSwoHJcp+AR5YEhYNWqJzOaXlAlfWzSpQBOsaTCC7LLkv0+/VHuNdOuXI
B+ZEsPUplr/rriBsbXSnzaCmxucLY9BJYHeGyDuVhe584VXVyNDBbKXBjGqqF5Y2jnHB1cAPYWlY
ZvW9pHk2Qa1nbPETffILkv+mxWhhP0oQ5Yqz9kas5A1BsftPu/Hl0RpA0LdDP2ZKfKBXMmk8FZGR
N8GHpuSjyXvl+E8yBtNqcO65svobHuKMvgkAVyjx5754ydCGhhSUZJVyltPqDCAzCvpghTzOpMjI
Qa+G/9eCW+E2XKBfzUrBL+t/MVSHuLjkn/u0A+wcE7kQ2FTwZ9IHvlgE8r36t38i3KXcETErljAP
NSfZke+lpfQrG6qg8EXd4hxilyQ1qYOB224bNN1sqSqlUbMxhPvBZXF3LUpV8wpYQtAgVvfZXwEM
oIkRCNw5enjeTVzlxgDp3v17xwkewEF+KJJDDQIQMclVLCbfsshAxNgpokEYAv3jj53MpHTV1ZWJ
rmiWlsd5NWCZAx49uivKgh9Du7xTMwcThiKA/D6piUZ0QMQmyOrf0ydu6M548icnaa+6B4fQt07A
jrhtQ+NLqOAfwiVzgYsxTP14buHaD0v0X31MGPg8Ddf1Swfffom19I43sGHt7gq7ilvLaWfiLE1l
soMTEztSHdlI1OsKbQvFg3cT3KjnuAoo1Wt58s5/oSc2qj5fAMBFZUj+cb47li7lqzzIobswJKr6
krc0qbjNJCJ0Deb5OQeG5erD/GN/2u9Ufnz5O92jyqgXWBxsf0EzPRniYHIOh6ZflZ5lO/f2XDmk
IsVoF2lHmGvsrYARAT4M7ZfDSvhxG8cRCtHEBwwRf09GRp20LJibxsN7Q6ticCPMP6s9RXZ3lI09
dw5nbTWy8ZdiK7OJPogtTSfhmFRjHUeM9UAL+W4kmLrWSU3aMlcPvRjaC/RF9gNTo1RfS4XhE05Z
qy8PBgSGANSbsiS2cIHOuHaZ0BqTCuKOhHBSSNTZzS+Bv7lHt8fdT5hxul4Lh6+jwVRvGxQeWL3P
3Ic6aIpFCaTBVViTkyTs/tOr32hBQSmbilOQ1MhNcgBji3CZEYLyUWgtP4VgJYaSX193xnIz1PDu
+O78XdL5ANCbAiKY5a60LSppNnfDkGp9QXUQWFKg6elqY3Ez5F+MMqynYd8QEB5A0CLPVyvdmSoI
60CkVG0asoRDBBQNykDJ0eakkHR17YoYxDNQeoyDFm37H1fIm8ImdyjPjs4Y0xNBcntc9/9XFAJv
SbUqc+6xj6Q18xS9CMSyFBD24LRQuCkiJ/cgc9+MUoWllFfnHYuoT0ft9YjM5sXOGx5ycqIK4El3
RP0I+D/uxJaw2CoCjzt0A/D2P9/oNnYtQL4kWYusZS0SR74dtjB9NYOgTHz54BjKT67oTpfiiga3
ppjWH3+UBg5a2QOf2msb8c7CNi308bpsbGNGmWPwkZC8WFMpFP1ywT2TP21OrurCI2zlLocb2zbB
2iUqcPgJeR5pTVp4fatV/CsfwymXBhEkh38g5fXgz76awemy6UyJcAs6bbg7PnlzkGlKMpWcOcy7
A9pZSfCPi7dmkHykVcCULxGcrCtVOeI8v+wH4n62c39E0ohvce+BBDFYDjznIOMrtimFMQxy9FLM
Pxfd4DXWffl2tABwINXLNEMi56fw+sHU+glkYC7KpOTM0sMGmKsvvaLXQgRgQKTJnMY3/DKRVuTU
Upt0EJEBb9stG+3hPDBnm8aGmq28EdEDiSWCwmgPJN+U61Cf0SXv/9U3SbvCB6JnxazEiYOYGZmH
ozqByRMwmlXFHdw7rOo1aUXg1cYgnDApKkM1kF37f01jRvj1i7ydq6QMoKCz3rwNg1POyM09e0F0
EyE7BRxevLZndPSehYtJKHyaij2Eh1cALHnesAiau6lIic/9Hhoq6Iu8kGAQUyNRPDUcmpzS5Xs4
Nj+UNAJTE3Kce1irjqse+daHFWzQSrSjwU0GJTxnZBxLnzMeMR7ikeDkyTa7wazIGZx/v92Ma194
2ujtbaXrOjRAaMCyNxNFsiZY9AuLFqs7tR2VT3ojkK9zBZseWG9UmOpiRdkI5W2VWrUhBXez9dwS
1W3J6SgALhj2MDn1G7VK2Q+jnk/GDHxAPa/VSMI7S1dPH7Ol6avnd9y9h6osW9PsucgFSJ1BLZDg
DwTV1LjE2s/NUOMo+euWTrPq9Ognc315go6Sfu/mquWaizLjinLx/wJvZduwTDhUU4XxPRITjh+i
0ZRdcUA2sGfFUKk4TnM5otZm9VDhoUcesboeE+Rk6UPe4jnRRxybeXIiYvT43FbAsjwy+PrWDIeq
bcn1s15h8JEsIG0TwNHiIGJjBlT3IXzlboMoJS4yr7DbvcCWnU0w1HZpoHGd2DsU1NLNgGw+zxvd
Ouxn89c8Ub4kfRfp+GZbuujZtNpd1yu87K1/bpdqj2KIMu73vIhFfCX3tCylP+Sc2MFrjow0eM6h
jGC7TIAvLKkI6vLAbRX6JbWF93X/NQ0McIVdVNPgCq/8T6Dx381MC2wST2Bte/c7hQsn2YfD9zZ8
uaIBLN5GrRQxQuNhnSAAzwlUWnxUq/dcMggqCFu04C9b6ntMuPAJ2VUOH85wjY/VJ2gOTMpWEbEl
fmof6tMetF+NuYToosWe6eepnnDzfaJ3VDkMHz8s/HMGfNBrle9/UhM96YlsjWw8IrYIxF2aJpC3
JCSG19TVP2jvXDMl08rcxff2xFbW5N5zjQUpw4dU4mFJY2uP4Z5MNKq72t8dMahV4NRKUXTekTFE
Z0Y6jmspzFk9CMCIYK7OgNCaWgrZujgSIqA9MZrm24cMpYDsDFomh71AR7ZAbnSRoUXOH99sjZA/
eO/j/mzQHxK2do9mjcZIH3cfAUpvJTv/cKEmfTZEabtnZY6ifUUhAucnBU02YivGjOaOHSqlws1S
nPlAdpxEApToLLqPYwdAgQjmbedj6RD2nQwaQo1uOx5ygS/lxI/JRWp9oBHP0WjDwn+rUI0SXa8t
P+9osW62jgF4tZqd9uhnOoJJI8JkyHUh2KvAz0XunmUGnQsY+VGupdJZ71f4Zmtv59xg/iKRnCM9
4pAYmB4YSDt2CdaJTq9ov0h/E87E0KgSM/6YdFQ8lABAg0RmeeW+Qt3Wf2sXc2u38xSzw7g+eWhS
XT3af1xwodCh9C8SowKYXk/WBwRsZXayYC1v9zoAYSgETrr4g/oP/rcEU3IPSrGepzTGPdwWFQE0
NiWrCFSSRCRbVpiKps5TeY8m14OQPVWBQ2iDosWZ4GI0AtJtmztCflCui0C6LiTvLTmOcKvIPXVa
5mrkrgVDpBWCA0K9Ykol75/5qaCsS3eYeynvnQr0Ls1z0nULhR7SNMYTjxRH7mMBJsX0ycK0Ct/g
5ya9ZRyS0+GKC2Suk4wm/8WHBgWbuVMlh0RdlMux3+WSF7cUaZHqBl5/YWRFBmqpVilI1PI/W4pD
3z8KQ110eU8/xDvGxucYFnSYVGjEBWx6PNKqvluv6Ue15vLyUWmQR0lX+3uN4zjBFIL/ZuxR4IYT
YqDP+JXbfjMdlTsFnwVxZ3BdPLU8E8A+ZW5j6i6kLfBhGyvpbCTf5kA++D29Ealx0/u2uft5QAq3
R513CVmryOfnX5fvE4IXeb+k4qK7YenQ92kaboYQsOzSMATktgYoY0qNRZ5MN7tUTVvwXfXVz4c7
RpJrkoMgCCbUI6nPvleSUqiZYtk4/ONH7sthhLP5LdPtmKbdFR305Gz1s1SEbPsqhMqJq8Z7yRwQ
+TEm5ngKh2A/+8Zuf6dIdjupzF08zyH3ESXTLt/0psg5zhsOYfl5IBtQBib6/UvzQrEhmCELCIRQ
XhFFrH1IXwv6XIar3vwOmUFhRFrTA8AR03Wdd4+38jnowjLjtSXiaCbSi3mHAh59YIW08Kx6/OTD
ipu+dxfCgiIUOWVP/NwNLWh/kCD8324z+O2Q7Al+AkcenZESnWQS1blQLyDMRgeZq8aO1YrMj6XD
rrZdWxkyi545qaFFpXbd/lV2sUD7BnvyfgcpA7qhYCXk6r0nwmZo5fHswPnAzz7FvDXS4A/s+vRx
c+WTfSKyJb2RK5Rj5epjrN4PTUhrJ6palQclmOu9j0PU0PVGJ3GlK0O9Zelx44rCnGMTuMh8n3qZ
b86VbNgGLQVU5HylCGQr3RZCmra7hotEWK++bFJpZT8ebcLZgQ0KsE2N2UcKlG5vf0PYKeUhBaZ8
Xdtxo08r7uyODpg8G7m4wN30R4KEylFdnq0oq5on111stQYKne68uKDt4DWhdW72eaN5K8Q89nUC
QuaWkTJ1r+h5o2O/ZMxKECoHBRQJhe/IE06kQTt6GooOcc/KGx3pyanT1lPO3Dkqv25jiTJEVWbx
ce6QUgzyHXAdjJmdloRSAqqCYJt4Z9eApTGkpT5Ir/sWwYfDJfIi4JyLqpsYo0EDceHouUufhMOp
0untyIS27DSfq8JO63D5IIUBXe8zGPJva77/oHMREg+cerfG8P0dJUpjSBvq0v23Xz3DTVhFV/v3
xBxU2r9apro/GiWw3EwfzIy1l/ui7eTCOdQ9ren9LLZ9zzq8PabN/4DP9GLOUT9zCZWXJ9HNZ3JM
kNg1wHOUz0Tz7fAWuqwFvsuYcWiSI3woOkwBJkDH2mhjyIvt58ZLACAhF01xzwXL7nZyaZLZoLB3
y4gJIs/PbF4nTWODeSsw347pNSvPTr8Y1YHbmGp7LbGPvdx5RStWrleWJR7kTp4NIdJwI752YWLH
ZVmILv6nM9ZqjfiBEYtlhNZtpnw6Zc8d4HI5Zmp8jEPE1uzK3qrXmK3a/lybK6HLhnrEegOqlu1v
03Kiw9VYRLtbOU7UIQapn2DFne8RtokFWMNynQBK3VlTCQTHy4hR5DthuEfP6x+RyyUk1u39R0+W
I8Em9r0rC8Kih0crDSuoZZVSY3HVisZ/jO+nkxolaSkFU8NHvFegi0NBIC/FurUTlHOrqwR59zhX
wO1Cn9dTNqHNh06N9aWTgjTxaOVqZrcTV1sCNh9OSSbkR2Oa6MHJdViP4cQCzPRAdnfmM47Zgx/g
FWtIHvo8X5bVc2ju9VqMvvtlQUHTxIx9B8jC0+bvM3rFPYNwZ8X/Y63oj1jkroCz+VLQSkt0Xmkh
fWxhNxRcf49ijMzKWf5jdk/MPEcdx5BNf0QFmADAoJu7dMdgyeqascf7GB5uxpvoGjHKDn/aK4pC
ennIDfGSykkmAlo5PezYqqchG/LKsQC0F89Wjc/p1sdFJbt8fjCtKmkk1GYTB3lQtj/5p31xVcHg
3EWSC5g5uLviAodrpE2brccNbu8Ca+GSTA+8Cbez6zJ7fq56ZJR8afn2tdPZmV/Lxeo599xLqORN
SR2/Stm3Kqz/bK9g3SoEe80kbxg/Pc3+7SZFMu5L54wLaRERZaB0BRVPes9KJMo84CTRQd3FBDOn
B1D/mdCkh3glmlIupdPn8BigjAMbkbXoxESdGrpzzsAcjB23p0T+NV8Osn/UceYzVHDXbTS+3syo
pdfbo/6zVHBbywGu4kViRGEzFaGqpaZPNgWhWheX2Vk85UHMsM6Oxhoo/Sj+R6f+ObAkz5duC8AG
YRzjKnMwbkz+/8YSsg5UhjJSCC/6YPVjLr9IvuuZ0PZSm3bWtwsfg66sqi03FU23fA3HNrEzOJjH
WPe6XVsMrVOmX8y2OIOVKSGN/w9s2pENssCiok0qxPxtd/sjsZPBq0xkcjUSrMJjI83o3IGvam5r
N1+NGhixBBzxPXRC+/EtVvDQbkGfLlXVktlRwO0ou46z7hMkO0jzLexzyoaDmv/krChpZJFxPpZc
lw8goN/t8XGH48d8+yeO8R1qojVeb4ENRwHdW3+0Qr3ISK1cosM/CxoJ3hc1YP9EBEnhPTOZVRov
KdRFQecwHdrJ1MPl7QvUJEdBHQ/gg1xQQIEvISMl2aGDEe0hnIqX+I08x+6BGW4ZzxIMF9NrBZG4
Wcj2zloc5JnaAPDKhNaViR+RFP+hkWHDv6XjQAkz98DnC9lnSTbjM5xK6fLtILIPnPDwFveJaYQS
HSBsttuafIBKyM7UqNjgXY0ooPkeCHA9GlAdlI6rtImICaygBg4tqbkSVxylfhM3AoFgWwjwkZsL
a7QFTg/V1Cpp7ssewJwqbzKKyRmu8RXGamSwZfAsPozCIT0nBVkujT17O1mvK9RvkLN5oRVZFSYN
4LFx3xaxjtpQS6MhW5JS12JzuorlPH8wV6J+C6wqjbRtrI8rkBi0Q1KG9952ejAdt5Kgo00koRBT
aakyEKf1tVAmLCkgw2lXUsiWtbdfSsj8Clswig2daigaVk8e2/0CHkqsfRNY3+DUTZbuyZnYc7G1
poOkHv6illzQXwV2kA79UGL6b9SpGPd1ftGZLNTMfSqTvD8BejJd+HQD23PShxYvW3Cut5ISdBlR
JM+TXT/BDVGRadW8DTEild8xm5ySGjsgXVrFfkW06udlenCfGENQ9/9JZ6Q7ic0ROJ39BY2fu4lK
H6Z7reeWpD19djtBzKZpAM2VQOBaIT6kvYIqvOGcDl6eE4FD4a6lE97zO2mqEA7oR3ysJklSbfrC
XbiLoNrBQxCbkKCjubgMJFO3rVgJ3jVUm/+0HElNS+0C41HrfKBVrr+AjUtU2iUbVgO7wTM3Vpqf
X3eR1H1kWCkcPy6PPISiAgEYxUk/p+AobGG3eMf9EahJjCqPGz0k7z/b7qaO1trEK4Z+L497MrBv
r23dszXOyYJD1pV1ek3IeZwwpywfygsuzJtq91die036HEOcw8DcYI8iSeSsdfD2xE8GuRugFE8B
EzC8ebg3u+fac+PvcJF46tyNWqVy7A9JJsdYYOIcFpvWpdrQM+a9xaPxo1XDByKyM9hY3nLOX67+
eLTJAWXFjtMkzxjJqaPKIDV6Xr+h2FDtQb3urWqv1Rjs4jJCopqZibIF/Y8n6pcodwsaoOBPj/LK
MHKAFAfMas34qNo1ttWUsuHLyqQJcmP8Ui409mG9EeIdnCnN2AITeKoB6fvx7YWGWkvr1OP5fMaX
V7HW2klxrFadFkPIET4Rl99vUYmJ11CU9A8ySHVXyNQYpfCkIr2DJFYnu4LOZE+83V8VQLaphPvx
rl7oNDioI1vymH89T2jUnkwDwXXOiVXy3MmLyI/Djc5A01BubOfP3xdbV0A4BKnldgLb1jWWaECs
5JiQN8x7Enih1CP9VEzxdk2CcU/QOFCiBACAwZ21viazwl/yO0oZAlkyevrp3yXarj3DhXOlyW4C
dU6MndAWtlE0sfPYFMpJgAphbO1ZyOupingiztinDdXdzH7xKKaVLuoUlyTXzKlUmdWkxKaEQ7Lj
SSzfp4WjmxtGu9HtF7s/OabqdCEpZ5Ei/W0ePN6s8BdLJlOFM8gHyjNWs3dyNCqzsHYDPWM9QYC+
UwYGaFzKU8jZ6+q2vpUjYiWdDcxiYf9kIN3fejk5KCtIfPQSH6u+dJHYYy+XURLbJfOJMdu+PFEH
iKXvhMP8xFpl5iWhonnaEbKAyY53iO/xyzdV7jFvYfmuJqu+aEvcV2NHU4dSnq0f+Uuf7HbufVUl
qPh+AvDAo/mVsHfr/M+fXJH01LV9qDSKK5+a9mLlvfTQYKj6WhNXTzF3Jiyo7SnrjUSG040yhymq
NBXwNrRAmb15rV0YkIuunWgZlhJL5wugWAHmke7gVyoUa3LooPmx/PUxd/qQjQIGpLofL57KrwOp
BAekd3LrPABcJnpmTosAs/9jexsuv8nwMz9y5uz2w4e8fPV3sOVwCzGMtmUDs8rTNSMYdEkuw/V1
BVdbetOLD6Q9J9Vc8oNJ18VV3baLgpc6yumD8x1xUsC8WqGt26c9qMaM2YMuCk9Qge133kD+Dkg6
dWJjF3rKjAxQFl+gu8UAyZDrWEHnZG+HKlkXYUXR5Em1z8SurCcYZv676U4R0Y+g4QCvzkvo9WuF
sDQxlXA+cTYXmNMvzF+LuqYWAUHzEnHePgnlA1h52iupcueR4OT0kDTUW6mxBhX3kSCfH+ithS6D
Xb1N8Ds/3YjbkAW8sUsHUS9elQeo9XHXl58fJPTe9t58E59YMSidVQ/6xW1W1G76chwAaxvhJuMI
eTNxRIxxSqegfHQHwDi1aYhvUYtFae7tIvyjePmpkR1KyU8nO8cw2jy2+g8IdcoawKExYbvIHwbK
eggoZ1sdFWNU4dtkGDjxMmSv0DwstPxg7uUNETwqlXj6g+3okLntQr5zNZftqFG6EXwueTE4uR1S
0S7UNV8jbjj+atTs30Pr71owSiApbZavth4BcB8phsBej/4TSEx+5gRuDt9w4F5Obm/kFhUWyAco
wP/bf00a0G7f0lBzM4w8bkahFIm090ednkjWxSbodF9Om18DSi0iP3M9UzTMVtTo0ynYD/Kvf6vC
UWP1+Hy6l5R45Zr5116rNieCKwW0Y+b3PQ6cCJVd5FCyovRFPwyVkGy7GIQEgB0paf9dXCDT9O9Y
NnbRN/aC7yjs36vrcyLviN5LT5+bGf/HQkjk4pMoUFIABn6WYkzrSTzvBtNS6HC6P9R/6WC1eiAi
5gI7JZnixdl6/FgheEqPVskwgGFAGTbiHEZBDw7vUt3OY7w3GNWVwhOibGdc/1LH5zQbvVI9L+84
HX14xbAOEWjOKHV4PhsNCwzAqzwK3RgMO5DCvUP0CH5pQEqghoKf3k2fnPlNdxjDPupJUASPoe3N
Q3r7PE8d1Xg2hisBP+awPQIXRxMO8/w5y4aWRwGOxjrnIvU0nPnmXtx/4ZKb88WlVsiMMFyokYzv
ye6Qf05XPQ78qf1AXQ/b6k5z/m9tSyb9MxIYLeTWJIgq3vR41yM7knefBTRwlxiytd/x0csy+oq2
Ck3mi0o3Fud2410Lr9t/wXz3KQurmNq6xUZ8m+j3PSdZ+p7+KkPB4NkAeNT9Pl83ahNMH3n8Cfyt
e70SmCUx/UrI7uyh1doODo0pEBVX5xdUCQM90OZH2whP/JuKbZAgJs/p4Ubg9hN1T2vGiDUc7U1e
TfYRJL3Y3tUos+S1xRfXTPDfz+8CfpauZzC+a7aEvScjJQd1FKIYLnCATOUNfPbsuGHSgcmoirH3
KBnPtl83luSQQab/CibcyuBoToGTq2v9JOig8P0BI9fw3Wq8ePk2Wul/fysfbZtzjlLXP6PnMU9w
l+wrfGEWYfcmq6xh4b2QQ0TNKOXFdcXOdMfoTPoObdW7G0sS6rH1SXBG1zJZW8CCBEukgUhu5PGA
ehBYnaaoV6CjNUkTaqi004d8quSY134HqLojmrlvexn42X/Ukmc8D8WwU5SEONkUg1kdXJGIl7PR
ydGf/1ivyNhP0nbnRYFSdAMH7DfC/f+7wGrmYY4wWAugNADoOm+HldVWMJuKpJSaSLcLC3iMUyFP
aOJ6y/e8jtX3d7vQNLZX0eXwC4gtmJscTeawvrYs7+FG8Xvm04D9a6t1p7ZAQhdWdU/w7tXc57E2
tX8QaD5DBj5O+nSx0Kq6YvqIliwYTIldFSkEa+NIR9B2xcGHwl9LdKwU0jGJjOspafYkqYdeqdP5
xaa2rj3HheBCu/DrnJiBOO/2zeNcFHgL/nvO/XcXXNHvMcfMOlWF5SkWIZtYs7IxyNANSYz/O0D1
nP5cSzA1HUxMeN36STFZDdV9grlJzRZKnejEEIviGyh7vQdb6uDkKQ5Xe44+q3l/E5RYLR+7HuS2
yzTKE3WYPc7eDkrqh0bk+LHqdVW5nlyMXlWjkFsUlRcSz3sQpKWswG7T4GLnFI8E/qu3R0QyOos2
fEEjt8l4iR6bzSjxY8UcuU7PeFOR5dOuvjRRfdPrgMgfJkA96pf+KlfmPeCeko+I0YoFOHCO4Cfm
1v76qSbt/59yNsCOT4sd585FyTHsd4uQlr31mSB3/c5QolHxpEYFSymY/j4eowyjJHCKA4NaJTOg
EyPeYz8a7HhHlFb2LquTgZOxL+SkNa01imx44A72Sd7PkrbfUcmvu6KaO6H/ijvcCCLNdU5yASEx
xBpJo4S4y1U8MoDTN3KsDoFuTqqSX1JgtKCQ+QuKj4ybWeqXi7Zr3zhBrmTHnBzfpKRXgE9uIpF0
rZql+Qa9npum4ojMZwuXaQPqyKs5WFbkf5tdT6Phw4hOhZBFRQSaRm2OYyjjcBr+4c5hhse2+E9c
fjI9MAC1of7HAao/PN8/j3mRDhi6eI9Y3zSuMdZyo4XAMfUh3E1HYGRwaKTgTRLKyXCrFsxXNtp3
B1ScFNJMgTkp62HNVs1Q3P97fTaci1l6oalznYFP9rMCPxtt+mDM2PLJlJQ6Vb3VZaa3mCLrLJIb
wMbRbB0OXhpUgBeyTB9qUMpgwB7Q4ZkxXyLnl+ysKWqM7mJkoCoSw1Q8M7KiW6hMTVnnAkE/h48O
BmNc3Btn28lgOgamNOZsW4MGdTxQ6HbPM5FoHrlMLOOQbTrBfTrZJexB/QwEVd0/Mpxc+6Wyl5+x
82iRjEVVxbkDBQ3mD2HV7OFb72eDYu4Kk6n7C5BjvSFJw1Pzaa/JQTishcbP9I++Hit0/gRlpfWm
CvgQOVwKJdhVmaBOpLfPRfwwUBItJFuwRdhZf0A0VxHFC/75CItckczZdjtH1iSbRGiNfqkFLRZr
max2HS6pXiIa2OgxXeiDK6vhgKLQjUPO/3Wsffe4k3fVPefYYpvm7KVyaIs55vwnCAAGjNhfIL3Y
Qz22TuY9HBMn0DCYzHfP7+DBnoiqUS621FLGJkvcPqgDtzkr5XzpPKHHIKa3nPai/vBfOotNQ4lv
EnJO4Hsx3CDdytcmj8unXUqphQcGc1bNpWHSX9E3gnxYe54h84odHZ9pmPLlMS++F6FmFqNEATV4
gzttjFuUefKu+BcY1lRnPHFYmnC/eA5Urf2W6wWshaSdd2qLnsZ4eHYtB8+qnhNuUsNxh8NF//9x
zJLZX7+uicP/++ZkIhXjjv4DCKDQBTcWCxvQHrW863syD4cnVjZ9bj01bb7VXdl/rkFh2gvI3fjB
Zxi87siQLp9lgRYFOomIqkC+DL3DLVp0vwIsKIX7+gNOjMVBDwKg8gwx9qaJvHFdJxF0qBgrgbxq
rccBvBw/9kWdGW553FJ1ddxTRpvF7dYq7tMuRGUcGr1iXobmxOj6QERVSW0znkFI2OO8A2PHD4gu
MNmpgpQdI+yKPe8YCjRlV24APHoKSm3xneU8fdhf72E/fAVbAhrsbjJsdrwGSpMFp3uL3Ur//wnZ
lfEvKnEFxkGT/5JK5QIO5fLNjI0Y3TM6WnhpRYTuLWrh7m0Fjr1tloHcad80pGB1bCW5aNLxk+S8
CP8/LqKZel7sdKs6K8MDyyV2okeKx2zgmNv7wEN4CZhLEb2wwNCGYSPxS4Sb4HJ2Wx1cneEtGoNn
ShyZT+IhoNfvMn+nk/NZ+R+1bL7olfn4H7ECDSPgBi/JQJa+HSzf/HPt+VjxA7sByGx7b1axaHy1
CsUoyG5zlkYrZRdIEaFVG62CFTgELSbXy41NPquyG2hRruWDqzTKwq26tpEML62fX4O3i14fs2Qr
uIpLpxiSdE61Zf8MzP5KlOwW0Q+kwnUEqvjjOPnEWBA+dq/3m/xxxWxGQQvAMWCbl84LUVIqCRHQ
U043XsXs6XwCMrYtODNnAtd9NIvJ1Ocmfx9ya8XyIjGTEIX9GNA2IbLK5bwIW9m3tYoz1O/ha6Y5
gWZjAH1D4HdO5swx1OFL0/c85zhClzW0zhqArOxfLW3+O7MJOf2FNkQUitr42YJGIuIUoyfvF4nD
o2KjbB1HOm/qd6GE/qdJXJ1W2iOKX3FGJI7dDkGzE7vQNucyigbV7abmvROegL2VcJwi7k7ZTEUB
raNlswKito5owPHJ1fFr31tjhPBqh7wAGgY8YgLiwe13K5hteNbA0SbmFEepBZcogxzgN9iTE+IJ
PIPPiQPa4SrIB3gwD5aGw0qmfrlJxnii5K9EsvH7YH5hAMxH+HGjgeK0Rg1+EMg+KFB+j1JA84ub
AsA7ENqkxsHrhYoo2Ql6qaUEfmJL4eesknKT3ZLUR6vMGbNQcg8Duxq7lTqWJR7Z5Ero0QHXNWQr
F28vPlRKvIwjMoB23G80eyqBM6cYcnm4K8GXRAHfiPHaOZC61aCeDcd+RJQY1oID/9XcWmMYHBLJ
NvsvdIC3cClwqo06hn2gMweeixVJClSTLDtNIrmcCw7h99ZGxUf1nDW/zVC4WUgOyZV+KvgztJRN
fgAEWtjkOurAEeOhHGy2vgNE4geVTkIQ1hm6vGMWwkGc6/ScZhIJmNbWgizJNIN5p4HOeWUHTnPF
najoPwDez026yM8GC0OGESjOol5TwXUd5pUac9qfhhdObScRQEG4Iw4Z7PvYGpiYQWB1ByuxZsiE
Euv5WRdnd1SVhknnb8XOOGOECAZoZgqOCVDp5ld8djxBJqmWFVaQ2z+7HkzouP80hiIl2pi+rGGS
2slcpzRpPuVebfYldibekcg7JmgLCGeHmAlgjQw/wAjNRBPGvD8OXp9hcEXvqcB7sNICL0CT06ri
/BIqfhZkQj5aZMGJAq8S2EfVHPNx43zi+88t+9qFbcwq0/TWtB2M+yOdV1vzCiPMkt5moJdlFC/k
treCtxpbU6n9lC1Sr+OH9lE4YTm99K/Kun2l/VZtgvb2qtcgTGBXHttMkcS5Y4fPFvoLfi06gjHu
dZEPB6WuvFwhvElFrbS8t+XjYGB5Y3wxGBuzOvj5k4mV1Pb+Db9Vko2tjMSW1d/mmA0ySu7xLR1I
d4Tjtz5VlbyWZ6/DRQOJtb+l3bfXHn/vuJevtacM5pYCB1CkOQxIoCydNwRbpHefwLPuRnL+cNgO
9SKPdkICMyq+ev8A+peDlBy3xkkAjG8PF/Zv26fbO5gw1tSCgQc4/VGHpzrlehIz2/eAyt8cmHyA
BpXlhagyTnb9i27YR8Wrqnnaww7evQ5hs2QDgYFi0rRiSJJXLwUQ7TIwAJ/I9JEwDixX3gWqM7hF
cklai4jMn3IAvFN1mHdB59PCxrMNzocM8xY79SgzveeozDH/dDhMX2y10O7YZHYiCv30kkJUQu+3
mCJA1FcNaOHwOCVwhAiIsdMjOU7dbPMb3CEMyx6nrCof83NWenLuHsFCtNKur1/Tg0ctZa+MpZVD
HtJnGM4YgpTr3QTg0tRNwwcWiJSAN0+z/kSJ36DzyXrfWWPWjE7YdRphJ5Nq57jQ5c03CS+POr5/
ZXWr/89C33EG9gxCushi1tYA2S8W8YmluCVfzoqHu5O7xM3oJ+VwUtLdumWSGx2uP9Ji+r/lUM/t
uCGWgF5PZYYUI/vQMTRM2BsNgB5SVj9Cwl/ldytmwS1i5itLyw0+54/+9t9kf0bItPtSYtrix+Xb
+K/rxRoptsEERSDIW7PjPG/IpbDsVUc7oUax2u7q72qgfZs3fmfjqxcoRIX+eVxXUDcFiBkUyWom
cPlH7p6sr66dvMJWoZUa3RBeSUqmc7Qj7AUipfO/05reDZ8QToafqs2tla7wwVGBw4h4Wl2+tPIE
Lrk3AD/h6ShaKljN/I4HNjCtoJyBLREmNxONjE0/nmXayqubZfHG+T3Ds+cG6BCpi78jzBALIo0p
lgjLhV73DPdodcPliEj+dy0+IDFT57vPgKqbMLTpNSq4jCYhEUsop/eaT/904ITVTpAc7ebnIwiw
JKSDjx9tE+Cu9SFpSClMVQensEY3fGQa0kdic7RO1pzrVtpXCRPMb/tYpy6d38SE9v8bFj+cOpoX
URf1n7lIatHd6/F9NWXb7dTB1Gbu8R4KPCX6M6hVIJsURIZ72ISTg415yh2uYVcDaeQAkewJau1o
9ZcncDFnzoKHgPWrf1+1aTum96ZRFfsGLeyyvdWHlUsrSsMAHT8eI9JF59g2K9qVnV9eCPpfU70R
E/gmzEbr/6dmAxtHvDvvDFJ/4ZYOuJQI/lYB7ismAKGGgSwh5H4TAh/BWsXS6+HzVuU6Y0Vsd3eq
yfTDJfB/el1PPUprDj2PNbud/ofkA9Tl54iS5MDLK5VVrUwohBz2v2zMItFP2cJkSUGC5P4XEXYh
1zU935O09aTCCiqHuoeButwnsLPbfyS1YXFKFkHTH9XDUH/++pk1hVj/OmQQjDYIKk3U0zh5PzaK
q47KCprhe4gFZakZ0awWLu7772RByxRnVFRf/S9RVeG1dkhEAJ9Erv8lkebYiaKzXgarBReGOTVE
/vmkvglr6MC3/lrAnNBALL8F92TrLoPKKGmyFkzAqpxh0KqwwqDkddico+kvRzd16dAmMgm0lxm8
v0r8C4PsOhDRHnmuANpiE00htuSJGy09Arow/Z6NJiHhBb3LzAG6hhkvlfd09BkE8nwwimCb5acl
8xfawYNN02S8oRFWfmN7mCRKQHMkA5a+R/OVRvyFlyOzZsbadjTQpE0oS/LD9suHu7l3M38Ug6jb
N0Ji6DoiL1wqtZrkH9yfuBI5mRVpLXRNwHra0Opfm8Qs0kpLWNQl+/E4V22U0f3zxIyuXnvJR2wJ
aFY3L0vO0fQS2ieTXibHpnRqQARlChcIueRG9GtJ4tfardBiDX3AlUeGWZqjh70RCKKm24VCX/b8
UITKrZne0az6NAFkeTUn1dJAQm80/urQ8n/MA2Lj8Jqf2VjRQx2TWbEXH+HAHhfNRQo2krRElZUo
B0gjfGOLDt35WBKW2uLwEoqSLBc1wyFw/Su7fePQjV7oxgtPAz/vFnBDcdDdwzalemCVj7syGSmw
aJBcV/DytL8WIx8DDbamyS2UEtkjexLpkoqpx+8ZOJsuClKBEWQcO0jMekLRHWR8iVCHghssGV1N
U3LeV6iw/jp39Dx6s7SCalBlYFZhGn05b4WEfWBJcTXgVXm3e9JZSOcMDMP/ierTVy/zD2XRdbIO
q1WAIoTptXTgQndBNAVGCNZpY3i8ofMIwcwsxKYPEDETRx9hBcCw5IC1FSyg+aHV4hAMXpy50u4E
JQH51G1CUrqfGmL5uc37X682biHjNLz14537iVcXjY3G+iN2d3w7pdtE8oSVvES4ck+Lq9o3siy6
G21Zi4OOVttGlr8Ol6uus2IJaDRuy0nPZ8EhZfFitYtrUuJ3ljinP9rG1Zo+2mc5aVBIy3RZLmsM
G3U2uHN3JoOBpm6kDaNDj3Xs5bFAWG8rpsAfOzAkiRnJXpDBQkMMmZaIfm+zgtvPBTfyLK6/5MmN
vdIqGs6Y+eArEFiVYAu4tvlkWsHA1Fjmt1LEP19KpFVgPQNIwlTAvRdc13z8+Y7sGtDI1GjZYo9+
I3ZFTzVBbDSnb8VvXLimCaw1B6SmJbVlP1VIKUZvqJTZHTTRn5Y25MmU2MQe7y3YKiomR+HTUUu0
9qKkb+cqGzafpLkH/XFt6vgM8gw9lHgAulKToZp7f1DT9u1cgayITy8jTGudO9ucIVoRtg7/X2t/
cXsqTrzcHt2eSx3qBtN3mdg79B0R2KU8d1Eb0oP1Uptxb7m1WaArkrHmR1y86d0Q4GsddkA6/r+O
iPQnv/0ofpumTHVYN9NpjpRogRCxnEjo6GWqedmHmh5hMWPJKdzuHwB3BDWKWZYW6La6yZa3Q5FP
csyY4fYezbHICsBQYciOWvl3EEZqCSbJv7MJFn0zDl0ejp6GQPg4qyMKjMkS8JCe7m+0ZOct++Th
EQjLEhxdziheWoYA/V1bCM3Vj8I6YlK1FDcmAepIcKB71C1tn9k2rfEAXi6C+QlBKMGTAkZ+b0UY
WTl2bhJgt6DiM8uIhxWuKFIeSrGA79GGDN1UD0do5U3O9vJm7sTiblQo0ucq0T2kv0ToyUwBQa52
s9T+H6l/cnbHXURv1pgmtFcB2QAWqYHdYRJo96tgcVzD5zHzCLwlN9oeKl1Op5L5hHzKDl8nKgrz
PiQ0f8s2AytYZkMy3gHS53y0Las3Q+HIVSM6zLXFrnyw1c1tLZ5WOGBEWnd7QDjYWWSnh5Ul6DEu
QB5cj33fTyZL4NEtfwqT4MD4lgOzj3HRwLu35UTIab+cdm51kenoGkTMR9cEclGlLPqK3PjhxDV2
sYUk7AcZ5G7lFLMIW2pfIzAFyBKhYbEH7X3MHzi8ziPYK6vXySmPfDNlBhLffXcht/FWItfFBvuC
Q4GE533x3XXQSA39f/+nxxQqAHeUO1unxzDxxfNfffETIfaPPL8LJHfynePUb9SCDQeBMqR7+lSc
YfD3O+mlrywMUfsGPwOOfZwJR3COozI51IXxk2KMJKHorYfF0TCp7ztav416sDCgL9gLqymALg+U
HlYDZSfmRV+t9W0Cihi4nbRW9rjEPYR202ukmvnpl1zCrSUrZ47pvq0XeSAEe5dJ7C4RzJUyLI9l
O+wueQkksaABM5hZwT9YDg1ijEmiEPrrB2cwJ/n9Do/zlJUMWduccbRHCRPsW0LhR4Mt3v8hO+Gi
euY6gal1aCP+XrTVKP1dpfBD5OJ4MfYi/scYkX44jjsNsV1CX4ngjBkJ9jDuKyUq1INHukRK1xO2
vUNssvl4Wi5bD9lZ+eWoDmwU6rTsFNdijRGxx+qIYfVl2OmYreHvOXxVOKRv0RUUuI7Lck71uc+9
6XE27PEcGe4akfjLDFljTyxctqO1hkTgtrA0ECHc5S5ATdT48uOEtmKcaOgdu0NpnfCA3vjiTnsR
tpWTWGYiDU32OowvE6DEIE28PSY/VNBwVpsGObOUm7/Z/i1Z2akj3SHDjKVfXCzgAI3gS+7WZXKi
PVQ8qzJuDfJmyXKBYTlhKvoFDh9TQMV+sOM6/JrKAFSBRLaAZ+j+KBS+eM/mzf7N8g7oBqCa8iWx
GCNLUYv7/FCu1SrrJiIbCG47CJd+1aONSzRuqn7RX+ZLPSjWa1z9pG/HRw2hls3DwYbY1oWagakn
qInDlUToDElpmpf65t1gQgT1xAoaAs8aBq+m2qmF8PvgKINDKdJUMl8+eYhpwEpEG9DZh8PkVZRG
blMSeVF52coqL28iByyjyXEzrCKnBPc0DqhgGBZ1mWaRtugnQjUBG0TOaQTmTar5b44dwHy5WusS
TE5/Lpd69xEHJEHnNEB1S0xnvtdBT4cb2XYB9XIu2rFxIMZ/N/mKvnlhW4mGGBzbITlGB7Bs044a
uOlWJe69C7kV7GR3g9XD7LtrlZAMfiiFUGEkblUbJpb3S+PWeer/E/2/hFUZvHzvfPkC36Jv6YYm
EW+Uu1DjIAqd259gbR45KLnIqPDEzJ08uMGSYy1+smzLd8lkfUw52ffv/aOAXls22iRpX8OQ7nCG
s10W9MsRJY/z5IHRxQQgare9K4I4qdOP32XhwvXTc8Us4Cd827TiYxg09ZC7Xg18iz1o++amVgEb
SFcqrWcniuo2Ejdd3tbQM5dR6loILLAvs++gZo3JuCDUvPLFRu88oLp7YPSspj/5aB3cQi0hDVBV
gqMfhViPVqEKq4fXRdZmnnnJbmtqcVH5vv9Ow4xDQm6JbMKC9Q11ELgVBG6eHh0aYDUKDYiIE6tC
+BVJCE1KUgmtgBA59TGQW/91WJ9KqZJmWdsGqRhi1audIh8ptaOTikrT8LYBhMsWLsHhSlwg4aYo
kHMVyj/v8v51urebkQ7Trj/MUGbgr0qUF7JTDCyh6Iz2a1csBhl0SVdJCEWDNzh5Rj6DGsP0w3bW
+6lQ/H5aQqKhBgsmVsLfApM05UVoV7Pu4n+pJpluz5RkwszA1FU0ICfTM/DQdQeYYIdZvvIjpVVY
X7aKOjM6gjyjSOkfROnU8FYDKbE7isZEUpORRutj1F2Z/1HVFF0aq19irXVYAXRzOMOS5136RTT2
vsQUho6IP613sxVTWL7IzftnhTJUEylGdiLDuciC8MPX99YUAc8ffLnn5iEGAFDEEVqMTKC9Bx1g
nzBYivef1ysEHil6b9KN1ehcmOPmZ1fnErH/VmJh7zVlykZCfbXGc+u4gInzKhUWqFKAdLgr/gPt
bevETICPq6qk+/vPogrG2DkPmpfOt24jBTbUtYu30BLOmzQt2Jrj6BEc5p8FhIuCiT8i8eQ2eev5
0NcFf6TqwanjXWegHdHJi7OStlbh774vExBepesSMqE7Zd5Q6Tt6IISo0WcHLeOvUO3kkJCsGlUi
2N+ma1KXpGuDVbzTrzt5rD+ugP4v6f6buxkITKlqrP9NM9gSapJl1UtJGlRvOW6tLqVEAdOJAgTN
XB5g6QUTMwnPx7jVm7hEGwu4zAiKf0GYn78EFS052iG1XivjM1nDgcNrgRIalYeWHndy/eSIxApT
su9WUMkMTSTQFb7wOAekldvNb5F7ZQxsiacde4urf7sG5DLIU1Bee9LXbvFVw9Y9yfZOpiFFrSJN
MmzmvEgqX5FHu05wy7GVUFO1MV/MaIxBvwWj0gjQieqs8r77q3ohqoXXD9VA8mP6YIVFsZ6DIu59
VA8ZtWI29EcE+rcenex+lduLFW4BSbKN9NUJv9PMAzmZim7ifBdtiWmYGBENSBi2tmpLBVS0qgFc
psa2o+IOiMQse7VnwFk8ckyrRGgFsy7UII2hC89OoscCgtiX2Yt/khJHlPXIr3OpZ89RAhdhCg4P
TBjLCbc2dE73F1Hri7LD9icIitMgstMqkiJEFsmDfTCm4kmOIkPV9KW026kNTDAyLLWY+FIVdMKD
vDH3E8ejWAAQTGZveqYjKqrRGofuWwFBpNfgLhyi04XnWeepNPbnmVJgAv+21hFgHieNTt8LXw0g
tzAXSZUpRYVkWLc3GRj8XXncPSUXM5MgIUcoVFzpjNwSNvgQLVq2VVhr6oEbjJzQFL81MuXBnppN
RUeuwnqD3eX/DFRoavByjft9X8wbX4uXpOSH5tGA+DoozE8gR36M4lz9etYMH0B+3OrAitV+ZWxq
rP2Fkmd6HwgNvBtwNyNQZs+UBGC+UZFQRR85ZU5oNsudiGLws0dGjOqb+/pn1NHtesxJToiybqOH
fiU2pM0XIilcSDx4l7kUpyOMINhb523Rw+TuihM6HBzIZuM8YvhuKl9HO9HPs4BTqSqL6SuhN6QP
N3BTLJXz5N8hMB53s7w/SVYPsDGNxL3f55sLiG5/gdGFUoHLSjgwv6jOq+YD+5se2UyzHjHj4MQw
/3q2AeW/rGm+eZmrWiLQAHA70nmLQ1uw1NlvEoP9QSAcVf+qGIzH0/wNuPgFq/ygj+3hUyeDE7h/
bzllo5m3yXlFPuJvMscwlLDW/zVbjyFeOLY7laSYZmlPqaxb4Hpnz4e76A1t9Eq43jHMTaK93FYN
p9Us3Qiuy0BArGVonhOnwciW77rvlm2I0gsZuUawjd2kz8t4ZqfmJXB7dSzPw8JzkpY/EqixKupy
18J0Sh+EhwTPUG44A54TwclDvBkiwiEMlqUeNK4TiYErik00+5JiTd0SdudSer9q17Ik1KnJ+t0n
gipyYHV7LenwGudHtpCr9wOD6oLdgGsjJLazek/Audb6r4mNaLMjSBoCZIxi05m/m0Rm8X5NLeFh
MjiuZx4KSB5Vt2u5FMAv6Da/8/s8Yh+DyxZUuMDR99z5IivABBKovpaQorV9kmL2iC+C7wr5D8yq
8GloVy0iAHVMZbzsiDq6m6cCaJyvQMQ/SnxF/eFzHUE3pb30We19SWRaC+seHl2FJc4lbFozj8t/
qSYpmhdTOse0lslS/iPO6oFd2P1kQU/YrGTX+Z2WunKdeWPZjUoBmrQ1EjQFhJKam6DvX+ZJkdWt
O2cYPlSrAsiVHb3HaFambdrCqib2UEZaL0rRMeaZUdt2m/gf9djGGIXnkyN6oI2vmoNXTWiTeuxt
8aXpq0GG5FX2BSUek85udUfp4Vw83T7x77n5JXsURrWqDZhWIORDS3BCF5LVi5J/duh8dlLpTbeo
xie5rbbKvYMX4Nf1Yrv+wUND9C3K4lvZbypJ8lwaKGhIiwAXbky4gYPU7ikFLOBjwmVmPRWFCo13
GgySSLLP2pQsV57kKbgsL85mtMK6/cKb7G5rmXZzpW+bQnL/hNfAJs+snMSKgkNCv0j2QWFJD8ck
OvWIcqXU3fB0pqwGdeOqt/tCa6HyefGzQYSaQX4/+FVGXpBq4uL6j6NGThNsgLRu8ty2Xbb/AcWZ
/kz/CyP6L+FMyvFUcTQO1VgX/e3qw5XM+LHSdnQkeCmowVYUi5bIkwvN5GH2IIj/yh+/+3jwi6ol
0UDbjsXxAxG76xYnPqx/xWwGMUGWSeKBSMo795GZh7xnIxmZldjG6thoM9EtXOkRqBdDh8EvBYZy
pAS1ygRKJY9/muF939BN6PW02iuXQCBzoILbDOIeE5b4RUzzkU2WkoxON3z2LZZ6ifKJtG4KsGT3
BPjNWrxcwyziNWXXJdEwufHsmh2R3vwP803CEMzGaRp5KADoD7XUkTcY+DFsidUYLEP+4wq9GV8D
plSt/U6YOXKopfvRWTUBAq40ueR0oFwH/7FGghOHHttcSsBe/KLMTCewm+cx0pGFvAmibyt73zjX
8vNazUzZ3q2yirO3GTXGh4GC/E+7WLxiGwHlAwdm2QhGERuC2lLI7o3jCrifM3c1re5ShLQHK7ym
xnClodSulnxFfG9q+nEBCa5SdjX7th0pKZFOGs1B7U08vlUnBZzz7ty4DOc3ogqtIvWSQ41s+Mnq
llveYmNTKPtyWBAR1tO68umhtmySIWeoW8/lfEH3Vz7ZxSPnkTSq19cCbziG5BS7cn/+uWG1lKfd
EJYohqSr5RBmbm085b+B7BfOHzGWlPERWubo3GrGtNX/xkIERBW/gbeQvauC5qRGNHRldR71by/T
ha7d9/yQlgPZXOEEL156xlYU6/7T2f54BEYNDvLHwiNpMGGIKxnxB9ELuBwkJJipRg5bTODdJGke
++gGJPF7nM1NEJUPbnIk5B1/TEg5bq0ClRZCSa5/VL42+1EatJZMj6jxwUuzcqDCxKrErdtRdNBL
y0FAX5sJi2PhoALwhkIBW3loSupcwcSQ43gOWEBH0vY1912KQvRminMkozU1TI8qFbJ2fp2Fkt34
wrYGZTh/5VHqaKWZcRjVDoWvGCeLlCqVinMZrSOvHais89XNNXTuX2p6/eLdTaUxGEPtzJc7yX1Q
T/umeV1sFcleSXNgaG6R8M5p7wvyZe9I5VLvsbuhkINGKw6/qPCsmKJrqXv+pCbzSNc0XIb460lQ
hKFfEqpO4SbbnjoVjBbmrm7yKStMV8DaKihPCIK85R1DrA8tAhpvKxjsbp847xw2Ai/9ggoYyj7h
38w6BhKrjx8JD2af22lpZ0sD95qR+4NjPjhH1V99rQKJ1ZZdJN6gSdTfzlThUXm3N0ihfO3l2izI
xR4AltoEoz9uqirMqJkAGfPwwgfYD7TuGI7nWZAHmb7buhH9vWw24Ea5QyM+rI0GY6qvxiEUYODT
34BeZLCgpPBlrB3EA4ODw7D8UdWHN85ot4p3jQuxGo1PADDHsdfNGagW4adyXrT3nI6Y5SH/HwOt
ylI0GjsNQSbCCDCl+6DGozLsm1kzAPQeNs7OCafvC7spJeyilgoZ8GIBQGUAHgokMIdOptiV5sTY
RShq2pyiEPxOXBC2NSA5omKAIdPdWcZRkbnh5P+G/CSE5FIo51tdyWY7/F5cS4Kq/RllEgbmn/2G
fofdPFvCYl+GhWpdm9kwZ0HH9BVcUJArNgAjnskO3bIupzB7P2gN/U3fRiIDNzvAvjxeCp+BfrSU
EQRQfr+qpUhQmfI1vZrBUidr6HYj9Y5tGjbL0csc2WjmsgPxTSX21r4BsrW5owKzsc5iNq8onC7Q
YNnCd1sVZiFQCBnITuyM7mDfT6YYB+MbaWCXQfc2om+ahg+THazKRvqlLVt/pF91pqJafBZMIYcI
c+lXzB8ogmRETp/moWovG92Q52Zkx3n2EgOmEhmjK+2V9elCIIkIK+hqpBrCevsfxWPfMf3k2K+o
f3vW1z/2pAdzdLZHAID27VtRTAu8X1uxqdWGaNa4JCRFQDUKjpmzNANoeNdhdTQKaf9lVYJlqIP5
TDThNszivUj4o12KwgG4ZuUW0QtkfHrZPhk+xuiwYSx8N+27pBqLiMPCb+dLY3MiQm28ymSI9QEB
NnItK4K67MGlXaLg1rCmkZ1E3krMJsMNs8ewj809VKwBkp98gaaz4SeXyzIccfl3+mk+au/UsSmu
yQ4asn3AjiArnxwDD3q3xMYjR3mTbs/WeKk/j13Pv255yYQ//DrQNymIRj5K0rCvJjZ/cZxqLsQF
vJfhjbTDamQV72LJUNKohvlmuW60Q8R1YvBTzM07yWPdlcFwDVjkZc25sQMeGD+rgeWqqf71ztu7
5RfBNwLnYdIWmQ/lzwbVmVwWoeawBCnvfCBsFzPW9V425zjFfQABuj1/uq1rOig+cEYJt1rJJP15
1ALq3QUTR6hoNbiYO+D4+sLPF0Mb4kjyv9u+DWjGf5yQ9rfSJr8o2mSSXoNMySxzxwMgTHcbXdyp
QwoQEY8+hbEZZ7Zs1JdbhUpGtnrn7JNXU69vZbkSQ/ivDfZSfiXfumABR13+VCSrifQgbD8Ldyz4
Gz95H0vzG/OZYQf8GJkxMbuMEOgBSe7o+OpmVxJThkJXUq+aOdF1//Z5GnCQG7w11CM/L5IAcswX
YaIbIS/3JCFapWHEPgq80KiJk2xp/+q4Lp9m3g2OUx2Lvq8vFVtWiGGyQtkVnFruEfs5Yo0NZCZf
iS1R6hEnqLmV2j5sXafurOVb3IZxfNxipz+2Skjkfr7qe1KJwpnXcUmdsq83ZYb0coFGxNJKnxGV
Bdc1mFBQqoMXxt0B0RmAXLJy1+BZx0xWBmGKryrx/MZ9mAftZUT7t2unNrVaDIYv+nnSKsI6xpti
aK6Ydy2a4DBh9uNDzOa8IKLf1nl7apR2oyAyothy8cgywJOuthk7/uj1v8s36LNZBz6tsottI0eQ
EE21gGNlI/BBKXNbANma428zB4e5Yj0tHC1B5OmuVt49/kj/6A+S8n7N9o//5mPNfTpLnxsBYsNv
2MMLDUkj4AGRNW+yDoOEm4t7XnnTUctwe32wm7fJBvflxXjB2fxDaksH5JzbyxAVzGAxOLRGs4yM
NVwhVRwatlBTvd1DjswA7SF2PkfnTmuTCYKKl6i7CbeeGxY0bBFuK2fYZ4LOjNudjIYL3vJ2ncDu
VUEZ1gzY3cjTkII0BDUv9zr2R+0CQrCtbLUL8y4XBB2o/wgGhmFUnKP7Aq/v7FnhdApxo0yzAwvL
n7AtwvtXB7gtjeqD74PHuVTrGoERZHXJFGdeKEkt2UtqbenByjHOfnHJQNAh97fJ6cP8fjI3qegk
8O3oWu12ZSjgGy0oVxnMUTItu+lRjgybLBywS4/jnXQRjc01rDzeQPfiBXiwOwXXAi5f9wa17ec7
aRdVMLRhJTqYNIbJPDb+R3aBmvNP6/eZqWg4snBaLYtlqSQVk0x/f7D3aIne1YeGC1PhNXrF7k+T
HUU4fAerLYA/Q0JUvAvWKCp7bli9riK4pb9SNwhTKwNQqX45CvJnT89Tj8Bn35P9LrOXjK6qp2m7
wGS9ub5F4VX9YFE4PMjxmSIMsGpGWcHA0Uq3cSVGvY1KjGOiwMxgFBRTcTUcr/tpE43cdb1djglf
3hzZFujCtkoExMXVh938nzroSea1ku80tomXtcgD1apIER9J1EgPPinnf7flCyRyU/sXwL88nL+/
C6YQfxDyuYw7/ITKTSvK6C2nqSHnxJE32hoWCjMmqACCLuJwavmv/GDefQomSXh7FO3/jTZXhDY5
cHi7ssJqlfgjMlhj9mvsL1JtWJ83KY4UxzfD6ZCcxCAeFFdhhZCil9s/Wre7RQd8Mt13rEJTpMTW
pIp/mjeyMR3A7BbBQkypNrXwMpHHAvq5WXRwohdte4ENTpXU389yrH9sGfRJiXfZtfjh+JvpP8a3
B63PwoZJwLUKGjvQOB76T8Q+sz9nIipMcgBcrdb7//VvhIyvC/se+DUPRIQwgNOF0z+UVJum/1F5
8/Px1LSiyyQ8jMpGX5qe3i2G2Xx9naoMk71EteUIElxQBu31Ml+ehz9b5Q+LLYB22qCXxDNZhsMq
Zdi9rAxJOZkLv4bKaE/ENBqtSyQTaMHZbOcFJlAqic6B5lDB3ToMFIHl/GohHO1RS2QLgfEKb79B
htfJJVuURY/2iQPzg110OUFkYcKVRL9wvWuOc2VPqTRN+FSmzDM+MIo/CEgZw47Hh2nt/BxKeDB6
regdAcJ8bFqQwqcDjOzOjNfomOHMOwq9Us+OnEkYvUx8jXQ2ot/BlI8mEhcRhrZHIHiHal2nN+Bv
LQxKdHt5kjyGT2EZi0cI3Tj8ZqJn+c7uXE1XccCjHRuYTdF8/RfN8C73YQuuGGLaSKZ4RortLt02
IyiWQJs9dynahQI9iVKgJZLaHGes3YFkyD8HzcdNhSl5StizmjY/7XfXQH658Ihs3wk+sQd3zEBD
v6EyF0QxmDdQzWOgUKecTJA4G8NklslSHheRE+EKQIQ8QwK/k7sm8Wc9X/htK4KyvLgcFOyt/+CJ
oIX0SIq4PXbDwxp0Q+RiIlLAzSESpgjam7KRiEFXcAy6lRLPtYp8EI9lMyEmehqL9dfL93TVtwnl
3flZSwWXsusWuwPdn2hTM32eMqOeHy2aVosI6JBRdL7fnRIGI2te7pCPDecf+vcRfFADghSt9XH9
tDzVQcHRv814n151g80sywZvWtV5OOYTMM12YFo4h96i1eWvuL/N3v6M3HQ49/AqRCr2qX0DNYJT
q30rTg77edE/xzspdXgqGDisIY1xu1oaEPLtechGid6/OHt1zZgV3iCfxcEm3iqFwlfh4WF+3P/X
MvpOvhYnc7WMSBR6hILz2lrk+gGfdY0Lpx4xt44mcRslHIzPKJTp9cwVFUOcgKy6fCbnn5K2Y9TV
GPjE3GncCcAbG9GOgXRvORgLhwU3JBuyY1s4tLTDaF1YHtyT61gaas+OBxeSKbhEodNkC68mEqH/
VNeJ4Lz6qEONdHW4aCLWg28vDHXcFQROIZxRtkqGq+lQIDAvzwkVFfdyVfMt7WHaoicupxqM1i5F
e4BfBKgMRMXMFmbotBn2zRBReMKdP/1/NaNQc+JEx5TbpkD7HFGkjMaspsYqcZppjKyjl2n0WCbZ
LZM/u2/Y5g3PtNhmDa9uC8KEBURtStH0XIotHo0Cl0AtHdoJwE85ov/hFIo6hcMfGF6AX/Je9hkn
HPD3MUnyFIrYE4wm6lI6YW2IHSTnl+aWd8qN/RPKRZa17r3WdOcwU6E2n91HFaNcLmE30iJF8RGv
Z06KQeH9hhHlQyN9T4zjTdcfU02EAZxhTF2kK19HiiBTv0zWKY3hJml8B8L3sV2rMKspFqcLiAhi
77w/OYO2fDiUY/kk/NQVOcz+f+xFUB0p94zYvipVeABtbGG+6UoDSzJIFJq8i/75nhmr0IXm3ZeC
mMzhNW0PzhZ/k+QL/h+POsAve5UTc4FDCh2oBHLpr0FjQxET1W9BHCvPaB8SzlUKK5ua5rtdw7X8
zXboKPubqkFSKEd5CPovT0DZIgaNjyQ5gaNKoyZMia4uqggDQW2y2jHyQ9dMst4Q3OnKFbghQwcu
FcKhRnNX5X89xjt7lZPZtXOefEliA4vN7avh50P4Sz37Jqw5IFNlWU9BjnRzN14hkNcecWjCa8y/
ZRnIFOEc3IVSYHwuFgz0FS45uinSf0zFp9o5u22jqBAxa0UZoajjIprpQp/wtAmDZj5s7t7jAWWP
jxjG4XWkegVvufHrCQNrn3WZz0VVmKmslgN4D7qriigT5hGqTw1ffyhvjMnTrF4AOKOczhdtN40p
YbQrJqQ1OMc98Y6uVYUEoHwjbZE/v73l4JuKqmAt6AZWLdCxZLflNssyM0OUbnJRx7EaiExxkk3z
D5s77LSpSWPS5NBykfR+c4n9BICcwwFSCpaa+LPBuZSYDMQ4WnmuS3GKTlYKuQxtN89OB7I7Aq71
89tvBIEiMNGWAN79ZwtOEmpkC0Afw0YstJjB188SKA6bM32JA4OQ/ikIPp+rWe0vE+qVCgFK3smH
ayXstocy81V7soNJdOlBNaAX518PnEnUSW8eJdcQ/4/oyKN6R3jQOOB2RJ7QlcWgCjiy8cbwi19C
KhYg8RL1CB2rm+OkSQT7IlRx8CXtgIzgnJk+lkzYTyLHbFj6d8CeSMZAY6EZ/CTsU6OZGm00zHtR
q6l6XrhWx+DS8QD8A6cM9hPcbLNNOmQxoeudy2oXAqhDewH+8Bar8acfH3+suRB46HFaiE1fAqp9
1NQ+lXoBjRoFnTPWgPGSIhaaWc8A6ZUZnz6hI2HZGXHs6ODWtr1UfugT/SyOwU66jYHecexC8ApX
DF0taAp3rL4vzVohxi1Iqm6GfvyJihJwX9QlmDezAToZNkVe5dI4oWYX3keJN3JnfV2Bo9PTVx99
r6wD2cNF8jyDd8bIwNb2tUAP+Q8b9L5/THyxoXPrQ8JIcUtfMHi3ijKWZPUbOYzeu9uOBqmpiiaB
D+sfKAWbeUIeeVeXmyuLjT84+/rfZzVszuF7yafdZzJUmY3uz9T6Wilxsjowd++hE2MpgnlfPDvD
muLt40XCDAg0pnzoleVD0WQgkpPmYUCSfQDExQVEDBrWidHOEFZPBBfZxtOREn0XCfJ9DZ1f2xTU
MfwoE3sRjLyO4T5Ja6vSYzE58imG5GfdHTbWyroxVU+tA+wFtP08R0hqP7M67EtXxgxGPkar1QND
Qibu7+rhgeBP3gQL5/Uoed2je9o9cvFZKvVr1eiUyqYUHCwid74M9+lwtmGzMradypJ9tqkNyFQQ
kf1sD0DKGUju83tDwo4hkZy47ZnbvNnVS9tcz5FFXjWEmCc13OiC1HYxC6FavWcgudT+cnHGiqsT
6I2Wf0YKmF+cMLjDCT6dWrU/kZ66Q0Z3txuGoJ1+cHzHieqsrGzEFF0ox1jbS/OPLVTNTOTs1vSm
hik/AxLajlYv2KbfiChDEYTU31YqmUnu1gApBPM/k4f5X7hKinQ5y6yMGgNZzji0XoBrdO2cVmPC
NKuIlAIGn4DwOYuFKRhtv7cAvmGTCDW7+UHpsIUBm/2rVKdv/xJlKqEu3cME7PbFlvQvXuhp0noh
39wp80iZbZNOcW7tWcMMJKhBDp6Wifmzo2qWRrAys03gaK+wQKLvN6CdTzZBFym6pmodlA68m2vP
QAzlRHro5sW3ZcL2fdDJMmfyzJSbFhCIU5wZWv27S9fK/oIiBlWwoRTbqt61hsaUJ5F+xQ181hvm
Aob8PkI7Ri2bBAlGrsC0a0mDFlcVmZ19EzQFmDrOPq5jyA3BB4PlCOGSBmEl9GqKySVdP4jSGf6r
wBiAKiS5ji+QTP9p2sPJDv6Cpv85bLf2WWVfmI2aEDI5VZ2DM42UAJOPgcZq4hYIKAaH71eJktTX
/syiQpljWKD89sYGEv2seut4ojoagMBHMEkJ8giBIvr8VMWg4WI/Gt44OuBLKt6kIBlYNKCc03Gu
lvKlqSbCmmpUzCUoqNv0Owyz3Ga0SL0SUhZz+FH4QfQi8MaPbW6W8f+lgiJHQL5xecVV4FU+Va45
dlIYFLG1wksJ358fRZ4wNJFA6p/c2lOL7/4VuB8CoC+Pe+oOdTlqs6puD5EuBxy1maDO4hJPd4dU
31Tpvdr0RAz/eUp/Ksgpdku6+KBIi/9A2XpI3aePfX0kE87srY6Ldy5Ccv0YIIlJaz3bRxexGhmo
4KaBOB99kra+9FCYbzAxHALxT/lJP2YY632KIlsgfXtKWrhX+Wi+SM1y+i3XWWmjQKE9znOAPSmz
lAu0DiTfK+xG007frvhFiojcXC3z27OcJvkbd6iTn/BFbYQ+dAspnSw+t6NjZDMS+td7j/KKEHGl
MQRLL/RLehWgURm+7WUUiwz6SS+xF0+lSpoLaQ/DHEaaIiCyRsS1QcP6lOTawieNlHuR38nCev5U
q3Mlo4atIAFgnNdcVw6FZgIKfoc3hpzul9lwlETOD72rSRLOD7w+Or3mEt6sNgQw3hMvOmv0B814
vyUn8PZza5vLQPkwQ8sYx0ncjJTexuQg/dLZtVMEimSzgEZdxi5CFnePT/bIkuBU2ANQcdVaDDbw
0my0bCgFsHKZDXiQNBAhVEU70BnR7X90LMl9MaRCSVMvlrwBxho8r69FIpnsn8uDqmhApadmhP3h
er3SWu1CLqghzbSMUb9rL0pPXdcRs3gb3Vuw3Mrx0zP+ELVrhzPG8dwUxSKi3NcajySEGe2jkMeG
6tZGXUwqxEOOg+eRW/Dh9YLkyTmdSLGC3EZFK6E3BogCP39tbz5guZC771JXuT8bIDdz7kr0cBh6
Qotx+GocnNUrDc1i3/F8uOXlgeMlSSuWaFitcA+5HKvgy1hSEdPoXmyi7t6IsWCA0QHkmRzgYvmo
TcKTLeqc/0aKJX4kA7cVK8GfvLmUFdMZb9Ut2EuwXKij4V/fFvDy/5bHDAXuRo1D395R6OhWmOzU
lhSNQIV2wcRkBjT8XHYhEtAtOTEN4x2YOqcXV5N6ol+jhW14sToEq9gZ+jMaA0vmVO2nWnVU8Cc1
My22lktGqsHH6JPvVlBWI0tgTfAzR0yZbAQKy3Pdsex9Sw5E+iyR6/UKPZ0tk/pfuqTrpigW9vhf
zSkF4BOpg/2ZnJwn1+D9K1nr3/wI3V9BfQ54FUxyzOhr8UXlVSvJe58C6MrNoDT7Ufqbo6NwplX5
BtZjfu46VeNM/RlzolvdJLbbGbqIZyEUll2QHEH+4i1OOWhM7MTSGeM4I4+bWS3uA7JEbZCGCli8
8Dj5woQUeOE+4HfxeskVLWjnMHM48h32YmE8Dg5lT9tIULzj5S+1AK848XWZucZ6P3XdeBOrWm2W
IUQ8Pcw0lkxRS/u0MADlAVILnByl7Vuu/TE1CSZe8u5uAqmKNGkYTT2XUmaMNwRCEs+slF5ti9n0
3023wf/UnMFRIvs0mBa0WbqmFkQrL14RFzN5OmJe08eOQmrhudUVz5gHLdkFgdA2u8R02JV71o1W
W/mu1xO4NkoMlpsLwhAr1nMlORt31i10akh4xE1x1z00NU2dNhTgKaUc73m/DWIXOixok51t9dsw
/pJtS1bkx4vpboZB5ThjcQYFmyfMgt6af+d9gnU5CoiMxmQOACngy9/Tf7AgB3uTc93dKQ321aNd
dBIzEAkIjHHSstWlFIItyALMlHejN9O1XLFMD/Z511BCr+nLlvyxsYXFl6JUT71zS0bRRp8KFMOn
kGelC9dE5XAPR4rgY3y7zmUBOcnVSQwDKSgQmNVZ0OTMtRyoOUoAKfA+tBOPEsjStdIQwnOp/BFQ
yCug0k0fl+QMJRNw2o6btYOgKg0aHZHPN4ZMTVDUpGavq32t9d6FjuX9mRYZAghcAV0iv6y6eo5X
3i/UPvffAH0a5Vu5VgD6UUZCVjfjp0VcgkhNdRVTjTElaqFCuYrjXIMSwcPOjjQz2IfHm04PRbUh
feZsVAHQnuEIcjXeZ1QYsenCqR8+zv6Jri7kmYIaLaAfC+XOz2Irq0q7H/N4S+WyBMGTLq/HyZqu
K+YHWgeB7F81+ZIMKLIQJJThNAj08f/epGF4Lckt1uz1WuIb4U/uklajyjB+fPvqrRVXQ/CSSUTP
PHNh7o4jEEvAkW1P9qejqbmr4PruPXMHWoSXHcOX65IgOr26nNhnRhgoH1y22iGj/SN5muFH4SJm
Z2KkJNWna7ssb3927M38oKWw+jLCq8LVPWtq2b0S3qlK+pe2JVlh0/7idPR/RnSxHv1+WpQb9hSA
qePAXjL/KIDNMeOzqTUnL5fzEHDtwdj7RJe7KW1it08WrZC+CzrLn8tdSj/DUPgO1Zq+VgoRL03V
ShE1ZExlKRvySrwc5Kz13HPxyD86WpuSNnPH62V4AIFq7VslaIAtbScjWLbnqXFmAvbG+03PyDFC
LCM34zuYG0LoLyPEvufzQAZDhRIBsLfScuAnJfIFq/kM/LNlDlOgtlyBoP+ppBLQmTPqSIrY/QHV
a1h99BSE6ox8tWUNsKZ9/FPa7ro+OPQhbpUsVG+2srICpCmiLk/k1lncOPEkkzENLhb7nWNskXmL
whS5p1mqJ5x+GObG3m6t+mofGoGbnBLeCliXkj9ktm+nUgR85Vi9Qk/p9XUpGcmgnSjxckya2gsb
WgsP3gigR6APwmIwsCLir+FRm/JJVOX71HE8ieTxelhT2R3kOND1VZJXXs4+7SlkE+7EzGcoUsUG
bFlqmA6jCn0i6HDnUKhuMp8vFsi6U5h1FvAKqOpfgWJXKvxZeWIqYpNSfBKVHJmQ1hHS7iv4txfo
O5AeCk9nnWp7mrrxURR7oHzvgnkeXS0PTPiKK5OeEPOjzLqpuelNkQHezRsFpq5qoeE4NhXtdEby
vJ3tdN2/hRFmUWMoV5d02uzCs26dgjDHAgJ09RVrz4zF5rn1W79BC5uSNkCQpDC1AuykSfTzHIL7
wom+Boj+E/S53O8lsMgowEO/8A1Q+QdfUYZ5pu1lo/ApvCnbys66QskxqksOWmDYB3uwXzWJjYgW
1Rntt8C/ahcXb95VOR8FQWwL/nKZPfcbRe9/E5wtuCjG7W6UtB6W6u64+4oYr7OS04OeEZYIEs9G
LMfK5mVepz86vY7xqV4aH8BS+Rq2hEwdFhBgCCXsXFY9d7fXa/RHwgDEX62NMhupZOvOw0mb1am/
EkcOju+mxWIkEhHEfoQwEM9cP5U/PpK8T23QtLDWtqpbEXbQ70Co4wPaW5433jQopu6+hptCTLQw
Mdlc/lG1kt5do2DX/xC6g2GjPdepvaDF8cBmHtQ+NGl9PV28grBimzLQjv82DILzmfY8Yt+RxePv
xxXl/otDczlk9MOwkP7AX6ACIbF0qbsdJC/+yH911WiMkJfqIPhZ61uAaK77RSx/03de9hqAf1b5
VTp/Lh43MIE1F01SrmjalZ0P0hWfKJSKJTFoGfQduOmYtyDoE+u7qRsBJNGKdnIl2WNkS2qyrrHk
lrQ/PBKjgjtsryViY7Udc1mmy7Zs69rOeDNtAVKIAFGp9DZsiCXezsn5db2TNk7LtS8e2Hx/gNgq
xYHU1rBwrWm1zI1AluKRPRaI+ZPOltbvAcbTaCBjk4a8y/EbaiE4rzHk0xzvyVZjiuCJpPGxLYm0
WFyJjPRrz2ho2qBm4dBXUo/4xRyI8U/l2R9CsWvjTAUYOyDJyRPAfvxTR14zFxSwiRK71jRrFjy7
u9P8hnFAYkAOg52FDpoddy2aHM+ZjzBRV4tXiNhv2i2kZVQLFELbg1zJ76mIpjUDDuMvjUAj3SF3
f+vDGo7ythH3UB/HH55OlN0l4ndCGXAfzz7C7beULVrX+PNRhwlQ0IVkwZf/7ATZKYbuw7IQPalj
IaxpKCFpquWCU6NIfNEheLiP/y2Yok+xi1mMHX+vG3jjZqekwddW/g3AYT0XtU/YdUCOSvUbbO/z
qjItMXD7rvu1nZqAtvVU1ivchaqNv6nwUEVcceUfrKZ7YtO5Ef3oz1C9G1Ui3FYGMMJIkR88SGHw
N6PewD0PPH+Rd/gqcd+Nusi9RLeX+KF6+G0QzB3uRO0KBBLzTb90cLnd6I0JKGQ7PmTkp2J2EkQu
Cymlbur9UtzZL1v+CP0ix6Pmro20LE6AfJCMCLgwIJHb0LblYb7++4YFZ9TT/6Gpyc5boprad2ZY
ELUS/HJKaZCDY0PnC8MJAkMLBYShW/Aw0ryBRyRONjFjptz0Lm+FOiUtgCKP/refsVJ+sLhp82ng
piyCrcbjipILTTAy+czNKICYaoYpufu7l+lihBAqKdvBga5Xp2nZIcP2lJBhTDaeqyxR8YDOKuHo
baQBJ6b4Vclp7FWvTLrG9fktrPjYo/I3w1k41vA4Kc8/Fw4G9l4vC7DmmdhXXhgUFA0s2VICnrkm
sIz+3LS5kz630x7oC5ONH17LSD1Ml2hLuHbfdo/yhfyXrO951xdB5t63dhoOU84mK1fVgg9bcYEd
gFZxZgwBKPcB4iaRjpDUUPuiCrdxMVaoV3G99s/onexaoCJDFEFtyDjLViWod/x5N4H+FdoHFR6D
ZFDjTSlxdcjjHn6RJT96uC4r7/GbQ7Bc8JuBwAzOcN17+gFhg/foLZhzc3iQ1WY0gtRe9bNboCsc
wSluegS4lVnusJRZckyw1LnILFttKRHKlp/NvE8phntbZwC/aOlBqTUe8hVGYgL2TehEEiC4Lv6+
wT/GBRFstD+XE8m4hrGWouZkHYIW30uEfq8527FATzY6vDSLjqs9EnoDxlrMd6fEg5T5LdyjWz12
MOGBbchYYMHBtScUtcqAAFiOS9Jyhk0wnNT5YZBezUZ70IkZzyEGGXHjLBIvyJRXDVmNz1aQam2v
KShnZuqreO+A02EpqJLcTcBcuL6X5ZFeoBcWZzn01m1t7qJuYjX47pX9qtmxTwIaM3gQC6Oo3cpZ
FOv341Nda66n7H4ZoP8ps4jWTEoKL3cZfSp1VNfVe63qBWCNdD0RyhoUeyuHl5xXCaw/KdvBB9Rt
LutNDJkK43F/CpwFAw8RdbJ3tsVliED7Gj/2f6sWo83j7WQQ2tw4/DJW8HQevgKCSbBOWH0bhC8/
0idnKa+v5t6I9kfFvLRgycH6rIy7Ht4tF1NC4NsoSlg1eadS0of4vnMmexFVmJzXNe2w2oiXYlAe
Aq1Z+sA6FE+p8zSarDnnONFui5GrfzZNUG+ZpvMtP+03Pf//kB/JqSDSpV8HKxA/PJfmhZ+pDz5+
g/rN4KP8t0QHE13yqpspASZrtGUVVTYLJaN4hjTssEeffWWfBviitGoBSBpaalUuYKg4Yap1bOQL
JdQEmyKmJBHD8lJSKLgiI0P0+AxcZe3Oa9iPqhyoDf9NPxwMEjbIHfg9sJreek4jH22uv1jfUKkc
BiG2VagYVtKvS7KbJ6IhTGAOO+x171j8rZUXVuLhj2XyQ/ET5Cn5f8QnYVxuK1nwOJB+GQmc/uMG
Wfl6vVsO9jynlexuG0I6w5EpOQYkngQhRmTx3GO0EO/jv6ZJzdfZlr8bUcFVmRudlfaZDmmW6qJe
NfE1sG28GI9A1iO8QIvw8SkCVHLsPiNmUp3t8cqCoqBrd3pYmkFKt41TSeeIgzEvgTVkr15n3gaZ
dNu0IM4yWKmYBBPIvq+Scxon7Zva0K9Hdt+VlbN/oKWeFsI9khBbpxuR7W5WSmqnQXWqnBwaXlPZ
kZkDDRFjZFFKgUu5106LaafKPJNlJBRVeq4SaHD1+ThK9sJFn+v/AQi3axSkqrGUnY+Shao9f88k
hgj6l7jRwoLftgJ/vuoJBJ08uLt6VW/vtvqeVI7fkkKRwMOXSjCQpOHU+EUUFM86iK8zBpaVtrvP
9jW7knGLrsPwbiFpgxVBjjvCBeMCnDtUcXI8eCWEhkcAP0LKZ8kpNHrzVIdLRHWybZJ3CWIQKr4c
IRw3pTWJgvz4NCS1aSxMWAp3xXUuN77LUg7T+ZARFn5h6qb/TY9knTjt52WToZo9gsHuv8glEmt3
GK+AYiWGWdglP4RA3M+mdNi9jL+Z+KbHmKU6xUcNeHT7aVZmdSCPICO9x2RyjjaniHGGNRtLK0Jn
Z3EUAixN0tEGEE1aPjikMpO68WfTepQH7mZBkOL0tIRQrHrPVYaVH0HztSvqISBx6+/MjSQc5XWy
vlP8rbDtOIqgfN493+KztsrXMi/rmxoQif55vLXq1IyRyTG7StBV0xsYQQZ8YBGF0Vc5Kq3vB+uK
8gu+SkdYehcR5rboEmEH1o4gPAYBZb2Fl+FVgms+eAP3GGUNwqmF0d2mrfGtTMlCOik+0d2u43uO
GA1hibs/bLC7Zax0bkUm9xvWI8HAoTBzli0FI8id+nzdfvhvtd2IO8uV7hXrcYboXiQc5WVZG0R4
7ih7ga/AVNRjz0bx/WM2NGHYeZvZDAL1fna+GGf3PdCoq1TCVSNEYPRjoOfW6YhRiEERKFdKAgiG
ODHgLnb4ApM5dh+KJzniUWbWgZsBSoS27wwkAYY3lXAHtMPkcFMiOns3z5kG2zPdhtznbvv1KMpM
sqpe5LUkdMq8olaCeUnAMFad9MaZSLQ3E9NdLHhKrwf9glW0P5D/j6OCJ+vwSXgHpAEcsm9jfSYW
EfQNycYgWlRBczOQGfIagXv5g0vF31/fX0l48XpL5bKGu47Lgqkkn8fUb4rtJihXOH72hdmWTtXA
pw89e7K7kTWpGjK4FJ4/W5zzWaEwHKFV4uSarvaKLzErodto2t/p8fK1UbKcpGXUltKgVrK16mYh
Wz3vRJcspcYGf88JtO9veEff/OgHJ1xCU7zrA0JOvGCzXHNR/jUMAsVMTq1Fs6c1vEIa6+Ju/Saz
5rUe3ITB10n0ifC651s4qkux6FCYHaE8gaMV6Px7V8qNI/kI4/Jrame6NPbIcOikiaOdEYX2sa15
RpbuhiW0+es+AOYgTovot/S7gZJTIxa4hl8V96xRitjxCEEnCZsGO7wNS+aZaOPvPmkHS/rPmxJX
22B/SMORCi3fP8X2LkmCyTwFGR82QNl5TUaqifnDc9436kYaOlsfHRjPVZpZpbks9CwN59htpXxe
FNrpqSclfMMWIR0BG3ur7JL05RGVO6YOX0dHsZRgPbO9ZjGP/JP+y883vzLZTHjMrdGoWrYtyJ8W
Qmtuy1E1fxiqgLLh4/e2VWTMHOdbtSkf/FQ7baNexJ/LnKBUzJj9p2jA0VRk62ugOIw1v5WZmAT1
09ceLwP5oubJmGKrQcaiI5AbUCMATeikqULhk+cHPnM5lcAb8iszYnH2PTArKRFc2XsJ9yEXOGq0
3t8RUD/ThaU7EjmYf1RrQ/AW7K6BXYGexWFVzFAf/UovXuRc/YTP1jnmscZDKr88l576PjwXQc93
mqm0FNOlOYccbHGMeiALlkY5r5gueXpCpvOlo2W6CISB9qh/4kBilDgjWAP2rc0GlK/lfLSZTKTY
euk4PYtGtlMXtBVZn5v8zVmYGB/Qn29abVajFwBcF5DHQFQDqu5eXq4OX4oJIjnmVDx7D0jhQtkQ
pJ+7qavNxIfAfZWr4gAQUx82iTakECSv6baA4M41A7S8xF2sFOizUfopOgWqD8Y2ip+FouexUPW3
73CcqnZENzyEpK08xbMocYBv9UrSO7SSwC5jNFtSR9aEr5hTLtRROboCJL5ffZzAaAla4C1Ad35E
E8VRAKQ1h13797i+x9BR/eSXM4KWXOBIZTYuKHqFOTAd1g17dVh90GJkLAdGVnqIBwZZe8OBHsw0
3cOnoHh6RXqgS75hv4bmFuX5oCZfADsmDYGckHoEvMc8VR2bk1SXHMD4WWiVKljMtAbkeJRNB34U
TKhsqK4CRscUhQ2dRmZz6pwD7JYoIZi9/+chPlElff2MeVtUWwlVu03QuZrv/qQEv6s2PBrbrv3u
36K1SwwfpaCj2PHTAeKOQ3rVpoSX3onX94DtIf0qcWjQoAuDvjaMskxsUDc6+qgx4gQisD8klIy+
a5tUXdrLdgC7TDdINOHqLtqDmBn00g2gDoYxg6EwBSrIOze3ia+9nR+UWcw4hhjPHPWVZZ3hlL6M
l4DecTgWyVVx4SpqDprcqpHJ55OV/OMj/2s9Mhp4T9fw5OsS2Qdq8vYz4F9IWXFpqU4EX1sJbcTa
LN1ozxbwp23f9UBwaTfEIs7Q8RAcw3qeiDhGD/JUQ0qo1V6iDylAtJqILaI6VGMMIiKW4wosoRQy
5oPEaP1Y+yRqrC7WK3pWGFWD6pAiVS2As3IsuDB2oF4gKbEDi6Qs5UwXr0u9dIoySFOds7Kic2Jl
HFOymCrTAc2g2PaSApNW8FSLscgDvQqEsbduqJFcu2jQVlaCTOKmCGzaiKSSbscbr74gNLV/kloY
iHNNBBmzwrgoI4wIbxTPWRGy8j8x/vA+Jd8oWiB+Er3yW7IBYJkyAGmbe3y51xuwGSizhvKW4o+1
9xTR22eMgo9GQbmW3j+WY0N/FNhOvfAGrdjyj/G/9UODXFZkn6bdA3VJzYdYjfo/9sLePVthQR/k
VeCBKpE6DholBsqHTGpO368m91lg+3PKOyEywgvpjdrPqQ6aZAxTMbg5S/wFacw3a6c5SxXY+yZw
vceDuGzv/99V64iGAlz+Ao28OO3boyRN6TfiY2xfViCR45weG9j7kQDT6mrUWcM2OvGp40HWoUAj
0dBN9twTPYeovqTKHorVWvoi+qcWD5WHQWII9jlGM/FwiOT6aB3jtxWf9pJRHn9musnC72RcvYmJ
tqvR0wvCI8UeyJKe2AcKwEYBKR8DdQdO5uFNn9LqeVzqCy9U4/EpsTyLcndlJEPEHJSJR9J7A2S/
HyA4UEZroyuLt8l4vBR9ULnC40x0p0GWuspAjqBZnm4YrvFPgc1tdoLTi1PpnYLEnVfm+mSm6mis
7l1yR6Hq5rJN2Iq0PXvUgr92+ItSWsKiawHJ2vBd46mKmRcO8V923FhtvnkttIuXq9IB7IEV897A
ROLwuoHIDQ7r/tmZYtDUKxwLeORmTztROl3OUwWpL5n8B98myQXbMnr4OzDIaIGWP5BscpyU67sQ
2tUvOQ4e6GTgxNn1PG0W6OIo9mdchNynB+wb5+NRyu8V/mpeWtNQwNlKwQBSicZGbjy08O3EICyw
eqN3cO6RlIHRsMd84vFw/neX786NjEZVqO9lTrB66av38b8onBglB8kxIrPisvmUbVWOD1Ny4VG9
TcpaVPFtxg5sfA7OOu3bsEep9CQWYJFAHBWodD4erhX2kb2Skzx33oTdhncj5YXiJ+go+3lNhQwf
F5GkAw36zkx/VuycWGyywshh77dLBditIQsL2UWiGngzghvjPT+/q1dZ2U0lskntS+d1ORpzqWxd
wS5Bv4R2hNkdMiFZKgY7GPoMfXTfN7cjOrvPVOFCYAtKq10acuiCHE5No/uDHkPs0UXJ5meg3m5a
C1ceO40OIEfWxrQLP+LyV7tnwJ7TKgLGvurHoSL6HLOmRzekKRqPxIc7l/mkfSFpmJ/kPEnae1JJ
oXRVRpRv/eVDD4ZQuSOzE1rXUH9VXEcZIbLy0BKQ/Sgel2VEaMd88E0NGAMMWkackyDmm3OcA1/4
hY8BwSMQlIZfyJEQ95LwES70PXrtwOEmX3mtO7RYZ7B9kQgpiwF2Aeux4tIcCexE9R/RJWjHU8lC
CtwPMD0HJDCd042jSzkgQbdehxCvY3fWEp9vy9CeEtvnW9nygFFof6SOWEH6gKUVTtQhyLFKBJ/U
cGEyabUaGs2C0TAnBt8Rf2FW9bQFvYIJ7MkGOd/OoB5sSpY2mNArtvR7PNnN00NSZJ2IQUwbWYYD
txfvb2q8BVmej3gRf+8f+7y/yOGX8f4ZTWEEgfxapog2biimfjVoY6Xh2FyXoLMUrECjbOar5Wth
lfjKHAGaXVMidEg1gy0tHjsMqSwi8Ri62oDGuf4RQozg1t280SUhlWZkaeIkUH/9SDLWd6kgSnqt
4DES4wrbubWBQ4IMGyrx42NXyJaPOYFtFg7ikt6wn3YWe9hqKqulwrO9sA1/+scgz3kJdVNPCqYp
+edTOIeNgGdndIq6CJj81oLsL7IKcC0j3X9yOcsthzpivKszyDQ+MR6c0sDMQE3HbTJZAcOT8A3A
Dk1Ra7MNSiLUDQmQLFbWlL76oXfixMpXIqyzH0EUibAaFTD2LGNb8wtqNM8p9h3mfEw3xCFhjuJV
QaRxnfqxljExCSbLc5g4yMaQvC1gHRk0+SOZo/Zzd6v1zNOmZzJDdB0WCg/M2ArdHYyLLyo8CG9J
wTXGvFgEY0Fqxahi31sJHJ8Gtqh/NTllJ5ebYeJfB8HF96CSv7p8p8DGnhb4F32pPwrBIYvV0YKE
ejRKLtXircii7vI1Qtt/l0aKH1rIq1Ju4DtaYQ+D9c1D1mbguaHvU5kgPPy2FrcVlQrypqhSQcWu
UTGeHZffVH6HD33CyVTOiRk9XB9W8RpFIHKNUVrxSDzd7aXidTCw3tEIwvw5UnjRkDuIiCU0JnK5
L/tq6ejvRMH6OYU4/L616b5aamiUELKz6JVG0gXiyKMbQOyLxGzc9Egmdqsom7vxmTVj8wL8yvUH
Xd1VGJSUJu/xHMBtcTjHoVUOZ5tnKkQLJuPzCtjWgPdrYCPa7cGVne6d1HqA4cgtjdgm5Mh7ayWG
4d2IlCxcm3Qc7R9uMguZa2Odn+y/N3Cngg68ELSIS+qzmnReBpw/aeNe6uj4kUppTD14PcBx+0mN
ZpBj/9d0FT0zkESRjdTiGW6J/pAAqssWaR3ty+/D/yWqCqBgsKyPoPXNXWj9bvxmFMDXux97MdxH
GqsZ5VTyZc6qcKzEXXLp7MJR0o+sWO8M0RNH/JpnWu+7Z8B+WEm16YXt8zIPyJqCdHHIrCsskVNh
RFuaVIgGvSjnBUH886e6QlMOB+i4mIhcPapudTPwvl4xrxcDd8lQwS+1TFlx2B5M59YYBaOe3+WU
8eRAqWVZpEI+eSb/iI2Z6v95tIC+arMRhdDm6abkxaZ4kj3zbGz9bA+3gKKy9YlSA+i0jd+xuDpK
s9gRltrvwctlLl1bDLeAb9QY3j41rz8jbWh3di6kKlLiVV3RCA19wQSgCsIwr9dXGU4VycKpxWr/
a5rZFdwkYEjHEOuF7WVXxPXR10VRaLOM9lRXsFPyoYAj1hxwTNMgfYax2+zxTywDTJxpMNFEeHBU
hDSF9A+Ypx56tmu1lntvVe413IvLF2j8/MxWFqmZOaVQSidwM72jyEu132WhSBtd0vX2aqfLd2j1
z0YP7obaspCXlc5B2TkoKCG6ONJyjvo4lr8uxqYUYOHUmZd0H1ovLZRaotm6C9K5T5bYPhKvD3B/
KEnaN6uPyG1FWZ2Uf9W76zPC2AkbsKbFWAFXG5teq881mEfZyzKsvXUyBD7Y66xsyKLbIM46AmQu
0qIcai+hQ2+aAhufsqtZULM5CAS/uzLk3EVKaJyMd3apamGxIradiA6LC05VZpQzexZcmWI/AIaz
xvuPIke8siSMmDYNobf/AXd8IZA4hD/xMTT5QZiaHV6geHZV/udjkTQLHcaktHm9MfF5RW7b2tLv
diFh9KVrLoDlOjGthg8HK3r5SA/W6ehyd3T/0fUhaVqqJ+uFsjWLhFkRbRuP1LmtqkY0HnHIombC
qseOS5acChdNi8ifWjwrVmOuZuM3m9snYdjPho/2w1G4p4WT+A6O8yE2+0m0HF9yidf8EMbnKy/b
b6CLysblju8bMGSvqH5Zg0ohz3+DcbQ42JvO9Jo9tkHd3k3CHsTIAmNMYb6C+RQcCUlpqTWAE2B7
sf8XPrZKvl8tke7+zGXTIaDj/MTAQ0Moj4uY6N6CaGfcPMbdTDvXpYn7UZm3ebwQqqEs7lQPtL21
XWEnbF9y/egBt1VPmiar4VMeyFZvVPcKDZOAoyQaK/GzZ7VPzqoHhybDKEl7GO1T2aPFK0nWp3+J
wvdAdcDsk6FlyB2vKzdnTd1zjbxHzJaGloelH+7GaXyHznqwhVa9E22uU6vUDAicXoJnE5Ojm460
ArTTN4mvDfx4CJiJm0OboB/y2IyoV1wFms8fST/nVUZ50yjaszROBlmgXTToSlrPZxMLZPZ11KSt
8vu2AtCrlVPitv+dgKsATrV4qBLisHUjilI/bQlKRtVRoAxe4pGWeQmvCNtQMUliNziOEcd2A74P
061BEKCOfhhAhj0uHd99butYi5TJpozUDdpLCMcblICqbFdGo5R/kyVO32dQQ31YPRkmRIykymYH
wPHvxV2VdYyuyWVmDnGo5ZtIak5VD85k7rLdyWkwq0n+cb6wg7z0/lMXFosW8v8i3uC6Ba8SrzEL
9caj1oSvrksKyDYeMMsBzPGuXJ9BZRlVq/1h+2E1N8QmtsY2ZhNc7BrPNqLHCjJWa6eet+apqAU6
t6L+OQx3dLK/BbCNqbRS4dXjwCJZKE6qP8T4cBjLy15PPjCUGdWkh///Wz0bfeQO3HPSi00iCyIZ
2NBx2OQx6wSXAq1G8TmdzlDK1NLO0mbDAW36lVUCRRLxA8z+yol1dJPNjrChNOOaS8K4wVqHEErZ
FbVVhT6XschGqrvsO/qHSedMNg9yPrOv0e4hJwjB67yPIuaSqyMbwRBFOEVVTRzpicCW8MPQyKyL
6cP7l+9hh78dZIZSbw/4MbPw3j/QfRzf7iQKTawi/UYM2jmmgUgKfX9OTvjGPP0Ckg/ao7IDZbJ2
lGo+BPlEm2wVz/MTEXEBtAp1yobuPugxo4B0K+HqMO3REAngZ/1sRk7WhqENITVAfhoI6LqAW8Pq
NPdW+/3Yt8zUb+XFGaA86G+BRB5ucQDIABYbpj7TOagtA8c88S6fXwm5TS2sc2rrIcenGF0lD/TM
mvB071IIoZuLMW2hxs6Vhg0ySYZIGEU3OFydIMNVnJ5mZVf0yZDA6kY3QT10dYp2wKKH92bb+b8e
oFWrHj0U+7i/iJV6QOmO/H1q0JN9g5Gaj5Wp6kq1DAcjuNMdARJ7bo/yqCsyCdW1UZuhhQLeqqaN
CrdXwjIfGMHfBPEmDc4WOqqky4eropvyIBMHUSlgriPqGbXNNuS5AYSL9uFFoAGJjNXNEYAPKNf9
A2ResNztG+VcQgV4UCYMEBqBwNUawlRxVoIW8Vn4GuK+TiBeD5IxL/8tVoLhnkl96XRrKD7y/2yQ
wphhsym4fSFSZtpGN+i4HUFmmZUzh2f+9H34E50Wlf1ZbCn+3ERHITiA43mA1yCqZV8Qg4IhbvFP
oC6L8DV4s5377Y4pPrrN/qkT5dRBE1uAGuFlFfQ9tQ6G4i1WLBSRl9wA3leiZCqpzslCo8ZGzCFH
kbn/BcLrowhgKEZKnJRm8KEyTpLXU0LyAcVke8mXjIzrU58gKBdZn9rIcE83A/R1VBTcQc+YYEV/
dVzd/YLR9LS5SO+cGd2EJkBTgx+ad9n4oUSnivNvvlbT6Iatni7IkE9eRhKFvd9gz6moDCxGN/Su
Nu+RwN5WAJF0VmIP/q5svWUrYAtWdrGOtsY/A3IpgG5SK5dYr4yaYVjUGBDJMJ2ptxxZyhRveaMm
THgUy3BxlMtEPj3RYuiAaIG5TCr/rA/MB+Sg3oDrtVBvf4TAvsvmlpKJjn1O+WqLRLOasbRtNaom
HALufcAwRygiW69991n2QlPCpXaJDhQbbKTobaHWJZTSIi7cKRDXAtmUDvsG2LcuaQH8KFt815cS
UQqvZvXLRdF7kvcpEBEgVD35HUT9RBnizHTHebzQPh8uGVIGMAhPO2gH52UzYlc6Y61Mpz1W8aBC
R+snetIa+MCgsWjjJ2brEG+TncD9drCX5tr2bXzhqmwvjXYBEi5/bOZ+xzS/EDJF6vO0XWymOy4j
DmTL2TepYdZhwzubo/f3NXakEj+vnR1kyiIwRiQqIPNzdzHuNlSmGytKNfhCW+eajgns1b9aCX5G
Q8lwQUHFPcofbZoh/omxdEKBXrDk4L0dlVj3tMODeOTddpXX/7T8X95DsKE+2P2Bhsa3qwwZcL5P
P9VE8RH1RJj0NerLg+HG+sVJ3kNGYsI92solNui4Hqbhcrq958fW8HsDpbdiAtAAsqZv9ynHQyBJ
iWIN1AabtSFNAwlwd/YGLs0DPt6IrmfOxjUXPsDdjjj5T53z8qXBKR7rhYgpjdY5k1/9vcWpAAsR
Mqy1dNhijPn9lifsaaTwvKQ6YKCz8l6XUiFiU55qHgQlFQZ42pM5XJqRyBWk5myFk9VRM15lLNJb
1VuwC1SbOkIooxojoUjYTNepQInL3sGKitQK+w4EmiNR0KxQTDFqzacJ+j44j9xb1ADG23mw/OCa
iprgZFNI+4jJdZryn1RO7O2k3vJm4D1EK2WsSLQrojTlmMeMLnhhDcOrpomq1plIKHLmhEBTDlxu
ZIVakHCVzO28tmsK7Ms5334hq5gBpFeopg1U2wzsDfsmM9HOuoUc4biZ0M2o5zZJnlP+znhq9JPg
+ZCPWK8Ya1taqX1nJylYnNdcp7iVMn2zSnlQcYW16zeJtb8/7RjuJevx0+SO3evD3nJXC9VcHWob
sDyIlN9aD/vt2+ABxHsVKl/u5RYdR64j76/9BtTj2gCQ/abVdy1WOnBk9MHRO8RsIv9SXcUjE+Dw
dwM7Abbr64K3H3XR+0846fuSl0USGjNVoReGnGoNQdx9oO9ETIUqOBh6DDHwDnPm77o24F5+6WBd
tfkrou0tVH0tOnyQphOHNhR6hN9E1FB8BCqPbwisFL2VuofKOw09C4++JuODKIjMeZJDX01NRTMA
VhGJArL30OMLntPnbsY51f9QS8JDOEY0OX1Fcm97D/Ssrs38ZAl03KPp/sQiEke7dkLquUFirDHr
QMicDuBCPQC8ZDb6FZ2Gvmo/O9iLBhwON8Akl3Mst87BoHenPOJ9QzOSyimHY0whgVOzV8tfrFIK
qaJ5p/jKk/SD2FQjay80jpzFnOA76xL6p4qgv68JpLX2umrgggW3nsaLkT3NLf4Ty56GkvzXN/M0
43M6tKxYhnFtCun+Y5VrqJvV3eg9tVNXXdb7Jk2BZS1efJRRrunuO0hdPBJPRdBQh9xlwQ24thHl
25nFdIDH10Gzi8z439aPdD6oFL0BsNnILG55yLrRzXa4JJEPskA7tgNz9gLzBfZ3z9iAUwjOHlXw
64YL+JYL4lF0so098LFTxbhMIta5Tfatxi7gpRAVa3xytPxpE1Yr1vEyL/cMIhzdqXRx3PR6uw7O
ql3hN8DFRvB+tm3Bt7f0mJ40qeFssStEPA51rwicPheshI74UkA2CLNzaLEM89DDeDH8UN+/gcno
W6x9zLQgpnmkQmu++IFBV+W3Uv2ay/H+5YLdM/ebkbHIhbVgmL2kdaeQdw4v0Y0Gx0PTdXpyswCY
+TNipzf+40emzfC0iDjszfldACzn9ywOma8kp4seBqNwYHjzVtGrwvqEQPpq4Esocksgt/xrGjzv
4xQXoz/zLEyTtgZh4xmlAk7che1HC9jO7x7cm/egoaJel+TeKBbSPNGvUaLS2obMADoFDm3O1BfG
DPx0H0DNGBqdOA+w1uaTG1kmcrx+Et1JdweZfUjNbFuwSIDr1UOfagBv3mFmZgfhdR8cMzG7u9E6
Ui5P1Luy7nSACiFX4YVeXatiA9I1JwkL4EGa6wbHwKYAJjtg+8nIA4CFiKspUlU89frLpoPyC31Z
+w4VGY5ZD29kIKGeMQ1JyV6vP6gjDt6HC3l/FsAEbT0HF6vBA7XlFMDdmiYw71IxIvf6Kv5szGBV
0zaDFW4TN/8vawCuJc2a1M2SLZ0P+DT66e3svQUoY8RlGx8PHApSpu7Jw2SZ0hrLL3WlDDNWWZaJ
88l6OI8mSMdGh+fRZJmfRScvW1PrIJ4aaRTT853ipfqDiVcDBbmtfoalqfLuRNebrfgsE44W4kBm
diJyJ0S4U5wxPzMBSnY2Yg+biHmKneMc4MSBeFv1B2C83lns+YtspjrfLF+/sOpnsUmxi6LbYZpA
6yaS5fqVXGlhRAGMANGaxBXW9oMWPmm8WP+w+gCV3fLw5fkGtLukycV17npm6sh3A3uWqxprC4ZG
encn3fjjKKwiDsOtsIT1a2lVEHB1t5OS/xwWJvsL33LwYg+hqcoKDy/+j5udJrY7oATyXlo4nbBt
Z4OXQaJinS0Ekk0M7qYvZtZudxQWRXleAS9wmIb2thqoV6M2Gjwck/9RKcKn7JS3GOC465VoPTCw
xT8fz/9NRb1ktOeGH3I5eRRCeMPKXibHOSBJWPLgejvvKinTNFyhuerZ/C2Uan3x8MJOL6oP1fPy
nqds9yYq8VRGUbG+YDhKP//hQZTlpt1l5IsexNNaKW+oDFJV5Uq28P2rhRu0Fekee0spCHkgczgN
M3wiH4DBXk1JLb9jx7JIbcemJFZx3tZf53rThDb3KWmW8D59Kncu24MsfH8QZ9iQpNo6ojocGSeE
Y0hXg4ubM1w3oOxgd9g+vBdJ9rDGxmdctf/TzXHid8MnT+vtPcXJY+y4/+ioJWvELUBQUKkjZv7W
6ldbGs45n98YZ9hIta1I6UoQbbLYasCkO8PzFAe0SKjuL4+fFGHmYgT5GyHJTs1pqofuNozp+1f4
cq79iK8lFZxM1vbatWawmfMEJKk+OA3SaLB5Fy2bzzSSXxY5+Bm20Tj+u3E40b/xNY7RQWjjj+vi
jI673RtRnjkCKIwjzI0djhE5JKT1o8E1O8HYTWuew3Ns/UXJd4MEee+QW2G93PShNrROk/lHAdV2
PTWoHkHSEa6/BYAM8C8CdfQaIUhkbsncWE3L908VwMSmGa4zvsN84F3N+ExswVO303HMkIDBdC8C
4vqOj9IUerfv4PnHu7SiijTttsdHcta2RWMGpHR+f9T9Rfp103K65wutV5H2PFVyKDX+iQtX3ays
5DA75BiB56HNwFaM7a3qdqrGXNCpyzfAT2TUKHpTxf++xggpEjojqoB9uylDMvfPT++j/K04WCZs
L+97SO1YNTTWFvsE47NsORPC0CeBxYTuKaTRk05CclC5Nppgb83VYV9if6a/mdtcTV1myIxmKNg9
eXX45HPsu7Qdqb7d8tzBgIRmujtWMyjL7aCoXaVkb9OeyyMFUCBq6dqGQ9/53kVSZevA4Uv/oOFP
gGgD2fX20Qsi+SmNg2NPZNgerM56vANv7Nc5XCyr55uF4fzd3kYkadHBXAWEtf2PYu+XiLfmodPu
NaZseHuzW9XKC+e/Adr210B1G+VIjmzLPOq0moNgT/N+g5sAHY6X63b9RJ5jUlc14+BGPzEOwgVE
lRtAHgAnTkVBeYE3JviTc/iqquGt7bppTpkvnk+GwsWs3vYSMSKNMAaaw14Z3KxXdz4/8T75KgkM
pk2U8eNTvMfaBS7uU+x7MWOBf7yYnEUlGFy34neUCvJla7qqDY6WGB4mMA4ntcQzWBm24BSBhRR9
bOGmvSKhpqFO43URZBqCyW7lUt40ZItSg3IW+0O4USaIacyzwB4HzmGCE28jflqnzjRe1V/u/AaH
4rKo1ALlFjUoZsz1aqPpHYYOAM7eCE2PRlg8oO8RKiQyqkwxHf1eytgQ+C4kOQNd3JyVEXYmzMBJ
AXewev5z8DYLIVu2IZP9mY10BKlOxjE7NBLvk+Mq2yOXC/zbjqQXjGeAOs+s4mzR4c4AbS62wuFi
1L1AyVjr1qTZu2N9fijCCtG2SdHxRgL0EC4B3JooDCO+7BnVORQamTTZFKk+KG3mTuGzL8CqkTZ5
JBHu1PaI/RessH4wZn+ndsbFKdTYbaupKf3YaAjV57oUPRosuerLSaF3MpsM/EKpXIXbbx7a3Wja
0R0ytouWqplK3cbsrPJ7+ewxSCYi1UcIrNFSAftt9LpUlhMEammzDWTwjsime5zEnnT8jojdDeDs
73kjaSYGrDiiiap7Be277Pt8kwI1I77Rq1ue42+H8leHnJK/LWg/LY8hs3C9F11qrIYZRcZ+TML6
GxeGstniBEbxalgJg1asR7M6Hegn7B199BzqlZsVLvhwW0exQ2YvXjiBUmuabkYTeAPNpNOz1onn
W+ORJHa55WlNJ3gruJnYNImR6YMPedSOi0ldXZKcRxU6HE8/0vF7YVG/mlcVGBOOFJUw4dHKqTTB
R79PVpH4xJh5JQ2Xsx3qYE/SQA5/Hj0modWEBrAc7OfQsMCc04ex4frdOS4a1PswddaYbl0/E1FE
ip/qZQ+iD42fraf7tMaFU5pKITM/Yih7GBb3tKhW6a6EWAseeqnVe1u+Rgtft0U4WbuIM/h96ang
AZIGEi9T/L+VB+g6jMNTaflCdkU2RaPduGaw5MsZJ7I7pIPck/4tZ06BGWd0OkEwyW/WkJsI6n+2
ddm2STfGPOGL3oBxSGeKsco/ZAm6wM5izfaw8QTP8frF5vtLBF61iQTANTSEvJq7Qah+vhGgYKG3
50vf9eDNxaGyFr57GB9NX9gyiBMgxn4HgNUjso1przzrjos9AjkUrgD79a/B4yXZoEVGeeQoJUgv
L4Y1HJixk84F5kZTND8wWDLJBocvIE6GnzoSfOWNiVMH0KeZy2pK6jSFZsDTG9AnDtgjuKD4xslh
uCF/IgmqDP168nWH5hdesBzZ6i9oVl07+OBJveXMHl9/A+MgBK2mtsg4p2bcPAxseirJphpyol4C
QCkIwKUcmKlozrgpo/XrVp/6TpEFRFq5PxLPq5a1eVvsKD71YSqzZUmAbG0R5w/WezQkuwWWg7ci
9n45u/gMl3EsgEUCsIS72lq4RmZs085/IyEgX/WXfZJ0HfaWIpAPOzL7mfkXepq85lf/vbjiAdTD
6VgCQL9FAmdn630yJ/J4fbI+fpShgO33zEQ1OnGlBUHTTPJGA7/2+QrQ2dAnQnehDbDUiKk17Uea
u+ocjvcYp9Ny7+2rs2tO3WgqJh9RHudrUw4qpqF2c6NMyankxdsUXD430RvydKxkKq0n/ThqXq5U
daAr+jwrDg+Y1tTlwrgaVpTcxZhrz1T5hgbgnDKCojkD4pz+SC8BjjC5mW1n+gCUqfCleibMI6jM
yEf5kMBA7MCtILaHahPdQcuy6QBXIojkEJpAjwb6GatfUjt9Q+Fg1dWSnclvz9UuEnRyRftMg05+
kXUbnuwok4yMDsNnCbwLg2Ham3zIMmmbOyNtKpzwJZlwqopopMemrw5mP3mt//f+1EAwnsUbjO41
dw6q3fFkOAZ+VcXNKpUc6PN56aP8UuQseU2CY6TTMJQsqU9+ui/q1J177za0zSNbeFUfuXH8etru
We3yK2dQdRhGcA+HLHd2D05HctRUXm9HCHgSeiTLd16iUYGrtfoKFAU4dGsQ07pjY4F6RcF+KP+z
QzZEFAXM7MKaZtGc+9OQ1472ak9JQKq89CfVaU7ggXxcb9/6M9PT10SVwgzxQ7Fy+UayyebXAHyP
WYRJDy6LYvP1zajlOArr0AhcbTbEeRfqg/oNas5klhZIOm+EMK+3j/4Jt0QyctbeAKNF4foLd+gH
mE5Lv8sTSOSIkMjQLQE1Vtlkz5MAUWYyXVsdLS3/4EKVW+FM+8tENfIH0SvVafk0s1lFlED1UZPM
VYUpEyNfzE6P3/ukVWO3fuvMHz+5HOvHu5+PM8rmSB58+YvAn5+LtnfKwiLOEUUFIjXdAF0Fxud1
VuhpNHMN4mHEKUBEi699Uvw5jC81tcD5ARvzRzbKd3sGJgXrjLZH7FZbVHaOOYf6gPCDB0rCeOFh
yiNio/2dEUduhf8wwPtu8UZSLwBSnCJ9yFTpFI7NcJ1tDfieVXrDNvVxXD7D43bGTV0tkci5CDVP
EiN2Gi1PXpvDNOrt7UYaMAbDRr3J2bg6i/q16SgS5EjATJd61d1hg4FIsgyW2uhH/0p85DgVhy3i
abC7F8gpNVnCnW3NwkkN8lYTxB4giP6foSF1p2y8DDJyKXit9V+0ZKfpK62fuuo2qxJKZeLdsQwI
4bORghCQJyhi77AQjnVo5DXafmFPeE6Vfo/MGhhi3bSxQRY6Y17eTJAdNlBPDWB+jlU6p3uHg2N9
WKrbwN+PmKZopNnqfdoXFxJ18ZFIeR4lrSgzgfq/6hFG2x3YKUVhWlU+32jij2v8wsu+KwukobOU
lKZe5Ai9Iu7SvAiPdm8gSaJOcXSdlDvrh8JKKHLHpZvOBPgUTkruWORMSnozuR2W3fKVRvgjgmgK
SQDp0Z9aUNdpt65f35muGNBNoLt6erCsz6/aVAOE66uWKv98k6w480bb82z6i8yzesXKSJNgfiFm
b+QVCnH3+6JybwAbAvERClc2bvnssMcPg5PsOqTuc3AGJVKxFRHL3swdmAHlar02FF9zxrsB7BFe
5k1q671nWB2/j55k75GnaxTKjkBSLDfU7xraXzL0T1PH8W4NFpk6tXz5qyr5o5ebYpym9nNL+5TA
ViRiiwwepGYGiFt1QBAqrrsmzm55kYWBKEEKOmkJrs4uiDoZ6No+4c+w28qtaKgEd9QmJm/RuaGk
TcHxOnTtz/xC7qURqC7EopfS2/gL63Sii3/EU5MD591vSOXkw3HtQr21hq2+BmRNmNLi0Clu8g21
506gxDXPFKFba/qfS98QG3xN+Ovm/Hq0P1HHAIdJNviCbZ3TdkdbBc+0leQl8A0kACu5o4ZV6r4Q
tebnqzrJIV5dRKxTOr0ZQwpcZWt8ho7g8VDLV6PGnIbNnooATD0XWmJUkanBwAGx737mpkjl6Ti0
FvPZuVjP0CUQzRedc+ezoY+EoH/tKsJwzOlqYqqkK/J1wM3wI5ogGm0sG96WLe2TE8OuB4vyneqe
QLRMG61ckKF0dfIHXGTybVLTG2Ki4KjbUn7ROWmwAY2jLDei4+4utttUtA9U1fqioWgUtOIHsXQj
lzF4jtLWA3kbRhPoW6Aulh6J7p1g+T5B/67MMZ2xuUPRVWO2WxyLu9pKi+8QdmtTzbfwHbg46UrT
dHsXmrfkCWaGa3ZZXYDvJDM/AYNeZFyFJmAx0/8HypUHoAvlQwRF1+Cvx9N6TQBdV39MJxUDcsSm
MGjZRpob0BLNj9VgImyUo4Q3+gjujx7+S1iOmMMCmJwRUChkQD8cQo7TPARC4aqRxMr6O4SkBVhd
Ra1BJK/+iysCsw0aUx8ph6Ytsc6npLFURLOLwh93o7jK/ju58xTS1/yU/dV0HLYVKX4efiCKQIOW
dqDJBTbJq8t6SzVjw+0lDPQyTE25liH4bEqmx4PrC15NNif3hi5C7+dUdYKz36EdsALw6reoYsCd
kAocjqkNSRT0M7Z7pJgncSBixSS6xAUSLA/JI+4e5T5KuVJs4ZNkj5iP1rMmizhGOlNmRExA3DeV
a0uYLxDQDpCzYdlrCeOlesgw2athgmyySMapAtEQQfmt/nNXZ2mSIAOGeiGVp8QSY6lGKrqyTs5j
MsNnhdpNOvTQD7zzXob05yGLM1SxclEaJuP3tWYMKG5m+rfSli0Ypco1WtkVXBMDfuB8fM7oUKVV
dSn7W9ceiqc6nIVPT4+aOECXQR4OcZRO8bVG/DvCRV8FCXeHSTBWz+QJjPicHSU7FvxG/Z8KYFUi
wIajNHjmE5U69BaZIbeTxZKW6xwx0HAPIBCQKdeeTJlBocGqqs4sjjecC1wgRFnyyXZGb/HOQABU
D0kz/HXUM1Qa5Kw/G7BVzuSFKdkTsFakK/A48ImPAkw+LYHHGEbuPqYTs/HsC//2VsreoxBRii7i
A74XD8v5yUPnrALHY0vjRuuhLw84ghNk4YQkwH8zOCZxZ+rQsZ8YRpwF/ZBUCrHmIbnxGBO5CXTW
QS9hHfU5kIEQfccoze4SEJhQJ46HuN5SXkRt6UIUvNhIvveDWv4Uiji4o1uF6/7QPAGmEc4c7c6J
KMW2Hz8FU/AbHv39HF7iAb4RDphHhRfNtLrEKVg7syjptFXLBVYaosqXDUAhad7U3CNaCCAiWQkj
CM9NSTuTu7fDfHXIxNP/qi7NnpujWOc9Q+lXmQ/98j00ma5LLo5YaCbkPtlykJclYKFJLuI13BFQ
Gc6m87DBR/f5I+FUdw0QkglVY9YJbJizDUcu3QOT64fV6R0Ngna8OLtktaSOXEQNJv+vPye/wwjH
lKCwye1zd62Nb6YndsLpPaeNWx9ankbPpXyK7u4LFOMdqRoZpt1mOhbeBPBBTH8NQ3GFkcUaikZC
JPaNYLVy2kTWH2OyBVsDU3RHyz/XwrZ2f1Zip/0anS4jq+Ztl2NLkRBr4jBjTOE3bR+8wQJmsqLg
10y4KtduTeI31RQ6tHtEhLTnPEE3fnSN+GnsQndw+smh1kgz8gMFxvzNuBJjpNzaZakdG1fm3C7+
WtCxrNJsChT9TvHEbwbXee0GAJpBUv1k16l/lir+sAIplgeBMUMwnGk7dRVRfVxnvqXs5R8yjShi
rdBRP+RjbxHPKo/P6fTJNHlRoMsZqumyJiuh5GrDcWdHtHg+U9bSd612QlZEFEVSQGJzIz11LUsl
V1k8h1xj0X4MFOZfmbJ501yqOXgHYTgrF1gmb2RQwWydq9BMoQ+onfwJCzkR3vK3fTVsGGdDosUy
O3E1qsdkdwrFyRJvy4/NW7IK/fLpKK+8FVlHfByljO5tyqxvvQFWW9k1T5e80AKutj/2RfV/r7TX
6ACwoYVBQKpgBrMm1/8tkei0mpGsdhyprJJiD5K8ptVmLi47OdDgu1qi1uJWd/Z++3ItTCZ4twJM
AQzY8lrVF2Cc4qxXWGYtfopjgdIFIO2lwnSJvzeRQPeffqOu7b49z+WfwqOIf9ceyvhgV4LsRjvD
pD+BrnhVeiyWY/YrCnXhmOeWPGZavdJ6Zq11Q23vNTf3PSh7Mm+cpTFuevShUOLk26C3lq6C6UBV
UfsfF+RXx5Qa8NanvM+gWJXOyTN29bXX3XZxWt7qlXw8rVWd37DYzfAX0CIH+yqmhkuMbkqJG5j+
+SLyj3Uu3Pwj5/z2MzTyExdQVJYcI/oSSDmWptFtF+SxBk9iNOmQF/dYuNfUv46hdBYx5AI/iTGI
7CEwFYOYwIENOYdtkS7hd+RgexzlM4sOCmlg6VNPKRNR1MB0XLkhQgtFa1gPWcaq3Y2lGVK1rSnL
Go6tV/hun0gKqpbydtD5BsVEthnfA1XgCxDBGjX2k2CxKlWj1CUXSdGyLrLaYdE0EVJO8yxp+DLQ
3t+S8CLMOgiOT6CxDMOB10oTKPaX3P3K9ZOsF1ENA7LQdxq1OrWnwcYYKBanISLI02uJCgv9n41Q
HnA84mk8iJCWSUd75zWi+64c6WUkW8yN/BghFLzdA499XQVjE+ulWB1SDCPz6GiDfeWZINSg7Ae/
iF9kjlj4bMEh2t1sEuQeMVDhX8gTGi/lxHaFRux8YL6BinHwOs3AkRChlmMLo9LcjjUnanDrzB6Z
xVvJpcjzwt1TEp06d0Ho75L0js8wEfSHUTvosb54sGjU9F79zxXhOXgswFVu1/mJGeF8NrZFD9xV
nKPCRIhWEQaonURO3kjVm9bNsMcerMC5qb5SMy6F5LQiCDja5ZU+ka1WGqiuw5hBhKY2DHPKRzhR
BuBKvlu0M1rDn8I351ZKGasSAulhE/8A4Adm2SELcvCvnnw0jEV7a+roEkyu8mSSbMWTpPK2j21z
11HoPT67FXihMXCxbH6nPtNknjNAWtekE2R07NHQU8lFlrseAhqJklvTYpLbXUKWLE6ESH+Xrb+o
c4bzkDoKpqe6Pira6DDctRGPOQF+675pst9XfZearyObSZ3MsJmIAjVUW+Vv4AqvMzZmud0zkYug
gmR2JiM/RlHNIKONm07CBmwvQhn+B0fPrS+ob8Qw3M3dO4tSm9dPrTTloOHItUWFnfbE/UKIw8lS
ubKjjE9rfDrvINdNP3jLwyfjR9eAyvc/q8avniDiTtoHY3dOc5ibBvCMS1h+4HsVDTGDY5T0FHg+
qwawrpzlJjzuAC5CEBQg1fnp0fgs51eEkbPQmtjo0KHnwsFtBWcgbmTH1hTOslUdNv2la+QIHlDN
XNYdxznNxpD0D0z7u/Uz2IGOVi5Bmfdm3kXrk0fYlAlAiF1eHxO24RTsf6RIvBYuYmj6DCMdvIQS
wuDFaSDp0vG0N3eClc7/AKpschyZs66sorcC6ziwKgNqzVRnzcZ17e3LJru2McylwRO4F9cl+r55
eTDDhnZVjVU0/dqrV3joB4ouJos6eBI/jkaWKXjWccvnRTycyZVsmsSq4saQspaSZqed/sHBU/mT
sPUDZ+vHPgSMR+42J/4+AjKzOtFdkZ7O0/TtrwBCWbXyZyHGmhgvmt6Zl92CiftMt1yGfpeceFOj
jGkc5lFRkwQewEyQ+N1IZV3uXKrdWDbmH2k9yzEHP0ko2k7ustlkaelT1e4tGf7zYpNDKE6K0uG6
qozc12k/DgrScWeeAJ0jDkxN2+nCpe4g0fc98cpAwSPtyxWsvO7hPwL1Th9Bo/252NvqbbbkSKrb
zejl1Y/mYBGcuc3/V6V4GIkqg4Z+MoC96Wrp49gIx2GoNxAzMT5RzUEtCKyB2UIgT0YATiUBq9bD
56LXSrJRFr8USdtCn2oYYm7+pUq/yf4X1O++B5LZrmwjqhdLhLdj1LEhKwytUJiOGplMSOMoogOB
oh0sOfWzR7v/zifSoWKphUyczElq2iTHjmHioM2oXvqz9s8zF+OlD2winJ8E+ATFX6MAEN8Qte1N
XGo3jTf/g3ZFeDvXhMwYD6Z6T+g0jkUcvn0oYHKqmMl6cW7Kf1vDtHPb0wS+Fzae7GY29oI23bM7
q/UpCjRxcLDwZ+cb1jfcvPV1dl+r/PIPhKb2opxiFajwLaq4hrylthUOoIMjiHr28GKprMDhgk6H
1dKHTaMk1QA2sGvYdnCMC0mKs2vk0peanUcNS8I4M/IAPaPBozUph2OaVqegpNF+rnVeMWcbEoQE
S9TZ28hQw0WPsHgFDHMBXaTnog7c85SVT/LwxjUkNNN7zpxUTXk9yzCju9+Vg6+A7vWKP0uHMqwc
ZJ07pyq0q19LA18dbOLPkFK2yFDmQFO4VXyVVSOSXQwK1d7hdUFhZQKXPibIqOvzoN5iru56g1M+
IRlPoLiZIwIHpBqvsRiUz+kxegaJ1XjK6PjcY15Z9ZWSWH8U2pfa5Mkqlkoq3SYAUKfGbI62LRUf
HxlBJcu3np8H+X/XJiq4vvx+u4b5uK/ZhHS7E8dFuDTaNSIYT90c3CT8TvZhrzwLT+OFiRZfZ7uw
2rNsa6V4jqXMwZn8e6vs8LyqFvj37Zs8QsKgs5FXexyCj2qA6B7B1EJ4Qnpg0w2ydIGPKzG8SwLP
Y/FwU/xl7B1aTDXt3ABhK4CCoYu/9kVCI9U+eqqIlT1lSCl9C/9/JgTTnKOgF7QNcwrpQHpo03mL
9lH3LwUUmprXI02U0rX9XumS7ctruIhDIrHA27JFp6okrUsgnoPvk98TjnWQlFk0NfS55hZC2I18
Ii+rH63dFk6FD6pww3WHO8drWzYdQPiI9rzo8MqoqwAIa5EANg9z9Ixiwfkvg6wCoMJTzH3aaLBm
azX48inPyQVxawPKGHpJrHNyEKbSTlQhaF69jYVuwkckyMdqu7qKVP7QoAQbnKsvi0p8o4d2UxQX
YAP8YXpQS+8nF1flyOabj0FWLALBLq/fPZa80we7iazbXJaIcqgg0P4KUYSvuRzHN3wonWAaPeQd
rBpGqiwkCgql4bCaA4xybZA3nKz3fqc0MrZ5G9z1Pq1Do2pxrb56EPNGxJDnxSu8X21aGJ51pVNT
rPdv3D9At2/yeohZDEpEMl5lsdeMauODqU3jaP6tU9O7+UENFXxmHUYmEcSyDifUvZxvzneCbgaP
yWdwSgGiCdkmlWdm1czkfGTaMYajcoH/nhRQo44wEeh/5WY8xDWAfEkbDOIRm0Olb5EX2Cgsd8ZM
tyPR0Qjjnszc+ICDzpkwRijT14W6V3CVtlC5iGNry9UKZ2osY8PAmj02152t2mvwB24nQy05zuNo
l84kLhbV5/p8Nft3+T2wup1RMBnFJSSdZy0grCuuJFrWa1NIWW/Y+VLA9D4BZ6eUgojHMjbN9y2A
fKTgLLh8HFnuPVAyFovC20P9aMHzpqZHJWZqdpy9+e9LSf0qLeOx4LlSq1nSIREZ8upGYGPmAuBc
21x4+w0W7SC/MdVMI2VgDWxZMuw2fO0hKnONmjdgohPQOCb40WgclNjf5srwPgSlCT4B7+1+AcHJ
ZuEu8ANXp+qPMjVoVKPMUKRh2Z8PVH8i/hkvOXp0PerdiwajjvNj5Iecxc7fHGZlEDuWzvadckTF
ORyiaXLcKImfXrTxV4l3su6zIcbY9aRSXoo8iHKpON5gKldC0R7hBZh6aYLeGgQTPeb4mttlKyPe
b28FhS7xTciapixiefi4PAOv4FTQp8wUqTfN28ebzlndGH8o81Dqita+8YV1+/1X7EgA6MdN5uUv
tBPiZCrtgVANjRSGeyOCz16xO4ktPEc28CZFy7zZrcYZ7on5uArn0lIF/lN1hOcQuM0p3EyZhvNm
CYec2hpqJRfXDlk2AQbCqv3vDCWqukQEJ0QvjBS2n5z9DH5bxrMtE2C2nk2FtaEKEVFX5U0br36M
FVrW7b1jLuLMtD6bpGVmIOpnojNNL+pNaHR72FZFFejO4rzgy8GlRTNOja73Ljdw1gj5sGtjzgHW
PO5gmL5wh3W8hcC5JZ592NDX0CMnvUkB6FWf1g9XfGHsf8DCsQ355WnTeYP4qo+dTPP6ga40KAak
0sYpxKamyYgH+Ya8MYJbQo6k2A3ZMbH6QbbcfCLWnrbpTnx7kHoL1GzqHPRrTh8gdvzcVdMGlOLi
Mi0WuHtYT+OMdS8I9h3wyRqyBQf7TvgoOJB/BMLAjf89CfdQ5cGRIj3TSJrFdsN9Chq7uIWfTS6O
BdLHQ6Lc9hpdAdYlEqZmqbMCXW2Ok9sJOAkygIZVvc+1IZ0uR2mW+OM9tg2m9hdNVqeF5nrW/n8Q
A/RZihBaXZ5n40k7X/WeKPQvFNCDInVf4I8K1G4AvwbDBBaF9W64K+VqXhX+YgXAR+yVEauDSk0x
+hvy0yzSQtJE108oaFRxRR/nGo9dsS8yA9NRdPNxy0fuEVLU1ifMhYR4obRiowxIFgHhgSo18wKT
/JNotrFF4u9rFlUZE83I5fHkHbmWRvJFXhGB0EEGFPu1co0pZD5/71DCkMvdG0uHi3m4WiZBS/0T
ST5A/eL37MVt36mgtmOpnNS41qNE94MmUHKh0Qki9wqxRXWimBEhNfwojwa1KMjuzeTjwP34pNey
n4sQOgeEhJNoGGDAvLMsQ6M9TZpnwC15LcOws3NKBmYnXipieGR6DYfhnte66FMjmYExE/lCNuDq
wPqhYOzA/bw1Pn1CmBalxtW8AJaVw1pLzULSATkTZTvJzP54SrzzqaWHcUWEpJiNCxK/f2eCe5xc
+BIBT9j66SKMY8ONG4DoQdmk6m9W6MREmG7QcJPWDE6JATrMkFfttO46Qzev3Dj9pnzRfUDpFUIR
M6sdlNIrLsw5XkAfTVCgvR2ubynYc2soBW3FKZGZfvv1+aFMiySCgQXaT5JJ+yrKrw0esBU8HhVb
SsEaXv2jYs6QE0psaEmoV1B+4DYqXpqBRAMc3noW7haVIC1b/uQbjCW/32mtm/3jEz+wYpU40/Pj
0ov7cohzQvgbIqHRBtXUZKkMRqLBALyRmrEpltnzesS1J13YVGBy4Ho02sL+PEYj9Y3ZiID96i1x
ljgtlLc3bkhCyxndqNeSKCtJSDCXUJW4rUCEKoVSOT5/jRW0XfT3YcG5OgfgJXG7CimKphrh2NqA
3hz9EA8D/QSuYB3Avjvc3zMZYQccagJyZ6QAqcNAMCGqv8P/lCL/hWqOmE9JkGc6VFyqXGxGG5+9
H0DVF6Ml7PVk2RdpDfIdhH6vWJS14QyERA2AmW6tRCtEx+7OW1XgA4cSCqtZPkXy2Wd2FEmF8+mQ
FN0l3EO+n3JcDEHoYufeXBU9yHxYZJ/ndsgIU4Pl1v/zcf8qaUpPCsLIwxoxWNiKkisJcE/E0jqR
xp+T3X0Ee3H6T/jWMFiPIydl8NnaVQ4grgp7NqpyVK+w5czCLKon5nr05U7qfvDwwh8u0qoHoMWL
6hIW3xTK0n2W5jbkrVj4gnY68OTrbYP0QAl5Ztg4ga181z58K3dpPqtqrcTOJhnQAiUkYIohH95F
rLJ+VqJ/nSJJKNR9bdut7ZOkvNU7vOTmVRwrV24AHfvG08wLcqdOmmPKG3roAhUg/wMIFVFox7Pr
LP6t1CS4rVRZg0WCYm4PqXgbbZmu6tpuqq/CTgXFpYAgS7Qp065AD5R/tajyxRMuMmnFwATT7VFY
kqWjA35hZQD2jT6lkW51ayswriP5JtT85Av2ZWcyMAUHT8XVm1groeDTj302OEYlcJh/hnHHEWWe
og9fYKj00Caf91C+hny7tym2lPyDwjo6C9Rm26wmqrU86tBJDsVWD91JfMod7+uPWuMfDNMMkWo8
9xEUd5crbUf6WA7ETdP9lCIpWtYms1dsAUb+N/fc5DpmZ+ynNlsPWyBlOTOvsFbZa5UaFQmkwtPW
cPz25JzDq/zvgLb6JWYc2r23zpYK4xeVkMV8ps+N4zlgQpaHsbP+qtXy9BBE+18utsJ+mLXUQoM9
8VfPlDPqTpw5qU+vtng6VpVH4Zl0XuksCt3wwwZXQ+o9D14XV8wnCmZuKyjRwhX66ugsjNrtemN/
2twMJw2K1M1eWYDF0llheYjAqMOGWN9u+yZXyBvmuc97JHiWz4oiuZYu7ssF2qETUC77P5+5rC0L
tpMS8ZMItXCLzSzAQY8Ts4JY1XrZE4sJzSfHiAbJYT2ubow3ZFUj1fM0brSMopxuezxs03ktRo6J
nSI4GH2N9fwi0pO9Qy3TVOBsoCnHdPbC0o/Pf7sWiL41EYUm2PEO63QOGhXSGCmmJa3pQXGWA2/D
kKEt/UDDi+q13vjYYSD/4Iq4WD5d++3ynAOPojmGSvAnPZ8Duyl85O/SANnoAgcT2C0v+JcOw3HP
N28pEWDywRToKFaVQXBiqFOEoASXyRBj/xmqYgJXemEpurGoM9jDr1o3f6O4zC3amGTMuY4gGGo9
vcTWu6re2+ZOGYdBsNgSwfTDRCSyubwetD4l+Zk6LKwUdKsasXGJ6JLAMaV/1e6Ai5O1RcxiuQBS
Q7/XV2dPRFMRUGgBAIrQ5+1SvfzMw6cw97S2nPq7dooD3iG3jkEwzAw9Z/t57klTuTPtISbPAJfZ
Ga4fumC6QhwiJ7aXM5Zbnzyto/NvAxnXxcHflHJn7/ntfclRf9C4yG5cha5ypFN64F043fr2hFTO
eFV1vMQl0G3xG7xWZmpEzRD8wsR38r7dSfjxxCjJ4/C8HMRkfPuq8k3XdcbWWbh7jcsTS/hvtXm0
Mq8ymAscbP1WqTUDaqXbTdY2LRysTv/Bm82MaIQrV5ICN2F6PfbYa/azG3a6ZVNgvcJCKSSOEY40
gW1LZ6iWuV8HaAqu96CQXNgFBu7E0R1PYv8wgijU15F6mesvz4foXJcJs/l6GKidZAy/j6NpoPfS
Yvy26cpi2iunGh6ibMb0noP4NIagZ3j+sYCNbJRIEnmy36Dt/otD6caVNj1htWFJC4zQItRt0lFW
k195KbBUtUgKslxcn9dZE9DhgvCA93NsBAZ3NeMXWdpIoB/zMiMbs6fFstDmZxJ5wssrefrPbqmy
Lip8SsSNWH6PPMy0aPRHV2vGKLD169G9P1iTw7OpznHaXAI6S5G434NwwxBl5BxsssfYlK5T4N7R
7OOrYL43ICDNCuynH8GMbM6favIafxR7URC7rQq4NJI1aFlJ7V2QA7eajOJFRqdl3Gr6BROShAcC
O/+5X7fBF2QpdtZ441q0+o5Q419cWbqb5fpyNl+H4I209s0ZDMenfg1wbYmhFpF9XUES7G0w7FGa
vTW/tU03GJezWXuPj3aA404hJIwHa6oSEKr5TSPjWlTEZL38W2pazSTjm/PZnKJ8rmWF1UsCj/tP
HvQGadWAaqDcvxTqbziTjUDp++Il2kcnszYLZ/BVgrJWLbc2Qc7KcTHoYtkAE3oLn18Roam1XcpW
XDOXOLpCjDFdmV6HpznlSlVbKPXDgbqpbz1mSaV4dJz/KEKEG7rqgzcYFrI5YmaoNUiwT/VMmsxd
JLSShSjpLFtBgQtL9iPQ9727L9+43jn9UDCPxEtN7U+kJNtJmNimhGk5ceqDwvxFf667MuuspOju
gwwbOWZHksD0L8rqW6eCd5fCOGGA3Vhzcfwbl5RmxeIg1NFMePbl8ATZNCdIJZFgexsvK9B2qtlj
tT8dJI/OYwGWuQdJ8tkJ+uJ/yHuXVKgnGg8N+eLW7v9W81hYyZYjC+cGo0ljnd/SmoBF29V4gKl/
gHHNY58eBZvjcjujeBunmVdfWezih24J6kUA6eUeVKIrZRrijA1Mx8Id0oq/sin8vYVyHYJo/Ihz
2bSr3tw6Yh9nlrZ0qMkD17CXtcG0Nwne9Gna87d3yO3vIqxgBtudoCJ6rApO1q7JGdfdYwT/L+OK
/U/Yxuf9IrIZtgU5HvDoZV2RUYZDc4nAeI+iV2Kfzpg6k1M+D7pF8hDeMuhtqltjbMOwWJXdaZXy
Lx6O9cSysF7Hfz8SlBYfZWd6ZAcyp7tT8sQBsCRWya6d2RIkcwrhyDEfn43xngF9+lJge4kuNMG5
KVx/or7VyBmHXZsPYjy+mZGfs2K9gGbummkCEB4rBUMNyQXGjFXpGJw1N1g3vJeJjbVCWITRMmui
6ir1EYva7NnHHV0xYcBabJtX1SciIwOJqffHLUi92G268K3UbyiL0mzrG9c1isAN2RGo6KMGTrjo
wRR4cE+wIckp4mrGcbCUUSNj8dYmOTgL5nAh1AWtfm95Zi87rqLhp3Xqs19RtYjTsTifJDZWMJ4u
kp76to9jCKMhA+dKlQIVrStr6dK7PbOUIiXoaQLH6ssvBgoCRubCW2bbU8L9Saz2OfNBcwCyInlo
/X53+oA3Yfcs7HkKVEZjbwohbCLRmn67gUyqpQj4ay9J2Z67zQQBtH7U8d3/px9T5+T+otsZkFTM
OqnRgF988qyrqLoe0hDU7BZBv0qyV8WTmFPwS8yC6I60kvy8ukVasRZpvMCLBslJIvLh5o4PRiV8
3YbeygVdnGCa0h0ormPRz/ah+ALYhkPn6Me19tmMirzGfNadk4LHgZPUDHN+tAPIAwBuIh43yLzz
+tCTeI/L74FgUZa7yiAiuqSOY63NcwtAdefVwx+EGYG159u5XZzlRpoDF+CjkiKxeX1KrMvD+wlT
mrWD6dzWi+hrkQ4zgSA8i7muHcdFkjh6UaYfMEuJm+Ndn0Jma/MbNcTMwF2dQ8U5QnLT19SUvsbb
KagrsPaLOOjmCUDQerq1G8FidffiM9EajacBHKvPZF6A4lYe6omIl6EYW/v9D4+V66MXaHkvN/7F
0dTQcEXSURDOhrQ+kZpDJhmhSkcNG66N1L3EYmU63KgkMc/tKh2LSoriqhk1yM1tawaIrcsVcfE8
d1vwU+DhUVcgo2gDLV741ecFo/8IWa85kOFKPIEJmIXGxUsvVtdMfYJsnwoVQ60Vwc4wxrrdzU4Y
y/ZtzKlW1Z5iuY+UPMTrQDVGc0xXgazIE4xo3fl2NNESye+NsgXdm+k9HN3ducUxxR6BBsdE0cUC
vh9QU0VDuYlO4isYvlu1B/5mMOSQdL0OMHH6Pattgu3/e6zs5/Ol7jCwxYgvp+1QFLk9QVC1bspj
57BlfER1ioMPzJ0UOCMakb3xW7lHNuk4L18KOfB9SAa02UaeBWdRZIoyFTTAJ2hqyZrUjZr5VbQx
UORbGvHLjJr0ew7TWFYUuAioqsFgRkpbVlcG3j36u+ChViikut6lsxbXHjnn+6ZZix2Ta3Jqr6Vk
36q8JwehVd2kzetaK6dBRDCxJS4Vok0MYQx/M88RNIcZg3O0mLThh6bEueF+AWm0UuH3M0Y1f9xs
8eaBBKZ5S2NkP77ztozexSdNrVtIeA+pnrQDaDdEixX6Cp43RhtBjclPvz2ddYJrTR3Q70REv9fW
Prli7jbuyqe40Bls0GJsJ4PHCMV0GyqSaf3DEpIc7JiM7//4HecgWgcArGcNRAzfj+9GWXFDVb6K
XnR2fSTxpz83JWgJUyc+bfmYkMLKIt1c3bRIpwDJFBLAR8RWiJ7sbJDm75UonZAxXh0GkQINj+Es
RkEwc4FJ3dq6HT0F+JsoRLBEKtJjLPTmHXsHV00mtZGIGSlDIrxeJutWdJuzC4h55Td6+Br/WWr7
dXyqNkNCbKYo8w/FnA3sjDL44dkW+b09hXj1bDlyWEtX6/rvyCnJjPsNRS0W2BNeW9NMfJZOsEN/
4H0SlXjxkoUJzUQ+z5fBIsvPLH0qsmJSOoBkOmDVDUrqApVy0amv8JE1rMZ2Yw10K9c6kZpmMfWT
gUZs/x2ooZIJ/Fr5w9dPk5Oz1GqVwQf1mMnZX+UNukz8M3nSO8VHDT9pf+eiQwvEGfl3H360F5sH
7qoYtXwMUSSHoskjKb1+XlKwK2qHjjctCc7w0GiVW6Cx43WWvQ48FrJAQxre6RYTPPF88mSyf9gj
+KCQjjRS3vVgTEIzF+ehiymeKAmhZyl52YV3zhOnNyDfVlobQYn06qelXg8a4yRmyqQfBVyrQ3yI
6jJBKCixSMA4+Ut+TIDN2kGGgW3swoGi/B7u0UVHyjdS4LD9rbpMqW/MU4TjqN2452F282gJvmet
KKoDdJpLgD6MwiPbOA4YHZhqx8OV5vJrSsv5YLr3OwV8XSfCRWtF1d9ya666BtXgxo6vnjOZ3HOP
wM+FfxOfgO4o5L3nZWRsAl3/owsBsu/BvqHWjNjQvzIbOP0hp9ASNknYQBxNL1tACk2QVqzTxFY4
nZA6rtEcYSocub/6i1SalvmEQYOoZT6SftPG8NnX7R9AQjem9lpYdBvl0PcnRmqkAOB/ryoWYL8t
6tPby0eke4k9M26yezybDtDGJbsKvnGpiGpU3wms2xGTOrtR2u4Ynr7UaqhMMdHhjswQubOh33wZ
U7N3iWW07Z+f/7lih1nJcPgr4V7CRTYovxORzU0Uk4IlDiEyOdAFwd2H/UgCtyHTNF5dyOUddffg
wxG7LQXlZ0mcoSpJ6GWb+qaBLtlKAYiJPghSkwgxX8ThhWu7vl+26YrNcxwHpkBeXjS8RqaUL63X
oS76vlFj8N0PBBic07vSST8OIp4PfPv6tOM3AKaW30muiQtv79QC8Lu00FT+T2w2tzsQOvHLD3Mc
GGNPxhbpbhNbLhv2BXspB56gWADQMIH1oTgn7pOxdOt7Duamm8XUUDQy5T/KCSpm3q/KXTK1aXl1
D1EH+xC3CX6SyH0DURc8sbRe6JjYmk30BpoH1oQpEOWR2jl6gUHJqKnRoHJQLG4w0Hf6XckRxNzB
i8rQtBPyjtG9oyiHZofX1MW2yiT8cX4G+GahIak+SI6c679C4dewg2O5OC7LoD45mu4BUABvJofv
GVp3CGxYAAaIAZuAXHVnQFt7Ox7ixRA8Kf7LL8FSX42XsTDrA6lIT6qYuTiyjFG88D1Z3WLF1FRM
PEvTIDhefrQ8Hzn7xnoC3DxCfjuM5woAquY56zZO6/Tc96f8TrZ/gt425PA3ky47EVpxMki/42C+
MiTmt5FNJZwqccsh+ziY9UJ2lNUNehIhDQxJzZ+IMTm+vLvph3sdsi6SZrtq0rY8LqMvPTy5zBdK
aO4+Czz7iNaMd9j6nlSNSwGoMRW7arQsztlMg29ShJdUpV20Xo6YjMBIY/Xu+DTYGRuyzqy79TLC
L85TcDvEQeV6VqWKTfyGxlUZIsxbSI6jpWoA8HIpxmWQxjJR/fnAKYIF9AIg4USwHpmCYSdqTcoo
ysDwH4K3vhhj3nw3RXIKMcu/KBOtLyCcpfhCOLIfgCTiIETlcxjqqWY6gnSPtsU7KWhjG7GbwqhR
grBUaxYmu+Oyw5+cSfqWuObJZTfHvg5zUucoPESB7CgKv+8su0wfGKTx1Q2UXSlVovdZadNs7hby
MAKV4mmpo0lfpVRS58kSdeWQErAyXvnXvXNucoKOKMwlejRSdyEY4cFw3R+QfPPdG7JVUjo82F7z
3igZUG2FA9WLp+oDc2BHvYwu0s6TIvyoWJp7R5aTLC+AI1TwbuFXO1b6QSIAFPbg8vl9JJJnQPVt
DfRbxRk7Oy5TYnYjjESrgt6M68WBukzRaiDRiyqkJrWoLTTsdKEUvo8JLLtw+uAUCiOcHOFbDBXp
Uo3qkGVyGGtgCH2n++NZZWiufG6W07Tcybofu/ULscBxw58+z4Fb3ZidkOTQK3nqKIDF7AfP7jl5
RDi3QFlIw2GQ0zLaBDdKMvL8eCUwWJVvj0PsE9haDkuadlbRhobWaM2b6tfEWde2Oy4nM/LL2EP8
c/xQ5pk7t4nJ62x3lPkQx02RfDdC6DhSRokE9mdmiyAgk/fz4SxtGf4LNZy/RCh/yjhPbIZxgjiy
DdhSqwgKU9BtRgLGu2fHo0BSvyqyjJ7Qa60k2nfYTgp/wGLBjbxASmNhprHRIwOrOTu1aQ1wTnCo
W2zKSBfzEa4zJINwkHTuUAmUuT57kalWMVZHG5P6eHpB0o81vrAtqnr1ILrS/D0IJDbqZR2hXOPh
yUJsPJiy/LlzxgNAlvSapaqpLsm3szLDkLT6ummVJBtAetdoJ0UBatdcD5QKttYnyS3wRimr/vb/
XCUHT6gOq9PPTPHWAXdmGJs0DrDF2lcLY5okiAX2FdFdVTA4eIrks1Ue6HO2oPkSrd5H1Rih/G7g
BqrOYodRl5fExqcQqfeDyWYrCXMlSQVW1cDBT2Pnx0t6lTk9iLX/GHUnOE15m1PiGb1Oc3COw7Bd
o7t2+kswtBr/fxpLePnhtHGERHXCw8+zPMfqC+ydZsvxVfNFW8Y3bL+dTO/dkMc+9kIlLB88KMY7
BoJvrmNUe/EBDGDot3Q4Zn1nxwaJHaJBSRiC3YHIWF6ip7cQpNnVPmqsFx9WHvi7S7NeoiVSy6fc
3og+gxdhYcAP6rkdWFerdwm/iRwhnNcSe2hQwgDQIJTxqyUM16jdAqikVsehVPiEr1KAg3Dm9gLN
p3yAlmkXj15QRPjibqsWI6vAFrFoz7E0OUh97T00lr0GN53zZLTswNb7Ae7B5H5NgRaaNF8SBiK7
aEVvNyyzRHTK1qzffEiIRCamAl13g2r2G24BqQYZz78D40SjijofQ0QRYAwV6KpgA+4MZWSjKUH2
meWct2/1aNMewrgYkE9T2/sz0mM4U3Fl7eWSflyH87vvw08eSn0SBAFetZWbccnNEzZK8+BKBF5u
LstYRBiAbMTxSkviwryJBfVPDBAMFglj/KB/WwVAlSzK6CRMlIVH8n4cRtkeIIcOE3KdLI0A69Rg
DILtf6AUpdbFNiN7MunIJ04pLNGsAjn9401knyXUAGE9L7cLh5tTQACHPQTglNeUG2gHsWjbVfVv
EW/+QZ0wV24mEZfAF1eIRbOE2CU772BVgs2MAetkI44DQP4aRMjuz7vgPgewcNpwkErF4QxFtqRu
e0r2EKisyjThMDnTepHfYG2AOB1ceI2h5E7cpp1Jt1W+Woe5QwfSCBpzgPsNmlDJVFuGTPa2Ur18
5Vp6daGwwW11iAGk4X2c2zUeNp8xv4Eb9wNU3JoGSrAJbSkMznXftt6busPFh2KVJhPVYMwZDs2Y
MFnUOIpmqstTjUeeGpQ5x4nguURicLf95ZBXIyPy8aHz/eDndppjGmRWd+m3IpRjbaGfSSXpOr8l
JEYDMSXT6cZL4WDsPFAKgdgBkR5+UhJXpgY6QiwMr3At/TjWO5+tdj4BkTK22SAZWFYkLDQ89K6x
prgruDR85j7/tDUDStm2Vluoc3Ouvo/hK7x7vcLu/+UN0tQwBk8TQ4tZ+pghWybSlzZuVlwynCLv
A4/chc8hzi77VNLqJpNAFvMFVVhh/2JuqfgL7gF/ZToQ9bLonnYo1dD6EAV52fse81O1aJkjHDe9
mebKArR9yvE/ntv1CJm8m7xaeKBcM1S4b/P89uqO9cfMHLE1haI1kUpPxcEvWQudM8iFyRWxV+YC
6Wh9wVHV/f3JB9PuvW0msg61QCQHPBsf8HBYhdTSrfbgqfVeLqo5MXTPUI9DHDgmpqmpWBUAnHUw
jfIzt+sbwtzh5bhI+yQaeyiM+prqibcWV9KlTUebGTZVvOnDnnZhcmCW/Kvk2dw4S7sWrEm1epQw
gTxzDopGy5xWDxC6kXLg8z1yQUgKylBpRLq15IymD5OpX6BYFdXZm95JlYK/KGfjDiSmJh7j7j1G
/39L+ohFiyBIVGZ8lz0SNGUF2eoHsINp2tJhdXuwfnE1ZZVxqyN1Lye9jaFLEGCy3qsRc8jeDMDx
RfWM1zspxAi4zEKMpMJtNSSWw3BwwaahY79M3kn8QDHZ+wlIvmG0tJ7z+o95RmU1EmGwMIrK3sse
vux4+dyDrsWsNRMMzJIfucbyA9VjE6BFTQHc3tGyRvA0QO7/JaEn/+PVYUITIAUetpD/tIjHhv2n
QFF1LRlxXX4yFtTh0puo3rs3kJN5qNEYbbw8K0Vdq0mp6mCnpr1v2fHGvHqyRytVUpP3UFvOxZqo
1qtjPcBDd36YoDfgSjFI5DZkqGKOMQzxeFCpKYvNcDYM0iVsnpkHk5TBRRJBIfn5pDJnYCXFSJ7N
z0v7+ZCLTS5+HC6POs4HD1toRyzXuIInqmU9JASMnqU627Y7Owl3sv0YQd+BADGtU2TDCqx3Y1+T
DoESu1eDyTripjT4isULFSgD0/D0Pc4qMooZBrHM2UWCddKG77X2jc0gB0GLSIgrdDbdZa/4P1NQ
KZveh8p7DB/vfAvVNUtMunhYtK6+LCUvt1UoGfJKy+Q4ias4GlFyvWhRu9VI9wtWj+YXP9BkAcnk
0eh5cw2ksI4aZzaYHlmNJYbgsaubJNZ7POwloK9QLim5EjlRUPvo4jj9dAApMbhwJjHH3WqeVqdn
aJ4NRMe9eHhR23scN3wTu+UVLux6/BuCdRC4hBGOhUSMNLySv8dEEvqzjoaQkPBaEZr9IyphsWqd
Jyw0Y/eAQvN7AtDqge3gqxCBvbdlKVvnGqLmBMKwmmvCwfzkhZqEFKoxUOKuJcox8WjUxBiuibbx
UV4buMHDhnD34pbG6uzt/7VQUo8mDp1mDnG6mfyXfzGN5u2TRRTHvDXtSD3h3FXqrLj08mTJ98Ek
4rosGIodmZpYRhJpD/DQS/g328ixhmzkEr1H65SiIjIbFTsG75Ca1VOZQuyVSqdFi3v+/RtbEZF0
+F80oYUYOLymdBY1qbLiW2mR27PdapVC/Xsm3Clhd63FqMKry+w0fheHXplvNJHKtZ80H1u6IDCQ
tXGDKgl29RwFKzqGDPO3CGJDf8xGSsxVTz3cniv5y1VETQIFFt3HUuZOB6azHYTXG0BiVdYMalnH
Ix78+ehVi9HjMG8ifsWSHEC2K8Sdp4OOPWfkQq/Ea0R8UUEm0RQ5Gw0r6KERk7fWmIF2pY1xJb7Q
T/EOxEDMJrBkh7H3WOPCv6/whjCmoMH0TLXdIV5b35fG3PlFWhtb05nh+3TmfNFx9MNV1zxbojY4
5yqQ3pXiP7ZxAUUUfXq3Ygt771XPh69VHSUnOMJOVagIF8+FpWL90SJ8b4iCiURjbk5L8dRCs61U
t/0fiKsNDhczCyRDHMirzF5CPTut+3bAk6Ixds5WrLc+Y6J2SnIcgLl2Ij+x+a8aiOQWTRWdv4PC
mXPCp9VRmxbcrkkfPvlf3mAOy/b15j8Zd8yWZLEQMBjULCwwAs+D65rmlsw7n7oYZtD05Q4WryOV
uALg5OGfar+06LqP8sM2H2g+ZIeSUDtOg3ql4PbBmNm8nHpJBaVYKwS1t4vtPSfYyOYVCeipb81I
XYhDPD6NvWpGYOSsDFeFQ0VF9fejWmXE9K9AJ4D+NPvTOGCWK1poGTheKLPTOwwK8+JbxCAyyjud
iC6kCOvAQ2vYtcZ2Tw67HUjVkTUWwUEpMSPl0tI+o5O1ZESY5cSR9mWj2wcb7Hg4eIiEZ5ssWkJa
UzWybLZd760ymNs31pmfY85Q++A3bOyVXnNaBnzApyHFLkCkfIfonuZlKQznjp9kKuT+17UAoJaF
2v1vjG3X3Z7/ZA/QQTIwwnORW3K0LqOaZNCla+aIncmr0WqxQs15FhQnTAmw/3dAOwl0QNJHC5Ud
e1eKou0ZR2PKhcznzTD2N1dU5cSIXmwrfW+zI65CwGVXM7tsdQxiuWPezd1oWRr1+H5TCI8gVQjq
xC9akeJLACJoh98t63GkvKtvJ8sVCbY6snli3FJMFmVgNqNpAoMPW/xMtnsy9LoJIS3IkECobfIA
u64Q8A2wR3tN8DDq1IvL/j2jb5rdwNlGqldHGaN5VkhyOLvdVu4FwTerkmXwqtbI58/Xvgnqe9Av
2Da2zY0uzid+HEcL/t5p7QNvPKXHgIeDAGb4LpgUTU8G3Cu3kYiIxoYu6GqmuadsYjP5qkf9Dnrd
P0aMSlyDttR4husYw+pO6Q3iMYbhQlcMHGm7M7QdzM8JcIQJ4MZ5bE97jhFSI1naIZb+2xGhtpsr
ZHOM9Wj0gI/itiCocICN/BUQWTgYpwsPaFcDBzkxlAKVoepAktrYm7tS1JDHy8Hx6sPQyQsYIeZ5
/6KFacMhhuemFe9Ku9MQsBmCSP49lQvfnzMfUHwucFvLLWK75tGrFXIB2FzmWDF+A8eFa0eygdaO
dSz7mb4XfCng8LR6CdJ8qm5qVho3Sz2PnYo6yNNenrqTDDJh13EUN3DFBBEkTSED9MS1jLV1QcsL
NlwSyW9Ie6eDiNJUHv+VzMJ9xrt74WWx1akDoJsCcUTLdWqQ764lw5malF3N23k5HO8q7KCuf7vt
MdvhfaUnJ3PhudmgZrnRG77pNO4nPkbWIekq4+XJ+vd9szYEC7p/A+wjDTvBt44JIG2I5+X8RFlB
pk7DJARfPRitcVGRNyD/71t6zEcbtF9m9WKraChFvTPVTrzGHPTnaIOXZRtWMXfPgcCXaWUld+60
I1+/5ku/Ap6tjI/MBM1WZX/no3bR2tjRRT2gcaMLndH3L+BBmQ4cx09ezBe3gSKBlEen0acoXdMB
h2KBNITAqhYtjZST/Qdn3lIOVjHLXysxmf+J41h8soCj5TqjpTxK9eQ1ViniQGJPPpc35gh5bYZl
511S50ZgFIyts2u5iT0QXyWfFkB9LZITufSZtjvDwYt8w6x+geRQieIFg0gDceXv1x5MmXmhnrDQ
vWDDYYaTfJp7VmAR7lUG9Nw+vCQMxuKIHdmTq3/N7yhAYPThe4pqXzuhRmNKk/NEK2RyPbs6YMff
5D9GJH+qao1z3uzPKFkGLh8eKEuiit5bLdGrCUiGVqA5tfCRQPb6VdnRkS7a66vA+uA+T/sdVE+c
fz0GyuR5UhkHLGEFpJsIfqSGauBZDJnppLTeo/KvleZr0wYB54HJGfjXSR2b8wILKC5CJ9IgTBlX
6ewVkuEsLdzgyN93Lx2M3kzfM7NcHcwoAdAYQrHyRIvoZ0YWNX4EiZy8wh5rR2yd5C2EfpLg+NaB
LrpV0daDtthpdkwfSSwLi67ZiSQDH5xhnR5zE1PLCvSiCKgG/OyU9Bvhv8AUp/fJcvId0PrijEyi
n/F6FPyIElYbKwEY/3LIuzlBuTIkbyjvME9qjQRB6DeUq1rVjNrFTSjbGTh5956AxjZp6bS3A3Tq
/AmVzKCa8cbEwK5Jbvk5DfQEBcLk7LrnNzp2NbvZHCOnvH1por4Hi0V6F3cadNF9mitwlvH3nJw9
L2887fxUUkz4INYaEUJMaESsSAJrGO6nDZMVPIVuGWD1TR6X2EXkANRc9+NiUErb/wHpDfHu8oe8
H7drihmVzRWBgGiUJAbjZxtF4LY6svCwviWt78pSBoNlzLo4sPRxeYTe+uXmfYj/LbfyeRCc/eKl
9gwf4k9kmSXQbCnomJ5bvFf3uIKUJsAAIwsIbPDs5tS5KiLWejtAGCyE+lgJC7Q11rU+kthfUrKc
BC1b7yt3PpcpDMUOfiL10km83GbBz4VKC7qFHQwQzVrlRmyPWJV1dCDHQCeMc2+etVtAwNtM0CJm
itgMhOQTfT8j3irSQ1IM47SK1HmCcrUvWcoAd4S2i5x4hFf5za68ehzhT25ZC96Xi2V4BnZYV8jV
8YucF1UlX0H+lM+ciruStfteS99HoZIzUllX44Njh5APOj1cmSwtx9XfdEF59ImJ9CefCc4A7mjD
E7XvBZoo9JB8KF+plAKLZshV5axbXbH6Cl1B/FrUlpuWp1dzHz/A0tVOYXjmujJQR8ATpZ5cMjRh
7A8Vz6Kowy7SsGSRsYOro1pzIQMe1qLkmaPRHAyDhMZC01IpnKa0YJozkmmJSeGd4yaH0pk/7YpF
D+KtIxAA/m3ARi71N/7LrZIFy1HplTO0KECFvbZJGniU/ktNT2XS+iNqsxefjSLIQcn6Vz7gUWC8
jaBcXo3zYOo0pXsoceeZ6hDXpE6WudF0WoZ4Qmp0DKfsQT9ggFgloNTtWpb7WwSmp7iUfHS1N425
+02uTJGS1OMayMJz9GtH7Z9hTZ+CaNGdSOU1A4AAL19VW3Lvbgy3cWxebVy3BpBsKeK1gvqg6tht
4PMkITDp9xHV3YFCFOvskY/6iwuBtvyUxdBR+X/lfn9rYlYtRh/W4UhBcrycfDZA7gnd+vyR7LSn
RULD5FfzfhJRpVZSwmVvBrYrqVaibqkW/WjlH8aWGTjdscJ4b1sB/8fjJEpYPHoqHzWzIUElZ3e0
ShSQrRkm9L2qXJwAfVFOCkvE2DOMf9j0uF5TYRuLxyasuTndn9jhZHiYrVvi8YFRUPNxVD/8FO/i
8GhT1nqiNNbD5K0UClEt+H89lBAPVF5Rk3nfIbWeVbzAmVcjp+WhXNtiwtthc9gDosgF1myAaHHY
hkEWtodE3ZO1cHuWLptnYRUGYDcMP5wcyDDNplJTqZZ7LIxIXU9liOsKscyzc9rsX/jfgfLBckpA
rTyyMKpYJjy9KvAQoeHtLzN+K5JIWVG5tCQGhm+j9LrLnl2I58ObtGjP1zsynfaFHVX7ugE8/BGc
zmJi7q7zzHngXwN6E7XIJGqGff/eGUx7wQ/W+vzsA0NmQ/6WHNYMWzUPeQhdwc0JNP2xmuxVWuYL
7oknKWHWYXobPuFuAT82ySNSxnrM2SpBOBFKYRhVP+j3UdzdVf129iOzVo1jLvv7ANAWN4X4WsXA
mugn/8+AtjnGMgydHL/oKlrm0bSMMgNapOLPXYrnKr9QxDPaqEO1FFVb1ea653rIMe5zPwt4zR3r
oDYsVFD/muLDMGYbWreWm4aXPg7wAJtMkAQc2z/Nk5RJnwxfZJpkEDlGFI9QYpC9263oDY4y5u0N
oo2WeTOEAW6m7ko9B+M77ifg8tbsSd6/kD69hGZyBveGuEy/9WFYEil6l06j6IdyDtDqy7eSh4GB
sqGJNIN1xcPbufTdf4GhCEctYQ4ti56wAgrJ6DaqePIqDovj1VRr+zVd9gAfs54hLw7p49tbHOAl
MAEcYwaB5phmCH38CTtjXsJrRmE8jkI+pTBhIU8D3GOSU5wqKgf0q7jfl6qF60OKKSYVsOSQ2kvb
mb0VD0CV2aEYXFdH5glUfKwhHBQJgOa/pjS+Fq1lyxqbLBoTZyn3XCs5Q0QMB1RUgEkSTcS5d6Bg
UCgpqKbe8w7PBgrAuJ5mAIS6VCuri3VWrrzy+g4+0tTQUh9RGykcPytctAcrrtl4AWx0q7c+lXvR
yI4bt/9aGsnsaZaAQdAHP6uZkDP1tSoea+zcdV0wMyf/u/Na43Fjw42u/uBQ7dASGMNIosL9TILq
340luc1hpBd+uNLwRbdYfaVieedbReqpoIbSnol/dcZNcr7YIzdbQzOqXH4tDGx9i4JVxnMk37E/
0HSMwc0tkRT6IhL+qvcpgYqa43DczjbEqhMr0BMzNNe5G/WI5vYa9T/jzU9RSkj+afSf7E0OB2wT
+sJyxzHrkkGlUaP35xIAyRsq2v1D+7GgpGurI1B3bzygINXYgAvnuEUCJ0dzH62p9adoqiVk3ff7
toyw5fdJP+UPlLdBllDkUzxsNyfiAfkAGiPdtjEL2Lz/djD1xl0NHojLnRj0BzGhfgL0KTP72/Td
VNxgWc0HwM9RogzQ63gZSEdtwqm5fRbZUEWvHY6uoGv1tAt4z/mj2BnwrsjJwXRJfM/45M2aF5sb
2e/ez2T8mcex6VcyOY3IF0Fd+ROZ5KoasEU+5sdhYCmPWMHZK5poOG1xms/R4dPdnVKJBnGEieJF
EpJcK9XXWoQVAUqcxGJGEVDOlNLb5NhSp3/Br/1A57FGKU9VfGz2zmwxFJyuRnDYjevUcOOnlLG9
u0bYOnDhjmTFyX5NC/asmacHKVz8WJ6y49uZJ1L8j496da/m1KMOaM78i6gqbZuVKxQsGVFbZ5Y5
4GZPWo0s22+sb+nP7ERy1dithOrrfsanGYuA1EqxLpr+nsSNsIGDKnGuqI2ZVxwu9W0CbQ/zfXgf
BIQDBZ5NZrr5yeKoSpbjjV9DiwWFMT5K+dt0ovFsejA1Wy+GTELq9HxGcbBxLn1Vsb+Qhiy1n3Rb
FaH4lMdxSnaQKEEWKnOx5v2T05RTeHF4r4g663NgovvI0I9EZy830AZuVa8Lwx1l3phswDZUox/8
fuG46k7lvo+I4JOVusD/nJQOWmkWaCkHI1oUoUgGOk8PcInHlrcjtu+glZTHmVne3+KPeIuGZIP6
JsqFdyxk/2Dq4fP3N7/q7BHMj2YbhKAn4L6ZqWyiPnIlCTrq7Swrzli/PtiYXvc8ZVNp6+Lli916
h08v6hdOZYMf47j6UBa7uRHgWKvl2j+kuhAKRqFcyWjTptE/9bSYlw1fjQgUSPWSt1nmL5TqEfVp
H52J6mMsgwpbsThCol+TczlHVB67QX+L6y2wUd0IUJ+9IEqfgR8lZbS28wwXViSZQGON2HGqeNBx
83eIr0wHt9J838sC12yhwpSNpXOg+6y1v8cj6mt2vV1AfLteF3JDrOUVjsCuEzVVj83MpHV6mvJv
ilfSkkptd+3MuBfvRlDF/ZTlz2tu8M40oY4wzJ1QuwZA2qwm2G32dJR6nyKUiGr+aFLtguyMKAuy
pYqFoX/RAAwZ15pE3Eflcmn4aDRs/P3Wa4BZSwIA0ggParseiuPzHrixzTquPC5x9MPzyjPfp8pI
waVob7BFvHkNTTSxqlQ1FM1VI7jaAAwV4L60H6lRZ5dxrNkB4h68AIZ7bB5/EcVfbdkF+zLuKxEt
w1CjEM1/qsdZy4GdTLPiWIwZzSRsCj2aZIQ2uuwR0oa4cNMi9mbc0ERZw7+xz2MsIveuXErmFg+/
nrInAPvGdzaGnSPsdcbFyWG9iIisMvM/9m1a9zqaaW4R6rZGzc9MniZDdHdypLj+/EEvqx+GLX8t
SSIExmAMnw0HbgDEH+3OPJwMuVXdZWiB7MUYXesn20c67r84MfGy0zZu+rdj30sh8YeBt5JuN7bY
9+Cv3Gjvh1elZIqHKijCLpouDpR3m3wsVv6GkHHTclaODNPlrTkHjmIyJ0uMkPFGiDSkRk+fyeCb
rUFTm0JStP9KCNbY44ZcAgbRJb5PHqWHAuawa53RCck6sv/T5/MFFbPgDmfS60Bz8xHjrhmTL8Tu
ApbYI3J5RdCGeoqlTm5PJ6BHtrfWQXFJFmfjI0RyVIiMDGpZPzJI4GW7/D4OLwDZDt287T/XAcGQ
uxnjPyxvPjn+mwCxaYNnU2eDyTOyLR9B4uCAVV7jM5N7WCG9ZOeOL07IhpcZiUNo1pc/6Z0gvLWa
SMZqBjofQm+pqDIFRYOsAxDQCtRYI3A4+UFQqWg2/xDwlGbt0RqiQlj4hUyEcTofuiMzULv+emwH
bLME6w3zJ3iAzg7cKXWRyKDYQ0Z7MJgqA0A56l4g2ne9HYFBCcZTmH+UT33MwEGxnMX8d6+C4eyi
QY1v4oDamoPh8Pxyc/OvLW3brYGmtF1pBkXknYOqVxVzZMM3lzSWBAHzCThsTI67+rBxCABsmf/P
tsVb162s1dfT0iQRuy1zhTfR5PEtdIDDK4eUzaGVjB9wbsBWS3ewbuFa4poPvq3GPx2ipuyS8N2j
RafCM0rDDojbwjnQ3UjYNZKbjOYuw/hAL7+p/a3x5tsCqbMYxLNt45Qo4XDQiLhW965XfskYONpc
MjEfnSRDjG3tPljpry6XN7ABY6js1WiEGZ/jgwF1OpQ7QUklxQNeFyBr7zJbLykBHk4yc1ryuC8y
AjDlmsm9N26vxQ420L1cSl+QFJJH8Nyd5czz8C6PUPHKpmo9jLNIdNJp39kNrUTLk2EtnO7fliMa
VM7NCc/oTDt83yX94bqt5Ycdr9GaAjO7Rgy5Vphj+eOH3uxFB7JMKgjrEt6MgrupsT0hVNOvH5Yk
AKYjxM5sLGC8+7yF6hEYVzEUTWbaCHto9lRwBDXV4nz4r72E0tyVeaMs0qhi44JDW4J5l8xzWtTi
VuNm19cvW1fhZzraH0LJRNXl4o7cTEDPBMQcg9BnSdW3vg3OPHHgrfrGvw4O/kTzwgtUHeWsEvL+
WKJlkUjKrZfkwPkWCrNDReNajKQCq5W4NEzSIAbbw2iP5uzEnKI6Z4DDCGqmlXymKqHOdnSf5cgw
PHIeCNvqEGXQGBGgIDnQLqzyzazJAcDctKi/4Av1mpqqakHiehP52D2t8uLZ18OVfGfbTyhoRYTb
LaZZRZhmuVJcIGlxMpTznx8ZnDJTY0S4Jkc+KWeokkkc7kuE5HNmDHTG/sCK9+9k+NF4vsj4Dqe0
5qQs6b2TDMyTTGGQUufq+SME5T9l/FIwiafKMO2lSBV/JhuMHGnIIiUWt67d3FA3RPzFV0Mm70EH
03M7dOGxRW7iHxscsePBPuGEQWw7AQQcaa5TVTmDuDD6NmAXDddY6IBrOm+J7F0ii4mbqP3inn4m
Yt2TQ3OAw5JFlgODlIZobJQqDYqTEZRmeXwYPIul24awtlo04pkolj6G0ugUEzI6LZko1SXUXZ5R
8nA2EsQqSP3mOU1hw8F8h7JDqoVXaLbwqLCJ2b8a8ho9AHhljfxoU7jW0GlA+InExFJG1cphAmD7
FMKCHkcGxpBXXJu11FbY6hzLXDvADGYXvb5nN2GGNj3xzr41BWA4WUVjICS7Wt7RLF09EyJvepdm
rfFp2GebQhbWOXBAzf7Rpk4CQPVTtz51Qpat4DN+TFOI8xkbAxrhVcWfP/lJWzVmo7kUEH/x+Q1g
K3YOJ1OT74/Fu4lR0JjPJwU6kbvUsv6vhUR2NqvAUgPAld9tXLRYohyfry+PthZKWLLGVexNQw+L
cbiHvuRzWYtWblFj0hFdHG2TmiipOb51YRy8WQiujJGNDGQSw/iWjHo6nU3iHUR1rHo59L+zCYnF
If8vLUzr57su846KOWO/czx2I4tHIRCgkuAKvsPiD8B5HTVZwkcUpiPM4btlVU8lJblKSkyJrVpt
azdfr7XR0k3bm6BdsnUWxyOAgh2MlEyzMP3RQc6mdeN7YZ45y02Js+Q6Au4irV6IEr+T2FTTdaMo
BX1rMS/P/vj0Jx8B6hgohDR8dGosMNhhb111KzKqvgNh5hDbZ9/9yoMhTXW8Zi9CENcpUrpsYzsu
Amyqka/jf4N/eHKplIWsQaPhp3U7DNTZaaY61gkZGKFEfhmHWoDZs7Y8hKMU+I8+W0wDS9AtcfX4
bOLna7Q1EqG806VZ3UTFa/gUU9LPl6zoknnwnMc1f2sg7o/uRfs1xqP/kHCyRQxIrvP+2GDjvhRu
a144gd7PVbTtP3Bex05UtOhSfKPthbJxMVsiWYmv7acIAVqxG3akJvn4yRcy3p7ps6cQRE/g3wJq
9LKjjqPRLQvwGWDLlwalbhA2puEA7JIjgj7r18krB6IeNhv2lQEM5jQmHfq8u2LvVh9xgoPsiAnM
VKFsGqYavcWQ3Q5q9G232XRQMEnuknQ1G2NVjoJlK2pU4deGxkzX+RPmdMfR0ulB2/jZrHAmRVBq
cx9Fuw921xTmpCms4VNsDMSe1i9cZ5fXZzmsT+zBX8E4sInJgAQcyEq8sjuJaWSwZb3kBaCo6NQ+
zTmR3BnxUwNWpxMI+IRA1phlN7gHQzym+bs6ipnwqszShtjAAFbq6Npxnj8kj8bcbFO+SaXVYrMi
uasekAnJsAISANjHk422uiOWcEoAIcCivkm1RmanPZLt9k2YaIc14AJIogTmFZgXIN8aSGc+JviN
vri96n+533IBivfw2lie3/YN8EQoXbhd55i5JMz49zbwNoRKDY36ReQY1MZyaPdOxrU0h9g7JhsQ
sXapFQ8xnLsCjRaqEw3nD5insGFET7Lv0xWsrUNVkeO5cy4HVpX+7s8uWwL6UZ6d47tAWGVOtfNy
r9W/sUo43pohrVsI3/apS3bDmUMxqrk6za/i+1o9ayYwSI/tTQh825H3D777Es85kfq4invo2PIX
ZmScTbNbMl3/TiAstDYVlSpUwIvTxsBflDFraOvOunY0RLlt4DxR+CEOOIFWv+TWx54Wdf1ynywh
z6JU+2xB41arecGbMhGa9zzhtxRVbGhSvBK0luku/5LzKLlI2Gdu4YiO6BEmDJIIQTdLDzmZtvSa
wnsj7pYjMFGFqOAdOTVCHU0e5y76hEco8D1L5OeD7Dvy3CoNaXT5+Gaxf6Ah0LO7g5q+BWO/pCMR
6PizZ4KNB1/VjeCVO/B7vbepC7PEX3zVMIZarPou9Z18E2IYnaJKZ68kWeN9AdZdTiszB2FnSP1t
v0VsA2lSbhcSZPsdB+CmRWP5X1HKVeQwKogfe6MzTtHx92vTDLcgwixN1IPTKsXaWI9B08YNPnj3
2AOpCwFCULGlI69eFBxbFQUHUXJ3RMu0QDFV4h++YD7vKNXT5BgR5e4N9F+zXoPtKKyXO6s9yNtg
Hu3vkknLJGErKY8UpVGLSMPwkMKJ+iAdYovm5lHaJlyKbQdvYvt+T6beSQ7WhmCWJLsVsnskxwzA
BhlzZ0Kr+C/dptnz6u5r7MKAjfmiNmG1JukrlatGo7nLCT476bwP++GLJtT55wflUPNdm7hUjYnQ
3DPMqz43qE8GDFVoIaRs6lbUuPxclVQLo5WdMoxFwVo/IMPZd1P7UOJt2FaK4s7iK+FNsLtz1BC6
OdTRjXQDEikB7LwrFzqTedHW0HUEUHPJX5H8tGTfn1qsLk/Al6+4nKUJuJCjd4dcL+86/zGNzE2a
9Qk9GiMFbTWe9dre+iaqZX4Fq9zimXav5iNh8UvMPZPGYvQpgR85LHNs3hpHIA6TPw1AcJk0ieae
w1o4DEuWCnJha6D80Zr3Hj23s0RPeT5BNesBghiTHc60xEfszVlHYRIFJz+8dPougHYUI0MhOVZm
ruPIhZdtVZaq+E595LSxmNDgL6pJvmsUi3pYOwPRpZa1hRLYqkMkbqJvTBWLlhOrqjn4wiZM9TwA
oowDvlcwGrTr0Iuneis4Oci9RBDqcsw59WIyhx/wccmgyFwzCccoxbqEQmZgBsh1k577Y7kqniBb
aIFe15rsN1xtyShDzi+w4/J4PfDzpSc0sByAGdZRZQohjFxQzHvG3iNYzV/dM4cB88uS2mf61twb
xhUglODatu3q2lMdLufIpTqad+MGum4RCQFXE4w235MHqi5qdhV9wZY9LLgHg6hcfOiy75Gr3UwW
YId4wofZIlmK6pEPFRN+zjoCPC7kIIyW9yc+/Bs8bnpZgvlXb/s575NIiwIwAUInHvJO6kyNVBQD
e3VJ/GgyvtCJlKR0qrbZSt84uGiBOe90qGu83GBfvVs0w3hByUifKoHEkkHGW9bLCC2A37xzAVrv
Owc48r3Kg14dcLdc985wOLfOZg15VlOV/lKyuks0lEGmSvdRzLe3IUFw0VxOSglRa69qxCywC433
gb0bvv0ks01O+skREXqcfWx7I+Mn1L1K2YmLlHbmuYY4y9oEuP8Kpox7FzlI361Uq82VG/a36s5g
y8ZZ7waCBrddPuVXPT1Wy5HSeAaRdV80tvO6pMEbbF1jTFdpmR3r5szFPCpNLoScnINJrPlnqqVv
F3Tj46CUud/LO7rqYRaNxRAn+XFvezTeyK0wtqSPSSYYAnyAJHBU/U0UQi2C+8erRxtX7crLgaEh
n7YtLPkwGMsXMMumPiiJyHa8i3XiQG0szhcFRhL6TikB/LvnR7G+xjPDS/33sZjxli4J7t/6MABe
rLDQdrn3FG5BWBJS7lmMQELvDpmh0ltwkw8Gu/60k2WTk0/emP0W9Ptip6m/YIXqdo5J3aelILlb
N/NSHDkOncyblv+QUchcXGKWEln+jCZNPhBWplda6w7KyrcP7rBqFXh+Fm5kpkFMVaLz2kfwUi27
nqJCvLJkEN3fqqEn1FNywSHm1KjcU9a4xyiQRg8qB20L3Jg9JKelcWa3JWb9mgiIWB8tcTi7SCQv
cV5A/xLLSBragnmZBzrSvQqRci0n5LrXk5U8IKXhTkC+iKna6OzSoUikXdlK0LJksf+lNfzER9i+
PNYHYskkhsEs0CnrBgV4qeTvDv8X46F5/56EDJiU3Me3lSQy47ojHS6mkbf5dNMPygSMwf0lQ3HX
s4yqDZPVYTmiV9OP3yTVbEH7pFKucj81ms5O6coN3JwpRY2L2A3RsVA3TQkiyxX3YGt4+WT6v6gE
RI0KJelV/OyQ6l1JUccZdoMVpEKwOA/bMfGXPCPSJGeQukMaq48u9eATmwxfvjXqOf9kJPeayo51
ZkiazADpCqSMcGWpjcNlg+X4MEYjOiD/iZ5oE4VYhZBG+yYsvyLyJHuwg/vOyF5QVD8cP8iMsq0N
3XwvEwAQQ1hlXlThK8hsBvPBKxfOfpSS64mo5lZ1r6Jn+hc+n+wAMELKjroTFluTPAla4x43cEL/
ELyv0rzrGjiDIECu54+6S2BR/fa5oNf3BoxXJBRrn6+BcI1AAOehk/JmCc4pxsz3FEFE/LY+sX/3
a9W3HQwtfzNa7EN/wDAOtM46AVCbH/kWl1aheqAPueAvKXKyq6dwXAmk2b0AitLcImwHCIO5iPNs
7/dBdVjZUnTnjzeYIELuENKUH7m+r259WglP+PjjLa9OApPLxDymK02+vbzwDKlAzYHEcJH/TKg+
B+VspK6HK7IBfBYCyRwhlsYZBKt70AvlCzFc4XLSEZvAPlVGHfyj4y86s0PjNgin5/hBzn3Qs7Tg
CLdAAD5saJxD3EfGRJFIgtlo/O+beips1wvnDHEQK16U2mUdkj2DAPscGiU0bxgAn72iIRdeZxuv
Q4uI2fRz02KtmRxdVbg+n6ugmuzAiNe9mT4G5kNft2sg52URzGAVPe99UhuQOZYaVs6AxNnkhPtk
qhPyGvC3410qrzk6mbP1rsI/l1J4HxDZ86YyMdj2hsvDtl3psAdMgKFiPcyATXdAHNsFlseP7+0l
HQczaBME1jjs2AhO6u072s5nskC2Vqq/2/8qUCaN6gTgqLnAj/0YfALhO65OBW/q2+8TlDDIoV8B
2cge5TOwqHfJ07sPtzYXdJzIVh2szsHo7LlB36EQ985z3ktCYn17pWSc0EMnZTq3FTb8sJfw7/b0
oIfVGFljBHb0un2Fwy+ccwDZ5BsoGhGNvZKQoaTvxnyQooHqt/OsVXGaB+uoK/DauLQLdHRjXlV2
j4PgLBQff1PoqbpgXaplzDciTxe0hmClhD9SdHxnnKpDJpEPM2pBkdAaRnhTB8dFMoZe5isqD3O/
dg346nM9oQsuLVcmN2UynQZpGzgpiK4AfOEanM6V05/wFhzr9Gz7rPd8OFYDGuR+nUOEMVSwXTad
2mQmYG0+i/TPX/QRwtDjCXIHOV8tIfvuI322j8Fxu75m7FZLjglO4z+8GCtn/Z1EAOxnguLS0fmr
iDv7i94vjL7F1s6tHO0WnLKvZJK8hTek58E7yDuy80TwwebuJkk/CrZVtYie0Bosarf0SBBtr/zL
BeVyQfrV1h8y5l2kXrAi1b+SpBh3mcx72/SuOVkoeziN/xNpcTVu02k5jmWAfi6i0uTDVfkw7zuy
Ua7vuQX9OJF4ByT8qDC3DvPS5FSgUsyxd0YJhdK4q5g+Gqdf2cuWI996CXPTgt94ejarVva8eIdj
4oNzfUCzvoiXnPPL4GBtmaVZkW9iH/fTj0MGeXifPql0GKKvW/kCKm9y+gtMj7v9/rsWrqOsJcJJ
s8iTsx+E2oTZfYBf2EqMSD26Cwqb++w7oJhejIR2Pptqwrj3mUkceCK0zNQtuFJRuJAVq7BsYgDQ
ATEHmv8JccMUmzULr688yr5qEuJDjuWKl+6hH9NsG2Urh2zZP81bLhcdgR2KTItuoKzYP0LQ1jzq
pNjZjhL28fb1wWzzMZeMMa4dNwr9IeaJq1uLHvHthn1u2H5ej9K1PvfYrzzufgXMRbNTVigwmTBe
w7djAWnQgApJREL6kMlZN238meyTChz8BKFhzjbCBQwzdHfrGHeEGgBdtwdURTCpggLRWk8HpLzA
mXyMg7WNephpdH/lSevyLeIFIGlmS4Laft8ZZwW/al7bDVp3uPsRbtp22nFYjiD1l9eXytXoFNyh
QpcaD1d6453tTKddjDBqC6u4x8w8IsFFbAgsWJYXHH6IDyUIEDUg7ARdButktD42alWz+bYfWld9
U7cM+LbhiNJVchtqwT7LjZE78A/Y3+jzBHYTsKqLYpZO0QktXKsAhYOBTfbYbMMHiN9pDMHd2Y0c
LYnNHy5Sm9MUBHEUbNXr5COk2jcRqu8Xdrckum58tiRp6VaAJ+qwrF3jiy9zBC3jbCAtEc+wWM7Q
TIqxDvsSUCes+IyW4Re13PTqYkH7YH4DR7jKETrEeOoEE+rqaauyfhsLslXy7YfosqxXmlQgaNdG
NkZznyMEUshde3wxOIFq72TlhbQ4Wz82u1il0Ogtt4Ngy7L7kRrebLwn2IqFdUV23xrKSZqk8IFB
sr5K2NzrssmgYtIsNbNnpvCrhxyp7djlmltEPaXxixOx4JjELe0FZm1wV/dQZ2SqHOWQBTSl6rk/
USWqK8pEQd3AZ9boC86xI7LLxo+NNsa4rXVZsdevSIjVQqyzxhp2Y8u1EuGL4REa37b9DDvVW09a
MPa5auNZn7JiGWqDVl7/7Eh78tV45kYBuadhY9qBCku2AgnqHNfgEHka6432boUCeVfHnRTedCyx
xI2LjQIG9DLPOPXnZ7hp4NSezher+lLnN6TD7ZBTc23ejXxgXQX0MheOxQvQinkHh5zhBZ1Esf+9
NRRec6GXWYlCd3YViNzx7F+TXhb97S0uFWcYiCg/PaQ6e+JI5z9wj6YvJpp0ZR0YIgOZXDIFP8cG
SA2P1sTuLb+2VwpwaqiRx1NJhJXwmzondPoNYNbEkAg1D0oqkQo2z9gEqCt6gyKB2gys7Y8niXOx
HF6tkAMr3uYrUUJjpb3rSVbuWKuZ3tTL8dDqHq9SS+bTarxUJaRTs5J3Hu8UM0wQADa0z5XE8R+1
I+1/AMU5nb3d4gw5ookKdfPdwyt7ZqkXTFrkUCTaOOV68ZJeTEgKwOYbY+aDfv/bB3Ugw3qng5Mm
6KOV7BRosya6lbuVXlU7wNe4RDpQGSIuejKhhrlHX9rRJhR4IEhNwZLi3avU3YU8gjQK+wRRjc9I
hK6OVnfdRquLhQod8ZVN1jhpAov+qHDFTK13ebYNrEtVnuOwwpHSQbSmBza0I2pQe13rrplyQhJU
Fsb4W6Q7cFA7z5StTKWT2ccGPbEm1R5fCCwGSCmrODNjMB1PeW4lkWiXgl1hijQAQo7FnTgHZznD
x0RmSejhtWYbSJ7vOzVGbGnw40bitqmjFbtE9mScyqphmsogdzVZgDBp0VTgw6PggIn6hnBXDogI
4mJojvq97EnTh/SpKwGWpyFzEB/48K4SbdT+8ltIboN1KUGaXCy7i+ClDQnemGJCg+UxGdXGcSHk
+4a3NLJqS6jDBKXeM8NLLNXsGhIDojbfJOQxpUqxKUPP+TQBIzqr3BBawDxrdukNLgzoTLNzfZHC
uRaMvEJf9/6zSn084rKd9kTKI+6oz9CkFNaf9QKNQt0SL7g9qVNiz8sPYuIuct8YxSk8m2MDF7+t
BRtuBk/atiVUxJwf1KumUi8dXxLFHWGOo8mhZ2kmGSWZpnUJUWc9HAiQ03Ryh9wYi/yRy4sbcOFJ
xIv6EXuMLNgblvD5zEvfNcq9w3wdvQjvHK4E28ikLIAKpFsW4IKzGJiYf7PB99T6ZoMHId0OE+0n
sRejkrevAqo4uiU2w6xxLR1x+LPL/aRwhgSafs4B8XV1riy09RzRZ3HGXacWNXbfJVHnsvUjgV91
TGBP1qORQsUTfCZIxlCR89tWFElRY0Qx6ASoOUskL2zGcHbmgxytb9qTAmIKf2K66c5m71PKpfyb
f58okIrX5NfLJeqnQtyJpnYZePduQ4IphSHLiPZP3lrRJ7CMxOW5uZYfNAfRtCsfhNlpXmkfH4re
ZTTTcY9O2++0iXOI+xD/bSoly7TNkBi0cRyWM4qKqAcwbfhcFT1YoVFhdNyFWxkfFGSnwq5/TyiU
ZwtAvDLSy9fhSeUJjoS+xomHuxzyVJuwWsum8BLjuRi5a3iVAJsYvuOv0jFZn8fZbIVgzWZPXj8r
tqPyGvbKFdu5KfSpmHd/KIa6dbwBwrQAObpoHNVX69v6y168P4+eeAZtc+bkNQ6R3Rtwlq7JYyGC
jRCtFR7kxMTgQcKgh4oi88NaH5gzBwL1VSFnOCshNnwRhgmLyH7H3sBbGL8zVqsyxyuT18kk5iGT
UGHSfhBA2gE0fYdmjvbC5jUzo4zb9+9c+u2Ua3ypmVSXGpi31mnnYdRwErSF1WKWKlScO7IWuHN6
iPfeuKSgjINcQZkFm9AgPyAqps2TNVFYbZFm1pcJ1rxo6lgw25fotaOTKP4ESqLijwYIQleB9HC1
do1AVqm3s2qxG2rx2oIYU6HBNm64tAdDgf9177z3hkgyC5Ebd5AJIqUKHLItEqnCkrX1mwVHjkM0
2lwqvb7SXzOnNFZNmlRTbBluzWXmfoyAQ1lQgf8LjuBOblClqe3RMwxPQ9IMIrbg4YA+cuw7Skod
VjorLH/z6bUCWKwTnnDAsdoHvWo0oRHBDy6OVZNyL2Oe/4P1E9z6gSs9FAbNj6fY32Qoqc+Qmjmg
gPZXkzaVtuDSC+A6ngiTplx5DlQnLL+/63HFHmwiUsggmKpbFFfjDgaztrBqql2IG+IFttJ1dy6w
h42K8XXCx5WiKwPvHM9PAB3LQRVC0KhXxRvrzZojDCWg3l8PweCJ0UATad9UNRka+O/6skzO75qK
JTRGIy2lXFiXB/heWXn+8vHm6MiGEUSR+zpT03+yIAKS4KbSiJEBmGHU8KMrjgNLYfOfTIQDBv6V
5x3wrHhc85x4bAPhqtTfsa45AD5KMVcFZrcVPRPhz0xit7sibGfaMI7TeHYqwJVP3WY1vXVBdj16
Ix/yz8vHdN4Z5jmbzdPvEaslsb/hcxvHNDS4iZDdjYxTcfKFmw/DP6iu93QdCi/ohJMzEmHX27n0
DhDeVAVyukLnokj1JG6dGKcMtKQGlA1DVfz3X4CY45EJOe+5uL2v4njv7u41iYMnItl9PbjqVxJy
n7+bZEQn1C1JJAr62Ofgp9SQ/GlqcrHoGak9YQvVM3ZtinKV4qF6z/rAfE3z9id1vpTwJQSI112o
E16QQSCqcgIZj4XSbfHKgZQtnI3xbO4Ixgw37A4MthVZOXrWPLpes3S7iJlS61oxOEvNNmHwj+zr
zfKnAZ5pdx27tI67VsaAasYeHTKaCrWX7UKDf22wM9owY83qOWMraZUPVa7Qy/osyjHN3Y/jEooV
Lqf0GDL5p+vwsuyCXjyeSMY/Lg3heocUvx+AkI3pP1MgUzUpi9TLjV9e4JQKoV89zJPkeQK+MFt3
Tuq2H4OkygrfHF3OEPNzEGzV5FOKA9uAyNoTWTpeRvmtqqxGgGoC0vDU8bLjMUgqo8GIwz2WbFiI
zMR5jasRDjE2t7JPpeVjC+8MJ6ntGnSyGP+oBqdgrMst88wsoBiqof+0/SFG7+FxIIBXfSINDndY
tEWcf/IwgNNAO2janDdUlB0Usn5i/41CxizZoVhP9USqZOPmi6yAm1pZpfH2id5SNd8h9Dlh1Q6t
331xF2BP2dZ7D5S+1lf7Wh8N9RIFMgwqQPd/9o9lJDLqXwaNBvS10j4wuSzP+huqMXkkWqQuqARh
qNVCDj34XAvL3ojDO6rF0qUGDTuByi1a/J2U3psOx2QWHjofIjUqZKVwubD+5mMIgRcfbho2Ts9v
Pwo2qF5GaBVbIXZWhnjxzPFYoiro+7HHfOaXRd0hngEBvIFltz61UZGVqvsHLQT2OpXl9pdc0/V9
PWSJJqW6XScMavumfhC9bOFgIPJMoytgdCqZU9pWVgTkj4XRT8258hFYoy6WCPoleOfXW+xIKEYF
1CNJYzvrgU549rYtr/1MR+m9YB/51jnBpIu6V1HP7bSz8t/ECiWQV4ycvSXVUqFBI7FMHIHFUAhG
bu6kD6wsFEGAmhDnUtXZr4GFq8534GVHt/3nzyWUCU8ZrjGzNVT8sm4Rd/XS9cOjCok/h/dpPg0W
eQzXfUQzgZe/NxOhpli/RuVVwTdUqslJTme7iZAx0F3pD2KWn0vr1I6i6mWui2XtkdxtmLRFYxYS
Nk5ouGYcKLhDBH5m6ZZBVokAlWmzDHUxvK7W2ZDANrQWsFw7EjDdR/JcGNZJAqw9RiWjWsnRRnQ/
Ib9H1fdFkUWyexIOMiKoOr+fk4qN1ZEngiYO/l0mE7DwRXXAtX1G+X3PoYvVGmp3jKsCt8scoVLG
4SOBBORH7CZYxN3bPye0Sm8WhVou0kklIQOtjxMPVHnvvz8p++ceyLPzxJnbxEUu07C9gN2JfrL2
2ReMxlxg7CzKGvqfz2ATyobbclqaPA1td3KNIvjhEX2OXmmTHRhVXsf4mX40zn8tSsZO2ieyOrz7
HngC5WNIdIUxypQ0CmcC6m1ljPLcnOyKHCf3VrUHMV5DXijxoYaraenbpJKZf4RXh2ep3fC82iPA
rN0RnIgyloUkk7FX/b88i+Jf7t3S7Iiss9G04a2EDTWj8WVht07wKasXtXvcSzhyb6cX6kUczrND
uArP0sTWrygLYMMbpIiG7PjiJL2J4ZJymxaXH4vJuCetwFKhIAriWCTkx8ifCL/yC3O3x56bLUTH
xnRjkhcavMaUEfb9XfwbN3bxjIZtpzvG+nBusSeDyVGYrOIhRD8m49BNJahCulxiczCKyJnGBP3H
wiqgUg522DaONWT6SmB+G+f4wcFWaq+9FbJsPq5EDFtchqv+6GAYY0Wk+BXl3DnExOCWiI6yn4Z+
SSYj4qi6K1+gnsRlLOKVPopT6+rLUSEX/0/e6PWeIbgXujpGDUKz+kC9uaZGyxMk0kb/vZsN1185
Hb/56zPk7K6QfecD+c0VkbmfjoXLwio/8W0CsscSEFxR8o9UY6uTZl5Oo0cgoYa54QixhUuAjTL8
MVdKe87WePnE+YQi8zJhOW9u4hXSCVUdx/DjOZacR/FKyMiHANCUIoMZG3h1YNGMjhYSi2BE4vYT
CUQGoFrsYFr6/Tf02P24rHmJJ4ERiG1Srkyap9N0p1LdsBzekgWRAnR3QaSeewaXsvCT1X51yNl+
Cmo+DNE7Hm4iFHTQfq7bjMyPJG3IO5HDS6cR4ydLyPTbVSsGmtOy2qyfLyJw1dglBp1bO7ysUyO3
zuke6963O68foSN5mv+N8VfI+yaGMnDP4DFXcCAlp1i8MkGrS2jZE2Q6VfVfoiaWG4+lLReD+eHu
ltAcvMfMxOLPEEMhRViaobtAAr2EhsFdQgi1k5tXLD7Uye0ZooqSnoxIbQOOPNakXDO/abiqUMzK
B7IGgArpPEdJbBqb8EWLaXu3aUc92jPBOSbJicDHy2M2GxnCYRvBug4ZQD9KYbDrzL9XCmxtFDYn
CxjUP2cIN8uGk2TefobsV8aV2VvgREAaabSYxwvpn2riEbEY/ZoXIId/SUmGwym/TBAg56K6+MZw
g2Y2KN6IF0cR8ddHKT2XthnCgA1sPeLDyQdfl9uwqLlT0GfRonh56RGXQZRPoJ5yFpXZDjQ+7Lar
SBl8Zc2ITY4aw4/PkHTig5EMBvK72GfBfT7gIGr/Z2DP2ZKMtAA4RB9ob8BD3wxEeymIOeALoa0Q
TF7aFyAN+yHO694mh1R0gCP20umbhrO1bGza8/ZcKFC6CrDneaB+2Bj2FHM4lRkOV7uBRVWKjcdd
BZOXv/CDjGBYfdZ7Ur/fp3gxLRcesLGXw/WflbE5b4g5hEDGvULfQFkLmk83crlAk8X0PjqAvYbU
R7HSVtVaXGVhDjtcYA5OJ7ghCWd/7OTVDmiKnbLq8U8UGD0+J+O7OB4PtVPChaD7V9uIkQ+w/hlz
eSMDTIACCLqUZXGyTwSyQa+TWgT3DB5qSXe57FnbWZJ1hcgYZII/RaVJV4lYNhZXhJWGXxEsiRlg
NOl05OZKJS090+hb7Tj2cWkq80Mbja2IzrXI/6ShLimokXnqEFru5GfI+YVKqgcBk+3hw3UeS0SQ
7ZGawQ2YbA0UP9HcYK2ruWmvcQ2GPjw5U0beA6OJRegXiveeMX6btzAT4eJWe3PpQC9Rg9QupcPd
jR1NE6vm2gNDtWqg9gFAyoXMSHa+rYqwFQ0ymnyRb1qGt3RxwDdqHTrfKThU+/Vn3kHLaX8a2QuE
kHkzmD4uTnnpWNHpGxV808fMA5pRmUn6rwGRFer4xbWgwcGz/Jq8dz7k+uj8yi13CdAjy48S6mhM
1Ulxf1uUQzCuu2ZguzlE4g50Io9NkosrDRTI7N6R86k+Blahf0O2x/8WMulgKtzkgvaLG/X+0Ybv
nLbZWYNgC2CWrLmL/n6O1pQIiJ5aWsW4W9tG+z1nxatStoYLV04qqL3Nbyj+5ECUsV0Xrv0fnz76
lpA8qFCt7OOEAM6Gjzof2ZPvbzwaVjwr5FPK78/RQ61jig5xwLuK2LcLBdOTAKRFqnwdmTdTHgRn
WCZvICegltrlMFpc9R96MNS4L+S+wTGedAIZLln5df/Pi7DyaV+W9u5fQE6D3Ty3QycXqbr2c0uj
dRBiLgTBL7HuJZtQBgAkHXClqYz3DAnoQqIQntmpmc/Er9yYUtHnLbD9okWc4Un04b3HNByoM7yn
CRiyLay9pB4Cuqs50moRn1rikomD0pBg/sqtaTRsl88cnyETqZwuSsIHjt6l7FEqjBvafP9WHAMS
PtqNm1jLlcW3n1jubzUOcGradOTNOxJXuTBI/bDn496GA/kETSdLEDDxmS1pCBRkNMcxml98BT4Y
khwjUXjjt77TCbxGdJYW2/Aj0lw6zKCrfRL9j54Ic2qhxqcTgBO9rvRgONzRAMlAWXVn9gwvG8eK
54zTcvG9psUcLEWDjvLujfdmWMZ6xYVtrvywGENQ+haUOC3/JqlQde2jjsyuHqb+/ij2hS3FE+NG
BR5EEET79dySelkV4Fm6mwiRCqP+qTnGvSyIEF68WTDbA2s2YV50TyDC2ciZg0qduVv2aDN8WVh/
tCQS2UpngjM+KK0vxbZmHNwKrVpDwRCorn4rIG29eynVZBYiRUkt6hMDSRHlo32JzODgTxZIfmw8
s52BCVcUqY1TGT+6Yh1xTQrmPlbOvEuTjq7MCY7kqNk7Rz8gaYfneqxc9t6SIebTt0/CvX5AV3Gi
P7qbTYQ7flIECoCOHC1RNUdLqINkfA5q1slrAFnHmEtDNDq9P5h9jStIRuLujHV7ZVR6ayl8aiFU
2UDeAjyBAnfLod5E4P9MNk0koIOBFwQJur92brvRRqIiFbewiZ21/O7+0xME7EPHyinrMu0cmXHR
NWnP+t3aSCAAyGjEKr0+qrxAGlksI9xRAaxhVW2dt4Dwt1eKua6TlneCuuqeZqdJE6viLUCvH3RV
bTPrAaq6o7KZVnKr4/N2N/1TuoMzblC17ftAS32v8pX2IF+kQnKuX/wGF4lzP00oELCun1nVla1R
qu2mQnsgL4ITL58RXU0MqfWEOuffpPNY94ak/xxzOxvJR2hEWnyW9eOp6rH631iizY8lfvy+npFZ
UeFFMM1FLuoIkssIUAoQiqCKnZaR9wOmU/BUQLL+23um363WLR49XYZ8l7/Vr+Yb5u/yWRwDhDju
WCLvPAd4beqIISON8SPZGFcuro4tOcb8jdniWE86xkO6z2pDTV5JVq9RuwChpCEf13xolrtYttE8
Wl2LaCKB9m5IHRLrxUlSwCl60mZuClwL8ECPTnR3jTXuQdYWKSjorZJbnG30PNUnSh9QE1oMqazs
PqbZssOvSG5RRONr5RlpOBxe5X3mAIM8TJUDUJ/vZjAYsM3U3ggkpGFQzypw9GOhoMBIcpWANBtv
uL8I3cozcvz6s7N76lUSpyf4nUOBW08YQajhF9gn8vSONDm4dIDngq07qjkjKrMxYAWFDFYP4wSr
uQjvX5T/+9Cq/ppqaQcb2tLLV8B06PcFj8+NpBaHYe575nnnvr1zA89WcR3n8uGodHKRX9O7KICu
yAkmnMOoakd584jHrlBCiOd+fVIuZo6FvKQxJ+YPQ8r9HuMC7x3fcRZcJhD8DoDXMRdrLfxaGnU5
Xp+3KTZ/SEZ+wL9WcM2t3KzuC/VT+gR2XTl7uE//G4Ips/a4Bm92Jwsj8I08QCFUVtBb1kEogwSy
uVdVzgtCjpHOOTv2+kRI3HQFbLfxseipc76CyGpttNeaPUmi9WbEUTnglt/it/3/Ozp14/SnhLPJ
7icUjew1+Dh3e6CBZZsJ6819IrvSLARKhpxD/IIg/I6ZQNWHdR/wRzjUY4s9o67JFIUcjmcgG1FB
OCc8KGKP+KnSsBmyFZMIiT+GsVV6zrjDEbmY4WnMvfgw1lb68zz3MPTvd8zcqgqnxsbw6ih1I2ye
PzkHz15+DP9iS+ZNktfX+JdFC04pPEvQPf9QUCd+fdjFbCdoY6znbQeyGQIGeMnpxGrA0KEyXPNU
Sa6w7QUEnDakzqZgf9vDrqh6E2brTmDS8Au/LsZceAsoq8zj6jfh2NMOg6hUxebx3Dx9Irg4hFHL
7xn/w73ud2GggLXXUvnQJVrAjDd0hjdKz6NckYiHYPyRAo1OvtmVoczGLhFrdBjs4KAEu8BeeH17
BIrUrEa1In+PoGM6stzzTTky+ktYAikXLQZhdrwyuzNVrqomNrfApdEL/NamPnWpuUiF7+T7WEBE
Ij11XM8Hbeet/67gHMz51yFE5uD6Ll7gocrelBJ0ai+xzRLb1DRaTsYJtw3e2axiRiKqNKyCeDeF
j5YieBi0HlQysOYzOGx0PEqUOQxL9i4PQGg03O5sO6Q/5cVwwtBF2BzZuHSvuOGh0YxFBXEY4V/S
Xc56P2O12A7XP1qI6rXRWaJzUWFFN1GavTH+EzPLmhuT83PdiSZo2txAgEzyglgz8zcZokIFb4cc
QVX3EUiXrjzpQl7as0yas4bzWD5UQxSl3FTs4qv8jDGeVcbiAkAPunlFjrIHmboJe2TcjPjZnBFL
I+XBw/rpu1898e5LodHX2c6P/x1pbIVSPCYUC5PYwUXJPTxyHdhAMlZVvEFubq4q5ItGLF9MnbZl
lIR2o0dWvxbIqi1WdHpEJMbsOWzw5yvWUYeck9EHkRj7vVl1ZYSYsIgqXPUYmBqZq3XhkVUvWWHr
mtOhePtujGFd5Xtai0gez3Mct0pwfKRDOW8YdTATw7dfAB/02iAODuUN5MT2gAzqWkYGWaR4ZY/H
HX3i9jJ2JdC5eWw2pqVD5f94GdxVVk5feM6QnrdIRw6paZ/zDHFgtsOYacGoAHkcM9OugJCEzvwX
S7jdfu5s8G0AxOvvw8RGZK+uicqYnZFeWbyEg29cQiXevo9IXMXctmSjVDCkkmyKQnnGa8WbaJru
GfT1WA8mcFkEY+PkbKJ1c/U6AVS3lFw5+BPBAoMhyENoDqyrjT5l8TQ9HqrHdCC0ZbOZsgWjvbio
wklQXBRmosvUUvnYlkmzM/OaKMwrtavRENsa4iCXwV6tBiMxP+enaRwvLy99NshvaqnCw93olCTs
Xg2Y+WlxTEFTcz50gzlGLYMN8/wCHgIw8DfOwyLf0drCtGqnigizFEDA2wB9kb5cK+X765XRcomn
n4uNQm6HyCZdy4/L0FCenzaf+W3O0ntAhNJIRH10XNA3oWLqt85DQNtJLJvu6j+Ofn9RZ4lZC395
OexOGg513l4PHrBir+s0r6kfR47FvVVjF3ZQ7EZB6o6jhofOlmqGQihVCF0VqpTrbVBvaeQA168Q
gRPs3PqYK9kyjIg/sTXyAvNE30njpWq87wP3Nl5RJ1G/ykOKHt8V2azYim+DJQ61kAZ1P2y1ooai
w0ZlkUjQLsiMfZ4476VJyGwExwDNH01c3CQjyiSZmZ6Yqhqqn665o7ckKdBhOjILclFcxd/8r7ZC
gnVC7o5IlhAby2l5Z5iSBs9UfUdpoy8UfC3VI7K3TkhPK1uDRhCjyH9zuqXg1DZ2HWSlMJI/mYqZ
sMMtgLtWiRmUeMImSlp2Si5Nz8SCx+oHChLo7C1JK/4frLSptag75EtvmXBSaBXHnvH77suMFbQ3
Ur0wetyBER7bMMBrLcuHHPglSaBDa8mU+gDG62K9i5LEYZFECxHYbyyUVu8lxYoITZJE+p8OFzA9
7PV4SWMMpJ3EiWydQOSSR/Ki5lNpvkDz19u6GdqAXZnsA3G6wjttJq8JFCx5n7NHwC08A+VoY9RT
IbooIUr3VTKcP2JFWvmIsGoHkudxGWN400PrXIouddtCS3+PTgnDN1st9pye2pIVRCg/MtAEt4rm
Eg3Fo8rXcKk5UY7zvoMrGErkhunIqwm5VTngr915P2uzdD4/3SIi3A58W3fyR42KME/sDuadbn0b
cPGwDFSvBQ0VdGrMVPGviwLqIfkwa6gitlIIQ9ufJzOMrznLzXSux9Az2b2jkAWktWaRG4SOJYaV
EtFwWBWcEPfA9HpQEp/7WJjyOqbrBqV/U9Ub2zZVYo0dhhELvtPXuatsLhPdrIRKT4UgGzoZm962
rsaiOIB4//ERh6SEfrLCJAiHd1i7KfVjHC3N/2zxxti2kBfwqAC0Z7u3BYZUbJGKq+ynqvX0Tugl
xpMFnq06BQhghEdzMdBwKkmB4XF9DY5u8cjmQc42YeL4/j92YzlAkt/RyMGS8Yg1/wX2hyDykI2h
mXrMacmGnt3eOlKhYlvIySrayUz2+KH2X0i7cGHDPXYZYU+mJejgVxoOA2UvsOhnggUrO3NhqWv4
CE7u0gqtcgVPJj5J6VBDfFgd05F/wYLzTxmcTCeTCsciFd3eFSZPl1RVrhrBDJ1Agxv2itEkiF5X
Stny0KY0uuMErNxmxz5pWN9Q/whtqIowVvZ2W4bUhhs+hca4wxhG6ehGzxGX5yHSHhFHqXYhoYTG
9IpWZK56fdqYIKcCF3A/K/J2saHXPeNKCtgutRAygc9jygCkAg8vmxM9K1iYc5xRryNsMPscka3G
gOilX1TdB3t14CqM1vW15Efzpg493NYS1BA/STv7M35RW+LXio5KuAyHHynwADhnKOVStf/uAgEH
KXyrnb92xZE4kSkjzRkNXTHexq5sIVtmLcYMAhospFOUz24h2X7KG05blkPHC0g3lPyCn32k2vt8
2wQEAgc+KzD09BKUOVtTkYjpsGNusZBiX6t0JhgCl5bi57ZL92fdKiyrtQ+i2/iIUB8g0hUazPcZ
u4ECEHNaYPvugnrSA4WZoJP2JC1eBXyMyiaLJzI0RsDmN4CkIWe4+BF6neC+Wt9oiQ6gSj+gUFy8
LKpPRrjzpPDzZGUtMOSesBGLOqDGD61p8mdQiwuHo2uS3uweCr001LnjFSt0Wlp0L5jlVd70xLXc
VmHaNHfzTuIO5FtteAnmPt1TtWq//50wQ8SYx2H9GCaYEIKxV/eyCNSJehpYBLCrdul8vPjKzxdk
UuMZBjau8vUBtZLzlLZKQsZKSppHnr/grHb1J8Y1/IaG4f7XPBz1QS/bdthZCDiHKyH6iEBPF0kd
sSvpeBtyIjY4H4ahkPB3XEuJLIWMF0CUEv0aqQR2rJza5zONFu0unArC7fvq9ie2n13OCBWRye9b
4yKNHga9zabH2P+N/ndrh/XjvmiZHafH3pm7SrfwJI+aFkvPi+fAFeKoaVK8M9FwnI/Li1NvISz1
UGkGRmEPzg162BZ9fCjiKV4foz/dJwniHSFArDujmmDSqIsqI11Awnx/IsS0ZfJY3KQTJXoDfwqi
EhIpc3vBntfajIHQEy7CmkJOD92iH4Pk3qfS8F8quBA86/SPZi+japU7cgNXDlSJW5A+FlGAWWNu
LgJV7zvWrl3zKVy9W/zwVvSeNLbTZH5VUazwTktAW+GqzQkD+v3wlLmDv6tRKZUANrhhc4133fyH
/3gs0YLh5PgzbkSQxIjJjamx14yKueYQw2NL8T5OlgLGfwD+GKBE+IPmGSDEcBRiPfjUIsGx2Oy5
bpfGPgrIHVM4atRduKCzjvNl+l91DvSnlBA7yJf65dGgful2FjBIIKOhVWYBadH+0LJQyiNNT2Ps
hMHxhYRs7k1XF/ifwIXq1IPcfyx731WOQ+ODNGIVVyf/IMFrtysXJ7zh6xLoKq6ArKSqtxB9E42k
HDkFy4TFhmhlyt9QkVikVNepmeH2z/RyXTm2OVlpWf8h1TOZijgdEINOC0L7r/qB4VQy+872kuba
IOebYzIj4dP3XrErLFL+7ojeSJAvf8P9FRIHDSsbTfjHZ4SzjgUYAUnFgR5fKLpkuGqgj6CTzKFp
LfXlfBzVkR03FzOdXLxb0Haemu4P5IJQk+9h6YpmHjyWEaezMmpgXBEJxhHcvHMFWe29hXT51OUe
1+3pKi1LStb2qwyTZIu6Yn8zKi/XWcl7CNreYKPXMmAkx1pTbykYzfvfO/lYeAm8r74E9kpb9VuG
xs0TDZdclfwNRHPjgDkjWoh/xH4QWg2C+zOdEJqv2rexPnbncZ0w2uu5ig9jo+T+0PmKXB18QQE3
TTxNsFB+O269rgudvAgTYyhrkIZ+Vq8f6qrBLYgQgJDdUA3JrU7csKori+vyQF9/GHCdVqjSiJBK
nkKwBBVLDwtl5oeaW9jUwLv3t6C9oFBotVC5V/bX5UGcwlw7l3tp0efrEbDCa3PmFYltmT+uaHGL
BMnPtmgS8DKVIzZtH0RAPvJEhLewDmW5Z6A3+g7Q4YBpgUmUgHOMBNr+rUTB5FeqKxrOTCXMwOYH
Az61nrxOomU9vzxxgk9tp4y3p6JnkyBEPNIcflEEMUytPOi0uRs1lqfKalQ1It7568QkGHiPJxk9
1NJmWTxWJQgrsc3mDR34si8QXhg/Ikz0pg+qRmzqs3mnQljnO8sOhgGpyA3ZFDZqIe9KNVxcy7J5
Mx3Xk5M8nDQEaO06TCcZscrQ090t9Ce3F7zmmD3Vlv9IbidUThNaegK/fEgvCD+iVSDqXjKXrZUs
LxFjgdUz01OWN4cgOkxJffGOZEhasYKn5aBa37l6iwrwv+n3bz8+1lmBZVWYUQnt5JAWRFiTvZdM
uO/lB+efe1d69tCglW3WsOWew4DP41VRXBBQ5wLy0NyQczDyvZJ+w5dsYfFixXA7TyBtMtNBhA9N
rl48voYnLQtubBLWSeIXSdlsQ3yHItcPsaD7S0g9oXU04gZoYNAgnnvE1AlTLoDa4FS7HqDDnJlX
vosTHNdglngHhSm5TZL+S1P09kBQ6MopT/3UW8bf3jU+yrE4D4f722qBsMSKvnqj3fKHPPi7N39T
0U98iAzZyQi53K+eh+hbaOn2gbPrGzaOE6ivKcG44sA2Hr6jYkmx7rQUTM31DhbmozoZO/sIQuoZ
ahYhCvplx5bh4h2QhFP6js04bQASbMBeaYX+o88w4zmToWPxIQ25q3gd03wjNdqFAV7Q4++BMx2T
J2Q9SoZOUEsLnjVJ3mhIY0k+K+EJubqSF5cZU4Q3m2Va/bbVJM7qGjjXHXskvzsYAvgcVMBl7DdD
ntm13Y9Eh3CWmVrnP6nEDWwleJ312iaBdYmxBXS+qo5GWdD81rC+CPg46gKM6bkAR84G8JtiM1gB
j21sek7QTVdFh4V6aOLu3Sip2iJQ2NaSXLT/q8tZu0kU2pGCHIUmrWvzcMSd3BKQzehOD8YBXktU
KutDvabYXXoUCo70YcsHC2foje2Gw3cgVBXisknQNUPPwM74wTbYVKKn5V31VcbzX6ZVWGsKDs2m
tmW83N+dvMYxtwBMgMt1a62ADQuezy3TM0yXUktsXLWB/hgV1eraV08AKqe6jfL2rx2fK8BUG2xe
Q6qODXw2hJAAwyDKLcq8eRXNn4PvT0j6PxjgUt5oprTPIW3HXbe88YAkPvFmo3h37OK8Cs2rh6Ma
OLFxb5On7JfM/nia8ekCdn7V28ln/+c5leU2ySfgZ9IZkUWJkJszG5YRnNPDwYMTr1cvMHObbLFQ
OH/evvCTNL2OkfNyoSczXpDz4UTbWYNh9GWsAjn994QOXO7XKz4fEMH5yYydjFMCi6l7ppDf3ehN
1LG5TI3YG9czPDpbizBKk/SorWfCGlbXcms7KgzgnzK6WwAlRirv2BS2ZsGx9FWJHPRqNSLhYUav
eE9c3qu5dd2C7/KRpIvFvf+p5aGhvnW6FDic7SDcQxUCKgbBmKexjbgMD55qVW/4RCczJys58uY9
Ooqy7fMabaF6EslrlU0w2U2pwYvABSZjj/UFHbAq6jXF2FlYV8xOmC3hVebKP8FyY0Ajd33jXCar
aEMTCmyCjGh+nhoTYttj6EbdNdmAdzoYKRKgrfNDtTtfgRtWwSnIJ/F1KVUegsRzfnVicW2WwFUH
v1kdg0YdsXTyAIOZeCxjmVNtMqJfYsOougqdRNIAZM/JMRDYrh3t7Ezz6b2KsY4QM1h/kfjUh+7y
NtbLae5POtT9rHwDjIh+EpaNqUigPxDd6KHtSRmVefwGTTLAbFlGdGvmfgo0u3ngp9/JTn065cn8
41XyaeiS5aoH8zZWhPXBXmG3z2csVkKcXGmba55K1QYf39CfSQZjBklr1BIvxfGtH/o6AL1/1DUU
dQTtaG1zc736+Dw4sTwlEQRCgVlMVKKn0MsnaOlSF8x4B5wjReOu2UnuA91c8I0tWtX0cMlwPqRf
A/wohjZGhAGysCnOimuPzEOVFh9F1S1hS8LoWCcn8hgcz1wZ0VrraEoYpqgacjT9lX75YLeDvime
77z6RxWRkEyn6essIMxJgsates8M4QKOjzIa7DOZPWbi6HMeJz0Xj74S9kZMSknL+xcB6acDMVPs
2ENhVwr70wDNe+kqRHlAVkMiXU1Z/MbqCA3kdm1VbrtjfnATPN+gR6F0ndHWZFXIVg4MBjx2ihDr
3SeMQgWRCvjUD0jReyzFXEmxBp2fxaDKbB4Q66+rPnabFO96KWPQ3QJIQZ0PBTrjxe67J2I8VBBe
ENaqhLuNvPjoXeljTN9ttDnVzd/cULoISEPiGVIJe4NLPlvM5VGIs4+61fKXaKC1nwVfnsPXkb6/
VhyZKML5TatpygKHbnexx8xl+vO9qxP83Cj8jMTK39yagnEUH7mxL5uIM8F2ld8IUrzYezmOuazW
I3hKWzy3+75fpyexdOwmJvz9fnRGj/p1u8jtgyd7ImROGFYTiysjjMjczYGidjI4F1ttghAj41/1
zbypOYEAYtno8b+4V0MNVDJnJqBI+ONXBGFCR/bk+m2wyL+lHbe0Trie0Tf/iJn68igmfNhFXmQm
hkQd3S0aZtM2loLCeEy4XRe46kws/G6dFqSC/3bBv7wQpoTVj+FGljrRBXMP4sKY4fSWpQtN5dNa
byyUy+XJwLT9+KitVrYj3q4BbjabjPyYZivAJQf+ZTBD3GSNH98RkTiIHqc59QPs56FOA8J9tzMp
45hRLNC0A048RhScQ7vhrSXN6y+raFl/gwFbZxBKd/irgl02p5PMF/1vpLs3N7o+bdmpRVDj0or8
dlJJNCZvBMWXsFeh0qJUiF93TCwLtz/ZIDxGDgNHNHO1F36QkVVwQ+jpVsyBlFgFWvetXAf9vLYx
LjnvZ7bpxjw1LJp5nOJTq6RAGZM9zBH+EApsoTz95smLMaa4tfPy8LDkaszD5KF0aJw2Xf8ddLK/
i8W1ZnLDwl6b+4LDhBwrdpaA0VixW4ffsSEUuGAYApPHHkoAFyuvPGNsNlAgrramc9mdXTmNi6U4
q4tpBZNepsJLsv+Xu5W0wAIAuxDH97gQfKuw2JVXrFUFU1QV3ZgacbEP7uE+3WB02wDmYMcFvyFY
Yi73oVFk2MJ3lC2+y//GnrZLYT9WQN+Q9KkRSQ0cajJGJnlYFI+vkqjU19w1u9uWtLOUZJcF/mlD
xXkpcrF9t0Qv1ExHJ6w78F0tqaot7pizrJia6eTUlF78CPdslmvELvynqJ5oX7EJI23ebmc2dEhM
WAYPwi7LMhHjq4/W36oqQVmSRftrI5RHJOTnvh8L20TmhycEvXwOjtYPkGGjNjw903nYcXtgMk6q
djlLje3PByvQO4rp7EVmy5L+++UWKadNt4Djdd5kUH8js2RQnIHLArq5uy+YrOAqFjb66WTHWz13
ZiQzhjDT3FKweXXoL9e6iqmHCzVZqjRyWKyvCkZFaXZad1UoFEAazDkfv0bjj+tiFiJVxK06Mr0Z
qXr353qD/AGIURZg9ZCtL7p1OHmf2b+wxvPLuy4PUFgU90HExG4AD/r8MA9X6uCiD/pVaVrHVrgY
rgzIEKp4YCrI1vghDQgjia3YLFTyGzP/4nhaa+yCklo9sFq6oYSPt9wDF0dq3HwWeDzEcuJPX0Cz
JK/Jz7KbItxbFvemy5x+5SCJTzEJbVXhTh+52BO3jEbam+wF+sNEpdmGmQVxMn8cNxqJxYE8oN39
mSmUxA0UQ6XLfsSARTj5K+OHBdXAWkHYcnEOqpwB4X9ewi7jhEDVUNn31NrrKl8EPKnrMQcyqiS4
wxZ/oNMNwn/KeevA9yIBTG8oKaK87BHbmHWWDaLHsdGexyJe7d0ixsArWPMUOunjB6EWPaemqmAn
NOvW3i37l5APd9ZINobScB5ZSpULVZSQlnP9DohwGFdW2JSwCJ779S4ympDZdg8Z29QjeYhBkF6V
xzLWaTzZqG5gpDtuoqnYvYhtKRU3UxiNIqJULQrVyBO5dw4NCwXkJlP6XMyBy0Xo3jFNDh0I9KiC
Jf12AArbKPJCGs3FdsVasatvh9d718Nu2buOQcOyGKZi8qVPdwsfJghcmISd0ixYs5VmGymbaJOf
KJgkkjtPOptCwXjLQ+5j43idCcYS5vYnW2ivGWUN4XlxQylHUOYIqiSkpXuTMpdAnQKOepM/ApMw
1az9d3VFKQ6hc7B5leA8EOkP37GWAAeU4kS2VlP7m4mePE1wUdXR/sppTVuejbAcxmI/uUFHg73I
zwurLRFC1Rh33Q0FGNneQh4PtSbUgmbClA3+cA3bv+mgMeoZ38mhyMrHzWE7cpMxTFkBxwtmyrKB
EElrGWy0dgh2NN3ATxy6b5gIiDqXUTGgZiWgw8nX0261CKnql0rxzYpQRFwVz8DFsznTPaEV21ju
WW0bwZjuPlYfzBbxFV+61JvdbQIxvgZG28yzMideO2s0nawN0zQ2fxkaL8XfsdZLLtDEGe9J9JB/
+UmyWpZz0B2TD7Oy9dTSZwvJ0t/AnyTDnke/4UNypQUbYVtDTLf67hsNIkaLn7DcTXzFMePynuof
0tke5M8T8c0n0YrRLq75UpqSLDVosvoAKpfMHSLQcfRVY1Wk82J18k2V4hER05g9uYwNe4NDM2NB
MX2cJFNKpu1emCTB4dOddxcNQj36Y+vI4iV50KBdL6fW6tjoumrfdDgulIApd31q5NcdMYAiDJQc
a87iS63X5LHD45y9MuAprHF5GEQBlb0bEiZ3LbRcebOsSTufScurEQrDyWYJVW4IPItx4PHzQOM5
SpLxyY6xFkovjLdrtkzPEl7TD7RQKIsNXy188EYheuM2otg6W05d8hV28Ire1qW1kw9y43BJoDNe
rSiK5Yve8IbqPzjgx2GtLqdZUoYPEpqCXEEwACh6xgoczYe5zXduq/U84SjcsTG9VgLvgpRG2C32
UVF2UafF6rGX5ysxL9MRsW5qtRyS8ucSAUiNtmvbRFAf/NuhO7p02/1uze3NpycxGzLhMsZn162f
MB4xlCavkdXzgDtARhfzSHAGc9MtjIWIQacv4uYQjYn180nfqc9D0kugsbkYkh8b8hBxrK8ckgDQ
H5/NEKmiVf73l0U/HkVRhEOfcYt5QCuIb9gqFb+JN6kwq0kjaXHSwUAxZTR/tHB0ZeVzNLOxXdkY
8m+s/1LCgBWgzRTegdV6pMRmLjVDfAzi1aPMaiT+mmFaz/iDGeKp0ayeG/3EpVIUgGVZPRRhEIUj
q6Z0rhH9tapRasoM+ykCgbnpkYwxlnf6EzgxWZgJRbXQWCiC6zH4EPqn5c7i8JTplciweKCT+2/l
b96pRFFvarL1RsBTO7p0FVLnoxJBd1gbcSIMODIurngOKh2ObWJkV/QTf7KP5DR3GlLZVUpyj79C
L4WLY0Z0WAOGjK0wW24VnQOnNH32cr3xNxVy2DVEXoRt5tuKAp4eZfeenF2TNiB9eJvDEmxsCtkL
2D8eNnNbmOygMQ/t0cES7yyekJyFiHCtG7pFlSSq0swswxfxGFZu2/PLSxfxRyXKdRl2Hq+lz+GC
7EDYaAr8GdNkU/tdtGAPphObE0X2TjnyOfMydaCe1RGn5ncaujQPtB8k6Kvu9bk+eHN9s/grQz9R
ywzDmLbUpD/0Cg3ee4hVw5Lfvlfv8NsDzAVrHEigZ3sSZ1X4/6j/UkBKVe4Ru8IpPJ1/MWYQ6HEe
ap1bfkw5o+84fCPzyMF/EOx7HDfNfJKxecRIi/gCtb9+7spz5fGy4cxKuKppb3r0XnmhnvWCZbUP
9w81TdXsvnJlNxdR/uwyPvPpXH9UBgId9QhJs9yJtnYCOhcsCS7Qx8e6nd/Z9nIcgHbv/UZC1awM
KnPjacLiZNzdb/TUkStUMn0fmOOc7kcNd2u9aMou2Rm6/Tru201hXEgVjIDQhJPeFm2EssIGAz+Y
AVdQG0sTxHqHOUuVaoEqtor7IDgEk0iYab+zuVdsiSq3UffVMg6WkbXIZoQJ5xISfLmxI8msR7pb
xj9P7A8DM/ftuyN/fCQy7wufLJWelnVLniiM3n6D9Qm9xB4xq1H3JF6jGnHoOt5rFtG6T/fsWBhM
1H0OMItzkYb0X78xrDowntVLaUKzbHaUd28+VKvaDr7m59wyx8khu6adoBG6nh+kZvcMccfgugo7
JZzVbxmo7iEn3T2eVaLQ9ilWQJxfTVODSgDdunaDvFUIcDrEg/hxCe13+V8NwGS9+Dc8RFzuGXXU
/sdOH75mQBNH+Ye7AhLYmuW8gFtpKG8mIrNHi+bSGV/u3HpJkK8QT/tyAee2hOQeNq3s7Z2a9PE0
cDkW43CX4UP47QjmcRNSPvdpPSXZCfBMtk8fXLUjw88Z1dJeacyw6dryTzsURVGXOD5znL/ZkShi
CRelvw2JXJXb28zFqIDCRwz4135ghJjZymXlKRHfhp2uvXxDTQgZPlMVcGu392VHeDbkOG/4dfe+
GqII02c8l0nkFGp7YPspc1zUt1Kc3yFYoQ+3eHr0i09kqz1oojx+ZxPeTC11HpMqa0e2NmbCmSBr
zLPLBnvgGp9HqvrKSDQ8CKTOSQb9eWgO8JDj40ivH0Z+r/eASESftXnlBT4T+AVinavBsIEmLhcs
N869aBDSvBrQ4mU784i2WF3YI9fCLJ+PCXx9+iM7HTNi6z72YfGFR7SbGcha8ce+X1sdLG9PxD5V
qmtMRxEIKwBMIEE33rKfQB8raDU8FWCPFYXDiddVzu++4x1N2Md/gAlKX3rLEXT6OP/gI1K4237X
5UxCnLDcf5LBHvXB7xjqGqdmQ5LRrxHivKvPBRn5EAY8cfgNOmIz0Q2v1WM8PLnxu44QZRG9mU1C
yHOkDw6vhNhitlx4ts7Po3n2OwK3LdqFjgA/eYGV5RgBi06qpGTrBUgPNusjnoEee4lZLc3A3nmP
u9cK0XN+DKYK+2hMUJ4mRHB2SC4CK5im7Csk+9vkDEyd6As95UQVor0sYJSeT1JcZXSuJ+6yx8Vz
qJmCU6S1osILi+v44PPyZKhBNvluP4tfvv8layUMUtGR0iR0avJU9ZnFrg3MwgBzFhdUReBSu9NU
YLvh4RniP5fEFKzUP76VKOzI8z9CHapoeraGlFQ72fu4ldMkL+nVb29abj0O42NPzwBq4v12JYoE
E5lD1oDef3vyNNtED0JO9kFUlwQil5Ttg5wJZ4uz8c4ly6Se6lRPXAPQfFb4mZO9qHbh1/O9ro/K
XunsnvLtnXCfbNAJd5oPGNS6Oeoa6j572T2DpyoUO3loGAv/vWA6pogMO1qDX/PmXkma40Cu0jNT
vAFUfGuau8bKkRJbWvkpK3KSorHuYSF1V5Kc+tIfLfwfWjUecqnXaI+Cj6HmnrO0rehBIdH/2Nob
FKcb/+GtaxWpAIRR+QNvFAKejATTerGKmeh+eMrE30X0NSYeUHqXrm8URV1nE/7YqEx3TkHV3dnq
peFOzZuFebMGCY7pljJsS4xFbPUbsmK7+V0lIKtMUsQbLdW+DGW4uc1z9x+ZlUkuLgdmENOfvq/5
JGhmEuFAOwYUqMgF/A94UNa2vw7BRCrKNsMk4aXup/6mTBPOSRdwUD/u/IoDubBiELqM9DctNrvz
LRPzcfTb2EjRfh8LQDNlayOM1EO7F3GRfuHo29YDd90eH8aqRIqEv2RzMFt5VJ6PvAI4PKcDsY7Y
o4oNDB3yq3SerlkmFxNRnsHegXeXcoG9HvH6PPirFfSiNEQnClHbfmrfJ5hfVmkIT+T8qWkjvWde
xQaQquu+CV27xAxBhuDJVTAQhvjFMqXRif4cieiSksfcPyOUl3XKqXf9rOccCrgk6oeftbtTE+Ce
9kcYUgptRuy5Lt2lhqDg/TZYV2PiCojSdrHqReXSzMsLJ0tIFSsv+2GNwvvp1HTvL/Twhm++9WPV
kvj4QnW2ITX/sI6YJko8B/rk/VsaSYm1XdSsazOETOeyDjp/jxAOBqhchZNOJ7MxS8dMt8JjGS27
O+kRAzXTTFZsFP8BpoYwBB+ckdt8pJhEKC2IlxUCDoMdClOmnmk3aPxyhp1nCk9wBGS57kg8MPVa
HA5nPz2ARiEYkkFuwz3ms3xqMUv6EtjoNvPft3RI4C5uedZfklmk2hB6qZnWIjWR9yYZW97Hmn6R
lNgiHvW3DMaubREvHUCTYF4L2kU5XGSP8ZqcTwCUpS+bALh/rnxHiY7BzcHCUiiQ75b/FxTt9Kqd
wGQyJOXIxnII4+S7K289nhe3t7vg0JgdrkEX9tLfikYWn0jLA7OqmEg478iRHi4rz2Y1bIe/7zq+
ZKynm+6gUWBYgvVp9Jc7VO9oSumvpC+8PTvsxFP4LF3Uxtttxb9Bp9/mR0Z6tS0OOalVr0q8ndaV
zv7b/rIuQSUKbEelRiobAfCP83dE6T8yYcyxBYFHun9qSLwwpf1dMwAwwAPeRR8NppXSC3OwG2Ph
brb7dnE9uEH9dgJ2rOqvjT1ZaWkzJzbAA5jFXXcAuUlN+a1+zoOu5NhuUx2J5apXe+hW5HLB3/m2
lzqiH74xVxrS23SkaRXcAIqU7pe21Kr3Bl75pyCwd0Lkm4cDWM6ATH5HR19hyo+dkWBsp2Ug9Ap5
hKowWsUstTrKLkagcWR1gVXPP/cq0aG5iwV0ypN7/v/olFA4z+wwJnYeocF6QXen18anePXhXO27
6bxUCQkKmv7iGNYcr16Vf8BV8QiOK6O2EhQIj9GE2I+adtV8pAa1y/V1ibiiyBcdBksxR0IQbkw6
xhV0BhhDbcoKTLvXMDfdPY9weI7cejWverIrEGWSDJw5v4pL60cBdxN9nIvSkqU9miIJ8zXdgAiH
KaUk3Ovy5mFxtF2qM8w5gFFQ6rQUp+MH8gG/y4Sr3Wc2QwdyotE6ebiSEVzOorP08/orKx6O45e5
Les/jQQkdd799b8jkN6T6ZZtl0Gd6ipCafOHyUH25RJaES5ngrXQ0m0th+RSF9j1+1pcdVR9QPnd
rEGCw3p86qC3k9zxTZ/YWT2e0Vfq8xwNOyGmiyaMIiqv/i7B7Ze/UwBiI2oAr2b5XRNCJboRi2dB
Ntuy70nPJqrxuZkMxI3+YeNk4eP8eckKxIdVAKaPAeq8Hybw60HBeda37uDWyePmWsiIoGpkxq0w
vnraTk5s6lS1L1GUvvkDGD1PhIzJfegairL3e33SEjNU0e7q7yaRkI6Ow/f/HsMGfg8PvdNx+kz2
/R9JERbcMZ8/RMeH7YsdXd2cMtvPetfpsfXyriRczMu+sKWk52XzgsrzbhVwi6ZDCIkT5G6YEaWW
IGUViQwKaLMMdEcFUvLnqSmFW6HjxLY0d44XBpRdg74/olF10hBXd9L7Lp82h4S9Lr5pz4PpARPo
Dl/VzbRw9FoSLoYcqtNrFDuofthhtR2BBPjV6ZwiZw2aldmqcktLAnkTK3WRQLJeH6SepCs6NVa1
Eh2LcGFfqBAqnYJJB22FBZdhwlAmMcJz+ZUXN/VR7vHftQ+7VWdks+RO+d8CrU/qP63eV5HDeanw
LfBTGAuUNcuIX269HyYygjpoKKTob5wyHQjDtGYMC/rhILPiRSOwA9b3KWBlFFPA2RkwW5rycNnJ
iTnaC0gL6RzETrNDOCHzaqtZ2Ay77Hkofj9+OP2AxyXkNhOmQs43naC9OY3eh5vERSRoRwKo62z8
bDoI9A+pm7YtTyCIDdmXNSGbpf/jW6kqaltHZ+X4W9JdzRlBwUzbCsv670RhjPUTQURCxdiM/xK/
K+Qwht+V/Abj0ycFRZ+6VVCRZE1VF/82eWmb1IuBvEXDaIj9R2tU7tT2It2IIQvvcvULi12h7G5Z
u6oM6Z+CeTQze5Nq5SVM9yW2RUqxUkqPn4EndUGD6bvPMk203DS7WxjjY8roqRpMJZwLRMuy4EFf
jSwk0i8GXjTyOg41pNYNylQuG3WEryuIIdV3FMokJl/KH9DMp0F8csUkBNFtUt9ljIYY/7qFkIRz
MYKR5B+PspIg6QeoyoFYROGisN6nB5PG09NEzkfbv9vjuaEsXIvFwq6JnwIOJl/d1Ei/5pqn+QP5
9270KZm2YYGSrMpTWD1JeG+Qi2+iaRKR5zYtgr+JBpRqAIZOgAccv1btlSIlk3nQZt8OjsmtupGL
hx2OuXp/U8rId4XlAU/x6FOHiFSLkiPNLehz6xRlP2SzdBdurTVsl8+e0au4lbUsC5mWuTT/RLxw
IbhZ6hYyavxlMkHiJxad/nwiru22JJp9uHw07LC18FtkJXNddP4/GGqiEGoSXakLZi9dwp3uJ/kh
+lh/Iuwgxo+dtkkk2l26pxOS7qKnPKeYW8NfdzAPSy/8NSZKNriL7exyyJriP6X9RppJhRTGajNa
9CKhWKkPgNac3cy5aqzzR1Renoh545Fc+gO7WePlfO27RRPIu3O9dkM2aukf54SjRxZkHhMdTqYc
HIIm0biLKKRtC5Fceub0E0klXIIfxW4TiAP3U028T+VFHCyynsA8pji9avJrgCbt2e2ZPRfT3JJF
fx/J5J/V6beVKrRGYl2S7nwMy03U9k88tkkWvlMKg6AJ6tUT7wzw1IRSuLqqNrjuuQV3Z9ZtVzXt
jfCFBMkqqhszw8UTY3AlnKd2w5YtB+Wx3vBWyzIC1P3EcuKERtCSx4rziAgeOlrsx7m2IAPE3aHf
a0fywq5DfN3QW4hwAgZPcj6R4Pi8y8lug5MCVOf9DGxWNcFXYhP3/PCWREaNtGITfqpxvUftzGR/
EWh0dsXRNOaZLv8NQzfXK1Np8A6sU8K2Rr9jdmoBwITe7ewUWZjetcr5QrKCxDYN11yzwX39foeq
JgVtYuCqvZQ6cOoI2DyndwhliRkmH0iNzYoczgt9y5+DujDmfLfe48AgqA8FBCSzDC1zbQJ5j30D
7TyNaq1HZRDALVFcKi078mGcj0DIexJKXGcHvQ5QQJoRofpkYcFnVvmxPLteeQ5r4mBAWBeHzK9k
e5jhoKCU8enQ5HctI998+wQnyqYO7HNCUi6rMQusSseEynZVOUXFBRZt3n4i3Z+jPrDAk8aG2+QL
8GR8mcy7fGU121xzwSqG3sxCil6gxAY3+afYwozOnAbCTM1ECrJFWFAZUglPl0F8tbmRqaOBM0Ya
K6wLsj8+AZvrRI0OkVyTouB9Ti0I2CCvUla6Yt5J+Jl2iE2LNuzlCw7BXQMC9L4ASSAEaTnytkvh
YcoAQxY1xAhsorzXNCMnKBvOeoA7Nk84uPujeUHqV1LiAaeLTLZZowXfa1IGRiWAiPhLNctbQUN+
/tcOgaX7IQIIZV3RqPyFMqrEAV0ltdQB7/GgzJqZdH4leJV9Hib+IqiPa7Mwexf0w7U1dukE8JL0
Lh+Pztue/AzhaJfj1R5HuNrApaCyQuIK3bo00yUc1sg1SypnTQNNRsovNXpRwf9GBQbt92CwH0My
9CJL3vOxHykVfDf7FEU/BPnhiMeAhUg6bwdj9g0P4ZQXeyIO7GeN9yl7gda6uYQw4vsjdRO8t3ZS
rzs+3Kd8pglGcciZ2wEmChScHVUgGfueYbw1kdUbTXJNDNKc1LT2U+BN8ivdbjTPUICGy39NTZS4
H/i0vFn0LukaWuYe2bMS/ZC6b1ZRxiFRJUKzytD96vA6obJkooy6mxdRqVvvndsYiAaFlDJATmyb
3xtHXaBAFubw7unOPrj53WVHQvDU/DLypz6ta/9DVahcRxPyR6OXSQSfW01thoSWjCCp3JJXz/aS
mpEvy5VwgEkyUNI3SG5Vp7z1XfuaLw9ngcPnuCNEP0apMLHDHzMyuJ7flnFFFoen3GuOftj0Eq14
t3+jYBdn0d7KjWSXVrUcCMWFS0PdW7dpkkdNCIOIYFv0Crhkn7vvtOYJIESRf4m+g+B/THx1DvyA
f5bifR2J67dRc7uNPEdn5d1avBFFzikyuZfFhXwAcSp4gepcQiF+F6a9+7bRJ1YaQ44C9Eq9Py8Q
Ywszsuh/CTx3LsD9UQTD1x7I1/vmFBGc/DLzp8Rpy92BSToTxipJ5Q91C3DYrupS5x45QAMGZz1h
4xx26xtk0NSfQvEPIQiN61WboGZoeXth+eTK6W26sVqQZYGv4jiACueP8vFEAnMJrRfZ/hyyp0uJ
EWZdwT9sE+d/QC6L5fP4hUPmDEut1Wu3WG79TIFUd/2pl9MfeOwR1ZqqLsz4mFhISgW9q9eivzOW
VPix0uVhf7QnsD82czxcJ3O4xRaLKvRJVcwAfKh9dQHkdFW6itEz7X+nIk+AZx8zkRJCdbjAm0Hk
Zug0kN/IoOLgH7k9IfzEAXCHcPRLzdkLW2ZV7RBXZrvvhnR6zy+tlHrQihcgey9RCJBNiSfFgQj0
cYtGnzVh2UwIglpD1owNUx2PywmChHTUEHzAVQGYk8pE+435IjJxOAbk6jAOzH4PZScjJcNXvAbz
hAJppx7nruIyeMJoIjT1Qol3R4och+v/I8PzZLxo+vDIcCy8GK5WEDq+PZo5Vxa8kLYLIrX0XrSs
M4tJcpaMB1yUbsqPYAF9rAV1LdLQHen53+rQjtbxmAVobYmgob6myD+7b2MMkpigc9UU30+SDan5
1ts1EPDdNqcTDnIq9QLT/edmXzTbFPB789qoRf5nA4utVSDq+D1ftiKjV8lZh8kX/1c4rLJstULu
VQ5MUvmxV/4pR6WDsEfB+/B/nt24e8uQFvodvmFtedeS9hlm9oi9x65LGuIRIz3ajOdKfqJjIpAq
yYEsbK+ldxO3EjOrZeTNc7nHsr//S4m7XGuy8+IifFjZEFHd/uun7v4BsbFG/ewEW0Vtw9mPM4VE
Tqcu8hd8zsPE8I8zgSACj5OEwudoYNfUf3r1+eBHfY0uk2BIeH6hEbGTjXNeOswJ2SrHbxJ+VPqv
7kArWIQaJAxn5Q558T86oQmnXJPwvOWI/jTPbd/UR+QJWq3XXn4+jwF4ZTatj0U4resY5lXmsXn0
qaDB+5GmFre3gc7AHyVjcen1AHsBCAkClAnm4yHy1b/RA1YCpIpYg7Q045OpKRt5MwuG6jqiRc9B
36JpcGPeGUQ+BCFbImmBpQb6mfUOHdFr/p1u7FmC9aIiR5cEjxq/WJNdr20kMoVgHL2jTfKeVONX
6vKaor+CWSGdcj11TJePzo7frpkBEVF7BQ4rhu/jHlUgZ3tAYQQveqO6/hFhDzRNntb7ukKy0KgI
aNysz3UGs3ZDVG4IMg37wZV0645lCWOFGbgVlAezPPfcuMD4yk6FkzK+LcxsDF2tSbavJMoKHFTQ
l3lrjHbjqg9GlFL4VqNWFWmZKOCsjcT/eCHd1pkeuCK+DwzOYSEGgdAh/Qpy45rettjWAydns5kh
oVTU/Q6IqImNAIhLy80uldYSOOHvT6TCpNY1EqUqIynkTqoEtEi4/s526nAOfmXr3jGR2ghhL5H+
d01mQgqmBPop3+FOHAGcvoaqTy4QC1weNPtM413ikap7ZDSvxUv+AdiUZQ//L5apetVySLzcZcTi
HaYZ2JJxXOYHg8zItm2RhSAfvsQ48YiWHTI3AKuJihwjULiVc3A8L9HX2b1/xwRMESJMmORPTHLu
L1Iwkc4PNROEFSCXa7sM4orsi3b4yTVB+JwBdxOn63fwivxY7HRlpIkq4uM53bY9JSofgR+wlyqq
h+7L6uH1VHbpleQc/WtpEH63tGlGGNkVaXJhdZS3NvfEewyPLf5ycqUjcqm1X00sS0u8N3Ny7bN3
SK/berNSKCKqkpPDQ2DCa3U72Sqi4gMsD8XRcmHWxirZi3bIavbVnIhxV03HNzSRRfIzHLaGdLuh
VX/z5P0zC/cmusYNiuVuMmIt869QtZ6lLboJEaadKV/47xfx02OfJVfs6TvDFe6w5FfGUZRGt/L6
XcGaNX3sYKFK6E47CzLA0VnqZrwcKkTxZvybr3zQz3tbl7FNpoUzy1zMoFTDLPXKmcw6O4FscaAX
gB5aP6tiwMM6rDmLuOIHhAjL0/lWN6MJ+TrWOZc03rlBLBH02Eix0snwU8PVLk/aE24PMWIlkApA
AH8hYn8ig/x0D+BI57nujf2MG7ZrMG9VkoxuJkfx2Cqc7Z0fvaRcbiIlavc8laFdfyJwEhQ2mHF/
PEK9B62q70br4Kd6o3Buqqe+f/G8UeMIb199PPRzuv73t8IO/0zGjRZk2AgttjQqENz4rY9ZicJB
Oj9YU1DsR3PqQB1xjFclzLuRlMk4iBFxC3ke/6I3TdDFdBWuK1WmxSiUXhmb8Mpcym9sBKqxB4kp
QkBtsNgYFbsGRgMReJCGBarUTQGxGNZjkGWkKdOLaLcCsHiuDIe7yaartful+w1ReYZs3knnveMF
xmR5X35/pOFYggO0vcDI/lXNOTFqvvJgoaQtFbz0ARPSOavnQvwLfbOOnA/dZ1ngjHqMK9Vl/8Hm
VTzlJa6laVHjBoC/brcoMmdCZkdfd1YQRDh/sfP8yt8+WxKMMrSRcpvoDCFs5rTYwqNSzHmkxixH
gSUZIpzKe9BmK9GOWH3hWLAjtzXgZhHJwImP92LvrR1V2kPzw2Tq90GWfvfzxzvo4CmmpfzJRxbJ
Hp3xUgGOQd1JRsYOMF98f91QmRGX5xSh472WUpUsnI2r2bdZ6AtvACtMl/jOd4UxCtzX8BpAKg0G
w4yiSBrfE3OSm4E1Xy82ZiG/JhkJP7522PT//e3JCjqmSctRF4ho9V9iGk8C9aMptooVhSw0ERzK
a1PoecqMV9knvaBnP4+oJ4GBHeWbWDy1UvVWRLkBfcVRxsdKbFaSW/RyciR/bTG5SbpBwNMOcP2C
wpSeDSe+H0H5BJYsuyHdtc9BGL+1szhViTlw5GZ5sE3UyeRoDjQWf0TSQbQW7B12hT54JFc9I8qH
DtUN2wT9ggB2htvJc+pzBkt6aNaacGFtQ8YL1g0hubSi0t27E3im+YcvPgXIDYVH15VsEsUe+94e
w2Vubyy/G+d4cwVjwyC2jgRU7MiSvIZoCkP3VKNxVtqnuSxkgFEgP/eqnvzuxUO6BXKjegqVoyIS
cQV3gOwNdn6h/wTNyXKGsaQE3+UxDHhBcSkbl8Z98slnoWnVQb1CcvUeKCRUqcKMvaWm/7iLP6GX
x/zl/FZOL3z/mJlUNvu1XXkprdtY9BeR41yMFnpTx7NU4CgovRYjfZVFJK1bDGv0YXGj2Q71DtWC
F+LypCBV1bXqcJYBotIjj/tfF8eeVv4UWfR4JhNjlglABNuLwF2XIb1v0LuggRzME+zeKYIyfgTU
Dw2xYqyBy106XSf18vZCdRs9qQW5uhqC7d28qZg7BYVlTTokpFb9qhiIFhL47ZmTFnXqYWkIenc3
mWWxb3JIb+Ktt/NrpkYCIJSHeBdBMaBj/3DZHvmLffHvrZr41Eent0VE574Zszykul8a6BwsJNqk
TPcgLjLvQXwX/JlSHpsW9dd9O3jq53X/kOa8omP7ILxxiYaFzpJX7T+xU7QHa98s0Sch38JnfCDl
xQhYgLC73HsurLH23ucewUj/EHWQ9klEJGLlU24QsGb23nKm+p0IFHUX+hSAx8xgLE9vpZ6zZtP7
Hkl84kyUpU+FOju+K9rNdm8PGyBa+6UdQUO8N85VaEvR2a0uxQgpx77Dhy/d/TplIZVSAyIEoKj7
nUroh0lYdsmg6f3PVz8LNSlWsMAM4kO/lBaYmg55poORVZpdREo6xGUtP4equbjp+bAyUDm3SSGB
a1GGgh7+gLbVRmIfSBTRIJidHTWqviplTVqK44a4PcBm1FNvVztvnB8kifV6bG9ZUmYTC6OGLwfo
5oZ4c8ATuM3FCwJFIaA8UK5uRDMLJjbMtzG32r0hRZ+ejnbiQqNC8kEOgBAYi7zxPsSM3OvkEH0E
8iBTdrwG6z7PAacllhzEmHvabqgQWbfvZAAq2d7m2aNGuAeqQf1qfyewGcyriYVxaM7WgIR1aeB1
y6Qlpk3/9CmRL8LW9ylmvBsidP7KkmNBe4vqgn3xrUR8NoWMrdH+BXr952ssgbl7uJDpU/NQ+i7s
FAkGDA7yiYphpzHusZobuKz8YrGTpiR1hNwl77QVfjKWmBrOyn2i1q1K8O4WoTP7NZGlk0ezbSQ1
OTovmACoSU3VvmSQ876qqYjqO27HT/Sjh8M9b5TmtmHZZiYuG2720uhVtUFkP06sUTXs9bm5Q+GI
BTKPEqt937fpZpOEoX37o88LwmwZ/NN4/67Rqqla1HDFUujEerREXq8RFs41Acr6+AdFU3CivaSl
QY3FVw8shfZEzlm6WU0kh/ekBBUHP89V5qiRZ5SiHqxsScug7zQHmwWtqAVD10H804e66900g7CD
6AW/029CPPgKjDif3NIFicRZR87qDhZFCkdUNbzFDd89KMgJn1sgiGp3Gr2YldhixlygXXNT31nS
+m8zc2LatuwhEZcDYWztOW12R5nOGGTz+fw0rZGNbLNcL1aWPOlO0CAE9k1McGgT/GAIkJ5ngZJc
xeBUy0uHp0uckCRnadqcksXa8AvB6Tc/gGttZe52lx8H0rRzLGxB7ieAhbbWY2/XwXOzU4srtDGg
2tDHhd6Ylh4wHHm9yqEJZ1tfbmWl2sRowdnFtndSoPfnSxgskNBlZJqyl0Q/Wgx2qhSmD09vP8d7
gjNer7/i6NA6VjOUpKa37fxpFAzMDmi1Hy1rpfSbPrDVD1p4eJS27XIWC/mCRCh3xX6M5jjYbiH0
WNt0AWQb7rP7O3UJupW14qq9P7Y+ae4Va2EhruhfyY0gmTB2RKiAlf56zj3LF9u+s98B7rvMsDe6
XghcypaWyOfLSOe40srj+TiaAQGHwM6/F6qcaAyot/34XY0+KSfYE5X7vTyDgi9RCY400oCWZCMd
rbMYCsJkGIv3/APs5geJqAnaCVK3CuN2+QzhOADIvGKDXkKRSJ+nAjxN01ybdEHImwRGsdQxp2RD
R0uuFsG4wa/6Jj1/Nqci6RghfcLATTnFYMRjSUfwfkj++kH4SCvpdmiRP07/PfjE2OdYDEMB1+ni
Zc7col/utAf5Yv/bMxyeVSBNKNC7wSUYPqGrLhN/Hlfz4XpGX3KRX7UliUjBSVK2HdEcqlohVgGh
YV4Ru4xPQbx4XdA2jfU2nTJcKiDlHdhx9RwH73F/tawX3meKG8a1wLy53U7Jsa84GhcMODd8GDOb
lymZSyweim3Y4id9Vk7LDxfduVNYenP/+H6geXREQ5jdcJc/n3yKUJkKeSwLnIStyY93A8Au2GcU
ZEA9F9oAqzYyLnO174ZBF3xcAO65RkTmXjEs2GMWhaeSv7FRwoIRRvENJ/W8Bq0l4QuuT/xwhtR9
6ZPKTt6OC+D/fX+I9JYn7NlTEMvjZ4s0xPvX/sIV+KgFnjSqFyle8AKASOq+kNKBjKjiBNeV7mxJ
WtUX9P1/B0tx6rHTmBMwlDIOowG5FFGqQPdr0vgdKdriZFFzB/6Q2JoTdKsbFGES63OdXclOLXNR
rDnYHz+gfIgtcgEUMesDeG24ji/mX65nu9moI2K8c4wZ9b2r0awPQu71zeCRQPUj2veCHw9QJkVG
1PGdx2vwuJIyMdGsM6NQU6pXuU7ylxnzYvK43rkUDLE4gFWfz79JybTGSKc/Xt9luOHwXoBvSOi2
xEKi3vGxoNaKd7b8Sxg5MyLAO4EPgBmahuCZm4QFT76FY98mZElb/rHTDMYKavr3fQ+qGA9jxNcS
7eYRDv/RTlESdqjaoHY/J4F1sdlqGkIT4X7X2pWxT5SUOU2NTYp8R7x6sCAFQ25LwCz0GiuUikfj
lZhqUzZ9fYfjaRY25gP2ZrjDsLB1FwUqRbepWdvgNi+keKRXlYnvyZlF6eYWTf277VZFZX+QFtHS
urGGgSFf/sCN4wICKp/OrfKddgwD4jxhOkAiZSJPeTet3EjMypbDgBtcDlvWFMRpyr+tvQJrCACK
BHLfbrHwzFvHXyZ4zJaoW4W10Y5tznOEMtWhqVTRBjgIxAyLq2si8UQ3CRhEnh3GlthEva7iVmSs
Rnl+3sEwytSX11b3XR1AG1l1wAdQ5n19PphsDkacYNdh+gt2WCf1Q2U8rge4mfZ2AtgxrlicW5np
iu+3l4EftDNryG0C4q8WgSM+8mP1imdAPN8p3kaAtD1ynoBF8/lUnItRm1QfGTgcH5s0IdR3iBy5
NJlAQWTV+c5W6vJFOHgX7AWx9I2oRlB+gXQNugGH2Pfm/NCmxKUJWM2ExnN7Nn9T9varYNrBUeUi
2MU3g6ugwEpPen2OlIjR4cldOh4/Y/gTqEKKCbLHgyPzOAbInUg7pnzEvrHUceDRlp+pwZNJAYDp
UpWau0rTsAGEt373GIHi+c/C2hG8LhNJmg9xoF68G23+IbvdXbk8ZxDd1cwQIjh7oGbg/WJ6BGwJ
1LYVWMY39rYvvFqjrvEUfHjcEeLrWdOVP/ghsAjZcZkpsfk4hDHX9tNJIMBkqcfvEeynVKXuPUQt
6tr+xZjuCFRrB9PZBPok6Kvjh8Cwghx6iFtMsy33SDltkml0okqETTs9zE8Y8ev5S7W6293v0iup
sDhIczoR4RSYeQuAt7ZnRYinJZGMK4+uIG+OM+l2dypo+Z/PcMBS64PGq+AVinqqPYueWZ3IAT4w
kMdrlau2qSU7iDNsAawSa1JZ7QTXTBj94frjJSSDJerGf3ugsb6WasHnnHwkcrmlpTvowEmX0FeW
FTyLCcwbiNeEsSlxlbFsNxz0XE2P1HvnwfMTr+HKDBP8HK3FgHXGPA5UXFPmY6pqGMdQGiEXHuUc
XnpKcHUL/IdMssPH6CA+2FrZHsvdb5PXNbaxyfhMVhSXqz9XRt7vd/+XDQctDbWre8jfNcX00HXL
P5KvtgTOETibHF2xveEeWRP5nXYfKJjtneXk0uqC0wKxTdLbXYA5/2YSK69kwJOhCT+P5hbzHu8/
RPT1Rinp2ZmFCGwNxnWLOaozelw0K/rlZv3q+IzMnr5Mj8LJ9ZK/o4peeoxkaJ4vn7zLzNfXLQDQ
fUFPduJXJEnIoiZfRR4tqB15Qo+sWyoRv0A9cC0x05vmtTE8alR2fsZcwaRyUCMvHZnD990i/uNl
6Ud1c+aZdFo38BK8cxxQ882Hu7bsBpwY8Xqe0REP1s2wPOsK7D5Jw/63JnTFOcaW85qNVgT5aece
mY4Upx/uLJmozvmg4JQ58pcgXRrPgBWprOXBTDNMQfPFi0QuQ4lS69Mlbth92m+MPYOsLNjNSMjN
luI7IaPKQIIpKeZvpZ4PneV5vFMG4uEjyYIJX6mX4CmqeSkYSt8f8WqkBUabXbotr7q4y464gjuk
6Y+ZF6jKTictPkLjHNvXlEr1A8jSfR0WcIESwxX2vlDF7qfNHLBPpSnFFSwPuy0i34p3WdiMxyPH
37LuHA+QhnxZF+yN+FI9ycdD7q5jcN3XCRWD9hk+4E8JZaD9XQA/NlIPurtDn4tiz1yu7JPZ7v2y
nGAmUzTRY350RvUDFZe5TQIBM25u3L4hTtn2ziBCF9thhc5kjRBh1zxnb8hFEpvh82Ms61JRww8/
nr7aDbIlGCNPXcLzdpRqNG7S7Aw3EgloPzk2julXQ3N0E92+opxwBvrWDRHIXNjg0M7Yny2+T6os
Wi7oy929wTCiH6j2pKBiPNTW2HRQ8k3FXI5I1ShGZKXJ73ddz2K+tukMyzyYN4lTCUkEq+C5FVoK
vH1++dXdb6FdmSnMyvpPS5CvDkUTNfqS/8w4887ybU3UZW+xJCqcAi7Q3vmY1vjuE8aLD/KVGimM
eHh9RvDL4fCJ9RMSv5wL6uaXIUAkfuY+n5v0SXdxS/o/IEYb4Hn0wa5U1Dujn+3KrQSJpI661SpA
KJdLvWTzIiRIBXEdNXs1h+dax40Z4AQWBySc2DiEFpzNRzrBqp3iasJA/go/eiAGmVAzSn2KAqVj
8riZ5SJNmZ3WQ8agoCBaMNmO8b4pW9N9xm3JEVdrr+IB/Goe1JdnRUM1K/Mwot7ix31r1rGKQw51
BH+XS4tpRXPLlxoGQRxRrS0FBLJ6YwD50xyCjXKne4B/XsTm6KHIc+DPyQjXJOAdPoTH/B8eP0eu
n5N3InSNqXMJerk8DzJOxtZeszl9wcrFkHRPusMO0X8boWfhLT0tv4xCnsRYZK42likh/mz6m1Hv
CaYe2EiH+qTeOHo8MObHo0Lt2KRJotkA399Jrhie2y4bmTV/WrjPj44ruMeW3rB1wEvj4UrTVwrc
VH6GBFNnmF7wKzJdNn0WDS61IQRbFmRl2rePRt/S1X6BdtuXL4hwb50reeTMUVWiEjHQMbtUEMXm
7RTwpCSfY3tPBDcHOkoWN/gsPStMG/dBi8XrILcT7+YMq4JYNLDJGLB/h9TXEPuLxrmyV9QG0zEr
f51RDLG93LalTxwcXUWjYIeziweWq7mnPZQyvt4OdMLqqv/LTB9vtzcfQ9YNw1HfF5rDkZgPjeKc
WMdeB5B7vmYwKfCAoKF9tcVXDZ2O0PSadGMA0uZu5EJUnG6KZeA34B6nQcL/sVsF3mgVZEJ5M/0M
B8Fhd5cBgvC2Kf4IgL0Gla50ZQme7CfvwLAmJLfFlCzKtPfvE+Q2TYrpk2ijSS+4RJhaYzQXpU3c
bsABomSF5yaMo/rJmkiFvyVNbgr5G3IX19EseYdfNJAy5LZHY+m5YyLWobO8p/tDMrHqRas8W14+
xwD/9ueK2xXWc/F7dYQZV3rk1gAEL8OqPry5yMArTuFrJie7cHiYOScwESbAfuS0ld6jC4hIElUf
ZyT/OOnwqTxejRQoeluKiqcTw6hmXlcQuyEyHumm+HAx9Icj3zca+YKDv2JcE0uh4+HUlCHw6b0z
h7PYcHWuDYKOxx+XkSfs3KDf2Pbg9dHLBo6BcukmIKwlG8rXtK0853o0JylbG4O/vrY1S03FUBB3
d53xbbMdAciQS/SZOHpV+nnP9mJNlbq/OjaplA+LowRJ3GeJXeJs7IE759ctLn8e2VePaOb0lqqg
NiZOC1+efbDJwVum81ikq3Fn6K8fJkqMX5w6WeCI1Ru1rtcRbDvJUyogXwWuToBIJPwgAFf/1pvc
Mpu+SVYE/h44jvJxoJL3XsFqbViB7eCn6k8l4O9HToNr7g9Ju0AsoqlmSLReJCEorDUuAyxdIwMc
x9srY+isnJ31bk6Q5pKHgRYvpmMLRDrbJNzZjVxpvDHNbQ0AmtbUnw1pwZuWpKv5/w2nj+I9MwE0
X2B/Ha73MEWRNUKZJqeV6rmhpX7cAFn/EPYmkPI/DH2hxMF+AYhCjjWqLazXnCZxPxQsjb+qJtwV
nfNtq96xHzNZq74qdBvJWKqn7CdWym1UjcNy3x2rQyu81c0FcVFnows7vOjDIAcQyMbpI7llMYRI
4fhHIgpqPjv/c3llYMKz8Yw022UUBlJu0GsH1J/23DHH75j6Nxd3MHPXIV9CGPnu2DSNZELg/M/b
essM7iUw8O9ejX2bmvMvcaV7pBVYbluF6vNm4tcbd49iz03kczOctnrrjpLiNuMdjB2ar34CS2st
wVc7t08jebslmKBFr6uNESD9Rum8CB0oPIJGTJmUaKarOLzwZfNqn15vkoRoeg9n8rDEQyCgIeXy
hrw7rXIrrlUXdHgLy2M1bsv33s+/w0H6J2sV6vkG95VBkFVw8uUEUvVaJXA1rsa1vcfgOMV8FmjM
ALzZwgLqwN3xApHBsdoVyfZ4kSw7oLVys33nBCmXaSxo1pkLksgpooD9uuaYVEY8kEy+ckSpyPkw
1zs3D/wDeNiQ1lnaxzwBt9ayIdm18YyadF/tCbmXxSJn7U+ueDZ+OW9+tOM9KLlFK3bgfQmHLv91
kycSaiWuZpQ2pVe4Qi472w3ca9duLty3CtxlqBujxAwfgVOSCrf1yDCyKHp7Sqqj/wHyz+F1YO2y
TTvGIqDqb8jha1juYBpznQ4aWQeuwk0g420q1KtvgiN40QWTmcTix74N1wgzQ72fLWauUIWfQxNx
Vvyufb7/r2/VbkmHRtWaiKwvjQEd6zkTtOvCCko2vwgC48LHIKuntE2iHWvNXjKsarv7lgRQJUS8
IyvaIhLGJJIIkQGkI539LqyDSOuV7MslDr6jYPW8FV0bZbOJadz0bsTRBG0kddq75YBqnil1TtyC
kxiAYmohpyHpz/z4Qrw9sHMxszvwow1lMd6kQ/xzfnVopMyxNlCNhICvmGNx6Gg4ZbB0V5cBJqFo
nCjnvfnnSA99PydnrWe8SC5e2nBdno87as3imsNKUxy09VdkChw5XVFywA4Emc0Y2i5YwhVZ6RyG
rwC/cBXTfT2q9DJEz2nP4YqzcmIhDihPvSpOrZWkKN1e77frgJvDr50Qg5oI3zTk+hEIx5B2YlFf
maVl0qbxVnUPg34h1h23bzkYRHAlaxHJ7UkFL8kv9x3OZ/Ty2SeS5oEGjdkeyalJbBscER7hoQLW
KpJ9XjX8MmpSJw8FX6EFCFGHAUulPw2cHc/eFNky+xh1HsIqGx8fbWQeTN4lzCKWNRPjGJw7AM1B
toTRRMkcGKWuO6LUTTPZBzlYgBA72ffkMrkPO3k0A4e5pOt9MxvAN/VoKjTeUJD4esteJTa3x1Td
5ss5/Qv/RjJqNiszBQHxQpDl6xpkJn0XYK+6axtbED4zKjcQVuCxF+0mVTbFf4RnbNPm9Q06rMD/
66hD5Vmqzz/hAwVLqu3dWpJ/XmdzuYLbhjw9YeRCS9w+2pvMtJ3D8y3lddjc8aTjB8H9D5FeQUda
U96hIuQm6puxZeJ06wn4CzdJj7toCV3VUfcy/EZQa3+87Gl83LX9f7px5zITFuHI4XOJ8KZBU8sH
4UP9eGGZrdd/lGdC7dlexkIcfJacCsGTJ6Dcou0ZzfFAbuk7g7lVKGe0+zd7vckOYR2NVa3pn2JK
01MVJxYgoaiKMSipIB4JCBGKMZ3QyROjn+409ZX4CYg5WeIHFu+4T4netTv0ncM+fSLokfc1KqOb
HHFxVo1tTomwA2z4N/+S3mknhinGDSjDqDTQn9+s81syfvxkzhsZ8XBC/42ePSwYifF3qmaqKZih
z28AxiXs/HDOIA69cYfcy5GC0wze2QCmo0pFfiXtVLZre1NaolBUZh7qT0T0lv93n7OIjfRxUm9n
IiPfrMAP/Lr00ylTLDWdHYL/9Qco9v87331q6slUHvRY7GhNH5Bkwq/KFUd7R79maiMrpBaAbjJP
WQDakdXkGgzSHKssYIm4wZcA2rPHejL09sV5Ztfog4aYuG4bwP7VJ3IoH9Abox0U0Gxbr27wwqE9
Sj9pTL7ffwzHBPWTwqi/fEIH2c/eTbhF9XZBbY1rW1iBXh8pDXbtgNiSO5nQLzo/t9OJHfmuupvJ
Q+D11gS/CEJ3mKjr0NZvQFru62s/H5JfBuWHIweL4KfR3z3fBLlqclF6DmNX2GBfmmBgNSEADM6c
UscDujJIuuh+cv7eqbCsETGAKOKzKiCuxFqjA/YmkvQ6SDWp7uX2QwRwbiMcrm30u7vrGWZJvnjp
8nPkXXutVMimeeo3UNMyzNEM2Vs//tE/O928fjSVsVDZ+X4TcHawexfXLzMq6EaXLEau4RijI3sJ
g1Vh53O1oFkZncEaLPtSb4Bc4mRe2xnYZu6IrfT0JixvU9Ev/njn5bRMcG/q2O29ocd/JYkD+txi
jtKvv5lEWIt4WjVcOduHYX+gJsyOAAwbDn8Ubprzj5OTZEg9SIMjyvFXvyS4if6A4GZNWEMIJoz+
qPayZmagrD7gAYf75SyPBzCFL+JDtmUVrBl89Hog88fXpTbw4Ft3zjpbIp2hc4EZAXEadj1YsH8s
NQ2L1A4sq3b7vorotri79pcbkaWg6xXaabdnuyHNVQSYuiffEDHUhdSBCaK1fpzYpHz1TNPkdi+j
1MgnVYgkAZUaBGfLXFRtoE/5i3FdvvjggrHn+EzTgxteT6m6aMQK9HZIG3gzT/bK9XGoph2J73of
k1f4lofdG0SoeG9YXWRqBWLxygLaw72+ZyB3/sONMcY8pYguE76Z7ge4vfqMctpEG1ddjgDk1/4i
d80QNwiWPyzQo1jyWTn/Ius1vFQ3gy+520B6fFACo8mHrgao/DQMvIQw2ibNp3xTJH4ErLanZyCO
25sW4cfRoRiKI6Cwu4tE1nMXCN4mHqr1LT2xf38ffcnDiFh/RLCAijtDh7OcAMXIjCl4+1XT3twh
EyWvE9ulQj8eKrEp8iK4spODPKawTsW+OQNG0Os0cVMh7gQQxAjdEVJfyPJFYroC6ncPZ2KIVmYV
AaiYdUhVEU7SzNCiBoRudacB9f8sfzO1pgdj8FRN3K9CKxD5eG6+It19ceAk5RXLsiT58p+QrxGD
Zz8CR3Hmr6NBdYV6chO5wMaTg5mfm4I+0Vjv74yCFdHej/L6aninq990gDJmH1LKFxWuI/tvOKLc
kC0YxL4QEuVDAHf4lAOJV+UqaFBlap1mfGKT4LMx4/5EFUdwoZ8JL77kpcdb4C2La8BWFH251Nt8
XXhIEKj0WqO0nGobzFXhcHlJ3+o9BW9t7V9wPU7yfVyi6LUq//bU3QiViAsZxMeyTHDZkzg5Bkxw
76cTXaNLo7sLYiCggzila1YW5F3mOiEZH182qK01YiQ7sB3JFlixifgvzi2WEhNj11VNDHGJxd/b
a1R429e/Igqd/EcD8n4mB9JRRkFVUbfQeaSa3KtyZDoP9d3LqSLzK7fhWBUljRRpQi9VxXNRn0XD
6fsv7MvPIrjMo/zZ12ImyEY0+ZFvUXRa6ZqoPtpjTmu41A9w0IWSLvsldQid6Btk6PMbrxzmsZQw
c7Cebt1o/vYGwCgqK+ivFUVEjEPuMX0FVWIqrX1Q2sqP1mZTiMSKvU+mUbwDgakwNE6Zo5uvxIRT
IqvvSvc/NZlgwanaRj/gTCMYkRRGAyt0SLWHfym7WF6rHUNZHtNxfhmHGpLb7jLOUht+iw9YQwq6
IeJih3CzRZLEdyavRpNm6Lz2eL1GkbC/iWVUJWWDMEdmZo8n9UM1IdFSPupV7P5zPuDNpND2gG9G
4EWsZOg+QUwCB5geYTp7RDbOQcRmqkkFR9Un8LIqeKjPKvB1W2+Oy5ZScHVcU4X+UtBYL7a0mGRX
CgQiI0ZE2SNV/x1JYDndZJ5oqZ+8AVQmFvj5NCWmseuToF2bDtFIJ+ZYtR2LEVMdkXeGTp1azEBM
5FOw6H4Y9AbaoicXMg0vlOKuIR0ZwAjunq8WTp3vEJC0/dDDTpQOI0y8T0klby+jz5o1VIH1FwgG
FKXaawkW53udn3QJK5khgOu1ge0voGEqD2fAydBEDY1cGu+GFS9OmWd41/gJvSZ9wDE2o3Mj1M4k
uhGfYqs3QBhBmTKLhY62mesQ+s8GlnJ6XYDm4hXrDge//vWWjCLxPZa4bZSjCQaQfwlBGU//cEQt
VOZnaLavYqDzz+cZutPmoFbRLoQJSF5yyZBntUQQCHcMXEUpug7CiJrtOuWs5cx3jcYnglsYm+kC
ce7ScoXxZMfcHxlcU91b6CBAQVm32tnekZz8xiDoxhVp3S3U9Tt80fpx0LNwViDFDSKKy6VSZ0+Z
qNWmSHZfmO/aBDQtRR+UO8Fk1CodjxMKr9HSdLq4R/YzV4Xix5/yH5tVZ/o0D2DcBx+QLhGJgVJI
lXWef91Xor+lwTXJ5lzt2gO4ZCiYbp7Fv0z9WsxwMelahiQyzLdP96+GA++IO6kqNEffe2khJhCy
gaIBPDZPazohVSYQuit5EGtudnn82CTJ+5hxtHJZoz4/qvefa+8ofVZgOtHOGkz7uzVTto83ZbIY
rm+4pU6X/+KQHERTDhP+7kpHDfjYiuvpEoLDljXA/SSOmPnvs0LgUck5rSdYZcY0jkR3FFuUEbXF
caFasYbK+811sNHNTUfIWrfju0irZNf3R5lFC7U32EBUeL8L6klSUUg3JvhFjsr0P2MjTNHfrEWJ
xXH4zVos8j3MJPmBoRjWOZWa2IbtNSkOj7oDzysmexhPHxOmEUGBVzN4fm2QKxanz8DaSaj2Wces
datZKGMqHRuXuzmA7H+dNvEuSuFwG7a16b90yUG4HFJiAUNOWz8iZHEfkcR1QIFpgNN32gVlZkFs
J0a+t/aS4YLBMgkOe4vVzMRuPC6QaalOVv/rtorBAUmNjjIVmpFf/QQrvf04A6/BRNqdBxA6xloD
K7V2JN++bb4oiLl30CoOzmt5AYcXDKUmJ1M+eA/uVGM0ZZ7OALqIwhnwniWuKl4jvrnevurUJCLV
JVOhwEL1XVftKSrEDxMxIUUu6RmEUorKeXEBfIaehyt3WyWfvbJcM2yXMKbzQ6k7K4ifJ1Thq3Fk
r23EM1cYNVTz4H5M0+cXGKxLlPe4ngrarPIINH8ZTFy0g9wzcejzsIoeUWXX83MsTIyeZP255CxT
M5bRdNwMRmXTsML6yRZoe9BTraPpTrrA7jjw5IVIJledZbvuPxROlsQNk/GFflRlEAe/Xl2mPMfB
mW9hvcHI0gq8nVtR5+EtnA5FRr0cLoVjkmkZz6pF0QNeSwr/XPmR3CH6pi8eFPp1azgy80gBqzt1
UoBNulf767MVtE8clh4+EeprYo2qg7cZ6uRIMvhuf29rF9Agusq9sBnAVVfP8XWvlxFhdfHVIGM3
Otvw0vC9QgySEkOMd9jwOzsvSVBFfemtI4IJJh4VgdL86dW8F1ieOxa67qI5Q+W9tg3p51BbWzt7
6k2PZ/fKzFCAO0U5eYca+eCfVDxeGiAzeO6lr7Gp8ZzMyvcD8XgW1aoEFuXqP31q4GWbCLUmJyXE
M3f4OptbqePkhrDcliHtNnX+t5ZnX5xKDbZ1+RfPXHvawV/XF1hVAXtvWiJO1DmWiSNRoUXepLus
Dti3ilPipf/0MV3XqcBZU6Hm/SckaGx4NBmerhko+WQxze63DZzxfviHzCsoeFNeq9K9iEaSA+Ha
Fcrc/8anvJ4wN0blQgBdt2NZwnZulx2a9fHcOqzA653EQJZMXx79L/Uuji4Wf+n+UWTtarZGB83C
RAZinUy75t1nwx5S/1VsbP4xVNM4sSCxITRh6UCWEy2a/W2sUX6xnQ/tOE6IpXJvVRIjJTQErN+Z
0P5S5B7IXe3/w6qZ4ac8wBRt4JK/qOePu8TIhoHbMARNCS5+UKVLmSGX7oYwN3VkHOYLF9rYLcoy
wEQBlMUDXu63qiRQRuGA4PLNu5P9A/PJZ+9xkSPEfkG2T4DEsS58zPFdyKc2XRMR8q8bfXY5Np1a
eImXlKWP35RYaw3mdo/4ksoe6V/stUsfrGqegEofUUHQ0WqNApUcY1Ah+kvmgyUspOFz26OCK6T9
3kbzAUN0Wd+C1xzJCyjiaM5o+PtkqOAti3L2z32ul0qLl+/V2bcf0ortyTA964RBG/jcfVC2PN52
O/CWsDrIAQ9LPassOhhA5+aVIInOHeW+0WzZyAhn1J2bAFXlM4J3ivb5ALOafiUprlegBsUvbZKs
ytXLKTYf5zQVsEz4FKz0Lbpy/3/ZBFuc3RfiQGThNF0TLXrxNaw0wzTXlNmwQKXWnN7/bssHBoI5
Mi1vK2Mthwhh7sBqg8l9GvKbMMOkaWpS4L65uOF+UTLwI8eOiE7qMIrvuObsp9ROiWPu6gJ0sA+k
RNrrmcCuvOaHrjcuUqXOBfB01LfS+yPk8KaJpjnGbjPA9CnjO3vg3fhKaNBnHfUIXTkdr5WJCrpg
p/eh6kbWQsuemurPe3D4fXwTumhdRGzYd5Krpj/N13ow8MmDCn+cnA9Q5Yn0oatKxNZz6/2/TYF8
lbkVT99oha8XRLlrVCGykZVupJ50Tm6Zygq2gmCpXXTATy2RkYy9Poe2XWkdYjB94l4SMXYOgq4W
+mSc4gkw/MmHFSUtTB4j0ZMbZ/ppK/mi9TnC+gT3KmlaCaJ4afx9Pnw5Yk3L995xr6swzmf4yviu
QMFx2Z1GxNMhm3Ly4UiXhrvpGuM8h/6ndhEZwbZE8zQywRMC9E5gXWNzSnze9hvJqjP8gs1uo2r6
0hvE+5pY55OA1NExDAWsCtG8Dn6EDBFuWCQJFdVwkc+Veh/z5pIuK+dy5JEbOAuZydDnLF0OqObS
11TD+xpMBHDWqwvA3D84sBa8wIO9sxzIxy6dKFEdlPIvT/EmuBdfSApnh+vBWyKYCMpmNrKUS0DI
4eTrkYSspQwKWRh2AGS6OEvhmdH3Ois513z8MYwGv5kKDoneVnsfeRATGPETQcw07sijD3lBe921
76tITp05wYnPn2SoqP5u7veoCFYGMoYwYHipv50O4/gPuJGrpnOrHLw36AEQAVNp60Er+TUuEx9c
Mh8m4WCKb07JOdvwsUOmxw0sJH+By82F6bKReqIfEulU8VFhywfB9Fc9/0bfu8WXhfY/eKHagccy
75TR280luzMq7lwhF1t+caejOlIrW+MS0Vck4rytCYQe974Wgr3fUVZ7fVtuOf4QZHGMTnm/IcYn
60mcGhLQoW5+qQoKX0uGqVWQp+pV2KPkkI/13ZNJBb0Pw/BOqC/asafQI8JHAHqp3Unm11D8apZA
iQRLLDSl2t8eNvIMpZKOIZq48cNWeM1jyTOLuD/utF6mqpWA3HJH75XRTDq24Gzdr7IkKJWVgznN
0IDpb2r1WbwycxwhzP0NhuE/rJpokDLwgimRWDgMFL2EbIcaxT+LKOsLmwEKiWBeRgf0wb4GxIp/
GFTo1e3vesvYMj8SdH9A9ZqUEt0v+2sWPpapfAgXxmdQwrgzxd4EVSuSsbmW0ZWhyEPssgdiNxkC
H2+0mW2KPnhRECjlYL0DUMhU07UPZrSARdDhnfsfZ2MaLqjtSYISu8oDdE4OgdQk4LNNZ4W+caWY
g2K9VMV9x0/JhsnIEpFUEFiL9r1jplhEsh4u6gk651XvjwFa8GH1LXnBVN3iyq1dSodcGqSpXt3X
VRkELz9mfv3GDY6TMTM/hdGvgAAFe1iAIraOvRg51Kyu/qBvFP2nN1YFEK6Y8qLHdRF49r1sQz8o
xLASTblq0PxI53wNInukYE8YzfYePqxiay3+R/VYaMjLHZxQFO6nRoD708SgZcgWFljusfo9tgx+
5mNQrMoKe5RQCsQvAlXfnjjK58FyUeVDZMZbdAbOtBlUmcUITczSikq743NJs/JEZP6PkcTW8cRH
sz8W6ZtJ/+rgrYrptd3QW+UVqzixyvC3JqrmvJI9IDG4zGyJSy+TTuHFBjjDzK2+2EwGQyaDTzOs
liWhYBrcBdEzXfrZKHXkNae+P6a1ougmS4ZI2iL1ILX43odpP2mABLHCMCFZyuMr7DRAjFmsrp/Y
MgZ/i6sQVXoWRECE3mg8sXmGRabGBKb11g8UNFgkThrKkyRXsYDogn+/mn/VRWS84281hG2RLgZ2
YLMJyv80zOaX1sKCvJfgLSjW7wHTorQpEweDUM0SF9Y74lpjQOm92Eiai/dIGKImAbY17lZw3KD/
Pu2VNUZg7NIV13iCMrJy1He7fC3WxhmyTPPtQFde1PjIPgQlDwTQ0Xp/SQDGYxkwgWvezMhtD6lW
WuqNL4cOFuocb5bkzCqQ2r2nNh/xcNaJoJim9aUQaSoXgpzxdwLV95Q0HD+kmifnsAZjEKOgYDY0
+SdQodBxFh/3hD8S2E8zUzr1FUouJUkO2VOphzjaL5Jo/+IUl+Lt8dFX0piTPmSnozCiqjEv802u
Z/TQ6piPpsBn/2V//rtv5I6Co/MzStMaHlxdZmBkUPO45B8xVR7XzNK34qXClHYq/RMwe2RmrZCD
srtN2Fr+nLyIE2dPEUAKzv/yYv/4+lXFSbYYeziWZL5c3ozI7ZAcY1XrvQYwbDewTp0Z6sqATT10
/HIEHgPDiYksWoFMGW92GNKP9jVMFDNtGRcF7dTzOFPVofyGaxkBrykr/XeM+tbDFoC7HLWYRRlu
KxyuO33ySKasvcYqnmAgMcU9Pudeob3IVY6/sG3OJlGo07otD4e290RCfRUHTQntuOpdDYjRJ4Gh
lUyU9UXaoxb6JsqLIjPFoq2Sj/WNJqI1olLklxtvdZ3drrMyptJJ6OSvhb/JnBX6qslMFGrR3tQO
jtgYfW2LG4KjJ6HxvGMOxwRsjfsOSZxGXxW/aMiIvhSt0kusnb4vVnQpVqxIPsa1v8e8W9bMOlEL
mpuD9a+k+OuSChav+Mpe8X/C6cMef/0r0XqStaqYDwYGf0gkwp8nRX479ffu3fRO7I4zvFG3gb0H
pMf3eUw6UiTkBctEL8hcvWZTJdVBhivGiUjq8jKA0QcyTB9Iks4nYkAmKyv04Uok16fjz8nwHk7A
tGXAXNxDf6BG/p8XU8Dl1q2qburdWezfVUH6I3TVbsAquQ3Eaar4XKUrGA+MHdFB3GaPFRP/NfBw
Me/YqzLSvQuFMAuOQO2CWR16FpCbR5htNmgGRpZptXp6uj2Tt04cqZ4mpFp7/C+tuxRY2VuGgy1c
LcNBnFqqqnk+EgM6cOCtxvUct6K1dlHQ4iBlWlSd1PnKOfJ3XhlG/bu9/jGgGyih054E5XA9d3JT
mzN4A3B1qEHNtZUJDSasHj4oL1DUko4Ga55UPuWQddMcBQS8Sl8jCf+CFq3oX/+N7Ic41KAXPfTf
vMD/jmEf5Eua21azv0BfNdKErZqdKgXIlVDRx0v1bfbKdYWaGKU2Oi/aPknqmvp507ch+xjBYaLP
efaOJ4skTiCdXa3Ggxx0T0znvYz27I4WXQuaPZt7EkfKLk0Om2c04PzDdY6tzAC08rh57s7ZbOQ4
T/MblDPgDzj3P+/z1RkNGgLiYqAQUNlY7Zb2uYNoPU04weqKcRDvL0fphc7OkZlNx558ae3kGELG
Yun0x9DEhhhgLWAg/gO4yh4fu6zkIsTCxjrW/TZyQslZNe9WENLRujLnSVEULTVUT4g2ioqhbcvV
uCIjb0vXtfxKpr3isP31JQ3Jb2ryWSl4+h5f4mctEs/9OOYRfz9p5n8grOcTLQkMeEM4pzdk/nXI
5/oYgOIdOLX3A+Fhew4VZcczPmBPa/NZ3Cwqav9VNoutjcViZzNPzzU0z08GvfAyekaTzsnE0BtU
jwBj/mlUuww8XVhb+dKDeysoqQNLc2fdVCONZon8+TY21jd5MkqDA7bMxeOiUBi6kZ8JuoZRiDvO
DjYUDnWhtTo7+C7uLLHQaFOznzZqT+USrNxzEVo2tNIiJTc9oDFQReNL5tlnX7Z1SHYAMbjg6eQw
CPyXmqB9bvO9t0Rw056q3x+M42GilDh6NwVwMrGbVyBSRBvJzluqEcomCTr5Qd/o753axNdgqLOg
+jF3T54ui1QlFIPNDcb0R3aya/dY5WW0HPinKevZE5OsxYQ0hi3WVQhqo76VoJs/OKV8cxdBo7rF
pVkZmmhoF8vLBQGUU6lJQ8QMlzUK+7rRq5oVCBUEFfQhaQxOTYap8uqR6LZKs8T/OzJtzchRPMcA
f1jGig2AkAwYJnqYiSVMRtMeukWfJcP2HcrFNS0RY1jF+DnU1896Z3pAZWZrI9Ku9RAhIOyvTL+U
GSyggIFCXQ9n3EdtF88YwXzAIcN5FYTv0untY9NsqnWmBWgsEUPxDuUwCpys4rx212FP+EZ9pglA
G4fsRS7wi5I2xDcIi5Xp/ubGiMEfHVP8sm3RA5v0GHlduMmKqwCTE6Nty8TWWOlS4GMb0tO1pBZV
3DQT+6T3M/4tZjsKXVwCz7ed5k84XdCRV09HD9JXRnSz2YDhaURFjGeIwlLkPT6SirEGLkNHSUhD
fosRgK2L+DON2LoiP+N2ghnDs4XjE5ElcySxSopyWzapzLzJceCdx9mczgltliPeUbkvTKbMDHJo
o9s8hPtbHOvQR1yTH1FjGAviNGbRrkgTgB3/QpKcwqFR6CnOfoZxvJPN5MpliJJopDD0JLIzLsy4
G3azHgbK56WUj1vztdJunKN8VNJIP5uvJ7ImK42Pd6YaJG6ATAHHQqsgrTWImLxbm54mZhkimmwW
W8s8+lP/w6HtZeXjOSTteyu9SDYXFMTPjCbRTGCNPcLoln7Y+Q3TKfdxYYFPzi/uigA9Qoqo6zbe
aFl5uZiovjETaFBcOuKQdmqBdKghV1hR7BmkpopYRhGmwHB1gk3IJLqZAgLOoXigOQiIEY/JC1HY
EuKEp8qmxmohQmG2gp6RKnI6m+uITqrZ67RKE7DujFi6MvmSX2gB1NmaHDXZEY/QQsohUlo0meSb
8qQHpkT4SI+hF6l2TdfshUlsUL4agQjDFt/cFcwuCU9WQJkwZtbP/HDVRLTA1PXINXFYhAyjY4X7
JrhrUsJYvIK/o3PK9q2+bHsWrRdBEN5i7rgpyhJLU5nxGZUYq+OkF8ECx4NMkiuQyX0tJzIH3NPG
5BYzHAELAYqL3Su+6kpUVd5JjPsWFMZP9L8S3ke4msPocXS27X5AqLgZlh8UZSnO/BaIrfOHQ3Hx
fjwle1sNRCviQewEfx7/T/MIYnDgRK5421y24+0gP0zz0Se9KhPgVL2k3HQBAOzZp6UnjyrST2IV
cAxYE0EXPqE/5s+HHEjXoJ2n4JBNBwMkfQVGJl2csbyRgUyDBbeNgAAeS1sYZV/hhVbuCUwZqt55
Gw7A4Bcz9AzOIATKVLuMxwYn32QXn6+ktMfMn6n4TyuxWLbvUtvxx/LEuO1SY4E9/PERvUCrkgUG
xyns5YBphp41ROWkneqHdAH/Z/p7ZXWlcR2j8dWEgz0nIbY8Cud3uJUHjq29npZP8Jba35kOaJGA
X68En23KOfoz5WPfY5gvNFoRpxc8kfQbylgpAa77lueJKZbQ1kKXe3+X2TRrlkqGDGpv5lscIu1o
vWuT9vPz0cbgGw7a7SFobJK8WkFRnoJry77n5EhuCoUmWmw04KDFiOMa+6EhYm+Uy+5PInyxusWa
BCzDOeETxFRNBs7cG8W9t6G+eT5J/0XdSyOwy+gFbeYnygkQqy7U6TOY8WTcdf/GIA8urcS/z32C
Jmc5AG93dR6DM5nl1Q8efmogQ2n45AOXHTBIUq1bypsvdDVi1DriwK2wkLPH2QxWGCJfousOsXkH
PUCrQfYGU1daTTEj5J0zvsImwMOWw0nh6RFwDtkoH1vxxdsUitSq+70YFWYr6TMZKnbJDS71fUcf
Xq9iH7sFCVLOVwPh8c5Dze52qSEaxA9VQUG6Wa3G2MyxOeEF3NMBE7OZygfrBSxmYKbo1S2RJqqR
+PvOpdrZRx4aHX8h3U3Bai6GCBnaWl/BhKYEzKNeE2OuX3Blu59GgK+B6xCYHD+SSMTIirkJos2a
tX3krubcrVgw8LZgfwAt+Cwbx6cGOVU3nZ3CE3MgSOSJKBxEv3I6fnP8FypAeulMy1ZDCfdQXdeG
EI2nDKKzTqT3or9Q2YVwDKACMKVvQa65Svy7bO2If9LKXAa7fht9avrrWEJZo5eDaNwwW0sTivVV
rNkF/YeNyaFyiwVDXYeHXWmtZZRL4FLdXscix7ZGk2mwv9thLEHOMivOo/ltVsbXDiWov8CstEvM
h+WdXTnO5VkQvr+EHdF6L+nmDLQvT3gmbFmOqrUOb037krOcSa1yFfbSceCVrls7QlEoGoWSyLwj
+jp22hgoUoeuJYcobsKKHiOQ5CW4llkj/3ZSAD5TCUNL9H/Hg3wPrpy/uRrqlmieAMbp5ILKFDWE
ADT3yd2tsGNWeuXqX5pficpYdxrnsbGZ1jNOd9zkhsBHOKXF2jsVMVDI1HHHIPU5QdFTDU75BthQ
WQrId+HXYgA2sJvce1D0/LLOzB5v6xACbEeynfpF0PCGnUvPQHH8tT17tDuWg0PpBAIcJyVJ6UlD
E6YHUyTpSJs+dNVdrMcrphJN8h227TdDaRJbyg6MT+OPgjmgEza8li8p9T8H50BXBe2yy23N0ADX
dU+2fJslhdvtn3DHWex1dHXfrexQ4wd7LjH0K4w2VDJxSjaigwQRxqECu7rZmSebTyFDM5GZhpSC
YmA6RkD3fwmO5ESG/c0mWISYk0eO19LBcS54Jt+C1ez9Y0GKUUiCV3ww2I2T43M+Z8pZ26JxXej2
IS5Mm2dDbAD5Raey318c38N+suJ4bTBgX52Izwh/FDfXv5xGmwk7WijbW4zeN2ej1Bicqz6oJmHK
DG+w1RiKFva/grJGccvMoTepTdYzYr6xCxPk0ifWuFAkiLooFOYEJAfpKU2kVWxxsRymv6Pc5SG9
gTFxh9DFp6LUVvpftjUeQgKx47Z/fIq2jfs5MxOLGeHeFWUCpmfOg3CYQbB1pwBJ5IbHG1QH3yb4
aDts37gSZrcoJdDEpMh7ow298tWPgqoycsjYz85VBEbnn2/TPQtUqNHMRm1BRhJ61Sed8kTGvJ6E
8m9VdkeiKr8szvabN9ibEEx9w1zKL4PRU9d9pK3yz+retpcMu4VDKVPi9Io2uBOhcS5+EnSLZ/pc
c2WjGS7Hs0ndOBEsGPTd+RL8eFxJBPiuPnET+V20p2uAl1lUbLIS/OrRc5HYvQy8niX3OGffsuZP
OVYheFnxgDPji1mRu47Oy37aY/taMqCykotjYOVwF2RgY6U+6eKj+Yn2UR9X7CFXeWZmrpTs1cZR
LRiTtfqxHV3nQP4is9MGYbAM5jyQ/8Y3QFycHfdLMSR6DeZYxdSf1Dd4SkYC3HOeLMlOkYJckcI+
+xAkwZfxwAb/nFpCOKLiMPapAiyPu4VkPtvt/5BD/sL46dF8oCaHPEB5hEwRf2xUZv8wzZF1LXM9
IEaLbDgi7CBTHCJyNJRdj0Lehw7X/Mu6aNNloU/zrX/CELoVHfECJs04jipR4ylMj7XkIZ7eHGfL
rgY+8kAdzTtqpr3UiInAhnYK1k8/BMEGUm8fVs53E9FGEyxpUMcpYpE0M50XnIdX0UGxxaJ2pOyR
HFV6x0X9EWcGBUA7SQabwEX9EPNw/Kh0AaYay8GbVPHFX1D8FQ0OqavNEbJGAn8HT+MS9vw8TCXa
q9tnd1lXagIr4ALDId5PJSjBuBcgpVow8GL63jL/CwL48pxpNjiyqK+1L7QeuhlbLKwBbrDxJYu5
iQ6Mabva51bFmMfbeoggzBknwYsRay4zD5BpSkfINrIsudjZ83DPa5nEOSmFst7gaopvOBqcPXHA
tAa5d0j59pu7NkynF+7tzBR6Zka9X9X2HeYMnUgySUPmoNS37sF8AKSJM1DTVIiJWaPQ95JuMiCl
bzUhhxBnjnn0loF4LG7/929QDTgzW6YecikZ9HPYCZaWozNvtbsDvNbYi1Db1BgBgr4VgHlRbclB
zZf+dULuyeFzUq6/SbHyiYaDKgtb4cW9su3AQdhjSn+SwuOsM6ca/eqFMNyn140ON9CE8LrxqIbZ
gY4hOQwkKu0RdtXkOh8z+EDlEM0WejHMxQ5MJmLgtx231mS7W0hNoJq0Z26OLm1db3GtJzlEEP3p
SUxEq+WvBZ0rajJQ7h4pqGhnt1/1Ahl796eubR3GIcb3JKzKDruDUJvxxNFjcpk2NLKOQOTZZK7x
USCYOGMi3aj+lJconxO3iFMuOaU1h7ZLlRf6wnvok0BfM4P2StkY38fBV8ZIDLFex9bHubnohX8P
uUUAOKRfEqNmv5d7GeWaUh+1ihp7xzgNJhGCMmLSVKcmaAudJUDT3KzesqiSxwlmB/eqIXDRBIpt
MFAo7jtt3k5Opgn+CIOgYXpwn0RhygMWqJzCQLWZ7wZYsPfQvptpK7JCj++YFuYFe5OZylE46r8O
dtQQ9/kz5FV8d8g2Y9WrqhxRfTTSXQ23+gSjR2jK1DdfodYnmYndQyntBhRunoVsBkPniGeGY8cB
crCLXoazqksFVt8Cs5SdJI6tqRYQt/x0D4N8Ay1tKH0vmJdEP515H/sKSr61NxW4sodGAGZ6YjDK
KFfGcBMA1IusGk264MfNJ0x31EmfI5fLOcmdmw7xlkGrWrh4/QnzWAv+3frpupLOr6tDZUAUO131
Y4SM2fi7lJ800xIdVlAJKFFpLknbG2WS6NDtHcAz9Lvh/UsAHqRsUq31dWcFwIfa57Uevq/aApV9
fNq/WFSCGkbb2n20b/A7KH8IlY4YWAPYQSv2efPJw2eSkHSNWtjvUxBBt5MACXJpFAbTc3IbuqmO
+H6zmJXj2QfpQ6RkZmPsokxkXQlLwsAJtDM+EAnWT/ShBAxaTAxU1FKswF022B6MEl0OQ1uTeaaI
D+JJLeACM7rw/tNGn3LdHJmSXmywvd26nJwZHru+BGRg6JKAMOPrP1XK80m6IWtO91owsg9ZkY3H
aMefcms4rE9E3ZB2Yp+a6I0UwEsE+2nf4cRdwdU8So8ZJvbpui1Ez5MMLGRfUyzEzeL+4NWX1iJo
87WhwD/ZJlNxKrGmAvMmq6B2B679fMlOeL1c4MHMXHJFyTw9rxvSyDWbXcxFFzXgX1LDAbudPzWd
oC/qhddhDfa5iEtM5FvBPiFSl+UpLZOzhEJ4OhpIceNI9DP5i336Ca1tSLgwla+6sOuKRnIE6oW0
xaRb98rCxWwoMUUZsaabCgNnhUEBuKoiDzRivOa11hLcr4TH0j82ws3zNfSjn3HqXZeIkYsU/HdN
j60faPxE/LoEVk0eGrAmKCaL/IM9AO9GLP/cTwX3tJZpLDwWqydBev34M+0n7ZZD9RsHh0ygYQWM
esHd6y0RgGH45YXzhUbD9jjIG76p6XkiwdC+wbGCpyKw9e21jDFADKkzARdri2j1yR9B99RszZeW
9x7Gnzdkcnd0hv46RHAaZT1F3uquyyoEgrpPdgyCNhnBylfN2UiY7w9q6nAYj9gp916PHso8YPdH
6vSELlgVdDA+o9WwPW3y/IGKL0RzQKSUf7ZGFqMTEDBqJTnUPsZQ2luAFSHbXlyvLwqQa4M07hNO
PtYIhkkKHQfXR6/t9iJILHaaIN8ry/TYL38Otmzk227MJdRAihkEyAOkm/l+m6kp4GbBtlN8vRlS
KUA/1Evgd2NgkNyFD2oTNyN++gdrgy6bvO4qBsH4jCZ0js63Ei6dxsoL7l1QYPvKvZkR72ID3j68
40jA9CyirtvYJUzF68lEeeRgX2u2J4U64otDuArsKqx0fHOhvjBSDCzphKeU8VgVVufE2RnuKY5G
TnvfueUrGADv2dyTJi8O6ldNlpaEZLIPrxrBNMGP56BnW0Vab+SykIY9ALLyLI+EdWL5xBoVyH4g
/9FjexASMrDI9Yg9m40D3XNOPYXfC0ECvIMx79Qq41yLFlqT49W7j2syEXVGjhaLpFQilCjHQfrc
ywzmJUpXYrvLKTNkKHPz9aUi+vHte6U9qMGDW0nLTGZrZ+eqfImnbzhKhyvidLWpXkflZOMeWx3z
rr4sdtbFavpigI70CIS9Hbjufz0O1uOGQrQosZF5Teip09yP34/XmgQV3TyxFOoMSQmOi6nzjHjn
H6Hb78Jkat7NNLxqstCcGxd5p3wFNZcoqjeRf1iswNxGkN6WwsnN2idKfDI0UJZCvnNVXlz04ev6
RPIh41P1wvfVmleW3uNDMMiE3MGBXwv4DY3s0f7YOuOO609LVGC9OnQg5zfGSWKAeTo96ZQO8Usb
YIN2DIP91AG4TQ14u2BPR3PUCddWhiMmQHn/GdKgSYExyBWCqhqZVOgieMVTnO1nQIw7gkBZw0l7
OJ9TEc5zGJVmCsMve0Rw0r3IGnV9b+mvaEpesFFnc+kbh/NBxg/Z9dJouLslhVL5MN9C/+yxk80e
reUFm0RBZ+O700jAChxWL+OyT/haI4kbmTyoJGffmsJyNFAGl8JiK/7lH56xv/0wb1wEOpb5TPq8
EEkZWCnnMYLTz36gMidAINPgt2OFivVdiWSfRqyxV+GJj1C/Yxf6Umfj4A8krPPsyVm/63sa5I++
YgqBqKQ+iZ5E/Rn2r9pAmdQqfAUZLcvoqUTE7OXV6T1hJ3DMOEb91AMPFO1uG9nuUZTqrBnbTt72
zNlBouZLGRqPjpZJetwfiemRkzRzirGBV74+rjEPKGNPda+hnGmaY/Dptc+D5UQtBqHBrwNznTDZ
LDyVVeJFi0KK7dKOV8g7PfCFEDRfmKUpqd4QCkFJ+x5H+u5tvGyNpWSh5Dikm57pgEv5UX5eBgy3
NmlKRa22hcUACvudnSf8QeN0lnlAEo8Frwslfe9+F+XAXeGUVI/FxjV4He3LZ2eZKWr0dkjBJoT7
4tDhWlJAPPX7Y3tW3ncwhzIpn75v3Ll+qAurEpXj3UjedgI0wIS0uG9FSK0nXde3N5HHaClymi2p
uCV2ALYD/BOIN14CYVsLbZKMJ+hWo8FpvHQwiAplLgyqPo6J1YHPCcFbuHOktCnplLKpxBC5mzRh
iyPtYa7Ca59nXoNf/ptvpINymHAeEh4ff9ci39O0icgp3oFj/9qCajHBt10K9CujwqUV/XGwBIRl
BS664L/QFEgT9HQp/9abqh8qAKfj99Ry4hg7U9vwp+6qLBqcwC3znBNiX9YeovnoGE12KM/9o4FR
q6HqbsW8RDxpg1neHs8qIH+6Ikwh1Z6y4nbtR8DQX/h+fms1J7gaKJUsUY1ILUMUjdPB1iSA14Hv
OSnetQl7E0rydLrOiYZA1hiNOMNmI4/w1QZ/jiA0+WFeh5CylDj+mqTNW6Z8KEmM834kUfVInVdT
ZZMT1LImwCcATeRRqtqyhhVwAQV1qOWT8ppv+6BDAIRnS6RQ9afwth0TSoVhrxhZwTu4xYM+ByAI
Q99ZLOaJr84Xq3mvb5p4DwrduzPbx8cI3qH2Om+CEEl/CTJSLER58GN9OqUeS2p97K+E8VqKhXAR
KeJXVq+heI7feEjIElK2s6f097Mf+XvpG34yg8ymUs+3hiR/fh9AbETmvW7zeCienFkhy+QrnSen
EquGSm47oP6xY2pXhTmYLwzEjyj85onYNglJnSEoQzocDzjKUPWlpktoRR2xk8hCHpepcfy65ahZ
A9oI82zmRJOpJ3JvunVVOhlXnYyTibJLu6/5iCX9UmE8SePECPvtd8ii0MoR7/CpHPtGcf+urvDy
bfKAq4mKZpjisb/pRwQpOPIuDjmbXugIDQ+rE2RXCymnoD5/hirY3ivwm9hZrU0ArvG3dRH5foIo
dg9/a9fZ6MpEty9B0YO6i2p7F/fria1veTs+G/RBsxXf5glIyAp+YsFjWkZQkkvBG/EP/GUcMjfF
PGs/NGxMzgW0X/XRFFQpJVtp4Fjf+2TRm502G7zU/MsS2MiXx5elomACVDMgkWIvsGkQ/KQMo8YI
unQDFUXKueHzKzvMotW3agqCs2hIQ0/Q5ZIDk4dH+KOIl8D/bbCE4dXs7+BXa8JZEOF9nhe9c9U/
YWPhzU0WFSTNbesQFZYvC3OQiI8l2Xzk/yeG7SZ8JkGTmZK7aDx80YdniIMQavvOKKtJDe3JSdnz
BgxV5g0dHHa8YLc8o43QMwle2iCOMBJrWSRlyWsyGoPJaPlYC56yO1Z9T6yHjIAAZzCM9wxJBDG0
TRpRaQmKVXD5tg1m4mfx0n6ARHn8YWfwABowRRXj6AngC5gfpkMuhSgVFVVj4wxgBXT6G8nDstaA
L+niTU6E4USvD6sGkRIp8iNJbdadm05nLW7vGs/CncPdBNbd3m3ejb5mNJkt4u1M/Uz4YiS1kH2b
fRKbxxC5NhG34Qh7rROtlQ0t1vGCXU7ca6GWw/E9QEadkkB4jmsqZnTRgtuH89AMhlsT3G8AgTal
3Wwc/6CG8sGDuzk4HGlazJ601j7PovsxWzoRBEL0s/0EQlZWXbRMiiXFpHzstQkRtgUY4a0Z/0Cc
Ff2lz0UgK+Rjei7q1ulv0akrQyv0oql4FdrYkpLDXF2sBMA9zTZ+1ZsuQlwe11h9paSdwiCKCZdm
qEzyeHchbPs0Fy+BBfJG5YUMIubj+GbKIpk95rqJyHiwhZxjqx+GWWvmbBPITGidUOtbeU44p6EX
iIB4R6tbJEgnYVQPS2qjjgTthKXILHgIavLcUMY3lboXNwBUSfdLs8e4wy8LT1GsdKWQMrxi7kfl
4/9vdGOVYQ8Arxj46/zAMk0iGlUI/fZU6Ldt43u80bkKgSS0TSmOaUmKZf9SqKexDS2fY2GqKXOu
nLF6GWGbT/j9jgwuwcLOu2Q7Bj0KnsVroLVuZHekpgupakdRYQWqizgtYsRDJAcBlT0QajSzbB0D
nqpXlK/nrzVDnhOPQZ2WbZnGqFXZukTmgpe/mGIIYhPqy1c2bu61zEdmdy+AzrQj1WSJZkxKOhnU
ij1b1XwgNh00ggCi7G6OHG9mL0QWsFwepXv304Bg3HjO3hkPdvf2Na1AIj+RlmTmc3iObP/bpGgI
RJ54QLz1K5pxLmzWnOVYtO7qY5zagftok0EO1cLp3/cS6QrG8GZSs+BH6s1wySXjd/t0QY9kspKJ
AwPO2WxfEn+NYLfWv4xCER09bglCygCgTczRkr0r+k4USna17JVhPyqRDMpQ6RDfA4PC9nSA/mAf
Sv8NmS1OXdQttqhV5uzlMY72CbhCmL+aF3zeMiIuUdS6tNkH/9gVBN4NkdElF/5c62Opw47hnpSr
dkEE67niCBeidyVQIWo3E11UwAi8R4BBZkKgMF6nyFYQw0QcGdDUldRBVijjB9O3ObfYDpH0a3uk
7FwbF0kSmEOyhy0Ee5/QBa34k08DA4AEgwR3ac2KcD0vgyYYbKLYdhCfUfvp7I05Lib2q1+P7TZC
gEimER0Jr+8HjsK4XoGQi8vDQ8Gdo39uuy7t9tFt0C28Qj0+6sW5xyuEvgCpbKPAmBhcOBCa19pE
nuFKSk/Y0ak047G0iVZ23tRpXs4aAWQd9ZrJ/5QlfC8EvBEtIvUh02zVzu7HEPgHevitaBL4iOML
a0BoFqJEuCR/JZn8OHz0QKCHLRTfeAKjlAlV2RyqioZ2heUBiBNMJMRvhB6xX78WkGWS5hoT3Dnc
nv48Gc+mpL19BrKRt5SOcjfa2G/Ju84vTMDBTgFehHP2W2NG5SBzj8v0FaoIZjdS5TMClK2jS8K6
3eMvnZrzNN2ZfEnNOyRkVCSq6iYM9dK8vXU13/l2KGKBQ85Q3UEp47wg7ekZgnRw59MVzmSCzgkp
zPmDrEH/2bAP9E2Wy+1Siy7eIgwFKyTASQuD9IEgHULLiffq5QFswfQ+qokfHTIJ+09zGw9227u7
K/BBb/31t58VVAvmcw8KjaH4Z7xnA554sQUm8JytGTrdCuXe6remRX+t2PS+9kEw/xGezIrR5ic1
yVL1J9g8D8ACeebZlr/qFq8uAi4cPoPr4iiNNAbiylR4OtidRr2Ddr+tdZkGK7vlPGJb6XRLX1qi
dI5nEg+MRSF/KDgGcgcC/c4xlS4Oo1H0njvw5AEBtO3PpAWIZW4QGcEXHRVueRqoH3+zBooyYJ2e
37xNO+fHjvwv5nivl5ciXgKJW8fVvaahoo95XOy2B6+ViZYaRejVG9qstVCXYn4I5ACKkIMydSLb
r6q0QH23cu0JjBXLC2d3cPi+vg/3pWmjmU2cMVRFKXs+k3/Rp5zWcsRkP7la/LHPluSawINrPF+Z
fmjiGt9FYDIg7jj6pb1Hbgt4xlQL7ZW036df0sVMbocjmxQPEd5YXeh9qrOhfeplBkutCchvVrf/
18CzqB+oQCLX+8JkGqejfpvRKBJNHOx6zjrb5LDmriRDPH6I1Ie120Lv6AHx01wX9rhOWULlsT/G
/FHJ4lK6Z8D7YULk9UbYsmOOEHQqv1JMlsWfGmSMcm25kJBN5Y2/gc1odyU4mJWWeginAFaRZ+V+
wMxeGbS9sDRSO7rmFitA8W/H0ubfWcmwMp8mDvuisttuxxmwNv9Ku0WKTGBqZPjCNTcUiKu6cY8O
b8VRrpON1csJ9kcSaUDLOCBTTvLG2MmJz5zNeylC8oQzN1zc3wJvrbs/MCtC8jLaXyEpID0iYsmS
jgwJM8GX9kfKC4fdrCHeDDHv6jBrT807MytMpqxLL1wY4Jfj2ekMb8rbkDqJuIkRrdroTIWEYIC7
O8i9krhkZPdqn1Vmuy0pTBwKuFbmQfez+UnI/s/al0y5rl/LPFIoKplqpYMb656nqi+bM6x5BERl
hjH6XqcczHbQMEHcBQnb7hRjVSEhrv3Tg6gMDWGRq0uXkppWgdIAbB5QNF8HMYHnHl4a9XWQegsu
+xZ1BFeIU6DRGJhsjvLSIKRf7pjxEvOeBN1Sj+mG+yRhEA/oGOzbkvkF7z8tzM7VBHvakbAd6VDT
17lrxd7GQbTofa34xs3VvZd31+NkxS6ihNmse2pTsBo4ICaHd2jyVgNMq6BUqaYwXRNL2m8nsZjo
1+KP2jTs9dByF410HPz5qCcX4Ksik1wjkwvvzh5V9JVq8Xhg5zeTKkd6Zc+JWfFtVWIuBdm3PZpG
aURyi1XPHId38Xx10WgmiIPkkg4lV9cAewgaEE8x+WdVYKlSIBKxUwsUlU6kDrUY+XNg7fC0p+qM
Fm+uGdoBXmBmt8ZHN0YK6n8B4wxvKXF64gODXlAoLMzSzYwNnYne4zMvSCCqtnjbPvvXsVRX231E
FuG6EZGgGZcNraR4vUykumSPfU3MOjdKFVhnfHJvXstR3MopcHa/1vVMkB6l0irhPB6MEKdp0XkS
LbNg97OuGiwNrmof8X+CiZga+a1A5NxmQk0x5Hwv4x7tkoSVFh8lORqJsqL6mbAu8jQkN+oJRke6
OCERpv+3YPc2+44C1qotW4JIpv90MsJJ5PoJp5wlLrzM3TXkt12HsujNZUDOZKM5wPZmK0KZOXot
5/jPrTMfyeGOleGFhtqzMCgxjoSSvjQbsJOye1Tw2r7z4C6IozXcgs7YnR5EjtJWWEfzY1vuahel
D14jjfd6DbHqgLlyhJwSm7L3o5B1RB40ITgPVjlQlLOTT1lk0vQ9S0JPIgzDVkips9Hm52VzGOv7
HJ716OdkOrkXxCZwodTV3Fd1olxStpUzsk69Lq8aTusED28o4mKcNpA5q86ZnUqNoZXuJm8r2cWk
tw0VktLW6Et9VuLFTsxcZZXJxIKaTVH5DzMmubmju08DLqIhGwNON3QQEk1XaHtUWX9p83l20YFP
tB84aE2Jxy+rssPAaDQt3I7dSdZ0BYT+c+YTENgAMU7BFvklzspQVsjHBBnquaejbOrrlE8KZwzN
P2bR7P8P8CgryOzpUGnzh93kaHS9q/OcU4nzLo5ecOk8lfdKXCPJxmD+VMnZ1QbjZ5ZFItt7NSjo
HTuqe4eOScbxEd3mwxd9cluG5VP588V+p8vMOkZro+7g5n7Ngmd7VAsUeAs0lxy2FSGAas2BVMFc
0pDJFmLoYOEvFOEUGt64ChpjWHRLCNfvvHbfE0yJIV7nbC4LoGoQlr2ePKr9/bND2XdLYI6aIrFb
UNekPMqNcSbBPcuJ1lnSSJAPcM7g5LdqvoQmoIRuIus1qhlfHj5yB9y4j9SmDSTESAlN4fzGAKRy
7Gu9QIIdqSxnJ3zSaA83n0J7iPI94MFe6wnl0ysonVMy2SEuLil+VnnoV0+0+4OcXN+OhNLaEZD6
Mit9oG+LQL9uqIq1kj6FD48xW0YJ7WVgc3Q0HlTdb5gGd7XNRjnqjNINxv8OtXUi9e4dVvXK6HeS
o0tTGIk7BTkyjbpKzoQBoLPLUgoS1roHyUD/JsgtsWjW9jG564C5oW70kxxJYATWaxKhkPOjO41r
wEFwm5R1AFVLrQkjjYK3vcUqK7xlRTrlLzuAU71BOwfHpJmnWnNOKhvGr8B+y7RUU1t4kGzJwnJo
11xaGUIxlWEe6sAO59K2Olt6uSMz2ofg311aT7tQ7sM1oMRQUyyMfbqsnwK/R1upzWWj8g/kp1vV
LscGaU5KT3LflTqrGI1lKPOo3Cf5o4fEfLjIup+ueDvqEDE4SxKPhc1CTRVgg982Ng+rfOgOJBQH
Nu0Sseg7RX6Vk0iwiY/XU3wP8vlurlLQyma1DC+2WnOviTjpPcElD10V0xONENDYCPD/czI1ENzP
gEFY49ZwjOX1xEsnNaTyOvNbXsss5mkM4pLUcDkN7q/kxXa64CSiX3Mnu4ZEoaeoJlV2BxOIkXWl
XQCRwOCaPwQFKbUfbzkWv/ddQ7s3ViL7t2mqKZYVM7vOuVTktpKNkkNflPtgce5QWWs4Gzq7Mr5/
9JtMvNI/7lD1kd3EC54LkllVWJU4SpI9CVibnbmAPrOQoZBTSb4spqZDxkA1NVGDNGSc6Ncc5jNT
bv/7athhGkD8UUy9wUQPn8CdrRoTJKLXx2j+ocs0340Kp+sfDue6zhmRrscgVodsjLn5wEe9bVqB
2F3SCKgGvJltPvfktjiCxIsx4ioIRwr4FnUjfTXBh7O4Xwmf4nqPWH8dYQhVq40Sa3oMN3MorIbe
oeqcQyRrX341f/EUud1or4JF2qgrWtfbcnDTfGPi+nWbDt151yXyFdnGk5FK0raVfsLR32K1u0s+
Jq05EWHUPM0BpPfn/v73PYdxmxGDuhgGPoR/NRXS0IeKH/xHth1DFVsoCa//QV/XrndFNFWGTJNI
2/+GoiXVNS1e8ac497ZY0eF1e8EXpBoTvUKLBuF8hX+zP6J0ZhlxCwQdEKxBsZO+Kk4Naah1HazE
eO8Q4hQ+cfpf3OO+/wo6yXhQtnqD12OjN1JdjG6Ul2oO11JbuTa8JIKJhkzRDIGFz00sbxwR5iXi
znF0XtCpHhjoddkbJcwy+Wgu15MSHbVqXsgoSSlcarSK73+Eg1oTNb0Q7LwTZnFlNdSyf70jXGro
ry8MqRW+rXZXnKSul+MDgX/E7K0UomWePPwDul59SHJN9EUeBt5a3rK/WdV9EKePc28wHGXoX3fy
rW8RrQAnC4MtMnhCnRelAlQcOw0kx5RQ7ruVZo3Rtn5j2q5ktEVpVnU+6tT4fnKFojoE2j3uVe6R
YggYhJFtfeQYGMLvmBEtrUY7kJ6FEC2YYdsJghLwt9mLJlebW0ytJcDxavCF3CGMKHWWbQNe3fqm
72g7CDtjldq9QhhlxxFGNAX2IWeP5B2TxrzEQqGWL3N/SHneOnV1RyC5XtXS9niu2mqnOmSuVG0Q
RwMhT+8wgKBBBFf2TornIchVoXoUd8MgRd2p2Fv2soio30+uKdZ4A/LXr+hlUGUVsBHog14kLjbm
a0knIkL+onh5njGHDCrUTZfWFyGUs6A+CelO+5r64/raUFi79Ra+2gzI0w5fOg6bz5QQqQYUY7YO
k56lKkCY1ttJtUGahOh6BgBrRFpfnCKP6cfQW87QLuuTF/ceq6EdoLuSJiYSSYTu69aICXLZRFPi
hXBQkAX620IT9EqCwzE5sFh1Cnfugb9J6UX6taDeHdeSP3HY3/L9cF5UFVn+Ude/55Wrz/UnOLyg
xkln/VmtyMHxqy6wWglMV5NSYf8A3ZFMJRbAoL9ae2Ce78usHWuPK3ZbjlnMj0v7Sd5MvhnzPzx9
2ZGXXgPpgtsuF+eZP4GrndI1mZazI6IvLFFiyBqUirkyZoxrp0uswW4pV/Z4p8reyaecQM2z8uKG
+4hYEqFfbKbihMLWYD0pMMOdcILnKmmJyHY1uqCtb74R2RyPpVlhCYCwj1pDAo9fVxzuyqO48Row
Qod9wS6ed/Km7mxlrmQXmPbN5EhXA3ptfhhKibMA2oTMW/bUcl1y9JYm40ixbDAEvauWDDQMEjqA
mjNgLYIvLNcUcjfXXPy2qAFassgdgtG5UlkT1f2f3aTFn56oPs6zUJgx9LyDrfvLweujBidLxMD7
qiSaTGQuo+Zny9meNlkz08KJ2SkeiTA3WXkZkWtLEFz+mBETTTupGSbgNoQ47YI5Y7G8lqIqL2G2
HXHbiCFPZjK30RcGYK+/M7Rov6cp+xLOBTk51euuWyVjWk+yocbkuVlt2jm5rars+hDilOITYolc
NXXRM4y/0Qw0TQ9fcAl+C9rIMGnY+tizJbXdcgi4nKlvG5SNR4u+tKCoVPRjooQeGXbGCLB95iSp
IiVf+s83+evafTu8YWF6Q3yQCSYNxt5YPRzcXzrl/Oz+yt/IYzhR77A+0UtMZEizvYYL+AsR4kED
qWr6+vCHSnD8hBs1UWudO3b8dWLmc7OXPWpm40Br03f+tFASny6tibgAW/CW/Ntx1ug4WyOd7bhb
YDdKEvxwSu+33xYAoaH80hy3pqx99IExDllarDP90Z9mI03Thdpgw39QUvDrTHWOiMvbohdcI9PA
BJSLJmtcnXX9S6UpESi8kBGfhMdvdez3KMWcEUewJ7pnuSy6GHGpJKZ66CvsxMErhxc1sYaJsL1c
2sBRkIbqz7cFLwoPrgoFGE4yv1jaXk5JgCxt8PncwMs+0Jn0l+AtzeY3Gfd2yHoxRqY/iXMG1bhY
ALmOU6CGp7DEaTyLRwvDzCk0wzhE7j09KHWi1hUHfVvCppoxTYXRxEahOwHDTPT9ezDYGuDJWawz
LYsXpB8PH43FHtOEZUUcG/kV5BHkZ8ViMsKOKC4kFXR05+b0pOdMDjn+kzuSxqtEWRLao4tSnAG5
Hxy5SocBIwspEkxAksZlUthW6FyrbGcvAOYRRrrV6zhyMLwGEdBvmXMd2zBmv4chk+SNV7+WvtUE
fI3H6Oei81IWP4mBr+RmoeV9dqIn5Drbj4bpM52nIZHBHKSlMZS/LQu70GoSQK8Vl/JkizEseUwc
IZOK+pUxTMR2Su0Ovk7a2hUxRq6/dWnlchAu4Jx7AEJdMzMUrQFyH6O76NS+sb6V2pGL0X53xKTH
ivKJMh1drQF9A1Os8Dva99BNiP998fTtUKHjs0JR5oHuiSP+/oQEpqB0AG7hXFtFBe+UAqxWSu6l
2zoNBJP+aN2V6i6GipRfsvJY2/x979Kx5Ju1bH7OvIGw3aLxlhP5uPAzcEj0kJGDIb1lMS52LKBp
TNskZ7woAVQraczpdSCi1SU4uNpm2qj2o90u7PTZIytzMEhFGBfSMsipp9B4UtbgGcl4uY6ZD1Xi
OiFmPjDjHfzbCfqPVZjI09Vm0Tc+Ix956ZCSJwXjG+Ys8ErlEMVTf0Ji9qfaU3QKOD0W//Ir8EuB
MLUBgocZulDrEILCGKVYsJV9vPI0Cfi6s/2hqhd6sMQ5+gIXgbS8Wi1Afd344DHHArZFNK89S9df
z9wxgVro6PvnkIC1giJCESKFCX5++3eYDW2tMfpXp13IjXefIqCNQvVdA13r4dN8EcRWwg6uiq4g
xeblGmP2okVlWYc3tkWfhwm/USmHCyUvIWrfPFYkzDbKzapg2+14zYDYKCgrB3odE7Acy0vghvOZ
y2VYLSUdPKAnPphn4vcJlR/aEiCdLq4vljUbd7DAf7YX1UnIADY/qkMyR/appB5ak7U2Yk4rGw9R
9yGv8CYklxBX7736JQ7fazjNx/ry1peQji/cetAcWY/LnunLanVGDRefqvgkyzm2Rj1icmP1Zvju
40YUvF500mYY9W4lXVX1fop5P5/IUkwxQUXUVN4Vo6orOxQ4rZhQXLFnF7alv7PkbAESg9GRZG4U
B9iM83WiJiouP26ERFSck5/R4shRl7UGO8czItIXG62ip893+GmErCtIpoiCH0nzxcW4WUEdgi2H
PtfmA8LOFvUGIFuEkUX6lEBYyFEGRad1hrzdgiM5htsh5jtf31zSH2bSpYBCr7O9WyQigL5m+xBp
CRGqqCz1h79ozPTkTUfGHIMdyChpXm8mUE9r0yz2Nw6BvgkRKimtWMeoxi44W7tP1e3pBfJxQa2t
A1q8mrQWdAX/efHOAh2iVaAXZjTDdlYPRXRHeKcemojDN1BgtOOlDdAd0EJ9CYMirtD4xP+lx/DN
VCd/xuB4BnkybK+Vozdf370qklW+1/z8e6eZdBCGPumov7h0RbUW0f9qe3GZHdMhpWLaTGwrGvJy
yUC1lXEMH8bDTCfIoIyiv6iikSiNEEKOkbWZWCX21VQNotB/Hj2Dimq0pPy9sqS24nv/07L8zRVY
PaS6nPO7Vu5nJY/RqTFIqkQNe9ElupB2LdimGd1aF7AsObI6NzwNQ0lpT29p01rZOzOjQOrDoZ30
agoNl9xtvnbFrEvRtSDflH3lKWVtE0BymFast6Cn/VW4vxjypIQU4SPjbJ52jpFoHZQXhKkARiGm
5wFxuF/Sgv/S3nfllczpVDa701GmjRHRlvTJUkwc952d4/y3XvcqYqVC8LvQrFl9aO8TrjKf0XGP
DM+BczXhVbVgv+/2JnMvqcngqcBpcp2uy4KWIHz7gY3U78unrebYozImQJbT+z+O90JHy2F7PQCn
k88vzToxEXOAYS4AHWWLF6Gmv7AZz2vJzOor7SSyAjquOWr9zkNesaVKkRihG43r3z70T7m5rMdV
ak0SZUdlw2fIvDAcWakoXEwa7/jwrfsEMUp2/2hdDfoSpEvLw78CFIAKdAcq2vTJkJRXX1Ea+xHB
5vGg7axbKnS5tl0YJxgdJUtE9NTvKb5kR3NnXST2J5eObkumRAajfmKIMUD5tmV5xFVIFdmHnnw+
H4qbCl4b9lfAR1d7Z9NFS1sS/FeJ4gzOXlpPtahWqWkzPAG4rPzOMFMGbgb9NJ4uRyPczIl2gppi
yIlwoqG0mW1N9xIx/kDd7a3sMKAdAxugOiFh4lPhzXrnn3DzkyZyeO5C2ftHQ2fqWRc4AWGsi/fi
xVs7HSelagTa/Y3AkOAI/N23A+i1MG1g1z+BigZevosL/RoTQFILsheArEGGUv9pm/MIDMp3Rw92
8bEBctIhDTxyxtJQQAWWN7x7O2aPRls6m3UYDujFQh0nVqY9jUs6nchOjAiJcbNuz2Sl0oYr4iso
Gda4S+k8cQMM4F/5UAMJre4hK2yf27Ljhnanb6KsSbRONfZHmoLjFRCbhkgv+Nr0i+yjy9Hr4w9v
d0KWLoocpPrxE6tICyc1LNcirXb72JxY+q+KzMyWeqlT4REQGdxhIPHjFnx5gwfKd0pRYk7lkRma
UdIEZcKxXvHaqB0VhDhS0+I+V/7AfMtrnlNqLQolKqs6OwWCtMHJikCHGHm8HS07bf6zHyg6Tp0C
wiCu2O6gBhC3xNyIpIUrXox8Bhx7+Z/uLiZAHDj9YQXZg/D4SOXqLG6GMr0lnRkB1x+5xlnSzPPK
T4Qwnc/6RnTzcsJgPqxKkgWWl51B620jWWFTRAgoMlIpVSvo9h5qV3ZioR2SD3uNqgL8Sd1PXb0b
wBmiIATjm5IfNnmUKLBSdcgnu258H6GrlhL+9PAIdM6C0SVYB27eWVLhoUa6vgvewbKUFvMLTlZy
mgFGS6S+u6o6Yy313umwJBx5TJH6f+135eg0/mIEFoSJfGJscgDmxE6erljMn2b+pjGGZtuxwva6
j7o2kAxEUqfBf9Z0G/02/rDHvFYz1edXSYGxbSH/E47BPivHhFNFu4RFe2MsnrvJ1vlAYKvovYk3
p/JwgnGQPoy552xo3IW7WtVjIMJExUI66KjXANjfzI2crmvICDRj101Y+FukEcJaw5cMKZ5b8xgs
L2ajUgmyyDPO+aEweEotg2Nv+JYHsZzEJGTKnsuZJG+NsNrkwmG5DBeSfvlVA4B3yxM4mC5bT1Tv
lr+d0+EZb4PmKif2fcXTscl+ss3VAEw9RbtkZV3LV8uTyk6eZElo9km/HBw7RgQMZcbhBEVs4TA2
VLTmsNR/E8q6v/1JHVVZTcHhlrNmgFbETX5Nfa2gNwoN6CssRT3HAg6kvyfsmO67PkvwZQ35uhdm
81d5C2drWlT7g9KDcMZq+KT1xe08JqgEharl19nmP/5QFsKOIbogJyWZ0GM1HfOzHJ1hYfG9+hbH
FHS7KyIZPpAnuAYdl2TWTX4rTb94IDVfjDYGGcBZFnzpdlrIotwjf+frU2yQWbnJeMLvaazz+7Qu
Q2zIyTFCR3eJQflzwc2ckehfNcxSOhtaHlAyVjF3hwDO4bTwUsmIz1myHowOyBT5gO0xajS1TxLG
vjc8X8wzHXStPd4LRb9qVdDFH0if7ivHd6ieg73hYY9vd/jRPsavte6lbwZHq/oLws1qp6AVV9at
l1kyMq8Bl3sm4YVvK/p1/dD7til4zs4ywf0MLfi5Qv4PYSFqW1r7qXDTgR0NjV6wzOLCDlExVtd+
49KlFU9ugJjerrmGAZn0DLl9UqDslR8tc8dgVpxjdqGl5hz0o1YBEu4t1qoXudwZndRO7AbUvGrQ
V/THQjfgHUqB52UlG4WG5o98F19RI0V5ZFdmSu3GOhMJlXJKe1407/XFxjff2XADN3XUyF8Z5iOn
v8frKyArn0NKVGKOpr6JYmRbDYHcLQj9nNie+fE/gxXVERd7Nm7mAjaN9k7dRHN7bALjuf+fzppB
oaJFfv1iozROi2UQ7GsX7vYSqlS8VBGBvftLEZ0YpdBpQOGA3aPLTmuOcho+gAECODVzUjoRoEvG
CvXrl0EBB7NhoWFI5hSe8iUsbSsQqKy4Rkv4hMkJN90iHm1qjZVK+wcpEsJhryv9Ywu4TfnB6Flb
NAhctjnATmfE9FkrnFa8Ul5l7pUxDtDYHRHu4p1XtG6YGoqiA2Zso3KnQZVPnBquLhL0cDjwfdcT
KVwOUj77znm5jRLS16i+qvQvFTB1vC/pGG2l3GsE9aEQ1N/96xLiXlmXqYuKYNNXtdhu31BKBCX5
vUqiZ0ElgQ90byIEoj7jvGShDScWYPynkZo3mNvHhYDT/vJenkIWEn0X2jQgQeEZ2c4BWdeJeRF5
LofBR+gAUmFSLGnnnGNX+r+0KyDjlA5dN2uY6UlHDjCWN471Q7P/8BfEpK4jq1Gv9QRc9DSTanmY
aD4yIU5npT8IF91nUu0xwuzoq3BFAUpJgwpNOE9N6NS+xGRXGJuFpoCNO/zvhOWrTAZ7a9/UWPNJ
x97eH+rCQtZWHVDq2c9NPX0ePxbUISp8KUYL56/1SQ7hOwcmKhpBpcAaE2JuujZEytK89fqiTzi3
xx6isi4qUJ2zzBn2s3oW03BpJZHG4XvYC68jUNuqR7fntb8SxQ4qo0j3rtr0YQHxt26WvbjefL/O
YAMeDqShTIks25hq7eO1fgRMdDWAtvmV9XBQ8YReRJJImCgTXxhcQI1Oqs99mectg/wN/X4GoLzi
mTxbn8DV6D3FXvwAS+8RJ+kZHSdcd6zizwcj/a5WIg7OYz00zslXpZzy/pnhGJnycSzyAQyIimy9
SpOZ7jz8Y6vqVqspMJIEk+dP5ft9TDz0OqXIa/7cNoRS4cO4lmggkjmDrvH6NnU/2+rb/FBHpJI5
MF7zLPzRdCl+eEIn+GaAmZ92MgGM24SJjCYBJYnffCxklm1DIlPmCO/StR1oxCySXbeGX8Y4qE12
KWHq5DT9wVha7w42uZzUlLAVeJPtnf3Ys47g/JKNSuA6WGaDqU8xTtK2ciWuDMiVFIi8g5lfZ7t4
+7rCmV0mYA6qgPa6gipkVsG0pNAPAVOdXUzmhaSrbxJIcrb/hj5oVnhBgVmtmUjz11BcZ9zJhTeZ
90xNBJrzfowtddOg0dHUtDhw8gWdgUXDTbzI8SpdfcOyvTH63nq6xBqq19TiuO07xUbZpRVUVdIE
+KkEui1RWv7AlBp8rVO/4UBVbglBIW9KKHJBxXzQ6SV3iylKbND8kBoFdiM/r5iJg72iGukfqhXy
+zhukdKl5YquuqHmW1I90HU/4JShVn3h0+QgjeWyV2ynbyC1/+fH1CuQR+eM2EUJtX3LYnHqt7lY
jU2qSsIjdRDxAOhaGED7EAnUl7JG5nyJDx7GWh0V3o3Om0FEjMFChviIkQisY978sevomTJhgYxu
YkEK6tDa6HS5+ZLn3tfwBLL8MqHvyCDtxqPnHSPTXobJPhJFBvZ59Clfizvup7nwJqDTUagp6zeS
w6ZOxROYRgGzfaSkO3Q+EGUzykGO3plWfbaokj192smzyEs9XFTUFTViLffsHyFp/cnrbAny+qOx
chDc2zheR1R99Msr0dF2cSNkk78ShU5JzPbzctlSuku+n4Y9P8oMog85KlcNcm8vSO0R5G4ICD2Q
3O01o5m+dHGpxl3GWceBAU2kXekLOqkepVlpXZVCcoIExFhL41QQflP5295N2nR6ut5wWOIPEwAd
WiyAz+B9YF9MwUrapFxs/pSCRIr9gFOQitH6biKwoXNEfkDGZF126+GbVqPrMZwmG8LnGjIB0fVX
ibnxP0GBWl+znnkIIyY2wgZKfA37Jm4ErVPnBOkj3pld6mpRLPl6z2LYuBV/2j5aXwlzhovYvu+b
xIWBgE0uABdV1r/6ILO6UMZageeYfsj+d0kDu5XOCk++wOWP9mJG5XdRJ/X0DlqVgw6IduB6IBo1
MfRs6OE+yiTmKMo8HcUCkEzbNE/Lsi6W9tzLppcyHouWlgn5xr4FdYqFj3qgzCvzAAUPeEv57Sm4
iQdpB0QzxQZI5nqsrf5hAC8cKLAOCmTpI5i0oHvmvMrwBLHGRqJrQSBbYVvWN8ftSl6v0blmjQ1+
h49+QsZ4FOKLqU3iGKqouFhwNGmD5DxsRUpkNVWc1b5m2D/FhdXaTQCefmhPy5UJPtuKgxDG0WyK
usqy/jwK0kCkjf7Aq3iFUoNYz2+DUbZjTmAxrQSDOVAYOTRySwtn/N++6fEh9SFkhj1kjsTiopaf
5xqjcou3lWjjgDDHBD7hTknZDn4DpXvv3dzPMdZLB0rHGiXGhbfl1dbOoJArNHJ77cqQZWtYoxWC
cGQCPdYnLRUJt7sR70L4Bs7Dlt5+trwLPm1rbkDsUiop0AufTKl/uuXCSjMRHTYeKLAESZg2PUE8
akNlhA6hVhJyQLSm1tBm4u5z4ZnKXBDxHxqgRuDtjp67z+7/ih9wjTWeYw9rwSJfLSiddxvJRGe9
ozyFeV14TLo/Exe0kk5KbQnuerRiAxhdJrhjAkP44YYY2Jsbr8LSSl44TH+QofKcpkRmcB2zlWaL
OCBfW+5A2t6z4ZyFm4vdi5DrMDLcmvk1NOlAf8ydiunL6/yJ6vKo4JGJzMHKBmt+MxFdeQEiprem
QG4JmabuW9daA+dyivZziLlMJ74Y6PWJPoHYzxbSBRFhGCboRZd0ZrO55nY6fv5gNEPSSWOHg6mR
CZP56wawOYhzQYg+oYuQyi7GzNb/3QZ1a96YrYi7GifLkm7FIAqKjIibEqY5fpjp1t04t5nmJWlm
WV+bPwUVQniYxxsqA/t1JAFwBDsRJmEI6t5kSAQJ7JQ9CnWM5gfjjr+1QbGTBpctPPAn50JgI+VD
aFdFtMtZoFux4PQNFpQHNwFatlC7smQRAiEGgfHQxq1DOrywpx9VDvFvxt67rOxIqN+X7P15NGvH
oW3ii8JcwBxZm+gEwAY0I4/0coHLuLJgqCXSCPZSzSP0H67+qr5QmL8trhb5ZD4g7E8UK9o258iQ
98NQbScKogxfIgVRKFfwqZKKkki4hkQ3ZEum8n5BkbYiXmuBTeJlNafjTwYFrG1FjGRofVJstTrb
VyKEYaItMueu3XPtx5UeTM4oRM5YrvbqPkYEXUDpxH6ZL4qo7FLwNpXAPoJFAjyC+abmNXd63ZHL
BtaDOe062jPX15osc1r9jtVJcPmPBZ5TocXumxJSs0ZsU3Hd/0S3E/E89POE1PEfO5Pk/2AxSI0k
UEQDwN0pqtSan5xWMUuztKIAowY3M44C+K7zzz23IIALWSEBnI1iPS4q5g90DqcM6GLKeSy9C6zU
MWxJbH3FU/skIkZsU6jrO5BSIBFtXqy0wwZIn6+ojwNgd67Wk/banSXstcR1KKhPW+RQpXhMb15G
fqJx9OZyhQZV8kIfSnsH5p1DeV9CHKpLlUFFWQBEg28X7NlEZnOzAkbG4mT58W611uPnDc9V0C/p
owR57EdUvn4fFjDYfPQLX6wjpR5HlItsV4sf38ij76qn/h/pjySqpE+nhZA6ukVeHlVLXS1lS8Yj
z6ZSCLQyumL/bJczAomAffyJW754/IOz2CATNLGre82g44RKg4bvfOTIROyDaAOVmx0uyyME4rMv
oeSsOq80Oh8Od+Lrl6PleP0LZmriHgbLdJjYvBxLqQQU0pssDaK6nwGVkRX3KZ9jiFMiok8rC4Wk
j8gvr63yDbZAdOEw9nNrE2uFnh1DWS0qd4g5A7/7FS2sA/S++LpkqhBLGCwQY25w2TSlBYxJzlip
3bBjUIfzHoxtIaYTk8fyNQMcnJGLXk/I/J9qJD7KhogvxEaht0FT/Ny95y/omKUFdV+/QqP7UclI
fvik5Sy4r1X9MF6Y2mFJOolcKLtTf/7rRccGsF6pidVjFt3d005Xpq6KPcJKXDUEeJrsLEAbrGta
yOgPeq4ink8rOSS3UEMPMuaBVaHSZPmbeNse6gJhJ0TW4pFa5rrbNfPe0iFAyPMsFgxM7L4zimgF
9RDGeTDOxERFUGKmmLNh4a3rrEeAVNhkVzdNDUgVXJY1LNL1L9wltBxM+ou6jA/htckCuwAg4FuS
IJ7Fbs5j4+WTocfNLAjtLXpHyejrhzZCZul9AycT2cio5riI6VwJqhC/Bz0GgkC4qi43g8Y0e8kJ
BysKAo1NFReDqeIUuen7UrVmiWXcY4wNmekIj20U0U79v87n21vDvvwhgbF4j9nss4jKGGoSkzTE
A9CphjIKKr5e7MuSLha4tqg+2+KdMDzcUoSAIq5MIdxWWMz9jv3JskNxyqMT9zGyzSMDzedVX5Vy
3NYQBBVVK+vDCRM5Mul8LH9Bd3te/VzdHrKKOaT/Gv6gHkl7XjdQgczdK3PCphJjr5RhuDF3cN9a
8PqnOioDfZxZqMNnPycJ21qK2m0pMXir1loeyFf+EapVdvsCVIaq0zdJASm6EbEn34J9FoZ4s0JT
cmq/mWmCDxTtUMYxbbnQTSF9WgyNgGKH2zTgDiWo6H//FZXxWe00k7eEx7RmtBOamRFjYJasj6Zy
zJMZ4F8wctIRFin2PXyarSdJdiNCX8AaFoFZ4MjbA7RE1fv9SlsKv865CBWVyUcx3u6p6qCWH0Dh
GWmDve5vWBKU9XVmNQXMahgJ7UpoRyT1WIPKpc59OYFg+LWPJ+k48Hp1xKi8StazLghL8eFwb/xG
YSYZ0J/dqglHJZK90r1Q87lhsl8DdQIIZxEB1Ypyq/9MyzXGOyOTdC+tIL6ZBnJ9h4i86M3Zi1ZB
X4JSj99f3//VmXnCuZnTwd5mnEPfB5ZSrCsOSIFmb9N4L9AX4IStGXNj9hlyancK0o3Qt4Fpj318
oxVMr5LGD2Jh7mp7g5O9050xsuTUNnN6OEjNldgmEbhPD51L8LWp9URecZPRZGszWLYs1K3Pszmg
RhRcnSTlPelO0uYpx/hQyYnEz568Sn3UP9DPOjIY4QYfKaqXBzAXbQaDNrNzd6BiJ/hGBAn0sKDq
ypBPDY66Yeun9bztN/cX7CsSu639wmS0HIHPxIigPRVM3HRno74UMEcKSVIt4XDCmWHueCK7Vt2Q
xFeLU+cc/r1ZSXnmZnTvIpGEGWK32Q31G7nnDT0ud54CTtbRQ5MXfpcLbCu1Mkd0aprBBpEY/abM
SzeOuloL6rtxfFnipCPnMhNopTpLgk0LJTJ00Hgqydsv/J0vT9HEBZe4PcwEyNJ7oqrmuQJA3mAI
ErRLVCk1XVmLDyJiDQBd5CuJt7tpY/iaDsOHeybRkyfCsf1yIRMmFrAJTa7pqayJwItxUSAOD+T6
SOPjadIHKhyVN6AjpBGL9gWX99H+iN0oAKPV953U5b3GG7lxRxxSOdihBwu/qNITmU469G/7r2eX
PBJdAul2TUfxH9vczFnz0HcsxIQ438wRisUNnWjp99ZLFES8oMYtvUZPT3fAWrbahjRcmI5nRBCt
DcfLbKs4e2fWOjf2JTm+S/6N6Fxmu1DdC+tkFTSFxU+njRZ/FEOfXDhifns4lu9SHhZPb4sJvTR7
24mZ6liXEMrDymKoC/PyqqRYwXrHocrKg27AZNzjNA+MxCqNahH+SgJuLNxPWh3H3kHxtAhSsjXU
EgT4pS0RDzu2oXqxqkJvljAhvCcFTLZOSVhIQxtJk6uwW2qZzd1hyFCeZAI9vjklCo9BcXsZFHeM
GciCtCAKOflI9kego94TINowlmKWxSXMtsPWoEg7hP4n3Df/P5fHKQbcwzEvYA44zyZDGTBCnZXm
iC8G4AK0tCtO8llNT0MzkuxzyfVqTop/swNI1yhjzZqh0bid+gt1MOF2+2Xi71knO/YECw4Dj2ZW
dFaQWyFV7KPsoEbVDqCh4PmN40GOfK9a7FAx/tlRavykFbadWvq1KjrWTZ4daTiiydwFipfFXJKV
29TskM4Rv4Pp5e2g9Xf/5s/KDyEyb9BeaEISYuoKYodc7NeGoYItPvIVUAatVXRFyM7dweE6qzWt
gP8HuhWaDVHi/I1uhZZw/7HBIA2cHFUMkTs+FXJbmx/ieOFKvY9yeOMfllpwO7qEFc7SgWo4HgdA
0GDxHYYf3Sf+OP9I4SqKZ5N10iVfqeclPE//6ZUE806K/VI3la3/5BrKkJ7B8oO93k+xOVOQnKZ5
8HlSzVatuyJhwHvDYiuRr+NhWGLGEzbjXp132rkKva8n5qaF1XHzgUlwHNN5u6e17ne/qJ7eKDOj
TLQ/joskk2KxO790eYCQ7sezqmA/W24xATZ6O+epDLnCML/4k2YmklyJd8kQRtedOWxk/fVdyFQ2
MHYR5XKsrmExy7pzb09ed4rdeHVKNRDZg0B3Sjy1ptTirvlt+qSSS1iH5+4qSPZ6uNYCxVn8QwrJ
MxL3/kUbCI5eF8cYCJnUls/O4c3xVRPUN8lID6KNPyLA2j8eGA650+hp8MvNQnmP9kJ2o15c/BBJ
OdfHiHGgXyL66uynUOqa3rwghkngKQY/r2anzMo14KmhcmiOcghFnuk4EN9Xwz5b8JBDzlgY07LW
xbcuyxXE/aTpOYLSVu76jnjPh0vTVjEeB1yPaycXBxhzWkBpGihx4yGv6v45VJrcPv1XIf5bNWmN
h1IBxSVm7qI+RDOQuILgWfqumAOlV7vermILRiygGDZ5IAmeLHa4jP50LfbOg8btEGZpEcd7kcWL
KlfBmcOgbhHkbPLMnNcazj/1K6qZB2PYM8LqM76KVPItG1msX9j/TWnE9Z5t7JbIcFJDbhcDZSeJ
8M8JEXbLn4owtg87BBBSjaIIFcYsutp+ewhi3RCYKjYMGmjdSYiP/W2C2usdb3UVaGJ/ootza+eM
Nnxo+gni+uczW1GzDOqrw6Ky4kx6uz9pVDTYJunEd+NXYuKdoI2bJOF5W0J8nCBj3LiByfu7CG/E
8G7s+krq5P2EvpPudua9khMlv3r/Ec5tJ5OTj/+1GXdGc4vBWy549Gk5dod3mc8DTHE1WDdIr8+p
7YXPgvZQpwnuecFVYqwathR+gvvZHZUuLGySNl2anFbYmb55VO6rc+v++KXePxjCt3nKiQ6PN79W
+9jS2ERn8U+hwg+zqPXm2DF3eP+eE3rDGz194C8OgMUd8R3j3ekXKG00TLiPl6uPaHc8hepGgA5e
uBL1oO96h8WVkR8FHoFgGCIT8XVA2MqUdmydEdAKmbTJb1ywBPObTDyr+VOB/Kr7dBkZHi0Hhvtb
OlKX8PbWeRAr/xWjMU1mEMSodA4c/Es32KHKJhTuVisa6q13qYCuDJAjMBHvsWxRfO0lH/7kwZHr
4odpQr4N1AQ9mn9aIGNVUcFOd/3WwHe8kq4JcOk9oteUReTjczPO7l8DonudbKc++1LPirLYWjlS
hDNR9OpwpVIP+qggIMb0ocYYPmzucHWRIR+Jbq6AIoJSMAd5N4R1279Y3CTbE8Y347RPTqI7AlcL
lgHo57qccEMwndnIhZSPisMS2CP0nwIaDT7weaxA91kATUpf5aKtO4ZW7N/7Zc7kNkxBFOCjYSTP
/yoyuY7XkflrDItDirp0oaidvFtmr7hPtJrAx2QsCVOnID35Ff55PH6ro57POSvUqB5AuJPFhiF9
/wgqLYCbV5IeEHk5MzsnAGwbMgzSUbrSO+zP+aa3Oqba1Amik/M/rVINtWnjAiWY56vovTnFofNh
6HBhUFtAWgGcxg16kT4N8z81GZEBH6KMp5/p+lo/n7+P7+qgMlj3MnMsrrHiEhloGEA5/3X0CBW+
qWEPbs0pq1whwVaDmjDEpkwXpIkIU7It2M3VxJLcvw8fH4yc5lRT6PzNvPjAcouG6gJ6whSjnuxa
LvEmnqKONTB8XJ03tZrpYfX/8ghCU45ru4W3/SEuws0oMbRAsd8ivyEkyJKhRaAg1zDhZZShwGml
n5K3suyl4pAeRx/RTMjXASREmBol4He/TAW7Hh7fWx7xCi4EWnYHYr0KbKFlS2jcewzNsY86XpL8
foAY/DQ5C4WpkWihbv/JTAfsWs0gvMXtgGxFWe4AEeoqiJHOYjKSpXateDKQOxuF0YgJsR4IZR1Z
F3YuWzqr1h0CeXmflYDTw+qtL/fDb7Ag6LJsj3OIklOXepHeryyCo+np+8kQHyYwFGy4GrOQ3Dbh
aKGTRBX9o/6fINSzoKZ1YekAtG6er/G/r3oiPOxzl5NQI0UtDSHC716Sf5kifx6QBQhx7eOEcve3
C7JE45honHhOWqxJSHPYlngxqmiOvn+WW62khclEW82WI2GCZOiAgJv2rvjt7ictzOPomxasSSJu
9WQkr3XT7g43EWZtAb5SrmN/eNsNWfBdNPEwRt0MsdVg8jNrcMcH9cQIRi4QXykQc2BtWzNqx1Bh
UszNQI2gjTxB3spF+fJNcXgA7CMveNT/YQH/d815a4CsRY3YxcJ6XGIXCUEnMGsDQY2UcO6eGXND
qRjgHvjcYL7FSkt3B7WEBC81K6Z2gI7Zx3tjSuU4utorm8GJwc2h1gGe2O8V5Mi9fWwdtA/f2l8n
egwkZBTKWdVA7PANn8eL+PcSoWCim46/KKqDx5G6mdZxN03VjSyqKLGUiWwUFrhBEIiYo1wHffd0
zDh0u5IgiOMZ13XBbMOrvAQ3T8IovpXZbbpi8h336MKPR6vA73N0+vhEERmBvT3I5M5B1g5Uphyt
El8RlU5pSYW7J4qAjmK+2XFLOtAoOTk/7pBoEI3ztcYP5RakJ9gCNaMNK66teeVFYMuGsOuGGWJN
62LBzxW+nuCwwacwFBHZYDNaUbzm4lYTEZ2Ajo0YStbwj5Ev1CEbQ6qMVtu+bMVsM21abfBF/lsh
jfvk66cWiYgcAmZn21eZRnyEFsvgifuqaV/zoDGJpzND9lPMmGSnm3eKnFHt2uRhfdAMyYsTYEIk
rIjqgozhG23+uuP9eKlWYPehUVF5a5xcxXsTOv0Af86LMPVA0rp9jS5LWok1yzlsTzD4h9H1LiB7
BIikOyoNlLmElCZKstT9vTWVrDzURcNQW2yNYyycQhGrl4IYfL8YXh+RAg6FrP8hysHuAYXJq4VV
RHjnKTX2SUhVFMkS5dPgDH+TF3q7W+xwh6uzsEsdusyI2AvVu3IWvxsszinbsPbpHrgeiWqo/37r
gjECowTn068ZJA8BdAAPSX1mR21L+DI9ek83rrIt8QB/K7ARz6PqrCeI6pfY2uG6zV6y3rl5MOwj
KTaQSHwZ6bPknkpXbpwKPkOsd0WUYqA7dUsgT+fdqatPLDiW7yOh9jF1w1RAja6v1aDh6vMg3gkF
s6PheGr6U1LLEEgXV30HhFIYgC1x/ZSpzzCIPhr9TEkM3wDQOXon222kGyZLFidlyAc9PUnN31O7
RkJE+GMwivE/toNqvGO3pmbSXC0d5ih9OIDWKm5SyjG2x5EzkBOXya8cpKIDHRE/E17VjFCUI3Sd
h0/a27nKzekT+TaukuOw4ionsUaM2DQMmHXb74gSllfc2i82Twh+nGk/UaZqTTrcnZ/ahbPTJfO1
8/XfA9Ghx0L2QFmS8kJnq9sJyyK7l79zTl5JK6F14X8xnn2k0pvU5t/4aM9VojpUyDeTWjIRxgL4
+BSQVWa379Th6oJrYCEeP5MOTivHXpkqlfEP7ZKfCs7QaAulpjH4OzFMUtxih+o0ZjJfMdSQBHfQ
hde9kEdhkOUM9Wow8s17qODvTDUN4elh+WUMlbQJomK2O5ogpAcQ0z1532Rum/TVZ37gcK7yojrx
is93CcPQsjw+WQvO87yuYzOMjluOw9gLRF++nVSaTvBy3gn7eHNW8wAOfzDrqIrl5Gkd47f5nOfd
cOCPmbJJC5hxihiXKod0lNAkfnWu1oIiXrLaYvkax72Av2jFJUVYwKTMoeuDTY48XuuPv1EHf3qu
3RrPeNDuI5MOYbxYFZjwJ5+XF2qM0fWWJWroAxBZuDhGJIfhBqnnwjTksa2s7w9IA0uxQnmk6G0f
up9l9zjeDY6Ra8NPNfJFnvKyXPEIX+bFlZYyB0hR7y4rJLKUC2wVhXoIiYakKXcGXiKYkUxHjJik
yt2CWZBMHQ3WY1I7aW4+PlOBgRU6KHfRWRAFiUi4h9t5F6B1KFNOOszGjkxJETwe6V3eEFYVl9Pm
z0Y3mg0agOWF+Ugf2/Bwtg6Jr9Gyx56t4tIyGC1iKHuoJMSGrplJ4OwHYO5I6jTbIwLlUSvRCKgW
YQAEqt4KC14jLAWLQeRC8g/l22ivLwBKEvN6kJEKcewqf7QZM2jO2z9F/mmLEZPuMAWX3Y2PDMMo
htr46Q+OK6eq+DzZ5+04q9zwop+33GbabGvCTuwImJ4zR+QOZGmRIHeg9l54UQyROfmBu2cPtt4f
eES3E2IzRdUSfz7O7QThPaQLqnSZ1XAKmjgD/jEQxbVK/nlJ9bk1jQa463ElvRwL1lpMQ3/RVYHY
oI0DJXEEeWdmrsEKmrhXmxLcj+6G1saO6qPINOJ3AukNgHqHRSpF4oGI+uaWYNVD3S6Yw3yrENH+
g1IcXZzw+WHioOcm+g8RGx0RjdvsKLvYpKodRMEIiBCAuevNE1ibL5AHnRbfUohDiUWLrcIaZhKg
mi7yrKYzmu8rxKlidkTH+O0lW2yMN+qxdpx3QGrTVyPbEvZp/8lSV0nJBBRnIOqPHDnVUBcM93Dn
chZY9OYipBlA6oQyRVDHp5FghPsZUD55/ZfLPluk5XhHOEgdGe/VFW7u6+LMkMw9OPVzSSCrRCdc
rVgbYAW2n/IvRYQ7gGubSiDX8EtPx6hBJDo8ZFkUpf11qy1yB73jYXC/yJ1VGtMR390zYVfnq43i
ryhMVgIrAAntc5dqhXFPjwisaTFaWKmffftP0HsOfR9Pt9mfhL9vjq0rSrBeQ1CX8Jmq9+sSRVZx
Bwsh6i6wXGA7kb/5FttZX/WJuidogIIIe79c9CeEsBsFZk5SaS0/Wbl+pscmfZxHm5kpiVNhW/7+
TkWTGG1VZf3dtIKIyi1eg8Rnd/9OGHCYslMCLaf9oEpRdsmUH9W/RCm+8t7W9Nr8FE0HVdwyD1Mf
QErNy6XQorAnCBC37z4TxIMaGUc2/P1JF6FgdEB7PURds6cBprg3uHUX/4Mhw3ZLxmNbUeQQ+uAm
t0VB7CxtzegOfqBUdB/uOZRpfJN9cG5+oSp0IH91Dq39TWON4hN2cZ6qsbD24S50S82KHdZAN0xM
Ax1zej561HIaA4KVSEw5ZBL7M8Y0cY8sfafEARsLy6VKGJ8w7winFo7Fge/+sAXNV7HPAk4lBLfX
SLGYhKoRlGtBgfHDw5gUnlWyLjVcvlzqq3WBnxzfjK4vjTnIfE3K2B0vJpQUAnFtJznWrrZBTMIi
+qsWFCCSKUU96Y0XkPoHVRNP/mJwFX/m3yr/YejbMaF2bveZ5U1/I26u9ul2qQWgIUATmXdGPJ5i
AoL72iv1+3PuS3qU8cVq0+Qf5VHIPSUAb8K8aQVTshD9Vk68Vch3I0Va/vPU3h8pO23psZS/8OQi
PaezhX9U4xYGqqfRCvTdBG8ks0kYKiN+2hfXpA/WKuTmTXxDRKE2hU/V/k575IF36H1E2AYbGthN
BTAEv8hor6AQ3OVYE/Nty1rz9JsV4ut4N6J19F7ADf1V8miEKmUUC0XnmDmOiOTGktk7rx3s1jB9
DlgGwT1Ev+L+W4exunSqaMG37JfZrayCZCZjm7vpXKejYcOzex1Ny8HFDJfhaMprRMvE+WK1TSRl
1g37E5Y3J3armriNLdTNolWMBXI8VdILEVFqyvQopj/Idmsxn7M5lmbtVfAhqbAlmW7fYt3FGPjk
PgCaBjSDeK2ibvw2GcSuSH4Hd1xkfLexP60QFZJ6ndJ3l4qjij7TLdr29uSGlJNJX3GkjAAzMRfj
H102vtvS3Ny7HPBWLCRlXghjYYFBaBUumSfpb/jeCKalrrOSuYNeLE/bH+fGEATAB34OVam+llvb
AgeDWXOADk7aaOba88Y0FlOZqUt+GR1SGYaQjOAWk0Y/6ieuUHtDnKWIk7sQn3ArapOwj6LuY7F4
Pw79DqCsatJnoVQjKpS1x4stYlGlHJFeYtWg5GfkfGPqxfo/Ec5PjzwFGCandNUxo7gGh13N4vW8
GMvzOWF66mhDz32wJMrtinAThu9dDU3FRTa2mJLxcNczwWoiKLeLBfuPeSiG4l3sGS9AnnYw1vVU
12AIjTd1CkuTPu22c2GQEV8IPJCESI7mNW0gwcQDkd/uII7RkoBF0M0RP5xXR1630r+Qy4whggx2
1QQRPOnM8cIF4jmzPUU2/z/XUyAuTYNavp0cmyp4Y/2EY6az+7XQzH6APLVbAlGlN//C5786HLNF
8dkuGOKZXWb1SBlF5yf7imTSbHifuo7PNZ/7scKM2F/QpxEHyqo8SwwJlLWCf9HdKptM1yQc7Ewj
ohdtRbf4bX11G1zAAFyUPlSGa3GrwBj+knSasypuBLWFxS2T8NG46UG+8ifKgf1VNXhJxOJIGBKh
vCwC3O4gEV7AO+YTW9NoFTngokYGm/V8mrz/3LvWsTspc66dpuMO2d13G55wAAHx+CYfTM3GgUx8
mUFesxFxgl36N6pBIboFRVjcefl9/iCsR7i2QRB/QTqQwhzuWRLVAZXI1uNA1erT0hGVWhteFJgR
xus6JYJJZd8nirbITOQTOHEG5qeFPvyYAiyzaKvmCSlNTIAA0gt/LQuNHS1iJKBuMoE8VscCzNMm
DpPaGOlcRO/vsjW0kYI5CuFr0V9y8ac1OlQ67kC9DLQMpBHPbRs+IkFi5ZAxPvmVxhb6ZHbnGbBf
SSSOBRcV40NrbjZ5hZ4ierhRxxGIFygk7vEw1J5VBDkdYkZ9d5kzZt8eSfbt8yw7RIzuk92B0V8P
0J3FSpu2gKzeeLh9nZG/dIdksu50pf7A9dDFujAFM90kQ2UjVg/EebLImFeM7mzNbnxb0EcE5Nkl
HQd05KabpU3fj/3qQ3O5TjE0AYJ9MYzXYXECxsn6ymWhGzCjGCL80XtuAVb9qHKdTmkn3EA14pb7
cRGKC6obMAJ0FXqq6t4EAqj5NXOE9H47Zu99ZbSmkPVA0cWBKolp0/Gjn9fZa4s8yZolOB5XtsZb
wh6kww5SN4TL9QCVHX7e1jp+RE3MED94dMX7APkdAP/okDr6V4w1jClQZaw6YzG9KSS01JAA1FOh
70nAZtwlufTnzw9GupMK6p7RSoWjWYmnKOq70YLLt4ED14hTRs0LlDpnMbCZ1Vun2VexkB3rHvL2
pwcwNic/1fe8UKrAsYxAUSOlvxDGoVG4L5kG4CrQKls1pHLT0Pzo7aWk0RDGBsQm+VE4D+cocOAO
dEF3Y4cldINk54S9iPxTPkqpHpem2X7e9IXq3B5rBbw8kEOAo+3mDI24YzOPejO2y00jhUjapWaW
JQWJT4yOBUY+WN98QzYEh5hdtTCG6jLHlQnUqOx77vg50tMUe+MDYDvCLS+z8sYut2QYK4C1FynM
fXa0gBQ66aSLRYDUcUCRabGuOHvfPFg4F6i3ctDS7FlR8SacIw/bs0nA1y3scwZMmJEfCIF6pnzZ
Gk0qQ6Z9bFrijsFZTX20ep5Odn8yI0ZGb3XuF3++h7/wCvxKHmqSvSdP+Hb0Iyv8x4jIFyQwVmNe
XDMME9DDtAYIo7NwUqR4eQxfY31eV08lc0GxALo3aUw7bcNjtmGS8skRHkgbEd7CM/pbYv7Easjh
QTmrdi7oGWM+jBDtZtEoqiBxza8j9AuxJJ7YLmqkgTDmaUNSqx6ecSqKzFMjyNrtCPTfXKVL6f2t
KYXSDqmtEVhx1FSwdRuo5/R0q20dNhOqDktGBG+axzzzWFaLLRcLSFGbt4dRWuGMEduPvcpMuodH
N1tngSZRAYYYIlvKkbyC1Gmkww6ef/AO8lZH9vBqtaaLXNeAlHCrBUcTb1gKJSPvBasarJP5PrnI
hgh71bO01hpKJ8mpIzvYA789RsdxB7u+6lR7EZg3M5WPnmILHm7jGirIi5RQkbrRJ3TPFiTCDS0j
3a6dlf6N4JuNhhPK0Tr6oOtllusNpTpt9owiJLnIjRfX4mt/4hYd29danIvfCdRF5ez8mV6XBWyQ
yQmcYZ4otfyaPpeDQNF2oSaispQj/kmK13pcw8TH4Lo3Fud8QfvpN55prjFUJF5EKaqdSape1jld
zIm/lJgwZct0V8cRmJfXBwuSIPzVmYibL/PJqbYJYvYNDMUvATn8a9yzwnQvQu83UXxGxQr2KNfO
V6lfT4PoXtge+6zlqGckaoeaqj2WR+2twm3y5vftMNgbg9k7G/ekoLg6Q1uJN1WxMak1je/91Efd
80EqSGQD7xxGNAIrLo3CCFtWPwdw8eWbGkHEd2jlaL9CKiO2ApMiFAbVQgV8n44nFpdNvDmF4fQ4
RCkNItSaC+iz8eU4DQer1uGIqiw8SqLu9M1uxx1BUNo/5dDSw80O91fHDrCQOPfHZ+z2UrlVjf3+
pZBiGPQJFuoMudZgv0UiYVhU0ocS3Y4qTQYN80EOo1YXX6p2YLKlyT+k55+7DrfXVV78fq0VqEWU
y0at0GAUGRjZU+s/WP8eNz/n2rOM8ofzhin0MroJjvytCveoWhdJ/U0SrBfqAQtJ0Adj/Yof8tmi
Zrxsb86UVzutH2U+YqL2bftOgCwf8zyvS6YUKaVoibQc6725Fni+Ok9oQkwJoAWNlU83JXJHymrF
G67BZpzP/6MFX6aWTDpko8bBO6SIYaGTdY4e95MU8577mFln8HyVqLzgOachZhT5PcTiX1drkDxY
LMdy4mK4yzHkddx/lu5+WFldxJTYiDq4r0uD4G+HKTq+sLKw1Tbn0bAIVLemrukVyPyljCy1asSV
XggcvD+122hEV/vxZ3z8FdHtYWc+33hmwG642GbJ8Ul9laXmjf7Gu/04k+WlatUtx/Ys69dC4zp8
Re7/fIOLvavd6LRXTWVpmTllZVTMPVlAJeAb0zvXtswfeE95eaH7xQEPNA15bVREQmxdRaFvASvf
brI6Lsj+toGvk9JG6P9qKWhGTU0yn+Ncii39FjEaV7vE+4y5nubxv7fcMdj8NIwA8ISvC8RUNETY
6M3p9Qe32DgwCMkZwOmm6LYMmSbD+MidIWuLBPpZpXJoddWzBUqMe2RjDDZkFcjJrzOuCwgjKpHc
u6AnvZA8uqgwyAO2qp+fEW3B27xWPG+qNrAH+67FfgJq6XGBXExmkXkZ/b1ND0d0E6NoLGUrvar1
YdvfD/sGifXh652E/wjVaqYrI0Z1R+4pZAjvWJPVNUpBQmdrmyUl2Ko1qVClVPGzZA02vyd6pkhA
fDjWUrwZEeO2NXt5NMro6fM5dKZveXvq8hPIoMaB4BPkdDYb/5sIYGX/Tp1s0VbuDhc0D14sorLi
5cNLZ5pouYlmYMac+OH0JGNRp3QA5dWn7thOZrtyBtMJrQlGwqj1WdezJF/b+sMxAXLxkugPWvMn
wOKVQn4EdU+rjFZZR8Zq5+UEPAzs6HMsIYXDToaXc6cVAScV8IQr31oZ8aIc6JzCiFuM9LU6vcmG
EmITu0MLpJJBH10GeHzuR1QWw8tETF6QN5NSuodfr2xUOrssP+JmfCJFFaPxN63GPDpboxzDocMw
sT6LtNtVc8+7FxIo6/hkPtRvv/lFi5RbZiMqzdemWnB485zfvPjwBvIbQ21YsAc8vWMQr3UqYkLP
tDqN21YNl2gsQ77RMlpAjzTAi4EQncu+F0KRH8OfZRoPmuMFVkwJNUK5YmgcXItGW50+HKz7uWk6
iFYrlwESM7PI8ShT+ckiswKzrG4Wq4iHZa+j6a2ARvsiEfDjfHovruHtBPLKS2LqNXpp2ui7iVex
BMY14fcJAYaaV/40Xhi6m9bUoApoNigf1/uu1AZ/cVT7qMuQgDYJZAohXeGcR1qWwUGKXW4/i6e1
gXGg/FrRnxLUjMzZBgx2s7w634Kf6tL2Ud61XgEYW4KWoV1dDSJPxzsQJjtX4Y3wWdiQ5dI8xeUP
i3V6jwxmV3q9dW+pWUiIGTbSEnyrvn9vPJbqZ7I53GjqTp2Cgd/nxKFzkxelgkcO618v54XCRMcT
iqGfwziE0kgAIVqpegPPUqghmYTjaOnwm4evteJ73L9yhI+uiNLAJRXUTDrGGxg4sg/oklIttT1d
pADmHWS+b0ZEiKImpGi+bFsXauLM8YdKYQKYQ0Oxd3n1d7JDaPbSSGOPi1OLagNWYSPRl36KHi2P
zaFKDI3WjLZnu8SOJo6j9vs8krlEneeKGbaSjZ5T8D0meudBYBBIS+TpGtfZdWL6Uw58nbwEM9bT
pThTGhCq59k4+VrH4Ifb0oI+wTGNIjEmHTMpb5BDCC66y4T3NciCONHUeuQSthoz+MK8EPXqnuZo
oxkPH0pr1Gzu/PY96lMUjyFW+SODmoPerQkSRzdVC2A+/kFFKSue0GzUqaj6VvoAvhRiELSlK9oC
3/B4ygLIWbT+7GwVNIziUsFfKCEWagmsXUEAgWgz+wrOIMwxxY2GqRIu+a23YwOY3BEhnhDVPtU/
08W+smA6157oakQPajKIh0AYMyVwKCqcvjboZIEIv4ASZVWaJ/ZL3nc8wis71IZF+z62jfEjCjE7
PlybPWitiJPAulr/pQt0pz4lRt5wSK46XZ2JymcMtws7mOGBTdJx1VSE2wAhHZ2mGvk0O67saMHj
3EZuYjY94Em+/0ah6846YDDkyNmElK0FYP29UMkzYDemvSKsGXcSD7F+OQ2XvOODTrk4dfsk3Ia8
NH8HepdStCnjy+tis25Smz8rOSjcwTMOHYryr/U2EcaU+GUvXcPV3qyHBS7sojzwqy+ZQ+RgZQBY
3LHpp9vRTvU30dP46rKANbpVeRhTnoqmrYzVEHKyTVuKf1apMREl2g+V0DL3TiyKH3tyAjYvapyc
+5pqYyX614SgbIevcJBkwFVpYqOg+x/8dLMrJdHBDSqWgxArAhv8BL1Tq9QIO7U706mBaizjhI9v
NiOLHp/cdWxbuAeoe2nyiDKTa591vJyKvHtvtiprMR/CFlgNRuE1P25ZqgcBXFrsmspauia+51gs
1O33o44p9P4YGKmEVKJpSaPDQIy6TfkG3iKKvCM2VVNhuwSi9D30XS9OloXmISEYTuW9ZyQGVWxX
CHPKuwqclBxjh5iUBQQ6g6Cl70vmlygXMZ6MdebSy1e08EZBi1MYd02fXr6QCMTHUU8H9p2pX5ib
Fbtq7hXtHWBUGcOE869lv+4aGwfi2RcERYVU2P1JMa6jffYqdZFZ04AXOe2iqbbGVdIso2X/CL0D
BiaatrthMJtI9dmWONT1Kaal8lWp4EL47ar4oY47Sx3C3nXeL1p/n7Y9By3KYtxjwwLGF6S88OKL
t+n89dmcgop5FvJbPxWU4wCR3tdbq2d6EYiRWDTPHQqvyE6rNL6msLOFseoHM/Xlj4zAqT+UQ5e6
VTqIOFExmabSqeyI8dFPyWjerEz0bDdYFviD2ZrbBLC+Y0PkXsa/JdyLXWzSFZnKBJH2bvZSihl1
vvRFDv+Gi+o4D9dtfRof+nWP5pXxcwxydH8knIgxOVA4Q/jRjpanIeSXbZi9NZegAf3ubWpQ0xC8
h013K/Kpw31H8zo3zDr1XnPZmdxWf/62GyDyhWX+UVOU7nOzsgDrpZ49MsJ3ABeMsRCMCbdBkDCi
sxh6KsCCmQedNSMPYED9ebw7TVdC6ksoPXLOti7JWmtc6z4knuqrEJ5c2W++Gkjx1LeUWLsAsPi/
xDBW2XGtWu66PrS0fQbzyUmOpmQTfj44HBpsnB3w4CTSSwY0lla6QeueMbsVoAz5/62+GZAL5yl7
r13ZGSdQ5I/nbUCSHbi+SJtkhAjAucN8p9rTPsXvX/MIkgZG+4gndVGmaN4Bnk+1CAUo7HGpP6l+
WO9/D+m8E0kgKbPVGrjsqISsMKl7HEw8g3FTk1+Wt9bZE6hgQ91XUt+QDi5TmbZfN+b4Uc4CzY2p
1PyREj0P9tbB6Np4f3ENRtcZXnIAHYSHYJ0W1THKm0qOG2qGZn7rR4ZP+vHyUUU59n7e1xWr+S7T
L4ZjhfoHbwTPQN/FMqsVmq4stA9Ha7WYDWrIj49V/f+g94rsEN5p1f73Tkg5i+MqfkQEnNPMkOu/
hLu6v/Pa7aE/eyiWD+yvvDMS3SqTY40GGvpINJ5ik4eIqnp86uKRKP20C1gXB8QIADsANBpxfXuv
WaTUwr8EQNf8ZDXfRb14iQXOHlo8b3tzsTNXiBtJM5HLB9ZSiX1i1QmPlcLoKEjrPEpttZJ/7/UD
shHs/aq+TtfYGeVIKLMpGXtAN6Ih1pHQPdZ0/zf2cioTsTqgi/7j6pPzAPPQb1SVcnCGnk9AF/Jq
rsoe4I7s2m283m4suAMNl9qdmUU16z26DKKbD4IVAUx+z/tQuQyuV8KxaL4e/TJJYUTfR/fEm1Vq
YjN4biB1g+JSXZMEHlepYCuvKXp7T9rz7v9xrYpEh1TUYiFXN5+qghZRQKCv8knJ+6vs1W1/+7QO
GwiwlqFT7sA1ED+Zaff/omfUpA2+3z4rA7exAlxqzqzU3L3P2f2aQ3VqNbXIXnYBCekjx/C9nE5T
jwLrjI7WSfIQOw8Cn6/kAgNBfERHtvbZ2LBIIo+lvWD/3c9ETZ1i7ibciuJayK7dnRreVxUZ0C6U
QstQ2ANTrq3BHL8/usQAYU6OCdt25K3ZLw+UhjvqjfUF3/q6fZQ+syGb7wN9f6EVUy24WvBJ3vz1
Oh7kUlFBJHG7QlWBKmXxxnEOPqmF4NUUItD4tbfAwyAvqJRoyI0vSPP4ca4mevlgDoLsdpM1EuwY
mpb7ueC1YcVgwBvXfiAzKMS+MC0Kt0yO8sxCA/qh62Rsm1rLFQOmSxRF8+LZOC6f7b7Z7RDrFIJw
HP578A7qibuQ2F+epaQj9jSbP0EWcE7u+pLEMhzDtZpu4S8hyzug6d48fxdIK2iiC+XIdKtR1jPe
G2Rj6sYLl+6bAk3OpO0tpNLCT4aB7XZWBB5o7EStCJy+g9vOzqJTI1eXO/fGJlgn1qKJBZSVVjQr
MWCsczg0sIbHl+WoJXyMYxRQ8Q6dbu+7gInjUlUuRz9x4ZeqqJs4QYhReSS0V4iYRR6mi/rablkC
ETsues3Qpw41YR0Uy+M402IKw9sUmto0i0ZlEPyryNq/iI7SSE1Yc7LMAwYRaNGzIezfKJJ7Ni1Q
NrOasd3EFEhqnE5pmIypadPYmwsNHe0zVo3lVcIdjhkaj4X4Z+Szwf+G1gtbgo4IcrTHEs56VW4S
IC5K6YuA2OThuv+I7JgAA3O2nFELsEJGMWnHnWwIHCdet26Exw2VrI7ZIjDeyXsNLnW6fv4+XByh
QShiQe/9hHRKMzaRs704ZEvxrGAJoF/o5JqzC/U65+MSzSsycnTtdmbvsmoQgPxvSP632fSJ8pq0
wdTK3sHdvwoP+MVxSWOqt5eBzIKZePIA7r7Gupg48SL396Q1Dw00J6Jo3ihi94da7SxjHSeytwUv
DxpUAqaHK3FBZHd0/KRnnJMCVMq7OB2MT7uHR+9rduZVwWnvgU6jCuMquvbBRDJJKR8qzTf+c7GE
vFNRlXkuiS6v/Z4G5QEw18IGgxvWRyU+RbXeyw+Dlwor8vcvKkC5yrNvAghbDWdIRywxu76kkz0G
HEFdWJ6i62YkhE2oDJ2KOXn5QpLApSGf5HoDJ947LQ2hdEfzTA1ufT/OqK8cL6jekLSAogQ2iYv3
5JQTj+nKHck/JFF2H3vKbNfBX6m63RDypnGz9TISjr1AK5DNDOGNLUL4sett/DoOsddawI1GAcL7
Do4qSTGWQjiQKVFc+9D9OzAc9zO/Ua9OBMfG0Hp7bcThgkQyIhc+bZ4sodLp0b/0bbhmYYdY3eeH
VcEtoVw6vFYn2e1hBzLwuU+dQo3r+HM52RblTGg/SZI5fQycJEnlsZ2ZjCh8joIHuMBNYaY48UZJ
9hR+t5gsMtUgrwMYPGp2anmI2V7KfR0Zb1GBwbvara9l3svHnrlh4DuSFCyiLvum+XYV1OnzqZmV
v5xH2e/+N2mS36K8N3tHmC7uTAj5tDCOaKUVVq9JtxQbl+n12ZviQ9vHXOTcdRe3yPsc8Y5tYa/N
hneelS4O8vTW9/qNAnf7OTohoQz0juvSz9oYWzTKYScWoXjRqcZo2E8MatedqalPjkdm+3A8tgQE
Cp3Qarg/62yd/5WXrIEqqR+lwYPu4p2H7qDFbTSJnq5XECIOePSDaVyU8P8QfjS9mCZmui3PvE27
t/5vTAemBhJR+VtzXBpbw54ljgDBtH9uoS0Egz1RqSClQ5qbw5UXGyw8YW+mVTs14bgpl7r9azbf
6BJ2C/xyLxjDT+TTO0pi/CXEyyU8oDEv4foOkK52WKJ4/b2Zbuwqj+2UQvWdMXeBJMtthYU45wPC
hCOrnpGoGyUye5U+6LZ0E1CKJyAFyNEha5Ib598suthGhHYY8w2hnx/5ClOWTGqRfZw5G76uW4PI
djfrVDthiHgmaK9RSfTGqKC3M7BbsRuYayoWNLEOrEThjs4GS/C9NfdEgpD8FgPR1YG+SRj2TOwX
EDZp2UNJbyXN7IWf9p1KCpFn1aFnFwdbQDznWs/ismG5Kwxg7ha4J2x/hTrZ0/cRd0syEYOapi1C
ysker5xg4KQltU/8ZOtBaeVPS6LV5z69Gj6rGS057sHVMJss+upLPSWidwtYymf0sQVGSOzwFJ8X
silDHj/VrHqPdG37e5P2A4tMJCzuy459jl8klH3nujYfOkpGjAlw01cn7LrfLC82ZAgB09jNNT9b
OwSh9po0l++PIM+sI5RtWJC/O7kqOYlhOMH3QBljD1fzxVvlJF3fwpHv5OISGT2/q8TRXRhYtuD9
WpPxO2eII5huSDdsksGvutg+1wwkY8tjLY5AIWfEpovf8jVsuZQpxAtefEyAgDvcYriCus+stAvc
rsOdrHjVYAXrVLoujNBakMm8CQ6Nk+VRiRaDOZLhpa4gnSY/IbOqtxdrip5UWHVw6eOCg5Rfe7IQ
mMhaUuon+YVmBur/C6XmGBKRbuOtQViDnWKDvsXa1zgQmVzNsKGWKgM39Csko8CFXRjPulQsaZ5U
P30Uhgo96f4YVzM+tWP0F8sAXisiddSZwAKzzuVhfjo2stmYhH5wc2t68znfFiZZOjLFvXCQ/dCF
JVPvMUaYdqDa7MfHfQ4dmH71yLYIiFP52MEooa9rgJ170oxuSWR7Ixx44GUMMM3HTaaXlcpn1s+4
soy3a7nOPgf24UBpuiadBfNkARUsgZqFvO4AeGv0yCSIz+HwPnrnrMow5wegFGEgmikS9I4A2NgL
oqF/Y5ZIpLt0bBY4iwnIEJVcguSc1pMS6uuwDyyGOc1Uu++JZ4dpZxuMjswToCdRiY6+4oqpuDTW
pUJYkSrcmjCdcBSlDA8N5Kkp3ylj18+xkTJ48U4iM2Xtp20BDZj4XUI7o4106WVJdXD/OtYuD6QL
0BbXzlYq+ubDchfLK3nASv9vh8KTLTOE6JtzHExiGJJqMnu9uOAfZmRbyPorLyFUeU1qWU/Tvbk8
u0AWQ/r6AISHD82sVUyQFtEYEnEVgiHM/cDwCwwgaWkRp1Ci0w3a1wP7qopFjcPWqcJZJDXs4/A1
LgSxlGHeVr4v+IdL4Rj2KjiYk9DeL46jBJFcofVa9gwj42hyC1Be6UaozlxiS2GVs7Qz+Yhbv+z1
yp0f2KrxlEo+8q57KcOBddWmo1WZvv4KXDUoe5rgCSZY8MS6XH/QW5x5B+lsajGEBuB6w/kMvoHT
Kt67nsn3tHIzxoHzUXn5hd8dKs7VSnC+JGJBOAoi8bnDDDmR+Sw82PLBCGO8huiBdgYT2KHy2lRO
oq5aAPoZEXLwhFIkcKUiRrg6zR/acJI0axIkhqKv0nfpCkxVaGT3TZ0u8UGsRFcSszrklA8hEtQ0
RXJiOntPn6Ip4sI9e4Cq1Tv7c8EtO4KrX6VFh708ELRb/KVpG55/K/UPt9Ks1iMg+X77/QDn4yoP
f2QbNxtaVb6mLtkATs6XZLgM5Vh6Ns9lDo71UsuITFHJoEEQ7GpDed3+jY6oQlgxHnyyaiaYPBkp
DKoS/wVPB2iXUxTvbR08jFL1bBURFNdjdS9DFXfJFfPE5cP1fJJ9tNi5n7ackl2nstRRp3S5Pzfd
Ggy23TcLhtMdoui9teiHRYuOptnKOz7b/fo8KdLfv9MzXbL/56H7Hizj/BHgniCWCcWEgVTYbb9+
tNyDwREEjuVnkZkIZktRxjbKAz02rpYG6+5NJ/yHO8/eY3rrfuWAzhARgLBQwyRuJzStrHddLl/f
t4LTFLVHzdywbcePX0IYqxDKZYixVT8FEXLm3mxt/baBj686MNkAMh1PoD5xU6r/ot3H4xn8MdJu
GjAmB1+N791WFtkqEeap+qrxOgWUc+Jg4x/SgZQOXfgifp6guUj9rqfvUlLZnV6yqOdaW+Ro8WtO
G7GaIjodKixtZ1KN7qqo95zr02QDH1u6ch6rFv7xXi284UyTnfxU1BcICG96K0Ez604Cisv4GW4D
Nng5M+c7oB9un3NBkIVBXaES0R5JkuJUxTWbXaJ9AFB3gGNG+Q2NQHN1WTw0c22LpAJQTtzE8ucD
ZVnSaXUZJj1AyyO9ao1aXaRiFYzGcNvQpRyL2BmD0y1gG7mXnu6a+fhDi6GpxpniSWC07jesfQ+4
fG0Z/8xSBfxnpIWITugoD1HAEkXbtSq0WzAhNy4LwPiEB/kGs5Wt4Uf/wLx1Es6cGG6F8seBNoZt
u2ZgtBNMJHeSDRtJ1EkFqu0rftSfKNENKiXQlQNK0ObBsS66cQeo//Qt83+BgPmkp0d8eSIfgmzA
nhmm/904YIjNaZidQBOZ3hjFfF1o1LWrJQXiXOzN3E6sxdY2QpSv29hr63Tn2ArQtD/+4qYgyUNI
vP4QnW9WcKfmFBXRVaNFF0Cme1ZYPegnRfKII5gL+S/Q0+Hfrf1mLQjZ6mMYpE5XFDLzduZBNa9D
RmsUefEI11jZ25Dx6xAuLabuwwcnezxya4FsGPWjeMcoBLqar1uiR6HElXeAC/aFuMzoCrTFHpah
G1IMDc8fa3/BaN1YwhqZ71B6oYj2AWElU+jikRmg7Y2zyNe9x0PRTYUc1WS9LKbTWmBBA2D8leWZ
ZnZObhSf3jUXknn01yqEefNiEy+jWHyNDC9FId3j1Xa+mS6EdAsnZUVhkEZOGzHrjptVYRK7a8Wy
6mp+2wj1GGXutG9Q2G3pcR6xvxsXet3PG1heteJVfR+76ydwSkQtW5qK6hIJAqzbXDLT1S2iIqj9
qsh1bURFzF1A5mgG5aQy5vOXBJahR/O8Uuxyd0+hxEmXvBJ1ft/PSPWah6HZXv40g9IjV41a27r7
91GiYsgX5YhIntNHALU5LSQQBEC9P1c3O46ynOJtQFeMoTehpTg3soLAW4Rk/d2NCl8puWcauxrD
eFIFlCBYvENHYMIBSzTC1UeUstYkbsG+lrGCaeGA1tNhVFvWFlgsG8eAeOcYaDv+gJ3xtKS4aBrI
1eaqT7EZYrkkNCyzDqoNE4p1tKLwQprzA6u33kQV0RE2aBPvF1Xdwsnw4mX6trQr809MX7QbmuHg
ReEcciXxncoJKbHZH8BlOCDNdE622eHp/m7Agv7yrLb94bxqZGoO7G4P2myjMl46tKuLBd0fSxRM
el3Sn+cirGW7QKSF3pfWeBXcZ5eF6RWSF5jfSHmehWjJX+VvMmMF9CM+QOFwgGWKzA2QPFIy/s24
Cm3fbRQOdFVKZ4Vi+MZ89bi7m3q97Vw6RcvivlMr7TXOE+E9eIb0Y1mCt5WFuW39dr9C1VlgN33/
dJhA6CDDI2OLPgIhZzFs9Wou+RO7ffvbnJs1w3YZHZQ3KF7d4wNPzpyY8D6X+4bcjxn59IXeusaQ
bVEG+IjKrp19u+0iCr2Fk/exhbGeoUmnJvcPKXWpZcgUYVPqFxmfTT3Ogx3tbZToafAxZKo1uSF+
6xHxqW5A4jSEqmxoQlDCyc55y/DCDIn5Bs0znP8+yS+vU04Ei8i5jyE8hfxdrmrWZnpZIhjs1W6t
/UEgY7M+2Hn4FXTDYxS6jWgPF8W9m9icuy4SHYLU9MaBjpIb0sW1XKM27KYZDGhiB3VNaTQo+EsW
kVuLKx+ml8hJv00aDge1koLLEztoEpUB97xS5Pa+4THuIjmMFaWacuJ0LN3/MlCIeK4U7fP056D5
SwMwAwV70RUZuL3fXTgcRZmIw7TbcdpN+Sdz9BMdQikRx1Nceei640KgLs+sGD/BaOiD7L8YjUwp
NpugbPis99PKMHrJMeviCtpM9Xi12okFWm5jGmASpJ7o7OHtXCXK2tKPoL1cFRYata4+aOWidRt6
J7ibhJbSMqLQxJHfqN1QneC0EMvWVdaQJEZUQRGOBMc4xL3+Iz/j8GyYf9kic1tFctImmc9oQy9D
ZT7/Bo1haS6mtNBqfcs1szAqPxRj++Qg+Y1ZQzlA5o2TG/g2fdErfgt+szN9sPvootgI6kzSgBiM
7cQ2vImPMEy/JuKx9rxz2jnJFtiU+ZOFRtrEauUZuZEy9L2AMw8h9LX2xgB49JuvAHf06Uq+VYrW
B5QPwBxAJEBa//1HH4kLmfF2OTaBBfPHOCHgtLed0zY1HUcmULKXEZgrBx8z5xjn2Z1OYlZ/2K10
g+Jl4cZIrWxJu252lNC5q6UT6iBVAtYKA0jy16XOI2qb87IpVwatCCnb6R45r2s04MPLovZ6j1W9
vZ/+0PU4k/UMLf5hVkMENjwhZF2ljNqooSbc13Yd6ZlBzRgBnWY6M3KIl4trimZH4BXEL65g3FqS
yGXRUEDtn96ofCwa9arF8FNWUtiCNWWKFNnzbOtQIVN3XAtPuLtCL8WwNEnfGYZafo5cOEI+ZxQK
2J2HEBOQ5eSsXOkYHl4u4Xfbq32kG1xOr9f2ZZLw5dM4CguPXME2rrJUxD5nMrqHRFmJKpjDnJXc
H3oxcvmz6sL1KfFBOa/kp5DTbUqbk/cgqtzxvB2+MfofWfe0PfrrHDzySL/Dj1ylWhCyXLmxHp8z
EK2OI8sQ/SUpsqftD1G1Vr2RmmVx7htWu+eY2NZ7X47Flzn+sy8qOIlSXR0D2/lsw7rqrg5qI0+X
1d08YcO7/oPEIYP36oGb/tOmrkRd7asRNNnpGLWfhMXKpuK0tS1eqXTG5yAZx2W2u5z/HSkzn7HQ
YUKhrWMdhr86zmTUqc5JmeQ2uwrbC/4y1DEVmbmKLV56lnScHX8/lOI5zYzPge4HXadJeDr/zo/g
OYgo7mWVJV4GUqg1EuxAp1Yb253ypYoDxhRAhMITjpGFskR/Sh2iiXdEziEeYZzBGS+ICLxS4fBw
EVvK0p6EiX4BxDJGeM8zclAU4y+84pxVLxLjYSbjSouK/H4cZxcIkGLPY4+DUM/V1mDRpnNuTDhA
7VdmJapOt9TmXUzD8oxEP6HQJ/UN0EcLLgCodfRJ6SueIMWRLy95vbsDSmzTzQbc31z7SltePQry
RCU6pvc7ii/QAC7AFLIYvfykPPsJ+0LUOBSpAMFt9HY/ooBYdLv/81SWpPs5qoq4G7SPKwJ/0opy
h0gFgJA8zwXmz7K5m91xvq3674UHNS4jAy4IOzh+QhQRtLy+CMqvvOlAuHPm+t1iWyUfbwz0ZlMx
fMSzFib6cF3cRY19XvLibM5erL11BcJdVgwdka53JAbKERST3tSZOk48IYUNg1mG0wyxz/dhEEQp
qE3J9My+YO/1GBQGp/oM/AxRjfbQiePVlmUpa2K6YxJlmbqAK10gG6uU8czekOrDKeQR52jpcMcQ
r6rvNEvuW5/FXa/Kf9agHInHRXU4a7Jfxt8djT8VgASkGUFtCqTd5u1TE67JRvGbg8WdHdR755ws
r8iqiB3mhevzKF6dyZw5b3NWH3fDFc+gScabR4LuLv9jznIQHmoUlgJp23jkGXRFEoCpmgDLSqb1
uWFIf9vNHP7p7JAP+/nfIoljU/83IXf0uVgSc9EI1kFBpSQ6Q7CdbdkmcSsX2kKPFJvDrZj1KGbx
opbXSMnzPabpzYXTXkpIbuSCFp5ZcC13nom0J8gru2+G4cSO+TZKUoVeMXh0Ig+LrJL5/tv53q7r
+BtsaaBRDbnjsx6H20gHZ6k+pcNoXouxkgLix9tQ4NwNKF8cYBRIdQVgOAkg0PUdD+8QZKg9Csn9
mcYl0OxGEu54gCzK43AUNPX64wHaDhjP0axA0rY5xG1nQpV18bYTcUgEN8dr2rORAB0DxQhWLC2V
wVNxvXWvxvozj8ecuwFEexn9r04nwOPo2DLsYt1Q8gqf6fiYO6pn2lCoG9FRB5tAPaTvxJQKkMh8
zIPIpvfCWVxGJ7vUnOzeUm4+ha47q4CSpoT0C2B3rhuNOUbmd6MiHtQg/Ubs5/NWCZoZlXGNoGXe
4D8blo2Otflc2KxhEMnbNVmzM8Vr7tkdG+vJSXSXCfwgxS+P71mvD03EnG+jCDHFLz7oezOu0FUs
DuXaEuDldRSQqi0/yP4a0chf+tHytS5QFCClf+QjGecJASy8SVxeCs53UYKuIeHkctVFBdwxOhwX
ELxPVZMCsy4Qmz2FkVMHG9ZcCUagSQw6UFDqkdnq+TbHzJiEl976cdsqM/91zvPdp9B2WHeiH5wx
h0fDES8YW8p/+UaB+7gjL5GPfl0lfmhb0hkABVeTXqCEyndQ2zyYSeFrwmnf/+J7gqQ09C0B+nVi
7vkGPar5bzQd8vK1p9QYnMuImaxPXEJZ2m9ZOK+9TRAjCfd432hAcv7+s1Jj1cv0A/UncaxdsRj6
DDwKqMZ69dJlMROD+1Pn+cUw7yy+x2IvmzPPMiHkK9KSXTb5yM/5ZG02gmBKRN0IdxXS0P8KHjwn
6559X4ZmwXD9f04c8TrspaJi8RztCSMiCY9o4p72ZcBX3n074T4E9R+hqDseje4h8g59r7l8jV+H
fBoCVizrK+8qfYP5z+gSbbBScF0MDLvzRYUoqPcDBvwk2QYDX3lMiNYKmA6K+FFbzrCZl778g4JL
ZRhjUY2Pv7eK8bPqzW5RbAJQPVyrC4mZHd1ixynrUJqmwnJC/2QcXWptybAwmykseQ38OyNfDZGU
4ihhXtQqoHZYkKkEy0RY42lGmdOLqCbqvG2Z7uxErccYGOQZPUrLUYcj5dWu/f0iGq6MVHnSjMkQ
oALUE///QVWl3yprLehVxfv8Vgx7QOCY+Jw7CHnSKv6ESm+85OeJP/fErRUI7pyA9K6VyVlSi87w
ZPbWZJHUo4bIigf4N1tP5pUp/eAc+RVfqvobp/AUTdLKWk1oGAX6KEFJON3B3nXNM20wIs4FsRnl
i260nSjuhVU1gfSeYocTTBBzpN28Agpa9Sut29+8JDSlCgYGsYda+G7sfrjdooMptZFkI/Jotnui
TxKlPUhfaSvzH914RODyLNS4etf2XCAX5vNWxH6RD00AsU19GBFgFu6vRVG4BLYOt23ebVSPAari
2F3NabB7PqvX/rKcGxrcwudbwPz7MAFGTyMI0PJ7qujMCgghxcG1n6+mFId8gR/mK8kXKkumY8Qq
qN7wLXCwrLJDZRMMfyNUW/MMRFaUGxqojuzw+NP8p9IBUOCaAKHkZphQqDJ+fBK+QkL/PWjSS8CB
h/la83UcYPBA2mLCjy58P72+Rge64MOhiTYRBMPAsS+2YsROM/WacvwUSuAAgGuYqi+kQ1MHVi6Y
lD4DJfYBVtjB+OOdGgYDhri/4KI6DKCBlR73cEjD9gmSGDA0S3T1choCuThsJkRve9kJ9lIIH1aF
m3F9ho2IsevcGKOh6aTikXRNHa6mnmMxAprCG8eeoh3LB4qL0g+WS1vKgXwdUX9dr6eyoLT5kv86
LIRl0moQoY2ZZeJxxzuRDS+6bBmZykN8tg3bMyKzna10Jn+RWg/x4WDgmQWnqedhIayZ14Tbb7VN
6hzvrFzk99h8g237UdKUSO4MCTjOymAwbtIY1xf67UZoeQr6fV/tER4hGf+OvGNEXiZvxfDb66Px
7WNb5LoUBzxa/YyzxAUPMcAlRYxqsajND+/TmQ6kRprVpusncrVbFzajalSNT2F4PI2DhD9vWvhX
GP7ixhpBTCy0fK3oZf4Kt6X8x4KYCYHo2L6swdlb/790hgi6ops5roSz0TEkLFWkkeSQKVR7Bj/w
UwKnRS50iw58CDA20s8fLhYH2dvGnIVsU2qxyUneh+mR351ivoFqp/znAMeDG+OlJC8bSCcK08Ec
LweT5jmYuPPgEbga8frt5CNBsehr+PujcN84uTcjKXB16O5vHLXitvySLq+GSKvj6XXn0zWDk+iJ
7eZSbpL1/p+nJMLU2yMeNAzGZDNmfnbY8qkRaPjCK4ihb4H8m41ruDX7Mxxief8ikXlO9WX5H8Z3
NONRb8xpwnqN0VGfj7aC3cm0YIIe5MZ+UkwQKgL9Uqjvjv6nZj7HTV3EQrFNIh7YLxAOpyrIwmDc
Cieyj9YKHIpPkBLnGKnGIHez5K4pEvC4/FhWXU4Fk1+78g0FogM5c162wEi0v5gymE6Sn5ILwX02
yFlB1obhpZ7PH7ZNx+ClKDHs8yevXwLWMNhQksXL+FJSukiFDFqnoFoPJNqy3mNBzJlkHCF+Q3vc
mUDKqgKqXuOJMxnvc40WiVfgbjXU5L4/ERzk75Y9wG0VVJNixAtmrrSABjXkGBRTW5LcEvE4Eq+j
8lN0szh/mBYtwbZaf1PbGHmq0FscUAa0FPnj6D1Ay2w4fiFyQiLHed9smeVf3876fHUfujDT2f4A
kI2X0exNihJ8Q4z7M7JRdYPTjrKEZNRjE3YYfYQXgG7RncNZX5aP1k4lkrgiIUlC5RPOGOCqq8oh
NGm1Rf4wtTP+TNURHzKogRKEkNzfaA3KmboB6XDMUCrgAC22mNUpEY5Z3PtTrgJeaTChFaTElb6a
iAPbaWPYmqswTecjiQX9GTIh+MqR556UxWmoL9oIZFgVAcu4Zu+PSvo2e3Bi8rrSL1axsxt7sWeS
rEI6rXRRKftiA6g/KbcUX5b3x/NPLAhAmmeoLRMDw/rBpSdBkUjjXamTI40tGsOUzhxhcc4k+5x7
NEG57ve9RXZTYulH0KQwou0JZRiPfnp75eiimUZ4e7MwNR/3nJtlN+j3D2fqgz3TxdEr54ljVj7d
EKYqyTAFG5oenaRf4nBWufVJKjEbUuMT6pbmJISyq+R3pbB6McWPJL+Pj6/PS8RO5NFgLGki8Mli
QOJ3aUDm20p5idcFyedq2ymITO3ek3ctIOIA/oskO/qy0qhFZ78c7IK9zxTKUO9aO1XmMYbL1ues
GI/O4Nzk7Y3Ih8CepukvM1ll/RNNiKlmVCq4H+f7MHWs5WqOJmu6A8QnPw52nqEsws4NW1VtUnPX
TOZSa2pXr2J6oXKs50wrjtteZfqgnBP2XiQU6mZc0DdNwbAJ75gRgU4DFDS1lBIlKLzgR8ZIKMB1
CucQzfVlGtWXkq3tPztwSYKovYba/1CFRXzZjJl2SlpzUEks5McFdCOtqc/brmjpy6k7/myIbwmf
Mkqh8QSNm92qCYt5ee3R+zcsNgG6eWEH6CMtmfWAI9OdRFrw+GzhdM85b8el/A3eQoMboAAT2N5z
tt1HTncKmEbSWdTwm2H2gYAtckgOL9m45blc7X0KaXe0QHjqIdj/8aUb9lnqQdJoW8cjWbIpHGyr
Ztt2dyzgJLDMdUxufzL44LT+1vY1IPODnf9X5bJ52t9+HLToYo+V9AfkYcVXw9RmLbVPOmqoN3R0
4vUwHcMrUFDznbARNmG8II8iT4RHS7XGxX0S+owOobEYE9KGKLx4X4OKexAKUdfhgtG3tyP4FiER
RSCeJ267Vu9n3N1W5nZ4KKc5g2MpHJuTnsiOfZksKgWkCB4KuLztHV2FAAicD/YEDiHQiS6x3Q+i
iCs0JhRRLSlPb4kldUPKmK24Cd4O4Ue6iPqKmQ8mG+fw0s3t+RaTncb6ylgTO6FHUZ8/bhH86Hjk
/17v0BfYiZgJKttjBhNe4efFhOJvTF3yxeMeOe+GM4n6iw+eDYy9DVZ30TBXu6B0xHM3TDSKV7BE
jiiGmjC94rRLCXbdAZ2wXj+tOZjvujgKfoUNyF8C6iIb/crFWMyTOERDgtsudzmiGP4pDHW7eKzl
DMpceRRb3UB1VEmagGrZ5C3vltMVKPi0ZLrw8wyW1pmSazfmzcx26PqzF+CL1xYUUtuaGUkvj/DX
puuz/MiG0mw5nGVSjiq6pNY6y0/EYFl23/km4IPQOBxFSTxf0V4kE/yiKm58cfIaJRA9xmyHZqJ4
eedBx72j4xrDPRLPwFc0wCbnnoqecID0FlkmHbzNPgnDFZ5SvtJtTvlLHSF+erQ/qZ4TrdgSmcKG
cTrRbk/o8xxY+9/fhNSaQEaHchXCiw90ecW+gL9u4hfRSyeAnzjAC1UxfrffInxSq4316mw2hXyD
LhYYNH3h14NORUGnuwHGQRWb51JQxU9MvAfO4/jdlbAyIxm1bJV1F5MD9uOpy0IGFIrfiIAE5yV/
IVdiP+wUfXQD3/dLQOON1/RNHiCeo5DcE2kFvdfhG6cLQe5AYTmNWZhqstn/XEGCWzRb8ieb2RuO
qZSMhI8ZnxcsVGf3YmyNW6PA/pfyM2JXKx+EeK/gZX8lHJhaQx8U0skz2OsAC6JtD2OyGXz2KE/h
FFpJE5SH/hDaHGdnfYoUT1IgOcxnOOZkom2yXhDf08ESSRXAI8lCpXqL1GUJlWoP96a0g8Ha3+Hd
JW0Oq0Iybu204fn2bZlZwTdcg5YJs4Ohu8pCpQ9Jr0RvNc5ycsubNafzvgI5fL8QTrq1NM1Fx1LU
XS64GDy22dE2lKuuE8D+C9yTLgzLvHfOwwf2wE+4fsQauJhHaY5WDnLj35BEZzp2Lk8ulRklZVun
nDSJ7sM2nJdUfKY2iyPnaXfHVSYIdcib7hC0sfbY3J7RSws3qztf5Hx4v9/8kBF3XcfsHF/2ueha
p6W5wWzFz8S2ayPIHcxE2lEFm3Y4a1ejBsB8DqU2gjXtNTCk/evR7Er0AAiFsj/6YxVQWWN2bBDA
EU3YqaheV7Z7P8CK+jDEV8kP3GkFiNj7zFN8663rAR7LoSc4710BvW10dVJ4sm20O1JHLQhcvB2t
DUk6P5sNyAXK6NSD++/qxqWR5QyjSYMNzIVDkg+ewIovCZ9lQ/JfPeyQ4+9GJzUL1ASdaOuewoZq
7lMAk0bHujkLGt2pcnHACLTANin2Pbo8w5UIaRR9/X+0BKAPF06rPlpKgNeEnRpfWfvW5nZdGNdz
k64pOJYrgD2kgyyVDfhCSwUVI/xbgXGj+VH9qC8zsUnoibZmHhjnYQnRtUj1amvq5Yunflvogbl4
3VMabAGobzcZSsN9Z/7QdCIsk1bJDiFvZc7KSTlUgTT8MFgpMQG5wscKSvFiXZfdqAnMNITxfcKZ
exu8KOfMqK95uLUpih2H55+y6wds+sVaq7bjl4m7q7mcwVsFOdgB1bEIYM7R+dLQTXHN8gPHrZ/P
SwEUKxJJiO3Z7iMJtHdQP5+8g3kqYQOVpgk/zVeXlJ8VMhe4/A4HZG0SrKksbkjq3e9oaFSOxVmd
DggbKlksUajNZHKAhGD3XdcyiICntR/tOL6mHr2qkq/q4OCG4ZyYzi4wBAdg9jSGfJK2PslZ9xcD
dk45eyYB25ENMbx11ENALo24ZGMGr1lzsMvmohEQFnmY7+mpmkjI11AP8ikWUo0sETBqRBqShuCn
U0ybA7nEfLpxv39BBJUcpT65hJCmcZPhvZ4wMZCMjMeuxfFV9dzvhCOhsomeAqzMfbuJCBBzAdCN
d4wL7s30pggeJia2w2F+au7lUhsQ6Qkzce/Gxif6g3TgA0FD/M4T1Aaelf0mi9PAZLWLX5NiB4fU
vgqsMFywx2mOw7S7smDpBy7mZF1fcpSclJ7GPrOsZVrBrnHo+57lY3pcSMf2i+91mHNrXBIRXgXX
00BcZ9wow/RwCdVSP51y9pvl2qhkSYmKvY2cNovNA42bJ6JHjgiO5DP4GgI+Vrn7PV8ohk39/CM6
38sCLhdlA6LcgZYlbq5wR09vvWdLvK5rGfaJQWkTjgEF/KmRXkbexkUApkG+/2Yc4na/8YIUOp8a
oT0jgTOrImkvNPbJMGTBdPi2dmhZVMY8wK8ySHktCkPQdI6Bue6Q1Gek4A/NKO/EH3KbRivpjEXK
QoM7b3GKWDGZfpqY0rRpIhqJDBUnLOXDZSwOQhnmNUqC92Xd7kB1eaoP2gfYATctefYKTRcKlOoL
tBmnda4xULe/AOH7kt4FZSd8o/A5nXF+9TaRxv/+alBnn+eeea7Cb8tT6odhd6piNNm2qc7Rk1eg
b1Km9+HqhKOgbEiOb1lzQ+k/J26u2tcrxLUO4tkPS2O3p+st7oNaZGPCWpQNH+plmVO2iFnTMCwt
rdWsLu5cRXCY0KezJ5V9e0TGnZJnxULwJU9RRH1bAf1p58Gbo4ZmnKH64cOXSsTc0gVwWijr7yjU
W0Qo7jhTMpmo41aQEh1Dq4Nr4KO8wFAjtt/YSV36slvVrlFaCUTHMjKMiKGy9Z+z7TfEApHYy6/U
9lnoV3EYVr7Sz5oLiYdBVsUrpI/vXZ+TPjirtW4K6uN7gYSFnAW/uBWw4oQ5CNGcUFNHspQJXmmW
ooBL8U9sjTLtROJOQaijnmm+mH+OZDUzbN+Oo+mA1FtDNGOpMtXlR6N0biwk0HB0IT4GEqhRfh5E
MYF82mC9nwE/V9sMnPorXHkhggWSokezD22yZeLrCJOGdUeWsrvnIGUweY8W7EK625uNKoxImJ1R
iO3kBLAOOyxHntQjjmSWOBcFxwKnb0OMf4xs977ddZ+MzxM+omR/mfELspL2NKifs/OzeP+T4gwv
IEx4nZyq3qluoUQrSTSQiPSopoETqAiV4NAoqQXlOaMVPhN33loi/nLWSaGcgBXwPpOUgJByOGlC
RvScPIeRsgnooUJV1vuVYsLosTJIQLbkljKizKjPGTNoZwYnphPy0N0Fu5TdAToUHE0nxpe+aUsL
FsP5Fgv+/vHbWfWJ0Ytz2TekKDN7y7TWxajaATw/BEma1uTj0qe5ZBSvSV91+p1vsTcTEEJeLk7B
QgQO3uVg1Lwi2ewfKEpCeB0PPPHniXJZH45ERq9eSjMGQJ69cW7564lBt2V0ZaSgT5hwT6fN6kdP
iqn5UZReGj2KktPMAB/cV43Hbu4DenKcROukmpAQhCzj808UNJGzm9pzXjitfnv5ZKDPkIuMaBYu
73e+LYyxXJNSih3K+RjIgsPq8RLTsA8xT5j3v8ZHPpjZO2QZPRO151cVF7UED8lnFq3EUDQuvcGz
M4nSgvio0ac/1szq+smnaLSrA3wndtvgTOstUCI/YWjNBpnGGflRO6m37xMmKzvtLA92qhvVtCvz
mhFOvr0ZrZ/t4YtuwPqfv+p0/RDEInn/7GqR7BM7UfIuBW0ZiLjNfG5rPIX5tnBovIwSAZmzTP1X
MIUBDrJM0/FvVP2G57vqn+XFN6X9nEtbH25Zpv5d5HSI87WCx8QDQakSYwi9V8U92CABrK0HF7dy
yuaMW6skX9VZF8BfUPrwBVdPw3BaXsxhE9KNSnwu3J5Bt+Ccb108guigsmyUnm5pPP+zoZ2Jp/6Z
2GhIGb+lGFwex+p65qFAQTBkzicA/dKNzXqPtN1DnXNpA2UGLXBZ0fP09J/CnZgvW8sM6XpwYdjk
0EeCsWLmJF/wLvcloQiZJ0wW0Y8nlGUisa/gWvxU5kJ6EpbFietWAA1mThjJyhWjubx73CvitiNg
9kAuBjMjD063bUE64oewd6nV51CkOIgXhDsDnucy1khxdeRfW2rFisqxNt1TO/vaAy7chkjoWycN
B0a0VWbfV+GHSMqTaWBxODClAKXLTSiqUxhXKxEj00T++Hx7y6opvpmkn0DN7po78RxlCaZrWiGB
UJKApLHjx2dUQCn3NbcO26rXMdDakvaxCZ9NeAFq4c0JYdS668hzT0L93QfN9pxSkQh/ZNWFQAnm
b8YnfY9nAvOicBOSljjEOwTsxIguvZYsGDs9a+02hALUqCXCEPL8YkQyju/epECRn+U7CoGHn/FK
jy5qxN35YhUZ7fA5RFmPnmkwBuk3DUtlB/YWMbrLWaqJfHl5r4+PZb2N7JsAt5YRXZNqq2Jszrj9
wxU6j9kNURoFpCuS3IfK9OWfQwfl8TYoCKInZ1hFTwQFMKedTXtLE11mF4iPJUiZCPyvYqs1wP4R
Uj6fncwY8d68bFeWCVdNhey8svaZD4BjKWhVcZ6SL2Ym5WG8z37m961heX92WUsLWLxgT/0iVTRL
FETpyHWxhIlgsNV8Nqd9mpSV+LJh3fZR41tPIZSStAutF5RJiBh2e9N8x4+VGXhQSTCMZLuGUXx6
CO/VP2BifK4KuP+UwrLW5PF285GOgOLdivEvzLYT38yD6iQu9relk51XES5DyOjLmR8d+HRbK5dd
2CdVVJuSATS+S9/feyB4j2OuK25eQEIv19FU/87fwPy4U98NuNKfb1Jd8yYKBfxu5Y3NVzr7LLNq
itTtY1wMPGIcBjVrK5MTE1aDILgltZtDaqBNCdz1yka4VYa+g8tt4R7aOgJSDq5IKz+YSvUvjQTP
veR8imBd9W1OCgx8zuf6Ty5xd2NbTupSvqXZLZ3yrzxRPm/Vo9Rrw2S4HwnPMO9PIuDK69PasFm4
AwbbBrV9PdieaCUKWn0AogkSF5y2oq2qDiVBRVIhlpEd2annIM2qzLcs62CIxi/tcFLRpbeLWCIk
hog43wTlajTZmMa/OHz/NXmKv/sYnmPbdXhKZHYi2r7Li6wmBZlge/VI0nPpAwu7XRDeGndC4gp8
yfTgMJ47t74iPy/ZNXT2xwlDiCZ1hiW59mwjHyl+fIQmDZISk59JkVv5BzcWW1SJLpNgEDjhRPJf
HS0BuDuMVIJGldblTxHMuzcuc1NmomzF26JGuLH7qZzoVdlC5triMC15BRu9BlhlWHtbwzKUY+3N
aXbeebtJfd88jAcfZdLb8W29pJHxipX/VuLi7sZMSMb5NML+J/Q1qhhoXvR9X31jFDZkVnANw6Xw
yt4DDXpSApUbzHfMF/mtIv+PIrLLPeCkS6eP12f8zlLFYuddQUcAoMaPV3o62+gXddLaFvWuBSKk
7DlaUngB2YvS733cI4lXtQ2SbRfeZk3eGsZItpyPCFZrpDuiKgA16PP03ewCZQsTlzpuLfUDW3u3
J1OA5oeDJ+UUVY/UD28d+zk4m9zPpcxffgmdZX5ylhaLaC9MH3OT2syBUaniM7t1w2tcufS/0ZFD
X79HV0VqCaHPqm+VbiWeFzobWTTPQGUm2sk1tR2SrOGsESl+coY66cG0i1UjYM86AdDOYLUxKWyM
4Tyw6ZFedlIIEchcOBtZ5xdlEZDtnayOtODC4fW1yeWBVv3sLQKxJTWzL/HIUE7XrvppsVVYDmf0
Z9VoSczJo+i5t3X5uH2sTxa3vQkxhO4SFr6LixERgZt3u89vIwJH4QS0LXI/krw29y7FjJ/HaWFn
ycz5G/9NUiO3brnIk3xSFVJlkyAhFMMY/YP0OHWagjAbG+dhNwNU+KmC1jb4v2Of8mhITWYteb16
fy8g5WU+6j6aU4xdFDMJEIF4TOOadJq6iSJTb4TpPMOARZuDD7N57+DtcHuHUSc8rE52RrfIYeF8
YCFmcR+DoiVS8gxaCO0kq266xPMt976dVj6gMp8HHhbyFiZPAKCBlwj2YDYe72MYqBpQwaLU78Z4
3YZwtZ+SwqhoVI1i6Wk4vLlevYdzpGwYyd0KV2sM/ANCooB5UbeeBpfBtWdeWlS+DkfGxrJIrgzt
1hc1tvkQ8nGdnCMy8rtwqB0HaX2v8nHQ3OuC2bNXw8UByBxEjjxGHRrywc536bwdfzvNc1OKq/uD
F8qyVKXzYudEZYQoYqA1grjdtPUDotF2O+PAqPDNk0PbO53srabN1tqeeKw6JdAVgPd25/XPDH3R
YMtMOVtrOFNK2/LL3LcoVrmbsoLbD3vJ3+TzKT76WlINOgQmiYbUvREDi0aEx30tERH4IQxVPszQ
6Z5UBDH3TAIwRwTDcwSVVURCFlaYT/FBK1EFKuv+NzSODuoyb/DZCPy28rWXVuzymtXiQFiFcnjk
IhB30KpHq7C8xtaA1IZMESE0zUtpM9miGPyeXxrFavQ4LGXoXpWJT9lXV/xRsn/Cr8K+Y/7EJcJ3
Gi159mWp1V3itvkDj8i3vRWGkMB/NqaLbCtDWHXYMWf6OsrgBc2aeygdxm6EKQnmk8DdUPetxo33
kfEJpBOKvj/BN+LP8DMwELuFi/hw262P5C5r1w2OtSsDxWi1r/lSzDxKtpyW5yhBLqs9R/dd4nFX
qEDFAwdaUR4o1vA0mrS2trixfKbDEHWyPWGVWtoL2TiAWBM+P9yORyQhREcVbr8P1Tx6LFe6qO+U
K2fzhG0CsleFBexGoyILQDF+SGKSw0MENhz/0D399ZmVtiz3VRznP9tQbPdXCj9SmJ1+70Pa5efc
AQ8nXygk53qxXiH5dB5mDQSngtyNSzNTF9h0qiqL0BTRoLzOdqC8qzLBQya1Wxa1t5CM+AaiX0S6
FSRQ+C2A8oh1kmwI5xsetHvxzk+zWkyKCkDSzpv32Ro5yd5LlHmQCbUrhPLQsn5CKqG0SEgxZGJX
dxqSNELYcJ0uNkITxOaqg1kmeEonkEos77dx8LzxFYL1iZtwEzEX8205TSyB34vdBSokuldgRUMZ
N81GCGBZ11vCwYfcED3NhwgClKpRvi/g9PuEKOL7MfjKDiUV9uNUoyTntJSZ3leYPo9Ckkx88ocH
Js5C8wJqpdUh5tGTGWWqLH3gn1Am6NF5Vcb87ALRkXKY+xQrK6puIARQrsCx+LgohGqPI2uyIKLP
BvBCvx9FfL5SPGihIozMldEwNtEK2w7qfJsLgVrPUrJloTSqHFLvTRuCw6oczG2Eye+gRCvKHmaT
jXNTAS3W03/gGF/TYXcdh1M7DHo8BreAxGFqjIqzRVzCQh91rAKOFOc/GlZGnp49ozC4PxEOXqYQ
V1N/HCh23L5aW1TL4vKz+GyxpdQclxqNge+xvRX8UxIQhuvymooO54zrd8+BHLqkV1suMb3rjl3J
IxVvSyWbhcFkod2fqIqF+CpHLNnqI7kD6phSQp4152HzK/7FmOYVKaziFCF5KD8bagj2P/CChBTg
q8gai32o2iYPoCnwIM3DXp5MK3rPd4Mnrq9ioqmTtgZl+BMhdKRG9goUKvcGwybbwPHweGKP/5mn
bLphQvj4WDF/Ox4r1KV9T/sLK0kBVrowcSvrfxlx/CD3u6P+ZSeD4V5yRo6xaurkncZdd0R/W4NC
Z77MOiuhMc0qMS4cOkDIaZy+7jXbLDCrf9jyMHDesN+wyAECc+ibBmjkDo+xHzJMY1oYdHAVDsP2
w20rEnEXO5yt1zJeB5n6mGdB7K4WTU81BP0iUEICx0yDg1IVogEP1tm2bIS1dKW5R1zkMAcCXFX3
eFo+AAD0oBH8p6nSiDzh7iOTh++lLiPc9XPpH3bh8hoeFfXZgrEHWm4pj3XDjJncnh6btdnrGj1S
pEMgLpLB+TnvobfUvLpJVp5AnZrfoYsDqfLY4JAu0i0dMvjE7qejBhI0enUi3TLyBKt1sY2boibZ
rNQ2a8X3PGXcagWBGWepservrOreByKFXT69tjVuN2ZrudmUf0OI9zDqkiSv7McqpZvkpQxMXqki
ZLoNGnYVhGzIUJvt3roVWIqKtPIbmyokn1N9heofIXVpF9HQo6WbOfUgNgypFbJMKyZ4OUqEeMzA
cXXlpX1reJoN3u6fRgHipLGqeAhwMRKR6SkekqWavP84lvfGtOEU2qKhpDWFOUCYxSUFsWsgxb/6
8sh0tzCHM/gMgpdoEsGhVZ4LoVMFTgxZ2SJ5oeE+5NY+q/zYpLLh2N7/ig7TTKAhASuOIckPasJZ
7mJoLnfRT1BZVGANNp5NelKqGvXnAl2cTHtfya/W9lCokYl0L8rjxbHRN3LeKSyD2bWs8lWZa/uW
RU/NoNh3skqeLteM+BgohwUbJdLpHbzf+xgrTtCgOaRS8u9xcD4ZdMBuqmzbJcaUeQ53jxCuJ3cb
3U22wRWvOboCnjZCO2Qopgi1wyfX2HKkEH1KQNrOJOsaY8lg6Oz4bhh2qUOzuQ2RtKbDh85kgmdI
2L7qbbmWNo6Ycsvq4W8DidUI3yl96pKhWoGnNj1qGeDilR3OmD401OvPXbXRPpWrlElkNNI6aXjS
ksXi6+o7Spu+LzZv5/KAYjQoAQ8Bshk8bJSs/Ia/0y6A5/ptq1Inq3QMK1u4HgQ9bPgo1M2IWxSx
o2O7vNAqbxPh1F3NmIH8dAtaxQkGAuAgtlG0qUXScrUqLGS4fkxPMzbXAXiItKg6/mQ1rFR8LQEG
FwYRXiz+/EXEmm1BvvEMWBNqukVQ/EI40iob1kUIQNADwBDBdqjl4eFYCPMGABkxeQwOx6eDPItg
zCxkieSOo4e7SBD+PgfxaPhbADc+gfKDyZf0B10aFSIngHE3jLBCe5C7UWCol0Xk5BJinOS+1ZFG
N1YPy0918Kabq7Xy73PiH+GmErQMXpp7kF/ygepDnUJ5psckrZo2xU/0/OeJrXWvVFYKkzTE1k8f
+Vt3fVjcPVKnf/mCZ1/+ZyoRI+9Ryz4bSKEhL8hKdj9JIQGgWKTODVMHYyGwUdYX/m+/U9EpUzJj
XhqA0+31MQvp52qMW89x8a8vh3TPgaN81R8+kXFGAB4vTaA//Dk7nArsAh0pib5tOQCsgypdbR/n
qrxDts5ilx/KbXCR1LwjXQIYmKq8yIMENwMOy4eDy0EdQZK2r8GbLqP1eS7irLz7ZvV5d2KkgJQO
xx6sEK69PRV2lfW6q41KcrtIVm+Z2OXPNhFHOrOpM1fxQuwcPmokapUMPmHU7sp/Oews/nvREAAv
tKdYa2G4Wc3f5Kt+26B4K7BMQIQUnPyEhfIaXmNOnii6uISeNFaCckbuJJzzvr5fdOj/q0WX04vJ
eSdjH1I75YNPP6+AYna817Kri/bRPlolFdvM7mSUQhU1UJA2JlmEgtSZSUesEIpumDV8BDLq6v8x
gb/fPj6y97X7dO7vA9fzol+IO8azaXfQhBAlgFCB049FYLfPQdMJjdUwH/cIbkc6XhvnivVJ40NA
Wzs4PHQmj9DE4B6hAHZw70avVMXUDC9y8seS/w4QjqA5VjvaGQ/kQBmAp75vsXRz8cB+TFsv/DDD
ukgxj3O/VPeoha3etScpoaENWhegqrBpIB7VQPXPNt6qHe7xnCMUPzMIXj+GlFOG0YM2hJBa0Uit
z2GcBSY271BJZGTp9BVZ+8A3eNIkZlUvXArG3eKA7iMxixSrqDmEq/IoPk5iFLVi2h4XZPj2CmhO
jN7s0vLQPnvhgbEggFHsEYl97Q6BoePWcu+A+aeDcq5MMppZDjlPQUrLEeyKGPR4XOvr//lZsUNd
+YqNzCvqDmyIGiHAEF8s2HPqwwfJYHRpNwnLWh0w7iJo2KWvieBy5yz0pXBwUSUjxmjggLw5GwDE
DJnde/7oo5YwPDe6RzE9B6Up6b05ef2VSpEDHhgZ4w4hzJ3sJYrXlXuadKRaID1WWM4+EKbJDxcF
8sV/icYaYNsMNZPpZLnpORHsnioZ5X3VG+eOic0qwmX8MiJo/sB3F4/ncYhaBX5dVbCyFHZG61PI
Kb0EmNU8GVVuM+SDbPYlzinNz2Y1vupun61ovhMwuj3xi4TErW9PhHuFt9c1KgTaOTcb/S9l/Mhl
b7J3w+MtGzHYiLWsQGpTx+pkPLCAyHglAiLedNjW2y/3pYMprH+YHmgFG9u0hkVpO7YPYPsROt2J
WINXefjFm2ODkwy058U0eHi+cRSNg6QOAkR/lYFWc3iZXWjHG8/JpHMUNHwb26Qw1aPeSK3WWU8s
Lw/4HM1x62BThs6N6yy+smdlGnHJo0AuVHHz/SW64/CZtyGlYKm4aeQXBNK1xTsMUT2hkE4M0p60
17D07EhpaaAP3HG0T9chvGknlzhckeaV8ySNRmiWvu75gtY5W68YZR70eVk3YVot7z+IjJlqyU2f
vMK992GSgaknHbMzKdSPg6g9mbLNPA45V2cRie4ZC6kGatZLIYIurlIfIKkS20JKVGz96HE4ksrm
ffbYlyfjaBXtCz01POCsHPjGq9OdjodKfYHSBAqJvklbqxVfUoENISOh4V5sj4OvjBPZyE+VdvEu
T2/zP8A9V+7JImFg9QBNKAZQelPW4qWbd2etagZmOxg+vfkXPMN33Jv4WJDSF8H9tQr+p01l/2q8
kUQrkfIzW90dRfsktTkHErEMNlK4pq8+n/uqjehCFv5t6qw8KKFTK2XbijhkY4UDWGK4JPectFjJ
lF+E+GKyGS0+YcpwlxRtuh53ylYVY69ecMSfEqtjKVEykyu4H4nPX0Upn4Y7b/BGs/CwD1hJFtkG
X2v5YiJenZjOLXzi9xIBcrrjKIX4h4tqgRJ4yUAM3NoIHjjlMznlnwq6xIUPoF/w91YM8IQZHWI5
UAWI4u6woz/EuK6p4qD1F1Ig060TNnZlY1FUiigRoTzjTJZeiRCyhPYiW/WJSnARgcRIIylsLFcG
V1DJoO2weqgy0L327sHYo5YAPNToONiEYOR9axyccf2yE2L7RPJUTA6fAvV9qQqYl/mTOSO7Hgzi
V2MVGBsFIYPwDPygewaoUij7R0iLcUpZAM3g00sAtDKlRqBJ2hJhlSHZdluCB7FPiJm249E8yVlK
nR8NaGagxall6K+2CVXv7zYAmETfTUbVCWtqBWMRlgvbeazw7qeW4QLm9mIXZKkPxmF3wYfEqltS
M3l+Lsd4V6zN6SSrCJ2WIAR5Nkecs4ayhQZUInce+9poDO9waPgp/6MDUIoGeHHNlceSZtIdFM2L
pGkDhSaSMOSfagqVq1Vou27D6MKwnGFrCzxA2oTRa/x6Nym6uaeQR3rC6NVDrBOYo/3cyg3o5yrt
i0TZ60+ITcPVR4fG3Ez67/VbI4M/LDpdjyOnYSfaETqMGNkVxYbQRH+9q1tYlKGLmzCHii31HpEU
F09ZXE+uiaU2D+GDS4VXos0KdhlB3yakQ2kQ24kMdniqEVv7qkdo9Cr1+1g6FwL5rdWdFYo+1oUF
1iWPkMK7S9ZxxsTJu/fFyvupYRtPNQ/cQBVlprqpn/TmrymQS8tsNI38awnnrB+ap21nGiTWQsnZ
EakOnnZDuv6QRljHme9OqxnXxkx6w/VWjqj9vCSCDlHRQxA+OwVoFJ5gizWU7CLkbPHESwO4o1/5
7mEsytjTSKx9u4/i6fJtMWP+3SpHkts3c68+X2nLp81kXIofXEY/Lq/TMjcQ5P2psNE0CrXJzKJC
sBnphaTJk8aZbvyHXNnCWA1bxkviJUm8cAVrsi7yYh88rGpQvSYdGLzNUrgiT75yxS5Qbf6Vq/9P
11F/bQWFUzqjsA3mFQN/7lev++ykE0alkGjatx9Y7Ju3Q5Y29c3rifcJJ/z12rm8II2LczZfMvV/
ykUeOrIhssbpClndh1kvpcyfHURTbovEj3eVbW2ZMibZdzcgDTIM9OfQYfvinFfWE2yko5Bckv5N
p9cZjucYpBMZwBzr6bb4iZsNBBle8WmkKqoaVIjOPB7kbIFhPLqwyZW3jZDdoXGyg02JKIOFkS+4
RMS6XtluDkjPjsI9uV0ktRegtj0eRZf0neizLmNOlcMHFpafswf8R5Ep2+fECjsBX83uz8j8xZbS
+nrwD3YxIzVH1jM1G6l41p4WJYCTUqOGByL+UPE2nGkzs5OoLDanbElA4QmgXHflOI0v3YhxWmPV
hDOtD2kx3KpTq109nzphfozc8RRdmRsg60XvTs68OlMWWuEk4cEtCgrE3dXfcmrJSZtNK4Qkcsuy
W+QmtdxpGQgvopuAOz5DAa2ISu917117CZBqKqc4odwDpNZDy79kIMsddZgykKs6s5o9Wjhq9/8h
g4PhL+hJoUBUxl4Uao5xjp6lwlnsrQXIOH2MrWSvOS/4DTZc7yPov3J2Sap+VZsaP4n2M4HyRIKv
Qv9UXdcIe78wsuK7ruHroK4lqh7kQDHW5l8EZvi0Amw/51+cdG6b4F6wVkZ4nmXMXNd5MFtYmDJl
8vb96k8rssCevJHWlx55KPBP9tR4fOHcclAz8j1Y24+hFNQeHCs6rz3wwjWW5TrFEffuoOggeaZ/
Q2CcXpZauEOTF6BiDtkAVWlYOsYp5NmdbHoEEP3hQ1VMkNzk+SMBSnhWOKXqpPEGhlCwhofZsm5+
+EOuDwFofhPU7rVlP7viqoQd1yPA6ERbkhW5d2qk2QUCnD2mTdQb8QiCQxGQn0UqN7qjS8OShC+J
t1AKKfcEKRATgotHpfnwQodo0eIhFiLSmbs55i1uvo+u9yRhCuUiqj2CKuMOUyAbTqc5QxIlF04+
pOzIfZ8BC9GD1sGZYltxI++9kd0kMZ/FBafIaEFgg0HpOhKlZJACCdtEb31RirRWqMDPz0QXo4A+
1oI0y167gL93V9WSXWmdHK4ZN6y2nihT8k7owLEJTZaRvzM+Ei3KRpHHZr13xkC6I6FLqESzD3Sk
U4C+SLyGLvO3tVNkfJ8l2O1fQerH2Ew2u1Tbz9Yu0fNxQHb3zTsKpZwVg6VnVJ98PU13OfpOSZWX
HJiHVuhKp5T1JBUMr8vtK9LPDQTqlAdEYkouEry56btrh2GV/1WQzrrLoTCPRv1In6eGhCWUUrSH
Mb5Zw+MiLPh6HlBKxy/WeURQMSE24wJtOAe4uu96KsWKNs11prL3LPL9ssLp2cV9cp2J3H3hD6Ks
h10rbyvpVDhZ7QcQw43Cug8cNHQYqY6MqTvem6ILThjmJJ/lCyze49ay7TKXQVWi6IU9vtuU5BAT
eIIMkk0bx3fD6GYhUgeLvb5phRNHEjiqHaNRt+fcTuDR8Rqw/cpzM7+ART5QZ9u/CdKibSNeHb7c
l9HZdOnzcReNauMaF+hVpHBOnUwwY3GO04OwZvTIGIIgbK4+1b5jIRLDODjJkOVloaKlk/s4qQ9R
peDCrhjfapxXS9d1aZPcmEpgEUZl00e660zCvJBW6RVicZWSU85TLjnahZxHl26sSiq+bY5TA1ah
q2jEPKTx64dmJaxlMXc3uBJ3Wnf4U+pxTN2ecHIkiCJMYtIO4WDX8vnWjVx9gB9e6TCbhnjM47rZ
tEKF0J1oL/LuOurdGnkU/8JCUejRdIoiOsFJQAE9oKLtcRWJr8UP8PUUSvBAe+zG2bcpQXcEn2PA
MayLbpwuFJdxewQAjBi3cKc5oEgkIDFZNbxz2PMHS6YhGvtYWFtK88M//EmFW3PlZeuWo1WTX+YI
TCUuxgXcjSmEfbefgndYOelGiYOK0fAmRf6DrQSYD0Ir9vTi0L1PpMqtI66TFd0bR9HF6Y+Y1bdK
ZtsOiBbNlns29Lb6KVN0I9wwqGD7Lmdr0Y9EbVqDKqYeNLQ1wFYUjHwxP0MHScbbUWNDs5J8tIeX
9FaD9koNdg/JnySpciW1ZFrhRMy5QOOCrTTKFH/7Nju3KI0KZ+kwd2G68xmfn8Ci0Vp0nF7LUwx5
7eYTGboOd63gMXgiDqEYMaVANNvYEprUJStIj+gG7YUoPO9v7lVwbeBAVhxNkgFomwOxN7Xh0Ej8
2TWk1NWm6PcPe01kr5ZCkPyB7/n0WMb+7uGLYSKRMOQobJdULms6z3WvCzvdHPmPkh5qfG8KeMOs
oMnlb5SJUmnlKm8MBFslF9A5Qzvk9Y9ji03Ai4vnkV8C9UU1K5OwBsdPum4BDY1ur7YlgsdgsNEM
rPqRQeRzzQRZV/aMkmcO+/PZD38+UYCjtWpmmHB72xRWXgWBVXmZEOUa4DOnDBRQYQ74OLoB8zID
kjG5Ov59+TGsYkqTp6VbhwklhEPe9D6q5tSrrJNue+XXp74/ShXpgGiTaW9pYQ/vlCcBKoyBWh7a
kqYYmXV4i+6G3JpefWaDHhnhOl6X6BxZ3BM0Abzl26A5iesnsZ1kZsRCA7EKPOijFa8C0HOIe7Lw
eEE78Ifv0QQkYl1K8NHXjROVMJPlIFzVZpZX7unkQlVrc7iienz1u9Ih3hE7ma/wjVhGfBRJrp+e
fpyOYT3b0C43t38zXxzwr098A6bGNhcts9JtDXEnA3kyAw8d5FrwglfWK+RbGaTwIGMm5BXfG1gl
s1vxHwDhSQh01+yRpdJOOchvpalsOy/llFc97AtWAJ5QV2jItj3hY0J6tguf4vrAxgT4HfBeZCl0
UCO1dtwK8JgE7bVvYKqm6Fu+gzjltMDx0nTvxQLTVyGdxUvcSuCxneyBC+Go3eeDYrjMK8rl1KKv
1CsrJ5vLJ7QqDTggefECpgwIZbAjJKgn2wl62OiLZZDm2Mr7K00Z8Ns/bQK8GNSFR+wMhn7RReGr
zHJ+0c2l6rRTTQO2qLB5uN1t1e6rq2vFmtzNlknMfJs/Je36E6gzHiFxftrbMWAnhiuH5cZzm6w5
/Q1nHtuCeYmi++UiVPxRm507oGKJf2gaQuwfkBwUyDcaTE4fdHG3WyKrgmJYfYuYhKW26XEW0PuH
/14wA5f9O9fGQ7/uFZ+MT7yRO2nTHAO0npu17HHcHkEbrReuzs5g2MAWUwRoACbeRs28JGXOcW5s
ZEt/FklQbKVxdDM/RVWHlc6Ql3VurKjJNnafYx2iCsHXHI275wzKJrzrjmQv4Fp5s0uaSKT7usQ/
isSRiKacVKUAQMC28qnFdg8ac7UGPe4kbCpkq047m5MPBaH6QD5+M2Kds9O2yiR6g2+1s95HW47h
gajGyTTlrrApuqtH+nszfbeRmfiCxcLvhIvnYp3cPeysox0fuSLeUIgCT5tB8DVNb+L+8jReb9ef
q5qeiCd0bQNinHoX8cjdwCajKyTlCB9LWjwGhHdD4nIeqKqlAXHGQNKvCnh9otU+XqgvLMnhY/Ry
aTpUJdvvk1a2YcNJTZc6HmkUnHjqmgKfqVWKnwuXXnEV/T6PlBQpO5oxzheOkFWUOZsNXAF4lCO7
+tuXRtCmq/z5VcMXxVZqxdXmDg4G3twawcLSDYExoucg/xRdSkKNbZqD4r3Diqm9dWfyo2YE3jJc
4Kp8LIDMUg2nJi876ta4ACoerp04tFxXbdgRtvRkplt/1Fcg3c9XMEOCxx3TR+/hOqoizrFLeESe
mBu4/TeXcrq4+Xrk1uSzg6cfGufjzWr6k8xayGrf3pU2M1FPCoOtdSWoBQUhG/7ORhdU1sGgELZY
eqymFPnAO4Zv/jwcP4HK++jSbBqV/5Fpuy5EqD5QZum4dHl/sAICs0qnok4KNPvOr+quYje2Q5ut
6UguhUY44Al/fuBptEnagaziWUN/AJuezgv8XRynBXn/Rvsx4XNEz/7HKsRPvkjy+OicVcvjr6h1
8B+JfmTc1IaZU18Lx8NJuo8V6endQWdvOW+bB8dphEqOrAuRixBKjlMga1VGzgIndt/F6zfp6UgV
Xha8sCHnCQjl61pPhKmpYvgk/LzidOK8J8yF+KMn1r8WhLGqTlySadd+QCAS06hAO578BNWkmHI3
yliorG9owVQPR4VAxfk8fcyI7WywwVd7sdotSqY9CySPPa3rvQlDIq9+luChDfKU24BmbAVPt501
6GvLmYz0a+U3btiG547C4WAwv5ay4hwEtsUjrckt5REDFudmrjsqVQf0/RtkhvODx0RUvZgGtBuH
0mES0LtRMy6UuDKAkh4me5J+TS69ps4G4c0jU8ETkr491rtOiY6rxikoBhxVBfizR09rwBlSnjGe
xYNgTQOrjjIQzbMJQnEN+af4caqzd5Dc2wyhafF3VZFGXU2RE7gziWxC1FoYYe+zJ7ReTX33ZTPj
jXBog/WUl4cC5QRNZAQ+tiX7oJs7sCsEW5FD9zMUYmDXS7M0CM/YvWwrjOPGf3SgnMp6npqBJnAm
twtI/jCxGvfMxsnp4R0gcKTf3RBcKwKZDDH4XcFlgNenaef7RgzlUtnplGcNi61QY839gTkevEqP
Q8+80g48fzA6+7zsz4vX5wiAiqy66Biq6fhQynWmTISozG/yP/Q08GvLzuf+y2bqCqjcl6o9k+9z
OLYUVyt9Sxq5CcDrBPw/tSOLuFYkS95byjHQcv5hDQCT6Fbe8A8fKVei7VnhFSG0koB1eB5ac9Te
cxyuNO08vlMcLAmB92kvAHlvZ7Ii7Tz0s3SVsTTkbu41uQr84asac+1xe8O0nGdGcHZOlbDWIl5K
JjgNNnK89les+FUufJr06kJJg4CYU2lKR1af1G6e/Qa+R31E0AscadnUc8buK/TCo83toIwT8lMk
lYdnLvlaIj3c4dcKN/u0HlX/SobAt9U3kaqFpyd51EL0FSJzrphvDnMdArQIzjT6qNdWeo5ISvwF
Phtk2q95vDmqvph0CdyZmWSQ52F4Y2iZi1NYXAw54LgfWs6W0ky6mosXpSY72ZRmEcToa+Ss6Fco
YOTGAcunWyE7fevYp12Ki+D3pZWC/dknkySKWgKXUeb18wi6i12IyVdKYr8ey4iVyIcmdhi4Jt4p
mWE8lFVJixo7J3kW1Q9ZHOnzN3e1wONmt8srSkLuXsQxhIQHVLMC9GO8syW6i3JMHr1+fkcgqNrX
Ah5kLCCj/LWBixRw2JhtLF+VyN7z0kd44zXcsPiZyRKW+k2RzfP1eFCQr4dGujpRKrguT/3RqTfJ
TGwLWDeMBAiFyByplzqMlkT3vug74GbU6XojMn+pxlJPmB/qXEUKiIisn+qypfhTz/Y02cY7PNj9
XFm2rDfftEec19HIqBn4VXJqb6DJk2oEVjTRD134znInG11537jcydqhhZkq0u5DBsPR4mcyfXxD
RIyaK94h9Togy89Lc4xJZS5XhOnvHPHRicRU1Y6jriSyewyqZ+09rA9OyJ2oOPwuAhf6FO7c46RV
2vcpOJo8rCLunHa4tdm7qhHxjxIz9FZqfliWQoqYyyZcjxaexbQq8sQKkcqpAbbXxL3NodRpDWU5
QoaVD+7QzaBPS87USFGqlHn9q6OIpiUo45zxc4xSX61L27QnO/Zh+FRPxB/zqW+WfK68cyib350W
7ElBtt3e7yBMMn+OYF19hC4hh0qskci9d4NlMkdq+erPmbx46NyXs25913dknD5dW0ovV4MpUiXI
nSci7eHudMqGNK6CoTj6VhP4zXuRdwp374KwQmqzdmScFKeRB4qWAbMlpGhT2Qj0gbZp0JSFkIDA
4JmV6VMMPZxvibXt0pELv3fF/IWyXH3o9HUl2mt+ICdZFfW3XQai7NFPlk3BssdN6b78aiPP1/NG
0HVio0tjMwqNZQibYyfPPlUiNff9ewmMU2rgYjEoJ2OzFZHK4cWK7Y+Xeat70tCgd/zQFSEUADze
g/86ybu2KcJCm2iCdKP157xifimLXYawQ5CKtaRK60VeXQdpCfbLTImBurjn1LBlFA3K1Z3PMr0N
6RY8RQ7KGpgnYotEBXQqws42PEFG7HjpMEZvFOTUwOa0TZJbuE6lRaqARfQzNVZIJtq45GQHc9Jj
fvx4723/nYrpU4py1xvk5mJiv0FXeyYTOz/qdsGNU1ipMkxx9udl02GPcg2MDpqxGm2llJzDVYx3
rCtByFzxIr+cmTfNCmyNV4ruub7o63LHeAig6Gjm9hszFxR1EZzx1vDlAUWEza+Nq6tjN6DunM/n
xTyLMtYoFHidlt67ee4jYAjmTwmgereWC719vpDENbxSQTC7DgvVdo7oqOtVlaYcpaKGUfFaRJpC
bxGQIsW/tkA1ccKqgJGCzUElmaAKCKvl0g3/4hIN+2szlp0COjRxJwcMPs6qfMMvctuDrHjHqYRD
FJbfVLNcVQQUv4tMvBo+uNkO6ZauaHVdK0hfdHcrnomTpBNHK+b2P5s8tw3zALWKrQ4lclltR+6z
YcZO+KchEnIlgzzx26bg2mVdha8ozl5SYdKuDdAFOJSU0NNZrH0wCdQEpKR5MxsEA4bBNZWTMfqN
HV6qJV1YdOWLiMjJqXGbN+aGVfc4JMWB0hRNqDAqLizkafZvZIYJHFH6uUiEtUmDuJSnGO4NlM/0
CAHamntJRQtDV1biSoHEjqCuB3l0rvVqW3tBDRqo6cxFHeX0bKo1gDbF7Q1qpKpDZyqNj2fN14/p
OmVAWIoYi6v1rJtJoDlPcpm2Ml/1eKZ3s0bihPuL0JtbyejZm31O4taJ6/j+qKyUQu7i2FyurOEf
DXyycYIFs5WWjlOJXx//T5QWnJpSDLsgBhWJEdcYYFp/ZQL7TLm4f35yZGswz0TxCNMyvgAWugnB
UY1D1U/qW93UeqDU4BerfhhnExQDCpqBo96kJv0E0en9ujPCPQ8A7j1AxFZ35lOaUaJr0V3mt84j
+l1isi+NfjhBNBpLc2OhS28q6hxBUp1qqa7DL7TEQTNhalCCQwOk4PMUf6cXUgZIQB07dWFn8evY
kJEzR2yMzHeI0X++/QOQsOkj+UvQw/Ry6VR5CMy2i40Qtpfabh0hP9DfOwTx1OoMChrERspVpr7e
0vdzgirbrADQX/cR8Q4wpGAqshqXFOvQwmcdQLICMe3CYnohjHwM1EuKi+0O/ms/vLuSc3J/SZi7
pBNW7H5vlDBeQgDq7nVxYkXoHmK5wzySAoGJHTKUjVHfF98UnNjASQ3VWHx3c7JrR7pxQXgs90WV
gU/LckbuONQu3OOYZt3MHUwNwrEgOlVmvvxDHnuDVjvkJlo1cYXEWnzmaHfMZa80aKYHpAoKpWNX
39h/lGhTutCAnTPAE6yMeww9+Pn3zntCQ3TW90Yo5bI8tunRAOUGPBT4Kv0kR+mQNKBdBGjheY19
z875Z0TmE2O3ncVKhw2tuFMFqxptva8v+WqodIwbuSpc36YA7I3fsz0vC+WDlFBo3yfZ1WLbnTnH
EMPurkw6/JWKWD1H8Jv4vTBHfayYeI4zBobPUguiHVNk4an+qiTM7obdkW729eaol9K9cUF6/PmS
FL9WIOOtyK5W2g/0HAndBk6ZfaZjVHPEJ7CQNDMKmIjdwIjheuuFdDjLavhssFq0J9/EsvEnDYYB
hLFjAD1/nvHuLxd57xZ0zbfYKxgEp1QzuZrYpsKzIJWujiIXIXJ1oWgHyoogLGeLWeyP5/delh7e
reHEPd1ccOifLsz7DJ8NHQnIhszKHIOQGfiilbpyzdYyH3ierMewurEBurHVlebR9K7SrTrDM8H0
IrpIM7qcQkr7jJ8FFmHr+mtVXxOe0u7FFRWstCl4cUxMlgU6MwBn+6VG2xdql06nBWlBPPBD9y53
jtpQOPhazFTg0UE4V4ceGMJjzqL2zk3l3VXYVo7OPBde1fp3XSG/ScuLuRUy++y6WhBzj/C5b8G8
e0U8wwlgsvo5jcq69I6LGaLH2mbI22bpix9gmOf8Gvdnd+4Kr8zSL7K8760s0fYVBhMSzfELvdIf
OqJksmOrq8R0Bd7B9xST+Z761gZxyqivm1dORfnU9OVHaF8Fj0UE1g0khQ6YZ4hV4nyn5L+XgH7d
hK1DnG+164Oxt4LZgip9ubB9kDw+SZXeiCVO+XJKzWEA4hisRGjQ5pdM7bUluuBLngOPfusNTW4L
FLC8ahbK9+Y6rhkEp8O5n4bpLCFV77ej/mHPjPHDHN642//9Hod7rd94q7ow2/AVWGg2HKacwDgH
nx5bun7bkOvvM1M4l7b5MhAsvvdFaDUv3CRO5WSjWI9ZLn30kyZLdAZmRrLJbSczat0J8dMf10oO
XPlWCBTiwCiH86J+Hgyl6Pzi0EDZA3M0jBJM/dXARrWX3bBob6yCwmTmJKExe+ydtturcb7qHCmZ
4z2NK4BWWoB22uxjVKXKHc7xSOJ20aYbuecf3OfVvrmhGGgq1eoDPCKIUgovqeTgL+uWvVI8/wiH
4wtGglFSOBf3eSxDrTJVefk+STLwKZAGHcVaRqspNGk6AAvt+4Ivb9p/jpzhcw1VA9zWmp+Qw1ZY
z2/l4RDMxG8l2S1UNOH4mgGmwom0qlb2VCXJ5d9vk14+8O3LVKzyyNTqokZlMSUdSN06dTMFRf5F
K9lqD0dNInsdQfb6/hrtSC91jn4nSc6kqjJVxZMAwRlm83S85pypQRB5HwZBh+5bgqt6PYHc8qSl
nKI9s3F5NGm5VLctX+M1L7ZBevNt3R4hLVzreJWRxQ7buh+aZdt4m7ctv/Az6UWLzVP+gErxbznp
2Jru250jUCxrAzdwK0v7fvGcJxwF3bf5dM9L++3esyl0XsORE9no5y3GxJSq3d5CH5uyKlc3tuca
dnCNZVHunv2j05aQsTZYtyflsJz76Hd53z7ROWDKL5zdQ33031y+WxELEYNlvz0PCAvVBk1/HzBc
AD0sxsk+A8azCE8PK32EIM+SeNjs8+P/x6b+bR7TJdMc6mGUFvjq+peYdDd2rPqW4il4rgCCI3mW
Uci7VdhtqCLZID14GW3VDF/SiCUetFaseNIYaM/ZM3Lmw3XIqhJ8+P1vFeWaEgukepxZc9TTvzLz
P8n1GTm9QO/m0qHGQSETMss9eL+nvRD9Qt8wWljpWmU5fnzfqdTaG6rq0XuAjpKQz6/QIyDUh8N1
m+v/PVI0oKd6zBmVMG6w83r6vuo5HATXZSH98gaM99NoxUfpYsTK9EatgLsjP4SOrbBmbf54+vf1
3wcqdo6iUpqiL7AG0B9Xvv0jG2/QIfJiqYWHpsgC4xyFmVGCYSh9Fu1b01D3BVjq8DSL6lrYaR1D
1eIGmcMmdBjhDVe17/mkZKd8kpBMXRxUu7DuSh2uwIrJWRweioAuGoqJgrsKVvwhz17A7aip4I+l
gXP9D23StTbeYpzA12wV5piX+lQvbehxaDH+leECrxewPC+71P1GPH3Wx4l/VLc+WcGLgF1TOfLy
t0i0Ca2KgJxA2oKE7vk85Fsd+nL2uQWAYW1CoLPOydhpjdWx+G+eOpFsYx5eqxg6YI5YefIBudzr
jrHqG0Jvp009/fE/MOLhzmhUn5IEq5Yj/4Ue6iWbl+IAT53bAqmXp3OvoMFxp2Lh3D0yvWdWU77p
DtNGB8gG6P8CT4tDNHLyPhXeKlo70nCC5ITD3nJotPW5xkMhB2hZnCRpSMHSxgQwwCEA6T+6PkRo
/DNSoeJDmiq0hO/DEeVQ3Wji1kQU5K3/8cVGHNIb7Z4HvJaiRBu54CBS+EjGqc7m7q5zSWnGTb8j
hU1LD0z9hZBu2k+LGfM3+zi0yeEDn4fY7D4FHiqjnRdCIAWXjNBNwmb4M9Fp+10cZnMl9Ig201By
+bmSd287X6kMajWvB6cD69WSBPxCL1Z5rdT3WvFwf/VVCrXd4FMDzrjbKRysG13AGXRnK4FuPDjp
YMp0/UaVGUzBURabNmn7DSVDLohBcgO57HQH6gSHc3gsI5IItYt1iVr/m8Y2IHnddyyS246vNDRL
gkZkBj6MIGZGjaclyzFZsfqcCczZ1NwRBFJOoLXB/fYx0TdJK9a1rb0UbOvpzRl49Z9MvGt5heiM
LXMm3GrY08kHnyvcgULK7GCxPyTP0wBMbwKdOCTZ4P7UGNhaKJVPsjSr+MtsikPpgSdgiAdkkEBo
jlNXByhTEqRuz39aFSPALIcctH/1pZltfKeiEdyninAAeUlOlpt4NOEW6vUwfTZkMMwU5UswmMNb
RVHS/ZdU3UzXT++v9/zatefV8Pwk1MtpAtBRT3uVVDyw87VR51in3lkO9be7HiJVzdxG3pXtzFBI
8lHkUmkTI2eEzW9VFWiPoW5fqyoUZjzV/Y8sjNsy5eIBLnP5UAqUsx8+ydnTS8USpHq1WBN7gYwA
fRaGuWYzcHD9bX9Wendov3RIZJKLRmSwXDj1kp5f/ll0un9V/0SyNxRpklVpTNEh6gIczZq6SVjz
apRXzp0KnDtkJYT0rKRYvyoPf7TsDdrPLlj7U7Nu4H+At5lKbvrYsuEaH92P75S4RTtb7yZdpcJI
lVKwwtQmWhbf3+ZB1ck6iiOZDYXchzdo1wTCfYHJvwEP2OENBdqEC7RRZKvwdj1jFZYRYTlnOSut
j5NQZ6AJa9wLikTyJYmJ25xCaTnA947gpcDizNNs7mgKp7Xci1TBe507MmYu4RRQA6x97jr5plUw
L7p6sEgl+zg6FA/JeipMh2xBV5vyX0ALDAv8yyvFpZ6IOGgX5rIKyP1XK1WvQxfBdbuYdEOakE6t
zwThJQ80XxR/43yGWag7h8NpPeC7LqtJXighzAFR848m6wUQXfqMumB/lxuQipe3F8Qo9y43I3rd
mQSpHNhez4dPacXTxuRVgn7vCZ+kupNsQOuJVd/21N36d5EfnbyvEi0x2W5aKfCcIpQ/Ri/iW8Tn
nCaIeWBUwdnX1d/Gk+AuoGota9ndolUePniNcsER8aCyLD1/GorzdYIF671nRDJBMAW1ahPx+8m/
qD/mvYAZeva7Xub5nwDj6/Z+3VaYxJ4tLClXAHKYQmkqk/oGeOG4Zn1DqP3+AOqYsK/dG7OsvbBN
ndvKsRJX68sYCFz7otLIVe14h7U35e8NC2wWQGtAn9ZORChSznZP0HbjRUqnk4aTx5B7gGVQ+Rao
wwvB8lL7prrZmHf+AbYS0Q0qjBXUYXLsWVwO5k/kKUZ5WzBk8R9d9qUYEmSyBfdRpq6g3J/HonHw
7ZbDiw5TPaed2umMy0rTwmS4v6LuoLtDDs158UG/bwjt89bTFlk78AlAuNIaD6xTo+7H3oEuKhUd
GAg4f5GO749dr6pOyjTUq33haXVkRfb2oZBzJOiUPSl5kT9w8+yDq56uvtUJv++rZ/1oAv1cql3/
fcfFs69h6oeRYCWqCblUsXSjRxNDwmoBMu7/wBIr55Zu+GH8TVjqOashGOhBGMTAiTJmsbzYGe6I
Em34yFEAZn19P53el6ehFbd65GHj0tyEvYaeCAJb6vFgRGAqPk1HdpcRZH1w7DcphYo936C1dlr+
m4dnMQmWJ49XcpAoS4iVS1eWVB/P1S0kxAXVuKdw2pz1YuCyniUj2POwPmkuhMVYtfPdabQHOHdg
w+jh6B0WPkPiNpgmA9DKnSLkEQyAx6OyqBarZTRyjRAXj06FAZtFprHTqUIssY9QLCpWX/uL3Eou
Fp8sSohiJ2hW9k4e+huBuwN8fUz1YLYkNhuk/snYYrmTyRfmXwMlBymHMMUP+EYfgvguZBNWF0Ye
KTn/A8n+yiUNiGMp9l/5v8yXxzgB292Y7fKk1xGZVrQ9tEz8QgoGd1HeQPyqButSH1sw4/f1ymHT
RmGqLUL0eDhZEqoc3OCba4dXGOx4Cf6DO2wdV5YemfqcBndeyOAC2v6/a7iJ/J/Obfp6jvpn6Uf3
a7nDYRTJdp5M6nlQwYSpw1Pg9dgvXjCAwZOAJ2+xSOzr9Ex2X9wyH/Q/71Kr9QOA+t9JJDrPMONQ
EZU0zVU28+B4d9BwPIf2ZvhrGa+UMIHQ+NOWV6Wd5WLulqH8oYeb+fq3kbPsozihCn5N6yi3eqUH
WMy0yVuU7gWrqm/Ih2luFumkWA2gnDu7Oz5ozYwTSVK0WIlOdGrT/aBQTzWmudoXkBDLNE2BZudW
bWeULhZjgS2lf2X7tD6BRNs2N9skvGOS1gH/a8Wt1apHoVnpeibJ0aRynzOENsr7JIEvDHi6QaiE
iQ/vA70MbkLAKhdWUSByChHYmWjOqkVLij2e63o38SQXuiT3BTBT/yU2wHy9UlK0aJwJV/+99bxB
X0nOhBfQMQ2Oc6OO2vPwvr8oy2h57kN+XPf64aU1FcNmqqO7438dgYOkFjvnXguUtnILRbjM9NMR
o5z/iRd4b2rwKV+NdH4HW6A3RLy2kWFMgIb5mgBFgGKXF4aoMWUgvb+CGN8HxOdijc9QZsaH2gWB
W8w5hFfW0KLvUKmbdT6jHvKS2VHMRzkS6lChWLOucnQi8Nv2LrBZzwWgWz/mzorI1ZLtjOYJSvBN
tPk4ruPBYS0J7bn9H/WawkuUjSbXANEtX45PWXSSyBKMl8u6nwv/xAupGb/7UsjSpktkW8xBxeW8
miVaiHs157mF2OPi6J/01RJRAtehUi5IlarW/im/tK8INbHylnkS558ixyLJcwr7HyqnFiV6jFp0
hbNrgE9SVfr5DPyX4d7Dg5+a2XDtIEIHI2MS+MiTbBsNDSwbu/9wTRsmu65G8XBX5l0Zt2s99jyc
MyvhMeTGvrUv28s+RyW7nz2UmFGM0oek+WkPvMsQwd/JCuQfjBB2PxBdD23sQ8enOBLNnrXcdf0c
l0ilkeRBny4qCEU2bVV4wKBTw18MUmUfIX/Hrxcnm/ANRSHi2tFagww3GdE1iA/cr698O7eEVzCZ
9kh39SlSmwqCZRYna8oPj/dp9RcdRkKoaHcJBPxA2clntLdU/NfkqL6y5lIznfcAh01VKTM9w1qL
suYW78hOKqe2CR/RV3jJ8hZPPbYPr7X3o2I2c2OcKQLb0P1TWRcVxafnPJR/eI3goPLfgDpvwlCH
WbXspeiyYsU+SCTwsyy3xqJUILWBCCo1D8g/18nE8TvfvIHAD0aE0HiTE9ZHhJ1WG4CJBwRm/I1a
lobPvuAoOjh64tJGJ76rKSP51nPnu1iGBh0H75FkAcoI96COCJ6k+953vZw5Z2Qbq36D/sCkeAuR
QJZgcKtQlT8ovxPavTVwE4KaijjvKLKVCC1UwpK40wIfr5TM9MvYOl8fLn0CZRnzhGXHdL1hXCvk
U6ctvYLKLIk4OL07eZDgGJLud7I8W9UcnoObgokdpGa5w0Vo77Bu7TQmL3lmmmf+YzHZWmv36Vuu
8cOK9MLRMVP1RHXL6RXT4C0k2WFoie7kBq96wuM6XweHJqjut/mXwJH1klhQq0TCarEU85XC7Fxf
rvME9Yh3WQhgLAm/21JmXvV1GHOPtvjV/bQXYrOIhVKcb6n40Sj6BQncQy7aTz/HkAsi7/L3ksA0
18WMe6ljyZKlxkp0Gh4zH2hY6IWo3m+e6003u+aR4GHnmoX2odElo/QWQf6i/IrIP8C8zzS+mLag
9wuK4b3k66oxIy1ki2hRE+0WI9kTGlX6kx658y18OHfPjShz0MuKG0T3CeYNWdhyCggmDOM7h3zc
cDKE02cstmgZW/xJIRCSM5KrKyQQicNxA4E7M8ch7V4umsrPoJ1Vg0rVFBewDcwbRa+/y4lvqKHN
VnUZ85d/G/pgJiKhE12Su60SRIQbpDM7ISMqQFgriEcmRcQ7oN0om4hR2l7rCSIoDkVubvFYUXaf
tb2UmORxP/cMDkfkkzPFpCAuZku1/cNzkfllHGTQneB4FCwplMVYcNzfVo5vG41bUhxthhFpuWy1
bXvldv+z26xE16HxMlpRUTMIESIoezxcquzo5w+ieYK5QwGy+jjgntsReFdJlJD2AbgawjJ1aMY4
MNvhCLmxKCK2XRhKsysb0lihEk5L2S3DGvaumYyVKfbo8M/zFxS5BWSGm66/iyCTZyqWde2mZ4YH
KduQ3sm55XHdmvr/okBQgiFpiSjoNe5m+8QebRqcecaFE9C5IOj7CmECmKQQw/qVUPq9Phq3xjzo
zaRIzLFDQrDV/X+Z9zAeHqeRuwlOFgdpKeb9sFMqKtc2mNm6MZeD4/sUsa/PLbkvuAlMRd2e5Juc
mCgssypsMHiMM5Rqu/WBgInwstCbsw4MaTjZgNLE/+PXpqCaj/oYqq3rm7zqR5/3QMMqJkoLI9oF
AQtoFylhgqz3fDhGcqUikGmdyr/FKK9PtkgpFu+KvxcNHsRiMoJAtC4Ig9f6zm11a9gkT1QDzMfg
SB6+xedq2N0MXCHY++Sm8U01phoxd59fWNjuoAlSunuA880PZm4AfdqdyPZBKWVGfaWr0cfrt0Ei
9fTJHS6DlLP2mtuy2JwFkP5Q3xd4dDDAQErPz1QX5eiLw8+Xpk7ZzhkzWk1dup77c7Ygom0clpfm
GlSonbJxQyQ/lRkZnPuicy2csRzzExtSlwUkEMCK4qseXGA/U+PI8gAfV3ZwzDeiqSof1ZJZQUci
c6fHgbhxLFKdK5FWD/+LySUXqQq+ZsJ4wu2W+IHh79AFHIcG+aEzqgCq7hA7hHmKIv+pkZbWKiZy
c2q91bogxHEFIhBgTj6rVnuEWsaPr9a5pIj2Uzf65Unr7lZYrFV/ePATBgl4xnmDDzVzuLeY3ek1
6YMzgp7UlZWYA+Q3q3iSLaKpFFO44idfVTRKcerZyei/IdUL7bkHrpaUp+PHTkkH5w9+h48FBTVo
O5gEhUj+TKW55Ar3TymQbJryqx3JLGBnpgI8LfWBvV9XuzRRNSXvzFMx+t5N1EvKbcphLAzBqqkL
pIwwXV5l3Xl6ckKLaQSADrL+NCeX9a899JOka0F/BsmO5ayJr85e4rWLv3MeR65PxHB6qD1mLtcj
1WPnN5WTz6LcS3f4EAPRr21vNDTks0Vhlu4PpH4s+qoVLuw88OrwsCYyrSxaRNINPRzfzoxs3Hid
UuZr1WyA5bTZtWYkwnzuOQVhh5l8ZA3IrIZuzLRxlYLk7v5S33XwBtpPttzUdbt9OHMx+BoM5e82
t2Opd4a4Oa3kKsc4k73glMYq1rZrHnJ7IPV3wSHB8z/ssp7X+gEnta77OEFB91iaMa2FuIqPEzfK
XU3bm0bpu/WXOPmLqcv/ntAzyxi8Bsd63Hp8wteYjD4ZxDg+2w5PE3Z9h2/Rcsgxr6xbHk59Qh+W
bDrazFNZlFLh0/8WZNPEXGL8BGDC4x3RGnDBuPzLXiEskqgdsPuTmMZepB/93zmZUa+3ArgkLuYH
9QTgPak9VZGsdSCXivztmP0Bp4AlUjOJQz/AFQ56YH6+PNss62AjQD6rDK8kvSXm9A2oGFUIX4uQ
xV01Mks2CQVCyN6AGiOMH//WOviIwvLfKTHPzZGHROtjlRkQ7b1dEkf81a0qLpMoqlBrv1UOewO4
OEtuvecylgvdVPS98YLhUn0Ac2e4U5Ds0fjj146rDdqBYfu/oJ3GMQ441jCIiyozI/e36MUBAmEk
HH1DE6dHYK7ylZLC7dEsrTLuUsGqRw/8KxWKxtGjpI6pGCd/PqOJkmCeugGmrs00sntrxTchVvY9
RNHQhppfsRQQsoFxz29pJVs58MQPAjyK0lcftrhetqK/DymkvJqVLDvTyOB7Frq7bLwfnzSQ/EYk
iP4nH0OxoMyutMGvlCcQV1Cf1VdcPdvxrhw6uj16k/L2bHugWA4NsPrsiuCK8ZMk6lmA6QUmr5YP
nOmhYrWt7cxcN4XuA/XiBCw/+9WWZFF/L+QxSNDzbQhMO0h+M2fz3+9VNhbppSKxwGOOyhNxsG17
uJhNIIZp9SDdO69Z78AVdToWXdEplFhNiDWFZP1YbL6U5cZLZvWaMglpapNlhFA/l4abkUmYak+z
BBU4SuxBj08Emyrn2h1AgvL3PebIB3+4slWVOSQwVezyLGYSd5aLYwsxF3qy9yb/3+lJY9ZbbfcU
1y0sblwHB0LrhG/unXaGZewbgYBsI2V4H42nsvwolLZ58NI2kz4YSxnrJYW6Va9IGUEya3FDnQy+
Yiea9+JFojwNf+eiuWo7iW3B5rORfxfX/4juAMii7FK8cjExc5KVDrhFDobcYTHRPW3ji4/Ls586
P5Wa2qnz9DtE37bgBwg41gkCJDmUXbjURysdj0qjooRG/6xPRbf35OoxC9xS6kkTC7KeiDQNCkHc
IkXcjkM6j3IfhDoIPua6YLhqwSOhpO/mzFI5HktswqYaTjXTtt7al1oT3kxUad72+8C/WXQXp8lL
LdGyKC/HWuCd5crFHMzOH0DlwcStrb2fIWTDo8Jh7HBjYajTmHvqr5VR7GmeiXepr8bBhqMVHpiM
PYGrI9xmfb7KLxGRZPr5YG+J0MbXT8NeTXqoZlOwHPlf5OhH9koklBf8A6biZiVhVb/A6e0VuFKt
EOwjS5EJy5UHYcpLoVzof/QH0ea/he6fqEgdkj53f7e7M1b7BmsBUA2HMtCc1CuyTB2J1tGFIChd
5Khfr3ZDGJk3gNza1DLaPbDF9tTtvOQxJwVAKBs5J76zgnKVTrDxnVWTdddNBjCjnDWFl7aSkiIs
/EXbLlPARQgQAkHGdkbdgkxVXq4A0TE0aHyI/MIkyRdql2zQ/9FQiZyw0J8FAsL5bNngtsn3P/g8
Y4neDwFMRpNWaP3OM32XyRqq+nGuHuoS3/svVcT6HQjU9Vu8vRnA5B+RUgYLmnn30ZWDf78rPqvw
XlrwND247Yo5KOFaIKbqzqa4wmTcK1M/Cul1v6ytcihveKJ6M+iD8//ObxywZKZl2C6a9WL0hCqu
yeG4nl9ND9FObU3IjClBhaVawrmgiF3+0IN0Rr50bOIcFZEkmwQSs8yEUb2mxuAVCkFVyUdJIrYz
pTKqv1NHItujhTPtQDClHketqSOeFRw+h7HP2X63Z3MfBcSisYhzNLXbT6lE1PiqASOBLxotNWep
gzUspOYD9E+fI9Rw4IGwbxqnQREFn8QJZHbUYo/5UggXUXOTMNCTfcLM7CJPRwcYsPz7xUEfdltS
yoYovi3PVFWl8o2osKBEjQfU8CXVoSMGPf8GCmUiCxPSyPBroiFN5s0BiMNA16ukeIxzWYBieCwX
IKBnzrkAFQ4iTCIJdsVexlYuJ+9ue6ozKmIVUT1QP3KrCRWudLfGI7GcsaQztcKLY6vfwvmqqjnb
3lW3jTXhm8mRxI/JQ/gpWFvDCYuTeAp9DlDe5rS0FyvSaYZpeOODKu94Op//tzfGe8CZg6rUqT/o
p1c/j9oYAPNzwneSyTfbHjlcvzLyA5qn7fwazk6MqapmxAOUPcruTYGDsTFbDiBk4XJulTN5qrk4
YcGjQx39RenEEdTUSYpWRrMYT2mIw2Mdcrko31vAsMd32ZT7xLuv1ZbaPuOHThbRzfK9RF7KxTLx
yv79cBLItcBOJphKXEvxWCyUj7Yiv5m4g4X6nBP4SC3d1C1BMMhGr68xFp6m/E999dqJH7Ck5GZA
8ybf/3t+m7nGkZAQ3lzByEFV1QbNIzf+tE55t/4uuylQBAwVqifY++djcv/UHtKh91kBVIo3mp8p
IaiD+BuvDK9Yi75k7l6uUq3OF2jSIPrv7qhcjDzelzxvxWbXHI8kYeOUMnKffML+L8nWf4ptebny
SNSN1qcNPL82+/sSTx8jJvv9lTEi0YQXKp2CzMj+oT62tgiyap+wiZ6Pa+6ePAEo8M12W7RZos+H
K5wsNKlL3Q/wSMT/H1HmQOIRg5EUlFH0YIPY5nlsqB6DgRvVpzys5jxagGLmeeQAeIs18Pg59nfw
bTqqW/z2V6p3Uz8aeT0bUR9oIOXidvHcnO1IzOcrXVhQ22tkPjRWA/jDvuCZVBaQJmibsGdxr3a+
YECAQiDVyCaVuaSW3jr0P3O96ND0VTewY/CeJ0EEy3UbshVvC39tHlsByD5FzS17XszsgG8cwErX
YUB2SZGbRjpvH0hck+3pFuntZW4dB6YedZjTDDznKyCysDQGmvRCuvnlbPJflRrJ1pqUk1CmaJP0
6dqdGd7ZRf0+MNV968qUUnIMIqNSt9UM4e8oSvArOUVL6CFzbzA4TUsAzb6vfTshQa6rR3AACSVd
j+tKj3IQLsfaFYp6Ok1o0fzUW2nQPI/LR4eWvFn1RGLp47ixvJQ6TLCYiq6DebGYJOKJ+5StUF66
AuXPTdsC3/nxmWDAelQVm+iC9Vjx4FJQgkyGFiplJfgYGuhVsePnpB/wS+pyIQspARRjO3/LLr+S
0roGTDhBuOn5o4zPLIEqrdRaI79seKYOuO1TyVzVOxTwCBcyqDodUrsUCzJ27ISajx8jFklS/AGS
zYVK0VM4WGYl8hPeRfgLtbv/q6cGNHpbQA3cIdENEfRPBBSDRJpZGbGO4awcBUruAc0nwoMdlH+W
UAzRKJCe0Ten6T8FuWtKyufgqIAPXuVNihXTnd7szKSliCzB4+DBSBI8X4LyvYBt+wDDO+mIVS9V
XxzourXMnDJWxWnwxNNDmEXK0WHIFot/pB0l/xKkHnGMhnBTjxLp8/q4HmYm1T0lgfTaBZFhxjWW
MwlRol9dSaA42xgCSsruBSPsr/nsgof5+ZkoBT6/zt2l0a8beHdOssFYR1kwknE1msI4I64n8JK+
lN8vuHr77a2DrfplZNCHEGlpp6bn+oha7oXwNMtRnOtKRncsVqDPMjAn0XP9oilETQmHEZ8iDWai
jata6uRJV+YeZCYQkqeI15Gw5OZMY6MH0EMzA0ghPN80Zrjuh71vHVsmzV0j7G2lvuR7wIMX+Bwp
7PGB3ZaXV3ptnJztiwN5q0P4+MSF7yPv+xxzbFz51Etjl5FDfXaMFH4WPetkwlhi5lF+TXeQeuVX
n3zdbNadbo+SBsklCkwa0/CmbwpXLMFiHFNHlW63ovbNN+LlUzrQSYeW+zBflwoG3lFAYXZPPtN2
Qzj4NJ/bvl4IXP9Q0YyqJOH94zDShTNMqG3tvu+f+HxC+QCedIVaS5AGfc5UPuHpjmxBHsPE59Jz
y8TxG+WsyU6jkQcMTivrWUtVyXTiiWAo2CG9vCmWeHsm+u9rArR9ySZFMRZRDjuLcZQIFqmc+ALK
XHCy2uBWUnIDZ8cZ6Y7yEHNDH3ZkFz4VCc9rIlWWSANbxGRIyGPu5lm/lKibhJo1sC3BiQH9El4c
XOvYTT3kJ8vukeOzv9RNRPDnfouEZrJzPxTtRsO0qPna7efYy3vgyX2sQw/tM6LMh3dvPJjVuzMN
E3WHqQynsiMA4v256NiCG58GXCpbNHlsaiqGnvYXyjZZAeEbjhxKe9ZrknBbc1dmSARjpkYX27Ph
dBMjSmwgcIyJfZaaOS3HXC6b5xa3p7A3wiqtOtJPBTnnvYHtUwOA0E0GXgdWqVNrYalKN1VaoVDr
7N/cvO7MV+b5lfwhB6UOUsRRHmzCi80CP7Dhz3y3jZOSXp+7bRESIAWIoo+zPL/667/n9mDWJQ1/
KpPBzu9olysnoUKGlZgz/+5guPYPzFb3mPC7i0dWpTUHYxKmY+RNJ3/hW2LT3HoAxoeGnNa3NkhX
eboV3/927Q3bXRbqaTtpKzkZXQVg7opGZtAzViZQ6Y2JZyGAuTyGZ2z628y8UD0Pbfcl/trIH5/R
58GK1f5moqJxNjUETSlIWURhVeNzsJYRwH6r+oRCkfIfN6O7xvNMqi7tnvTravvNrayQL1Oo0TML
SGsMNVzbXBCQJP/jwOPPZHG/EzeaS6HqZ0YTxexnsaAoopD+T7ZdQ68k7s75q19WnSQo3TyuVoBN
tvriLhLYoTu3qrfVfN8diN77ClLLHgwVaesFVCTGSY77pg5aAVgEx6UKbz945vYpn1sfW0wtMBAG
OvJRX5yePT1c7XMuEQkb4LdxWhHInONhCzwLE/gfjlQpbFWhdMhy7uhu3AYaK9WXfuKP6WeRq+pl
D0iKuoyuLWhmxyx7a88X7stdFxAP2IFUfGgOU2OJ2qbuJQegrnBJ2ne/+j41YIw8oRxdAZB16x2w
cM8rS6Fxf7heKyivs6wxFnnmASb7m1e1/uUzl0X3f8XP6qyRSYTik8VBiXGmSBJSHR8H+SzWJ4sB
OhFGm6bkXx4AqALsacoCInYCi0enW7sO1lKLZYWwasgwHcJN23Te4TgMZM9TVR64TyDLLbmiW0Hr
Fhtr1nP4hQXjXaQq/HMC8C17jIIQ34w50TcvEOGThpbJSReGwI5kNFgDwtEKGN2CPCCjTDKFV+Ff
/0Xb/qgKuU54qwcQ3814WJpSQWSMmBLUCai+PM1tOuLyhHaNwDV8eeVq4h2uU8g/SaiutXIOFKae
L6n/zIuYww4JhG/+XKxiNY0hTPlRyD2hFSaVdVbwpv1wa5Hhj/HbjVmgYXDiwwPftqWw/nm8MHjB
VFZ+GnCegFt+h5N5b21yEwXe4HC+pq9eR4QQg6s4ilsIdDbMsvMsN+Fs4mCXpJEQs7DOcIcnJQrr
ozBFE5rWrG+JA42PFT16ZGy4Z3kqmRFiII9G6pl/DiFYz15vaepQxcMCSOC0md58eke6lsZemQ0X
Sziy4qEE9vs2NJktiCPYQ8kq4TOEABEc7gHbS16+Uu0u/zSenY7JIJYJlQAKX/WyyZNwbuJWoIAL
Vb7KL5laKa+C71AEEinxengGVbo0Xo8NyUsTmNc+63rFXBVAFrEM03fkNBAOJ8SPzV43ve3e9XuY
zRT0BeEURufQHvxBezzUC+sKWf+L5s3+JrPTy8wCMmwuOpftpLCsIfZz+F2A4pCUxyCZRa0l3Cam
K98nGsV53rlk3GCWy6E1yZbYcaF0zZvO5FQzv8PVYm6H3DtdctsB7sG3fAYxFtOv0fHjXa/d8XL1
udXA9FNc4/kl+lF1ArYsfUwjJiMVP5f2KM5jR1Z6+hbrxz0t7MC7bUPwheNBdlgsc0eICRvQly7w
EYMr+KV5QMnEVvgoVcMbTY1gwmR8XuZHqEtCqd1iLl7sPGWWU1o4TMtR/ZycdE0qQ5bRXPiHndJX
NzyCexoZvSzjLyPawORqalEU6KP3Nopob/IVCtwm3lQxNL3ZT1Qxe51+wlZLmwhIXJfE3aFoKY8W
9ejgIytcUKozANAI4nygqpLWhM80IWgT2hv1WeQEGtoxHU+F2/cMZpoaP0Cw5NRd1RwprxpQHzra
ERCjIkHsTql2X+ICZMguACpkjOTvSMDcOk8eJGm6BEFNIz/S8q/CM9P4J6qJULsdZ3WO9HhATg/2
JIKeFqWCTgeLshrm893BLpF9wxsm6xcaeYoS/ka4KmhEuMQJ27mL3RBeKlqJ4c7of/jX6mHJD+Lc
WsMvBbAzyHqbbGCGQAmIDCABkW0jOIlYbKbmCF9o8DEq969QT8Rcwb/MM2KNjSYTbsKJ1i/7V2fb
7yhqHQwGPDFn4OMR1couDUFPJukK4EFsQ2c2ExOLr4qxBb6kp0ZueaoUMRu35x+mDWohQiYM1Tm6
gl85e1yrjZDWx9ep3ooOZZw4x/OMqou8IoakEWyCpGnoZ+qtEjw/1BSRf6RFUNtFTxrlms+6kTLA
Ao8WFxD4DL8s+Jr7gab+Wqxnj5FnmoJ0SvP68pGnMaxYDCNgK2WcIHgt8yXBQVZ65wz7xl5gptOv
M5yAJeutaJ12PZRNuT8lQxdQDtZlgEZtMuMwjcocE3uuFDOWhgIUBc2zgMqRjY6MP/FQGlejxzxo
v4rF9S17Ic4yv3MYvoH2qRBiAdr4sDL53Uz0X097McBNFDF1yEiLrWvVhNXqnyrdmda0yP+lHnu5
T9uHlbN4Hdl9Atxj+al0Bua8chTmpo4AJxC91uaH7bu8InqtUaNLhrjpoZCbmwCKelW2/pzvIpD5
EpRbfeRJtSY7QpwM8gjI5KR9hgn4U2Jhc0qllEGdLXmhIsJOZejQDIlCnYcUxNwqmZHCJJdIp+M5
85JMj5H3JzrJ/ihN55TpFga3ieQ2VaJ6qB8culs4Tt1g/oTI+3K6fajufcjD/XM/Xs7NDpw2oqyj
/MBINisbGwLMZWCGffJxa2d4xSRuSGQJYlcENKeax8l6d9RJSQRnCpz9mZ57mipTMT7K4mtQvocV
zeCE+4In4rNfBWK/HUxudgYKxCHiM9ffrx9jfAyyn06wuemBCqkPV+xZGbi4peYQqJuty4e8Q1rH
aqt7niODwMCXEpqsDBwG56xF1m4WyWpqrjYhjvqkdhcgUVSdpv78vHP3fb9/fX6ENk1wWtLoeEzl
NnUKPtG7LOhRqupvYQUx9+jG6R+ZMtsk/oi9vPS2DNlUj2DL6ppMlx/wTKWjQlwBGCtSZy3i9+pi
Nv3g71KVOLhQ2dWAzbOvFl9Bpz92mpYONG/PQD1cDqqqoSyfscID22hIhxbBNCGVoeMSVvn7rubS
3iCyaIBUU/FSY2cCtPNlKUnEiGJyOVMcsVUQQs6Frv0WPeHtRcLzNt/a16oQbtDeZQtay1/Osrzw
AXHL66Wg28OVfNzXG6eR2P1o0rgRT19OmAyUT+XJzsIdBrzsbNGKYoQMQbq5VMHto5Egvzzns1wG
Jg8fy6FDnTdpOXLdWnVlRoizGHL4ZMGJct8euOhlcMuX3cVe90ADIgElYuKHwypi5IaKo631V9dG
+qSLDhMViBzTBCgc3HLgWl/c52MDaSYwViuMS7ITYZcoLfz5XWi3L1G2TPoS9wk5/o8SIgkt8Spv
tdexFg7kGonO5bG/piyRYVg1njZhMj4yohYP2VTNm+0yoqV+rwL8QEQquVccblqxYtAnXVJSWjtG
BL24F5wc6L5ydSwkGIu96+ByHxsZeDEIZOsBv4iKFl3Ddmy435nfXvaFL6jVeR1mP0dgZQ/IQRC4
8YMm41vE9n4z7B4kmo1dNya56TVSEzhiiIsDuvYnnxbuj7hiSy6QcxwuRxCqpGOD376PSc2G5z5z
WOmRWTCGs0my9/OM6qGRGHBpqEfqm3BsbWFoLBQH9JxwpLTTUYghWydpmTCKN673bIwpLpWm6cSv
8AKWJCrqkqSTnavjPdCtA4tDopkBqEqXjsaS6sCiDXTkj6IOuJiztM/uieij06tuGhqSgE2/uqa3
YMWbR7nNZ+cIhRqDMtzU0Lcas84pfXsAmB2+27QqV28YcIsCWOKlX9kVSm1WM8Q6FWf2PP9e2XIL
ozVhLraG1XxZOLLooFXy6Gzh7hqcGgsWBcNizAXb5SR3pYfGVENHbdRu0M4dIXHRAU/2wmXVW1u1
8W6SAbELZ1sz1bwF+VAFQnhxi18jx/NWS7ncclnvngewofFtAE7J7gHpnMDO+Iu2Ij9hiXc2byFU
QoJl3+QfMsf1pTwelaqMWyzVtW1ho1cNOUTq2Rt/GNYSBg2ODsjgyolRMyajd0b2AuC98us1i+wa
X6W0nEfoxp+SJfPTZATUdRgEjaNAwApE/YKy0wrzBkDI6kxuYTAi18RpUTDPiGhuQ/R2yoRqLjTa
oZ3B2BMZ4WigIsGTd7NIMsIym8xi1cSTNc0lGeN1otgSOjoH8yyuotzjfdUFDRmcjOEgUD1Njkdy
E0P4N3I5ktvwsqVAausZWXpUJXxjsC9A5CKQU2n4x88IwAoP7uyN1B5BBYlF1VO+H+2PFaERNT90
R81yUf/5HbpZedKE3IO2hg7+RKCOpQ9F7+CoBqyhs/frkAk01EAShBWGFOFdwLs/nClEI0ipCO1e
W8VcHFOUgXnBxQtUO2z3EZ9mQg3fCgcb1VzfxnD0c88MI5PRXdGZWDWqm92kkO4n/mWjOZVDvY8l
GkAe/hu4t60PFtcVPGyQbo7D/T8xqGnPj7yo/4uYWuijn99Mx1A5V00SZZ8HVg7w8N9+Ee6ISt3x
516eVkCzbzAc9D9ennYi4by8t43lnkJoQpG93tC3lLeg/+Fp3Rrhk3hy27hZd4u+q27Dj+Q1/I7y
sQIWiKXMJhjpTluCVfUMqAXTK/Wpxvh6s1UrWDk9v4Jp0XGYYJuK5GIWot+g1p8fkHZQRMMtcYvI
si2Mv3LDaZiDRzavhppcBzyeNxg2GwTfFf3rn7xk/22g3EOZB9W6qWQA0l+yZdAaBPY36nYgjzfF
RHebIhnjL35eHFmjk0GDp37sL+Wz9vJal/JtgsMbDJWw/Cpg3cEMkR8g+8/qphzRfxrPCU8t1GPN
LP850rUCcwE1toYV76BUjLoaoCqrDJpLTMC5N/eiyUg0UyIwGVqOwm3N6dV10Q7MiCd1kZ2sGqUP
zadpREnq9LQpwmskzS70SfIvpZho0R4FIIYLUZq8AxQwfEYhd0SRJkjx9JhVRtVOpI8wI+gNr9LT
/2A9/Otm4RolRzwWV7+L0L/wZmQGnappjUN21ZTKtvw/sb4lLCaYuQBUBp64mgR4NUadSw7IW17Y
AEP5E90zOkXnN5cwW+yXhX/KE+7YVwBkm4cbBKWTKcz9Ke3OvdR6ugzvEjr6IrarY14H66jIFT7X
/Pgz1VjYQ99PRmuEzAZmUxVNAMHCrVoE62+PJu3MwOQvMycTued7na6/sE3d6zqy0QtDbTspEKBj
gNEcdENw0F7pCoYX1CH4sF75QemrMOO2GbRWYJmbAVgLpM0HlFFpzhBU4aY4GvTtnjnlgbqEQP/4
zFY6RYQlSVuR9+xD+1QV74SW5+ma0MP7qL4RUMXBQl9B/2hl90p+Dz5ef26wK9zNRjbxzrWXRvbv
GG25q6mWrkdn/K2ra9OiAi+us2xGODJUMln6e+VIZiM9flqmEFzFZG6ItszOMRcUOsyrNVxh3r2p
KSb/jm25jfbZLv1enG0fp7xTOtMd25a2G+0vgT21Uejh2TVNJNtFU/m00ErgDyN33aOT+CTM3GEn
1dcsB5HRv5DotJGokhlOnopiIGywf1uUAcxfjcOdYuFKkLNYfGB7fLpRXszoou6pdcpOsfb4QTE/
QvQ6cUhDBpuVo+nxujylutyVFg1+tYry3n33Ib9sah2VkuHQ2pyIWr0hi+wMCuEHN4z0RXSdrwt6
QYsJQ5ah+cwmdbIy+MNmgWQS0S70lP5+l/S92J9oeOqW+83ZqRC7pXoZBdc700+dmuYT9E5uagYa
Zc5zgn3uWeHNl1/LdBLauVweVMV6ncnEC3Bw/1Q5pqb9E6fXFjzpwG4vLFFngZU9CdU0tvrW/xd4
6FQPt281Faws+rwTZX7wIovuQ8p3x380yC5eunb+JEieP8ccHnYK+x5YHWzGN1VFZGgDcPjB0k78
QvtkjYo7eeYT/iIZ1R+8xkZF5rGhVRLgas/RpamGG/ugcOS4cEpvyEXu4Rp0Z1dO6AN6EyFJqRVw
pNoTXhI0oRfE6UzRBei3gwyVEogcE+o2xlplbgQmeGGAFWC/yNXlyyD/e8aHZJVkVWXSO/lxV5tO
0IY2o2Wx86qRlrcy09WHxXgZePpD+F+Y/Qq3CVDi/cew/qFOFcI8atiIm+AytB4sHp/TUs2RXQLk
FiyxhyXVY7EQYhkWSmMDpr+rkud0BAz47t86j0Drtqemk1F0F61W1IC0lSIEqCRuU5zMfPW6lWx6
xqm1l4cMMV2uWyBVXktlANNVRqkwS2VsreajErTtaa+3R3QbscY7/dkofYN2wQgEF+36T2vCiZ9f
XFaoVHclHmLD108YXXBPC/B84RArmysb47xrA4/oZxm5mda01aM6Rqc7CM+9DCdhwQEJSTk8phDL
IThIVWGdFFvg2Kw4YxMgO3V2RuSLpTz47hmTfo0Mmh6mE6g+d2ebXQ6zfZ7SAwEH8bs0eDvezlFR
W3/O+2n4acpA6nGxTXKfjZmpeuTQwoeG/B5+Ud/1zh0hvZ7jjN6fjLkjgIiG8taU+Lp66V+kWM7l
UHVD+pw7T28h+x/0/ClUjkJZvWJwm0YplkuN+paYLcS96KPIHvooF8hYtZ39x7neSCBikeTK/fb+
oN/jmbRpEUyARWDeC9HET3/dDFubsiN3NmkCZ2Do8YKtHkt36q78mST0c8WH8Rv8b8VSS2rKhLk0
MF1SvPljUpIU0Sc2ZEnSm3iKvgmG4bgYZl1DHJl5qXV5EkbqJUqJBgRQUUkpdgyefDQ0SSzv0tgJ
xvpaJ+++SaFWAHMQ9nIxGPmStj2nJM0MaQ6GDeDZWfn5kW1kK4mxUBOjz/yx3UJ5uh5o7Gls3oRx
WlDnINrY7wvbvhCU91OvLdHNM1lwWAAWfYgrI4dPcj7P/zu2OAPF/42tbWble0hbn4aUCmT5APCN
sXKKkqd9kz8D4e1Lu6fz4j0+iapSTjaXA422OIdRHF6qIh+5Sx/GzS9iEATYZ/AtzHcepUMZW1Jj
/sFypCn1rFcKmBP1IYq3jEGbX4vSdPKO++ZcLaJWKzt1Mgijqa0/2D0PX1ByRHmOcylQs9u6SpT0
PYKG2czwt7RVtGRW67HcOMNCJeij+kQxrTSKTD/zvejPUfsDPkb2ZLEXsZVkgwO//aoKKVeb4630
3/ZbHStfrpl86YQw9yJiFqtydX/SDTpmSbRLWypVk0UtH/u2JqHF50wYz/xflc7Ie09HDKKlkd3N
+4E3RJdOd7LdN9y/uiA+Rbgw7ucYafRVcvCilASU6WWRW0D3mW4agIMXqtYqr3VJUSFI5TZxy+JP
Lo1KT5sKzdxPyCMZWZ0l2QlUtcLOzBKCyYmk5VJ5Sn+jARkO39RIu/rTCXAWVV9Ice/9YoSPj2WW
Jv48gEfieMiyWTW7ILmNy1OE79oetXiFOV72xstSxvl50uianJjHNjXebKJ9bhkd5zSuZc9muDQv
FiI+ovrJ3NMHX2Jan399UqOn9Ls0OCTgE0rMtg26pC2nqIdaQD1kUfcSE4hL4bCYyqTk115OjkZU
us0AYgs9FJup7lbEwFckpGJNYk6SGjAR2/lNWPsQzI7lLb5DiUehMajlXUFAL+7aMddkkwVzOtcy
gzElm1a/ih6rzeiw1Bym1CEYSD3RxD4ZecElI3jkjs0YNL4oHhN8yMAzSgujhSkuMTfD+ZiFkixV
JcdOJjCUGkmLwHams2etsaWjUpjltbUY2loa79MNMqEn9f/DLCuAAblgj6jq8CQAQueFuPrK8ku8
ZddXrXuQqWxW7UI/8wwJi80EnBgtUE+AZbwcg9ujxLsrSyvXK/QsJmC8BuHSszcYHstArPSctldi
bi0/d3WhTzfQrOZ/ejvt9oKxLwNDDtJSqciwnQeeSnOkoV7AIlDQofQNYKmR6hpU3lou3UtuFNwZ
B4EIeC79P0pOyA/C3DzwZK8eJQzE3iYIYQIYGZmf9MqGJBmmh5HUuERM3+V6gE2hAP6F1w9alZNF
oJgFMf/kJx+ZKpRQFD+toW1vdY+8NRLSH2sURpZYUVEqT6FsdwugjzVoGwCNlsBqoR1xL6OtFJbP
fg7UmGg0a2V4i71sY6bWe4JXhqOvwzlcpAesis1gPvHCmj+s52dgQbOsH+0mUqRvR+lTpU4t00oq
Nf2+1NPegBs21QG36aE2JaCpCNp4Fo3ktYLIUpYLQyoG5Y3VhJefvSpgKNiAXcwPmFho62QKqVLw
4lL99zbgyyPXbHAyhBLtc4JlXNYGDVWq6580YnMpkpbrb49FmC0HeypxaFzgdKqeMAKimRXkjLlP
mQP22SU/7PfOLYkIrjCXqCC27Pz5ppkkH9ms3Ypja5XCa8IKW2uO+GOkKbv2Oz3PoolSKXvSTKfk
mHVVQGsiHF14ooZX3zXpc+fMnohbhKwpmMqcJb35yTRmiNmZKJPsScU+s+S+A6TedGCL4bmCjPTO
mR70/ig9ucU+jeezZKg+60xQpks9CGvPlFIc18QGhO3e3rBTOnQ+uEbxf+KiylhKW9geWyU5tZZ4
2xCnJ2Qab/jYWoLfj2U79cf1JCu5fSSCs13QRQhW5HXdDsCf+bYFi6uqbkXpzbt4QXx7sllp2/+w
hqSqALXE58JcKEH7z9aflSwNosucPeN3peKi5VM4N8cxdyNFYw5AW5bi2R4IEdSTdCjnuCgduuae
c5k7iOZBz+cawyERlQMmH/A5lWC7buJOI88Hi0QXdNV26O56NHPBzMz7LqEeLzjba7ViHLAMKMV9
08BYJXCS3A7ja+tX4EQw4v7Mhugf7vpWpZkwIO2pz7/I44Xw2XlXQKvvr978j+1qQC9MweQbxL36
K0c66xZQvUHfo4u50+RuN+1BE6F27Ctdit79Ioq5yzr6571+sbgRbVTd7NvI4UUXe0JygZHUJK8T
QSkByH4Gi53rsOoSKk6FfmMelFPcmlHmWC4g1NedAj5YEQXC0/bVrZ47JpRC67IRyXn7oNU1aMw/
YBwq6SOXORI7DXKDRbJ/7G7jfIII7n2srlIkCrT98p7lFZLPHMjEimd6JX2HmB/xeqE79MaCMufh
7kwtXp+xhTMZmu3ht/jfVZE3PXipq5ybT2l/tagtk2GoFFWXBnTyaGF4oQcYLRaAI+enWal9Paol
GhcgvOLFr2xVpi/nIO3etIO7bQg2nYSmlPbqHhwqMCRHn2kPjHh73r0SG40vPoEIyl96UyxTMo0V
cok2EGGIwPG432mhzCvFPoHeI2EASLI8vMWcOmo6XLIsTyhucgSlrOht1/Rt0I+U+w16xzUlD9Rm
HV1pmXgm4gQQar95NNGlX65VTg19EtZM7Johvz7RnJBPkFa+Yz02JaVk5dGl3VSvFOjroP6cr6Ph
G9I7hw/i1312p6HebDMZLWJtstwVIRTRRO71NdzNZ7hYrN+QdSvLdutk9Srmu3j8lxbyfS2KrCmF
DWcnooDIqjV2Bh2N5vdd7Z+7UMKIIivefDx63iC4EOJQC/eSqs5BEej7NTAsT9swYgV63BpnbeFT
GMtUmypWYx8jmIUh7J3dWrx5uCdz3x/K3fykxuONn3T1veX8icMrt5cfGub1b5gq+uewpbOExR3r
hiLpYsl6o0Lq9XMAm2yJrbqtBlvlWUcXCwzyJGS6qc/3TJtYzkpZ+QsYKgcNIxrUgq4a0ubcu/Ud
ctJRYjcyMCMpGnahddE5W27bGauQbfXMHkJ+CVBcvdC+Qy9b+k92GSRrVeyjtR/4whEnuhHVycn+
1SaJqo01+8JkbowuIEeyp4ErCQFla8dyKJzg4LlGA21faiN7cg3bTUi+/nl/JsDc5TGldn51+AOo
/S96A+14QnyJolUv/IEeNEISqQpWhI9sDp+dpwFt29IfRQ09i5VCG4CrDqwEdFbtHBfGccKned4S
wrTVlV5ntkZ3wTKkQB/qgZcBHlq6OuEgk3aB/w9cWs7IfX3eoRGIZ0aywxbOLvEdAWOxB0uO/Ix0
/Nfawd+1zZJmlapQ9iPJy+PfsmBGKdE/YCcyBcs/YFKvk+GU9Q6VNLc9n3azt7IHMcwikUd0lD58
Bfvsx4GdWkEgXewRm+pbO362NeQtQ7gy8GS3ymFrkFVwkvufahbONgBiEJu1He/Pon4mMn6BbTgU
4yagrinq4YBBlLp4jv9fKXGq7BBAv51ajhjP0mvfo22KYrVP3cD8e1l4k8H2KZDx7toKIMydXBGj
LDYtD1927xIZ9Ud3puDaBS9GMlwn+W7hacPlSO+/obLEF3xNGVuivuRi7V442vMjr+mQp/vl7/Dt
gZ6GxPCi7Cg7mTwCkt2k5PxlkwfFOjAKC2bZ8hA19TOU+jHuy0oliclKy1naa4ue075oM2LvQ+R4
29bp6vhAldYJlMpSt1QCb6NGDlM74hbksYsAqMWDb4gmUhrZ1sWm3yuZYohbBSMkycg7fi+anxE0
mxJiPaEosXZ8euN8PGhg9M4eqXiuLf5rsn0T6wefSB2ncCT001zF7raVm16jb8+zOGHsLRpgV43n
CB81hWibDoXdtNu8Gu6lnBFzMzr2noSg21mWwuvAcHskX+B6nhpq25f+podbcqElrfHCjoQ5xtBI
KIYsyV3Ta8uGoQvrUcXIQNvKqF8O1KP7PHPhGSUalNheRfbOP/ofqLXu40ZQjyzG6wjSDRYK0bp1
klLESw9uXlrS95SI+JWFwfvZGX9mQIi1gaSAJyaGUgiw7W4nAIVGBZkFtZSrgoPYVofGzbSa+7F0
EFQRG1nEsTVtkXIkglAQDHV0ViVvGtKyuOSJSEZ1ZuMpivF084xhNwgfd+1eYihxjd8bSGTRYWhc
ecZoJlWFP89x/mw8MpSEgjLYRhUEo3y1abMfTFJ+pgwzsX5E7agfGK4uiVCYge2wbP6l5GCI442I
ZgEv+onJJyGmZ5pUO9yLFLB5MHd8rtKaH9eHmZL2EKUCzJAfyyvhLs2crA7cIZ6cwwS2BUAffP1+
mUo8PqDeMqBHwgNszZIrCEMbwFQLjtBtDM2zoju9CsxV7wnkVlmKZ+r+zUAiHsazK7ZINXIqdsc+
qtMDePYseEkm8TGKO4ZiHrU6NX/2JrAFxxjX3AHric18FOhZXrx8f70cJQ+rTMIf3zPKnksclDfE
JghW4weUnIt1A7qq+OoHqrgEe4UdfxMMz8wrStmnncNTzGaQ94enOPLs8wSy4BWMcg3zQsKK5yiy
kdynDydj6yJuVZfZEoYP1NEPhnAZHbJTmEdGYWNjrzltqEfQZdcdqOJKlGTzgzHNYtRss5RgTaJw
UaWjC93meclhK0exCl9eg5/l1iJ+Gij1RelzFwpc+gAtRwIl2Vtt8ogxT02g+GR9kXhYeSVVQ9O7
jLcsIxoF/6IOq1WbZ98boOak9apCjPp9aGHk6+9i1LnUmUxrDXUysRzjaR+fH3H3zcTGcwsWICdx
RCZwIxTm9l+53ROHZHTU77+wE5UPkpBnOn3Qipv++HOYJZgDkTNmb3+NZT2MoLQN6BAp24cOXZyZ
keleYjm4nHrU+Y0YAaEwbGNIzd2zgIIftkOOy6exLrv9QdmhMG2vDvREdfNKKj42zHGdyBBqK6M9
LzrxNJvzAeHzoRoIVqUT0VjzguWxvkjbyxqsgdxtTJ6OB7bE7f1qNPRqsnR3zRmWm5Xjda0r7nn8
1uUlpp56hB2d8LalKoJd0xjJFsxAN/Wlt+7yp7wObV8cEYSd0MDW71lDlBcWsyp2/rWxFVLqI5aP
vOUuQ8t0fLUxRAdfbnzkMhuWupok47gEDJBIYI/7+xQa0/v5TGA0XDseLRg5ilCXDp6YokrDj2g5
/vmLXgdzcost4smnU0hWn5OATtsicSyB81T5d84zu7BaoqGO4yfeI9r95FsaGuRiSYNx/x1emq6t
VKnn8isK0IWl3RAZCHGdrQKP8I269gQiEKxvUJOEQo4xLN20R15/VQalIJfRocoxI8WKTdNairU6
rgnID7uSQgO80mr0yNkkIRlHDKpL1sZwsD3xJkqBdmBi6DoRPcksopBiti2LHmJJ7z/4ptQssGqf
PElHCRyV0mIfu6a7ti12nqS7Nzh97qhEXegRzSSVOeL2qFptCDx449FzNSp41v4kr2FXDBg/iHYY
R5QsoxZSBKglx8BNAMXGZ+MUymlWsOjVf5np7b9bbUXFXkNZUmtFGRNe9TvWg35Iu6tf6C7tid+Q
gA9pid7yQaAd53v7ZqUMSpYB3EyW0+kuaKW2B4LKCsdZqD4ppNrXy7VZreoi/c+lg5EMRpZv4GSM
Ks56X4F3iKqBa7ijluGdBcuZlzeS1tH2gfEA4/yJuwPktSimeDcN3UqN6oMI58Jhq+o/fLf0JZp9
dbxqhzrsZmnJdsQDqbcWeL56JHuEThodMEFYhmG8036Cb15YCK93eU/gTl1bMy7iQOXJC7q01yI5
35ZfNN/sE0Xkxa+x7nYtOQGMQSvqyClcp6G/zY6MpS9A190g9iqBnOjIoMagtX/39kEN5hY0/uzz
Wy3ZlcvxSJ90xcr/DfIAoMSggwlm6XjOgIx6I2ccNhmr5YazL8XcBOk3TeweLXSVLMntc1jH1lRv
cKZG3CT2REiDT/gFjTuIqDIc1+WJai8+QWJdewswN7vBgqs6ADRhQZNrIuLQaLgkdCdwQzrJRAcQ
tKagr0imQ5zJ2ikPdxXz1sf5NHpT+pSDe1ApbvHbabGgoVykfZo2UPpjCLlXGaVCKcrnz73SwK16
jXSvlDVlR1/ND+pNOn8t0A6P5ou5mwRtaj2nQZwfN2H0ydEiDTngBBxz4wP+69bKuB8M/zki6BAT
b8bU1cFqk9feLUzWmgM/wpF207VdMqiwqkakupCbUgtD0ONhovV0YTghb8XosIbW4BlQMKb7x0qI
h8KszybUwUB6pJODKnoIA0NSBu1p9uCKUWUFuES4Il+nQ0ZBHtTc9iPfS6GkdPmyGgpBpPPEUsLP
iZz9AsW0pFTx0gXJwtFilfoZG+Eeudv8AIC5enfiC7Okdq7CKCSouGv9H5iMnRI8DS/pWWel8170
N9JKYqrLCl7nNRGgmK9M6vCFHuff7nt4iLLNJpXbewdU+Q9gyEO5f03v6yyqA7yEzCTgSbfc6hXO
aa3jWOhL7JF//Jh5NCm3yMIyMtSi8P/mTaB69rC/9xvTthD+F44mBDN8ds1cZBZq3ZToCsyGFrRH
AROJj7eWnWlOcV1kE6NHCLrwvxWPQNyjyUOXJt9ue7RG8EyNAxsydcYy8ez7hObkpzORU5TuwK16
uy3Cm09ii8bTm6L1B2EbZL6IEZLjZVVQc6OHRYjPMksFo4dYg8l+mvSxbsAz2MmLu9Ikgawfd7y/
iElbZV6AejoB5qelJZl4lwRgkO7QSSErce+Yab/CBAX2DU3HOUjXK7RusxRDJXvbcdrbezdkkc5n
HcivjgzHv1DMXnZkJlMpH18H77jI8d/7WsfMzHUCoUyl2QdL9SaSukZ9S5gJMdgaNoUG9c1qdoWw
DiXYxx1YtvZLjFqeU56P6BFpcozOLFwjxGZ5NnPsOIzTd8HPMpSMLajdaVpoJCLZXtsroGu2GYk4
nuLVcZxB5LmnTWbThjADn9p8lpx6Cjqc2yaS+dXqzEKTQV0jBtmCTUFWUFbOVBC9um8S1MW7+hNu
Q/y4SxHWqRW/+569RQ+hXEv7fqWcPQAj1hVcGKjA+ONHBjD7GjF4L47VEauMwbiE3diRFuv0xJ7l
D/mDGGTDEDRIepLn7133E2DshwryHfVzp00x6d/bwn0Ho6Hu+DlLeqYzWKgUfHJuQAc5N4vWKNWH
v0bXXcv/MghLfBmZqeqIBiCJbTI2V20nF4veoW/J33638i3Uq88LI8tQxe2KmUeSpPs6VXd/ZTIg
5G8lweA8ihLgtKF93LiD5oLOUAV+mPegY/RG88R1swCUCvk44dsQAJnJ8Jgisulb7+7kzqrrWcNA
TN8X3ZhfkwmFmnc1jmcz/hBz4fGDnuplRTCP3e/72h4DId+T35hdFP6VJPdmI2KaNXYi04FfGNbh
XCnlvpGnIMDqVzYh5VABC8zFM9hXOpIBDlccSIH3mdyrp1f+ZA9JAPROwODrzbppDob+saNugooH
qja0PmBtXTAgV8VmnVewqA8UFten/7g0KWXpMxPa34g0WiNqaNBmRyT+y6LMN5s/1EVTAzBALTiX
QZXzxitPMKlurq5vlWBmmLx3oFzAIoBLf41ncW7UPjrfY5+P3sFGbNt/0mVnG4Zj7Cw16HqwdToK
P4Km36ryEaIogolA4YE8cr1QTtQp1fD9aMgjkMyXdTDKdGgfuR5E2seqjPeZK7pJvgq+paIvtobL
lcZgc4Omolq8giP/3iShAcqe831StcA9k9A5jPjco0eV7T6HQvLO1nm1TN4435mYfLxhmw2BsgJX
a8GEt6VHS3gy67uhVvWs8+h/CVfPryvQM9YNdPPyr2ekSrdXujPQc8Nvp/rWaONHt2404nruvXng
WqJ+aViOmOvjgQcgt9ikFz8AHFuJrnf/E6wcf+F5aY8IEEB/yqQrya/xD1lqCAiEP6+85/T0oZBq
T5wXeDuOM/b4NPXb55Pq7wjuZEExHFEHUdA/dtXMA19ksM/kDJ8hl/3m9/jl+rmlUr9gIcFdp+W6
axljTwlo1UejxoxNiSMvl2SniC/2ZDuhcWg+QsvZ0CCoec+DdfQJqNe8j8+2ubaaM4Tft85kdLCz
yBi3nBXiJlYny2vPxbenDF0hNNtNf0HDzGoc1hJYN/VRZuUw4DnWkKO864WO3M+2Ai/C5lUaA+O6
tbIfU7/hdGji/vu92AUOK93GKAe/HvvCUtZZ5ENpQC6kxD7ka8JV8hC+39kcjsDcHBu+6agu7ZeU
pdZb9zmTf0VGng1kIF/97BKsSuvk/8GsafuThOn9ARtzhBnwJu+M0+JwSmm6nknRI0+q/LAjUU9X
95E/R2fhAlK9n32xkXppHpAiORECBkUv1p/mkrE6cEfW5xU8a7C71Lmg/VNpEb8RZPbOC21HjH9A
+kGbW2X7Suc38gbgYV3nPQ+XtiI7UjOrckMNx/rqUuzPs5WvF9atrXLN+9CJxituhIdW71siQWJX
+6DkqKMUup95xC8ZCd8V+ucD33ev+snbgbDOvDQykyLmTJ6z1Wa9AwH0Jpqw8k0HTg2TT1+K/rsQ
oz49yLCykHNUSps0T1i5YlE9c2k3eY8qU5Vbj+a/uK3NeOKGef6Z19KC0085EERZjWPjBGPgncHJ
gZcXUSXGweQMekiUXB7f4GZaYb+I3o58zL/upNd4ffCsW60ExCi3PRpmIGpql8/Nm/pNM+MsxXyS
yIwRJGLp5ISsQ4W7P7mraSPPv9vC+mP9nITVB992tpGsKgCs9ZvbaW5YjWco40nkHC2DXs9FYoRR
k/zg1MHDW1CKH/FoAoRpBDe7efd4JGj62vaWSNgoTJ7S8l0HqESQIzvwsoFj9hXXf7vhPCXQmW5y
yxEvN3U41On32sR5ocO1yBlHntk+/2H6XNhcVkG9gk4pU8IOfgIcX7rYS8cE+QWOgngvTOIIn4Cl
/1sgiSuGvV4bOQL/7YfZMOHKvJKqqg76WzPOBdB5SglirGTSTo9jyXut1OKHf1rqDRE0bnYkhCLX
orGvu44ge9AbCCwRpqSt+fc9S+7US9ZkDiwUoFqsJptSM3ThZhNqYDyhNjq6CcozoFQLKdhBVwel
JL+h/zRWTaiC4Z57d1ahHTV77H+/BD+1W6qAGpRn18yo+yyYxJWXWftXbfAhUtFyIXfjLV4txcPD
i60QeMHd2Mf1swz2tANfDnowqkrrDoxwqLyFXIbaPe57hQoxOFfJBDOVpzd6lBr9xRDjoerGOrCw
9uuMiQFBpIdilihYUvdvR1Bie4649WE131aniqEbq/HZkVBqbT3v1HuGX2LhIkP7tzPTs1MjW0bQ
C809cdPFyB6hmPNWeOQNgoHIJ1Ig85S/1UJrmqHvQw/N+hfKBVIKYPiuSkNfAkvyToGXXfXWXeZV
9kjHoP476oZzJEORNhlZEmtK2XNRT7p2L7h/PQQhhHpTDr1VMgQB/JoRLmC3fUvJGaSGhE4G1RnO
NDB/214TUOZ6wLiTQLY+jOHbkE1n+ZJRnoitfAZOl1nRnsfVMMdS7Dl5RvjS3b1Aq0p29+hj1t6C
YfufnZOYXI+4nbMasqza9q1H88+r7dR425MzNO7cFOOULIMDd6jqt+BXKAmd0OnlciDGfGEvlCcZ
nm98nFtcpKcMjBa6HmBnqneUsNsoVlpVINgBtyC4W8TximEuZ3vMzMzy7d3eNWJLiR0Y8OC/sbh6
ICS2gfzk+4n0nbm1GyeVVleA97+va03Nu00eCCLs++nxuylm+Jr5ba+dSBLE52pXEp48Um6IC1Zb
rOHd74wQuLZHOitIizSiSgIf9Vk63FZbaeTzHY1bsvhssUZiySo646XrEsFdG/rIH4Wftjh+MNfh
PxSpLbKYC8l1as9BBB/Y/lnLW4vH9TDOMn32CqyQY05gq9D6/12i2wAUogO8tTu4a5HPeIryBWFk
0qCJ4sSQjT45vbvgLZAYirZWloBSYAaL0TJA/GUb3n0r6NawVJwFEOpuBrbvIUCWnTNgVOvU5oV9
UUm43wsnwSTElE3wxEKEgxFhGPr3+DPHwwmk6x3pAccMgBOdBVvZbLMzp4hB18fXueDQBRqEhQEL
oZN8bzr5fre4DOWQlJBGVKRp1sRZ7hrgakSu9LGLem8Ng8uo4+LJtvhQMfjj4zXnfCJfogYe74Ny
xFsiEZEsZkhuWtMn6Ner7WIIQaK9rU3P4zK9ZZMlXcKJsaNSV6G5yaMko9YqojlophKzyxpkV+mh
Gehqa5seb7nooJtmG3RpaWE+iCaPB97z6Z4ef80GLbN8ArYC3RHY5n9zXUMBIFbqHumN+31m+aP2
Itis33r7E1ogXkHC+P9ynKDJ/F1vhNdZ8ntTfzXdiBOTwCoO0cSPssvoRPh7ZmYGi5tn/HjjlISI
XJpvwKAKmQZfu4L/KRdxxB+trnkcgJ+tlIe20bcYidBn77zghDbC3tZ3svSH0FN4YKzmBZSXIrOv
03sz9Ae2O9svwNICWC2xiJ+Nzb/GsYe33ehucvld2XJCrv3Kt61KkLv3Qfjnn1HiMhJlf2qHMga3
nqAc2Q50sm5slhsOkbk/AdlDnJQJB3hyFNyGUa+aR+8M0e9DNDkApjL463KWTqJvtK0fhTfU9MrL
L1RI/Me8R1rli33tn1oXs1UWN1pDrD6R7tc9sQbUmiqOxxq35L41s/lJcPQNS8dbQVvd9ZBRFXQn
CfXgLDL2JeTv0lWaSumh+wgdeNhfCDtQWP5cQw7uTja75BAI4c7ld4yg/VgMGnPWy8VUCVKIdJXX
xCLx/bWq6mTUihYDzaP7TuJLDJyc8gMBov4hAWN+rSNu8m1z6gQY5bgLr7CBVm2ltseitXdaM8oS
2vDc3AS9umxMVD78fSYbGz6fDbM8WABH+sboOfUgyrq2RuxThjgI+//DTvYLsWSgZT0pvMnZjyKQ
o6c786MAal3zBhgSbTLZ8s1zMyhMTExXg6O02xVVLSW8gd/8sBK3hFaEoKDya6Hy1Tkv5+OgT7Qf
UWV36bYiPpCJ9w9lQISC7ugKC/fUpbaahtJDmVe97zmUxV4blNOEYAn3vKHr1eWNm2sUU3YTIwKy
E3Mx2+gIkBiQhvC6qqsAwQg/nhWsjrjMt86moieMgIcxrvlBoCKi9cOmux7lf5vGBu8sH47P7nqH
YUtvV1OuPv3mAH7oxtdMtyBoPlieaB9SU5oOlzTyyPSG4lq986NlXZlMEl6evKejlxF9bnDH8Q+Y
JN085KyXsAFdGkGM14OUtRWs1al7saoQp2v+3xBMjMwJlqCs5mDnUpehVSYBUtciFewDjmqt/ax8
HUsZcZaO38DqIZ1bhdayH569VnWWnVAb6t1FMByTDqmR6JocN+OYVmHXpLqxxMRJ9ajSZ4LMU0+E
n2qS/TFc0EUD2kXtSgOHHIxeLAT99mvG8YwPIabhEClBZAbpi3HQv6O+9CJJsHB70NeFhyGzGhyI
n1FlSfZtHLMt32Ry2P6FZ/jfpNK4tAgGqzeHhe85bCfnMrP88Jr6fspZ7Pv0pJdnXV0rJ9EZrILn
grk9x3WZrXAzvSTv6gLixi4VGDIsRO2O37hdZ5xtXg4L4MhhSjGS1UX3/PDArK7VPXKWrIJV4CXJ
V5UVIBIHbVTrLep2P7uZF/5B8N0gbdFUfbi9zDHDxM4PT3hkrog/eiTWh9soCJJCUZSwlT8ULSWY
Q/xvnLVr6oTU6U2GiIRxB8z/5aiMVWKLIESyJ3L1NFIC1pZlQs6SpMc65X23o2i3wUjWU1m79XGZ
fP8Z9cnY6mkn3Wr+UKQe26XKOxnzGftzebmJH0aT+UyKxGDTWRISctHr0VqWJnfy46MdFEQYfV5L
TDSRVGTNrZHD4v/fox67fvsWxgopZf3qVUy8CkKXlhDsHbT/TS7V1x4v9Mxq1WcC9ByYhqVOWN6t
Ru8yfjU76cUMrIOtZyEpEB7xllxi62QGc5SKNQOiV9llLwQPddK/ErQV82mzQWzThw+na3jKgWsC
t/UA1SkywAZZSBrsb8Gw9Houv0/Q1ANCaT2tppMTdnt0kgi8fkYIDtwd+R5F0u1sOydgZ6a4pGf3
KbwxCNhQa0aMD3sqpTKmATThC1G4fGciKS9SFu/IP5WXMNBImqSBYSLu7EwDfSFfAlgm82/GSzlh
0n6OevDtho7iZ2tTZ2O7IFeL17VErBp+i/dnV9GGZnjqfQB02WO40MKR3YOmXI5Kn1mn+eXtwgk2
CmhsvUXIYa9COSuodbpNwPP0PnEs6oYswqz8G1Zi5+JxNjC4e8DU9OgQZblozqstpNm++UX/C+vZ
yTrGz+M51MsPkbRD6AMgrxmZQYWFwm5DUQ5ErdFCVpPHyH2An/aS4RbJ6F/XT9a/XB6R9DTOYMwa
6RvZTBmIqX/pMJOID4Is5bWSXT55xSKbG2Eq+m4UCmX7NNkryRQ9OVPNe39OJDSJFC9kZDXgUe00
wLbWvbnGffo50sGrEz/DJi8ral6Sw+/RFa7WFUST4lw9zZUycXHvnJRlnXI2KNgGuxgQWF0E9DCx
My2M60N5DDw7L/++i8mv/lK6bplhcJiRgEszjH7NasuiruwIgi1qyfCyyS8E3rGVDVb6AZT0Gi8q
GwBNvB+DFRHd6UkXpziQsDtemvUabhdfXpM7CV1anBOpSdngjHSIEisg245yKB605MbGQZ+NJW4D
P3eiXG7Ci/ekY1gLpzMC75DLiNLnRUUiBitSwdOMz0nxEU7wDzpnCauYKwZfFimzmpX5jOJGY6/E
qQ/6VeYAH4pKpsv1fN6AiaJJVWvq00fxHqFFVHZorX2MXNjG6FnvYkG5lDbm9Cl4YMR4RbvcxlYA
d/pHcYFgDULc9sXbsoEC0mFqxrSV1Mij3K81RkwQEyGGpVqxoHW1LK1lwtWxNODGO0zDdUHCVvan
I6tEB5kplZh0v29huzlapx+DP4SUe5m7fyN5oCjLyqSoVhKySVqj0lFeNnh3pcYO4qQi37A0IDl2
5ZwBdZKYFb5pObViSC7gsHCoxKdURu0GrpcK1MA/f8G5Rx/JSs1IvnvxceA8aPxBEdlguvqfnwlG
q8k+QPLKtYipArb2JE6jsQPkMVIIvzBmqMuo5o4A3oy5dtFfVO5Mv8Atbqd5Wswtl5SJd98s4Yyh
t0am0zJPEC4l6LFM11AZa7Qq/LgBeMGOczOCL+KIrMyV3Ko5N2TE14Qd1D3IReYIzYjQ2WXpYxhV
xII++wQZVisvH0YrH49SiWuATSFmVWUurzIs8Ve5lV0udXv28sw7G+FT9ImnjmwFM9V6gfkxZ8gW
dB9MWzN8CGNl8zuKQ7/zPbrvAwcl8B52jyPmSJuG+AkYBrqZeYfQ7eIOUpIZfXuL+OlMHnKGh8cr
uXOxCVAS4OwQTVCygQJpTW8N7/22/F6BcDdNZ+WhGf59b+8QBe5zyxt6Q3ld8MMNqwhje4+C4pTS
Sagb2MTGw0QNfzHPcviKDsRNdkOmfH8zNPrDWbnHk+omkmxDmYVZJGrpr5ZaSnBvay9Y9LOzSMtg
SGwdJ6m2Vup70J6UOE6pUWXau/zAYp2LtFUUr6nCUD52xvS1MGQ9rFt+Z+il6LabL/ltIy6Q23U4
76Zy8tn/9g+h76B0pOC0+6h6j//vZQC2dN1MtSDj4DpPI8wBmgqLEA9lX3k37811hJFsXcGgLoiM
1AawTpqTZxZGECwcKV4/pDr6DHpOCdwgT7Ca2jV6fN6vL6jZN0nUUgwtdYO4p4TZrkdsNfR5dN6w
Rux7kmE0GSwIwoeQdYu+Xdk3XlJiM0KrG4DcmIpONn++UiF+Fi4llvcNl5ARAOO33k4qf8FEdwI+
oiZugyK5x1tXVHvHL79OQsN2MyMUQDQlIFbSJrGUDIEV/CTx8qphvjnevo7EDLIuetfkfZMO7UJO
ED9ALb2T+IK4zGKoGdRM9YXWUFJlaexOU80e/EqHGLWH02BeR7vQT+j41iCBk8UWBKO2WFVX5Wbn
P/qw5+wyn/xszGnAD91bqpAgJRVVDl+SGG60ZNCSK75T+zBmKbn0B0h0hs4F8wPU5G4zNZK1xCv7
E/GcSo6+KOxJe16T32uGLsaVAiXOT1v7FFsJcO60G0/s2M/EerhcDbns1Y/2HRjeq0x5r4KedcTw
QkYL020eTiGr+7vG4/Hh3YrsgtiCeCVDoPBo0nbzCG8uzsJBaK6vo68eoRMr57SXu/jHJUQcReFy
WKm6hAbPeOoJ2D9CmYqPpcFEOW0nVsnBMdYBHfRzIo6qpJJ55mICdtr0B18W0Pi1zdKqvVH3PJBp
WFyBrbcThuomLvzcr1j4fE9Ss0D3Q0sC+p61gAspkGrFrLbNV3Za9xYcIRCIYU5FCntd96QMVPr1
znIqHq3j7N9pWVExyBHUrw5Hk8QaHkP8PuRTfLss7s0qWhf0uQ20r1IMnNwLfBK1PmB0EPF0nS46
uEC9php+SJ/FzDHCw5duWw2VnfQuNbm+O7C/ww0X8K2adsPAnFiLWTSRKXCqdCE5HbjMPcjJVH78
mtVKkpkEC6F7oFeMy29nsgilYE0UG/Jlc8PBgOSOJ3aRmbd4hp63xTm1TNfK2tdPKbwRexXMEkgD
+g17jjf7gxp82/uqw9MZ8lFYJmbgcMO4HhqXqhMmZCoAZIOEaXTQhZQD/aFee9xMvau0l+7Lq9Lu
77PnXY3if9je8pcDR3MtzDJ7HKYyqsgxaOL2qeyvW7wztb2Jfob7GCSCB+1auUvTPL7s2yLYwHjv
/fO3HqimGiAc92LSVQLZw71qDB9xD0HxDfkfmIO3s9KU2xq8TDk+e/gUvjLlZRyfkzQW6k5NLRWl
E0PNb74TFeA8f4uZmM0HiT/QcBw6IqzYbXnlg78B/z3+5QD2JcySjkv/R5SAAx/bo0XXU6+zJ9w9
yXmt4wSs/DlVzXj+VUIF9Rw33+5Otiv3wgAYb1SZFApWQDb3GN9VdGoNsSmKOsdihEjj2BzjsbtQ
nk638C9eLI4QiyUuBO3zVZEN099z0ii+cFca0W/SIPrUhMw2gZGeEB6MWVZq7q6U8zBcPWDrU8Xo
aFIHgc1fpimxLFrRaWIsI2E07uZXxV3WR3dodg1PwUToPR6uLnntbNNyKJmtoo1hQKccOFpcDtKS
/SG+NsUncAK+q3fxWzq+U+rBNYiyIJWYNGmqx6uqnpAnjwMJE4Mwb/3J4YZErFGFYz/TYoxr/W/Q
1y8vEGry1gq8t+1VNOcl0rufbdMus5HtOO4W18/jrqIuJw9QxZ6ju+dTmwBE8yjxqAhc7qNCwYiE
PwUC7OTfj253BbYjWy4PrhV5HpGRVOYmRsc7koPXIZ8HZNDx7dXVPwfdpMcbqHVWN6/KQdcwvVh9
RWq9hgp78Ts040dAfR9ZCNPQFRTZc92T5uCDN8lpUq1InL06CNDLIjBJYcJSbUwKx1xaGTeHIrOf
BmvW2WpRIwl/uX7kAFulB3vKdPAwuMqFZTIXPTPVkkuB41Lz/7IFdiluTo0XB37eSf8oZW1qtDTe
j5VocbKRIUPrXIsXhrHlp+1w7crBBH2iLBsC5loQRr0XgO/OdRleN4deRZ0NxOY94V6VLsf9sc6E
oS8+d46pn8dGVBi7qR2HK6OYq72GpJONppuCGKcjJdXBzZjIFFy/M0AmbRqRdn7VfJ/h8VuolZIQ
8Hen1vTrjOtkUT5SA1lhB94dGyEQQqO6bx6BIU3wsXcfeGiwdMKeDpETxKZL351LHNZHsGsTMQKY
tJcOK2rLUAPLp9GXPdzLI0ETRKtZ5iQNKuqtFqA4lzzu2dIb/rbbpUV+0cjXlzR4GVYluvxmGP7F
665Fe93eb8/I7jWQC2AM4DO17j9rPdy/2za4qnS7osonXr1bvX8PyUCo+2PpGtDyuIyHp98Srebq
MUTcNAu+kxgwkps8t1TCJqhi8RvbcY5dH12ZPwkm1m+p7y7+H45TgWdNaPr7z7WzhaAB3Epu82/J
FWCZfAO0LVMb8HkMiGW8orlzNjujOm6aqgGFIvRpTqrPLvwcL5W5ZJN9cRHt1U7l1lY9MT3r6BxI
ZUEfYDpBinD81IpcR7zfnTwyezS3jDGWPPWlTN6lc89RimyFTJiSP/4RfOftkomtPuisWpXWLw+R
+8VXsdi0gDckRTd2zw4SqFdSPc/4hwbIiRejGoeKKMqeMq4YwUDgAGWbxmSUI+0/KSOTGfew7wMR
NhNSqKHWdNCz11R+I+CVFXtB1PIoSppciDk01wflgTpK08Chc9St3Li6td3sogkVo2J6vL20oR8L
6mabSb+JYH1V0RjChxbP0GDn17ThNJXWh3ypjPBMDQ8evCEKk/yo3iQlaXgO6QS4O+Aaz5pG/8KJ
D4y8zmDHdJj95JAY2Cccf74Y2P+re92I1jLy+YTem9PWHZNzQa8w0/EMMgJ8AYeRdIowNp7TOUyz
jz7RuRpbqBvL4hEyIjcnINgyNANus+UKgpRGZ3U1xBVk4DGquiNe9l8wLhcTl9dBNGEJAVCPXaVm
RRlXsXK1/Hg9UewIDW/mhs1Oth2TNyU70gWTM5FcEtDwO75KPkARpo5glFJQU/cc9WW9pRIuwPlj
ibkPZrq5wh4LWjCcO8EwsMZbQIXA03UUirnK9VreXzl+BuMxQRAB+nyBoBgi6yDn1vQTEihRIDZB
tg/G4bb7DaEGd7OnZrNDVs4HV2esYriSRH58Ul5kgESAcUArVIGI68xmDtT4adBQKAVumRGu+1ui
CGdSAZ/iyehodyYvc6hFek+rFEFhad96pMMa+hk8qF8zk4mS6aQ9YirCpSH4n6hPJNyL8TYzvHiI
C3GvQF2KzyoNPKyGMYyx5wOuUpm+NywPtR/nvfofhxUfVvSUl3Nyjov+/mqas4gfRT4GlRDHrdy7
BcHllJVHdj3w5gtA/Crdf4MygsCa0R/HA6ozAHPprAmguA8Bev78My1wxKUiiHDklaV35TwOC25M
wo7cA87KZThOC64nwT6+R8Wd36DcBDNlz/dx6ODrd3ujMojyk5zJDjxoBbzjU+bCHlQc61YQClgn
UHOQJ58q0ejjNvJoBL/VeRuwZOF65AoQ3abYDak/O8P3UYvjBt4eWbCKE1QptBsIrnJd9VW8CAVs
O0CLiwdVaHBlnlOQY8jHjBYAuvQrWug8d3KZ7IdL8yub7aNnDDjVzwH3xTsGfmWivuEhR7gmXBtK
7apYKmD2mN9cACcu5DGirLtx3fxmyNUcqVWdK/0mdO2c43cXUT+aIL0iIuuN1ih4Q/EAJB7mZWwC
HEJIDFuGiXJeCohfElBahbM4OSz6dMGSb+jZaJEGym04pJP2pNrUQ4IvCviyO2Y9PVz6GaeAix/i
0aCObCP3XioBN2JOqea/VKbWi2UWgSidGa+LCbS9rqPCzokXGFPEexR37dPKLRG4Rd73y4Yp5CX0
XHw51gmYREwy6O81xU92UxoWbsNXSfGZS8UTAhHGp9V7vcmu7h5daxJMgkZo0M/Zf7bnfVIRp96t
1tnZksiycoVi2JuCxeLInNPRQOJ3I9qr5P1Z9MwGrbEpsa6UiD570xz2Xb77Rdz5At5pjbZRKO1x
GXbLtuMkQVSXAsGmspBn5H1ltBLRJIIF2fkw1yLCLuhF0lR9c3TwMFLRd0vNEJBGgOXnhhwtlS0E
GjIzn4w9IJ54C+lIc4v0reCDN5dJGwnEzTcWZMESXr0qQv27PMb9Fs6Bly2xdxejFBC4pmyrA1RW
H+AnC5I8UYFKNso56TrNGN+OqDWLTaa59creWIchJaTMueuB1kxPJR8uykayDpoERH7+xeV53qsS
5gy0gRGA9CD+Xdff6i5ddqT9nTvf0Vf6HpWpu69n0ApwhF3xYFfAITh6nqdQntFyHDJ3rPVapWw1
zFiGkysdNEbQKpfVKpWKD1wh7dfHVL74BAcPJ0+WwOhQbjkEQR892f0q8PxMbbTgOqQuVN71VXmf
f1aYDXHbYLx1jsjumB/hHl3JGajMcMSpMBulr/5ObNquGva7fxzT70p6NYOg2UWbmBr1vfDIZWCD
pH6fvKFm5f2oLT883b/N8J8p+tm+3BU/ALHQjo+RAj07zrfbc+bl3KqpPP6U6kpsGEIreSzRSGH6
LDv2PBb8NspmlGnzKOnNKhftnqKLwheJAph4UOWim1+C45bHUDHkU3NCwmPOs6Qey3MV1RzFfTjO
aalzVKdBr2ag0q1a82xgtI3Cv2ITbBWzN9DRUdBPZjAx1E4sy54nbWhVvcQ6/LJwSJbILHAzj71/
IPXrbvFChARaPTgRqUKN0c4y7VJ3s7KhK8TFRBp0lyY/TYSdF1TDCStZXhNhcnERRB2IL3MBYZyk
GbDXFV2MDjH35rHXITL6EHOXZaX/e5aePI6Fgtt6RdeuMkR1r5Nh31WJWHw2YgIW9NoisE/oc9b3
VaNnxKIUVrA1JKKpDjjPaUYT/bkE2H8+IadKn59tN9SrfVrSyClTEXqLqzOWuVBm61YRN1A9UI47
CPb4fH7SrSAc63tkh/wgSSAhAXpblQEgEZYZFpmaDmUZbr6w4wlDHyO+uepcnN6vD6VShK/vuIOh
TVpGbg1VhvzkpXnE2Te/7TgivQMMW+Sn9EWXjUIwpuF8tAO1uYhSjRxB3HdbT1fugmGosBWixqkw
qoyBpVVQ6Em6FykNjK1uK7wqvEQFZc0YMDktQqSiDUGyQuuKpGnMeFdFDQWZOI05fxclnGSWcEcs
cTn86BxfuCGIJWkg/MwoP/0i4ptkeS5xeFhcp9XOQcOD1pkYVqrbF79SZCopfbvSYib9KYBH0O7F
ZR2LPa/rax2uXL/m63eUVJeXo2anQKTajSw9bXXQKPG7EqVYFLZkGn05g1Hq1WtnTH+ov9uG7WA1
X893Ayz1CvNT4Nvh/jaJESarTRO9srYZhwraqRInY5dk4KNK0Mt1vQjaU7j1cTckAlBZpSB4tr5R
VA//tPMecHyIyGFaIN0nGBn5Q/Hpe3Ek3cziDngLUoEu9W8xN4Txx3630o3qF4i/VGvL+GYz8jKy
eEZKL/BupZnE49sVpNkLqfats+E6eMhhRhjU+Ux4dqbBz0xb69KDQa5taaHS1FXOt2LB9ug6Hoih
l61s/FsAiHPNGJ2G/jTBdzDYbA5KOmZNh/YB02d6h1yj6kZzP2xKYcpC4RWrSO45bdT82U2nt+gP
o8Kcs00Rj0kvWQACZPfx0KA74AwPRc+rS89FN+ZjLzXZDPjyTVJhfWtE+R2bsfZYVfLX9HvgzClg
xB5tcfB566a1K5LJYvJd9DRuU1qlhev9RGzbT6jzZWsSRruAnQoOgFEFVz5EX4MVSXpCU9AaDE6R
Iv1+/OT4t0mfftsxm6h/45a8623WLhJESDzjd5x7JLesg7anWH034j/h7anA0InxTzfnpciqVsxB
TkH5mo4ySpFZMDyardnQJfYu5bHNKoxGS3Z5It12xZtMN2x/L4Fmir+oxtNUJfi8rnQIifi3+cpt
BOAc+hfwetak6EFZdSXcWV5EdEgzqLpdtYJrogscgmT/nltTUxKX8p2Cb29FbmHSAIzoo1AwokGs
d9WlsIiJ/sPYJTlkNP7kbJ/Ger+bje7nNSBXDV9g1YhezWU989kAIHoArJveVHyh7eBB/INmrus/
svPIxQ56MzKD8fB//Qa/DD704Oo9qJT9rr+KqegJkoKZuWgarRtvAMuU6T7s/eg4ziKLBiZxRZJ1
62YT5VdHHxDBlN32ntzQfRp9250BnUn1aiLChAmvWoxGXRvveOYBrjOt7pDcqvb9cOgrUUg7XN2t
q1bzRHUMoarm/5NO5dv0U1qyNpsZW41QuDWWteLIiMUJijifzcBD1CAhJtOFhsJpUJ6kQNT+2TUY
IaBJToBf973a11Yq9GvENPfOjJaVBcF2xh4HYcVrmj5sP5Nvm9xtr9dBj3cHGyZGJa9c9hkzvWIk
aJQeVLu3tZIJuik3Z1o22Ni0p+08XLsdVlkBMrqVOvNzrDSlC74NNQV5QkF9tzBB3iTjVolrSion
aI1kezE2cd3rPYu1dhCf+w1amT+WWBZ2mdWIgadEv2GuS0vaYijWN3HOldIr67hE6HwaDtAH4UfU
aAtmWgrLa/rTzU9hJRaWumkSje+Gvu7GS208rM72x6rbhk0XzQ/t7m9rc23zWEPb4+ygfq1TdNe6
ERCnfeOBUmqEeXgXVsHwP7bUB/UcYMBHraBtSaleZtzlv+ekdxGStGoa0rINu0KO0PTcnFMesGpI
eOK0z/kwKh9PO/kkihWPW3qiRaHERAmtzO0agzVnQjLr9TjOd2+fN8rsOK9UKsoF3WcylBULV+7v
OPQK4yhkU5RTsKKLDaMz/jzsvLl78UoLdjQdOis0rLUhCoem2JNbttr14LwCajrqsiCLrHOXDGR+
xmxfXm5jTTyV+5AA18F8VGd0rhCWiXqiJR6qxndHfdRfHeFQ7X97G1zcK60XuOVGLtf0hyNFewnG
NiqBYHzZcONTxQLP78wU/RAKrnojZEWh8kY+r3gyU0lWxThbMINgj1tDY8sAs7cPnO646FdooV3F
1EthpRQH0h5Zs4DBJMDJrWnONwg4erQuPsvUfRT1eSVb5b5yUlZg1ZxbVJewTXYt9OB8XvN+xe/W
UYOtMoih+mzdoC6flBqYFBzxqygUBzdZxES5bFrQOMxupc3QW9HJ0tehCLMp59Oq2AwuXWgNaRv2
42XWmIBsKOd1k5tJ0oiqEPJPa7XXQUmHrY9RC5kW1AXLZqw763WQYhLJ3Y0ZI46Oi9liQ3WGxktS
BZPMVDtxhhyVxaOp/gcR2/+y/N2Rp925j2Yaa7u5WXEZ3MK+8q3ISGpjyBJyw2CPu7p/E8Zr+SjM
yNNY3H6YzPKIIiDzkcq7S1okVxgakEzW2rKWHzUbZkuOaDErTF3+DRHcdOz3uFkd55i2+aivhKkf
Rs4giUAOu3fcLCCNgDoY1c31T20FDq3qQMM/cibI35VZvVbsMyDKkTpZRNxHq1ur8KKvpV44D78o
J9NQzfqY/R3+Qylo+IdZF6VIl59ctkwHEFMdHz5CX9UW3o87JFfnEBzAP65EOankw/YUIfSLhrpb
v19jmsHZDNx3yfOdu5esELz9hUsrHZZtQRIKBSyf4ypLmZUel+GDZCUE/WqdgbHLFemqgXb3qa2/
j3Pa8Zqbd/TUDr7bkg8lYFHDNMT37uW0NC1HePZPdD/mDCvL6J8CTZHVku6YCCIQXyGwOOhayQow
sLz7NmAgonmn6mRlckdrRKyzHbr9tr8lucqSESaSIrYxPYXiKs1Jvq5X1a3u1nVGoEtcGkk+h1uo
k7fthE14xS0uC40ikLJUgDE2CPQ4ka+RZsoiUZBpUFqAPZ4/oNxu/NBKbx04kEtaUYLqrb2sUS2i
1jBL/09aBrKvDg4qpMcE0N6qL/zmnXKncnPnIkQHEcELW3m2JCattr8hq4dB7//uLvRswd+S6g70
ZUnJ5096/TvbZ2uqaadMwYODnfHyx0Cww5AxbrVDFc8fi47d2bsNN1dzh4dibEhMvXyWs3jwVEtn
9ZxH9w1ocmH1V9TLBBfGUj6D4y17YF1K9VAFTPGgs8Tl5ffahqNV7tyanlmRMEOKrSZNBgSyDFLZ
OayCqeB/44s96h8o4oPwiUcwEImnRQ/wMTiWeGIaE5zuana92KrKvBRVEu0I2d2rod2MoXCc1tBF
Kg6qQQHmVB8CxXx8QkQAa4tY0w2W/+muY9NexeauzcKs8/88uSG0AWfTH0b5zfXIAt09IbuXIkg8
V5JQt0c5CnyPMg6m/MK5wrLcK05o2rDcOENTH6VKku9bA9hv4/JGfx7DC0llwDV6c81vthshLnBI
brL1UYfdcwSyhgJSTTk0lA/63Dgq5kh/pr8n3XnhP9YGhYZtqTGpC11lufwP16Tsb8nG/YdRfPI/
bCuEGWOp5vUcQjF69Cu7udzFQLjuDb6nTr+/kOw90/qz6Yr8aqpxQ0XNQm0m4dIXY6KDnXfTYhve
gQsUv3+RZSfpagBK7sSU3jT8dUzHeBY+nC1S7KQSzU7LBi+kmEFT7SZkQUA5I5wM2DR1Lo32/GdH
HTxFtOr3BwR2QcanfWUQ6TQqBZj3eRpZ5GmT5pSn8g/NEtCurM8t44blv3NlggAXprx/8X7XFQ7A
n4V/TMitc3i5ywDxnIuI2VFv0Osz7I9p4MWQELTYJTyMnn60+OHL5cdaYuCLUVZ1us6ccCBCyf+L
HnBup/+1RT7JOGNS+D58t04dRqK1siRLYbaOh559cHWv865nTan4ps+c+lF9ddAkxkNjOOhV8Uhe
1CwRVZduAgLwa5hcKtaGDjUWJcSD3jYaiqYqnz/po83+q2kh2ARP8Xi3hosxvVX/n150OJ8rZ3fa
ixq65HeyvegPCjhLUY87tSNU8VTjlbBKhu5KgkNilbDhlz2he5TYJj8R/AqCO8dMEU+QFbWe7Mgc
7RIhTK6CJJMwbs6OPniqmCcGScb9Jj9dMZMMH0pcunTNOYXRJQGQusdleKjw5eNFlUgoPgDE6lDp
vMsHgZHDdjO3j3NYP6ARNu2CBQbS9g1BdGl0HF1WZiqhgIWuE1AnWP2uZqpsxx/vVsL/19w+jLaZ
hplrJEpD+m9V29/K7dZTFPVOaJFTopOdDpfqsO5F9rdFh+5wwV3dFvoXlbRPn8VrqbeH6tY1odA4
DUIlFn6oQOZ4/T+/zNqidyLTTVg8o82Djp8aHrdzRDkIx2XgJDuEe8tzV2ufb9OD5zYbUC2OZuDr
YbWXhKxQK4Jz0lsOP1TM5DLEk1Js1n7IPtEcdocZdxzRlfA9c32CKD6mFSqScGunL7ic7cgxKM33
NkghJRjxhKmaZxYqIQ1lVgcXzpLKKWxCvz1XnGrBE/I/4wKj+6SE0wtHjEq/DYrfR2x2y4OgmNRL
h+ftum+XSjs2f12HOUOR3Mh2MSXSb3fGEnQdxgAJo0LN4mts3OiTOMAwDFv0ovFNOWsVDughIS1i
KeR9ubX88R7ZbY0B5c74RtS/grEmRXkkJDLWst0CVC1V/XIaG598ZJFzaVgHOyaVTUsjGUhNPcL+
gEV5mkp4fHBv4McP4iaJ6Akz3oP2cu6JQ66ErwaaFayyHmUIksIGtGx2Hgf9eyWiZa+qdmnyrMwN
zXQ5NNklijOSn5hQZWI2P8UwB72hH1KXIZLRwNBI3a2Q7malLXWJWry2bALQkYR3tmpnCH+KU4/U
OyGSsY032O0+fJj/InipPVU+cG7U5Qsqtl6EBhWwasWdgq0PyR2SezHGuaXgxcwr4MZuuf5qFIQK
lbP11f5qFnpRKHkMtEHgKnPetbqri0haRAOPm+WDLhMose1bzSX/uGAXe0qUVUvp8Tl52Fv2K4LI
+gkID0vFb7MCvTiWdLtebX1yj3VDshLQneK0zDht3NKGuwGAPyjOHEw8tBwlpiLvaCih8Pk1TFyf
6bRPcMCTwbhbGckCqXIz/8D9eJUuJDhR3P8aZN53XvodI9drBtCHD6gixL1oGg1AFc4koGt38OCV
sEWZjTi6vkd2meJ4uzuOwBGl7Itj9WuvLdnr8kl6r+DrdkbeB4pdNNf9OOomDjE2cdRCUV5xIcl/
ay921xVUiavJdvRLEndLofy4r66N2V7CHOC9P1V8KoGf7zpGIsAbcm5JefcjMSDz3VNHe8RXEGFY
lt9sA+cFdYB0ATsKgiIsee70lEwAmPpvQMVFLKj0KSITbgnWU768eXWsCdA126uKPO+SgMoDda7t
O+x2yvWBybEUJ4nEeozYKaxYW/bBdCMkZOwlNmybL0VJTIsXohhmDTfbagjHuxKydFOP2eBwV7Uj
pbpVAK/otReF62RrjEPqaMgg8VvJ2fL+27oTL9Ln1J4tsTnZh/qp8YdK43Qsm8h68j7mbdTpCzEh
6F6YOrvqMrMteoI2V7Q0LN6WyQGlL7q6NuKi+bth5eqRH5tVqOYS1HABjETVCMi0qDYS6Pe3eLCt
U+s01d7eBN2C+VXRSqzjbSTRU6IxKB1L+SAOrzte4lf8WBdtNcUMnShl+w8oxwM8XQRwmQaRHhn6
L2Q00jboyVt/VWdNpMJxq7cGwuoaayNDVQ825qZ4PhRsgZbJAj/FTMsZ+dsFG1TmT7lmQ/r2bRTn
mHOSx8q8w1AohQJujKZERehdZDe2uNurqHlRpMzM5uUmKTYFd94ZXglRXBkh/QfobCF3qf6hVTxp
ZUjK4rUhf8PqiTjzTC4Dt2UK7rLCpJHO4HW/9sftRgyo6OosR6UlaHS61PLRu3CnT5RIuhcF8pRF
JzVmP7XDEOzsJS/klHX6V2snT9htwCQnozVvOIyGHKVYNyv9DgtaEbJ6qmq0OpOTZ9BkozvxquAN
y0Hn7zjkTbXoAI/UFA5e9vrjKiD9OafpL0U0uu3F7mtg819+nQAWmZzraIhIjFAwpps5MigDxTdb
jSV3ewx+M7eSa5DTRrAWhU7awWt+C+OWzU+uZgLFlvjU//+6umIiXE1GHalZ1JsfoaKolHd4Rhqy
FUbTapDqVdS2H+R2YdXNZ64kiqRpvY1fdTGH+lpf3w67MDX8BMrHVWYr6BFEdXyWMHqoB7PQf0Zo
liaVwwI664795/KVbAl7zg3BS0hy4MkRJxH8l+EUUo+VfDIY36w5cTXawopSmMmcBbsqdwb7WJrr
TEYXY0htmwh9O+G+Cx5fyVWpjv7nJeA8mvKL0towajGoDeHRgiZNTY84DAitmXmCvcOcdDojzry7
Q5MgsTIaXfyLP/WnkNhpvgGAkyYKSEtybmSpxYwvYYxcUUntCBtR5MGF0OBxhZy6onNLUhH2KhM5
Y5rj4OATlOR3WrQeDa3OFUmaU9Qo1jBrvWwqK8jDq8wJrbjhLwjM8v2DzztdlsF3zcffyLOsj/tI
QqfKa/t+C8obrA7mIMEp/EgL2KMbhJG+rg+Md9hEV3rHRTve2j4xLFgFTur/sPe1UGfVrS4yOm+M
2N2SesnJLPpEgSVrJqvGjht509vHQiNdDrjULzosYdjnTjdoDhmK3XAyaD2uCwh+FPJdc21cxscI
s4mFnAfiTf0Lck2o/STy1OAZMNvT7RVcnA/B2FfMAopfZpjlhuu6tl/RkXupe0Ys/D8w9BmYhuEP
2r53zB6Fwm4AgIfzC8ZkyT/kbMTVkQsgSuCDnsrncybEY+jrm8dfylUHqCMTbmxnNSZa1Gti0Qef
KgjDPmt5vHhz0ezzkfxl1adZRSL1VOauZ0pDbwY7NvcRNohxx0cdXMZCzMYXeiWgt0cEVFrT9Mr9
cRnUoXI6lyc1MQJ1N+VtSbDHQX4DzpEnpRy1jHd41r9nzBxtu0aFYuKCEG7SlO69k03mBlgodA7o
oUtHJVvKrt1iUZxF+5AVeKTy5IDwQuvwujT/Wos8G/P33FHz6luwZmKhYcFSO4SSRtZdOQXEzTEx
+LaZxrbuMl9iE+U4kjXTLLyr6fVpQOjwky5UD8YuWH8kpRfE8CEmCLxyLyhHnxJdOXIhyyyYH6NJ
YEYMwgyhlSUFWAy9PEo5glK+Hz5/ZLcwIMt+35Rvc6BRzWzchVTQKunR+KJyOHh35G4/BSaA0uNB
KkaGSn7TPi3tuEjDStLYhLakopu71XNnNIpnThOIyAGLHVAks6C/EXvJGFJE3DthZRneBgpE2JBY
xUdVhxXgsT4ViD21MdtSuoV4EJr5LekdEXpfy92O6oiv548GLluZLOmFyRPJlHt5fDlKd+BSMt14
pbkOb0gml9N0NtykBZBrQgfljp1s2Lr1qzSt05eyyk+m/JG5m5P6KMB5ZkSfeg0C/nzJd4OFzYiT
QiV6okoPlq3YLnrcHFGs7OKzclpN1Al/M7SAbs2qloPvVgmRT1nRCJka8Qpj+sYBcfnIISJoWTJj
Uy4ROX4SxvrEj/CKZjNmjhbXUH82NZ3rbldpP8SI7vMT965esS3urZIyCq6/Yhy6ush7B5phPrrk
hQErhECY3m5RqblwhnCT0LIsRYpzqhqyVWVPRK6JTFF1V/yxm0N4X0F/cRAv8wuNlcOMs13WS7JG
+yS0JvZOnaWWUyMqdYePaSwjKRDGQugeyQxFIXL7shlCGA3/TRX+TjJ7Ckg9SJvfv1WyTxuIJny+
sLyh5wwR1TgrikGGyea+MdaWtHbuEQjItyBIV7mMyJz//4kY0fYX20AG+AD9ZFHFl3xErKQsHsV6
P9aMs3bitWtjQWuX48WK/Qm/ZWZEabD2wnUzSkONZDAPFh75HSSdXYvBxKN0VQI4KeXTnU+irEaw
w+kcHcBNXpT2fhh/Rc2P/iqHmUdO7GGS9EwQagdUSpiUU4/A1q8UPguGUA5SbaSjBbTx7L9hyXYT
N7R8pIEH/hB02BXvYnjU/D8+r/xbOEer33+hP5wog2s01aqkt6GzHlkHk0GWlvKApPuz/bdurIxu
3saSaBsxEBYBdiKLY7TrI5BhPXVlUGoc9EGfV5NIPIQNHrf1BuKzU+uZ+2SZWM1ATW6BpJCXWtH2
wLVXVPV91rQ+zEEbNgVUt1VsYmIjwRNlM8L8E0YWrPQuJtdfLayyyYynxAHKiaUCcoxfAzxOejXI
+IzST+IsQSPKmp5Bb0V1aVslGygEXt3Nerunarl+Lphu+hghFyZ9SA49j26E/p8+mq/AE6KD3+BV
hQRd8sKWciGC6i43Clv6SWncfqOpdO1Qf+1DpykPsKFFAFIwkTIkFgnocqX0oCzK61s4oMx9cocb
avKWKbvWrdZLZkxijJ6BSbrQQZml54A1IHAVoJg0XOCXyum1ul8fjrWOrP8bK0BRtpPh4E4ngnyh
MuGOWK6i2gF5fC2fwgEtHIvGmBvMfhXZKD275yXO+d52XwU0pWZK/dk3a7nRwyFBxARYwvdp9P4P
4pfzh4FNFJ84xNR3E3/glxdfkzCoz4JCO0n63CwPjmzUbuXYlMhAGhtq5cNDz+ePMlB//vu+1Jhb
1C55adIHHWFv1WM4Jq8/GqospocXpCgK9isbN+x+ywZsKD//AgvoW6YKQ+vfwnx6W8Bqwh713ns+
oR2bn6h+MqYdQirN2kOX+hy4ZyltILDURpHwxGbyslPfTm0JmNxLNc/Y2reSZsF74kvTiQA/9pfY
2N7ppqMLzzdDBb8V4tzGByH+glogWPOdx2rdOu+rjdvrs76BPpEHa2gPVGJ1fE/XisxdwtstBeZb
SuuzyKusIVo+bhfA2PQ4/J/VmBfDh3p+nFfQvwA+gfTz1XQ9q0U/iaEwIbnExcBKF8rJKrMwfnE6
IDSq7dy0RCnfZvnWg+jG3QTASn2mImxGMAealn8LsIhLMbVfPGFEnsPymITJob+Vpful9IDtrmTp
g5AZW2aC9ElOcE6/d9RrZvkLAaZEpChZl0tUQys6ztysQ72ESByJ2Lv2RqIsknO/MWamOHeZ3ooO
viuwA/iUtJ75PqVEeYm9AsEFK86vk6cwL7OB47rROlXfd5bdhirkdIwXrxeWlUBW3aTc1WRobwDm
plHSNhQ0NDa8n/CpddrkGS10pHeHf9YkrkcIuQmj0q56e54mYXeziqYvVhItAf1gW3uAyL6YtrHV
5fVNC29wFx3dFpgtcZh7OgiUezefhYmiu36d9FcH1ff9FZTyaR3yVbSfWa5M5UiaoKeJdywLXUDd
hiYa3EOPl3anj/4A5F9fYd3/KWYXVSweNeBe2QeKy5IA0klxIekpjwnVZPGhoZtx+Q0mXI1DrZgi
yiUXVSKw5XVvAo1O7x8sGIj83rPKN6dDCwu1eG3ytiycZnA1mTAGonCPi5mSOkzGHGQih7YN2YmM
xgCHSQjDdi3PHuPOFWbeZp8stWgLv4TZBIojXVFByJebBOWxeJi0XOploEV3gqmoCYai49XbIscY
MEHC5/+Tjy2xX1XamVldWyMtsvhUInWSXwrCa3ZGPt9ZLo5xRepH9wwZkMtuDWO5AiAU9Szc4fF9
Bh0+mRgnH+kXmcAiAjSXxayjmAfE7ibZeZPfy8XCZ0nDI7KThpPRGoR10L3OCy5hZaPdLjxb5GI8
wut2WPVQGQ594mfUPZxZhtFsVI64yUerYKTCT9660QwkhYWGYvGvqt/NX6IA1P+yL4DJUWsOm74V
9cCrUHs7Ap4lfB0a0Q+gKwinFt8xh4ww3nYB2NF7PSAHDJlvQQHdQHz7kzeFt9P2Xiemc+gBLi6H
xyxlC0JOB9v9hgs1yOtRZ/57pwGXuTqvdB5h24b/sF5IEYOkLS/zBIRhyMBqcS3+qq/M/hkfJyme
83C0Fe/wYk6J0A4zGHpkuJnCAKNQLu+VvEeqAPMN1usfEmp48gPPfC/YUg19Clebj/qbKMNJ7e/d
4wfsdNNdHLJsMXYaewFQS3aaHAxeinL/iARopvWyz94U6mxGG1jtWYLbr9KoHp11xaK8MzMg5AOt
IhRQ0uxxky8IaLMM356RjihEqhypLyaQtmeDo8LPkWHrgnisGewSNLd8Eh89KzrxwgxS1REkaWFa
peqZkD4ktzftqy2KN6/7MS5K+bzsGR6NvYqVL/527Py+i4tS1Sn25tncx7bmaBe2p4IzJvCKJ/mO
u56faW6MKn7JZ4Ir1qHwx9+wKqw8VKycDPNb7+KdTmC04rT6c63DKYpqzq3ueJQuJOzonSB4OpNG
QlkbdSOY5Ls8nNVlfJcQ33U6aTCLrh9usex5JNf5MfTJ3DeBGxu9B2bpYFuUDnsiI9xARH4xj8/s
6vG06GFeDN2S3UepShH2gZbjdaAHx9rTyVhhkQLXBtKpqVJhsN7gLqvsmd+6q2G1mVT/+csob/UU
wUjBuTR7RwbUcnPwrZ7Pg49kbjBGbVL/g7vFWdovMbXu6p5+gBAspgQwM1rnSL9gU13mr/TDBFlB
1znDc3hM20rq8QOUvQZk1AM/ZkwM2gLdbMN0EZ7S7a5LvvA7qHKDhhXsmBpXgnD61sRJlItTb+EK
0cX9w7DdIBUw29vxPJ2cHI2w/p05qk5G+MgAytdfgSnKXE4PPfWr51rB+aKG+3f9UwH1D8BKvuxU
cC1RlnfVTZ6ynh23570vILnTaKpQw2gtCzUO8HmXTwXzM3gmnJF5U0XIP2m+34gUjFxQ9T3cZ4wQ
aS41N0MkRvCve/3+UWs/vyi1VUX43yxeWH4DkfS2AREEqyJ43YkXIwdTrAMtqFy7C8gvQExo6yzk
Iok3jEPWu0vi4WOOXMwvk6Lzz5WPldoBsxPlf0sp68FiVIk6+X9ZkqLAKwXVZuJfZbCLchTizoKb
J4uyJ3IPC++FZStpnxxbXOLVtaghLeb6Szi8mEPWyW/pk1fvWzE7JieK8jbrap629vSRqCMHOBDj
NxOmWx8L1VBRcPlm10vDbehS3gT6F/9qp+AkMyAfrSriFZ1O41NhpFxpuvQLXbNxsNPi9CFRv09x
SOB7ih65RqKQMW6pi123xgLQfvKQDPAI91i7NUI/WHgRdN63O7hpDScJtnelFfnaDPh/FAobKyu8
cnDxDa9skYNzjIuuTPK9d/CTnay6crr4cVsLwUphUlt9DEamVIgv7+qVhbLuv4mGlWuJ3llF9MKH
KyWauc5bFDf9sfA8lVQOBGoyiG2ikhlcexGrGmavMIOIDoGRQrP/9qA3jTWnFgKI8mUlfHe4eJW7
BVCwPLPTn5AaxIur0B7+Q6AK1VriED3c70sS8geKS+QerFcEh08aWO4wvTj5SsKuH40NIvgWqutG
VmR92YczVRhFpzLbb4OxzUkxhIVJE41n0sCodbVj20kHq/0jTUtHHacMS2MrkuBRI+pKGeIp8tf0
kC/j69dG+uLAP0vox23nBwn4TcFTe5gciNhDo5O5dcZWyTqEy/1dpum4HJZ4i3kCgAWHoaUCAY0u
aweWsDsWrSrWZWM2bcMo1Y072M1kqczD/YclL6me/xx/nJ0CSMkfFQq4OduhImTtlnbdQ5I7VXun
1Cxr++Hsk/Sg7sbns6qrU6iqOqj1kCSsy1oceac0QYWfQjxa19yrHhZ3z1Zb++2H9+bc+GF9yPjV
bmxX/j5/2d/to5zqTYn12tjJ2JyuD0pna7QasJh5kCPTv27zc7PFl2bt0T0Zopk2fHg9ymcTZSZX
F8HIUmz5dtPH2Pi0se5ey++kWQC1N2XLLXuuX3czSz5mbVOxQdsYlG0dsNGXMmJPqVC755MWL/xV
XHYtCG96rczFrVjVL9lpRF+Rt2cSlu8gfFGg4Hp2gu4SlgmcCvXIDOdcvW53LkIep9Qhm6vvtBM6
d1vFm6eshO0GvbqLrDXvjL6LnBFLL6UJVHniB4q7/heL3vbjiN8Y0Kp0loyATlBQusfz4vijXcj8
DqCNPwIUfxW8SHZIPEr1kqaUSeqlC2j1elOiugGSuD4tQRZ86nUM9LNgj/Q1klqYB9fM8qqR/Vjp
rshzXNvcieeXBhJa/htDqyXxnsAA9DLi8uDvRe8KCOW6ZM2r5tlydyJBWplQ5ttU8oHoKNxYP0jP
MvsV4Sf3Fh+r3HginfuGaI1qZGFmxOGf4AbhiP9PjqyNJC1+ind+Z3ENytN6VcbWQmmKke9Fcogq
wYm/DHLGHNNsm1eLSJsSa916Wmg9dtMv5eHMlxvoeDNhWRcCZUnRST401jtB6jf+h8ne/70kcgZ0
Mj8tw5mY37QTlJYhQX9NKPjh8VActvWc6yn5kBPQzfmfRdyPEAw6G8jQMke30oiFslJ2ptK69Cm/
XK/54vq/xib1lIwQncMt04dLEBYrghaTX71RuePmna8ceCo2dQLGqzjc6WyjWyGzCig73oVjeGmJ
UxjafhH9y+HPf4iaiUmMDIUu5VVf/svBClmZufNO0hlpiMNtmEptX3zmLMNZCNhWKtrodI8xZXGw
+s4vbG9aTO2MBga6Pg4vC4qFOzJa7yc9bQTJIvZZh84df4cpm9C2yQZvjOY+bz81YYpFTyJlmel9
XL5pEX9tkwtnw8+WGZWwp3yjlBlmRd10n+010g0oSyq1FZwFo0xwp/dm3j5BHntHCj1XZzPHhtIz
6DiILQ+nXUKXv6Ie+nyMng2Tbc50NBBXWYQ16npmTiItfDSfLJ9YrVaFJ2OtY2tma4/R7YtJx/Cr
1nCdfX/ZObxiSPr+Y4bOpmhWAymJqDS86pMYSaEVbKaPSb7lwW5BiYV76DorOBvzp/BBZpD2rfDF
oHiaUifVLPZoE81oORFVhHsVDFB2th5rb/AjIwzhPIxmWInkZZ8BtzRhqHzEJQl6Js8uXsvAewaW
+oeLE1jUe9qqmU7Gyoj/AROVSmZTuz7kvorRehUdWLKsJNrU3FN9dPXMJsipLwctj6RnRf1Xea3f
NDrLl7p9k2QCivGPSp6RPwmUtI9nyQ8KXFdMFky+Ri815mLf4KyCjn41rFTBhE1ACJktuWJcIYzx
H12m7qC8aLqgRwC0QUd1DGn55IUcKiJmYqBz2N22E1jd6sjPmU0FL0emb8AgmI0inmr2OzbfJKA9
cRMMkHOi5DghTsSAmHutPbvSf7KvO38rOSnb1iCm8QsNlu3aD0lTBVZhKJAWgOpjf2xGPfcRHgir
TptXaM3/WxIzRNHoh+alQzAfJXolQ0LOzH7l6c0XebHTuOGGUyuykHr3YDkY51yIeK9JXVKauyZ2
m5QpJ2OXVAXbEHLXKG6Hf1uKTIbFZLz/8BwRAtKKknfM6faa9YDsUFu7dkdi6Xh/UmBns6fiKzqs
OCtvdcmF6AIoWzETFZRb5k6q3uhSYmfEwlPFZassHpKPpG3Vhcp6aG77ERGsyRkgjgrCRUFDw8Yt
05zddlZJ16hfqEMPZcGH8m/h6gFxg7zXcSzOVNTLd21V+jPEQorf2xSsZX1L25Cp6zaUySXdRl4j
/+8XSCsf62ZXSf0LZr8Dk4yWaWsIJ1R1Gcl3DOZldxAuwxfpLtvpLqdlJ/zP633fMzU6tJ4TPXVK
MVDKLXhiCG81MSqFqWSnSqFyXn3lStZUcDwRDCV6D6a1ncQOt5pV+Hz0uwg2bgsjbFSMnazM4SNf
YLpfKVNhFQjuH0em5aFxAO03C6rhCsumW3wOofSztMQXVkHa2PUaQC7ZuhZp3Fq0SqIbJRUq8HO4
STX21wlOHwh+G1tgjBPqbKnSnhO9HmHSdXoJJrG1/sNIEftR93kSokOHl0U/EeXFPHi1KPWFcEfM
lhj2cAZ+fjWI18wmyuWMM/op87JHEZbcaFn8D3KHIc0tL6YRGzLtHWNbucGWZvLJs0u+JXMZOPqn
CcEXToWexMtOhBI37f7N+TjRiQ7IZvQLG0sLMWzm7MFH6s+tPSRDBvwXXSyRD4hDdB78NrmBwPj3
MYyZ/BAkezsfgD6I+PolfUcSgc5zPG+pv9vv9xu2hRRaw99R/FbgScYtvLwvfk4J7s6vRvXMi3fq
2DsY2Tq6hVpE4TDxVru4Hq4zNB8Hcu4dW9kzowPU9w8dNCSOztmZb6Pa2zlyfoVdAeg4RRUx2/84
2Cpf59Df42IcNg82LTsBNoRML7kq2V5m17Bvy+L+mjOljyrepcPGZ+LleUR8/Ghtf8IfhRhzygXK
Z3BPHPEqEu3D6DUc7KiS60VtXwvNSanaP/88rdazQ6Ki1yVUE/E9CYfIL+Ib5nUbt/Oduog3q+Sf
Og5wxPvYHD0pSEOu3xA0Wg1R9bLBgHGGIv83kd9A/dCEsZO/xlD4PV5eq640y6aiXX8EwvRP0Aiq
k24k3ij6x0IQqjj6XMu0R7EaEetJ2Rl5V/Ef5NSMVnLTQ7fVUuiBAevXUpMkt1ZH/seLmpnmYjwi
oCfcXUd4r2rByvmdpMEJd1qOSYR2VJSyCDy7NdkwL+xJxAYYK08OZKrS1jZBNGiDZxZ3VaO9fZLi
6N+ZLl2A0NV/sSsGwiE75VdfK9vf1aFm+1yBV/XNFqypl8n6JnyKWAdZmLE30sVxqROVfKUqfcCz
nRe0SC3sJ+eTqpnyhlP7nw+O9Thx9hCfP2sLzKQZFbXUQdC6eeRcX8udEHa7onTE2dzoj1YxFsvH
JKksJXiNIFTdHhQI/680K5Rsw1+KbUUGnPmOPCvFxYsO+MdjUZYtecE4wVulUmkyS31UGtrcGZJZ
T7u44YPjV26sB6nKa6kBLf+AGkG93rwC3wB26lz9R6DIbPT/hBwejz7BqTkaR3D6Fe2u3Lag6SN4
LF7ovn6ff3BpuAE/mgIOBFs67CDjpMzykaIFH9+QECUNOX/zPdQNyiu6yJkNXk8QdqGz9oBhQJe1
dX7/xg4q8SJ9LnhX2fmTZZweni41ad1Eb2mihtq1cFDR+UuUYi5oVRWjjz6nSVpZOiT1KRrzxy9J
XzP1OLLDX1HGPrUOt/udwgOQ3488Mlm7ZNq/kWuLTE9HBbCOZdFXJ6D/hWMYqRtXL3IphhsAOEcQ
kLR2J1RJ1FhAQe09MKvHjeKxolMKPWypUWOYJDfMG7RRLYXdHnBvci9apUP+qiw+LArf4HYoYxyz
mF2XAo25v/tD950XQ5OtNYT/VCLRxDAdIe32yToM7NzQueDyJpEZKfdWSpvNhuJ5/nc2fcYPKJW7
cgtGJnCpkSWFqsrmPhG4dSoqTjJmxpudi5xWDnjNy5CFnTxQPYjrxn0eqMzn+mz/qvrJP0ZDaTzb
x3Sfq0Q8Fx0ynQXsw9N4JAywnrjY8vAHpAb7nUVJNvKlPVE6Pdr51uzolYgJspl6csHq1Z/PcAlA
m2bA7NLOXPbv2TFtPqiNP7TAyKjyXf2IyGbuJYCwVLV8e9kqAQpGjaBzDua0UwCrtP4O15VFMZb1
enj4a9thUEEJsqb8Z8UX6Pybu+t5g9WpHANdIuzVjKifb/XAI20tdoG/84E+0qnmfzjnLOSQ8fg2
a9YA8GyEU1ZLERSGra7Ej6rXm3gHR6WimTkj8/Mk2VgfctqZlSpq1b7wG/ttJc8xbUUNJV9eEBni
k48aoo+j2A0Hrqfu1QO0sU5cCnUB2k7lnMnl9EBSuxEzBgNOZ64qGtlqXt8+XT35uU39/CuWs3Ye
StCAO9VurRSuqama1lAOicEYH8PK8VGjPMxS4VgWmlqt9gjoAoIXNjVXT8jeJ/BEp3qNJ70nUlY1
ofIDFHgub6T46RDBEF8/2OwYTLCdUanHxZh5Ac87GeXi2PgrFvcq237C+mKu13TMwbS7Gl3fK59N
YCUjujsswKeSG18TnUpb99TP9NfOsZE3F6w45DgHH9fAskbif81lpicEJo7jXY+oCh9ukOT5zOin
ikbfBwwonTIULiTltIIIvIeb1NysZNY+eK1VqybQaVkYB7rZThYrCjRwgqtEBzVBS6fV1g32VydI
zNcSan7H+hQEfU5IcIRKVdJwzX7AYbF6kEjsvhfW+ZXLcR6kK9jlAj3dmDdMrlkeATlnuux9lF8S
Bj11u6xRv7lVChtBLJjfPoUvopUx+PsAPPtni8WDAOxFL+TdFw/WqXaSOTIcv2FL+mB/s2xlB/Io
rOcXt1TEYOBrMRJsfMyjaZGUkA6TVarcD8vPH+TEuN7q1QoZ4Fi/IqOyZqZsyLRuJ7881c28h8BP
EfBWvHiMUKFBoWFWXseSN8kKESLGtNcCw8qHrjgfIG+WpzUXDKyhlPZLgxQ1Hlsp904FLjwmxUl1
8Nh+LCSQtUFik1WB/a4cn0o1pqzTCozsCCzehqCTawP8KKlHUSmssbyToIDI9zU886yQp5JRxwIU
ESFhnYC4dVpgFMwS367Jdxd/uEWJgbBn60NyH5RXT+Yv46IA0z5sP0BeMIsp7pPPvcagAJ3+xOyn
vQN5vmWWC8a73ZBb5DPTp1v0zKJrL5LDKjPwg+mjr0NWz8mciktvGnJebAvyetD6Gi77AKjvMmkz
h4NxyTNlkUBOBxijHMNB6sQtWSfA+dD+OiQ1qQy8JeFYjbxF4hUi6UPbMxHCvCkcmR7Wavj0x9Mv
voUHfOmiGhA96FfS3Ov4XXVKN/6Bc5Ne3miKD46GyYc2jyJJhEi3ch2c1O7bK1FrAos0Fsozedm0
945xa+CnySFpvjvY61cNRvc6+eKPCaWcxILegiffqVpWw6Z8mavi0xhpGn2CAohXQnBRjQitrpuK
VCCJb49xh58q68TPlTOd221GLCJibTql7vKBcpq50PChWOHti300Lhnk6RVG6B4HEGF6j20HXPWF
rwBUO5K13jwJC4VKv82FuvXupVERIeHw77weVvEA6eib+yI3/9tw5ZPSO2z/nFcN5jkgZtBx9hSG
rsPrMF7a5hKDRNOWMHhY1Roq51JxVjS74k/dK8jYcD6lLF9ncMmzu18lxKEQ7UJNbV0dnk5Hfs1q
Qj24rt4MPGMzMl+kKReiPTIRi0Jdrm40gJ2TUmUywtWlazyLJFLdVEjxGQLwoJthewAynvmSBneG
u7wWK1tobtbiSjs3CHo5B1xdrKULw0PDOk5bBfmA62BVSfShHvzPh/nyWXuit50cGs92s3T4Z6E4
20TTt6Cngap6TNCA/hpAwAdlwl4POr8MHDHjeJLIx8Zo2bhwKYpeIKb4/88DY5AgwJlSQ67T0Uuv
n0Gx+sKh6XckIq4ndUVNAL4wQLpG/8OyHG4DcjL+iTz26kzib519egGOBg9Jhd3MUGLBjCscYhaV
JrJqS3JKiN9zRrOqnJVzHeUGsqHiTxGoHNEfa53PpzVuWbg2SPv7v5TioMxLn0TXf2WAzzkuQty4
B8DntXOEm2Jns7AVc/h3KwvLiBco1cxc+xQLoyaaMOpsCo/24Kft/z1iYz2btfwgkeDq3H/DaNbY
oNrvJZFZgRb5fS1kOxrf6rXve2GPflwplUsglC/Wo5e4OKN0IQO6LF17jIkEmqdTnsFDGqJHopzQ
xncyC68tOz3/q7YoSTM8vYsJ2fSoBoMDoJN5Y6ndPB+G+uBRlqJxxHnU/n1ON91MTszN1OhQz8p7
pHOdBpN3y3r1O1ONdbtzIaHPPKxt51j0JFMUQTWxL4TpZAGWRdR5GyXtcoLMN3UEmJY88wwFHBzw
HYjjAv0fd7dqNHWZfeO0/RtRf3RAcWaJo/gmV0X+YcP+4G7xjqFI43q10qiXzS+YT0XAACa2d+Z/
vTGsvuQxMYc3HNQLlc3rgPCMLz1OsAPv+JRxyZNbUY+akSXpDh/JqDyQrsJk71lNI2KiLpAjtJ6Q
XdG4mcBUs8yef0bkQdgN/0HLFAFd8/E/qbiBprm9KAPj3i8MSer1MsD369m+2X8SRdqMBxgqO3Hk
VfTys7dW1+NU3+0wr4ZBhqfNmqHLNQCcpE0k/DeyeBahHcOia9bXueHnttmtpF+7MQxw6+9EapZ+
iu3YobYgBTxu3PFTRW4SziFRyDoAPq3eLxte9VvczrlOLYGGHH4cLPT/NKLfrjkRs4QNW4SfSvH/
Gz43lNgOWC8G0n8FoWlsXtoBoCi695mccyJIIWSX6aBgZnNGF3Zr/KO04idGHF9XTR/IxPlCAE/O
H5PKqiuqyfNL5JL4uFz3BREsX3caKGxgfiEGI83QR0TylGHZQGmtwFSq8hYyIQJHh4hFnRl64CnM
L79kbyKCGLxNGvMuh/K5SK3qg4RmF5ld48CpqzLXSKYt0+aQ/QuOjfBUAXd5bEqftZteutECuaBB
tqXJT0XLNoMc1z3z6u1fjxi+8W8EWio7P98LmIuX8NvcxDBux2Ve2QxDEKqOg3u06x1kPAHy/W/X
Km5aEavHqrIQLQ4WhGJqEtEgl7yAW0TMjbz3VuRrWmP4GQMxsFgpp9rJj0IaDAH9zzxHHmDOOOOd
h3tRH9GMlBQhO/nHpL1GaCc7fwH2tkrsWQkLWIYmMzIQfyR8m2fzcMhVU1NTNp9vOfAx8YWcnTi4
p8RV9MB2E4Z9TPxQ6p3X4ta49IJVIdYUT0kMUq4LKqoFCNt70ZNc4FQJvgcus7XjlGTNGT7iNTzo
p/Ir2EuaMFo3/ZTXEQ/nGqiqPCN2cXdHdAhpRoXPLMYh2oLNNJinyboYMupTZwy2V1zibxJJseZG
yOVqHWSY8pBqNlPuGo0Cx0vlR2wDKnbOHquIfSopWSFex2UwN7dg5dtNgD6Ev468+xt23u3WLLbw
lHYTSh3vC/iivR3oj5q3Li7rDYd1EuH/ZyCc+TB4asRwAFhI4MokajiTPrBRIcNk1OOjsnb1ZmlG
0EEQ5i/YYKlV2awUDx51kHfDZl7+79XSHrHpLoeXr2kEb+2Na1lkfKVa8mvOjdJziwHtlzNDvoEh
pa9IokUNzjJtkLs5MWC1HpUaI65UxdN93ZMMeRFV+uJXCu1SYyODwgOVMxcP7+rfnSK6de873KKx
ZQzsFfBnQkVN/whJwPiV6VBEvSpUqnXa+bc1jeTWyEvCbSarUlDDUhBJAFJhzTe6i5+eLRCCeniP
bGUOqLF+GVs4Y6PD2YsUkEwPLZ4S/5Ri8mpkcgD+8kbOJ2YbVkuIb1A1rSpZlvT6mreutXOd70BB
ejU1URIs7vmOEu+65n03brvOU0SVop2yYdFn0Sm14a5TSNhUKQko3NOi/1J+au8v/Wzb7QYoWMZ7
otCz02Ke/jMEbfhBIy6KjkfzxdhCGTYYbkBb8FXLsYD+3yMQt216odhBzJNLlzCBaFMZL65hWKYB
PjXjVqzcTWL57t0Pv9F0Cw/5/cbnMc7Hcc6KZWAeSU+R//u4QzCm0a0wY8t649y4xzuOGRMuzTeQ
2+cVCgfBtj/ezJUeriW0vp3XMa3f6d6qh+/WsHTf+y6M7Nxh9UWItGjZFGfuuCOD3Xxr0MMJ3x50
yDZn1aT6gDuceL/Ft7ZtnvgHjh5zRvAfpKGWK8txEWHR55L7YV+sggCBGCGTPF3ShpTqT+w9OcMP
bqDjcPVY5O2eDj4L2ra4Yl1dcOXBkggMt6f4pPXgolojKSOonN/sHED0bhVvTu+OGgwfjFNvHRlh
IX4EBUNGB5F9M/A3lcSNTkjYQJMyQ98QTycUA5UB2/DxYsQR+4s9eAMAHqTZRNfTlaQc7AQMg+Mg
TeNK2YYj6BGMWZyUOV8fY4CYq1Pp9Y0nW3GB58QrgW9X/98xQZX5CCXYVzTsFhRKqWLU4UL1IOpP
5wCLbNMgQ1nPV+nwDz/s488J6rBOZ7oZ6ErIsQt3ozijUNneTBZjPfkbzfDN41CLozutzZbYwa94
DMWDChIVqn7AJTSzhkYwko14pw9b3BafzyIYdRUo7ynDInZxtb7gKu3XV7qhXSAWQMnT2Khl8wJ7
dpGu4cZky/5IaXqOKKGI3u/WI1QB3Uv71+PWQIGmA5vxhWgBzslcKvxyYvXeCC7lr6KwVyfRCt0P
ITk3CV+ss6d0u1wbXx45o89nTiCYTCnMh/SSRznWlWuCYKjez3NBCSrS5qzmeuFszAp70+wTi99X
qKu/sh4NVuWtp/OveFYHLhDPxStV3UD9TpONjH+KPP77zNtldjq6Hb56J4hTkSzqWSdFyxcKFsxe
IVhaO4oZvo4d68ae1tH2okGDIMvsC9hLF8ot0nZYcreHq/VLMrcU4UP+UNwA3BxkXiXP0dcn+tcr
kPE4RWnLdYNQQ8D0D+8n8d/yUKUIIBksQxgdZtxnxcusR4KWibjM4ZHwg8ulXMqnPTqQTMlFqv2E
iyLuzucXwOnPNDjuADw8HLuj3+pZcZaXQk6yoQJ6OpeEM4fo38RG1exU+zl1SrJU1/uvg6BlfeN2
b8vQbRoOzSFqDtflgclZcwUSO7OwjMLT1HjKygIBz3bjL8UqZuwXO0PfuCIDd2zJ1ZI6QrIaGdfg
V/MnkKR906gFMqD5z5aiou+KCCrpI10JV47uGXIybnNdwOPcu19U6VtU3JKBUvvhLQKIwSFREXhv
+28iFnhqiijTJd4knNDNmmEIMg8fhg0QhFakAfvLSZCj+8UX/fS1Gr7cOLdz71d/09cFArcoZwoJ
hdZ3MGAnS7/SfQhq3fmm7HlscvI95vKkmqxlMprRIDxo1PnpWeme57Z4oYqjho4MQGl3S50+pVmm
wGWmfdVa4dwfhsJKgomzcwKuBs1LpDTey4wHLFGKPbqrkbQw/0WPhtdzn5K/ptXaOiwyLtASo0Qg
S4y6AIkhsc3miRIQyMITV5hea4XzN9DGt0Gg59ti0sVA/8KhCH4xIAZlx3fNUE0/k7ubw507i7wb
JN99U5hiMQGNza/dzOLkpsCnMDKZCaU10JHwlLcAoLbEfbdWu9wVtdFZwrCqKfiVu/WbXjbVOikd
f/Si3Rv2u8N+6wczfR1CoasyJPUriPrAaJuoUfTWDHY7+S5QvPp2qEjWCosy59UYvOeN5Q82bVdf
0RFYzu80l+c8Wil89zCqxVgjNMjgZ1sbau1mhnJneBcB2kQ7aNAwqdwsPO6u9Y1I5rMB0tdzwQ1U
lV9YDcbWnekOpr2B2Jdpy3jQzB+FQ43r30/C3MyvGxxJn3gHhiaFXAygwExDhJpuevBXYbAaHHsK
PxqmJGDgWiqLm5VnyZKHPs4K1H9J0O5atHzaI/ggRcNg5XAvQqeKik9MqZj4EGm5r+GB+IrTdPgR
caV0aprsSGrxadPOzVanK8ZZz2rSFqQ2XB+8dHt80IaBBIBPZRRXLrqeC8nfqIzFb55DzKpUHN3U
sYGiwn2Kc/QXgJRdM0swQ1TM9Rn46HNM6iuz7PIgRHRJgvwXwcOvIveqSdfdhz0iorOTyZievNGN
pcHyMkBZQdQ/w1DGwdL16NMOsZqvv9NubjouVTXcWG0hrNq2O6ZZu/Jt0nZq5AqSdu2myVzQCumA
fuo/DMu60CT6mjB99nyZ/Q2mrloAe55oJao5fhvJTxrApko4ajz6+QmixT3+IEe0975jODN9UGIy
eOc3jFkKBa46Frm8eZqC4WMLZzlCwoMmSZ3j5rLpybGQJN3EJKI2YbzudZ/wv/HHJKYgS41hhfqv
UBc4swm6MnmUR3Bytx0odKUlYS6Nez3YQrOLFingDD4sOZX5pTNRpbUSKPNi2WE1bEI2p1krzW1b
T6zm17CxpYspmMkBteVCrf1gzP0q7j6jUzWpgqAHJWXM1Hh9BftaNvF9en5juM3jm63/x+6AN5dQ
bBhr2A1J/0YDmmmU8keI6YrCxcI8u5QN9aqgGktV7csD93iKziBzwlBhEZ8ZK1C8/ArV75171d2p
4D++lzYOkPWm5FTc4vDL1pp1h/HgiFOKSjPjA3PdTLF0C2vYeIr4q2voIxsarenMaxhuVwxqh/Td
+VfDiiRE0ai5o4sho0LKCMHhXTjhCaccHFEJK0ROmBAA0VINIj+p/WbP2TxgdflvBPDE3Fy+xuN8
6icf4CnDsBeQd+q6kSOfDN53LcUqZlTTXI5L3AAyn6Bff724rXf0O6TOnSjLQeDvSuuM6fNf/Fri
P0w/gWwg/DWVZDVAdH8rUoZPS8BofQIscGrtLbsS/bE73wgqCOYKCa51mNur3WlUg4IM6ApkbPoV
P6O94mvQunyqTveakYFYJsblk0cuzhyN7W6SyXujrTAJC/QEGO4hCniYPTctXF7iaeuql3eG7sK2
FKoujLffhQBD+A1cI6GlIY7ayCIFSEWdWXD9pRQTw4+mJexfC29iWJH5VhDyvwXil0TGLmoPjr8i
J+SNskksbPZol782Wvlj20VYfwVaF7KiS8ZIh4xZ5SAfpAS5xRQwsIjyBAIZ00LF3M86BFgO/gFG
3v81YOXlTiN4QZgIAmTU695DEqUjaBpSlYz5uzQVGH8SbjYaAswNualOCHiQ5i39jbW7Iaq8MwGr
ZadDWREnsUryfpmpDPPQtrqr1DzQJNmswKjLg/El/IpcyGrnVle2hgdHhN5nWgTlhofgcAA/F9Dw
gKR8WkuAEL1pQ2r0ckzj8UwBBYAwvUV2pnFgrsFdNvdvK5uMmDzTXckEEcbaQyfSLzx7361UouvS
xFeLb6erO4VzVGF0ynLKgDZMHojFcl6MKDtyj7ML8sPnVOsWdxTRQ/pheuev5ulRXaJgFJYQbUE7
4NbbrbzPCf/bBo/7XwWtqaFsMq2U3thPiw6QXokOcTkHFic9FPCI+771ecfzKwSzgnOWnJ3lbukw
sd7Kmf3VcOj2bo8s8K4io0+12Llx7uXeeEMPh5j0hC+kaFuu1bQNn1GZxjO58/ReUYiPxCk0/4JG
kKSM2QKKbnwkXTosFisRGZT/xk7JhEHZd7cI70tcy7KhdPvDOSl/2xcpRQOqsBg0StOzAi/fyfka
2DC3wzuaVWjVY8UvuM6HF/AE9Y6Ysjl0PwTzBnzDoDkqCWTksOtCj6nA+GxhsoxXcJARgBE+ZhvB
nS5qqrALQygNVEeVB3qWi3xVrGN6GTA44M/pX7ad89crZmtE0evTaon5DV111OtkU4840ojx050G
ahZSFeuvY2GnpWKE/Fk6F8XTXKhFMlfy7kaepiHnyrSCTKbcDuXgVYbyhES8JpIEE3HwV4UU2Hvn
35nRGV/ktPnpUYsSs8pUF8uV4ITSnA/8MD8YGWaDSOD0K3X0bC35Ns3M6L4Qtmrf9ThV3NRf4y8E
OUtAByVu+dv89PLatm3lMWdqUXb0PWkroidfsodEFi8E3BWyyMMWSu9muhE9IRgxYqtysCYTocU9
e8zzkh8dD83PC7dd9QXQXZjxaeTOLWUUyX3lX7E4YI6rXcjkiglujH/Q8KXNP1G7CBbNApy5gEr8
tYu9QkctSZ5etC+AYYzLtY4mQaWTStokx99f6QKiYPmPf0BOaSmdsLSB4pWePKU05UYVXs56Oa3r
ZL6FLY+6QckMtnxd45CNRyaDxQzVLKaukeWxm2kTRIFjecNiFb8785Bzru7rAyzmTofNlZ/lSeav
U9Nri9bwT5Go53yHm853QCno2ODPkhN4WmQibE6QrD0dXxQoSTBlqaaXl+rTC3CpCFnZ48joQlys
z/KTWSMK/q3kqiiq6FFFPIEJqK/2FEVh337BhQCZlrKBt/kcO5CShLoaksUPYx42065of5r2FXdE
CvztMO4juXqi3oz4mewSnJIj84K0qUcvd+STvDuRBzn0JKBl7GskndVNhjumzNMRkvSEPom2r8Yr
qDmaECPp7WQFWp3XJvVj5BrdC09C8xrfRd/Z9aHBuXiOW2aehvtCT1HSL+xIVlWyGxAIe1Q0Z/J5
K4iJcdRbJJkYTmbiPcOVz3o1T+rFKO6YL+1g66s6s1/RlPv6klEujvTAzTlycun4YMveG2d20VdQ
fzZSBmGKrK4upHRuVH1jJla9mm4hCbZxMZjhDjaoywn2wbkaCdCTwuW5ieNtmBj7j7PdxHcz3WYn
EK8uoDhyxZ1HGY5qNlQO6l0SW1ilncTm+zkpQE6JArz9ZLv7cY8EzNYkmIg0AknhzFYW4yMVtkIm
E4DcrIobUk/yr10b+fkpRiTe1fUqxxnouoS6tjOveWK3rM5Qt0neLdaLRzWdSFMTYOpFVWT4JDT2
xmgk1I/avOMzekCD5MkAtDBFCYYYxsZO4LhnLCaFhZYELW2bFws/p3C+VexPRTgHINGEP1Y0Ovap
zfMktQjLM6+1BHh3wjqtj9mnXN4CV2NpzyEDnBgKvU1isIKEbGD9IPpa+lJNvbU39MT2bF7/T5X6
dTcqrO3vZkkSsQ9hhqrbYUrjsSiT7JyMwEhMqLBimzP3zMMg11fTiw0ahNwlN0huuqvwOvlOV6Zg
6LC5Kc55eLdkNNFx0TAzAZI2cNi9nyoOPmjY7MbqMESqRWH1x9ePwsfH8JnV2my6PNrz+cuDIccP
8JWyr42+snfHUwG/P4CuI773AI2RX2FlAoNL12Z8LOnK8QpNIwgvyIpasWD+2fKPBDUFpdJI/doy
R/ltCI7o1TXBOsvMebSmpuDHjgSnnnHMYXeTLGO8b11H9GxKfaP4M0LL0dDTwECYKBG/6Q//OYr6
/zWSoTABL5znAqFFRZZe6BCrZ9ycO3ul4dddraRRf0V6Of7AvIwEYerMxOAy/WdhgEMEimJuMfbD
u3CgH48p72u5nAnJchhSGdhVQgChREXVbZP0O1atWZJcJ89VOwTHgrhkpPjAe2Hv9M3yYQUmZ2Xu
yIyRUnTQuLW7wEm9kzX/KwFrteDJpX5FtfZgo/9gfcv+v0Z5oaraFAyw/Vo+7IfSg641A06XMnST
nyZGw4vU210no6x4lKb2uMY2rJyaVk8exroyMJZ43QKEcdc/NXEPaVFuMFqQXDrN1+VDUhiRLsTh
rim5hTYUZGm8c+m1UP2SU0v53k0jyN8x0NYwJAAvWgjP0nwyB0ALnR4ECuKM6GsqV3NOvBitJ2UC
ZKqpQaEmrhSjmaUS5+L54ugSWDEWxwpEiuEgSgAwmbCmgqVP+YArDHTZP15OXf0PBOBZ6mVU9q9b
dS4eH7ckvHRdnh80+zpAbLkDWm1BHRHMabNnKjwYOMoohjpNK9q+bxMiiuGAfbDGhYv231QWHbfK
Y0yTUgLkVCAIcb+avgYFEfHYzB1l2DqsGMoGFd/i8YkhTClhGVWpoInCCJ63h8rLnkM6V0b6R/K2
oypz7jKWjXqX6dxW7MH8CQ8m5zORxiILN+j19p8A59JSH5xaRWxbyYXoXjnW3h9ZxAjdJfo7ohdE
jQLklcXx1HYDnjOU2p7erN69DSt7O1q76jgjcqToZeYXUnf7QtRFUEwB0k8+Pbj9RFxMRqJya7Lj
fGAXfkuo7DIBWSuMRTModpUdOzd85gvmOcI1OVL1zkBc1yhmY3EQYaKpXhXi9mgYx3RSTAVLf7XO
OrUgGWVZ+tYN0Nh+vAD1JZyYuxvgo2URfEpKC4L4ZkcZnvGmjlsl+15fXwu/Nm+KevQEz8h4qLOP
0gavF2sq+2mvS368/NYk5/10vLgj/S3tk7811oVVhmjb7i5ITDyKXYIqkmuXH9aJsc1rVte7UnMx
7s5qlLgdrXx3n7JTy1eLr8JOppF1ubb5tKLY8fkWiVQ54zREcpu7lqWVEbFCz4TxHO46GmkGq/kV
CChK0Y+yTCwu8IwFbZyg17js3D2YOhxePsdnl/9I2usElfAJp3jMVZLoEFvXskh0WqL6jJ+RLSu0
7hNyKT04vgFq0bcZ00mzw6ENAWG2QjQ9YIivbEhFZZqn/E1ystan7msbB7wSYiUTrnHCdIIPUSS9
uXethGeNc9Up9LzlY129ECVk1IlRmblg5sYigurN250yyPLKSv7y27+8xMgHM3kjc+B55PUHn/ci
uWpzQh7ECH9TmjO835B1cR8avUWtz/BUEziolfLtP0hopHacTc8BAFUJ7yFMWEAH8Tw501q/u4v3
ClfjDVaQa/si/wEBBCbaK430/3O4sXp+rLrOTr6kUdfIsSZ3McWsFDpqlZnUCUNFosaPPf3v7oa4
dfeBB//C16U5Azo8ND9ADH+nMaROMRmsnAWx+0aVrqxTMCfDRlGCfzli2RE11anxuCdmcsv/yO0d
zpmmYWBeZzR5ep+sw6fkrysF/iQqALGMIajsm5NJVvEO18LdjlrbBDEQpJ35oXTXFDcphwARy+2r
x0My/5jQwOTcfeSF4wEcPfrh5gSX8jQaApIiRDCmFJEp7njQcWKrtC5QP5D7auNMjTi+mLnpDWfu
cy2ClUqlp9AkEUgvDs0QPaXPvBlGgfTqrFv1Px/o2/GLdX2YHf0A7IrGPkHFDY8Ibw8JkJ2AZ+HS
sKHybzAPiQLQZNF5/AwWeF4XFUvKCCp9sEbTu0z1dZCyKwaPcX02XyDLEofMX8WPY4veAqH4AojT
QitXeGDfVIXKPYdgUDmjUUFrKNui+WiKB3h7RkWOysLXz9kKtr2u+xlGbWgw0fp4ELSPpN5thuX7
87dI+IyLnMFLiXiC2OqfZl9LapttqCaKerMfc8GWbDEC0irtCU2fc5s6BlX3QhYfPZxmiSTW9wE9
7o80wwgdwocVxQygH08kO1gl8NjXb+HE+KiXtDFx0DYfyBqFgYYNg7irMHWXKSDAmOSpBnAnruBu
2YZ4YnF7EShTCbCLNbS443THwxFBDXESwGkupt4b2kuBaHLJKby381XqLZgBm6c1kxWYDKKAua/a
my0w5z3mW9r2+EU9ri9Ua4UwpISHdStw7iUbtj476T1s8lXYmEM4ffohbg/Z2A4996mu4UyLcwGC
w9WtI6TRqUtVtU3ecrr9aC7W3jl4dZOJ+FXVmAKWRo2kJXwy4hRWJ1ScwXkjxhsmXaqIVnINLUdI
DZxjrQjOOsUSdNT1zZIklVj3yV9xgPvsu6pLvOs91wG84EUTrcRhXSii7mfV02CbysiunRWXAgiK
ilmAgLESMOLezO7/1HMVdDXGOVZge7ZNwWqCJbbU+dt025DZTsSL7lK/89ilR0EL4w4PAbhLoVOu
YTFsopBIE/gF2AMjY6+xc8QWoDmrG6AXs6K8j2xiOMq5mPfyWVQ6jlJe0stnzp4gyDbtI0XBRuq3
yyD3oHUsI5v8wC25f1Vc0AsyKyuWx2plTAPzHG8PmtvGOidFMLA1w3Y14qSod6snXGRie7gEvS2U
4Q6XM0JKQqZr7QTDWxln6Xv5LyHUrzm7HW/gdEHGqdWJdBYXk3sIRrs11GUFc+LrlrGTBFGcsRHz
v+g+v5SlzQ/gBH4lwPSgB6haRMNOaYO5q/8WnJnjY6YHnImBWQPnu+mER+u9I3biA8mZyjqPU5bo
0hSnhfYodqoPdUPH36AowayJvvWG27osOIkw0Xc2jA+TqEiwwFs/3iBfQcSuoVOOsML6r5ZnoPeL
YofGYsk8ZnY6wqrupGZ+cOdnKxqpPqNb7wO+YXle6ZYEn+EpGweoo3i0vchsvWoLC7Pp1cX1cQIl
EcuDxYQjKgPZk+Jf3t9G8MXtJvvUcy1Echf/JqyDiKHHqJASPdZlmL31/HI6Yj4TesqfE8GpgNdZ
12Q5nRnjqIV3f2cwk8YL1ceO65EwRk25PF5bW+G2TS6i1RihFMu6amrgpPmfRawKVh8fiVzsSuRz
qFEapWVxTBy2ZbvGXGJh2KlA3NOLpABm75M7+y1baURll3Xs1hZTZVWoyN9L7dC6iadKVZgApbAT
pxB9M+HXeR5KnKPFjOtISG36f6pkTRbcNgEpx3c1tQjrUcseWZOHIeilTQeTiEj3Uc2HL9RCgYjO
ho4m/BvfytLnH593KDIDy8/mahk3ESaQSvM7PpGapLKJyyWBilt4NejqfVzHyFbPWF/1N7FhQXej
68KR/Xk1qDLZ8iM9UwHYLbh+ao0YcKH1kL/Lxy6gZ21TnhskAANx9hel36mOSsk+Rt7mUwJo79Zs
bb0eSc32OpruYfSAkciqN9vm4HwqWVXk357uZMo9H7KhgGzGpuFhsDDTIIC1NWYdqSlZH0WKVmDV
O2xfWuntW7eRl1cqhhPNmkbdtZBc6wvG973AKF23hRs118GpiHK4U4DWWfBTpUZivz47ACNYh3mW
6K0rIDGtpPuxFGI3ZOTK668vLBP2kUYb0v/EwkzXhgbMBF1n6ZGAngHM2UvTxn8s5FPEUzrvuWYm
UB9sRDWR9BfuJPhVVebq5GE+Z5Ahihioz4gDTX0/z7jQ7dnBnl9f5Du/FOzRrB6mnt8R6CXglMe4
W/1HLuerd+8GGB5MgFE4RvgzjzPvXI5bkp7S2jLRrjKZbMuQiCnD0yE06YeE6eM9Gu98TZX5JAJ3
XTDEHpz+j9miaA00KtROgjLHBdrvHQYno4hCM80Xsw4bjTIsE1eVcTcu39XnF16es3dW3835y0eb
cSnMKfv6bnJg1g+/NlAqgedf5Uf7axaIicencwD4VopXqcP68siy2vKIZ3RRU3Q+vTSUNymcbIlp
V0K2euG86SjXPl9O8vt8NDiSVhtlRPUT9BuVB5ExydqKfHhluupQ32RDt6Sk22xvj48+bf5un9JQ
uiqUxTcxfKeH5CuNgogmky/vHDqMueCXuHeC4/uhN2xjB8Pk4L9tQKhuDo19Fd1MTAhmik+N/9zZ
QhQ97GBA6IfvizR+NhDQnadl0K8aa+Lj19uvTbss+LxLJFJnpLwAeelotaGzAFk50NNP97PJ3ThL
G+wlVeMmJHMI+cSvFHNGLxZ2WrgBA1MbDzShRkzbUBVveaOJrPLlINMVAscef3VbnbCPmyZEvPEX
mB0DfaCC2cQLptpYSrHS2qgOYxLLR3wO/2Z3Js4WxH/gPx2bHynkqu7+YFibph2A6ruC9gFRePec
sFP1wcC/TMCk1OQgPK4CdAqswsWKHeUWUEdA5VnKhO8U7SzuSoPDKYUgM6w588TtWTRXsrHOhjFN
PWfOzDCayndf3fHB55Gx+FM+SShGV/nKaqxMx1CQayW94WHRHW9yf8P9EpOkJeEh1G3peXLEHK7L
AXGkF7uV22xwqqK31srcErUSO/ruM5Fj2XXZpnIe4yuhfVTN36i4Zr6LwbKQDB4mi6Yb0miEGENT
+1n3GerMj1M3mUxyRS70xpfDmLu1+SPEFeIdAjWm6j+T/dA6FMjnjhQlfXULlRs4L/ypSKGbrCxN
CvrrpFauaFw+gJJ5/J9IYW4Abpo4s+dIZn3A2PYDQGfKIembVeVcT23xB5WwBgtdFt+LlcXM2aol
RR/dfiL65r2oxAaB+wWkITqXJLL770zjMzz7Ae4gWKM+cw5pdRY0FYY62R2P5QMY4Bk5cvuTntQ9
Q8ay2nG7PkXJiDySRiAO5w5xC9NSQL3W2CSecynRJT9oa6C6Jqe87DEz8erXa9LRseC1q9hXoUsW
793VoiANfaBUZGtRMVijVakCXYuSJMORqRh3pFrniYApWNnn47IKELT+3qWWq/XTkeoniS8NvCSF
EYF9P/cL0XXb745RUi7znDc0iiIUTU8mdl6gZLVtzHlWdzQ6yFMBQ8faYQJPK9PIIJuRYNZzbXRW
wIw2qh73B8WEOpxOsTIYzXtgVhN0YLSmYmoH0oBgFqs08yIM9qn8DtjM7PEaD/d+7HFeJr5AEzri
KQkryCPVADMUJ2bFRzC8D19Il3n6VJoouzJdDHTXnkozMFEGUxEbmwEo/O7eGixPfg4iP6FjVxQ5
Wj/o4yhYStZeCmqxzZy6VOysCM3ZVazDqUmQ8KHyd6zYFg3knpg+G0PQcMuIDEq9LLhk3WEkfDzq
6hmaazKU+0xsGRTvUgVTit45ided10SqTb8AqhrKlx9VgvgoY6b66IFEuBRSnjHgcVKWl7kLvBk8
r/e00rBFcUVQouENUQAgMLuyxzLU7JOuO1G/85RBqqKf7CkdXjV35C+JgkkWhfrjBzAMNaK7xWwK
OK33+TSd6RxW85vldPiLivY7g4or8oAdvrcoETeEKzDyK7/HZKtpRO0ao785styAF4CcC/oAaN9t
A9bUKXSqdjgptm/M1Ef1K1Jqd780jGC7ba2pI73DQW/E2cEg8Q9RVh//rsMHABKuICA3WMdm5TBW
J3HJpyCN1I7w04VZTkkVwy6ls8Cc9tN/S9lTIWPGWs3umhkFJ5TwKSWp0tv/M18ku/p/lKV7Rf1h
KcmQWUb/WszWuBKJZLzAJ9ejP2uPvOdTH5XsBCv8jrJ0TZ7oI2f+uuG8MbKwNc8/xd1vK+D0hY8o
ijTX0qj5JJdooTK4NOU6jWv+8UhbHwg5pNpZMwRon8dyOcqlqRKP2byrS4r3mzgAJEZTODljYa2x
jYatbDXhlhnM8ZsNZtqbmPuL/SWq1F82d9EUGzhRHGRz/Yr9u2DFR2U2EdyyTY5dHgvuIy9YPEUn
cwINYerSx4n5AnFV9tVhJA/WiaeIBOMc96HWY2A+HN4aN/AOlsj3mj8oyzB0muZAKdVUKyqTPRwN
klLf25dt4VVA6kseqUrhM+ttCVBFeinGMBtsxDO8GGIyw1s4SR3wzzv0RxEfMwTNERjTS/ID14PR
Br7hUBPmqrgJ3llSN22/XtXlwMspmd5RrP+lCmdTeyfAwpYO9Kl+CUYXTiAT2XlRgo9fsZCu1uKi
a6ZdFEFKGPYgci6xadv/W4fRCHlRrEAl9OaUlWFuTq5bHpTEccX10b8cRpJRjwj+aDvCdIipXds4
igJggXbSvIgRkzKspzdcN6fp4T191JrInVOqqs3eH1+Ksy284vPjjRjOPKoe+Wnuz1ftOBkIuBc0
JCEEGJqdPge642LQQr3GYPJLlBKJe+vmPTBJWDOwconpzrr3vpkcI4j6qLvciQOigcH7o2YbWaby
ZnCD41s3mOzZxb35xAy1tfNm3V5CqTzEtx/qpxAhBbvBWApLXZYkiTg6pTGf4NAaL9zLMTAXMHLv
hExkp74rpc+EF5H7Wfo40g0K2fg9mzG4h3zHlaSRoXwUSwOBgoCY/9IaMn8vmbjQ7MkwzFFKVUAP
8hPFg2NZ2h0o8hy6aU83aIx8sYprhUjLLLwgJlI18CFTPpv7hlNZTDux5VQFceiC6nJcCsRPhwNz
irXhU2IB/7HUw8mI4L/XcmbCeWIZKbjRmaewRN3Gkbox3NzXvxIMKLkXxDJP/hYsMMCWUDHeTmZJ
RH2rnA+U4WtdC41zNe6k6LhKR2OR3MSXHrgW1kstGL/1ud9A4e6rGE/LM2MRiRsXk99+v+EVeihf
Qy/GW/gLRPVqspzl2KGzI5p5yEaI6EnTSMY729bLIun9Gyeldd6nRBL2Oe5mxUBJ3JeDzvLIBIV6
5xtbKs1Krx+ljY+qsyGZC8J+2M+oV9zknd7VVSKONWhR3gpIlxBvGiEmlrYmPvNB3KzyWwBj2aCI
SuPYUe1YQeVQO1f7AeFZIR+y+07vlzUxVKpmrDVWQwF8HfBO8Y+kr1vwX0JTfa5rx021EZ623Sxh
ww7KP6TGu1QzItP9VRHQRvGz7Wo3t3i51Q9Gx2wgzr3t/7ZxrGRSZNErhJeg3A2mBk0BPZoTCijm
WDAsMnaq78gO4jgaptEooMtPYtK7H42o0IT67NEXJ+RQYW11C12DSKZq6FI+5xsPblOOCV4Cp2ks
KKvDuzaGuHoiX5V1nIxRaCMaS2Ko21kibtjnXdXhIDifKDsubz2OLyfzp6BAgAs39ZPXHQykGT4C
/AokAM2xWDZZmnzr1C7a0blVDE6MqqmySM1s/gbwAsm/llRiuO1AGQP4ZUnPKlPamtv7tHBGOzE/
fARBWmi1Ys8+K0PC3jT2vMgV19pt3TMqDfZ41+HmRqaMs5jFzr1WvidNjTUf8v5YSdRbaqNz+ViX
fjT9zgg/q1oTvqaR5M6d63mrnNdhmrur0utCAeDuua7jV4DWj4GU4etn9UTGatr2CtlS7zX6W97u
PdMHkzMuoXmcGRdTRjWmCV6RWUOH/boYb//PUr5Au1iVJ0vthM5c96rCQUEXo+E40lvtGDfL/iBS
fid4SMKYZhFJPWCEb49ZC7ZD0WKW22nByHkNAU9Cp6Ly8AjeEKP7rokmBLyfn3AdrPPXlwnldzJw
Xlkuk7bJujLEVxvLPsgEAm8huqYaPlipQHxWZyvkWBAoIgI/+5emL6fdA164Zk5sE8TUHGY3jfuD
XSrUWxNVsZ5bGmwXgePZW6hjVa6PbTpRpV3pXnlNSs5OeUVuzibBdT5wFpb8iEJBkvhrJ2udeDPj
AT+eROzffEtyMWJyKUGMERCPPLigXCCt9N5rsJWsmkQ/KgoVol/jXEjOM8G7H5wM1zWWNRR4nRir
cqO37omAJvtvpCVY6YXtW/w0BxrOvI4OLP4lPE/9FQA9jmu6Hn/zgGZOK4iiFRwjqXwY8XIYVQbY
NDv8xvUu3NZnLRQrr9IBVwM53XmgMA4E/zdm3NDQ2kNLf/W2Pe337m3LRI5VdVlk0SZsFlFRv6qj
kXayD9q3QJvq8gmMLx84kSRP/H23WTz6GXJd4c0jfFst/KUxIOvYEmh6QbQasuMLJmN8xo4I5i0P
W8y1WrQZNCQnaFNCnudLnRmw20mMKZkWhzmQbMx3m5w2+gdRG7xQ9/cu4if8wr5hjnFTJMbPWI5D
llWzccpzFui9I5cCTdnzl432KLsc/uTPlSfTAsnrOkKpD0EIUmcmp3+o3DX8mtf8TdqwjwFO1876
kFkCwVEC1tYQV81iMbbSt4kb56RO1vhaDoUh4TCNIxn+OfHoL9x2NkDTh2HRiuwnMIbGM38Yc7LX
eptWuVP40YL9FL/ruYsP8HftWTFrnygwse4JLbLAso/g3j5OdG468m6Jbc/TmYi5JSjFfI8zO0Z8
9U1Ct+f7IWIpHjusdel0h4V67V+uhRlbMg8OWtT2s4GNUxNfysozdj/T3Y+pP+VzwFsuSPeu0zD9
dNPegjAu2is/xBYMKVLHTpX+aazs4scwrMjcvOz0+nVLrHsErPPkZA7aUXlwEpPevXgpw8jtJ5zE
Lyxmvlxs1WysOnjMCKS55MVgusz4Cwf3vc79mhsbWUDMmK/4Kc52Dx5nv0PCtsvX/iMtoOjfWcYt
8mQKBIRN+AWd7rs18VSshDq+SfAdFO/5NcchdiMDlNCG1j/NzY27UU1MFkrQOTSq0xW4GVtdUbNC
t2EeJ3PLKhBVSusZ+dDnxqU03dlIbag6T5VSQ9uSJkGe66IwwbW2MIrQ0UqSmp0wDNv06LaIdoXo
BzGSTs48QohZYNOKlli2fK+DIExk6pzQjZMVRRUSlIjzInm7T6OIcTti4qqoLXLtV1nrhNm9aX0d
SdCCIGkAwRc4MWRTMdAXN/dIh0zFT3uI0hcyjOkLRNzv/4wOFJFA+JPckB7hnl3qa4J056Nl3gvV
mkRdABHmmwK/ONpN8M5sKViIh0fwQjVBKBfgEulFJ6jrVZMWMQ74gi3M62HZzGonwCklzwJ8wSgV
S59khF2VN1Q/a/wZQMPMTZj20qyi0+NqEwU4QAvWjypsuu7F4H1oh6iQ7c35p/BcYXZTi46AQyKc
KAlr4vSZG7cLugy09itcdaLn1oaVXlje7cJJKOLsL8er6QHOnEVOE5cLFt9Zm6fmBTZlJ9oiu3FR
5J/r7T9QeMp2gkQkmY1wRQnz2WgeuwaXMJUqK9H41X+6jObgKjwCKlG6x5INUIjWCXhdRX0J1HCJ
FiVyyaMVZZyUOy/vdBDjZjLbHWDVmCqI6mUR+pPfmHMYbFjnXc//5M4e9OXJLG7qQyiQ6h898L8d
m1EEiHAUW6fZH2SotDbAYpnDdfa+kyTeDJSmbAoa8XUl32nppE2+DOzkuQD8aGxFT7194aOMJgVG
m2NH+h6y+DkUYGNF4pHlzHEK3FoERnSRA8uRzSQ7U7sGEa4juigJGCKCkNB3d5Q0s9d0ZkCe0y2l
TkjyjEnco3ujojseB1qx+3McvGpEoNjX5B8GZX4SbD3ctUBD3iVNLEUBuBPY2ChYaJB8ywYQCE+Z
CCf517mz+pJi7IiRZZF2iMCS3jeb4Axycm87XLAQWMct5MvFGrvThgJGUb8yhCa730jPo/LYXNLe
kw93d4hv+4usiWygdHnxm5bHBf1Da7kD2m719R2YNx/WK29jz96PVgeO0laZItoKNVMNHuSLvOTr
qSqvTBycX5K/+OOJGsihp1Jl1/mdsW+7AfiLiQPdsPaSWn0c9SI/7NxqKYpWaUj5q/z/ku0ywtEu
4dNvOELHBUWUDvgP9UuhaP8kgFdBGi2K11zoPHsbLuhbWbQGNY7H6p/yspAUrEos3s89Kf8dy+0K
2hHfKbaO+4JRhMniPz5gtbDWbApybzrTucflsue4nlyBRCQGel7lpPMdmLEjUJlNqQpeMlSI9IAp
cp8iSIU4jES8KIzswVmYi/AmcB+ZFjCTKUhL8NcSt2pJtXT7h6dYeT8HUtxkz1nfTYynJOAhmFWX
z9hQsZeJ2JBLZM9N0HHlEBQYyGACVoZpDzi3U4UMT27/PFe3mrPn7VQWEhKKGA0N/x8vcxGFEymm
9NbKMhg9/RdqE7cRwtNpjMT/Yedfmqx9YHmW3H1GP1MvHv5zdEbSYIfyn4uz3iIaMkyshauo1EFa
ZWrXMOatEubImcDKDBNrD9R4fpEOgxKK/eXp/6vuePqvXW66iUHqHQgr1T9vlZpMSedqKMCJ2c67
mSJ1QrpbK9UvoIii2AHcKr3r3tSUtxhh8Aw69E+1tXUcnCEG5Oho34VY36FrYfH8yEs8wTRW1euD
pS847QNXUry2dlT00K5WqvUHWKDchT/bKC6/tSSVapRHXIxHSlNyZVo9T1VnmKwyHbr6lLJAV0rc
L5ha4EWMCnLENWNj4/GkU3eWAiJ2GLbWcC340Qhyiq6EVuIEXmS7EJiyrrtBf3aQnPpY9MYZX8Ut
b1ovdIwGqtCQxNuVH2urKS8Bn80wZl5aWY0nPkRM9JaSLDlkQL5M21gScOpnYNnqzPDWyN2EZ3Cx
LSRTaQKK4e/6cnMQQ6o0DocpcT3k4rhFYqK3NhgSngA4UIMywMquno4dWBlD+y14hq8WN13yvY0N
NQHJCsIgMwLqbDaXEIX1UOsnGzzFlJuce2tk6EyVNkz93cGs3Ec+ilGcT0R/pzFWE2RvCyoezBcR
ptEF5BYfDGS3tVXguV1J8NJ3nRd3gR7j6hJVZhvDY+B16/Jb8XYvSuHk9+f/l5V6s/2Xgb+qs2/y
YJHKk/EAihcUGbQEhC/zliR/SqoKwyCd6bgdoyjqE/9yTc7xKlqJ1+qht10V/wxM+/fqqlyWR1sx
PTUCjkDbHMr1XuBk33hq8UGPgFzJQZC4F+jXmKnMYTQ4bdLbP9k+MPGb01eJcNYJzi9jKqJal6fj
oC/6z8lU3BHxEPvJfr9HCPXgF0NDG3xmkAiwEyozvw8OZcNwD1gcFJ1aV37gFcN7JKwHKYDAkuz3
vzhFSy30szfbLJzop355qXsdx8BGGraWdDxNDBnHmJzbNJbOaft28JuH+Lf86IJT/k3FHJjWDVXG
eh3XCfN5m0Tvrx8KKehLVmJiVF5C3Pw/Ppo8eDpht6N7wcXy6DQML+c/pK0U2jr64WmwzrJH7OSR
efK0bwdJ4c6+kXouRGEgYqRAZes80/UpghdEs+asUmfrfmdoE9HwE1WIqappEBROgh5g3u6XIokE
rUAWDeuGuucxXLIEG7puaNrP72TXv23WNv8lowJsqonduqY3JdfUQUz5Ev0ZKAvjoogjyuHRFLJr
7vzBfA9kyPWRT2Ysl21Ly1Obfo9WZnnOgD4xbXGuEylZPeMoGYhte/pFU/VQjl/iqzPWZj8Spuh9
JnNQgoshM5RgZgdM5pR5Y6lksbZbu0jyKqv5XGbvPxgqr47LVQv/Nav7xbWM+ku+EzbmeMB+xlFh
UhXtReop/9lqEOISG/bu+Wj46r+z/er4TJg6QDr3dEziPwY+EqQQU1SkkHYHT5T6GCR1p97hcCu0
YfNIJwuWdaiLSHB0kgGcqqo5rzhPG2LuM9EuMI1WqWU6T6ovFAEsGBVuva7afeaMbxqKOenoZIGX
lrpdiLgbqhL3wDj9uZrx+/AmIN08VMr7wYbvu4rp2E3yMhn9HBAv+egX+FzmATAe1xZl2NtC32H4
aBtMUfIp5wdm16CSKku3IcDFG/t34XCCclzWUgZJQZDX0lgHdwK5aHZBkta8cFozYf52Td/J0uSj
f0yyzbgcwb5ZVjtntnzLWLtvN2P26i5fXWNbHAGqxe2wb2Y3L6UGDRW1ZxgGKjvUWNzj9ySWaY7k
vVPmEwCMTiGBFPcXKeaT149UGA7s9SQjAmNiUJlw4+IfJJMsE1i0vNS9AyPNIijVl9SQTTKXJfH9
K+/hY4GhJc81XuMp+Cs/ZTKQWfZSfvI0lIx3gkXAfPu9izSlKfn4/8/ttM/Lw92miLdLYgF7CY5+
JuZmA+/J6pEq2bq8QCV8UBffEwx653MHkK1TPyFdHwKJoi98NCIPLqo3sKbyu232W6+QzCvcO4FM
j02ogGUW17hwyxP957AMFgDbVpzRBnlyrq3TWAvDAzP6cvKxWjPIujxmKqX79T9L416NuRjuhtLK
k0AnPs0d0Xidu1GNoVbBT9GEmfJsfzCWRKx9JJ6Hj+cujNBCnDzzD8hSq1Zud6FYHAu/XN0CH3zg
urOJ7YxCeIXHacftzeIfWmhij1i8fRZdwDflzvyiBLQlBrBpRaC1euBE2IuT1y/8nyc6aQiU1vkM
IMQBWB4w9tiPORmdDJUQ1o5HGFyJv3UtMndQoTG9wZiZX8f3d3kFRHmWTL/byQLsPndLLQVI31SL
5fpjGrgiced/UhL+1VVLwPRiwjauGxkyz/GNfw1lFrlW7ntZhw9xPzlZ0lkvHl3LIqnVpaQkWsy4
LMaLK1o5/LMFgm7LfZkuDQU1iEb2VthcxkXvTbeXJGhHn7c+BEjMh6vpAmLGGm3bwdn3XXcU2iWw
0A2EJ14njd0rm4yFjGdhI7BYDNH3cH41wF1HQ/Mu2VFcCoHF7WKatJHV4crhK0Gyem78Bwt+FgNm
gFDVuaNNls8N2A7zEMuZSgjdiO+PYpxMT/Ny5aKH3TdAWtF4nGO11KhvdMkrsGop8iPnnBUJSM+Y
YEmmS4Zx9NcG9Fb20GPb4KpLnvySjZqzdQFFNXvIzFtSeIbSOWoa+j8dpYRBdkgK2fNEgmjJui3R
CbOPU893SSQx5IgfXPVVONDcRNRK6DyZrZr6pxBvYoPbRceCsEPHVOkr9fRi6RpmKf4LTaQxHMpW
y9sYfIxg6jece3OfB6dOTA9q7BXpxbDVPgvVYgfS4MBIj+NKWxlApTe6uJ3vUmoQ1ci5rXi/6t0e
8peHFNCeMnHFkIgpKq4JelfgljnLk8V6e2objHEdHlddkZSbvGK41p3Z4v/pAKGU4T3o0iwFJgl1
BJHccyblsh+y/GuoOe5iWFNnPoLuMeiXUVBGmSm0I6TovkfnFoz/r2lmPYEvu2mYb+eDN/W5SK0+
Y9/JNjFFgptTmYgheRms9/YkbOvV5Z1u7U+pNRzZ8pubjcxHBWjyzAWOX8DW97CeSzSOdOzGM3Iw
OK8HDOwWvafLBwQUx15qd5563vQDaJt3yOEAsQkicz9mdPCicm28A/YaiPWdF5+PCN/RKk9VCvYK
aegyHDUmo1fSwAf72SuaZd8wXLIoI2NBXYlXoS8nSFH/hcyqfM3U6+ngjApYT7NBPoajsHIEDAXT
xeY5fkutTbljIXZOvZbc0obw7iU671VkNTZKeKlu0osGvQgV5eaY9UnnP/LXwlU8nwjIynCvFMSG
7J3qQSJmmnvDQZk4EteT6DDKjqMFmHX4OiLr+TTBLBFuzufqjNGWPil3xE2NxsHGbAHbuD2PNEIh
UX4912ropTNa9+/DokZpJvNBTRJAOxECaw7gqVRUsAhZp2aBtCXkItc7W6NIkViZ0S/1qho5nMXs
P6joXxLXYZCQVscj/+fIZUYBKcGMp8rZ5P5SDpicBLsMaHnNGZJnFgJiuAsXbJsj4XjwWMm3EOzp
gm4x4aHILc7mj8AN4msI7Wj+VYdVfeN8UvPeKwBedpYOM4p495tAVAk7wGxcFhYAJysGSnGGPi/f
qg0F0HjC/yEhLf8K1eNwxJTBuaujZmRyepYEfS8EkZipv4+7rztDOms6V3YXYb0fIyk86cVPX4oo
w8L0LHJY8xG7TYLKxAzhfN0mKsohp8hEqkJelyhxTCweBzgBdCnaEH1ev052dbVsazV41hKqTRWz
8ABKCpH/QjXZSB6T7ZdKiz0es/zzzPeh0ngt1db5icjbyMlcTC97qbIJxCFa1rICCbli+CLmsdq8
rz15pPZynYfNNf+jrgV77khjNJuT8x8ELjbW/Eh0xtnbj9xJ7HCnKokDjPRozH3MJ+ZflTEDkko0
pisyRprOrQb7y3CuICKvh+XqwpsyKD90onQekhZneOXttbadCLp5uaOcLe4bCB2tZJ0yAq44Am8L
FPwF0aRTqN1QHHHgVZgIrSWAJZygwlvZsSEY3EBcI3GKtd0KlMbTn7cnRVt4c6kNNZqKAmQDObxS
IhflWI5n9+MmjeJ1uzp1ysWusus4K+VcKBoUue7ReEoCzcFzQcUGTZKP3avJ28kn8guvcCS8WIVG
OA9mvM3Btj7nQ5ErYgPFj1TcpcsBjmp4XDR7A2fIQrSjrHySbzSRSipH0JQLwGobiG3R47suq9hp
pu7G4pc2lkPqWm4/Pf5iizAFOUreRIgdS4NfqMiOkkNva+p+TeLGtghIxjRREZlfd3L5h0eDtPqB
pt36hjOsZx48tQRNnB0vOlFVn0FRqIXzNxAWNMd3noW46iFtJKRKi/YT297Td4ebwYbNkanAOjb+
JfZM5+tO8r9U/c7SvjNMVwL4tgb1e4faExYUNRrzPc95oVx6OzO9eT6XtsCByKE34T1kYrpYAxd9
rUR3TOUvph5AC0O12dKTwLGFQxImcsWbdTN3f+GdhsxcvamvDdifvB0UgV7MbezcIMBFhAJBcMxU
izNQkhuN9B0wxM7/7zvgiRhN9XJFqwPCoECCyGjRIxPWGpTIQ8TEvyEYAWOiIOLT6ddfKvOZCSPJ
TLHEcT8u6d86wI/neZqyKMjVJBEEU3axP1oEiP3iyXlZDecCTdCibUGN150Dwh6srQfXW9x5NLYY
S9wzUPkJo3gwOs9JuwJNbGXuZ5ILFaxIrs1wBawvHNQRb+oaeZLCJqCvSD1uwPtcf5csEGJQWOXm
TrI3/Uq4M1UEyQQZcpidq6geUF1kHEb/9aj9pOSl7aiOiI3IEhcQszMom0xQ1yVs5axSnatrIP23
k0p60Yzpvk2zFzQe8HBy82tJJ+1vVi6jQdUwLAjnrXu9GcSWKeMJMRxw30Ozgpudz1sn3tQFDLHZ
XKA8Pd5xflhDEwQR2+IwW9kyT5+tyzNTSe6wBnx1kDOATXDV+qjp6iNhUgdbBe9nHXvjuRGfS6pP
oLKkAAGRi0DtA4SrlVFOHQiiZNuOIdjdyjzy0gt8DyO5j3wSbXv8s2vauQR702aVLFt8Y+Y2FxIP
Z39sC41HkUrCVbSaerg0qiN0CKePxcnwGkuKfTFV82Eeh279GVBS5Jbf0oggZ+VBeVqXzLgrPqaZ
q91507aJrp8SeQE+D4kblT7Fk9l/UHX67gCeU7cHrumeBpIF9xcljK7ADL5GB9V1ykZ15topD+Qv
a1dEQtlDLAxxoOVgUMEFGHE/N78CLcKtfXpqnRFgbyi0eexu8kfByiI1X24/4Vd1Cmd9QDiNrbk0
AxDFpjIWaYt11w0FXXyNAgjk9vPFY1YqJa/1p3nl1pSLWrGYinPxOMbdddRcDGi1IRg505LkJEc7
PD+V1/+MOGvIvVsqBZwndaGJotwtTZASB9rFx6gcmP0SZtmbytx9zZU3AxdTpU2Y9dLoueedsjls
CW3mKyAdwUCXmgFdDTlkm7+/cFgOSCEMq3XbzHWMhzuTx90OJlOBU5+NPiix2woKeGmatMp6aq6H
5C3CGqIvGjjWIuVqhYqpAIZ5g1huhK2nn5LD8+aaawCS37Z/K0x7g3YFQOJxF7YbpvJxsv8xZbqs
MQr3aAVACuIzxg+YPOxo086+lJtKFak3puQXUt/gLQQ6ZQhwaXvrFZYJfKbPy/UILqKjdpDcZX5Q
MqLZ3hYQ9VWAdFYsGaxmpTver4PFHk4+j2HodWhIvb5iw+jNa5wB27eFQmoEq7LhnTnhF7pSXSET
OzBFdS6vz6FS9qFAsZk0M8wrm/bOchyBJ5AUyl5e8szJTQ067kmfABiYvyq4SPxGEC3IPtRqE0ek
yKqAnzjm7WdjHb0ePyb9enJwe43aBGBI7CxERvuF3RbQj6o+fVo5mN4/eThF6Ps/7n2FkMSMbOtS
sOeXh8kS7Asbdpk/9CgQAWdLviKBCucz3oD+BE0J+5vr2eFGpPTjjvQb3MsULV7PRlgDUXPn6LwD
S5PtpkzZepWQV9wZO/8xUhxDQDQoz4cK4Cnii6HKWJwD3k4511tWdFsXZhmKOnrr+evTyy+BIjyN
pxHyHhIlyk9FnDKvwW21X+yjH8D70VHjxk9ptu3C777s/Fe64B/UcX4TbRcq9jl7oZYLFWM2kMuQ
7MZdfLqr5sP4vYpgUWP4uFaC2tA+qZjawT4jD9CA79xq0IqSUYnNQvbkjKqkXBEdWk7Lh4XNS/Y9
0YQiuXU27944v5OROYqn+qoULrNkZ8COfdaYhljukXjD7NH5b6Mo/SqOTjlu5GBEiO+jd5PRUwrE
tLiwWrensdFjdrtAKr4HzmEm53p/4cE+Tet+zO0fN+TFxaKyB6V2iODE8u/SULCVpHMmNaxqjGcT
c1nqitc58jeUW5AF3y4EpuPkwA/TZrKkg7hrm22nSNLk6MPSjM1+5PLZiwDmdBWbsuJfnizK8rf6
UhOh86oXdOrOZgU56xNTtj80ZgOXmuS4VYMnryH+iF+doOTvrsic03Cnckq55pgq6l0XVmBsgSSi
4pYY7Ny2wcqpiKQtMMqBRTXFNEyIn/aUsl53k8BzQ00T6hF0cNrEZ0/F68LGw35x3yLmrOGmHPXi
tcVHoore9YmJ4sr10Ahyx803haO07+vzZVdxxMWcpPQgOzfnwZ30xgtQc+/Ay9eZZ1YQGiyeT+FD
UnetKt+1CqcfqZHuiNqA7vDDxl3aaS3v/S802N3zXIp5Y+uPeAT9DZIWnyuA8coK0aXH9QfU4zRg
FMfoKq4b3CYsV9OaEvcdrfXiJqYFdYatRCvBGLrzakGuU/hpEutufVcVs6q/kvWRATqpkQNHuG4p
/yDs90nwhp8UIgJcPl0IPpYjRqKynvfXKsfuQ78kY2B3Y3rptWsmbHzek7jP+YaRRL/lD5ZM7mFo
eCUWHoTf0KcZhhnGhQ1ftcTcJWdGRhcaLXMMO9IJRLKaU6ZHEfM+hDrnPxDUzrxFJL7L31nQwqfX
KXe1rJvwPkUWXeStHil0PsQQVHINZXkd9nCz0anhT0DiYI7N8EmS3Z/xn654cA7IJt7AStpRK8xh
g8vcjYd4DpXnsgz2eoRH7psdkcw0+VP7SKbNDEi5CxfKhC28GQwvGJEC6gDSbJyTA9BZkFVxEtDB
Qhf/yA4/D3mxFIqBjSnQ65c4odgY3YP0RqOatl0T/rfneoXBqW9YE3c5A4Nae378zaGCtetDUeyY
m1efyK7G2euVQ455Tsb+aqy1W9ySvTtUOn2GoyF7jtB00M33alya+x74Z3EtIy8WwGy0K2XBKFEi
3G2pqLa8GmucRhBuKfyPdydIz4LP2QUZFT8RfGGOSQUwwO8H23w2a4qGS0NOcGEViXOBqTjXPBQG
YJt1nEQNWJfu+5DQtLwxYX/LcxsiCHWZiQDyN4JmnWDcOgFgBX2MOk1UHztLDw4GonJBgEcFCcms
4CrqBZlXPxYmg+dF4z91uG8hFm3N2tzzrTunTy8q0NxQ8fHJfU0ODe1rO9ZmaB4XutxaK/dg9oxi
6gxFu4GTjjLiKJ2Wj85xzSWTat5zSPBPbm+UnmD2vzizuMRRYmQEKTJ9GQcwIz/2c1r8gnCwUjbW
6bNWhuTtRTjPp5UQAy+9AaqAZvEfa8eukF2y5S0+n1dJIiUcYwXmRDjObNpgwb/6t8o6FP+pErSY
lSQNXSXCKIAkI8zhqdt0OQE2U8URNh37Ao+kGsfyw/srzpGYtg2UaBGuvOxXfJpLOGuKxSmhvC2i
Z+8tZwWSB0VLgtDtFhwoU1b2KdsZwrtnAGjEArzcX9nwTVDkllKMkmFYTTq8kmvjQWhwNmQPcDWv
wA7XXi+2nRHp4/YJLJSULNZHph85T/0E1FNupEqOZTy1Pi4uqwRxQzZkAN8XZNRRF3jXX2qaJmAA
tHf8ZRNGnnhT6BpeV+zdXKvCLp0nXbMMe3pqdXjj71Nv3jJIhACKjLy6Ebd4I0JH7ap8t/cxeJQN
hVvNKrahueO80b4HIlk/02qXsvPq0Gc9HilfAnEFfLppXpHnlqp1FDhcfCSSUzXaBKLP1xi+B6GU
rgUD9iuMUFkBOr/UQw0r4TtI3qxipCy6GRfOWD1pe69NeJa1383sTNrL2A4jNULqfJtV4Gap4V2D
ao4dzUHQiSPfBfjp3neDm9WEZ3EOk20fWOuPsNlcXrev2uR4agEE5DSDFIjC8Kr8JKmCzVSNLWmM
LutoHi9NY2OZLqm3ZjNTt/s2D4xV7VrxVHmpZ7cZ1n+nuxxLIT/9W+duwD5u7e/I7hQlF1da3qJc
aFz/ymK37uJiEvPzUZ+wuMdaEJ+15kGSZ2g0wC8cXo95FpHcboG68MwtLZT4hX//FrpwFUcdct0p
VdEnBLcimpy38EK3LxUR0wHFfb4ZTuWKe4eUbUul7zy5RV+Tl3DgMQelvtHjVwqpCECUwwH36Tw4
T09gXPINDaLDg0EVhKWdyvATlVOSH8WsRZWwSs6Q0tkCsu98Vccg5KPcAo0eTO6xLnV+EbXKL52f
3Pfxucc/BwOYUkopGB0E62sPwgVQ4Nu6hOuSlhbnnXdzMXvzTDq+z1yjd7fZQoiMm5JD02yhLG+y
fEKQEzzln2aHPmbABTsgmgDw6aPPn+O0EaQdeCGSz7b6HeJBr02K/WLbYNQlV1lmZ56jbRuEjtJw
Tnhs9oT1Aa+J/5ZRM02TWKuSNMq5WRid9kpdXqZ2E8yZkJCbZo2qUacI8sV/5lslb2VsbqXrMuk3
PwcTTtJaXvKbHp7NTx7YRZ1C+gnC5n9eFwW5bR25Q+wPvbetBX1iRczZMP2EbwEdbj+1SjZ1iLYc
E+SjHXt5k6r1+D+9tncvBqHIdXonnEOIgRx6U5dlM+egMOWjqMEBHYyoSo6P1vGd5+If/5r0BSTm
C3Ovziy2S+9yA3mfGwUGd6RyeHSvuuDkByf8OjGMR8OHzLjvw991wnCy7MmbWNeT6FZOuy6nGxFk
M73RKEivUpn69DS+X9N+6NEKgl0MN4Cx2V/FNnJRxDNtL9jTHiUzEjzVP8qAvcyjB5epSp7mDmRt
dj1Rlgq+1LAyQZr9c8/u+CgXCTmUVo7NMKn0iTKsc9r7IIO6UZz3eTUxDNNGl49JMl19OUW4/DoV
bE1EjNkZwpn5QB2nYbUwHfhdKLrwLz9iOkgH4nbr6oJYjw5xFThSNc7l5C6nn9mb9+TR/5Fmhwm9
CmEytpY11ccWiUYJvBQ+RdzshuJk6kcsnDVhcBc9du4j/9qhksxrIYu5E1uZLYo/0W4p/rBMITtK
glyCeTvggMyqD7X6IEItK4QOYcuHkyeaeE5PoeScZBax/i2d26se6mGyapnlk6xmvnpIAKkC0dzW
sNme/dZkvg5ch8vkv8uxpwyldFXpZQi3UzZBFL+ax8e5Hdyj5/AZ56xKvnH/w34FL2+4Qk8BYmN1
b2WSbkFxn9KQCftgENPidYu2TLJX2eXWZ4OicFVcTcxEoEzGAjr6Ye/EMidjznvlRBG+OkbHgPa5
NQqgFHzRAsdIozme69sxuqDemgf2Uf8iIj33Qe+ji0AaeHam9asslfcp6GLi79hIH2msVnhrfH/i
56yM8WBJMP8Hc0kL0myPXoZpJZFRtMZ5y3+dQPyv1/BItG4ReNmTCMksZQKyFl47p2nATVK6FLvs
WAocluHYZGq+xGNKHCnMHjihY/8XOfsHk+0u4rfPn6C2Eg1Dx9FUB26QMMH2S6PIakotF9fN+E/s
o7nkiXfX+pMMoJg6giNN6n+bCunlwSW7rZCqE5KcakiWhETLomyl5uUQetfkQLYVzKhxBhQzL9h3
0d3INisAoDUq9FxzKr36UpSUSiua6qvMzDU+Z28bIKKk07jHFOvMhR1F8BZyQZ8Vabwm79rQBpH6
9D5KkkIwdxn5RX3gsU5/+s6KCVC7muN49+BG66+GFEbZbtSyhmZ/ta1qnQ28uvuL4bpkb7U1kVlE
hEi5dZyuxP3TvNSav+t8AQ/9Fm708RFT64w9OI593E10zNIi3XSJr+QqmMeruhyU8g7nBSLMzc0M
cxk7rMB3y+QSe06g28O7Mu5DZQG3lKAKvpTPkQMz4mFe7tNt8TtpPkmi7X+RPMuGpyhPK9WhtquM
QlowuRRutrXHB39GD9iMSAYwaqg39RHOtNAjDh+NdMkJDtcugDTtUQadGoYaAkwDsFddBPKESERz
WVL8BWJwVKZ3rci556V0YFtl1JcHXKpafgMjIu8UD6peyPqRE+AS5xoNJqNwC2GIRphBWR/X1f4e
OiQ85dwxglyBuMXw7T5yC3SRhuXrkcvBLLE5fEygHnWXCM7kd/yV18cfRLzyWwsC4iWa79CO+lKO
idXbazjTdGnjAopFj6aebHMUmcTCjyfUWIF8tOXWLLNoqEXfQ7Xq5a9agZHQYvSEckHLYupZEGTB
/H/DkFHIwfJIHrOJIBPMKu/jWMD3cqDz/9HAMngr25hYsAKTQHmlA8w/r05qQZYgOUtUt0GZ//oy
jvT3SYUznulcAww/fsLUiugcKua7sadff6GeLrAw98eSFrAa8X8P24T217MwaEEKu6zCOMxDYlOT
nSjpalKTZi6FeW/RWs4nXdtxxbpvZSFACwvXT7xBPHJbd6POO5FEFe9MCt4ifZ5jJ3TsK7kFSPp5
yQN2sMg6xJXzo2MStom9Q5CNhnN4uIpHLZmI5Yx8HCP+h4XAHqWb5lqpX9/nSxGKonFR3+Kqa3mI
kYxN6lRlKZy8Yd+i1LkPAn09fKUqWEkRvdGV/29UZ44ECSXbADTEFP30Dm2scGgHzc7l7q4I0Y/j
JNtFn+HAWxU7NQHDa7ta/Ti5fQcq8r+WIwQdcbkLaZGAPQ2UCxca80d1tgaxL4kVAj/9Bl+2LYW3
3EXSLmIMF4mt7T7UrnyYR87TwfHUD5pEdoVYmu7GdB+fAzNGl2tPLfNt6gp174vPYn1iQ2RdKOjS
jtX4mET4IvCMHv1iI12FeTApBSecB502lQCAd7o3as7ybAwU8WyRQlm0SMHcJqveCs5c+XEwf+cM
1kkZbtwCI6YF+Nefos7SxFSxTBQsH99s9UlKPkBujIvLmTi8JC4d2/+9f9d/xnkuq9uNWKSmPLRB
7QS9k2SEB8423+eyZdwzOcDOICQ8JIV+ZqY/jBgEAQssS9P/7aH81hg/QPtivtttb4Rkq3IipnOb
SHrs2IWUtbdpDQlywWo2ezzZyEqPNuvrC3s0bnjgHKIOIjiIeeCb1fDUvD+KrWOmCUcC0nPHjUB9
F/VTSpoAywiZwvVMTqjD5BbJ/dNQoMTJnlSsSjViO/6ueUbGQd33MnuNDe0KBB3YztBma8O40CYm
o6KfcbpsdLRhSbR9xnnGNeMPQpM4BFI+QdI161BkbEYcet/eENvhdai14eRyYymcS2wKXsu+OjLB
9LvRHcjirlpLwpk2queo+BCgALOR197oXWNwaGBq4SSS4LvyZpvE127272ycEOhQiDPsrZSsA5Kf
V8wAx2sfoA5mWNb6B0rRPE0igQImWJw+sQy/V9nz+2uTGIdhrbUauJOFOMD5GlqF8MuZ/ZbdNeEo
s8GYv1nRwHrAugJAEkFTFj6Tv8QVweGdrioYjIiFRjMGTOjR/cIsLOU+0eOMc7PMkdS+ltZc7B3U
3xWF4napM+ssEmthFqjDlXhqOYM9RGohjt51U4Bvqt/1LHgmguE8/7Cb06rclzqVQXT7235Vr/IF
fkHJvIc5LhN9K/6XyApqLLLg194MEZXwfol4EGToxHLdqK4eDU/FLP9wRCpoMrPQdHab0nAw8GDK
UnhS3kWsb5BP/TwE/VPGGmqEl68DZ5dvcdHPw8BFvTt+LKE1Azqc7TKHVHsUBC/+VunaxlByYPEG
LTMyEq0uht/PYCbWgNkjBHkVghKT6b3yzT77Y4JfItsQmTxByl8/806zvGXGXuUP/g2VMCr0xDBf
qtpaem5OkTGCp5GOc99sKimjYU/+ECN4v+5gz+Gg3ohnjl2iHP2tZRgQ+c00NgkjH19KKL5XoaEc
R40ra1v9aSBBvBtVUZjUerfqJ4IJV/h3LhpZ8J2wdBrxI8WDnRnxEpxTShZPI0Gr2pddxpRO1L92
GWFS6zlax7i2s365aaTXEvcYvo0SYCnjL2U8m+w+L5RpuBLZ8ftOISZB8OcqyL/y6Bm25GnHyTCv
Fyh8SfCeZysSUdwiJ82AqnQgr+1+mPHK5upz9FfxKEj2odLpxRaqOkwnIn8iSEbMnbQnKiqITa8Q
H3nOrp11cE95pq4xAVos57Z5FxJSny1BbHILE1zen2ltwYMyW9rawRLxSzBTfkynzY8Mprn9IOhJ
G1nvOd79/d30TVg/WwuJYPJhs+ltNjUYmGrxHy1RRqmL6D3r9coVbyl0R1aTB2JfAO/i9LyHjbpV
NRMGWDwpbA1cBry5ro2FKHDARiJU8OtDb+FhW5vHtKP77binK9L9YMvfCsjxarotOg8OStuR29XU
12Z6ljtcRBxzUenAbE0ZPYxdi+M+nN1aj7hbDojfR21QImcCDHvYUjHnQQfOUxSUpF+GzvD1FFDE
cGm8QHYTCjNBCs0MJt4XPusiWu/CKh5s1ahNqm8bJFlZjQdd+7XhXJKnNdKc60/CIqTmc9ufBjPF
balp51XtpHIF7PHmZzyRiOo8M7Kxs2Ljwkowo8Nnd2WBlp9YX3Znf/Kh5ov2NbZLArPkP1ZOlYJ4
XSDDLAc9z8nuX+/2DeXdAR2KiC0ao7dRH0kLO/sdIZtu1Ul4AiC8YI1bAdAyOztF6EfSmvcWYFxB
tLfWiXPB0TlvgeXzVJrR/8uorWiKnVYwUzoOLSFcUjF+AamRUH5N1614dORoNShxGmXUkvQCzTwY
a94y0e7Y/EiGVKl6MDwWZFOIWxGdwnWUgosx/CVU89ZZw3hhpM1Wh0rxraNKNsz0tqG+9qA3yRUT
mAD1qWzKa+UQGFwB5eRtBEyuaWJqS5HNqugHy8mTowwVH5a+Fsmtn1JSbgmD2a2GGlbnY9thmQ5s
LaGSfFAZuUOOlRnF8bPq37bJZWQ47UOIWZQMiEEmr/mGsjVTsPkx67WYu+h5uqJOMOiAOa7UEEgX
H0EPNEF1FIT4eQGFG9bRsDd6UmcbuBCBjhWjjiwTkn2T/V3X/qN3+jfGLB8FMy/PRzqgaJCJjlmE
vJCw2zA5UMmZojK8plI0/LAUr0ZBceiYSfHJFZXlMnKUL7Fz6yW92sUE+8pAmN2kogEZAkpjlany
0QnseqH8HM55QyQxq4tM4ZL6nToJnPLE2j/fKTIHgqKUviGdkGRC4V1GO1MNEjFnkNyPeBNd3kkk
HOWvMi970TG08HTzn6nW7YBEzSfqPPYs97aSHQKLP3GhtedjIUod9dQyIP9iwzO+dFCgKqCrqkzl
2UoI+SA6YXAo+WM2oVsZuO+dlnf6VO6JVgtY1d0e2kxBcdlR6lZLwntumJ3511qLk7YJXHMuvY24
UCfUMwa5t+bn1T0QVk+DW5xgXBvbNgoOjYQl44Kn/Bxwjvkzcafrth+vCJjviOPmMkNfWHAvn/hb
hI2hLSnpDcjEJIF2QMBhotKg5vApfSWq34LwPOijk+2Z3hjOMJrYupizsheATJm5bv7qgySKBuA2
vvMZ40dCTVq+rlDC13rVWzThkkIkLG9sZMQxtKpNeOtXsrWF9ZEWyafOiTNeEvcJYtAgM2s+cX8N
iOUjpAlZ43lOH3F2B800fzyY2T2ONuvz/sf7Iz0e/f+pdaIrRqAe8C27i9mKFSkkzlX3gC50CgMw
Ek3UenPbcvw64k2XpTZ5uiAo6X5Mi7MayZu1Tkb3m43ccOpZea+7xpiOUxyDiBGDtf+AVqn+R4Ll
cWLqeCohE6YqEZlx/Dbrh2yjrj7uwIhKJSj2Z5P8zuWGx14hwd+UHJC1wo1VrAALaCDCYWQ0eXx2
SFT356cPwEqth1qIOlkFjDur0+MYNYr36j82P4411pFk3RyDRTRXg9ADKsOezKh/qzW5oUsTBPno
3dTuWcuinSZjoDV02Jcqz1Lvu/DbEShLUNS9qJdb1Joe9AMTDZ2/RRSEQYdqNa41qGt41hbjNaTU
to+xMl5wWKZZW76eFDZD/2pZr7TRB86M880VPCWJTC2nBfAA4uiSYHuSDRARMUSia/4A16SL2Nek
C725FJ8LcMDHX4Lv7SltT37Q3yfv/7V/GCOXi8NVnBkzz/z4cABjwEO+T731Hl7NHKjjnbJqq7J4
bdAkK0X8rlhSkMC3B73M4lBmnHdjSDDVJeVKtGk+Pgg7x5fgnq2QVuWEUt/QFfn74/i9LnzMcUPD
juvUW/pIwuOBNVv9Oa7T0+KM/y02y7zvEgVoY5nJk24EAEklt+Gqth3NwRanNyTxZsnvoeoeo3M1
ChcC1vB2o0kz0GbkdSVvUrO/JKdMtcYM9fv6IEZ7ygaONT+BIkd5pY3czB9CpdshxMK681mft1vh
0ncSv8dekPdtvglQ0qJ0s+FYXwkrhXzoGBIheJdFDr8Q8Yd0lKbGU13eOoZQuYbrVeK5XyE825md
pmqRYo/ivBaFuHOTBR/SnPv0nrU8ZxlFX82Y+A3vjWcB4FoDAhEgXtg/poQR/4EXlvFWp7jtebNt
dHYOfzku1RtQd/edwkSOBkm7HX67fv45zAkJBbwcSvGNo1s5o1/J2rC7bq1C1d+404W9hu9SIbco
RhipXG7wD6zC1RK1+c84XLwEeXuREqCCvnFGs0Ocy46zBn0iYzBtPImvN+4E6CbClpV/WPaSJ3nP
FGSgZcB6UvOTRxT1ECmhrurAiTzmeMWM3CwAQvWH4JuivK4IZeDZhqVe7DT+bhMFgUChphQJJfbe
7xihjsMIbrYKXE5dDkBZX5mZ+P8Y1ztIp/COO2RJ4JUNRh/sAkhCe08ndatZ2JJIWmvRwnKJ234M
esKzmO1JUpEKjGni85WyO679W7dW3cQy/ym1PlpQ6opA+pI371R/ZTjrB4oL2NJQMBZVzYK71fYT
A/K5mrnjzbVGv4E/LxF1ac2JwMea5qq5uLujOsz7bVE5xxWHf+wLm5E60wa84/XuWe5vDDIngQhX
9anHj5kaYSvQ0qkkdGfjALMVBR752GmuoX3btaco7J/urdpRAXL2sVAX3fQYbS8KWupzGjsuBF0+
e8ZJ5cXEYm5d5WQvVYRL8vTMci/cXXfeZOdHEjjwYn1jV+bv7mDv5KZkFmHf3moCJsbeiccwVhDL
qshR5JHPeMGoF5GWN9EBQwDO8+SHWlWmzO33LUUij1NUn5GEdC7tBYBzAhs9WaJTl6EZn5tjuQAN
AGqqGkU5nDdSz9xBDyIq6kY3Vs5zRfgKsqVkEE6sUhtLRz/o4rvYl+BKqOYFqS03x8NYtHNTek3X
y+XZwBccKU6EVXmJ9nTapjvBygwF47HMvVxuYM5SzkUQObgj1dYpwx8juMPzbxqxH+JyIG/ZpKpn
K/lYJ/ht2/vSdheIhN3pNdlDOYdoPVV9dVLPNtel2wE988+7WTo7RXJIb3MkqoiROZYt4fTOrouI
FIcU0GMea94oFKUDrrH3yLTt+Grmnm39tYjB/xG1Wtv/POKLvc03pSnTE+feo3dWVyjORt6XsgXb
VDgYR0+00PgFbDSe93fDtrBfjJIO/5Ee0xIMOqvIy3LRX8tsH9O4MzSwwOQdQaPJy/8hlswDwNn3
ZrltQhbttQ37hK93pJyEpPsMt0ScFArqITGfFFCsRldSKS+CKIE7DiokPSc72fMzUjjgs5uYhfKM
ExCSz7SVtupljK5/6No6OPvfSgxGM5RQ7y5+yyqq1IqxAvHlUDMg6dgCcKi7VRGR+1uWGDgJ4v7R
VNdd81/JryR1QnQ5D/a5BCteI0WPRCpuqw8zJaZ4o1r2u8EjUTyQC5G6KryA3OCeNARbqcCFQAI4
PfPeQYe675o7LlkeIaNxTvKdq0EFNNXQLRYHTPfiG9u6iGjom8BEwmi7oukGI+sVlTHU5Z82KLM3
cBKayMyAD9XXQcygtmVPFYm6EiKLAlwiaTLZPao0cGrTskyhshqpyOo2VEIk6/kO7QIs71muki6j
Kz1H2Tvb9obTP0utmuMiu9UIzqFck46YlIkh8WhdmGaj0Ru8EMaDfu0wnav97cn6LPRlug24bl95
cIR9iOqY9Sfr6dFnr5Zv4x/SQjdtTHbgazO0tX/zM+Wg+7P8X3uFjTw02u3+ndWcnrwRn7MbNwPQ
IlJyGiXz954D+Ih/GBAageH586cCS8yCIf0VFjgoLCX39vMF5wmKoLieS4mEBfdqJb9MlKYG5PvJ
eMJuKmfqjFlkJjzvQt/ZAZFxXnJ16UUN/RalAnWhjpzX7j5U0o4/jA689YfH+6ZOuEEOUuZBqf85
3pFNhCilF6WUn2Y46EeKiEe8KYtMq46c9BzLWYtdwWckixaVw186IPh4NGURxU+QLy+x/U3MHipI
mb8q+u7fCfWJXbRxp3zesK3SrC8GwmOzscQPQ7Lfxrz8U7heH3yC19D12+rED6Az6kSriVFnQ6K1
YKrLYBXsnrMOZadBKavZWgAb0G/ejwJ97NKzaM6tiFvPeKzG/F4nL+1um7KYt58mgXcrx4rCGvzV
qk3tqlob//OYxfo/lrmM2GjOEp7GHarsd7wuE7MJ9/ms4wOSZ5+P4NkuB9T3hgj9uG0OejjFH3jM
DlZi+G2MVHzUV837vybxEkQkjUb1QKXro8KD5exTgQejuWcm2J0UIYhhw79g06DNOFr8uqOQD/j0
feMdj6rwejd1CtK5001hpe3SGEa/t28kjdH4npXM25dITk13FCPHKL7lvhD2UKbcaqbrR3jD7w+8
lthYUkPbIltLV/k9Ge0ALO+FKtESPvU9MiBrHxKdjiys3OSPMFxPxZeB80vT41aEC8HENTGC4tMV
WQH2qSG7pr3bvgnedexkfFKrIXKDl/q5C0UNKhr1AoX7ZnmrJl45OJIeHDZTNvQhT5nu+SmCfveX
iBuImK3DS6O1Z6FKsJhEjcgPd65Q95jds0wBP2Swd17FmcjU6hdKDP2ec0NDufZGlXUBckroNWis
hksAO21gWHC8iJ+V3C79wunl0l1WcdifuTRY+qOENdmZzZNhyQ1kJrmWf+6A8YmSJu5BKcBYqECT
3VfOJfEz/B1Jhtn38cTU1soYm4uv6eD9UNTcZP4/COQQgOkPS7b52SsPCH8n/+GX9jwCCZXXJNa9
OiLGzh+Y2R1P9VHCfBmcPQeKmGul1RtXiNuADDgTRdJ7x2WR7tuXrCGPj/MrKibBTFDumqwckjvq
8VquB5y280sp8tICspUrBlCB0OXTJg36CK/gMAH04iRpNiWzYU/bit1vdqCVxlAKl32ERAKdACcP
M8kIIL1sgMGlyBS9RJB32dBBtICNV6SXRaP3vJEWO6N2jvYDcfXhkiQlvbvG3OZnJ82uMM5MrRjv
cW1/Qd4FSW+w5ycHXe6vXxGaoB3ckXe/4dW57y/QbwPu8GvFY9YdAzSksO1udVXeDwhwVO9ooLNV
eSzi6DE1Qvbyb5drwHd08V79gSGJf7Pr9VpWRkIqVb5lW+tFzCjvBeqysS+CD+nvx6VQnywi7+ep
qPOXMqlf2/Bs0oSpy2TpXtCI3l7el1s29DAhqztKBCogfMSXKsPGPxrXaq6odkwVZMQb26p4u7a4
iJtL/xZ6I6SEfMWhw9+eriIOxP/PLCkLLxRScIVNgRY3sItANz6p4LUytrVDZJNhDqqGlVD7QNTE
Nd00bUxo268VlbL718PJSFqAKYg98hoD++ub8KCW6eUhALoxRMWPFzgnoXFahW3oi1bsLOgkm1qX
M1ZPv81tQIZjGw3o77JQEv2me6o83ZXbk2TvIxKeEZ6+tFfl0LyLOw6eM7TdoAPxKY3Damg3zrPL
zQj4GImii4rxf5tf6OApFm1iI/5y2JskxHfsKiKAm0abxZV8rN67GiWXkZ8JKDWTQxTQY/E49ANI
JvIpZaQO2vAFv8Swun1CHym7+koxYmmfRbtFc4XQgCORYPkN78mTd6JrpikB/v/JTqOZlr03bEAU
fwuorI3WI5wMJFndAUE376bgT1ad6+MsoN0W52sGufpY06Vfj6db63Bi8ALWvUB05rnFWxNEMVmP
z2dBKpdfocKpVOsbjDVb979CaWgxsdI1LnoI5Px50VVt0SkMV7wBGYxsProqE9mOipNA9l/de9ID
68C03twTaUYaOBYIyWlYKf8zq67tw79tFv0mcUOYCNOsoxCS78J2E1ForZmKKSFCKgPcYqPPGoGV
rYsX77yfO5jdw1JYgzV3yzYNtRZRtfJnN8yP543XyeaIs719RWXNmmuYKmoiwaUab5NhSr+dn1Et
i7JyQ9M1O/yx1aAjacHQqR07unjsmsV/VBQMOriskYSDtAtoJ1vaw6hwQOpbXk0nAHrkgVUhOqrq
aLalhC4vafCheI38hM2e8CoMswiQxEOi4yGWaT4GG+fF9kX0vqBIu0GlAvA18xdZOoDpqUng2qj3
V+QcU1d9ULnZGSOABItB3H9+8JluozEQs6gUtv70xMoBnlTOCd+nVSTrmQEwv4kGqFVlfNWQC3bB
7e6LMOIxkLUePsAuZA5D5zkPGbXV9yhqn02mtwrrBXrFYdBv1ym9gMc5757aczdJKo5yO/snvb49
qQebrx1Br7TKibmZmDPaaKb30SMSoMrTmhyxCcPBzEoquVzGh6xuG2vLg5MGa+ccqJtqBgKxSHCz
zYXXf7Eye1uqKau3yaIClruBPuCWqujMye93Je+8AIQEb5TqEp20CCPRKhg12rJeXKevBVmxjmAy
hv0+bf+qUbbKGmyW+q6U4kRHlN4jYfwNcUPtBEkJdWGzepSBYDIV+MlSPoR6FfaPk/rPyR96fW/5
tyi84iGLtvzt+qnOtHBzxpRr+kJ8YALzid67eofHtb1N4Z75QOvxB7aLDAs9+oyC54kJEHCO2Vv5
TxYB9YeycPzbrGSsOSfOImiit2BrwMu/WJOIizHSXXUQFknIjE/AhxFVuLKN3hvlNIz53y1yrhrg
XQN5OgOFEN2foTJqgUVrZ1bVgdYwL63wx43b6URn625IpmA6/6kOp8znZ6rUp77AjtdqnM8aiPXw
QLocUlzL1NoFT32xFxZgnpMSf5kiaY64AYP28JO32DWsd3ozF2vhA7TzPK6BTV4x15+5x2wwjJP0
f84Od/IWJBi5QihYHjuElq4PCOY5i9uFGHWTVTp4TekMw66U6Y51fNVM3PMwD8uZt5h7lkFz4UcR
HR5vu3t9r+4wmOa6IBZ9dhnr6duEBy4LqZxdtj6wt9ZFIlh+lVHdg9LVyINykj3awgno2MnJtx7x
s6ae9Q1xM0IQHh5VBdj7r+lJfPIdCiQ1ehposIc1/aL4a9fnc4m7K7YSd5XY38VeBu7Q6pMHTZC2
5zhuJ8W4A04AGmCErDXL76zARMlEb1226r/SgRbKDyX2YF9nkwkhQL0fYuDcSzk1/4Z876sAlUZl
Ot2pn47nTdoRtji67LpFi7PF0CK2zf9KjDbT9fDFk+Dm2xnwiXP5GYb0Mrn5iEOkBp86+fnFC8wa
na3Ygg1emjr8AsyxSp9xOW3LqNllRumevyw70+R4DY2M6zTxbF5ZnI572AB6S24kCe9xcEiwfUkv
WH4BV7H212Jm9YeEbDthz4ZBD9EMTpt/IN/dpbqxM6xOKVXHDvxKzIvrcgFCq+tCAMnyV6U83rTt
mhwTRXzLkJuw8kwifLt2kgBgBY3WmT3PbEp9J5Kos3Ht4lZxJD/gNvs9GeFBOxXztvfQLflP+tPf
MjDNiUJzl9MGjPiZRyKY7CKTRrOhZVwCXW/Y+ep6ctMGS9hUXKQTox7btu7t4hqWMM0TcEb4mvtE
jjUQFflPD7TNzDRM1nbsmKv0JNcaF3+fqaO7wbpdVSu7qwQlxXpAD1zguFbp7vr21MC5OkcFwSom
X4dss4zkvpxNw0lILVqCyeZV7DRnsElxyhjB3RtvY9KU9Y94IWIeEQf+75K80b47n4uKJG0FF0Qz
HNeBb1p77/y2ZGHauU4xcFTMzlHQotIpiOn+0GJhPWBPggUgRRSYOWiMPI03nhrAjDF1LwyKTvTI
FtKB7c87VIjQH8cZ+KXAkRrkKFL8LzK2+KV+TBVzihcl8jK/vPYEHEpzsINGirGvOkoHu3XzGA3S
PUFIWCHzuTj7uqxmLEdMYixnJEojqxbEsHvwFkji4GpnkQxAVHShz4CfGgbpxPENqzSBmXOYVPwW
pbi1IWloTf2o7ucvjQ0OcNhgqGa+h6tN+HL7hMvj/9xdny0wPZjtf5cIGRId4jB66ZwRG/50oCRb
Qc7QdXlLCLYBv2Ih0BXnBFruZSDWkc1BDDH7Zb8JclZfcLQKBd9CQycqdu+4Mb1eziTiUpDG0xLX
NC4/FOR1HKxuO7jojFZXkVIqB9XgIKTYpoumD/JHY1NQh7EUH13vTdX2cnoQu5qMeKs6X91K7KNZ
EO4LhlMvlWDb32ynxO2IL7AUk1LmR/JnfHl5C7nl0DXn5bz+p4VgbZMJwSYWZdp719bC1JWwTF3F
UqQHP8k4JO3LffC+lbxXtIIuUT/VPQ/V79wi0WJd7dA6fp3761TucK3h2rpzXSBP3dalMj41YYLI
SrWrXiBAJuKzNoFOeSWfVpMcNTBPRbw3uw1Iwr0tWyPut0pJVhL5P1A7LiRVmo9LLs1ltSxHnGqp
8rsl6ARiDWMnmGN34b5ybRNLXsmSIVK7VZu9JkYf9bAVqIOHrVHFb9MnC8yG6Sl/OPMSLmPxcq4t
wNkAONTmzHGWpVqpyP7K2KdKXuFgy23Uo8KAL0i66Iq77mOZ4RYfnuFJADcVbQ8Bazm/ojl2WaQO
xsq7MU4smB+w9ClzZ2QJYz5h553cpTd1CkHYd4eMMX4e6cBwJnq8JmkL/z4v820TNAmXvBJ75ufa
nNJFN2EkN8019NVrkJdjE2OLmJjcrC9nEYuu+jSbOBMwm5/KHju/3kzek/J6tOVN0a8bV/AG9lQb
NMjUEshZsETZt1JFREJfepbapkbFPMcfGgf6r4ln8wj2Xj/ySmVeT/BMFxceofFibKntBIryOm9n
HgvUa/JkiWlpv/O9+nihSBhjU96vj6G5CYmiYmeuHMzVyNw3Dib3N7ydFhfgl7mbP2F9rY2zcgMU
Vv5JT9oHKlzNDLR8yMBF/i7stzlILXvxXgPmM4i4CdDsyk9Pohmfn8M/gpPd/AoOlzwPOM4KqK0c
wh8xcsnPyiNxZ+veOZAvcwa6bAlVFMz65wcC8rknw1UzyiV/NYjuc8pLMm5p5k2R6TNAQmxGsMCj
T0PkWVbqWRgk0CQ6s64GktWVKpJvrl9iuD6mzBt8IADe5F06JN89CVT57CdxrCZ99D+L/e0xWG9+
9/J79Yd1nstPH/rXu58sF0FADhojx9y5gQLqN6FDOgsmuZ5bTmYy2J36lDSD3uzxOAZQ5pTpe1lK
8Jtb5aoxtRk+4JQgcp1nQ6OoWoKz0QRxG2SArSEQur4Kmo8D2E7F7h1xbTzvC5ND8L0YZVN7gk3Y
+hoqAXaBJunRz4hA5SosoO2br1RCp5KTfjg6eQlB5MEEA2G6r7Tz5qkXTZf877vn/7ve5GfRAGGk
0U23wrMcv97HbTExYdi5oxjmy4/eHxS92nsEfIswDaBirM2ahjhJb3wQzabf6IdJtAnu0PMNmMg1
WlAsbEgdmvCHdGnttEimz4UXGA+FShSpbsN+2wW6VzgJwkH67sCVBV+IN47DENq+yDPcWvJi8wTZ
SyA4ZBEvsNN7TxmNLz9N2Wyh8I+ynXUzGC56fbQ6d6ZlV+jWOPeL+804JhtHelkAp1utr5Yrn7zB
nlL1qP9ST8a2aP+pAhndGGRTPM89kjvICnRlJ8GwFZBk03pwOnyVs+MkZmCBMZ7HnFDFJGIQbFYZ
7+kr2vZSDixbsdeM2P+u7RPZwx91t/x6R7C5oH9RmIdmDIZXl0UJxStueHND1ZVPl1BVOo2sadzB
h2V9NpBV5Q80RrJl8LDpQ7D/k5Ne7+7Tn1aUr8KPrI3qd+IFgYrZ8QvzwgTz8fIAmOpKyuInmXzn
3h6lTrU20ow4lPMsXMKMGoAXNI0temFk3r5H5PGg4uA9/tqoiT2WLpx349KxyPw7/RxqWfqVdwyT
B+vzP/IHhfj31So6pK9uI2vcq3S44x2pI3gsrmio4J1Ab5p0ox866Qd0pKT5nh+wVKJt77C1fjTV
pYEUVHqupyj1jz8UwDJFXSWlzfmHlhYOVZnTPVbPOPpT2F+8mRFczXUitKaK9ogCfsEJRj12Wqnl
qV9ERwjN0VZ/HYUpxh1HG+AFtDlk6DMiinIoc7YWQVq3aTx3o+vQVwWGzmbhEcCboo2m5zJHIuWM
QMqDgv0OPZfad3YLmhBxb611mC7UuR9pEApsD6kUpXOmmNSvXXA1GL+saJBGl/CCFb38ePWrbHe6
hvjpsggVhTjzFatndD1w6V3Q9da28KjEDJvIQ45uwk8fTApHd4hbN3aTDArsY0H4j9mI6jun78T6
U8y29v1xfDMfvoO2AWM7LVmNZ2hJnzMbEh+9Onu9l7XGhHUvw8vS5ColjxjaQuxrA++yjca4EmRC
NpOeKAGEitf5vONAqCXtfZdC4iUIPZVeDgMmdHHlKk/jRpLt4k5yS4t26DIoWUXIbfDAzTL1iBUh
eWyDuHhiwFe+eVG+jMAOjoh5f0+18iLbsdxH3IlUyiew/MEfoAEXjlnlKKdp1ARW8YylePtmrwB4
zoFDgCHQjNrnEL4G+K7yNywfG2s4Ik4JTtT2eI4L/YGtbPocm+TTE6Ednv6FwLnCFWbUO4lmyYuv
52dRFC8DwngtCffPqoPHO/zWniqxD4O7Ci3fAtUdvx2bVHwhA8FicQeI9keM33kZ7sIH1bAiy/GB
gKJG5H/vkOHAePx92yg+TO9sVSWqF1Nxkpuj0FiAsGDsbbWF8czUeHK12Ln8okSOvtnZQ3qJJq6N
OONdDqEnxckkKjxr9Z5DjLu/ph30w73NjheMgMFol1RXJ5dsJmIyyNGi1+ZBSCQPjr36KVaTlIoy
a5mIAUo2ERT+X6pimZWbtTGPLYU3EhK3COrnxZrpF2DvrB2Q0XTo5PqIUUANIyW4mB1/UQQH6NMR
R97OBi3ZE3JholtHvvoRuFLJlCWudchwKA0QuYx0fmzOP5iJsR9zPbeg1EZgDkjgI/ZRT4+qfS49
+sK/uWZGAflH1dkQOT2PzlincRNzgCSgmwwM/lbgvJ5m8IfyfZay4V+oOoJs8tYjpl4PtC4Pgltp
xDbgbPUlcrXHSyaC79id8p4WhihD9uHxuYEWgU0HJzjKqfHkehEQ9PQl5sRBnQBlLx2ljOokjjMt
b5i79kWmJVExX5v/2QiOD7FAGb5B1yB2HNVamk+UD6j33tz17WZiTZT5kEV/GDPghpEXmS9L7T4f
3ym27xbXHNhBSHDBsw9X3MxUxn8iWmt2kTvKTTGfsZdSo9JqTfAmnLMicdkQdKLhxR8lQy6WPm1a
fA09Nnp5XtwhodM8Y6N4nRD3EC58QdTnmONniIMLVFA9w0OF6bYNyzOa+8yyjrrQpPdshric+SLu
UUfhGVSFQ/W5FOCOo6OSTTQ7NAmsDN4lggIPXbH5fXGmjrN8+aFn2qFe0AqwPpawxyR6GolA/xSj
bUoHQKGnOcpIqG0qKWVIrB8bqt0ZD2a5cw9j35XRgQWFi90cQgaC140OgZ/qWneAbCbuB1fp94ee
LZ2MrZl5697uqSroAjL52z8yN0vO4Ypxq3kMzY988CwKIWEFOlxJxDc2HP5rZVx0a6JbepRzRJXk
Vm18FO8gWPyE8jQ5VIsqn3Hb6gq/qt488JaOc4/tZPEeba2lAFhoiwZs7s83Q3JpAVvZp6XsOnBW
QtUm3DZgy68NTC4Fmek7SvRXrPM+W9OV0pZBBn/KBzcdKizs6Q4j+l9RDv5pw8cLFv2iOLVmqh4t
exCsSirnL59dLMROGJXJtmRVe8o5DKrgVziv2YyEye6qt4L6Uas4869jdg1Lzc9TPgI08EzhYeXq
35EQJMY6mInF9CJ+1kmrmdcheJk4Rk23s8hcgjCecQMq4l1hcMHm0lAV05mnY/Ng+hVCeOYrRx+W
JjH9WDJlNXMlTYcYSINSbz8R1C93bh6hEqXmqISqQUYHjkv3Xs2iC9cNjTQUKf2bCrw3orYnu8ti
1TMrMFH9ATrLodaIJ8/l3aod4SIIZweaCVs6CszEHa1FAU/HGu6rNWodYWD7ckHDI46SP4GtVtOi
O5PIuCu459yB2cW2tIiUjYJ3sctOoZEcxi6LhqfRkYWamAkg/pU3QglY47l+eQpdOJaHvubh2BAg
1F5tawV4+Zmk5RjVusecV8CqDfz7bIoQwDELa6F7QzZGydqDdkiEekKDom0AT1JwN79XhQF19XMT
rwyJBUwTjeuUK5ne35mMh5xcbM3EAWrjjaJIjW4OSD8JpdPii2ItNZWByPijQDI8xwA8OUvnpak+
ix0KQ8VbL2+cbbHQbRl5+XtQJZFRhqBDkLAIVtK/Fau7iXB08hievpXmbv5diafJIiq23g/rde5g
aiLsWToVClyOPoEw7Y2bsAp9sWBsK0N1jdDmgyAQdzqsu5CU2mfMkefv0w0B9AXxICoq9bHif4/X
RgbQzq45EkpHsVGzX33Qqm4kntwpTQCEO/UPMc71n/s88dz11IpamE2h28jmVjOzxNxyJDigSqJU
yA9mYbSCjfVuJwuVuEDHJpNcVgDgDHwvbMg6Vd8YzWYuI+TjIs4yCs1K0aHp36awBNAdhzs33UAV
5z8huSfhVeasZ2sGDWxqBIiODp52dRjHwFPrtLmyVnz1+bkQIigZ4DkLv6DfB5X9v4AqIlW1wO0f
U/5f/3igKpz6M3hhYs2mcAb6052VeWqvjv+wMoFUOfrgHX0Xl0rPCrJ0MCkNkTDuisPjfjezzzpf
hI4w/0KmRHleJWlKCWdDMcwksT7opyyvnxo+2YKocPY2Qp+5ecKv7RVyMx5oHsUSfxYflgNG8uwU
WHLKIxzfWncUlLuLnPBEoTx+qBQVX8TFmsdT+ZMVNOqzJxCXeY/Zv8kn7VlbtMQmBz5G8uEd3eh2
g/NeVZOVhofBMY0X8C2OZLyUHBKyIFLfjXqfsvtA/yZKvjhkHhnRYQYhXJUs+Sdeg+UspKbOvP43
LvxQW98HGjITyLRaTCybuXR8xoaL1LoCpRuqHb+Fm5WjqgzxpFYGDj9SnnNPjRk4Yd6UuXn2hInO
JPJ1hnCeAMgl/g9xFiU3+Ep0c7ilKZz3rOssXgNLbgcf7H7n8wk2mYpgwRNTzSFep22EhQUPCGK5
axzPV3BOSIb1DGp3hiMc4xpV2CG1WApqNF8WR+wUoEiteF4m8e8OO+36HEf9gNZW+pnwHMEe20Vy
cJJxI9hjWgCBeZMLoYVYpPsA3YL7CdWrSA9oZOlKhfP2w+s+yfN2nHMy75JTHudm/rBAjRT865Ax
0NflTXHHapgrDCuOCHyau4FM9kPYbqfuy3a2k5Eh3sMLO4fuu8tF77BpdE89pK5llN5aACqJYiLw
eG/jAylsXT0ju3U0FmKiK4ADtkXb9sMGvmS52vZXkfJctxJiW6vcAoIeJQ00f/kl/A4rcXFDAwFM
38Czs3CNAFyFWn/qAa8CfeQJlwb1Iv2t37MW0P24XeUHiU/vEWDJneQwN5hMOwvsVoY7XwLIRXCK
353fs8LgCFlRO0OXTqZos++c7ocGnBkX4esQkDtONURUpB6Ai76F984pO8Y0QhPt4IMmN7n8UbfJ
yFWaDY4eEq38NEGdte8aXQi1xxZAad+/Cm47mWXLumLX3yCHxERi4cDptiRaVKhTPP77kqs+2Y6c
mxJvJYPalNfltLk6ukGdqVPCD6H86846v2TIUGE2yQHHKZwE9tw4zakr4Sm4KsSgEIjt2L3kT3qB
zpKQmnUoSpoxbuIoohJdbsBdqEwtrmsPpy1//zOtWsO8WhuPHtHhNvCjXZFm+DLI9uHR436n/w1V
/nCTBuZwCVtVnN3VbzpUrSfzqKBd9r/vbZZOkJ/ownoXe4YziXLcLkzd9FmKI96K85WUWChaMvLm
mzrfVYSbV9yKQFWYYjXM3JxzEgTSdgb99BvdQDQftMMR8TAbKkRue11HG/ZBiQ+o2zhMpijiAqJy
crX2ezV4z9KAhxNlPxr1bz97iskjcqAEINOH+dgdXIaYReaJTKSeuL3jDz2yMmawe0jYWWuA8YBE
25PcU8DKvuG7GsLBK/pUjTspscLGr82pcLvkKQAIvlRrRN/VNTiA3LB7WXhZDj/OEIT5lounn5wf
/gV7E/9jQsD3BbRPF4+rl2bIaPGmymKUHlPQL4pewDbZ4SZhRPkHDDkGVamnSSa0EydI4FE6fnXI
HuEJiNZVseTKXRSUjIrvNL8n3N8wn/tqS422BbfmkCFeGW1vgdtVD6BE+C86ue+15xfjFmfGLtH5
Cl2WjkWiMNy5iGHaesp9WL+BODDmAI0w1fpbjUro7iCbD1D5edCuHbWt5/UF9hDWI54woMc/bOE3
fwbpOmmHlKHGXTMlw4G2TucQ8KW2PPeWIEVvdvhy6CG36LjXtaeeBZmQCCjp0Yf7mOA2qxNcXNSv
LY8w8748lTPCx02LB4L6wxnv6GAi09IqeaiO70RIGgDAGRv4EyxSlVMbfb6xv7V9n0AKx+lLRRpW
EMLTcN6alona5pGpKFOj+ev4NgrDr9cqvbbNTP8mLwMzHnhGtzQ3yNAz/aOVHOhMW1nT6rRI9epI
/RoiQ5DOdS3Rm3gMAaehE7wfr2gHs7kMaNnt6Zv4+hadiUAdd3U1Q16VfALcYH+LBcKzQlNO6SXT
YL6hK/VPNIVAaB0heF6ooYk6+b7cvzWfDRaGkTfdD8wIFx4Ybrj9kVyjK9nFv9KTDZluGbnPY8YE
59jvzO68jo2dSo5qn6l4Y2GOjLmVaoSGMip/SWGB0fpcr6F6m2UGyXArPPi9nbEADtLNejwiZtK2
9LK8bK2yiMndNWQkSVfnnNXpa+o1RtIkYXPAphQyW2N/E4gNwu5l8qUV+zbCGf9ZZU//lVPaG82g
k6a+HqScNgN2QMQOl5UyEyPPG0k7aR2y48pGjNU6dPIkZ3Q0oV//XJEzBZ40/SoiZLkJ1zcX/bxE
PgVYQH3MeuKJ/v5YrIcZPDY5oyESyJQs5xEBpXR2yb937LvmzxagogfuBwO+l1lX5I+yN3t2Q4Pf
2LPqHWIFRNlJs8vEfg1PvEsxBCpurdLdJQn0r/RSzo72THc42veZ1xjmNGvyYf+hPlY1fT93GCrk
+Dx26NJFGkVUGGcgLruhPqAHjXDy6b8/wpNhCJ2zvslsz71zA+C8vmlOgHjIg0wnQtHr2RKGEsku
3tydTH9fxjYDCRz/NAZaAR+UY7hfPYy012X2GPk/td2uzG5VQGS5TJGu7FfTJ/cVHML1VAJ/AWY1
2Aor1T6KxqlWNT/R/H+0SdgPOe4nIP0CDkYnzhrMgcnHXZsKXdYBzuCW5siDxRpA/469uOhyO14N
/QVUAfG0O8uPJvydcOPbSXBD57DLZbCUoa0h+JoXSdQ3HjrRJbc7LqJxorlvGl/ME3YNPCRgAj8I
3gZkUwdEGAtawkhQrKT0ZTNkjci46s+PDsQIa451a3JrrxLGl/kppStyPHyfSSzemLFheLE2H1cS
U9YapAm7hqOOOM+Y1RuaGMML/4c+02XFfLqELkyguRMuGbMA2JMjG08jT1E5epgkx9/EfU8+wue9
ezojRteMtxlEcCRGzPdxjKNl7uwprsQvVOsKp2HPHIrTSUCqjkVfTzPpSrM60x6Ezy7aOPNRxe1R
Frj74+Fww6uBPjp1Hy0VlzkuwwqeCUfnkbKlH7YcVQVaawYvYWnGhHiFVunPz/R0fiLf0Qmqocbb
KvzC/LWj1q/ELaT/TTgRVfC1prJM6D/EQPUis4jU4A+Pgp/UpU5Bp0849lvjT/bnwsFkBgpIAazZ
c9nhlzMp9ZBEYuwWJIBSqCAvT6KutgwJjVyDrw2L41SyD/XiKuJ4RIGUPgwADdHPZ20lgFqk9vuX
WK1dENu1OC9FhmkiPv3KAwYeyX4V7rXjNDTex5mOd+a+icmBopV3GTgwMoQDLmnfcu5vaO1OXAQZ
ejTVI/Rtx4bZ4M9AjyQkx9yJbR3bYsaBCyfGl3dbalu8ZFvg2yET24l6hNKWTBe71jq345QFBBL5
+Fu0EpFupc2JAHlpH7ClD23dLxsH5SL1BGrAn3GpR3C7051hPc+3CuldGDSbhF1EmAGICqs+HP1c
plp6Hclozqfy5lE4o6oQSeji/Isyb02wIsjiT1f1fxJJrOIWoUVdtU+3wGZIh3PbrChg09EspJR7
pHHfmaUEiTyM4GS2QaPhIgytO7acNtk0Fi6p9ZzvzkLsL3zdbYJcaAKdU/b0jYk1cs4Xsk9054qn
6z4Xs/3VKl5Su8wegqdrDFZZCwRGe1aC/RDInymgn5Ba7qw6FFBIiLxFa05d118RUrxHP0FaTMWY
t2+EBDUaDMi6UXUL5nO6Ua77GRvXoNMQnPuTkx7vluJmKU+KtQDYMYja7bN98jZzxgK7nRlFmbHi
8QTQ0XdPFYx3prl7cv+K0cqPRhpOC/iKY0eTO5pDMbUdQU6p55mmCDCXVAkomynNNYWzGROmV5mK
HfORpBWsjD/iVpvCMmbk1JvVGjmXGkj+4WeOt2tQSwM39uQ/JwGgJcNKNujjoXfeJNI+ReMaZwr/
v9kYcGmuAnn7am7VJJ1cMvEs5oe3GV7k8cMn7z1PJrsz2tiC2ESFpcxVvTCVNBgOXwf9qsdpN9K2
aML851mVYUiFFCmRc0xr3OiKEQrNlvhAiXCafaASYFkn0y9tPDW8IabSk5Uf4CSxZRdAcpRosSgX
5FJ9HBv0OntwhkNQsIRoFw0jM+YYdelcDr9AB6rBMxPBZ87HdN2Orooka6JXN8BuudYfO82fuIuc
IJkXo1MbUdUyTNScD2gdrqhU5k+tDBSUWE9bGdRu3cZAfHx0+Vx12jqsl8ba7bvAq5clpPGym2ne
kp6kFJzlicZKEs7P0S6fkPHPJMk8rqXkV1T9Ul9/LINtyafkJtUMmP5sxF+dvhcOAj4Yvml6dEvN
7lxCeuUPFi5rJJiLGQcVZNLVk1qkTPE3mL14II2WV64zJKZ+WUxjs/2Kis8INPZb0MdK/HZgxeHw
25t4QkPZ49jdHx+Pxu9PfUYKohHK+aVju3fkpCtGhOZkrwnzvrafiLjHg+5a5LfRYikdujAzBE3n
v5rw0f+i9nPQIT0TDfj3XM3K04tvnjZp/fyAiaELETVYUu6dqaZMnL3rgSl9daGXaPiomEQCi+/k
ITD84t3xrHERQmCmLJNIj1tReTsBtoKwV26ljtZzm1FN1Lt1na/LN7+e/fpcUr9dGUViVPdRIs34
QJPbIgdJdIgXyXPlAktLBSGS/0Cfu9dDsXFcFAuNYFTjouHtnCgSXcZtFLR2BfcCpJyCw9WOSoU2
f9CQbdVc8MZECqXrFIuW0G5/0UKWBrTv8B+2ALSOoHuGwZnJUF6fmARgkOIaJ3M34kzcqbzPu2jH
nIR8T0NBW8KhPlGPjHuETdANVV7EAWRndGLmguIltvfSXyHywUowTCqVBqd2suc8ckeo+F/OHPDA
2qe6Duc11ssL3y/Q+nOjLx1cCMqa4hkQreptJASZTMO/LlGAOqcEzrAjf0iaW1m6N9GiO5ufSMwb
ufNoVy/24qKuFnzaCtYHu8Eh2E+NA+1VL8ghd0MnFsMEqLjoameVafL1xE4LaI5HlDUQ/c/HxG+r
0aIxfKTj95ysANnzUiCnYW6lgZohlCjcl1a+HppMZ7QTh8S9O35NcHu79TCYqbQBc44kO4lzCF+b
G9bhDGE9X0TTLILFyWqcpSbxmEFqODU+g0Wli1SlVjCvtl8EB5sRMTrbsd1NlNUHB9XXhfXnM2ub
/OX3AyFm2Xxrw4dHJ9v3MDAS/XLmpKclbG0rqER3Tw7fI6otGYh+c8/FbuoBOmYT5PNHuhLJWh7H
rU5yvBuxsfT1z3mt4QwZGZBInxETl9uBP7nNOcziZeq10lkNZg1aIRS0RrwN4WZJ0rtz7mMnp2W3
WgTBdcyzV0w6GcqznoVUTx9TIxgBrbZZ0ACk56s8IFP65OYjtlLGX3zorODqRBb535QxxEqumlmi
jVhLsIPoxmCrUcLMD+MIHPE71tQvZOw7PoOF8I6XQpTeZ85JS0LosUrznAYJxQydSJvW/2919YAx
i3HlXzHq99SqESFYhm13R9B21wfGZPW0mhagf4u9rAov6D1bsOM0FCntenwwY+x1rnWoDxfr+hS9
DhVougd0AsK0bMrtSULdV8N66f7h4srBNHSp78rCwHvghArVZFRC74aOe4oMPcUQGFWdkIwxAika
dMc2AM7vngehMj0BX7kbzPUHK/n4lZbnP1FXGbEBO9Qk47s0jkxeUg/3Z9+8GcvKZGm79m+sKYGX
DzlwHc0NmVjOO61MhyIWnXKz2wZFbkPbWNIFJccQsAJ1xXkxNXzU0pdbLyqnh+u1d9hmGZqmeuxz
n5eLOXoCUn5RPqIc2FkSbxvuvCSeSwffErxateRHnZBaArIDRL9lOzPOnJkmHASOFB+sndMS+1uu
VX5Q37nDYBiqLNBHVQ10VfpBiS6kTQ1bknecXg1XmFSHMiVLicdx2S8yuq97Lw4f2HNjpHxZ0SFG
gTYV5IO3TefOxRpKqBjT/mnCJcoOQlyU4Fmvvyt9IYk+pInn2YY/ZOZps24r0mAJbrxCIWbFWeRU
5yRR0EHanI44fnEEezjoU4dkS7ZqBm/J8y4INOujAmwG3zt6bDQB9FM1bInqU/S1AZKxp9owtswz
ITjWmuPRMZUK2JnB18FSJ8UEBcXRlDW3UKcyoJk8b/aGLnKbl9qQk0QX/kjPnWKkJeGSWUx0v7am
FU3vjU7N6Bgh0pApWTcwch+u8W4Dg5/35NWf04S+WG11ve8dC9zeGQv8IEKICfxjTa24YHGGc4gN
X78/hWIsGBDhAypIcOXpVibsCuR5BahUNdjS0OwcYLRI0CbnUUCchPq9N1xYNBoEvpV8TPCgmUJY
PlZSC2UA0+OjCoW2EpkIaGEjQYXE8IjdLhy1BLdWhN+U3eu7tvppzL85fI+dACCUnusB10jnlMaG
3jJCkRE6VKJHQG+2zv05vI49AlKo6soAZolvWgdt0fNeP27uPRYn8kRrBWsVud0KIekJkT76Krfp
g0NhaPg51hA86zE+dAev5XTjpcPjE+i32TGhOCYLUscsPWSP/pdyTnlde7bejaro7cippScOEjTi
oXxdsnQ4oErmDxGiAynVMN+a4oBmcrM8l3hdKG0hepsykCuxXpZ6iqewnKOlAmbH8D/CLBxa2AKP
ybdkBRDb9esrsKw22B1LzgHRdBkIAmLC22IztPlk+bIf430dWg5ePUtmcWh8qUzl7f9e7SaPA2eJ
ZOxvHaaIAlxJkkwJ3NhZ26R1vJTgx+a47a+z3/eMDJTew7Zm1JHFR4zr4kmcD4fcYwu+Q33JGqOD
zFniL5ZLNK2B7yaDIjxIVLCloi3UQqkh4BHPDWIBBVokRqEmJGcwuGNl1i0gMOnj6qPzibvKGlwP
41JrgimqtTHpAf6kVizrwCTpYgMLbV6TR2oCFD6Tjf/0yQrBeRfskuoJ1v/0ZHMkOsuzJ4liE9yq
6f77ak8s0OeFYVMVmcmM5AoT7rvGX54JTZAiV41B3MhrZ/ZbsTPN4sAuqQPE6PRHdkdebldobHKF
2JpRJbotTNh2X4+1cGLluClp88YlEA9OZukEfUhUMTCivkywoewDpRNJ1/QyM3Nq8t+++5L2aEuY
z5u5Q9VhHV9EbW6lUaDZH/14B7CFxLjoVLjwh2ntOa/HFWkRQONd6NWa3lv6WEikc1wxGrvhyGOF
s4jjvALo/8XCrbvodIFd5/eWVbLqMus2xlE/Wz6Qfxo5FXHGjuFJoJxrlrh6Dl/nf+3Uj7w5zF9H
AzjHVTjYAW2HeDJXV5A50tJQUWNZNDa+UTpZkm0H64PlpGfUch58r5jK7IOpfxO1+DMwV/T98UUv
BYb3HtrL6snmxxWKEeHFfIYEuEPUqHSHI4Y4a+TqRuB9ObVcwWQi9OVc13XudiORzt5IwTMbIWcl
c/57yKd0iF5+E7cLCpxlisDWPcRcuotzZUevAsgsJxsfIHyqCi5S7T3fDBeCyZII6HzlBt4qfunm
Dxu1cSIfdqh1P84Aip3KFZ/ZYIURNEhQ4W52bumSqrtj1Ec7yVkuKsAPeuaAsj5eTnFhiI4ZwO8E
x54GotH3tm/0gl+2dqrvieBsrzoRIOyzR+V/gEgvG7pOKFGh2bNenNY5cuTDEmsBuKom7Q9UWBsJ
i7lHnbLZkm6scQ1NdJ/sMyEMHXncInSmUb9engiAxxXQIelv+9w5lf8aUBLkwyEkNHjZTuWZEzx9
+yyNT4rUzSxXX1fDIFCpCAGmPjKyi0Bn0DXsvjxhj/Ed/69Hlm1QRvp0L4r8+5bFV9X1OxKHL5Ru
066uk7fjexlEC7/i0vOfTlgPCv1ZTG2N52ckCh9pHRzal5fH2Vc/SsWupKJlwkbXO9gG7zWlUU4m
A7hLQ3nipjECB3YAeYkPwSaRwRjvzI0rseL6EpeeOxWRftw+ciu8UJHvd+f3fRpaSTjHKgbkR7Bs
6nLnAODir8M7EUbOnlrF3ChmWRo9/d5SIzqF0QInFHOd+S7V5jvciVd8O+RS/qAKymOMuMnaZYq4
l18U2s9PpV0NPNV3i/URd3hG6P94Q5tRxMdf+fmO6sxquYRZotR7yyOzuTdP4+L8FOD140bJVA+a
m9SkAHzxxO1rRuqSysGvpiEClAi52UxMCIPOln6MCCVLBod1EGmRKX0Yqwa7CBW7k+wcmo/tMR9a
N2051Nb76aJ/NuD3Z6WzC7JBg+HysEekJvC8B+WKnzKVZO490DiKNWfLJrJISHao4HOJO7XnbNoC
HFxYgsp1SuH57h2zqLXHo1bABPi8jCXZThoc90/Q/yzW48TfkIO4PFem3HOMg6IXK+vtuWUdVxNP
GOffQFctuvWStH+LdxDC8oJfCrdnzZWB9UMBMvRy9RHQmk/FsCitLDrVyej5mwJviu/sN4Hpg0y2
37FMWy7LXhmzxpYMFXy97CG5bF/KLbKb0+QpN63QdLP13WN2y9rdEQmUUN7HsG9SkZMZmVxayUwP
k08Q/ximiPxdg4bVH0mJrlVIKvV2RgptjrsdGRig4veXD8yTgrQxL/XbSgz8e6YPne9Wd9mLKxIS
/c5e+zegLTHn1qZpA3rapKAkRMnsFxAwRSDp8k8KZePk1YKfmqIZuSgSIdJPaufZE2FtxCK1+akD
2WznSy24evGtN95cOZ/9TqLMwYlRtDM8I7BXxUFSgq7b2UtyCekrjYrHDnmi1AXTy9uyDON+L2N4
npoB6H5ZbuNRwa0eNFXSvsvUvwpHjmBxesyU/WGZmeC9CD1X+N1yny7X1Q5pN/7p+psTMIZ9unib
oCOMRcE2YljxWABSzfZeF9S2QX5GN4bN3rYCOj6x+daGy6kOjfqN1ZBCAsW1fnUtMhgwp1qWsfPh
lT44mWsM8IMVrlr1wGqhWRMjJg1KvRfgrYufTrvjQyz2NL8wEbKdUH/d+pL0mn7fr+gEdCr4WeXw
AQN24OOdsRAQ9iZdeHunTH1GnJaCwfV4vnyylaXuzdEW/MlzcUmJjxDC2r0pfAkCKdOMokMH3sMT
6h59pda0A6SQdWFmSEECSJdl3nuiRUsn8intDARLbkNFUjuVMe1Fq6MtgMj7RjFWBBZwKiE9xaCF
xDRuyHnS5Sg6Xlhm2dg3aFYefmRIsVCK4syrfyBYVPa5hU5bhM2DwvhaDEAXOO64ObO3K9cQQmBY
YrwbqwHGCA9DodCT8UresrsbrN/E8RWnJXAx992UkgTtrRjyRpzSVyCz4afsLp741X02Z/Fi8UxM
2Xm+rdfei+8ljHyMJ2lZes2evT1bxaWHWK9fm+vwGe/O/iKphoia0scHymNbU4tYoe74Bbu0LTlv
K9MES00ZsEG1elMF5oIbvbsK4BJn5XXSpKbS8Ir6NDb5e6rHKBCWDix/RV1cVDq/zNybVTmEGzQD
3YmbQlH2Ak8UP2LG9Bre1m1ae3T336d2JX6eObjU017tRCtYhOnmbGdKuGyvIGD7plCkwfNAkS1A
b4BZG1D9Wip4AVCHC6ekWyp2hdeQICNsPoqmBsrGJrm6fTzq23DOvnRUCGlCxDLNE/tGhQXuDE3U
UJ+9YVnRQozbL+fziRPq19Brxp7NCkTwQvlDS3LwExxDHEFCZ9c2SE6p8P02zetFYxc28DR5b2eH
sM6+EYFuy4icB9pU/t8rzynnM4iO0WtRUIiW/bF+/UeyanI4JBEaKm54QL/7/3wiK3VuftPSwbKD
Wj1sPML0ITJG+jWkGoNrsVEsqPjzajGVeESOz9gMvGqrU01GL1Vl838LQrOoad59dEeQ+NbGB3Yn
jt6JSxGTh9+L6P7A7JaxtKxsjpaC6q5Y9kxSPJDCtszuzAqeLEAk0L+OUkjGq2dkYcA1Rjp90tKH
RcIaSku9IbYIKxBN/1MzZgAmToMvnfnIvS7uC1hu0+DRGlzl41Eh3ZrrNRqhpTdVQUVI0Vb/LCHZ
j46vbpJOwfYRHhyDmUP5TLNrfEICiqf1kGSthALhevEtNHUmCbKghm3mZ8Fxf+6YCEduSHSuAxi8
uUWFW/BtZaKgcX/HYScSgM3UqG4IU1i1m40sWbVRdEICht6hgdUTPlT7e/Uc+MtwHUgynwdPWzHR
FJxb8hdzjZOy6CCiSPcj05dhZJclIC5vaOl8miAHRsRoqqSJY+Q1cqrNWb7+x4Q9ZHPjq4SZ3nLS
IEJcQYSDnf3TWF6pVq8PkoGyql3SZhqmL0xi1OuZPNmk3sdkinvufmIERWN87az6zfPxJC+z3Fce
BW7cYxMy/Y1cPBHObF81cZAiI6/TPSg2U5TwzrQUvGye4fcCflRBr58p2Dfk0IDN4S3jvzhXGKLF
Gnux+1wGxp9TPdAosfQludGsX11UoNeMgrS3lp2yH3U7zAIRzF1oYiSSszMbwAdTHarra3dXBMk6
YR/VOnRIcnh/Bx/xhBIZCjzZDNFueDGpzYdkjVJ00KOGF297RExVDhYmuXOxYli+7vg+CbXsjD7y
N5dfVhhNBRhih8ASpMvTR90S04hVd6gAFXqhs9RVGaTVRnhiqupJhhq3CLSrdSX6iABC5b4BHCz8
tkp0lyo9HAW+tPIlcoW0jLlpKKQBFr3cw+noeZu6TL4T5LEqyPl7+wPcHQQ9LMxAS0/uztRlqh2p
5D41cppUCo854WMx712NmjSNhuYUs/t27m+l2lXddbfcWL7jmq0tbSxiFyum/QEoCUmrUiAiOJe2
rxW4YqpNY2WWUflZixEX5Mu43Ig7GCUIcg0BJUy1FdXm9mpaBJgaPyP/v2O/HqICqLKNqY9JPhh4
RV73TxAYBGhwK0OJMyHtusoYKw5YVyq3CGn33vKzfwoBQDTF+HIay85GSFMblRxl3QdsbvLej88u
+S3yVm0L8oLtlHlds7pSE3XrTuym/v7hSawIpdW1gtcCpAnNzAKktL+wTbT3vYIkLP+ahPcdzgv7
Z+6DvAmUbxfNoCX/9iXq0Po6e17IadpgMMXlPBgtRYFMHo6E5vT042M2F5lXHip7t5f5lM5XFQTC
c5QxoGJ/afwrjrqlfWsVpK42Yq+cXlL9Z8S8eZrFBJnG0xb9xAUALQDwmj6wbFZ4C0F7fNvUfA0i
pI6VeU056k7lSXNgSjOskuzHA3a+Irk3f+d9aoi31iJ91LgUDaXjvUrcvEPAR8ZIs3H7xll90fpd
7he7LvFXKWJBrb7CHu6eywyeFpzw3H762XqD8+/kcrOyxgZxyIr56mYmlBrSYqWZIeymCvBfwuJe
ZKN4HYSlAlzN8V1hR87gwsmRYru5kw1pkfJezNF2V/mq42aANbnK7yBrzmPmVncOQ2wsb8KIf/hr
02+Oys+YbJWy+ce0zur+nNhqClRd1DL3FvlbNvySmH4GHleUgryWDxFjOJy+I3b5BEZdDAGYubM1
PCWM8zRZLy7KYJoetNQrfqWNdt+PwEFmIzYx0I7pJf4SlIeooyN61DkLFvw1m0yp64AmNiefNh7o
f0ntqqlAX5ks1LJzLsuKOXcRB6mDS7uD7fNF2Oo/PuKseSVasR9PtL6ev6i0nWD00z+doEB3KZ4o
AQhBWdAywgitgu9cEWOU25mfp6A3jM7QZMQ4rDXDhIOMqH26dA66YWKgc9WyU9Yg8mU+xiX3D3tW
S8v0LpzITbSP+UgAn/VSsDGn1QxcvfH7KKNY3kD1tdlE76E48HHJF6v9fXZpfotKwnWU4d9PhPKy
ouijOxbKg0WnUUDMPd9iXOOV1JNPE6QBjfPRQ6P1gXvWOEgtCoYge2VZqoit6owcvreGnH2YNxz4
PjOuellzJUCla/xZTki0q5e2mI5pQf4UM9qv8cnztpW21mtZrpMoIocqMB6SjHXuNM6cgztRglhz
5G9ApSyxc4b3rLGCfDtjUGHeguXB16Azmn1zc9t0MziVyd2zJkC5eWtn55Fo4PzCuIzR1fDCdPjH
IIo+uN4cg8r5hBBbwYcFwd2T/5gh2Kp28cwWmKtjjISNJIvVSN+RWS8X3dQw+i+ux6E9k+zZ5q8N
tnU2TvXU0I53pO9XSG13ixLclK3jFIptpCpjdL6cGELFOmkjBXMmBkXo0A/o5YMUqp9gnFUG5zAA
U1CEmO2CzQqS1DaVkW4qRw1u1pxgivEjCTkC2zFpZGC3m1roMnyxXxkAdd21sTUgJr9rkjovbjxK
ESG8xUnkzTNZS/yO9fff9srpFO46U1qM1mQhnSXyjql0k8O6yliGZmgjJ50UhuTn2u0m7Im9VUjI
zHDN8gRPYD/uaZB6CB5u/RJCEzgaHe2FSfLfnpkf/ZWa+cT2gOmIknuYBvHb4Y8wiZRuF7ut1gjB
ulc8OmSzOdGkKvFxvsuy3qR9lhUSm/XDPcZvn0speN+aYvzMPMbiVLmb+N3Ndv4cgjfLTo/epiap
qu1P4gWsRAih5GUkfFO1kHj2e9fDqnDIkDqT44nN/Y7dXVwMX63zrXDueXSmXnmR8TgaYi92m2gL
Wj4yMOsaPLxemvUK+vgryDK0aMpqVwTlz9VXmh3D9jUHAlFG1bd3ngN5Vg59kSJ6/VmrIVMtAX36
F7orLZCLYUPT8azdvrHsEBlpk/2gITXjhHT/vnDr0rulXkaIjzCvaPQy6B7jaiuqW3Wzlf1XXqNv
7Ur/1T8x+R4Qu3RnPqsj8cwK5cLe6RJrwwYlwtz4GCHJR5inW3aYJmP3UDTX1oSEgIIe1LJDS8bq
C6YcxChyUcTqM84eoj+fBnwDo68GOO1KMIUll5QSPr5YtRVd07OYjUskjjjrveFtRFxgHKAVoEC5
0jbOGxEICbvo12xA8sd/+5B1M8nWbRgQnP+WoUTxNj5zFK3fNJx+qehbl9wg2DyS0DqdZcQVsALG
HnmaBo1Y01pjS2XRDGy5yKTHf80mYDDOJ9yHvKR+e6AurLKZmXfJUyZ5xQAjLdeOm0UMcy9X/Gye
wgzlkBZQ8LmPuSXefXd1/KfIShq1P0Ya4h3Jup5HVDkvhzvx5P87uq8oR8gL1Wn4h2xCf/SDubt+
LKTKSVtn8hChnC9mO8B9BKljRLvlnYIjAsc8zviHq7B6WNBRvA7WH9bfmlmQrdYWBbCnFSLd5Yhv
GQ9/A93FZzsk4ZC1xB7jWmkqZ8A7IiTZ8wtrIFADtMdU6npMRl3mLfPF5wNT0X+o19Hy+tRd8XZL
qAoMfenkXKs7DxQzmVzlqZ9uRGHj37QelzTushkWI5KVOLs8oqwgqIMgoX4MXeuf/81uVNd0mxIh
qtYiKlvLtme9fKtADBKW6yu6rl4qZ2+3h3m3LIDi5mp6MOlghhKfTkIptE55vWEYmsm0wHy0Xbwe
oLP7oqFt2WatDvlEBsJK91h7w3GP18o77JesjiIipmmiXJxzlyzaVvVQ0ajg9B0CgHwcmGfkhL5u
KNRT7sqxt2PV5gwyDNxFwTPgRKEvcfcmHtFmyvhPQLrD5RqzgezbtKQilC3SxwFt95A7dJ1vcW6v
X5idAP7RC9RCecYYPQ9VijcLE0ToiI+BFsp//AIZV2vyDvrplLl8wOOBggQ4V7PtfCl+68Y8iFGb
bH3n5aRL+HNdX8tMVp+70nV6c9xj1n296xiVROW+1S/wzfwl3Fgylh01NcKgCNs1IKKbpK5bWRIZ
4AiH/rZZYVpVf8dP5kGZv5TbgardJXOcQGE2WscgUcXtk3LALSQiH0fxnqjsg+ZEugnmrShkSujg
AMQKEKoiU+qb59R3WyKoTwj08vgznbRYAXkUnv6JXj9KNciF495OddmouU/kpMnmqghQuHCyGo5D
zdXEzsAZ/nmTsFnekNfQ7mKR6z2aFjGmZxzhxKH6RhJu8po+vHMD9oiRbplQGEhDJABaTYytGRzg
N+de5Oylrm9q+utGiV+8zpYfzo9vmgUhOzEjCrPff1yL8hURnzux/BxFrDvEIdEQxnAUOm1zP8E4
UmQtXBSupH01sBS9jwGnyR3ZR7HHgZv+uWRVwBMs/4yFdkfyFu8+MwJpBZdoq5Ypw57mQ+T1eScV
vuqfPTfNPAgAdvMBeofjAV5bYfJzw+lCqd89MupV0SYpKkfnGtWEoQ0tanwN1A+QXCDnRFfu8lKY
XzZpK6QOH8/kGQ7KoojDC+Y2XfM0E512CZEUbriSPYrtDMjB3x+P20LzzbYw4P7lKKQGRocTyxoP
18bHe+/U6o6qCDpQEyD5je9XhmDicwPDssimhsdsRaw96cRjGlfIL0/VtN0D1y2HrHmSC6jpGEoT
aaZKHau170XkUKNT4tgFGPcyEK4ibgJj+Yzpk0OXSt973LitG+fFjmxqETaLZY9UyL2KRYnJeuzN
g7/bmkLawT9NMHn8W55LjuOejRCTk50cSciwbfJbvZ9qLq1IxyN03qMjHmd6n/2t2zBbDtwLDPhV
P+bPfRc+dElyLwXWustvtwNlKCrC2sCmOHHnzrjLNOHg5+qYkGzYCY22Bwcbzcoq4Jas3vJko/DM
t1Uw7cpMxIrew0hIQmd2nGtSScJJiRn860hHuhn4Hmp5UzrnrufaNnNJsmYUHFQ+c8pAEsL8PYFl
0MBc2w6fM6baVBBdGzvJ6ZaaAGEHLb+tD3eF/YviC1ZIFPHWOxoIXfviGPTI4Jw8hbT25866UzXu
5BQtbfXTS/IWNp3Fx/IzBz6wpQq87LjE4JP2dnbmyaGO+kD1ZYprwS/ZkHiU/as0muP/P2Rhmg3/
MYKZG1wK5JBBfszgGBJvdhHC8xmx90TspfTMUN3PVNMtGNmi/LT8DqowcF+vjvzq8qhFSkWh16Yk
5uvvjfZmiT6X2SsGEGWZqYu+RMZ+sDl9iMvrbexxvzF6AYn4bVSwK+DTe1PoiMkxDRN9Vaf2cSgr
0uObtOxiXjfxWcSOCc5vIS/Z1IOKv0ZWP9XWMdjmwohjpE57dPnb2YOzmMvES4PGv6HTGA55bI2x
MBFFNOD3O3tSY8kBm/5da2Hlw3VWIhrqBj2dYq44GDW1ums0DB+EC+ACYadEHV+ds5RRE4vx2Ecl
iVpBeoJBgY+tmk2zTQOvyE5IMJ+/HQcq5habBZwBISot0RakuitNxp7AC/Kysz/84tOkzRfL+xwd
gc/lruXbqE8kinTVOf0CLN+FF/ZXoF2SvrkcNmTMt5OH/MnmguR2vrRViLvYMc00VpwHUgtKeFTd
G+oJwoYZ1bxSY6G4Cj2mtfRljnRxrcbVP7pPp3+dcJaAC9UT953AbNFbJ1vkB9aCtjqEovouXsye
Us5PtwJk14RsCXHGOOjQVVHSBfVrRsqkrPVH5p6hKQ9NLQZUb6wpzyTFMFvReSc8fn/kCT+1ij9a
J9+BPkYDsBfTceUNLrzPU3jCxLgQV47d8/ZCErwyR6YsnfqRBnSTWBtZPC4JCfwgYQO1B0FwUPp7
oJShrqL5ss4guOEnlmov85lXBRIBtdwF5GVGdtrqypSj+vzLlpQq25sYLoWpyoBtnPBB2Rv/Nhve
9bTHnv/CK/DYHVXdv3O3rozBlg83Kai3cFZoxPxq9ZGx5qOb9oNQtwBttVPsMf36p8idviGviRGD
gmG+AjDp6uBunF1v3cPC9eVfit63cLhLN3GtOveDpQLaE4pBKLTxW6RRD1u7dBWUYzAuQl0FilcB
CMX1/aBVdm3uQi+BpDDdZcB6YIjIi4CF8xe3KxcjX1WW0/d0NSmTicdq3zgIyAe2hja703TA84Dj
rcaCfyvxlxEKQQ9VMbAWkgyEjqLy/W6wzKnA4gxD167X1EE5Sb2XjPuYVNvOTHKnrYHIGm64UNit
Fuz5gMyGEDXHRd43lWClIeH8I8LKmUxcDnoGMm/juXCInJzZX/7/JWd3jyaF2Yfz6DFIbzQN8gr8
kL3lij/gI1jodxTye7S7RXzTzv/8I+TWJz5DXb+P9iPgZcPNico90fRtWCTVVZFCoMRi2SI12hjg
6eCPdlpb6TuxsBSrCKYvNgInTtuZ0c6g40dUm0Oe0s0yMhcnXCSPrv9tueMS/u4SWKc/aQB+t3Py
4mmX7eWfzkApzg9/18HSk9Wh3TkLtJlTkrbaViFOqw0wvavUJ2eUFJPfGZXV0sqUV1o6xo1D4YgI
wI5QjvteYXD39e3rDE1ZW5CTD/qIsSkfSU66rtSKCR3ah/fiXUAYrJMII3zdI9clZbAgv0MK8ybQ
wCKhhOgZDbHveGRO8NQp3laXopmwyEpTG2FQ7xaIX27L7OSlcxy3I/gdThd56Tj+fzf4edd8mCQF
ujmJPtCQZTeJ9tm1+5Mf+79v05hrY0Sd+V9AYEPcylAKTnCoZdVYmSxE6dptUn2ctqZ/25h7y03c
I3ttjslFci+geIIjVLRAEkPyhgQu8hIt3wN4o7txiXR02JDBO/y+EU0Te8Pyk6Yf47w9nKgx3JmO
X0/lYMuFIrXSoUovjFqDkVNK7VJ1x0yKH5kYcqgUBPvj+HqrdhbNA/Mj4Nsxj6OYaT2lShUB/d85
ayNC4xsZhp09MdLi6iVr5cbjwd/8l1Xhi5fnn8OHlohW61rZ//lhUXrW7BDkNHJI6DwNajq/fX6X
w+/y/79Kb9+qAlDprYGNxfgrjzMUIymhkLfL2yO+ThOT9kHLb/QqRBO455kIGH1vLv/oGvqWEbgn
++VFqoy93bvZL2u27lIzN4A1ubbOx7VNnAhs6ZdT2NKOfG1vpVlEZbbgP9UMDfsBWbhe/kW6Nmcs
pVo6F6F2MNTEZ1HG+0l3OVCh+pbHns6hOene4sgA8lTL4/IMJCnmyKSpccdeB3q2YMqsBn4+0OW4
Fk+eJva7nX54BlNhmhL1Kh3W0tFstw+QiwvSvTDBFUf/o0k0e9Tyinh+PwbBxguOwvqBugNlNmUk
yBnS29kf2lGAtX8t47qFD77gtB2821dRVU4PmeF8mN3PeHiJLfWboSq7/U+J1erKIJ4aejkCYY09
282CveiIICk9EdBCHo+njtCMaTgjqZElnd9P7vIJK81BGXqYRsGm4RnivZ85ieuhfOVBUXS1snjG
qUKyPzW+6b6rIFXQh0MNu74IfQpRTeUdiHOZXvJ1AvLJ89rHJRz9cbnzw1SvDejEf20uGeoZMvWj
TJWd0U9d9nWOQW3Ga6F4pHkVUhikaArpu7j9HdtYJUbJWMieZvAr3lXrg791JBqcEEkV47H3WlEd
6riaoCC9zXNfGDvXkvQGeawXfJubiOwNfj76Ew4blGFjumR0i/7b6E6NRACaUPaTdTLnuDe+zsO2
WUM8GnIzd4eU3GCYsOYmO2rMHfmtcO6C6hYoC2kcZq5zrWJ+njDA33eItFK4vZS79jh/04ttX0NT
HyOwZsDl4EzZ6tLbXF2WGQ5CbWyHW6K1in5UbcDiTI8usSNQiRSOsAIAD3MeiMb5AoInOuHdgC4d
/LKvz8mRoG4b8MIZfNw/KwjXOmmx9nmkRrSvPkY1teilVd85oK5kAX90zTGj6ua16lLSGA6ADfm1
090C7eXG7Pysozorb5kzjBYxGXlSnyHlooQM2FAZVt14DBIjSbp95XgXizRa+j2HyEDP92TiP+rQ
mJ0USqfPsMUvE+nSInpFqZX9CoZgdu972w3SbuBnY5TPBrIUvl05XcXTfYvoEKwf2rQ1kisoH1ze
+d8zluG18BrufR6cAeAhAqwZvleLDFH0e8qLJ/Mwvn8tJORCHQe4iwA75BZAKIjVluX3pEDaG8wN
ABgtUSQ4BxOc6W+qoUUADuUXPKbmz9E6TtQ8hgKc+R/URvQdhUh6TXinCph6p41p4f+9xO4aM+G2
wGseivxcev9zgZDl+i1xtJcegeV37zjsJv+xOO85hGKgJDIKB2yIRJSOtnTH9k/fKaTtFXGCZRqX
cHukryzNZzKyPqpeVnhhA3DFoGARTAU5RITaYb1ZTZpKjNkN1r/XP/y/76R45UtcbBiPbA+ncwWy
9roEf3GLhwxJyYYv3YEEfK8sW4DGlr6DdE3LbsxDZHceB2M7B6OeBEDUQmGZz7LT2tlqJ9QuXh/T
OQ6+T4jZxAtJqzHWg9y53mt7ZO5r5tw4hTQf0MX3PMgUn0Upo67ty7pfcvUcppAf9xoJ5J6gs6Qo
9nFvYVWZfYjlbAooVwUFwGc4qGw009u8yrlFqFfqTInfEN1VxQ28IDWOs9qFdrl9HqrMatEq9iof
ECWMoHOGSYLO89HyDg70TG9g2UxBOXx4w0iBdzNLsP/kZMx5zRylGkCKDCmdiXjzcxtvuLO7l5mX
/AecN06JI38BjPeK/C2iBoYFD+ivIZD1CwS6xABKqSDG4PZzZef0953yYJwbPhi8i1u7YUau0X0J
QixBfBv8+c8SedZGg/K64wQTiqNVEvw8jdlFA7BYwl+TdBXTNQ+DEWAmuk45sHk/L4mfOpJ4L+uI
Ypad02kpAyZm/m/FErlIvemGQidKLztEBhMaiPqUYwoFDiV3+srcO1Oot4zEMPs4GITO7VGeVmay
ei633G9zfJ6QN5lZQETqjNM0YqzBgBPLYyCSyzf88M+Zaewgm62c+kzkoTO8hO43KKMP7fYS0idH
ck0jgFLzYbgbfaAmAzRPgeX9DY8CzKCzEzBTcivdchmTx2JaRwurY8JHbEX3BeHJNSHaX6dhf73g
LlMDBxX6MuD4TCnYyYMUCbCf+laFL4WaVsHJ73U3A8T1IH6t75TMjNdUitJPBhDNOmERbnohALHy
ijSaBb2GwiSVM5s3vJxaKWyEG4P04c8pCXWqvsobJ9IdiEKZQzguvgWiFX4eqZDQHxllqjZXbflZ
nGpflhMR37MAxyLBQ+ggNlTOgdqDJOJR88EnRANQg8pIin/V1IfA0FPanWlsED1Z2dDv686o6MW+
8Jfe3FcnGtgq01SolqgJMm1IcKWIT40OJZJ0foaFwtXgu/DHSAJX13nbYfoL34a2699nDGo+EW1L
QLDAWO/IMo/ZjtXHNTkWuWjBEuAU7U9Sh36hIaIwkS+CHhnVI0QvdD0PNKLm+W1tJdoXc9RsqC6V
VdGzl6nDhSu4g3llKYULtx4266uSJBOCgKcn8WyGCgcjn/S3H5StSPvdblflzIvbVsXs7C4IGNzY
Jj48mV1EJ8n6ObSTr131cTEajuKd//l+ram5vJcQu7X3UHuSPEe0Ojj9G6vtkDiPtzE6FL7q5gX9
5kJYuOaRZLrF6S35o26zJqvK0IUDjE7H4xdXuGP2l7WZiJOtKqtn68I7LOpVYhPl2ogYnPkUp9MN
rGPTLaas3TgAY+5Ta38vRygNfN8hCQ2LKWjLqUhX6Cetx0FGPeK/6f3tAsVDxnv9nw2lgf9GmMHV
FG99HoT0mZJdsppwhWrewEAywvT0AKncu4mIYr4OpBuNFw5uRu0Wqg2mAN5Nt3G/3Fe09JMVd82u
YwMXzU9lXOBnzepWcklXV+Qjq+BO+UHZInnG86zoe08deblB8ihMR7mFTqq0avc+CUXhSwXJ03Oj
TvKuKXHCBxnxa8NPMwn2n/6Zs4KJxIUmgdsuptc0Rs0ss3isi6kZS9EHBjYnkHclKn91fu2bK6d3
oJoQ5GhzRZf0+u+lh1ydFPUj6fGOLPaJ3L5cl80RvDEG0QdYTYguBT74B/WxHLT8/QMNzJGBz+4f
Q5BBdBmofPrG2Ok6tIP3p+JdHQP7rBB5+8BLE0Qg4bdbWauYFE/f2/9ly+uHT8mpA2BwX5xY0Obw
VZjP9YR/I2VdGyo7vPUalSUju4T8pAAnEmHSEKt7fyZdFTYBeD2uLxtz9Umq0S/4b1BkJYC0Ujyv
/1qQ9+D/KFbdmOBGH5U4LKYeMFjhrLe2Zq3SoT9shKOAb1JrViDKJm1lXtNoMLdnc0rh5PIXpi5g
yFu9TqQquRaFRSULGXB0SqfKxw8FFtwVuSdjPHPqqei84232BXaY+dwIRhClB1xdq6RZSzdtid6X
9UNcP0bqDw9sK6VHrdm5YbsCjNSBm7fJZ2YX/7bUfwtVKkFH9EM/Zc4v5QFJ7t7MX6R+L8ABQL3q
2VBHRJp3lpggiFBvO7g2ucEXhcVcLZz+mWEjTFp0sVKO3YbBK1W81t8ZCoYt63aqlyhgFqDlTZqd
eJYxhN9p5bKLb2wcuDbdgSz4hscXOLzlADCt073MRYtRat54bHinJuCTPl/u+uI9ZD+gYKRfHKz5
fYjNjqKQQ9dteaBufWMK8WHi8z3pLJbIknvKzchwGlAYxJvqpqw68rSmNlUp7Wp+u4Liba54FaZH
KKTTnnTWRTOsKfhAj+Z0xJvFUzxzrSz/uPLBwAGMjhWuywFKByyLGaJ1MKl4xGgqBnVge4/DcDYQ
A0v/9Tcq8hwQ4wcDa1ubpilJAtHXhShm/3qdDm/VO+Bq8DCCVrmuyrHVHb6F5toYjsOzX08n6QZi
IW7U3pD6e2TQ3RuYJIj1+JveGM2kobeUdHc3LZzFcRoE22X7raD9V55CZwmUnFCNqMsQxhJWFid+
3faomrK0yz6U/61rgzCTBEXNSRosGUaz5DYveJrSKPfQtmnPlJxdESsv7Hgszd2OSpQ1400mOFSp
aVM54l2bGlFwYKsTMG/7gkgi7/+c12CuUQQQ0THFjmW/HYliFijt08I45qT1r01VXmGr8UQQqR6F
IwvQjByt+5Xt43lOEqDwn+Hk7fcdSHidaWtup/AV10vQF2YTgZR//lXHmmAOcLz2ubBtc8U/n+B+
ZqsuQW0IzRWvVulNwoPhOcDUG4pUW6a2fZqLlRFLszDgrbyoRMO++nS05J2XLKTARzMJaMlL3bSh
pN8qLgby8MaSdgYHCZkvhxEHMxavswbDW6SnsrFPrFy5tXUVRKCcZcoE9Vmm6Ne7KSo9HevBJoMd
/Nu0nGg2j127fxcN2PBhWk3Pbhh+7NXC6xMhsTVvmvLCPvg+5mV1iS/hv0DZu/kRnx+eFppXSgdp
qvf8WYQFQGNevF5i7XrvAgD/u8ExFGIKIIy3mOf0AiUuyZdhByGdDbYjKRo/sdxH0Jzj3OOzMYzX
zm2TqXWAWb2gQ1BTigpEdjy35iUg0pnbDkw1zpgKH6vDo3l/10c4/U77KfOZychbc1VpWc3ShQJP
uw965xMEKg4bBwTlXPd75WsZcb+P/V1SGw9Op1V48Ms5TUoX4E+2iMRXlGFwV9MP2iKxx+Eyh0y/
yANYsDtvTTHqh+AujE+17RF85UsSycxAi8RoQyws8ie9nmVcTZwhYs46UJ5Y2PU3fNkq9PTuNVwZ
iDe06JWt1y/q1+ob6S47R2mEMLVA7GX6WZ13Aj7uHETH1e/Y9ff0t5lVM/WYwDihVRx7m6jw6xXQ
m6x5zT5FLW9od+9vTAb79uCXhKvF8/K3pnLwc/PqPzbTDZvDlbVzKty/Dfi5k0eP/D/5Oe44ClhE
k85F5NyaB9ImoiFt+2JybbeWx1LBNpJpCwRnd7m5e3jlLr3WoP3Kld4Nx+09XVjwggN2+I3cZ3RS
48IW2g2JtMEll+eUqIz86fnA7kMOc8ZiiG/QMgFXSEv0g5HXw4sjX0ZoOHjnT+F2i/mmMl5e7jC4
C6S8Lu1mlao4+q7y20OM0i3x4Ht67ySQUZ6fM8GrLeoBcW1mHG86Q7QSyfx3As6bzks01GJnbAef
nPEWC7b51DMUkmhzEdEpdoSBa9ZmLO+7gxQeiH75NGSvv4fRn6kYuP9yYQJ3k2PuEfS+nVjSCDi5
mHBNDK1zTr6qOCDJCFSX55kixoLCQLh4jDStWHFAq9V5nE9pr/HJ3UqONbm5gkQI55FQ+l2JMtt/
JnA6i1V9CF52ZZJcP+Vg7yphPqrB+VYMO6ghk+o73CNHD3OzuozmyWjkGsqjrJDdTXUhGOGp5GI9
169rQelYbm6ig6JaUe3d19+kyUNgQ6ws2F9FKlhKVAJx9bbrv7aYaEANz+GIDaQupa8+v7RR/ag5
UXmLemizAXreld+BW7KDYKDB3BIyoLZ7jdNriZaITPfmkyNeSo+g71vBZ8rnptSc00ymqJ15y0Os
fUWm2ku7A5bqlniqd6Q+0ng8Ku0hUF42sRUgZZx5a895DEDkmKopdnS75p4FxOhUaNOyVyVCLSbd
bSSxTPQfhMMtrHgtY7oVxUInrarm4BH2d6daHcXEBxgxwSMSVEHzb7eXjus7f/uUsdtGIkN2jipL
Gh3NEN973HuY2RHL5HbvdoL0/R2IVRXeKfLmoqVwaERfo+f0JUT7B8Bi73+pvRixwXzHJqHbPUfG
WSpg7QJKcpi8yEvWl6G34yy1DxMGIpyrOm9MqT2XY+F20KMmkHcP5QLWjcooHJdbiRCNFoskvAMn
Az+M1rWKZizge4Asqi27KDnubY58AGs33F7laekMQUPqqKL1L11ANz3uvCfaDyZpAahyofcmgcR4
/nGhFMfvIiM1PENdxxDfuM3NGgZnzMYXJcfw93SMrLhEJo2qX5ZYTF+fwbP2SqDRJCpnZnk/1VE8
mTFQtPSlYIFeaJDaeCPLB2O2g1/QrUu7l0MyCvfqaUvcubIkBKobIJXI5et5tJpmVUYbTQRuhh/y
3VAA4tEAEDkgrkLOu961iG80AyX2DXRVOaKtryZubPlUfP78xfvLZmlenbI2uJfQT2nj05yEp+RQ
1o3lt81w1UX5tKGptYsDxq8t2X6fvTPQBi8nteQj1IHQjAsAStLO8T/udhHyIY4houYw8V8kuB7j
RxXZ3c44+LZkKJ5g9zercdLFuvO/RlaK2Ln4Xj87Zhu7aV2q77iEtTQ6/4wtwPrUmYurs24zkIr3
gcGrM6vpbAZVBbclkItOG8e1TBUgcE+2sbStkfHQfBgAf4EaiTSJ9sacH+yQLPcFEcE9gD0syi6M
WzAcRCnDLzB8ONaqHZUlj78GSSbWWY+bk/aSVpG0ISTTSV8na0uJa1Mlb/JIECrrwDzXH71Bwyqp
BJ/BQ5GbTfiGH/2woD3Xk5CbplDwpShb2V0LvB49hxWCCaNLB+ULFAa3xPs3VQczdsTAsbyvUXd6
tCggJAKRPypLPeLXijwLZQQvd1bxi0AbWvyY1HUxC2DHFHrFXWIb+NsTKLpO6S14G+6mlnOcjRjK
jU9ojzBM+q5iSu+clCIq1xDym6FErxzv9KYJa2ss5PWokpSYxzckbPWPZlxdN65coEDKRnig22Hv
OFf7bIfKXiP3r9J/lGCgIqhwUcV723XN6e50vfnQXrdOkkRinF3IFYWzXqFFxszLDwM68417Qq9l
gzAOvQsSC9xD0lNo7Z52NLM7MENvYMlPpeCzo2N63jC6UWQdZ5mbzL2PqhmAeabuJxj0Lx6N8Ds+
wCga2Oj2RWRYVuKX1AuHCHLwYSCeNAUKsDY09CXJ0TY9wx0BceKmjQ9lgH+9YSjTq9YQCh7ApsnJ
HIbzi15KcYw+gHl+3vhowdKhGio+sXLK1EPzye40zHuwD5y0Tdo5FF2c64s9yN6BqzimB5AsWDJc
Db0wWWAptVilfj+uZYioJ/Oq27ynEIqZMo1UpE8bc4bd1eJYbIxxxOt16o7YJ2Yz2d8d+ide9QDL
fJ0mCrLYJigy4Tdra/C19UKXwNTQKP5l3MIGt0GMqCsm008aojCLUlsCQvPivQPZHNXJy22IZysN
k2YWnAk6vLglya/s4mGloRtFBggs+H4bIUzB0B+x1QzUVuuoXPgRdz0cDotQLEfyoV4FaRbK5s1L
TUn5bLywCUIVYaJjnt2MTxPqEcO8OLEV9pnnfAurJBQk+dgbhWNchIXeb+v6Qb4YZBFG3m1P6IHi
MHLXcGTsoTqw1A6xMk9Zv9OKEXz8rh8kJaxBdlNcWP7/cbetXGsOijA2pS9d2YNIZO7vx1Pqj1uj
DvKHam4Eusgl74WkjIirxl3Jq6wJISa4siChJsX1Cp/fnpwhMWsZOJAigtzyDlgubS4qWiESydD0
SLw2yjFIB9Clgb5frMdaqxpOZ4eBRoJpKM0XfCHPCmZ7qjb6SAHzEgmtkT31B9mn9nVpKWA6H2v4
78QF2NL7Nk0fITdTLBlucXPGp0pFfpl2mEslwNZgbVRWgQaJimPxtC9tGWMzsvRo+o+bIIm2f6le
MOxKYhmDjX81JGeExm7PLMmbX7IuzxmhD77vqQ2yZP/tJ0C+mnCmLJwr0Xk2yceSeQw1AGEYoujv
GEry0buLsmvn1EMZm9hhg2bk7HI9B14C/3SvxEC/ti29vuUnkXr9VJp70vK8YrXLKaI38QpPzNpE
zvkPWUzCowy1WARx99sQoFQXtYiWka2czFja8Olgi5hWdflMrQwQ+8A/xuBauQNy6xCfbiGmBsvL
Qg+llOmLviNLSq5QdhsKsm85rPjdjtO+a72+ybq2XzzC+aQEM8SFYRboaZ4l5Z0P9YrRpoaMOMZG
bB8my2Mnu2UDQScwbm9VQjB8J3TYEv1LUR1dg860TGnDDaPUD1wl3wuu20pu4GiXdBGNIVy96drj
mOkVHrK7fzz2TSVUUZOfP3SLVHbbYSKbXOxiqZzR6jtKLQwc3N818KIFi3T4QjD8zYXD0lwcX5BG
OmqAeDPoCDqo2M4Q2SEKDdWoTIDOTBFvBPoGPgpFXso2RlPgcWqJTY8w0lOTGjMw3OyDyCfzQ38Z
XbAXl2y+Cby38kOyVUkIKzh0ObvLb0T7DnkMel7HFytiSBc9Gr5nKzcEhKWCdicSyd+ICGKzq6Yu
CQgF6zaBBSzuF8z3UYGudj1c7ypiV41H/mcFj8YW/cYOEDGtbQW1emb1He3eayiGRtCOlmHhWeWN
2PeB6JnGorocpBOoWD8DrMPBxsRAlpNTI3sxAMr+E5dswlUGOvXiMHXPrBQg0cg8OMA+AJ+BFtfH
wZLUhEX1jPEw2JAxPZlx4/rqtp4govCztBCDmaXb6QU7r1RvHC4m2DcjNQkhX0GDAFv1CBrehcmk
ZKLu5lCol5A/yohRSLUjyk8Gfm0JCE39CfFQlUX5nKa8+Mp8F31DbQPL/bkFif8+yVRViSTDj3+b
vx8uqDJUz5dXSUYVYgmP+3OGFP1JWc/Zh9oiLeQ97D/iz+PHv64naLFX5VOWpPGmcSnda0xiobf7
wrducfdnX29djPC2F77Faph5t0Rd9phGZxFHzpsTLqborv3TcREmQxwmycN3lPRgrIVnhIr4Y50U
Tqwj3LFaur2OgQ17tBh/LsC27lSFxjxAx6Y85SRkaB3s6Mx4rmYzEUgJJcsjAQ4lodslL21hMOhv
oFNlphKJYrKsnAQpSN2kVZv04gWSS9KF+HL55p3Ggt/R+A3/78k0d4gM+YSQBFkZHAyw34vr8BHj
QaVg5/TECz/pkOZPfoKI6Muz1naqFiX3endv4hM9Y41l2RYDIQTf7sqZrX60IOlulajZjB80uUhv
QkFAXGyt3iVOwaUFfEiy8mrhwCB8i9G3ScvofTooV1IStPJ6CnRDJtwcTWc8+smxu/2n8giYYYKV
ieRy/omjheFVR1xD+s9Ipp6py9nH9/T05iDEFOvN3dpfUh+kvFr5WVPR+g+4EEtRavmV2ql6OynF
p2refAC/qLdimwy7kFkTDphfbGLj8B8WWOm3QOlBdxzUT7al2QEEU8Sug207BLCY7cxpeWx/rOLk
HI7nxDvXw1B/2tppQacEoWTufDwCe7M8ZD8mVuEeH3We7UBejFEL46T0/sJleUA04VJXX5emd/ZG
D5gmPhNHzdiO7gll/ccWjfr8PcYXBqYyf8pB1LDJ+AnOFxC2QvRgbZ6ieTs4k3jW0P+CDWgEbO4+
vu+D1ZIqj320i2A9UjCXNkO3twg4OS0LyBw9qs3edJNo9FvOT9aeTCQaTkhaLgFIafh39jt8VQ0b
WjsDyluSvp5Sinwo5s92JE8E4obLtHNuCBjFXw4wth9TRo5tKps6dzAsJwo6CWabgIsbZ3mPrE8s
5SnZ4qD73nzDCg4FdZn3LQNs0cbzugsmhh6tNFJ0PoUo5iQQpRO9h8lEuOdO1OAnGiUUiqeEQw/J
eKZARcmaibOqHEADqmfuL7BgJNNkApD/Znyn3Xr10cg8c6HkU9b29W0Iha/j0ApVaxbCZ588krZR
PfcQgrAj7Z/uSvS8RnkPAkbvgqTuMwl1UHG3Jx0rdWR+a9C+aQyQsCbdHcoBue/97nuRRqMKUQRy
Lcg/NcylhknauvvOe9NJRRXDsJ15xgdIi8/hW6O2ISCy/U5vvWeXLJ85MXbRpKA/L8U/4n0EvEXT
tr2GqbWJktjOiL0aolO1ViftBblWdcxNXg5qnw+wiwuNgG0Ka2TeMCQ3o7hWYuTl8rTuMZ7BJfWg
a9VTH1naSrgaXNbqi/XVo6CqbnOB0vCHN9inpUIITsj2XKZaCcFK+qQpLJH7OwO/+kF1P8HlDgh2
SAvH/ihhuX2DU/KvpSrEZzjl/PuXFssYbHxOcL6at46cF1Uu8hcsk2O+iRCtMOaj6cKxRNo0Ru/p
SG3h7A6hr3Ee2Ewdnq00zNKQnxN3qvglH7DsUz6OK7OlgGo1ENjACdUuXBpZh9UfeHNfDFde0Ja1
vvvuiHzwmGF4XNPg8/yJeAaZS0NGB0zdN0sypHkxbDw4Vqq6q5S48l4ezqHO0FMPl59TQmRJ19w1
GC+62w8+ng51qfsVDqvEdLbVxA9fLZoaqzx55MssgOa7uND7vpdNXsjc3J/N8xswa/NfzcviWoiW
O4h0XdWWHCJWobwHepyYMfgLPLP4hInXuTBy1tpvi4j64HjZQYeLPpmLjC3ZvnGw/1doIqS6uG7k
CI5KkoUF6PiUpnjhRmGuUrW+UvESESvXIXrGOrjDZm2PcfrdE+RNvCUA3NEN0x54DLOV42z56FTk
0Z1v5Nx5qYKjaX0GuXSIqyunzInujJx3kSk4jQQ7xt3YlNx0lpf5ZA0lFoGjjaPdcq5owGRE4P7v
2IZNNIBof1C7b0LnBVKapx04Wq4c7NuNFFdokr91xg6b62GBzRWNFnt3cSDM5lle6E2m3Y9sgj53
bKdDS4h24HG+H9d3jfJ2V4Yj/n7W/3w8Hd1QKWT7VHIE6GWFva2cYyvjxeklP0qRun8fla160Qqc
9lADQFp7/0ISah8gzo9L8IdOercgx/rbhyy52nX0Ev/nVvXqC0J6WB8i0oaw+dlRJgkMeWQE7Bv7
VbPxdw0M3tXcSlJxb+1oNKITp8vNPesO76YsFLjs9tDDiPQArXQHGqUCCWi9Y6G4lnfedTnYsZVU
tFoPtgYlJz2ntZajSJH5Ey7kz/u6aIowGSM60iKc8H9TksmPyyvwdDzmP/xlsInprx3KX6xfIueI
uSygAHgyuUeZvW4n113XzKWA72ZMHKVQAIVg26BPYc74ZpL9ztmVlNcln7jIFka7Jjz6hcRAGblD
+3ftUmK4HfABYDa/H2rRs9ODtWakRHcPU0xcEtH8wDFKmVnELRfw5NKrKpBMl5vSybpcRxcXzJw5
J5KTlVLAry1FZLqzNnkF073n/MxDrONdAJaMZeXoOp27KQo+vmiLO9KAuhzsdsH8F7aBUJMkeofZ
+BUw/3M8nMGxXa9bjkKwP/fp5dyTxADEdcYYx3Vy4n/VDxHhUDeWLaSCVdHwowvHqy7swRvK0P+G
Z+tI0tSOzDsA6KgkJoyP589QgOoKf4uCMvm7Sg+/7a4ZRLelp7OAP/r0XukVpYAyguRwHj80WNwn
0ckJxQwEKeI91GUOP/ArfBE1xjZysFAN7XC1zxQU1e1D2btvd1jQOhmZtj5PWPM/lZBPeMSFNuuR
JvGoaA70QKi0Cmg55gpkfBASXVo8NB4HqqO3sbE29GVz0oJzhvXiL3naU56yl/8F3OUDGuw6mUts
THg4XFaltydYMUkkVOJuBu5KHCwno1m4uUu6z0u1apJ2E/5QHue4vX7W+xVGxGFCp1/U0NmlNbmj
/p2CxC+tfo6aAB6sbfEByXR4AbA4++aoL5e5s9Vec+TRx5zZSXYG0+ZFRINXk328GKYag7BZCNdJ
q5XcP/rKATR6k6F7mpIvu2mjpz/KEFzFNfZRg3puPxY0GRPf0obGY70CBcg9u6lLElUW/Mf+SIrl
5/VxRqFB0DLqs9iCwrV2Ua8h38qjEFM39qCu85plBm4k15godWjYubwYZ5VskcU32q7KdZt71CJb
LPFbuyVNbmOwPnKC86x8vIuBe+Iny7F+eW7d3sTnmv/fXiy7yFyeJhvpjPAylusZpwQbtqPPjX4a
ll+1nPPKifCQU3BF86/mlxQoHtG0CRbzb1k7OQpDImuyI4GvFxXGe2UIlF1wKv84kNw28rvCm/1m
vxKz5ZHuywf3M9CeWH4K6+SSfHNvEUj023HDo0Ngit6BdlJER6PpGM7+c5awvZeMm04YzyPeSV5H
u6AFCU+Scy0GO6c/2ju6nYzNISkGjeYHDSBzYFBX1oKBSzMa3+r7t7G4wv9WQckquVm+hmEwMhS2
APcZ3SFyGRS4aJuzTTt4BWeeI5zJ4Rd3vc72K0TmTtJx77IsmBa2Ih/kzxOTy782NLbGlcI2dzBp
L6i9aq0TeqTBV3cDLbrcSTb/B5yQ9OPYOifEA58yfy/wOU5+Sb4MmzLgo5q5TfYgA8HEZVjCCvyV
0xztdpfRFH6Lml3yJ7ZF+5nicGNa7XkdAEQpY30hmTFIjOdOGWV4CobM3Bz+U0570dGUXaC29s7z
8UqYAuC0Jcrv1DUgdEcuNbPzyT1exgxqMG+LNr8koGf6fBKkGqx8jFEmVlfVV73JVxb3M1GLid2v
Fr8WplBB+pL73bexeK+y5cRqJ46wF/c/O0lbquJ45X11aSC+uN2992xIKpz5lASNBrSwSai9euz5
F2uy8ybq0QuofP2vUSZlFXa46IcMsZnCGKLL5BISfx1PFVphEJwcsYWVSAMKkBRO+pZZid64hJ4p
VWusj13xglNSkTWZ/MyNVOLeq8z15uBsCJNI1VXpEpZevKKAItYVi5LjNbrcj1csEP+gSlvChmDA
ZURg/JOKdeSaH/e5YWdFPnmvbmc7YwqhakxRIlA1wa/0Kvez34cjveKT/pYPTKS8rIDLiYvpLla3
9eFtheZql6krj008ISs7mGz+FOu7Fk3dinx170iSVkupMJAbLw8gfwFN4tPAbkSNAgITxfDSx5gD
B5shlETxpEbI8Caw3VPpfdtpSfsRrd0srh6VaGWiQEkCxzUYUNdrI9bTrDJRj/uodeU4JnITuIy5
7O5XOjmU2U3+PJLuUT9/4kDNUGMJ6kHcVwkgwgXQdtQvBcJjA9Gc60c0VKyIYru8JCnzM3tohzeO
38rTCwlfY5qvUg9KEPHVhwGWUMVj8QlMjMJD2OIxhecIeh/QjR271drs4yrWjcKUJ+CaGwriLj/R
5373rayvHJJLtgesFNW2jhOQIGcOEocH8IWoPlwvb3YTy8JiLgv+w2zGYQ1IwvSA35LyUbmhMpVY
MMze3hJzVDm5mY4H+lizn+wXZxv1sPYKo0Ew1GDsfC+eyiuByiBuXuJTLaCTDnxJRLwWLNs7bGdd
I5V5Hv81Bn4kZRvdQl2+adBHkEcdoVZaQew3eN3twVonoFQT74G3du8Y9frgZW7P+TBd909DENiE
lxDFg2UmKtD3MqJD4uwTwzD1lEur8gzy3EWZHUg8nNb4IJSNlt5Hqbzj5qOxk6flwdK8/MmzyMCu
Qusym+Hfmh1H/aR9cmO514UvUsx6zvbVx5vPQMulHrmwphhjVsLGD1EV+9d/A/cuKR6vl8u9i6D7
NWBvfftLq+j/z1ndBxNFDN+c0aRTQ7HKukNRu9NMx9ULh+kAPI2V/vd5xG032xEcEoQtO4azygvI
8q6nEl1NfAkvwWAi4IaKtMUbupFe18lfoAb92PKApGjWuCg4OBaWGjV0UMIOHPe4bTKfKvhWORq/
vSTkWbhT3jNotsHwCxWVjohnC/uqDJFg4KMfNbhAuytC/s4ylR7A4uclp49hupJJwgBhEMiOOoUo
pHMxA5Q6h2tDt5l2iqMo721TCmAAU4P6IQwiiMcA3wz/hOGZVkoWTHFveYN7C142Zi2sMRcI++gW
DJWmdT+waRRfe0eoCVEtQUAhoUy99bQVop4mmxzH2jbiXraR2qrr1udPpvUnmsNtKdiBi06liP59
t+opSpmhcUkCXttaIHLdjOAVnV02mg79Oi3eBn5FPg9aJekrFUemYZzaQ3qDW0Iw3ZH1YX1WLpPh
b83ORDWQG8nSrq3ajZrWKRnR/kQIj5f3X1uvGT3qKsn/mRwphD6tMFY+BeY1LspTIc5m9/vLMfcn
hp9hxQLzllySEoR+xAZhLR2kr2LrBU4GkxXb1r4BaaC98BJOtdckYtZYAeybOCqAduJtSttIMToK
wRvuZLqDeHjNqGU09EuhfcfDyt/yes+zpJ8RlP+IdxdJLGS7lArqN4M2h+HSftnpPbsI8wBXTkwo
fb0leq7O4GP1xyRX9m5ZLzsekDSRCXzhMX5+tJABs5wEUNfvQ/ijNfUy/hwLHIN+CjZjweZjTNCL
LUcJtBc1iXdzhDFLk/0wc/qTkFEqhOlVWMZEXJWdFEdoJyKWGWG6XvYuuWxYjRZCG5Kei1j3RusJ
+VhJ8srg3vNhsUcumFsrioWBOv3/i69JdmQ2+QSUs64P3L5a/hGF/w8zEv4eU1bM0TYkzvrFn3mG
cBr/EzDEjxuDDAafl40vVt3KRYts0/crIr6Z0p9Y7aguGHagr8/Bn3Te1DyUUZu/loJEPk2lqXzC
qd86fZCyS2buGF8sRIDwHBjDXqNXFruW8zIwXt1n98IfxF6gyYeDBaZaEtDmg1gUwTBN7reYK0wn
M/k5Rww3ni2Uzd5So6fzHrP0I0nI27xhrnzZwlhCHOkUPuinnmXUAFPxJfLtih510ULMUBuwxcjR
miyCRmvsDUXUqQvaXwg5ZnrZErf9Q5pa2cw1ZfgDxM/Xoy0vL0FaiL6m3aw+MPPFI+tKbdAMRVPi
tk0JSw5N+NI8U3Y6JCSuSU+qeNaetNcN6a+C/f3hMFPodqJ7t8tytdb7LwlBzIqwAJhWlev1U50t
6oj0Ff2/9DVFBNiimXFgERGxPDWBa0x7knmphouoFrB1umcwTA4zw+ml+eKFwqczfUtEiuuO83O/
Cm0W/pCg/R91x70wIxiePzbG9Rq1d9dy8sGZ2ujRnHa0ExTHJbAldp3fwC1zphuLytMepFkFJvuT
oyVxPdl5v76WI7BIYTzw1ueDEcZHd8DMgUKZNmBc6M4WQQpkeWYD8nsVooTnEdp1eJyKotsl7WMm
silaj3/T7t7JQsDUrkx3HNne3b+azMssf36Wb/wPe7yknHkDYyzyQ8RPIw1oKhmEnm5Tgex71UU5
tDwgJiAcoxqbAmLs/Pdqbxjbsx9sPckoptDnnuDrCrBwsJEbO53Wg8lP6ouoJ26ZPoxH30DIGxI9
09zPEA6zXOF2rSGAwt8sitaEL9xliEVwjwGgs/Hv+FOsv2P1Nu5NL2zMISeDKOiXGYHiEUIfgi5G
Wx7oPzMWDh1dp/K+GGODt6xs6dHHBqpg7bbf3C7BM60i4P7oOekZ7NWtn9J6L+cLj2w5N3jEmIqM
bRTX55wvAkhkSqKqwZS9qUY/jhnIgnCHVvxMndJ6vovpQWa8fLoUOKY9ocRNyRujd+lxGYMs3OOC
+jdZGk0OfG5Ycp+LfkbF6uf6edGWU+/TgB4AaS6g0249pmJE4wpqsJZgaGpvhNJdF0p2cTonB9Wo
XlylqrNPIS2rd+dhJG/J5Q7Z5XhhRTDfdqU5E7AGugHrinbezK9Wd2mFPb65THn+B5dIhV2DPlgh
Vhvktnz5Vb6vfMCelTh18X0zMVVlgjP0138rjUeLk6DOyy71hVLOPSGxfcTJ82WkFae8pPB/TiKu
YbOihUoJa0wReFab4QLlyW0PUyKBMV0hVYFb6UFiq+kkd51ucNiYRe5sdx55DDlS9e6NKwNeYy9X
ei5McncldPvQKBgVAelqPgFQ6qC6NhNcjJvvH9kCtoHVarr1jOtdG5ryWw8UEx+MFRB76bfG05uB
FeSrYQMFtBiLZn2rJjZxQocY9YNROGnvyrxj7KQVljTEMhPLmFCbB/UPxgupsDdQlEFYqfdkJ93H
7xio/hRF1tMt6RIvafPECF/NVeqHrjHAMARUp26jaeE/033sAzq8bfTXEF1zgWWmuD3/aqVbftov
VTEw+EkOq1UvFSVpJbkjPyVMXGqU/lNQ0VKZ+kHl4gWt6uk4YWqCPdAZSzEeBNhbJocaYUmiEPpd
UtenBQyFyFppvAQv5/5q0MyXJEGMLvKds9KXpNu7qmKYohj0irDDWjqeaYqqh3AcMYueBgYFTNS4
5jfl9En/Mi6RswjAEB8oa6TKxx1unouHOhfX/mYPRJw6JZ7nS2l3CpDsD9Xj+AxwbDVW49EiFWsr
oSR8tuJxvkp8fplC/5blMwjY6effDFwKoT8Dj2tu3seaTuMFC4Qkkz0Alq6Bm6obxbw6Hxi1BV42
Qt2ulVt2KCAq3YJdBc1Ur+Z0uqTOgWtXQQnBnjL12g+QgHmZjMbn5gf0rqfd4JBAg0xsY6jtppZ5
VGZopwaP7dGZi7K2xhkiKxAfGTT0vUK4vwAP8C3XycQM9u1EsI+1EBxolBzUhDLGKPv6Zvy+Hu6T
Me/b/XqiR+bLEf4P1YIG52PxdhRJC5F0LxDnbfY6+hpPNgFRoPHqFfh8NKphIW03EIaDshGHyjtR
bwvm4Ku6B0wWSOx7XyokL04kJqangeNUuP0zwxU4aEFNCFc2ishB2XERLwUmPCZ+/Pe6Ij1R4iSO
5mbIbXDcOfYoyLzAKI+PWiiAybC9AsgUTEWIFO/QvvAS2J95r5L4qhBwQCMbasM9GvfQhI3VvS8y
u1ut0EG3muSzIeJ+bC/fYHGsF97ihfZ0h7yWmn9pF3S8QkkfG/Jx16eHd94HLGplXl2h8v9qdTgJ
c8eNvR5RNMaLo6svCDo8tcqRpYaSzg62Z/JWz1xKg36TvtC9qsePNDokJpbnf3bA8WYRJX8ZQNf3
J3Mo6sDwe/DoCXldUIws/OtRmPpC0p/LfZvDKU7Bxq2uIRTIeQspgOeYR5V8UmxdAHk7Sw8mesl6
Ep4eTBB5V2sxtGbcIs7DvgfBUK+Oa2b8r73Xftbk24LAe7vadVY7uO9Z3FmnZGBXYFeFjM7qn9xp
S5JlPymfJ3IwX3cEsnM0W+ZMZLqLx96I7lPamKaNdQhwkLiMzzTOmP2a2U2QoI2kD9hHIr1rUsBr
Qt3tD7mWgzBt6JUtn5izXsZ+nQPSyUn5ymhQ9x14HfeuNrRBDbb76K4EGCKZP9TM5UNq8OgKI8fF
8f9CRxrYz2vb1IILCAWCjQlaJIR05+nmLk0ChJSyYUGBpGiPv/X2CBcSvDTeInLIBbcgBMEY2w4I
dNj03+bT3gsiE8Yh7U0sEZGXr/skytO5i+su+aIRnvGmTZW9CaEGJnYo2ymGBCZM4d2buw46iVoH
2ZoeHNky48SICSZfh6psNJCuyQ8vVYR9eaodWNhsi51eE8D7pTYxeZbv1ouWYIIFElHgwVK7aThi
tdrWznup7ZB5bZA/J1GKfnIIvCZpciKqnGR/PcysOnPffeG0uPxFYUfh82MBHX+btCK0UkeaFUvb
Et9ZRrBRx48ETU0QrKrLXLutzSF3dJQeWa9KmsjdgRYrI8NbmxUkobTSoXhjajLson0L59jtJzMd
x+sBWNEsNK1pUy9+A6K6aPq8QnHKxLAKrPK1wpleotVxhFKGazj0mWrdXafh14G7vUvXDFVDQBHd
qJUPqrubVY6zAt+uX677ve49J/lB71KzLOexmUNjRl1BeDEglQjzv+5vBFJVNTLUYtWvUUNyCqca
e9o+d95wl2byGo2dutzKNVGURu5Cf6HUWAzIPQIXsDBh55VBcHbYjEXvyRPam9waJlVv1eezttZv
D9CHWU9jkRMsMbLPeN3ppvymYVJQ9vsuckaS9BYZY0VAmNNX913FhiJ4ijASZJ6EMNPq1tOVUl0l
NrlxoaLyBV5L4/V+IFkHl0R0kO+uKhSyoKrkujXP3TES1WEqI/3CxpeXDWKHS7lstos3Oy7tnivW
XkLqn2HeIeeFIpnWyNk4HJV/SeLMyRqb4k+McrAgdEvnV3YKBDvHYe8R1qrXl7z1Voyx9Gc1DVIn
WHDgxU0yiNntd3p9oWDuus9u77zxw+lYyrgg9URtKcQ1g44l2S+quaIczIx/oaR6pyfF1QBM5/9r
hheBO/ifxO2dxVmFlNweGWQyrei1ZjH096W/g6jGAacxaQJGeRgNnSz52CLIxDLJOweylrwrgfba
br94FkCB7ylvULPObRi04d6RkRGZz0Jk037WoPHGWEm0WpGVtYE5BU8HVakRUb1CHbNcECWUJMfv
9V+jAXz7Td6BJfe0UOqQtgWMcAxwK/gjNt6o1aE4IwvQuzgsBzBagUnmFxIpBtjzpkcpzDcuunte
VJPgj40KPgEaAlxhqbXsG9NJUQ/f4pVuiEvqIH3sRSkQTC/pDDQftn7M0JPijUMBKGFP2G2B32wR
jKvUfZnLWWjjk9cqJsbop1ATAnnkmB81AY/eHKuZ0+y/erzeKiMSl1v5e+f3VmDbZeTxcNKocZbm
3mQYLPe+lTw+HZQnaNah2wnLQJDiweZQGdqaDj34DFTgSc5n6PWFqPL7Ps2IUE6xIT3g4vXL4Gu3
EGA5+PIhqE8GhWqJwPoTds4OPakmH8mHWvtgg3TUDdSS2VI7+iLJgqpa1T83h7F78zLPh+9GISF/
CKh/kJkEon//xlMWoMbcM9YO65AP4qNvG3mtQDPCfQFvtfPtD4lJpdaD+bWArIOj8v+02Tyuw8cQ
TFoCa+pDO8XCV/2buXxZU9YNYpeyhKEYRHpgzW+N68oy99BChug7Rx0ddmXvj6uRH7q5cO7fIyiR
oMbhSnTt9teoXIxKUqpLwymnTos9s4lex4VXaS+wVRKQPwhCNHVTpfhV/POKi9yDcX/e4srxUUnZ
z3Uv396qLp8MBmlt0QwoYY21GgXHv0pzBR0e9X2FLswpmSmThsJj1TeOxurG9iFWj7geBBKEOg0l
eIZAbVN3lnREZ1htc0I0YDgpJK3i7DZt8dgAyWUZGAAnUS/+7pKDYfcrxrwyMR+goiqTIeD7stR2
eSy7jClxwa/MlNsn51R2S/8E1SoP/9I0QdT6HRIgfZOcgDjx1Cl+2cTogkHBh2VbFReJ3MmT7KZ0
oH1ifrixDR4BZMOxak46HWITvnsztl4ajuCfJXqDMnJwsTqOXctWKLHzgltiwbmFPvZwqm+syKGg
2/0rvbNLCxDRVGxiGU7Qynw2JZaoBiovsooWzio1P9OdX7HQ8PkHYd4grXchcWGgPietQbrchzkh
E1kz3TmgmcU/eJ7p5uMwVb5QzKXWRWv2xBOchDUkYV6BcbTRSvNY8AEDNamgN5E9QnMspTh6zVrg
lPPMy2SJ4nDrFWDMctjgJ4NtVV7nEzc5aIJc7dnzfju/x1FOBvcN3iAqvJN8LIKT4BgK1LHi3bOj
3/lh43a3ccuM0G71B1lFpXEq7CjU/vGgUVhFIMGVw/wMlT3LB/iJSjKhO+/Y4dcAKj0/hyILCAoH
nzGPoC3B0QNK6n4/7ylDFKjcU7f4m7ih0+3o5y9ZI/z9zSlqj4qpfFXYvTibmZXfqg6MGDVBInbQ
JWwRj8WJLpVbSRy/ERXhIKuHpTR/3eo6Ez3sSqQwaog4aL28qWx9UaXY9Zynnm5loRSD+cXYuU0g
8CoA/wH1pNC9CZJf2+9oC/OD66rQ/UBnvhPI8PxeAoQV3a4dfyukcpUvZ+1Xwm6wojWele3sNcS+
AL8FCk9UDC4Y7AYUzMIYKPtIY3URQ/FwRGy9UBbl58UTgGxELUrx+mdq3SzXl0LZx/maiTq17eii
blFZguk2nwiMqyZcOfvZLM1wBO8YXERVPXh4T/dP2vJpszk1IgF+vdh0ZqIzz9N9m9Flm4K0zdkC
FbVvfFNH/gpoy6QDgVYzfD4MsQV2VHSymV+Rm+TRrc32byr75ONCcQKaS+OGXJsuQsyfLAVqL+J+
Aqq42Mp5TG4mLOA5v7QpmslvsI7FwScyUEmkIHg5vfhLp3D6t778fEO1JAs9OPaBPiCRdAbejtwk
ywqdwplC7CPwQMh07PfzNBVUE+vQFExclJ8E1Q8ifP0n325Ba/Doq/Rw58B0O40jSYI6kCB9bZwa
nMcSSPG+fvloTzmmQNERrFt7XfFvTkHI+eVNSCug/ydG3IjmXy34tQU8MPlfgqFpPiOwQSTMcZLB
ot2b3xFLEHmmOroLv0H4ZGkaOxUBeRo1b1RVNn1muQ9R/3zAEQVEigv9gv6ISnxdodrMNYYrPBa6
pdvscflpXtO8w15czXCu28eXug528QNmvzL4wKI9roHSmWPSDCJNN50WYY92lVmYsp8KbsxF0dkO
aukxHJrtk5VQaUcIQtW61w88oMh4yWsuo48SPeY4XrIjk0WzAbENVACsUW4pdK7bXfQdr8T70UWz
RbRiUYkVRn01ujXD21fVr9PZsNmEvNKUd9R4Fml5Wfhf30+TYd7cbLe3ULusPPPhDZz5rgSqpDIY
ax36RifsNE0ua+iYkj6Y6O+xzjZjWwwxcz1JhhfISa8LhJuVTlJ1SoR3qYcwvES2qFaqPwxUOuI5
8AQsREXq1vo82MViaP5pmBFb/40scSSjahqXZzCfLxdqKs+Ox8FXaGmbU2Y6zwDiMmt+5EAfXqiK
Gjs4m7lLfHtAbUzN/wv0lD6SEp8aCc9w8xonkx5BZB71/iAVgB3nNLboyUf8c3pX032bQXdnUhKK
G+jImJpNx91eWH0PW+rIgpzRQJeSWdiYVRIfxrBxBT8Ygux16ViKzWCqp6BErEmCnjb7hp2IKfxK
JVZEKIt/Nc5kuJbatDr0PsaimsntZTw2vZADoYGh8kiom69Kmtrw7N+NXJWoDqoM2pCnFoFnx8xW
enot0We/X3rBqVGQDZ7iXZ8qjUVt0SU2e+2OllOLaDeeVhtJCbpXJhq7DVEaAyuXkG22yzMQkJd1
+SR1ABg/SC1g9z6uCRfjxLMytKh0bUyYq6gnn0uGSCy/YxLgtDgWzMUhqUDogNqHGd405Vjy2Mtp
jt3hmcHPiBgEIxEN8fXVZSGF+V/cYx9hR4UeGpm/j0nlMkGMCPFPVa0AzHW5ZitxgMU3Hjz8lFkb
MQyE+NY3ddPCpDAFl+T8PmmYcon/IsLBLXzxbhm5Uga2Wvnm+TJx75wyCbQeusEnvHGbf8IqBUiY
2JCRALKnPcFyULY2OuJhRmNJ64adodO55C2UUiF+ucmrpsrlXLT9vKiiwrQE1zk/ia1xVRCka2H3
Vr8WAlbgHVsYlOYtLDjk7UwUMMhiYAUL8UXLCZltD2IOpt/zbdW653yl10PBTH3UMpYwRxhPEYPE
orvdCwSmopJMS+D2vgtGL4+uLa66EeHm6xUPd6+Ctdz/IyiRzuKb0Reo0H2vSL3VOSyJw2V/vBOh
mY+VVdbQjAnt6JN4sVAaSqj1+6H9w02JJ+5+YmPmJnoGHKAG7gujxvrz7xXj79ysmaBWlMNC34OD
p9VujGd+Fkv2jTDTdJSZ4PBqMC4gCh5tkHP4lUnVVTNInW36wdOpJQD2bK6UcHGA5Bw+xEXbAnd5
uKesWbAJUM2ReaPmi6sZGqbc+SiksE7XgFK1f6zr6KJ7JSYBbAqoq908kSuEMXXY/SAQ2S1tZReV
XAihAt9RMrHTZNxjdAgB+xSP8+WMt6C4iXY8XRkXXqnC9ZJUvHJ8Vve4N6qFlQVtAMXA6VoF4Ner
vSgWlN7FQznGu+9ZEfvbrq6JzT2luhlRHa6Njl6/Fw/vj218UU8BwLPJalGOd5+iHTd5OTUondwc
t44oaq+HmuwqnYSCq6fbGtPVDZAwstA14ISffIwKamtV0zp8AFDtvla3oK+XGF+b2EGqB4gead9u
jX6HuuuUwWWq2uWqH5+V5xBLnd/N2X5kc7uGvYgY/SsrP5LQW5nETZbiJYLiai3ZTQ1jmY6kXuLO
QKvSXpTHq10nvTDoQVa/Dg4xb4kdTO7KMZI9VL1s53M6tykEtXBswelMcjO6oyyYCD9GDgyco50o
UUL6XlA3ty6ipvdbqlsRKsmvaGdpFFdqRQ2YSscQHu1ALDdzWyFvlxag4NZjWWZ4pynda3tZ+L1f
S2tRdaMmsrn/RSARQO3oEj89d4IUBc6Y/hDQIwQJB7xIeOQ+cIT0YelOhup09LpY7DzsA4XKR+Qw
rSSCco4gOk1EyBjD9foV6CqLYhh6uT4QsmkSyEL4TR62TotVa9lupzKhnrfWs8OmtWLWyfrvqwUc
DT6vbC+oMAFckQ1S85RjER9aWPX3d3V6kBPCsLcYYMGa12KefMs6fHFAoEXMCpeHPOSsR8f1PEzP
oPq4oSorwmZ7SeuU4kxWRiviiFfKnAtji16pHGEZmKPCLlNJohPLJ5RSZP0yHXn5bnPWbEywuHPN
2q1qRHa5jw23AiQOi60QdK/N3J55m+pAEEx9Gh8sGiryxjCIRXG9kela5KszwSQ8Q9VSjAG64P6V
6o8ANBp4qJmD1yGbqVBKci8T0jwLNqdrlEyxxpD9F0o6v/oLHp0GrHHN2Pfima0+1exmtPJBCBcO
q4YbIYKQ9dmy5x9ysNbCCuFhGVt6HJfCrSraE7pho4Z1FZQfZMDaiLtA+dRrrZoax9woX1fHyjXw
i8rJuEyBCQiY/J+AiwTqkvXQBJPDI7z4FsQ8FKTTFokEyMZ7vbsWJR2Ho/lKwSDiXL5g2oqa5lK4
z9hkJU2SYBtHKL9KqzVhSrCOus4ZDRrXCBmQdH27A2qj0OQFwGjeJr5y2oH7UlSzynN/d2NzxNH0
XlEn7EbpzX3NmuG7VmmFQBcySVJGf0XW9bvbOxGim7S/3DVcpnEMbGGO3nprqe2MFKDjWZ10g1iz
NjbXWsXbAlpS1oXy4IjQyC9SJ92xk9zI2YzNv/Oee9K1VVFlCT3JprJGIwjQWLCTwnXVgazdW6Jk
vDvRA5O5Nch998EN+qfLjkN6KXvqiKOVFH8QIZHYzbTvxi044aiDJ5H3hx3TxhNysyXoqnT1lCPw
PGwgJNVU2aurNPGVFGxF05QGWOytpZazE1tHz9ljlubwJYE7D4uvKE3E9ZpoZZyxGx06aXadNmOv
LEcobfBpbtVPCuo3iAIRY/O1s+2IeCwevoXwyGbPuIkVk829FRmuauNYSVg/B4m117kjQDEJxOwk
PL5Cm4bogiOOClel/abxgCV/r1PohK8w3uFCOqpo3zOZHko9142FzaMrLn4ewOLkwvRI9/DPJDX+
KnapRELDSrKIL+gk3DZzHSNOaG+6IUPqMrDxAmj4ICinstm9iqafE/4LGDqZo5WJT2Pz01e5mgH/
rA0Bk8Ykxi1U/H2SoV5MWiG88O1wMLkBcQXeUAoq5UwUTIdIMGH6rR2Dug49bz8HNCaAoaBD/wXJ
MKpAVgm/XIZmOSSr1hClJPwhlmGiTJ+9wkW3SpxBQUlWakHcBVvxoJANsjJEINVU42DqtjSb6XkT
HRw4QUl7VyHxtWX+u2PMSiA0ogB+UBT7+XgsFE+OhewyUozu0cqmvm9CxoU9gOw8hMWrHXuD/hdG
E5ZJr1k4QorhTRxfGUqhri1t0XGw/EOPLIXdr45QOwE01T1i1Doo5V+srgggUwYeJJKEjz2NpY2a
VqnzMARldgIJjeVejOJZHkN0K60t2w+w04F2inAhznJns6oR7up5GS+lyYenV/r4GMmvwUT4kYsV
fSjCKxwkKEz8KCiOo57JPVtDtTG1MVcdsTzL+ZCmYyhy7JfLzmuRxHhiPzw/idxI1XppM7X6pZnN
4XrutsmQAIBCTjHA3CGJ55KqONKinAbikDQpSkjfoM7JVgixyT+ehZEnLSpwk1IJ6KDUd0liYATF
JlF3IWrC//Iy50aUpFd8d93jPoTHi5Zf4sw8IKVys5yY3VlmxWt2u4143zohrvGr4pk6MiRJsD47
wM1nQQBWwvi9d7rRPXtrWdoRaX/eI3yD8QmVyHmYHOaEaON9j1/EubpJBE2GCuBqEfoiujWxZtxH
ogC/pm15GzYSNFEqOeYW6+yYIoCligqEUvKh4fJTZlx136rF8Te16DqidoUiIbc4+098qKFxZSSp
YvjVLN5vz6u4UcuMX6Pl/FaDohU+sJwr1AP5gWTv9wBPC8Q9WmoK1LN/TXyY8LfacA6yU4dgmAV+
g5M8ovW5Yw43hys3XhLgiVCHJcgjneDc26H+t+Smwk0UQgXuwjgfNBtgqn5nWInr4Nh8cyFX01eH
RAhgMP05Bq15pMSDLYWkOHm+RYPbUZy+CFbHFd+y1O6RCBu+wZCmTmDYOWJXKc7qLY9+61y2Lyql
YpMNM4Oxp3+SE/pu855seZnRS/FsZDXqRTGFoTP5p8lko6Qb5Q2wBDmqvnpDh/pa9XvP+r0S5pdL
/3G/RPGY+93ZLizdwYXFoMMI8gkelt6DeMIB5M0Ky16SfxIMJGTSF9kPwr/CNNuStRMLNBkwn3Eu
EKzG8WIMD7WLeaUYI8K9xBpWw94eyt4eMApYVAAvyHc2zTE9ernSrn6G04OoEHLgkdA7iKV7y6ON
7JOZ2nRg2jxAzAtbDB0xsONvIb0Covo1/yV26aHaM+Qu/pkuTorGLVk7bm1F1mzLwu1wwONjSb+K
kkWIIYwCKg/r97BUe7ioV+f7jd0wUENXmAJhU/bLsASUoxM4H5sBPIbASgVISSdpkc8Jew0dSTiD
1B60r1LoZnpwwFcCjCf6/qj15Zj9l2GA9M+15lmMyZp9robWAVhExnf8DIkSlo6I33DBpijDcB1K
rDhbpqTBFF9H4yT68LAECAlPjFgCQTjMnztKSY+dvWAIDt90OvXsKE/xAOJHT2SOq9J6qJAFF63N
xHrxicXd1aCMHI73jejU1tcXWmdSgmWnKn53aHvVOMd/fcAmp6YqDp74zizqEDF1KR/z/DTITHb1
fLd83hBKBRdm7c2vPR7i18PnVkgvbQxijEjp7W6M4YePyuhhOaQLmqHI44Wons2fapCqZpISB1wR
GpLv9SAlE65jwsydgDxYNSO6nNdhMC70RYXUg1xtYsdio1T8k/jcxHLxw7oScebs2nrZCyqBE801
yB1iwwjvVbkUO+oEI20RhuaDG6+Y7K7lOEzNioXVvLxH5KCvOd80WDD/jP1nED3qfmluerl8AuWF
Xmxs9WRKvGg+5J5cr2+e1Kv4A9suKxKK/XfQikvWU0oB9pIPn+JaFtWzCSoPz2ne9HYsOthPJJ+L
FhMY6r5dPPDkb02wc9nr4an04xSfNHEUe5zbBGLbAa9P0EGcBisScBG+Spq0S4o9Dww64NmBA+bP
zCy0zklM1ONy2V8N9ZefO5AvrbQ9YNRlje3kk5vr7/vbZHWXpmR/6WggoSsUMHUkIWhEs07y3ZBU
Hi9jpL+4rQTJ5l/rsLJOHW0wfiCD7QrkKR0xZXN7ltDr6Bh40P6nM+T1dajmddJGzxa7jSm4ht4v
xzXYl6o7GS3T+EnzGtrOQgb0lUPJxT18ZQHumQHu7Qlhk4cH+XNx7pGcem8j4EXHVT2ZeZIqhggy
FqOhUMXI5uAsTLUt271Reqgr8hA9JDOmumQtZQ8Vf2TBmnkmy5IgH+4FITzyHU7K1dUVJ6upooM6
mCGwz4jnjdpJsM7c2E9YixO4U0Apzx85BlWaaEmBn+b5XNMlweA9/pkQrXcRCcvGNxRRjXucAYDB
mG39Fwpk5Hujx/P4e9uhykf5VsmTzyavEyw4ybvoLLZ6q7Ht5nDf/onnp2ETWiaQikquRpjVKY4t
hMDful5EiznSFa4in7hQm//8A1KqfufBYRXlSxPYCi4G0tEyvoewy5CyfjgAkzB5PW3smoNyQXVq
cVwdLDxHiOwXOOoVqHFFMWbvmykPIpo1QN1n2S2I0bD1MyQLmrhUhW8/IP6R0b72wv1xTX7IiOej
uQs1YGWgAL4HIl6oBGx0GvtzK+7WrnD1oUh7yrq3S3z6hHMhf0+CUPuKDOkc/ywOwQMIlW804M9V
JcL5ZZchQuUrLtZmNNVxhngCB7V4i8ASOxQ5Z095OIOsDC4fdK9pdpdoXV8h/f0FzMHQnUFr8DiZ
73Srex3DeOJFeMMqs4ZWEjSU1s/RkRzTielzqoHxEJPQ9zYMTWWQBgGCLE3JC0XLHPCg3DGydmuB
m6DlUHpGeHDx7BBV2n2IJztvo3dIOIw+GIPVITjpKyfTxLWJViq1+0kHXKq4+3wiD7EK2ksxK8L8
hPoyHBMBR+ysxkhaJeJ1OP1AKuNAp6UoOkByqIpBbrJm1KA2db2z2wKFZqWxo3Gixx8jAFUYqO89
ZrFYf57Ly2rE4b9kxyGe76CU3cZiya9C11/LKwoi+6RjiCeRhBt2aBKCi/9w7+4p8TTcKIa50AtN
dVE5rqZTqn7L5UASgvM4TQlcAcUvEGOoqG8brwMd8xhv0kUqBcj7mFUaAVOOEMdvzOmx59/LrmWB
6HL1JqNanGEwN9wpexcv8WgwrYy/OAjzftq8YU9n2LBzwJnVTCaRl63U3dYkfEyLYz+vyHaEvtTu
8cySkB84u4OaDj4HQepDOIJGOwW+cHeUekp90/IrHYLQQNBt3ZA6IJb4xUrPmCL3V4+Bg+jsQPMn
/gVFbYjFzC3BMi1hk7bEyQvUG4h75iHv0OC+je/9DGWaxKsH1cXEFREjDgqSFudHthtsMcBD/uhm
Q/nq92T5WS5/f2gB3ZdiIvf/XmsCmU9uxTXNA+71ool8heStVQDPr4QjgUPf4DdhPXwj+VxKihn0
aNZRhPEzAeYMekfC0nuM8DJEJKulwgBkZnNR7CcS3u+q83OVrBQutFgmiD6IOs01POPyhuThvvvI
3V4+4AeM8pGBemaMVoPNWuRTTa1q8fn/gwknZvN00LhLx2Ehz9jb+8AqxsB2EwoYvjavVfxp2OR4
YSj77Ef7nM/JVZaYmTFaP944pFd7BbBewrt8M+KI7mpwbs0YzvPsLjImJ8k5CwXEseRiBTkuM7Bi
Y9JD0uRjP1rcWrvpPxY+tdAAuL3kAibc8RKf5e0e7N3Jkqlsm1C/nPcEIWMVm7kV9IMvfKoIrUGz
+t3NUu9ZRQciAFndhOfbO0oMEGXrDp5aMf2ZdykG1bgLL7501YcYMPaJM6v+xnEk3FtgS3n0qGiC
slNQr4hnI+L35C5O/+P80td2uwJM/J8Iqs9p5KsYYBe2ab8PS8cEGJrGpDY+igKA++4U/LElLcXY
e1jZqFHCFCuddTL0Sjx+KmR8iAYqIFayiMytbEdfRcglw5Aliyr70XEvnaNqKv6CN7ApWHCK8mhb
bfihuC51L7crDr04bncOPKZzhOrz04a5gk/FtoeV1Zjcuy6z9Ka+HHQdUfsVmMv4ih/GzIst81EB
Ug1PLrfKUD23rYdw4bViu7NEgqXIWlVvMWIKGbMTwjl0U+sVx4XjYHU8UvJSZNIRwF2gbE/Iz8FN
AT+naBSZVLXZemWuMdTifji6QV/F6UIbQoJVrNM/xCtWMrcbp1aDzDm5FBdAoZRhbdVZYgOV2VRF
dboZz1qU2YZXfl+2xu4l37ojwWKpGqamdtw7jEJ/9z9yhnbAsz6litcqeuTDL6pWwFzPT76M2+kd
znK3SQ/C91nzPbj3/gymmRc7hGcmIC3Ier9zSoCJYYSc8zsTeuHivJ/R3RlYZiW+zsWcHTmPHZ2L
cUQ4Wxs6/J5HQpUsrTDY42X34ykHMM1DueT4BreBwUEnR1dIdDQ83QGZXPGtAU7IAOgJ761KvrhK
u5yWgxssV23n88F4qDsbK0JAlixgDI+AugQ6cVlMC6I4Rp+ZsktoW0+PvxPOWX1T0JL6h20oMufE
gD7wRYBZIM7wCjGcg5h/lVq8iQvzOXUzymfwzmFyBApWMo71DoPQYaEJkVHc6feKEY3WXdqbWXXk
Cu5/eg1KEB0rKlUzTZHmJlrxtDRdzcfx+GcdUB6G5oGLTmYr+RNfO2TygGUZY8CsHkweKljkiRq/
qT7sC0oY8+McT0nfnmuXNnFAWsJxCOXsAQID8vvYyc6bdhx3SwKPXrS9Vx9xcPMpwzzp5gXgc7E/
YpPbrEvlZKFRUUGQeWJ8tdjYJS/m3CnKkIKnsyOZxZ/FLde0t6YKidIBnCbm4QPhyedQ0ocRj2dZ
lK7yHsIdCNPMg53gcYaWA9h6ewGgKahMpJf33SqgdSw5m2xS7kLnikPFLcY7/fIhGwN4bwqeZISF
9T2p8NenIn0GA0oIQHjZWdT8E99Wxw5jwsqtvtihRTLW6f/KyZ8uibx2PSYgqcOLBxOufDmyiDZT
I7cZnqRnhOC+zv7UxZSrAw/N6bgjyRk/8ugmKWoRsVtmXRaso6ohsjjYJdBNnM01o2QL+F0VljJE
cpvtTZ0wPxtQPs4JuibdgVPCpf9ekN2ueh5Snlobhi6jhZzPGxd5qHz/f4wfPy7LK13ACX+gE+8N
NgHuxavqkCyn49jQ8kdidcURJO1Tcw+XvZirRH2TTnun7CdxsMu0NF2omAMONYnCQOkCBza3MRdx
TJ5WK2RkhrtHmMXqDcwRZHUdYdaJxbcQepp2R78jNpQBVKHC6VWmmTb55VdMR3wxMb09hQWbA6XF
2/XlwuqhKvAQ1LQBE9zab/cZgyZDC7jVRfA/x/JWe42vHuCaNXOE30XgAOy2UF8kEqNRnz6vkD3E
etbbxfruwIlGZ17xSwHlszpQicHVgBCrnViHoY3x2jVHFpxqusZd1GRPKxGUFlP6FEmNS+p3w9KD
zAlzwkG0EARtckcOZtVu2gzcgu7o7iqYj79Mwt+tWi2Rla4+wWuJkC54G/E7fkf6kynvala01kYl
porVMne42vu7BFJeg7buhNyZnDIpwrcQKuo5xfhXRUVBlEuxfsdi9OZ3Q0CtwoxJKnVaJTXeAQIP
XBJxcC7oMbXkZIqZD00pPOOcvyRFQEAdegLmhlVLap3bo3G987iakJtMxhFrKOuM05LyrRpEieXA
lNkZyF7alE2IIg54JDL9VsuvzRgvBuqfSUtMoTeh+talweUPaBYgjDVm4SHUyAy6Uf8ak8FpH9N4
lBGmWwEK0R57T2wW4XAKOWgdcgO7XmOLei6ih7qt3bMjl8sFTAL511GtNWFjjOLBBTgp1/n3p8D9
/Zxi6n0ceJkbj4fmGZhxt+HMxXxt33Kb8MqRc4OYwuja6uYScQ9xzjajrpskkA+JQK1d1eVAqTYP
REzj4WDKGYE6lhOQ6XWuEYYP8pnUkk/AjXdipgJWfC+YQccJkJW8UYKuN2PkRpkyOk6frigIghFj
l6IYe/aOgVh+3XYa9VTYeW3eYNZfX48TiL+d4CDL+3ydI65wwZS2yQVMtqqR0wQF2jEj5GP6zkI7
fw9ElmB1Vw2WVS3euLvQPPseNzAT+JiSCaYZQpA8dcl85Cr+WtmDXlbO2Wvv7D+/FCXdkKLS4+tj
TNWrZVbjvvpskDHC0fNK4eXppoFLELHu9oXdNpSgHJifdiKds1jpSCzixJDHwIHaGSjSlSv5xV+K
HiWqLJVZ+6a7/nH6P5SoBaHpWcSYq9RFgVD2DqO4QOd+wDjV8Qj13j0kgypmDytBsJ9MlHfvcm+4
8KEDgYZhY6/1/4gEYlWjXx/kSP6D9buJBZ4r4D5CQz6OMFF3KQRyO8DQ6I0huXeE0vyqdXDJr3PU
35Hf/GfE/l33+9QtHWIsHzbeEai2zcwZMzei0zekFSi7lk2yVjchQBlJ7yiw6sL3NYjgUPH9+P9I
Q1RXJpYvEgfgOxN7fLymwpfxzXSL1ZW91/vgFV+7sJnVSKPgMToWNtP9bYNnGwC+fN+7GP00+rXi
0Zata2yxnkowmX8ihCZz9lV6xU8j7HEedaAiyjvWMZ6MMDtwYhOCaj8WQVQRiIPPPuI3yW6UUE+C
6YDW//7M8EdP4TwQlmmwX18BzsF1yEnS+iWmM4gf2ITHH+DgN5HLrm/x2EbRZhnEHgFj/8WKJJPl
jwo3QKLVNhNvuTH5m4OVKye48W5OWk/OgRPY/069CgPWrjfX5anfqyJFlncLsnhXfccRg+4Uc20e
GMqUC0Jz1zRLor4Q8t6BRE1m9UCi1zrxDaU8g3vQ+yA5y0AEuDgJTeFcmG6tZwYli5zq5vMjFWs1
8c3Q+gJQ2YmLHJH49jFXTOVUnB0lCrTuwltxI5E4Edj42SojoenlYoPMlmSUWFdwUcswiHHIk1Lf
XHDjvSF/HBDFotNUUAM8r2qvw1PTziGHnewIXyZff+MC3+pESTYiV+qvNBkeDe0igs15/JAsgQQ8
E0Dj/mejrvKgnIligbUQ5y/lWfrgrO5W5Epcb+R2Qh+w3SE8Gg0ERKAXjqkL6i0rgDq/ESEAvAgq
XzzySWxGXLGVcFgo52+dJSpSwg6KW85DdRI/7RXs3OmnqE0JHEQ6ewcCG0mGLEtUJLcmyG7E6fjv
2uRjHHh25Rvvx80DyOXIFOSQzA02+VhO1lAfgXXvpo8l5hdwEPkntfOU7HQyz6f1o+xUTv0nZydu
5CQPl9etCxw6KuQJHkOIHUOyoIHztYJ7i76PyC4Ip+cOk1olWJTVL0rDDlBTwRfnyfzdb4V7f8qs
OH6we5UcOpPlyWw+JQy8W1CS5Bh2IP9q+ohHrKnphdUtM5o/S+KgnLY2J9Qj77o+95qpQq5ANIM3
iLmqzITvSOAfhQKUFMNAABWNRoVFdVfXt+u2JM+ty594RihIoDF+kSurlkB+YmbQmSrpq8XSGLAi
vInZ1PCiePnUb33IKtrMskNXzu29HGEtsSq3vH5X7cyNGYSdVfGb1Eu77d8MfLM+6hxbJc0bNbAR
KfFKtSjfLljNkw3cLIgNBRGp8lRFUYCBx/NsHoQaY3AS4R5uzfNiWlEjNNKBq3v+uuUojMVpWpLK
S8cpHnGkGtOhYIzn0GEQvKDEqnKpmZcKaW3S8w403YQJKsd+f1i8ZttWy/x/VwWz4F47oVle0OAP
7Mun/rPZoxq90rG1yTASDZM/G/+OL+PgJIpOQ4JQagogL8jvmntzyCPILSB0ThnzbGWsdoKDBKr3
6080vHntdaObllRhE8gS3c4N21wZ2v3w+G7zQwTXLHhxZnMnUYc3BLGG4jgTZPj5HTiLxTwjMPzj
0BiCtxTtAoXuGwxNLxmRv76d/EDeRO6Rsy0ezi07wQQ6EL0sbEug5q8lgNmADEoZjcjJFVgqGiJm
l43srSx+1U7+ItKREZ1J2WJ3XBmVVuYtI3dMi3Dsr+33Ap88iW8Sjc+Bgvtd4yGaHUu0+YIHPapE
Vqm8j3QBW/wG/vCEd32Bbr7LANu50GEzaqcPhN3MjFROQU6YGS6D7MadkgUxUpsraRfZcOrqvq9m
tZDbNGLJ3tNK2BNrgSo2lP+VbnsAmVCPJlotzW3fJIpMj15mZz3Y8qO8cLlDNk9V3OKkcrcx3r+4
p41T9qP1plFu26blEcJkctmqetYX2XefEMsVhGQzur9cwM4EcuskH5vk/qNNI+Du/6mt5O2aBtBX
Xjcm3W4hHUZCLx9F1buEvZ4ncP84xzXk201Fss1tJ43fxKF+mU+zUFBx0UqltV/I2NximndMF9lP
0KjcuWgPvM7waEqosiueUmghaRsQyMyD9j+NEa7pc4mseX13fI1v0+3+GWUKRPC9sl0ZUR8rWD6I
K/kMKtI/OZU6gA9IWg2Cworr7mzy0oPX/Y+4g+0ReZItYWZOhm6RCHk4aF+TGOePDxbZgZZa4RIo
xTjWpB1r8Mx6LpEaf9LBBQK4WVL3OrqApwImhmwu5TukRqjNtfYqBcSdz2sN76PwokNXAo8D7/K6
uWzIr2kqvFaI5W8WPWUUEJWmLlYcUwI6EHJ74qxhxXcESHbYJtGp9J/ePJhBx1dOuXeI08+JS9WQ
EwWaYCuoyRpdW1TTjTrmrMfKJ/hLbQv/O6Ovu9dfKDFdM9Tj5z3m5WIEpOoav1u7t6Px7YJEwn+O
R2uXc1jNumssLEQsXKsgrJ9b5KQQd8be8G5px9iQ0w8d/SgwkOeFlCeVJpIJpIIlmCQ7foEQG4KK
2JE4KxErS/PyQMGBUVYvxkIM4+qhqhKue3JQyYdRzIjONyzQtHjl0k/UbZRfDXcgUMrxxX51/bSz
SM05phgA1t3z9sVlhc/z8yOC/Xw9+UDjRYIgUInGtDza7dgzvOUdzzAgqkMylGPa4tIg6Ykyfr3W
4O9hD6Ikf2DBWK6P4Qsgz2E8qa3xCJUZbWAG570mYVYhx/UJht48c0abCqCqn9xcTraJpGPlF0t4
RiSMUw2V5rB3vXOJPEK0fTUyljbK/cKV/tjPyIKXLFIUnLdYwEip9u11n2fJMQnApQaKQBvttNrp
bJxQL/m0D9X4gRgIZywM4tvgA0GKPMg5jTH9yOPtUxGVNjNr0r6zCy5s/E9fmd0Ej60z8qzwlfR+
s7bA+rqXD0pHKxK20svsS1Q5ZZmMPBRGdbX53mdU1ApUkB6fzoJN5wJsvRMBB1xC/dBOLZA/RGz9
zrDQ2YlvxPpRq92bGKBk82cu7ntTPqbB7125sXrviv4lzwPXJJKEi2dAGZKToA7kWI1MsOu2MVdq
Gte+eRiNTNq/jdWe1C3kmSsh96S//y5xH44nFzzAx8sg2EtJVVc9qBrDW1ubfYEbtZYUhc71bmp4
a1m6d3R5fQxBPZK3zbe6yWgXZ2iwWQwGClcAYvqn1GFFjE2aAYGG7opQeET7LpFXgbhT1tWFPxYJ
i4kHLZ0ULugUuQOrJt7DlRgY5j9GQdB7uUrUgbSU3cuGtv5sT0noRsrOlq9E9pkH5gKxd4bUuK9Q
xxseY5nnX330xMdIq1RD15UqivkaNEzXYxuvmKSlKGliW3/0K++HKRLnP7suE+6EOwCZhEeq9BFh
aGR5p81S3d9dAjyntMTMptjqtrPkR9aWzrx+w5/vdEwPsYF+fxSfPAY+yDfSn4ZiDceKe7aCDi5d
1e4t8lA4ecBenx4sChRbduU3PFwqeJBtK9rJwq4cmv1VMhlkLJXcO4U0Tz/ZrxjjKqztFssCNEIS
Nn1uC1gnTX2g+tlZLxfHGg3APvHCgspODqpt4sbhf5JO9P2DGfSGy66x+W6NFHcHBC34/yVJ3Z3g
pyonroTszlkzJZVpwtq5o8CXg/YGFjEpRRLItETMZU77U0ypb7lD0w6jfbGKnJrhRcvg8SPF6enu
58yUbX5rgBLO8wZc8+JS/aHtpfDj4RhoWjeUtPuVcT0SP3QJ5IUb1xm0aU6uIS4pRbZhklvoJVnh
Z5W66G/o+VF1rWd8AyRGDnG/bDskAV/77teUoUYAfwvm8SZ43x8SYuYXEi5cVK/Oan6+m08TYKn4
6Ss/l5k4UUkfv9GC53PzgUGzaG07aV4QgyXke9hrQpBshf+Zzh7Z3VODzXBAmSbF/9ZnGC3neBl3
V/1aXOrzSYRb2VB65FvEvWX4+gy13k+LoGxZPlpCIKbiIVws8w4w3U22UkrSLissAK5mbzsTzmKi
hkbou683GMxJIzokfXt9QrnlP8I6/dcHo9QNdDm+Sjq314RDwKt7o2/7oVNnAK/ZUelfBQ/FjkL+
VLZ8jXOSsWWnT/iaJW/3k9Iid0DTrukPDTqOt5lZLdzimD8ypk7OvEQMpfuleYqZClxJV8F5A+1d
5WFBnqengm0yzX+u/O6DpyMugMU1dgzuIuu8A5mKzGKkZhAhd2tL3IZR0MHYQSaYsOg6ydOUM+65
fJ77iUlVRdo+SEH1lRUhVY8/njd8QrXH/1CGTT8I/0MGnrQoVIbLWbbPb9hbPi+H4DZJv/K059at
dtGf7AuANPv2EQCkGugTghw2XJfJLGJ02NjhxDPQ3XjMn1ThGjaiblYl15nQWr9VBuoAVy9uENsb
m1AMYYDc+tNz5Vcp1diBs1KzvgoZS9EVHisr/qu+tF+0pchm5cfuRvUOUy4w9hpH8nL/ij+j6XCZ
JvS9UEPJmZgz8gbOCJRfqAaGqvIMWrMddo2cjsxrcZNZ4L1BhcZWcnSAp1AL6NPKJWHHSHtsVhRp
HzE6+ZASRHYGnaDf9hUhE/1GRMX28FVPnHW4zPjvVy6fQnncW8J8MBz7SlsH1j2vgnfOOegDlqEj
mqPzyap9NvV+pp+HV9wBi82M5kmXyY0q0usEmdwqqQlWWiEqpkTE2A5xMYnw3pBQqdG/WglfNQ09
zqSQl2YrypdT8eUmQoqOg4aQ+n3+CrJGcbV6wZud//arr1TA2U9nYc0bVg+cS7t3Dy1B/dgF7GUD
DstsD7zfbQQJVq5eMRoe+5qcVhymBbJEZ0el6XHYvxE72ubY6JiONxJQEzlYfE/6XvpZvnO+ZNgV
ioslWVyd2gaSEbYRtQIEeRMCHRErPF+OvbRejP43SOIIIe3y+Cfh4RKwdorkd80hYk2MWEMEfRhn
qGoh3lp2XrbioleRUiGPXxiIQVTN7KOZPnrBNHoUI5wAV6ux0BTNXUe7rCaIeZYIpENNTIZUQSkc
vVhGm0nvYV0majfLw/J15cpSrREh2S1E08vGVR+fCQChAMh7ZBZZ+K6sJt7d0P/tIf0HBIec+3kX
ni82fl1smdBNWW68DYl7Ni0HWg+GCgMAMzQ4r8IvLBiKtuV83EwEjNmfwrfkdw9Kzonv4vjmpGbh
9Yyv5UbHzf8qvruLqVAxu5+isKRBgM5bTc5sc1mPxuvQN7s1jZF0sX1VB7Ba1RJigDBhWSH6DDRu
Sbjudzt3kfTDBua5/hECr++7UTRpmhOBqASXjL9mcrCxzNMaN51zrh5qPDS48q4KV70kjgkGwCEn
i5/emyWV7Ri0O+8nCC+QrbECnthgVVzrfX57RAihiScpw/8B6axUkYWvlwmqSwK2a/bxUccAyKK4
QYPr9iZ2ZLY1+7DC2MReJuc4z/a1BWyme5ROcalmhcMIA6uHOorx/JeRtIzqNYp6UYRFDfuHK5b0
u8jz6rM+JkOOavIiy6/hz8ZuXavua+B0IZ/MHseR8BwzeCm/bcq5g3ghWMnQd6SK+d3rB6tJfyMk
2iXU1W03PlSQhjVrFojBMCWie8v2+E3Lt/UYqXdSNHwophxBJdc/FQGQgHZ/UEJlle9Zf4jQ+xCH
xuDLiOEV1gSN/9AraiW6RETs8cSUewUXhtm46o1n56ObYfpVOiiR+BLmF3oL+ia2C9YUJPQVgn8L
rsF68Xby6hXuQy/XPmjD/HmAwG/BVp29GF37pccilOVDOW8b5JZfLpaIFe+VrlR+wPYvy+a+7Hb5
NU17GBKXmlgnvbpTaXbfYkq6/hvMAGiXDUV8pdwJ89tZ4KbO4YfpN+Q4Oa/KPHAfffEMbJR/fMo6
MIlgAwPyIXcqNc2vIJDeMonYUkTy7u1mxZHp/bg5tnxEaV8LDfSLRXHZVvPby08Z1DYRQwKUoFyE
oGMlwrGR4xqBsu7nCQ2JZ8q3561deTLv1cSAXAOUX8CZMnhVKKq7hminkxAYEchFR0X5sjyPm2Uy
TyYOWDmOyCuUtC/bOE0iGjzNKY03fBGiEHd0yRucs1uoSJTVqkSBoXqjZ7xG7FquQesc6uaLEoAU
2ndqrZj3gRFI2/neEImd8if9aUm34+Yetfw+R0xq+69eSibhLFTcz0iy88evBVM2ToxylO0N1Ifu
FsRFBVk5XBb/BC6S6ioNpzY+q9CbL6r8njVkOnjrlmkz4HfVcHAPGdjCXZajbWxB8oB4Zso2TdMo
Fzw+jrjgHnyXTsP81jo2L0ROYg5A1eBL7R3eeFHyD887FcXjcboGL/gG1kGyJlrfC9QuOGQwOt29
wfhn723gWB64hjAll+Yyonv3Q/Hf9PHRj+q9hLj2goVCtIUtvoVYZrTU150pRxuaSfR4H9X6AC1Q
M7HlXWfsSNnblBe84ELPAX452fFVniKOyjwSDFECCfQxAEZUQxDSn7IUC+DuLbC6pENEjmwcakFf
w406EU7Sn2VcHBvKk28eqLeimP5+fqmCAtqRcdWOSFyRTZVmyhuOEb894jJgMHISHNM8/71comB1
jnX5V+nISLIj99VYkZb3yQ0rKD6EpFgkUTJ2T6muqvQAg+mXcJXgRTwa1U7v69NGHPpytEKtl6oh
JeCtgIB3WStOPp9AMC2xxYVFYZzRui6K8Nqg4SIGRDaKNjD7DIz855YdYZSI2h6fQo8BOrpw1bAF
l/c2jmA1JhwtqRTxccuvKlLI0TMGUPtrNZVYKhI03Iood+OwP2BELWzkbITck2SsoI2t53/DqlB1
ObjE/6ls/GMDleI01WlTX8VQifCCwQEz3Gj/zo5SGky54b2wcNHOk/uxtQjiFJhZOVKcadAtLvfi
8hVcFoRTZNtlj2D2awIW/xMsyMCVLcqMKWFEqumWAYldq6JQm5NZadH8JOBxNR0LfPN5Ojp17fUo
XuCys7P8FUhgHghPPVjGaDaYcNPBFIYe2pcmP4Xp+RzlyTZ8adchmFeNZPlb0lisTzqVKrCQiiBp
Omzm+LnwT343fEhgF45E9athf/FO7qgbywBOdrrQjO2wAOLpzONIDD9dZleQOxKrNKFCgUh3d7la
cSG4GjLzY0X4O4huZNZ8V1zFe0+nI3bPqlL2hzuOzAdlzjcoHUwf+SL0TJYedXtv6C7em4yn8eY0
IsoDHas1H2RD8uVkPWCrMzLdb0V2WixsMmBCIXnbASfi50K87STp3hZyc6sn3W/E3KdNpaPBGzj+
k0PBk9jK/DahA8KintqGej/EPipD72TSGcyejyftl6DZf3KEJHb4WTEeqe2KKVrA7WlcuCtdV58W
gJfJntL0uYyg+nce41XnDKKQ0+CJrPEuCiJ/Ov6tYuKlCc7tSc6GmSz1eZemHujdCGh7L9SkAOtt
Rqiest0KaYp1oFuXqIQVYqnAa58WbR5yvNTqdjCcDZmBxggrs8KCNxCUiwxP9ZGPOc70yWDnrP7H
BmflRRcIu6h9xuQMvvEjHEnBzbnFsvl9++83NOfPglk1YJVoJzfTvo79pvepcI0jzx3fdjHJXlEF
aBjlE0M3fcUFCvRmC9JQTXqUaRsYG2Koa9ZpURUmnTCL2nN89rZft1l69sMEaVoQ6b1/FQfayTEr
sf6fsPbrkFaMqVHRTzJOulWYA0v62MyRXd7YjLIRu8dmG7yzl474ryt+gmCQXAx/mTi/MtWO4zA+
w4WPiXrF4q+te24RBi6z1TAhaJIZcd0dDpodCjB/b8A38QJlwSL61gMT0B9DrSSb4fsLwlISWc0M
Kzfp7GkzCi8KF6OavZNVc0Wxv74fLe9mWTgP7taql8xsKyUajgyf/IgpCBLEQrDilu6zkN/8L1QR
DopkXgbtTeprSOgKtfR6SvfVFuf3GcFlYuMl2fZXUytgE67iLhYJ/hvOVuM6WdnQ8WUUZpxSAZzI
E3LYeWailVOJV/m2Zx6JEU0GydkPl7eZMivEn6TcX0Q9PSUzOR6c//pu2Cg7A0/eMyVI0EgxYOrP
LlEOP7YDH2NdmaiNuFoZPg9S3k6GmWBu/2olGQoK7MHm78US/rAJdEjApRWlcw1vbRPknETKHUws
j8DMHERDTPwPMzJgrEs4Vln3AOdxs283475jAKkwE3ad5N+OHd/vUGuRRYwgr/cZ3ktnuZWmTbzL
WASev6mFFWheD4+F6hCNM54ttjzj04cXPsU75xUMkjdLOKIiSsRtw+KDflPTEqh1+6J4V0o1T41I
o95mLtKvGSXX0qXOS+4xjPlZwWMnccCK4GFWGandzbyDGN3KAau3bUEWTVf+0kBJd+Lff6IVr3w+
L370DYtbNQquMInr7LsIM37Ql4yPP0nGLUjCOabeLuZLfY3OWKvDt49FJvS4TacnE0MvY6gSrnFd
GiFkfBDWY4A9XBXIQFisju35Mc3DPOdVEarqNi9K6opwHZ12R1y2TxRPyj03d/MOjVaSqjo97gzE
RsdOi5XJYvAmisPEwBOAoiXzg8tYJzzLku9fLh3IcX5STCa6HuLEubAbFTfzZLwgHAKZriM//TpJ
64yMeSBIOyhowkyt44RzzrapNTfNnXVOIv2cveMv63lLcZr49K82paAKnG27GZvUt3SIiVCiCNtv
14WuGTyb/K0mPZAlOuWMJWdrDRhMMvI+xWaGiZErNzIg/EHPze2rbfM4yShAtOwMYibVOETr8o+B
TSr49kzaIBS+wiahvOlph1LCFwbZneKw97olPRO7RNKVit9JZVzCPd6SZM94Fcf+4ON/gMeuCdqf
kG5lg5GQiSZMAlRxNOUQh5r+1mpcdXV6lS3G2Wl1SkDOsUFZ16felxwYuT50WHlh1T9Q3esQdMaD
WiBNmog/gDtpzSj5BVwrNqvX5p06CfFSu5pTKAWUSrg3mcTiX8SORawN5qjIJyKByGFRlLllAfud
XdZssuJpX3IXXPvHi+ynm8I8OX5bd3oswsMIHcUW10e0H1txdRxhmdY9SIo98vk290unzZoRI5IN
/Rm03E5blKIiie6uheL2hfDQg8aOjn96wue36xodtJQhKromxqhV2WDV0ORyDk1H8Ob8UfErULYw
uNsUB+jaP918grLunJFvXph8DKRDhJrDDkhyHs7RJB6mGwzE/NgeoPvXlUfBlgyfotxAaxcvKlsI
gONOSwUFyTaFiAqlyrvy35aYIBDZpFOoOV3ztlX0XafeQmJFzHYjryeZaB/EUoQu913SKnzzy48w
R5Wi4AviP/M9GqX3+1njlmnKRgFBiEI7JF/23dFV+WcaRS20N4gYfdayiRdq+xfsLNRFqepKLqv8
HPIYp4UZeNPAfakvqHX5gjP7k6s4pWDyGTEG6l434jPNvdHzT3EG4D6wC7I1nP2WspiitDcWM6vh
uyle+0qvlr6iEhN1IX1EWr7NDRht8w8zM36wKKO77MiWp5n1yVWM0IEnnLavZogE++u9v1fiDaUb
50Bxxn7qolPaHuo9y9w9a6/ZB2aZpKqXmnf/HxrBqeKnGbK1AZbCgxZCX4ZzQqdDbYnmL1T/B6fd
kULs9x2Lo3ci6vXCGmblJaowY9An/YNu8lOFQaUd2a9FnLAuaoQqbZ9ntIggGcFQJJRF38EMx7TR
r6fZYaVnniiJyYhyY72svgj5PejW9XXOK0RyOtfRk8OJjxuwEeK9gDDGqJXeWJhnZ1dY+HvvAKtz
5dMcbfra+hnxySqr2Ms/rmdV+26IycnmSWM1WZumwlC91ZYcP4egwfJnBSsyV1rwJNsy+GWS20rv
Fx2u9U98oP2MTuT2tzaAD8RvmLSsiAzObNzTfqPEbnfQ7paXQW8eyWjbTlI614HNd1JJiovJs50t
VRKwcJgmvNFFc5vgfmEU1WYNKFl4TdRTQqjaKW91dlwdSxlBdwlTSb0sX/72lVZ4sOPJEhOqfrMQ
IXV47bGidKd5w+ok1sDOK7vq9A29oYOJmDOPfiHXBMTuD26D7tYSy7QaUPhW3MeKMgETrBn3exN8
C/TmQ9l+yPMLDcbV/M3JvaAwBE/sb2YsLHfQ7Pd7i2fQenk62KgHpzY2qiqZqtb1LezxqEMDZBzB
6p/9RkvlYdw57e5G0B97/q7ve3zWlK79k3iG6Bn0QVoV8Atnb7JSYMS+Sg97DAGusf4BHhK7yWWo
AHMBt/0gU7aV4uwoQEnnwUXPsKdN9xx0Ye1L2uhY9l3zC/+vFypGFaes2GaSm0T5mSfmty7h7Gw3
+0y3WVMJ7XPR/TW2I3s+K05vWWc/Wr2nWYBljTXyGgmxF9shxC+h7U/Dxa1cLHnndjv+gk9ZYTAq
9qlwKLHdQoZn3Y0u7JQ+GTy440YkEtPWn+IXx4HWQZXukNOtsrmqvmqAC9HMVuoKewo54SHZG8/y
bsHSc6uXCY0ZbTJN+3a//xbIDFrkm5NJpgYKfbbyj7Pl3RiOik9hhFZvpi2HVapf29RMZIXPbxW1
pv0Wj1suA8dpAUQTJkHicJeM/vWIWp/8xXNdtmWTENGGanR5YpAqQEaZbLnRULqmep/u65RYq6mT
CIwsz1ftteXsBlR+Bk9F5Vyz37x7Dh7pV1d89G0xEyvaLepbAZLWjQOztbQzJozkQFxDBjAtXTxW
q1ta3pOo1sFnEZA23nm02i9cchA3xfd4MBRlpCTnxOMU/N81g6IVGJQb0UwOEBjg6rlgzgpJxeQJ
lL2wbotLLiK/sfwLZx1GqV1CNi7VJitBmsFPQ6JGl1bEoDCca3EcEZPqLkL126dVl3qyDksAfHsi
sCSPwedvsV7eZuImBn4Mum/O2EmrNI8Fa6qg5Ou9d8FOuJ6bW4/xuy92qcc62Xeo2KHE8tJaHht1
Cl8fGU7kkY4pfihh0/HCdlF2grOvF7qkkoS6NpgtZfPpe8Sq8oCeJ6RpqVvHMxdogun9qU/4yS5k
v0n3MZ3qF0y+DbGmY1il0Le2+/z0sk9uf+b6KBBYTBqvCM+ZsxGBCD36HRczOnRZge351CGhOaP0
OJxp3+43hbMrdVzc2Y1kUYAndw2Q+Ao6pEdzGJhUpW7lXX2OeCLd79EZ2sFdrcrIiqDVDWQ3jEPu
sKwJAQ3ADPut6WKiT95kMh2rfsW6Y5V1hQ0mHqwDW3L5cYA8M4QjTKn+iSMUdDaC2iuQXKSx3GtJ
H323x4W/pddZpRZoww5SDYVv3aW146D7lPfOV1V2EQsfb4M91qaA1EeMnxPjTTo410Vyi/600pP/
EyNWwCvCbgWNxJNPUyPGc80keSlkAq8AS7be58YEmBeta8kUmk/hHSIxVza4PESVMy6as8187Tz9
YI43ICdsp78JHAhryrQ2VKaMZrItXqOiE1A7j6yTjyQIdEcqvRbpIm6VA22Z4L0yBt/LYLzjpUGY
0jQlLj/0ZXVyrEFj3Gf5n7b/qX27lrMvEc927egiJfjXvbWgrIc9KG2u1F6wXv+HffY2dncn4lIG
mFVOC5ukcQg/TIZVA1RVcz0HovJD1tF/vmWJAo4Q8nwV/fZSa2X4YvC3TiCc2FhieasoQswGn5cJ
eQVBTGg/qKeLhaszFyvmDWSPzE7wSz9754i7q++Lp6Lv0vDED0Zm+bkP5ZhnhnY4onPMIRbGTiTL
4UM/0WUK9It0XxOg3oIAkZ48S6XUaHU3DItiM6oJJQF8XU4KFijZTe0FiuehE7V1y+IXplEZAZ/O
4QeSEUufmxs+qPaGhX3SP72ioyHyuW9UHkA9z5g5vvpCoy87xIyrovqddDBbYoPZzcoSSFN9TBM1
G92j2mNk+xra/xLZPt1SLmhDtbVMcGZNjLqPX0hCsxQwrMwweWmdILDqqg6xanc7W3VdfN0pGmge
0pcXXkp+zbB55WnR4OaG6Cm+tPRU6CvlRkuGPD7bHEixizU0ZQ/7R7Zk5rp92YEmdYFfrFYsyNT4
6jgWMpr3AH8J05yKvfK3TSLAO1zdPIgleWwTc2/XK0/0fyUfoVphPELTvnL2+LhN6KoT+hZ/zkGc
NRIkPe9JeX/lG5YxlGBArBOpg+EjLuBpS3fcFx29Au7DqbTezSO/ttd3lM2PVYx0ds21Tu3gu0WQ
Zm537waYSGogyu/LrAUw/GPEnveoZYCI5lrZsyWlOmqMC3azPhIV3vIgBhKdoV1aQb5V5q0dwRJF
jf8oxOoQkgR5SuW3D9zw+dzfVl7HXiHVNPaQKBL24RSVJoXgz4C2zZNalcoGrnO6zfzuVyYiQzrh
D+8bybFmtEA8vU+u1REIt6bu+/iOdFRBKF2RS+CEiRjPWvz5tf31c5pHjV4GxSrLepJPMYzHRFI+
dc7MVcSYi+4Sx3Qp0Fr7CCZ9XGcsC2k+1ViONRtFXHUWT33fxd8HIv3+PoDHz6giE7ZOS9mD59ud
vxzIkqnRor8mTz4DV5bzo5QoJmIT0GOUKWMcdUZmr2n31Bi5FQNwX26E1ueFnHqh0C3KA77Pd45g
kbz2KJR2ALgnePy+0h+ryB4qFtlEJ9RiuuslNEfe2d7aqKIxHATboJXuusf4olw3yXqJmNBx/us2
6tKgFiJowGoabs8qBqj2GavGq9Ej03I6PxEzclk7UrgXTDHqyLBOKZc99FwvgmxJrSPHT/z66yEB
N9m5AYegDdg/kxLIBk7dmqkLu7s4uR2GOPIRUJeIQ6b4nqDLCHPB/p4RY8agynj3YX7FWZPco27W
Csumk8+of6NeGrCTf824xVSUeZ5XFB6szBL6h/UfiaB/wh7DfLIHGS3lBi/rbJcSJLPu0HnX0vPd
ZuDhPbgnfmcCtXYIsk1Ah3leZKuURzfw6/KA1R6nVpu+qgULM4ocPYpyrk92Hg4XCPeOIvCSCaGQ
fgOq1lOw75HwTs9J0YY4eMsrmEb2hojXt+yIRHTEW+A8zPr0XOqLQAgHDGrHY/2euUk+EQWnmoIn
0cw97EXMwfZg6gWKZcgcju3zliRPNqJ2uPVTN7ESrkyeJV8aXalTDr6MQ0iXZ4BVDZ3/gYg7DmiD
H6ZMCOLE2ZLucj0wi4nKTqYPiMPEj9xVjoyWNjmRKkHcqAW9/YaCJP5ygaejWNmHib1WgusMHKnm
Rd3fsxITWKVrGqry7QpCj7hePYw9Y83S+oYegUqOV7Tgg6QUZgM7UEkVaPlddU6mJrCgWsPoSoRs
vMAhVAagSk0MuyTwzNfItD1UOfrO5dQaaiwhixmV9uxMG15f+RN6oW5/MSiOFuut5alAAmrUxbbC
yaN939Ewuti9i/ACxXT0QcGCFFfSI6eatjTIyxINsKRpe53VD/UjwXuPnv0VdCPbJ1fF4KtNdso/
Z1L2ratBr19u6l4xEyROLivevVlj8j/fRZsDQaWS22Z2Blw+CFGf9ROFDfANQHYBM0yZ2IaAgGw7
943wX3s+SDO8vLVUvAtdwuplMIUzc6j3UyPO6AUKdHAGtfId9WvOKmKDw7jQ+supXhReuYN2aNej
ymyj65+Jub6Co5sEiKmT11TJmR9hhzhkcA0ksV0ifs0Lp8KsKHXCj1t9OS1RICUdtaaOA5OsnuCo
qQEnW1uhxFWb4ebg+79XGPB7PXP4WDzDO69Hom9vAvd2l3MVzaJzukUdBMMOykMkVK//Qsz1fCdH
v0TAmCN+/vi7bws7uzFMKLYJGm2yH1ZQXp7TxVztof+2EvQzdAL4pp8cxw+3/0vb93rZ3Ktq9H8Y
NpsDxrvr+jKRO5tOPrfvH25b6gzfj1EghqgW3ilbH8NG1EvC/KEzcBKaknDRARdZOTpxiOf+rR5p
BC0Hm3PjlU/gtL8QGGnEguTaB29eWj9lxhvPLs2VwqjX7QEYHdlTEnNrNKT4Pdo9AdbXrb0Uf5rN
qTnDEYDVMCg3hWDupfOoVRt5WTz+RiieKiNqhODNW8zT688RsANYpAFVY83cF0FiMCCFxIrtj1xA
g02zQvxZTab2BGI6VKvXK5v8yShSRTZkt/HU0001cYPZ6E//8xWmJbmIwcJdTh4IDBMCQy+kF4v4
DBHs63tz7RsgCF5go1mH/85UWRztXbqAKYrihizrFVzZM/Aw1y2dOHNdsl0WwllxSryfRBATySB0
9aekUBVh3Pqbo3LuRZRBwr1x0FPVCwjJI1m2ZjBlKwcI8aZMvsyFflKc7Zq+ITClAT+qsNrgndlx
h3bW9ku3qiJ/N1mA32/V45jlmjz6PfFwF3KyqwaskjvyFndICIN+F3VVzgpRO0vslVEuLkzcVZuG
+NpoguFnzd0CTrsaXapXyXM9H3EXEM223lNhDEY0KDR96bb59PT3lHP7Q0vE/Qrtnr/klijqymlk
xC8n0z24dRrY8Qtk54Vk2u1dsVJbnPKIjyxaiU+YMsWEB0xnWxn2nVDjgUdv4ZfUbjv20f5b1MNH
J90S5EZ6Cj3eqYB4ovqggiv7mgD7UkNeBOcs4UfzpXq4Gpxf3lJA4AmxQpCRB0IMWUjQM3KIsoze
3j3nBAxkDZ7aimnEy0BesYe60niVpvfHmixGYswTg79bnpNoITOFX+nG/nbTyyAHQDCcbcU9j5TO
9mqcyrI7rMY9t4yAafb108G9cgB7BUr+6hvPyVyZ/PlbmF1okWpFYW+85FlcWIrYgaRrCSklEQyL
KlJF71jkvotfPI+pMJssEp3gnwgJNB/BGtKuciyOTT91MrLqHW/DK5TTN9c6QzCAKC+2L8Ig9ZzJ
BuuBLsOjec2FSScr41tkSclo9cB1+cp+XX2tV8x32uaEdi36m8iNBvakj8rFj0NXkldkWrY368k/
4WDHyh3uBj2m9eueQ9K1yT2OZTgcESAjKzIAmJhLc97zwG0Dmo+cXHZ4ZTQF+MhxJ+NzpKGAI2Mv
tRFK9EZgS5ac9y9SMPEQpU+ZheM3eLlHuHoMxHxaSTU9e8fNdWz8gs/CX+RZd/voJ9p+pero8KXM
BidVdl41pv+bOJbJXTiD2KCecTC1ibF5r0RCeMfCUwwj60c6B91br3Y79qqxtro8r2XCqKOAF9Cp
0+HK2CX4YgLdnCCcN2t0a0hyedNB/CSro3+ajvGEuIKaAxSbDLWL1925bypUvb5DHXMOBrCpQ+An
14xBfLh18IGqG3QKfMDpjLTGjW6UmL3MV/BOX3Ih3q3WcpIdGwsyG5enC8JSHOvRPHulppgOSW/n
4oiiQQ1+J8ObGu6nWRBRJCSI9nCaiIpId6IRxt3suN9zi5jQyCMAxa7/TabXEuetJXkpZGBIbojr
jJakw2/k7Sxfv6yu5jgKboysYLC8TJJsQslQ26ebXepaFasIJ9e1a3Tcz3BT27vGPTk7mXm3luen
2avbWw03y/Zbsxy+9izR9d/TQJvJyHwnDQ1gBDUnKPzwgXixQSg91229ow9Zi/A9Hvc5wVqYIQ+k
63b7CgD15pdB4aVbRqayoJE9TubQfvlXSnIJiXnx2++T8jbvxNMxXElGTzyPvJbmFLlkcX1GjKzG
HUIsZxBxPD061tVMKA3d4TvbhrP1NYO3ZoVHOfoZoURVXsynCc2RCsDWMWQlD3DpLbOrG4v9EUVK
fDwQpzHxmtiM56JdpqJ0a8kxD6C0ixEa29vI8TKfswcYChyVmubhPkiL4Oo8pBp0TX2klUeJNs/E
8UWKM8t6uvDf1HxA0ewML9wK+xiDiAPeIyM0uahklSPvF1T3a4h0NYwK5BtCklhx0W1NvQ47wdYb
irmeNRTD2hPK4jSC5S8O88aVIyHdBWR0lqZFR+dUsmjkMSoCnVNSacSfDuXfuyROa9wl3pFZHckI
nyBkA3BXcYMLS4IkjjP9yFfvsh4U+NQ0U7xPfVlb8jrF2EAdsvSM9toR4VuCrMRHHeRUzWKVaB1D
UrMVNoF5VAQjIkUmJRPfkcODWqvRSM4VMIv3P6QF6SWiNDv3rxqpB0NguqBPoy9+c5JXdzfNSaBQ
6dC34qPCenP5wWCx4NL7UBQYaO0NOpQgbP7X1n7pGUhMiA5F6KdeQuDi/6fh7AorgRO6ihRDE2TL
dmDjTrMnR4EJhPfKkOAlqgItVO6Ajt3vutqD5ppXcAzt++kn6luMszRIUn/d2uZ++pYXCQPcwQp6
CWuGzvBJqbBYd6YKtciCNztrSABmv41U3hxrei5y+5k9C+xWasF2CXPhHMHd7gdJ1/nk+C+9d0o+
yMnAkv7Af7C7/gnvMiDxqeF2EJdr+8ueXtE17FwXfImpLOY/2tCDt3fH6fiiTDD2pRww0eIYSdTp
pgIgbtggKg60KiT0T8R/U5Rbvlhu4He7hGNa7tbBj5md3KjmIJwD3hd8HSwpBZe+wHuAIpxt3mNz
+2gENLqM7GWO476M5Q6FZtj10RJUTZi2MGX/jrW7iLzH12jTTRiajtTVvC8iYOhqxkDx/bPdpnBn
HhabPuZKT19dapo9KGhkCb5EYLnE8Xd1hxlmzx9IMW5Yo36suDF/HVle992UTlIicomECEmYbTeJ
cCN1Lalqcly4yT3NhrIj/whiyK5NzIjkqvNcvtdD3hLyx+kZn78t3fzQdXSl58TVXNQEffqZy7gS
irDlcpy6+N2bzZNr8dB4kYF9Am5CbqN7JVKZvok0p4xQmLm8fyAiKGN303Hz1Ru1f+VUMFqFscsA
wwq5qpDlanOTIPgcTcoNZRCd3Rxn8201Lnj1kd+0lZBVqORUUC5bg+MihM03GGn1fu+JYTs1pmuZ
OltSxg7IYnlzLmsbMbkCNDPyTJPkdoQP10S9h7iMNMzYuLrgcKpfZ2gjXVCqEkWueNigaS498h6o
ek4WMuDzfLXrFzxHMCXXhXmrk2KTrz2qGW5DsAOP+1xBjConcfobBZ80cXv30wOnZGk1Ag15XdGg
UhFL3wjrUexvRgHQ4/gm5BjL1/EqLhV07HLSbb0nZ/esJ7mnheffBsiAcT1FrNk7omrgr5e7htyx
ZQeVbqzxfSadFfzij5qgFdMsprwrtZIvdTr6wYJ7/ApP8LX1x31fN6l0txA+MBbpRf30pXUMwJGJ
ZtETaYiu37Ib/vrWbvXSWKCQzMMCmImVRexO4poCj/ueX1sj8vNh6OewmeO4w2WKbbjn+fqu8YJ0
hnM9Kt5ZEzdsBRtQS9rpiKq1zIgP9U6XKyGcNY6dja3K6tDE59J3/PTn50Uw5R5bXoxJvEN1vhCM
5ac0ORMSfOFsLJSSjw67dT5JbjqqDbggRPPP3qK7stYo94ODy2U0n5ypOMdwrN5not6tg4dar904
PJ5ZoRZjSzBzP0tFbQEhzCsx+mdEfD6zbDSJDng/zXyMpgogEqDE0/qSb2stUe9ZRjvvcTGeWuuM
hdfbTMdEqRq9qe/DVW25pISQixDj5tLHYRzRG2dxQqXPDBlH2AbC6zCrUeLjilbTvWfbg54UjpaO
lbb0o1+6tHcISGou3azL3EQWUj0n2yqsxh/qynCNwvnDYOd4Z+AUFlJL4/G+S0dbFPYzPd2nKjG6
DbHk3IGsExmQ1g8eVEzmLlOdGwkvMZz7ecqsyzR6A2BgS1y6FMJ5OWnvYmhddAjAic5T3BYyM2dy
pkaSMApHs1t+aDDN9uj+S87I8hTmgcPQno7ifBntrWdG7xhHMSvs7HPZvl/AXBctNDV2RtxAS0qF
EN42mKen9ySiIQOYhbxLDfZimq9BuVA3O/WzZ7RLZXH/He6JnitJ4wFga1c7vPGBDqlMDpeomcX8
xp/dawZXrVqNGgiiqPWt5dPR73tKEM0jDvEeaWvwkuU5UbsS43jbxS6PQZr4VM/BZ7qJnmE8znG3
fmu/2oSejBA19Uij/rK0yPed/8kQvdefZF38WXa7HIR6KnwZB7+J5AlXmY1iGrlbu+Wknu6u+pjK
xzyEkmeCJSjZAM9P95byTQYFRA7ko8UjPgEuEmxAbgEOShmxr9HbVHVyrb+vRFYFkx/jie/z957w
TV6IHRuGqA2z+tMqBrLEJctapfJX8txOBs292E6b6LjxZ6D/qHw50dv1RgxBycd/KLA26MFAEVge
P8QLl8939RuZ11rlcA8kvCpTq5+CtyysrHBqnoZKEVqNKuU2W57zMKDt/Q5AAy4dGF2xzw0xDuGx
coADCiUOsGcX/q6w+k2BhvxUc0qI6hSW8QK8W1Jx2Kbrd9opxIOVKath/e2hgRKkW1tW67om4c2T
YtsQRPHXXM5IqRffoRxFOZh5ENZKlm1Sjk9vuL9eIUI9SpansDde4YRm3aqzKF/1p48oxMgoj3s5
7pCS0F4CxlMkBQCflkyK8xQ4L4esSTUDcep3sZevpShOChL/ZRa0X8hhd7Kdz1nylBYxe6XdmGkn
aafcQ5LBHbCJAijvV+a30X2rVOeTG4LHWwQOfFSwptr1Ymu8yjrYriv7RzHVLO+VhewHVrHFdZ5Q
Q7BtwOn8xdU/0WK8QjxObFHXpm3azmllfjizKTmqUK+s5o894XlTQJX5wypM2Vsy2oh0bT89lcmC
LinluBOjA58rUabvNLFGMhmA7S47CaUBbDZ+g2Fg4YUyUolz+LCFLOatUD4v+YYQSeBMo/K6pAH9
avvagmQQbU02n/JZIOZ4cD1kkFAG3GcrGfMNemsc1qe0qH9eKgZvSRARhpQXY74JxKokWYcHlOEx
vans4unLo+6pxmRZIj7NL0On2/5OsZ/01Koz4ogGCvXk7rijDZu+Fa77HhR101jVa87LVMVm1ZAv
YBGamsPfKG9OOI1FZE77CJluba+7g0H9lrcQGV+WaEwlfPkcVjTor5Md4lsC9rduZ1/FqYEtCRxH
PllVDTCBN4+7fwKa93a/0mnUoFIj2ULUt1nejcCak+CcHPIv8MkzOAmDIkwcjFlTcOnJaGqkksnz
uTdgDX8cm+giwp87eZ25cWz/Iyd0sFeoxhAoDGZvFTISp5sKUuH/tt3mNXMgySGXaQkzNcYna6NI
7vW6u8rk7C6TzkeONJgTRYMCzt7KHkExQ4mOIfccz1zU8/wLjzbwSCLbL3zxr5bVaNt+8eKqJwBn
O1e2lykXom6bC+WVkMNGECFdIM6ctlPP1EYlWB8c+YdWBqA0VPnz3N0sOSHvunRItJHqt0AbDMlL
t2POKCMYhyRiYytRoZKeGT9ZreuF4p4j532fQ6ISSfRmH5fzDv6SlJeTVqVFfeCOLDIYbDWbUgia
HKgC7rFzspWcPKrQIgAoh/8QnVrJIS/oE2NwoQ1CXFH+jMe95MOo9AoLZQe3e/7FaImLmgh63gGy
hZb6wUZYn7eQ3pH6X77jtdyoG6RVNU1ANOo0+IP4fzblQqYaSCmbP6Gbn8EzW6I8gJAmjdKk5tqN
M4VmtiTMJkS9NmPnCXhIfzNpgLTCfdECB4mcehUtETXbpfp47sEMoOtKlcO8KUznRxl3PxKP1ra5
i85uDxek0lcXTK+x6sWNPWy/V4CxrElr9yjhIS8Yyb8DuCvjLDyi8Xumn8EhgMcoUYYoEuQj5CKc
eDaLaoRHs4yn80K5Z+vo/wcRoaRWPpupR8XJr2p96MJXHKRDm0d9dCYq+loAnyIrCLc52aKy0R15
UxCdTySQ4psF2AJlUdQrwefSdmQUyjhfmC1tgtwvVQOdXE9v6OdMr66JFZ4X9+YPB9YuLAhyOpUy
YfUYdVGLczvnIUJrlCANS6AARcN+IGSqdqbLbvt/YUs5l1WtmNPTKkTmmXComcbxvwDFkGt2MZKz
3yj7yCcDdG6IChsgB3rqIasBZUL+1nkbvsEmMB2tGE4/fqkFnI4k/4oBlfJeng/Ip8Em9SCVS0rH
wzAe0DYGc91UR14jaWdt0U8f/Za1KS6iu2AmfCHwK2MH6wugix82L1AlK1zaqteUErbmmKpGHwDH
wefOYUXXbMNSNEki2wKhQz14rtsWNbE9OHlnTEWY8dEaMr4e8n6vOFGnUCE7Ppg8gu8VTDEFWV+n
SfJEzwXeXkOp4iuRyZsT0znJri+pF5HY3htEm5Y4J/Cq3ae0cf7fmWyrKsGvr73qBIuGHTzCGLp0
N8PpWqUHJyxBWPoiFJWAuunK0On0lb5nkJy42RrIKCWpLpIVd7Nw9/r4N8KX0EMV5Xdiw99vYsGI
v4qpMUKrgc5J51Fczz5sfAJAhCCXaHaMNZXfVZ1beAi2MMNE9jlGawuS+b2WmqpzvrevUhu2sQ6G
1dgeBURE4y9fvzbUgHk/D+Cm5kmR6P2j6acMlYpy08ReN1Im7mS5IsEZuCCNvkAd7aHBYQIrp45j
X3z6KduFc4Zpi0OYdKx+EgAYiBLAKm44/9Uq6tRLoKaGQ+t1O52wihISuvyB59R19ACcl+TZtw25
dU2NPEQDg8TRWa0zA/DkwHuQzjhPGNtyiDkJdqPfyDqZc18ajkiVWOLxGHiwz2dusM7LqpTsdhdr
Bwn0PjW2yTUOsSxB5Js9QOxV2kMABOVUDACKzE7x4eDOl9YZ94/B1qe2nAULZa/FBgPYXp1f8Mtd
ZA1i48QaZdokPDW8PqdgfFHzyGGadzyr1gyNRJrgSm9/5rvfDxezUqavX6hdQ6+Nt7U318umELQr
d1EgaJywFAgVkUEidynFaiiTHNftMKsOH6B1ko8ASONU+fEva9nKf2thaZ3+7MdpKyibRUBPRvlJ
wwQmCaFhI6d5IhsLCbwZVVq70nuh/8mvQkpQgDwedF0hVaB/oXy4aRHwsBrMDr6Eu7Bj9AOU1tqm
ROyvsZYlnlDtMDOkQ1pa5J3RrAHbAsYQZKNolzMy6owGneY7CnblPd4/5jCmYpPhkneuHxI9ZQco
Mx60yXLeLR6OKqWnE1DYxkmPOEmcVwT1B9E/a90WZWv+EKUApz+GR23g6KZJwU1ewdwVixB9dKqC
MuSSuzywdn0EPUeKasJpHPTe71MlMlpY4v4kTv92qwwo8giVdZem5vrP2IF+IH5vt4H9pC547SMy
oipOlv+eLlmKJyzPYW4z+Tlq0xW75nVMA94q5+SD92zh+KopUvQU5b9Kvibf48o7l6MMFqQ3a1A7
Vhgh1pDvJgMufXenc8HxOsdl+T6fU2O+LGNHEn86HePtB/ugww+69lRkfGPGjkQ2wxfOR4qTuNhO
0+Fu9noNmYTfIshFvZxJYI2ekuioGM69a888YTzZonj0g8IezCAJ7ZD8YMY1SDiuFFb2T/K+2BBR
Ux7vZ9fIVd4pV44UVBiFTq+rSdLAI9FAj/ph09MnZ/klz1ItpSWt420hH4OGefe6t90Ie/3HE7sF
PT5V/IFbnBnthFD8gJBoaJb+LlU+CMT9SUmbmzkoqY/F3SYm5HKkWIcOI7IUOjocEmX5mUnRwCxt
xieesdda3EqCsIjlDVOkXVQWAOt/SgB8P92ywKX7kojyJ0qa/DLw6ZDqS827eS+dBehek9SO1qaP
2ICV4vCAFKE5MH/zXTA+fGhcuwMnrT85/bIH6gY/hQRYa84cZvkGIbwYbGIeMwgnpsZR1W98mUZB
RohWcXqpLE8916oqTJ0/il6Pn0ZUNFXm+AeBgfB0DHVvBXZoa9RA8Skp+5xjNmTw+Z37B1UjhMDY
vO7BhVIuIlKakx562w+B1hD93P6w+BvB8L8fbKbXkW5Jue14Mps/dvdi4QGY5DtCOV/nn6e4pfa0
Oz33wREYPewIs+a7rNnkF+x97GoV1DzdrLQZ8LuzrV9m7arpNe/Tv0A5yY0GJz6catxBjWgnVlHL
7tYZ38gv/Ah699JE4T/vkUAXNtm2lITPKOMX8hfoGaUdBRxnEQaymC3FoCQ/vhY98EcXgGnREuhP
fVV6sY7j5SMsfOZ+sq7UpYu+r0Ny1Ltxw/Mc5HLxTixOV4+sUa7e/7oPBN+/p+WIWa+U+f1SkZpd
uEdiRQCpc0cGTTsWN/qGxnnRr2OHj7q7tWNKhwjhuNFap/D+ft1YbBdDKkQHfhIQA/vjatWGd3io
8/2UXb+FLi92yeMyUVBsKxVyy3FMCYczXxIIFlovhSOmxUtWC4FW3pEGMaN3Vje0bMf/iOVNO2fX
obucmD5ZXX9p5iCrHUQupb24/emnnezrKL6wnbqi+P+NWx3UVYZ6Rh9e8T8a5MfI51DcuNkMgAxV
62bfqIhjs7ecJah9TuKJ1TLpbemV6HZs0ggfudNEEtot0UKd9/JqYJGTVi5tLQOv99gTNJFKIh3D
vSWNJBp9xOQ3OXxhtPgfDMZpGs+iQkNFJy/B6yVhE5TtpbP5J4zNTQ7HL1HbgFHeDGXbAGR98ECc
L8cFlIG0jx5fs38GZ01fHc2ITDaRxoFaOzA4EctK5MMv7rmfCjFJYmUVMtUPS1NUcj/+8OsJ+OZr
jBcthhxibYCQiEeOs09AD8T4mfPXPoPtZvPcuVOol199K3V4CJW7YBjnI+plTJ3xW/t3a4zJ+Vxd
VnKnKoPb2/XiFPDQCftDawtlCUzuznP+LzOpDXxtPPuqk3NUpGGOOWB4MU3JQbJ1RtC2G0POnNWR
xyGzzWn0CadY7odToGZH4AuzIwnIXWt+1w3DlA4ve4UEnXy8+ObOTVtCtV6OBJaTSC7sD0sIIui6
Z83dWYLNxgx0CZ0zOAD6ZZi0uf9hC8W6Q9WGyCBHbHyHBMq/7HoXCIby/50aZiQ3OvmIiTUkBmqw
OPDUWqKb0x+V2dOKdgpE7fkpaObC8vt0eaIwJ9yuUzDz3mR2H+j8i3CfDQZmqpShPFIpn8oy0rtF
xhJPREtJn/C0QvruObpLfRkjYu8Ed7uAntF6P+nKVfUP5eU/YX+NAbswnu4aBSUNXLlvpN9hSM/Q
yKGC6qYe7iZWUFKDanJludAK5BUsbR9oRHzhhw1yjidUZP5Om50e1sJTKJ2lyivupiQIHiFDXCxm
lf/GScRWy4GlWTsILT90gTax+YSXSDiYUP+iazo3orlw6qIk1W2GxBLK/w8svBsQzsCElB7BO55f
x/nxy01ORlOrmPGEKbisVGIQlGkZpCXtQWhHspp1caYAz6NsBK0grJsounzuIkvRt19L+oCXRqQi
9hf8Ro+Y/KHRQuQPkukAdngcIlqYG/8dZCFLI9uAtNcOe5mM7s1eYZ7TceFm7oZU3Lso5tc873Hv
+lXA+UEJbca+TkxzXIAsNqSoh0Pqq/fG7KIwYN8zpLNx2mIJAwDIgfbDQkO8f8bOZ064egun8oNI
FSr6FOFLaBgUvBvOBzDUmVEFeCYtpLwVIAxacAvwgzqruAHcejMC7K8rQVtx+3gfmzj1c8xOLF+H
rBfU4EDzrp/QsnKYRBSdiddW3ox/qCP046BBXG/YU33yzZTzpGCZTZ/J56WzdH6XU9yQa0JapHpW
nUkyJZgh2Ziocy4EtA4nW6V97dngBnAuJrCbKCa3B/RegVHptSCm8hm+yq67FPii4hN8KyGABcEx
GpEyVeEIgmF/M6PYAi/h0RiNke8ZH5NaT0ohH0yWxXT4dkGdpFN6anw+3F+V79tIPTqGcNw+yrhk
BbbI9VV4+pOTiSszdjlL/na4c/xil4gWCZKyL+UUu26kDINB3My2LW9MWxyCpxtYDloQhV20h4OH
ttr5dxU9mto8Msqan1Cgva+9aVkWTr9nsykDgTmGavaVLx4SDtDblILkK5EQ1abyULneZkyYCBht
tfnCNdYj6yymAjuNH0AEXjJuoLAFaXnMrVyn9PmxCLG8zNK2yjdp3D3CzGiTvss2/fndPE7n8IHE
kx8XzPpMoFcdaRhsv6YHYmFvP8GSjRnmDGKCDLDdcTAbrtcxpnpOBHB3rmroZq62aXWO2p3juehe
I+Rf5VcuLdJzuOsJyGOV9bTYHassjdFRO90EnCIKawvQnJND5cnkJPtsUSZlhUU8KbNZNxPm4SpG
f44npAOf0P/ycJlQuVV8Fi8mdymqmX8bvoArliRYjqWz7WPCUXY90GLcd+xmLiuTXkfFQnpNFPho
TjJaTVup9jm5KT6MYaBT9kOxzHDxHinURmlX4fdFQeGcJOHtwko9fSxM0lgLZr3jM7H4GuyamUtU
f7+PpmjEYnnwgp/ccHV7TYwtYBSv89EMMKkUpN/HB+GU/pT8z2njW76xw1C0eTsDw3iXgdPF2/ZD
ZGCjl17V9Z5ZoEnr4ZSbdUTm6eNlvHzrZMQ41aN0WiNEbTxK7YIiJntwtM3KuNCHrryQu5bSIexz
6uoY9MxOIP0uF/8CSc2TCNnAA5H7cHDjohT5Rd1LS44zjYR+NaRS3ex2Q4LIzlHJAFi4Mq4wMJq8
VdFH91039u9JgdgHuIZbjPYnEXbU1HfciXGZ0F5s5nHBIziI7dht2ltx9OHv7ldi7Rj9dQtF5Sz3
ELKLf7VCtFSGQUdFuZaEmpjM/kB0L/KHz5bQnuUb+bzVXLTPjAq25TcU/c2eGkotYYVxHfHECZ9E
EC6c3pPCv2rdvEW7mqMFvTK84I8iw3NTGKqzcKYLGSJ5cIzFvshKWE/SnuPhVQROp/MWsiiiz9pL
pjaxSw4nP+100/Nn/wC0pWQ5iFQovI4eCi1OL/kL86B37tgEqzadMyO2gik7DiZVlq2+tIBTIjQ9
bSXqhudbHLXAK2IYjZIkzI1easankkSgGKvVmmCEhY9WQOciAAREpMx3p71j3YNk/Jpsc2tYkeUg
nL9cL0f3NaGDFdZPEgSo78sDtSW8Pnws6ZRsg9q+nol5QdhJhXC6UwdEF3YN5GdHQz6YnMeclRN2
3LpMriQxUMhIGQDCTc4z5I/yBdFfoNHKHmPkjKJNG+P6fO/ODNsB9pFqPadPu2LH17A7apsvvsUu
ZdXkPfZtGkauVPZT3pzag4UhcDiiLavMbIhqHgoyITe2aZYBLoQSjvbQ/sxOeKQWetSurxgOproH
4qj1Z4cNMSu2/Ptc8H86OHVi9ZBwEXfiwgpqLkBX2+YhzdVFoRH8VYsJHXjjlgRkrrigeJrX3zrW
Eaoe9a5mVnV7voOOM63CWTUuAouHAfW6R671vBv3IW+8mg8IaZcQGOYrXBwNWRJNln40LUPAjM6L
dXi9OmZfBBNQ+oLRTUuDg29ccRe9uRmjRHRsRt5Kbsk1jKzFo7D2bVETDBwMrJk5ffXlPaO3H4mU
SfQwifV9ODK26acvnxvLEfzeyGDxp/uXDW0NFlqzgigtTkycc6uetCc8fHhZclddz3EVEXRh0Zyk
BDGiJyP08V+XmcmPXRerEvWEGVJ3CqZLzRXKqjqaGdrNwYt0vMtXtwWuLpkSkH1gbvZvhRJF4zaQ
v4yPWzWDOdwBoPPIyinLBrUvMRO7G2rjEgEm2YMZnPPiDaMB10bWX9RYGZ133a1vZ33w7HslmGBo
//RQgpSoEoxb+QuU11gpmXQGFLB6WLk4NCvofmE/ayy5/HuKEiS7frvaS5z5KNsknuIxlg3PV21i
4Lbo2OySqWf0ods1IAhhQFxXwoqRSTuFoBEoNc9HqA9gBj1kR0UIR7uH000nWHUmxjzEctsvkJq+
wPSrs8zKaTJP1WGZZDncRxqIwE2ejWdKiN1NeE3A1V12A2XycLRW65fG/5wmMeRRCogvecabkPjS
IZf0OcCN7dbyKD+5SidqgWFI00lJxzirmHi2jPf7gECZhZ8l+gPYpuPOQ20yTk6kac33IrqtNjEI
Ne6DqVFxTuTfFJl/d7o02PeoO4hIOLgoA7DUD08p5yiO2SpXAsMBroXFK9ZlMRR6rWnoavCC9EXu
6NMigayJExi6NcOYlUYpRmn+5bPShdyC0t1lE+Z0imcg3akeQ9OI6Aa+REOh9FsCKjVquU3CEzF0
7/L4xAJVTu3YM75dZxaYOTlm6qW12QiajgkfbmZ8SrNlQxCqia3aYbqarD7KdfZQObn3Smwtb+no
OIGOLC3JuAnWQ40oNWjlgMttDJWlHK0GcvIeqCtgTHOyLQ+ZNOeuqNY2qxlAEI4DDd/eB+uNWAkU
rtt1oLjfT0WMCAK9+jXYGKDzgJATK2L22sDPt3gvfXooV/4QSLIJPtb1eBjusSqWu1vE76YmWkJI
ouKkYxMCDhNTSNAkXQXvNh+aZZYZ8/BvERImK4nBdXcKmsXhIqOIRp1vdrJGjoZp+s6a/PPrbGqS
jvq1CyMlSHB815pbpCg6wSQ/VZ2BP3kQgg+JLrgqR/s+R1AJcXfPTZn1TXfzHhop6fY+P27/CGsZ
uBqyw3fByUXQyi0GbfArhRVofwBlrH82CO51q8T3a7ZOv+p7PUtCfrjZBfdXXV71P2j99l27GAH3
92Hnho3MtfcJPnBxpNy+4FMuTrNVT8Rm3/5DQhwoCbyN5uP4wtAPTTSvrwGs0zZHYjqcAdahxGG5
LGx3P347c4RdiLqhfIW3wYI4Qe62x2C1WDNYhmGmq7ozAFAkrNmc+y/Wng6FvzSl7hD/ho+z13Gs
0qCyXi/kaPgPDxBMONW49M1AfhwA2eUJolXY2slyLuzGk+KmjvTljem0qzV0X7mpFXhs0OnjQwyf
8+JHGLIXGxY/T5lqL9FJwyClMSm1yNF0Pw+Q3OtUz1oetDEBP75r9w8k9YbZHoFElPBuH5jhwEuJ
MUa8Too/Pna3Yp4ztGOEBMmxmIAFDKmhuu5Fg9K31Z+MH+1tAYx+kMdzeWZGZj9m7Qllv1BfADvU
McAk7QOUEJVJSq4YCurcesqCphl2VSo742P/8nAC1ffGjfpY8NDyZU7pUpua99itdI6SDHk2gLyV
B3nLqre55mqN+Pllppme6c8YRH307sHqf7ZwRsx/nKRlpNczEsntm0Befbq49A2sMQ/G9cJ8r/q/
T1b2PTG5eeCOA+hTFslLt9lobWm7+Owk2/c1DW01ZQJ/i1pbJapAIQKMfr/umfcAde8QP+tspL5B
Ahb+Lrh99gyTm7vrb+U020nMk08CPOHb+BysUhImMPH4bzxv87AxJgYvqsGD3kox+T4i3Jz9Xv3d
5wCSN9C4NTGyAQX7yf2yNMUY8coZvSyDFC7F8Yvzx0ecN1EVX8bAPR0SLYdSGjramYGeaPjsSumR
GUS6+c9ukpDkVNK2bAl8lUZZLvaFrzmReQzUYLw2Otvk52DUJeR5NH23Hfdo5Df+rSzW9tcR4gNn
eF7LpVw20YtQjA40Z4/D5l61bT3cmJcN0AfAbXViDKnlVo3U5crfOpWx5BXcxBoVfRScBiAT02+P
HCUw8IOriUd+tdx68vjtwsOk/XlUDp1z6cPmFbV/YiQCbse2RsGFJY7qhZbjsyAFr/+hZmnbjfC4
a6qwXD8Cd1cxzlgFO5S10fPksEduA0gIo6oPMdV8C5IrH/dpo/MTlKbwL+SQtjWzZohhkFTT/0h2
736JOK+DqZl2fymNn8Rt/Ryt+wRjjzkBQ+K4ptJdVNINEw/Ec310sDKiePj9uUFSeVFVaDBOGq0v
nYWCgLJupH+WwgBZ5ggKseehEF0741CHzz2SK7mAnFQjuK5ney8gQwpKws/9Hh+c99tAvQrofK6S
E5lP0yzXBOuMzQTNEOLg1096XYF4O/TykD7KbdsDNO6NNGMcuqrb0NSs2P8hspk5Cwc4osTkL1Ya
U3zV6yhnYwjncFzeLE2mse4ectCHsHPwNU5PlNQo/b6yx8QmcrTCtooUwjCYrIIPdZJcDSVPPXX1
NLtK3fdKMIkAG9RAVoMdpVBUsCnxMg0l7mNz5LYUy852N4+GyqXMHKrPz6X0lqolH0rVzOceaoW4
K2oLaehA0DBW2HSJhgBB1QQ4Ozb7Y0hwd57TB/g/nFujsLOYx3VCBOmOCxcgKxOP/psfCnGl1hSZ
FkaRtz90g4nwb9sShoLBPeAkbLgvKojZW/7LcGJqvZj4wNyOuerZ+UJKCy6sH/hpKTnqMbBHq3N0
ZMH02i430TfCoSluFdUcVMTQu7gL9K0c4dcafIUkoACXwb6lEbfx3xlewP6qme6juBHmtZ448DGk
H+ZQhTrFA1a/u6R4uxh+9gVRRcQSV5wxRT9GP2oOlggde/7R8C0DueOYRoz4z0KygiSPIOTIF7gv
7Srom0VU7IpcLo3HgP8S9QaaPlA8gRT710MIT5vtky5/IrhhvewZ9L1j/NN3uLgRO9v5zgNJew+3
yuEocFzWbql2VH3r0urA8YQlDU4CY0585tP2XbklYJpSQiTt0WnvTE/Ea4+55QL/DxGBBN4CfVSJ
lf7ix5Qv8pcW99YdZi59ZHE6Q8100vjaPoZCgQZe+GD095Akf7G1xUy4An4Q9O1cpZh/XYLtLjzx
t3t5epgfMywMmdiDCW7n4a6xhu295uZQynaNL4l+mfUxbnxQk4EeSI61IVWAWsgM6OJyxSYh5c+c
k8YXgtsoE1Ydzz0IJHDZFxBnNFDeQ3vbEEZnrd5GBMehTe6cInfENqCSkM4di5INLZyZLTBg8YOf
L5+AOypqqqr6Q9+sU1yQaPDyamEDvrXNzF1o2hl54D7nZVYmuV9k8yfDhR5ZGL+dqPdoL3xg+nLl
3M/C5KIcsr9TVFuFbrYcuhEXx2li3LkeY15rIu3T9JpKm9aYZLqEFrh5UaTA84EdIwjbUVnkdZFI
UWUrbtKXdQMBm268sEp5piwIuKWJ0dTH9K2DCj13R56GOr3hmTdfW0M2sx+bZXtj1/9UM6cAO89W
va+psHsLLz605uFHnoH1U4R3qBNPlh7EGk55EHa/I7o+/VLa3H0nlKKM7aYjWcWXwOY/VPjs6o7t
NziukL4hoFGO7zItlPd+N7W9LyXq62f4nARhd/JbK8HAwnVrv4voCzOrQvtX3+gMgnJxTBiAiNMT
XxpWUmWUB97E7rb66A7BI6h5LjhcM1ahPZddnRJy8zTNxMn6T2EtLg9Naiwrjp+CwlcxTuzLsE2W
wB3Vb6TJywUKs4StkFjm9Hd/rrFTplaBfCQjByMYDopNNSHL4FqGHITKWRTOoBuFE5XIIZL7Pxak
oeFPl13E7IkSJ0aHBRV4jvaq0ahJB2A5wfS3IcazgZi9hMElBzb4QPYc9jz2ab428Dp6HW5q7+8f
kgIypuIgMj2cQNLBHzWRNo/OZOLkqmb9PSTv3ndPbWjUknZAa6Nx+xZIAokU7zVVYyXVt8MTqzwB
AcSzakZ9MNMyzP9pLQr8DOmtjSSZXcmQQbflu4OLwMwOYCh7WCCj6D6io6djDFLCBb1DUbehAEf0
AYsbsDwRp6NsAzboIESMXZv8tbXn8LTdfo5ADgeIFjC4NQAh9qx6u/pd2PeqEOAkEmkIRqPbbiFk
GkK+0/K0zzEA4Xo4ybdt/OEELzUsSmj5dlckYnb2X33Sp7F/G1YIRNf5/JE3Ynqd2Ta+AHr0Htrn
OYDy9jZUxtTXJnxKNvHUney9UQe7emjFKflOkJ8CT9Zisdlsh9m6Ahi2WSU5zHN1YkQhs9DOuBJW
9GEdStGxhINFLnClKiLNqXhWicsVzE9QeUJlja4ZtqrJsqA5r7H5SVc0z7vHCAdO1IiqnnGtPtzo
7Hgp16J+oRyjXpbLdqxPuZFLBCInp0KeW5JwjOYkXL6l/FH/GARN3Op2AW4ZiXJLjf7GRGdRHukB
rrb9BDxkjqWQMz5ProE7LU4pwuP6Rip3851Hx7SPAIJQBm0HKX27FUUiHJs2gbvOvO+DP/H/kcPe
5KqKnXWTB70QdXaadLhECuMoKC6LMvmODoGs8+wL89iqLbw9wEMe+DTF2BWDp/MjEnC9zGdPF/wM
OdHr1lmhToBlAwFlj/mIfjyyqaiF6Z0iQVrdNWTYHY0bUhrKxLO2RaPxXFjJUo96RXTWePrp6h4Y
2m9FaLpUDvM8QylnogrBViypydClpcThA46KdL3XeunGJrno1NhPZPkWpYFkO6Qjeng9YEEocA0i
ksNnhKU5a7TbwI7N2WvzL8VTuXCALPa5k1MvG7EFRBT5HHoHlaQ4FwWfCS80I5d+2tVPIbci4Ug+
lSOh7k8iCpfeuL7duPnPZy7XzpPRfGCK1QraIG7DIHWaWDZlpsT/JCHVMMGf9PXTrTrNRGJLeGC+
uVfcIfdXc1Fs7DpOpl0x0LRY1OabuM9Y17+3ujTakIAGxZj5aqAx/6NfMWo953KQCtVeTzANLl5I
LjOSzQ7w2WvNRGk5leMoJjtZLzNiLV/1PsH1gsQKS01ncz9t7lNUVCOp9micraFpThqs+K8w3K2E
2naBmzGu2GOHUVRAQdLYH1RlzK0HE5IEfiuTukqqWl5m1DaqCRUXa1Jcpsl3PBA7tk82+akNTR/E
h5+OK8jvjnhkDY3kR9Af1M2OCfAlYUjb81++X6yquuwW4irPGCTPWqOlo6rcEFcUj1ItKV8AY8NB
5BfKGlrTI26CoEri7AMXrjz2qZWaEQruaojZkNTTMwK20qtVR5SPlnaXETzHeOrEg6TuzD+z0nZQ
THa3c3NSSDSU/l2rxa7Xt8w7u3fzT8fBOYGuD15e5wr88GfaAxuMZ1a/G7Hag7BRELagHT4V1FaX
l5KyXbng8mNqBg8aTatsvivD+ilAQ73EV0Ekuz6lO/yHTsC0uEVgZT4OjqIzsTvssH/ssyvE/xXE
cRsOcVXa3CvwawnO4/AjxboSL91wTGrjaQYYOX7C5QHTsffwdBGCz4f/fuDJ37TF+k1g8RbUZTtj
USbKx+9CmFwFkXuqbEGQfkl2DCQKThtPxezJIzcUBjz0147/Hb5QJW2bpDgG9GmsB9ufDZ5QT/pm
kNETIA0BiKeXa95bZA0JehjhfK6jgCTeKRjTDTWH10lQywy06aoYCEsFQ2CDcKdIXaDT1QlKLqGi
etsPJXXhOiFBR+mQlQI4ABfQJCgGoNzvjC36ma7FHl6eS29walhDciuP1MlIse+0YTokZqF02tdD
CX4cJJXFfDsfba3eSIM1ubmPgx8e+8nFNN6SIwcKTtrsxY6eiP3TabBxLtAzcFiNw5BblIQ4Y3zq
W91yPK6PvlL2RpacIdQttP7zTtpd5I31V4Bd2ZMpjaFM2lfnY6N2QbuNWgmysDnMkacI/tYAmMik
q8ALrhwidSu7Yy+nIqg30WjxkQlHlEdUTnNgA9jsK6kM1kGOI2hMh6qNWhY6ll+nYDLrRGzt0nuz
Y+ktPJt49OyhvL/ytEUIvK7V2/XJkcQCz5v89cMLfjCRNLbcvuv3cY+n+3mSxCC8PWR2O8CZPyS4
szE80SC8WTSsrXvLya8fXUtrxtJkYCVZ/Bl6DzH6BtCl+3te0NchKCMqYWjwHINtDfIinb3K4OdZ
UkSaP9T+XFubfYDlPiHgMsWFxHm3zK0sUj9T1PXoQy/FmoVXzftdKQd9NxvKX23HbtvxSt0e+5cR
aOnrv/9g6QcQx0PUz0VNLOZ7ZmMZ4Tu8TXrIo+vRZAsygh5CmO2pVTbE8WDk4SNJSbgq2KK5gglo
vUPdSdW5OG8CbvWk+trIcJOsfCd+gmCSfj3HEawFBQDeOsWcCKoiblsHdNVkr7m980xMetRLLldF
Kh+d2C5nmWtCoxZsPUhzuIMBBdaBE63Q4ntxX/r3qMHZezYgGNGJ/b/QJccavqIB0gUxzBjNbUMg
hVuN1ULMmov3QWXMwkNzQyhAcwLvHreT+aLa276c3nOcyVXiatBaqkahzMEDGyirgpD5KjiLbDVD
HlBwRQGZW+lPtdeK8aexZTuH7R4IC+U/hiMutO8hQz6nTkNVICF1Yxc6qSAwW1NUfsI2cLHNde5Z
sksyFMvI/XNpjhxyCZ0aqxoX5zhxZvuJI1ao76EO2rUHgg2OZD14fJi6wWHZYoQ8qTvs0wU65B+m
wYw/g3NAFqG6O3F708eLeOpNXG8hP7n28Rn5q7E8hwhd7db46VXBZ2ZLiIskCpsgyBe3I1dKrtwP
nc7yt86hLPkDxEXNcyejf4V2klYqVBqMmYkCFJVxYXZtgboAvGNxsA84Jv/DvZPP5JlRteiOS2ke
snvMHsnmRAo8c+Z1tts3qlF2CnEY9qZW+SYOizQzOUgKL6d88Pn8DvYoe5T5GmvH0E/V1i1qabdk
2CDuVzOh6DBsyEg/G2Anr2K833GhrOFM+eQrv1QatHPQyTj295d/GmuC/0rjUk0rzhL7xwhHW4Ap
2u86xW/VKmodsaqSc9VnniM8a4QMDQuL/GwY6hdA7yfeD+LC/gC2vb9ZLJ3Pw645xhNbZ1ofD61M
GRutHOJ6kN7ZhSH2DTlLnxYTOrDwqYsW7ll48A0fIVqT9M33xPkDxoqtTVRO2xFyHDKvfPSzHfCf
JQ4PIJ0z5lWFpZ6gIbzqC3jCV5mqT/bOeFQgRVcCdeUYY3pxnFkf7gO4OOm6x+amGwWzQ+lqfOh4
IKRUGHekUAZ67gvARIOyDIZsgul025c8KjSgsby+1a9n4C+hlJRLXd9Gqiu0d2k1bW1zYjrPZmK5
lPlCBVwme60qjpoNTioFjdPeeIcTOlbwUjtefTvrCXIb4ReOdPM+u3npydg4e6u0QqmL5K5e7CVw
wihmVxj0EPnuf/ZlcGmVUda19iEiFyoljjguJYurKjx02Y4iaZsWOYf0iEzNgcEfB5fQH//Ab4dP
oBufsqJXJhEQbVXZu9JI4ivsJz90z9sU9Vz1joCrvnyGc0NuMMFy6uGlrOYnyhCBr3GWzAsbCoCp
TwNW8ZdWLxj5D+f8q6bR+eltH2PpKwy77WqR6WHaATznzsrOURE9bCJ2sKs/dm7V2izJ/fINNp98
5bfIu3vhS09QkKrCmyiRH+vIw5iyIxhGrQvo9uCCsQP+sIpPPDdwIKpt1S9ecCoogeLWE9z5aE1S
jg9y0G0CzPZpXehdaZzqmYyH+quoCPYduMfKsDOxxvuH/OvnAr+RQ6R1kVk+oW/xmkwPz3FRsRBu
NMTqxkdVcY0RZYQzL55EsQFpUIOTXQ+woRocRYI54W66liPCGhBBvodRYbPJpnIm9tNGYv8ljHyt
HSoHB9hXOm3+0qPkBbctUsPhNub7ROG93xkSop4lNn9kgnoZcqwl+762x3h+rySY1qo49Z5NRqOR
edCmKlUe414C+d6WM9+LeeVEEvZb0W6q7bTuFezpEOBSzM/Ct3oiEl6CWMfLIUJkhEgOfwf/dl5O
T+MtohLriGNiHw+EtXDaygp1Vkjw4VGsu1PQg662TM7+Qxh2g1NCR1qCVmsYtr4LHT/NmUxb1Z7+
/PGIjbleTuWfJNns5VZoQ/lf/Z3amq6lPbc16GgRoG2UKxndhw+ltUbrQ2CQiDbA/dwHZc5ilWNf
v3iy1DEqXP3vghBTWQ/EYpfPVbgu2D6Wj68LKeCk7ljFsGPRrOY0YctkQqx5YCeblSVx1PVm9M8j
I8ikPxKuS9SiH6HGDG2qiGn1OlaWqy3Wf6mYNTWT446xb98Yt/TH8c/qQ/KpQNYH90G1Sypufj6w
pskLSBS0/lHN8nTLSGGgz59x5TCVXMqjL18HlMnWiBE3RzfixzZ18NxG6lksz7OihcH+iSL8f+rB
S+Aysds3OWkkt91eo9QTc7Y5S53i5ZwuqSu2cWBnmdkYXCIWOHhoA4R6xjNpEd2LDpC8aK3YF0wM
ql9DTZCrp2sD8lAh5dYHQYdaSKb7hj103i67tVysTKSH0kd+IxiMpmH8WDGwHMmCE2WnzU7LhfPV
AfpIuTqCMzLXvNdM5/b7dLunCbeU92SARAQJqJfOp/HZG80elc2BYNhUQMn6KpONXakn3P3qS0Vn
7iMy6Mnrj0HC5YPJXmlHMLz4uTrGWaCZwrcpcDnmDfBavl7mt/tbiI+2fCi/SigUFnK+29LJSDvz
kzOXn4PQjzS6uRoVjsa6QS+YDJ5DSMuJ0v4Jve2UEeH1x0um/EfqfkV6iF2dtBJ2LYwRyjjfEyTA
qEqv5eB1LF5lL5OVt5K0j52UkCvUn0Ba88S9gf8UHJbbA81/bqXvCHa68bQ0ZEl6gvpyg3agHNWL
QLLERCbseuB+p/S+ZFaxwnIe+WXIKK7xmm3/22YAmlmR5BZt16GD/7dv2DnqZIR9MciYk3GKqKq8
6jsKfRwp6fqNylu0/3vzS6hFpjCDQhC8ESn4dCPNGrz0jMWsv37HfVT4tG6aW2Fw/j+Vu8Jl5Hs2
cZhPhfudt3qpk+El+fo7InEQLWc7ky2AAMnDnhpMIQFgFh7iC0khXA/QpjTJv8diq+ws1eLZWKaN
Zbcb/xsua2cQ5Rz1WkiGmpEgdRN8EXsvE9bqPRCKh8hEiLoJBmZadIbMJo4BVDwBfY73IuWgHxgk
dPAU6hdC48pi0Aoa09wpUh/rToYijxw/kMq5GyrYpzWJN/J9HIeQCAE5vkqtiIIamZi/1wNGbU72
7KjsDtX9qeEHX16WHPE62WYt+/Wx6LMlA4RATgDjz/gTAPddXW6i+Mp0FS0BMaA9S2enqrRjG/xp
UaPKFVUlKX1m+On2Aw54OcYxMCeqyyMaghYNMLyQde8vx2z4oONXA0s/AuBtkOiJpRaK6ynst0UV
6+jgIzi1uMX+qpvHKc24/CEOsgHIFsmztDpTwQCehzh4ZniEIo57jA+YT+u6BM4fj3geRSTWRVLU
QkEm+Eq1OwUrYcjvBXn67+sVM2gTVMh9Ikkrf8By7kw+CIHrmZz4NjoC/vl+j1hswA0uGuxrqNkq
sVzbzxqnmF4QAL0N1djzpNPzSdKyMMeYrndbYWx9RC0SkaAuVd4jqiaDWQkIDfYb/I8IHJWUNGAB
07f5ymXNiFwKNDjpg9QFKIoZGJTB/9m8SWi3KQsJHkb5x6aA3zKduSdudSUx8FcsBR7FYB/yUx4S
1XBhHuZKHuQkpe1bCU23fb4dGlCyOthU9iPvvSPeMlPhBhH7CWR4kjGSVP7I2ou6XQQdpDHUKhTl
2vtCKbuQMQvOhWNNW7YrBX5lpTyc5rZmT8c5oX+el/SS9OlKosF1U0zT1BjfG1i8jLpOJ8UfsWvh
vUHxl8umHiRJOn8F1babGTWaJ8mcIsjeXBHBYVofi2+tgL0oBXmDg+vjX+L0y+4PGLVhRAcb4pyS
lGD/WT+tRsO28nmZcVQYwGCHuW06Szbk3OnX/9GkT+BzDrddVFrJ3JBzZ5TMZKuDZKlO+PDBgAr7
nL3IAhvtwmk7Lo1GKI9k1LhWFjgPdzvTSimfDgEY93Effrx6aEEz2l8WxvG2+6a2C0zTmf6Kzrbv
mUB7WNOYSLOna+CDPPAnFYbPo0hjb02Zxa4Px7HjZIXFpXq/qzaV8GaXbUTghMJgD2br+e6blves
zhehAcKO6X9ZRKphg5MxuxuBEyaTrknVbRjxKKJt8ob6zMboLW666OOZ++QiKylII5woOgDoO00n
cAaTlbHMZ7YS77aLxoswEeqFxACtaXs2NVXd0gZJxWAxfmHn1Sv5/zGJiAjuGqV8WIVeWBcy9R7A
4J7z2vbJmLUK+V4ob06r6vw/LY1cpP34FoohrNe2heWRMntotoiC2v+iqcREo7nhLP8mgj+M1wh7
UeepSecvoalesvhrrtbjMte18PbYkdloJTH8NpQTjWmP5Bmwz/OBeiicHMXVw6WXOPo3wdvs7FjD
Y6sFudGhfliS/GBXMSBuTMR3URFshdiZ1glxBUIxiWf5VrT2QgPdn93vACUdq4yEuNiLu3fvXuCr
GM3R8Js5xAfP7QPhwsNt9CGCxu4riw3trf2Dl0I+OX6mcGWOUrdyCbkZSQ9aItQyjxHoLulLd9nW
EriRLj0hxPoa0Dx+gIli68Tn6cw0BHqGr3C2mZH+A+xRtUCEB7yqYH7+IrDPscyfqhYDo7z9ktmo
N7sxY3pw+oYwUeEfP46rS7XAX1ZAIJv24MOrhf0zP5PzdHsa9BvK0UOzJK1z9J0Ujr1/UkmWp3ow
rDZBLwTc8M4tB6oP2z2Qes5q1X9+tWWCScDiqcr8LRfm1PvJKR7PoM1IeCvTLyIx24ga9cL2r47j
8zrX6tBm4JcGeqqt5OQpNfD7WOZ/DKvGbyKBzsHe5PI1jpCzJ4sO6HL+ucmCVlW2wCk3zWpynCP7
N+kOSTHUsY8G0IbxejveJZO8rn8VzhC2vqg9j6v3P3vYgsmIU6Tm39qez7AGZbcGt/2GjaD4RciH
YW/N18m+C+mgZSBheRIlzo9FVwAcd3YseaWB3ul9hEABXXfz58LTkgusPpw+QSmFeNKFm12D4LZL
dPCm34PMqQC1iqvmzDfJe/V42gkhD2VTfgMWu4nl8iPOMaJEA+mnoNVcTzPRUBaZgzzcbJtDh8vG
wXGwiIibZRzZim9NEIeaVL659gygAgvx66f+1H4AzDR61MJWDmFqnGYeoELVgGrmUOLp/St519jx
PrYkq+umfSGdQWFshMstdTlxON6UYYftDbXRMzcQyikoUCrAQFXFFzczyxjBNsKxwXMzFvQ7+c2L
XX9zy4q2c5gReVAHO3AH6biTTNXrqdIsUoY5Ipuskjaq9khi9gTc/hrBSHlDC1hZaO0zBA0YTwLv
TUBljAwCmFOPJu121uXP5sLWv8GC7SlJHEvcQ+xchXCz5WjR0m3cM81Kmno3J2agXsZ61mwBid9B
lJ0e316j7ZuUmvgh8sYsEwIFUsOwQQA1DT1WS5PC8qKeAIM7Fa03Dw39lR0Oqea14zUyakSvQKl8
uUlyQHxMgORK64naiNjAl3I5Y2cysH0yyGq/uyUy3FFy+lUlpSexS6jGWeABQ7zHs9X+Sr3bIM6G
aBuJSWQx6DeJoqlOiocXFRT4cX5rdrusBLgedQnCjHlkVj97F2ID0pf6fS+grNV8yLgZzymOHG1J
mE0h8bhbYw2BFpBXdhWWMpcZQ/KE4VeL2JqK280xSB1WwdT5cO3GAPZU24FG9UcuuAKvdZOLYGxJ
w62dJhLXLZbJJGT9xYBGYQTp7X/rEyhByGlOnxXGTnFYYoMNiF4VO9d3rajz6gVi4samFow5X7qn
aGZL2iO0qTLjzL4Fo7a3SE7NrGvQ5zDc9O4iDe1aLrGwZQOuSSJ65lLDYm8lIaye0+/S7PAi6csl
6SPpRtH+bhxKYohqsQxRgSJn7tMOetxuA03zxrOe6rS359bp66kooDPAUi5QrxO4eMxMuKUnw24c
Ykb7rXQyw4w8rA9H+dY8o1hqJP9SaWlD3lGlcmubXVRHM2IcXmfnOt1J8A9SYIAQ82VQBTtj/oYf
WsuO/mFWSXWReEzYF7v97GidunCOuEtBTTDHMFkchuhQ2s/fCZaz9Q2WaraX61AaJ1JzhWecjZK0
PQaH/uuObW8n2w82eq1UNuhfm/cD7ndsB3FGSBBcCykKYpFvp0pLZ8r8eGdF8Ndzpoy+Jlzv9pSt
cEE7yN/5LmXUn3nEJrAECA+0j0xKo3DHi+9yATqw4RKeWc5OmKIwB2wI9CrhOxhHQYVE8J18Bi6Y
ZmU1xQydesWHyO1F+aL67We6Iax1v/Tk6LzW7S6xCxnDH+TYa+69YpNhRNEV1svQO+MaqauEgMED
US5dM06D0e6nrjkSDycRcHuPQNpyCNhsPIG9r/9nK5ryg31ORZXPaRG1qbAwi7Y08d8d57W2Jn4A
ZyenMeGsJkyJ/RQKeS+MzsUpmxvgXJy8fuzsuJTsRoLdcBAaudx7DKmwK40BJlmgcLPvJoSKK6Os
fe1T/Y+CpeHCLUysiFreeSCesXlfMQNTY/HCUMWITNu/ktga3fJ2zSUJJHW8FE5UwelmvAuUgnmo
/FGlYs4Y4szftvVAHHeZzykjj4I4no8wFazjBk+3syIJtFYSwRo+jK9qIsc/uQrZ8knvW9w2tDpj
cIM/0uW6DgP8W59aIRhhZDSWSFfiq7XNiDcfZr0Bba4jpx1OPO0efDV9YdgKEIFp0kxR7r9UlVAR
t0e0WC2gQdd0pWYItn0dOsYgir0qg3TsJyjWRi4gOpCI/iBTblI4up/+tcI6HwoSq8FMoN7Uy4GP
bwYBQ2XlcmCNQDY31m+ullVJJcPuz9XXOi4X1hSsYKxc5bJeEbx0+9ETmzTSljjc/1uKYAGds9Hm
apS1p1ZWGNVxXJQBe0NAZRvWCRTA5GD4efNcK3WhZe6NczGolRyo4HZS13V0krJHPz/OM4C/07G/
kd7KdHq3qY/1+4awSmTsf1Q4zQmgMHlLlK4VyG7rbP0PWGUVHs6kbBhwp2JAn9BWUl5Gi8pzVuaV
BFnuJfeB6Z0wGxAWAlrj0TKvENmV7wUW5iwvl8F9HZJwVVrvb5S/JN/D6eqAiqhT5pFP0BX0b5aL
BGrLy9FZYLRJava3AvgMB5ky3CWuQUB7cy5CZn1qzLG+kA6dRub4TuQAsJbahZVDjK9XISb7xGte
Upzv39FG+8uTO2dOMZrPAyRvyUq8y0KnX9ncHFJAMwl/3qFHfqor6N9o9a+UHHQN58xFBsXgQz6u
9tsPFdtLYQzULD9XNyJ8/6vjx9Xc0LYn2rUNnMzeGJwTaUr/N6lesZlrdf4c6stLFTADQGS+WEw+
0cGryQY3ZMJ5S4nablFt8EP9NXaKGPkU2/2ObxJtK9wCy/HJv1t9VcjSw42NmeQOT8RLRPRfqSK6
P0bYbiNMQfnpUUYkAE9JlUT9yNHLssdBPOnxoNc2+SwtcrTaS3u401wjCWyUh3PavOpzRnDy+Dju
mpErhe+BAtIQGxZxLLOS4FHQtCbdWYdIL3Aj8bVWlEYlvUsee5uHBM6tzW2WMqyqGEqL41YGaMPI
HWXjaTBv+PLVs7KJ8kmXA8s+1Nzo2v45vVX0X5gD/YYMksZut1EBRFwzDk+iTw+qstf2U3DLZbg9
hQ+2lEBTHi3NS2QzG4oQzBEIio9S8eFY7awxM+9Whytt3IUDn84i8Rmq5nChoN/1vmMLGHUb4py9
iX93C8HWD1v4lbzrOjCw+dKkVYEn3euzsdpqhAJAJkG52y7SUhZX8hPbyxlfXrIwfNJ8pLS7U7M9
oiIvOqIJ9HZZBG48Csf3Qb7QfTkTNWIsLfwLobFshGWyc94zzMbLx10zLZesCEg6mn+qmJWVtr8j
6ZZ7dmVCnkAKmRAAeOoRiOmtJbNjXUICTuKohQk9eU+WA7SmWSRf/8LJXw6WXFxXH45AzksVfpEa
/9vnTSGi0a1XSu4y73UayXO5iBeFOFIdpPXFSYXMXXbg8f43QtU/dA96jKhtoI4UCjITWb1GUxwp
yj2yI+o15vGzg0LZXke9p/L6T1MRCD0PD1YLiFRt75TIFJP/CxYVapiheIHP71Z52XUma+twoCU2
fIgUCkhvlOMeQJehm5f+bJJeCLLN1wpTTbSHW33U/oMtpmGXbv8HE3Z2WoV69NBXSh1PDKDhQTr3
pFx/CnKmeARo38L+/16IdHn6oyr9g48Fz+YyCwjwuD2nFI3MbND/X+VXNyk6IwmKFDCTIJBt4JmQ
27aNJZLzNv58wpayg4oEWpjpEmkWJcf7onTsDMRTOqKna0jCFEur5Je2RC11PQ6NnphhYLuPUCOt
U7Z2YNtYLnJIBlv//92bEUfFCxbsnxyrMzFbavKQgCJTwDFqMpd812addB8cFLq0oOq68HTJl90W
Xrtj/tDiZG8wmFURYPncWgF0ksY1gtL8KTwGY+uS+ELvJ+37PiILzPiKAZFBSn/WVjn+NOJTEvHs
qEEycEdd8IyRvr7CagXUbOGp9gCHGjTk6NgRcM/NAqJNrf3+snpsRFD+UzTJ6h6kgtNg/x+Uwrzr
6lb2usEd1ZM1enaIZr4nsxTsaqsGbr3nmSpiIESRCH6xw7BC2ZQgjfETb6U/fxuWzwB+utws4AQH
+HGnq7co2EyJ43HX18XDae8UOpFmMhV0xXoGGzpL+6DY+2jdhtML+HH4ap3+fjg311gbt9KLtetD
VXM/5GlXCGSTxyV6T9e2znuqfnWw1+aOSGZlSulRUgAWaeQ+w4piTgyyWSJgQglNnkic0q8VvL08
n0IjeqoNPh1SqQvK7EnLHZLRXFtf7dGOHxrXQDJ+IiNJgutN2bF+lb75DIbu1mEUFlaYQGU7f04A
/wsXN3VN9cXEJL4MqMbGZkjJYsuTNS590QPmab+EedPciNMAyyCEmEkrHht5d0BLX0CehxO4WF8M
0XlCQaAVTF2j9jGhEssOSMxVN/jMMuojHMUpJ2tdep7GTsaLz19siKEzwQOBnEMTRUfPCQhbiAn6
pMBV/j3qMnCnoBjcpmLu3KkRZWpXQh2dphiMD68UaLICgc25ygxMVN1yvmAHKs1NhJncXmtegCVu
mj6XUxsWJM2mK/zdS1AfdmXfq2CD6O6p+O9kr5/VpCbHNJRB+4Yv622YTPWQLwcihN1YoMzfPR4O
UgmKXgAUnhRFuonp6LtxmyK8206PXm/qG6gb6p/g5qyWNSR2mEPSbe/9zszAGzs2UoAVeNQs7OiU
XWrraEIWx0+WfTpo9DVxRRorQ6GgbHa4Nuo2cEeg0MPSlBiwykDcK5F6wCNMZpjR0cJeFuGKxN0V
K9sZHqfXmhmO8jiItju/x+ts8Z98JfX3vSqyePaKcP+fc3IT/2ZoMhhtRB4AuHtg6gvFx354uQNQ
l4oylPt7mzEHF4ba7gi3K9gZIIYBkr/sz3eeEyCHLBETW79YlW9R2FUZokb9BmfLcRfSxP9cerSK
thclSSSKqbDpuwhbTlYVfw8Qmrrtbx8Ry4qpR++tDtIUlRdJotJGHYHT89MyjuzU//OidMOI90gE
bZli45PJK4dXLSxlw780J9PKeU0Z9DY63l66P6ugEIdqU5ULCa2YBSejE6/u5t4Xen3cyupL47dX
s1djsA0zFpeBJTdbJKep9chPkLjkivRi/xD4bs5OXxfmmSAKHlMAk2FqjXl7KPfmwawIeeZXNWLQ
VK8+L/hH0+zNEATGlTrZz6f+D8Afw3io4EmlFpbsckQ+IEjqlxQAjxKTUZx5Qxa6g15jJUrqN59F
kHK8HyeDDexVzaY/YB7cQcXF9NtHiPKEi9E3NFtZ7xuWXGkCrGWF8qqGdlf3ctkW9/8hP1mxhsJq
LF98qtQ0z2HtKIr68mOHo45pkvgw6JF4orqGwTlBRaLezKMRQXR6+lcBxt3G/DkWZKKbLbWHFvFf
MQYDV0FxOu1ykt4h18nCjk6rFF0x4lpICng4IfFMpFnvMjyuyyjUcWjI2AvSoNtxr3El8UrszfuB
lrmGIRfjkOOkSufL2qlx5weTImhYB1UlKIyEFkjo9pkt04iqM3R1Q+jHUcrjrIMxNNQijkWPn+mq
C7vXnpbaJbtFFPYBpk9IzJwXY4dEVj1T2JJ+dxFXfEL5mXOsBjQXtHogDFUG936gVaO0KvCe+YPo
O/d/t2Bv5CDUUcyWSLG3Hv1Otc72WNNpeFMOZ3A4bhIFtkSUswMAftPJPisBagE+fIFXynDDgxqO
mXMw2+u9tPTgG3/SHLNmkGz7Gbwi70Tqvga9jCAaU5gkhwoRp/ae2ZI0Dl3WnQQzmtnc2Rjycj52
IB7XMvpKnCRIkmHszU42Kzoipn0/TD4sdm27Uk52HW3NTgWMcDC+Ak44bspS+MVrg6tshx93b8F6
kIOZ7bbLt0o6zxXvnTNT4NdJMUsOmRT/rAymhL4JWJUgnWFmg+HwGfAiBvP+LHHD1JvsFZrNzLKC
wZi7cBewRcp3QmoxKvpc9ngF1TCvze+uytgOuGpeMDoBNCpEowHNayUFmWjqjPY2wD6B0N0aNUSl
SWFVOJga9D1NvYliMCcMs9Jf9R64eb0Vec3w5C+Pk4rK/EnmqFd5qPwQAEgsxG9PtmTONL6TrssM
32d6YLnNEemFxb+UD438OSK0F77sKR09YA3Ud8E6uGOlHL73KQwADRJsM5rzG+AOOL+1dry68Qgb
C/yLvUR6dv2F+CtzK/EjvwOinKa1YpFyGnpPzu8Hhs8cf4EDOTWjS7HfrAQA/4VCH5XcZZAjYa3G
H3CRfc1qolV6LqIRPMD7DqvWEoJzejPSfrYjzfIyXCpNKA2Zotg+6n/Gm/sGZjGpfsoXeRBSvTIg
Q3yQS/dqbjKIGit+MPCSuRzGJHv78IiYKlZnGdw2xskHWzHw4rWHeuyVOPDYzNrT5uOjuFvBoV4Q
vLgkMWZClmUQDDxE9WjOWlPV4ev9vBlxitR9PHftpsIog6wdakLpiurw5TFVjsYcHBZnws2FIreR
vlMniYuzp3B3Wr7bUO2ck7SvEFPzOSDe9Fz4XWhM8UxWO+ACQUNSvxpUbgBeqeAx+YgMMctl3V9D
djcffmEp7fx8NQJTtT9AGoizFZIVa92xIU1rGlSlGmzfbK/WxLC5n3rtZcWCJqpD+cmuMlvJOOsy
oUN4cQC8+wwh6qBL62OJlKrUkPu7rHEnXIzbk+6zOP39hTjpIvyHDWg6f4oVs80gcc+Hiu+JWICq
yOcwtVe65prCglrjwKxNA59J3KSxRrxEf4VkyRG7eDZPuT7GuBJnFdQXZNf9k80OhI+J2hjs0z4U
w8Gx8nKa2H2dF/iuVGK7DZb4MiDPZMZEQD9AdWtZbkigMPef83aOWPTc0mbtNPuwm2mUK+kWTSrd
+4Ds//NC0+EvMl7ClxYs8rd9QT9Eu6SJzrj6haL55ze4fs4mEpIE2UjKblx2a+U4gTxWwp+F90vm
5nQ2WcPHWD9ITvKas6LGdL3lG9vCGV9R+3MeCIdSbObakfP/H1svBcBV3g5e09vLPwyizSz7aO/E
z1u3DjZusXwDgPgvsGrPBpZRIAJdWM877JqFg4wFngNvsv2g3IRJWKgLkurgu7t9Mp2PXVwxfIl+
MxmhWIv3OBEgMjwiGLe6bPGyKEilZX73cw4hC5IZjkg0TilhrifpIyWaO8NyO7eRB8fJXBj63bgp
AJ+GYKjP5NAl39XPVlgU/evbgPKj2D8Ip0aVAEEYC+BlcfhfJ82WjFsqKwRewCxNbNPM/s0qADHz
hsy3xoVYYV7neScvQtKzXERijGA8b66rFidsPSdr8QyNfajt5skv05tiuIUJRqNVaNRFFuX/zpfX
k+Qb5cOwUi86u4FuWiDhaujLNeLaib2dVVRHmiXaci+rhJ1FeI5Mt27UQGAHUE19znQaZzxSrN6p
hrvEuWKLGuS0tW20BgsRgFaUDxNXyBqX7ghlpj4U6nC7MP7EiSHEhkcqxLCArn5bSYsUILAP/f6m
NufqgxrgydXXv68vs1U5Uwau92OU4ELr86o0OTRE1qBtwtPxM23qp+blo3Ly7HPLh8f2D7q9p+Yn
Sd7z0epAdUaZbFXvHQ+oYBA08h05QVHI6TUJa3kIjK2qcerbuY9ERduQ3TVturb0Lx+ha92q+Zrx
koqjbI86O4Y2r/MAqKZY6LPPev9QLBq5qQdSM0PW7oSxoQso1SRLHBssBQ8DC888L48jSLxsefzh
RCKsCfW/yHUWCCBYPSPUmAQ02qrF1YYKo6N+clxpbo15htvDvUcBOeOfsl99mZliezCJaequa6WY
IxbYWXgYXxD4jMCksazE6saxQgYucUqzvbG4ck4WspCUS21M83915wYvoSwx9PaBE/UN0wRRU7+Y
sckFoQusAnwUFIIBt4YdDYwPLd/Jq9ICLDZM3ZCxsrTSQGxOUzogS8SaHjninA2dfdmbuSXxD7l/
pdgV6URxgZ6m4mGud9/aYdnZzV2/I8WCsK6pAYtP7Gyj4yV6ZzxvUUi72t3hp9gg3s0JI+uOTFpc
2fKK6o3vdtZj/f9tHDKu6/X5jkYw+vXsAFtFEqMuy9b6e2LuUoKfcwmvvcT4K5ZbAgcRXf034dNm
Qn2jXn7Q6xiXRuyngQv5MiBn0tpe7++tcuxO1h3Bpt0spzb0EbDwobYxYS+/MbYkX0TsUQrzG9SQ
1/UXjE5pt9yBYX3nRiIXQQ/iBI7hvrcsSrWCPPVN9c+mc9Yl45zVrAigPtPxlitl6rS/tHGw+I3Q
ATt1cG8mVeBjlqLzxAYig2nIB6q5nw/fcWtKtLGwoUUAB4ABvQ/UM+LjE6OhVpLpWuSnzrmeUvN+
ZwNvjkbQ3P39K6wlCyc2nFi4VHbeni8y/lDRiHyjc2ErkOnolafk4Rf/YojaXr6fV1cz2BcV5n5w
jeoZtphwQyMCAS5+y9g+Ya5I+upBtc2xUkZRXetEmqCyLWoR5fDBL1XA8uyIkH0Zo3Nyfw9gLIkC
uO/sUBUjrZzQZ0BvDLx+H1ZADJhgHZWl3ZCTKwyW2lJW1+SKDryWuKDpCr2CA4K3ebtV2bJy4m1t
KDRp9JAJHQ1G3ynN+2EJNmMO62d0jSTowqKixyiCeq+Y837BK8TBT8i+uJwEW/Wn87NiC20X65S9
8I4uWZGo5aqAHKBc71+0jYHfLG747jcr5fIqkLjWktwrjnmWWGMf+rX0MUezGrrZJTp7s6RWklc6
MHvZBLjdjTYA8IK2/ELzdBxRfk2u29Ea6bigu7oDl13LziZya9zNryrjpHI29s+jrHalEfwPF5+3
27gaSMqWC2RP8srV/BCrbcyqM8xD0zzSh0rvCZAxMk9vJ4mOOqDMe6qGF2YzWl7gcVzyWc0BUJiK
4+Xwa5sd8M7qPmB0E2OCtdMd4CBozogKgb2m4Tvs6E3RVzc/muNoAHPLmTDLYjpHEahGY4sar5h0
sIWKl7II5Z2+QPmx8dbLRkwH3vBHa8Hqmf3U9S3SNhzdKEo4wrLgMUgvC3oflLU/G3D1N/92trXZ
OK9tgvKUdbRKjqxlaP+l6AUnaaOVP+k1eLyIIcfN3tjQm6NZUvhlhLGnqra1Z8Bfj8ANikfCvV3E
qwON+QqdKfM930PH2/SlXSZn1e+Fb4dg0tdbwdaDjUejVNuHz0XUuvpxERHm7+mlb/Z8Jf6a+GuD
p/zktk2c1oF1yTCmMzab9LMnEi8oT0O0vt7RmBhFpg/eu25KuxDlVfUeUYZlUnykbW4qgquHMOll
o6YQxkkg0LlwC45+H1rHRze4Ea2Do5H6Hu5+xZQkGQjgRNsD6t0MJeS/kBPMlZdCcPRWczc1P6fl
UOgXMyQHDhdLWs3gTh5fmtvQmSauRJa4+8rtNGwZAaN52GnNtD9g89tqutocUcOyEmYPYQwx+gmm
l62hj8nkqDp80S83Res9VbrcTUgkUME+GhLA8mSx74Wx1eIs8ZF2WnMWVdDaa8WRUM0f+TMEPNpj
LcG+Bzw9y4ZXPKb6SHIXMdFfAx2MXLioi9eqTfDlix2tgYWywW6DNlngcSFm0ffjRtB5AsPUr4dr
gVO88JHNr+f3Cwbmm/zArgtjMAE/vhjixTbQtHbtvRF7ryiHxNfXnmGMbnC4X0Y8lx3N2fewDOtb
Ojh04X8/NmavqCKwwXK/YdLAgxQkk4x3Pes1l+RY131KcY53aQog7mVjvkohzMBmbl8/ueXRGk5Q
GGUvxEHdB47vktlJ424yYvOSMmU1gf4HKORPaJ5mxHdwPgTbUPXidfULymgPbbkqJQ2i0lsCc9oe
ZvP8wI26R7lJ8MSsXdSb4aTbrUskwaCQTU1zZU75vscTV0oaAW87BOS7BQK0mHvyIZ3qO7ffuyqy
45/Jz5Rq2doBl2+7D8dYglZQkUFEfm2my7xtYrpNioGo0Ift3UD0DWGd6A5urqf+7QT3NWh/rLxW
Z8AQ8Ww6y23WqlJoLXQLapQjFP4HHCv2O+9FixP7vbWU6NNZn0vwD1mkK0+i0Z5V6mhWVHNHfOq0
zJEaFOr7i59ZLuzc9Tlh2nW7ThxSPhFAlR1QTdITSwlV0fi8Xdm2nistluhy9it+yW/5eJ/1LjuY
3zHbDOo138RjDDx1aN5Iy/F4uQZpqnXWf/5v3Oz9ctvFCuQ1Wy+n3ByVbU7PMSq1cbut2GCwYcZr
kRrVM7Pyn+uFitAIplHcQku/tMHqFGbzwGBSJJe7PzFxkalPjFlDprEWASMmpN6sVv0L/DkiWCgt
m/a462LPOQPECLBBkETPyPQdTXc2A/+SVEuEuhrVyRtKupJc00DEJk2nj1pB+PIsgDFqDg+iwxYY
4JXd2UQfP+0X+fjzt39vLxK4YUAk6Yrc2ZOmMniwgAnuPG134c3obVAoUPxpPOBYEblWqfwFLXVX
XHVW5h5EJBXMtbBww5uBPxhlIDOZ5ZE9mvytMPkaUJUbOiXtGtxuVWk4+qSlWwUCMXU+P/m31ao+
cr4tExVqlOzAg9QvfQaUS6zRxFHy8R92D/mTmkbeBjdaM5FOhgkzZb8AYFVD5ueeTvupLYk3tyuM
OfnAY9mT3gyS5YSQZmVnscRuwsqn5Th2qlCfrqN6WH9fH9xyRyLb36+MyrgwB7Nz9JXHkkV3hcD6
dPy51tE/ns8Kdll98C/ZK92ziJmeV/tlGHJ264yZhJ3FQ5vKN6uVNnXFtZx76x8/Tq520/J9n04O
0HmYwWRr4VF9Aasi8oy6Ff5S27neFs/jSBq4N43ecQglPOsWGwnkSwyBjxoQcNGEZeImuomwyngr
o2ffCgwGClVjkJfVyHe4Jjl9BiXXEPpW0+E7RQugnETXz2F/M1yEnmAAKmuql9SH6H8qciT3P8YD
o1mN3DAOd/hbCbWuFXCswcpPmwGwTRAm2RP/ILuRszoNgped/Vs+tXMZ8hh3LpRWCHLqC4j4ypuF
dGee4m442iN5q4+KYkfuvFyrAP2qhXPn+XgJYwel3gPZC9/wLEB12BuaT+vs5AFMEv2/DV4AxDou
Is9be0gt1pv6/UiCMJ1+ItyFTJEsj6Hd/zjvbFt42Z2sYzo/PzM47tAf7r/VbtIoTQQPyEuT09kg
zKjfN7FQaj6z34Mppp3ZesWM8YKw3ptHEZWpwVbFlzSZ0h4WIiOPkwG4kZl39W5zF2/5AmfkMxTV
c2EAJzM1l3I2wu+diBcFnhAKZzfwYf9XXpVhPJ6p38rKwo+PuiaX2nGfsl2Ve4qgqIHd+iRdNcSD
9Z61NVBEim/iVkyH9muL8wHNYWvfBpleFGvuJ94qR25NvQHUXzbRK552X0qowZH1gfw6/K0WYnTl
wFLUsE0YQdgOK9qu0kyn9cwan+y70X3ENa7j2Wxv9RATKANa3AIOpylvhPcKpHk3Ts6ejBX3YifZ
thTbMtpNurw8alWacWqIKeV1IjCQbaIIvdIj8OsMWX2xaPGcWJT9Lb1rbl6YwwV953jfVzU/w/mh
SvNgTTufIHO6YWKUX2huIgNgwrWFD7oehRQwBkRkY/z7KsvLCKw+zqgp6qXWOSQ1d69JHfKlJndC
T/q1HlkChv/MAK+bHW7QIKnQE8zsN32SPahA+JilG8fw1eUwqJ/P7Ecvz+dYyO/V68ZAg+DnGgre
YD8iSB4t+WulVT0PhTzq11xk+bkSPzgSwAqFHSGBkCcs0YJYrAC/RL8UNSVEZ67tL7Dn3Vi4mwHD
9kpKx5iuZSIHj1k1F7RU4dT/ut3UidjMgtFr3j6H9MJM2+gj5IHwHu57chdo8BDYvLz/WUt9o8Dk
raEMBm+IgBdbx1wLGKr+Lj7IkZV7KqwMPLtaUHkYxRGCrWHqtw/VuBA0tn5KDUTjqDwYJmk975Bn
gdWUmYsFvGVG/oBBdxTngY+pxcEF2TtzRk3JzvlJY/g1RMZzJpTW8QSmwYeHRF8FBKJ9GF7pi4B0
4GpJrxvH6K7vIg5DHCPobSAXtORNXKvS5m8e7H7S392w8cNZaW2JfyPYqR1ROLv5kprRqFXYgN4g
2bczH/KWgEbDqK11ed5bpxK34ulurPf3HH5y79M8GSR1OueckXnQFLRUMquuPhSmMFdm3FJgJuip
lw+GVRlY2rBGdGHTwrDs6pSq3vFSykTRwxPmmJ7cPn0/YL6xmh/2lcCF1pNZKXPhWIcKd4p9aHsP
Q/hC7PEACTTAPQdDY8K+GyK+sXsEVkV3WBIzsGOKJjyZx5syZnN0Y4vWBkQcl4mkrDmFbp252o0D
IT7Yefex2RFm8KP1TF0Hu9OH4Q29scAoAs/AQbZLHxuQTQBsyiBp/Oje/GUsKJZAJRW1vprR8zK3
qFf0xEm46OF89T3TH4sjI7rEi7SAmJ3N9HJBKDgBD/6VjXKc2S/rzgCqtpW8sLj9y7yFIktWKQwX
IoLzDAx1PbGKhCcMd/g8NR1EG/6wgUqzhDA8cJFCXwZeZbj0GVhIYH4NsVsRR3iqifsAwlfk8UT7
yRbkr49fuuvgrEbAB9aAhncgZWvGztqDADbrNkmsxlI7WERZblyyv7iNEyQhNWyZ118DSoMpGjYo
sD/72F15b63/+6YkPYYWcC2GgxRDNpkYUNS4vRlP80B//QHlNGfw3SApJVNyP+P/QTJVSW+5BBWV
FUeIpL+qSAa/U+2XilJUINMv1gZHDD221aV/cZ9uTwEdet5wrgrRqQPMVw76Kq3Dy22fk5vCpocu
zZLVrA1T+MymyHtOo4SKCJPoJfhWLur/m2hvyaNupxuFyAJIQMD6RIBuEbLdP1ETPFo2m2SCG13/
8drRL2NMbLTmdShPJkfaD2LqHK9SqXbalLgHGfTywT+o9PV/0eJ4FyFkRKKC18WwVgb+b+Pqt49O
qhQ1OFshwaGnDmU02HSmQbtUiQNJBFSyCPXFJ/eosWbB5JeYVCioATyvlJOfCa1CGqZo5ZdUGoe8
ZBp8VPsJ0a3dxRahAo6i1rRV0n/oolLusQBIef1km4a+AJRRec3UYI0yRo8WQ1pR+C9HSda+rjLY
KBggVZhbLWo3pm7eznBbohGqvlG07mL7Aopww4rKSLfcWJTidFkXHh8Pjqp+6XbuPOcsdsmMUgZU
/sN06yEH4OtF6ubA4vJP0vkqTA9lyhRxTsgqrGnaa64B0xTM0uUc5fAxvU2+qD26NF9GCf3uEmIW
ajr0tAU987xl/yz9A4wv/j99w8Vwg7Dn/ZBtR+GSDPnTu7PnlkGyi92KQyVfjDhSXGcDYMjarthm
rWhBECZ6IUgn7m/5RjUqboITi9rmPURslbt3YPd6kRvHVxKHeHYTXOeVVZqwdUs9+vsk9NRn75of
IK9yZB6XwE0zBWKEDMvLakYd1U8b7d5Rd5CbQCgO9slxRc5LkJ+Uw3/YmAwgNo2FWodzIfZZ+QEs
dM1KrY42Aeh0TrgRwUcU2XUuSVxJBRDi2HsBADBGqx9doMTZzxPsrkP5xy+PusACRsb7rBHAJny1
p/GU90Ld7Pghw1RJVzP7O6yBE5YRsOw1nv2JaKlnIwXZsM1R/pIYGA9iB5ldgAcSNWxIGr75a1Y0
DxTw80VjdJXyHdNU6a5Y4HF0bnMT6PPIXXfisy8hbyU3kCmyAua4sUv4oJ6iY+qek9oRGYr2q9HA
9nT80kSBFVA+/OKqTdM+EqeAdNtYAjRfNAN5HRFKB9RP8wpb6Lenx4hsBi9Uj07pyHebO3vW2oFa
+Oy4SiWNSFm7gwsWeXh7exZXsordERj5AHKzeB5d8L6AhInfNKxp/PzNdJoORydCkGCZiFNQKKD5
pWhFJRKO86T+Jw+GRSa4Dov5jeC1wvrLc7e9WTWow3437zrewWMYh+FtQMTTtejtMqWU6MBXsK2c
hXzeJBzAQ1kT+A1+HeFCCv5wmaeGtqgoVifFcSFRkxqmFXEYULNN64FofSh/bj+Avuu2gmQVo9Vc
G+or8Xta7hv/iNW1Tr/y5BXF/qtUBYler8vP1jMbhYx/oOdyorqOQ4DgkXhG/lytuPyPCXAYHGxG
3A3s9eenCvTrM5U0D6e+0y2hIiF16rJI1qR9KulVGkeP/o6o3Yp+PBBhjt5JvyXr9zUYzkUXydiR
InVdzyi4H06WHy1zgvMB5xpdIzZg4Y4/tSk4jJdLPSccI56+2y/pNsvfdACps8pb3aXKyyCsTgV6
3cNcnMUtHHhWJG2fWdQJZtToDCO21dEPGOJt+dMo3Y43h4i0EXB2oyHsIKa3NnjzAgnT/XlNHZXf
mdAlodN2OOZ4m/42wOUN+tIaFqCI0ddYszsIz3KnkY6D2756/1dtuRp6Rnb4aWkO97zh6j+NBQ2v
T+oQGQGybSHCAGQ6XZ26DNl4numiusoZImCUrQbW3LZ3B+b6xfOwUyN3OPt2vzYRuZO0n/PfpmuJ
c6MoV+aHTbRFfE2m4kCOhYUtyfzoJLnmgjb47k/so1hXWJi0DYeniq+peWZiUgq6WbEVioKwdCDD
PJ00DVAtSfnuKoJXoTZxobSrZTj24ZRqClMYvvfwDi/8SlID8wCxnVm0kaSk+AP649+MXvc8acJK
LSQBmhjsXBfASi9VwXlCPWxBj11TuoUECqGZT1riTXfA9Cgc8dxRUedrmsxrw8HcwSArmMjVGK7b
1O5aePL+AcbKA1z1A+mlofBnYRJh/zRiyfYr662XYVQM8PsVycF5ZbYLUYuroA1Y1g4Nb4hGY539
Wn8+T7zrNSvuCt5qUc/zc2cplVa2Qrjop8xpDUqkHMi6t7dETwI8jRj5kxqfOrxdlzeMSJ3eoLsf
3j2y24+B1hPqISfNeJCYw0SZ8PyfWfhbdK6R7yef0yqdu7cxbjtWkb2iXbiMN/g2p+NLL+izP4ZN
Go1A1xvC3PsWWfzqEXEXpW7hAKVbu9tTiasxOMjcxmfr9mgpNsdtvC4Kn6P5H7LoLA9Y7AB8cLMX
9ItGT80/aDgY4g0DTlFelK6S5ga1wkqvX1IuXTaswknJbRYWykd0+e5v5yxidTM6THJ68Mv88rc8
esvGf2BAyaVg6/zCPYBIj56RhgI/PN/zfqHEdrwz84zCjUDoqp7f2M5TAlBy/Essz3W9n08y68US
4iKpUUsSUErCOOsX0hA5YNfFLPWqoT/SoqgoLxMdEgFDcE7If+XQgOEVEron0fhBoZJ03H4BtJUt
rjDCFnphM7J+ER7yGaNKXbvrT4YlO5+33d1k5nbm+HMF7J5UA5JwiTo5uBKDaHREuNnfnFA5liDZ
uWI78v3UgNYxk0jzIwTt/HJqai3myq9Xp2ndHJRu+yNXWzKNcmMdr3l22apD+8zYBdO2IbU+v/Ge
2YuMgwk2mg7C8TjuRsLVect0J/T3GTXqVvbMVaBRTqSJjgMTVsoAOwcrENWwDGrGHJ5fdJ4CCUeZ
GlHBiJak6YiXRiSY0WhpTOOteGVpzoSGcrCd1EI1bi6PYVnrntnekmnGrxd4MAXCr1pDdC0+80d3
RQ+LoMAH2w/qM56eZtsWWeQlFMdCcHFqflPqR+/ThRFuphrmCdT+6drzNRA4HjOMwis+PuXrH3gl
URLFhFMDtXo+LLJqZAZBQrFIJILImPSZm/+jDj3ahch3JHfzE2l0yg01fG1kwTJ3MpqHZ3HxTitk
WwKROxL7RgHfy7aTaEHA/ZP+mZhXt0TXXdf2RDr/W6V5lkpBJLPoXD5St51DKgoQqOT5k15rpJA3
6IyLxijDWFvbeha+1Tq3gp+QvlpFymUEbMP4XR1wGmSDktMyR+9bvzVO4or+0tkjK7cerB6xs3qA
+ifiB04qx6hDLrLzPAx96TNEnjn/ktOUFckBenyNaW8WhQ/pyAWeNI4Gb+p4zEnzsKAtfOZTYXL3
QHKDc7+Tzq2gE8HQzwfNE5JHufZspVGHbTmQ0XYm0ZP9s6cfMNy4dDfbqsU2TUNQpJKKnesSkKWP
uhfVU24X9gbqJ9bHPQxB2nL+ty/Ihf+hcKvM2srOYPSFqaOIrQrW7zX5ZT61ZW9HrjfziKq1XL8i
TBThHWt+r5hap/xnmoGNOR0Fpg082DEJnoNOSIv4qwK683AwV/j3KEqVOTemisOv3HfnPzNjnzG+
8sbKyJeolV1prU3FDGVOLlAupxf0tNcFAeFzW85f6k9nHV0kH+b9qSTsp2uyjXVZAdnfuUoqtzxN
hSO/qrViEJ0z4XseYFDVFRxpUtm4HawxthwUulQA4F7i3dG06c+NOSi8wYzW13rvLq/X2h4HWIXX
Z3PAGDUUz4CUzKSXYpJsmzqIL062fdxMVDASV4yL1li0AmTd93svE+OswgB1V9ZQdgwRIv2XzHUO
iCUGelAvQ5qh0PhTPx4xWG6xJzbGwWufwSeA5mw5GDTBf8TPVOlo/HHantAq8unuXpb4jyLow8Ah
G0r5uw/uPNfuod8lXi4hHzBcyA4HWfh4g1zrtP8vgfWmUamTxE/TJP49vvQ4TC2bn2b10a8g4GRW
eo0enChN/5gVZYlvJ6o+CRxfTiLOrHDlOG/FJ/tJbFyFhDhWCMIlaVgKR+KCsHLgUCgi70RnvPZU
/g4KD2klwX0MNatJEuesoGylV27lsxYXFjam5+yPNZ66J38eaiYZ97raED1CUSOMUms3siDOFQh+
APc1P/gVSDhumhWf3ofJT6iz1Kwc05PaNyL3GKlh7pCEbQPAh/MOWVV4LDBvw7yjBxxGK2actB9w
KMCv/AXViBT9TRspk9TKbXJhX2v1dwMCSeipBZSkK3Nu+vuTMt+FIQybchdsXgLu/32GjNqJLjW0
iN5qePSQfu7tafbm6oTIP+yTq/HgRY04MEZfPOIlqu2lZrleRLHFuw/Cu12q8rDGS4m8BKAR1tCy
aIqo2U9vJ2StooxVUAGXI/MWBFORlV3nhG78kQJTMLWqzTAYDSp5+DcAKLeVnR7MKOoE+KfAO0cg
6/ixDX/s+IhXyrxaLjqqCktiB/69fySynL7jDcCGAODrOjrCQbkZwKPhBZUtumosK3KD72A+9MGl
LHLUS+/swD+ktzqVAWw2GF9y61sBTtf1PUbSAkBW2dCxhQmaQfr+amIvl5SQ6GQUSttNVKTXtPqM
D1FsOAUdQk55/cvWORq0SZwozBjBXYIYWtglpHoqVyo849bTYX3pvwI7is5TIF3dt6N0aPycynjD
zkj39IScUZ+fpF5ojwkcDZN5DEJlyKf9UHuyxCeXiRBi2fhSofhBlEmjNMZ+jIdRMx9cBrwPNpmq
CTqzifKjEpo/BCwytU2LZ4wkzIz1GI+qjd0Wh7bWQ75SSpKK1i1Ztr/Nxftx4j5q2+8Spj+q3cK3
ZmWOPiK8dTPFwG56w/9MHbXKbeVBojzdpIsoKSBeCGb6YSQPpNxHhHzkVtj0pjOOrJqLd4M62oRP
INdXQ0jFGdwtuPFNCoPEJEx48l1s/C2xCdEAFalN8F9k+O49Mie7bEsTyK83ayrpC03c1xplYiqj
Hx8hS9J2OTjdFNesqBcu8wfPNjfB5TCp70EVSVIsPbzqAD0W+y2qAQHBT7GhUei2vUsvyepJ6RR+
HGacir49iedcCijfI8HFRbcojbvNx0dIrEDEQ3FqUYdfdcR28Nk6wo1m86Jf6lEeA6KONfFMQKd/
p/ZalaXtg7o3GsBmyLlkLjhrzgRWWPypvh9hg+QjwcGmPphfwe+e+vBYeu5qA3yjHVFgD6P2Wpuh
o4l/NeszjI1BV+XParG/a3GvvU4tQceVzxy4TLBMFepvQHMkJF01qOCPdoXrTZhPf4+HadiAI2RM
TxntYAMbSpzgavRstrnzEVZd9RieiqE24jGkpKcPf3nguZFLtqpBa+z+HhPZSiMi87NChCaA8Ysg
1KnAr/l8CGTLUr8DorKEe9Ug3uUucbH4r/Bll1Q1ZxwNEharBzEs8Q+/89ytG8zFaJwkCAwUtSyC
jQmBqouh4UcIb+LSkmgK/CyKXy5weYXyLvKtbg/hBktGgeNl2IlMaZH7xBMb23iSA/Tz5hoX9jKJ
2tbRM65vOR1JwPrZc1OTlht4Up7eKFBTDc+ajmYYfXn+ivmj3QMLg3q3iLCs/WKGkZS9xrr2PceM
28TXq0OUFbl6lubLYpa7EcEUe9F8dt5jPJ3iCpkHNjOPkWp8E8V6Xg7iLBq4Ic44b9TvGapc/cvI
QSO3lsIxJ0cwIazCg3Po4Z5NP+L4xUwNqLMGjQYgzCN+2r7gTNdgm1JZxuUuMgp5gl0KjAc5XXhb
GJ0ofJr85Aq5iSKEbgRV93dzVLjs32fYJ1aMBu67c2+g8e4/fJ53lRAyKueFYClOOvAxTJY0jRXL
2Sg6n86PEnoRuCDVXwvXtjAZmHju6M0qWcXU9H5RuMS/1zADAjbA1RWtipj+O8EeIhUQeMa6uvST
4alZIhnhOku4Lg8DdDM+6Th9Z36oafvS+/dbh+VrK3EuZtrpsOo2H5yivz3KhZPyI7uXnIuru5+e
ErDxM1oc04HXXdhDMO7Gb9x5Dg/uWNKAqzBSlxjS/SwPx7kYeJiX8203Zn1EDVHEJPK/Mz9aAVR+
tyISKVf5L2HE93jG6rqZzQq4a6b1Txkv9n5ciID5ifqSZ9aryP6i9JCH3W8ANflm+Jwx0ziUKu5F
BKotv4T45Z38YxnauQ9/e8OeNs/vMrPQlY9d/19b5KKaqO+HOJio9phUdiDmlz2NQoD1pJDbU99u
l7M9ybpa2JuPIbEOlf0En80Qz4ZAZYHaRNnOx8BXbQ+v7oFQP32tIABAQ10M1kog5nYOfcZB1PJZ
7Zn5H3S/eCOMeyP2Aa/+956merQkV+tavN8h4piShDgXblAypkn6CZNj9JeVfcTlXf/1YA4ZT6Uk
eVEFqoAElDxQVZCbMVsHxNt7VuvvygGP5FgiUR531f6w9BO2biwripRihlhZaVl1qDHPFddt5JZ8
TIWYyqe0FyzBR/VxwZ+ZVfZFd7F0Q0OLqRVt3qotTC20ZwmUXRFsQijJ/EzkEa8srYzro7oKST7y
vZHA0GUEyPSVtllAHw8N/zqv4exEKv+655rklzFDJ+SCzrmlLKVBSW8nUaQe/Pr5HgvdfGcEh9kI
eMoYx0iS8hiOjZNfJooO0RagAT/qK73TRTOJ4uhHzX4wXmEEHpP47Gg3DQXc2TwXNj7hc0FTLuyl
FPk+BoLTB/EX1gJ5esyPlbvYDAgMK5V8np/7I/09h51qS0bViWJw60qGSUrTfp4bZOBvuKED+1cV
Ieed6NXxhOEV/mHzencByUqGvF/pJc8RkvtVluGuyR03oZsrZEvcWKy21h/zewHVG1+th81kJxER
xjHtjQ1AU4e25Aob4i9226bBtqa4D5e77A8vPuHWZeajeZa5TsLSkce4AQzawxwctweJ/fJsuZnu
FIYQRP0WIGkpx2dhffRRypF2yeDHizAWVFKr6ElUhUX/f7nhRNtUtYn79oBI3ahvG9vs03w2fERT
cJE9ebrrorrBWpZLeHtjJldY8XNaEvFq096Fy9gaEvl9eg74HAynThmrd2CdkS0LD62a8vx2dRoK
QWPPSTcTxm44AoCwgiZHEHlO+FK1U3ZgNRN8cr722KWo6+67jYIpwQ4fjgQgqOtIz3tZDu3zt3Tw
pnCe3b0gZRW6RTEwK+snJj/ZTMvxEpfUpyZ6+mNn76f1yagh9uQFXO9RD+RFj3svfEv87Waa4Vn4
2vZ+oIBnaECiJG5KAXDT1RUI47OdL+ALHXHAdAAgcdrcslFuvQLxUBcPiSdDLxTbPtL297Y5Fzzi
/liyLp/mjWRyv1WppOFpC/yhadGKoQpNQEs/ST6YRaFtNbUKSBE50J742XhLjIOBZB3PbuyDUZUg
yJY8GFvJ1BjZ5HdtXcwCxB2bE+T5Cro2fzNdjB2Z89TmuaUY6/1teBewfrtiQJg2hSW87qSjKrgU
pPY9tMogkRY3nqjSuGE4mFqR0LfwI11tiQ0w+ZgG0YNpZFhvtcPw+HfypzKs7Z+0wIUq/4Fpn2eN
dXsyf5cuytbWQUmUqrCDFQCGreaZtF67KvR1UuJgLSQBArQkZ21LKjavFiqvr+48nSccR71tPX/q
dgCyzsxsMpYzk8egXOVavgufmBB381k6cwXRuNOQgDmnh8TjEfcXJNuN6wFJTl8Q+rMJjzpsE3X3
KYMD/KLN63xsaZrNp4Pj36PNniAHme0vMQZ9oZ6NoN08SdOXMdy/Pnx7siKwDsk9gzxdqs364GbS
+XG6IJBFki7mOPJh1aG1dR5adi5EcVlRvUWieeGb14SlWdapd8gjBvfDg5Nv8jlkfcLIDBOFQgpp
F1z7BxJsS6uODkBlep4RoxW187s5QpeaNaW+Hf3BkKQPXIjeAmWIpjwgT64GE9C1DJVdwNGg/jre
iyWzu/R/ktNdV6e2D0apgp3E2ShJ7DctOZsI/PQqBThx/902SLoxywubQ+z0LcLAs3qNiWz9zjj0
4pLcxTnGBeTte1lj5b+Hyby25vkEHTNTqvNp1j4AY0LHn4jy51ds9B17QzsIXZkwaslVEYMjwj5R
afd+3bvE85f+IsI0DDXfOy9HxMtw753Y/75lfwa4l6xqP8PvD07PQ5Ucg7nMk+hu5ZkfoppF6FwF
Rw81qqie0OvY27Sq99FtwGQcti4axkhwefZsccNgdyke4o+fnGLOJCe1+ZjZQ4BiLjm0Qg5PrQ0v
C/TMOeny1HS4XIh6R2CkpMLPAHtSopxeTSDSnc3x8OP6faTiIAxtNDNQlC1U9xaAXsMQAb/fHWfn
xWEQ6hwYqb/saPn9NHeXqZVXEjF6RwhyWrnKC8iWU0Nq9L+/ms38Xys743Tha6k5vQ/JH7VtIAxk
TgP/R7QQowiZMF8EZgPFXMehZiPquvnswseNct08q5sEX0o+6MxapOd5Ca8UjNGDlI1P1LYMSD0D
sv9+Zuy5ZVXs7WWjSF7F/vcMePaDDk47o1izwXX3MILCGbpvZi7Iyu+GCSxivtKSlMcQIl0uAVO6
D8u70F3yXm3A5i26HogNltMjREjP1e8hDQawr9QdzYv3vlny9aBvuRHqDlCHEVkWIQFDS6dncxsI
/rWYtNh0O6eBpp7ndvJgK+CvAAVGEWOFVx2lVPArL9okQbbKyJ+NbzzCDXOUhgFhliaShte1Ltf+
dBYsaZDEwO6tEUR25tBRwAp8jVRfBDDQGmlZXex7HBYzo4ZLjRKzBg/OHACeAs4wz6N0UmUIGPsL
xMTAy9SsnCX3HW/cstEBHHED9uqB908dFaKdfSI364rf2RAYSfO1y6pH9jJCu/vvybuh4aEatLus
56tivoy0CJbnZRmr4BEmal+asxmKoQRZlTBnAkr1cJgRowVP7waeVC46ltNg5Nb28XFfnqupiqOD
qVJc0nqoNJ3MtavAQHLFjZa60aXPFmo9ACK3kKzmFoRbFG9sKhdEr84Y54vwbcVHxpp2JImIpQSF
fN/KoJ/TB6UY9npOqyzFoQmG/rFwMA8B53gtn9/eT0m/CalOkNqLXJNy4bv8UKne2XK2zhyrJTaG
9fE8c9bu1zbcu++8xF+BeU4CBT0hvsBuQGxTjoprEX7fVJk33cPOQZOslGadQsTLkELjnDMl7crS
jAxduAhwrojYHGUQlVZH/2sHxAYsDQEu/zQf5CXQtnr15B6Y2YNT0Jb3UJlHypMp74IhVULSHw8j
sijhemr2F5FEZPjLNC0Juk63+atdv3VvQRvLqdoT0WiY3oC4AqL7iqldCKJcmc6Hri8E7dFlA8nG
Q9WILEELvaX611Q7RTNO5G9K5BeUVIL9g/9kQnxNr8fXlWDG3vz7L0GNNBTwkUZlho9jRCuTw+d2
C78FiNMoTcfwaT1lSan4xg6YJt5BwSEN/Vnj1OVg2qe50pVx179MFZ0XAtDdsnvQ4Ehl3nL2rqpo
W4InY9P/SlgOZFyKqtVQTkT2G90bHBb3L9ev030moQJInFM8hsNNL82wdxbiA2QfrY6YzU6pLkHt
6lOdUIpEFeQDTFiFm3cxqBJmP8p3u39splfS9ChhUdSM3IqkyRd0PwMd7EOnt9sN7Zd0us/WhPY4
FCXQ3eUJeBYJlyJUwWAjUg0SgMgSQokW0q6o6VBs/lKY14SiOaDKlS7Yp84qqXgzsnp4Ng6BFcny
9U7uyOUSk6d96gZCPfCjSRprlhEEl+Bri7jM1bo7FmNHs8FHi0L3K+69HgMssTEYUhix/fn1t/oe
3YMUmWx6vFlJjMeByucz3ljFLLDaVjJdCADphWxSjXERZ/3Y4ddH710I0AbfSIpqe8/uF4QdQjrZ
C90QxfYrPwnZrCnqe5+7ujiCvmkZq+0Xk3Jt7lLpA8pO3fvrokRnhIYXzZFhzov420yaZ345GDbl
RMYZEYbmJx+3DFAOwkkst1zFKc50mGXKCWakktTDMbZZRZdRPI9MZCxmWq008/vdMoq1aa2OwVkt
V2vseVdqsGvUh3Kv1O7lu9opyWt9jkbLz5irCeVsJmQGWHA3pxhuSgV/Hd0+Q6kqNv3pTfYtBfiZ
HS5hMAgl/hdIWIsldvaAdDh+t/rlG02jOP2I7SKPj8mReG+JEbVuMqsEFA0QFQI5mRyQ1fLVZGQh
pH7FLqN3TaXgV8yGtXpMJodC1zmMx+iZmEhRBJp3dwwbopOU6oT0YVV11e25rT9CynUVDuTDKOj2
7sXCOCZonaQQZL3+7TgqGUiOu5CKzIpLS9RmBQrVPH80k2zMAfiBDumEAkp1ZJ3YHVyZEGJUPxZ8
eFPPm14W0qcSN+G7Xh9SNLwHW4L18EAnz790Qc3Da6W6Wmbef8bqUkOTHT65RBQL4TN+vDWKtlyv
qEbgjCENx8LHfU3M+JGTdUiVa6gEG73/slTKb62uhX04L6JV5UuqUC8awqhGnYwqG4YpJPTuvhq+
zVJYoSZ6PwBTylGVq+d/2euyeFuxwy8+vRYNEryqS599m1fPAF/EyRwtQrybkKKexbTG+xaIIMEX
XNy72/gmv4HoRU4T0APEoxWmorOJXulZsrRGI58yNJXw1gy6EJCmofYF8VOAyLebAmet2v1zFM2F
kofTQ4y0vsA+e2KYYHqGT5PTmLpu4U9rXKysqg6mwhp6jXBcT+Ydh264Gjq22Rx+d5t51v0ZdlGZ
n3XVx4Ou2NILWTxxOcr/h5l+Bm4GoFyc9QDEmogST2J3S3Sl/OjY6T+cIKCtTF/BchmSvxq8ln1B
nZwlLHw+24BfU5FJxc706Ao28ObMjEqtkFcGQ9Gyj/1G7DkINRKg+/kcYbJjTVnMcfsCswkTm/H5
fGShsfth2YApwvQJLxkTho3sr1KW4KiSMu9fEHgNqdDUXmLKLAXPE9O9PQkDORi0rMJTIRhnB+PK
/+pqYisAfXJ/ekc/HJggff0vPBXUyZ/YSnEsoIeVyhznkcnmtkr5JfCO2DtnORMTy4cKATSlcSGa
nr3KnGq/i/3rrpVnrzCEJh5FUe2BMg4R9EjC+may8YfP6zPsPkpzqDw/DQ0tqglghNXWVT/KcR/R
FF9pM/1zO6cWYCFuTa/4Jh3JHd6Ay1Hs+TCRpRLWclQMrhNFdrs1gulNU0cmlyPQM9bL46aucbQ5
FAdGvLn9EWM0/ccQeIsqJ+zbUaM2wRTb6cvL+uBL4I1dIJZqbYRRXpPFV+MJ6SX/fN6RodCvWweX
EwN081oISccyDFhUQN2IcoHw9BnyUaGRG3mf6nj62tpyPmklROTwyckGp7GuJZKS36KlSh+zWArn
zWTitWkM94wZvBY3pyHojtP/HQj2ZlytVNIMBVE5wL8D/wkzkJAkgc5KORWGZzeftP+ei+FTiiLm
zN3az2uPfgf2wBy5V0dEIaUIMk68XcuL4SKL1r5SKHmlE/U6IlEgYwOmep8EppSJRbZ3bo9ji1fT
pg4K9lYvJ0vi0EfGnWcpKk3CilSYBvijztZbANpt0Phjlca7qaVx2N21ZfnBkwvdmGGdGT1Xqfkv
sTN06XeOZKjK0e94FjDfD5UnMR2ZXJM0yANhrcM6HZHFrKcYb9MHwAMk2RNjtPcaGf4ZtnlY3aKK
YJuzJrlyjN70Lif2jRA6qqmTfdqLrhuyJw8tfwfqHymtwRPuO6WKLltJB2IOgJQAnPyJYYFEdJXK
MrL2IhqPneasVER60eD1sR8GrcMnIa4P+P7W5dAlaquBKKityT+GIB63rgFbhj/3r2+0tnUe/zfj
vBGOpVkIMhF+8OP7TPI2CylOau4tX8ie82WBnNknDpY6hKshjy0p9qE4zF2BQ3lGv6l7rIVr0yAG
eoEI3kEoAHQn+azSfOzvlutT9JoWVBXpG+cCmRRr27x54Z3ZHILEciXtdn/HIH9FJFXrVFuQaxk4
uWg714aLeKt1P0UnvfcOIb6fwrch7zvjxoR3u6Zqx+tHIraMg34kYncxcqP50ixxa6GNpHUFfFgV
AxPDHxMDRxAal2vK6e0iAUtNeydQXlPba46kWaxR4pNBjv/NxadmeP5NptNqYO87YOk4RkwA4YXN
L6uADlUygBnK/ZXHHDuaHUu9isqeQSOPHEfZhf7Eg/XBFrAcOX5yd7xBDnyBwlA+Skf5V8VurN3T
t4YOca1vsKXRWJ2e8hPzzM+DLBYDMrlRD4utRckkWr4aHSVi2DM849snIE7bQNUuVfBDNz9vga2x
Vid7GilU0oS50WKbrafNNho0jmpnm8+olIroV0n52Cx0hGLQQU72DYtoGnxh8tuyh6it5QgIo3PD
5en/n2sHH19+JdTmFVvTli4cl6iqvvx4/YxH+wSZEEWKckyjlB6vT+ntNH7J/fOrKuojZQAO09gj
9G/86vSpRkIsc44U8KoyvAftBBJwGYHuU899srkuzHGuEvgC7uG8H9e8RgDxZX+XNkmBWiCA8oBH
7cfIWejF6hh2fDdfvM8ajP7zSvpqL2JM0M8MzjU+ATDK706hxHJdzwy80uGfKCUStLeH/hwTPw/R
aXpYORYTVGJRfHatpp3c86IoMbO6Vy+StUuwviiS0HmCTXhqDGa+BsdJBUCw35GpEMbVs57Otoyq
UzqtafN41ubawVa5J8i7MCjimSddV2WNbSdOc1H5gTttgGQZH151B/wSfIgsHH2j15Gha0LnF2jr
WVbFOjT7Pi6rHbUQLWZIKQFXkuUNFEkhs87ky8IoFsX7eK4tF3TwalpeE/5XHAxOyABwrBIYWRrG
YMu1O8LaQvInU/m3ooThzHvzHy6W2bQSK3315Tp9PKVShlrBa9S3x17o4J1Vuh83UkfFTRqhfRvJ
7fxS9t+rMIY3uic0yFgtvM2DD//U+O+qtbH5UZp8Pu5ibBi6IAfAmYwxDKZobDlaqymh3oDq54v3
0WpLwxvXXptVBA+HDfVb1LhHTV/23c/kkXK4Tm9fycB62JpIlmURrq6QiCcIAPDQb9e1XDvk/o10
17zno0FtDh3K3gtcYfYrALryJtyJMxGZNPbi3LobOFDRJ61MKVcxuaUjHfXaX5yvUhvdxklcR2Mn
nEHPvSs+WO81b+r1/0f33v+dr61QTWpRwFL8Tw4Vft4b+CpiP6e3noOPz125fl8ROhvRqkuCVyA1
iPPZsLAn3qIhC9iBSElenNi52yVFyfNhwo29LX2xHQ+c7WAFHMmtFP1pps44XbhPfXXOArkyZkNY
HIWkUsIcvYrm9DRj2q2AHMumJPBcisJh41CQEJOdrDCMGsxh7Wab4VhOBawQr6uO3oIKBDMbHDSI
kO7Y7nOCsCP1EQyJxAxkjKzU0gKlsGVlH+FimibG/+7caxM/2hJ/+GmIe5S4k67hpI88MqmbSmqQ
ozYkU1nCxpLmXkrfV1/zXjnTtXT2/DcIoLju9OjvCnief2ILxsA16PbRdgM7oYx6tp4MHnY2AJRn
rNYzX2G/BgjHiFYAo0EQM4spJC5LL1VEh9ITJsw3UseezoZ6SYCWnsFgQjCnmXbK8Lr8/E/nZt3B
lqWV9KvhiOikXyui+y6zJLqjPZDMLoh6fK6+CJRhg6lU2mTiWx3leVcLYZX6QOhLM+Q2af7NcvaX
DmEqmcI0kHz3K1GTki/FtqHnj7EUU0lwRGk/kFzvtgDy5hQH1QfzSu3yCVgY23y/1lY9gAxdd+jV
aUfd6piyrWMcny9aeKsX0RbOlIGQW+M532rWV8F+ZSAveBKLMOJF6VY915yejjNySOLzVlfkZQfX
SaN8nyPCPKYvvz3bC1B83gEYoZRelkED+bsN9+5ZwbUlkBynmAs3kK1vfITuBR2prHXTnvranGrN
KuKXUyXqpyfUNjpXvJZbvphkEJahW9aI55F3mTVYRl6kw3Dshia798h0A3R5AWjAq07umfyzWS3c
vGpmEIzlglX8fbXRbpf2yoEmf6DjNtdlJPFtGDRaCzdHhxSlGPi58RlvREMLZwkiB1fCrWK2vypx
viHUVqkOij7yg5n5INwYHJoWvWogCBHR/mex7kKwP+qC2hzH2ZtAZRPLdD3ZukLG04PbtdmcIdnA
P7KH2IW7mleDk/D9eLWVqELZ/rheqyJQqhTP3zYJS/iCWKGvafAcW+V1+/lePDksNhBLSoolntxG
8Lkwk+PBJxkGVBbXCt+/I6lfZlb0Z0jK3YNcpzHjbk1uo5tGoWkFRGfQD/WNO/mSjLsrcaVPpyC8
8LK5R7jBSbofRJrq6y1/Ku1GZPHb28pspZ/SuSynbZuiItyAzuaeVLe/7Cb461j7jceBqhaU0Ad0
XsqkXFaKJu/HTjhaSMGy0WJG6Za3YT4MGzaLyypWtOypjnj0J1OTxblrIutoa+kOBmSu6nTCJ4RQ
1o/0fmy9JwrzCsYdjyQAewHCjZCe95ELJA5dVbEEtW0GtCfdsco2QMNgGeFP9BB36eJturaItkPF
CWrotK7bzQ3woFaQyV020+bztvJrMlREj+edoIW3wjhiYylZ/3DgtV4dS7aqbKssYKqQkO9di5YU
1wKLevWffIOIpguf/3U+Zx3l9U6ctNzzGIph56nio7qdX8V7t/agAE2rkZdcpg0V/c3L8FUUc7Sm
ZIwgwBreuX7AMhcxliMvw2UvSv6Mu9VvkpoVyISfQiAZUVRFsl5poQnxF31CioWHQog2siR1CP3P
OE24CHAjNPsXkTNZNTac5spDYB2NxNBoPwyP95AsTYVA1JzbsZ4Qj3uQ9kncqHwGlMe773znU4Ln
UNC3JG0WO0KtzJmGikn6n1qdB+XCmAMPZqGfdcy8FzkcLLztq29rJdzRoenr+bq11rtDP7hAf9Hz
YavhgtPkJhnM6kOXvvtoVWxw817yFWZvTbcf08O/0OmuyH1KOjKLbRczoNJFJOjDeWhGmpf78sVX
OcTLWq4b6MiSCJFoI6l1lteHrKKBChpKJNluuOri/xIIoNH4q/XBTMKjR+2Nu3f/pTxmw1eBHwME
ukNqa8v5TfqseYZjoDbUsO9AUP0WZx5kg2IKNpUVK7W2mFTL3n6xKxWX0iQPdGwSr6yPfG/u5Jk5
aLdUlQsscOgDLi5S7i8OAS6iyVExG23Gy+VoDjnLXUdRzCObmSy7dbPKRRexDZfRrAKiCDKyWej0
BNQM7qI3XCw2f9qdLYBCHP7hgeEkobMgA7fhVRt2t2NDKoqXomP4qMtbzF4USS14nWF+uoAF0o+1
rDMwyrH/jcfWdgMBQlNXv5OcLSpjaIr8FOs878vsMoFvmR9i6vkBDy0NoaH7Broszbk1S20GaqCC
JYk0gH1t/+MGK4qAHd3kQpbUm7rlOd+svdCVV+XMQ0aajrASo307owefZVo9IDvE/bbKbe/X44iP
DRssUcYl1adI4aNA6iAwDohP11ZjG/hkLCazoFDt93JPs3JiuuUrXoz5wVCUcp4YFYe8SmNBmLul
ziS2JpITrqMytG5kj18kGOXH0UTm88R7SBQBLAX/gm3QsgLsD2+4vzfC9DItyWjWxN28ZzehMlA0
n+IFud8x8GamwQ+72iJIPUOcrUtFLkR7YQkUH1EtwxvCSfNCtd/4rAWmFL6w43KT8yq77kprVXi9
JDvsDKggky1wmTK4uFQuGLj6UwCQJNH6xTdwpsOUX5Ru3VQr3FgtqaowjeEeJmO+BEr0W9E9R1a5
cK6EtT+shdBxfycat2/99hVgfyM+9a7LRFB2/+3N1ni1g34ThKIOO6nWMrnvE5jIFH2Ef/A1gQ4X
KV6llp0WYF3QpR6x7lP2gtZ3heF6bWL9jeHBAkZ7qXLRvz2CHyXw0h+o6kt4Al7Y4b9z6Ut0y3hz
HydurjiufDnFMVp7cW5DIpQWH/LIQ+vAmb+m2WQXkcIpJrepSHBN7U4J7j62W2JyuybqOVc9F+aw
Zq/rcbzYs2/FapGtik3eUdEEXy068J8OvuebAlBPfBFscYTr/QRh0stg5TBqQeTtAFZxeSl2OHPC
sPjRNMIZPt0bwddjVLQGakC56DPslaVp9hlNkPJ47MTrWNjFzFGK4UL8AkZISjZ1UCGDMjzUapFV
rQfpnHrPl3zDCBvELgeHoiv/i2swphHKyfIU++vB169qVttd9bWzmsO+OLX1SQEspDco5KN4Odc6
Cyp50cya04pOTAZoa2UhHBcfj310p9iaBWOi5ZOP4R90AOTi6yDQu2XH5sWg46mKbUf7glW5IVC9
Cq4ZWAel1ZeLBT882VEkFswPl9E7jZt8PeFpZ2TfvRrPCZ4G35+7SZxiSBLBHdjeHAozAaajE+ZY
fJ9CRezHGPUC6GMi0tD48jAFpTU6VuihEdEtf/PWqA9yy9oMOe/fUTrPcm4O2ymmjvVL74QlZ/MK
9XvEHOB4fFNKcyDWM4Jh9x5BVuYDXc6BVvGW2rnNueLdfEWRcr5xAOgkN3lSMp2/BvQ4x1YD/UMm
lmcF0JEvcJn0LjepVbl2YFs3VEgR+RXjvdAyQkIcFI/jZYy21ts1Tc08Ls73mE8pX9W0d3ijGfvA
AKUAZoWfu9+vbxIRrG5RDsiej/fbiMPnfHD5TSTJWIgMiRsrksYxvMtxRNu2mSJteCmTy35Fy4bF
k59FuD8dC/bLXPiInJHxJrRZ/LAe+hvceI6JDPNI4aDNdg89nlvZsppAYi/Hw24phgLKTKp3QGHP
7xtR6aVKTQk6a9CO4c4Z53yXrj+TiquTwaf3DSGk4dQZB0rkGXbV8iMlndEZ+3gQtJGU6k7vJfqu
Sse3FmgnT0thnaaEFE/fCLu3ZsvhRVC/JxZIU9n5DCkcpuf3Rq1ByLkoqO/N+8GGzrN7PTadaZeb
j3W4WdNNL2it1+4OIyBvwyrqt0GxfOTwMlU8OkmYq3kIjORTIeLUfmzO/jYCOl35vtSc9XGK3kwP
pnr3jsnwDD1wiSlBR4MrhXe5MAMn6oZR9znlIZRW81dcJxONHOV8l5mRGcU9IuPqMhvcAQahsAmf
VSJQbOYbFhTS0Enf2Q0CnPB6rHxuZMFiPtCPofVBi4hF/qBTDeUFVw5XlnMHpM/4nOhGUMV/v1kR
pcVJW8zrzoAB5msC733Va4uzMIz5sZWPiFqV9ToTrNT7wPAwx9yicwiDXNG2qDDEXnz/hxk+0Ltz
wvduSaz7nFji7xrYiYyjOIHJpV3yLhRSPOwUhiGNsyNBmJZdyFx+SXnMB78wpDaO6/1h+8syXpnE
BMylucmxmGE4yPkFn3wG5A9EdnGjHvcfeTEMjiulO6ZUDGGEh8BA6S2pkXmQEMkLkD2aJ4dKrVlR
ifLDUt4BMv9NYYF4qT9b5f3aBxVNdANjG+BFYoPh5VpVWS6RHf++7CKErJI69wGN0wTwrbXlSOhl
7fKbo/b7r9Cudo0jg91hmbOgTBRkKNHsH4p53B4gi6lzFEF2NhMJ6wLNfPTcefg7O8D5ATakBy3E
ZTq6oToeU0HG6vz2UWFmTn8f9AcGwSuwExuu3458INqsWP3fIHKhpp1CoegFD3cqMsOXekdjixcu
zDBQztwjWVdio4MkHgrAOC3NTjs15UFAOZbtywHJVjw8PbzeQdh4H4f0nytl5bIyl37o0luPGZxh
8P6ivi6kQdFDghVBE6gMCP3pK7HrOAen+UMKkmrDlgmi/OKJCAFymqU3aDV/9jY4oSKg/ySEHHq8
gmfAPZ2hvdBWlVXZZgz2cQt/Trf8KNP+wwiQsCaqWfinZge4eNR6bNH1zi59P2Y7FFdHx5GJjG7t
cUoCei5CRO/QR5F9jRNEZ68lSlfsKUUud64JRMQqm9nS6mW+oFo6wYmrDyiGTyiqcPLcFZkLjzQY
lylkRICBcS0uUoFbH2RL7RQUEynjkkkg90WZ8AXgR9t0wUd/7WiJgBoe3drEjGhRBdbgbXBspjF6
iBuxGvXuoxNku7qWK0hy2kbPcwoe13AGpPEIlWEHGvqVEf+yRTuGT44oxEvnShUcd7GLrvPa8zli
DQC9HYHBSGIDMtkyPGvhQiJa7J5BZDNo9E+cPjdY2aYuUANNkUSHjMEieXvttngdcZftqtxr11K7
dk7rRakDfq1Gt1RnuKIlE/+qrAML+Su5g7uFUApVTjw/eBf1mhvx8s/G2Tsko/FeXSV9Z+4zGd5a
dH8BUpcjktmKRvr/iAM4x0wuZVu2P5bo4KIsrX7ShnIdKQqCE2ccn/QDcJcsgsJYH2/f1oaF5CSx
spUfL+stOQ5bsr/TJ1JUC/MPz2BaV8m3DQ7UiKKVn/i5WxWXPTnbuI4lYsONza3CH8gVbTDYmZmN
x1grVxPQHbD1mptOi5w4LiebBz1Ero5hnD+fYR2GmpWekXWFyfGdfa3jS7nCMlG8c7ZbsKlOY2fE
pUSsBMoW92UgEIdPdatduMbnEifjV7xdmgn1DVsaMH/ShdCG0pdUFsCYtT49QOGQNIix7ahvctiw
pKQJvWyPpxk/nNs15I7QHvxYcFIjes/H3x+B37hDtc49cPUwTd+uhFbOEdhKyS7NP6vpUG5ktVjs
ZJNSzvcOe+afAHJtpdLVdK37eFQZkxIw6LDopuIU2wmMJgO4PYMBQMzIUDPFdrQyn2It3WUoGrg9
m1D9w3cOensw2j7MP3f/P6WHbyMAsxoG0wuhmO8up+/+9do8ELbv0Efn1BrnQ+vdYUvwmChspeXI
GQnMpYLkm84H8NHiYwfERmtjg2f33gYDbhA4rvADqrhMwL6ttIHdEDY0C+AFBUS/oaz81k4cJdIv
F5IenPlx+81wdhToiPCgrXWCD+kU6CVdIv+OsTpfJtawFkPCId1OjhX5WfgnP817l+MUCH+/6ZlK
3YsLAcX7gA4gm8L9AJhz2km+8mUnNh+cBvreummLxMaxt/Dz+mjMKnBU0X/vle0BAaFDUDYJvP8h
u9ddeD1rqGd3JHB8dj6R1i0WatroLn9tlZtywNnHe2uyIrk1em7k+ea3Stn3+vzdzGxs5r2GTSmX
CPglXejWs6thypHWtFuqUiJRVLmGlcJEJ4V9V6sLYAefue0fIE79/OdTqS/1yi2eNObWexZTwAau
CT3jCf04c6dAXPv5d9CsOEtWYS6Dj1XXtH96K14CDXuDVHpZJEmzSgb5gSCkm3ecm88Ylr+QOcWf
16WniHpebdx8FXrB3+XCel2d3s6+pDBU1J65fNoa8RiE7sLYJPIw/0WWyASzk7uEbo64e0kXAgUA
bX6YTACc+jpahdOwa1SaT2YzWllKxXn3sh1SQX8/OyoHgZvUYhpPzgUe1YdKGZuUqp43JB/bUasV
cPtJzd8a7NIpcMZMGCh080moBnlDnUtbRLGLuXc/5DcKCJ9cNQw42Ju9XWRAPBViI6S7wgXjOeGX
NqT7lLpIV98uBWNsuMPhgLNfEWDiJqHYYBMRm7+F4f10lU1G+pqnvwz0aqAVgdDUw4XBd4TFo0n7
d60x7YNM9ULvA18Y9GZx8sg/1yN1FpnxxeB7WGbrO2c3Bd3lw1f26p1YyQ7yLFMcfnJGYt4Aev+i
6bfMS/L9nlNn9d3owb/G7jAIIYBjcgnMr80Puhy29zlPBTlO7uWIFl5z0b4SnBl3v1BBsMgZuM/M
DJloGmgylYhO/gtqxE9IGYar+O9aBd5JiJPzNI12f5wfNsIcqXdTZCLanY6Xpjd7BVLcFwi9ugNx
o5OxnjOKcLZLEMEIcNgiuT0eiE3M0aKSshU54es9nD33ScGdYZ0cBrKRIoUMIy49/+r0xuIaNRRD
/Y9sZTuyOBaXEsqU8X7VYeANDH5ZCxG4O90+gJEfhQ1e4VP2nXypiapsilu6EBIx+u9OpWvL43/M
JbKxrtGAChuVQeoKLor4OFEPE8ZDK9fQAT2+zup4hJz8H6gSjELqGbzcTB8sDyQQQIv4rhAAFwiO
qlfLo9uhL9xupukHpjIOWMz5xwQtO6sAIdFSBv1L++ifSv8KXG7G243J4sJPwVyIspzHApHbux99
ZDCsHbFbT44t0tTPrM89fZPG469ku4QAIYy2lr7LCIDTf6Ck3z9xpwfezmE1kKiC2SVcup0HXOjU
gtY8OCx3bzR4dv4Lx1AXlEvBUTxhFYPXQDIRVpKSB7z8e80n2KwKD1vhGTzczq2fq+aevyCQu3Bl
5lFFRSuUSifPJMMRa49Dnroxl3HdYLJXvwDaZccO+OuS9RaB9HvUBSw7s1np6HmeFQvsRGGVaZr4
8Lb/VM5ngTbPeH4VLfCg9lNXyufDj9tIPudrLJ+y1UiJRo9r6k01lacAegVrt0Ji6GQ7fj3cCT0n
m8yp7WeQ62jNktQgtznPBNZMHHTF1qqdKnVfkrcAVSCKdOqgCv/PdqdODzeZduOCuMy3U2yzxOjO
fWH7XBLr4WVq2/0b6es75KhyVOJXT64W26nqcsVmvrAo2hLUfzZbWPIm5KUagDWqShr1qFaalK6u
e/pB1P7ynbZFSZADzFQ9PfRuigRnJABiYctlF2SaW5+VO0s+SAhy4SXnqjYHOKQG1oZEWpZHGspH
1kdgXRAOE0JTqdPxMnNG7Ot5fH1Lks7McJARuPV1pZIWf06DQddeOgQqaIcIQZSRc0MKQaUqpSjz
wxwWUVLt2bpcaAe/Wl1SMLfB1lIVe+kLbiIkwh2ATpmaPHO3VCAFVodOeZ9auxZ7Xiq76GE3r9y0
/rxW/M9yO1hquJOqv9rjOb/72R/7UJFsaOE0v91bA+U26nGIpzYH0NlqZd4GkRNG8HFQehdNEILf
mkpmjgTpDDiTQ4KAuSrAglf9kqDFOuzLo1CfcdaHVJWK568p2z3zZwXdFdJ3MfzovPjbatB5I4pk
1ZQMhDf2YxLNeshUSHQc1ebOspmBvOFNVIlUAdECvRlr3e5ZSgasD6uwBOYHni5deBq+ccE16Y7L
Dpbfu5ZpGC4AK3AZ6lh8InQAYVX1EezD7j2fopkpXk8VQipROP5+cEXfFUdKMeWbF3SafXJLwqn5
glDu8nj7IxcEO/WYt/G7k6Vv7eflMR3VR6vpkxcJwo3hnRHdmVH2Rt2dtXJH2Jy510yZ2eWdPZGI
GFc+wMqljzbzpQgI8afIvzIj6AGFNVyaHShL6T3pzK/0J0EhDbugYttoYg0ijDZg2pibH/R4hUOm
9altAa1ZUlh6gWRU0gH/XlPpxPFRn+iuYFAbfD/ZmT3AQwKleJkVoIMmwquChl8z+ASMpV73erNY
eOq+CDtVdr+VvELWGLTI2G1Ux6ANmPLHwemEinIGokLSyYhymmcD8eriiPdpQHlmGZ4s+taJY0RV
lj5BZCuSpgigGy6UcRwfLUzvxPENFgubdk6mfelWj4nce7LS/EtnHnOHLZRi29XbW5v3mBGJZnwb
CSrxHlt9hCREKR/VStgR87hSIv+skL0FkO1e41RWowgnuUKkXPr/+JZhxN2kVbHEA94Ep1uwVf01
JpRv9Ar5GVIvh5zjmlmdwKhjZCo8bWMFG51egCYGRnu4r1NI9BioEw3lJP26Khq5ehnReQXBuU/N
5huqDLyxayESQS6gCIygpeKER+Vn3TqIPbLd83iUCLNf1Phb4BP+gVSL5DVlE34WBEg2JHmTJf5G
1WtnsLm0MXek+5Y3uy6/BdqixASzmkfr3n1p0PepypdTTm94Fn0RXKOx/AbGc6jxpR92I6ZVmO7V
/kJ6sokmCwgp7ytBPjpehH5DcKyeOzaNdNs737dANV/IM6RyUrxEnkcmevlJMzx4yizA48biZKwe
4S/uYwin8RtmtlM1n2f7mLRgelE9C0K1+GZ+ywFovcd+PkwqtzKDLMdM2+ZXK7w2w/EkKl4ZB9N8
nLh5AHQ0pq+rC65s1t5ki27OTnD030wpnIEG5CBLmcoBU+76sLVKvYyZeXb+Q5M2QBzL2tfJW6b5
iSWptkvMSgk/0NsA9Ju6vnCaTKFdrMnJoSdhqsioDgomIiQycXJaR0iCPwyrNRAKdkXpnERXCaEj
C+FIcnjGuk4IPan4qsYDnLHOxvJ9j7RhuYC+hLwuWTzdstE22ta4PhIe2QAI76Nz4RQ5bc7voPi9
hUv29Um7MDZy7NdI0VqGZKBvasin/yIM++CWkqRRVg0YY/5fIHfoQKT79EQSugdjB7k5ZxcSwga2
iBiG4jgQd0qYtqHODjGa+H6gLmulFHwkFE/MDdrhNyxUkuKVGmhiTZl6p12EvZBpCytaFp8o4tIb
ZZKnOVFEreIoYzwcoonwBr2BH0Cj5K1ZUL1w8wNtAPW/Xi5sNTDo4KMzWlIrVa5ez3otZdzHMNaD
Rw3OBfDqbWJ3QK14UTlnFyt7ThI47nfFWYE7Pbi09VrfrOmtVKvOkO4nUUDEyt+pSe7Gt39kfSfC
eElZs6y23aCBMn/EJqNrIolqaj2QFbGerzwcDagnT/ryeJGznkSCY4/yId1WrJkhUHrqrT6OQwiq
j+zrOO+hJAfnL6sSf4/Gk/uGz+sszof7Cu2Rm413aGtuyfbvX4Z5qn7Q7Dq1Gr4EbeeQLEZPGe5v
WabXf1Nqkn1ZCiIHuqSoXBqn1OXxf8h1bac3hy7XO1GNI7H88QE7HHA6tD05K9lUZaFXsP7lT5Yz
z9HDsW1ic+JO7Xo+/4CDL2ykGdBZ266YZulv+mmwO9skPlBwzGsyZKmDguRw745ecAk6UjnPTCfd
7dKLCV3J+8KXd0IXcAzz+m5MSi1mm8QAiUATnV+Lp2thsFWdpVRSTuU+m7UjJY8EX6UCTKwvReiD
6zkX2PbC81aUIh4iRjB8xfAHiWnkkToKh9RNbpcA4n4cM5c1o848GIB+KsvGGEwZgmaqO5XcSnPX
Jw5OQnCMqmypG4JjOUc+nyMvwk8eXuJSsXaPIG40YpPuXrqcRx6xCizbqbbw/FtERuhVhwDlS8NT
Y6WW2yhf83ZMtUxounSrEGU3a5k2I5XAQguM/8mzn4XfJE/y0eWq0K3h+Hm1W+gf/mBD6Fmr51ra
n06D/FMQnxy9BeyahsqIIHqyfDfmyyWngQ4mKWO8y2TSh3MOiwkoefTRwEet1eWaCxHS3biqH5ZW
sjhVLiIhj83sA4099dD0tBivjokC5/dzdAiAnqshvTFiogRUTryhZSZMNk8Yxla+EnTRpaPsgbIV
vv7eU6euKWSncGSMNx0IdGgYCTXXOyDdx0bsCsv6wfzUCZ73iurvGwnxmUhrE6PC7XsNMMTPqOzs
Zdnx8vV9eGuhESylDl4Ss+e3tmM/cBH8Ram3nxLrPqMuBB4mM9TMWm9nXhi5WlUsvwFhpLEL/GvT
7TrjmOtkRWe3LgUCUctHqBGQK1pTfsXp05JzIITMD5uyVbfNwPN1WKbdf+m6SkT1ver+6T3vsWde
qmCeH8HuUvd3olR8FS6L9KjqNvywckdNzJ002cZt6XXK/x0aKiQU7xQiiNda/aF/vIIhCLNz2MkK
UE2w0IErf1nnIT9QdCKlcnPmXLL4lGjMldowKEczqz82M6bvM7c6IHMJH3Yp7G13ugkC65Lf/ETj
44YBMgiwP2+J2xRLPIc1imltsaIFjn8gjLNY5jnFUkKh9oPp4tqmBcZJIYTXdfjwt5lVwmPlqTZM
nHPQgbXO/SxRmRjTYDG2KyiXZkkXE8XV5AWWaChqysWCLoPazs6cIJ8lsJYk9Gn+3TBnQeUnfcqd
3suI3V3kt11r3igJr5q2AdLh3dYliHSWIZTE60AeLavvQPB4sjMaWUOpKVnO4xPmcKUGS+sHMMWf
HgG0G+OF4Yc8TxgvUcomYf+H67BjkgHV+eE78DN+hOfe+NhBBW/iU79OT+iXu/AHDkTKldMSmgtP
2EenrFAcoKwvP//VjRZCekWELSzLpGPgkZG5TH0wBl0CWXInyQm6OD1QAZOXCzNEnYI93+Wf6dB5
4aVj9ZWfvlHfQY5D7I0FuWd7fiFUXS5XKIj/MbwPFaMbBzDsTinf/JUSl7n02iE8ybZvdxRT3m3K
FnpahOVXJ+fpEYzqvFV8dT9WvKlv/eZH05CRxRl2s3wZTgqheDIMtHyZuMfNl8TJV1OVJjdoFTvV
OJ2+5S3SNN++gbfo3c7PDujMT2bCf+cofJML7NRbtDyKpXGRJNlk3rqeYyGsgonaSmpOYxK+V1D6
+EObzTQgQCprcDxsVnhjkm26J8tdboC99xjTeLG3L92+ueGBoBqfUYSzNZ+n2SjrUVY/LwVP0Wc0
f7qQpFYd7E8A1mwHDCxE1Coqmroqsv6z6lWH84OkVQXLfXqS/ri/Uu0CNeC4CdmmZdFTFAdvmv0h
LwsbskAN6EhmLvv7G0hICltFeu+8HxUIBqJ4qlnPSnj4Pn6+tepKtDkQJvle14nGR2CuD0M2V/lf
tN/xQBZlT8kcswD7fR/FFc5VAIVTQd/9ce8fUyw55i1BA5QZ0WxMTq8CxlHqEl6KSvaJtfm7k4Y1
VC6KohJFOWOeWgXWUm+MwBa2/jQ0dBYrc+fqsZyBgEPS9l2igK83K2eUy7juM9tdC8nmcpMUZbQ/
16SF/PHCyjJO4HBMMiHGh16GZlgyb2scpOgX3AsV3uwJPg2F3sHc47AhIlpDhvAF3quqYB99HgYg
plLlmUBhZWfZADR55+BPyXBqaUik5ioQsuBLB+fWmHCt8vhAiK3HZn80HXiCM5O95SHtyn/yiss7
nSS15OHdGsVl/7Fe6oPSUU9TeqZ+iIKzkjurOuuY3zxYwWjRHXAcw1xOh2gDpNMvIMggu4yJ7cKm
gBCD5Cogn0me4G8xmSBkrZSXhqF6pcl0x88dFhKhUtWsDKnwDIIRDOcySu6SBZrUdLrOMP6HWH3G
1uo+YNpn1K8ut4b1UADcjNnkm+ToFHT0ysVpNDHvL+tj4vOxy5dVvUkysl7XDy6WCV1JXXqK17MP
PmYIB1I6VJTrGP5NpbRYkPuI11lgBPzwWRWUA1gMVbAE6JlSIv2kKLVFvTEQS2mHGEW50bo61X07
UqB5vUGDWCkn7qfHxSzgFd1Ai5UG8d9vRh1Mp+G5wcuGTXEhREBhKF3ovwZFl7yHW8PDt4w2TkES
sOUXvgJIdznyHWhNq3LSgQOccvi3o/uWMaabSi6Fr2C9jiRfGP2UmNyujvfnO0EreCt0UCO7lb5P
E+/2gHSYq/OFwFOr9z2/nNErA4fYtkbziR753096DnqSpZG0ZX812usQb6t9Mq23CKrxcNOZfq9O
1jiGogr9+cmjWVvsUJMKs69OjPQK83qiduS2x6tW1B2SeYWQMdVvjlEh6ek/LScF9opxANpM2ye+
g1JCN3KG0PaYQ8uXzf9PM3IXo3nWPtOTD5VR6heJ9h+DmeerbgTkIZqYW+r/mGqQB761MLHsPeuA
gMxXUNddsntVKGZm4gOsHnKJsuYVl4RVnsOtN33o8BsJkztPR0R41qNIqkZa32ACuSkPWhwpNRgO
0Q/OtpchF4Twq/wNo6goHO5TC5HqL03kv4F/rb4EzDvfc7oYQnOsOGg3lbDqwO3EdRKMNX28AWAe
9AIeRJrc3XnXlEemPEPCz6zXZ7+it3yZJ55Ug4vug1pZxAOPjs5yBj3tKdBBqjU6vQIEFKsS9xkB
BbM4MSyaAdaC/ffWckRKGyQoodVhuPUK6Deh3d4d/XAwfYqJJAN76STch/zWbz1JkV13yaLqhP8k
avGCdh2MqcziqtRUwNTemf4V3kR5LHmuGwIai1VoMbyvRJ3JRiHWkDfGpWcLmndOgHkm8USDiQUc
GKapPwTo5wxybErXTNjb5aJXhnhv+G8WW9VqPJDucxZ0NCjW851VaBmQUUhsnPH2Xp73I+VIwu4y
iF4TjqIJKCnm9NVzQYqizqSiiZZzyuVuGnnXku8q+4R4LtzH082fHiIvc3Sz+61cWcMlo6XnEadp
B8GXmMvdAveev3XK33Mvsl6h56FAWx2ToOll3aMPlYyRPUYcrouXnEL+1w3j70j9/zq2ZESCSJ62
vcdZdXnM3B7nGe+Xm/g+IR79O4+p9f0I2QBBzagdIPoaWbt+T7VrmwReQnlGGkPbahqrVuTnWJWR
UPS2EzqcfFh0aIQWxapVLy6Zc8PKdoTxz7mo9WbcBbWJTscRRt90+cPmgrIKjdfuwVuCBqzkO3Kd
sr89EbZc0UQZaByE0DO+/kitsXP52bsWXEj/Kd5GbF8m0SJvqBPJbY2kgjwGnU/mtfAmmXE4moXW
CkbtPKDTYDAN8aH+FF9+cuL+T8pzcgufgxrVHAFEqqKpNJhC8PbCs//pgEXH++gl+BpbJhwXEwvn
2UclEpjFYJZWaFaFFABWOmnvhjBBPJG00EdxGxP1vdQXAihrHUU+MapsFpIZTmHUOF7uXh7VeVDm
5UV9eUTuaVQ23VaHbasxz9UFDnTTtNplj1a66qCPDFNa1YV6eryF/CukMlzN9MxRD+NOWapw3+2L
usjHCjR0rIYPWtKLYgrcN+xZClsXX6g7Y7g3dfBv7o1DxZvk3RiE+MFP5Htb3Yl/Nc8yu34ODN3Z
Aoa+wUWGsshvHhnxZyBhU37b1oyi1LwabcxKVAqrvPrd4qaTYGmM5jdwgQ03fBe2KumJXF3jhDrA
cw7y8rBGltFgrvPU5Q8S/sQNg4vUUa9bzQitdDz44rqDJbS0s0vGKJsqUxPPcdt5WoZC5ag4oBb2
gcS53vKQmd6y18hAH06vEl48PXTbOHJA2diItElHvC7JwycJeJf73L1+/hRCxavOoOj3A+rPtKMt
0MJGCAvfwCrwaBbiAR5Q2dwvfqyI5yWbiLUj/vikxnSnkGFCdZ/zmq0NP6WnBoq/kFJKmXs4o1LA
s6GxKvV+DinR32zYM3vAeuM/KNqF9EdgZh7ELrpJ+kdjpsaujHFQPBItHJKvR9byuuJOW2oES1G7
mw+El0zpB9nhBkvET4RlH3O8DKKjOsexR3+GPIFWI2rkZkEumvmUAicu9EeNcQNhlrW6buOhqtxk
jJOk0nWKNDP21kTN1rvPXmycIgla6Kh86jq3sI1VnBhUd6XV77saTVNnVfXQmga08p0p3YVbCpS4
39CCdMIQDUHkYJWvQTyTMulIRJeJnrMwX58UYORM5YMYaTwvc9FtHb8aClRbfsRy2ukixjfDB8VF
LSSv4LKdZBv/Wgb+zI7iD8GPnpwQJjM5e187mjCfmdUO+deKmO7KDeUBz6mAyLyEdXENAR1TYPEf
kfW1RqdEqUB8ce1aK3lesU+4KKMxVto5JOCcO9c4QCicvvOi/vXK8LfUl0f72p/P/4PiHKsxjodS
kI9j47YolY4gLvAt/gRckjEh4ubdyUo8dzEBX2djW4XmyB9TEjm/klheVjZerMF+QUP1S5X5rlqt
C3GXvhXXIIZyZNp7xPe1dtNBcYtcK51+j7QbNv3u7X2QRH/WceqxRsMOxrz7Aagt4ZvtmgUaU7TR
ORuPaViJK/J8AV/vMUkd4C8ulAcczANstd44T1Xyv2qEiGfA1dRVFZ/zWJu92IBoRJz1MqoSuSF4
brAqxkQod8W9Q/DGxUCNGZ2H6HMDF5aB+1cq8hDffqiylERYjRGJVusA6MY9ox98cvZ0XL0ozbC4
R8drSGQjrow7gHuT396JeaPG0rw8LHNistI0NE1s2CWKj++ZAX8frbPiYAGKHU10NvIXsj9f7t2F
jqD8sCRUM63GXXbBevxKMBmLdwj4rrcmidgPFQwUVnw/U7MGB9ye1EKxxBzjLxFApLGGj4aD/gHN
T86qlaIwMWUeydeyLxGGY0zpiqut4qwUTrAht8iNACxQsKnObnx8tmIqNleSpMjxrrhELqjzfAmt
hIauJfE0PMf75DlnyaHLhFdvb2LkuH9GwYPGyubqNK/tEiSPLFBP4RL8nkas9EKZvImMt8AymDh5
3bWCOlHeEpQxQ3AkRiNC+HnQOc8Y5qt7sWYkNsYBzueklGXVypmRXVT1Ri+21/+1Swr+lYJ3JTDq
PiGjnnLXtpo1eqznkFkCim3p09QlVWJE9TPYrjfYv4gGKPNRbE7peUhspK5U6vBnPvhXvcEBol8t
m3RvkBFjFLFb2Hg4/aIwO6HucC9Ay2koAH6Rr4NO2swOtIhvV9FrOSJgFB4ol+3Nx5rquzGGvNQ3
CADxEUaZdLhnOtpJR9pi1uFmsm0Uidv1MGN3SzhyWpd9VsXFJglxW8DVQDZmEJZ6Ldvwf9HTdyVR
BTI18pV+6JYi6x9n14K56LMM4+VnxS1j7IiU+B3IVTPv2c82I7yckKUlp5NMZTnelcYc++OUsWBC
zb2iEqYl8oljeZNiwU6jf4MzMBhxQai+7wJkTH6jsuXxxf7aVlufB0UidFxVNk4hjXtTZqxZ07/T
4LaTZJt8q/VJDULNwBQQgRqa9Vz6oR9yVGkTu2SZElS/7KDqai11EOZ7dP7rFbL1NQ9fI0rWPTg6
j13UELZ5Tm4IeB5N/QmgwLpaU66UYJowv0/SL59sukjdcDYI12ZJ+dC78XyrtB48u1khdXD/61/d
0RQBV23arNran2Mwc9PvrfYlSx4H3vLrR9LjAKOeKO/lw9drcIga2ayoYlldcHwEA0+DasvLKjrp
SKz6O+f8fy8zr4IBpdX8/KIWL/C3QhTnVwZzg6q0aKqXmQuad2riOiOobOQSLHn6lx5X3dgWm164
nqtUgedtke1YIM3CZ3+8vzG6FT3iPRbGFbF8zs5P3lNTEw/NVrCVg6RaXf33bms9X2X0ByLGupmq
BROidN+n1HpNymcahFcR4jF59Mdtc7JYImtDi88CSdMMrRidz/KkO+ap2aFe1SXj1sATu6uONXYB
HP7H+bi+3j/TEMzN1t620jAJc2FIxjnfs1IoMA0RyukCd7lyV9PjQDTy2um46bs+Lj+v2YO1Eqgn
HppcE6CDXrPxeska17PW03+Fkxk+yhNKikQ4MqvcTAuF2YduoWStmx+jOWbIELlCAeg1nmPvpRIT
SxeeyQ2CsBMN84lZAlDjZ2hDW8BWNqeLdTnSAa0hKzoGU88WTpIBBcYOGvQpW4lFqukWl2B4mVzf
CyouMTu9IQlvMc7pG0l+pOuWGuggpUnpoOD0aUIkK8vrKirX3VIcvhmq09BFJ/v+AL5X2suU2S2N
sIGl7a6uDNAqgliUOIp62RSGajSHXUM7DlXkG7vNhm1a8EEyouufvecKjLC5I7pfzxQYcl7Fx/fm
AfdFNPBVLt/Z5SXuNzbbYWDtH1h23fe1iRpnGUvP3w6vY7Qn+cYdSjfGhjUCGAXz5egN4nGhBpW6
TeHow2Bnp68rOJuXGXF13+CID1W35eIrZQvq0KQ84oBHQwKDHOAjxexk0WNHVC6msmQfD32w/SLk
rAnXdgnBKyz+uiBJszhUwfW08nG0EUgfumyly4/tOxKIkUZibRV0p/knwb9BTAbbflV/DG6XJG+6
dKJBfbWmkW32ICl37BGzTHenNUTAsKcQ1fg+vNo/9q1nsnbgixtl/Vvxm/4rB8PNWHZzAqsbb8Zy
eI/mQAWd7E6i+FrslTrB8mJiazrOB37RhJ+sfC/m03YnFh2bSDCudQpM1vVzT+5eYpBm4TSalAGq
EGUbKuUSozylzZ5m935x/vXM7BTaXM6LK/8evuac357UVbjajAaqiaqDIbi/9+NJUMJPGpRB1t58
IchoqrBLOQr42JFY/E8ESfNQNaXHLGZivSOeXeKwQ3pb38Tlg2rL5iFfPBLjKcKJfUnxq4DEsaHU
mu225dbokLqdRkxZ2knIqv4GJkDGFFFmkT7XYDlFscieKblKCq59LUk6J6NYMt8/3F3kCzfGCtI8
U97OciLuy8fd2zONQohkcffUYMeQfEpqHmK+lgtQ3qyOShVMjP5AE7ZS3V+LCddeLtYtFxvLt/mL
BD9JXNG7lomQjpe+EY52pQsD3kJ1rWtgPWSokrE/igymMxtCDgz1M0n+newTHIQZouUWzGEwnQPD
nFYR3Df6PPw0D1z7iBoBN0zcNaNizAUk9/zos1p6j3ZENDdE9cVp7y3lBgpcQPB8llLqzXj5Oq7K
8R8BikVzVfBwLTdPbEPP4VGZydhADHnMUOyJhlp3ASCHoAQYiTSNi4P4uvH5gymbdszJsDwvuam3
CVbTknLDICL15E6QQ48pdg70q5MSV2RmulKSHPNjp2Zq8qXMo/f40exxVcwKtfj5TIA5fH6xdHlN
MgIIv456THs3mTXCRakiZ5jsVpszy/mTBPwv04I9RJd48qQ33O7mqhWWXo0JCZmd7X4PxnI8p3HN
UKuT4WQQKS+K6ePFqn3/uz+z2vuHJL820k2dSrJX1k0vtzxs3sl/pi7aRjp5ZRUfjjgJApAprrNn
X6nwY7WfWaDOO+RLnEUZDvJDwkgWKz01CXpZmvJeYXElphuiwP4TVlXzMEG5LzNfhVAaXkKZ/0ue
kEfflvcZi5R1+t0ncYQMGqOpO3uQ5ATaFiRlfd2LJx8r0krAl/mh+zaM/KbC48Ot86xSKXAmD4Dq
lfxRtUiDtGPmf/gYLK4wWy1k+/mvA6k4K76nhJYxqzHZlJ0VDQr6nUqHgFlkUR1xu4kFuX42A7q6
SMgqQ7AIH8/eW1WOYa/+doFE1j3bhDzxzs2nvZCmmdHi9kmiWqw+X77Y0By6vAixXVeDuJf0OAug
kH0lBKZ+66DLT+BUfxT4trSsiVYVeDpa6rYzBm1Lp+a/GB6hupsfOI1jZWlg2d1OLJ68q8+6voIp
hdJAxK6qekgB0jIfYTR2Lcqc4r0kbr8iKxDE6ykZmnajBVeJyrctUp+SK8acKqq9K6TI4yH37/hF
Wy5AI10WyGJsCDCQLMgF5fiSCy3Y/8WnTJH4JxAwpi1rZgsxeeTATBM5FOGl45mU4aRScM1XIiJ2
TQgAVF57fifvqnQIXglVhBmybL3DWBBbDF+iUfFPQXUfpJn5k1xJ77AopzCfrfZGeF+xzxACcp63
OfqYyM2r7qQ0/6vyjDU0J3B1B6I0O6BH4+mtzXdtE0L+agxXWdRAnjIB+mKS8z2JhqrjtkNa/vKX
pT7XPQc7l5VEw5kDS44TJFHfy9mvNwu836d2K8DTtQuPw+letUMljzJmVH0CasoStB1OtG7rv5tT
tS2lJQME2Yk6SWwUgP3qb+4wMjFBGddzkHDbkHqjOoIhmpKNTrOds1SRiSctMq9J1PPI/FToUb4q
HeJGd9BpLnne0d6oVXW85LBkTtQO+/NxiQPFeaPGZ7fcQVvp4NBC/kq5qHeLwR8nB8of52F3QOth
Jco1xDVwTILw6gu8YOrLnfQtJeCb0GEp+6mdqq+ufIYtikp7j87DvUXmZ1CXDGDcDA16QdmvcwQA
+1oyKdv/hknedpRAakYGQCtWqT1me1WAYq2Zsqcf3G+LBBjFLS8VU5bHOpl2gauyVuyE27ROWpYx
6eTIkb+H9XMmTHwuuGP1DBH6X1Cm39QeALIX4szCPe/c+7ZsQVbwiV9PUavk7ZJXBpyp+LZViWlW
f2KFaLENaqtiR05SVCcBLLAY/99xf+g9TPdkzVDqpn7SkxvcTalxZQnIBf7RpZBrNAU2BbMFJWPH
kKlyxkopG1iXrA/2YsrG2UkDLiuttMkMpVH9L4KuJqvStZBcPPK0HFHcAOQx7vp7gcE94COYOkAK
HJMmeuaLH3p7Ru16X93UEc/xBHX2cJ22fiCvj+S9Aeip9+VTPzJ//Sn7qaGwjZLM+5jkShn3+7Jw
1Q3I1zCD2qpGR9YSqHdILVyk1OYQk9IC/jnoXV2+rCNdeRZ8T71+cW1KaCWcUKS3IdWooo30z7cI
A32ZTMIrnTk8dVtb8iOaqadi+yQPlEr3uzFCHBYiAFapxRJzVjCaVLUCOoqD6mHLawtH3SSmwsN7
ZTHqXPQStBywDWGUj+MnVSknLlRRVxcpXrVeI2GEfXfAS9ezp+uMHzyk2eN5mMA4uXjMECveCpmw
gKxQB3qnn7uSg1SOUyZPR2qWg8G/iK4sZx/fYwOXE9xsn5oWHlrNwUH6QlVukhOFQ87O+UTbnaV/
78BieyUsHWQU13KQEQhMdWENsGeTL1HXLDvvH7Qno2mJYr3k/HA92xwzfPVhZV1XOBl3wrTXVnYc
Y3BVlgsc2bF5BvqT3bBf0c/GJ+SZ+FE4eh3jAxliwP+dZlzfQp0YhSf341g1zsJ0+M+nuO4UkG4x
EmT7PsitTiIG4dzg7syjFEIs58G8vPZo5SQ/cV6EBWLp0KAVSUil0ZDvMu6Ryyl8hBYjzw9jhGik
wpqFvvpOrBvbPA2j9mghsAYLI0bHHUH/oGRDDm3mNIAMfCtxZWMKZ5C2RNEkWu7i+F4SSIZ3Rh2U
1oE8pcORVCBKK/VTkOS+jQqIEDNS8SYvFnJYc5qhLnNLOjRlos0iOcDzYZjfepEt4fLcyCdXod1y
f/wqMqS5CzheSkHFNqEePhkxftX14TPKmQpJwXmUejvYJ/C1FDdHP5+nOLxXnBr/GtZ+TBdOrgzY
+5vK6tQkzmX+gzZrj0iIg3fuCx3N+WY5Zgi7cNNr/ja0Un8e3DOYCXGBMeY+LAtegkqeajLSBSeS
bSEOAg/u7Tk46sXjPiOQ/Qh/JCSPHAqYorCZwNjdYBGrEFgQVZoc/GFAHICLSUUzrA3zrqJtpRqH
nQ2xkmqAaMtdN0wQnDzDEpoluvXIRKJBg2Ess5YIOzsOOmkj6ALBmqq1hb6E5IERymVknrbHNJV+
ZQK31X/7Hw3ZZQPOt22UA5dGbcNJYoh+3le8ijhoBXlYiorBsu4mOFVCRP52xM6HGYWYhZQRfBE/
0/jJcbolsE+cHGyyXhly7awnMmh+NhU8QrY+Fom4i4K9wgz3E0cN7DqGFo4G8nmks8oT15hf2K3w
UR/L2m2JJfzIQ2/6nC2Nk6arKfDlerOZVFC5J0WQYm7rWLpRjuRxN65yXmFptK4QfALs6cqHIt0W
RMbRNqSs7ZaETU2kyo8f6B7f4dMkyt9Djv5RqbSdshr1SlZHdBdd3g8LRJwVDM6beLTpviYmYbh+
hgtcuq4jti0bSUVChA+jLdY/yPdtov4P4tvGOx6J08YMGc2Z7gVS/5o/oC/WEWihTtSBPX7LU113
SGAr7yL+y6oEFTdxpu+Eb2Qo9sn+PConJn2AA+TkUWhRcw6R4klwPnOOtD2GK0Qo3D3YQmQvjZVb
6D8NHRb8CanmDYFA0FLlxWJGByeGYWfsKH38ptyG7+vGm7mFIAu5cnEwq49izENtd5GD+ExZkzeB
392CKd/iJ+Pefuptd6yzkQVGR8zHtRgGDf3o5SwbCsVLlHaCji2yB0aMbsWmXpAnNUfUIDlKZ6Jg
cMxReWDGMdmcXlFT+lZ1Yrub6PJ/vp9V7vUnVg0rCIdM9YM3xfIaL5xzpCRD3KYmRMgm3kdCCecz
wkCZj2CbMw7Q/TjE7GcVpU/FxkjRQGALku3+gI+KZvE+Zf0heDJruDK3WjqAxvuz+eO2HnNfai4J
TQxzqZbfB1dxGc7+1oufnlb0ASBrxfT0vKwCeph2MXgDmL8DslXCUJHWJmJzhCVfJn5/iG8Ug9G+
AhStB0xxi3hjUD26ZYCnCtsmGjjTe7oNOb4nQYUtD1Uxi3Gdb5N07KwWRZIzjFo61cF1EGtf45Zc
sjbT22s0eihqCQZAbJBe9/1G8FUyrEjXTOygayxLJx5EH1v4pgBCI0o6/hjrFmhI//lBw7Vo9G7+
nVUApANLaojsdRG1X/ANF2kp6D/L3DZ2hJR5GhVHQDeiCKseKL6PnXaVMqz3SzDo+vCjkmxpf5wO
+jc4M5JBFZ2zZTZyDv/VJ9WVxsR/XcOQshRUfIsUoSoi7EayfrYeSnJiLzedNcKLcMbtIBKVseMd
0pJez7PY4qvEBMJZMP1dG6WeKW6KXkZziCxnEuSSa9+1FhoHXV2GALFesNK4ge4e3J8jr5yQsz9q
zZnufYf3VdQwYZZ548cjmFnx4k7buykvM48TyNaixQzxlF1c5B90uVrBtLuWrULOJ2QyTF0/N3O8
2NjZF71AwxigHTxVbwKxY57QehmCCS9ibCJVYRVe+290i/rRtJx43F0j8acThby7PQumKwfm8tV5
A9AP1xmX4OBcROJ1npzNdAqkw6urvjjPragvfiBDvSXS9kkQ+51DmLyJSYyVdaJNHjShPk4JsuXV
kxd3qQFk3FiZJ9AlTF5tdsCyVxJasfELYOGaApeQsyV/5qryFHgbmLrkOa4A+YDJQILfomhvSxqF
4ZylNMH3ZY7AO/DxpPALL/mxbefDJNnAUluhhef1xHLo/R4darPLTKgmWJRQfDDko76VCu5orR4z
Lu2mUErz+ENpZedTb8ElCsGygLdtsw2WiFR95GE6BJMlZq959AXTdILlOSh/VTnCAv4rCEdwCX9Z
zO2RAgBUtzJeVvRYW7RfamMUpE42hvoljnHv4SsI9Eatq7lKWoGhT0qY2itZWHzzyewRoPsChr5t
WAukthCKEtvl8S9b2FvdJ0KbWGtkfTuMBq9JnsrlNg4V+AqOc7ot3F9eRvikxZEWQqfHgCP2WhX/
3xxaduYZEs+qGBSkCvxSEv/o2CgjuC1TlvM8msHBbopIjq/R1+tnxo/Ogs5z9Y8YiZwPpes8kHAz
YEpZ1TYw2kfyNM21dYiUTiVMvIBP9ZmmhigIlu/hZD8pup0yngyDCVO/AbFYAjuD8JRUn9ornd6b
zc2EUQhRnBoiWBlvYuqNOmfiXxEgPzoTJNu022qZOaZD54cKDRufjcM45HK+CWmu7Lh8dKkJ8a2w
lMdx/D7sQaKeJwVlvcxx3WhFjtX9aJknXiBzCVRcraFS5es0Y6eR9YXcG9id3fzh/GhZ6zne0B1e
eELR1ScEu/bNuLFhyHHMgEbm3MvcVKkDOzXzYYzwzNToZ58rlGXW4hfLaNJPq1CcQUUhlestWvtV
wH6oW16gdQNjVsmfwWL85uZUsqSFsONrvXcJRIA3/YXRVCyhel1xwk4gpPc/bAkpkBLzCDsCi9Is
i2G8bP7hPHvUQd36cJad39uczw62xB4kH6Z8h0x8wDk4wbmcn7Xo9NItIdBI3uR4MplSCd7Gwgo0
eNvdqIbFY+pJ/XExMHl2zEGL+O6xxaMR5UmPz0mes0zMfbeEDiz5Ql1B5gETUnsqBdnWchtVK8tu
Cim+dHx5PqdztKgV+ZajUyp0ZjvY+NGfWZ+wEHtHnwBRveQs+EZ7J2G6rRrMFSq7lVfWMOuB54DC
YPz9F0NStRG0gN9NUkEfJsm1wbhrVVYupA829RmApJ4UZkaKuXHvh/orgTyrZGTrs2TbBx8AYKrt
Dr1t4mugMm/rYiF/4XVLxqXqKKZdMpJAYthc6cfzS/fFmQaVNiuivaArkrarPZp2oeTRddszK0zr
NZMjNChOP/ErpWGH6sUAG2omxkKDG5wUpaZmPBcIST7Yxz6Sokckz1BYmB+MS70OBbHU/Q9HYEez
9lBEeCj8SSiwIeXTpUb1nFscDoiat/7ysotQNILsHglroSrzq2BqjnIB/W1yJ39/oQUvmUtyM1dS
dfgJzeqVkoFjU/GTy55JnZOrDigJyuO+uhXRmeyNoLZ+QAycqfwkAYaDgXYOmsAjJd1HqSByuvVR
6LN0NHGKsgTcAOGn+SGioYAXfrRj42eVaatDlu1+JZPYEZhhx9ymIQ7gR0NlG/v6APhaZJ8idTwO
7SomKKD0jhJuPz0YLI317LVki01IMbQRgCquOJsbQXIBiDrOpEE+4yzxNkOEvd+X5sDJaRUFaey9
FEIML35US9EAlVWjvwr3Cx9PnjWatrH2m/vy0ESfnuH2XkAP10iBCOP1RrC76Jb5Mz+E3yb2m47h
OSzZGfAwmcLR+p3hDL8Z/X/ej3mFFqNDaAQviy4pI7oFPDc/Lg3oa44BsmXJxcd/fGRZkFhOMQ+P
Rz4V/X7H1xiSelkeCfCJKdp5XXe4hwv97mcGT4fZDpGt6Tug+O61OioFiMnCDVk0m1g8FTwgrTUC
fDas1w9MWMv7govD0bhTkV3zG5L68YOB1v9nT5/V/VPNEUo3VVFCdIOQMmHxh2AI1EV4F1hqFboY
QxowruPgass1f+KDQ9XEZhjn/cRzI1VGNaXpxmAhQIWIncm/qoULIm/Y4e149Cp9VlTXg2cBxiJI
lplgVbustJugBjZpJEpqS61v54PXjNyucWWu0yW03bM3AK/8KC+XETrKDEees54K7gIX9fpLNGfG
aGAORDxL8CdIe4D0uCOJB/+0QyP0tY1yv0+pPMt6GsJu+PPvCRcZY0wGMpbERftsPwlc6OQqSotJ
m7niKYF9xQZwxHwE0iR3iQLuoHcwvB3n998HK6WMOJSlK/GQ/1z6giQmdkyoHz7eB9sIl7FAXvoc
hUsmbR6xyu/QvoI9damaDQGCEH38csbyS1pSwDXS2DhsxPgBMcPnmkopVz30bWgi5UqkQb6dbcGz
MzSQZa6G/Myxaj2tPvTGilW1LQkp0TW7xT45V9Uz1CRivn9jpOtmoW0qwLy5c59Kvi8HRGpNEYyI
fueawEox7Z6T/gTxiQYbRdgsjpxZVrAhOiW6lJ0222hXvLh3VoDNg141bY4IJHXN8mO7CWQEMXLG
20FwznRuklETEcmxd3/TzoUbW+xUoX6T9IUqVhbupEIpu8yXZdT1HJTRuAAlDxKcq604KSpzA4FM
nXTIFFfU5KxK92oV3dTvWD+yFXdb315I5+8pbrFKUnZdY3tVkNTWcUUOJVEGpzYYOogsxhAmke0H
JN+ppn5J0hScis6LBW55MyWMpTndV4KvVHJHuQi1SVuAtypjlhx9OWKwv0KIFPDz98/I2bSk7vtc
mhBAouJ+PRnkLDpoWLKj/7rCSyLTrTnhntqLXW+haEWL+eM+wZpxsEPO5+XXRz4LA4IXE1u1GCJE
uO0fEk3k2pVAdCpnjXfzZsZ048ywmWLQ2wnkBnQ6Vh5ZdjC9uouBm68sXOPXWPalBgV/+1SP9j9e
uKiPhklycv/7ij02tCvyZxHPPp3PDKKxBD2bctt2lBzVw02Eqpwj6buTNAZBEekxId+4cHXdxiAf
gY3/A5lrHt7uwdtyPHA4xajVo+Ob+scmOgGvenT7fon5m1OtvMls9Gs6+vKh2QOyoMJ9lRJZS/BQ
/RNTo8Muvk0t2rvYQHLUNP7znyIUB77S0U+VBoVUJrUeFCmqMAz+oUX3h8qTaDs5XH1GPavYsuMc
c2JtCHGd8C8UQq3zpRtWqnJgr8xnupjroJqlgnnxIz8WpE+QK7EAeLfnDsUftmPnltd4oMwU85wu
GP+TXzNi4O5EDriV8CALJNb+8vu/bTIYaDIPXHwCTvaMAZGOkaFDmuhmCclgN8oX45ocmuwKlHM8
0zZgfOaUfCJyTislLlOQ+5D83l5gfo7JN1+rio5ViuWEPEfCwyLV9UcAzKwJc3ZvPqYTqC9dsVEr
bQfxCiCW3zp0NqZMGrX6TEAbCJqYubBcghAf61jaIC8l07PYSeHNGKxNHVtoajAXCA9H5Nf0XUTe
QHBpZaIkoa7fSGB3c9zhtBMXwMmpCZLTYSjPNbIZxcKUR0bK2COYt5djHc/wf8IHTKAYB5vBZJGR
rOJvlgMnBjqO+iRolvWWTb/OlKXmDoiulszQD0LCqQrWjlrg/qNqVOf26oROevSSCnvhcpM3hqlA
0KMBh1EqEVCDyvPw6M8byO4sD//oUZCA6rW0B/dkkc/UIM2iVs28b/PmgzYbtGmK7IC6brCisyuc
EkPlBjUzY0F4gVDP8QdMEJIwu86WoCYk/iJ8h3LOzXov/IjqpuH6nA5opkL694nYteYxu40HkoPz
LUA2iClySX4cg9PilPnGp2DoyeCc6drHTnqWqAH/aO+lFJAZRZEDyn647SQeHV+6SdkPIRpXw3lu
NYkeHpvrhDPbzB7ofEq/Yt1PNR+9t+56wLWxTzYXoN0+BfKSIwD9qAd2t3JfYtHvXZKL2P0HWNwG
a+PE8mXKf4hyG960KH3CPzOVncFsOS1W1uP4Xg6PECN2Tdt89QSNoQ1UR2s/sbSPnuW4Df8CN13t
6LixSvE/Tm/JMS0zxdI/CXn/2LOqCdnDCSCqXEepTVs5zBvfbowgKOKFu0Y/f0M7njA1dgDuQMGY
7WEmX2ksdHzxtwQnBSbs+4hDO31moGUYPkPWarK0XPoBoRAJXhI7+W/YfUJ4TM0/0btThynEzFuL
eHSphNVKBZUpcihSJk+FKgzbM0iLA8NgrKqifb5M9N6k6M3VfmXdcFyPGRSvtxZcwNjhcVgEsUJW
a+dOkqttAWZ1DyZvabU38A9jTAWxEO6OZP/vQUYpGB5Qfwrc4/kDfVYhXzKwlJKZsE7+lmWiBrOf
mT5urwSttoA8mgzg2/2p0mroM6/NgbJAkGg+WqxMHJpUSoa+7vNUmLCzWooHxpWJYsGZxKL7P8xm
xwjmd9e0RmPvpZE1TN06fsDGkqH3/IbpMZuEhvp9k61Hw0dE2gRc5uiSBtuAsqswbMT5x83vthnz
lj9Wog1rh+gOhyXrYzsF5wjeOrXhorZDh5RXctJ6iRXO1OvlYN8ozK2OhcmKlvJvJyxbh/Qe1nDV
xKrkWiSBeCrdDIe670qOTkOQ2667WVR2TnbJQXUuI/3NAqL1gn51K4OkHsrL5KnwFzAku48spnjo
KtgJsW1j35H9dWVA/E5zUjMO83CzGTQShnPaFOjbmjLJZTxGQsT6+JbRoTtG49AQN1mJ6ahD8ghu
XGr0sUj6JbuLgW9BKTpuKgvpvlSKtoN0GYQUW+lSgn/hOFcfKUcPHdq/h+ufbXYtWtqIQB/1KlOm
L98/y9YGA8M4wl3SZemtfgwga2/MLZ1kBIgMceMLgpP//Cm2ZWAt4yZvhPI18Q6jAwQ0EQJeUUgi
sxW0Bk30em1LvnEkehUii9yNa7vD1/uTu4wHpyIVlSAmE8wx2nMCskSX3MLBxbFTE5bi50KUfarH
vF/O9YQvVtUTtIkO89ughSRv5rK2FxqMyFJO3eszknA3F++RHNVQ5k0bn1MYjgvB95lBSADpobZL
E5JxGFnl27pqK5sK4RTsuibA2ibAG9B2EIczoBUByi/P2lSae3y9jxizH6mNzcR8Rv/5dTct+YK2
6/z1xbbI32avuaiXhDoB95+Bb6Z2Xc/NWm6oYaqOteSw+wl/TYmb+9TQZKa8Ed+qHFh40CAE0WZd
gE9d06kbDmoN5FLWt+HPqVZXRzRJgGO/AKMlBNEzdmJwCF6ctkjyQCPeJWboi9vRKCvT0sqzfuDE
xrZH+UOoQmWj6s7TLAE2KO6wQrQ+P1J9skjBUwTNjoHYwpQuy22RLSBaAYWSZipY4iX5JV6uP7wc
OxhvVCLJfJqCosKO8v3gDwcOnVrQf0ni/zjQ7i4ePDGNMNTk7WoshWyHbCaIwLZEeVftxki2Aa03
b9xUGcRPWJq0dZBOKvhP+hHbk4GrsZGdz0ex1W3pAek+HLiGwAygJpc4NsZ8ihS+E/SujD52zFkG
+NGVyOMgHJPPjNSC+UU/kOOot8Eo5FaSQ4WvToujaKCRsoPwCoSWjOv5YQGu75F5qf+rYs6Sp1ML
dYhhdDzrCVNnsEDWojznZIWK2MxBDSlSj+GZmKd14dRx9HczMPsLwUFkbIV3T+Newp2EzkiPBwvp
BZA8S24RJKrttZh+3ZDjtpELjqJvJrajmPjjxhkd5sURCEGmQGxfrPzz0+DZlVS5c9vGHs81Lfdk
5GsAMZw6eVPAtyQq4UjsacazMApMw3jTk9Vs77mRtBEutXQiEHapXwu20YyJEOrgzlNq6lL3UKcC
atRvzUTwVjfPU2IDkle1PQK9ScRNAtFWg2+jasISckGwK8Rm3bWBnlkvIvBDX0p/AdbHTwRIj8ak
bN50ywLBA9LDMHUU1B0g8NQYhBN8CgzNnSn1QGfSh78w7X//byaJObLD1AWee+ML/i/+ZCsVKtiU
CWK4zbxWgdzvxzcDcBISh9I0q/z5eWuEiVkhXw02/HCcGPHHx9l5LUuxarYSa/N7jdgd/4DAYoGg
eTMZV4gzLtG8LVHEJZwvCWL9sEykNMpDv2sE0lN62ukXZyBIS+TyEEntasESOtxFjNzARXTESHKw
QiNlwVLDjml6NgTMIMY3vBTr6eEhHR5/4husj6FfWideGXr/B8KjKE0WKVXzWh3fXdIneAO5qWxs
Ow5ucNX/9DQtqRhSiP4JAfwTXS60cM9AkTHeF0unNo5qlnhfmw1yeTfySm7DDBCmSYGcuSZBdB0j
HnrfrN07bg0CpiwGLKUpVqLHRAcPARMcq6ZzfLUpezzGjkidm0jnJ9uK/y3a7JTz2qn5J0FvHbUP
CUXJ3UerwSw9vqOrd4CpjIzghFwyoXLZ72V5SHJpUNPsSCBD+o35TIYyo2B/Dy8T5i3aWDf2HI8m
QgK7J3GijcwAXquXMNFQAUv8pi5SRjfPLbAkArRHTifmfIIU7ETBFgdxJ1Ml7UDt9A/EBS7qThrz
Njxku4W4MSWTMFkIbL28ZG+EnnCboFhPfndvuwHpf0ANGhpgd/YWND3ddRSjdgK4/tq2rX9gOQXx
2n2FsBen05QQWWUgbCpOycWmj8P/OIS41KBwdT9F2ed88meyPFPDhOcCKsvPMVk+cGuVj2/4QTZr
pm3ZyZkBoFASr/t28YUEXzYpiYqcgC45MuF3tWw5bVhiQ/xcjkdPY4eN70SOWMtrNkwxo2vgSJhb
HwUzhxPdMEFdYklPtz5eRK/vsLPwfCDWkAlYEqY3xEkemsche6EdXJtrfxdgRV2n6cVpd6Xtbc/X
/KYsPaPsM0kV115QOS5dB9G0JvLAvJ5WxsjCOsLjXA8GH3iuTI2qBpC4yA9APguGLLyzGoApBpQ+
QnnV0G7Rqs4xrSJYAnHLJvKkeX+ZojpHPWqfkh7Y0fYthlvcpRZnLOuca4Fju8H/paUm7hlYyNIr
y40EV/OHt2/KghXQL68+W2Um0Q+eP+yc/XeO3JZUOXf9J8XqCLszydY402kyJQp6t9VAwp1VQx/p
yWyE9fub+K2jhN2b/J7MllnNoFeNVZJtJKUsyex5rqrBNO3yvSPv3iwmT+BUHvXLOsgWBbpZ3vAN
PBb2i1mt8ni+S2n0Rc9fCLZvUnLVgTIdKyBJ6Q8NGHq/7U9SdEes5XW0SnFZKTJIDhHCtU4GiKX1
I71TXb8z7WeTU9EIGnLvw8pe6wLjQJyBMqzcYHqyFLPhS3XWAqslzJyLK3gcc94daXR6eDrhqJ7Z
KDa2IBy0gQXTpJ4ehJVGj/1qupMHvJ3m+DBQjwa6DjodLFue3THG0Z57tXFZHiDjpLQHPNYgkdLh
6OuefF6OUz4KWolSgXbqHX/HcPdNSrQZ8EaFkgx+2CZK52C2brK+UZauUlR9tjWrHDrXGN/kpCjv
naec/0ROJm4J17tmdkK6AqpGP+DtU1w3l5J6EjabRFM0PIOzANmgU0ASMjCY0V00m51f1l4+lMbF
pJBUGdSOBZsez8eZ0VzagU64jXbb/5vZVeAMwl3l0FHP7+wAyrT7YH+BQZy6jAEVCzM0gF5bAZpi
V6DrelqM+Y3RTaJhBnZyHzcrZbmIuWoc26mcuQD6+pQSKhCUaHNaRUBAdmzv5gvBPiKf7hRYlbVT
Zk5SjfH1R4mR8zBaxLoAMNMIRHgZWMkrjGaqmEib0eT09sAkM1ZisIvkCo2ZPjfWEsgH8rFZFw/z
sd2W+fEHMMcJhTYpqIt1/7OX+OZ9o/7JSKcrMZiPt1RwHbJlkr5L8mRqQzPYC9ggmrsrhIBhHK7I
Eoju7qB8ZLvQMb0vUMGBYiEo0EgWM9+bepB/X4miSjdskhoP3MvNBa54BchIg3lBrCjGnydgNxme
uiJ292lhwBOKRP6mkgDDP5UQi/11vsKs/o939z/59sHd+A8o5uK0CT5azn8G/vT8qLRBtA+PYwGL
h5sUJ0KgdrudJZ1fDNpMhGvFOuLR7B3yHR8bg+IFaY9xJWCh+Qmb9rluq+YxzgtpfXydaBkR4Gdv
tGLfeYxo0Hcek2E4SRcGZBV/b0p3PxvVsA9A18cNYNJmJyzNCVSpaHavbx3OA7OL6XeR3ChrXw+O
AjB6qY63JogAvqx6wYjXS38UDBCJ4f2QeSqaT6FlOk20pnrul6odxUriYJvS8sdlModWf+AI9oEk
9Nybq0RHBvMs6W+qZ7XJAi/M3foMQ2tUm9svJfXvGvB71c6cwV+WtDK+mtjcZXAdA4MuhMN8DGBk
yyYLEMgHH4HIYeGzA5czy7QxiIKz16nBnoiR4pexxMt1FDnnX2ojeKzeqXipf13VkcLBtgVW+3j6
ZmRae1JUCxCyN0vPpoPABaREUFq4MY6fRhLcIzVAtjbW+/T77VDs/eUZcK6YvTIkEvAN+8Y/Jzgv
TK37A7EiqRAd5oFN59cZVO6GdQCpnCGzSWkOVEYPH9E/aMTvnXGApzvusCw2XSiqQceCrTFG3jnm
gXU7IkiyHUUaDBZrGPs9LUvA2C64bMcNti8JtM/CqirTOEUGShZBALfIRKiEmG038MB0V4BB5DIv
7wgz2gyxVQf2+03JYkw78vC9uVdFtaixnFJPMR5t5k1fglhFiDMJ4Xc1SdZr/EBflJdMAtdlNgn7
PTiCSVxNq/pnommXMpsD9KSeNRVnz/ulggZXX6YaAsGnkgNE8D2Jbo86bxlEvTl2sgSuRhYhoeIs
+VaO/J8XpapL16/FzAto/POSX9QnRCqiiAYTfCHoXyy7NTmG2p/MWNLlL3zLbDf5aboGeTpPg2pV
DdjQEJrBQk2rhQWtPYaKzf7fGppNV9AOgCahz4NJwSu6CUmDz3UyD1sBjwVYxBp9qvacPvd+CXQ4
Y6b4DNUrtRmg/zvtFLosB3VvDcmr52vN0kQqXZ742jxE91fe4uqkJ0L8kwwFlyqikWUaVs3ESrDe
x01FaLetJjZjMC1wqB3DbsKuubuTO2QZODJ3sxtztsrMggm/3NKtq7nAMosTp+hVUycMfTXn5jID
tZ4L6PAZoQw1Vh/yIytKlcXI6WD8vzLldPK0NbtsMaOL5yuwlhZAOd6pF5IGwX+K/dhA4zATw1UC
2oDcCg2Pg2FMqrAo1HgV0WZTyRzR51kkvjMoiAX6yoz4VwTE2Foyl2kEIj9kgTWVkqnbRcGfzroO
uBVKeRHON34TeMzYSpg277fH3fRu5tUJBtSE5iYwxbFzXtuPn07RTxo6kdyT/guwC2sAprDSNGXL
1uWtCBlAACWQUGSD0YNwBrIKEAVx40rdND4yjWH8yNtyXfkQ54n5ecAsLyXkbBgtHqe3G684dRm7
cLE3r+2KRKRy1lnFlxDY4k90z3didLDmjqglulx1PUMEUFGT0ibmyq3kHehzK5dSeZ3YBMgfQtff
1RZm6kwq9mh5h8oYrrnbx7QuA7L7HVyE0UffAFOJzdQzOL2TGzs28GtAIxhFadXvn8MF14XICrhu
QHSxjp7LdSciVZKOCNuWfuSrP1q8JAzhQtwet4+eG1r+Mz41yJdafL6X+OKD+PW5j3nS7LlcGXBM
KcCRK7XApRy+yjxVEkxL+n0JEPOuclIhVnQYZEIPdHVa7QDtqyjV/W7gnu1bVWlq/sLJsi5iMflU
nQKj1ivkUgeMdRhojbMRsUYzYrLYApbb+j+xSVTm6zkzPvOZ2qjDfwDQWvCf71R3nXWBakz6pCQP
Io2t0mQzghl4Bv1MDP+l+kTXkYN4I7k7Sbn+ekCr482EYdD+Clw2vfs5JjA0GtjsLZH29zMDZ6hu
iAI0NOzjNo709NEmKFPZ8k7+TKI3TGnvW4l3YozDqvLOMPek7lxADVECknT6D/ZZ9DHmzGS55h2a
u6sSQDPHok5FnWyRnZC7nmeSt3HKrgpYgzzQJGyYnELByv+9Hg0odWUkVWouQj0lEdtak2TC/eqo
zON5nkElBkY7hvAPIKp94vgywbcvlTrF9J/at5zCZewyqOHrl4UlqspeMVegFmqpqz6vHUkR2qhh
P010++n/hhSxRQXr820f4uXmqysFiVL/Swpp9mNFRO3BXWcyNJEdRCuMVPyH5BE0KZBDKpztttGs
/XbhCHY+kdn0rxyoEKMatRnrVf0ad/BqUK56i2D/mzEehWEVNwwA4XUXLdI1vUDst+Dt7hidKa1+
vJ/EkPc1o+xbDLnGhEL9kg+wAIp8uHddD/33xBSO0g28ghxOjGPnNW7s2U7dYNebxXeortY6SV3D
xWh25/ikPw2sfAOXHAlILl7l+4LNjdoBKLAouqpD1yBRd17LTNpndGK8FMzUAR4ZhQsbBOEaeGkD
Tap7kEHp1Ww1P9fkFu3ESWF0bDGP3ZJVyqkfZ0lZeaoLL6YWaSKeAxuvejDjtEHs+KBCKQ0Da0g6
JaV2hDkkpkVb90NQphSekigKb8Jl8LX1MyxLQJYAbQXpnVqbeiZO/WiMEHGGjmrZkTjQ3uIZEp3v
HiZMPmZHwBxPUdgeXGiQHN8JypeX+uy8QKYH+sYWrcph/Wdcqm4kJnHtSWVi4G13ifaoFxc/YS7N
Rhl+GF0PHsJoUnSvzFPLYoueEEDks+KpL22A8vHXECuC2uZboTkpVvGJjce23klRSfK8gsW2RsbC
F55EDUEJcpneZdfV1UTY/K9uiW5IxnOaj/+E9YHB5iGKoz5v2iHNDL2SeYdzM7+GNPUdIzSE4CSf
0FTZN/y7HicZ4B0p+o4WTdnfjj7r57q04K9ga1WJ8AqTGX6JeR5xAEVZrHDpFgaR0qtwFAPRO8Hk
4L0tGAPzqjeVfi0PBh3o6P7zod4gR7UCHziFfDAUrXEKbgEsA1mGRX3BWHUYCmVWarOPBRTqdgLS
lU46bnE28d8FkPiNQ1oNJNHoOvnH/U+9DEFiZ4odxjIdaaPpOae5YjMp2PyHtBjkhfDgVFVp1qak
EnJrKMzlSq3WoD80yslhv/A3ZxpnJBxRC/cmnMGEd//4bYVWU3NbAbMV9UyL77KvzBMKxX5LbIRQ
JrP2mUSGRxoHuxApUPp6oR+7kiFWoXPsK5Ii5UTIn/A9OVPKOjgqhkpv0osQzrrONF7hroe/K2Og
xdeMWjbhHimoLpltDg3NIUNqlf414At+hhD/66QciYFyKzRnMu4mcpVxcYkckn+UQyTmtCDovUaW
RAHSuKgPoGDd4c8xvljsmD7Y396gpOwHry0S2jWv0jMHw0MiSBjzQVrRoJaLQEBZebtxQkU6iqRO
eb8JS5ZhF/Kr2egWFWBeiDXHUJcUwsQjyGOLWedh5+q27KizZNHb1wuOt3xd1l7yud//saKkFBZl
B02Scday8vL4x4S+ZO29fH0Z+F4PcLlty8bvlvQ83iE4HSxeD3vjPkxdVX3jcl3iW3VVSkARAX0c
xLBOq4HesXLC1c8vh223bjQilGwltGSiWgN/mg0zu5K0nRfBbmg4AhJVaVumFFe4Cfchk2C6KWYy
e0sv/9tkMSupR5CqzGrlfGdjw3IjpmR2/B+iBJmQxa3OqODFgpUgsXUcTjppkNUd1Z6JJXI7TZrW
KmyUrm0HnQTu2IMaEccliuvZ6ODoAIiv7VVklE+ROOXtw8zhvveQJHXo+4YP0QchqIN5VW6DnAIv
21H3eSWCwYyrpFwoTGRKTDZHw+OwVuSr5bxzYGWHaVUkIiC5xHCdmjn9Aty/cQlCIvZU+yuVg5l3
RyfJcGNqh0TFPeOPCgBcB5CSQSW+MTzvpQnRKlhKnSlo19q0KWIYNpG0PuA0lAnvVScP2cQti4y9
vbCzdXvJaJjXUknk9Yp43uVYwNWdPFHy3ErsYSJE6K06LG83VP4uyR6c9jRpGFvcPK5gqHYPrqZb
FCkn+Un/KKMiHMpfsl7qFYuYpPMHNBA/yiuBaqikFuzJoQ67EHs2hdH/wvW8gHH2DMJFQcInkz8J
uMl4dLFNL5RJLOrUdiZomYZWJ5aeUm6YogO/IoI9pIOJ4mZEl1L619OzsCE/07pCJEo9638zhWW5
cDKneqN8392Dlyci03XoZom91mY5aBAw5LiJ61XLfcLoFyf4sK7owGmUM/CVUJj6k/8vNPYPAT3z
aON5qv5RykiFVi11xmFH9xAuas7F41UKGEenoe1lFBWB0Ucv2FMBpMEP+TcmoE1dyOaafez6c//6
Tyyl6X5F/cX30DRK4plpf/lIDfVKU3loOLEPx28/B2HAPJfDfo11cU4gGjiUdqaMkbqNQ5hzeRTo
zGgIvMKeTSz7G/80zx6BtuADZLj/t0HJ/heeYBoMc7n6PMNZmjhr2CteudweEn6bTjBBTJ1qu5Yt
M5RVFqQhRpD4YrxCfh4QjfRlWOyKNjsDkeToh7TA+De+MoiD3q3BPqtUv33y6zj9BPLgC0/dJ2J7
6W0Zy2fOWcRakqGFqJPRwh2Tkd8sEuPD5pvuEsXcwxorqUr1jXnVM/eMBsbKVI/m0bAti7lBIXDh
g8jl84GXr4qm+j764KABf96Vm3DGE2SxpZ9L4LEZ7xJGOVQkVLFiW1VvImSyawRN+tOf/ObC9+8K
uTNW/lqoGh5r5FbiNGIh7bQN0cQMzBmH7Wr+AOGgyN0u+iIGULonkVwE/VrDmQDGfIvuDO/tEVDI
aBlkOMwSJMkeY+znBYnwnX4NOr6DMgJNQGe1NFM+AFSpHWjLWzmca9nH/NYnY/6YaPD8MzGdCGxk
fPvfGKpy0We89i5qYZZy7HfQp87+IDtkSzg+Bu/RJ1uudGMmGpgv6q+7ob3E9HvzmAvFI06I9I4f
UHH7WzBkZo10YbH+h36DUX+Pf5pM5GnKHnHl3g3ZvGsrjb/tXBoF3Gasyw/xy52hWgYw0XxF1tZR
Gr0ZB2a/XAAlZLq/FfMUVS7u1W0z31w4oiJb3Ci24mFqr6r/W/Da+ErDE+gc0U8OUaG3BuUeWTaL
EzFxkX5U4qGwZnGOOnJqV8sc+5KTAwsDRe5uJOasek+FcDsSgq3xANV+pIlK3f6opXBeTfDtuqhZ
QmGlVJ8H+zqA6SmCDvNIwqZqdn9enhK3dqmhSijvoeZU2ufQhtk5PKsJbdtnQIzG1Vq7E1GKyQmq
uQZY5surIFC4SrnNw/aq1Q6S703Y9hRIdTtgPsjAAf3LVSxXXHzwOzi+PZRrbXYYTnmt2u2kjVyA
fT9XiQBlayOeTAO9RaRaLEtjA2BR9wnVbTBEvcgC/Ot+sOEJAvhAWOOB7ftyLo5ADFG2AnYVXDsv
ifaz/dg8kaJMpi5i4FtiRE0kQXJmJ/7jduv8Pn4xmTm2CE3gmFpBxQ4OWaOFjXFDN0QxLDxh87oS
JQM2q09sKo18YQGM9bkfV9gTlBTb/fsyEruCr4TGcmxMilWwS8EYpF8PhAMxdRXSwTVYjaZMcCyR
CpoQEWGoi+oCF2AfoUYL1IO3laO3wwAOV49ylG3H1xhNR3321asSchJFF1fYXYxkN3qjoYZGCHcQ
9GbplC1AeqCUCp1eJTnX4r/JHy9h6oXvO8sYyVzu44XWYnrUZYvxtYOKNEudM3YdReyMQo9X2PwD
GJyROzhkuNYEjm9Xlin9PogBf8Ajj72fSMtn4f1+cP5er3kYyx/TYeLUJP4PsuLJtFY9y52nkF3X
GbXTggZynnIHit4T8SvE8+miLLHeZhTHuol3wwtjCs2CR3bbx77LntMwRFDNpcnojMHO6Ub5ZrDn
WuzquWnbxR7dCbKtGhXk/15fyQGj2uwrCaYTFE0EPOHeB85BVepOn7RxcZLtsgNzZxcwe8qUQJCF
ANz/9mZCuYf1Yg3bk3ylvEeV7zFAp73taLau1UCz/PbIBXloIOxOyms6rR63sZ0992fhdOHJTl0B
8gsF7S0FHqXLZtVn+N/jBxjgNZx9i/gxUP3XSEdN86ZpvKR0v7GKqN/xCMn6qu6xdjW2r4KJlWFd
/rTD3Mv/KwMlDM4PTxB2s30zWG9C+uP0yhr9OXDNJa0X0NqKaU1x4gU9q1DTkDp86qF0N/mVJeWY
k7I9lz+lErlD/Jsq/oi83e+vzzukeyjDq7LvaOgu2JoHv8BN2OwL8VMiP6Y2CnG74UT58NOlpMbZ
WaXSdd4QL1A4eYGhXJQ/FvG6EYVHptTBYq1+HBEyKHSHjEN7rEgGRCk8Ne1SALSWV77ELm6aDWcs
mzJzKNt7WhC80RyVtR4wn7SAG26dPglp1aVVbHfLf/VBc0f+pwQ+OKK4HCYMjRrd/Av+Zr0e4sT4
gRcRPrJXLK8coCchHjHboLEdHlmMggMdrtNa3H1haX355Ot4LmHo/oOq+G1L2E9tC869MCHryWdL
5tAE6VVLInL60o3isJO7JvbfDnHXWan1WRCTwbCndiP9zmL+AO7oA08iTKylj8aqdbLxEuaZqAvl
piafq/+UzWmJpYqZbwHzvygjwTcE/Fh03w08du7Gs/drnp1VAhQNU/09QnJ/zZ7fDQDvKhR+DMkB
JnFpsNCCZd91qOJ9OqSG/gvayLRexsm9JERTAO4Ee0rPdDNt0WZs0Pmo+FffR8OXPNyccx2gfmLN
n6WCc4D84Uo0+pEFXthYvCJ+6E7YF2WN9GCV74PQbZ7GRexXppizlKQFwPLHDKXMfwJAeBnotm5n
wciY2fmUOmIMEC8Aif5Ty1ZRhg3eJ2VUqkG3GBjPdIzD8XxDpXgUNh6iKguV/CItV0tCg4SYP6Pt
J5qfHPiUbVpibLUM1LvjS9MZDbC+HCw6Jcb6JKlzzGsflSmfGCoMrBdnF4mrZDIAh0AKAU63qC4Z
BHWkmW5ZZJ+yu1B9cw4ka8vyN5KYs4Vi3ksZ97tQGjcFHI53/8pyuPZPwhHXtZT3tP1ArLZ+NiKH
JNxfa5XVIUEq9vYXyW4pemL25LrdpHGBDMvOCDURgIrQ0s+zVux5YC/tWMG97uNtb2zoolS+qSXa
zkutxznmqdkK4qKQZJL04dHoA1ikCKeU6J0Q5pOezbg+PSP85P0KhOdbg11m+PoKdALvKHJtoLxx
YrDPtNBVwXmjCxDMQwaSpOlmJ4Hmaw7M7ht6ieak+l/V6CL+/W7bIkyJqpWEg95L0sAVRhvcUT28
sA0tmv09l/gLq/WSi1K8WadnPA6CQRi51rAGmbMCU8Psv5PKlHk9BfzfSFKh4yDMIuLVLjf8jf3h
GuT92eYpZkiHZ+v0GYCvsVYtRVKXWypgnjUo4enRm/6fPUtHEBneve4LdpgFANXFlbVh2VjrcTAj
1wM69QI7LYgo8+gbJ6BTLHfQRh4R2jz0huszQ80bpIU2qcKvJ7TaWJYeS3GehtsQpRXjwnHaSRYl
NstUDy923HTQEfMHmoUgPIvCqng3uwWon84d4gGorHwYh81tGEr7cU3qMQ05ETLImHfdrCAnDHqk
xD+/fiLsVjVDheYJHLTitpUNUwCRs8k/UKesLe+W4rm05zywlxBJs82VhQihhsyhA4mfrbD1qUQS
zlTefVz7N6Xs7zee9WC2rkhoDWz9YsTs9e86oKFiIRo3nuTh9M2l/g7CBJDSfBpt2nR03exmcP0N
DapHjb/ktil/GHJMqjBAvK3+oGRrTg/OC+3XXuYYs8kDoXgJn3eZ9RTt3fyhgPaf3iCE94PipPoi
SvSAzQ7mWM1AxuQNeDnswl4FYGOyd7mEGce0H4+pQF4KAfCWfgRWSaYroXEa8np3rlUCc5ZLL889
SUbJavBo3aRhw0VLPNrglZj63cknaEoUVF+5HCMomQJpblqZzkwABZwn+wfQhb/vzWMCtkN1w36v
dgFUL225sPKj7Kgf//6EOl2K5r1ZrzcNefBaWbJSybnt6S5wFioMSiMfRIEHWM3kwxPTRIytHksq
PMH4jL+YeDBKcPqtXChsUYdISMkO6na6l3fjWc3aiTWbpF2VUrkFvth72PFBqeF7ShwFjehobSN5
C/JY0LCVLa0RQJmPhG9pwNFMPgSJTWOyai5x/XdmxEbzpUKe7fu8iN9A62ihdrKXuzl7U2/0NbZU
p4oKTyNtLjF8uXAMef7X2oBHLc0dBK4OdEzWCzqjaKNwlUVe3BDBTXE4JqQXvs0kLqpGSx3rnpWg
WEeQgszXHZV1nOIEvrZiz5+gmUI4P7DjWfZagovFgiqP+l4ekBD+JvpQH3o16yvJoVH7ERySLOCO
tvcoONm7xiLItNPYa7fjBTs3iPjC2D/rv2doXviw22MpS6QqiCwV7Uosy818XQR0M+A//iAffg06
07zLZ9uGya5yG2n3XZ0vYrewoKw5/BZMZL+O5y8+CJlfJrBvPuOP6o2yEbAG7MalkbUlpxI8b3nt
qN2IsYyC0/40AmG8Qo9uqoieJmdHHStuPLVhzYlfgjAlvr2BWCSFiMbEv7ZWGArV9TWeJZdGQfpH
/ADvpIDOogPs+HQTvOWQKQVvWmkVF4MwVNXdQ/G5QSN024WOUAPtYmtF+IJ7VE1kDXTUhTqtdtEj
fUsDM5/mltXjDOnIpqejJiFmOTzP2mvA/4wzx2f0CvFIWKkPhIezeR6YkLWchPKX272rXjJ0eryU
Q+fPrvvLliUF/YWoAFPIwKlOvvnj5oPwCr/oGkWWJ6xGpmcD9pZi5jOZh4Oilg68kGDNuiTiJJQX
UNB095UZiQpbHJFvPJrm+mUoR6dK+cIUqarrfzscGzEWOgGQIl7OLh6Ozrqiqf6FCR1cOUxDXZqv
FCxZNw0txu8LnPHKPWSDH55zBtOGGwDM+zH3EcgA2XB45rl97owvSGoTCYLCTHJgpH3mNF8F0T/h
vCq3hoj6ATKBa9IKxMKOG22tjpP9+OZw0amYmqmmZ/yH24rS7TmV9s2GweqVsxX80gp1ThSEGhzx
2DqIfbNbVhIKXUd5EJwQTIq+1RUo3XT5URKuCW4ofevKH0YZIJTbVR9jXXmptF2K7xknd0IJOeUo
hto+Oyq6qIc4G46fbRUFB5As2hbN9yiVt6qmRlu0L90kYhowCob396Es3sPEhFo2hzYiVDw2BC+s
JEiPA5awwpIZyL4lv5JPnnrWzFFIbaQAm4ibVYdTMklqbcXtC2BUW6J2dzU0TWZkGn0NHHDeToDv
otD8ZON5yAbcOFxylL/7BmrB5Xf2rNmL+M3x3rYdLkfgIkTrYWbqen5KMf/1R9eVPrh4BYKnpQBk
twkteS2+6+J/H1o7d9ggL8WIl6Ol+ErdB1GB2iTUq2W4YENaoeLe3UkH5xpDrCiOMoK1UgWDgu7G
DINaRbj4GFyFX/39x2ubd/QkAipM2tvYmigso6Ky4el9Y2tFYPItppC0oq2IV64RT5p5+8AfnVVI
ZmGyHccQ6ZjavGw7h9cJKIa4LeimVGQCFUJh6gAHTP1ZptvsNm0rnywxVuLlmguX3SVCkZ9Y9ZnM
N0wr20LYf/fet/jFwsJOfhW1sSnBF8S7Grsrq6tFDKRp9+WR0dhkZkJdz57uz0wBuaR9oCb54G3i
95w2x/K/sJTytWCz+8XFv/MjVniwnQXn75lGgr7jGswYxgYgcIPjc8ErEd3Vts1k5kwMAiu1s4AN
PJbvsMyFCsL62A2VMXP+1DQXVo/GtnddpMSJkywBwm8nSoY4Q8OtLngx1ijzXaRX3Er1Ho/SMaKx
xOio9SmgSjydpWQA43aBbvjiKQKEekyXtCLlaLO/+F4BiN2BJ/hSeFBkNRcqrhG8YIqp0PRTuVWB
5p00UMU14XlNHU0X/kLhJCzuf0U8hBCCUymvN5ykicqUd8P5igR8WpewmnNsOhARqaINw1+UfWIf
byqD5QZoRgmS0KeY8BzRhyRPYwYJFxwBQ9VjC+xFnPwt/p22zmWrkk8vstvCQohQHqZo/bWSppF/
K8U6eMqK9qkBhqrit6EbrQ4J99hr+ZzK3UnYaMCc4FablqLeI0K3vURXi5qboTuqcVCX01WYnw8i
lUVubVn214p9i4bQBUWekg9WtcHLnq2HjFmlFnNPSTq2UWa08FCqzqiQ0s9QQ6ZEKdLCP0ONaaGk
KMBxGRQTa7gumI7OwxbI3Cic3vSdHudVxZJVsBCgfhFaXoX5LzKMVNui+VjWbeKFtYgQ4O2pu7pP
OPzhcbehVbZuzDvCOzsceklaLInDdDxPi0Z7vTmPVn27AYsmVsClgExxl3+2Sa7xTjqSi0NubbkM
P8jCO/giRE4L35Quw+s3yqzDcomcoTc2wtXLX6eg4+qMfeLZtpD0Ubbx+YzV+j7oKLG0+dY4yRNz
jEKJ25MA6xFqrQ9b9xo6QUnw0zy6qI+YA6nikqoA7wm54hay9OK3Z0Xp6drZ15WLMAdyVRlTj8pP
s7nlC5bu3xUveLqGylc9VwAXkes4raoc7sJXKDAP5YC3vm/EtZ8gE6IufDKrlDaa1DXCWqQAZiES
0v2wjhTz/POptaXwC/S1xoxqa0ZXrMh4PkBW0Y1+PA1yLhUxswzMci/u2pQ1e09mi7NaPB/p8IvL
tigD+7e7HpoB86atjGhB/WUGRcsWCxzuhWfQThDSfc7EvoerGPpx7a4a/R4j7INAe7aXhKUhd6Th
fg1wU0ofa6mXoNNG08ktBduwFn3O3turkRbNBVw1iA00YepON5DcaI+7wmN2+qTJOdlNrIbw2QNa
1tFLbc4eCbAmXpSBWWyblQ1FCbyfScu4vfyE0el/PpA59qk3nFkEySq/pFyfR1PdXFZSQVv3sYVA
y4EuQfhxISMa18OgrblQ8M537sPHXukAzh+vHz5F6l/nFD7geHvY/o5EIkJnfAYUSZvP8xwo7Vm8
7c8W8eZBLmm70mHUabFa5LdC8wQpwV9QeGmuOhr4ehhGasDZm+NncRhLpQhkqrArbZa6QristY5d
STW8Wn2NZRY1PfijV7EPh2C9DgSf/UUn0iNZZs8QB22BztK9M8uwBS6Fl061CNTxGKF0annf+yTF
yJI+H9PojPf2aX7a0tVQ8OINoAhivUmx/fzVDE6nOusD9FJyjc7mLgucDQDCQhgLFEsrdi0fSOty
8Y0RUGITQV4Fi71Mzf1TyFdVRz0GYxU+pQLbLbA8M52wer7fRl10NsHTSyqfBrN7ng4raz+ehgXj
yu8IjHU/pwvU1b9uBscZaQmvdRPUgCA9AzJth4IcV9Dcsg7n+KCVaCLYmS/yoQgtZFcLA/PHietq
FFUIZ4BxS7qu0SVra1rtVgTZySDVI3L2z1KMMA8Zl2O2QHwysD5eMww6cL/1MK3wua38D3m94vde
W84iylnw0qY136w/lIXKaHEhq/PceGamcINPwTXIZfX8337hZKkKA62oxW1nIQfbqF3RnW5eM3vs
WOIXf9H0e+dy/x2z1vrp/yZSWWokuqTzc0EQ2N5MLA3LwdwfFGGnditCeez+LAAtLpCKt6GVEL2h
aKFps4lmziaHoS6ZtX431gKqb23NyQQNtfzMTKli0GYWgneuTbT39vknFKrmaSTJ3Zs2jdnu5+Fa
g4PzdUGXcsbwgqsvgb2CThjc2MGnZ3e8ehpSW3q/+uu7GUoGUyCmfPxS7zy2EJemgtYldIJQbKf9
gjjUNObXwt0MGAwvGEDLkHydU0DiKYFpZ3gCW0bt/YYLN96O6lZgn5IX+8hlKkm1HTn4Bu8GaoQD
ID6/wTxdDlT24qgJc7tNWJ+z2WhxoM+PoFLCuN/ewFpSNM67AgLDhVnngeKZ0DLt7NVTsiGr4qP9
un1BxywYyFaoqRHLt/RIubaFJfz/QejOjOZRmbp3LUy0c1vtaEUrXw1T4qAbLNFeYzZwo7kTO/gR
37i7OUIN2nwO+dgxEQkioLsQamsjsvoTrizuZIzTaTrS2rVlSoOK/4kVAD9V7Np3NjBuxJp8kEQa
vwO07yyZmwA1F7ChbBCM7JNzYFe8XUEGt1kTCR+6inkDrz63N80sAyJ/rmPflMxKVBtH6cN3JH5G
4zDXFIhZ+HEmhSFk74vQZjC8OBpLHahA0GsZAxqY3Pq15n31Sb/pGaodoM7AHAiKp6zzRC2R0ukk
Kimu13LOObVBU5agK4gUp1HvhZ5//YZvyv4o7y3F9F1QySjvw0IBmQPgO4JNp5VhPlYsTft1TjOp
pC0z4efPK53F63T3ctqSfKHfhrxSYhM5xB4/LmpAhPHiEK6wXZyIchLP3M4pOGArqHgtteg2hyWb
sora6JYFdXKZ2l2pSfd+OAFpyZPuZIPVE4u+AOHACnMz9Glaa2p5+0/7cr1uwKiEP2kD3Uu8FV4m
WDjuuyvvLQX6I3T34Fj3+aWQS02EcWd053BdVmoABIhftPG7NaRFdVKs6JTyQkZdSQUMFESDUuAM
p315qp9/6PbbrHdwqeb0c4kq8iIVgFAGdPSuOFdBk+ADUvRz0yQOJK7AZ00w168zI1bX/gRZN0sP
nCB9bQU9AoYC3Oy5j+sR58zaxXn4IlU2/05Rvz+j8GvqLMaEygfplQH2yIHralAGVJpUegTJuDkT
/WvynoHLqa/mgEZARgT5w/asEXBaOcS8mlMJTbSY9FOkYTe6Vs8OVVW4TMEimCflFFgbPkLUj5V8
GLOlfGwgSINw1JJ/pOWqBa62W77i+EuEVpryugKU3+kDHIU4hqakkuTHZZp+uK3SfNFTZJGh2eIW
PkQlrYgLwuuwOVzWX8RS/Ye04emf3jr/K5VTB/1wSnrZkt0UtjlLbGf6G/CjLQWj3rFNVQiv2wd+
JJlLmx3WBolnAd6OScUZwKSisZNQjWV33ZIzIJfukztdwf5o6yUZBt+D2jQF97e/7eCtloCYGIbr
T3tajHvvvcg/5DibUwUZ4AgSWL56ipMZ40IFtyPR363BuEMBFwOgffEqdhiSITqqhWWOJXxUy9Zg
/cTs+7qYeqs4wftLE0dPotnbIdxhMeMR74ErN0OxCKZP3OdL1JGO4Amzlqrz884jEdcwKzHlTkYV
ylOLy5G55CEWQtJkmoQvpSgiLerw5NCKMG2Ba+8iN8WTrtqf/qrki2kWC2omPuJvcyLd1dzXavNy
Yvp78CIw5XIVmqjoV/RDCB69O4lRu0YptizXUe0b+zW3970zOU9qZlfIQxLzQ/FxeyJ6TOcdpF8r
RRME5/pS3eNd3KyQqXJWT5+NlUDCI30TZVXkB6RbetgbNSzMsl5Hcfhus9X284ewnPdRjj9QW3qV
y3jAOkuNG+MUs64iQlZk2FXBhX0H78fL1Y8NEu88XWr9pYANQ2qCTci/Hpf9edlNb621EmiK8Zin
r/AZQeeF4+ALQL15Dp8iCM2dY7iaUc9NDcTZQDVqh4AvIsg6fBhIZQgXIzyAb9wtOw1aT6MuPnuu
qKmdfFhNXrsC6N1RsJeQVWKja6iT7gu/tzMUS+uYBL6OZvvTBc6oB8zMtg81Jly7yrGKxupZpd6F
5AY2TIMZejLZGqxcycAMX2vkhliYKKjkwIhXwocHd6u3mlpktemc6iav84VNJk0fdQKi7TBccUM1
lHgJnKYuM3AMty9BuD6As0cq+Tdazze7OwaT8Xx9oLGoxxbkGwpj7OVu+oj0lDwGRX4ianJ9gaL4
kwElmpmPM1jRJ5IvjERDt9ahlo6eD5lLOsaO/cwTlbYtOYZpbeE5BCwW8ObAGt4Fv0QwePxrvEyi
olZJBpIU6fNuQKFJC/yE+5KqKgn+bj2XqHQorMTkDYrBdeMGHm9+5YZGI8ZO8TrWZT7PgVI1HJpw
vwJ4LZiQ5PyBOK9F4l9YslkpFTg8+n8Bu6EkBDS91ArjoVIZtfLYRCY2YnXOF+7JV5gOPqqAtLM/
ikpeBQdDSF/S9n3YqKULXfBTKFpVyeB01qYCRzIMSTfFoZJwCZdiGbLAkc5E+sRwBmCjonBJ0y0j
aI7zy4Edf5njKk3C5cVqejkVf1BplJqZV+dW9YQdrxuo/eG+f+Wlcr1dkmoizk1CquOsmNBNiXcI
uJ7ugt0Tp4YCWwlDaiczAudAqSnnZJ4XS9G0BFxH9LyNVt3JmhFbhwu41QFWrWXKWVPNFd+GNPeE
PnhPelNX6BRl71Ax/XlHA14BcDrqxGUhq6tHfelWWMP3IYDcCzNkF+UEc/vImD1yH7LWgWp+4ecS
Chd4DcQMjd5rrQuNRCr9tOI9rw2MBdMpuhIkRIZ6PtBoMfRfqvl/ECb2NuKKwcgYSbBSqdxgrPD6
IMlgDsPIKYJvEVbJMeiDPQNp/kvDyhRK9lsImgbZ5l4n/1fOxSFDxd/rinxLk9A3CBNpOP9zGwIf
FenOa3r8DDxXinjmgOQWvLtdwBK+Uhcg+o03GfoYle/RIEulg8ynBFMIrhlu/65WdjMYkiTno6ru
EAP858E+Nsr6ae1eVQMRtAAp6mMsCOjVWbOLLZCP/N2RP8zmAAKMkN0xI0lH4gCGS2rqrQT8uDJa
eGuufLmQorPEi+oKs+XP7utOexh9VgdWMNyH37O9gTVuPb0fH5KZb0uYw6z37QtQRx7XMPorrFk/
3ExtT/3FxpCrCel2F6iUzgXq0aF6XcLisYBSYoD9zDh8D57ZkZ7Y5HqY5+ygfA8PNsmuE5Kt47yE
FNC/0H8UP30C+MsJeV6G/pSI9hCIQFVOLobCbdjW6GrB71kTiOGdwmPUxNwVt07H63USsvTraBWQ
BGQTyTunY1GIUJ+wRnpL6vAghvbC2IT/xXrStiFCQmqw7gWve1kuj+ZtkOB/GWTq3KgkKYdo5itJ
BJWkZBwZ4KTSwTBgh5E9OkrGnyH/4SQGPaNW7qh65o2HwZtILTY8fW8THvMc8kobQbpOwTKqxG5s
NsvXRUq2hmboTipJ1VqV4jtjdI/aP3nisEmM0fmARLpKLz9lD1SHTpks4CNOqXZpGWFwXz5cMgbX
VdLGDeGcpaZ1F2R+coA39fi8wnG4JZQXu75VBCGWvfySaGb3e1jXzOdc0Rq40m48VgrWApP23onp
1KUDmYzhZt3uuSKWVfP7LSZJiLWBTe4Ay0PbWt4u/rgcOx9t73+FXw8KLapKVGnLI48z+/woJA9k
seXTsZQGGnpXRu79HcAPtr6f+hH2DpBZGlm4uuu6IVBn9xekUkisqB/Ge578hLqtC4cY+Fp96Buv
wDaQPzRGVfxQG1GPwm8jWB+Zumyn/CraYoQFjkkcuyjeviMH+2zPzPFYWxXYz24fHUWfxBk416sI
oPumS55z/UxCejMaw7O/WlQIl+EE1YajOvYg3JeNePsxGChYLQCysMWnECAmcH0VunBFSho8mdcz
R1J8SqUVYblJ53lItA6iZPjwuioQNSY0U8APGdT+J+scTaOmROBEae7uciM0hRY6Yoaiq2Lr/xRu
l3JiepwQ+SenksDzHjlhZ045RpkFVaoNuK3dZtl/Q5aW00Tct+foHqmcYIZ7AJHzF5zEOYHWwSYJ
8+Tn8gCQ/QtUQHiOMAue7wjDEGQH1stVcpcWw2m3curnideHu+FWimkNPe4sej8Ec/IUcD5RG/j2
J2xWbP1dwjnz1i+BzITd5/jqJnAvAAk/esJJReQRL7bNRyx2IMX8N3kIH1vSBJdh3b6p3FfChF+T
EOROg/bs4plnhZlp9jFlMa8ThJ/n0qheMl28KYggDB64Mzbaqn4GtBbS5N4xPWYY9igea7733rWZ
F811tpXWNhZgXLe+o26T7UNe1/px26053mAtpLkHsirvExR9WakXTA5FSiawcUwuZfjlGMENa65v
cLozeiayjQdhnr+tmIQulxsofFgkm+0KuXu7QLMChBQMVV0+T3etMSPgXjuO2qoxDp7QTtJXfYHh
Ha6AThQ+VXewpleuaV6X5t/y5vM9eFrJ6evDBxUfi4+AFt3u/GhA6AxiIe96jfI1VnkMxJIAYeVn
toT7xZeClb99C9z9c2O7PyKuBmdkxra4Zg0dERkWQWBlGimaqum2de1Hk3QDszGwUNgGJPY53fpO
0HEdvY4AdVs9bFmx6Q0kPCe3J5cUzpURlALfzydF8cGEXvfAR2jLeCrt1EDhxDv3GCZosNwboDv5
/Qcm2WweIJUy6dLncbh8CYcjklVSR+Te5ghm0frzT6qzA4oJ612yjy75b6PWRWliiTP5NMQQhyX5
4Rpr980NJRqTNyStZeP4vz1PDYEgw4BYjDrcHDyLNio5PW/VAqThty2b9ajOe8pMOBeDGn+VdN3b
WiZHQdmiXCptlNGKvlEQfKRcLDw99LcnIDfCVsnP4MjW6C1HoPMXEa3ftbw8UjhRKQEpb+eSSMrH
7LqLokEi3GA3odJAvlBPeDkH6/i2zsuM9CDUD4f8z9TxhjDRWqrHJVJsGjMlFKhOeIgWzqAN23qz
PXv3IyZTfY6TIwV1ntkOe+OiVLmBig68sQraqgw4VzueW+iSJL60YKTcwzoU4AcCWFPaDhuzCzPG
sA8x17+64k8TAmhI/FlQPMjq6YYpnZwFml+cqweDDfaenNK9PJCSzV1JqrvUAejdqNXueUZ+9AX5
8bf6++nV5YJ/zg1Bn2VntbC1e9OsNfa6R7rmEaQGy3K1TwDBUhFItgpIN1cxCYCkZmYk7WO1o71o
UMH5ANUv3+7Kj7nEPozssHlVKYXpilaqKyYhMiUVAWZy04X22u8qxeLbGus8LBXwk7LkpSDntVN1
zc2rI9rO7HVVkdrxepg4NQNl1eV6VNXarXQlj3/pRIJtNM0l7jeARfDv+B5Z7Enb69nSW3jR9dgQ
kKCf9Kxj/aFNXh1EABiZBUwxJkhqwqunslTde3kE7YpKgHetlr49t0vyfDP5rbx2/qmCFxodJS0Q
QT7eyevvCu5hWikHvJc+3Glpbp3WhhlAcOPVYy0+7x+fJw83uOAUcKokOSUXMshCewbg6j4nriPw
RkPWPCVwIOvgkCBtnedaZlZ9DyncEAj5aFFkLaSQDiPoxlUbJCL2EiW+9dSjlk4+x/OsN9Elts6u
i8V+YWFPFdpqn3zu7TJQoUoAhByZnzBnvuOpe+HN5xxLjALSwRb4J6XTc/L7rGINn9NOeFRnIG9Y
v3fx0zoDvH+XSecKs9E3JlnK2XHOPITXEis/XIyB7VJDCPIvoX71eanMuN7FPENOp39/YOExmwB2
/lHhA6y2dHLJthmwVcxpSATXyMNfXoXj8r7KSVBWSWRWFyL8xYgVIv6QExF4kYAO0uesvvlgMxZL
BbnNpuXs1doDBEJYTYSqdO15iHEiCaelwuJXJz8wkKJkM/w2iB0rHKDu1x6MIZy8OLXcNUErmFOs
snwKHdhjft/Gn5LlN/HnYGLQcIp91xt/mXgJ5TYHIhIoQkQjZkcCUazW2yg/ddEppJToXekHwtTi
mbKRRqsn55ivFCv7AArKiD9wd5FbPJxfDlLEeZ+PXAQKGikjsilmzIiXzoehGgxNMKeQRg+Va0Fi
sym53wBJhFl6wmnp61Rcl/uoQ0xW3ze0+KiTl2R5E2ufp4F2fyORsrDcMnRHCJckoeOK2MsrGeId
lzgITGcFyHtm1A3KsnaUSndyM9bZimlTnnchE66fs6jZyh7ONb7dxOrk7hA7rNW0TpVCjJ90FSdw
zAbq97JkyPQK8PC52h28RtSVrr2GSyPrBU/BCcaJFmuYUMPUZVYnr0jxm0sUEthO7Zch1y/2lUNl
ikedMn4ZvZVqZhWWyvx9aYSiwnKzciSpPUxR7LHvtwf0+qK9s0mEhiYNPQTQ+9i0FnMfgw7Ug8OO
oiiYu1P8fBUrwr3o3DWguToj8gZW5/pvXxr624beDxVkG0kJpUu3IoT44e+dA483p19woVerRIoF
KhDXk82gLxT+d0aEvmm0Mpq5WcXSuKCGzjEs6Lwww5jGjY/NNnOFOQRvtfKDSJixFVv4fPuJa9+0
9aHAk8yWl6W3NZX5bZkERDQ1PQElvwQ2SizJMqFvFTxFFi9OSK7QHUBtcYRMJpyqYjZlrERA+BOO
AD/aSFmwbbdNmOVumg2WTH/hAT1o+PFRDVH6Cu/kS5Anr9HO5bg//K6zsod3+sxh+C2MEVmVUHDO
SUximYMPWkdC36K7RvYS4k9Jeok7QbB9r+HYBH9A1oHWDGo+EwmKTEDC55sBPyyolV09pjfEwZF4
4PXjibOACsBu6Hq8Yi+GIh2hWtjTAxIViI/MV9GjHyqbTQo2CRO8E1X6H9Vnz9v+RiM9DGkrS56p
sDaOKPiLrkcHc9u+P4APtoQsZX4+qv38wiZY2xgaBpxTuOiEnZLRgxcECmsEAxi8JhGDnHWmCFBM
R6j2GWweSDlrl7ofnNnt6soicN9XOQ+/rMEL+cVgMG9Cy782fPR1J17waQ3WJceRc+XbgKIkGTQ2
CWDFnYbLKpi6D+jQ1HnU4hFgv9nqUWebrgQodCt4QzmQGA3XbZZ2zFGWm7F4NoajNO4IN4KlZ921
y/uKub45i47kAYZj7BIsrfvN+iD85ltqAgF8SdBY4R9ZAMPKuiZGGSb0bRqQB+MB5oymXCbsUgoo
pC3Zh/DcYhOlcceV6tQvnL8AtqlImdxVZ9LvTB9IG6rq3iQh0REWjnGZu9PnzhKDbkVf+TUuAyur
32tAusIDpwprNgCBnj4rTI7k6tjir1XQ3uSgEzPztlyZ0+phNzdNs+X6qk/iDTL9Mf5l4d4chSui
nhRcfmdldZJGOzFNx0dOHTlRpmL5YqAfbIF0BF4BL0U1qhD0oGCeaEB3fjeU4FwK6lRtq8EXxYCf
rGW+HywB8Ii0k87nQ5uy5Sf9LeAjiA+RUnkMtsntch5A6s6MZyuiGAJll3+0OTTMG0csfSNZPjT4
+izDFiy9KnObtZdjncemGUf92ppGYKGhmqU01kgtr39hf4Wzm2gmfT1mjtpo+YkhuFmBvGw/VaoX
59hznoFSlnmsLjOlu1ZRZXEqv7nee0oeHEZa8qRQSkmfHBO6GstAa8XAOzH0Q1fFlabL+WnPw4Rr
X6tIRXPqFB/ho7EHC6mVofgpyRGTGmpidIjz+ydFrKPWu5r5JgxMr+XQIk0nrL6v8q30ga9UngD8
OtQXOx1gQPeUwSMwGDBoFjJNICQDP5IWYO76aSkoEcOodDOoTPoDT6bRT9Opym3+VOObWevbcQS8
Qs4Zwzvy6J4CAS0/eljs/XJA6kzOVoPkZkvjGvzUxa7RQL4gyRwgYMyNn8fz8w0KQHG0KV1Bvru/
vHGUz0dMXKvFD5CcKKuA89PnzROmGiubTTdZENaEf4GPTLGggtIng/uM7ah8YHfkU7AZDqheZ/RR
p3hAHdl4utk0flxrfWm2G41mJ9f/WVY/ep+q0BopP41vzK04ILVmpgOknNn2fFGFbGVRo/Z31N4q
ekadaN9ZwRxSK/t0bLN66qXKg8qaCltXHf4HDopYn/0zKkRknrAtLkTQa57v3oSGyIUi0BQNs96z
djVN0fUygSPR2F0MXeWhPOkZivjW8TYVwPBYlQnb/o4fzWdwjgQqazLKWO1Ns6cXL6G+APlRq5h6
bS8t8WIjwOjWxGwXZcc94xqssKVPlGh20JtIsoZecCGX/OFMbw0zxEvokOBKx64BbQW2Fs8BLvgE
04DXzAeorS/qL2QObBy++/n5b+ExDZXLVGv/KSJ62t3ghSjgYUOyMkeQIpNzqv2y7KDUiclLcU9m
DLzkoUZ/H06x52eHT0bnQhnDE0OyZON0fV6peYE2nUD2C4Rc/nzLblldP81oTxYG0M0cCtPjQC1b
X9VqYDBIOH+jarRAbS2RqreivKNEGnixVIIfQsOdoibaI+qm9AtRwE6qu3dpdkVWXtosC2jBeDwn
vJpDlshRDrIXQQWo/mjz5Urz6CCY3/scXlZdauhrsCtCu3+/+ehnmI4iobncUrLXhxrTKUkNMEFx
AVKGZqSpHBM0tTF27W7u4mQI3vS/X8bwnUsv8UDVyWW52Q1ppSmEQv50LEKb+iv4bZsbhhqhk3lX
FrTFkn1xNu1ot/cPQ6ETtQA3o1L/7bk+F5wuDxF927XbsCagE/Cwph4RVbOFpY/QiUsrjl6rQbHc
VqyVnqDNrqs/PU9sU4Q6vU5l9HwbB1tGcBRcSV7+KJ8VoAScyAMa3J9r9X0skZ+k8FerrG7W+T7C
py6N0CzOfqZmSOICxhaUsFcEVkt3+dxvp74+IL12EnQQlwwKpic1hqXrQFIRYCuwlj2HW65JdZ36
ZVUG50M9xIiwZR6BszW5+evYv6aV/xRxIcM1AqWMPOu72xGGMdKMGQzqNxiUxigSShjltSEbLKTJ
0LaYKCuUBuMXPXvjeepWC3n1AKQje1CBUHxzb637eiyvAIOJLAlN1UB3PsjX4dKXSKRIqwvM4YkC
3cMaWaWddzmViK6460a/Gt+5TVgK3Ov4eMqt15UIS03jFeb7vnvj0dIh8Yk8NXcSq9Gz/Sbc+oN3
3w9svC4gRrTT5FNeu2K9PR3F9D5VL2PdptatHr3Q9mZ3NDOJdf4OUJnYWgJYEbmrpL+pNU6UXRUs
D2x0XaFOHzeIrdM8trX32an2ALQXdiUJpgh8mnNgbaGE/txDu8XeJg0zLfcFbLcsRB6PvagCXZ+X
tepIoxaSRru7QAbg0C8PTDHFqgEbFMj/PmgYelNQOYINprMj8p8vhsVXhHAgEg/o1XyaoNpCbspf
EPPzDG0yaF6glZdiywfX4RxjraJPWvIMVaj0NteyZ+9xMvoE5DZucURr7+sRRPgGx+YoabBKlVlx
B/dAWRL0Mbqs+rw0NhANdqJVqAvt65hv8lvCg/fSUdMpTYGIFDy+7qzz+b7dBpCxoNCvwiJrJdP6
MgeXtDSD0a3TUMD1iSWCBygDQRlJtAgxMhhpxTlet/O+aHEm5w/OF4RLrRDpXvleQf1xX7VR6ZSo
z7BYZ7Dl6X0IZz1h2f5CmZgF0OGqVK53Q2SaHRbbhprY1CqNomrnmprhC7hm03qR7WKPb8cB5VCN
AQuuDY4WS4jdI7dKr6hFT10NBwbYL7KOvnO47p8ahQRUVKL7edDuRj9lhwiXNzvOKMbtZl1UWDs9
hMhv1YlTBzh/kk6uV1rAe8jFFuBkDIuZ6FfOcamBci/SLvqMA5Fj+bBCTCIk4EMJyw+imrG5AzIC
vNOSv5Km1J8xos/e9pbizerDbHC61p5uO2TX1wn03g6VXbB8VhyujMKN4SY25qfyRmO4aJRQLnIP
0JHrW3T+MAxO7K1vuxTpeo2dUQhaUocK/+iSjgQDe/13Ej4xMTQdg3xD5Xy0oSRz/ww4A1mT7GRb
RK4cE1PdjA9dfCH1tx0fCQe/9Zh2QJ0Nyv7bc72ARYdjaEkHw/9+ibz35HYa+5u0S23IwjVVZUHz
5pD1J9aRg9qvhHl4LvSxv8azEcZTHVB8rvTwi/I+yV/YqUspaN4YsNvamhTY+FAYquvgXhqrjVf8
xTLTv/cKMLATZ92DkQsrfTHm3+5tY87++NyPgAyUIrj7fSeR0mtv6mwiFeyb8b5Eg0yL5ESeWQKh
W/wPKI5JqBx5i2RbMR1ZtGZP9J2zms2+7MXeet3Q0L1LVK+xi8hsxVbltuNq2ctxPIrwDC8u8X+r
a5ZaKz4YK7ZCzpmKJU85fA3zxVxWEDemPDY60rp9u79JB4tyBn7SGE2xtC4uZHYTHddeQwzPKBmK
7QHztpgkPMYLUzhbXktY02JJ3PDuPSK/22Iu41YGMiYITB8nrI4absXnmFqJnQCUymmHPMXHdwtI
fiAZ/9bGtk09sfKvULCcDIvIQGH7IuVBuz+5K2c2ykPtQaXVVGbtGPSqDXdUkAC4esEs+mmmhh7n
/1gxp5Qnf1M92UdCpuOim65Jmdg72faL6a2QFMXqfDyMPCpGrXe2iQHJ7LEXaGkAfpbTETjZqNgh
7mrPMqQF2kVoxQQG1bH5H1QJ5mvCr5QyudDADM3vFyS/LCwVuU/bIhUuFALEhauNlS53GUZh4B03
EXg6hjP3XWSf+YqM+gLTkPG66/TC3XHXGLxVZjjR+7kExlL2WilDp3yADnyMQW7yBKc4wnCy6tKm
89rStYDujPey/eOixTf1wycdUnbFN8hRDQHRfnM/X77p6yiYorjmJPVC7rvObvkxIqaD9Wr0Hvgz
cevBPVIxJKgL+aJoe5x2fte1AY/rtx4c+LhrigwrmTYF142t57jA/pHbteOykM6IXsYhP4WnWivI
Hhari5x1GQ1WsgHR7xf7zBXi1i2vK9+/HfcSUxhL8/kvn4javAfCipaRjxNVADet5UBpBeYzTL1x
jlq/Xk+EAJQOFLSFyNxjW0gZp0Q7lDSucPL/RgjxwJUWqfm1hH5xLd/WoHv/eWzOwngE8kX4Uf2M
RVKg91PrDeryB45CUjdmHMU5oNkRMRwVuFGVDkmD3/i3K+JtaD/XxhLHqgCEjA4smjUFJRU02abM
oktGdD0LJWnqxQyvUrZIzaM59duPnfUer8l+RRVe1RI3Bd1vU2qEY/HhGiKlp5N2JP/tK57kR+7E
PlnbnNckulykKB5XYYCdSUFx6yX2mZExyaX0j4LpmUUo7bd1vTbAaL80g8RQtFEcx35xjswzDDzG
jBsddhl77hhSHRQUtu0KZA4feGlS3bnIM62YhYVfhfYQ9k8ef6mYJqbXSVB59blri0CZwH8ts7fb
6EWeu9Em/6X5Ff/Y7yaw0l+Tz+w3m9jmqKZ7lWnkAKBgVllnd3b33rOhgpna+z5RM6GBS4GK7fe0
yudNH/bpa/+tnCf25q0eph5VF5ECQBRFK/JG09/qJW4bnke1qjus37v1D5+xzBzEL5TBR6EqDi3O
wTLlYOq1gBIWc97E9AiiEmBXX4jJ5spCkGN7EzrHpN5j6l9VZaNMMBXNSphSejMexQmyduxWifRN
69ARbmSd+dY0J0e/5LcJ8al4bxNWHFfxh8r0rtE/1sSb6/PwQoNtnWw/GEZkUZVETwwaK24IdTlA
p5c44PLbst0cUdIGEcxpXAhvAg9rYiqYh1S3SgTgO6m6ydi/euuwH9tL5zd/AHwZ5BU/reR5UOgK
6kmlqMEl5H0iiMQFQSgAxZBeBianAcCPUEVTS8N7MiVlJDu1i/cW50biwszpYZCRRCWUDRO+IGC2
X7qflYD1/Prr396w016668Gt44X4kKcPqUGoCkInG3cmot6p1si7gMi8+uFcIccjC1cClRUb0KC2
cPtdrcPhyUp0keoUtxUSct1GgeUS5A6yf1FeGrdl/P/zvBUc0ch8REXtp/y6r9L69PaNuenyuzdY
QOTRi/oevdZuDX7BsZOUc6rKxFEXLs0FoPPSKWFSXu1P5YR5gA28M95YoZDsZlCdpZssdio2BmG5
fJ5DVbUpEhCdTBO/KGC6EWzFv7mW2DuySpRoUaMO7XKu8fKerazW+xcREvL0KPeTtwuN8SLQWlfL
8OsUQd8DZ3p0NcqhRjDPnpwGdG0ZQsvL38kEtdZ/c3VIThzBSCOIGJt7s7vCMSJ0Yz9NFIZqVlfY
bYFAz0Wzqd7McgGDiEN0F8AIkWUGEYe6sJmbPNEk3N0qv7wmvc31pBDu5TZy+8iLLKuKHSPx9D4M
f/XUcyE4b3bYfP1sdxluuyV6BQQDvhYoVHJqTftpzCQDJpnTQ+gHjqQrqJj9yrGTDipvOfhcoPxe
jV51sl3ko4Al7vzYG71v2XcaOFj4DZdp3ofhxAIlDRAPiAp7v3EHu+tmqwTzWArDoUOhKVYdflhi
mS85yANI/XUX7nlULMzwdK7nrbQoEIxn5EhTTWdvdmKm7QDy8nJucZunxBWmj7WoF/FwaJVLfcT/
s5WS3k8QnuofZTV942upFgv500K1CpDzOD7diUnGt03KgbFVVAwWUBJVyyeUcjb8qT/9GNbIEaZu
ahvwp+ZR5AU5d3bXYF3Ke5Wh/GyRFn8EXCCvqlRmzgpgenYo51nPHDhQ5nj0ebYfLXYRG9l++6yZ
65/PK2VWAu/0qosEY7aogwHn8vProHWvIlsX8uwEfW0nKbtKH5BgffFiL7RwdQiQMnByO5EwnmmS
Lc/so/d9zUVZxE4JjKQ6wE61UrBnuLnIPWLU26Uj0ApSflnEGEl1h+oYeiGWOVwBwoHLK2x35Nzk
Kb6w1kV4kVlwS7gYRmSxKIwWo0rzMPBEHK+LCzi/cxYARiMp0e7nc2z2ykTyFr3Ltm3z9qJ2+pL/
DMuSTrgbANBBCe19pk0RsnWwWJusWxJfx/v2w8on7wdhJgM/KvYWrNVcH42epTrpsk59ZFQuUZCs
aL5QQ5JHJmEyDcQmrijVXrWPFowlfdwBGKNl8SrMq7BXQQaf6gUNWcXmefowDxDYtZ9dbrWm2AYS
KwXBuCIsav7Wpo5kq1bN4zDk5WcUj8XvGs/mUlxu05DrXa/M9EatTJRHQW1DzN6F1lNRZ5MRZ9Gu
BBTt+HalguJhW6j4qSvSM4N22P1SjFvbP9DjtNRWDF7YMxak4F8H4R811tOjs2zRS6sywcM8A5sa
yTRrugs5wgbsFCvhPrLRBNO//UIPh3iDWEXviDPTphEjEkb5fyHRNQh5w2IngGlOqPDSGQy2r3RX
FHIS9XxSD8wVb4I18+4nlm3ladPrJf1uqh4EmEtEMhZbBVplSyzj2az6On4+gpIlihbWdoh7dboC
xB3fIQl2BH395ECmhBY08K89BCJe4Bcx0vKS9DGyYWM5NXr2buE6+XZLxnJXjXpynyP+HaFevoDA
L8UqGuHjHeZHQtQJiwLVUpu2n5gSXKMAyEyF3cMgt8UKKzL9B3LszNP9aFvo0NLOzR8iyNbiVPYZ
0QyQ4r7wy3V2NHCpnf2OdsI62NhJwEFep5YTd3xtHqOn3PycbdlGA4SIj3OD6GQve0Qg9gDLKYsl
GttIZwAQkHn3ax0VqoBxWFMo3D5RvoRnzVWbTKbUgfALEeen3aanslgkzw6BE/KvaCfxhUWCvN/J
pTq+xSNt4wRdH5iAsZG8e6oA8xDwgqt1P0BCQ1eDQmLK1ItvoU4Aq5mVGL9j7Id9YFIQaUhuVUjR
xW6wO02B73BWhTcsJy/hjjBrU0vTPI0qcD8/Tr4bFe1MP0vIkVTWPIvqv6xiMlxS57FeEUcD74tB
qywUpZPb2V/z903UXjYcTIa0lBei4O6Iv+vD7HgjBGU51MKzcBUIkcNwXqoeL1jugxu0bjGf/s2U
teu9U3KuvfgrPTVsa9vYLW0khWToWo+GM1Zxkr0CW4gqjGqmUG27VBNJY7zLQqcj9Hg0Ockl+zAV
MKyn7wR0+diU98uMJa1pJU0fZv2DuVaby5+CVllKizmPyFGFGElgb26cForelN8DgNDmFcF7q6qy
ZBqKNMFNRBeW/AnZElrqJRsZ5e9iuDP0PuCB1TM7gTMfe+UqpXSn1cJzr/fjt9gxlWIBS2APfrA1
xYyBzU7WqS+VprgPp4rqCy8EAlmeTXDeFnUM5c6ycu2fo+IMjGB5aVMtrbHJOvWlaiFxSmRWcs8s
x1GNt2GeYL8Tb4nu9JC3aDoMIGn561hmkCRLs15L+4CK5wFN88IKbJt7WTWKbFkoAOVQRKa0slBb
K6eNoAcrdOAiahNR7ByFg0dkYHyqd1b69Q7Nw8Rj0ifT4a74vG2rTB3I2wfYWjKTkGxmsPXjJz4T
LwXUFrh0SgKvVJRGDHmiDNTx4TRIq2DXTXHVADuiISdU4H9Y71NHKVdHvrdnXIvxRm7XpBzXYE4s
mHAJnZ+4U8ep4EeDoQ2alJLhT2pxQAdhS9K6LgM/dgHHmtcl2iVMBxkqaAcJn4jZZb3SMcJ7RWRw
hij7FskzYQ6UX6ygVuWJFxZnnlFNjw6iR/mfKWrEMO9OVKpBhb88uL5lEJcG2LaTuuVxpIv1CBtZ
FP3daB24Rp7CzaU9PwxS7hJQrWoYX7f5wzc+m9hR9PzDGNhPjAMqaJYiXWFLmafas2Cp0D6oZ4fU
PoUUmeYk3r1+mLeh0s1bTNMKQNwkpedVFT4PAcAuW0t7egUxVkfCe4I7DrHVrYDUonn/fGI/dmqh
ifMWepMA+pKatw6O8UctOk/07z2Kr++6D5/NYqRPKjVyMcxflwDyNET9uzDuz4cFJV0cXHmA6Svh
ScAQmOn5FzMPnJ4hmhk3BZKVaOAsWyxPw8oB+B3agdT+Cg4cpY+S7GQxnbJ8cOLCx6A4iuK66iO6
rz2lWTHowj/lIJN2pl0is/qaueJixDfAAOYmmhzCumpg3OAmVzNrf1+v/rNe2XA5U04LgTH0swmP
ot6ejzaMqRceh7QMi85SkPd63Cbc8KjlpjLkNE5XfS7+SmoQLactuD2/BTUkstNxE/NfWtFSokwV
6suSuCDxL4gt5M79d91M8xSjwhIfpYeAhkk98mD+iargIJK0DIXo9FTG1DPfj/1Ihw1fdHepAB3g
sIWn8UZF/mrROiO53ndrHGuR7Ofi35MNo3Ho290EN4KK7n6oNiooPjAuLpJ0TpB+r9F+9e6Wfcn5
cv37nYBWA2UJqmrSiDSMdE8ZRnQNHyTZMqdKQwj4aPGJySysFupuLaLAy1g/r9OuvHN0cTumNRfo
5tTOAz7N+Dy4sbdAdUtLa+b451rNcTQUmdoEQDnVdDe+/EaL/yWv06lGr3nMkBiG1NiCzcjt2vI+
b6K3TIejDIXLj3umCO8pQeJFljPwxYcOfgGd1zY0kyWGWVwKtrLIcYTUFqmYcI72wnkZnciH/aVH
fyyrzCdRnuiNI/ii6AEC2QPyTKSaDtQad31AthNOBfx4wRPyfIbLc8ED1ucCYmbTikiJUC7sgWRZ
r4gQMJ6BNma+OGFSxeDTfbs6lo9DUEQ2QKwal2kzGztJ8YBsC6e2cSJwXWMEOVt9hlafzDOgp5G+
1FM6wUx4IV8+JgKBTyXYpMhYMe5mLfzOcU6J0AX14b3glDnzpiP2zGFPlbe0wr9aGqmGNM79VwsG
/AfpyopjxxHBAVmHib86WwvDJzF39CzZSQV7Tm6nETdrUv1Dhhak0HJxuKdEGua6U1zzF54eFhr8
ZfNKFmNobRuEK52cdyIIbSxOGBLu6RzSaU1gYfwFbSJzhgUlqG/NcKH+T20UA17iz+lqAs9ErxDg
7oRC+Xm628YtKvexbccvF3k/w5JNPPin4Q01H46gFvYInUmdIbtEsK5OQHDJjBmBSrs5XpcRw/bG
Oq94Bjykn6cQFUCNgjhCvfNLySaetvDwo2UOHQl1QEFzzpwOJlgjjAtI/xO5dlWpifI3uWTvQB6i
XtglCeGcBA6R8cjc4Ja5pi3hcyTYn7yp1ItN26HSzc8I4w9EeRj5yh8TwpKnvcOMrd1wtVF25ieU
aayDTmvWNcpxHEQOPsEofYV8ddAR3nbeiCt++yTzoXAjk9rcduy8O/y3nhkDNfHp2mHWzDoilWOE
bY0tAtZQkMKRsk+WFPrBtsIMFBkhCCZ0UIC2c4VFC4TbQ4SpWMHuTc1Q5ovp+R4r54+HkkD9Exg6
T7yVIk3NT7TNZkWejHM0SUjSLbdahfaoEICsfMnR8oKHyeQbEuRcQSAUyuKuj4ofFSK+YlBMwSrG
y8Ub7p4SzDLofEU/aIoueScbR6VSO0F11fayRevwI4u2GJhD7U/V6H9qsoyXmUidcxZsy+K3BeaC
szI/mXXI2eco6QDz+yuE39YBzoJWyf+KsBnhAfKQFDAaehXHeK8leuo7EGOBaA6M79bho0i//P0U
qCBJurqzKQqxzOMrvLMnzWwuGe8Awc3laykjbtsZocrbOFh8e/vV07iExya7Vwl31bCSsi6OeX/m
OsAIB9ZKVyC2S77oRc/O+ytSG8JvchFGBNxZqics9KxrOTXbT+LUMQHaQbgfFRGb/yeNi6vlu6ei
1HuUxUD7lUum9EzF9pXQeIWQkd37O+zL2axkyWl/Z+wTPrcNNV1wfJjo/yByGhoDZ2EDKqd7WkC6
D0E3FMnxshOkNIYraNFivtSA2O8ZQai6c99dSia3l3dpJ3GLYNtdYR2OM2ixcda6fpUwzdlFrPiC
Hj65UQmfetccejIPstRGc6o1FWMONo0DCA5BKgBEcOV14O41M2JECjEfssVSNIcnFO9n0O+1JeHK
ToxjZz8uQ2DO4hvL7IAXWxxKf4HJTI6JiTOD3PtYQfmai/B+hzoacCexTVeH5Kgmer1BRQleoxXj
vvLEJRBIHyA0DwbyOcxaqypuGaR4nNVImMDbRCgJqN5aCArvJFZbF2PxE/Q6x6rAi06548JsDb5m
Q7DEuRTmC0EqjPy71Tuire7l/vf1HYh0AleeIPz9ZkIEN1+A4160uuRxOUDgmXB3KBDUIEJNZfIB
w30X7KXnuJp778a4rJ6v533b8OwuZ9a+M2jUyUvzsiSb+YPWrSuNTwTm2tDtV1gXkg13KNeRZpQI
5kk1tSMkif8lk2JMUy0S8umF1QhEgvwRvNw4g2ZCZebaRDSDi1QVhUSdSPwtEgHGxVfkJlrwNfiQ
scpDhI3UX4Wfa3RP1FKekgnFmS0zchVUBSO2sIMMz9E56tciYRUntBbDDpdl7WVVdphi+pfotUq5
l4KgP43iirXAHLdv2HYDmzqy6K3Ggns3wl/RpvVYwOme60bkhXXZDt92yLgGPItBbmRmnKE3uuYN
XyCW0JsDTrSvepa72Cfv5wdszX7c9ZWdj+CmVosI3DB5SnolAe34YocDaqrH78b3kLwnXW272/Vr
weUN1D+7Y4h1RJ7LEV/NCpya7mhoHbX+r4nNwqytdKft2e3ed4sQLak89ZhYty6OVKv6X7kabXQx
a1jDYlRTBg18gfDpT8TDYPku81R7cviBiTEoEV5hwke3yQ7c2cR8BkpXJLF+zetYe6ILIUbYZ1zE
oDlHqCQpoH65n1/wmnGfXIp6x+GSgF0MuJ4+jIHKDZLk9JAXoX5g/uSUqePGTyihaPZwykCuGPFM
16gm86fJ1fYuUSP1Usk4HF//+Rpm6mw/KSmKrcFsBqxQuj1/usoSlhntewpeNkQoxwimRPMV5dcF
vJD2p6z9ZO6d53E62AcSnJ3SqUci/EYx0dUzbjLjmKo9lhzsmbRZ6WWueppS5gE3nW8e6zPXhRtd
E8BdhsYG4fThuNEwyptFjT8yAv53eL5/I64ERw6SFoNKbkliIENU/JAMU8hvkCMPtOXbaC80CRYy
K/4wpo6OCJx/S7ibP9sPy/ZdjRwps1QjYz+LPgRa1QfO4sKkXPgChR2FJe4+DUyvwmwkwz99LY20
XW2LfB2L42JHKhCYu+FmFtY2xpqA5ykZpkc1NrB/Gs3JS07i6uau7ymCKlfureduThWTM7ZoUWNX
ISXQ4JaAyurOdNfsZbSr+GZuI3FiEyRq9keA6zpqRnW0YwmubPy5FGHFA6gIr11VO6ER/LNr8+3E
2ZfboFyY80PRlBqBwVHPbWUTsc5yc0cAIBo5eKFe3pNMXeelA9fAnfJVW7+UzFoNAVamupW/xnBT
PCyhodrzvoWe6ggzCMsFVeBlVUnbpQzFIWoW0+rKFjDYTvPwuwGFrsX33hDrXjhLflVe4ZOclkvh
z+R1GNET8myhMvoaDFcdwC8wGQPboPYEfXiv5NI1PszAe/a39QT+WUt+C1OW+iEOu+nYAUyQ2Y2W
vDFBCH+cqcYmhxW4TC4VkQPk+DP9URfD91NwQIu9XafEssUHtdpmxLbhm559uNfS0TrVfW9OKF03
UOBvp7e25aRxQB9rviVAv38kYMhe5sr8/3reIxijU3GefuHrmzMjLWOwLkvLjaMgJ0kKq4GYN/86
L6kt40yevIavXtLpaodGQgqYpHxjnxXB0yU6iwdAMHTJABRkeg+ptxVd/VS9I8IPAG6L9zTwAiea
/pk0aYDmA5K7h5dI8JMnK+CJ8HUsV7hZCLfQxDS/OpHo/evYPxm9+gzyNKio8d+fSYgDHMnF2/6T
QI/8ky5gAowgEPEAJXBKF0pDM5YMWugCjUAm9ldt/XUyLdNi7Oh9KWUvtFlHiPsH+3OQhD9gr8Gc
O7Eqlky2pNK3K3aEuotmHkIY7qxGulAMds+PfKrFtNwZyJ+tysnfs/IPPnkpafVJmTDAuk2G6FD8
6C5xICRf/GwdUxZwXcPYtLZK1mYTUOoa3eY+tQOVFUodabu1u2tbvTV9clc489zZhrWrIsyP3GMS
dfP0jOgKnk0dQHj31PK9VRBLGrPKPTNUvfSS4DMYWpAnckpyCr49VEHPSFYatgu6dcVc02EYEtSP
+x9Yc0lOsV2zQOglYeFlAgJ1wrlrwJgqj0Tdt9A/iHRUUfRptIBespJkrNA6Evjo4o0yfOAX3iFo
ddqvuysRwlHTnMYM2StHYWaIe9hA50djkCwtJAbZv1/HApwHWFHf5DHCfE6Nlw7tUOWQ9v58gG0e
tpxEQBnQwUj5NCPxiLI0n8dNz/VdidjJ5jWIgTqSrKyQdSTpUCBLmu/eaHhY9KJkatndVVdD7w4K
u0sOGcph3ISvG+l7LMEsl8uN1JrOP4eDx9C/pjxEiX5OfxQIAhLyO86vsLcJxNHqULmZV/ljOxCR
RA+oKKX7uK9DshX6aGLSYNDgJ08lw1qigmplwsg8n+43GoumAxkAxsz0fMtY6yzzZaG7osP3zrND
XJ0qs4zOuM8tV7duxvXfOFhWjJ5ztkKzQpkd2nWB+qbQj243/Eam5soyLK7zKtxfX7+uQ+kzAaiz
vx5rwPjsQhG9gZsnaT3rLoRzBTcU99Dg0y3o4+4sNAB46etaBHpEa6pMcSBiKHTQwUK6wWYMx1Pf
hbFDnRLHQDtqYtWteNE/covtB5up14trSCXhgvcQ9y+mcmI+4d9NKq9VS6i62dHpfXgSBTVp5+MZ
+4oDSTLAarjo2aTsPARyKWYCYp2dVfkNEhOTQ3S5EkKj6cJXZ7T1YhoPjmkMYB3fgjTR3eeF6Ynj
w+zpTcmmd95WBj9WQ1pal5sdr7Ou1drmfOMFBWork0/vni5YjmKOHL5CyAAGUOYO/LYbApu+MHpi
rboRdOa5cN8FDL78+BaPI+akqq14OxofwKfDNouo26reuChy3TJRmERt9c5w9XtZ37lTXcrg/IEJ
qkhqMId3RzkubbujhRpSBZwZub+TkwofX57Tki6fUE4GeV/7ikhfNG/6u28iUdfbcWFLVKd1wmiD
cesxyyslODS+y5O2NxXOd7TFfsXhcv+73OmLcLi+HKdfAnSBwiO3W8L97ETp9tCVMKgLjoaEdUfW
j/6QfNo5xa1KqEx6HTr601cB1L6RGIm9G7K8qutSuGqRyT/QQQWcFMHqEJ9BLsH9X5S2HBDMhVaD
7z8mA/+fV/Y809f3ysqAhVPJg1lWoaUmQJWkF8hHENPVDt8TMmyA+LTpYQZe4NR0Q2kqrZEqoizr
7fGt1ycQ03r0fRQPCSDZiNzSQm48DY8t9XNl/YjbQdlGBA7OPlVDqOolcv6INPlTOxEw8hZBnsNe
qnuuBGe94KxNn5oKFTwskR8OdXiGPlL5s+x9FaZtQfIwFQZ5dIJJq+ITGtN1lda9l5P1Cjzaf93z
G1z4kdapf8FRnnuZNuoHO9NqKdi8EktHec20ODX+bT7oUeFlIRI6/jJmes0I4sxFXUakBu1fqdf4
MWXQ5tRtS2w6QJXCHrcqSd5FMFawa2swYm5YkfdiHTNMIZpsJHuG5P40lesUS/3rviJ05QuMVhI8
s/i75GxBb+Pck7QRftW6irTX7g5OIws5dKxH+OtjANcH6y4LQa6zjyHRoBQzcboSONWwotbjv48L
Y2aPF90pVQbVjG+ex5JE7ZfNdMK4wS/pNi2XR7h8WnPVE5qHvcN7Hb7bsAa5jM+FoSYM0oJZ3H3u
MQYumYvuuD1Dx3WIRirbMEaDho8pvUXguWxHsWHEEw5JGxVGg72ehX4biZKykiyo+/iavlJrI1zF
GfhHvGXtNR8djZP7jiI9fUCtuhXoMl30y+0FdMkisF5dQGFVf77Qwkr0uahZ5nO+poAMBtj8UvK3
LLyIfI4X6J6KUqvBjAd4/7wY2uZEdAOnKTl4fDESM+RtwICvtaoOnzoDr8t8/9jet++YYFC4lfJ1
9BcmKNJyK1tWriEBDfruI0cwJtEROWIOuaHm0lwBVeUG4ctuekuGr73Ol9EVb5Lqpe7LFos8qOGA
V1Xup2IViwkE6ge9hWFYkqEMM7+h5taD/jT3E5xU4iYgO2XgwO62+HsaQZoIYAdDOx7pjpV475Tu
0bkH7+N0IKYwhp1J++yMVKz7O+Qd4MZ8JGEp6g86nzgeZkPFr+Kz5r3e3fsLAmU5dub8O7Vx1Z4m
WlImBnG+AFSmKXlNBkds6HbW5oX8OBSikmNa3jO9CH+QvoJqZaFm1w5GyNCUSJpqzJlUEriDxYm5
C6dKzvSujkPgpVF70ExPgFc+wk7zwUcyZ9t+9hkhjle1Yx8c01wTgOHMwynHqTXZSgFc+eqnOSI7
huwdIMReHvk8Cc6c91J/zEW6bLxgfWeO1TwADiS1AEJDwLI+UiwpvhJJbkOAhhfqgk9O9VdjE+3k
kW7kDs7MnOGtpgrGtdld84BVVAD+tSoqiSvr61jr3ZRsvcQa/YZtCFcwnGcMmdhy2yGXJqunu8dm
ojXBEcU+2Qeaa6uSqAn1CyJBzKH4Hv6n6s9j9OkQ0h/wnDDFsQ2XmdAL5YuCE5GB20D7cL6WQCl0
lb/64WwVyx/eU46waJHpyjt8wDsl5PmTbOYy7OW6Dir8AfRwDB9Dze2IEjKHqarOuA/ceeWR5/v6
3qRkbqCvi/LhV9DjvqHpYpp3mISLF9RrBaO0GAtZLBUS7ertfewN2cOlhUofjNeWc9lKiJx3Aocv
FqTq/I9rFJaiM6zC5tVKU7q6gk3f+MdFtUSNPGtxYUGBcCqufgJ5vYJ9Nlcdbg61mi0Yc7kLHeq0
zp4Botkto920PmZ7E506hI83/R0U+ZsZURLYoCFzRKUOrMV1GqyZ7NZMh85YVW7u2I72aW8p9HDr
CokckZaQR01R+mSscnQua8aiCdIuKyYoO5gVl+QwWUhPK3qmYkwq4J4Qly5RHf/9VTQ0gP1G6j2K
LUU7+alpCO50+nBv5KzHxbd5niyICvANfqHy7x/K+ODb6QODOYkxF3SFHe+Z/SFREfFt0gFOY1Vd
dQGPH8dLFfVXXEEGeoo2HX9cZGe4gK71CduMSnPsewnCb9AJRgNiEU6S49Uldb4DrxW5On7DHIIG
TOJu+IFVPivX+956XEdoihJI8CcPwP/stxARhSoJptnFVwbAEola6H279di1QytnSpISiMue8NPZ
0gJcAM77aHolQjYNMULcPFpWjE9pg/md0QU+uEKa9CF8s4BFz2x8BAuWkHphfyLQcAxF+sl51sXo
jJ8Crrg0jk7MpGJuLn30OWYKH1++fK+zTydOqPSVCLfEAOLywVkA0ttX2ZK5of270U816WZ3G1Xp
lHPydpoO0rCi8oqCxz3sASyk+O038ZjQnnLKLRdzlppQS9ZQUCzT0Dwtr0eyMQv2bzk8yRc9vn7u
SeR3GmSoLoOf1UVT4MVTDJMLyGR8fRup+tyocsNkKC84geh8lLreb9LWArfZ4JFqgQnS8wFg/UOe
lzKGC0KbDNlfOzIS99PsU17/jN6n4f4RznKmJb+LThpRr+o2wF50mwqWmunAJzWWHygEBR1ucHGY
N9iaqzG+bU0cJh1Av/jBec8sY/MwXgBvaMjt1VvsNkD+YTwUI0WIZCAhK9Gek126SWTJPFcBZJ1C
AwmiVIrfUACMlmt1m51p9Dh8BgyjwNbiCNHJNaQAOL5BnZAyxpdgkKKoh81+8nibbWiHLXv7yBAy
QNzfIS04z2xcvluIQPhgNyUSd1DyHyZxXryiTuvmu9erL2v0+68LVCzacS1GTH9F7OHbWOhF28IA
yTlKD8Le4XdKKzL0HJ9QukC0dvcxQbl+FXGihTE8WDibwz8IOu1X+D/vE9N7i8X5/Tl3cS09EZ+z
nmzqWtcTA9tCCYnTgHtlICl0PjuLZ40/OyXH5CgNJhgoCqX1HfoKGGCgzUyN9+tGi+yvxbQJPpjF
nOVaMe8l7inHevB1Hgx3BSGhtZu20KoZRHHXeGvOKQErWF/eedpiwjosT5eKsWL1SaH8u+cABDMQ
UI72aObf8BTqsDeF0Sd+RLl2Q0IfKuUuFe/Fk9Iuw/3EjUWex7V8ilzXAppvOf/PCGxA/vyDRdWt
Z/YAFO0Sttz1x9/JBE+zNW+rfohlW2wkFJ3EtlL+olZvgd4VoLfY938UDZGqU6bWcjV9fsP+7GLM
6m8IIXdRsERRpqoeqoIWU/G96yVRhlAQoYHBuR9PU7OoziZyaJ58ixEwlGxPVOik8MHkzkIgPg+X
5l/F6FDiu7ay5sMl26v0/zlalfYg4R03uyotxteFc2XT7Snei6c732DZctHwhI0CScRqyzzD/uDB
cttkYuyJWGmvaH7fATJrhn4SROdrJ38OIf3ZOOPt466HSygPyXq7vc7VJmY7KfTR2W/3UqcHYhR4
dW8h2KU5b7jybhiyRdDJqnzRiT8EcKpYWFE+LuJhODF+v8NVKm/KuO1pchVc8hOM6nWtjfApEioU
TmSekDW9n50+4yffUlkGA9IS0W/wjim2vFxPhw+64hr4gfJEoH82Fmw2Bb+tpLHB8GxTSyRXK353
XoVmvy2fJv6568JjKM2oz59zVTmN8cTJxxuwrzUGTCVc4xrwERS3dlvrYBl1laol432xz4yFpkzF
ilRFNWwy9Cxy33gkcVT3O7vmUfnaby0/nJxU0WtmBEukf3H0GlHyESG/SqHpHef2hxnXX+tYVkAc
Y8JXTB7dfWVLEVjTcB5rSmoAe2cNq+71XYSwY30y72qeFKoVhAn1ZttzvhwT/f0eVdCoQKKDTHF4
OfRdHXbjL7D5KG2qgt7ENExuR+tf37+FHHyGZwTCxuQv24US6PP3SqIopGWWcNtjoQdeQ6eH0mUd
ydCfJXPIVt4NL089xInqqyOTT0wmRuUE8PrkZbRrSaFnGwCmJo/UA+p+pI9xC/4PB5IUeuu0yoVS
PVTGRzXaXcoDCSLEFA1SH4eSFZWfg27wE+KdX9hCtitu1exljBfXGgJ3kueNIx+ky+ru9pp5bDJF
giU59ep50OtPsQeD+XQPrbk9lHaYH33kKeUm0AVA8x/uv413m3a5I/ErnpekT0LkI67mpIayw/vx
7VX5GidJHJLRpykH9nprz9efcCBoeTnEt9R2Ud7pHWRQ3yKqqjU5h0dk6nm9NyHliiFmNI2AUUdw
nKvGZbWQ48dVL5yjNX6XKTcx+s9XZ4nPtP8OslmJaIsaI0bTzs4bC+PIcDgmlxh10S6vDeJluN2Q
T5ODbUA9Lk3yOR/3GlVtGVXhNl/qi9qd3CmS+F39Jx9jVZtCjsdBz1lTQ2c6/3FTdAoMO8UI8ghp
g3nabSv/SY0Ih7EGBeeE8ziPNy/FdKkYLvxlm7i4pCwjCPRbPLfXmTMSBG/eRcDL3VSq7ukf+D/G
lkAnVDNsOhihm1oPDfLoEkJEGOn55McPq4Hnu6v9dVXpM2P7uJ63IHk3ZP4BWdaJb7uuiIkB4/pw
tFLuE3YiZZnHSYxQTaXSQMt6F/bdQQNOEJZcE0dnovHenMz61kfOjHs9uxICE4Jru6fJFnpp0p4N
BEpGBVqUdclWjDRgV3PHq5PJNAIOfnH62CqrjbtJ9+Q2LfWPROuEiUJZhl0D0NHypD/i235UFj3v
F/OcEpPypidC6l9FwaS3w2JCvFPzf4j62M91SiAgRPY3ATnhCmXPK2gDR811AZSZYAunRpztLhny
bGOhhdpT7qP8HVRrbHiGRXggx/uHe7aDAqNuVWU3i7Q7282gMODQoISj8VsjKNM6k8EEWEa9v+j9
D6YrkPoicfV/8vdvf7g2NozyQwY1YKIBROiyZdrDFFMu5h1BRR9LYxk4kQa1F3aMPx+rL1KF6tv0
qOju1ylSaa/Cr+6qhd+Irv0te3sYY1KtmOrATBIhTYV1o6ryewblxNH3skx/pGXb+YwUqJOJyxtC
JZI14kZKkEjplU8XftoZ6z7M0jWn8QcvnpLk68mV8pQU0UMiDH3a+zbjNYm7wBPS2df9P05VnE2o
rhCS7XH+ENjlvQs/1tw2UeCkgXe3wTXSfg5MYc/JFZls71jLx8XhgIZA8a3cNlRNeAcRuuyIGEU/
padedNZGJJ7i/Kq7xmiH+Dqp11in6EisJUU0Vc/OOsLdSgxp6NjfpbXNLM0jJ2zT2Ddmb0G6GKCd
3rphtp308bM0th+Uh3gDumJFaUcYtxdh+U2WxRFY68hMD4PtSl3aYdc7I7FL7kRCeYDLwTLhEaUc
yBv/ts6OwgxOuSLTWjIx4W4okhkVubDCdoNna/7tEnuC78AVTeI/zo2x97GfIAuL7/Rcb7fYgptP
jYsKh8b/xgbAfMLBIehjxVYGKV8M8TTLed4CnXoPCfRK301Lytut1pb/NznfgBMTK5PhLA/rm3+E
wT42bpSt66s/MS1YnxL+tEgO4cWVNpe9GVhzNrU4J5geXiN8uxmUAgl1FO03xdNawxMV2nADuxrI
pLZAfKCpeWGzT2P9FNMlkACOuNzZhXcEyX5l4Vl4As7i24GgXUFlSVbgE66GvaLD3Ack2RvUSwRE
2UJtBRrEnPd0SlUC24YHfcqa1uSjBjl5/FbRTFvhFgmQuLkUwaDgN4yCcFQphYXlvInUF0jkR8c2
uhAeS+sBE5jqX3+7BtF3MstcwclRTWS32b/owigh910Vd/hlzGl7jalHEIha2GkXmfDHOCqRo6D1
mb+BJr3uMTmrTlkJLv8wDAUY8e+38Yoyyac8ztEED9DNr8aXIw9N18gg20UDjRueF3OGAp1gMFra
yWh9foUMvzb4oPM0dDC5KcPVklRCSthgRrS2j40gsIoKB+zyEJVbI0KHZZuJ8VsgsJ3RTHIgsAGt
nE8F7bopMR6siUUmMwc5meRuWEAuWvb6D4zDA/YaCLfjP/JrxQdOz4fRtSxoEPHpTNmDRrZcWT3T
gSqkivuM/qWjQRM0HnmEAubX5W1ecq97oyE9wJAs0Cj9skwwxmLuzbhP0+Dud5j9YZhi0nzxE60K
gBqrmhZlX3DRiPwDMlgNix8e08aknRgPyTPl9ccHVu9Kt57rHJ0l3q/4lDABg4fDyNOmv4NjzZv+
PmsVMhullFFdETg/g2aU+vc4FwP/yHj2ODgpJjhUlBTCL4xlqFpuq0ATvxf5tp1kMUbscRe5Q280
XZXELepf1GwQQTP4zFFoLeWU9VbOUM0Bz/P6QleQCKtNL+jQvHeU72XkHwtB3CYlbUCazSZSmwKm
lykxvMQz2lJK5wOQofGSWKuKRl5X1uB/ArMQw30hbhBdBtlxRpSe42kBHSDBnARVpExpz436ywic
HXL9Fhss/xVYgIPnbZLrD+bo7jAASskRNL8u8gLTy5C/7Ukt1Qmn8bQ7iTjst1Q8njhktp2Wee6e
FvzKAQ4oqjXtG/qOXpLcbG8IStiOsz6Xsgo+J05zr+JTdMGPBqRR7fAKROGwlcwV/lIK78vzTqdf
z1nGimwei1Gq6dItO80uGLkzEdoqPE8M/0FXZNM6mTJZ+WRfgRAk7n4cSWZA7qGztePiDacuoARP
SyIgfIgVpFsiXdLbB6tGEFxzrs6e7llJZqOUDN4Y+s3W9siFOxVVrKa1sKdCDC7m8qlT8L/NFecf
/zFcxQult9WCyiYXaj6oqHsi09dQFwU7gakhbQhQ+XUB0RversgdR3C/+enffc2Jg92JsyaMipS0
+5F2w0x8frQ44IgmyqMCsNlDe2grKOh/qRXHqQMH5fim6ldVzRbNKclVOrE1Gdd7NpI7ONF7JL28
M0DbeF3eFZKrDrvQOXAeWqc4WKlhPR9CNDXZ+4vPvJc9lom49PV6xuaR6ksojmqoVlP+gHIB3rhE
bIzRRuHvfdikztUCDFfN7TueugLd1K5oJHSZOsvtJwqoGn7uSuaLYRIfKoJaqPe1qYO+NfToZEWd
Ni5LYKwoh7IEfWm3afp4zoWZlBhW8JVEmIZXJnuqwDd//DrmM9aXv7bD2HZmU05E8QxX4CLqBhxM
Fa7lxGjVzQDol8xCwyjbBKnG8qd93fdcCphma4Af+7/3HEuGqAM9P+rBTKFvXtykOVwOpN+v4jgd
+15lPzAYhobUEBMNISi5tgdbmnbrD/YXJRUi6zQ8eIcyHIp/zwEQ38rsGhn3knSfVOZGNpeW7LA8
/BcAEh3GmuIu7AcAJX+GJZ68L4muyE9vJG3Ftnl0jV36cYtAK7VMlEZBKGjIz1WkXNRO3jkxIWSs
gpQJ2MBqM9TYWCRWFQfV9yjPiRmrOlo4aixq0v/7TweVSAd5UrDPwCSwUR/sNvIggusnaXNP9QO1
IkSbed3Stc5tJluvosTSQnfBTjdCUEEYjzIZiHy2KzEF1m99ukFKBQTc0XdoKLuRyilYzBypWLVB
GB7SsF9A1azitjiPmyVnqPSa3C7cgUwOnTTSbF4+552/953ZYXdUP/Y4NPogi7L6DZB9qK6rdSaX
/uXc1kUDgcVnoDMDf4hL7pzjHaxNbiKDxpDuHz/4Gc1WoeLBasbG+oePn4j+dmm/tjzdrF9TFHUJ
B74j+iF48dZnzVv3FXSOvLpTUtBX36FilosuYse/W0cYFCeGvJH0175NANGIIjuBUAszKWWjq96n
RgqPe9zrPjWApTnYNYt6cSiwH0kkpp/LxaLo8wT9yF+Sa/qy8ifaPed/GKOGUyfSPDmxdeP3L+1g
Yw93g08xhhx3/i0vsSVKKWMDaHKg4qj9H+7PKUyd5O7RQxCdGhFuwHa5SL/zqJ8VSIbJKUefrVtt
5KwkAIJAwyN/THGqaE6gcDjM6MiyJsImcb1zOE+IGqPqSzDuTFd1fJ/BOBJ7SWrwtiFzZD9/cRho
JnSu7hCbVd/kmwmCnR22pud9WcNG3eLuymTwl+Del3elJX9K0iRZG2FkwePYHyjTwmJLQOpBGG6/
OCQBxi5JC1rpnNm4eWh84Po0kcJalrK5Zonxr2fcikWv5fxFtb/AGtd8C0y/jT4xs5dCxX8fXhx6
P9IUisKM1jwlIDMYCRx4oMbmjTRRPp/NtR00l1NoRdLZta+XKDlpkAOjB93uFHvuc6ohR/ELPvEx
fneZUR+kZ4S6sVIRw9sr/k4iwE9/hisJKFp/3t8G58OMqGVX9IoU3gSAN4mXdvD08VS+9ztI4+1f
4u9Q9ViLZmH7R09aHGLLwxIbDTfSFdLVXrBOVHppR7kKtRDHOoFCkKXbGkB9NFVlRw5qEM+XJnJg
3g4eME5vJrrtGKCa5awdjo7OeDg2FqHZE/dG5Bu4Y94M5o8o6R4/jkEgVkO+XRct2zjmCIdsd36w
GeGG2oprB6sTeSmxYkqLmSg9T7OEj37XQNGp+wrVV3e5iYjzlIiHFjmoORK/VpdkSdAqGCUSXphx
/JW+EgwQNqVEE7J5oDEK+comw94YsSJHdNvpFUiDXhxGpCGVdFR5SzvMqQtCWUBujOO+7Uk7MYO9
oKHPZuzU26t+fyXWZFD4WqrzRth7utxa85dkMRI3A0C1lQQgdAr4u2EAEPZ87CgN391za+Om/Bfn
+fokzNlRtkk6eu34/4x8ZggbdTRF4ShZ99TkTSBtS607yYbR0i2aRpFFrUXSWI9+zOq2i/IghfdN
FUwRHS60rdClBtZmhddj7azB1VFg3QYdNpl3ef5CdjalfPeZGiCcpG69B04XGM5t2G85UpP+q0gB
07q7zILlJcbgA7vpvGgT48Wptd1lg1GCeGSTF7TgDgkkg7n/UEEpUTJ8EGGb0ayPU8sQTSkbDahv
KfQ44/Flg9lfoFonnh6N7wvy3RcwhlZw+3nR8CbGVYOcRHuu/CH64P4Z5G34nJAlRGnfqpC0v2OR
rqBLzV2EPrGuHsuz6/AnmxhK3TX5qEjE7TCnwlOWF7KEBDTQ9mhc16dTxsaczBCfkBeXBcqNNLqj
Hr/P79GB5IOov2L4ezpNzcgYkOF4OCgUdyKR6RwquUVPt0S5wP6IJ9cSL4EZ5FJOExnuGhE9aLg1
xxAg8YeGWhGui788aolAG0/6eESgUCJVmI2RN9ZEHpPfVbvKCSmVMUlaa3Up+atBXifjNpS+grI7
HpVUvTWUgpiS2dvSMmowgiv38U1Ae1iFNXsgY0LcGA1WIV1pAHOd6nIOr3y6Wcr6Jzq3MyZsCh/n
MiQVGF2X25LZ6/Rr5fnXNTRKzWBdeFkZYRwh4pLiGkaqHOsK3HDNIg7ZsVO5XhBkQPxPSy3E/Uyo
ANHj/xW9bMOVNdZeA/Ngwg6c15ZqnIGXWo5TTblDHzVIXiOCSmU4fcAtEpJs7nBdiGGIWOkZpk1r
5dmqJb+7n8/AQT1UDTodmfHEmPt+qF+IQ2d5CLVPXOq8PRMbPk6SpT3ebvtRoBr7JTo1jSdFII0t
PtzXjzPJoDO/XTA2D1EMo4br7LsYfIkm8CjhcVHv8GuVcxFptBgPpyErzR5Pa+swoAcD5Hdqv1Cs
qaNwzHa3tvdVTRPl7C9ugpLjrOAf1jIu6JayunMiTwtYN7r9dLpnFgfrMRLHjTgwFkC6qcwqH54y
zVYZVtleg5lv+H2QL1ueLzq/LpRMbHLAkk/ThwGtKsqn0AnZATRgzsjI8+1hJDg2ZqpGfZ0AE/UL
iKJj5HUlno6X57JKOWM+h+douknQGDpmKFBxxkggihYcv8OXGJn2/Ee5y8S+wElgbrObMJ8lTRL1
NSSyp5kQul06f8j6NRziG/U1M7OIjQL7tQoB1wrEp65SZZAqZ9rfdWuN/0CgmctpIBdC5HtEZGj2
ZMv2rtcYQkulWAN8UGbV28eVvmihPFLv/bRzv9xuNgpxPifD0xopX/Jx7E81SiucozPH9BMstqHn
J02P6Th8bgpd9NG+x1PQX/ZHLBNAPkmBP47V3xHw8lHEBj6JVr4OBKQT7EC+I0+MQ/m8JBlfCdah
z4I7oiwp1cN3vrAcwNlIm1SjDjkF8KBhzZO/2WR1ndUw+TQrsYmc/xY6M63BCakR1fbEVDKmOVh5
mZPSHdQEwjl5knzRmitfkd74OGu+rvvqTPd4GtV582bV0tARXcbfZcWAp35dLLuql70GBHR7zUGv
69PS44dXB4Sq2ZAMRPcmeBVTWks46LKzfxUkOCla0Q47yd+OHlg6lOmN8AfjII0E6tKxgJ8Q7svw
E2TjlXhu58Kg5xIWpfC6XUV2AN6XrQh24zQtcpGZKTyMo+OFbEEdzmKxmY1ciqQ8rhDe5XQRhCF5
H9sp+AqqkiVlJZxqMBwSlU3ruFZ/AmC82se3VzEmvonThYy53yLA4K0rTgroQU2fYzuremZ61F52
dmP3XXsBN+dQBQ1wkc0KSs6OvLb1qf2/9PeC9qjxt6T71RYPbhXIWc5s0C8pIJSnUtzPlUje8dGs
wFtWu6yXK6WOwgCF0YcR9emynb61oebDFAo+smpjCT9UJZGAObkzBdNCaH4ubRaNy0LjuwfJPRTH
+PUzBTNKi9cQqpDgkxX4VBw2ZwWrz16pnyqxpb8d4e8/PVFVc7Kmc7C4/35S1iQjoPMmAx7osKxK
ja0vS9eEkDtfTyaxeBsDSP2tOOZigt3SGmoB8auFNOkQEd6zZDsaP9TqSEE5jIaNVD5GD2n9PISw
6/EWEvTVz7Q8b+ZOThCdFCPc59Zz5NYb+pkrSQbqs36ewu85EEwxrHWT1EyaAS+zkuKCcw5BhjRc
VbqOL8akLogXFl8P65YF1sqs+S8JOXJMVtQvb5AeupJOwuugCcK7dqV51S/NlBKEnkjnelmf9fOs
UnYo1aR85yk/M2dRSSvdJnupFWjxg9h6rr6KsyfLpmxAXHW3t5gRB2+0KaT6WSwkNcWX5lUvidlx
QIE372JAs/TPGSGFD+eZ24DbWgUodHQH9Hv8CEYkFuSddMF2QuNsmdOOpuRJamL9ELZSLtFN/YPa
0HicQ4paBKFtEk//Iy1w+cDOSSJdSsqcHja1MHEo9fMO7MWqfUIdzKtRocfma81q7HWHGFrzazOL
Fabxm91swsD3phJVoCkVHsZCYfIzP54wnnWBIBgvdrkHhjXka9zsN6YcXgwg0N10Q6aevXzOi9y6
+TmJNcrU3uyZq9Yjp1Wp8ko9IfPIpBEwFhozYSFwLYnTtVTONCpv/AlcANRQqe+bOET4DeRXIZI9
U6OVLQIoQ720ZjCP7pVHpSOZsatJwm5J8XkLujIR3lwWQ+f9tx48YjOHKaqQJ/7wiGwSgBbshkQ7
fJQTCylT7//breuG36k2BEIMVxgC54B3caq6QWGZSzbvSlndog6NV0dZNhCJDJEI/8pMAP3k5VPX
WX3HlAvUwtjR1AQez27dhR+4JjeMGWKHdikZl1LBNaGIc6CyDmI6VAvzMtlcTM5bOWUuVLRwGKpd
Ho6Ja50IvfhlzddlMYd245iOgfBIMF8TALqkDNOACjB9A9pgmJfU4K0in5lh6mgk7ovOSmapnhU9
EGDKqNdQzzg/J9m+C6yLAzkRKT3fzaFZ2IwrAKXDwJTh+VmgQdUSJJ2Jwr+vgQdPz1uZXsbopNKc
+PBDpPHAHsbUeAkC0l4YDYFivuo0VZAT0TQqaSCxUbcCIjVL/C8Up+UGQEV06JxwqFJO8xsek4Aw
BN7NpLpAbJpPChCX5Eqqt18rW0pvbPuGFVn9zfHAX+izodOULpaTM1+OE6ujoBJHDk3SSc8P22Bp
uT6BxUiuo07TMJ0B5LUFrGEMDgnoMMzY6qzfvzssowSqm3LwSWg8/cMSm4q4ocFZJV1bIdWofV/M
xiF8ZZHQwwMzLxmiIvMB1DbkHlk3STwJfO/QxDe9gPXBH/7ss67TFk2hDH1Rzk4w4jfG4MpMNVma
fG9MXZL1QQWhnq4Ib+SfO/xovFuj32p7LykavXcnBDnZNL/GGlF/iXTsw/fEmm79XWoCX748Cyed
h6ZU4+Rap1q99fvL9cT60S6eufdUN26Y0F5wzLr05Cg76yqyE3Xq9QjWPXjCo83G0FX3GBmbElad
Yx5Y2BCRRpenMiuEnqCLl0aBjUAaufbb8qUNXIjj0CIpCpvueiDKZpHdkIibzUjGH+gwj5krupfc
B3tlRQjlLTdzLKOlkhqTC6puafErChH5NSgBe98lXh21KvujI5h1joAZW+kKpZXkTcsuemUnZwRV
E7dyNv8z6+rFG/q74znSSiimbh/zZF+SWBlWPbPnV2/QRtZvDFPAXqXAMi21aqWpSQlBy5yvMNKk
ZcdAWtEmvUUuwwUbIHplEkAsDKButTtkZA1hUf7stTjoG1MNkPRgAAjXqGPJqAqYarJJQ1bToI6Y
d+RXVQJfUwML2ikak8vCqX9h68pOyMeG+FTK/hQg0SXdvKhUACu3MHMuPgY8dlDhibH35uiNbtjJ
4r1bZYCQ6WZ7sZDGW5apd+Wlz5gCicUxWkjdr+Rfdhk2IDgoYtG4gw2W84IJ+7pGOquhwhSJCUDY
8yUexzFlnqM0+wgFVXEoMblSlt+DGkJfbbJS7hXFC3tdBVvjbLWpnyi1/9l9lVo8sh8SFcpjb4Yj
+bcjIldWMamG3xuN0tzjyM2vA0j/3r2+Mvx5zvc4t2PPrzeBOk9Xhmc8miypVuXAvWn3dIL/JDjt
OExzUi9A3lSldztc3XKCoPc2p0eGFjJp4mVsnxl5WA7FK7LX0wrkKow/y/o6D6NuQGKcB8JdNfEj
UI2vxpaK9+EtWhMUaL4Uv6YBuWc7A965fH4yXJLBIKHGBkCyzNTU/aG1hjMsQ7fLzhoRnk2C5PiK
ZmX5tP7wumuszmp2Mylwx4/pb7NvHwLuB/D+qK6dnVKSeZqQC9MYhp5VFVk1lf6ioo/amMKebaFr
51t8ligxnMGNnWZlK4ah3ps/Xhf4hyJrisrrsu2Z5RNswsjbC4oy3AfY0mSQZcQmSTNWYNO3AFXE
oYKWUnTm7HLcnKU5lkZ+NudJuue6encpzs2PyahIwHa3HVrCEinMfM5y2NUyE5exMRxnGXWbbsU1
MtmFaaoz/7XLv9eijElytmnbeEv6llMLBoJAznGbU0sqwpM7lMhTNAWBepClKUya5/Tbkq8Z0SHM
jJ0ndpQoxAsSkbymkPlD7psJfskhC2AMeX2cP+d55WrANv+1Kaks7OYEj7ImAgWVp+GFzrU/j7QY
JjuewHrAE0C+P9M/0de+NYwXx4+yUJBAnwtCqlhc9G9tdvrjCKQALQi34oQEes52OW9G+Gj7aTg0
+1MSlWUVUIoY3Yb5NqKohUrGryHtnvsvLbaDevxTb8xzB6BCL/Xwj+bNXTHar6WP3IiT8OdPQbFz
9tRGrX/uK1h5hlljhuDF3Yua5CNhdER0RebPZ5AgdMEryUinNU66kadKnZCSjbYVrMJ21RfkRGKl
RQ6h6jBNh0+2o8dD7LHg7Ay+T4v1y4tFhl3Yrg8M1tuqY/+XsLadXvcZUHZ10PEfhLWACQXh7FDc
xcF4rFJ5MbHfypfKJqAIc7+5I1BKxCzF65FawAfiVrYLbnvcUx98fzdr6wcnk1YwJ5CH5OjhzW4f
bG4d3TGLH1AoBaTg6DYczCLlP+yQ5/EayFpjNATRcNQyvfpp58U8ppYAvWjsyIzXQWWFsQV9zk3y
JZaDdDnHPuDI6290BzYPD6XZZkOpCR5Ys8QYKfl0iB0ie3R7qb1NshBDkrY6FjMzmxU5sniobcFy
xGGHHfFz9NHyQXG8jgg3x0DRkWIsfOAs4TVhiSl4gM4Alg3bB+gyVdTRY0UR2Zfvj/UfY6CIGxKZ
301dfk8JDkwyTiR3Ox8f4DNR7HUg3s9S9d0xzioFk7dKyb2cSW8v+qIG8eEoKCfO0RNUGYbr+0iI
4Pvx1cJBFKXmnZMbnB27Kq/QcG0hbuZQebLTx41WjOENuhyDT0x+yTbicWcdFQ6z+7xpQcgLCDuC
cVVykrW1m8GFBE/oNF0jCFBxAx3MgTQGZwvJE7HoGFZ9WGenrb/FN54vXpCk/Vy7huAkFitdwUuN
KCtxafeqY0O7PdT2UVlfw0WnJUI2gcef20dgIfKuKZkFe3xC+QoPrVFAAFNxkLtTrKqn6hUAzbS1
YyA1q8tekGyEyCD76KUiVYYK2wEnooRRP+oLTdfzXrmAcFM0rUaFoiUdbUF6aZXGWZa8H4vJJ27R
6pvywAjU4wyfSekFgRvG28SzgT+T3lKKQBZzNkZcW2NwjX16SBfYeKxgyq2O6eqEw2ORh1Z+Y38S
sKa7ZMDBeO9QldhdwCUHPf6IC0EBysCk6Be11SO1UaDNcg/rbtgzfJfGjapGssq+FFxra1aJ+mKn
nYBOPAWXv2e2pbzFkR/R7nAPrg+gJMbC0Boeg7mmOCMmuRhgz9+mV5VBOstWiPTYBvodeaZku6xz
wEvgFhkweW2IVHq4XdjAaZmf/5jQYH0T7rC9yM63o1th+GItRyw2kNdlxYH3vGaKEdvhLqewr/pZ
iUPlv4j8df5i5Vmr5V8nt66BPhpCoSg5CjcWIn5ZMIKqzeHy63bY2GLy1ZxeuSaQTXiM1PNwMYsW
wDeUqQZ75Uu4WBmPSbQ6LKRBm9RZTYf2Lzeown7WbdGM7AFxgZSVCOR5/K6iWnL1ozIY22Slje2K
tDjsl2qDGnVALcZHia7rtBosg/lwMP3yyTSr9Nd+toDpjHUD6ko58tSFEW3Nb/uvfmIcgEQLQIES
GC1hNrqe8mdb0oVcHpmPUop/PhiacKivfPKoPR+ar7hKAoPlRGfgsVSSVbGPyCg+M1FmDVnDEpzD
Nhv0Jcr+xnFzKq+PsZBlySrffb9FRp4M7aMuYWde8M6yO6nYjxwtqqMmxkjSNgAeYZ8A4BnGekXS
p2b0hJLpE4ACfvgEFs+g7kv2z49qztHRXd4DUCshjDf3oa9DgnMlXZGY2kM9b2KnE47PjEj34wIs
iautYDsxFfsjF+lass/RYZxIu5iK18Lb+Qip4oBX0MwxFsp4Y4WVLLgujsm9C3EModLkPGkW5pjz
VGBBkOBtFjqZDZ2HP5JJebx+390DSqizAjlHgJzegRtMIjVoEV+A1UjOfVRsw1S4QWpKNl6bCSFN
8JG7oC2VmQix2GfhC1Fje8/6LRZgVcw7xA1I8WJ+osFgWdJiWRDJbAc612471AyZzVGHS+H61xjp
z8QUQaxj1hKB18lGSPbgdn6T+IN6JFwSNNlQXh7HiZndfV1/6ZCZj7PXWkngdAsQ3WPhI+CIBWwg
US0WL7h3K2n+YUYoBhg4CCu0hD10L/fCEIYG7e4VhFd+8OWCpIwKNdbyLGu65kFAzci+xAMYhmz8
9gZzEn+0yhr59QmrgU946OS9jaJxNJjA6EN2bYIcB/AH0PvjupyKE1RATA5g8afUu3AYWMp6J6C7
yvk+zRjXU3FCti3rwEf52yCLekTOW5ygxmW4P+wnZZtkdgUoq0WllQWBFG+yLe0PgwOAWtrN7P3L
at67oDUbM0FiO5K9QZlJekUucqpzG3ZrykHlaUP2oSYkGwk9jbWMZt6jcAOJVcsjOrrzI0sQtOE7
+OcLR5fS5FPtrM79jYV8s6KiIDZ4gL4RvcXVD6n62cEmVXN9LQr+OiwGzINaNvqCBAjDYWphduqH
7JCHq1HMHfTXkp10FKiJ1mwFWFAE+kXx0ACVAa+nrPgR6w+uav003VtAl02HPzzV+tDathDw4Vxx
RgBm0NpVbpR4/kKSXMChHjUsACgBKtc34vheuQytym+EYZitffs0rSEpSN8DBPByp5WT9MQVSFDD
3zDyB6ECsSZgPg0CUEURi4Lffo+dyGEzwlBge2nBWqOFCPre9+EnpjnYqBzDErg/FOc7tzwBqd7g
8PfB+nqcK16rCLUHBwbSQcR7NSGOYegv8BhF10k+Jzpk+tw3RB+YXEKIlBJmyjlQgI57XDWRDCx5
OppxKtn18CYW8UX4wWHxAr+aIyLRTmKDr6rjpU5AOuGoQ6wJ1VHKoAdUXA8KtDpw4A6RsRZDX+t0
fRlHq0NwwLwgr2lOt4h+MJh/w9WZwjITi0mVTz89yuJRpL/v516Fh6sZgA29RwTm+G5sEYK9Y0dC
ICgMzS/pxYy4X7VKL5gXlt1ktJ+vO2+NXzLgUdhNozpYZcVwh4K1Uq4bgLcBuy++qsYf5G9qJU3p
Ear724OUeN2ApAzL2/Q9Do/jrbgF7trZK+HzMOKFeNSeIyJ+e/vv+ieacm8aoz/CsbREWCb22kkC
grX45x+1Vu7gsmWG+nM0569GpFpynB7p9WpNOMA+jnR0c+POY7fyOmg4gTxL0pRmK3BVKWOak1Mh
4z62fVCJtoILteA9u8jok0ZT/ba/m5WZYYjlw5gAZ+egaUdU+hT1WcE3cHR1a41VyusuECWbvGZc
I68dQbZiJA7e36qzbyl2QHytm0843k5hkDI28EFHCYdJ3XX24d+j+NAJ3yzdEqDnfh/ow0xayU5o
5qMiwqG+/wqvv4D/tjA67YaCxbcawyknVEPahCTtq8Vt1t41kJkGZC+yVKvTRLoPmV7jGl54L5H7
3LeoDm5dRH7eBh/E1XHiV5lOQLlu/w9hJ9NGaw7w96xsVHM4z6WUKcy1rw3iQSD4S7MHhFMM6UmW
UzGIvzGb5mq1q2XB/Rl6PO0rGH/YdM15tMfhCtUo/ZpVLBr4HSOqwP5ljkzOeiA0TgJpZBRBgrY3
LRfcFW2KrzmUDMAedpPau24rihvKQNAPIA4WrXVwtfQAFftqGNEnD2MV3uJmWjAFBdhxfTzVRtY7
Xkzx/KQn3ubzwckXO3JoQNvCLchX0ePOZzIDyb0Wjl51Y214suO9sEmEkkRC55w9MKP9pp8vGWTt
jwwcOGA1g1Lsquy3syogGkjs9LS963wZI1/odCcNt3kwqvBf9iSIlIr4Sz9E6GY8jexuyoVbzw6+
knbdHfqdud9N/5LtQp9L6O4yxY+9ACPRU017YlP1JUvVYrqlPmQ4yAGms5+vX3mlRIOmlY0mnpTz
H+utR0gKMqFbJnh7MrQtj1UbjX3rNXcZgmv92nzMAs1tfnXZNKOVFoBsNXlhpQvVERWqWJVvHwXM
NeSYv9ofkKkqbaVNMP0QWCb3tc5jcfuiclXQURnMBG9B+Hwjp0rxl29K2DvM6WgOhf6ROyjAk9oC
r8zWIVmmylzibT731KppBtGfNfzBnpTQyC310qLCwSEvPosqKlVY+zEgUk+KUwnM9QuJRcXVjhGY
cJ5QBiiae7sSv05QHz9zsLVdt8Y4Lffh5Yx53iMq1biws0AwAw4ZexuOxoc2HCI3mLJ74fJQ0u1q
ypVMvQucuK9uRGT59PK9mESIIx/YrqB12tzJeFmbIp+Ou7k607nbBORphnr+jNKsyKWfwb2850Mq
1CiTAnuc8bmX+DMStuUQU6It4lIRkGFTjxdwtcZcrjM3gyWyBkfZKSHacIR0mBeTnCbri6Do8Rhh
DjFWskGvpF5Zn9wYDaPPcEtfPKA4lTGnLOsvXnys0HtxOZp8UZsvkGeAHZDZ9Xcx/EzKgg6JRN3b
rsoNx9E+zuHl124UcbV3pDqyY8J1tZMMlR6kF4Wp6cvcynLRGlUGOAPGlZvrPX4ueXvUHrB5DV4I
wwDZlNe3rt0gBgb2dsU1Aw6gNiLZKv27CqY3tT6KOGDQI+V+tKhk3ueavxvJZ7bz//4B9hYI/R2A
cdeJ5QmFZezqvr/gQ+iFBBG+tO86RvmOTnvwkkCVObrrJZQffJ/XdqtoF+j4QKXwgZSnKA5pUnAB
zs0y/2Wdk+o7jPu7zERTEBikn0aP4vrf/jRpMhclzLS1qLVmBagRuCjTz1JfDZ+PyuQF+jf/69tp
x84kIu09Bgp1IitOSfYpGAHldzkqk5aWWCx5p/NflX88x3tZD1/Jag0SQlvMXVVwXnvhzPrwfrhT
16A8/+nTg+AtHYfTaIXt/Ea/Acp/g7GQzMn90SgE9sbBEealJqPdSCgCYB206g2L2Y7i5/zY4Ol4
c2K44oL2Jv6CSg87BNI3mx066jFFVtYH/mAxP0VKzuv58iUulICd7KHz6EFfC/24InlJE++EEEHD
UR80n1mRU1sQZYvNp7Yq1jivBQbk4Kl6LLIF7B+ImZiueyFV6IdC1mcxvUvfs5sNRH/AKPdFlNmY
4t2+/GH1/lyTfyKUMgJvGZlE0KTx4YZ1OZzM0GxMWmQkpv9d0Cg15o8uRRMIcrb1D+DN8JXmKv/j
v2egRMTr8qgZ3vcLmnSMJMeybeDAItqReA/RH0Sr930tkbvdHhMwVMIEIzhL48rC66DvkFMNtMjZ
JUEqvDT+EGrN7PB5QvYUpII+7Z5cP9gq3c5ZbmR3lh8jNnlPscsTyp6gdGn7QFp0bvyVDZMMlZKi
mIxJNLg6NxS8QnSCMFtmpqw6iM/sVVy9RlZxH2xqg8dZ3+dwsji2ULJNP4Nx9kqLlupp+NZ0WLYJ
2lymBqtRE/74DVtXvq8nRdptOzTN3MLeUaJJqNmrieDsXCuelU+0+kJUnP4nbRpKwLsUQaDCajs8
uuUKcauJMDGbtWEPjwbdyxbGynl5z3ekX+vrcdj8m+NHYLYN/4ErCEMBJISwAFkNzRzXRzWL9toT
1ZxSsEXpttC50uwayEfndZt/dkr96CXsiAPOpdjclMky+7/rNkcf7H2ZnTykbUIGuc0ELSY3RMy/
j9jd5ZgkIPOMNgs86EocYnQrsT/pyn/BG8w3FH+KKc+g0e+B7KspxnKck+t5PNlQByWT1e6cjJuS
0l8e9dDyGd2SAKWkAdeVNiefD0ACFiisuVbJLn6grg/ytSWlxe30SdbrKatFuUbkEIoznDmrPze0
hFsRAdw+hrbYztDNntWnyIlcNlcjmsRWttf8Gr0WqIWCopF0ivupQwv+3WYrldKiPzKRj3XiqdvW
G8PbMIx0YsXt1XmicezVWKIfhltlv6FJJ2xl21FjYnPBCgk1kde4atRM9WThpEWqDiYgaXui5y99
wkujhkhblI3u8j1jwVn1vIKnqojVppRkGDllwQrsTGDjLiZ2jP0RO85C3DBxY3zMK1/kneJLts9/
BB8AoIwYAZaKeaIgeC8opNlHKVEh8yOR5oNms+lZZOmPODF7j53fNPR6J6PB+TuHJrxBrnZXEi4J
E4unsyjnxYzWMsUz7kDp7lO/Q/o59AROOkO8f8N1OX7BZlHCU/Jjz5uqfkS369yQV5NVsLY81jkY
DRl/OinoYAk68+QJdzNAep7yRvNyyTa+o+YqSr61k99HiHPY1nsNT3T5uLJmmRc1tCMZfCbwSsTu
S8DOarhZ9YGcjhDq1f8lAHJAOyFYMGA0/J2HhO4+lHlWQc03H3ZDVc6fUGfcRyMK7O6XBLWIkLXw
flXOy/rv7VF6vF5+7FnsZDCZJIS6h0tne5+G47RkIG95//SQRuoV2HRhIH5mCRcT62OCXjkRzX37
Mvy7GqOO3Bt6CZ3Mfv+aMnaoZwWAIOOy6tDSwNX9i08It3pMMom/RjlET39w9TWIRiVfGvdBkJFz
xpKxyBLbrdtYuMk7r/EQ2sOo/SV5nIU9z5hXsYUb5KUN8hVFGQftqK+NzjOq6Y+ibFhmMMvR2H/k
5Afz9ewbayXIKkYqcM8p6n9ZUYOPbpsUqgFLCBL4PSa2hyYcU0cCMJ5VC8EdJ79r1CdPOZHGLOQ+
QvqLy3RDnwFk99wqNW9AMVckQrlP2IjOeZ79oJFRMjBpjx6/il/WImlyYdj8SQD9B081cbcvHMme
2XKtGFJZE5T1nS8Gm50vT9eixeA3t/ykYE/Ixj/XTEUnsD/vHIfDI4V/atEkwvySAlvrggD1Js5x
tuQg7tqzEmX9wVuAOA/oz8LnAGfP30ba/lybnG7g/ayZuPfLh5w4MMAO3pbO26EEFy1u7CbmBOXf
Sf3hLOLqX+gC3IaudYXIL8WRqh7BPBLPVi5Zy8xSWXP7v0Gt+PVpFHbTyzoHODZhPEeHqTPWVpqj
MIfOXV+mFfNoTEeAvBj90fI09+TD7WZlMwNq1ZWozRi8r07WQac7OcaFNhGEmLS6L2eBM5MrKddw
Idz/+EvkAOT3UEEY4UXmwb1oJUQUcQpifAWWnIPwJjFhmAf7PYPoQUswZQbQgymlohqM6T1fff6D
ADF8QORuwVmYrFyHaYQcIv8H1LDJZpFskXG0YTjRVQSV5JPgnztf3Ja+9GmTQQkUuVjiOAa9UHqx
MMlUd/+9zALcELoV1blq7LQ2t5RC+l0qPEjbVRpgPfQ+hMnnVUwazD+eSgbrKwhc+UIX3E7sdahP
r7R/gU/n28dc4Z7avsZYhPo1q+s2n2OOKxYI4D56js6UPdlywNythnI0DZrXSNhyVUWMJ9CGIZwS
e+S6K1HOS0vW+O8bpCzztvc4E79lX/M9MDUKeN352Jh539odf2Dbf7wPzd4bzHNLg5k3bFCreGW9
sovmDE2F5ZTecqNV4WIrXUqhufkjYsf4x34ItPQCFmWWywm/gzZhhNdPw30arb6KdMsnAm4FbyGK
9ESIDvxf9fyrfdFni0lAM/K1EbIby75dcI+KOLTK2yTHAxSb6tTZRcATqQ8W9HGpPgc1NMQtFE8S
zrqZp8uKJsvOHch+7EA5ZTIBsJaKxUNGOaXgtM/7kuZ5NgKhoycJg4PVsM8A3By/pWJa2kNIloNv
lhAufNhDD7sxSOlBKFP5h7KUOHZxS2SPfpd8GrRJkbVEJJFoLglagSVMpQYXfeA2Dik29/8pQgQe
eFiGDP6D5lEr3KQAlA5gWWKMulWCvDgR9yuTcumaqBPFvQ7FQ+ZaIUjNw0GfTxlsDDGjD9kRyFj5
dFcK7w5E4JK/SxgoxJuBF3qCmxuAfDiXqotkkE0/l+p4tEHGMJJx024i2OcUSzwES4EUqsBrhah+
fZ2024KvTpvh34EdxV9bnJ+W6mFBZd7gXokClzjZnC2q9jwSfSLVlHT4IHks75Gq/G1tMudZWwpf
wgu7jtgNxrGzViJ/sT3Sojk6nAl9oIkUuSiSoD6A1D99smNjJ+lo7lePPR/6ogl0EXdWP4H00YgK
4tYQx5aXMCys0dIvp61jqT8SlGLnSl+y40SCTFkq2aQD3FqXwqv3Z4E5FzygFjlwQGzE9JGeaGZm
LZ7W5qlerQxn7z4AVhxcFN5g/tyZXSNN0Psq1zGbqW8lGRysbw1JpDkuP5KZPVk/S2tjN4E+Jy5F
RPftX6GmMi0IAKhvAQZtOOe5qiE33ZRjG+lH9py+f/vSqygJVDh1Na6fKyzC+mPcVNJsCgFrZEjH
G1kXdn5A5pWIgrG7gzC2qUSNF/ELwpWHHoulWqmu4I/r0v89K9SK8pM/Dm4Py5SxXRzwz+8yB7xs
zzvxrLBT0HAqzLniA/bF8T+ghlpetNWgCTD0ljUZkoaeqGkhm9RG7nA1tVElT6JV2KdSXcGW0NkV
UcXDbD6roP2L1GBefMwCkarId9vYk7AQWs0y1KskSx9nZjNWCU9MS77ZKRwI1pY9CjZVuirospW2
39QL0AKGcdOJAUUOlL7xIl+BZXX6tvopwvY/Fkw8lsS5V+bmOKCdMnR0kxicaqOBzWfCjeRarbN4
bJ8wxsQ774bl4CQE0eYGovkFEwNe3IYrduHSshAhPzX93vd0F96HOv4Riz4Dr2py3Czrrk2+bI7U
83hdrvAZfrIypUeyfyTHbr9tXF5sCenw+mLNX4uBdXmr5YqrQLY8SGPSiHAsShgVsoHVDJB3O9oF
te9dWY8WFfBKcQ/tFM8SKX363+BfS3cSWmDweaK9tbJXqfnVczJHtz/87YrRk1psBjunlT9o1ZZs
zcL9hxP3yjPmP7nalGYIkOKIxHdOo10dWkXAPj3OiZSj3nZnuq+T7raJUAObjKp2lYWRwBcN0Ph0
SY8VLwc26Kpi5HqZzYmbROXypamrCh3zaV8sZ5d02Rdh8PwStztEYGuw5W9rlg2/aZlmg9F7w1Q1
9Q3Emb2kci7rUxAvQCfdDiriyOWvm1ABmkkdI8YhDVjEGMIzRcxl+lY5/uRPWDlHNXq+1+AfJa9q
4dWV26f6l7e7vJaz5XI6UUKC3pcpnkwC4nmKYW51nCgFJTFazyBpu4TAwRrD/LdqQB92cw4ef9wZ
r8emCCb8bwmkVzghgzJHBZurRQJKJivG5CBvcUJeBH1hQQCEURrZ0HhO+78J3QpJ1Qi6lXvpWrJv
G3kwgfe0qLM+Rdx9iALVtbvWJ45cB4PHrjzbD2P7gWigMfhwVYEIUgqyJelWUv9XKDDb303qH+b1
idPW9yuNbQZcc4TEIE4hsTqtf7SnoDNrIjdz8Br8jfmvmWce9wHr4KmEtqT9gBrMv6YEjxT07iDw
79msGWR2DFHaTpgGLjPTmv/MciloPqnNjRmleOC6AlJ8ixK+XgT47+ut2PwashccMtXjxwYjIsoT
L2dAFkYM+Reoru7bU6qsWPt7BXpIhNwcIIcbjzwH8GxVtcPzPVmZNHX/Ibk64EWVLKDb2/+pNbg6
cuP/OfFQUAyyMtYIgq7cRC1q123XVCy0yeyf5EZEx9AJOVUXPJI6xFHu+Vw8l2FNM58IIP/oZHoL
CfW9ScZOw1qR85uQJv7Y+XtUJW7bBPslmJKxzGU9ypbh2AjNHyFmmsDw7Hk9gEgwoi5X8tXD1vS1
ZDJ2+n/KoAOOHnInmoyKOeuEl/YeCgGKU0jkVZmJiKmi+d5yT22/eDltImkBEjF51Fmj4ApygcCm
pNkiaqUUYn8pmPq3ssmM+UDiVVZ1j/fPkzd+eCnMMa4xUkvp9wSIU5TRNYc43C15nazqdOAJLZJg
sTf2IbAUQLEy58H8vb1JqRRvfWGoL/U0BjHT/W9tvu9IEIRBCm2+FD9JxKHgLwbIxCWxjhrBwY9A
Dq1WaHo7y8Xxaq6QMnZkvRZOnSI3TPHYQwVfBwHFbtcb7DmJXIewoPTyl/do+jOzorE1/rx2Ffgb
TYWf75nN+d/Fm1IM5KayIiP/COZdzpE08UoVnHqw70Hcbge6TLLffxX7NPYxsity36d6A4D/0NT8
NQNgF16sqAEajh0OmR9PisnXYT1otYB1uQpna/TxAFDuK5fUdvIguGx8JVudhq+2E81+CbtCB98U
SRcfQWEqkRf/kvw9idTARCLMk1IgYfpCU0ZFBhlvegKvOlzGgBzT8dywMvzyZYSJFXf5JBxLwfLB
1f0uoyQBIS7auokHHNS/4uwQld7G6XFu4O1Y1zQUU1WXmR0lJl2oBWJLe/Zco043NBxUjmv2zrEd
cTYz/q+WOIGupaHqEvXIxhx9Zul35iH49mPMVYOM2L7AbhM00tSotH1x4yRWphU8Kqy51yk+2pYd
YqF0+f+AEPZLTZi6uNuTEVjvfRhi8l830km2eWWgm1hnaE/RFPQVqC9HOOLct1fec1B4ArOgCYla
5fm6HmRFZEw29oI0wmVG28FDTF1oCJkQBwRqYh7e/CkoY21ehxPi31YvnMyLVA3YdB+Rczh6tB2t
aqBAJFokHNbPxFea0PJgtmTgVD4Tb6zcmw1ajExNrAcFIdIV8aexU6JWbgt2Dl/R9D6A2GjFXO0z
2zwgHJqC+EqFVCNOpbYZGIkKNcPlnnLTdEWTeMakVh+BeQqa/M+x2L7LEqvu6Sx9yL4BiJf0+ZoW
3mwl35qgtCUfl1sXdsaWNc5p9YbIQ47o0HS1jWrSTJNdEVFQSiaNzmEACC9Z8gFycvCRB9mKcx6B
174cFN+I3N2OUMqy/ycHa5ftpu12gb1V7zwkS4ZrDFhrCogoFMUIaPZwWeJt+tPwaN+WLScpwjHS
LAvVq8ECbV9mhFjshSpQU3niLfLlniYzcWbfcmKSfPn08o4a0vffDXrdsrcUlT1Q8Qft1NBR+0O9
1p8BUA9V1ETD8MR3My49HPy8iCg+UkPtD0JIeUWgj9Cb4t4jmLfx9vsBajh1iQOT0zbkwOXIa9Bc
gFyZrdUb6h1aCP+UZZrTS4RsMv9wL+AP0+CMJ+c/FfAJD7te3yh/26QZeNtVSShPlUYOXak2hrKa
aObWfFqDUAfiIStexAh9xqbKbyJyNkTdDqmjVi+vOuVlQ0S5i4caFOj3mXBnQjU/Ns9cR8D1t2ws
SxlElUkLzuY+31DSY9VmObQ7Gj9NQRbQxn2Re02RiciUVJyyedsi2E4z//Uv7ZH2mZB4Drgpgn/7
MeKsvVNDpdg7jYEx21R7zjDbANfu90rPnp5j372/L6SXPpleXkdpBfgEJZkSLO8G2wMdF1E++lXP
o97nCN9jeeMPNMxy3PhUAVwmwb3mn/vx8eiNagdKuvKdotmrf4+s9jQ+XVhSBPDhqJ8uRLV0QMPZ
fSBRvbQygfcSAwiE0kETP9fI5UEV6VVv6MNuhhOT7b2hNkkS3aQi+jnF0wgT0qBE+H7RWTOM4Ihc
1HbjhrVIOhAJdM9Q+Q3ybGhLM3UQYE9W7Hi4F2bv/LuRYm/eOTwLPmFFRM+6wOBTthioxR4Gf2qi
lY5VYUk6WRb0gaHNBhP6dOUWYrru/jKYKkM6Wlczh/sIJICrQ3vayF6nQehMQKF1h+As8gjizY8s
Xz6HdYIRqf1rH3R8oeRR0bKQjPiNozHsFXn+gMJYfOodWJ9wSS8hQiB/C93hl3qlynJozLLl3s63
JpsK7ARzVHZhwA1O8yN+HxBpxfDWU7Bpuu2Tl7HaCdDiZvtR251F6dPuWseEayzG4GJcpuqi1sXW
gvEGsRfIGNO6rNekugebTz2p/3WGcXduVrep7wz0M94Hvs0s36rBhFRsDtj3CAcMF2xNWTjA4yt+
GjpMrTnMvJJmlc4u7I+VnFx5cNK0IZm0jC9PCsukqH08uaCuBHREWvayvzq57RR8+KlBgZ7WHmTM
hUY4z8LHbpeufGukEnzh+xoIhHrPqDOQVQheNYw3zMxmsF9Imi7pf1N6ESFsL/01QKyyoagJrpEQ
ky4YCFBSjUJs2gYs0/o7SxZHN0RFjag728bU6Xm3OeFx5FXaR7oIubNTUbxHMegTOF8nHfJDdWpc
SaVhciQNQ5XRyQkyxQUdjW7rPtIDNYSaWiKUTk3RoSFbxa9+NvpOEu99J1zTuCSxzDo7Wj59noqp
BG85U4iSV6lYxi5UoCGat+YCId9ztc/hvemOFqmvGlckgW1/8mg0XMcygwXz+F01TQ1c4T7yoTLx
QdqTLGubXZPguyIi0D7i50AVvt2Klqv5dOeU7t+PxU1uUN4wHJnJpzgH0tWrXHZF9BJNOahtN6FM
dMvwuFgGFrDf25FBSMfzcspXaI/3vOhEJAa5mAHqOaxrZH4p3MBb7Gj/6LmQPlzZStovnT5ytWy4
nJuBesM0GyQnlLxOSYAK76amMwSt4QlfAc3CH8nJTx4yfLtFlySjndKAD71Hs+4QgqZ30jpSVqa5
Lztkl+VVt1A4uOsb8xWllZnQq14xt2/qDzFAIyp3z07pqyQeQYy58dB+Cy2342N/HVwOEnnsKAs5
gx3sooPNII81Pv/WPEslng8tZWQuqSOa8rA9BH5fqI2CjE5AkJ+Q0BcLrjNU64OaSiMVBw3PTWxw
Mkb9cliudyAS5S3gl7PBOecL6yVPJ2SaNGRhzXqGXA3Kzcl54KQmiyU8p7HmUijP8SWQM6vm/Cz6
f1DYDLOhryWMqALYXTcuLnopDwyKyfvIqS9AA/7hI5962OeZ27hDZClFDUrjTPVVxYOHqrEKt5y2
YSIgmdBXz/0lkzeeQxRi043Dkc7gVc3BZHldjmxemF5uUZVn6FWPzkHFd+36JrUFliELTiV4xO+M
8/+OPExTIQ4o/0xTExqDLGdWrvhzshYQtueGVHist/Vrm28uMBZQXpLocT6TJKuU45k+uOOacsXZ
HVs1V7w/+16rBBHO5j/7fImHCjCoO4wIeBr++jm0kPkXKrW4ZAkbYuDuUwmi/YY2MoiZUS10GtFF
0zaSPqIxOpzuGbXwwP+UNY5l2rApajAEx0X95Sh9iwj7jkh1UaClAxrYik4aOYcpN5dF9mjJGnsn
JePu8dGIzKD1vXU8MM1Xcn0hrVIMBSLDe3gW3409L98F+9QBK7rMmxY87RE8EWuS1OO5zB94P37e
d1qWwng+YbogXa+N4hLI2EjyVth86oypW5echdPmO0/vGEHXIdZlF/rcQxCTaFUdQU8/e0TuGmG2
gc9Hz4YvgwdtTFkRW6FRHIX2eh1JzjdS3TnHSLEowUGEWFeHdiv1jlDKzACic9wXvuIr7HrKNkuc
A9vOZUjB9xL90v+mlDkD5NEnnRVR0683mG3g5Gic9EK8OxbxBMdQ36VGlXmWXQUhZdfQ9XO/0PjN
64HkQZyZFdXd4f52VcnOiDG3MO5O6BOcUaSbYQy42+x7mdf4KM1V+5uH3Wj+zI+ypBbBk9p9+1fR
Mun9bhNtL2VVlMifgypZYEpRhHSCRNIiuPv+aNHPn0gL+7F1GyQ/x7au8hIEMfmsY9Bj4PAuUwAT
evGKSQ7ejm5mhsk9HDwdAmH5ZuAVdm9M+Cfzjo1KkKQwahXhyDYGsqyQsOKzo6vFJYKnrOefztan
Lktkc+4j6q9cPFF9Pw5gSAKBlz27AEaTKRy1znDEy/BBrju0LCOUu7g+WGBuyj4jCf9mr1NOQTZz
eOKBhqcIjy9JeQ32uec0T77Fi2WPHxi3i/EI3ZNfn36nqWTRR4y3g8RMIYIj+YPTQlyqAgKrckYV
ocIhSgBFthYQsEmwtwS8jo6BTgnsDf8J3Ulee1b6+emP5oNrzzj4mxcDkiAoxzVPasszqkUugDkL
FA0RjN29Ohv8yTx7O5n967ZA8LQq4lJ7EQzARlToZeIGZVNg5pny/FtH+HNk3bAqMhrJQGY0gOzb
y6VCY6BoDHOL8tIosERbF2wmdirFJuWsQwYtyoWP9UDHQGU2PjPgQD2QCvYiLnMCoh0ZeoJEqMJo
CM+Xuheq3b0/HWNWErQw4MnpIlDgvOgxPhMLprgab2peUaGRQTAQa9RWRP5npJMgaU+KhI8zmQgx
RMta2lTBUx8krOs9uX0Hl99zkaLTA5L2wEwPm3Pz89Ezezy+g3MQbrkVdumI3L3nodkT+2mZ74bj
loKZ5KC/X0uAlzf1U4Nbomn7pXItgv0degKeQ3yqjonSyeLwKycGSr+qmUPXKv+72gH/6GddDiY3
omaEG3pDHizZqYakBlC+cSXZOC3RvJBK+AdePZK0rmJrZwmNLCG8E/vUHjUwCERTSEQpibapLlYc
whv6liQbdQybC3YHsIin6+EwN8HwzsDvtxiWdi+6+qARqaugdldQMy/+EUD0FTY9Gwz1+uQKumM8
K1m/Ri8SwT0aBV0v++SSUalodK8Rk5YnVeP8fpJqaOQ1uCuCCgBFDIb+n0uc8etGxkU3BbtlsPTW
0nYbr4Xo6KUQsrS5f1oJ8jyUjqOs+js0RXfXmU5rpu7eSfZe9FqjIynkWHYGCEbRAm/Jp2o5wDxy
mjaV3vyybqSJRmF3lOwVQXXRaFmjE/K6gSf3mVvQsz0irEdeRaR7YLamFfvWd26KqXe9uuixSyv6
BP7N6UduxRVbQVlEngOhcWkBU+erd+cSjU6UL+fbIQMdd1D4BNbWAA5ME/KVejzmFO8a5QmGJYC0
p+hHuEKXbqTFoz961MCsGs0LiDa/9+iXFFcWFV1l2AVamhFZS6AxW39Ifh1Zdo3Vs4ashyK63Ucl
6TLyUr6GioxmunLcrAqAgF7y2EqRlMBOIygsWbarKhpT+Wl//cCt4NXsX1gR6xg9DSF5G84fUANO
bhC2g5aKbBGpnBFCvu02vKZ5a1BCQa7XmisSNfttb7YWkg2do4TS7E9Qf07xoCn5lCikUi+ul/LB
LiQNLILyzCBYLWXkefhqZaUunkmFpZgBWbWrBLJSHf5mc4cmbBKlpUxe8DX8vIwr4ND2COCl1D19
1V1DYr3+3tPx6XbhKHh1cj8hiQ/hqopifdUmJH+QKUaI33Xh+9wkuEhWbvTyIbYlGFOa4iNrmyn8
wlOn8RxOMKPJoVj6mUcxPcrXi9HwCEoGkahxlQkIzfJI1IUMLch2hyoWp/D/UcEJDilT5SmG21aS
l+pTUz9xXirH9Ujgt9XILHhKz5/yZeV5xHKGq/N19CVToGZ9/Wzgk4fGxJAszFKAKGWarbbpR+B9
0N6rxI1+EGR4Mk/FQIcnjrfbJVaJ3zAVryGo4HQUVtVsFEC4R8baNLpcPgeXzm/n941//kfvEyhN
9YcssScLfRDaiFWNe+GSFyZ/6cWaeYIxDQiK7Of7h8hZnADA++9KjxLoaSMzzQRBNyoW57wnM0/H
f2B79z0j+nExAyD2Q+4x/rWK/FttcgLt5oWXXggNYqqPM5RyDEIhKtHac9SjhUmxL3gj2Y7pAqrS
K/gn9m6VhSCAvcCemxP5YS1bQJVA3W/18SDX5wcL1vmme4trnqhE7aiknCmrIjxRP4c7RF8B1aG4
oFHYAGw3xLUQi3GK0xwSqkbDy7Fm5FAs/9+fs67KASLAyxPsnwwVVytRvhKPErl8GblMnA/yXphu
zzeMbNzh+SLR3E89Lj5DYqHgascassukIhJ67x8+9cDkmMlNkRy8lPgr2DZdWVVxmUdL30GVI1Po
xSPa+U2ueteu+etxCHJ4gZHslM11znIf3djbh627+rOL3GUjw+c7ugtDD67KaDpVWOZdjN2hAZbG
UHWNParD/ioZrfej8WAmJSEGtVMV7Kx5LFCQqCKXh6AuB9BHwN+u9UOzjpghiCS6/GrrNv5Ta2Tb
8tf1+SUIuiK4bKu1zOZmga7wCCXi736RbUKcETinNNDqkhG1wRPC4ntwx18VzTLfP3EPBgg0Jb03
VZE0+PSKQej0zyVrzHnixeHGln9myvOcul4h6QWqakrXBTL4Yn5yq96+J/CFiKoOjKmTmfbeFf+W
cumg+4IR9N3k+jn3XLsWPYsQwgsrOo1t9qqwXv+SBw8t8mDasx+/0KCQitlyQcEr8upVNAWY/klo
uvLAMgQqPtvoc72Fz4PCJPHbalmNyrcJOXra4rS/TRO1wmmr+WsVRvCHMz3ff8ldK+85MXWcx4f6
GWMZUjrmovp1T1Ht2T8tMBfbbUzl6dIOanQbH1ULTjmnOqt75pwRDTpO37lNh1x94XwsTRmO5Y2o
cnQrAwk7iMcFP/p1Zo++ED9RSQIxxyD7sUZQpSVL4AiOyV60MWmNjto+JN1Md4ZjUYqTMs+EA3Em
9N/i81B/uWG7gX98SRN6ouGnSqbjSKLNXP2YpRj0Kx4Vhf/8w+oc60UoGPpoxT3E8nUwWZUxCpgb
XVttN36W58ZO6CZ+SIQKINWFQxn0z3LQorE+qQYVW3Yye03RJ5DSqpdpVpa23aChh1690FE9SSUx
+tvmv2JcLa0gVuM+1HHKnBWHtydB2yWmF3vtbPLg0IAhhx24HmFVmgVK1NrMNJYO5Gy/0iYNPSjV
yZgMWRVB5mFglo5/6nJbre03yFqjOstln3ovHfjl7mZlZnTNnZno47qiJlVk+VlJjIdhod3eTTcN
hQtOgc8kNNcU8nMaBPuwRAPHzrceykx8aBJX2fnin4dLZ9aC5oMzhh+QOHTb01/oJqgRaPt0jiSF
Eag8E8A8hupuruhRE+KdrauzHDv/IRVeGmcpgjN6wzxKJzCAofHxLd5fxfOvN5juhPOPIgLxorPD
C+zhBjft0lq0l+Q7pJxU8QR/fwj+Y7VxUuz1iVn1/5isOchZgSXHQPpb8VmM3Nlh3wzQBytG8sNh
SrSc5ed3CBMpqApGM1WHhhl5xGZMY7tqZLFDWMdpEOBjHI86mKulBAUWyG195EqMDwGKPy5PXNE0
ozyGrn+v4tSYKXRH3M3Rh6swioEnKrVeDL7va2HGK7LPTzA7j/PK3Uc4rgmyp995uVColEe1+54A
JXz7ChBUbqPD258UHjZTmLb3MiNJNQNxUah2OMpvl2SzhhA1vB5De3u66mlvGaytkb8p1csJXX69
GEjP0hHuQKnhTzNzkrxx7xswfSfGzKWmzajIns6dIEBlPAgCkuUl+9FqXR5FKjBKPPNHIZPdCt3d
80mgULtWWeYYJxaEgLPBJAt10oRVc/OYSIEylNh1PXPt2w564rIUZIRe0HbNpPMMyl3h00wfJRMP
AoidzsO4vdMBHwv4ZQZ8g9K8UDMqObFFO50TFPnTfcnRq2NDwkpx6cStF72F1hoo5QZd+IcZsaRA
lLDf0s6y4Q9HkW4FOcHPwcO6TKFfgf9YrrMVMDdYmDB23QA3q5IxiXH7p8uKMhYzS59VWhJZW7yE
O2LtLq812sNSWUdUhW+I8LdCzqUKrn3RSucuEWybk1jE6uoVs3Ok9SEehB4LmjxHjng9+CAQPVPt
xH3IQX9c4jwnX7a3Q0RN/ER67YN9I1no7Bk16yVp/yST/Rhh7ZyIUL8+GvVpN+yhJ2A5OvpdfIxs
Chb7tu5Xc3hCiWqag8HjU2+WBO7VrZu32unJOLQ8KCA/X14eftFMOYPmrereQwmkLbYv6SPHUEt7
ayUEoNhek/XNVh/Spkk/+otgWGtJx99aSnGH5K6Ejdt8NO/KUf1ggWB5DmA6N6CMd6Uydwk4VQ6k
20KE5M4JWGkfbJ/OVikenAeKtwu2C0Ew+Y+jp+Ew5wTwjPx524SFMoN/FZvWnkw94VmViY8hNFEv
BMmJutijyf+ilyriINNBHQT4crvzpBzgO8KJY/aJfTQW/0vbSaS9ZYbMGrRCWojwyGrB2MAuMmyj
/Hm8VYT68htwr+4NSEVQkfFsZ7awjeAaGO3OKpFaJyGJxYkseqGyofU7+Tj75tYgjpkjr1skonAy
FLElfnppm7Eyp2Dy/1xoItlfhn/X8G/CNPy3mFFcyvxn6KrtNMuV+ppwT/a99p2sqaa5keuhB57m
zwYLYfWCXCuCbz6pIdQCc7Osd5c0vzpWlm8DVlYFDHnJPYVRL7jSMhRaFPceWiiEiSGKNDUsit/U
YvKk+nJUgA7iou6/HFs/wxI3HHTXSb3jPUS0b0DouKX5cmdcDfK3HI2FVPz+eADvujIkN3LgJPwf
zfVrZvXKhqTq0QCeegmtel9dQjK1lZH/H73TdoNxhpig0p+NVyXRFuPE/gECcSeYEXo2EaoFWYW2
t44BSW+8+sy8ncefby84+DcXj4jGBs1GoMxknLasvXGFlYTlczVwfj0LmBM1EXk71DLQB1Djlk4O
iHOZgwNDmE6ewZqisi8C0L1RlTDUrpe4zlNMJoe5fAwfxP/9SPnfH44dd0/EBRostIbQEsA5zqzv
VLZLE+AlpmFizW6o9+2wyB0r6lqQaGbmmF4T1SMmwhBZNuDqCZGelL58xoBtlro+wp+UZngyWlwp
UgRyuyoL2+2b+O/3KmhOHQX2ppQKNCR58iBNj0JbF1148k7Nj3mFxsoZ1LE2YtwA+9mY6EmzXoQE
dbxr/dwuu/N1HJn0Uu/vGKLhtnQwWOYLsPWzX69INX402in9SnTWndyfk2QZ2epOfWWbkBi5SYej
P/232z3kcBGZEwKZvPMS99OQpeA/qbPUQmS135pj0+XxzFcEo15mpurFBk/QujkNDIg+MmwlQU81
3B0SmVduZ5iznEbXPhO29vIMIAaG6v4wcG5srWIsbMRoccCoUfaAU+IAn4YaCZJNISVZxqFyPMH0
K2wL7jLdcLZFyoWGcnYtbFJsZ60C4rjnrwheopm9vypSH22C39BZ5wFwg+bn8gYyib09Mhh1/xeX
GzkfzL9Srb4i8wWqL2YDq8XWJJHZ1Z6dQhtYFPB1j3+jRmnLY1FtpvbVe+Du2S0mXDT1UecgQr/7
t7RLFk6O1AIYtnVRnmH53VG+QEBUsuiRHa8XFtZV69TtzupiLMS/OwFBfXUHgbPYyAjG/a8xiXIr
gdw/Y3f7hS4uvc8GnDp9v4W0qEPKwKpC019TwS9qiRq8ccTILRmVJ7w/DegpXrEywaz1+ajpfbI3
+VTtqXIlT4IvbBQd108pS5x2Kwk5O5tIXCr1Q5w6BqTPcQdNMtlb0flZLkR2eMNjW7HIIW1sgwXK
Emv0+sb7DLCAjrsaoA0hX5SsltcNEh/+4rAmM8F5bPqohE/5JzILo8W0AJLA8jNnslhOORvt4Ids
nm1oZffuLnD++tV6ZNN/DRD4NygCYmhgqbfot5LUZLGHiKl7gg1JRRubnXDpkIpB3DJvUQfTzZ7Z
dyHvjotSuddSZ104HuyEvfPWK3VhbMKxxvngQ2HqhHtUHm2DgjW1VjKL9fJCsL0CS3YrVicP0CH9
Ms+D1sIZs5/9txD3LpaBj7cQcGd2y5Y6x8KDaJj2PR0YkxKfgEHatxpSOgeepJToGNMV4RzFxjf+
t1EDqGFlFxj7Iw4Ry93EMI+C2dQAecRpUN1vT+2OqcvjjSAFTOdVW0/uU4wy1cWxYPHlVQU/9/IP
ZQT3nUoa6C6fZ/W9um9M3gAgNEWzMMruvDRZUypvkowJM++9eV4cU7cFXKaUGsgC2ixhX5hARDyp
pRkUofSitjRfTzRT6L6xC0WC04J5pUg1fZEdJcNOQgEgPH4CXXnKnjUNot44iQrBMT3YYRPbI2BD
dw5ipwNoThSahRRSZTBTul0BvleadIfH1KWA05wiiwV1K/+A41v9H6r9r/+Y/DrD+qPfy0rDghuO
VwJ/j/E+v7wxMGZTOF92ymHHZv3f/Ut6LULfB5jMD2LHWIO0EDeCIc/HDWVpgL49cKv2q7GvPKBs
CJglVP8kMPAimUBwXvDht4uQ9/fZVKyO3IbMuntd8Y1KaUGwpV+UEjH1Z21g3Kx2Kli4upJ8PGtK
+Lsga/Isr7EcwY/p/KycdWzlHa4FbD4FCTOGDc+0iqhdbJG/NohWaYQBNC8BEzOXJrRnf3mdUzgF
w0jdt9idMX5Tq4B4VjeMy30hgElLBwL7X85XBvFYdTLsGjHKLCgWG35Cokw+94Ih7hH0sCmEM/oi
UOVbl/Mc2/rlBXOaR1broNbkOQvhJAg5KWBuHlZhS8VPIfm0MdVj0TUrM++63kAtn/xi/zH1qn/M
p4HpqaqEY9FtT4qjbpx3W6tl3DBHMph7sS6479Sh0evjbfK4bg3yo8upG62+dfFDykBH0zr+vidP
neAypcreXBbft/2BBqW7giUEbxrbxmEUVFVl4g/NG08aJco0ezYOkHkc/4Q3UPNsE2X2nZ4k+MQg
XkvzB3s3MdylIvj0+MIfhxAjC1MuJi2aczQnTsYKHLxFsawUTNv88MQGTxxNTK980trnwyJVCqtr
1TckjM1neydq5u+HIijrW2Zw+P8AMDW/DODR7dhKK967oUGUNWTHSIOnh3hu7PlwKcppjipXQoIT
SJhdKSds3AYjOqgQfctZLZ0lS8G8Ast7K3dLr1Nvyff7rLzRhfzva0bG7+WjPnqo7xkfZm5taAzu
w6Z5WhI5wkEb1D6FiHaMpu4e93MI/pSne+lrbbHHDTfwE/clkFwZisn/iaKks078BjOY45igi2sQ
vcGt0QnREfMuFkA95Ov/i6Xs+lxf1hKZ+hFCACpPuo/D9WVniXMqKBNzJTQeUOw8Zwt7Ciaffjwe
vooQBWX9OBPqJ+tBr8FuDzWoOPHnDwwQknIJCaSbokrn85iRV+2OMcSN8n0DyZxZH5B95FORduFa
XQpzifpEaGhMXI6VwyO7BBYo59XC/WzeZwS7UtL3F1wT36n8BQ8SijQdWqgztNNGQtLx0dWaAE1Z
ErjqaaCZaTsM5Se26mAt03joU6cI0vlRcxG2hRLRUiPWuzg5HlSbwMeX1s0Hsi7EIVC4ZtWY5FpW
TlDfWjcQnRjBksNgMAuz7DVohEBuir1CSL25/0ENyxl1O8+xewptNcIPP88IzE53uzkdhPnSToqf
7aTrsENAuyDhM/dDzG8A/+TClu4JX4TYIte1XJR6tRh9U8BjVOuKP4au6HusyN6Hmjld2048NRIW
jb1zRAzaey4m2u9t7oWXx66TuHKESld7ZNsN0UocWHJqdNTqBSXFFQ5td0Cvp0CWTg0gmHN3B/dj
yhdGIwx0hqr/6Uu8Y4WVg7k0fo8s73D7RoxExJFhLQ5tuCxoeGyHodgdd+c7slE/OI5nFbQRXddP
sTKv3egX0CKSJqzyc6g2u2ZRiPaD6C1Mrw+82y8EHNDYmPsCbWrVBZ6XVKOTc9FNcSJvDGOZv6uL
h7mSK5M+L8AE51tH4r4zpbDcYlOIvxLr51G9oTuQnmT0Y/JVAwYYWFe6vSrA/PicUP4dNZpQTvBG
g4J6ZBpNNAAnwfZxmXS9s89PCMzwNPyEgBP6M8IYOhvNlmeWwjwxbMJK25OZLHlMivwlzPcq01bi
iYEQ82W5l/cn0+DSvqvCNCtrJPpnFILfq4ruSIRClkeJzslTSK+MaG4+uNFroA4H0Ox19Qk5yY6y
C8PBlDCDnzp+Emy3DfxDpeRtnplgoKZ2NnNO6jpt7GAPqq8DFUDyQABbe8LJ6L3ShFQYxcqf+FIN
FPhlVt9Tvrd2QFF5d6CZPsshp1Wroe30S7HSZ9maG/mVvFcT5S9pUm3BelYP3szVlPBtyLXfbY66
yVMDuYoQVjdEfK4WviCQVajtafgfqfvrmF7gXcs0lT8+En2aURYwVgm7JjYF5iiRi75SArw5MH0A
wryIiUQ08jsA+XMm1MNlvsjFAqlfx6/UWrjzJJOI864xJmu+YyQOd/u/x96EbIkfiLFk5ogUIKbH
sJ9G/36k+5gqU7GdpycDd8LinpCmcY1t8SJpkp/Tr9H6UdtwfCkXTNpBnVoz4xOYgUCev7mqCzWg
Lb/efKqWFl2cc1YWV+xaB7qZw8GO+9T0Y4zWsbkx+GbB9M89tgBjlxcfIXp3BJz+hqdk+ooOL8nu
x5iD2DCBBzVteL22zn+nHORpYBHWMAyUQI8ouKPfEa5RGLACV2/hIEZFYoxdRhaSrp66xjVV++tu
YWVBXq+J6TkGBam+m4TUgRC739w3DHGhCu+bZTuTuJWn6nzvzoK0gJInwDR9N43NM3DxlNS7nTrL
crdwnQMvrr2QyB3758/cpNe6yXNhJtVPznj8WfFRy/oIQtJ+MyOg+sV7eafnK6HAPahOnQ2bjvNK
4zPEugSaVbptW0DDd97VeIJ2PoiMXXhQCMgXtsLM4xPgRTHgw+J5SQ9jg1IF0y0u5Q1DfdsxYHQb
9GqfyQ3jYewjxQtMwtClUpSdS3JSCn0p7Ktlzr6K2EcF4kuur32TPV7Q756lcUzv9ReJW/TkhqmF
qvLzoP7EoJJ2Wfoa95fizEyE7UzFsIH4rnbIMwA4Pa75tMKIHSLUle19m/MPU5lcwiB3dR5xJA+z
SHEpMaSu/1Eaf0SmZZ+7d/oG+aHpeSW/9OwLuLU229b9qO0qKRSpWBrff2ktkt9ilQJhaJ/3v8am
EaIrA0abGZkC73rjD3/Th0pXajDVHW41bRO1K2DlZzQ5Yz0z5P/CU1M5HASl1nhIQfrvY3DQK6yq
vTfmzKhNfPN8rqg9aA03aW99nHEB56BHf5wf+sJsIqwzUF1SzFmLhUTu1hxZtdp9/cxYOgAGDMdU
TIEFUxFNToeUkOxVfRoWD2vQeQuTd/skrwznS7oxih0bnH66tdSZtlMDnW2BIqdoHyCE1UpiSPLD
Rb+OWin1IqLrDO4g0TU2uAMvbxU/sY6UOynP8kDu4PpHnnFmVuvijdrraKfL91SpS2bosBLdASUC
L1X6wawX9LfaEdQRYBq+MEl6uL3YH/H7MTfT3AXaVSMyJh8iFHb3CiuLBjG0KrxEtv/CDFn5ocjn
yJNsaXfVe4cLe26mhHK7C+rBEAaDclJISPm6qoKgh2iqQP9pezEMsPRoegu4Lfj5xhPFRPfc3vF/
SxvTTTa7o2dQZuN0YZ/AFOtybTTRsqGx2aDE32d2IU4Tke9VMaG4bCsDMbbilk3vmGwUCjZSH8v+
u3TDQW0E72yE5f2zCzefuHwOMi+LjVve4b8tdUSsmmqyZg0eoVkgS+7aQmA/9dtX3TWV5pOSqcZJ
wdkeEr4t5dzsXRlw1LMwQz5gZxK0x/zFup3ANWDlOSODaJG0YJAeX3dDxX+4Vz818U9FQbipmz81
i76xBpbNeLaz32eKp/bNK9OTCAIdREXtuqqwyIBFxzEXiBvfk+0h4f9KwgEk9h7XFjjpl8ikFM6L
kggZIa7o0c9zd8TeESxwACaTa3MTvX/P7sQUNOeFY6HCjsWStgjowqtMTRnT4h7vmGerVrNzlpgp
DlatQwShcTXdGJmqaj6qW2eKiszXXstF0EHvnHFn9C0BFe+Pd/EgxIWlkHOKPYCGMIAgZxxZrquf
PITmutWCutbPVrsFdjEP5fbIqaot3DJE0OofJ5jvTd5gt7af51uJlsIFr2bgwaNqKZUKjiSaOhjm
UwF7DLTGtL3pzwYTqB1jfvzle8/QR3Sfbd0P/Ztlae3BUAUweMhCs0JEirQPJrhBTSHId2SHLtjH
Kv+iTeh4dp6ENJZSOFeOkFR3AX1s1Tj9prPXxa8ppwLx4DDU9a9EI0AdCBH0/g2aqiPpN50c7C99
egR2lfmuwy/EMjMdoNuE0q1lpvEuWlg9UL7+tIYcptZRnmMjldycdfqN1wBGDApluJm2/+oLI4oT
YD0vUqvA3M9XJdzEs5+n7De2Skd36gPD/VcrUWuic9Wt7iM6p1bWtoYqBk8VexI5MKTQn/Na0xL5
uvzO+cdznmhTbnMpavbWevWVkBPVfq6WxvLIzqkJJNfUD9J48DuMcIhVLXLFdBz66ifSgVDfd2xn
RXTwe8iOhBDUz/nXF6BFnuywUoVjNF77IbzcjRjvAo5wSoC+tq1OmU0Xzah60zCya5BaFO6PcY+k
Qovq41jHhfr3wETjQ1nDXVyUn04XuqWG5kTbYRu+LL418hppaiLgsfBKUhUfbaZ4kTR4wYuWbei9
VlSxFpKaFye4GXSovO9hqATct99TKvH6I5/tVuMCgUz3oDQvEMlDUI7ebX3YyN9E7pGu1n7Hh3kZ
RpJA/GdlpEhgOSwvROSe2LF0T2EQDDcIxMNsEh8OKbcvCZOtGHgk+96FQjtlgSyLaDy7HdSMhJzM
BaA2iWM6iaXTZBsRZ2Y1P1W/HwSvbvlW43YAiIOAlVuJpRpsqEmgYYEQ4E8OrFX/PbYIroN+7fSJ
8Zr1xL7pCQWR7be9scq1yt27gQmzYUCbH6DvhP8Ch3bDBky+wXQo8zpk5mZxuQxtjZFsJp/Moprl
RDuigAV5C5hfca7CWF82LkJawLKzD/g2meRYrC1aG9XjhCNfrYvM5PL9tr+L7zrLz8YnCmHPvUzf
ql8UWcWhgzCP5NFWp40K0dwqTSepN6mPtQ07bFleZj9xOwAM4TxO1yxVvnUsv9g4+NUKh5QY6gDJ
NDL3mL7v5MKD5shg+Ij+8HoD0kDfrn8Yuz6jzGk8xLqjZ4D4meC7j2S3+kf0KAJbci3FAZHOd9bu
lv+D7YnDiohb/jsLDLdXp949XZUN8spZIBOX7JUgs9WNntYdZDKvTNt7JvXES/f2AYj+epid+iKB
rIb21aDZmp8/5WDM6StBhZe3nvjz6TyMh0bXCtHUsrU62qaEjl/KBZBtFMDU82iBGLZKK1RGefE+
0r5EFlgft7ecAku9pkuJKsKHRMd14303wRhBE647cUHKkAKQsqsDNio/cGzY2peckSi09ku1S8ko
OEEjBkSI4Rvx2zTJiZY7SqMAdqYny7AnnUXT/rGQBQQZUrfxveN+jpKabiX2soXcqC7aEL65si2h
Hon23FpKrPmWo5NrHZg6j5sQTbM9tQG3jcYjkk+GYnhR3YyLrLe2AErRh1Jg2ofynBi8IzfhHO+K
07aDbWMencZPST3hHKzGDJ9v7WEVtZ/D7A1Ze8aogfdVW9pNmQzeXTHCmW6Ht+RUZanI/pFbqNIE
e9ELgZYgzjNFp55IuMTE9X4kQ/mm7m6BYjkUPYK9aP8RBjyyKgvE235ttXnenq9dZHOO/3/nx0Gs
18/SIhpFOuj7OTvKTyYPIKf2hEcX2hlprgYqCFsPEl5GwHtdx1LnO0eYqrVu7hIx+sbkllUIIzwq
f5yP1Kv9p+RGGd8YipGAhX8HeyoDmmCNXiFIvvK9xxZ4iMGap6E/4jAmjqh5wcyTN5eSBCpNvgDw
3l54hTrLoyZCMFs9ohK3pAohewd4ead5lbmv//lzfilzxf6T2hSjc809esw6BTVgm/6YtkJdm3x8
0lpGqUwgyBnMU6H2w5f8Dt61H9S+lgVMG9kFngJvXSx8/Xz+HXX6b5KKxEZBvf2Alg07JW+/awkd
7x/IvZMSRm1yGchB95+21D3IasNyBoFJDWmEjbqxTq/pz6wN9q8k0WgRjs5DFWxLdrvfPKZQf5NP
pFhn3U5vUxfflBHZlsGwC/C95LgLLR0EB//SM9mnfF54ZC85/P31+nupl/QX8pDc585y0+c7igJ7
E5ryVkWn+zIxxDYLOaQDdcj5072OrcQdzTgTWvIbeGLKyYIfXjFLzZOQooz63rngzaspTpp+u5/7
Y/sdUv9uXNxKY1X7+rp8Ae2WWsv1MKaOZrW9l4Cm7AMlLoxdXTMVR6CU8+DXOcxjIuuTZP5ebqJB
Oy/DtYi/fPAU+OE7SQ2+zJh9P9VoTMKfOr2UDG5hDKKclJmQy6Z4ySX94zKMPmLQuf7Ddz/pAm7g
ea72FUHaSH9Jx/alfYtX2Nh0gPpbQ2y9WzVhXNffUaax9WE3bV7E2OvFHYp0gIBiMVBK8DgHSTTv
P101lJgEYXXc9ApRmVDCcjkpFLcgu+C8geZOYppSdn80bz3GCpfmMjvN2h+Zuv8QPvnp2hup5iuk
Jic1NNZ66vDQ6oyeshC958vo8I6yNvhcSo5mnkW3lslxIMe5DKbeA+4THHtUp59pPgt1kjpkPPWb
ze4pfVvTxqCySazsy+QOr18Z7Yq4Jvtxle7dVcYW1E0cvUpT11hNa39V8py0isPklf9ryURTR03D
j1ZtB+GGUFAGc8RoM09hqBZS3cAxNPJrMdbS3SCHoxEdXUvpNEY4/GHO/tPaMIfiCH/ThW+MDKG8
BonukSQvzqEWrFxnvV8JZbPe3L6JZhN+2SvJ51jJQXmftlvEynoDX7RuB0mhG377rMpp1RFnY2fd
RXjVinrX9cs0+LSzm8yNqXpZ1M1oJqk6h9MgZfZxUes35rpc1t//NvvXMcf1nHjjV+BUzw213YQI
99swUtPG0YbiZlkN4YkP4MD1ofX/DqVetct4an8caBu/X+qAsRvOzwSmwolYMHsGpFKeD68UBwBL
WQqUELnOWCrgTtywMKez6VazjHzvDirTOS/4AcNu2te4khthInUZTp7VoED9ZQ25ROhlkHCFTlgy
QKt33CBqegt6hU0qN7VcT/c3lDw58l0ARoevo9G2pQAFcWsDZoFsGrKm8ZYuDV8uR2X1YUFr3i76
9skeyGpgXZFchp+BuVtVydkNtUMLmXckdxvvU63EbQzxLFWiTD5kOU/VKydG0V0H5dV6UBBy9iEj
yRzTIUORf3bjXNMDxURmnRl32QzNi98T2QcBaxvDzUn8tznrjgt22GtJa5ruYw6eIakjdomgXj0Z
FqxgAJQscHRmvcd+mt1bicLh7jRo22mqZkvn/i8gVjTUWVEKI1LipAif5SNJefbPBNmVOSQH2mBe
clEmQuwDC57nrXuoYq8b/YuHzRoF/eSgW9qkNnJ8NjYhKiPSQnn2WnKmVbPWusMtMFBHQGDWSgGA
JVEvLYs4/faHAgq8Jw+E+wa/w2L7n5NjhmzxzY8byxdcHlfO0dKwtRgIldwmK6SBtmo38nqFejUf
wrNl7CbCyuLL/EGEpnj1ISBcAiUX1D8le3M2LLuSUI9Q/jFSfBnqNIrKd5mDhF041WbueCHIi4Ex
K0kwfUUa14w3zK/WCewb2ek1OTcv9w74tPM8sDNpvBlizdblojOVpkujsM4bDuAZaVCaMzPfSoyl
lJpIoQCoRdCYdaSNngEXn5g8Z1wx2yfzrlVWQZfKYYV7AMs3HYKCR8WF6N6yJcAVcuhQIpATgJ2f
GiEJb2WvmfMfm+f/hAMSxy++qlZkB7Bx2kw76aO12sm34pEh4lb1tqlMqotbdYxdyBdLs3CiD5Ve
AQfBANnOg5eroU6Tna9zR5tdDYn+Jv7h1h8/GF3fxs1mF16TH/gs1JCXRiJBSHlUOM8sXguqUybS
k5k2D1xiej3CaYJ1yIWqUGwl2q9q8TTISZo7tKJmkjo7kV1t7ez+6M5FD6lvfLnR634+r8zwDBkT
kqqF8iUrPg0G4tFWUQgmvu8TRBEiHQFmDXD2mpb6lvNreUz1OgOavOnB239v88ADWVutqc0bk4sC
2q3cSKktd4EyZiW8b2PYGUh4WjIS55+bmdMRrCVSBDe1/kPFc5w9atudpIpOWXzglNOs/W5awv8E
FHEN18AL+tVGWUv1vFGkeBhyiZukf0q3qRCuqPbKbF5dq1UwyJujmd9u7VU/FASsMMAU36hKR59c
q4UacnXaRtsBsmE9D25T8JAPzJPyXnGZGl3Iqi8x/+Jc0QR1N0s5zu5RVsiyM5V3th+sbULCUC4W
XoEGDbOiExUE5Gf5avnS0SVw43OcZ4IqGSYVVCi4wgXJxIoufl8Exn9f1rZnj0YfEvsCU4l5r/TM
0X5jSy4iWFAo50wwHqI5yIAkL16QHnEhdDYRj/hLEJqbRnvokT4pVLAox/mNDZpx5CMtUkhPCP74
2/NV5ppC7wo/yRjMFCFnbKOjzW43CgjErwb8elWqpeQk51zbKUh7/+cSF1iF7cHqflzncdMXFseA
IzbTZccvrnvOvz0bBdx1vCAMeX+Z1mUVnINQtknozJKnamnM+ufHc8pbgaLy4HJ+iS9mHuIkojvH
/p4SX0l41QiVlMIOg69Fe6pjsh7t8F3Vgq+Nwd7/S5I0FKAAnaGTsRFCGPGfs4dHMsZEsrq0+xUf
OmgggrWWI6G0todH5qIhivt6a8nHa3gwq+TdaWVSJIxhmQHX/pgUqXFy6NAvH2A68eQRWozgHKa4
uSGUfyc/Ti0aLV5L5Hti0g4iK6DzPuKUHnm03mkaAAGqy5mqkSgi0C2Eb1mFfVnMapolr2s4n03P
XF8SM042mkPPzcvu9wtPuEQ73KSKhuPW+U5i5m1xcSSkPDZImsNBFqJcn7UzRYNMWDaiSYZmlAXB
FLli2QYjReZc7Kf0/dTAVsKcDUArM86mkQkIfiN1wKR3+Qyt7AzNi9J2oPHej0QQ3rUADOxBEAY8
J/lo7Q66L34E7tNUsHBR5YlgANJlBgT5pK43o1XnqU+pmHGYHO1Z6S5l7nP7Kh6FWUfmIMIKXjRD
fIlDF79LfTAkpNmwX/I0D/7wPzJapEYT0Y06Dhl+qtAmkPjKDB5suhgc8upNEqANcA1Kad3K4mfs
Fam562gRpLsJegvI8qvNuGCPA1NnnAIBczSmG8RO0u/KJu8rAfsvJ1HQkxV6Qs9w5ZL7QCvB6fIU
/p4Mw4z/uPlUcGIr+8IdHFsPOfHHwsObAvWKvaE/zAU+xExGSXpzQQli+JTWV/UuC9RmKPukQavZ
SMhdjpqw6qkD/jfG9kF+TGLIldVn6d5X/36c3OW4OO4Y0FUFthNUPARAvfWA0wxUB7WJjsDL4E/r
36OPs8t76j9lw0+627EKSD8R5FbmIPOun/bGUoxtXxUUfrjvMfsTiprvbUJZeTtDk935FsI9tLzR
bvfSE45u25TVldE8agEiXpzFbVL8f3nJxAuobHTD81YTq/3i6dIz1Jdpv0Z2LmR6MdA2PjJNRMP/
2/mZlSKYxY+RhhL17uvTPntP7tdbGePHDapatOl2aWT0Nv87wo6j3Or9WAGhj/Kge8awL0iBBI9A
iIxCv14XvSnhUx/mUJoSdLVdrduCuNzR6aZrI3q77j/tac5t1ohfFAyDYV4rt5HNEUhWBhMuPnbf
HPkYKDNaiFfE141LA0xLxYgFIfGYCm8opsEfP3WP1SKBnbUxz4/viNqA25w1NyB7u5IVPHEii9Mm
Ex/4KfHIAdwzF/xuP0OTHfhK4HjLPJGDGzMBRIJ44dLMz1hlOeZVFm/kCJsIQZG0REjaD+/LFtFv
FwAJU9JcXrY7bo0eXF5hTXgR0J2PGvAK5SIj0x/jToqmoUlOoNANT2iapCmXD814yo96sWmrHzyI
0Gyen/XXbespGWPB3Pj6U5BAA0V8yNzopobpK2ndNcM5LG3b9QL1TmUEY2W78mkHLF9K6Kzz5J69
7s9iZSMdhrNfLn/UD4G/v5CYQ3BVJDG0+IQkPrr4TuUK0VV1m9nYXOD/bph8cvvel/nNNmVzQsqx
OKWEJ9a4WgSJNeRFFcTkmJFQg6SiDOSrlG7kI29NeC2SJLe8KFYNod43GWPitBiZG2irZfmV9N7c
AEphvUS2Xr8zCaOuCNZM9E0/ujtmQkOBvPQf4ebvBnELAUMj9Ur2hW+zlLRlfu93VQUSki06Ohyl
Y+VlZAJtjaaCmqGEuGzM9UswTtdMtMRB7vnHNItcgwIr1xJbJ5k+LxhCSOSwrm7LhMJaVEWkgLty
XPskrpGTFlQkwwBg3vuq03OBLO+eJl7TP3b4gy4aZteCscNeU2eqak92V/LYFQTVdlcM7RUh5sZ2
k2b6HnL8PxHMAYQsmeuJAC+tp9eDDaiN45XeWGTUlrY6P5hDj5741Yx4XSq2AfunCnSJhFT/oYML
BixrFohhujJP3EEAnuwAlqEOAUPWUGPG9O3K4QiQR72q6kyDdqQ5tuiO2SdG8rmMUGFSqEbhOAOs
qSaxod8ba/ZGLHw1TqtMV/mbK48bqZ2HSODPGSlqfmURF2OuM7FIxQTpOJa365iQyIIrBuecCq0B
80woREFziv1HIwEvr+gI5IISHsnL7D5MsvXMjV8abmuzKSoXDK2RGuaxPNIuNRXvdsO0pBdOkGgZ
QlFX/OvbnlWyWi8/51Ye3TyeEYjWbYYdf6euqAazOuTMj9hasdBiKuYhshzca2xvOyRntyHVkc9M
Y0k3Qkr26d8rI3k3MbaddNZkLBw89G1vQl1q7oPjHvbIg69a6Hi+qmUsAZAuirzge2Hep/Ggzj+4
yS/1op1cyVO1811CLm6Qxj2ZIhV5c1a7nHbV8DLUbiwr8XsE9TGmLrf9YRSoK/4nCKbx7zxPZHBE
jWPhVH9zKqWKM8U+XpwdGIPqhSyFRnTqbUnUslI/2aRdsOB6IRNJWUNNQqus3ntw0wKITkDeBU0W
xiKLsrZQ7xAbz15AAKTXrrpbzkNoJ/5hKMGK8D9Hbt3lZP5nLwfF3GFVay89/lUE2yNHDSVEo7o5
m9J5cKfHFeeUwUrQLOvEUpX4W+yQQO6sSb54CArhCYg+0qeP4bGCBKpCaLf/k27hf/kDMMTZADF9
9XVwAINNVIsgN6zXNww8XNx18SkddaXiR8YrErw054PGaR4PJPYW92e4/trZqDCOIx57NkCQJg/e
dbiWAai9qGs0znKBDvEchTCVQZDeUNQRqm/M6rHBAwR6auIiLiQHzdWLleTukFUkUgi8yOMKPyqp
+GNPTj3Ji8juXP17LKKfjqe2md4oE/2aCDRQxfigufjntAlcr7cSfxP8zxzIc9YwF1bSx973gCfv
SEQ3UaBjo/nRlF2a2Uc/ekwGyQ/puE+09vl/ycVg5H2wwYDXTiD2zjmlIx4ptJMtAHQXxhnSuRqL
fsUB/s8dJotSUtfdSknP0c52sRC+FHn01ZnnjS/T0FXvcbvllswE8jG0llpWYW/wOcgo9G/k9ldP
SXBcWU4NAJj4v+KsRNq6XyU17Bs+9ER4BdfX61SNV0CozBe03kzAitEJaWTcXhPtzbkfwqo6KfKr
ZLAcXAeEThHQbR/534ZnGP+cmQTnR4t9xEFNrEEKkCrs4bb0t6DGyUSNBBIjfgon6g2MTIrhQkfU
jJ9k+ihcfePtmXpsdHyX/Jrq7Tikv/XUfCASZ3VoPR/GNLxedIMHw7G09ylYrR09UjkOsa3P5FFm
CP0k9q1KdVwBYIXbI1iGIAo5ZPNYzT/R+54qeadV9nBqlOjS72WaLMsDUNfpQM7ZHOZ7A5EozbI5
1+Wn086nYmfp41g5QwqfjMkD8HJJb0KktFcTRJnz1HKkNdb73MI2RFLc5YOA6cZJUZhEd6Ahu5sD
TjuQdAhvPAPb7kFR/8SYXHdPnMSZHqW3yx4w8kgoJcqPqlY9SuLRq9LvmMjI145ojhfO/3NFnMsc
x3eL2SDT0OsDXPXYdY7nbzJVhV4zV3gosbZexZyhunTh9vZMZXBXYDkrp9KyCoDAgP2K64AfSaaH
LwebGaDjCkAZ3DjHawczBJOionHVrFM2rL9eamdjLdUYYfLy7kBgBx3hmfaNFyGbTMoXmAGtaBbV
5e0f6iZeqP1GAXwjpxp+wxCwwnDnYJBEswL4DGV4hH4iHXvl+wFnf4tm4MFnX1slmPpsRTglX9i7
H/8po8v8bqD3oUJuoO1oUfeTvu6AdJaDMzfvBL1CT2cS2kDoEiirdOpPvU1oB0Y7g5EiCnlwanJ4
xMmIhYSMM9jNlunJ7gpWe43dxCTkfaqC/VhIvZwA2IAlha179AlrT1Qbhh/XMdiT9sNa3/UiTto3
ybKBrqCMaocfXlDd5/I7ZqJfgCPH0Jew03skeTKwmPJbwA+bHsrbjprdKa4ulo2617AmwgIGGcbM
hLT8kFpaaYXL9EHk9EHOvcKBUHmI8PNC1yYAeMOwR2Ewpzxbi8d6Z496L2z8S6zl6K8NMYw8txXo
a19RQCSzHP0vZWTZbIp+gc2CL6KvcL2ANLkTEIeuWjm1UM/+pCVBvxZLD+JpT8w7nu/A3ZVfdfeV
5gNZfhgCZH5uRxfsu/4+v6j+NN25MsX1XQ8c92J8+OOLkFvZG6KOMmRhwqmc20mI3SkMHrwpV9b9
jY3jEzOET8dxcqlp0zgLrSye9b3lhf49/DZdaCXmspTht1UBrwS4Jm2AyGoA2nU3vjLneQN2d2cj
q+wNWyhkzzswPbLBwE+wZS1WWL9vToVQM9L1WlDN1GgZC+ne4P58XZRdsWSvthKcqOiNPvZnkiXe
TL5rFB9Iv6uKOi9tRAaZOZL50HP+FVcrPXObDtxZDfVVYVB+oJ4uKT4w6yntNLAsP5f/PW1EjIf7
E+N92CTsHao+fHYTjR6+ZQFFCz0icMZ3mOMkZ7U1kxXScLwc3mnItu6Y6B6jxN/nNafJxLOTR7Jq
P+mmEuyUDk2mKlrJaxhLsKOMJn6zFuLCOw4HoKTuUjkG0FG2beLgxQUDDKBU/ZIwWhgKoeBJmyQz
9nKD+4/9GUkUXtpJHGCHjK94pKA30pKBWEYkA/TXkh75oJfgmqeCnqiwX6O1Bq9hHkLMD/TGPZW7
hfR24Gdd4aMRbiuboYURpKQAjrPUBFDXRD0JSz+PTa5nko6DKqVQVBNwjNENdtx8jfcIVQVcuU3J
MQNQXNkmMOLzqymRnkN6CgvtIMF3DZihXMTerrmfpg5XUROE46eiNdVhKVFlZ+wgsrB6H/mM1SIi
1NTY9G3WlwWoC3DAE31WUqRKOp9MrM+0DxHK9bdHiuq1sl0N6XeURsArRjwOKafhKngk00dEzQYi
dac3FkHmhqVICmUxOEvT07pp667Ea+NtAvkfmnvg1j08YM5+49cpHRCKDeIGjbON/L7jzHkWgoY4
qWRkANm4hXlVKSh7OvalRTImzZddq/iZ9qcyIEU72JC3P0aEsAzE5UrGQ379YnXVQwvR19iVam86
udEjIoAa+kAkDF8DyjXTMVjpxkA2Mi+kFt1QZkLuDngA9Yz80VUePubsbE9FY9+TPM7Qf21G/kOm
fg61imnMBgfYFJb/ILKwEH7qSkRfDdo9TIAyQnNheeI29UjJEsqpPFxUqnrJIU+V6XjyJp/m7MPl
8LlEoY40bvRZn49maBQ/Ft7LEKkgwQDE/43AVeFHDYy27siEMmyPNAusXAa6nCdynmlxkf2WeWu/
Ima/fiYF4v9WFLtuXFBy/KXkavnI+nW0gC0XE9Cp2eUlJZXe7AmjtRmZqoOXgdb+ulzD0dJDdcER
u1u5reiZYgXnUzjMuWv2Lv3mgyzY5bAjSq8CEZYN5xmlawDONsHSVk/qgwr8Byp4qe33NKmm4+1N
X+EpGb9Pqr2IXTN52S0g2VKuPJpi+882s7tJ0tSfVafEpLCaJ84oLolKPW6xABsDBxDwW5LDlQgQ
hH1mKA+CEW4U7ePBpEpT428Kwtc5cQCaI/Dxmo62D3G83BoG1mnrIoXx2tSX8hLB1RO8zBIW5WZV
3lsp46rgpgCeB4j5pGtDNAS1h9HohCHZkt0jVwLIUrpUQ2HPOlwaH3ir+COBLdYSrdeiyIFOK9ge
7NLIB3E0AwFKfKHvJyPOrgWymU9tq2WneFXJ5ZxXk9ooPYlC0VP5LEPeBu79NgbGrGPVCDL+A9if
jsq29uQCEKlE2w9ohxlHMQdgxUgW27r9vqPtUI0ur7EkWQq8itai7B108SjTpfomyOX9BuI6cn74
ybhgSGUXRewDSKEGxHi2NLgOTjI/idHRLQXJoSJHgX14l8eRUM6J0m4CrjlxxpJfb4LEWkZHtJMD
abLB1wGFwATlUsWXEmdb0KQqadp135kgOTcsK/5L+P/g9M3KhDNkfKxtL9lHwqKl7kzWLx1E/nIZ
5q8DOAml5a8hifCtfI/P+oyPVm4GoYV0N0ZATBXsdx+XdTaDo9wW9W0jfQ+acFHshxDblcQNHfAH
Y4vSFu5xQKv7hKgULw3/CHuxGVMgqteZwjRlG2/w1TxmhgpvBqeV5Ns+KpCGyN4zVQ/gSezD+gvP
KeX0Y7bWoWerEOeqZQ89h82NzUYniUzW4+/uB7v2jT5qSP4J85ApEu8Fu+5R9AaVHwJTsJ1dsfJo
EaSpBxxs8MD/19HMxLy+V0mVvr+qrID+Q1Fx9ao6y36dS48v93sSJN+Ut87PKaPdD5x/IvZ654kS
rzoIUAe4JRd0UOvQh8YJZzOEHARVPK6HntZUfIyuVHVlCwndPfRHmVVQtSlnCj+mGfWgteRFZg9M
3vV2Cqm7XRBqUuIQSw+J1F+tQnklUr3dA9u776PsjucdtRxP2ME6GJybVeH83E03F/ZotH2rfFP1
9J76abs/IEgTez+eKHBgEqpiUG1IteUgSyRz14wVGakTSvK8nETIvyEv7vkh7Siy5WhVlGDjL/Gb
Fsl/ToHlYuzUzRLtyR/1McnhTl6odWNahv0+oPDamXjIQVAi+9ayMmy5q85QkwDWL1szUIh+VSrB
jWZFdjwZARS81gEnlHBHa4pJfaXhcMhFYeS331zsoQQtR3FOlYLMU+PQxxolP6F3zPqebNXRNOsi
TbxXwnwwOa0Oa/w0JWbHk7xpef3lvByNkBjKFf0jFrXnCHule8uz49HHSEnxPwBvAn19gwgaeMlX
ZbIHiJ47+T4F74DCxB0ZlgDjYS6ULEnqmQGsxGQC+fuAbGcPBYsIBaB7Qvxr7HjLO9iElEZXRTpJ
CFjV1vfZLyoJKp/9MHN2vBLCUBH2I99aOLz0oAGm9qyiTBCmJUFuz9wA7U8NGr9L1ACMnmVSAbyj
RV8oxGx33/mwv61JhbyWYkl4a4hxkSJUExy5jOkCeOZRT0CcTc4SX/SJQvk3L1wY2eiKCmzxOsSb
iDByqCFKtxMX+VFIHwSD9nrYOof8JOsGmkB42Mc7C0F527D8BwBYGahupY2J5c+8v+xoLUCowQi6
ZoSEquOYjiJmSgUoZ37rUOF76mqUbFkiXHPqKoeDJMFGShE5e1oOjrVx9HgcboQXNFjgLBMmmDxY
bItgUc3bLtcjTTcKY9S1vFEU4F3Ytojy8qf1JkbSh9M3qaE0sn5Zu3WETSb/QRiej/k0V2/7jTZn
xUmSpLvi3+peqtPfP8wi4F54cDurWrL2MdZvwdA7RRv3+BIVVZOgMrsdAqH5r+aroltgozblfuST
kQmaFxtS8i3fYd6A18IPYfvsASwTf4elfANsqWu4OHR5ZGLllKVj8/xCEll4KLuWniyQ6aqS7ePN
iVnWkyQjQvJjEZnLeGp6ms7zLtr82y+J2E3J1YsJk5iWBopHsHXORu7Ma8fWVcXRzHTPpY3Zkr4o
BRRajTmGCYzn6ZcAtWSmd5psSwkKVXo3jf5OBxpok+Yr8ZQ7o3GcAsH0o3QSlFrJ2wBil/H1VKSP
QTt1w6+bHwll2ESA33VVe/eJ73Odu+LPpZF6eYLyvbiBh1cFeuefTDGMXcEyEMFDlsOjiGOizcQ4
6vRhzrUwcLEfaD636SbPmue1pfGpaen7VHju4uUS/YHqjnO/6xnJvZE7MJnzj6xw4TZc+k46pKuR
pKri+P0E/UPD1SrCmjbOLQUZ3IfGccEC22qR1z9Nlq8AWVVg5qtL3jDrmPSkCG+/O+YQHN0I6vlS
yEAb6gCnFUTF4IcX53H3PW6YiovAHZkz+wxLl5joeHomwTPZ68U5aTogwNJ8DP2QrMRmqo65vl7z
MKZxE3me4z/szYYcgvTy4DU6Sq7RetPL9F992KVY4dSLQbWgfvKK6aebTJB04anOXVDMbaGnbi2x
7t4WA0/AbJcNBCcmhI6/jpBUC/FAVJQHIGVbnEswDkZNjsNHib89fUpoPJ5jNSvZf1T9C1+aLBwS
ymAB/vxgIonhsrS7xIDb8vklf1UpOwBrnTLtCIvSGU5xADiJuuWfgxemP9ij2egvk8Fpkda5V3pu
7O/0EsrFWwZsdWlZMR1VM+RESjPHSXYz9IDOIG8qdvHMM+XY0Fl739OVDNwHYc92k+/IfAZViFSn
XVXn/iADunxGQnbn0dlzt0q9EBWgEOBshechlO9K6kSePep2LimSYsBAP3DsZwI5LQpKS7FlrBBS
Q2G57sJWFeECZZSFA7kUOBC22NUaQd65b810JJgdraLh27RDgFoG/TGoAw5v9XU92eeBxT421BLP
VQni6a4FWLfu1naHhrnsRxfC5tPhID/WhK4J0FQQsGX8o4gQMwJ8jr0EL9VSS+NPJx3X9kL6NnGt
skHuR7NLazBvBwKZJ4v2bfPdBipgE9f4LvOTL83U/IkIT1giF6nlfUph/jB62/WMx5vLWdcG1eX7
kgRb8wTJPrIfx+fOQHH9bbyRHqbgEdh2jTRdBsW1Am0ymRuK0HS3CfnvPskpEeKDmtALh6za6Gug
QZ9PxQAMd1EpHKVSQU94qiLeJCesFvYXc+2nBv9oT7uYzqAXln1i2SrOIu/lr4oZIOoGOs+eVOgC
0UciiOKIe79RAG3acjxXkF8kpPILU1giYsBSzZNCQ3Bv0zQUv4qumGkFSmx43QvEOkJFwMr39U4G
1hdCLDo8VJVUzTkb2VGxYfTN60wJW9GOgLKZEAiZRodxYhjhx05DM4itdGJ+5uelZh8egBDIvlTX
I5+CjfXL5bVBXsHuOljde7/6LzANmz0CVNOKc7OSf/X+SVyTegUInZnk8BEK33VJkXegFJed+wb3
Ndo3mMK0iPaHjzQa+AJ2rATwVGXgNsL1NTcoCyYqtzhv5EEbJXprR1LUkDltBzt97uOJMprUTiyn
Xt/TImnXlDANKZDkDxiV6WkxcMso9/aer00DmNfbb3ok7nnQrHleppcqzyq3o+jVlYqtNdGIHbFY
8m0DD+ctxCCTmzE/oTTfwsLdIVjt9QHYDt8lOdZiP/fXgXHhEfJiGmABlg1hzRMeeYgmHTF9sGH9
tYay6W2AN44eAOGvVIzs9Ifjv+Ruezz5lcFrKvNQ96wlZZUh7uZ9geWxBIR4STcfHdn/wbKu6q0Q
xiA1vqLsrUV5ZqsCJcoyHQ+7/0/OnsSB8LHWL1qnQYjUjBrMeRzRtjgP1qu9qStSYkB/DedKaZAi
etq9vhqP/hwJrEPEsZqrgT8oyJSsz+B1JhwWgRwixhIUMRyPvGNtPjuF0FQqfeMkBJkCjZ/esKKQ
t0/qBmMovzp3aJpuvG9l+4ytcAno6DKDp46GGRIufirUGQOKDXOON5iClNBIw+m7bQsre3HC2NH4
oC8bZwsIiFRyrHiLKXdF7iIohOs8bKDfKC8jcxqGoGf1mdaaUyCgGgQ1d50+eTazHN7jogsQJy2Z
/lxqcRw9tLeVaXTq/5VzZOU5Q4VbkG1tuiDTf3a1Axm4gS4vZlF3SOMVwEyhuqQC75D5ssS4LUSw
j2Qpi3QAxDsGT88gq1rQnRynku4Zo2Pxyf9SaQcxdjOMqeVQGji/o/POMhrxsKel2lVuRK3elYkJ
k6oVgs24Ys9dAjGedG1dBvGC/+yI01K1FUE/Hytmg9byEaP8aY/wVB7M+lt2zhOOfHX8cjny1SmC
SIX4TA0J6Qj/5OBEHSipx0DnLtCOvONPgulWCgy1fm5iPRAhINul/1lYP0uaPX5ABuR6x30BKvpy
Y+nsrtWDFWcASnjVvz9MIO1nRejEBjanEwbGT6qVqaY5fOtIBIGNTDYnnSSJRJxQABzseQGyZh7U
STYM7RtybzFZJHJNwcxpbvS6e27ZG1PtpvHmzaJ6Abm0XnqOVUZusZylU5EuF7nfajOAvEWQjsu0
5pFPElORcvN7ylIiL4bIdoMlbuQMzUMNaJmw7aq0ffRaS0gNJtKMirGPAZDZIAyXI1zy77JWEVOj
Wj1jKhJosGYkfNmR940PgLoHxmqXIOFYJq8DXuzPyq8New4GynylkypiK5OjPK14WzItmJL+MSsK
nhuEo/JyLSS/eYD5oV9C3QFkNslmmlD4NUhDm8hNwyS1iOt38eoM466Uuml5qEw1DNcPBsKLhFWt
yaq7dOmjx5noqH+oDnpOmiJeBDYXx7LvlWK7a7aT4gUt/HGyJk23gUXg8KJbqMnW7MDqTP6xQcpk
Ygl+9lyc/7Gah0Nu7EGXn7xOrnne5SvcintBc5Q/AKyApel/fh+4R+tP+8e1Rmq3dxbmmwspjJhP
OrMbJSQT29+it7t8/zUc3L1nqdo2S5uKigRx72Sch3SBDqjfF2GmohkuUOEVy8LJMUkWaVJKbXch
upcQ2ei+OkxrGZi1G+YWnKv3iC3Bizi7c1ExdCY/Ak5qqcMytXnwjGH53Ed969wEFF6B2Gown7z/
2FrmWMkXQ9ZvV3LpYQFDVP8x1yGDytLTtpk5tRk6O0Qa6D60zE+dzGSSp53cEK/CtTsciurz4ZeJ
kV+Sn/PqZK0xAO9DeOSC5JZU7yqMf2dlQNEDWue7/NmgZEQUbUgRhXpN5+kuAWIZnUaT6XitPwQA
9FXHF7BsSRpsXVvphoAwJzbYLYzwR0We3ndEySui6OPiuny385tR08FbdjjIYN9M50eWRfshYj7B
DDDTn7P67MNFA/Q0x49Mg9643yD4mt4bTj7Wj3Ypt+TfV0mGXhwE0qL99ZZ7h25YQlHZ3XqwFyQY
4giGFsj3gAv4SvJaoMmqNPQjolQcrBEiSjSBtRFLC1xmes3cPuBQir55iSn0x3Qo3MJ+Mk06pmRa
Ss7rIh1SsqD1JRPGfAL7tnE4gg3v/IlEzkZeZmxJm3URON8P9dYI0U+iOnAKPSwkWj3Dg7IcZ4uW
1acYLSFDtoJu7AzoVDX77CvUXE3m4Ox2lHVk5NZbzQx6MXVvuaAhsFn3tavvEiGutDrcAlNBUEpm
2f8lOd9yltYQDysjlLcSzU5u7vZDyUdLAzIYIgXdVsBfizqAO+DnebhzmsOPYojghf51s9DNfM3v
jTDbEZoA7CnYw7+kfJWUBmzHs9dDGua3YDI6yHjPrCVcGzew25AGFTewlhvX/3XwUCOIWVBD85xd
TYt37MBCJeW0NRLlbZtqGn7/SuKfSVdZYn6K5Wj/sYR5AIgUhIF+/uBq4LHTsSvfkuEJgMoedxis
lcLfmLPOt8Ie8G5+YDduMzbd5lXaEzSf78e0oXEVBCU1kZ+ZYUKdmQxSguQLCj1ELQQwO7Vj/GXA
HrzfKIUt8sUONLzuxtBmyI3FbtX8AeSkI63Nmjmw5l8I0/l7Ox7oxMR5bWfulzJRrnC37gOcst0C
Hsu5/G4UrcmCQmOSs8nVV6SHNRn/iLh5TNFkChgZKEqKmB1vuH/WmYkGpWHpVkWQrJBddKKg0Mpl
zc4mus6r1CSUiBOBZ4rumiy1OxFJQyFAoUaWl81fBC5AtBYfWjal5Cv7z7mCWhSxnwzVSSJayCl3
cOvTJbZWTUX6w6X9CJB3vOzUMAu/PJ583HuUEMeAAYFHzU0Tr5WF6Npgv3ohbx9jl+pi5vWLwkTc
Z27AORx5GeVny0eOdHtjH4uGCH/TOuxvRlKKTzsVmYgdfZ64WrtZafmRJYHb6MXdWhbHBipuauGr
KzBUfwBis71sCTggYPzDkBioiglxeVVrpjMvz7kj+aGzQOsxFwQY0deySYLtq1z9kiSTPEgP5HVc
Cg6vlMG1XI2kvV9z/ThedhCKZOk4tdL5gS+mXjLH+4bNa04mNh5ex2DZteeze57KmA/kaQ7hZXZ9
K5JPBRXbzPAz1S61/PlMO0tOHaRkaZ/lsFcfmRmr/2Df+NzonJpU3UxQ0dB7okHMXTxhA9xyoqW9
wRnPuSk3Y+dx41xlBGd8tUtlcpGNpcgiANy8BlP7Ay8d4mzvPWlyZHxLKP9MUG7miYF+F6eAz7LZ
FIzse8nUoh7/bxJ0+gpQAyoI3+JsPnA5DNu7oik39aoq1dD8gIijojTZTI+lGFFI/2oRDNd5HVSi
5mWmB7dfgvPGaEscEhpQY4Vy286B45074u1pZ2m9JUGU6kHbTMhVUmcnT/gl54wRm/iD3ol2qGEq
vYOLf7TImHu/IZku8bmk9xh1ZMIR17zTckjSJQVPd64g7JZJ/oEkCdR1A+iSHUSdhV5d8KpLMLdZ
0alp4Boq7qAOSGwvP133Kd5Ef3Klg/7VT923rCTENyKlw4KAKWlbthFHexXEN6FYW2EdWJX1HE+Z
OvypJoOQXZfW4WxOTbn4zqWFcJluwkbvrWYOkdWIPqt0fXiQlQNigTSJxwmEAqCa8qEy5SsfzD62
aeUZRDrmmw64up3R95tAlVro+2CXMmFLMbHS5eREAYQ6HOc3j3TM1DzfqpLfCc8Hz7faSFl3LV21
nWUzJqfefnaetZbt87wHG6zR45rcgTHxev8xO0AskOEeG4sS+XUyaK99h5jncr8H+r4lIboi7E07
XMw0eHa1pp9HU1icyJFjXjntq4x6zxAoRKxPwRcJJ2q+HOMr0qa4j2Xas4ALV5VbFp5NKeT/PjLG
sTf1ZN+Tk5t6cRnUA4oj2vIVX95GxKVU/Xx1AhHd3T0ao9oKJG8BubdOX/VkbQNy7WOigqixwmGN
m09MLBhkBwLH5x+q0UJh+4DLWkKHAaxAU/67CuKkoyL2pqGj3qvBVT6eYMKICuDuY6HTo3Ane7ke
/HEmnWY+fb/LGo34AGM1L2sVx+YOTLVh5nWbNPMaf/04JT6XFu7iJRpBbPnan4Hlv5E5ccSi9sxJ
wmFLxUXc5zSmj9iy/gv16R5DoBbMC2QDCd0WxoMc3H0nWX5gUDj8l2s4i7eiD5/lknJXBErWHAzK
LZUrCv1hLQmhYRYXmpYZF3LL53YLqZpQ8afKxNVZdYY5BzH8LBr55qJZTmWTYXMwRDtYCUFbXyO3
JZdefNOqIUtEfwAdvITKRDARa2F7dNqdV9qq7PY/Re6F6HoTtbN9ab4M91YXzR+Nft8SfZmBcqMQ
BEkWnVWzQxWrPnddQgIq4qhdVCNVOOHnFC+0bHOA//9NuwxVsOJ8l9htgzaRQvW/mQay8+dTCXfr
UPh2+6P5gUQkeMtkpNpb4vBGfG3ScmTU/OuY6T1022S1bmIcaktFELIrfkG6qVeX8m+iwQkHeE9t
3RfEaY/jIVvFpRe/49allajGelzQsk0uxYN2RQ5DYn/xFMvMxO1wgxcJ/NibRB+LFCDMm65HLmza
oAH4tJ5U4gFcbSxI68EqfBPvQc8/ZVqlKNTRIDpId+8lbtGnbI7/fPuSv4lrfkuAxeW27Glj75bZ
niUwquPNqQaB9vkbmrPouGgKOEV03fcx9dZZR3ZjG9Ax66sSFB5HlDEHywHRuk3NGXb7WHaxOBqI
ZXNLP0SY/JDKO35L8uLr12CLHE887tEmmfvP78xkT1Xy4ooSZGl5H1DQFs1Gn98zlI9Pi1sLDR+u
BsrsSq5gyVAYUk39HzxaFqRt4aYL7/zGOzlCTGTpb7bezFgOjWPC2EaZe8hZvmZfGj8fz5O4giTl
vp0/LfUOIysV2L9YHx36v7l2ZZgSOpri9sBduLHvuRR4xP1zpLzoo9MdJLlU7aSrBOAtho7fX7/m
dNMp1NX+5ApU/NfqKjYGNlNzQfxtvA63iZR1AQp3dI4OxyysbePzkWMkDM+jvZYOuvjXN3wK3h0o
NSDXyDiZqU5XzJ7jF3br/LqF83Khdg/tYL0ObhLHg/xDCgFiGgcRKDIrZ6Gf+1rXrmY2fTXhlDm8
ZWUJe/t4/xVTYzGDAteKBF9xGuOP4OrF1pPjeuL7k/4r7EtENZ0vRj1G6Xzq9cWcbrFSJaIX2uyk
ZS20j6BheusxeFMfDLi4n2Uw/Op1G3N3swbiZPWm0C96sTlbAT5gv3HLfYSl3rhnu4kNMY1wm8ji
+YxQ2rbUpx5NhVfZ/lUxgoHOgV4dPsSbHqMskFkVKNDRpGFraCflwrXG8eSdVzVLnHmYKEN6cZrk
yY0GgqQUFFHHNT9pSdS148/I9iu2wcUn7V8q6PiwDyL1qYht5mIHVoXmBWl4amVS+7CUDHpGdlAE
q3JrO/cM0SM3QRQk+zBxVWDjtkiuf7qeyt6UWl0Tsq2dVzQs8DH1U5horwTWcxlvr7cMZrHAhjnU
sNF1vsESqR/lgq2u2vY9QOpr1vmmYmt8TzC5xs+Q+KvoD5IEXU/5a3F2mBq0X4BBjnUbIP5GZsAX
DyQHpaAudCCkb6HI4PRlOIdZvafD2wqPIu8hbnBD14cGrlrN5VO1iRZ26lfPG9OfXg3NvU4R9tHj
t1+hCUjZlOfAmaRoTm0s+ilwl9/A/AQT6c0+9gv51f3Kg6dSd8md+fyElBXxKjsBF2LtAm3+c0OT
bLZF/YVtOy+RCiX93DC3eIMtY2TSCmW2oGgq4TGrjOVIHDH+5AlRbBsokDMgW4akqKjVfOQNMmyA
ViO11cDnzHeDKP0qPpH2RuBsGCHSZtouekAcalkBG3sImPx3OQftx429HXg5ij34FjcUqwvYhjoP
w5Vj2l8KDUFGQdNBmD1THp0pVJak4vjGH7E0e9NmeuKmTQHMO4GSTx93UXSsBDyZsxcvD2ahvo2e
TAIWFML+ZpUE6SI4XIlV8BJqcmxHp1c/A9rxPK0aeayFD7frhC7YTU7zgk088MXF9hhV3+Q5+1uT
fJy/ZFJkQGgXj/Dr/Vs33Ei66910vdBND3G2z0g7tp6Nfu40MCWlTbA5PQi11E3EHem/4+XzubkB
2nr2IQJ+JpRevphGTWzCQTor6szTxagdZJBh4umYEelacjw4d9Vmu7V3htOGn1Xjfo5wK+e+NaQX
pn78eZsvWd7yn7mX8iqRRSD4yNft/Lg3Xifle2KpXO9vWKXvTGBX2KqZEWjYK6jo4yZfYaHLGEl9
rZ1y0Bwou2O4do2ghDfVRANCEX7tiyu4memYG/5A8q/AB4f1im2iei/DklDaTB93pQpI15OZEYTt
vnnyD+oSGEapaOsuKKbDIHO61uuy/ocwpqQjPP8NWngqLuo8UjVsdLuEDtSWl3AwI2SNxVnpDWNw
o3OHxVnZFR66LpGscswi9WZTEdjQT7KVAgJPEqGPDW8spVH2RzjiuRaHpycKb+Jqcuixwn+fi7XJ
8QD7inrGrqCU9BfYOiRsf4xO2DPHXMDTdnTguOm+FD3qEpvsSsd3DiieXF+l15mSrmdY//92jkcM
bHHrlAvU4gcc2Dv0edOAaZFZ9HpBA209EWY9LRfzmQ6tL5t/2XElqdRka9FOCD1mjG2yFPVounui
X/5SjYOZOH0OBPxPB7gzwj2SAYqGvy4qIVPeWC0cF1XZsTWskwthaNW6mJa6m+ctn9D3z5jtz6To
DxY13GLTO0oQM6MfG5O+W0sMzg5u0F84kyS4EEkF8wCXeCRANS0hzPkmywJeJ2/kD0XQbW1LUY++
dtGhB4gxk4dzSuZSmURbLQL13qbaaPRXD48YYXUrgNSs0XkoFgn7KpuOgRU+S+JH/XgGelZ71s2H
UHhLD3pNvFg6eYyxiMV5//SumyooK6H/aFR2oJjcAC2z+APf9g8NNTG+JZA0HWRlzcVYnn5eibwK
X1zOsQvZr7j310e3/sRYp24WBN2+pjzFm+k3VLzG1BFXfyNJYmxOSfWyVE4uRaIf54mguUx/op8Y
jd7uC0Tr584cCRrTWcZceqEfhAm/SKj8fR/KwL7FklSPGXYPDjQBBbPez+p/gRTcNo5uOTn1cQ1h
p2/Hd19kv4uLrJb2KZ8WmsEJ+c77Od4M5cJGamy2k53lBbnM7Pdj+IHxWtnJYOndL1DI6gh6CbR6
/fHeLOGo4by0RaNJ6B7Xk/8uT1zAKBmgWsBw7yysq1hktOcsEr/gZdT6arL7XwApncGC/XK7BHZz
jK/Uv/DKWF5B6F1lbXyh3lholJ5nkTGti6FZ9lvKVj9HX8NjiP+Ayziy794tcPN+VD4YQZiqS7CY
jAtxO7agCrS3cAnWwGNcipQhfoBQnBea/LRxjZPPKtAc9xXvszLqKXpwnvlrMxhdlzHl9i2wvLNM
XbJ5LZfqYdY3lkUUtm3jqaQQLRQpIxg02Bri5vCc+m8j3ifIxbwqhoX7OYNptNmRaOtzekiUXxeX
lv3W64WqgEgsGFQ+zGrZSjkJrs5Vi9Ga9OeE15JKyXsoJQqwBhRtq8O8e0bSITRh3+bGenlNEoen
bOLC4AFUNCsLmI9MZSYTj/d1akn25R94V0k9AtfDq6BjYM+YIYmpAhUqp+iSbwbG0Vvxf8O5018c
MKT6lbhJn0HKinQ7bUsmx0zoyq3ppPS9Smo5+gowaCCdpiH+1MFnqH6R7XOljAtDfzsfpWgW8pfb
0C65NjZbBkOk8XUtAiFBCP6YA0lxFAOURGkeJjXcviJqSVQ96oxsZpcadar1zoMwYBT+Xj8QbJ9q
6eVVYJarNIlY+7SMeTBq+D06H8rATQpc6IAXOJGpGoZIVZcDBb9r97xM1/E9g+1b4XkUoUhIHL9h
pAYj9x0iGAIJRJx2qJ6jD4wxm34QfCeVVnH8Xh1ANFZHvvp01mpdiq00RVn+2qtY4okQZGykuEi4
wwqpWjSGFtPjre2bQ+xbydACrgDCYKjeVAAU2nqrd0lapgADgo1GEPqH/Ra1MkE3tZt7KSYlLd1u
ze/N153pnix+rTUAdmIA9Fxl2SAvF/ijdx5hrz7lwaPPFax79T2ML/hngF870p1wNSnzhj5MBIib
qAcQceZnbAma/LK2q80lMTr/pTcm234aBi56efZjbj8qtWXNikMM9DVbAuAwYmU/FDmpmDV3VUNr
jDhD34EXAwLrfQVmYsoKqirrKKV+mTjsrJfXuwb0G3v8HikCmbaLlDkR8aiEfV0AiO1oaAIJboVG
mcmvI/rqvxacgEQt9WmfVbegpiZ3ODbjT0GPwOOUbdr0Oi4D45zHwTzYsQ1fccfMea10khDd5guc
3L7vN4VEWFxNU0EyFq4WqfD/ehQCzZNRppwsfs9xE6gXUHWDZjgK8fNqt9t8cLDQ54qPJjUddB5T
NjyWHtkGRgo8DpL61DsFK+uqrzApkWJKZENhnl3Ym+MsN3Rdxky3FGNfv49Svzq8W+hhgs+NQQD1
hFCmZ4+VadjiGnJg2Wj4UuPWp5OTAzEGoT2oakomvNBRnWmocIFE6oY3sPFVD/bXYQ2kkoljuVhl
EhK6zaeQTF92ljCZJS1Hsj700l9zYWOXfx/3WTM4BkquojMpAh63CMipM4GVV9MnCXxoF7Bwj76u
jbvTttNaIvvFScILAcX0uYO+NKqjEYua39OJA5VK5UfcZFOEu7p/ITB6KkzqnKcyPO6Fj1qSShTL
WOPfF2Vs1ZgX4a6+YRysOFx/InucGC9fe3IPfIxCMcXeuZivZuhq8Yqj6mGM0oYI2a9sVxX3rS2v
u4JobYtuvBCmk9O5NIzo3ME4nVwQkCwiOURyLMOBJVYOPYUtro+IMSmBDYLbnpgADaRdGxhFl+Gv
mXfXa3bPJFmcS8GfUHg1H5m9YKsFvEEjU//ZjJZAULX9ocPN8nQ4i6A8K7TEjtsyR3g03jdcjFDf
qXYTbpZrSeyzcAVAz8Pe+0hFSxb3+zkgOY9Ov0uWtgfkJQU79fqWiISkMk0rQMdQC0u3tDjUIBiN
1Rl2JmLzUrFiaLPvbmDgFmA6IxseXMLUUgovWmXZNaW2Q1WX0xJG7UrKdbsgto/Zb/EFcykgbqEF
YIZCLHmkru2mxAXAHo2NJcQ33aOTpf0GfVnXwkACrNKbhek6uj7S64wEEUia6enlmCwk6caX+zVZ
THvIfA5fM/TFuGRxH80VQ5W/nhMlSa5w8RZmbPoHran5xK1Lnl3SIdYO0Vze2Hwf2HDjnB2AM/uD
jmw/nFcTR2oBmVrEoAZ85DzcuQuykbb528RPFyctW0hAOnMwCoNBj/0GVMAjgOSLkMxaZvlFSaf3
1rCKmxS8vAtQtoI/oB61fs8cVR/QISGOb03Cno3Ue+gfIa4lByuIZUayal9JvvbVb5ExMBYI4g1l
kAVOPmYnvfV+J9HV3unHWO7HQmoII5Jdx+BA6N3rwjSG8L2J12S0TBU0GNk6L+o3bpZlStaIlqFI
mdQBczO6hZBZFAzzR8PSCb+dyLh1shpQk/oPwYQHehWQSIu4miRTm6hI6FThZgeaQ5prKo+ZyFIP
oTZ7D0oK2xo/53mgTmtNudtM1ojP3uvQLrf7+WYTaKiFjWW0Z79f9rEKXQLCPpQCNvBUuy4drgAs
UWLJR4AwxRZ3PnNTnHYP2HTRmVFfLIzTU6lIzmPJbSsigjzovBZliwUO3xyJK9GFIvn1J9sDDzY3
xSXp0S1W4NUTC6BOiZH+L5lQJhCF70t5jI9C7NAs58MsJpGwYjzGRUUQJ+zNLbswzBTyWnXxhPnG
vw2xV0ne5tMKWrinkKgQzScQMFIDqsYNSHYksWmXp185eTbP8euBECHcarKYCi20cgs77DVdo7YN
a+XpX9rN5onRUhNQpvitRm84MqUzB+SdAQNFVJ8C4AyEv/B/JqKpr0gk3mSOsVvwTo0YtAK66hqF
PhJDb9TSn/RzpTNe8oEWEM5gpDXjeTb3QlF0/lD4cdZx1huwktF/MQgbiIuYekYYoU62Ic9IbBix
RHKyrCEVDEeWlz9mxxf82ZgiwcvS1D7yPvbr3kmowkHFDQX/aPzEv19F8wTwEngoDs1wyWfdKVXV
IB4jQCVPRYVWLW5ZBAco2P/NQeddlwaNs/3rL199XdledGic7gjuhitj/JBlyEJVb+MYb0I6+P6A
E85Wyu5JzyUhMeDL6Ozgygmlw+WOo4Q9V2ObIHfVe5BvD4AU6ZyuTfw5OFvy40OHmrexvglf6f2i
yQs8KPvcRrXyO/QirluT771dNPgBckeq1bFXnkFjKQkMKhid26m3jpsa6d2pYJpskKn2TZZq3eRI
BaK0OkO8lpFvJQDJhuD/gnaQ+g4ZzvnmTS9QqylcDRX/oag/sfW9dGCLsN01jzUBfdw7pQsOqFkA
a7NUzX9JxAq1q/8N5DYGWbEo3rvfCPAtOql4ZFtv1nVDXPcaKwzrtuWWDBQdC+MI8SiriivXo4jz
yQr2y4eS0jGXv0z0E4avZYafywr1M6C/WNlnZpN8RnLA7nMJu7Zz2P5tYHjeX2L+CWSbqnWih2mz
8OiMd34txn4tZX51xnCCx6T1gyzf8XWcrUjJy5fDAJWarDm1scs5wtaTXguxoO5g2QWbP3jrWjNS
4BNk8TfLtnDTV1DrtUS4ZU4TsZYi4Qk8wfvQfJZZOW9oc9uMqFeNZSGKacab1Rpey0uTa4wObHfy
iepLyj8QkI6GjBdzWuPiWkNvk9ARddRAScXYMv8ibr4U2T38c5aPDErUwwZVIbIY7yhLOXpfeQyh
DUWqV0296qbfzgfVS1/gf/iYI7oTxsC6TMaOrQyDbtYTqPIG7gYlAE1NDgn4WfeJxp6wCKY775IB
F7ToOsw2VM5WotKh/2o/jzgzsi2KgEZdK2PXS8+0g2qZZvycepFfDfISVcZQjnAg/ymIChsz5XmY
MPlxuTTrsLKkhukxdB9Sfcq/A5ZJdumhSX+hDLlDpYSEt+P6v1oUqVzAXtGrzydKjHFxNTvH8sH/
vLTEUTe1T/ZeM+Hq4Nvtsdt2MIpcn8fg119cTIfOEeVIEHLR8Imfa9W2APwq2L4ZnpPAlU3San8L
e0ePwM+d7sqp1J5D7k2YleAmoZbyf8T7qEs3N+9QyanOnkAELxPoy3Xwu786QhSMroH7I5neZDb2
PpekfdL3clicLGHdTr9YG1ebgeyC+ibLYJCBEkbE8le/J+PPQ/j7pjRN8QTEGan3wTNgTClKurKN
D8f7S0pO5r303K7N3nX7ztIV2Tq59CN1DZYl6OG/Uo/f8kJUyM+9P1svSzIf9suiyFPvP6/0H00i
89YavCp1DuvkrDFg1NqCe14/DQzY+QEgK4a4ROf6cGT4tv1ZCcJUFvkL03NLT5I1foa4M99ni8yF
QErUmNx1haGUuKTqDI4ashS53Gor8/3Ehdlub8pg2inh1WJr8rmJfCL8Y5+HRDAN5DKqrx9ejBV4
rqkoi7g8M3DDkGERvlQmkaxirkn/jPbq7peywSpN0+nNsD7vrI4lSg9hguG5AvUaZY4k1yFg4cMs
jQr6b2qsEsLSL3RKP7lWYJOzKkxGqTJpCdyEZShHCPFdEbDeh6NUbeMwhu+mec1cTw87sNn9YeD+
BZsnI7FxZ/iW6FZ0CudvXlzvR2gA6q4j/5TOeaNDeLtbt/Ae584wjyLo9pcaAW1joWlMEYtVWm1e
BSD1Iaak2VHKxj1SLs5HHhu1yc6C5LMnQy9HBfUo4kjB1vD3UX9xxa+QJ8KDVcX0QoTM+u8BPdMj
Ca/1axFlQzwBRDexRWkcgXYC8JUBM73YytAfIEGHlPfvU+2IKnprwJwk1vQDXklBri21CGLk+DSb
pD24C99lSe1QF/FY3sEglex4p/+qzAHejEWLw1IHUKRaaSGOdbhzj0hOdcRQwI56O2RhI4Xb/CRN
DD+emdhiSme8UywoYZ5CTkFhSsrdkNsisjj8tIR1SynIFTGIu0mauFndH+Eids8r/bDIbrcLlAbO
ovTlqgDyIKYjMMdT/t56wgAKwsbsGwcJO5YO//Qj4fFM26zF77/5LvEDvkrpyWIXgAOCLRBw8zsU
CTZ0uHJsSrb1LyQGj531GlrvSYYb+uqrdvssn5mKeGPdeGmYkOUiPjukdCtFFnUoywE6Z1PfxKdY
JWOzw/guVghatZrwhwpvPwtwcBJ+V/PQburVAyeVluBvoDworrQqP5QnSNstXdb3N6+ZdAS9Va1V
IBsk8uUvkIUSlwbuKW/s/sJEgPA10gu/JuZS39uetRkq5fwL3GGgSdiDbZaNjuAHLQGo75UEYCkl
8p5qrMVV7FWwzk3e1BY0j3isH9+zkx1tqwLRgMFaDs5Gve2SrDmtoAfVhKuzbfN4A7nWdvdgZN4v
hjYMzdKBe53EZHQg89mKHWAuzxYhadvToWPfZI0+kVeFSYYIBMuNb+AD4S+I9G8qm8ufngwMfAXq
55Fsb0x20kssNqx3W2M5SVUXQXOq+9McgQ5jp2R2axDrC8xuQFrI9bg19sQezpootaoPfbQWNPiQ
gzc55168pG/hazLkBPGxhQTbsFeGzNUJBegPBhU5H/fGHnkp/uGledckkaTsF3+Lmfx54wGe+soe
X/DhPIx6LC6It/RH393IwCGrIcGjB6mDMvt3pyME5Z/yIsvyjKpPn0m3ewh4UAKedbjA99fScupS
O+TeMGrPyye1N1JMbbqb9pWuzdM8rsbQVIn6dGCPylHjiUdTxqpxKkXTz+f6aA2p2/UiR7TJL0PV
cM9J2Lq+OOBkt+YDO9/yIr/j+ISRN1L8/dnybYZeKrlK/o3TKL1jdX+bISOM9wI2Cbmw1aiwu+g7
6opf+lIxKRhfTZpyt9tD590dxvUL+Pl7ggDb1wuo8h7f6PmHuWAbF7pcLpLZLaBnhNgXDMOdTQcI
EWeiwE5JFmPcEZacbCDDXwjpCfvy10n/F6SjmAnaCfMA3uLHwdUzvrAw6FO8IRvqTXmYJgyfgD+1
ypjCojl8jC7ZpwgvO//f9t7ohA4xc1EWXM+e66tp2DifVjqT7Y/D9w2KTla16BpXCAewvnWocFEE
8kXQjllNUVIMVihtcFWHMu1Vj1NG45sQcKdPZe7kiY97+TX6GiLPtkNuk+96vZKuRKr26B47aTsR
656EU38fn9rxAn7PIgd5kOa0gNzVsJ4F3Ti5oteVHRXP8DPIcKlhCt3MWeKU549dDCE1yGqbvBvf
UriearXBIZyD4t48IwNm6VjGFTPCq3fIRAq9g0mXCfEGHnuBryEmUaYv4lB0vRaTf4+XO2wW5+Uv
LN+4SfN1zO7EfUCB/bkH0H6eGZBQbOnCLAss1k5URkdp6VnVRQ9UsvP7jkzTW0dxzz2eUtmWSxK6
NGOhEb6gI4r6tCFRb/v5QCxrpGJwj6Poyk85bjpgTu0J+chJGl02RjbIo87DURtHS4suEwffA8He
WK4EvAzG8aRMkAt4/Hlb8H0tYXDFz59YUsbQgrWQ4iTOaLk3tElP50YC1D2TPBbsgSxrMjVh/ojj
qAmvX5rWxlUbNIDTMq8pMJA7UpGs465/xCUTi4thbwXMQrUEkDhkqw0SgD4kiNVVy2U7XJm87nkc
O2WXc5JnmA6S6paxQVAJ3Y6cUGAXwW+CztrYb57yuKL6Ua6yCmO/r8DbekKnFw/7SPA5Ld5KC3Pf
XU9YvaSNAmqAnqpBfgrQsmvNy2Cw+uIcvQpySnHDltgerdAPnBuOnGehoYhU+aXV09G6XjTk9qbU
0cw6Bh6TpIyErfCrxZQ9j3K4Ldyt36JL630uv2aQK+dGCu7geXTpOTy44+FT8jYpob+owFZ8pISR
OhqIiVDvaeUbDYWqCXwNbG6a+AgZDK4LyglIShg2PdJLj6ZTESmw4rJ1XIST7cUeLzDH+IKyo0c9
2o/mfDGVsJiKvazF7auH7+mfTuvkhQO8L60JeYwMamrQS9YRozxy+k/xUfzHtoM+uE12nzKUfbWN
sG9Yr84RGvbxVPqrZnkb5x3PNzgmo+lWRSsAZw0HU1dLt+0QFF+BxfGd4IVYyDkUrwdCAgvr7lcR
f5O6XknFm2moG1OW241NkZ0aMvXGxSQXjiRgXPsxKBkWuD2fyLaVsbdOcGNpbQCO2ApNsbyRrl+Q
Zf3gV6pXG2bw5pIES7xbwoJay+yGUs0zHZW0X4udMZCh+V/PjAF+S/s+e5lsOUppphOyU8bVn26b
rXMowBVKt6ek4gi/fcshtWUz5WXp3PxoITHyaoLeCaX2yb9XMcnrHwlDFijFqqnCdJeneP5ISwcy
xPtb4PUNhrc41cFwHXuzo1jc4cMm0L3CpEQ009bmx1SkbZycQ6CycgkLBKvmweZNjaHAz0aWK9Dg
++qSz4yopSt+Nwv5vAMvliHk0wnyJB2fY4B12FeXOVNNn9/K72CcA/WHcOzQDOe4w3WTkAyVmxa2
HCu2pt2BtIDLyZw8+oQ07sg5jyPWLR2DuKlo7HDfGhZuOYm6LNxWERJ5N4hZzz8FcBC8kHUn0uTk
jCkC4PEqld+yOuy6fuLjAwbpCJoJcQR+qugqA25ryMXdoBrWeoFmFidooAX+aiDGY+ENZi2Kp1SJ
GkoTkRzpdVfWApjDVIVE5OvcxC9tRy3+ZqJASZGKFCJoOamj2nf1WtuegYqLvuwOt2XK2gnNufGC
K9xZnbE+zLJxBBGcMRk0KRJwnsFBrntANJ2ZnZW51YXZmL4JkinSwA9ej7jdOHmu1OjXaTHI0BjV
+aC8LtEeVpHyEcSaNAQ3VS7pWWa3w7uhEgVSFrIcURfmEN1FRiexUyv3RrRUJjZ/YB3K9AP3Sd3t
0IyRJJ8wQPgPFybdW/NtBwUf9jtCTdC/Q4CfIdwU4CLo0UT6PuQbc6a9pC8ZoLAtOVR7lxNcrr4U
Z5VUr1hBYJi14vbyi5IROWr36Im8/04cNPnk7o0YuPIC9Z7IEpjXh00GpmCwIokbe7eCkgCLWbkM
wPNyHYW+S5B/Re0cli73evRP6KGEuCKIyidDwDH1DZ/l66J3Yu8DDWuj+OV+WkUgtGEpffkcUl3i
uLF0YoPJTJ038l8YgBhAoQN0Gs6y/u/6DtqZkXBGUfUaMR71KC5JycyZ6jXlYW73iPqZI/fLWdu6
UlQ8dPTywdzVqdqhQHzo6/B09S64Y5JpWk8JoZnouR4R55NKKnYy4bWhzPBAJ/v5rJxkmef5d5aW
NzoM1EZZtw09mnWHMZd9DeNjWOsik/q1llJlGnUmYmYgEe85X9U68WLzBgdw2jH1Wrq+q5arUFiz
/aJlVwKJ9t4hsKcGEOh/DaA5OEcSb03G0gBTANvnxbkgWsuYuFeJV95v37HZs63jsMIP48kchHKQ
0lZgRM63tP6O7XB2tOyXqj0DWZtDbMul2gRpAZe6EsuYpxS2/bGuf2vyE3ZHlnw06tF91G9LGd2A
crSTkjTcX70EoVoiRgNe6X8wtMwZ6jZwTN6u+BmS0CgWxYiY88MEdfqZ/4QemgL5JIk9W9qDNq2L
AXnFEyjQRAjChZe8dlTZ8T8LxndpPTm+27WyZoHI42fgCBzy2m+V3ZWNQX7xsJu2qyU/Yn/IYdsW
bqe5+mHzfkIAkD3isH/6P0PH4VXW+33jcyNWSg455EX/227EuvfNh6JJXV8MUC8nmqeBquQlg8CE
nMPyuhD/x6w9SD/l9kjhWS7aHn1Eo72DfbUzVZbepJYDumFesR/VC/+7rk3MuI53IVs7TOL2YELj
Ax6dpn7QDPE82IeJ/RMp9WcP+X84EnvDKEbZOqqrLGrDQjh7uo4+t03BPP6BgPgcKNeZj7qxR1OB
iblpx+zEn/x0HPPIhQnCTevC3E11uzKNy7JWisrt97VsOxJ3/uiu8iRIWo8TSzeNyan35y5Yi5WS
Pn2JC5a4nFHVI0+v22SUWRE2+8fULurrgTYHDiGzEvoqj9U/D00kzjRYP/KJVcSB+A03jVX93nbI
Dt6XdPlaOi5UnPne0HF17ZmiFnri4k6FgpkHXIfUWgJmCHPqKl5qNokrSwSH9W/lOxdfL5+zl2nQ
SuZl5xyQQ7eoHH7ym7i7qKfoV2OzPRqqs/6I0cCULNfp77NnaXV4V1k+ZF5UFy8seKY2uEgOt7XW
zRK3Dk1kI1la3h3sdAiliXYGIRm5/Tj0JGMd7YVFjjyxTb/jdev7qLSoNbbmBKaigwgVRtwbBeey
k8wmDHoCguca0PpxZvWPCJPb61PrgRoW5IHZHyNK9QxZa7qOA6i38d+1moe6UPEiUu8TBPlHaClj
1UqvGWFBsAcidFhG3JtAhmRcW/sRmdfr5KDa808GB2FrD9n+JHZ2ZEj+qWUHmLWDOnyVfuqgfL1p
YJo5oZ0EK8osh4MHVr710YAU3Vqbt+a7vlx5TQzf4BM+IJGgKiXni5VeysEYdmvPlTQ7Pjw8D9S5
66wL3dsbyN0iR5Il7WV46jkfYRkSknd/VPfWBQWcYnrPHHockTh2N0nIma5es/xQjSbU4elURzGg
bSOjN0It9vxOz3GIpVXM8PzFS+3mZxs59IAmjnQcfTeJd+peq7sO6xV5Ohr6Y7eVRMNqXhRCH+h+
ut4/5SRCeZK9YmuuBMhV83568CvGfRTQdG2H2Yw7uRnfNjAqgJO9rOvCv9WtZ+u6oq8V1PqzpIHW
BD1DZLd3HTyR+cEXXtkdmsSmOsLjGLvs/lylL/jaryC2xq7mBTLNjKGkeSaOvi1+1UjEjI4LtE+K
UwrN7koYHjlILMmyWF9lFI+LqbT/dYWWgxqQLgpXr6BAPZjk1eByEvlHXmNTiUyWI06PO4eEmmbW
bS+Jz2aWYrjggdqvJpml1DI1ErqyznrfP+1WnhrJJvYsDyuxypMFtE8aX5eGCo24SKhdRt4ALNeh
Qxl4HP1i11AMpkH/a+1NLdzz8Fe2Ti4xLkEO85PwNZZKISiqm9hU0ce5/3lGGUt1ktRQuJA9ihun
hXbofBQDF0511mptSBbhJkgFyHYEgKzVV2P0SY6u2nV6eB1hX6AaFUoldkWWVu9kikKzvCYQNjC/
RI0nDTc3JaHkeFtz3Zbbt8EVZnjQikSIocqLil8RtbNSI1DnOyzc5LHicY9ZotVvntaLlHo2XnnX
qDkJFHTtMPxfACqHiOYwF2cvQYJP0SnEO+aRoY+GxF5ZpoWbEEppWFVdi3PAfAMadO5pgRYr68Ax
gBP+nCEJkoZFJe/Whj9C1V9E0og3aRA3M3B7QFQ5xpTDNo343tat6MXrYGQ2LTtLeHUvseHIN6tE
zLM9jbSbLc/QDi21j6Usvoj/IjwY+DI2SzRnOkrPQ55MCsvbaPYrwxGp2ZPk63Pzvx/V0CxYvnNs
Shey8YMtL3szwRPFtC6lQXrZUDtRj8+3oexfepGM2CZXzyvtKC0Vrvas/6yT6/ykk3bxFZd2owDA
R3NNkbAo0Gu6vuq6i93d8aL7/V8t4amEFHtPvr2WN5AYV+2tl2M3CoUqe/tIoTpa61CdafcTlrlx
y5M8fHdUc9Wja/LCX8wcx5rcIH7csSnUJYQd4q5yOpNY+uXNhiUwgHYbUiBKTer2aOg7/z4diLDT
maxc0NfOxHCt9WQhOVHPV4cJ/hptAZmFabf0Hmnf2UNNDxJvIxO0Qy5+IxKlq7qpnmt8lzzGZiou
0zfLF7T0ageD/6lymSW7JlRxc0/5Hcmptb1mCcbBhdo/56J/oEHtuWQPZbD+hE+TJKU2D1SnNG4w
oVZSOyoJrw8jA0sl7oI6H5DzoWXFbXYav8U0GKx6mK8lGp/jS3SLaxTttDGN845vLv8ah0Fb/wPq
8c/azQ4eyU10C6JEdrzTd5KxMHi+1pwKbEBN8l6QNvlL1MY17xGzv+bmYZY+i6phyKfBOBtQ1NzA
/lBwlxTWWvRt8RLgQChucgjhPfTAKWQKhsgbs/fqzPeHvAep19+x7bJpH1twt8YSoQTBPogSqFMI
bDnIpJhcvNOU9yniQ0wAg8h/Tal36dWKYJ3WRpVjC5NQAQbZQKwn3DXnVreYsIVEc9w1JFFUQ8E7
+zkR1kgunhS6Jd6uxuTDnxfsD9AIWHVS/NyDdylQuCFZM8UQISw9uX6GvxZfbJnFe3dKsKcWhGAk
fBhM6aAny2OSYsNJXHqtNmb6oGBnkb6kw+eP8+v3shLN1NKqB0xi68rjaRiaCb5sy8frCwaeIJDE
wvWgNpN2KXpRwiGlYtNbzkHpQI1SnGEVrn0tKjAL6Y1ULSt196VkRI0KW28+xz2G+5CescYyWQ+/
1LI1ak+hwD5R7/OkeLXBi/j7YHGHIZag9RfXl7vQQeh7Yhoe9DmjylKhPwvWyn6mhGYufDoh/0No
BMfzKVUnNhlyHicQ7+4ui+vhA5wx5hj1VWjqGtroZwglIIqmcE5R6dWLPCpcogrh+FSHOO6vEybh
189wFRiAFvL93bRguPmiPDdDfvCyyQDis48+Ll9uzhCfQJzs04qvE632rqLKcpxGOrAp0NpjYwaM
pgbE+pNg2E0HxhWZ+CUvoLSirVRhoZi4lRsxMl/wV1haXu9NfHpK3/ty8FvVPglGb7Hxq6aMO/wT
7v0a+2hq359mgTZ3gwPfvEU8tIswLC+75i2HsxjLlluBKt+OqtAGPCN4MNPGa3wm2KPh0dzhQg8U
GXiBVYSmXm7sMV7MBV5O3rqTUc+80xNHs4gpa3fwy/xUPI+rO5C1GnFTi2htH00E+ViWO3QleYkg
wAJFLpbxKY10ot9N4KcfOdLjKu3IwBnpUIBjtTu9R8a5CmMA2JpBTG2u8xktBNT8scD/vCeIUmwF
Ta1MjssIY078ujYOR5eeMKSIhnDVGvWviQB4b6YnwXtzMGz55w6R5/HeOASKEfUl+oDYmCTzbQgq
tTQuchpeB045H7XnhASrSpTR2oogqDhqu+GViCx+h52KM/T03+Yo4CvM/oySc9mMsRDmlXxHvXhC
KCZsOeLXOCRIGlxVzWtFUdruPfg+4GUElnbtTqlqzBeBlmtemDwN4mWU0KiWU9bP3LIcfvYd/mAf
3wyyTs/tDP4nF3I2uZZGqsi7clbivIdRHtiTu2IaR+poqa9tSDS/SLbJ6JtYns7zgqUW1ZJ0trK5
7pWF8gbnHHLwdJRLrms/1npQegfz0EwNT3JF/HsdtqRAewJY5YXsf+jZbJHJmF+xSBwZp4Bf7AlL
H/k8AIbLy4IzNC/O2oCQEwtiybPJhGZ9udkJ9MQsUf2P3MFPf3nPn+/eA58jFwQfam67UUZwJ8V1
nkEEkeqdGUp9Y1iXVHBPF9gU6EKijkyNTqcbBNMaajiPyEqZV2ElWCTL7Icc7t8y86+GGgZDVvPR
5PRYDrPhz6VyvxAhMX0fZqVT3Rl4+mg44bw9Rp+yEYlcuSdwdo33+eKPyQ4VznP0lV36ghf/bSpS
sZeTxQQLuxee+jRnrnlOuly5r4aoebWRsvBeut/FdUjfiIJXcr/MrocRoontn0JmwiTynFKV/4oj
H5b+E7pgWDI8WX0IWDVWShSNRPs3Pf33offFv7W+qvEIXPN91oIsN+Id1aHXoWuwLJn+U9fOVS2k
V/cpXPD0wNyPi/35IHwRpR4vpDc2neGxH657waLmvX6XI8uX4OykRX4TeL10aZVWIHq7VlpsVnB3
rnBjK2E2n4IWMmsWB3BTSZzDzcmIsrm+d29BQXV/R6LwkJlCG6m39Ni/G9d7HGyd53CSuBg7h4wI
D3PHNjof4o1yyNzWFMXj8O84xQSmWlX2xEoo03pCnwj+1NGGl0Jvva5ZV0nvJgiXUaOdN9Eyuoak
SVZbN8Y4CSnIUjkiGpC843mgsPyrLtcGKq1tjdiedqKaEO9eKIhBR8VmxtP1L6QRlBk/pdSGH12b
Pv3kd1ohaSARwnLS0JBpWvc+hkLB4wJENYJZBdRxIrsajbNd27kZwKqyalax+6fAc05YUJjSku1l
+XjsoZf0apLYnqQnujx2ATFIxKJzL7CTApQPMa+B9O1VSeYJnChbRYRP0s/VbkGmRGWrnypnpYX3
uQ2cBd73c1Vn/5PE1D3zt8gj0fRR/57MtkDtjHOJ5UdGztV6y8xouVLVCPQBkgBqHyijwwsxhQjc
u9yNjPjPO6TE6EPFW2sz9xTzCw7xq4bntLfa3QBWUIqM25DFvztuSrCkasMfjQkaf+z8l2mnvOcK
kkCZBRwSomlP0lsU2USsng53FSyxARUnWm6nKGVdQXPvTZVv0SMdiJenrNSkkYeoziH+57K0LLR2
BrtMOlSow6By0MTrOQMIASv6e86PWMwqEyOLMFIeoky/2WFb0/H4QegmsJA2qcujvEiviSfzCrCz
RAhmsAbKWdqIX0kquJHpXfGSlK/rUZDEvIdyrKWBWvNhAks2TALy6TtCNKMVEt/5O4qlYuOCiexc
80CtgBEmUKftTKZkD1INQit6h+CmDEikvKCp4EXc8/niosh02IxM0X90zeXu1Gw/x0b7kKT0lCGz
D0Kwr5u8/UwicCWoSm5T0vFQZZgOzFqFGL+DoWgua4UBzXajDNBGbaXK2kFhudwcVRK2OG++i6j5
XD33gK+fIn9km8yfU3e6Qp2T6hNQhzVNnCRAnFPj8KKHBWJaZe5u5ohZUkNCigikFAcALP4y0OTc
X+6fTCJnmsFrqmsjX1oRWBrjUuH2JwAvkxAvkVLFxVeHpZQ5EiElBeGI4KePtUYVU4pKtrASK/dn
ukZ5f9rWlvCmCeRJXyJAAO6OrJPtVV3IeX2yRay+Vjrd+vsvZdD0uG+ie2WEJb+Uz5y+Zc2GQybt
RIHFTFRllw0LGFxfNLXS6gcjFQMv36zwZ8ZebOUo/bnalDOJE4aJALkWN0rU0EXj4rT1sl9ZYjEv
ZBhhWmkGRRcOgY2yhWREWBUM4/pTfSL3rj9hWi4ewQrFafldky19Jfg5rsh2y4vDvVwSUz3L7vMa
ErmfYgsefmc+zrn1dwZCmUEYBcB6cLCwkIcMv02hEcRhyeQEb6BHlt4xtt0NQjrWXCRzB/Fp1kJd
MQMUL6lPTbjbJM8ko8vi9ck1Au1EdJV8rk2Nuaemu9rW8IV1nZsXOl9pYumNSeU60s6TLhnWJS3K
t0yroTAa5GEQZvIrIkNIqVf7jGNK7pmHfk9XRysWM8oydHCcWQ50VsYWtWUAocjfUevPnVn/h6iY
J8y/BxvMqX+hdBubP4mQKcKnAfOAFoDYtbSvPJhljTTekPAaWrNkGxJYvsUE0Hn/Dj90CBqNLoQY
b9a6EAF7LC6dgBA+pPDDKb9iTblVgvl/p0BTajMRuM/YWXb3FwfT+ZZPhQPzS5haqqU9K8pkiQlw
uWWdcSF9TU6CSRzUN/IwM6M9Vm2rXNT3liMVLKo739Bdit7iPQMtDA7Jx2pjaQjasNU9nDbSGA3e
7792gdNVmLQUGlAH4X2tUOdvo03BYsms9O0+NHqDMqpzY05TmOwYQ/QEJxz0kaRilSLoJ7K6A0g2
wrTDMYS7e94ll+41UPf/uFOLL8g0x37qwJRhdJUtwsmiv+TLIO5DkYeldTgc94+gchGiJPWuuEPw
U9T5YWhkDnkelB2H9NwF5kZn7dfwsX7KfujEvykd7Gnv3zkgfA5ogBQcbug58RqBleXNw1UcU9t8
C+3MJuQQ1S3ERXtkQsAAljvlCSgdaHYOBYOsVBhVRoassuHYSOsN9d270V3Put6C7Ek1VWEI3RC3
wL7GjdFrtIJyNKNqdW8/OC1dmC7e782N0S5bkAyfrD+0FvZkFH5+puM2b8z5Z8ICiDjcOjxOiroU
UFL1Drc7JrNIOQffMi9JGOaUm5ehTrKoE0gRuhxpee3UwHrm8zEIZ3e6trBC4Kehu08+fyG829Ql
3vKfQxtlmQLicMpeaiCUtzetxbFrKu9SA1eF6lew3++XmIxBLxxr8JEUW5AcQYqVx+NWntXev6Gx
J7IcnFP/68qdhmY9qQUMjymno5Y9kHL2UkjC47KkUFMz9OoS+0Fa0NdfEeVS6hk/qjgG3eOYmZnl
c3DwaQPwuLpNc/MRcb1Iinywlf177FQXakf/21I7bHksr6qkW8z06yEf+uPs3kCfS1Brle2tMtjH
XdjEy7f4Qz/6o/JATXz654cFfFHgxDZjNuGGcr8SAme4jiywZCKFqAks1ZgVA6VAFYWnG+6yBGW4
q6qpNJw7iUAsL5JjpTdBlqsoqPY1mCSXRuSYK0ArdOlsXhkvKEsHXcb3AJHAPQCKpuFr8UOqHuro
EYjYFjMFpwOx/45KZqENiuF1UD2yhZLUkuQSwNg0NXcRbaOFXsCsCceLUE4tzT9r27UryvM+mfdv
d6voaGufSmH2CPSnG4otspgEEpLltSQHuEpvxQSBXUP4LkC2ZJViofKuuMcA1kL2DL9ntEVkqcvg
Jf6NnHgBxMRnrarDlpv2Ojhe6JoNgGCc75+Tfxs8TTTldKrcHXu1FvpABo2L7p/17dKyGRjj2LRg
tIapKuKuvrMa9xBGF4Dwb5PzCRibdETP0mrCqLolhiar2lvpKoa93KAdfgYAWqOno5wd0UabUkfj
9eW2b6/wqOfDW7eABX78MkKk5HmW71izZDSNycXyK5EWkI/DhVjZ3Nvas2hPT/CyrDhcBYhOcWjX
4UlgbiiG/fNc9nS8e2LqHsobLrj3/bwyqcxQ6vAJcxUVRhM9Zq/qiushBRWwMggM1XSHeG9hJK7T
Ux969m22o5H2Xg38XuHgOr5T2mDuNlJUChbX8lJ0sKiIaksqZZI8RO5WgztYE+9dDx0pibpJ82cz
1XiS8GQA/2cvXM2h4eYLMCrDbqQkW9EEcDaIwDefH1Sfi3fqEGGmcG5U3IeuZhkfSiyj/R3awVPz
D/5UZDaYNsdO2fVE8VFWd0Nxh2zUvTD9vspuVrFWcSUGs0B53A7ToUVZQ9UgGHoVFbVeJP6RtRKD
LcNDhiPIhmNo0GoJ0OLDHJIfAaGwGdTcJmWd2Md0JdAkzi5v85qfFSDPyOHWv0I8QTF2J1I1PPKk
RhpzYU7CNE/lZToQ5/YKIQv8uI1dmo10VoUiz90HwmWYf7nGvxPk5C4Vc0Djtcmb0Xud3HQoCyi4
HHMXwJInhqrkkn5vSojhhV4mttnImUYbdMN/nye/uuCQk5Ax/QsUxCgH6RN8PAA1GWkiajGM2qc/
64uAia1GSkm+2hu0RwQ2w0M01ZrwSIyCRrERmCI44F+8JMQkv3Lv1oHYZbRbrVLaYGS4Uqa+yrir
CDZHgyhsqlmRbGszwXhYXAH6iS+hiZwMGH7Q4gwERnvLDrI75um/rncL9z3VTPJ+yrHWFG37E6QV
p6+5+uTvxiUneHswrT4ZBPI2qvh6UmpBq3RJxvIvTvkJiHxBIXaMvmgyUWIyP2uqnyD6JtCIWdGu
Xs2gcqKksmq8qkE+DPVOKgU7PSMc6ON1N80GM+hPfwhcLQk3pra5FnE/1a//hqiD59l7ppPJEnG8
J4b8Lq0bMs6scEPG+ZGGYd+Ebd751NjWpcA+T4kuFJqMiGASkhZHAUt+DTOm8wdQdP7mES5doNO3
kzVOB+rghtYzn+FHjYSXr3/WxMYCceI3i8b+a7lCzo1Ea0t9RAMSLM8xEAcdih+pe/qXqImKTr1+
D+h+fxFrrkO+iZqn5N4QX/RUWPxDDohox6/VNwFDQfyi6KCks/k8vM8opxVRncFpgRm7FmYFJiaV
/U9h3DoREozAj1UNyM+gJ4ERyq+s9p/+BcxPfzOoYC5+5x/CNLmURRJs7tieVPGMu+7PPmt01yCE
RuM/PYstJNC3BUxiZIdeiFXYgYvo0nSuqdMLbXog24Tljeg0+7DcTUb8rl5Ui9rueoYrAd/FWPrV
9HqGCNrhMjAag0415F6oCd0hgc/XmfN1n04taCvd9Tl78pKQQFTwh+98oVwVUdiZDWzU0F1Bv+OY
31B/upsC0mzfW0pshG62pP4NbBK1k75YdW7yQ06SrEZvYGlQDwyjnXZO/1cbxQWXOnbNoxjtznAq
P4rAXPemFMRjO53qNBtGMYtgSFtQkPfwrrXt1pqeYHEXRoxIRevcdxDsBF3/9v3zrIHTa/q4UFIi
ZK+fekHZPL3ga2MDAB4KwORx+fNJSyJ/rGI9BUJPi9+ccPx4DNweROThweWZnmgst3ihs3oFV4K2
ClZyhA4AaRJXEEkCFZkasicovBS83XCxgalHCJAt5HfCvPCgUDtA07rq6u3no6xEGbwQeNWpT8u9
Cgb4whWFGV6uFEqJKqi9N6HhyJSKAFoFZzPnDI0andJz0/AnUJAPgY9kD5zRqm9ievWR2XAr02JM
XZe8WQLhDk8fvyqCHsTbKCUkMPoLDhY2Hu9vlmpIBTo0+cuhuSY3l9NIFtu32m09C/qfvs6al0ld
edSz9mlO0S9tDf5q2moOmKtV3O+3exP4hm/WZfViA3rhnshZwJdHW+RkLsnt4wLfLK09lRq58JQ+
g1QJ0O0wwyEknU2MvrQxb4/h4NSU9bWdWN1ejR0dG3PKNKw1DMeJrzaTcjbCIm5I+w70Lt1LEU6e
YKsTkv1pqPquUxd8EbVLSRiNac0HaktX8IyK+an+VWMn2IPHw7pS2EDE92BsJEF7lpwcdqHGXrtI
eUP5JJfDWYv5njf6vbeFenoEsu9ucpRKon5GOYpXE6M3sASEuRc0pU99Ub6ofUT95z3L4ZFftaCc
1yCpnaYDoDZYMsgPK0T+FpS8tZXLUs4HfdPevnI9Ouzd9tDQu+iSEHc+THLNiziXOGOnrRdZuvCb
keco97TnTQyV5Mo/LAOyf80q2BNe2cBInkGjnl2SvfO+eeCrn7Rb1bguzJCmeUMDbM6L8vYR7j/l
JihCHuMLeriY2FGBV+U9v2Ni8Af4z83S6o4HV7g4WJPztv81IypEu5Ek2Gie0T5JT8PiBShiJLsH
PObXR8XYVqpyVHZRSAQxUSizDibHUZ5SOc8aOnW+bWfa48RKHcWsw1EW64zri3oxaB+M83ziqT/B
sbm7pBQ17RKndVgU1FlpyqBNz+iWkqNmkpN3z9pKZ1KhjPohawIIdusFqYOdivlGUmvhiEieGOJG
0+7Qx/ow9ZlwbBqo+4BziWos12+s9nKAHe0Bl/LqAReQpztRrkf6MycOKVLnWDUaoff0/j58CSwU
FyN9Jaob8rHsPIYqIr2Fb/5eTfyCrkKT23pAoJZJyvDlU0C49Ntpj4LngikzvCOkQKgF21sWTd6d
IArTMjUhIqPVkxwks2Xg4IRXvWmIiyGQeIf5ITEiciS5UPq5MBYJT4jtMXR8ep+t1eAropD4jOHt
4J7/fa9YLCoywdYa4AyYGXwnVQK96zcqDiB/xFXSroWw28ksaxLouEEMbO8BO2Mi0rJJA2v56gag
hR5t2RnOHCDbrq4YhodPpS07EUQ5yi5a6Oj0kmmEpQ4vfb05br9ZA6dFuFcPL2TrwCj+OGHXfP7h
46q+pDP+OKJimhAbQGTjZQed7NNrV/1bROLSh/5Y+8CU+EnIzs8ZiL/A+vBWvlPQOj/tVAf9lz5d
dhGxmuWMcRN8JnEDMmdggleKcseNWclS+PZ6pWnM6mEG4tOFaqBwa1Mj2PpGA3W46JqF0EsjFkVZ
I+FBG4r4setSs4acJz+JNmuBuj7IWNVklZGqWJ95l452qOhHqAw2FhmT726rlwhgucVMtBASkinP
8orF6DOG3cqX0ZxKXlleh7PVMVYW4P/FMyUKet3VaJ3uPV2GlmBd8BoAj15nDmKNWSJR3jBICI5o
UW9i6HIl+kUGMaDoGWsbhTyBZ+fD83RF9b+v4aVzUWLEKKihkBJjgsjBmyrsH5GikBV2Bz6PuvWa
2X2GWxE50kOWCOkvFT1QNT9uX0zmcHqqvCLOCRzoTqLFhIH5HI0CdpfauIiy4L6ovgO1Dv52DFzE
Y5R+2KdvcjDRYWAxMnQShWhmOFfhWt8d2qnL5E/GGGLtj9zIN5NqnxMXKBYl5RVzp4bXpOp2MzAZ
8sMWLA8Vq96khq6CWAMlnQBWplNSpSueR+JMfxPTPOCTce8H6b/lApYyoMMQ8HhAV7z/leuSPZSK
Gp+6/Nzw9p5R/4B44rthGGsb2hG6kKl3fSdoe3DaJ2vMF4In/lHoVEYS5eK6+dC09OA4ntb0/Zcr
WPj3qMyZ4WRrucsobSqOCql2oLEjZSSM/7KQFYqhWstgf1WW8rSwHQS/Ov1Vq6of+QnOv4XxHviQ
Byq4dv3VY/osQxen68ilM6uiX48a0sUlE1jFomQ1zGhDeFNKjLGLuORtZMSiDOpfrQt6CPtC1/TR
n7e8wGHmqxz+/YA1kGa6oPyPrb+qVtlCENUcjqTpTS1gQAzMosOFdV2/PS1yPbs0wlojsFeCR+8O
Ky7pi99mq+bRirt8YFbZ1U7IWs2OTVlbUI/13EiR9Qd22k6L7Y8m+z69GYa9yyNQM5k4IKwb4v9E
xu9+pkniJNwtSgCd/B+KuKak3tr4EF9aEkBIfImwPbAvFTthh6ssBlGky9RJGLTRZHvF3FaqgHWa
oGQy4O3KllR6NTPfrY7zKZcZ06rn2KmY9fY5XF4Ve3uRO/7sLEpbokYPVKG8KtHfZbk17ofPRF5d
zgsV3nfnN5h6B0plxU6iRt/M53em8/km6WAeS4yQDvNDElRjh2qPuBwqpL2wJ1ogpJwS8aeVUZ4c
n+JF4ogd1Zy7IGcJpJ+XpivuEv2l/+tXC9SMGFmiLLGWyb2LQc+68ia3uRh330Hg8rWBV0A/D5/Z
mDCMPwWGx2hvsR27vn/uS6qwSbWmlGJ7VZwCj/paGoW5M2E3ngJwQ/RzCkjyBpQG/F8nIMZBXQv4
W+9PoDWCqVD0fKw3vr1gsfNVqAaYckF+D12fP78o7VoxlHDw24tsz+K2idXv5pFlwVTlYGpzJFN/
X9AVcB8M66VtGVgYtvEemDwqJJaqT1DMoeqfsq6YhRiZoHwMNNnGWI6IrJ79iFDTBlx/0MongqYP
z9X1QYXeuj0Pz2C4otZGAbbzGpXs8RCcdpKKJ9iad4M/ur7OEeMFcwUyY9cahqJ+I5XInJxV76Md
RnOFkWDFzhhmBiqnPkqbgiTqz6bYYjYwhyU74SVD+G9FBjqf4u+P/8dZYzx/ywv/cuOs1SLzkVYM
fE2WaqJ6xE8XjaV/1AJvy87gbiHAICAl9C3Y8NQXbDOJglrcIjYaBUCD+A1UMfWSH+BKIdLd5Hqw
0pwn6qJ78cGbgYiyrdGi0s8GsMXnWZ1GWHG0v03LTBeaiaKanHYdC0NHGrNoPwykRkbuSyqyYTEq
Wx8MRQqLC8xklPU/AoGjhepFt1Nl5uZvSG0Fn+afHqSHtmdn/7xE+ZMP8DCsfg96Rz+An0D09B+F
ke/DzqG8FSVS+A3qjWfhYnEzQYWRyTBsdcZuJ1I+2SWveSL/wjbxYRDRUA4DOUDM8FMFH8tyd/0D
+awtzR/pryyjMDIF30kQ6jzICWNjkQ9tbcNJYPx2UYn5cNvF5LpTUPRpSRfWI21rwK9qy2VaOPPI
3CRaGJ5j5vnr6nkBtSIrJxUrCBUuN8XyN9var5BaJdh6NSPD+HvsWeL48sZF+AxE8Y3Vd+ZldbmK
9ZaF1CFBb9DjTq+EI88+uLVqped9TdueWkUcFsf8olpbpEXTx7IsVmymHuDYuIWw1eDSfZvDoQJP
AVptHvYoUlJg5dXJ7hF9JupYb/YQ0Io/POCUlWkjHXv6SqnbSaZVR5i9inRcKBTTf4Af3STMDRhd
hnN+glqBMi9laf3BN+cDkSEoEJhb9MUHVeLWaS+3+V/u2MN69++RlLzmxsEZLEaIUPXX+Le95i+F
hxcP9oXhzxREXvsfxftjFMES+yFfhhbUcRhHpEh9aWx+mi22/V7G2ZVGQEwmAVfMgyEYPE0r0veT
B+ib/VPF7H7loHTRNbyusTvtEpqzvBmVNNaYdQ7iXFonfOr1atXIFXVelabWTbW6s5GrrG5JmoUc
vvMIkKS6X+6KI5a4RI0IQIi5XD3bjyVbjHdvLyMbkqzcLQOc+D4CeawfnaZ33mr3uWSiZRRbLkAl
Hhj6j/+kN36JXSjse8qNRUExrN1eJvoVPARn+jlkrkhNlJJKTzNAT95e4yMO0A61Sny96Kb2SjwW
4nU+V8xg4MFp2xEhmxEy0XvjpfnmY468vyalJF6Uw8dexiC8rnLPk32lSV4THqerTYQMyOPJsBat
a3m0f6az+YC1lQn4dnwLEBtp8UQ1vd4ax1G55rH6metOTYWsCBkrjUoAtIONr8WU0ofIfh5vfkVz
cmTJgH9k6QWF3LjHJIYnghCS5VTNDL7Yzx9ElsTJWAJkDsrjTF7KFn8MvrWPDp5pg88B5leUHIeL
hYvLoi9ZGI4y2LgGoIrDoB27neIE8fOneVDzg+stQc8svQl/Hogd4yeBKDx9uSLR0GBYQip9b8zy
9rf9PSyQ3Y75EqrxULAV5PNHEgY/jNEQTLVnvfSYDry6k/Z2zcMqsFRP02Xz2u13PhJyOo1qJfMV
NzYV71qWE0aNRZsnk78vy2Ukl3vbEzr8DnVMScc0DTy5hyGXwKSl07WueTyDOWXtVXy5BwkAjDyY
9nMWZ2/uEskUb6/KXjaQkuUkgSRvCls+JIDA8U7TXsjbC0dmx+V/1pHO9Y9iCrpGVLJyGM1cvLFu
9LwIWZYWm9KLtSdV9eiv4I492ngpTpwmaLI1a6hDH6Q1ANdAgcmnkVBFoFN+UfaIhN21YWxniDcM
eHOhoQDNQR2Qw+b7GFWMsNmsU8X9dxzSfXBuYSTHTNqzzNg6b+AYWx+HUe76o00VLVS/EP/xxYFu
aGNvLMaD+Xv2kj2lS5GurNgzA9cHnI+342swsSE9Pqvsfov7Gv5m0FyG80JEGqxwZv0t3tvYJiB0
jtti+APxFobLYgmNluJ+9MDkdUtU6N4E7b5LC0pkZapbzmnyhejYwcV1CEVTFFlgqk2xxWfeTzYb
xJZctsmLzAiPqMj0CB16u+66X7PHYRbmIUPpcfINCTtiedg2ms5c3T6FzXYFDl+d7YMk6RW519CQ
ChGx2IgbEgU5leuJwDthgtRJe1sCqcasmmUGbdRyZW1DAx6H4W099eVvXFQBaNYkcb3vrRa9+f59
IVxfzy8vurfdInlVGEsJzldF76XzISgJcJkwasklucIlFmvuDjFpK48p1P9iW9eNl6RQaooqNkXB
JAGLr4ujR6IeGCmIfaKfeJn2gS5XvSJT+UNw6G6djchF3SeY/EQwaj0/Yrw2+riQVlrg4YcN+HCn
qSsSicvrGLPRkj5Jh3LoQulZNcESQPRKOX7UqHwp76y1bY6jd2kIyKJuX1cq7x7ezRLS55hFj9rz
fwA1k2FkQH1bGcRraCoMY6oTdJG2X6cs3EwFy2Xynfk3ETkY8sNz7dJxayKXoyep0A3YRLMe1QKo
zHX0D/pIblXRc3JZjJ4NJ7KgpsSa6xjLYoE0Oz+IM6wmuGCfrXKkusBcHW1K61bM/a/9Mt3cnS5D
jNIE0X4QE+nXSs3Z6hAIS0WRsgVoetolOf2b2UjmTbpCz0sPO8GcbxCdgb0tSZfUuzkIMsmMP6bC
juUTh6eRGmauGNfqSr4WP/SGJfea6tJ1G+zW8/8fbY23okry/EmUcqYBCRDBfdxs/2XKpbshae4D
49Te0HKgmBT1L4p2Amas4VQZg3kLYd+dQNpguwHcSbTpupCWqkkoAonif8jjWceBEGlU26CM1zCi
noEWKqzTMaonssJ6ktGdhv6L+I+7bA6Mw0CizXMrJj3gTHcla5Z3F2MCNZP+IZ91SH6WprfTycS5
MVY6FnC6wdrsN68Sga4rfSrbgRuio4mhxzHL/KNjB7HRJI3MyO2AJJciwGBPsB5B8EIlxNMtP4kk
hsfBYdUJ+Tegd6l8tNX4J6dZgNoWSOjdzaM33hCjRCoCyVgaYSWmfPIwnWKZt7VBrnxmsnsKzn/O
GX424drOpQ3BDEwuzaCJZGE6m0SSaGdbFc7IHL8W6HsgjVrJSw2KtQLMb+RvgsPTodM0s7d0n1s6
AY8kRBb3DK+48yTzNG3Mmr6R8/799i9BfLBmaw2mF1tMHzCCRyPO1PyC9jVEnT+4U6ZPNu3Y3+Rr
goBjSsNcdXGN/VL3s+kDQ5bu/KLrJJOX10g6OJNNZSvmkDb0DEg75pKeI1wwrlu+WSX7QVc/1ELC
PIZYhfoUuytBZl/dlOEM5FIjm4Qz8Z5+7We3FmSVkPy7OJgKKiAgdDCPWLhIZazuGCUfrtFMmb0t
QehzzY11FsttbNuTb9O8XgJsGQ7va/VwvGxOpIZ6scHQfwvTUCNSEKxGedAXGkYU8VF1e5IuviqB
8q7Aga6JCZ+Is8baycYJgBjnvTE8CA0sZyZW55AkiZ/RiC7e1A2z/+D1v4qezks/96TT9eZsCUZF
10hMACdSb+lChC0p5/DhwlzZXoieAx/p00sd31zH80cSucy3thjDjm/YuK7THDL+ibN2PkiAlK3y
njudMUdtgNNuogSI2/DOEJJLSDcKJSfo+gFamfrbLwSUDFYQJ4utDs1CgvoxfuMMYz4JMc9Xve4/
xUBfhO0ndWyt93hDOV66i3HH/VkQPPClQydkh7mohj05v24UeJs4YGrxKLH5tV9ua+RPhvqGxLJF
Gnr/1yzfK2lYqNuizFiWC8Bc6CEwZW2wT56U27O11bvsLPU2k4pTmxFMeVx9m3zC4LPe802zSpTh
J0EAiow95DeAUDeev1SNX1q823au+jDubMa6AUlhMMu9mzKi1vg2b0N6myXHHw8uMoE9GLPoMDED
wqLh4wikr2KRaLkgsC0uXyYnCKU8F9HJXZXS2amjm6cgBZcmZpQBNpx5PIEOQEV9CVPq4Ga3+vHN
IuTLDZtQ3o718QR5ko+Gcr4oG3w5eIuI3nVrYwZLBnaDAYYDBBrbPqPu8KOowHRO3eETHtCTGYM/
4cey5TpOulrSn/EARQRtWKbcZ6Glpxf4ppEqJH4uRz+NIodztRnukoglAAAVSb1mnlmMP7L3qHnz
YeeQNGlswXv1oz3pbuI2o1Pn5nW+GqlFiK0v2yoMd9xRdX3eGivi10HWpAg1M18D+5FDJ8HQ6RQl
oTx2xCVFlFts0G98msgUvy7c+yoot036B4JnAjx9Oi4D84FvGhF5vjjH76c9XFDMKPzd51oGywIw
xQH+aI/rGfuz6NQRm4FKmo/eTgNvFDF4u30k9uWN+m2MU7a/u1gTQTvfqaAl2aSqF6fX6tES+eho
u+xOAhgcW2sO3ZQSwMBeRq2tV+j1vKshsVBD8HhU2RmsUuFHSyDbEfBVbzWzEnRMNR57It7jb6ac
rSHrjRixTg55nirPaqKowmGLCbW4yyJiPG86c0Fm3mAXkrr+cVZMO0BRZJSKBp+gUCSo8pzl/Dbw
0z9V/19SXWayGagvTLh2uf7HurjOG2vpF/FfQKwXrskmAH8egTvBRsowc78FLbnFEs+7e2/1o9By
bUga0LY8jl8mw4VehCtwUWIiw8qsVbkalk4Fuf2odOp8lThuxIV6X8env1hwei0+Fpi3Z52MxkrM
3dEcOFaHPOILW4XSc7rXNHTBVSqFuaHmKqALUfNmdyZLcfRhSsz4AIOsyO2gi3WDQIJwG+o8RWCH
BMZO1YMR9R3aIP1wqbqWxKOakDkuvH1Fv2JSLorNxyZtoZkAxUGeXNyuUz/qGOpNQNEFoecvsMfk
5LC65i5LCP9nL3uFA6VaPPj20xdrzczLQEcN+9M4/N5zThvSW4lQToZr6bLS60oZTAkOF64NHqrh
eIuiyBKG6DVsW5jHeHYez4BBE0lxJUIDsw0ECjsPKjANWFK9g3IVQXdhdaQME5UpZ0+KCb8n0sR0
mzp8w+qp9sN9kkg3JjoKiaM9i1NuCFa/IlmgwYpAMnNjREEk3r2dRh37G/Ai5HO191E3LsicdCi+
XRxrlLhGML0nSwKSHc/XloJb0qQlN/xWfVlGSsv7Mr24MGLqB0iST1LJbpBnHHCJUpa6B6rRd6uq
1jYYvCgaTtUdoX7OA+ybJkwiEFh/nUgulpmncnsMqBhLePDHbQ4lneDVytMlgOOUGRmAcuhGnzL/
ErkfuQU51GEDW0jr9iAaiCUBsCAi3azPYNN6JCUXMxPgEuH0fQZNoWXKlAs0m7nY4L3LFscu28pV
ubup0t1dP0OJmFeuJme17/L8xAMK9wwwufp88qA1NkscAiMfXI+fJobpYF3fZzV561m/RULYVIWy
0tA5GjqIQQWMJUNVvkzqAQ2MH2RyNZ+ApHF2vEGbpV4XKwj5fBMHLNGx9hjYvY0MvjEQMQ0UeRNF
U6uEbJJgDRfvwcAa9Ls+sJLg9x79WMqKTDIvqkmx87z2UcYxRbiFnTlCmNt1vvM9mtVyfrQ9BG0I
ayBivQ1vBYZyXrU51p5bPca71ku6UvIO7a3SK/4ji/9OA/nyk/rxTUtKN239GZPy3eJj0lbuVtXy
wpjm7wWs/7OQAeH7zdvVUWIo8FeLvrQUou4PrvfcYX3W0JyNTda7PYxGso5BR4HBNqYlKnkyQYPo
rVOkjBFDAgPMoTIu/wx6qAv97iF7atrnXjiZbueB/r1g6uo07BYm7rrVaJGE+LBDCDEfyvSfbaXf
TjL4K65Fk+5/BYnUW3Oz0o6kw585GBwbW0E2B1/yS75KvtD3mPHyM7bMOLHWesrPwnZmtE5QaWNi
OwBKiM+G96colya9C73FzB5pIg+MZ6rKqNXTZz7zUw7ora/Rrz1M6KPfElky0lc/EpnxH81VAQeu
Dji3C011cfKjpjUQdtA1La4StpevNH6TzyT+94a87lMOcp8fkEyUKTTqqJ6PVGyAarmhCvQ5HxTl
MWZaszYg+P04DnXZ2l0uEjoZlrKGe36Eb0qgt2EgJ/vPDiP+MYfXHGDJPQnvh+duwnJiYACubC7M
gVml8vrURBSe39IJ3PIP1JIKsFBdagi3vRAaPONLsWQN7WQk3uSVguAOLvRdb8BaYfxxbwKA+1NM
51x47dTPblDG7UkhPGjCErjWAEH+p28uoudyzGBh3FmaNmro3iCSCbjJzzGp5N4BlU73EKfANNfQ
GVyLVzDspkDtol08t2IzXME1V5AOLhQDkCbbq4f0h0bMHrJriktsY1NZeD8M1vO0u/PJjMpe597j
nxPtwJhaxowzYocbDwEB28FKfTWkDsQQ9Hz8Duh2iSM0iUUNBwmfInF3Uh/6VpwgIKYWVXMqZMI1
rlJmQUWxNibX0F54p57qEQFhyaxQALoblG2VIYGvc2ZOacWhm/EK08RmKLGLGNYEJNTs6v78oRAP
tRmwNjeDuS6Juakk/yzqe/g4FhRx6OoqWSSYphbFZv0aJicR73ERj46ldK8JhM+h3+KhYjKpDmb2
VJTsKYGZQVuXG5Y5tyZIHQUNtsavGMwBp7mAdHbGYnNHpa1Lde0H01xmG4l3iFD4p5mXMsze7Ycf
zRst0oPi837NHq2xwL2NpMW0hNBLKeJp4QjRauNFiPBjwhKDEf2KMW/PXplZDOYME8OqdK/WxHhr
8aN0pDSRaiAF+CWtCVHhZfkxC5rR/DBSKOgIK67+X/4DAfumINLlk6cYLjR9aGU2tc6wTrlNqOEl
P1moKT9REu8weMg1TSw/ACuIhLjCWSb4S8EhRsF08hfna3fMI2s0DCwypKAm7tuKVLDE6wirxIJR
XN9AaYLsOAcVNoQFYm1b6g1xVTKcEm0iq6AUaGoSV1XGCzclBYTr5quz6w+Rn7IgZcURvUHUCHSI
IdjwdG/fqqPzfqqWX7qVbuaaszWyR5gn0Wxz8GrwXWCdbuVjlV6+4wdPK25MBdVaP0m3HVy9C+4N
uTBjlujhvP/Eftxz2UMs41eOQGUWUVav6DJSH3rydXD+sy4cQO9NwbghjtGWBjE3BoQVTIJCKw5t
DZna2A1q42SKSJGKMSciqhuS76gB+v98aYLEWd5xNS73MobZwu4E4/JZPPlFjZfCNhVguNZ2fOqn
fTVyowU/8WWmfcGXffTJKrsHIdQftXmpcPrmNZ9AN6OFQS8qjpwuGU/UbPg3csshfwwGkuMQL7HM
DeGEoF1zK24Odp417NVYkkvbJY1gwhn6rxEHIW4qxmTeiAxBgF068z0oL2YJJqbgPzBCLnamcm5k
Mn479WlzeokqfVoqLPS6JvFx6ZCYbkfn4elGu2NGzsEQng/tWK2FTFQvzrfMZsWk9ddlfsx4o6yq
LWjCal+bLJD3XEVnkxPOWXLdqZZ0S38qBiNtZ9MtQRpc64l9chTn6FihjoethVDH+EnqPTc9XMyL
TKe9Kl+06FhuM39wBYnageKYXW3M9WyA6iiHGtxnHFrypbc+xdwZMyVejINxb9UljEn1hIpG/EdG
JyGLeFbfVeSiCTH+GP4thbIcc5BcgAY1sFtlbgW2+35Fo+26hHr++KCf7PO4GzTqIMY0D3o9fnsR
efKUgRVMExjZDh9rDm/pPE7tNsh5Rl67rAu+QFXgu+nh4rQ6/ttixe2D9mdxCTq/iYlhWrUa/jj6
o8x2AivhoiR2Svq6JRCy6ZdfrY+aCxPBaO88JHsQU5pCgFpdKko6r1VlZMU52s0Nvwgckku4SOBH
b9rfMEOHLAps4iCYUqdoBDS4b/vzpkX5LgF2CDNDB+o0wVh95EEbNXLQITCLFUzBAlOsj8cLKygT
c3Ku2wWjHtrgvuPUuPq90RpzDvNVScuw8HaShGoepq3Kbg0WSoRCtGqjVCKyPGjjftsYtOLAP6PY
MdxYzJGCsvhol6J8kfvUkawPZGpjzdOxPojvKMni5cyUe165+CHCiFWhGsudiBbV1/uAUHQPR+O4
Xj22GPNg0sfkjOCbSvFSvEIQ5hpIbcf68R5qo+8NB855oKobv7NgL4iSCtk+pLCsOX0cMZTstKbL
a+xtuzrkH9mCcNtOziTpqaT1bEzRgJvYmA44mbstXuj0YHFf2ub8+J55lcPq+pqbOUyzXkq6Qi13
ICIL25fNogIdbZlPxwi4XfrbLhTwqKHnGvdhyqW8m6IbR4HF6bue1GeFB5MGHjaI1Qt6Yop6aqyF
sh0WjNe8JOk1XIE0s/kxcZgPA7n9+zjDpUKr36RERep99EwfCAte5RKQnYIJeoerj1SbFMVp6tet
bZHDeR9hjfeyn0Ok7RSSmpmrdz2VdJ14hjRV4OJFPClol5/yqgpi8ilxzm/MbnIfVNkmY6F88QJh
paTv0JVYlluhXBGEuB6a2MsUM1An9nuWoTVBuAV14/425j8QsSHsxwoog7/BrSGTI1RkVHy3RvTL
y4OWlyugw8ySlUC/ky4AZGbgdlCnVLhb8Yn+Soyjzs3DnofNdGt8yYerCl/keFL0INN0TiH7INNU
r/dG8oYQwtOxJC5LEFWLtMS1NViVU8CY5m+6im6yfVNajWpkia470HUrwNsg3q0kxA6Ehxfe3v8z
T9HUxZJbpf4S4lp81CgaOJ4KMk3b24aTdZlySYrNcrzrYAzW/XyZKwisZG7u3FUN74U0iBL771kh
eW2oGYjYLBzHbSC6eY9zMdERDpBHcDPBqAgbkP4H2XlS+Db/sbom4d+HIr266eePyg2NpZTRf6Ol
cfMgJ7Jf5CZtxbJ4nGKqNorqVfDqM9IWlSq2XLlAxJbCAl26d8fuZi0j446fkjsjBKIqVB5S79e0
/7K9nI7qi+gcDW0E6XIHO/QTWeZUOTFMDAAPPlhWLkaR/Y6Ygq/Gvimkw+Q7Z1OiDSL1S/uxO0xx
GYBF9wohONTX1hpsfl7vM+Bn66/lDKTZ5BrsbOGsk9VKZn2fzxBOpovI70ZhmZJj6qUeafRKYaXr
xgAkanFDzkkJ62i4P8j9n7EsZbY63TGKEjpN1qLivI+vPKf6LZ3EriZfuXSmDFBod/0yfupQGHDv
+WWKxYis6pDu88iXoEHQg3r2A9PRa3DLrYCBZoNu2fJokba3EafdbIoCtFuJ/k4VbZZjxoQ7nweY
kMmKynTToxfvikoJO8E6e5BxkJfUufzY1aPrWnt802eEvn5Mvo6qZYPHfKjcVtiBqt8I0Oy5u9xU
p17ETy3DYBqkjKaFROejptH2Dcpfry4qKBSnS7A0ayfP+6eDWsgq9BMVt+FqvGbx1khMAoWrmjUn
WHsR9ZHcCOlSOGVoRUvqbRsc/e+j3MirtIgK+xPNPUNhg4Y6veOVEKU7an5CMom7jnul9jFehVwj
dFmWdoVBO6YtYHjf/fsUO9I1dQbG9RbtMRq1izrKBCfWZk50ufeUZ10V0pmdvygH4fwggGbJqvpU
qlbViEJXZcN0nBx52aBp8ayvBYBQDtClvrMFc8tLNrFlrfRvn3lwgLaebuHphCPQj5xCHKOzRvCp
GYwZjVgVaDVAWZPJtatDLnucLJepyZZSSvGJxzFP1C+OYDRoYj3Nrd564scuTV0DTN3z0DtDBT0L
J2J6fv5LSFef5DifOLtvJek4sG3Nv6Sup8hWP9n/cJIYAShBU+5ATn7gVOfDdDD0byiMerKkd+43
gQtVX8K0Ynv9rjlwUA+J/lHw2LfHUS8i68jAYTwxkB9cItZm/BG6QDXhhBp11w0pF8SoXu/EvOpH
0HTm7Dj9HX4CApeY93DKbUTK2Et2HkA5W0rkOF7kCHw6eABcpPJdE9fbKK+qlS2CQYGhHMH8jrfu
IYwK+kcFkVlcnyUzS1ea7KkCvQqmToWO63HomjFGUgsbdJ7h/JdCxwF3zFxlMmrHRgLGnIWhA//H
FtHTFzyMsnQtIySFcfNEyXSmyYee6FQOV7ov4VyI5+cLj41dKIoecEaILWqyBb0BwiRdJVVS/dh+
sQH4UA1P7xQ5r6hA7GLWjpM2HWd3yGRz3Rpy294xm0itipXWar2rHorwLEVA5Bs4Q2nnGDbbaInf
gG33Uko176cKbdcWXm1WTwnIWt4XNp/h969gL1575rX1KICSDH1acOh6lw831/UOMVX7jnVqcERU
dClLypT8nut5Vdv63EcDxWEmZXxzuLLy3h9rq/zArdebXhEVwXRF7AzCEEgdkOE/qWfvtQFld+B9
4xaHfqo4+X+PS37aW4EVdQuMgVBTa1NY/tp7I/4Ke0+P7raWeZ3z4gNrVxobVZK+nrBXtAP2j91r
Fxv1Fq5mulp1f7JhvGPOd+HJ/77kLW0xwSwgyIw6srjzBaKpMsiRUIL4cCv4M06AiKTArdRDWNKJ
Hn6Grs5qzhD5XCGWpb8Pusxl/LhlTXcVsvF+4VOi806OahPy5Ezo8g7AcJHK/I1JFA2fl1fwuK6u
VLItORxrC0N3OiPWx4ErEVk3fXPjLRJQr34y4mfKBUNr7GALXmG0sSjvkp5NgF+JJvnrO00HYnjY
hgI1pMOmDnLdF4t1/WJCALDx5RENB0fNFQEJTOK4n6zEgeSA9EVHV48AeBlqfpDlVCLyMarxOrU0
XdJ86VbQsnyKzm3LcMCyvoaYCiVpHGJxql5Ac46RD59UG1IvB6J/vYXN6lA9asEPgebo8enwy/Rj
mOKNa0QvgbxChQpuvUZLFJPk6rwVoKfwjgZTY5faLEMCAvpp6Io6o3enicQ+1taFseaUBpM7gEpy
fwTEJEYSalBjJNTchadkjuw6HQTyZRgqSJkRkbP1Hysxu6H2NscLQUziKCmtfldKwwLHMIYXHJ4F
c1o9Ik3RHfHfoIH2qP4B6d28tRpAyRfoNXQw7t6mdXDkiExMp+mZkhc0k+U4eO7+bLFMuOPi9LnX
Hu2+LWws0RlKfgogQ2LT4E8UD1Szs7rrUotaU5k/QrQl0vJ1aL+VfIILRSwJuxFRljrnvVWTH4Up
27t0WQ/fzrH20rBbBZRlSKXEw5WBgLTyeEnDBgXmC19qrsJi5ptLwxVRFI6xmqbXewFCk5URnkvr
XJ7OmXBj674D0OLJIHmoolCVP+r0AACGk8dz7Ggbtuz71zM25xLzebFNM/d8xgpETUAseBmtNXbM
9xGuS/96jHSg33XzVgcnpxgkInZiiACChKdJUS9/BIPVv8R8xOZame3NLZk7xxO8AhQBVsdUCt+w
vCPq57w3TEBmNXyagzxUl+F2umVTc9dK2r4JI3ag0eAKf514JiBIEb2kKI4edwox2UgHzbnqadBo
8c4IoxTwXxNKegZN9RZHtrmK1HAjTiExHQ95oaohMKQ9g8R8yGmhvXea9xlUhDR6UODJb+fQ900G
x398SvGdchEr+gy6dklUWulyF0WhpGgF9a8/uJUpgSGOoUS6sSi0J+7P4Egqof0qi+pBH8lmYbBf
N9M6YaA4rYSySmx9VzT+PjRPuY79gZGKHRzDJwpCWSk1qN0xITj4v+zeGLC5eDWK4KBDMrARgLOA
VadBqzagaJQMi45tYWads+gG5WFM+xDHXTg6OoNTGBFIYlMCz9jMBhHKQLeq0VXu+HafjIu/sRq2
9QBMZpAzVne2TNLqRhCqVZMIrkM91gn0V3W7hlogT2+mo/hal7NxQsrkfoXWxivGDDECE7jjLs7d
24QtBsNDdUQ7V9Z0jZczQwy/qxwiowkqgJAYKNaC2dxjeFi3N996LHrMVtXhSvmungDcJ5bbdA1s
XiiFxBrrMQf3q5KG5rmWjn1xwp1xh56sNZGc5nZ6GqLVbzPMlvbpdK74QCnRpY3fqSIMBAnF5pkP
W3PrFJ0FFmoaL0ox5YNNILw9G9O5ls672rzwMNWBXzjH0Uz2krtu33H/gTNCiV8p8xrh9uWiMEW0
v02+EkTL3QirxSfTMFivIAAemjVrictZkE0A519V/Kn83y8j4OIChzjpbZ1t8HAC3CdEuhNITtsU
R75+6iCbDI6LLf0XM4a7nJm/bvEc7WWP3V+o5Kf5/20kNTkQPD1I+ly5Ln2/t/4mYLfRC0hpQSBU
ophacg+6OORKSi1xa1N8PJQmy4ChEjNgIsw5BltERnH9kYu9DBKAcKAG7N2UY3C6CcTO1ekKIlfn
UFO0rvNN/T5Gv1Zr971KdivJB7VqarFvU1Mz12D8M+6hiwZBkalWFCQZu5EnYHPVpamOT8F+SgFu
rNKzOmQg2f7jTx0h7ivOkmDUInAH0t/wzlWJVHZ3oJByp8B1uuzxEFJflpiPZcSKmBGePnC8jlWe
swV5B9/YAjsTpZz4y4PDRa7aLWRI7r/EV6/VZKiptjhrwJbdFd5CdffFkCzGELnWNhA4J4idcHdj
AYeLfhQN1yMwWWCtaajwnhpdWCvn35a1XqvUXKuvB40VEgVUwwBdDrCIlk4UTKFGUlRmjEs7j5J5
VTuAUB8LQqFfhxy3yAsFC47wtCRpm4S0gXowpgJqdVOPCJMvEUaIenzmJXXfOWyo9NAyb+Uc9Q+1
dHM7pqYrV33uviwefIXxS9s0cSg8IICdtbE0t+o5+IiarkNYayubsMFB53N4YL23nVjHmT6+e+o6
Cqdk2vz3mIjn3t1pxtxSKNNguhvbgstEjzvKs7q6WC2qG8sMwG8duO246wjchT96rQVYoKiSzK8K
/MCh+eqWXmddi7SBwR9puFgSE3/QfAacb8GnfU5ysQthva1Ferm8FfcRMSQiUmlXqAizl/Pq+l2O
JFEtzgZaNsX23bR4MyX7KuvrnuZuq6Nw1nU6xDqFmSkz/F5L6keX17hZaeT8KhnpV2Q1eaGXHDQD
jnVfk5dhstTfdjqouQHunPEYVlYRVhFEaUKzTQ9wNhINGqrILygQ982EfaMVFyp95KBIsv/ArkmA
/yRZ6OkWc+g4JQ6j7Ml6MCsPY9pRheFm63GYlkuuLZcNxNbdm44WDWOsY5eatAACO9YsLUCF0Tg+
Lu+/gKrpq99JdwZ5tf7yPcXGefPA/7McFbJSN65DUillA3coGU5QZXgkQcju/KoijNqMJTDOpb+B
vqN5g19uFyAYtpE/jA8x756KYwMfI9g2gCk/JrVVpAxgUp2Rowwe0sct7qM+n7U17uN0L9oj9KZQ
/+Zn191HhYF9gSd9Xm5x04qeQIWbSkK7C/FdBSX+OyEZeVK00TXuBB1IgfrRaA1UGfDaFuIDLsG2
rd9sURWCNUY6n+TqaQv8j5IpJwH90TdtlgrRqJJHPuyCS2k6BO88Md+oVfCthmt/yNFxmOtHd1A9
lh7u//M7dOjiKieGT//PKdRnPzImS7o0nW82635w+LEIiAsEz0/f72LXLtORrZ1yLvL/1whrV6fQ
pjCNXfxKLmPi3XXg1XqnaHdwdEcG1GP32+rZKebawx2C2BbCf14yfjSqZdp7MZkLDbINrEqxt0+G
Bfi75t+xhuIP2mea7HGLDiXlgS6rF06VpwiYAAsnJNzXFIS1InAtVcH4G9h7nPzdlvICSe2KGC2h
FFD2pefoO+FnSAE2QPTkGKbD00plbVTfq23Ol3Y5taMTwR8QJt0RQB9bvNmd9NqtX37ZCcUySCFz
o1XxA5TcwLPGvneoAmhT4t1YhUXwnnQunB860sAUQawnuwGUSd+PS2M8nG8gqS3STH3ov8aIUwjd
8EeFn01twx3BvueXzMY6uReLioMcfPToejTLoTKAm1DpOL6dliGvl5VcpqUt9zvFmLor0SwaMgwb
whYtFXXxSzCRXBTY5HogjI95Jc53rVojesMx9T7TWxsZDg+qbFkyERgKZRflnR/ZXQwukKfpiLjT
nJvUDtA6cRV174TszN6MMi2TwFcsajOrMKKzdiJAeIiS5IlTKM5DdrQhJIb/xIdBS/e8Wjde4MRk
oPHBMARb7RXUT1MtKzY06Rtgm+URnlA38QscXwZNtq1i3LBe39rMDTvjYrURQiDy1BHABvCmK4lo
aqrSIY4C7PUTg9FLtJqrjYKpk3Yq9ByEDox9n3/i/bI9PkJPuiwoPQVrxLQh6Q11GYv5pPXmHcne
aiN2oT2HIoySnv4nNsmKmUWubieG3EhVyQa0CpvEyfR90ihjlgv2J4DCzvQX8YZbQLKK9I0L0Hnk
FQhsB3Y8iUMvgZ7uleh1J+IogEtPOvsXF9hJv/qhMZTAUhEHVkVT2DtSj5t2Vf38A3XNBp2SgSPD
hvhVJo69YEmq5d2JfzGv1VCeVmx2QGvu3b351FvHzUMOTpGuKr8oicLvj1nO/tqReFCO5dhEzWMw
UVgPjs43gN4BJd+POq7V+6eL1dquvwHiUi3kXC/fz8JokyN00zcKiIq6w34hPi99/aRJw5JW+6Fg
ot5v7Uurz7X0y+6g0bdztgDOKLYMj2pRjVLVYKnBtrvMf7iR1mPALDzbWRi1pXSCEPKcdTGKv2tw
niJMQ9U+K4G3X4ZOOc00VUK30ot+lrPKiDX1q+Scpc9rfOm/wg7dfDMmtmhXtmVvI3exhksSoayj
S5dT8PFq+KBkMIwQVvNykRme8NBpVYRwevMsDoeinLUN6LJDXzM2k4MdMZ44hodkI9qHrrsnhuG6
MnHv/fxtUWyAm8D5otWBDFKHpO1qCEeuGSScxy4bdssRVGUyEe39ikMHJd6q9unF4R2aL+mSXyeq
LdHVvT2wFui33CKYK0xQ3Hg6Ig/pR9HdvIMfx0C0OyzQ8zZ/KK6hP2tJe5gOjDqIqTysNk2J/g5M
VV/eWNTekClNTGU/HPe5JPl7k5cxouB8ESxeNtPuYZ/7+h925W3bsW828w1IJaTFvhizHAB5ZhdU
kuRd6RmCBrBe/MeC1ZqXp8/4iDPST3jkRZ5LBBFuVZG84PhN23zhK1FgGcQ4qqKFKge/qOnYj+D9
uEV54SL+yCyDnUVLbTPKltLRFRFIvbFVbs5aLq4s8uKZhYlrRMF5EEwy+OzC8thxOKz35Py3BX++
ndmR06Q3i6xFxOAzXfJc3H08L9Lgk98a3sfWQayXSxwN3MDlhgcrLrlgIsRaPuPoBTaplqY1vdhQ
a69aKqGmfn31YfI9qGOEA+B5sMzCH5ocQf3bcozvZPwrXR6FMfpnAF0xDVmkSoCUDoF47QmqbU7U
oW5CF+t4KdjdODgmtyJu2I5OknQA76Ah1LtkEy7X2QdnnLhNX9KVcqg0cOJEKWLmGgMcNFb8x39q
G5OxiUnl/bRTkZ1J8kP4rDugTIhLFF9n0BC1KiHjnbHDBk15w3YlOANcgZy7HlvfgxPACie7QWw1
MRu+EQU4G7O8SEbxuc9BiNiXi3ZJLL7rnjxXlB9HOLlkmovFHEvMvAA319tckdWfqNOSt9inocHn
bAW093Hxdp12kn8Dbr2tVimdDxO0H+fFxn8D2+i9js+Qp3acUwzx2iVIhYjMqna70hWPsipAKHQF
IFFgAMRrxXsk27/LzzbU95K+pTHceIALflj0J2D/381vhMGbrMIF2HkGVmE3fxQDJdEEGERbGBGH
zzsmV34ElVp7DsbAzt3inccNtBewASJAtV01wSIH6yAyvU5lMnm6FaUuNyQDslX6+O4SmI0xSMnx
pV+BXXBZWgLSf5SIzsEbHrSh1kMQsTCOvUv/H44buPoVQt+amXX7ZFsB0JDh9uW9TdbBuqKlaq9w
trcHOtgj6YfmW5cEPL9stHsn0mEw0maQQKZn99QXFaoM8ZpGPN5OXo+IdExcA6SYpdpyI4mkFtNp
Lvvl5ABts4B5DxtsFm5jVNAT19ACeoEFF7Wc33ZeJrqWamB0U+mLf0QotVzX+URXFsWJGkxwWARP
5e8LbeuQCeEy7QCeLDplQmt4bMRPYLKo4dqfK0sAlZT8BKpzDZ3T6D1dSLC5qf1RhJ788FSFYKWL
6c56jwuhHBiR7Lc1IRc6dH4u2gChboLNhXEDEeKltQbNMr9McbhFvYX0yZH8g0+BC0EksjhEjMbR
u/HeJcInzt2h8PJ4im7DvmB+Hy3TqjZGG87PoRNZ3G//YpusfV2rk+I3hJ8I1UMICMMAv6F2Wyig
6On2+zyvPM0v7hH9a2J0BZM+y8hXZdO6eZPsF4dv1MUpP2LqjOBn65FeOdUjRq3wCRDeEjZueVnB
WlRgN5gSUXqx7MjEy81QjtREciJhEP3QDr17oVAS+FF+/pP7VMv2GtvCEQI2e/LbU6VtUL78egAe
9RzmQ2hH5Lzpp52Gd/JVsfB8KU0rCOONm4/JgnvPVRzSS53beUCPhWODXCMpQ23T8wcoLtFH77Qz
RKsm/b/Mkkw6YhB6gwd4u8Im2An2WzevvXWXWLnF7RthBUN1oD4ngfRqQDYOi75vukWx2NskTXSx
QdTYQL2vyzS33MQkiTM8JeCKptVcRdKjKJzPh1Ir46uJUxPm2PmQWe4CHJWeKj9dYqS8CFk8YSc1
q93r/XfEJH0BMhCJg4YaiQ5ih+W1yKfHYQWRswJNkWzmlw1mlRW63M9hJ2rou8wtrjRYLiwwsEZH
EWafat3/AGyW3HchdAPIw2tqMBM2repur+IQmwivoJZqpMAIg47d2Fg1D3WrI6Js4AlKdiwnDuga
0Upe5Ck5heuE5zUlCIiveCjgucc3yGgodIMjOMnfXcThjGafPAnpHk+2dk4YoqmQpvB8/pduNIvG
aOO3T8o4pjP40GAPTZj4TAQLS6zpkTQMbgiVlTKCAU4tXCha5mZiF93D9CNjBao5z6D38RkHYdwT
XdKl5oxZXI5HRaEVGfLOJ9UUz3a4+vQfVbNyLQAAF8A/jKWwgrmj+Agc8K7PgYZxkPuROOwk65zN
2BDEy1M467gJ+WFlsd2kONAfYkhbq/fx2Oi6NaJ0j+WYsEP0eXBloCb0P2oViS1GqdpSOTQ4onD/
7nXB8KwHm+C23O9nzb+pZfbsaPoUhPfbwqEn2Qk3Sy+HOiEJBZ47WKh46HQcHxt/NQqvxM2VB8CZ
C+rvPu9oUtvEhL5Nj0ltKVXjU/05HqlczYchgXMhi4fc49dG1kk9JcovHIfLcfbjehOJncRZyBQ0
3oRax9t2JXYqhfSN/ibHeqWq+zVqBE+ZwHm9IRzj3kpQSdVvne0MT4fX14vrvscp57YVi9pUck0l
hxdV623ZSmOlsHc3CkvA0Xzn10vdZcsi7r1noDclI5XCdIXrvr2jYbaK6XfkUdK1+X+JPcfxetby
AvgbFo5neNa1GPPveJ+7Py/FkS32pvrEHA3yVRoyjUeBY8gTYNoPdyvjs8vBSAV6acXiGUEo56JG
i5x76xW8NlFAqIqwbCsULZ2TrDh/uqsfyGZGgv4PAWV/qXCZKe87qs/AYsTaAAlYy156VGG0t8+/
k4ab30fd0087bjRRtQJ5pQrp6Pq4Rb/gz8BBbK4zWpDhYATyU0P4iawvaIBwFMLy0kbhQzI3Bgvo
KE2bxdeu+6+ZS2qhvB/apME6XC6EO8jBAVIWydoAL2SG21NgDhwaEvOH/dwLErl0JRgwQr1gFK34
0AuMRBMPRjQAjf0Zd6L7A4aZ3wu3TfH4x8ZIOHBBbat+3QhK+Aeg2yYjYYVosieIYSB2fHUQJ3t1
f5qa4FYFBGOGgykDM9gnpimQxDrFtW/7X6Ickv8+xyNQ5Y8/aY23oo298UUGb9dyBogiA7r3qBp7
VNxmCtoZilnYrTTwV0J+o2C2yEu0EEZLb10yoTO8Vqsds1CmQ8Ik7PZXkHHXD+XNC9EEgm7WxaxE
c5HAjRvTYMAg2CWAQaMx/by1s6bNsoaC1dPKZPqZvlb+Fi2o3M9dFkcTTDMavG6CkPOjfKI3f4Mt
gNopD4B0rQX2GeX0h+fYGzbci4AdeaA4rcoTEPTJx0TpAaFPGRry9tBNYVvOI/q7nRnE9i8PBIUB
53S3LUv9cy/oWNO+ViqBdMwNCPTbPtzBilwCunfrbcWCV0kspQ+CqZkHFAaSkP4vsyU3b+R2h9UM
LnUw/TgYF7fbdC4XdKem+wj88a/+VXaEOP2/gyxZegR4gy7GAJ4cIg+nfxIGFA8TRmYtH9Cn0pZ+
Q10UlSeft+yu4uCkwjAtaRX0i6+RfLFBmc4jny0M1j0YgUxmFP/6oQgcA/ihOMaifLsalYXnFRdN
2HJIzXw4cnJe3uktoFnKsU7mnBXChsb6+fpsaZxuOqPi+ZlrDLgE57ccnp+sUdUceqzzXNNoAnAG
hMqxVLcvhPPG0JgPsjA6Hcu3rgQKubPXKYewrJYViilwRxKiU1MYssmDky39bbCyTc8L3fAsYnr0
yccvF/UZOe6iBQ+koQiGCGsqymoUmlYop7yxpGgeUQe3FteTfP6pYsB92lPWJC4VpNpVPLru7mj+
xTO7RIWwxg/bq6YtzcKlddxcB3Let4Q5PcfXZgXVPrIqpaDMm3Q7jm5iTwhhbdetzGrZq/K+K1g9
/WbpVDUB6siOAFKZWuIDgcXLGPExTaakA+YYe3LLSBZwR0n7HIiUzfC1d+WMzMqlvNjyinqCK6ev
Vq1kFmy6eTj1NRWqcBOCpmsn3vwC6u0wpgINymsuLaUzurgo9G1OZfA1pqjOohZVYpAPlNbSp89Z
hiBp5Lun6em9AIZAnARoLx3oLq0AbV1me8NFoY1s9UOcZWFSOwEmXvHY/E+iw/m51UvA/jvSo23O
OaXFfJypHsuhdQm5N27ETUfFWzJEZFOXFR78WIp9grpUhaEZRxrhBBAA11pJtNLTpntCzu04V+Ra
n6QhChckvnM8y0NzWS77tZBTxTHZMZp3MNDrMRaN8Oa5xaGTSUvdE2YvOVUdBH3FvHp+tmjbuwCG
NpOX8jD+qN0/HDu4fapGyKFRdph6hiHwLV1F0gnbYHxmFhhW1DvZ1B3/URdDBinUY0X58GP6UVjk
3ILLAlf2JPQ3NguNoIE046aRG6Cwr5iBo4gaBRlJWMCyjKPg71IpBnY/+BWGrLdTUtirltCHtzUU
PjBuAmoDxrmMK1iF3W3qCuV+UOHGcI+XCHcCd2dfFppA5Mnowjf9x2XGaVMN1se2x3c8TYuBd5Ka
+3kSuuxW9R86LXXYTbNTVpK05KDnA9ZkJFo8hqJJOTLv05cGaQ37JzHwM6se0ulRE6V8F/SYKDlW
0WAEPxioXe4wMyDtzYMd0xFwh2Oyz8k6kaCbfoQyGhVoDGJFPjxeC93rKv3KODqF+prQ1fXFL6sg
0FblqOW1/D4VMP93ykyqxi+YuBw/gbD3ktIQ4QBuJdPMJcYxlqAEszzF/0p0En0ldbzwZN8/a7VN
Hb0WNE5jf1DZuAcNALWYtctbSygqDM2aF/APb8IQpVFOgBxQOp818OGJBdu/2eVr/FnGMd5x+raR
wza52+wrBtNEGRWqmwhB+ZfF3rKG+gehbzgxNTlgef4wqlDj/U0rGbPhy1OmVdx7eunwguDEYCZP
HfwYr2qCV37nrsJU5LpnGZMCi5hIEmxRFUe7lrngpV5nRA2LAMM3FaLX03l3Isvlfj0dLz88Nx+9
jwsmSXWiUUMDVVhQGmb6YVOp9VoMPveP8+5LaxiBaNtxXRjh0W35kwsBbA8oYemkvRxH5jrhFIO9
DtXkfylOoeDJnPfUprKTb59JInIeyp0whBqHzXs1PLw6N3JI57yLZ8ft14JqXMVD9GE3+/Snf7xr
xL6hs24P854r+aXe8eIyNF8lnFHnCZ6+qIYekkyMTjAAlsCfsMvJx2O7hjl42sl2i/dP8htnmWM9
0VmGVJdOnjM23EyNRJ1Tp/AmkpONbfZAlr3qik/IytUGF5ZmKST7rkSWAZMW3M1CRlitUA4Y+J7p
Pv5xJjVf3ULvLN8o1LrjsNg4Ic/ZwRP8dAgBphaHBpJrL0bqg+IzHanlTZHxhJ9l5o/Dz+NEMVmN
XccRAGrPOw4G/br4+RIAOzA41Tff0woW8+uuSvLEaorHsjRjcuJLZ7ghFFV6sWRuizwNvxtMyVcS
FLjqHZDE3zE2gUHGnYd5BXS+kty7wthg2b4XuwTsQJmP2bopjmlfpiO98Oppc+EqxiO1wZ5mtt5k
U8Bn+AD9iQBnWARXkqw7WhtJ/saR3uSccdSDUGk1mO7sW7jTZsmKdor+0IaR+hiJN+C/yBEAqdtO
3JoQ+djBx9uWrZYcpW3SnhFIoLzrcntR+xx7rIA++x4Id8uPWuIrVphgNaIZ3eiB/xAaszwdC9GU
W2K+pSee8ubQ1+310rj/Tgr49yPC7ht7OOZFVIHrSLcRm1kGH3OX11cZPoYNczu84PysG5PLckVj
+BvVHVoZKcOelkwR6DS6eHPaZk7ef9/WVCLaDI6M4cwrmM7D8U6tceBd0P2HL7t+0t5E9Ov8yvLj
zynFg3XZY6tgFLI6l00KMeUUSqANfyp/mItXqe9wsolZ8JuIKlM0MfLfANB4BCRoLZchYE+z87AB
iExRrNEq/lPBisI141XsOxyPn2utkvLg+btct/tiOMazEyt8NTYJjOd+j27ZAyGzUiwOglTp0eFQ
cwBp0hbZ2sow0mRA+3EsPXIH+XMmGmIJuJTHA8NCU00Q4ctUxMTzJ2osEEJ70njrJSZgrHRGfNM7
XwaWxgZLHnS/iAq2OOsZK5X289CX3F3Nm1RPzwDjaR9ZSRnPyTsHVWoGWTUMjyOQ5GGeORxp+qtU
NW8Szuj1v0EpXsTrKZwrPTpWe07TwESDVsAauvMC2WHyUt1dGAhseljAIkHJmlGiRmUCnu+ysEu1
+Mxb3KtenN27Evd9Ft9PslLPgMeUc1JY/heYJtlVyqfq6K3nmYsfAM4ziYYC9dMsKaDX8ywS4/Cj
Bq3pXuOiW0XFqIR1kSZalm9wjE7N3w5Ut+T+48MF5y24htW8d6zEKg+n96S991WHXgb2kARpPcgW
360HTRCNIBAOjJdBMhHvt//jhEQjsW6LsBBTVP7HZMcCPqlH1/xDOBECcbkGZ17KOZLg7ICtHx0O
poGxGCe44SVhu8zlr362izimNDNZvQuQHI9qsdEGJEccgvxQnTm1xDob4LCB3c7eQUsXycYou4r+
m+QnKXGZ576Kx5wWRvrf2qiaO4GapOm2zcKvkhbmzRi1PRhdJfqG2Jr3pnp3+twCJmQnyxYyGJRc
oANBd7AqlaC1bORDQFmhciyGm43BZ5q5EVdmbriEof94bbVxkHEOpJMaqh+ACJVWNxdZALHI5oHQ
KeXOmYG0Wb29Iqfr+ZBEzblPQ7sbsYTCLLibvldC9ST34rE17QAC/ZbzF5FqFB/reRyIFR9nj/Ta
eh+rhcJjbkWQOan9Q3bBCT4Nw21rWaM38oegHjgv3fm4DXjfg+m1lrY3ahOu8Qs/owSa3OwJjEBU
M4cK1aXbagD89HwiiDmGby/JPJKsOP1Gs74BCxqYGXiQxEuAOJ54TK+WKgn/tiMy6nu8JW1TNyO/
/gCbDxZ8WTeiQ+SWKK+wkDyV0SO8LdyFy3afqFskbuG9RYW8JEwHb1a8ok1ArsVeOrbhNyX9GoCZ
VmLjr+D2EFiz72SiEg4/b7wOOlQv8lZeBwGKCtZuq9XJ7ZnyqD3/nxqUzW3QLdxnXmxALB5K2m6l
Z9zThGphQyZBDgDsHW3rj6YsfaPUe7Cu+rvcK+DbumTpaXDGDmApOgBGGn4Y4zYgXVcWei+xWj/5
Piz8DvRD1jWWpFBd1k3DV/hGYrc+b569cvKL8o8w4cCgclTNzfPZEfzxmfWqFOxLLMrXpJt1Fkit
+in9e49XcCi3NNqDsfnxCOWRfUUaTgJAhes85rBxwksHOpEpyFWXmEzbVIEito+3qQ60lCaDLwq6
K1fcOpv0EHvRXvbB+3l9xOZ4Dxc7g9Y/N3qMZfPkHZK0KgGxL1SzA1Dv3CW1PnfyEbv6dOnSIfnj
OGc4aYDH2bjoV2c3PU7/1Vn+xS1XtxIbLlwrhMHj30I3A0OExW0Z22pi08e7oV5JfcGz2p8ajIQ9
8+llFznPsPqTPbgwG8F/liBKEWmn4Zs5s/ju/D3XCanyM73or0kpq/cR83dFXOrgTnrcJa2kzUSl
RJHIXxdljIRK+LUsOMLWEjQABDjp0p75ZuCt9ZrpQkBnRm6TySIjpmSkd2YoefV1eDqPHKmg9gmI
4AGTzoJIKj2kBQ3TQHt+t29EHYmocfKlSCbVoQsv0ofcrtDuJQ6NWoBHHD4OQTT0O3uLIvcgq/sh
alzRCLk0nD6XlVLIMNqcJ/hv+b8sS9kIVD0y5Qgyj6ColZeAO0MGZH3tnnMCUk/Es/WOn9Gfm8lf
famBJ5i/puOKrCriLhXCMyyGQC/D3Scc/Cf792s0gxsIJ+ugOeH7B48+er2acyq3dQkFC+kGANM6
7Ak3DHiGveOsMt49/ci3HIgwKAZpUAnQbCJwsVI1hx65X+fj5JNhh9EVTpI5dl+/R9tUuM7mk/ax
djK/Syeo3siaVyjUBqgbqN8GHPTJyX8gsn+CIVF0MV73019PatXxFlBOV4LK8xTfTqJwW+8ijanI
cU5deb+lnGeBeiT9WxYcKGys8/YWdo2QaOPkqnwyFKVTQTZFsm4ysT3uUNKH/OptpP6AlWmNT9aT
rxMJ10nx62EMItK6ieWNoXauQtMVcn4M7MPPCqBAu3FqEXRrtM7gZ7K6UDDrykdzYcLz/XFF4j7B
vF6bTsrDI916iI7yuxCXpQe7/gHK/Ik6Cd/Daitw8xmgEgoKGDLsDEEG6O+vAj8F91A7KkNZv4oj
tek5Mgvx/DUT2N6BkPkUUvtmqVHonybdEAVCptD8Od9QXHDDqt0qNLKtsj0xfMx6e7Gublje5eV9
SkaihQLNWAUq88IHlY3awGpJOt0ZBaghiFg698YUfVCUJYelacf+Pb50GGpgrJnTguPbkbjAGS+9
U8AYorwF0wJggusTcZr2TOf4jpIrQOdE5RvfmJfN+7HAtqwKftICvj91ArOdwEpyYmiwJZIZhk7w
ANXDlcGojpy2GIhi6uf5xkQc/aHg4Tu0sCOwNJRS2hOmwTqru78Jfi0+gQ/G7BmfYLsIXU6PmbtB
64l3mtIKQMnS50ozKDJqBvi/29TccHGV2SNegQnkzhmO703S5rng6MIagw94UXoyrryyGfzEXu3V
FqjeDYJQfTp5qOfI4BtzBx1wNhd8JrX3fO+9oPA6/Two2l3E28kgi5DsziZMpc3rBI0ROFNms2xl
fTRaPIWfbN/DHLxqs1kAxlrOXPwzLqVl9fIHL+IGComL1bvlZA4DYYks/nxGFsZwpYyeG82uzuI/
D+XwWD057SYZd4pByJ4eXqvZeUfFPQR6kSqQ6EyAXDT6BHKjZ50K4pj5v4qJNimTVD1/maGI7PIq
kbgECXBBQdllQodQ0lDFnRKFnMNeNUbMY4RExsdtCykfs1+wPUhoki9po6Wqd5ocYu1nIoPrRGd3
ERkv+qYLGjXlIvjVZ4SeYjlyJZrWuuCOKlaIz2+yTb0exxGGj8lKiBjHlP0+EcxKZHMdJtiSv2tV
itRypjqxNzl5JLsQI9PL8LyvvWGlQlOBi3mqrPS0axiCfjTB12tmKSwBisYtteSoKPmXI0PEUOjR
GSw/DArGABliZ33Lyw/u/JjeFezAehHNXo7gWkn16FkF/+iWpo4vDsfVZ9hxWfVpLJcFqOevzCZZ
C68eq24sCpC+l73HlQr1vRrC/HQCIecYRaX97s/TRXrxqhv/rL6Ladj6bDJpuNvN/gJ51wcWLXaw
RZM7auP3Vtmrw1vBSQkfm73Hzgi9YO2JhpBTsNLCL4P2yo2xNizftardLGz7qVq0Vr2qK96iHxDL
ol6EGvJyOIXwH5l+2pxSNw1+QdEMu/qe9DxIgszpVEPu6kgOQNsXasmwI0nxF5+om95ebZIOBLEz
0lvYQ3Z/mc9JErguMdsXhr2e2TsQ38Lx4zY7DKhwuemnIKXlLUXpUUz4LW1s/8WmpvrrdP33y3PS
nJVvpR52pHdeyZCZONZ27ct3akE/S0iyjhqOdYVwJP8iN7ywUCVQtndFx9Si8NVYvjickKlWmrXZ
xy745Mi23vtaD3m8njPPyLtcuhZnYqDxphhxjtO5foBhHmrrOrgm0FlO4SPjJxy/36+2tx3kD5Tc
stMUvH51wYmtimITXwd/b4NSOWwTPiuHal/ZZmPDgQeF2vQXk016fer1svH43WU14Hhwk//KLHQb
tQbLpjGHnOZtm4I6hHqlOTuxaS3tDYaNoBYmBmsM0NkrgdERb96Jo8yN8o29YP9j47ObZ4TQi06r
SCDq/On9ehXLVVlxoiSGZIaxctUTL77XMNYbUAk1TNUhC4a4jlCFd1gepID2DJ3mMHGW/OZab9ub
JGlzNZdKBqeXmGwUvvNGNDW5XSZZ4S1cyN2P11UniqEYkAS8KApMVXjZ8h+hNtjapOw8zDoCjSAe
TCKmjKgkTEVKmWcob9Yd2Qu3K7A5Yw79F3FHxaUXYT/K/GnYde/bqbHAHJsGLcxUno+TbspFOHqT
A0FnqZtsQ/qD9avdHmo4pC4tG7LmuzYJCZuNZLgLUAOMgEElQRxA6x/s8s2bPOKfbhxHKX3VbtGX
bSWfbBtiMRprioCj6HdBb2lQKbnSlXXpRp35OX7SPnFVbfsojRZU6rZQ5K1M9iGUv1sKMmvXjKKq
r2GmfJ8gVB0vHUIo0Zv5LelA1E7cKuVS9lvWo62QSK2J6ZCz48XwjGivdWRrEWCrmPEO24Ca8/8J
6ah3+pTJJ7zGFAKYMXHZZnPMxRDCA/gB7cqtjQIgCDbIurG5iC2MgMfFuYGsqGXWO9udBclp+8dm
0dUpPRfn0j+GDHYv77hW5Kag9Fx/aRA8xZGCEmIjhFlfhi1EOeVdyMkKcIZpY6wCicyFqdd7O+UG
tEsempGsYrO0fvvkeyEKfdufaYhNIEXaN2Yj7obaopn4om3S+NzboJYwvACq+YsTJesxBDIoZAOM
BrtIFRfxneExNq+lCWrK1OFyAbJx8QBwYTvnPtp3Z9w5Vnjp+REG0J8mPVa2JReQJAFmHHDoDZqz
prgEx4bOQ3vTHtHgeKTi6Rl0QqMTCwtH3wu1W3douDSTSxIMeexbfpqH8FY9wqu2UO4THcLCm9gv
5HRwdR2wq63nIZQ/gSGKT52LtPoik46oUJJL57+KYkjBk+ylJv2nSCFX3MEFaYedEzlzho1rPLLj
vOTwOMX1MMLyMCpg2x8/3bOgE8II2zGSEnER5UlBC/RAz2NacDYHVNYTJv5z4FCjRRsPJHKl32zQ
ASf1yu723Ag0zM8wbbXoJCEZp8P6uYrlDFbff9srMIxS6rTxuV1Y+WcdR2d/hYkBHtI0qqKhhhoJ
qFEOkDhqvnABXjL2znPAJbZ0fK7B9mCjTX9k2W43TxYZcEtZrXjT+gechVIW5iNci3zPTdfZLgkr
ifqIM53kWUA4IPnHV+quqBT6u6ji+8mI+eheopT0nRqfjxixb7xwp5mBZZKEa9KLu8focFb5Onbv
hX2O50I3ws3sYCwnfY8pGp+qRY6RQjcFV4pU7+OdebLVGVvP58iniPsnACN+1NjXhwbY3cQDOYnA
u+Ca8VNpPOyFkLbeCZy89HouFDn58nqW97dYv6o9ljhY8oN1E2v0kiwJsV+VLY3t1SYuVlqNp1Fv
9Pwf/dLeqKbRgHJ1t9TmySac3A6Gtk2k14zxlIUc6FNoK+Nd/OwIdlw7sNEjYDrb1204s0Jr0a/X
1htRpEugayJJczVxYgVlFHiTZWHWyfTHiPHH9EOGjnRemG60MfcOky1HaTOEqKORp1qMVw/9BrNe
4NOE3sJJ0e5tJJR3i8UqWhJoC2Lm4vJ9GIrL5z7S199NAJxfSTIJth+SEVZjpRXDU/8WfSvhtih3
0VzHnHrY+pMIoYNmgwzoRshKLSyd1PzUTIxFwEsVxGEZG/kZeC2Gq7l+AGeOzxH5O2ZTC1a3ZYbE
g7L0hvvL9MIFxHmPsrpX8loaUmELmA42WU2qf22KIcMGGjSzR3yVaOtKmbR3InqI/Ho4NeA2BUp9
jBJ4D2K/KFwjevtqZ5UDGttb9iKod2m4BFMrxIUeEouYBbS3bA5S0pI6CoXsGMXExy/3Y5Q+tsfS
I2Z5APZUq/86uLpfm/JG1/zL7xrup9s/M9nAWi76ydXgS1QcEHnt8cChAHAqdTY2aHxAXY0j+j4v
WgsGAACRqpA6M9/bx38/xgd56wUyogkvDCj3zVfb8wBryDv4E1Fw6r0+NmynrLXnW/LEvZx3/lR+
jlQOVEg9VuB026Lfrsx5ljZ2XOuZAYxzLnqsXVl1Gcm71/mzBiaH1ls1KsMwiejb6docFaCdVMrl
SByaLRQcyTu7xS7PTjVonBeP9ImCYqw3fIpsKPFOvoh8oqqgVdYcHppyTNXKg34lJ82An1Xe0taE
T6CRz0Hoq0bVgSbOh2RWHYIsLPXvJ3HTy2qZKCSq7Dyv9yJ+YGD/EEwk6qTUsQCoSu7vhi6xndXF
gqU6LW2zdtIzbQq6fzzgZaKU0eUKvJWCJYoKzrtyn7gZDefI1oq9s1UFxffv1ZPWChoIVniNXScO
yDQ0jRhLKbkYQBY91hVlH7VkyteRJ6gI7Moj/3oi7DCyPIhv7gewsFM1BpnVhbFQhR6lQd20g70J
03kkHYK5g0axSZ1szVIGpwPymPIzOfNqMTa4XjJBaM90VRRIlodk/Scbv1TOvEkQuEun+40uJfrO
Hvx8MjVG4ouvH5vJFK+Y86pTnP/xF5pywk16GEic/MB5SbJZV+nuGU9z1kc1lGA8H2Lj2tARJPFL
gkAU+4ViJQtxOo8Ets7tSSDYaGEZuBT0e8QX8O5zCLyns6tPEsOP68qo7GYpjR4Td9MVhpLnKbNr
lPEp29+4wDDcHm4blua6XyyHimAwfhXCB/NxAkrCI6GhxZLhbFVszn9myNS+tdLHE+JP3Bum3Ja8
bgX40EP/9pQ7hvXkhUmnbtnGkhfvWn+tDOZGmwtilYvDKQ0qRR5t+IP60A2NbutFrxd2gQeWu0Sg
lTk5l7Lp2VJrl4JjxyiKi300yXVHphzPk4te68djq9Pg07TkSK+icZVhH1DJI1VZ87vfMx6ax3kC
K7Tkk/hbf0287EmGtpoMyv5+DzoPv45aQHNu06tZ5zfSJye8HEV1K7ggQnvBzFvIOqspjZEnDTBt
jJFnvk00GiGhIKmsPxWS4wPNFGxstKDwp7dt1vCMTUJ4T+GmbPI39T3R54mOcA+8aDUEGWAGXnJs
ncfPisNrrpuz0RBZ7qEvr6F1/A5x8YXh8acIY79cosDVOlSUjKM/FVsFL6JokP9Tqj+9VFkhjKD7
mC4eiEw8crayIX4kbIT6yv5ZwvrYkhClaowfKXZfd0QjMnPfU1W4AuIO5+k1A/yikBOlXDlLDwWt
CIdW1ZIY5P+kgochNDI/A/9oHdtnNd+bipNFSm1vAPeZRsLKoaGHJG4mhKmG/cT3pEPhfwYMjIrP
VmSvRd44X2E0f7S/firnLlZTdxnFHdDuy4Y9xNYUj8MWP4uuIrx7WTbc7nW1tCgQg1nGOfSKeCMI
UuPr41sHbQfrkurWxRVIDO4X0swkYsx1iOCWvG+dXYA3XRBjperMmNM0jJxfILZJhnZm19ibER74
RHty2LNp5AVJ7Qc1b+WdNv7acKoieRtR7wxhdQMXFnAurBVSif+hdps5Ywxi6XX7gDFZZv2HJfMr
7/YT/tI5u+NHqO/7k0Kljleteee1pJlebKXyUrI3XCi+VJVtbFimEUl+eYzK+ZoZIMGP/hsOol0W
qjMLy2gvHafIV5+nKASHawKUZJB36+q37zMyxjkQBHLFX1ExVb/OdRJhVo9WaI2bwJ9a6YKg3E1Y
25V+90Uvltx0ZI6jzmEm2xZrROZUiEETY2tyPw+eG0M3CrIFFRZzI0B0vhFI+G6t+A1YJifYDug/
Hj8ZQ+FW+bBOfRkyO86fhxi1pRM08Wdm4nb8JOD38OyoV/zSJXNv+RDKzKwYZQFkoO6qa6zVu/O6
EN20lD3lnSruN2g8oGnR3xgrourlf+q/XwrRtfZ0opPY7yrek+dBDgiJ9PBCw9Ixek9PLtP1Kmxw
L+m0kFMujaf17hd6nXJpRIUAa7PJD/t+efDHHUqnHE8jMaEJ68JL3djVi3e9sIO3cf/rjuhdjqyg
itj0KAiV0g/B2JU8xNe2RWQBPRVdUTsARLRJpP0uNy09dTVNJCMlPqkZEjn71zBr+I8kLqGBI1gm
BBF1IaPF0vVPnoTxaSbSqyn1CM8YnHvy+iQ7Gx83HQWX+ajbzLfbHxkD5SqEknq1ql8MoOpo94Ti
FdRGvu9cA+bagv1Awdi5DwFnZm10Pkvy3oyzx2PHz8/tWUHWufJDjVeqJt0T/bJOu1bL/wljB7s4
MADW/ulioXVcuxvZJ8jVWBv3w+zOSb2FNr88iedstHDy1/BlMQqESSe3+ZRNcY8qg4jWxbjdAgt0
GWxp4+2jtJqwEkbxY/eMegaAnneqs3BW4V+5YtnadyZSOIpoDRLyXSgMTZyByr+Gh1upEsw1nhD6
42zEsoptiv7nCEEJGnXUfWEza3CcaiU883To5Sm0nA6WbLm6F0z/p8WWNuZOfdw+1mlp+94/KlYC
ygAEdikpvd+CoRk5cRk/973lWJ2trS8vlETrQAtSM+dCsT8c88l6lKqc93rDo7wdacaiiHGrsE7k
AlEQHrg2ZCWF4+Ku59UanJw9EeEmetrOvNnpbNtqjmYAEccZm4qNjM6597rEwPDjssbwa7Rz8+AM
s21LBUHGGtY4inZ7ScxuI7pDH6XESmAkmarzxg0uBhrYcYsBSlfgkxGugP7/FnlsKeAvKTan67/r
/7j1NHFtWRBy98twBR48wzwiR2Oa9HihcudJEdvqpS/2EOwKxwWL2dLUYDD+b7MkH4vtCBIvh3Su
8a7pVzF/Xaju2r+bVltZCAZAppXSr4n5X7ABseX8p8/gcy7cxA6wJhz4JBdHeOS4fMtzAUAhLEkb
Qjc/EdfQxa0BySpA3MQLjCImud+bAdV56byPsxs1klxHsc6Ma18it/XsIbBNaiUxen/u/OXYpYSZ
H2naiU1z+uC7ym4/OPFXS9ofP0D7tC3+x+3QlyxWnrc2DPqee8bZQAo+QAMWjfJPvIP7hs96lWhZ
81Yzpawi5atI62FtCGTlSwFFSi5ApX3d5NFpyPifqBwXT+MbQtd1P/CRn9Z3Nbdb4lxdPXwwqAZA
V8g5VlvVv54Fq6fNokbM2Ho7y2r0UdAPVbwrjsZhN9H9XNuIOw5aEyEFKLHBTWDb4a6rBwBPRSTr
HUDqFKwaqLrHXNEcYPYKM5S8PxPd6+coDCxka+FPHZOzkKG3qWvQVht5JMnuD99Lc6Hts+it5N98
8dlaK2U+6qi1siE2zwbYwABhS7r3ejmtnOrlN/JVQ1wXZoz8WRyqt3fyKC85Rp2qcLtxbOWpBPy7
HpnxRUo22IJdbk7agMvnvl32EVlEnqjady5k1gHnLPEWVCU9hvO/RYUyZBWqihdkn/sPyqRAW738
aTggYo5Ykm3mwJItmVyWePUh7gK3DFT9xLOht8JmAxBY5GT6/ARTivoh5Kn7LYzUDKdouKOBo24H
6itDdeRTjZ+PaaLy+lkDTbcxyf9T1SXKVfc6RAvr0mL0r+EmlYGBJ/p+gScAtgvurMlS9l7lfuD5
7XMxrjb4rZpLEpeIC889B9I1kiILlurO3LPJ1+nWR3XFje58NOD4ZjeRI+foQlwklp5B7x15Dek7
KGfDNAzzRdW0x1Ks313uuf2M6BSBynYrEZxmRbd7sIjC9zvO/CqOnUrZ/9yp1eyyOntkoLMYtBOJ
Q7uZbKrFyLv+gURtSniDsL28bMeol5LGkYZ6xKsOoLlJFLSiquKPK6PaygPI3rOok/mov2v/d2xW
f9ktBMWw/aK1jXfopUQ+VC7k8oDiViG0pdvJeKF+DnakEvMZE0mw0mwO/Xm63XAgAS2BFmKcF87v
14z+7D7iQIxjiV/Kw1sTEpJZ4/ckTdMFArCj192TyF9j6HMDiIXbcI4HHDmlNyEDXpIOG0P8bAOK
yNONxx2BzAVb8W0aX8ICRxUqCaPveZEmT6li79NVfY2kxM3OHRaI452CilX4QWjQBguby36/k4bf
uLYc5aZc3VsNwMRS0Ul60YAiPddZ03CYMOqbAG+OC16ruGHdImXmTurlYS6CNUCM8SEQHaBkf/cV
CkXxP1JjfYNv2nMPWBiOBL5BGBq1ixwY7hVlcs5C51OCksijkVCrN8e6cwq0y7EsLoyD3NjPs8n1
6r8dLI+izVMhNs5+UMTMW9lNvwmqsvQpAtB7e14NYzsn5pqeP7rbHyMaWID4MdzQJKcSqDLI+h4W
lRTD+IjdQtOH9kWNXNYBDC9win9RYww4cyu3cEeF9454VeIDoDJdWqD1wnr1Cw8yURkBBH5aC577
MMnQlh3QAwKbSK64uupmDh0hxHGjlFNO8vZGEPfSzOahmTi2qX9dfbJftZ8b0GZUFnmhAw6PUfQ6
cy0eclKds/xfWzcSiYSjnmqHYJmiUPHd/MF2CEVLO6I5Qmf4l78+sqlc0FtwC+t4gewxfU7XgEh+
BOaUUpgf/n1qfVGm8YDx8z5uF4IWb4aRoyU6zVxeDwCqT0B0RvopnLDu9V0V+Jgiy+SNyiwneRpG
8ratXf7Uald3XDw4ej0t7BruSmE1+oF3FsIx7zCv0ESuRBh0TbUwVXqUJ4qmWCBxR19aKSkUR5yU
dtl/zDUqMpTkpg+Ep7YI8MsP8kAaLT84ISHfFWCPrlJUrUdCYOlQruDhPFKc2xdTaX6sL7dnKe4M
z+oZghWn72afUT0EY4xsPFLZiJMOyTXbBgBdlVGjnsSRZ4kIeVz1D92wHFvD+yjx49hHRbtL5JFj
uVT5fc8XAVpswno6Z8TV9XYOPKGr53FfTnQUFM0/etoQbm0vlOd8QZmSDDoyuxMR3Pqa+U4JyKAQ
QBRPSgJ2M3vgV4Nzs5JzjlCgcd50sAt14ddQSiZtV7ssvTUNSbD3mLUii5ZQZ/AcPW2F3NLocDVp
ghDThCtqlOhUPtrESNw83+R5r449EtVskStkmgWNWuEvS2hQLgr1f8zpv2tttppmlW0hdIN+LmYR
CxWzEk5MjNc35do1G7OedaKpTuo+HnnO+ucglIvaNFRWZ8PNiBYngLfS/KzM6SvtGKghdt0xOHsC
S+qwmvtCJPS25UIYEmHDUC3+C2aWzaUoZ6lzQ6D0FSfD/rNy0vZE2kYf/pwlGS9Duo9ssMgFVFUT
INRxDc1jp+RxrTJxLFzKwI00uZkT3m8xcMn0BMlOWbPDBbcMBNOVtpT5IRaxf53DojwHHx6IP9IP
cAObaBFOim9W/7OWC1BhtOIZWGpCb+nKiBRHD+eNvKJMuJzi/IqhiwmyriLEpbwvG6yKGeb9jrEK
OzpeOpV07kAk8iGr+hBj+0v5EOIcS5RG1p35ApV1ov1/NyaBheEoRB5WDfkmwxbtH1C3sKTTX4Q+
3WvzGDFv981LcxMhkV3uKc9vyrb26w86JpObcoR5STlwCXjTKP+Ix/+oboA29zMlGRFko9nIYTGd
CVwsLrQ7HdCW7ttpVvv4eq0oGzDM90Kboqdw7QiYprueBKUf5VlBhX7Qf2rhUDYDpHgKEWwtoGrd
TMBv2ZcoMXLHneC+MFy9wbPTXm1PfP1kvjW7APYSrqr8GMlQ5G3uzSrTaPKcv8awMU+chWB8/91P
6zGxtfGTDWSb1keVrD0NFFQoipKM7eYpu3CA5Eo42ejsbc8QGcjpoU2Z52haf2iezWIQSX3OesRV
7XTkMm7lvXcM1Wv990Im+dH/IXjq5NyCLbUJtmCM3UDyEBeb4m05tND0owHSDn6jHWpgYe7jw0QE
MLQK7nzcFmuHasOBkbNwM4JOa1uBt3LdrYUUiizLAIOU5+1Chm47RuOC1lfP1ofKXcLZMg4Zk9VS
N3dsF0Ml3WfiRXhEtmU09i00i4H1fjhE4nZs6l4OoqAa46E9fQnyILh96gBBJ6dCn1udU1B/xbgR
44F4DPxAxzo02iOUxUkPU97CbH1Ih3n3lJlWJ67ftng+J+GPcm/z4Hhw2+icvtcfXlk6FNEvrrZu
nahgfe0RnT1VzHcefCcH6JzwfZ9GoQOXl83yrmlo7D0oMLspRp/ivlMCVErzQzeAn9okZX9SJlQv
WH17d3IZrBEiYZv3hRD+CdLmU9Dm3K2O3ecU6kEwgvg1yyhedFO2wPZI48L/LFLeD4cEDRaiKnTN
WYhRGc7V8owi4N4YQOTCuKe/b4C3iKubarWD5whE6GWtcKi48SSaJ2x72cMIsG+8hEglp+R55Kut
1BRRaEaKJy0BVKwTN5Uj/uFNqJrowJess/I2WKNEco2aDXVDGOaPoUrV4zuW+z1VaIlD58LmWTVc
uFLhQqw61j7/5HjtjQ7WYLEmU3vt6FuJnn58tCAsBLd5xwgvPcieDC9Z49bfbKFASRLg5lYkKLQJ
5DjzibQtEbkKx6HgRiXFQoX/3Ym2iDWWa5Uk0edzFiOrRQRnLHFOQXG7ClQyMML3CoRAyDkHoq6t
6Yxd8/6WYEkfgvtH4X/6DCpsHQ58RK+RO0Gab6F+weG1BZsYxvK62o6Gy5tf+TYcUwvNqzWLqBfE
+EZW59Bd86ziP4bUbCfQLovC7/jd9bHglC75h1sZFKPfrykDbwxXVgKm6wsPxAHmc3DB5PFttcOe
qxKY6TUO8Gfp6UmvqZIvHfkC/ym18XR34ufKLjHHv/Pcks+IBhrs5O/D9YaqCk+5jee0/YCJpIcc
vlzxF/Ep8/C+HFFdYBAHkjkxGhXiuxp8A4V5jGfHcbJrc40erP42H1HDCaVr83DlHIzcvt1fR11w
B6U6o2XL2Mze/5DlB6MUcaobGDlAd6QBYnOj7WDpM35vb9gBFJJuWMVLp351ClNjNqwhf2/bpm+u
frWplmmWiWZ/6BmEJG4gu07JoBclhbStM6JHqYr6ymmGlM9Mr4J25a0AnXdIOaiZNZXjI1FBEl1B
v3W7EQ6aaKIMe1+wSzuW+C6rb5pzy28J8fMyPPBWLoJdtfwQHPUNPf38PniRflJXeJIbuNaaerF6
mTTygTMA9/n84ENzqviFkQhY2clYyNWeoFLcIr+mVOsMx9gQJa2hqxYaXzaSFtiD6tdIAtvbB9GM
/ROixVCyFUFrpqQRYGsTkLkxPlS0SLMlyRPjGjgUZNcKdnw+fzV2+qwXXAIEnUsowiUZwlSMK7H7
rIVpM80Ncz6L+hh5G2XIuG7naSOQo1EFo87jwXlk0YkfTkzSHk6CaCs+h2bPKjhPgbRwnGB6x3hu
Uu/mkwDSuYBn8qxmyIZSNVdmp971elXIbCOFnOPGT66+cvT48SJhQPcaVz0dvruCz5U2U+2Hk1aY
zo/q7TJe16xTc6qN68+yofivsHmOeTf1cMbHKDO8eG01xI4620XJ7ONC7pdT4lusiOUp1gyhwos+
bSG7flZQjbeFLgOcA6WApeC3i7xO9KOJo9wcjDkUCPX+9aOd24gfTQPYvglZ9Gjq3QLGLC9D4F6k
k/+YPhg8gU/1hnzwN6ZEWE7hRQ5hzMDQmH58QDFWKzRGcjY6rr3MVtOsZzGxtpdwq+tEqQOzGiHE
PRmkGEnkhbSyQ+fscn4uDulpF+P9H+34gVxSiIpBawEr2kn6aQP3unqifURbGSDv8IYDXxXOtuGb
eUxPUGqh+dMHjv2g08PszM1B8/7FGtD/QRvKmmae4XNVelhzNysepGWRv1kFdv+Pka+lnkek8Il2
cSMkNisMUgt5OKvMhdYnYIomxFqBR/PtsMRHHBuJV6pIu3uG0tXnqgBllTAKs/OAzlb35OadLBYf
xKpTmLkdFtg1x1OX7eW8x2TfHHWNXH+i5EHcsXhnYY6Ffus5IuInEa5LF3wsIi2QNpJg0h14PjXZ
C7dEj7jf4PLaA5Thn54Gm8U+4vLxgDcVLnCXUbusgymHCjaEQMOVXPwIXUiCEVkFd6Fnb4lA2J6i
zXJTmgm6jlsP/ydm4tXKLXd6dCUWG4uE597dOJK/lB2NifZkJ+SoacKcBLSx+p3SSSg7z6Bi4SRu
409C6Yi+jSTLtjok8h36GFkm2sDPzFOrpAc0n/0vFigXTSLxxdhC4mnBdW77LpHhn6tqhQY5Lrjn
ZcCcLMOhwr82QYd5bxOjygxsnR/3w1RMfq0LLOkNDWNYudfEoPn02p8mWPi4aRANcEK1a36ZZE71
OAXvqoiMnXu1c2Jcl5KEXYHM1dJVidaDOqHKs9MNC/2rvNRTZP3cphIEdiVuhEGefuVdm4LJnp4v
ehZ3nPBlNymJ40xJoCVRcweNc5LF3ErmYZlMhrBSfO3mqkNLiDLR4W6cb8Qn2zIzVmDv7IOXiV5n
NUnUUp9jyVQyBJbkobH/k1FKQ3psQqWh55HsDw4xKyud5RAzlYvgeXE1bMm/ZlVjheadvGmq9lrD
DPjdPM33Yru6MU88+9jIv7SvruyBcD8z402Tphw+V5/5bNxF831c/V1P0bJUiDD5n6NBm/zFYmgr
K9EKxn/GnQD017zZZRgGHSftRY0CVCy/Y1lmhLVPmR3QOaNpmzeCSnyOBU8vmNuEb3e7kYMa18Xe
XFMQnFXfKWaUyM0nfcHQgdgszWX5KOJtJynF9jcvJ7YFRiNZt4hzezwOZNgZgr4C6JzyzxhxileC
PWjwi3fGlhXGe+svH5XCD3GVCpB5MtGYy3Rn1IRuNUZpc2lz5CNjeZORfk0vb/wVzIogJvSuuGxL
eanfYcyQ+1M9sNxfpRugEcqm76/fO0srRcb7cJ3pxW981KduMibfG0tQHFzmdn2Pi/sk4099k5DM
U0I3HvKY/WiO+ek7d2CBYed7i10eBE9kdwZOvEaatZIIFPojD6AE/93ran605uGJPjT+p+eXEWlm
b7iR9Nl6v+n1xmzIlcTC35ksSsQYt1LJ8SrHy/Tak4eYfBWBwAAzOjRef/uw5mz1926hjzCZuHPB
0j9eGfH2LkoZUQRverN1/E9U0ihD64s4yvPPh3iZyhD66TAEk2RXRICpVrvgp2L/UGGZHzT8d3SG
aWhHm+1uxEPTugmlDAo11eKJdSfBrSQhMNDVn8AN7mLM7ppdoNsR3TfBL+cxt2UbLxRa/L5nP2P+
oQNe9ta48P4dgxDxHroyE3pzn+LvRnYdsCZFfA5QB5e1hXdOAIZfwvbxvfndgS2W4qoxMbjHjRnJ
SMuPMWRVJSo46HN2j6/t9FFw509i4umUeN8gaz8klRzB9j3EDmiU3SWGuVgkDKqyQjCVdzYaaAjM
jmcNL4n9X4x9kDy0J+dDoVkG4sw8VgP6oNNM6Mgl4TCL7+UR2+vLkkftBV8bvyGueWpTsSYdBZTt
jutcba92Drm8rlIMnAP20ZHc3+xHv4xnU6Qn/dabnibKluVIyecFF7gKywtlJOof7Y1XCgW5hZCs
Ho9XJ40HrMRDv/WoBkrZFohqrJvsZ4VZrc+EVbQxt7MWkJoJ2N2f3bax8Z8v6iuhZXxascexkQl/
6BtyT3cAiRq7aDYaWjrV+wn582ckNdn7lxS72da2a1VRW+eTo+S92ZgBZ8GoV+z9RhScJeA5tHt5
CF7Hw8ylwSHger2qWs9XxA2eMGIy9jedJo8VYR3y8VHaUNhM+M06VEgDPLKjDVUhs/bnUWkC9idA
awCwEmz8b+z1nslYasGjFZkl8nf6h5pNWBzKuCIvVLSfLWkvlwslE5YEJsMwszdNTQ+PA0AYUEPa
+vdUZEHQd4ducUIV9QZHJMUtl25P5MNbMaNbIKInV0mfQsoJ7DvkUj/lirEL9Y0HBq/ySwYozCcO
t6DANltKSCyM4oST/4Fmz8QfaI5ISwmk/yu7iXPrRLvNTwygljhNcjTL4Cq/iYv2cjI3pcGP/1uB
2FH8WUxcehHpjoQMlLZ5HrGaSN0fa4ttZAiAURuF6/ltT42nEiYRcqDe556oYSKIwwbHusrq4J5A
dMQKbJz1rYr70Qfw4d/Gf82ubuJtbvU1thnTR7+256HCzi3w+wF0u+sTrBM9SP3GCnKozcAmE4Fj
5fZx4qLyPMJlWQD1RiXlNkHJhyvll5epQRC5RDUEe05ilSuZG+P8adtTOlwnG2j8QjIe9xGqG6AD
aRJwjl5G0SjAClAy6LoADR8oXXrcQ7UUWGIrldHvP10ggX8bh73koG4U5Fb0gpWWxKwsrsefnZoJ
+h6bZBp7uZFbrzQGgiJkDGdT95LVBwAluC4uyyEJm4tuCKewq4Ry4HbHwIe8wPFOqwOHmK7Z39HP
sR1BZJKZ3BsCvulablOBZwyl+Xjcd5tNjCbPTk/PL3Eg44Nca8aFcMWTSnjGptd4orlUhJvMIqKl
zkoZpB52gU7FeVQrhnEZHnIurYekhyeq59TSrlH8hxo8OcjI6lcqvBWvDaBqPiJGRxAtIeQwUrPh
958YrP4LMTI/7z2M226kfU9KNL98jcy/Bbe5ImEu2L7Dj5pIt6hOFNJqfnZV4lR7rmGntEcyh9Fx
FZqv1Mhir+lBaarojBLvp0hVe45C2/Ax64P6IHe62AD+qTYT2kJRw/0j1aY5bbW2Tq5X2hMROmf0
0ob4oLBjjq2MSsgz5fitAi7NrrYtKs8NKct/V3mS8hCSGUeD/at75GwFDeEPjBXjh61nY9FtA0v+
fZjv25CjHmY4NmQ2o9ITYH8Pwxgc1wrRqo9bqAfuTlzJ8z+Ysd4TTn2j+DOvWggJcHA58L2rNcwy
p98xhW6ZkU+PmDEQUE/gUeaojdDdIawZlzVeZr76qi2zhSKtLrW3wQVjJcR6YIDZgKUt4qzkTT95
M3/JNKEVUnybEP+/0yVYf4xoNtXR2ngOttz3fBrZrH2ehgqb30BBkpjpKukCsM5Eyp8yqDBMSfVY
hRzvUijdg8AEp2vimyNPgDjvwyi8bl38eIDMWE6A3vsXm7UcrFILI4n/G3LoQn6NAVNndV0hb2Q5
kE1dRjC7pOFwAUQO1rn8VSqp45LUzPRM1vVRrwYkeSp/KMlqVM9PUnHd1a3rJ/BZV39AyvVRjQha
FrzqAuBaxA/c51oLNVTwaaUxBnWxjv1+qNVxM7ISkB4z0MqLrIV56euKSV/YhdlKVJiHFddzeZzn
yvU7l7McdNTHIYuuNBJ1l7yTBouLaoA3HgnPSUCipfDMmJrfO5b0E+DHxyzPpbFq7AQkDgRgYOXm
HjRQ48VNUwiEp6MN4vKCBot96X8qZlXWoUsqvOC3FKxwTkYFweJ5rkGFoWPK6dVIm8T6AIijaQCj
Z3gKE1yhosIbarpFfeTiquGjB03+gXaWOlk5FnInFmQLZt7/J2nMVlXxJj3r3f4EthMvOIC5xAKv
SqJnmwi1e6T6X6S8hSgLen3/7135hxbNp2UFpHd7XlSfxDdEnBWYhmXXJGTekXgxDjT1b3i4PYLe
q4TSuFVnFIIdjuscLmwOikVh5ucH86HD8jacpMq/aq7nKtbziXbecpl6h3XU49HN2cecFBzYRs40
S9QOHBWlfpkYeDNa6sMvfnuxhYOporfiQUV3YfqI6EVzhjN3OwQx7fPbXViwTgRmoIymwlDO6vQR
bwQCwkdd2NjZFJ9R8smCwl0hHbJFiZvI7sVvOtcbCXvCLZbg9OfmaZ8JSyJcNNxbhvScsiJlhMMz
rB6OteVUJq7fvrZYY4gcxAiAysb/7Iue+n8Tq6pPcULODzaxxK6mC+lbL8kOzIGVWObSvB+7MsqH
39fMfmP5hMa2EDZkwjU/Rxy2F7oqS9mJlNGhf9Zhxjak9gABKO3Fqlp6akJd2uDWG5YW1eVj21ZS
dubcqR0SsL961Yzryb8eiVPkn5a4jjIGDeG6xoGoF9TZkZgzK9tfx4edXox/rrXI1eTafAU2xKeR
kMqwjGGfPqdwT1WJ2p6gDjW/Gx34+jRaaP9B/0mcndhnkDXvIZgwU1v3fasy0ZocIQVNe9pFTKdd
tsc4jZyhNWS8Cy0bPuleVgvXXzmwHrB5GhPjQ3NI0+SPv1xS0BQjCQkaID5vsNwEVA251OBg/PdQ
fB/I1DTqqWBZK2wOpsCTDLX6ZoPFmoFYsnuc64KgNRXb/NtrTFAFSJ3fYBX6YGKnvzE4rRm/MLaz
tv2ep+xVDyXnqIKh5+9B+6/eWYKTknztcvLT/lciZyo/kJ8EdFQaNl3tOYYjTCxGKJVeNB6B9rVQ
+64HqRaMQu8PIzB1clZ3CFasXmLoOfNCxImkskfHRVd5ohA+D7FCpfVdNboVi4UrmRnlOGNSXys5
hGMVxsEt6sqDoiQCNZAEli+Ts4Hg5LULvzWy3bRWTBFOh8C64YLhb6TiZro6eMC2W8jQ0AAPodX7
JDTFrJvWk5O32x2XANrAbSHsOBPtrp/D3vUpUp55Nseta0o8zBHwmHSA7ZDUTec0iXqhIqiMoozs
RBbB4znFOK1hyc62Lkg241EgAt9so8x4hp6awdIB9UxzcHC86rajLCK9VcAsjyAASGvgyPfBdh/L
CSlQylEgWXv9cH2FYzFxVVM83iAsgJ6lKc8e3/LvmLSrgTAzwsBzI+2zzibhNNvpG6uyL8iydcL4
JVIHkA07iRRseKSwQjo+7HnwBvF3WhmZJuIBla1D6V+feCHtg/Q4OzLJvhFpxa59JueAnMBckOzQ
mDgf0UD1L7dZQEdvqVmdRv+C3EaamJFtLqFbSXeUHbBWjaNs/8uUb5YxSopg25gUwxHWHmyiAWTf
pea29vMbLdQPnHyTCB+cK7Ts3YxVptLNXpGvvJoysmQu6WHhKpjck9iTBzOJlmcsNrwhM0NgYkl0
3a8cYTwFEDwAGiyz7VfFQVSQ2ikYvazKqXDMjTMncMxbR/75wFFMD2CmzLI4Qwr+VNzoihEc2Ddi
9ZMVuvFqksaNrGxUb1G1sOrQMhZyooCutuEG03CcH8eqrHI9bYyTjZVHgAb8HxFMBxEDEuElZcXj
ZioLrqySdTTz7DPj1X9+sEWBZEM4lyb9+SG2VOVXNwMMpI1qsHx85OTXMH/FQ/c9NXjNiXMnEYd1
FYRcFRSH0HjLtxLn6Tb59YghKd8BdpdnGR6Cc2AhDRBUbOcdTmNAyXb5ga1nS1iMbjbME7O414a+
363JuN20K6qCyLbT0iQABlwe64xe0MYRp0sleeBELKe5bhs55phRMIU2UEUiA3Zs3N6Wt3zgcYCE
H9T+y9ssoc5L3pjikzBTAK2ObAxYsOGnhQLiUUlYdHA706DzNeECsmqmyulo4sokC7H/vnc8LdXu
lwJVYfPl23hS/JFbwUvGejRjepwO0gUch/8Vs8FybPkfAxc8ENlwyJ5jcjQkCGb/Gd3fcSjIEULS
xhYcEcx3WTSLfZvLutDWvzkhhNAWQmU+W9LXGt/Har1e7q4Tqge0NnpxJCM13+w1Rc1NDBsf5LMy
vwy5y9AZopsRg8XT78oNcGGWOjZTIf8PDZmwYqoTYzWNAl/GRkXlbZp2etd00669q3F9OUQrkRMZ
7h3bj+tZheD3TvY9ArDdGRgiiuSbWSP1OlgGtZ6GuRLHxNS0efIiYTPlEeVCMHZETepkNLVJQOwk
Q7//UCZcbPU8yA4sR7cwFaJdXIa12/nBc5p70ZUxBcT3td/2ofwygD2z53xrP3jzljqJ2gAw8Fht
14qtX8bCZE05mICELALZcPnVxpBOgQd2iTC6CnKh+Pf48AQf6QntVMlGtLLBE4vFB8KbKyW2sFBb
9xtoGm3UzNo0d45bFCy3TzWXWbkvYpLY+q3nRTQoULICDZGD7LSlztzuaUH7b6X9nWUJXKlwM4l8
4iwSddtrWJ2qHmyul0o3Qt9FPzXa6YpcM7L5w65aJDYI1xcupC0gss3nJvz/YcDeOYLiFp99125W
TX6V5i+bviS6ek9CPsUQ/RRMAGnN3SFNkdZOEviGMpG+Ww7pe/UfPVdE+lPKHrbPOqZbyilnqlbm
bNvCMqUZhN/567wvIKrwJp1By2DnqeGvpN6d3W3o+XwjRhgZTds/kccy1Je9QKKxSGQuJMbW/0WN
8pCREotn8iw4n/upcfzpY7t3L1xDozQN0CIn+dNFniQ91hzzTgyk4Bxo5YTLJA/IeB/LFERlKfrm
fHo+bhvNdJt4276Q3A4R0tGZ3/D5qnv6REgInDxNGDxdQLCWn5C6JRJ4En9uXCc7SFdqK6zWwojV
kUNmQzxIMzGYYAQnhkjs3Pe3s+BQ5Z3gl/4ZzkUnCpvJ594EpVo7JbbimUTDGfVR5axLr0HkrKA2
4lIrdIkeFPFTkZdTdafiXsToFZZinGFsQ1gLmiG+/7DVsCTD4Ug3VjOy2S04l5VLlpiFeRAUvfe7
NXhe4Y4SnNWL1UBhDaPDVbrOIJ2I2CvoZmZbf41nojljPL/u2xhUoz0UOnKI/w6+1QQSEbFYGFQK
FLWr+6Cz+0mU+likTUIsk+NIBm6SwkHume9fLG51VWVaumfAs8Ndr+9Zo/nd5kluxKBRuANPpP+e
C3m1+ctAGQPrhj9Qgw8Rba+1IO41LxXIabck80X6yXE8e+Zz+j6jzGLu41vJNDCUl4N52rNn0gBW
lhiVZtVCnVPjhk9mxn2nu0ESbxYdwVy5OUVois7tqxBhXHKDhbKpmj+YWYxwOEvk3yCt73hJG4c8
4nqw2P50P98gCAt7Vzs7pZQM9qjIanVxj4UvB8IJakOSDovTNhC0XYCcKLBf3OgyTaCr5IpY6yvH
v05wGub3brd9gjGE4RzBjTETee/6qh4RbEySeo0RzWIzKKoCxPZ/iuvtEDDZ49Dj3IzlhTlLYJDI
a6VrbwZkBKl37kpF0hDt8CkiPqRqwhy3dtgL+5+KYJAiYox75sIvwdolfdEikYjHWSHb21QtgJlb
vimpJLinSXLopB0Bzc5JYS1Hew9LPXf+Xxrf1xvrFoSaiy/HzdRIpishY3SgtokHqOzR4zHykteu
apYf7HAlX6pjGDaqvIUaEE2fiSJiB6PoNozDFW1zkKrRb878oY+msdJ9AQXuvaByoXHDYxKu6FqD
4VeOTroeUYF1eEh77eOjqS1JmupYNF4r6ZSUM13RXp339Fgo4GtVW7WeqQN6ZD+oeNYsELZZ/Mqv
EHPFpQ8UnmrzvG4plraA0upNuV4JwFS/qbYD27/DNhuWQE+J4AEph9UL1l3trdGdLXEU3YUFjE3g
r3DQ1nUPRW886M3pq+//Z1+gJb6KaUSZZ5oHPiXgKbjxlIPcEK5+l0VfmSC/ouhAIlIiEAQKvYtx
R7d2Yx3qBlpZ6F4xS4Ja5cIAKNGrPYh4VTwkaSyICFVDa0XcoYfueh8Et2tIa1NA4IU4ogf5Oyzn
ctoLx2JjSIIXoXDGT3vFC/xLX5sakxd8bT+VEX35o07spyCa0OOakykWTyscQPNxc6BfkC1rECln
o6jNjdx7+GMSCjkQmt1MT10MFnBqXwmQSzGM9T+ylBGBS4l0aMzXhJyK5UGP8W7ZlsenVW7n7eWL
6KJUfX7hFYqI7vr1yHApsIqMgNfE88yy5kxfKwRcNqS/S3Ag3MPJG7fpiyzU5khzL1x9zp2sfSMf
Sj/bbOzrizJIPQHJZ6lxLBhJ2GCVeFyNW1JPYsPCJ/rEUuGafFgZBOR+ojPbnbnCOqKHz+oqfFvo
bMYYT+RCSNLqbQfl+1Zpau5EiLx3JCBDp8ryPt8ABquoA+pxVAqCUsjvDSiKbitffgrlmVEp1qRu
MxxsUF8iuKXgrq2TKnisRMS0AX3g1dLuli4o8btFWpqpSSp7AAbcbcZ6eS+H5VWcAa4dPSgl7Ksy
EbijapoA7pQBY70kmLgD8pjv0pfMllPLC3YH+D5rGZYJZ8lJ23O4RAfqD1J2vwTDOV1o7nUeKhlW
gqMVKW2aGCbEWgFAAGCs4e1tYUiXVQ57yVlm+H7CEIxkItNwakq9kyuC0IWN3ydpvyGyh0UoHLjB
G2kgyKwgYiSkkXhwBK+a2OIPmRSnK8NeZ+VOR9mpe0Ws+2xMyaZQh04Z3KBuo0+T6uMwb+AAMASe
OcbSaKhoCeoEs/yXGaTLYXZJdI4JUme2BpyQgPS9POVdQZEgc97A1kEzBIyvVkb6hdMyMFUY5VR9
T5d5iQT/j/ouhJSuwkgifyGC31dkgpcHtDeQu0RVQx2u/1qH0KCi+9A+V1PWij6NT2Tv8uyXpkYx
0Y27of6CqNIfRklnW5xi5H+EcOq5/EP3OMdPF8vAAB6k1JrQU8nhYHulRZ15bMejrublWuKuOKWF
ZrfhoXEse/yn1XutwSeYLGdrWIhuL2k9uczbFxEsLthndBFQyA3WVSneOUeyBFMu9H8rjFzF1H9i
FI+gLjtiwVyGbjXIHQeyf6oqCDJZ3P/3UlDkdc8mb/3eNElf8iCh38TGFA5KwYsM4CzNDYxGSPzZ
8/ropsut9aQFo/FzkY3Jw88aWciOkS0hHSO1p4W6Qe9t0jTBE1R9N4hs1ttD/LZ3NZxMAunDT0fE
Slood0i/MtGqeGMO9A5qzlyt+WEnyVZMO2sKbCxc4EtOJvgKRu3dM+G0nIzxx8OqJa2XuH7CAUMJ
to/ALek9kdj2nuXU4IqQIRXFmUTkWCKd07EAQR/E4oYoozqn1oWs73xMvU4HJyPvocn8pcRDA2qK
I5MWlUwqgd4P/ZeidRzzM5wU4Ez12BCd6hV9bVhmT5MFMJgwhDblBbna1qThveJSAnu4PYyHY6K4
a2Aw5MbIRRWaYdoVCiivwr6tFrJw2CW9lXM9pYEwHN848r/hHhuzbjpQx035feITZBwQ/84j6L8k
gytq58f6Iq5sa2M0LfAF53+Tg4rBf8PIJ/a680fr+NqZaracBgdLZe8JzcydgSyKuElvDZCyUJeq
3FQMjEp7wv8uPNzKxz0395BMoZ7oAnlKnW/PvL2nv53fdRT+HEg2gOdKmdm/QNJlQXLMmgEOBWbZ
B5lkNMBLDyaGMoXam/fx+nEsXk67ggdY0nMmefeAwWZNsfH06xpG+EF8D7FUIelwSVj6Xcwy+eAb
HtuAwC+Cktom46QO8oEuyZ1owYw4wZjo1iQ4plDsHoPEjyzrtuLPSpSSTJX/0GOU6bK47/aAdCki
/6yZEhyVuC+rioes6vMiz2PvYnmC+f7qiwbRfW3BOtpxduGzy6mmaAKR0PJ3KKn9Op9CgloqEJMh
6qdrwfzn/sY4MmrCo47X6aQfcnfvO5zuGaCOSRsgnWTD4rbwAvlk6v8W5GBtTayR+F1NCMa98AfS
D74rk32J0iK9uDGflFDgfTSofyBI2GlbGoioE/BbGfCwe0alVf4gPyWiTbfsKZYjZo5/sHaKIV6U
q3IphTfw4jPuUcsp8NpZvnUaYbLgKK6fo3bV990mgOJo0vDde5S2+ZplgLPAumP2jVzDd1a0qD0f
9HqCppkhTL4HRnUY0H24EYbld/WbpwtdZjiCVQ9q2vJZSWxOxwpSp6zCFxPylxsnAmkDTRCgS7zd
bZbg+gkow0YzqwMw8vtJTNz15xH4eQaSKil5IKZXBHbkbr0lhuw2bzdwknyDrsrZo0OPv8eS3F5O
ci4s/8jyU0ddfa8/kPkOOhQQGimPZbF4L3qlCGGETMrknY200OGQvid/DQIYfIVV18r0G1LjQhau
BMe2aEqUU+diEdUYfPIRdGENASNNdovjhSNjgwJJ4xCdBnu55m5GEDsHs3z256EPh7mdGUTghv+/
Cwg+RvCbxsj873TwqSBLSgZNodCTzghbUx8LHxNf+B1e51/ZP/Xqpj+pPkWR91UNgPE8Ws0A4e5T
RYwKir6lmc5Ug7ZhHwjKknfoAigNW1LUXULXM2KsIKTT4l142wmlFtnERo5zmlpjcunyan+tuLOf
HNWTDfrVue4LY+FRGeXA+KXSmOLLOauyWzNoFueTPjc/yOUaUyvEKQW4lZS5CY9gyv8OyMw7q7Rr
KHGpqYaWHg5wexQgEtFnfUHD3Jyl3Y7bNsumEpkDkPBNfiYDUawlk8d2QW/+2kGtqtSR6k8aO+Sa
khYBtEQ9yBmJW9Vz++4b3ENLqK26tZbQA9sKj9xs+THZko5dzj5n3MZ4vTzr+7odM+B8KUTkUAAw
mhvYFyjswWaB39PX21xRYUymWdwTw1V5pbR5ZPek3Yz5Y3PE+85vvpgFsVW4i7/jY+SgqSD8IuWo
zqxFaYEPrgctfcqd6lIyhx10yv6b2G4uP/LlG9qKIwd7jnuJfMA70tXpijXBBn9isZT9DtaRecd0
z/X7omx12lV2RjpilohpMSPU/H224vC9BHxApccDiaeAWbBJX81CDbf4YvdIaVm/hQxDxSYAy8q6
PIi/UaLw7JQXDA3sGDn8CCAxRQg8/XbgUcqrDv5MWBfsIaB2KJuBPbLuh2hWwIBEl9WFMelXJiRY
VQ6/4ngNCrxn9L1cX8yvhV6rKuXgjAzFwFwhjU03lqLaB7WLXhVtU/FONMYlC86GV48ek+pwlJHU
P3PXcgumpFKgw6DllIqvrAocu2o8ukDIxZlFIAMNTm3uoHVVSDpTddWRGNDm9WvDHXEbXbB/55qg
ExO75Dp+hJf67rYyEMk8m87hbBe0xD3Hw8Jz0AlGLU1qSvLFPY/nF+A4V6XB7Uld/KNUEFsFVGXc
NBvfBPECaDtMEhU2pxzKFRgQLxNNmPTuKRvWpQTa9uCzneES+IqdSdf/Xn+EiTM/5rEGi2ESvtPr
YiclDpEM8BHaNxBmV0AArOb+Zq1sVgKkqkMunz/bDSjzaI0nVGGlWSNpyGi0hRguTMvyP1IQS3QX
8O0uej5wL7DYT7MRRxdPQZUBrRnEZsOv7mjsXyeKg7ruyJdh74QcRMjOuGFIGpfoTPZdFcp9eljj
8/2wX/21vLB64RKLPQQ0xeXz1gqsVi8rCby77rH+QsbjnWDsNPoXna8ymVjrCrayKf/c+UMAGtA0
LbG4fKXo7gj7IsmNRop9ErhFvGDgsjlxSWFzEIvd12BNGOJdwXa3HxHPKtEvOezxTZ6gz/R64bGv
D/8hcqnmofb1cfq6tu5jj8L0dNJCX32tE/XPXPW7nmPRGjM/zx36kiBq0T1JJynjcZx1ikILsUFh
utbKVT1H99aWOHnbOf00VTYIL0BvWYe+GAYZRq9+6qij9G4jKqvNAxzzUTMR5vCCvi+j5UuLhSvJ
+SOHyZ7OnVdLaORlNXJHIclCcyfnPTncz/z3MalANh2p03LbxtfdLvC099NBvTgeN1bEvELhbjGR
bWzEGpz25qRy3xO15BozZFGZ1V/SZNmJds1JOjVZfij6cQi66I/h6IoehxOyA9417NSnp0+EieZE
jNSjMSsgI7UrtH0WJMf1OE4xvcoyXdPdy997taUzns5rkQf32bumgJbR+hzo4SLCjawi5Px4szsf
XSeF1+qYAarWyMkApH9qdBp26Ae/mE7rw6HAx9I/2xwu1hGMXuGVAsmhbhxNpNLb3um/Gia4JkO6
dKgq9M6HTiBN7OFKpHSeAaFezujSNwqz4NUygt8S1tbfU52/ulsO2QvsPb5B2IM6j2Px7lfmLK+J
t9Yy2ymNy2tOGwAd4HcdqyXCrXIT2ZoXo3YwguYr4LWHYBR8eDN22nCFV+lmZUfvBL1MY7cJvzG/
BgwNAsl1MxACSj3iVN+WP9bHMYjRRKcz6z2ZRc/vN+2laQMz3Yg9iUVFziA+O/O1sr+QbBSOM/XB
R0mACTylXWlndicYNNLbbavpJVhchsJ7gpoCcICt4O1RCX83IyLUMXIxRHI+jFtEHxffpINefj9l
hBrWTobfR0VW0kl7Ab523hTuyoTz2FZ9t10RC7JmMfEIxeg7XCWW3EHyFt5zDQ6hTEdhsXcrD0YU
eX4M8cNb/sbqHfqI5uNxzR0RRZqxQakWntwgk6U+qbN0M2dgTKOtvPeh4U3p0RPI62Hz1n0QtWqm
KI5hmipQRZIxrfe44YeRcvZlwwriqV8Y6kqscGOGubdCntVj2S9eAC+3bDefP40nt7oF1IrETDb9
TFBsOC4MZq9OJjHhm68uR9HEj5cQ38ag2/4+B4VBAhJ4U4ACHG2yElLcT83to7TsPks1y6iltI9l
/WkFNRhcoOQns4FBMZSNV0qQb+UTn3n4m7WD9p52UEOaPFVdcIDNEqRfnKNDX/hTs8xvtfhtUPM5
btvAD7M6uOlWvlql32oH/ANDKzbuUjnz8x0HIGRRNvhCM3hLJKGVVEUPpnHBe+f1bR6RVW9KVElM
eatfj9IkQr0ysEj0LrV6eM5X4tESia359fKo2/sSl2gaF2VJskXVsqLI7osqpBJeBdS3tCgqsu9N
JZ3BinGPc5CUN9Gon6pJHeIpUxaB9zuHrXqcT2YJyxdDX8I1fppjRXo5+x6W//tFA/mVVnEvoh7r
sU63o66A0uOC0Ang679CVwrb97FH2Dk3f7bKKh0kdkzqflPqGlizciiY+4zJOpsEa63rxdpBTKTC
+1ZqeWc5cpvZMBBXdedkSLFzDAjBcYO3w13RE13M7AfKUu2dWwW/3Gapdw6vUvcsEsxymHTC9Bec
InyudEkYGFYwUj7byehL1ptxMsmnK/ml0+b5DIT8IGBsBjuw7rSDvRYW9igLhA9m7YrzoQIxVB0f
3QMeeQhJDqtjX0vF386wHnlf+S0rjGO/SBIvjizYZwnTQjgnSpBOX5Cc5xhnzwYOBi76fMx/P5BC
cgYrCE4GVyzIKqCGQR94Wxw8/6NdRvbqpROm/FuUuF1DNRQdDtBHYQDQzl/rqKUKV/W3e0vuS1R9
pa1dwAWAotWY+DazTtYbVZu9IejpQaeDU0iVSVCrBtrO0E0JEsXnV8xRtfXph6Ux0YqWIz3B+VZE
dT+m4VectwKoUydpxG4qsIyKP7rxcLYbjhQQe4bOtXotiXowSGTV+70pDPSD2XphCAwNrsge34Ox
MRzlHhGgCazp8fPapj2q3vHyiQnw+xZJb4DbeQ5UTL6LT+fv90PWV7WJ2GS/3UclVcQPXH4j6RXL
jsD2z9OAh/9wprH+0vgyPKpV2YPNiT2NguBAcg3k2gBnCjqyMCTkGZYgSNhdCXisH82eZfgWpqFg
sFX9Lrye9yQcGS7IzyyLefq8qZsbYqowb0tVcisy2R/yTSMotfJy/B22aY3PFMpII/9UF2dOvug5
vKh1Ahl8US5pTLe/3pcE+W8sO9WNpDa+YOO3mMc0z1bvpW7RQciYql2yGk3PgqueraE104/fpD6J
4RTf3yp7ZQX/4bsWEWFSk8u2/9F/MSeRWNbM2WflYm0YyAN6nZv7lSy/S5g145KVn2Awj9lW2tMG
5XBjKhoXBt6jQgipfaKhH3lvWqU8nhOqn/1VIldX2lAhapLNF9EJDMmMaxdLhiJ7ZebzgXV099Li
i4gKCyp8aQZAuM2WGq7pPUME0tEjlrF7GZ3IrKO1tJkD9NbpM9ndDy3xbMJNTqqqNSSXMmP+CL8U
rvwIpw7SrhkelGZxLbvr4mQZJHdM/wGQ3iEyaZpwvvCNaUh9uFdOBKmr20fuYsarjXPxBogqy9ng
tW1xnjotyZQjM0z6tkgdNDmGPy2btvCihVk40ND9L/vN/kyUIZ247+cFs4oRCxf+AlwTYdrYk/WG
h4jQ89JAeUIT1ed9Omlrcze9jVWV3beM9s/nkj10NOoSYKt9VqinncWW0eRoOQge4RzJbrHosr9Q
NahhUriEBfESIyJYcEWXrlus8uxa/yOHgw8pzxPO+/uHeha6nyWjYHnHAj4gOgA65sPAbDeMgrbv
U5Ea6mBYCGa8e+vQCFTXphmLECzl1a3y438QgDVqXSGSv85GMfCdSMQF1SU0uTgXdjsLDnxBpv/t
CPO4rWYxhIR4X+lkO9Mu1UD64UYnz7zx0zq5vxjDbQh1UqIqkDoRC0oD6N58QPhXjbSUA57zfufe
grZYwP7kBsodbmlYmsBV1E2GtRDu4/3/2miCdPIZxHfHIGlthUlHlC88CJWQ9Zc+XpkS37D2/NWp
wQ+dOBgZMiy1nhyMFVgl832DmCXU9p7LkKPoabADnlM33Z4Yh5WSC0tx1ZvUQTS9+aKwH0+M/k9Q
nrrqqz8eR3964BUs4d+IIQP7hqqGGVQKtIs2ITF8wMf5kwPdGWxxtL3sNCh6R8YCCuy0II4hd39h
LYIjHf5vPXTko6yeBMoKQK1tJJxthCpO8qHZIfTOhAVWt0e1/+dYCi2WXXdxcMRQ8XMKbatLw8KY
8w76OD9GTXCivTBMij9LPCmYc9RYQEN/mNiRegMXKfCII+qVx8aHBPGDVe6n8IyazipqzNU0+Ne1
jliesT+iu0GgZ+eVuoG27qtAgINgDQVQI4ZJphktCnjI3obkn8WlXZ6uxXLNuqZ2n8jHrZMkUzIe
OW8mNaYSwol45r2XQ+kuvzmO87zQxmgvmuvGRG+u8wgttAaQUCIh9J+ltIZt7VkyKCKddLxXBnSS
T1oK+LMBVi6dTH2BX3HfcfEPdHkKg2BJ2nGrc2KYtwUmrPDmGA3cyfyIIFWk5p9h6Z4CwMmgSgzt
q+Ip08elPFtJJZGvQxfmNS2J6M/x696Yc9FOL0/2YXpP76z/Fx6x+4NY7duGRnwIOL4DE87rVXoJ
nhtHyGCT0eX/agm5uzyxAOWRIyoM/qywIvXF2DToFYcEpDwgHdNh/MYxj7i0XnYur64Z1nNiSt2T
/e3w4Qg3XKcAqzYrOGLkVyRXtdxLZNA9RoV40ULvZtwagfWuL9/zHgjre5lrrGTqVg74wxs8439B
2JBdmlDGFqoOD3WZsb0phMCuXXuC7t05PKHILnDiTNGGx/jjndV+Y+4wnePkRP5FQ4Brcao6EPkL
Lenof/lT2BPgykHCF4NiYSRQI6Mhl89P4UCSmi/6fyg8VaKGVjC+oNB0KrDPVfsNqbBjAyugtp0L
7Ce3SJZCpzxxwXNaMYICYJWSWCjIctZ5UFREOE/pBTcGtzIKsTkLRnV/EX7+aeUFSl7WEstACJGI
+obrJo08ruzGxAdL9iden+E1SUUDhV13JqV2ReO+Ht9c73qR6Tmxn3JJHclDe3Y8l6jzirhqMD+C
K9yh39iQq7nGxC4lWZgA9RTi8QGLi8o3SfnmXGwfuvtl0HDkfuIjjLzPO3wQT+T3iFGeHbDAzwse
KJ0HleGQbHGzKk8SluopzpW+0W54Lt7QUyJD67Iz32jgVRqwxKc7ucoxAJmM19DUTnNtZlHA/x5m
ERDro4eycuQTIylUei2nEThRTHzdycs2hbqlCLNXkflDGjS6U9hgeHlAjZvqb8KKUlBluAgHgFvO
mo1Ub3D/dDsxhJX9ZZ8DF4zeXJra6A1BbplMKBfVDXItIbpHH6jtlzeWaThzo7VmWzr85vNswTo3
iuMHxmAPzw+c4zLrh9UNmQ+rV5qL8KMzKnql+cUF+WxU+OavsmtTMt4of9nqK0QT8mD63jtnPCh6
Aw7i6TqUGEbI5QlHPPxpOKc9JVHvIF4sOposr/vyab2TMVC6v9laGkpLiLwwINXQmVkbQFA/4qYa
gGxUI81/hxBOKUgCDm8nCiBsXpA8lp7nkIH+OtfrZIW35PdJBBGOf5HLHmKPxk5jbPc6bvaDk20Q
Aml9nNcyEh+gWfB03jYPhMCK4ZF7GrcguImFz9hTF7RImMpSy/vVsqJuIrveHL2WyRoO6bzqhA5e
RwbE3uLSRH9MUzY+cLMeRA/dR24EJpy3e53Tfu4UVzX6A+Kd2AVAlm1Oe83RLS2IDX3ZSuPlfLD2
zv2Oj8dROwpDrXty5UPwtVVJsREfL77OtNrvjTXmduh7OpkcoXZtNPX0tj3rZ0QDpLbjzDOYHUwW
t28Ho2mphzveo1kOfTFVOvPY1PA5mlh/ZzbNoYjMEhDVHwNwIWdLUI6+Ykg3IuuMoaNeGClxgiwg
cTtbVe//wPYwASTEm5TgAEAIKebrt6BQLI/vJ9WWNbvwuS0hm/AsEm/HslJqARZzOUPEn6XMce+j
0k6OQc4rynByvUVnMJdbAHps8dBh2EmERS/9DS7p9mhLbM9pDN4LcdLTkTYlUxElxl0Rz3KuC2Ep
aZzQOHyVqfQzow0YJok5BEXhP1hXGmEViKTi5ZzD9MO/gijHkEeshcM90Z2npnDKLYESm0gcmyMS
2pkMxjvYSnCIrqkqy7EBfKQ9g2WxgtxV30ADctPR38FBIWU59V5l5By6CWxiG5P7lp87s/8GMhfO
Ibo4dqTogK+sYETKgWlmeSPdduDsmqXS7JnADG3ctvdUnDz+tCEXjZSGv43kxxjCItmVmuIx532s
C/wmHk0rzpg3bHBSvX5L5rizQICOurPU/vSPvEUX3q+exAJQtzcq7EUZpMNEEkdDMLqiQuIL0sJs
rWeXMFtfCB9QiHA1j9qw9DOX75BOI0HO7IEEJKde85/HYSAZ8hK6ECku40mJITULOSqztE4vI4Vm
TR1CGraR63cpnN9JdY5tlZHVpOlrJVe4A/wDWidmAXCYqxtlMOlzFrXmVE1oZ6sipUPYevRsjhJY
Y4MYhC9lmi+rOsDilQlAgvIhRW0pQUMJv8mkAU5ui1RGY4SoKxgols1OJDlfSUvDM2IXioivvKyZ
5T3m5vBgnsZsgDuMaESn0jwqiWoJmyHAAKXBk67qdwVcxUstL2MT1taqWdCNDptw9hJdVKA3tNVc
5V+91BMfGeRJI6F6PaiiUbf9Yk2FazQn+2cOQGJb8nB4Z2Szo3jz336gzX3PGMBX2RCOfJ51wN0n
7rgyO+Cdo470uN4iA6r2GK4AfF7DtVachtAsD+aKsIoGaDC0WoT2fY8JOcsEuePOswiVlfYcxpnJ
4rYKcXJTArf2zaoQrsrhVnb4B+UJBb5RfdgtvL1QagoWoqd2lZlujaxN15rZt2ws9JJv/a+9JxCh
a1JQnKk30uRnSkBCllF8B5wu8HUnSR0vKz8BQ6KkuJihA8T5+C6ffCX6hjwF+ZrVE4O0YirMhKT/
7TtQEEYYyJc98yT+QnBKZGrlrQLV8Qo5+l/5nmcH2rUyPgEm4nc1b9MKgl3Qif22IBA0h6sKYFi3
KWJ+e8h0I2y1H0uojLrH1CdNBfBxRcB6HZxWnR1BQfKGRoxIq7hXfeyjMENFPub7zlXVCjGS55A6
UOMKWnRv2/SWbFFA+3yz7c77R6bQo0PtBHsOxhUsVgW8ZSs95MPWxg04yy6UVnZL64ev1k44SXqA
Ckt3S1uekEaqd3z459vTZDdCNxTIk41ZleWs++hLTjjsTvN/ng4SokrRIM8YplMpTrU4vqFhqEQN
VRcQosaMHF+/A8F6hMytVQPEMIt8Fji6+YwyIsjEpv7lHPgNSuLailInnqcK4Gk4DR2j31lbcwgQ
NFVIsF98WiV45uxJULpT+/5U2HWb3bMr6BCjv731BWyOLcLFlr/dIEu6DTtRvM17fjByyXJ6kuCv
LpvAvQg891o//RLOhVCgFat/F4m01O1U76vc7RCMHfsWxCLvUvtKeBfGMsVb1wf87DjHy9YniBh+
u2E0HisP+nwXX4kt63jd7Vc7wMNAsml+yD8+Q0qJxTH0zlij2znvhHDvnLgN8//7Ei2HknW9zzPe
c8elJSnrpdhILWJbtcfyd9Uu2CiqmqkomFdyx2XOLSrHsknStWsjxLsmOr3lCf+IVW0wPC2Rj6H5
4MqnsYYdj09D9YYPECn4hfU6PGTp3NfV+lSJ6/9XI9bGHkssk7u7YpAoM+F1hOM4xMiy3/5mKb+N
Q/HPi1O/LjUfYIUMX3aTyUCWD2wQFBoRshpTPlx3eMm7FKzkVGkUsBSJHkQUa8ZiXPBd+nOMn+Tc
lkhysWfO8TOlP7UJvqOr1VKEo3mKEOIdhPHJXYxMox/lXhUHyRijKtMeA6/TOBzWN2ILG6IwQ9BG
+vAgmwID8hScuahHvPMJiPnvFPxVOkmGHIaR66M0aObuprF20pCAAaMmJrwg8YeAJjSGX6R9ULr5
3a1bVvYhHUX3kAPCaurvd8NUfEeOED9EG2+0+d7C4+NPIHJcRrbrfwdJOoT0QNhrxmQA/y/I0VZL
a9HjW7egSSBN5Y9WAFSjLPckBD+IbHLO2yO5VRK0uOm2DlYIiwfIND2h8MNO68HSrZSFPpPNzopE
3V9L92tVeJKsv192WjqwmpUJNnV/P+RqGr/toQjNX8Yt2iLPM9wBf9Pgtfwh3i3evwnPDpGZx4al
7+iNkv8b+67kfEhOEnAGXb4vRqRlYR08mVpJsAtPZtMIeOaGZXpjhUPJtf220HWQHduNJtFjJaue
N2nAi/t/EbGNSOg7ZkpfX7bWINQGJ6psC0kmXM6rmjT/+Ju0hZ4agY32s+3fJWR8QTSmPO+JgzUa
qA5naqnwInt2LIh7Vqzee4iZwFCiayHVCiJQy4YB1arJS1Cvb5zmOHQkQgDdbI41ReKrI129oF7K
Ipra1G7WjlmbBkw4jJfs81EviRKDPWI1aY3rvugvqKy9FuP2fXkKL9EiGnfHzg7rcxI4VS2/BPJS
ri12nssyh+9Pm7CscuiDJMLof9eA+KfnqtL/Sj78vRSjRGjnRPasGNTdxEeZAbnPD5PqQn4cGwiO
Dm2/s4NU/eV/8q2eXPE26j77MWKFaRVzVWW1dee/rzlZspvO+2Zkxn92rcO8Hhj1DxNqHbXO/Nos
Np4eyQLwUCpi6r8leFYswIk17i4GqkeOJs1PmSWipJYOadyVPfG/pcjcX2tco+g17FDsWe+6T2rs
HOpF5ycAqJVWsidal2KsX3pcXO1NTaCukQtTxNR+Poc/iIY+eRSBFDa0XGn5g0MfM9EmfGZ0+Ltx
wHF9HOmg4V9fOa4JlLzoDD/l3nVEtgp18rlODMsETohoEf91l0uUHY501db1bw/ff9vF20PMTbFY
OlHnV9kMu5DjQu5tSwxkM0ychVE46TRtrPMTeoeU30Kv4nZNkqJuWD/Jm6OWHiNmmxvAAUlR8plU
T+8NKPhLvfkiHCQkXiYHzZxbYtfc9IFQcpEwuFsK3qyNQLrSusUItC29FpLezKqR058Ri8+NqK/z
oPI8ZF4wLd5oAmwn9Jwlc0KrXxM4l7k479OxGTRnIIsibLmF+tAWmJqS2LkCsh/dWEEriKnFEV3g
XZ2Z+D5lAbniAEqleiifjakoqlBDVWVtZAU5ke6J+LAM6VH3OD8mSVanZ5kI9lafv4eDAFlfSIM5
5/l5mCoaAsbeXYoaHGCGufDJfOgefz3UPRSOm5HoSb2x0KGZU2xMZ55IthhOPX8IbDsB5O2eQ8CD
rI8HTDSVKkbb4BWM4iF7Exrjc9Ex+3J0/REGn+Ze+RKLba9MKQbE6IxH4KGka/yL0ERWOEptuJIG
WD/gE481SzpQLSONhdBm5h3Zafyg7hgaXtwOGXlIhXzfVHM9AQIreAQesD0L0T050vTiZUs6bSBt
TmvaxizlV89Eh684BNpelAJiFVNAniBEBkzKTmi+qR2pbsW7d/OHw/76Wr45J6Ibx2kiOXbHIALN
Wlu+pMs3utdTrgZUdzEfQfnwIZOelN1kdnRbagi2oFKREqOshhb6NUVTaSFGvuMbVOVGCJFq2N5m
uNF6BQjEU2t/jp6+saII4vE46lsM23FOI7I39laU0Efpn9OeeBVVQnJyhpAf/T4Hu/QTXwc+YGIh
FA4+u33IlcoDCsWyuYq9K8OKGnfwByOSUid0e52UQLrggQduinMAVi0ofIey30WHdeBGfmU5LNJ0
/cHuZSplTeXTKegUJCHa4DSUueYDJFZe5D+Bc1FuZU3AcMK4do4WRz4LKR8VhOYjVSwBgv4wcKCX
ynZXjzsSwUs9FpKXYUNcvBC+DHIBp/P7pLuNH7qYZF9ycGj+0S6T7er9arLFguIjebgxGXcEhuYu
3lb9F3k1AXxbJd3rvG7EbYkfoFHRzIV5U7Bn42D8U7SvQGsipjFZ+HAzLwU4H6ByVTyHSvVmCfCH
9pZDon+11WpYTarkkUXghzLYWFl5ZpLbkvL/ZEL56O0kjwDdilqGLLTJPPp7S+oo83HqxdCwh9HO
3IakF5Lcnpd3oETQsJx6YKeGrRg99lH4lCRE/sfhSOzqblXf00kon/bXgC/0hVnhYcipPMlaaRAm
7kIMhBIkX2zOXRlh/UJqAE23VKj6fs3ZajNN+d9aqntTqNJkQ1HFmJuiNrl1L3FIg8yXWNSTF+ic
jVy1ah8MOjQpASv/HCYwV/qvc+X3w0GogQVg4w7yRzZ2XLtlhr7cWQ1T8fUaonAQJY9SYHt9Pv/L
h92AwYNoFTR+aGUhaMUiyWeBeIX35HVnGUfZGOy8TZEO+PFaKQ/05P7SPAhCN262PPJafk7i9MZV
OzUDfAVYLNXyWfTR6Kk1lzYi5wI53e3yCgzmYDakI0miFDAES/q0FxjVkDId8v1kFjlYn7KCTFzU
C1TH9ukWD4HH971FYIIdvtgn8VkGTsiT5GjGPQW/5old0Xtm8K9Ft3atxx947opX5GSC83LXgGZc
FSJ+Y7lf9yzkCLe2Xf9CmVXwNEptIKQSbWDnR8daasbYrFM/UW7NjfCKQaeaMB5qZMvbgp8KA9Cc
2PTPHDZtgYSiuGdtXvfI2bTL5QgUYgZCmq8L9YZErGoxObC9GQ73XLn+xEJ8yCFSaGPNzaBy0LD8
I9y+vJXDRLY46GCK3vQRMqtviGsua64s44a1ly1W+BoAAnSvaEwAQt33pQ6nxi42IbmxstvaJ1Rs
oXRRe/1N9UhW8gzWOvJxGTagaMIiFcQ2oDHhnSvjfHDkJLEPnWi4y2XxBxia+4jb1EFY2GSlhP4H
w9nVceaafh4iH1LXZn6pRxPiQN01H1RoQqlzztYPfo6WK3NIuwnVcgnMPxaU10OUj8vQ6PMfRKjl
s7/8+T6mNwMntAoZsXxNOn/bkyjCFvIQ6upVaH/w5+mK1dsCoMbQIervndTPgFn84zOMtVoVphel
IwzP4i1nvArRA1DMl0xuTylpeGK8jMoNtA8/3nA7zyDKIMgKhoARPitLEqSoSCl/F6JgX0o0RPNd
cOS8BgGL0Ub494cwyFQTqntkXRAJ9APfnf3Sbz3c64LUfTdy6u9l5lO3rvqmlWliGpv7z2un4kiZ
0AIupijt5928SC4W3JOW0wGVfL8ifWR1hHMx6mAM8QnuoXDVs8qdNIYTGVpfaCI3kIla08jKdh9m
oBL5Hk0cJ3dYr2Az8BM9U3bUuq9nyy/i1Xe7MzQrGCKvTRn6DrnjRd2EZ1mu2nk6+xfxGGYyqTRu
xfFvJyPKjYolJP1aaPXG6O9u6QUeR8lH1EV5tLgZpsNv/TYCpDdPqz7Z92zIobfgRMdlMzAeFS3t
1gLUWl4gxlZ0UD3PUUJ7xz9BkNFQP2WJT4tHlaumWv3mHZv3w9Y4AWHqzKkft+dqIj7sukLAqLjp
80Xf3MnjfE7b97htTL8IHswwZtK/N3Czx0a2NBtd/K/QzlLPAOIM+xj2i9Xj1uGgvGj2nJrr8wIM
HW6Giz4gD+yD+X0sH324tU2lphYMNxtM32R2Cjm+4w83G/BkNHWxtNenzVkO7FyQjybLQe2zcY7V
cBY/vpvQRvxSgiDoc6AOjYX+PAib18e/BY+AYi4/Fv6Mauc1ev+r98xsEgXqB0ZYqHGZbAalkd7x
oEEni7XNttnc13IA6vWlKnNeevm6UnhlBaJmqjKnnnm/lzZc1J8xWQs7Q6L0bq4L/XgGnht6c+M5
vo5jbjRtOGqsqdbJYPN5r0OWHeg3Y8/fti8NMRKolF/wWMTedeXd9lTfOVKrwxnfwuycybp3V+Dy
F2IgutmBbmaQWwzuXFTxM96RQvsrPwsGAatdSH+xOkTUUhV9CecdAclPM2jv1xkNIGJDpeBqf0GG
KsNPXEEBHHj6Ei9WAcT8JVJFACSRVJdw/wK/D81WVQPqGoV7onfwUk4MzE35zk8TOkP2oj4TNk72
c3a7Euh4ns+8/1bjAndOZcxP5RULvn1DRxBnAKbubj3gDDreM5COdjljalphZtR+71guQlTPsNXR
kjF6v4V28DeX/KoXZORFeqoLFXBf3p248eKNfISpoFMoaD6dHQNEOvmMCNh/8WGm9dKsfXaDYMNn
eKyt1ref7twQnZH45cCGGQi9Lmm8p0GsfW6jGrWtd0QjRuNrjUMGwQyuAzIoGjuBSljwoua26R5d
cNAuFP6TuH+NJu2PH2+4jNUgJN/3VU4jr5efoHwZ5WAsBqxEpy4LwYa55Z03A8Jk2uG9LaYFPXl8
dTFaWLa17DktqQpv9eX6WczKDblMX/oTNQhrhad2wjv3/6gE+T34NNRgT+at+fMQsun+X1LFc93Z
Fd3qvdtk5dqQYKcYdCwVqmZsrTk4f2WYwgMOLZgrBn7S9Zb+x4oZw5MZ/2vIY9JyNLrSZrsGqE0K
8BKuBHeNK6c+85ITc4OJXJtYSRMha35cNx+ZptafanJo400s0XCEjOkKQQqzf83rKKIhA+Nyl4+l
P+e83NQc7wjdHA8TiX7ZDBb5rtEWVlwZqPYbH+FfYOw3Ic2WKPELa6wM8quYnKnCbvRs5LsP3D1b
Jtp0YY/TsswqrVtpg54718ETsXmA7gH1FYOYfOe5A8BU843UpIsFI48g/nWswNvu/SP1YLXVNMj6
3bSKRdn/QVPD5M9tugcSoCXW9nyPyF9n/x2xPb25vXcKji9CY7jJB8dSpN3XMuWYfZNul8YrIr4s
3+krTkcFDG6JBQWhMnH9OerL70rKzrKfi1X2EEfVkVdQknJA7Z7QvKdns95U+j1L3+Co+SFwfgBW
LFDY4DtK1iZZCbxguScqbF6jE+kRW1BjETDLkXmWAQjKr1fqp9KjcqbAa256TLPVuw256QjJ+XBu
iFrGSogZbsroSws6yzorz2Rvd26w8Mexiid3dFoGaLbPSJAd9fOIh5VMKC9btw1dOrrJPh208QCW
sl2oubeAuZQ+sRUFqz6H7f7zHkUUfn57E2GGJdD3wUXH6R8dR9mPXk8Wsayiln4s2JmDEntZdwux
mlB+y+ayMaUe+Jr/+ggy8bS4u6cW7ZPUD7ueqZanysmnU4jvRQ/rs70AM4pCBxz71s6ex8tXVhSZ
4lVHKDfqT5dLjK0ERju/PMczqaMR9YRJLJkdNEJz+cH0G8Ac2ht2mquKsZg1SVwy5sr4ojc0tDw0
rZOM47pe1bZJYvuuSh/v8Z5C2xoIR+II5U9GJhkoxHDW49ip6BHijQS8q1BFWv8WFUcuAJgmP3b5
1gzEYvJUdbdqcFb6+e2Quqi2ssR34L6qIzP8FLsxhzByWo6xDJTe8H+KF4998UdFdKPRqlq1tMaZ
NX3DHCmWsjOiz7vAFUYTMpu16w9C0xm8diU0UMjt6OtK2IHe23rfV0mLhl2KHz/Tup6wXHW1Lskp
yyalUBndkw+V9ywIYf1xdn66JYDYWN0olQrLW9i61EHTAhQ+BHitCOD+D7hIN6YMsbIOiFhEwjY8
j9+OXYnOd9SIurL4XTo5a+SrClV3rX22KsqtVGmC/GWUB8wSNsGGjQL7sQp+cauK8cHxlNjBF3GV
TyjTvSbCY8vl03sb74l6Ld+GRR26k+7jHtN7mcJEZtTeFHmv01TFQf21ySb2aNvGHxIRqNofc7Rz
7zAopaCulZU9VEr/Wl1suKZaj//GY1Vq3kqz9hSxTANx/ZQAmX8dKgFQJwTTHUq0+y1tnRlDDYOz
UWx2aElw4DkfTInJ/Vk+gDuxlD4oGQzPwZccjWXD7H59LwaXCmv/FUUuYJg9Grsk8iCMRUfSwalt
8wkKsMztq/M2ApnnrpiemGk+Gsd/wLoejSFzHDEoUL8jMBBvzAtLpnH47gBcll7PtTG/0kNapJEM
9RhNeCC3Z95z4RRK1Eerk1H/QXxFvE3ThcOZTHlVSNRErlDR7eI2y0mEhFg2woJXSm2pwp4nO9k4
XAr9b0IGZeOuzf/omyiQ3JMKZbPGJWpHOvjhBV7joORJ0SFvqLG9xmbsnQrLi3M3v/u8M8AyfN7D
/Z2/I/XaWxxiydKSWbKgkEjz5OF+pWMXfXI/1Dd5QY5PseFQaTQgWCquA5P/wtRGTvJydUuWwBOL
5iD+PiJHvvEH9Ef4HmVj0/A+28JicFAR2BLwLkdsKyUSIxdE4KL3fhQ4+ft9NAW/UVZozQAlXkzE
uNgm7NNEqKUmrrsRE6SqsXXjaxnrIzQJCNvu2BtaHctQ3+UlCfW/Y6GUltgN36BQMW4f6TWlVoDT
YVG2iJzAyRsYqMqSXO1LtFATfoe+JrfB5+Hzou7Vq/75MyUCb6lrfGe5EgUnKx0+ZlxYFNeO3D2H
jKFRhdVwI3FookB3tFjd+ygnVBXkMxu7HB+cOVC7jJHjv8Wrvsb8A5akm2j4z8viRpWsJMgQYtxU
QnU77c45IMD0795sZW99rDeXeSYyl4gn4EnsO3rXdGNDMDdmwCx8f+lHhCbeY9FiqVItBjWjLkLm
9MszkSViAK09GbGPXsoY63md0NHgZb3onojAoIWh1CbD/nFko6F0vfnQ/3FVY/gDaOwjA3elrAIC
X5UwScB7882zasp5hkxLqMtngww1Eu4AY40BUD2QJwiF5xgh6pMSp/UroTZQrJP1JoI5Upcl4Cdi
LSdN1rQ7Lpy5JxoF0m9KF899rEcJJFvE5+Ss3LQQKT8lOTJCaenYCX0MgRD8ZYrhMvHGSajMBav8
BpCHlRgDEoYOCpPl1rqxgnAKUSir3lr7kwD+PmNhfPt6DRYD8i7eebJ5Cwe+uLa5J5iYWxExtJ+T
KIpO594t7iqs1I/qtQ7pY4mw8RT0VBR8zB1U8OsqD82vTzGmJakAaci8trVDMhuHA5XNWlQSC3s2
VA4ZWm8CGT2A050FjSST8xRqupxzcAK1f5VyWnJ3cAnYvJcUba1U/HsxYwEC/rBlnvAYmgfd0ANk
f+8hUVmzi8khrcz0SBLKMblDt9zFaHXS/HxYn9CQbSUp0wXaPN2KNVB0id+vJ+n5sIGGvkCD6Zt2
bkPIBDzTMXc9Fo5JNnzQm2PVaPzAQBBD1m2/3DN0gRA/Q1pqXqG64UsAHnmdGYnfTRBFEPs4Azng
RhvylOVHyhtmjT6GQbJkhtIzNV2M8NNfeICaFkt5dLrOOQ/cCNS9IJdsq6gEZoo+VaNfWyNN75Ci
LZy2uCDW74QPxbAhUBGfUoiPC8LE1ZcC6586izFMK0B1HLN+Ej5sM5Roal7kkeh6Z4+aziwi1Fkm
NiHoqY5pxZtn8GZ1vnue3hFRCxSebY8ObEfFAI3U7P76YfoX4vR/rNjshcFlxsTnBJpWU6pCeg2M
Z3/WCDoMwPbIvmi4lboQe2FTOYyGMQIOJnIg++enkJoSwBRxVb3ukQePGdogHMmsKtB1rOlLO1n2
2l+qNqxR4C6b4+x2ygMu/zSGR3DVQZ1Fyp/i92gVLHPnnwM4EyDAHWiDXdAHCuAW6Tw8b0Dc/TA9
cxtc+rJ1IFrwjR89sdmxG7LWSenrGnU5U4t5rfT68UftAGLe/E22Gxif7Pq/pTh51ON1Xv+SYadb
6cUNXmR+aFnpdfy07Ct0CIuch2piKq9+5xz7JNOXp0ftJRqcZ/yq/L+2/TINGJCOGsa7nvxjDPQC
UgB2QKZ47Yo0IseRuau3aKeRpugohjPxv59LaT2yPYbOe3ZJNpPt6oeXf5oTaXxl2At9To6yjPpa
tGlBT0x6Dcuxt+0r5NQaC1GM5i5Sw9MzclcFKxSiXyPTWeckL0GVu2vHE829oaw/rTBfvcqkJmNB
5Org2axfMpjofmBd3WMg3pwVzY5K2Lt6ZKkPEDFli9S5SFFNzY4zK8juaG6oOzxoYeZ0he5f1aGO
ZbpLVGPvvsGShIpj1a9+rHgaLKz93HgFgWkxEI9W4I9Qln+v85PpyesLjqt8tzkXKjoyo0eZIOLW
9rqDJj/F9We2U12Qfx0ud1L4ovkL/TwJ74vQPFLZ+7Ppo0me0GQuWyBWqt/qHjLHcFBj9e7LD6qG
217dT7DyCfVGYPH9As9Zfdqol/ZB0JaRK5lJ3fsmmp/mQuq5UqMO3SQsHco1XaCmsIOFbALb3E0C
/lNksq92wSUZt1uLmSfAxjm/0BUL1loXnZBRVc8JV0L5MIX6gakOusBLufd5+N/rVtCCCPpnEl2X
kcnIQDDMXj6RTzy4m61HQTXGvrq6/douiN/Rz2AWWxnmBzweTnRO34K9iWLTuY+kSSso6gX59HSd
al/p9ZIUizaPQVRWemDp/ReK16jj8OIPkFqcO7mhyv+BjSTHUojKiVNyNMvradwfXAAHZRYhIcVr
pdqa80HKuUc0AoLrrk3AxrE564zVvIYycrWr51TY51kv4nceGHCIS+OoGxIdecQdUVLmXTY3nLO1
yl3MCUrcHxHWYBwV2N850Vgnmq+uO/ubJClXin2dssa4qhh3O7XbFuvpH7qsyk4boc7PuG/uwwYI
VQGkpXQI1ks/s/KgeNlzQ00MvvTTzHRF17R2n8Qhna99AfyOk67ptKddI+M3AIinWv/sEsz8/QTR
w6XE2TmycXWhTpC8QCBJ2ltwKhvZIIbDjwaVRis0CiVzqzJuopmdQtapIQ9ndKrOVloC/lCxNlSP
s/4ml0ftTD9N3kUIshwT8XKaPh93sJVj9+H5h4AKslU1dYTJxSb5GOrUY1N7j2qvZQzVM8fOodte
avidfEC48MWNCL8tySTTC4/aSuCt/tyR+5aFtdS34VQI7gmPEKnwHR56qg9xjLIl6hnuBsUZrzSx
Bhb5o50KHZQv0UNZur8eMM7vQrnTSNxf+2QWF9FfdAP70L5JJE+6ZvFSIFzfW5zpSaUgfOdvsMvL
uIyhwAsCn50e+O6XSzlOcMlc6FOoqTJ7gI7wn4PaoFqPDGXiI2rgDREnhogkWbWKSI5ATV6kTmYy
PR4vFUZKXP38o6+C4nCztUZHvQ1yI0d56zaS5/jSlqmR3opjXXzgHGBicrINIfNNA7CHbctp036/
1G5zFLkbxXoCrC3njr8uRWG4kUyHVmWd/AeHkpUprG7farCt6QWHysor1XyouuQjzi/LmJTEpuqI
7MnjkT+SvHy+QB6LxHFgBDtK0BfHHiOmiA+Xq+ryiPTShfhy91HJry0tOhevFzVjEDfhblNk3+3z
cBDJOYXiePlMxbC7nXVIyvWfZNzp97AUy2pvd2OXkNmxTEC33v4J7iUYrFk7m8SHdAH9bjlda1NF
26aYsAHiXAeJTiscGc80AId30hAT7tGMajZmo74ZN5ChKuxmKkBW+IWUAJWkZGHVd5rW0KWfM/Jw
Q1K8tzYcgUkOtj+lORdsoFYUTcjHSdYT0+35+cv9MQ0N6U0jIFZ2HUBoOrpRkpYQyeopcXrwpby9
TLkiuQPYCwmuZgskzvjnSDfZ9hRLzXIo1BUzX64rG3/bjljPUOL9qEp71e3NwTy7UD9Pn20mhoIQ
8hCn9e6BxLMj+0owsNgN4C4os/S0gQd4mE+qiEMM9vhNoKsLqKokVkUcuisupiRFmrTmHCe+ttzQ
vdnZVgfzVZn3oSvMCThQaP50d0GxwN740okPx4O22RKcVRSxM43LN/+3Qf0o688wo6Kn/tOtZ22G
YfcSdFMQE2BhO/Q5togOgMoKHB8K1zC7FJiKytYTaMmSmdtYYPT7chIhkyLB4L1kFTVUTIbWqpTN
ao1khj2QH5KhgwjfzsG4UBCPIq2YhbFgQCyhoYDBH7gW5qw990n4P5KFt7kS4pdVJI/5YV2PC9vZ
hZzhlLNY5Ne7u61pkb+Td3FJe2/CZUqPMBlP2tCoRP9IzXRyqyfHi2bJ/pNclggxxtaP7APZUPGO
rx1/+fEWRBVu2ZtEJ8SMx4JmxcXy34N8isCYcuau99YWvwliJxS1ZEWblNer8zr3ZRGYoyx3EqCO
WO33pu/U5SE/tAnT6TFCFVwqRSRo+6wtNqcuhTqpqil1h/RC7iTNa2du5GQeUSd3+cATmgbEyePv
ATKsnXdF3NqwyObTppYGSiKiouR8DOhOFzJQr6bNozTtdoQeG6VaMzmuwNBo0ysFDWMFGcMFM0Og
pN4qRpcHOV0+9EHOD73C83WZhjqJUF6przf5COplqIGqob+KipJYLig7hNmlBdMk31Bn7KBPsgIh
PaTX69OAP59uvROIwX3gOw97RY0wAbCUI18822o8UP8NG6dni2AjU4mMv6jdrvvajiaPCrFfL64v
5rxkx5DS0j/7lIJqcMvpLexC5jsbWvJno4taQKH3pv+CBBIFXS7Q8lyNdKGuqiWwQxNjH87ggBX7
/uOQvzkZXOtVgK67DHIoVL6vc5zkyvts4GBVtoHpgx05m47oEj+A7ww0sDmano1wlawzDedMSPZ/
WdQBaX7TW0x8QOwEzzc5o6sZOHQwQSJTFZf5s54uCWhUXhkMRsXvn+4UZSMP2LOLJVERI0kwDGwL
Ll6XJyBjU9w2/yclthrYjZzEuEOWxMXbeGxOm1tWzs1uuvm3HA5vlb/DAp7NBHjw+IKcoCuvKQU8
BKVbaxHVbt/eQ0DbepmwSAJ/ObtdfJmCtB0fGJM8K5Re85kRmpo2KgtLNONhRvgar8SLFKCfBlz8
wwIyhLfnQbebTzF4IlH2ZraWm3U2Zdh08dcygYejLutFODER9WMx3OtA1PPalRB91DmOyaVF684R
/eZmrXwIvc0urZmdlk6uyjpeNVTvrqIHNrNLxOjKefXMFlEVeElgVlV7YqHzreWtSZt8Q/6kqQuR
WTqNE/5wmW8BgNesZsFeH8JbmFuCZQF9c6kczzSenyxOji4ybK89E/ahVFb6lT8mU3+et1qaW0AO
hubcat9IumaITKLq0z0FiMoxs4+ANZqV4ot42p8eLrNQcShhDDQ/TtfRyWP2XYjiUnpGczkhUbY4
gE6/FpVq6ljzMQ4KTbMOFqSgagsjKOfVqGFf1hGjdrmFKm5Q/OWW6S/LC5jzHrtBZlV0VJ1LDL+h
U/Z0pK9iJ12Vqf+vWr+at+7sudBl9jt4ll0boGNhp8uUSUg3psQLS8vIGXWCFFrv2jogVC2Vrr4i
UPByo59K9rutwSV3bltT8iIhh8587kS/JJua5P+U9QRydnHLxRow61btt+3PkOLYP+dHNBodZDRi
iFyJcMjsMKqGSTxBX8qMSeaP9a/ODHfuBC2VWg8D80hRszNUJOpQrNnKEsAcwYlyy0FNKUHJpbB4
HoJuW712i1GRyeT1jUrZooSkm8yzZajCEAEMEPZPJ6H94KeoAJc6LEGsY2KCdp9sVtLbXlKfAFzq
t4PrBkW0OmF8bZ1+M0jmicVwn2FO7N2UfPRE7sbpacaTcIGtZu1p066dSEbJE4yX4JA+Vm+19Zwu
dYDpkVemAXlZBegSNYZhmgzqi1oRFsgx8cBZXIpZfjYjjsZHZuDnmZwGCKVzhaPsLao0sB5kPARL
1hOiGSyxFj6CHqz5ajqP6Rebi257env2KnXJ3H+prTcsgi3Q4uXSw/isWwrIFT82UqC3dwF/jJ/Y
s5QVB5ZIN4MrY8VuZVartCGGp/JK6ABx3neObfHwq2WmhejadxFLpPjygMMR3yZd8ANcBxCA1n3H
CFY/EkDnqXJX8ugiiorL4wnDXIElGIIVeVHO+lhAjNZye311PPd88b8N/JPpUvcn0B6LR58FeSl2
XImEEnp+PPrGnJq2tQRxyjnu1SEo46GEy/NH+PVxHOqzgWdytDC4N7tn9axriV7JI39ykOJa3rZo
dI9pD5RkhbAFN+gEOvLTsqtBSi1MzSt29AFDuMWiqSm3de+ggGm4008sD+tImYRte8hqdOMtNoVP
bAT4kXzfOiTYjQiGY+8S6i8jCcmX1tym7L02anJaVbqdp72jKDVMM/K5xd+g+t17oBwd59QMn0rp
jPnW3viN8C3o+ubwdQf4xzJZAH8NTX8mJNAI0V+CBtHLrf5kQvXPkMJD3MOnH9T19LBEgm+mHPZ+
BIVGtAC1+gP7OcsVJcxv+xGEMLpR60LmwDgKaQRUnvlELAMl9i0bfji+TZIqe8PAvdlI0r2JwGsT
e6doF/pxWqGfLTaWo+a7m7Im/xOFgDc6IJ0SZsoE6lUl3d3Xc1KCwL34s77KZKXO1T9dwBgkMowG
cXzUwlkpA68MfMZ6qBD33N3XL6SF2rdSKKzwZzak2D/Ga5GLLaYdJFIm48QT4+9oJ4FQK6Cqa+rP
nqzV8d9h+gKkr7mSYuALkcWaXt0+hzSB1pxx7Iv0RMCmjllOGPFox4fyk1OowkvPCLKTThJZOUCa
ZEr70NbaIc7x8DLdBwskntccmFreWsOx2wvtYiqxIViyNat+56mTy6cnr4mATarEXfBuSwEEuCry
Yca1xcYRHvXP/lsoSxELpqRzCtxp6KZPYF7NQSMYj/3OSN65MxpsaCF9a9UtdhtfnTTk1ONm6G5m
InAPCj5Awh5BMZVkh6VfnwQDy/xKO2G645IRNGXX/WV6Hb5loZjVbSa9umz3tG80/MI6K2fFYbJN
MW7XDCAvcKe/pXEozfs/4l79KSpRqI0qFHdnznIwOmcVOZ5kZ11HxtkaLPVbg51NlvazybgcSiZe
vGHJVaQ8/36k2lpsIjocQE8k9L+TDnTETqCXJAdvRAD2m/vb8ClOrotAQ/4GQ6whvGN8axw6Kme8
MdtMKtmTZF4pDPXXInopibJnQtGpgViPc1UQ2QwGmUKz2bUoi4IJ/TFPIDQaZeiX0KWj2C4BTG3i
c6Wa2dDHD+4PDG21e/iEkiROup0Cw5hQPQbhP0rSmxRPQJGRHbtzi8zaOFqpJfnC4JuHm2Ika1ne
LZhNlIc9ctV29un/+gBo7d2HN3cl5G+Kdd/UzylZT16TKSlnUGnOoqU52lPbtUL7fS+yQotA94Yc
FIQoM2KnZcfErYjAxlaun1SpmUUESgmW63jNdq4xd0Z8K8oqrTROxvlgYBCZ+IIVrG2D5VLPPw1d
IqkcxgVs8/s4SmIqHL0hiV4WjczDADuy5I7EH7D1Gg2o52uqvRTthX1YmSeds+I6VVE6lWwKlz4H
vGNv1/v6JWkSdWuRvNEuJLWFOCXWYbaazEhHLD6XYaA2zGv1GTzzWdalcOuN1CHuI82iO5pfg7BN
Hs5PqCnhQzgaXUBGVmnp/YhuVqyAw9fh4gzL156ui3lbfne8iKszws2rT/Eu6vMWZKKi8tmAWHt3
yXeKUDbVqL4XXlV8Pvp3wjKk9cZ/PznU49XRMjmNcCX5xckQus0OnQ5QOLgARCGF55w8fMVx5AeR
b8wq/x9rWCw4R+oxxYgm5UeGiD6n/RJXhY3G77TYWz2xjQzv/qcAUc9rh9SamX7n1XypX/C580G1
jUTXuGicvf7q/vicEN6r2G3lgekxdReZHYrlJqcxAO6jlUPC6TdnHEIRLtyrpTjI+T8gzQRcoylG
qdhmohKxa0k8ePuLAInVMsrLyRMVUpuzyrbvfY7/8tGXhqFf3IXn/edx9As6HpTqW/y8SBJY2HjN
lD7tllhQ1ulqdvUdSnm5VsI3B6ZuxoQaSK3JAsDRmIAJFZH1AC+pfDhWvrNGG1m4pfVko5sOH6X4
K0tzX2u4TB5RJbxI/d945Many5IWZNnHqehTJestH2C3MaFzzkzM/cKtfMDYvXC++ma4dra21BmE
wHmpnUgNUm/WNzieb/EhCqeX+uNCys2Dpxmkw/TCY1dRh6IveQ0Hvc5zrhdmcOaU9glgxLaMZr6F
66Hsspxu9JTzlOxMJkNKsJ6U8WK63ugvE2ShGcqQ8VeYJyS4l4DVlodsWNpApHVnWJF8Brqeq4ZM
LYH/1m5Yt/l7EpVZnRPUXleYOldsKql8G/goSFEHVze9t05O6hzrykdryNzu6A2OWzOrdFU9O6i3
4+1ub5POOMJn5cQh4DUCxH7l8/WYCm4A3zG0fL/GkhcOwcrG8LQXbd903bo146fexRRYCBKmrBbH
kWoKRNR3TI0RUpuBcS5rhRiRjZ8NTGIAUqSOrtzh4xXNVNdrY0DZM4jJuZFffU4lgEbjKPhvtolO
rXP47rDm/0K+qQN43AcCXtI3JAnmGt3dVVHckFTLiVQyhOd0k5Dg4NCQgFvjD85ntIZEd8dCA0U3
xHeYElOZYA6cH4i+yxVfPAZa+sTGEO0opaNHO8rsSLBMcFSeZOwh6u8Vlh1S+6x+gS7LoSkJ5BFS
r88T3BLEroUWWDLzREgzoiM6RO+zKtrSPbV6qgJbiXYek/eRZmxKsfobdD68B59WHf2oP0xjgeQp
j5tymaYcRAvF6Tx4cYlNf74mEATkjFVSGy7EI0YyNdBTJAbywAOT2SaBBJDNlRDlUehzN+jYR4Uw
Dnga2o1jstkfs+fypEeZ08KwJMOKuzYwDyX6YaYdNG+qyLws/uH8HmH4/GSr0VpK9uW1u3xmF5Fn
UUHyTGPznck73UduSL+pyR3IiF+pfYRE+1G9Zdj2U+Wl2pKSP1eU8nDixuXDQ3dSy6YveE4B5PBQ
d/TW3kPmdZ1oLChoJjtaPOevAgZUrCdGJZpjEJi4KghDJwROMZ4390/G4XMqsZzDtrjUEYvsIqRm
rrYJzZ3PnzFWVqi1wKIqz+Yvn0UBLu59sL3XBUoyg1/kpqxRY5SFS2EqR5vJxNtA/9npn3DSjcLg
Z6AEj2mIf22RLWiqk2WOCIR5wqkzRWcx77l1cNbSghuIT8lpIAbd6sbD2S6Sg1b1B0LmvN5muv1f
8KV8WoTvJAMNu1rSROAduPYseplHCavKmvgGhNwPcvXiOpUKIds1tCM+wk2OnMPbdP6RAmpWaM2m
MUAts9eb3aghG+x92TtG4qV95Vqf6BfCCqqqTjh4KCrAaUXvhllQy1Iixv/zmMAGHiY8sQkfVGnX
yh7CDD6WaIjh7lxIwX82ZXr1+pTrn9IbiTWWFrwNhhrT1YnQ4aFn66Sbt1aN+SU2VicMvsr/6TeV
m4QfaJrS8J01u7ejj+bwZQAk9rr+vTogwPYwWDAtYxnfsX/CtJrfeEnvgsRO/BvelGqHX9gmFvkY
jzUCQWZ/keWXKl3PMJmE11MBNWEaSnGRFGRTTmuhu3jJI7CX6IkzIerdCbzGbaeaR9Jg9rCJgzXo
9zWMD3c0p8lJvZbFf22EK3Qo/WisJtQLTbfK/NI7fpz24vXFOqnfbLNkwtRmWG45ki91CAzRPSe9
sUCRaGxCciYZrXETeDyoCgDI+Z+Rt4GeDY0UWijy5+0RW99bdmkOkHVknHynQQa7xLTYLY9OYchY
NrbxbeiXQ47RpOA1gaONa684YtT3OuHki+x7IeVwM3Xxg7CksByeiwv2K5N0zL5UYu/6AHVVrZK2
oNGKLVDvwWlU6ENHEUjpgYoVc5fmFP5NUXRmW+idXu0aPoyOA64w1YKHCA+j+miarjOaaFzx8c1X
zIGOQbp86rV0YAnoaUsV2CN6dwRPqUoJ+pKxyqCdS0UCe7uYJd+dIX6/we3BM2KtLFHzAyMB/bJd
AxDi+4xeEtmQK+0fijPw8qfBSI2MbRGAS366ygOnFN8JttgluGtZfiZB4WmUXGp+7lfRVnSUJxFk
U29NsJcgWfdzo1gaL433eYWAnLRWStZaF4l5xJiaGKnPtC5ZoRg5t2SjybhkRTdaO3WFbi+kX/A4
t+mfOjMjvhP1lHtMdPmI+YI2rgdN3aunFS3TFd8EHJWQMLeDYRgfb0Nxz4vbDj702REnQeuGRPd5
BpiFupxjJ6gzT4vTytIa0PjpyMwSal+hjIMNQo7vH9yVzbe1VUGnOq56VS9LAUxcQejyBMCCrU6j
HChx9qdNRtnapojVeX51NECCcm6Kbl1OfsYJ42bL61PYpiqMgQe6y0fg+ckHZ7aZckKcN6w2go7c
eHxZN7UDVKbrGF7dL9JniaIcVu5Pacodb7CtYnju2CXepajjlqbDlzApK5Ugy9/H5tv41Mhzwk29
v+fm8dIHAm95uMCt9SoZULCCP4t4FqtvO7Dv/v3bD0wgsMBiT3JFEufaeEEGYuuhk6yPMqptSNUT
CsRFnClbhUhHpZ9vVmM+mS5XRMvlurN46msmBWvc5pWs56ner/71LcRbiGHE7SoZF8anNkQYrdN3
r6pnpkIZ3edRUWWHvqE7PdZT8Q1lcHcMjD6XWSBgF/zsxQghMa8/sSde4Dq3Sa7Dzrc2v9RO8ouc
1pt2A9uFLP+rX5/wFcDx7MFbvBJbkOI0gvPLwFjZNWEyHyUeSuDkLB+NolzxfdAhOjIw9+uxkZVa
DvvDoPdLIga6/vo1Ibuaz6c3wYT+N7ODBzzQLHtsnd23/fODdtla3VLCp1kjf5dUDSNHr7dcBRBl
38/9f89qHwNesLqSIlE+8AYgP535Qri9kZipRHAX9QNX5eQYFGI9kJpZebw+MOhploSPmi2LhPDq
YQtci3fvTVYSjoNo/UiVKrAiCZrpamYFy1Vw2zG8sMTcMIBkW85mlsEYZGfOv8MIkHYwvqRS5Y3I
XbC95vXlE5R0eM/2f2GUU0FYAjPqqcW7zA++bZJkltW76onKiInzYhc9wJiN0Xupys+ab7WXhH9W
w6o5EkuRS4Z8pQfeaAKsXgOqSQtxeIkPgHSAfPnrptFFHPwGSRwG3ymuyt3fnOcxMJyZqT7js1u4
Z+ikDk2CR+ndztoRML7kyB6ncUwhxXsoF+tdujgrVChydBn6Xl10zHyF7/wizrp9dlF/wkrpPVc/
Z1fjNzKHC9qZWnFeoAlnagQ9mqm0dsDVjAFNuA5K/OovVu4SgSfmNiPpfotiAeXtCTesR18ilKZo
Mm/znLfj2zbMj3//GqbN9iBzsdJHNZjPm9KX2kjidCYJUB8FdE27TXWGvZb8vxMX+GmTmEJUMlBe
Dq5RFfay2+PVf+6IBKDwAjlwHjGLdJTdCoNUxvv8cAmu4Cp5JlR9I7Bn2tL/xv6xl2j4zV9lOpE+
yCj2xW5OfUzX1jrZjS6LTwsdWAXufVC4cC3HJj3+wJeaoSfVEJxj/NvY0tsfoUcQ7vhHOouzcB3/
iqEb0V8MZUivgdwaxNS/3AJ7VKT+JqNeCxjFP/8GxQlONvfdOhU9KiJiQjq368EBx9js6X39KUQc
iSOe2esYD5fPf/wZxW2QhEw/pDC5ot8YLITnzgyxAmgmUeKOYjmUWrvDI+XiBLZDscMqWx4K9NDx
VC/9ud6CbXRnKiNuAbZw+JrYQxk7BZSpr81hwQ8BjYWAQApHd1uvCDTuImBTseSpqKF2xS04lXvz
t66ePC9Q4fo/t1dOR4T1wGIoOM4JWjSDAH74rD0LpoYNlvi0fRB4NCxQv+X1rouY+tBSX9IXX56V
tmAlPKGW6tP/mqII3PUNyBask1/ZhBR5gQOguUXmexI9vigrI8+ddVY51aIMpj1vfeevLxl6+3zc
FZgmUeXWa0PhuMw4fh6JGwFl8Yqe8bzwnjafUsb6vsAm6UVKBpJNWAliajVMgdkkeFlaKUC4a9OG
Fk47OJ7JMddmRnlgupeco7Z2FNIA3YowmNPUPQfhrBzgpQ/0/KJyKR2d02pykVKxdjug724/eIbw
PBbh9V2XkozWVjqRuR/4UZQHOnwGvK22UWR5lZdDYi9AYxI1Fj84Hm2RuANKldfhg6fvCt+lE2SD
YnLYPAc3MxaghKMW8VJ3NtFvoW7xylIaoli2JoEFC08jZtpRxLuP4eZd/gEs5Zw1QO2EpZvMpG9L
97l6AM5LBLP8aRxHlN4JDKafzLw3SiD+n7gBtUkdQfS78H/mCZqiBdrjv/7at9A3idJLSApxHhim
dA+EyXndvu+MbEf8kxTrRittUb/pHxBJ6pWhT2QVf5pH8wMYDwn/o5nFv68hJ6EvF3pH68qPWejC
jwvCMrEllM4eEHWmxeaC2mLfV4lYCy2TJfHJI94YxFQlxcQaeUXYBd2cOFt6Z1/vJ2hUVDEfjZju
rXogEj5GZQAgioZzsuExCDRsVq7zDQf8Aj1+c5kjdECXkzLGjvDCrrHMEkn4KkEYot2Uf3lrsZVn
NrV9j0/fTbzeoYmBU2/NMA+PqrshjLGnBV5Ag+oMOhzpMTgkN8Wbkg5BmhXlEgSn3THImuclJiRH
BEFSxBgzylp5w/9FSacpIIEflh7+9ivdpUd7ObYLdPV7Q2pSJmebo1GwYHEnFgWNLWZxPmDVT5SP
LV/UOoahviq179i/QXCYgVgeb7DKCQGRfp2/VCx4hHANDDvSVHWDO8oXqTeUljvq9oR49D1483jR
r1gYLnX6714iYEo/FO4sy+RnNqkn/MzmXgvF4VP3GqfbtFSbyvtVgp3KakuDPXeTCPM1oUXblTfk
FQ+W+TqMAS9JN+9nsehkRVW+t6G0HVhU+Lard87EdO0m+dm9pIT/38qSupaCNRQXFlw19TzS9i8O
e7nG/3IkQgieTxhsXDYKnpd8BWqNclejyvnxGG9Z+mwGnazHkOuMXGN/YVJJP7A6xpl8KQTua7xP
dbTo3jUG4Y8IwZxIIeKpjtp+/6BVGdOU5qUB59JjHG7aGQd1mUghWWV4/KaYAttPuk/CKx89JWx8
/Jb1BiDfAE5xuGRqn+E3A/2JdOoKnMCmxaHtVWiUCGDgO75f1mK/uOClkqmFB+sUHRUoGUYtVGYh
ipkgyaM07tXcW4rs8ozxcYwfHmQcMutl0w+XGLQFjP4rP7ULDuv8PZywJyr9Nms0LZrPY8lPnElf
+P6OvYpEkiwch+B5dd3jsN0L/WR418GJ150RHbttPEX3CZ0aOwM1Kn+lZsySix4vbw/+2m0V98J3
kC4OuAgoNvmQwmngohs1xUCK3oGnzacryQmb9jWkA32T055gWyPfnoDOJ1ErKPwQzeLg+SUnfFBp
IGjEKdrWImDtJoP5C1BkoCvHin1uYBXNYGSbiI3CrHFUIMZ5gacvhav7NOyfaOe/mr9R08heewKT
71tncPxLFZT5CUPuAMp1bzuffO7sDCSoxjgysGOtn8ljCbEDqD5LdJ+F4BNq+MHsiu02YlvzwjhU
ZQ/i9w3xtmHGe+Ss4yeSwTCYd7Nve3kvkg/VPVckJ1NKB1WghknQ1AZ+tOO6KejNnN/dMqqcSVT7
8N1tRA5YQ+vn8EEWuoHEqUjRv4jBwzQsqn5/Jm+262SzWgT6NZ5hsyeiZiLLLYD/WriTwR+WftBP
7ezkKlWLndQa4P6rLwdZzzn7T7crlIQh5e6abkHtXn+pODw6neZ9vVLWqJnksQrM3bv7uTTxlvNA
gaey6QZ8bC11fcFj2D+Bpfgoq0fYLme27PL4lboJAXMZwudZY11+veFqEXnUb0bYlnfYp2zY6JCR
3ajtZO12KXjWkDPO+sKpN4J/D3QJ8p6YxgJvAvuaYDgcJ22etEFOCPmMtvTtXl8PCGYk2X7s/DG9
PNOrR1fc46DL7qPiC/m6Q24OG+S28mwDBrset8Yek3ELd1ppRxJG3l7X01wzGTOdya+nPeBZCbTv
ka6C6DsH5k/y+9groX2vwhrRLLmDp5ZqO8IzVik52U9E5DYgwf9TAZ3iaKHuYxN6mJbm+2pEWA1P
Kh+3wTaD3kG6mpPNezC20UZFhhPF7waEq4RC3bduag1wAfHxPDbxPjdbTfidPoiT970Bug+5ZrMe
/x13yVYkVou3vUojQOyHWkt/36BV0uqMxwbiFMoVQ085BxnE5zkhASIT1RWhB+JGqxvjoklBfGYC
Y+cVepKwnb0PgJa9JyIL4UdZI5Ab46lY0PWcULXWEpfsBxo0S5MLrgJR1LuAcvXO5E6tWvHOBq4K
bttRIyauIuIE09oN8zd1iht1N6NI3RoZL6lA0oAS6aCOfPbSfjNoVeXDhlmb1s2XPVxJNUjmh+i6
w5gAQgSyZMaItcSIg0pWvy4lzvmXDf+ecBLe0iP3J27VshtKjud8orN8Qzi4ty+Ms4M++Z8fSoqk
1ZMQ/8lkEpro+oPWpbOokotXyd5KjodoNIBTiFZ/9MGZQzjcifOGYzThkT/MJCW9aUjWmRJ3Wn/g
eP10w5HO4IB/2qmhPC/z2cCC0krOuKEtE2X3LfxLvDOs6akNbtEWoaow03f79Erkae/znk91aboc
lpjLbv6nY0IJmpQxSdDsLV3dikM1knPe3jkYw6RVtKzlZdt49nSdOABTlPgUZToj6lDAbj4CAelX
f1SGHY5HskB9U/D7CGCnTWc0s8nugOWXKrSumvANEDvAdYlaNDzZDqyq9FsFHb9XPPCwXFJ/NQmp
WMAj3hlV6NGciWuHEB6zZ1TmAJHr9seNLlZb1KjY7D+yphuigMjhhRVXjQNEItQKm4+e14ITcHLU
Egz9K32n6t9ovkK6TXCQdVLVkm3LtxNT0Lv1wRmer8oY0z5OnF3faTwV8ZBPZPR0tE/v33bejrZC
wDfKQengUlI0R5/pUX8p8D7UpHAkrk64JCdQ+qkNJ0BKOz+TTLmGuuzA3s0AQyI6yQFV0yo9iwor
UGQhaBppER1oGdR9boZDlcsQO9tsImPWRi3i3J9OkxxVVRfoaULSuA8O+fUimUDcfWiDPMa1o+4U
s52YyE1XUkgebkpN900PLTymdqE5ddVT7lVkQ9/86h7eiV6Gjl5ol3uClL9VNt/ALguptj8KUYs8
JSsXQnbClxt1U6dNKLiVSea9v1oG21pE4cfmgKKpk/W501W+8ziYdZrCwOEBFPzR+JPQQu/ueNJe
WMCjNhFcas1EO1GfG5uk0hYMG22zFUddmfQh2aC1E33q/evLuPqWG3vzwR7Z2RBJv1oGJYUjdrTB
IArM/fVXwWnsqggDZE/lTWraK6wHmofSizoZn5hTEpkFK6qHFApNI7lL4DPYJjWsymT+U0x1FdNc
BzuXW/dV7O7V129dB1N8N0cfK7O697Qs2MyiAQA6ZQ4zeiszmbRMvNAnyqszmTvTkubwCJUoJ/hu
XJXWazoALmxkb23iy/2i4qk4di0Kxtdn7tCoHa+SlQ7h8OLGc3O+r0GGtRtbQ5v/5n1yjh35dQqu
5g0dGk9U6TNZVq2KGY0frR5ecLqrDs0lqWQb3NvP3qAEPc5MJD/5ba9lme7PvtyLZADVkgBHDTiy
bATxhgGrz1UzIcHWjMElgt5RXpUhFOnAjUeKKwTCvME2jAT1vWI2vdXSEXS1Lm/wPbWsNy58QmUn
Dthu+Hl5cDChlwbXWK4eha/r24KOdQ31DcHYIeFIwfd3p4rLqrtCbVygxe/Md6B2P4QLZ+s0Bwdy
hjRuA6pp8Q8cXNuvlp6hg/mFY50TOfm6HhtGH2luWanvsQmumAP11SC+grPbHsSz6QazclRMDqPg
AcYOgnoH4e7Bp2PpzahgALPx83sKZmXs68acA0im8rXZD5/Oj6C5pJSBQdsl8RawPG6ntO+IAw64
cik21JZyMiGoo9fMa1OwVUDMrbnsp/rm0/4wDbeNSSKWbGNmarURxtp9hWv0uak+wHupK8gD4KkB
b3ri6c2vmU/cd5AMkvyqiBLDI5VV5HfX14dQpQhb0eL0yGDBuXTEjXh8ZGaVluR2GpZDOyykoi7I
EW4KlvHJzd4MYcwFS93i4ijix/y6CdnsX86AR6QM5cKeIVvRVIQztrTaqzobjBJ049o4CjEoFS97
+lZk6nAclthLuxYhExVNQtkBJLzUPWkP0Hm/bpOjVPa3sQp8dQ+Yyo0SALvfQMLz2lhecQ4K2y9U
tIImvqSlpgoUTPW8nkkbljqqqhrzaADMVSxadXzHl1eWBddDp8uXTZdFNYvbybn64JoZ7TvEVPiB
mErN027ezX0cxlr6OJkds+fZ+5D2gFjgLmA029BGgOuTqWlNAk/mrr8c4ULEjvoBkDnZES+HaCt2
iHczRalRnFvLQFmuv98KWMVqCG4AwE5lGR0JJg3SQj0DTqQa5tDR7fh6TPaSTbsiT/Ven0JehmcB
H52M3TByTDYKUKYf55B2BmbZvLxqhAp9XWeWcGVkvYIQkX2/CpTU3mCAv7jXMBGPwAYNykX1Fpod
03dqggbzyWCC9nt2b2ehWPswmyrlabURiirbWODFvGo9cMtd47wi5thWxn7Mr9RzMqVHEHzD1lg0
QTvN3FFKQqP6/jf7/TXgBB7r/MuCTMkiyKfNKwleae2WTJgBkCgD12I5X40WEexNpsb1tFROULls
u0GZV8lhmC+s4/FeBO3uW+otZguljKjpCmERfNwINhT1x4NZiIIQv1A4cZLw63zjz56kML8U/I9j
lBk7aqYE8HG1YlCf3eb/xM0Bnra2wTLjbPpLSK7at2+w2nCfz4gAISEL5RU5B/hAwL4YCxujHFrC
ioPGpffS0BoOacQue/9lzIKbTfAyM1QRH8KZpz3OWT409o8fVSgxv9/MR6Wu2n74x7wyqG1BiyJk
Tzyn8cxTdpM6cJzkvdeTA7AIm4m5lTkG9G7KfKpGUO2HLmQsILAI8jzHamQKPlE2Fk02rFZdRIQL
Titvq3TwWOUVXFLOTxLP08eb0Brz7Oo5TFMVHdt8Y8RY5tIDcey2zPX7SzjT3LSlVO4NXDeFjV80
7bmb/h/YM+4dFxHYxEEPqKMI23No7tn7Cqbu24uOJvXqGHSdmDgO3PHul0Kps0ZQFsbHwNmy+2aS
z+N6vM/7r3SrdXMIUW5n4NAVkLuKeelVPrsZ0NSsu0bp983g05saEQxCWPkKtxqdQ02P+Iqiwp21
elLTEa+k7+WXRMfU1lSVom8IUInnftxmZw+6TYOgsCUNfwVQ2ntewEFPAO/a8WEZIW7KIa7gEKqH
M++cmRdq12Oe9n0Fj0OEo+HXD34V83yW1h2uKi1V8ZFdSrN27R0mXY8RQ6OCT33rlQ9LVRQGJLz8
PVTOhH52nEK6jafIFSHob0EjCV/9RNbP01jknqgmEBuuosc0sges+PLURVAldYBkgs3xGaDoFmLb
81APaE3/2K1J+RedVDm6Tr+D0gHEI+jwiYDqYzzT3KHm3daFeR8zS+FFHoBKpwVdJaQfkPG+nF85
kzfjz0nXe6hfN1OJFwm3hmnld62bU1nGBpAx+e63T+F4kCnjh1XAK4G0UCShn5LTvbCDuuSAG/rG
c14VA0M4k4CeGLAqTZ0iybhamPJXAr8pJbSqp/SElyINeLv6/PoyCps2RjxdM1RG4i31or8gJOMd
UDjCp+66YUPoK3wkxtomVLuxnEVhlKo8IOyEGCFuKsmfbUkvAKWvs4aC2HR+e8Yw+FNlj9OzljF6
R1f41emQyWAqN4gxiXJA0wsL/3UCc8A8+Y8ZFgAya9k/DM5ggiJMFDVWaVaH8lLoEnvw4TUg4dQt
XPCJmD0LqjucpOkpEab6KIWktjVjPapGmPsFzxDGUcaLHXUFEmeHhnW1Wo0HfLDNwCPurguN9oH1
K8ptQf9iG2Q8nNmIlcUsaghGOlG3/HJhrbh40UBCvgafKD09JjByP+Gzsd3ZMwXrKqgCgJsl0yzG
3NsaaipeDlbyYSnAnWCFzYuzFZKz6fXXvLNFtSbAuZ+7/vtITIN0P82L/xjBjyFnslZYxzTVGeIp
PPrTlA8WeprmSQCee3e4SaoWINUbiLWCKUcNS6pPNv+jrdikjE4cijpSr5dU4HnjYC3MdzNIqstM
Nm7zdjbymNUV5Jw7qv1nL7ApGr5wEiXAdQJO+VorK9DyuY2eePFy0pgMg6HouymO+8RuxmElWYZA
dhv9rvV1QSGePlADqXycT4kI9rovNmaK8q/IQ+F1/kw61yQtbrIKsh/+obMBeAw8YzpigpXcTgkB
fI0ktk6NbEBigs7xnQa3qwHs/v94hLfr0swWGpvIfxKUGQBH66jHhAaxNAzNIp7DsWmNhi8gsuE9
KJ4+e8EOynxOu/BCI3ObajCdAmZcNbeFFRqmkj7k22dj8GtASnumYZ6utq/JB6Em43Zyi+XH8Owr
mfBtiDZBSr2SnN7QeQs0QjPcU+c7kMAgXYRwcaf1Ryc4e4sDSr5dvSgSyeTOfe8+mD37rE6WYRCy
0lR8NvnGAfKTpPepsIdsvOH2is+lIypE+RnHLSla5DqfQDOcjDFaTO7SZq2h/kGaMry4a24M25sc
P1JGEQTedgKEA8iHc+M2Jef4MA+W1Y9EEsw5Qh4xJifwidtwrKpV2FzVb+9An+THYYdJnSvOAmML
PxUvPjmhqaVmVP/59NDBZla5Fq+HC8Xlfj9DKLKre1wPCG0OKxeRrXu9p03p+YqdYWNO1hQIc7Nr
0/VH7XoOab0KwQ4ERW/AnXEHXR+wtiRyTxBotblo9dO4YLtZX1o1ncsHrWT9Fbg185lotNIw+URO
uoW87o2J1DJeMsBDH4D+LWYkHv0APhUNdA4PIqUiGLHy065/2oGKz49ANrggj1s/hGmfO+e/IS9o
2o6WYCistmUb3EIhCDLDL0JOFYTt78MKN3DkAlFJKjvcwGH9G9Gq/RKAa/gPRr5PgK2yUiK+XBuc
C9LTpFTqt3rRHNq4eQSJy4nNMK9a1RAwPqRO2sdriaEBWkWkoZReSDzdA1plURpInEt6yFcbkUgO
Ph0GfqS5+EiisoCPDUhpvsvwNLST2Uns/hMLzo5feH+tTB3L1RimyBtdOh+iCXpZ1ythHqjI5O/X
Epucu0weywKUbd2m/IN+MNYVH2SjlMCZIQrrRLisnoPmhQO7gmWGPEJ+UZ9O2mkxPk9zM0qLn1qe
Qh1OqsoR2QARiRDBtOP3RDdfz7CsHd2c1+co9xgwlx4vUDpD6q0vacnYnN8fHUV8ND/ZfSIp5tR1
6sxqhewxVfa+RcbrzYOSrCB9FmeDJgp/OKIUiwa4JbXezydG+aGXS5ASj8M1WcbLabtcFeCZI7L5
TZXqOF5g/itFNLC9c1aTfVcwh+aqA7ambD1lXFhXD+6a6etF5dSUMD57rINcammJQOKBcCkiQV+s
F8rN5ZmATzPbsuQm1yPUMlgixrdmMyz3b74zm8x99n11BojNIN/LyDLjiHKlRQz9ztRTispwVA6U
xOq1mAGJMj0nDzrmrUQD+qRvh7qWdA5p+GUz+VnRerPHVShXTVkmdGJ1oe51cBk0aB0NyorYDpqb
ZFRW3oq/6UZd7tX87uxyitczonszoP6LkJx0tvC1uC/PBNO0uKQ0Hq7Bt5Mmn7Xk5IJ47gGD9KT5
mmr47B9c2FKCj+ApaFlAJ7CrbHUOe9HLtjzsU50t5aq0va9RCz0yg6+FZB4k7nDSZb+eYOWAsNO/
XV1Qvxgd89Wjy7fAJYw1Jsqr6XmlQWe1t02Nw0nWRX/MLiaEC1ix1N19F1arQhHz82vlagIPxpcL
h/6imqnA6j7Rq2H1BW5h2rfNCYctmDk+Pk8y3yQfDEo+If9Gh397StF3W0EXuB/BEa44K4b/5R79
2oSG/+nPSG6mD8anvyVWrAMC93WWRUKOPd6eas1CXQGV/x5Bj22jbPV6qoTWcbl+FUjsyoTSKo5B
yzxshxLT3wl7AdGH3NbKVKkcRa2zoo78TWJZDRFZlblh1vPgXD0/wVDrI7iBzxsC8CjkIVx9HZ2+
wVhLSTheAgjtfAiADc+i4YIslKJtNE/PpoTCtI1K7OGlkDQ4104buWtKxGbTWCe/u1m3N21ezSP1
lW9AaET3Nr2R9k/36+XSwHF+3nNu7Fz44St6OytFM7lNfZq73BRy8aMOhD0wppNg0B/XCIYHCkhM
HKpKqfwr8JLpveyV6Tn6vzgCn0nooCYb4u7St1MErJhNrdAcoJc2rNPpZpGNT4Z5uQN/RNnu1l8Q
kUukpGJXUqbPmxU0tAtEIwXi81iv/9Rpgk1X8SeTWfTGh27ZwH+8xhAMvysBX0t4EbMqVgLChNNm
4wcqJPa66T2Gh2ApQ9gyyRlFMR7iNTAKRTqZJRB8hKkHVmm3GbVDi96opZLoabU5KcSGLdGsSBts
DGfI56fCd1uJfp7f45i0wAmXEmZxiz9v1KOX1pLMmqyLZz5sIAP8n48Fl7B3u/lkcDBVyAvN46ew
Iveg9cND16dtIhm7Qoo2F3YcPP7GNn/gm9QM8C6HUaQHI6lLwxTP7Qjy7r7ThG8HfcKAH3Ng1PbO
ZLcaeV3fUUKSwJpo5JpGx3qm5wx5ysOcMCawtnUNjlMLIbf2BeKt18pPV6q9okdMJeK3EtBNlUZl
Y2HCxLs/hVugHPDS/WQWkQp3c4yPWisDAAVmhYtDonbRSWuW/so1amv2STIDVK8YQvsN55zfDB6t
IzyQ7z7arzrzphI7HbysfmPBjyJNILHTyMQTg6HOesXgCw4/3E53Q88c0v1z/ZbeOsMF+rfA124i
Pmo7Vu7nnNOsxmrKeJq0WdnIY2Mha15Q5peJBO1CW5Cu5mI3S30/tGMTLkBg3PSYAUMdGdOYWK1j
OeEWhkMS2q7KXjF6/C5H+Zt2fUwaeBl2lkiqft8EqLueGhPfFcwhf3vPpkJhu1D/5krNvgr5N5yy
5OQoLlAQNcQcwnwsB2Rpp7tk7HTztGT8lUVppprqRSBwRnYftLKKNVStnHMjV2YtIBqe1dfkD5oZ
6HemtNxsAoIq494zdEyP4lS6nrKXSZkeqM8Tm3HG8Z1lBtpfHJcy24tWkm2AXd2pJHYa/CrhOAzI
5+cC42kYhlICklc6E7duwCbjgiK09OL5QcuGAUif+3a5NNCbBPb6BoxKS6DkT6oAYedrZgolU6CH
jekgpIqXwhwJWYyM1fsolU8FSR4cs9292b8Z6C3i1C5vjWMDjVxv12EvuFOaX8EQHTp9MVa4CX9u
bAGpa3PzUJLoSSsGKAHVhiLRvdtbsAMPf+8PZLmSGcX/MQbYtNxdGMwy9HQBgmup/edcq2ITFm17
AvV5UUWRq4R1CvRc12rlkXCTtzq7Vo4JgT3VJuDd0qcu4tldor42YRWDaDP4tE9W5HfaY7a05yzd
OrySvEEQhLP+wZk03jyEfsUTeNSlfzDKk+Ix11FhLN/FkiaZpZlhdU3c8jRF9OvkT4vcfMj52yiu
OLMrUP3fFRVvaL10+gMmkjJKzJQzkyZDoQC6U2TV17uOBYfQsjuPdtMApmohEBD+6xCj0F8rO1X9
dzgBcexQPKt8QOYFraAyUy1o3T7lkct+Y7Hpgw1MlNZGHFDHYvFwBqMAXAoapuqRSGPldAqZOJrE
IwvuQjjF4wprXWuX7oytxIRQc6W+97qQ6YaYoPB+nbRa5tTTgzWEBkmZikKRDBOVbRSXmm6H/fJy
y1a6763T0BsvtktewJqH0B0QNjp/uZKsRjFrIx0EdLFOuVlJ24u6NWZidCwojXa6VXEP6Dve5xRc
S12j6xktYb+L1qepDkTUgdbx+JI+R2qYnR0QeY6zF7MffZN9JYNadO3USQhpntW2Xmxs55Dswucl
jbQipk11z1e8u9d89F4aCMKOSrxrHLsYOFW/E+9BIofyNFSI9EqiQRi0vx+5NjqeJs1qLHkzYfzV
U3J02YsYRHwQrBOzQnxTDoJvQBq6fHcADeDerdgrkuEwkuHIC0y9Kwo6VEG/Y2Pw+aTE68Hy6KiQ
HTahvFy1axfA7hf0WlN+lmlZ63zq3qP6tvZ8THS5tmXpcYFSXgh+ZvEXeyALMLY5t+3ltArrXyeN
+LfR/VMfQlfIQRASVAfFbzLyCbyHE/AN/oK44oq9AO+NsJcXJh2p2tmT4ZI6+BcdBqvibH9f6A+H
KGNgmN2wixPOS4yBAnVMldzagbB1kUGs4e1iCA1wUP4n+mu3qtN0REWgadiVxY5+AClMeWEQjxXq
HtkfouN2Ic3mX1cHPvv+O7PaOAMtOp7O8BP6oQFq8LRo05Q05VWxA7J3zlLsir4l/p3bph5pn+Mq
JTwxkFYJpYKctamnM28bxoUZgdUHuMhHqqpzRVzixCCwKrF3qruS6ilCn5ScfTcfspfwyd+Uf44J
xIdJzG1fBeZAuvaapUso0mFo4K8PnSyxJaGQ3LpXgWfI+P8BvGTrcEoySfvopeYgwQ8/4L8I4P/g
w04Dx4+179qb2MguqzL+vTCis+CCQIoD6DD73OcdAgih6UDuQrh7w0P0M2whhEHLA56F0TTz++x6
nt2Hmkazc90pvYNALfztvJ0FlrL605LjWYWryKmsT5DUVKywuH0GbsD0dd5U5MH2imUsu1ieJoVD
QoULXzGRL8zCfs9TpiKu8XE0+dows8nMtjeE9CKle3k9ttDVZKf1H13wTlFo1I66A8TdBz3gcioR
tX5Xw8reZwfBOoeScW4syDUcrkNRHa7bfWvmiQ3HXInBxrnz7cmP0ehzxYFzTc44Xcl5jg7sSYSz
dxMjSsRYzYRA2M5ANZnNgoCru9oXpRS7k7Tk5ib7DnoFHAlpHIdXFHNdqo3LTvOJmbWdgrwcJeR4
e7L6qNgw1lzO0LrVfo8DysCAO2JjtBwxRtnZ4gKBxcNWjgXoEphTp1chL1oankE7vcWGYyFpaw0A
vI2gwYbVZzyTwGFwGIWrxMZwdgH+sN7KYyHtReYzP406Bu0qdIBqBxhz2nXCc9SQdrbQQsYLM8D+
UQ61nUWkTtMl6MYmnNdgd8S5+w8B9o3weVOhgd/vZDTMkSeaqbTOAOYT0A/xYo1YWc8kKw3sKqvk
FYfLh8EEuQ2BmwLFxOab+sx4LS+ZGYi+ENcIPX1AU3t2rbv4lO2VBU2b/ptoAJgWGoYRfGYuuW5J
/gbILbvU1gzmpbAigwiVJnprqGlzzxZ3dpM00QqTx5KyPkh2xlTWYvre/EyQzg8Yxt01WaI4vp+C
mRWMRp6ixvfu4Mp/MUGie4u4kyhgpcRnSYVn6erNmkOLmrxqi9fWUWmLo9StStjHOakwS2ewchtl
B4Vu7laiWAUZknrkjxyKGMQB82fxTSuMTjUPESLcIsuysp/dv/Y1tqD5aQqzOeYEzEFQcmRFcsAj
VBfEG05QjCDs7TxR087WvtU+uWHLSgXNxhwaFxPr/3KlKY0hdluXetVpR6c13Sx+UCTCzV7SsKZJ
c0I9w8UajR9ZAX+sx5ptUrIAFOc4vkxN9njUPCIXXE4m+fvhrkH+g56Uk0XUik+GByoWsucNX6O2
mYU17kNBzocbVKqhxai4Oli9satq3agqf7mYIBQ1uePlkqITPOZScxxGuIKZQYNz85Pj+aHuItBa
VQjgS5hLnj1YeX1CLtw7vecv6Snvq0LVGgAJ5r/BClXFd/+1zjpYNtfmiPjCVWVMlkBkflVi0iez
8gy+ZrDtQItldgfEpokcrkY6nOqbCCGlQX3BBhTon3ZaouL2LvKBFbmSUGlkBR7LerG6XrRM8hvc
46dPSdqiPMaczTLu19rIp68r15ho8eOI6aC703PYmMwJ3FylR4S5+KH24k6jZ7cVhZmz2mURxfZz
gQ8cKGydd7ab8q0DeqxklvIXMcvsbJJSwbQ/TV0+YFwzwsWJGmscIMr4cnz0qtFAOqhZZFetXAOs
Q9ICoqiul7e4VloDWximjhjxHCFuh6dQ0j55LJ9VhUC1J27k0yrSe7Hj/N6grFgo7TNTq+48LgN2
/3MBAbvmCpxMNbLcTM7mihdIRRzv0khodEckb+YyAlQ2Nl7Y0Gsa3WBO+fa8E8dHD18cKje8Bo8c
KYT10Qgac3U57UefEvRg/lWkZa+OHYHCgSNZf7GHW4cLQfmla98AUdwAua+16NULqxbxcLPhorGg
mta6ZJV8DnztZHFcXRU1STBnwYR0eRn6Wax44x1Ymsi1JZ0cpHTESyeuBOQkQt+6LlJRMDS2mUhW
tWhY8n5AshTAaf3FQB6Tty4tn5SfLWI2pneTRRm4NWTTB1tUuKKhmWvCTs4RXEXy70lmCk2LfJv8
t+huQblgu0G82328pqnqXPgkGYMYedL46T0oYPJc1GUJKuwTxboR37wsfDlLDdK+A9MmH4UeceNC
QjlXjNGUxTnBoCwRVABr+NsavwfbPtzTuzOzFu12poHXCTDvbNXy89V0bF+KwVa7aaGJtNVDhULy
QOP2FatpCDEnxw5dF5D8h8/ji1h+sLk6rV/pd23YednAyvh5za5xg6vW9HKXEitpWLDa2eefUU7b
G3zzjSO6LqOXZzRKSA4baqVZ+k8R76mo89SYg3245ODSqZfpnHJcm2zM4P2lZ5vBeBPymYAno6A+
uT2WcSZNifV6lXmkfcJyJeTUpqCbI5IXCFrInNPOL1K0Rf+I7Ib201d89XPhKFtgYTRt1kGObmEn
XABOTlun6RY3MKphz8yOepvCb7DSzV2zq+w3r/hHyFiYVA0qd91jAxh/QdISL8Axnjci4iI0uKGJ
dCqS+L0QFqIuGHxy005RcCm8R1Ml4mNsSpz9qmgAbmMdi3ARuSiUhfNK/RsubSVyJE1pmVYJKyR0
y6z9IsHNbAZ6C2jlQ8eQWsd9GymTZlAIsWbMKKfWLI4QqBRIl+0I7AReGd3iwyX2gZWTKzF7WW+F
kGdAZ+AZAmiD0kdefMAF9zFdSUt9OpsE4M+ELo74SDZkhxtoLOWJdgVpgkwNUJUrvyzWuxOM4AXk
9TZvCFbShNqlcSq3bNIvwvpCy6178ZC3n9/hCp1shI95LmvReEYXBNPpaV3k95GtNSyf0HhZ32gc
RZLajGCPZno0RWuIDiz5PBP7hmILgjqaSyydsMVtFKktpXd4a7RlKG82iPWZXcCmiRzblNp+Pw0S
LhTQibOjaQS0ElJttg1/DbFVjidP64u1Px7WAnCkyfzALnTja/Q1KKarVG5iEHURoYQMkj9SiOmD
b65PiNR1GZHRVlWMowbZpbs+p6OCMJXoflC5YtRj0vNzoxwaRKrGLgtekp19bhcVXuyd3C8W0p0J
Ty/MKH45BmU26XPfWQfCJxW+ZRVyfZ4p2D18p+yUutJBSb0HaPqok9n0YWmcsnqrBVPPmc1g58IJ
d4pe/i7w6x94YMh8aS9jY9eRK5UQaGa5Im+jMAWSN6V82xwn4z+0fteiCJskyTqEWvqyaGZyLE1r
OKL9C1cypIhKA6LuWHTUQWD3wqKXyesVcCU56WREb6WQ46gqNuPQYfpGr07l4UPWOoi2pSquVr2Y
jXCvtOxqS0JLi6a8beGFawlHtHdnwFGPL0hE3gXbs7+di6xEho2j6oe319dC9MYg3kn3j5c/usDn
vmO2sBV6KBFwq7tXAT7mxL6APWN17EYB0OojFU/YWEvjx1nYp2dX+wD8sQfu0IoPtFCG3VNP8PZ3
SMUsmXCcIipsnqnmPzOQyOw23cm0affcwW5j9YmHmbg1FmUwfDPHwitqS2V+003eUHEjzDKqdAQ2
DtQT/4UaufClRp+4HQIQRLsbRtH5wcYfmUKxX/hzUSl5bUiMs1KfPJVFRjrUOcppj0jxHTPNMF4X
kjnrrWE2Vns2yX9Yf51bAUa8Ec0JTBald9SjF5big0N0dovi7dL3xF65LTDivJh7Fez8h2s6x8dz
005B8NeDa8CmL1T0aX3+E53IRGUz6TdxqneCtGxkcZ0A7Wtrg7iuzPBQPXV9tAPMCynpZrPoY63y
lw66OC6KVhrfCApFIj4h9dnr462N2rUUq11kz0IDe91NAXkhDSfq1KcxYOhK7ikXfY0OYIaqZpgV
LSaZY7poTKYeZtewqvjqkAblTC0qILW3gg7YJvEso4bLpx/xEzliK2AWbDgTVQzDGJarotYfvPLS
Dk282cTFfAMFFENNanCmk58lAAzwI0dx2J09hBrgwRjFgqoNqZQTM31oip8ZPJ2+VE5/FEGQUQ1H
APUxxYGH09lc0GKIwgiw5UwxyRw7K7y4pVygkLrlF1Ksx0QOvIYnF3hmZxtkTIc4DQCAwQd15/nP
M96SF0xIRUqn1ysPomOmQxNup+/TVuFE8zudiIhdi5HFwc4vCn4W+eq7lRG/xELWb5sBvX5wXgeQ
rPUlPZikG1puIBpPv3V/JfLzV12vGYf5C/WAL4w7LYDBhUdYQ7K/OUCPyAZJ+7TapTGYjuWJK0n4
dR6To7RIBaDNSwsR0xlS8pVuS/GAy/KrX14yIaCtPrMhWVZMoSmpwFswdwiBE0Zue2a65gKbxlgv
ehibJHOvXLpX2UGEXhp53IY/axBB0TkBi50yugg3TP1qq5y+/Nk7ThOdxu797I7lpP8ewMdu60Po
B0EEeZCyJGnQbgQrAtvn1ia+r/MLtQcMX6mppCeo/T+gwC5k6KmPZcwqisLHFXYjujRAZ9aHfriu
/2QPnCuRss5vC+yiHtKB5NtkWGuJr8B7oY//sxZKN8qUNN9Wuwkfbqhp1qMXKfB0IFKaRH5D5XS7
DCuAKzlYR4DnaVXlrbzTYhX4LveIhBqAgGieQrgvpToS5Tw1TeHABTd8jMDHyKDLcO7Ho9rUqfX1
eMJBm11scmH/56Kxa4Gu3SGKRbUy43tjAJgUMMbpwFv131eULzC9pqHHYDuRU4gKS1oAiOfk5r7n
FqFUx6Ku4mjNBOxrayggQ2YD9T+A/JUANw7qdDpqFqP2nTVXwMunXuw3wl9JuhS526mRFI2Sw0Tj
enOPNSJGLnpm5BnRCBITdWkpTWbR3nZt4X75rf/gRvcgqLB/ETKfbYWw5N9nBtGbOEjjMBYLx8gg
GA1PeZ49Dl4TS0H1YgHzW7sEJau9vtyClJK5msHcxWF0EMNE4ivOJRaB6MavyijDYihqbdxCNij0
02Mr1eOW4R+Y8ZLHW/Pqh2cro3zaC6vxk6qy6TpBKL+ues7wlTHXSC69mo3OPOXqdcG8U7CMHhcy
nqca6CxNp9wBnxy/vOFdGf/T7//sBYTk4dB/1/ytMPNNZDkeaiMLblDhYE7zPotUxxOLE+b/dLIP
anWhgZBMThAAxPZJNOfQxpqDVtq21Xg4MWhnZeZruT+jMaE9trsFMKPWALW/STb4rvwTxbPB4hdK
1ejHYTiWCyn2LOgq7j8j1FZ8WNeYE1wZ4QYw7hkJt0T/H8rrNFhGu1IYTK3OpZtSqrfvgR4ISHNY
esa13lyRKEZlMq+rsJQLrCzo3ZupAOrWSV5sdSCAkTH/ZunZcYKhEmExpIhDm6b6guWK5KGNK7Jo
IQUCc+dukDagUuYZXNjxLdEZYRZ6FVCGgjc+kuhFta0fg0R8cdxBj24tiOiasKGb9+zfQAil04lO
6IXM6mkzPw9X08lbfeVlM+TPGmS/7z9tyNdMsAARA5yKCkELFq3Rc67WYWrNgmk/KDWdcYHleJHW
7tAQ+uSntQrwxBAjBmbcl8QxBR+4+al6wq8YmuNCzXtksm5nUyszUKYAMBxR2qbBYaOjP7cEOVlE
qiF7N4Dpx9hnbxc/6TO2uipELy+/HrwzRg8KTYuSHGsuTSL+YcBiTauUPCA/17NEXy3nMS2M9O4o
Ye29t7Ge5NkxdFJjrgS05c89jqUprj5ff5VfxXyuq5AqD7UmyyS8dHp6yl45WV9hSP4py/i0sk+p
rlHCB1ga2mgD4ka5l0qb6ok3WApcskkjU17wOatcdfyOGd08dwr/PdeRWmKq4uQBkipmFQODyOoL
RKx4OCfhscJWV4aNYOGB00o0zXY5xsvbh6qx0Y9wi7t6hpijAIqTyitCzV6J4wpP3sDnAFviZR4k
JrbjyKVkL9konMHDmvMgQJkuDg5aBhYiJgxM2sFCCp1CATPd5IIndKY/biQlNDYg8j4lyW39+P9K
XQ50bM+9CoFSxVHtBPCwCfIkOaydY56PZZTozMojYO3rNmdU2B1DjmGHREBTZDhx1qWocEu6g9x4
QfiAQnMHp1Brz9i4PsNCBXijhj5wKPkkKmuuqAXqaaCozsv4Tj0uuVopXVveRYfaVMJ5GKqZmT7Z
TFLFgp5LzUnkj8A6a+4xALKbGBZfqgm0LRPM5O8Y5Wpi+YDo19DJAxnvprGvpXNQRfBShUI/KKDA
qapK5s2rFu8bpQG0Q7+nsNDj/vd/q0Y+ZxY+6NdiZn1zz3FPFCVL2BK0PvaGBSnLkGRJgEcyWTjj
RbA8ZaAXUcRhj3y3MXVFJftZYSk1ESPzxMsqj0i//f3tRDyMPOyxqlvynyOMsEtLis9r2Osv780b
IT2f1QCsbl+2tTQO9T77fCOJZ5Yf7t/vN3KNSYaJVcxwjdDGUH9SzXwyOCZQYou498MYN7fW7uCF
mC0Y5eciZ07AyAK3hwh39mUDbGDpjjCnRDUoFFkTQ8pTF7lp7L2fKabih4nmo0bcyQh+rP+yDflO
EFukGsi+pcIVgUV5OPfaA45ppyJ1nDM9aLRUsn+5hqokUJuQHLWZznThCNlBicOFdNRj6XnOlkLY
h9cQjkK5CD0ymz+xtzp0tSmA2rdZ6Jp2hXMskkeVej9Yc1JwTSCpkZ239/UJSMoFIDqz0ZdL1aZq
4zVYMwFv6PF4Mgi8WSxU5T3EOIQ9drLA8DOyS2Gvj+N1hBmnaUQH0gwDaD25FKjOrAaylI6uSFCU
e3q2vic8bhlRVG9QbnxiMLja1XigQas6VpY4ChNgzOjMskGuVaCKayTuIyhkIruSuEHUdb1Vnnyk
8Q5qqaYHqXY/kiyc/KT774gbvZfXnL9oUQZyfmMeS19Kkuu525qEcWVJ8PBEQgGMzvrlYsq7AT/x
Kf4Iy7owYBmJ6PzamCUOiDO6hE5RADEMyGeRJblxzEjDyjRbU+y6xbpHutMcjWirj1MVr8I67sEy
1eLtVZd+bM59FCCB8ehEr8a9BDVjknkYSUZFtmox4uQLM17VXh0twV36azWAY9dMzGv2kkpyBSqf
zROdMbJwj5WypfWqCbm1joocgssSS69FPhhkPHs2VsWA7BbteC9QPJ22zeE6+Jc/E5L3+GGPTEKh
tft+c41LTNYqVdF9fE/147xHEtmnK3D5T+NUVY8mTBEGlrjgo0hqhGhBdu7fHklA78MHr0/epon5
btK7U4+fjGPi41rQWlp4tQoP0aKjD3u6IO+Y9ieVz9px2tDHIWFXWbg/vfroSUFWqc3ZkMHRcK4K
6ixZiHoxM1Dz+nzlgG4SoMOHHm4RJJ2pPddfGEtWL/S7XFuRwkN5rVXG5jIBJPobVdW6lhJbFt7S
bYH9NP+3dxZE0SVsItk0wbnDQX++/N6vYf2vjjomRZzBlvI1ntQjt6+ARj8I8PhMTGm4O/mykoiN
VQURoSikJ7THddY7PghH08PJlvl32NASnyQv2s9/2rWYC0CvoZ7YNq6rX9CJgKMMtznaEzPWHBrn
qo0VAcvSRVwam+c+N4RiG78BD4g6g9rKn0RPPIYijI8GfOZ/gf5k/kTG3WVsSwEWCT+ZMipbtS8l
w8EBkM5eBiDWu/5WZPuE+7LsetBBL978n4+VaBxjLjSCy3lzVN1BE5tHMG5vDRrhbqCvR+JDVvpL
GeJJSWuj1eCs/xav4RIdGebLbNuLUiQHuL0v5D1H22rOGqWQaOLDUeIwrnjktrqHrpkPo4+Z5ETw
p8T7AuvD6CeNbVQfEbAe1tJxBZwvgXe3T24qvLpt3BLTpYql0ctAb3WqaYCE5DuMZg6b27R9B07f
QK0Jv8wqPEiDfw4+PEuJsjNN484wwAnshVnwHwAp9pOkreF5qpFj8ud1mBHJGojrmtKBDCcbnLIF
Ne67ut4y7yb5Dp408lbUzACHsFtrSRW1/vyc9YDyn2/Sh0Kyfn3GNXXeSL31sPXBibzWoZS7LhMU
MX/Vp2lIR2l2IlrdjB6Nn7+1kWFWaeoTt7ApH8Nvy6UK1EoCDQzs4JtHo3WmmI39t72ptNynn+N+
GVr+fAowsLbEX55QguCO/Ts9trB69KHC+ThhHA3DU0ur0yPHCwa6n9B5EP7w0CfNiel+pi/yqswN
LR/EOj0zxhNH9LzCzD6bYfdT5R7GPEIMZ5hRt1vS4kDDTnz4qMl5cdWSHH57FQr60Dscx0Z+F8gh
yqhbFUI1q+4rZE4ojWj0bqKeTCmLROCOxPEkIje1Rzaia2tmyfAZFFR31oeC9aowhYs5nqpCIIKy
I8kIR+F73jqNFUJh6w2jLY9ZtbBFPEUZh3Z74N45YQZYxnpsb4iXtUMNoRf0jXoHTNkm0kSm3Phz
R3KZ2TrERH/VJ1GkHdf9MlSlyMdBksfrO6JOJ1gVwULPAH0aYtklIyb32Q3o72FwI+V7zqj60nBS
L0Zx+f4GUK1DLAlwY20it55fN0jdL9WdPjmTRCpVV6n5dDpGocjmbzKdhO/zMnHWUiNs5N10DdAi
j72HUNy8NkfPzs99K/xTBcdwJAu8RgMbweCjbl6jF8Jk33ZH5gjsKQxVq4nQ3Y0+w1DeAfFIappX
c91UltpCPGe/6gc6CsYJplEze0UKeO9JQm28SiiyaIP6pQYM52SyoZpXLvV0PYh3S6Ir++6zJV+s
qrSWZtdDjoObyAhb6DhNzzAYafL3CdkfEdDagCHQqLRyaABmQ7VtDbrLchBIKOKhSY5O63MCdauw
O7uR/SzhG2zrD7wwpZ3FVN3y7gZ56JObDZDAogfAgiBr3z8t6Knkb9voQAWOzPVNQPFUXfsZMt5q
BFQufuCC2h93zc8CJs9bx3ic01kmTofExgSoTEIs3spkQ32SExPetkvn2OnLOYpVImmBIasIVMeD
z01EVZ+dkROldgy/H3gZqPgtsPJjjtoa6Ar/kjQpSSJrnV2Bxupubn7mtOiH39A04FgDtmriAvFz
zoIVXeLKEJH5epCQr0NuwqczvGuiid6P8O98AjUVgIDQI1dHhmKCi1bjfFyYGCUsSdYy/5geH+nn
N9MekR0ZnODBUSW23d/Er7PbhLbtN1BWayNFqsaqPUwtBO+5hgQ0EJxj3D/v3Mtfr/DUSIbHFUdk
wyOZzN3SuNcAeppj0LnN6Ak8T09KpPW9d+AYjLqEsFfij1U1zEcqinRhdN+joJFy1Q1Pgy2w6umD
HHFs/O6TF65Q0Wf8tMlyMUsziRql4R4YSQwXqCpx9HvR8BpVjM1LT2LGMXb7QEvRgLhxrR81heLW
tgY2oJfAZLMrlfWvvh5pDlTM15gdH5ICgtHcPKfMiAh6Qk9nmkwQzXXpkcpxa4X8zSk2wX/6vVHR
gfI79Vhqw6g5cufrgzNVogN3wpPDPoOlhRHkgDuUdBZ0FS0rZvnnKpwPPIZ53XTTav5HiPkRphJJ
vb/Pzdg/FisqiZgk9IvXgYTioKYNUxLDodCQ/vWyykNA0/786vaboKWzuuNNpv0MtqZ1k71VZbiZ
ChKITDjx+/hS0n2mzbN10kwbCz1lY+ZHyeo9FM0HDf0TWQ3qLEUtbYJVGkOWrAqF0nd29uWXxQq/
h3PaZI5FLjfM5suz86nZ0DkxAyktdZ+vGle+VFThyncdEop7pQAVAKUfuVNrVNv3a7OI8r6fJdiU
hFFXyb9x15L/FIVllIF+Iq+FNe7P87irDjyOPHArTid1jXYuUACoZaqvn2UTcDqEWZmHAOYt9Z68
Hm7wr06Kw6aVN5RMA4fZjO+A08shXwcdedLwdqQMzJVGM3vDpw9ztuWJ/uw4b2DFA+nN+KHnhkGr
DntPS8VJTITA9j6q0xJsWRaZJ1tm3ywcwRlg1VzO7q1mKIwgHYqZUBktVFjh5JiUC6o2J6wc5oUy
GvZ+WOiGVb2MAub4lh8F4L3K7WerSaQoIz32qBb1QzzgsBiDNNhLEL+CvKuVt/objoGNG+c2zR/3
n4hoyMznKcwN6vBrHhVQyzYStBWHSUdtVcRSZMYtoAwseLM+AL/97100llcx4rU7Oy3Unvxa7ZKn
Z6R8a3WwEdoeqK4gj/6lPSZcIhL24bO2CZdD+nIecbiujk0rKJbBXIEzwfY8NFTJB7taJVW2hfho
NS4FdiEKviyj6FgQur9wTURwWeNuyCVnkLaFW7R2oyaCi8TI2PcWw+yJfUcN+rkwBM6YyfePq98Y
yDYLZgrViBkXxGmJ2Mu6Pak0shYs5qLjVBNItPPyH7o4kb/Ta7r+0sKId4iBG4uf6/4ZJElGuvA9
4n23z4h07BCxYqHD+y0vPs09LMhCEMS4nJzBRxT3VIa+1vQvFk5zmvMPsvsCpyL24tM5r41mx2R2
SULWW2VOEsYeDtRR9z+wcbXYkIsI2MOyKbuxod2GncA0BPpOGJCeNVr66sBpNNWAiURBVl0Ey5VG
RSqI15GZm5Dx+phm9jnbMaFy6YejjW6qz9NwDD2Q6WKC5ZHumBkCONSzrqOsr7mV6SoE1g1X/pUy
MAuEWs8REE5hOQyYP97zOjv9mrNq1sc0Ilawwspxm3m9nKX1GETWdo5uY3RRkA7u2gxEukbxk9E9
pBj4eGXBx0QqhY/u1DB+T2DW5JUxYnd+HlTYYbSaQMmcJ3CoZmeAiHNR1iTv63IVeic7Oef+xP0M
Lg7SLht6OM2fhHh7+2wbeZSKn4n8IZm1u+yt/03+9bkRUWY26pqzMl6d6bUyLFas63nDAJvTahot
SIheKezS+3gJKE/rlzSspvDKCW6cd48dWaguhdnDmbN10SEe1nnfpFAnOHrniZ5DeYbj+PCGuadZ
aG/p3RliAHHcSt+HGnlH4yTUjvJDy1kpRHfiJOB80OZ3Ta4heIyh9rCl+nUwA7K6/ZicPYPkwkhx
hYhGc8lgg7r1BvEHSNHv3IrNiQKGsLcAwz/ocd3ZPPW/zSwzIZ7VlTr+vKogWC1pGH9zPJLboqI+
F6W1qo+KxVWNC2TEK69jrikAWW11QQsMdXiznCtzwGQBiBUYGHRQZZWgKhRb8lRmJWAFoKRz94kE
ZCpa0Gcjcy40B0ujVY3iW66iU00EjquE/shZAKLKQBfYRue5NmRXgGJX73azMaFj+iart8++YGCH
qhR1EMhlQ/xOMgxZMble3qIIqTWXEo80bWJ0EO1pk1nfpNviebpcpjQHbcMTz+zoakDQ7hxJBdxx
9fKiDAiLOViYHKWDZAX6EAbi6LwbFpYDlnhzlS+JFD6jIWY59kDWdDBXlOFRAupoT7Tw67TyTn4O
WLd0Si3ZZqmrIpfWr2rao020itkCn05qOoJbqZ4BLh+ACCq0nRgp0A3lBfi+H7SVAKNOt35Jv0rk
uYR5TsPnpydcOWODpj/UYb7mScf0oY3Q1StQjtzsE7QmMPw4Is8ZSA0NFJEj+nWtM7Ik9csXoM+m
LuHQ3oKGxCYYaUROxg3Wdw3GoPpUGbxrLlCEPDRpxSMv7IcYVmsDl6Rzk/o3jugpXN25Yf7QXV7E
kAcezJaJJQt58ScpNq9VgoE6YjM2tVNurEFHcL2PMEN5PmpoPmACPcVlTPXvXnx3H7v2GQMuFe78
d79El+LVPWbj7crHiJLyngb95t/tRC/6CH3sLdc1U/tT2tlkX9an/m+1BturMKI0DdKuZ/Gct3Vu
RMcR6TZPVYnXHtRh63X+y+isiHTX2Mz2wG8F0Jxa/rEG4FxfB9s/UDIH00/t6Gp2SXhlSJZ2yj3Z
ufo3mbJkipfRXtZ1y2L4GvAudBxBEbL4Ke4nx+Z8ecWIOfDzVsgrVxzscG5eJeibKiRDu2EZMMv4
cwTiIcbRZADT1rHMi3LT3ZG2hPppL62a9DIgqXYZnR6HWPkNUiQioXQE8gTCrNwWfRPJG8U3edif
Jp2DomF/cFJPA/nV77+a3YlMw6a1pULA7lAPPy/NzU0bKS4iYzvLyg+3F2pGg66O7eB1chtljUDr
YBB0Kllum8t5p/Ia+GK7ini3efjCkRZ1H7uOlrfzuBHH4A11l3qV+GfX8/LEU7/3aa96ebtmTjF9
xsRt0jw5iVkT3epw5pCx+NGAPUvlPA7JVp3pTy7vg7QTmM1Vdg9aYiXJk3J4gYCxTQq7hyXRIjwn
RA5o4dxVw+O1muMW8Sb7vPwAFlGaqN/eDWm+3LacmuFuG2x/GXu5+o9ueEwjfX2Oi6sT0qXpYc07
RnJMKb/w/8pKb1OzBGjyMdyP/DUbMjRH39MmXByFXcg7zQRZbVIaYIWrYEqMUh+xCjXD1IW7QkZt
axzUfxXWM1NMTbTpZFkPZtRitv+PqpfssXgoqSgyUrZH8TXTQjhhp1YLobdlJQhxwF6UeN1KIIEy
U7pIH9kF2eaunCxiiXG16Cq6lo4YB2mxz7Noegvjjkb6szwnYDOOrkCwi97OOstrxWmaPhbnKceU
aPMfK4r433O4aKzP7/DG5GOzrT1+M+klQZecf/IY+sMTlLjvfSTsAWQdqB/WoJBbvUDkjyNvUzTY
IC2O3Jh2/lG2UHZTNzxXbQTcwVJPy1aezalf1wC7dzEfU2dR5mXwzpq1LIIvbfWUwSurCvv440la
1QsXC5UvgPM2Q6NRJE6sSqMxwG7Jb9jyKA5cJHrF6UM1Oc6TAwP/a9WTq0lipZqS9ZDnrXBpY02h
pGhwYKbdyOO9Oa0PwcZgJj0CuabIU1g2cmhGIBoFpQK9jGNy7qHurtMkFOqrhCTNhVxd1JhvZCn8
Af0kPuD3hu+sfvVfZ4X92FyPnEdcsjhnde52PSKpak3wtY9yp+vZBfVl6QQr0d+l9A3z+6Z30sCj
gH5wsrMtvNPZIVLc3PiK8tHH8T7jkbITwzJUQkvzhi4xfk2/oRu3kP1ga9zRMiFBVszSW53NLzML
HpZbW1vSTIPe5t28gFsxhUvDmSqtSrUoo/yp+Edl9hLUt/AxTaOt4nDz9CP+KfuGpbI3qTZx5v+p
AjH51ad9Vh5Vy2jNSXSXSZbkmUq7iEHXdp812Wg+/XPVCW9murKbt81Hn4wDcFgrvurDZCEZCbxa
cPv5qkiGOMBzRMZ7ICUeQJum1DQOeRI6w8fLvImYeCEonGp79plew5JLydpjYHzc3iAODaDr6yeL
BW2SXA047gXqpMd1GL0m5bY65OZiOUddv5nrDhyyu6kfzm8ADXRprVZogpif0ufDnYj4bWRIPhug
dTUdhbvgPK093Cak6OeqDxXZWkVhphr9nB8eMDUU7ZsCgMnI0Vl0tIoSD9Amxd4Lwzn1ytQRYPX6
wrBVn0SKoWCx1NamVP6+O7vfhok32kxDQ1qfyRZOixLY/WK+h3fi04NPApxtKTLRLi9KVuWxkk8M
XRGXu5U4pB71eMvY3Hr27Aq0aH+K2Nr3BGwbrEhjEjlDQ1+7fzfxWRJJ8tan0EnVwtxR8P0qBWQ0
tG8sTmuY+r/PQNXtiAoiWAq9g3RbdZ58IyfILKxdtZbjJoKT4l1DimW7lZGDtjsIdTebPGAl2noI
SwISgtqN69MSLMlshdA9xShk/Jwhxqtdpv7WFZg6YqAH3scX2KQW5mctb7Xg/hNRxm4iXvPHTlru
QTDpEnTPVSRM8L3PfJ4CoCMNstLt6GkfVQ5eEl8Ii3sWJGz5iKur9S+5rwd7IW4MZXPRyMMAljbm
/iqAPiGOOTANMwcbq0Mcq/3+2ESZXW8htTbwwYKckHYCJVwtu32+Bguw/RuRW5H7vI0clHjWuBO6
D+b4h7bHxvb45x60Ryu8SMuSdEDsAZFU64L+tWkOtnfbXvN9JTVytKRLmxmrKTfKUq06SWzNjjTW
fo5cWntrZKuppHEGnKbiTvPvMUMzWSgxjcRRXGh5N00epgVVwTwyEE47dZjyStbGSPImxLSNP8tg
zS7JKfheAaYjDEGU4pTzCrvXowp1EhJg/aOKDSFi3beSgwt5Uf7AXu6a+KTEZs+xUzsCyYd3jabJ
c0BdARKwXD2evUn+NdqhKWqxm1pka9MD6nUNtJWlqPHyyuADEsu+/xD4cmTz3nG8w4yRXNhHrUL3
Xm+yk/7m7NQKAEhhjqM0lSVrizdF5ORS3aU9CTUJviGiNp+rJONkDQ/8aaQXgL+jHCaPrNPWl5di
Fw8d1ZRpcAnQEeef3MiyOFuzcw9AzcX9WhfFod/F2WgdhnaqKmCvFA5zUaW8DacluoKL2xx64YwX
cdnbPCwBMebx4mo4Ne30VTkpcob4xBk/1/pe/v9RfvikMYGRSrifgRIxv1tySmg+4h/AXph5d9oK
kBSnIs2nrHRpWAx8yT2i9yABoyGvMAqQsGWY7zTN5Rxx39Em8nvHfg2PjmpCl0o63xo2sLWed7RV
qNL9N161/tiDAc2s7fT70OVS2Cxa8PFDksPTH2sPH9NpM2/TY+AhlnfVbrcI9wtwlbonO2e89/lT
/3I3UxEijpt4yCJ9Ws/JsQCPAd5VunpPko+W0xo7agsMpDdiZH8Pf0+ayztV7Iy9Jeg7XoeLS0BZ
O5N9Jrgfmby8qHo8mf9foJQRrDnTiHyzikL8Kh3E3vpZf2CVyOfzItkmeIMsEDOFwOY5FSQ8L7DJ
PsxReubAworJv382w6YzBDBLeaO2BPKxOkdfa38RBXzPK73rlNkTzCFs2GF/cnp6uSrEsM2yDQRT
1m7pdF91bsSAbmYxWaMcLQVqSh1Cih0g+sS/RCeB6+igSIC4UcfdqHWJvOqrxFX3yRRo4Szw7jv7
YKuxMHiHpOsDprYmO+zirQ7RXYGRj0z8SA3C9kXC2nUALNG45YVdmIx8k/PCcsfbK4w8fXThjOm9
FjGZBYmOnJj5tol/2HHAv5qm58ufFvA3IKZJFBCNemURxJ98OrsZLHExSzMngjwG6lyLuu7e5Pwt
04G1x+XXyQmpTW9CSeHh4TE+bJgD3nvvw42KxdvS5EsP9I6MTDiTY9ji43TcUeiXiXt6H/IOPWBR
tStuKz37VuZkfNocebt7NjXzVKwsqJj9RgUoDiRjbwqkHadNjV3ZTwjScDJlL9jVlN6OqppDRURF
tOrK0gtaHPxGcfAr2mYXTsc2XvNw9k1te5eC3yVQKmtle9UWeChyp8CIKnhmRrlVhb4qNBtMfBQY
gNnCDE4cs6+HGyzAgXoPvzvl6GwFhiUvHgAJCDR66fTyi/q4u9aZXQtsZFWaLhreApooPS1pxCEO
q8N9+PLP7p0Mv2nX2ph04G7MIh0Rt1b6I9J75deIVOMHLwolJda/6ykF0Q4FdskPNYjMpPTvoPd1
1c5D5GpqvdosSEwqI/KRj+2zNX9Ay+hbscTuqhhe2Ncp64B07KZc0zXYWNAAeStcw3WWlQW84vl2
7qWKd6D/VYBOxGqIa/R9a3jj57o1bQjxBrNvfQ1lGt1H4ApA1HHv5lExJE/glAxWG3EXIqJk0HAj
x0zr7hDsiiWv9BdEiIHfTDrsovtvW5qNWPAHbvCYRr91hg9xWQwsCjoZNZicitEDDzleKy+84Ztv
gUUJqFQklsCPk+Zzrf4aVPT33E3xFYmCW9Yo89VmdUQ/Pcx8b20UYC3AFNSqj4CU7Hu5pxcD1eVz
diCmzPg/DRQ2GINmlvkIGcpppcXsMRm0HK+dRYn9oqYB47XlN7Y1zMFRxNd+1F9H+wnR+58uYwEX
3cIwphCfLw8IAI1tKbTjycdAcjFdUTvlrrGnfQT6o6p0KjzQulMJunfLp54SLkvCm+NlCJREBgwO
iohyX+7PEZXK52Q+wixHAtmQ8H0zxORa0toyQUDXEdmlnWAsMC0Wm+y830q630cycHDZWt3+GDwO
dV0xYZWLf+lJPhXLEsOAdS93pOm4aFqqctZjxUiQHwbQ/q53LvaYvL0rJIY+wsAMW9f/8W0cxktX
JBw/qEMqejE1dzMNxCkGxW3RqDg4UJEmRrb73idb61Wku/D+Eq7FTClgUt0ciCOlDHuMW0JWxBHi
dDtK1p+Ugp8/Q46NAn0ZjazN1bd6r68REudFc/LjzSh1f2JMsSTDgUXu5K0cvoXVlNy9+AlgwbOK
gcum1Y6eEH5qdEu/YKIuSrZn6uYr6aBRhwLFhT/UU7Nk4hPAp9TUBFx5PzDS+VYDpugfoe2wLW0a
37ZVkSqQZBZk6qbb7nq6Jf/nXd5SMYiSDfWhkbr/1Sj41N0LHrIwalSqA4o8b4lmgFjTzPsSdqtG
L05T90RFQiJQL5L4nCa+RvQC8LMtRdjuBML/eSIFkxKSE74yN5xI55shBo4QaaYb/lEXXIrXzzAH
gfs40wYArE4ftMOzV8wtn5Z5xvWZN3FndMivRoEyBsOwwQH2uax3UW7BMM4IF2y3UT3z6xovnOlD
nKFKCqIC+sxlvO2AoXc9Lklx4mtQkw0CRmb0IjixuZ+YPCb3iPUbzMephyaaJUB5tKDe932NlVrY
Q++piBgFbD24VxKsk77lVvcM8CIosHkQDcMm0Ioa95ndd+lIGfdxrcq2GUUNtVPfwlGjyPilqQYp
q2McoPZbLTH9LiscgZm3O6ffseaNAENLt1dekEZfyoIGEWmXYPwcfWEiVMkRBpmyqns6iqnAlSzt
fIQrxBOxDLIYGM2PMSiLlZkwbRWqmPfr0SvQTXz4Y92HD9wlarn8M/2GjIjq9UEww2guUPKV64A3
+c50ldisfpf2nZyU4uek/SIwrpQKOQmBcYROcPy3B79cpkXTkwGLRx7ogo6TF4yIwdr0BSZ2Hhfg
QIwf0phaB0j5VoME3LKyJFPV2alz3DjJjC6FHZer8joPm/NbGRWUicT2Ejlu3BaaMCDcXHjNZqAb
u+itNKbHqS5tm0XzRXa2FOkTM1SppvVO8H4uooJ4ejlGNW4GlYFOs/yFpHDm7+XNG/Zn/okGmOuh
hcrvaj2pWvOn6DcKX+fj5cOhBJQ1F5X8Rg88OU1e46wpHqqj9EjabSf0lEWjwAjd/8p8NeXWboYc
fNrpfAvYNgmVSAt8d8sgf3aks5l3nVq3ylFRCcwfDDK4pKYNyvcHs6wxAqZotzZwC8WMEfGT0+G7
ggUF+Wvywy4+liv8i01VaEOjJdnvtEveUXVlM3Jy12dtBj705K9+7hg+Dz1NevEObqCi4HbHvW2d
iPibo+CWRu6whVHuHxdWxiGrdV6wvCVJq/a9WkmP/HgHo5jYAi+LTixnPOMrb6+riYuXNZVQe361
cKq7qT9skqhuPmBNM4FCOoMSd7hNof/3raYfYMaVjv+b6yKiygDjF0rRGSbBQRGd6VL3uAuMUcWV
Nv3BWrBPeoo2v9xSxzdb54l93LBkimf/giRSpGCgcqrmX3C1/Zy8aFymdOd6rtOzrxFCHXKFP1TY
biKBwuJ9x1UYOB23/p4lPAWHjzWvJqNI4PKnKDRM1oHu83Oyo+SdOEgcKjQZVA+bAWSNLK2rFGcT
Lj1Y9457Rizxjznxudj9A4DP2mcC6TZMQ7GdBcsPRhl5u+JjOEmD9YVLBA8kh07Fu7bU1zNhdVHz
mtyc3XYd56NUzRH1i48AM7GagZ+C8O9v+Gc5vZGHsCNjDT8mk7L799X+7so9dSjmX2eQcBQWw2Lu
fG3Hk0+ngpn/zvmD64e7EjCzcGZY1GmaPO8Y3CQH1BUrnygy+7GvWawEhEqbo82+I+utK9NhE9L7
CAcFamzXs9foQpyIPn7kFa+bd6Cgq03NcUIIGz4sXlcxW31CoK4E3PutGhHMVY8CLyWkwVjvuKui
fe3XsmYQ1GJRJDC4T1KEZvuw+sntk2xYtcE1apq/8JwR9OS8x73uYY69JoDhpLf+lWlm2FSsqLv1
29zAXQk5jECbYOlUZ9A2KAwX8eyI8+D8n8obKJcVjwwN8L7yShBsM7y6fhxUeHMrkLsBayNxFknd
i1/669f7+Q1khCpjSYL+uPjiNvEKAQYzJEB26O7z+/CXEdnI06HjYrZa0n+Com8X/YRnIwdN4dfv
9Rt6EtaTJQVWEsbsfBr584lkAvxXIEsvWqIOvNN+SnHGipJxQoOEU4TqAnKd6Cgqp64e5ii/uEqb
dKSgpmrcWSaAbLRck0oI7QgfxK8FD5Z/Pj8vEoERth7NPCm9D8o5kGhVx2O6rzqQTreH+OzuGdwR
cBOfDQc43Gh0Z7MNKcCyCHUbEbSXm++dSeAzBGBy24gQGcZNbi2tmn7kpcAPnigKER32tgLZQTIE
aUCA32QkhDO85O4XckPkyZbsuuF2Vl4ebGC3N0YAf4dRwD76ssQlUrQEP9nGBFITnsHFhoRZJEoz
Kbe71OCP1zkD3ybN4jFoHcymLMyV9KTmanY+0PzNYSOEjiOkh3P+suHHjHxUapMgOe0k8zzxHqQV
kNXUIgr/vnneoQTvQTWICDSrF7Z9vskapPU5/NFKPD83a02VB4fFDajb6WKMVr8VvQS0nNh7hC46
15gqtrOKSrkICv2/1xI2rX27BDSeacpQpXMFNTG+U8BXf3AnsoElh1bbGW5lSaM6HEyXApaHbvGP
pgDGlAYL/OwDcsIXD8P/eHRr9msPNo3Z2qQzs4vucQ06Ej1NrjWVZqkMhASdzvB5FbEsHT09pG96
tqzZe49bD7eou9ces1KABP4oewvvkQ/FNTtrKK1xl0iHWj+UoK6YwPq+nqx896jZpjauGlOEvEh3
wOaCDDYg3f4jzSmHg6SfDQbWSXozqfXTWMGv0kCMShDCZ0dfZx+e/gsP0b6NETJEG4LInpqjleoW
YgLncXic2RkzG/MiqbjNidZ0cnuC9u6UZKMkXIK3+CIdZBVQ1aKaLE8XxkjBV8JZZVlYzzGqNPS4
lQz0Uydk4qNoAdbRvNhXbgf5zpeVfMmtLxkWFdjnN0Vm5sw0xiTwK7zGS/PDVq5TZqXzx1ryP3jY
2Blu0zw6tB/p3HYJE54eYmaWQcAn6WGfihprPYZ5iaYBy4EEzmNYyGB/bFshSJZTdkpct8561QLt
28/vpFK9XDpx1T3UKQDY5UxVb0EcwQQxTwk8zIWQwNbldfrNfXdRaaqq8ZaWdNqngEFTQAG9ISaa
oyRSI7Wbk9mF/z1ycVEOySGgFK7NHU3hddWMiRYYaP0lFcVnuYiHin+SyTJQOrQHzfuVmMGT8AWN
LALn98WwHuX5t2lFy0ueFbfOY/ViSxfIdewP0nKQrciKI0U0ItE7dofAnbjJNbpVBrawhSHXwUMz
FWKjf5Ri6Xn6uNyj1kjSpiz1H1chNOwMJxqTqBCsOLD4u4UIO835Ashf2Pwyj9syZ43SJGRuUHF1
zM0tYVa+bU8RZRrK4gB0LsArnGp34KzSkArIoykGpSd/vRr0j0oT0lyotkpSIlgLHmHFWzCjrCoo
pw5lMJWk8+PsEdPCW6MtCKgrec66fkgOjTeZi1tmPfoaXOvYZIIiuksMq2hEbYVlwJYkhoc6o8ON
Wnskhwbg2pnrijBNg0sjX3l6yf4wg2pMrwLLHmVqHE9x+9aNB+k/f8PJyb1uTeo4Olo2eJqgkPzW
Crm7U8fI52u9XUDUuppC4ags34SCeooMrcqzWjFQlbK4b1g7piORI/P0VwFbNe1wDZNj4TW//Kpc
2tKtsY4qriQVD+OcJnfN4glAzvzPjAzl2yGjQOntqf5srn3b9Amrc471FVnMs3Dp2Q+v99VHVcl4
v51/Oii7vAnHHceNb21MaoLrHQJNoNAl//v9uRpJet9scSu1wRuRKPkwfYabmDSH9GBspdtTHYxD
kY5neI8iXTeiMuZUYkFAPtmZJS5gJaEKoDLmbEb9wJliGDnQbfaP6BqDamvdiUWdrCTadugTBgwC
lXyumuxiRvcQaQshGofzYtF7jlZbm38C+nIl1kuWdzSHRklC2irbHc/J+GooLSZ9DzfwJHscNrSF
1S+Enn8w6BouOSxgHF08z8FqDPp/4sPmgtOzXf34wSmgi/8T19xyZ5ysyksszI/mJErY5gVRhXPD
tnBL1FBbAxO2ed/5p/2QpCkIKlf4Lz1yMnLNNnzcfJ+K6dUyWz7rGl1DZrJjDPQHU6b4pTaHgup8
7BgRkDh2vR6N86Q5Roj2ohNWwKmLnDIPwvKT8LOHJMVcQR6W+QogahLFn9OpbucJLpfNoEkBP0a3
K9dLOaIxTZcWCZW6UzBzvKnb8G7CrjylFsaD8Hp97zs9JK4YVViETiJiXlkzrMPvqhzbtILWGKNE
++k+sMPY/QFv9AMJqzQKuYgElfmhhzNy7P5WcZKCaCWy0D+K7ZD3VD6/J/8FRdQ+LGFwJcBho/we
NfbKPSuafFbOK771WyWIpCFu94gqqq9kGraMVaLBBbjpO12o+OSsVVAgQ2V20GDGqW6vE8jn1PEY
SwH9FdgCBaQQkyrb0vx1qU6n38LjS55Nl9iO3y+JdpIE419WPzOY5jtBNQ2anFgU9J3pNypXOnDc
imSUhDMG3mnqWwWTifwI4mj44WLEeGINV3tnw7PLNU/6qmkJhzpoxr7Dcl9LcA7jLRhi/fW791pP
bgxOvfs6Ha8lQOYdO3Ezv1tg0E9zWejf8Faa4/ExjBTw1IScwjfwD/787PEn5HThytPCLj1DIq17
Ok8qRscDarGt8fOwEaZ8394zUg+UMLW14LDUBejzEF9YZ4M3ioOlvWl+qDU/fSB6VQeURaa1k7cg
XzPq4Bjmk2v93K5AWZm1/Grt+LP12eOfhyVhphT4MCnSM6UaJR4JxncEAaUJkzDKXSkYOnghZfJS
mhJPHFW7m4OkbLCgZCMjfF5C5n54e0luIYtTG8UX3F29dcKe0yZlq+jHj2HPx7SY23RmVZeqtlJ5
fjqY1GuFoXnUG7msPwhcigGbDHHt+FRi3AR7TISAxgEAAjnxuT++sB8+5sl2qZBVNdHpmA22N14u
caCDKmi0b4CDNIJGgz6PT7xO6gbnor1TaiNbjZCOqDmUWZU2SITMvUnCXOTXbirdtUGvBg4hfCbi
iQVyFDvYg3De2FdQp5nnbmErwKgoKxa4aCtSE+YUna5uxfxHc4YQduHUcc3Sqgt5+y0O/1wiOKCd
DFJAnt3m/olIhudcEK3yfeZkpunf8g1ZLnka1GAugVOWRRLRXl3xMeRC9prem6R5ZrEsC0RIWLC8
iTzt5bkBXQgGAG9KLJR4/LKMfWpHg+2GGyQw2NQ0KQhwpe8DD9y6mamJQhSpIJOFAcwYcUORTcKD
ugquQFY0uWMgO7kXM7gsMWILcG0sSS/y8nhdpTaqKDlYjuTZoJ2NmZDvI9w0vte/3j8NuG7oeCut
pHm9UHJVg/sqyhGAvFSX28XYoMo6Fadj9f+BWN3cs5H1Hux9Hx/djy+fRBvKcSQm9HtvGt/a0FJJ
LnIw14SNm1BJjyyD2e1m5qSq7cfNYAnUeeO8OBSVIJQHBUCjeUohq0re3mXkUQyICULaqqVTewbu
1jaF0nVPovbK13t1uXfNnNad0NMUTAQShce0QBpfBGqGQjJ/P1+YcjpLjtoE6s26UvBXFueiv05x
pWD8LjefuB2vqe2Gfh38Y7EWa3N3MBluwUQOy97JB577fdMW1VWGHYV4Tb4hK0ON++eSdSkzL2ka
h4b09K6t437gQUh2B2YUH5KQsiD1fF1okuGIb0GTFneGk86LLYLi1+EgeTVCOx+zHEFZ5XAvFcYk
Qi21Fxs3x210fMr3/Gn0dKhhH0iQByZsuVBBgUDrt4tfGqE2BYuyXeP6UDqD5o+FZylr26twanzp
Jki5K9KPwSsJq30vgv13O+oVZ6lwPJx6eL/hUBIDYQFO6h2kiix+Je7wdr5NlxArAJH2vMdTLeKV
QToJBiDjkomZQ0ugU0W7LQ6hovJg59dexYayBSOLe8krUjBnWr/1pZ3mLHji4dKNWDcZ4xunro8C
41gqM8T5UvQmGELTtkxHONK39KvSm4D5k+BajVyXUqy6ErX3lcdg04TM2ZAabZ+QQDB8AqefKOcS
GHWj4cIrkJOVQ7XgAHLACSsz7sq6kFOKoy4VxaMjIKSz6UUtHHwa4+uGmNTMdAmBfdzvvtAHegKB
3OuztjBJwQQMXxvfeQm9LmiCoPwICnZZEHSvHnu9pG1h7rR/OieD1oqxuKFVc4axaCNkjzKoTe/p
U50yB5uh+wAy9fU14zVNTklHLOcBNj9fOOMiy6fwY2LF8Sj6YBQ8Aez1q3mMcJ5vDWE1Ew8HOWfI
v6cEo3zknWih7NTSFP4YyVuH0tKbVki0qL4yqyY6rjubUoOdTSzwX8KhoDHBteA0oJPzr6fJ0rbA
+kUxdpNbscg4p+KkwEfHwNTI+ZlnakrqS7oiOcKs0B1kOhTF5NxaY9a98DduWkXSWoRktVJq/hPq
EnXkQzgCbyLn1ZOEqNOlm7J5ZcX6wmgrqxmvRQ0G06IeOivPGu1RhaE0TyeQSU2Kyr0RtWACofIZ
OpF0JOOt4IKOQ+3yvMRarui6Xm1SdyqAyIf77XAHciOhHSVaRGF4xR0TsA7vEAo5jcojQD1GvS5X
NQeDk5xiqJyX3IsB5WBRmcGWdgGdZ56hnb1yIvdn442oLdANTlZMShpw6daXJKGY9X0pS8Nqz4ze
qr/Erf3U+Ka8eFkDgRkU8tEkFJ8pf9hl+H6/gHqkN72KQF8dGSSbNgsjZS3HxiCllT0GjAt03mfg
uXqn18fJ3HfV25q+hUVxRXs3KJEb01uNkaefkC/RycTRs2fQnPsr0l89u3DKD9kDOpqDc4RndOPw
HMAAt7t6aH0nkg720zEB9kmZP1Tek9HQczmsSkoSQSxPIp8mLBq5CMue0JO/MRi7CZ9YwomJrBeU
g1BIZ2LUn8PWTEI5QPLfoXizgwqJA/gxv2rBeS0FmHwvl2iJyTTiMg2bzjeRjZj+Zkjnit7PrCKJ
xkZ1ZLtDVZXxHPEqzWOyHf0pQzvHwSt7WQ1gAAq6worpvRuH09SJauc5aGtA/JL2Mdoe5ibMP/mm
aE86zCTSVtbPNBIIF05e3VhqcyjTpC5gRj2mas4bKxHmaKuzjSt8UjvRdCPU6CVL1Jke2FgK30zA
MyaZsuOk3SaYjxJvY5yjB/1oQwD9JawBKI7V4DX//jxqkm2Lns194+MywPaGW9t6Fz88CX+IpRrB
cKh/XAYHXXeL2md6MJzKUSZ/ScN8zWd+QHcDE/AeD/m2NLajSehyF/MohNv6b6dZ9SlXaU6A3RvW
zhpA7ABeUij818SEw8gCOtkbfeT/UTWONeSQ+o9+4QjgZIMOx9mwYuLOtNMBl7LzodhIvMYf9PXc
Evd1jc1GxIhet5H2QT7uwlyk0SbDgEf2IXP6ff+7FgFe8//2Sdd30vwumF2j7ml6TNy0+ILfhCdS
rAbCf+iZV1KxrJJd4az1xTvNUwgAxGOsieSPAIaINmKGjNqTnHDqk3un3o973ybLQFMU1lccA2b/
6K9eUaReleRkTbAc3zM5BPS8Qq11F02JzDn+pHldbxi7Qck8uiMg76X9GsOk6h1Zx6LkhgkbnnC6
YEjq6Kpvlfff+0Fx7WrN6ts6wPaAMKYFpkWoapIPTc/XlJxNmR/MOw8whG5RonlYx9gbrrzqpS1C
Kv4Uet5076y2klRq+V5Oh+brN5g1CxU059scaIj9r1ABpNiMcRqSy2i6cL+kxcE+raVVxz58uOBM
p6NDe5R0DQ7VNJP9Lm9fIcOafU7y34dWXlPujkcCYhecZrCDb8PgRJdPdtsQcwib7DxARc+yWfE4
wpp76Gl+WkyWQrFa9Wt79yNk3D9plAnrzEvskVU2kWS38M8/i6qVmSKLKX4cHUv1Z3C/y3lmnio7
YbcoCpQO7xuAKQrSdj7Qt+G33XWxevRE5N/ikAcOp3spcs8Vd0ystYv27/j5mXMU502mQS1l+Sdl
iRFDDMTJv/yovFMGBYFVoqP2o4w/0mFlmGbPhbqycsLFUQRJU3wmKP1Lea+AUYcv7tJ0QqS5kS/z
KZyUQmxsaCqnsaHKe3mjAo/OGVi/AhWZYH50U9thXJcnHrh6CApW4VvYJ+veFZtZn2Oef/NtzU5T
SB6I/UU6ewsUIfSJsBoaCcgz77gY4yh+gV5t8/+lU+MuNQo7IJpopGtBZvs3YY9R2BXZpo4lNW9B
dFeP7gzuDhxQCDSTnsrZtb0j9DYkPx3w5rKD5c7zRXZrBM4QE2UJ3MhwtZEN8vrGBIef6gCYxMAt
SZPZBhvhaRWXqEZCjwtqBUDoNCHfctCEPvGk60Ho2+7xfaMrA0GlLZDabRqqJB7LwM7P591jUCSz
xkth7n7yAv1pGKFloZGYsDNkbPPyevlHz7G/dA3il/kwyb5I9V1MrYUmEzGAm1R5pZ9xMYYa7MNV
oUfFGNvqPBTyLK9NhsyLdAjpyN3ItHJU0Z4iBu5kz5KQTgVTlccWwnSTQSls5Q5YHkDTr8nv42ej
DJgooRvqUuaPbwL7iznznuTW73mlD7NTJLNAWFx0xP0xgBgVqip20Rz49epcUd3fxlCE8tELjpds
NCv3yrajglkMvuw9EZDePfppMN8Cz6DhdtU1eooYLAfPvy2qqFg+rfOGortPrms1SuwvREiCPneC
ZGm0bxfAlTrnSq+6t206BeDzLQP49KciTCC+pGTjHNAYH6AAgmOK9s8boJMbgADnxJs/1MBwxby+
mRxYfWAXcdT1KjMx0go5XNPqo/9rC8G6JAZELbA4iIXTXBXI/UaAGm+yzZuNilBBV4OFHVOiSv5S
L8m4yH82I65QCaM3lVFjbMaqnY4V7rjsvV+iP0MwYT4gg/mF+p7YCl3GaqMdk0E9cS68tab7Q+0V
pkQzXowxtNJZeWXBTxpKG8vcC2NsOhVTEMFGCL5auNw8Ek2nb/QL0y4sBUYWlJDJm6uo5EVFNA+F
pSRe3blT201sVYMC5z2DGe6PkcKc4gGT2R2KpovO5GLy26M1Mmzb8VpXxYLZXazOxceM1Z16WPhV
FlnqoJkcQdcuWOTIeZZFCO50FXIMOtSQnuFCRgo+WKvyZ4SkLbSAaj2xsIcIv/kgoGdDHMVH6U+Q
2w8Jg/ynV9pErb8oxPSOVXa8rGDq+44gjioSCDzXg+cJANnAWlhDSwuqFD0QvLrYxDj6tI4Odml9
fwaE7nuBR4wTQaccl5wEWCjOhXobq8OkCFqFgf016JOWhSblasEzevfdccOu6008iD0F2EBBJBVS
YHedX9M5a7sfX4qWjyLegKdv1y32WG7IUokEeMAWd8sDIzNr3YH5rbSzFPqT8YVrdHSeraDZEfMr
rHM5fX5hgrxK68Io+4V8AgCBGegNMEztLPgb+ARJJd5o/qHw5mIJc3epypA6n+3nWDFaBttAqTpb
tl5fzzOUqqff2HInTL7Z7mn7g/yWMLxM67Jprmibsjq5qOZ3Wcxco73HOsHj5loBY1KSXBG9Edp8
NueDoYuT8Iwu1lRU1UquEVCWx2JXi1suuxYdx0yMPoSqlVUaA4zToifpj5WMfme/oYLrdjwtAemE
jiVDdwi8jlhkTlC0PPCrEFEIwmiy7cuLBhUaC0/7t2NsS6pCyt3FLXXmAEL90QkGiIpGxVfP/iKe
fgWU0W6oATk0K1F8iZR7TJD2dGvo7Brcc08s9dUThwivq2SIuCNH/yjBL2qdviLRq5+QTSyKtAcg
b4f8bGiwwGlx1xEn0HC+Nn7Er1+cmlNkm67oZBSQCNGWIP7fH7vU87i1++6e+0xSMKpJY6S9VFL4
tydLDMLNtWX6tizF4mtYMUDNubP9EdyiCfLA6N88xb5cLZKyIv3J8ftzN/tqXGB+sSj6mFLbt91O
KSdtAYYyocL0CI3oI7W4MFLylNyfE9+ADgtFD0JvnEbFRbUPKgf41GZ6+uRyxIbZ2ENsga1t9mN0
u25+S5+d8t0Kshjenq4YgJMwXD8UV8uDm9YjFfsoJzlnAnv3CCH8USx4X0b2XkAUXc02gS3bBqnf
D91R9uk6WwhZ99fZLdEOwb8vm3HikmaI0kcY4Hf1HVKlU7zp6S6SlitK6nskaujI2nhRUPvRVgIh
QNtkYU979KVHR9Zih6LcxpkVWQgipp+EbgLW+2IekFwUMRaSNeiFI36+BkIGUR3Pzn/ZWHneQNJy
hP5qH67IxJ8zUPAIMpIZyRbSxItYTgt/XaNQTBs6i9ZUj2tNRiF45a0toznetnvdgHmr+as4+w7P
HhcwRhjXibkIZ4cJD/5DyjwUsRwem70TsWLuH15T0YL7GJusXlyeHznoCa6mGgoK1S0rE3FYz3ep
3bOliQqjUxIugZVIPpVJUqBW45AGQsiKTYY2VrSJCaGuU4iJul7ujBIku9rmB5nIwqwCWS6KNcl6
41o1j092dCYgVmZSR9HsZIeAjX42TLjZrgg1wXHi+Zc9q9zpt0Wq1CU7rKKptxha4BhUm4/Usft2
P9lCiiYBHpb/71mw2AboRQ4NiMJqnYm1sFPkakVXbT5RtqB2nlxzs1ymRF5qYe+OpV3LOS22EUZ+
2vboqZr/5a40MyDaKWRo/Xe4sw7FZP8HQ6Fdfbow0amGGUMsNyZ95hur5Hl8GdE4mla6/YrcowRb
b54EtC09yQEoR878KaqHSDfHPWrxuiWWb9yve2BqRk6mUHdoI3z6l/nvUj4DzQK5P/GNNsEk30JT
CpaAybPYhpx6sAGQqTsspQzsrXkm2DXoXPGKbPrItBbXQlXiTPy4KxTTDdbsV3KYLLZR+65n8snz
Qcpd/245pHeLJ/ni5qQVnh1QqInuM3ziYbPUJNdkctHfP3QsIHclDPSXa/++46cUqumNzwD8Ckc3
F93HgliV8mqInVhr4BNtPpBw7MEVXN7HNsX5dCdg7C9LeqiR7EWe5qOtLEQ/2vl0xUzDEnhLXSD4
64xJnycfs01/jnV+8Ni9GqDcQXVJjBsBcOTs6tNGgL7jNN1RVYCUzTNsLmQwEi4tgd8qLqWbQ23o
diz447rKstMWPsSEWtpeeINf0wmA8CzBlK5uxXKdJcO49vSTNSJgKZfReKR6aPNuGXifWEeJLtZh
4VOA2xZv+bwddnM/BIp4gBvIHzQ9jf4bsx8zADIy2lNnNH+eUgQfhnadfyMNRWqd8jrpyZ6Yt6kr
5IioEESKylqjTAdtCtQHRCgmBui/9K4+Lb2zWa0rfYL+xajoLyppzJBWdPFi8BJTpPAxDur5kcIr
7mH7ApzfdQk91LqDYPfZQqJhTGL+di/MlEMrU9A9p7uIGRYB7NlEGjVoOwSNvfsQw+81+eYQ1izf
TCpW9kJSj/P1+cVuS/AdLjx8x+VqA+zsF4uf9x3oSmxSCp7v9JqdJL948zXSVpwHeROLjxIJ7Kpt
rfiiKLe8PNkft7cRg3lSsFp0KmsKAURUsQ9XCpQ/bN/O7nbyU9w4W6ojtYigZrga22mgvNWRbxst
ISgL67YfbXzf4GnyotAdV6YMXJ1BcNJxZY82L/MpiZA13FxwLcD5fUQnv/5AB8vzf/WQAoFxMl+w
4DrY4O2p3sAXdb4P0CRCTR11GcoMqBi+V/OKgh9+rIQ/WYAE6137LWg81gPIpybL5T0C9x3IOzC0
aMLdh/BMHTttdUaxll7xsBj0gHUy55O4tDMPmNS6F3oVWzDSQprPKMitLwdcZ6OQr44sjF8fGRm/
zXRfCBue8s7oqEyQ6st8deG5wZnkWB7LW8kBjon+Vb1nJgsMIfBJQgRR1uYu69DSjVibCCwBOFEb
kKoJh5KK5A158eO5WfKso0ZWuWATGnzzing8FpWIC56bMkjim72ck8GkruWbB+L0CKn1eXkhcoCl
zYhWOcLzS+rTh+6ctoQYsn9VsveNXrH61W3x9yzEocG9BWZArf9jd7mX8zZtYZL48dQzfH+HPaPd
pVIrf9FucbQnk+3l9SGiy/aANgUoPTFal0GGQNcyslZt/PrewDeYW44QjuThydKrYSsOaTDGRWfy
C3tktBl4I95OwB9t7VdAT/u22plkwZ+VxZNaT2/M7063OH9yDX5dn6DebEEJxdQuW9cVUrlz+KbC
1zmAKsZISdBVntRwtYvp2En7MQXr4v2k/h/DUyzW79hdD2PmMKzzUYRGXoJUH0+MIQzycT2j6Q78
tu/r4bVpeGheXo/i0Sh+e5ZI/Zem1sNLxGrrvAjXVVt17p7aVxes/K7NMZxyQvIbFc6jDqJX7lQM
PhDXVc5zL0VgKqYdneBvEvxCbWR4FOW6isru8TnOTbEp9pbKBTSXmBgSduRZWGQptaf9oi1wMP4g
K9o3cnQ5oo+c9gortA0KG92JEAcfSw8aj9a1YMQPA5Inwad9EFaM3Vun54z68Q6el/WcQLzMmboT
C+BvQwxfGaw7O6gt03ohjGn2Mr1Zi1yz1rUGpEEfPpcBfcR3jYesA9edxm5SdtuQoWRpJ3DG1Bzl
zQ/azcM+id3aRiPHqd+zPqDBpdyqYdQ1tgINQSYp6e34FTzauoScKtOAPg7JKCspfVX5E3H/c118
FqTO1UxwIpAJpIB/+R3XtLZJUn1fsTYBl6sk41UHUggJaWAZy6PoxBYeRGSbjbND8PTSejWyLg30
JjT1BNWZOYo1x2AQnO4pIiiQw0+C91dSu4SkauAOuCwkjxrMOUCv8FLlGaY2L4z+z2+NfDEBFU5m
u99QKYv8tlnbd7Zg2XhAJJ/nuIxHaIH9l/x5wXmR5ifDuB1v/dyPM1ftEnJzc4N1Uup8Wh3m20fa
2+D3m0+Xal/jdN87wTGl/C4F5hxHdQabBg3PqVHdV97+zCw108voZYEALb8f8DJ690IHBa8qKMR0
iWvz9vudsIoggAXUnSS7tc3+vmuzGx82jOvOAu+g+7c9J3CokW974JZ6O7+d1nOgKZRffkhHHY8c
NNvGHEkLhJWXceZ19u0wfXE7LbBrWoq5edCb2vZekntWGHLiNQB8tGVgsl6lmho7HHNYk8rsm1Ex
ga6+/3sF6ZinMVmMNXzqYrHj46PrWIJQAz2EDc3tTUwEbWBmaIiioY6cJauMUPbyvH+CN/Kh8mXf
lHvg1zQT8NzdB87065WEwtk3Y21m4btIQjvofDngAwPB6/jvnx7+ann8RwWdMbcSEl5o/nWMQNCd
J9MU2wqNvuNW6NntyjG+LBHk6xiGIngU5HveTb/Kv2S9XdwEzQqvTLVncE2lLyRhmURuQa3sJyin
YyEVvjeiDsOmgCKTdhpHfSdL5+40bENODDg2fX2rjolmrtl5HLpDb/Ah9EFor1aZsUsD9V7zxHMH
3Zg7bZttuZLOYxEt5r2BE/fN/R+JI19LAsh9K7+hyywTxk8/PFdL8xDlh3X0jO3pqtn6MEOTp/y5
Z4o4SllinhcsDVSRRNmGmbH+5v3AAWFIG4CH3Hw+00QBBJBfMgzCq0FbB77Z1Iz4VN/hzcNyxRJV
P65vLmpDkMoKCK49b/aDYKyOURu7I9WQ+fvlFifaOiF9Lj+n5kcQmpt8ccjItN5aNi4fuJhxaAs4
OYDnKe4E4y4hvuyXJl5O4qAuiwNOTa8e7WBSNzXMzCnI0zuL8GKTQcFiJzKqaBb2VcMSdKFVO32W
iogmilrNSGZHs9H/V4OZuoEdGOzkNKMpoLKFtCXBmhQ2Ve0UFFLhEXlNYQiJm0IO3YDYC2TwmMKy
qL5WQJjpuorg7k9Wx1J0GZ65K3EHsxM0FvYLsq7ArSqgIJ8vchorNjEr3NH3wYHNC0V4005DKDfL
9uAyopyzT4GhfOlP3HRXJ5yk/+wyE04fgKKgS3ieNzARDUr1K/pEcM+lwsIhw7557y4x2HGD+YL5
pQxe62cvlZ99SIVYmxG88Cr817IWRW5hEVjot6j0OZUTdugKSVIkgRgt4UqsQF/caLJkCTdNy9LW
ctrzftG7hsvH9DTGZhRlZ98JamPOnUvSir2YaQN7svDgjUOaa9edpuBumXGqJiDlAwFwWMf1t3/G
O1olY4JlWnlTaT5p8zfpi3dNZq0V87+REK+6onyEqarj8gT4CBCcUbt7GV/zIAMEiBI4CaWmIg3P
mJZvT7pAzJ87PrvxJiYFJJ17/Sk2AlyUaV4DdcpX+MCyWX/q2CslGYDZeT+F9ze/9zhoeUzA7Lqe
HOon4hqskDoDRX82MkmWAuzp7KfaPEA5akxSGVzihH2GQUHbK61QErOvluClP3SfUDgHvVFh2DFp
t/y1lBJyQy0MKLAwXob/5lTDxYkyKw6avMlSJC8/7UVbCZKTfIkdFnj4Huopeh9bPLLQ0lCEv87k
qdY/OMHs/Wq1DtgJrOZVmL4fL3RaOQhWvolaiMUMD+RRlLhHQsSwuaUmNcLys1oWnh0a8ohRAZW1
C7kBxWux8iRHNbJGNj22u7E55y/YtCgPf+NwDqXL50/XWXHwy4h7XpbNYEILF4dzJI1I2os6luM0
Uo5xEBovEr3ypCRHIO0SS+Yvnj0ZVBd/KkOk2lrApkFbY1PCGigjqYB6o/Z5XD2Y91Hg/v2XF72J
ECk5NWo6JY7/MIWRoW1+xnaZP6TYmYQhRLifFeFS45jUf1U7Q4iqCwtLbWwTW8+gwOSZJhJDMwEq
0bYeb9PVS4yEq23927KLDbG0kc+bj+IgvgQydregydz1EevF7Z1jX/pZYNsxy0+M1zb7uhNkvGb/
AyAF7ig1Ies51FQdFqIZJgHHO1QyCwIukV30t2rTZQYWbfL3Evy6nYyW99a5in3e8jShuz8S8Umn
TAtz2zwSBPg6yrI1z79316N3K4wnrUuzggHsYlStHuRkA6G1eweotkfZNJsUpjWLMIH6KBi6qLRC
00XY/Siefu3zzctq9t7gl42xFc1fMH2khoyk0yw/wKV/kzmc5DVK/x3JVZXOXjwAYmJVBxf9hjMd
/J8JFQJWC5Ep3JnYwOWXTuPUxcQo+uUt/TTEVKiYvge1nhczlk/xWkgrQBo6uztgO1pPAiIN6xNf
EuNOeK95ukeUyMBSosHHQRhlp12dxFfRo/6pM9lihtaqYD2aGR79cA8ors/nPtyPBne6SXpss9fl
g8IRzWEOoYkygqaFEWhTxGrevA4MM0vcE10oKnBnM8kKzKx8IFtH/A6E4VB79DFHaY2paKVkDPOv
sSzteE7bt0aQp6yTw8JCCX0TQIXjvP7l6BY87SldWyw0SICoYJvDXqHps7ZDfxA3ez+15edA/Ek1
a9+aWm7jb7ZCEaskGRRQNCq63yx306b8WfIamfmr7tKpHWHzUhxgKYjkOamfdToRQ/TwoDlvJjcb
7y6Obi+cskOaZlC9rwiqu6nAxbhHok0ko1ricQiw2SEbLXgqCEgN1CVguxJ5mSDX+sB7Ikk7h1Ic
1cjK0ItKbDA/eZRvCrdyEgt+7SxEQyi0d01I5rhtMIrB0g2tzkTqIMoFsJetIEv9jRqGda6FZak/
t2nuoWE+azgxrJjVV0wjx/8lfAIMpDKhrpqT6Qxya5ErcomPXLIcHh1ZtwmGQqJDevYFKxswcYbJ
73aXSpp7oOweX6UM6U+oap+h3X7kykQvwHTWMVcYrIZiLsBj8HtJcFbl3j3U4wQJnBEfQvyipPOD
18eELbqc/QYTTFOV1bDR2KGAZdmmMAmm9mNWgL2QkgkquST8NeUyYSRYT9KuZ3hyPbIXbtYboNir
LB+/OS6eojhkFn/XnRyegfi17t5bKPMf7ARdPeaxlxBL8WxK7Pj0jzDNAFenmUm/GlwDnGXnMfuX
o0I662jJwRibaPDpdh/S7avjiRIakcWAdHzqA1yK/5RGxKsY+E2gm0eJJasLprovMKb0IH3gucUt
KlshYjOkcQ8EQRJsixxLHBz+kVZ1HvCK6sbcCu4U/BJm+MngnVBCU09NAfWZU+F0gOhH4Tqa9B7r
JvwqsYCYIE5TOlwk79Afx+VonZnPGtRBbRTZP+Ea6KDYs3KPcavgA2jm4Dr1DbmHi2vRbptUiGdy
VfHkIX7Tywfcaw0dBCiwW22yxD/7jwFwQuDHyOHqsL2Zcvow/6XoK8pGzZ2/8LVn7VuhOYdfBSvY
Ywypnb6LpIAW9ImSN1U1cDZ0Fq/1nYX9j/PZo1zg3K2i2tJlzHpBgmaUshK07undYYx08KHL3+C0
uqrhnRM08u5HdcU4gkQnDw+5dllrhCf7EnB7yCmq4cAk4rnNT8id0AtvISkY2XnZfPhAdbL3h1TM
mMTQIqPwGUq1F8yqDtH4ccOwzKfQ3bQo+avh4IkX5FeFSicMcPE4egUm39w0mzPI2ZVrPa7fKwIV
+Kariwh+FQ7UWhpYKpaEEFJT4uuisM4oZU8EI4kQ+iGcveRWL05vHCJIQMVxzWj/NlCWhqFw5BD3
LsbsJ1Xj+U0vlPAspUFfn5l/RmmqMgsNQiaZ3WDNjO5J9oPk8AzyQGDSgmmNGDilFSRc9IIVOQB0
HlJP2BI8k3LEhQPVKGYOpTlMoWwxOhNyETT3Qb9/3JRlJS7xaAdaTs/dKFZcbfv6QKBxFPDV4/y+
JAVZrcWwHRxOMNnsCnwwspWWMwOBDvCCkqchhIhVfOodiX0FKjDgqfiyTCceQUWHYtQVgAcIg6Nw
NhZ6ziV1nnJB12rIGPBR4nM1npjXNBvLszS8AnJxX3RtqJ3M0hO/H9Q/Fmmga1fAHAgJszHrItmC
3M1kk8JkfH/dV+Qwp5aQCns3rqXf37rp/qF2eU5lfqBjTQI55Hj6cm3NCBTkVJMmBkMp0RrtWNuF
JxXCYMKRwi4ZIY5JnRhM86aCVGRyyX8THi9QG7EBviIoegXxKOg9aEx47HGhwKgLmjXJ/uHP0xV5
RZvST4ouY+vDsDPkma1xuspWAS56nJHvKOCONLXEVq5/nZEjShGd7TgMUMFDhmICT14w/+R728Mg
gMPgmVqDeqsgIuCaYW4wrE2+7SLMc9f577wBkbqAgrRxFsXOYDB13cZr/MB3lvdQ3khPAZRVPGCH
JdcdsDktEaUqm7TPfqu5GJFiS25wSqKFo1apLvWYEIwS3p1a2jLMpMdevmmOnyyhQdymQRGWRRux
5TGhwpupzF8HnUtcmgHqEuJ3dqowTWogAghaEtUyZpFvf0HCGvCHew4yleDcbJnbwxA6tkpBY31H
6cucYTijpy7rliodIRYTO0lbXOQino4ztarfz5xIhk0tufG85bqrQ0DyRjnx7f5Ll4FFhucA6vyB
gKgrnMpDZZTs/5nqSlB3Xj/L4kFG9pBvUqmunn8HzTP2zBbCB9UoIieA608itTc/gnygR45EjSiN
fJntZCnKydCwZYSAzISnimmnuZeEGoxrNrF8hmFZQRlM/vC/zjrXagIK96But0fWNjPpWZisMqGS
9ESIRJ/PLESvB8kkxpD46TmY7CGEzTuhWoFjsFRFyBek//QpsEFA4WWoB3KecM6J3HxgxSmSiTQZ
EmYK51tEG8PlQj7Ks96fK8/qAEifR7ZaHO9nL47Vhdftcu8/XWAb2aaeplW7PgrJkgpqZWwKif+J
Zz4uoMN8q2FzqNifFd8dpg2kyTS+z8+jIq7br3eVR6eDEYM/DWc6H9CJFe0ebqpYSgpOmG5WNEQo
SvztM6ag/mNWkkrD2YvaNOsqp7aUk6XCMyhCGV/Guu/n3+ZhxcXWSA7pKSYbnzV9mKjT004nRk++
bDOE+zn0HXD78lSNdaqoJQCPB+bPzlShzJ9JbQOtbWsL49kwON1bWHEVCCp3NYRZ7thMMpg/Bj+t
eSVGj/FVLku4jZIg5UbTf7rnCzxFtlNI8Y+/Z4qtjcSYGRyngtqKIoXHzrftZmsjbKAvO3iDu5d4
Te2ys+1MQbS3iwLZx4K22xGYcJMfcIhi80MqfwBkmxLZwWKAWvMdM7vNEpQdfezgE59AGxwrv/k+
sbNAbsyhCog82ut9R4br5asDNkKJjbv/07Dny33LmKAKKDgeJKBpPgvb3FABHHDbWWCWS7nvY3bB
KrAfuFsMy74+i2Wzmzk6H41FfYb1oJRYUcC25kS+yPhCbUqMSNLKVMr6uUXKaLi4d4sJJxsJjGks
oISxsS8IIPsxmoqVp8fSA5xOLx0PknBrJQen5UaRzM67lYgaFnhrygsZpVx4gZZ4Nvm2bwtN5BfV
63DT25me7MJw8JYPw7G2dR3uiDCkQDAlEVl40OUe1hK0LX9y+Bs84kKCCP8/5fw6Ufj3AiUKydUD
cXdF8PlsyU/rsCXMbdPNquxx8lgt9eMumyFBQrMVwBH+obq5ZrRp2o8ZCrK4/RzZxS4eHbXL3j5u
qq/iMhj2OauRDyMkMVDmlSqVkJ990J6wmEoYm4qb+EITwsvrPM+QaSAp8j9NpqEr7Oq4+s14VQ2z
+Dkwo5/WkqtPudSgCOYq06tP+OYYCBOH1RCFXBtztjkmckB9jo+irl+9HTfmMmbJ3zc6SUioSltP
LJGopUKNuGRWXw3ob7JVbBQMcMzWwKUWtpj9H3w7srQaOZTJcDM0Xs2PiImHT2/oEXYrVKn0ER8/
jm3Yy8jpi0+KZc3Dmc3jXIti+r67B5j6TQRLUycwq2HGJbouM427EQkqdeY/WGiK6GztN5H8ZU25
PskR7cVWDbznsFplr77Im0w2nBNvtrgYkicDRIpwIbUE5ts9F9gqX6VPU56S70kF13Jz0MnU/xkU
rSojDyDgsNiUpc1ZfuW04LJ2blym6hA1o4fwk9yxLtecLLe47aXd5kFwcKVdpDnFXFeVKjqwQptp
JR7fm+xuewGS3OLYwRuikJEN+enAAF1cQT4em3wgimOlHhZNJXtsJQ33MBHEiT0jZ/VxyTzl+sjH
FeOUfXGCT7GXTzVv1pyVV5RHvl1in8Gprru0/TQxqB1b8WmeuJkZ19bsP47W8+RcZvwmp99pLreS
oDLZZuY7sryYOJit0JvTHUxxgj2/ZbUKKHSQQ+X2zg6tIaqHhV2WBp3exz9BBa0ZrO9nSott48JS
r0pTGBpWHMbtlqHVb31073TUCEYd0e7atcmXMMxn1NeMPtVc7AQCwRUvsiiP4s/To/oUo1TqwM+n
hFx0bjS1xFQGJkSaxB+XAXKRafUSkwMU8I2icCFAY8SPpFD0CqkHLmO2tW2hMi8BKTW8jUQOwTT1
jAc0cOgJEwghxa2v3bG/XDr7PWYSNdjuOVDsCxBia5pFfOfjEHtEDyEjqAn4PaS4nntQBspQtZ/+
FfDl/wcL0gLxUbH/XjGIqltfR7GHrnaFD/FcwSNDHhLkDKS+T0JP3gvAP7W4Wpkc72It2vJD0YCB
nl68PMbnEwVn3O76+hJVDnP9BeAbFDSJ9GBoBg1Aw9OPyys5z4e4U+WnkLyz/K1QKSftXDYd14eS
JQSMhWobns7m9ttGrXhJT1Pn3Hcp6xN5f0suporvcORU7pK6w265zdL228gUZDRvqDeRLygwYLFc
C51gMjezTpzWoCLX4vxyedOKgyyuHySoRI5QWpBVqNppbaYGyD6mzD+px81aP8H83iwVy5fTJ2xP
Bash5UTpX9MAiZSgoGTtg7a9KBYWWDll0H21U4954T6mNP0mDDQThTh6RUp+ct93NVYPh5Ot7uYM
OA46TUXn3ZEbjb2sVcZU6Cxiy1WK2BvS4wStx1j0hqo8C9UOAe3oWgF2A5DsQb7oiNUVjcLdr0k1
wob+cXurgAQ0eFnYZQODKbsnjHqg/MBxFhXspF/d3wi6C5vnssrvIPGONH7npBAHRrECyGk3psgj
S1ln/qvLT+90eg2hfPonTbU9VwBGZecdo/0ynIG8nC+Zb7VsRpuPMMpfvlDV0WB1nU8lBXJaagXW
nzXRjgSQHQBnf18vGnaIV2FU+dcJ5r+nB3b8iVw9q2LyLQ6Bo8xSEwkKTcYEfF6MGkd3jtYBfOBN
OBwJ9+W6DIMeP752mf6JWrcksQiW5dsBLhZ8vi24nMp1dRB3uTZCBLUEdzjv0h1G94WfIJXKU6PU
g3n5jVCS1FTbESnHVjrKtk/JGiwW0We3mZk6ah5jpQD6CBQ8i5Dp2bxz5dNcVZNUeLsEdBsY++AB
Dy1pAG7m2p5qXjBLkT3XMolQhJiiHPk1E43rz84AreC8KadYaaugKngK7pbu66CM5IFMb1eRF3Uj
4kUYWt7s41kLiyowgf8ogATGn9HHFGjgL3sbf05xc3RCtHqmWarR+XN0n1KtvWViXJTMCv0nHVh/
w0m5bC6GY3yWCM5kvJztuFw6nDF42maAWkwG5b/kBuKtD549UqHRGVVglLX2xz/RTYIAeZaEmxrK
7rrI+awXTkhuHzzOOMfLdmTNMcA0cBnaW6RsLzqdYK6PNzsPNjjbISu98cxvord7BzIzkyujE351
xaCY34FaYtx9S11zsJIDMPCBA3ObDF1BbMAYKH+7xbRZKKTroruF/wqjv0TF3fCHqPEpKX081xQR
v4JXV0aj1uGglnuhxGF2ayMoXc9pTNkvmrk+FADotyoSsEtyGC+xwMBJJJFFygaLFGAQCImVYzVo
VJONTAQzrYU7tiZgTesrEc+THaBdnVErt6G/6wqf04YYVQ9u14OzOOJll8AUP2LXHkWIxh4hSs3s
P/9EfZee8PnG7BdQhpbAn65AUEk+PpCse6oFXL7VhqmkJAilAGnaWoUJLeeu3hLk2Bg1O678Rzlo
M14j+CS+RoXVjEElCb1XIQUU8G4fIA8Hwx9fX3NpjvLcGibXpYyspNdoWPi2DkuhCV7NTVtPsS1R
fM4zAEhbSvTcV6uK1DCN/8vzXnaqtp47Vz4YX0tndwFxZknsUcytUxPSckvwf9q8cXP4V9PsiHRF
mo52WBs/05YULO71MIbSXqwphjwvG/vZchxwLQ7dnCk/f7PkJyY246X1TaeivtufLH16S+m7NlEF
xRYh3ZfmB43Ls0yex+l9SSdSXeUXPOgW9xzGgCR3t9/ZHjy27aOTmFHw93d+og2t/BdaUPxIdlp6
Li11K/MpkCP+RWWs8txPhTCzX6/mbul/8PnWbdnuZpJ9bmLKDehr3x5JY90FMWB5pn3KKd42ch5X
hLGfNUcfL/Ozz3zy3LBvWsEf8h8WfELtiJ1Y/DvvjxHweQ7pBDwzhZseM21Cd8Nh7OTHyrDgZ6wT
0/wZaIWIMbKi16Tk4QM5avRH/LWHE4p9mfPxjKAPp8nlfYzHVdKnzJnV7iIGSF7kJnmPeoNQksy7
1rOTg1H0bg2U78frEMvt3jP0BNWLj6EEeeN+A/B3tnGE2BMXiQE4r4TjBpRk2zcdyhBo55xTEKa9
RQ9scG3OrXRX+DfKErLDJcDlCCgmXTfFkiymdXQTsQwNl+5tmGZPlvK3pd0z+v1KHdJeViGhTwrt
sjIa2iT3TyXZZjlR+HAQI6nNkX66xq4aqUY9FbMUD1yZ4GPzrH1ofU5YYh3R6XFITqMwMiu2yI1G
h4SXCxW+spnjICqT0gTnlm7J21EKRRdoo6gFhYFyIvu9Bvx5bpfo/Y9dQAP5dGG/OcLDaayyDBUI
UQ/anACPJyd79s/816ymW8TqITo8ObzouOj5wiO0PZmVRszNgl0J0/+iGhoBFjOXvpeoM1dbNw/s
YeRaFuys+vvxK7VDG0ThhU2aPUeB2roVZFj/YVCBjKvQsZ9gLbfQAWQ+9Db3A5BsTA1cY9i3FpFm
M4SLt1dOGs/cpPMtrNb1LaUtudXRcXxiQtTGDNH8yO3TrisfrFuXgoisQ89XDjPoh6Hq/lJxHmSF
P3mfpmbrF6uUZobQHGcCRj3vghQ7SBMI/NMnXIFrg+yDta07JgquJc9b4JLEY6EjWsvrIqloZJbB
I3NMNwqRu42/XWB534COE8vSXe6bFBIim/UzXrFOh/shZaqt1xWAeHprVQSceZiIOU/aXp0JfZjn
Kx8tlw3N54IPpOCPW7pFf0PuTv76hQwMsyX8bHR07vdLdnrRafomLdNAfyUR0FO9dcuY7gu/N3n3
nZCSfhO9CyG4rCj/3pdVqIqmMpvD/0/klEv3iDapSyqna+A93LQLwqi1BLNifuHQ5Ib122F7dQOZ
TkdIsj0JTLcnHiVwJW40hhvzslJ6UmqS4qknba93+/ocxGQsDuRGFvsXG3TJ+i8/FRjjf0fKVj/m
CmFtVzqCOOnv84qIPGgZa6whvBjfFf95RhlsaRyekXi76rROts7WdnDwQGsPr9/gF5awhcj5HBvi
Tw769DGJFvdggElr+6DAai9cVLBXZH/mv4DRrIYOJ7bShyfd7Mb8p2Jd2DFmXc2VfpdG6wvwClo+
1d+rSrjBRLezyRvNVemb+vDZekbaEu3V3/Y3SJEjfadixhY+BUqddhvTJnhysairqUVJyeHEkOVK
bpE6Aiywe/rELt38ECRvO7CnSWqPp8CfNlLmlkP3UTzQkfr9is8dxD7rQAdJMJ+/UJCUEsIc+Nhg
glO+s8sG+hKbV6Q0WUx4y/H1YKSU8j93X3KMzh3RAL/MiaLY+nR8bhLZobcCO1ZZZgtY9uzdLHFE
L6OqJZleURwWjagFVtzTNi+Pth5Ihovwn1lUVaCk2WRMUs7CD/fK//5djw2gSzwnyILRQHVTyCyG
SqxKUYuQRDNo8bB2rxKTkOW+QuKIHr8hNlYxNTkYzi15Wwry/yOH1c58QRfCtVopBTgPmwUvkjqs
q22W56zadx5LvvGCLSdlIvX5fj5BlhbPl5Z5E2U66TZ9sdssE44SrKD9if3ZqNr3tski01rM1uTR
C0B6nN4iLyRPe2ek71yfhWY52n5EdEJr3qH2iGntTMOxfRUv2Sr8Urm5xDbL1PMVypN7UYm7bC3X
6FOXAFxEybyyQmacFMIGLvs53TpjKTbxMwQaeaXUm3PhmyCPsc8PgwczBFXVtpv0ZxDRPEjJ9BSl
yJ3WU5XewW09f05TxAW8q7MBUDd2v+ox7/9hT6AI/vVmrkGs1FGp4GG1s9PGHvLLU68n/M3fNrms
MA/HsWZyfx3y0DhBpdJcILN+yyIOfwYQXm/k7+QEf37O6veMkF99lGiiFDpWGMjYD9zpXqzglWcp
w2ewZG+wkl1aw3Q1Xar7fmrm8evd0TW5Hw1SijHlU3yq2FNljcc1i74UUSWncneWQnwirM/txkQ7
e1pmqJKVmduoJYO95Ai67EoEmWKtpc2S5OeShuSx7nnFILgJpjjSK5Z1PBW/OBRVRgEF3CgjB9JY
DbARslGiD/51OVhJKrqzduXS8pS6s9mLi4oOb9d39IomH43B4R+gCB15PbWcALg75Wxl4rQVBlyC
wfbpK+PuiK38HCL8jJXTYHZrhOJxBMNGAcChuJIu9axhJEdV4fSUMm+cqS5M4cQMV+k+5PngWV73
gniq72eH31TPh9+VsJBjQfg4t0+jObOrMlVzStyWe2riWwl1C+hbkMf0wMtOyHIZmdlg7xE4n9cS
CIwWB2OatvbYcPVTnOd96nc+u+ogiS681nCP+aSCuFrnd/GGvIywJKxvUCutWrUoJHjBOX7M2Irk
HT4TbqpEvdtoknCCdvdj76uIIpKnpqY3z7HZSKn7nBe6AXTbmT48RpNiZ90qs6hwbwzjWX5lhu+8
L1NAOKxlxX7u6f5URSBvNqU8pVIUF2NveMyIamI9P13IZwkNp+WrG+JPjfHL/369sj4NlydOQQJd
AQUKXPY/XtbR0Kv19U5L0MRDR499Sw0ThSomgPt2i4Dlx/pdcE81Jc5H8I951/fU7Dn297MTXj1v
J6mHOYR8tftyfeY6IO9luEaEp+sjrzjuAD1S62zv85L7b9v8CZntc3thh0V7ZVc/nto1mh64BzSX
xr9pXYHpWSxxeB1QEtOtx1QV/Bz83pXrICqEapV5bThIeI+t0O3qNWC+c3k2zU1XMwLtZYG9z4ik
B3tT9QFimA9nJUbfmj66NM1DAbEdSjXrTaVNrFzEtZGzD9bhwDX7zP0msfxcCn1EFY0Pz9tqPqrx
1hcP+Kvt7SkHvbcTc+aKCc4qhDge8xtDqHkRpenB7y/GMnUHV6OqW7KhT9PbkyvsD5sOuhcdRbPq
kL2Q4wqs6YTINLMbMJIqvemvMuF3XxXy3E1zlXisRpl5QVogxFP2Kcn7/oOy9viILWZEny/C+y7s
QhbwVIbbz7k37X8hlTcwNu5NZRsbPxI90VYaCVgBSkOJLe2WUPsoWN8lXR6wE6/0PJD4pNxy2SfA
H9YfITzPHSJXeVLDZ4Xs1dCcWPG/ncx6dzBEJRAqUZCb+ncJCunyW5uAkJn6TQWa/gCNK0t+vGSw
NY2UFfgPkV2+FFaQEume+1LT25pMjq/YKE9ur1yqnKG3/jSeDgX+T7Ymkbst0xYeRmG62ozPh8QB
j/R++pp05G+CfHN3RRSjguXXDTTb4+3a/UyRTqQ51hEtUk35zxD739bFzThp6d6qkBJgwYgqgnev
hLmpG7UZZcWdGSgCKGTJYMRfzuK8IXBWpr1c+krkfaxaQ4rn1vaVhPiunoZkwqG0BKDAGDvIRSRG
XCYH0THuKQIut6Sq6K4OAGirxHsqCUnvIZLif9h8kOnXzwdton9AviswZHuwhdub2cDwnlhZZYQp
97lnr3TiJAkB8LbjlxeFc87nQ0itOseziT+XccT3zm30/BflUfWv/b6I1Gl/NSwsaMyNSej4JS3A
qti1kZwuWLx9AE1nf6pcfoxDkLoRhM1HuqFTGGHMrXJ9D9PAyLyxgFNd9tT0SLKMICbZVOS5NuY1
F03z4XHxJdsvhpW19vEX24tlLnJPRnUrjQ4fD32IZD2dCApDlQI3JHIS41GnXvAUEXMEZbpjSINj
9PacA9dvWPo2khegP73IFYbV00bewXHGaKMpsGSS3DFtM+BVDFnWfLIaRxQs9YqWqYvupoPCpEdI
4R8qpOinvj8cXN2m04UOJVg7h2oBUn+4mKDJ0388xMCKSFh87hLGeaKaLzvMl6P5Py4wYMwHPvOI
OM2YALdiu0DLIM4NncCqjPDynL2HM32Puu4t3Bx4tZDuATgWt1xf8bA7fG8Yh1hSVMg2lZIbnI29
RU1X7mi1yA0+EYagCsyjS4USz5p/kzLIZHc/Dsn7a/1E9kCH5xOVG6MQoiY4Cj8Tu2SR5+bC/baR
WPUEReKWRKa3X7V/RG5YWQWjrovU1AnYMCTg5HIEJp/aGtNOLZ6B7sDazIlTtKmoI0J6GA+zeHAD
YHhHveH/BISLUnCl/vQPq9Jq4uMGFdMyNdu8nW/DH8pcIfwwkfSc5aWdFFMazCHkjNuR1WGK4UWw
JkzAoZCEuBHcGbSdMPrkRV7sQylaePPNVxwWschVTYWpmwXTDQiXo5BIgkzwZXq8Y0/7W93QOsRd
Aj4hRZuz9Q80Hua3QtnvvyVP4pEVOC23Sm2RuZRWSZhmbvSwC0FVHL5Wyqj3VtRshTh7Aj0WsEjD
JDKOhjAHXjeRBVYac5qZ18tuQfhpEjXof2nMzkD7D70PGjfnTWUeT2+1H3DVJjlBsgAv2T6As93N
bYkv0XZXd0DIUjZoUN9EweTUzJ1VJxkk91OHjI5XGyzY9wviFOahVP0mXdPq6zKHgr1q9AhPyKV6
UV7el2Ms3PtsFY1sdK8GSeZMYAZ4qYA6XbiHCOP07TOk83UkHW6gu5e1iiHeu0WmGKGXkhSWxugV
VDBcFENisLCvsndjs5cyTom4XiiNHzVKhZL6gc02mXw3UPxrw0OSgYLJdDqeqPuPS9OnITJTayhq
Xx/cFJDDooXazT5cbK4r6j19vO02ej7aF1/er2UfutN6fNaygWUUFJggbn12rdAznvbA27HWUQgH
7wWSceNYJB9qPLgUUsSmszZsUpse5XLdtyZ0SL6Z0H2UntoWEPSl4DCrl/OqUb5Mk7sD/viJS+L4
xYWWaxH7/Tx0tsVX4CzJ/UAtsK8EK+/IR2w4+wQHYE9dUVnfvg2wi5rJPm7OWhZ2tpcSTeNj0C1d
R/7E3cxtLZtIetCrw3tS5cSfRUwxv792OPbmJCNTA/kf5OfynXJQsdMhetIOTL/sJdRFVV5tjTcK
phmRontHMwgR0ydV++sZ4U+VcKi4vQMbsgfry7ObaILBjHHnZOzW+PrmJvfHgHRoAblrZS8eXONF
+gZVSfzc0iFoDXhqqDvtXeaRIOQRHNGZoFxszPn8Wiz8iPTLzKZmUS+LCY4n0KcY+RVw6me1lHue
1WK0Sc4pgtVxWY2xFrT7MEI7zxV5G6t38GGbxoxr78QWU7i2Lu0jhlXo5uPSr+7T8nuECnu9rZ+H
DMVcnJILYAU6r1eldFW2DoyhpbMnuJoUwsf97xoadyYFkc6VyjSQY8r/VLEVmtdhPakXFcVviby6
SdP2S3b9ThFe5yumI/Y/TCLMI1JzQIDLDZjUWxPzIFjN6itTmAEnMnjSkIGuCzVacn99udyG/Mso
+4r9mSchQW79VP+MhKTL0iDwOxVGcE0dv7tRZucO3Wi/U7YuTgzWps41upO+F0pG9Z+KGAVb87EQ
xNsBLFcJ66BQvtQWNuulHksrKUl+JjkxyYvsKTyusikTx7E7V/OvUn4p5vYDRcfPzQQLuHuOE5au
ZPm4djfwMusQv120OPumpqHmpdLTd4U6tObkkaYbozz/LK3TOzcd+wyepB4SGYTAw1fjqwPr1TcG
JmB9qpRp8x+ZTZef/vM4ZQca5l536CVUZKPMXa49tMk4RB6ozZwdyXHWnse2+HpDLyF6Hwc5EFyE
jQMpmhnULFu6GJ4hlfHmhImk4sn2x4cwzjdx1ivXHGgkC+97WY5uz9i8iB5Qs7Vjwxq2R+RBbTIh
qL/utEKrLtoixEchlIdXzZNpqEay3grCa6f9h94hsohkU2L6txq3J8qadCZ/X1/QBggJy9QRM02N
6mDAZAefEalqo7y0uU+O5VwDJTalBoBuShXzwhfApxBP46Te41IHHf+rUDm8bEglC+LNCtZHQR1H
OIXpyDvr6AznGkcWoAfj6xIesZMG+5Cn5YpqyfAyiWaovVUsCfL5K7ZFwApmJ+QDTK6yHIovAWbs
KsNI61vXy/C4S3AGJKV+M/jia3jmcopVQx83UKNnjdpR4vCpMmKy9btXwRCpdFBmUib8Ayy4z8WU
58Ii9zI+0neAWMuxrli7yfXQxn8WPKASA6EiG38dwrlCZbbd5PkzppkrHMrHmOBxAV16dTPRS6fa
K+9lk66A8aUl9KL6+VWVM4EPU/iAWVvfr6mR/CrHkAlTGy/e3UlAGYtB/W7sSxVJYzu3qqiNYDiL
Ix/SMdB75wX1b36gsHbzaq4/RGmipe9L8ccxGxxZdyaYx6L0fPxB0tmTDgnCxAau1/JghdR/1UfY
IGEB20F5wtMKefSR64CHSlWmYIDSmbT275QzKYs+umBfc5FqFLdZJrP+iVfPCMD/f5QRbnSE9vu3
mGfmpcHAsDUoIh4GUMO67asBl16CLJjMY09SIq2zA07aSD5qZaqiXQqOZlblw3X0eBYofuSBAfcm
Z0odXzRUxSVwxzJzRQdc9HkpQvaChxRDxKYHfqgtC0Rn7ZcN0/LfuSOPbtEMB6kTIwDhoLV0BHxo
4WUckUYvjDVdcd/0C+ZqsuMzFoxV8DmFHhTzUNYAQIjJvnBYPFVSkn4+r6vwPWMEP3tMrG3ssSiK
sslq4uWWFyyMUdw871rm84OUh40ttSK0i+dLju9oh7osZO/njd5qzGZBrEqU5o7f6WmXTXQjh7DI
2Ynu81r/AXHRSiRViLn2MRrAoxvg1ZXTaruQUIhXWdklrDsJkIyl/YhIvNdUaDZR5AOLDCQimQ1O
HzxbtcPLX/BwC+a5mp1qfyT/a4udMLGFovdi2SbL7/9us85XJZw33iDpDrFKmiU3ysXp6b185koK
dFB0A27naMoIoNRoq5brLI+REuoa5MvCqafKkeFlTMs3v+Di2vJh3SfxX34NO+ZiJ7J7eWM49QPf
+UeaEI7yd9OCov6jvu4A2ZlIocmObBbSDwTaYU6R1Eeeo66UysynnP4Jvh9x4XvnuQ6Oq/6JWWsv
vr76b8mGbTVdfzKJq6OinKfqSX7nfq6OaewCFMzFeJK7tV976XkyNB1n3d7TRcJNqJAj+vCqCVOP
hF+wpOzNWyXRVl+caQE7AqN4Z2JjnFxtF/NB/H0a3R6H20CXzCcERpqF2WtcmYOKWMS5HsvDjf1c
Z9I8jXuS6z98wQtlOvaXMogFqw75oumBO17jocZLZYYzXvQYYwFv1AgptiA1Yp25gHI5ClH+J12u
9+cRCVQIf0u2/0YQDtiDcN4Wki7UcnWML2+QWaXJKNpfC4CDvUybLpP2tW49R3pG+massSAbTmhG
LkitPc2IimcGjrkVg1qz0se1TA3Ud6K/Y7YlKv5RnN9nsT92N19fD1rELkM947bfIZQMvsu4NDad
Jcn0SYMqjlNN9yVpyqBZR1NWQAeqEpHmHpo6BwG2Wa0xFQMe05SBTBh/9rg+FVBr9lT7FeZe1z/V
N3U/zCfG6LbgwBMm5pDMMaQy06bhhPuCZAA39yXPrM/ltWfJXKY+BrsHAiOZXVMW0ByY0B9uzMTe
iaI7nSko5IW6zoVgH8DWZxzz2DUp+wbbByIYTSxnGQ4xS2CFz22OTGeSUrcOeRxDGK9Rwr31K6IG
AjMkHpSiWbQZa0aDtPns0wj+PcDCgtQwUWc9iTBhedvn2JhMlclSdy78b2zBcO3Lft7EU/36j9A1
w+pxLDG0/BnmX+YIFrSkuP2AGA6ihdHJqGKHnUzEJ1eL4LSNlgXfZApAlSVN0I47NI5zRUXXJGab
mKL9bcrd169tPGvLFEi9n0dlkYcA7vjuIptLOTSt69wf6M7W3vOwhkj30TjCg/i7/weLKU2tYad5
vg7dP8rk2u4mALYABdpkuxuF18NUiVZpeyDb63JGndCYfXENMddMaSqQDFLGepXBy71j5FmoogDy
4/xWmwyRxsZ1j8mPC/gjKSTUsOU1GrRBp3mrM7Jklwlav7+wI+F76nQUDVrD9a6Aen9fzVLymL47
ggwCSwaafL+GavlyCZsyPzx9NUFAsSfl/gP6djcIAQe+4/ItdFKVvPWZx/IhqxjiMQP3cpAaUtjl
oDPcbSYyBhFQ4P1jjK9fzBzmTyDzzVca+VlBhnsHoz5aFPlqxinlh1kiV/LBmea6K0KwcTmHq2Yr
CSOScJ3A06c09j/vipFtwBeGyViVjhyW82JPddlEGlbTlVzkP00acoq7/fz214t9ZFW8uW054/f4
DEFbcpNFmpPGwOYP4oGE0HUeMCZlYKZ+dEFHWMl+L0AhO8/XtQKCEC9l3XhA3KeRyOGiDO8vvU7V
Sv5SC5unGRqccwZikI5duBMzX8sjGjLc9loYhqBLNh9le0OgFylNjCok0pM51HXBjiXoVrfCqwJ4
PZUJYoICGPTobiv+wqFj+Gzf6O/hQdCe/ALO+kVtOsuq6zqAWmJcVHceJfz/VSDS524MIBQcKLIR
I1AUS+stDqQiPQw7n2l3lfoUmSIXmSCyclZ/DhkZY8PsmYrxmuwJaw8Sa9MLU/F7Zqh5b3wPeXuv
hwFF+dHrAHWqQvv9dpd/oecDfhIeC/bknHPTNHdNABKLT5SnsiUSutenDNQtHUUPnP+ObkIO1klW
jaS225ieH5gkgvlLZe0y/2t6zE1pDuy8Y+Il8Ee+rM6WM8QnUtf+0VVA982z0CDR8ea+mIBKJPSv
dYUMYnC4nYeLnKLuVvLO07kS9bI2kB5mQSIyaQOuoMxBNhT650layxz4tWV5hIpHhflfThSF2pjU
H6/YLZ10p+8ffrJOEIyQLvvGgzHoq8PDgZQ5QtdkzRCXefeNELYQn28upeqV2FHpDTDGxoAjZUGL
KrdDFFKlbzFOvhSo6926DDpyU7S4PrNK1S7d1envaXwkhlg+6hTKMfFqFTsMLThqzqCsXM68qaA7
DJNWYnBKqTUjf8WcnSpgFdNCJCaRodKuGsBKBv9T1EHyQ+IpciR4AkV7BvyHyIzJKmBuUzFRe2Cr
LQWVhAP8Zw6K9bIgrypGeItTDFpW55oZ/AuEuJhvseMA18dDsx8Z+LveM7hihd6rUIorTpT3RZ7n
FpPu1S/WFWQEZF6CVcKytHfKHICtORN85vPzPcysYPzCPn/XPP41n/UhrTIQQZ7AknIJHRDKmWKo
Z74mwMKRAXtHLFPZUexUm3nK4wSqXJARuhVMkE5KF52v43V9U6tIruYrWbLq7yw+uRIkU6q4vstD
TG9f5sLV1oVZexdeKalfWr82nCPnb7bE1JPp7bIGh6iNTtR+C7q2cBrqXEbHuIUbNc5ln1hNIamS
HKa5aOcWSpMyUFezXkbjdpXL/th1VwtbZ54uPCZrWjMNO1Qmb75a8CQL5tIIQCLPneJKr38veSTK
Uub2Eiq39rEdgtXVLakHgp0EXv9yeyxLCMroVyGkQUMvW4jZthoHpoEVDQUbnAgMiwIuvh4VVgQq
xg8es1oYWxK/5gq83WypUQ7H9qkmhgOL6636JxehQ/LWxaKlc+2tO6ROLVGr7Ae923HoCT8S6fSC
Cdr7QmFuvlOQIW3oRCRbKBqyg1FiXmV8pMTy7evNrUJIIMSv0NfshD7NKdQHH19O4wBm4gxjA8Nl
Pq6cvkHuLIKU8MKKuVoquyGlmPVLtK9OBh6e0/Wznprrfbmj8G/Om7bi2CyhtdB/yorypDRS7LRo
Cq04X+G2PPGZLqCW4bE1TSYHCDwNbbK91YmTiDiB1Mw8B3YAqBA3elJ1qB6P3RD+vavn5M3pW3dJ
QqCfeFaP8FLN06u2hXjjttNY/KE0VWvrt8wc5lm9WT4ySPh+kbQwz4KGieUNzLEDRI/P/bj69ajt
NQx9PUVOv+Yyv332SG+9/Vwn/znhvslpjnwlHuvY17Fy1sSQ2jAJg0EeL1pVr+vctiBwl+Jv2p+3
E1Jz0GSXafuDZd6yCB5pprelGziTT82+Zr1W+vdSbLN8of2c+26NA7b4TL1DrqqsUn9WtKiCVv2y
MGaPNOwvULpTxjbmvSlydHYQ/Bm+yGIbR6mGHoErdtN03wDYhCybFzMsqAk184MpBJmzZtptq+kI
7JhXl1Y3p+P16WqkX/Y/+xzjhRMWY7u4YkGJA28CCKIG78bMYm9AGLj4lIGGm1Wqg2LFELlK2EZ8
F3KHf5l4gb0UpbrQv6qTjiOa08ZmIRG/KZ8tVViUd8ohw8pV3iY6trOMWjyKkHngjF4LbJd/F1tG
cl7YtD7C+PF7O1oqSQCYtjUjPsrAyJRshY/UkgCGbhx+/sioPF86kNoNdNk4fbavtJVIJSebJ+SD
dcb0NSISmGs8hDXmtntikn+FITcqQ4qBwCjqJh1H2JP+ja/Em5nuR4AX1CYcZlBr72qeYMy+oX6P
ZNbynAxUTDw3psMn0lqNbDDQcD4DzIhND5zXKAyPKu3u8m/Me/xDlFxgCuqzCARlrX9OEKq/KoTI
NyYAAK6N2VH5r8pp7vKMU9OKBLHE3YhaksU3rGglA9EHo10N2inF+nR7NcgaNkKXSXsJNCDvr4r5
O1ubo1ZKN7rgZnkhR7dAHJqqEzQhdzfPkK+vawiaztLRIL8Q8GLo6LqNP5LseOFpZX7W2UWiulY1
5SdcoccHBuIrOUFDWDa2yICCbZ1BuRl4eRKpfwNMTOQHSdD0Djep0tUAvW1iBuS1IFNPCkeMLBgC
8pjJuLYT48HcNlmmGhYbo73ckm1XfG+TB4lpfePfT5ZLQ8JlK206cv87+NuPe8tKAdgAs4qBPeyi
jUv0MefKsWqc63jw01QcW/h/27uz/LlONxSu2ZOIfWLJeqjwjfILdHQhYx5nctuIlX9gKaFI2zR5
7BQyQhyed3IpOyQBIbMKl1JR+mNK2WLnIisPAsr3fGR0vVc09FMYCstpLou0x73fi4Bhu59NA5su
Hr6B4MWNO9fJk3lQusdj6UWReEY0D+XhgF9jJz9VqDsi0xcNhG/xgzUOHNhhxwhfC39SVgQmAmX9
XOjuEW6hwDTMQ2TQQBKSrItRGGtnYDSrNH7t1gnF7x/cXwUvgmfQFU96BlEhC7RcyJ2jbesOeP99
I/HdmvVvVE9uC7yaLtLkhCmqP3E+zAWdoPZIkmi4Q6T/tqRRKlnVHtrtRvgRiY8+dDXfd1MhzV91
btGvDCK7PS7F+nAPi2hwXxvRk+ZOzEDF4hGuYqg+WfNWpzQrB4DtT7FvToaem0odYAc3EuWRW9KA
0MzMmkeacyQ4u8IFdZxDMXKwSVGYNoa7hZa1UQblNl7PcRM64ZW5h9VBSOFMvAFCsZfy3u0CuSON
iKfi4YWf3nPSJrYz5r+4QP8xMBEJJbITiReWkGsNj1j9NMPE/zsatH3BAdGeNKnkJdFhxFW23/IF
kj6ax9FOKwZ3qsWLIZw59KL956lhIq+bHyioTzGCPW1DEU8Eq0LvgA7cQMRmSj/ZsONCKX3Z9W+S
yGIRtLigvBLHGWlAqnLV60PaKEx7ppZzPoZSkzNQVdxutMOAmbRB55Z1/D9/Isa7yKMnpPgVkryk
gZbT5+d0AVey0pWhys8u+mAKaloAoJI3U6tkRbmJWEHBUI+rGzMpK6/GAOyBjOZafcIpwYB6keoN
ntgc9F+iSdsDguYyRWr4k5nguuRWbSIn0xzbjjE/dRUO4KQS3nvtP/3rWF0YwPf5ksBAkHLP7uF3
TUHvw1SuDTB9cCUbgE4cjFoDz735eDe3YFaAZR3E4YuHrTJtFPqYfz9cayqDstjMu0xT9xnX/gWB
Jd+eX+BD7fqqvmueDQDdy7W4GRTypY6b0YdP8HfV/ZYxx+0oKPK/a/Q4V2Xzi4tEn9A6BvqodU4x
jfVKXCWaaVzvggK173bGj/mZL6Fy5UKsEzgE/QQyDurMKRoife1evCWdr9praXRIk5uBdebtBVZL
rF/fpNlAxfIDVeNYQQbw39CVv4YxGIGRMbjq3CySPehBN+cMsdVQ6z08UM0b6P+EKhIOV5YE5bFh
mFS0KvjK/qBrAwEU5cWKVmgljeXoN/U3NrIgs4UmV8xVoRPaqj+CiCeST4Q8LZHnZcaXKU9oXz0j
ovR+YOpwmwFr0hNEmwuwE7QPi/493fVitKoM+FCGmVFyBnViHkchn5UfYcE7BN548H3uU3YdBDiY
4QfNraeer9NWmPctYSlvkkrEHf10yWPVUtdd/5LqaMr8Lm51O4ZDam9YAVt22ZTwSdiKGQjSGRsS
zvAZ/F526Tid5J2gLaWX8e2yOY8g43avppMUw1FYOEu17p0Gx1lofI4RhDMPEqdB2SzLmg6uMYfY
Kk5ZIg/RJPqezkg2nz+XmzDahNjg/d4tuZd5YFV9mGRMTwTRyqVP3O+wOOphpHZXdQRnJ3JYuwv8
9/nbdqf+6M1nNFXb5dXBUwI0KSfWtAmKuUZXSuySHZ//tQBcaDQvBwyyhIeZipbdH8zyZP8NIPHv
cfUkLv6LmAhI+zr5i87QOjHMbax5KHgGgnWLbROx58yHVO6GmdXasY/EgVy3k6HHwzG1v20Yygea
pLl4ltFetFiTqKaDu3dms7UfcfsFSaqUL2l5fyM0IN/bSYOg2wqNZKXfbY0HB6BnfPlEozxXvql1
Q/DZxvDNrKT18iNocxrWR/q+hQ7miGHRb2H6UsWs03qdH2u5eg90OAgiwwCXREfW1CdgvGggRwIU
pepujhL1d5rQLRLuhKSfVpU06fh3Q/E7YblnOxfT5h+hT9PhokpBaVRGdOhi0pK+dmQkSim5SUaQ
8yDpStWTTdivmFfgAHT4Ca/txfA8wp7kCKhJHXOWbBPqh3pfaQlswh/uW+Jh9QJswZ0THamll2/c
Smu0Yi4AM449YDpC8+i1c63IL3pe0MnwZ37BJznGDJZ+bdyjYgqqQb70uuwb0CxtH2N5JHg4GxcC
IuHC9Vd2FWDSAWNQ1ZVzdM3WE19kIQCJAngvvA4a+b5BpG7tiQB3YMjjY8upSfRISpeUELfpmpsb
fI0vlZasO732rD7VxyYBZjohENNkiGgtSjzXymYGFU7jelLOXAmzs4mj35owJCtWI0GGu+ylXmyp
CnzZ2hpPpruTZLQ1WVjoXtgR1oPUUnSV8uUOfJwhJEs4/jFvsi5PktokGtaQMwlep1lTvsqbKlL+
DoMB9UvJfeP/SQLIBVksB+3b2lkHRReLpRs7/YDi/LOqSj4LdZ7qR2YmDCmd88uiHOH57DSf/XpU
R+x0WgkaWXgVwdVYvjyVDHrcS5ssCCM4OY3qNBJ/anmvbJVuKGfDM7yXszERjGXxdAW4ahY+UsLj
8HAhW17pGegh9GVlB5687Y5oNhx/H06RnCCIUf/+RpQN0NIZqwPrMqIut0fqOpeZW7EsXSOW1dUY
CCjEuI3YSgJFLZhOX0zG5C98JKJdGYfg1UvHyb+7DuMjf07/HERTEwYL4wgeb7pT50pIFhbeT/m1
n1UCOwIR9+ZheJWLc2+dPfZYkGYA+Expp28/1XzwJLZ0F6Pn5c1RRBh4FAi6jhCb2jltmSwxbhok
m0Ipdt2Be/Ur6OZ+m+KmJNOmY/xJIRKdvgF2+2jRFQFYAFrUMnefS/rPPHisDUAZbTh5P3d92Nx/
mPGf8lhQ5bn+arJ9Jh3zNSYSs0+q4aA0sOTRPSjo5AOffZBZDIZ99nbFpe27s22RihI2IBvUTYba
BQkFfTPSopRaB9MJsuPALAmTSKY5if+JrINCLCknckqV+xB3lW+38/PEvcG8/BVJWOQ8rO4pih/j
a3vqpF3E7ZxgtksaHzp5LpjW7hdqLp9M84wEoOYmA4ghoqQgB5zrod/df8JkdzCEd25lOZ2ZuisP
+1Qv5Fg+NGFSRdOncQOjrsKcfEphTehC6iQtvVyexDzYOlH07Xj3JrXyvNnvKFuEHa/DcxzEzpeu
893V3roU3EbJGX84KGNAxbzfqj1BDXfVEDB66of2WC9hCkh/Mt01niCCM5ArSkYDjaEHBvkBagYB
CNWaE8Mw1SRBK9AwEOtaj883mPRlItnXfMSzfkrX1KrpZTEQi7/1W80c8y2b3AUwkZhttzeeyq/3
M8JFNrjhMPWOX8YUbloWYKyfe/RQvd4CXw0nFjP4QlYZBH/xZZEYqqOVLbsRZrhy0ClwLz//KQMX
B5ZiLNQTUOAxtTGZ1y/O4BktFlnW0dD3BfHUeHq4BNKczSN1ucErUpnGg0kDNdWlqSZzBcskFNRJ
3Rg7CSeeqNJXEFb+/czqUA2LDyRTe5UL7Afw9oyG1VncLvo7qCC8e/Vk3eXLICYNpv1s/oy2ZOrF
YsFQPCKMa1wbKoZFwKggYFbANJbtrYjdr4v9h6T9KRTlSx+EFTxWNggYOSXMy+8KSvwolafiIp4Z
EldbHcnQ5VkuBjSdgsU1PwEAQEuFAieXUdhuSd2wN6EMh0fEFzDDNLlLTpwYUFv0OxswZXK8cMo7
wSDYYFNYhcMGhF4Xh9UcjUzK6vkoO4fQ1FikzRwiT7jhRUP3DAjfGyh+FkSpjbdson5+XtAFZnci
kZqR9UHMiLJfRYmpP9h9JBmUEoKkTuffNKAkL5WGeMGvBCy/5wiyTE9gUzcVC+in1sZl/bre0hm5
AOVUzu7EWQuEpQlx6TD431H3QwbyzTrfiQm6xoj1tZw4z8PxU2B5R7rYadYW8C2/t7xF/efcH2ux
fKAN7usKLVrOGH1GAIFYxMLcwAsmJzGs5X/HccxzqcAFizFuZFTxOMSjFAlfSASrzHOqUEIEygJj
cnjBbQnm8R7m3DZVnumll1fj6SVA1RyfNmR2McBH5tynujX5tmaBnrm6yLNrMcLmEFZ4cKyZ3ygy
HhbQMdoa2wBH3PWqOnrFnZartggOT3aIkEAMIA1kuOf3eWPKY3RBCwjUYWJdS7h0sBWeAkiBoQtC
lH88AprDp76esmotM4BQ+x1yFMhxj/JN0vySNHO+eHHcDRDhrzIxQKt2ntRDQuNb7NHE7EtiFWDE
HD6SWgHnHXofX5NDGl6P7YDl7H0XtZp6tBvwK50nz5LfdFKxiEFuIAt0N5U5rRzVbPEIocAYqza9
Dtn+vCsFNvhzWrSTehsfVdBHjVGfX+7xEHG+QqDG61Q01h0JfM7PF+tQpZTqq6tLjBG2qBoms1Cr
jO/Hl+L/+LtiPT4GyiM/C6OL5oeL0HF3VbI1vGgscsqmSaqcBACuMWl/q8wSHKGIASnbb2PBP5TG
30BsIwIN4xo4UnSsRZK2iTRLCrSnmVpZZzXevrSk702sm0QW2J9KEARfq2+dIn2dToZFGDodf55g
889mjqF+zrkYlkaDRgO9t3rMyHbMzRjueTXyAXyxr2yBYzvE7hM3cESPUPrB4Mp3eQFBvj4GOuvL
rY9tLpKRYTCoUeT5xg7/8YXoLbcMXGsPcKFaWmnBfWdZ41PJjiBR47kmYQ+xCi8WRDBZMTYOqxFw
8oZf+3TkLI6k741lVevSw3IWMKgtMpLGrsnTs/C9VU0jkfA2zdMAQVs1YQSId9Uh4+XHQIRd+ymj
riMcsVC2SCbIH+Qmb8+6wOUD6bnfajVmOmcKHN2QhdyUEnrl7IhT2zoyt0O7eJU7epbHZxZPQAT5
1PcoWpcGe0TjMa6335DnDchSRNwQaFrZ9gbTIDlB03BM8TZCcvZtmuOYrxTzM3PNhaVawnPhNyfj
59wn17rVLEpRPa6yJYaqulUNgt5QfR17D4kcbf7oj3DNbTGU5PhmDSMUtLr9sQX2whFNmVtBnZXT
BYkPmTfOPSzZYVV2Y1GxnkwbvfbTo2TlVoVywttkw+CeWDyKPpI4eNkWRAHe91nx2oE9ul3diWt2
aq3bGbp17JJTqNiaNIAuXkpkkG19jZVAzk1pU9RzbaJ+k5vxp5WOqvaE+z2zirf9P3xtheKHgK4S
H3xSY9u9AP2s9DdfFtKZeJJihXp7xbde5KymEMK5F87qSLwldQsIdfySVc3L0iBiSDYwR0Dg8iQh
hL6vIqoEJTvFt0MpNrDUmcFj3N+1W9ebpScqtr1Yja88eLEVXaimIs+IREeF2bUxQjjdpuS/kzaN
Fck7THZ1bTOmjP0Hwd4V+2O7LnfmXUqBlu7giNreoVphlEbz4bzKK+tr+JbvWkcL3HUGyiJwXwtk
5XKHMP7PWT+QeZZfNyKhIX0w38K3vQS1aAdVKpTHqYkwkRhaDtAQl1rzow2p9pklKqkP1sKd+btG
dHzc4cYuTVcBDWmV+Ihc+17UgCgo1ozwmGBje5TLDXvPUzXFDkumVnj8MJr64mderJJuOTtBvOwS
azd4uHKiLTaRBjmw+eV6baAgQ62TAMI/YB9AAUiuJyiuzleD1rbv+/c7VxmzS5mtJ1BBhuLeUT2x
eOaMtsTNK2D46CA/bi+OR6V62jyFDu4Qwg1ahWkK8w6fr5tWZATmY5Lgd0kzVbyvxNkrBMDUJI1P
/XfG97G1ze2J0KEg1KaX8ZkvQ8xuFXS6sN9giLrGvglILluNgLzXNZRKXsdeFASLeIvO5uRPQlYe
Xwgi+WozQrtrdKxid9NNpcuzaqM8zL/POL4DHtdAOSfhtFrFZQlIXoGJQW/CMNM5VWkPHPnkKhVV
PnSfnVqJdsLQ5S7MPZXjlDpg87cOAvGEqKlBxE4fjXgroOCj0dAJNTzdGn6qlsD+UPxUDzi7rOGb
vKDhKlh418wVWYaD3po1bnYkfOeHytNBegDCeeHI9u383uThCtFz70XTAdRnacjlndwGjuMEWw0z
8v121dbIPqxPNfr7fLJwWR1jHpBbhKDEaRKe8yfRBqpd7rPye1b2IqluJFVkT1qfmJB/l3atkQZd
m9pPU2cVqGvQ2xClFM9XYtgNOjseDv2DjVRg6XdnfU+dEGC9CBsKqQeRVYsBwGEIxfW8SsIqkhut
r6yI6AVGEERVY5xvlZyL2uS8YXSUGZcriaUTGWA+9wt11iEMVNav4yrvrnZbaf28z6nrCHCYtMp6
RRRr+YjmCq/nfykX6MBx8Q/gIWEuPCfTzLDfbQhsglqNsuDpWC9jTjf8y+DJ340Kjn8/chgc12Kv
8Vk6ukKwjTbmMTs1567trpziQwU8iviLvaJhLMBUz1r2jrPcSN1yKA/M5RGmffDkLWyz0R7EHKCA
J/sOvNhECw59hmX88wmRaUINiT0+BZkP4zR5NUFaD1Vy1f0e7spzp92/xhEi9k8dHgAB5/vG/oW5
1QcLe/PLFRpTZRoTq6EprJN3Ua421hwLAsd5bgColUZDmGgMBeXZENJX7w6KRXcCsd1ssZa1n5hF
EGUPPwudgviHsP8yz8mdpj9A7ZV7/NmWcYVdD/FE372l5qs5iVME4O+E7JO1xYyUuspC9KlUI8Gw
Sq/3rN1kunrZD+Kp+U0Bn7Tycq1Sl9l8obNa8jzBzifYg7OwzTOpCH0RZmyi3fx7CGu1xBjKa45s
8wbOG1vfLbtE8ksNV0sp/FS3a1rKqZeYpWfLgIDK1W+YH4ZXgYaKoUi/lhijuZbHs4YTsZ6R1mTn
fR5SMFR/4C1+GxMf8DMgLrk1jGWL/Q7h+jlWqHdp5f4v7y//Kk/kHkCQl/bWRIxHIlj+IDr7IlQL
C6Ora1JYrXj0Ff5y/kaZJkKE/GH9PQCRsdeb1yLZVoE0gg5OjM8MBHNzXJP64/eVGVd7Kh2sr0Is
lh9Uc2g/Gltc55Ede9IROPzKccmdDUr+9tarhpOQk5gsLvxa+oHhzqFCo39pjBVzSHQyUmtWxXzo
YagLFI5zT1Va3UB8nodYvjL7jqjopHOzSEQnZrSM5zOu/+/XmuXypk5OC+wkzZlCVdFc7pqIvCff
cWP17F+2hrl8byr4GHlo5HVklB5tOtXzygXmOxXkJIExIVHKRORNSN3Ert/njpUVlR9Ksk5g1hWY
aIbbO1mE5fZHZYuQTcyO25hs5SAMMU7niBmt2qdQMwHUUdp5k4pbQG21zBnlJRVLzuOX5boutCFU
2uIykvsTSYzkFpDakEvuwKAZMmFIZc4z2Sjs4ezvaNV4QcqwA1rriWbKNuCvrNLV92GMriyerKsJ
602K+emt/6GKN951oNgeEAIs5uGP8s69tNbqWRuGp/jbOo468n9Td7LT0Vsp36241WSM2xJ97xdT
udwxOFUHjHFnJaH75T0Er0DeAjiil8dv63VogOMt2R+ngaRkEVKX1buoINu2iTXUvsU88ezxlMnx
c/GF8cgk093g/Goci63m0PhDhy2DFlTJV/Z0WbBGfPLxeBXKtd2giwNJxFqRANgU1410CKzahakw
n3Zb0+R74fNAbYH2zu8qwZRylmKeIwKRZByrz/jPfyA9g5STw9B4xetA8OuytkNvkBRGfORV6buS
WeEKuQHG8btSrttutJs19qprVeIoWnWVZBvER9JrrAiaH365YzboLkuwPH01qiXJ4V89cXeGXvUo
7YPOMw6b/p5K/mv1Ub2KpVhVQfInKLtlX95AXE90n1/4dSMRXPsh8/ocylkjx6BloFi1mhTHR/u7
A9AeBH2P4fzMKWHib0XSKea1YR41ecFdhZ1lG0YtHhQkHgGtYqhJYeAPk+Y4Yy/L5XYWj5xlMeY/
zdOe3pzOOnH+rWXHT+Tkbv2HI8tuH8Tq9Wo64zYimXgUQgvyqNu/l0gC2lGc2x/FtWryHHCakSY4
HzL1MBb5yFFGIDhSYuJ5JcpGxqq11I6JNqut/sxjnKyBImZFk1Gh11XV6hs1ONyXID+wSLObJamL
mMidhNYaeEQHBxZCt96mw6+2UCckB9E4XHQjsr/coFUM1+Fg78E5bOVf+fCOPWk9sR7AEf9dOCl8
45x1Q5e+H1jDEjiGDpqclkgWhjDlsDGZYWawBmbLxM+mE5VtjZ1ySjYWdbo+nMQ/85Lf+m2pAn57
WXisA/PBNXwPoQ7x0ixDH5lFF1O6szGuB9gvhLOjJyxrsb662KcWgOceqFr8R24CYL32v2nmlEsf
fzNu2RJTCzTg3NiVMRFTUbsfMqQqKUxkQpvQEetanGOItyBxMHUQS2POeWLc7nGPEtMZ4wemENYu
eiYNe77Djws3I1kak96AvSd2nlr7iedNy/HFGvgT2kIomjoCy+fUJkFcbb5Iqba5TYWO2sksiwEY
pTzx99yyIEhX9W2wYXU9Zgzk6MUwfQOGq2C7URgvauenTivII+rWZHcERvsu7Lc/GaZ8PSsLmOZZ
12CxvVsc+G5M4h64vehfPNK/MIxlbxMDeRFgCoTqqE7qaqCWm27VkllWGZmPYX1xpU4tb8xIUOAI
psgxu6CQ5Vph8vYAf4iOVE/UA4updlq/Vd8qJrROXFd2LuNvP8Fh+lyNiPnayMco6uLF9Zg+2hpI
BrYG+XrQ3Q+GHZJqrLESMVQX2PdZUWN8hwqOB4u7F7NzRSplMMnF46VHUd6cnZGqRbqh7CePiCDu
zS4bUFnEHj4rm28zPMTkqdY7DuEyggPVR2uFldLAO7SFzOWvYvTsPWwipRiuXy/vxOAhZehuwU+A
qEPki0XimgA63zC2Y8z9rYp/LZEQR/ykhwN1RMrAFm8Ylo9wOH3re2HdCZbbMUh3mTYbFoSGPksT
9dVU4IzdU/bQvGl5a/LVIn9P76Fahzi/zzHcYh0s2yTuvqaW4CyT4FP/+udMf9M9mEnOpt085FOo
hBEVjVknZ3Cv2pDbwHV1XfDx7My90b7FfUTAG4qP19zKSW7ph18YkoE3jHbaIsYx+6Oa7UT2FUBm
Vos0fQYByxmFNzLhQhLgDPGYgGbwS3zXiSrb+Yy6+aqXCQc7EI49IGlrJBpIpOlu276hKuYPArzy
5hXNIIouB8ePWMhOf8sehmF001efDnZPvYkc1pgjOUmHrk6hAUMrL8rT/bOC6hvtUhVnsYqE/U3s
R7V3kTHqEIbx0RqfV0m0C0aZatCAZoO9lWBZ1+FMq9fj/tL1X1pyXW6TfMcGmdPlFbNBPTHO874Y
shmRfgp3/XEpbzUyuzmsgXjsgQ0uYwGJHrAiR1zYIKb1Lh4RTdXHwLsJ64M+B6dVkNW/JBFKa6tF
6G6I5Yy1lBMpQAaqpDEFd7IxUkfL6lWMFTz3Z4JgtAmIXnaD4g49WDG+2ak10oB1xnVk9JZgizsX
jGBVQKFS5Yci2uQJkSIe9eMIZwtOHo7ROuwmPAFQU9paoazwH5tDT3lLGKc2ALJBJQDzuGKQvGoS
V/Rx2VPN/tw1xTg9PUtkfyaj6Njq1ENOfdQ9zHvNSCivJc0tmScRLGYrhxAwjfalA6g/F/buSz1X
d5383nEluByaCsem9yy1mlyct0rEEKxXlrcH0dNmkR3soWVKmWM7M+jw7wwelS1zKX2xOcis1er6
Sir75wDEuz2YNIRjAhF6cphyCXCgeGSpDzmG5TbCLT18AhvnO9R3kI4PE1lio3rEafPIuzsGRcW+
GmBg2h9RQKBKPMuafnohwZpbFgb6DZP1y4iznf7XQaGHK3YeJLPg4Yye0GzXTmV5dX20X+2a3vxk
7S9aF32V2n5uCJVKEza/NsYQMKdCO3WIJByTzOYdOLvrUydgEldYq27kCJ7oe+OkR2mOcf92mUBQ
ZQSjwY4Arrs3vYpubnpKMm7i0bor6G0Cm8q6O/yE9+1nNg7s1e/BNhi4hbdpjB2MrWcP4pXEGhAC
wWUCLhUsJc35ngNYSvn2mW3cIxFz3T7dM5emOiL2G4Mtj6dwg5ruF7LLcRT2/KyAsThhv5Q/m9Ic
FtHsJN2K3EHThM/6iD1vF/xAZgJQNa8cCdhY6HnKiG+GNHhqb7n+veFQw0E3ume0XLXGYBSOZqG1
9u/FtY/CXtOD1PdAFGpqUy/cK6uRFHg6kgYc5WBCqVJFbou7KJESdutFMcbzamS7+mQW/lpaWjhF
5a89CO1UGnVjMsnkr+n49zcaUOXafr0iPvrKFlmeeE/YKyo4i9ZOTR+zlC/kWtAYKsafXGHZwUl2
oI0WYahhzTx71CGMStzkxTNcIQ1c8eMKoVqVmFQNSq6+g5IlQUs9QuuJVq9w0sWkpibb0Rrpis0D
0uIOLz1VTG236ywpyMXTfDuTioRM0aD0FVGVyVE6BLI6prpfRArrZWjAv/zc3uwfVIyK843JzjBG
CrJvl/ye8b7/RP7CjgG5V/f1JFHCyfB4Iq5650LDvLGk952i8NYs8ijgjznQw5GNYZs02LPusB7h
i4ccfVSVEpxjsSC2I4I9ngDElMch8zGglKGreEWpeWSoJmnAL2VoDE27OgvJmE6YbTjyTKdtWyS7
nocsMzDLtBGJNbpWSBdgSE/YWjSTVOwuKmh9ei3UmRHjaIDtZdjYhwJKsVmTjF0iUfHS0vPDAMBT
5iCf29Ne2UMX0ht02Urlq+nDBvTK5e2Rn2KM3jJKEyDWoFtyyhPH2n3vIUT3Lffqb5L9UFYx9Qt6
H4wySnR0KNds2wAx7Po5EUjVehdDhX7Unfy4BFNB53Ow8JZ45+zUMabM2udLoH77B/f73xxzDVSA
A4DHxY46I+fUzVaYyi3YmId/UvgNzHID1D72mxTcDNRzrsUpQ+u0hrLDCKsdZP1voNROSLCdcvxY
KwxGCIK/LfSybFiGkGujKqVfJwRCR9xvil7T0TUDbI2FtgK0PsidQRBxYOtTCoZP3jR/fonzBmxE
5nMQmC0ftGoysZdWDI32spPJV476zp9o6uk8+COFPBSR/kF3R+slBdlSBSg2z3krDSRkZR0QpPyc
mAXzOM4sLfHzveDqSxJ461H8W76FcJrZXJN8pe2v+ji1JCraSluebUPGNTKR5/NQTvDJ9YwTTOVU
/g/IoA2JCJumRqmA4MrJq7fwWi+N+VPcN7Zpi48VXaSEbm8nBd7YOC8jILBP+ZafaOOZMHTsrAtA
Zpa7tUaYM3UOEhu4+096H4zoFKaMrMdZOrrsEhYlOdGSVTEI2uNbgu9Ff3PMmhzCDiVCm34yH4di
T1Xq6H4ZNMZe9LnykDZPfzORmPFwz0Ory6uyEk/RpeyJUx7q74c8jYNejqWgTklNDnUC+o1oG0Oo
1ua1h4zYTOkgYTHk3oPdQTK4ajBAuXpADJo0qzYIm7IE0YEXwW1KHMSFAEaMjoYeTrA9h4VzFQiN
iHDsB0PDgbKVyrGdbd0oF4tXWzetvLRKjGz7QVUtuf2djED/+BK3J3hKsEb8AKo2tDa1J5+3oFF3
bNnEQOExYRIG08sEOM+l8NYpkCKKR6thfyp35RIYobr1kaioBKrfdv6E3hXXpeYFM/YrhTIJxkKq
KnA8b1P8YaGNIJ6kFNxiWELu0b28CWad6YVjI9sJ7ugSDqv01gZeLhsGN1mk9XO6TthOrku4Rkql
3MqhQVCLNNsPfL9aM9Mnt90mqmdPL+nCutnMdL34AU8vCM0ZPrPGYSa09Qi1/Y1BqpdKtxsi6eeK
iH1SEW0zuE8hE44+ckxKQR1q0lYuL+GvGrsyW6GCzZDpX8jWVxDx9CfNQuN/hkWtitNo2A3Pwo89
k4Z8CEvJXj1UoCho3HE950ZRYXqXD2sxcCvM548ZzQbiwOo+ekUA2VWK5IhAWrkJuMl71YTU7PQp
Wtvsiul+yzbIUyD/u5/j+Ui6bnlAcHCyNBKKN3kSozHcT6fayuXPAr4l3Uy8R223Ue0NziywE0hv
TWulRYKF7dIbWl7HJ0p747GELLjvQNcefQgzh/YuKjvfHttGdV5GBMowjw2+6X9BQXJfSY9CJf+C
dFvRtKYmvFtFTn5EaonfNtS+ANaunBwtiG46Jl8ru8XLvvwLQ+v6qUGLPb4uddIDHhmOdRQkHmL8
EhqCITbmZckUuphSaieLtpw+JrmzZA28Sfn0BrJrC4S/cGfgytMrSTEdEx6gf4vuClNmIk254iW3
6buHA+hbSVqfmgJMKrsh/Cla7oLSPYEJDo55BkBl3K3ZazujmWNbaNAar5iQUUFVaJnskeFrt1Sh
qicIkR5H0Wy9NhS1/OD+hf0AqJIokaH5j9Ae8G6EX9Ltrl5ZGeQZriEa0uPmrzyGTdpk1hPgTjZ0
fB9FV//MZpHlCp6SZmS3oRFRhTAfvz9M8mPe+8Vka+2m/GSeWz0Y2HEdBj+zfy3ZCDNLv6z9vkAq
CqD+81Tdt6viImtCyn4J3vd1BK7gt9SNBCsXhvTrInvsdgG77OSj8BkcKEAQ0NPlSY44CSqpLIJZ
sKHEcwgDP73pKNQbSMcN9mJeU0diVrjOaQvc5EbCa17upkCAnvmMZH3Umlgo19K39HnPhkmTTcgv
4go2tnMHXmEpWehIBPl1oAxvNnr45mur1DmDFWBUg21WRWPVh3kUyMvttSWFbp3b0PUPKpn6tZT1
wviXKEd39eLq3LcWZd5xXimplbGpDbVzjYo4x0eB58hvZ/NzzIjyFuOVKWjl//sXkCIZoh8mEeSp
kzE1NCFj8SHlOkHMvZydU5YUntc0/EymWV7ETKDDL15hitd6ghOdBRS2n27L2KaDwOjo/trvrVzp
3RvL0hcPcf0uKSR6UXYilVwCPMCd2KegYIpW+b8So/S1kmanUQqynJ6MUgfwlNNiUCekD/cJ+6/X
qIj4wgDTV0xiorMp5LQWE2bOGOIuWm7W41yTCd+ZYMGWDa9NTj/D9Ttfw4rtoAcBe31Dnlq7EFae
pDPbbzw63QGf5/LC2V8C2M6AGtszGDMHJ7wH7u0GIVjdPFhvyoJ6efQsRpVPI553CXAMBZ/M+fSV
CHElSDBYvFyqJDxtignFBMZrhU5jOf/RA/kx5y9LHl9xLRC0Dhre3J+J5wHcBo/Zb7KOqeEBR0DB
pHGISMyVvD3wj+KsBO15aSwhecs/BgNeHvs9q1grHxxWgZw16RjvxIGOF6A0u6ytN8cbG6WdUG7m
zcQlnfvPO8ywzuldC0vw7YvCp9rq/kl4QLPfXJ1cmKhXqf6QhWgykNZ9Q3W4WQwEQ4s3OyE+w1Xg
NFwEfDsFCqCcRV9ifgaIkDDfYN1SAtk9i7QF/SxeynBlej416427iMx9mjOcEKMDnvJeBEKpFAzU
F4pxvs+xwain1JU1bcM7g6yN1SWLC5Lqmv8cQlywZJHvgL5j3QkW/HU0PSLhwfJ914xUo97LDeMT
sJJcwNYXnolfXdY8K6cxIHSPU9TYQMLx3xO2JKBT9e+WkhW6c8OqMFpZeWWpfGzEhpJxbqJLKiHK
Yf1sETptfQOA5hdlkI/CcNaa7h6eknMeEbrhxIsvPXxMBznjDnl5sbXZA/CI5+eWKDSRhKcFNTh5
Te0MlgllyDtIvpVWRSKYiMBiX7hSkFe+aIpk3is1hPaJjQ7S2BM57YhIq2Y+J34oJ2ZMZgbNwst1
S4B+SmaNczSNKp+tYrI4Op0V8fWgXhZQHvzy5wINfsAoH4Wcs8lKM6FtEQ/41uS6akxei2WDlEoU
vHPf4AIVX3QcmeTM13HSKIIYoSi6lI0zCkMoYIjP2ly+xtJq4dsxpKm+BLQBPKh3sAweCjnigsYP
Ln5xZaa5L8O4DiZa/t/28EOZH71fagDXo+9Xw6tmaUtT87us7ZYzSmwPV6xQny/CRnnBrSYs92C5
Ye0EFJ1UTmohtzFKgAeujbE9TxwYV+OGE/M3awaouWjgDjfUD5vUk1yDta0TiYLw/6dcLQq1T7Ee
6FgDDRlgAY0YQtcqiiMicrvBB8k3ZBMkOBytPiByiN057WCRko2Xm8JbTKRbVwJHi53ubU9lGAEr
IMmQZxEzOxiBcaShtVPLlZpnBhgsV6uf5v4htbfAGzJvhDlXdNJszBjGrHiajcuhyed7TuHa2f9y
1dHSU0ZiuZRnXGSRosYi0apHcz0Xq5VQfbD8wa446NshFOEd2TiJHsXrMhM64Ng8WbAEyFBSdEeU
ogI/+y5T+XojzNEJk5IahO88SPTMGyFWrBHh68jD/dKcNinMDJ2jF4QfqocVCQ99X39tCAvfP1/L
dDADuVYTw09QfL6FYEzhWvkuZLr1OSq7eu9rbQTYvufL+5o4/LRDT4iMSGqo3nkKZHTN8JyDgRhj
28HWIo8QIrhP91V79mmsXN/xe7js93cqOB3f/wpe3ipuyMapfFnF7r13whykQo8YZW2rxJXe220P
P/yyo8HFENhmwuCWm71e5wPrLe7Rfcea2KJJnzDSSFRVcd9KD/Pn5i4JkpOxORv0WHJ305PetXcc
tzneToWrdQ+atkQqTf0aBbfIyvEgjkDNLd5KaKychZCpHgZp+Oh0ThGnf9CguXPPt+mBX4/R2Nsk
D1v1UeKtiGHHXlb8YhjxacHhL1ugiMgI0TLWmBok8SwLUD94k0ZKulHex+y9nF1MIK1J+nQ9r6pr
Fva/EPnV+x2jg/qdY5vqLT5YC0Ov06SqhdFRljpv7CUPUS4nIGqlsmdpAPiN4fS4eoKOrIkr0Mad
moCgvwAIPFfUO9R5ORYuM0rHUBJy8F6HS7g+rJhUy7vGXDmtRJ1ekInGxOzccKD/k8wZLx763QQP
HEuxV2NSRuquPZqriIe511+IoIOSIakSmsfEtxqEvlx7dnVl3v8PYEjQ8qBky+RStbaLhbx+zETb
FN6m96n4dw3JAUMJAMS8SQ2y6yw7vX0dWUCczTijO8l50v/0zOfe4yC34Q11EibFvdX+O2fywvWY
56xINJJhKlsIcCXVe0OYHMP5OdHQRXudpRpt0BXBmWFv2Z/AD5mnnKJ4mOu0jFke7jRD7difH0Fz
1lneSDP2etNCWr7tppZAfv9P5BC3dJZ3TwmCAskfZcu5ivbC9sbw0y3Qm9bd+RiJ4CW0n2/A7bro
XBLKm96Am0j1AXDkCbQNQsC4NG4bnxqkIiW614sQMO0CQrmbj+2QHRjFPmTUSI4Ne/BndEZlMfJ3
lg6gpn+CNMngUUxOyh+KzSx4CH4EI7NtgsLc3Ofk4/s2PniSLdj1UfA2KmRcDMFKQi2jRL80ja34
+LCwa+G1XJO+x22jTNPw3D2K0QqK/wvzv6u7CLhbrMjHN5wPGMSiMUxMamgHz/ci2hc2G+sZy7a+
3qrzJb5yKOLPOpo2HgwQi8l7HEIw6EoJj4Im9OmyiUBXvXoi6pfioj7QqWt2vBWWrZyAwOlg+6oE
eIcEIS94QgOdSAt3IrPGL4jhqQl1gCwD5Ekj7urIfPvvMjmIQs6Q0fL9kjVyvKAje1Dw4Gdl775M
4ZigK+mqXe5kPpsmaCH6LU5QDHdGTa1ZYH9MpBaJvneTkalGAmENKZEvkFwHE2dYoseBOEHn5Tbv
KGC+b21bd0z/gB/By3JxnTVVZp8vNGH8vmMlKaA9XeCl09c1e0mFYDfEWYNmJQzmBk3ZOsOrqJMx
dsstVlcimtiATCgD3EEWM4BkKzSG41VUhFTJBEnsEihFg35WgffeZz81dUdkJbF2Cj94Zm65fvjj
dFd88vv4lxS+3qsY3IdD7CniqVtQBepPGIFxGP8+w1q51915Fge9QaCKF/eXxWHdYEQ3XFc6t9Ml
6MuvEc/IYva5naM5QObcw01MQgBoo97buzVMntYGqP01IRAXs3/b4mx5INb1shP/CHqKSNveZ9Fx
jECsDAY3NzR/0ygLNtlaVv/CPNyRgQbSLh64eeu0hf+unVfII7Q/qT89RNScp2S8A/R+KqfhYbWJ
HNBp/hma1oY3kxIvRXOuYmjZyKjIMEOr94JDhhVpLaEgOF4s+oZ98tbu7p42Jm2gSFdcgyPMsa44
MIBiz6KKFq+iSzhMoHK04ADgs2tdQu3NHviRdG1LAU6I1efqO5Z+HzHbGcJwBEL+L6SdBmmIlWEz
0mAy/8ASYB8DJ3Zh2lxQbxd/4RRQimMqtEJuqQ84oYnvY4FntE/GwZj9Fjq+kgihNcrqQN+7vhg+
EtCQJ004VZCURrF33TW0Nkf7NBPkBpxDIe3+cmPBvTUNxwu19iweuNOUTAAD6scipmD8xDLAiA72
I2yZAQZsLa2tyP9OgabOcHh6F2EH/PldQ0I/ESDqk75juwrZKe7R2x8TEgx4lSllAq7Q9lEORISJ
zINXG8CEIuD9ypqhAK9s6h7OWISrHwYOtQWK+iEMqfmykm5vkJXZxDnBcljOA7x6AIHCcifqUDLs
R9EuG/1JNeL+pUa804XVOSfQw0AgXQgIE5dZbnK6icm9YGzml77svuDoLLEzsfcdbFAZCUo3Si3J
+R+gZZg1Hb6+5SRy4c879pNWUXFXS93bZD0H/P918zX9SHAenGiBEe42LXWGLMdrv+1E6ju3V90G
K+Hhk2Au2z28HPkYkrF9lh6pcZKjEbzZr0YhxWxbCuYacJO+9ZlWM6tdY7EbToxmPyz3mJBnCuTU
TVjgXnD0J7CMkMXGB9QyHykQ0to3ZuyKpgyrPq5D7A+8IYdjk4aunDP4xS2zsoGtqqj+jSmbzyIC
+eZpkam0F65gxMKzZjTvm9E7X/QJrMk/+BsmAqZltxgtP6efCsw8nfAilikVMQLHwEffd3rZbhMM
40jYAy40TFH4Mz8tj/0iX2d17FcBxFn4cBn2ayV1oGKdjtlowp8wW/SxoGrIcxvuK6OTka4IkrAM
tywb/ccVEr9Z1BYYscYpCQRpxBClMjGl5Z3Q1rPSeQ5hi/6Z67J+tlU2K+tgeGKGkHbeK3+Z/fLm
ZmCgwH7btk1e1Ufo2U/5+aDfCX7yuMPqCKvccYV/kECvnaMdaR3012wky1jI4RSDuW73jtYDTPRD
4IA+F8IPeuTz0U2oHxT/KKq1B8YHbX85xihQ8qt3HGTQKkpUwGwjn/eXv09foAMoEfUEfJLn0STr
5cHbII/toNP63U9/JBdsC2zO8MwAAnfcfUTFgojW1GNcQ71Sy2p663dAIEC1GdsMb4T52kqIxrEu
ecLGheLiiRtuWQ7h6xly7YLq7Lv/DHOfAZrOXmauzg0zvrk0jur7smpn3MIH3ZXIwLoKUgm9hOws
DQQ8BzXXblLfm3hDt55L48uJflBqxIAdMR+6it0cfAQLg1GBzPAIGM9EvqPB5Nx25CbRd9Yip6BP
19fw8O91Uv1YcIIduekl8i6NfoKvyRH+mAVaRKDfcQePj6b6BMLAda1apcqgnXoiYqbV7G99GfHO
njB9mShgx04UUurInnjQ+8vyLabKIdRflL+6THJlj6a9A6BEIpSJkggz+shNPwf6nCph1WY4xADn
M1SlqKGTLiiOLyDkVgcmtfYOY0hrtZ8PPzQrbw0WxTiG582LfLrasWyrgsJrSjy5GDIdfPFFH1za
ko3Pi4w3eCWIaX2/T4Qcu8TheMVkQKkD6I9+doO+sBQkqL4GzgS4u5cV2WT6bjeANy6FRTSMPCQ0
b2Ndr4KX6Cm063Y4VS5378oviaohypXwL7w80NxPgkprCqqyxAjAZ15HRAzlPTz65Tz0u5F+ZJ33
vp/LJzputJlq2g8wB/WQi/5URsAI4qYC07r7fWjLT5PP7fMWNBIturnIW0730tJiyeOPEGi1BtRH
nIFD+MAqoAPjTM+xcR1o2G6xm6jiuu/rnpWdTondTaA3ht/QhLixPJ8JHJXL845oUCerceR4kE+V
a4hGZ0auWQC+1nFeUid74kjMPTAz46WjDRpv5gxBFT8y/9b4jqTjlGFSzSvAeCgfUvpn0XuaTa8h
DyBQ2c/rcZi5ZdB3npuL+CKBn9sRTlSC9hioMZFrI0gcPtUIigWAPeqkoC20jCIgmKXjBoo/ypyC
sVmj4MoaUTwyxEUm6E6o4bJACVduGJu6ZRofYPPs2oU8IxriNVHsmZldjyTLO8hmtnlLHj7EF2xw
PfB4SnGK8HXEusH1WGwZxOU26oNbottgnhiFJVm0FY4bGmVO48veOcvifPDvc9CCpjMoHCDyUIEa
3hLZGU7thQIOMdXJS4hFNwq5Wh4bt6SXAKB+NFDkxOtjQcJ8DX83dYT/Mk1+V79/UeGLO9QccDt1
WM1pAwU2HwHu1gDmkCo5l0HzECvh5aBlYNTf90GFJCjT1Ymmlj1UwWDmnphTWq8JkORgoddqcrlV
PJjVsCMqUSAoa6atjr8L25+UQZMi7r8GsAzkEnWkWE61mM6/amwAWu8j3Q6fXrM4UhEgH80vXlsF
KwyHM9Af2TIKhvB5VAxMfnbaHU8AgDudsKx0Vk7AM6ltYIM5/dGgI1EwmBTLm3amjIl+vAXakG0V
Vw+yQKqGOz5jTc94TQmbNLVPjs7HGuGrQ9kGQpIg3OYH+3R1lPcYLTGn2wzl4l/b7IJib41BPWcF
ySwsX9vH452AEvOr5z9t1w6WQgXF0gdjgV6E6QVIrSecnaVxeqzw7T9FAy+bVfffvBOwc1bs4NZ+
J4F71EdJ0YIgCHcfQlTKfjWsfgUhv+EUFFTCGaPiDcUQZuZ3LJOz2BdSW4mTfNQKisjoE6a5nfHN
l6iReDkkcDruT5Bv/JfnyTsQlo+P4lAgaKOK887x39oojAsLQHTKnCgY/40a/kJA3Me6uE8bvorn
krr70gDeSyzd2SlXPv++HdonACFQCgc3+tmSAu8Y+MJnojkkTnHuwUEnwWbydEOeg7F5Fr60yS6t
7V9mnRFXKu8rF6XtgyXKGw+Ofy643fNsuwNUuhDir8hCGp4EV6wTlSzOhfTY6HVOy5MF1B6gpJHo
FobWoJEQF/C57azlcJW/xKEWSupDYY0vyfr/cnfV+rVC+FV+mXhrG0+nRpcewSe1lRDuICBQxdFM
6cxRF++jeDTIVluYZniVeKn9XOMDh7G6CkCYNp/GQksMpHAxq0lJRc7YHkUQb+4G4jJWlMTOUeC2
uQGnO/9QqMOqzUeMNL8RxasQU5NR0YsIEKw/R2ALjbyUVD3B7kl6EBC33Uez2OXNtWH6PSdpZ76X
eAwaH+B/g5LrOliwE5NrszeAMcpRLoDM5xHtUWEaK1/bCuSVgVNxmzjq+tGCOWeD449DLmlU9dRr
BnCO8ElyKD+3h06xbm0jxS56A485xNAuLaEE6sApHkhvpkEt5DicwBSkW3vEZRAkLHzU0WeTH//i
v9Gh1VGl3SAQOHbuU6ddie3sZU0lBg+NAQoAlTy2PTbGPdg0e4Q+WthbwBggqlv76WhCxb0Qv8HH
TR8skUfa/TB7vpkWgP/jqKtQIWXct5HbtHL9Xiuk0vokGXN2xuQTxRKmduzq5zzXSOzKS31DV9Pd
8ZSCGEM5Zr2zCHsywfNM+xj1G4GhfGQ1MYZRNmVed/yXxpw0Iho5LXvcOM+QHikU2VV9szjoeOEz
lQhVDLSh3kSDfqWinmAPEHK3FOWqfLmr64JXYSRdcjlakrQmzVROoadnfzmuwkTKlvBvnPlJ3Ni7
/RFclJo1nT7+8+eAkIk6F3FFTdthLhQv4jyvhQDzNaGNVDlWlVCdspiU+WNo66JgbinsJ/nItu0o
jDypZKkKhsPKdl/by4QmQehx8hQUDiLv8mRcKUfMg9Ah72kkTLfcVFYL50vhlwMpw5w4COugxPLP
BdvPciPVCBBYYE9s53dXzZT0iXfYTnkt1ipmKd6fy0ICXbIUJoFZeFwTYJTXtb7PkT+7+wjj/F4I
P+6mAYucssuxNHR4eP93LxlipUtdTh/Jt5a1N1XqOBHD38W9G3dcPQJUwB0Ualni9IWs0v3WpcTj
8c/kOl7ZfQVfgSG+JKyApn5sIaVz0fzLLG/EP4XjHxJPWH36BLKx4gf8YH63bkuL3pPzd5PqbFBV
ebUf4nalRqA8C7pgz18kLNh/8RHna7idxkuT6f3i98zXH2CCLxAMYS59aCBDWwbMaWFl/tQQsKYC
uRlIcslcdRmi9nOChk8XpdHdViPBEri0FlWmxpCtkzuv0zW8ZH17ATN6hjLLGU1apVrVi7JH+3N9
4+KCPBVNXLdE8uufNGiAGeSC72IijvHTeVRn9HLqWSlLptaTiJnv00yffx23eywTXzKVLiJEUzdJ
qLtBdcFN3/5R0dCNBWTkF/H5uCcYQMXC4s0Z7HnzW5J3TWJIkAiEH0nBvB61QcT7LNBJzoTZ43kI
O9gIjZUBFm1X4fk407RBLNbM95PZTNMLVBSGuM7Xit4ypVhrUf09CHrWVIr9SxhSPTxpdAQKjUpw
IpxAEHcTNl1GHsSdroB84Sp6OvTB3vW9ta3NYs340qH1rM5PIUsCOgdN6lSVndX88SsOpEl9XxMi
rtAF6nMvr2CCWRgcx5iab+G+uf2FAUTY6sfHNUQ2nTqf1PnlxNMDtEQQF/ecC/Ll7XE04BfNfMDp
XEijzpff9MxPaNyyj3mVD80DCbiCPzvmG8/eBRQ/oB54pXanziOPNTWjlbIl7kQ2X9GXrNh/lqtp
U4x7LkqRitM/bOiW7Cb4oplBUSz5kgnXYeLntth+2X/AQDAHY3DtTSs6qI7rFcWtD3sfAD0DxUWz
7kbG91JjKMPtlfJhGK2iTklwhom2UR21tN0LOqRppvMgjlIzsGBTXtXzoYH6bgEttHFChNVtXJ0y
7CXf0cJXV6ViAzZaNc/GusDYKlbV/dEncFupj5mnrheL3mWMsiW2ylNUuOA5+jheSYtWWIk5+MMg
VzgtPp47evBCK+ZZ2TOFjzkjTwbWmd5tqCapoBnEUjEdx6eiN+uyvK3kSiqsD4YYCjtbGFHD2UWc
XzG3Z4gGrYQoF2R6wwqvfE0litrMC8veIQdAQ0B/hyKW42Inrf7oL+1uhn8/PGgJQ5eNQ+jWbYQ8
IAKeMwd3T1eNrkldODfgfqgzWRmjpnMhAbleuA00gbWmnJTJgnzaGF3zw/iBJqqzhFqvfuSziKo2
jjQERYFSyicJumOXh5OEOSCNEij055JrvlbLPFZTtz35eFio+DC132fNQ8m7JQ5ABqa6og0Tz5mf
ACtXNCHVtqm00vBWHRm25Mun78JPgYtf1mw+IaUmQ509WI8dYhmP8puhpmPTMmIlKXlUfdtDyLV3
iUxiwgrksyivIcjB4b0ZbhXvLFPAsbx4iAaSOjW4AQ5BUKnExYjV+zuBDd/45dLWAbjaagqaTmUF
/OAigTcNT1E+cOmPFrp/K5IW7zJ5v5ztAsi/GB9mwGLc4yOWD7gs/8QHUlUD3vuMKbOFF69IPAxn
LnUnp+pG9PuKhvAPq0oEQHwedz/oEvq7rk5doyfXjBqWJfrNjICiy7QrBDJD0dZGeK7hidWtuGxS
J654SGcvwuVHrnCquace1ayheHuT8/oQk32lkLjyDbdJEkjaIQs5xwk9vGaSbnOgcLrO2+HCIivL
KG/PVhf/C/08p/QsaPkUd8TZQHDPHtiwX3Ba4lDvhTMQmKtWlmY6/vHAyU1O5yu0Zwz+ijiQ3ZwK
6vlk3W/3l1Ko891r3IyDBiAqSZxxX5sKF0Q7o6RcJrrD6JLjQtioOwnskoXb3HksYTr3NbpmQhro
2A6BG3TFLxm4u2UojFdAHpy2upZXDiBekYHmbgFLSd/46hrDt0ixhjvEFOHZ1Zsxs4/ybZ6p91ye
DQPI5EB+A6KSZ6AbU9YzrShbrFCPot/7BftrxMXZtTSt5cKdu5YyTJW1ulH9RTK1X07/ZR76WzzX
Kueyw4Z0JZJaXVH8qikomq0Pq/xhkqcPwd/go0XNyZNNo5u/VZuNYmYYnp4JTGfk+nl+KTpwAQ3R
kWEnU623LROYfSLGtWKlmTYOADN4zDKa9Bbc6APMgpXVt2Cvm8lgOIpjjjo9FugJz9ASzRsLxC0x
yDsSt+umKeR0PJVMP2K8hpwGGnd4eyBjy7svi9l3C78DgVMxKNnoqxtyQ+UpUcOAiUNQzmpaeKaC
pxmkgE/K8rJc1bI3M6+Ssqm3b/B900Fn2J9vuGuoK/85VVECIqZMWsfCRxc/xQFjXeC6TFx4qUJS
3hsdgukNskfDiC5bMcXU05+NsFShPh3v9IC7T3MDkascbJr2ZH8lutG7QYAlhOu12XlyO+JKlhSz
h3ktSA6d6cFMBGAUJ0Gko/vzY8AgpWJx/1EV3vD9l+crf2S3AGdkvJx6IPvtFMA4sp7rz2pO1lxF
E1eePD1+GcxXiYHRubQm0SL0pl+HuAVUcTN2+c60Ng8hP/+UV5fx2sKmVLdvX4fiInNXF+kNrIDL
5RiG/VDffwAcEFC9RfnNSPAwFIESGEoc6X87A0b3alz8C5UDLFFypSCymxiTbpfmtJFxq1f61q9g
zS6QuUOQdLVPduR4hn78wznDFrwVhIvWLalnxWCorf1sxuF+GLy8JlV1T6MgF8k4mF57oV9twwsA
XDcLRAnaC1jQKZQwgmE1AB61JpuQOJmMucROLWC7fuaH3zHF05P2Mo+tzqGJEWt2h9cXiZkOxFYS
we1Fe4QLSD0n/iku5A7sr/SA3bxDHb2Z6TdEncD2U0QtDMOxafeFh4MNsqG3Zomn0DTN7kledhas
9IfJRA3ubGZFtxm9uwGPEeXiMrhlih55j/ie73H2GSWzndOUN66bNda93Am0VzkxlwWlxEKwPVwh
7g1LmIcvCJrPpYXeS7OvvtvzlK43APd+UYEiDFa5Epng3DQWI4wVeyr/BlmfYBxv3qgyx9UCz2VY
9s9D0U6bn7SrnEGgl6PKiIXHKC/NmsSQouhXFcO8TA+yjLMv0idtDbVvkPVZn0qdAGeL+rnxthZj
nKowZ6Elsx85Naqx3+BZkdb6ADZf3GjybIJXF2XiSZF+cxJ+A6n0GqtU62KNC0LN2raYfdDrsQqJ
fgJ1YqMv9rBxNyYEJ6Q8DAEOlrIkLbaWxsu0D2FCkNtETOvX63fAL46DLm0p1mCHUqxeSC2vZR3I
+Hu9hTXbjvbt9ov0VdmoOF41ZxSeeKrj8YA2o+lGL5VpmfHQGmOhWvkK11kLjZC3oub1qwJ7TdAW
wlMs2M4BywoCd5M41+5yaU401kcvEk8au35CTv0ZSd2ReFaFPNIdH3XMcwOLNGCBSxVZEgEQ2XW5
irH4xkbpaUzbxLhXQmiRd3xEiNTLm5Z1qaHV20Nl75t8MlpBSMjp9GQV3IPoryEnYIhdFHBTwyc5
EaCRKpA08Vh8vauGXvUS5ghXQQW3zS+82ldfHP2xPjzSZEP01jHpvZiqmoD6VlfbBDT+Fr4dzDPI
2LccwBz62kqQegk0Vk3IG9UlXieZKvOLFeA+rmfsv96mgMLNgPc4phXUgoxEPrBbilMnBEElKWrx
x0c7qgolveoBEgV6f9lLrbvD20hPcyWGoyfzzPTRZhvpO2ovZAIeN8ENL2Rs1Lit+JsJjVl2Xg3w
fzn02kc1yFp2qRTNRQ78mUC0nyX6GsWVcDz6QCrD2Fa4hlPHa2aY4B/AZQ7cZzIh9LG+6Rpsfltz
imkV4e7ZXI9MZaxUXoDk+U9ipT3Z8N9NSmuKudD2irX5QPscVrSTQGNcYgnvCLfG4ZsRDHGQXvdQ
AjsTsxcAhsQiv9YIg5a7ODhrstmkguUA9c0GU1tZTQNqXhDIsjz8mrp8bwFE8mYFwpWQ7USNrUkx
u3OLpOHQi64dN++LWDr+2v+3phCz+FqfMUvuU7ZvOcAuX38FTEW9gDF3ioXhjruMEXEemRUtXP95
j4zC+S/Yak0SAmoIkmwfY+rWFmAMJZRLIhYo5nShaqA96GR6SjUujm2wYGzOWNJzqX0aPhr9ss0y
zGFM6LMdl4RGHrgUrUqAgptCKvrBBzqE3Xye3dmyVHa1X3EMNoO4U/8bHkWbpAnhH7tOzBU92nD9
R4eMqGENhXZGcWzVYpRhF34vjfpqEuleu1MLwEsWE2rAqYvXYUXBNcTwVjbolnElL5TMVDNvEU0Q
UfmXWMdtPC/KUx0YHehSie2BKnSGro/UN0FQIpuEyLlXoH5psOE2Vh35ct3f7RFjd7czNoBYj5Ai
F+TxdA9eEqLQ0oMGvsh1gjdlGZZORsxfvGb6caEieQ0th0MtZ0esFb6rrHaUG+GKxO1x4O8Yp6BZ
SA3YqdFnGmhW9iqIZq8aEa439Andr60sTGnlmsGbqL5tjRKkml1d8fPH6PD6YFUtmt4Qwn4jKJZ9
/VENtPVe8s1RpkrahFInCK2kUd2yfY84ayIUTBot8uYZcKN83QVjHgV3sYYn4T4qmgAsLVhPYiC0
Ervbpz7zn8qS4UY0njKu0wzrsH9SGc5zJjxwx1Za9C+Do0bhGgMTPwqpZVB7R1Fn2DZ3YfiJiOHK
IH4IH81L8p4qPIMTS6NbEky9V0ZIOutwzRGCE21zWHSAmtl90g4nb+/W+tMzaA5Y9YgLUdKKnRXk
Jr0ThDY63bF9+Wbt+ffg6Hox270k/dr6Tk/hhUFZLTEt+uI8kUpb/3EDx+76OStG7GQh+bssMlBl
d3y1t5twYJMbcFMJcyOoCMBiyAxNmaayttXq/pwN+m5DXwucyoI5birqBuRtLpsajfpfxRWCYEQ1
tZUZ3hTtSzRPaMUY1/xYQl7k5q03Q+ellpxz54VjK0B0Apy33BvUA0OIloKYOOn/4Gm3Bt/ktprb
QL/GL7MEoLFJUOYnGCRu1fzWHUNPaiXCqwslCedcdI8x97YZkmmIAfPob8Mm/rbTQ5T+tyE9KzaK
gBk378bQmqZuRhId0C9eKtb3wXDs6EH3I8MBF7NRAlPq6AO4oxo1webwkd1F4kPVMHU1bXI3AsuF
UPBd6TJv/I/D7WbvQ6ZntF0JQj1s/oeDD+UWBRmJXqPfrIFCOsIhlVmN/dAwsjnr5JvdP9/HgcBL
BmxFHREol7DVj3Zr7unUjsdJflbqF7Yew+ekSC8TPfQNOYnq+6T7r8C0IRETtrLRd2iMK54kiId7
Aorcj6XdqUNezM42NZvQ9T+cJwabHuHWuR8pqcQgUU3kk2Ta7ireCG7e9CpaRtv766uyAVyf2Pdg
EeMCMmpzqNGHgVaV/RNetUr2DyXr82KEo6NZf8MlaTJU9FxaiZPeDpT+vNs7IpVUJTPGlFX2DUJX
JZzZmkQWWckJq+ivaSVFIYTMDCikGswGH9uVklNeDYe0nDB13HnTS5ryQvMBbdDvPwqNn+eLytwO
hBr3MUQI65hyZz/bpg0zwWOV0CAPQ1ihwJEMb79EPaZVn7byTT8g96Xbgvva85F+Ig/B7Ab+qzcl
wA5bGUK3znKENx3bghbzrHudUS25gxXgCJdLkFVi3Hu32fgfaWNEkj8ByFov9+R8+9+59o/biTBd
xVYwSEt/fkrqthplSsZq8/pZ7On+NgHglMp7c3sS/B3ge4WHRRi5yhd+jR2vWrJl/LxcffMc6sXP
Q4qMgurc6l4vD1G40lRqloruPiLXt1W3EcB7G7Uhw5U9umZmPCqgP22bds392eQJAIe2N/fEuy/6
3BLK6rnzb6FEiVAXmZmCCppomtVgcbG3USIv5bbLLJ55bqmRBBhKTNaSbx/31aT3TT+WSZnq4Nz6
eIO5wl0G8GliGX0hjlBb12VDR3/SH5fNyHSwCJlZe5M1ySpKKmorhaZ+ZQhXDBm+sDbKP5xZtsaD
8Z9jM3oDStHPhrscKn6Rvfe51xUlbjMb+07iex+vc3AqSiNYpsnHbZ7mPprVgJ3JG9DOEeWPrUvC
Mo7mAjejhFBFDKG2BOfJaRxjpH0+aEj6d3AZ07ZWCRdf7dy0eYQDgtcMKIufZLDGa/TZQpMxJ94N
W5rCJrjENrmzVMYwFsInHNPCSV/RBqjPXwtFE++tRJFyE8IcCXoXlwE2ldCnjNx7ElUIojaHVq+V
UOtr3My7ACdqlxYDPC5FW2mLzyCVa/uVxBFxki2IDMp8jep/7jXsNdYM5ZWUp5mQumtaPQYgrepi
u9PbQQlKUUB6uvYlLoE8aM+Yn/mcEVBRDDnEJFItUMBi5LGHvGLhEBqnsGWP84vR7rGJnsurE3ie
PqvFYkc0/8uNPLgd4nO/RvmOs8ERDSOcXawLOE4kfwV3wmFcHDhFFLIf87suT8S/FPpawKhcT9jM
uBVbZMANeB5WlB2KLOPfHuLRu3c9KS78xfHsb6ARpBfgtv+N7GUAEHoYjRfiP5D/DDzOeFB2VYGD
BPd+BLSJGza30KMCHcAVzDenKWs9tFeWjyquGuuwIOOEpHMccpFmdUIm5oXt/0pkBnYCl5dtNKFN
hCOmsgK30l9u/yop1Id7yjZqADsPmrNlToyKE2eu3xpkm7Z04BfxHp4aYhVpkrj/Gtw4xJuqSqpA
lVioqLs7eRiwwCuG7+hcpGaUVNX9Q5lh2BMj3XlHWgXFM0nYVJjXrkOa6YDsQuNiRwo7YoGjsMPX
4g45LPMXc5V3O5ZvCyAbho26yAcK2wR62wQlkuMWsBqFUxptrsocBPoTuD865tmzfqXjhDxQ0Lig
AcnKmWXkZvZwNmR6VkVlPnFngALzhPL41BJuWg2ijNgjnC+sU376tBFDiD1e1kd+usXXeJYp6PzQ
gCVFomEAGzaVBPbHILhm6clAuGYk7clS150tTGSM9axfts4szt3QE2ZMImnGWNddyMdvP8/RVgy5
UWOc9Eb6x0uQJSfTfNomJnKjIVHuSDV1Y493fEmVl9BHhwJm8rr8/THL80eUVKHKOoZgDp5iUPXw
RzTKvOzpq30+WR7eZXHAjMsJgh0WYiSWRgnJVnrwTQO4RWLcNlulLLZVv1dmUioR19qZc2vmnn4f
yFN2HGcLNCBGLuqo+M8YtyB87hrHHE3IruQcNgsvMMsUU6A/j7b/TnyNrI2iwLr4NvfVnSitDHl4
VtNp63Kb6npKIpN8g9TojU0I9Q7KT1kPA6iEvcTGzxUAFteljA4KTNM3Htis3Xz43DkGLxp/vGIq
Eb1Y7FMX1Ireyb0dEBGl4AhXAt//1m7WLuvjeNcmapbgql+GAE41AkuW0T5haSM1CMHAER9OqBVL
WauTeDDfKs1fsO2VVfPl+68GKPo0bUQelsfhf6pZwW50mp3bt6elIWOcVBMe7xLNEM/gYjqy+CX6
xTMdYmq4iKBOGB1187+dBqQ6euKZrtiDM3KBybDMV84eKauBddpNf981056X6onA7VKzZ7cbtCsR
dit4GLbL9jftBf3+XvohI8OqhjIa9HgtftvH25JSw/FVev24BarpKk6FSq+roPKAvC9eyJGaF0C1
v8wApZYtCy+G1RJzEjso5EKj16BszrXz4QSbirlLC41NVSvlYRNn0UGz3zzgczwSTqrbIB1mOHKD
c/ngVNSBTMN2t06Bveh8afv+L7eCr80J3xWOIGccf4CKvoiV3KF2UImUocHiV8qum4wo2URW00wp
l9DnQxZjeOykFLMQU+WriD2GLUuWYT2nf5UNC5cVl3Nj4SuNzeLBaTlDPDmU8NhwQWTPcxJ+yFa4
E3yE81GwhEZ10kmVqQVyE08qILFdDF1LZMrYGfds/xQ8En3ahojQ0Tv8Vic4mW8yLLCx4CDdHsjj
tx0QkETn217S1t3uSggYx/inyoucJhgbavmRyCbEeOpZi+WD65tJGJ+vyXzWZghHrwHWqMb2jv1Q
dGNYJLr/wRaGmjsWDdMa8xVViZQxBr3H8FDmgS7K+6NrO27iB5nplzrH/MPn8e25JTPqoPyXvNOc
YYgxefcv+I7JdEWrRK3eiylj9eA+V34OA0ik+S519WNqo2ii1rlEsuq9ST79efQOIKokb8N3XQUn
k27INARH6z96FwypsOpwsDy6Xj0bZ1PDxEFp42cYgDtoVmNn4DM9tI/fIayKLWD4kwC+qBNK3EUd
+ZZ2tjcMrSZoN3jVqlpSmnvOA0B+80swzq4ehzgvXhj45bHqEBGVYb/jTMufL0EGujOkEqmk5WZv
h+IuvCrXDJBEDxo4wzniCnUxVbq3XDhnvg/IKqMH7TERfvyLub0+pgtgl3xaZ0TxWZb7IGBygf9A
OovlTs/6fZAWXwQ25q0C+8lmv50zLzyJ4N1QNdRHo8fT6yUH9ms83pCc5tpT8D5Xz9lpsFFU2B4N
+gSel6Atq/esd+VkRSE82GHsRc6fv4zAv7v/8v+t0K3R7s3JLMt3GoHhMe4OSxAntGFE8kl1/dGJ
tHBX09VPWIZLekK3rtblDEGXCAKu40MHy4ToX6s3RfNjxLlabXAmzg+3/Yp7nqoIFncgNdP1+oEu
pFnbBMjiZMmQ0qhyxK/FDaM7A04W7E1f9Nyms+6OlPrayTFilVQmkH0mF7wUBsUSV2S5vooCAu2V
ymuv+a4jw4Kc6XBHVhXAkzf0G1vjUFbhPRzjrzZLJ9YVT8yaaHLx7ViyLZAgHSufY8I0JN5N6Bvi
fn1QmF41iAyVDNfCbjziaU9+5s5hSoOvk3h/TvLl/BUFhaqaUL1dLfMhDx1GXMI9ZpFlYjy/OgAp
FPLcbiPhopsJqkmt7yD9+3cOZsmOLSnTsUopQi/v7NVwoKhYMznDUSHJ1YWDP7O4BZLk4fxJNECU
XWBLXq5wzuPaq2PmP3eVxZGw2mmS8LXKO70erX8EJq/DTWTUCqj8Q7pIZh3vVOajxUBDoiQWLxz9
6cjt4n/VL6Rioi7lF5WSe4mFZ0Ck9WnquFkKCKsa4AfUovE7VT3Kuhw7BQo2mQt3X02LoRkwScf2
Wjeu7cHkFtovEJCHfGXkVR3nkWgT5KRYVMwuGS3Kh+g3ZCrR5aQH7czQ1+SME9nOya/1IFtheznm
dydOn59vYgBxdJEY0Gd9B4OBJ19FxR6i+7/+tL/3aMb4Y2YZr3DMR9VowerjMM6LtAi13wDL+ose
0m5zFSFkM1hKYXp0IR6cTngiKpICW1EsZ8StiTtDIuJb32k27CQXqb7S4UH03rPrW00htkuuq8G+
PgbXJ8GACjIuH8wnXt63h5UXu4uMij2/3dh1CL75pCWmVoGWu/Di+PMrwJfbxrStyz+FWYfmaXZI
JSHQ4dqW1Glq/84ab1JETXjGcBOa3ROL7OmLC6U2naeaQZjiwDWD+OYamGPoKq/LLRwGVYnXtv/j
gCaVbTA0LPLJ5xsKhtdlqn1L4yKk4UJzZpdshKw9NkeH471SQvexyhFkBzaml63Jyi3GhEdILVzM
UyOKGD6NbD76Qq8d/JXjgSizvCzoNQMEEY0CAxDmu7Ixu7EaVh5ZXbrk82OjTTOA8YrPgTPcEnH9
0/OaAsergj9cQ+GZkQ0KMINS0epzdD1DWWDBTTGFMIvW05SOTQs14IvLMbKsSMp/emjdzvz3UtSz
nDdCXbEIS8sF9ywmJlzFoGGyhB61gD4b/xz9dRIVzEudanaauxk5U+DkvO5V3zfYqA9mHpocQ9Ky
I5rUerOOx44Ous10EubLnYyZ0368eXIyufy6rvOO+O2ht6wnqp6tQwhA3Co3VHADRBhQvZCyEEPN
W5OjXJYh1RYuT940qnE4ZbJ3ln9QycRGOV7GmrTw0luTFcAx1ZHL8grlwg+5ekTC8K/meyeQ0mo2
8e18LHvyEeggRROzIzK96xp3uxE1ioOpq6K9xxDxPhuVsAwCHwFqc8EwX4q8ERraLVKZxTzHjoh2
rB6Soex06GMcjY6dXK+oxypA3bBLbAKcr+Wcsh9YXcVoeg6cyz5apU2SCgEP3gc+EBQ2WzmLWGZQ
0KnvBVG4cAjpoCZxQVyAoYSicMLh6e1JV2D7jGgSncdDubBUDXU1PRX8f8nqmpU+ExDt/JmtpN5Z
sDpnVL9xCDCLnzFaKu6oOFxCqkRflRp0Ujutu6AsqyYePPNnARKlmQlmOR3mHdpzkt/r5OTwzOxF
zpygWlp26x9azAnE07VF0WNUnePdg9l9yVOiScdWCMSPdtEcH8entaHXMuwX2e2Y/JwRt6s4dicm
Yd81AVhttxtS12QtHiMUu9+hwEfTlRcx0bA9HgGhyMAcX40xRmPIZCrCxLXRhQzi91BwHAZAMjkr
PiIYpC6hSxVKI0w0RodLUFPGnutRlPJFWW8wRCF8bvyJGkp4xPHADC5YqcYG0BDpn+je8C7J90XJ
5bYiuHolhYiv59+1Zqe6k8sLFu3oOwTT1XG9t3Eg/dzzKZwu1n0GYmqwhc20lXgGEfmaC/ElyV7F
tfYLkrDT4v6xfwg2pK2p7JjGAotSkzI3KJhOesEZvJZgCR7d6CPDBVD5TQlze6iFTP4yo7YEwnZn
joCtnvh2YcY8kz/kMs6XNcIU72iThRSHd7JUsTtEVySWOQBsqWtEX7D8kCEFHcHevdPm7cpm6Eco
hIk+Uvs+CKCg6WGo3alp1JggjYkosvPA05bitDjqNNuSecr562p8vicTjqDjvZCVvsDhE7ujxJv+
qJcxMQzifjfHgq7ib4jIYqeluzX9bmfYBuK3EuXYfiVZspNvPfPUxu9bDKnEgFTlfervjm7DkLxu
hCcWDxViHGRol77279uPieyX3UFsbiH3zxoeVi4t3K2KQLUrxQ1Q4tZ/LrUoSaHiGH3IArnfa1Rs
9vZiyv+N4O2dXQ3w1z56X74cSrZSjwYq63Ee8ayOKuJtNHMKF+iJc4Z+iOmLet//d6HjP4Acgk6D
mMQO9OmTpgj+QXGwx44wiMQeV2z7caoKBGKucJnKyTZyuMXdr9iPeP5Z9xMetJP/AE/TqF5SYAsQ
GHOGLClWRstXYZRETxql6F3JO6qX1WDIR63OEOR/8sGs1ZXGLIdIq7KBNN7H2M1pHbjoMQZxK/qs
AKLINQ7bqMnLi5naAz5kq63ZK+m0BIgaRsH7vkp7C//Tq2JhBMP05aZJ/251E5Lf1dqYXtdewKn5
J0PPQOY7FvEsxQDg3RP7ypzfCV/C1Mk3Mt5z73vdSRN0LYoiIDsXAjmiWSFuLNi2W4gowdwkfXR+
316qGbtOEKdJLDnum+KrVXzWjosZ9hs6fWq4/U/mOf0CWEfyrWmbKG0lDzJrYxH5DoaVGtVez+Pm
k5WkF2jnWornf2Q/PBwz7dI1d+xiWuncZO6hYNYLwyEDk12ShrrNTmvgsTDfGcY8JiuXDu7O4A93
IpZ1olr0IFr3jbK8nk3/ayoKAC+QDBpd4mb9yqtZWAThn8DFOsRjoHgoCAl0BcK14Scu3NhOb/Bv
tHBigrO9hh2IWNEr1ElPohVC2M0xUSVD7e4fdbe00JQuDSv0zW794wzM/daKG7RTLqk+Y6zqwUP3
VH/xbCiXLZUYX6lbNbz+vYUml9th1xV3twIP+a1G8RwSr/bfdbxOERdlZwxgzqstV69Wu2P2opJS
btK3M0qKf0XtlbN/WCYcDTEwimaI2XEkREnT70P5ZpA8BFENJbMYD8xPicjRgn2KexGXc3/LDCod
5ITLKzT8+IISoTIgSA28F6KEpmZdo6tAyhWoT2JAGYJr+vjd3FXAgW6mfQTMbC3fYAg80jdp3IGB
NQyr4aqDm64lXsGKrAK1vrP21PnZoJmVjLC9VCQRUBOT4IPPQ3kaSlJiMph/d0D8bVaBJojjuh9R
sxYRPPzXmWOX/TX/ImPszWPHWJ0xt+Vsi+MJysGSCbbKrjl7I5OKqWCD4psTVFwu8yphsf0tswNQ
+DcSQJmNz1J1l+6zazE6V64k67W6nXlvv06xKmW76XLYGyaSoIhizWQvhP53rnEcvojVzyrXKNNt
CCVGIyka+2UkLMSacsUpQT9xPqFtDrrM86V8W7EnuazrG63FhqZ+krwJ1mwrgY975hEtIF57mkGk
xUf4hYW6wK3wj+WSaEthUC3omE8vzCSe3ds7ksBtO0buGiBO3c/u4WwwchtkGAkD5OGTUUO0mVSi
oDOjdx+FHWuAnMUw3k+6ffoxL/w0+N7LCtLsaUuaw7wUIAgqqtMZChYnrQi3fHacujJicdRNFwpZ
EnFPZcmnYJ0MSRJDth5JyKS9nahzWO8aP3/Uj8d4Ehzo9vWr9ImLYCJSPgDeivJMQMAJigynfc7b
lBs9e9Wh5P5QIyxdYA6031Sn/5NPk98IjJEEcCIVERposXSdo1GzFDCZrB+8eD1/raUIp/uaUAr4
OJ0BGG53Znpo2yfbQCJ+b4d8m9hN1Dn3mUmvIhM5bixtX1ovZ5R0fHhTqQsiKlb/yQKbvL89GeG5
mF4Fot3Nrqax8I+MBmrP1xckg9PuOyUND2BHzKATjdppi0XtuYxoSi38chRLGOqUIhuj3TO/ZGfm
oazdpQR8r6VzjmDR7wlRBiqp3yMMOr9X+c5DA6Lo/JtVybG+jPW3WsO8c7n+eophGKQBjNO0nt6z
D3NSIPzKyQMKc2xupOz6IpY+bwJyllqDUW7XpW0W/WwHq9soUiwz/bgt/GFtomN+H+KunIjl702o
ZGjAWejL/I+UM9iUvLUZH4tNIcCxGEHmLFgZk888o8DgF1oCiaS7LNcYeFPOORWSY6EvmONwdSKe
0wWeOhJ2T9Fe5exckNvrAweRArJvJ+AEVgBeR2jLsXcXMxEUb4gmNsBHtPSXIe1NAVOsgUvd2885
+CB7rkE9R16z/AsyrTJDuP0oUt++xo8bwLjtw5xtX2YOhRkG5PEjRFowlQvGUbdwa1yjB40HPc16
V6E4oAskg9i0FU/0tkLyix4i/RY4zPQLZWtZ18ax8VZ1cduZUT9w0BUJakgKgZpx9w9xtOnOJxb+
Ib4vcaMkcses6Qz8sJ0GxylXMcB/VlsvJJy9uC5+UZeViYINJXpLot5vy+MsraSkCjIU0kIT0LJZ
ouxp0Z9+bwGQWbo0uNdJhG9GUe9WWfhK/kq/FNTLqhdYij+9ZwxK2qOhkOzpz0g+vy3su7u+JR7O
PTyp+CBS1ZARkLUg+HFl+xr/szcfxiX9HDdh6EayXAIY4Y9aTHB3fVC9lWmg8HPJU3jHZv+mytk0
Z/4KIfNw7mJdMuJq1T09rZ+6Fq53DGibEepLwhdyameHhWxf+6VvcyFfvV8eV4Dv9porvyg/b63E
e0jAR/LTaQun0sD4s8fhUd9OO8KvDtFRfD+MePL8dd0+WoZRNbAWGDsihPLrRrRSev+4eQx6411J
XE8DgKMeSzUBZ8IMqGfdSgACxjOKHaO3W0ZVW1dqBEC/pgvyGenvzngYQeLie/JXFij85JWnxAhE
7iS+qEI5vi6y5XYlqXWekgnaf6WoDNduiyNgQtWtdavjsh72a5FT1FrLIwUv6b+SwWKa363Vn+/a
GojT0DM/Dx2RM6lVCQSGN4TUkKHav9/zhtEj0HgAgiBXj71gbeY3GpEWzZn7p+j6CY6oTPIcNH92
gAjH/9w1LQQFoMDt4K+LEITU46v2llLVzOj9nUgEXQD8XWJMKwnVOPGgeOpQXQSC54xyXOcrg/0U
IYK2OxvA0FSkvdEQtpGSZNvKhDLoB0HtvSVJ2pfjtlObzIgYfzVz72dRU79yA08WNVtofIVK3foR
iIb664bHvbr9M70lQEDp2+BmQs/VIdbTWyalPNlzvv7ssRYQQ4lmHJe8Lg/jLUpRtvEVn11VY4jO
KW46N127aYh+yqetXYfhZghD9ddnVnhE1lwVZCw+lN/zGIlF2g1G1lx86SJDFaGnRgH0WVhNrsTW
Yr6CsQlbWj9gDXrFj/ljnikJ1XniZCESb7y1Oe5sD6auxyBybonuFqU0cH4g4raFk1+15mye477W
Ks3+f3v0KQMaX2UQxixRj5ClbCk+SfeKQR2afXXKNRGKWR5kykOkyOYVJPXmWyrZm7//qKxxqoMP
VKyF/OvzE+05yI7w9du3Vo84hHd3Yagy3K0bcIjIuv8QTdxoZn5DgfitzWr2RQXqYBmgwlRjZany
jD48WhfVyMefvM1C6+wVAijmb5QeQjzVAtAAHxSTZD3KBbZROq6InQOeggHoUcSfx2kGDdpndtpj
GSaVCPvJuQUderFb7/1MzXx73c2pUhO72KZdg2/EZpdYYEUqArkYzmf8OFP8nXrOkOhr11ONnSJ9
m5zdjhKY7khiHe3C/KZmbDsqJqP/lQk3aqheV1N3VadeYQjgmYzbjiUD00tvruNHAB2+/Bv8ysUJ
aiBo8lDdlhdpwWD0GisYrToeYP0fiyM7dtwraGsoVh3WXwxjEDsVRbrJAuMUzAaLJ97vl5w+Ui61
eN3+Whgj9bltScoxjqiuDUR1oKHXG+IM7nz+xEqAU72uSZ+8jwEbdXDRyMZvOoMj+Q6hGCdz3YT8
uBm7Vvpih5yY3WsD3Fh/Uder+73gugzWdQEJ3cxJyqrTwL5Ubr0ywi4mAV5ck/3W2X5Z3nEGT2i2
w1T3kZea56LK2YjHCHLuTJOjNX6QuqJ0mVN14WGORLFfeZzaeSpdHMXka6APcR6t5Ff3dtfH7OhG
FCpA4cHzQA5uy5EfX4rwQcPWiEdjS8ZEY4llS72arOfhKdzHnfzOAkxBYUetIRg12m5k8p962rlp
DaUU5AZ/pc72ALlFFWtgpviJUO6CZHjIWVE6wfbZk2TiFr6gxfk4jHZuz6atWmRSxpaJsADORu+e
1LViqi/czyUY5Tun9cqWhjqdYPRtNQSup5qXEnkaeYF2FF6/nm09w5+Y1aCGyWrguNMdC70YI/v1
VjYchN2g4QOj65TH05D2llbjakfkGYIn4GniAxKkls1gzDPivQRF4o6Uk4RI7Rzy2Fd0Ti1eP20O
zx3V19qFzMrBUqTyEwovU4kcXpneRPcENb1Afoh3gch0lVdX2WCAUnRyuZsfRPRanYYi2cbJFmKg
iYtLVxI+Kqj6e9BJwHI3kWHkcbC9AMZPznyVdqwD58pOfT+bwizFq4yG7nmP71Z/NYQ5Y6H9pZW0
RUAXdwh5cfj/nH4+nD2XJxvGd8KjNKuYg4tg6Y0nk3hqs9Ku2vUG7LsWdF1jP0Sgn8G1RmJNVkUF
8M+emW+hTY5HcnoFAl16vu1HWSUAdEjbbYemuGOIxxHtdSURwJ2r2bRqhuvbCe+8K0eWoJ5OlOaV
kHk/F4V5dris7p97LOXNfHOoHEVtaLJTzMgh9HB8CRAoZa0NAPDMOMAxqe8CTPSkIxYE25JX4AA0
S/NFgaWhXq3nA5NyIATYC+h49lt12CUX6Luii6355XaLpw2R5H49WW1kkeBoAXw6iOuRyd7jkE3h
8S3ylnyImDukhCVXmiQSRfazcEQHYUzysfcvrE5hr9t5Woo73tNpENSF5oGZJnmO7MiPf0rBNAac
2OX0XHpLQge5821Hz4ZXGuhB9xPu3TWcWL/+2Cv87HiR+CSFCbkFMs+XHtjZaWqL5aO3B8aNuWJQ
5P3giWC9wb/Y334NNuIxMlGcrRBn5iqUT5txwXF9mWG5pkfkxH5114khfeQOkO8GSrZChC3WB3Qz
3B2b1JCtSUUgGd3/kUO8swgmgJTD8n+Lw0NT8gCeC3GZt0nN7K/838GH47Hgoge68d+jTYv6g+mv
HqbadvLBXXyokqwIDaoeFLAp5CuCfbDVPN1GnnnmtnowZYdDJoSqXPorDTFQajaPqaaD2oNIktJv
1Z8uxuR/m6g8GMbRPnsJ7t1m3p/7lrX8WGsLU27KePxqtf54FNrebdwypP/fSmTvIE5E4Kc1XKDo
CtVA5SeFTR2d5ezK6H4lIC81xeIbV2QC4GKg82tRMynDVCzUyETZQsnvNZRyRC4cdJHkW+JGA9fn
PW0krCmnChxuN2TSOIP7DUIdlfdALhz3QvI/1H4eUHVN0ILE+y7iQZ6HW5+Wc61wFcsRVDrzd2cx
CGo/xxAJr/9I+vTPPFvPe61mEmGQ/UTv/Pi51xRcuGR3G007ZolROLOBxaH6MSq3WP/cJwG+nqr1
LCa9WWqtUWiiMbGJYmhAA85mIlloA//iRY56o+y3me1aQRTqyPcMffUKnjV5d8U080A/MyLmpPwt
6hCCfaX8Zp5vcKGSZKbLlS+HayoJYZphisYNutmLTd9osw8B+Ev6Ql1VEj+UFzQWs+45hupSByr9
ow2V9GYRllTUIIq95+TSnraWrfwSga7QK4DOiCyqoMRs6mnY/6wAFJfHGjDghU8W+t/56G/owxhk
prqs+riZ9sLFEARpxk/vAihJKRCLb5a1NO9CTO1JZ58OrS/H5VknamyB1u5uJ7I2S7sHD7qiU3Ei
3ddcHVDdhs3BcPXT2CdsKLX0Ndet0nEwd6NTkj2m+G2VjaiHtya3Z5UDYVF2rxB85PjSnputsL81
i/HgB9ivsmVB9PRbA/ESzwNAP1L9jhOiRewM+VObRl2qE5FD88RNKDFbZUXL+8qQ9tkR+5B0MKx+
oXMNQoWwkveC4gWU/pmtGIDq2X4SKuDlfMvDyG3kcCzPfXV9uwUDEVMqQ7/tjqjUsOra5BrsWVHy
mraERB93mC8uH6zO2tgdPVb+05u9LL52LOz3qvVe2nmK2APvNz+V8aOJvIhd0tDuj8cX7+SFgwc8
VuK47pDCqO3pUwYd5UODb4o8c88QRvqnZPm/fdFaa7copbEfCO7/sboEycElZcdEbDg0gslSYD4N
563mJ0Jq5a7CuTrJZRbYXPYBUuPUzK6gj4/EMG6fMS7ITXgIwvhcyB8TT6vEVllAYt7ylXLAv+8i
k7qBFwu+uhgjKH15NYe7YvdEeIzMiPexwiSEoFaO2hfBoEqdb4vvI24fCjvNY43pQwjQuIvGp/xj
l89qMKfXOlioivmPYXrdclvjBi6zAuQmySXvt2VIRKmoTguXc8qqvxZF3/g2azYep9DpzMwrglOE
m+bUT/pc6eunjTh+ykedKj5dhaR4cWoMQXmbz8/5BsTyCsMUW2A/5Jg7tk+/taUU7rQ2vGcn3QRA
jkO2rJ2G/CxzAP0UGr7jvo/nx1vKzF4RyAz1E42O04K2Uvw54FVApgQC+pLk1+GFObBsPEfEcLIw
Ktf9uvt7VfB7FASpQ7ArmfLST6godMrbX26UFQsQJeJYPIUcUvdTBk/0d9DGFPsK6rxtIz0dR6IZ
HL46yFl95MdZufIA51ZSQ2iw5NY4VqNZ/2fHx+sKPjOt/0Lst6gjB9ocWVsGa5V9neW84EO4jpLn
T1thYPo0WBC9qU0cKwLHtwIn0SiiIA1LQhg46pemaJesorav/il62Trt9gAHVvsqZPPqeSAo7C/6
yi5+3CVecZHwoUpHy/sdGe//lv2LFc3jETB33v21ZdsY7R+loOjL3V6ruVuRFJ1jbTQEzJVVUN33
DpNpPm2ugMCtDvYk834bWAmeyA5Uo+FLk/sYu53wKL2zFuNsSOiZvKs4MkHSl7jM3bsPLFL/XG3Y
41U90qAiU3WmY0Q+cyfcDGQ5obbXTqlD2tDfApEl+fWr9msKDmoy3P+67AmtIGoqegVGLycDlVBx
rsEjDWF8noEEHFUC3DB/2k7NsfYvps/33tKXDD/T2lIXEd3pLBMkV082LrMbwKalKcrEIH3UqtV2
21OVa6N70lNKLtpMF0zaWLst98HWNf9SVxh9hoLMSmCELJo8mmGU7o2EbK400MZQ3KMCEEZ1je6b
rDEd5jB9JDsv5hTlKS4gEHC0IOgPENYHsFcHkIGJePYDJu5DqjE5YFUNHDF29LyR9bOy9Jx6qdEi
UsRc2DxqvwqsiHmrjMh1av13YvB+5ZsNo7jhCvSoo6MU2x/Q+Ry/6OfRp301Vw+a9tGoh53INDSh
vFfVVMupwMIWf6Zl+oYqiVow0WouueG/oo83Q15FsKfg3WVGYdBvU8Z1hOkepYzjr4RqZqW++RXB
9rkKEkda5qFRVrKtLzy6OX0WORJOVI8A408KUkPXXhq+CDCNWHkfNbNZGKoTh+h5ZQG0seZwombe
APSmoJ7xml6Fzt1CdwE5ZzQJiivxYs441L5t5h6APYqcXy5jgjHb745cOVsRwOMvRHuIyNrJBQWq
7kVtTrqrMBUF91bckUuk1bEdcULoYza3+tzFu2c6ElB689Krwcpmr5Bobhf50is7OFLgbPBu6Sni
h7dVgV9asBeCfa7EhcUxRbHRqh+jifyy0fqMn2vz8R9aJMEpKc6kU7Ks8AX1qBkR5bZWTkJyq+RC
cekBnxDC/e4K6+M6/CK841vtomX1NIsX3dQAt/VDV4KsidR3vDDPLZHXocOPDxPDFkdxuP0BrSTz
8HL9o0jqnDgn++DHwrdSp6DeFoFWiuEGzkjUZLHN8aPIJsF5wDWOzItRh6CEEy18mLHDLTBH8xS0
k/K8LNV8d7Rx4joD3HwqXDQiK1l7TIkqotF+rLAkh3FWJjvRNpUBMfbJvxKUimhAHmYu3r/1NO+X
+uYxPb1/DBWvzn6Iub5AuCKwOiycwqx7kF3cki/xP/Ub688E//BI8iZjdT9HlMJduVWknDDo5dP4
2szJZ1j9xIyQHthEuELOQ6pm2QwCLb0qZCx5SF3C37OabFf3ihoMaaGcVNUzB6Y7YZgF0albOEla
thq01S6PBwD7byg6tBlbTfhKAiPfkX/J9qwdx32eP6hkF5Ckab63sSXqHNuSiiZsy1m4qQaNNosb
TI7l6Cq5q12hlnSHVTx9yRfRKaF7clDlCHT3pCPF4cs19sRZd/nb/6lMKpgSgwA7emwneQE/HaNM
sEl1UrOuowDmRUR/FRUulrcwVfzJhw5ak+IZ6JoIUPI9qZ0LwCOEElZDIanQmMFr3oAWgybelUIL
5RkKE0E6syyMZGVP+ZJLkdk5FFmquNpPogjeps0QLQw5FJM6A2S9d9oDjX7C8FST2+EMPQ/GRdGO
labWxYPLxhtIDrmXT27mfiMozMw+mN+pMvPBDjaIDtsALhWKlxcVrWb7TYCPgMPGXCOGzhpAXl0b
w4kHRzeTpmU95aIpkFOuqGmCjGSRT8r+tTNKMOdKjRUugKaLsuDwRsh6h8HhG1ZhIxxO+L8ao/zp
HrB5vDqfC5JP9RfSGyAd+pXEp8h3TkHeMFWU/NgdQQPExcs5O9l8fz17Nc8mUPK0eXugHCynJzD7
c2D6+TE2XbUHptJDt24OAT96ZlYjUodsDiGT/D/j+6jN0/Mw/hUyQtW0nKVI+15kS+n9iE6qXu7U
VzUH8vHDfqbjPm2nwmFDvEzAiQVSiq+pDii9xlRhuN6FiKAbVluW83LhpdbsUj2OjzhnKTzXX/0+
RxjC1aPltHqqaJYDq36d6KPyQiUoLkXfz5dDAIzbCl3EFyA2KZX0Qe9X8iecTpFLp4m8f3v0zigD
RT84ZZfzbw11iqfHFB5Qcei9daL+WnXq803OdWDP5zHsLKycRjeKH5u3IJketsLP5+BNOFTzXfmb
c50F2deGpxFTFV5jgILHpRUREpKUVjoztQF2wty8apMQ4tDqR4kfdAPIZptD1/OS4BFF42K8x1eP
daOzjBIHydNgjUjQFpU2c33vpvu4zJzfKQnB9Zu62iLm/iFM2Xh303rJ+Zz0A8KrOSzueQeN6dy1
IINFo6NW3Zn3IlOd/r5as03Llu4wEKlZFBjsrodLqhz5CrOMK2mLrf5gZQDHAT8mQzJtqPHbDjLG
EmFoJyScfIERprS2YARtIrKBB8eCGirr0eguwbAJ9LNvKcWHGy8vDzt5varaK23ZsKT0yVaZ7kW/
D7c1ZfjTEBeLGxkqfirg099roE8jWnx809H5Og7HcAfselMQcph+7JL8MfztrVRmlaIUsctBRkkr
Vt2kT3KfKE/rwcYqDZuIPQumQ59Cuv+8sWMQO9mpC+kqnfiSu/Zp2TWi6Qf+lWVmqFalwdauyx/e
ZLPSjA+nIcCvZBnn/kri/DKk4suT1/GiPIaTGZruzNq6Mb0PNQCfIZ5OlZcMnBWqbcBRAx4mBoss
RHrMSVCKbMzaoToUWBHu9+a2eoISMI/iy2I6GU9UjaQM/NPRjKusavrrdBjvpVA/1i7glw02K6wJ
ZPR0h3VNBOu2jy5fPkFncGmqFSzDhM2HOGeNwozXZmOC5TUmYQiQcziAiSZg7BlmwF9ER4zGlvca
n0iOh40rLCAk7mQqfzMV6uiWbMivcwmlvhTso+kKFZg6pJnCNQEBSaxH+TbMAc3WqdTqW3yHyXeU
H/qbuW9bFPtvahIsaPCzpdHq1OZOSUFMlXxO5tWehg65TahEoXWcJLqxXHF3eomEjYB138byimRk
7j1TaRM42p4/prK81X0/tsUfSswFBN3TBU3oG0seM95xrXPP7WJfdIZpHrul7pDOOi3dsqNKrPz3
emZR0bPbeWsm6nGY3V988+IBTcti9oZrGAYO1Vy66H3Ol2DhmvmqMf81VFbQHuOzgGc+7rK59Y/X
IJ8xU3FtsmY2qHCtE90+u6y/ixyBYC5CqPlBa4V+RT2Q1eST5L0m1C4gbvNNHhWkqEY2GtFYnyl6
+saXYCeJOcQFP8UcEfqJKWSlI0pxejuYQUzXgEL88tBF2aQQrZJSjgdIdA7997j29fxukAnGkatx
JsDwofxCXyqEh1KROVRFyJlDm2I6H9wVOQCB7Ux6tBbXjVt+8QDN0Odg39RvGISpZ+Iynl4dwTpS
B/ccCj8T+TFHkX1tDHJYTYyaujlAJZS9IWEhOJ71mNgWXW59WQWpUNha0pjx/ks/CZerQLpgEYhJ
KiVZn8fTngWA0LrEQYyGygF0RGYi1B684q40PRPxzqyW+iacx9l/s2nFTvOUDM7IbJPDh7yKB8Ch
SKV5SaoKdf4QRCSGCDFqQNLyMPevPxPxFxEmG1i72lTkxSs1zgg1D8EKUDJCG51P5mIZYsCVPamI
p2w9LtteZAfgWeL+YAp+Ui8ju9rG+mLHAAX7RS2y+LPW1V1hm0pVsnYhWg8fwB81Yz1OoacKnW5X
gIhDvtiKr+gDbH/AZjP3Lt9Dzx+w8vlMgv8XXDzYW6Z06DAjzgNV4hAzdzGbgI2ual7e6QXEJoX/
OA0mzsa0TIbXWPWzBmZaah7vBJYcAAs1JKIBuBpSOmu6U29RfoFpfySCfIIjMIxHe73bdViuF05L
UNZqBopeyhwj5b74qUbFUHwunNE1tbK3gx+2k6RCAihmuJa2YecjTbzq+syv0dZ3ACxZQwaSfrJ+
fcOulH5j5xVcHs+vwp9bTSSkWnrO26g5fYiCKd/zzf7d9bU6fpp09oWe0txu2LIuiGLkUl40dgj5
C1wYeO3jnHheUVwkqPfjNHwS+8LxNYs9+t9VQlXJ4ghQSDnPFq3dhryj2nT1mGZm7Mkcfn+qjnHV
ZlZq3fEktGDEOHKKcuvCgbMygSyQEWbmcqVtVcNXQSUCo/JBOjVbornOdevhG2e9uE6JZj/fXT+k
qEHrgRzImMtJZozli5JaV6TLz4pY7P+EYSgHrrfwrtyVxAdUZQ38HLyRo+636CWj+OyrpsveV2RO
mr2lx7jOKNXox7kKu2stpy8qIxG1h/gB9eCyd8grCPtyPlpbQS3NqBZo2Ow2w6EWOwN5n4Ga0s25
wuojKmxr4rfRYuCqrvWIUJfvi6vnWCDKJFDPfuxUJ2OZQRFnnGWmEG7HiajobyKJCO/z1lmFXHVo
ObcXZl7AdjT/+KNl7PDVH8g+Oy7dNQ1tSshCX6ybh54v/stRn0wGMccITgs1O/NuPVVAV9PFIySq
LH72wqRv17sVOrDfxmVolwaPs7yumQb/zAAStlwx1QiRwNAw8ZLBYwC9AM4DS5k8kI7gx7HZ26wM
9tK7KKA0MoCUsRMc8CdT1xfn+vDi2EyFJZTNaUeS14Gd7Xt89ou4C+8g1y5f5M3H+QN+Vz7mRj1G
3DpMuVQq3h7SN6zrbjes5ayCv5FRcTU6J+QAoBF85MnXdYedGXJONKcwu6m2qC/mAnQhRyYIwTj8
LiBJGj8WBM6umADLpxGtRqw4PLyzepe9156lb7FTykoZuAzk/PSNos10039B+Ogf/cvxL/n7moB5
rK359fhMIQeJ3+lKNHHNuI5LAqnWEUFE5ChLnILe0qNedNoiRzmdTL8FVocD0kWBlGU0IM3ILZaz
m0rtmrUlFl+x14nZR5UBD0bNFQAF4V5f0iGBDHeo6KC4dvPZ2avftZ/+71TV/M9fjwyIOcaCKwQL
TkVueg4TYqrBsMblNQlx6vO+g5bVbBAsLqjFJx/ask3G/4SWTBEH7DtXcbTXLMUvxgHNOjcmTBXU
z0YW069XQ6IotLhLcCFzYpT01OFqE9YPoNAZCIH+sCNNbHs9ylaqarR/OuYTmzC6Ddrs+L6qJSXJ
JJk7uTF5wHmfq9D1/PRMMCLtJOvNjAPSTjlSL6QUQoyqXcbVy9IxOL5yJuUt+4TLVojO1AbOAwx6
PAIXwCsVb94FbdQNsMhUCRyft7C2EXTNrsV7PapUh6Vn9E9L7JstrhfQF6SjipnoHKpVSmRtaPyr
PgvM97ciQOLQcuV2OSRKan7KP1y/lgvsy7w6jOQrRudkZpLke3zv28SWAvVS/HK8r2VmLkaJ2HDW
OUttWkLsaa+VPnrhYhNFTVmN1zN/aguuz1ImzP1OyVHhMTnkumriLgiYYKlshMEJTREmqVV+vQpz
0nFZ3rNOra4D0Wch6HJj4ccyH65rlwxpfEf4m8L1+eyRO/SNAZsyqeqIORdpVv7OAyvzVWxGoN2K
2uoLrmROD/iTwvw7NuJF51z2bDvhMonKG+SfxSm7A5prXw8rfg2eRb1i0G0Kk7Kulw6I+H3Ml3++
P3MNJdD2UXzaVSYA2d9cIVLNhsc22bFFU9FYN63fQ1DaP1i3Jf1a7lDFjh+VU4rn0ecdXB04JzA1
efk1MgjkmKJlwD6D7t4HqNCUfIKwnzIn0azuypxmyV0RIM6p7ndeEfbYtRFHup9pGMg+kVMVuNjM
bOR6h241JCWGdZEUaOBliopQkJHoXED1KvNUxxjaB8Joe3cQMLvQ8RveBvdJW0Wab26KK4YhU5/m
A6Tw2AZyyNzf9bxTs7rh1LUr+BH/h9+5yhgCUDTyHbTgi7Y/fClxiNYgHxW3ERoGP8neHo7rd65Y
WqjcEepoLptbbj63MR8fmfvEfeCaIanbJNI61lazuP+MHc8kMtNp7EzBtaCd9ft7Qc+CXFsE1GPL
R9yM/qwVpKivJdClc2FAM5gc8TQEtL4D/AN4vuwajdDJM0UTUdQRVk+mv7kWpRbzMjtMCSEmCKsZ
k1VKEJBwpsbGS0DL3lzZx5HhpUNYQxFaXLwOnOqFVYgIDfWYpu/Ga40fRS4LE7bp2SvJ55tHXiby
FGU4ToCVWgHjWVed6eLsALudwgDfRiXz9nptq2mfkY64QdeX6AezOKaJEdErPgCFqHf6zso6zmht
8WUXK9lJIeKSh8cyhx3Ys8OZ59ZAb8bUcINOK/6jADlpJbuw/GpeoTBM8jQ98upGLjnNJgJ3gMm0
zrnLNm/oo0zsa1/gtdllexs5bkYGqJdNcF6d3+ls8KkLCsRSKGTYVIWBVhiCUyXiynPd0auKCEYL
ZLAIGGLdxDac/dC/YO0ludF1PEnn0lBUHChHQbq4VsX/Vw6zDfXkThjfLZ+ZuC1IcK1bOAwgpPi2
l9BRtbkT7DJb6Ng8UgC1QUJAg/1Dk6Xp1AC1RehNOPc9504niXpLd/16TRpQy6umofRiqN6r4E9r
bE5XMR4sEOBx0t4d6qEMfwzLODKmIzsgjx2wKQhS8qpKB168E5E8Ds9F73FUCupCzbsVmmQUilS8
68ZypJ6P9jizK5DDUvGu7k4RSQNBDI2cy95goK/IZxwpoxW9ImyYIjpkGM2KNM5sF5eGg4Gupnrc
llr0Q5azHHV5wzSVawOfJKdTl0K28bp6+cCXt4CRUKnGeAoIeh4oeYP04p3zpnaP7XkB6K6Q3fBy
oEmoUfsv/uaUmiVyV0bxqW0LqFpZasAfFz46RSB1ZYBUQ/Jysfk7S8qvG8ZfTM2ipJUg7ip6Hiqh
Dr2Cmcf51pFqCtMoHqX73L3Tl0LunNOdOkQ2hdyKAlq0exVOwH9cHvTrkOijrY/A/5RxfD841+py
a8dKNjHgJ+5VApVPSq1vFJOPd/iRZaHnm0FWBxf2vO86M9BESPUEvZtooe30jNSCUEAzKfN+5NVc
I+GGBBN0btlFVBTEwe9Rc4gkXREygGI7c0TR0nugVgra7UqA1S9gZi2rC+k7FTCPtjlU4PGTpzAq
RkSt9F2m51+xqgK6HnsznBn//NYkn3b/ORx9q3HSBlvsDhaeJ6OYKZ5dvlRRyhUj8bEkthrO1R0K
Vw1pJvIQ7V35cbE9BEEDKBGxT7m7TRcALEs4EqgGbyLsVtQH4Otb2qMYmrl9z9MgNTqNeCi8nyGk
uSGzcKBVT0pheZLVGk8livPHq8goEIPe3lE37Si9EEUURb44PwLlMcbLJVQrdnWBgsWaNFGfCa+z
PWiwljL4BMSISHxxWok3scnpgYJZt9ckt1xvt5jMhmQxkDwLXDsiO2A7xWh41Y/6gPl3hrXR0WFC
QueTslDymuwKNlxRr+XiOdfgHxt7ZU2/2kwzJai4K++/NuGqcO/KG1Uas5PdyJesInv5gFRnKvTH
8rReqinZa6p7oJ03fCEAARDcDoGMYzJdMGcC+H/Yz/UvGR4d+tXg5Qds0EtFkvwKRRzCQ5WVKPa9
8SQMEDF9v/XPKzVYrZabQkSyUgSZJgJHr/jO3xhUGRnruHuGion3BKoymjT5CgECmCfWDM0N8vUA
EfUBK8QZ/Dx670vBk1g3OBFfz3zLkr940R1c+SrlQwsYC2DItMGGLVUh8krmJ7TTtqCiOqDK+Axn
TFEDXpXkapa9ws1f3fRiCGVZ7xBP0GmFDhwytGUro8INJfn44pfLq2W27n5K6GvCtxbeN5+XF8Qg
Mw3RLifJOvaJHcFSqOGneJtZFxeXDWoNwoicGK0QWb8coqRvYpcY/LNkr3CMpx381UyzLDfxA833
UWl4p95we86RqZVlpgHiApp3Gve9NCvctxdBXhkUYTy2AxUKa8twQrYTaMXKDwnjGvndOC7OXAgW
dY1O4lFRrMXcMWCXF5ydyrh5YFFhdrFsl3JPRnd97Kugfv/VwcK2nxF+yJ9UGN3l2sYl8ZnG0xo7
rd9VWT1OTuTx9IYp+9A2fYmajNu9C3/dsAsyuiOVCe0kxuRhltQtsCc8iV0OcBVGjK6D9Ko6jaBv
qHqDmfkgiQTwZo14UQHOgg0b/RK0EGe/Bdngo+Gq/bZ1sdpwGbB5PY0a4LYr0yl8pQpEJNC6uTuL
uUCx1WOZgmP/FsAzOc7zrl00t5FkAMKrQ4Pf1ErixLdRCkVEBsNM/u6Dn3pLRS42xgSbzD2aSNpQ
GSh2O4qOgRry7TV7f/7Hhp6XXTGi7nKo40HDQCSC8mWdetuFTJVf3sqyqRS2zZgC/gscV5Z2OrWa
tgRBFei2AGOwP8VElS6415eiKCQc8FUFQMPx8Jw9nlzK38/1n5NP6pLQL7t/jXZzrWfENQjpGJnH
MI8qgTSjLJTImrjKLNl6Pbc4+y0lAD3mbwG9iFj+qy/apgGIsN42iTh7Xpdbpz8LXcKloyd92Yrl
/IoznfpIMRGYVZ2Cvh3pEtr/UPfvJKMulOSK88IzZ2CwpVejq1bS0hrcYr4CqemzS861AleNchC5
3jKbKbID0be1SHXS7V2DHCN3fz+3zZncTPvDdFktj3L5jpMxHSOz/noIQGror6q+rJtAZBxrBxVq
UnoFwJ+SJLZFhUQhRgz5CM5FnjADtlbDfuckA6snkGAYCuVUPkrlz63YMnWRX+gUUeoVrZaQ3e+B
jfNN/2Mw2GMU5noiN6nvOAB1q6xQl07kI5lNO35pQdkQdxveFLLbNLOUkh9eM9aGC/e+2Iy1UTr1
Ela2YAA01cRrg9CXfacTJRr2GKsueNH9wdgFxlaAXyjk6nBP3z6lgbduF2A9KFVSFHgqial+gO3R
450GWMqp/POtzBuv2zYEHHqptxQ6LeFUiVHfEDlsK89FsQ+Wbxok4QhcMYSGB9jxV1SzMLh8NEEw
Kz1oHI81UyQiD9aFjFPFGik7rjsO2GiKXtMmFpoBKwUXdpBwPWPmZG5kyhiQ7EgPKCBy9aF2M4ol
TvkizqME/gksrhMzWr8ijO3v8FsLutNYAs4y8t2+RTJF/OXI2aSt0rjqSVi3hdwWik4xgFdDWLn4
caY8ojU45Crhwt37xUXdXdNg2w6f6h3gIAexAzE+deiAOySqDnWJTnBViVeTKYZWdcNYLXtgDGz4
Glngcvewd7jHHEawmfhwZq5q3pQzbOLJySLvHV7aCsS/CkiCAZFKIJmdSHjzGtsK2ydkrB+86e66
oiBCtlyVX9DnwQx3OUNl2OtmVdndFNwmHSmg6LGBO9hR6/SV51pFBtpdYBW0ErPg1tl6B6OI3cKs
Fcp5hBgsTlFfhf1rC9yKFkC8XdcSer1g8TfehoxX7OyVXJjvUuoQ7xmmrHCf1u8FOFyarGhRKp0o
01iI+6gb5NSfV3FuIxoqYpJD2cH7OXEQtXIthwYCGrRNvbshvvLkP7HXGrqCJ9P5/HzwSd1YY6B8
3LVytt8g/ppgQzNTyq/nGzEmKHyyPNbmprTbp+LUIhoGw+VRTovnUaVhkF8V3Gyd2tfaO4D8qyT4
bKcA2KQW3pfJzFluGI0wI0HkgAv3zugeY463T076rOzvSdybb40l6qW+s9GMCt9YVnIhk0KrveZy
utCkfRb8potOVmu/kDWt6GMqP89AXsxIzRVjAbyO2bwTL0GR2M9o7tYrrSjLoYSsd4RbTT5xmgNN
csah77GdL+s8vNL3Vl18W5m11r186aqK0v/uouwaUhigoGML2EKFrUw0vnzE0HLf/nnNfobirdho
LWU+dVDeF/l0KRlyjTbpVEOIq5pfH6v/nLjlOg1Rt7ekqMEsxRU+w/jE6lgMLWKlUSEhNXehN2wU
QUjosbuR9GXuYcmCqzV3Ga+pvjyXnv3n+66Bo+cSDmvatMvvOZCr0x4QflLZLrNmUFon/duX3tce
j1WYpW6EKyfmwllvcy3LQo/shjbabro4IYeULDsG6cjh7UQ3iK/hlSlaesUsJLl2gODYhX4MJY6m
kDPKMW9SsNbEwL8wAc2ruOTotZOPDbG7005EiFz5Y1ymeuLqi9DLiNAAVMs0X9GNQS3s5e0kXpvR
wEPPW4+gI/yr2A8dOQ8HpmsPuy8DvuSCG8MeoTTBrsdI6nIuVaBkqd5Fmcb+Bboo/w1dV1npLtvg
VSKAQQBFJQA81wbpYubaWbeOJpy7nEkWOrP+Itr3wiSmcuqRPq9M+/Vhdnn6tBPdbQDHlOATZ1Sr
wapXU+cVC7qbNVfIADH5ntMuNWlZwH5Tw5/GjVDO9Qmhpz/zJUenpdVfMkJQXE9ksVMWswQBEVVl
pxe0rz8QZuQEaBP8fM/ZfC46C1tQgZWosP8vTALkIypyWBh2g9Z2q8HDpG30pvUNTDRJFSFrAlJ2
/08BScG3bH3XffOHyyE1jWBP1m3mHbPzSte+wYtcsfLBpevzTETjtARQJuDgNKmO6I9HSA7W3WBg
Gzj3vwYsbTWHQpEfCSgPVGl7Po6YqrgYvL5fDJJdEqFYsLWQg5YXHZCCBcx1TXiRUSAztSdOoC3u
KDsjmy66RjmS8V0aaBLZ6dhqnpDUSi8MP8gur7wuJc05MK0kGVnHi6yvK43eRVqM2JHDRX1nJ3QS
+1DcytLu5DGIeUW8XUvd4iEI5Tdbdaoj+0ivbtdKfDGFhy195tGy569QX4DksU8V9vE25Hvg9oIj
xsum/NVHVy72I3D7CSNYn4fBQn5hlFSwokxWyTgL0TPLqQ4BSjzckduZogvzTMrjPtGpxRMh3hbu
eP+IbaezKOG7RHskeCLI96wVVTpZyMy+yRGz3MeYOZ1sO//ZsU4qhL0cFRC70EFJ+H3s01FbHf+w
X/dLD2SQJWGTv/bfqMl9mfmYftgFyjikB7oZleiRLXbCMfQaSiD5myUIiQsiAeHOJ6xXLpTPxrKf
30yoJeF3zQI4q/xHP+jqORvZ0v0G80jnJiucNMVb3+Kq73WikGZiHQdKtoEkZ1HtTR5NFMS0bece
hDUZvE19ZBGm6dDfS8jkdMsYi617UQjiuC431GWrDFMRFVJQrvmy05NyX5ScgbX0uteqdTlFrXTs
AR8+zqLu6Op/hJLuEIPGhA0kbhI83KLCF36RPOJmjF/3wKUE82W0pAWUhYxx/GJg1+kCCYk2KOr7
3VsRosVGV39IWiC+HeH4ndxK8lYzqoehaP8uxNawLMZtFu5iIw9ipokPf65hEhXUchQaj3ikAXRQ
X4knBBUzET08LwpnudSsQAXUotVHMOBfvSMIZBvpKCwSW7+2CMOdFKCjr77G1N/d5FvdiEheDNGi
Cx5lpjFzCY5rKtxTUZCFa9fvD3xKLReXyLDPj7m7UPTLNXzFI2IKutI4OFqQ2yj2sm1pY+/A63tH
PKLx4r0CsLG/eKF6Iifhyh7eSD8bGfcI+ZmVFK0xLD9gfXZcyu1VP8WHsaDyDf31A7Wjv73jxgvP
gYkIvRwn4L02TAtdt92XYVtgs2u0waEV8pc/gZfBdYkXqgK7ejl1e9IL+HUKLEY0o3rWjKsfm5zM
i2fWMWz8NtTBjDZpXFhoj/DQ7pjOCmxTquabP48psSiLbzbBQSzXfG3/VqM/nLB8rnux+JdZ+7xy
3lQZN7Wh1XpAhaCGdcU/5wGcdF2jHlvRUxTlHWTNHc+eAaLNpWeh7ChWRIOkQnhWYEIDk+4v7+m2
zW/FnaEAaZ8Jdl48NPNkplHcgltmXDXUPzOe/Y18ZU0rWB0l6fOnHIeP+C2ohaEerSoF/myPmMNL
e6o1DD8n2vawao+hDnBO2JnyuwnxXkfvll2+ELRQwll6bepwTHZneD5gsF3o0V8JLa+OS6x+SL6x
+bVUJI6fbEIMxMw6yhpjmBKbYleb/PYoahKsqz2DaHb6e7zRXU9oGUdUWQHHAwnFcLXZs031Uyjg
2zV/cCz70aY5h0k0eFZXLL+hfFzcVN2L+eMv+qYjMk7+0MIr/sfXJA9LQ/BaKLAx5lzoNtwOH5VV
3PSEFKEsoQiOKIVdp6YzJAVBxhlA2rv74qPgQaXgUvAg87GvyT6+ig9KulGvd4htRyr/02Y4BgVu
MUE2LRlBN1VBHdm/Z8nvE/gWHW5zKsNIDNUgC8BqOs0vP0LR0JzheuDzc3tCqJoLC9ZbCQdzruKt
EOfueYRP1X4LFIDjk7HmohYiN1tokv4jH9DGRmdz2P/k6XekmwIrwlEtQ0dx1ec393+kZV3yEw+G
s4MW1Rj5JoGXiAneoUMA7THXb++s6cJ6hM/FtgfdwgnJ3pIezY6jDuXoxuPDUKcpFaf1CUNjr3/+
IdjzaW3PYjDhUcIY9+V+Ojiq+B9XCjVTnuLkAzyk0fmWKaJmJ5Wq0dtSwQI50cL24TjbUU/S9dkJ
t9eVbt4Il1aTVV9yU6/mrpVCjvltKHiQwVNzhqMzWJ+XYiW1Z5SQNT3V9Id0YnwrghOI7TeW+wv0
jR2bR4NwFXZZIgQ6EC7BYoPfXlTjhz6rpPL4n9ktB21bkR0MMlOv6+qkEvr2i6xWC+AMJ41RQO9f
BjYQupF+TUTnEFdP7LlfTWtjJmhREE/zvCpK3D0aXMu0CyY+Qx9eUOLOm0SSfl+enIGLt7LARPkb
ioaC5anIleqzrxD19ETsyeFgNUhhPO1BTGn24Cai7ZjnjMkHoqaUadLShCH6w0TyNjrHuO0RJe6t
XtcR7BPoW02a/IwPIjSrAfDnKIzDpwYsK4O5BY+K4Blr4OoJ/RieBLCMNx1/0Ec59/p/99i6Glcw
Cdb6dOVGoLJEAF3pBkPU9fHOy5/BBy8nPN0uHiS+mzh1mMOg+7oSNCzbLkW7OQ4Wn6oMASeRT+M/
qHLz0bEaUb11aaI/gV0t2vtc19QLH9AEzdIHHzQW/7Pct2OMcPxq29HXjZd655UdPIeaSySb6tCC
BX98nvYfw0C6Fxmy9fQtz60KnmdildRaVuIvCPeQU8L7Fn5ejLvnRrKcX1mfubpvT5FW+Tvrk6hS
urnk9Szo6ZLnrcNv1Aw4EVVCaz5R9PbjzUbz4fi0XzVukTA/8zBXUIQ8vSI213CnpiFBK50HCVYp
HJCY7klwz1vokjT9u0RXBdqKBK1dTJrbRBL4AnKz6Z6lJUwaZbGU7cGX9j2pFCkynVcRIyfPgbd+
sXd4q6ZpKjCjcdqNWAd4kbpekb5sU/nluTb0lWvVl4xzyErOm73EppOf+SMYeR7BPs5Y4lz5nGGi
VrG3Yc2U12aZc74guuoAx1SyXKn1QS9D2id6z1WMVWd0rD+nTNzY8+Ofz/Ynkp4FjJ4lC7owQIRP
tWl1aF8jjFcEPcAv1eX+GHTnVoMDU0P3ZhikN3ol5bOJofcdzymYRbjwSrpspvzDMhHei0fYLkF4
fiRjTiRqi6/cYYIzAAxaRX33O8tTktErSVgqULHnu7mEEvKMX0WyuMo0lvIs7pQE0yeYEgR8BqrM
8A2Na1YMzRl0nf3u+Jdomw9grhWFmHDw+3SraWsjTzU3rn6evEKO+Z5MHt4lyM5Hgtyf1ZjM7S03
Ywzs279zfCbItbEmU1RIlYTeiwE9rjK+nXBjxi1+oV12Yd8WPXvPJngz/xH2I6GGkDL0qXWHxkos
UFXHRDTgGSyhElsN+pH8WAdWeXHU+Tm3E83c59p1fXE/XvBNWfkE21Ukm+RJ8zdrSbZsmrjBxs5T
2Ka7yzXhsR1lBZmmVzX36E4CrUlhTvcjkhB2cfGbSf3dHBiDH6cn2W+kPLMnxzX3MGlmWODBKsNO
kM5ais+0PU7LSRPw0rHeB11n5IdNYBUkWo04s/cjZ7o+3EEkUnzqA9uorrZgYVpVG70liRTyx3id
AUP5v43TtCZxu7XwrmnKCFDH2/IbgmWzyWdnxJrX5LAPcJ4S7CYA8ievekcKD9npbc/gidSG0mBc
ULvKaKkLsboUImj7zQyASR1EAYblwA0SrGal8Ar4dBi/GapibGiiAgu3jp3VtJl43iT7/s4qgKhY
3VRQyjIAoYMpe8jFl5AGjSBz23zKLqSikYH9kSHxsKqgEOj6n2RROuR4PKZWJPYwPwoKkUgQdw5F
/XOc3HpQ2iovJPzF7nweoVQXFGh4IHOSCPbG6Ri/QFv+8bgzdIRIzb5lHU1WtEuciPsHhWtkrBLw
eCWim21wMOFgIRJu7H5uFw7nWmz4muPv4dYfh5f3YNm18BiSzqcXGx7J0TqO+x5TAwTIBSsdx7Tc
8lUPomB1sZjPwjgcw84FG/ozwoBF7sJtNzVDDwd9IwKOmOG7uB4KdNAa/+psYGPEFUrNyVW3zBNE
yWNZtUPHTVGKsBPMUusGWrLWNYYZUC7T8wGqU74vtFWk8rHJdgi2BbsNFOA8u6MjI1wEha0NFACE
w93JHMX+Cs8UG6FAMFIV9a76hXmJb7z6YqZizYBNJxd7XXyTMpbgypQT9x4ZyBVW7S9r081HhOBp
EDAxKhB/u5FRPUNkM2KaSiSKi1klhzXlIntJh8A+BjRfgZRCBjmfFL+5N4SqkcZycYARHPGgkBiq
rl87SgYCymiDpjJNPx/ldOljydteEA77SUm+Bnu/HdFt0OKfVEVkFjfMK18jJwH9go2jSYUYTsz3
1DXxz2nUvi/X4yW/UnHFn8mppLDnhM+ToJp7/GyWLZElzRBwUuk4/9Cl6mRKB0kxvLXclnReNAwI
fp07ysWv50qXbcdvljcZRxGZ1BNhfrcq0AEU7FvahbBpqmC3Qzgxcu9gCXwVQ92MkZ0cx5S2JL8J
RrOns/H7+WHRtoTt4PLebynSxQYo9W3Gt5UAZTPVvyA1AqvDU9F9r20LJGBX/N2OYO7V5G0WM+ci
EVCtPVWrjMdEuJnqgZwNtTSBTZN1D72OE/lc23V7J6VRU11MbFGnHrWaQCMsssMjgOWl9vhnR1/2
Bkz01yPiaUNMyM6+eZcSXUwfAOPD0Mt8RNXpwtI06Z4HPv5gqd2yRLdkcn5+euWUBG86cOAFBqWQ
jmVJSJI8pB2/5uMe4XuKZoItVcmAnymuKdlbXdqDZB7nd4ufIM98E5kP17YAyL8mp3ofDRC6y57t
RimO/UmvUmPhVdQSC30Gmqe1pkuvqkq8Azty8JtU8whVJkKR/xK4L8RpXdH/YpO4XtnYXOBLGWX8
MSEPRVihimL93bg0pe4E+qebmug6AbixdPN4cQ9ogJfdh3yvP7atj4L3UoR6yaov9Q9alg7FGXo3
XJW86mxvht2+plz4QW3K2xcgqas0xPmfAorxxE/6IuKX7MSiHwYqlx5geOZIKmJofH3jhrSqfXRN
zX5tL4/Om3Pk3bMKXbuQ+Ge0znsoZTIUa/fx9iRG8Jv00tIEXRugC7yJmkleHqUszKrRzGbdVzhl
g1FT+rYgpVAPDPRrW1q94loXqRxs6bQhs22/G4bnpdz7XTHvyXNKYetF5n0OkoS02soGMG33KlR3
QMSWwmho+vA+IxatsKniLXmAF02hGCmQhCBwHMrzT18DTF3uXwM9VJX9mFe5cWY6fCMjghGptv5n
dnvfHY6hwNFn2hqjqmBdPkDcenH1s2y58I+e6ey9sHT21BZttABH/WKQ4iTzbdUhNJF8Z+X0H58v
avV/tVcF+tvo75Q6eYB/f1ZFwgOV7dImKnahhXhDQV4Ljv3cbKLv25iXMZ071IlVPRLGcSIyRFkr
J+IIPfJGBcCq1OQKYcFybagtgKRttF5AXRsuYkIpVuocsnGuZijRdn41EfTtQmXAgcr4Pw/XX27l
S5kYc0Jv/lCYwDImfytDdDI0ZYkmTcp5lOcIyzHLUhW7QHI8c6J6tucUmxiaK6PIS35hqGK0rao0
RhDAP5V7/OFZoeqD5ciGdpE1SsBrJAwh47bks/bTeFXRMJppWeXbhFF6telSRCnm0VZ8uN3hz1eh
DtnmQpIKrD9df0ifSB25gkqX5XkbPds886pF9qpQTDqc/YmWpxcPVIk6q1CyhXsabBugIN/GRCQT
AScV/vhR6kd7XOKqy1d8E36mfHP/nDHjDR0Keofhi8zCS8pg1GvI1B9IssqVtvChC7L1uIMcXnd1
u0ICEvUf6Cs9qecm7zpw8cLGR675OzkCNmYKNjoLmdpIpJJhsEoYpcXzJ7HhQoG6ClswVClh3q8i
ts6njqIKYl8WwhKhjDI2o45YTKtefQVy4JXPC8ovtqjl4U/39Psjc244Y2wC3NZY1/qkp6335n7I
HN7dKQc7xaL+biqx9aY77P6xrnrVIBPm4H63hopAZYOY7Mu0m6ZyCYVaUL5zEZP/xCw6TSxuK3zW
Q+JOjnCDi3tvIzkm9PtBAdoqUpXKrlKENgMVwVKL9U1KXFOzOMaTd48nYlouMIXeXFZ72MJtJVLs
qYq6+Jf94/QEPySs4Vl8gm5w5w8qtI0ejrIcdDQzoLYyioYPrBYtTy4YRJ5hqeneGJ+B5eh5PBOK
iYunBnRLsXCNYwwOG/ej0fYEUTuO8ht5btjXQp4ZeJl3m/ZZb4kuXMiTKEd+JWrFHSVbLNOaGD3K
DVSP4V9bpH8zqluJLhTY0k+QJyDTWlIqZwgkMupwOvDrsdBMaKPvJ20G+daSgB6NiMcM0DT0AHFG
hk8HqHym30en3AxrgKOm6WJ+Y8lcuVMUzlttGy98zXycY106lydNjJ8zeYXitUOe3anAC2bbOxB1
HepA/I1LEl3i+nIaJeHj9HGqRrpkwIySl2ymvtkpSQhDnKi+nWogZxmIgI5KRTyrR4D9v63eqPRr
VGGKT4ZLJGSclFdCJfzVCRUws54t97mGGwfwd5S2KYYRwxRoA8EMzsISyyauF+ensDmERV4uudtb
El/WkwNY3uDB/0UBEGRsRsvNYdQdIh9p+Sy597pbh/vZiB4kBul4rnypjg6NNGLbd3qoBJuzB8c5
gAeoLew+io2hqb7DKy1t4+wmd2N241j64tDv94VsE88BYLsxNU1Nyy40T4LELMs2kMUggWu5nzfX
sLNZnvqnRAYq7ojK5S4XCJTfhZAr6dC+0wmn6pammIXapDGzwKHiARSFDF8Sp3qkBXy2xjlvVkwU
tU72+hoIt7wCQoYiZkJ1YDAz/8LzCOk15iajVXD+JYrF83jAoPMkeVH8Mk9KzDVMx43bgYQK3/6V
hsIkOmW79G6Dlv1Vt3NwC6N/zp0mxUcbbyyDSo0mJLGi8JECnOmOBZnhPfdDXNmYUOu6lvdWpOJU
to2bM+agb6eWjN2Svb6heej+5PieaHGxwOsv3c46rhV+z5l4E7N8Dzaf34X8IiYOTKVBwU3ph8IU
2rSs0nVYlRCjLQEVjm+l3KwAIE8OOxgDf9NFmH/61p8GLXJ6LBV7wUaNfOCF3iOCX5TnnoNVQ7l/
57k87hwxfvsjZOz/pLrOf2UtuaIbun/AOf1nqUkMY2yZgbCox3tQOPnOYN0nODVJW+NAsmnCZGsv
9NJ3hoih+iTG5B01MOIARrVi528NHuvsvcWITcMWLwCZYzCB7yGfZShPCYSCzfTRPyQE0AJAdbV5
ZxKb87JXSLmcn9hGjI8dIyTVUAAt5qMRw9L4wIB09BL92k4Br4QTUrBaTxKIF/DXl7RGv90luiQY
wSGMpSks7jwNC7cDT+bJqrWrKuWcxLDzJBq/cdeh8xqjov7tpt536ujwklVbuk0deEzDvszIrfbQ
pG2pGyJXYQjJXBxSo8SzZebcGg8OI59syq3gCXd8p7Wi31T2GiYVQXFfkY0U2B6AhuohnIsH5Zq3
/UqNH9rIIaKkrKltwhtYnMOuWx4sRgyettEFi0PWN6yWyKJ5v+5Slw7F2HyUJbBo4RFSQdvQpx3W
ncx+nfddhP6sMGw4Ah4mzLmo9GGiCE8FykVfjAWvRpVsJvah+OfKKAD8hmbLAVuFhyOOlz5l13yJ
wKhjA7BpYAjg8Nkcflw68OeaxbQP0Z9bPCXJ01R3fNAX0dA04nHv0tT+Yw3/BkPG94mKKRP3vlvv
cqGfi+gkMAdzlHYAXCr+MrmCW0y9AC7zqbaMpfYxlsHV1tszoUzNSUYMaXBD4TkDIW/2Z1Dww7ZX
x8OUdfyo1VZRk9IuuGt2IhCzK0gF8vXm+FOlm5fIGQfIazisXqBIdCc99w62pehd0jVdSxWQmec3
Z8AzMJXjDcqeOSAveyvi4DdHbGvrIiGJRzq/jIxyj9MrjXf9yYl8CaFqVtGVL7iMlJkQT7p3Et6l
nj7lQREUlVSC8v/wuTJCHo8Z50Oup7zz8qO7IYwQDe9XjgDmHNKcEMotLblinIXyI0DHUrH0EUAz
/RsEkO/jVMHrly4pm0aDh7RWugKRr1bu1B0d/Hgd3Qy0XaypKG1zCSRiWp2cUMoeH7lCreABjI9X
Y7IwLhUokj6VH24Rn/pzvQ6iFI1b+QoCYUFsRRqpar8/Qvc83GW4I79cpXtHDvroS4ImG2+6iXgV
87W9zrL1loK9tcXn1l7TsTcGxduoeuyEn2LNCV8jYLX9lx4+QNCLDn2AnBupGZDIx1msnwkSIDjW
e/GlSbWmC2jEviLQ5Z9wevZad67pSs+a/5EScuQ6N1XeRTMOEGgrr4rfPfP2qPsMzOABhQw38kYE
FrFAhx/IBIPiH0MfVBkzuyicwEauRBRLpLXyUCRHQmykPHTjxe9ECEFiRHotiDxZEKsvngEsbmbs
xhiBQtKRjj/AJHZ3KPIFOnbYdjNk4jAnDle+C//3K5schr5yiBU6nu+eM0ab7zlf/6Iza+Zo8zTR
7YR2Zog0m44RbyXwkcDNCgiTTkbgjKvBA0tTDFjDpKBO0ddj4nY4N/528C1+jtSvHkBkd/jcBEZb
noARqgVH47GfhYubM4K/QYAAfUqsziGX3bq1JhsJ7qiD7onBCkuul5KvwIpIQudZEUsVF7PHwJz2
63qlsbN8wYIGm3cYyuKRVn+N5UFgjX5IvmxosGyuJ7+qEadzaOCMrWIPZrdYY1dnuOpm8GttVtno
c8lQG7/WgZh1S3CHuM3sbfK5F2ZoZI82ESZlm9Esk0nyLk2OBOPRo0WGBAAtWowx9waXyi9CcItf
Jnurmuh8sdR8X9QSFPI4SypfmWz+Nff8+cSd3gyTa5gzDdbqiN0UtOxABVa0/0LfoWw2oK+eCuvQ
exf8stRKHfc/+kAgpay+2LjIO2fL07I3VS1BnLcHHadXxYmMVMfWZ3/al3EfEB5YA7xtaCinbk63
Xb7kF8RBFKN77phm3xGVonF5iwBV0jch9jD96P//ICQvFciKHs01xbIr7kspFtfErPUm/QL++l1K
Fvm2PufCjN3cNYv+BWiaGhZ9LxK7NAq7HsZevQug8rKTCEcp/1tmy95HH9hI/AT/y7jhtzp1h9Wd
u4cvpBFJRIxLlfk6ULR3yA7sw/PoUjuvgOmdID6A6dimP1vNvzBn66nQefJZC135idMY1pKC/PIi
TqZlXewrmGWGO9DGc+tUsJjkCE/u77dSnfOw76kJBAiOOXKh93wr19lz8I3HDnniVDbZHufQllxU
VSP+3lBFaXMxPQg/BSYpAGSgwQrIn3unjA65fqagfBLFOb6On1RbyawIJX1tVWAgKSQBvhZXd/CL
5Nev5U/vSkGykqwznKDJYPxbHjhVO4C7WI974GAN2v2J0/4cAojxCxvBDpoE9N6OyLujnswlfvGS
st5j5pmmaI8O4fFrnNUyo12uwbVQ+vyhnY3yhxOwgYBPoqxaqxgQSzrWSr7OrLz+mOMMYGdxeezp
2pvgn5e8rcQFWTTpz73X37WoJQuj7bYsMWC+9bTnHlWRxPw36dCFcl18KHdAYxuqVafqI+NtE/pM
+qewGbtqt4gfbGHBb6GQusaGOIaOTrYpq8Jepuvl2HWpl55xM/JFzizw1BIokzRl7lh4s+PDrVMp
rmC0CdGdo7FVrwShs6hRvW3pzniRsilm7cNXpAe8WMiK4aNnaTiOVI+69Nl6r1FcdlQsXB7t2X6M
EgaDE67SQM0G37ohSmt1uVqZ35s8DHPv6CvVQ/NJXMR9j82q9HCqBUqjPKh79unSE1eanQDA8Idw
peb5Ehqb5wOxgTvRLmNnF85C6SZhCUm5vB1oedXBJ9quofz6dD6Cj59QNA+Y5Ra51v5R/gCxhE6L
eISp/W4GPWJ7zFakJGOaAoMvR+AixXyr1VpFDfm3I5ZkaAxoUpI4nYqUtBXH2byolsPbGGoTtVkY
dIJf9GEL3+fjsrw79QjdO3VLRAp/RO4aYshUcBUg0Xj0fnS4bvzpiWNaDwXUUkFDRZz97yjphQ+H
by9RNPxZDYABW02lEruAYw7btKO3k0iMKJzDpKMoyBebr7a5RL9ymPBIXMIj45QEJsihv4ZsqxaR
tYv1MW41Pcryt3UG5ATNF0uybHN6EmBZT+PoF04cRC7fVKS8h7xceY0xRzsf5a/RhJXLDPGugtNA
af2h0QLcty2YWu1+QqoChJ+iH5YyHpuqetja5MCoIIyIej15+r17XtT4u3/SKpiRr/ZkUJachmZj
jnL+D8z2utZbU2kV3Al8EKNtCGhlH/LVBbgwT9HNinrwRprjhUjXNev9YfV38ZxxGqtR+7ryFXxn
r9UMUwL7Q/kFDNnC1+51Pbwd9K2cipeza97PfzR0C0vpMfQbomGhLTfIxWdbHeX75rBSLOKsOyF4
wi/5uP6hJCO0viJaEhyPZZ7DxIH1MKSOoXH6kLTQFLX1gP/iX9UdMah6AS2W2dB0GLzdpU1exMY8
Bqg9NX1K/48OHOoByBnAH7sqS7d2/WdvVdHxzRigpfsR00PBA/jLXe/Ia3Hvrw3AoENQhpr4Hp8Y
HJQsdWfpsoxY7vBMuEr8reAVH8NLc4eCw1Bn4owmMg09peqWlrjgwssJf5HEe/1VCJSL+HtdZKPX
d6dAWuDXuWF9yIUSiqzGBWpZ62uyw+aLUsgC8LXhFpj1n6hIvJXCR02HHXltMymcLxwFsdK135Is
sZep3wPkQb6R/Qug06/d1UcoUSLJsF2FjHdBUw6G22d0TW3lYXh+KFlV1lUD6Si2ybjux9U50jLJ
+hnHV/Njxp3PcQvjR3KWRrTJoqeTfGxNE+F6W2NyZ1EVSMkb0hhHnrcdlk6xPIVfWaGOoegb5YKi
rhQ/ohO9dY4thgsjPDZEhZLAe9CF0pDLQm9rwQEcKMQWKgAVfCOYn4qo4u6sM18ZzPNQje3iW7WY
W6j2j2b6z+ITIRJjw29801/6zlUCMMS//MZJbA2RnPozNhG8tny1HNX2degDusFiY4EqEWcx+Lut
/eDEpF2y8KI/JW3MWMebP8Y7Xi6fgrlJEQfYaiWRkCjHze/JTvwNF/JVpUc5qp/I4bxk91PRHAE5
JB1fjkGA+FO/WjjWqau8hOPTB46y/p/2fltJkMPPiWZuC0EN9YiPCKX2nnmWhqs/JYptL1cjEtXr
WFxw5N3zS1e+9i4Yv5qp/7bHfY2QlOTFbNtN60u1Oat/l45ScJWYN0koYP6F2dqpU+7R8HcE/mdc
ha7fQLHuFsMGJ7epv95x/okb1Yi0eGuWJEFPaHd7Sh5sSUcOLfjNE7N5hRITUywaZ2Fonf3iziHS
s2rOONO75jqfKkGPyWRDiwP36tDNkZvI1ad/m6JBgJXAQfk9pBrepZWneMK5LsHGqUIhc0uyH/5S
ufZje5GbZK6bMYqccr6iO4JU/QFT50XbdUTW0zsC/Gj0NNJz0JegEoNnHTk5MmijzykjbXI2UcJ5
C2Gw/oxXFpbiEbu0nPTMBe0YpKxigOzPqO8hLGGWczx9aBE4xRcbnY5Q/TVcE39xyzL+2bNJhxx4
AZ8OR0V+WgdfUM2YVe6ZGSKlJ45h3LICWJt51PXA2skbqR1iEEj9qyLANkQo5CzIwomS640/wdui
3yZh8q1NQM1EkAnv42tNwKcSNQIbaJcv+UEvgmlln18iZzCgP0maS6Kva9ySLvhemSlaugFyq8Py
Vp6fKQuzfEyFgArPWNC0qmblkowpmXUBGLUc63TDn2k0s1HaIoVfMFSdJfupwiBr1dhKTEayz3LE
7PrfnPSbfZGD1c5KYkVS0oSF9gK2kX54hcWtO2EPcc1WV3OmD6mXXXi4+uSQpjIU1DEtBzW0qVyq
A6Q57ezKQ1Bbkv+OpZMBjXGySIXQ2JG8n9lf+I4VTWl9aWNHbic6RefVv7eHRK3r0NlW+SfSWFhF
qsybG5fddC9flGiXufdp94/QSpfEfzlU5FfWW/v54wdubJXFk44v0HaJ7Wrg7JG0zaFM151revv9
rvia24hrE00wB1mrdwqPILWZc53yYLxZuQHp5VIZlvytIhGQdYRLeGGwY6GsbVMXgRwAaQMQCK6c
tbmNsgjhY+nykcBYgKf0okW7c9iTeADNEh/r2FuSWT22mIV/fWHOm49QK756nj3J/rls+Qw6xf0P
T3q3SH8xOHMGp/cW5AjDlifSdOwnoKFvYOiijpePL4QfCDNfv5HIMb1elXk+lSyEASDPrkGpzJvj
f9AybCGm6hZmJW6wzs+5JkTyNGMlIMA/QLZiHI+46aaXHdOsEoMZgYY7TAUoOg/yCnqPyyHN2asG
9CUElxSPEvNAapjVhBMacojp4L3telMGpL5I5Z42QAVHDJMbSMODsyjwu3sRWUuSDxYtiTVY0qxM
S3jp8EN5m26bzMlr6p+fUr9Rvw79IN4IUnyhug25l3iyEFhbnzk6Ml1loVGMy2RSl3xh/qVt3Hp6
xBsSenDv1xFm30bImtlXLfyO6WIeiH4DTd0LubnVo5/w036YnfebcIqPGV4CXWbbV03qsXfSSkoy
t9fXK7wg8KUGTrqJ/6pdmEywnV1gEkb6GeOIDsx73cCUvWJFL4a42XopBBZstfuR6nuysnY35tRV
M0cDnGV0AULjpvCBdIDi3vzDToFO5lLoXK2M0fiwlLWcD+gPYSuA0tsDOYsr1BB2W4JP2RahiyHV
t+smGsASKccmHXM2IHJdLQbJtu1yuW27U0/PptNzauSdZ4fF04D/Hw5/rXmRCcuFBB8n+fFNRmnx
1gDk6FLzT+HV2VQ3rCTq4Q8PfKD7QH9PTQGTpMQR3byul/3Tppp/PabuzVGVsgFoTa0p2PqW6hwQ
88GuPMxN3u8L9TYE9ntCGeM36Ipa5YfCuhDo55hSRcgvJXOu6H+OAgWcU4bkohDiND5nYlCMjD6u
MJtfQoQ8o3YNg773Btrrh8i23bv/T9Os85/WL3xT16g5o+upJ9EXhaMh6MCy6RxfGNfhxVlMd6Bf
kDlUjyAEj7VuOFxsYGM1Cvl+I4c6SYl7+xawDpkIoIbSRAwzkpgSleFqTsLm4GkbgTw7Nb6wlH6n
O8Z3imtrHllPqYF5Pg06rmFw0rPYCdUG+5YAUGSTV9kcYhTsVEbdjt5o0tDrQIxLBuzXXGBan8Qv
zFP2CYAynecz1KLTRlNpZVHLO9XyHuOINGGqUUHhE0o/+CWi/k0bOzu1D5N9/YI6D4MXdbKtfI8I
I4O3nD2yTsJlJyo2wh9+c+iU6FDjPkSH8A5XEaP/ud7KCHhJYFiWBLtVYNQr+QCmxlrEAJozCLgS
V1Gm3mi195Ft+whLkBIJX+9oyfZuNGF6wLmjTB89dw211nANg49RzTCTL2QSOMGz6SUeVjvPnSuB
mk1yrTBnp8SDe7XoEH++1Po8nGpQIINvyOH+JIf3kIHpuqrQmolS3ySIM4v+nL8lWOVGPBYd5AUK
rvELo6SfduqrUAMSRbniLOourUw+SRk22nAuz1lLdFvyhj9ans6IdL9DJGIrKd1iX9gfFv8rklaF
H3GAnplDXVdBzvMj4IlC8FOV2uKCPDYF6dk12TL6bjOsBb4rdfP9qZFDBrdBCcx8a8iGyOnH5sgl
RtGhkk2qSEZz3w8T1kuGrKnM4qBhGDqjuMPmAS5wH1wG9NXWcClqoaVpo7SgwJ2k3d9t8K3Jci5T
m03AWKArF/aUUIeBnetclb6cA93XN7/ClaZus9QWt1ev0bpQ3BLIWc3Mjkjpnp2hegRkoxFlxg05
fC1tMAYNAsaDgSDJdqK+iF8snNVqhVPpWLK4InEPgHoiLVpaNup+AttzQ/Y6vj67kNXKA+AoE1Wk
Y242wKY5ZyJRcj+CMaWhF4xW3OjLSHR2jl1MMaAwOj8aReDUbTzc81WT6cUDeMQwQ6m+L/mG4U0U
dEi2b4JuFwrlE8UKcQvK++ktVXElczd03ZT1Bh/5/C+DdtE5Ud0PodYOK7ohHTCqiEnoBx/RBxtZ
nY35sUACucBcQnmQqtcSsk9G0CWrueF80yKkzq0iicD9fpIPrXrWLBYcw5FK9RoGywgAbuza9R08
RnoyneMLZVd9yS4Zoq3FmnTDIfyp30+taoZOe8t5fN+0qg2rWSorMIcsQyBALS34AeHvTDmCdE90
VmTl50AZFrhsvaUByQBFGs6Dvusl/ZOPKS6/bpUX3KLUwl8C11qmO77exE/XJjT8iOEp9sky6NaK
GsauAihqe8R7k6R8tcZ/GkFWpTMBgYL3oGvBZWfbTFscKIBKB3Nq3hPv/nDQwBwSVwEmWMJLkfnQ
WNmKDtvszxdw//ZXazow/QiYGOW3dulnHTjaQBSHV7Kly5WJQg3EZsrczlF5EbJPQQijJXHxNJo+
wPAHAnybwLjG/07QCqBO/FWK02UwC1cy7/vV7qYUK938ihbfX7mNHy0Gk/TSLTMTUuT31pWPeikS
Ghd7Nd7oxjtlX5xxRgeU7Rh03ilWFbFx+wQkxXnBxWJ7u781ivpkwyP9YNsGPdCEF5qYE3dzvBAT
mb02ddU8qvMlyZRSWWwpHTb3yN0b2J96dv3rKBJB8ANKfK/UBDo0lCM7Xr5TxNzQ06foQ46ZhYPI
5Zp58YH+0f6D9HVyCWxM35GZ6PKNv501dAU2y9z4VwAb9eTRy5WrH6L9yFonCWKRvx6wCYi0JrR7
kCYbDCGdYmjT6oXSXPdpgtMPxlYbk3NIfnlaqd8+Pp45iRXarIzSPEPFIDS9vOVg8LNFqUHUTXgi
AUZ6ZmId1nwiGLbw/7zV8P5t0h9PEohCx6lJTuwz5cNIXS2N9lc4CrCNv9O0tVxyf+FsIwNYnldF
PrUdqee0IDN1kmRJmnUf9YvIXbEjllg1ZnrWzDKOmc8BNJThqA4Qiu4jt9S01Y3c1O6siQ1L3EBH
zyzR7Tm57dpvP36x2B+pSnKmlC4fuTasEMa8qJpkZFovuuWlQNoeriV3wacmUJZdRRoy3aya5Nva
ivE3hMK/2DEmQ/VLvlJhi8Typ28QMfjiN1IW+FSJY80C4+LfD8OGdVZ/KxfS2gMnqzIRDE52nQsu
uogJ7BvmElC7QLBeYHGXihguh1k76Dkt7KnLMadT6LeXU+F4+9t/SXny2izb66Sfhnm8yb/cix6n
zPiNWwQNXA9EoxnkuV88t3+hQj/IWnxLxu79CcSungIeq5eUKW37cxgJC6s0oCex5HdS9ZQEh31p
Hlv7TDhsJ4wzkodOVjJPjsQJIDM6WweVw5JUyOvnoCZ1BrEoxWHBqjzUdQfrS+tmAbY7cOX+LI8O
5a2c0KArTqMLONbVdGrfRQxPShBa4KouUxeiFoW0GXtABQ+dGo3DZk1DxTCwcBi+6MNUCQS6T15J
g6kQKlvtjvs6wVe9PnRjqa3Tcr7Yfgs4fciB1PBehwRhJkXXS9alyTRuS8jt9k7pet+KJYdjSzdl
rCEJ5zs08QsaViwfrpHUzCsSn73fP1KJvJ9SwdGEgML5zNqojPtwMEYACvxKRp7v8opdAFj+t5tb
MBxM+GC3bQrwlpS3plE8Qm0zkaKR8ulCpCA3eY92IheVqmNhea1uXVd59rnP43GoyNxjaOWHBWXH
mJeP+/tjKW0yCnDV+W9UtaWo12e5hV5xPzIllGO6C4ZCFKnUamvyUuLwpGH9NFofDcRjUQ/s+yu4
KtOMD67oLW2Kw7pMaEHwgcwdeWnkO0DEA/Yu6VoYgofiz0lpI8alnRKNITiYhNLYTEIOSDHoM8+Z
uWGDG8vZE7V9eNJhGXe78MTQDI9CYBvaI8h7xhWnf4DtIgdC00SqCBRy96ocxvefzZRkZwF7xZN5
bqKesfDjP2KT6P79q5Z5O+1fYizzj2yFh+tFpbM9k03T/IKN4WtsS9YwKEcPcbJA1dXm8uE4MfL8
J62I6sYp7UW4PXxM1ujtzQ+2MRc5tBv2DZjjexEjwuB02Ud42uUViYJjnO4fQbezymVnJIOfmEov
/ayxaaoSK7PfuOuJusuSHJ/TmtiQMpzXqyJJbTelNLX8hBzO9M6Lh7xyNWcApPotvGCA0SlfBmLm
WTpEKCgCnatLm9pjf0Lmb1Pg8ikrh9QvD7qEEiwQ6NbsIT/5yRbz0cqPbC25sicPnxmLbCgXW0M5
SxssWa3kmT7MThg1f/OfTwk6nqjG7Hdh4cDd2zt+r1eMqBVWwuWB8vw8Vn9fhuc4IYRfs9NCg0P+
SqVCxGlrY3GSELcbuPOewZjUYyha9vFX8+tMxqkEnIQzXvN+PQqcienrmOASOtBFU1dRfCvnt2si
y4AuBFCSftnRtAKEJnpGGAs14VgGbnDhf/mrdKS8wJHsyixcUxwxPhMbeC8rhrfg6+nTWGi/Wc21
q2SBStz/+EK+1rrsdNlj/K5VSBv4L8xNFo6NOOQsIgIYmwwCjftCwiveyFwYSnkqAOS6+Sgl7Sjd
HiwIPnm4K/1rsxeXSYfpv0/67/1GN+HBDvQvo9BbROMeVl6+uRZwAcTPzqV4S/g5REyqVCsvKoaw
jobg0FwVm8yNSzGaDZhngZLg5C/PZ/kUrJp9UluXHh4ByFz7+tFZWc49ZWG2HtNBxf1LK1dXT8Lz
5fR1+LZNUD+d5YBd6HseJPVAkQmJ3AMAyPV78sUjup3Sn9b98V0AUNGzFbrsoPN+rEpLIMH3dN5a
cYITqTPg9DidY5zQClrcOOaa6sXtHm+iyaKPi8yxC7jOMsI1XAOwNZ4uK5OK02jVk65pk81g72tf
GVDedU5bJgLbdS1yLX3pOH9PgaohCM7fFJDX3Esu9eVfOkFDajnd+bW5mMrPd8YIQTMAzQ0Qv6Jd
PxozLhKOp9/rHqx8wLURujmoZ+8HksN1dVH1Hhq5VG8hP4fyRAsyZhCgWbQH5cPDYgIgzguWlIG7
0yW+C/9gw9zfVr6kyA8T2qoZckLYxB++HgtQOhyNjvMXi0i72t4wosz5q2q7+4OPLeRWu6ocSxNK
/oiVS+aYPrjSHHI7d852cwj/AbXQ8rGdYUoIY0jt5Fw1kdl11xAuh0qvF8c5yGX7ZDWquA7ThtwT
16pgC37p//ldoPJekdLxgIdrH/Xaz37CLuxzD4mAtCXAnS0DOnkIPi051xPUIWkL1e12Jkinjq2k
1oCuYWvNFTix3OFd1rFexmzBau1cUyEeUYMyYHs2JqW4YLRWh5qhL23P0K4rtMhWMkAPi4MkyOYv
NZWaDMxw0U96ftRnz3hIxwLHcZJxoQ/puALkDVqY6R/PnYz32SM/ey9CXpR9UXWBtcju3cfeL4cj
dRw+xDYff67O5ZRTMiv3mm6LX3wVcg9QWpiHcvjn8z5JTF41WKaagQS46KzbL6LF7y7iVFfl3zL5
Y1yQHw3aQJjPnUsKUVYh4FBY4a0Rw0OZKp9x6O2rDbnWJ8Jeeen4K8ltUOTWM+KxJbhDRfF0Bfwp
FfkcD7MwMiwIw7QbnTT2U54smO55YXLQ48Ja/XSdPGTjGoqNrcPqcCPRk2IZ9V2eh7plFdbW+/Vd
wVaGRBGl/T26UEjPwECWwqVAJZVRaB8XWkNfQMi2MQvNkoby3GtZ6rWPcncoVWxMZytZP8lBzHD/
HwQ4Htcv8A1wCz7sKB/Ad/ERvkuzTfKDlexrcHZFzhuPG7RnD8xF6DUMnKjuTyXvYytreDwyM6st
gG0EESsOITGTV5mfTAzqusyIa9rHDkUlCSoByW3fYElblbCjSyUNkeO60sFOpmGK6FcJEwZ7Q0Gc
mcjtNZoZIyMGlxtx+ybjCqK239pAWps6H2D/bZmKsblk8868pOM79mASgr7SKH52zpezj9aHu9gU
xuJ1jXZQCUuSicz0byuTiDqxyk5RVqHuTbIeJKWrnoumJSLTOU0zA074tqjbEQjiTSsExdVFgNAf
Okfr66viBZkRJpx1+OIn5d94kLBFfB8I0oiAEVC41NcjO0T5WLNQ877H/zNpGzLX4LnjAcOBsVuN
RV+P0XrXjS+pShN9GOWUKN8xTImafxXBh7qaaUvIfLcpzsyEstJw62EwCzHjPZa/gdGlmppx7TGd
jKyQ2E6l/g2Dpdc+TMyLJM/p8pjA+nytXhebKkYFYWutTmpaj5R+WaBmgXGIaKMHCLblRG+/7mTD
gPPdd++7djmcuXZJHysr307FkGtfCDeMDdM4rFckoeIypHyFtBPOgS92N3NKAwhIQrLeq+MK00OK
EYTloxYAPyCEJTBZoRqUBFwixu/y+5dxISvLG5FxqozJP15SIbLYj7MiJSI2vwmgg142IkQFxStf
ZACa9MGEE+Yr4CSJ21DJWqicVwbFK5nylW1cWTMpdbQX56fmxtsFT3JcaQKBvgj+hHsDLgFKZIoD
1/teKtXSXYGpdYkSK2RHt3jUdA2uqFP/4KphSA7e3uoP2/hFlYmpnNGXhZzKncACgtSln8C5upem
cImmIpbSaFVlvAt/4fV6ukx5RWMVQSTIEuxOqRA9QokBRy29CzYOM4bFbrSTmrstRt81tfa6nnB5
C0gEgulj/j9MUEqM9VNDR75qYS8bpo/WzQ6dz3jINhy5U9NPzIjFGyfXkPIYv5Gd6gBI/nk4a5jT
IpmciLyXSUXqoM4tpsxAtGNDjRbfBkwsL7zmESQ16K6BQ+U/zyu5nAqdyJCpesExmpuRlUn7KxQD
umrLModgBeQ1o8yITTinIaKrrAQ1afx1hGybK+iWjwmXWUHSvUyC58M+iU+uOU0hQOfZuSm5UXIt
8FMM2LlPLPgl6yZKUVBKYgJvO8gLCke15A3D95QBGwe2oujUY2kHHn7kG4bvSv2gOBXEMJandXh3
ZVpZ93KXoNprPOk1/ZCo1efwdlBrHYFL69JjW8m+4Z+rdAtKQwomNohhNA8dOaHSFApqXM7xj8i7
N9KrZw+To4Z7XYeLb8zNcDT3GMwfdwwwrJvNV7sQojLMg96xYv6ta4qXgxqSGqjAUL3cRgUpa0q+
/zhCteRPCyZK8iiazCYIcq7I69+jlSuB4q2ag0i5vSnoFc3MshFkEqL8KHvugjLJN5oRPDg+AiJ0
bo3H5VxWl9K06TukRb1fIttHf6SzIn53BI6LPWJOlWkGIhc49svKpHdttkOgPbTFXBTaDPWhXd1M
13oPlLs9LIlkWZYodp5I8mvgghomwYhxI6JZfQ15MJ80z6XckZ0y6nGqEKGiIFfD/14IfKYcxDnO
0wk93K+qtdCfElz3IhZ9sgAdu6iA6iDJ8usRNBQdXGXcmHvjgOTVGgBlXrqVXijhtdMACWTRd9+o
1nEe5kw60ZnUg0lKQpraw24O4liQoNETA7YmtMlPue1zPkucA3A1F88y7JpHcT9okmQb0S+NmXKR
4+sYWS8BoWvl9chB/pdXAeRZU1TigxHAv4GLl0PfOmmaQl5oMgsimkPuOHtCx1UBpoxGFfqthQJS
BtmAP9Qbcx5zrvf6NjfA3Irl+30ewWIQVtnu2E8vCsCKmM6qRsI9AheVqPNczZ1/sMc339Vs87fG
lIWPIekbk0c0264O9yzsV052vzPcgEetmk4Tf+PGZ2G+xPYwiq4BT5g7HCCQhBfEhiZd0tESabpa
Wh8jgbAqXqK7YWisVjXnMhUYa9lr5E0T2L8puuzPfIY1d+1Tg+zAqHmpkq7lpEZxdZr7YMedcxZr
fE5rCNBJmyKpaJyDvWIGBLWDbV3CbdTDP04b4h6lbl8Sl88WNyTFG0adGUBoDOFgr9wievfwM2Cp
z4VBEsXuI6Q6h3/wct+l+eizpfM2zJLxmno032C+PXppYS1qRcoWIgsPraZiG7m8JzlCMOIrzKDB
q/04E3Nvay1fFkUi0N0eECZ6Ouxno2ApSMJXTCAanIqdQIGQJ6hqdGBfj/8E2JWz0qmR/2ctVA9T
KVm1+xQ2BYauLxG+cvg+30vt4yMn25xyKTkbgnit5ybnvWmg1YjC3Juk83LNfiha74njwYlSQ2EV
sAkww6VQ5AXqlyGunfM1g39twP6ZCitirbNqW8v6r9n2c9PRO5e1Eo5n/erTxAXvZojPYMTuAcwI
FiRnWGFQHFcmlrFh5+svrAOEAH53sLSlvVoNUo4Pq3Tx8SMxNBWLS5ubT73suLAEfO/Hxkc13g3v
pPcmHX6/1ftuu4HPbiQsEMv6ll1T/3fXWkOnhN90IxFsI//GGg3X6r1FGA6AIBjS7Y1IKoilansi
Pt+xniIP85VanBue/2rZBsoAq/EaqdtHys02Ksco1ZaSIVHOMirYRXlxCv2nCvPDpWZlIB5EYsHW
v/Uh0XMIfz5/JgRBBnTav/nBQKIq85xoryJVHDRHEd/jPyQebCkVNfH+b2tCymfuJV4bvgro2HT8
U8Rnji6ct6Imk2I95TJD7bHvpb/csdPXkuJw84HvZmgQKceWAeQA/aHXNyBrhZYPzZISjSqKicDv
lGuwpEHX7D/lskx5hVamNhq4KqlaKuz2UKbQktjIJ/5yRJdy9563q1NQkefndAcZXkPzCkZSUV0B
eSWi6FSVZ8+vhjIWfdIUR9FH4LcIoXMJhULfoBHsp2EUT5TGfiHOESE7wPUSP3qXuCQisrz+b/P6
qVvFIC32Nmjb0iqGJNmhw+2sdO9Eew9K59n93HWW2x5pxF7fNLKN7CDDNSsWbP6J8djk9Pn6IJKZ
Gn6O5f5OHIAK7mXM3PA0K6NszPiKkkLPRA1CsS4QH4A4ye21RB76m0KYwlcp+AoM2DfATPSGmBfr
7FGuqs8j5/qgXxzLpBYQalGjY1TWJyjlxa9m+iSS+zFg8pbd6hV+sXfT70bcHWt0dB+wMiA1cIPc
6kgnFmfCRcsF3ykfsHTqee5/hZSx5fs15VsEvotOdt6OBlvre1qbMIPW6JhKv86bmiVPuLxf3ESV
TIidTHhtN6nb8LJxqUqfCuAKsfUlK8hZa9IW4Vt+nhc8WR4My6mK+y6OBIPpGkfyYz8jeScptLib
tuTLgpeqauYqisPrZELY1PnQmK7xcQImw/kGi2bucXVXUe4LW4/iQMDnfmNFqsrFf5pnJHfBzS/j
ypqysB5QVvH18Wh6Gor8ou1W7ggrEWKnViIYxooM1IShFG8utMGsKFZ4j9316kGDxcAaI4dAEtH3
p9n1YqolYc+Hii7EG/YXO17Smvmdgc4tTcfzkgQTDfZr2WxgiTfZKFXJ41pY0ZxIFW/ZZ+c3GwSs
Qde4S+ODtrUDDCtVjn9FiH95tkUfRXGSdIZ8Ns/WxlycRxkyD5ZjI8JFqjEdUFwhuxdDLdl5EM2d
Az0YSy3CYm/n+jVBFsXtGDavshFxkTx6GhhCvQagXR8Bn9XdQv2tahEC9dAmL6RybXMnoGqp73ii
zOK95gQy2KO3t0RsKX9nYcsmuZmgxdVcBJgCoW4vf55U2XgdvzOPbUarPnVetjzkvKL73NYaYvD9
59ru+yCmXFDT710GH1YmeyPaEKu2rt3g1V75kQDgrZk4empor6L6zIyQgIbcjK70ynkTBuJqz0MP
r2A61XSH1MxAsiPNqDPKEhuOeF7cmO132PVuebX8LZwxg3sEdcGs57y+FgFp2/+12D6JDZkZtgFF
RJOVRhLqwl9aHPq2SfSkeT633FlXZ5AuBctpis9r2xXatYRJhTeYKVQIJAOS35UncVKbmQUsO5dK
15kI7zkLirPXLTvVGCvWwXJmVOqSWrRbQaMr44tfsc3AoRRav1TyQFKBO4p2QwxLX5eg0MMaqwMv
dz1ydLP1XrHPGzdNF/OtaIxmlR0VUSfVcUxVjLSiSuGlCR5n901ut3gDgg5YBAv1t+KStOe/UIDg
CSzwNSStu4gAnKpAGMVyA8wPQMjxZ2WuTSdS/ALJT0tM9/PbJoQyTxB7muD3Y3izMW+YFdIxYsxI
xdHmZdXcXG1P3zIQNiBsAFjX3aVThwrp9vmNn34v7P6C1KiSgkI8tquA5YoCilg0VnsUYt8B9xIt
klmzo2/KvjNR+Qunu1HITwvinukbz6Ix8xjlqWCLTrazHwrxorx7B+24JhJVn+ZIJnKqCzYjsEDh
1+zuGNXM0pSBogIMu2e+SiTjKbQJyLjJrq9C07TQsaHOzddvXFkhgRxEm8SRJVhVOjlDKkMJq0Rf
vVE837+lDsumFeWUioM5gWo0WJyhtD+x6sbDEiFOSZF6+VzRHUbatFN73haDrLqBiuFFcgFArMsX
H4HBd5Z+XC42OWcHax43pJX8x2es0D3yiOjEskyysLXyzc/JSanDezTUVzJYfP6PgZXdeeTuHR6W
xn6ghg8UiRI3ruksm//gnQf4x9xgf0+HVqqrRmQuvARFeliqQRXPjn0IBaXwGCTRvjVbgCKQUF5W
xdWOAgtteFfnrzEBvg+a7cwjTlTs0MYBdMB+SRPMqj1WG/SgJ3TSNpUViYm7+oYgpJNZTd6Bfoer
L6+B7lbNPLpXX2awUhPgLQ6eJi253Jhu2qJnGmzV4xZATue9oDzmGl16vIiwO/2E1rlAGsQbq6e9
vN4oldHY7yH2Ixkv8DlZEsUcuMbbLfas7i+UkJqZKJmdQDBs+A3HgtWrw6cSuq8VWpTkVnLSrZMO
bdFCY6qob5VbiGFABouuWDiGJfBCSg4ItQLoZNnVcL2B0r2AJsmoOSd5yPcUETFNZnETifQ3CF7x
zOhlCcUn+2rFpZujyyGKFCgRHMhFLtqzy9LMfJtT1jh1mSePBH3tGD1ETtFuQH9bLC3EkPMAQ5P9
q+3bN2PEjbQAOxq+EQ9R9dz8pK6ijcHXxFvj8qhvzNMbxVP4qCPgRQ1SDuNJfCL9fjyBR9yNuleX
9z+4HTG0qI+N+0T40KdlKpddnCHyCRqcfspe12rIjSt8GpGkIa8xI4qaKsnqemECGdQpw3vE4U3o
/bB3pcdu2sRVlhK+52H4D0dnAc7kXl+tPTeUeEZ6/6FdPTtSJIiRpnLFsBtNz4NKNDNZrR30H6OH
VQZUbjN2bE5maN+3Z9lnjCLAVsAHSBeJ0fxCjcve7B8Q2uA5975nRKLZjDBNU901n9HY9eLScC5j
0iE0u/c3qRNhfiTJq64rpa2KD2tqL45kyzZR1c3f3ONWl681iMfgdcW+X4xH3AZ4u+Z78vpaWZnI
LZPE93a1z0vYUuOJhDWEMUbkMShx+gVJ0SW2bY9WBVazVRWln5G7+JA3eaCTjHaF50WWxgCqeoH1
16UTd0Naz8fQk1ymZMmB7nQXaWqeOoK/rx2R7GvifDbWJqmcll3rfULdCxlSHNCY7WM+mYZnPinY
moNzEe/jz64+VnubhrkrQ4vSXNj7HQGuO4r00kFKgOzIqjxInsAV6xvcuWiTpuG5yLbfJ8DkUbTU
gk6HKIAvsPyEMWWwjoApdZ9bwMRfUzUDkvCMuz1xMRrCLDYMg0122a2M1qYKiqJaukW7gtHpqysh
FOWM6mxHDrdZF0hbWqUKe4xt2gWcGRT4+RPuZk5HGZ02Cb0CbG/zYg+Z2HOqX2FTLY1exfGCpZaz
vfkZ/pflfabufadk6T8GGBMk73c0Nzk9FgXjVtO+61hyLV0eyPGdBH2JsUCw7GSWvnTzj+NZ5cVo
tg+L9xvtX7Z77U9hQJef/v2yuqxl0TRutHaDNzZCnQc+a+BOM1ESxd3NFBRSqdEzJTw+KUPdqX/w
l0rI+qvwHmPp6qO/61UpT1mLK4C8bmw2u7yG5hTnyGlxTA75JpcrXn6emjl8aWhe0WE640N41J/Q
bCvLTihp5jU3KSW6aOXoGolcSztewCbhzM6Dhvg3VcA1eDQCztah0ktTvMamibzXwXoBcy8z++US
gBwH2skwcgVe2dk9CJZlkxd2C1hcc9sij53aM0Yz0ElaZNkHKq0dt4K6HfOviAS7T8LX87xBWN1t
Qzv11/BYBXxNStsE11ccSrFRUaitw7qscOqOydRz86MiUqSgkxyjZ9eHLXhj51ld6UNrIF51+R/w
/acmLQIzBJ3NWplhqwYxJEZXCfHQa+HRx83opZ6xJrNDZVvWPorBszivEcvcqb1eq1/lJ2aKstbN
XXV6XUz0jfoydxHpVpnFpPXBzSflNPM/bGNbVmQJiw+lQmyuHt3PVNg5Y6Rw+DXPI40SNqxoLug8
njET5glNOY9U3WTc9FLRFTQouI81ShC1KLT/brad632NfW9/g1scc2V/FFQpxoczFz5ll9hTuIVp
Hr7y4pHtGj/IlPxwD20rxm6pXeoIywuv+RQPpuIh8fJDyF/tofczrl9y6Nc6qgMSYsTB/rnVhKP+
emW8aq23b6V6qdglCCGFqHN5I+Hf5TMP1LoTYH79bA2MBlJprblN6DwxDygMDLfBdve0jw5V/9Ml
O9uhksaFFSfhEW/rskKkunZ1q078UEO4+YzLFNDQtW/dX+hDiF5tzI5kP8t4iUtJByAS4bHfGl1K
Xq6doWtP64A2hPt+JMSMfrKTM1JiZ7OwIeuFoHdlkRSdtSF6+5v+mXDHeIlMFniVXk//ePA0EP1G
4A8aGw5qdsxOQpVyL8V22uwUb6y7CG2aqLp4w77d3B0vkoyCPStxlRFgyp5b6u4CTXIW8lFy85wk
3WzoSbNCKZd3SRuJMPfNssSyo0v+tKWuAGVBGdFYf5GlLh9X8kB6x+9gQAlnGI9XBg3EN5FwpWsZ
E3bZodnn+Kbh1mZ83/6F/ZuHq+BYdZSuxeJR/97lUoozI6AFiPwru9d3HfU5mz4ucM7tKqYHgHi6
bQuo9m4k0dx3Miar95GpG7rFxvnX7LarY1dgJ8NVw4Ld320CozYysA/Z7MEvjYJB1UeXkADl50b2
IBb4NuCs5mynBJrpm1N4Ftox6CI64soWluViVsCzkfFifbRsELT8cMsLA2pFKdUZFKb2l23RMw4i
HSfS89dYfPuavRRynL86aWBY1rMWRzf9IEvO+WZ3MStvPP7eOd3qBuIgHYccxTNzu6+iLdOXb4L2
i1jph0chIqmhHTuzQYiN4BR3krymetDcljgIt2bvgtsXt+jY1AJZ2QvKpsJmyHm6l9bkoD6DKF0Y
dgnEgw7LWCT7jn3YMeIyayI+DuTTd30mQSg2MyzVof+MSwgpSgDFPV28W0AJbFLRJV5DJs/CdzD2
SZRkWxCXH98cCF2YNlsT8C6oZjHVRplAv5OY/ek2xw0n+CLp4tPD8JB+yTc92asEw7fEuDrvC2JE
rA1C6H9701Rml2qiFMPQpM0NJG4lALv7pdtD4tqm++4D5qRTiPkKqjSjGrG1L728DA1lrZgNLZpA
JEZNnQkVJNcaCSno6Fy8T+LhOvTiE34L3gVq+jRM7BuufwPuRA6XKdE2W4q0wOcJR6l2qgBMIvnR
U7GK5ovbhy0gaT+aOLFBBhjoEoyfZkcaLvII6UWkHixJmOmRNXhfW/ddRLGhRbcx5yd3qySg/yHt
4LjAqBNzrjRgou7chibEA3pYmi8Kx0CxPlRg1H8G33bo61ZASwzR9SyojWg/5dzSvE5zJ2HKqyGs
6/j6ykbmyFr5zT8xGmzFoi/39xIFEUT/fNWZn2DxDb5JJ20ktCsJ6k356wfFPDPd6EdC1KhABaYa
kM7GF78jwjJlrRUtQciZSpThN9AsV82FFMG4e4JAZwvMvkLeBUq9nQPA+VDwfYTyz8EIWXcbRY0v
DK7mdzbc/K9BrvDzG15gtIhVJ+ORfmPRwPqIxnZ+iNFnZaPD7Bml71KTPL2cHo3LCOHiEw8S8KYR
NUKufp6MqC5EwuFvzfPYO5jN1ingrurRvoOPDRnvds8c/zN9q68ieQwu4ZxTjTnfaBGWzUw0Yjim
tbG/899FJou+6XDmBG87Ar3x8o3BLQJ63EweneRwToSA+aKHCNceDvBXWn4V8Xav4U+hBBvs0KJR
vNns4AdZxZvfuomVJ24f8zyAxW0N7ynz+BsZPYicaCM8vGhdozyk0PeR1oPBuCGKT4PnFTH4Zcpb
OauTBXFlO46ZC67+J0xmn2yJ1XEqj7QZjUCERA+Dk9WJBNMzGh+ORer61V7ujpVQG4EzDvH1aece
/ZEYibiWQ6+FrNinrlWkVymBlQO7aWzb7ORB2KolDRjPdfrpQ8P/TbiwSu/H5ufSJWuT4drenYJ3
2TqayhScOxQloY78fGKkCDjelI+ccdKB/yMvfRaOISvAgnS5WSW65M7hzaiCi0oqrjQ6CSYwfzde
dcT8dNv4Z5DT6B3+riBZJkuiLS2VeHql/IAcj96niU55abeNwea0zX2tDR79k8blVS7U3B2N2NZ3
J0wLg5nLUspqjkyS/bTrTM1KBKQuhZwOLzmusezTjxPHqfPRi1XZLgShRV5dh/WGW/jKLfjf4hdm
aEHTGBPV1dcI8G4AkTlcvbJ/EFcHewuA0w/qRA7ALfZkH1XBAKmqrlTqvZ2i6owbMdydME4KrGTG
hv2um5Kjc2GZYaIXAWnyEi1pSbx/G6qRx9Mec+7s16yHCxoSAL3E0IMQ7o/Vk+QKyLVwg2WS8yij
3OQRtntk8iCoaRqKj09td5+b4IvgcAgAJvRTUVSKcEEcqNZXOfwewIx5JrDFkr5sutVvaPbdK6XU
W4IcO2HCLHq5Jockpo5K/BH2itZ0sjkLunS8A/4X/vrL8CNyGRa0p2Xp4K3/HwvCYkO/GIvLb3pu
uqtaGGZgmgykGmikzqQTt2UWX/mYWzOgzxDWOb/UdMKUB718nrAItN2SNKNt6LZM8OOEurqbRwIP
UNzvga7wxz4DQEi5avC1Oqx9/9voIaFwC8u5Ge/2IlCKz+oUFqxgoXKY5LpEp0jFSp1uUWLWr2TV
dbCNsYvnKuXJh8TWhx9ZbBQsx+6bOA2ch4412ZA59JYw5BxxkZT/KnB3fikEz2zYMJKJkX1LzZAv
kUIlOmO+RdN1/M2ChIUKa1fae+/gn5Pyv/eMvBJNw+ZgUqAg9O+Nn2i2rIjUyPm/qneSs0dxWeP2
+/9EogW+6WQGU3Szw0MWi3iOoENPiwxC5HQM5TQ8aERix41lxEy19jn70sGcTfv+6LqOEHXVbpRo
eoP32Emrc2UAV9f1Le1W3Vg0FLPkwRCMBtLTQWT13tt8FdvKP3xK1rjDVWOpeGYPts0rScZQtMyU
GBwXp2SPLH4SVY+VSSRsJybq0BQ6eC/oTSaMNPlFx+enPpV2thiQjxu48/u74we0IFi20AD6HrUW
vB2FJLE+FmrrfB88I4kr90muPTFVIYFA1sv9ymzxc7aEYUetLYLVZiQayrNsITUwqENRccf9Pyz3
SIwvZBdesMhscVTSmdVzMmUQaie+lWoLubBUDyNtcfs2dr+yJjSrsvQcD1VCaAO8KhUhYziCsFaW
kHFtU3v9Mhv0mWdUSYWFF+LSPqNMPRsGDUORlXXTYa48DJel0F7x3dnUssoPLTWcu5Jba2t9j2iV
+T+dFLg7t9oOIk9tiljU1hTVIW4QIhierC8XGa/oJfgQIyjF3FiBJ25jgv+RSqrDflnRz41IAyBO
akELOoiYmzrYMkeXmvNTyPmcJn5AWj2wZyJAm/x7BxbWltcgO6BGwNzJBG282xpbkfJEIgbSHrsp
w7CTZrioCuNa/5XKTt4Qbtm+IDWeo0BLsrHY2e7s17E7KBMVlLEufncsKD0tn3NMnmrVDiNTGQLV
0eoN2ql5G6zmSXoD95Z43hgD8isJvVnAFaPJptcNNnVakjHcgAwm2KZTt4BgZ5xHblMKEL3AiMgt
RY4pqeUhk0OyK0hZyh3D5AhgtxxqMSmu5kDhKzQz2b25JqJUJaUcLOHNDUTjaiASXYAcvq0WlGWW
lVddGvyAk0BEDZlvNGUKunraFtjEgzYjkTYUulB9hPgY+tCfIrP4Oedz/xkF7nBN3Ge9LdU0s36K
QRs3ZoIcYC0HdcWHPGY9BM1qnCtKddwQzQGMqlWuHLKU/F826IsgW5uBGNfCjYjUw6uiEKv6M54w
oOAV0LYfJYaRo0mJgKBAEQVZw9gjhKxgf9QGMfaCG22JlSGUdgx8yxVkjC/7r/f+8iK/icIlmze7
UK9/86qu4Fx9xB4dsqQ/ClXOW3lzDoVzrDrBmD0LGP/tKWvFn4/eqVKrUTnAfRr96SfYHcWkhXT2
HsoVF4yRH4C4re3gCvBMwgTnbtzc5W0zBs51FLp849O7vT97Mqvv6/20b79gHHNRyrGLHK4FaFyi
PO47zHFTAdsONvbDmE6bZhHHOAFSv3bN5Rq4UthT/WTVdP6+WN24pLUuSIZVmadUdFUk5FoG7iCS
2vfPpLJ1xeAFKPD5Y28gBjQC9Ir1PrTlYr3hnQQKUbraHE1QYNAwd+1QNXM97Y+zlZW6DEabud98
4m60vwvVSg/Myf5GwMd9x0VmAf16HUEv60AnVwemT0afMl4MNtSO9b9XVfzRbDiJTAC/L92o+iBZ
MZ+YbFilyx1nAqabZWsdhJfFR1xdA0QlUmfQedKUMIPe70wSugJOrZ9l2vmw91cXSyqG0ZxWP1Ry
daWm31rIU/gUjF8veX9SdjXAKGiJ3WKiKs5Bf+zNuixBiDdX1UZ+fP/fP1GwEZ/yrzwFi9rxcF8Z
gP7lGX29hsd3fr3MC4v6v8SR5cwvRe//WyEMoAUJipyczJf4ImlZio9cmWkH07Utapa2kVwBRz0w
JFkX9nUhy4VcYqH3qUT5iF0ySTup5rVRIGznZDdo7Xr4PE1in+cI62ou3K0LRK+QHl6/qPbPRsHG
zWY8paKxqjausILyl4alPSGERByAYf4cvu7QAYqDhACfdNXM9Wbn9kI6h3qjjSnWR9Vsj5EtBja8
oNwv7wj7GSNkhxzL281tFOkCDaMcGAq/K4tam/G8ZGdqmEB4aGz3jfYsehD0GAjNKL7odoQcx1+y
w+dM9qW/8OZdVmV/pPitpiIw4qanefSzndksYeDME4CRwnOMj0Z50jEC2MV3UPT5tBoj9+cI5kQq
RPUjQiCmu8gS87P9qVIXIrvxVgyWHlH+8TRw3IZRVg+fp1moQSf+j9WWMVkWSWq+b+GSO9iPKl1X
D1NJ/adB+RSW10+VTK9PkFEKgxppMaosT2XTX+d0ToLQ1zq/xwIWS7S7tVMoGG5SGI5I2OaXoetp
w+mB6FHRwI42aQ1jGALwV7OIN7fnbZGYSLfC3ksCWDs/tLbV432eLE2RXaB61AgawlxroRfV//Hh
1TRNKU587UnmuvBM3u5GeWDUsTTWdDzeExYq4oaRo6+TvY1VL84uOm5BF2kVvTKcL7As92+8As8w
63fOGqL6TVJGUEcjACxnx3NP94ggB6JBBigHksDYqgHl1wXMhOntjL1rfROVzvBqxv/7Fn23qgry
UvmiR1gRCsl0xRvVS+8fZi3hsa38I3xy1igkP27+UFvA0dF4kISfgkz1PLJaQ0kFz4GBXfWSMjJH
8R+MfsZK/WFLpF4V01WJ5dePS5zJLEiCyfZiNNNIub6pZJu16S6hFPcoesG3PetDKB+G0kzC3Vl1
ChC/vAJ2e5UQtso+Ee+5dfp/oxIepIKDyBO1GeNOZl/Xm0u6YpHoqiooZ0NiE3NDHUF0S+J2StnC
RKNRaMvHs7AfMVrgeX1vLbPbIFanuKNlPVjHBH8shX23WMPp9ctumzINXDp2ijkGn0/gdGbyykJX
5w2G17+ooYDr45YTM9hY7lmrp+IM2WfWvW9EKZ07vQB35uSczvMtqcO1mdPvr9OAQhm/85qdIgxD
alKohzJ4U+EcjbbHh34xxLLJbiOEMkYo0tYG/AwpzOpc3QC+lm5cAMqNjlnhSfrCIMy8Hx8mduLX
WQkriJj0Slu3raHmskgZ7RPspX+uuJuU+SGXZeJP1ZeXrBHjp9/CAY++6danWuP92iD1+/opsQM1
YfAHRvwwI+i/mAc9CmNIiX7I3VBuhOMUST097r4pGH/K85vo4VE5aKaAaVKeAUiqE2C3HwgRYFsU
wWp9v8vPAhpVyhqkGgUxXP/t6kNaumLJtMAs2Bz2UXozZVfmVTSabCfVZTWE9IT52s1ME/jNVVnD
HhuzTYOBqVPrHtaN3rgGqOF+KQCaeIO6tTiZHf9qKWxZlnCKlyPkSPKCl8G5hYNa3KOwDfyINhxF
qvSSU+HqflSi4WDEWREbO1y/RRKWOwt4S5ILEx+PNmUsUj2O9AAjWznboLgKrGHsJaVQWVufbuj8
epwtheLvHgnsfRT7FsCxziHTqpHgMuH8tQiPLmROGZlsF/S3lVJnffkORvHr+/zLhPiHRm+1BZie
ZtMIW+P53jP+9/+31EiNWfumRXY6zxC+QTBnYx3/VaGexZAG64a9d4FEb3jCHmzmDeS4mKyKQ7WN
gr26CcFxalwlvYHs2Nh5ZdleYR4AmQ7YYNdItP9+vYj3URdJGLhoAWrpezWzst/Yko5SlicI2eh+
PlqqhFIb7VHvspzf/3mENgtI3KMxIC1e7LrwdNOznWnWYbgE9gG9yhh9zsRPUFdJRMUTFpdxT1Cn
0KpEOjRB+nsh/s2r9CV2rYOGY7Hc3JPYmAWaT4SAVOpOKZqHWleUaMrZGtAk9yd5V5oSa3e3sdp9
YD6SqE6DSxceNip52pgZYubQUnhKx+JGyvX4p8fVy2rjavPjLEa8N0432DLtPqwXtVuzpGEk3ptA
/n2s/ikF2ArBkSYzlxFSsF8Fnolzs9WHun8aAa0Bwc2ngwKOV7NZxNkIoftspTU/tCakKoBw6H6v
TA85+kzphm3qR8T0kQgx43YKn/uRjM083RUw2KrGkVec3cTCLVEflnhp0biLRFJCf2dgsPMUvRZ7
Hoxex9TswSWIEnFUm0q3bbkdog8DsiZiCydkZM6tBRGijFq6ZKqge/p1wz/qpQoQyyQBjC+mu4+G
+ZG0y5CKnZwQfEOvRAfTIS4zT1GhpyWz19J/j937JGpzEz4e57SyZlrtUCX86QX0Y2F3Jhryeo9D
7KNx6oO/cjA0yRErrBLfEWSMaTAc1GhYx1xdPUQhFY/tG/BC8vFG2e4iaF84aV7WtTA/a1XQQu6j
OWMYtD4B+5r16iT0MVPMUF6CMdQlQoz9aHRT6l2JE2iM28msWFpmMF3Ae0meORR/XCs/vMRBqpgM
cEQpB3tGIhqdFQfik2I4UeakZiMvCcx6rDXgwcwAvsh4nIO7w2cmbwZ5WzwuWPzZDUFI+On6PLWR
50VEcMm9n33z2OgppUq8oFBGk/h0z/HULSiWRSy8LVm9Gxe/Dm9kRU6DMxbm308g3RuNpNI66+Ck
VMYou5zt0mMFilIiX7rg8zuKC5ODunTIEan6DglK5FXp2T+JO+BA/Sddi8tSja5vrv30RI2Whad5
qEWze/QSm4CUeEaMCjtjy0pH5bT/SkBN/XD14JlzYJdkCibyhYts+2b6kbBvoeoJ3YkkDoN5p/Qm
DbAndk1iNr/nFN/Orb/6E6mMBxHYusL0tEQZ176COd8vGKnbeZO/35uK9SB9jp/TBuvPTspj7lfD
7mcIVl8ANWFXtqLanNov3MQY6CxppJteg1EhTgcZ2qHSjsJP/vLTqs9ynY64LJY4mtFU78attK2/
At6ve+VrEKf9elh0mKG52acsi1+Z9MLsyc0Eu1GAwML/B18/TvlUoVIOqFjODaxEDwF+Hx+oOWQ+
g2R0gP2OFocJ8fRaOGPpI/nah3e53cjpTI/W79MZXcTeaVEL4u9s+kaAzeg5Ee2vsRo6BfJALtpl
Y3wnxFwbLLcQIhPvRbIgM3Pr1IbGD3EHYRtxcDAJaZok+f5Kkw+iUgZqNo4Ok4jOQaJvqXeJTFxZ
0MOCqqafSAFsT/Ok6D5yVS5YcfIKAYAA5gTAV/LdOdg960dBXwe2xT9uC/n5ojF9IycbBUJJf8dc
wAIFjrFmzcPhjVw8yjSsGT9NU8av7NJU7rkAUnSyaWxsKkbtSRT/DFcHgz62FBqz7PPhfDSOe54z
iJlqUb32ONJNTMW+BNak+pTQq5QCvTakeea5hQ554M66oCxWa2yhSd94jZBUCacZ7CCWIiGinWJ7
3JIDLYqbydapX50RVXHK+qJaKg8HBXgwtGpdh2TnbSCxVPXoabJqPZHPrk3ewCrKNjWIP3HQYOvg
rtl1oSGMb7qR9OrLIL6y7nINc1dVW7SxBgSbmhBfzZAXdMAI8DV2t6ppqATfWSKUZVOMAv7Kzv/8
7ZH9ymEK9VP2N3hsVY/fMLt6ESCvmsxBJobH/oJ6Vrtf/D9tl2EsBRIsJ2A7fXEAWpBMyedxyvZY
q5kLGL0Q59e0oIEekBas2m07752W0jBU0rAy++1Og1XE1q01lrumUr6aeK/0WFimqZrfiBx3FYQk
9B/CLCFjnAbTsAeKiVIhSNENdyT41xXsrDN7On1vEiTuxLd+I0JVTDTEUofhfpNX6qwE44es22ZF
SmDCoFPu0XCw3msrLLCYeGfJ4FTUL9kibhgFUgNz80pIv7QofoYe7KUA1uMlwP71C70M8ChFFQRc
p4pFnO19fHo5brr7PeArBsJs8JUsu25OxJ1rXlPB3nmMIoB1YXJZMXNeNliScJv/ZCTrw0Rkq4/0
3r4eomcR8SLso6/PAnYhqSX/fUOxxTaw7R/9eYvHSd1SvU+aSEXSJaB6ULHLqQPqEVxjFYD6lc+9
qESoVRVcAzgQvdc03pVAa9YGiOPhabDV0MqaoVDZIR0EJZ0uPFsM40NKdnQRMZSiHifPvhnYSrPg
NYrA29basnMoK7cLNHjQVE14hXrEfRyHz9wxSPTnmNu4OwCoYPGTtK5FUJNj7f7TPpt8t8NVsqrM
NA7Ho5NFbmiCKfl+X4I18dqJGPjLCnbe5k07q6wPEiQ9yg/QVhg6uV1fEn1mx0uUmLLws2Jljg/8
wqm1DDfPX2bSOddSDJJthxkyyZAhfDPW5ZWo0IrnhVY5WrUmAHUwn+JBxG1h+od+vQ/YHZiEzjR/
izTNfrKx3a1YW9J2Zha+MYouy3so2cII5IGFxa+3SXtLtMmJvsfWVib2cS3mOv/xMLgrnN+DyiH2
tFV2DiVCb0lFiQvd1y+kb/5QNATkAXKwyH0tJueAfvOOuwlQQ8YBBQroLswblDn3rqJFZw5c3qIP
oUZ8XTUH9ISWroYsPzAjrNxBJSWDGd10PPQi3TqESWtKuAJApuQHSyvPUIntLCIG8jehFyzg2YjT
Ezd8KvtqrQOAFgaZXpcYC6eN3ll81dACKe/JSruFBXgNsyA3yaJaNt6yy0cpRXCuBIMynuBEFdOM
LRbohwuoC2Hrl+241dgy+RopgvvL+ZdM0I662L/ovX0N99qt5T6Hv+ShCYegfRIO43YMPjojqmPl
w6eRyIdQb6Kqb3w/2GYW8cScTDEAgpWE8TKgVPBartviiPvAqsyuUmPx6DGLb+Jnf5XrUtLIU6FP
OmUcP7yi1L3jIoF8xu0bPMc/Xoijju9jgW8C+CeoPxxhlvqjA9BaCsWGKtbI7SNjjwPlQcQdrQ4O
NPAmtU5a18kKiCIlCSlXpwlhLTsE4XXlhK5mSD2KmJ583mlyhx8AQOnpAXhX/t+BzBiDaO3PVhxW
hzWzxuxpGdpnNEAa7vNtzeRcGPwA+VVPkomSF6bvNCNSPt0Pn7AXsbmXAJtXRi28Fau+2TtfKLe5
0fnIffKKWSCgTPGqXSGasnJ7U88N09qqOzeaHZAYRXcbUzIx3YarFKYDcxe7WJcQYGS7z7smzgmT
51uaaQDDQmigpZgTKckW4+O0ZKfvsI5UJkhoRL/JSy5sr7DYGq8Nz/bRasEe8h4G0E0op8jnfNmN
3uekcjzwSyK/S4FlepVSRYmGeiy4PkHFXHKcMFa5FtcUbqDI4/4sjxsy7jxcyPSfwGmxAK+AW1VI
WNOVp58ccmcd1fAqGzcAfWNGvWmDoO8vRF2ac1P18cCtSHf8LdPnHBANKLJASVva2Mp4gJbig04q
S999LS5IiMvAiwettEpUTgjYLWDJQ17EyF5rwe2f0hVFDgamd5hA6fm0XgU8iQsbIQydq2Zend9u
HVVVrIi8cHSSe1o05XhYeufpTxlQsSSwlIHpI1WhBXKMOVYKlxcU62GLJ7nZiOry+yuI1iu16/z2
fU0OoyNclcdOf+J7rRnRRm0DLCVYZIWD8wX47VGUqrBFSd4DHlMBBjMlB7AE6U5JFud4NNzsIMje
FNe4WmfOzKhcQkqGQhlCdVaXrsZY5I7Kj0dJEMYya6iOrxjK3cJ/FRPNgnZEh4ttPs6HYy7EPAuS
HfMEWXVT94o5tuH8V25EXNZnKLXZh1e5gyP7aGY4YvZtJEAlphZVzWGBA/qdwIFuIBbEBIxrOnYm
qqbH9iWr+u1NdXDbQAVD1MsiCpHhTONLvLHqmcMMbmO3VyVEKvsMBUwi4XdW4s6086c9PvP2AIJj
ZpbD+OaujYypgRWSLL1aKARGDppSvu+t8BXOuFCsisd2V2HN5HtEqt4CC+S7WxHbXNyfs2+nMsPY
SjCJNFZ3utjLUpse2YrbaOEEMrjki6dBDs8NcX1COCsmCbZ20A1giEm3as7SkChY9shCNKwvrQN9
944bniyuJQxqGZKKIxCKYrsJhsij5kgmwe/XQZZK4mHTIXt4EY8B93Rh1NBPiOHok5tUZyIYnqhe
aQRtL4t/6jeucELkOGQu+a8F0lLosOB1yvtLNG51RQG6wOzoEfm7u/GGLeiNIGasGC+HBzQ/Cx0J
Rwisl3c666HoXMk1lzqCYXwdst4sZbjXcsFT+yUo2CV6bo5bvTXOHYfoPlQLLwSf2WQSfWjtLw11
o2QwMieMetdHNofCnMr5GKZ24qmU7c2MRMa/K4dKl42ivEBeZyLmDTr0kipq9/retTfsLbUnN3ki
fiKxcWAq84s+PusHrryijzdNFx83gUfbUvoQsNDnjOJX/0ZYkuVfTRuzRLBsCu7IbG8mJXF3nOjC
yoX8tg8IK511Q43BwNda9EHwDl05UvAKasEt63wWyb8Fg+rtjGjDaE+Uc3M1++JCy5Pqcoyw2BAA
6NYYXfAQmYO+3CapBzdjbLS+nWBV9EBTzkNYmLKubgnaPo4I2siAM4XLNpZt5N819JNpwPe/RStC
AZpvyjJlrBfAB0G+u3hGS1S3UlQKorYxHSi41u9FJCc0b80K/dnfYVQz0E694k4TBP8z949sdMTY
nzt2aSNOmqHt6qT8hlFHrtKgQkq8AHEyoNTxEcb1GEMXBm1K25QX9gts4Hz1kibr2bcSBHdMmsxZ
AhEmpHoIloisdMHrumqZTnUt0kQnOf+xR9x1qbDHAVlMXGy0zJkO0AvgeM/jGn13N5Qs6mq7UA87
NSotSHFL/n1LD3iWA4QZ7CwH4dhuEo7S6VO0AbxgDlcTItoOK5Y5BQWRqptY9m5jbe69RP4DBGAj
qb/qiyOguHm938UEcJkqyzGjZODbQDxNe+kAfomEf1y9R3ED4lEsoj8/aFSG7+CWUkNa+JrNDr0/
e+o2eEMWe9IXXgQ2G7uAR6m4GicgK6Ir58+8PUH0wO13UmQhbbmpSB5JawW8DopZEhlK2J/31Rm3
N3EXuObeyY0bfdrrKwy57Feb1lhHGzhbIKTLRuDxgWmg4YPGNRrSNAMbM/lLk2e6yjI3J7eDjasW
j3tvgKxcBR1UXIVrkqfhSqhWZWLyqwnOi1t+LAVsKulND5Kbg4fg8RBwAwfo2SqD8HCTd8Nxz396
x5lX4tYj+O6FEz8fgkxqXhmojHDfEwI1NH2Os6mSGT7rp0eBRW+0rpP1aHBBMBoE3ECcKzm1IyVP
osFME0tIr5OCLSXXqu7XDnAHJ561tvE8YiWxP2j71N6/hePni99n6Pkw541HmvwuV8upylxwdasF
EMjLw/L5qk/kK+3NEPDN1YsKLLG83vjYQj7THFs62jg7gxMGmAhZ25wt+W0lLvsLH3IlYOhgdyTe
VVpAuBpbCIenrioLMshHAg9Gy+LgKh7M5YQN0qCFu1F3b4OG9ZAwC6EQ4YAL5Pw0hboOm5FiyAUO
NB/7qyYHYab5qdJwSehGPnTPKGkPoazYzF/rHwSZllU2fqaN49btGgBbBTSkjjZgirmXLJp/EX78
d0VMYxANlwqBMrLuDRZfs3nEGZP1i5rQerEvvB+icW7XXWKy413BN2+uzWPik4ONzuOHEAwinaaX
bGMfl3i7gPL+3raePSbijL4/NdH5gXJkAEpeOBWwTvp4gtIUeBBPf9n+8MhFAAjBZkabHCobBuic
A27FphrmvOQS9Eqn2ji0SLYWgtQ+lnM/+GhBi6QxBETighvSBQPmcC35LfMVN4qDYUoFCLYI27Qo
iCcQk3J9XlcM+HP2HvjPxuglnQ2BA5GOAIq9g7PhsBKWeXhtVytaUfGtmv5rZvzxos9hNyzN8Zjk
ljLZzLMA2pYMVu1deETF1AH5G+BSU0cQCoxiHGMOYPD/K5RVRXpeXHatgCi0N0gyZdQpEHKs7EdT
h1hYYMnjoXZxy4JqevNo023UfAPMGjnOwQQ2yWyV0lMuXetHpSF7wSQfl/tHGXNWW2i3tuCNpGTb
qTTJWvyS0/tYWw35weufOhVvn6ctCoppXp6dA+w8zW1WAPFQRdxfyFqqY2Okg4iBOczHxE5V3m6I
HnLbmO+f2QDQ7P0Zk4RZBOyDCDXU+mgWB2X9l7Af0C2vCfkZpHnPGjTGWQHg8ToEaAuLHqzUNxm6
ill0bFEN/0rcHEJk2b7Z0Bx1STdA+jT/XYlTE7NRvXP5BTatSyiY7YdkDtpSrtIDRSkFSsqrv5Hb
4koYDA/a1th/MbcZVgIyUsa1yKnnVLX1kEFbYNAD0K0TO8T9HHZ1ttj75DYMXQe4kLKHS8tgypwo
njDZIhoWdESAbdmpU/1voBMzBDFVBEBzAyyNbRPswPVOqqnyL2E0SxhA/l37RDsXBMuKGvAX7KSW
s442tjNlYl5AtkdHAIx9glJg7dm31V3PF4SmCAZ/KRdpNHhQ7Wfk8Sd/RzRgsasRyTURI+fYuc36
QMrOjq2A0RXzzmPSM/JXIdXtl2rkj9BslRHwmZuxyE9bZuytKEv2ltvDeWc69LBfqF/wa3G0xCrC
0MtPhm8YUCUixT+vZd/s3lwauTEiIx525HKlIVEDBz2Ohan0j10CtC+yNkxgf83ZIRNOTIpzoDBl
U5aXRZLZh9IfzDXiuY3EvezVd1dN7aA05skNR/d9lxMUMOUBQdMf2b3TJZdwMuLlbHcq2bxrXyqb
1heuY6i58m+z4Cr46Ca67aqvvXBTcOj8L2R0f+usbo+cJClcXl7JNhSnum9NlADyUrp86MOaFRSF
LKB3eepzCVJEnuiopYr2s5P9WR9BAvw0TfaKHUZ4tDP13fph3vwFAT6yRgRz2IgcdmLmPEBcxaSx
DOrzm4ZNFhFY6vEF1b6+ax7CjfwbXfvW1lyc4mTgybi0qKubo5IvoDPmshLHOMvQwnLXXIOhd516
+WhkJYdIRqqHHzE0xBlshK/69UcmRC6FWUkALbapebM1NcR2V9sZzls4m/Uylv4fpJofDYYt+9SG
yWJfbZg8cyBTONa70FhppWipbXmFwtOgApMOQDYOZS8yv2PouceLlm87UkkPoicKEoA3ArRiCXhm
/VnB0EzNwPrNosa8VeAdFM0vIqw2DtaFDUEZvsSilYWB/kU0csmPuIP3hJYmaEe7qqv6/Leyvzp/
VV02eLWfcDXMBY3MOm/spRDEbSxjMmGOLZHDa6RPLKR/5ZozltK0NlXHGOXHAkg+EPrvf/4iKDhh
OiFqjws0B/skbWqWffMweiAod+Vdcm1WAHZEktRmoYG+j8+d9OoCI8MUEdKPQMM6Yk+704Hu2q6X
wKvknmBAbAX8DgosVyqVbVEH8mh8axXnx2O0x+lqeguPyzMh1/1hl8D6zfHY+A/GZFUZCu4X/MzD
NoFiO8t2redtRNcCkmkjTYo5IFRDngln9vF2JWsX/OwIedupfRggffUBJeZbx+a7rOC/wRfQPvSn
6fXP9LopJ5QOlJC8+UsG3cqanCRh2FGvdmuTfm5tNginrdhUHvpuy7RXafNowUl8ClSmHP4rthVT
xgjmVxLhR5wICeLrdL5C19FeMQaq0JP7zkcB7q7VMec1mdHOR1kznAHSYzhk5iT4mxnyKgyCjnrT
DYd2KoVOLcTzSSBP8a+5oHGJdlaHxICbHK5P4gS+NHCJb3H/TeG5kFTtCZaMEbiZYxKgQGW9BXeA
S2LyQkAZvoQuVAQdzkqxm79++2rlIBaFaWRcB40VCUQSwdZ3SCNZ8kX8GFBbSze86+2I76TVsHJ2
YPPweN0X274PnS+tQbeopzovwBxMJQ3AG/6RQD0No7ZVO5A7NFs/6GrfD6IErhU+Z4CkutEg8qfL
G0ISMn73UVoZzaBABG+KGANa8P6o3bVfy6tbsS2vhE3qLf2/4H6+V4gYrSGFgS7HWQ47V6rTAdIs
qol1rOoW1+NVoP4jYWiGn1pifcxdOH9iPNVQYMcnvWbQN8iwT9Bht3HyPtV3ubEzrjj4JcINQmUY
NFmmIscbUvkdXu5cpHdvfhnK7oIanCTrCh9chGoayKmRRkkrDZXjF0kiTt0mpEnBrUmQ8QIi/8zk
4lBvey3aicMDl5HMe7Ba8fUNpfNjyU+qJCdOVI+/kjZQOVE0oZ/5U5b772n/OrzFvyRMpolT50mC
F4iGUBnXeqsUAKc8C90iDXMjCx8qzxHwGIejb+GylGsme6ArH/N39j+AuvyUwi+oxU2pjFA1sp9W
ZXfpffk/nqI71OymWFOQFiK7aHdQsfcfYHnaQPdsfQMqVZKqXS4z0a/vmlV3ttGgCxtR7uuppeK8
d4fcAU58VbO8jEDZDwbJrUmOGDTtig7BN/SrBAxzKM+p4OlUU6rlDKxMJMnvnHNoJcwZmfAvzZ3z
l7YR0XY6OvzwTc1Nx8cxYYRZsFLFNSYDJQab677ev/pjTqms4YCbuHzKF5z3EJ6f+hqMsxzLaA2w
9yD3ZbHPM2X2kVDwZlv9i4IOO5YvKP3qW1N8GMZD+Got3Hkgl7wBE0HKXNwx/HchTRRQV7fP/D09
7grWmIjm0qStikvSktRmKBkNbdpoEU0KeVxcj2SJF18BzPge+pYTcZi4qGCWndp+GjIuFBb4v0Wh
n/Cz9U6eCxW6Ca/JvKF9JF7IimSEdDYGLRZ0TAzx+r5BBclsBInNDL5qQ8WmJUkUFNP0YZcV0iPP
qMFVhYD9u9PDHHaNXg4zNCoID363Ow2X7LWKc6TcTxMKDAFpthE4SdXiOEqJ6DhXj4+sXuyji3An
f9JYXrYuHtLpJ4WcMkPqVrHFQMbg0xh1ghWigifCeT0RacPbghY/0uRe21XMl8uI24nsbnD4SRQW
0E+vNHDaqW19I5YdgJWvy1QXGi70J0CH6sSVf/+kx7n20qSGexhpX1s3HJDmW/o+Ohg/pldM/Hw0
bORYHYzKFbXXMoEWYQZHAkFt6boycqsosS4mvsF5t7I94HNFhb9VH8oUqlsYC8QlXervJz925lzq
JAGiMElEP0nOUEy5/9P/ssYr6JLeNDnyhFXyPgN+mpcaNlaWHhVyjXjqXnOWMtUqozQApM863Kbv
aEE07WCDIgMEwpCtfJoB5gt7MyNuKwZX8JCHFQCr0+W1HlzjfIet9lKobiFrqaauk9P7rEeYqW/n
UOwaN2KzEElfLN5mGhl6dveMbq5Vd4lY9NolnEah25w9qUB+C5g661l09nxhwhVV8K186Fi4jd6X
b+D75ZPqhOZUpYWxmNnnDptzSMcyLTI4xUnDP0G3d3Bk/c4je0H7UBnrKDW8ozbQLVCIl3+vYEV2
xAlDQXb2fI6uQLg+/RiAdNLdZWWzI0YdhtUD86zC+hQR7OG15b/NPQdVJXD3GvUeeZDmMay73bo5
2PYbWqZ/2i0LKC3ezwDWJXi6psgB3aOxQBRbuD1muJLirT1AUMItcDIwWkHms8xmSy40Bmb3WbIm
KN1XWCohm0qeWXjaAoR7YXlCVhSvWEQxPyElcJr2DvtvjewEqYIcuhzEJC7jn9RmI3/vxMiez3aG
TThQ3iN9ZZMkJemf5JHW6HL8qqvj4LVvSZegkZbZ9A1Kib8NfxkT5JFeccCUAB41wyt9OrxdXYAH
lzH5azBljT0a2dT24MSacmw1J/C3emqOsDsbYh2u5oV4lIj6vJ8eratskpeC3mh1NSSyxbsi9vUS
uvi8jdWjb1oqPFdsDU3g8lubx/BbGLKBQYFa/scIRIRIo7H1wV4FkYMaR1112MQGJdq0gc10eGrW
Cz1UXVaFfCtKx+5R1hvlUZPG49e34LfitbHMBWnwmVotLtX68Fq1KZCfXmqmhWHWaBLN9CfxJlQe
atGi9svGT/Ya0+WYnvGBZCwuMW89ti8vdEAPdWo+6TXYdixbCcXmfWPl43+Cv3UyFvIATQ0zgJLQ
E/aVajDTRXtE0TPp6vQLxx8rlry8OsQI+jVHmugOQiNX+ce1WxVTsxYGszXQEolRbMTxObdZIWmJ
dBHfhX4/Z0k42gPyc8OCRB9B46P88tq8ynhMbK8rg8yalZDHS4tfjcBNjAM/FZ3065YIY0K1vKmJ
1akIVKbEubQgPHL597oUneccQ6ERxGx4LmLmvTzXZTW6il7YRKYZr0Ai3Vrap+eqRlyySqKHZSu+
Vl9tR4YcpLUKNS+tFKZDrKGgjyEEDyCXysCeb3TJsQNwxpyj+sbF8jvh7z4h0RwKImiSguxdnoSI
4KwQ9gmQV37rdsgsavye6MdbEusQ+wh3CR6EA3Hhe/p7CPtN11SHXItAlOXxkoybFZLD8uhu55FL
GC3UU/9tKZ6WmCOuiN0TaElyWLDE6ooQ//giu8OCOA29WXT5cRjZ01nSFCgJDIZ7uF5S3uhjgscM
ZAjpWegyvotkmQ6dk61K2NLj9bAzjuZ9tIAmYh2dApFxPFQBQKt7g6f+m4dskyxnbATO3IsfBbqW
xMfeazsWhXuAVVJsi8kG5my4VHMt6JMtsOz/jD4OfISY8G8Dr5WlUZwVVEoqIQMXj0WAAUhuIT4B
QkWpWo8jlsJd1D4msfOBluaGMNK34OQDknc9PWpTpez6uujZnCE5rP0LuPXuxsJsCTBD8qaGZYUO
jwMcw5xtnInVtk050RD21GorPorAsB54O8lon0BOwhRCmorM1kSBUYWhGipDj+PRTprna9DDdL3L
t14HAv2geKf+fbEGH1wZsS/wEebGtFr3RsfU64KMZKiB6b9U2fEUQv0LNgq9ttshKNZ6rPxsyA86
BuSy2txmOYpjFy3ibKDKTMgDzBCivKWJ1iPQ6YuQCmzr21vwky+cQojhBBIKHJMw+RjLqfD60HUp
cJ5lyaD6Xy1hednQ+9Acn9QnnNgfHavBJ8pzphKIXfWtFZTUeYreRy/OpNL03XVVHV05BNbheBR5
/r8ApmVvWbmqU4tkgJZuGtpXCyAduYqwIYpgZ/tM53rimSVQ4QmmAHhb1rudaSWcB3Euz6jPb1vb
HKiEwv3WPxa+nR/RZ1Uv1Tc/GP4gmrHlsKzpLM5WYzdjD9/+Crd7K5HGOEovWW6I15vfQuESpFA9
hEOXAstQLX7IiqwXhZ4lyGjGomgBlwgujlkKkbMen6vke7kovSfauczF3S1vLuh+EXGDNQoJiLKi
W3JLswdjIZ0iHEL0p2cwrKEQegx4gMR7HH/xCqc+njQS5/XmSrGnnzD/Zj8jAY+AuRC8u6eniJkd
iyKubZ794P5F/nAyjM23ZPHa2GW7vtxh5Q+krHW03cQmh/ItA5a+KnsZ/FFgGcHaA54pDEHiUxYS
l6r38AXKP4YKiTZ9hXFeCVyQto4t8nBjG6+H68PcUnqviX/EUG+gzmc67Wjqh4hUAxITOEvzBuvx
XaerFw36jVvygPtGAoiSCSt7PyZmgUBa5Tfy80n7hIJVD8kuihvC7m/v1EmpiJ2aFXiXQHE+AH7M
RKH83QboLXEtPVsrzNNqqWVQQ5HAUNomvnzzQD3arJy1QTHuPwQulVNJSEWHsDCLJB6YbSfawReW
LcjEHVMUr6RYsOD1OaZNoQMHbqrioubRZ9XXCks8WPxf1bJBW9qdkKVomeuauwMJXKE8bDX3Bp3i
QTbfrFXzCQqWEwESc/r7ue6KQCIAKPf8/OKjJOQhPBYo9h0YzHCPKUKmE/o7ILdCn6WcaG/o7/+n
Diu3sKkxRWPVsjbzbRE3bAGKUPAKTGMJTbAEzVe65o9tobvMfuGGfrp+IiW5eJLlWrGsKQv6DglT
WgTwGSxt0Sfhb7E1i9+PvFDMT3y/F5Kz3O1XgCllUMM2vJ/wHzJ31mSVLtICU1uZpw2LzEzM0cHE
xKBuGFunBa16BLq/vJMEsxFYqbUrkioeCwwZLz14qoG/Ncuuv4R46Oh/U1kcFMf+D2+AZK3MECZk
6xfh/K98YgusE02I2uoCu1bHBYu212rl7Fy/Q/U/3J8idQLHbCfg7IkCZarySIGYW0JYYwcrV37B
t8NgF3yw/j5NBn4Oe3moXXzqpc+GrFNe4bV1WwDHR5nsnfa4kxsUQg7P+Qk7/LCyid0v/SW42LH8
kx7mb/cC4oWQxi7lhGWY+S2x109VYo3BrGczq4B868U4mKYM6oPdcEzGxcbwHid1U20t0iH/WxnF
vadQfSFBgjhL4j623jqj3E0PVwV/hG7QxTP39jb3PKlG7oLN8HYn++ctSnhTS9PwmJz88tZ6BZpP
Jv6aPvT5gRCCmJuBIL0n9iKcUxyclUKAtpPhFGF0G0fexgA3AOLjH2Cg4Kt5lw4opHDwR4TVxItk
kOFvZtnkiBkoY6YsDcCYvPO24+RXDAArCnhTpEnZ5tupQQNqX4J/xJrnHvKj5vKmQAlwH7zPcV1z
wL+s1MPffA8nDD8HufQWWqt18EHxHZxSfE3JL1GrZZqtjve2ChzXXmPK2q0PZLHW9lCW4q8o+Pxv
K+VvkxzKdi8Kf/fuzhiaQgs1D2OpOmQcwe/lWWBrSgbqjn8j4u9RANQoV4CAD+fuePpyBtXLTS36
rKWAozV6o3FDYJSqQpDMeAmHYP3WboHBIr/Zj6ltmHTbwlMxENsgFGfeuOYDBdferteYdswFk0Nz
MjETaGlNPOPbDfUPQQzgZAaE41AUf8014i28mq3Cv7EtsXW9YJrQRrAs0Rvd5QfhtxtIiqcnOg9N
RB4m1SlsUFncC+StcwZWi6CaBZzxrVPw4TdPaBeQ4cDdSFfYJ8u8DUVT75Bg68UDnuuv3CJCADbr
U8AD8caK1hHppGJDIH1vtW0szle9tNrX8dN6WVoSk/VANAmt/PYpAeJ3lsKRTC989qP2cjgFu9d0
6OFa24EmWxOGzIiYci0uPxkxjZbTKHon88CW5uyOmu5kIBO7HHt8gwyVzxzil9/8i/yXLer+WSSa
084xf46TPWWiaTxSqOuEflpEKB6hCjXkNLb8QVTJmK59y5LrsMVmwb5Xxg2bS5zzZVTjnB3zcTDJ
WZgY/qvpunoPCcQB0cNmIDc2SnjUB0U3qcarZqWpqfaopXoYPFlEEBzHP8pOAdCPa9wU5ztiJK9x
W5OvP4uZOGD4u8mLhpoHM6FgTVDEb+vaaGkKkeXs6foTh1Kqa6KZlGmqhQlmlqji6k4n5MsOiMlE
WJmFwGbs3T0JhvnUqpoOLYv7L2dYzCMhrlJaIm0xl9QcPXXzeqIQG5mMEo1GuZmK5u03pnG+UDqm
WF5S5/sOQL5o9m/h4YMhPcrlUWW0GcG3zwI+ltWVhKXEXMcU1HUHn7tjOJqm65FhAcRYu30qzsEh
TO8yuD1WdgNzXRrl5b7FkqjD72vPmHw637EpPcttoRNacuYrfrEgS4qydT0q04Rl94MK6jE7Psc/
BXfJTx3sgQPfb6RyfgIJxJ1LgnDMlNGUcJljrnfiHSlH8mq2W2fhYSyiCtp1GfgfJs2xJygMH67z
xZCSfBnLfEpdn4vMVqe6BZWmK79QMzaMeVMk0fGF1CBqKBzzoVOGW3D2Tt+/njOebl0zAvwmF77y
qP2UaqxdHAxdwiU4sBlef91NwNu2BJcjZ07KoAXbjsH0JM3WHaP41QTe2eE+IWG6kPomUyUMYsTg
9z42sIozD8EXckErpsSR458iKHnGURHvR5qYd63xjOEKkQ6qRveedP1k7b/jAnvWKWyC7SWsXcej
jgckxpIRrP8jTXj5yoWEoBsuN2I1cI5KfkhKSmHMk+8ZCfyNVaJ1gnB8EBfHOaR6kgbBQ/7wU3iM
EHQ7THsqgP1D34tREaeuKaBMmgjhXf7UMTWXZSsw16h1ltWK0tn6lBVCbhvKZwBTteblX7+2ejRh
ED/JlyWtRK/SmoS9KJwj3ne2PDP6qE+E5eoA/+kQm/dHnfi2DOFFEEcKkU48nni6Om/grnQlMiS/
u43hHwMloXbN8oSSC1AIPWYoHDGBWjGySn62UbKAIjER0/XmzG9akoy3uV+tAThXgFefI+MFrT4w
VoT6VV+Ou57cqyNSjSOQtX/tc8jmp2BL2Y1ATjIsgM4k8/jIIwQKyrSo4wf6mP3wltLIyfSQz4l2
yrr9yVGf7bVNFF6CeRwJErhUDeikQwDX68zupCzc9RRJBq41Katvc/v0435+dUtychRyCM69NFNu
MRsT22HtTDoJg3oewVCJZAE8EceLwutuzi/Pu7p8AKUjAf0smxE3DerTBITFlBXcSz0MESBkrno9
IVH4zt+i90QdqVAY4CI4Z7epWwuZ6l9NMYj3jEeMMYmKQxDfZCEYtKvxnwiUamUxPUZowj5V8BXo
dfOJWY+krXo9K/UosvQHVDAQMI/LlFnHNdhumQeC4Jlpy9H++c9G0AqiETDsf28rsAPkqlgF2WEF
I1Hc6ExSwEpDvFRH8V8GwT4vgp8rrXAVw7AOa9mWgZ1u0eJt9ZBehZ8sDI3t5D5oCZUzg2Vh1IBC
h00YWVFlSDBWYyCtCsOD/2JJebuNAv/iR0m0gDkqBifzm/HnJL9ADoriiJ9MjBTB0vdutZMy12s4
ybAB1ufzswaqMYVdIeZGxR0U1Ix5L3jbtdIvvqhxMxjGJd+Zd+L/VG0tQFZrbaKICEIyWHZSP31L
vmjT+iErU9tOjlaeK50jC8sfr8ekN2soXBWAgNX4AO/L8fHJK9V4zKMBKL0SM0Ky3/inOPTdj8Qh
SW0FSobn2wuV+e8SO88eb4ldALnrWA79gabg4cFgVXF/hzrpFdnudKZGToiRZV6ctP2EPhkzgqkW
/16tiZFlFsfSeHwZIXAEg23txMtuKhCEdaayimzk5aWVeboAkvPzHMYLrfPqbLdm+Ju/93EVKyF+
FTe4aqGsePnOLposdWwOGR1De3Ggm8zcItdSlWwMs/eTFbufZumK7Zhki1WPCaY8y5RSeyhvyS5M
fP1UgE54EjKynzaVkNN60rtl2KBmwQAqVYXn8pAYeH5PTODclrYFLZwmWtTpYfqT3L/fH2jjv4HG
mHJuJo2Lfz8hgQkJCjPsIsAhTLfbUUJvC8xisCp9CTKTKw2VkPNL0kOru08yHbeQtPNFzeHIIQQX
OJKAV20u1H3767WbkjF2o2lOEPhU3wehT88+4gSGlgTOYxugI72XLS23NqcscJ9rO/yvH7Ky/OCA
iCEA4COwfoYIbEm4ROzFKK+/GZOaZHTGyC7Ypz571Q00ajm7LodzCSmJbh9Xqc1qK8PQuZCf/elj
6zy6MXhvnKLF4pkf5hk7bhsJ2WQc0OExC1Thcg1EFzPPZx51LwYeLq6uaGmPWXH2PlMS1tIjkFVQ
iSuydV/lQXzE32SqCR7+Hm76Vn4G1HIECJqIqaAUGrqHGZ37Ul61bm23fxjBhPKQKcsuvkkT+7UI
z0LPEFxZUjGw9SwiiH0DcyeOrDkSjJXS0whreCEYOJPVPGBo6sdLQ1eAvtiLQ+cWOHp9TmwDv8x0
k2ZZSnDSgXxZ5dU599s6GpscQo23bwftRSPnFLg9pbETAzW0NxK6HWdm9jUFqi34YMpVnRKNIhPO
/T6m/Fft0xBlZ80NLmukdCSdmgjcDcNWjQaFQbJ8PjbI9gUKTRXlRPybMZnINODrAyIOR9Jmunec
Y3DX8mS8jBb5tSAQrol9R5Eayyun/Vp63UQTvL4mXJ59cgAk12DErjFvcMa/W8T5JC1jb6sBX2J8
n75gKH8FJbP2MSqE5UUOFOXvLq7pPpSbLOUV6E3GL1GywzJCjT3xqMYH4XDOaNWrU7ZCuLybXmFt
Hq2LnZ45rLSE0h6R902fjfm9hGGI9kjikpNRw5cKS0J7gLPooz/v1eEvOlkzJRcTqI/Mo61bJ0Q6
s+2nDdDNFTGkPAEvTvmSqbaKpkgNaALpqyDW+qJ5k8ScFGiAZC+hFWrzWzwzOlMPGYPS3fHahprx
umRlUUqzq2T+zLNTCUBAUw4vR5SOX9OANbeVzNrrXQFMN8MTtvcRrlE+8ILfCMSaC0uAro1LSAnT
gEUue2thXbvxrN2pLHaHKy05NaT+aFmgn5K+5Kwe1VAqmFLwbLtB6dWMPGHLNPOlusc6rCFFC5lY
InIIpVNdBiJ1YLMG1XYOi/Yh4OBJcFI7uvAC7ecMylgV5RHfKnfDbhYFSsmIEYPeQWZ2Mlgza519
3EKOE/NMTECYI6kaOSN04kSsvZKDTGBJAdvxlq1BMde0ufUYuSJnXUaiYEDGU3bVpFDfULZop0mm
hU7aH1CSWHTXwa5c2+hl8kXUb1QS7I8wU1hNK7gtnktFxsG/2qav+VoYKy4cG/wmg/Ci/U6o0gI/
9OoIAKkL6IMO2rCXdPTzl3Hw/IHttSsKRRgyBS4Mv5TuWjSC9gHnktogzEbOOlyIfx8f/k0eC8Wc
M65Y6WQEij3mq+n9QiT0CF6Ls4ASBF8ynlZmFnkX2HvWNrGK2i5CB/wRC8nE2iJ6SP+aeyHr4Ydq
hFm2cNd1aEfJE8rI1Cu1+8K+6BKVkns1g4AjPW2MgoF8AFMzi8cwKP50Qe0Fmq5Qedt5wn1epTds
9gNJweBrKJYKSfRDBheQFZnpjRYJByaA+EK5XOI7Rb9ayJ/FpijzvbpcxXXhwBFLm7iAb9+sMc+4
lJTDf1usdArPZ8ZaXNOyEVOLd7CXQ65HkxxM5+DR8kusQEfFv6cCb9pvriy8/bfjolnyPuJp4rlw
eAFejKJhf3NYg4NOKqziHVZV/BtY9MRJAien1ZnPwgNWdrpJGA+dUS/gc/Se2Znhy47GHuGb56+T
G7/OS/SrrpbElH7u9IBDIQP0TKWl1lzLM5bYeS3O7VQVHUIrAT/B2nwAee+vJhv7PrR7QCCdgctE
96iu3LLzi26loJHUP7t1+SVr0TOfth5v25IgyqIV2io3VbaZ+Zg85mFEqFS4RUrcbi3QNd39BMmc
YmJzq5PH490EY+z0fvX3ieiuLr2kQ/l6LJEruj1OZSNggW+vgb7PodL3vdxiETo2Q2WO/1DFcfpC
QrZu4C9Y+iFolS1Mndb0eumsk7/771G+fuFtcrjIvJMDfr5QVz/3+oh3CjgLLsqX26KhGG5NrAzF
dgH+BHePLdBcSnEmJv/G44l6doaU2yBEv6pKpymfdmb+3BnLRbjm3bTd4Cby74qgZ28CxscrPtsn
hknO/MwNZLE1is5clYN6Ro/KFZdbdDF/546W24SdVVyvzpTNKLzMYH+BD/85ryouCf2k6JBKPYgS
xLqRaxjsAvEHXPGMzgZOyNr2HXzADGTGhRnGOmyF8tCP5gBc4Zx8lB3svjS34rOHTuxXmRPHc/wV
cdkiFDCRjYVm0Z1paNalZhuBKByUaZl5x7Qzs9uGfr7hn6TxNhlG1dXyKiiMob+ZMcI/Qj0XoIpE
wMHQuvvDuAv+GpayhuCU6Mg+OqmujDJxFDyLSLreHT/yHcy1v/o9BsfiCkhxC634Z0Vh1QLhmF8x
28Xec7aC4q9i93RPDFi7dx+3/QW7QRts8Z+Or5bVVRUHfMJ/Tx6cQIWe37zp+yLraIICwA7K4VDm
7/p27I42UHiDhpfO350CtlWqrV/O2MEk5oZ7ViLYPAojomoqJ3fWAkdjx/ZD5HtsQ4Sh8CaiKA6q
JxQbDfoNIZwwPtdr8QSpx+WR7cm2wh7NU7DQ9ekSMNe17r85ChBN/uMIQi+oVq76zwrDFccmDXhk
gVDFBprjaA5mWiUyp7HtRo1TROt9cIrKTikZ5M5e5QKrtIf9Rou2+92YxNEW1Xp/GC736BIm4/Ac
ZJp98BXr+9VZa4IZqdE6l4ih0bnqryuzFkzQrix00lulKvDz4XvetJhf9Zu9QcFgGUActrvYPwlQ
gbmv04rrP44xwjxW91gvaSf5VdOXagbku2b7fzhKpiKGCPNHT3Jz+JGOhsdW5nHEeuAl+vAeJu4Y
3WmW20uJ4lu2rbVReGy3sXcp5CGidQQCSR6d2pYs7cT5U7/XjDzOCUGwCDBwsPlUaNoSsGHUzgBR
b80H+XmX6xy+r+wPBP+jxzBGeFtwRoqDQGc/w6A005nMWoxFfZ+mUyQXTrgRkAAM3NfjEmu6gwHx
g/2NsWyTCopambhRP3Rkvv8qEpiJtoGoLVFVW9wBYFBepXFOkvDFWK/8c2j++/wwj02Kr7UHEj7T
zR2RV9bfhMKZUeEhj/1Tl6qlVF7rhhdcAjhRceOraJfrniIVTnTnNhQNWcZ5hQDizUpgDkbJVmEu
oVjTwoVOEQxxCI9H95n3FKh6EJSpS/h2MFtIgtW/yfXu9k/bFtveBXmM5xQKNqdHLnaO9nzXnQAN
3H2R1916NeTvxetLojMLeeCpDMy9lGEKWdeUabAMTJyhVluaNsxF4CpUjqgbPGJfTmeHM4a77jI6
vLmDJdc7z9QKvVV5/6p2aGl14USA+lvWn3AP31sDMHIzigZEJd5zrE9QpHoPObGvvN/mL/rwt44n
nRr0rj+l71m5FLTJ7InVQrvQIDIMr7kzU5MbmKlkjeRLLpO1OA47eCUqZXVxbndl8ImcA+yaGGPS
WcgusBifJ4EeNruBpyYzK291JxJMu55HFlLhkB2IcGStmTubv0RQSSB0GhGBYlJ6ejUU3U76SKxF
WZNGJlKNP+vZCKX4aoKJ8c3rreUkdVPQ/4aAFhUWpEkG75wQoazQgDeDvuDGjvLDj+iL/nTpqRSv
hqxaNqim4NcDoW4fd03NzTF8BHjmW8QrsLLAzjjTmgqQ8qcRiDQGwY+fFXMS6yxZJMlHHtEAOfeS
CjQW6SyP1jJ34UjcBvFuFAbGK/FrOWIQqJb/pKJT1cI8l009FvMuO7d/JC182mMtAk/dopR12uJL
4uJSdb4rqHtfqPrpKzR4TUH1RqbqTIjBPV8PvoGiFacZmUC1bSX1vd87/QJQ6gecPSLuR2YVWUup
KxsKPQKYQpe1KjDL1Fgzh00DZ5I1pYapTB0Nf+3BpDo6pupu6gJakYw3PmkS3AnauRVHztP7kt/O
HMmZKOiMnX0kRMgtS22ulYAZwj9zDuMtQUJnHxBcFKBWC01rxWULXgfqdsIZhWiVw3nBxGE4y629
Qm6AwFwvJC7hEN/gwFje+Zo/+g2hbyvCXFPrFqfQ+LgKNh6J2O+05pSq0jUIz3TQAlOVmd/nXPZc
ULKPwt3vWy2dDZy3tOxFsPxFlakyaobph2j1v0ARcnEv6vi71ERgL9zwzVUKi+qeKKqJzPTPfCC0
Mv0XG+tg8EQglA7yPN0MhckKKrnwMeVbkHDWHMrrBAI4TM5DeiJAgEYxWdvVTcRdpesTg40hCCUH
SVf51mw+wfUFJazmcc8Wdh59YMYzPMuzg0TJw1boozOzSVdE9TgnX3JAz2W/uK+fzMj4byBuGUbJ
jzKKlJytqcPJPlYWlB/R8GdHS4Rt8ByiN0UB2RXiwJoiuuIWfjIEzGK3R6gEKrGfxy1NtVUlSheZ
HkQ4qi4rr1WIgqfSw+YfLEdFI/c+PbAtqU8mPxHCStFuKSvXcOLaH6WSYZdGpQXdJEckeNDdp7Fb
MwMK9H9+Tts/NM3TKKcdlhQzTalNfOmj9xeXBf4u28Z/yBEYe+en63EnPPF25H5JV32t6vlRGZy5
O1MZZS+L23n5WgDqaESNsd2Q95jXg9vsAAif1LUSgaU9/3XpsKRuvRkX5X4wgKoDJEa6o7IKw3nD
szc2KOYjpn2sUT5GOKc7epBZ12DbnaC46cjdacwF+MyApsoXZOjgXfAJyts7FS+AmF+VioT0f3D3
4Nxl3oZZHRfNbNj7b+ZSS4HcnGQgmKixA30U1r3R8z/hPukJ7caVm5rW86U+XZGxDw+kLljaLgO/
NvIBttVL9mCTydI+7ZnQ9P0is0oAg1Wkaf/Q12DoWaV9Ibe6F+kpo0JaMQHfiLHr82BxuCLWfLQ+
eI+jfKyCDTAOH998T8wZtnoO5WBzcAnP14ybzdnj1+BBwoG49l44vD1Rkk3hLZjtWwQl6rX314xJ
9u8GEWtw/7nour7muFh3mwV29o3+YhBWYoSkex7EQeC0mQ9qlXzBzOCL4cowF3bzI2g/iSN9YXx+
5PpS4YZmIk38rKxT3rKaOB9bixGK9lao813uIyTKGu1N+leoXYgwCfVySMnqqFmkJ8WKz/9eXoFk
Xf11wm5wD6FMZKIYQxfH53zaUHBAlcNM0z90wcE5soBlfPjVT/gaW8gc1VLde2ba8SCImcUtc/Bx
L8I3qSErzQSmq763zRiTzGbDZH6FazvGnwza9YImBolD/41QJZO6K3Wi9ZdvHP7u2xFbH3GK2SE8
Z78O7Gq1b6X7jt7WCdvRcb4wKSgtqs9I30Xy/tHpIguePTdezSzgLoO6gjhfSVZQnQyMCPIVgo1U
OHDqVi72UeUv91u20Te6ILq6LyyY/8ARizeQIMVTU+d4BrZfhP9kkFDy2MBFFmQcIsD9QFnCRAnc
q/82drlOTvczVIcmvuOFIE+lB+AulxsezpqmvXN41gug1lk+uZWqyKM2+lM/WcitD4RMQvvWk1p7
/WYdAbbuYUGOTJPPONEu30HylM+wJm1tjt2Ycr4mdV/DVCEPhjqvMCtiiMM8YyJ+26wBwiUboVlM
ObbdBHUFtml3CmiG6b98tzBDP8TFmYQOSNJJSexZl8SHv7bTI/DJNeR3VT03wPexy3h9AkwTBAC4
MfH5jwrSxWJnk9/+JbKPZw+kgt5PnIzEhQzgCPwoxFwd7bIlXE9k9js1wVEBq3HiWVQg1Wk//0M6
GsJro4Ktuj1X2dyKLLb4EAzuEUsuZEeGdEPVHty4p75Ok6ndOMd500A4GZaTc2TMvnb3wfNILH1t
U5ECcY7WGge+61VL++qh6NQG+eAOPgWe38nrLwcNtKL60syOW/uec5fXt6AmXoeTO7CbJ7F/0WEw
1GOUwBXYlQrlf59D0H571gwDrVnWbcLhzRou732wU2QKO2hpu/ucwTgsXAqe70vZYsaC6fZ8sJ7E
uDFOul0L8ekDcXIHbRDh2h8TGCTf/76Vj9tCfnh00r05vGUfOINc2e9kfuEyep4t+qR5mtZkx6G+
kdlgnKxCDEFjOpajog4yaqFn+WgA7nxI8vrMCUC5LUSJFSTanbgzrwors1pXR5ytSAZgckNdaMGN
KWTGl83veqUeKbjOWTene1nr0vE/WoVp39vYCXBuQfKiW/NjScu6fl6bW9rKnNh1JWs/C8KquRhi
uYwD1vUNFqaCSP1sS4aBGQwygMyclGohw7EjU5K216ld0/fVe+0sysJyCZbSWEtGy4ttrAp1/UFc
8A/fG8wKi6VxlNqB+NBcfPYar0a1NNGnGDwM6+9AVJquSSPnVMWNz2YcTVRpUVLFKMYJCiPMA/7Y
i8AcEbrTV3n7H3nGZhRtMS817CPNxXM66MtjnnMBfB8L6QwEf9ddIN2ql0wHSwP+ow2qTDdkoJeF
NePbCsSH97ibKqQj1CSKPd1KJGMdh03edMCR6ZuLKkuOgQf3yWTypxIZW45zs6GIfsn99nuvmHBT
eHnJNdhpQGn8XiiuoYU4GbmazjFDjH673y9D8zarN4DyjCMS06rw1FQpFYDpIfKyV9YVNBh6XQgl
gLSGYzBXzQQ1WCdUr6ItUIuCzueFkWpn3HTE3kauzOgwL/Zp7IyaaCxBU77APZbIffotZ+pt1XVj
dYj4PCSTdegNaDxcCNhGKcvuQplnaQkc3sNPstbkkDITn/Xp3MgGeHT77O34nL3yxrTDvAjLaccq
O7rpwzj5IWZzfl01RKKJD25uCqgFbtRM2WZElA1K9I/Ux02Hn3L+VvWBzFf99+f27fBvq9re3bW4
WPX5KGBeaMwKLRP3LJoWioPQ4Wye5tzSX500zc1iajY3RYcaDN8UZTax29uOKQ0lHTJHZgVLKI2D
1nCa7X0TMHHRRs8wmGG8GXT5uiYV6Rt+9d2C8h/BRk80KH5IEo2cuc0cRldxi66L/ENbnCy7tDQF
hBdYPaeQm6D9v30T1uCv7x0P9V628Ry+C9E59+kYU/w+xed4LpmD6VcWjXjiDiLfyZ1aKvvc206k
tl9HJk3iOqzxecxCdcAlsAPDvV7VblC5FdtNpj7o8kSwUR/u8MG19NZFiKR3F60oq00B35c7ictf
ZG5Lk2e51P83Nar15wdBfFr4XBVHWeT9VRAYm7ABKqRsK+mMaHpHOHqaGsobqcwY5R7jX14PICgI
3pSttEXZZpGLVSrF3XOwq8JrhbV54sbaD8ttwkYHOmdT9wzm0QiCmesUzaUioIbIUSQUtDHdQ6wd
Clpjo8kZglU43yEpRe2Vo4lO/Gys1eMwVLMZs0f+X68DyfLUAt9ZAXYUUl3pCqEMjrASNsYXvWeA
fnWBXzDFxWwyxHbh6bGe+IuvqrNJ9jzOJxlcLTV7A+vYBcLZLpWS28cdzD8G0UCIY7i4ycSuiujm
r4Cu2fgWw404taEVQFPcC8d9+pBKxUajaC8AADvlU9GkTrEBov8elNLBa3sSJKmHyBk6kk7TxGod
zolsPw5cwrhgUVvRhLUNFVZRVu1veFsgn99GLsgxy5XxromKmUPc0/NebSFCY2eJQbHVBG+nL+9c
DzrhtIKvuD6fKVdDQDMbwpOR4K4b/b9s0HLBtEWSAcZZMzTcpmSsDzT0lsmTWIIhSs2vb87Bl/SJ
Eo+y6QZP0CSAK/YBEQCUGllBNsPMpas9WSgNdDtYCthIzb7JFwhVysUJ4+9qIOSillJw6ca4rDCc
tFAFnU5XNQZ8xQdOnc1zbsHeucPtg0JuVlwmCJx4z0LKSI0hix61zcFqyNSLzZcMM1YhVlNerIhQ
lMoW4LA3DMM0MagNC+jt594QKj+Cnfo2Rp70Io5TgnQEJ0k2j7er82jyCqbg3p+RvgP69d2Ua9Rt
UIi4g+fInmhhUwjDO5qNQHU5sjThhOefFo4yKZXeEsBQpR6yR6A6cq+T7kkBMCVzxKI12DXciYdD
uHaVDYuDTnSArf5hThqivURIlWfDS7qE13uyyQZnx4A/W6UL82n/txPwn+MXkAeC6bXH+PdnQ8jY
dGd+HyK/CJh5lqAriiqXvb0KcunIM1pxZEupaZONgdOUBmUipsWUh79SUuwvmT02iUkIY9es99vl
hz3sGyfQSIiW8SLaZO41/GOG8epiTRK76cl7dicfdbS8sts52OkrsefuDAzGNqE1lGPkO6BBbeHk
cyvAG1/pYtrMgL+iuOV02H8py6ZU4L/7LsLTxZtdJyUJRiM9E1/ual4VFmpSVKXY0BCXrai3HTfo
07EsMM913TwKGsSt025CXTV60xBN1yD6tfa7gjtjVbLbrw/NRlJjlpiqLmeNe/2FjFKm0LVigubh
IfCLV6FD6+mFjsl28cM7ol/Dyj2fgHmINL+I6EOoytJ60HK42T6Hqk8hM9o/SeObah3IJsiwvEFI
WHmKGg54Vu2gZRX+gn4HlT+J3GdovshWKb5pH9lfwInukRv/q/7dM58lw+K0GxMBoeZc+Ra1ohPr
TiJkGs8sZv60mNhtTPcrgezpfadNQV0Efp2kqlZlQhY9YCfJRqD8bwxJpMoBLaXioRwQwJNh4/kf
+rAbdIItACs2g6NEPcXejlxj1wMdzFYg3QD/8DqAfQ0i0iu117gDY/KfvDoTWLlBd0eJal73QNYN
oLVfMB5SjQi+KGVvd6dXWjnyIr/BYTV8VfZ9v90S9uJObmY3GhmkhF3EPPcSJyMivZ0eaaMoLxZc
3QZwm4EnJH/7IZ2IC0HIHy7pFcJR83ZGArQQp5InMksttS7Xlf91cBjeixMS0dhDvwsmSdm+xfpl
Zlic6LflunbTgUplgHSvfU0ypYuteAtL2m9bcgm9sVLjje3vemShb71rKRSz5kJddjH2ofrvlmLu
3V8ryYf2Vf7AkqCVcA5Ac08reMkrZeLPXQEOYG1nujgXSAiviF16hJIlsjvy7PxfX9VJlkrTWX0Y
bBh+rlVO3EH5mdRtxffludyE1OZ5wNbDNdbMwsUrTEi4SS5HBIAYx+AnLaNzdi34pJhEo6N1Tnif
4QS8ewjFTz95foCiOdqpTYflaM9mR3uVkZDkPuGhAN/PjTN6/mlaWkJOIk0LbRQCsutgARFTEf8l
wFmFqh8rUiTY0U3oE6MZPVuGHgSRW1wArx4qnGh/oySLmQO/STljHOlj39/aFxiguAXxxR1gyJC0
ylpY7LSDU8zxzJZyyVkQiNQ3V5WW8MyxdBsMIUp4s/llGjRqz/TSzOWHpG2eQbVQUqbJPGnjOidU
X4qplZxKRGaqDoQlOLINM3WfI5Whwy0rYEQn5yo60dKopP2VeQW1/op2kRrvHx8pzzIQujdeSsNq
b3tDLX8VynJtI4UiF9J5BMilOwTow4I992k1/aQnVvNhaaFJGgP1D+o6sGbnYOKq0zdeDBLhs9yq
33xetRHAk2DIhRcLqJqPU23p/CqSvI4IdGfjX0mX4YafrWYMQih5H+1WbYQUy8h18dz4itkS3SBH
6MEXNqRBsk1/DyHBkO9/Pfd/Oj32ywgYLO3iUAiUlKoaKgaZqY4ISLJMGjStcb7FrlS+UHUYWaNp
+2aI9TLYT5mbzOTMLmcPu0APQj1QwNKxfBZbuvz6IuG3JhI3xEV+Q6qpG7ZZHXQRnYPCUSr/qRSH
4qW8V5BvTsY5ADxHnSmXRDJAc6gjTyUnjWPAiWZvHp0dBqunf+GQ9Q5dnHxRjN4ZpIZeGfb6wdgp
ubx/w/33tWJCPG1C9LUa7gSmm0DSrCn8zYRZpLYSUosuCFGzs00EoxPcBUx3rJAvznFIMXrOhzji
q2N8WfJvalmr+og6hkGw03GIxRTswkl4ym6rV5Bs3jAt/KPuOKwqOvURVuyU9V1tvbXr8fe5dBXc
JUCsUW4FzCoQvGBXpirBOAgegRliaevc4tjrZBSJEcLMb57DYH2/HMMLZJ+1g5ytHilamKX9U5r6
X/WP8cbTa2qms4AORmBj28t8oGr2Ry3lGC5PFKpav/YMYrziMUnCMG27nab4ZQlvzQd+Uw5J4vOM
feh3vpW7ofOthF8bh4aJF4r/hBdPIyYJkjAeGxjJB01w/8MwyGtnsd2jL9DXfN0A6VJVbioq6fkA
0KRIFQDsXSKlAsdSa+ULGTqGAkeX4v0m94ewkA/0I5xwzhwKurHM+b1e80sQ7THcaruOGq9ejMMF
B2iyt1NmDtsWv0rGjC582erewg4Fi5aKiIFhU39XwMXj7uSp2jrgZfkYEJ2KCvbo/STO/e7LYD2w
owR+HvX2PzgnPWvYpsT1vUUOLIlpCydrCAeuQMGG4IF7DhziRS9Eeo2GBw3ArGzdxy2K7zcquDLc
jlek56z1vOggHdVc3yXjk7fmCfLUBiZAPNYh4yGBrs9Akpo2x49xhpQ6rhMVk5rrvcyawdb57FeH
Q31QBsnITJZKWyAwTan2ns8K7zmsVWLyjKYUOajK2d8D3LHogWkwY1R3z7Xj9c0d8TujI/KTQF4C
8svbWBK9qyrfpmHgYY6Kn8TYA2T0vusOZndjf1lu4ZD6w2n+ouNGE09iLENrEfGXEzZz4dSGooee
NF1F7ZAbwH0iky8olN8W2BznCoXC3ZW1TbBAaoWa41R9PcqC0w+/lcBf0T0sVoCUCupQOyB4Xrwl
U2gR6jMQalhhEl00jO+00m0pX413/BWCuSexuENUStHAfSPB9sRUTjdgfca3Yfk4c0DepEba5gsI
HX89QsE5rsLickUs200Ld4KEi3iVSUAasNDdbW6ARIDRy5HvUu6hyUEvIS2aOpOXBrGxE3kbGO6K
D1WSA0VdGqHBKPUC2I4QJuBhOq2X5XAWNN9Kl7sODjuVl/PtUCbn+L1YZMXrRG0iBhRfUMwI8XGi
H7BOLkYXC3BI3cW3fvG0SOVnR+xcteW3jI/zWoV/uXymq99bKS4vedHX2SmSvBIbt78o5am8k7+F
WTV/mFFxsAaYlOTqmZGjhxGqWNrcNplFbHmWpHVZrgDAEY8cE0C7m8MqdVyUDJ4QNJLs0fplp1fp
IfFEjwvxTnZ8SK1iP6u6GLg4a+XOu/YcVyiRsqrg4uf68bNXCp4PPGnKKvHgcPwT7rA3h12XJudJ
pT8MXHTZM7J4NwVXpc9xl+3uh8kC2epQZH+bxuKonHk4FUpgcbNRZleipXrNMiNur/SdMbAmTTrm
o09GtUYs997/FzdjU3RuJVhm2GjKy2788Mgqzg4TmVJPegKa3qXatxpSFM19w6vZKfc0sIunFQV1
zZZqH/A10LycDK8ePVjAEhYAcINvWAaBkxJG6eJUgEDnEAEg7wKZ1J3sddDNCYgCCFTwheObBkkB
i8MQbRY1o8QTZXxKxHMWxSeujizGXU+zQmSfxPfz+zpOHtHxWMmBsm7AH8NAZGHs3jjLFiHt8GMS
VfUmHLms5K6UVEIVDt8iVBXtTmM5UcH1LqAs4ng4AoIeEOX+GZqabCC/r2Zc8RiAOkM6A1muBBgz
s321oOXZtcSy3CyBpUg9qgDFK5Ui+2ymDalnKLjW3vdf/Sphorx3X5MgQW74azSXcZQLirf8M2uM
8IWydu0a+BdwDjf4MXyEgAnYeNFKPrCFdRQKz2JtcFkHIcZLfJEIXiIOuaIbWmvovJxyR0rlrgLA
dxNNPR+RPS6MUkjIkL2PcpiOQKrfjsIipgilLJq0khfuzjZKnxz8ewJeNalMFQ5oUt45yiH0g96a
6DweyQPmmUpR36JnJgoCHzq+84lyPhll2cQZ6XI0pSME1y5jbLFLOAo/9AsNR7TVGXo6NPXCZrLg
9W6TqYVFTtZfNYdQMEOdZf73IcGCk0Rt+Ane1oWhoi7BsM4ZK24kvU1bGdcOUkav7aMvdEjAKxLQ
/R4GQy0HVV7zpwLdM/rWvV50XaSkCWoJ2adx1QCmLkriCAQBLUZItF+8MTwJbV3CH34LUixCwlT0
mf7I4T66ABXj43rHQYLXGi7CfkEXCX7NDYnSOaJGJ2q5tcFz8ZbL3hTdCN0RA+9P+oNehp52qohE
9I7djySoSczC3tbCx6GIg+7fJTLUoj+NrlzthkjffWh5a9x+pPJmM+1Cp4vPiIyoOQOUib58r7aG
SvTciLvZACc0O71xdtkU1OXpFFwSrviNeAV+xV/ae09kF8aPWxWVDXD4npe+OWIyyVNt/aVdDPjL
a+SHTmwAMeFUqPqwnC0YsE1A+1TyxxY5hDC+HaUnhSTTcnd3VepCLXJm3yXuOziIM+JQGATyPw6j
f6fhjDrTcondX7hkti/sJWrIoPz7Fk81RIbiBzoE4aQ+KPEwAtnSF5zAll59npwnWkhuJdMbF6zq
x8kCpHP15vavGQQY1+E1sndKi/dzJIpmGYzKYISQ8Qix2Mv9D7Mv54PJz1ewCTHYcblVtxdavoDg
BrHJz2ydNQwPgJrtWAP8xh/QNO0utLCml4vB/ZIVo3ckhRjeQ96An+a6LP/zhO8ITGxxws0Pl3Jp
5QAV5xoFCuC9bLlnTAWnU6xTz69ZrqIGJL0pZGzeE2SxFtWOoaYKUH4ZpWcMiOY+ByOpetWcTb6U
MTPtmpzHhIiV+CwOgLu4JL0brue39MUZ63Rs8Nt8L4YvMAfeg3/PEw8Y0oTP4M/TUD5YNmHgb1Y3
8NpLFwv3hdfu4yH6Isp1SF/aRR0qwWRp7S2mRA3nDGuT/Q2anVrTXt++1SLSAfHCuAa9ub98sJy1
G+irxL5s4+a2JpGJ3QIbieb8fu6Xllj4e7b37BFCR0RgjpxvyJ/9+PIcFSNcSeebCJwb8xgoTzFq
/3Y9fK1FEGRRjUkc+aDdX6MheqtZxB6F07vEalTW94l52KWqPyUI885cpNOcnPVdAk0GXoVjhpgB
0xW9axZFG+VT+yAnP7byvcHl45nkuvXyQYu2e7nAg0EadLlMoP4l9vhnxTnxgIiY84K0C2lXZFhN
TE4ad8hXjNINWixDTXpkqaQ9xeM0NXtpgzyzmjgtiOWab3sRzMfExFQW2/aIseWp1XihQvW+l0cD
qQ7DJRIShXsLvl0o9HtH4o351XmMa7NwoQm3m3m+uPYStTq4UsP5VeNtn1oFmPiQr2aO6OoovGCX
N4NaHV12ZKfVcyabxBMZn/d+vaDt8pctv5JOzsCmnWE5353ZYrw4lKRkchD3TMMv69rm8o90fHdI
8du2208A1/WACsy1yV8XJ0LEyzHunmcd08BXa+r+bSSB+PTYPODHnSYt0GSJZE56j4uZvKJL4Egi
3X7pDNFejOSBFaK8grhO2QjihpgvNhGsdTx4EXvhghR5TNRw1NWR1PEfQ3/g7niqJRXSurxDnmHu
9EafmdYhuNCBGpIQDKcY7oQ9HfldHBRc1b3ct8n+OicuRrzgdOzgYpO6CStzGVwMo3RxaBHxktgF
Yp2z/4TkBXVfSGKliMpILTlufDCyhzMNHNuIX2RkQl0osvzqp5WCYkp7PRPJW0QjEeHqa/I5Xoh1
RYShHP2QclXrvl2LwK/JrNfAqoBFzHd6DlGWeuZrde5KBiQR2ebBoSOQHvPlasK/dOUEAPX7ZcM3
Ik2+i6MDp46vLNDsmUmP6kpMXPIuHFUHc2m96o6fbAWVRgpJa8zSsZpkzRWXslzxuW9UMC+AkG//
8FbbTLBtUWb8I3TlhB0FSteHpjEjQtOv9ycv8BkTNoYDDPBUQ4uQZd5uKczkwGJAb6m6FmbaZ4fB
h/P9dZn5xaI8IF/0RYqqlPQjcukQRvvMfQRg30WBlieljG5OyJY3nrvm73bQ+egQxPVLDngf4vmF
58Bb90ivHhWJIlG1fyIE1oEVhdKh1tVsOLynxBcdGJZCcQr+MZy2hHpPfN8qXFwtdo0TPuRbu6bK
RoCUdWwNo7aSxaMA+E2ccO33oTx0dQvfqVVgL0qyLxcmNkF6aQ1myxl0xJTdRXpmiUQfSHVoXhYz
XTsdfJ1FqjcoBH62iGA/WRYgDDHLIXhn+2vZ1wGuqm+aU4N/o7QvUxeus6JB3PzgUf+Fl8MKAUuh
2w8H+kEsNKqk2Ck9t+bpY4iqlBPToP1+H8A7ToFHoVz/TK0cKRwqnoIw2n1q3ROfMv5V0s2J2rsl
jSlnROvxr7KH4R9ifPPFqGdNWNIdk4pd819JCTvTdiRnYC/v8kGGEXFeAK7pVcM6hYtQF7M8J5Te
NpG9ZUIBQ9YpymbsaO05U3ApwCtECOI9LfDlbh5e0+yk4mLmAt9G7+VyYdep0IL0/krL3zfc+UFM
WJQXS0QncXYHoeFOuECLFh1yr/6ScnFTT1trxW/629DVPfsTtqaP99rJMmMY/+iT5oMI8gwjRUzF
SItfIwOvBvODEKhgZqKv90dFNoquyil54LWGWyxiB+20eS8q+5CgnG/+42twDx52oJi/oOKuJ9zS
V36WDgN3KPjQPmvn0XEQv4SkZO1Wz3arRE5BKXSLbDjwo+lnOgqddq4V5OnjxrsbeVIHebSlhj54
bN8S1LP7r2B3Z/82bqz0zlB7+Cgf87T96k1WUn4OuyJyMm4FNEB26mPGN74uJHA/F7nOfKhaTxTg
LOeQ/nF32FVO9SPnRlXemRTb9aA/TYC1JrdYOFGDvEobs0z/q7AZlFBafeHUbGgt1vWU+f14rYiq
TwJ+SoLM1QMZiW3Jv8uoLUGxaRZf/7dfatILV4+N9m6kiagK9M7RYNF31XDOF3RjgpIh92h/SSN/
ROmjpUPJ9w6DGuNHxdvk244cmbaftlFmLAGbsWzNWiTG+L/8i3CigWdU7QIZhDE9aGCWbK3voVyI
X1mt25m41HSJn9hPQCMVxSfy0gpWwE8aDyIUWUEdRVS1nPwsORpBDiP+7uCeqlU260Ty9s8C5FLv
+s/BgSUMOxR4lSILLH2GZvDi/FOSJBY6R1b9o6ehwscnsg5YfOq6WB1FX5uW+suFIHhzpSdbp2OZ
47EtcHZxUQGy7+5huTSEcRRnWLBeFAvUCwaXaSV9oSlxfYMW3KbeTIbflqkQVjvilRGWD6Nd28Wi
4ns+gLKJUFBQatiM+spXUWRODfIam96KztfEara71+YO/r0bkASBjoatKLR0XH0lr2Jj7yiT8Rxk
DZ92fUV+UL0jUugF4+qFSqlDUQeXeLwRfbeAkSYiTQGlepoV4eugCnJG+uWDbmT8GAilZ6Wm72dk
1amlTAKkI8ASpnH1Uw79odm63bc/ufsGzgB9O6fEo+LJ1yNcKJibbK+K7oiz6vD41xWPjmr8LcuV
sWpoFbiBsU5QUSXW0Fovr0OFjORxlo4CI1ZYdylnhQeom9IJZipkHr0/Dn3Jsff4BITwU+LoeyC5
Sk6mGvI/8jK83NcKZXwsETVqo2aCbosoXOYeGCoSjbnyGM92QX12vUtah1CU7pCBdluyvbQcQJIr
okrj/qq1vupVSzuE5IINVZ1W0btKOutDCG0bX3ZCokg/al4KeRIYNTmt87WAfBD4WVsKsoYZNEyi
MF1ICtRCvPIV56s9yN6ylHlRRayj5bFWLWCn+M5+Of4S672nhBwgQNq+xp6i/YBeMg48L/t9DQ+w
3uw5xg28xqaxyPUpPUtMZYueNAgL4FiqwPYmMMP0Lc0uRDl0PmK3xlx1PHkFa4ztCVOoGlFheP1Q
drEb7gSL+NpV/AJCfNRDmLlazoPu/UWHujBd5oy7jMUr+MWPdB2qtitqyyEiOL7GUX1NrPmfHRjk
5CXwbPhnuoLJMr9goIfDaZTkPZExtT5M1xjomCNRdYoHP0J26yiX0nKACWi5rWXGFquLB4Qxs1kJ
tOGJMifMkWWgOUMnkfZCs140Dgdogbe4YnhhSn7VBqR0COqIzknfg2D6Tf1vOZsGDnfW31v7D6ag
7DIuaezg96IYERBtytcQXwBrOz1c60tefRDCZ0fWIksCfJRoHLartQ2vP6JksQzFcwy2Dc+d4CEO
yVMFR6MzGAcxxBibNLUHhL39TACnKyx6QWWgRrCHERUkFoBDjDZsoS1oSolDG9oHHWK6+0Y1UGmj
axeESisBVGQbGYpj/CRa2fixMwuDxdL3VzVf1m6VPn0MWi6l9FRR9h71ll5/Zz3Fvog1kdqwhC1+
6wUJcqefiidT9ljMZGfX6BlHWd7jKn1ZXmKXuLXlHx6lYc1UL180+BpIwd1hD6yNVoezgzVqLMcL
U/ylzQDAAH4Kg73hbr1grTRXJO9MsxUEWVYso10YToDllAeg9JDIlL2709hVGmQldGIDmrkEcSW9
Imn6KhblWlw9jqSPGDdgB+a7Aos/ZOhC5ot2bsj3eXGnUnlxZD9nB9NwH2dkt1yB1/uzOyt973Wi
RPjGcuZp6ULTFoQ+hxqlY8fOsfACAqxz8NeDJMgMPIm1DAMozivOP5o7Q/ejZk6rul2F356sa/oY
OUzv0iB94J2VS1zildqItwP77hmdRwtzp9Y2rWEDUcT+oMcbPs1BD9Z3UEuovPGMCzV0TvDf4Qso
6DuB3VjYKPEJCW5GZoFhd5ROwiKz6zmbp2OLu7wpdKF+98j1QbxavJZnl0UP67RhrOTjMw3t+BtB
gqplzc6XnqwRQrM+1jCZYvm2CUXN4PGnN+BWohVrPvixcVmmbv4AmXIrmFugKgrT6csB6VeJQ+nl
YdQIjCouFV+FGgc/7unx4fRx0iuMDzx4pcIQui4s/GyuW620BZDB1mTIPFDuio152nakLRh21Gzl
guGHpa5qWteCcZP+NwHk3DSnUtN2FmG6NzPixuYeM1ngFqpBlTTPnEzbYAgqQU1k6HaE+DF5/uJ5
IEBNxc9LYmdXBAr7p9njqM6SWIOWpVl4KWq6b2gNXVVwJ+1huqgrSsU4MVUq1L8h4PraRLo14cpe
Om2BBLEtXgymgmR2Povl1c97sCnQ/0GGrDwWbmJzp6xPDcoynrcSvtaM6B2LiPatN4bqZmd3nSs0
+OftvfZO5Oi/UslrvOEJyd60gFhwFtGUWFSaSg4qwCi0uzCABsu4CnOZOkvQVPwf20BMCdlrA25C
xXPkBqNvEVJAE+UeIO01UTw8PJs9aqbhVoPjgjQsVOuF8yEVwYdA/XSoJJ/eDQ8/cUXh23lGG/vM
t7xe/0ybg5jNoiseh2q5G0JgjgQExMRhUOwjE/svr7/JTfxdhJRpCTnkR6ZBIODzJ/rKEizf7G68
tWy4UWDgL1XmdMC5VQZobcPs7G4hXBXR+gLKbku+A/4w3j0dhw9bzJ7TbgRxR1AS/on9THfhKcQL
j7zFe+JN/PUVosw1l51hw5OI1KjALivEQdGqPDTKeik6aQ6z6GyKU5Xg9iCJfCb+qCv1nkM8Edt+
I3QHdcWALqcA1iV1USGQWLYPtksb3VIafyXi6fHAGtoKJR5kah+hzxgrizV8yZymdsZrb6mMK7tD
4j8JgW3QeFRsX2WL1MHQtPKEtiQKESbjlq0NkIYV0IzKRLHPv78zelBPW7eEf5ka/CaqI0p6CFbZ
7RfkDorHQDG8KP6gWbbKpkkrsOPjdA5bgssLcokXm5qmAh7lpLiOIp0f/Kcc04Xr8OLcK1g4bLM/
+A2DFnTwnyKDin5kZ7xQ0AXuJz5wN/+Cd9hX0GFgpZyA0GCE1r+V1gwEZtM1eFd8POLq//qLpCXS
etR7o8q/6nfkpdmzX4LxIDWy1Nl7cz19nqOhGuuT9luLv7z87kNZge9mM3Ag18GJsk16+VEAmn77
mBlwJHK88ml7L8e+4F0X1NG51TdFA5CDTFeEDMRSJoQqJf5Po2gXBrEnOIwEgzSBE/aP+ZLlesdV
3FQlK31/FdQGoHTGdFZGfIb4/UJXiedVima6X3toEMmQsA3iwqfjcitsQz9nZAq3FXi4sIRtsAKD
tYPYgO34otKOq4gm0S0cROrTy5NaixWIR+aKNU0226uelbRvnTaI7Bm9gqSqGr7ZYdKupwN6aHG2
jGVWBC7udlNt44AIk8cz9hHHFG/11E/zVjfgItDouqcWQ5Afr1HC+j1y0q2PRpLtanD28UEOukQ4
zoVnncetPRfFOxN2bAR4AdhQBPLLfcjFaXPDcZ8aMYGzuP5435RQ+SwN+ABjno6VP2p+P9NjAVXg
0mlfZoedS5UxJPjvVNqrMf+ijmkGAXn1sANrdPd5DrtTKGyacbSKxVHdbBtWTk3GRCgFNoenOYQH
6p2hMaWtWUSlFG1PdgaC25AHXOFXP65QuIzfKfRxUNUpVcExTn3yQko8KgLI+ArzagGaR/+R7C9Y
0EOknS2q/+PvRuNHLb3Xwgp7UcJvdGIOy//mW/1szgE8LH7Y2zAsys/q/d9mGhCTvRKcjIsLTdId
ohzMsQKugQX5frzdAgA35C7AYaw6Cmfnw64BwAk3PcQDtmfMkgxjjFpos1qYdOx+84Fekyftej/+
i0I0KilLsWR3N3veyTS0n1lEfKahb1gUae/xPNPQDzag+iVaNG42qrVjz0c4x0gHUbWQIR5c2a2e
COo1wQosRvOT9LZhSWJVMRePolK6qhsMO48UAu9oEikUoyvooHZoZmUOyb4GhBmYlXIV9kKybsCp
EdmcvUsMph0bSn8EU4DYcDBoEh3x2fyAOyTSGiU3wPA2mkzaZJC5/kF09Oe5u5FLeiyeceM72FP0
w1zFdWWN04u24t6PYAcwgOJ1UN9iYXWydClWjbJmwV36DBagsOub/m5lGtBtNP7GHvzZtSUhG7BT
T0lomjTiuHrXknexnsLif5sM8Ks6cf46NO7gHUzyfDL+zta8ZdflHz/IpCMmsz9c6JWBqkZBRx7q
f2RRoBlCc4IIz9lMAYg0psBal34bSw3lXpXWr99Aw9hfI6PiKTbHd+2tWAKyEAOcDKlnZRy7utfZ
Ypemukcm+PayiJtXLhi1br+Vk1LZ+z0sClZlqSU6kUzEtIyOI/r5vJtPCMkkHXFKghexbxIdU6NF
jrYJxtC1zy6BaARBhvo+qaq2+KdxEFbaIjnfjoXbk/yJtzCIrDtr1/fnHSH/snVN06PxBIS2EmKq
jUNNlG/y7Ijb0YsoPGiJVN8sEBJV2PVMEX5koDFF9LdeCKkmky3qm7QyY7DVuvpvu68gkJkf2Gwb
04jl8JWkS5rbOa7k+M/Io4eBP5cdifyNT/eEqcYvJzl9G0h62QWR3Hfaj6nR7ArHF3rPAuTvgdu5
C97969QY7KyOrmDCfJVWoWU23DPJNCE57AfD6OP3aRVcCf514qrHNy2EUHtVK9IXaS+Tj+lH7iga
QH0THwJ8iAj6aqqt2C26ZYWcvSpRfOH1mdIClh1SXLarwDzJBQ21i2rvcwJab8oReXGof6jG1mZH
cnavBiMKreucDMqHMqAiG1V2MxcuIVLm+ssDHxhj6FTzJRPZFiAbg2S/zbPt/EXLoC1Ec385mIY4
8kNmvZR7g1QxL4O49zB1YLHMN9GSbGT629jhOZMnmQJ7xGnTOIrRC09GYdWVzPhfYRrPzPZ25do9
I1HQAiXFcJb1pCwIy883JJbPEKxE8SfdJs/SAa6TlfQdUWa1jFmw7xLhqxF9X5BBZN6HdZNVQgsg
jO7+3BvEOW40fvfQQaq0KuX4yNvqvEtcqPts2NgJPQcq3hpDao/LoeXPVOPu62uK9RcW3jxDif6v
gM7Tin6IpZt9rVD44n0tMZaTQ+b3ylrEeKu+xubDR/2IuBhaBFoa7UyFLd/+MH4yw95Zmy8a2G/3
JD5q8d19UCHO1IHHmLLlETYqO7lusRne3p2YjgkLORTmEFxjMCt7Bs+DO594pYrnqwyiyl+kZ+1I
bQTI2SYuSx/8Sk+7+ByvLSCxz4pv3T4b9OdnydA4+6FuA37YSMOxVDsIbKwuzHPH6MdUlFPKSxGE
tf9ipazD5o5r3aDD5482Eoc7irlrmozYm05SkutKKpLRoN3Ae+pY/J8TL/KnYZUzUbAbvX4Fynka
g4qFjd/FOXudLZwWrrduHw2P0o0yMGLgbdSIolACfYlytdRq380vO9mjQcMO6tENZvalRHn52k6J
lcoSYXAkc8cwCmYncZpVk+i9g5RKvy+Ymo6S03+sutUMDAqSORHl+3Bp0plUQMBKcEq9penYqq8w
ENZf23wFjQ+ryXTziyNQFsLGT5kbMPOV71SR85Lu+QX0h4p6aYFEYNpsAQZnoAcHLSvO8X/trhDi
6Y+3A/zQxOGwIM2fOulwnGJSAc4uL+ISFibeoepThorV2tL6a72hx9UA92+JmEp9xthL1zSCAUtS
zARzPbPH5EODfvEGuqwmTNid6W6qtnp1CviuFyhi3KMbSeOdhhQi82dGAsJnmxyL4R9ZIeP4HvSN
TLf9Fymjy8No8Rm20I96EDDA+WNqnQVKJxx5goeJIGtzSzQfcLzspTFUHbVCGrrnP/6xIBkYuUv/
lFkeIZI19neMr0PAI3tB1U0xGorRnhJHp1/5xrwtM8IHOEKPthb2slIrwZhtEh8nvchRrhnu4i19
4zB5oSJW4ZkhA3lZF9ixlD5phN95dp5C08Xgb3QvAm64heVuPnoNdaXyKNpYxG6hrrYxVxQh3U7f
OAHuf9Z0PL0FfZ9zAIB48KGM2SdfIsdGVnrH1KBD5+HksbF/H8ZL70d+hUAyJFC7HQ2ZoBCcbqyo
lP1IA05TcTHGX4SgADlzQGVUFHh0YfiBPTZ7pxPR0mMSogkjKGab6iyt/HtpbDu8kuRtmW8n4Peo
E3FSbHJ5sM0E85wKE+s2YqobiH23kzvCclHAml2m7C78wIOpk0h5sdi/XGbA/TvZ/fZPK5iiBDVb
SJVOOe1tWSQaZ4AqwwV4AMBjg7TTvPy1Wta1bnty7URf0PoFQDsWwUzhRdwEd+VIcFjvrjznH7+8
UKPm8xWz7ZdRpE5wQJcrEO/sWxB+WAMXnJ/eAA8vM7e8dovXBhKeNAiTmwaNFSVoHYsYLwNXUY1i
9rKnHVY9U8Dclj5VzT3GRFCicESlApGrFLALu72iffhclaIJjIt2IcMUVAHidSEA90Ab2YEaHzlV
Lyez9lOUl3uiQd+nu0vi/a7554OKhSDNaD+u3SUWsnA4+fzWkpYZrZE1BJmyKcLpHskkwhsqCenM
pziyB7GBvTh0IRTIpah9+Hc0CZ4XWAtw5jUeCwPNc6C/00PZmq64KUh8RsYxHj4Py7nR+U7A+hXI
IIkR5mtGgzY255+kHVqOK+d9jQAuqEhLAGK+AcYzBeGkoFatfLaPnuH+p2LriiIJDml/gIXD4uqW
MWD8VwBXt6QjNYqqpmS6vk/i2Yhbq7hxM5RR6KxbN7QQ9r+PiXo/QcFSRNpQuhLW3GFVpqyureJj
8DodxjUjzwUt5QpFszUjxdVSV1ery3nae0cWvqkWT839gUifGWzjpCT6pcuR9S7Qgm1bujEOySfe
dll8Ixc4wXikj/o7Ql7UPqBAFsvkQ9r+yEAvzm+qafeDKlyhUriZRNOcXw+eInEWF0nfPFh1QjqS
2wymWL4iU81E8raFCtr0khwkiC1yc+2kPZYWy5Mc98fy3VxMfg0VtC56Rn+bbeMvZkSNCDqbX2+S
drVNk6zD0zuxGxSMHSFWt1NHQ40HPYLuFSwMcHlBDW8zNzrtbZhgB5W6XFG0seuPMgYt76vD+dM0
nba8/kPuy6M957J7O9Z1rsqJQNUXt0r3jCLhRroE4vOnhYspaGKmWXGfb8Ty4Tw3RvZ7OF3xe7QD
DpLus9l8AdaOsFujPkJlvDP4zOov6oaPlzuWLQPxR14jHJxaVUJyIViK8xjBpMHDJe7yj10rO+xe
CntsjWrVtvNB7W1DwpTiNsDXmL9sq0v6/31+pcFO9vENpNOrC4zGpGkhD4tmxq/UkjVk/gyh31+E
GaYmo8+zPS782W6B9vZa4CNrCsVjnS5MZ3amhS8/MReElHD5Ah/fYBZXbKkBla9Aqh6ff1fDBGOv
OmWLwE2BjeQDVjqhxE+0wMvutNBqHggwJdYRTSy9ss+ffKTjRMbYenBN/chVIBrx/CnRCW0MEnSj
ViE24E5TXxBFXJlYRzHHgkpNB89j3jtbivOPCM8cOE35CxmLigVSNZivqaxgTyi+iWcFpLi0h1/l
cJlTW1EPfx7A5CI0dvXiKucz9oOraPBLrpIjKbrLfmvaC5XjEGw/0Kcvy6RHOratzMGbKPMDK5kb
0ZVUlzcGlPl6sVIANk679NXHBoeJZKvxwci3uD8FlWl14hDzVn7Tcp2fDMsXCJTm0H/S30bUoN+f
UR5Uh94Ck5AkC8OWWY4Gx0qpC7d9D9RFUB5zjRopWxhZVh8Oa6jbW/xVGud02K7v+nVCc3AWsydA
OQP3F81BlCSEqeEtmCP2dNQ45s8aYtnP/GYcvQ1KlzZG2fwQlM+Il5q4ln1gx8jq++cQghjc6VbB
4kWPzwCKXKrYLJkfx+72MPwc0QwU5RL6TeEwk8rZ2XcGW6zmNcGCSf+8WerFXiWDaC9KOZ0DBGqj
oDHBK6NeCwN2ITiuYru+6rF6mJaZ7H/31h2fv0BM4JIaw1vI0t4fVEMmX5t+HGhuhV7pPb/Md6oa
AB8LIDm/zrY4vaFnInl+pKSRZRmWHcjcIVlZ5aqtoi2BFmWsfwm9ZsdyWfEC/1WJxlAyNq5R+xTj
cTuVRCYnveh7bpvLwz7wJec4A4hc0ujce+jazb2wVjoyIj4SKFxvQvFDFIeAJ4zJbuGkTLJX/NC8
8+PuyjjV4vzl2ujERxavj7/us78D+oO2HiVZfnR4qmd8uPjGWu4CXukAzOzRZxlH4q9j8b6a/wc7
zj2O88vGyRzmpFL/xeIjIgvrZvsnoAC3Bcj24Av2s6YXzucrfXdLBt35T/wUvvu2FBOjIHF5ag9M
Qly2buOuHBIbPPLK7SWyzgvC4xj9jBVsGlS+XFQelAsRW01Azg/oMFqYG1AWcrfbBUoKGOr4Owtx
9KPbUvcbAr3S3jp3Nn1tXLFjGewZahXiZQth1MuyoreeNhThZBPduZ3bwFin2q+7JtF+aqLKj4it
8JMHmvxtXnMVJO9QdQsJb5qRktGWB91bZlY0ifIbtyyBizN6kasHEzmixUMJfKTftoWvoZ5mOSCd
91WmJGbL31g8/Bs1MfbrTjjG+z8zu1q+UQJtOQ8agRmZL90PzCZXGsfW2mWP4wuwe8zgMhhf/ROo
w7meJGJ/gLQRp1k468zt6DGOCAXXo5/voB5SUje+QV+JE3d99mCvpI72Fuhn1/SFemEL89M1MtMl
CL+ZSEgULcg7ThEFgNSyDt00xjl2VrWynBkPY0p06BV9ypvp3WV0E+jHHDN5kV/EWGC3N+CwhfFq
RKJ58RtRhszmWgbZo4khYEfMV2s1pCMU4jj+YYna5tv1bK5UTINYPoxmwnkemIjuIqFDJIed+5NH
a93H/gnEqxJOAiCHXnr9eJWb83t7tnAvc0dzhmsD0FLMsoCw3kelY6gVFATaEITdeje/qok1Bo+T
x/kv6wuQU2Zr5sM5T/xPUOrGdXh+sOHeVaQqnKmBJApSK0AlC15OXOziCOfem+CATeOnm00Q9d4Z
ubEgTNzNbKGCuun7vw4vSW3rGUrkj88Mia7u5sOOpQKATlIHF4BpBcMMNKS5Y1jp9Yh8w3+ZDU8q
uYLml3zJT2j/h6aRkCekT4A4zR/wvFzuonXfuBpjz4bJ/ZUWXR+mk3IOsezE91aLlofia/Wi3mRc
9qkjRy5O0drbN2uOxUtB4Go1n3ot6VCZe6ycoTXzY4ZSEmaqdSCLAvDUPWjLIHvFJNX7fqgcX/om
xZJLhSyMqqK3do8cKhGt4NVGn/0ANATkeXGMy9eEDlIXW5e8RE9iK84McXi+ctdmAFangfaJgYL4
anDPHKZTVku+W3Rk385aXmuNQZmsBTsxQMINIeCfsWHByhosKfI6I7DpGIVcoFYm6tuO2OspMbAd
Gz/xidQ2MgV89j2HFTK0cgBKiYUDa2EtESjtTKwChly1Z50XB6S7b3OT7Rbdiy5Q9ZN1lM9LRurW
koAENeTvQqq5a9vQwmgP65G4ujkGYGYpXcW9YnVBLHWRST8lnPA64u9TXY89SULv+p0HrPLG6a2M
rOiyQW2MNF6HPYjjTFUCe23GYJaCsyTUxa9uiPmpfTCND21H8bG/AOM6z80PeXrIjBU/NlIgzA0c
qWcuri38iXiETyUdS9QsTELVyalN28YkE7MLnRaQx2S48/Nvb0EIQNYjalTBljic4koIsaaOl26v
9C3ikw+ljYN5cRRBc5GkhTrayhKB36EkAORMh2e3EAMHD7SoHGvdwcUbL0ykoxJbVCGvH1qg1THR
1lFIGdrpC5GZGUZuGCNnaSUqlXETUGA+4OqkRHKqSMUvd3cXNvtkLtAb3oRo2Sjzoz4QTCxysInX
cQxIE+G1Pnec13tfGGgMZ59MG9MSqmBe2hx8iZuIYF+/5UbqWhVwAt1XowwLirmzZvXE/Uk6lPLX
zLB1QGthAipsMARIacw7cIHAPJixT05IocDSYnWTsR4fa7SZWRcu4KmVGRK5VWRS4xFshVxx4nTf
KbzDvLQIXMe2dhzvOz+LOGo4vxWb0sKL7tn6FtyDZo2DEfE4s2Hb3AfJDpOjMqJ5ubkQ2qxS6i+2
93XfzZNJVE83zm4IwHIuZFqrBPvKNIGzxTZrQHVEVijF2C4NE/d6yvysL6+Gms7Y50hokNdfzuug
/c3EaWVJPdlelTTRIxdWAh9tsadcdDnzIsf5ak1/YWhB04wvnak0A1bHSO9eF1KeVoerkEXwKLPQ
T+gPEWW2XHbLEEQQ58GGT+i2XKfSxtCu4yHVOWq48WixLEndTiYuwgCW/uTO/47MhmEAqFX5TLeU
w70RK/6rb0uBft1iIW8DIpYGNMP3d0+EeKKXjo0rjMZ9k57NKVfSFPoQTPuApivDSOTKaHnfmSxM
zpM+KkaxUYvddFfslXhwufRS+GtLjyFi8TbfO1DPd9hV1BYunB+R9JNPkyWzliWViyNe2H5met8U
H21HVmio449fvHcJNGitad6XrQphBBYBW1x8K0VAZOKFYA1SBKJqAW/obFOLELKBiAXuJZjbF4CR
E9l4hzq3O7srJKqc1C5v8RvpXCVZsHsSv0gGfdOsUnN+zrWXO8/pQ+8gSTg9MIL1MAdJ6o4qdnTC
ZwEHgp1JFfFn0H0mteH/isRsS2YSIkM75DGXloa4TGpEAwxh08loNdkJ6E91vIka7egIeXBsJQXM
onDBZxC5qykpkUrgMSwpriwWNJz0bEahGPwXRUdiiZMolMTlwaf22VRySThrX0ZTcy0jFHmO8jZ6
P+Oe45Zw7kJSrFc05bfk1Rjx2+7nrZf/7UxLiswRZ3uLE0Q6/r0CIN9BhOQiaegIuyTCkx3QHg5X
BCPqZrMU0ffvjR8SPP/0VDNa5n4+KPQVLuwmO7PCdM+Xa0/6iiQi0NSdaT+0La2NTbxCfMHNwQPy
IGaBP4zHdGFDaqnpbAE2X7MhauExvNn/zlEFuP+cSdtAXoXASvVbs3BfIs2aDnIlVN33nCcsu1/n
EHG3PWL1+E2tInvaq8E5CAWK99rGyKRQ3a79W1hPcDX7SLSsogFR4trJ3N3QyscCcvtKs4gdFDWW
sp8acvZOt/W7Of/0dFEUNl1YuUok6o/+sZrRTwZkWL3SC4GCzdsoPO4DlkFWfOQV9vHTufzRQP/+
18KRqwRSQktVC94WzBnf94Demtwuik7hF8w+1P6ff153LSB4qV2lEnBXsMzBUptkjk1dyDWtpUd5
eTRhDkwoPKyweWZSNNiWcU08qzbYmrTVWoZDvjhTzHTpXf/zx/+xMhBxFK3X9m8XF5pG7K+D3DvH
lv0wMwQmPmARR9H0rFIfMCzKm4Ip8+Mu6qOXiwthBEX/WiVkIRl0MkovGLNqfRbhttnPd9LPY6jJ
JDPwgA7dM0jkFHZC2Sh6zJAPQxeTboP3B+If366swnbMRvh4GQvlm0/Uo9SUoI1iIT71uLjrIdnS
axvGnI1e78vvdvvjt+8ngC300I+UCH98BUhZ3RNrXTWteVpUywLgydYl36V1nnJUKS2fXuhBaeQR
pvzeEu+YWHx2f48KsGu5REezjtt/qMulwi62GyA4nxU+fAGvXcKpD0qDcbZiWxKjzVhblEVbNFcb
aW9lLfpsV2bGx7m+9ZmZV9v0K8Lrftxy9JCRQbnzKLK5GgMpqLjrO2W+tVXovQpR2bQCi6vdZ+Kq
h+1RA+WAO60SkrLVcz1vuXdGBHtZa2kiIa3T/LAyqWbEj7KQTJdFzyDbRzfzDLxILe/UBJ69MRDI
ztVp2Gd5KjwHGy7rg1EhbVYpYw40kxkliR++sXcyQqAMJFFWTkLbOJrE2NYvrtBL86e/UaSd1MMX
19svj9oT+oZjoNWMdmRFI1epEb8EdkQ7kE4r0EtLyEhnMYwDXOKgPvpI1VFcNXn9X1yhWsZdciND
y7ndW7NCqu97epBOXqZnh+uBHGIWHOcNjii8Ky+p78eHUIPRqQ98mxu3KT/Yez6yrSzkjvo/PZae
69B/6WH0zOM5K01yseVSZ21SgxPk4cGvfSicuuWaYNSwApB4jBrHw7LqLsYwRs8SzFz6YzNeWsBh
XzhAceapFwCKaCKn6KbJFnyQO22W0zyzcgGTmL+6k/xijwIq4Emar6kTGwolsU/Z1EwNOXGriJWB
E36kSV0qxPuj9v4/MtNbG1g6PfEFff1KKHXcC90NBHQRQBIfSXpYSDkQz075wXg5QpZtONfjFLFQ
ST2qB5/YR4mBovoyErNOxwpTOQSEV5Cr83CsqDhfXEbhgh/v+3FueNu89W/1WvgizdyfPhzKRZJM
ba3OFA1pmbQOgTiLiFC4K4NuBIUjV9P++w0WpME8pV+iQ9ZeuQ7tDF//RxtRhJmfVOO1WHO1zFJ5
Bn+Wx4r9D5z0cPVIfwol7gwwrJCdBMwdWYAJWW4q8RdvpHtKcUpge7+OOtSH9ZVyQyXvSOx14/8W
sud1sDqGh2m15kCxcKDCkoxOmHsU2CFf0yZ8zKUpYT8zHBEvCJiGhTshd8ayB9S+P4oTKtoV1Vwn
haaqw7DRx/pAMFKdTF5xc8r6OxL4UUBVDXctN984cxD4ckESzx39l0fAEUB+jfJdFZJPFf1QFE0c
oEczxGB5YH3hGZveQ6qNhHrtednigumd6y/0l7jyF4a1uIWPdfPKpJQFmZ+iSlgGZ2gbXMmmIW0O
u4klQg71H54anXgi7ECbNCQI3xEr7+VP9biHjjxT1kXFOzTcY5Nc7hA0hwLQaYIVzDQm620cFmCn
sE+tK9C2mT81JiV65SCa5u7vATs5UhJ4lwa2PnUlEv4cxFZdRLYSjkWty7lgRdFePfSrrzVrr9J8
t0PZgBgu06Xxav3HDcBJOQpymKOHj7DWCR/EHPaw9erp5QaUL188FOR6K9Ue6cjfsWYoinVcogxI
7R/emaV6owB2PRNTaroiFHEOgjC18OLhkheGTBWz0AJPrI3b9ooJmmdC3W/kcdyEQ978u4Qz015/
mzZakUNCaDrqfAH3iYhRxIghIWakmHD4u9TZSftEA5E3IBJJy3bkRxyb/k0Qs8Slc8kWKUn/2GBU
vIRmnC9kPokFf/TbkrWxClEL1c9YsZi76VdCPz/0tr6fGDCWF2Md7r3/w9O9XR3aG5kwQoC+HWCI
Txn9oxRzMOwCA/77n8+dI2L1iCjuHxhWgW4rQIpQlnrjkqAFJDe2LIeZ3LemmQ6H1edpPMd3ugk/
kEocQ88oIMy83lydfcWWobyAFXT2xeZ8V/1dzijlmBpciytr+TMzohAKOB/cxWtOymJ/maANTEKk
q48dzDu7SKGbj0Q7bgb6+L9KzYa6491NLUHJaLzNcY30SQc8WJOW/RXThZFYfzJ6RC5Z15vpn/zB
EhfhgQbl4XXlL2K8cqCaTbPaN1/O2dM5sHqYZTpe+DqLWFyxafYCWGyJOS0oRCJFSqhC56/Zjkjt
dmC09OK3fU1CQ3PphaVMJXq4qFX/qIwh/7FiMy0HH4ZpDPbLgXS8irOB7jSJzDTQqcOVMlUlIcyr
IRf//02sVmjZaWZ5ABEPvWhwN0h8WGuCoDypkBnvnUoGG1YHqalgTx41XU4S6vz8yzDow4eHVtqI
qAPiFVnEboipxokyEUygzvHaB33r2QMs/m+xGixsIh2Q0aR8nErmv9zcFHLEoeyF3lvb0vfzfWD1
SMjqNIwez0EE5RXPoJva3NAgCJm+xd/1z3x3jyCLT1p4UDNAkrvQhQQaA9OpLgsO+EtxQQIkO+aE
eRjTn12/tN4f1q8jWLo23rqZfOI9mNa6nn/vza2USTqSpqqPXt/pNMBvCCHcZcHOyS/DAKUZohHR
9SHebnfo4Y36/Zv/5S0joX7lo2ORgz/2ojLkOFoFNa2pGTLPOsB1FyqZO2fTziSpKZLtMhAr7wQ1
lYw2eKGlxqMWZvRFemc2ybMKmPaD/pEGNcgM6Ol6wdi31FMGTQt7bhjFJGke6Isn3QszAU16YqHR
mS70De0LJ79ZFgCP7QMGEW1v4n2ezKSRq4d60GsMH2dOl3t9KUXdfBMFvX8y4jKlhYZvxo43BBvd
9CS+HZusML0UEtO9ybkGannf0HBOXWf9QhWoD7fqIw4KsdJvoLCukbfOy3HsKSJO/ae98MoQ8+iT
gORmEpI5X05O5UycU957hAu+ZyYnN2EkgCmMNF2wGdPV5IXW+Nog+CeVeVCP4iwvZik6PYQKlflB
srvkjRmQ4ZxSo8XqtGkjDklJfGsuOMkpV10feNgu/b5LM2GJQbw7N/+EXtj9tCVBolcy58hhJQA3
5DUXUTNmT8GCZP//knlewPiBTnZoRs/N9gy9hZI6WcxXrkSyOprCZqjEDNaqt7uS4meZf+je5D7B
toCW64FkgKA6E6IF/X72p0mTjwoA1uOaV90T7IeR9GgI1hLGeGSP7NhZRH6hlzY6MU5WhqaXEClB
DAR2/b9+0bgc4c7jnceoP2gg7nF7e4NKiJeTc3jjgwe9ZqcKMcAGyN3A5ckeZPqtrh0BJx54QzpY
Bxinj0V6yUkZa4aJ20VOY7xcQmToLeWEYtneNj9BsnbyEQKbW+cuu0oxET6ZEPEpm+pd9WtxcHVe
1F3NIkxnW9IuXa3mW6Zito6/fBrzbuyccEeCDnROCz75rCcixkKvvPdzm/g6gnR3l6LO6cPba/Bg
jcNcPyyyMQUmiDoYB6a8yxqx8xOCQH6rdpAPCnKP93rUK/VaAO4Ydbdqpz6xMUrUFvFqmYbRJJ/g
tDj3dWdrWM7a11JOU8FCCJUnhMm5j90Dk7Xw83IZAhPihUuZhMPUkUHl5La4TYZa7+u7WsFKm8zL
oPosmDT5Pzm8TuBhdxpeu2S2PapsQIm8K1WU0qiCWEWSJVCjLaMuuAFe/EAiDYVF3npzdF8ueVcu
00zxuLuK79DBXqLy87nkKXnnfAriUEib11ZRsF8XHTqOp1ufknEGKIC1XFXlb0LJaL2PfvddU6HM
Nn8bsI0QsyBwp/4BGi4yjzMO52YFwzsN6QjZ9CA9JM7VybpfY/p6TeqMpjnHeD3DmytLYbjP1A99
JFPg++/hhDysqbHsf0ST29/kMGne+Ed/J0wFq+IlLb4/GmjLY2PT2h9/y8tT1eGdpBTFueETpTZQ
XE56U5A3OMqQAADmsnVQ3zcQREL7AKd64j/skD1lDPfcuuic3hZAsy0yJQHQOyJ7zp1xpQOwAZLh
2YiMOJOHPZKePqXWh4QbKYQ9rtmfcC0Pcx+DWgSBVBYF9shXLojAY/KjQw8w+uOIjqyBzEcfLBkb
xL+wsM6IGyABld06+9PDG+M15ieGnxM8ggkwWp5Zy7Aq3RhjTVXOdoIDljtGRX0CPI83oAo0vxaU
E6C6P8dO6u8OLVCI7hxflJOLo4Zm9uQu7vqIl8IepTid24x0JFNpaJz/lBwZmdLD8w94Odzcub5s
0zf2UM5e4dVvv1YlTJjg5C/rt6q1U437FHBjH6Pk78Uv2NUf/FdFURl1KDh/RlFWQBLgEgn9q1JH
UeVs5rX9FzdGQmYqjTSIQy1ooDLLk6SDd68MCu8YMGDT2rx7bYGgyy93NdKrMBeYw3lLS/y/P8os
VtyD5V/z8BqLZRTzOjRB9tIQ81pf9l9hecylJPpB1KacKkImnSCDw+enSQgnfmrhVcDa6+LR1Orz
tKZ2w6bAkWdI/qgkryXcXE4lEINzPASoNyfY722rjI/Sk61YTB5mauTPeTneMb06y0Jkd05byUaz
gzw/6YN57EQ0DPYwUhkLVhFi1RBLISUlrToVCJpn5oTretH6MMk1v/aT0l9HYdjazWpmV1zGYq18
wOVXzHNVGre5y6cwyqC9GlBGNTEDGM5Ltxz5UFfSR7q7zQcfFqKzxI+5wz6h/z68fdlxu01nFjIU
cH++1HTReviORpL98agx3cv0mnlFgr688zcWp0xJizOb5NmffSoSI0BNJQxNdMId+frnSfW8+9Kf
hTAm/VLsPCW97GVzYQqAunRfNQD/5wzeSlwd5LbVRH6yfq6kLhjvwIZpx3RJMuuZuCOj1chCvmd3
1X0yfQaFNwInCpjEEhQsBN0+0ny295+rU+xteDH+GkI9y4zcIe9xpaDkX8+PRsoKLWZF3E0aAOjp
dxZT2l7pbhbMZAzn71cTNEmU0C1SDouv6uU0/QJuJ9MWOg6ArMv6eZhI1zI9utCD6rEK96u9Eo8D
qo1wFhvrJX6S+0Jlgu7pQLY4HzJIiveFqBrjPa5YemdX52+dMoqsZj+Up2MKs7MMljMGwZrSHbGn
gLXbroxMFECEKim4WnnlScTkON8J1ftgq6IeHI48nJp51yV5ak8D+br3BrTTx7IIdcEi1gUnlB5D
99oOzmyE14ChrkzkFCJH9rrHycwjIfk3ZzPaC1tv7UB4io9UjpZu+ouS1N4Zze4asJY/tMaw/Nll
QGsEfwHzvehTfV7gouOAcDq+M408i+6RrzeGxvUwUYe0+Ye9Y77DQGxS27CHrap66uWgTfAMMfQJ
bfaRs31zcrlxf+vU8Xsm8vsKHA95cvWelVFhRyC9JD8wu4eD88pDN6VllLrPTLKRGvAj/5WFtVkA
XJWvK8TJ5W8G37NFu6xJamo1rOc29WQCOWkGfs7tA4B0aY9SvAxupz3ORefge0UmxuLuNvAvFHbm
vMDCy9DLgarmHnJMkKFe0xQK9OJDHtgEUUITzSECpulgfAupfnAcdjfI6nJCRXDqxnvVxi9LNwLP
uEJZ1F6TbwFu6QTOy7E6NbN5E8CADWcYaOuVk/x5VcWXz5fXNiNY/tJKOxVSqyVeXJ6wJA1sXTIU
sO7FqLSpzEGaNXPZDdRtWZZ44T5mq+G6CbLvLOB7HNYlnGCQNIKaxdeDbj0i2tbszGoIDNiLEnrH
SdsSphxOhOAmVcoZHyuU2au3+Ah4Dmk3DxXO6Pb0ZiZSF8tE8GHmDQl6xUMj5Ovk587hAVXOK0u3
90Pr1E4Vm9DIk6ms8q2oiE1nlok0hUHP/6wpfSZxU1r6jXmTtTT9BWVe3I86UJ/bDPK4L0iXyhDY
qmoM4MyxEW+JBLijqsi+nBBKn18vrnm2OIsCuBYszqj688LfYaSrnSaPOs6gL/aE8KW4VaUj2I+I
Fnqc82W5q2UNPAptu4RZpZ2CFqHx8Cy9id4da+V83u8hhCKwl3G6oDB+bS53MCGjSF4WDGgmyDqh
UHDEY1Rfa7DAfsERRPmDptNOvXaMTYuklx+YLsI+LXzLiIyRIhDoIz1HWvLGw1fwm1jZbB8VtFfV
7xs12fUQkxZvhiKiYmH6xs8ijDGl5AgEgM6IY8qeWAL84U3cPfEgFoZQVOBwDwC9xd3Cuf54+DYt
KFeLJ5NL3tS8J0uu6LcaYkxKs9hyl5H27FedaOXQgTZFAiJ9Sdeo6aPC9KuhL2O3/ye+XqWLS0J0
x2wEufgmZJW5fGCq9k/FnbAMptNhfSud3k9QOcztAmh3EW93N14VMoJTFUW2G/4Fzc2F9fTi6wfM
CYC9hd1o+8bEky+RvBlYJN0HprzPi4pPFVjob1HQC4TQuc+Pmj3meL/fWCZkQU0vO7buHn1n6yK5
eEXWxFBcJRYZBucYiwnW85e75NkO/fo5sx5XCQSC953UPuajWV1yCV1LyyhPbH/rBuxTeCGI0e2b
pyTAOcNgN8CBuUNoSGumGRd7DJA3iEaFfJI9kEvtelvUSoFIWO0YWcs7uLHxYdoujAvJb81SMxU5
7H2JYiVSyGREzIEvBr8ojLw+C02O87+J0qyGgWhllzFMaTn0RS+y+9uHPia6P57X38MtcNWMQmO0
HFyEwOrHnlrB36yIpAFLjKC2t58r2Y3cblUIRh3+6x12Z7YPOyB82XQSun1EF0Tf0Iq8e3XOOunD
Xknsl2WBPkXvvOB9gci5fnPhDnkFDa4NfD6fQ1faC/vNMyvyUz5CIQxuxK7txTmSlRsWWGyAZNvT
D55T5yodlXRgcFEdrX0BGhv8NhqLxM3b13anYG+zql9/Lvaew4LtTrEHkIrHXM9lrz6jfjiifFgL
xnfAnMDNVFvInCCECxZCpVmaqu08jMfXKH2O3PFH03tl9J++5rFmP0+U2HdjYtTuGWP2dyQxBSCR
taEB7eKxltwNXu8CCMKvFtGAQJ5Ahi+Uwja1IDd82+SiUvjIAeyLUGD+3u5PNUBVAHUb2BWzfJIf
XuXZsgzdmpZEuyEh9/m0PD25fBHIaReQGnenHS0oVkeI7DjN1HrG5UnjPygTswgMKTfGpF4w65IO
Jd5kmZ6YRcrSoYXWEuYqX1TfoZ3STIukYW2tTy/Ur8NTc/VGLGhGYfUD+2rc3WSr7EvdSXd7LaR7
rtDy+7d6fwv+rYH9d6Xk/6sWCdnZiZBd5v7xbQb8Q1gCeQfti4ekNNoLmdOL1RU4ZDe786vtWtak
hzse4EUfCZ25azfnyWN9wUGpTCgFR0WOdFxZBmOvsUHIbqPCj8diaEqHNLDPFKp+shmQkjihb7lZ
AftaPHYtPccCX4D+FiYCcq9zWo+k1vYo4kVGROF5VIgpzSQtRcmdJ67OjmoEbD9JvKLvvpONKrkj
GNNCdJ8IvK7SxDqTdVvBuUDtKMVMq5EO28vzh1q2VKkr9KV72wAEJ0V3sZ7OPbbPUnxhR2rgKWxQ
i4EmDGqxos54Zn7DAcEDoNeWXS2QHjAcc7Xtj643G57KORy0KgoG0ph1IoQ/zXkMU/w9PfoY3TsW
HrwrYjcUBx2h5/XzEzTGl9NJCOvtnhzfzYxfFRmXB7bFp0lY0sXbyTwDeOp22qlaZB55Me5ZBU2I
nCQI7UPVntC7VKuvz9igqucvibV9iywkpLXtz4mOLUlRthwTb+48MvQmWDcoRPfeVYGS1BCF6z/I
/gemF412pRbQxMxfb7Lr97Q52nkLb8evBctIjpvoMRZ1/u5xES5oIn19LwRI4DHeiEmWmebvynPa
q8R+Z9835cQcz65N++YUxZnAy8XI3u+z9cq89tU+2oWO0kJcVFzuIT8piPQG774Y32rJkwyqnXX6
yYTuFqp4yiRYrPyo17+gUwuJn5sK6locJfuvItdAr5anvvZBi2KdLBZQ4fU1BhHlJl7LWeXXNZQm
PKS2aSJDqmLQBSTDgWZuAthpTFKScQHyHXrQuRRNGIFlQYFpzm6GmEcxXaaVmbSo5uJKcpRJOAmt
Exmc1R+zBDRK0l69GTlMqW2HCX4yWRTNco4o2c8rJ3dNCrgENe9/on1t8ns/Z26ndbHJvfE/CaBH
uhrixJhkm5NKQ/FSn4YU43XuPNlXhKsZf74BEOVvmYab9JVQgf0XWRKO4d707M0g9Qw5iaSU2r8l
gijpb7/WJePEPmfH1g6tmzvTRkxZ61TJLhzo+oQxO55kNqy/+74Uf059nL//viM0nRVxA6BL8VV4
PhsF/qM6wTFyPhY2M25hDL4YdVSJEmzg4wHch22tQy7GAE0+xTq0sffgYuUG34FZsVTbMZwednoO
Q3O4rEtOZKqX2sg+Y5Cl6xl+DNr1sfGpA+jKo39kDjxu8Uo3E6fP8YVx/tR+7LUMsxuU5zVmGcZ/
hYC5EZ+/JhB3cnA/PBLOBXsijK2xJBagsix8IxHrahwTuv4fGXaMVOCW1hSKPlLhbWwBOUbUR7mC
IK0BDRQ8HFJOBlITP4DK2ns7YXQGkRBnFsu08GcTWDi0zwD+K+UoQGuf1OA8qu0qYe+hpqzyKtEg
blTupHs359aBmL8x2d5n2Eu3XT6xsLCA0ZEJKNoMW7sA5z93pztty3P7J2NY+smFrHH87MzXCHyh
/29/Mwe6DZL+rvpaXFgo+8re/D15b0UD6ZwH7JAMaoipiCuQ17CP89zdQ3hgaeYVQlVHugATVupt
0zdnyUHMTMMrgmZwpeRRek4EvH1vQKZoWUzj2lT7oDs56mY/Wp5C2haxgaV2OCW3rs/116VFDWeP
5pN+JUnOCc3uRRtN/31pfGM9uw6cFhnhREjl3tB/3Nz4KcwQDjAwZdf9mfgEFX8FKWiZsL/D9QQ1
4l8Jd7Yteioqw622HNJBF8byx+3FucKxSsdOnLd/cPGOdVUi/6KkzWnSkjUaeay2OyNA/YvNBym2
7ELOtMq0QC51DEp+XhfIxkj7nOXQBb8XZcwcjqKvC13cKaPf1Jxl28rLUP1hcwD5V0v8e9IXCQug
XmqfrGPqCwdp10yTF2E2BEAX+1cMwGH8A7uMwdeGpTIyORoJqA+97niracmB3XwzCSlTAhYXyVSz
JhKAFErXWORK/wYvIuyrFFTLbSei5szpbg4Uw73HcIUkAIy7q5Qu6IXTZDrkhqu4/8nZQU8BOhsN
5w7K2DW4BazFseTDs6pKKmtEuZT72mZ9BTWRtB7x2NSqjcXltzlQpLWkD3pBT/NLLwh8w/xQJGEn
C/iJMdxFa9BdqHiTePx8rqBYNz4p3ynM1Z1NHd66LqFwWLsVCj00P+T9j+RxZcGDJtL938oRXzCH
bgxYIxJuo34NH6dz26OQpzwcEfbiYVFZ6trB33xEWBljpM2kySJQiU9UuDiPI2YIxbBETk8sE39h
rm7YB6Ssyf43JXXsluKm0TKNo4WjbW68Hc9/O2Zp3fia4XtssTaRRhKan/U3dwN5Hfd2Djkkxs1D
o2yJKh1Eem0fT9d1JtpiXbO1Bmld0jmRmceOkJDit7cd7qALyRJHe/OEOQPiZFZuVYGloN7rB3MQ
/kg26rXNorHLVB4sA8jrbCrceQXsnBsfSSqc+Pt9JX8WdVnLemne7bE1fQuG2J+jQSQJ6QGR7oXq
Y8ZqALdahruQLGbfkWXjEx4PO1S+2KrloMidXnIGTKae3IBPlXWsR6I0igdK87FGDRfQUdCip7i8
oGgHqNCCnQ1FmMgrK5aUXSQimG2/r+ZYLq8vNXXL3fOXIXQ6hKiSE0cdjrozu8gBJ5uO6Cf22VWC
xrA94Jz74cerfutRUtkUdQhRZ+60L666w2rwhsIJGIbJD2lfCWCzxaOlSZOIVXWFQ97F4/88s0Hr
tBBS+n/vB6utjmbjaIdazIEtCMsVzfjjPBvSy7d1/Fw3kTn0QTfSzRTiUucR1EG3lIkWJgPT3qwT
PNes92LN7stgeFgYwIpk58t5cbxPRinZe+n8QKIwUJvzgJM6tiOOL1sZ2lLZ7IZB91iX8OBC5ZQH
F3ZNv5q0394s2eNC+C3CHHxd6ArzWHej1/UYG0dTm62SQdh4YjWlXOfM+HPvdjmp91hGiv2OWF4y
tKbBbQN1EWZKOA82zE/yx70fIW3zbzkeCzqFBjNw2lhqkBYw754GiVVt5DjzVzDKka7U7a25ZrHj
zn0NMYwfn5TLmA0frEYFnLzgx90mx8Un2EVR1F9TZNFOgLK5aNWzZB76Te1k5bLWSl3xb8KlrO/4
hHYs0ycnalgw29UiDibuFM3KzNfy+1MMJ/brGOHQpMFQ2AR4YY5Ztt80sgy+nH8bg5QJzgRVPXV/
HZ8mk9Snz91/ckgaHOxpY8ZWLsWJyLVm2OzKYR2OYqKveLI1jYDeJ5uyX6OXBQOiJ4doENOcdWPk
b2tvLdXavAsqFTT7OcgpZ8qT3VMScQ2w82HFEHNSz1FdrSrqMRoDtVNMeecfOhpSX2i8vx6AN8Nd
cHZ9dfe+BLExycaYFwM/ylXgkGYrb58dM44HuBVomtmmvAmT5sipzFtN6mdEHAeAmDu9HVB13t1Q
4XjZUtt6oihlMKKegWJgUUcC+FMnSntz+nF1HXx9B8AwjRfgy7lJltH/7SgBku/HW3V6LWGD9wP+
jz6IDAcO8KjPWi3VmnOiLKAco+t1S19w/aVv7YMDyy0a/fqK707RSnFAHxdsa1m8Kmqy7379G+7o
+M2BxrnuDm3xveLdSH6hFh6JT+cNI720YTbEdXVBxBVdmb/9+7cGwiYujvsb74K112H7va3AMup3
vCEOtt/WS1g6iZqYhNmnbtL2ZyX6avZHz0Gqw1qtxDXHOSzXHVxvasMPphYRxs7slmWXRsSt15bZ
b12aUbufBB4zsTzg8Stuq+E8krrgIUT61dms6hlK9syk3l2WMqUsbMOo9vTjUhWhEzdEJY6fPcTN
+bA6x0Dg48S4/nkRB8yQVclXCZavCE2vvVMAZB4vJScJ0mBTRcXxFwAy3AqY6pLrMAS+LFKrr9eJ
8QiZDKoH+ecijiWu4HCxTVvL8N5AONfyxN/dPU1j8j2c/Ohn3D1vlsIIPmGC5C61bW76wMh35utP
kbv6VFeAXKRYogguvVIwPu0JS3RVwV/8bhr4OCZm/Caz3D9xQdU9Yt3BpHyMe84WD7cbVb/1kcaO
LlnusnDm2xQJEj9V5FLWhmIk+/jXBl5xSs4CSXTbt/vVyhFMibhrXxGtEkMgopu6QlQWBcbEQICH
8BvjnAt2L3x/jgvqaSuM2g1CqdNXCzquTC+8xoSd5Sh8lrtOAZaVt+XX6/t8tuXjbfHnrIKLec1d
zBQamQJoOl2FWf99yqKfS7sGEbjN0SljYNy1neQxhWUk9CgLzrvkNFRiRGmTYkckPU2Z70ENR5I4
FFygFf+aiXsBNIj4XmvU7w72Orqw+vVt1aGa8+gqK+zHBSN40S9wKjO1KzGrL7iDNX+L2sHOpyjl
EesWRDCIYN33XCyPhpTzgS6GhdA60LA5bRGeISlvKwT8ltyQpkMAxnuiQGpyBvmtDIpQvwHrRMSR
2bnj0ckGeYvJGCg7vFCVSfH1nz21ww/8+VbhCVDNMoWMHDcLNohRBAML2l837PpuhGIU2WbiYlJd
x1oydkMv6BtDX5B52fPqruFjoZtN/MKOop6pKfoEowrfGInOFGDBkTRxoJ2mG560fnjGa0LRZTvj
bZenqGLKDzGGVgm61+5k7vh3SWd3FJL9yodovzhTAKAC8frOhuhsjlQyI8d+r+/ebqJ/0v5NQUJu
bXTHiYRZyC8nH8KtHDIu8r6tklZzR4IYtviQ26HLRXuTW5IU4c6tlICzQtTSbc211LGDAxFw9ayd
/4BKGPIX6CyED9oUrKa0QgCOjsH5xaaqxN3i6rsAH5uxh06yVGJO74d0GJEZC0Lkf8LVgFyYbCKh
hIqodDhgyXJdAkOxVtwoWbRXLjtEVfUQGzvZm+juM4Hh4HSH3kH+rtZGJNqqFERdluoFRKURzzAe
5nv6UgOLcr5EtgSfOJsz8Q1AR/2sRVCFWGx4OPhIqN5BL3s5SwmNnQIq55oIhVnITdsZFC/m+7sQ
k6xBoKIbb61zdxl9PtCwgLkTn3BSLXegVt/f8RMH6RdfYC75Z74/AzBq4okF/YocOzltyO7kAp6B
buR5VHthBdv1EoRvkoDA+9zanWhfsifncIdCUE5jXEa3a6F4ealyKB2uf5oK/chWWgmsFOX8Zuln
ZhAia+IIAn8NoP6GJukcX1tuwkl9bMl/sD5Oqg+3Xc+jlYC+uQm7Zv6yODjIwDXQ/kaO62ZkXsjI
iluiZj8vZhZwIA4oriL1uAQk559luWrvX2jRU8g5zRi8zwrWCEo7ZuQs0HTevQlMH3Sou0Ve+Yh3
n2FthQkivP6bgP5wmkf3rqgQimRm5ZtW0VwY72odM3TOWj0bdHuyOvaU5+veNx5HfUJIQ2Kxa7k5
Rkcc+AsCWA4xTqdQdXrUILDPYmxt4iN4yBTbWGsMreKtdalrHmFYhmcuvHxtDTGCOB401xRwKRFj
wktcKsJD4tcuPmz0BpfCDBFwhVpXBCMPjf4WnbMyq+ib5j2vXkSlRmzd9lSCZ+tqzZwuGX6ojgcR
YJBEZksGbQ0epG8R7TIfJW2A3nciqoAUTf0zWxg+pW2ifpw+jCSo5SHGoSecrn5Uk2clWxfkvhju
WFSLXHycYsKLI9S0iYSmOdDDZJIwvVz2cME1ccuGc0cdVWVtpqADll+15c0UlZMLOZG6O9CkCNwa
vilZw9W9wUVsNuuzmvrqrZJmt2NCGgU5MiDc3ErJfNqVFVVc9wHWlf+qrYCBbCtW6mc0aSCbtuhQ
fAbIFayss9NayWEnLPTjbh63laL+uofvoDkqDyirmE9NP0XzEx92b66QROkhT4UwFNRbx7PrYOJK
a906Ac+22RymyUbd3Xm21m05l9SWshpKPufodYq89pWNpM9r54RjCWr76qC+vB4XSn1ixjuEPJS0
brTSYzS0PeKu5clqhDLw8Pdrbwym3kB/EZHg+sHuDOgAduLSDXDGogWU1cHYcVctYKxAs6++4sLL
SQxaw4GLtGq7ivd9ETPdKoqONmrS++aHL6EQze3yuDgzyMiMOpEQSeze7aiVqN1AFu87IjZuZdZb
7wzyXzzk+/o2UrbuomY8zQMVsojlcxeUvrG8o9h5woDP4yrF++jXtMgb7UFs9v3pl30nwOSCRxm6
RDGgiKZUpbDRx5cSRml46ZXPwlplmk4JVh37e3SQ/5MK7Yoh4dEgxytpbh8/wE+37x8gY31MfvS0
hnPg0fzEQcVhE9S8wxX6M/9LsMWHkkE5rHO/w6VtGF0kh3e+xVp4mOGXAV7fHki32w16E86PeMkk
Gwsz0cPf1JckzFO/GGcpJdj6Ewr0QJ0GiW0OQDk4hTWOX6CObs3dpnb7dDa9+1dGAABvDi/feHpJ
H+EjqNMfTrBdaL/gK7gwIMWKQ2Zn8ezgdxsUR7PbNCcNipoo12nkLphmg1bjqHwguwlspU4uaN/Q
t18w/wuwT62fevMUsVr67RaFDPomdEibIZ68g8FLMKfD/nN1vxv9/Vs33ily9p63RcmQ3BJOPEJD
x6CXx8jvj815vEpNu72/wISXfU4GBAQCAzRq5nWfgZNqg567CYd94x2Y+84XbYu8CjmspCJ/kHsy
PBoOCzlHZb6cNIEJvDlmVRw25GYLMBqn1UQyrYTnKKQPkQyNrtdP9gogN0zl51d7ZfNTKYDiH7en
l60VQS8tm6iYShJ48F9ku8TxDvg+1RY1a4jncg8BK7BQcB3lRsjkqEitRraAV50jWHJ3hr6upJvU
ROQdaEmDYPSF7+On9cvRQ71QDeU9Je5z3N6EBKumceoDMqw9FW1L73SK34+KMa8S+kGkXwJjx+RI
jnMXZDVBAWhWjxw8m99Tsb5+xmC2/KPy6TU3wIHBdEav1Eqxwdwmx6cvjueBLDuWv0/Uukxjt/Fe
XFlpDbvk6gdUDfyuArCj7RqlI/wS3OsGvwsvZi165mK8IJngzTJEkL4j+mMiekKm3WhM7MfCbUv7
1ZLbz7JLYIxIexL8mcHnAce/T2DsHVXPdP0RkAbsUyioPmCiUstPg1MsF3pLwH76jj3Gdv4PeVfR
hTT40UChlysnxdO2joWobk1bTOrsXfiMRx3NRIGJu55s3aYtIa7oAa4LcmeYyN/767dTGE0HGj5J
r4Z3sg79kaDkvgK+vkTVDkG4imxuwcD1yRn0fLbWCM2P0FbxNWJId3VZQal0Al1BOWXvmdyt4QaJ
+swL5vRAyjkOdNtLXLysnZ5o37Dem9mTouLdgtEkupu6ExmlMxHBI3AM5wcoYMpW9FtNKnwhqoRt
wNBswd/UBtBSirksvN4X2Fsn8DOXpci0EYkIGrft+i43aKPL9mW+N/FCMY72irua2bsncY+pq0zh
kW8e1gcAjWQKNbpcqPnJFB533A2rm/g1ZjIj7KxRsXlrZmVV2YqmQAh6BxYDzZHBlsefJLvdjgDY
zsPQon6gnb2BetrzjQ9IeH68L26+qso8uB2mrYqXy0SbThfcqMdN7jvrTTZutVfFLn/Fg35eE1Tf
eIxBU80Eurue5BEu0yWMnuGgj51S/5WM6Sgm8s6/rLX48o4eNARRWSFCNlNt1tZXTpJOiWWeKMvU
k2bhDaNuQQOVRp8ePNdgTeDwZmpH3p8scU7bxCVD4D0VPDS6cks1lbjesk28M0GwwOq2dyKEpuTN
h8yA/lNhnbJEkSuagLHAwQl3qWfg4cc9Zbzfr29NJUiE6rEx6up/RudCC7s3G70ICqYFuju1TXeK
0rZZG7pUb1aFzv1Hjm4+JR8QHBLXm8bAzorieWAd22Rir1dlx6S/WduJpq86XAth/7V44T4AnECq
qmSnhyHAhDlFVUZ/C1wIf+mfrdA4VavxZr1S0qmX5+Lm5CoI/wC6H7PNUGkA2EdqHStgM8dVU7oo
Cum1Tmj83RDVrhzE6OkLGzUAYbsF1/ZnYnY9PqCP59BBb+P2mYhL6hKCHSoVpMcYdV0jAMx+PAC5
6bXq+PctmnOhhq96YI7Hl0/Ydak4fhze36w4G6UP36Mcxx1QhAqTAWccjX5Z0pXyHK3Ns+nNDtpZ
nu4gf2Fjt4AXCBgMhk+wUy68OIffDOsXI1MPHq9loZHH6mxiubAtqmHRy+g6ykU0B9ZDicd1TRWL
cTEnB+Pv8fLvQGjFZ8qy10PEokD4h2Cw1Jq/ufga3JCvVHEePTMNTkvh7dNrhiYXO+ocfGSmswp0
Eqkq4OzqQbd+2G0c0lRm2ToOwn2orxLY2YuUJxmpQadlsxxqXUBKc7RjYm5qo4fDdmMUC00h0Sme
FRcTKMO3oxUxS2XbrapjZs+SgWRUf3UYnM22tonDWUUcQJKEjKvuKeksHZF449ru54KQprbUz8sU
MYOmAorgS8FlCT2Re4GK9UjjYbobEemlHONfGYIc/omdCsEJ/6XzwPwQOOFq3F//7mQpvHC98lQQ
C7FaJ9wZZko0YlcwTn+pe5K013D20dniNXz4qyQKuMXajfeX9/ocGRetLydxVTABCfVsTVTZYh75
PiFpNA0wrL6OvdTxwXJ1S32yvkhMRZx2aoYATfXs0AEaT6jIGPe/pHWuz747UHG/iZU7TcRM9CYx
vTZ7L+0MvFAHdzbsMINaNPiI7TkpqRlFsITcgNYWvKDVO7eYMVduyvk204QsBy8OW6GZM1xyLw5u
jCZ+8+kbl9tXhTKCAJ9clb9dmjtcQQL0Ae/HfP2znas1LhzLfUSsnx2yHYiWnVerINUtsGPn7sUL
DpZVtw1a1sFV5dLO5vK01hPpKukf+igwVfqdBSesi1tbCc6oNuUX5Vm5jQzL/If4yhHRpi3GHz14
xpYL3AyyaZFt2Vv7UvqgnH/vkL37/tzQZ+61JPspZh6fBjWKWKdQFdOn5mpwKewIpTYBrqNSWP5l
QN61Ub+Uqu6o1WisfFWRgVLft+bRzEMrsUk5aZoKci+3j5AgfuS7HhjXUSOrPwKgvDST56DGVnle
gLoGyhOTDJY9VRZibqvrwMGY2P97Kw/hxNZ9eMD+HoWieBOSG3kGWC6zhnWCK6D3WLJqmSMWr5Cx
FskYCFrLmI/LaRYxq3C+evNs3GGNx7bShEVCHTn5SV2+7xQjBUVlPiHqbiilLzbsoaJqdYXdraro
EeH2MK2kcXK9F+Xaz38N7pFOi+PrNjb6Cs0+LP9URgGNlGoO7uVF3ZwobC89lMI+xaF2C4lPfLq2
27cWau2RA+tOp2cbgEtgZFZVvAScb1IfH3UxJ4tEGB3A5vsQHiNVu7PuTnKR+qyM4tLuIzWozg4P
Xinxfnbw0rBFHLFKk85/zcWkfUBkd3ajEFcUyqWMFP9ixMbStovPMcGbf5JEovmBDHHnmoWbYuKI
eEohc3pnejtvs3fEo4m1BguitwepiG1cWanftAVSnk0j0LucFab2TqZCuqE/igg16orrSRm0QXFc
ncteOVrNhfevUk14vLtmoQ1HFBWTV2iS526KxVYpnuIbMlLeFbecnTh3kr9U7RweAPuZL3Z+HDb7
H/JB/USUjkIcA/I4rvxqQnZnb2rDkZQlYkKPVwJGQC55vDGOMkGfGwrzmLVcehllPyHwa3TMwmFo
LSzUNVOjFM5EDMJMPFzsB4ljjjmiQJkXt9ScEdFZYPlGyb0rw7ZvWFn8u0LVmH45J0HWeJGOhVHH
ss5W7GqsUfR/pUrYEgrYOdhi7p1OYY55wSzR5C3L9XmnqzEFL+g9Ur+++kdV9GdXp4TbetwHq+T1
nxQgnXznKlYHa2X//KE8G8CgNuOs77cg37XCy2EmKElUvohBWoggYtYV2one3UBMqYb6k+8wCPxL
if/1UD1oU1Ut61Y9QxL3EDWNVsTafVuHUha9kycuXeFU2ytB6qrc7oE5tgjUjTft8G3fH2xiqyhR
U2yU95rEAoMZvMqGkF1/f/jriAcPymCcbcZKuP5fmAytsf/uKpjaGO4+n+CbxZlnls3XLMpONFOl
Uz3Hx5IdLVmrbw4MCxBi38KJwWwOUnJnNikl7zfyt3zCPszMugFNJQ38n7OiQrUm6QwrtrAr1dvO
KXpsmPmx1O7v363nkIGHTKmsBB7ybiIKQpMh46KYCziS9HHFA58n7o+hSjL+DJ7MrWQMM6EjTQSZ
urU1Y/6VFUKuqbpVoaIULeHv9FVz/i50wcLwrQMOKFkTcgXkV1GQHZyLF/qwH2H166DP0LipKQCe
ADzILnlTC0GP/RxhxMXBC5ljzTL3nm7n01WRpun46iooETZjeubwR2WZfCxQK1kaIqhsfRUOa1Vp
j63FQarIHelCRmVU4Y9Onbmi+ssf8Uk97U/6uFZ+g06CUpg7nQHawBM8eiw/FDG7t/YgS3uRETTU
YsH1QfrD5L0DzkhcCVsMfswmqg4RBPDcVCgBFtmekBfKoTMxxCM69b8uH2nTxfCDMFY5AaHm9Q42
LEHGxreXYOvVuCTGTfYTywxALCR+4mxgADsqdKcdgXsv2ZK9dggmoXVirgz3WBhf8lNC4bKhehzD
FvhBm3ioVzfbj6ZkmRy1IAzorao5DWfwYcyEVvkpWcHOutbQLsMpCXskMOQJ50RfWi89iMy4U3SE
u8MujHLzTf1slhN01BXwVZbq7SGzo0Gft9d7TVmHff4EZvrOtaWJtZyn84dg8ey614fLeE92LWS7
LeUGgiV/76l/Q4Q/PO9QKwLiE9kDbdOcWiYSEkp6W1I2kk0V3kiENqXlYIfyzXOEK4/L2GDQrmuk
ZOmHypTxToaqR/W9HR2bRz+L62zrekUn4ROHjBggXd3B88xUT1Czwi3HVwmt5xlcSUGlirwePqBV
Mov4XhaoA8YKqw7wWeVoqu5ENDu15+kgdteJcf7fOuIuKhMfOgUMD7zvIGPnD3d7JwlOICkQUygh
OL8yFWrA3FtSwKOWU/laQmTgS4nCB5QDgTiFlnvvXrEaSTl/Q17A9Yk+dXjLW6hMjJDc2dP1r8bs
1hu4ce72VO5GC44VOCUd9PkLFeKDIBCSUnY2XJj9kVQRu9U9aUhNQ/VpRsaXoZKotQaF0GqQNhTk
F800hpOgM+nnO1lD+wT4612Ugnc1hOF8Gf/zeaQcZukhgu8HkzXOi3sSST5SqPxaaKfsPjR937ch
skY38VIl+LJGKuWCwDIUuiaCTkUOYWaSH76gM1Knrh1DXxw8QmWErmcPDwxOPBXaIT2OA/s+FmJx
Vgug2DTQSvU6fv5uOKbhVMc1arf2ZsW83lBpE4vpZIYDa7YqlgzLzUF7CQJ0BetjKl2JQ5+FHr1d
58XGFO9Tb0kiTQUJAO22gVYE6E10AOmqImfwot7NWXP58tUr1LRWacnEUXJbrf3PWDvBQ4DFuOsy
EQw8JqgWZU3bFyAAWfuFQpnsUzBxWQY7JpItRJWAW2DFGCOKOkdsP3uu0eHU6jQlFqKFGbxn6t/h
OkwrQWvxRbW6BkCOcPbcnf5j1277H7j+owYzZgrwv22R8C/f6Z9fUZxUaeUXC+OI0mPP6tBGbF/V
bJvWwQnExP/I7SgUnNBoGXVY0RNS3Q4XqDk8LkwdnVvLXNORqEfElB21/fxCIy6jnb/cpuIgr6gf
OePDdh9tLvHuds/CexWmdda9/aWBBiLSVclv/K2gW4GSQQOnsfHt5uOTAH/G6as0NRx9aEGvoauO
1RVR9s4a+ex2q1QPPDcRhRRzHu9B+4Ap/D5K7Oi1IW68sd01t+8nwrx2exUTv53Lr22EGsit56Vg
MaNopgR2H21wSPNAJQoleJ5eL0wsKMXHko9J2N+mXO0y0+0mjxy9DyKl9QbOnYpEymBWmfrvCPLB
n6bM/MA4CX/swLwi2NponCrJ8eAPZoCueeROZFBlz3uLJ31e/iE3xUO6J7nukJbBoSMoLnYfLPEV
MBht+aSznoiIUnE3tcQM7H8PPyvFhxRwi+/3Zwu5WjPfyWlVzJAwX16qsI0wiOA6td7gh+WcBkwH
PNOd3BH8xCc4MSRBaBA9Ifv6fdYWkRQ3KNlDp9rqdWYXMcfcb1blozRybzMXE9gXAYQ2l9daI4xW
zWouqp3WP+6b3Jb36DWjRGLItnMliJton8QvTgRN+yoJeqFsIs+2p+NP0ndNFMh43JE/M8twnDRn
1dH8deeLWTdINf7ImurXFYTmifOw5k/KgfOVCbWCXVmtr1nLZ7uvI1SpesLdpsRqBlpaSDi1aIBE
MQUxMvYNe79LGadOJoZe8oZfdKPtLWkVZeMRBy5p69BbFgDagryR2FUlcnWe4wrt2+mWafoVhlIn
GF6ZjFsINVerpL/+PMjBIMwBNaKV+zXMo8svaJGn+AR7CzpRdUrKrAAiFRYm3wnBQf9nJiYQ3f7e
wot54XRZuA4pTkCbc1yyxph/d2ktHfEZM/Qq+DhzuTvRyW6/Qdqh1+oQGflxxhxIzAfee9rPJfEj
BL193KOfwsEvBXC4p/CmII6hFQkJ/Bq13DsPVS/GAq3LzGdhPgZR4FGX6ia4To1zyiwDLVMcuufs
z1MsdhFwwyzcoSWU4phkARYwmNAWzzjbUCRsCqatODlXxylERZYM49L7HpKsZ/QpKjcGjKy0oojV
qF5oDcnszdRkpgJZ1XVsk1/ipqWcIYrSYcgaI6oSo2deayYCmYxV+1fbvrCfaYpAQJ8R2mk6ws8G
YU6Aw2QXlXpX2N+/zUuS4HHhfRqYlOr3WGAOcpB6arrx1tAIzfaLrmDyTGSXMiRxDpp27l4AkTen
fXDAGqm8NGJzKfzBduozqmJ40raB2HIkWXmoFnx5Z+Hk+7ifwkNg1splO8A15e7CM28ce7+iAOG/
7k8rd78iW0KC4vEdoslL5RpZ8o5aScFurJ3r4I714FsnmQAgFQ6Fy8Al/mwMO8fydSR1DH27yZSM
DTmyIgJA9w9A/sk23adi5iLSdXcTG4NtkWoebYhMU5Dm9mefdp1jeROW6HYsI+yF4LfbPXC6iYUN
nhxZh1A8dbbnVGzAM9OVHojo+I2Te0oHXVQdFujLZrRdT0jIKASr1czg3wiuAbPebCfD4BALbxAO
EOQSbhlyk4UQzljbY2Ip3iHo9qdRBkE6rWmSTgf9pbEhBbgqYc25sE0s356J/kIVtyvggrlKRv/C
kPxCc/84ZWn5kG5ohqRIieTDAHx1h0KU7yDGrIrL+vqhTqAj+2PpBCurYXYsqWNgMZT2hF9+kTnv
dYGPjt2NjJ6/7HGF7m+LRhgM1mqgGVBRn3VxACOp9Ko7ZOhO13TksSGluLqFYiTbsunboiBaHGsp
taW+WsbNpOkohgvb2aZ9NiO0C5Zusmcty2BlHA59Uqo2ta1qEnenl9HIweHVwMhVaOebHrc+hna+
AcRJDu4Xe2sj5Sl6/aYfZGmWilca38Xo1q59uEKVHZymMr0Xc22M67nr24LeE+WhAcxWasEyUqYT
jaNtsrAcZBqgr4nDuB1As/LRmpcxfWst2C+SZet9MXAEWeY7yB4d8eiUs63a/6hrMekqT0z9uDct
RHbd7vyxi/kvh4K0Kj0uv0NUyXy3hFDp0A4ePdebsRlYiiKk314snApu14KMsBxEKudSx8QLwdQA
YeN2NQEPsKbaQXlaXx2+ovPntBawv0unXB2T66dJlagrUZeIjCY64iEKdhKqkqb84TLPzgtr1xoL
Jtp/uYRv+RXmH/37ohNWyIC+mrl7ITOpXwAi0Si/MFfkSnkUFj2jiJogwAACQP23YHKoKTQ20MSB
aean8mJBr2SsARg2a67D3hsQ3K0EkZLryN3EAeXCVUrArqhGMdakx80S5VUNae6FekyZdyJEKNvZ
M+SZwxD4Sn43tCGTracCUM40ex3pu+FXzQh0xLon2swR9AZXe6YUbMWEh8J2yVAIQuGXFcA46Na9
Dxc8gEQ0p5wmybH1j/WvsKjXswkNAqcRjgFMcPkUkQVVzuw+grsfgNyDmORXBGdE+cA+anDUAcoA
tvmVykA0xDDDA33yHIHgD6NhxW3qhFaG67fHISUiAklUTWh+Vc31uJXVa40e+Q0SB7OuQmZLtLV7
f4MuWnVHVOmouPM7pyQXmd7i2xW9ysLXKRSJNY3LEc2PpvL1DWVBEMXzYN+LEXLsi7pcm4pyzx+a
3Jhnks3vWVP2//0HoxlBiBVqH4FA0JEQDhOfrOe4K9iYCzd4tEjF3bmjJ5ZMcAiBY7HSsBYxcXih
gcQ2DWF9++fX0oS2yVClTXyS1dhbZ9wMtNHfYwv8/q0dWeQOMMZIpdflBn769CKE/yWMhTTyPZvB
OZCn/Mz5q7tYG4K4GxD8X/rRwPezWg60sZB/FMSCX1UaaEa0E5BYI0+RZ4slgoTHatolL4K+9UlY
jVnOOrsUHqmCKbQjscJtRTG7haPJim5mk1HRRXL7dx17IEEYy7GmoR1GQMcUTnS+AgwKmW43aOrx
unE2I9U4suipZLtM9S7v0l8D7+FyS93YBxyBxnZmzjyjRsW+Y6oB+j7QYzHKADsB9v7vl0Nxd+gM
zY5HRUSXLkz90ebkJfgQExXTpvFavbNCJ9BTbkKZI754060Tf51wMeZgsW7kCfQppcvmjP76fDNj
vUVBX73X1+IV/cK0Pl5N3Ct3R8ljg1dFPeq1aBxGQig1Hk6qEwlqTN7trGWFz3Gvuo/uGzGDLVXv
28vCiQAlFfp7Wb94cMSRoNj89LxlPRmAvdudFUae/Y9IxP6xhQZ7U3rU9MN70RT7Xc7lBS/N5JYw
RvwPBPaeFg81YZdWLh0IrK+FzEU869atF937fpSdzrvfLTbdqMm7QwscQoshVHZfwn/9lFXPiP5R
xFbWkYog3qa+E1CTjTn4qjXyaZvhcH+QNdgpLLWqcirC8Zt9fgtQbHkn4K5bGRx2DY2FHzp3JAYV
k6p+ffYiH1Odnbj3HhD4FXenDnbazePANbkF7sa8qFajb9UBvNWItL19vfXmOWTjtTHwSGmk9leg
denHvjQ+1O0AzmaH4kKmqccgJOIx2AKbchPQ7f6KjgwTlISeRnMj/P9ADnZ2VZyVSr7yw7l2PfYZ
hphw+d6YAP/l8tf+Tjd47svzEVqpvgaH3FlEBjNIfXRNNTHoutM617HffGqy21bsnyuQXfAMdp4n
QHmVwwnwyl4DM1PuwumhdAgipb0cyNehlGgga7y9jS6vbCH5xTyrmIF05012cgDXEzYwb96fkGuC
l+yLjSpi69Ek0bs+RjkmWS8TjJ9C2DLty54x8c85DAbzxCIE/kb4KaphC5pO2n7fiKi7H6UrUKQ6
Vmwbj2U+KAHgmj4ew+eB94Vv/xwxqG5iDaOXQTgmRs+vBi2aYYjxo59S4DqSERotgM6vqulIIqzF
fZ/J1E/7Zdf3EcEc1+w2AKd8guYHhUx8pxgNZ3kve4vdQSYdp4BIJibeo2aYDjQTuqso1MdGvd9U
0o7aA0tpKoZSnodeciaPYw0UzSnsK7dvnHqxdPM45Z4oUVEONH72Br4rwLgB2oma3LbjD8SIWnDi
QUDcxIqsZiAYZw5xivMVp8ctDbzEzyCx+uTuG85UVQPGJnw5GWuDSFplqFZ97yFZz/dMDhbKv7aY
x2nV665tx6DcOZhIpkcSj+ezkoOXhFIcaNeMRzyFBnPMXLT4s5xtNWHWriA5G/7g3T9YDPuX5Aoa
e5zZXM+DJ++wc++J3pVwRlhrV3il8jDUWnVm6ffrPEBB3gyg8Ip56tJQWlO1RmYgtkYrl3f/SZ3v
/QqSJadGjkSVy+9joQLWw+Ph9nMd0XHne4AjA9M84cYM0XgaC6u8ikXnj6WhOCTNQN19x+GjVzYw
256vEIydt5JASw1BiXWNWl3s5b3Uyvn0CgGsWMAyuCI1x3MezCL2WnosZ30oaCMlc/iEt9m/x6SC
eSNzCV4dWVcZIgO6IZ3wkATsoqR9oH+5jZ6rfosBC1cx/s2bslAWyFwTlgkSz+E4CuFvn1mnXRaI
gZSQGL4voZ0y9N8qJChkbmWtyI/l5Xdvo42SliN/4appvs5ro0394h1yPXtdvOxw2dHX2QMT6/cZ
wExNjGjH+X9VMpZiSvVr5olNV/QWLLeknrEZ5mcih3Mqr2r2LB6xmFY6FM8o6B/3KKpEcYStPTgB
FTiDdzM5zV2U1OHU4gtJuwnSnjJuBURVpKhV+i0zhVpDXJkohQsoanQsdbvvI6AZqzDrucg8tjJH
+5EE6Y7UjMPywc/le0gZtBJrXvFQgihHyMh0Wqtv/E/fn6sP/Z8GIW6XY2H/1LftDavP4v6oJnqm
2lj/13G6m075HuA4DvmhLv3lvA3Lxqd1DFe84q9Gn/u7uDlYfGIU/Hur3pvcJ+5VbZbpuU3Dpq1c
MRGUHxiLRPO0AQhR++aubSEWKY0D4gZ9X34RZbg0uq7/gsdWC6DBvhjw9x3StG+F7GWFGkR5Ra8y
VfyKgXqRzA65JuB/HFFRIB/uT/vle0aKtYd8sO0C7NvkrO1MSRN9JkHOdQc86x6VjLxLAtlG5Ccp
D/CUByvC2TMvVtaBjP05CVaPtcnj62qXqgJCrK7zNvixdIKz4kGbCthfgq1I86KyGjjHaGht4m/J
yfyXZJfF8uOXSf6sNPfjqYUhypRJZmNybj2eoxfzyTlcUtmiQUKbZP5pfdu90qcopEdfOF2+9ymy
QVnAXDrhc+PcoF/JdBugIePwEt5/xlBDpZgeJ6qlLQtUpsYUOJK01X5ezvpm+gh96twIp/t06nr6
5+5HpsSIsPBo85q4UYGFqI2SvJ47btvwqNtO4YHg6kzj/D0ous5Ue88RwvPbfaF67BjHrBeEnOLK
J6hezRMSowtJNw5ni3siNkAz6ZK6vnRSxOylRMKB/AFhTAcnJldrJpYcAul+dZfxwb4A0QjoMtDL
zhjrP5wV8i/7cg1m5sU+scS44dnhVLo0CVHGi4zK3BB7orZC6pYffe/goqaUQZp0DOWCtid4AZzU
Kka6QaxeLQdAbA8OdaQTYEfwVCts4QLMDlIQhOW9HVxjzACqWireWWhKV+5NJSow+J7UtWhSwkzu
Vb+LjB4LI23D23WYsgqftGxU3Z8dknYpRwxg2Zh/o1GwAkjy5bfYwtqRSK0VijYR5lqFN+i7G/9n
lLLlRv2dfU5lZ6XSOGzYRE6h42Tj2VMf1l5yOnRTulTma0sJ+MkDpcgG2dpiKuXoUc4WuZQSzdg1
AIMIKcRrG1M3KCGCnlGtDxLZXRDnU0v6ltsKlPCJd/2tfXbeq4dc0CoS5RtuOCFoeYApaDhxSdYF
qZKf6Q9P56dSBIp6nMKRGWDiBxxi/0I6GO6Ah3gTeD3q12dRZGh5Td3TQIRLTbCEA+8sgltJ70PI
m04Bkl36DHx4clUOJ+8Db214lf6r6W0AUJzeHKt16UEKBPoGNNaANPnBvfB/XbDhDRGDaQtgOv9h
LxCWlq1AwciOKOPu94uC7f6XaMMx10JBh7g4LnnX2aI68qthFhbE7L/xI2i/ZQpSsruX7TI6RREM
Tv5lxbOWEQUG8y5AdoBfsn9RmSBIMAWRebQSfyCiVKxAcyqNOI1zRNxjGeLrJt4kbAud9PucsvQY
EhvlefTkPUPrH1Ni2d+uBpSqlQnmJJIX07FWLa4WVkvz/mkj+IIIe9eTgFY6HWKA9jPs9O4gyx5D
VfF9We5nzZ9kHeFG9lZkMoR1COi+cmb0JA9MunUTEzXeUqMoMEB267Y68+ckIGAHOjG+FHoKk5P4
ugLEX0X7bLKUxzAfryO2LYcVVRa5lgbNiNFxMEqnShpXf3F6+KWGEt8hV4TMZ81DK9ew8SoEAKer
gIr7HE85WwgyaP1n5c5OiXsK4z67BmUwTmDdf1oopjEreeSjTZLNdNhWcBYNyTb0te5Kj7TNYDUy
niTt0/GmWcFdiNJdj3nMuugHlqhoXs0QfB/v6QGQ26uNydoya77Llm6tVSDacs7l64cm3DYGVHui
wPd6IcyVtolgzurd9Tf2C0riDgdSzVL2kcymOY0WXiUwFbpQ9iJUm281XVAeboUKT9F0TQPXR/Bq
5X4ylQb00anZbNNGWiNcV06bhF1fQ5FjKDCzBIyfPIE57iXwe/aQj1T9YNu0INLEA0f/sQql5/6i
ryAy8wy3JtsiM9egemJwFVZti9CJNyxKDHfR7tlCUklurIomIpY6nsQganln6esJAiDkJf8qRCCM
cV7WuB4SpmmSTH91b/557aHpNIve5Vjh03xu6S++WuuKSiigtGIWpM3hsuyR+mxqaDojBDYzpSXj
qwbJU5RuJSdEeHHkgS0ogO0zyojLUeA8m1vib+mUAmQR96D44Xf3MEnISMKrV2121zCz4aQKJYhE
akx7NRzF1TbW8nb61KZdDuSd+49V1BVU3kgo3u4lzriDjE06roRNCea7P49Ckjgyq+Elhpj5IrWX
ETmuOnxeWUETSHoDOZvvasFE5Ttz9STUDER/ofktqet/x2aoe09z3Y9nC8C4SVEIY4Yc0dRHGo19
BtYwbUCBBFt+1sQr9VOMcamS6wuVKhtXWBqr72jLRv1HAXDWwAFA/HDSCma3AJV40fK5PawgjMuD
WY0uyLczw1ue23j3QSstu+8+3J5WUrng1C9AFy7fTKdyaJuj1d3gYEAWTsuCvGbOgp6jJRs1uUUw
+eiZh8Z2MaS4APz6iWgXYZdS0JIa/Smy4U5vbXp+iB0lcsHXMcMrRtCZL3nSEY20jiMdnpPTh5i5
x8cGl19l1DCgot1QMGZz3z9ydfpBYVr51ELN3yCerseMiBM1NIWjyww6NHEzofWzOh+2PNfQDciQ
k4fbI+9mSLfNTiYtgJPR0areYJQoo44rEXjFXFycv06811RCAopiQXBiebFkchEcPl9YJFf2BJuW
ATO8gBRRv+/F93bWrM2eU1d1BgXf5pR20mfWSGpaGfO8D/qwcXJHMjtim0KtzfPv5oWN8DNJGaE3
3VO5s2U3KhoLuclAr3iSvvdjpAejHmX1ieELca6CRJ8vYbE7SisgsZHZ8CIJSF6z5F6zoTpr2CyI
4gmbu1fdOHg9OQlrv61o1laD0KlIxrxHHbf4sseWcIPhazkwHazAuoDyR4GK7mZVBadwZj+ifUA5
qrK34BVI+5Wvvp+0pJD5NDuQhm1O7tVu8q72+R8PlqR3rYZfhHMP+I2v3vNFtOSO6NgLuqD/YkxK
s/N8jU6XcZjzGbh5pfOZwSPl5MU6NipZUr+dBtho/0KxwNOdpy4w5Xj0OxvwoNveLPRGptnG1eOt
5Qn1m9X+wOEFrvvwJNkw6QMAaIDd2gHmyxGbn1m5/sVa+8I/Impj9PBBBmP6nRMmG30WmZHRhzY8
J0lgu85i/MZ4pgT21K0cmefBCNTm/Ve+KI835KgHmP+/dwT6zMZfIWWQL5FKWFGnsC+Y0h6Yyd9D
tjB1ruWTuVC8d3XeY3LNJL3vG9Vyh6oSy8WussREzk2OsQZuhJ9sP6f4D0mQWUNnfxPaORzMUyQ7
uoJXILI+Ie46Ak1M/tt5FXRURm1jH0TmMQArTmBnRSzJvvW8bLxG6XbP1XL1kEKVcJKYkVvGBuwq
xvyv5TcDHdf4EbpcNpbwdB34we7RbUSNRJu+Y9qtjfv45wLpzchbOhlOsFyfacbRwSmK2FgXXYuy
kANnyBdLQUsdSm/1QlgOt5TLjprRaqyUAh8i5LFwfDu8FWLvpZMlQhf0tR2wE50+BbfVuseYQBC6
Bg4cJFMvkfH24OAGKmkxiI4zOO4VobFhzw3xjaASS3ANFW6ctUNwYJEAS/BXVtlKyO2na8i9+guq
R0B1B9bPcgCrTVsNDn0Afv4Y/tCYziB6ar4mFEfmyhu0N2iXA0bVfwmz+T1YjavPwRl7lCTGVJME
0xjoHE8DZex2LSi/wrq2XxMez57JpO7WF6vT8nE9LGFQK/+0zJlg72W1HDHm75v4xo/nOnHyKy6y
C2gy/T3nR+UTm8HMdAjrnu+pIS+CZsXjH63fD2AmBSDHJLDMXrk93V1OuC7ysSmmKh694Nybuz7U
IehDfKCVkovNu2nmptXrLPTiFb7XJ+ez+LJFS+vgt9xHvr/FRwoww7fhms6pymDYFQalVuXIYJYK
uTazxQNjJaQIIeUjYYEo1JETA6V7WpqHJuybknX5/cKrJKh45dUvBQRrJ9Br0xTlMWof3RLYms9L
yThVIe2LCpIkXyH61iEtnD1XY4kzvw0F6bvic/bnPbF2tVkBxBE3fP+KuhvdBL9u2+4i10Y1VW2v
vg3JBUMBz8XZkYcHAZlPGZh1SQg9zbmLxzOIKx6TqZW/pF1XwplWGvo136mC4kuopeKkEmiI0U3+
WvXFRaD6X6UjMuu03N6JdGWJJYD6Lf85VonV/bIFuDI6Occ0Ok8+wVR9QIi54afm6NlbDohhG35v
jYdAOxZ+nRluRzoQhd8HTyJxq2vyCZkgahHtOaheX82iSOhtyr4UiFRs+5umKBJIE2Z4EbvUS8GT
K6ETN/l1oOT9l/8fFqPTaM7utFRY8dce19jNb4Oo0ndhI7XdrDDLbh1D6rEzm2ze5/BRx9l1Ddsb
hAPhjqvyTXRItRjUYmx4Du+3sk8R/E71+O0kD7dkOb2IkvEE7piIOX0sDirf+FGOHAhyMDOR7BP8
CKoHwIrwojUWYgg2t70dZ/JoSOdJ4t10GHzEcOzbsOc/F/Gq8C9sF18ctxHVoP+CFZU03BEdPRNo
KgIb0M/+pYfLcaI5WLWz+LGbn/0HA4TFzokJ6CrUkYkVvwwYD7ZRL4cSaWszsJ3IVNtNIz08vaVK
WlBPF4uO4SX1A41yaJoVDhhjWHOeZQHHQa0sPJjfefkaLEdyplw3LWs9xrdEqq5YYmJVVSYTXgcE
gUfvFx6t7LxT3+bKfccxMjnBta2C5tCsvkRPOxzfPj8xwvB7YO0bm9Yk5Qe1Wd36JQRCDs6zAchT
BX5O/vzaOKOcODh7iAgcueUSq590LBjF48QSoPLxN1IY1FCCNbrBRG5LGHQKskOMMecji6lR0h9H
gKSDOzsz82i0M8LH+E3cLXPnidXQJYJW8RRQ0j9SPMnDsWKWNRwVoVb7BfM7KgH0g4dtFO+HOeaf
Qp18l507sGpZK1Ok8PL5lPWt2ueIWZT7h8sMdnyddNAp4AhG+zQhGu7FeTgofTh0VFAH1BnR4ws3
4ndPHOtIoH19Zo4rTPEfknNSBsc6lljuf2ap+CBVESPNQZdCLJ9AZcEa7GVsYq5UCDFjx69tFmk5
N9pRsoEJPU03CpSQt1KMxaZUWUUrUuZfaE/mqF/dVmn7JsMJ9TOQxx+InCpL5fI7bgXb7wPixGIO
BpRTDvgrbQ776dydg1ERI9i28JAZYAZxrj8T3yS6vFkIdxSlNRVHWKd/hyBiGGmB0wHXDop0/0kA
/acLvNykXSfHpEJLMg+kFkPCdCoeOGrmMByt4NcEYCLpDCnXKSa+17kVUAKRdHVB+4+UWiKPZsPM
hDys/fj87SK6Qh2kRJ7sNneYMbDWlBmsz6EBfUm2ARHIpWr/T7Z+lnHy0wwr0LpsvKEPTtdSTxZs
eqOc6J9+Fx6QqD4RTePwYvfTdV3l67WTaD6h7iteZJ/HNvfNBf5CAEpQboc8E2EF4ojvubNZS6bV
oSAmy6emzVK3BgmWY24PXBSwe7l1wxZbadz7nnfGEAKVHv50tMNok7d6Z80GbQhitiKcXvl7RcEP
HchjtKE50rBGad3jNU+Cz+zmxmoAqxKhziCnloDaACofW5/wjNxMvBjNbL87LxyQQghYggAWW2T0
qviEP4RS2bV6mIxyzTTU4l4NdV3zR/tsw5J0HiCPuga4EqFLpgF8YvDEHasBewzmz0vkEKDwyxWv
SZxRfyzzkNWQpw3DZy1kZlwesBY6ZRAk/Ga3o/E1xaiKmLFrzjQ2AwmVIqedN16VcJ55+FTElcXy
fUmbb0OFMNP5ZLTWenfeBde87d9C5RFcJsPtB824dNDVmtigb8hwbKZtUDq3/MZCJeUx4cv6baIl
zvPDktA0VFDEjJ04kmkviHiuw3UTR03I2ySsj39hDiV0dIM5H0Apztweed5ZIuBNGioihTGhKVtD
Ll4IgclHc3/Zj8rB2rCCU4H9XD9R2jNs2miIPMUthh1W2mr3UH6m7NbHWvSL2fCbqImckEmW+AUR
F+1l8e0VpmlPCBUtajf3hpbp6MnXqVjf1fbvRBeryran9p3nFx9Mu33t1J1FcA+vdEx3pce+/6cW
ALwMBIPLbDdSmd17hHyQaY/wGiFMyGWkRiZIOsn1tihwUgzLMkrR4R7kEJNUwzXSvw/PWQayVa5t
YglI5zS1qSqUYCfTGYMvlPU923Y3shnOjItH2Y26SOATLQd0ZbatmcsiLhgZvNrtaTTrZC+weEVv
G/tQqGyoDQlVpejodNd3/fa4N6m9lZCVq00gnsWBb1uE4np3X7LpJpCRNV/bmBSzNL01AbZwUiYh
6JR/aD1bw5dl9juTGrg9cTC2eckgFxgi2ptqfwXHwQfSQdPaqeSmK/DcBXYEddK3QXdmTsj7fhGr
uAHlViH2hR3q1wQzjzlJNELnCltjm3dMRebXIdERpq8dT+t/tiwRuFwvDRONROxbh8ftgUoDsNrB
1c9JHNbptIpHiQI/7MTZ1J0TC6EOW2K04PjxD0Nu9NCgreJNZJkWW+Q9LI/3OVpHKQdC5S5dhvHV
LxCYTZoyPvgVk/gn1b37g+B32JRSzifwfChUXqHaQQbcaHuH+TryqOnBEJpw3+Ye4IE+NO+ky7oh
c+ceAiuHmqZY69G0bDjpTH+1XYzyX3FA+CRqx48PAOAaksTKsvgPYOAGv9WHqxUPV+o5IbRmrjKU
pxJrSTb2osvyXlF1ExhEdTUujNATYdXRcUtkXBvMMZuDqxhtlkHlwAzBJ8G+9Wv9UYu+zPgxpTqw
JU1k1jrve0SfILoNbWdEau485dsah7aTNdmFdERBpK3o/QqlfnM8e/ztzPYiWDFUP4KylIQmMxIj
D915LCjuqhmfklwdKnSh8qZxxkQb37McLK6ouMJR8069eYh56DP5uS8X+e6xHFmdTOjAtA4xEdTs
YdLd+4wuE+2xh9yYcVXpQ9flQUVDDhYzMPD5MugC7eElSgIF/TFL+zPCn0OuPyUvyCYX0j/FMyTL
nvRnkpt8gGT68SrMYEKVZJeFppeS/j7ius3aglHdoPpgA0fuGGLwu7mQfgXlD5EhpY0f6E4E/JEr
0jpFetRI8a843zaHQjEo+ZM9SQMTecLFKfX3vcPGXF1SRkblq68/HNRO+WlbS6y+h1KomPMfO6Pn
ADJtpFuoc8uBCgDeBgamYOxXXEP+I8Cy56G6Vgz0PKyxaLetm97t4sN8oe6oFU2fcELmlBGdKGao
xf0aZ0i6/0w1L+cwC6cYTVvHYFBOOsuK1sr6JUafLVTOfW43fClnkb1RhwSZ6DJ5q2TK79/OdobG
88zKm27OEM9xeeqS8JSRG4K/ai87OhqQmadaeqXwxsvg5vvPhcqwALQHrzBe59GJqjAuocV83e7J
dNRSe93fbvAiNT7U1UnjpVS/OFMG2eJVP6ZUzJSclQXeHy6rcqSr/PbnDGm3zozUVFUPoFZbqlHs
xOeUbUb4P8Ysw1xgoAFHGy6QpBGLRJUx+VyT61tMD95TZP1ZETe9xBYLILkUwmJyGMuFIMJyK28e
2J70zMtOARSJIm0ukWe+R/kc94Gke8pU/1KPw+eJQH8q2WnuK2wAbcPPEby0kYOxJ+Dzviz5RT42
DVNfjFTOCjhTa7Dm+XOw5qqVYwWmuAzq1X0AIzWzEGaOjPDDi+tRfwdqC/58iVffeyeXiqLMS6dF
+U78LrjUl/Mx2un7hDDmU7u14fDhjPzVxHyWzN51UajG2AN5GGanZPjGD7CsPK6PNx8Twh04iwkr
R/3CNOz/yMJckxKXX8S5ytiRTGQvqrk8J+s/tJOVRYdDqrRV+EwB7OZDYQbBbSfzJUD7ForEqKQE
7qEph0p8zU6c0EQ0CVvsxOyLEpMHqA8cJMI7/PhgojPAwEFwJ2A3hLiL6CwNZF7gcJyXl6DQ4atF
7LsXe/zfUDSu8zpB8NPg6aTnv3jHsLdNAc5Eze11UH2wZdzppJuIUaX6VDQto8H0WU7FGVHaNqnR
0f6CiMsNKZvVMK2tVjYDIrkbceddw2Gf/2AMPNEJ8wu1RbHLs19L8I5dCcd1EJTMzzaL7QOi1dQb
u/7pZhbrfbRKlFQtSyGwAFYd038pCFWm8hrhJkpbmE6cCq5VXC1VGeAH8l1nzxFtMTN2KMvb7xOw
eGJOq7b2i07W1zlZGANKnQzNusReZ7MgG9LfhbnaneEpaw/BINB2ivDyXD/BvTb7aD+xKFuklK1k
fN5LCSaCr5awrnL7R+Jeqb7N2yzxEx6JUi5YSyvFY3uH+zf2Ny6eMRV0zbhkyrBd3plvbOZGBN7n
bg6fvHqBRbRmozX8LLe8t9vAq2TRp6WwdaCLDEaupiMRVooHUPNjWEdX1h650fUoI+x1JXRVlrj5
RlX2fEPvZ4IwnvVACcl0JsQtdZhLOe5x6QEdpWCWrw+cag/+88aDFcC3ANYYZpNREkE8kmouCakV
3WyCfzD3eXmrKItA+DEYkdpB0hZw0s4jPqi8Z/6qd4rPeUxF5SvOV2rJP9Zl0Nko635S87u43rbr
zmuhQPwe5ZDUa5akcGOegVRObbfG0MFvhDScTSo9JEz1dHubZEx2wgU06lJJUnLFiQyTe0aRgJXm
UcGCK5IRCJKMB+nK3c+gq+bz72MlPLrw9J8p0k1PJ0pQQGUnaWY/GnQx6r3oljy2grkIDGIxqtBJ
iZXYyi1pFG5IQ7rbp0TxtIEm1ru3+YuM8T3d11QAH6OSiDeOuzb/jNWJ9p39aKLCiXRqgAoBh2fd
ALBLaLGbsronGO7uW0GmtQ/ZPL05o9JWQF79iS48aGXWlup5zS6PeUZKtBv4FsmETGHFS98QKpmC
aYhlpy/l11iLiuxJowXTVQZRtLx5D+BAHkXIkkLDgU/WOum/A4OUF0i4mFO8cjKoLfAwzEQ6QXpm
mCoxGw9NyNqp3ShFDXRTne5xgV8vbaGaEWC7h9+WkLJyVQrqCdJIs90CihUH0yU4uz0wc58cnTPn
A82upugRiUCF5WxFyRsyb/1Ygs1l7zDuiXrNe60hWJHvwuT2b/jBeHA2h4tBoffKBJVXFpOzync8
eo/GGiUGZK0ARs8XdD/dhUFvTwjrbEgCvTyBIzWfKRf0l4XR3DxirJNA5xcVkWh3rxY3P1LBwCEY
hW6314judhltMycEn5tdirmNHnIsF4tqiYUZkYe0EEeDpKVbBD/pQTP5KH+x83szoRTHIWFxCXy7
B9/yBXDrQNori1LohPo5KxKrCL47M0UTboHQTO2EsokvGHhSsmb5luIMDuNwWIH3bEdWR3pNeR57
9FTRi2aQVevNzQ9HnLNzrhyqdpi7VPUe5wWc7wu++wxyBS39gJA9JuA0HCRcWtBFIJ1hqq8BGIRz
KxFPbCpaJ+YK35e8XdgdtO/vGEfkwV06BEDzL1m9f3lgvgzv7YFF59SJp2N3TFFgq6yNz8IKcd5N
ihq8nyD4wfKdKUXjMFjmpwVk3AwHk464Rni1OfiepISs0QGHdbZUq4N0RLGcZpXzr+8ibzzh3OOq
/reae3KD+ul/n/ajpSpM8kqr16kmMO2sVBWfYH4MTtcrhYLHgJwr+QS8TY8RF5+F/QTRZgLCQ954
flBb6NgVt4iipyec2fIIY4pfk/3OsU+ZrvidkRq9/hAvnesqEnFD+t+5S9quJmwkhx9i3yCQ+TOE
MJQQyR/qLwie5d1pqPT9M1N1UAyScNU4XEE5bh0zxhJPbubdL1c4TvNQYfDkDlNl1O32CIa8MbXA
qim+CVFeIyQZlMxseeiJBL02knbDNl5hMgsFtmiIKa4DeD0jzU/khBup4CR5eZdU3FtysQgJlnkZ
ABfOBg1oD4R8GRHURXbUk960ep5nmPU+gZLC09oliDuU9GAJgzq7dOMctu4JY1mwxyt7Z1ZinALw
CCCfQGhJ42pbrPHHlYAcF7FN2prh4ou+HRfQyOpxszwcHqzQpsX9WVJdCe46Mv72cwkohfEYabTJ
Kl7akk1BAKWMHxB76bb521z31yqxd2sdwZZHoGrknFlOdLS6ux5wQdYJ9lWyWckgo1YTxq+N3Uy/
ZyHJ0szK1ahJmgGyoZ9c+YCkCc9YK2ujFXIdLMQ16MWJbIk/6swFZ4s88oU08fucaUI4PbAZtfuK
ggLRfptkOYrrEL8zGcqwbFAXuFs8kidjVwXeMs5KkIMJp9q3osQHrEJdJ0WQQzRkKmMH7qFvgYjK
y20u1iY4r5h+V7kE19m5k/yxiL4Nl/WiY+EKIoItO9YKwi4zW2H/5cjwKM6dsETKYLl8OSQq9iN4
f6Zfpnk4Pm7v0//D/mvs08bIK4AbcOBjh0rKOnul2oi/wmGbGIzHja67+qs7g4Mj+MtHF5edSX3W
TVh3o08t2qaJ8Q0VhXha5r0fUMgAk/CZZdlRoqzMYkq+H0t3mkHwn1Umj11Ev8wj0ke8Cd0CYcXc
vMOG4/mgv/TR6WYkAmayjnAQw6C286b+DyA28HFlTWvd2pRQHc/+6AFwmrpWU2PtLMTfqvCbKAJN
/plrrc8VwelyVvt3pZL/VcB/O2uiG4k3M1IgBEdmvKt3P/Znrk1YcZStZphLfPDYq9viL2ouXZd9
JkYYo0MxBGiXID3BBBqNGYbg2M627Jo1NU0itbBrruOV22KuPmvHuvQwTfLFHbRwu3d0qkbiID7b
hxZCd8MJJHt+TyE6egXUObGbpcaVvvDXHgE9Zgl0TcKAyw9RxOIk3WN36vwFEwIXFG4FbCAB5Ksu
zavP0agJFACfuaht3YWXtxt1rMzQQvKxKkgkpcUNgo/qL3Mjwmq0ZxxcqbTOi+4a7TstkLUW4Wog
JUSX9PImDldyo9A6oPS5sxMkyRjvmipelgHLMktPji71m8nREftqxI6Uagj2hAjSG/RGcW87/1ym
WZWOv0iAEdrn++zvNwfBKypQACQKWaJ29oVICBgY2M4AstowkprhKghFrxL6ecSlNcGuext/uicf
UYvd7vdBOeP3n+qmzpMzd33kkhRbmIfPblZSmxzfVx/223ihNL4Vw7mNE4Z9Tsg1u+zFRAjc32SL
vAPSMxsBLyXcA3gytrf6YWibDNAdRyCvfYQCabsRpXvMwUehoBUrKKok/NyylgD91ac2078/cAN2
A5FnP4sl+lOTRo2Ny5ETPM5MS+dpaGSYQ0ZDSnVDTbfMgW5WpIl1EcR/IiOXMiI0viqLrwsqhBf+
kWesM7lgDLTXzYqVrzJwHAofsbMfWcZEx34TTaY9T8c3IDhmywpQhC8DnMdAnFbTwdY6QrAJJH8w
XqUffwj6STnTjx04D1yDkcHH4UAfftbftnrANKJqdGwd3KjTa41ZNsFxOy+5G7/m9xpaR1AF/J4i
jvyYExHyyvftWtHAsg3wJ2vENssJSestLZ0/Yx5zN0WGvjUF5VQmKpqg2DnHVxwFFjRovEs+NbSu
lUyOWHeG1/+rkVnrww0ycQm1+qMs94eqMkxf3CGZbglBpcCdBqmSq3pPDPi9uLeH/GvPAKEa1/xC
WJnPcOlJCVatZLSRGAoF0yOFiqBJ1Vutz04vE3E6j9z4YK9uxDuLLjY4kd0caGYrqfdDcoGeaD+3
d6wCmxpp1nhTmJCdYYdL/Ehydz8HQDwqUD4rTKypv3iVfHI/0kgIY6gd0IcfcADsy+qxz3ifklm8
BpLXZ9anftMWiBY0d9k0vHtN0CcJIr0GJpIkjqVzaaHRsdVnVhoIjlM45tGifJTWBtcnXTCgjn36
JBvhkwSMtVYjUZB0+FXSIQWd+Am/Jn+HdR2fKSQGW9fRHb4DbwMHDMpZRlOsPqypgRNeAmhrsHDc
KuZ3QBIUXZzNQDoZFMN5oB7y54ozKje7e8NdlURi2M/XiaJ4Hv93XxgZ8KQhLEKFXclo0wy/Q1jP
ZZHpeWbCAcF5cL+gahrKggZihmV6fd0qEB+vigwamDR1ER+BygGsmxyAwXMIeNf8cCSjHR0nESGp
zd4YFGjnS8TRkw+GFrIxW5bumrB1xYLpdl6fwEzDOeOOjLe3Qdh5Z+7qiKCklemPJ3fqiYSQ+8F9
NoXRpPG7IBMn0a6mVIMwykRoPeg5UVPXArzgj2hnXhA1cR8AsWwLyV99wshp77P9Vikk56FKlIHy
VG/IAXTtiEOc6qUgkDMmw0qXxbmUAdSekcOmPiLlbw1CDZqAyBB+xYwW/I5rJPFo3NwuYlHSCggu
BNTqmcyXj1mtMzWMtj+8OYn7/ysEnqNPXq/usKQIfxtC2eWVinVA/aTaV/BjgKyF19+nkXU39ZmF
lGsG+oNC0yxZ5ulsb0UWDBXe55rkrbmjTFFhITlSkyUpfHhYdYjGoXceebVPw7wt0ucrOAlxZIp6
Pn2ZbYXVsF/+EOIJV1/MFw/4nyoyuMG3I0mjxqSlpEbrWZwT/Q4OQt8Y+QSlB4DGTZj8jfWdnVWP
PLMmmYWyXCc1YkRAngCvhdKwe2Kz/fVREhVyGtdXtCX4aJ1qLlF2NykjaiT/L+dP4pxrH66MQ8SC
wpTeKkTv5lVEnc4zDIr/pwkkeCdRH+6xffetbAMD3KnLgbSdP5uFCT3jeBAhO0G76oTZmcC3sw22
ertr2/xlSvsOFL3dKEmyCHj/1VB9QQ9YkVo+tduCJTTTph7hqRX7DmiGrc6iW8471Y4v7p9VprV4
CNykBvioKL4HGJk+eYfNELXjr7uIVjGiYxIi2VnsDBqgTs7gznIuHrvK6jJ5PfhY+WXNlQ2FbxjX
d/R4coAcDm5yJuTOp95QNv8x33f7lkV0YpSTkg4fLUQ2/GED1M12SmhWt8JuhH1P7MHKBCzQk+8f
Xz6Ox8Vdq40zDFBCJy9OgYwYCO15LlQWIOB+p4tPIprkFfNzfZjY/3lKqkz8G5t14g1nvnukBUIu
p+dGzUjfkcYLnang8Dd/+i9c6hdYET5n09fF2uveKevPhfE9X2T794/fNClY5LGx+0+0LwCU9X03
M9kztWmw6MgXhzFf8K52BghzdDGuRPm2eETJ63XEBUotf/vBn358L46DNu+Ju5GyvSQff3qS04OV
y6qD/LFsB8iPuM8MMepgkZKjmxvSKtal2FooZd4lCFTNgmkqBLfmj7m6C62lPWMH51I9i55QQDH4
GgPO7ZCZOVgnSQg9jZz6Tv4imD7qDAL0k3TPe01zYJJd5muZwGKvD54rgwNGOqWOX6SVC7sABKVz
0bQhFbnryTFf5AByyeWp0bpRQ2vhvQwjmCUbRKX5qCoLdUIjT3eBHhM0Vl3GaVJ7t/NXQwTefnSJ
P3/JdGKKtEuqYeeQyIKLZa2q2gyNdrF4nwgm94HaJoc1oM8hdHirtB77eIAxXwKEu8HxRM5wMtrB
HJgM9mX4uUV8i3U+dRCNr9eOj3831x/kgr1qORNLtBUAD7jTvONZj2xJQn4Me5KDvRiG6LUrh+VS
GoT2SZKUUDxf5vBTr7gdqhsxKEw4sISe0p3Ztx0796Juy8cAgvlgaR1wsI6qo1oMNrp0lNkDsyo6
TuxtXwqDx8KMRn36h4r8wQ4mGDz4dFEK+Knc7wf1PFY2SQV+BdZQ12ZEh95ZH5YTnNZIY+kbSh/v
NtT0sspDcFjLowZ7r5KKb8q1vl7FZ2CCFEJjtrWQSKFpe8mFXYBtMJMm7IBIcSH8jhzfFXLt/qaW
ndP+53gfRaVUsbb0Zo+VUMrKtzx3Ho8xl3NraKXni4GzcWH/E2FQe4UqJK1CHbR4J7WXQHc+r7qm
VxclWqUKZOkuEkRzyrwA9CmU0cmxy2lO1vQYT+GeVwri+5Q16EAq5tRbLoEIHuUK2+XHnnlUwrDL
GTwAO1wK0f1BuhPy9GN1grOwVxF9KRVMeudq92EPCJzkgHDzp2vFT7QOAvMnX7lBMazz8h+XivlT
GsUqUZ0B/dj/HToZ+w29svXxjoALBLAcCH2CBz+8vkxlgVNzo3V0Mh1ceE6OgVKFVS9rfr905qIJ
gTO5w2tFzhM8PbGCax2wAqvOrFBjhOx1wIoEHzU2KN3A4YNw+JfU7Zc7VjYzrSoIemZemRxHlGxh
IiAJDnl3/7iIblz6nnD+JkbIBuTPqDoKWRrUBnYxS5PL/Qe2rBFXEMRGK3zTgSsZ3XS+ajf+mxMx
RqJZWeWioP6z9+9WI9y1i1W62HqBevLxEUrIFzwcn7L016pbmvNyo0UsCebfi74aYZS+9rExkqo1
bfxP1JtCb55n5OEKIo0CAAP6yeZowPR4r5kYExjrnLHn9CzDV/1RdSPvClM44T1YdP0zAzJRFLWj
YxxGpprw3xr7rVjfxvxWmQ2LNrhdRNdjcxU6QYiuPzdkO5X3B4Uh4SNbZtmt/IcnTXuqodJGlfV4
TtDOx4+SlKJCjrbAezJyZxygHRv79Ti1u/imAro+57x36SLfk9L4jvuTXes65NpNiJoDhC0Le3Fo
6XxM7d7yXEmxqDeJw0GTA2HMOOd6lbBoZspKRaHuAXphPNyR2AaXHinyCImLgtjnKUvA40KaNRmp
Gg5E3WlbfYTom1CrJQxQRQIbxMeHSvQfYzYSDz7IjhpziLytQhRjwHN9j5BHuEF9HHd/OOfOFQU8
tH9JAD9JElzkxxnzJ4QkDVEQtu9JARm/PwhaIscqSym/HZYpZIt6CvoB2znRbeCSEvAFYqBPItEK
r2uVSnq5FHw96tDziAS6KJgbC+cNltp8a3w4/Qwlq3IBAiELzxEde2TRP6kcgLYxHLecXZwtnw4m
2vVVR1ZT4b6/tbMES02xUySGRy9cNV75hl8EknICWNyKw6oxzbFwzDEPrwsjT6Qj21vRdm6Clh3s
uUgK0K+oBajCoW9La1HpkRQXGvguPXQxruy81LWSLrWvb59FpY/7f8x1Pz6jRt9T8sO0hTOSCTHf
NbqCaDGJ8rBqEkHPwH4dQdTYyMbHyorSRDk31Pcq3DpkAUhbTd3rwbQxXtU8rKCOz2Cz+hgV4l5u
LVuvhLcDzgWwEjbtUND1Izv9EEgOI5pCxMdjVcQKKUJQiS12B/f5WHI2ieD1KWtsYFjn4GdJ/wh1
72f8YUOpzBtvMxAm9Z6roiN14s9C0LBy4WDzlITOUibrqGM0GrDe409olg6qsV9R9pGQYaV4Vsjd
q69KZ1VEWrsN00ZWQXjB9mZTEWfIapNo+uY21YqXB0RfxA90G6ofQD1vqFQg7scYzh9Uhh7ZYFE3
rSTJneVTmrZx7l+2f5LvaEQz90/jbA/xENtr6uI6JCgXsb+ioS83MIk/SoApUt9JaKI3XIkgrQOU
UdtVQ36CD0WLrLFVHF/u1zOp4nbxDENSL5ZBHXRXH9eWlG32R1fqDCwWNKf5O1VfzjFui74XJjzp
uY5DNIhTbmJIwrsHmyyq/cm42hAH+B2rS4W8MpGQmUuFl2HxHU+GYmzTj9ISytG3utjdVGNzqL36
OCrQPTioDj4HX9aYKTNQ3voXUNHK9mMXsFwWXi7Vu31b30VfOlmRzPMrHddP/6wHwnNifczOMCDs
cRb4p2mJeR3qJ5/zZ4iCy2hFLtxcLDK/kJINIEBwrXre2gpnK05QnQwXxauOwzZf3v1PoDygfoKU
/eVsfLJFmo9c2y5y6PXJ+0ufZBM6Sj+B4Dp2VXA/Nw7Q/Q46v84XTWucmWvrOQii3zhsdVgbxge6
UAkhQNiLpl2TF1imoxqbVcDnu++1QvwUqihmdyQGLly9R0P7IbAYADVYvPW+hIXcPesM1EUZq5iB
RGWdgx2qvTwDAefxL1B2/w9YKCStC1NilkNUHb2DrMt8vqc1ubsF6aj3tAbURdBPSultXQTTZXIe
rRcdK7zgNVqWgm+FulYjzrAMiXCe2zSMGImdWHSI4yLXn6wE4LpKL2SXdk4FL2DZal2s4dKRicOv
GaizGMn0VRy4DxXxKPyHTrmzdClYeDXRWKFPGbZ9C4OfKZO98Kcb6hfBOTdNfD6bQJDMsSRkQJlT
84yYANqsh0zKoiNgVXcg6whDAN9nLJrHm8DqU8zpDXEb5Fyp8uJ1x2bccD6bVsHjmpsaBGooYtJH
DhiC2ftniHREHhUJ6J5X1l33REPB0garztWgnCx/J08QskK3EvG+LifAmXgEwMqIwR8rm+m/W6ez
axG/9GuGYGRVrVLZ0zyPgeQWiEGyGt3K+kOCgM/1R0Z9t8NGDuJxrRTX1zv6cdfe/ywT91+shi5m
PpMpZY9Onf/Sn+sDk+Ipg4zNqbS0p3NnJNrA18pV/EjhyT5MrLdmZYLxvbiaSQ2xuRXmI3bqFnlc
6z1WfZflEGvscqFZElqmCJjmKT1/gfVGXgXxdbQ5U8mWX/xKKJlZG+SUZu+GFiTHZrPm/q9yv9rd
xuU5JJbihrho62dYRoBsHRJfBWsHZd5JdzPMSWmfYdPf93gZ45/rSS4LigcgQ8jmmV3YFBfExRMD
ksff9CgE10ScfJEj1oMXxBMCUdAOitgM36vR9UtXnOkvrnpfmypUcD6V+7g3i5qcMaOvQ2wYGIM/
UcFY8i41q2vvBQbsCavE0o0Bmw/5AIW2tgQmOIxPM6wnXn0twqDeLaFdWcPlH4J6sFb9jKqJPDri
117lSMAH7tiyqq8P39+wnN3DhjKaYVzcj5uG90gVYAt0Zt7fMQgejIOgkx4NDYaqhgH8UScCdwmk
NGLdzPXVj6Ch+F1wyfX3JiRLWPq0CkEBVVEZJfYSkEmqSf1O0QpjpH9DYSqjrqHgn7GGbXdNKzrR
1vNA1T1SgCwrZ+L1HOJE3FGHOyXmHq/wovY4y8/Ai4LeuZq9xaYGgp67op4m/oaDoqbgIpXFcgZ/
GJQIOrSFPBQed1sjuDtA0ehBIiBHIXcGrI5QgX2N8JCXTOGcfp9aeTG/Ei5OLneAoR/7F9VCL78j
iFoolsfMQ7e1sb+rqqMrjJc4LfszdPcOR6Svf2WsgenqeTfFr4kT666ipj4q54/qOE1QR1O2g90k
BxzytGMMlhSk7Ks52uxEQt3x1Gxd7wdMDnXtmcx+m3hsWs4ccwCcJIvBMZ/BNmqiVU7glMcD806X
MOnvr7H4Fv9EEyT5/pzV0wEW+xKsuxQ1HyuqLKFaYDLXJsfomKNEWGqGAF9E9CS0KgbTRm+Qm+2S
rCwmhm7/lr/Zd5dSiGqFNiH+39BnBmxtSmAo7BiSBha4G5E3QvEzDVM3PlZkBkRt19URdjMofPrZ
c791uLoGvpzKy+G24Z5Orwdv8VMaYNj8INddF4jy28t9khAQMkTm58wH+lriSzSvZSvKgImvJb0P
RZB9l9HG/LRuKiSo4kGj6dsFvKGKZP2BhjG8+71PrgsPsGBItJWvs6Mh0goMwldu12p5dKWmPoqw
DyrzxaddHJAPhS0XJ6wSIHxt1GF67xhfcmXGf1ZuXZbWPuh94VLmDb7kHZKF8Nb/MFMX+7LrECpo
ZQpVJHNB2u9e/X7m6VtWnAIe+OhcFHowCrLF/Ive+R+iSxqPkZrTMK/Vq9NaPUZE5f8rP0WSof6p
wPodJmLlP1KvieZKSYQGlm7k2P42amg63SUD1KszH++8ntNFvVn+ddWU+ZGxqefV/RjpPUCAShk0
t9KQJbuRKbW0ng5sSzM0Ctncp2B80n9ZKDolIlVut7GUdsq7r/SbyaNTjLqjivGLe/1LcAFU4TIh
naJ9VwTm4q0ZiVbSiaie/ZuflBpsGhef4opdbqXI1MlVvMydBzVKSgGmZoxgL0f8xaok/2jX+EpN
fxadevD1u6QJ/hT8nknAgRxloQMSxDKxfLop8AjOex2BZBxu++nf6O1jCkH4v6pCdt9/VhUMAfGg
VqGUQoSVZ9bcw0OHNIgtnnvYz3FshURktytfcTWyNnQikA1IcbKvsODRksi0M+QXB2BRNooYMABz
zw9/qobMJtHLah7Tm9j+p0mei7jdjB9bQ1bKNSMeS9OHM0FN2VfTpIuXfYNdWoYmQ3rsPalCI0W/
PuSoGBt442qMPGXjp00FlFduBQS3Zq1k/8JCPqoCbPJH8B3j3qpzKrKcS/y+KQ++ExxC9iKGafEw
UjXtx9DyHd8c1je+LtUxmXQ8D9d4x6wwwHTIX7AGwaRWdbp6XkJPcxOe/teQMvXltqXjodNrFoA0
oPM/ZeItXbbUGlygE5L7dzKNIc5I+KNV6o0cQOn+xbYwDmYfcRoDBGQvkl6S5Hvf1xauH25Jz/Ym
tcnT5I8tXZRsP++9vpDYNwpLlgstyz/FWvMWZJp6aSk9GCYYVoP/9pR4YTMY7GKUHc8VOB6Op1Qe
+F+HolZ255ifhZc31qz/FzBl/tCIbXSf75ayscYf82GlVrMKrPouUU0GuxH0/SgC1KjqHmWZrj2B
EpUugG6ADvNSZg8CS3lADkJYkHlkOft/jgVztqrWiQC0zAkSPfUDOcwxlzsTboeQuTi/LG2QED2U
akQzdTXhTH7TtftyDsL5xwc9O5JU1WaIWoqtTFiV5xzuwPEbuhxn4n4060WSC5yiDt9lhn2Td0Pz
QOiFH6J2tspC1/JWO21RpsAmDw64/HXv6eWjnWLEwkQYPovEmrHayAgzPhti5JPMLS48eloOCINr
mSG58iYhfFEPdXXs+LWMq/saoXkHjwv/GOaQ308hUIuKasgXNsSQHrL5Vlaj3Nq9tjPbYIZgz8Yj
/ZZSTViaO6Ryq86VlmGoYKDB0jtlBCYIU/y+/Kw6pb0eoY1ryTOdsVQ/gSN+PrPkbkIpU+Gs+T+s
JdxTaFl3phqYk3tqzKGegc2CHsyXOy+/b5Tj3Sj8L2e+T8Xaminx5QaGWF3m67HKZNCtHZVeq49I
BXhjyDt3A4NVMauHPW6xgqZ5kcoYyZReBcdz8bDLotmFD4GRxubWhy+iLH5S2rcBagBQNGZyQTn8
e8vYHTqNjbcw+fSYGMZgE725y0n/2GHcGim6dbI097Pk4lNYoxWo8P5KVf9V8UsyDX1bhLa+b9rh
GVqgQ5VWJn6mcHfvUN0iwCVZrdj2/CAYmsZURV4ByjjJ2uJijuGSemsuInrh3wQZBrS2wbmCm0bb
b3DOrEzwcZtPjLqWymQfkRwOV7nRX1A68lEUKtT/r9k6554wJ92D3aUJ3w8P14iuGtDR8FUOHPx8
ELIZwgQ5aSOKCQLgj0qGyDm1gV677iz75z1Ddlh3GY0R+mISOV46QdyFM6sSJS7HT3mmUdOdyFvb
UBclMxrek2BBS/G++yRcviy3VnfJnI9RDTp8+atXMnYylFpLvykZdAu4EYcPhmmYoBP0PP6psUXc
iVxmWv8no8HcvzDBewX5Cl+vggYy4uVMNqg6RI9N8gAbpnwhOSOI2aHqd/k2ysvIxnL8sEKUYtNf
HcASIYSxbKgCFmhMxKNy3hbW4jnq5QJMdp9iTQrjltZX7SN81dVSGRrmM4scRYNA2edboYNBklyO
eflHz/B7pEK5K1W/yvHU1CfPo1L7WkxvAw4LRR87A7nGVLhmFom7AJYuC7aSZkZ8V9Zjam9zG4Ks
1SvHvLrwf1KB5peLYrfFIj7ri4zgiPUBDlbfvIw3KZonoanSNous/Xm3uuMhJBPzGFGu/RAM9JVB
TYaMAVt2auXGnPCJ24G4+CY1/zjmzki2wLdC9AcOyEkWc38ZlWxqEzTQwuAtPZpTUCIkMPymGe1B
bO0p2jml1VIUBdeQEnSiEAKktTB1uqUe5puqRkpyjfb5npRFpEX8zJj9bzSP1So3KYyk5IoYZZuI
uC+zLm2l0PAaYW1WwF4ZRXnBEahpLXdigZlIagXZGk8tEktWPaH2KqgMDFlkdqniVoGDdTQTeIa4
D0PE9LlTgIye13VOHWmosdNPmL4OfH21dal8gMCTKQnRnpoQGMVLM5LA/KVDr5ItfS/cbEZ/wwO3
8QRzb6HZfxTCgA5FTkL+6IzM4oRRAFGp26CobjfMeq68DWg8b0b+/Jeh7T7naP0GwLaBFhGPs+Bm
0yLkR3C/19CvetXxAhbUvpQYd3p8WjD4QJDn5f0wrDLKHhdRYVt2kch3Asaesr4G/Kpqeq9NyTCL
d0HOHmgW8BS6I2/H3RL3NeEt9XHPNE8T38/XmXWcBqedQ3dN3EKS375KCqQVN9RLw2O3i9ptLiIk
o8scInUUnMJVIN1BPC5PsxCggoodexBYZ6y8PA6iYTZxpESL+/4QIkg4f7ZWSWoTt/RO9uXcJ8dE
oinWvg3YtkBiIlFVMmfrDBFecIPHxs5Wa0fTwn9bC4xrvowG8JAtJO/+bEdFebwTGxNts8qp7ws/
cxriEeFHKH6AIfLz8bEzInmbe/+lWQAJX6gMMWxbzI8hABh3Ux2EmvgJHG/GOiMYa0eUvq7HFvcv
GzdnvFC1PjZUxRGDsVio61lHYcqGnKU9ZU53oy5u3lFfMXjNLNZjlRt7IQSUuCFjDtFsz97XRRtH
CWZ1hHC8SEAJ0TL2mrGNp5sjbA+xxXO/o2Tip11mHfIxREPJuzF45H2UDdvcysZMQKfBje1eBXMg
g7Kxjx/pVXjHAWptCQPgeei+B2jhyR2CWlLeEM7G6PS/q+ImnxQ+Bp7zDYQvy3DAYHEReuh6tcVu
slmBe4mxVF8yRqtX0WBdj9kzGvwYlqhZiOylkaX93ctWlLhra4ljgkEaFBXazTC+5nC0g3cSLb8Q
1L6QtXjUKGOipZdKE2p9KJ1y0uTB14BRtYVSa26kk429tCZfjy0M8RppCXQ8UloOJz33WUzX3M7c
wegLJ7xs1X8GMyqGM8nyEKERoeCZ3oPFMWVXW7mrHM0B02baH/lwHIz+sbuPpN7tZk0EJLIVWEjc
UBfMZg9/ExJ7SB1njSyy5FdkJGp6461zYA23BNcU/c9lrw7RMa3SJXuH23UpXvnFBqCqLah1uTQj
5VTo8VkRTL90YceYiLhVvfhapqiTzaoQpBSX3A7yDLqnjCYrXWV+6sEU6BHzrNl1/HA6U8KF117z
5DrxsD9JEAOsWFwxYch/KB0I1WYU9OI6u9jZPD1zGxS+KHb3PYMbGGEg4wA7unorSbV9/3Prtzxb
IQUG6UBn1OozQf0L8QcsheVuqQH91Cs+X0e9HOHz+VMZdI/lnrIHLHM2wW+H6CKcScn29vSVFNlJ
d3gF3Hn+4JmIkqmU9rk4lkXWlnZhQufDk5J5qcqbhfavqJjjlQJaNUg9Oo1VCtnp4htHMXyI0UPl
S3epFPlZkLS9Lb7Fsd8VrQWHi3FuYTox1uu/5zzXe4ujST2Y33Ng2+2NvSzrJoZQslqhVnmqbGHB
F3Q3naQ3lNWo7sf21nYchcZ7ncAfywA33WcXaVPCWphAyzakbM+ayBmfyr4ME/yQCIrE0zXBk5kR
aTQSpFizu0CQZoVxaHaru+oHhu95mA6s6N+S8ifJMkxujXSM6vVlq4suD7U883a0ut6+7R0z9FRQ
jI1BDUHbuUTPf+U/x8bItVowptlwjmlwpMV78bskfH+VeaN9bMUs0h55dTLUDeDdMsxq7t1dUVZ4
RpOIMf8NKNynW1BLhvkOzWVj8/pnyXYAf5oN+XGSbVbxdGMnf7MbHumU2n5sHJ59W6Ov+7hbnHo1
NFV3Cwy4aRvRKa6vSXlAEZGmzeZk3gMyiBKscpDaD9WRApzt4++IehCLYQBsP2KSUX6/GqXMcARJ
EhH70hknfQrmlkpnTp8NqVvHCG0D+Lpfq4E/EQ9+yryz7Ta7HX5QSP5diWX2t9AO8SVccNCleD1G
NXykPnFnLWgYCF/lwS+kp8ca1rDEAsIGPKt+DbnC5wJq/rwYU3smdtXaGYpO74KJW2/MbHmB2EA2
YXq9OVR2tEnNAEaUTMLjkJ+dHx6IYytGnoQ956D3vJuUN8GNONXli3uIDlsdLYy+3lUxqOnv0zQt
mgQ4X6nA8W9e9/NudXvj8IlzedoKe3asN1GrL4Higrkx/+uO1AeNOLpvWb4w9JxM9REvsRdoVMhN
ArryVA4pmp2//JNTu9FIc5QyHyWwCUqbQXItP+h1L3RlRvxPUY0An5md/7umh9cjqkScO+yCNk+9
tMonsrXrkNHs80u1MZPTb/c5Pxw/UrpeNw6gZEgB1wUBry9HFBE9hG1704KffnL9pQwmbI0nQKib
H7aSL4aItUMJSoI9OxOhHtXiAtFHFdYbolR130W5cBIkL8YAU/1b/G+obZ7BZQlunOJRzD6uuVr2
0KmqwpngaNEUlm3pwIvR7OP7+w+BkuMplqhZuzsU4gUG6fRFf4sZyWDDLWCsD9rDf7eSvL3WIduB
sws+hWi0TSuqvg+IkITTvU3NkSJBtsHiAygusUAK4j5bK7IzYbYp0xC91ku5cSrcRE5kyxNXh19W
zqODuqQUTW36ND6YobNVtG2BWzdE0gb4sNPWV6Vutca96o8a7j3BZfmr8BfWM8NGyb4DSzEEGFlE
wpTDk/WNXol53QEgPcKMbmVAtIl4WAMJ9R+vNkgrDNMgmmDntRiY+ozf3dJ0m4lsKRQePMMkq7VP
mIvn21sbRNHWRBYYBekvwKzxBT8tsi5boxzNleaYCAklp/D3qGCQDp1uMbBytDSvU1uAASElZIY3
oLd/zG8r6tkBXpWTqU7Ca7qGM8VsuJNBP7Tru1NqnP1qkuDq8KLxd4zySPB7lAkEkRRjTcBOlSVu
E+OONrb4UDjRiABe9x3KR5pdDyChv6HMOLchcO4StARdHM8NRySAWEkwCIkhu/uy3WbT8ytAivG+
wFg9F2vUGhdplQQESacmJaP1eUMmp6HLvGikwKrlMziZnqE0XywrBuuaEvwbji8L45KI0XV7YP4P
5divig/YyijDr1s86iAUMBqzua2zJ9tEjqvtGiEegTig+uxHjPDlCbXpKck5fgitUMJuBDurnU97
AmPWXzchj/XrMxfDYXYWQBTEJI6nXbtVrIH08JYRvoKqZ9Qzx9JLBdva/5XjYEEGHlNxb/ao4Ose
BlXW6fHI4OfO+p2uPy7+NcYP3kYvSuHb5V3dagNItMdL4lkNA70W6wgona5Dm+IYH0xEYdzrbSHF
vx5DfFQ+7Rh1LxUUGVf8CAWKJMINMsOSpImjnOThxLOkCoAVnG9wkzFkx4GOFGCpIjs9D0rtk3R3
uhJdOmEkpF9ebNC+zeiLd445CXcZ1GDajCNipunHjNTdgIZdo9NGRnLDfvKyGmVmpbD/f9tWZLfs
ZrOpuz7ZElGKjVILBVwFKtGJdFwAuJWjDzezMSpA07uLVi44zyZD1AQG8STye2OcWd2OSzDxR8Lj
/fnem8+zGbu3+UGBhaTROrN7OVJBrjOjmzLzkN/uwhsvP353/EPifsVJQCVX5d942jCi4IETHPVE
LANoJzRGvXS5P7Z3kYFcIIsxb9AGs6/FquuRlnM8a05Iqm81+p7WD1anVkWZAODv2aJzsIVFPcF2
LuyXBQUbQC8RksJESJnaEAnO5yMpTrB4zcQ/jGcaxaWOI7iw41jXk0ue0kVK9oxGR01vXBeZLWaA
LqfenfKnyv3Mru1UiXuMCokNqTVz9rrAx2wu9yVmLwB56I022+mtj8Esxql+2LIIQ8ZGhGHDRvDS
95FlB2RQsWQKfNS4brZVFtLEkAmHo25o5hRhJi17s8ApdjiLICmZoEnqBzfFdcwN+rAuZbuhaVx6
XkoJjd64MCWLpb9nLDI2x+lZzZ9I0LtdJvuQ2ZTnEC1xj4DhulHAOHYYBb7SX33RchC3VKfPmNc+
EmRomxDrU4v1guBfGjJtbf1BDGZr0Ls0XiDkXEgefveaQHrdgPADhXDjxqqSfF9uimhJpGXs6E3P
6EFr3P4LSBLc0eD1D/MUD1qn4A/d4f4e/f1DoL1uGNE5wXeYnpdmgAgnoqTtc+J8O+sXNgPdEigK
KNGPtQWUPnnsU4KiIBn9Xj+ind4ay3sTY5B2l0qmgq9/V/UulgmZLQb+KWtjgzyGTKRgFAIAUpUF
lqKwIaCsUMc9X9KnV0M16UdqecTBTpliEOH7UqjXIAx0c39AvYqdkFvKlDR6yhuozav4nroDgJzG
+0z6pyyreKf+By2WS8R90wnJE2KfcSIY8Zf34MxM6QsArEKUVnDhkHLnIBa7H4jul1ZKANBaVfL4
X6b5FO46RQiSsjcOPis2bhp60Qo5+03vnzHuSVfYSuk/pOPOIGn5zehoAW5mGkf6uRL9oPPRSb7R
o//HEVYRhe0XjjQh0ipaU/zVtG2oaEP5DWIF5psmT5jln/levAhY7ddASjUqpbTfLqFBhHzOZdJo
lumupSpxlobJDTAELtRiidJEgpxEVdOd3fXN9N9imEeW43ks7EmUDtgol95qw0Q+EsHxcoGKHwM1
acnpm4Zvkafz5HDsCmxFUrY/EXxEIHYYjb+ctExOF8kDsPZtlhqRJOtUzIkiSV1q3w6lJcJGiFge
isPxqXjWJEJVnyf+3PW7lUmFpEnmCIlZ82r9l84p50QLkbZ8rcKLoqIrqx11Qo5mcQz+Pf6AYjnj
I+j8abZ6bA5Una2YQSVukyzJJfCLfuurluflxoqKAoBAHfsnBpcMwLCwYDFn45elg/l2Kng7p/Al
mnstbh94v3VbFuBe66MIUjJqX9ciazKremDLT6ydRJGhhxgbUA4+eIlScaY8DEUXc8wB7/LxNZ0T
zbRaV3OqGuvbzRZJgrdcR+9qtU0jlfZymVesWWM5bEOJE161iCmn38TmO26YQQqnLVzPEq8RHVcH
gi116qPzGILbMoouanyZSUTnuTigPjFbpuMak6Z1t/6IUHHjF4vNVAAyvjed9r+NNaUOMCu04f2x
Y1VbqwWHa+qiJ207pz0Vc84mcNmWfP9EcE5+rV4EUSrpEaV9DgM8qzCACj/eXqj3OxiksFeeZGIc
/5MCrgcw6UblMTupcyLSJo2ZTS0OFeoMjqR8knYsNpNQoPAFAXvsDDoHksFKrfvMxvVN4enMqThY
cxwDDBzZPZXKkvHB2y+k4EseJYb5Pt3phLzjmDy9Ltlso73VMiLo0PGJRX93EDn0inN8heBIaAKg
ef9FKL/ZRSexaf0graPE7FeneKGKeXuldLaaTFNTqidDKZuVhzXA1T0B6LNTKV2dA/YTto5sKF0y
t9nwpZli5qLlc7N+DcgH7/gGYSjqoPQ/xKiGzSObSB/ktyMCirJ0HV7cPSy9OVx4r0MCHJRoINNH
RN22cLsCcjtJhpG7VdfiaoQHQwzMuaO4waghLlwp+e2qqSuBcVe/WqfMCwk9vcXqtiKTMDozsG6a
c1BzIaNy5mRya7DP13oeydknN9UV1U5XXrftvgStVMV+NHPg0tCq8/0ZQhaWKEMsCFryzYUCDP6O
+741uX2DeQEjZeiil0XNHz0l54WYFWIjrXX7DTIGjcChM/pXrUP6ZcbiM5mYCTc1CT+IcpMwfXoI
LOHNEhVZuLVqcISOP0XHqZnj7OkgrZjSSZtBz6lU21Y3neq57jcIao/Qk7zY3VTMANi5klLjNpw1
e/o2LYqD6O2/aDEGaxnN/8UZ7A6EAQ4MGJVi9wUZA3w2f/PbVT8AB5Vb7UzekV/TnRWno+KiFe5b
3G1/AEaCjodQo8c+aB0KuWuCq7QbvBOfp+YW8RsgS0byMq/pp3z3SPJr/rfWnn8fu/OQI1n2/DEZ
W9Q9xxwU0RPsGm2dFSB0SCC1FKqOGLeX0E60uyLDvGOEw+IgEqi+Vma/Mp7J9/UKDqxSZLvKHS5n
rcT4T7mxIFAlszeIOfQsPh10VJ45PNxXAzEShZ2ppJ3s6ZqgbXcYXcdX8M0i6Ar4iPI9Nu3o3Gvk
GcOohRRrlMU70N5+576F3WOSHD2lPQP4yQ76tCjEpGJta8cZO2s47zbUldqH5plvI+NjG5n2G3sf
ceP4DwI9woHv18udqIJ1CjcVt6O1Qdsn95XGh6QU0tg2HefIFGL03pR3Ge3XbF6h/1Ochm+3Mq+X
R90ZJ6scAY/qtNRVdUcZiU/dvNEPhGoDpAtZ3LLkva9F7WXIE5mglYQVfCnEkKMl6BQFuYuCP12w
OAQe2+ROlyzNwGYCKBrSxFl47wu7B5juOUPw4PELsUILObjx9VLUBSFcvNnad0p8+9UNeu/1Lnz2
JnkN3XPMOGKwAJ2LG/cOkaoIgMVMM0NFla+tDrEDNS2tNFu7niNNd9LWOQHJeWS5BWiAUw2F4Bvp
2VZ8F/3/quVQ0nQqEj9e/JpQPj2kqKNSVG6iDZ2+UzCGxK1gvC4CxO7siHl1E2ARQYA2OIevJFo7
x8zct7Tip2tI3emep7zzO33xl74n5ic1Yqcc2nVWSiTZYPGi3li5Lww7BnTAsELOZKb5myKR9iwU
l2Wa1oAH2X+EdRTTyMkrbulW4ldqtsKCEOwKtDW+A6BeYNMMIXtpOdWjPVidIsouYshkV1KRcc7z
rP9wPHV0AFKmYB+h1oc4hgkFoaWLCHICIZUcS3BqtafAFV3c6iqfMvsA7ccSId5B59tEEW32mTdA
Zrpjjyeig+SMDFSRZWntafEGz7NnyYSPNB/5ap5HuMJwb1ORo4QJIdE3sDY+uEv/CV+beGdobeg8
cgtis97yjS0+4JaRbjY4Y6PSmS8yuzgRIARIYpqloeB4TzSC4xCTaQjuKXxU3NsEwznePcKarsQZ
s06ZWtnCzPfBtmGYhDhHZZFLU5FPK6Rdv6sDA86vzDw8POXWBS62rcY2AeLP/TQVAUSsR6WAKqso
h5g+QYvuVzwXx+9X0X083048V9txEF6oNisFcZulT1YFsPMFL1M4X+bOUCAMcfJf/iMczruxEJKt
UiL/6A45qrL8xXac5+tWr/bry0R4M/XPNskXUncULxzeHcc9mmhOm4v+KnKd/MYhP9MfxM8EC/gI
4ZCHlxxJZ1iSK+gBcsdqaYEqysKl/QKidCjGMVxLEv8oM0QFlsvZLlcEYJwlAY7pRJAjNK0n/hVg
Q9zZaY4c20hEDORb2TGukKHPYYuQyjbg3gO8hro0pScgZoj2hChqyWVf7oODHC+Ld9wy+4/vHTey
5tXHYZMR0BCUKq2JlmeJYDAE3RicvkMkH/l16s0fOrJzCKf/RPpGP7bYviiLRC1hdNUuV2/KTVgF
u5GYb25AZ0alnDjNNZ8GbSeDD0qKlfKKFjuZdpU9/3UVV9Zc+U32t8WCLhhJ2Bab73SPLwa4rcGW
9k2AonZKyVB6GcrNrEyAV3oV8efhqLj50GNgbo1971HuhOyuWM8Z/sb5iwQ8f4hYX/WActb6QRPI
37D/ScOf5DlpFSHl/MlGVG7nfG9cHAstj97s4b9yKNSMjjIvdfaL69IUoCBDKIPGTW+hc0iXz4AP
/pJs51IwHwQEGlG5a3FlxPB9uWud3EMmi1EJbhEi1ZtQGkxW8ci3J4i47n6uaKnNhG6GlqQtknQo
xK8FXgykz060gFpoR5KyF2lCc+Mxyc2Ah44VJ/Z25aP3EId9XPZ3ArjYCBixub/gktf8jC3sKS9N
X4FkQhUtwXUDLD4hiAN36WzqTled9ZMNdXFyo4MTQ1KLrPCigsWY4bHrfYfqMs8gM4YKO1REV642
FCxl1jBMoSQNhNl8YBdpSK/RTqbK1WFN5cU0z96DOzFtTj84utE783zMwONWeLngoVZSICY+fUC4
+DP05MzNiytvM9SnAB5jTdfDBf6LwlH/5OAUXqxVcXJ5E7O6yY1iAS0DSVHTX1c7QvF+ghhbsyV7
RAFogEeqEChLvsuXSmlR7XaPyq4KxMm51eI8LEEX5J++13NRuvE24Z2vDMlBUFG4IAb+sikRw+p+
YqGNNmr5c0+pZttUrIL127xZmwKB+ZURIYR/utoxL9IDc7UX/eLl9RrmL/WJFncNfxb5D+EUTxok
6odPrivE2AFhwyh6wASOhnkz6wjae1TEWcqvsiAXM4Ji2guLiodBgbt7yGRKbpcuWs5GparZjHET
Ao6UTKQF2bThSDca3XGqW12dAluDg1OxIJnp1MCULYBG/68S0GBV9iO0lD3/0yTKwx01WMca+s2y
+AdnwGTlGijOlk4zewAuItvGAYnridvYhhYXkLIjiQ6loQG6OKg3nT/VC0K7TWkqlj5GLvcfJ3Vg
ZLKcueRKSKWbV8pulO3zS5Xn3B8s3P1aQsqQMBF0YEmhR7E9Iq29Xi6BAHEjz84zOc8HNw3bBsYj
KIJ9ha8nBD46yl+GTphqaaiQKkKxdBlGlVwbjJmLu/EC2trUEqs4t7YUCpmNHGvjTayDFQjuzNU2
I+pbdqLjRgI3sT6fqCf7Zzj7pATN1KLjPTmE9wvYc8gz4zKOuhsF7ARCMsDc21+BkRKfXkEPh7wX
2p/+fdTnxrPHHZegFKrLun8qz07E9cViR8oksJI6ps/ex9tSLoGb2z4LMno6L4wJk4qdyp2OGS+L
PR4+X0gHmh4Mji2B9riQSdcJmNtxSJZTN/+KOuttmSwvi/d7uiMCmjNrAXTUI7sv9sJODsU0l7Rk
ndYjl7T5Z436zC1jxwahz+sT2WnQEncozAopRDLson5GMu37J1r0wSRJPB1AMrLZ4tcNdZmhlBBe
vaNt7Z7cbM2sATF2fuT22mHlCyA4ZFDAhSCBF/M432smKptlDoQ107SBKDbJTuuLfmqcMfWKdIjl
2ShdqF7JUmIk/tjWWXygJNgp0kxrX/kUoa7Mzp//Dmvm/ghyeOjFLJqEDz/Lv62PJYc3rymcxU74
NN7xZPBW5ffMSvG0T5XT8DwE4SJuPtfXBmV2bVCHqmzbicB/icgvVTEsKLZkjsPdFTW9wuQ/t5Z5
+kM/eCP9G2uLWzB04dY5SfrfzbjZ0fvk0HwCc+WEGQx1xMqlEkukJkCOXgeUIxaklcnJDrIqYM1E
lX5wwqcRAHFVxoYCYiyMKIa16SC8GVLU7HSr2I3TzbJ1I4qHosiXz6PCPGBh2o1vQjKn9xn5vTng
S3OBQ0wWT7OWft1yPcq4zPdakocPfhsy+aYy+ZNHUzT8DmU/4jr0H0EliYcTcy0N9fYxLv88R7UI
oEq9LLrdwLZi7FbpC2LIZz9c0fG7F6vZAhlVuDrnV6ZqudaxHM21kQl9gmgGg9Dv4dbCKcjkm29D
zQmo5jEy8WB2zt3s50dkj8fp2bRSmaWV8b67qBsgnR8vHfbQlWSWTnT3i63Q8yUdowsWSLcVI2Eh
zw5TiJ8yUd1iCJQoX6yXc39diRGSJrztW2XKUMMeutBbjXa9yb96p/WcdD7aF1f8R9c+kv74I9Iz
bXFj357iywfH8SZ2k79Sfgn4a7AFgUBn+hODWJ7G0jAdVMhsuivF1C1Oply8o7e8wUmiBytjPVzg
ol57/qhHcbSp8xS9m7Mbq9Eu+5ldq/I91Sec0XFao/Kmk6KVc4SsDQx2LHL/vJffakyiZzuP3KVQ
7WyXyA2XWeYSs4Fa88CdjU+dD4sHg0d22bid/Eo5tV+cOL7j6cpoUrE+W7XCwLfXjy81FC6d7+iC
S4U0VvsIq/ldyXM8NggSjwUsHFjmQZECgMrrhlPFH8MAszGNsod/gnB9LHgSCS10B8np5BvhTOmw
7DrfmXiwCY1KCl9TrjGiF9f5VnYKDSCmCc5INCsgpqVzJpZ2Gr2QaADMXTS/SYKgWbiv8ro6HuTG
fXeGQhxPj4BvRWXulkcquUAm1EvynmWeWiuYADyzrS0QktXBOPiNNoIe2wE9mipCVvONlLUnkfYD
FReAgj0+ybfOE6LGrdbm9Dez7kwXHRmo3vE+5c+vcVi1EW3zFmZO+3BWdeV+cYF4YVvgEgpIfcrd
lpkJpoaLk3OeRS33dyqO0CO+ZOaFAt+xebE9Cs5Q+sKgFfuL5fTaVu1TvNd69JkuI9od2x7nJlKQ
Xq2ej1PTtuQw46ibBNk34LNEKnDXHkLTtzXcUxlHjN05SvBUTZNg/WyA8ZL4BXB2311mHvpUZsHz
KmKajNG8cM61lvlsDh/83CqKdVOWuGSgyEy3P7PfavJvy2Mpbxaw7zOdS/8wXuleBnTC832Wq8dn
FjvII5Xw8niz/ac5mr0bRXnt62b6NJcwCDStpZ7u7pc6Y4LcnY1qYcQ08xG6PhXLUF94n+OD5XAn
/BG5UFEB1TODUg4nI3f2sSSVEROuo4gMJoGdVtUayfVTJdeopl/58T4DWf2ZCv0vCCABiiD5joaw
KIUmw113Rt+4NW+DRiag7riuMAgbe4SxV9jMfyV+YRBUdux0WcTT8gOt8jhAF5khr6K5YuUax9DV
LHk90fZVizRBmTgy8CO8EK9SYDccsxYIYKjeXO/roaEZZgG7mRz+zxaJPSRNIiBBW7uHg5hVyYvP
O76eKeeTCHi+azSI/sGso1wGGshrZQ0O2VqZDN4qExj1v0xJjIC0SaD1KWGneUC38tRfvj+9AVbs
AFyLnyEY826VrO/pROoKU9UG3k+bskHPqorpPHUUQzKelzvl5Cx7fhAJWW9Rujer4VrCvUHbN6bv
tw6xjuuPbXQLDsd3BoRmFHdIFi9qoo3v1Cxh8/4kf5UlmD8/guqeiq5Qd8v8rG5CqjlMR7+kUxfH
GiOgt2TVpMWCsBNztW2ijdZ70sgqJrdL0kEJQY8aFxgFBmIhPhB9XwF7p6UKg4gSLKa/clp3bxo0
ro9JF8mQpvMPa2UFj4opxridnxGPacM8HMaEjXUzlI4Hu5sifFlBiPXc6ynfvHHbT9e0J2zoFtK6
dFL94gZa9RYiLfubcRMyCMSG1OVqBTkY/X8wg2jrdkO6uht1/gRDqexhjrr2KF+XzfHjIJjHQIii
D699v/hP5jrHGq+Ru9rN/7CUC45rS1NSwRu9dGojP2v99pixf7kR5u3+ZuiGj0nHcN/zZaPbmCxN
E8EOUJFM20dllmiaX3ZydgylMhezTeKniXfJ9VR0cVugkynXGkoLRSkCFiMleLCZiJ1/ZKUNuLkF
LSgP0H6Nzj65vSvAKYpSxX4ZkBgIpHbguqpw/C/F7N2cvAVnMTQkpNMBj7ScduekNY2XPtZKdZz0
0XKwrN4ioTyVf9RC0mifBGbIFRONxelAgsBIYHbTMC8E5i9GaaXmIMb2Ok+P7IbTf92DkoSmYqRQ
tHRGBdo1VhKPakP9f20Jx4Fbj99WPAMXXDgdhhaBn/cs/0LCwCe3JZaAxEc+1o+A9LGFZJuR348v
X80xxQj+8Hf9cJLQjhwCKXRoM0LdQVFSTmL59y6PsExiTvGkJi93auOOWFMhN18dLxGZAhgBUlyj
KALilFS3vnM5k1TomYMxHtj5hjnXWQ58FjGe3kIz2KlKLoTSmFaTDp+ejsL8DB0KNuYN/RHMJSJ5
ehnWjqy1eCDNaUj5uhr42FY+tGYx3rCZj81yu++dnEsQUotMNuGDZaXA8n0eKBwJI/NJQdjDWVob
mLS/QNmM02bIgpF+HYkPOqQ1Vfdx/zvo2xQxhv2nAU9QLj+QAJxh4s2ecfXfOzzcKTFL5qERrCUY
S/ePihAndb1LcYshVoKlJRzC5eqnl+ean9QtWnCjH48OJOxwWk6Ngo8oA0rqxm5Py9ymnPS1Kc72
oSzFSEoTYaoZXi4PBOOka4keTEp0tlSQ4voLxCDZt1Q8r6+vnbxQrdz+QNVYUd6ftbGvLhCzdWsT
Jc88ePuko4ZePQCuDm/AyDeJpvAEesJctOTpOwcctcNo1EQ/a7T4L9QrusulMFvhX9iqn5Vy0dqm
OY3Ew8I+0MmCZZBv/UAFaUDTb1wYUbdL3kLgKFiYO/hVm8rMlCEGe24M9Uoi6pW8x5Wgs6Et8ZoT
onMfhaYxoKqagEQ4Waltx6t6ZJhoJRaJmOLHi4UEd+0Ds0b2g/5txP9VZaHr761k5hOhSrVf2/hd
th2AhPgTcwoeTeqbn/P9tbzJlIlCZp3d2WV2yQRdvBnQed7ZBV8lTGePV/vxQ0CBkcq3PRxo5xhC
nhOoigAhuZd7RaA5xEo3nbh9a9Jzb2j1xNSULo2P3T+xXj6mGBzxtTyWLy5gGnIWYtEClnhBqzMW
QE6W4P2twnxzoPum/PzOt2GwziMzot6P2Tk90K5xFD9i9MDxHrSbwS3A5eY/5k+fjcsbdMt2b9nf
m7jyMylEhx6ugX3JS0w/eo4HKCUSSnZCkffGkXoslrQgQzmVSbj7gKxG0oRGTgPEIvY3w4JAjQ2K
EJJOScZouObqqALb3Gfj2TUe2gt98rWoGw7w33otR2VfZJvI8LJ6QeJcS7zWMLFVhjiVdGkZnxaU
fvchlIrqsC35FrZbv6DatSLr7n27lgHsEyaYvmtgGPp8wSN2mGNtyh5ibAa6kc884k/MiFDgb72S
RkE0V1xbz6iwpaKL4N2mRBw6BQu7KycOybOA7xSnk56DBvwNpFKy2AdWu5dHS0hA6fofyP+yIOwF
6uNGs2dw1+kEwCwVs2PBFpkURc8ktX8RxVOatkUNLvZTIIBqjhw5DvLS80lGr4Cd83CHWC28nH2O
/r8p/m0JlzYLtcTAC4xkWFI96l7IXgGbrkMe3KZA3Uig6pOZ44P2GWaKO4grEgVcPZgVOrmdp8Dl
hLXjkzN63wnLxeG/jWLbzoiGBtITKkXncddpam9tdRH7CS1BoxY59J7EhzsMEFy4P61QzmNTfqxJ
ujWACj+BEbmctT7Lhu6VVyo/By/jPrtJ4PjYz4vgqLtA4/bDUyVUfLi0oRxBT1Bw94Vc6gcT8L30
XR5fqca/JagGOyt0k0D51FgR7jYXNTEr3Jz4ddbA36WsALdZggE+qAo48vNgtNdd0uFlfs5YUJWA
ctcO1Jkp20KwI23/9r6yyy9Hi0zZCoCZEsSCjXSVJ2+ke76O0S/lcY2yIBl6AVGb5DIJ9RbPRGIL
EwnXuA+/vA913R1IAoUrzCeMAKC06ttWIryph9FolSXS3bRCUUFycUt5TnAxm4gcj8IFmgq509o8
RKNGz9DadVfnZ1G6SaeTJJTY92sh7QkSQJRKj3k/W5hyHMjmjyXItwpAeNhZ9e3+N//8pN+z8rtu
Lsy6b5PYINdrsedNTC3i+x2ELp7Ij0ZXeozsLq5vYWTzpwr7M60P5nJcK4rhQ9ODp5esBsATHWTS
1Z9l385+U7mSA7OOsIdfRFSHTnDq6RNJPSU5i5HWgQXmTWL1mSzaZExiGP/Sr1fLL9IXx33SvcsC
oYiI0Zo8LYHfZBlqsQoi9MXtM5zxqia2ue3wTmUTsv58yY7Vk5kQJfGSHaZIU8iU412AUotYMVmy
hk0cfXfWaAm8FwODtg80St3iKZG3mgyNgYF1zGFGGGDOwj9/etBsvE6EsVpbHJmsBOnm8GpbQXXO
k36LyUGzxRx1MSj/88llSjQUoOrfdKWbteRjAP4cnoKZE1D6++Qa/Woy1XcyRQhSbXwe/pTzzg3U
WQyEbU/4KUsZhrvA0mKcwuVR3dADojAWUxSqDxTyQY04Q54LsHtIcIEcDgDs8NPY4DGuZifGRhMY
DPEiwMpUaOAM7YNlOqX8JHgiFhbFkFhtHx2vJDT17qPIez44nc2LieJ5uYUBP+x9o8Dr85whG+10
VcQXxYLgRZ7IUC/WMtHwFLJkOnKGFRqJavcIpFMNQpIuncPUR2v9c76oJtxhKNmXiatMvWBlfHNT
/wSyb3cOc2P2d1lsXPPxVC495RTMfXpCUcpM0h6WSfCxhyo3ADLw2FE1iYHLgRw+CPZ9Tx6tixmv
42eFleEyUaYVaju2P7yuvfbO6BJF3aucVn2UePjiOK5Jnfnnpq2GExbbsWA49k/cRsz/bRRI+Kc4
y8JC1tavr1lW5Jg4SHKR9g4sDIGzCgchM3r7+ej4bY3Nw2Ao6eekMLOItYmfQqz+0GNIek0W897u
6JWvChBamwcekNtJSdw1WUeS00lI36U/ExyLwJcJyxY6HbHvQfxEw7BJffSvdCymUh/wD39C/2Wb
bekRoYnijWrVgYuGPqPFSwVgixO04B19/BD+F1v/xn+heenkkiQfDl1oAOfbErpVB+6wjj8oSbLn
gTXFbZpa+ciejXKUbFRwfBM5XoTuWNOcq8oJPvyjL4RFQmlGZ4wRh0FuPEmJr6Mn5rZ0cjkb9kgB
bnpxcsNozNNwT5ZqJKJ/M0hWGgfJ1W29AJSMfVfvEvOGOzG04Jwv8fze4t0Ek3APsXAZOe27mvNW
bHZHMTuC7Jvi8dIML6lb5WyxJ2Ob2XcBH8bGF6vop2KaiCDIZbEHGQja0dYUjr66XrwuY5vwwc9P
MoyNZuzhnOBbQlIL7FvvRIcfCDA2ZCjg8nxUVtKD4c3Lf8S0uIh45OQDMx4BRzzpJ9/Sizyqdt9q
QMZ3QsuzoNq2Jlmmi9uY3WaUCTlCgvbnU+INAjwB5HcvxZhazSPhYgj4V31fSMuhG5Qa0VFZXe8r
EGX5tOMSent/qYCfWOLkKeSzBStwDZzVghV9bof1no1rd0W2PT66TGcDN57rncVOibi7ANZ3dnEt
FLuxPrkF/3WqRgJlMTgc8ZykVeaD/vXT4zWf4T0xt444O/t7hEkrGuymdlhESiuhOusrU3PVqEys
4SRYk2dX67GbF3GaBJKns96vQHP27aoVBP4+B6CQsDkIJDgXnFe3lCQMOSY4pALgE8kJYeIubQoc
enevDwii4B8vf5fpozj2QcOszVJWYBt1310yr52X3OAaTxXCWCMJVdM3z4vGGXlq7YgzN3J05dbV
AI3MI6q4P5LdxjXU/USxD12nFzKpejRP/2vWrI3AE9yn2x2t8rQDcy6X5wZnAK3mLUYssYY/xPQm
c3eKytnFBsprGLmXuao4MGJ3MF3Uqq6KMkWWCBoksGultoheHtfzApU7I/jWxHxMYNrRLKlYfqWl
ovabW4kYNxy8e9TTwfqZJRZ90Zp7cTtzopKyl234z6ucLanw+nyZtlNBrqTuxRRPEausu8ciSL3y
OH+SmrQNStbzFf+ijOG4BnYdL0MiQMPk1iczgfiRpM9mRLSHbNCwpvZ1furQ+SuLOlOTLcdDZCbx
9GJamD3zNh8/0UWqInqNBp/Xp+lmd3xDDxZsH9muuyFTAGIFgNdH48dbyIN95cjM/nEzqLVFKcaq
0MRUmlU2xpn1WzluTDuhXNnqAHvNMCQc6PFIXircnPI0ozTFqQYF9DxvVnsgvowYt2g/x/hG/6yn
TqIyHwPha1LYh4BPETHTIWqFvZIX9Lyc4JzGAkBzP9+bYgbBFmkE1kBHFo0GzA10i70EdKIruDOf
duXLLW+eo97OQ7zS1zYPo9VbmKi1E2TXIfnoip9TLxm3ZxYx/gB+syyLmKk90MF1ATFzkbomMrVW
YHcZL8yBzsNDQHYnJ5c8q3MjoryYArvoJs7Y1Bq3H3V8sQoV9675EiNU2eYd2IRu7CGVGcjvHi6T
+YBp1EpR8IlgkJIEVZ/M2W9vOWSH9eZ5pnWc9faDKyvHx+dLYi5XxGNKvAayP092cif+ZdJ/gN9l
vmZ034vaAmIYlVGR4J5ak/o7W7+h/LYkSptHYSvSvpwHTqZ7glWupw6nxioRrTNdyrBUV3IpwS82
WeW7bYMYDz7j0eNuPr2o9rOkdrxChwdGQYWN+Q8YylWyGTyjrOv0VHRGiQkmNIbdXSfnIX8f8Mfn
WB+Vhe/snay9/PZoqs7vKWBITH16od2P+JtduzKZoneE+x5MiGIy0fRp26k5gpyVvJJyOsEkJ6qV
TxeULR8xwZAyDlQgmHxJFlatmPfS86EG9fV9i/i/FvBEaaYed5wa1DPAKSd2gzKC3VOfK9DENXkJ
dRywJ2NsM4GLxlK/W8/Y8B+JEUQ0mI3vgI+TEzoEWc6nCGRpLIW/TonUfw6PrO6A780JI7GcMPLH
aanydm58sh/sTmRQCJs1DbG5RkpnkTpnaUwGgNaHjJKPMOz0LLAoU4LlllJcfGwLhZFnMc16C5zW
4Kk9+lUg2yVQPY7AsGG56PuEbNm5By7+/gEnCALw8VJ/GRy5ReDrCIm03bkUd9bOzj3vaebvkrB/
48eEHFgWOt8vJ2AT/dEEI9D1im1Qr5B0aNbT6iBM0aqOaRtzF3n1mOR6mgXwD4lXu+aoxPBzrkbe
1bnSXKHQN7tPlfASKnEKDvQpeZJ4NMvCcLrbP/gIOSdv8hyrcucc7xxnnaC2qNp2jaIothc3bpi+
cQYDw0pgQFVbkVHYY5BnSOXF1quY8dYIad6hmEhAJW5I2x1Dc9rnP1/VPx+BG/14gc/ET66nVv64
6evwV/QHzFASFWKvWo5ihXqKQidCkE/afTA7T7W2Cq8+qqSTA4E7rp5HkQ56iBjvAcQ5GtDyjGSg
ih9ZSkPrxav/asZkeOD6sifbd5uv9WwhUr/V/a8ytTeth8iPI0rq5yxjw06M/FzGHxwcyJLwok4J
DUMUySKtY0PVRjdmAmkIyxJcp2ma4rzrG8aVPBJvDDEZ0T2XMe5aN5LM6TJSijBGsmAXbtfH7xty
j88bCAv3DcdH4KgfvaOhEZPs7J+w/szPpI36sYg4b46qhNfEndQTJs70zDRhvgABqrbx6lq5IjTw
D8DDskledOLPNM446zJHXBoZhV+w8I/sN0E9ALLrkKl18nZRbHO1+45AvJmRUtd9aczsqgOmOzMl
1DnqyAvXT5NcUMvyC1oCVJ1t4KalK0hCwiV9fx7q5fExFpEbCAr+YdRVq7IYmMXlqJP+0uevlYBS
NkW66t50TOAKBMNYSjlsgGGoxN4lHx+vMdx19MOOERP9oQJzLNYymxmXmo0q3lNxT+9P+CK9CUqX
Qx9JG+SISLHUFQT5iig5f/yyq+jQn5fiyVAyl8rq2PWzON/qF/v8dFMdil+EfF/dhM8i1RwljI5X
kyco5GrQky7KzYfekpyORw7m6cdDAEGVVHKym1KihfCv5rHC+7ttkG0jfdncNYfkV1VOEZNSptdK
2bN3rWmAZA6EK/okNUbq348voA4GpKNNntcu8sYADK3PL7yxVX/CcGOrhLCT+OXqQy7Okg+R7N/h
zu/Mq3yj6htooFK/qxDRixWx6ecwSvZ1Ok0xcdEIUNLc07/pUt+QhWKjXL6hYPDJVVKe2sSoOFod
UqNpN3YlEGTtYAvLceNrcSHfR5aVj+J06mmzC01oSUdBAtanKdS2DEASmrfItcIqX8j+Lq67N0cf
yFGsbrc/hFoa9FEa1fJJD+CWguSypNlqKzs7fChK5HbQ6N+2UxzTf5HIlP0pz+G8W37l3WUji9WJ
aNZJDOJM6xeeMnMQyVBj9QK4f+albNoXy0xKiOyIie8pZMXhI6OoDiP2ujuL6InvgA0SNqhWBxjo
9aIPpnhegDvF36kR0ZNlruODYiwCTp5+iOtzDmEjJn1UrgFOMqHMcwtWLv5bYhN8PdGH4bGJaHm/
LMjvyKe+Z3vlU61phVbw2boL8J8GXAOa7oNLn6sIMzluOjMh/vwoys4ziV9DExiTYl2CErU7rXjY
vMjm4ma0sXuaBERhTzntISnRmJWTSpVmmQA39MlnLwgA6AEpmGCsdvttzvq9o4JceYgBLs1Q5syI
RL7MPoE+H/zrKv/IpOHEctDtCdvQnla5nOv+cXwRqjT5mNns+QfxUQWQ98FfLkpostbAzG4wUK1W
j/anVA1zsPpL3CtaaN1f4DZJ3C4lOQPC4WzTwJhZ5OOuzX6g9/5DeaA9oGvmj4kr7kAsEm8VMjTq
6pNLdGqfKByUXDbnr8NsOAZcUQtX6Z3+cDs8DPEyAMk+WcoEZ4dyhgLojXtSuuzpj2ZH4iu2uDbt
CDLXp9JO2RrnpwNPdR6L51NpIG6xQlh0JZOinLtHDLhmAvnbfqadc4xX9qpzwsscLhynRNooEa4u
QENJbHILN6rIQ0U3AgaHED/+woYZNcxd66P60tqPBg2UVE+mN9wJOsGb6YqVvr25WkDzJewPGFiV
GY1bMB4F3xVLWnnXxzBl16kD5gUOtGzWrMQz7kBhHjns6D+GHzVpfUNCg+rHR0pg7PvDAOvWjzga
OrMeGM9hYZpeO9tgPF19x2dqBBELD66PIXyq/57H2Yb15v4NX0YIFqyuaSUuRDmPMGbzyTUIkZmV
SkAdiclFf3SrU5fwLmD5YTP1U7fXPlWWV33omRP2JRbBs9uH+frPqoxmKPFV7/Qe15DG9ZBIQfL5
iEvd73NnfnQDXh6kSG83MPokBzcGTjdWskz4aaaLtewUG3r6tSbxXGkQcTGANUqeQn9MkSdW8vKB
BMvbiOQqNb85ivPeR0XT4i7OFm2vPSnSIwzCFA73/g9I0HyzFrXLRF0ZmRajsfc2STEEB/LK0TVy
VTFal+uTSWdwkNmLDQz3V1E2RDk7yZqAPBF2T26CMELPh49YD2K/G/DL8mqevgBo+AKeEOrv21TS
395wc6QqyY8DAetf7jXwAvy8ugKrTqMsn24qAvyxuGW6CHeHpUvvE2gA6bWrGq9+atrVzmmSDc8S
+LbrohEazVB5EMfxoIVQLIZGBIC2BhlELjdS0qSs2rofMUyGLWkpSxLqs0vJEV6Io8vEMOTa/vcH
YRFnryEYGnIaYbqCiBy6Ek2muiRMQx9EVkvJt2GPjRd+rn8XAb2MAw1KCJCo1vljizQQVmypnZvk
CLNe/cv5gZhLijw+1byEdw/IyPhc7QjnuDjCOl1rKMymah/62fD3705iQ0BUOwurRDU0AIvRtCIm
eLYzfr1UglM649JvYU3CCCwBMdHsC/lCHTTGTvkiVAeeEgl09SqoHQ6H4994+Z/rTbwOl6SGzEAc
x+Bfudxhr9b3n+oT6+QQZv1Ad1qBZPeO58mIqOREC11AKTZreuXnPUazT8MzXkDWwEhUqDlvmwYk
CbnFKZ/tQH7PdbcMpjmyrYuOkHuMNr9jDESVhHwGyQ8zjGEcohGQH1t67V3zY8iWfs9R44MHKIRy
YVCKFa5EOZTWrXmlzkWbz/91PKnqI98IIMo0iVHj8BX1PVdybN5PHupXsyJSQ0brXUtzLg4rUZdw
T91adt8vzCiPUZnYimEggk2S/RDlDmO+P83IHjUxTq9RSWWe2A+nU/23Do7gYPUUC8l6vtHLWf90
OgnJ+THpwqKPCRIJl4v8x89KGVF5dzK1flR89qBRYAm9ztWQu8rgTdb2s1GCYKvLETNPcIk4C4hW
XVYuXTco/Qw+TWqO71nRceLZwbPED/CtKsL8yQrMsh2nckNEL+i9SRHQgxv8UITarYZdjJSCd0U5
GecP0v9dVnYwBZ76P9qqluTuPz7IYRSeAlYgO1jvql9XTmbY+30VDHqzUEIczP+rRySXYw03ga8m
4i3Ps/A7ayMLB6J2Cc+4e+D8wnVIB6QVGYUZQkOP4KO9L8hiiIIfIJURkf4+uW/AEYqLdvDDhQKY
2YkAq0VlNPb1zd0OKmU+CHgYFJhJdb5/hoVNH3j3dDuEaD2h2MKBRNTurMFj8OhHQhs7y9tMVBS8
c9DdNiESY/vVFdiej+0RA6VIRVpAb850AEPD1c6qzd3sDALJhtTfpRWivyh6w2fuZ7/8CUYFYTy+
AsYF1ySIhj5oDSHuBdUCvGW+GKl4U3p5MXUDi8r45ZAjZlDYG78WO7GCsoz5TYpXgxgECqGXz2y6
5DgTwyrJUyQbM99hOLOr3Z2L5/H1k2P0LdAB5mkftFq/6ZgyS0/myC3aeE16LaLRgQd7yDiU7AcP
Mkypy7uxGqnyZ+5RsVHAk6RtJxgGR7BwIbUaXy6sB4yHfaY1drleCcIaD0RX2A82QIRvk1pD/S9D
ehVW3A2+iOyuVLw7jVndfnMKGBU5ALOjFI6CIM8zWaxCFZ5+HEe84XItKgx+SHIQWaF1Zln7pOxB
zIf9A53zZicnazvzA3glG3+ztOogPmvgL2pM/PqazkkIE0EsOjIcPccv9lGIX1dvLORWeZKpQEc2
j2mr58YEMp7BJNXh2lLAyOtThfOeB5LIRk4/XaDsaPoTM0we38u+acXyItBUbvbrSvQLx4RE96q3
frlCwbzXYWcVQpTMIZ8kRlQ1Kowvou1XhT6g+I+D/DjdEbP34D7bR48OvP1q5J3GyZJeKGhbkIm9
REthru8VUC0cEPMVnvQNGnjdQUXgq8aXfIUS7UNKTUhAINehvyJU6rrWZVzV1W/m0W3rBm8NIvTv
Wxyn4qFnOYw9D/CFYjLSTN7FVmOyUZIE+htEbq39L6DgGqpOaJP/LtIJCFpwWeQchOGf0nN42BEg
Tis+CanKN/S4ygbDOCqm7wPwMGWFWcwrHLvTESTQjnSn3tYIOh1NBSKMc0kP6w9vQQz8yy+3GvUg
4iBVVExu/Z1nR27qxuAYRRsBT4KcEbsDZkBx2JUv183S9v7Nv9/glrGznTHThqRsDyWify+DiuVI
FYHKm6keK1rINk6CMvN+Aot2eArKtcEMu0qFreJAs9+Tz/VFfP3Luh7HTf9foU7tb85qbEZC8sQX
lzB6w3bEvBpd79m6RE35IgT08ZD+2LF5IKCGB1d0vzSB7BKhW2Rky0HHDeFLpy5XDjtLf0cTKwAg
ayz8hBkc6/EM4TakVNMDcnimmRDVSSiryE49BtGGcXAQVXl6pXZtdwEHsmf55IN1iggRTZPQvdMQ
pPo2vusQ/X3cEYyTghXkmPg6OGvVhhE5YP1BS7RGo2WGvfBsFpitLy8yqD1zlNCCebIvDBddYmqM
70qvOwdohKFzsbtEDviKEDwQ5v3Hu0JMuXoViOvyyu/hREgd5tO2l2NE3byyP2noTprcuW9PK+Xr
uxUiw8JeQkifEjpeoaNsmxYLaYz7g5aXoPWu2c6eFcU0q+OoVtyl0uW1bMH0ZzYIUnmW9uvUtlTI
0lY6nj6/MXV0x05LYAKiCsetY8OaTlwWRc4OvfP9kcLH3IYeSQ6ZCukT+P/7p2EQEz2IC6mJpLmO
lSyy2q6BxgU6OYojCb2nrGgNyuXA+NjswMN2pM5Mpfx6Ij85RUKlPsfJznuSBh9BtPKGEi00Kuwf
EywXqvPzg3dH/2wtr2Eo42lxZz9JBAUBC8dHyMLKi9Zi13AMt3THh3J+Sm5gsFXkoIxCEw2IOJ7b
L1h+brro+KEHPY7gylhSYC1rYp52QmjRLYYB6N5v9FF11mi/1OgARnmGiaVfbHgoU9lsw9YYBYjn
knvEma9pV5AuurQIUhgWJ5jFnkDw2eQTi2FweBH+9Lbk49+FffcSFy+ince6MREMi+8rfZxh2qFF
2nn6rRN1z4Hn1BS5CADG+R78ECRZAQwysNZP/lDZNoponck6vPO3fBt2PHglUtoVlRw1Yb6vI2NN
2dmkPHcIqyEBsjnklL+yW3avYjTRzq7/qdSH2Sqm4X0VmXA87TH2cwFHJ/ZwrVjuH0vkg5J28ia7
FJtYPAW2E59yLqARm+shDgClNlKIZ+1rb0RzDXW/dIJGAEmF82jMAAujP4/ca9oe6jBWZSreT2Fy
TDKEoz/ugTXu44kvYaDAyGD8SxLHVuWKhaxPZMf4K1hMFhTRN5cJb7Aq8VkqD3yW1CZyJA9WRoyj
hiWlphYIifmvnll3cg4VOYx4ravlTlp4YWu2hIs4bGhW/bjDEt9MrcSrfOi1JL7FBOSCOPuBL8+Y
9WX2CbkbVOvCMrhMncKck5Ouusg/BkoJrnbD6wRkgOBQUNZba+idysW8P9PdVHU4GNs9isB8Oyv2
UdMxOW0oQj+H5KCK/1beeTdQclFPtfXfadwA6AbrRN6mo5vY8b23q6G3N3W6o7omTZIUNPpnqOe0
bJ2695LZFSTEpaaOmXHt6m0ruNx6aoe8TEGFirbOLspv+IvTM5TsOZIMqGIZMLlz6cGySW4o63t3
jsg9UyA0JMS4+k8HCy8OB8JOFpLDKQ1cS+w2xFXRA/i9PpDhZk13dedxs1ObNc44rNb8cjEiHwxo
N9vymAA3mOyZvH82/Pmufxb5reEdfKVk5NpNyk9B9kMwGTBoohVBEi8ZLoCscKi6fy1YHNbX9rfy
d90RAImJt/b/hy4waCEALoaR/UxIEko+0ZBH59FsnR+Bp9MmcbH9zm5meNy2GWrTU9wwUdva9F1e
ULcbFxDV9RAABcMo/psGUzQuqQafvjV4yI70uwhGbkwCx1zA23Xol7zMFbk8hyzYkVzpo8QXUhEZ
08Z03qNgoULv2vSH/j3CNT7cx5vrDrvkzYtzoj4R8dySfbEOTu1utNejW7W0aW1FM1cQY2919zII
gvXg5OWwyLN/4xoErLD2elVdtXJYv4lx0BSgMekb4smydYGHD6SgsVC6BCimWi6SFpC8wcJf6qYt
24edM+ATeNu81TQlVzzwHVXlUNkqmHn9tELAToBaSIBslI8Q8+Md1RnYtBc4hKbrBoCNPBr5ggrs
PZoiU2jJaPpsJ98JWsBUkQun8HPkTr4jjpt1BJmi7Z8UIWf//4bDYEGBea6snMrUEt19TN4BQ0Yr
pFm6NFwCcpb0G0VOR4awJprHzQ98Nv9HyuhLooHYZC75SYfrjBPQ/a8M7WPrV/ISOKYFs84iM0GT
DKw3Ug581aHQ0dvbdDaIpcnvrAxDTRokDwlv+OJorlaPOijeQWpxrmjcDIHPp9cfNcJutC3OFHaj
fYp0/5t3Zjxo0ezGOZWGrr9hMx7Gm3PZ2udMONVCkqVlvvT9+OXM2fdb/wgblDJdoP5AbkaNNNFu
nb0DR1SCwCdAcRa7qeEzSvN8pFGemx/MjwST+2N2tgde2WaQb3Wea7kGmjvg+9z8ypd9UuFsJdcG
1L65pTSStVUZESmtz61s4Xg5HXJv6GxIQK/RXwAGA8iNxQpDT05W/itqpRaxbyRDrhh0sD68sRFZ
cSZ22zpnysGzxyrO1UdyncP3dMQzu790yKOZNfmlLWKCkZLo6uRYnC7Thz3JB5m12ymBHnq+Bytk
v3uJiGagWMs/PxKHYgFG0pS/I5rWBXgpPBDNOdlNE6gW1rRA5QnSxB3Md5wNFvSJgAizYHXx1GSG
mx9lMgoNWv2pOESICZAyhT/KUFz4xC0vAebaVhjffE01M1dcoVLtby91j7JvtwSGJ6kilVFIb230
Mqg4vLLO1K9HxSg58/bLrYAAa03VijhmtSMLLGUOixcYnpx39FYmk2yITT15SNTae2s2KN7Z0SPB
S41Imc/kkSvlY/grVPkw2YKhSi/olcsytB8CGmC4TJ96tgwSgKGOHteucD+5vWR+62lRVV+CfAxr
KiFT6mI7FhHpT4FjeeaTZHRS4qIIl/4+HKCL5m7DgctZr3cnaBRUgBdGRVZFh3wQirP6Beh4ilHr
oDYqRdm1oAUE9vy46fVnoPnA41Pk0zm1DmX/ZgsEiHJoJsNf9bMibrV0HAfR/UqwdC1XAPDAjm+E
v69DNySmwcXD1UqMG18xfvp00MD3+gLuorgqViZYPx1xRPH5hVUn1B+4clhYHAwQkApNPT7JamIC
/Zsmz0KEHnAg3gLRFMk46m+/6J1sLNhZZVrPJFv9KQIHh8ZsT8B5+r3xYZeWXLV3nhXftbeELaBl
VmfjPi4vUCrcuQSaJhHpRY4pgEXyXIs8RG5UQ4LYcjAheTv8Savk97RMGPfmCBA/Cp9Cksp984oS
xP9Y8kc0U85odttD8rY6iS5Yo1QFcT2EZoG7qnWrbuLRgY2vVmP2tIFQXvb108X8ePYXJkib0sFs
0InvMixOXClJQVi+93c09JWiEAR+Yhb5n3tMFQM5Aktd6zxZiTeEgdeIsEatu1QFtUyYt4F5e7ca
ocgpnaaiiProXl/x9uyizB2e/Ll86IyQ/jltKzyz1jsBfYdAuoNMxjlBRGpeODaEq7p4c6u79R+T
bbA/OFHY0HtmR9g+YRaiIXGDHbnGgwBvJVFV8eHNAgeytUWIDuNL7KqaDoQ0hGZuhpu2RIkHQjaq
liPfSs8kiB1X5XDamgKG4eLcXMakzzKiI2BqMvp+Mwg2J9khRF7YZsPSX+QxW4YGcK+kzynmKN87
7pNPKlyh9l1mWnT9TSurpiEiBSLEcDGwSQpY2Ss6OrVUSFJDyX2Rg/71KhBaqR43cCWKjSW7FXiI
OTRCMl33HLDSDj/mX/cxPWCEoK6Td85R60rrui+vIBnBLwoOwpcp3buPrwf25GEZhvaNL+2QgD4W
4GIzEoFtYHVH4m3bmLGa+Li3Vdbc364f6j9SPIp93yBx+jIhVJScIFk+t1FPAZ5KGdufJfJDImS9
MeRtVAKJ7npx2vswFiKlJ5PCIqARGo4F3YQgsh2ej/4qfSXJrP7ahbVQN65jYcGPx+SqGT1x/Qq4
z2/lJOWkj6mBAf+7vLULASUQrRkM4g7SLeMil8DvedZqZacEhVdyC8BcU3o2BZYrAh1fssEBsTLs
uS2Wfxk4sVYjwu1UeXN8oy9F/0sUb91wMAFdMaOH9uPeNwhE4Ldm9LAq0jwLfZtm3SpufzLWzO3C
08mtAkzYZJD5aInOKRjBf0Vtq+s8T+wsg+bA1Xop7jqcOlQDUu00u7A/Dr+I2HEuYfg2FyLYoCUb
MuWj70WFyApUqXvhN/1HsisGxJNEGh2NapDqzYJQfc9wb1MqkGd89vCek/mRMLjuknWSaDi+EOg0
6R38DuNGVY+HR8HpsnGYgXWyBXY9AOfTs/8a7O9E9eKB+kUfwLxZV8MKZQdSbGt0gz4EOAs/WIuw
Ook+DrwhwmELQdmZdNakt02dRKsRMgb+tp459p6mwe+vHmf7JLv4QNrhsXwUNTvLMMqV4H1QZov3
XE+muHXW/CgfIEssORlsZbURdMq1NyYGq7D5BJ1PWnMyMcOgzAX3vMF+urRBCgOI+sDE/bVVDpx4
veib6Z6hWbmZ5ML+8hHFne+WzfLg+klZnWxMwYre0JQzKUt3JvqYwzvA2kPpg6UO5MEyAGzGO9CK
6KHSSxTXaBN59EKAUwshjKCzcLj9grJS2upR9PHJQR8Aoo5HeKjJOEwIVT+MA2JSts1Bwmt6peUg
dMVY/bp4UcP/hAAtf13uzawv+R6jjrrXz8gsM7kaEC04v87KtjQsnuafEKepspw/l19j75JoCgRy
ng/B0LIwWpSB4Q86VZO0FnQlfyyeZ4hBwAQ6Y7RcQFnU1wtTjEAuye/Ek61nAlQdIRSEzeXa5ki5
JT+RLhFKrCSsZ2TGhQvAeif+o2ukgS5LZEMIYreghVu8ZqPOSL7Aewsy+E7Yz6LsvCkvz7cEIjDf
1gZ9TJ9YIF7vF1MrAIwooSuMVA5CgNQaVMYHXYLMQ/lluBjRKTcqU7OOOBKjzn+Xn58Azp9uCOQK
7ivkVH4an8LiaPFHsHBNkBGrd02EsG0+PpCKBatQ8/B1OF0LhuyZ+xcFoYd1cqRU7EE4Kpr7Mdlp
JYZ4d0xNCLyQdLK4PIh/eewDYaJaXE0pMGRdDdsaIa/ofONMMPlCpRGBw757trTT3KfOYtwpcOa3
vd9o1YioCh9rBaWk1IgVtLpqedlDl0QpprkK8y/VNDJYgTAsWbesGF8dAxSxBnq2G3Qm1/XRir5S
jWfYtQoENoZ9sbpAvbAimMrkfCnGYG0vGdumSydfnYTKvfijs0p6NU8AuxXL5bIPKrE10rbUsKU8
6RLJhmytbfy0zaGB7NruivIGxxRhOgkXvtPCaOxGJuUJc0taN3e6914FwiNOHzX160pjcd7yN/xl
CBJDF21/JwIsACQzjh1qpxpBzic98VpaHEVwZoAy18bmmsYFvfWsOl3Uw3BJBTF9Bl4FQc1axcXz
lj7eganCbhDj0TGhsYfRcGXsgDq8TgpZbl2BrwnWtaigLLwur5Zsg5jN9OOwbd9V81IyxpYwu6Fi
qKnP2yASfiYELlLNzZlQ6xCYwrUeOJSjhuDP27h4uRoOyYJvwyDcLDMzVaHvJnW0bZ8a0k9bTzba
zRh2N7vr7vneKwR3LTpUqk5//Xkb4YSJZJAeyHA7loYDz7Fzs4FiEN069d894/NWKXAFNAIZuc//
+wy/V+SOcruVyqgQBhGe2VP1QPu+pN4VRqpnE2IW7tkGI5uGSqbqeG0gDIkrjhprTWjcuzwQpSEL
fBTXdMkRDq3S/4Sp+t1rHdax1rCNiwm5XrZ2UD6qh3ozPTBffJgIeO2oAFmknKNKwdLRg7zwfYSX
7gND9cGFpczCm+3klsbXwk9LthUbCxfl0vECsrsG8MLW2DUmerRhyHfZLW85WPSLaNUhTk4rwGTI
WUrd6Jw6NpPVRoz5VmBWX/aTE/XmD1iYdRAv/+0WLRy4aEcOFPLszRX4ZSN1F1Ixy30EqreLSd6d
slXVUE72cCeJ6XqPR1KYMcldJzbihxJtx5bbImudGIgS9iDHpJC+hX/uyzy1wfH24quLpqI665eS
Nh8ZKJ/FI8tWgL+3RUzrhFeisxKj9i92zlqQXzOxrLva8R6JNXQRi5E7/D4ypPEuOQKtjJ3dlnYP
PBcQZfPUvJJiAIfclz+zYltWFEe4ZvdSV/epJE+654fHw1PIzEK3Dymo1g6J6+HtRb0ZeoxNeb+j
hcDOOO9hk8+rpi54T6gHPl4wEBvvg000Yh6nVm0uEiLToJItOGPUPAwpjVmM83MFbiW3BPCnSPZ4
85Uxq4NTUqXI3pnIAfZmocz4aX98PfgI4VEFWl3fVif4i5k/6HEh1S+O2QhrC3HmLJpNjedxV/rJ
SxjATk/4MdX1hI2M42hzmPACoxjgdERNC5mJXGqydI0PzWyuO+VwViLTVbjoVwDKocIup9R298ck
52/i84aVKb29PD/hWwSW2/KrOtaWl3d2c6HqlMmlXaxZ9oDSIyaWURewKilUdRKZT8srcQtm9801
1WjauQJBbwSzfoAim84ALJNNO/Mia+UManX0Fxly/o32SkjLofgxGQDMxTWFNFUR1o61C2pIVTmT
2p6RLEuxEUEOLngSZjbCiwd45npoSTiWSG3vizcI2PpWAbidKpEYBDkol/2VA5U1CCbJvdyTRE47
THPmDJzl2F/3yHxQFSaGaXYpUymaDU3Wdrfcrh0vbWLJ2ncHOUslN+eZSPwyUHGl4MGwN+Zpw7P/
ZC+YhrOxVr8+CIU02L1xp0xsDkxr3vUdZD9dAZvXNg433/Ua5oyCkCHDkIJJQJ/NsiSYVYFS/szB
IXjkHhxohPAYC1uI0jyoX2t8fw68zqAOcoVTU4LYBmhgqk8Nv/hhD3Pe7FqSaQ57KlWaBxou6hTT
m1EV/y1u+D431AGria567qc4T1ToKP8ya7X5LFf9gRq5+YnjUSWSkp4oQH6cangRvgmxNpAt8jfT
QvbkRMsff8ry4C/Qv4xW7/YtJdHt5uAm0TaHDjDLhrQrZTX1muZkHvihQa18tzaMDsTmJX/bAeqW
aL8/qtRQUhovjmWIbOCp1tK5+cHWWZOyaApE9+rUGLk/HWzm7U/Q2lkzHpniLX1+R3cSjZT5zYl6
Yuxf0Lj5wauMc+s+MogXfquuzdqN/QT+RbmnwAXtNxeoSSSlumHiYDQk/JkgPGHG6t7UByBha1Ml
5bZMvonYBX8ebxfmXvLxiuEE93v63gesc5SBf/hX22O5cfGKU/eJiIuTqcYB17DU6wjXquliCmdA
BeKVepQBpcv4Ml7wNwciAhpssWpRjdEizRBB9vJkezKZ3KZ43nEkvhguDnvEVhBE0gpw8ln8vDRT
FTT2lkgO0CXyvHnvhbvEsWus8+/HIEGqlLpXf+5pLxnlbB77Zq4ajByV8cR4OZLtbDxWiYiJ+4gU
wbIFxzFdeLJn3Z/UE/eh9bceJiUHIRGTUQyZKOU5pIAeLvdL1QqbTaScGPLmTbn7n/TXqVj1HXWa
U9ZoEU22RpVQ6fPO/xhWZQSarC6VvBxDKA6N2h+S3MZym6oyZoleL5iofQIXJjKAlfcnUg5oq8Eh
hNZzFC24pFGfobaX0k0U9GPxgICDlPArYlevAnxgHEB1yoUBQUhoomD2bdMl5GIiaO/0BqDuOvoO
zmr08AtisKg84eiCpCODnMaZjPu7XjwtSxNXTTEeNqWko1ZRP/QGudFYEuh3/ZawhBVy5uWBdFHv
cDk6uk36S34G3rp3lMt+dRkXxiCvFdItxb0IDJYQyHWgNk9MVKt8EVisVWJEl+Hj3ocyHmaCtTa+
NIspmnm7Q+nq4F6s9984kD24jytnFdhaworW5oLEt307jpNqlRUo5ZLJfn6UIV99CHtivJRYwVe9
7Kg9lOOHG2bPOuMy+e9a/Y2Mpuu1+2EFV/jNLx9SCGHxd/aEPUJvSkWs+J9cwWxcPPvaakFEo/4e
HOS7sLxu97ap+kw0eaKEUW12OBoW2xHiQkb+rzifKNXeWoYvhvdIPk/ZwpsVyiBLzS+FKT9+R4h4
RJ27VCEiBvX2rIpxq13QVr7xqLhyc5ZKBNh+AH5TTJrX4e5b7VxaTwfbYEI7AGykPKFznAVsVmaq
lVwnpY7wcapjXMDAIZfMs+WI0ZLGOXR5tKDqr4fcc0rzbTfRGXOv086v2SEl44ab+ZQXv4ry7t3c
LdqZLKT9RcALWBxHz81NlMCLiYOVzgxBkracSo5d74QkGyPfmL/BNaGNaGRxxWAlnLpTY1O1iuaU
3Z2QeMM8g3lZ74NeN9OshWOawW1XGCxrCmCsZMFngc88EryJ2f19ZduqoKD3OwyncF0ouzxF+1GJ
2B3fNtnCnk2cwN5ak30rcmIv4vQVxMueGYhqx7j4MOdzKvaLyI5wgj60t2BxSCSxxbc0VL6t2woH
O+pz1LxgqtS1q+nsut6R02Mn6MGGcQY/jAFcdDKmzK6gxmNv9KXwMRXBQMKxoMDzIHLXDqcAlcWN
wwP2n7Kr884wV1pu9ndXP0rNq8YeQpkribEKVPWtopW0tbhT3Czv0QTIkCYEnxAOxpCqTfxC5vS9
tlgHUbv3FUCX1WYC+vZCtsbUkHmyy/sADPhaVQ47SdlSQWa7H7nvu6Q/cbKuVfx++ZelZVH5RT75
Xw+qLjtMWn7FEDr7+29qoQ+dizXD/DeJXdP5fYGLStDdQoie868rgneoIY4t+fiIpAKmJrwVXPgA
3gRHd5q6aYmSmSXCsBtpjYZPRBy7iYfm+EnQv6YqnBjJwqF+tEGRH8SUlE7lsevT6k3hNdtq5pzY
UmsFgxp7UPBTp/CyLeubua06S+n1n8adxhP1ff+w9skZEr5Th+N/biy6jvuqMsRsx6/v/2ZzFlmk
DTnsH24BVRPI2tuXw5fWLNIL4nN2waDR4YS2qt2gyRZWcSAKifYfCbvkTG/fSkaWtJ8S2RFO44OB
2xxPZg2dgaMi0SKsi+29DYOfvfKUuSgcPZsvhqjG+4egU7ueCeAmkZ8KuCgyIXjxkbN/iq1shzwy
bVfrrG/Xjzyx7LdnrCUmffwjyR7ON7iYWzSSSfxMft2aB+6GoVtBNPRQFkqXNqby05CrMDtXNhlu
RA6MlGHLXrdSPpwJ5v2EwF5h09J76tr83SzDVA2GsDB/Yg9ShNmCLdeqdtc4oZIULcQ+IkxdXnpU
q0Y2wxsCGs61GEDWEY1BHKbgl5sBldGpLyCbgp9YGV/V8rQPPe+zJyc4QFstjznnya/0j4yXLzWe
0k2dgDeq8O1c56VIYL0zt4sOKirIGYKNJrVopK3Y3sWTjkX9AqP228vvN0pSTy5CC4QGFaADaPWx
vci34xMVi1FgI1nEFPO+JV9KFZ95in6W1tpBzz/Tp7RkmH0vzp9WsaUh95ivmm9qFg9xiEAGvt6E
AUyFeSVkh9mxxU/OIympq1Yh87wIIozXHedIB38oASy4/jjEvuRJQEjYCF5gc5lTbscHbSDoThLO
1qopHuUy2uT5UqmscJrriVwaOFlu5IhMPFhvi76jZFemFWeJm/W2oF9y3aQeWyqfwIszpCKRS/AT
m+ydy31Gl9l4TUTyNn2yV7Qk+nnyTI3i2PtvxfwNKY9bnpcu1Uz772UjPQCGl5RaAtnfnyw0OTLK
1LuWkdywnlzvGPqRF3KdupEOfxFoPGk0/2pgYkAAcFPMZnMv/nuDqLdPblOJpQdgrPd/hYD+DIJj
aF6NGXmx2fIGMSDteyCyPYYF2+hujRQTmfvErlkCXR6iX+X7IY7o7PUuR8j9WCamfCXItXubzd3a
GSoLGK1K63PDxkiAdKPgoKmTo19QBTvRX+50ExVWAT29Q8pcWxMGeW1vc6asJSmrsA5WTi4/23SE
PjN/hgtJ2IK0/1bKkE3QQT4p1HQ/Uc7yDwsdwbzJuSW1u0urjJ5/xjatqgfdsgcOpzqj6GS49ESi
tMxq13Ckqe6mZrgphmo9jGzEuxtJ0nrFjESbnAb5pJwgFDx5CJ03C63Dwb3DapDxyUCo9iDTnwQL
Gb9Oal6CJA4cz1jZy6p5+eSsGiqWToee9BU5FczwoIyL8fIuTH+KjHcYhVvfyrZuCckZm/zSpYR9
scn78/T1GMFH89aWahpvivM8ptYGb5NQKaLFITCsuKXFunEmgIK73nh5QibYXI6a3yIG4vR6ZdIS
/0r69NGAcmMuWqWttDswUhdwvFN3UiorOWcdU2+lSoRSad+QtI9qiW8wNaT9A+PYPfDXCb1Cp2F3
XWiP56aUArKieH8F6reHF2kzuf9dlwkYhcqVHjlAh58I/jaFLaBplvni6widg489IHn0WgczVj++
E/DdYw1xSkDdkfQKcvvfCbfRMtdVhIUOB7DZYknas8MSxfrG8uf99cT2sJvocv70XR6vQ1xcgqvB
NLSTYM+8Lv/0u5BUQO4MwHlpF63hdGPw6pKo+I/d7b8Ry5xNlqFrkVgLqHiT/PFlWcpRJqx3Fx5m
5H+XRrWBJk7KLBIMk55wlzn3ygVeXMjAFaiiF0Rb+Yl+u9+jgKEnQ7Qi2KyRv8aWCDl8QltrvkmB
5+IxQ+X8pf74onffrnFsZX2/PrzAoQXUnC3Qz41akJvlWQI++M0o2MjiBdHEs1MKRCyIv2LBZGg9
ofc0f5k1kK2Tv/6brB9NOkwCoQlUsG/42p+9rJDwhDRdVAAj/zaDecc420gDocSxvveiTuncgp0R
VTxgsrki1rtYhmNfNZPB3745Wvbp63nY1Bp2PjlI0G2f0BoCBjJDJRg0dwEcsnmgbIE0rj1bGhpF
886wJrT1LJgS14w8o6x4vjxkZUVB5Dppsfeuq8pIW6UeuAMnFx67YldzeL3xyTEvqPMH99VroG04
1UNP4B6l8O3VsinRRz6GKwuspxdQz+Rnp56uW90+wt6/jxgj/F/eEytaqvgVtUyYSXSri+EB6SgI
0HunTUSRIkAXqjrzqiwDtVTJsoBLMomuPlPgZCZqmmgzL1LQUQhildVrCVOidzrTfzCa1hyCbcFs
bAcr1te5ZZfIsAVOci6STtFKeYL56y4AkGWsg0ajxwJjLNZ9SeGK778Ng+dwJHKNWFPa36WMdx1y
bu+W28tevQ2w4pp2SrUJmfpPAS6P9WLa5DKtAISyN5JSqPFxVBJE92ur4n5JawjZrTLJOHmCxeE/
8ybCeoa8LRZVcQBbE+H1JWxUT0b6+17YyUDny6tYEnoYmYTD6j3d3aKIS60ex7BuEr8lcEZfSIXv
j7I0eSZ5Qbepnsf2dyBEeauufBUvykzpRO89A/pndnimoS+cA8keTWdvCmzXM3iM1/VCyjXdHveX
3UfLVYigsroQ3LthhfOb+7CNhgGA3ExIDvSKyDyhE4Q0zmElH/8YeC6C7b7Q7exSVri7upKanyyC
cG3KP2sLtISltC+qFnV1ZvWNxjDfRD+pHe9hXeMnswHeAUlvcTndPcfQvLG7tc+0Vl+xZNp+yjSN
qEMR3cm/Xz5pvpfjjM3KTvNZMbEn96fvYQuIHy6VVlXMYJx09E3HwE4IzN1vav54gJw7hvagBqSn
oMBhIZeC5DYoryUy3PpbF1Sjo76AnYzw+APyRFC+sEUcny90L2kqq1SB7lWtbyd1mkZV3klVfz+c
DazSe+iMOewVyB2IUKaHghQ88quyfUeygZV2qBurRo1h76BjfMrdDysa0M0OO2G+Si3ja1eHBROa
VLnWVSHLVLU0JkuDsR7YvEuXYOhXZU/weHHUKhgjdD98AkSr4JnPiuGDa+rq/Qrt8OGCLxglyxMB
blua0ZSvK4y6EDaVKOedHo01hkO160nsvmax6hfqyuTBsCJDJH+SZ//QGLMcY9wQ+iVM/VF3TneC
DTL78GQPVHcKo545k+qAieqtHDBAXloRoGbQI5xs9Akbxb4kM+8s8UUv9WfybMTM8E1U/J0uomg+
4ZfPkDeAE6crm8iBfNe+itrbsbmQKhoXIk2IhBR3gWAi3qi8iWuIN3C29cz3v35X9JfM/ycj+YRk
zdOKm/bWtt/OIYL5JnvE1uS3TD5MOELrmFgdQpBVN+ig2Hh0rLo8J8KLu+sPUh2SZ/u3SwAUWTGu
zTk6qJ4PAhEhLoYytQav4geNDclKE7kuxNWdS6x+Yzo63beh1Tf+wurzEG48Bi0mmlWataFOgqNF
Vgp2cxcf+CZ9ai3Bqpc95N1vYjtzZYjS2OJoXD+mmw49+QEVWwrPEk+8vTvv4HlagSByvFlpU6ka
pEuxax7pO059yPBb5DsM2mxWjUPux9XsAoIvCP8WBG9GZt7NCvQu51Xxyj3uSPDOm1vBjEnqLjIl
1tR9zXDCJIdCQtrlbZ8SKZyjxW76Qn0hbHAp3RpgDAE2Jmd56Z4jZ1QWPFzRLP9uPfxKeRn9elaK
NNmLfZRLlPy7Gh/EbYC+y4IoVdJpHvj74OYdc9XDAoRgqwg1KqQRWEsH10bAjafjAVXyAKlOucpW
qeVaGhkt4vaIx8GRyySHtST1DKmkImv5KFSqMgZjOCfN5UXY66z2ODY6NCUW/RWuW5Cjn4jXw6wM
zzjIAadse9a7n7JkJn33X0Fy9fuEGi4HNOeSnblROJItsmv7hbcZu+LDOzzwY564JtEtvoZWQ2Sw
9KTHoaTMCEV0EEBWZc77v/BKHURxth1vkfEb6j0uekJgoUjgYet3waVEcgPgHsM9GcmdrgjRrpSk
CIbj7BIzv9emq3+r8ix5+uT63PbhdKuv087u/9Z0BW+gRSI3clIBa7h797QPuG5DLyw6uA9iSGrv
0fjoOA9g0/vSDSyGqCxFaKcOLE7Cj8dnoSvMITjkfHNJtWv++lbtBR3JqCWIORyFpcy77Oo0inz7
xrW7gQ8/tGu1AaFvFBimghpM1cnC89QXFvCzLw3QHapn7CtGaSwn1p5gFR3wqWdbiUjIQI4zDr9w
xRpbPv3z/VLnVBLnUABBlJ1+O0m/PeEOlJwhWpe1TWvcX5mhaGDHTjy1r3KjcQ5n4/sw+Ay06xto
ZNEqFHnQGnZ4dil4gQnpyxXwmUTgC5RvsQZa80LvAAS8H2sLEcc70aLrVun4UV3xx5PXuyff+++g
QgpS8H8SZ9iQVjsIwRCtvAYcb3C5AVd4a0Mh/d/qBipmzwbdxmUsyq/L6uGORD6lnHTuvfkpThSm
A8jHyKqmxunN27feKO4Y6NQuFcEM7n5GpMZnlfwKPUFC87Vf0AUYjJiwwYEKUmdwL6NMzQeC9UTj
vGPfKbaKve3Brz9tikkBqhimupb64Qd1fFCeco/CKn0x9MSyXDZc95veHzCnORuNyA8Sfti0RVGs
cavO5fVrPlGqIboaF9jwt8A+0fnw2zGL7BR050EKfrDqkm01UT8dkhao63e3K3p54WqkGHYr8GFy
jK3T0zHA3AulRT3ICYS2Rxxc0RFbuhY8BrKi9nMWqnPxiDNPlFOEItBDxDEwwMQveA9ltEMLuHNA
6tgTGif6x5jz2HDhK/RFRK9SYEyBwNMLqZEvKgpmXwcZc2QTfLPrf1FU1GUvSm27LyNTedaFq2HA
j0xylVNDyLosfqBG06+I6+YmhkZIUOh9IWfO4/RyMYm2QrV4yzQvXYveFgK2nsY731pAbtt3Vwsd
1GIzAyVak/xU3MdXXA1lz5/eu1UgX+3RYgKM11zAxlx+0K3DAoGEvNMr1dAlk/48kMaE4iTvv4xU
JJWLsDwTwZcKc56JZ6zZupO7kYUFPqMgOsaE+YCnRc5KSXOn1I5j/Opeunu6n+7vidGuGmXL0/ZO
w+dndiH/SMXOqmpEnr2X7hkeuEP42opQ3J2rRkCljS/69thayff5PijfrTL9M7sV9aqHU15nuu5f
rFEHQj0CpVmUMxbBjxBS10ExjQEDl5rujOs1GztXAjUbsXiX8O6YBQrN1PWtearuYVtD4WMIdYVT
6qJqCVzhcxl03rnWHSRKfG11c+soRozdY3xSdKHnD0qT49E5jjaW8TH+e8AcoDPaJXqH/VVTvrUh
XpnTpWSpBagNgj7NNbls4fPeNzvnvy+Fn5EiHcvyakSBnwNkOhm5dLBKjQjQQMWtycZN8eT7b4n+
wp0u4vBuYOmoeErhu88IDdTT1cB5QzMN9CncHFmwXbttO5ZUsAu3s0w9HLArBCbZHbhfdCfcULwX
qwVp5nct6pn2RYYRWgVX0jfHMmYTnQPUywaccHp66hW70yJarETl4fV493f4olTQITRANUrmV20q
I/3CapZrSG5Jd+LFnatrC38pHlqk3kxGRIq6nF1w2uCu/Trgt0mveHoj8ya601vNpmObMAVOZrJm
lXbJ3Qx9X/DW6boR+UNMbghrkjVKaYk0aRf80MF8b4NlvyI74DQ++jJY045lme2Q5Rz77OlnWwUO
g2hGcTr071IPSyC41uDYfjKqcQD5Guaup/jFddvumDjoiddqjFpaxtHDy5c96fjmPJFjZDhvgxZV
KDD7IUr4BPcQ1JQ/1y9bYJs029Bfn2CarAsnbQ2KZI4K/X7kPibI2Ga32QSdLwpEFNI8oakpfhYl
2p5dkgL+WbFAX3FmuKE+uHR/frPOyEr+HsW/ba/E2rqmkB8pKJkmqrTvWcTiwjssRcBmOM0I7B4E
WckfScqsawT9xkh1hkKhzbUPNv2GafYi1QTu/AlL/4xXH6Q+393WdKBt1MnA7v2EGVCO9x0NyZ7v
SNM1zO+fqgF9mK0yRnbgrmTC5zDxsNW7zfeA098P8B15PZnfIOXD5SmeNPJkJsfAZc7zYJprHW3Y
8ulAWIO33G8xDAC9WKmWvjuD3orB5FV5x0YCuRe8+9Tw7azI/THSeJXo2gRbIqIsmDMHrWPzXXs5
PCfSF3CZa6Bl3oXZhmg9x+iu2mdK9gyNUKCkm7ALlFB+6IR+RLiCTzqwr/XaKOZl57Bsn6lWcU90
mkqDdvati1gqXNOXKOoJxAj6JeWCm7qdSV7WMKPsT7lem5M18AWbLyUyk44L2QKQMmlMMowsZ1jQ
uSoCaiXbWx9iFqDwxlK/h7Q6niJ4qkLXTwZhg3iAWmNIHcRM6NIG2D1DK3JKHm5y38N7qvFhV3p4
B2EYuQ0WbY6EWFmcVDX0FD7Qte7a7+QB4C3DeJK33lXhjqmbivEID/RSjGmsLto9yQrV4blyG4lN
86eEflSJLARbkrZzait8ejwOLeZ0sdmY5gtbVhSxDUoNJOzCkWRoaBfLGxCq1GvwNh4g05sdnlmN
DEOPJrDyCsjONnUsx7hN3NXWRfQqaj/K9jmfR1SUVVfxpUpod3txnsDqJE9K3SPN8Y9TIlncsesc
hhEMrGzDA/sPg8PjRN31I6Z4u6Gh5NY1s5K/vy+uHMNpy265/a54k/ES8qJ0USWVysAi5V6MLizn
YJ35R1KAok1PsRX48rNbl1UCLdmnZQjghFzMssMs8VGWIMf7R20AMA/v2pU8KymADVfEP4AS2saJ
5dNbV58ojCQ5CbM7Fd6IacwHBQwTfObSvXcHBMC9dTFp40/jKMlIyYDPT4vbVXSZbJ7c8NG4tdt7
6maj4+Nzd5nfph426TCoMnezmis8XsmKeFm3YXfnjuSGwnsK8WWXpiwz4+sOxDPgjCpwN5CW7fyH
c9WZ4C7DPptyj6VW8Uohfd7PdMyza7VB9LCvVC/3KDGO7029AGvFyvJaAqV7vr1I5SeaJSNVNa9G
X3m8Mr8VNdrOUEaZys26pzQARhdyqCOouHuzquZhzuMaP/w/qYeW83vNrAhl20icu9RFLV4LyEEp
cAP5LFFKWMDj7X9FK/iEIThoXVTOkoC0brzSBWQn5uAoayqJ6CfugtLfuWWwnMbVueFwZAjmWy96
m9IYbD46LrjeSYa9v8CNL2iaqNHrwSWhjsWVOmjYypRJsIqF9us3XzuCSg/l30Pw5sOM9zJbti9I
vsTftGMfoPqvb5eh8QuyVT+sbHs6M/C/iurPFFV9lw7Jkc1A1FITRFmPPzXDfk6Ol9mxo0yldoRr
CT72bFL3rwd6mQC/Knlfjay0cfBTZxWejCvNYprd6l/eP9vuzQeGrE2P35VkMPZDbn8k0TPBtUKp
YsL8GM3gN6BIz5lU1wU6nfKUnSVK6ETJqw/JBkayGBDZgT6i/EaSWXMvov4POXCL029Zt1YIDhV5
IvlSGGVWPOGbNEpVRawGuS/ClZsTIRWw+AXForMqrlbhWui44QIcXGh8G2bATGHKhGmryv1Px5o+
ILo+gvhWqgzX7tY4JxFLBU5d6HyfywVdSrunjUZwcMhDhOh/1bTSJXuGofGS5ru0YMJe18+TQDgp
H8/5hC1wrYMmLTC5HWndATjAemWCwVgV1XbpfsilaPRT2GSLClMoJjsHcNMs5mUPSDZ6ebaVW+ca
MmU2hObvcIIyCBAxCPeneBB1uWhi/RPNoFHsAOQl9X7Tmwa971HFp9BQCbBp1IXv9ZecyDgOazcz
gbX2GuPpaPypiieIsQOBHEUw2xLQaYlOY38DvbArppt/zFdbrl4/doeUHuYNnm/uM8nsfyu74x27
v3XBJ3vxoV4OCY0dcwvZDSCCNKMuBzg+0twlXvZTaUl11DbX6zMarPBMc4X44GU/8sphRflQJUZ0
wGrkTI9B3+Ejh7WxdiD/QvQxb+C7BG7jN9H8fUoIxlRT9wzGQW+kc7Ub6scwrA+Eil8btN4o2dIs
Lw8URe6Fzj606bmywM40jPS8JSkx3diDSqxCmJYfpnI9dsXZlZPJzWycOGJhpKf/4FRof9Pdzz2i
17B7RvSuAxmmwg/ca3fnd55F6phd1HUPAy73Rl6x5GRWhujYuvIct0AtBX3TybxEKu+cWiLTqn9p
MI0D4M0is0fNbQE/0Pbk70j5KhS5F7ciyQjtp+5PBjWmVcWnX+qTlEYiXGkcR2OaHwXZ1AeOUwmm
RIxtbsYqwqWFYT4Yddl+T3HRwMN2J0prHlwnSCKMuiIhErFMzLugA74/KzeC4rikhVWK8M6m2UgG
DxF7qBD0yICpFSvsZYB7s/usWZLOJG/SQFt1Z9pDwabI027jCimhSFPmHUP3DXhj0QqSTPBX4Hh5
yzj3PFrHWgQ2h+6l1yRTEGxb+m1VMSLjuHDVSKq08yjlqgqjIlybBX5KHIy3aXV/MaI+MblgyExA
52WiXzk59nsOy8K0VV/pujSzmE22MIRtiMwgbF/EUfThKmRHAGEUwUnXow8Hlx4QQe3+3CSdlH8x
8XSeuhsCbyof46LufJB44wJyLJIaJ6yyPYi2szpkycyya5Fs1beBnHGwpkL5Ydl2FjQIqRrv5Sxp
KcyaFuyXLjiuY0huWE0rmQTuHUAsDN0h1LI4+AmySDacGuw0Bxro4+8JQYjXDgITDw6ADLny8lDG
UQmoCgsNP7b/NqxP93AXaggiOkA7hFIB+diW7YbsmRHR/gI162YhE6xOzl0dSdRFiD9xDN5p0y+W
SZoxDRzxaEc8WAdAofGBtOTKGkIC4iq9lige8GB0BGusBTs+ME/wn/bbCz2xiVvn5i03ejEUpz9N
xJppfzkDl+3QgVEJfvOoVRZqR0uz+K2pH6M9U33YGeyJseKiPAksx/l0vMs6mGIj983b8m5vf7kD
pxI+20VXNyB3299rHyzBqEUK8MV3Bk/WhRiBE/4Yv65rvUohX1E0jgNUReBFaEStyhO4SMguaH/D
k/tTsbBDPUiE1AQ1P8LDEDHky2jBxAdQFwpB/htW1xoIROIcNJrbWjwGelrpIJQXBUMUHnFzqVIX
XY3PImAGywNh8WjXAgx+j5m867pTivDtOWhP5jwk3/mX58HKNz/UqVIPyBi+K6NZvD0bQeXurWI1
eVP5zDzbbNsU7jidRvt8wUGac0mAj8cYjk3T2n65jF7Ou8p3gvgSl3tkUKw8dEN99J+1r1thIUOa
sUU+oRiVQJEh5X1amilJEQwiTnAIszVm3bMu5O3OjUhyrL9UgErTsazW96htu3zYoieWPwwM0Mz+
LXikgA3qN8qvnhwxco5HGtJtDDH6a675ivyxWdwXNLOhKbbSfuQCiUjXJVvsWMQ6BbKkESpRUxma
EdGE5X0eB/jw/Gy4bMMASS7Y5uj4+NHuV+D0IXKAJgD1f20hkivSyzsGl4R6b6pYaR9CZNjn2HAW
ORHEHbUpUjkS54nv3vuLC4sp+WXZAdkNZfO4Tt1afL6qIziHmsG4tBgQLhMlA5XVkSqiAgK08lnK
6e/NMu4QXr3NykZoQHsI9WL8KxK3cJ+mfuO40GF1MR03e8uEuFA5AxVNvU+4y7XsY1byvDq2OWZp
GZVTNLXz88gH95yXMAQm8uciGpVazzo7ovhRHs1SnHJo3TworYCFQo3v7JKFIcfnEap9UyD2SV8y
gOGCToShmBMguX4rNo2NP45COmrbsLSl4gMTJRRx3Fgyl0SLp9Jx29ax7A6TfCPBCI32/GYlSgn5
71xCi8kWKeZOt69KrpxEcw35E/R9vuh6qH3Q5usbJEF/SYDZ2mIAFS99u5Zba1jMyyz/bY3oWDBI
ercLgGyBOyEsSDJyKoPf10q3P9jfERPwWsbQA+JRUKh0BieZKjQMvgybCFjg9q8EsIva3p2oKFNZ
os2gr7PonIzbORMV17w7tHGY8Cqt4eKP5UCRA+nRS8ToI7MumpT406sB4KNZ0m0PdGeR+P/UhzpL
W+F+7Co4E21sCO8ittlW85gszrJEvTJuEgf/KGEOU5zpBme8XG9rPD1n54Psd6yQ2wPyVs/Av+DX
VTc0K+NGdJVOnU8KQJwYdD2z1tAvK2HNTvhcr5W1hGFXupEPQ7MxzckS8/aCE7ZyZKUWbCDKMFTe
teb/yeDbrq+nDsHP8GvaQKrnRS949hollB9n0tY8ZUbJNVTYb7GxodTTtskTmJlqlaOBu0srdl4K
nuzDC9PpL+lHuPgKncDqHtybkR+5T5hdyZXz2s6XkGZPttSfzJvvJ5mNMHgmkUO7+s8EcfEy7nHG
YVGv/bEeEOCpd87jqQ1wNdGn+nV61m1uL+xFFmDwWvyS8683A3rS6MqTV1saLNvq+V4kBZ7tuzjf
F2AVy7ABCeRcV/onWTqyRYU0JkraS7t5hNlRbmzgJJN1E8hC83+KzItxypbmSw9ITFRLwFvLUtqn
L7c03Fx6DhdBzz1unHMtaF9Vd3GXa8qA0UEFUBerm8onr+qXZ3s0Exc64+TKNGmCpHa+olejLPrv
cIUps98nm2c5W2YeqXhFmG1ZFlsipbHLn/jThlQQfRyIJiwqIRdBE29De4gPXUfj8RBTRLMbUoBx
TvISoKKofjfvxnnCOUbU/qqm3IwrafLBUY29PGQIcmVbzz0JP7vQtkbZb13USXVGV4o6CFHGikTw
BlHDukVZuELeozNmGuxZSVHKwYW4ZA5L/97L7snhVtJow3MDAm5+93teDcZhg/LsNOmm2LOVhqvN
1/u6+SO4HpVBCTYEM8QgdGV28yY4ZFIqGfHZKhiPXQTSuK6dj1uMirGP4Njo5jn2FNHWGegXh+bN
VsYNGPZSmbrjTedjwxNFtexvD/e0lKF9ITq66xPqo9Y16PmnmgHSvIujNFu9BsCbc4CXw473ktQP
Sd+BeoFTJ/WLY4C0D/IOLAQZ922+aewpzZUP5I/ZbH7OCPbT+k4UtckXAfPNHafjZ5tT2KTZBtF+
Dt04sh+0MbIi4BI2w+KRDpeVj6OXGAlCVSDfkfM8S5iOkn+PRUJ1+nvQz7XzqTTZlpWFjF1W4AvN
/s/117Hk/hwNMqMSQnHAyHVAMTprrE3X0Rw/KdBe1pI1g8sKQ+eH61jOcvjlDF2VgLKX6HBhiaja
TPHbqDfcduyTiROBhguk0ECx2+e6+dO6awfmfK+U7Q8Hg7l6QKnGGbR9Dh2Aam/JAu8qHCc8N2qq
zFSbgoCps/L84NFhoPrUTi0CIZrRUbguEcjMlEGU0P2SBYigHLnMY2KPeGxPGnmaOC/b4BjugnES
oMlKOAbdhN+INrg22mPfq9tS0MsQtnB1UivGjJr6mQn4BSSu+iMQp3Ty8hpoafashKQg1yCl7don
Y7Y0a+RdHZ8yfye1JFG3XkT7MTmeuTKyGJAEGFpuJ0Vn3AWsvGaSHcOgUsWCajhXKr+WFf2bjU3v
BvRW1jguxgN0yvzetKwLuoSTNHS+BWhvzFufPT3SCpxRNkiU5QGRR8nkanvEih4SpIzy0u022roI
07zYU3k/zEvNQBdQ+vnmzu7UWvIjXFX1+eL8d6K5PUtYwJ61x69BIG0ZumSW+hTnZTxsfwQQWHtc
gJCL0MNtG7JxXyXoQ6nyqmYuYQ9f16K+oP2LrHjdD3223HeZ+/rJuuPLZnNj/eR8Amh3FduJNYq8
4H3rD3LDLqo2y07+qQ1UzKWYO8tT7Lc8n1859p5natUNpGy5SenXNu0kRXTEDahSp6htFLQL6lZr
QjmFhgaHyCEcK7syL7RNuGDdGuCOlUQa1H0qfw/wZ2Pw4TcPBb4NHUZH7exFnDKId/AAKujrGSaz
JE6zDd6KpUE2lLt4Rm1MnnpIX6CLIKL2kWgLONg95bM0CrD/v1M++fD9GY/vCEs+59qqyeYEcgBA
eeSqtejOYBXgBhSUxmNWfX8/bI9T8RQwtv6vlf524ESLsvdzyzs1JRDjEInBywB7VfvV6pGb02Ck
cQ37h+k8xtHtLEnYpEPXcMX3mrgfRdFOYPvwDaXpp5ZGd/qTr/2bLWfl0uTvlEpltWDSk125+r2N
e61HKOvA/D6jJ1xi9hp/LZTLE73rf8dFmfROq9Em3eKy5dsueDjEgBOuc8rbtU4M86faHNCeaHqc
7um2aViuT1fTTkBhwg1HT+3Njw2wDSv4PjjXyC2bmIjcY5UEbvcvWJYGxlOzKpMd6xYtt+Zc1Xtm
2jVsJo8kZGKiUsu72eVqrLxtEVRcsQmmLMGMUlhUWaymF6HwMDOzCtJ2rPU2Gw9bNw+kjkKshKo2
NsqcXMXPhp1F5baR3Rq2pGHQxc8qqsocvRWyiq56DA3dyOPZk1siRGC2PY4Rk7vsGHnoZ81Do4/X
bhpdKFxrPB5zCOtbA6eDRrfMEFR9po60gIcxXIPbB54QpgxqO1EDpRLLwet3xeXD/9H9JlI29URS
ZOUuJsOvmlp224FOQXUTo0a/8tIiNzYFTITg4LO/LS9hGmywsqmyU4BAa6tC5TPBc9mwunrUPd/w
qiAPo1UqFfE/4ElHUXBRzcGECuELRZFKfLeYylYu3gwPXR7WiATLHC4UEL9txap48qR7MAby9WVV
Qqn7Mbj7KxiczBsLwu9kR0JZnlhjLDo2zA238TX3/vv1/K3MkQolgLW7j7gLkTz72dNuoN6JMbnv
lXZLOSZ/TkRdTjoZrZAHxo7zPPg5rGYUi4mEikzGdKRgy+VNaBvDtU5wjKIRtlBAY5E2N6KCVLC+
st79mqN4cBijYf/j6DQug/rDO9+wGwAYAIWGgBM48j26v7bT1BePbEKSDyGel0bnWpsFZlIxRmOj
/LyefbnoOOJwr/evA+Z8A3JQW4wm4WcsS/oLdzK/jqITF7TwOhxE309D+3cvejJi9Z0mi+RpaPCO
0YZ+CAxcLAFAtt+iwcpjjV91Axrd3RmR8us1s0hNdn1s2xHMv6uk6+N0UKrC5vX6/4S87XNEWZZt
vE+5zXzj/cM4GaZ5BQV4rROGxG9Fh5biiCXhPdrZ70r39FYw35JbTKE8DummZU2OghE7mssoriiX
dTejlbBJ7Dd/0td3mJ8sbIPIKtnxWINkJDI0zPHsBeAHlV8Xrg0Iel8wFp4DiKw3oxxdIlTOcGPJ
vnRs/oWhXSlm0HNG9+eUwdvq9fPOysZuBcFBhm2jrE0j3JPdTISeAWbEYRHHaV2IDO/UJQUalDrc
6nFtxdoCG6ZnpkYz9VNOvnsd22/NGVxw1KJS2PZ8mKFJ04WoQ1H2wNIR5q08emGsLIf8twreY4mD
S8Lfpth0IoW8c03jKQeZROkwuXRYWJDbkZ/xtFBEEVIKdljbmXOZdHDIE7pG1iuMGbzq04ErPo5X
Dw2ox0szvCTQTfy8sFAj73l8ZFg9haT5sO2YxcQ2DiLMK7PUSknD0GKtfTnnzR2G6AFx8cmzA1Bd
1eFIXU7UPunAOih3MOyjeiFTS/zFf68DcbdpwlvdL/b8twa6ciAGRhpGre5/dNnf9YJO9onbp5Pi
bT6nWTdVvFdBVMkcQlzM2Fkm077FJqF2qGstG7/UYadjiuHCiO4fhscjKG4gCKu3rKgzPCGFVk11
fA5jhC5tzFkbPt6a0Ms6vMAYTcq6o1UwyUUEay07moEqcg7mX1ia82j3/a0625clWr4U/1yG/tn5
KAeL8uIEy2L3tHaEtrN313uOjAo8sfMu31GOwUKOm8YGiMDOWfZPdSWt0ytvlTl9Wb5DrL+04wEM
RwVsIW4mDPjhuBOALOiunCCswgEv8gMmK4+QUretUy5MXRy2bJXMbhfJn7g0rLCiv/4o1QpjMnB9
PEBi4giscKmAl+7dnkVAIViHN/5brj5o/3hBZ1xZEa9UdixHxnXsI2M/cCgYsHKPNnSrMJoD/Och
CS49abd/Gp0L9zP4viwSVI+HaNAV+fE1MBIi/HO0vi9kmagqF8ihqF0to+bLGG3P+kvZMgKzGwFA
sMmzXv8O4/OmSXDbmKnGp6lSfYPnVgwYxKLrp/0U4/sBEygnjsUt5OJS5J1ekvYIhI/AHYpVIQSN
NGOoQIEJmcsdrEDu4+7ysiAlobU2L9T8wLDzrwM0+HKNygbpCymVyRxLtodKWr4CyDoPchC+1IoM
Oa5GI9qJ7fVP1xGWkBhBEl4DEw227gqIoJS6XUwLg0WQOqEXJqEgfkWcFx/cTmo8VwYTJXUuOKrJ
a94P2/MmzH449bzZh7UNmuVodbfg12EySnM7S0NcdvmrxONrCqW2+K835ZfVBOVAhlqM0nkFtQ6U
hlNXj98NfyGaKE0tsc628CcHBc2a8GUfOtfJbv6qN/XczTzi78UlK1mcNrXfLOt1BcHkbJKohrnX
UI+yBgMSqOHzVXKHtoxohLwd1I4vLisZZK562jWMnkfd5tXD9V8G4KQI5kxV+62v9Cuogt+f6Vpm
yiNarSA1UWg+LfHpQ7X7EtLDWjQa/JYEfsI8vvgru5hATPf3jdF39pM2w0NAi4tJU+A2fk2P6CDw
4hiHAG9ihjsbxv5NYD/qHNsAg+zs4Wu26nRQBWDfb3PIN6J76ej61JIJeCc01+yA9k3zXVnwNSuT
+wbpuXBPHDPmWP+N0x7ZlPAzT3XDYAaNmOBkpkuk95H7edGB5wDmYufjuN0mtu4/gfdm0hAOQXbO
2fM3ThnuUe98F/CUl9tk4eALJQt41CLcFtBq4mHXiz0wDhCJ0WBugD1HGF8J3UFTwtOd1BKwrkVr
Ozdh90kh7pSvHjKLBHZtimv2UI5E0+aoncbTFtQas8nvGbioFq0xH1UwipZofH0DdfqA1CiP8FXc
rkI6XYS1XjbsosbPtlVNForhDyln02ELfumfk6DOXQVRVptaP05IKbjXpTZwRClrrUt/sXi9kwph
sDna4LofURyTRm3E2oafvRMnuMtf2hLLXS7YqoXxemeLdpS/lNqbNb2JjHqxpklPKXVAeHlVoMM5
ZUYMQuSI33mO+coLhhwiBrnjTnNfGg7xVpt0wm0Pm06zELjKp3wM67JJ8EPeKxo1725sT2OjNydL
nsCKmkyYPgEvCNLmJOPqzv+pWoU3D9khfhq6H4XMebvAz7MEdOIm++BFGLNRv0KhO1SrHUHRS7cV
jQF2lWI/Wxr9hsajEkZ3zI59wnSTkRM0Qvr91WBC1+wwa9fVMZREetXRsH279m33v9HEZ6W5SujK
s/8CDvMRRZ8e+gy5frvGePdA8HSEo52RIZvYWgESNT7EO2abt/Qg+lHchNnD8I00w8pJloFKFO9u
DrCxp1y32CBp8DlxNIYwlZpGgV69192TR3OJWEwP4FJV1Iot+baHKjCdEEAgEhKjzpOlKOSuynUZ
/AL7VQa8FRqlVPUiyXpMLLiwCE5y4vlC0Rx9q4B0aIJrhBWMYHpdQGD+DtmuybKOpHfUWODPXG84
+7DLPiBAbAnTjkVRV5oGud+jCrKM5165zJpdsHowU7f+senyo+uDPmouoq9GM9sYggl1DZycb84g
7iMHc4ZlwSi3uqIsewR/T1NwGLz6/EtUawMucvcIr3t0U3AVOifvjw58M4deL1eQIWCDMN1Cq6YF
3tyro5yzWG9Kh3hIEKYbMeYCOBoj1UauiPa5Z+dXwqMycF6cKheUf9L7C61LbhyWkWKU31rVPId2
jA6MsCqCnv5zaNpzStBKSeG0Qs1p1Ndmy+Z8jxeLleuuHEenw4KE8vkDN4bxAoSRUSnDKASaCv7L
A5bxVSOpjIQeXLfXpG2CoQwMVhLTr1Wmj5wy6LegsTWkCSCh28EOieBSW3YjtHDzKnbOnqzM8FMZ
pfN6C/S6O7jypcqUOBoU9v6H1UtmrNzZtGund0hg3c889RB+CWhKGKPilT4ZNvJumRkqqG4HqaCe
lv3nWVvxu5SrFpg7f3YF7SD4CQybjrNZ17QVb+UD03UCWF082E+ZUauRo27q5r4p9FHlwUp6Z5ZN
abE7jWpsnT9NkULf1KO6VnV7C53zIkKx3mYTfIFxIYp5rPufEg36YBuuUxNH13J9aJktu4Y+olsz
inAQkDJ7TBU/5y0Cy7UuEn0oC907dUrwtr/kG86BNxL/BHnsr1x44Q7qE5WaCgPTUd8Qprz9GA1o
SofcSpxaKhSNo5qgiDWeN0pB4ieFzqBUk6S3+bPnrcyubHdWdcv7m6JeOWyliHO3QdDClfj7lXiW
w+vEfdZhUFaxMlMga8fekKNIXsMalPXO95x7uNl7hpzjTrijwYYpRmcmwRfN1DtKThNCiXmdgsZu
0zVDqVUtJd08M3th/x1hTSK/9CkM4mYJONPTkz6FLH4EbxLGXqtjoeXVpHw96NynIm3kO+Z41Xo1
clxSNVx9I3K9xhgmcNtZb3AiTDs3dkoxNdE6eA33Sv75xJvj9OYBTKPnBUxPUXNlyxTXAqJz+CCV
eQEQjC4Nybu8WXBy7vhA8/jA1ClzHXIMi3YKHPL0K/6NIqdo6+2qVaPpiuvSoxFSdCMisln+4OVs
fSDRwSNj+icE1trnJD9O027ZYmdvvfWhci4EOSw6NFxi4AvetsXiEA8SGNd3y1fhiVOHLbCsLRVU
6Q1hY6tdYGQU5tj2NWbaQyTwBynQz0s/IQ+csfdJfO56Fd67t96FriHD7tavfdZFMVQ5IBOQ5V9H
+/N2FCYWdOwwVd4l9cE6/9tbySMMbEbYkTUzkfL7fm/3kkjhE5rvL6X7gDD0w/KzSIB3A9LgRHes
5Nq8qshol5DDRZ+OVq36qnSS3VRcs2kcBRzd+vt7H067fsPnET7tg07fitBnHs33rbTMQmc3zWt6
McgI2xN/s7GxZ0G8G2gJEJKhrLGPWkaoQ148X9l5EwiPdRCAwRcouAlZo79/G5lH3XZff6sIFC+4
wQ6O4g+ip+JFMcKfGR8AoXf4Ad0y+zwitIw0JMjgco+V4BFcDxQh3pK1fwjBkwTKiohkSQ7t6djh
G8wSvbid7JT3PfxXERGCJPHC41sBqcK6aABIUn6oEgKHFjwRu21qsJomcm4BeG5Axw1M4Ogn231d
kjvigprgIR/1FP+ZLf06DLWBLLFoVsWd0k4JfQusAZ3BcmcHUiOVCLQmdQIAYmWefOLEePqVqeB0
/Q+ilazOVr3TpWvA0G3/136NHcJiWc1rfuv/CB8gXqEFbffM0Zcdsh4O5/HFQ8Vsw0+gJponnnsC
IzUCY1YuVcGkjXykuMq0eTIHsRWuXrrtuZEHfH4TOA5XIJkPjfPgXjfFeOxoDNSOTxBZ7qgEzuJM
O2xb/xRe/twEiWRlVCeXgT94ciNqs6A/r5/W8PGI8uSH69J0oL7x135RG2SG6ewO2fCxq9xiNBii
gA6PQD/oPH1F5dt4FqPlvsaWeYmZxV/892xniheeRxz+wUH0WBuXLkBgVZqDJZNoipJRyug6siVJ
Pe1VVqnB8dDZoymnHGA2HNNcEqWkLKYBNz1kyML7lZRqvA2+el5hT7Z/lteyxtBEW89+Hi5ck849
A/68DQmh4WSLJ+WX/F2Vg3XJK0ChWIBiO/nUety2MuQbNcGB72VNMxhLuMp9ByqdyLavg6y3sZDr
aU1EKS5mkIFudyP4cBja5e3hr25cMG3r9vYUIGanbF4oVMezOnxzuVm06GK7fRuv4dyjilvRXjTZ
eWFufuFoKMwQCRVTd/YpjsUoFEaBMq2d2sFEAJNVUWJmCXeNlj25PLUgYQo21Iul5BK/y+WVuif4
35aJKDHtM0ym5/Ky/tuChbrOrSyGpYQQfVAduIh4GN/h9oN+goU2V3zHJcyamb+YcBMU32xTgOh4
tVjYKBEtTCzX+qKi5L56PDN6nnsD+wkIDSkytt1858z72eQe3p23oDQRi0hajspyG4JFhjmTlr7j
/zRkICfbjOzpdx4oas2xV0SdnRb1iLAAIZnVWwFFgfZLrzyeYQBe1a4j50lNQFtjU5RWux2Zix9K
p6yNi4wNT2oqIq9xtp9bGVg7knYDDuhAjtP3dMegCxPVFZ/iHW5T4MHyUiS0sH5Udby+qbZGtFY6
F+BsCN0PESMqTaJeosLT9obNcA/ysjFtLe0V/rB6jI/TAqaYBotDMynLAg3QrZ4fpXWOcdO5+UGZ
W4uRtSv/yTmJmMg0gsCXNA5tLuhOgffaqYSyQzbYnxn/07BJdt+lOAPzV27quc31UKd8UZGekC/c
QXKvG4gUcE8t6iQrJc4frkNRytqQiNMYxRDumlZuNZIawuF1GFsdnEk/zhc8ka9cRWRruOKexkNV
j8NirQL7rKLQbMYSW4+E5LM6WSI48QTpkmUtKWcr9DMXjLi3kZ4dLZmXsiBCkCgwFMBhI640iQru
rcq/cbPqTjAWRVRthsse9cRCkynia0/7neSehJd4Kd3zNyLfy+LyZNXLfEwhQB2vUt1OoHv4mu5L
63PpIx1GDyn5P8CqP9quycq+LTuyKu5qoW0TKyuULEPz1WXJhpMboT9fdDdZT0cutuN+JWbObiIX
K9DM6UxMJWkgL1Sxt9TMTURkh8mzmlo4ucBu0G+moZrQ1s3ovIB7o8XNIQ7Dnixyybfuqpq9UUf7
LmY8edBzPMfoMU+wsraR8vnJSEpgIsckjBnen8qBbb1xROWIgTl53xDk0NCXaFmG3KrteYJ3Nd0a
fSivJfSWein+95QJUvzUsZMPSq6h3tjNeVsMGH+1+yKyhSNdSU+TKNT4xO1JrXkxHcFRScBZNx9l
uXhtZeSB5u5py7hsw1Uem1k3oTBQ8fgBaK/XSS/UUUKU8ZZ/11E5VqrQyqhpL4ETOjvUwAwMcbBO
5ZGR7eF4IHlEfsTiYjl/89njnOaARt52ANSYn0rJO5g1lmPDjGiFDAeIq9YgXL5WgyGRw8XNOjn7
yuOf6BlFW2KAd6mY1YVx/h8qXCl8gfTNly/FeeEQELJ2lKDW242Gxrkjy140OnyX0EhxP30VtzDL
GI936UohNBxU7LavI+W4anEPMYb5eS1KPe9gzFq7aJlqvdXzZvHtDcCZA2w4Y5D9M8BiEbydsUnr
4uElX1GJ/gQmtJRVPyd1/ljhR6D2RIWn5t5S3GVrMjLI9PwVn017v9jszuPiZZHCgw8L/uI/6CoK
g+swTNXfFXCmGB33zK4Pjt9I56/EiicYi18n3eCSp1BZB82PyhVXOyanDHfReCH+JcDhaJJ+rYNh
kc7netD85G73x1hKQAvKKoVkyizY6hG+OsMeFYkf7L8Pj3XQa+bLwkg6FIxFiEhNTwrRLEtpQkRr
V7XYd78c3ofqfIyo8nZuSqLaoSycbadlYn2cTNLwamYzSnViHgtDg6kclV5OR+nhiSC94x2m/QC+
fR7PiqgitOjEQnSrzFBMdiRNlbwYakb+pYDr5HqkqSN+SrJ7jKkT9989J7DQTOwVUTTOPGacATjM
0l+AKF9EZONz4oG90fyQpv669cdLRy7aK3dyEyPA5UEuGNetoW8j8fx+eNRCLJRztlHP3jaaDTJN
nth8GVCW88CiajAq5HcQ6lSmH4e4Cp7tSjDaNxIIRyE3tiGbLUus3jTDhb3yD89NZIRmsZQUkW2p
Pxiu1+dArVaiGVfL6im+4xuNR2WtoYdPwvQhpHuzJ1IQX3M3G3qIhd7BB6hjIGtuFVZuyW6JY3XG
W1nGReqo3Xo3hinkW+1MXI7+WaS7GIX2T6yvVwD5BNBHlRgdd62wkRTYVWIH2eAQ7ksb6HtdXWgD
xB7j0Z1KxKDPIbGQ1sXQjM4qKkwqAsaca5A+m22BV507XfyERUjQvQlH3Gzy5f9dVuUbspcGyli1
wM2cUfe29mIehdUy2vneghOcmbw3HdGRbmZp420cPyHrkWacmYcF0Gk2iMBk9fqTxptK7x0Kc9mC
Y8w3I2xwetx8tpiybHBS/1QdouBBkR4/yJHL0g4NF4v8Nqn/kgZbHS8gXSDv+wApfA37pJyb4Wpq
E3Gy8PWSoNKhd1VpSLjvxbdWFQbtS/eWM1uWfR6INSN+DpCvGNVKMl+kmVBjlDCsGFK5Tr6ZRWvr
lZ+ST/dsgQ/+Qj4j26zMAttAaVQYlqHjj8wOIb9xzJVM3jOoAaVrJCP8QtcsGib4DZ6Z9YwLxEZC
LV7LNgQgwXQ+Xy8k4fBM+F/DczSx58cGNV2Olnr77TbmH1FVNBNDrV7SVAWFztctLnPql8/T+hx3
XjvJrfFNmz8xp9atMJ8hslUwSia/evpS8pWB8ncdEyOn2P0xzg4BhknfwkrN4zkuIujImO29jdoi
oDqQ0tHDtUaxZ6sTEiVQVOU7yrmZpuWtwsn1BRALEhRhjS3ChBBqnwVwmWy5SXAEtGM10WdfOTYt
0z9xBv21xJgL2gZdhMljnvd3cVkscJLwKetIEjsyw/MPAXnqRq8gxLx7qn+ggvAbwJo3QwGbeaXQ
l05Jk6GviVB6U3BZ81R34DhrUUDSXXCG5ZgIlGXVGFg0OAbQYOb8mQKKxRsMAsPzLN24OU9552hP
vwtSbEyfViGbOuhghDUPlVeK3pPn4H4ypIJChHf9dcmcr+V2gcca417EDeD28gXCnocHEn89voYS
c8HUuVFqZ6jyfFbzaHlHIclHlkuJFqDTc0T+XjJsUUFkdD0eRygMplEVC2YATRoCK79ctQsnyqD/
tFYnTr0tnEss7kgmp2CsZ6zcofQxFUeBX1Kxnm0Kw1SnBd7zXfE8UGGWtyRyLnDuWUK2Awc61/9I
5CpOQCwI9rb6r+YoVKO6KUSeSoTtSimBj0Frx14iFYNk8xJJfr6R80+NQhe2+sbPlF5jZNkxrjxc
3Rq1HNOi/RQNJh5qrdud7GBDI3vXyVxsoZKKxGZNF4/w+rn7OZKVdQeRDveMBnYDviU5OtsOKYR6
tZoOhD2+FYmwFYF3YM46UrCx0HsVYv6HNMrcN59fXmoBtxPQJ5JID8aftYUSfERWhDuIVrewxSPs
CuwQo76jbMvqzF+zVv0gFrEvznevPUfTlQcDJaCqmOnfCPOu+419/8/z9he68kGL5GD0UZ/RIGR1
kTn75LBlyRejNWcQpnUa9KLX5RoeWR0JDqgzicdrQ3zZdMHqaLZMqTj2gTC11Lf3Jct0WMc0iwgW
tqSqsYT+qrmv8OBVz/jL1ML/SWliG/oGmlAdTHA+9u4uWD+KM8aLBuIfpe54f2M7XbUP03e/YNh8
pskja76779R6rK1fl9UAzv/N+bjars8nUKBERo/OdxQ0kz4Q2Rcp72e8s8uFKT5u4EC//UAbINkX
XNrJPtgRCAPtJ5jk9iXkk27fS0zqajL6q9uB92D0v4uLquF9V6JgNPOqi0NpXPXIAHW6nncWipd+
0M5FJTU2tSt9VQTygE9oUx/zEcQygSgUmIMt7Ae//NEdHCxHT9FSmZQ18IZusVgeXgYogwrOlCgo
N7UqRAo/OxXXjt8uBna7pUDxHsMwqxMBN4kRmqVVhLAti6kYYcFeCzN0Rvn+mwofdZlbEVIbK0WV
MNmYhp0iOJYHG/rk12eNx1gr96wOR53bIfbefnzOgmpG4N56vRWqn3oH3c4iug2ovfpYrLGU6CvL
NHmsd/dIAxKVk1vkXqQeWtJfsee9ze1yq7GKXXPVRQt8Nl/wg29OooisySI25mDb0nShXr3S5m2b
eE4+CfP+nBJMLPyDfPsIrt/Cwyi/DkxRqwiFVXhrKQkBPJDYaX1Aa4dWG3WSFf4nSgX8nBAWAeG1
f6GjxFXAXla+pNOxKsU9hl+rqesjxz7ppQgc6WM4LDz7qAkCLrFKT5xYmbnWen/wWN4nYTqbk29U
siSk90WXTlKxJR0rhPJtAv7DYTGtVJ1wN9VjD7rsGhJwersvibWb/UreMeDO3K+Zx+YqKW2KNXHQ
lUqEFcf1IChj6qNfNZyXD18LKDeeGOY2yd1tBmK7nNS2m1a58tn32Ugn34Th873mgt46NM21w/zu
P20jndoJ/GVPkOFO0boUv6L25vn6a1feMz9iTQWuEzUvnHu3u9ealUn9cWSsICIgdQLpBRu0cpTX
xHl//Dm9FXI2MCBYaNOijT/gSmj5nCxIczFj+d61a077b5F+ZLoBg863/q+qf19smanPZv4SDkU6
ASSjxQPf7zD5U4D6G5T+ikecDwTDyneIG99x3a3WhmWgPVAlnjLK0wczmLv0Txz4eLKmc0kZ6gQO
WtXMDSvpAEDpRGp7AcSEVSHBdRNP5u6wapqGXSFDb+lNGcarwplnWRTaSDW2rJo/iqUYoDGK4YeH
VQDmrg2f6ckCuWrZM8swuAI2a/x9QOWrkZaodiW2/WPC7yRaabgl2yGR6yTzby460OyU/r4NMPfV
Lrayoh/j+KGG8y5Afvk4gYk0UJ69pAS/xduQ9+HYgvF92ag4iP71PkZvPaQlH42zxtAzcw/J/8v4
+7zvScT3WuSegw/7v19EGVL5rhEkxbSXh81Br2gZfI6IwQ+oBNJQn6GJg/zybXJ6fDfMHmDdHP+2
I8Go8AB6X0ezZy3sEo+GqGI3vsXt/RalNv8hxlKtGJ2JRPKlmV9Irx1q1FtY3EsiViW76xD9UO5A
uw+QEqM2tINQsfqNtR98EfPFw07pFKV59X7vnBZwqfLZvuBVWEFeN8A3HyI/Fa0qPoyYTEOtn6ST
NbYxPWGquaNN8uLmZzHSgV8IT+DvwEsE+lMCjvE1jxnDoH642TddK4LlMlXcAt+7QSRslvOLAVAx
zFBiSDdbuQ5VpX8FgUPJnmBWs8IX/mfCspjrAg7VG2+Edle2mXRjR9zIpdiZk9FnLjWT1u009Pdq
L+tj2mBmhqpEdYaf2P5de4mRQdC6YU5tmrsJXt7VRXHFThy+ghftvAo15XGfMKSYzbj8QY/Ve8mS
wwnrr9nz5MnhyUoFAmu868USEqw6ECxp8BUxwxxut04iE5JxN7BIyASCiI5Dq6UFvD/0FCDbQ8bb
8O3BwC9zTWSxQpGbXuGHq/VcONr2xF17p64KBGkIYZ92khvXYcU6Cbar0LoF7w5/Ha2jyy7bV3Mz
Pcyscwuhg0aGcJDvm3D+54HLeaPDwy4kCu3SvWZXS8oEupqB0MwuXYPVVhr//PJwUkPJirBcXSyu
Px6YE0eqMJw1wPrMPcWLkX1o1oB1X/EVXIl73L/zTImnQFyEIvzmN/Omfp5DhuL0VSv3jibZ8n08
sh9UBR1J0/jIqc+rdodaBTTXrB/loAfRsjdWYPbs60zPRnjHabjKMf5D0wrSJnr/EUearJTajwr6
WQbQ3pQoj2d1rOaSDwZtLKfQLh6MqIui0MQvnEHMZxUja/kVwMZKWLXOaUN7ZxCfeX3vpnYzDUGq
SO4wcn9waXtNra0Lz3fDkq8fys+7EdP/WBJKnBC7UvPuGXglWG/RlPUy0Smx85+MqkUVCHSpNkY8
OoP8REiVXN+PA/M+/TjZ9Hjh7uVxdg76duqMEXIhJWPS/oe0Hy+Cs24qlRryH5xgLzuX9L1gO4Hq
LvuGuvEujdiC3DgCymPMQ8KsAWrncolz4UO1L/jLhtDhsmX3em7+rU0pxmaJefsXXIOc2KbDkypJ
2Vdtqg23qEWoiQxgWT7DewyAZxkf+9NK90/h68hy+lXgsZsXtdLcfq6auOVr/yzbChIKRL7IqjdW
bbE1jId9ArCNr9V+2XU9fVR/iH5Xm5hbIkjqQs36zMU6LECkUoOCDmWBFBkFeoAPETwrWv7u84ML
FYDtitgeMJF2sifaCJADkzVkcAFW/9tvhc56Jm06Oz2nkwK6IcFWn5TAsVHp5aeVAancNRHer6Ed
ZCV8FSmsB5DO+7KGHKoCdg6+dSmq/UZ51d8tIUVCT9PmELv8IPOIRKeb5BoiG2qSsWn7q4vZtBWb
zvopE9jpEH1kM7PbEGLWjDsXMgp312sOpvRs41Lwt0Cai22BZrFMnLbVjyl++erqbNTC2x1HVeAV
yHaR13PvKZq2ABccs8soNy8B1YpkyMpwFcYbee0c/NwT2My2Z4WsUUNamSLe6xBj/TQ5/s3UU8SC
vahwdaTEJgqNcdg7WQmuvU9S5zXNunTmIosxcMPBYEiQlmokgHqpAX3e+5Nb1h1euAyRFmNGnrNW
C5jVCDfOc6JRUwwCLKsbDqUlB2hQGmMvq7eiWL8Ah0tYQViy18mri2ab9HdqSvO2FTZRO98urOOP
94xXjrUoXbZrcPj1yX9CLicdRsGz6iVJylucEDdZNsjNcYZ+qwb4bxl2i8iWCHuIcdJcjLDj9ss8
qC5aDB/GFKJoFqoBRMLTTKU2KTARF8CTbt80DcVYYAyTWB2nC8IZgOBWcsdBVxZctA7QxgKvM38Y
oWmCdGaVgfz9dWsxgABGrcd3OXbg9iQhGBdiYKY9eG74HM/0CcYdGIy9VLux8HTb3HvtlPAy89gO
nduf3SvvLeBkgTHuxlk+j/zok2zC/2kF16ilyXO8fL6BORlIuVMfK2U7TgqKFBkAHnKnG1S/CnKS
qOfYbJevqt8Mh0mOa+LJwZJ4HMyVsI6T2Fy1EX8yOPVM0ZwaElc/MWUbtqiWNo0TaWuT/OrlXdlx
PV7UNGqvl5ARPYM3LQGB4SGQjeew+6MHXF85K9jk5kG6x8FVfdonAwhMowpj8O1eIhgVM1bdrfOc
OXvBavWK9PRK4IjUO7TiZz+QNihAgJM7jaTYxIhvX4If+UtFkPq8+20LzZT3Cwj34yPcsR2rYbgU
9yt1HaNXnv+awDEaxOOREnocouGiq/PGUbyfHywifQGNc5f86gU87JWiZpD3Cxh9Crwtslg+i/aj
BCAmF6CCtNoargVbEVdsKcAmbyhakSXXK9DEKD/v+hFLuDuheZFmOJcUjXkyvP2yaWkJS6Tvm0tm
bQG9OimBIPbzdx/VCkSEwyz+Ew3CPCcjHBoXO41lUzwhQtBl1DZHLlsh76lrSmP7DUHALZj98V45
vtxqWJMOXcSWylUd5nHJLjWxWVdJlwqJzSEP18rZK4AUhUTnjzPYVLWArOfQDm5agU+EbjFSalHM
vtC8FhX8DCt5g4TvJ7+Jf8VvarVD2IOsGhu0Cnme0ewWb2lqvRNUiEywub31vhJwQngD6ruyF9+4
pi0ChcC7nMVzogfvdEWSf+V1Fq8yNv6msI81LfbKNTis4zmEzsPFjb/NB7+omzu4ovDaSjjV0WGy
ZqsqfVBJ7phVomhMFPk9JstOvcHIXII5+yT0th/zqx5F0/m1CiCt3zvmps3liUl0QE/3acRkS6WL
dZNsKQeXa6/kv1GWg8ku8TCCIok+DrkW2TDpyfn4ibO38FhkUEw+rPNuAXsyZSn5CDPQX9w+b/Aa
l+G84R/l5txPJtREglbZBBk/x+apTr+5XtTYvXQ3t+C6pf68yeBejQI4LuTqYKiVB9ovSYG5qOre
JjdZBm0MpfVTiX3nj+YxKg7KA5Jkr7wbkVb6VVDowFrN6Mul7sqPYDHW+BJrp+hkw7Bx4lUySD5l
VukgPZx55KhIAnuICzyscF4tFDtl7OHZwPtyKDmKgCz1VkugR3rBTQfeSVsaMDAUw8cAQzriJ5FZ
b4V9NWcUrVk2uiUIV8KnoSRVXjVYqEOCqN3rj0p2mqJk42ZgE3huIvG1ldTCrxLO/VusImeEeXtw
trrR2dB7sTnqrTytESWy0UuvJS8VBSRQ2DbpsQWxWoQiXBdqkKNwY/r6c5t2/xt1+ZFatw4iETHo
D0toxFSH6UUvF2P05XF30kwdy4nXoisWu6Cgftzo+0Lb7bZdHvcbFei2bqCyB/i3KYHxFF6Kf5+R
fJNeb0FE/kHi5Tvp/YWYNQ5c962uuZ7rfT8E2mh6qWmvEZj5c+EhCcScJN4Y78nxYi2JakBq5kxD
KXw++Axef7UzKgRrvrGJkzDg9Uf/anS4hMh57DK9caSJqbtQG4bKiGwIssPQffKoYi8gLRqN5tEg
I3cvVUIlfEAneJkywpWTmtuNuFS4lDz6do72JqRJBIVdnX/MgCsDudzhgk3zfK64ExP9HvKgOMnB
Z1GpvFwvd2QUibtKL4w1s1GxKSrCsH1Uy8RELTzmZjJh2yt7clVIJ68U8Teu0xbZNKZSbhMmgjl2
U6EhB9AFkCwpJZxTqPF8e6hE3HaZp4L/6x71vlPchQuRoeHa/mWkZ5jg7sZJldWobantNy0aVMLc
EYLEJJqzGS0ZNtja0OR3JHDrA0UR9MNpxUJJNKmLdzFyMUsu1fNa5qC+xewXTsSUEp/Nyxo2V7lL
vdjdiGPJkpta+LP6jYDhKvWzAGC+1pkLMmrrXgUlBHHzKr3zDpfUl0spbvmx5se17g0hAtTzPYyL
Aa0g21fltRcWA4vd0gAiYxJsja3BJbyX1pcmMTLLZNZOb5zNm+aHmodkO1bUblkkYc7VortxSwp6
itqUSYW5KCKZcOIBg6RoWeTJT9MgVg6cbGNCvKmRyKuRtSXVCc5cVzobNQt0qh4xVatDsJzY4467
hsXmMFgO8xcwD4hYLAOLraLVp+btkPWzzO2I1WLt+LcFXbD/ymvjcDLDXWyWsgL0Xd1BgnfqFNU+
GT3xR674fdouclFRrorhA72rcaMjHlf6mJs0ZmuXQv9jZRCjNR/0yipDs/CvrmAEdtdSScAgARrW
VThmRv/KgJCh4ren5pn+veXCP6ELN1UNDEjIkPRgTLrMHYxLjRWQRpIhtgLukrdD/toxAS/a19oi
1ow5CISQl/zEcdcB577ywoduUOWH/2jXYzfuCf8svDSKAW12sLi0ghrsAYy1bw4ZfHUz9t2yjnMO
/CtFIOF4/hekNXn5SmWySXZQWi88kc7Wl7F877x95hHQiYcZIuLSqI4F3ETOYod0OnqSCr4fXyF1
Ax3O8ImoduxcomZgXLgMqRYsZNlCC4Gd80Ud3cKcvSK1HRA5Al6L9HdW/pNjyH2Y2bUxer9wP7qu
9bnrCWHwUr1mLpw1B3yaaG/qterFuXsAEU2HHMi1UiB3iBlfHF4DceCrPPgFq+1pDiQfYkaklWQX
N7cVwW4Rl6hS3+TSRpGRBCYM7PyEhNo+9wJls4P2uEcBcWkNjuNKQOn2HOS0T7kJqjuHrEwGMJ8L
wqM2m1qaEvEzDQPvZA7O0TkEX4IY8uaJHSi3KWhmtFx+eYUiPMdRTwQuTky/3K8FLl3dDMc6f+Ly
GPQfZw6v+RMWGKmDv2FEkfMahjr+xev11Ug3/H2IW/Ms6kJjt3tj/LzSI8tKtysBOFQcAEqhgAd6
JBgNIAReJ0X6l9quu6mtOyi1L+6r5XnqR1eCI5X9FTj50SRZ5t7fad9iVZ2amEVSam3MSd6vcRtk
meI/HHj1kbZ++bp0CG5mZCZJlB0SmWh0umhJ+mizNOqpzUzBX3/OiU0uxbrTq2dax0p39IdPfsLW
6wxkmo9eWrROiS2wJjf+GHXJkdp+GHk7xZgIJH+5n/rxFQkC8yF1AJ7wB8zw9+UI3v8atikbvszK
RdbhGSKpx7pSm6CbB87V2Uw/JXisB/Af++qVpaD51pX9f6g6mm0W1aZkuBARyFk+5RlRTjHY9XOk
0AeCYrPuTgwoSDD0g4k6vLSCwXBU89Qou2X/BidrwLzgRxeW3568oo70Nm1BqI9U9CnBEo/sT4Ih
D0izR2Ehj4fcaUJ026UEFVDNb0leDKwwIJS9o9OPDQvnyVMYq80RVJZoFqjKb6S9YtEDB325Ekcu
Lfs5IeY57Ipd1kEoziWKLYpcUpaIEDAtdopfFOQGZ8nMxFVZwaJnFjuf9hRwtvstqKCBad1s8v4d
dAqal+JDHKdKEoQqLJtjS0QCpjsL2HqFFVrF6DIgUaZlZf2R+K8ZQfECdj7Q7F9v/Qpve0Cml8VQ
9YuhdZ0RhUUEBvxxMXPV8EMx4Wbyeof3Ky/Y7Jh1wlOdv7zudxROnVI5xOZKg51sy7fvBu5Y6oq8
vncoxMzwb0gjWPP6YVkBAXwHfGqVb7uWWI+WlB/0ES5n9uzX/OdbnkSRS7YSmBNZKUYdMkwwjx5D
558mVC1zcc77gxj45Z+RmGXaMCRbL+8vFmYMUIOIqq1niDmmcqRmRneCqkQs4gUZn+TgUGnHfSgp
Jc5AExw2b4n8mhKU9oqzf/bW4b3JKW6a351ExMMBXXbs4zfMzRJsNAEKEhHOW+cY6IxzGjNEV+5i
yP+GQIzZL98Jqu93HaK213MEzunhvkgO6m9riywWomOBe29GYYfXDBiRYUtJMlTt95Oxmse1/YF6
Ej1WJg2RGBx7CACcA6uraw6Xh6Ska5TcAc2mL5ZzFdniZDlMZeUCqoQwoxDNyBQnzf+PnRopFdtg
9aglmHLBXPUfyWqmgQNlJP02NUF6XdZWFzHqasu4bhhDNh2XZBrQC+HHfFo81NsrKo/MX68Ds4Eg
ssDfz50L4ceLryOZhT0+pr6ZPFH/GojEXQa97tBbGFpSISZtetVK+cyp5b9h9Z2pgW4NGX5C2BaJ
qNltKXjGNBEYw7uwAx9p6Hz31h/AOC20QVanXSLaP21M/ARFLlBzjT4ZA8DjFQ/cDPme8aEDW2NA
MRXZG8Ndia+WFK64jIV5QTAOyW1KHS1r4YMColIiyx+3FqnVv1RLx3eeTQbZbaamFOnZ+PApwRLs
l+Zb8vkrtw0645Y+aG7vJ79z/GF12e24BjKJCIAht++dVzO5r2SzlGSg374h0m4QbHd8pjyOrqSI
PmWfUmSs9KH9RfyZByMjfedHDA9ig5ey8MH2GkgZCFcr4EWroI2ukSacufyJBOdxQ/TTFrycSU65
HJk3lSW440pZdIWhfh3QI5PxUcS2lhMipwsE3pyvwIJ+7cy+rKPDX1tY8PmE0PXvvgiezDVeUhHN
jjel+FwipSS+wnUM/+pRX9IJFdTm6GzwyDKDKkNhiv8N4qiKrSVohmBInRQt+xdb4Kz5hLVd6+OC
GIXFERkJI4zu5ELoNcBX0afmrVCSWi0ZxUqDiXLbpOiVgAH9VTzKLrF+B5uXWhekrGxEnBtIw1T9
DQH4JXuBz1TVaAyaHPrLAjB2ZUgmsgtTy9enmsehapx9GjCqZbf/jNeTCqb8YT4Vga/59ETm2NZg
XdS6lwjhjOAscQx0A75FbYII3fSPNg0G68lZlrGbRdmTuRJSWlflfrD7TPBmxWEHGFa5omBOcFYJ
W0RRMOkg3y7UzaUl1M8CZtb1W5qkq2ll5G9VXuOFw6y4EYzm1N/Yd52QhbGY8Brdaf8GrkLZp81C
kLI9UIdYMMasu31PxuDdnGADBl3+6+fCWhBpnAfinfM41643b55B7KMzLx8p3rHFeWa4gbU+j8tv
0hr2agCA/RjCTAf8U0DD1cGaHx1/7xCV+hM/wp9ixG2sD/OqM9v8uTcPxmn1zhkjYD2+BXd0T2It
pPSc4iqWYIan1+EwLN5w5nBx114tVRK0LfYDvA49oEvWcuR1urnqk1RBaGAt7G51neUArlttefGm
tXsHGNwMsds8puWe9TU194FCFnoPh1J1O9/EnebSXYRRKwUbkpDph1jaqAsYS90p1+6cG+a4SYkh
qnrVAOwyCNSP6NqMKhhzDLo49Smo1/p6DsxdqWeu8BLsnyvCfMFGE7ENA55bTeRZfx3EVWS61g7o
VI8uhqVOlnogDIaLVOXLiVw8F2Z+q4UeMUNIhQ8uIMpTfZduUJ7mLBLHRCigtduE4LCfPnetKnHs
OHATa3iKwcKPsqIxbYFBEBPQBnGK0PEYlzdvV1292HfODWoC254QgtHXXKyVZYRu4NupEAERnVvP
FYMOvoO+Q4GGaInrFByZ7HOW032KP364rAcLxNFtFjz4rPHxoy+QU3ua043XS2l+Nza9pSgh/HV/
Q5rZgDuSU2SniI9yiGq4QQbW+GoOL+O3bvyKXEVqfnRudtIccIosM6NJIXLkA3McAlLdtBl+wbli
/Tukm2eQfJHfDT3sRXfcF9Uu68zP7UuVeD1BvHAk5iCGQgg0MMFZla+EjJ9M+I9T7wVvkpA1mibz
paSqKz0KBOi6PZ43mn0givOv2hQcoMv1mou0NAfsALzKQKMFY97OcVXe7cYxHGhH6GmR/f4gy9ld
2sp9LLLDdrUPHwN/Nwr9Io66teITHsxJfyYmFa1x54MgryVlzRigsntuGOxvjC2Hdxf+DC2s5lT9
JfLw5SnPI2wr+Ot5KbS3kH30ltN0qNyx41tHrF64zpLG8reH7JnP52G1qxYHQfRpLM0Fea4Np9JA
LX8ElLLQP++Jp8JSwdyP589P0z9Ln3f2QAGhqtlJ73jLYmc2we/cglOxTesrIA2boktqtM4oNatS
9QTNENSPyQXyj5ETd79vX8LNyFDl02oIp7/lwboix0sZpKZRtITGXqI5SWjUMLzd4k7s1jrehQbm
aniFImpBTdhLTk1KcBfl2nZdFrUlvtWHWl5wUIGNdXnfqZdPD+GlWodWwRciC6rlPvfxfirpQXiL
7HDSk2nFFacfr0vcucGwCXkBMEdnUrSF68LpIlVOD/gUVD+ZdJnIE4XLZn3ikaU/TOgTP3yepMT7
vyBZmIYu8UhvfRkUQ86nDYMNESg7x5xmsTbWyhERsQRxpmNPySmL/h/lfuw3UoRuCjMGM/B82BuV
7GubE4+KOLLjHpeQTk3ZAdxNDYlnUDOivK1FLgdzLFmLlWUu5eDfte0YpMSetihr7XvMsinBx3pZ
wfNxBxM9VhNYIseFuFP77C7D1cnM260N7FrZ25XyROT5bPY0XlGpH/rxA+LtyVWNSP96Lp+J3TJD
GAUQxuUWNMC5Qxa0e7/c+CHTsqWU0aAYs8TDkdvl36n7LLeEeeTl2IhAfgRWaQ1oMJ+sT93nwd44
hh3jOMtl8KkyUqccnmCUU2vjH7+D/kq6DeFQHrvQeMZw8ye+ZHzK/sTcO2v5Jbzz7Lo4YGVntVSo
epXg/qVaZ0DuYeBhb9zNjEzDTphIg/qpuETyovxX/bkRFVLhiz6wk3cFqBE6Mq2FzDayV06sE0bC
kOPkM7omV5J0dVNGQn/ZZacIqmf2oKYLbEd97Q6wkyIqhVPQasi7tD/Zeav3Y+Xh+3eo40QYU/wS
zlzIMjgkvVMGQ/bc18BM6FQr7+aEZUVIQdqFEM8K3q26j0LHa+xHkvg3eijw3oaleuOrKe1dj0LL
6Zm68Ed/30a1guxHiIryVATqxzrA+skqW+0E3uaxf+wlTAmymuHut8CJJ/Xc2natCWCCBpl+0a+U
hfLgLA7Q1L5gsKzdEHqfgoi0I69yOL57Q8L+wC+wJBL11lEGng6tN4gOiD5ScsaLD7WxBLPdnyXc
svXVBZ6tCPB2sTv97cxc8b7QbiqwOM+Ap/SO4xqBpVd+1nxKogzWUOitDQFW0pb05K4lyHVX44y2
zbN7zEFaT9gbq6LdMzjTQCdgQE9hbCWqUxjKwxRsFpOB43CQYWMy7a0pAD7fmDMx+kafE6VLQkM8
7G4ZuYcjIHkeViJy75rOFz4b35stnf3Ib7L8uyzE3p730jJjgHpbo67xsuiZ8ZrW/KllXxG8FeZv
AAVEeTwXXQzRynCo5DnIjAzleZB5qa2PK0T9TIpnK2rZxoJFhyhho+2JaA42b5Doy2F9GlQ2g2Nx
eWhASX1WyyJYjrcrIed02Z+BGiCoXxecV4u8j38ISr9vdgfNsnfrIjJY2yiFv6pP2wKj+BmACcsN
qGUEkxthH8bKccgbJ9mI6wn+oIyooJDK8C7N+/6qgtMHjPlzZcCRQwqeQVWYG/cS7ue5e9VHRw5J
A62aYMj/lbsooNeK3uldTgV9i1smPmtI6I02tsbGZrMvTulBPxvfm0XeWGr4tCYBuaNYKR0iet8F
dFv3jFr0AJ8bYCZ9KUdITkqJ0m8SDGfLQREItOILxpAH5BxLDd1+V0bUosUePOe6zHI4ozoi0uD8
VyXyep0KdDnfstkXeRvQS2c4+sqy2y8TJcJI1x91F2DwLTACk5SMbZVCDWvZFvG4ohIhCASMViba
MtRM1E7aNimuHkkyF9AABc1Z0nkzOugV3ukX8407Wt84pG6kRINk4aoBzKrStRCeCnHqBJqNE+/H
iih/BVTTYBMwzoWwgGhsgbIijOBRX6msp5vZAHLmlnZysyfKa5Bgu+vvOSUPN/JH+hngM2LcDafy
t3HWo5I/2kb1olwVGBFEC9Uu7n/yeCUG/7akIPK73y7L1R3Zqm01g2iPKlerFtVm14oK5ByK3LGJ
VrjvfgcpB3xLDnXpFrKPbfX9oMuM+uOPM4MK164ZTQC7BxWoRWOY8Ysg2wcI1B2w/pzJ/bbR/L2f
QRes1LoJRYMJ8XB+xD4LlRElOT/VtVRFH37KscZNDfYAxAqdU3WW+StcDcpwrNo58FTUhyE5OX6k
23T3NBvOlGooci8KA6vZwzamNHeVWlMcvc66B1p1IOghDVPFSNoRtiTkclWkAgiUrm4MA273tYKZ
TgJfkWM6Ec2VwdYnMdzm6r/U5mwzNnt8RPDe4HZ1F9Q38crkQXf2XXA1ZquDjawXqbwtrjLkwyv2
bERuteqFRJEpAJotYOgebPSLH/E2vRzsRPIAeyy88sZHEySojh/61p+yXuxZZZdvbNaxr3EF0f+b
i+/8GOZ2JEBWpBBmtqMCCoe/WFRVMy6ib1sTTg6HJuKmeOLgzEPHdf04rQVGBqGZ+M0H1b8mAsZ1
U2fAtG6swI4EG7JEPWDakQT7lkioMd0YVprO1PNhxbk/MJwdywYd0mYxgjIGb43IAXGSUG8v0T9u
PxI6aet3Z8j+cI0qIrpzLG8iPkpbkc4xFQ6fB9oIS2Ljsqlx6sXbDR68qNO9sI6DrE2/0uLhlZ3f
sUrz5/i1YD1W9FgJbBQOnYQnG9XG1E8lG4iV2LTFiLzpoivucVHU/tOYUt2TqTGsJywEer8/fYTj
m2lMWcqSlkJleRtUHbyUEXedNHDXaTpba8Xe4S083uonXEqp3QV/AOCfNv80VXEwGout/dlJogkx
jZosijobdqc7Tdv5fK73JgriciqPWYMmaf5S5kGkN8z/CeX/70u0ePhZi5suwtFVIsl7NhgMu20u
hnBCxB6UVJSZ+oOEjb0rqBumwMRjtHbbPhOZd0FOjOunGDi/bgSs9z8MyZYWnESMZXBb6uyhsjVC
tyMBvmyCv7FV91tlbA2BnTiw1czH1b6FdGixNySaKrOUITBPOcg7Vfr6QXvdgrwpVByK2wOhb9kX
/A7EWXDST5BOPojE8gPA0WuwcGYptCWny9DuZtPgTDG3gEcDvrd7ivCKnLQl8Kwp0RYsVoufjaCI
k4URorNrprvIJzJGyfergg0KJ4m8SCsqJoB0I/g6Tm13zayAteFrFCUbDuxkVhjM4mkTROSVKW27
sD8X3oh6SSP8PXGSGKViIdTl2eKRErNsUYuQsyGu1YF4nhJKKs2NhLSHkExNMH0aHEwuqa2bZfIC
ho29zd+ZY5JMkrnRpfKPNyWc9tqT6YAnGPhcK5X6IOvDH/wtK6aIE+6POjpXcHsfta52VkqW3oY7
dH9PPtLjb9dy2maV9XOuu5Onartrm/LRc7FcW++vGfGlxsAcxHhCNRfFwaVZo0gPGm8GCx7uz5t9
YBufvNMKaWH6wnQPqQ/Q2L5kMyeGj8FW9AiXh9bYE8t/CyGZp4NzpomyN4xZ1vSScEKNIkuLl6vT
oyMwZuOahQDNqIVNphCaHjb8jATscw27b0fs5kMVn5FIRxLe5i+GKOczaknK814ZY0fvJzH/3rN5
vgHy36+6tFgn1G3VD39VNR5as3cJ+3FA9ty4/lVZiK2fz0O2vYXKUnIwEWtgCAs9aWiQhrnMi32B
WcEgJ0axoMVRM+XojVePb3w7SKjz4L86awfu1yNzJoyBX1fWphtBB7RdSKC6Wnvz1U24+0utKBMG
YSrBcwjB0AdtHRhfMlTLBX1QQlsJ0tvPebnPFuhKNMb+KsFJK8Q7FOtmVuUkMXGsFPDbnQIAhNfi
wjsgkLBnVExD0FKSNJwSGws10HPUoA2Lm7CMEh/v6NCYyYeG1GplV9xtPrRtgtYlgMrdSsgvwGZx
4+LGqr3wQ50/3VKrE/KZ3N9WayyJ7Ouytahun7GIVNaeDI/bqVDcecrxEPgKQYc567Bww9I9rras
ocEpmmAu6CNYg5POGoZYeNzNRJll+4N9TNOCHGfzDQkGjxc95Ij46erh9sOmmlFzSa7ekBPFTb3r
21vTLaNdO/YmJ/E+sbpy2zaF43qIYUHOSgIW5spNetdh3Nspa3UDXpgR1/INwFZtMFmg6Q9EjciK
BwQlitDMSf8Vk/EAbLUo699xwVOrxwWePuDsJGsmBKdNhtz4pp5MWpeG2qbVCLwbnxIpO7rwzy+/
dVMkz9KEeB1sqykrrvUeHUolLyHuU5yTtfSATHYy8OoegXmtK362YOSR08a90MdRaDBLw88RWcX0
IYW0qkqsqZrSTSiqS9le058jS23WzSkIBFOY6MRIZWmvkwttEpk0DI4VroOitMOzjgORV0dUG7CW
KDMli4S4SRnQ7pNMwN5IXzlJXQPQ7Nq79evESvhqr2nn9pFgcHBPzD+0Dj6HrYVy5odeHiYblUZG
g6GnGTdg5fOM/2vfnIG3MNbE1caZnXOZYqyBeR012CaqYiMUcISHMaITIWjfbTomodUN7srdMemM
bhG4Yt8a34De4pdcRYW3lO7yzYnlCYceaMZ70KJgnyHjh5jx9CxFJ0pao3ImhsCZQrNPMG7o6YYk
y0Ug+uzcVoGuDXRqiP8M5+Rwe0MOft1Y0dPF5QSwFEs6Yn7hGHJD/KV4KlPCOmGfMPp0KKqQIvBL
fClFYJlpJixpg7An0rXFPyHvKtdIN0IlYkM1LcJHjpUUb7wKGUZDDpBQQQ5iCUeSwz4SGlAtxBmh
sh5Qzg08u+yZ13QrWU6ShMDWMbp2RdLeD4pFJ5NdTiw04Pi9IzzbyLqgfVdZsU3WllUJUDSTseuz
P3l6jJNgiChB0EOsIwnvZ4F98/qoJPXyP4JPCdWiTedqpRDH3aaKoGx+UD+gD6ERFKu06nPEbf90
MTNkXGVivlX7xPiFcgJGDBF33QHAZDzTkhtCJiSp23PjTJP9oAn0NyoPoLp/0iY/Ebb6Vu0BeLLv
LBDZPqxKin5niCy7JNB9mYo71pjREXFwDwKMtQWI++vivqnDNSen8EGi4nhdQsowgSdzY2iB7XX+
rfdKT2yHQiRPY5lVgLjdW3vERwx4zhlmCYN8YSU8NN4tj04ketgEj5RaTOkfs9jj3Rpp/f+F41ua
KoAiV0WCICLPcBe/EfVUmJOb74LiMAg0uBpGEVD/A5aCZGkcBi6jC7pHLW9p0uGyTKKAImoCGFGa
V9Wdt5rZidO7gzKipChsZiYDsw87slHEQ7EY6Po9GvIIa0rFy1VFrlTOlNzU8Gv1t1vkMBLM3K9F
hx57WOWrGZP6Yu0jxR+Jwxz9ZOTSL3UzpHvKPNbC+dZbKlrf36WvZ+CIHD8AXGqBDmFolx8HkfZ9
PKjOXTC0KDkYENrGRhUDbEze5to6px5wgz20k67YmYgsUY7P8zGzlh0VuWneFDoWRO5YlRfwClnr
TlqKh4TVN3VhXPTRJp7icnlCB2Xd9LikEaOV5z3ja1G3tKaaCEYc9xmxXcmzi4scZiO9lZdi9Ip4
DRa0IX+/o9YrDKmv2MHds5SBHHl8JwBN2AeT9/QvqwwUbwrdBJuWZkTNn1fzuQ38lH9kfIWeGP1O
ErGcyu0MTT40DfmAATvlJrqpMVFVoAIAqyY5BmiU/iLuxoAmV+ZrVsBqU0QvJpxVm+zVzpiXKNRn
hl5v2TyRDEf3xH6BLtskvSpieERbjx6PHMhXeDytMzb+AVzDwS0GuY1jT4Cihi9S3AaERUr+g9z/
tbQWgDL6TyALef5n1UJMsOeN/e3+1Pl78AH2g093Rw9rUE+8XRXTfUX3dyqiBLabl1ytuI9OrLtX
zJLbHUhaS2p2TYPm+8X1iVvz7tk7nsJiWhUXMzCNnjqstc+IeIj21ahWE7aA0K0D60uFbg/qRhSn
ACo3eceuH5yl90DQ1d6siZl+4sE1Ukwy/JuaS/SFD+fSCPaurNUqByOLlMFczGVBWJp199XiL4AG
afKP4FvJeGcSr73sXGfHAuZHo27qMP6JTOEkuLkkFaAfMM2MV0tLTqrPl24c21wGLyC0rUm6bGfN
SRGqk2WtKEiPzRv/B3dfu/fBBtoXxlfi/DN6FOe0xFVTZdEtmqc94lgB/RgjhKHB5Vnpvi45y/pB
ER1RdJDzsGfu/IF41AqUVWenixYvv7Qqf99F+MyWgPQ+c4qcQcl5C6CopendizGfcLCpZvdEzi65
m8R8AtEzRcWpOu//gTpTasXbGhbvApxF00z5Y7FMnu0+0IOOM+/wbh/DbVGiqhF7FyLdfLTzCXgf
rqZ1pTzJbxvOaPR8i14ctwzCzybJTIrP2Ik5KHgCoVKGM4POk6cBymuKWolc+39gDi1rcLXh6g5Y
m84ulVJlbB3mEhwrU+r7zNNZPktx8wm1fC3t09JPZA6yELa23Z/G8gecC7tfnyAdpvd0/JjiQMHU
azgtS1jiOOAfeMsAsrb/p/RRyck8zCtOs4yIqcYB5GG/+YaY+ymg/t7AN4CnzHjl7v6ycg2VUQFl
qOlTxmLSOeANKc7JPwZC+z5lJcLy6GLrqhKloOsclZmdvd7mOxer1izo/TK9g82LrLN5rR4enkEF
hggIikJZ6DazY0nEU8TbQv1xcyUtCro8Zm2XLAEKcVVUW0Xyn/GTJcVboLQcheQ53J2DNWtkNmCT
07oYX2iHqnzZxq6ZAvu1HYDDg6meS+T+cqmtPRp/PL19KZdxWwwgvzZrK2EFwmqgXU1jO7/Q4ATY
UFidGpuk0pk8wmxXASJfeF752oxXuiEFdMceJmyToVdW+rtyTjNJSE06U+w0QNUIUvRJmqqcdPGM
kEKF8JQ8/D4mfgMFQsdgdkXlDX3eOoDdFKJ0OqwP25R9paqybgxeBS+GjpYG6bDDW37YPBlgVoya
CR5hS0ouhjWSQ/vnBPUrDlHO5JSud5VzgIlOFD4Mu9PxMa4WgASm44EU3aV3Z/LiwCHOxb++VjfB
45GINpkx17jz09riIRLbXQCkKpewkuplziPg0W5N0wZA2s7fL/Wm9QT1AMW+JCXPpSKliYMdVoFv
PjxR1PspRTELNFccW5qDJxrba0MYadprK0AIaUN4JWZldasIMeqZSO59ABZtWiIss+KloYu+3Bj2
0V5JNe8Rc2i15aOfif/0d1rwi+JbLCsFexu0fhTXgF7YXWBnGMEoJFVIGtnVI+8GJY99P1uGBiqD
urBNt7ozaT7D9G9aWNRstpPQkcprdZRJlJyp6uA8JLC70OU1swhSnKmn+/250icdoX7euEil/nJb
m+4ikWM83kqg5vk9JCiW28Xi2RHD5s0/wIAS8ABPqYYQ6X5cvkm2ajNkRFNTAWu39tP5WsEWeNc/
PSqNli2yfVuniF6nABriNJ+wPxrdCy3HXtQPSWmyC/jzXMjI10n0gFqO4+38+NobVSUm5vEDogpb
QYJxTbOqTD4sEbCFDIRVNlhJ+GDal+f4CHZ7KYOV6k7fTtPApvO0UQ7dnMerKZG090CQF1MPQ4XR
+F/UZBiXWQXxHQi7jf6O6311uXPkBd76Uhp8sK8bLzY2IPnEzhCaTra8CYEPl/jmQ/DZv/nVeKiL
qJwYC4U81sv16LAz2GbY77fLDAixFujHcwVsTJLWG4pJqVYtAxh/xdquXYCOwAxT0NG1og43VRq1
/vIcwsnd5E2Lp/ezzJBL4d2PI/2RLA8HAIAk2nj2AfFcXBy80tJx1S6NiZuFdrl0Hu19uAuMXfUJ
/XhA8iw3P2eUykTP8829hMB+DvvFt/5zdg4sJ9+wgEVEwtfg74yuEol6R1KhNHAqFy3zElVeYqkF
nsFte/GYtKpGJ81F83k5+5IqDWCz07IWyxTqhIXseg+VEkAp+OGQUnW3YTVELNCsqSR9iM/hfAHJ
6/q0VVl+va5kLptUsGCp1DjPUwSaFBewTqp6UhOKib/z5lFl+hx3u6ikpoStBB1ymoH32tPW3iLt
aMZ1kvsfYLfS+bGYWsjl3ilrIPJFmvhQ4Zcxcgu33vW0YxHY48fBmQOIemkRr+TwC/Sh9kwCgEo9
v3Rvw1/mUhN1agNoogBSnjDSZj2a0uo7BBZGy/MJG+kGxlw2GyIriY000LoFZAxypLs8WtJ46F6w
2n0fhCUATHxGp89M1MMhzcVsTA9g6PtP3YDb5yhNJzHsJEjTTrwR8sFgyPf45PMCdUyhHCoetQwf
IgqKN3c+akWjavxLlL1Ck5PD3neJ5UdLKW4RSVk6OsxcgtrNSvve8KmWKcvVYXKbd7JJuW8m4Lqh
Ae6S6XU23t4/P/dLmba9o50Jn35Y0LqiwWBgNye8H0jKsbRFdM8QRGMmPd3Wi8pk5k2yIHwk6Hel
fi/BF9Sj/QAPiQ1AJCg3w7AxQpw9j82Qtor0/bUbk7Geh/5XCXGOg5jbVoQqeK2wl3rnavhayGx9
8CVwTC7f04F6QDrzm2hFwKque+YdtSHe58GFta0G9tbA8AnEEuCTE/nYnHsX65cNMZIMn+upnN6B
LV032vD81WFMKHaXW4WRxCn0sCRGqNww/jBTngYFI/Xx8DTJOZMUhyu0Gy2b1gvozbS5xVGsJP+t
rw1RrtWGBaXn2T9d/zaWYbwu+wtG7cb4a9g36wnvzel93X7zm6Fi19OyQMG0YvCTs+YZr7B9Mhok
fxojeMB7kLQZru+mVok133etsB6/sbz8K1O7auPgBgC7poRWjgBIN6H9KO624Rh6Tg4QTDUh99SU
TDgmDHFXkfrnddthWtyfYwDCqirkenz6OGw38NVw2nzPBzrqZP++XDXyBrF0UMZieDlisdhIJWz3
t62K1hUHjse7qnH8qzpKMtweUXwK2DL7nvbw88haiysFE7dFyalijadQdXdo0U4NHsopmiTBk6yk
RhCz+235Z0z3ub+rcl9Iy6k0jyLPS8EqBAq2obZWRrxYkbLeweu4Y9b/tdDrSBrB0XhZ+tSgqSFt
/FK0kZ+4UG02W/5BQn735ySO0m4vYwH3vq9JFN0v7EBhl7ofA3cAW2WN58otpBgJef2yPWNpab3h
9eS6p85HufL+eWPtdQuaL0zxYlC9fhBGRebO0HP/O6fyWxpu3JNMVXBnt18jRfRL+TfW4AkUoMmD
sv4rkg6A9Xqe6EvnSgMoyspxel3+VVKTbMEFzpJv4WE80AmDTEbfr866jHp8SOKCCMJY45ZTpX+Y
ITPwVlnu8nUB56un5xCPRUQJu/Iiu0h4aKlYHEz+IPtP1buGLTP+62iz/sysm8lJyqVMQ2A+eSJv
b43KD3S3Hfv7+LwRK1ArhY6e2WlxP3rbL6BUVLCewoVbmhVi8qxv5+9LK6hdicZyQgapdvuKNwY2
B69l7uU9jIMVOQG5OAL2NLX/322zUjz5VfoumYVXdsl3nhA7tkA485GShDF4rfCPth8jTw1Me8gg
J6cqA3TvjdEPp5rFVO8/bejeBCpaAdsqgT2hV8xayjVXXfcv/YibMJXIVBRA+glJDvdAF2qFmeHj
JkT3Heq9RCx2LbJsoC4MqOmZ1H4xrE/kozF93DmpbQ1H7wvbq0ch8lyU4urpFvLeHvS9dT6h7/wl
cGTw67GrZhJBIX6cTBiB+343ZyWE4OPdVNQEA5caP7YYMvqnjsodpqvjdwDN7EXXFve1U4rfqmL4
NHcXsOyn9s7qfQyjH8gKu7yqJsRilNl0RkkDFjy9d03G/dTUhfqtJSCmed67bRF4848g28XUCAi/
E0/8BF+rmuTTXfnqmLGwu8tYqx8VThBfb6Pi7fMvgBzGUNAn2bp8sGSMBffO1nKx1YqtPmzOmYh+
9AddqAErwXdojnxrvSLsb4Six3kY1s8M7UVKsDCmPCol8Hq6BslkpLj/UGtFgEUZOH0Wh31jBT7+
HK7C3Ka+7/elL90xSEnOGIR4ULUoKy4p9skUGoPffcOWbadYuohdhmWo1MXZcLbRA1p44M4ZbEC3
8FDIaHJ525n16tWJS6gdAGxmMacRARa4itFT8BQk2fQ0+06KuN9GSDcnVkYRiWOXfREnslmivErC
AVDhUWU0w6oV3XC5OD+ZDgO40E0dGHOMNVGt+5gpA9Jj4rZ4UaHRLHkhirSFHmAAj5qHdgsXJqAR
UNbliLIORSH++E9U7V0VNxLXJmh5kWLkAR/vVvmA6UuJT5qdqgshbPWtEb4waiaDuTbeJXvGWfet
npOvslflTND9a5DnVwhco2I6yVkDp09SJ85iY/Rpx9IkRpn1nKNckf32xLADqO7hgeMJL8XfTGf0
2yP1TyD2vzdsAsuxz/5wczkZxAXzg9SSSwr12sFs5ixmV4vjmxVKEG7m/SyOewm9YCSllwJKhwqA
ZdUGDWQCMnY5pFshzCqBJRQ1aJRCboGFKAaQ/bXyRWsuE9CaI7U2zNg8SM7/fR9y9pILziljs/Ab
GNABVuyeRkQep6hSXZAccTD9514M971hOdE2xijOfXZwaj2fhLWbwAgUD1rShgO4qdRaxQ1/Td8i
n32iQWddT7v5StzKpApt+kCZJx/yuboVSEwRKzH+hXTd0kADwJMckDE2dVIRnehxEgkluJ67qvD0
McASCHMitjsl3Y49jQKcfboGLdlYEnW5EHCY4h6gwxM7dI1TwwwXGjL1UMHUyjM16kpZk+iL3T39
BQrB/YH7+6eFTbrbLbbolpRm2eX8e61hiJRWsZH0qtrvfb7GaA0YhixOSd7USpjnYg+eceUDiSf+
klnZ2ZXG5ZjciUwXBS9g2D61rlOljEXQtrMcvrbWSsVJiHvSblJh2/Olv0P3xGWzKpUZiT2qbwiv
0kz6awIpiYQxfNszoVWPjYo4tMxq0ZQc7sov33w/YMUBNdYGIa5DEuh6lc9hNgkaRLHbABkvBe9J
RKe4iXq2rSCvNX86HLXAIxBrx1vp7Rm34apmJ0aelIZi1Qjq8KRt98G7TO4wvODTY41Y2AXzzf3K
FOc8JHWwv/YLc1gxFhkEP+IWnct0gLYSvmw1BZ6DcwZoHz3diz7x0KQgbPdjAnHEVgVUdnKe3xy/
h0htKw7XYJFRe6c7nIarDlf1dOLSzvGIkszQz8i2zGJDAU+BPGYvh4r+LnqMNbMazNA5UW+IMgmm
OAqxZBfbsE1vP0WCWiZJA9iw+tp9evrvx/W35XXAhD5V/okvhBVs6fBAV0OTio1ZoaCh8roWh8z6
s/FBm8ygGBHxAHIOsjtH+BuCzOZUDnwA49U0UraQgFHNhyFt3XF90LQ7DvC3JGEOj+q4dwoo20gv
Xqb5KZ2cwq3TZDRBP+S3S4ange09HagiEvYIthdMpmeNPAn2nekB8Sbb8WuBsJpig0Rz5Cf+jn7i
IHLLBIwru1I2+cCSyWadzwwrgADNDv2AikiU47caCgmin7rYxcoSskOD63s4rNLBMNoHIrMwIdLU
/J+gwgk93hMbAx8rogHYy9XvHt5OGYMyq/N6sgrcTQAcC1eqoS0cP/LMrgf++/N2+TNp4dsVb5Zu
6pOkXKI96XAQfMRkO+HeQsfExDq/q0Nai1gtIRiVupeq6DHGxhryOU5TmAHHZGCq1im1JmnMimo1
0Fvz7qjWpqxU2jDTtUk0GLjbqJ7GtaRPKNbDf/hdT1ungIGcDC/BrNsPDQgVlPwYH7Ephhl69vcf
MGanvPIb0EBL/WpK1ot1w2U2GU6lEyl1bOIFwV8TssDflYgGHai+2+TjmaKWdW4gLkpJTqJ4ryiS
dY4YVxKnnm4yL6k6M/iPIKD3TSZIASs0XVeWI9nFX2IK+48S0hdGO1Qojmn8CvGnoRxAB8BpZKsV
XZ7cQ1hIh/Sclsj8+rGsylKDWsTcOLm4SxTsWyhGHydFiCLePQz7ODKvpy1/ooSbJDxZvK5vjC5V
PgUVA2R5YdY40MdzH48I0dNSMUitlbmFRyfhB5i1FZlvo4rgpv3x+AGD1YRAeR+44LC/WKMudNUr
RdpeVt6LIhaRuSPumwDdo8LMjeuqHrVsaCWz6FNxSfk2K2MI2pWqJYbwsCdV4Ni8rFxUrWnsiZpe
ogOBD4SibNdHxcCMepdpwXr/7Qatblqbdp4c4YhcNgIRYVcVkGDDqQy6lJG2wVqS4MmbBrg6Gt6t
5bZnebNk3C52S8pHh7WeCabM6xw6Hxvb2Lj1jgVybiqeOOwXujAbKwZhZO6NaAjKDmDHnTUJwoza
QQGqtB5MfF/qCRMPZ4Gayv9e3JgmirsM/9tKdsKleQq9bmDNE1TnQpIzI29Jyjseum0go/hKCxtw
T8LQA3ZgGPdvTO3L+J3dsgJSll8xqj+5t3kwR6J6iECWAbh+gRCEJUzmAlKt96pZ+f9C+7KwBIfC
8Kp0JvCQWPsTEMGcyAttX3ReqNrcLne0ZsWu3izBMeXcHL00TM/L95+VY8k8Tkl241vFxffz0oRJ
FhYyH2ShVU/RV+LK3YAJ8u607wf7l7HVpISgw6C8usc5UWtes+Ywt5RHxar4Se7bnQU/wLxOHlFU
q73o5RKcI3s1DqANRyBTxzpazuJicWka7rp8NPXcKMfXEHQVponHFcgPUTdGhGLN5Kv91r/GeZTE
7RCKWO6Sp7Bjs74Wy9w2+PXw0NXAI/+6mQogMkgdt1DiU2m5gR1DExgYMyNaFlfWyvHOaiiBTSVQ
LuTXgRBRIHv5D76pq1Kk98eTYx1udHDPjPKCF8fwY8sS0mAOWP5zo1xxWqRdDibmpZ34TdXh0k/x
PULJW3UHq8Gv6CzT5LATCD/klGcmU8CqkYUPreouKCl5OPtZfIgoSagdrMMYVrAocVDUDafriv9q
5dCQO9mcf7shdtUnJ88KNG5NJQGGIEFMHH0ViasxrR2yHBSoG5jsvXMWqhynSglgnwI13kI7hLC2
Ik0NrDXcCyZ/CjNi2IbSwJ50RqDiKw3jN6RxUBuKwI2x4SIt6/q7CbdYHqozeqhDdWEW8SW2Y9KP
kyGg2QYuW4sEtnc4PdQxrgfMOP0J2/OIaUst46GUyy+GL+FzMYDvSbfcETxI9LFTSCJyBGC66HSu
9dCynzaXOCJcE+l4It5/wJIMqCDUroB201yOSQC6JVeqfEzE21DiZBNsqu8K6S8lcXPSgpZBWPBK
jEse37H/VpDYOfcU6awO/7nq0+uXpfVuFJjKMNJu3lRS4ODQZu06OAEfybAQudYLnzepKsk1V8co
YkqnhmnleGjtahCDd42YxqYJj1nsInZkumCCYTjAar9T2SVvnjUroleHC3pNFAol6+u6KHPjEQii
M5kG36XKJpfDwDFKvFypsN25mkg1ypgAu08ajz7CTeRshh/jUJL8Mi8SHoT5KlfG1zbTzhIcoouc
zjmGllDLZJivMhFBjFtJxoonIbLBtsi0IaiSTqlRjafhU0yjqJQWM5unM8LIfsazo9I9eV35Bh9K
JGGXhhmbx0tog4hoeyTQ1tSou3dDaBxU8Qc0GLR75UGGJDjzrIQV1vFSUCcC8tHdy/zQazIulSJK
1FgfG58dP4RrkceYFqFyF9no2VAiHaZjxuBWFZqwrDjB8y4tg84THNI0GSZBSLycUUyOIqLzw9xe
FY9aygxybj6wh2WaGF91qgYnhZLAdsIi/JBPbZqeBUpUZgu9MQFsRqBLHZf7bhpkzUyh1RFwZqpJ
+HkrFFmr2XK1pmsfGsq7AKK/x3tCauTSWP5KrvNnG1cI1Vg1UvNMICyixrn6NaAxdftigQpPmFrh
JoZye5HGChwYv/tgsM0U0qo/taAOwB5KkX9FR6BKD45UH2pnH/eDXVXjB+X4hQxNvmNXQDFr+3kX
8c37uKZvNyjVpB4IeqTDxapo0Zy19HVXcZ+6loHqpWwL8kJeaMGl6nMA3lLID3mp4QtvDWJVQ02I
1RWHsOBtgTdzqTlqXbv9Ey5Rm0Ip5/Vqp1UcbRkYUDileulCuUt/QpjYzkSd8RiOk9nDiVnFoZIu
nBMpuwSUBK1Ug19u4Ltk7NB9dPgqUqtcnuPjeWOcufx7ULvKUTkkVrQc21vIRSmqSrjXq/NcpPr4
ey0VRv1FlOh70SR0AG24zDphI4P3SlljdFflAuZYQ7/ucryocyuE/ZETg5s6UtXcVoXk2Qfg+e4j
QrcHMvjAwkahVcRtDyYsBEhUXxiOFTI0RK1rSDXybM+mWNYEjE/gBmHkjyMC64UR9F4OjakGCS2q
Kw9uksNhlciY+oWoY+OTP0UlL9V9dxELYj63AY7mLLnluDl5zPWJ8B/yHFK2MIaIl6o1So/0cxRw
uBMbgDsmyvGSLvI4yc7FV22pTRdT2n6oLgTONsWi44jbprwGqRQ2qUR2Q4/CQ9ixEj8K0T/kAWAy
B5xHyrDAyDoGBTuMj4WUvEp7KfVX5ptMoqQ1ltTyCNeyYHHUxEBgz+DNVIdhZeEapypuYt4B7t3f
1fW3CbVyzTmUWfHoQi/xLW5abRTrrGRN3bNpDBHM5s8rkwoNpksvbnjZjb2zuFMPsM2tUiZXVM0l
pVegbXQB9Bygq1OYHRPum1p5EKnmITb5tGwvDp6DyRQ+vKkHDJ8LCGJCarqDjGAX1mPswYbsLXHz
7L2NSesMo7RzvnHTee/HLRvV/Wh4RJhvCJ3RwM/BLN2NcdIJBAjNcUpMTyvYmlKUjOIIDG3ZQumT
riSjTNzk19f8F850ofVlzjafZ+wkNDPcFGKHqV4rm3TMOenOfTXFHX2pvJM71KNcR2YyVR6A7S41
mmWA4Ji5zxoMJUD1N9NfoKCaT2VhDxtdrqEFORZG33dEP4nWvfk66ClA7asVrfdBECO2O6+jQA3s
qtk/BkNeoE0DGHXabOS69eutVKc7LTSxgzwVUOZNsO3ctGVilf6uAo4O3gGMRb0JyEPZy/iyLBgD
GNVcND1WRhcyjsGD8AZtu6gBtE4NiufJSzJ1VboML+QMKShbEUB+gTNJOzjrS1IjE6xAPUEshL+2
2o2Vwpw21dKt3KPCMwFz9rgVHTCASMOvvOilVEkPKvJYJw9YeOhIMGXRGSxCBqvOn1nSX9UXzCDF
qez+weVN+069MqQnzcQz8ue1voOxINRHOuTw1zVX6GusfGbWBHKRNotr5CyTGoh6sFP/LmK9GpxP
Gj9gbkbLQn2g0CkQv1UPAAKKDy4nNaQyL5ZmQ3/xpJOfofWPhcSl3bfxhTNk2lXPqdraqaDl6TQx
8CfAbKE7Gqz5J9V+4WvVVVZl787WAu9LRzNa/rg6/67Gy7c2Ld+5FXeecthzx8688DRTszFRd18+
K3YLWa5WNBmkQe5+pnjRBzxfYxB+NRIpe+z4dDHfJhBhiwv1OW78JR0kR5Uv+J22RDnWliGwGvrP
f6H89Uzi35q/c6DPKFWGr8pSgyKQoYk7zI2iI/O4WTXP0fefwoyjMBPtcadUX3gMpYBe91Fz7q4c
RDITthO1f7PJeRvP9+sljKaRzGbf5t7N7zHkC3wwJ19/7YwMRwwV199CGAOTWyvRkkZz4I6P21mb
ILsiWSvK96YDD4ECqcU67ZNoFhUdtv2z99yyBwWDEydp72nHpiHWWs7NWI2iluQTe05vWGTZ0EnY
T3FcJVgt9piFwmJuykY5X/UIqBDYxZBDYM7UcC8buJqjtDdg953VWp+mGkxr31joakbITs1t5TqB
TfvPnR6iO8voV/q/xZJYPeTeEpnpWRl9HC6g5f+HaWqC3Xreuo8djtsUKoy60RR+xhf1snaz0OjQ
npUs68roY9eotG8OWyqQ4okgdo+CtFdt5kZ/UqZtNpq7H0AOGi794S3O8e5ql537XMEbU7j8weI3
FKR1ZGaCuNl5Se+LR30ZdRqBhMp375LHJu41FxAVd69VFpeBHX236ygRe3FoSt9HwvU9AQ6JApBf
EFo3ziBSfgVFiop8bW3HdYl9bIU8q5GJBT85KXINWSa2FH6Cz/GZXbj0ubEWLn2idu4GMXRGB8+O
C+oufkSfujd4e4j5ZHDM3wKFhsKKvfY4Qfx933YoAFlV9AX4xHLqY1rD26wON2cRAolx8MaJhDxg
k/Ao45Cnr2PrI9vE2RtuG/4RNMqttWvItP3ZAkPN6DZz9QDyKlqIIoGJgnp3sXj6lx7WSVWb+1TJ
8/RD6e1tTLdRnoeQbBMzXNv1GoQi0ZxeUkB8ZCGjLb83qrHzzi9peTgxfQRw3X1gdHyt3gR8bgZj
RakqHNget7D9iTqwpASo6NRoI3jzmSI0dyo50O7RU0D7Rx5s+UbedA0v6esVCU3rQXbaYsIkhtMo
FcUGNRqYCZvYuXuDQP7WEYHmwJsqIRx/dnZoXo5+oeoYY+PF3kFly702TzXO78m7C4OLVRdEdrOq
gSx/KETOFgiZoku19mTT9lvBYxtH8IoTb8dlZuxQpIAA+mKfwrXZumDA+590lzHTIO+Ypmr6SsIs
JtsqblVxNMtph/Sbg+mKgwWwOixKwEPaf4lI8E3GvwgSbd1e2jAWxBwM2LrLyRxz3W69J2BYVclU
XRvPsdkQb7CXj7Gr60OTcf9EpykWDAP3LoL8x/3RbgVBevp7rgnkYq64S1R5A631cgtYYhf3Oq18
2xt7uoY689qaij55js0fLEqO9AKOh2ZeAEfmQ12BmpSvKqxeOvOmaaZazAHn6opljpzZCKCFbwon
ZJ1SmUxy4Fkje17naDdSoKRVjQ1xL/VqchQxC0nEUtS1hlTEMEFqnzyU9SPnhC/m7z2SysccEpBn
YivDLKYjdeSg5itbYl5VYuqmomERsuMxUkpg1qtI021F5kfIhVjldxSA0hWH1vc+jRr+aT1/r1j4
qVwkz+Ek4aDYIHXGl+CL187PZRoPpFf4s8bEmn5Jv9x1VlrvkugThY1n+B1aM9gVCbPyGNfJTJDS
uys4+pivk4wfOYwMWW0cBauNcj/ozBf0lFEAPyeHpFnwVGaFviMcfRWO9adT2G0wh/RvzcxmJRpb
1lFbjSoVU8pGiL+UXEnOoJQntf1/1yD9cyp+2JL8BPcAMDA8KmEXhldpWCtNAmGn3TSz/NDFLsNN
OvNUaKhgWax7tjY+vPLyIWXiJR0Pk/3gz44umqDSx+YKl04wfVEp/9zrCWqXR2Ug3K5o76NddpG8
ItR5V+Ao+H0bLm0mn8+P6YLgRgtvxzFAWvs2ODe8XzPih945q4QJ7UliSghdeV2JctC3hc2VydWD
MoWwsw5s77ZvbmyasSZpW8q9CzfkrnQYS9JDOIpFlkL7ApI8Jzbm3Q1Yc8NZWZV42GWNZTn4NSBM
Y2Vp8vFan9tjadJqq11kPFbPa+oagG7mArZmxZlKQxjHQyfgXxjGCn73u/XyANt41GM9yiFAwRZI
Xjq8wraLpCrT5BW2pkxV5nRbQc0vF3JesteODg+O9eq3s36mPO+dpig3HaCw53h8eRB+adVgxcBO
Z5kSSJ6oTqHSbLjo2HjelCN8H0514/RfqbKak56cv1ESlvY+4UPnZ3m10fTBO83IyOA6I2bnxYlF
mDTmerjep5KG6wdqEgtXiheZMKh6yr7kI+scWw0JXXHE9ugBdgI1sKMEkiUiKn6XqVhhbO19Y6Pq
d+L+5nTpvpAN6ewPYc5yPpkAVjcvPH7guyMwX15P6OYHnbrErnHbrFLA08nfCAA2JgywvkH+lFSd
xX4Ab6M1l1iOF2inTrv6+r7JXAEFCRCbB1qR8WkOEs086hHXbLgXQqmxInIdLWKEIKVp6OcVkXwu
ej0QUaAYxJpJRpoiBPlaOoFkqVM8g0mx4otoAw7h1cHJ/E77bHPzzWMaizIyDhXuEJYyo45cBhte
deB/SMecROTqgLk2pBibG//uwY/5HMsjYMBccC1JYDdmll5KSKYoTYRQsOUce3+Vxbux2hYWa/Tk
FEn2YhjtvsdTC74sZitxNwuvd4AmrXiCqJagGO6za19Z7cJI7XaQQkBFACuQ+rJHDW5w6zRfX4BF
PjLZIsH46cXZLRHuxNVRvGrtXLkti0GKOFTDr+dP2r56AwsoWpTI2JtgbxWHhHGcMCfdrWbAcwBo
WHozliBd8lw9jXhlcSybhPGoTOgC4B6BSaYlHXRAHa0iHF7GP+HCLAlqHmwbfcuRJal4OKxRAItZ
z2+IOE1Q74bCQF9heUq1SqnQNfIVx9ajBtnAmru90exhRcgZ5BtVmhdeDb5u4YmCebTneByNn2L2
8mktTQ3tlMrOWStI0ay0BncqKrykrrgMhJfB7gEWQwxJkwQLe81EPd/r9UpuV+ZEihNdax+J88O3
n8y2PNORSsNpCX1Uf6SePO0S8Mn6Pe547KP697t1Zrh1x0pk/gzRCT4Imcc69mnbpHUjfHsvbGSU
SRUB8+U0Xy2L3FA7iGAsJxRzsc0LH64unw95LBvQNn8pQvE6/3n4A8mQeZEx93bB+LmhAUxGGs98
xQPTjdpob6oquq+DnBrX0qEwhUnE+lBrtI0EPerd8ScplwU+wu0+5LcR8ZCr0oAjWNN7PZrzKK0/
PCwQHisrpcdWhCPo40NRFtNo/fqCCmDnxYy/hC9IwAbjMxWuBrZf5IoLJ7gljcFr5TmEl+1U7u2N
Ymp9OBY5IMUHO2/KvaaH+l3IHrPvkmg+I+1oTE6ikdcftuXhsKQB9zBGYDoZv3L8nFFH2msv6jDx
FMJkyS3a1HyO6fhuhs3XJRUkxHMw+8R5JdcT75g/NjReN0+HemSG6Fr3MlcQMszEb4OixC9EkfJn
0ariyP5BkS2ELQTkjL2sm7DkrXpxxMArjFEIYsKG1PbEycsE8VvuqPT+WPRpdrTCZZJjw6FmyDvN
CrMNEi0ZWCcYJs+HZJWRoc/RjPFo6pP3bn974fhH1Km4tJxZ7dY2nAv63JuKu11VekCNKczQMFml
HI7VGrZQNgukv+DangC5jF7FiYgqQ1WNF5sy7rXL6HOz0kTP0pfI9wxi5ZEQU+RWB/ZoMG+K1Wsa
oNmlxhRBdPZbUgdHtnzmbiDfjGazo3xpHk8CZ2sAGwXKyezWfuADUkV7OD4Ins1mHwBDcECa6Zpz
Yq10PaHbYr8hyDOvE2oZ6ZcuISDXRHJIhuypVh7YWVeEGxKwtHacR+RTRedX1+cWEwsyIH+2Vk7t
Sk+Pwryh4GqkDwPSRMZBoIhz1vBbmgCdPp6blSSM3LZEKdiC7oleMyB4tSGHwkNInu8ODIEsDA5I
RKGzgT1OptoM1L6YfY/+gWgjdrldF0Cn6HkWOJ9aKNL/kzYjynQHRAg/MexEX+CoZ6mH5gtnfitR
GLwy/kFo+WCsM6uswL+git0mKTy2UX1aYDCmFx2F1qPwrK8vsE3IFn35fStxD7rvqK8Xs6Cppkrh
418dMPQeuQDpk0Jprc4m2BikJo+KdL5UfEX/s41fpNV2lUiYvr4eP5CORPBaTekeKQ1eWOmxteng
Dx6/FJH4tHnsE+27gy5dzb4mkkfzPO/aujaGn1Ifi1i5x0cdc8gvpfmF1CdHRbz8kzZ2OZE25cb8
+szX3xDrv8O1aLdhdwUWQiEckaGCQdX/+5GsTut8++bylxSgOPuHgYH1ZX3F4e1TvdWWI5mwyqm8
2U7XAdJppK2+u63qxAwGxr9H+9DECIuFl3JPJOoiMNVaz8ojoKgJ98fscAWc5xa5jNSTvBSvxchx
cGI7YtJKbrYvF5VV3l1l/MeAV1n/JFuOBK9tp6KEkfFjzWnDZsf6+QiSPj1l69WrxxZK3pK96J9c
hLjr3zVoNq3ba3kILtiK39bESF5+le9CXcbqFaVG2Zj/kyZOXLkxsq6yG69K24xCn6uXvon99GdK
m0f+ag4eorJ91mz39Pxv3UE/NaLvIlMOJKKxQgXghEn6Z7+x2wyDdJCtB3CvzKaE94RK1OdASlpb
yRztdC8g4X2kynFot3OAFkktghiUxEQcMPfOrf2Nvr23Ycd0rkCaj4oBM4utPca501VYLCV02Tf5
fzTM7jNF4y+fO6rGs4P//TlpJAiaUSQoWWDCWw0cc5twHDrTQxZybkQ1xEgAVA8K0P7JXBQNPDM5
jd+igsRC3BBIzxvYD0HBtCWgg5+NW7IDBDhlDnEW+vTfijBuih5Tnf4Tfwtd9osiLthIHwQQWL8F
+flClzv56Q4V7Oe3IXYGPJMwtLrD1vM9YegyJfLiWMdEJWvqNzmgbk6cbDGRZIfqXmXtNPgD5xEo
f2tgV60T/FRFK5fUyjYdAj02KAtKiw6Hjzp1I4ik0t4HJpFCqQXGHXbAgtPi96AxQgXDtLv3ZG9c
GiVa1/s2+45ts9OZ6BoosyVeLV7kIh0RY00we0rC8ARtEsxgMPFTJSBKpIqkI/3aNmU1oNTdJEJZ
by4Da7E9wbP57IP/KTQ2F3ysA5LNJxySJrwKZaGyyY5h0kmKUpTWjlo5V3gSp6lrEbyGinT//EGg
1qOz6fDGKErlEo/K4WOgULAP4KlRNwLZERBT/1yCdQaYFtrd3QNAofCvcMuUgQ4hhXREL6GuKylH
Y4fmzrIXbtIVB6MtloTWnNCTJG7+VmNCNmk1tWUN8qH3WzAefAjPjbK3bvXbjRhQfWxjXUggaDjl
vC7a9nNL83cdpEcXy4QCL1oPwCD3Q3GwY3PmaUukZIZgpYEqtLKnWRKwcGqHTuwbOAZ3q7BFZ8oA
1U326HNvS/j25t8K/Nu2ri5Cj15Mn87WZ7zhyceulXqrIkDoaFpnsYY+MlaApyeg7cyxNnI0ZGtP
AaY1gFWWKL+1noyUAyXrd+4+BxOV9ybYpEJ5DOVZ1O7h5ji2m0EofnZ+JlEgIs6YSJ5I2PnINu0T
rxXItQHTdSU39M7yk894mVX+boCQjdR52zueEigQRU1mJEPj+qY21Y2zDuVgQlUDQRzrTG2fmvn+
GVHXnKFSEM3Qr77MIOfg3w5WNs2O/nN8/wEE4wHESpCbMEi8PVPc/wLvQBtu3QT5NGxi0Zig4DVC
FRo9NuZFcIkOiW7Ci9aqYHn6dJx1bVnDavVirhaNcvIo7yWmi/8HufMMyMG5GpNJkcdqhLUG+td6
Wfl4MDhJOxR7MRbMRgMxPwco4o0UfcuZ/Gfj9OoXoqoEAFk55NhUfpcYBuJ2O2XgyTGq9bUDEL00
wbLc32Qa4YQXCc8bGg9MGeyq2GLT0ii87aR6yqUvz2PyNSgPZGQpPkZnNDs8tttbeMP99mbpwU27
Kq0idkv529lXrtYNEeeGYnYwOdOivDF/JGfdbOilkVLbXosk/kNvDn0r25MV/VefA28U3Ph2djBy
rQk4bKYaoG7lF+FDJ2LVxb/v44JDbRLhvEiwV4R9xJXDtteQfuqCaFHbbbh0gOKBL/pWAzzylMsc
pZBLc3gCp9sOX/AQ/+N2Wn5fUpPHgBWgVtSXas5+ltcbPo8hBYbEtb2ee2Taecm3GfWtgCaeZb2a
mRaShHLRgn0XnpgJqYU7E6v7YoR1eZWixbLL3tfJbtxbseSuX1GiR+HWncp1Vst6oYT9U5VwrS1/
ZyFds8pGdHEQX5G2PXZb0MGlNc6KQ9RZLHApuqEsDALppcPGG+tN6pWMEJE1JjcVwvAoAs54cvQ/
/bcqaoOwNYbFZawJRoAZyXDBo5PHtMllr6Vk4ayawBNA7qdkIGqaVApBhQX0c35ZNCYLp49A09hw
4ILHNP1p66Qd69bYaaobD++aztQvwFYOZgRjO+tf0XJ1SFhojwlzPoGo+7R8ebHgENOmBmZGpIaC
fOB9JHXOH+Tcico2QR53jqTm1Qi7R4n9iub1LLhtngE0Db5eciVCKxv0D6wF7zrcyXQLNLrLb6mZ
l+jeh9aiemUEhP9Sb6swcrnW/A4kq8DgY9NqT7FTfnPVtPBgtfeA+QDQad7xMEp/6j4wmLpaq+pp
8PlTE7aUQy/qdMV5z48Zxi9g93qHXw/qAdCxKxc2eiyKb9F//Myvqp79HZLWbS4F48e1CUSt7SfF
ZBbpKNPfREjDvPo7+HJ0+STEL9Na3plMoKaqUyOx0d1P9e4M1NRva+GEbYTFmIroVzL+vAgCkRyn
Vpkjw89oXYcDxsyPYarvmYDFNmKat+1WmpsCH+qgr8RdkrDGoHF6zLeAnI7kvgKDdlcMdBYockke
5Jtc9TCRKw7K8cd3EmWM0KJNj0s+9F3nP7DxHSofctUw++Ul1C/rbah16jCWaqcCLevUe+Il7u8R
J/Ndv/Eu01QuJeWHWI/a6g69OzNtZDVWS0s6iuySbCG9UmLiVezzcjSYyv0lpLwUVKvCeJ67Do6D
JY3nfliGRzArwI0gxBYg9HZFbtQ+Kt0dh8pOI+inegHDVbI0Md7/5aMB4F8QPZ4a/fe65fP3q9x7
04dF5WGzq22aPLgXWu1hWigjqr8kv+u5fO8NtIG/szPD5kJ4nvQ+dE7W+FMhPNfJ1lEwJLnDnJ7l
x6Jqptr5YU0nHYXUjADC4MGCEbTbCIHS01XPk07fk2mO2fJw5KMWBxI0z6I1W1I6/y5N0cC57H69
yuCKjnvP/gWXun3+4IzThucV/n+a++HeLeLeQqycYUH673jS8Lm3o0FVnP7IbEvE5L1sYh4FrIrw
f6ssHNmzudeQHRjixbNiH/r3jMmWq+suQCUrwkG1Fk2qBkLcygc4s6351//FVgj2SUCdnIq1GzAv
t4YWyIlJGipplXSoYDKTE/TwO/LvX61ii7emloOUW1EMYJ350fMnblvP5VrblAHcItldYwg9sK6d
BmtQINfDUNEu81P9pyODZy31aotbRjVA0+WKJJsnUbUFW+DEh9GAia88Og8tuj/zN4UB7vudMdCJ
TrcyK/UpJVE17KNL60jWTiEU3jzU8RLzJ1wnFBHejtsnS5Vx/lfR2ehlySJjnrz+eZSMy/36li3c
bUrDjw+h+My59HDht3nwcqrTVjQEPASCsYm41bOADyrVkZjHf9jOOjNmuJEqOzutozOMRbWI6HIr
1PbGo1e4p23qBAwplg7MEI4LYwxP3G3LWDm5YzC2UPNOzUvnMpzUKIsHKGeFSTqUVH9MT1mVZRvE
aqCVYh1FqXwosyC2d6xogLaKpRBKuIzOycWt80TrZFF9Jbj9aINBPU7NewsIrCVawii9H3YsfHRW
ul69aFwGs1kNMTDJCxm1C5bCisi5zIVZrwlOA2WgTNda47vAkoxFscwnTVNob9X0JlTSV7pW83OH
zE41lrY+0H9+z8060sQRmMtmsFlv3Mtsmqe3Gq1/KHW4gQoltxFIBC8CdV5BlqIANwM6QDzkL5qQ
8mVcbzrbD7EEXx00efWvZukb8dQ+PPUQIAMkv6ST6sMcxyq+jzNEviGrpWz4Y5XIBevap2Dhqq81
yg2V+abGouEk5k7lEWwsTJpvujQHZqjhYcesrCKk6J6s1KbnvdeZC7tRzjZeKGpEKMn2UoFZwEvd
+bmgz0T9EgzLv2bAFoPsPLYAKnmaIwowmw6UaJCeiPoKGELvyyDfP31ke3THZdcmIEwc6ef2iy2i
YUNkneRCLcuPCV8a3+kDTtl/xuNW7pz1+rNd/vLE3+4LnGmGckmCuRm+1VQKdxpo4JvLkiGSsXMy
RR/PguRne72Zu4JPd/SFWUZ2Y6DFv4pSBGLKfirsqEcC7ImawKj0US4+fWp1awsmvQezDIrSVyRu
pMN5tnVMd8VcSCW0jKu2QA/joHvt5nG3mQBlsRiY1yQ58IKI8m13jUCXf3niYOMs/9gM723ro34K
xceZ+/iXVq7oAZW3CDsKpDiG0wpOYQx+XdKq+hJZWxwp9eW73IU6I0a6dGgs3iS8Ukg6ROSJzAfW
1pXLE+pjje3sm9SpNO7kNOlbxrbahXBfzhthA8P3JSlcll5Wmb5aVV3DBJz/e4ZBhWFJPufrGo3G
EM6g25XcrM1Iw4urdg6qP6tQgnYTUcL2h20jbmo8q7O0I8qWkp80ENBUqtht0I+UqUXItUZJJl3i
e3CfTWMpyTPs3lfT9PxawaoY4WNbqE6LM2usY8E4TKHaboz2b4FpSveqx6/z4Jm1g59Qq3LQDR2Z
hIzoQ+2KdVvbvBEN1cczPAV+JHccM1DewOJ8uMNNDrqYSbBeBhpOgVJOQcdmHhdxKdwS5pdREsDs
rh0zPdbhHrMV9U87Onm3/p3vfgQ78w+aODSCgPYpJE7lde6BINrD++sTjp604L6Xj/FI8a6zDVhU
WluoecoPIVsiERLBXI5PAj9zEZbgyopLBIUWmC6nR4RdanzWRXiMWfJlB1GsQJyAEmn6gEz/C2Gm
zpU+qRXlVjDo/NLBhSXDu3cEmZ4ZU3JCh096Otaz/xB/x4ps7vPK280s9kGdgFfjnWJOtAty7RtY
oBzCdhgi232tRXZdNdSJOZXDuTOdDV7HAWVzDJdoaCW/Xa8aZ6+xHUjaOtiHjThU0yzixuWJJt7h
0co9rp6oeJxE31RL58xf6FzVSIko9PEBDJmfm1oYmsg3x/IFPr1MhKKmeaJqLGSErMPctXuNQSLZ
auyS4ADzxOtIm5ulsAZKkhA4inpt1anzHa4lvRWgYgLKLjHCdr2mWthjyHE9u27C8yj4My+VCjFP
6R61oAHxAyDhg70lgWi9xS69SUanrvVO9SlnyDHZblx2te2/rUiezUmn+CdehvEzS/VG1DI+Txkm
cf+tuCda33Xu5VS7fX9erqUI2ABaXdz9VDTaWWkR9YDYy93Bw5pL0E4t5hTnGqVPEmi+9YyJ7yaH
ac+tvVh9LTcnkuPe4bVDLxW/UoxCoSUX4eimR5nvzKXtdCqkCyPaEX9MGmmdoVObmLuRJG/uGSlZ
WCT25j7F0E8WEcqXm1EG5Yp9q+Ouq/kHxBBf9bm5LJKmpA54ufxD5Ud6FDOikMhpNvIXnFTm+Gld
zAT5XamWEt4GhHAbAG6oULD9P/XKXbatIYMsMWjdG/ATuCETExdYxfPuuJRhxKXviGnp2WtJPBJ+
88hpx22l3uL703HcLb8lR9/5BJaL8cd8HmVm4VU+4QYQVjCp5d/KDme/lzdXN0/+vOSIj8r4tw9/
ZV/bzCdF/Wdp5ixakCkvwP+YAuQNX6nf4NqW8dPbhqbU2Ixkyk/9FSHPY2IjiR1XkSshBHcmZiCJ
DFVI7lvegKrbxL5VJM1vCGYnQB+dnBtGVlgllNQzglJRHNHKr0vTO1ed33EXOlVsWysx17Tu9tei
PGRPjQJk72OCgGQbeeuOg/CsqpFutGNTEwS+aMkwWsgLseKzsZZYTjgOn1S/DySg0s45HOkN9SOD
1yLbZ250LTA/5j5KzF8tTyEJyZ+NmoEXQNFuEm6FHNKE+znHGpmS4Rc/MtJuYoIXFCJnVJEq6A/h
RwHuiNrU+sGyusx43O7sMt8QfFEPpILXaOGJiXn0Cqn5xNaTwEPyoNBBaAS3xwd0ecQD7Beh2Kme
rUQyBIiBilWKukwpvnyH5WWpwywF/TTEkt6otyszsb81SssI6z3qDf5wVv7NKbaC7MpwiBhNRSjp
m3xhNQE5U1lOROuWvIBFrjRAljMnKy/fJXX0/xoAuPicu6CBSUC6kRQN3sq1Vjt+XUsLTeYkKJZM
qla30ivO9tpJi2iAsVrEsq4eQPgSb79csu2M56YD8bYkW9+Vo5sncPh5uJ+RypugS3hw4sZtbo6h
n82bj1U3E3BUsAtDfCY+5eGxnCnGjSjugT6DHG8XmVk3qpXM+AnAveYKdGusUHCHdowJOgjEpewz
8qKZLV7iwsBYmI6JXpaJCBOTYdJtjIDpCYe8iigG3ZemKf+K8TAvqJqZZPmIvIg2+7ZDQsa5chAE
7rdozgN/0A83d+VJXTpy0Fzi2WEAmOu+7/C/M4IC1J5gV+a3/kQJlNm2nLWMBT9WOuZHymE+GcMD
6ys9/ibLztXToUaKFBbyC43b1yr9JH6Wc/XhRiex50PNE3sx8kCHjl69mup7nRft7y66EjI1ex0L
qPyCFcZDuFK1O9497Q0BFVgkUjnqTKt2S9eqktsVuwOkSse9nLpmg1m25seIs6OZv9qcdWk1lkz1
KSy1Olo9vQ3D2eXJ17vsHXVUCBDU8NWjbL4u3fjKbvRuNwCI1xAWDvU1J8njDZS66xrqZd3J22tv
CDqBwZ4cmCTEaB4qxdyy+nnVd6xI6JjxMNqR9ZE/aNL/utQRyqicdq0iSGOY/Tzi+jnQQYqWFWI9
h7nBxRKUNMWRHgBDxJYKgq33FYK8pPiQxqtPE7Nw9Hcu8Pj2zkjLpN8fdfF3bN5tI8LejPiluPMd
UsVXHTrC8b85AzHyRKQXxMomPt7xcwNLC8mqs3KRyjV5R3dllubazQ81+YWpc7K5OPRSgaUudHKr
SYwM8Ll/FIHItc/g51gu+QOh0KSdpRIB6WVQFl1KXbGuO863sO8r8k5wWuyvfZRMCJdietEatuqU
q0J21pJD7+KjDXAocAhQ4GPhZLJ34x8WLUrR9YQW/pWjvnM7Ao1rXhRX1rwUBGB9JpcQaVGUFiwy
NGMWSr0YauC3edq3fOIeFT8yNisOg/0yp/uPed1zbyica3Mihq7BfnXiJaBZbJWv1r2HC7aLLopk
WPVKLhW9xklXjwiBWZqtYc4Ha1P3dHhxpts5HvPedoe3wV/jknhIOtYKKsKHj3wR1l+Uyg3UiSi8
BuRfDiN1maHbzSxUrCyldCyYhT0ygNaOQPu7QgfV26wSbJyjNt1UnaRbA/6UQ12JJWInXLAsEs3p
e/jqFipPU3y8bX5jl2LP1ghW43WJU/Y0/mN/Dj4icTSU5+iyDCCc9ITrv72Kh5ZyafunvSWc1qU1
+3LSbIzMshzogt2klXAR16wMdEcupQMmDh+hoxy6SpOOlq1Kr+fRLs8ykr8yZ05P27G7PGHN9/VJ
3hOUb5n5pf5GlIYO2+pEPeCOyPjsgz2pZXKPy+xiLXRBEY6JN3alfRrhqDzEXxD+GtgSoCr4smZl
+QgNMdXwJ9jJh4BsBqlNq1pm6ZUmkVSfGCzJHj5aKH2+O5l7lEOGLaNVI4y+OLiExbJunfbhQaa9
Gj2qbyIUH5fF33UH269SeHYzq1DXo2PkKHB79bJ0MSlJpILcxYKu5PZ8EDhrdkHteveLnUsLBJoi
dBVPhow8EkOidZl1us4GSHQRK8L4wbknKUma3LcWvRtGK+rDBh5b1UmraVv2rzaVe/HWJGYWhvGq
cnZhE2xMb9nCSWkiWYuTwVF79hlSGBVSl29HdIZLoraFEdu/8AkwK9Yc2kjTJq2SsBdsVZnQUIe/
Li9s4ymkTjpUoC9oEsnCpVukLFl7wqHwgHpacN+7Sgnkz82HY3aPWtBvt7L36PSmPgfPedpC10Sz
RrT/Xmy+Sp0xM7kfbWftNs21vs8f+DqQlt+JHCQ6jVvX9via3/JQhmXogN72Bodzw8KHSHGShPKU
Q4r19Sy2gaWsgPOGlfT1EmWVP35RNH9af+sL3QoRb8scvyf5DEjTCqBpCYYBHSUZjXgvZ+gm0YsY
IblYOVWd1dxsykNkk6TN3n+iRd24DIYCukdS4GuPe4nPMsSlYpcpffo7gQsIjVGQjKJvuiL6zLXK
8kQhdVFQnqte6vFC845E9AdSSv73Md7d/nxOC740pwvIChawq0zIET5Zh/yd7eiRXPsX628GA/hA
mu/aoM2U4rbVjgMFxnAJEt4Jdbsv9crt+ue9AEneofpn17LZQIUKAsTSjFeq6pWVpE8g96tW/boE
NJV4dAKrQcVIgAQULoku94APefzPaGEtjw0R7t9BBgArExFcn5C6hSZm0GSz7OtZLW/8eZoIDxSZ
X5Ock9bcIwkXu6mckHADrDfcTTFN1VQfkJ/b23zBA+SCMRdmPeDrhBQhOc44K2Xo4cmeAdSA+Oxt
Mfh6XvcRolqnGjlfK/geCly5SfLrSTM1MCDP2PFkyn4n2GcMO9CzORYTM3fWCGtUzvnzV6rDZLS6
SEOAg58u8PMTSqH1+qnFiDEklviEsMOZfpB73c+1r2ppnScZPzBWcu0ge05yGWdFpo6u3sjcL3C6
8hbnZtTbbMg2+nyWCfyQkrx7dR7w7MBRtkZZaxn/FtP9LNzS3rVvMgdB4kauSg0ScI/HHNVlvzc+
rH9zc7tDmPvgR7ct7DyCGV1jJbSaagD3XfCY09Bb6sOdRtLdck1oSIQSvRr/vapz7qS+nQVGVsH/
ZhpJdwdfggg6TgsjLvDkG90AgLyBmyQZIQnaSoVvT0QZeCb78Pu41uUPPi3NXwzz4UNq3iraUhcn
2QgIefjkFny5n547DusSUtZbHRk54ADumeAp4OdIvBQQAhK69NXtMfV9Nkcg4j9x8l36jgQgLv4V
tQjy9C/JLK2c0AZCgaR9fwlvfL7ooA8Zlx/Ie4nsaMYyNV9sAwUcxMabGTEgh0S5yHv4rE2FXDB7
6wfrBRAPBQvLiDlaX7tyE60Ds2IgIcWv7AbOxwoJ1hqD0BWVHR9YPoFZlLmtcBu8KdyJ7TrThBdY
QJc0DeeuvQw+eSzV968s/IzFclsmANw4b2ZgtXm/fmRT6jbQOZ3EFbSJd+oTTfB2r47hmq+B4QBl
EKNM6KWmBGoJXeAcVnWNSGXFR0Dx1WIjrpuLo4/Rpez97aufbHoSYj1DfijIzNu5RQ4hoxAkcopR
f+enb8x5tduslC5LFrBOVoHgt0BZd3bGvW8elEB2lAht7N6Zkua+i36tw3YQqokQHh4V9ymboDcS
i/CG2guqRYfaYWGNaD+J+MHbHzLXD4uP8GWJ7I9NFIF1yYFdg6m131GULv8tw3o1JRSuf5B+TkF2
uH9yuHLCjrYUOtcghdxC71DqB2iCzavegQ353jk5B7Y2LQVrUALk880Mw6lHrZvG7a+7ILx+CUIc
udr73/+2velcu93zBEfyiytHZVEU4anea3VJzc25j+rFtSPiWcJosrmlvFFDGPcbiqgKNi5CKFoG
1gsgsN7DGowPevJEhbtFVKjP7sx/tw9p04EDCUr1J51PRQKT3aFOHa7xZrhMjyRVGM6lamvbfFMT
lI3NmIHNpYACUnT694xIdMcuc4t1R8mafWtXr/QOroRyglMGzKDQM/ipPR5bjKziSe/Ibv3zSIWe
nfY8ujtKGaKiPBZElk8qVlPEcylEvCH3+DnwSj6Vg+cBy0ANcCxdbBXvxalWPe+g42cNV9CjDB1W
RmO8wUB0y7Ragbr6z8PNhXEAjaKybTh2zqtvEpuLQdC0d3fgj2MyuZ6ItPOwIaGZ9gvKWtif4ZRs
m3GnUlhRo/x0oqRNACRXGhrKRb/cKSXbToMPUW4Ep92jIw9sq6euQz3UrtBV9407Yab4Mexgsl8t
EBi8+kCUGRFYqbvnUN7H43IeXcpzbxLXAV9E1m/uSUcV7lm7G695tEMcF0AvIf7qOLr6mcsKAy3H
Dx2d3fC9LwZTvQaVkSzbz1vDIxdcB8Yl5YzSwoEv0vmwH+DVAp4nlc+9r3JfnGnDUJxqqlWBcB2t
nbqqr778PcInUhu/jeTrwDhlnD8cK2EzcnUk7jtEB21CJ7fL/f9NmtY4cDy8uHVMlassHXQtY4Wr
HTLUoTX9DqrD93HnKOmOep6h9A282uFXDoAi+1UeW2JbwrbZrbcsXcftG8x4mJsWJmY1x1w3V3d5
dhxB+l32GBhqYynaoa84XKzl4cOuQJ8CVtmIeDrXzBJr+wVdRLueJ+gk35kQy20vxIny44g6K+98
2GBfS771uRR5qGMZ6rRgza7faulfBNCoUQ8s9DV0FeQsgFW3bouBgUWPnGUJ0JHwdVcCz+7WcaSC
z2XmBhRxPqY2mPcK2vK8CGi83MBPa3wrrIZau12TjMhix5HIAtkvKZ1+W7BDTMaUI31Z4x5DRU7d
YBdedNOWg/Lv+84U3yfDWgEYubxETOHXNnhy7sdF4bEyRb1dQxPl/gN1FgldRXbJg98re/6fwvbm
duR437+Xrq1E85muy+LqbfFK00iVOSFS+rbUf+kjVKrIpQxYqPsCKZs7BdQHlOoX8m6TMsCmoYVG
pF2O2K8ERhTXj40bkhHMhx4fAsMktgHheZmoLk0oxLCAqHFMx3p85SIMvt+18Ddzxu5GCrRzbSKD
mjnOoP17vUw9t/qPVdbI4x6w/w/W9wnHNyP/PtHDjJ0PRij6SdUbf0v/ohCaiYIJhBE0DdnA+ZF9
yY1vfE30metWk7aoTPpTyHNtsQkomDYWQyNNqyosRvjWuajJBzXqMQNcECxKIWRgZGtxPeZjJcu6
S+6SI3BZeaFsWJ+aZ6rPy+PqhVKZAc5YhmUgdmnbe67TcBhYoLyW4gR8aTFkj+2uTvm1lCW3mE74
7EOZ9u0lLytOTiCns2m0Jd967MWDhHaNUw+saRVT+D5GQ5ezX1numddpxXMxuKRvOipdXjUHwiLt
8NpfPK6w+TOtyZYrlndEaCyXvB8X/VzmmEcsXrfqWY3orVwCfuxi0EoggXSk7uZudwo5gBXJIX7D
8ncyZuKNU8vEe2dEWgxzo7xpWbwoGt3Txj75SPKIwPbpRxQxz08jdlG4sq0ppZSlSIzaCzUAz90X
vT4dzog6Fw5LQYTgGYj7Xqj39P6gXVSs4sJBtoT19RHuCktHe+NclYfY87Iq0G0m6V4OwMLHjzYN
urknFdeNgN+DEnb4KEELGbpqCcvaBfMSgiYjQbl/g/tbsRTMnWipA+bd6h8LiTqNgTx6AzvgCXLL
xCePWRFZX9wH1vgs5QajiCAF/oFcFz5CY49nh2Tb+QcUeRe0K4rsWUCG4JyoWDT/qNYr/BY3LsoY
Z4jIw4+DHpAN5GunemKKrtC9GSTiSk8mEHLLYzAgdeUinkS7vIw8Eje7qHogCfI33RgdlZj3jmqP
V/wg85/8oqRCvDtpDNEM5eeo0VG1ZLS3hTMkPkUcftY5NUEosfjwdD0PPmVJ+QhyfvzQ66nZSoDa
15YNF4XhsDVahtSXZLxFa1A2kpywvRWXMX4PuUFp+5zPQAcf5oLJIE0FCpZx9V7IdWe3rMz1qfbY
QgVqtPH1iizZdVdiM5l5GbFHiuxiUle5dNLI/5BlzpJZQt3pzoxSvVeagdGX3jGhXyWJRhTzsqT5
2+8kAn/CVHWOpqkIk/p0FJx9STIbxy2gv7RC99mMLtB7ClvC/kdpF5KLVaFV6XIEaeAn2OYmlaJb
HtomF8iTlP7+7sHgObD0YYoVf//odt8CUci0DGftwCB6Ziinl5wdmCmYX6pm+2YoGmf3ShdhB5r0
ytI+EJXfJLvywh/mkdemlkZKKhRXUBmUkXxsNN29EDcJQkD7W1yfIoT9aENalSGdDzk7rub6RvJm
HfJqYalV293vPtZfXuamEKWwFbWxTLW3+wuADtwTotrXApFLT8nEPvInTRJMUBYFIcVouO6VtrqK
ksuhmzTOUVVMfvdUOjlIahtHfyMb4Bj3NIair8rlQqfoFG4A+/WtJBzNXJxZuo1l3zdea/PShmHz
wh0c9ulMhv29WQPNxk4lmYy21pd7lXjHq+aEE38DkIT0G4ICQs9uLKuko9GSNLdnos57aa0l+6/V
lrSU98ZswdIzDpe3aKfgkUDN5iD9VYMrxR/rrJ29SgCMLeNipVmVIPP9xktZzX8tz6lxm8hLDqvA
D+WkGtDcEtlU7Yt05YhBjEvzf5ICY4W3tbL9Y3BPmlancWJaeOVuN1m+OFV3RW5apbyGzX5vSahG
lSzq20LJiAex1JMvL6zCa/ypT7hbePUF/GGYBfC3Q3RBUFFjrsXn4vpVr42iZDPUfRXz0+RYRFiX
qeR2tu4zmiEwD3kb07S2wA8vKxqSCyZ7reOUSZI/S6R93q7FEYhrhWe8f3EGSv7lrUqzyEGsAycj
h+UX6i6XeMNVd8v3IWylj4+igoGjVhLV6YcSIOjzIfUMTaXkKiCZpy5crzDb4Glvs1sttMISvBD9
sLqfYR0t7gLKAWsfs2eFDzpYYyL2nP9PPplfFZPYwvIf9iyOfsx4VTcJW/mvFonl3YUzZAicFMlv
CkmuOdQKMHxcxsiwpUljPReEkprZk9ZFx1eGRIm+Uw216cDuEzOyKwbac8SQUGRaumlX8qAkXqY4
nAoa/iAcYo14333V3oD4eFP3UyyfVJpuolLypzIIB+UWk9HrbwmVNXsVBTtBGTIBLPkXDV/eUISY
M9kvWb+5G+HqgyjDn9ELzzK8XiDsuZslBUHTXWnkuUDbmElZtupBDz1YNAvZB4BqbtlHvOl1MPZG
NJzVbgIGz72e/U4LEesMkBqeA1TLNNjhyvEE6RxC7p6gcqTU1TPz0aKChC7qYVIleCyFo7b9rrsM
4TviY/PjlcXkVgzTo6sJWvfjUkjmCEzejE8rogVPlSk2Eu7jwiPBZJ8IMosjBUHL6WtlaXD9rIHA
FaHcGXVAMLcWuSt/lFZqW4d+VNssPgTr7I0vFaI7BKpw+sc/JJzl8e9RZ5HolGgSjTEnqEL1kPVd
FmjgXeMuDeIdl4xttAb40s2+z9b91053yjZSCxFtDVRCE8lkeeaY8VlYxZChP1fukzVjN0F51P5n
yF/MwRJvADSYn93cOdFuUOC//l+SoGHeYpKAE4RETeCrRKwPWSE/54BWhz4qhBCTwnYXCeJzDly9
C05bKiUiy6wE5+NcvAP2cUDBlqwAX2vET+PjRdkMO3wxdRsFbBgb2UUkHrc8VBkxwnFOYno4Ppt8
1B6FGHRcPwJkVxodI5UqQkgvS63C0oNp8q9WTk2YJNswDfNXuoRPjXswIWY/RyIs8jzfpxWGmc1d
Gi+GqzMy3kSjgzlME3WBfWflSuTw+OAGqdhNfO4r6FvJLYUTeOuyRn7cNzEFIwNiHg8FpKVNNH4y
sMljxuc6e6wl0mwaThSmpsnaILBk1f0hg/PKrIjIJvWALzSTF3qe8KiQJzBLj1HQWd0aCVeDJt09
lBpKFBC22epct7iVVCgtJEm/kdg3m03t6+fRyTAvLNpDzcvefy8R+knSU311MVMuSmWKQ5LVfkf2
N7XBu9D4eprj5vQrsJtNQ4J9Gvl0Y1hKmDfYvB8rdtBO8tCrV3g/sPBRTUmAQk45U0KFosXUweyq
uY98JXIrSDUVHfEDjfvj25NUFwD0GDWfgtWDKipWZvPPgpdNAMCDZagAeihCJ7BHcIGhX29PdqWu
IGDB0A19d6aDhb5yr/vENNpVUOC+TOT83l8TyAh5M/B3KwcvNgWDENGRqoTpdzXCn+sVg192uCBz
08hwM7DQzPG0cqKcuhug4tIs0NDLXaO0oFAaebLnOfBFlWo6czVOCDH329is61mG6xwG1z+X4pv0
0MlC8XerhyHOMCE/5zzc99aWucXbhMEFzTpXdaMNRDQaCESIS3VD5CZlNN7owjWMFwJU9xTV/Z+h
+Mj1Ehe6t6+b34kNPt2iOd5eRRZUTHfe6Lz6x2OSG0vPqQlqhGIcR+uD7/yqYvZmhO2wZpHQ1/G1
IsOQPBqUH+uSVZetuA/DhhATQX2JDAvhswNAYlvThRpDL57qei87UsJxCyl0cRmMGFAKiSyMeUoU
ykPPPDaS04nr3l17gfATqHihX4Tf4sQqRw5iX8aJ6fWPsXaz9OSDS8hhWsNe4TvFOx0ZITWFSbq0
GNjZI89PXZpXsln+OYMFLRUHoI21hfch1hfbGv1JUC4rTeVsYgNAzYmRtruPupsa0gMtqIIDtNQJ
hd2vjls5TxEH61fn4iWUCszgYLSmvvn5oRWNHrPQ1+Sn4Z/GdPv9Y4GqNTCrxn5WztQaPcRpL4hL
NygOwLqQWZs07BQfxyfS187mtwT2++X4A6Ka97gDRkYIXAJwTDkm/EEHtcWDwCWE2XspkY8NablS
MqIlr2AB/wSx0xut4N5aIAjDzM6Mjmu7KPdf6avYjTGqF6dOfzUpFnJU9N1oxCxdCKdAvmm9KTEm
l31mk1lbf64z4+3sqckHHOwff4xq6AwIFG5yzpsm9/Ui+mfQab/C/+s8btf6N0TlU0n2A8DNxKc7
Zrj/HIhLYq/dvLVlu8OQE1z+bjqCO1142TQs8GoZJZbwUgfPcblSqg0F5CttdsdP30yf0vVVwyFg
cIqttLscIIlXx0BS/LeCr8L6NjRkEmvWx1OIo5eZHdAsZirlaokABcTveK8fzrOU4g/QfMx64A17
qDWKc49aOQFSCZIDDiIjbx/btu//hK+KTiLt124E9us5EFkAv9YdyQgPcewX9amMOdkm5zCfrFnN
0LJtRQyzR2Gpj83XFgPbfSDmeCX10dPkQgvd6l2CFme8KbzfyE2HJM6sxj3ATUG35pcKUywWE9zt
0wL4a7oLXH6Oz2J27ehkPCmSE8Cdj+bEHwmzUQtfhfE+yKogc7jNR/Qe5llWRJUArtoyQWRTocJY
4CpONbVIojrxGRyfr/btV4PR329roVJVu6GVxO9sgvaUn4OMO1+kboavtJS6aF8nIdNdNc8yz8ll
OBogBe6Pyzm9h93VTaXPMLvcCQZpdh06WW7N482aAe4i+3k09aRUpqs+LisJvIuXm8nrbveF2CSk
nwWFalzwToZX66eliZLXl8P6RK66rG+Tw3Ax/8tPgRCm02xkPIk7/+w1OXLBqizWuby6R0juqa2d
T5oONokjCBeMOEa2bMnvHG/5+qg0I3VYvVaikaQjdWLygXZTDRkjU+IlEBtZZfacqpZNxWu0Gv7C
Oo4EZ085Gea6unUH8pqrbIrQgFt3hRHkgPnkzmRNdMm+YZXj7UNczGKgIko/5B9vH6wzMr1Xr7Ra
8yAiDUHlH8ecsAGMKW5Umtc3wdQRgThG8plHnN2urqf7gjx5Xg/OzsbOB1c08eaTMFokM0F+3sxP
g0akr+EfjC5BNFf+5AK9nMQwg1RXPCzvoVEVhEvTbTmKojxHqhmwusn9dHxRDfamBbvLAZ9nkrzV
qgJWUEG2sTBxzAoPVhTEoGFpDgs9TJPBfEy8q+tGhffcCOuHqyaIHoR08Y3vd5QO46lsV4yR6MgV
71V+2ccGoahO8yfX2vBEyb2yPITeZfxAP7uPdmad9Y14YtZfSXj2ScCNeBov29RJvSa+heHW3Tlw
uVEMvE4zhGrqxK/oCWMXDD1PGbYOS4G8OIjR0V3zBwSlvWZmbwPTQlagDayoY7GAmF358Q3onfyb
REV1DKDOO0PLTKJvenKUsY+mDdLVZePhMkasjUG/2j9z44MaAUG2KhFMdQTXpLLQS87r0PWY+/qt
lsuBrkKgTH02+pLZgKMrtlOL8dpmLPpd6yEbiKlO1zzDXL0dOm7hC6E5RLRvN/1iGQgd6Wh0KJOQ
xXIJb2i/1jBY4u1GDHv4Yo8R/9WmEbN/wywiwdmHioCC5ZjiWZUZLBHCTXwLyT1oelw/njhZZNBw
coOWAQLQAv+Wxd4v8cbN7Mfj/OfY4aDWOKOmr9jue8iad6c5hO+QllS0Sr1l6zsD5sXsReszF6MD
e6t+mSfGNxV9Ke+Fw81e8ZU+TVMFn3x01NK2CbZg+S2GBzYSmcIYA2uOlgZZnmjNsd0m2S4XRCEB
GfCh2VyuQ/j6Eam+rv30+5XBzrOqtaZaCSnB3I4Vhc2Q+f2+9bXRFhEpEvf3HJyrSnl08WYtxLNS
4REEFxOaFIIbhxU1wDKg/p/gv+REclF316H5VcsHlIgxUFE5fEfOCJqifMvdXZCOLCa2tFFP0iKf
AJbl2Xqp/5T6pxPUM7ydf0WjvKD3X10oIgUvDAPIysKFZ9zxAAWDlui8ewei51OvhEaEyGCQttVZ
CllElfPItlHuTEoLAUkLXOheHaDaPuizcUj4tgVwrwxK04cTzf7f5uitMCWXfneVHYEKTDd83AKq
x0GVCUJRrp1WrsGIuVBI1qfr82hDcHn2UeVeNaDtXbGeGlw8FV6Z5OpgDN0ZSLWoLMSffqVYJmEx
23mChboeT7xWE2eZgdtfUmB8nK7JQIawzpy6mLWoU3Hlp7l7Zgt2yDUcbUhyWRgoqAPkWuHTLgV+
7Eip8uRE7kZwVVKJ2RR4DA75q5PXYg3cETGqe1zmBlVje2pRAiY5uBisM9GW2hI2zF3sXg4I71j9
MJwjGuKMeIywC0dmjHR3Ne5hTXXAE7rHUkuThyHWid7Io6HGOwJNNxrvwUPF2zgHiFN/Rc6IqaaC
ji089ZepP5B9DaWn+xBbPcJUrX+iMqAzTu1fbiQx7RfpVpCRUql6WWnSoX9K9OfzN2CgJQoHNxbA
woB1mjC/vHHD771Bx6sfmFuwnMVBCxdvhMynVxWEXr760lrG81FsdXVmxUp6iIp0YYnV8aY7X1AU
spjoNbgpkf9M4nkpBgGwtAyjCZduOZQtmsD6QTyvdUvlrPXBOAjDbYZHIsIlnvtEsPEXd6YUzmJr
igO2zBpHT1vwp+/bR5nOE2021wjXv12OpzscEHxdxOqYXMiZ/siAutP/P5r4CBXqoXFIyeqG8qV4
kMuSEMPHss5SvNzM15fCR5Jnh0GLAIN7QLXKFeb6mqWuTDtQcPc7nq1Qo+tw6vaWXRX4Bu4izCgW
jneGKMYhG4XskGFlTYJ03WntT8k1+2aHMV5LZ9eH6HLrbX7eBO1bZntUB2HlrcS/r+yf3oC6hyYG
XFvJAXHkYeN1ml1z7L5lArwstSEvbXvb5myIXaqezbZ5Qx/3kgMrGXt9X6u3PqFCuwkTTcAHnDFO
OyvZvBNWAJnOKArVQG4NocSmOUyHKMfGVPOsB9g2cjQOSKp0GkhPCAeh4BFIuWNqDoMcAss5b/WE
2p63ZRmZnWauDSan3SmnAINmgXXtTBJPTLSsi7emv6+XIdMgueFhy75rmDqf6lrBW8lcqu9mL2DE
ZWd18nkWoss6W2uk1BgnGrf7fYJtA2m/zvw5gtzBuqFkETjPkEdzMhByQ2FgFnK6p6TBex+eiEjS
nu0e+dbZhjsXgxHJ4GMQHXfziZdwDZ1tcKnLSKCKe85dLtvYIDItXdwz1Mfrhtd64Ows2Gy/TWM3
pwEnkS9WVMnxNWD35tpUGl1tRFUCq7uaR5y/f+cq4hah13xJeEE7R3z00xS1vYBt3g3ikIQhxzg6
r0YzijYGqM6hbiX5alX8vdxytLuQj8eUuP0IPDuaAYVCglJoAuV2UsuWoLJJrzugF7E1X59lU+sB
bdpHzE4d2G3GXTL2eI9cLUFGGMktH5Y7mX+9V5qIaoKJcNn7DeHqPqy/on9hKPqGLffztxacfADa
XLtbvJI0ejgNmi4nPcZCtBNc77LHI54kxH148808+nO/oy5yBF2o3DHg6Qyl/kvQlKzVpSQ4xtar
JpshqWDWYMTZBWU95rEf5fdDeo7q/gHIDXn4rFDQ6ccEE6fK6Ate9H2FPnIXrfoVDKO301TgjSIU
BF425aC7oWrBCnXa5WhyuAfkJihK28ANiqJg/JJS7If4SN6vwkfYMLjyt2hU0DbbPBVm3hROFDQN
obp947y9vzf0I7lTEcHh3SQUcycskpN5EoTVRVwTASJpQOiSS+3DD/joBjCS2xeT8C9tdktT/SuE
knT1GHUBTHGiRft1AQh/j1UEdGoKwk/ZbMPpXlLyk/qo/NLL0ylvTVUx3nSNwFNw2buFX7Pi2yPC
L7MsL2h0lafBRFlxKh6YTISWwPPcLHeLhsrpzYpZQtHpaz9qiLRfnRajrIHNP9/LDSAwqP8em/6t
8/6yzd6sw0AL9GCkMSiOaUGtE6dQblWCFbLfdMtsYsXCN80037WkqmW2F29NI2Ry5yJVHQLcZ+q1
WAf2SBxBz1aMIE+G25T7AvnYYt7OWtEVi0+8+R3QyOT48dE7r5rMB5p/9cDrjOP61WpoBz8ta19R
p9GJIrmYB6381zuFrZ3RUb9GLHzWx2mkCTdozGFo/0FnwNNs1OR+DAYyJBJzEYqQ8YXqu9TdYBUx
Sgk3IyQ+pTLlsVGGMMGP/L39zH2GRPcTbjlvObAzoHZJ707BMTLBAod0nyS9M+LOM7gkZw7Ws8rL
aOhQ+IlL25jzKa12uIAVscbllpzCUrodCHSICy+JePTxow2MORb9f3+X/cHsHoIkSqyt1bKSXg+Z
3vYYhP6VVUj1FUy3KoRiRA5Ju7dFqvFyI1AINgV8NrSSB6cSa2GLFz9wQQL662g5b50hT7dR9zF3
ElJLMdPaBofipRqlbKaCpIoeid8nXd/4SOjRUppOfylJaNjEWLr8DoqAu8DKDPyven+XFNYMDd58
2ocvRczgORaVejy3VmBDQEIE89CGDZ2v0DyNyO6jOtcBXmL86uMxk96dGEBFuhP3OpxyWUdUI/of
cjhtUErz+ScmHB+5dwNDyK9BEwcp+eTppcqxpdti0klgKxWUCCjRwq3Yhl+jdDza6RJfdvVsjOkh
glvFmaL8AjmRoaVfLyWx/k3DvPZQzqLS0or1S9f09uu4XkN4fREb1NOrLx6WO0VojQyYo8CYs5rg
iv1MYRiDL6lc0JiwdQiMrDjDW3OI58FyoGV6OKOfuSL2rEosePj/fkaB62cd4W+fYuEHQlnKT4Ex
Jx3yTYvVnwStFQWnrYnwDcD6G81MtemoQKiwjYsxHgkhCLr/y/bgQf/e6St6w5NXKxbOj9gCGgld
e6Tg7DH+3bKC9wOR0PfHzdiQpV3pjDeLRWHjecxIfilcaPxubniotIkTHMioF/92J/bW6nWllbKc
N9nP4bNx+NROB4lT+Hpcvl+nOr84DnLe1dumHtf6tRSLoIquwqVIWhgg+4BeAdNOzeOIKfZazYOS
NGVhFc82gGFMHDzM3lLpx8cn5gLkjJ13GabujTssj5ZwP41MG1VUSGkRxV5J2HBSNunH/42J7fWO
M4bTyvxcMyAk6dv5i5P5Uqhw06EtFYIidphcqwDXMxsXL042kNdlcbyAjVjf5l17hgEeSqRVcfiA
nnqhO1RfdttR96KgfcDY5yzjTDJ5OFUO1jRMKZ1PICJiau1DtvERnCbfVdGg6mkSwjUgFO98R75m
auopeAoVPlwwyYa35tJ+PLK6JDArpNx+17uIKE2DU6GerWpGKusb1iq4BcZoxDssWfrYURJWhf2h
pEf05Ufjku0qf8jVfuMs6Dar6DP5w8orIhdIKArcajCiai62JgN/CAoYaVMbx9iYOQ7KeVpmaZQo
VzCKdJWXB/yStMbseYebMJFCVLHgIDbYH3Gbgd+p90z9dfr1o7UsSv6DP0r13WBaCBH21XriMcCV
gS5TKxKz5EpYCgw9+mTG+Osd3bJ/lQeEkUEDbAMC+y2j6QIG/W+Vv205K5VMthO+ZUH5GuhpEPMH
TF6dss6Rq2ruyo0kg/dR5QJcH+o2DbeXgY7mNNm1aX7vNn6296b3igS4xyY0UrG6Antzxe6I9bcp
wMOrzGZ8MNMprdR+SnWm0WxlzbKlFPC/25O+1FF1rUM462yXGZsdWzXS+YkJsYfiWId6Nn57PMoa
1QwQW3TUdYSeMHEC0hbSunkqENFHHScz63APERXkG4xge2X854QV+mClZ2k5sMZS8M9F7ET/6n35
hzuKC1yCkGR9u2Z4N+Mro2PIABZni+pQEI9QO9lrEwfA/YzVU43BTLiGFD4OehIzylh1iBPIO5M/
kEGNOF8Z8YuDB91Znq7DTdBTv8snKKdqTPpmWrRNjYuyg2mKwUZHtgQUrVk175Nci9jmRYMthDhE
M5MDOJ1yomATSHcNyrlepg3bQQTJvtFx5whaGYuyOje4CSSRuRF8Kq8QTe9Heo/3etInVYM81nK/
AM1HJ724dTAShtMzAAgT32VDYp+5GLVKjgl1O86Dt0nk1ji4oY2nLBIlqkWYjzeVAb1ZcN2uLE+Q
YDdHGaXyK34dJqDEWBiSFVyl9cFpR88l8zRGh20ZtCr+SUln/xdMt3XdUe9vB+87MEo/VFr4jyVm
a7Uo18lIYhaOg8wmrY+4cBoCo24KD0QPvqLYVV1rWGEjC1g1wQTJ9803Tzz3RZ6NEnu8YsXE2+5C
dh86jDg33xh1Cd0JhS2oACKXhJ/lco9kjk4OwsvHvRFacYjKLxG4oKNGIhkwDxB1i6vc9O8weXJq
Nx/UvQskOs5wrkwHa+FX/w5+N/t2G0YPeoBiqkitsayP4aK3sFSoNjuNLxxXGzUwesFwp4BpI4yi
Y6h4sRbSFejhuoGu5VOVQXTogpCTZUSq62qaF4EyCd9kOGa4grFcIcjEIn0lAiLtmksunLL4M9Dx
AZClbuCtcqJIjuCNVnuIXMj/IB9IV5yN3Z2hIAcGRvr9OkF3QXfR9lteILslRPmD1f+jgu3u6cFB
K4/QmyNcDt3uAF+OpqA1b+oWikR4jLPm9Wm1A2khnzMB58n4433RdI6JR5p7u9FJ9s4FQPoZetKn
BZ9Oc8OimPjEgZSAA8+Uraj4lL5AZiiYc8PEAm81VenJU314FjUf6EicfSFSgg6PmuWy3qvo4Gjb
hynLSp6n9TA/eC/jghustPPk7pVuV/nZw15Oamz/SovMBippI0LrArQeO2htuaQ4oq1nqn9Dl/zE
wrwMIwLAkRAanK7MEuTUZ2kEhU7O5kCTAYiGLIGbUo+8iCVV3jakUHHtRXyeSZBjTQf1hP4imxU6
BE9rqOhiOs3RMCUaIU217RdiQ6JR9unjStELOHjL+n6xLAozjvZqdEXEWteFp6gn7OXjJPjLGIJK
YQOcW57EnFIB1PhtXrTyy3v5Mzkz8TWdAEF3JZ1ebJStJeqcF1Rqizpcbg0O3qre5oh7sI05SeY3
RheQqrKUExqeGJQKrIpJEfNMtSue+kwZ/tztRVgwuloJZUqD4FyBs84ZatUl3J4IhybzNWs6ZakK
BKmNrnT65+qi5ioOXGRNy05BoxPY9sqAwkIF5CEQ1gDgBc/Qau1h0UiAxeQoOczhTV3VZF74Rxw5
xTk9fekoh0bd+quEtVoSthwQBLAxDyIIYSR/q7RGnjFXoNSjQSrgpsjdKJ/Mx5erPjFbAu9let5y
2avqKwciSswWgUhCbnXZ0Y0fTOeKbnPN7SvHuRSQpMTp4joOSGRF/BmGk/WZmoydnkKs7UvoGW+9
+6PcWwrWxt2xIezZennP24A5VGC8suI+Z7/bi4bccw3s+Xg5n/Aux4Rm8egQKqL84ciQo9jjYT9f
fb6Ki/UtRcTCBoyfpGZf3qXpVfFK32LSvD5MowOyNoCR1ga3rnM/0zZwjUg/zddYYxwAFNo8mk4H
zqcTgMcQNfGB1BnqCk+odR7E2XnvwDAKhxZbyBiKneIWSguerrn7mrOTQQOxxX0ZRNFhraVGMZWr
HHWylJRSBkSbUtbkG/mqWR6XbKzD4cvOH82Xquug0IXXwPTvA0UNgsNpeh1s1tk2OxS/8yG7Rd/J
63WXeeTZQElXrbphAwcWxasx3strvBYGV81bnGGR5PAytm7A8EQKrTLu26ryUVnoi8mewGOYN/Mz
7IWs2OSD+I/Xi/rrfzt3Bb/RUyEdggHOV0Mf2n1pZ6HysFa/CRT5QaBmRhq36fLr1oBe7UrMVFVW
DsJA0hjJ4eFRSWGn1QIT2F06c1dy7O6viRIs/R+G5cGPwMrl5dLArr1K8eoUTtMw0m47xL5xGHxc
+t8F5zKnYtn1eeypacksM61AN5dWOuFdzs4VO8irvDK0KOcsk7w+lozobgvuAkrmi0+BdCNMXXkQ
dPzCo7r40FHkPYtIB6k15jqAD/yQ5k2WdgmDzxcV200rzDwCwMVzWakVRuAhxeOPN5/SPt7pZQfj
VTu6V3SVxtgA2AQRPnubKvwhVgCfE5pgltA5h7IG1M82ZzdOjUxizgQNiJ2/CrT/9c3eTQrQ64B2
E0jOzwYNdMwe1EnF38HfCSmDstXauipIU061xQsX2tO+l1712ChVYxnw22OA/StXhyj6i9BpBmmA
k5kQe0eezQm2kbxh72TuHq+vbef+2eLksplmtxY0Wn4J5eJ8cPfv+4tMXCbCGdzy5aVWioEN1VaD
wkoSd2jc7CmBLC8Pi+6oBjTzin6mctIBd2DDy8eEx6tCIWKTm3k/7VaDZefcjfprCfoc3J79CxFG
t9LAKBxYQiHSKfEYhHQvLdxGwcEBFHq2Ibd8ueXGFNxouSzDWYwMWj9O4EEvLtiIFJiLDZMrySxc
HwsxSObLi9PMRKAd8wSMI/DVmYhq5DCEJHjadlxqb3rhFrhWqq75d8tThGv1vKb5gMtCB/GBHeqw
cViOIx0UbENEuQcOEYDHbsR97zj4be7MXmDNxKAFGTlOtbC3ASbZdluY3zMmfMar3Cviv0W0xW5y
KLkAnMoBLWcZJFCNfyJH6SvafICmoooHfdr4TBe9UawjfRYxDd3c9PapwJP6ENRtqY6qQLJX+2SO
kH4EdA5NJ8ZQ5+JtsWeYGDgo5gGgP4wkwTdru4mM3SNqRs+uyLSAzeg8n1aMQj4eXdAGvaOd07Hk
JQYUrC1Px5RG4TfsYamvVBi4p6LM1uZyHd6nTNZuul1nWEzZnVNU8Cm80aXG5SWWyCI7nKiSPUSC
b0lok5jP7dTMTBrs6keFD2Nf86duDX8AOmbhOXl+AOl82hOE+sDGPVkAwpFqGcRufnVFj4KaYc7X
9PEqL37JrlWPpzAo6mu4joLvSMVMWBLJTDfsBOGKeKlN1exLuLmKzv1BS6Yf8qrw4TtPfOXtTfeU
qaGDSZ9XtCtu4zD2HGsVGUwoQ5vQrN7xbXJ1dEm1oO7rfbn3+4zqCWlOsC3q1hEaMTtSGYTdlLI+
ds2htm1lgundiwYIjX2O6Q/wxNgTFL9lYIDzQ6YTx0mGXB3zO0mVJ+3MTpr57LNs+ETlb3QjiH6v
nFMI/XpQFEn6B+qXascGUMd75/OfzOaLU4ogCQgGJnoxzxoENdvW3hNRJ1cYwPaMzSyQ/vDeyykT
Q3MTqoJJDzpJCypCtWKBQ5liRx5zm+DyhcEubpiAkWeoRaFLxmHs/xWh0cb0eqbIcQOeWUgcOPK/
tDXHfL0Xc8gXd2x8lCeifdyXfhW5bqJl9ypcjmk2+J1eiWy3Xvjo30WbQmw3i0fzTBQ9weYXK6/K
/RRgQzXW/fBwvkCmzujPHiJZVCZvd8Du0B9bGh3epaaADpISolAXINfGamPshtxcZYenAXqqCfM9
OyHyhKDkdUG5Uu4aq1Yp+aMMcguUb6UhGh/iR1GR9Osaid4gigxfa6zvCMGkpiuysVCB6jTz113s
uod37UFsALcEOvqx8SPahmxsFQR6WbRVWV4k65bkv3nFkume815Y+HqsOLAA2jNjQsrTfouDwx3q
By6euZ5D62a49k4EWOmfq64FEJ7bW5cRbUbUCF1MLsyQOhvmEbKYPoC9SyVqvkqcr5I62tpK+SAb
BF18chSTYXeCr2Z05Aw6hEXDzSz8bqBnxWGmutY64kYFg7u4aTfPXYRwGDny1jhf9vwnvcQ9bnKM
tdfKNduIKJfv3bRKsM4fJVGzExXkiITXOs2YwD1YyNaM5w5rgtPZga/SEq6IkSg3O8aEFbNHvdU2
AcKG3MuplZcIoaGKIVJx8DRgmRt2+am5yl6ibmdEjFcYSix5LltGklj07c0ajRnnOZTMdKJtHOTx
VSQjeRJEpvt8Ie9pXrYax3GPn4i9BiE1wFvrdwoKDKL2n3QTl+w9J2pyMgq7Z2gyYYJesnEP6gv4
fkISrctQK5+zBx0U2xak1r8xTIhWd9j92ri08PpDUUUq1FTivsYcTjgJ0g0AFNjhgGPhsBVwHG+d
aRO1JlaqBJhRqBOUVr5rPYvL+81TA8AWomEI5OSjmRAAIMxCHC5giUdLx8ErcSWilY95JbrovOt8
ORsTi7PSweFRi4GbdhZ48KpqhOKquIrXHR0mZmdhT51L/FvtQEaq1f7I+helRlVjSOGJUJOiuDcB
7B4mDYxXFQ0WHvyE29nxYB+LhBiEwSuCddN5OpeHxrEsjzqVl/toqUSSPYk4zrRx10jmQGTlNibD
WhLlbCxcfdtmTHtVB8qkSGKaAm00HxjR6vvgVfUakqm3OWoL09CehHWfvBzZWZlXP49XpQmXl9X2
rceGNkT4Qp0fWH+fUGDJXAiMVSEh8NRmMciSl4l6Fkne8rIXCIqbFE0jfovoQvk6TUIYytE4Vevm
ENt5wC/ZAuQo4xlpSUPtWPW/jzbgb+waeMSv4vRSzfKNHquQsBxh805I9SQNCYgiO6WkFYizd+X4
EhbQX0OpzDl/ltMKyaDfL2q2mGCveI1OSxmpxl1JcLOLTMGOKLj8hBn3aA2ZzFwd2D2+iAPwODht
8ieQ+X0e5jQpj8LkXoOivnhfqFTS15fd6kfWJ0hKv+1EEra96aDCsi5ACz7UFQ5P20wUyy7TlUCh
rCtMf0zznudih4Kc5cG5FMZwEnCjTffH2cxdCMPjjAW/ze40+JhPnrP1YR9fn9GflEpTkr8JglT4
KGQmASGKxF/fpMDE0102ka4jzrhWk/Zopl0sekw64Of4chL7MbebJtG51aAfToiCRs0v/KCo0BVv
CTln18ZVlhzLnnrIrc0Zupiw7Z2mBXTtuOSppfijDU7R4D5UCFsPTd9B535+WZgFkLUrYPnCfo6+
vos5nLySFnEzhSXByDlu0HnG5rAC1h63QU8ginIN2DVZ6vek8JhVEUxUW3PPUgrx/jWT9byM4OhV
uxcm/6RLGodEOK236bo/ZNpBHeLKrGivXaxPWZdogecE3z1ZnfTfQJXPCQIrmcDqXN7RPNEjLvm8
5Wr05fd2kdHK/ELi55o58RypFEcoSx0j9HCqJ9NA4K+z4unQSImideynAYsTN1P8hPU7NeOP/YSW
EE/BL9QalgaYRWA7u8OKc/IFRRVRw3c43dVBl+RbK47Ill72JX+Dhs4/33GseWnS0RRQFAvJOB24
hFDxlOy1g7Ym0OsruFByVwrbsqnIKyEwPstKgtqvRNu/NNskd2EhcrYauOL+LsddeEzaAzgH9mke
JKK8wTcAh+ZAUNh815dNn2HrpcOjQVTxD+qsBQqNgYPQrqVl7AC9/DbgPAuc/oO2czeowgO7p/Ug
icpbNfExqqz6bwcT9bitZjBjga0aNlh2oQrYEpM2uTPk0bkl9GLfjpvhmYoCSSWRBepjETgBtWfx
GwEIsmJelCEDX9UsAjYWBHi2rrJM4cUMHMqZZ+UIw9L05mYtDdJ345ZSv1bP57/Ouof+YlnRoXhX
RH7943ECD+3iFrXXE9SgJ26ZLfE4zu6nn7TjNe7DbmNFJ6ph6Osh9AVxaR4ywIAOMa4QzLfu8zfa
b5C2iTyn/3f7LNG0R7aOLe6evbFIRvFQwOpzhPQzvDxCF1TgT1lt13EkdymR0wPhyLI7FbFL1gkc
6BtojBvw7GV0jU2gkL+wCidFsgt+td/WRGo12EALZkbCRTVLGgdcwV2d81HEjjHPeL6PBN1GWDIY
Ht8Pe/i/XMvDDglxjisLq8LEvHnDkNV1/hk4Jvnviaym4eQAfvAOlWg5epEHSwGO1nKlUhdtdcoN
HDll72qiFltSTrV1fMkwTdNjYXy+ulZbc7r3pV6uZWOTP5JdPntwdn/kyEke6zwVxjhUfgJjUosb
WhlBtLKKipsVAqAczl8THPMXJ09rD2oDZ9kCNgrtu0bm+YH8qe9VufgObOjtLbuSsw543soO4A2q
1R6e+DU2WYOStbsEPPty1iWNhfTQ0qZ6udn43lwUPlnp9pIs3+WdrVkc19SwJHtYKGKi/soXH9Am
+YBoyGUjr3oF40UDfatgmeh7kU1NfZ565f9h2ShD/FT/6kGiJ6k84ScKaf/dAHbzDJ4XmQLZR5LZ
7ZFUUYVoI82yZiTWxZUsQfDfIDvgSgDn2bPszIL+bUZ3ha0BDaHzX25mqV0L/ly4iAIVZF38T1Dx
iRivl6vrn83Fvf0K3j35CVhCJ1xJrPYFZQ5ZMgDUn0WzZb+Snph3ujGkMYi6/O4zKYSJzZG7eFU2
ExiwZtgRjCYgC/flZqMqdWiOxXvt1iZzdaNO9a2tFR21Z8r+khZcekatYK0bk2YKKER5MwbBFO6X
xhzVydyjlSJ6bhH87iRkJfJ/cYZdIePZcS+5LbCc2bi5zDHxM0iHjN92lysBUBTTgXJUZDbuexaR
FRpbqJQxknKc1BJnLAH7pCqv9GDPf7V5ElQawuM+Sz9zGrQf5WP5az+KFD4AhusQ6ebZKb1cYMwP
za9jS0R6dTci0IbzyrzxYJHi+OcsBly72lLfpg/uADeWu3JzC3zU2QscF61laHQg/2nrCiILkrgT
DwHlS/UQpS5GmC9EchJwxcTwWVucEB14XID/SRw6MqMDEny2bPPFAoTk5VR6j8cvRQOpAOs0X+jI
9i+3G6+XK7HyCXj6V+jwWaO3Vuv2xhQoxQaVJ+55K9QY31IV+Q28fhLG4Wi6A+aIWfri/baRrL9J
wk+6sA/QLaXGDK+jiOvYcnLXBYYnHZai+gtkhN5KVRQww1YgB4zLmoyvWebgR+e0+QcWrUkjN0TI
jsU+/B0UNqdmyn+nPXiTUx/rfZsTicr4rhGPibz4UYUaHKIEKVFmlEx1Va8r7y7hi53L2ZHYtogO
crDbIX2bxpGkOqMI77hL9clPtVrtaSItxfecvZRIsNAajMyR3w6cl+jRwdRr78MgcUwTBPjcEwbn
f2+NlfRcEffWQqlHlI6Stk5PRDCZd+VL4jDX+N9CNK1Rs383nmx/bpBUa0USpeBa5pDEZNNdSa8A
lCKnfG5hLYGtRGf1MI/unVHyuKRTM7DfCESn2SV3Gdux+/jbWr0eWEMgynHMwoHzJ5fzspjBf56G
FMMs0bCiZSiS3REBvLKpl7dpmUhhNxRd8F2D0kfRWqnPov565WQwgN0Ae1r8xGm8ksZaoRRFIqLl
eTXeVSNiPrnMEjs4pLyh92dujXwzwRnZo+Ja/bx1U1HQDCs7dp5m//ElU/uoWtNpVqf3J/keyo8X
aIGXHAZD3+Aemc48Vq9HbF9QEdgQUgKl+xAdEPMnQFHY/ULfCEetjFGPrjRtrtt8Rv0IWr5AoOEb
K97MzCvVFMnwEXLcXI6cxoi+X9tERHs2smiRRqQLsxuCiw9PuDLa6lK4sO4sTZO9wqjs5De/r/Nx
IJbZBxoUWf0m0kmq/7pSb6TT+uVrqf10V4qTaij2J04WYiyL0DKRCdELDOnf5iDFb1J5RGLcpiuf
FR2vFRihmL7xrTA/zkcN6tvGxkv8H9NvhOuyDsIjcYp0GoBYZ2RNPXyeuypN+ov9mgWWGYC1A67t
CtFEwXOxnKesMiGyK67Ik3nDN3OyedT3+/ppy+Pv8w6n54jcEYf1PcrEXIsB1JukqOY56+hcPlD6
cbA7vfLX+YwMvV5Ktfg52xQOc+IBtw/MIxv5fnBctm4R2CNUdLW+1UGVnt3ukiAptFDpdcUGWemZ
6ADqu9ioR0FGeHcjn4YzDYQ8Rz687gKfNR8a/D6b8AACXWwQamI/ghTmXCkHAzpFLBySJWEl7WMs
lz9YU8frec2GHVvd60TLzeJjU0QHU55LiVVg0AMggkhUWr4gIsN+8YCeLEPfAjBDR9FIk/KwsFph
bUU6k7cGwctoGkC59KlY208lvFRIiVcGRg/CkKLjKMFR69MquQnMzO4/jO43S13qvlHuPm5n3ER8
cmeiaVoLT8cO/wgXsvnTySe4hueNRNMrM2e9qoytOJoKBB09ksJ0kcqUur6nA1dALVhOtd+Z8PLm
NHs5Yf/mhn04dG1exHyZBvoxSh03QW2420gY7eIedzjY+4/KaPoxL15DcYdpfxIWzY15sz7Rl9C8
MFMo7oN1SNhckJummtVMz1tLgk+PpEsyS0jqxFdYZkOJJPJc0mHn8lS2o5DNHxcEglb1sCRzFuql
2GSRjPYQ/WKVwiLKN5+AxNkyknLHOpUSkZcpEATjOuSg7yuRczJmTPInvaEbICbxO+KMFMlvNfIx
owmtDvjZCpv87sLhd+wT5aotmvR/9Netimqn4pS8L9wMeT4snqdz23iEdAS3qGObvYfSTOWYjadm
PNETbFJ7KYJ16wT4bOdBQJ+jRsTWfMHm18bjjLgX9r/Op1YAez5tKUnyQwWMhUkUNbrPvzz/LXyh
8Ja0WA61vXlCKt+44IynZA6g5FE8+apICJDQM6umX1jYjQsTiW7YSoRT9wV5+b+NLQmTfWKG0Q/4
D/v1Jvbgsf9SRyOYZtFrMYopqhBx+ipa42F7z9dZ2w1ji0yd/HTENSBHneC7eXHVF65/wFdFGEwF
Eoje3M0S9Gemy2a/FVL+eKaS2PALUD1iuMjX+IRRWe9PQ357X3mjJDVsqNY7BRnrcDqpskSIV/OM
qd80rr64gwf6Y5iSuamrB51yB7o7PdWxNGp8evDz5InQPpGaNa3md3yNHT51zMTBCSY3RyWgmlmv
YLezPGOtr5hwwQy+i/ywAdh+flGymQhTVJFBz2o9UyLMRP1R3suzo6AOdsRjLbrUO72x+pBanOMr
owhEe9kUDJuVwmnkZOZhnEdzyleI+0IC6x0X6/tWtVG5ICYxAK0AzEFLN2cmj+ut+ZjZLrnZrIfe
96A6NILFyqNAveqeFaAaiy9NecTQYkR7gLKTJg5SAG6j5CBRlcA9Djk/7m/5qwPF2GyoWbaWMWei
JhN1fvIWIOoj0MM071cPO6J5a7al5+pkBKzrk5sWp80cTuZYe9rWoGn6IWIcq8N8ar1tHcjGtorX
/akqgpfZPo+4xuMNZrJsBFRX2ZaTdzkmJdHo5QLi1/MpVgTLJE/SikVrRc87Ra+yNmFjCob54Ii2
7nj1f7j+P9O9yilMFfkkr4gds2GnqdUl+g+lgOXQbySZ+uH/jTatG3Kprc0+IZb3Xxjzg/FlF0F5
QhT5x/GH4lJPBRoruv6XstXdt2rnZWfHwt3o9+ifuIVBfK0Skju8aaZq5fsJz9DqYppjvf4GCB4r
rlGE6mvU/ahr4rKmuH3QY/ZKG0SYE3AW9CBrBD7/tmYOJjK30Gq0cXa/LWwtSy3p7d/+XTyD1MKH
zFY5jkdpUUh0Pxf2ucacKWvcJYI43RHckAfMo7FjfN2TN8vsvzFEvxrc0v6PssRcYUgFlX9cP+Q0
ezq0sq+BWqqsGstq3eKwfmzJ5Un+a+8HoGm+gL3vZoDC8ECiwo6/Bnuu9Hrn1lWTA9wDFzVJKU+/
bOrpQZkFhDbCDWTQwqODcEhP42OApJTxuz1eqBIpxDKumWGxiBb2RIv55arDNRnUIe5ogLzFGWDy
52VUX4Dw8neN3Cr/KIPudYGUfDEbmeAWzKm+zzYY85zlr8TxC++o6yQUfxDhsaV5jAapE7oOffgN
azYo9IQv7TtPvyjmf0cT5DAfsLT1bja4rKCYKa0u2v3VjrM5hKigzkNsA4kyOsJ0K/SaJdx0QW7R
fhg+GFFcqZIOZ6sYfQbX4iH/RaunRns1vGoiLb/ywC9GYkInrQpz22HanbYa+B2gwZAEyzPGmLxY
qKMv+KJ3TriT/PwhLzzP4N+HE9n5ryXwlrVsV9e6itwoylGnHFceRYx0LCBMvWQQZng6FhwEUAFa
Dd9+VvPa811UF4o+i5p+245QStI5gV20JN4PstlaP9eZHQkIZuvK1h+vktMMgm4WJNR4HIkExO8H
Ob9Dp+IdyUiWAJdE3Exv+zcz7YML3BcL31aQ4IpxHOIlPSBXaSskKxW+lHcXVwfwsc3P7UP5K0Cc
oEW1RcJ9cYvkfR0utwHR1Vfn9QRIqtuMybxOXWEVleb1Y5Tgdh0iIIBOZ7I1LEgau0fhvOj/MN07
PQFVYnHf+Pp7CkbveHRq2WsFD+eyun5CZqjWD1NEYejIzmYV08K32VaNZikqMlYFP0S08gqDHiXn
JJXeTvcy+LFn1vXSEuyvWSaFzV6DcgWksVi5l16Qh7F0G1eGPtxjuDQ2RqkyNZIFL4ljXjxmRLsC
5mpDrEAFc+MO5fDCUoTAxoEuofLFINEvoiJufNm0J08I68fu94GIr2qkBNwPLqQ3xz5tJItfqS9v
TUhfvZvmS2/fOJUbzubZZ33BpKOUrHzUsVMvP2IiQN2sSS63pFRIz3tNe1q3ja6bnDMsj/QrtFpk
X9HeBPWgAZvs1xFf9Zo2wHfn3kEMqifxBZnMky84CJ1QDKyUfHZhNQchUiuLnnQ6yPKErwYlvRMt
sHadm5I2BGMGlCdDoiOWys/DsZKDpLV0bpBby6/niisM1HPz0r/RrxxA1M40wnRXQBEyhaxOkBuS
US8VEVvCB6UNnc95OUT3LREQaJX7SvKMNkFDvWSscgtfBZbieccIbn563rpvKP2BwurfE6vTz4wJ
hi4NTs12wmVDlbIwsZPHhHRQ67KyZ6SkMB4E5ARlYX245QZMfz2dxsBnnEnqxQ0YVDm4Bah+DhD5
TprUiCR6baadEYMRCdp0sejMgQSBxfzQABUpndXJMC9D8zK9bVcCcKEKWAijVPBS74BuKLuWgWZN
A/p7ygYYWAuRsnM+9CyyuOZo1zhFMp68Ye9coVPoHPLjyJQl9go+8NLUHwxYxr3iJlwrLhzjU06N
FeuJZ836Z1Yr91pu3PWeFzIVuNTxsGjmnFsiBqB6SHJe8PIV+3iuKjV/gfUv2R6gPn80goP11D4N
3nc/10FJ2ApKfLhm6medeUV57AZUdzZJOyQPGJA6MXjzJkBSfyO0OYzQuYv0AoPNyDMXZmI3swz5
Z8FfZkN01xibptbgmB5cfuyloe9xzrsV+ebySUoSgt6cneeNsr2z8hymHzbCwuPHRYiUlJ4Sc+mx
ONAeM88m63NE/WF79XhRpORFRjTUxSF+qmvdvM4IpktQ5NZfSCp5ZSZCl9D9qrascqWgBfCxhbkU
Vwn8ThZIdyEQnInOG60GUPTods3C4h9xAy+3z6T/8jNWfEQJTAGGTIpPNY0GeUL+NjMUMtf7vowd
OCHIiR1Y1Vx3HdJ1dJEZSp0ncg0F0x3xKMtNu0HdZh8z30ltLXFIcK2SkGVnPplCHOQQWfAihC4V
NWO1RpfpDwQzRNpazB+xqUjyFhPPcP7jLBdZYDxRVNxkzwiTAZSMlgCQD4u49ag9WVDkTcCVpT1E
ZEdZ4MkWbsRluUY9h6qlfCr81O5wvajmGvI1xf/b4zvd7FWi+k2294xnddOFrd7W4joi7zQ5Fbd5
RIybXuu53Dcim0J5wOZN5DCSoTedew9T7is8PvxQQvLNnW1ykqCZ+/cwMXraFb31uMFICY0qJAVx
RLn3po0RjMmy8IWwmn8mQDECrtMWZHKYAirfK+pUAcTL5aIutnsz65DdgmWnq3dNdNYjUiRBxqYH
iYqPydIOmB4n9WKdw97vkxd5Wil4cJQt0K8y0naqkEsfCsiyFE/g1f+30Z9MPzFsnbNPatbkBQFr
JbZI3az4J+kYiI2fIxfoLP2YjikYEVIlfGbLOcEzKGksrpj0M2SXEd7gP52z4/CbnIbEyuwJkx6n
3na9H+qTS0IYhgp/AdCdyKRVEdWZZMM78dJiW83ArRezV7mbpmIDfelBLZt/xY/T4gxWTDmoW93+
fn+lRIRHb+sZousMbA9yFdSnW/B5QMOG/Pe4rQXoofx/a8DBpDMoE/VN3uy52pfLLEAYieUgKTU+
8l4SwNWrJ6XVDi8asNYrWMP3s9P2i4uDu1r8wSHuM32pP4CHjyhOIKX3Y/+bDfwdzIi8RdOwDxTp
5kSxjW7LsEYMuL0dM3Iaep0VtP+btnyPLQKiJIN35LthM3FSeQXo4wBca94QKS+LD641JV+aXIT+
T41fLb5setFshBMflafgIRg0kJAOelGkFD55LfamojYQEGGzmlKfrsSQf89V+brpcHdJWm3TaDr0
L0AVufT42y2WRUfhHg7xoHYgLmeLurpcepMGAnJhcUQ/mzx8uqt6UNpUghtYwVO4I57eLGQErbs8
Nih42k1ktWjL+9LyxQ64SV5vIrWtNMdpbnXaR4YTWnzvgCoi81nkGpVvxtWSzN0/6fG3MzSHC1sx
bSKP9poQqQaHBTXAeAFv2/aW+62FkvfzBau5uAqFS8HIhhBdfSweHGpjWx8f3VZTCkH83wEmSWlf
uaRNtZaI31B0DoI2gSxDf1mVfoAP7ptxNZLmTp3Iq9zE34PGQncdrC2TWh2Zi2QBJ79nj99MtwJJ
KBG3pz5kBDriucNvHVeHAYJwK9PC6ljr8NBI2RHTunnGG6ccK3fconO1F94Ygxla/iGsmF+oaM2j
RZqh9D2WWwQ6GZ5hC8NVVebP2mH3+gIsxltZ5LnyMUFObDa24W4SjJuT0mrdoYsqhlTpuqWTGTPr
3VBhn5rTYgHiIB50EFmcqBqh7go1NryUlNZjw4tR6FFtscU5rIZRSbaqb0W6WTSxBRZSHAvfAD1X
2ZhWFajhus7sW9xzpGWf8hyn4Hogy6VTEV7NlAEB+IFp/0AGPQX2shkw/kqSc/zaPGkvW86LCUKu
Rsbl3VEY7bhY/J6lqyAaucKYphOtjmICUmFYzxn6ft+lSAR2WNnq1bU+z/Zy+DKulh14r25Ae1b3
IeMZEdG1tky37hV4a7rUXa7hGDCqz9pIwlaYdujQmKn9mMNZUDGbvKIqCvziLX0Yr8sWe9gYjFOC
wtYaxOrcXP9VM7ZoWz3XbkVYzvbftdAvc87GaKRUCOb9l6lbRM/i0vATZK6HCvnr9yGsxXtY8KEr
LUmIVtZWv8wdQTCvfJLfgSPn1rlnCHgAJdhk5AJepxa3Ol0nhbT0HYn7FoWMM7KKIRZf3yqnh9hv
1JQafV4jSip67PQr0w7ovDk1ldsxCBqP29gHQeVEyhiM7JihxdrKhrAhvObWgyOwLjuoksu2Hc1O
p/3XeuvTVXw77btLyLX11JCaWhI6HfHbrxTfwPD38b/TH346uYG6t84FEi+hTJBKRsML6Re/vTbY
qIif7QPhg2ssqS7vAtXHtdLI96lNIJnhwptWVdvtcChLG/rJGFQfs39Yx+PM09+eLmnTkGUgKTjQ
UsF7Qi0ZWP2cMmP+DQEbcrDQ8+2UaTHUuu0/CJzpVhs5vK59DMBwJve277z9R0aW/vyKNv4GweTW
vLkDuBfbus57iGbj4s+5bQUMgKwfAP5qkbhjg/FBSTZOBoWMBf3sRsdvMezg8ZNKiG0eLbRlgwcp
qrZTkmCo8T2CiLY2U7yf3sEVnYvWR2beQnqpKx6/ZQledqbMgmsFsGBcOwPj+7z1Qok7K9IxSa5k
Vn8/HSku31e7UE4O3N1ScawUMVrY0xYapK9PS9rSoCJO5k/t3/fklM7OwfuDIqWBu/4F/wbYijQv
qLhmigMlRfdO5dUgJd5RQDAYb6L1nsh+mTtU5iQj706wdqLjCJ9g8p3V0ecIYWkLD2ZFj6kEUaf3
YMPIW3ck+eNBhSEe2GVjJ/4upliw+y5r/Y1OZ7mpflPFnNh8IYC/1nXYCY9Sa5t1zA/Hsfd62y2N
9QmellXa/eMbeneJBdq6rwJFloKxEqsccC+icjdib05b2gVW/z1yWHaiwvXqQOECr6FI3rPmjK94
FOt5Ee7YlIwbxjqdAyVqcZrtU6ferSdyZvUZL6j0C/DCXKYhJOa/Lz1RPUgVveWavlrVN4wMgJGA
cgTTTNxqqsIaiQwNLatCiwi7B0CJGtN9xqNfIW2vV5gvsiJ4JuFZ6DrxlN9X6d58TUFC39dSWLGm
WEF3/+EZKBSHIdJ0Vj5AKUPZr5ywcdQUhoruCNTcL9q6eb48AxzS+Trylf977m+hOj5g4TMJqqHE
ZGGMQfcGdJ5PlrqY8SGEYmZfDSUG80UX1vZ6hGJQhbbzytHnH/nmRUMIFZPiF7DxcJB87YLPUhnK
rH45x93QUq/UaQaRmnDzg57xvx7LtPYo840B/9DC6rUjxlHuTg94qnlMUMhW6WC/wvK7+snDE5E5
FOTDDkml/RDFFeTxxNc0WXONpBHkdzGJR4STknIoaTTlTDBYVZ1InS/RcEu2Fd7PSyBNEv+WUT1O
Z8wOw0aw0vAEFGPAslykqeiYdd2yQEOZWUX8XqDcK7dG8PnayGsMea8sVY5KGgeUPG/2V5vQW6lT
EiWyhEO/O8uP2UIxYDkl9cdkiRZj63Fotc88r2eoLOp62XrRz6BM+ybHlZKdp0hyEPQB2f+uczGP
/SSQyxO+zKk+yp0wtYWLk/P0YwyG6Ui/BKXErF56ZM4PEuJ+QSKEvnf8zwTS1XwVL+CDozLzWtpm
UaPpQTdG/nukP7VuWnLSUUWsqEkOsLv8v8SSxBIrWIBEdE3ZGo5E4jA+Sj9uHEOaAx6e1M/PuOna
L+HmmLb9GMCM0SsYriebFm+kvyAuMlsSe5jpPsoyLfjHNS6X6Hq0ucT8UqU9SSb7nM9svexRxSHt
R91KuJARy/p8+80bER9ha6tNo6GGSID+xpDls/lG8isni3vo9GIHMt55ewSbM/gVomSKqhzYko7W
dA92dKoAm65MuyRU6Wa6fJZR4GRvSBJZHz7trs+ReWQxeaMCDP62SuJfJPzQGYhmCqSGxTqZxEQT
yqzg4V/NxQM5MXNFmWSHV/Y/ub5AKmZG1zngi4KDa80Jfsuv1MgdW9aiSjBkNkYd7YBtocVqpl6o
sKCkbmWmZcLpS46qZhpXMfbEyQBzyRh5cZDU+7dRSp7dmcl0SK+htpYxS4H4etCVZjvnQZgCQsCv
teSu7Jb8khmBKAMVu4lWJKw5bkxOu3Y5kk4uXeW2PKIplTywlfqugsZoIUEdrbY4pbZty5z5kqv/
7sVer2a6Y75m0hw/8ji7AphSOOaTA38dRhj/dZJZKX/snX6DlwvvowOEx+ttG6jQf4aS99YKvPwC
pfLSlYYJgxdHCyR6Q/KZkOEebIYXLogqslji1kxtqlMI06+zvlFEIAxyPRoT3QPMKCrjWf7ogw/n
6sCxTyhwXCCAmDQ9hSqPRC/9hcKkq9KVEtGiFYp2X6hJnvYiHNqYyzdGsl0+p+aroH1og6Xa1vsB
LtrLsuVyDd1kwWiRHUb1rjtY959r3wuwTXkuF7hMVXsiCuCP85dV4SyuhlXcwgGigbJVGLDFtBIZ
qRCFO4LOieZIsNCn+RWHQAn20rQLvDbju65Q8zXAMpU3RHvh4rVNAk51uG/7esmdDZh8PA6O81nM
jZCdVMVauvFYTFobQ6fQlUpUeHjMy1Ctd9Ap2letP22qYCvavkbMu8K7IskwDksKYfgz1Ne3HDwS
YpAz4XC/NCeYFfWigCHL/GWWVrk9Cg00n+G7wsH9LGuTSw8+sc+ea2zxmz42Wmbpj40zh5bdhEpA
ooXvPaVlXCXt7Rsi/qkCgP0P2NI/SmSZoq7RsYYcD985fezcqmXbKHBgrK2hMr5W94KojWrztEzH
lihKySHjGSRtOEl2FVzjy4Ue4f3enBGNH7X3syZq22yeeKY7tGIgQUzWh7e89cc6ULYVE3/5Y7mZ
EHPhlQ10gG+QtSwi6ZqnPWpD2U+/rnYMSwS26lB3mTQ3BNkTp4K91ZWca9q3R8DzmFSW0zPiVi1f
tUysGB0nd/WMeEPn9OrP12OA5lejjZg2hm2Nr5xkliYbiw5dMsyFFYXGXJ9X5CUNFRF+t+EX5+Dt
twJOwLSAK2+COiO8pVoyOTnMYLjLwVBrLZ8gwt4U+GSCN/t4tJ5QyGJGdMyUFr2OzZbq2Ja3v5s5
hUnb+3+pO/3u6/pMtRofzkOGrv9JRMfv3VIAV/s9w4Weq65dJdkqZKGo0KBAY5fPogghupCuobhM
NgN04V6qgmnXQbQ+/cSEzYVfPkEwJajWtPx65FkBgmbQn9bCDxlU/QWKUXtbdQIo14ADqEenmnS1
XAqAGI3izg1YVJP33dPDO4HGKGtTHKaGSthxDTLcC1czxX4aDRpvwa8jX3uacyLu3MTnSdzi5gH1
ir3+IyK9t9mgLDLOWGH3jXmTPRIPpebuMSB4LhsEuoYOG9iQl83QAGQbq1oQuRCZrhmYbWy3MJ4V
5491fEnIEO5VIyV7bYZ85mUejt69TphyCgZgD1SrWk6xqrbzXmhjRVY/BNemnD0r8JMXBDahQT9J
sjhvjeblLrLvxDU6EnoIpPk0xVhv9XFqQCa+6J3vgV16KGIhQAmJHhWw1PriImTbqL5wWW2Y77Y1
u/AfieCv0H23uAxJBWb0Vna2MSrrh3/7TQbUNAWnQy3uwDCgQ1SGy6WbCAFykaSWbJynEi8qfxjI
sjKe4QDWQyKlxqH5a26Nftwy+cj5nbdlgz2qQB2v3DYzGQ6sQiNx7SwtiHFmVOF04onNLcnWjclo
R/kVwyAozC6suRPGR7UKAj4wHlvai2w1qLvbjNnQrEKlaL6rrs5B3XLW1S06LPGKzKVrEQDfYwGq
sLpafYjCdKORToXo99srQZdXBCHyPOxdK5JzhJwZhNTLDVJ1zoxG+b4LHOCR63QpUCQvOOjniyn8
crYNc8fzLwf78L6g3skZMuX5ut6+MY84x8XoRIOQbhZofp68n6YEANAslEgcEydtJlAFdUVOSsA9
ridopyl4BZgqT0+zbwNyg/83UiQppthKgKOY5mqUX5sIcfVbp1Scbf7nMi6VqTOSBoUamWvokX3h
F5yT6+jYWtpD0U2FYyScrvDMIdoVHz/9P6R9gfhbNP1MPP8T3y1/nVfxotPez9MMx0DUwf0zvBW6
9Bi1Kjqm1bGKgN5ygzRiLAYU6VD1Gf56bdRCEBZTQ90xj5CcKZ6JTIAyrxHTDszzzppZe/ZS9d4n
yfuuFCo147LreR+ilrNWNPYRPB4kVtYP7dS03eqnLgekrE6qyFYjwQSLed7Yu9JvFiP5meiopAK4
PGGfPg2TtqNSH+1d+XziXjnCfbSkYxfS/ufAz22HoOrbNV02PgneBcno+qlvOsPyayYpQcQJ4utM
utzVO6OHRzkTDHuvl4wxbLH1wNZXU0udFhcJJEGOn126yVMQtpcg//ed6/SBtVXRsgkL4iMkBIq5
yfGUmIqUbDPMC+ZQRnlMDYsgZJ6oAuR8Kp9qKAEuYfNKeyv8qZYYytD4Ezmo8D9iT+ybtAJMVxjO
MKp0ZwISKQj4CKOQ7MtMEbbCWFtVrhByJImkZsXFlkvr+4WDivD1sJ8eYJMJShC0vtNtfbUhtAo0
HJ2MGk1MvaL3C1idK0R+c+4glyLE0x37tETlhQScDUndDQizyBY0pCpmG4vX1MbwLCMyaKVnud+G
TwOldZD9nky82CQ43ZLtSeaGQam9BjoCgdRx7cspsWO5gaZWZqPd52yKVuhxwx3eadL7cTrlf0Q0
QB0d4Hirgy1skcb9g0ynTJCcGZFaNGeJllQkFLtpgtuMvQzBe8x71ESflDfQ2Zn33X+bITdPbHNt
Y1vUtMGU4dLnoJxWwk+hXPb0sw0Fugwy3huC4Bkn1NiEDSPl8VcuGvg6gIWA2VEFVQgm0N7kJPgq
qakvyXiG2Kohy6Z2XVP13qdgYGSBy9m1/mtNNA+/RqMFlD7QzMqalnTU89VHACQqkQptWQrATLba
Uc12cSQJ/l8C090963/y77wyYCm4VR90sgm2MUDSnHLZWIV/BGabjr/YXbDBftiJSCWsm7aGeEKK
cOFgC/2TgggemTMI4PMJOzcenU2fBPP8YQgSVzzpuTvdossAC3QspwMq2Kj6caEs1bdTsALq/WPE
vSZqkJW7dbJZpU24D+MhBZ8BEdyytEnrRIaUWzVq6TcNq2JrspcTuiu24TZcuN235RgD3onJmH4v
s9SFur6f7Eb/20IAAxn9fMT7DOAGbspjax/un/RYKqVOOKvm7ZQ9Qi4G4RzPt2KboDh5ekGQIxn+
gfvHZj5MWfK+G1xP+Os9XO4rvY6DhgU1C7Ah8rLHT23cn6iBGdQnJZpyadA5pEPPBswEuY/4yNVH
BQhoAalm2krT36gHpdWDokk7IMZdKeGZKJpsf9q0LHnwsVlhVENNc+y5zCY4s0pl2D0ZCgeFRYhG
+4vVmTbG7UkK4fLe7ktPRTY2/lC3bn5xKPBUodDPgG3+pLtpAoUlOny0OZ6JH/E8mJgZX5FP11Ao
73y4HhH9BdA8jXFMRcXXhH5b3KLLKRE0/N3dC+N56B3JyxtlV46K43FXrelyMVkj2zHfRjGJZEws
1n1P4abLMEuVIoI3t9onKUBnd9HPsigTzxmlXpmqwdFc54lKW+an6dyHo/B7qSKQ+h5j2MNgDAOR
hBcwYIv9MxI0WsyLdBAKpA2IZ12GqbOpaR+apIL57lhqVcH/IQwo0kiS2TufacfjJFuB5KN68fUF
5MRk2dx2CAh6GGVl/rtS49UkTDVj8YowFViDtnrCR4lPywWnV1WEiZ0qheFDGF45e6BrLA/H0lID
7dDBHbAc4JmrFW4M4Nspl1ckxTbwSv2JaP25+ZU+liRToIhewmrDw+3P1qlohgrSfRKZx9nNkpuh
p2BQp77a0vHqK8hNEQDARHFb0RqhQBAcKirWlNYWaUNHKuCjV1i1qqXwb3b9mNS7sSyyI+ex6af+
/6y/A3MEyl28quBc8xP79UXgaiavXsIxDtKITE4tQtnRca4l4kAgcT/hX8rntZ9bDTF72FCSbTO1
KN4SA0KlzY4/uDO1+AqFzMRi/hnWJc13dzc14lGtp1937lkQJUlRkImbc2MimvaAyyErmoFwkzIj
Szl4VRBek5sOOplmoC+utMjmSxtICnUxoigxz91KlS04AxUNXijAEvrC7M74XHQc0/QkEIEsGxE6
x21apEeapaIndDzsJqkdRlJOeqArW9i+SBoO7xIo4fwiSyeJ4oZaXFQ2ruuJjTyNYaxH01Qx/6mW
mHzLjyutGGUTm5EQZ661IhCsI18msEPlwUBwJhf7ONK5wNgh6x+QmDUa3Ico/16frobShzixVFQX
LWWZZqHoHk+7sm+hu2kbvjJpIlX60i9ACoU9q1HiCTcnTpHJpLKFTYIJPF5cexPbLb78t9c/mXnY
WUBD9UzRZCFRnv7HPOJpwKT9KYyertZZaIHEzc/ax4iUWQT605l3mlS8TldaIWACCrExUxvEzMZp
YLQAV/gIT/5GRi3vKa13zFyP+eLU/LjPxlRXJq9CPXskMJcrjNmyuP/8iZKs8rADxgoRI3LdEknh
28HFABup2Nc0436a1HUWjPcxvB8nOgAVbFUjqWoKwwTKllDCxrbiXExUY9GTeR7qe9mDpn3ADZYJ
zcROw/v+kSFYyusz6f1b60ypmBqX8vlmANZgxDq8dyeDO2KJ17ryhb+zAWnSuSMWVwtTVOTsP+xl
UiQTOx24M+tJNDLbwnTplTt/IoHoflfbnmZyQYzd6TdjrZFFddyzELOi+eDPLAAdDeEwzNjyquQ1
RFHMfhNP4VyfQ3KZFO7yCJXkq9ZMXupASTeTe9DMKwXO+OVjDsuWfx3d37jXEwiWViamq6kazEDA
7yhRVjrRVfE8fZcfqkqGzyteboYQeqjS8NnrdNi2JYUdlk3zzwEPaahe7m6yS+oVTmhBRck5Lk8y
aLSTorDgE19WjgdQc4w2RkBHjK7a6JNpQ4nED+QT+7N/SBSYoCN9Lxpg+sjBBnh2J0Oorg5xn3eR
RPQw6zjjpvs4HHtqWxwpeglWKuSEJ7dRhYJmC2C33pIQE2rh2z1h6cRQdI2mMwUMdbHgn3gIq0QQ
bpoloUFSFwKUQ0M86qSw20tWflHbNwUlbgh7sK+rmp+5BdtRz7umXMHnJaMdmyuEVFTLhbk2Xdkk
oyS4DIB9ksMGrstzdFeH52sil/ph5BWUYu8USYvoRMKK+AOoL9Mti+qOTRbVeB4KQ3T4tBHRZ6CR
EKuSc5TuMtfYbbL4KZ35PeG8zT6kXtfu4eI7akFzUsI9TEY0bwBhhXwa08Qx+10u8WxeY9WpDOqX
WHz44DFkzENSKeUojwbROJddw+WWyUR6NgM4jxNBw52qFzqoHZqEIpNHUKoFeo+wHrS+SRD6ctsS
DN7miKCviWSuR1eCExMEj4UfPwXhMWIEt49iKYVYrFv+dzMaDnd5oE6BMAoh0BcEoFTM9rRJGm4q
2vwvbFEhqqUxaA1w2CDuPzmXtV46p48nTgPig7S+z9BnOqSbDuB35ZtyPsr4NQy5MoBp/udYQW/0
ibmEqMlRLdDP7z+83FWNopVHwW4VvwhApjRzWo4ovkTpJD4zRlp3oJ/y/U5AiwDOI3WA2RjJ7T+u
vHlo/xEPz/RfW/vZZklie7BB/QNmZg4aDOEC2CAAPznNuIl1sorPFarmB3UQskbd4k6oqM7jIom2
du1NU3tXN9/sFENmVdLBM20B2xIvkh7WX6PRLV8pavXAHG4JmXy956lnASc85ar/F0+sor2H1+XP
Jq9rOU90r5MbETpo6xHHsHmUgwAGllcBqAFqwo8cikMqyMc5eYWpsv12m1ICM4sWQG+7t+ZvsCAV
cKH7oXgeE03olAinCXD9q3S30br8kllk+l/gQqMVXK5vDlOC69Tz2tTWyk96mddkgLpCIYHskqiA
JVN6P2YzVq+1lfGnq7ByhZxHQg1H3Z8CBPa42vfuKr2ajhmnO+JGMZLVnaB3mBdoWKdpoekfPCvI
/C6YUZFNpM5VJ8pUZxNQoxBMZRl3xlDVSOx1sT/LvlO+BrtziJUCAsTrX4ycqi0oDEBhCxBKASRX
Jxoazx9zHyuhHoGeB1rtDgXJKRyh59Jgfgyo21yLHsNSPuhw3ya8Ft7lkyeEe54dI6OqLQMKnxGo
xRMh/CLQ6AkNnD3njAEtJKTQdBYBZ0w+k9ssARopsYPR7Yl6Imqx3Izb+tlJHXPjDpity2HQABdj
pzBPnHr/nYsxGX6ZyqDSZ1JSgAuzQN1Ulvm0CE3UzP3X3qGI1Cp/jXOw0+yVxwPpafQSVwp8+xM0
ERyT6XrDVT3ItrBTNPrDQgumS5QSSpHO0UQOWC62CiVjJYLX5Rq/M6js0HB2Vwx9a+BciONFWwcB
q+8TqJUApsv9gNFsZp8RiMAU0t//zK48CfbFUfTd7Rl6un7L/x9vfFtMDwvshL4ns4Vi30Ji7Zvv
1rF0hjm9yjvOZoK9hm3ebOaBU2cK0Zjj95zgia1gXGxT5cZij6MvnuVh4vPMyfngu1V+eKt/vGrm
M6Ato30Wr/UwqhshAmK5rRxBv3Vbw6FzEMQhmnSZmbEQ+ypMRFwh1TiEWODMwRkRB+COhawnI2cy
Gl+YywGjo1vqFUAifrBUnA2aXDT1GLO0P5WvMnuGBIg0YV+AEypEhbkDf+NtuTzVyF+odCapMo9Z
fAcRcyAYDDEGOJQJTd548uSqBsbE8D6gFnzXrdLHEu4BcWGpFAO/ACbJY4/M5lD/iqCXMkpsK9pQ
e9bY4QtKe2gWrjyv4qee1zu4wbFa4xMhPA/Cv+1qBHm1SJYAe1pVJnp1S6+eFMPcX1NLEhRqKXbF
WaE+YKn+r78dhSlOF/os7zMM2hp9Gv5T4OxdLtB/B7It/ppgM3VeaUrYrJc0nRH/0SVx3ApuDJPb
KzCYltj4UV75p3A1wt4cnbL30BYhFAgBdGCqviHtdcdpqUcI+z5qWcMObpLIXIWNcKv5kEQuLqRh
8+bQd1BbK21E9SssQI0iVWtTi9zl6IOF7MgDiaujo8JIZfp5uq9porxWfhMECL6Td7oVL2q0MCZ+
URQDxNpOZ/TfHxIJzViDX0dzyrXLZKvYi72Y4HraO17eiN4ZykzMjsyRGLiIlzK+l11Dx0t1+pjN
N9Ot/KFF/XFC00pjSr5MAIBN/kIg6CXA8jOc3tMG7YQw880WZHoztFnFD0YSB2ef76GxoGALVFK7
YqWfRsa4xmnuvYlBmBb32swUtCb8PsVQpVeNr3rP5G/GSB+Z5RR1P4H36HXOALlLSl019icEeVJ8
3SVZdjvdgoyisXND1GuaF8sWo9sATHbhsCqZnGmHENvMMGTFQDEOsLJG0TN82BHQSz3R7NF3yFBB
EyxNsYrD4ZMEY4BqzQ00vc9Igtdd/e6YbwMQva7sPeoLdgL79U5qyn8V236VzVc6Zwin86aJcAyw
8VsBk6r9xpc5AxzaLzPLCIrBc493ZZIntE9iDOmQNJ86n6v1tatMzOeHLi+I0dR0XWjnAF4DsOhI
RM2ag5Pfzko2N6S8SE5sJpqjdVlYWeFCxgmaGQ9jqMY1dlryKRg7+HeU8oc3Xau8ckEhBg/dBZEA
Db9FTBbY8IH6SL53DRhJIpq3tlQvZrWWHquuxpxbOpY0NqO1ILRe7VqwhdTSmdnGv0NR56X8RKYS
1S2ItiO/n8ihR0N3kTlcirOrpGNVRB/yg3iFFedanqH+Fg6idD9VlMPqo58tPeClGFSc29Mxni69
CTtJ2ghava8bxDaNe/twvAstzLDJbtICCfi83o78mYuKqdE1UyaDhXKoSJYYxYn0roLjTBFw8PuA
NwMyR+T7dEC354raklz34knTrFOrJQeXehukGYJLaT4kHFFqShaxJeL7n8w/PUajD/bV+CmWWiq1
o9tgrzP2T3cecuaRNRjAViiweuk0zmDLtIrAoJbVzUDeFzdQAo41XM5hWagMrZRQLMQhfTi/2Kn+
1eaY24zsLqhDgRGvH7C5CFqHn52oU0C0VbvRxxk+BKrZ73y9J61/vsEfXybwENexHfvwSr0W09bn
HYG1iXVh9FHN6fzOAj5AYqXgK+CR7gcExTkmHxQHV+9UEL0GA4CifMo6/HiQVsKvWq7EbpOxgGs7
YrrfkrP3ZmvwbHCDiSkGrcOh7tUl/ucXqyz3zAU1Ag14/RuawDVCXuHE9J0xsyCOzge8gO5CK030
hxmGmmajdsmfFmRfQ4FiNyyQ39BP7eHmleBLBit3Z+bH4nyn7le8eK2VKYjSzAyJV9SPsZsTvi7Q
nebpaij0UYG0LOAAAm2nlYAJ91YGYjrXuSmIULzTtmEn0zS20LHM7nAar2sP1nGUYirzXWkXbyQJ
GfgAYCWq23ufzHGSD9HZS0AXoyOlOtrQMc1A+scNw2CEdkhwUcGgXe179+HQdMKislz/MbZ5o0xd
VWps8WU+VyBieJkd9O2lKRLSC+h49vm6vh5FLmxmd3dUOQqZie3mvt6K0xhW7ZBZxSwI2wRNUC91
0lLGPEiTfFnGlyGhgFoY1wcsO51PeigOiLAwFmvMoKlvjsUlfROPcAgCtpXZSifE2Lw/qtBfzpoB
+1b0TxYw1tSKV/OFA33gS+OxiWe4z/GT4TZ1/FFPKtrWdjNbGj8tW80S1pKxv+rSfdY3Nm60gCyT
cyIIYOcMg3jh+e7ZIrVekz32WfSJgo7/REjH6lavRjtDtXp5VCoM1VQmujk2caNCdjth9MQaVWuJ
frqFtUsExZg+ihdkwhDYIgvw89WBO9500Or1tUtXP78BD5PECnMKd3bOSeWqudSsw3c2qCnjKkBz
PmaVq+WkMDysZRcIJlD24VpEh7lKHWNyR5xuSfzn1Ugn8ecCS0n8HIwKCRORYk9y7WV+w0JA4Dq3
9jIeT+Py+crXp+8+LqCHcupxvnzz3b9CrzQLrfx9y3ivGKGd84Q1X/+BDh8Od/TgRW5Pyvcba0m6
6XoQB71NtmuquKY41UB8Bmq7Ph4xk1pF008pPLxAC7IFmV3ePlnWNog6aZuMiR3ZwDJZiY+aRPbQ
Dv2W4K8TAXZrI40y/eb7JTumIuY7MMiYrcv8eMyAfW6JvhKCVS8k1UGIsR9cYKZpD67FUI0t8Mb4
VfeqeIHq7JG/uhNw7NcFaD3M4530FSPcgaST7Y1prvKpdrjOhTFrwMyiJfrXV1B+YCzv1QkGM2Ql
0PIOQs3iGvBoDvQINLPXcemammUp3k5FFB2gWRZc8FE+YbeZ0tyvv+pVh1NLTdNbsFCHzT4RbApa
m5jf0ZA+4DpYXNSHXl5483dNCZo172G68drdqh0ZBi9oZgJblafOEmtu+0XKY2l7xmylgk3URE/H
+TeMTG5pglQx/hPt2srgKHHOLKaIdOoQ7vsMjZEuBlg6y31W1CZFnI2LsRn9SGSZbo1uYmkbkrJF
80J/bN8BQlHboXmIzhWAk/sHoZT0hv6Ka90jbYYyXVr6VMWyUPBCcKhvcgeYpGszJABqoq/IIZYD
Ki0SAntIWmPhbv5kIX/6DISQNIrxJiHQp/7+iOwgpUtN0mnkW8+h9gWfWPd48EKsB67eMLe7/dNi
II7+Ontfge1tTOub2dqjyUE4WcTRvrxlrxeISxTvcS+HcQNtCb+zym8tr5NtXX3i3EsFDaBDvvnU
J3/BORZivBoP6Tm5sA+okQ7Dnm3/xZ97AqZmOJs+/FuMWaeldyrrqltPC/jcqXbo6r8w6wkEshWb
RQzYcJheH9dPRH54NxRAe3q8GGhIRIguAfPS7etcdObpY76xggOwJ+bc3ZPYHUqBA1bmmUn4tb3i
4WyTu8FTA2ITL42wqMR+ZjtMVfWTVNGmfd7ntJVfIY4RjWeI/H+YIihsRiNyyzZXP5x+fQA5+jAx
N+S6pudH6G6Aqm9DD+wzndCBwtT0xOqEnxKwt6woI07c2WIsFxnelrG8wEvLYJX06XuqW74u1VIT
DQkGePJ1FtC0ef0gdcVFFexRXf+oUKcZafx8XCrbG/6dBtb5q5+OIE+gcQx6D8KEhubvappNDS3V
/ZCnCnWQJHdLWIPgvuI//Bq0t6bu/359eQ1fbdqbrjTRzhQgvds/jXyT2ILwlFtGJ7nSXluEuhaT
lejbd4XzmsyW3lIv1HfeMIWA37q10qns319dcDxJv1q0qtaunfn+0JfH08/0AcuZbqdqppeaF5uD
jThTMrTobHokSUTPvf3v+CTzry7Ngu6ad/ThXj/q76dY/0nfqORPosovVf/YTo6j+1g5IJbeW0O+
Kw7N577iutYGUznVIN+GN8LF/BmAgFEALuB3xUSLURTMq2h0ylE2ikp3u34WgF/ClsUFB3+gJuzJ
8liuSfpp0f2rVbRi4mK1qq3FRzr+yca0beB6c36dYczirR0X+qc+L286ymw1Vadnj2TP+dTlbzk/
07ZsB82kIH8sXRavYdWhfS4I99R3cvd36ZbDNIREf2iXYc9VwcnemeAwp7Z5MqrUM6wT5xont/xW
XhpfAiHZJDXNqMbLxYndNI14eZCa1Hsu5eCoA4y1hoDVLZ+dTHgi1ujn5BOK7iSnSQUcmk89qXDD
7QOPE8xZAQMXIiGBm/X+4YLNeli5DN1BktJrs2NcV6uAOc/Bbu3g/zjpiekWFG65T+f/OHcxvlmS
Cgdk59oGsl3y10uV9ur7wMFtiorhQdAvYb9SGTQgJ+PkdHcQmLYHGKQFJswhiW8JAySvU/aTq4tq
qtrJ6Xr5TojzGhxZO8WFqc97zPoI5SdrP1gjAHl3MWtjc5MRKCoPh9zz8BGg0noF08v7o1gMcxlC
HbIYfXW7mdpGSwtKX/hKOsuxnfuCdOCbE5YHttGvFMVwipasn2d4SpcdkJEL4LUxRxDkn6FyHfP/
dFXOrKeUiydsp3qyYPvlW5zBBrGeGKLXKH1yrsdRUVOVb09xRvrZnWdnFzj/YyH522MxVWtWXkIF
ahwlNr9SX72sg+0qJMUPHvc/FAXGzHyAm8uQMwuODon/IWuTr88PA8D9dLHFOwlZohCjlUqYAP46
p+yj855vOHTVzMH7+hIOW4OYAOLO5CGX+J+/E91VUQVwrlU/6xaRAqEamHTlqEfy/sA1Tu7ESm9G
LGULI0xSUl7CSkR7ElUCQpL7lTpknxNEUMoItO/3bGET60a89zRI7hqICFGgUW4reF8RifUX5hVP
F3DTt+hVtv70gpBg4Jbk+jxvYpkXG7zLjfjE1ZfyVRDtRGJTSh+YDvNK2FX5OnixvDILrEp86PPW
s91fTxKZoifF5KhgcNcZ4O52xy5xLWsFh7BjaK331vde6xv0Vg7CG8AiEtMdp68xmHJjm4ArtQfo
u6qXE7K91yKaOmL/eACYLVoAEB8SvJpZexxjIjW6tSbRgkHfSQ5nzEkiRgRCHKMy0/6k9YF2tDtg
YJWJY1qLY5/mtKaa9lA0HJRV0jwmuF6n9pkUPuMPsRCpQOC+Pg/QUe0+2Wemomr+iA5NeyF+sHDn
PSNx4nTBDY8tPqUV0JpTLG0OwnA6utHPHkNzbKgvtZK6cZI8h2WL6f+0A6W1vXnJyzLvGaIhOf2s
+qM37XfC0hnSYYgxfGh1as2GT2p/OErBk6aDvASr0g23EjCtGcWnZEQZWr3Ey0zoJp2amPvnK/wI
nTaw1+wqslzez1Fl6sCe20RMq9bi58JLv94rbxadCpsY9+zattUsLt69nRFJfuVJDRaEmizQA2Ln
hl+PESNxYK2HfGbZI1Y33bF9VfvPPB64Iug9jaYIZ6suHp1MgAysLGWOoEbN6mUB4d/kHzcAV58Z
U1vT8CXoPHJJlwNcTU1x9iTcrbCfEdvWunyrHVFRh7MWLP3LzE3Xcv/peBv2CfCBqu8eL2M3VLmD
KQDQGS5VoE5Kjt0EX+Z6HPepTqgVKX66FTZJXG0TWOt7MT/Yx1L/4qqn5ADnuNGk1WHhvW/C46Du
n4qgYmbZPPc16dN7ijqsygxYDjbrpVp0IeCLRtcRc7SnGlHaXBngU6ZEKSgyH6yXgN8WethVXl7F
CJzeC3LKjKRrutFaPJY+jTXMJcRoltEKFqsye6laGd7xh7QOawpcSD61EDBYZRsYNWAuN2/+B4dQ
i5s06t9FUm9LT6uMKaaJFtG9Pw7OcAj6vRwZQxAErETMKph03RNzD7dAolH/ESHe5vOugCmtHE8m
ANwyJx3sJ+hLFbLFSlQuSgDkGWk1nPG5P4PaWXDuRnptWstTGpBY8oc8cqtFDPASiVX6XZtP8szI
tv1/z7wIBYK8aDW8yDKYwshQkocZUpTZJWGNcHPV8VKWprwGB72bI1GljYdcORJRZkzeXDBbY4eL
SmbnEyAGnDA+ZCYO4aY3sKuE98fvfdj79Yn8bwqypuBrClRjVc9Z1NgPoq0dGnJ+V0IazOtYQFYF
PVk2MT8NznveaDP6aEdO/dCZpLxVJo9bEqYWXPR8D/J1iw9EeY9J8Eh7XK3mFYy0Zye3k+7/Dyhw
QcUSXN+JBA+UXV5SnX4xI2G65HfCDTO3tRVn13pwjVYrZ4mL77S4UR4p03X+scv625/AcmrynwKx
ZG9vm5iBJCiEAoj7QEhOMkk7Ku+IdblcsQ7aWpOO1SLIOuO11zQuHrO6gDoPuC0HUCs9gi65zguM
eWmkdNqOjqhypyeiiTcld+IyS0xyLM8jXAxL2pbGoXWE67BiYXKLimFwPeH5HMUcIb9nrpRurVi2
pEcO2YV65h5CoHicqnrg3F40FCa5efQx0xUFSh2sRDsDoLlr5gAAZNNqHdAxzxmSKx+B7OvOXvKX
YFsV90Bh6y5ATLClG+5Jiqrn4d7/nCPdUt0Q3uGndihnu4nT4dTWppuK6VPjwP1fIYHbn0dOdp3M
pReQAMlCNzswf2ja8WRWxYzmRPX6qy/nKwR8d6tHDX1ipMJrndDeZQO4JYjKUcM2SDrAVMj3/GO7
wnJA4z7+6DWqYlBY7SLXOi/VoODh9Nz3Qt4r+LQOUDc+NSUQdWuMVCTOVxAeVkV9kO4/jWaxyqVI
ygY/B4dncY0RX6uknXXrArlZIhEgBt2iLuQfabEvA6KKrybNAjJN/qUgEeW7ndzFIzoI1u46YI5S
I+/R7g6xgjXKGB2KPEJzLuLSpIrwt0Rc/SDreUYwA1nz5sg6EC5J1Gb/WKPr6KSw2hmW0sYfTqrI
gn5g7aX18SMkKvENLWArY4U8ys0ykH1JGb/ln1W9h0ptaKCXapNGJHtbZFftf+YW8FMEMwIzzM03
LnJntuFwr82ElWzC0BkGILBLh0XxAeuzYkPLZi8rSio222wcWYAIKvV61hQzOkGYjd7+rtXRidF6
Ijw/LoqucYm0nTHGnNjkksbkzwBWmwzSd3NtmW+VepD9oyuUCNh6sBizsdJP30Hr0ELOFaO8Iu6/
mW+TlnXNBIL0NonUFD3J+cK+ZssSaIDy+XyV5/YU39ggQpPGq88LafhF2DQOqSHVSaaT3diJKzQ4
ethOMvvv2ySQnczKbGH4xoVXP/rh2BkK7uoB+7dCVtLBveR9HhL1p8ZOuCjfcHLiePVSGZqW2xYh
EvICatJgguqydrr+DTCN5dC8hQH1NfdD75qY2PoF/89IK55jUUAHtv3VIhPLBsRSPf2Uuf9RTeTh
mBS8vzRF7GYIwdzu8XVDpmgmv88Juy5TZAXWnbqto38yjkDZEUbaoHoWzlvc5RORfjWXfjPhkAYE
hyDYqPaWM2QpU4AsszodDYYuckjzoq0Dwic3mN+UfCRFbgjx/PZ7bWk3W96p4/ewRoDdP5zgwSky
M2Ro5CfVQeI599VPEai0o/vckhRCNmVZcI0ETPifnREv7btVuNwfyFJjIsSPSDKlL1dIKDWqclZn
83l+cubgypE78GmO3fEwEn3gRCz55GdrkyqDafJLaZ8/muDYsob8MQmA1LQnz15AxTbwJOWwPaze
w/9tSgY9pFLXJxg1kd2dISk7EO+jbXlSnvx/pqrCAbxu7CkYhiLKC0rtzoO2z9FNvO+Rwkcg1Aft
6FNdABeS8my+24nZTyU9c14KT9TmqdnqNQlWcETJiLmj9vstd3nEjI6oMvLkn/URrjfIlOq/xwsX
/hLf9vSwb0e3j5uPqCVUjwm34ZORD4wPUMtrtsAjJ3+/9TDEuUY/6rCMxVhuPMDPiIEFsFWcJv/E
Cc6MV6pqu1+3+1zCzaDuoNy2wngpj6or8qTLEySouQvFsvp/w3yd9q2gCjzsomC6NDb1zvMTBV0T
hK79P4yL6gaoRsGAybX1RkMpySZpq/3632fCDn6ra1Bro6qjPUQ0ygkwHeNwaVazO5f85DWGLY0P
LShU0/ypUOm/bLorfQ+HtZOPLR4TN5d1TWpRoj9TZwBvaRH1coCHq3Lwr8PAAPu4pndq4q+h5eNH
2lWPISRBp6H5nQgupKXr1DxjGgeiXH8F1DvZaOtnbYyeU8MEp+ker09lcvIqgBvXnnqtMWEM9sLH
a7Th+g9+5CFYMHAkBso0tnjzDn1k/fLwlgrVGu4tn8ubM+9Wlj5L+j1gxbL2GymcurYvRBRZL6sJ
xIj/KayB7nPp90heV+yZMZQ6keI1K4jliDDy0nsT68ZkjG+y8bqVWHw1fGsuJW+8h177fPZxiUw1
7BIsFm+yjLOp+AIRXSvNKVX9HY91ud/XzUyhKBsBUxY2PBHYFrch8i4BQn5vjiruh8WkU8zGf6sY
Cgz+IuicbGkNOQfE4cU7+dZgiAIqWTaBN7NRdxdRGdEFIYHg0K6KtYN8TISP2er3d0UgAFJ59AZ2
EyMCwFvyGPInCoh0UOsvKE+uzK804L4TBAY+0Hv+6ZX1qrtWBi+qk8+OFk+6hHUw7nD8j9/CRPId
IU7hP+nIEe59NAKCnqH8lnSFM8xOxbzZ/kBIHAEO1tn1Vri8NheygYOVCR++bG3z5T57R8s0wumQ
qHOaWPd69sEUkcBEcTAdGOBJ3zbb0ZsmkuntAoES6XVy+tt72XB+aBkmXefzLvGuNRQ+k3ZOoFTS
kGxpkqhdMXuHieupAMAg3ceduQe1ML4Np2BtWiT07WgTNlaTm4u2CK0Ln5LhcZ4ldG/SHFEIk0lL
2+sih+oOT2ZKvlVdaEu4L/VELaHWdLHRD381leZJ3XqZmXvsbQCu9vuwmhr/vhHAS8WFDUadWLw+
c7Mbg31e2PfDdK2zOHo50WDOpQS8to6voULynG9mzMIPGiEUTTE9Q26/mYallTZ0AXV9sGRxlibE
z7M/S/9MDU5rpCNFoIx7INVT9Lj+R2muEf/AacLoFA9WpkV7Y8KOnGaZql7Y8G4mJPTY585CWMFs
CFnLfoHycIWsU9hube+iPnCt8ajW4GF9vsx7PEFcrvDxGC8nQbNI/a6CKAKCzxxCzSmIvvDmqwGq
eZn9B1ELeNE6O/ytI4GGSPYH+7jhosYR1UNa9NS3lhy2cWbiyYY80NShGojaEcS6xraifeCaxWQA
GmeVjHHWIY4Npl1DcOsMfvJxuwUqIPcXB9Oafp/VnVG4Fnz7GUL7JdjVInOHuC+I4K4nTERNEXQJ
S8NAi5nZvfcP5xjrerkO2T5ANBS8B6TpHQldeuJXSc2ueKYSPFuM8Tet4UzF0V/dswQRyTt3uHmd
GK0eHd9VFVnNi2DXu9bAz9/zDdysBPmc+0zGmnai5BSUparGbpWhEnRTPUvHPdlIpy90uTkfg559
oZvepYfa5qLqU3QluyLO3VRW6qwpMybIWKp+IrkmWfmaPUOO4x8btRf19HPgkaGok+7I9XvGmzSy
sjrBnXOVFZsT8xY4U3gfUAXCfumspkfX1MJIloJ1Oz2Cz+7D9i3b8nerI6uK6LhOH+LgLsJjeTwZ
VsXQtnSVZs/zfTVRV6vpwIWRSKjo3umLtwG/ocFjAH7n3/rZzWxphHIqt0fzj6LVtHt6D9ivbH9k
hjGOViRTyYd6rLUuoNM7gAS40+0EHkCjr+B7OAe80BfOneA2lYnK6p+B+DG/GCir7y9quOMmUsRV
0HkPVXyrVTjUMLBa3SWWckpoONKp0/2UlM68ZpZ6KJynJiRPHOWN1LrM0S+NBaQB4OUjQEANOd4/
Lg3yCJRXtfx1DaT52EHv4Y5q/tIEGujnSI8CK2NuFX6TqDZh2ND7CYUSztWPckRWYCmhLjQKrmWK
ss+MWcW3SRsy9iiwL1jYNHctyVJMz3WK+OzYek1xlMqEeHP/0JGIOip+C/scYfdsOboVRjQavLFw
8z0Nq3taYtXubxwaazYbLD2c4xMtpFhvWR2eUc9N4H0TRxc8WErkj5mzN8cNJgOYxU24p1DPM1+y
GAImDDvI2c3aG+vPI9C5IXkr9Dsva48xUghk2eWl6jT4R3femp1S33rMhmZnv+3+4f4urGvMHwby
pEkYVy/Z0WCYA3840LlLG10ieGZER/za29P00bkfr6tYfzXBp8MKbsol5jnocnbiwuX+7q83QHAb
xBC0pzGV4LkXuXln1FK2bokUgjCzDuPD42r+xtZQbzb2cjpQ/xtCo4dWlFnSE2sbTbq+gp44hnHN
VJ/92Mmztlzgg16dFb4qnlW92Jkyy78uvyNJWXxfTbfc49tjVJbuh5P3ysVNTzFYTV7OxEVuxlIg
54nRYCihRHkuOO0zN0oRU154mi1DPVXcLuAkkhTvzjRq93wjCQBFwYEgCbquoDo4WM1qO0OmP6NP
SHy5Dg6U3D4ETG2T/lfFhOOnz4A2q7+4mi6s/XJ+T0ZZYLR+w1ltfYtLtM648cRuFIgAJ2xOf+Ax
qUwIfsw5G7n6SN7JsnKR5n59Wc1s2dSGS+Q79uZDY/Y7MikdA3sKCJfVG0zNgPwqqi1H/edgfSLr
0ySmced/piwrEHaE8gApoP3bOS1bSB6+k1vuDXqRN1poj1ymZFXH33BWb86brRLY5L/7TDknSAV7
Wmv9Q6Wahe1zec6PpIpMi3li8J2GD/2EMdzcGBc/gfRSF4Mg5WY1TL42ClwlUMfmCb593PCHncG9
89d5ROqeauhKqlo22fTYgUg9dZ6Uv2hYAJfaO6U4Y8dSDdzXvtQH/HjJh3he1ucAQ3S2oTtr/Shc
FWIx6Zhose06C9Y9adN5gynhQIS+5gCM+QVkTKNdsBP4gIqiR1ZwogBn7ZPZo9utX7BbulYISZmI
wdNJ/ieyqBbFnwrjW8JG49oYEFTZR6oCoALWUyAG/4lx9qC1enrA5/95t7RxgCcx3cBV4GSGPbHb
jYd+tIU6G56MY8GnhdZrlXpNAPvkw47soAt7TrplNKqYGTW7hHkoPN164Aps9/1oWgyl82SKUe39
4uniByqquZPz/C4X8pMSNHEVB2goDL7+nfpyXUbxHBMr4v+4sJQ+FwZ8kRjg8dq3E2df6qJiNav5
xZb4ZYCU1lmTvK+/Dv37yPASET4rxpkLLkvlLyn/3XPgIWJnwx7CSa7GEJYM83TzyFLbC7OUCErX
5QMBYKuLmWP1ETj5uLmj7TzrfOLNYZriERD5eoE8lT6mSAaBvBt6X/A7CVE412CMwgw7KTeLfTS7
MoRUhlmab7FKzGkg/05JSrir5i9jsymYn8bHZwHjMjjNdXZ/S3O44yokdP9Rnc8bL1knH1zdNCpJ
QOdlfEUz5ETIGiQ71gPA6JHGg16eUVmz/ozrdXH5Id4nyZhYexyaE9NmNe+mN3n+hrj4h/R1wzfW
pcit+AHMnJ99sJwguXqHe3vAI1b2D/JZ9gmNb3HA6NXc6kcLoWEhk8dU6iFRqcEiHXSM5VcD9Ivf
IxAN3Gz34hMH9/P8w3rlliC9cPlGGmYxkiOY3b0atcG64mFs3kuKV0Mm/Tz1bBWn4aDFH4caePtH
/t4XC7qesd352K/NAbVNVBV885IHAIJ6QUfkUXlftoD6GpcM67CDZw9K0/7XqwUIFkP3qF1gAVGI
Mixz8srFGKqxHTwfQeMSaIb8hRFlmeiireX9mA3f0LvO0XYtIIhW0X0eky/SDzCdlrZbxu9aKGHh
ik2DCMXfcx8ff7UTGtpUCupXqBXoTKm5RAB1DQ8h9rUL5VmHnXtu/iQmbt6TeF425ppkOzRABkIJ
elegS47w47tb99n+B5w/DYsV5vMcdZD9oSuSc2NvQnr8/9J3t9iApW1vjwR9znvcr4TmxD6mNyGj
MmOdOAMmLVUNi+nETreqM37U6TISOb93gAe2Lc9vTJCc8EHAfULHKjGDBmxQXWwGKBc5fS4k0uYy
F6C3FPvy/vJXZWtsFhpHq1LTA/V6WkdAhSA9Hhw5A2BCyznHMRmWmvzi53QBtXHPbOvCx3bW37HQ
11IdCc/oAitYdyS8jXCL7AQSjK1MzE6ENdANoSib4UbahOnFD8Sly0Ft640O14HJv2cKYRTRc/yy
B/SQe3MRqwghkUWPODav8PAtddWiiv63lavw1CjYy7bjK41Bi2X9Uh56bScP7XTRAQTVqfV5jlBM
uGN69kYsk+nM0nJbJXDWE/us41moyvw9PvRQ9QcGvsldIGa6Xk5OnWA7Ljz3UCmreP+tY34lgSlb
1HSmVToOFG4jRc97M/YW+SUtIYQ2PE2uxgB4Rm9pArRDpz60kYjYoh53sVBsQkJrjHbJRHRljMJT
v4Y5ts4rxDi5MWFCEoN+89pxEdRcRQ0gMgvIaGjWZbhSWq6Hp2fhBX5Hikj0M6VVhJ4kfyQ2XOGY
EBX9rtcIJwpyIP+CKS7kfun83pCROHmQdQo7Q/N69nj8ypSF0f0a2ZFVFjuB98JNt/RlIe9PW/RA
AqtGFiDp3zIhylnA1DuBBFw5KgNn1NIwGuBLRFACKaqFjlWcgHVx9QzonRCIZebbw/fS81WinfGN
iGnoEdhXWwW/UIhTpP0lioQ+F+5ZDHlfMMWu44R/uQnqRVUALvZyoEyg8wk0DotawkBRiluI2Hst
pG4uut2DsSqQVCsapV5Ewf3WzZQI4KDAaH29ml9q922Y/loDRg28AC4JZ+H2ajjKWXgaaBJ7DAMg
yEKDi1BNcZ6waf4qcKpk6f9SI37I5WI15W7FdgnA5HcbutsyPI002ommBiYZLC3HEaaAd/elc1MX
N+QzVPhlttkyWfBxfGv40On3SfiV0vcSJhXc6LjFMXNqa9wYz6AmtAjnN2QK4WHcl1lCC4FTsZ7A
uYLtDXADJbMlvOQkCIh2rTBpzKURDE0qnzweoOzy1FgyuFMmiA4abbvkcnvFJeH7XU1c/C8k3umu
7n9+WRlPOVR4loCXP6JvdP60QaX6i+QIa8WPWyNC5jGyX9Yl37+Js1am1sLPV0rY12DKFr03vly/
Rfe0IPeLPyixfdLu4YGZIiE56qu62roarGj0Qa/3Vc3q82B6ijdnY429BuFLYUmh/dkzMMABLwgH
+iqjhUIMOKpcahD2pQ/ZMmwfFsz+NzI4tiRoTbvSwjVe95S2hF8BlKZoskiEJxgPWKdyH+9Qv5mp
8fYIwOeJiDWNM7mfpN0YcxGRJIrxvDgyieJXkAGHH7SpK+kr21fConQ9FK+EygKa1ye8Le/gdpPt
MemDKZnudCLz8EfSkfwVGQZThUhPGB75wsiXi00LXKigN47q7ofQUTL1EzfYVvgxrrzrEXFpXAwK
AeAO00X6Q9F4BmBco/eflxQKgtYxW38fMnKibLZUBY6wwaLMnOZ8oQP1uC3GUDT2COgq/sxT14YC
AJ6wYThXxDagu7jcrz/MSIQFA8kcm4XpbvLXyDZBPbk7kQkHytg6Joh2+iF8Zb9cyOdf452nxogz
sbegX9OOZA2dM2ianck3c79GcVreH9raN1hGNIOSJYWtPo+1ndjdDaWt3FNDdzySW6SgsCc6DeDU
DoNlDmQZdtz1BZE0n8ALVEgd96j9Qr/dJWRtP0tm7RHeyAJiLbaP7uIYCkIYCiZXEQ0M0PvMXID+
7nGjDo4Eid/5zHLgy+xu011j4WrclVpz5VJ/W8CDmDTlOIJlFPPEpX+rUJFK6xpctODDMBQeYsf+
nEmNNEeu/1WwEFi4mz6VnHDtGCvRqR6j9pSBfa28Pq2cGCfnRVRmuQ0ev57Ux7w7sQr6pkZUCjDM
VhEko4bRA0NIRS/YhtznETs5Q64Lv0uT6w0OWF5OHC+sCb2cFFlL/bzMlYgX3ZNCesjDqsuqb8ki
XyZvshYHUDdVOrjyFcY0JEw77T1fWlZJDRhwjXXtjh/3tustymHLmfmEcBSTQroZ3/0yGMSvQIP4
AO8K0WDsDeIMfolMQYBSk9ZvbKEGWoLkMcOMp2YEnLvJarXW9cW4+Q/OcThVU/77lc8wv+c6ASUN
6Smtf5YEn4sgGHAAC24LzzmHiCxe4bpzxptLU985hJOf2L1NtdWxcu71WdE2GjxJeCvHlk/PpcVf
Mml66ktL+5v4TZYdAjHQ4w8ykPREKyGO3yrmXoukjIbsPz6csOixwiF/OGPqN61DIKCEPECZtMlx
vFDqbmcROuz1QvIab1H+JE75UvXI8ScE24XxguFHH8BPxl3ZD1zhmLPjmF0XV20kKZucIXlxOQBt
fQkTkUPMsEFLybm1/cEnBh+3uPyqpzK2B0Y+hAZuoAi19e/bb8jqiYEDrT7MLKKFKbgdOc1RSxDB
DP+kWTLZqhyDQ1TeNnfIwy7HfX/rWbx8TPnDCsBnruMvEA52+rhOiCol6rjA0jZUCek9XzVaMjPe
A3wJRi4bGgA4h5t+dxYcoUQrKyQXsP662afBG1IKPR3PR1kLML+XFKMDiWBEYXR7prXpFBHsZ9tL
r00oRoamHxRyE1f9j/joJoSlrdztmlk9Cf/0VEAMH693UkBI5507MN9bCodbbB7lmTFcwcc/SfZE
5VY0RuSRIkb5Mr51TWd7SjL8ip+3MpdkiNYtte3IgNeNDPmAyukznuoDm461MJhdkVsNhaYpJFKl
YInKqPu+6X2eSfFqjlacyLq5pPC8gMKFpwlllaPdMuaYisZTPzbNVCPw6aC7vuqvFrEsOOy+RNO7
pjg2Zy0pPM6LE0c86u8MjbKOujyAYokfnT3Yd2DKhjy3FQIuKVPGiQCZ5iBdKfC1/m2br+wdiW0W
/VOEhQcxquPkrm9BpXYwRlfeJvSpN3VIcMlwJb2SwbDW2JVNhBdzZDggTtVkeMV3swAR86WwnA6/
kQXpTzPIlb/nCKtiAx7axjFZVLciAsjhxNE9ZbX0f9WiibNTHVC8fn8S8pJZZy5CQDBaU6X/eW5r
D97q4JVJGtREsy8Na9ctNFLdl+lyd5yQUVJkMXKiEwNZKADO0SD3DZQfsjIV7xRC7F48jejR3CGi
MrYm1Ml/XKe8GMBfM97Yx3CcJBnVifIQyTvK96Q+nOGwVewbJQCMNs81wH90V4fyVaul98D6QSuQ
x7Gqk9HhzulzHtk/EjUyn26t7EMIsUP6J4Kxykku8MGQIr5dsjt15FvmLF7+WQdotMOA1CwmNSIp
gl2mUUebi6e9sE1FZwylcXKGvnBzRPBeFpvKdrNkPpVAAo7k+GAt2MuKmZxQAnh6dd+uFdM8BK/+
Bf3mJ6CA7fXSFb+uh4/bN694u8XdwkqAftTB6oT+CKh0c6gE2EWjiIgafjSE+6GhRoLvgpVhJvpk
pMHj48b1jV1gPoF+K1RjKOcUR38ypgPzYJwy7H7nRoYy+SfV6DBhhUv0EQLPTlD43+CYO0C2y3Aw
gK0vEwXuTdA7EdSpgOM60kwSrMRf8TR0OavApoorEnmdHZEifQHTt/O3+uU6iNwX2WNqManZBN4u
LV+nvMKzI48OBPaZSO+KSIKMh7WlZJxj0AjvbirEcl5FfimrpHO0HYrlOHdRwKSH09QSk0SZhf7W
dbqRoTuKBlEcxZW8dclTCjjx46YPUNrG+PeyyKZoicktEcYbmnAED14H7Imy6bGdLioQAL8UXuIe
3qGu7M4Psj5rEth4qyyzy0shimssJkZ1yo7/e9H9FOV+3EUONrnWJO0BZwHEu6xH/ofhs+Z2raQh
D6z4q9P5A66ujxUwpXCcIXt5XbhYXDCtPhUzK2hSvswebcqXKqIvkzRMvChiJChTeaEUtELXsXWG
A1Eyto46F7Ppwwg62o2GCgeETqcU9/mVOjB97t0QAyld+/Wy7kRpqakt+JH9mq/t0oMOH8Dkbw59
Mfapmwa0tAJyLHRPmnFG0irIrGIC+SVQKRn/k9TICpRRzuKOJKxjkEXC+tsOEq1tE1a4Gr+Gp94j
XqAk58cH8hplK7GZsLGVQKiDY5iCXLsPGCvxp2ZIc2QN0GX81ddMANgn0h0twKGUwr4ekBPmf531
S+GjFbeYNuK3IeK0D9g+c9/vN4/F9mg/zG72/pPKHiC5Dwe+tvdDPr0A6118wrI/OQjMsMAOnNOT
N92P4igkEqmoz3XtvZhM2PlAgK9CDHCGspIjjsPW4CHAtKAYTYk5iOt8eX2eACnO2syziilc/sk7
DFTIgvDApC8w8nRVKIIbZ/0fXf3/6gzNcYRfZRVwTOAjN7KBqR/e8/tbLDP5FNEPhpF1y0dR6s0/
JwQzN6MiVJ0UfHOPmhxqxmFkYLTYGsGzNMj5os5+4xdRr/xvg04MxRHctwYxt7D8uiPkAieOkv85
m+ke6uacPd8n1Omtk9oGV63LzXXgCj1aiexos4mNAenbKKAJEHhUG8mLEt60fPUaAvQas0yFkxIB
BUmQvq2ErrCnX6laRWha2jESrObXEDpvZI+tVM4L3a9JNX4lFK2JKI96q8vn6LQBFUDKbktBZB0R
Ra1s+jP/x0Dyi8RKa/eJyM0UAXhaKgSitf58v5BcW31d/bu0IUpdaZbL2GdEHsQjacuNq6jSmOKJ
VDELoDx8z+0eB3rftYz6za/XmDWC6EBM5vdY/CCbK1Y6xfHmNhZMkLkclQuKjKy7VTN+AIox1vek
PAfRYDoQWPiPMtHEWT3T2x2IG5P15vZ1CQxbTWH2eSPOx7wGurvlS8r54jRv+JsbA5GdyWGU937l
+ERAt+TgjIYJ/k5/j6O0NyUMJuzVTsGT0/BYEBAUHUX3ERMBdD5qCh61dvCo6ObzfLi8f3uOkjq2
gzYTJm2kwBedMwPmYTTrT0gC8J4U6E2PP8Zc4VmK00iOqbOXRBinDTZkKWNx7+I+wLZVvt2hNiGt
2NPi7dpA9Kq5wGRwGixKrC49tlX85RD8EMgdh26TOksqyHN+z5tjtchVNjfoRrZcGYTO9bb+yrrv
tzsRquQKGz9RZXh4AFVjv9GIAZmWYdklXDAei/Ze+cGjRyCxwQOBNNfXupliVvKSyYs++aAQ05D2
+XtZUBycuYcTPZzLTYiqrJSqsTtWubfSqEOghojdk9VG32jqjpx4VuEbH4R11CReQn5uFmyuk+YS
/8+U6wJ8SZoDiTCFyRZ8y7pPSEV9hd96YRu+bxrNdDcT+WcswjmxH8TUBtJ11/L7M+mKf8oBTzwh
MDHOV87DnH9zTMy9YOoKNFzPPa21jw6IChp26E1G/ytVkQEIaLfnZ7Gnp9A6D3EMhP8bhsn+7jhN
ogSG1eZ7aQ13hjKmsK4vseopFFBDwjikFNkXNy4+QUO01SY+hsvZWEcOChF7xTkYuhUzTLkcEYCv
FhVCNeZlHAEe7bL1WkQllBFp+sOMA8rkg2dE45kawQaDgAgkPZMshqSM4u1mzWK1fclxQ56Fq1Ai
HJqCArDbiS0ttb8rcuy8rn6vtiGbCYNeui2Scp+2QoK6sYFILUqPO8//tLCE1sGyLaxef0KwDd/z
D8Y6MSZvDO+kUpG8gtmg0f2HiduvSh24n4X5n3gzcyGlS0ZRymmw9rwaOYg6qQ/CqMtlWyfivVTh
UnVg3fQq9UGIUYoTNHf08fGrZNRSbViHHAIBNHa1D24J8dl2cK7RMCilYlJY/7RUxMWacwNqhGj/
4Mr+jADu09nr6v1GFeXGrxy96TOwfB9jBaAkQpcBm3DGknnkwUJKAFz9w2aXooXZgZpKOiyIKoZW
FY0Fbk21uiVCfjPMLT0cky3BHXU12HHF7Qk9FlbrMX0feCQQi041zpLCg7SKEN8aU5Tgs5TMVY/m
DyiHuD+09bTYZINA2O19CcX53Ni6M9sKNa17Yojcg8c5As1z2fZymcHq5mt/zOayQzWujPqTBqQb
SuUjJD+j6HbfhVCnXpxHQxm1UGtGpvbE6dt72dT3P4GB3I4onxGAN4xrHgkjvh7HFMGkEwOz7es2
nIh2NbPZFskT7uRCIPXhmiW9HvHLwdptfiIsZC1ObA+lr0uA/opa/6J0TvXXvcQnEBQtWI5zlvyx
eUZOa1nwhneqbn/a8J9JJALNk8Zx9uZKfwb3piPtbYuV6n9A8NfpOa4OAa4DnP9Bzc3hUF/GDw6Z
V0HveAKN3VdLI5F6ZwrvPHqEzxblyyi36NvQs4ytySLlB6dV54p9c2DtqUjXzEeV6+KUyW89ZmNE
TrjeOosHJj4oXP022XjsF4ixgTqKMm1bMNAASPL/C/PG7YG25tHgn61xlMXezGDivaRymIy3bpnU
PewCvSLZczq9zIDYD7k0jHnkeJRn+JyE6NNPRzXpy3Hm7EXeK0SYvC7njCbdtAHxkz6Jp/GcNYTN
xBtTodjRtk3uCpzQIDHfKwffxbAv1Avpfoih7x3ApxiUcaLzbeq5yH/u/Yrhq3fimTlt/NrlVJBt
2lu7BzWFNMmTMiQTVwbmeMmw2rVxglKjIWeyF0PYA6EoeJjqhzz6JwbW5RcjDkOC+YE8h5Giu14V
29N1RiQ0cqNUtWjOkpcXe3Avf8ZmG469mEQBJl36FCYJb+GsDbEQLnPtNQr6tEOYtctj8NEHcc2P
sdC+WJBdZ0deV8VPuDA+qrYgFxlKcoUi+tshlAyrz8AjF+nFhvhl5ybP+S5z95NYkiak9AsUqwr5
J6iFJxFW3bDnqkA7ceth3QFotbV9ms5UGy4No3OuFS5gEmxbq6tI4NsrkqgHFqLNO8QU+38nwxIF
q2iiEP0OQ4kJHKiivZll3YtomrRk8bhQtM42iBFrQHEEGXYdj1Y3FrN170WBxyopoIrlM5rUxkeG
bddcZjyBv3DRfdyGaKeV8C+TTa3DVs7YMg5VKyoluaRzME+sVmYw3M0JnEZesFSB/wOGFXSu9SSn
j9te011++TXTc7oRc6dGpbge3q/aNY3nd3RurUqqO7p+xrL2Xfpy5O75TChNZIisbpwjP6iWoF1E
TcOGUruiYts8ruKL/BfUNb4/J/XU0ys5soX9pQTadUeih7PcKUMbOuDxA9iwktNAqIsevJXmkJs7
SJN+aOfv0NR2hG2hx+WedqGL4ilkaoH4PznJKRfbq7ppx+dBZn4oMaNKU5tuULvQwHtBUcQWC2Zu
qNEEodHQLybmUM2dTY22BtftQIY7Ya7SAko2GCdhLYlvo08HA9935iuvp3+mtAlMjgdBBNprDGjK
YryXTsMWTxRl3Tmgbe7ZqslL8TevDk5VnrGL5UCZ6RxdEGD4XEZhx99ZQ2sK8wnWlvB0fHmkJ96l
nXXaGEIBchaIUiN+dtJzOVgLIjFuRQoHggR1AEfqf+1FzxN6q7voWJnUTQgZYERDgQtugEFluo/9
pqEcgEnJuYcs9xlwXnhf3/dOxs3qV5H52Qfh5oNoN+bwLej5p2D3lu0Aw0gJ/fEVakP4QMtWV0Nu
eYpIu5k9+BgyYiuBusfnPDZV6uThaf7SrjYXw2VKFX6aquXOhhfIehf0+U+VpMjYHW79gVLWfFHC
E/MRCAPCZgvO/1IP/LRp0Hs26ixQ22P2EgzjClMONeqFcq/n30GV5QAv/hbubAPZ9Ng9nq42WaMp
11OEnRgJ7G/u2kI7PERk3k2sC2VzdjEbBW8B/tvi3u0s9L6Aqtlr+tor5XD+BjwoX6kKcOD+iKnp
RawTSNqm1uvnlWmmKjnCqndZr6V42CRty+IWVnG4//yNOJE8p4VVDT8tnAdio725UqCLaJi7Kt6F
01OkczQQJsJBTxix6LNp41uANVlQ+SAJ0OgYywOGvCvCkdEqg1Xqp9/FdrNkYlSLFAEpAifYVYGj
QG2ZG+SMpwibH7fIo29/tkq+PZVK507IN0sajWgGnO+eugDDiS/r/1l5y4FNPRszSwTIZqG5wjKp
YiqbmyZjXB823FCCadWLwSweiWC7I7s5ouXFrp4YyCfkO5dsWzeo3HBSK1/Ie5xpBSjZ5YDLAzY7
RDsGR07R5RsguKZh1/zsPESEXq87g0HajBSGFmGeLxv3gIgrdL3BVAtBTDfQc1lqTaUt+QOkxjNz
j3oPMBqsz/D3s+UwkWvEWu10sQzbWuI83tidF9peYwD4XSMbZtfZ5gix+kK+AUGM++c1TL7qY3Km
+oUDHwxa6kYDObkNQYwdN6Da8J3aHL1JzIfzYbSnQ9UVyh9HiKgMhutjuWYdU+sUFjI4ZFQJsAHe
u2LKKQbHkhXe/3x2U2HHCTDFcU2PSYnpxSWfWXSlYop+R6Zsvm4U8QXsLNUCM3BuBWlMjQwt4MgQ
2LcjvuI4Ufv7njmJJGAgnWo2JnFbd9XMawEHnZsw2qGrh0v7AJOeyHEyeCFwu2+ZuuhtZL+PPTel
aRVKl0NT4Mu8WJPO/cgBlmFesjhqxQqjGjz34RP896lUcIXQnhVrELFUKYeBp0MmebE7n79YeUIk
dI3icHtPpsbbG2ywT/rxSmLs1AlMxtxLoVZaYx+d1bQdUcO7v/YkCuiv2RAKhOJRrlzSzc+UVc/J
cRcin9tSaeoYVLDuDXN+s5BKjpI4lRM7H41M5m5LOJzylEpWPkp3QJ2duxYxi3afoBFoIcxWyhh5
2j0fq1vvh5+vpxBRV8NV0LrWsXmkqetx1K63iQHjXvD/qvfRXiBqXkhTk2V2OYCxRe3K2KtOpZi+
WiTJnWeARoR+KSOFkPILoW9DGiJIAxRIvxeucgDbu+Lr644b66RakZmI1J26Aq8Ht9Uu4d2FP2B5
BJZc91MA+SewxBnvwfEDOrkU6G7qQ/skckTzxbieuzQG0TLUneuI2JKjbL1O+SzCueImdLl+mM3P
t6l3/I6oezjjOpizjI0yRFfgL1APzTHFcp065bF5vHgT+onKK1VDswNgaI7/jEM7HSEJcKSIBeuM
czckB0C3aFZd2tpfL+wIZTX9Fc6Wq5afbws3NcFAdbPlAnrxhUSw4RCjqddpnw2L7yspO34WAuPZ
P8sIDnG/LsAkPceHFWrl+ZIj07WGJ1D4hokYemCMQX+Gpa5dBrgMMUeUGIo0YGN/4eRhmLtUoLlt
64sP2oYo0j3TV8k4fnvdYbAmLE+2waodsE6nfH549C06knX8TXapjgYw3AN6w6UF+JTFJOtWEEcj
YSJFzDkkDUzsSoYMXCM7ZtIi+VQHBazBWK6pYNRYewL9vpjmHjvuC4jE39LWdGJmwmbp/lEDzNaI
c1WMI6RsZV9UZR40T0Qyi7o/CC4XkiMLmkL6c8bTjHWp5DBX9pV0nObAJDr22f5FW3uRis9s9aVW
tSaC7o1ZzRvw0ve/yKHhNS6Ik6dILN86myakRFsX1G6ID9rxPaXSWdNMRP92jm01SiAAs/eDscu4
ffm5UpmA3zIvsrWloUP+41/ClVmFM+Isap/kgh5PcgcwFOZ3LjygtuJGpQ4EZIg4zDo9zEfOs7Ps
QGz1dCHJWrNNfPpNktLbsEWTXojQ2ccckwuuj4EvkFJ7TBsMj2Z3Nihh5Wa3TQFHmeiePSTOLjik
80RRHut7828QZrVlKpAfmbKMrCLTckPNfG9uFeLy3fZI2FAdvs5ryOgBcB+qo3QI6shQEhBryup8
L2oRo3kULopnppUt0cd0HLlHjlH/37smu38Wb75f6uIO/sMqh/TvxXArq8oqAqlQ2ubjJ7Mss98s
PaHlHa5ib5jQ5JvivQg/YdovgNLApqDJCBNn3nApBDBe4K3VPrFPWE/gLZLMBC5uuDp+hocnBehE
3PHBYD8URTNxb/uvsB880mMFTdNRgX88zbb1Db4fDEvEMpbbNU5tYM07oY7W2KN3oaRDFqtlWdfw
WWjAupS6l4Nq8KQcAyWJruARTO9vLFWxJq9kVHra9LeZjGIdDk80AieVkyoWcNFIh4o8t0ru+5d6
S8h5RzB3UGOVKXrqPK3LozjF+mdmosj5XBfqc8S8N3aPbLKHQCj6mTlw+z5dPTDet2mKsYkNf9eU
g2ax3se4p84vNo+eQTeADZQ0pzfOhiE7nDk/U2SpIPbnysw/+A7sXTP5hTKPDqJJ4JK+UyftNNu0
dSs7RiBH3DufJgt727QOqoOjSp7FaJKEx+i8J1pQog6lBZIQ1YXsKUE3HRL73IJCUdEn0H+NDt4n
7QAD/pxddhubrmU6/leukcfMSTZ9VjqkP/5+xddiydngtZ/hUe5PN+/0gh2kGcUuuEWG/S+9zCR2
eUh9lFne4x3KIiyaGEv2Ld7FkjtaieXlxCWf/zkIt6tk4k+ma7+XElMnm5CfFsWTdXJCtItkjq32
AGvhPn6dmMc9XHLiZnlHxvA/yF1mXYg/AVGVV8SbgsWmLLZmkj7j9F81nzQAoSdO7bLT51XkkI2h
eGryoN+UCDF/ydjCeUSk5FIBVJ+/VRLL+p2mXeBt23rufxy3kuh/pY9sYw0X7Ixrq/jj5pnA6YlF
9pxJ0ut84iIFFj1cDbD/cFf96yhxrh8Z8MGsSHJLWh2W6PJtU5eIuE4d19DHcbewOI1+O8jp0am8
aRhLa7bg/rncUqTNpz7bcaw4UcT68WsPeuIILVmeGCLulGvShmp5zS6cwH8i5uCwsDWi4AZqE6XJ
nHe0sGy4syfkwf7Wo0ZboEgrLVUCUIdDNwjEhRaOhrTG5WPSYR72EJK2L9MS+ZfMlxfAucrTQsPE
Mj4nc2qT46j7/8m3Qyw+U9NQLSbgugZGUrL1cO5Eji+Gpn3wI8cljHeM1N18GzQ40G9sHD7GtZLB
eZjwoK3lRrVDtfQ8pkfUcPkMJIv/nPv1T42DwUjCm2Dn2/phS0JDgB89T34M355rRsih4Gob8P5o
Aedsc0d2aN8I10UC4UB18BwlWeHhiOSGP1TwOoR2rDgNQBfnwuADWagw1YwG0eZhWXV7wSbCfujU
G1TABrk1ZIVs3ix6cx4my3rWppuJ0Je/aAIq1AvDALWDA5WhHhnGMNgl/IM9i7B1zruw1ZmWEcdh
QvfDIaQ3JipLlPWMreq09WjvHy5MEaf3gFXz0ISw8LScA0WBBur3E6Tnk7WxNxaIRT8wqCkvfjpv
+2lB305JoRFdoYBUz4kXlrckfzlQkD3mjpQctt58RPmLmWFIQld6WvKBY1MBkrLthCdHBfp55JkC
QYdBdvEJzLCuV1n25SRpFEE42NoHrqr4hScned1ShzMg05T+hK8T+CCDapbpl5EmPKtqQ2aFVFAu
tr+MNC30vPuhJJn5BoTTtpYwywpPiVgVWvp1ugP1zjUbDSvvaW10vsz0MApDZfS4Qf+sCaDSWWB7
jk4sWDdPWcGREVWt19+wskS5NxSAbxKim70tY22RMyx7gCkF5Y0KODWUg7me6zm994DoTbZCT/I7
5FcTBG9YpVbnMFqtxOD6bHIWXXkiiNUtBK2QRmTD8tTeA700oqQD7mezixLIC5FpS2qqcbhfu39e
KuXjlANI4PxuvbyUXAs0C/asLvj2ZS+9jFMFLCjtjsDzoOerxlrUjT/ZMq3K/EaS0w/B/9DEGAFq
aWw1vULzCH53vnoPZ4aEyBDJFqQPQPGXUB3xjaPcd24UQXqHrqYExTn85nCqSqy/7G/LhXx78gDW
gux4JuewNjoaplB/UBW76MwitA9JBFJjUu3F2YXZscJgQ35Q8ZsMZG4cxTld63rmecFvOGfK9Sop
A788sHlIIv2ervCVifj4sygNhQ2utebzIYBdL36n82KOn6ytzzx+NxByMC9RoTz22jwTRVzS/NE9
e7Rvrv5GMmwIXCBvURD110ZCWvogIyCPrCTTOzDlj+x7PEvtpwQzREqU5EBb2dfPeElb2BkNDxmB
JZY9cYz5WaM9CmJCHSPtW5ArYQ00BiLAHzAI5vkTKEqQ4l5zc4xFBTkTxloWnT7FplrpLv/G86+L
h5YLqkCf6R5YVhpWoMgV1Q/RjeGcu09PumkvD4VjM7K/WbxhWkx/BkMvmOhUirkYfO7wtvKMUmU3
28QFC59wGAS4o5dfxGPlAgYSDG34Qzwo44HW+gZtIQ0G1zj3N9B5D02lapLzmGOV/Y/7F/qhQmoL
3bmRzncr9V/f0kstaChRrRmFQpFqHAinJETR6a4Tu6FUy0StV21QQwRdmHP/r7A8nxF0E/JrvG3r
JJzpeiHZ+t0H+/nSDnloJKVeDv71fSeh1PONtUpueUYJwUT9njfhunQ0AdMw9UCVMpqWGyrhRjfo
b6PUGUzcDjtO7BmwtvlPSpst+LISXRy3P47qqhquLh90Ipn+neJI+LA0Id5pc4UELEFn/N0yK/oO
SOFVAWvE2sSrcjwX5GlZFgHo2ZqYhoYNJdT0DQ0daUGCvyrFroOF9e+W7mgqh+w1vgkkxdB51ekB
vkhoDa5lE9ZMc27F/aUJClv0xc2YGUVrvYLTn0jcLg6PqgH72wRAax6jZnB6/4uoy6MX1H/oBx1/
sOMkoFiwE1QxqocwgWM7iOG+W3DoKPzox58pZDWKCm3ssHBEIo/+hXEzndIoOmS8NJF9SJ4tKvqz
yK8nWDDeqfJHcxq0syiEq42TMYwr0u8fhvzbspZXiS5mFssOlGyLqqau5dcsniAwPLOi0raeabv0
iaoDpzzUwO2hYTxcqZU2pOveIjfWN/gFh0YK/JDDAsO546+wECuVaSr9qO6sBCFx3QzUVuCR3weZ
TVyIX6zjExk6zg0AVSoswBTBuZfn3CKZydFcaRZsS/iJOEtot8z3v6v1aLVA+57gho7Gh+OIY0wg
fL4zyx7x1wbIs3k+dGR89jvAxNKXgBWM9a8CQ4sIkp1UJ2U6nfzFie2AZj1UCvRNrIbXEJ8Bszpd
D7oUB7IueuT8iH+O1kH8y++zF1enx/oFDyjHsR7towdMFjSZL57duJfGYWqoExEhtv364GEVGhCF
pznVHd1LlKzNPFiFa1FZM8KeDlq5GhkJksYyFDgk7ydCXjn/zk36dEFkW7bjjTQlSAhB/YRute9p
bkDL8o4p4oEN/aKKwwGvYQ5cOjwsauxjbX+yfH0g/5JinpB1hFyVBwJQGq0XqeCLWMtMvyZCZxc2
7thwy+OaaMDAAsbWCpg7syaP9B7q8GWRVA2spnL1LjpVgRp1mv7arN5mVH7DVhOOwSfFtDNbVq++
E3bIuyY3fAA/mANVcOjbuu8jdce70MsI7GmVCjdtrTpe6pHzHPUAWaHBE7jxI2HlnEPyN1IhnEuq
82//0284RClsC7BBAUXA4hVFke1Rg7oKQy8pcRcsbyBPvQQ6ulidRDV9qGSefJ6YGHFjf7TS7KH0
z1BV6A2s2egm6iBhtEd2vX84x/0WBsIpRjDzG5p5+52nt1lcEZFDV2Z/1FwrpOCCOqbd+FC+t9g/
3d+J3EfqZmCmMnqQKeSObH/zHq+LPFLoykTGiAw+lJTG/Exy8/+xj/qhE0dPizQwUqCR5XznpHRD
Wm9oEi0Q/SGQPZFLmLYL++2PXyEZ6ECssHHzx7GC50Qm1JimxX269yAAVIMsQ2B8GxSeChou7Ewg
RPGEB7ZPnEdHpM+xv3jpaeXkTZn5o9ddwcdnsfGf/9F5fq4octFOTL68PIDng/soCkjFbkiYxQ7P
3mvXD1hZ5m9UnvWVpksoK7R6+lyOVtx8OcADh7O39ix+jXS0U3Npd1x+cOjx5bV0I+7mRQs+rfiv
2GbyB6AyAP3qRcpy7M5h8oUjCBXxNoEmesmwYbT2hvEXLF9wVgEitzgHRwp7YQ6WyEWsuR/pu2Qm
UlVHpQt1ohsw6g28Nlpse/zD8VZ8XIBmwJPrUwW/f4+oE7ZQBDZDYgExMKZzBnh7FhOZzrFAaNPC
o1//W9CKAJzkrifAYTElEoBZY87IQBA+lDcoIeBARXj2uJUIRW6SmQTNnvLiJOXAbcg9NjJ3SP84
C995nBxlOmSDU/0wSk5H4akmkppaPPR6durrM3fZWIyOJgaXGzxIaWluMpN0Fbp5D9ilbDcQtxYH
l9wzHwdThrfDkbirDluBVvn3dT30VSTbqWTYjvlXF/ro4fE8yyX3aqZo+LeNHuqd4XYHAGz5mwCh
3ZprWoByDH6VWPA14IdYrj/V49KaAPHzRUfRSZGQtUAn5ATAOVPeMVqpYkFqNSa9XXUoYCq1ne0O
zJIIf2pOMFHMCSBXXwRNtyFwgfFTMsC47POo4Pgsi2AvkJSLoat0ptYN13BJiqQtNVuRTXJI6L15
k8d/oWbXKQMxBBZpi80S7iEF1eYd8D/6LkcXq/+K316p8xZCmPc5wkqTheZwwHGKiC64KUhsVIre
XExJ8EuMwfEjyQttqetidlqoEWr5kRKi/BaMONIm9ftEgaA3g/NmYpgHTrLiyEzRrdHtB3nO4ugC
t3lxeSIxzFawlP3ho2lWQZSux9oNWjUhr8VM+aL5ptLSmUwOJUyfXq5JZ7+YTXsY2IHqbvoc0Vau
9FjCovLCoFtaWs+daj/TTwlqmCypy2b8ag41uHCHYCeaPmtsfHNZKEQp2bByZUSjMqRGgEaHgFtu
6OawXhPhUDK43dbaDN8TO+FxuClDJDc21Z0+3Xrv9iFMjNWNfH9cfRtP9Q33GoIawAZN/HLnNvuN
2xuQGfJccudKOPoXoFTmhjYoGSmruqHCvYWBn4pvY0YTGxTkKYEXRM1NJ4X5jbLfryDRVAjgbyTI
LyNWx3hIc0C5NPn/C45aIIo9TAzsss79rhBQjYl/Yo46pHvzlTJt4Q/L10qm000vXf9jMwe9NWsM
5/Elz7aOzsvqBTBDTNahLhNSM3NHTHmMWofa8+gjgbZQM5qtA8hbtBOjgFtbIbv8TgAih8jIeQtM
pM1b2OuIlTxVs0Ps39zZQET+YjaR7dOs1fZCikmC0N3xxU805nAdtUW9+4vAa9iHdMbSDsexr1sw
G4GkFzL391C6lW992W8me31kJtEBBeY9Dljnz3020qgc8QkhrCR2sYWrOdBMyLXEzlr4BSHkdg78
G/io5P8edPIJCIcnZKbYzlF+KtHXdDdHXFnm+TvEFLYrSGcI5wr2VTTM2pkIavl4INAk38OYfHlh
9/YgmMn5AmNgBynetiyHtE84P1ncOIC7TIPLVtd1Bm3sO5UKGFd5MWHq4LGBNwGSeanvReAFXGCN
TS9i/U5Y3X23qgButle0BGqS+n1Pncgw8KCpvSdCEEGtiogSVPjKtxkT/ip/MDfxX693BSdkLFK/
zh40Sg+WAX7Odhve5Z9FFoJXGScRGq2sNDlwOb0J55vlwjzeRPT+oI9sOZHb6mP1zJpoLldxHO4s
Sy79WrgQ/zPJx6DDM12BuWOjzF/+aormJSXzJprDhUaYyoGs64SmiPMHs1Mgh44h8RiibqUSpIsI
75rPdwQ2G4r6Xcq+Oiy8+En7xN5M/XIGlFIXQ22iu116fbe+iKSu5FNxd5ioAjA6SQlsFFTc1llc
wRxmiMdXoXICPKGYSjRGbu/X/7Cf0vOM+DgkUH4+n45vh6iKc3yzQIaKLdKIQLw2Yl5wjpC7c6fr
6Uu2qYNDMEFupJ5jcsFXvvnyZIOaYDnLsQM0WKYOqfg1CjlrpPCV80Bm9yNB30qnBxaj3ugROXet
jyRNdQiK+r2VHczhF3YTdqYI4t4gdAPA5EITcaRncL7w3X7YfGzJ/TRhT3ovd/eYSBUVvTkvGGvn
8frDn+vaqW/Vchlj7fnyLiGkjImPBlet7sCuMe7rmQAW5wwilirrKIpWiKJWL6ipkZYjRrMq6sl9
c9gdvJBgtTIW+IHSF7eWSWeJr19D/BdutCPTcQibVrvsgOUqeePgXFMsrUtsv8T0s7LpGid34G/H
JMbpupz0TWE4Kx3x2A5/5egKVhOSpC930SGRoTd9Rb8uYQTn5G9iT2HUMlkOsagFoIXOkeVHbiqi
A4uY6bT9MDVlU3A2625mh9MnzNyXuhF9wYZHjBhf2BarR0nY4Yh2X07iVMD/0+SyJre7C9wsWmSc
fFIEE7mCzpdhW7oc5TqT7Hub3G1T53xRbm8+CoC/7jRD23r6zd4OooywvkbN+kBuc/nzpEwU0Odr
0l0kESXYfQ3dJ0oDmwD8B3DCXKMIvLZQli1Z1ogV9PaI1BFa8pnR8JuwzrUYYqjqcNcXvGPJsx7E
KBt4Qkekcn5Glr+wnweSdJVSQKP6tazjysylhAtV1/BhL+7SAnwNnK8sYuEvO0sTI6QSZDgoVCn2
44DkTo39qeYgJDrBkXoxPWZDD2chD3SfQhdZdB3bHNEDY5JP7+Vx2UOD3thBqhGun/TfU/oBQDy2
vmIUQSQ6Reg4Raj6U5sWt/PI6wHjsUFubkyDOj3wD8e49Nwotgc5s0r70D0LSP2BTFPdaU9FoNxi
SEv291RfUXl3qrnq6AF4MGSmSkT4W17PmC+D70KqWcrMweOYIvAx7d9ftwCGVlaKYVBzcCeNc3cm
LkFZJMoccz/LZpM7PqpOUJeHdl4YsKRXmt8K3hoR77mxCxXwMhk8o3HhqTfuwRBtpf8Sgh+qqRLR
BozQN18AbVuTiKcEdIZ51nnjGpgPx6tciTvZHNhL2fONaS36OePIQuOl8Ph2DrNxD7b+fM5/fRvA
PjACuECjuI9eEq1fRPgHZu1V/KhgUILWERDqHolSgs7SNvUr4oL7j+bxOzQfm+ocNIQ200FWB0KO
lDLF0/ywoRBlrrvYxK0St5GvTSU/ZfufxbXUvddMQWHX0rk0OPckRNwlVtE2dmNJmQKNgqQO7bCS
wN5jrNRzutvOw+W1tuT6JHrVi+Ih/Mg4vnjvo4Rc2MiEm8kWni+lsk73LjtntibJR42VYQ4flZaI
7dmVGqvMGoyTGSiomfol31WBP+br4UcgkZyTsUFHXbcVK34jIH7YAsRrweC7C4i+2Zk8eDVfr+D0
2XvGXtMaE9SzjSkgDVPTmPRcCBSLKtKIcwymCit7p/Ruw3L754AiB4sKe+IRy1zxnKzdT3sqCcrr
C3YF1hVvtBhImQhf4bTqGELWA+vasEwzw5424j98p4dLGcpFBiVj+MifSefLm+qYS5dZ9Fnox6nW
Viurvv+X8FTyXHSO7EX4JUkvLxYUavFlmFB52dZCUK1eWaJbSr5KQJtbaZB+spJt5lEpbfeok72Z
dDKopDjkwUmnEBzhwt+/T9iPXlZlhuL+5o14nES2UFpnn9AElRcBQxqlj+9CBAmWbr6ifHjVmmRy
PVvkT64xE0qaORQKfFdMJLZMV308fGlH8+BfJg93NhzKZ4lqU8sHaK4+nOwkEmWpMBeyN5rlRFVd
hwQixOZuVUKS+GufZCLXs1ouwh07OvALgqAo4ixJrSCsnzxQSMfa1yIOo4BaZj52jKfpBxXiyEZF
0zmbL1n728D3VbWO3zt8WNNYo1IEP7qhxF4mOrPcaBVymZUZyuAo9NDr2tcnHQr8a4eH1KLU3FJy
vBedRqYq6Fj/l7bDGyCc6Yh4iWGe6hZOhcTLrWYGxYe2/0SN1RE1+z9+BO7riyquUFjXCfysgKf+
AbMDUGDXot3wzD9fLLmWL5mmhkic+ecG2VeoWSohNCd37c4weO+rvYkocNbpXsQD4CYFP4WaQMMQ
vCRp7NeXJ8FI7aYLmqZ+bDPBzCj9QYXG1kI+SddNL+balAbpgINYhwneV3BQCW0sFemyJez9Na67
tRWcPg2V6crmLxa16K7BbKAPBZrcaBMSGlWnevLH0hGNNYwM5GBPKNQygqakEHK+Bae7Tjv9/klp
I7/tPe1AVkUHPLfhVUUzYbdjaNYi50TQ5X4nyUsCqFgbQY9nlEIlBpeUEC1NuzWsWeP8P4rj0bst
7IGCLAkO9erNQ4vt0yLohZgAKZx0a8c+dsdVXkmOcr/S86ZBl5PJJ21oeu+TSipY7quP/XcrMqpB
P+ubBMLKgdRH+/0cJkl0HUpibWqHNWQB5gMjQHvcEocfP168UuMctYDdok2VH7Zd+5FsyqUVc/Vw
7UqrEvz0DO5RX7mQyirpOMTCjHLADByLorJGQO674lyd2cFzg3VdJOxh2AmnlNKjFsZVoAF5mlz5
7rRALXDE96wV8u77HH5yZ9Xu5t9tfziq9H+CUN/4OCtcrujdA7U/bjCLmXsxtWNfXKbVaQqNrMjx
179t9vN2E/xkQabhE/Hku7UoJIjYap9A3j8I/AfTUuhFakJ/fntJsHLUBLPOC0RyocPWtTkvP1Tj
h46A7w6c3fZWPhMk/DTArBGL6FpxCcs0KHBPLY9Vl5r/NVhdBXPqZC32TX0Wxm9WKhh6hCS42+IM
yWHQ94AXiUydf9sa6lT1bRxv23pvOdzZNUODu8oFcMIkqPXEsLWLdbwaVn0rA3cz4mKEBQhr9F2p
LW7+2us50iJd0d/9tmuUk5fa3MQDQdxKUqHBjoNXXwliEihVwofWPdbyursV70lL3U4Eo1mAfipa
uTzitmnXqpawVRcqCMNvmTAIjgGSwqgpFluEtvbHJtCFox6B8ilyCZlenZyVNCVOi1BftR84oE5g
pvhqinHETFclWozz7xOEt+2RHPVaTuCrugaMAm08k0SV+iPSGRnOdIvF0DznQ2ndm11INZKuxMd3
mP/Rozk0wUad05/GKCrwfmNt5V1nwEWoF3v4FNtOBHGsFEtCNsu7AZZL78yDz3Vh/eOgaQ+9zhwg
M1Zrxejq6d6Soi268PlpOJ5cPgku09v2hdBFZbHY0U8xlUz46121Pp5Ln7vr/gPzlcm9qKIwWGSx
QHyU/TMC7+WoRzV0G13gCXL6E1Dr5ioZnDey7UcJGxEXFDaTWP5WEtndrYuAvgxDGA0/QgbFYhWb
kmZRy+mdfrHozOCJmncAsEVNvNGpgKRLmNXc/NSqp7vnhHm4tH49koar5FCm4BMaIpYpd/GOUPzG
MUERoSb5GmiyaOYUGEtJGnp+AwcT1BhmsTT02IPpxJAdGLmQxrYuejesT1LEjw4R+LAfAP0z02Ek
o8t027YFiYFeA6A3FK/i/Wc/S5r8U6Ap24OOgfpKuh2d1DQxWCN9vSbpTGkt9WcI1qbqlJ0DJtD3
A3dY7u8ociwyCs3WOGVC5OLrTjV1okuqcr4gXzHAoyyFdjy0XaOuou8jO7gZiCXmsu4A9CV51tGH
dlN9pImB8jO0+MLI2ECKU0DW+5FbJruFODCMxtoE1rb39CEV4ueBG6MH/DeWBQHr2Aj7MnNkW4iX
DjRLfwSkGZgzThuIYi+4zc9W3FEB6J1MKxuAxStIPeNDyGc01YCFf7pia027BtCP/lxu9350N4eN
sy6DuxdAEa0vjBnwSj3briTaeSmjdC2TAQHrdPKEZsYA+rNe1rmaO5Pug2UucZLec1i7XSRU25Wp
Oy3bfb4hvbu+k6h7G/xfDyzTiobiTBraMP71xeAkX+m9NMw3mFTSNFzbzrcaU1UdCzlsIG47FkWD
ZGNFFir+C7cUZ0rV6HZGKTVVEMr/Z16TAKOYleDqMxVxknG/j77d0+ISh1F24qszadxQPX6vo6Ro
hsjsWYxotI5SYeMvaHh5L7NBwU9bnjsHh19AeNQ+osgDs2VEh9VnU+i1KUfobkKgR7Un54fmXTj4
51kPCtqrTH/mvcAcl6XUS6cgEYEr2Ju1JsHI5pDL4eN9e0K3d/BjRUhBSdBnSN9p6jTJjKdye9LE
x5ENkczIStItO4UQrIwqkUCjnUOcAlr0vIMV6nrQH2+k19nz0ZdL2EVignQxZtkv7Gm2TKkuHpGX
PTiyBmYab2qt+mYEVISyiJLow6JWAV1ER2YFf+Rjb4tXFMIRs7wvqOhV+Rxr5NEaB2n5k+XgvqiF
VZYOYEFOZXkE+XKNqWSHLLlfes/2wdnvttZNecWIPwUyptHb23ph1V3ZShKZAqBSMzT84H/ZnxnT
ZFpCxtKjQUMvqcV7S2EjOy/1KD5Md/9WpL/5t29KfJrkM8jlbQuLpvn6Lscus3o3gCg73BPsMUR7
rmo9noXxHb900w3mpYf1fG2wvUh2J1oj0uJUpXKvGUAGx1u+nQVlVbagITs6XpCY52p6kqGsd7xW
eAoawsYtzi5rIcapSpBdvnzqGXxWfrgE+a5gpap+sS+HUwYzLi+JAeImFedmP7J+pbrsqYBbvBkE
84BAmxh50ZQKAtjnVr9Mj85msRLXjewPrLSM9WVC8zfsq1sedP/X+vNgIeqFJNFaNo6bYPMDfmxl
BH1fMiyM8LoVfwWGy5YTbC+vwz8L5XD4VrxMs9c+z5BG7qAWHA42Ev5LysKPethQE6vxmIZSDFTk
2TD/2a5cgMG3oosp9ivqXjZZjsVbDS6nQwf2nyw9c7N0p6Qgk96JYWz0GMdlxOpwKDTgAl8euH1I
d605AoTL7Fl3whFe9PGUFSKiFsM/yPlLC95sqdMMJhKbwuKuVN9YQl2jZ4yIrL5IndXREXjmKkht
yRoqsCcEQkVA6mK3CIW+MsRVvXpiM16W4p86T9xBk8epHkwuJQz9CeOSUCRur4FB6+gNTQIx9XEz
y4nZGyU439oY0d8YjUGCeKRlcJTmL/OyfWCJVGbqfhR0fQqjvR3hEOiWS1vFOC6c+1zWlKUVzW8Q
jHCgLNdtem0u6xbJIwZJ5lUhuY2Oo6RVAWwqWpoeTfl7P7qczn4JwE/4rn7ar1J2vTX2YL+dG0i5
VhANR8eSHpoLVghdIj3rg81RqE6EqCUwJSNPafwBLhXGCFN1yEPnR6jHV+9fmZqkfaAjg7SOVhc7
HJKUzQUSqCeCyST7AOjL5YuE6DKmKKZxZN8gnX4P96VMWtBpCEGejAlLStYl3qbicm7dGnxrAcZn
GI/fEgdQScdkY6ftsdXGE558QxaLyU5rhW2AUSZ0IdfdXelwVHCLq53NRqz2+tukUdQ5kuCUK/s5
HqA68mtFYcAvpVCAxM/fy/ce8iXZfxEwhwi1dpzGAil7zckAu1fCsQN2x94uT2+xUMYqUDTYo47C
G/i6vGa9JuEDE/6wQoq4TBiQXoYPzsYPxcUuuae/r9mkHEZ7xb5yMN9xeOuCGNY/8PORXkEJc1y7
v7oRmJ1mBhgXQsa+xrDub88128QtApoXSx+iI6X9LFtZvoMHtw/02n7dsXfW4aY306Z3xHiaZDSN
vxG+gYt3wgBT6ILANty5K0rNvZsNqC2Dsn8QeJs4PboPj06DZqIdROb057B2vbrfG8dbA3mw1uSa
gEN9gmEEhUIddZKtxx9awj44cXisxM3ttUN/8mP1UgJRV6ZKAfdLDpHLT2hlzhEJMiG9SHhRgcEx
dUCcNCHzYLN2wxaBXe+bhWRSG7jQ+iTJBWOzWEUts/N0hFSTiTpeA5WPfSK2MZmamnJHk8w2tAHt
VKFQ+WOY62QFRXji8q+C1Mjf5cQvsWKQiHKURzwOIWyBf/ye51rwYuW9kC7E+ZJ2NFrlyZMkY/zr
h3E7gct4djtx2DZWKEjXkpdAypgXS3Z1QaiKqQBLYjc92I7Lobgkaq09ES/CUApZQ2JYSWHa2AUL
BeeUMWRWtwHOtC9TbTrW5Erj0BQ7QirMjeKrJzrqHv4WGgJwC8h5bCNekoy4/2l5L215uqiqA1X7
FqZTRF7KlH4Yies8P9W2S2rFMINgrqKyE6nVDSK2sAdT6Cgb1G7A4SUwaJsote2eDNdRWbIissYG
JwTkMctI7dxOswgh5nlu2ZRMfnf52LTifEJNaZCsE4LpMgRPm6GSTRp9PAtaknK/NNb6skba4xV9
ZO4yTGJ60koDBgh25UDeafKIoidHyW9qDa8JDtXLoidiAkhR09dspiELLaLVmZ5ljf4fKbGlFFIJ
AdWUdtiHoM4UlSI1A6rd5xb51ORnKorPmqMfNTAtht7ZM6h1WD1qviLuQTJMgkcMzoLBFqSTgZwE
gqyXrs6FI5yKpUo/IAyFEame1bEojRbjHtm62Q/ZevgTp6DiD1KPbSAE0va7tHcVgxczAGpHzz+X
pQaWoCBYZ5MNgchx5XRHdyniFcCJN+zXfkVtxHYy5EJQUo6z0VsJpG5ez06MCRuvW1wHQwaOKgsu
MifWu5/wVCgzW1Br4bhp/GtbXGWN9w+2GUV4uCKfPvco6Vc0IZIXZKeoEkLLtEJ0n/XH7YOGB+nu
/Kxv5xqMKfJem/rqTCP8MacyZReu1trrxolb0Lg2ntKTuSrXTETr3+xwFk64LTxJraDWqD9EmOH5
0ak0gd7fuDjUkKcMkY+653IrJDZp1xncUu46Qf3Yn7paLtgs2RdkneJWIYhVGtRjwztAaDbZmCmi
cZPdI/OMX6q9/9Nvtwd3bo2y9W1MBA9iIHP0DE7wT8dB2szIOmbimOJ5PNcIFO1cNBvSnOAQ2gSF
VZoAVKkq5S2emeWjnownXXrsvTss4ogpra9DZQwj/Lr+QX/b/Wkefn2yuLDPCsesVwOptMWacbCv
yUEGrSNP2j6gXeTyDasobVOaMU97y8JZ2dF8V9HmAgVPap6UiclYYQxiTnA/AM1CMedo5UcyqUHt
aHc+/MlwVpra2GUWbhBjQazsRhxnOWhH5DEBPfSSv+CJHbrhrKWzg1D4P7YSmc0tobtV95DYwI+M
mcFUz9V9sm+pgAqTEuMdOa3XMdfVOgzJp7/snQeuVTU8jWcB/3C/glqBHtiTqh3azzl4wbroA9wN
dY3PO19V8WEz8FC86J/69080+hBupnMymxLuLj2XLp9MfTzct/BAS9JvpLVH6ITvJpwTWq/Zq1GM
AdwU5EOOsb7w1FjrxNBzljXtlW26Am/+YjOKfFs2ah5aZ3e5J//NpiaBmK/dGMkAcSDrAPd3IHaY
ZtE/VT2w2exZ/LnPjYCR/7SmHmMaKqvpVKG1iZxK+abeiQbrgqqtZJ21F2gCEkUoJC6taoHAq97e
AYow52pEJ6DAwrJDzPiXggj0qsQ8YWQvDRrwi3BUD/rv54h/1o17PSDWt+zKPbrMLbZCs8gmQDvX
n87lzqHwUKhRrM1ICX5WmTuZPTUBslx3OfIcFIZjeJgXC41prPTK2Rn6VOYo64EjkvgWfbZ0NopL
KzWHqz6GXA2RlHMVzoQcHBBpiw0k4mf6vw5Efuy6nOf9H+Bszj9/VawPK7p7nKuxPf3ienD44bwD
BOZDCPUgwPuWmF1sNu0SLJdQag0OnaxbATtFAoj0aSXdZ7ajb9puEBIMzUCVypZOU3BM67unsNWG
4dPmiSKvy1IMqnH4LPC6M+jdwQD8DgEXKTj+SJnIqIQIceDlPaKWi3MLRoxGtC1eMPdNbVv2BBW9
6qzaeASMmpySK+h2xDRzDhJ4osXGTMXuKsCWowXBTSNtsSkw0NKIXHXfjyybZRPcO5fSEl4Gl2br
yU/fJn0iHlMqhNszUDf4LNfMCoErkyumpOjdMI2o0tPkeKxTan+LzjKvlr8QTkMMXTjGx05WlHfc
3At451iVPbMyBV3xNMrFIVPzSBRhce6ySkaiCopOkIzAy9t1ceXe9MBCv+KSSuwb93LJXG6gZA+G
p/TDQL04EaZb6hgsiRtzophWg+qFGo++2C/LTnRRWfpkg5xDjW5WXqjlUESNB6cPbSSsOfGS3lja
if/i4OI/trN6/1NjxAln2pe3lvVBMSXFymCVRtuTmSQvd3vWUVJBzmvNv09NMzqVQmEjoNObVAKA
b332YBKruA7tKElN5SN3Ka+Oe98L5NFBO2kYoNGbriFfnPwsZF+qxN8TD9PDWByAgEGbyWlN9S2F
XBJdJw7VmfeuLqOWPoq7erjZyQA8i3tBNvbKkit6Eo5/XoROXBf+BSZBOiYcpwPfuFU6lzpu4/OZ
kxAbgekvI2ColPa/5K2n1qJ39igrBpsr/hq4y6dIV8dL2QNySxtYJybhSOysOyG7gM+GcbQsqH7c
33qvezzLQdHOXpwIHebZyuR94ZQGIwd0IB1YCFujVPwP032Hpz4GQouVypXlwRIMzSiokZkQktL8
AsiyekYY63a0NyufT5hbT1Nr1lC2wPurxAiEwtPm1e/Ay+xWUjioARbzItjSbo8ZrKvNqK7WNQ9o
xBfLOA81g+GxLmTC+ow3OWGIUOgE2/mkQU26DyHZPAwiL95DcheiA8Kn95BPbrGQHNt30t28QGaT
v1d1bMHPdsqKXTkedxoyUYdvHVyU6fDgdtSf7WMU4ibS8d/5/k5aPXJwxR6Bm9ziNzr6fShbufjD
arnQCofOZdQAthW5KBOz5Atzp/VOegK6xLWs+XgFuq6j+8HRlif8Sbsa0CGZDHKIbAh9RRjEXYmk
8xDr1JAFRicoS9g8oKtdILJ8KyzxR/g8L/GSSDTKZXhxTJB4G9aLMw32/752RpR3sH+66V7lL1Nt
M8DyOckp01SgDJKT/eD2fsscoDA0LHRpkfZGu6mbzWmU5llpEHrMLQQ9cyDVNI+wnLZchSeP0VQs
ZrIfd9knGaW4OFGD9y0leLGyC9nEaLTuOrorUxXLWUTrA6uJnVn7Ikxz4p4YelwflP0tqCnzK+6f
7EvfaxDhmTvpXi+G+sn1G4QsHpsNUApYe5WOtyuTNuSBDpVGIqMkeczI43z7RmpCh2sk3bELh4ZV
KpeXWheveFhwOTALFsc75jyutezm2HtH87yjwuFLF3RB9u4aR3p3it0cfEjRscqQ5otWdWJtzFrb
8WhCuhO0lNIFJ2A2BpHbkCKnro9KalWVvrNO8T9eTs2eu06J9Y8w5EWjpAITUpN+oH0LwhoyGyAZ
H/NskTZfBsKeuu+32MsMlPAftNL+u1r6XJTPHFz7Uo1+V4q035C2+UUSYZbz/SN7wt5za/JeX2rj
892hKjWn4k2fDChOhuKDuhpebTPAC+RTohrh+eX+5OuK21RiSDzTmhhZCjRw2nJ2SWFiyJuCKofd
1aHaixGMPisjN1XkW1vq+oTlWyClIeTH+QPivgcCqVR2LlKoaNchB5YMWWn1LY30+YfNuCBitxOr
KJHSXHwdGhsaaVNOnPN3CpiMK5oGV0qTUlU2z3j8yp9+ljZPrb6BfMmDKgSIWL0pJgArZdT9VdCa
bX0aTXwQU6q+4/cF0uW4PCrsUO+JXwQPmvFRcypmtczrCSBPMjO0x4d+1+2mGcGlnPbTIrJYxA7E
zS9SkAuMNPr/9SPztdygxiOBCAh3lokIDjhcLPWxOWq7JNWZzQ0FoBett+P6nTgWJe5gv8GLtsvV
DpDHOlihmSiZ0u23v7CkTXadJBU99R7YnlQ1WFeArYehGJ00NGdKd/NQjW+zYlK0F0oryk5RGCHZ
+MYjrNWEJL0uqcwJCxC8HrUOffg3iEJitTK6zfQVEW7SvmZYZ1eod4AUPQuw5XCmz/qMJrYPuhC0
zl+JnDPsoB+//HgUI/x/Ib2YcFANIVdcvOmC80aWdwsZVTy6khWEj+Qitljog7prtD23Z27oFpo0
bmmgVgJTUmJrxevUgzejCx2LvPzP/Bry/G7lTlIpAFwMHi9Hmwr3CLL0bFdIIRO67PpWOTcu1hBi
IJa02tOO6bEebMcLX38BqgmJUaScAZLOYmfOs0dAVzky2EJyuPcTVIDgvpKmqs96ygAz+q9BcRQg
ef2g1Rq2Qv6UOOyEOkrkZXZFvvfQrGtto7WvbtcPIflwx1ASX7BuY4lKm1nHYOAtNKvfEYMDmEa3
PbnT1I1f1DybGVjpdGfzMS8c5XjsWBQj3PX5Ij2Lxvs68XrOEpvsgOPobGyQjMmQ/KjmOZnsZxDg
BS+zEePbxfjgISNxNIM6djOx0D3XCqw7xOqGOVjtl+shYNd0lFpbcdYyUSvNEu/mu+WndmKqS5l6
83VaaDhcaIsM6ry4FN1J1y1I89uRnzpCCOHsxVxODBCjwtXcxQsBL+LbZv30dj75knlKaP+hkZ+Y
Po6kfXWrN3jF1kytS4LQMuPCahoW9DM2N+EEuVrfuDDSfbHZEQWxRJ24ALODxngI2hIdxVFgtiiM
J1xMnqlqaqivDnVtaC+a/2EL0atRYhaYXEAh8FxDf6ylbMHJ5r515vGWQq/PoLAQWBUbFfT/wz27
XV7kgSwh3TNwLicTSYSi0vCCeat4B+zmWYyn5JMDwsWuRPjSkVT+AS9Etv3D7izVGxg7+v12RRgC
Pm6co/pDUeobDfaiPR2s/oB3KGDfE4knfQr0uTQZeJFfec61oFPC8OVBimQgH7n6bwilSfA2W9XH
cXbIent7jPP3D/fjKSHr6W8QhL808I9XrtEwBbFZ+1C6wwuolRaU5QxeCADI7HZsEiYnNLrNJMVN
H35FoKxsCe91lVwHfCXHUBgGvVZipPU2GK43hnzvaubQY0TTYC1WTeADQahpT8NrVIVsKre0x7rv
W8YIpWz936lBrjvKxd9B8iMG/KoXp3Uk68zDwrurH5C+Lryyr/pHbyVp7ML3P/s+sckhwjzXFHIa
9iBy3SEavvIMbSO4wvHo6ioW++rPrVDcwf3NEk/j6dU+jIWQSzvcsG9JXitLUN6R2+IUs3aN7/9u
f+TzwK+fvv7cplw2Dxw/yh3FTnIguI4fNt3siSMsij21qxnqVVrdj3qlmXpoRKUkmg7CpvKsQ+nD
LfHsfrJxnU2hL8oFnv8alO1b68IGvhzVqFNEnl7IDLseDNy7iOIY8wcfQPRIBkeV2lml5P9zw8XA
bnNH92lXUgCNOSHFhweqk60dO7m3k7XXSPVuU5kkGVLoAzB1ZV6tbVS4g23Ekrd6h1LRmFHNAKss
KYsxUBCScqhJXcgUPmB+yTL6NhI0TJnRUxnQvQ8SmPI+fbzRMYYR9cwe0G9wyUcEss9WaO6pfeS7
bjNhVccGilHWEo/SVpuh2xOOZckdLHsuR2hctwxYifhEmm95AREu8GuHqiZcxZk8IvP8NelMRcJb
wXrHodQHt7PO7QvA+24sUNx+VIWspuJf0/D5xdM/q5vYcSEgkcqhvIQlbcSJamzYj4O+D8AY1cdW
Rdei7w98GUHBczOx84c2iqY9yOR9tUgiKyzp3vTu3rF8uWpSyol/8BL/RLs5V1LQOdCuk6AXGLDX
y+DuO93qAvJwUOPAL541SzZI/WKdGeBNbGYgTbxHbt6KUHxZlwxLbUm1GoOgke58afTT9wZXqZFg
2Phro8FyRpCNTyk31BZFaa+kJMiNZKa2oipIlHuL1TThx0HWET2larCfyQLx+wAJy1KKVKZnJJqN
/VyqFExGyP5POFeMfVkasir4ggQ9zdGbwEgn1+XsOtuuj926Jjnz005euND1rgo4AWCxyVdnVaJA
krrDv99bsPs+oDJywveESr/C4lEYy82kW7FYsmWQczVWb08ZsWLxj1rQ+C+3NYl1aEXp84yDrWcB
/cnzQJAOmSrPd6AvOOMLl44Blyq5WmvDw41ty630Z3rP5Cm5RAKsyWIh3Y+WAUAWdsvUzgg56AS4
jc8040Uc3Jn4hfXoSk+m637kLnY5bP4hIcWboFZV/8R15vm7PxQI4p6cqidJpP/uH0yqJaJcUwDR
hPqMouUUCEly717sasdj2QXUmcPsacO4lF3IrVhcw9YdKsQcsX6v+9HbUvgcktfH1OBDCvE78mXA
tEuqExhbymdbUJRgOQBfg5i9YLQ9Av0gD2QIGIRDXAtfjAzNjAxixMjPrUKke9Zq1PAK7E35Izi/
blzT7t9i0MLqK5TecFpujajCClbNyfMKFBG8AHfLGIpps4nkL18ky6pHYZu4UlGBEywogfq4gF9u
7FPWQ9rNYxWnD8HAuLXcOBOYQgGtMl8iHktVnccJUt76F4QVwA0MlnY/CX185V1u1uzmSflYbr4C
XdQC2LWfO0bexQKNVHyUoupZsNAg0eloZllKOLlPuEx9VSJVk1hR8Rb2xVWHVZkGx/dkXv9arsmj
9sQut5wq49Bt9Wsy9Gds7Qig1w85JFBVlVrpb8PMbmuQXc4tgqussWBo2LzElvdWBvFHZMTwkq1T
dRQEeiSSISr9AcogTnq9LhbHhkwobrQgvgggsBKvKhytlpE+AGdUK0cA3gk9gd2QfV9XVV9w573i
pKalHOVpw5bm1eiNLwFfb4gaE6bQI4ABq92DLmPoFDJfR6hoRV/kL0Vgcdb4eOyoG4CG+n6CArhz
l0H8Qek4XdSnulIZUWzDGsnKhfU1QTGbjNqCCshyHb8cD1e/M3rfhlMQM5pnv3meCguC5XnOwCfl
GxV31RIu53JZEMprnLj/1+F6YXeWv2d74sAvEImrt9K6aa1F6P6M7dQdAHNTqG/KVx7lkRlFU0Xx
+SYX5OLNt4FrQqxfwNEvuFYrgrUDWIjydzpeDjfV6bFWYr1yZV7DzIdnfa9mpGJth7RJsvHZkO1X
FBxKlBBGF1qhG+Hf+v7Q6aBLmodtPBpS1n5DJcKWEfcrUKzW7ZQeyFc1ArusO9qKsNYUL0WQRRHC
Sbp/AykT0v6ofjvMwHFtp3IZm6PI4BzQwAJ+QxUWiy1h/lbO8xl3kZSxq7/RO+nGfU4+iUexO+Vc
j2CBVBzLcHkpViNDXYp6Fk2HEcRsBc5+IHQ/mT09k7lCE9TNJjfhxDwa8k8RLV4aGmyFPiieEWh4
3qll9FwZrGKb8eLsvMcs8Ij9zr+YcOJ9uBCuMmhem0pGBiErgUJ3ZbGmwC31XL06/jN3pmbJq53R
fqese/NFqw/ZA8gXuhk7oMviamdkwP4/B0CeqQ4S5QPcAx7BW3sfp+swYiYuXHzhEW9SxkRET7ut
ebTcrVkK1BQciB/YmHZpVMsbS3RxgOjT93Zsb+EUcyQR9s1P81Ge37lVnAvWYVjwGCIceKpCSPMO
gsioBkQ5sK/VZLFe+NrCEoKcix6UvSzJFJMHJ2aT8dnCK7J0vBCDp6oAosrRx0HlZkUSVJ5q7+15
qWFXZLavGBUdwoIqMHO028msscamBxIlZxs2t3BvLXfbx12lZgqImQFtrNed7xvfKRzurBp4h0yR
Iac+V5WDEfHmaePB7wvyiIlwXq/nM2p//x2ZLcSgzKNmFNw4Bml+/Dwpkjef9hzYBcokAR2jHCYo
BgNAD2jY0VQaL4bDf/CFpe9ixJuZY2u/l8XrN2beyEFOZfVfIjQcNFyYW3U30bV0FRMkij+PngSg
pD2Z7Fnkn7JNA3hqj24CRxgjMfXTqEuwMENXfjdY4d27rUP6nYyiKqRuNK9v+3WriDVZL8B5+v2Z
hXST3vrg0hg3iNtr8hYH5IbgCt4im49Tnof88ReL099AMNFFkFUEPcYGbEMC7l7PleJBdn+0YRge
fqszv+oiDZsA3nr2eI5TSXKpC8IC6qermIx3OkwP4Vaa1cJNm92wbA3LBJUUKNBSMpxBtTXYu1yg
HxNXXvvC/jiYx5jER7PwSFHf5Si/8l8UIhD3iuE/wruaQkhs3HQpyXb1E/rBZxP6BcIcY0Ucqij0
zEH8OPoKmYT3NAKwwShdnsq2yyx2vxZyIscGcHaUG1DKRzC9u2nuqJAxoHbhnJtnPuFo/KT0/Uir
eSJ/Frh/l8yuOYfGC0Qqc5J8Xe/BE0hx4NZFvQgXn3Mhd5H51OHpvnB87g900cJQuTAFBFcpAbX5
VvuRENCJ3Xoi1p8EGKJLcjocBKHlS+PCnTi0LM0PwRC19d+/Xlc6w18/anCXVZMj69TM5JU0uRM5
iOfVsBIOfVBmjM1d5XqElgyclO60hNhToy7x2IrpBlFbg1OqfevpblgoDTIHPg3Jr3DGyQZziCvm
LtoUxjaR4zi1de3S8Wz8IRfZ11/Pu4g3wf7xS6yK4By7WYTmA61E+HIcZr9CSSIVEogpnLbSdUuD
qjVwd7jX8EDMMY3+KIKIGj3STttsqDyHexWpDPZqpTOF88+GISGQcnPm4surHd7I6Ub8YtlUzc9v
wu/ktkCLzkKN1omKLSCN/Dmnvzalzi++ZpUmN36F/HeuYv/7/MCUcJ+A2T7ghzExNzmC8akUCXEZ
CYl7nWBBcM5856vR8WuXAB9lTxf8R2wMsFwwQyIj4iNsY2752TN5Yz3uhgT8dDyl5Z2ZRr9D1WMd
IR3KO3tdJWWX7YbOcKQbaFadnCU1SeC7t+gssN3KCggA6D2mQ2IXiDToeVDpTsaorAwaTAKz2E8N
CrWSuXD4IoNARn8MIYNO+YKr+qZLD9v495WL04oMakgi8BJOdRv0H7/Rsvu7DREVWNGhP8ckxr9S
pn0FB2XCx+KtNL+Y6p48NjGg4wklYEGAzYytg7zwz8Qmbzs+m4DfbUR92cz2vcVIi40pZCEitqkW
4/Ml0icUh/P5TnU7tFSQjOfMmZJ6voXYRGtOYYSdYpbxQBhRNvQlh/v9DUY4Yh7fP8AIOpAiDdBh
X6ysfuyf+qkr7vSvTDJwdB+/0cbUtllYI021v/F1v/rfZ0p4UvEDai02kH3AUVedPz8UNH/K5QBE
qaPGy50fPugwAoxXs5YzOnitP/66Z/piOtC4bbqgVGo1rs52ybIh248Y2LPbazLHopdh0K9klEMN
xjDO+5jeiR0grVcy5qYPDXZKJhsD95jvz1yunAY99UrkrJOm4K5IMGPln/SVQPRg0jWSZOspO5bY
Z8M3QHXn6gl+khiCOjzlmPIGnb9t7gWSN5SvJg1+4tHJQEKr1dHpUXQ7reryOvnDalqtLbVVV0Lq
JToQSdTbjguD8AQ+u06ubg5tuWtHWHKcmnOPCJymf30chOlw1AJDQmKu6SnKgaIHhxV9JjmFKEtA
/V8PrhRa9sPoxmSf6eEtisI1nIes1YO9RZEYtpHmYj1q23FaETlu8h6Dp0I/hA7MlB+4LD03i+0M
kuMo1jIdYAuwTaLQyCcy8FtHBmbUTHJCDnvh4KngX86uA3g0GeTJaL5O2s4hFEoAvUr/m3Xp/Vvj
IIRwRS02woDQDY2fh1QLmBcwumW7GihxJpVMIgq7KSt8mSLPipInVAzXdWxVqDeflSfDrCA5ymPO
NWqj25KPtZoJ1zEduYoagglAMhhlGHkuEs7KuOB4AjWTdxUVQYqtE6UJt1Bbk+nAZtv7lOx2NqAM
jbG1qHT+GaGt0dIs5XLvLGuSlQsuQmnHuWQRmdwFfUepOL+lh4oOwccKfHtttAPgxJtNvVJv0tHF
zpkOGA5uv6hh03Zs+PMHl61ZAExppX1bRS9jQ+yAZQuzIL4aI+cesqpu8fWZEgUsY4sg/w+CGOgl
tQ32+PHQjY3CTZszXE9F+c0iBTk1NNtM/CByABwqMs9mLwmWUwZq0jBGoik77+RoWGxnzv83IaqY
PU/XWVxh0GWwZdHRn+hXlLCifjKcIQZC7i8WDCFWkt79E0Wg8Fhs1ak7gcsXxxK4zA+slOceT1Gf
z7OpTCWMjmvEkX5GZIaSqzxvgyZ2eewqFcoocHwPUWlxhBLuqru7pXTQ+VlDXx0dPjyPs94pPFG8
dIqLzW+uLxX1Zy1wov4+ZmAg7YZVmFXlZVJwvQbseoB/1Q7IzhJ0ZpSPRTqCKpQDh6XjapDfUQzW
FAoHRgkghBWYFjN2H++CLP9H2Pfu1a63p3UsYWLr3aJegerTGddl8reOn36PzWeLcn/59qttQwZY
ZO2jVMBac6irOwwJAyyrr59nOOfE2/pZBUMWqhohjDvJPj3mygZIOBu03VJE05qOr1fc4FbRColp
B8TzPpY81Wi7/OqrId93a/zrHNe9OBpjE0/5ZE3fimY+PQZYB38zFT0LxXYJoZq8YJnHef3Nlce1
xYhhUCF3dGkjcctGnlzXF/vWBS+/f7GfsyGEaPNhO8Rqw69oZage9/6RuaW+KM8IyZPITPf7x5Ii
Fta/LUUD3u21bB1K1nhaujopTTQh3eF5plFZkbxtytRWsQG1vvFgTpTGc/DObS65fV/3gH2V23tf
Dvgjd3ZZMmuNmgQaOpale1q98vZvBKAWsuqk31HNe3KifODz0X8+lza1eR5oLSnWDax0OULkf/Yl
UG5BUjEHz2Egw8SqNe+LRLoX6BkkogXxzLMv8x5ZvAQU3M1WvcXn1WMdDRKsPTM3GnjvziAup7Vf
dO28TmGOko/4zKwiT6RWSgBqYow77KFPH0Qn+CB1YK0K+nHAt++npiSu1Ubtps5f0Tms56g4Yocj
/d8H3JjcJJVvH3H2or8Ybc6K7QG/mIg8HWB8OFcZNuSS0mrQTg7HAmjmiTP/qs2RX7N2Z84QZyEq
AHzdO8W8la+lxNDWbATNFdXmncwvyiFJQkPU/W0ZYU6pWffvia/YQ4kNfWlMTW9UPdefBs2cstff
jwiIkSCiG9KOm/302rIaJttdvyJsJ8mrltlK9Dqg9ij5j2CQSjlH1AC2WbkBuYyfH7woU3C95UnZ
QFWP9njRSTvGR6El1h5WrSzLn313p4KAtARobKejk/AMq+GrxxafuPuFC/oZPFgV+7QkaACsqEBZ
699fetAnzEEwNpfLx7L7Y2LOdqjw1K0ebALDHllcX6+UJZCVfmkneMiAB2WcmECqjQ8Wqn3DWoJo
NYuYEsQvEfRkS4I5a0X1iBDDOS65/mk3O1u3MQlCstmiHKqbBM8LgSGCxyGkDJI1i0rNSA6hbPRp
cxpzGlPa2ibK57NApwRTuIBh7K9P47I6w2FxjuZHxi+EANxiCNR31IUewfDGNg36MQU8BVX+S+q+
0VNlqqOCCkuyyK1t7DR+NVBAUN2Wuvmsk6TvFs43eP8hOBgE7x4vsKeVUO+PnTaTGYyJ2rSMhKOZ
uEKziF8RKKdjg1GIpkIc1IbFvt1zsLd8Bd87seAR5FdT7snXkTb5ZjZQ6tnUQWqcGFuTrMRU48qw
fFcSDQZ9gItpsSA1iLjgRehImxfgL/PEkhjReqID8iE13neq1umvogmXxXrdD6C3vlWygCmDWGc6
BvrSrIwBeq0LYc5u971mAi5rN8XudNkdcg96ztJVFxK62QRWgjTh8mAihtWR+u6HPcq9FMOGmSco
vvTHtK/BW7e22l2TuG3mq0Ij6I3EjNYspsI0RruU/efXDbRnNghqasMrtn7NlRuJhSePwF3tQkCW
gwGqMjnkLGH1RLGDldhm+g66Ph8qFxHCBhoT4JJXyr//PLqQfN/qNRwbpZUmDi+2nAtN/p/LTsb0
5pjU9hmh967cfDNmD1qKaN2ZvpMqU71M2cpIcKs0whq9C3M0Ub6J3cFO2qsW1CHiSL5aziCNfZNT
pt0b24FDgPGokfiYaGn8yRMsD6E2MCIiu0295SdXQ6Mn6pNQ3mJycD0mrwZ6tqvhVfDForfXOHNW
ncjDx9LR654fuU7e9Ack+FBFgVPtubdkwCCoTfgysUQYkhwzjJcG/vDuHqg9uVJjYuX1u3pwfTRt
S/nyd4GvGESYKF3GO5PgUqGbLQYCYVWIV/klN1BAdYznLhGVFB1C7T5adkWGAbQIJCchp/VAWaks
VYKIOI11kQrjuRuJL4DvK0ofCqkT9zlxi/d8y6QRQAi3h82BJxVQq/8KNIXt+wL8NXNHoi6OJR3Q
3eEUBtk+cUc03CHvZg62Zy9DVXrLfBebDpmNKcQgQCwWxfYlAcQoYX9aKCErinON2ONcqzYBZKeU
8y4O+Dh8us5Q23T5f/pGy2Fr0jLMIbp8eBz28ytMOxjGRsznFmFzPQOG/+4Ozld/MDKCq3g+zc9J
M6c7VWyCHeec2j7afu5emLlpgzGbPszh0RjKYsQk+vZfhD+3Ht4bJ1PSaQiUAXFbWoh9ltxueHQe
CqBHReQvCzZA8X7UIjMQ4b84z9HZP2g00Vs8KIU6Qa/t6E2Ul/1Qt/qfwQZlBAawsY7wt+uSRA8U
RnM3+LWJdZQQJKanJWgO6rdTnWEkPH+kpgQWGZTPHTvWwkt/FbOTLyD9k37kzgnY+Wrke4G8jnyT
25Zz7cRYiU8thBtMejWMWwqd+CvPLGaQn++t7bnbaxsuTfkVnHOUns1gvxp/JyycWQ/qNu6o1bqQ
vsEI8gJG/SopmBPpv/KgwuNQ0Ya3Ug98PfrB7brFhjNWYpuWoJ//DDnKI5DRxicAqOlpweIYhOzt
NN7d8czfX7Qk0C9YkEqRqDtypEhK8NtSSyGdiN7ZZkhLtZTpib76K72eha1LZO1Pyv79tzI8OkBQ
FaD/rDH8fzwG6cC4o4s5Ec3wA8GDnBcLXLKtBsaLtBg49h3qALMaLDE+xbcQ8KT6akjHRrCHvbCp
hQyLbQpCrygE5PK3e1vCIu57NrsQNEvuepJgqSSd9alc/kELuIfvxqDPD6Az8JOtlxPpoIbcAbCU
7/BL6Tr8zmH+KxkW+i3adpl5hZFjegYyp39VJUB9YRJFmb2Yu3laoi4wo88Ap0Pt/FW2qs40B/UQ
snG1T65GGQOIBExFAQJjD5pQdZHVHAK1Ydtki76tXuputIeZ3Unzw4VpQWi9xODMJF8PMQjqXNfh
cBYNfBs6jwN7osGJEWx4aMsb0rni3cHTQzR+1gKeAMAuLUtWIIvZZm5ga8LLYVVDZ8Ze0e5iPrKp
ArnlX9Q0CFY9jkFG3ehhxM8uO5Utfazh3a5EhMKcR9oTotRinZbdC9bAc7sQ/b3bad6Cf+yIdbkK
UHvJCxA9JrkYe3a9J20jnARCwzPOT11KSvw9Iw/SUxdwaG2TuAWMQ25xxdym0HGqiRhwiDmmH5Y/
HZL2peAJwG0gUrStHHxedOq0o0KMfM9Ty+0AadQ3Slv10EnTuINm+b3Pd2AeaqmwHYOTCxeiq0sr
PLYWj5iF92/O+g95eHK/PV7L2u8SyiFMlQZRz5oqrTNNkVjo3WycmJzHnxyrd8WZFwK4bEe8bpu/
WKZ10yDYtXYViliRI/XhnkiVWfL7KQBRi8XYfL4sJAuPAP9Po4cc1gopvR/9tsv65VHwyX6q5HUK
FIdGz+BbFA3AY1pSHthUlRG3dUHgxjSBQDmwuQR2D3b5gbeJ294ZvlSYpkOvHb8/cp34t9ZdgD3k
iU6U77E/HLfuS4eyvWicwoPzHyPPMUBdlKt4Esv873OCn74txIeFvrzLdUIZgykDcaDBPg/Ujhl3
4wOpbKyzLZSJNMkAFmCF5Hs6vAyY96pj3BME3XCk4NjlqJymjqMXi3AUtEpOxp3ax+VXY+wZfvrG
gz+ueXFHXSmNb5MkLpYQQc88ZzWzy/TYJEK0PPMrq93mnvM2clMDP9VED7MuCwNCX0AI4tHW4mFp
lq8hVMIn1vlaVB0mFsZiQRgJ43aiqzSHKU584XxjL6zqZdQKWvKkluLUNavosrhKn3Rzx5IzQDKn
zlvRoi5splCMsR+JuvvZXLislgAzD0UvQxGnZZHhoBTninAOBKYxbwYFC//oe1PvWSd3IHN5uIRO
FXI61Xw0YfNJqqbWqariJbmbz7VP0jAHE22c7j0Ri0TJiWVDoxeaWJvT4T2WmWR3Y0EVz2C9l+uT
M13iZlk+TPvvS4lObsxgZzBUpfOUFiWfDy9u84kx6urXd2CowYdEN+kVKg4n/LoiXd2YgJZiOaFr
mzYvF6kzMUuWcRikA4Le8XcDFG3uEkSFpAHlGfJELvZw+V9SKwPR/Lpdb6X6pEsr8FVVha7ayfBG
zPK6C2fK6NHqhF1NSNYxo6xlMIyAC6vFKZ0mTLjjdClnNHTKaZf5NzjtCgKag0pNDAuIPuoKP96V
6vKZN3To+eMiOVkafJBgV/oLPFaEOGJeYUtyUPdxYzYYPaSC5rj08ePfnygJEc5lEXCJsAG5cKE8
vALg3pREzIcILQfKMsgTMRSmNvPmlYO78RRD6D8/TjgkFuqm/JntRFaeqvDm1u7uLl3Hb3+ZHA2+
29HEnfXl0U+zR+xatBogFDGtP/wURp7QID1V6MG/b5eeiRdkVkW2E2O/3ImnKgrJ49bB5GOO1eBD
5UUkU/uREprPCgQDH9cjiYpgj1zov+DCTrXJOZve4GcAfrUx8n220DVwOTheJwv4MgYvB1RuTjtS
tYCRM8FMP/FrwUOhwTwfxJeOSTmFD3rKHexL7dtNWqYfxFOTWWA5rVr+9wnXLMqdaXqMUvvLU89i
VVch1l1ygK8UZeU0OtlMGR5pFkYLoS4ZTrcoKna8OJqRA1jdnNCtCpQmeovGWpjKyw9Cm5pBIDZD
tAwVwq1SoY+AB7XNre1BQbmfiQBQvQfWOEphkpab/Vk8zmWv9iaC3THHB8hVHbftvqBuLAQqiC6d
5Oe6unawK8uFpw4pHkCQqxMgjO9IuBXXWCCwCHtoVs1OMWUUuO5epm6nPBdgiBI+Ab68+nuomwZb
evpIJRyOs4yKp7+zJ+0FEMBfO7Q=

`protect end_protected

