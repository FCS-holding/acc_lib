------------------------------------------------------------------------
----
---- This file has been generated the 2020/03/16 - 11:19:27.
---- This file can be used with xilinx_sim tools.
---- This file is not synthesizable and does not target any FPGAs.
---- DRM HDK VERSION 4.1.0.0.
---- DRM VERSION 4.1.0.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinx_2016_05", key_method="rsa"
`protect key_block
vroPXXcL0qezwdrxLwgPGR3ghJ5UreVjmQbhSLg6VGxrzxP25HvYQZPWtXUiiDU9Yg3hPZXN9tvT
gsO1sVM4erXRSfB81Qo+p59c/0XS4h06kToA7Z5jHd9eillirWWbjqUGuqWQ3h5GqZQsLaHNRSTT
4uMQJzDhyvaudj/S3QmOehPbf3GjOb0YF0zfnsN7pecstxao3VE65k1rjbvlDr1DvXFoHHc8UgrL
XMGnAQWO6PcYvhGKoxjPTVbmccNTIhd1KCOIQJCTKEzil/UGz2Qx0SGLQC+YVssEMMGGT/zRurvc
M+c/Wam8QwP6hLh9HRWRJwJXiY9OFUd7Fn1J8g==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
sAuuH+uz0jP2CYLhXPdz7MvfOKIwX0OVvmmDIgwlKLBfZ84k4JC8KBFjTcfUcOnCTf77mCZGLkh9
3/ORf8SNzScXNVaeRUxehgJ4AiRZJj7pu+Fb7SdX+VYVtdRWVi93AOPB3saFwWaeDdcUepJbMDHp
xByNyWzEm9sqZeoCZKprpOKj6ubKPkNQmaHiJU5gcayxAwqW/VDVdNfnHW/WGKzYVFUQ5iSla1J5
2PrTJZIzf7KLq+fTo04iOLujzybApvebKDHVzcRryg1t4ZXDNHW9VOD93uNbnEVDS7lvCkQpmTqx
SAsC5AdXLMVEGLvOAkZzbDESSH49+nfm55OodQ==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2019_02", key_method="rsa"
`protect key_block
aLvLH3AZox35NRJNXEawgD3HvvreL9gpkTol7bKEHhB6Cjnf11ZcN8eo+97EunYjr+0NJdRGwVam
FaM8yOktB2Xx+6n0FQTatE4pQeaRz1c4GWwQ7m3cgO+dWjuw4sNEvJGME26wZyav2DcsDeKh0o0B
DqNVdamG8JCFuZnLzewXDqkKMv8wz5yKH/Xf18UneWhpZJpYTFvEO3m0oJmNQfBtEN7M3mtCgc0h
7oUUOCLSzljJzTglOBd2n5WfE2LPwvk7YR+z5mCTcVudtYcdAAxuNch2eYeebbNApsycGTqm5MBw
2pH9NwGPA7k8NSiAu67C5hLkoYN1hHgPcrlt7w==

`protect encoding=(enctype="base64", line_length=76, bytes=836080)
`protect data_method="aes128-cbc"
`protect data_block
vXYl3m3JsCUGzWcCy5MFe9YIb+Nxdps9zdv9iAVNb8ZVLjEabBWwbnT1oWBPEODqP+cSDL4K1Ax9
du+5AMLI/apmt1E7VWvJSD2hLQXmwuYNc5e73XeNqzGmxgNG7uGORubSlAwJLdA/Fr5BS8rum4je
KDngZ0QIJhmFsPZliz+Vd01oQ81/pnJ5gHgO/rWSOQCBNNmp5dXXyZ393H30QoLbSNYjVfR2R8Gf
3JzywQem36kjBuV5uWciFrluAcHkrZXV7JrOBqlXRX/AROh84JlfF21H00S3idAwOwEjhg56OwiY
NaYExdhYwXRBT5DvJiSDJTyMzdewpB4ZqjdDwuPV9vswJbRRKuwWIZRN0hIF7T1meik2wJ2spjz8
hDbzpHJH1DAiSIUxxi2Rcbz6pH8qe6S1gImmYAGX9yI9MFnVz2qAp9Tr9XmPfnhuujSz3nubhA79
kdZ4jsXV/xmANlZ5myBsqXoMFB2GYpE+aL7OK3hOg496lzHAAEHrxGAHXfPijxNGyleOPUh9aw47
jI9uC0AzhkNVFbLJSXzWmAwOLOWG1vdvjFuwimZs7z0M6UGY9KaTx6DZafX88KMG5fShoi716HFm
C1K6wUjF4mdIGZj6/Y8kVaVImMxdcItfrk7n7EJjgUAzrvZtLdy8Pn/3EDKXK906nEw0GARyzY1Y
V1IDEPyrxgUG1SBl6D7tAbOHFQ34JRO4FN/OtzCingMUkViodg8HFZdcp+IfzpMiUrpeezclQ8iO
Vt55I11TdMxIuJl8w0w4a8h14ONn6vBHwm+knaBT2An/gRmiFaVNuYPeguhI2YTbh8m2FrVR5JYj
lNSWyYAtRUL+YhgzjFha+Dlz/RngIsTYJi7ziLv5rFQU7BuYYIejUFg8bsdSolNEN47O9L/oINp7
FW4YcnzR74T8ZBfm3jLJKn/yHIIXKMp+BTDysmJ9LFjN51YeDrMyRoYm2qZNRzxkhe2b063g/z0X
7FRY4XBykdHbSza7eRDDHUtxkfwWQ5rmk/oFDzpdtU/w/3UmWvKJm477nm/Z86oTvT6xiiz0Vug1
tYL5msXXufZtKhnQmeiftUKGTw5aq9203rbGYy82shuvYcc+jvjI9ODGKAmJGPsalpfQKRuN4ZAD
gnJVUIUmEgMGNm8ec5awSvvZonDbTOX2A9NONPg0RWa3lk8FxaYHNsOjizdO1DhffxtRsluLAy9E
IPIReI9c6ELZp+ZHXaOj9A82Wqa7dBDaoIi6tde1xmeUxRyWiThUQh1uGYJGBUUdxBMn8nkAaIQI
AICJGmQt/xIAQxaSjoDg7R+DUUtLC/BwnVvCozyRLGkFeF8d0XNve1IZc8ywaytmnPLyLAv9lGEn
XsQtNJtAFfVPG0erVtRh6WXGvZRixpRcHG4ickiiTPGB4Jn+QdwJLRW75YAGFMKjaUq4PQH8p1wL
1HwoCspOXo/I2oIrThdKQwX7VRHaIZE2aXKEv/M+ZEWo1bWcvNNPuLCbghClC+dVcInEKOgk3CAv
x54vVQygHTM70l/gB+mYI+1oq+ZKExvDjlAB9TFyPpXeS+XJQ7Gd6IBTzvaGZBKfcReiWAVvhT4N
acV1kGs9pV585QIBr9fMQodlFTDVe4dZj7ZR/RouzumfPrksvqcCGQMGJQD+xK21q11D1jnkraX1
mInQ8VEtXrP9Ex3U2TwuYk3eXA57RtCc69rITmxzsZ07PM97zfdSJvN6jt9su04ifjfITlAhPOXY
0H+Wny7w0b1KUvMrdFq0Aw0wGmeugc0c9yVQrvOMVxxP+d9K+sgcABw3l52zsxV2jqzqcLlNc82f
YN1K+REtBroQTQY3vsb+vnWGgmjbi4YLYyav7CE45IS/AAsrzPGoiCRPK8nD39lSUONphqynuqzx
2pXiRchY+UfteGu5wo0Oeuv7geijr5ejOh/vJrImHFogTGJtVPWrFBAUgnBTx3BFOmQJgBUgkans
TClcZ3QiTmo4/u50VnpvjZQLZQQ7IKkmHlftLcWfmFwzflOqSkJJScyrtYeMUlnNV68QqVhUYXaJ
R0zMqgoyiGmYYFyPpbDK/IXdPI2Fe4qaPgqgn60E+vl+SBLp84+o6J25bSodhLdK32PdB2AiFtHJ
d6Pi7EAIi6bUP1qU8dWuEzSnxv+qs4s2uomaCNXCLx48jez4oN4pk8wxzrcWkckCdDkQ7qaBV7DB
TCoUJJMuE6AV57Hvk9FArEpJspqfXmbs+TM522s+tNYkxSC3tiHLbLkRIP/k0lo2lqpBHYgLmpdM
SvghwW04No/zdBJzq1YHaOP1wKfSFinu+hlJXRH+dGEudhTxYLC3wNFThDOb+gThzDQMyMLuLiic
7OINlZP0l953dPpbT3lu3MpjGAmdK4ruz3t5to/EK5K7xX0sYEhKQlIIP2e3tpceCUm2L2+1rzqO
memV52bjxUpzKoOSthokdnLnG266wMY0LvNCyOiZT1npS/uqVqdFBbHBkyCXGMZQlPICOjG9B8WM
D+Dft99UvmtBD0wU7HfcQlH64JoYEvVZwDBRhtt77FbHR9XrRbibSPZ2QtTJA2dVca/bA4oOMpS3
snG2MdpYbJMcKOMXAszNFCxvED/CpJhGVsHyHPD3YoiWXetbBa+dF8d/WEBKDn7QWU8k2/uRFrGa
d1DloTJCABkIaww1OKv7F56Lu9EF99KUMOPLkuT4OOLPJ3Lup+WwWtcyS/YF+aIBkEt6e/vaYjdR
JVVYCAct9rEa6xuB7jJ2BYKpPCnadyQFsG+7eCKiJSrB3mUI/okR9xwCMmMMkmX1GAX8JQjzhNgc
bAjShWXEzrJF5LjiAT3lcQhHPDjMZCCfX3Srh/GtRWrGYfJKIVKeBolfHW5Km0uSLTaDfXTbm+4o
pyUPvyqCRUq22pQXOV/9SzH9VWxtd2c0vKjik+PEMlmoruS2ggrjjSksoiPUIj7VvAUmzZ1DBcjl
ok2r1XzhGiM9YOnjxvD/FBW7Yg0nFgqtCzNBbh+BjRZWx+NhUFv6CzBZi9ewPJPbV6vzbHcnvBUI
IqU1VI5gbfY5isH0lH4bm43hyLXo4Z2Frg5qcbVEhioSAaektlb4nwqxR3Gt7iuATMYBFnv2fWUe
D+xLdwOc3OS6EqUXijLzCRUYyvg728uRmipYuj9CaLecFlCqgmKPsMrl2v0o3geIjPdZ6jXISdMU
AOgZiFz5yHFMRFgygCIzaCwjkQ+O0HhvFQ7wP9KnqaZVeA8+hPiindx1UeTI9DRRLBqUMwLYVNAU
37uKsMEio8/d9G0fkbk1qrpaUcC0bRHPWCnu1rBnZmsRI5dHbC/9bI3huQ2qyglInd746MM05VQU
UZde5mSzo0ZhPT4ChdRgHIG+NDgqHwrk5iTqhqCRTXRQcohMm8I1gWNPhokJFKzMEkRjvNKjnwMy
Q0cziOTfNq9WPGKB79QW+GJOhvK3jzyybshSmYvjURypdssliY1h/N1RcFv6FUrR5jFUixznyZme
JmYVVhOhwm/4t5gfPbLVINteouE8qH9W5bnWp4DqLXoZIyWaVY8hIPL+nSqJAYcVHRoJ4qqh8p+n
YMxgUanTCovt67OnEKDLFNl3ZfHfZ9qQ3naPDEmpF1MQNZyFdRfDPnlc+pZwovME919UkRBY6qdK
nXx1lbQn8hkp6DYuVGpNyuDQcdSCfQUUYsJrW9bV5g19v2n4vnk/LfSOYSBfM9AFeMybhB7hN6Uc
qIJ/sq7t4n+PZkhElc1/zRQueahspppebj2ZrTe+2vnKOr77B30kW4lOFBM0Gu1tB53NlrXPZn77
pS2efmyp5x2PZp8hgRAFfaMkjTj1kvFjVsePdtFflnyMdyLNf9uGiRJ7fGTugy5kC9SIAD4j+Szo
sYgn43tkTZPSfpIhwhpNjIlrwvvsBYkgI7eWC6wv5QtVHdTPhB0Wz6Nuy7OVI5KZYket5kB9FAa8
ReHPupPLuHFtj+mdiEpoaOv8R/FgRkwr5SA+yAu2Dp9NXliD1h6sQaFE2E4tDv+7bSTtj7MPg4U0
LB7tIlHyQauuRlBzOxwzfb2dbFNc5DhDkiFVBQmkI4NlPT6lCpIX3vfHHxMObmd3DI+Zj+wrTYht
gw1XyyuxIAiRK87GjaNJlL8PPfMnx1IfmV+0vK7Geywuz6sNeQQceC56maTlCwXN3gmz9+py0o1s
cAOCYp1s2cqgFKVvpRuGK+8RgKL3e4g6TEUJM357HZbSjNcmeFNJiizFb86mUcGHsMnUGJ2TP5B5
EawH+tWadyflQJmGiKBVOx0vmgUXjEnKSfOkZUY4QL7tTI3hlZpIvj3/zSnK2jRdK6CzwMwRWtxx
Pyy8jNXyzfeSu+MO6aEC5Lx8DLabVweZPt1Xasy2WVC8ApIz+SFPFnRsXMr5irQQetnBgpsPp+I1
JiVN2svyF0ShB5H/2cZqjDd1UHXv3eIX+2m6a1tEywGm+LihQRd7IsrT4VCerabb3VPbBT4C6G7A
HrPF0lMbom2MduNWWd9yoNFQF5nwf2dC3HB3gXnWK2DwCdgIQNeQFJMNAKjhmhDc0kTE+WiTrGXk
cn8dd5HKHls33ucdjkfuGWteK4wGOzbRyKT96qECWQJ3LgfRBoxHJBHgktK+4yKyaPZS+GE3N3Hn
DIFp5PTKQkIavefGdT2KVwrTj40eMqEp1vI27zJait3dDpRq5Z0buw/s2DdLyQ4P+zVxuhoIAjh7
czvQj0XFNtwkycy8M4JdWviVLfN22/xFI1axQK/7lSext+CuTnc3dSqHM2w2L5qlkZQPdQrtFs5Y
Nt7DsEdsSgCdAHfXozHXQ4RBaU1HZ82Sw0E16OfUO0XMSamuMUGvBXE8Am2+tWvlEhwCArcSoU7K
fJQQiSp8VUUNzMNbkXqNyLSlInEQE4IgENKSrjzaL+Q5K1yltt9Wiocy1bG2cuFm8rrKGGvN0dfM
kAungRdHiEBxq/zzxoQIAf4/GHHUQHfYEKRid3p1R9DFp58rD95AQtOyNoYF1s5CEO4Hz9sfdyAm
EM1mM08q+XaBl+xo8v1JKN84gfGiMeqJusXYROFEQhsmcsvSm//4f2exHS9UShF1LTsFS8n/oauB
4nrrs4HYtwnjkBluPE86eRoBgHyJxQohgncIDnQKIVKnmqYRzPsG+XxMpr1pnNOEcrWzH5fUjv+C
41dQxcYfLf+1/utlxgbjXz1T5zgKC1vrHEFwaHFBDJUSRRzHy1vH6RSrWuvFbGDecxY8ENOfMTv9
hnTPtw25gBabOXQD6/Kc0pk5+H/lFZRz29uPk+b5VV9h8TPEfWCJDDb6tUAR0DcupBVWawz8UBUT
MeIeTv2oLSiuxK3E4dJ3htT0vB1XqBDd8Cc0WJ2V3rZxP/hUe0QBtYqKvxbL9i5hEiCdkiMBAO8x
tyY4wVJkktD0lkDNbTRhB1oAf0HatCV0kbTgxFHYtYTdS4Sw+j+H7qGryw8vU62uScNliWtXRS6b
I4C1sIF54j9RgSH6+/ostW6NNM+it5xQ4Y33WoekSPhUEMd2vYZdN2FlWr/wOQrY2e2LgDprRurT
tTB4a/9jYRZY+LkxymXzbYbTAJuH+fHU2pl/K1mtAFPwrjkbSR4Ykk2eV23GGr7ORa11N1n+dunb
//Ki7PIky9bybJu50C3Vi5fKMsbdcYkARn3rrCQ4TAJZvsvl4JJ4KEmlnuc1yR1QvVHy1hFrbZ93
odfH3Dx0AAAFTIa3+PVAhaNJJLVg+XwynwQsSYF2pOkx4ehJoUlnDpZGNXcOfz3CsF9D5etSOOnR
ty9+lsEQIqkeRVa95mQFsun6qA79PrDHpba6ARrmqkEo9/1zBs9uK4ycUVCgSXUkyFZXcpU1CV2I
G0pSNLYSku373eyVwYXSuXTeqQ+OFzAo5cKa1yFgiyDQIwNQLdpnzIuwFncliDR39ViAhdEwKmJj
jUyhlI4r6xlVPgkWOex06fhFAgh9YWUU/uLo0fqDUnx02XQct7nyu6UXDAjmRXrzxiLMVL2CGA6I
CnuWJX5OEnGX1MCySPEBtonqWjhy095VSSAKXpNn8OhYn09Issz+amRzZZoTqHVbwRCA3XP94iCG
+zO18pKPQ/1gRquoQa1A+Qypq8Yjgcq3LPJj9kJx/Smc2xU1jtwgTsqyq9OfbNbRHqUOXCWvQY8W
wN/DcI985uUfU4m6Ta40dj04TQv0hSj+ynTmAtaFVEBTxt2D0PBz3lgzHO0TnG4Xq3fMfSwl5C3X
gyHeQxXZBYO/FF+hjXxO42MwKGFxv3F422+sIbvPZi5BLJnDGNnH8qdOYOX/AZOEX9KC5Jt283FI
hYGxeGKyVM2Ghiw5luT3iANJN6AicCAp7iAkldG+yatcEC6QfFAMgnHVEqzxCMq+7R1E09npHo9z
EqHg3HRLtqH8WXEdFjEwy4GQK3z3FFbgBAH3MNaUn6zEbhh7EuTVgOzYdVSne/0PewkdwQEjLoxZ
SWdwzkyFkz8X0e6YF4IzVXVbIoD9fXNdqrhdNSeAYiUge2OoeBOJyrioOv0rC2KsWhuy8jhHMKFX
4Ygh00LORwgWZJG7+5Sq7Q3Qg2xZ+4r5/uCwNH3/leQKcaFjlwnmXbPZ2czkQ0uF4gcktAEPPbcB
2a0K8Kl3Z0ydrJ0/OA3lg9GO74Y17vyRm9TqoEvwr7mL4pZaE77r4qEOGAKDcLIxKS10sy2uCb80
1XWSFivRmEVVsYT7VlnhFbkHtBpQOsaKKMJJE4HuSpfRyOPIOerzkAQ5HOZxJGa04f8lvLW3hDLs
DXuqZ8M+716oxL9xH/lDaUrLd1o4pzFLQDGHE9dLCD6EH9JxvdPEQ9M3A8TmaxwYnuvysYTBN5mC
7YbkgAzcbtkXFUUa4yHCybXhcZX3aHk2FjOzRlPqESsPkfqwFmQOJxj6kw5lz3AseitRMyuExJXp
zRsR/lyqE4fZhxt5os8oU6pfmCnaV/i2UGWmtyDyI+Agud77t6ChkzyzDkpJFh2QJ4A0Ka15kSC9
4Tb8McxSeMHroWdkBYrALTCxmT8Oh+gt58iQ885J2peyuBUbv/U2EXmZOMtWgO5CqKjRyNIeFbQY
ukF6TaoXFhFtlA0GIolapxSMwr1sGqzrmX0kAnWJrL7n9mzX8z/I9IwG1W8lPV/E9urdfT8QW3ts
32ptSR9ndMbindTPnTIlAgJPNSLNOWtML7vr7F83MSMIci/6oeeIflBKVShA612x8oMaCWnh/Okc
6mgoMd/Ov0UvBKsDzAT/RD4lSIAVMIdsQi5r1fQSZUXRdZH+UWPPgjrsNs6UjokJ6jOaa8uYyYJc
+AbAGU6exRTTqLNqqxhCWQ1PBBkT8mO/5rkp3KwM16NctEkWbMUN+8WZwLg5631EEtDj81J85Hxx
4AgXNp8cBWv6rVIjlJuve/v4dmqBzveU+o32Tw8beM8NsExRjGLYlmLC/72D1wK3I74wCHyfC6Mf
EBTnovr1gfVKIxjMys4d7mXk5I+RJQYhGb8SNZZSWqywVg47qkAtg+g9PLqQvnF+ktzqCYZqhNg+
O+to402Y5HJgoe0qiGhv0v9FnFi1T+ugb2xSVeDfSdi9erAn28Iot+WwAhtMXR+mth9la0c3GC+8
g+nCxf3vaC5M5GTI+BIt3943Uo7HBFEs30xAy8+Q3rHuLuGpIkPc/YHeriGyrW8eZskp1ka5h9qb
3DuVRsLmmsIZFIyjBIaNZ16wLgeMoCrvP38bTUgrC3pkq41NIan6FK+Eqs0aIb66DNFem/LfT2tG
UVsyX8Eywlxfybl5NdNSbOdEO6WhYhjyuKCXE0Vb2TeXCVE6Xb4wVQkeFiMg7ymCkoqgOGsDPWNk
7SQzUxI6B1Hivd4dT3hyeg+tLlWxnPUKLU/yUqtewiTDbUmp4GxQX/xP418EcvWKrMk8lcOMGjv4
RCPlLys3i7qTA6QHjfotWqb71DJQwawRlp7sxpSf+BKoudM5I21o+tc/plC1Mpbvy5IotWBNeIsN
U4EJCyWUMVTMybI6Kt9NVP4BeG8+urBbQC+Fu3dGKTtFDcWKRC6MdPuszSC0K5b6BUk6ooubUgvg
qKSmujYtJey2zWUoI1tgDJkCiMt5D9Itl2dcr5BowvZc1BPj+WH/frVKJ1aM84DNKmDCBHGs+Sfx
tzajweveXXuV+omiLZBn7KiGOExq8BgrnbQZmlgrxJ7hg2jAtOos1hAy9a7VTuZ3uZDMDXj+Yh+p
Y/bcQHAUyGP6CcULuPujEnFKI4DOMSDe7dY4JLqA5VN5GisWb72539gT3O4JIhisSs28OL1E1Iv8
CwnXG+ThyI/ERRIHMMunpoD7UBrdbREw1v8NtYh0u+Mr4cKoaf8OxVWEPIgwBbxM+vWt4ZpKEcnq
oX30IJgabMb8NPbiI9GaOjRgf/KN/tZoGKB43ABd77EKhEU+vyBAbujvl5NCSxtB1/rwZ6HLEIw6
+1gk/oV7uNAdarrPa1LrSqJ4SadkWEuaB3X/2Qgzdi6wbcCYcVxBf9lhMNwMR2AKHBL7m/HjaLIV
yw7WsW8OUqAW5PdUtqp9rdsbRGQcymPSOBZ3yIKZOOQRtEcIKZw15CEB8Pfxg+snS7tWbeYIlrNA
NDbfL3OWxGAcc8ZHSLvwdKP+hMsJstrG2CvuZBkgc740mrt+Xjvjp1MgUJVg3apn8Io4FIjk0stu
IW2JxRo8PYpSsaNTEbih/buio4F2TP4HSxRliGd8KUJcm/XqGu0iaByth37hlFY+608PeUVBuQ1m
2zLh9j2KdydWZqA4NB93AWkr0dAc866uMNo+PfbeJ4gdz3zYbDbmHUL4/AO919QIW4UStC5IHbPa
qVtpSXhc1GIZDNK7PUu03v8pb91NATh2mkWBEBNWF7GxXpU38/os2b5PiTitMVEXixJwjS5m7Hqu
OjmdBzzeog1Hwc0q8gTgyY8vh2QOJFm/hFrPaDN8oGOtOpjoE80S/dT07Hrsht/8t+42G9XAYSrP
w2pmZG/fsB0EEWiU2/VRbBSTb/QUz2SHUgowpKZeDGxUQO1iejDbJAe5LT1QTLCAYPpnydlQssUk
zpBsbw0yC29iBX1I6UijP1BhNJURU5eAubaQtsyR9KMTd1OJQqCnn5BGXhk8ZyiCMcYZHFjiajJa
gx+3I1bt6BtcbSI95EHxk95sa4kAumQjvqdYHP5XFHdZ+HaNtTO9gzj7M3ShFwDyUc/ty7t7KKTI
uxgn4Z+dNp39vaYoAmREIA56y8rTihnvYVjNx48r6rDyu+ltTUqRT8oMFz9H0tvdf6kyIyWQO2Qb
S8w2Q//79JMzYVkJJVAXDUhX2jC15Zp6mMRy98hv+CYYNXcQy9RICz2Vq41jDjo6WO9jKa9591fk
2kg1aht9OXfvGs3XfX/hguZsWmRJOSfY22sfXMbyfzkrGJZJIV2Lt6YdQrn3XFfo+PjXYrKTACaS
9lX5b1sBuKMkEqcURuwna4Wn/uUJsa6JWuam4/KKrUCaT3imyZgrMdKgBoUpNpf/AgPJNT/Co0NX
HaiBZw6KxxGwgFUEDig04mD+lMPNT7Zr+3UhvKSgA+SVt4Q+JgGeoUsc5i9xcRnGbRIqiwaCw2dF
lArHfGWVucA9q95wA3/MvQVd1mLTKW7fbBrbBorNaWXArP3VmnjzonQF0TBgZW3SugpxwPjE8EPd
7RtwftysnY6LJIm+aeYtjeM0/eN6L3LM7H/FbfoW3vI+UBLq21qV/nU+Znwqgarfeql43hAZTEky
0IfNaBiqNsjY2McxmaCzAUsMT/Wiyj9V0nS4RclWEHmFtT81S0dUZ0bPaFlaQTFcwq3EUQENiTee
b/YMwx8Reoknoo3GCDXR5pzQYtmqXNMwf1fRGYOlbT3CLuIKk+ro9Zk0VbwDxnu/ad6diHjSez9T
LghtBJU6kgCxMDuWBz5NLkWcurHZb7GpS16nCe014c/PJslxYq4wxJhTj4ZvBKaP5AE8Hp2IFofk
PV7HnnGNJl3yNG/sVtU5IuI/YbmrCvhwVdJBSzQIMRWaFHcylJ6MwjWfKBUnVtXrFvdzP99vt+On
x0QeqIyQnUDmptJ253xc1EfA0ku+jKUV8J0uTBXTIsOUIR9yDN43tNoh8gfamqFUOBBj1PV8yPds
VyiqZ3BkUKUzXIAXF5Rwta5przAw33njg+xk5J8gv1fGVGReIodd0tUUCqDIdFjHoB2rZ6iX7mPt
rEg8ZYAcef4/HOVBP3PPlRcxy5T+xwAAWPy9BCyzXb5bxGeMcglhvcgk1uTgu2fuJur4jBXr1MB3
1n817i7KRMNdCsWWYZYu4Ly4kF7ISpCHT0NHafLuk74G786cyIzRL5CoRgW8819O5ChB9VPJPRv5
pmWfR+iwxuIxGQtWWxjkmIVlDCuboeGYwH0lXZUryvkA2incZ+3Mli+3gQTQnEY6zS9YI/DFOcFZ
adIBKJ+uqnM0cd9iFJCjWNeUqucSDDRBi6AIWs+RPIR2GGOK0U9TXSNDCtY1L5Ik69MAcIWrl+mJ
8Y5ZG49e0Y3M6NW8HDiI/cS8rr3sinTAGpSWW2Q8gbiQHYBtLevC1R6WFDhcolAo+A7gESZknguv
+1bEEgoRrMnmY0jYCyvKRiTMg36ZpA40MShfukU6tLSkAkGvIFBkLurKmQh3YyNqcH9o5HchjkkO
vZfOCGI5sRlF1jW95RfU74pt82UPUuyYWh32t6yKDcMiaIhSvoAIjrY2sFMkIkK9U/GxkTaigpIu
XzZQVFI+BYJiRnV1cjCSgpOBicDzMyhQmqyJ3AGAuiF1Su6TgV2RFVkkTvrRdAoSzXvKnl5PzvHz
drrWyF8p2ipHeQAqpNgEhNPMJ3D29udPXz9sM6nQkisilPqpPDIPrM3FTP35aA1Chbn5JMS4+r1z
ncJzZhb45rc/54paevInN40aCYR388O9bh4ofXqimwCOSax4I7ckYd7bY9+M71WO87znBEcE8gZj
iaXiwlpUUuLi/qG6Ly6EA13m4alDP29lEZeMkkx6r4b0XrSXTQvTPxuz8dlQDAlsI/y2tiDb05wd
SCO3IdgniObHkV0uCCbOs/9BaBQ8tBhiBZ+h+r3dHMQBldBEGnPiOaScjg2lcoYT1UyWo6gdNbIH
kL4CcjhPU8Sw3ue2+vAAr7oaiRHEIpxvT8doIvAh12qqF5PhlJ51RGCs49hg2pxsqrUrEPi+OiYs
/uST/WSZu+bXNURRgmO5m1whCQvQh9BmD+plamIs7jUI1worQ3WweiusmPovahH5agCf2ZqLpnq3
pQuhWAQh7G10yUMQEArNzrbTijnm1hEUSotGsLIJJ5kTmvZYsAjQ3xWapl1ngtjxtN5GVOwwjq6s
sam9gMieyKq7Gw+fG3wKQflb9c8j+Hjw+9gH0eww5By54JS31ph9LYDDDWd+2NY7kVjMwIyH4X8X
EU02ygM1xS+kPbgU7lnmsdqLpXiZ66vkhrcAN7RRL7BB64y5BEw/gXBNTpW3MoPKG66UpEpLLSt9
iKEQhObLxU4EX1nDKxcRmIXAGlfr8jg0Qh3TpSM96IkYpXDsZwRFS7iO8Vu0iSYUs4QigZNJ4/U6
ylDH+fbsOTfG4U/QLhzRG9Pjws+vwH+WZlttC3rqKixct8Hkwa/QepExFxS9c55SwxmdOv3tbBwG
r/9VKrGBTB6MTjBCYRXxN4RUi2r/AFGAmTts3Bi1Lj15KYpcfmjPPlctzLrbBHfMiFksWiFNZi/a
Jk+IVnbYLopfc8XiYAejogIc6ZAxiGTfFUD9pig+BHjqqnzlMzryOHDSUVzrzTJoGcydwbZC5Vui
xmwXJQW3GDlh41sHA8PEWRZ2rUAxqOXeaITPHYlQTOwZd+8noKjhCTe8lG7W737iPhd/Cb6p+dlv
6pJ3r1P5VvdHYVV1K3w/inuxbewZ6uos2S0Wno0OAkaKmFo/iP0IkvAAcZfwcvK1QBm5+4whsK3Z
fqGoy4AIv7wK+Q7QIrABBvQW7FJNE32s2rmW/otnBVe1Pxhkr+zZ+yQqYBPhywijz19cqklqsGcM
AxzceRztxncCeuT9tc/zdyZMlDTrLG+WRtN2mfYZMCsEUfU2DVcmWndAvPwy6bHSbUxREGl3FY7n
N6W2EMRYmVe5J9Z9+PnrAeJ4vMBCgc6X8TwZDclUbUuPBXmLaSe4CBs9TydWn/i+LcmW2dlpWFqa
O+xakFIuKKoRLBabYa5HScjrk5AkLcGNDdklVtMU4xpzsPG+3a7YO87selRxFg10533FxEWE04O0
5aupun/8WYmKaRL45b3P6SZoCL2RTHLtIdVZxyqs33V9O0POEDdIEJUoGRMJw6qJRTLEnAYpOpq0
wnt/UM/7DmyxyAz8FYXjMKZqKgRLhHWIt61Ld6UaXCU3j2oakWqvGTC8FsCIQuiWnteKSZKP0927
alfGMHhsEgYcGunG3fejWV03VSUdsE2dRP71ZZv9OeG7QB2mhW0nHObHi9Gna59nnF0q/Oh7ZipO
sVmic+VareXVtLRT2cMuRnNTGvQi5uX/7hCxYFvenYiD8cOAU9DP2v/vKMCC1FjMyOloD6DRF9tw
rFzI8kQGxTUNeKT3ji5m/44aJR1KW9dWfG7/gL6VJLMCrXITdDTx9fGdFScNcnK3hnvef4M9C8zX
hHcKsuTinQE1u3C4T77OMf+BcQGx8IOW3XAmidrN126drR+ijTZj1ATwj8wKaM85wHiczeO1Kjf6
TDIH6+gKY3FScIKAjN+3KbiHw1v4C0ve/rN9AxUDXT0KnKs7qXJYfJqAM+rJ+YZM0+z/VBWeyAVY
NFrBBypUC8rThz3BW/EdCqejUgM1oBioPp21DpcnWuLBHk1bf/xWu1h5MQbsprQBUZtaV5KgUEqW
DR0CY+ygYMuK0n462nSOJ4XLEhEqXeusZJS4Oi/6eU24HvD5CNZ5eflf0pd1D2rc6RMsCYva9ATT
01Hu/Ro2HyXbJMGnZyNtmLp9TUygr2KEC82ppfeh8WPLJYKwNvLVfdcDVxCdlUF1hrA7q9PESJjB
6K3eEReFGj4JLrNhRE/yhp88pwpaHH7UQCDqwtVz3padlhOcAegWfPBVpeEi0l6LBRebUQhL5p0O
fYzp3o3UL3epTBiWfU+F9Amu8cPMa2+Ijc+aC6nyYUT0A6cveVExEdkYH+AyxUJIYppIGrzVY7iw
1XkEYzLgnMJZSffgvBNCvySHK/yd/Im7TJkKi+mRWcF51LxYxc5WqhVwHfclvxrMiK7XPlnjoC3B
9vBPQsBH+BnO9uiV2XCy7khxuraQ06wwMNmcox/rbIzzn7FeyDhvquT7YZPZCj7feBovFI2mPimU
DD0QZVrR+ZJ1TY59uW6QQu+RXEsUsKQWGiXXyOXe33lCmHxoN+WXYBIMhr3wCtyflDYgnBzSB5rY
iqjc1+mL2rRVt/v0e3mEq8XVN6jAYV1g4o0FyoE0seYTiEP5ACqbMfPS1kWfqsjDnrCUCUyPlCny
b5Xj+cRs7GbMcFz9ydN2R+ejMj+YnK9n89BxIvuuNywaG7Iq1bfLeoqEYcBVO0aTVBrKwSO8VL7t
+sPdmoELdtCDwpPWcTiMN63qKx7fmqHHhii+Ico+JLQUOrA9PObddzJp2ekJoudxVh44LVR0myyb
ohNiH9O30ElXc3QbLcDeaVjI8nYt1VWAsGbAEzgB0dogY+12YEf/n0Y8xGLFqwAmhGswf0B9Beda
GI94aExn25e+aozun8WKDs97917ZlnQZ6jWJbBbbbzSKYDPF0LRkNK0h+3iUiLKp8qPYWWG3BXtG
7JTWKRRCkh3tT+e001jaCB8hFWq1Nwcq1l24zljD2kxyyt4Ra15bB3X7NbEQ3x2apMIsTtdGr9UW
Gn2vy/K9YFwE5wA14tDClwQ6eLD5Gd8Kyfjvc9HHNiCaxRyqYyDVPOtXil1kwpYocovGWyk/In5A
CpXHbPwTn6DbgVWKorDd9jVaIr1SE8q9vGRdtLwMhhvzNTivIGbNJGExppsqJChRflieVqpVUD8J
xno1+iAQcrqxy+IvJkeaszYr8UOl30CFoZR3TyR2MezUNtqUe+bffhPXhes/e+9JObR1nUVtu3Hq
Yd+Gsiw7y+vSNvXGgDQtFu2cnjQe9/DztyAuBWUobVdxWlHoArKbD2Y5K8jFDT6A0cemsAWv2hxd
nezH/jWVKFAgnnIXZmpUrau3OV3PeQRJi6Xt8A3W7nYX2lzeekib76G8ID/fXTtjC355BXtZ6zwY
rCV2EdELW7latOJcghoKsyxv68W8yl2BYiKU06/8VM/Mp+BUvHEiw2XZzjJqEFRqa52ncCeY3ZdF
kS6XF95M+GZ5wk+INfMndZGnPmciNvKLq+xS18uek5qlQ2xDnXth7hRMVdywtWWLlk63JSuMIk3u
GavLQH3Tli7XeKnZD/RULeHsUliFTNI6E2mt8FlPUpl+PJdAD6SvbCHrhShn+tSIVBvCzchcj1fz
LtXsD7KGaigzWfJXlVngfKrQCMXg6mzmqMqgT6yJdzZ9rAGbeY7Pm5LauhbOhdsxzqvjKFWPTR+M
elmIsfi47SWcE3VEU5DjFcfspEfrUaWo84UlwdkP69O4PE4UvBmAm7VaEXJ7EtLFXMfpPyrSjUMG
wusF98AkuqlUSg5P4mlkNMTFhTGenPheckbH3TJ0FKAW+nkkBvIDzH7bNU+CJ1iJQQ9ZNh0xRUZL
GuNOTbAFG7V0tmQbzv4FkVgsOvJJxocWIwC0a/YTZpl+QS6m6+3hNpwQqSxmJSCh8gBzZGiNDDys
7T2joH6kX49J6wD/yGcsOB2cYauMm8P2mCc6YoOcxB6lii+51rWg7UB59eZmJGv4gmCs1K+6iwpi
4fg4/0DOhv3anQzLVwY+FOs7WPCxbzy5wzn1cW6yMqU2gtdIhbpWOVr8uz6tOzsmVSMthZFn6apj
1SHNaSxtuRtq+AXH20Wzdup+TYaAFiYrwtjc8nSlVAqZtsi2Cv6N2NxcHV7wAWVJCBDFQ8kuFeUn
CkQjmeIk1gZen4n3s3hBcWMVCYYL4VuI+J/H1Sj75ywwOt4tCq9aBiirSyFNAcEH5LrFvdRjosYZ
9jN8msLbqsNa2FhB1UqBsvFCPzkHk2ftZrtcxhwLjul51EkeBg7L+9clgZ5lPdEtyKgaw8bXFuSo
A5lqEkxg4uqhx15w7TmZH1I9bZq0UTgXSrMSS6I5B/j4QhEf6F8FoJckxx/NfDSfDzwZlNMzdPmy
EyfKHbY9k4CoRjTg4Oya4p3cZm64IFDZhVdQER7kSp36ZzpbEy/+KXTWmBqrOEkeHdyyv4QpmYAC
XJxFx35Om5lEQiVNQTjwccyNu7w/M1soRsiC7Ls6i80M7FjwBzx77RDF15US6APT5pYRny9M8C82
V55/sgOqPFk24FpCirN36GYsbs7xpxlJioiAQqGpEn8pHZSMUjO+n28YHRDJp3AVwWagLUV7p1u7
XhNVzL/bWcVhvo1R5yzUIodgC0HLYJODOueDKQqkKI6FBpz08xFXRoog2bPGBSn/b9DWZrmgDBId
DDNntJZwZYDBfeK+IkIagCOv1tgc4aBRfTF4OeCeO4EAA9VtgaP+B2r1nHtkt4/mhBSzErJMw/t5
/f6zjmQJkeNkjnM3axeVPi2abpKjDsO5r4CzDbu3aENSHVxhYkT8oZq3YjKnrQfrifjRHIQzNDee
BY94AwJL37g7/hhwZXijFIFD93IiJtp7QIaVMZl6lPlHi0ObybLMlZ87FzgFKzZbZyfoJZo3dppL
m+LhEyHHyP9E0aJisIOVw+IaX1dWzTZvhhVHsWQbfssX0orB04as63ha0H4cRX3dD6JnMxayRKG1
O80lWCdDN3prlAZeKZSTOA3Vk53JQi7Se2Ozu0cJeT9ceiMJrrAUfkC+MnSPekE3PvPZ6EyAyUeo
6L+C2YSL0a2XdDa70Ko1ph+lwUXwWDkSqHay00w8FNfhNRsxMnokoXcrCG4kf3J9RaGKblrZkwc8
FbgA++hze2zDxMfLiBNIxJWxgnRpi/mIsPFtkDUbxvMHlwrjTfu5xf5Pofgbd0OznW0xe/Fqpa7x
mhzgJGFuB/WZtANCpErmdQBoQSvOfk4atZANUx1WxuiM6N8W8AYipcY6VsKRon8GNghGAZoTxuvi
AzUvMfNERJboQrkFaSD1NdLbFzZ6sL6pUzhlT9MCbe9CLtxRqmhTlAn6sMhEncwILggwB3eYKqqM
4uLDcxyMD/p2YVWb+EAHL4MI7U/Tbx19/Hfu1/rtcK50ZPSntEb9G6vd1shYPqimAi4UvdTxCWu+
2ubJph1w04iIriFiaX1jcc7GdpL11Wh8vQGcKPKsA58SJjh/sw0r/ECRT7j2sMTfBGwKP1G/Y9lF
dJDZNkpyq9vlwb81rb4V/FuV2utTLAFvm7jTfyLMDfq8JUKBRkKBGAbr83y8ajeydeCn5vO/b/jU
HM7M+4kP4ex06/c6eaqIvDtASMLRRl1IYm1kgQKWGvOZugmYLX/akyVjz14FNBxktB3AVfMmMiMp
TXJ6MDm6I+TSDh+vrmFZSSqLEWeAHR7vJtXrUK0OzVSl0oMJzsF7SVhu33myrCgdmI/l4iABg4A5
2w8djV/hotdDG/dfBpiouKceZ3l5Ezc0qC06fV0USCtg0a7cFCC9W68Yw4dj/NHlPsR3rKQVEZ6J
J4XnR6TkUQ2WCQi7opAsaxruXSTiex8phuoO0RWyHwP8jDDtZvbQJAeREBzRJMdNlezzarwAfIoO
Y1f3VIK8Z/rv266zOrka3i+B/MMdV3kK8ZASM9G8s9zpmu09KQjraJIh8oRbGtxPJ6Msjerv/RNQ
4nfGnV9S5+gWcAmjVuHQQwooQA+8jEqNIhKH4sl3ExUXr4QydkLCzO36lFn6+ldDb8Preg/7nr0P
nZ5ZRCIB7vLZxqs5ExprQJiPVsfepKcgR9uYNMJKja73KRoWjhccictLiKwpF+b6BgZWaXFEm13D
KwCgwk2F/4Wpz/HQI9KJsUgZ866Afg/y3UWItUz+zumB5aOzkxqK+MCcYnPHHiPPnwaSqxN/zM0j
vGS+SrySgN7q34KfKX8owxTixLjybz5aJb9UNmyGhR8sB4S8Gk4MxkBZAxf6qlNpPPq0fa3z8Wrv
Z4NuahjQM1Anz9gYUGljMxTkqUg0qv+FfSvlPCZNs2DUSL3cJrrQ5GVyPKpI8aqjaYmGZfCX7p99
WFrz/2QovEsLmjyX3bpcwfGjbIW4QLD3xLqBT9tpiygAeOruHvjGTl40D92fkvBYg27quGtWS+jw
Ui74rKbtYn9ruLU+cSkOdDG+Zlh7Gv557E7j2XtpjsR1DeaNv+8C6YlkagfqWW5iJ+KwY3dN0Eas
Qb+ELryMbS9J7gpdX8+3BFdhsDj1/NLv1lH+SBo+UlEIFOj+r3msuopKJdA95xuq1icglskW3xY2
CIIcZWdsvGAdT20LL8DQbyrm8DxjZE2acaIyXB/elakadLBjxVBH7yPiz1IrsR3LOqoceambk7E6
T60FmZvi4D/TSIrTW8pf6r1OgQ5Koifc/II0Zc6KxCn11HOuXXrqp8P1BHdr3cyAOCB9noOvqBjV
AUz2WVG7157Y/h8cN0I9/7UrQ8OYxg19+uIZSSGaOynuBv/rTnubkFsOZh79D3Abi2Zhhobk+LwC
rqPvv06gEN0TkN30CwG4WtVi+2Ew8CfiU+8AT7JpO6Q5qFgbcxWKWp7O8h6ikkaNLwuwKYb2cp0k
9+yYHXsxYpu569jXOOyoox3ptWccRdZiOpaNNxunME+bQTlJSlENKu6DGRH3ag15aUhmmtzPGa9A
D7ZPXX85Emo7W2o1eTjkMdXWGS2jQt9DnduL5AcrH5HWsRYvjxM4K4Gdx4zoO5YAfu6ZorVLRijH
ZnhbBG4meBC458/hHLf0bL2kkzdvNd6V1LMgOtXMSITIPsMsbJP4koDFQfqZ+7L35aax/cDzOmoU
/CvI6lhEGmQesgB/pQOZKXVyA+7dyXxnlx8xp9CjEcuERN4Uz3sxmHeqHV+taTIb/2TLNGofAZmu
TyygF6FdYFrsL7ft+t26AaoYG1rdyO2ryq1PYchR/b7B+n9gfoR3V8d8Qr1Y3tAcUFxD6MOT7C/0
UJ30PqVTjaOeo1P0xVETDTs3bbMeLAaB91u+QfFxKniFm8ZReq3hLR0yVagvNEsCb6AcbxaQUclu
Ct38Zlay473i83xF5fZKPw2EfLolXbGtr2RxbJexPeo4gOPHtlCugXFjDRF7QxgR6MRZqCGerINy
Y5VUV/xmqP0b1QfRY2aQzKK5nLjrHgchjWYYpKfMgZIoZyxMVT89Bk9xthIYWYyKdaENiZtbaVE/
5Sbu1TnDZdYgsqG/Xh+9wxM/C4oAu6axN0OkOVHL1KM7BsIWlNDV9ayirh1sjLUcSmKvSv1ATSc+
ZWUsY4xXM47RKjWYHfrW7maZLN2lsAoH/Ox5tj32T/VDuOr+NfpV/m5nm37EOtXG59qvgrEIrH1s
IUrhhNBhkwaqcacxfO+aum4W+fMo0iitBKSLoynBYqajYyunvg2MaHhrDLvI2Oos75Wu5fATLkj+
u9sC6V3MzJUs3V6BawDiYNE2GErrRvHOZAlSgKlm0aCwvc8+/2SyvddRj2IgZ6iwRnrqAAHvIAYq
hCPXN3w5vxfHQjTQolfVDpkbAeJd4nQN7BQ6SEYdyy4eQCnKk1ssc+eEx9OI3mzZ5eWBXpm56hZo
w1o+BymIq5FPgC2d3/2vdwS3RHMgLhZlyDFOylTs4WEsFZ+HLVaqwXd5xOabNQG2VusTJw//KzYi
IoXIoTX/YyF1/DP8gn1sVfb5WO23JiRjQiJB8mRci4GUs3nPOoa+Nc0w6jZEnVbzIvj4vlU8NXbl
xi+ge6ICcYRiIQtDJpiCUtNJouY2+spW6Edz205W3qcMEmwc26wP5rmUkFJyJ23ZbvugHti5gDQy
PvdWlwYmTQ+TTgBFhPknXciDs6Wts0z0hTr/MOZPSfsVT0NWG8gRDhICUdHS6Sj3W4URznoTLOHm
bjR9NhdRyLJG9AFU1ePB2BLlOfh27tU6tYthRSRtL0s3WtXb0uVfOtO0IUjW2tjurWL0FAOiO/LU
dQJX6iauv8HaGqRJN8M++xKGERCqYNP0vmZ3GtgGHE3nwti9mFphyj7Hc8uz4ivfAoYiaex6EXr5
K+xkym7BtivHyEfZ0sE4VWKzJnJKyCo2vYNor5QRvelEN0iyLTCt6PnGXQv+p5a/hgpRkIW05y9M
laBrpuR33K86tNRpiuk5VAbOXaWp9flnJtKdFwzDluDObqFTGwzruUBYhw+YjbSQboZWMXxurjj4
pffSKkGeLis1n71VIkfhNzMBE+Pqkch9eihYHCn+Eeew3z/BpTSKzVClkVROR/ZJBJtjYiocS6hM
VlJ+ltjTMZN+NEX1Nnq3KMggck5WaQP24t0KInF2HVIMdiMP+UaaCEHHLLUb9g8lNlD+LviSnkph
uagwtHO7mpmUIHNvfcptNB2ZDURb9A3aP3C+AW2X2Y01zopsc0jJGN8M8MYCAL17+MRdhes+jsBh
xj0D6Usf9p4d3OV1FfKGl/5oI/53246SaEtVo2Trc4GX05u88JEIsi4wBRjTvRA/VKFFEy2MhbkJ
31B8XwHv0BKln8zqPzNT2ejSWuEj1PQ/fjtO+A+cPp2PPRgu9edo7ayZO9t9YpuhI4DD3kPLXLWv
RShBoEEVJfHWQ7Y7whPV8w4ckMbBess51H47FhPUI2Fqo4Oov7hFfByZVvtprAU79IhEjbZPUnZ3
cimnK8IjG3XpnWlnzaI9AzUTbNMf5kHpdBf8YNk6el/Jky2mfTZIaqJeA3sDbykD4Vs8we2WLJxv
PMY+ihCCtHRRMgRzv1mHV1u4u0cCzqP65uSY8nT7JuQKoPVYL8MxYHKAd9drRry6ndNPP843M287
FrlxYkVhynIh7gqtB+1EAN6I6kmpJv7Or8cKRcPjEoHO8i5WZNesnNwylewnUj5Xx+c+BVws8t8P
lyOOtwZs1oUeO6xq3X9N0z+tlbWHUgld4hXXI8ehiQzwMMyQVTOFUEEyk6SUhUlT3GWdozazqVe5
N+Rh/9YuUzopuGksYUZcraPOokoajydU8KMO7UXfrbYkl3aNFgahmMVWQg6khY37Sz+WH1u10tjm
Hpg8GVukR4YG1QTM64mGQJVfuqoGjommP8DdOIriTLYI8KKiN19KArcPuEkRD8hMj2xvFQXedghi
oQyG7J4vNpGkcryuUnuqZIXjmKpusOvIwoUyP1KS+AdSSJ8P4EFyMZlhxe29SCnru6jnhFsN2Zyk
W2tLhsIDZ0efqyl+RkhIE6GF5zP3flz9j0Bg8s5tkbGSJ78mesaD4Z0EelxyRFRnCraJUzO6iJpP
MsYXd6nBh+HzhuieUFuuGgUrcp/BjumaibmCXnflYjoZtucpknai/o1SvH2Bk+6c0d6+cJKw8GVK
WLeeMIWyd1MHi0nNQl+q+vzQR08DlDk1CFFn0cvcJd3CBtt09KMqX2rRTjMu204yrtLh5OHtwIft
j/ZrJCIea0YD28JvdcxYdKpFomZNVEV56nvjmHUvRK+YB/zA1un4TZCUms8QWzdSAQZhm+TpmnEZ
uw7y2mJlmHFCvKH3WeTOINTrjmLyzQM7nliM8OnUI+56aw3WAEGAFEkGn4o8oaYHfTHDNJuG7XNH
DACPyVtXlA3iA5cFXCV+Uqmqm4PPfwYKHe4hx835tfN8bg5ZTdYbWGDeK0aHIBZzUlsA2KLr27OC
7Xb8RCYqzpb2gaUKCB4nNqCNG91BDybFAPyvNrjBTC5ZcfM4UKxW6EufCs4bRWdzctFMl9DPgEc1
PjwpMs5GhCsNcGuys+gwZWnq7xXqW3Zp9b4GdR0gKhxU/KOqenLb5Nw4PYf42ojHmFtWP6WYYGtq
B2BAftsSgMdZnJR3zl8xVq8hpivY8ymunzTnWluW8KMF2nv2z8eAOpjc+d9yA7u+ZIYlBuF0Ov2B
l8mwIXdFry6DWoxjSzOJMmBkPYX7eI4mvnWDGKlBWmliKtnYOtV9SKaqFY3GLLLPQzwcqm19YNfh
Sc1rxhMNqTGpES2qs3cJbAqxvAZlomXtRXXsg3G9pxiSwUFJTTjuPP0ZzC9jIGwJqQfbWebDisqE
oTUV5qkxj1o4aQlPrhczM1UeX0Lq3Hqw1gWIrzmF+oIoC64NYN5N0IFo4LQQa1I6FN/sqv0PyvRA
rEzPsIBomRFpC9aocDlAii5L59oA/9sTJROc4usOtFfHoGA56fXXgTAX5OLJ4KGo4+lORSA1/1pn
AAxgtZw7JeEP7apOLrC3ClLzEED/XOI8wxgfg48Rldf2JgX7N+X7ZQS4gr+PVSugkRQdMPwD372O
/1jzOx3mWPgsAhaQ8/jn1of6twoJS/KrfBwDxf7orMw65g8TwRnW7bcZhyOw44byQyUf+nGoApIY
ja5iGpB7FQaqlGBhK3J2BvTdQPZNi3310e3DOfsR2LsODxqSQqTE5mYT+6Jt2avrZ88RFunWHrX9
XTYzjfS0/MZpTlmOVWNko2TAAph6fXFM1iTbLhVNOAPc8ukp/jigKEJZqTE7ChC33dyEhUi/Lcqj
eyOGC8ITif8LXR0zVVzZUa20RkDAle5F5X2ut8oBPCn7q2a02WcTAXfeETvU0Z9zonJcYE/6AtbM
Zn2ph8ZN1sOyn9LG30AuFK2EvE6Z/jI+R058vcYVyjtD6EYIhFbzotpzdNmJqB9HGHGIQcTXZFrd
pnP8bqXjXTgmrgMTBDI38O3CnJy58E6RzUnn8A719GFfMQ2OgUJYBcJgcXJj3RCxZ4WWhmYSm5NZ
AI4Wb57rKB3PH0FF+g8TVzpd1RYqrciTyaUJi7/W0FArd6WB9jkheq1uhRtJmUj7XDp9LYzqBkYt
b4BH7OPz4fjvu3T5vfB5g87IMI9w8w9uK3DGgYW+IBEQrcM673OXujsrXUDg+JGMRZHxJ4MYEIrT
1gMp7qEdm8G/DrX0igZy9nu1ezKWc2f2NT/RGlxctPq35NcuakbInU1Uv7ZDZzvRAQl0kywqHiTc
LIZsZYgThHOYozrTfVVlrjcDdFqGXeyD0QPz6XIbxbZ2FquOZNDjA+LZN70xe6q2AWYoPgI2veiM
wIWnNsZe7aSEvVG7uc6TyiskvxDLS30b2IS/SB4GGs+rxYwSsYAK7HS5D9oo65Oi66k4kzBQ9I1A
zrFqUIvURjvhK4xoaIfqVE9yGFnA8G1I85jHkiagktCB4foXiDOM2HyZhRMB7Dl4vFiM6NPiA1cM
2U9llP5qDGUsk2PqQbDGNieGg1c/XiXhCi1CgLQiIYEwNC+l+1WdMOTR3HswZLODXh5GsqJbk8ic
XB5ltrp5rcKQvcTAY/iNUWTmqZuPrFCgW8/sV2dT/G6vKps6v01n7k6O6AwC5pG2zuOgzGIXpHYl
/qfd3cBJg4PIx/E0MxpktPApoSXTyuwFcOx/AHcCdEAwkBMtAFXzZXcOXBW7mI5Lzny8cGiJxjLd
1bB+dow/UaYB5vFWYmdt1MkYQ9enzw35wUy+UAuCnQQUX3wtYixjf2OGMWs6P2aWgSSljabpSqbJ
Crdo9rCFARvabLOZJnPiTh+4vp4rqEsGVkBJvD4ezojk8vIS9vEAhrsxOjGRHtw0NMfRoHJY3ESZ
hD0KyCzFeSg2As9yOT9QnuOiHhLiIExSrZ+Y3MRG6OQExeNrtIKaBc77RD9nhKPVIxgrKGZ1H7UE
ZH8/beyHc3X8os9+Mj3m5y+1ZlsIy2ytrvJzLj1xMXbltlJrtqwMgM9cDorkUxWVXTpz3Cg54aou
hY5pu5fFLC2boBMQYnz95FqhvAAU/G+sz5xW+p1offW8sYCHeOnYqF0BjtwxQX/ZoNuhLBT6oZLI
V3h6Ne8Wf1PIDcILjwDXhxVPEA7bZfBvyHq0q9rKrjgMF0V/UkINXUIs87AYy3IgLxB5tCFYeboo
m87rQpLMiZmKv2/C7FOqmVTa5/k2LObrswq7g1UyQx7mzNlttwOOTq+ktgG+vebhTMuQZpThdXZu
DBWum+qaDKIIiGQ23SNNuscMQWRACNaWNYWlODilcFAqSKtBH62tCyAtbilnrscjWFsquHHlG1L0
DlfZkTh1KAfVhupCYJnMEkBMACxg2JmFXyzB3ee6l5/u9svQfNHfGo11s7ODfAb9a9pZnEpCjNOM
Nm4n4OGiybOdaJJbMEcKJs7i6Zh1OVcJ4VUjwAXgqqDZ4niYv44h678Sh+Uy5Eb+KrshY0l88gzv
vXroDd2SaXrFLUGtOS35uHnToPR63rHbrSsHMHHnpILPqzrV8MCJoZmveWAkJyrLn2X7q5b5cH1K
5g03GIJs0OfaYVyfsbu1rAniR8CRxVH1GnFtCnMmZhJ8fejE3CS+dXPCXBOkNuaXOf4466MZRxYY
XjAUIagajUWk3fCS5Sl5VuieAZNgYnQw96GePOu/GkxrDLbXMTA32TS50qZaHmR16H3OGecSoQ6o
etsMXRbDyC57ONJ4+ZgwPuUay+0zsPt0t+OGN+HKMSLgAaTGaoycD5vcV/jxlAMgbQ5DhrXxeg1O
lutu/yKH4Z7g/qEOZxoWdx8VWRDOU4DX5r1WJPmVzSD9z7cqS0IhmeqbXceakVgSbo/iPsATnch9
Se3aBbAllZWyfeBmCos+YdS1+I6FybaJ7ed0FDRGvC9IjoAU+9TXHwpDHerHXIwAZ2XHWsqdInrN
cVHsqlcAHcDhi7RybZLFteh0KeJ5sXoslxuTRwqcJUeAX5/KewFOwebi/yW0T0SIiHgmbl9/glUF
4XmBjPvsZzw8CWt+xKy/MPcwn6tz/2R0Z1hfuLpOojkWedbM2q5Cc8Zy4C2udtavFNieZs8h/tBw
6VheR9917Wl105EwrKB/hgssMLMim2cBrOrexF1r106mn+GqXoEUKOcrlq9XwLJVADfGlh4OosOM
1CKVNiuPHmOurpPJpTlYsNOjkbFMcGSjSvY8pmBdLKLVqL8sEjBGEFtCu5TYatqSUoe0u25T9YEs
JKhodSsQeb1/CVT+Pv5My+c2DNKoUqfRDGM1m8xjvZ+aOGVDwZBHnnRB/77U8xyCfyosOrYb6+rj
xipVDhi3Ei2GHQLtjb416CzWytXBTVV2onXZw7QNFVMUIDqUtv2T/x0fzsjlg8x901i/GjM0nTNY
RTgKUqabK2Am8YPg19GMuh8ndhOiJZuibaC1p4cl0Qz8gaaIuRKP+QuHEhPg8DWC2wrVcr95lPVN
Qa2Rdnb33qm7HIw5DFvSBw0VNzi2q0MJaaJeK/EA1XO2cK7p9AHOHOl07KRnVIz1KBXtvxNgKYhR
FYhIIR5ODl3aKLwD3OvaS7j8AUam39AFi5sHJ8VdWJKCyofY4gylVMvkRfSd6aEVTV7SlcHKFqDM
OxTntxbbdukRTHmUKq4MkaWqY5jgPv+3BsB+baTH2CZdLm/Nb2cXrqfFGj+xEdYRfRkBWZ4K80Nn
2KTLai8mOU1lsuUoofxgQDjBlIImimDhuKr9u/XX6doxoUctPPY+9gtwjsh3VEMGdskj8bMnWW6M
XLPqm05uKrSmYPhyaQRW/GpA0W934yKNbUql73gq8wPQd1ML0FfStcuC3fU6CcwLbTjNey0TPz07
6So5LjK0u0hl+Iw482DLxyRvs3j5JEb90rBW1DUmfcCgRXUNWb5wYfNDg6fCCINrXk9YTweJ8rSE
Ykjk3bk+gu6TWpAtjkCUIwteW8l+/9qi7mHDCkQdVI3Cwcs4XEAa5OzQyUo2LWOgxNARk+Jpyqab
UnZjYO4LkDHA+9y+qD/o+nnQRX1kmqnCyx0y7fJtxusf2nfDssCfqxzoSOdAlMFdfQSI1Zi+PA+d
7NJFfWlqSTTxft7I12T2W3WyHSzoqonbosxo7Yfxj7e6tqZ0/acha61PF7CxAQ6KJcBJFN3QJTbP
Y3XRSeYTzdQknRcpL+fESv24M0ann8n761tYBCCQxvHSAh5dqyESxs1TygVWGyqP9EvYjMajqQ8n
jDLE05sB81O/XYfaNEY5GtrbtkNMBIfLX3XsslqZ6cZcw+7DfiGlr1wiQBhRZtM0n85u9aIAhUBm
WbDo4dqIDIbdDR3CCNCvV+/S2HHEjOAs9/2rYVbfCPJFucGskkzQpKC5Ln308RigtoFCokFey57j
pVjhxE4G7M5WplQn3RSIV8neEcfEpKTM93k9dmEyxHVIvpvuyK79AxPMhAaVieSAyKotzZrasiyp
FKT1+Up9PmfNqwtpcWKEt/TNQes4q2b/mNUkEUGdcf6YEI/HVDqDhVhty3lGTSN5qJ8jT2ybhEaY
0wsG3vAFzDwO6fuFCFD04+IgC4CPYvx2VuExI2cMdMceodIrjp1wmHkgdh0kZLm4rhB89NZhign2
rIEiFxHGatTq3S9jdzV/SEz8lCN8ZYxIZZwXkAAEnplEuj+sz+4qQrUsH7QNrxhH5GgslXwhfUXg
atSjCaqvcu/vDDFI+VSv4Iv8lPMd+aOqwMRXbLIDiv57sbTCjKDt2scbvcghOjiUPszKKkbhziXY
Ief28Jkn81JhoyTpL/exYshRGgwUkIo++x0pnYyLHyU7U6YAEtjbeu666rHugUdtdB8dyfHd037M
uld7HHjC/Xoe5xlQafyH1WarpPRP+5J6T6OHw/hDXg3/GYX4NUa5QHrU/sHAQ15YRAC7p2BiwayC
fMSzZaP5QIAnJtJF2d7UuQbO4J2DgZfoXhK9BdKiq+eCF2oPcp5FzjR7SVo2GPBcpdNqBzIbDspo
5Ydu5h4M87phhqcZy8mMd/4NlnyHouEPpPm8+bdvD0WsKhcdVf/lp2b1DwdN91+/CUlcS4zsSl8c
M2lEFzxkt2lEgf4mxdtEMo2MuNHa+WsnWhDxS9BXod2wO4K5Oc6qsiliBQlggZQC8Zwb5pAQRtDM
wptfu7JtZ4kCUHUDR06xpATOjogguZf0LWyMtAuseY43/q83XxbvcKghSHx2qwK15UnFDPeYvzM8
shGWUYqrFBeedecrckyaAxecPXPwJQLtoryVmUgZewBDwjRhGBa94zVKChxu7fkVpr1c4aPf3FFC
k0ULX5U8Lc4MyCqIngQjY8C/Ne1EyC8X5FsdKqZGnTmd0B0QOGOnxb0bgllB9/b0m4E2SSGMhpeX
nCLK2vlWI9g0a2SwyBWGyOD3a5n2O4nuSHRkZVtlm4y3jqB2J642VnFV+qIaXWRhdeyP+gPBa7SB
Fo75Ni3S4jMPUx5v+qMj8+F/+qTtCrVCPGDqGUB2pLHLigQGX00W8l69Ekkifpzc6ldyyT9Y5xRR
dS1kCQpnjIA8fwcmt8KpAkASTswjEP5WQhw3mCmQ0xsY59Q9AyUhVVFiPKcFPOw9gQRxnAHmwMtF
G3Y/oabaSGQv6POZp46p+Xu+5cYKRpAnj7VLEdyNETNGkWoIf9hYX8LArUgi4jcZf+TTe1lzmG3z
RQJr7GTNbsJsnLyQ6zFjVkjJuGk/oHVQYmp+ZjaXOW/FYEhpON5uAsSKqrk/TUtFECf+rOYqXxRw
Y4WUvg0w16nbgjVQZUsrrW2OJtzDao1ZiFIEbrPeNK5EquAJmGc/dbKz3bc47TqXgtqYCCTjhIEJ
5OP1WFkO0kbEo2Q7BjD9aRhJN4G9rakaHob13LDWiw/zW86/wONNUfstFsuDrFmTF3rewMV/q8vZ
ViWVpozkPjocC+pNM/pmO7S0ZlSaCcKXYd41iSaqxmM8FX8xHVhLUwWTtlNa8Sj6FxKCnG02mS/S
L1uIc1E1EfCEjq0FrbARKLxe6mnlFBIEWAe+rQ9/sFwzvx1IZzBqF3TIUH4mdrAgeobhoKzAMRPQ
x4kOJre6fxQQxeeDxRUOiwDJpdTkWw3zCMLpWg7zx7neh8o5Im5u/AExbEHX4gbG113kX0MUwOI/
OkLf5ey39FIB1WpawJqaI9RAlStGZNRpM0wciVuxF/0U1JF0/bz5XscVM9Zd/EnCwQcurSkNIuzS
lTYflIZtAcH+Pslx6cOBLdBSq+8mnEJt88OJeWa8hGvUQONuM8n4R/pB/DEnuSB3laku2G61a5OH
XgQCwn5jIEfKUBTV9t3ARANF4Hi1KAv3mhFiWvqHHImp85pNXuEJWqLevokQQun9JqkIKtT0Lzk9
3xvn6bvjKL7MLnFyyTpVYz2CwxhG5cAd8NT+bJNT7vRYL8e5J86lme+Eyg/DCjHPUZyZLf7W8tVb
i6aTJqG6gX33zqwNZpe4yFHyltgCqujAvv/BJ8oryYBVQkD7UA7xcKmHcuWUNZtSJeT4AAVkSJRW
yQkPPITXQDviun4NNgbx3xX2RT3ChoKMq7etfETbaRHZJLPBY7MrWksbWy2KQ2VFYVpwVLun909q
A14X0kz1WYE5RAHAj+FsDfVSPzzTmg1LK1dva4kSO0SzV4vHRsdM0BIpo4UZXJNRUlISTq1IQ25B
/VdOGdng8nLhwLUQrmxPmqfPIQGUqMFk9GiQd+dKdgpYlwV5vB9a5d3jJWbm5GauKyCSJ8T4X5OZ
778rCIhZSGvWk3cHGGvuYRlz96qJL1KFbPfTv9W9LDVe8ZWpVeYydfviavdzhJXvmoJW0G5VA/PM
bUoVFmW6CsbjwpTmhGfX9jV9ASVuB1i2+Bu0+/234hO2KMGbTuAxPGGfJVhf0GAcT3QiqqEEL+3g
CBKRA2onElYYgjs7AjZgVoaL2zhk0ULQVKIe2VBdiBhD3NopQlOHAJIXvQdu04sFFXF3DccBAtWj
pz2oTSW1OEAKgi5+PLYgwc2WwL/EPfBCOMCegCpczm0e5hO20bV8+M19pO9TvLD0S5/gSr1AWz33
bMCnG46B4Iay9KjKXMfMRAt1cSzExW/CNg3Jd3r0DRbXFDMkfZYenaoVvSc9XiBlCF+PgK7mi9qs
mW5Rn0s6Q6DOKWqIKucpb+Hi86+9FVY0iiTQWS+H+sJ1rQv7ngQ1AfspMzxyULj7lHLDyZaUzsUf
BwNs/RI8Co02GgHlAtDv455anHph2FMCkDATgcZXrGbMtG40/Mxhl6EtI8zbF7n+DeN0hGAahuYi
Lbn0+lhBj+f606PQ2nkuP996n9RCOU3xBDLYakU3iSyRLjT0YLhr1b2f9YGfiYJTFMZUMeovuJCy
BhmY5bcVZVGU2E2xXD7mt9MY9uJPJKmzZqwlD/OKm5bUwrFSEH4gBcf48XhvU2vG8+0h7U7Iu+Cb
8Xpm+zWnNNVRquMED0sobdhExnC+eq54A9DmAe6ZnQvqUzZiBbdHPBU9v4iT3cv6WuGZW0bSBDjk
3t/SAzQb5PDQ4d4GuSYvXOenfLQWTYMMzq+ydMhVXNZOJkxcXuzu5/IsgtCdwXecySsgZ0tq7m9o
Wi5eYm8014hKGiB7mEG+nipIqVXgtJi6W5jRh4MgP3601bF0IB7fmP1dXzS/U1luQmLtt2oBy/+F
GOWEbyXWaqStHKHtyPAaRVnaJetzer59bXiPmAw0/ydtsMyjKmK+JLkdDWNW8mRj+E5p9HuktnbL
t/OOCzbkGBjojsWsgJrZd2YKOY5TFwQbs0nocSsItOInNeMGeFWnfQlOd8Zm4CufU79YdZZ0jxqj
1vk0E3ENdKY1zoqRcE6OWqfOMoKccyC5X8oJQ04VMgtu8CBMkocXQSWhoA3+89wbQDRC4cydVC7G
Yh6ffxmDC+09VHcZvxFNRFSfTnI0aOnxMLwxfh2+eBcQFf3nPxlXQq5OuYJgOOBO/mUWIWQEpyGi
kRYLQ4kSuJkWKnli4HXm+Bf+E0H0uXu16cTPWvs8X2co2+UAQMQ/xsjg9mZRRuQzuVlKLJaG9lca
xGaq/bdXE/37gC/znzwUqkQ4IAlAykqPNuqEYwiFFu5RLrYcanN4v5DWQg0zpUh/I9KtWLU1/EeW
A2mblkREWp/69RPHsgm17W6XLfV9AbkiUCu675wznHlAJqmnCpfv+kzvZ6sFP+1+K7xY5uwTJ6tc
iKZX5C2/6tKfBzyM0GJQ+Pac2FeljfIndTamVaW/NjaM3vK9h+XHwKIjKjwPqzy+RZgm0WHASLfR
ovPKq6e27vnbx4eOf1nAReZlzESDp69rBtPNddMT5nXJYDTpL/b+H7/WajGJchNVxu1Ym4fmOVa9
kBRh+h5+mnEdKuhW163G8FbBmaFmk5DWs1Agz/5FoxGdqlzYYGG/OHaOE1+GweD8SgaVf/7wFki6
vnd8qkMpkVR2E+j+jzrbT2Wu4I3KXDmKAnB9Ni+3L3oCu0qFexAbO33G0vMp+Id8NmQtzKTMHMhl
C7BKjrjVpSqVmt6dV9pZtqix3dF4ilqlZ7DKgsG0Q0hzsRBHcc+EcBaramUzjWHIFIzVHCEBNByF
QgqDhc1kyjdslnNYlPr89oGW6vYFZzQtptQhG2Ff7Uo+WgKzPwmjWSOtrVmItBf037f26gCyCDaV
ZqsfcMZDnKnK5jB5Z7uNYSTW+UuwpoT6oUn39mKg4WDMeHXjl499wysi3ssIYJxqJtGOkkd9KxNS
EZe7w9Tln+wwFyhPC1CGy1AxEnIvJ2DQb3YgO7+nPtLr87qiiT/j2W49rSMIsUYI+ibOB68ddmHE
hN+O+HUZZsLLoEbTBTJCXfUMHODjTvLUQ2qUTetUIEnblUpueZertfy2yKjgz9/9VJVQg9VvT20E
wYqESys+THd2k3wPPStE+D0ZUpIDAIMIEpi5jG6+aA8NYp+Yw9I7myH1D/USTIpCHe6PSpOqtb9a
gxroMSuyCqAvYQXNrKe9L4U3R5kx1dsB63BlOsYQYX7ZPfYrrS1ha80mxXwAhmK7MrsEN6P9Lk3i
3izxXVMQirYVi81yNMJuFTgEVMkWwblaD3wOWAKoEYOaO7mxlslQAT8d6wgbjNymrNzjPci3YDMT
rVGNMFSQraTRHM1JvtI5NPI4MfLEAWoZidHEtINAyua5whpPOYOG+QVMse1zxoZrb53yDFBHKLS9
3DjpUtVUs+ZFohmZ4RtPNcSSJ+55Dabv6Pu68rawkQOD/EJu04t52OOTIPHTWGaT7EhR+2xl4xQP
cE90d+wyXIfx4mxkS3wUKLi0D9Ptqgu/Ael5PBiQrWtKIAc4ZW8vxwT2OnDesCEDrzRQqrSyrz++
nRj3gRcpWi0MlTNp5mjzYZTRw3bQ/h7a/AkrsQLcJi6FL91VfCg1jw5PcQhE6KFGJcAFfoIrd0nI
ypfEOBGQZ25sDhnbiAOv+/UDicjwuoyxhY4HKZ2UAWNER2kFTYlCjSGFs1btXdrLtUcuTNbzcc7N
gUAc16uTEZIOkKu7yKs1TCkkpY/ndchbC5qp+FO+KrrAUZxqm7Uh68aaHJlvaAkwD1gTydoAP9sf
rDCryLpSceWkV9kUzG2JpYFikHGhSgnM0uYFembpdpwN4ZbWTkX3P0zInsazEHpyEGCckn9Nhxmu
JOuokgjXy5SRqo+W0Meu2afi665nlIHTo7AxBbfubbfZk9FycsiLz5jPZpkW3ho3AT9mKYHYlaKK
m/HL6aAFPELZgPW8BlNuTsRdQ858gQWqCXfCp3kimlNQHuPABbEcQ7BbH0tYpqVIpj8g/LMNXR4G
jR34yt4Vl1bpGtv7uEihCnphIwa1i65xKKCZFAjrIEuyegS9WPSjWPbo/INBkIYtmJfN+AEZ7VjO
gDAvFqOnmxqUhH5qD72BuKnbzLove3eVUi+GHpJi4tEUqK2/V/LZodmrEOyABYSg1ImR/uvemlBN
syKH4joh/WY7rh+wjZn9Eoi1rpL/sUnVAVCBRHVyeqZtvZmthary3HIWw/FwoBMqimvhWMWQWnkA
pvOEuJJ6bo6oHqej6BIkjOLfVehXG6Eg8nnbb1X+FmYrWbq5WoL/jpYLSIpsAxM3mzfHY0OXgpxs
j/NxpYlslmQuMJSCnrBgCSS7KrDVR/A5W9yDF7FVlJjpHd94FGTiUug0Itb/23nTmizc8xZ9QEAL
kg2Pu9b+ngey0sO36rEsvjJfJm2VH3lFPq9S+DoKhGoIAm9Kxb6U8ftMvZWwGpp+hRdq/WbgN7Vq
aWMg/AZoVz+UiTTMzfFaNq7PSISo58lKB64VBvhNMJUwelnIfDs6xLr46nQD1PmJ036CUS/ldTuy
LOAzbliu1Gus9fVJurVwv1G/ngvlkDus7eH7UR72OeN+LnASewTBjNkeltjep2KAMo0jRfHsjkpF
+xRS/MKxUAlJZ+bUSbYktFbCR8TiRGZKXo8jd3OLNkbnHQ8sUBzeCOFcLlLH9cPQkkdGIjZIcGQs
PdpqKvwM0orY9rcdHu4bnd55iMbHEeHHvH7o8ud8dI+QSoXkZVdL9tBJev5BeDjZw796ZiUHSXPa
vpGqC9w/5H62TrH2aWM1+g2m3fQBAKfy5edr0xrcBaB7Gz44AH0MOuR1MBSnK9G3JvJBjPBc3kfL
ybcTK5ura3A4kvWifC0960RRocvZtVmBfO1dvFRnSruS+KaaY91q8z80mEDkagzZIB6mdEKVg3tH
S7PQhVDxg5ciXOTiZF8E70oeD1JOy+490jgtNEKmTly6xXVlvscblRfpEH74JkKMqBg5pWhD9RRP
2YqqjJKvY0iOB93MUsaxbZtlAsgC/tILXZUDz2tLAbL3/q3A42AGYAoDrAQpBrA6AqRbofShZEIM
huTpJFxgiUUgdA7FGdWTYdXVP9Km9HPZPqkF2yjDQD+Ni2rxQ8I8jwJiulzuN/fhHIaFY9Vf7Mys
Btfr3+KzRnrkcrJSGYfqm4/oVmLuaEPApDeWQ0Ah9GVWqbWq0PDGWATt8Wt+88frWnSv6KHAHV6a
PtJxnZWqLqPBQkU/GPmcA4P5v36oSZ8ObX0+pEZshsd5FBCC/UF4ygk42Y7bpax1faBXqgoZVsSZ
iUQ+n9+rm7sXF4r3lOaMQKYAR9vt9pTH7H0hEEBb4CL6Eqhfth4inX27wMH72bRjsA4EboJJVEu7
koXn8d5FBPZnNeKU35n8Uq6mE7i82HEXPli5YMXp5LVqdUWRsGp0oBcspzdRTvnnZlxed3dNUivy
aH5neB/klmiCqp0GXcK4wpn/oZrXc8hDHgCIBtQMgb3O8HDt2E2Yhk995EJ16giFexpCxlvREdaP
6DFnEUnirwVwFpEFv8AVlKxXWw67NZl2VhwoyBJfV6ze0axkozKEInpltpRdkfk78oopYPu9xitg
vVbXCQEndmXLs4AiOWt225RmfjVzKJlro03OuqKoGoLvIXOgFHfjDcHmHKiv0cGXdlnpqR6ea358
1sZQSoY4AArUxFZhVj9rA7asWvnUDYRrJNzBVHS0VRvyNTBF6/Bgf0OedFjHIA4GHAYXm7UvTbj3
NyOBGdpZfX0KN/BR+mmc4JabaVCGnw78LmSxPlbrbvV4+qbsdLmd1omd/lvG1sbe6h5jy0VU5SSq
loZMQer7xW6IWF+rRHCKoH05nKVlpgpvAryAH0H1zb1hBw6qRKqsnAHkUAyOdeMex+jqy6IrL6j8
XWXYACCs8rQl4yzaqkGYU64W59JpeLmoILcU4+aywciftkYgofcoDzCRwbBxWB+t1bHZSS1fG+9y
Bhm9VxS3tdqwTiJ29VQKSlYXSSagMbSCyp6Qr4ZAVypT9WuDkKIduMUvfdRVjGSHH/o+1gx59XYP
4ygU8NldIUo15pFHNPs/x7w4bGqn1s2wGCVoxZc+uerVhzd4bAm9xmabAH8wtadvvD5RUjBbdfHB
7JkyhrKe/WEcKUSWVZtpnOz2dKxK0fnQd54ZEYVgZcZNJmEx2sSeTRSCdoMLeoXjgP2YlvQ7JmLQ
ldrYRGxhASly9+c3unyL1j5v3Vre0gH+pKXS1QPn7krQvWHdwVlhTFOBohFvs1ZsimpI3no6hPuH
kAy04l3Sz25wvxGjxcfpI2HRJ38dcd0iWzY+T9FcD37/mHhJr60ivLsMeVENEmRVQ2EkMpGJHQIV
CtVSlKhKIvrHZZvwlAzVtf2NzJrBn7AJEePEHJ19MgHyd+rNs0d6l8q4lAUqzGImzGfrlblGQaPr
4djRmZMCkJCxoia//waukK4OOEOK9YueeMChvNE7bP71e7+gaP4VOgU+c7zmf6+l5FSNryMMZ4iZ
+Iq8c48JVPsVKmC9zUg6sq+o412a3KCoOX7JDX0sBIIja4vC8pLl65VAAOZfxRCuR+3NYnj0WoKB
SZjlvv/9k/iQrhw3BmMb9musA0gfEgm9g8FlnYYw3DPslDjtQYTp0EnHUMwWjlTG+De4uterWdVd
/8hWwe8l5f07F7D5GxWUwcUmzQzr85ADZnPCxESLXzGujm5LV++ofXdSydkxFIW7+Soj7So1rG4A
cU8WqSl+fBnLSYHqAbTc8RzT3SxprKzCZGK+3qfx9T1kPeDMd0EFwfw0uvWnCda6rDBtiR6pd4bz
802l37ApFo9DoTnMDz9l8K6aMRXVcqNr2X51wJ8PWCPqIm+0AgpPsmvCB+m0GFz0ne2SvGySnAA0
S4d/FfqQoBfrEnJfqkYrjsDvNxlGpsRJbBzqCu8sDbuDzr8D4j7Td8p1LzbnlRtaCdoygfWZfVSv
Q4qSkKHimjNxWGVZb/0tLSFfYlenwh8sCPz84fr/YkhonrpZznv+FlYVGG8eFmNMQgsYzOoYIy27
uNZHC73Yu+UIQF+LNcbLyx4TWXS/3qqaqzG3HzRJ2mCwF6weo758qI5M/xWSmxuxMmiAIg2eJexF
7hpC5vo3j7VerJCYIqlQ8yA+MXzl5Klk/VWT64/mzgNXMe9rXnRFWDkxXmV28hDJRwXbh0REg2/L
A9DMrWRhObIs60nuHqoMlbU0RuNrsZLKoUNR1sfgBgZVFYySuUdrp56Dd+u5qclD4AnkLNBQ9iNJ
H5NaEeb0BWH9S1PDaQ1LIcOM4CU4qSuiEwVtGHlkEh94KtIFydNj0SX1H3X+tCa/cvdlnfsAgqWA
4pNQ4g80TeNoSqAShw2wfzfHOcsaIkwT1cw9A7q7dAOoYuMQewHXzYhpEKKfBOxw8akVpUtgTE1v
+oGm3RQ00E/qEdSDJ7/vLGGO9iPHb2YHBBTnw0Y9LLjs1dgufcXIfK40gEkDESI3CJNLiLnkeG3x
4lAdXhCDwNGA+S54gXY8B3a5pmZKABy8qpCMiirFXXKtz8nJ6EVFUcpq3EZKFWRAYWEZ2xe1Slkp
eLbB5kai8kCkAzcDlniPVSUGvRyWWz50aqOmWmaAgn/KUUFo78Mg/HW0mQWzDA2OAd0lnmiKG+eG
0hMTR2Pov6BNlbTF/npMeXtxYjeOFeNyXmbjJcUEVQwfJc0RbvmgnlHFaHNnlwumb3FOdjbRJ1IA
wmRKJmmDJfaFwiWHpAiVLsgl6CiEIH+YxHNrWsnIaMNYcrEAQCbWPyJ/AthVcM+1zPEaiFEbnUlT
f12q6KgaL/Arkftq/VdqS0jkjU3jfpAcrzxHY8Uj0JRd2rKKAI5G4qjLi7XQO30/RAHEuYQ+zv59
7cplg58FcydlsRwQgfp4pipaIlOfRMrdxiWB1lgwfz2jwbc/RAsx4GGggnTTfLh6E3ZUF/J1mIQg
/Z9B5BuOLgB25GjN4vYJOecmfScFmmtV1Y6gdL35S1A9UTXYUMThangOL27eqlXsCTLy1ZXVtmJ8
wJGuzjEcnijBoVP4tCesrnJScMQDAIOwb1cs+45UagqIT9L/E2qNcRdEVe1VNtZC/M4rhTJwtI/U
dyfEqweB58od+HfUq2SAK9V+jy7bP+dFNV2Wss+0JRKFgnKdOM2Hy3SUbJB9ixs/IO5seZ7P/bop
SKixitGmX1QO/06iQvFtcl7f0OJ2XG8LgS1EcBaJznXQuH1ZUJFhAw8SquC42BURvf6l7Bbn1N7w
4KdcEXdHUWAVkgocDncA3l1NGJu5rYZ1zJaMFxVOnmFPXBkQ1inU/O6tVX1eJD0ZcFmxtLBs374e
2c3JjP8X2978nSj11JG4kh+iaWafTSL8N/heBGAwKPaZf2lIeByJPVWdcAwzNo/aVX8pX8NhVnP9
HCKdocylQIPGmSuBsgh6jYwRyVm2J7G6/MZpyhjJ54Aai00wEf20LyPXpgk5zuqX6ThzBwUrtCYm
DSpQucnZ9gESgWXsX/lpfwJJz9+H+29Q5x8Us4QWkR9XqooliSdfIF2JC5Ry3+3EAWoescKsD/2o
9kl0D1R32dZFzpyKAe+EUqFAOQ8Vp+4vhXUpRWLegfeX0L6U04qW9NeSeR/iyUXHaK6mDn2aXEDE
8AydTuk7MX/NV5W6QI9goqJc9TD+dAPgqD0abtEdc40hQoeA2HNQStx+B5fvNhCsQ5RI3Y2Ch5tU
3CMYpBOB6ZobEro2ge61T+GeYPC+5EtitK9944Tg4YlEwMibJQqaYNDgXYCZAda9NluXZLXS4mb9
rKQzKJeV36L6TyoBI4zpNbY56QNEJCTSC0NUe+a/li7aZQD5JJIjlF5snLlCGR9X69rN1ZMefDnM
kytWlHjOvkCyhAnhNCSj/bWQFHk/ZkMNwDFus5tYrMc6MV4iz4CwJ6QDMcsx5VzOZsHKOxyDlTg7
B6Bdn+jz9du4dv9KUCmwqg0AoypMS6NB0d960xMzytYEVfQflGV69KVi4DSyQPKd3FJ6XSuLBT/P
aaJj0ck3GBaG4qqeEdhKqkdhH+HAUHqGhjCXBZj8xjydquif57bDBu55s4jYtq+W4VS/LoKO2Cl7
VA+BnPmny7k7Do4T0WmyDIFAxwCq1Y0gidrMKJnvSr8eRpFSIJuzDwRaGNPl8jdBM7a+GXzvCI3d
A+Ll3LOt3TzSP155cgVtpADidPB11UOXIX6M0IvK9XCLwhn8EBRjyaW0oO4fIo3rrL0L5sWtDVRh
QxfXIfCjATfs9gqNmz7IXynN2cKxXFY6rI+xYEnjIu/JTs9KePglYeGMrSC+wxepYnrmVmVIMC37
OXQvCegEzBnB15JCqMsh3kHqx75RK+f5Yudlx7iSNp7WZ0sN7zaF/FgCIr5GtdXSw7c7owx85BM/
a0NnUqbp0vLxauRVS/CIY+KBQkK/tx8N8f2xsYFyBhuXXdHQok7+KwmLQ+ohFuEvgkqKHAmO5N1P
kOeI5d7kw42/QQABDao/eOEDD9xwZcNgreOEaBI3DPP0KBnH7uVnE7aY8DOMpv1dT1m4gZzTXZWz
JWPuENmlmUsVshVo4g0Dqt2RND3xWcjcyIGEBU8FRJxZHdSCcTC47DslEWSHyaoWK6h/9kbZL1+Q
Ev8/CSU145R1AGBuzMGRGz/Z8lc2IQwJ+24xIu5DdEo643qQKtEboH1f25bVr+CWJLo0YqBCQsn9
ln78MplCd9t98wEqyP5wXk2Gss9afpxVz++9Qe7QKZMrxjauGgXtyN79T/VQODZk+5HOk191ZW7c
wt+Z8fVbmT8gxgNM1dF4XTdbOpyZufeQgRGNMqKmg+iN6LDLX+rZn3ZLtoyVhtH17D6L2KEAXhrm
Yehx9FtHDTemYJTxM0zbsD3ieXveQkb5j9ue5MQxvHZcFLxUIG5sda+FRdhy6+XQM1LiNcpoNCKw
/W3wRoa0JHxhoF1ZogW79erlcLmuZKhR/2l+R1hYVntpLZbCWY7G84bZe2A4/Y+t+5+pbiO0uoVy
mZ8e7C0cZbMHlAiasLAJrMJCTsNQ7UoqPFGKqA4i1YvPw+4N081ktuZYJ5w45fyEKciwlAUy2Wif
xsRb5Y4dPHIhiZNpsKO7hzL5bIN8AmvpzCkXT5H9oiW0fIRub93KUXYlQHQGPmSuX3FxP9cWPvTW
Q91VMVlsYuC9ZC3DHCCXOLHuVEu7uK5oVR95C2koadTF4WJ8LvAzO7nTUVrMJHrPWndAINgSyYlP
/K5k3frd3SGevfQnnXWeKhnppLUJQCAxDEtsIma7vECH7U71qAHkTaRvahIMbpk0UBO3aM6Jg2J6
iMjxe3eiy2JosmdsXKlU0Ri8M2VqVYwYApBp7ILKLC063uaadjMmH63AT53K0hsueXx7dM1PRx4l
AIeKZ3qNtMTRgVOhju3TjSc3K8pHoKAy1nKa6xoCO2XHpm2dNCBDuIf3NbMv+gwb+ecSGwaDPa//
l8mcIBP6Kbrq04E/mqkCOi+pENQjndIAeUsN1LXSlv7DZYUG0yPOnlV0mpk1DkD42W/AuxJ7CSt4
LCJE3QH4c+gBTqlGdQBq6nZbSSxnlCZi7zs8JK19zA4bDmzII4KtdfUYFWc3tfZbArb2Yuhzz73W
O7X/k9RubWtXZcBSDJ52SfeSChUjksiuEbkVf28MgCjL3YI312ehIwEM9If9ELbCPNKw2womj63p
+LVDxazQksAlB6KN4bOSgJylMErUdcqwm3Jd6vRiNZLK9fdqaQuzoruW+baytoLMShXgHF7JAMn+
j7jvAFoLdA4jzfj9i3f5vRQIPxDU8QplwjXZmJ6NRH3lQNdlbP0s9/ywDc2x9qJZMcmNtiySIic2
b+W91IqW9Eo1RxgWnvBIcntrPb0UP9YvlQPblrofv/6G2/6AEaGLCTk1+u16m43COXrPKi7JPZqa
nxFwD58kcRrz5dyOudASO1MH9MiQcwNNM9746k94BKv/gwz329GtPvup53XkGd7lPLF/YDdmQzCX
DtU4z3uNeJ3fAjNuu0uYaAb51QCj7z0YUqnMjvcCVs/XJ2kiJbYxhXuZ08GUo/PJs8eNGQGz1m1B
8WLstRz+VaDsbRDBcSKkRTdQ3xXotTKuxwNrX6kdbADeX935tzVCy8KpgKDvvX79TIEa0I3feaBT
fvqbpI/CsaFVC2x2fMV3kziPfY26OOv/+vkIFhXxOtKYRhPM9PObqyyRXtRaQd/frng4s7BnUC2n
LtWyMXCu8KvjhC0r5EZSynpu2YwuvekzjXXEpEJV1exKhIA4A8fUB2XKhKZUw50ki9cD7uhWKjwG
fQf7QxPUVyxoRuddGVBXrKzawC5X7uFgEmqxt0hA4VhS1aI0lIcTF/yQmAcgLUjbRa+ydONFkfar
Z92JFZdheM1Cr0ELrBmL2YJyqzIS6BaInizHNqWbWkmv+XdAWuC65mkbDc0eOIt4nIq1TDgB6lxo
fD6h5232pXHXv6QAXWDNQKvsCz66yw28tWTD0lVahu9dkfK5EM3msTcvEDV85gVNnkQx3Lhv8ZgL
PmyclqCgUMmwhpMtYIrTYXMvcbmaU8y0DumAkJsWqbbKSu1pSVKrZxrpTnemkRqaZE52aNPb0FaE
wXa9qRXd02pzR0mm60TJlOyO2NAjNPnca0Kydu5aigP8HvDa1O0//B0cyVXHvyt8m7zTtnR1STp4
L00B8wm1kDKECMWmsEHls+EvXr79FsW9ZH/fvzSzrc95yRzssGsWMQ+iwmsuwKJYBW5wD2U6GHzk
yVrRGQIWbby0CCyTrJP2yhSLfrUNklY8pDD8j4Nd2A/0Z/JXhL6uqzCDra/iOcT5zCMSzWASilRZ
hFrlBsVOcU6QB0BUrxEZiLoeovDijD9NYWpc4XA6OZR3x2VUrbk752Vdf4mpVBYzUD0ahezcIAtu
0b0Au+fm7w5d0Uj39LBb2d9ao3xiAVC7RIemGu8m+CcyprooWbFaci8zjCf1secPmLFg5aYGLcne
IF8bS6w0mXBplH7VtDdkthYrWE7W3zjbCwomjtuhTQhowB2YOXhdnxWE7xHmZHGyXSoSV9hc4TCi
dx6uoRFoc1ze0dCj8vVbX561OXJAvD+cpyR2aJ3Q4CaE5p8b8bQJaf05HLrelgbZuuxPA1rOiwnC
dpQy07/EnLf+uwIm07T61XLqh91Y8wMFkgOAxl8+/lMVCdABXuUCyzQ0F7csQ/y5G8ZMW8ZxaX2Z
ap/q/987uRVMg6AFsjIKM4rKTjp2D51o4ys2eIgVKKsZcbtwydxy4sSbeK5HDPtlSlr/h4OHuQ5S
h9sG6WURppRw3fYsvU8lxJnsU6vxemsQaLkO4kSkAS7vAqUB34Bmoa+KEwp6ui07e916iJ2p6e9D
SwAgLG2SidzBAbGnWNq+prSm+pPwNgqcElx1nHXMtrUqE4CTH4Xx6zpAI9GMVlk5BnXKgHnmj/RK
shuHrUYEtd3HEy8MiimPyrVA763tXhI+LATht/o+Kwbdcn2yrGYwNyfD284Gt27K5pUNfqfP8Nri
qnfcYQogTQJl3rvv/SfQOG96VpDvzwu1y+/hvNNJZ+qvPoy4wG851d7KKaEfEaW/vsQbLT6g8L2e
NPnslWETOL7Rzkm9poqrk81jivitPwgCq8x/y4IshWgOImTZ9tHhF/dHb4YsHtjXNkK6LFenzhD2
pHSPphqsHO5yKK9MPbcGrHvYZEuDTxgKFRgSEH7aYlcWBDfACbdSdPSp/dIpMKY7ffJTQXK79qjP
MlkachOj/8hTnS3rO8sADT5IlDnzgVS3eexFo/MgJSM2MsM/VWpKzOcopfjvc85aSKBzhOi3zfh0
veUu/G+oTZTY4lIGSlIcrgWwJjGsHXhCcbQ3tbBcUzNmyLgIIQiCXeHBNFo/t29fHJKgP3a+nqTn
b7a7Z/luf2Fr2e21Fwy0x27+NLfG7X4iAzhRKsSIXYXwRk5xZ3IDP5TTMgPAsefFiBBT1tmmSEYA
/DIcK6KWHsSvEboeGMVcIrX4SBW++zSFtI4zMIFvKX3FJvz/o2cr5c2drbYZVswYP8o4qWiR0Ag8
bJyioXfWe0hm2s7yVE9NkQ580poDlLQjGFzUxrW9tgiHmSejvEEwJA6BDYkQ6esmltCv9Yt5PiRZ
Lm+NnDYMGBfvflf7W2EhYhGep3yYrmbhslZjb2tWuhyzAopnNg86HzX/tmUg30S3sxjtFtiVDM35
qJPMD+6PdnTyTAbc4+Z1HTiFeT7dN0U6e2glhz0C+T5P1lHAFZG8s7Jz8GjRSs0D6NzmccBmNjgt
nTMJEdRWRG4pcM0c6CH9raur/O3wo3W7faLejug0ah+wrL5eU94wOjKDhT9S1/6YPbWZ1yGgw92C
kI43y8YMjsvEWV15DP0vRJBC6fzRd49EsqayO86KjNEBCDCxOQHkfPhlnqePhMRrSt2oeQ3O3UIy
Ykf76BgHsHjzpEjtnqfX/NL2z4x8L2Be2PUUyW/fiHENh7w5nkLHgjOAFvnpn7u0CXbDWer7rdst
BbAEwND7vKbNg4PP57sDHC+uD+ju34DvaUNTJktNnmeACvqYmGjKyvc3ayqE1SqxKowKjHeGCSiX
Fd4vAtHNG7ERfoMriDlLx6VzLdUdj86s8+wnisco+/1lXaZh25Ivtdd+VhQaWM7rBYX8iihDBBle
N41AONLT6GZzZecGhD6IB0VZipTT0xwj/5kWK06YAAPCIIxhWJftrEpfpgZ3wVZs8zcKzk6SYKxm
/A2u1rhvTLnFRxBHQY4REMPJyFIx919EKRaJ5S6RA3+UklYR9fy7zENjqhywZjTITOtdYS0HzX9H
7+pEeWW9DJSFNRY8zSYoMz3D8MsrBUhLz06eVvYzrAg2sOabZNEG4zX9Uz1jpEtAzxFaJ9yf+xg/
8YBlnH9DoRRCDLTMxbbslK82hXoslztmgcOn7LIbTNqvafcg1UOSUP6D3YL1zGbBVllK+/ypFrp3
QEz+ZOTN4r1fPECgKckWehcaDqtHFtAgtdPR7Ft6TqnbiaVFiCXIsPLN3ibWo40DPfRSkjz9/zPx
V9po6I/Yj46y16QWFKXWNsRXWXz+WAIZWjCtaEwIZMuR/rIMz/K76Dj4Vfpq7dWvJVFbf6U10kvN
7XnknvVAZ05N9rcJy4UonQ7KD2UIfMj2/+8ccRePR+v9GzrK6pAglyf2+95G1G+bOGJWxcPdeUE6
USTQxoSwfseGOWl/Zjkqj1GeBCWCFF3YF3+iNqqX0JWp5N6T8k/w+cyHhcTqlF8dDQP7B/wFzkux
XH7+fHwz1pJw1dl3RhsQa6seaC9hOqHxIDiHuTP/n1enap2QWQQMITPEyR5Xr1deTw8XCoeXwJAs
MJPT8VwDGKbB5dtARrQPICldCZoKUi6wn5pfZGJUwi85qhQntGTNdceTkMIuPv9RZHLs0BMGyuuC
sy2leF1+rCwPVJl8Pwdw31QtIgOREfME9qbd/SUKse5jdzW8J8evww90EI3Jkva5NGfNd4sw6wgQ
m7YS3ASt12Zw1WaGxX0OcWnA4iEfhO8xF2k95oWAYvlPA4sPjvBif77QePyNScFrAbs1/VY2sQvY
VqBlFCMHXFMNQ5aEWbIwP8ezU8SXwWsolSlWjNB9obV/vuX9Px8CAH3cfRRQ2S3ifxMTfq9Hj2K3
Llze2tEW6ffG+/5kAwTMden2NaTCuTe+Pzk0gDMkPMZW5wMLd6aCsRF6AmlqFE04o9os64I2oP66
B+9JPua4FThtKtY/F6uyFeqd69cFgTpCkwl1bNkJA1goRHN38ADueW4gqZuIKhXb2X0JrNA2Vy9F
AkOPmn+ACNZb4vVhz0rQVuZVwB9tK+ZPaedx+io5fX1z+R/z92Im0GZC10GH0LSA4cwjhQNTy0YE
jJ6P2/bMkYrpX/X/8qDgVwlyAjyBvQthkL3rcWcQx1InXTRLWDzeHZaigyz1NOzHjnBpis/DeBDi
a3DXmyb3WL69TFKD1q+GGSVYj1B067lyp1l9kIV3XX7zv4WSlavu5ZS5zrHed+kJ1XtaewNXl4E6
Dxdoy9PstV2zWrmdFNjqkzHrkAIV5oJn0wXFxnTkdNEe/03pifhgaPbov4Ir6QsThY0gR2jjqeFa
SNGoXTd3Mf7BHD337TWe50K3qCCDIiaZ3/JDc8S4M6vuBfxzbTVfPQ7Z0uZsuLRwEjxXnE11NgkP
aQsKq6N6gWDugNEhksLuzI1OEcl4l4NfPJ3IpsD1EwsqQd/cmDDIKi+C3G4c9l2LCIbvmFW5jZc3
OntWei14OkGI1R0pW/Xo1lOw9eyrllW5CYE8t25dtqFf5iHOWaGVizx+mvrniXdEUulwQ4a6mId1
M7fwX1UamJ7hmCKazYtgFq28JtXquRXoFwiaYDEZ4gK3wmWvj2vzdnkderfxGobIxADoc1pNWHRc
8evKeo1nAG6wNyBw/dH/53y5GaOWoYGQXzruGqeLDZg9+lYTRTfc4VB1SGJKRrfjwx8Q3k4R7uA3
m+5ZhRIsY1IoYlSVqp3LOSD5OW6WEAnOnn5s05YAadEN1U84mSL1LJdAZNjdVFz9aw6FQyyiI01X
YQGb65CyJj6uY2pBbuiH2HKBcC0gkQmXBOk66qYrzQRq/khKBA2nx28xWQeEeVUhgEyNRy4YOP56
NtLt9xOcJPsTZaXyVlvJWFQqsafUvq2tokyIE4ikNf1IvRG5LjGYgRiI9TaoKAWC1UyWVQjrTCdl
DNL2/rjMD3kJogYYdVHarLwDmbjcidtJ1O2QmKRt8YHphKL+LTJwth+YVbO37DOpzxdEDa7FVm4F
zUt4/5v0o1n2FmdJQ1GwIl8gUONiDTW5czhJRTPv1uAxo1bCVbRveENOl0LWbgr9pZs7Vu30JtJA
+nBKQ9ZoNh1QJzb9LdBlE4p8limY/JYvunLq/g93YPgauCTvXxHCGuMM6vDVoInQhpMIpoQL6g2a
znGjwMuTDm1him3YfAhlPjvkPwZZcghTHC27XIsYW0EGrBy6I6lelT2yjKEb/r8uiOm91bLbW/QX
ShRzWFlTJABDU3TXe2jQADeNcHU7re9laWEb4ulC/6c9BqUZd4aUY/IV6HZt5TqIGl0BMSLIE2MO
4wZActYGlK1b/qqJNiB3sUajozZfpchz6yT37/+IFu+hqE+Xmi3XiMgIfhre1QRSmDJndDWQ9ZE0
qN9o4mScbBFayLSfUrD0VByQg7Rc5qTuOGLrkgg8tLc+ZwpKQOZbKh4YdCavP1GPlcDQGMh6EE1U
Hyat9dv2w402M0vwKNXnnYbFyiC79hhkh4JKztZJ+1AzWy6KDFjFHZ+E8sR/VpZruVaoFvJ8NDEn
3yItpepVN+D9jKqEok+sR3oB1vhNcAfj1SXxs++ekrICfwdu84W4Zh7h7zEBFo1U8p4BovulDzAP
zBkgb1i7npkHqLiogxnMGbc6G6zokHuB2lAJncDyvbz5n2OVL3jdYEcN1dUJ5lT0kfHIp/5XvrCW
aoInJKQ/9P6ixeWONATNToWWrQ//UbqRzWo7YTcCQh1Br3m1+u5i8AWBaEYFaCJDpQbaHyV0Z04O
kNsLROCCBTHqT0hBj1z8oNcBusr3ClZZ96JMyUibfn5TP9T1nino68xp0CigFFwak/gNKlDg0Wpz
IkcnF4g5t5Y6QyRKle+ydnlfpWIYwgeQE3qfyHm9pM3Ib7O5wE+GNJUiL/R/322ghJWNarnF7zOq
TK7ejmBmOvddO6xy+NsCl+ja27BHDtl6FTJ+BWkMjlUv3TjX++XZ2fmwaI1fw77TJNN+ks5pPVmS
/y6tGBRMX7ZbeTyFGz9KDHUS7IZQvprlOBRjplud6vFjogETobAyGRQyY7/z06DpiUOryuEtvYXX
pqb6SjfG8GD4TMYLzo83yHAQ5PCJdDgjJ/PQHi8T5dPXEJGW21cU72j01uv1fndJ5LZzgsRpWVkJ
T7wg72wl7bACbJq98e07j7zfVXxzyc6g21mqzB3wJFQPBZlFqwKL5BAWTKJs6oPi7Efh45uKywIJ
mShZFKwMKH22PuXRuIjqXOaPKdhBeWP3m+4E9kJK9FUsAzeoKCsSGugyDag9YdR5hYxOXHitox7I
bRF/yzZG+Cvo5m4mZ6CDBq7WfnpbPvmQgshacdxKUQ5UEOFbgOg1evjRo1bVXduhMk/2v9ksslkO
ujovWulgM2JHOB9Wa3RL8AK4iVoPMXwp02bCps/0MyRjiDjIP37aTOdUDZDIt4TKq0N/TILIlt+J
nmO8bFHSU9mHASzhW8wce7M4uKXN+GUNJhXGeTh1DHBTTPjjQvcmFPPml26/827SBv/n9AflNyxC
fwMbnsKAz2wE2uN4jNBWJ1BKYi8cgk5ITe08/EWDiAh3IkBZy73DxcMTERJ68Foq6zkPkhwyZZLv
yYAix2oI1TuyZDHr04S8Kn+kjd2YRO32ZvXH6s3/glNwSagGTJL7VrmHAv9GHXQUDZT0kaiXRPKe
D4Dz4nhrziSPkANINAFukDhMITVXcsy5RCcWcCb/3Vqb8sHngunhfqWHKbbGLajlSl9qMBlc14sC
7IQbdfa/o3YiNaN2H/6wluTcp2jfb4RPWq/BhTmK8JvyjLOpITAPnNaYihk26CSF2hVGnSNNwYDX
mWW84glvnvY4ZZsV5CxyOWG3Zo1u5bQ3zPBrBFEk4Vq+z7HM1y4IvZ+A0ofJcfRJHSZ+xsjQ2oqf
ZMfVzJdHve0UgmLN+yuaN54bN0V9wBCnXtFd8H8YmU0joZp2LuH1rpFO/XqxkPwPnThbR25KwIu1
+ocZcoZQga2sC+GHrbx/Y2DDHwljW9jqwxJaFSvleAzmOCspZhebCTa95MCXKVV87jdH4dALM4WR
njqWZ60xhlLYINom1PEXyR17usjnr8lKWFN+pufASzcbM52J3cfaaAf1Y5oE/Nlpp4SQ6s0rpEif
rdtMvAP0SFL/4rb3h4Fvnv3T5P0OET+dMzgMOQQsbztQywseYcQXuc7FhRSJT2FVmKTjlGuW7+NV
qU2q1y5tNfEyWysZ0EsPGXBmXL3B+haawgmgcn8Vu1FcCyflZiTGcjG0CWX24ONH+2Mt40hQS4+J
m7lf8JVz9iFqR8AHMfAS/pwByzK76U+QqAFoWSGGqYJijifR/3PYHMLMjmp399F3dzm3hpDiRamv
WeBxNwEbUcXoRmTKTlPnbIABpKy2Ij2mpHHQDJFWATXkz+46KRda4HbBzZD8LRZkbVrndBMzamzy
G9zHBzyI6gYrAfwp8K+trfORPtC5025MFbGItdYFSSwUdzj0gbr7zeiVjmgqvHpMqoH+MG6A3mBb
tgWHZCMpU6CgfoAqkAdSDkXFYNuhNbeDNGBCo3vYOMIFHDOKrv6gdiPgTeOIASEnqjkH1Eru7qYl
S6kLxdTrCELZ8kSnWmgaCF08tvhgBwQl7aF8+xn/AW26tzuzzcAFaehZ2Hqz3Ho18HIjsVrnZ7Jx
u9WkKE/nEUuTwktqxsgWsxtQ56NQ7ir2Hds+mTg0eTzaPUkIPD9DRxhId8QNSSgwgJIAIXqZokWJ
iaJzyvVEn+37EX6040PSEzTRXD7xb1tTu2hob5eop/xT/j7Q8HNqJCnwRLh+4m/bawZwnnsQIOl2
m6ntec1Onx6vTJfHGsKWb0wyiAYTgCp7jKrQ0aiulJZxVT+cOCFy8PLBeqU98LhBUmiakNh1ZCS3
noTTn1/XGk5AL2pY9pu0tBZDd7un9nNlpAlOTnT1CYNb3VeNQcTsfs8xC6vZa8eizC25t+p+jMSZ
JH4ZCoGWX7v51JNnFKgOZ2L7oADP4ODIIq7Kk9Fp6qjnnaTel8qqfonyqscaR2lzQ+6VgWhzSYrX
tWr/uXA4209AEfeDjyGwNdVepihCUk6k5Vyd1xDHjzcuY4P1i1SyzAEqIwsYsyeqnC79pNZTbcc8
JT9aa54t/XFW1i+ArowrmH/6z4IKoRCyoWk7INF+U6+Yq7Z0ZCozfqnN2pYYdPWwDebm9BQtsfUZ
vbNUL4FERAMcSnOtumngCDdjdLrAKQghKXuT5WgI1BruzHpq6jU08iHjwO/z2cQm8RJROSfbM4RH
2+ZM+hxJiwvr5wA5jt3gRe1VUn9wSfRoomgFRf+tqg8XSUcEB7/g68BMEesM/QqMSoLMzicCXTpt
AypVRpVxYx18DOyuAVEaqf7B1xxzs2cX45NEIWrHTyYwyuhlGIUD2LV/2EgJZjwVOmz5n12BZKCD
8+2ed3lm8pLxnu/f2oYqisNANxS4oenDjxaxS9fcIGvyf/FvtHt5P+BeyWmcMBl+lBRUyY5jteFa
44poSACCxUhfIm8APl+Hya6ftcwemF/JeN+QUTRD37KNaPA24NJwBNRE7NJdyFtCUOhwvwmW1bNY
xm+uaX7acvo/B43wKhy1ZYC/KgAOivY7HqRO1q3o6Lzor9yBPs0rPXQjBepy/nlMs0yfqdBt2ZkL
KlDE9YsfrNBQgwk/5j1Yf60jIRb4kL8J7McynYDtlIZ3zIcsZcfgHVLWVq/GHr5i1QLlBjNY5vdw
NswkoJaM17X41Wvt7tF5vKtFKPrLrufeH4IUgw+vTc0uqParr4j42PibpkWRNkKIQrJVt50CcVFy
/hosXiWZmTgNFIPCtB6mA0G54m+v+OgQU876hivsTPgbFVQNfU1velm+emkpG0A4iHNTN/nmzGuy
pYiXoiLcmmIqjIPTBu/21spRT8M8/dPzHj3r1GxIdEO5XJSqIWaVQxJvdtKhQmPw17IT5DcViS4P
pp0XjFj5zMYkc7QUGDi1KszO+CWrFXSZ1xWLR4nQlVxbJoxKcUqX1wvjsLL6WPSU08AcgtNZZVEh
Xr/XrJPCmKmJqlpZH9X43yVCq1spX4Um/QSuSpiiufVsc2iVrGuNYeiUd4kTqJLOHKkmA4MvtTzn
e6NYywz6zb6NgvYVYhuhS3WMlvpOm5hLQzq+wyaO9HHinjvciBASxpNM9n9qN0jxzRFfoPdMuxGN
ou4Wp1WopJqFEdue9fq6WZ5CwbQ2U3FxCfgIop2oCTojUBT5cQeZhw3ZuigWidqV8cNOk/NwdAeK
BDmr1GUMIz4/a/4feFHszzRprx1Q6p1Z/FJVjhxz9wGAy8VObKTRUna8uai+7hMbSblpRAzmzT/K
zV4O1mVpKYw6hQ8L44j2EY+y3Sowti/XeIXcJkkWJOluE90a2G9yKKOqLdv64BB0clAz8sWcy2nK
v20w9k3xTH4THO66SVAM8pLZrD3i/K82C1MZeAkLmAUlhnHye9d3wcOfy47Zp1AVcTgtiylqmfRM
0bENApyNrtQ4J5U/QJQO3pMjhrWM4uTup5olsVH2DcmZSMm9aZRwSrybZXpF+Y6YfkWBZCTRG8X9
DghZ8qM06tEN7+Q/+NFj72Y9kAmqHwS4VhwZ6Ve/8dC012/QZK2OIDEesX4mOimOmeb60Kcwz8pV
2sAkQhIn37zmHARoRX7Wljk9XXGe/HgCiV5XuME7+PshU7IlYtMM9Ye6EpDpBfDf2JD7nWt31Jb4
ya1Md3DP3c51VZL/FWW5/Sp2rM2hGhYwkjWoRVlUg1fmDg1OEFz7jpvisvRFzmHayzkvMmuwvrpE
JOOrxuhpO32RYDH+li8JLFHMmp7DLVsbDf0cmf/XM1lxa7PdUgXkfUTI/qfXBJpTFJVCbS5qpeoT
CcBsxLE9FxFRP4p4NvK3TjJGgqnL18fGNgWG7DFRExqqZpOGuG2kcHP3KzcKmN0EyUBhE88czpwL
7a74F/EjogTKX3nECDXmoWXVSde3VJ2C0gZcFGby/Ea+fL7MgOcFUoQu9fzbFP/s1bqSXAl2Wi/u
lwbY0MwOD8BFebXJZ0pW5tLVh9D5DOb930wYnB3J5Cyustx3ENbY85DCY9K0V5k833U0nPGW6vK9
W4gSGodwwAC3Ea6pRiixH84oSwG1aYJJS+vcBEAmFRVgKRMl0KIn8DsRl99R1Ijv0bQyZhaZqJD4
ce6k8gVmbnaWK1cn4s6HdTbiLvxzHyBZCpCbDtdbe2qnpBiq0TF1yjCEV6Xp+n2OmyHsieZ0YqE7
OTJXk9PRHQtAWdaisKrBH/rXFlnbNanIHmxnPN1D8tdBW+Qjt0vZQXdUEJUr4KKXb9WzWnKNMUQU
zt8WeP/cA08a/7toN7x06lyY2siMcPyUMm675B4ZJQvP4ukW0Sug0sBYKTxVol1HTLm1mJ799J6l
CV7Jbo3F4f1Sey/Pi+E4cJ52/u1/iqiNSjirDCgTgcNeM5vmP49KCPui1WdSb9DNA8T53ndoT5lp
j2xJwewSyZQmMN0K/Brhj0zF7rgdUopxzf+YGRSTHZ+CN/wWrVJTk78t9pr/I/9nlpgwfQrQ/7rV
Fnk7y31166A+noTN9ogP3KtLksH7pdez/+VDQteS+9S3FvQuK79IYQGTJrKayFSn8Z/d2RH4py/2
YpL9e6Ya2L7ZYkkVlgC4t3NIb71ELMDtLHbsClI442UW8SdPV8yLZYqETrmAiRc70Nq/iyL513lc
jIkwvKfOMo9EuAtDc+K0OJiPpu0l8wS1b9Vr4nyq3+HDqcc8QRHv2uoFiTxsntBHSLp8CcRNWg+K
dKtAMbjC3KjO/EFbCKxqdFuXWoWP/xmE77UzUc68DAnvlzU54smRBsHR6+a14p6+3ZkomLSQ0xAT
ZFhibw93OznMTEcVUGjmMIRxQRovUjH3rWJrTIlxzuTUB1CsgCg0YXHhsHKbk4epJYEag+wMCCL1
Nlt358akVdLyBi4K7LceErRxF9mshqc8vhpzn0t3u+4eghbyNTEGY3EodDt8vbvwUkkKzRDA37OV
9MXZA2fVMlc04YwZFupaZ9O5PJd9lxvLXpyxzKMhB7t+YxXoc9gBJQ0VHsoX8fiDdKRAgJSmesTB
Ur1It5JGA0Eb+nF+nafBpGFpZPnjLQTxAtcADfnqy7orvzlMJEBbqMTSnv7uXtQbhkpkETQyL7Mk
hSVK5BJnxxIXMdere7UHIHG3bLInH4M8JKB7lpL0pb04IKDxmvUi3hYWHyUusY2q2CPOm0afeRBF
BhZjBl15dnTNzPPstrFIbsjgqQ6iuZA5Zp5/QNW9Wop+gF6OWAAl4VAwhfQrK4brQTM/vVz4lzSB
BDiJM4VaPMEQxDf47JshbZnXYFkIB5g7ggfsy5xLnpIaWyGvMij+M25MqCkmIxrM4tN3eJm20uOn
B6WacN+AKwhTEtt1PeIAMKnPBR93Rhk0SyXN02RBexNpx22XceWoSYohB2AWY7WpIj+EkjD+CEHq
3jz3ZgEPOK2fpMPZNSLSShw4Rg4f7W95Kjq818PTGfO8+7/GNcY9rxKUWC910/QdTTv5gAu/pK/v
peNTqYarU26Bbk98SL5M4um1woMt6GHhgUqo0bp9S6cepgnY0+DXEmIHtOqsEqCvAEGCdrkHiny5
P8VKLwL5QRDcZuO3u0mIHaDs1ae8NyYhE3ifn7r0QmTdvCrgpr+mC4+ybxDj49EqXb948J4LSBV9
vzeIxFGB2dckxfS8Q9ETanMixTJypu9sfRI28IpmKola54aU4q6JdF6TKtK5kuKOzBZG+9zOZfM2
zYWrr886bA8lKs3ApC6Kq+/2BCD1thXyoBzJtQGO79/HqtdGlalq4+AWSZppG4I+4Pt+EHnH1IAT
pS/v5Kbu4AWbzNwKvGhEgURMnW30IuCDdS+cPZ9yZsfSY+7uurjIFJs/EDBPtNgDgaK/UjlY1n44
/9RtJ9mHPZeAZRlGwq3YMRK3ZieMyJ1I1AzSr86+hWzh6pkpEPFSNw9XY6A18AEqldmsCBH/kALJ
RhgYq+sdOSLsA29/flIpWwH85k9OdLiFEBuaoyEMIBrETpGdvnJ89rieSxgDXJw8k9UiWKk34mKy
qoYZx3qhRoEDZsTNpg7CEIxN+H/LDtVAQQ3gLiGGtuLgEGDjkDUj5uMuBc3S0dRV+La1ZjMwI7HV
8jhp2cudfxzXY/Rs0oJNLoBcKYkycrT2NvzGbWa9W8eGKO2DJLPmefmBJRw81G9aN8P/jT+dX24P
/XGmsSTZ96bT1ywcS3kpEMtoe7ulyjQKH7zFaqU+IbzKJoajoMOBbrKc1rQGNBnp2tb+bdPd6cFM
4iRLpsAVmTrd1phX1tahyZjUgHaL3sDMMDKKT9DQpFuAzSxQQmcULBjzbhPBponeZmudWl7X6Oj3
H5ki7QvoZKiJb0BgdXACRzoySSeXWc3BFs6yaSy0p8YMRVmx7QNNpmrJuNaPK/+Jmx1Fxo94QRzi
Oe8N7GXd6zYN5K/QLiZ8uh/bCECnVQowQj2xLSzPysveMPMfDweowzHjRo+KaMmhqLxsBi4LlrqK
K6rFC4akctURh1x4GSOqTD4A3HwkGN1yIX5pn8WbgFyPDtmQU191pB15lJIoeDwvKRFoYE0zYMUb
aQO58Gx5wxZHskePI078kfxI4D1DI+RRbH2GY3ZqimYlpPryWKI/SVferg8Y1GIf5TSVmUsAgsrh
SHozVDifDCzjr71O9XF8S3AJ/q5pKH1dwQGKW/HkNTB1WahxTrIq/GgDSZDM6mFw81UjOW8pSlrq
hWARSeEZtp+Eoxo9425Kr0tm7Jv08QCI9jzhfVR2augts2jwdI4mMN7jXu8K/6Wwa+nXhmzwaXWV
6ZSss2Pg4iARcd/NTp88eLf4S3/Oz3KazuNFfTbGJQtu0aZ9P4td9ad0RXIco/xuzGV2vPuofaJf
3V8wjYoMc3GvrEXajX71SVc7luGlkmm5v/oE6CwJ2OlcHMLTNDeDRU9TSTDRm7fUcN7twp3DgoXi
/gOCPuYfG6KwlXQxwV76G+bZgQ5EOFFB/YOs0Hpj+jKAdGf49+Oj3n0zyVEzV8OIRdHsRNn1uO0a
ElNZScnDTCdslUzszkaKtLBnmDmVzjraoViTyyyhE9D1yRHL5zqMV/bL3MitI1uoqBcWo3iwYdKu
5lQJdK48EfZhjsGTwIMF7iVLq/rprEz151VNfGTJ2AveECPToZklh5P4dSitQjkWbIVz72w7K+fQ
Z1FJYLpJUbzqQbU6GorBgF4/OVdE0si3HAPaDcoqB2R8Bpf5J0KG/DAYv1KpNk9zDJn27rv/JyQD
3Oc3xK6+6XWK+BPTbOjmYvFZFmaONAZz6+v3O11fasPJNKKAkO2c2YUAevijLAnIhH1Gv1CCa9Xl
WkDN/9+yn6qMfDx75fVyytMMnVwPcgpe4u2Mw/vkD7QeMqrdcSLz+KysHXODEXiwUuthhu+vcKr/
+PWEfWwdagREHeXGLHi6mv04jwpDZYlrFmkqVmio84BuZYV0wbfdsDiiQK2wRI5ZZjh6eRdUF3eb
ODQOAisQ3MztNdw05ncrXzhPyqwGkmXOrcOrHRZ3BmSJ2o6xDCS5tnb5Nv5ZtyHuobpRvd1cO2lE
mJrgH1eTCFuMu+6je2DZ5WsGnqcV09aHD2kHrkQh6Ml8gqGXtjFjFxktbx8gYmGX2IFsFlmk9jkw
zdK9Uq4mR1z0NQEPVnwlJUJzbgD8nB5OVXoVEDKbC7mWrvDzLQcq2plYavU1bO83HczK/erZmSNg
iJnqHGLGGV5fBh6aK3Mo8qxIEGzymbBnQkOlw8e0hyhogXpvw1sc+MvVjIXrB34XHR5epyV0+kNr
XnLRAIFiXmvSMLMVUVmFjgPPDJTlPqsXmjl2tjKOO7HLL8zH1YM8jAACjxptVYgOXNvZSw+oK+/G
S+WkzchNVeGDPldmePgdZtBAEYoYYNS547PHrBeFS6WWdbWEap04BLED7NJtogLPghlRFeReafmZ
hkuuo5D44zZi9696fJJUmLTHvGEjVKEzhydSojAEPcdjdDx2BP8cBi9UKJAZE/sP0POGKjqmzROm
RbjF+oHCt/Z4rGQ2kBsBX2HrYPbRFFZkqlhKQsQxgwcgBhj9HUsI2Y2s6yr0QBV5twDNqqjg690I
hekny2XzlX9P4IkgZTfWoL7qTDW+N6TeDNiIFqHk9YYHWXVO1sS7cfXFp4vhZKyaBQ80MTr6w91A
QXEvfbZ1qxwljiulOip9ETukFuhUCGdMPZQuXCRLqv4ZsQiJRPLyAXGzUkMy6+am31HwNo/c+rou
7e5/LbgkyIX9pd79Q/gAsqsRUbJT8H54Xk6Bi1NYsAtN+S+DdZ4Cma5KKOq2+UAiojwdFgcdHEzl
APijhi1brF7949mBlCfRHgYLrNunRafndz8PsCzTXLtwkG5Bw7f3e3fkNwkkd5TvYRa560U57XCT
4qfWun00mITKLWpkT8z5IBZiVrsaKdgcFl2M4AhV1byJnFi57zgZnGfb0zli4PlBmo50SKMATizv
GxPBqslchwbcs/lNVKd7m4nFClq0hLoc12be2K3o8dinTyL5rckayEYC/jEDsPdgQhhAEWOpBFs4
X5KMa5VDt+NK5m/6ztxhY3JwCO0FesQV1ZoKnh72K+JoP3HPsB3C6Bxg7lMLWWF/J33fyV4MWSkW
GGcSJygq4/ogJzC0zpzJZBZ/mtguCc+w8L8nDlH4YU5vlKzl15xLYTV8a+RhLAgsQFfnR0qG1ikS
scFQ8OKgW+jlxW2lGRdZ2iF5UFnpPPQSVeFw5k1FJHdOHL5xzaSWG6ol5qOASK+d95xKQ8AE1r68
EJz/YO9SWTS8N/Bah1nP/mcUTwsvHFIh1/6khVnCIxvQ0M/mLWuJ0KjA/Fyz/N8T7y2f9zE0eFAe
r7tsyTPdW6QjOdEhUYCEHmO3cgcZSK/SqiNdLFg0L6wNe77/E/M68Zk+FUH1+EdkpjhghcUtpzt2
6lPZ1H/4qqDVFx6VHvVo9qmcolGMhx6Mty54s/mZUrGAnfHQNCRdbQCktQKqTiUjC8E41C5nS5CS
XDV5QujnFB5jTi467GogpaicSyaxEX3hU7tIrSZ6eMb2OZ0Gu6wXdjQyLgUW5rd8/h2TPha+14TM
kx2BGVlN/73LBpayr+9s6Y1u3koZ5Jsi/aBIbUnZGmUWMIhniKZFKZEFDeKOThtpZKtfgqVw+mEq
Jygu+ZWV5HshBxizz7GmFXrnGkxJnD5PIjUJLRfJw9Gs4r0K5lfSdzli/LMT9xW3zXC3BwTJwtZf
qh6cRWV58kvN3WQfRcZMeWiC7BhiTlW2QIYPvB9/anwcLVqP5TVEkWW6acglDDhiJaVxZb1/sko/
V5rvY7dCSNmtKnfqHS1tyqhL7LSBlfIAqv1zZcgA1u6vyM6LWYXOkz1TLTgx5whZKospmAZ6q/8O
uCGVTa6n+hE2jDLT8edebayJrNNIPEpzIquWyFq7MTt8rVxZRMEZ6mZWwK0UjA2JBqtccia1Ie/C
RpyItc1UKwUx0RfAO76CtzzNorexJi+uXyd6SaE0gdh/rDvk3wY+IH/69Up2uQqhCOw1HW+4pS9b
BC3fi0+f0RjyFBJ/1ZBbuPTOB2L3aVZfNM2PcWfKYP5oLk0OPaie3S1//k6V5jtkpX65DYB1neaQ
Irs8YwcCsUPXCor2MiWcCabDpXw3gGsmFkwsA9C48bTNlz3kQ5Vo/uzSHs2LktspabqR1dYLyz++
iX+SA7lqpdOFhFawQ6pZmwXsdJMweLSa5mZHVHvyAulweQEKBHkzZLLaGVfmMIE7Lmf0Ofy1YDum
7lC9R7H6rilhCbDr+/lgjwO88lliu8PEzY6yVRYeUxy8HOqnlmp8mz2GikdcJ0/cE8I9MEPa9wDQ
0/CvSU4b1rIObijbCWpRi3vcSZssaPAy4y4G9vAKoiK07dH4JFqDh5PtIIoRQNpOMRwjLqG4TJuc
bB+JSQdisOaowXo1T+qV5y7iwL/uvXvPykDbzxxHRt+UjuMsroNWo1bW5Sd+J5g8xWrM6sd5aBOK
bu0/iDRRLd4aWd6UY+0Onvuu0oMaBzaNxf+iSJi+3XnHfTnPR+wz8zaiJApQfQCoYch2msGFfH/K
sxmiUGbGE7ujWfrbBPa9UD7anbXOIKZe4b1mpkfCPJ7dn9WK2PVfNVMIU1yqDIrri/d7ojSpYtXC
5l6B+DplVcbUJ9/kmddQSqBd4zRvcCUEt8aFxxSOD0KKlfjVou0lrmNWKQrAONO4OW95Pa+uuavK
1PLtsjOo1YrphN+MuucQy8A6TQSWUshR9LUt8bVFXFiHARyhqiOMylWIxK1dHO1XFN67oWDz3Wbf
GGJOwijoS6r1kT9vLHwocxeCtDyZMCGZP1lz63MUjT9JQ0IeWQQaCa69sOthDqVIb3Q0Q7gFWtR+
/n7rfzLYrtMfqX6ClRgx6qev3AjGiPUz6IfIBRCmRDBvTz4fD9EoaWpmGuw7OfWIxZGs8mTu0ye3
ah92FJzRD/cq0mP3JIzKqBDQbPEuOdh5xJsTPShpN7s8mFjbJgMmL1KVQaXgmrm1yROT2GP08Cx3
0TgvN1QXA2R2bCPef/uLg2OXJkOBSOOi4kfts0VgkS7mQg1RNnTU6o8j7tBgMDIdTHwG/Ty8Eob+
w6iGOvF4MX1z/loCI3Ypu1JzKtg3+wnKYQrct7xbdJaDseoHUwXkB6sG8ctsIaftyR2d+Ogh/Inz
SrszoqY5JpKlVpIZXZp8gGP4z11Saer7Eu6jbYPV/JfbnCkcXWSNOUaBk2Am2vTkny41bIkDwUI4
e6Qj1N0fgXYHkAX9CQqrfYvXeLtzUc/GY5RYpxCs7cPmDVucUxtz4gXNIFi8XExH0LIuDC+ZWgSm
o6ALMdYyKR/WGO27uORd8nlL6Y7mHpYiES4sNi3K8Agspc/9XgK2l0uO8Lbs1laGZ0MVHSBCI++J
I3cGcm+wG6jIbfFBuLw/E1Xem+r1EtId/s2EeyEBL5pDebmKpHHr7LHdhwGMI4RcsQUi32i1nPNl
dpPwY7DSRm7WS4lZgeDB2eBNaYNkaE5asgulnw20Cy+g1n/F098CO3/uIzcm+b8Y+tdv75Tw6Gby
KHJfE1flKll6c9+FvkGt/uWKwvKMkZBwAdfVNfqRmF0LH8UccJV3Qk/Wu02BN1zi0j7w3Cyy55cY
mag3EAeCTS1SoxHxVqnDD3+49YCnTfgq+0CWOHF1sVXsxuhggAfpFN9XhMPysu2a212mlE3lM6yJ
U/lUJSExP8YVvkuVfR9qRydeBirt13ZYJc+/J/j0oL57hf4GR+X/Gai1VAZAtjUz63H0oFlZh0F9
ASpQFg5zKhpEJiWZdaCCc7n2CZOc11CqCkTaCTSx00klO+qQcBsDGYPI/UDQRUJGcPIyVhPpsDmM
zM4Tra7PuV88gbRpF/Uz2V7pOH2qTeqpEhBW9aKNvCZ4+HQYb52G+88oxfj/FqyIK5LCjI1AY5oy
YqdaecgvlrpwcL7dlpv5PrrY1ldcd3zOTNWzoDiWN0LawDem1oFGPNqkwbLV+XNns9b5BLWrQfKw
dntZSonVGf9kQrASwnTdvfglgVAMkm3mbj/JoFcW/LBQLWS4ErGiv+lx793tYIZmIgjLzihWuKYd
OARkI/twfQB0XO354C+qAySFi24vpVN1AgweAIG+WLeX3DZcKCTe46A3w+ULLXxc1Ng4XzwjJ8Nq
WNxcVL3y+Wu1RiWkjtInXFbGtiEK2w/HHcmoMUcF6I/R8Qqm2xH4f/0dRsby6OTygkKQTdEgWaee
us1FAObD02IBuu+WIpIQCcBgyGHkX1Ff35Fw5GrtEwijo1wfLGLJewuOibBZSZTqgOvH9UOgMr6X
ml3BjmFkGXomxv7+V9gHGScoAt4e4jBS5ysjJ/2IGjh1mbqaLS4oUuP4F5HTez8EdreYlicKAkSw
ShraiZ0Zle8U1EFEKO8MEipGPlZ7+3arm8feRyNhWEl+L/DdMzy8p2HZMHpp/zkDyowbzEZ37sDr
fuumSO8vMLv18/T/Ugj8XxBZqP6V3/MnEhjiyEBgltXSVEoh3Glyrl7BKVGgE2g5jaAFw6oVElxg
Uev57XsoM/ve59DAytFRO3lXIYMGdajxGC7fX7a/jlsscgVX4wsHayX7EGqOWInHpSvqaAYDUtRO
g1ZsIy1R6QEaWS21N6C9VbJOb2higLvImWBzcP1MzEzbPAhn7zoqQ1lJt3Eln0ziJcb3HdfbA7vf
3GSMVfdCDavbtswgkSokzOvyD1nA17KM/Lmu6BYx8OD+0+9VriTl2fsfwxJQAYqb4A4GhI9x2WxN
DbsctHggdauuLAe9DHX1fM9Bxisa/rvZILAU8tzgPS1u2jhsZjC8HKE/PZh9ugPF8M3FjzrcfIlM
QDS+CS6nLhnUU1REj9VhzOs+VNbejexXRwdv/8+BXZPAVuQBXUTmJRdvjXAMexJjErkNmU+DN/jX
s0qRMK7xDZfmJwFXkyVHxzWd9DEJOsnO9bi1yA4EV4POkaKND2mGUCi8DESncisZcLCSR/yWGFzB
I3IYZMJiOJns+KYv6si/Wz1vj7YkNwHDMCNrsni9FE16GnYX1tvQXBXe6R6Wt7gFY/lvDf8A58cg
3QzRDuMdNotetIkbqLv97DNUOt/QSXxVhiZmplMface99/93sVpxz4xYWjHcUfdCC2I+EooKdT/r
b02qt8qeQJNt3w2i8d11KxW8gatdUj4LU0nRH2lowlEvtvos50BRFmUBvJxE3FWIoq5y2UUcQUpt
Qm/4EvfrUzmUtf4WfPvuTBajOQ1UJyCAU01MfnxZwg6S/HwvE1Ix1OYoLcE6zhNxwWCxcpi6sYdL
b1+x7lHAv/XfCIW/JOx1szSkI4cIpYdqKQ8r95Ca7KwwQ+OWTuhi7H5M9JDvP1piZBmGw/TJo1q5
dTNrtSo2dEcpIvnikdAiUcnMN6QSdwocjTta3a48hjvWWzOmQHlSeY/I4GSKhVfvuYS4TET4Q5MO
A/0WJwx1pWYXaw40relCVF0QkOqZX1QrSjr+QcFcpNEFMQSMaFhL00PR1sMEcHrMySRyvyLX+O5z
79vVt7aWAIZlP/A72P7KaWmM+ywAR5+YOGeBKFO/Xuer1jM0Xr7C3Uyl6stlzgohmMoFJWPSpuia
5dphLl7InyCiw4DfCqaceU3IJPKOv5EXuTYw/JF6sUgShDxw8YV0kX+LCPhaWEO2PLWrkYQGYbzo
BaZtQz6o0qYww8jqJYcAsxpVtMShUR2x9lieTDoKb4aaHuR1icl9v03ggcL8ZDYjw6xKPeJs+0Fq
Z4BVEGoJ48whUcprQqtr9jRfjKF9u06DAnH5gyHerIKsLeSNJBXo8scJq6wGMtAKSev03WBVIIq8
AMlB2OGC/PnIQKW7WgxsIrxWgb2JsCk7hTNH2SBBFOFJdPwkANc0cgTHpDz75K56eulAcSNT/nAL
umXRog0KbgRIbE9Q3EHpUSkpBWEKnUDfIpXBNAUMug+lFQSt8+imegrMa3YhiNzFfxnznm7BGhOy
RNK9FhshAAJaePoYJAU6rRxROxvFLfdjAyb/Gnd5uw9t2+82hsyUU+heqAPCkebRj5gpvUL0Le8P
blMM5UqpvKDS8bMLUKP5cW4OEtMC0YJ0lFHIrqqcOzy8/FlmhsVT5Vs0bL+a71bmvDxVjaNBm5zu
T8KEb2E3Kqljzz5XiqjdYJNbV4/qqWswd8Qd9TKm5FfdXbIP8QN1W/3qwT0PKyGGS6ErOWvnpB4l
tVkA3V5h9BQOtRt5Wrna21qbPeTk4yAxXy9n9eW0SF6eES1+qDOik4KtvZoEcB3JMPn2iRSrNM4W
70lQD29pXQ1EvfReuYwo4meTI5DqDPi3i9lR7PBRAPU021PsKKZmiGm5YfIdvP1RwDW2mvWF6pJL
AxMYWhlaeS4KP70qCff+l4rIB/YAU/8/cl2a5/yzTbbL0d0BwuKKbIc3ESBLZMI6FsipBI7M+PL6
SfQM/S2chosHNOGgFWoM9s++QDeLCi43si6MrNqF+vog0hZn30lnvWK1Qf4qpIVu4D1hUlK4wDdH
kLA68EVJ6ttpoj29FM20+W3/CtE31HnUDUgFjOg7cfhCRCd8IuAtCm+DXhKNHxtddwmgCC1v8xvg
zYJfIqiEKJaBhSEBvtlnziti3+wKMg7L1pvWrkA/KPNBq0g4/2/z6hJxLMWUrtqQbEZyMP3ERU9y
eNe2IrjnJ0Ij+N3RnJcdZ5KReuxZ15kxSCu5YGlFd3QSfp7xLNTzv1EhJMyk09/6Tq0CCPtvOZvY
I9NwEDYPZuKGNeR4IGzx8UwrH3p8jX6rXm+tazLkbqLqWpXoKmrEGhIht4VjdCJsfdd3I6hNBptX
dGhxL4PyQES3QHmrSeN/mAYZpVdOlvHDaf7Jc6To0tbepW1aAadiHgF4WvCT6MqCni9AnJHnXMmq
mjgsnyp9g1qBMjT7wtNUt2/0tS/oW120ZWw43l48jvNi2/oJ0QImuTFD7fdM4jWGej0eHc3F+6UF
O7Y82S+5LGosC08OMo5Awr6ScIMCyrABur1UTLH2GG4SC0eAcLdfpp55KHVDEeJWStBh6rKfL6xX
7c8p+OdFffGvCH0XNbB34LQtq8GninjXdURXsGinuPE8Lc/X4r2Lz/uOcU0W74xitqjdqBO4uEsJ
d/Dal9GHzJLjnSvr3AzNK+1CsiPmAAQjdiTubm8QI7tLetNvCa7lgOGsko+UDFzhB6zj7LeBgWIO
SQV/zYmWyUH5G9oLaVjfXJfuLJzFIXAbErvslU6xFsZccv97N1aXcYkRnhLAa34kd64k0TTlsd9M
9ykxPg58a8xeZmxh7XDAseL6fiSUtSKQtgzwhX/GU+MeCW2bB75EOCLKpdf1h8rHrB59gRZVD5g0
Tr+vIGDRGRQVPutp8lk/J4nk6VbwHDdw2/qX/K1snvedvVnGvdgcoQvF0ibIJek9z5g0ZQPSYXGh
TE8Lswo0INcXwOBJDOP4N1oPs8EBp/Nkvlw0rTs5BIg7CUzkgFBTB4INbmo5h2dTKClv0cQE3Nis
V2NzVRiQF0u2EBtCoO8aydYEQvlR7iqChZVHt77rMC0Sp+wiX04yY/CRAL32au8eERBkJE0zopcN
RMBB/tqe3GIbuF+t6HaUJ6y6hOcoip2tPNut2WzXHgznn/4UWuYXMZdIl2W90RXEOwfuUyrozmrq
7k1misBgir4KiA4CqtJl1QOvJkWgc/dLQRXq1VDFrVU9KtRXxPFEuO68YVmk4gE30QP3l3pDgY4I
tLgrdNa4LrlWLp7sIN6QrsvpWM9Wth+ttb9yBWQ8UqzTwvpzl3qqLjWw2e4nB79MqtXISbXWVa9o
3O1DnTOZm8HqRFqP9zVITl4pmJzYoluTDXqvoLBLblZ/d0ePFWAv+Ib/ioBWzbfzByx7X4rMnoUP
f7A0M/WBcwZimjQXq27AN+QExnhUkmE38sp2VDJ3YSOz0Tl+mu+02duTHqHCOL7mMy5iswHWv9Ii
b3t+R5SoNVBdKEogktRLTZw2MVHs/pMAGWKjK1LuZ+/S+xrwyt8G+ozYsiehGL9b50jIeW/vR/Qj
ftsIY6Tf5/XUyboBoyEYnKL49u3p5I1uMnyXzLI0QkzApnkS0qQBY/KNluQLVQkxOj1IeGjIUM1F
oYqCNmH2LHoDnTR6jjIkgto0kUTjT71+D6BTo/2UnM2Fmb2vQdy6RZg9swQ7+Lwexi2BG6L/7CpH
Ym6ARZOTvMhb1ma4LLTaorJiQgeTNrreVavSRpGJZXEeja/iD1OLVQPPzkhyRYP3GeHLehNhRTpu
8FYfZdImfkFxuy43mCNigAkREOfvT8lGk1o1X0HfrpaLgjrHRTM63dLIFuqraLp4xPQNLqKDxY9U
HNX2IzLApXw2UuGoPqYkObhNIXRXRgj5JUALjur2P8a+AaLAQmQJHWmkAwEmxAWmD+oHsbzx8opx
DpSX8dX/tzAo9NdoLYxPK7ed8bRLX2ptpaJ/c6rmsLPsb7xvlK1Iy7ngJJLq6Yu4CpCcCfwZqiKm
wH4Lzi+I2L38RkzhLxoleDAdAsqjqin5G4PZy2N/cTAvBsT1eAnY0VmtUbeT6NVx+pLWf1Q1CUGS
Fd9XPyw7wogYJwg9Dr6/JdnK9pHUz8r66B3ATpxwYIjuwWEWtWQEHa1bBPX1geVjpad5uYjHaIDh
seDYCMijMVB8DZMPEDtSOb4XYTgwRTe6EqRD/qHPZawaIIS8RSUooFZlVvCrMtNyxhx+W8AEu6pa
fpP6VODZH/0OWR6TWsfSex+7eaT9rwt9FBguk1gpsevO+xxDxtNqcXtk6Z0EWk2fjoePlw3B1EwN
w49XiQFzXPZ+SgREobQA99uz+MRQFrNGpyHlxMZSzhhqpOq9hmDh0JAPJvOhM2LhkzghC8hF+wHs
OlHr1+JLhaNzLi9pIVlKgI4ALBEt9DNj3hZrchh+SMZVHbX2kchLPgbMdwJrqaWp8nQS6F3PWa/s
04rzMoF5Cvdf3USk8WeFx1RdF7rXlCF8J9wYtD1Dfx1TxrsNX41V3fQ+LQu6WEKghIKHCoh1hGcQ
x/oAj/ja56W+GNodlKXJ1XWWAMuP98bvqFz1UFxOO8huyU508eZ0dKrr2soHC0gkQM/tsl+rP1Cq
BujMyLTWcBHl5slPtAUUTzXVn9VOHliOUIM3BeWCOEb/q4XL8jyJwTsq2M/WVoIK7gW1T8j04uDM
GjTg6ca2bEitzE6t/ldxJqON7eB7OuA0p3XzMUORXl8TpdlFSvRvdF+LJvCUnB4AMnApmtOJJnwa
pR7JDP8XMrvOVeawfM4j0H1UMPb+9foXP374IszlqJcJ/TgqV6Ek6qRCmHHh345jT5PQXpH2ZaDC
FquO1RXUtLZiPztJdhGKX/EXjnwiJwySL7sYTfb8b3yvjObwVhr21QYAn5A3P7vZoaMWGrI24qQ5
BhXgFQbAIQy1upl5ym7Gy4gTdIv1NSJdIIrO/eFbhXnXC0i1W91+4jkvDS5Ci/Jq/EWoDLkRsGTu
31/M8gt6o6f+zni3mEN7Fl5GlDNkrikr2+oPdI/KonE6VYNSNqbW23j4NsB5Yv4YDQkS/R1/OcB9
cWDP7NhVB0GcyL2bci4uH8IEbh3OX6bX9TSdjoGMNWTCQKJeUA9vliODFrRmNa/Kh1ceK+Rr61Ks
Sz3OXAeV3nsEDDjr33Q2AJlLKYI39FaCBAW8NeieWPppW16YqkJ6Htq6VzTjSLZ7Mbm6lAKXgGdV
wiytMbRiG/SWSlG9t9eYm/kysLrqKLlFkN7dSmVfYvwzCTbmVlVQpdLv9VFEO6k8e7XcD9zwftmQ
yqWsA/WMg7wHT1QQj5n3WuG8G1l8IdqoW2LE7FV9smFddFWDPB6jgnDQOVzj5DTBwG2Zf5bmFkYj
Cckn8CL432T/j3lJ1sbvyoJMLQvKNhB0TCVyQk9TelKq3KXkLxlchE0PPztnl6Lu5ByMOeY5oRFD
G1lt1KDCU81wJltBa7YNiZW6QtsI2Ce35RQszhGOVFbhWkT7fJLWBtJEkLmhqEn/1olhXzXv9xFR
Oyqc1JlD3mT3LDjRgFfClQaovQDAP/3z+tpolsFO0ymCjZ0neCgZpERnRse3cyIx8jEQbX5lu/fh
ZzgJxXkpEAcT/S9Ahc0sS0rb+4GdUmxNDMaTY9LxWpKRy8MxdDKOyvJfdp4mGlpjkXDHgNpCzV+h
pwuoot0LSebFgZMAf9hLnf6phGVbAF1yoKwOXKAhP0W7ponyN4EX+DSqOi57EnEGMsE9PbL6xxhZ
bfOCbqdO66W8K8v17eabXtK/QxFj1Kplx4b7aAZjTfOcLFl811jrOLRUfqKwsNxySz6bT760pg3b
Z6Cmu75B7CSbg9CuoXSONhSn6PeOVaRB+4FTR7jS4wEeZSponE4f6iSHPcrvOcMz5gC11KVWyG6t
XeZRl0cTO09h9IMnnsY9DuIaSemYKr2xXR/MIQ8DScFog5NA0Ic8ecqUO/tcOv0ejFbrlROJznbg
Gf24WTLcFjcXKGiEgz4nPLN3m40H35uahVdqiZVL/1jXucbkChZlG/3iZtGk42YB7Y01D7nqQRw1
LJ0ygFIlxH4DSuXmKPOTa5ZcTMS5gJUMWvV4sjNN84mPEQE8FIpiUqttu9uRx0lGQBEQFCtcNzzl
py3EdYySwZGH6NO91hdrdi8dMbjIOAZIZEyut+vBZE0ZBAV2gtNBkcXZ6RnxA3dxeXdfYwxx2BKp
ExlnR3a4O2CiOmBInzKj7vTVyYLMbyyec/B6b/j2Efy5qC9OmUxFUfeHDsNvP751kdf6sLYdwqVY
lPemlV3JPxt2Lvp2S6wt59iGGoP2WovYqrqrc4DUtF71tjvP6PNd+v/8Htq+4sRXXqf9rdjHoDZA
19no1RFYPZ7moZWUi9CdCTtXwoUs1aJiQS6ZlvklgLuJid7/1mMj0Dl2wIwZvXdpT+eAPzolJB9z
jAB/xwbaBqDSVsIwtHsWPSddqnzxuLdfDn2DS5VE+tWY3NpD1VaSqWxNmPku7d8d9c67q0acuG/y
4dQRFIZVI0GqGSv+2YokPTLOpuGnBr8elj5OY7VMVnSDsAcyZ9eL2nL8+xGnBIyGnhZf1yqituG3
yTdaG2RrCLhddY5GstTBigXl3rFDJHOUwDBLxwtflngjzQ5lKy2G+0lMlyF+7tsWHddmRYVuwljW
HQxLKHE/IETmr+b+URaPV2R/N/4hk/baGcWSxeOtq3+CC4kkrZ9+ngB00zN2hbYSGkLbTXgS56e2
amE9WKX50mroT9S/OTZZnMEPHDjWeARvRveiwprqF5RTAFG/QTMjtlYG1rmsvY46J31Bs1yAh5Vt
0RaCF9ozz+4FlwgNH1P8+S/Z50xVP7oWuD3QlsGz7kdRPN/8fNpKEu80r0bemziqGXf7IP3v4PKB
iCNYcQt92TFwCz2zdoacBDhRTtou73z+AryvJvEi9H2ngnp7tXUbJal8euvHCZaaOagzihOkxGIQ
U5XBv70KmEktOH273tw7E696CEJ4JbYW/OKYTmfE2J+qDDycgUgbDSYnAX+DPUMRsIvG6j4jnh2l
uHagVGcupivzqN4uj5TfrIRPo04KnAWFS0MsrX2srrhpyRzHrQDwaGNOkhEspdyORzDDb2tDxFxg
QRabxQMXcNC7tLvCsCGv4LjWXAMfYYcckmjmCRqTFmt3wY0olv7TREPn+7IcOHBvVLf83IM04SSM
WwWhyuYKKIHu2noEUIKylDi385eZFocHeVvebHTBRmTTk2kjzyLuadFzv2/Gca6S8TGZ18TO96HB
ms9WawVCg8gxgaudEETobQ+nnyKTUOWs+TCy3+Law9bJWwRDFG3mRCic/KuJdzR0QWj6fGANq2ZP
IHsMozobph8tMyMLcQ17lAclGmKRyZT6TX94F0wWNOAXqMqdNjR+OwkKZKGYEHwE7/xUU1HAQ/6Q
WRXOfsja90pUfuMiik0woDwOQF2WLBUnn1yOqyHkGub692xdBlAYMRltl2PgO/BemBL+nOEWNGM8
Gg4QUHTGLBwBDzfVNV94EGUS7YbZnKU+6r3It+3TEqp5kW+n40yLENxKC2j6L6ljYBYuWT5PafB5
JjRU0m1pWuIxdY/UT7L1hFX69+qpISevEWWeoZdy3H5AkHMbkbE8J5s4UYOLk1BSgLSQ+zqFmULk
lnCC54zFu73NIiOju23/AIxjFQuv0VffH2WBkY+LVtk3hJ9qgJHcZvofvgiydYL3okKMJumZmOHe
2NeRrSaYGf+jWfNBXSH/haHnq95ZFBUp6IP/1P1N6SRWkwfPN5B6viM1yP/ISgC6rGX6wNJbMj8+
i8pxFd90XyZYZ+aQ/Acte8ygT9w7Vab/TXfrB5tN2EvIkvWSHbfeh6f9sVi3M0Uc9T4JW6ZuleOG
7FMSQzAYACCcuOr5eFJ+w+Sza2E2/GA4zhG6XtzC3yt/3nuA6HtK/kBsbLT84WraRQmr5FDbslWk
f5pvhZmU013tRx002wsZE9NvyYR36a7EOJMNOIrItHY2n3qycdnntzZKi8VuxiO2z7t5FgiJLLMy
ts9QZ74MMILiYEsfvTLbPCbyg0zyTrgk1LJdGOJAtaKw7laU2ODMHI+fwN234wTrMsZ5WW8fU7w4
9IFVB5vIQpc671prVP/vqpiNulI6J9BXEk3qN3ja7f2MOo3snUzDqaqSqMVat4mlermqeBrV95+0
JsxR5nmGnHRq3pFwSmfrBwH1T80H9TEygnXM5qVOfNK+LArPaUmEMGsRrrzxvDdIfeElNncvYd70
LvmFQ7SxO76YgLwOFZzbNmIwG6zfq/NK1ozc21SkZJgSYtiScty+zXvFKIHUY62RxOmm1dR/9m3n
YldZQJolMjZO0loNbbNVGvzv2XXUBSZdvV+kkJSbpREnMV1CBu+zf4mRfuls/IHagXS3Fafr0cI5
6gBBEGlrv2SZgdDn6YpRgrYw2M6dqabiljIPWLN4bi0dZEfZl7uF59I0AWiTocmg2QffQ4ilG8AP
AZB0okk7uh382Hq1qwhGIUCxiJWxtJ2aWG9BXsef4Ng+6oDJQt7ij7/4cJDVFO2Edbv8IfjjbPGE
eEXEfik1Z4qt+CVCPDeO+OdVKDXXEgaVOLqBAp9yHVgYgO/26BWpTaUYh0GNm9CbINlptsbe2nHQ
ESbw9CS692dhHExuk0raJb9mFHW3y9bSMpCZP226Zi38jBjkA6ks9wqnSof2lP8iHWcz1jxrCWMZ
VAI+bYcqPiwAZ5Wk/jKYsaW2wz8wOMtRiZYqvPbk+wdELMOLZ+Hfth9OBleuMIFDaJuzXCu2rxbg
kG4zrD4AWfjUsQyBPQHemVYbCoKp9605wYk9bGtttnBOL17DKFfvGHSoei2HEB7EyVV+jLFU92dF
4RiElAmy+K5WHH3wzXk57REtJe34DsjeQJoAn6sUXTIswpvl6MZKFrjc//YxFzWTj2mH1ONfIZ2/
9hyJ5taP3Hg0g1e57UMadQ+IhhyP6sflTF77Mabr2I6qp+tJsJRBTmhV2cnRolg/MAAvvxUTK+D8
764J1XC2NVlydH4LE0I31YgcP/DhZedQZiOuUaanNWJFPsIUutkn+x3JJAJoS5uWgJiah52TeGtV
XwqwrtIqF6D9ce6mSnz6lqB0m+rdhoMmAOZ79ineXGzhS/Q9w3rSkGux80LbtlH3Q2LYSfljLELC
AazOtif7fu+HaHZq3kj7gcwXpu8N/O6vOGYv/YGpKELUFCGiHgh651Aa7nln+Qe1AO5/S9XRGTP1
lUOsMbk4fhY0x/gn9VVcp0yxEhLD737hsfiwwsEa2O+gvUwpy4tmf0OA9p8MsbLNxIYhKrODkTw0
upJhMShs1icvyc4WTupyS2LHTxkWSjvVgvtDvuansLWfs6lwNi4GkJ7vRJ6SFKzlJ6rynd/xSq3U
iNiiIXdy2+rLfRiX29fNcsVooo6bcuclp4f/oqZhzh/I4C1cRTL/tgT6dxb09+ar0dH/rOHu8dgd
ocjKEpA8cxeDUbIUVP0i2S2iws0MU5EKk+WRDWBdgfbqduZZjl3nA3idTKmuDqlH1mzmsx0PzsGk
Yzdh+D+enl/Mz6eO7PJPSxjrhWuTxaA+3At0ruDGr+TSNLV8M0YDz2ST+R5+PJU0Hrf274J2pJkg
f/IMSaJU6Vay0a35oln4REVQ/76DXfmT3M59DKgmXeb1XgQDogD/iTXj84n4GtK+alYQgbTiksB4
JOgCCogjUtCjQ/KLWzkAtbFafSTTIqGQYFRTi8z1dqZCl+uLqrIs7KUX/HOlsxTIcHMN5EgRILAu
JwexzLOCmXfXKgtnPkyRFgNFixs0B2SHa3HiZxF7K7n8M5AAPDt9iJFdpH2X3gV5lEJ5v+dI+EHB
9kxCDvWfrnyvLpDBXtPxYRTyR/91qR4DVRomI5dZoYNoDnSVvEiUX6gY8Cbm0FN6X6ABDnEGeGIv
Ws8yoLPheAFg7nBKV+SeEKry9QGkutznAAdqcrnH1ZLYfKEhqH5KRXUBb8CY3Dd4x+XoxkmAnrec
7xq+Ogu8cdyUpDVSpUxnv6M6Mecal/0IA8uNtcVbP3QXMis6+w8YgCUPkFi/au6JluHdwm4Z124l
27cwQQr+j32uMVjuGS6wTVm/HZXh3PQHftSwZbxm7vzv59MwNL6RoY5j3JvTut5hoemwlEWFJO+7
LGuDRbeugSF26NpOWHU1EXEemSOC4BeInKIRLpwL6tR7mxhGJCDOgxoBwYbcIVyBtDDbi1+Vx0wI
fyu0GTDH/kr9zrqKGsabsaxB5qmQ50RftZCQ3HSyCulysVkz2uhqVMnre+hXdSpULNCdi4nhcANY
FU4T1A3xVaPwF5Dvw5QiA+y7OetBH3gHj/FUXyxyN/NG4RK/aeIvogJrvk7IC3bZsUIi0SK3i2G9
F5CUwc1jljq6dMkpDo39iFZKX34HhnghffVE7Zahuez+14Ya01fJ2jjz4ckqlrdG+jFs7ftY5ghe
Y7gT2R+2V/cWXrj5pBNZEl/NP4esMwNmqIwSfM7WIJxMB9pAl71W31CWyp7aPonjStqwy/4gCPM0
8QW/qLkZwzh8C1SblFHRQzQaHpfnue5u/TdkmKG9c0ixBua8ws5HPQeGNnt5UYsP2CV9oolRwqd6
hKUKqhz2V/B/wl+ybSLVKKxU9y8/c0c+OgM8fsoYPbY9Yj20A8fe9B1L6+QYv9DXazsqV9czeH7R
WrMAjNDyocduy060e+CU5ei4g9Va2mdZzbPfdCY7qu72bNdvFMB+DpaUXb3s32mlG2MN5QgtMHhG
WdRefDpnz2zfSzaBogavKfFKnT634Vn7S3vBA1PJDQ7qJF+0uMnskJGkpoDH3o6CLgAu14IONpT8
BDxrYcIddnTm46mcAZ+11k/3sXQwaEcV8ln5AHsqoRCIMYyK7C3tXrMQ1tyDWq/Pe93ln4IQr70K
m2CJGq5wN5Dk6Uhx+Ui6xdSYbNJac2Ri/15oTGthEnED3QacFcBHfurVeNzRO3qjoUJXwy4OBbbN
8FWpmEJUDCuXXE0Z2fXnamQ4OIhTECU7emjIHQWwa+G/L69IPhhl1w/0gn/mF0BYvqr1IAe9tEGz
TsDvNBjMbmRJwyZpoo/pb+fjF+Fn7o46VIh0ZwxdhqI0RlJDtq+xtb6fB/f1kXK29V93LT8LobFT
pRZD3ZzH/AhTfemA97wHbYUfgmvz7XA9txVIyRMefV4/9mMTKK7F4uhk5Pxj50wcTwcEuV2P+YrF
8Uj+28NVzAY7b22B7DV0ISe4s3YPi37w7XllDRyOxGd3EC3WZitCRVnk9ilwfIVvnu614jy/utDD
lm+jzp0VoRW36xzLrOmA7lG0XoXHbQK/+RU2Zk2acfodPBqsTkVdUj04+WeJQFcfKssUfWf3RNCt
yLzjZ/aPtctufDgqvtVOGza5qwWt+r+G0P+4vPaR0Yya10nT5PQ01Jnowa65TB0il6SUtFRx7IL4
Bx/vm7PUJTuSwGvwBfd1zgcXZ+JRy/o2yCvzxuhQlIEGjkQjsT2ifGyeA9IkIaeaMBzes7KVON8E
AvtVcGY323ntK8Ac2jHpIxDzqgGquHSMYNqlpJmDwofhHlh50IRnm8rNkz7WCPYee7G9PbuwKial
OIIuAz0kYtbFdsyraqR2nCku49qCnRmwUVH2l3qML234bcDPZdT/HXRAxqQ31gjAaPqjmP+FdSFS
G3kf4/vQDxwEjIKnTSSJFJBOd+eRNluyFEpZ12BFrVdIz5FAgtX07BDqpcRwl/Vlg1ZqYwFgdYwh
gk91KNEy3reZ5EYE4IBQ9FM4gzjCj8nj3a3j7IiUGQC5GU+5M78Pgs+Wh0/4icIoHNrfMeUHOFmX
PZfeCbb0lKB7LsvFBjVVA45mCLGB68PAR4I5M+bVLsyK3FstGxsCkRzhxTDpfC5L4Cn0hTA8OmRk
k2hzkj/kFx29C9KK50DtryqDZ0Fjc2zGyqDR2xrhXjHjuLsxGT2BUeK1K/gOJqMMMrDoeZXy4qg9
FaXLKrn8e8iUvgG3Pbz+tVIEzcS6vHZJV7hgCz8XF1boe4y1DgAJXU3dBEDGs2gM/9NozDicRs+B
V3HOqfK4KKn4FReCxalPwUY43n8RaLxxs7wwIrHhX1yFoccAiZIt8gfApxx9ho81NiiGlqXQc5/m
w4DodUlwbMwIhJ2wo9wxuhW5xhyM+0naK2o7cSvkqp9dJX45VWhGza26p7cW4FzAoq6qYQHjyzXm
WLveOfqrVl4okwphfE/8MTe0c8NI5eVweRFk+tvjWb7etNlEkZrwMb60GOea16dmZ0x0Uwdu7QiZ
G7mc2ZK22sIi1ZjKvHgFJIxriFTbZtUMDlAzgxqXpiS/pfh3KaRgL31ibwiYgFkv6LyQjHRozgje
LAqxo+Q8Vd3uQW4vDPuftXV5G1MJGHFkr5QIWS+lbOpwKNCN6P4pyyGd/h4QXyElI5zviMVpW8uq
s7au6GcEn+P5eDnAoVY8LtgN6124UX43WZF1ISMRDrEX7DafH0HXZbgD5cv2qSygfbqW2ieaRXFy
jSNBlgz78Z/LHQsGMkFf87su9Uwak/Ium+2ECS2YBsq9cNIICQKntIpV5+MKTgsFz6H0d+adWCIB
KXddIIJAlsDl9ODOjpFNMYjuNvY6LUg6uWA8X1j9Wlyx8KR247ShxJNRJmFptsama4cbHjGD55uK
IMkAdz5qc1PQSW7o66Aqw+R2YIcKYpXAk0TtFyXEiRd04NncgNHr7MIUGGe4pp4QKS/IzQz0VqTX
IBUsR2XIzMaPsVkNIaXTtTMmMiKWyapGbDebzCo0LLsBZnuh/feXinBnKgsKqk0r/xriOelf0WzG
10ul3CQnzgWfrLwwRLp5jluI2K3wrEHOvlqsy/f3Mcq8UF3oKAY9CvQKlpR1ZmLE+VKEF6mxJF9M
enum94CZf+aSYGuCKtob59xOUw3AAi2u33cJwzbfFgq7kBSsFcIVuyBGIVhnnuB5n/s9NSCypUcZ
dIkbSy8X4bGOaT7/ayDQzaEWIisg1+jZP5iGUWXnybvZ5v3V7YPAQigWMAHMR7tReGXARa0KNcz0
rx/1ueN8dxOSYD2OYyFoJD8Oxm7k3b9Y38akGbi3UkP+5SwffnYfKOHvGJ0KtiJc6pqMFCelSi1w
ODnA8az7dQ9x9uutpvQMIdt20YJT5hSfgVN5+DHr1ZibVLZPrHizm6cNosM6m5oQGxabEwO4VpwU
gWql0ERCovrnimRqpCIgPsrY3djDe+v/HU6HnoyPStzT8HjZxiCImuruBsMrw459K2KhilG1AjPi
QJZ7qi+zafLfqi7O43DBbB1CUpkJ3Paqfp4xon2KhNRaVHoVnoTEewUDWTQD7irw04zKdEKq+o9G
a+nu5URlITQqHQds+k0BU4tKlSs4+8pyWtb+kfSOmzfj/WthQ2QUfkutVmoWEHWwYq9Mg9qn7M0J
YijXmyqCOOO34l+xz8CfktBLOAWxkphF2x9sFbrahLaCFJu5gm4jh4EuLIXynPWZOOb77FgXKx9P
jFNEl3hSRk0MjpmY/HVj1g64BTqVZeQJ/a6Lkek+bmsFuEzMfEVlU1vUsaRPHG+KHFspeDokiO7T
yAwkiSlAsa3dj0on37T1uNaPinWux0xcYoRqghrzrq4Z+Fzis2iLG4ugD3XEuf0O/t30zWdGrqjz
pisQOMJ9uUZ4jDjrq9T7+c2/CwcpetsHjYZd16PEqbHNsbb11pKLpCce6cfxiRtGwnbhzk0f/+Sc
TpBgXGSyTsf0TvmPZyq620HJwTgnzxALRWvWoBcL6VswnZQe/EJ/YDVjkrD2c3/oE03WbruHHs8a
0rpLTrwBVaFhIGW9ZuUE1ZiWKCVWNrwOMAYeg+APnFuHSvgu6N4m6khpCl/Kr7x9xDi8uWYCokkk
rbjNlxL3U2g/4t8UOjwI9ijw6j0Cvr4J/fkP7DRMCf2yRqxPGjqgzJGDbUKftKgVXHcQ7OamXQS6
cp+W1pMQsoHZpnz7xoawzy379hDPhtu7WJhKgpvmwiOYA2bSTJUAtZPki2brNaRLpAngDf2Lyu44
NaPE/EqacG6VsWDvbrQ8EQ/YCTnpyIR2e1tkf7RSp0YWuiZTZKFD7xhLUyWTjgxD3fZeL15pN45R
ofRmLqrjnR7Uk7nZu0MWkjtrCkNsrl5ap1FKrD3lZSMZPBrL6Z5Vta0zWUgyzASpzIS05vEsf50r
ldn4yXIdE4OCxxEkLCU0srTjFREFqh46PAoqh/FPzXtG9ePoRm7eDG0F9RhIFqyojkUUuAKlPsoe
Jq+wtv1RAxH5AZNRNb8CUgLHgnyq0xpFopPjxpxz858y240PraO9MoGAHyGD+Jo5WOLPYOMo75Gg
YGsO7ch5ldDQxrfxMlYU+/h6BXcq5s06UnaxOIXpdhWlXRBUmwjCglSAz+SPaXXRVtQ/85p9QGot
ee5F2YONwIixG9qY+uEjatmjhSLGTRsh46QQ11GlbMyEScs4qIqZWT0u5hrS8IJ1+W4BIjrkE4gW
VSr6G0NuYwTGDvQKH3OZMGbVjg9rlQuyUqCsaObAnrSpqUf20g0LZjtj1q2l0c491zh4mEqYCazF
g7Yun7YR0/MH4wa0I2QcI+UBkSyjJPgINFQ9TaP0BNi6pYEc2dS1k9l1on4qGOjaqJ1zaYP4LOao
COki4sEBMcDpOWKN1smwnScQUZTGBymizM3z93ztWwXCX0n8f6HMBFFrqwrir6Z+AU+V21uqw3nz
xyP+WuFofrGtX9PzCbQMkVK40BvLkNc+5bF3KoCaFnHlD9POGRk42vcnuLCn6kmCTdauvBX9kQfL
rFrAJcH+wsj4XFcIj1/ga5dz7kA7HO2bcP+OVGD/VdKw5XVlPzUtcushXNc6dUY+fj6hjOt8/N+q
ny4B1BAso6dXyLldYJSfOYrxTLTo6DItWnFouQuuaeBjHmYv4GfwZerAJFwFJb+rmJ/SlJHkK6cy
vxUtrfWVyvzG2X324WySm723j3pUcb0mFIbRwuHCIRYvwCWl7HZ2tvEm7T9gdoaLfT/LGMFkGjOQ
zBfJMlWR+0uyyOb3M/jSiecVmLx59gZmns0El6IiiG6U9dw5FeSiAq1F7Fv0QAyyRu9Sc6YveOrf
X1e8xIToVceiEBuRLtUs5hnwwh/meepxZt7EIgd1fliuNSwAygqT+JQZHoyR17GqosaxD3NQMbXH
OIrTD8cR1TeYosXj8agrbYigCuqJ9rTpgCdN7xINAGtI+4VUCzEmf6TeW0DoWP816fB+xH7Go5IC
V0qHbWfYmVhOOAgMdEpTvZgDu43Ml9661FwwQPk42yQmwxf7m60nCS3X99/vvkhIP9jXiYiaW9xk
OrB+FxOkuaIMbmSEmCyHyLzVORyeLVcuLPbZrWIBflGNlRTHSkjr6ClZ3nN8vFI6S1VzqpYheq4W
efdZYsEQYjNIJ3gMFZK0ObuvytKamJYNajl/0F68KM0Y5b7NEy1qudif0zypZJX3bHK8TYu+mnNo
oyi4GWjyBDoSkGEjLjAiRMlaJzockSimobq3zzmaHkvftlsGqOxYVVgqSmyRDaDXUIcLfHoiJOzq
KRxhvvnlvbIwvWGXmrLcu4r1oGsQzg/CJFscuTi/CDhz9exJE0RVL1Gw1iY81UYbfqZhRjWoqqy6
FOotiLNI4pymAjboNKOSi9r3JuTUcrMoalEDNC2tDn0+lOGeKC5zBflqeObyZuVjgw9rc49N5rYF
4tlqMn96CYBeBTjHZlkQckT++VF4mwa8mByfxilVeu0T8cn/SAsT3XcSGnEx0jbJ1X2J/M/dSREs
KzEsSWSPJXK1UE4vJTeF7t3oqZrIcLcLsacdJyhytI1uGwZ2fVaIdORjSIla9BSyt2tHorMJMLyK
WKUZWy+h0acoq/CZBHvqytO5lors3YbcSPJh9lSOcC4pmoyFX1NYeA7hST4PURIAHzNWdtovw1hi
bzkaFWN96YibeLk9sAY/oIGrAmTdfIGktZkaJ01QEYLub0haSiW5lgvHbR+DqzK2xAfhQdTRMjIc
o6s54WSvVgqYd1wODFeg2SPQxgqRstWvtRWmSaqVWlIg/TsGikHnKwZW3JtvkCwo2NhtGDxyrqcL
9saVvXa11sr8JhQomuWE0ubKXICMQQ1je3ZjZR+hWNdiqqEbd0uRngadeT9OOlAZh6JOY1LIygDW
uWzv/3yd8Yx+ZyxL7qjkCIwN1zYR+8t6JTzxiXy9xA6WFVsRm7TcjTaCP4mKbMwa0sw9VHkCnR26
yJQ6QujNjd00qAMqrrXZLWfQbvpo+q0I4j6A4w1zjLruhm46dldcLEM5gWk532kpdkKC1fns9tht
7FPIp8gXUCeSgPaiL/2dtCHq4XQjMFQCSR97ixtYA6kL6xK4K1HDmeXxNqUlnEoaBX45/EAdWV+/
hPJxjbjuv5oR3n/B5OtuNH6xOgxP5l03L/hWrWVVepNC3oyRMQNAHhx09S4IVZhUNyOuG+dxxKvB
ItGftM0+kKtUjQGk9tk07iN6kN7Xyf0pDSHBkEQrpbdE1bjdngV+Yy2rTDfDKkTmk2ool4UfNZix
t9Fe8dbb1A2Q2KEUoO0Pmrkx4ZAQP/Zb4TXkWcmTFc0vUkBLiU6Uu+g4BEjQa50FMe4Qf8lKLD9k
+QK8XUK4a1nsAz54bh47pLRdnqHU4vVkBEkHNF2bWQDhyBbrnvvxAf1mG78HlPkb93ujHlexKyOc
7F7nkehcXI/4GTvX1gb9ksHC5qnG2eJCPImRaPsdvWQo7X5YI8i11McrWZAWaCc/MsdQovWx6/7J
/VJuhiNR/HvjVqlGY+6tSOhte503GFSu+mXHs261yPGsDjAyshs43ZmGH8KLvMsIloNeR8euigla
kQviYac8c2WZNJy9OLRi0KPVQVaicgH7WJR2qhZmnQiRQ6f0uuLYUiTJ3BUtIc7NjcFFNFvt7GEB
o5unjyYbWPKYH1CGnnHc/vXviWeISGyh/zDCQ3w2HNeINoP2PcsqaNxnNo0pkNK+ohTRweuxOszc
eOgF3CFKSwcmd5Co93djEFD61zVz0EUgbBIu0aNDYjqbU3HFERGg1k2CH+khHAUdz6TURc+eJ6IK
S6TZv8sAZHpZGjGJHUnaF2IlkBR5IOl8iUjkue54komvMcclTnNAqeNsSqJRg2uifivlI1/ESEtX
XFU+UKS9mGbTi5ZKt7DK0KMts8mN1dTdAM2FkytP+gOPwdgykL+AvMLzQ1jkA/ydGQNeA2IOEnZf
UGvm81ihWIiKFEBO+m/RM3YiDk2i01GDCUmSnyXCMuPUuSqSuU11yi26Nylnxw7dHNmJeFSIP57c
DOQqpdCUJxF09LYbSwTWfh1tgqS4dLU2XfZCReRWSeo4vScWCaFo/pJ9lPZVoZSyQoPCRpdKLqhP
sVZLeXeFQ/7QWvGT7zxS5gNEmFVTQJCp9AqUrrKCeyI/fx3PPgRhT4//ZGyugfv3scGKtgdhx5/B
aeOhypPCY3Efg8MJPtFWuRcynwAAK6jEL7uIzWWZpsdQVa0YF5QvK1hHhlrhw9A791LzRzixLqzM
hCvrxb3UqomE/HKGYcf1+7LD2NAdjf2uL6YXLuWiWbHYwbgFdKT3R6lXsrRbU8e7h/d0l1G9agHy
wAoDe28UvXr6me6GdsTOq3h1wJvTcSlM9HavhR6GenBHYQZJPllPkQGrpcDB13Hb394ztR3zUGGT
uOSrf1R4Mw+ffxbOzhYdCyBLzRigv3wjd9NfKJwgA3td3nnPjPvtY3ajAfDf7XDnN3gZEq89iz3v
R6LeG2XfaLxERZ5CeLXIh2RwDZEM2zw5ed6TpBN4ZdBdXIvOcUVIkvOEr6HVlRAwTxpEpSsvGPHI
6MsYACT6YpN4Lyvc3qL01owIxlY1s+98EeIgdlww+F/RaHaImTv7eEn0RGWCsDWkNx7/gDDF9Pmy
gy+DeG4IHTksVYwLKTfldghfNFJ/P0iH3lZODTNI8RZpPrb2Gf0rT4N+2maudp8gIJVISW7uiQLR
TzFOP9cSEP2hacwVXS3vHmuC5jpniGArBUCv9j0wGcA/SJpJN406I6qenK0Jq0kBQmoXHfdXd1iE
UNAoZ+cUJ4rPNjqdiCEylwGsJcRp2ab+QfgflxWouYBPXnT3H5mWxWZ6wyuV/qnCLEWHDLRdJu0i
Yf7yi6tcy5UwdD6kUPv0L0HzT/ebQ6A9U4aDveKlCByBUpBWQ9a2QyYvuqNGxbalCN7RoHRhqrTu
xnsCyGDShoGw1e7MBEO8U42q8ebSQvswCBcVdBrTOwtxbz7qByzomqmeYwTg7m/gK9fE2I/2JRUQ
rFkaBxPOzg/AwGIZEFST9Oop/CpWUXQ/eJM48Whm6k2dC6xUvJiVVnbTwknvTatt+pK4ALvw0JL7
a3qoVNXXnuv7rsfLRcKQaQvoIYLJ1Qs1VKCQ/N4WMrcK4zPed0eTz0R8eYUrSvdPhBUc6ljhLHUy
nRIFivwWBWq+OakyelLI7mUgZ9zZSBmwpGO4eg2fyNxMMDYmZzGIQn31Sgb9sjJEr+7yDTJx3vK5
GSu2WQtGlwbJzRUBvx8xfNde3nVeUWEW9EUae+5s/KfFuxTTaiTJAEkzpPmAspns6t84ES6753Ql
Vfkn1a+ZrR1qv2V2+nd0W7iOZW8DD3j7tC+fqyzVndxMVtoAByjF375VNlqSxb61yJFPLCpOfvjN
4W8/VOETW5MI6tmX3p+IY6bZYdRHE36qA2F7eHR8qJkD85fvFPqooC3sGONS/+lR68tD/u7WlpPr
6DJcSGqFwu4EKBCBJheV0Haj5iM4EitchCRPF871Hd2ayOopkENqXRTbMxRcPT48ThjqBPy26jzY
IxgRpAN6s7hRhe6cjC9xEokP2JKp79ZdxOxYS9uPNfGp75Mo2obXk/kXAzfnvKvUPzsbv5ELJpbI
gHJsi0scIq9IF9xcnYNhsY0bptEMsSR6qbFy9cD+6/IB8zGxIQ65/cf2Zh/pyXdeJcdm5Tf2JUUq
EoVhFmWDXdu9y0t9rWpfeA9/qkqBfQnbMBkeN9bszbZeynAveuXgBQl/t/Wfa1pJeE3G7D0eqPhZ
/aKcXp1ig+P4xLcQKaKsCeUpkPIr5Jj6Hx3homPSDdz84G+HKhuHz8Cu/lj5IGahfOcbb/FzdwTE
i0EtC0KcMYpNMMwqtpR+HCKM01GbyA2wjSiCB/zW8rhUnqaAVXrTRRnd3LSsdCUNMldJrXHpBxxw
9s0Mrdfr4NHPfr8dQEgMTirciSVBJZR+89X5ZdHA/IL11UMNq/5RnQg8wBcU59rtAaYy8szcvnNY
2rKsdJidv6nD529FKqQKq2TI7TKtQBkyW6+aEyq9himNn5OmcsLwh3ie2DH3zn9D+rRL0IOV/ymU
1hGJpM3uwnGSkU0KzeqtQcmvS6jBvCZhjZZM+j+ranL3iSdpc7GvpONULLrY5a749aiihPjXvWk5
nj8JruhoUHjxn+qm53DQzg6honmFyCTdgnfKvndh14qMgVpX3bFjN7yFNjOcvkYEiFs7SnDslle+
+peLaAd8B/IDYdiCfozFS6anH4YCH7VREl5kAPiHRifaxxwEgAf0Qs3d9LfoM4dRBlSXlEtl0sfm
MfD1eUw1Hpt1xsT1dbiKPYesg6borLwHBYJa4N0PakVsTSpigRciLqC7lwiXk9Dp6OPCPhFYjdjK
A+E3BlMVPal8Ip2IdmKlv9NZRYBhFt/r6t28SKKb2DlfKHNPb+XYNs22EJFoGZc7lDe4w7wL1vQ6
BEcAVlJGBfnYQknpnwP8r55X4i+kSojulrAE09C6o81FGUuY1OhK4jIEJPp1oXKFKncoYGukYmOR
SKMjyIxltoZHQIXZCreZ/1XxHID+pL5iIBwyKh99FPo/ksm9RL7OOWLYc+O8rwEGZcYr0ifkZCIp
0IfEuJxVdWr3aQJ+I3jopEgqUYGBWz2k5SPp52zyRyHq9zRnNe0aLVdBWo/rgSJbIPjUidbh8S60
bvS6gM0Nxwhk6M3F1iTLYd4lWsEa9E1qwtHbdwHBxeswOQqgeHc/N3m7i+jjbHvPpoKnFyetjSZG
qEFsj3BdWYFWJ40VZLakaBO8txbBqyafkSyWiGgHBkpntNDeMzgxTV13HOF21/RRCaC33cnbShsu
+QN16aj08VGXhOEOB+JvUBI38LezNz+6dkiou4NwlFaKYsk8R5UiYspBnTINpqyS7c1YpTg7mrfX
G4iOSAuTbaFDQmtjvAgA9y1YU9iIs05kaBKRDIokOk9JYczE3RrUSYYAxFfBzPorhU1RtmNy4jqX
kyEm6WGAK5t6sHmx5rqCEf80F2m0WKj8l+Uni8VL8O41+tsS/esbSB4NmG+J89HAw55f9c+UClFE
Mppjmzgz2LNq6w58mCY+1tV60tRZETQY/69qj7IyUlIM6lQNBgAmhN7gLuBjtNGhSBQCuQ2bel0N
muwjlrH9JrEo7EJipiBymoXMpzJwrWlcSj34v07mm4l7Yj/rno2qBp3sRi3K1TZ3afcH+CeMk4S+
HSfyOBOfnNCpnx2xq8Ye0OgwCdDqq2UQSDY5K7+3695dyvNbExCtaV32ZrwpwvmOjvbrZBk/6jDb
36JLo/jg7ymyYKuAuhiidvO+IX5bRds22H351kQMo88zAUeQ8ZJx05Ew9NprNFltEBP4eob8iTb9
TEQlz3/6hApmMKrgWQFG1Gc/Dz6fTE5BmLq2Ha50LGQyKe4Ss2Djlqcapd09u1TVDxL6zrzt+eqY
EVNKg3IoQRygbvVKDo9N/hZjSJCpw5PzstPXRiqbdDByOYgKl2qhlzeN67ShH+tReFImKuuomL78
jM35A1vrAoK7COlwp1UlI7a/zk3Hf6ZAXqyQCo1DifMuiU3Vwomh1q31AjCIj8efUB7kwlFlJA8N
1GARqlGUDJyojlXuwzycPLH2ds1q1cJ6i575m19DtWugc5DwUs8fwioQrhsQkPiovs8Di5OEsHKN
OYCnTHnSxlEd8M/hbJFqzw2XEMFJc0fHO07GXc8vrlfs0oinxpnvAdyMqVn2nTEVnsT4RhlSqSQr
AABYKu3NbWfK9lbK7S3X6V3lwCgx9+Xn0oBEIbcXigoa5UXq/9aJBDsZZa9HNBz9xCdNjpavDN+K
Ft0cvZrwNkPXh1fNZCo/KE8BmuSOZ7vluF7OnYNItPGeBJAwjLTGzbnmqX1w1nwRKl0ZBNbLF73l
sKC7OYfpQCO7RnFUaVwMk62n5zq2OBGQ7uxgs5PB14gOOXf2NvwicacyxmF9ckL2R2ZkhSGp3BO3
sLrBFL26/yotESN2yCUssdnIOC8/M6/6/33c9BQvEYnuic+2EGhdX8G063Rby7o4y8z6/Aldao8v
aDge6I6eAzNuHJvjpto/A26gQlA+NRnUUtwtvX/LplrW/GXzzSbxiSrFnAObl2Tl68nIopCz9et2
YCVvtj4ENVqG74b2HZw1jmbe7NOwB2cjf3FdX6K4Wy02bf/jme9yWrFQCuPO236at2LKaXmzpz/H
38zKk5oTrGzWQH/cgZ1OOoPh+1EqxOeoMs7kpUe7/KP40Ze/ICpo65DDh2wHzpd+NJGwV4sg6r7U
cIxBMrh1plL2xg0tERraVmXXIfRsZujEVPve6EDWsfxZi8SYnYYzsn3SFnWKc4B4GZB6Wn+9hPG6
KNL6PqcFk2Hp2AJiK3BzoVQK6I141Z4WcswXgOM/ctfjYnYEhuC8/LwyzW4PKsgXa39GHac5Abgw
hKEqlvKH1xfs8f9KOKNULZJTxTMxWWZPm+ryUgpkmoiCpJ1jpEj0bV7uu3OyL0+d0/5xAsPRJlON
PlbU3ne59DROAH9XvWe+ma+4mMcfK74e+0QOdxFHBW3x5xiZmPUX1aowJ53TT++KKi05blMN5SB4
ZX5tWWqQHCtsaXOtz9CmOFJEGWINKvzdoDUdBGFR0BlDrwaENCBWJkSLHYiFWIsZ+ejR45aOlZEw
DyxCybpiItB6vT4SaASru7aL9O2F7/UOn6n8sDP9C9sanl3WBKSUi6ESYKjwOqxkgvIcFeENoOam
pq8TkdzcJyuqRSJXNvlZm6LkvslrWJI4uBEbGO1aANbpDtKZiJg/FkRVevQK0dlaRCBuXHWNrrO3
tzRhcyPqxUebVo0mroTTejW6sAqdSDz8h2IToATuoM0/KIKsQPm1YgOVnn6yjGuWl3HIUN9zU6il
uTu4gNDIfZZe80a5AsN44Hxq93BarYEnYC+wBxC6OdGNEoEr3kwdWz6zJG9mzUsCjbj5jKE0XsGq
XVm+gjBt0RdRd6ljAot2k89NfelIJbWMuVIACpagco3oka7lvdESMI0uXQ63xHNYMO+hZkhUumMk
Z0jREJIBSokjciLrgMZvHjNU6L8aIuY41+01HTdZ3SkCcNlsJSOzLglSr+hDvYuciFmIUyV/g9mY
ZXji07s85Jteer9he0ip1nAlEt9i/J7hkWlQgR8OzIUx/wq+uD36aiOD6JIXW6nZzXuNg957INWH
YqEekK3m8jXy+zHPDME4M653MFxwn4LVuoTAfpNaEsyq8FMFPMPCuoKrYHxB8hj07f769N/etl5Y
Q0nK9whGlr3e47UigSompsp8aP7tppGjPnPC+NoZ29fev+46RVhkWZLeG6g5i3hrMg/9ul3KhOha
SZYeufsaHzhNc/DGkFZhLIvKCVj3oN+88e3zCJaVeIBAyGmoHEP6AP75Fml89BFtcyZl5IhmFdEB
Fzu3s90jdXwJWKgu1UtYHple/E6K4r4b5K7yW4HfNano+su5R16jxMv3jgfvLsa9aUtUVMZ7QH1u
4+Jesu8/tam6c1u2ZvTfJwECjz3IUdWrV0lIEde+1UFmjA1KgEDLM03a/gt/DM7TwZwLNwgHuRml
VfFpQFkH8PDTwXOEr93R8jdLl8m7ED7QuxlEL8AAWSw4cYAJvQKqFmDd995yRYD8DCLd0C9GPwC+
4WhyQ6EE904PiONxZHJIo3Stndwt1TEYmq5/IyBdeLjKWa9zwriKpbXYMQvElqqUdQ3p5MGP7UE+
w+Lj2vlwi69W+l0UweaAvHYs0x/aXpgzLneSMDh8NVO1HBCyMU+8FrO7hPVr0sTccqYX94VHq1fQ
YprPoYzrjGAxl+PN9dr+jfzEkxz+3KRP5ghdDNcIfnwKEvjAFwYy/l2bJlwe+3oxdh/Vi+W7bgkU
Pvc+4Ab5zhxIliB5GzaojtCNYyu0RWjAa80ZZjEay9XpwGFYdHlRM7bvq6+03fIFuqDlXLHFTnxz
Bf83Nb4jBXWfiKXYm/99gbKHWU29n0oly7ytsHT8lbLCi7sMiSBiwHbQ4dHWYKkp4eurAHoxnL/B
h3N8RJg1+Snmclp/smdSEM34sLWnPrUwo79YZXUEI/bn/VVJtqo0YkYCLZRj2eiKziCZM1/3JtaL
duqD8ycLZ00XVWbfLtU7wEJUZ4hkYmZAhaijYHvSkya6zBBHL1qsYRHNGoNKW6U82MDF1IySjVtA
5fiD3jPEuOPyhCDS6jofyj97/IEirM1xkYLg3tUDG+ReQ3on+x1zK3vqzhiMjLtrtnveNhBZNZKE
12MmCANrbj18lHQij2kKSg9zIWp9KhshAl71afb+K1sdw073AleXvzWqsOL0fJET34xv1Avn2S1W
GjEhoSllyzWwaU20hGRczx14Sdvecib/jYxdli0x2+3vqVulNlfqNtP22Tg83GRX7RScp67vd4jX
pdlYg35uSt7Hh+YptHAs/eHlgEV1sjy1RN+Fyjwb6u30P2S6O1xyzVTaaI1EBsuFG7v9ZefquCgo
ypDpcoFg2yTfobrxRsSqqM+Gvy8I41RTYzAOn6sblghni/0dPdS+BTBGHHMVXE2EFp6Bf24KYw3c
T2xXCwnY3V6iLTcCbitL/1g3QbVIbAWULophvkrPqyFH1DRzJo/Yp6kAqIpve1YhhRIDRjo76pbp
XEMd3qXlm+hk2llFv3jc/Mej8WfFO6HILi2O2fQ4PpF9AW7hIH0wJwUfDV0h2stopWKcZSBWKPvd
MrYHiZc0lLJqQfo5GKu7m5JjOCCAPvotCwb5xeQCl1yhbVkMUvaXHP7ErZVNMeqwbvWmaHoy475h
ZjxJeTcSVSp7aDrDlaVtXvQFX320/pGtqgcFhjfE+WLwGe15hQy9faJbijIORtHmRlZA8Nirtww5
4QDdVXkO4mgGAFmNvRBWJv/NOwTwWsKZbJWzUMCtQVwCFx7Pli45i2wB4FluPXMWy6aYknG2J8Id
EL/nJ5XjUHGZlifXpguv8nBT1u+ZBp3GRApfaulz6pQ2IV457TswSvalDktVb94R9bdZdOXCG1ey
nURWZkR40D+SmWP0e5UqhQ3Mb691tjlCejQsrY9yQA5RV7Ys2JfBmkxDL5lwDbEffy94mGRpJ6DV
mH3khfk50pUVwH2B02RVnY2p/yzvnh20qVDLy2fRuJQ717f+dFM8l0YVhWwqy63cRuK73zl2IfA8
Wiyp1A5vHpUXewaxitJPSLzvufv4vzKI4wAylunqS7GqM8hzFRKkwf6/tUTeTxtW6X1RGhGbtpFi
InTBnKvdt94aqnOSsVgRILAUi8nXtQvvO6umNdFaxGKqXNWXUFDjrppxDEUNuoCr53Zru4TcaN3f
MeLFqQyPFmst39Km3FG2sv7jytPEmgA2tDjnIX4qAyfTtxrdLyb6DGYbYF2cTiKBUFJdnvp/7i35
ndPujr88MTWLVd3FEJ4NxkTJtpNsPuki6DTK/pGro8bLtlD5F1w96gQ7zhzuRM8Klkg1J65hD2Um
oXV0ILMAiDJdMsmXuZ9h9DzafofLe2bg3C7M1e7bZkLyN5r1AepWOtWO5dbdDIrZjlWkR7BeqvZr
6l1Pc5imjiqttcfdXZ9txatvuXAo9UFZnIPZFBoNnmDE7YTeE4OfhcOtB7PXUqzD2d+aq7ia+IdX
3Ftrlt7rVPyXF0uM/+zOBDjOcoAYg6n25MqIcr4X0+2DQeoftEXnNVwJb2yUrm+oXQWtEWq9SzrN
ounscwCSiwmDst+ISBP3vYJoPHfwlIn1vbovz09FsXClVjCuTh3G8D/0LIt+SXA6qX1JnQAXS3et
Ec5PsopkBM0Pwzzt0HaUUwypmK5qJ1NtZdgNy9pHU+5h8PeEtlc0U1h03aNzMOfrep7SuC2KK1i8
U9OHyc+O2EdS+5TXyf2dieHhmNeNBKEyTQGz/kOd33GSC8g1O5LGxJgO4uNddWCsJSAK4KZ7b1v0
toxg7CH8y71HDa5onRyHCDFi14/XVSRcrai/dYHKxtBluDnTOtHhEl0mzDV9yQ4XFH1UHJcYbGto
a+NPUyt9wUWfmLeb9HIje2V5JKtasuXeppshByr5UBnqPGdVczFvlYSD5cYKvfoPZ/LNdkU/ZVHF
MyeHvL5SEiY7fqbVg9a9OjxujgJG5sYV/RnDywmeoNf6Yg+SB5Q73PAvx1z9J0Ugr16rO5GQuvKD
udMj2HBGtbotPjAkMK8X9zXHgQyClAm40a/quVdT8t5bTI7SN36mQvShDwOsR1UhjoVu8rdmNfDx
I9p6o2hA5z+DgVBOSFtmNYCgOvu7dUPABTB91A+LhWkEYg4AhqnsgOsTI4icMh2N/YIurzb62jI5
/+kC11ybkYDNSkMnjoev4FgUUp73YAa7Ox6Mc47GJrFfCzuYfDSSohS8yJmEoEfRiAU7hIA/9yOD
CUVfMZ75Ovyj1w268/6DDhAo6qNeBQHpEwxb5YhX6EuzdYq37+pua9hCkpvre0JokFcjyRdTWOxt
C74DAWhTVo6WR8NzlVUEx7ataJZNqzAYdVQp2r4GqwNnhDCSyzTOgbiSTI7YZLr0NouEggxQiqMJ
wFKz5ZgCfefFCB5cSdPMuJ1dl8Q/P4oStoQ+SXQMZ56gnN7SoxLeV9TYQshl987oKj3zJeoRSzkU
rkCVlqHJfY/9F5jIWQPoVrBAENvvd2N7vshW4wiSLntjUVdMG5e4HCMOXGNwyxXYQPeEr8J8455z
JWw0NxWiHA3tlBsTE1TXzY/VKxkl4vWbmNQqfzLyMNWw0XUWYfKxobDHBs8LbbNxbDgnUfvdAVB2
MvjloDqAwprHqw9W6Ovmk6E35HgGe1bCyHbqXNImvSsYUt9/94OtFFnP+9ktLE+4WiAhfnKIRkwz
SmfwDp3OKRAf6Tq4H8EN2vmzyCd9DdQcUDOtN0h7Fo58MJWjIApNIkcUEZMH0zm3/VppJh6xtK6r
kQqNKAEONbd1i20RXeAKI6kXPUZuuw4Pcgd768o4XwlT62eC7o7Y3I2gs4qqpmBKOVpt5sZWTEcf
57H0iYJHMceJLkHWAUGp15x3/6QcGF5lDuQwfIDi21fFtbWZLXjfqBGw2l7C8uOr5BlAOlTvAxR9
Wb6L8TPLJfVs7IqHgd3EZbgqYQ+T+YD1Cl5PvYYzp0fH8Cwpgaq7QdUFhWFyxUkAAXJ9nUgAdv4s
rfWZniXYZgXuN7k2UrMxfWXbi4buuqKeusJ/NDHfqv60Jm7oAA/VdO+4jcBnxSNdN5jjreyBNBVT
xHkHK2aOTQVv29CTCSLkJzc+FHokXi+ZJlg9Q+oKCJThtWnMDCIfx6/yuT4R0d+pBNN9YbpYY23t
nXwK2vL8rjADkzxpsBG5sGihcwB6mtgMRToAzlpSeJ/6nbWZ2bcTjIESEBeqoP8ajfvggRQ0qz16
IpQOFkSgpeUS11EH5hWzzy0mRtPlH1GiPXvLoYEPNqcbQym4Nnf8baauLP8OitOLHNAiv0uXjswf
bactfsh02W0k/0RBTy6k1v8F+K7x0rd+WfaUf2xefH+2qiwdp8c+vPCRbykFfCCpemaXA4iLW3T/
Tzko0qOIdsbiN068ZqDoRGnHGUoMLn+5+UA5PQX3tav8a8cV72DnPOw+ffP2QnHwn7aptRfI/D/B
nSzCL6JxvcmciH5fmc6EbY70J4SuGE21EQNYFproYt9WitnK70VLhiQk1EG5KQlPReADd4bOT5Bn
T4Ny/NC17TWtZ4w6FEQrQVSrThN8JJyzye1mIVJXoMe0gkIxhgAalYx0wrb25kyq1FGEZ7+nZZ2P
PM/y73/4huK2g7z5KAt+UEL80AQhGKsVipcx1uHn5QODDPY/DAPIdlXV3xca8lTGwqfLv7y750TH
gem0UJdKq6ICP2dvWUac6tBxY5HvcRec6aDutJEKT5IT9/t4VJDlWtZ6f4kbmsN6HG+XliX+KlT6
dYxjxxEfXttmaERL0ftti5wNhU2vvf0bsR61blpkPNl7H0d14NZUAlQpRFVntxi+AnjA3KlUn7zD
jXmVVXiXf27Flmwj1l1jvGhYf2ofyW/qJiAjCaHVvXHMCK9Rn3kXoxIfT6Z5lMf85leid7OiAizb
3ab/TDFu0UWdWfKzLYVAehAXM1hfKiHQuX+zaASy12QIB4fMp4b/kAO70cqUba11GlwKUh7RsY2F
i9TywvvLOfxfzorQp7aJpgrvX2GsZTrq+FPCI1FkNAiO5d4XTNM+6RdugiPsn7xDGBt6K1bb4JHB
W4eTwOMlDdtm9aJhwvi6vl5ZkOWIgQFGz2LYRdV3eu+9OPvHyI3NKaiCUcMcSJsb9nOfukd8kF6c
R3Kt+VGeppP7FIxQJRHTEEdO2pgrbjc2AfWc7vBKEeD55oCivwLR7xLXfIHNrrBynj8FzYGU6ymy
XXQVYbXHB4o+E0Oxfkh7V1ygZaYI4/nu10Ga1UubmKK4gQtqPebeJ2RDrKV5lgywZVaKV21MEUxZ
0Y/FnmjhacLi2g7z50Rmpc4JKya4rb7Qt+CHZTs/6sTMQcoFfEg+SQbIQKVWT7Ko5jFKecAudm9A
GE/vaa9duSNE/WeH0go6Hp7RSbJPJ9qTZ/BVwJfOCG1Z7Vki1n5X3zM+Mb05H0FXebgoWdxnFby4
GkIILt8B1hxl3hIIGOQVdf/uPWf0RT/nYF8XqJIPh1/rP3tFj+KC1S06gMNP0EMrwxwoxXTHNysQ
LY6CQMmalHwGPhxCANVBYpMwrIgRbpRjob34DyqcqKo8PFZYAIwXSEF2i+xVC78z16NdPMVzWchC
cgg550+bPDddvm++6m9qq7pZ+8hTMWzB+faA/8LKSwclNfeYhJG9phoHzPVEJiTFrq/5lJNiOe/I
MeSQ2tqnfxUL1K34QlGNrYofIWYfJF3k5OJFwisxKZvk+58c0jfJ1GkA6eFhLxc0dY6vjgN58BmP
gEf7r3dyY5xVQ34oLRRvrIre02+iD+3BxAcXmL+yyDSgMaFVyCNQqMqAJxwYRTZh+2RaPSyFxQOt
NTP3wFObl9s+QW6tyUjnuCLYtWc+Mhm3lwMqzsvR/yW6WZvX3tZbjovUVitn0hzLXxZEvxpCXmb4
CkZaO3rb+B/h3fc54flELiZn6Qak8JhpxQSiNYBKfEG1ZWfskKcQknufJQ1ID0feG9oSIcjx95ow
rMWdok1ApaCXD9lT/r4x51XuzIYM3tucLaHyVM/q/4eeGE6zLFsoxWURjQ+HQEafSkLjULsBArWJ
iyeXGu09a6X6y9lpQOV73vHDAWAxcXz8rfAQbxEUOxBOSxEDzF8r2qpwFvjuKMnAG9zJVwXuPBQO
nzrHzP/myxgwODUrqQ9T70uE+ZeYUA9LV3PO8BZjOzbLk1t23wuVCAFNBjI1FjTbt5rEWR20K6p0
5ECs4nJUE0p1bArzVuQbitBahvPjSxI7lvZzH4HrzBikSbRo+eLNrWimoniuCv5zJPkCnocWbY8z
m9S8+02ifhvXzcC24w/iEXm/bwlzZeLuBCET2LHgwoAHaUlq5gqbPY2eCJbOakbhd4z1oAp0GsMr
/rZesAqlK7Pet9ctmnbHJ0Piwrsa6teo+BylZg71mab/L5n7CkLWLS9HB+T6f/XNuBZ0henG0xJk
+FeuQeT26Y5FCjLwCvAzuD8yZQ66+KVelgbNUwksKuzYsVGlddbfsWmDhg1pUHvY6sNyTQJV85YW
TW7MmhI3hBJ/acSQmS0cPhkiqmVUqfZ/FsIpFSu/Ul+3AeIMzMmXfO6aH+zvnWhdMFz7lXeoV0qs
7vidhSLyezUxFE894pnk/vFQtx3FQZQceeR6163u0bjNw95d4NK63m+8yhOBy95uTMRBI/GeaVzx
OUliQjdTM60HM6IyJhM8dEmFkMO9Jz4JweOVc1R3fiWLf3uwIEBPWZXFUPny9NXnAY39mligSGWv
jN3xdGY7aJkDWONdq/pxcwpfX0LBUO5i28wHUPlczgPnebbSiyonikgfCdpe1DcPqTwLcAc/8pfL
3dE0BR+S/VQXtU8+fimG9TR1YlSN8WeKMMvbV6nqvqsYnCkB9EDCDHcHj+K/BL2neub6w+zwVs38
Bu1JL1JdatD5mOq3XC43s3CtZjTZo2xUl7v+x33lmBC7YxOrBNYPvHd1FG004/MT1gDAlX1PGIww
hYZS7MCDZeXkfWIDLOT3yG4b+jqqiWSCvrUVMvx0gOMVLJfoLegdfFjMfEVjEhs5dcz5mSwqYqLE
aJoIszLs3KfwKBiQbtNpyxE+fg+EqAxH2R/9rsCP1wZpdtagqKWSd1Z5Q/3+mQeW7kCgA3q1A1wC
H36XnfFRIslj7nzIaE52JFnCvVErURIQbHLerFDt8/FX5EzubPsQYZZlUTVeB/MbiD5cQTdfL9Bz
BZRM/A3PUETgVkIJVzvzxKAn7mirQ/v1Y9TsWqRTP2RiW3bgbCGcN2muQzSVXM4l9AiQHTlMpPF+
tFven7RVCfqYbyEK/kcsjcp/L7T4tJ5J253E7HiUU0a2BrAPoP6GjAjwEmIExOObKD+dCsuO0hiI
xemzo4XcuoyFzPgoNNNfK/6bNld0OyBjvRZ7Dx+dTfjLsYQWFBtpkBgAjD6hcVZL0hSBwJyHrJ7u
JgiexaKogfofTKZtzkSY/nqjJKrGM51fL7Bu0DmYSgvBuh1szM/l2jYqJjNpEz+A3RDJ7uymDxGB
kbHV4n8CjICe+/TljdsPJiugtKK5MvicL6iGGGQA7r95TJsvv1fvSDgzSNYwKdSOoGv1zf6roxbi
oQzso8B7T3bBcOlBCuQv2SiL9JZlwlfySzWIsPGq+ppqt4wNsUFXhvi3BnQVndnT3elRF72DWcXl
zFWl7cTXgUJAgZMyuVmR5jJpoVVe9wGklJVDztTVF7+AO+RCA4OpHzoufGnGLnmbYi2AyKtYnYoy
cQc6PQL8F4hgpYxKhI3W5LrsbB5f4HZxrtDlXDR3ArmSYSt6rcCZEkPoo07zRW+HV/2IQcBRz4Tl
EU65xMxDabau/auquN5vJPNw0C8L0lCIu3b7vjYe8ktz8kZpz1KU+BDQCQi2x1FkpB08wvsJuLKP
BP58LUgti3meYw8g/eSyE0njWYhJCgV8xstgqAqNkK4CU6eSFtldqw/a5Nw/0cNOrMnbVpVTGX/n
zFandhLN8TZlDwqx65Lb5vmQqMYuIyPCA6G2slhMD8BFvRnCGdRuGjKN/JEHjlnvzln7Qc5b8nPf
2Orx+J09IGeSAOIAgD+uc62GlL4i9qQFAYaheRP/TSorEQEUlDEIiBxrB4692Rp1KJBvc+SHCNt1
hxmLdpupVbUKjsACmLwiuQb4/NZCZxEUpLlCf5OVefudXa/U3OjiWGk2rVedCJdpH+jz2sTusC+Q
2GM2Ud+TYfkLatipiwh6ABPZA6xRc+L9+f/nOcbQAEZ8UYoBdC0WsF1QPPi0wFZdEHVW9QldTrPO
hiSCfr4dpbujJ//ElUST3uC1dfykifdZgZRyK7pws+j3RP9YQJEkRdWBytKMhldaWcq8HWAqe3ab
KtTpJwOC8QFsGBVv07YHzTKGwyZRHvu0/FUvEF9DtEQruUFYGAVR27Vb6tbeXPfdpr6tfMGLTYfA
9jQ9H1jKGdXMIA1wSTahTo6wv9VLJbv08/Fo7vBqce8Dtb0cA07dpiS+r6K7syBvgjQVuwEV76YG
rx9DX5U7b9mx54A060htgsz+P58tD+e4zMcmmb36SiM447I8a/JNF86j1ENOyWz2RMqO6pwO0iPb
i1T6Cl9xQXujY44+X1OJpwDn5D1fG1CXUCMUtlSgCjW/iBnFlhoVfU2gyWImWEwXftm3JE2eQHpk
BZVnQ3Jrw3tQiHVSkKUjfUTt8cT8XDLunfipqKUhCT/neeDJAKrb5JqJvEyuER/3jiPAYcbZ/xOh
mdOw5BCilCfVBfaAHqdDOyajcjl/dWZilPqX37MatAuppusXZgRd31m9Xi6+xfpvIv6pZM8a5cTO
Y8R2B21QhNqV0Gf9sA7sXwb2qgG0JDyyVjsKWQGAohpRkIXCzrkyHSOmwbG0WhBX/SicEuDW4IPe
iPafl4wqaaFR2xae8epo2Evc0M/SjFhvQQD3MomZHTJaD5DDJ3uZeCq0jsImd30s+XKmN5MofL32
N+4i3pNBLa2TLSokU3pEa4zmO+fZ0lfJNWYZiABzUVf70tdzXnj6+CWQKagDy2BWG2zEte8InvvM
vvCbsG5WAD4vXAnkpQeZfDyhNCrp2ATspw/2bF3JvfRxXYZ5QNMf2PdPNhneD6uP7rQnjEdR67M6
waB32dincdE7q+VStIL4HW6dq37zPKB7LpoVrC/eVBZKHyjViN5WbbTi8r4spYnXhuuuaqh9PlnV
oruVbdOJBNULXRx8cMPffh3v5W2KbQa5nabSzybnvnSD5Tfe2rxTJE7Epb3Geac96vvYzfNcHjb8
ByuL/LCk/UbbSPycuv19uaYkIRDjLh2GegexADHEV7gMO0h2IpXAZsvjDIKQbRuHbd9iUtzt/qey
250Dlj6HXC55tvUzRHrYcaXc5KQ4UezTq6l+YdK5siie0ZrtFWOUMveopVgCOFgVL2FbVVWruSIw
TAXQJFLdGbswIasXxncXzcC9X3SsIUlNR+tJbKflQy9eVdPTAEcRaH31U2ED/jDLJ4kj1NLw11Zs
KcdoUbarnIFkgxURrtsJPTeqj5k0D8fdoOIF4r4IaidxDojB0bLh42Q84IRn3PR+oIAp7YEw+MZu
Yht7ISU/wIeY8RVRPlXc00SUuRTEAo1PO5MmAFsIAYL2Fvn/cB3fIc0RrSuwTHVas+sx/aV/tLj6
VJ/SPxKkvfYPSu1WaDY/SqDctYozkoY6v778DjymAj0sGTD9b8tjIsmTagUTOQEtapoAyDtlBIEG
iekRDIU2FnSMROFbeYQPz2Gq8s3zKjXNObwamDRV12T1Ty1/2n9+ck0fjvbO/pgr39iapaprT/gJ
CmjzL8gVzMzt/+wuHWEgsDupRczNB09RQrRKDbklcRpkvCQJLkbpOz2OUMcmF3/1Fx75nIZsTcKm
aHiwkhtZXjZVicxlcSv73Vad9NbkV+V57fMyYicmnU6pvQbo+yZsyEzJpWvyGS/OISrJ0b2U/Ac/
mDhZ+IdFqk6f7B7ofIBTGBuZ4QtJSmEAm9D/jDBYZwzP5Db/jf/FiCDtSN1tJw09YQi3JAtn1TO8
NWFBjp0B7P7UCHqbMASe38TtzxrvqVamcN4wxsNXdCQOgZtrBtZfdgU+6McM3xKX0STS8IYJAZug
R+bkaGjLXHpYIt2dyTWgKFIUtq7h0Mh1OOei1LMw7Fg0Wu1ulY/UF6FbLsyH5hrz9BFfWNkjFo0B
f/t22hLsOUn2dx+OdsNtgvVmuZC/OttEV0B47R11nWfqdyUe5OQRMuD4AJelFaI0fUZ89y9mCS54
b/WrXMqr+rc6g6ClBTmfsevzClZ5OgRMabX05BoQmD3DsDjHphZ/Avl/u9BfQvnHzYthcBJEpW0p
4v5HbdXcMgAMTJ030DRvAesB3zyC4HUfPKd1E4/td2HiPQ5BgdBSwewNGsdxYgurKKuvR/XMInxq
DKN6AkNqJsZ4xg4M6uNxAdWTblZgOIy33dRtW8CDro9lRPNzjnkQK908fVXHQpsOOtgk75JldOH+
VwxZsktx+cq98j4YaKD6ESUuxqrSbjQyTn1q+8X8/YnIWYeb9uFRc4EkH6sUwdmIryteahqczBXL
yl4tFEHS3y0JYG2/KkUSBxVeeVmJEiTnZ6CIaXyucX3qHCQkeNYKJh43TQSKvyYaL6tfPP7t8uLd
uPkR9+AufpUHWJ9KuO7g1lg0GqrFqJS01MvhItjcNTlGzhZaxMA/IM1rHjC+VWkErTIDfypGXzEX
SsHKDdU8ZGw1xFT8RonVuZwYr/iTCMwBfRC2GtJy1fV4t/IOO6aWAGvpkC7gqT5+k/ipNUBe2nMw
1jVY0oT2yGLzNVU1Zlx4wSPgyz+Qr/i8cpfirwCtLV+0GeNrMoIj1++LkbblVtrEHU/w0n0IiThR
kDYLNub6a2oJgx59R5+Us85tP8Wt70+d7BNFY9Ey99RFYmwUjY69eGqUVXYGz4EEZCN3gr3JeqBA
XZGn9JLlF2+pr23OKcbmeTiNbpIw5Xky4wPKqKgLhH4KsOzchDs6EKeoqma1egHeCZG4XZuK0BoD
kS5PG8dOZ4ps/3Q4Qx8KYNW7SM3eJJM9gHBLb2SJ7Eqq/p0a6Hl7v2WgeqBc3H83bUzD/aVGDjfE
ZGMphbECTq0YIUKzF2bbQ/X5JR7fNSvpBxwg4yBRIYpLusQN24Xo4vhMxb3l7GqVsiITW6a8Fge0
Kqypnc4KYNhTXzMft3v3fjKWKTxLpgcBN8tYrT5/C4oB+vs3t+cWTjiD9sx+4NvV1uBH0utoUiBM
WmpnBnvqjLAr0SQh2jCIQud6c+EjDkv4/IQ9igvfMgRxXM8tutny51qS5APwwY0Y3acVO6BQe8fw
02UxKPKVda8l6fBM/w/puui21uBGZ4CaR/+WMWOWMgc2G2Xx+vzDCX3/ybcvuwZUGMfSNt0yktkV
t2CfGpe6zGUE2x/XlHsAQbzobYwygoRkcRT1kwNzwmH/8jjWbbr0owpQq8aJqB8mFmSQ4Bxnv87r
mY+bF+gDwRAvGspIVp6nNZfqSDP2jXo8zXE9Ac/i5ZqGqQQ6CD/6LdzBCQv0y3NhcPNl0/x9gPBr
OwthPqLBivJGHU0Rl9rBmH6EgTiLY2go+W61BpdhWWE2CXahVJO4eRN7tmkIxngczbdLi++api8o
lZj7LBFFvM3jpMMzjBC8wVq2y2rzeYG9rFBcDvTIE8SoZZTaNJzfTy68x5QQm8egw9goM4mtSloO
+YgGwkpxIJJt9XFUuNqPasoX1tX/qzT++ILDik+ZC0x8MZLQ0FqKA9qpLC+g0yB9YmMwpJOMUldz
J3miJwjhdpwAHr6qrczUXL/njgM8duOTFmOxCjb2RjnvTwBmjtzjB8Hs1k3barvL6HMQnzeFuFAE
LT1nIFJxW+73qax+zeUAUYUC/fOIMhHcyeQfoNUqmE7LOOlQiy1oVDPFEvc7IjJ5zlnsEnzuLl0J
uIORbtHk/H+Yqd3x07QQ3MU/DhC9B0DpptmVBXTWx+bPYiNEnB4rzDlMdiCPFObF3XHpof+dba0V
Bp43QApg5M08cXqFVUuUXLhf4Sv9dCqjf+YDeg+oNJNf04YCw3KYIbQImPrKHZO81TlgK29TdASw
8EXjzv56JcRIXbLeSeGbCZSfNCU/7/EQ8qfJsnVXcOBUPBDPuQe9DH81sBSA1IKBhma5N6kq9zHP
P/w0UO7jxszymy9pSNV6JBemIrhI+NGLMtyjXKInhdOyttjs67R4QGW8gKEWqRJlmkaUju9D264q
ElBr4VqNkX4OYUFBLjNIouDJaw3JDzjXtl1VGakgREWWwJDyM24lDseLN7/LMX26ft2v0uD8BZ1B
JM9Q8nSC9ZGMgR0wdiQ06kvTfi+maEiianFwTnwXWpBXOlycIPdl35VJiLXk7fu3rjJ09tqGC+yR
6aQBOGat8AnnTKhAnBUqBNbAPzaFWQEkrpyci7GDbMyF7NXOkJNkfhWKNjiBfH+mXLdhfv8WQxCP
7TVslyBuz+N4OqwbTUbRN94yi1pMrLjLQCA+VuRR8ifaaXR/LDh4pv46miG0mVAdeq1BaBCRrY2M
z1w8DIKofMPHmYCYlwUR/CdQvee3bIx7TYwkQK5JDNlWG/5N19948RYf+wIHr/p5GKn66xPfyMSe
L0N7zTcjV9iDbyKp+rAKFEfSrIVeteOdZQwbRWSNmepWkWR4bsY8piJGce8RZAAdQjtiMFsuClvp
sioud/KTZQXY0vMm4vmLVjA3zY1v91O1/tu/CvF6CV/HTYtd/4cNRUUkanLAoGZ2Zg7FP9sa/9+L
W7htllU9a2OO+FuEgDrwt7VVLy3QVmXfQnNfwfE9iQTcjekxG/u8zDQfLX6uI1L6wiFrXF1vEgxZ
OrgJhlK1Wa6/dF2lTljd3VdrQwRDRMIDiB3KjFVY9E9A1tGNkWEPC+mPw5p+YI/SQnGiDgPhKZVf
Ua0RqCVpYoD3CYSJJfh64TP8+QezyzCs4xCjd9dpo0iCnufXtBvb3qnTRyu4aHcVdx2BnQ5NiB40
lt9fph/rFmzLhNr4pfkNQ5MOPsl3xHsLzm8apy544cRBv2jF+xbLFJXkHoci6lCkaq63K6EXvJCh
gfkmEUsgib74bsJfSTgPgvHoDr5aQJH38S8R0xdsXVNVUpjQNKL/QxaEJieaSpK/c/r3XpBs9yIi
uYObrs2D7XZGmSZF746ynKY6lZX5hAsYn8TbVyfZF/4d+kTD4L55gMxs0bZvtWfqwMOQojSuPM+C
wQJ/WNg5mPiukWnZJLCUdbHEN+HhJsiof0UjvrjS05uaHtAgcJaCIqVXPKhoQXSZBQQaQbenQoKx
wh5TZmnSU0mCtFBSEhMiqLyee5l8KmapKN1F12rxA1TPTWfcxBUXkpWBn90akY6klJCTUfO50hcc
n2L0G/BJgBqfNEt4teEkrgmqNNTL2csghHu/zuOXcl6O63AkXrYLXVWvWaa+azp2xX3VUoheNDhK
h4HZV3oJJNipI1ah1xJAUBMYlELFi2upXoNZBqBWwi4h15ngC2NMtxVxw/HNO0AP4DlzTI4ef1Kp
6qwffjNYvstGBV3Asbf+IRfKS+A5MsKpllKzjPZex3MEP7KHicT/4yu7DFww0YJfeO0hjWkaihRO
HTTikafsF++q5Cbz3bVCulrkkwqXiOVxqehv6UyCRI0VueaHwOT8TZ7rKJi3VqVG4wOqPLoCbY5W
Ikf+G6q5ElFBxTmsfHXTV49/E9CcnrduxHgjbX4ZfqRizdYLbN6Y+U7OnI24QbjAQ8RMDvPmN0ce
byyQIfDZhOQiEFdwKlLJyhLeogHfosLQsVzS5ODxJQzOLEJgCXFN9wd6F6FIaNFbtbC3+hFd9nE8
eBdI/n8n3dWpzzIx4rBLs8MrY6Ki/Q9NqJRblktmkaBhhiS8G5gQnXo4wrs0JMo/9rpa7pbR3B4/
otDaZBPpizBfwtZifinzNF46xUd7u+Tdr9kk+u7SCFDy1Zb07lu1uFzL1aeuS+jbl6ETl9e/y7Qj
JiZP6wx/U4NGSzXLvLlbcP+97WM6R5B5qBw0qpnsAd1BXLGiqCNl9xx8tsSizY98yEacC1sD+GzA
wr39WY1D7LWkORr3t379yNAbE3Q8uSKeEVS7x3OVblGRa5MoYIM/jGVjr/wFucisbBU0KE72Qaii
sZUoilk1YYSaTwo7ii5mISPUH7EiKu5uNHqvXEcpQcPuFiZgcHkIGlyS3UY9UT1yaXM04qyi1P1k
Sj9p4S05O0fL1422S5WopNs6zI8rOKrM8KpT1JQgrudP1m/0yHTh4iFM6hDlwhyGZOh2rhkjV5qs
PKmyFvCnzVjngOHhUBAac+uiub/JQM+thzY/UQvlOFPNVwpUbThzS0f+442BdApVJTRjE1akk4SS
/jciqld/UEuhfRADiSZkW7zgfI/MxN7X+69lnLrsh0EG3djnT3Lb2xwO9WpEv02Gu+ZRxMRx1MAI
rcsVjRxdjcqUH4ASGumGGihe46KRNsFDVM7lyDmzi7ZuKNs8HDIzjPckDYDrL236HB5VzvxaGhMx
vmp2CQxvmiiqNsHC1A/t1mrfgK4u/pL9zNtodPDfyBs2l2eQ8Jtdx68YTRwmxW3oh91ZFaQCu6nh
SEz1xEJnYnHdQ5t5xMy9SVuN52zLi5qEOuPEfAPrnjrMmiAS2fGeyUnVXYY4B1E5eVsb9UX0RZBo
lRwMdaP+bvbWfvzJkXgvHl7RH781W4Ro0kbFZew/rXMKcjNj5QrxNMVjmkRQ9s/ATXbz7/R0Rboj
2yUEn3gLLG1Big+ZNmyojG4J2LMA9SLQDLjV+dWpMWjTsinDJ/z1UyGkHIeVHcO0MWOWv/BHipmI
Kb9MxCe7jDHA+9ywkd7n45BUbl3mTgHED8scC/TIegvF/UDFKNB4aJtE7/vu65p8xBRlEQsH3NUo
rJoyZOnidUc+mw2aHhIOdyNXXlpYAzyjOhIz5aSxYN0GiDgznLwN7iOc02d8kEjvW6f+Es5a2Loe
1fXan4G+AKPd0of8TZjL6wDEXb/2WrFqt5uy3njmIuo9AoYmWBNUFx5PiSWSGVGpqzXcu/k4SXsA
h3ihXj70S7RW59n3YxAbZjPU0oBp1g/oCUQ8yfv+oW0j0MFrLorFnqf/hyNQA+QprLfPxVlgDDVV
TH5KUyskBtI4A5999iHNUNETGqXuQGH5Z4sNXxdD966Ty0zu/Cj0YLhcXI2Jrs935Zq4NwXF1OKm
FARV1GG9fPtnDf0yjgzYZm3x5lUNFJHaroPCYWyYoqUe4J8SZIyBKJNe0b/G07Sxzx6v4DOyvO+F
Hxuj6NSmKeSdwKpNcTP2YGDmNC/tulOuIAuyjfxg5Sm4Xp6pWCc5BhBG1B8kHo9Wq2PBNqjFwGDy
9JwyoV8m2Do98fGl5FhXDZJSuqpEQTYC/A8i+TrvtXoGl5ruMuL9/dDVAgO9X6wp2akQvEpyqZrG
gqHlht/wQVNRTZLzAGh6bpFKyu7toqt8twP6BEixKkUsX2glZYVcKqqo3ayE/vJxXkiuVVBvS/fe
8fXy1FH2BxwmMmqkqBD915yY9SGAXzoOS2xOHNOgmBCn09c3yY4MCAGP6E4y9M52rhq2EjMMw92B
irL8t0lpLUdKiM6kcUd+s+1vbeknaFh2LK4GZkos1jluXJ+ytgi9yJol4XfR19KjEZqQf2mkT9hC
g8UGdLLTE+yPhX7YGmJPQ09Oatgvb1irn0PfVh20FO6kPni6f6T/akObmDdnHNh43nKXpt8w/GOF
HeiPwk0JZHsXPz4hpEORUvcX4PnbZmAtF1LXWf+A/gu3UwuUDZjc/WUUifioYW2ZaTCNtf/joEx8
809HP6iCxpZYlHYXRYHIAmvnz9Pw9qXC2k6d6q9qaePXFzid6TWF2IZQt7jagjzMNflhURqkKElo
/ac/1hrNBYeMFs5ToDPF6nt/cVskjPhds90+bEE2Ua2ZyFO7THiM2nmkKoIdxBinq6t0IqqI1/1x
5ZYvZHc3NyXW738mb8vVfix9baPtqblvjNPImpRbfEmA/L1Lt4xhT2nPg40zfB+JTogRz4OawnBp
oIeT6v26SnPRcKdbCyL/P3Cfy9EYlE34/pmwMSmbkPubDZ+kuBRs+fl1O5n+35cT8yBZoptLGfp7
Je+y87CWguoG1tRQGirW8w1CPGsb0C7UOcPCZquoNsA5tJY7Oz46YPKcGPew+MTD78zLT3kMoaFs
XPg+9QPR9CZBfGh9A5iZhmYzRh21LQCUdlBq93Ypf929Z1XoBuOWtRwoeBEP8g2N6Mn9quVxbAbw
qS+nj3SxrBc8lo+nKy6Tkx2imjKjGfgiNRDmps1L9LogMxZ817xSK/phvlm176X458jv2U+Na4WS
KZNdw71LyZm2mCXM8d7FbHhM15ryKc3TzCm10ap/TH9D1Z8SR0mBfdPRwZzpaNZWvcTRGjFMrLTT
LpwIZZF2IKSRe+t24YVQUckkQRo55DtsvvuSjsoKCtTXbEz+2QBiJmrAYrev6Ty0JJXCkJAn3/bG
Rrd7tR4T3NIqGOaSb+i5DnNrxdRKG4/k2TC7Ve1SQF3+D/wMxs/Oph0A/IJ9DbcxOeaZwe7XtOjD
3XURTbqP1o+1h0kMw98IGA5tVdk5xidCjdPmIMMi1Hy8tg60ZXmmZYS+/+DWPy9JoUUaOj3VNExl
klrnoaUZJY7+JP98XFmzkrAzrsfjN6hC8/3GVdOywrWJszB0TMRckj2DiDYe7wcDR5mHnbC+pY5+
g4X8kxLN7/xBWgZdFce9kG9f1XFiUIMkMdfEWEzg0vsL6naN+0dEGnXTxYRJrm+LM70iNXbQ1ryH
vrOdOhSm7svWWSnOPGOzQq7pTwN9ry/W9C3872APRaSUVqEvVlgziq2pPdgsCANdGncKJQnw5Liy
QMTM4wjADAr20IL3qrNpj87p4d5SotbqF1tzLmuAwzhJv9Lfe/Yj349BJAeWLBS7dstzKCORAs0/
UjGwiXRVjtnYlW4wD3Wg/obnyqwj7wEoGvbhN6qcHul3WQpENXPrm0Fnux5iBE8Enf0SCn84ySbE
zQ6xbjHtlJ422tI8ZhRQT1q6v9baXYyY0+9fGTs4FDJghzk/nXS1qABv9lzYaAFnajcsQiiHX/xT
DPIyqQ4q6Fr0blwxgS6iRNwMeLl/FmzGBZpAoDN+L0zhK5WmXrnZdAkkaHxAR2Xs0g9wrOGhijWP
sK3JR2DClPQs9bPurc0EqG/V3Kc3XLRFw3HwktUdeCN1OnPA5yv5B/GcdRIiyCUeSh9N1L2fD1YY
/wBj4+lcyid1B5gXZkVMlyISJkEe/AisJlpEVOQbqOmvy6youDCPYk3s/3L9GwaU6TvrCJYzCRAC
d6oqcBU0/bM396ELiA+7QN7F52NWd2OfiRJwj5a7O/nm+QZald0IcCxwdh055uPzwzg+AN8qlUGD
zJ4QoRbKU4fsN7PXGkxPjM85/NCAUpLTXvrml0hP8B1J2WVctkuW9f1eloV800MpT6ydrIxk4EKw
JpnZqMpUkjjccRVqE7KAAIzQ0Y0a838o3FU3ccnb9wEMvsxmwFxHre5DFFy0b/DFmecSnQ/3EyMK
DCnuLmT6iGEH0esWmJrR4bqwKkizw7f1XV7u93to/eIhsdRibx18qXKmnsd+ue+33AcQp7hcbOI4
NVihUDkZp5N1NwFhv8EEHx8StcKHS+PonAKDYR+cPumndwttHmvZaEsQI9e5Vvcg7NVVnepjvC4d
PHAv7O+9YjzgeNzxNnox01nRVmKtfcIOsQ145Co9K/gndibfCTY40JJjoxNoJtV+DzgXZTljH24K
5vYl9o9YV0ac6Su67nwfWtuEZ7O5a8PWN7B0zercTmKbm8lNupcDCHxOvNhp23xl6JNfRgPL9P9R
VN8eeQ6YomCeuPw+cpixiOIppc3iNrfj9cSeWSAaIdxB9QPEbZ3gaA8/VTrPGLbVkWk6bJYcgGwL
lflVNA1fw9Rxltn7xvRU0drb3zMingUB8sYXspu1QAT44KuNUEELuxoBxBa5HLoutEARg+JEahRW
oZ9+Gd/DkPyk//WRdWY971+6rYpfND+RVi/ZOK7AwBgYdutyO1uJMVEJT5GKMElcnN+njfr6Pq8o
FKcgX1xJBvBpS4kKfZJuGxS22jviL15ZIqYL/Nc3TDc8xMAvxK2uE+0MSXHhIW0hdMHCKXhUgmqv
wjjxrcpP/3kP6GidNRw0PneBo5NJiIZipM/NZHgCjaIbH/xomlfgDTCX2c3HNgUzoJzbNzyJQH0W
N8//EcHly/1Wb4JV7vX1O57iNxdAKEL7K0/RbDbGycV71vk8MAZ2I+A++mGLJL+WPRVEyYi8OiuF
FGnIPZZuEo/P43jPIdyfJSItGgEJPkxmFTOiDt00Eo2dp/nXntzMUzqWvv2uBN/nL+zx4loTjaer
ArzalCzAZiqlqAC+FmgTZi7XQagKWBzqxf1PwewwhhWP7g3Fs5/6ReeqK4YS5ShWftnnA4rQ3NNU
3CvuHWgb0jHbsOCt9lpqi33qDRR9c5/Kstm+I2OEVLxVXUnJsl//NjFQCDL8+fgItbsV7R2DZtGa
FCifG2+3iUD9ee6uy37qTPjElcjwm9iE5VqIMHz+v7gsTbvVtEZx30SMCvaHMpBJWQlO9Ksca0c7
MbWnEUmhgf+PNEwrp/SRlJcvplHURzzVUd6gUhha54ov+cpTxyh7r2yEEouitlcqXqRqnpU4hPYu
7FESu8BhwzU4peHs3yJG1VeNYMCMdFw9fgANRqByYKGSjC8HL7bh7VPfv4pOvbpxMTriy7e8Zeep
pDRcv+aYz3ooFSQVib+iQxhezZpNNBke/56dwh+Y8QTxM8JuVw6YEUhmpMh2BO1us5Sk8+FSMx1R
4GlOc4f5LwtRk8LGTyyYgu43EO8yjflL05QY4Sk1aZBfY+vZWsGPSFLMkoKGmLd5dUCcBIbpNnmJ
lTZItFABysjb+6aX7WlUs1wFL4v/j5x5dAF0xCswzYmU4mM26afrmIKJPMFMAPylwoy/6bQU5Q29
tFmI4tt3qEpwVAQiPdw3fbTzxeEnS/TCz1B2DGPCYbGG9tIe36XSMpByzEbG8h/KKHxGvpcwV83Q
8q0xUBP/y2UkpDex5eSsWux4Go/g/he+V2oc2Vy1hRFqeIOmADZb5q7vCPDt0dhPbpafwpWwSQzC
q7agbOydEwZK+HuvB+M3+9tBm+wJRpUH7XDQtSEPKmgpBmTYCdNuPxeIkjAknhrEF9RC6bWfoxwI
c8xfYFkwqxCHmghQxcXU9ZviBMRgpKBLw3UOrL94nCkcw48pg4uco6O/NEmYlChAXy4zCxB4L6y4
TXMv8GBUypNjv0b2OnJU29zxJPNU25rsDadegtF9J1zsVxx2XX/9Tn29ZcPqi8YfjpIZlFb3M6mT
zduHWj5BNuNlXSi/E8Z9BmE3WedTVTDF0n7EzTZK0XKHACyvJwQDPOKDDKvLXRW4uB9l6dU5TVxy
w8UZdrkInFtJJAyPrPcnIn9VA83k1WKBlzNohTYThnA1ovcaiuGcAhAhMvtu3umgZ2WS2qixFqPu
9rnAA1G+qaO9x0oNBho4KIzS6hMHItpeIja/ObYQ470zYAszDpcT8gstjMPOSiAQ/MvKu1+jQLV5
MY6vUo1Bv3tEupATcJO+azpKVYGnZQ8rp66jp9ZlzTGNdxenXjtvvMOuYIZiOL8/rOqPvJ965npq
QnF/gnY/txWkI3VlqItpDWX81zpUB9jO7p1RqP6Hul1b2LOzS2a0Z8yDr9x/DuY1sj2mT5iavQQ1
VkYWYXgnOFIKGzfxb2x3zHDURnZqWFJfxSMv4o8RfqL+J5U6Lj/vvaoNL+UMcVquB1Sc0Mdog7vv
hd9VaY8YM8OG5t8M2dAorVXybJ4IObY5fJ+Eju6ANUuZNQb5VHJoB+qcJ9YE91yOpNcnn2ZjBbPM
SPoC9nKx0Zg5vD8f9ztFM3YZ4T/F7GhJIRbuQFWYamoVdp0AQZTQABTSa0ri2MsFYY2ImJeR07fC
94KAQXqtvA5oP1tD6TdE/UUfl5a79WsfWEFQu3WgBCe4cOnmFOOHp97NkDYFBnmPA9/Y6LWTQS30
EqPO+o5XXU7GldwrtytSQ1Qfg/MMdoDPSPXUq2AaANMCnlw975VvsP2TPKDmzdYONRe8/doKUVj5
5//N4BYuQLKgmCgwoGqUQJxYb0+ZsrqhxJh5lEjB9C/oMfMxrhRUcin9LT5YHBG7JAgWArcG/y6T
s34bGEH3J2u80cWx1wRUWUa9VJTAd8JHCJcfEOB01rsCTw5TELNND/p3pEZIt8GCSE2PkLCiDX2C
spDvik+rokkouWpILU9BTgr5WwU2/mbPilzV8wRbKC5p91RHiNv18RsLA09cXKBh8TigPDBO67g4
m6ymbq9F2VXh1LHa9bPmA21Dk+vP935vWzjAKce+22EIDGYfjncPxv0G9eKs1kps/F5PmMm9VwSA
E5n8Nz3dhZ1RLHCqfEwl6geA2PDSjUr6vhf04JWKoXDnnZDXw4dAGKcG+DIPV/RZYwzF6Rlvi0ST
2iRo6Y5f7Qz3wGnHhAyLl0QPOVJ2a+oiVNh7dfo271eX9sPkpb5CfXLMQGT3/oXz1h2AyWt7w429
jOv3+869O4Ez03S4jWBMhd4PKhe7ZpP8mRAiuw2UwOJ06CL3LorxGDbrO/J4z3DWArshm+sdywSc
IlJ5YZ2P04VI/H47kAlrlnpezfNtid2nVCXk6jmdQNht9R+h/b+8RMREr2oI2aLbvwCrsXqeT9z3
YUUcY7mXMQpWKLzoKQ6I7A2VVDqkIKEdaCIcmV2hD1tgh7ReDEaL/1ULeWi7e9c9bR4gYhPAGlju
ynDZkNplulD/a4fxGrxJsSmE5dMHechDl7f4qciWLLX2LLTv/caRpL1x+SBb6kGOjOEMgwSr8PXT
UDUeAVrZZ0o41YmqaMkE3sXDgt8fBIRmuJA+itCc1iLQyS25toimDv9V1/y6pqoa6tkwoPfgjPia
wJBE/YBVfqhfu1QzQwzgN7pxB1j0Nnj74GA1RR+xnLaH1RXWpN4ys/X7Y9McapPOAkMA+iz2NiuI
zsmzJBH5PsizgKW41tGUr4PO+GYWZbYis6SSgmQRJhRQKsHtOZGrQ6+7S60goL/E207Yq4gJ64rG
XJ+2FVdWYBuH2AkBnzYYEqQyogRNR315rE3QPLu2G3nicV9DDQSSLmsErcogwRGMXFzqSXuVcsJH
2XKy2TuTBLeVGs0HJZBg17uToST+r5aAt7KaEVZz5GGHFb3oWTy/TLO0b/h+ZC/XxgkXGN0FGGWN
MaRHyTtMEpLs2U3GsErWttR7wM3du8J6MEqM0e0CZq/ebKPvtHXypPk1JyYS/fmFtSraSzrc8GZ7
VO8lCAom1yd1K0PT+krAc+ykcnksIkPZPB2CNa0MJ6CTYIcpkfmihir6jCobitUz1TbM7a6zykCw
0dt1iB7KZplzJqN4WLkNQS9ltwuMYg3oOKhPhjavryIdZP6kBdEF9N5peoP31IM20IB4zaU0q2Yv
GKj1iiM37mLAvBOlHPXuvSQMFVSsm/JroHXqg8eSPKtnJUkGO/BoEyWrMSoVz51pB4uN46MatcKC
kRN4/EQB7LQZH0+Bu1rpzwLvPnwZj/6TdAE6hn5gT1MIYwwUfjGsGE+ub+4h/BPWhanou6yWEzqV
hFyxivDKxeo+Kd4/ViP2DtXeXclMaIX52HcQ8DhFaCq2s8ACyBqSl24CpxXs/AdMM/dZUD+5RG5y
ztsQlzTc+hLc3r73L+gq3+2SGiFqhBsTmRKngJCjAMxE6J02xdCmE4BO55LOsLNQZxqDXKEn8Owp
v7QAXDUw09MsyBTTkj44hjyLjboMV5R5t7lmfFqawMC1tMW/Mj59CBi+axu3eot6Ffh3VySzPHt0
Yc+dB1Oe+2UkhCHGckooQA1gm92qb+L5z68wHx4A7oylFmVYEUlFDDeKCJOITXYPEDgv0spFAXRD
ofCDm32RD8aiH5+bIEnDghLeBSs7tPq6iF+BhSU9ThRa7iXf8Lbrj4TbHixTaXhWlGlud99BLNak
5ieq9RFtLm/Wbv1o5bOfCpSn9iRbc5e6LjRjLQbxMuRqnWVvNwtvEpjreZE2g2FrJArZq1MdNMLd
8JYZh6vSdfYRwbcsgrpFaItsTmDFNRvfF4qV7v9JzbIc9WhNSFZys3LguV93lJwmzaFJXWS4iDM/
ve1mq8ku1Va0oyoOoMjMmEw8aZDIHAFXE7JdZfPlqqaKQ8xxJQbXalqCFImQNWrCv95YJ0KdVPyH
tOaqomBBEY5nHrXHy+UUpIjyLrqRmi5vr4LBR7X88BdbdNIDvfrKVFxI0QKglT3PEv864Xn5zEN6
tFVBV7OkV8r1T8HucZQJuAgq5ENY0qLi6FKFL+U2e2Ua2cjDJ+dyfiNCcR1IOQQSOcz9skVFHxqX
BTAn3NvUHEmVO3Rm+vYmtrXBksIni+zZKIrwu1JdW+D1Mm4pQRurX1nFcKT75NB3UjXlgXkVc5jk
xB68PO5aUrhp240XW5QNnDm+j9EGJCEFXRaIT0Lz/zThQ6TqxqKJZyLtNQriaDbCExbKYcxWcsGm
PGWCM+8HNUiJj3Lu5II0mTUZb1qVPMFQPBIKE5DlZLt1tAD9VisB8fMhl6B5oWeRmFp4RxgF3AFy
GPIaamANXNb03blJkUXIpw92G3mO+hevm1KresTiEGCB+nVXFwQKGf0QnSMt+D7RvbEGp5PgOO3z
0IJ4XDNVdkmmhrS/TnArXodx1XTDID4GHdVqTFCovy4oT4N1ra3S7KtKqMTD37mIyZFjG69CCUXt
DJ4cyQ0zS4UsBh97chdVJ/2orkEuZB7YabAHT1H4xsdOczmy+5r3slOIPQ56631hwqVQKOD672jp
DEoZeu1U4+V4aRuRHjQyRRsGogPeLCISWW+L1jS0fHLHZ3xa2xrdVMElrHWsM1LZ0CVMAInNmFd6
3t34BUY/wO8GUwbdNBeGHL20GtqetEVvFIM3rPTpKEjV3okaM+4gVCdFgK3A6s0SkbQakU/rDqv8
HrgGm2Ln2UX5gHXTroblsnMQR8zW2TPVizoMtoySfSNX8wJrQ9B3mTUWpsgvxwwiGoAXDsk6MCax
EkIqpHyDp1r5U9JOCS5xW1qhAFf6CLvwd64tHan/f/hgM0zDCtHEdRfB3UrJHYQh0OmmdfsvEYyC
3louT/4t41V3Ej/Eng04vMq2SSwzR8ve3z+7cyh2DCI9J4W0nOpFLIdIIJnPqDDy/1nn9+9TNcjX
V8ozHyu9I2FJ80T69wvWeBcF6SPrwgMvXiATEBKVdp6OZSpMWcJeawWQ4Lqm/VqCILJqg6j7jnml
R1zYQN7IZIPFbSGCclNB63YNl5oSpaeepMx95gg0rb31dZOkUqVup6+5nKp0uG1knV0CDGQd2gU4
DiGBXG3Ijy0CwazlvH9Fn6UZb/QXk4r76KWtGKVrVI+YArsp+0MPXCxL/tlhjVgcUzMG2REnQvrM
gqk5yl+1ggKyfuaA9Q7aLkHArfL2l/LPGU0s7iYassvzPMP9bPRIcYE6YUX8hAD68Dlz/NoPS+Qr
tGFuPPPL7JFUtcLSSdWHoeypemNtaI5D3+ihTuZcw9fMXua85Ge0bQjhsC7bFYa0VZ2LOFPgPtzK
dm2Dx62WYvcgnLDD5aBhb+oNWT/GiwpOJzeZp9pIKFTwfzyltVt9tSMhKSczmDFwTgZckgqWeD9d
FdQvZVcKfmM4zj0xbENYcSmuUdMQty5vs1pdAYQ0c/6iuZTyXTG2tEm05XHwsHkC0YhgYlv7D+A6
daCBjYnEAeuO3CIIiUnIgrOgtUIVyqLxL+cjqBrXLHKfLhpTWTWgb+NoFwn/r2i9KRWm9yypcxTl
Y2KM5uRlF6UgHcWhRnY9DRLS2OoFO+TaJS3KnXrlaNYLHiysN14KJ7AF2rgUR/DVxzvxTxPbvIux
FxiyroloKry/vdRH7m15YSVJu6ObBri7H3bonnT8R/vncsaFyqSrDR5vSEXzXSb3lEs8De8QlRQT
nACyIwImcAERYsNees8T40Dhs+ip0HINXREriupXJ2fVnDfU67w6LBetl92djIcNgxTJ8Qu/Zybr
ol30hBHq+/3M32o0z+37AWu19v0Eei27rLYnYeXtpfzQHBa7lrgv1w7T8lc2c81PoNLUWK/8i5l1
WbcSCldV6GC5GdRS6jjoHq8zd3rFzb939bEc0VXYZvAJFPrFUuMwNP8XNeLLHBirMAyM2Df1lpYe
A/UZZgx+1UuWy5B+ZlOKdZPJncZLJd3toq1Gh1XsZ7QoodxLuOfbeHTJbO3QsJPzVBy8gjKYREJl
JN+LkMEwxEBT2lT+X/twFFADOUrQk91mW7pqeAlWFIhgld77sldO4vuSBjsb1BFh4eIbwimQuzvf
B1K6wq0kjOazToF/xFKqapBxbH3ZGsJTd424Z+8af1nBI24er9VOE+GgrG45upiYUe2v+KhINf7Y
1WALAdLzMeIbZxX1HmlRgVWu4SXcN1zNJpHkxDqCohcMu6hBJO20km2bN74xaU70erGbIHy47X/N
u/lL0AT39dEifbx1J4eeaakS/+NZn1paFsxC6BKMZuHrw1WMk21iJ+6Wx/ULNDWfZXi3lTLo6kbg
OswBS4jFlCUyVkYFJnBpSP2oCxCljztRJ9QO0JcRAw+XXN4fg/RuuiN5aJcE0RoiiRbpQ4X6Klkn
CupSBMbITCyo342vm3MhMGG5Jph4mS+0AYI19IuNVf3vhvnAKFZXNtAjlVpTLOvcSSh4Gf1hoONE
ALBu/LXpSSf8+6LeHcKIU8w86WmxjgoJaFSNxN73HLPQBl60VwrY4bQ+gv02/IicUJqCzWIu30FR
+MZ6fcrxW74MlMHmKX1TvMHZyCdK2fYPn9nMTOEUHMzmRH+w8lyAeC85ydWf1fFy2AF2uVrzJhaR
YgKNHqu+clJVEK8HaflWni+KSrhdQoiLuJJYCgazlvFoJLOtRKnXLv2ATm852drtndjc3idCqFDp
UxA4shlWgrYtTp06kenDSPnOo7iTaNgS+9VaB4sx/jeozy+6t8uY2SBaJEkrIs+XxwvNbNr9zUi8
jjQTDvBwMyCsBSdV8+xxYwOE+Y/JW1WSzdyO5bUvNwJSLQ+leDW7fIM1GcmPXdCEqsVPxI5DNLGN
a/Qv3h35eSK+ivHr/njOeSUnUgQ0CRvL7KCR/PYwKjOQddHOIIDVnXCajJ4p3Lhxp494HsIQKxeS
EdlPu6u344z6R9xS3at03eGNYwQQfkt6ykt0kn47TPUYrqq5Gq9lwigJXZXUSRDgEZrK1xnLq2Iw
BOBmmWmP2zoPaIoD3wuHlrML0rO+thN430V9OzsWxZvXzzFhmoTW5+8hTDMxOVmg+5GW39dXIUZL
fcttwz+ckp/GX1U7k6fO/hs1C/InIAyIG5+Y4FmBhD7P4chqUp24OFF78SmiscHWvn6GssBHGPss
RNCkeen5DeFMW/lGVhKKLtHLf76n79Bf4ITqwPMgsR3ZDm1fkwSHAbX4yr8uPUh77QMQs/WSjWhn
04X4KD4L/115/sUSXXtvAx3bCtK+PKDrNUqhVcAL9afgGfIz3rTY2MvQR4A8aYDlntcd/r6XtgPt
FBhcI+W0nZBpRAb73+l5GXbuWR4fYd+61YrGPh/KOFsKepSqJ2qy6n8pgH4Bg0018YOnH3kPleN7
Wi7Yg5gcSoDE4BBdk9rC0AbjFVK8GO8+LQMHQANpo18M1BufP0WpxXj4keWq6YjGAcToFoB6dZE5
0ZuLl3hEwCDnnydIVBF0fEtKSduzNx3PnJSyhQpxcoppQFLNHPHuM84/LxaKS+H5NHOpKFsCZHGH
fkklKCwoN5wHA/XA7Y5+nJdau0mRS9yn52Xz+ATcMqnFyGG0GZ8yOT3rvaGL4JHYunNhjVKcdu3o
T3CV104wmtAN8kG4ZhPrFCZe+wK1mNfrJT//oqTZPLZa24f9VEMEyQ7KtDdFqSBFdfaZHlTNU2og
sPnHZAOM+LV7mLggaWheyMOBP50mTZ5LtCQT6K71vW/1GPVRlSLUR0Ci9CcYJ4ed1yj1mZiV72t9
uedeos+d5qrbPeDLmLlZBjMiM6HjvtOGNEHm+6SdKH/cUnKtt+LEgrGhf8DTjvky/IRbQLrP87Af
dpYRvlvMh6U1+WqYQHueRcPiE+Gv5uliBbXRYwCwut1+hWZlB/Gc4Haj6rziEhi5NhVTOjkxCt+J
aHVE02589nW7PxJv63dqcPHzad5jBqG85hjg6lkis9KsVcT/1Rr6AdqoKkH2hK7ihgIAtHFqWxaB
4otvF6dAF+JJ3auQwlvImx/vhZYfvWi/ITGjvbFKwLzYRoPJSKrrTN9wgOsrMT07hv2pbATfqTAQ
CqXQH0jDhykoJdZ3uiOlifzjo6S81zOC0gxSSbXXxdaseou/e9/p1e8r3FA86pn5h7s9j9LIeqh6
FKjkxCezW99hJP5pGT4+ExYTr+ihQzvoCUOzeXBN+7k7a1U9Nn/aVekS17MGDRTP7aCG2rnL2d6o
0xFvKCTw1JjonM9tuCCLNG3jFpDdbUaWM8Xl/xTM39N0A/ke1E8YvYP2HTp9Q44QvhXH7AS2T8yh
xBzCCe1VZuxpq6RL6fWw/jdZgCxVZst6TH1t6LvEMqH8XzDK2UZ1nfnCjfmMLIsHk74rf1FhOZaW
GkiNvgJ+aHydDmRqy8FnA5B0WlchpSO12R45znfj5ouU1arVSpAGDKTjMaZ2k9YlGXleRWr3ySmv
QOR+S1yT/BKtKz/njTggbSxBrKFWhWENRCnDrgJTtA7V/+Woy3xTQTGDPqcKrM1g1hvvbVO7WOw0
x8XjYrTbioHlwwPYW69rzVj6qHAxaQHIjhVzI01hdVcjLkEkaV8zOqIF90rTc8uPeIzJIQSFsTh3
NoPQGSQauS6LoTAQY661NzydI8XVI4lFfhOUddyObJZLQl63gI7wbuOePwXRGNRD7mqKe0HWHTh+
K785yykLn2J8/ndljXKEaSLdj1gBKzcqzNw2HOSDmcyMEKBRMjBDKhlynnZiQnUn2QXtwr4UONVt
M+3/tG17fv65FVHaYindNgNnEavgbE5AVYtW/Jj07JG4qYg22FdDnylcOVV8oOvuhJg07zHGbJTx
Ynnxv0IyuTNkqxR+aw4Ysqi91E/7gIvVWdQUoVqAadJzM99y24kAGcfAAlYhD7++2w7mjPWzvtgJ
4+knUmTjWnzO6NwGeiLg+F8H/KS5SlUMBNAzHzGzsgNN7uD7QNRkT3jrLJxJ1+r+eauSKJ7SjWw3
LG1HvVDYRbpYSptCI/vP6HBJ60W6jZLt7a0SvF3qXjPg9bc3KKqsbey/xBo2Bw5jU2VfcDmKX76u
imV89j6qSVG+hrqBXhLQzd5A7ZD5yeUN3CfXH5NO4OBefIBMXSLMcpnn7zWgTo2BTP17DhnMIHXJ
L2+LL+U1PiYWKY7TceA1Xau2DBmylXK/OzsPOzDaOMK0sXnH26ZTRKiTRMyh0DLCrk9yq1TOXMCq
ncbUL2JVc61H8aE8i0cWvKr8XEPHT+Sd3azXkb/kdzSGeutVsc4SlYjq4LZjfGsMWGV/b3dFI386
1Qs/MnFiloOvQ2jKSa89GvDhMT4zJayEgIupoyn+ZzE0xdVr/Gkf2Q1n0ZKnut3lnFlvjcxaKje/
tVp/zROIBzm7goQQ8XRmDB2lNFnhQ2FPSka+gnwC3mQCgFKl1rOBOoMMgrJq/UGd7whLjgGUOtwW
P84RMaXLH6yMnVTAVJfOtioz8UHFlM6F57bUYuSDqxMvCMoziWsFHfbCubDgS85f4/YhNL0WXgpF
fs2y0ym/gUyIPzM7lvu0tsOSstB8jBNZKhTNWd6+SE+k/JmhQMVxQE9i6opbxTnthiUTwOyJ9+3s
pMynVMG16aS91nMnIkFjAMnPS4ekW25uAfWiVckedQDUadim3I0/LkdLiGT5O700MnK3t3ZNi6aV
YstygEmS77h1qpecMe6MKWT+IvKkrhUogzmP8fsP4ZGXFAYnvTZwyaAPiJf9XBqnE5dzJmgV0v7M
FeeZhyo8CSlACms9O+UUAB/bUvW835yzvz0ZvTzRUyGT5N+5+iQOFpa7KqpsIduognYJmEaHEMeJ
M0xbSkrlLW9KkrjSkkWbiktM8i4BYZqS4MsQan4FxL/A0B4MeMt/hkn1UDSkOFT4QsUHFbMFAeva
A79s+fV8M+VLVEyu8xfL8YcdKyOMfKNisyS3bSNq+0Vw02TL1FjtwOIagiBDHtZrzxsrie7IAwOL
UWzh4sk/+25yeAO6YCSdsjQkCHA/ALJmg/KQoo6IaHq8wap/wZCwy4GPAJWEw8XgqT6WrXniLO+5
aMiI1ofbnBBezT3WfYo74LjVSn8EDhDty6L34cf25AttYlPsk5cVN/xq60qrnjNPqvLfnhP/S9rQ
t73OWWMXmlk86VddH2hxF+6RCGcMkbw+NwAvxnY+cpp/nT5KOQBL1FBvZMCDKgP4gnj9JiSprhg2
PhBnQN7YPCAxt4IUZtGTV6DE7ftJBYwN5gZDiPaOM5wyTemdGtyAJNkSB+6b24aOlqxEBGQBRJy8
NHaaxRts4PmdTSuD77kwCq5ybZ5Y4ciedPUB6il5biXldSfZOxYEaVMhFbs2FF+HQ7MNf9pEHJ89
viAk7O3dQlTy42ccmPuerLQFEqlwDeH8d0dG2DghQf+C1Aw9gPwW7thkPZLblid29whC7+fMap7c
27yNYSa4owxwc3KwSwelIjISScWD24Ub3LUnugB7TsilV0lhyKLwBCyLa+vENLO8Qbl834SylfZg
AzAmnbMimapfELb7jl3ciCHEn4kufg/YU2cEl+iCHs8nL84PkTV7qNz/17OJmms8IN3r0oIwdi+H
Q4VTBivn96yYqhiq6/BBm8lKGDT9SCjNct80Xhje3pWEgRWVYIqDZINu7H1f56gQC/VVIEo1xq+F
ZKh6n0qxVdVrqSOU3SdmvmrwKxO+x4b4Gja9HFZXyRuDRB0M5gH/WsLO+gy6ohNBQyDUtNyWiJB6
OSAmmalIZgXE0a3bDBDmOL7djNar8fUhoY7tMbfTpKKYnkTONMAwOTFFWlhAOIZFJrhSRuGH3u6d
Fnrl4nXtxosTs5qWkNvKU+/VUdx6BSXLLKLY8OMPXuDpgBsciarZgTBJYKedEHmGGh9bG2ZiQn8d
symG1m5SJSr52Pg28gcn/za0S5vNwpDAldBBDgSOSiKuFe+3F/YSPlDe8k50XONKdagxIXAXIgDS
4lX1AIxi3JCaZERn9njQ7OMXAjwaOE4Gl9FNps7V1JqWaRxwNi6p8kMNrintupO8blQM5Z34eYpr
uz4Ohs8dOGA0FpsRQ6MxaVWsYxIw7mb+7EweurHsPGEnn4EHmHvt0O3sgdctg75VR6ApLgARX/YA
+zyNPxZp2uZEttxrnw6x8/ll8BOBXeKiiGhIWztxm8A9ULNiBlBKldYmHI5xFeXh3mJiUGpljQbD
mAMrEUlAaUDArUNlnnpkeLtPy4BQtW55I0EmNgz7XE9lzWQStlFbrwn8fwoeJBXTED5ayZCJ1DSe
T3nOwhpb8x+GypxGKu4gK6YxRhpElJ9W2qZyP5nqk1HZ2Q5aMNX3FIYUWt+BF6Sq6Q25QQxhgxIs
hNyVuWapjqlnf5M6UfSoqAu5qNBCCWsAgDBlxO9j2jHG0Fq2z8WuI8jI0J8im8H+DgTgSNVWhAdi
13qPQEFSr1AY6nADnhfYHjpShz0Rx2oyhgGpCQXoyzLC4Q6TB1kH592oQinEXRSyepTOa2ZTt4Sw
2ofONdVs9WtAjdkb0mXo6z8qwIRHXx8/sv/fhRcUUOxnetfytfEsIufQ9Dq+Ud9AzRvEcj5kHwTp
aXbI18tqzye7kWaufYTebcXtPH0GNMNASJtLpL7hPNgMXUOz5oqIRF3r9feWGPyNo0m+erJjDep3
LalSwdX/8K9Yx0kjjtRXx/LPopvzm+FmCuKhm7NlFGhPW5XLKupYwNGrUJ+3rzlr0S4FzFx+SeDc
HtCWniqdlCmJiqpn/kJfgqFjiOLwiqb+Mn8VQdjBbeGcps/At61RoJikR5P8glhivOTeH6PuTFna
yAPUDGXOGw8JKMSZB0bGB69zDBAthndrqQ9luZTPG8+SKaAcU7x35Rqxzn4qGSiMk1t9rmbWx/IN
9ls71uZECU/ks0hpf0UEoM9dB3UoOOnvS9R+a3mHsOyZ3OyGn81PlKRpw/9rfvZuAYMVG+Reap4e
E+a2wE8EnRTTSWH1nG7CLnidPmX+cipRTZL2SQ6giEXHIk4zzQcjsDiNFqWEDvp94REOwG6k+PvX
6y/eq1C0+WnjL1NdUVdCl3ORl5koMeG/gyp6JMZRH13LOfEX3k2+nrE646QVuE6BTEc1yeCCdf1c
FtZ5kthVEyUVUiDo9KutKcJYifKY2JnymROL6uXPstECehnCJl9w/n+kM9hhKbduIXaLSHMC6jp0
7Day2VCd/E7WZAJRs8RaZvukirCQNSloANPzMxTBoQvxwJ2pTXKoaGsXlAgf2A6pNyJeLfoi54Qp
dtz3LPf6VF6776HvfROiK11P9oqp/lnmE81tR9n+1TpYRU83gAitGueS2flsYbWt4kRTAwee1WNE
oLfyZ2CMzHKT2Irdw3LLsVfZTtJz1bRuBHt+bGdk517aWqZi6Yg/z6v6+gw7uNOE3X0fnWnEAkEX
ANitPsd3txbbnkfJ1NvT8aVw63IkPPSmOh07KgOa2PIOJVV4EfZmpqxyP5P0cnD6WpMqPTbmNfgi
Oj1TJk2IUQ4RQfYad8drWiOKnu870Q8LhVSRJVGq5Reh/9KYmnpQMdI/yPr4qgW0Tg2ddZtQofAK
52NWBu44BuEbnAUEwheVthXVrXptwndwbmAcMeUafx2B10tATewPNLNklONdH3xY9/fNWfqx4LSG
krm+BJ/dyf5Mcwiok9vFSlS+JqLG7BBuJRrNL+V5lq8rhPB6g14/d47oC/rH1Fl/2o96+jl8UAO/
mSlxU42vCS+mwcDgqUHVtC8fTOkuTPsE0EdEYsw/7G+byWwkyRylE6hdRxHf5AyKjDQ2UXOApyu+
x5Pzg89lc0V7YqnA97iOiDn2UEc3u0/gyFuLTTtVuzQsGip4ZywGhi3HiHAs0Qfioc2pmKQiZoNt
aKUL5rlt/k/rCeeM7cLsriyO6ANb8b6Y7nh31LGfOMpeTCR9NEm5n9pXfCbFuLrqdyNIjMAejPL5
X1xwrtjIRGRzZMwY2MWotZ9KufoilMyewvbIhrnTRBwKXv+qUF44Nk1yaowlIermeO/CIIZV2YBd
mYtrooWoWZWD7NcwzXj0T7scAa+ro1hZ3zBtxhWLUl3r2z+Hwvwt16fhBGmo98Qx+rar1qlSQg5t
fj9uizCu49h82yhhIJpXdfejn6MT8cqobpHxwzruI/qKx0cCNFMKlQMpzDKXLIDfHrQr7l2IVssf
lCm4tzdwXk8+EHksXkVn8PWls3cUBFZiAIydYNiPapwC4rpQia04Aii1z9fIiy0PXp5+F9+929m6
frGd9w62b+WLQgu8ng04pj9p+A0ju8tPQaWiuO50el5JV8ljIbdYJJr/D6lt/DVaGp7sVI1r7Rvb
YOhK5IUX801YXuWgUSROPEZghamTs1TVNEu14lmGIsopDDKK1QKIo4yLTY79OGaBnDD9Wpqe+qeZ
1sLGFS3vNC+hs2q/5KSV7OGIF7yhjdt2FxJbnF/1NSj4kk/GKm30/6KjA4+IsRFE9wv5Pf1nSOKL
jDEbUUUSMH9hL/IY7iarkJxavDCKhln73MiMMOZYXDhNy/J8VD6dhbw1+FJdd06XKxIxgtB4ufdx
I5vK4tCpas6ASuCTwQr0LcZMUaLzozK8OhAk3OSzELqbkkhlMfVSsuif4aaIMwB03NNxQXC6DEkY
DuDtoU95H1Fdu1pEiZhqfGeJ1+nuM1Q/qhYEYp8WMcB4v0h24M1iZFk3ocmEDYJDqaBAAU3PcB6b
yN45J0gRgTd8yls33uFMf5Rkgl/o8LtnLDMs4whkjlI8/wxMX6uWFTjPJPrPNBGrP61vFnHvBAKk
l25ivV8cmcyIDuMq6Tr/lToKRnerbWXsmey+88aUAc0J8/e749GfvPxXdU7s4vM1w5aBSvIRISLc
Rp8rosJPqt1wZDEsnXnyqo2PcYtsK2rvPpPCRR9g8l56g1aUHXgkQE9x4T5QSETcJGsX92ZQhDjB
gQbD0z86XdYU942v/ZOtE00vew6T89GMnIyhYtG5jeOs9PZuloztnLI3I+3mgZCm256sf0yeAWx1
TGhWCUr0ZFty4jWYwZxSpG5lYH2H+C1JRw2+QpCp5B2PIIyF28r2NuC38BZCxNDF5giV2hKOguM1
HFuZSU8iyUcaCdqNN2j7kvZ8xVjFfxOUxFsp5SACDioVAWXeZN5G7bmmU/1S9gHkWNsxvvYTAFtH
Yj7DEEn+M+CMFScdxMvlbS4oNZN2valfpYM/rat7hXbO5JQrp0u3UkkQNtC/aDVnKWZh77l4xzIT
Ye/c1rEe9uXI7y4BVzEDon8QHYCz0wE6ATmsPPXxcD1uqzEITkt4VHflOKBlD26i/KkucpeURiPp
UIk2Pppp0Z500jY9Jg6/hw/N6HdJTFXWAdaHew4h1UVM/ECbg5KQ/E02RtuuGeO7mNLsNlB0Aln5
m+ck19RWRxHNMZA51QbQM0EOk0zHsbRUshxKyGpOkE3SPT/ggQteVItOHVTgGhnVmX3azmDDhcBh
dQeSctU9l2okARW3wDY5qrmTW3is7rhGhET63u9TiS4iz8G+5VrTkIDCmKjs5lKHnxs4PlXcTXdf
T7yUiPh9Gu+h01jPV+k84vkP91qYFDczvBivfWgkwfGaI9O1qpcbP2DpWPqhiZwjrbWM7NUzdD7d
LymwO/MX7OstiO9GttQhePyjp44MZRzp+akSax96s5cCI5eLcKeXIvJ1B7Vs7FTEUlv2cronM8j5
DHRYuW2Pp/Ft4j+VIb++zdyc+ljw30eDcjs/GfYTDRPJHvJ5Oo+F6sTWkJysFXaiubc3hznUJ3Q/
U7/eHCZ8Z81ap8hOU70NcuILT0s8xwj+pFPr+A3/7Oy2TmcP45dKmnBKOGaWHWAEKozKZL6GVvYz
QzqSPDpOVz89iBkZOx5bGOZkJ6/CYuBHXpxf9oz6JosvvgORBnr2iAy30lVsME3l0PASi2fXBpq7
K68EgYIB+RxjzqSnKH7+kZzJQ0Wn/47R3wu22d1lJqUANgEgNrEwfo2f/LwbQEjrv/LXAKr4fqtj
SARm7KV9b5kghNqDYDofVBZiqesRfyRz2EwmlAhzw/FRXbRgQiCgs9sC7b7cpCN90dq9ZmiKsc3A
316IfBMvCU3TUcJHhIXIdYYOZ8tBPcBJjNHwfvf3vU6O8XBnibJJh2kMUMkFfSSAAA/QvMuSlsTO
rts9JKF8zC5T6phql0l8TSGs02WCp7PiuDq6BMVNw0kNoTuG+NQ3MRTCrq4brTwKJwi2OJKVEug6
vzNI45zPL8NXja0K5INWSyRFK8WtkVHacBP6oqG18DIisASa2/3AIfRTlEjnPU9WPKnA3ikJKqvJ
8zejax2YYtvYmQ5Zz/LmpsvziRvI1AdkGTUsWSuxhK/vxa+kgXJ6HmGMpXaEn2qO14aGXqZLjnDf
2ol2CtWVZkZyZYUCO2PvgrsN7GKhHFK7hgb/HJCS68HzQIbsLhiPgAPM1hyXh8Lpj3i5s5TaYyFe
A2ozjILVHo1oeVYqB6WXY2JMRCHjfQsitog4od3at/LIFw0u6uixbxg/ZB/qV2bIwSbfj9/Dw5yg
VB/zxCMjE5tiHNFjNEI1O9Nb34gEtS+IzbIAN2T3PwWrkjF+foy7WKG9E1ErGk2Wc7PS10ufm+O3
WZWHi2rqAqsJLvH/XEDDz8QE7/pL2CkAtlBUL8/kGxY9fO1AIxTjobctA7gCfPMhKqMK7XuNTdCg
Z3ZNPDMJgKjWE7ypJ2yzScbBeRMQWa4Gyv3VhlpqlRUxWY1zqF3uUlVGDIhGgksbLI4RWbdmx59m
Bge6jbZhe69XM+4OegON0BK55qGUdI4Uiq8RDDHcNrZfiuNnJ59xMIC9nrOU7+iqXo/ux/vofR2X
B7vj29TuDXVeQFb0N/XWkVymnvgbehXP20jYCQ3XSYoFXbxnHQ7iQUNggcXto23p64ugsXP++Tmn
uEqbGNzTs7rVAKYMdjFtYaklhbMaSPBo0Pm5iWVsA2F64pa5brp/4i8eSr4oNyr/5LdqLQlfxQGe
deJaOjcfAULU5ICDioqXGxKHpuRs9FzaoV1F845jZ4fhuUHE0SLsFw6+Z7QYYan89Ypv4lAxiojH
mcPSCc1LhU2UpAeP+Rn3M27UEb/sMCTfnCZiPxyetWbIVSx/Kz4d3vQuT9AafmmwxxX1LlmfO796
wyodYM6sEySAfqd90lw6MKY2x9TnmQwpGuwY9hpzwq7Irjk84U0nbUVUK6DNLq7HgP2+mZaF94gg
Xj1UOEDUr9AIabECrlG99S2gSICX8sPNNA8kCsj0DGZnSHdHzUW9GOF/ht9iNNgvYbdhCREP1/7j
mzkEsJu8sjRwkZ5GA99OE6QshGmcsArCzcgMl7Z74HW8BfC8MejWZ8C5rdqOtX1qSBT08YI6jBIP
g607FnuXY49asfPr99rQqljGKUDVNoM9HJzfVvwMrCI88wRn/VYUgBI0+HRb8+B5S1s4nhFxtTJN
tHlt7tg9nFXTw+axvzW40+qpFJxy2d+iI4yhcD6duRZZ5utX6NkxlLmBEbSwnmNzN1n+4DoZvtHl
eCCDrV3xolPIKyM9hf575gjyz/bfPm7ByUUbVnf1tx2giwmSYcGgrrJKuXTuLXvMiWeV0E5jOVVL
ThbDGbHNJPISiHuJQoNwcPYzPwRmdx0rl/RuAiNu0PviD3HDkUkPWgRdCDcuawPfuDA7bcsiyxgx
kep3yroB6GfsKCo1uJVRfbDzT6TUV/zHRwJ6egp9QdAwQmeMIVkaWAHkxVBn28C1xdvuqPuyTdgn
utHBvd7zm6MsmnzixCaB/dj84D5oL9RR4yKpBGRrT6ivOFmVJRrlzRieeUEDPtuLbaGaEmvwXbHo
8eSczmueS5H/HFAs9iTUnLrWVfEXYQiH8JT6blHUSfSZjhrxHB4KaCCQyM71KDP6M/lIOPWUB7kR
FQMy7Dc1d7tPBAnHvVqhTM48ImfYAHZKfCdqIfmyCbbmFv6cl5OCMzlOmvyJIfYnRkv6sievGwhd
kGp4jU3yVXbHazWC43lB/r0doVbVx9IRyQ6+dl1RuEIYJvLC4hXZlh6j3XTdYOeUu5sFMkTsLd0l
50SV85g4K6vqNmAyrbLBly+PE00TsnQ85/WLcuQGDt0klMaSU6a8IKwmLMGnot9xtpGeqE3ljqtB
FlA0yMO00kU88ir9k8ZVqdtWNNSRbu4s233wkQftq+GAbJ26cH53tSKx8CYmmAVY8i6AHRVeLRBO
VCrNh1jigWxNblJO7hEbBydCIpYYB5frqb5LL4a+3bWWtvuwtOdJ4CeJvVwoqJC11ExtvOgCkOIX
ZmTntahoRZs7AqnnTgENWZAPioETqKzF95FeawrlBEvIUQjXrMzfVCVd6FYuTQpomC2G7ksuq+aR
e8HQ2gvF2a4WuRvC9LC2ySNNKlAxVxJMifEf56bIMixoWMGearn33Y3AP0L1v1HAIGQFB8ZFC5kf
0BySrExOl+q2TZCbLbmGw0Dv+SbQe7bkuR9hSnttw/LIilyM7ZPgGO8VTDJcYW+4LkmHsoKH5Pkk
58zQeDbc9w/jAkvZqwO3q3TzrDdQzNL+K79kbAP01F1GFTo/HU42JPE42Fy1WNPturdIKusQOS3B
L70nH7oNkiyUhWkGQEqt2C2FJiAU94wp6WHfIEeL7uivPFJNShXXoBGAS0/s1/OGXwM+EBTFuILO
M8vES1qkYncKiGQ5EXbKoQNqdIos/EN9B1GpRMTIp8hHBnBhagqEDTXAGCy9+x1SXoTLZFIIaQlF
aLl6u6g22OQtO6FdKIMMUjn1Dwh7QtLfWeafu/faG+tE2AeNB74/l58LnhwjjJ1ibkMZyiFRiT97
LfVb9/huUuo0pmdHiqMD+xO4VXg0mIx43LySjQasV7s9VqBXuQGmi0XHBNC9gdQvDphwtrTKP+oP
zpAs8FNoohCsHSQJ5Y2ArtsVAZtdgRLCaI1wk4KahinqvRXdLxPUW/0HOnnxAi9J2uP05ZfRmHZX
g5FDYJN072vpGi/8VW773J0sG9akZYbCO5YFvE0qqoGkY5sL3vGRdN9l02NNUHala9I1YBL37sKx
lpG1csI11aELRbmmnI40BuLmXlBYpFHs7cjirb41FMcqi6do8mBDCXUvGcpts9e/TTnX7+akE+uS
O9Bbfc6SRW9GIZyWzQaEWhHyzPIxfG2RTdY8cG/ZlCD2TmjilsMGl4uRu6lKbN9j7NCpZa4xJFHX
OlS61hZLB1RQXvcFmS7znuyf3qu115GRn5fnJVao6rH9Z3hhf3hPwIaCv83fW7W7gXLGTl5/Mu5h
ngEJu/cst43G77rB5oscmu5GoREcf4COyvkuEwahZ0MYiqauB8IrMTaSh/FwcZoPNrlu8ZyZ35nX
LW1w6xPLv6HkdeC+0oXRixDGhRJY3A88WeuE2t9aBbVJUBEADSmHOmNcNIGmX0WmTDFUTR+PqnQo
gu0zNiJP6EOQ2RVqCdOB2nBcjwo78ShoOZnHilWJB5slRuugFxn9l76yiFHDPz13XWMaGVg0UF6s
r9ubX5KU8NtWd6DRmU5Ia5kFFvtEu5wVCdaIXzXwHH0C0iXLOFX4z0NJvKHZds1mGyKtGgpLszNS
HSeI3aHlby0nZ79SFhBDT5KAvbHuTXbo6QJ/++88xiLWgeaY/OEuSrH7NidFcPj/AbyeDvek6y8L
dy3EjYK6khnJa5Taw04uDnxy+en1cUBj5Ra+8Uc8Uwi1+WNZr38VHDA3b2sAPFlDtR/eKvwhH2sl
sgT5xsrkQJvSX/5StSZ7j6QQ2YHqxfz/4kajC5danx2PzGKxQyfKNtpAeuzAOcf722embQoqzlKV
ipu5UOQLtycArplmdAPD75OtsuS/z5qOjEZTh4NnM+4SMPrCBt4HbCGlyyoRRG5z0/OGEqolypo6
SvI596j27TaLhA9a4smluV++AlmuKqxqrbuN0gLqUI4Zbq3Mn2XZlE9I+b8/7ymeXXEuiqQca6fC
rzwltAsM9A206rh1uYwIp6pmsAIOpgVzGp9aUUny8gU1/6KW0D8cTdLqmYwRcVvsJHst5FmjWfhR
LHUXd9P0h3z7jX/X+jI5+JeKWnLIBZMgzP+zMM+7Z5LXL70Ci1dYfT66LX9nhFqOfsZuBWhrA4eu
L3AFeEyIV927hiYVbjcw6lALmT35Qrrum44w5+9nsJmdbiGh2Hckj8fWMYE5R/m7qGk0eud/SbYn
A0t6rFLotTVOf4ko25j2wbtaaZfjffIFzftts6DnEq0r6CTKfiBqsCaCv9FQtckE4zg+1NFT3c6M
pzlhLZ87vFRlXYgtMYXuUlYJj33bPyMsbllmS9CErJwKL8YFmIrkpfX9IzxYUWcHUHrQ/mEyXeH1
aKEP1aDh8KE/GzddNrgQNPowOXLnuJ3xCyfJio1fjahUuftglBDHaoJjhkh67zbKW6grA2LQsr3I
OHcOn5kIfFafI6V2USjgw9Enb5WdJnumnnauyOy0AZmRw00dvAfBR2mNMQ8WxlFJ6YMobDwm0iip
HLOzSrC42ZTe3fktxZ6UOfkb3+ByeoPUIg4bl8mUOGSXupIRWh8f5UDsNOVCBLuAdpGHB/ZxeeMT
XsTnYW57v5fM7fRnvIZaGgu7n82TDcy9VHYFsg81o2NLnnvoliFg12vB6rSIQFDBpTKFY4HWhGUv
iKji29wO/s35pNm9MeSgvnyj1aKiOIwURbvj+bGvg9SQdk+FbI/oug8Y5M/TWq0NDbXZrWPtkc+O
zMPILv4sLrmlCLmzIh9mIAqihMbENemCNT4KScz8tNK1NRzgPUF1sOBtjseheiXWiARWjjTILMJo
l/+EmTHp4EpGw566ukRdK0DteRkjk4GIwhdc20sB/nOSpArO+3rTJ9a/AjHADyVKaZgwCtsz8pMu
aDsJaZJtMQHfHwobjo8X7MngYVSmwtd3DMigYovV4rGIu9sMtN/Kjw2TBFgGYAyYos6RKRwjo5SQ
24M5/yUq1QnJNbZM+92ueiDQ4QOgjiw/EJcL9rWUkOWhUYDZztXnEzTxusjN3krq1/Z1Z61cgeE/
1s2mXwCrmcVADgu7SxvaAA2JTEzUqsL6tUhDQXYwSslBPWdtN0AfbZqqlsATNjFf8N42JrTD00GJ
gIUMrLu0KgRMmCDOvU83B7Z8ciT44C4IHFCaydgZNzmrTbXhRO4CuctGuijPdmQCurLibjH/qlyr
McQP+JhdBlBgLVNsinZKhjRx7vrK4DYTXwfyD4j57CJlK6JWzPO/XEset/jZNMgNk3iMbu8WqLNT
ggcJSMKZcotDO6lN/eSIrZfJTL8E6Yrak6SYHWjPWwFjTD5gvS9M6QjgVknMd0Y8YvOoZn9BC5kG
IIrggXnbFqNmglf/YXWaXDQLIjWJ4JWtYZc3UP/asq1Vlz7y5anjz5p3VOUnpCMHLUSqSv18jJgB
CQuRBo8g908CIyA2QRPLd3U2lof+jbQbGk8rvM+vb0BSoshr5xfH06rl0EajzfAAOGXH5yNl+vtU
5zZ4BOKl/P3eMTgrky7b/5znMZRWF2tcL2bcYR/naxhavZODM0xHH6EKTV1z+UPI/+pTzilp5+aP
Hc11c42b9bYfdt8tuaCFPcIZVpBaIEcfHIqzHGPCplLZHmeEgcOIagNlOMO3RxmNShb8O3y02BME
KfXWWbH3V0qXXOf9FHqIcFJtNZ7+lScOZx3RtBG20F+Coy0gwx0TKkksXEFBcH5gBiM15L7GxZke
WacFMFQxma1uRVH/jHIVdtiUujK7v7PjtFKViV9eXSTRmrPSEUBBhjbzMTvEh4ndJJ5CKjTRfYJN
Weyie3Y9dJvt6L/9mKh0vArYMXRO/o47DwNGH41hC+rOr+x4Y4Mo/kPleIiK5K88aLBupB0JLGbu
toqbLtUdLZLlUEJdsbD9+yMjrUYW9407gI6FXxo/EaEgECXYjRhj4eQs0bWe76dQhgT88lbM1fVm
eOqSAmBaK+2GDvIZsJk5ZEkmn6t/c6aTKavilZCaXFJQ4KO1yIMCa7Z/FWVNpDsZzppiOGSLC/du
0oAyOjua0Eb8nxVZR2JkRp0Nea9i3jXF/fUf0+TDrYbvd9zNrh0Mzdca3p2/j6+fXTfSel/46e9E
l+KYvR1BD65LxruDxGcWEfOz3WBtD6Ut6TVHAdigm0DBNJUKbx2GZqbXERIJYiZ/NkAzDnCHj70W
unaEceqBUDdfv+We39OwIblWRdwkUPHMREl+dprYni0cAs3NmCxSIZ8+8QnHv7Td5c57ipopxDJi
6sOfPVO2kdSwlIXjsF+KEXuZzAvvEMxix23laNSrk7B8z5VhnzDMvhoTAfni5HcztugQR5LOz6xN
mqnhwbkDjlalAaNBjDrNiKetSzL67Y07UBTugR+wijI9JDwltpByc82eR/4KNP/adBPY4FXDDUk+
WMuVoE/sgKKgXOoF7oC5sNERH6/7H+pQoKgmqYczODfZhh84ahLxAdSE+djIwEmcLXPVP50wdDj6
yMNyAmAblaQ+nbBi81e6puvtzdfnJkhLDJETQLgWFxPLQ+N5KY8ey2o3Yth1qwSJFVSiughIKtAT
GFIbc4U+ODEkINAf+Z4+GoZ1CyCDE84fMEvr4xo5A7xU9isMHWSMcr8k6m8CnoKZke9nJUwp37mG
PtDKDK0qwMTUIRxR1J1CFF1owpnz8HiJOdL/py7J7fuHjkvOGn2++FLxloigHIFSlXDHyad8P6cW
JJl0Zy2HgR5rGbSXYBr+T0AdvQgkbOEpirKUQl4TDu9Y6W6EQjWG4d3bFe6xvGAdtLuOjSQSWl5H
EKelCfu4JaUWLzIcVHyzPf0ltjqXyQYfzfx+VRWlxGm6JSc93uisWY+dPaiy3kpvyYjvxMUEquDH
+N1Ck3JOwtIo+acNKGPUFT0N84KmytKg2VcUOi4fRPXw61dbBCI/DcP5sXPqTWBdi9GoOk5En+0M
I+B0hoVviDuJiolr3E6Mzsa3Eir9wto2/zdd5YLDKxZ/fJREXNdYLvMjHFQJzcd7wCp6l8L2HJ6v
jZP2kaFY7NR8IPYeJBG44hfLJrZbdxqZWek7LFhye6vk51OBbbIgBeCSNelfv5wn6h6YqFtJFMQ3
D1es3vB6wlZ7qYSmF1vxkls5Grf6mv4dfu+3goQH4am981e6dCjzFmRu4IUwG2g0NmJ4vbIEUphB
BpBAHq2sCWDTMertkyIM/J5Jy7jRJbh5vDjr2yKqs4PDj+QcVzP6H2bRAzSKlJRoYH6HHhq3K2xH
IlnOfi+MhxDi3Cfs9XbZKjvi0LMLQV650HiZjYIFt9Yoy7LEQ70+OHWo1Bx3aGsAcZ6svHNDuTvy
7pimgOQWJO+91HC0wprMnOCqwf+hA50tP0P+YPTafRo7hD6lEqmjfgoc7l8/AO+pop6ygOj2xidO
qrgH+OkEbdzGyp15N6sUSNiTJgSX3aXvVbMvs2cYSFf8NfKvhggdXpOh57aefcnU9UkVqKdsk7HT
Kw2ITodXPNxSOUPHX9EiOL/4UCqQic1J6B6n1CxgFXUiFUTBFVcStwiDwyVbWaL3ESMseDgGKFLP
u0Trar4AX5RF74xrPOVyrdZZ+bQQgJK/UAyt+5VkNu0/62vETAaxsS805Qcp94fejKofdSmf1kpz
6gjtMlZ78cDUIya4OnwCQC5elbO6IP3V2WGjNLjcbjLnaV9TNublif6W7H+GziTMQrt6QaoWPDds
tSNkozAIoNDv97UHFphRZw0XvV1gbebgEdPSRChoZYDsHke8N1rvhKMFE7Zpzyxj/sfKsHw/9l8V
bJCLl6kJSKuqyIZIXvcB0aTRylg4d+KODT2a4xZuqRpWqp/YE8J9rqA+CfasEXCIyOoVdASlPoo+
JtwLmDaPzpNlw33KcWgAzsVOvNAoLNuPnmvbArKZ2Z0fSP3DYBewrHGce7opMvTNyO1JEbSb+Rqr
ySzv7OU9tITGU7/aNjL8F1ioBStitKWn+ThG4cM2T24Gm5nWK11JXzG8ovguN7irL+VIW58Muds+
rOsFZz8IG3SzLA+NMLYtgtO0HjrKZEdDU//QTsS4NNmgy81P4efdoKUlPmaWttnoxoPggSfkwJ/r
MqrvVOSFHMkrNTkardmCBoHTdkqTDXv8oVzQyVeyOHIrHSyftUvCYU08B7J5QSqll5fkoe3A18XZ
ZwMvi0EUUkWTXbPEqntS6r5K8p8RMPRcg1p4O6SaBzZ+PvGAzEyjI+opN3tKCWjimL8tOFgJR8Iy
CLWRrG55OQnpXDgaTguwzI8pqu6Iy3Q+C78PsK1Dl5D+OoH17dFNpIrzjBLdRjBj/HEJfravZVln
+zF5WZh2344YHROaC8TOBygwBBpaTOQrQGK1dMrEQCLAWl30C3om4GFp5ummxR5l3qJ60gtnYBOj
GszZd1w8vpxoZmgj3gstdjehyM+42qEVCHVDhW9XgNkLdO56854j2IYIfLNxVftdh0SBBaQfIFuG
xrkusHofJG1SJ/pav6LyigqhPnNpZnBqVy+5dVyiMYPdgkKp+Wbn6decmMJkYUU2jBlvZzSCuQsI
G6D9B5VBy1ijSSy/QS7LMLnDJZ94HH3NxSaO10jt1wzjQ7TZEjF/rSaI2Y56JaXOzWGpYPcsZ23X
AL67pgUp8g8lDs72wrxY0N+JidMQaSdQwWPMbnMIE7V0Fa6MVpD6jNmTwoqlZvd1OIVWdE3Gmvpl
1wndlV32StfjuzE/gLSA6gEBR5KsB0g981/FjiaFjf6P0Ucsqdz4SrF68RPAx3d2/gEpy6u+ghT6
pVfDzvVXRw6WK77JbV5gkTWCgPCMl3U7HFfQMzKlHWyUj617WYu6ItUhzGshoiKg+3YenUHeA4mp
JrHHPHYMWN4FtpNSJnZrjOdCQ87to2s/b33BfjI8ZcW5Gtv83VJuS68NHJnoDwmV1Uxo4QLYIsYv
AhqSAoKeLmg/Uepn31KoFzqzdDLduUXl6BXiufddAmwglMlQgiZ/2w7gun6NCxbjmbOiflcBM+Vm
je528LEynEOXpRdFg5Lkx+bUPKGdgr2iG4at8+zb9NgF02uynUpih6Jrocj2s7LTk7w6Z1pxSDD/
0VLoxvl/AmI1bRDoCyfXm+sUJNOaDL+3kPrRdigkkrINMkt9zW2bM6jX1tTCyLTtG7mIeEPPIsNM
fdjxguk+qAbNJhRnj/jQ6sU5WoCJLpYoY+ruUuR84KrtGQDutmA5h9/MTSiXS0LVv08zvwuSElhE
6tIruNvxRpQqT+UUCEw4oFJvu/dcYKZQPzz+64cEI8QusL971wvdtZSboLIGiKP8PmTK1QkNYDKX
3PAu0zGJ3pMwbz1KM0Swivj5o68AWiSdePuDAhE2GtZv6dao4v6En+M4j0o4/ie8Lxwi2kaeQ0IB
W5HkzzHHQzshzl4GQiajqElXGt0uejTWPxubtoQeyd9It0NJXOq5QBKskECPmi/fhKXib4MZc+sB
raH1lN5Bsxbgc01s/uJTq/qpDHe09gpCLH9N3yC+8s+JaTj/YYvUdSEC1c4iVik2121VqF+HgDd8
9YDgejq7aIM786exNyqJa5klMkyKO7URd3rKdA5xOUYZE32Jhlpm3mtzaPmzt2MXFaJtndpMWnLB
kWxehlrj2o3RkegLDSiuafo6UJ0niCeXnedsXEDBDncF5N0PAQ0ljRxC2fJq0SxHUplqr7RV/1Gk
xUoFOonZa9vtXWBjDvOY9lBt7H0NFpk2fZJc3+VhYXtKvGz8buOJEsO7AvCHhHoYtXZjsI3xCD8n
icddBVXrZrLGyFNAo05LFzcmQJLRVzf8i0/GvKkLMAqc8WjSGOqFw0qocIe+bUp/Tcvvqr+E2mFg
2C+CYbmq+81HEfOcr5ME8+u2N7tCZy5m9k0stQawiTuVY3mEZYQNENvtW1jpvbTcbkwWVnj+xoyv
iII6VC3Vc0zpEntAoxMwtwk7s3ClCVPfdsUsdc6VEDLu00SzExcUH14rTRf3EF/k4n5tGdbFzIYE
aFu3eCwVSYtZZWOUwV+IYd5ozptJqBnCOuErunlqev1rcPmmtB1HcgMX0c9GN2nq8trqEwx3tpuF
so+WCbk25vS/j8SfFalV22KXqfkluYN1Ak4QHUPuu9W5+Wa6NDK5eokA6hODKh+zrdd3+P867Ksr
Bzhe8S7lylX4CNzjmq/pl4yCBMOuT/wldRl77WarJ+kIbGFpzvrJRLHJRp19OZhzxi5GmkvNNwxq
Mui+97XEE+o6IuMrb9M+KRRUizIWMJUqp98eMQpM+WJ4D293AU7KYy0QRDlZPZwqd5DlrKj4Domp
B5+wZXR8gUIA39whpWZgiA2qoEJ4FibgmcSkTQ0I3SAti0TKVYEnK+fVLz7rR5LkprrF/yMfwBeP
OuM1HoGP8MlxngqoKLqLncG40Scvsa/941pgxJOCml7NJCMUjJDna0fur1QFDNi4GyBsfWLRmuyl
jEloX/OssrUnZquAU9pQY49SooS5McBhVv22iCMc6KG3FA0Jhh7CZDhn0JWO6SSBy9Ju0v5GmR00
6mQS0UkxeyvNyZWGgvhTWExgLRd/2TSYSVZwyyzR0rbU0NyHuYalSFgrFRyxymrMLmvba9Vk14J/
sFGo6Z3uD8U5tdUlLwRy6ogYLZAK4J/mJm66WO7YI9E8s8HoduVrWcX13Zt6n8foHsc0tXkR0h4Y
ajwPePvIjK98WHkh0Yk7Dfk+bPaFtk5DxgUmDxgosb0sOsap6q30lhhUVGuFyHlIrDsbxTM50GSR
or4dSXk7LItK8oHiRrd8rlZq8USu8CVohA4vxL+Yr2pXR9fZoNDckZ0gzHdR/sA+2PW83GmqkCyh
IN7WzfLP4SoHh7cxbSqMxwY902iuJP30QY00gV6yh6HZQjnC2fF9pGoJJx1v2FhZTAUWlyV8VzHL
Q/zG0YBFP7juxzUQU2gng5pap0zAwCiD4wQfvX/atBQdXnibGY3kYiKaJhe8nvEAAFcPD8e2Xm4Y
ALPgjRneFhK5/eJ1lCU3dLVDj+Bn//vxxHD1dxqeGmWD5C7r1i8wQSmlPELt1aENyFZxyZGzbA6M
XpFEMaQkj5Boxe/Swq6nDbK65jwbWuirlcikOfPe+Y+QIvG9/0XeVs2JPm20jlExQVEtkLE85Mnb
mL5OB3kfXzdwu560DvliLOfGhvAmZU9/81gXqlTaG7oZr77acfin3gJx9PGBG9TjT8jxK9uGbESV
M9YNUWI9MAnHTLYtVaKTINcumCRZARhCKgaGkCpvKCuDyy+N1Zuxf5MJIfuFICExyp9vdXOxbZX2
Q4vI8GkCZkAZ4cRweDVdJBYMjNuulYlhdgGR1PCIWCXC+GSyudBZMaMxIOWQJ1gOiXXsMbgtGGfP
pSM0XTdV8iPy7lpVa3I2Oq3AKp82wpNN2QB1naaH/0y1XC9fpKEyZnV7ZK++WAyZEn+yZMLJnFTf
OioPfTVR/a1uaAeHXJ8kCyTsprwMzD4diwS23RGHI7OP8KtsiWNkMFRbhYF8RVQ6kiFIfFgGtsEm
JpXzhXYzWwIprRlA5RFW/+yVFiZElyZOMAV8/thAOZtIw4txPBNy6Rja7piqgq7iwKcdNNcbd0YT
4Dy4yTG4BXPzkfmFvGShng8upbVvSwzwWUpQbv89AH5bmJogESELje1q38spKoHHXehXtmY0K1z1
1emIgub0QtlLHeLIX8oeqJnKpDsCNx3TSSPphbzjLn7JAPD0amUcatNE0395wJp6cd3QtiJlFPSt
HbaZjbPy+knEyzkR7QEf/f5iX3jwReQ57xrgqPmH+9Dq7015IoSns4cVVsECI+ElBQ4jcdVtB6ST
uKUMQy6c9W7y28LUKyzXUopUQlAOkKVQr+hEbSLeCNnasKs18+3d6eEjAwRtAeqMaPIr5/95xhIg
wqJN45DMpEfQAvR+yrR+F7Bf40iEQJiBT1U366VwfzhAnPh6SDx8orOGen2L6ZjrTIfY2dsIZlcu
aXhegoSP6q+oaikxPmnzZwz+GlouaI5PT9vnytRp3oBfFzM7YwDRcr/l3Ar6IgHWMAfVOjq6vTl0
4FROb4/1RLCwwhmd642ZQbyni8ehws/vIzQ9SralWvnMm0hYLNzBI0wDM98ZrcyD6b2fc75x2h8t
oj03CuswgxcRWTieMxmiQlwrQs3bNF8wR29pMxgIjyHosDwPY6oRWzzIX+4tQMZdg1CxLd0A2nE8
BO5NQYb0Z0eWY9+O3MeHBYlCJOCjJMfjM+/VxlV51D7CDQdGp4xYcXLY3nTwY3T/v5soCEbPUYKT
vuOTcNGvdZh6nGy5L8DqdzKeYtzfL09eFNYIw67E/iV/A9EDJlo+VjEKVU2bavENflTAYId5PsWj
wsjyG6bZuO6i2efT0ZFNK0MiH7kml+thm3aQ6MMIXfMq0NLhXH8S2Zl+o2EjAadMp4fA6e44T8WS
LS1hgNeH4argZoSMJxuLxCS6TohheX6I7omePFtF0BDtRW4y+6b5Y/AmF/x3ifcwbc6S9WJtB74P
C2qpiH6DLYYvFpkfvKHLrkoIB99PPSM49XxP0b0vUBdpjy7T3JeLnsQmppmVK2n024MjupHkJOH7
8EyVGR5I2VDtIbK3H7NAxypMl26ETU19AizJj3abri3cC1MqqVSa0HTgaOTcssveceXWtwA7iUQ3
miZKNXYC+duZeqZokCEPgaQfr2JPzW9BXht97My3phUOXAyt0DHLxvZN7rr638gd2oDHHrAaxYtR
O774jiOup1sZhSMOsLbvET0isOuMF7+uKjRo6xGlIfQ2BXdCsyJonhDGnN7TNM7hOgwO+sBgYm+a
iFgwke6hRoeO7Pb19vi8ymr3q0s/T+4smdVMJ47L+CXl7iZs1Y5/QlQUQATrhyf7LyJKFC2ghION
zUaELc9EJC/mO0bcbGczCh2sNOV+jeirK9rdNQUi1idR1plcwDvgHodbEe6IKzupHSgXUrrferFb
AvozDU7DYiZCqbvm/zGJ6AKDS8734J6EyvXwgF5+ze/6YMfbrjX6iavpqWdNJ52Uqaa+4/loDEbV
qw/ZjjQHTVHl2TXOXNNLePkjvhtNyFUXrx1lr/qgDzfpTcvjM0EeOHmXIF6P6Xs3yKWvQnHgQ/4j
cl5Ce02DsBPFrBR22zf2s0SHiKvcW02brQXjBGHWLyL5rUi2KMTX+KiGr5z2UmRMQhhdS5Eprfmz
+AwTZ/ovyXTfGbii6NjUuoFvWNq1SMKQs1pdFyHuTDsfSNMlHf6jLLYgX3q8Aqv4i0hHsRnc71f1
CIQPT+AAe0AQ1GSAU0UBTWPQJjKv6O+hYRIu31JxhW6CAYexJeLMkOgwYefuf9aX3zehCbl7WohN
I+Gpe2B+5OAGIVIbQcYwjnN38SR3Xm+uVwuFgnwl15SZWRQNIlUyjd81GgtuDgEGGMVgYADvg72R
lCcpyYWppP80jqmidDMbDGBmJN/rAlAcUwpQ9bQsvPJwNAOWD347lkh0xHLX2U4fAlx8KAw1ue6/
b8LYJKpsaOi1n0Fcb/d3tubnee2NwSWFPwhN3jFNQFLBV0V4Hm7leGNx1HiMNQC9OLCdtJan8FKs
p0K5u83C6fnBOJVvLfBpeu+sVuXrM6n2SuvVv4398LERrqgBXkDLu8tY4Y5NFXHSDId7MzbUnKyT
gWAzdCQ5qD8y7pUXUmOJSAsQjxWclyYLndgkpLG0jo4TsFwGwFjZdT+vE3ABpyPJoG9RyHNPVTmH
WQei5dQWwls8QGVwgCvPw68WnD1R/EP5yLutB0fstf0FTQnJHqbU17zPIFFyN6sd6YHLJf+lRLK8
utmHoSJ/fDQ+ltJxs/Hz95jrVgOp52JJuE25mAL9nTyjwSVOgZqVk8MLjPWq+dJ3YnW4XMZAs2MW
ATOL7g4OSX5TavMkcx8Xn1ctZkPrJ2AcKvRrL4/AliBgsv43C2hNAkUu8FxASfZDqyC9x+0Wwj/F
PJMuQURek0X37b5TeIYmwYC53OSGt2PC6z5yvQUY7LfIMWEypxJo7UmKSvnvUumxED8uHeL+D2P3
Nm1w7wd9O/UmUYGNMFoHBYDs4rbXLzqJhTAEVCy2DJot2mzGfg+KWl479atN+4sT9YKzN7TtFv9U
RvPqAOT0FwbX13drc0Gel5Cx1quHynfPROPytXoEaV7Hw4KCNGmI07qO9nD/jW7LQBqCb/MJ9f/9
FThVaXqgIcZrDiKq4yYwYdHDXDjrfX3SVKBogLISfYNRUoedShOYn6AxWu9g4WQvbxwJPo9Ntxz9
mZdMm3PEWQHcIFnGLvYn3MXhKKmqWpFnVL1xr4r88zptHodSGP3Le27CP6tebO8oywH4qzKA+Y0C
RTL9VSlZOn3f2Qw4pmgvRvFVNfrknIft2M2kwqbeMzdy8YAeucZTAulOCN4hyQHq7QL6c+8yrXu+
zVBpm2Bsm6EGq5UVmTvBv4ttZ/HaKZt1+sUSPV9Q3xzs/D+XktBS1WA8HztCvyKzJpcLDULxfTcp
MZs+SYcywHGRWGFHSPw4YzqVd10oViZsZGnQMaD+s/05c6B9d0EWU1ZTJUj3uDF6sw+6GbJNEEtr
bgw5PtUzt4Ug1WZCcq7vMxlONTD8/EwNt2nlQMsbvHv1eDPLELwerJdS/Nn4gGIHgRJ3+/hrA9gP
tEU0OwzieIT4FpiCFoQZTUafAj8dv6TNk6YyNYOKm+glwQGu+R8dMIT3O0gNO/P8ti7+WhkI+dWp
6gYiAUy1FEJSYihjnaliROJxOvvm/cur/ZaIGUl66IqplcHNCA9XIRs085W1W/9o+sffpLsahAO9
js29NavXa6dwvqXi6jaflLNWhwZgU3SqcRgCVM6+vljxYTpDYzySkaB7my8dmzxZ42wvK16pjWLy
++K+Qs9mWyeSqCqeUXP/LvPicXb0MVfVk9LlN8s6L3RmkD6gpncKHAixzWzcqAD8yvk97sZiv3D7
RM+dXF/4YAYUW3lr7Tzf8qikGJvmziiVr6ozxrob4MQRbhshJt+xh6vEYNharD6MJYU43ZqADbDt
8dtcA5QWocTq4qR/PEEjKA0Vd7/H/BXKTLqmhvZR8DH6WiR+F6Mu/9rH+WAPsuhew6+1zbWbSYUC
uPJWhC+9kll30cUjf6alcT3GcQ/Q2tCxzaB5W+p0dTD+iE1SqGL2uB4tDR8C3rg+aieI3IQ8s9ci
OruzPQwFJroCXLl1nCZNvYLNb/xSqAoJ85wVEcCDd/pbkUt1TyLKuIG9lhndp9q9LoKvd4KVov3A
OZC21vb22fJnU9usji/Gz0qUmPVcxB6Fyj3Q0f2+n0YvaCwFExHu1W24UrJvwK1ojAnzETzNyB5j
2gshx3co0lrQMzwb23DrolgUe9rZ0pM0ASkoBgago1OCt5okm3VhqOn5NJkpudEJKUhHv2i+datC
Kab6OKij+I51L31h2G5Al3/c4xTVbdDMzXAhnOUwYI8V7S+XmNdZRXtXMtyOhIzx67WwRpsfkVa+
Zg80nstqWzhdVSs6XAaorA8WYjSrBeYGrg4qCXE4cg63LUEXvjGBogrdAcrb9Bp1GNNLu5iturk6
7LxEJVq5PcVPLoApoJM83g+fVrD7dscr9uZzbAjG4vZMwolGNhjICnNSuefPKrYELwBHabLnkDiX
JGX8mSthWWX/yd59ymBTfzT6vf3e0zZnMqJDmc1TuXgwHSdhbECAD4MVcWY2rC3iWuPQlTq79YmT
PNnM2aYVLZ84+1LOE022MifMX992NvCQUUBDxxwXj2ovgNmvfVAwXie3Qz97gaGGntNgjdRAbre7
9XWA/FtyeIKrANafiSwbbwKkO5LpoSyG/0ywXQUe2JDcXboFBKNSPHl1S9BUJ3oUXq3WZTT70+Am
FC1V5tRp+eMdIqAGsn/5LKdYhwNeuoXFnUXbzekIVKS3QcGYl/aS4ikCx+MqIm97PmQYMSBpXAGj
EMgaBKqkVB10bDZdMWier0KWo8747ZGCevATevyIwm8+XUCYvCEUK/+3ZwEBVuA3PnetjaD+PfRJ
aNrgP1AK92Ve9T1oMMZi7Z2rTlHccdlkYPP8e+qMHRk0ifPO8QViwm/ELZ1EZhz99N3E/SJyK8XL
HgyN+NceJtNcIt4qwnCEcV7L7+nITvUrDBbKBpX/qUeO5wGAaeFx4rZqY6lMlixfvv7viecYDXMd
XUuQX95WIPIKoTyyvVk9iATCuCu++R9HhUu4+rE1v1Xd65FXWuyeksgtyTsELq18ImqMYt1WllZG
8JVr8gNvFZBt4lXUGUjWO2m8h7Jl58Pb6JsqK6R9b8JfYhfcem3Opk61id1shub3t/pyfwmK6pEa
kwYpFU+sOc7J18Q5IMxG8Yo0CEvO94uKbBwHNWyPiGZuHUk7cLsl1NFSC9PJ9hIFdawmZrTF7Mut
BRcbLbw0L29CGWBXFZrdPs+fUbvBbG2jvZanOhhg8C7zwUI6WtDMTNUTmhRq+I7c4QQMcLE/NX6Z
JrEEmUJw6s+lMusXid94CSHbl2yMHPD/LuRjc7SNSeyBQT8y4Po1WWmK4I1hYnZstxAEA7qb8qFj
i8wLZQP8mLhFc4tldBNJyhFeJvfrshFZ9G8lo26qeM3TuQBOj/X9fHUfvld3Ag7Mcob4V7Qusy/K
U5HMclfMBoQ4G0Bau/XJFBedenuc6fJX6ZqnSjylBV9Y4/v3eCpRsyn/FqqctEgmL04pthzEGb2v
aWxYnX5+0Q99lE68r22z6Aj2Hzaqmer9nJfcP1wbo8WrlphmjBPYhTNfWdjNN5x9EHiomqR4Y5Gm
/crzWRqSgjLZJjfR7OGqbk2pSHAXoUBLejnpP8ZMCZusYaeMo5DGfzUonCy5OoDhythTxgKsMHOt
WGh9AF6JXV/l/T77uUljR1K6Zr22HITyUFDzL9Mj0QavInNB8e3f54epHP+8mel2sFzosaZOu+dJ
Cjis8/+KL+82wZKcGrHwVGyFZ2zAY8xj4fP78VXrnJVCGHjiFukH9xGfE4rueq7s5qqF+Lyc0lRS
kEYrelXXyRMbwC+W1XlFI1YMw0oewT//pBW9J+JSnhak6D1ZB3IEYFa0eU1W2OVqSFG73Mw9T+SS
sKTm5E4H4Ok6Bwyb2QD7zYUdooO8sHKJqZzl+JzbKLSPIriXZmzfAvFlBUpPWzqID0zukTYlL723
BXtyv+hkVrmFIv5nHarUhDTEAVPz32ADSO46qWxjB+GnPO7kci7fXLmKVzbNiY1DRqKluM8HQ1Bj
cQatGCnLSfNMOtvxN1cHdOmMDGcYBwWkKvy/mHXjh7jM9lAM2n4lK85J3fVQv0T+WX+2NtMJRx2h
72g65EAyw8f9towJjUCRP8bEEYUm7NZlDnF0mg7Mm/6zNuJ5VUGCMqMSVifi5QLVYE/ArvSWODaC
9VdLDTbrvEtoR5fa9jPTlSEupaY0M8f5SsFLJcbhORzQb4UDtaDkhucNKI+uRQm6uPNfKUMFxZLC
1iq4eBLD1eB+whlJ6mNfvpr6UV0J3JM9H6BlWPxZKLCIrk9fdzIIEytHrjxLyZADfzhDMNzTUKHB
BvIjIjKcOqxGBe8eb18Pt6soq27wDjCqBbprM2AvYsgYWh0pWJAyolU9TqOtPBdznJgofsRz/DG4
XqlI0/zcsBaCOtylCjHO1EpHBo3Bg/19UPv1QUaN/zHcCzLd81DekEbvsXUNcqOKElnKjHvrxPzE
ZogPm4Iiv9E+nZatMAZK6c+MoZKAD5FVolCZSRwW30F516hN1hugl9W1ADcWrfoUhMPM9sj8XEvW
XpBmuftW2sFrWY824xyelWc3r3wIaeh2Bst0vA9rJUH5/h1F03lNKZ/W+6svem9CLx8p3HY3gMGA
7JNK8Ue791b77VzXdTfZyool8voa7F+BCwK4aXUcW4qgwLBpUt0yzY2lmE/kQalHvBIAQXmuvTh5
xxlI0JzrMNyNVF2PBs9q9ccZC/s2ct3AtGgXz1R7E3vlQMnlmvMkahviSgghzgKFRYFBnGpV7dbd
eHDMB8dNFAUowPqAa0L3ASiUgbZ3yVHx/umlI3P/w0CrFY3cz9Q3XghKKvKw2TkFYZvrdsS394Dr
Y9wAlg5mAG6FElgUWQiOASeTRgMr1qFZjchDC3jbHKSWPESGVoc9a4Vl8x7Jmef54ym0HsLctlOC
fpbdIVW0uSWnBGgnjMW3x5gBS0prbSMYNH/SdOuRLC7LO2mGsvxQWoFSwV8/7cDyErDMxLmLx3O8
B3jKrsKoe5wTPQnxO/fLNTHmTmvvu+9mpFLpckK+fDsnhRXkgopXAuA3HmZZB+UoD1feQ0zDVIsD
yzdrkExRAyZb8alc8Mb4maua7tThQqsLWmyNkEKlojve9xUw+VobrPPTeRmvaguTyK/a0qI7ddtj
opA5BItcHluH6w7MeKePu9BT/RJSYRP3tYe+LexxJzXYMrWAdmOTUbpzBtdY5qXg7MSjJJvs/f4D
o31cxlI5nrtRGqnVQ1PDk8RsfncNMulg4R3jA2II4FnhSgnRyzQWuLS5uZmy4S6yDUbXxdS4Clrn
b/Lu9enYgVvLFDkz33BZzt7ZNMXjpfwWLreb+yMFttokqeImYjrHO5rSL/YWRG+1yWxkKgOjw/r0
x1Qf6Utf7NsNjHk/ILGqlYYXCpysIK41wpOoe+PVjhfvfhpIUAoMd0ksTZ+cFyOaXWp5KcNHrTCb
awp6E6bod6P4V0zsyXjAlMioV8L74Bxvun2460DJtmekRjS7OKPgZFKQzywpK4h8tvNreJCP6VZw
5BgZNQ2jPEJd2lkumiXyiZvjmh8Ss+y2xJlOldG8T2KEIAOfrLlgEWOPVM8NxMBeqvD9J6hNKzU0
CtDL6XrLJ9fQYuqDQQxbxCc1g8fU4XKHfZ30Gpunp2zjzM/xttkTOc8ZNtvfDRKNsS7aMwezMgpR
1MTPJsK4Wu7Ji5Xt2bLXkM/zelbSLwsMzOuEpfQ7p7nSixCsVBukNNQ3kjL0B5Fpci/KB9M2WqHF
xEZZUwUrUkkItFcJQLGL93QHHAAFxF16yt5v1ls+3tZDMS58VNF6sk4NxH1lc+qQee/MxxslICyg
JpvDl6ANetqp8saf4xBK1qivaxMOI4HQvcqUUC6QZXegHZ4HWq4dur5e35AM9PZNe42QPEubg++o
hXQDJfevZOiKgC0TLUHQWjW1TuC2OgAn2Ze0vUUloNTh04T3DyLb02LrQw4jSawlP+aNaNlKqaYx
Tpn3cz2cbLskAs/G8037/6lOXXvLnvdYGDunueNn/c9ltYhT2OrEB4skr276Ekh7ILsRSJLxBcn7
l9kqC2hiHm3+/GJUmLl+27WeI7K5gsmAOXat2BJy0vxAW4Z9EScpTm2t59f3CMqzFI3lCOov8u+g
cNpKA37p7MoeyeNr3FVb7UuoHFHeyBBtY3IDeLP0nYCNCueCv7sh/BCoLwpw5/5wTzo5TykvDPSo
UMsnkjmdHzMd+XR14SWGVpnppOiqfSsS9BcHHoW/OGhCJhdQUlxp89Rjnlhp2MOflxsvW+I0Ifs2
qWvPcVYBaEa60LN2HdkktPzrnYO7cb6c2YpDDiEqLyKrku/cPd9AYljjNyAdi4EYAJI9mDNFkhRJ
6w+P8mTf2ShMUFeRJ5tJtQ0fzJGkYObvp/G0VQK4G4AaqdiKQLJweTgPjaBX1NMD9H9sDWbnrJIf
31s2/b3om9mxIm82MvPwZAEsS0UoyO/VZPKDsvmKm6EJ89W1aEljvI7HdrdFIQKMJVw/Jm4zCDsh
AqW+SWHfN9mgsHLavSLoMa0AkL+1oPhPobJcmUe6LPIk0lZxPDHRS+cjILPqEXb/CiYAhtCqQaBk
/sK86MjvKdaG+aD370W1WHr9slIPlKBeJVeezwOHE1SSSFsmB02HZGShDEddUhfKAGmXpGFgdpJY
UymwoG4zt2P7aNeusjOymf2hSBmp46Fcm3Vjal4oOWxipozu1M/uTUJck/ND7/l8QJF7klpInJ1s
gavHvkoNV4nMC9647+Pfo309/TdUllle/5r4pq7z2Jy/bawypxCr7yUlWOl3ww1ZjMHxyDb2t9oe
o0A6zGf2IZ/TzMjFRcDp/PBxb3Mz6mfBUiN1hcAWT5/ZIP6wuBAnOyBNc6JNVD0fv3rw06cnxsjw
tC6aepWvsXBeFV4G8DmvLP/Kzcojt1LnqPm+7yPbQtXbyJpSU+G28OEo4D6mLhBiGh7SVv+w2rp5
CK9ColSZJNnA+7OPtiRTsjEKevQZyKjqZELqa0C+z15ZwEyG+L8zt9ud8ezqFkFp5QqNRT1SVQKd
L/LUlSTLZ6pfi6JqmEHz20Su/gNUfryTAquyZZNrmEqC8FUV2XuMNYlGR99+dPnT24/1OEnN+c53
x8l1qZ9DWLLE3yn+y/XMPbISxfMLIwqywuCBm+6kSkLg+RhDs1s9PspalORM5fTZdXV1WoqWXy9v
4v2Zb9/gioN2yIG8+X7SnF942HzfZJuGaIjK3iKI/IlB9yNB++fdjS+Qd6BkXYVGix6h4lrZ5/j2
JbdOEHz/gy6WxWZ8dMXwjUTN4oTxOPo4VP+OyC1ezMDqER+0QD9JKUHdAeA/Vk9hOd60dK2GNuHw
B3A3fZyVvpYufWXxdg5MwgjjkM84YPABfBoNg7irYNnf7HsOD4vqyyJn8PBXBzweDCdUFdr6XqqM
vTaaBxFuS+/17UNmPGxEfN7vGOpggtCrOefdXZzVy1WTKIA0rqb+mFu9tt07trczvQRNF+Q2/gGy
PbkxE5hVJIpigKRzaHgK00IwmtXZ3cQaQs937LkTE74fwePhM7768ySTF1z0AvYPm0jbWRi6/rMp
vI3Ms9XP4EwLPJC2FB+YyjLSp8NzBDUxHv0m3eXh67qdqRkQqzkhN9tukwLrwVv+0sHoParEajGA
v9nfgEYCTyPu2FSqeTioBxmIWEakHwhJYiKK+D+zwMnONuBpNxtefJKvk5jUT0LR2f6vgO2LPgUo
ji0CtiIv6+wN5+p/I+lSZBKXOUpHRW2mHz88/YwXtcJPnGY4qMb0PskMQtg2cUUySAbsXLnzYtd7
LdhgigzlIJKwe9/LxX/7NpiqR2WSJLZgm6yFI+2A4qeMlWbkF4WU0ng4CoJJr17c+wdjOsPhYZZc
DsXqCASdOJ78ibkNkQ4J9faKGyhxPR1/HisdA229KTSWeU4AnF9w+SfbqqiyDqq7xYkNs95Devyw
YEt+r4Zmi5+6xNiiGdnbgVLzYn3tZiwR72YcDvs0/lbMVz9PPYqozkwveYbt3gyP6YjIPPILYIwb
m0mBhNUL7mpe38YmAFzP2XzTNMNfMQ/PoojcJxQexQBRmL9Pj7zCN211ROIBBZJc3iYRj/zz4leC
1H+dpwTtM+gEBhRq7Rw85jrUTR3cmUkC0/l3Os+1FtRRyU9VDwfxD0Hwmgo1I37LsV2/xZVnKVV+
KqePToanbziUB71zcCiUKXit5IsZKdlQHPz8qwW47qy7l91yf7O+pnHNGxQDnuz85c2j+1MXkdiy
tBvTHY6KBymaGYJaPg1rnfvW0aWar7wuYFU77ykwR8u/Vc/td/4FjlJJLvF6/tyDYhIwE3VW2Z42
HUkEtVRTiHW4zfbDWo3DZHE2oloirkaNMw5JW1p4euDClNHYFgRaDqJbO5mMFOx8xn9UHBR8jsDB
8Rix/Sc7Gv62ZNJEscbJtl9gT2X+oGY1fNEB21RKPKLX3LFRlOh96pYgntcZ65rGBH12GRhV6lTb
A2mFPhsi2zoOpDeCHwqt85vz3P8gEkdiEb0O97lHKXTOPr7P3fXvKlALJQV4kUX6U7Iqau5K/GIg
22yu4RewST+b4kAUUpBZPESdELiEWDVDDATsGdbDWAfC+b2hPID5UJfYTPrOhUpwlRM7Xzrp/0md
6srD2/vPx23ct6Oq3yGHABsOmuJ208Jsk7FwGIGG6Ie77dD6m2tLgC6UKWrCeCJJcNwK4Sgazk8r
Cari05DHSY0Nyo6HKnBOF+5xbfG90heOY2b5Rb90e/ScPR+4rVofBLAseuB0WB2/sjZjfsIUbYW2
OvVCXgo3u7QXzsTM4//VtJMojLvUpppjZSgNx6KaGMYdGxV5f0Epliyyzg6sc4MJXuYhffSYqMFE
MboUC8JlN+Vp4OWn+aBzzJeLxaRjzdl8zC/l8zt8itZZPIdin7f6WRTC5Vs+RHt3613d5+egPlWJ
NXdH8XCYYOIfhAOq6q3r1bldWDo5wwCFdanAHJ2u8i6WVKOawIJVegMqND3kBBWdS+7Q7LvYchDk
4vHjRMIIYfyK6dfEP5Ae1hViZJxiRIztlj7SfbA5vtItydSsjBIMDu25D1H/3QjU7mS+LyyuwX4z
d/4k0oKvi7uGG+Qt639N4F+7lRN8OEM1az0DeROlmLx2wroDqGjzwRiO0erRtThYLCIYv+mvnaTo
bDpkjIJrKubmWO+kArpjCmodTZCu5aG2RP2f6ivrRExxRPL3y6DO/M4L+GG5rRGMDk+uKHHJMH0N
oJfokbNdOuorejTijz3HkDNqn2s/eTS+KkjeqmdjXWCgmP5CZF0jhHKYjhMDHHPYmTpjluQHDRx7
Mb0e8EFeVOMx300Bm0iBJPhP51GN6Qx75hClX2nGfPn3ewc+ib4d+MzDH04LLep0KpbiZU5oe/2C
RBmBFPIlK6Cm+2GpuorrqL+2Xzu7hDqgTJeN+U/UbtRbx4E4ylQO/ZH1Z1PiWn1U99BBkvFgqrkd
fKvKN/SB78OY2Jgz/4/pMyw7IhFgpioiMlXdO1iMKDuAwjHKlSwW0cjOzmqO5cQduITgdscb8SOG
LRNIUFjKtQ/DAvFU+8aTtAP5eXi6fanVBmae9/nqMV4KmN7oPRUIWgLqzT+CRjd0QgJhibZ3ohqb
c7BJ0xj6NxJF4TqhU93Hpj4z4ZlCJChrNfaFQpmJE9QWdt6it4JrAatnbpsQky7/fxSoZGduQl2J
Gqatb8opr2TvV/kN7gUC8juGFCwUdmpSwqjRi3w0dEGQfvY4N7pgs/ZFz63vIzwqpm9ig8+a301f
KQnoFHf+PXk3yZ0yl82Qq/rgwggvsQhJ5O1JrNJ/rqlJ4/C1OuLP7i5oo0zDOToeEUT5OQaTAEv0
yaEsF5LNQBksHGyVC7Wl1wVAJeITZaVLeJDhD3nd3Yx7zWqBiy1rzkmFFQKvQfTfczvLyzi27Y9V
lvgqLEq8sPzdBsYKkDbX7+CrRkAbdv8POIORHystttclTlBaNoui+p3MDw35MWJWCJ23gZ41KBZC
rDTh3GW3i75ZjKoPdPA2UQLdH2SYdcQqFy8UxlD0m31znWc4f+j5r2e9H8mvSg0sXQy5tl9TWsB0
ijDqFueruPcaWEhpJSgNOb4i/fG4Hfnrgb13+n3DW5djX9lVKeid1CgHoyzffQ0fcWN2CQ5Arkzm
FDPMgul6AMVqQRXUHsLS4bRBQBYhP5sxtGJvUbZbHqVqm0hClwrZKb7wEzF8LkE4qq/AZ/Ca1ayz
UlJkx22j/0IT6SEY9gXiLzoWd8AM2IgEAgF+fxoolcli7ve1T4bJNeBmFvx98FiBNQMbQgcmIJ3Z
YeAMZZwexYbIl4VG/J4+U96tXUIZMdvTzZX5I6lYGuHHtr3MLHpGV4C/aMlbAvwJlwTkd4KH5qDU
1eYRDWs6vp8nl3A1Q0AelV+oKV7r7eiPZZAB418r4uoY1QnQRDj8BRyvOQkWyXjTrx6Jvcbd1jnb
/8DqvZAf9n13hOoiCLFWbwp+vkYmIyZPS8bAAozpFrsyK8EQ1QjSo4J8+u6GZoespB4yFl6anU1H
PUXbAeT+npsvNujDWdyOW+zbArLxpv4MvSYBS+8C4C1a5Wp2JuYHEUwnU8ujO9wI9/i1wjOhvcN8
yqEeJIbc/NZFw9JUSHBAOWmlPWWBnMJrZ6KxEQSSbxk1XQLwzdEA6psQx7rZ01zKIaU5hf2dkp+1
rSCAbzR9sXfqUV4GyIKtzNeiwj9pNHqqaEgI8oGXaw982HnYPRpzo6V0EmzLfV8Wo/tZH2OHsdWy
Szzl4IgqOOyrh0tb6bo9U5CNcm/ppwAKI+wLfiMtXZIjTd4n5kzaCyYCS6SFl69MB/Bk9bWoO3p1
L3kShbsgo3n3kZ+K5zLbdQJj06vBA8u+7gbnKgNlMwK82hci6TTshRpBYtUgMF/wb1GvoCBb0Hdw
A7jvXtS790GBNbXriqMs5HpygyMwLEBWCTm1jrghTF+cTPLIX1LSY/ziSy58RAzac80kEM2eTZI6
cXdHDeq1HqDLjigMmMG7XyoeX8/z2GNtQ2WkDDXjWDU83I9/J9f7Xuk/Lh0FI08cBxWV2Unc4Nii
ZH8v4LBO+Qsht4fsEamHWwvjLpGpUd2tbD9drVSykRyBxINfkSwG4n9YlgPeJ3DK6KySsEk4ugyi
9N81epmWjWXhPApJt/9DUsXM9xSAQ0p6dr1MMy3H3SZneHymln2s7N8zQTuemVNsTj9XWoB2Orni
WhIdGioMOeHQrio9iBss4AdbWjSbsrKyp893QfMgm8FexyCgSlXmO1KlEjA/eECOE+DPWCG2Lq3i
efs+pDFLsEqQTw2wOz6yTh9GQSjOr8jBydPk7qr58nAvEt6KmtIx8TasVYQ1Yejich1PTzmbK2cy
1p41LHxUJYhyzobDGINOe/ZhfwMsXJGa9LeVC6gsYSS3aXVWjjS4n9ZMO54c6kozIWv1+uiYNc6W
GLcjG/CnEY2tSNn9BpxGa3cjMmgjx6jMoxkCT/Eoo4ClirHyj8wJmm3KSvvUuhoRTkHwvY0VflGw
KUgZMAmv+bUHnx9aqNwGXXHPs6hDrvRX8qaaX3U5MjWE/6CFEMO+K9Y5teLQtIcVjfATpGZlqtKm
mP1A4dKBtaWMHSuV634xKZNADgLqBKFyzUgcXSTI5r1Yr7jMOoxDUE9vXbHMt+Bu7dYfSfMxDBYZ
/Qjo+qlwVnENdJsTOKE9Av4oLtJpB+CJg19NOt5VqzAcodfs9Kk5ozGP4MGklaZOIC0W+KPLhp+Y
MHvJqUg+HQmPIP+9qkaErOVEreJmSUtFx9UOndyV84TnsDTwwawGy8k2m4tzBA/mChYk7x8Yh+Pl
ZYe8PgOJ8OAJ8IR4H1nGUzzJtOOzBSERt3M7eMq4CNQsxReTHjGQAW8yy1o9ZPttdIcBalRXPHOY
ALrUlaYr0tRKaIXgCNQoidjmXNgKU5T17o0qcwGTa3SYzbxsKE9/mhF0Xu7cZr6PB9+d4LULm4EC
sj5ZAh4Yz6/aUoAUEDK173Z8PiE1GMHpujuD1OL9khttH/4C17ED7VrwLZwAdlp4Z6wuSzBPqOWo
Dc+6nUqgelrIJ4u3+25WCLQcRi01c8D9MOiiGnhdGfxOkuYu4DUn2sP4BA3oFjFS2dh3JKdXCFuH
jpZgrr0I0ufiZcN0DamUgBl+V1kcqyofXG+WddLO5+NJ5Qdj5zlTt4uMraoXoDAappeKSpV6mW9N
2RRj5FeOnqaNlWGnUCLUqZn8ezXi9tb5SL+huQLEQLGioFQyly9/7GOt1qJMOa+c/fviL0yp6tQS
H5tSeXOq+8hyNIdLG1z8lOor7R4/XXoCKeXdVLo8jkVINxF/yHjqSEb2SpiZURreoxi6FVCKAbXd
OzCeaCjrr67qvFU15WEiFT75BAsXWpNUafau1KrLNLT3Fe57EvL1mDATB6MH6RYZR9pgZ+XRE0Ku
pcQRu56jwnEG+YvixfODHwkJy3iio5kVgML1jS9ImQu3Y4BNHcNfkVJ9sZlmsbX02zYeAIdEefVV
IHwODDD9rwTP3y8/ZUj2sNZ8z+RmcbKoyo0a4RxFrUlpMvC52Xb/ax5cWxrboJ5men9gb/I00UpR
ea2lhDBDUK6zVlotswyFbqBKaSttwyJ2G8iHz7EkPxGPCr1cw8VXnz7EszfXCS0uZlbsxUro9Gon
QYRUiSx8zQEuOAjpKxtZm3WcVdereUBtF+At7AvG7+T1szwFM8+oSdT65R8tNAPMHZjN0l/8W1sJ
yyj2RPCm/O+bbjRE24Eo8yF/PttBhFq1l4wSE9j9EDPGy5cTHS89oFi6RXJTArGFf02vLcP8D3U0
9Unl0DUI9CAj5xQSSzfJ648oT7QQG0+v22wfQRpFqQF4JvL/GWCViTxEwEGXNkxZQW1Gmk+8LjG+
PMiRo7F2OoQeBQCG9b1Cm9E9n50eoLKnP9VLM/yBk7bcIX5zJeBuWcRCy/psczAYBfQspFxkVxfm
mVTyP3dWpZeu0xtpEgw7pqDYZap1h2LcUUnAOVgGojdW2cnnzrkLEl19ZHegzuqJ6NzkRoIJbuk7
TmZnEfvJaOvPYvQO4aK7ADgkF79/FGNTYkXCAgYWwGxY8ovqxVxaNCMvjI8ejY0S/ucOqcNwj/vr
7pW1S0IfXnB9qP7UJqzGCRuLC8zP4zemZ1bY4+FBeSYByxEdppbufLzsVzOpykcNNyeVxxHw/IVp
GsIYDRqFB3HpPWbsU8hq6JdxDwFIkJm4H/ldJmrBy4/R5QPJH5ZM+y00ookywgpEZtrJBwCWBXvE
QUUIPo2UDVc6zvJ4OZjDJXPf44jt0SBLHonbEww6RxuoxCoBw8+QYprx3Bxo77K56OrCbXwnhkOR
KkLJVvvHFYoNVkQDmXpHMdeOjMEX1SCgEiiKSWHjxDb7i+Ue+NIs//DqmYHY+4MQsBnYjP05kQ4q
agSjr8v5oJM5uisD9Ag3zzp1omKeDBBhSsKuKSkmmCOSJMdTl16/HZpcW9TO8wsmTXYiOpXEjpVx
eGQHxlIDqDLKIB/QyUXS5DAtJa43bUtoW3DUjHr1iS4cZPweg9WFkiK6X1RSdTKO+t4nZRvoRkXB
rI8cIX/jtUYP42i4zt7wks+XwUeH7GQZJU2pgzUbCgMyk4vuWHMblgIeJQzYTN3b7ps72lR/A8e4
5xvMmO8IWdA9WMP+sYpuqoqhCp6KWur3Tpwmr9Q0QwatsDGlP3l7o/7bavPFnACgXuWfHBXy7gSw
JIxCZyiKy50IjWCQrvoilGZDLeT1iTGCFQNnvA4Ka2ISn3+DO4D5fEb1JrPlr8O44VrbfsG5CQoc
NGq1A9C2i2m6vbWlQB/uVwF245WM4nmUWxxnTa6SvB2PtUcV1Laq0qcqpv02XupQf9Z2eOXGUHbL
Nqu7drYDV8nYvH/70SlNvSptFOuGeS8sSxAqK8KAg8tMN3eLfjhTF1JgUM0Y0p2yOUbgHBxLUr8v
q1XfrQqIbcMG3umY2IgQ3mv31HREmOsgNox4lw5FLciZAgIqz0Sacy4GwwE31vomKwl7kG5sf1ox
XPLKJQpTTmidZVOsKV0Ewb86irwSwTR3ryld4WS30gw7ud7kfyEhq6lUrTCYgH3BhZOVD/l7BnrH
8r2JiD64zKPyvW+2+OG376BbnS7BaSbJhOZC3TrAQaLvK9F3m/W7yvMwpBHlGtQkqWlhJPNmNFQo
XUic1iSI7jEkoXg5VQZbq3SdfCVmpHh/G7TreUecRMpRRGoxoG1RlJEP/Rs9+zyNtRrn1lsdUkzg
cbN114OLI5NbLB6T36qqlcAO1LMlEpD7WqvbBuRw+Pro3JU0XQO9iYIR84RQernSD/BfGBKMVSBB
wAy/qNsb0pBTm0RUVWRPNMMgXrRgonbqG6LV3QlxIa9Jz+1PfzHOjEXzXA3wthxQ8OGPI3XQNTBq
t2mbOlMcgTuRL1O7sDF2yxARhT8XaY7h49/5ZMniQOsCsLymxnl6RLw/Xf2n125Pxy00buwHRMcE
HDUJK6R49aQOYWNOkOZA8TnbeaTklkgB+tQ191SlgXduuCJr7LdRkJR8JcJXfbuUqVtnEpfsezZ5
mc6vm5tvtKJ1hQg7qtkRNge5jF4sMXXCwHa0gODpK2QxhwmQkaaipk5V9D3YeE0sSVW/44r3okIz
KeFhadWT3jR+6YkYYuXSb4mE53ucuFUxy+M01iXI0pMm2omscQqY7nLBKABj+waC6Y/8jkKTsnVL
KW98GzWiqUOH1vPcEN5TSM4N2At6OcLCNRw65X82fQ3FjFkfLWK8KefGQ6u6D/gJpFr6+0azCd4e
8ZPvbpuyYbEfN+cYCS1MxmZ8uGV5OBf5BL2p7ArevEBO7VVpzFKIn7niRsKCx2eK1KBydbLgakj1
wg4oU7jvmN9UVt1UnI0HiJQJuPxfBax4mTi2nm60MOmNNaJp6SAZhQv4H7szefYHoq2pbrJwy918
FZvr/fX4tKRqf8AAXQmFyOlaK96YasHK4ZWxe0e2AZhsoYTfPMuYPAZ2ws+lEAA+3K3rk6dU+iTy
qP+G2knACz2SXG83N0FHtG7zsHlPD9zGkEkMM+Calj2eadfgnnjqOj68QhhDB2vaxn+Yf/oCK4CS
Y1MmWMMP1ypQgyNr6PBR7GHftSvT7amQHcG+88P3fNEdhNSUoHXF74j0eaanNJn//TThWz5Rc+fo
LB+khTA+0yuet+PEhe51DlZm12lf/bvhGDHRDrnvaPX3YnrXlGVspZiutQIFjov+uE2X9sLtQtrT
ApOxRzW4JTQZroV6JW4zfaMoURZ3JLwgi9CRyWHPJsJtQaH9XHPVRMdv4LbSgt/c61Xk++0oifdV
oITV0kaLI8nUDvetdjD+6Lkeix4r5tBa0yIr2tvq9hGJIoPdcpuVBTQCkA5Lne5/4cVq/1uxf5O9
JNz6atM2hpw15Bada82SmrIXYCOniS7tUKd9b3eZU4OG7Pezpbu0JX/+Sz2IwNPlzVNidFsLRLJa
mnUQaejI+ofNFqlB4ZCk3ONOHsbdjCWar0gsFpFmQGR23QwmZYqjivUSz79sw0oX+KYvg6+K53kQ
sO+vYIIVn8ONySNt1xZHyW37WqAJKiRF8Sn8qVqh/lVY6GCmwbshptZIv48Hj8H4re7E9GnY8Ess
w4aQQDNaL3WNoWqmgBUkcWb05scZj5s5P79phpHKBVKwnIE0o0TZIC/uRZBj9/qdH6oIcrGxZZPl
4se5uEcUH0MaG9apetxHwElvgX9i8kryZ6x0CSnYo+QYVLFmhKxCe/92uo48BJdkCqJ7Hv+MihYo
dQglhUNi0NGgwx26vaf1SEpcV8g0yQHT+BM7ha3oQM/D2Mm2TzvXPFNZoPwbsx0aMW2nN5xu7GWH
Ucw9m70JcYiUIKrhCnUHiPMN1DY/W7w3vfobSV472qKLPylLZQsfKk6OKyrYLME2f2IE0bfVJ3lY
wL99zgyQOdvz6UVnI0FICJNs4JpUyKVgXbcMlzhRlyRQaPS7yBn3JlhcN0Ukix3tGCZ8UEMs9eAR
LmbptE/AeR/AV83gBm65RWHcxSrmg8zrvfSW5ynjySMq1Nnbtu3dOK2jv4Lwnd0X9yyMCwmIsiqm
jm7+d3pvNVBAoNjvK9dld4mwp8VD9Db3QdG4F4w/XT0kxodeS6q0YSACqP10nZ17KfabMfzTJfpu
yDGQCVs7eo6kkimbIkpAcBgViH8yzQ+b2b7xkcOBfHtsEOBAoHiT4uN4qhYMZEyAjzNgHfx3GsBu
lcGz8TMUWhJWkuOeEIEv5JKiR6sinI4lZIvMXAqFA84b/GVrp6h//LcyhuBdq9uKr2TTNBY8VVg/
ieAjBQEcW/HqFKciexNUJc2P3i+O6j+1t/lbwATUobpj3rNxZ2n9tlrHsjZl9Kxu44EZzgP7/hD3
kB83DmrTtenhsAnB0V8qsslJogFgXBhScz7P11kEIAaZlnBS/T1buebrAR2ksDQ6nN1IVNHRBHt0
cB5yDza8r+4Zypsqp8pkriiZdRgOxBD3Njp/tnkZ2rZroeC1IqZLDVzivYALCoBWmAhSABp6V5zW
2jDUxD65WDarJ1DVtQy/19N2KlMBkoFuKZz3E5ugiKoYvTfurUpxntOjTp2FBXjlV26pdj+iiPPn
grODGT7Sl6nC660gny882GRB9a8O2QjEs852bc/AxNgnZvlY1qCTS51/PkBo/q/DOuxAOVuvSqfB
+HegpcbbJKuYn1hozm4rvT2ucV4jaVowYvtwmHIULsyOnYMtrNX9nyeHOG6jkGm7VD9r2DWft3T9
6mq1lhURFWabKzrUlvAaOJlkuLvWO7FcYKpvJ3O2+2K3usmv8XZIqFwxIdvqo6TDMYrAcnPFrEXy
TmuTloXCw2DOKXjghM//rWvqH9BoW7EN/5mbo5cU1waIEhscdzaXvuVlp90RGeDxWdZBWfRedTFo
c84k+RuUO/qdsfz1Ii+XZ25BPPzDl/5nWdy7H6PUdRdrukRc8xTZ9wtolvghDIQAfYJ4riTAetgo
3ngVYjVSdDmECGEyrPd7nL5FsY8u7BNc7JWWR/CKhBtVZjIUqtCfK/i2vL0FLNKko7AREuSfljUS
8p4p8gMTcoTpn8IFADCBovSTYABuXg0Zx4kLyNbbREFZpRK2YXv24jy0KwOjGIFNXzjMa99PhVv5
C3qAJDNCOGPm7P4ICvsRHlKEyr+Z3kqL5Ia93dj7jQweh6fhtjtdKZyujpKcxKgQW8pxCxUDN8JR
39rowuts0bPzp0kWOlQ64zJbHel6/2ZcQ9RBuKi6BEbn5hXVi7u9/ILRUL8NILmvPEvZSPK6GLrD
Ak0d/6kk3uGb0yNhsPec9qQENp/0ihuCNerh9LfPqsZjcw+psGsE6TP/omv3HC1KOm8RO/ZbMqHr
vJsX4G05Keg4v10TKu2wnNAIN9PRFzhD/v3BeZ9nTQflFYxwU6Q5vqiRzFV37EkVB9+Bt+Qtomkk
Q6SMf2pTE4p6R8PLIuWRczqOnUy/KhkYJdHUgOOxEvW2uFLspKIc80TqfN7/i6IU0OruHOMQJtwC
YyL7HiyuoMEJI5ybfHsZgyQQYB9t2dFuloQurKXAUqiSGbNInHd4o1PvRIvNzapcIh9369zVPznW
+Zrcaogpx+D8YKEH+ZlicBiyO2xQ9iGyhmamgw1/CNTVROD0S4mXecLUgpgKB8z/+Gw9cVVnY7dx
hq19xb7zLYWou67GqKN+F0lSOa4YyZJMX44uD/DUSmNTK5o/navGqT/SJoob86Ul3OhaDDLYwvu7
JZuM3eUl69sbPYf40NdPioMTMLOkcgfnOFuiVI4KElFKn2NQJusC/1jcLrT5F+Fk1YlLKr11lk6A
Vs8VArZ4O6yE89hCnK43eqMmRSFlMu4TjKZd72odeLyPdGS6LrA31YwH5OpV/nb/Wdaia88W/eC9
PISzMtKQI4FdU/pF0mcFE9Fzc8J9Urmrcli1J4v6h2UdPxBNNabMn3ejvXuNYPTrPYjxMrB2oIPL
MNWJqzUNqHc9yTLUp1vtsVtmCRsQ0EvAxMq+m+KwI+PKX7BhlSiql/1WVWtZTykW0h+4WyAl+7LZ
J/fF/hkCayuVpMguiwWfJvuD3IHuHqmEC0uG+xx80mgy6UmnX3lGTkWFfnCiyOOAsaYVuQna2yV4
602qL43BA40hl+NWwDg1f5Nch5cbqTMPLtrY6BN7Li4qX35PY31vkSdP/ObGgXiv6PrF/6EtL3CX
ODMPEIjGPIeygiyMI+EsEa0PA0ODD2lVdlHRjHe8lgAm2fyGRM6gDce9MJgF8UYaHE8NKZFsCCEA
pRMWVCzdWkAt+ar5s3gp+DGInYc3N9+aE8arMSW+15rZdxu16aB1V0HzmGeY0STUPt9XdzLdVsqH
RONhxLMD0B2u9zKlLfklSwIT1mFvqDfMNW102spA+liWedhlcM+LRo9ndAyJSEXNz1DA4/BfbfLv
P1iGULM/64uEjkdNq0htrjMpycewCi2/FxvIT+TxKE+CCM5BsO8P2TXM2G+hMUIyBkggwdyMx0uy
yu3c14hYuxIC52ckHyyCvxlEDGNCFAIpKwnXBqiJI2PHkyKxq+J7xhFtsAvxV2tIJ41BYkMH+Z4I
clzgL7Hs0uCBtwqElvAEQPfEVbfsEf2RyTQM9U1qJaXW1gsbxCKHux/1cTmbIiUyTgDwhd0n2U1h
yaQJGrI7lDl8bYfG6Vx5sN4lnh8YrZZbbUOLBRYXax8CsbJWeWALlyTzAhonTIWkO0hWenIgWLDH
VQhtcWnNIkR/x4w4HhMwkeJRl9RjyQMytN7tFlds7gCrJRQSf+6F08qmcKtdX260CnhUA8g2xRt3
qrHPjwFBhlnwIuGi+yco0m2cl0MwlmlpBPee00wgrew4eqfNI4wyT8WjTALkNU/i3+FC6hxFnz/e
D/HWddcwokst6TPj3jFvXBdOa2ooErTqUjaVqRIK1AHpuDKBg61PyPC7x59mqLULsJofcSw4T6h5
xRh/YNS90j+irf8410f0/ULDH7n39MNSwTF4yN6WaO+5tMKQgLpFJC5l0mi+aFgWFrwnuCkoQgrx
18kZc/6SFt0ffSlnEk7z5cNjr/kKiISlK0GQBJz/OHpxu5kdw1Ww8gmkgzyE9gORLVLMRGqtnyYo
gcFEwqm3YV2ElAG/CW1jvpIdVnW7CEq4sc3VAmvrtTn+X7o9nxQNn7gUKeYd38dFTsRf2AmvQ4X/
TaLhTBNOIW4DE9i34qwAiRJwjXIzOYnlReV2hMCwyu0uidZtQzKkmAzqqf5ySX7p7g668vTEui/3
9CeClTwGtdNps/aZmqprMYt0HGviiObMPMiNdz7hyfs381UaT9UmbDhjjBfLL9YqUI5rGflOdlii
DIKs2Ij45MV7UYRNZLt/6gHkdS6ZuEONh6tBi5UkvXIwtIpJ0dDK9fyRxDccyNq/UUkLKGTg8Tfn
VUCZYvyZY7QnCKIMHzAnzn5c+0QjfJ7J+L83QSs2iTnqniX7yrRIr+chJeYzKe1zAC7G/nSUr0EP
L2J4hr3Q7UpviTyAAUjqd7Rjv88bDmpsiYLPmVGqafLQ890aY9AvHgrt5tSr9rIVHww811CoFKPt
9j+xxUxZBfvp+hsNsNZ+roZtFK1+xNeRaexg3Jak8UHpOHaGIGm/k2aIi+3pgh8Hh1AGPQmN6Hyy
fIzH9JDMU27DyTp6gcUrDGyHMm0AoOastM92GwudDVTDbiIN0+DV93LXTOcQVsV6Q1dzcmfYazqg
avJUVYCemiBvTz41ra0B0M8v27GplQXK6Pmqcqi1UZEb1BKeEtB1Lqd8SI6IzQDR4p7jFKrt6EJw
/PacswSZmh1jaPhaMVVeRmwq30sh36WdxFpsXv22AgYJlmZTHb+ECURsfbCrzCO2dickHkNuy3Ub
R9y4ZTsymR6hBh7RHBY6tEluPWirAKuBiqKVBdB2VJRF6ORrbJT5QdkjSUU0f2ULYsRtP6kK3L92
o8/3MGHvPfVHYoHDgwjqEgT/yPsF01y0Lr1MbIm0oYFOHDJ/SMAUy32jQWkz/VDcNHKRB58yVchK
z/IYthPkwwIHF7VIJiFuDDhkhcO8zeLbDOuUICY1KtOuAr8MhlW3cePqrG+ToSXVY4xGVNUm1udJ
kDd+Hl0fTwjBl7wh0LAUgYvQqdLsPPlb9SJMt9XbrHUFAMv1wxMpnFsDpLoZcKpnFpNMNDSPITYy
J3Eqxjnbk/95mU+I99eoPFcDXjd7sKyZ13bh+I8l0BtxNIKMD2so7JhNEbLUblV6DME7k7TCgXTZ
QQ/Ededo057YVaLZM8cLeudvA3kwQrCLuXuhV35lSkrz0GXYvwRovjBfakiz2eQ0DuN+FYvOE4pR
Au8EWgiFnIv7vqTwIFVLAZS+LutrL8a7RMouJWmwotZuxYWDeJlrwX46gUjPwBCnGyW7z3U2/Gxj
ZAR4ZQXYyTTYrTanKBco+dAh5VW7mrMkcukg6MskEEDFAoAghPmIviMMFq7t4FpLC4fYPldpSYx7
4Lkem4TFjw2khbNGkOrJskxUvOVWgTpyiH8fI9pIhp8Ww2WYupkwqDHGVtmhbtsxDcY3jvBTsvm7
U55g570PiTl4sxiGwqkV1z1vJgbY6rZjgX0YvA7ozSyzaF3DPDbRTShfpakZZqYep4fGv12zYKUC
rXQUPVosCZ4kb6bGDulyN9sOuzQcoDYcNe4v9ybTU8ryuWf5iRSJi2SJa00WHAw4B9AfXccR7d1/
BbKiLlbK0LfRsFBEnIcGcRdcKthpCrrkVX9rPKG9u6fd5KTqc2yWhepempY15X1k1R/gUDK/fURM
bfmYH/hgdk/jl+agXjld3fhCpqPoJtP94eWxbNSSHPwZTHtU7E0HcvUvjHK7n1cp56g2BxvAtrS0
Fbgm5KHBqLpfGId1N1aO0CZSDAi52HcJa/52McMOsT+1i6SjYt/g3oxttlA1501InCH+klYTEZWH
a8mflaHTd+rdHlwp6KKmLtLRGNugXnpc207uk3dbAVxg6P3s076FGRgWMHWp0khv98cFxU3KB6RW
t1JR6KRqbFyAq2lXxB7VJJh/WWVtNvYA15u3yY9+dNGSxGxYw9ck3f/xiWYOoBGBzMomqFF4v8FX
oM9hHPQ/YmfFQ3KS4LRO1Uc1KXYBTB6ZH4QHDXK9TPpyZzHlhiQ/yDAT/UYTiPk8ctW0AHX0iRWt
tTfDWBnQOASO5c3PyIkrfSYmDuFyOl819hbzWxN48v5OVdGgShoXbBb52rHeQ2nE7toBl/RGUDfR
/zJIjRTUNSJ3wtBCzGOWM5+OrNAKsF7ssznrshK9qD7x+5x5+VB+gQtqTzryHsmAolOuS2gaLJCB
Z0japRJw4X+xv3NePvQRQfnmIptNSg871x8m8kDmUqMo2CDy9wuZoC8KtQnTeiLryaXxjKACA0Lk
THAHqmz3b12YQCDzcx1wCrnj7RxrYLj1akvSW6/kRBQG4HSCafkqHZcJVnRIINWOgzA0BL7hJQ00
YL6D2NdVpwE8i22CpNo7tzLULLt4EdMKN59utfUGWc2qmk/JXXWUZYhvHItmhWtcmoC92XHqvwax
xzpkY3rKoB1jyt7Vx0aiFG5f+DKvLjRnsPIN232hk7b4Xm+wYVv/HjsWfuHS29EEomoZ/3xPsWOr
/7Y6eHA7qqO+EcFBtJToTdcqdWUXYwa2Luz6++bEIk459l0gHfWzLUzRCVioZalnppS8gkqDAvhX
Qp7P3BEzaKODRi2DaUYp751OOoA3G38H6w6Ka7w/c2/AU7BPIGPUShj9coyYlEsw7HYJpeY9Dm6f
44ULwi/6fhdPDiZJuIa3M5mJMOt7Aba8rDs6TASH+tJnN/WNY2EhYj+7Ek/ABYRKOExncZjMHxeT
UMDq9P4hhvUVaz3UvOj4q0ap9pKQqjSJiReOGyNqoOm2JRPXX2Tg1QnmOOezfACcvVYljF0YrrmJ
lZFG9dW8lEc7K8Ntl6waP6LHRmLhVJ0XbSPp5PDmjZAY0NhaGqGquErCf6jB339CEIqs8H+abqH+
h+V8NA7lzKuFShad/6vGbLr/OxN59Z0tTOqK7AQIqV/ze52p7WMF6xpJ0bu8pxniC0ADpTL+2DQs
qP0rxONaUTFGr96KloyC6eeA7GsAhlrk4Mr2cKXWhkeevtwiLv0Z+OhZMct1cPZ4unxGp5dP9WGF
JlFdZ6Q2nmtmznNlDHD9asjYBjih8rmRRoHWZCyTLuVna+8iB5U/F+/9rL0y9mThN/kV44IY0wVR
nrtPlG7jt+ScimYGxs8id4Tq+lxYECra/TuuBOg4QLLeR3vhO7LN/UBUBXY+kmyT6xNfq1RSH/aE
jvS25WsTFf0YwM3K3epE2BUKuRriM2vbwQFAKHEaWsmSl9xh8O2kofj0BLQfv4OWlxHcVFuSOiUR
tNn3hSo5OCg2Q2jFu8dpk3HglTZY/n9C+7naozRvECpuhcOMDzZq5qq+ReQ+iqBN6rVX8jVjiuj4
2CKWfsepjiUp38VKOQfYhMStnr2FBL1URe+DsBlRo48wjnlaHQ/T7zGxTBPR88xGmTAnLPOupQiL
F0F4+zON2ynEhbrnf28VUhx6a6OF9Qxx6+AJf0qqcle72GTBEflhIstgipl91nZDRROHQRijh2Fd
h3Vdvcujrzbr948DjYPsbDieS8w14D5+AxZ6350OcPZGHd5mHTjfI+u/U67QnfKZkf5A1eqC+L3W
cXQ49WKHCxfdLwIcBKvCnbeWCgs/Jtsvu/nwsBFkk51OuAcADMCtX2+UQnUNhxhtoETItLkHBAun
vwlLIMIaIPD4b8gRhblf2IRJZa3TnIb3XlwgQYbgbjT112EOTrTqHmtnHbSBA7Fe8yrrot1/Fo3H
4WygZ5gY1oLfPI+5sJr5yWlSOJMJ2+gW9e4xTYFTEfDh9gr+AbygHsoTb6twtlqZsLFulhNIcND8
L2yN0gytX1W+vTo3AW99PxPpxD7KzTixHk+zM1tYNFmRcIYnY3qxowjwB+1LPBZLrNpBRThwPpaF
6SQZDGK0ZhkoSE9vxMzyrLTPu2Fw5WM5fYvxILLUFsl+/911PA2p7a3XPOsDBYZjLm0Jc6QQlfUk
/s5mv5RP3mMDhRgVnAmzoD1GwduVRvB6UBetrmc8OeDrIXGZ61ESVcIGMaMyIq3F7uIMH+KqXHmd
rdntPVaYdyHzebADxorkxMVFaSNrPTFG+RsT+Gkf+b7OSIe14ky6XPOuk28OOBpDMqNFK13JiOn0
jNSWD6F50gigt214RU1Lr77OiEX4l0RctL3Pt8hZGQAKvb6QEsey3dpMSuPMzfdg1zclpl9CqikI
Esxu+kkkoUE9QscN0lOQxyR+m9OoLz14jmPkx3F5cfzv3YzzZnqEjIfgz6hJljWrCaJM/zAFLhTH
v3e3BUH/e2aKubUaprOoM5LaerE8enNa1ae1+ZuyqjbQcnbnbHEIvEcvjsBqy61nK73AHAxykv5I
kcnzL6UKp3WNhp6TcfF461ISDFX1JcEhu/mXHOAoxSlCprmwv/boRyxipVCmDMTXw+puKx65Uzs4
6ATmj2vd0tlNd7ZEVtlsAiTUqMCz2eU0rRsoAcNXICgAh8H2MXocxOXLAPc9G5z4d3NlNvtovMq3
/kNytOnly/+m8v+5XsZ7mWGJBRqHTQlnGiduUYfXZN692P2DyUuWIl8S3fqA8X6RLfwRzuJraQ0l
vAWPHIead/3r21IaIZgjB2nNUSfKoPe+cnAgmtdKEo2hnQuGbOvX/v3lAvnn/1JDN9i0wP6FNc2r
Ru+JR0ysfhB/qLX6cDuWJmK8yNcA71FqJ7b+X/UMlxhfGumWSePBLEtUKMC+LgLRpe8GyRz31kPG
7EP3n4brO+QIFUD43VSEY2YKOtVD4/dxOsLiSxhfk4gtJ/h/7xpUOo+qruxqQeK5o/CvVTxxT/rH
9W7oZy9qPt9v9L254qeoXm+ELwEVtw1s7aPuOVcjsTn4lBIvWFmne2DCn048lntfnI3oCUN93fIB
OjUhPUUqzOuNRefz/axZab5/fJBtqTvCT2XKhXlv6KaOpsy2+ryGbElhOrhq5JffyteN4VgxJvDB
/Uui8ctPtjOKVo3K7wJoR3Zw6twDJHRh+2Y0q3zpz0aPpfS7neJo2ewwHneZIZ7tsDp826KMzEPd
R0kUaYWLxRS4GL/LVXlBPIrVEphcOZmKFR3OKQ/oikbtBSeIbrQgjDQhuiVf79ns/Hu8666sD0YE
lOuapY94HbK4w5uB26vbrNnjxFYQPy45bXN8+dPLVBSGRA/lSbYIuBIpD1onSW3KQtvC7V8j5sBg
uLHd9ENEw5FYa/xnPquJ551/S6ud2qshl/WSTlJmdD8JoxiGRye9o5WePH2Vn7mj+eiBl/OR8XBf
6nAHRsqpXs4rX3b/JeoEwUIxOth3BVcG8BLtajEb7lXb4/TrfSHe6Xm4jUNe2Hv7FwkToCn/j+mi
XVa0ba18RoWkAyJai7CFnJciCNblOcxrT5N4HU0Xgj4LM1WQ2p+GqTAirSuFyXlQzqoO75/eDDqP
JNfVtrJCS82aPeNqJY5LTHLNSkLNvwGoft6QXHhioc3qmAThACAXTJ5lWxFQDNQJyrsA0VuOsV95
LfTcLPO70RJgDT2alq8f4nUAESW+rfECbOKuQ1aWEx5zw+gIN9XXQdzFQL8wf0ioC35rvoEH7sZU
UHybWzIucZkP9wL/jVLNmVwerubAYXT7/Qg3PFn8E9lZamb+SkY/2rJizX63H4I0JNyXTzeVwxrO
TlSm+Qd1x/BxZW+kYjnIp4FhPmFF8q0dNsgIJuvj2PLMNvebMRb1/Rn3hmuNsgeUzZ7S5OtNb2Xj
kDEQzRbMLLk9OHw5f0hgVBBrrFWq/csKYAtgtZzLUUceVlsBwQ7ky9I5TnPMyvsxZd9FvPgH4L5K
l8nnt+ITBMDhBJ4k1W2nuvvG4PoSL++I7E1xrsIfeJhvQow57pTmNd1iTHl0tZ+KB32HCP2DPm+B
PRGUOnfUi1Og80M6hpoWLIv5kXq2Ln40sXCtRb6WyVKLctzCGR0S8Sru0iaP6y6USXG+vuvARHLr
VgYXFK6JKYeUIgdEG7fHXr+m/11leAo+bwvY6nh0xLp0m4VNNTejKsshjFKWgcPXlJTJcHJ4Dj2m
362Lt66GNYmROk9+aVxfHjqWyOV+liJ+LVU+Bg1AgAZF5JAC8p5Bgp9q/SUj7Qof2zjfn3wZYnvp
IcPc0Eqw3l6vcfJpFGxpZiPU7Ux+U/ZECGty350rkIVmE+TkCAd+KlasR7a4mQEaTtqVU/0IHYJe
OcAjahCMyjjj/2pL1HmpL3LD6opdWfEwhDFA4UiTjofu980+n7+GzD91k9MpoOR67azyz9e4RVAD
XA/c3HgkgECMo1VXvqzR83RiViDlVQzUpCK4R7Los5XJ9U+m2p4duipJfvBO61w6JhmiZTk8Tz+j
syfQ8Loa1ovWNhYVz24vn4M+8jxvd3eNsRQC3RMv4/Vz7UhavLSrPWBSZ0+NeyWdnx/DGKN/yvwU
18ZOzEPheWTNb+B0wXGgLoly1zLCxD44e6xnjUFkPIW2i7ptQNF5A8IzNzyNjLUWxjF28BZA8Djz
Uym1LLmX1iI3urjs4nAPX0CbEZODAeT73LpKutJsfTmRZaN2pnd/19KfNubVWIg6eXHP8ZJwRhdt
hPVivub3l3pg8jHkGJGwoIxbElQcCSRr/zMQgj6JSsQptUVFThSJulFvtyH+ExXeQPfOPy45T/nP
5RdDKydiffSIHUDgu11LfZTONlj1whjGerAqf1ThOfoZFygH5iFB5e0IZRGDuzbzbmGYsJ/DhQt3
AzwUCH2p7aq2KBt6wQq7TbtG4UHWls3kLThqu5RS7ebwBZjTiTPBi44ZDZ+8kuUpH6TUOimhjyN/
c7Na1ydKYGOX8XAemHcSEhYRdJe6gt0RTHCYxklhAjRrAVzwnwPtuYlq7UAxQ8EBCKDhUWeFLN/g
IP7focjUC+ktJkYz07LZ+VyB0GTvIgWoH1b3e4wl5QjplcxPf6Az8ODg7UmIoLx25eLB7QIIRvfZ
oXR9t2Dtpragxy1gr383d9oWMssMzDKnc2rWKalFtmLUHzys1Y55csqMJLjni5qH+6v+5cCLTAwI
gPT1QOyUgg6uZ+jVBQztlGm4MnSA5aEaaZOa5U2DaGoF6G2Sp6kzEa1UairZeLGxPeTFSLlzQySN
L4B5fPVjuFne6ohdKqyTLba2mJ2ff+lg5OXjEBPNgi8n9sGnHqv27TmTMUWbs/19HsMr4slWMYHf
wvY3ZhV5a2+c26risMRyNNdJizIlUjfPmRyknmTo0okR9A1q7FmptW2teacpNNTvyBPi6E7bFABt
kblOfMta2AexgMQbAAQGLssMs+shH70S09oV3ZIAXcaCcLz79RBzan5iTD38DrwkITpyRm3MNhKB
RQtAamYJOCGZT/yaYjmDTRgBmXO0i95R649MxtRD1rQ+MFQB0qYuWOgVDZREQo8na8fSbJp20f3r
/gaOyXcRjwhxyFsStFDuk6Tl2pQ9BnkUM8IzGZyNU9oEBT9JrNRRJzDt0zGW75jTxqax7gNvmFUq
OBbZMm3XNYSMJab6sXtz4wlV78SPWOQPzDg9H7tBak6X8pmmuCDQiVkBgPJxmbUxnGJceZFQbani
IzsUJAeMlpVgLhZMbwExrJoUBwm4X4qnA4vT2o5sZXoE3iwWuLMQzT8QzAeMA6XC7T0LJWqsLnnX
GhQ9GVvv+7KheGZkXGNZXjL3xWkbsucdERHohqSSrNLubLG9jnpxAjU97niRjdv88tlhMydSNbmU
EMJl3h2E7rRyxHtb8GxnFnf73oeQIQeOw5UoOjE56AAW0DKbWXdsTgxeu7DBjFfnUO3jEQx0VN7t
rnKLKCI90zxYIem+uMA3ndtGYPY+hU3QIRIbnxg3EQWVtxhsAkimt4DJga+oF41oSNKbW8Nwzuw7
1cjZmryu6sSQwCKpykuTwcR7FSPPmyJZmORF3OW62KPphsuqfAtGMYRrJl1BU3XLe7HHwbmaZHwg
fmBsxJLDivFq702FR9s48mZ8CruWe1/Y0of+ydpV26h+xeVtqEG/v9OWMthbc+GrvIl9Smlxj+2n
LdQr58e62Sllc0TX93HuBU9gkEu3hyvDltAI9UsuEoDZA0AQJSCAnNLGJQdlGKXkcPpjj+quljkI
JLLZIJhE316VAuMA4Pj7TnsKxiYGKuyenx2sCuj0abRjrGxbcHhq2zY6jjgtgnVG2hSsJHkfG/fl
H1mvHRVvpNLr2yEB5zXEU2PiHYCsz7bXm/LNE+g6o13ChC96YKcsuF5MbC0RM/WxLDciQ5pbbBLV
3mQ4FrQcZ6qUkjtVzTE8ArI7oonpcS+jeX7BMQkKUwvDqcRC8Kfusb/w0hutSAcra9TtidPcEapX
1Pr35iRiFjJDjuAsVfK0bwKKNKVXhrxbmj31vSM/gxanNDw4Qr8LltmZm9ROyDej/B48QembjEng
E1WGyxkYd5BEmSwV+2iQ5BcsE6n4YyoloyWDoP550A+lebr9F+VU8kqnnUUHbNXRc49/ox8Rgvzl
qJ+ZbddT6/veisiOKnCm6tDESGU9SI/vWkbvBntih3MjeCDeqAh8wYxVjrRQb4oHsQjhMU5ICEX5
b3gEHl4kXTSo5BY9I+HHoqPx8Xlz8PO/PfiEa1M6IIS3nPQqCRKtcYLqKqH4srOCe2a08rSH8O0b
kcBwP1d+LbTy6ZZCV6eEXQhh2WYlmr6Mssbr8AU45IZrUUOr60QXKe1aQzkmA8W2zntla1HGxNMF
eXgDsS1JdHOki8aZIRxsCdPo3ArncTHWdth4ykJC2GM/w8F9zdCOUcWZijVKAv7BimWlHk+yJBX0
sk3zi8IqA1PEFFDa4dGQX/0WXdIK9ym/N2KxQ3LoAPfG8Sh34Jb+Kx+60Vs/xjb+VA0XYA57WZF6
vpjLHSIOoBikkyF4qk3L68npnyWUjvoyTynxZpjxF29SujiPrYQFh1RfBXID4uBl+BfXPP4wC0wZ
3R7JMbzPmdRjVgIV2cKsL5qVsr8BzpmxIBHwXYE7MvSmHqzNMgdGac3/X/RRoCcBwuqbTA9fgNCu
gaKu9eu9UQ00jsJr6+rg1tcwRkFvt1hv/k7Ent0vLtqhTW2dC653JF3mnEmKRNorteGllCLaS04C
vs+F8v208stanDwBg+H0duN1R6OCy2pQ5D+Mv3qp3u+8Z4dkVeW0mw+HTUNdWaDvytFiQauPXUL+
7D5lmG7okC4wE23TJbhNF98cQhSMNjC3YDh8KBkUi5hYpMX99Rym3j5oGi0vlhN52w3wR/dUxRR7
ZTb75Cb2ZKT1jbrFVMYXat/+ewdKUfuwzp6u/b3bCouAnBLMR3CB4B0bQhGlg8Ukk1r04flfUqhM
Md4HTSpVoDtsTTopfmsvQKTwuazc+auBrHMGi0jsQYNj85jB8NDRbxR/G8LmmCpnsHOjl6K4AmCu
7kAMcDwi9qpjHxGkNyZC5DFjjNP8I9paFV0EAGfJZnfIP2bYwSunFMdv8b/mR8tTxHkN0un2Q/3h
ZQkkZwvqUQ8osRRxSriVerapFVW9YGK0OmwEotept7+MljOUmGYTjHZU4MqYLLeKEZOEed99p9sC
wlSo276HZxgFpSVDsK3S2OYKR6njjTY1ZInC8NvKW5emiFOvqINofoNdte1CPYtTkVpf8zz7cPpS
yeyj1CpV4nEwdmOYvfypckrinAQgaZ+JuERZn3bX9fEO6sGXTIThpnKTW1o7cwnhZO0HH1dn5sYq
/6tapfxbXvMiUq2EEaBPyfsMsCGbFIFsKlr1PrCNBLRV3SjN+gnQ0FV74vQFotaMZwE6sIhNKZqC
u+laoQTwOksfzJrMciB7VNL6hoPza8E5K40MTuOun4CvQpxHEaQj1oV6W9LIwr74y0FkX7ZRo1Cn
73k3aIETc+WeiqLAgIKkPneG+laLkLLfl4YmfLJuV6jZR43mLAeWdmIdqtc2qVqHGcxWNJSYutFh
Gm2wXfxVu01RZIJ2hUhfeGkqyHhALzQWdIHiZmTx6wXMPUIbQq1tPMo9lMTC8hAAwubKVNh9chGl
5ealrZj4MyREdXWJKFnjWC2UKfFuvrSUcgb+vWwQ4FVV8gZJL7zPs/39OYagpAgoKphm0JTtebzk
bTHU/sI5QA+ScXnnbypN2E/sw0DviynRX03hcMXMeaF/LuxXyGq6Wu7A6OUSPlWAgrSiTCPc2nRy
OGKwjV4uu+OIzBx+eA7XKDUXsog5RxJgHTYvnvGwYTzZieTx4Jl0ys6zZuXMuv3ALw5EYoGZo31w
BxfYq9Iv2rVUnk4cq3e1ZKwLoJmZ/66vyrwgBZr1D29dOica5fLvsfCicV0xFFmipX0+XNSNI56U
iT/v/0YqyNOw6SKgwsKHwXP66X+/2YHclZPl8O+/IS2Cd8M1I+m09p7UqBhmboUF0M8pcSa3QPDF
7bAmaGO+UfM9pmTE+ZoIX2xcxhaY/tvOzyVFvTI3Gs7VsMXtZoHAvxMNcK7ckl3eEFPtNoX5bxwJ
Fmt9+0tU7qy8OHQy5W6nQEsHwTzyhRTGUhLZW/El2TFFAyPZpdaHRmYCMP+IirXDFirAXTAEl7FO
kHjeWNKUv7pqy9n7Sar+YR0fan5FXoAdHhG1hpIme0YlpUp+FkT6FDuMvPKAKSyJNUp2r8cKFjTY
CzGlfw1smCUZVZmc6qGkIbwoR2zyy5CaK67YNIveuTASEc6ojPeGmR3JLpw8BG/SPtY0WrUdgfpV
9TnSt4qYB1YsFV+tEP6SC8Lwa8n5KnZ6qqtkYRoUCKLCuMuv3nM6P2EcfhNycUInYJT6t4rAHN1G
7deVnjIW9Oq+ZAtudXDguuT7tfQGQkpLyrnGozh4SvluXuhpbc7SJ5EYSKkMn4WVu27LwZhcasJw
rt8Px5UVA2ZLf/FeP7iSQoWh4h2bg5eGSe7k0EPttmyLj6l4YkcQv02BSmjlzi+7GcrUOk/N1Yvm
w3RdWaOvfNiMpdZOpchxy/ZJXZk7HKCAhWkGIDS6lPfHgZ7xyoeosFKTbaIKWXjtan2EvFXfLC/G
b9IsV7UrbJDSnmLlgRHmurw4R8mV6nVD1/wzivALjej04lbIIVBBbuUuMMczGH8nUwna3LQPTdHv
aOY5tj0jDn47LH8q9ICcIQa31FdOE3g4uc4h82hcwOgEiwtgp1UPA/yEuQp6rG5MAfgUuHPdgbct
i+76H+vv9/S0SekuuPH+JoCBXSNGSd4875RJ59rCnb51Y8uzvBjx9+OWSyk/4PkXAcVEIb7CxjC/
yzzZVIYb9+HxXssMzhOrcA+wQDO8+p5okA7UXR0/gW2nU3b5tR5nWCUBSHSeT8Ewb7DXgMKMNjvV
1nHNxaSURwffOpSoHyusHCHi5F57myMWzyVkIkD0bKjTdA1XtDk7r8YTdW5bG29I3Mm4nZt0bNj6
dJ1Zq+vvB0t3Dm1HUCe7NqSkDuAo6iHbZzvb/GmmZO6waZi1qJ3aWiMnmdlh74mkwTuyu6ICh99p
Bt8ggPMvdLYMSHGGCHqUC/gyKetZBl3oG/yXbfzNam6dzBArVQmmMzJNqU8eS+dUrTtIHNy1VLYK
Aooo3/9088H4V9HRy7VN3/A5Cn2Gg7HiZpicjUUfLLPtPj7/ZvCiXtEpIaq3fERJWv2RNvFEODgl
g0Nduvon6Hhv/59+7YYhvkzeeduz7cPiKNgihqooQOwpg2f23s6q01UUD1rsrgRWxr4wFH+UwrSB
7THbZTj8ylB+oW8qqRjD4w5CNJ7G7wMZUSPylEahjtj2OS9YZ8TBJiP47eqgk1L92KBb0JfBQdE5
M2aJHWC37bsJdTQ0bMvwwv5n1hiyHJ2mGJQuvnNOFnTxzVnAdElG1BGcHZ/ZaTiyKDJiQlpFOAob
lbKFxD+pa/66S9cHKooCcYMX53uW6g0VoV9PcLRFA/gquIAFlecKWENG242kCc0+Ooz8ShuQhIQT
sJ0ArabenLTkmpALgAC7yiQQ3ZesLAZvlIa6IN9yXXLW+1SLbO5+j+j4hPxDN9u0N9ljQSVGkawh
EZLNQ8Ou1kJ95ZTm+lkjIcuc7PBj4E+agc48s/9AmHrQ07tmtxy2r4snDbRvqN46fsuCzkvqrVR1
p86us4Utepn+sOMYbaLiWsdQT2ZQiJfO5rtE/W8u9Bi4aT59hpDvxCKU6g4gszn8wuKT7GIueTyv
3IDtUNCU/Y6f06m8PhOvvIIPS4t4KgRwubswuDgZfSjWuyV9FPytMz5BI3XN3vs8mRmBDmwEOeYx
AhmjemyZIeSsH5yhfo/n1QVc3k1UjbPCMJIkc0iLPNe3za8D25vz1Oxm2I/1/iCQVV1eBK9MQZmA
0X4hhr7jIW/5K2F4/hw3yzDhR4EV+9YLbKDRALVgB7MJf7reiKoucbmiGWSkhUUQo/+Xa06LaFTM
N2c3M/IBvn0wVlfB13Z9nVOiSd+vhIpiZJCIJxbVC9zG9/yatdGUFXo7sbV35Z5nvTScs6EJHy/4
r/+/rLKbk7wBY7OVWXR6CCnNBmIiAOtIpQqaKHJViLcZD/eQOU2m6TM1JN9sC5s3fyLW016O6LoJ
aEizN+l4/NVqg/hH/X3l4MkAGO2HMXDxRfS/Aun5nCCKpEDwsH+Xdzowf8vCdxv/dJpX/MsuaumK
Gh/wST6elu4i9cN+itfB1XuakOiPtyKVWPMunZ+xnKYobfHKFJ17b+4MgDKL/yDFzYBQipOYquJX
cM/Fd2/JWhU45dB15EqdwOr1Jb2maEH/Btl8MBCScGz32DkXM3X9LYiPpoS06gdVDAEdS5zI8NGV
cuWVLeZuZsCQ0nyM6lkYqNvUS7wKsobEpSomcGbPy7/Jop1w8/kjbeWwXvpj3FenZsBgqPsKxD4l
ByoQYJD0bvPYtl6VXNk3Ji6UEIZ4CIFYWWA5DI1BmejvdhtwmdWWV01Z5osZFOJH+me4n8258+V4
MRNqbsWAp+nnkJf/MVelRHWBiNMKWjOX9X40G91vhIBbe9i+XZ4vZQmiYCXdMJCXhevNrVzpC4QZ
9PUDWUBQY5HvFuE9rRiVR7nuEGuoj+pn8EUw01J+sWX7vA5Mxi525dEsXqDWMnh3gSaWBSR4rR8a
Uwf8M/2yX/ztvsOhVmyo+i0uUCKwQFnkdbzQZG0mWrUMxFgglUdTICWcVaq1XUZfd0b6Hb89YAKS
9bF7jV+83EQhthmvgLiEaBE59pfGQvfUWq3xP7fviW+cpYo+nK3wUKd3VOxF41iMNXfCTxSS8tD+
PQM8tQea8WjAwhjI073XD0bGtqDmXYbMVy87i2Ax9SQhyPL8etOS/CpJl+RmuSLGe1Z4HFzE2JJp
Ve8BrF7dqGeEl1R290IY6M6bjU5NmAvDG4fCvqVI8DdRUwaZRyfQz98G5zyAeNJOPvkMp7RuDnEj
hfA5eSuqArw8rHb0fOAt+MRNjTH97+yrdvbwbnOkZofCq+y1FSJUwr66I68mXQoE6AfVrXKcLbgs
Mxigj4/TA2fGKuLtAPAcOBFQQ9I3WBVUsxXJOx3nTrsCZtuC+4K+688bObGy0K0mklAt9Te2X2Tv
nH5PggNMV+hlmBssJ27gQBnV2YttIgaqWdQyRhoMVVYu9Z3sGC8ZZVJWooxIrRQRpN/0HCmV4hs9
yh3RZHU+xQEBrpOX7pYfExdtukG3/fMUhbvgvfHBCWV+bTXkO7WTW1kI5v5aRxSCGKY3z/T+TgO9
/EjOCWTGJopwzGMew//P3eV6oIZCRD5iPPBDq+QQPenB6suj5pxdp8eLZPxbaHtbfonVUckotL8t
CzmxhTB4xqFG/l3tBb13EhKoGsSklwzNXVRjtf8WBB4OCtO4Kd+3hdC1zn0XHIKRiDC8FOmmsOTn
dofR+NvP4dip7tsK/BeyFfLjLoiW25oBwLcVFO/g3Bt93eON51DXOxceEfE2vKfq0R8zprLiPljP
YvSPildsfxmjLPTend107UI30F2aV+7ue23oZZPlEzABABShMPvaeKNa+z8J+FBiNSHi11z8a5OI
3X3TBE1tEjBgnjeqvQbBD/ZpUQmCeB5SPyyGdY93dt/75+QVdIQtwu+yoR/3zKnw/1+HVajQjx2l
3DsyGkZUo6JU1CX+V+ZHyzqk3U/kaRIZBeA79j6yfPH0pFmuOZtx3mUIbLqL3rk7eMHFubSu4OuE
P03LXFxvDcog+GbjSlbhjaH+e8DuHMt4bckWY0N8+vGwceeUkwFDq+UMOlh9jrEJiiAhm+j/6u5+
az/FHXNfvSXwxAuVz06k4xmowT/CewPEYvP26gL1f5ndTi1X8PqBz7hZatRs09UXvuw35LglQIeO
gMhs+9vCTlkK6n9wc/tzIIpZTFY/5miSnlrDwoseLIU7L1iHM5JBDDCXrPGm4lGWxnuJ293rW0RZ
MvxqE2M+imfoshNuL3jpCJcyyv5d5I/SP9OQ+bYbiPEKOsUoluA1uSOldy8TJJGpfrkSXiFDpMcV
afyazUno6r7Z8NFlIE4CJVwygMu+aCZLPbbgm5eR9YcmgtydBkBdzuoaiq+haNGcVtAyGSh6Eni6
Ub2NxvOhLVFKV8onWVyq5+931eU/ySFZU1uLssOfpwkBJuxl7VWB1Df/eOhVGqtsfLp/oFxYudzP
oXQBEgPmL7JWLglzbUYhgGzeS/xzKsXaztYPJMq5AkJNcrN3HQKa1a2xwD6ZMWgrDdRhzoeI0nEX
rg+X0qxyQy0YV5f5dd54l295cN+5kvZwXtRYyqPSbrzHEDooMx3cM9E/K9/TuX7hDq0kLQKWIMIA
xWEuB9RFfv1o33wWOj0+ZOEGQwVr5aGVheGQxng6PcthTREe+nBbwj7qT0dw0rqolV1X1i9K29uQ
o1mcjRB2V3JWR9DN4DL5b/1JdgTjv3VheGrVLrZNEQqvHAdfZmiPbBZoYDfzWPpqsJaLCx2NHtl7
+pW1PNehzf6DLksY/FtQY2k49URlK6G9O2RrZfd29ArSAN9poUw8hBO/SOWh4I4un4zqmKjQVYcM
KyEh/OmusoFuXYSrHdMy0j0DC5o1WCFDUbH1cILA4yh2DMUjg0JZPlctWCzJ9e27+togwIAAFQKU
OXzSBwaq/HSpvuBAq/3cHee6+ZRrGn9W+VHTi0miqKkKqIzdDK+I+9Xzk+D/4+QLY5sqB7UMGuFL
bhz8p2Raihc8RFg6VTvApZ+EDvanZ8Eqt4d7RbBnmDwsLTS633uM1YSusj1TWTbUCgGbJoa+QnLL
PFaUy1SZfrmhpyQDzrrqPyOxAYGjBVtWi99X0vaHDOcfjybT7227KdXSPYbYAtyd/nhiiPR/6fAc
Cb2K0uiDIdU2M4niBGveEMdp+JnbYcyAXhYlINVaTEjaTt2R5scBEiP0h0Xt/boGdM1czvwvHj43
kLK7SS5HjhEZBSmw0rXC12iXvPVSzI1u9Iet/mt53t6YyKXx1OIZD7dQPjX8+SpKC9j9c2iZ3/1o
SYPCKS7N8w+a85tQNR+WbQ8YCkS5uZnLe3M3RmeDBwpDBVDT1+YL3W+wW7SrZN9rwlKfvDYlsaoo
H4hE3zf55kgyPFcXmEEs0etkY9pJsNrz/xvAEDn0Q2twbM+WfBexaV09UJze8w2iOuc3c/dPiCJH
hTORvzP0L0W/EfMzQZa6EQuXv0qxoNq2eCBpiRPbkLRJolRsMmkkMCYbovc0+bX/OAAowTdWTzPk
WgmIxmntuKNRNtwehtNkoOtMR2rXTyo2b12RgBfy/G79c4qf/xRlvpmGxC1rXGLoVn7iyuaCS+WU
REs40gB7UrcPhQHY4b5thU5ddlQR+7hwfGbtbDfGU3fsC47HOd60N4u67sJzz38RDLKooZ2YNUDO
4NOB7tH/IxT4OSWLnQ1mo04bKAmp59wUf01nHDYFWKsDQe+gzGaH9ulSBV9yymCIwSj553KnKS3G
f+lR7lmcu/SdXLclNXQpE7egee3TD3+28np0tZR+UsleVpCBKG7i/8u28oN5PvI346844v9U7mYf
1gREHJCjxmK1w/Em698CKH0LRm1T/Jg+ZupUbC6OMwwTgrd98cs7bkg/cj+arGkgf+Tp5ePnwSbV
MesWHvjy9/CnmGzYkq5ACkCjkqq4gs25IhkvcBSyiUVWXPeIxw8bs5Be7mHAPraUuK0C45VrF11j
eznBF0xMv6wNy29YPTDyo7GcBKaWfbqBB+KRv6bKEk61di711Z6K2wHr6KpfMwjTwZgLpzxsFPex
U351raXhHwroOTo7+csW8kefRonHC8WyLO8hXr4qaOFuD6wT/4/AGtBmD6S2WnhphH77niu9ZJEl
/5doOljleJLeeQdyKHB1huJQ2ymudMY6+1JBSN7dUodncRRa8FttyczSnbMxg5Y2vY67lSpJFW+e
glcZil6fiK70RABzZNqxVXZUvze9xjvDQXlVprFjQEJsYzZdpHWvr00i2PW3vB1AhURcjhSOpnjL
jqp42/rUazJNdptHvxIWdu4MJoFXu50ijb9+bVxgj6/osdl42lQSmYztwx8ShUmoVkHTmYXwzhge
uG+23iD06zqX32xrYjVLayVEfyE5VHZr9wF1mG4s4CVFvCvr742sdNCICWJ6cCwQpzrmMoUBKbED
HqaizgKonvfdqpRNkutO4YNlbRMdxzz0zonLTj8jyfBAynA+uRvEMfaC3yz2aBkYMA5uCrhXdfJC
1M37qxiSPDkf1UyUFnOow4oVOOpI7hAR2fZhvSMAODKRqF2uYmOHLTc4cUFwYanYHCFOnQGFGTWH
KdPbYtAVlI0MbvQscXUG0+HgoFg2dMwSnabwX2LZCCP8+2iuuyFiwnq9dhealCYOuSyIEXkDosRn
jKwhwDJLzBSR4rwFmGR9zp0ix1S914x8bTzMJkbWhmcRvCTKmsPYQstBFASiA4aOJPsxjvmRs8vV
XLSBkvdleDMsnWeFY8k5iHNZ6aZoHb5yT6LMQRQhkIUnJy5xbQjU8lQGkmkU5an5562KTvOdYCS6
pVnW1OFV7z/hzHrkyTypXoHRNh0EKZGB14qNJlrfnOj2HFz8QGvkDOeexcyvA4tbCPP5cGC9uil5
BkAaRxMv1oZjLBrgBpKFTgelXoLA6RGZKqUXsGXzg+kfq3GLDJ4Mm47/OrRJE3tfO8uUDQIMK6or
aQZ756+c7YlPDQ7mYYmoyDl2p53nno3Y9nMNKbG99UgTte/U9f06+5S+cMv956eSB1pGSlIA3Gi1
EdZ7+83Mrp9mD4qEhvDeIjq8LVY6LTihu64YjhCOnnnkqqQckKy040RUuy7bKzt5CBLoWT/q2f6S
A7WY6BqOU033HjDFGIF1k9gJ34CaFN7iQvfqTUUM3e10cNOGZykbacxhO8KqOWsyIMaCWXsNrZK7
qWhth29C8MNGyQkbUpYJr85cL8Tzfj2a/4AAT7d0qOisgu+CIN90JqZctVZXLdKuB909xKWEKHFR
HmUZW886T9hwhBRVdFDYPXvLUcZU8m+jON/PkdU8RrsIsW6GcuHrR4QWBeJcg+csAhyrKSwtGgj5
+fQQYGb5+tEonl4TXwl8VxaMY2aA8d4VxfoY/uEkEzXZl6EwX8qdQDjVfXhgA6d9LLbeDuZIvbR1
836pnJFghofdMvlAazKKwD0Oi2KloVjYAoJ5HkMoR5R2e9k75TtsIZ+L7+H58ClNBAiQglwf2H2O
XPpUVJ0Tn5THlN/R4cuOE6f2VxqV1E9ITY2s+GS6OS/L2FyZB6TSghBnFai48/8X2Cp5ykQh4BuD
bpSVRNnqM0uuAwEpO1mvKqaaoA3Qs4tJG3KJuiiYFGivUfvJoMRRyotLGewPsw/j8IkUdhaJLfHd
5AXWM15AR8noCwtQ3VMIgglbTPpZ2nJx3Ny4Y2XjSA00vkY8vAl5x8z4fjxh+GvcZE/gehHVhoru
LnhaMQPa3JFVkPTEfmKzJ/xeL7Yuul78pK4r+V8jkElskTz/kOiLASR5FvZc1qjkusuGodq9+MBA
N8IVSVnomYQ4HPxKB66g87FX7xXNndPfyPbtGYcmSnIRA0s+pRqEVMh7gKEwckxzT7xnF4ERacaH
c+IRZIIF9NhH10olTI+ej2oVaNq059bbBjOWQoGGbdgR65OH9g24CXXxq0EAHhDUFfDujDAATEbD
4vBTC4kUmusPLOflzV2ZhWN7rqZLebjKopiBE8PHThDCHa1hoCxu3kb+j1Pns3nONRSekRwwws9a
At0bJLMyC09ouwtsH/+tCw9QKuTWBnczsjzFTAWSRnc2Mro+v5Yv8r14vkO8p4iYv9ru2SRMsg2u
1F60QSsZNdS68vaIqZvqR2o0DPEWI6YXKen3L376Cmy57/Hm3x6Xn8cYC30K4C2Y9YdN9rK451p9
pWSTN6lRbyPurGe2RICezhNyz6Xy7X+7z98b8INyubNS/DrWarxFCIcQ4EpTsqztuSq1UdtdtvPg
2Y1z1fLtX+NQE69Lbe3pLOklPyORnOo5SfLkbWJF/MPkNdQYzGiIqdMViNh5KrCocRhXZ04OLmAM
X6B+rhdisl5o5p84/F3ZczGeIUv0ApJN81qtJf7f3dIQaVAdUmZti7KOVInj/vnAMrYeuzEqkgQv
jEpQiVORA1PUAZFSnHLJO9VFWJfYzZAExlYI+a8+zxBDvUytd34dNtueO5yTWEcvUBuKLXTwtCWr
I5/9L2ZDSwjQJ458VzkZT77JGCFcsAysWIZ2mblXJqcWXtOzTwMf9eeSTlMa/5yy5SPF407r1NJ0
Ll9pt1lGF9YmjE4QbgkE8QkBjEiv6JuC+mfZTpm82oyv1LcADu05gezmdBbtd7UXNRrXEq6p3aBQ
Vj/imvygEpmEce0wtP5O6tpyMRkSV3I8QDswuaWQuLuAAMzBrHeDmKnqCC0kQQogXeaZvpPKLS2N
wEIBlpkwN4DGvv2mChe8q7QCgUpKRYqVo0NqgjqmiViJm8J/k8BoAA1I5MQLoNlHpJu6D6rpKyX6
MUmiJ/iTy/6YwcJ4cogtmz9vDWVig56RTIoh0uPLPJ8OKYvMbDVMv2E19eBmbNzdNju6F/LXu388
JheTAhSDmMaxuT+A2rsF1pl0IcGLbKjGBhNx0lO31T9ttl9DMMR/X2/bIO2vbScBMOUaY/aqoz9C
gjU8Tutl0Ks1d8eJKPJf6YVpWATg91q0GY3ZLASeiyB4shGjdG+T18bfF4ZBPXDi5UR/4Ysc3SY4
4SOTjWT5aRP7BF+dnOqrXP7Gw9jVewom4WNVWcqnaObe/RQ0xLnSxqf3vueDJ4XNlQnR4QYR1JVi
d5yIwAelpuuRgo1zRKFjppagRsxaAKgdxVhEPbG9nJeAqBbJevp13ofswgAyP33jB1OgoA8eyhaH
txliX0VUdY+sSvYkDKpNKp1zAJ+f0dT6bAaUqi8DUN19OPwLTVQkZ0HqQTj67fRfl+pJjeutWzAV
JkyOExfHoj2/DRmCTt9b5yzwlkLz2YuHpZCZYv+0FQX6V8f7ui1i3tl8Bggq0yiT3DAlpYcaGdwv
PHee4hQhhHdgpQI4awevMrJXVi71BIeLl/HvuZh1k8I3QKOy7vgXdGjOaH73Yt6RSJtgVL0WtwRe
uF8uiPSEsB8LjuJdjQGeuHVbTpDFjWXQ9OGg/a4RQ9GlC2TLZVoxQBmw8MgFs/j6yDAkcEfDHtGJ
ua7Xjo9ugvPzfzPRYfykI+UXC3ahRaNf3BY75YddbgyiPrMxckFxdIe26u2/XwShuKFUrRRpq+/7
AsEH3jjCbNuRyU7jehg4iUbDxXYRVfNB7Jc+XohrrajQ5Kj1Qn2k7UyeE6UA1f16FMr8qZ49rAW5
bS0yldbLxO5ZNL3y6Vg2QdcuP9DgEla+1GvMPRTFyoVlgmiUqQ0bWW5ueohNTS+nSFJAX9nWGlcF
hJi56gIM2bm8tv3F+uW/SY29+ijowGFKEbQ18Eu+inprgVhncQKs7NHeKDr1s5eWcvbW2dTwZ8nu
QXEYsYeMlhLNvgn/Za+OWNlnOzVacQTFjWjaPITZ4PEUSGJ8XIA4ln6Jbio6o7Fz4vx0P/I4Fu8r
IutVlcH89Mzz9v6uHuCzmM1dUO6iKuNJfcs5myJO7zJJ8sOe77VfNj2e/IvsyEQKrf8BHcc893lw
ER6Q/3m7NQ8U5OPe7nP7laLwz8kQDSPkN8GC9f1VtNyghxkVj7ypJNb+WTgy/RUNqcLCS+eywtSC
WlXZq1dB1bhZwu4Tka+Wf8tWYTW2LOKMfq0Rk+v2YhGPzHxw+1/MTI0xpvNeMpqp9q6gAD4vqwxK
q3gyPGXPcaR++F7B2G99tGliVww+nk9s3P4BH0PD9QJ3ss2uxmHrPqRJ3AWCrScSDmAvNuMrTaP/
+2DnT8C06byUu5DJrMnS3RnXrWXHRxHGfLz0sbVNlimNCE0fHFGe7iH5g96koUZMQmkxHGg55b+8
n0q+exmWlg9LeV4LlrIWrztS/VoRZocHocyP6FGL5Mc0XrZAq4Ww7Ujxbk0x9XczP+cPxbG6x6s5
ZP4xmF0TEg7wbdWOmFjphOX1k5u/qxfqC34lEweTXuvO/B44D6ZJ9nR5ODq1L2tDs+QV5lWfPr9v
sgfXU2fErvdnfkL8tqZ2zNkcS9KtZXpR2P6iQa8H93JCQeP8HjMboj3WAn5uU0xm5jpmUz+K4RyD
+07jl6p+PiQv9Ufo9SKlDJpFPMgsOVOFqpY5zVXH1K6l1f7Un1j/Q+pEuEh9D9FiQUvBfBYfbJN4
rBR59mBtu3zurg4SOuTAcrIndtPvKaKKzbGqG7cXvsvcp3bkNfkqcY7aGsYZ/H81Qy1wdlT5Mku9
4IQ/nVh7KDfmSgYh4f1bOhTiZKuW7bhotTJgUR1jCxpa0okQ1974sGRWQKIdOSzLNFLG3Dfnfzot
TlVri0tKlk4uynF0dedpML9yJhu3syWqX1KVeMT8ZkHQYxdB+Drc/5H9gNgGuep9UGOSpAJjx4a+
buAizcLdH1ISRVAE0fKoQzVqjIIy7YwUhdjfEqJjqlihVHtdGZqrSzQd+B8fFHrKLgfSREoPi3zA
kmF2JvaVUA1Qm16VzN5nHjMZFcs9dumYlDsGREQ0Rg+emW2cPb1uFvkeH1oFzu96upnP7sWxtzM0
ozmtfqbyPhweNcOUaWS+d4i/NKm3p6ruzpAb2hdyMBtqymIJmv+6rySoRo2NhQjgg7yURUiBkFMI
W5OGoLIb4bL/+o/lMkJs+SPl2m8hHJthefMuTTs8IU+EkCelKYmtrcpzC6jsWI/xlKLs0Vh8jnAG
AeLuF70iWQ6ekrLzstvWxZcM/zrLShcwoikooEC/XTEyEautNoPgRxwjx4mpWZrgM90dwALDoXmt
Sb247LLny/utpMibzYQwWwociG0JWo+Xv3A010s+P/Umd/lSV32T4mMBtIqf5e6trnEAOsKHL1Ho
YuRN7AxDSyORWQL/JxCvw3mjtFSHVyT32LVNYNR4vBNojtyAqecA5qU0VbJDr/TcmKIVrHX6PhUv
X8OeKBUMUPPy/18zy65UiXpYdCmUvHQLwz91i7KjPALPkNzSco+SC4LSD5C/H50uRrAtf4RhCy+6
8acH92n38rpv2vnxb8Wo9/7NzJpF5PMBgXP0OvcVo7fr9km74u5ypwFHTqDLmH9DkLhXRE2B6fry
2mUb6EcRTCFAOaebFYm1oCF7Rq+ZOWEiIb7KgPRLXfr7ecFhJFrXYrdhseUAwPbkrSL3w2hvvbje
HmDI9ojuxMvKwmO0wJuPCScNZN5qRStpTMpOq9aiQ52gJjgsqz/yIFibv9dd1SF413Y2/vWH3MYh
o4Donbn2cXqa/C5NKdaS/gijcUDm01fARcC+zzFzmnhRAhtc9P6mkXgYrY/b6JxRgUuwjTf9DmM/
TQLFsV6zDrGKYjU/OVl9NdZgf0OLM4ZIgnBPxpd1jLTtgFp89iGu8Rmtyn5b+79fQWoreHkVtipC
yrhw4yuWW7hx68dApAa2kL2DKyFo5l9nLZSR80S3ajgTsdNeLbxP9SwtQ2zd1hlLMAGEti+0FyDL
FcfDnySgup8EBbS1hyyJW7TwIS3MM5CWPkNbztd18XptZBTrLG5CydnzrxE6Q+8hSE6bOOW+kRlq
xDhyzUeuqtTMTGEbsJ0UhHmPkLUOlC2n129zGHmwYJeUlfzk2eUIQ7H8h1jOUuA6peiwBCzwsWme
wLhj6HitVVowVVhzOfg/h2SxBRB5mhEHEtXrHkJiVZuPflLvX8qPen/p1UHfnyIZ/ZPvPxuWLXWf
Q8Qz9NVVWxzFLvxHNc3fQGzOiCbtQCoun/bYwdP/Mny0T8phq5FbQJplugGOqDsnO2GzPgYvfAVD
PRf2rC6HC+r2EmmJcBUFszYl77CgUOYfpnqv7EO/gOF4zTttle55bLTmbg2+6LIpqBZzWsLhFNcm
K60VmdTCfUoi1RC92Pj+blmAaiCW3Aloc03pdYPMWC759gdLhQun8o9vO8cGCrzYvURMSxckPSRK
FMVI8J1HMYeZQG7jSBCkCwIabLx+qNGVm4SfMgosvgOGmRHGT5bm5S65lnxIlZff9pVQTu7SJcCP
u3nu13AoN/+enrBff46JXh5FU0lz/yeYGSVRm15qP8eLvwAynfc4rg7tIuA+5/2xOLWi7tPjKE2N
GgmEz2fCjKp5ZIXYZnMsB028vbZmdpuRVrtI+YQnakFq/4U1wP468//hyiiurghbI7/cv1PY4vy4
uqVjrzHvJartzfvIctqlVAdQFnmoggCK/tlc6434IBRlylsYsc72zVEngmpES+31uQwiI1EETqpE
n/AZFlLiKMmBZllCFxraSsKq5FwoL1pLEwSjCJVsj1/Z0I8lSJhRvDPr53VpvyabiwhB0E0laOtB
yUgdzWP7jifi/mah+M8IoB7MWw0QpzAcJdlPT3JqLzFc0I+X5lN7v+aIsDREomGI01mSLJT7YMUa
lc5Adzufy9NHUd7RGxfD5QcIe4kEOrZrRPxIlzght9RXQ/x3uqqhmJkS6jwYmbCkSYj4ItJfGSy2
AqxUi6MWtexB9wx4KB26hxYf32jezfiQ4/M+BKFup6l5xryLHcSTVjxxuAO8MFbaGPXgPV19zs4/
NNFVCYyQghuE6ge+nmMV4/LmLUdeNXRlx4zgrjo2vH/YeYKfIUO8TM7JNHNvvmVjccEoZBKt8DIi
gg1eviEOkRG6hos7QQNjbIGrB1ckWRgCwzlgWR5ahKzdNl2G9g3DPEEQNJGuuaF58QzdU+qwjL+c
jLHUmggYCBBDuDccgIInHFJPmysCvtoxyEIbFqM2QQ+T+AaeAQ3EU7vOWaqL5c/D/HJI/4Mo5Y4o
cVMxeL6NH4JeR6dAwTn6Wm/QJj7+Sv/D1rswpIYb9yylkZ/qiZ4nqWEUvBcWrpfZkS04mCJJp1nz
VfHrj0yFbl4KdOWSYShnHtXO06TJireZv1Msw85kIpCEPW7nmYtXXOiaSPrciop+fTbWKDiBdieT
uZ909sLGOuefXTqWZ7fEtHIlYNBGtjU0ACDw1qqE1KmiJ75XPIRuoOcZcXb5ZKcJFlcZLTypNp6P
GgHoXLqyCQP4WAmKnD+/sn5wRYnVE87/RJ+EcoaxYnucaPeg4UTM6C1tJp7+8+KZveo1V4637d8d
CyUOuFgxu8hGpuO06raWqKnB/wTQaA5Zl7m1DB65DJA3S5+Nxa8BmnhDBu0aZDfcxSNtl4MoNxc7
p0rgbFiBaF5sQfVkuc/MMrtlG3B1RfA5+UWbaaziwG6zJaJ/IWj70fw+MT243csHJKQVY8ndL7S/
IHv0AUWPoDNi4KtcfIOc0f0orijpQpCuL7U/ckLNPqjvrvwnIrlm7vXIrr7WK5aL3duxSyjvLpBv
KBQFenJSjNuJsjB20qLIwhpY26LQH054VB7a35q+cGB0T8SJWT6vnDrywZU4S25JbfwVQLY81mgq
IvQDOBdakyEG9X9zPS41xqvwDYrp3RWFuG9RDabnV9K/i5ESyrBW8OPc286XphRvdQdOpV4CdrOj
GrMByUMFSWX/wg8r/Pa0EWBd8BuC4QIA9Qk/wpmzpyTQIA+CbSQnRWP7lUw/ms4/2xfWYY2/DGQq
V0lwv4417gj9RTirFBFcTNVMu1ESsOVnbyS57UnPsLmaYdqTn74jR3XRJ6C/PYZULbiMs99lNgWM
enn3TXwcx6pSL6nq+llhkUMSXgTv4vCUf8U5VQtn1tZTPTCAPhBgZSwFkSfkXRwZMWnW/Rb/qsKu
GNoWFFjYsRykutW35AfNBtWC9coX4+lcGtRcEJlUIGSMwjtvUG2m5NKZCCgwvgPCEkADMA8mIzuX
A9C8LJLTLXVUlasGn4YOTsXqJwDBanhOIp01fq05cdA27CVO6KLiln5zHP2AJHoUgg4GawvttdWA
ypgbtDkPhfH/N2Zw+IF1/ZQU9vCrp9k76p0FH4CPqdDOu2kZ9faia9PL+84RQrYZNRIb2ko3pvQD
8kgCWy9agK8hsOiRcQdCSzr2uP4l/JChjz40G04YyuvaFZZukOhAsR0+w2zWb7WjMFAFVzbxWVBW
w+3zX/CiSy2bbQxGrtcuv6VbXcGtIiKkjUzJz7m/0HJrJsvBb0PHJv3oOPo/o2vqkKkw/5DPiI8k
vyUUcXRGtwxEqYspUelN8VMw0GrUUvtctosCtHP7XstMwxOjr11/WgrGZ4d2uncsdoDh2M6Un84g
xwM6tDfSi+NH5w9bvM1q/I6Hm+O7DfKzt8rLYjkBJt2sxYOa7eqmHg/ONw0NuT5Bvrj1tPkmVC8l
8L13ThUMm/llWAVPoXw2zdA3yZ4pJUf+yqJh4JVpp5PgBxprMGPm+wx6hucOUhywUtOX7ZSxzwHs
OpcNURRTGYnha4jibCHtc+Xfh4WgCyol4WqnFbMp5btuaRsRN+kdc5h9G7Yq2p9kfOBZut0nIf9p
UnNi7RPpczz54LxxIEQqhQSf+AexN4ZlkbzFnlNu6MLC+7UpfcCMkh0s0J0gWKrG9MNKLNwLybaB
aUnNc+YfPjOPVX4QZZsuyKQzP4vxm9+dU2pz5hhBwUjRra98vQh+Yfa6+eoJJzQIeYFiaw4l3BgN
TGiOdHS8zbjT4Agp8LCgRS2NdolRKlGbg2huEbxdoO22UBiE4SYjTFafoOLxcU2AB6npwXw4Rw+I
eb6tD/KlDUopJmvh5kStBR4szkw0dqkZ2fctQqQx+FPwhthcBzp27EKigcYgFHsZx9KwkXzKWJ1x
Fm6DbT67ws8zMXkGYgV5wnK3wjJRsJ3a82vmEStB5jr8c60jGOZyb2/px+37R3dvpLsKWKeg6Sqb
cM1OW1OftW7C4rDvp3iyE+4DloLTPlQEQ8XxZR4qUJ2+4KQmDCinoTIi+dY+dQ8I4PLwR6ifEUg1
0ll5k5PWsjqqI0xGSXCXAsAn2R6X/ckDqs/OaBufY3gHk8rL6TSYpF93oZNgPTBvsUxgUszhxd/u
9ZssTPO5DSWMR14G32M8AqR8X8Je7k45XP05NjsmRE2vr3+/fjc4xiEHoDU8VkXYXKzAR5In6Zaw
eKQTpiM1WZwmf1UZOYSN1s8qGieUjLKUv7Nb1GeNLZWfZMtbzXv2oLtAtR4tbxMoACCce17nEdKv
SndGiOk6kkNwV5Jy2m0Y8FyK3RXwCzETdRGXjwDfT3TdWqmuHoQ7T0t6v3kQxe4fslnKWpjj334z
ETt4wuvQjwAqU7I6seyl5Lr7ff6YNjhsvDbLCzSm3jA64W+m1DfY5ytRM/KoDa0uD+pPlWWMJ9ps
/vA1GgkckEmEylyZDhGMtCFeeP8q4+C/nXP0DLsjDmiinffEFjAc50gSQlb5qRlrQkjN6wQ+Jc+l
EIQNyqaqeMbASJsUD1s9VjHejunhMZ+wNho2foTJ+lG+Rtq55V2hmlITI6HDvblknDR8bfavEIQt
BF4n6qnNf/QPofvB+FhjnHH3jk4dvJnnlz2VJJxnkKUa8whygmMmOoOH7Cgl0+V644c0IpedeYeB
67JZRVeGzAsK1Ax09BHGywDB6oywMgxX+5NRPzxT6Eej3QN9a/+zFLxFPqAOMNW+nD+nt/byEbDX
3lNgLDxmysQx0WOEYPv7c8fWUg4ybeQG9wckRLBXWg3bh9ec+XTjwTkRc1pMkwkWIzQiIkaYmj84
PDM8sZ8qggXGToGZ8EQL8vsuHMHrzolZbelUvdRKUziNN+uTwa1sHggreXnD3v97JaSoMWF2P2FU
4MWBOrarcQCXQ5gcyzZMb31gS4eLbJh9cL/hfFBFspwnBtWAyJhsNMYrU4J9XmEuagzg3daI+Zoy
rxlJT/JON5qcNt+o/91DQB9DhGEAG79pRwHpj91sC7FcvmxxXWC1KZIRLLu3iCPNRsTjGKYkk530
1N0z9YBQPZOESJkueaovM9p0MMKs9BFvNdnMPOOE54V29f+T9RERWiPZyUnRZ/q8TFzAujeVsg4p
Vk6dGQCmGo27w/emQMEMOZmgziKxmOpHpbH0UP8cGjwAPnu9YVPDjV4szfIHGlMHeR7cLiCfXQKy
N+NKf6giF5Y1EsbZJSnQ6MJ7j14l+PquwpWmXo9EKQF22E3nK0mQQGdB95NnuxHBfGd8evTwyNJ6
EHUmGk38BPT58gxbf5G/vZ9bJaJ+kNH5HwKVRHEufb428JmCoQwRe/EkhHkO95qkHCCopPPLbLJj
PaXe4e4OtFsYMVB+hURxftvJEqAxCAPQfTHMiBse/B+eb2QyflxGWm4T/w+5w+MPWutAJRYnenOV
ASOuLPTLRMbK4i6pfgVEzCGMEBCtmxC35BKgt7MnoJj3OzFAvmYmgT8c6OwJza+qXpStmNScr1r9
qcvmlO+T0SSSakCeamZt8/oKwW8F1zrpmL90FDdKf8nNcYP3sQRsaQqmsm6dE/UgeaIiPGd0czHe
Qkr4fsQ9ZqJlbOopr2XUH0zKBXK3pnx4PTf5qNFAuNRXZF2lmN7VRSWQDLuaOBjvEVikUwwm3SjD
SZACDvADuGl0hm3NgDW3P4C/sVuQ3sk0Kwa9j3yw1zkOAfxSIrZbYsDWBO56QZjJBFRPkEolsOoR
mCss/15tXD/WBowZsbhoiKFvw4EDCH7CHN9iVDWHJDu+mzh1mYn1XoylKlOXdgszw4sqHS/EwI06
nJgJJWkzLTd83Qam9IpoWazegRFZYTnbrZwHxYUi6krKlzjOhz8BXpp1N+yddHixKIZUr8Z9lzmN
mJ0HnNXPR256YQ3uoY3lTOK2Fy45SOS3iESqmc/y4fHKlBXa24AcpWJQmnQZuLiRNPKFsZYYBnoJ
XtqlgItrda9+8DEL9FwFPrDaPBcSEAsF9Y1iRrWYrt3TtU3berhqSXb40Gp9NPf0tDCmYy8Nf5to
ZVzwniYGMW+x7lMDv0qYiseFHx2lwUb4mTzOIDmEXkQrM0wgW7K+1WV2hYrVipFKuvwXerdy2uiL
zc4LZ0/t6SGD4o3Hsq15icRNqlGMSLYcvuSCPdPAOPJ6FWaWRnGQt1Kr5rpVcfVFetXwEgdCzTgc
oZF2wJk7/ER9tmHSOV/VrSJHeKnPlI5MGn0tg5aoOoSXdwVDJdSWgyMJJ+aZCPlaakeXXpl9Aorm
CkBexjOYcVo18hnrJwKIq/qeW1Q0yXhOPds3MKAzMOaG7KS3CrYuqb2PzCePkIJmXDEcKE8Ru9o4
p53xyK3HXFUaPJpIFpXMhgBLy3zv6Nl6dolQz+coJol1axc86wk5u3egjHfVxHFeMdKbl+eFq1mS
ld6rBIimb+YdKR2gdtiSSe4pL0dG/8GNoo/auOR5O435VamzUNcyr6ohDLGTLFKMBFSoo/6JdAj/
E07wMn1zHYIIG++ayk3JUE3tthzdN3ExWP3XUxlDsNfdFXZY1URbDa2z6NbnKcu5iScQEaE1NJk+
huLKmnrzELW8Ph3dKdIy+sca/oumkojyOTaVXrHgjJMxDbY9vu2vdt7MEjQFpQRnF9wttLzecxd2
2XS+LJVTjv7TcMt7GqW/nyvJWpQqHYeuvr55MS0cRTl5pcObHX0thScc4nTT7kNfy8f9tbRuyW8r
CBT0QnYWMOFkFcI66iaD5qqAI3U2VapOwaCSWdA5+vJ6ujSnpRx4WDDk3N2OAnZjy3pphu30gcPl
VZpxrIF1UagOkqL2NjumZE6/ErAiqlW1MCiEyGrBa+eupzBd+92fDqSDaBPCYzOhdrIkdb1l1Ewy
0nr/p5Q9m39K52SWxO9Dreve5Po/i9MlW5F3XSJQvVDujFAJXfdjGKKVSpLvtcny5dZM3QtTAAKw
mA5Yemsq9gKysB9kwEUYKeaGCkd5UMIK+tKYwrQCjA4A5bh1UvoEC1YezWuhmTVwnaSHmJ/pvI1p
0EjH58NVhR+NhkKrRTdqpfm3ff6+8BpWDNC1EqSXBhQ4cgn2/cH4Ksm0TXcLVcSB8G8RHlEiwfWl
u77AcHBxKn0COCKnftZMaY9+4oIbZFPFILbcKkyqUhjjwsi+5Ar3F9oiqP64cB/ZSeY+pSz9pJju
PUEPFvRUO26wuKt//gYZFkJSgdNm081WFxrbGhe3zTjQl3rCA0diK8/CP/W60NRjmxvzjpJJ4bLA
1RHg3hguTOJ9cep1qtyYRqp8db7fs1aMnKUKbViYNab0QKka++hgs9mASE+2coVX+Il6Udefd38C
+u3ieKkg8e23UxNf26ovxZkGjXLOpR3DAjxy39B7kbSihsgR336dCBpdnUmdZpueNAWUp/ECjnB2
VLa4zOPmJGdBQEtBUxk8F+tcBTH6N5+AuBOwCF4UG/I/IItW02yP6lePCMGz0kUxJWCRIlAuSods
Lyqd+LbarDTETc1D2XRYpLIroVDPCCaJz9wCWc0pnftTa6xkaU0eGYkcT3hGXxwsvgok31ofHFx8
srCzmQJ1GMY1kNlWJxG+SS7pfZrnpLO2JeVupZyUceb9CRGhSiJdN5B8QXeF/eT99gLDkYozh75l
Lz328R/8ZUbLpWkwsBHyDA9XUtg6L/HJzCc31Oecof8V0ShZWwZYZt2KNA6XmKryax6fZYvCnDI4
CSOLQpBf2LowCg/sh9Dxj0dAQux/a4729JukePvhZP//Z0rDLPSS371yRL609al/uHMKI4v0x2I4
x8Ii4h67WGq2cPB+ZQQvL8ZxD1j3hAyH/J7hlJAexn7HXZmZ1474WV1LUkVTW/fNAl4LKtVYq/hF
4NAX4GRxS4joRPgQYQhhcz/To0opHv29dsO1GH/alz957erNhWRZ6DaqV7Bj0AzPAbFN6b7uEsgQ
9V0zLvr0kV7XQXpT2ZGPts9ndJpXnzoRENp4s0POL5mfDUSvPcQvzogxxhb27ABv8BZ+NTmCDnzQ
OiTk3z0d3BmKx7/AgoIUBlR2yRs1tciX3qGh6TaCAKIXu4HCFeZJjTDAald2R0ppyA81Aujl/zcS
LvcdPTwECOYCqjGkHYmFbHWWeKe8mjR57X5GAw1W6xuPlJVCUWxm9LEqHbYDTRHzHK/RQ7+J3Rxj
69nLwhJE5fnJe5hVsWmz4J9f9wxpyzrOx3LTPaNaGTXInFBktXesF3RWsi72NMKqEmLW6j+dVh82
6ld0bW2QedHVDehfygZ1YwRRIif+DFgZ5GXWRRtN4mUkArEuzZh2o97YyA0yi7OgYX2dntTK6IXC
47DDWm8l0Dy0CnDRAmjQyhGF2Djd5D8Wk0QEQ0Rda8F/3fUsHAJeG8WB8bbXX9afX9FLWlgsHQpN
4xkg5I903XFMeQaeOVSIbu/wUgCVtL06eFbTCL4/qeCGaWo1gqWLHTUUU/G77yj0ajHt22zINDF6
Y+ijrNKwXXfvwDJ5VxDS0QBVcB5COUVrsZykcJAb+rx8uujXCbmiXVcz4MdI3Rt1mjVIfpiQYKqO
IIljrmfKgaoNajtSpOCcfXvBKvyINI/jQ54f4Dl3VHkGQSRpjdomXc3nLa9I0IyNzC6mcNF/H0Fq
bW6jkjTMVfyP89nwLTmEB4auwOuMRZlqipyVV3lOjHwRfSgdeGIBTnyuZb/v4wbb2tq3pKVFfMWg
BV6H7fJZ8AfAFT5QkIjVHL152omW+pc/MJEk8NiMyfYH1JAK2PP0QkKKoSvgUdsKMyP2cLWSqoXb
CYB9p+eyaIJCcbyCX7dUCDiEW9ag7WEugAwFmaKI4jdHvj1p1+dSge+h1l842RQDGxix5GrjWlla
InLTJghshmLPd8ubetxnvkn40856ZKALUs9ALvKmN5pLr+tYMHmtSPH3f+EZDdQFfFUuBbZ90TJ8
5CpdZaMpybwq3L0HXRzWSKVl/pOux6ziE6bPFsje+ZyXIVDLgBdcIWRUysUBeMyDtvqQ6FXtw4KJ
8zNCqi2TACOQZIGmUGRG9fk4z0uS7LpMnXJh4kgPH8VEBrHkO0Cvjjs9LkeTGpj0GOzZC5x2MOu+
RWRkjBzNjCONcek1EOxxSem+6YG4gUHOFlG3aLvWWo1hsM9wVT3L5khezyFOQXRbixndVHprHxbt
0Bb/QMgN25Bn5M+Sz9Q6N1qz+t8AL+0+5ERLCF+keRqhHran/BeEzO/Jf0vblm2BXaPf8CT3GprT
v8jpboWo12rj6k1fXphoWMiiWnw6ZgQQl3+Ng3TQ5VaWNiCUdVqGPgnur8lh2oU7AoszBj/uRWOq
HyiR8SSYHIKle9An3bD3nWVfgmUbfEigFcjz1BCgcExglyEeZIMf0dJoiBLZwp1tr+cmAtJqGHQE
SW0jBI+ci6hefxYhHaNyWdC239H3n1HgZ/x/Rpjo4GnsIRhAQqkjZt5VqHJw0X6JZPi0mdswhx+D
THTM/PzIgWC/cYEHwfC4Meb/rwBlZtLSqcEJ9MI/ATiS8x3GUpG/yBQ/VAW5nv9WvFJsfxuNnir9
9gLaPQ9jkXhcUahbLmJULe97QzL/uy+scoKqOdqdzO2sEHCtrgKZprg89zeNn7zub5xRRv77h3UX
PnaRqr5CBMOlhQsxcfbJ/xg2QFBXpbwoW+VYAnMc9huePC2oqdnStzKl7sXn8g3J0T9gnzF/+014
qX7ibr3I/OIg1E2rPf8VFhMTi3ldsGuwcZDS/Pz0YU2IdnI/BSF6B7DMfK9OWGS7aDQpPGPG4rhQ
Y5aQGQjJ7uDEQFzZKTfrpF/joVlPindhJJn60lwoxCnQ4dZMyekRxenGYhPCHU3uZirKzJI2Qpnu
uE9il8+aPumxqLCsOVTypN2Pb4VW2uL13SftDHI6zDvlzMKe4EkDh/ChSY/uRyJ3Ot4u5Dmmbfw3
e8+lVh0dc7UewDu80ar7/6vKHJi9j0fCdbke+ov0DJOjHkPaN5E8C/zDVPLoCsgsEA3GPdgJ9GWS
NlkfNAUBBXqDGjv+XSqzsRK64S1J2g4eix0qPghiBGIDTGirQv4pkCZTieR4UglKsC16/VRG15OO
taTwNqoWv8/2nGOwve2sOMh1qOvuR67Mjee33QvK3R8LjPiQ5GWpeE5JhA9mzICw+omm3q5evv58
iVh/YtrElluRF2oz7ys27kCfX7rPIy5QEHNF8omSp2gS1fnYqRnywV1HmnMQ14pB/43hydujXgM9
E1oFoyF4YV9Bwwpl9Qfr3YRh5vCasQHjNrxFFDjEsHQs7NHbrDAtXzQvHet445k0czOU3i89Lh8k
vGd05SgnJOZe7c/HkBdP+dqpsdw/U7dlql4oD5xUBipF2NaCsEUu5bzH29vnnlK7Ua0pXZ5U1q2Y
iNxC5ZkpsBRd3XWu4OsjFu3SN5XlQ8sT/7wFg/x/5C7oSc1rBMSiZumPX/14chp7wsyndOsGq8nX
e53BtXlZoNTe3siyegBzsWdlHN6rKqK9E+Z/nBdNBrwgcTjeM8+c2QPykMvsClhWEetqGSUBHB6J
9pjrD3wJ3OZ3lG92VRzQ7BSjC1UARvKYHz2gQth+fCLXaYRiWs7wY76xb8+TrV/PXF6cAXNSX4T4
K0TNB++Ud0EySYm5+Gmy+FZWPFNo1TyjfybmMmyc2hYXpNHGYfq7QhiwiFWOpIQ5k4gFrCGgsP6t
k9jEaVFmKTevqVY2+Jsm7jgbqc1pyfGayN0GNjJLj2pgUaGMqDeVvbi5fRLlqXDapX4Hux7SrvoD
EVUHdSoetfsgaLiMcqnT9tCZUrWlrbngpY8Dw7BRRTr5/HmYTdqvVmGFCUKXdWdiZycympT5L3+c
Ni8gSm2Jdu8XH2LWYeNkWPkTPPWtjgSKVqhMOIbrFI8rra+J82bsqPgCC8Xrc7y065PFyVVWDfWX
oo93xLin6mubY+vXrN4RiQigz/5yWtp/s0aQiGSkP52nP+3Ewtfz6VFW6ujT8OKw+LJZpMuD2m0C
SOddfDPLZj9t+xGufHzZwBiFxN2HeN8j8VwfA/TC/9gPLGwnQi4nOyXRXi32qJqbxBMIgCx0QLBa
rhNxRxsAIhjasnxECETxeuQqNp02HRZlcQge9juRUw1QjCyaogbHrR+eR5Y3EwiJY6znl0mERRU3
Qv9s/gh7kmrpMRWuEZG4+u6l2oXwkjnN1XRB2HDskcq7OLKkmvwC5WANYQsR66/n1DwCnzFcsJ5z
EmoLvwawhJZMV8P0OpvdR13bXhKwRLSAauRF0XN6vPU4aEv3GQC6LJR22qxIzthYomKveZlIhn+0
dENaXKw/aRiLoGL/cJaQsJPrx9OUU5yDU5YyCHwxPqoRTgIJABjpQed+1FfoGMQ9oKXmeOXwA4fq
HQw0aA1Wj/JR8hC649ArMrHJUVn2UJEWUER2wNA5ApFBiObeb37fDqT5gxcRmInQ06xgtoy9LGoO
oyQ4rthgFVxjiVduuCgsHg6Fi/zs8OiEQ6Ey8rBXHXhVH86g8FS77TYyyHA+hJOClU+4Mj4yGoHk
+6Db4fiwR/tToaomaadrRhueC/uy6/j/6rDAH0sIZ0ND15q+REJi9l7MBGga25bOINx0A4JcFcyf
Dw+xbqDk9UrDw2Im5v6jF3ery1Kv17WUgmHA2vy/ZFMrC/DNZBflXUZ7yB3Hl0IHBVz82bRB3g5z
9RjCWXrgwic9aZDYmjBJK9WRd8Cohi58/cqAtmx1BQVabhmo+M5F5zOmKygxk1BFuw1OT4z+sKwv
9OXwnYnYJqyUG1F/nfLUbZTJqBEZplQbUdvJSCKDRlbMAeZdFTGoTRGQGIZRJ9Y+ztbVjEK5bdq/
FjsweQrrfelLlaDDNfUA+ZUFk5gL0BG4npKCLI9W+q5X2E00wybNmpL6u1Nh0+FeCQvi90DovhqV
28XxvUTCJWtqeP9g5mChlq+sL7MXjn2+MloPohrgxqWi+mXdD2Wb8uD6esH4GG7jyt4S7gCqwvmg
twevZiMWOpWcJrYkBolxwpWSq3wLxpKpaltfKn4Zt/qc6ezssReTEKXykRLrG7I+OKaEiDp66zaK
Iz8wbzTaFWI3Sh7PvQMap52YxL+cwR39PFgCUoqY7TJNOhPCWOLWv8mOqpq8vsFEBB/0Ane/6scf
cH6Cg8Rzfx5nNhqkVfJhNBJDHFoGWGoAF0IBczxFc31s6kLuKRxMafME3HY/EKr28k3KgdrPzSoX
gPIe5VPyelWwWb5bl2vHidH0Ug2hTWo8ePBzePCcjCjgysTYdLswIkvKYOaXHlyLtOsr1XTdlP+D
CTYQGD2zKxoHZdbKHVIK9djioJpp3O5NLu6nwYDfCYui6WrKNvMPOyhovV9PymJ7iu4cIlCfskCd
3MOtE4GvulTdHbBrF/ASgcJII3qGRa6k++OTYiX6Xa9FOkBuBMM7bRegXeuQOBJdabh2xRX6GP71
O+pQUHv7aWyYjjY4s7QZXXb2oijarhoqnZaPiwx+IJb3aj874rD57jNxHXtZXWW9mjxSZQRSov/l
6ZwiBiBylD53L3Kt4iYTChV7ONZmvbYzlishoWwUOHUhMtfV03gG8bRIZoP0u181HqQs4KEhBjx6
1ynKU7SnnGWcBCvSry64b2USwLbw88miX/y1ZbtPka9Y9XHOSNCjgnxcsMwH6vPxLpOiSzlB84It
D2/nnT2B/88KxKWlk9PkcVtL68xxRCVolvpA7djoZBymlLhBREQ2WZ7c3HM18WwWig0HwanDk5BU
svEaArbct9ZyWRkFXvFhW7Pu3wHBbp1H3vlcwGtdhuyjbjePz4n+v9j9jwvo/j0vrlht4lUyZFU+
FNW7d7Go0D6GN2DKJSNNTzW8tjPyeSItV6masFCkPEFjs/ZteCbbxNGyIF2jdoeTbs8Nxi/t1wW+
Qt7lArZaBm32J9784viBUybF1K4EN0SvPbNUbjeCOOutXx5hsdQjM561oi2rdjJ4krvUPg+tVUcw
ytqeCRnjL/Q0tQ9mVeKt8CvtmTBnnC7zuxttvjuDy4kryr/BCskli4dkrBCeoVzaXm0wCRL3s7bl
qrOiq1H7DxxXLBcDVpOvMN/t2KTg0m4rVW4xLkreX20IIKTXhrd6HDzjdV3F3YHqaf+0BG5HcH+h
qNf+mCf65194oBvmiMByzhb9ZKHhn9AQ/Z2uBOLv+cZQwisz9n8H+M6hhxUoYfWtu+xdpjFNJF2j
WV/9wPnWRj6mN6JvNqWt3rlwkQWSqqUBjIsQ4PJ2MtkwR/GpZAP2W8qLFF2bzf/t80b7Kvszd2l6
nL6DSWMEg9NX5wKjLYZaCGrKck1CepGxobjQoAYlntRVjsTiFtWpdu6WHaHmBWWuMgnTt0qYoNPe
epghCY3whYZjOB6/IsTyBJYrzSrwUwBg2IKX7Fi+uuVpAEaqdyBKcY+tv0t5rA1H/U2jQm//a0mP
1euT/5XNZIbAhzjVhAffgLQ6ZePCL6LlKoRkEou6D9Dmgh8gH+4ZFTzq1nRyo85q7gpHt3QIOZko
yPRCDIGYSYdjTR3VWnMu1T87Gah0X2Nwry3m92CsKuUTVdVsIfklxDlJu9fP4NXS9Rn1LSwIJvGY
WqW3gVaaYN2kNwtuZWP1jzHy8VFaPXzdwOsvatABJyIZ1Ei3GWNFWMzt3LInRlNopPLPLcTVm9io
7j4OIEiChrtTw8ZelO5t0aDupRlNBN61FC7oF57zMzCIDcmS/Q9XUWIRqPHvTAZiFCgOU6QWjniA
1tltKYLiKkkQ+uqVMou+uTktEKJSscg+NXqCrwsaR4DNgzA0bPrM16cbFpAAnx2ANtJmwdn5Yw2p
7ew3bsGdvxsq2/5EeREipUb2O4pOpCEtPM6yXGhDKffexTPwST/YrG5kjRFd995Kab7DU6aaNRcB
okdK6Ujhte+28Cq+6V8lRLyifEOQBc6m1dHnaw7XTRDEi9birV/Z6wEu5r1a+T+6xRg9jn696/AY
Ezz0pMKz2Jum8RRZcQILKIenJafmuY+pEMJKDCszQFSLvtOF7grfQ5L5m3zTJJXgnEtfFsA8zngH
xm0ig+0FVJXjTCyObB2SDM2hEUaEx77AA+rs0iOhv0MypP1WOlXlub+bqimLJmacgeC3u5j8Meu2
TNxp48TbIckuACadSHnzCBW2LWJGDZE5mAscPdH3Aow6k8fyH53xhiwX/YXy73R1/uVvCclUoysz
FlrseUuORpnLarPQTtFLFCgtz0NC8DXbZxXgxN9JfvCGv3I6VVM3F7ZPmRmW7lG5o6lPXx/ZZU5C
MQRilIYXHbavdOObmWPRbr4KS6kB9w50xyj60uHaDKc7vmn/oaunhNSGvI48O8QFKjiHQE6M3Imn
drJLd1kYSYrG7zQYwmXUuC27JRiD6n9eNqk8HJnv5DjvnyqYZc5OSLnXdF4n3Tb/aZidLoc8u+6v
nUqK4yIFX9aYXW210DaFQR1x8H5sYO7ZN0H7fGiQf6i1Kht/tFLbood93zbVxYDsbU6PmYZVFWSO
zYbn0efgyEbP1GnhwAr199vAI3EVDjRPuplcazh0sOtl5gI6hqBzpGka4QeXfvD1ed76ImHgic5d
04m5IRMw2Tu1UQN/g5cf5SJuDBDWCgZSnUU9Wn0z51tnOA3r/Jq02GmP/JbJBphM80n7e1/01gh8
4L85w7oR6+d77kALw3mbBbB3kAKoKhbshC1HFan1ocU8ybkkZuIa3AXx4JWlWyyqP845jDKMpgBv
IIIsR9E4vwBfgD+C8EZrS2GVgiupIp3QUyVrxXa+QTQWy56v0wcyImAyiPQvKjo4dQDLGvs/erdh
iMd2YZwkmoO35h7HJObRCztVcK9riL1i+Y8v2C0xzdK9m5Zl6X91WyQ1Ybi0cgkcV4wsHEIoZNqK
kLWWlVF6R73pMCDlqsk6huSq/xBfORkOgP8OY9nunDHVIGdBEPNmrN7zX7yL/c71PJKsXcEfxGtE
CZ69YpA95wCyFsiwvcm3kh+UVZXArPLFN9REyNqj7pL/3/ZsYyoTjGC4A1931PIS7IzD2AfoYUGe
Sm1rSJ/fcMUcTz2a8/LF4MCC9VbcMModqGlPoicQIaw/9bgQjiMg82NagTxQowcT0X09cq1h9f1m
C4HgEabKawaarm/LpAFXuy6Y89MU5WoycRCYlhUkEgmn2MM2/oYNQgdYF7W+6fv3dr5chpYcgp3J
ZJfwzwi9qZRk4KPO/LxkrINB44Rt1IA8aQgufwhn6hWwVmH0N+6aDlDO/3hNCOa17VHDpsoB9GRC
AYvbQGiRTxz/tigetm4/3EYGj702zArbVXGaZQBzzpEdWHUxz+2DQJdSSkk7DfEhiPAuXK/WM6Fy
oYchFCN/eUjUA6iGUR/dz825C3ksuMPdGo/N8r/9cqaQQ9bRcrmmiDuFPj9ZsQkVe5oUZXWah4Ft
Pr8Vcw1F/c9pd15/EQdv8PeS5ETmqnv+Qp+nEnoxv7uUP7HnqEQmOXm4zewRkXlTURmjSzoqsH7w
CPxMhES4wXqnC3sVTcN5XZBwj7XI/heqg9MAwMjOP1SjqtYi1/5P/bQ2XBtV4H7FYyt+bVHqH4te
W+nq1OoIKrU/UF7dG7y7W4QbYoHhaJ07yArlSM8KBB08bHOOrsvVVPcuOszWMDlqvlw7FXU3J57f
KohY9j8oRoWsa+1MmMIlXFgXUyZ7fX7BvzrXZ6QEOEgZksZotNcfhCpjWqRjszYg763SfcvDd8pb
gG02ypnHvW2ijNQ7Fm5Qh2eexPhwILDOel1T3EOx4VUzw8RhNlI3x7BvD9Q6schSsLuqqt/VtxW3
7xeyLbzPJ1ll+al1j2OghWoYV3LImKKlzNcrjfeKcx9jbIKDERHPCMzRtd/4LclK1s/LW/KwMIDn
6GvBbAlBriuxquRSMc+0AUr43rRFLI7rsP/hfW4U21x3dXOIAySDoC1SLYzRb+DABkb93OopYEAs
gVfKJ69AbDS3UuUZJ3oTqppMcYNo9vEgGv/Zs3zOqdVLwOsdnWkDxNAnfzQnDOe/L8S82Ic3W5hz
vQWbwGYBfBDivhVAsLQnr7BDogn1OeLhXW0LamD+4DO5uzDCCG6bX+vqcJbnNFVluR4rw962ImU8
oX986/UD6sxpbUf7JNCu0KPa9uBV7p728ZqLD9ysCv4msuI5hvsycSTrbpe7TpZk1AXjl/vZ43NE
IPhj0rHyvf6SGXlByPUSUS5RZomK6Pi3FEpWNnp/VN4hIBlcLGeupQFAKpkrmhihclex3vFLsnoO
j418Ser94Hc7wgljzmoC4KTvdwoqiZxzMrCxtNzmxE9a2GXwSuXUnR6IxHyM1Mh9UzSQppGT6eBW
7lPc+8fXema2IYWaPOk2/MGzlpIMG8Atlp00ZTfQXIhnjMpVwuHz4H4mhZpdwTmiZy5w57WGK6IZ
fJs1GH87mCs1m8HW7inN4gRU7P5dArH5OFl0GE5hfqpe8+sbeUXNmO/oOSI+9UzBxh7C/J0YziHb
gy6ekuh+SRzSx6R8pZllPBtvTY86bVYiRigy34jXF5ui4gGLwXWVH5X2DPYBEYIS1iU1r5/QMDhB
zZCw8+PIARccQRxb/Ah8ifaWko3Mp4imy8YZErNgYZlklRpxyt0/M9kkBEO8hibTJJE9yaw/ZDrX
ayZNFHq2t7pM01symzLEJ/fJG/i1JKyo8blvLG9QB0kBzn/uf0WyQmU//nfxme+31MhzeZnxstf8
SEIzbpT+AUdPdtgoG0lii0wf4DpJFotSaUxjJ2tRxdYdOFWfSwfLEHSZtv68jEVFnIZYD2ZTf28T
HpvkrwMR53rznq58yfRN79t0MpyUWga8B8e3dO4CBnYcUNh11I2nniNuW2PoAUWvH1iS17Q6xo//
FxnMo5vR+2SWJ4E964RcBlqxHouEiKLRzmpK4XXaNtoqKj+xW16AX00vciSgVNGqj3k82t5OBpWD
/XZqG4lAS/KgEmSOBUydE3I3mRKI6HcxZlTfUhVURptlWcKaRUWlurjWuRTxYe1+GI8P2bL+k5fS
0GTdrWYuq6S4Ub+zxbVg8qDmAHiGIonJCHKUnD5C62191xBXUtlBFndBhUsfBuPNgO3CQIJjg3g4
qtUAXTu9IkCJ0uy/3bKRDOYDqhj9rYWqKZ0sYLKFXehlX0gTK7Z7kwudP9LIImkv+sxEbUsG00Nn
Rv1+USMEGhcBgYGCjeme043e+WYZlSOLvi3vSxGWft4JUK8ljF66ug1Rn+fQ/eLOqxJmyguhehfO
l19uODSuJ5aRi+AbpvziS47en7oMA40my8RYsGZ7rEauGqtbjRPJEQjxy1+w8AYLF2K6oQVZpGc3
15F+HDvV8+I4H/WojdRWV0F14gdBbFZ8TBNwV/6VbTZva9L2oDaUdkda0QA3f4w4AkMZIaObt5MH
XJmsv8J+HtB6DgI0C9LsPYmaP9Pqo2cNr/obDExubJIRGU9IlA8prGg2Xic+A8x2Vo7MsGD6s2xI
kAGkr12R/qpS7LSJbitVviUs9I01oIWRpUoecw1rYFEu2EdRTYtLBus6pIblj2LPR8U8Bt5ZtMid
Bq4xsKQ5m4jXhLcEPSzDASRL6hvU/74iIkmMRKkqSNQv+6fy6tWmc7X00jKuelgkJ7wncla8+YK/
EjZ324naQM0GQoS/WeVXU4R9dCsE6VTBIb2JzWUVa+GuceI76GokyIzJ367gOXfiuLHsulRyCxcU
xDpdbZNmulz1YnQc6K3qAvAH8x9mnKTwPMrV1aBT11yh48c5pk5PgmaUTwLzoKiFbgMki78rjo1S
RzRUdXUTjFJRPeL6VavQ3+PcklAN6IBkbPBETVLbRoughUsXHURlN4O0iLmWurOvRnwQpY5SJqcY
orKN/xIbXU7/nkqaB89her0ElqaoSPM8Q8ikpzUpmbQ4wr1nxydG09beAxjjp/PKUTaDdoXl3tHF
sT8V0ZNaswL0dxEY0IRvgGVj7EGzgGft2O/nFISuO1wM5z46hMa/M3tjAEf1Box8vWY/4No4GFEu
NCeoL1Jkfnut241hlIKdYmoJ12uoBj1oxFczKYYOQo7fzvTIw1goVtiQ6U0my4U1f7cSitUTnAPr
StOa3ILgPhfET58XjlzeRtBXGoPK8vcCM5a0hOqC88uPrWsJ1arNO4M6zBSoWma5TVbFiuyy48I6
pbx9dY4741BZMtZ2iGhm9w6QBRo2/SpZ7QXWj/s9qaWlNyVGBzeMmPaapMAH8Vztw4CFU22bF8OJ
ijWa5f6Hb60jKC6URde9OYeq/X9vBTg66HMA7qF6S4F/p4S7Q4Z+/mITAsAxfi5tdeH8XrT6nQDl
23l4NOoCtV/P57pQenYUDiKqk0Ltl0XyonZpLQrgnIao7d0huBWifNbDB8l3AywLjUPncTvH3EF5
3RqgR1EgTD7P3sfneGp5bq3Oi5akyAHzQ8cJMTkjksDiFQBF5SuHlmM7UOpD6qnGD8JUAJrP+VV3
DtZIQSS04oKewPet3acrijvcAzZsXZf9bcwqWJDJ5sAtsC4tTp6NUR/N/Tovghi0fc6aTb8gzK9b
JeO8NrVEwpqdiNe1cDpGzzsBuVCRJ8rOSxGHNCYOlaFeK6Q3vnrZrg0mKLKeR6fbrsaBL06LCoj/
G0Jm23juA2Y0lkmipsOZPkxJueqsySNS3hyRvt6RIDxeJ1q5VDEtyFBFFVIB4cuenlO/W4peFhoB
B1DrezExRvsk2cYcg82O/ggD8dL5SwQNVQm0EK9JdNTw9V3Cw6swflkfhPB72tzR/GqVAEhYkZhe
j1FYoL5r+AO+/BFpyPM7tw2osgGpaSwYBGT7l0W8jz9wDAEbjPfZPG4cKSfVsJsbxcGrnGFuHPkA
/1JXxu4Bkih8dvM5SvSKVrWAJCv7CqJZJtIlfiFkuDvjZPt+ruSTqoI8FffXoHMHpJJxaQDJBcbV
/8LZqGXwDwvPerqvwoIUYwmhDGXkNMv1B615qhFd63HAHA0m3T7/IFAT7iiZAj6DJO6sbVNWLs56
h2WIDuXN4sQt3ae6s7X+3Bwxvxli7KTzRp9Tdd5EDVYI7kmRYpdrsI9/VrAzhCbm2xAmiRe/Q9LA
6K53MXzdDW9p31zE4UoG4iDR2x25Qc5nVhevshwwoInD1cVIW+h2lntd7IChKuWbfS7Yvj/8u5eF
S1sIZrPzojK4AiirNwLp9Llp7LjutZza+wD4x7kn8l3IA7IGceXeaKLhhldbGzE0PAsLjmoRWl6/
9Tez7T5OobfLb+sO1FG984sjsketgtcv/RCi/NeF9UbNTF33ACAUcq7OoMbd7ytzl7sMUpztgidw
AVCeKqS4w8nOA61RxesvAHpsjFBMM6LYTf3gp3wV9M+ynGgY1jMWxW6EdAkAGn5nnlfXsZg0FELr
Ik02L5qgJYxjRFZAQcGvRlrayplR2hKNvUVa9wRhAI/kZaSYGUm4csDyOI/Zo3HcJuzbbc1Y+4MU
rRqP0uHLLqlvsc58Utg5vlB1nKdzsqNqoRoaL/B/fPzWW6ezvDJFeI+zXTxPx9Jw4M55NzrFhVxd
QwTEIiB+mjbvkXS/WErR/4Ss62I96zuYS9gWKMcJcoiFMVhJnXgSdkcyr4jqyCZi65MzAieUu0Ww
YSGrC1q2Ohlq3VogWBaVl4M/1yPTyxDBUNPMWhVfFv5TibhXOyVle45E6y0gYx9FUDn/2nXixOCO
/pdoiDUSzr5d+vzmEhnDl8IZZbTD769MnfCf49qaTQVq2PGwxvaRXk8Ge+v++zf4wYlclU8TONEY
bEXKLX7388lyTiXtH93mTK9GlGmNN/iyvKEui5CnfzZ5hPnorfD+UN82+SkMXJ8ZIUW1fsQY54QR
KkdR/2WX8iGvz4alMIXe3vVVxfnPoCQR4KtG+gUvtBbAoUjZTZGjJBTcyOObyR2LVf7QeGkWuSE8
wtIfXiLBCK41OQ3MZs5bCKpMilZIUgizZijAcUWi2xBKkqWrAzAC+PT6xcvXi8ijwn0AQPpf2U4d
s3xkWe0a1iHc2WLnrZpUp9u/PmDEKYXw6AlHjWmr4TftN2WxU8In4bbcF9QOZMX4GQaRQDv8AuEy
T6N9gSOVdT0nF1zEk3eYjAM4EQOJ8k+aTwvPnn0qj6YJ9LkJa425aNlNR49+TAaJ4B2kkVfuJqD9
EwdnFQG2MNY0U/0JU68IrUs9xqGf55tg5mvWnkCDkxS14p2qj5MReTHu/HRVIRb/Q8fYfWXbc1vb
6j87lnZSnk1XER4ils82xbRfb0A3eh14RbtGQFfOJg4aW2OGL8CZ2J6HsU0KEvSUfrITx4uPECPX
/XBCsLs+yVeUdwYubESO2HzYK//H3pZ+F8SAql4cUkQF0OZlxTnAcVhNdUot+2Bgx7FapJgPD6yC
5sB0QY1R1bOAnwZuF+iX6N+uWPPwVPAJoJw9KnBWxbkplfTySgRxl1oLd5P+yiIAzGDrS57tzmvx
LeZMS+159eNhD2P8BybE3tscqp/dgmJZFiw0VIZ586vh391Br2m/P/qnMH5zsG63zx/wlXRDgkOm
nf/qDIp347uXRe4GosTXRrQnOTUfhN0eUVgdKwIjwNdECFwvaJsaqz74gfxkEzk6rA31XO3ccFfp
IH0KSEnVC9cbnBcZnKAgQ0ZouzVvkPlmtqOMhlcU+r8ZmvjFkOCGHwEqs7zl5ZyJWCfZgskSMFQt
MkR315fIW48Z0GGEReNnvbmiNNBHNPRI722Fb9tEES8RyoWB35lR7TOKzO9XM7vSHXKW7AJ2O1Yv
fCK3p2Jnpvc4lRuv2xX40m/mDMSDBovTrtIoxsQ/7rtsClJmgsBsIByjAUtqOD2HMnYDc/KvgwXY
gShxEPXqPEO2rJGWvXE90dO4alj8HslA3js+ainm+KtBP4u2c+zMettawgvy22gvjxp/2c5xz9qx
H6nl1GbT4Zc503oLjZDHo5BOCjXveE04j28OR5hZ/45FFZRTBgqSTdaP0JZrJxVq7DkNvObo5+jM
FkJaxsSDln9qQZ215IMvXaBijKep08dfTwspOXY4ylnTQfZbmNKL7kuq2GEcLVr2AyQsyQ5Sv+Fj
zptxOuOQJgM6oOYRzEYA4aJLp2EQy30IkuGyg5NpnTx417giaQC3Fz98mrJOzHn4Y71eR1pr3K9L
aXMEWWdq3xzX5qxGwUy4N9tl0igZFHsJxKKHair8KVYAN9Z8SVODbICc6ydjTrfzt1WMJGx0g2wh
UTKxaOtLN1eGoTNksEXbOvhT1UctJjUfmKNJCo93ox6o+xtv3oFisg1afQ3XC9Le8Ic0jsVREAvS
9JZMByE0Ah1KQ4IZ30GD7jasxMQM2FQLbPEUWS0Dit0zTmEVRWtgd7XVU4xtQU4C/qc76jWPzFow
vdY0z+6w2BBByHRvwHHKTrn79EoBE7GdvHovLqPFYgmrQejCqxmZ7USuZDYDgvmi4YWz6ZsuPA05
OX1zn1aIzlojmIdb/qzzsbeDcrmZL05rot6NZYlJC6APnqp18zS4yDdXmTSSFI62/GNpZWgkRpGA
x3bk+X1QmWcWUcq2GnC5+QGonZcQNRFekwnRM/v/jZ03yzmHp/+N2v93S/SwXVCOcTDikFKRuEf1
ks9faC+aQTPXFXFFiGCy15ggl1b0h0pOyPvGLfQUk3rSPm7JLrYzmIi7OrzuuYMdNidSW+R9k3rs
F6nCYANw/mSMExOpcWeQeoOJwK4JjSoSq6ETedxRVHHt9GuvGZAXk1Juh9T2+vfuEr0O0j9nDniA
Frp30DgJuhw6Iufrqu8caUrDUsM4HfxrWR1ATH55irnQtk3XVlUAu9fffngLrlSMTJvQR79er6j0
YJCUi4y87ppAzMmOKepkmHaFjQ5X5yC3jYAUt7Nx55+3UTdNtpIjLqn01ECC7j0C1vVqiCwIOVoR
P6e7qQFowxgsjJy6O0Bmz2KSfN+VDBf9B3GlavWzfkhR4aJ6cAJTHkPLRw5wDYR0/gjxx37RvRm2
ksH40bMwZHoRMn0L+R1giOVvjbwHEXQVMSnOmlwwFxOv/VgubNh7oGO3V4im7pekhRTqWvPoYae4
fdL5liSLE8skpytQTy3c4MF1gYridHtUOwYnf9sGu0QR6X6xYpVT3NJoFi8bqC+G1Vbe3MMFIvEW
ORRHghNAzPRQS7zpFRHcAFfW3nukK8fLOYAgnHBRoqXf+UXW3vZ7ZFD6VtwQQZSUwZXTT8UfZaQU
b11zk3bJ2YhkC7aci5zET/9dwKOgXDyomCAKqdSc0Ih6Al90SdLTPV4e78Sson5ZOn6fJbdmFzEK
LHMGKpe5LnEmYWuy1/jtMylcmFpWXHVQbvUaZib/VPbe5afwIcACTD74ADzmiNAr9kTTzNeMp7GJ
bE7FmpI+tnqA1+mrcoXheeVu/b3Nc3UWHBzxUhNYS+63AvE34BZ+mWMJvldOtvnY75RG0jC71W6h
suc4RVCJFEpwRScXrXvgCWKyBWJqI8yuajK4AbX15HCavgG/tl4/DffwkbqRJtJr3sItA4bd6FzC
TCq/J++a5oA4fLjchEh6NTdVKzEHYvTbbMm9s/hl0UlNVFL94Unizm0lvhJD2W9cdwXMW26Eirro
7+F9l6Re5YctMXyn5VjsLvl/lTqI8tb8CfRU5Hz4EdikXNlMWrQ3HBJGMHSrebDkCEcf2kKkyvFP
hqDlKROMrpR37u3oj+68z4JwPQtX9M/q7E3Y6lGwk2Gk9LpQWk7dCS9HCqMUTlYma6YNaXfbCbgI
0s1sDOp81u5Fibtu5U3RIYzNj0OoWzfy6XZjgto6IWOIMvVEb+JM8ViVp6I0MdyKxRz0enhHOtxw
SBrGfkR/dvC6CEzn6ggLO5XQgJxV4cc8v97vLTAbJcFaPuP47Q2FpVDAYVADmtupWAXDw75ezt45
ZPzADijPJma3xXrGYv0aILpriTUOBQatgz/lVGZTlabF2HAof+8V2/CBuyOZ2Ft0ZfO71q7SFIw6
o8JTp+eV5s21NbCTdvk7D2XyKmPNYfgpeeH0WFXY6TY+ujTPK4F0gYkzOWGuGaVpL6U6kQ4sDbG3
a9q62bI+ybvA83+CpWfRjyTlnSErAMlh5IIPiU6zBcvD2ElgUInyhHN+wZjdNwDQ5+OYYS0JfZHr
sEinoClodyuijzc/S3a3Onx6DvzF0gv18Y4QlDrnDxr1pLjm5uRAZ0jasnfnb2yhnzH735xgQBpe
S2uRZ6ipg+ZrMGOzR7D7t5WNBzhMSoyqTgm1p10M22dSo0MVpWYCElRJ1acZ7a+LJ0tekfJoJDQb
h/sUmeWd0vNamS8loJ08nDmpc/hN07dBWfq/zmiUmhQONaV3IFaAmZiPOncz0JVaQxMgRxQ6bZj2
naCGA0ysh8GxqZ8YdzT9K/V37/ANHbEH6Ync8WSdKA07POW4SD5WYWrdi9TVp31ZdUF17oMWuP9H
eO3AZVyg5ddm6R8+iQyuB6EwiHgriHG97WSdcPtM+GHnIoKQcvpt/LaRV3H+opuAFuPRzV0/mk+4
G75+pyQjFTsSpBVw7hu8jlAPkDzSDnQ9BFNHe42F91Fy8EELJMNOpQiJhYRKBBJckUlDNmNUud4r
5udkD2R91j3wseKm0jPYGF1xMB5Da5zl7SkHfCyv68Cf9NAwhqpQNJBAWexfmpfnIdFNCkJgOsMl
u72v9B3EgoYL4Z47za1mW3bvDxL4YzyK5XL266rKgzKkmpYP/RCw1aH+XOtSsauvAOc1ugT5yeRy
PDO+o0cw660zxWPj1BVyfZUML/0aZAreYqL23/TtsnqxQqwS050jpHSgVh4VRMZLKgNTclS13CR1
sUcqxNI6qulB0EWmH74vm7WPN+EkMWyYFgM55Hu/Qmc5OjP2UIge9t4JLne1m1U50pQVkfzETy2H
elN0TUDwfSCXe5p9N/8SBhGkUBGT7oDBG7+alt5wbEcrm4ATCQHD+dRS0IGc2vjx8TARypn9yxiA
XJUgazKq7RogiyHgPrLL2+O3bm2ejTTdVnPLwP9lLVmxozmW99vw0AekabEBywqWdYr1VCjAUvxx
F1IQ4iedq58hvXNfh7J23nNYsx2Mf+UIcsMm9zQfsOxXZrsxHLu7YeaIPtFhVN6NlT16SZgC5O1D
/Arqlb/Iwhka6AWrXfxYhnTAwBCGKWf1Yc1qXZjeDKc7PJ2qY8cDtIpR3Gk2CVumSoTlEn7pqzFT
pXbyTdNr6TdKm7edGpzsglHnOMdKf+fXGDcd/XGSBOEsuThEBOzORVpb20Kg7eHNwT/uw6zHFZZd
z2NGSBeoGs0aZ7dIXYwbe07cQZXFKbETjbLy3jGlxbQyY2zDEGRWTiOTqAScWgkm6e+R6a0t/nMT
hXouxPwTZModcA/mSW9AREJjEhMh8ukdFBwau0sEyUg0fj7GzSjmMbXfHhU++xD/5+Ptz8Pn/qFC
kxyJGRaLflPfBkRvsYNOMn8a4cy/SqlJtsQ67lFfszNdzyjnqsYCIHIt6rzVQOQVqTHr3/YE9/CU
mfNVE7C3OgTHjr8WkDzuf2+19D40AsshSMyX5jFZzXr62SNRSDapI17U3tDYZioFWGENofzJRkhD
XKk6PJYM4LcR1EEDdInIN663gBBWP7BSs+bBtN4bkf/DeVBgSX6mzctKc2OG0VgBX7jMjOR6uRRN
DAGPaFTwM4SODhlLtO41dik8Y9nvNKgz99rjpNHJmFDZlLLrBgNOBCPSXRiLVMY++Tqbek6HvPfc
iytmbxMphW7mH8YJgKK2bcFUZ0t9VxrATVcQoSrhlaG+jSzBkBd5xI+ybzrHJrDYI5Fe9PsR7FJI
TrFgwxrwJrYr3lV5nGT743Ib+yXFxHfkT7zYMKnnqa0wOk/aFxoyepXTGhUGiP+tykgAoeJFo5Fy
Cz7LoAvSWCDdZ4H15xZljtxy9hUAEnZs+dhreyH0n4pzkqkEa8hIjHq6J+W0kXFGwEMuE+ft0Wzl
0gaq9Bq77h1bb64rtCFh6OgTvO18bGE3aDdUQkSHsrvPnJzye/m3d9fKPH4w2VthPzJSi/DIoaGx
3Poy5G/tsZx2nU48wxVC5BmBZMF1A3XilMF+D0yZYTN3rsBKhUGv2+vqSgAoErVMTWGuXn7uY69I
WhaNTpxd222uHTdv3poyWkAlUHClZ0KEP1HK2P5Ifxo936AoMEyqvOCPl3r3QtLerC6vABuEUfyY
6nQxhRj97XbiWTCFnBqxypUB3medg1WHEa1ABZhFWInFeRk8abmk5/BdUyg4vir0APdwDlR6qi2R
0saQx5+SXLo7Igarc5hL58CKHHzVJW1aCNfF/9WTHRkkzuln/DLedRdz5b4KGJcJCE9lQIqZxwGx
jX7pW0OvDyI1vF5Q2f0rk+B3dCoTs4lS+fnyBjXxtFlQtD3qgvFb7U9n65sP85Q7a7yjoeHTdT35
VrFuyR5HTsVi2ASKQ4ljdZTc7zpv01DvqSqUE2X4XCGp3FbBaXcHqmJQodTncxTB36sgHvUC9SvD
GfgmUvGlnUTx/qk40PvkJjsUn5XLdRMufxpnU8d9veSMxFpk9CTTa2PVUExyVYTIXMQSWmRQnNCu
3RarnCdvN7wXSPz7hg0UoyDtZaRVbD3DzI/uYduP7tuliCWVcpNFErkaaNdh1bWMbanYL/JKghqj
ztwK49rpRaj1F0OzzZekvJb2+dEjptc2VoUk4S4FrqfBFNjFA6t2RkV+PGlpSYX8hOhDAvITBLIy
qWkaGk5jJMKtFdLcROMUkD0hT1eYVZ+9O2HYm4cyuXU0q0PxmJAYq99ecjueZq5p5R8ExcgxZp+V
NZZ43fx7qJRNdTOLQ93+7XU2BYHnge5WVwPdti/0oKHMaS+e2X0lGmHLN0fuFDowNiQ9Lq4LKPRx
gBox0xUydysA5jlWKTym0iH1qiXZxMysUjY6NNMFQ6aH5Gkg0XZq1MXzwKilfb8ZBrBarwsWQ5Lk
MnuqH/fRG1Kvpf1QkMdGfo2g7PSi9Dd9jbjMpLCZA5M7KLpoZOYhQX6Itsu0Rcrz4yVb1UHrldYl
/QLMj9gkBauv/Nlw4tF64BmHEB5Ty/YK5AADO11PU6J9gISVkqAlNmND4wS9UftrPvafr+bw8OXz
7xMZBDU7KA8bYEFwS0FGur0Bwr8CzkyJAcXh5HdgLDemwlPVcrWjJXyvDd04GEZzs0S+3GCQkxRa
HsywX1qON7M+x+dzLwSRLO45zaiIALVowXg1sFh5oxL6hYsC6BPsh5YLyWJD/nI2FYLDr7RZWJ7/
u9nT9mG7d6R7RDnw8jRKYe1rWhRm07/SQG+nlf1LPOiOUZvdMo6s3OI7CitR+iAWRnb6tmnsDNAm
dAzZA7FvCGAhdZL5xzbtgI/gfNq4OgClFWEtXss9Ys+vRmGKoBkeMNXhKX1zeOghJJlTTkC0uVBI
oz130pBN1lzZFi3IeNxEYZgiuMi4d2IMk1QN8CEa0ZZBd7aUIlU0BuQAxDHVOmmQTlOdahHwt3iy
blHkmt7dMW3pplZddSHsETvrBKMF0zV4nB1iZxc4frVBkXSbx/neG/TjeZrlCNsJj01HQjRKoXj8
dEe7TySUtIx809GJfD/EbH185gmtEA5n7nOEw8xEpX4mbw2EJMP2LBe8ozwI0kHALImO+YWte5OE
6RDPqM6qslD2JfsHrApgnZA/FB2OFMbkq0TdLqK+GUDBDJwe4PQ68uc4AAMHK0QV72FUzBHHa9L/
dHqd3sd3FsgPcv/B/spXeVjxOsN+WfKfLkODncgLCE9O/pbefDyV/6hrbLgO2jltXYvdR+a/mXWY
Nuubhi1Pkb+QWGxD7gxpMT5I+MlV3hIVDFGEt/ee+fx9qZlGmqse/sFRkKE/w8z7Wip+TqDNU4YL
M9Ye6euCVy6YUlx+5sy9IgaOAPq8vUiPKiN6CtczylCxUNvHwJTsBv/UDGNZQBevxHg6MKZVLIDG
fCJm2ucjWBFbBQ23ZxMktTNRG5PCjrVlE2LefI80kD7s7mYusmJTTSOUrVcQjrAolg/6Pv1Dptg+
eHvYwb3XWJbadqHmSy9oZwJLpAGmMS/cRp6mETuyUMdt2FuRtsVr6Ps5cazrAduZ7Iz+Nv1zW0dI
6F0/4De6ECKl33ycy/48zwGW74UbES78AgseGbcvzFBsasD7qk3iZiwugb4HKkWncBqDN3tEqobA
Q8LvyCJ2bpBZRSVeQ2dBEnCal5F+Qv7SU/2ZNVRhP2CAtdq5mU9tQizdccICSKfOASZxlvzPj8a0
hiz5GXhquCDGI0uxkxybOb/RJIRF28s7xCdU7SLLXIc2i2namMM+JRS+lMjEY3dboUZl2z/uyR2J
2cL3PvLxdaSDbuiE57VKaw6IYdUzGt3bWvK04WFMJVAl2c3tUFm1Ysp2ZfIpMknM9or+FT8QvzmS
DzcspJSJtO7of1A1IE2h2Fu2UYbb6tR5TiAeEWRykHOjTfdOtlCoFQkNY4LTVN1IPr7WAArC7Bgs
A+W7QIcFTvJSkR5YLbTqLoHliAjCS3PPjhrmLjDCI8cI+tlXSH9cHYJHKWuiK+wKKRu4DuGkt6JV
1UYEWQNovT1CLvIcinjyn2MsI0EmTakJprPxzTDF9OSPzBFanwwc/nc49Cmhh4PzLEKMnlm0LUoh
bkIo/jlft9Aumr5kCEcO8UE8H8tJVkBa2ulz4MXyxKVBkq98jVtHqkxQrC8T7inEcCvCyiegkB1B
YEi0ziNwpRvJPq5RFoyAGxhc3VSngmuy8ca3RqdySue9YkNtuNVoJK29xs6cfXLzbUopoELcO72A
URdPNJTqZOQB1jH30kkjsZudhhBehzhS7b/gfrM2KD/NN+nRqRDP2Ivx1qAI+fb8CiTkXG7aJI2g
jFhvPzXNrE9Uy2dYEPHggGGYq4Br1MR+5qTLYy2ZEGJhjlRW4Ot9XqUPctGtshVWO1iODULnqsOC
x64T2hVXq9qkk9CUNvEq7uwy1l/26SNIXR9euwkGkO0RfQLLkwrcYZGLgyIZ4hRznryrvLH4Ggsn
ObmN4aQ9HeylR04H6kf5vAJJhP9P+7XzCWpRzxPAGbMayDZTv51ksiHCSxA5z69U4zwS20cuviRL
gCH2UPTULHLByCWg8zsyAxpML+fSk5Xc/Bie5QR9TGtv7C7j6Qzedmnn6D+LhZ/97gRHCnuw7faM
2rwpymN5ljlA9+N0A9a4AONuO6FKDuKWw9vs9xslZx06BhNUWZ78ZtkB7O0WlSJZ1dwRtPq/Rz6e
uY/W2GokKyFcAsQh0EkVoY3UyJEeieocvh6kbg4iKM3E3HWoUHKdjHNLT6YFmbV8Qlo2r+Mi92la
6GjSX7es0BNm5czgr57S1tGI4GJZzXIaRHenv/trN7kntJsmYeQS5Qr5fiIzlm/IarwtICoF/hpx
9gxgBt4gw3olECEawZnK0qUrGkJ4mCtOkMkjO5z6GqhAdNaDT5jU/SWfXlTdj0s9CXBCm9QPcadR
rHyimmJbDCblf5Te1Vgs9wr8Z/WvHB7kNlJ9e2VZEgJ6gE1z2pCi/fNXLH+Mb9ioQu3uMtp7PeEx
gyTue7ynnAymrSCl5iI2RZdHSM0vqArc1WVyCg0DSTd2FoUGknM3tZ0PZ9EAPz7uz5HamSNc/xJL
03PLovkSnZc0IMllWkzGs+KsbZXkQhDbkwRKgxX6s9usVI2qgiAOHEzgckZCfyufHqj8RtO4IwBo
kE5W8Fen6FloffoNt2Cr2SUgxnSTqxnGCo4b5ZGWFFZENjqYFVdtKRyd8eKFwKpG3w+rknf09YaD
FJW7X7g5pl9ItOVs8HXb6K68McjNkOZy6kVoYhMYlIl3NOXKmA909ywAeatBPpS6GkbPYqZVBVSB
XWuGm7/3vmPHISeOvxqsPL5oNpYF7Br+a/FWRSQsJyGmQfA16PaYIzi5VyUyGth9wQ6Gsk82uR8s
mRjvfWDYQM9VdWyyx3X3eIlLtEfz+9dDkFATirLGPS80WM3zmJZ2z1xc/acyh1V9QBMjC97i7YZL
TaRPxb5LSE0D7M0+Ejcsx0torXJpOU1k6WGCZVMYiMrGNlK46tmke06CQ3qnBCDST7ouUUALFaxB
TCJu9Dd+kw30xsKigZNVGD9kXfOa+L2gbkDNSOt9tuoIde8D+UHprbkCE+HhRhtWUfDp6UMHvYjp
6x6Jk1hNjejZ5VtKwkbd0OupZ7Cf7d61AeAM5tFz3QRUimvg6AKr7u+u1QWRanc56W37vZzXSBLe
aTwrTpt6/xAhXZdlJMNLD567ncS9nzNkE9/njJG3WhtkL8+t+sADR6QSZ6bswC+e8LgAxaS8Wi7f
JhAYHPzn5UpOp5AhddH1jNygjWWfzWzb88g5yuJSbM5ixG/xFG07JpGmJ8z6gXl1NYIcFKCSgFI+
QRGCindZTsqlMtOKpAXFwAjL14RKvJTvINd46cYEpDLMqvUoOhA/4zmB4G+Tk706YcpAuP9Ihc+c
+MD6uu7wQ2IKS2yEjAwpdpvE++hG4jnQW7DbA695EZMfBIV9Y6X/fQHKdxVaui9VbfG0uftZodJz
X9wBbTN6/7SjhghfeVW3GudmECIOeFOAW163X4S8ZRzyu8Rw2ATQgFUkCIHD+i64VeYGTZlQ2vKG
DEA+i/rAsGJ+BICxlijHyK3ICeuNTMSY5pP2IFdpEWvOsQIrPVKdZ6Z0AE/WKIvPMyQqaIHMQ1rX
nWsH96ml2EedGWwBTQbhsDrDTpwelwLWvbCJLpgMlzB/BY7BHbuVYHgAfA3akX4meNSPzPXdNX3k
XsyKFllijMiXYGhtSqa1MyIykrYdKbhodX6iRo7Q0hY7UPWDtEYdR6j1M6bHg1jW1sfqZhIK6BUf
ohfifgBqhHFRYeqsoq2FNMC8zo6QM3UjArzNMjk7q2DRPtovbWOjED9Poc6AGKeoKFOiG8ZwpblD
onGomApoOkThAQolZvpNNC+HGaV/zCfzhf7nvrw6hPgSbXs3TcB6ggsrFfMC/W/d4uVh3V6R3oO7
EwAPxY7mNJ78/gpiBKdRuu3kAJ9eH/np9e8K3x4NcC7dqBbMGHy2iGHowSWuV/XLccRLtGewZjKo
TCBG7gL5hFgMySNcKFg5sMNXFnphj2QIwlXXfSA3YEsVapNCe+itOBFagnM9OxeHeLy1AxDcuCre
Wy7N2Wc0JLK/hGJKxAvDXbAA4mlEEifaNagTK7WLo13OIhpiKuX2vjNq0qY862i8ZsSi/KvRlazk
cqItxqilip41LwXlserpctBpOvj2SV1+y6KXTDLa4Z+ig8PIDYPJkZq+HFKuq+Im5lngoFaWW9KH
1FIlGBgHDCPeyWXj+k1pXOJJy4MinamMaWBuLRk7qI0M8McMvARQZ50sSqU3RCnzJKI6dH02/nN1
/VJeorVUKt5nvcUShFscqtpBMd11w2PfFWB591C6iiHsHRAcoHURUzXesRfjWRDzIVdPCCIWsiOg
AlXymFyKjHwn0A+lKkDdlYxM2J6JIRTtW4g01S6mWbqC7pDlsAUspkrSCL85R8HpKgOPtJCU1twv
Q0pUPYnsyQ+UHxPvwmap1zfgF9p+GkQCInseZNAn7sKKQBCS1bbTVK8QJqwRaBGmKw8SvqovaGIn
bcvF/ju3fS0f1Wde1k6F1R1uhhx0ATevUtnP+dMGb6Lc6Hml43GmSfMKizXs3qdrj9KyZMtkTy5d
lc9P3VRwVe7AGggaECejkumeSxVZzpI8lDD+ekFbm/pUwdtekyt/rxhtfBvzAtwJ3MJZkIYwI/NI
vMn8WZNhPcJHMjDC1nq30wW8dgHqJ6OJ019IOI2TjRxexUdY0pLw57GZ7X/nMQfr0/2Xkjzuc3ME
pBgvBDy2vQJDuZdUmrtUHt5Rd5RZjnf+hvMx5rUh8wtc73b9CuqCwZMIofZ6Ry9ctAfVaC599PCL
vtSS0sD06NTW8+nEgT3OhuwnwA9tY3C/I0+gbzuWXDgFkls3g8LxCDUwxsEGj82KfylYtV3gh6lX
tIYWATtwigIub4r+q2MMYILEWNCbrSVPv1lAoRqwOGJudsR+eY7sF0jLzgE2acRpUXWKfG0rgjRT
sCblpk0END885jrsG9pbU81i2slg1Jk/7nRCQZzDl0BI92nIuFt+pWg+K56OhOwj2I+Cv4fTm/jp
LD2dhddArhlSfFeUCmaYt84wnmw8Iy5najCKkAKCdAuTlylT1RCerp0jCaefcAFQXstraGTTaNff
O+kc9HnssPrr7vBcjOVkEIpVAEtIvSLYKLIOKYxsYMAP7WbmhmQrJR1NsB/4by03eLF84VHfuuB9
LYe5mqBCLWte2pWVgpoOJhsDn6nt4YBiBwUz46tdDXlo5XTzvIhMdVPoHraj15fUZ5ePg1V0P5KS
WWbAcOmwtsVebDy1OLLM9JS8FMaaKwB4QZ3M9Eo4DVQSKaq4cDA3XfhtZHoGQxhgyV5jbr9BMY+N
ojsrELTcHEV9LtyI9G3o1Ah+vgUOFio9w21rISFKh0QfDYyMtTLhU7ExPeff+EFmAj+dAZP1x5Vb
WISV8+YVkjXGt7/JQid3vRefyNQNSV6ncx15DNyK5+MoM4GOviGl64gKwRtDNfxCgH/pQD0OdivQ
UJ3/nimXMZK7qANk298+eW9aPYCEdYF2APbOtwH7zWoCu7/ESYd9HHnO8yBaO0FFy+mCT5PDP11R
6mhjKQVVaTJRUuuKihJaUsMC7FdmI7BDk4Sdm0PJFJ/E2Z4iDnHXdXEuAmFr8tcXo9tp0V8xpssU
hpDqGTl5Qv4qbSTpEZI7nRTeauv7ONMhFfgFXmC9a41ob93L7gTmek2mh26MQd/rlb1CUJkvYkXK
UXf6H5UCfzCic8OArIDti2fIxrOMXNQYsH9brkYnMjR4aRX9en5V3iMSPz8YUlmAbJD/X0NylnaH
mFEFduswhrsjs66cFz2Z8/LrPCaIhlsmwFvMtnNCBBhtYA9Rmx9qd2bzg6DjDk561Bn8UMCJECIp
4UcOMEBQ8Z8GOtYXU4bN6SD1622dp4vaCiMRbehzCFJzSpyZGxByoi/ES7PeIQB5wJDHENycCIW6
3/TKP8MZwBaegAxEZVoEtNFzx7Upo/9JDPVgFLL0IFnVkwBknNCsL20bENtjoE1xsNCbPFx5/iOC
keGiL59P0+d5KUYZeDEehzhYAF9AhdB0eUg3CvrlNdm61xwRYRolM7wbCDV+sw69cwsISEuHaFsc
Gr3l4QWWWl0kx5NopsinALXatA1fdzjRdkcTnxKiinc3EUddX6GmVX0glUPBwjDKhED4VRZF2+sj
Dl64rFIRyWmIycyYFfdislDfPBugNO1UxgA5q6H3Yflbq3GIWl0mPdPy7cUMlywoOlfmxp14loKX
+hEYyjGer2s4obrrF8LlcxrVsiz2ntpiIopmVMdbPhAg6wVjA1D2sDd5uxSkDVBG3QJX1uu+bDsq
KKRin7LIQXksZA2g7ybtCC8IZMA8gKVGxl+R1ryuDUhFutDuOxa0E23EklnV3u/cquyG1Kb5N8+I
l1aKvS7czfjqEVgxJ+B9f403TDp13qBAKquMTdMrknq29kXahqjk8XfQ+mO3YU6QY0Fo8mojSNX1
1SsMg0AjIviS1IUjJqKnIXn+Z+rcXW3LaewrfL+UyO8MfmvRTzt9km9+b0cdHNQrBThAGdbJG0gN
gblJwa1zIofN+TGuGfwD1Cap4J6gtcLUvbTCFM0M22GDEbZq1yxf1nsv7z+x9F4dCmtP6fSNR4N+
cItiDDs7wTZzVrZeV8tMoJB+VsUl5t0gsJoJfhGt9SUCqSVRhSMXsu/FvmzFhYXoy5BCKKF7lO6Y
80RwfbExua1SZvHrnHKNB6rLH7pdVpakrtzHdp7dgas7Tc85ThpZywjJVJ/SpJeRvtWw863uHcWp
/MP5eA/o3ZRxTL0Sy7DG6RhaA4NnYJe0ryVfmbxH/uy77VG5Fw1PLtaGVFi4f0KbBX2AqJLvRoW6
SK1G9F//UzFeyk1IMf2hTioK5m96wJXDERfzejaDgXLVLtPp3uLs79iiAPm3Z61HS7FXuQ3tJGwo
8cICotXHdG4gjf52qxq5Zx3rQ/cxehVrsWE7tzcKfOou80WVrAbJ8xijASBG5OhKHlToiEZ1X3zY
UpAlX2UAggIWm3Fcuvfnu+TWrmxJPluaBpOZEyvin7l0YNnKKN3El9dWa6hk8emmHJozbuTB3Hya
OkmjzJ6Wsjt56PevJIqlZ9lJAY1ck8cK0D2+oAMF8fIx3SAUJjvhq089EMdtey4tTXRgPECVVjmr
KrvO6bJYjXBGFOgU6s63KyXpOXjdOHHSbYTpro9sN4AIQEldRy9AExWHKafHLRPiz0qqCeW69XrE
cT+jMm1IvCOPtt/Z35Z/WL/UMhxFPYJD4xJLv17GZLYkIuse2iQrWXmvJvyQD36AEWxjogFunXfR
I7s/E5mtr72USPqOQuHeyAJocXE2pXr8DO09oMWhB4OKNCjahCuQtfyXQPGsRuxXWJb8gwR3zXTO
xxBwS8qLJyDd2y4KLMKD/OdykLpOxxxbS7IEdAWS8OG5cwWr+mGCxai7gdK38eR1T0CDMjGAKJLm
cQB4sbKoePVok6zAbVT9EO36ytrt9i3xAwXTWZH+YJGnwPgmy5UxHSytK9PFi7cam99RDhjiVm62
9ZltvfR7eUXMwN55iea0damLCNnoTojAXuQkXnG/WiuVmYTixAZA9ERx/rBYkd5EMe8UqTk1bCuc
mNNJtGatV2GQrgiqwbK7CWEOpO3w5JtVn89yAlcUo2wuvmde9Etiz3m1DphK0BL1P8qZz7Ruzw93
1XM4hoDPLJbv/IYDGAXyUZNimG941pWVGm3qZKDTj2eUNWbmhJt/SfEicowcrowaus6EXsVXOFiH
QUf7IadyvE3GbAjG7+T8O66YxTps+mEWr+qqEdezjC7Xkp46QEnE467Mk+HTYp3kqN3Fm+uZaxTO
6AOlMFl9RHfcTGHK12I45WEtNtLLdEyrlNYM25IgqyyKfx56ogy0mZmLJoOLdtQq1LT2TkQZI1fz
Wn7an9uFaAYcVtkinVvVbOX+I/rUuKY5Mf5dvNGdZsoCK0ymSjLhDOHKDl4Mne6xUdU5fqQaThib
bKiyFw9JGQky21sMFEYqglXp47ednsMBwASfcutoPHtVBx1GkGQTtyHWFCQKJJ/T7vyOWIRsuUm8
Ls9kqNlSNIDr/HGzcoqVqRcNWAkbPN0HSmNa20x3cbyc0g5MXCTMiSrJndzLJGaKbJZzmh9Cnpa5
nqKZVnh90bAjz80yLQTzj9jOkcNkAdzkh/nTvOTFzVb2VSdhMcgEtFDvM8pcD1bUtaBvp72kQhzm
+mKJTIrr7zDLgogPb8FuwakycF8QPLkuwjJV8kuOEuGz8DIIShYPP3gFRia4ercdybjxt8sRDGEv
v7Hm4SHoP8TMJxEeQ7SCSZuE4dYUXO/oMjnYyBhECyFh4pXmF9Z4q7ehIh6s41zcLHs6FgEb/RV3
+ZcPRlRv2r51H9Z86dGRZp2OCaoiLUPqAkPR6AdC4HSKvidI7uxDDoezNJBuROK6iq8uMX59jVn1
ZINEDDWri2nSzCV4y9hPCXZDZTDKsz3SIJTBDp3768MUZ0o1U1EyYHTPoe/T0EYrMP5/GDQO9Eca
wvU0wdK9dXxstsFHOcHdTRzp98uxN1qv4zxdjo8vLggQIxcwUD8sleRUAgXKMJoq4jJuoTN2LIZ+
KTPJVdjGXYn4l6NAMOJgVnWaJDBfC3LKU2iw1cGyE7hvHEo1Nfc+mJUMMTgaPRYmIXC+TiyHj9P6
PtJUGN9+pX4kY4U1TbYTlUUzWXoY4bT8HmxfGpE/8Xypdb4G5cFJKG21VvZD+0hDQwT3sKphKRDK
3dHb3vkS+ZlKf98O2NJhXY8qsUGzB9PRLxt4CQZbQxnv/6vef+CqEZupCG47oGFp4clTfDmxaJzU
vIjybNfKBPe/iSW94u+lvzBddu9cOZf/D2IvP/5f2CX24xC6CBKUheY9Vw2yRJT8N8llfdNjbDu8
+/6B/gN1hkUNbWMYw898dY4ZIrKcEfEnJ8ivQ4nE0wt88lDTZ9EouCXKjBNh0iL9/DQe0t3XUNgI
Zd/azxCHANEPMc8pedInaT9k8Xv5VCE9YDnMkxQ4IKzoiLjhhouCxLk8u6Dgqn+t4KUSViQgwk3y
BgMpf2MBndV6+rYYtyUENK6dac9a30tW217BTpm4d2xdJ+J62Xaiesc+jCaK3G3RXchbEKrjTCqe
AFAJWFL7vnohlOjUACj4UoEonXMuHAonjae3MuNBB/ArfbDuU1DczJ0+sGidq4o+eLJBCjTQzEVV
MhI39mIflbwCKI6OoOAS3D7JIYSXpLZRSrlmrg+QkURH5vGsMEnRtzq232wxEPJt017VU3zcHOdP
lAxf1sCgDVakO2CCVWtYNhVRAz4/AVz7YdvR/mnojFdAT+OvwHQS1Fh/Iz9y1PywuLW2xJOHeS2+
R1D1ca/3Qgxzhc3V5oUJDqvRFJeT8mtP7TOPGQEjuHpSBWm4NoEx1fXinRb9FoRC3z+cJIN2h24d
LvwZ3GnD/Tg5vFd5dV5z+3L5rs3/hWqmCtk8LSwXfvLxgYVxDVjQ+F/0oVKALJAwk6bf9JbTU7p4
lgoMpOgEYdt8Lt281J4mhsh0/0DXR7YIaTinn9NxfNTN5LBVvQdJxr9m4RKp28osiNVLb/emiHFQ
TZvBwVpEQyFsc2ZtB5gn09v8t8fY+nThodhBH9Cp0fsYLVOZFpwmULIgEzwcWICLUOrO6xT2C6ql
oEDL37ClO8U0nnI7LbeSk5uFlD1BthjOITQfWxyvPHK22gtb5/IDS2xj9q6oK31H7Opxabq4wveU
wBKswzBOIN/YE+2aI8dz1a6YmFDEXYzU/J6il3ijtqemEgiSnNbqzLg7y6iVygUn/XMiqA7NXC38
1RyH5h9lzhhLK6lUihK6FvQiQLZ5mh2cGV6GmAkqkymPdUuhbsxk1M9syuxFfXxBQNhr5cQKh/xm
EKlRaBXXlRSRldreN5VC/L87CVrNiGwsRg17SkVlCI7SFGNQjPFuaSJ7Y2GJorfwoO9m2PEmyhSJ
+hXruZRKp2Fh29T2NlOUtT4UXPgoB1mXSY20xaV4tq1qlrbL8M2+nd8yZIoS1w4/pD+u7PgOUud2
N1LAVrhIOtq+0la9F3LnCL7vXoEsKsaxuOZ13tA1B4JEykEMXSkKOpGtF9GKpnQ9l3ZdsU3jBuNS
3MIyuRBWIL3X8KHeM0vlgGIYItmsRc6t5EpeFD0toOEhswATkvoSXtxxExe48VszXyr3heT4d52J
5rJ1FgSzj9Jv3ywgRw7QciUN0ejKUC80WF7ums+SSjxw6ynQnl23V+nb6MYjQabddh9DzGTXwSu1
zKAyxcxhPekyR3exINc98IFiw7jd8uDLOkN+x/nRh9wYJRpBHG7FC+r2J6DyANBWuKET8fGgZKG9
t0AleHvrfX4cUg+IBcDJlqozReSIvA5OiduQrWD0EMoivWgKeFmlCj10BgdJVlWs9fJUtFXIQpSj
SvkPvTmeJlYeXWknGQDW+l9SOI2ZZIXeeqCRc/1Brz0HSTjoj+lqWtN+Esc+CMmFIarxdHX2dVB8
jtsoERU+49wpGCwHbp+02AAlaG0zry0FxE+RduTmq7Z6kO6O5Z3wyZaCN0EmlFcwmN8F9I1TGZAI
8OKO2Z4mKw72u/nVKRwIyc7LM+APhMjm2a0iPN0I3ZQCL5rGKUE9IkbXNkd+K+MvgB0kt/L3yJKC
GESLGQ+dmOD4i1gUf5llHlwoESTmk/VM3KgozCCfM5kNKmGkEvEQu33j+X2R/nAJoyZ7B05zC2Dy
QoR2GANGtSDGjfq4IgTc1lfQQtj3aiUKt73EYiXwILcMbwTOPTz745GzD+mwxnhE4zLVIp/3IH8W
se7cvvrPcQ77AJVEI/JED0ytAikeIcsugJBZfQAFlmQV8NiUlgIi0QJEHvd4aMbzn4H22UGaWkx9
XxGZb1HaUyRuooinfxWIt227hRhhwy4pH6dRXQZCSPao6EyT3XafFdM9XT6/Ymf5FpxybltVBBRt
+hHqsNQyxXtwaH5rdcx1Xv0VFFC8PLFWwSIDt38QMU3Supfy5oQ6HC2Ir7LGyxkf7hVmySZ4R2IK
8DxIgCr580mUsXeqWQ8NIcVgM7CMBrPu+842kUd/jzmYBt8EyaI5Y+8ZU3nGgRXO14nDfvkYeR2f
muHYpvGfux38ySwhKLZnv2mPseHhkvuWr70KTNDd9clMT+B8ga62Tcv2SQKc7llhvBPHJUY7jPe5
OlwfuEiEJpJUal4W2d7NEaG4rfK7gqX84GxXT8vNfAMHfErEH2aCw7WMx1iC8IXUSJv/rYGb6S7s
sUmdApP89VzFLTokFb438ht2Ix1B54MYmZ150XILK4Zjraj4XmVjNNPMG3TKHO89ILU9JECf+8Y9
qpqduxCOLaanwITJ9rHrYbyWCyHyoiGNw9yGVju8DZdw7CUduB1LAR/pNqbff1in63BaXAy3Smhn
T+EHNXSijwGkcVGnenztpL4aV5eepv7C/kAx2VuuU+uUCY0yebVxiLKo5SxDnJTtjIRAp5B2EXQX
kBE3IxbiCzPAng9YWX/rdJ+CoaKz2zEtWVr8XwfnPmwnID1n7MiIhZtAZsXiOBjkawEfMLeXpIdl
74q6ZluD/eAUFARxouw6cMJhXF6A7qApu7u79Mu1EbHCMNoEi9kWjEoRJ5tVyGCqy6c0h4s5gKh4
7ipukmGIR8fYqEQDKEbGYwULvCh7eLiOz1v1d0JMkXTG3bPOAuiYypw4y2Seqa7WscVDL3Fl757q
Dc39+QxNCiVHqyCudVry1dGaZsYH4Ik4uRDpIsg1+06YrwGVp0YWNrnUDMKRHOJNm+Bdn5y+8Th1
sp/hu7c8RGgDeS2oQLoTSlH9EwiyHnPAxg1nOibCknDBxuA3/tuL7yNmeMdtOY6Oxyqt4w5taW2y
Uo4vRmBnQnrT7l21ItEyDbVoUJ8vyinn+tnjxtx15o7ZGt4KmpVVWscAakvo2PnnWuJjR/dMyxB7
VOr/DIQk+XryaTH6QwGq5wZ4TXbKo9IzntGc5s8Kgq0NZ2Dw9nEuzDL20B5+ClYjGAlpRJ8j5MuL
39Fu4A6abRKE/2aWoTiOKkml7Fn1KthxL/JvWclPTRb3f0cl9r0EEGA8nB/s7+wrt5vGm2iUx4qn
gMXezUvaK99D7aJcRSHOzUwAsG/Aaui0uW4ZsEks7kkx5hfCk/Ctlpud4ER7NKEkWdcwr2DBZpuC
UYIJSEHkD8LAb2IFCjP0AEYlgb5+UryRny0tsqGWe/NtG1vnZdOImsRL/khTm0UHavEfrG4BWr7x
bDiLWwTExcxQpkA1MAVvzk/0l2/RRuqquS7NsDrbXLu3L4KB0wCS2A/F27AwHTKTchQgOHjXbZPl
/GhJl6dHs2T4p073I0PhqR9YlMlo2sczwmY0oRUFp0LBoTVnpu0TopPA3cHOSqfXj/u+XwrnfRz0
u/P1JVP21RP42aORBK96a+hq5UvF2ifaqMKeTLv+hdG5+GexQZQutIH4LzQJvjFL6g2EbyXhn+pH
s/9jJcILBNOhtS228zYDfcna8x/i5XX7DSLQzftApTluVxrUIAaDLaV+osAPxaJgHT93HQZHrSB7
v0ZCVxGxxnAVYaqVyWhCDl2s4EcfBlTrAAW2c8S7ozMOf6CMucAofTzehYNwgjpgqwxtv3a+yj74
lx7VHHw9OhkCtengHMiRiHU3eK4NNS34eE6mJDbvIPtq3mTd19KQT3heeFpiIXFN5YBwRVmrqTs/
48ig6h7lPF6U9kLjuNNxCD1t6rKS8UJ14z/LnZsxyh0C34QzChY1wCw+UgpU6vg79g2wyeNMf2Sy
TytcH1QQXvQijgGBLETJikUOCqD4xxWpsLwzEzQZTqXxHfPJriHPupH3bfZK0zhE4usSLPICs9ma
EC7idMVlY8V9kN1vBuqfm6vw30XNwcIHRiE6Axcl8wtaQjJE0qCxI7/i3If43ldd1KSk1HL8H7dw
6TpqSwKDbUjsp2dtPNeYN/Pc0jei9CDBd2g3Fvs1cqdsbhORI09JyC/A3unuG7bewwxKK4PQzx//
JSrntiKl+pUrh8wp2dJZNRx++3zns68GjiTUFWIUZ/3T2q4SLVnZ/WXlsr5pJLd8W3Cab2UOcgCm
+uavEQQrMXv/AQU0klM02dkLTnY2RwJZu2OtxLmhXK1fz9d6HJ9npi7ClAAE0pWO9D5RLLGP+Wsj
m1SQSAU9PHaI5EE7pnC2Qn3bvyFx9pLtZ9hqvmiRr4OPG1G/OtTPkH3VwwIbPLAoA6lL6GL1fSp9
akWKXRgGg+5Q2o5YPhm4bPa41lZcFZXWPk1qYIzHdlk4xCFAmNt65Zl471SIbhh0ZjnyxGUA/od7
QFa+Vj04HaUBScMLLXpMxTozRjEKuVTE44PfZF4lP73LSQ/U/sISMGckC5MuPutDFyCZjYTElt5n
ZytAYIaGEhV+9qxX7lQUV2YZ2ka2mWGknW87Opc9zegyZJ4hS1M3gB6icYSwqZHOCLKVuTivmolq
rL82KvqQdsaNrJ+ZQrpzvFgJRWJ+FtC5KmZZNML2AWIbw6EvHJYfcpEEwDJyFeOGgPWtfaVzzyev
4ua+juNuAFQjYTPxoesnxO1VqWylyNsEOWw+DHLQsrlZ2TkFF0sWdXbjUU06ET8VwyS6ZXUdano1
pJwceDT5MaTlbr83SW6SSTgZs4GKGUi1ZJZFmDDcMtIUOnN8yuGXOXa7zo6MhRWfKhzLpNSp7bF7
rLTTESHmktshRATrbqo7vzJ+9t8SpfYzLalZrT3HhxVHwzR2OcftJgZ8qKizzfm1kzWXt5wslljq
/78EiieOzXXYTpoxhLvzRjSksKteaJDQMginfgcJxdMDSFM2yBhwnG71S0IwTRBRyJia5AILu/iF
948ZyobnWCNdW+vx4CohwS8eqQDesq9BKkWEES+xeIfvtecmMwO16NP+vO6oTtXUyIjHQrLNeOp6
aHKYHjD98GhgADICdtNVWSF281xKmptw6UBmWcSursx24LTFzC3aMYs6O9jqckfWUbOEVusF+Vta
YNClzOGoDtW4VRwTEN1KayrkAzZV8117/bF7aUUAC8/UJFtdJXfHgZEr3ZvHkTn0GD2P1y+RnyZi
BbIfJoXnALA6XpPeCEzILis1nFvVVP6QM9FEr1nR3JQ/tEg9N5knGBYdWcXVZK0TywUFxuePrSAz
6PmbomPMxv88XKYfL3r7VMpDo+rFLF3gtht0pwP7WC5+zptRNveiAjakKAK2qESfvAbvOF7WWKS1
cLsYR4+Dnpv9iPT81CY2ygnKsCFtwlGg93iXKO0oDFSYBNzgRMvPyNNKh4HrX96H7RBN0P9QT5Kk
71gL+DWIjTusex3BDgj/7Sxh2cAzTJZCSE7TEoKrbsDNch2gPGFc5oiVTQa1dPvCGBqWDed6EOCa
14u3WiGmBXs2Fuy9S88ixEKtZ8PhajRNNHYLQa7XzPGLRnVH4OHKGZN6G5J2pHCVKTSeQ46Kgy9E
IMD3FBztHzveKbEG0I8+LSvkyxX1560mtvA0HrM3KDS0rIeLLCw597IfrS2Z0D9xfGe+Bg9FPUxb
GhmsVNkIjq6CQseyT4rYSv+L8ijfMUtjD0XjdZf/XlPEK71act2lVF+WsRSs3p+MskvBWpr0gHop
D5pFJm0R/oFYA+0++DUuzRLwcrpNYUvURkI0kANS5y2edUrIo6P5Y81sHsJpllzXBH6b/ZrdC7YL
9l+e6zZzVRrfGT9jQk4q/sNLQ2tMrQ7XG2JQ7S19qEIm3YuNzTDXEu4M6FTFFVopYgP/rmddCDnZ
5blzVWYTCayK4LdtH7z4FFL7zZixmsCff8SO4auZUkcGCc3TtqsZzuUV518SNiGeL27qH24PaNSm
y3QAqGeZ8rBMJ3D3Kbm6J9kNzhy+ry8JxkAim6URGFTHizh8bdX57NGSnWvHjAp4ZD6b2M37gayU
8nyxpofKxD/iOhL1E/MzzMjWOoT0766tTp8UWHvdNJLbhPM2bFNAi7duqgJ6EGWYwrvJhqPIZJ8A
heFfkz/PvVPNHn1GOPuGpHiVRqZMP3qP86Zvcc5oU9ycdB6o1Rz0NSmlBYxC6YdWRTXmTmJTrGii
Efa3BVCJMByGmj9ojPS5kp6rxO2pT4tP991qT7eoxr9XC46wVdLAGonxA8XC5FoA9227NrgXHaKR
Q/NlBYPLRgCGjTXtUQhh+s5IaJzyPpynLN9wu3PIBBapOS/CW0VjBRz2o0+zzplbnVyb8dGiThTa
OPKlgcgrja/aD+e7dgiIv7JBY3GmAhjyUcDoj1/jaLNYlLpSzJRTOH27zlfyI+WaAC4HHEoM8MPd
xMA4PYYVTpToF5XGj9UuYqf0AP8M0ZKKfuYYm1700JPh73NMEsDA711CuboOk3Fdob5YghmjJYmZ
ZJkfitMOPbtM2rbTqeOm1d/XlL1EaKDxGccjwCReYI7r6K7I/QwvmiE+m+oSH6pn1C7hlBbXOElw
aMzy7vLUTEGbdHSZyLNtNkGJd1botfw2uGxat8ACEgaRRQY3dvTXY85Z7/YcotBh4zGCdLph30aa
eIPnZtCse+bMTD7t0/YJBhR8nobtEJ/OHjOxqLBMVc3lS5Ji5BWYXvVDePLp6ixJjE+o/pGaUA/A
wdeZ3jf9OxRwEBEXdn0+s+5WOrOQRzWzt8mYaPADB9TVYFO8ZRe5v3Cz16FQ+phkH1mmKweVeorf
1RgRpOJMCcGNa0JKv25h+JprsR8m8eyh8plwWqLQDzjHE7vZIw9WQpIka1OcWhaxr/ThO8rucWk6
VSRvyCrRbHJfEMEoNgC884/gfNjgU9bBlzp+GVV6uNqFgU96k17DXbK58qF/PujEPLIkOf48/t7m
fXyq5GPlz7weHdIyj6mYno5tTDMhCpo+UDKJ/BI886esmJlB9+BwgZlxIrYtVb/iqVj4P95nWMX9
vklCNhf3mmNkFWZB8fDi/PVfi3wTJfwiSyTeaLReEfMY26QeC1Aovpop8oUpTkVYMGQA7Lf3ptbr
BaxjAg0Uk3lLEXwnVSAx9DE02/FsENVI3up6WgzkkKOFNO2T/z96fFEDJ1Mlmjj3+XC2C+RlpXDz
XgUZRi3ucFzGxIQOjpfxGURZ7J0mymeKCCDGcVLva/DIO6hxJEFP0qcjYvd9uCeXkFj2FsJDEI9k
i3XWfP/OEBPVaOZFxSjM/MAQIYYrcrhwAultMpMu2anGCIgShqQf4C10T2qdb9W+8k0ArFIJ321L
K9ipA4Cl4RRudp+HbMxtxc7Y/QdTrguVRhNTazaGanV2S126DIwPEHjKy0cQE4vBw6cTiQty+y3V
XOQty0LKZt+MXWGWo0fLtFZZQQUtmx+vCZNM170jmPGRUnCXEF309ey0Mt5RxWdpeGC15e98xhl8
gLp1EymmBM7z6c/p498Akq8HMX8PGxSO32ZpQHtOxFcL2xuxZaYhJUMl2IVrvhZfUkS6kWD/elBS
bgG3mlVbXnTmoPGoMNs7SandnukVUHOSWiE+ScnxR/iEyaqavWT3x292ElHLq+S8RxGczI+ESDBm
j2RjXGIfJV+Skcf4q+W8RJqoF5+1zKeNglZKN3JCGyV/eiye0mjXSpapmKWljqX2+KaHI5uFRGSB
KdpHZtaEg380Hgeam7byIyzNSkFQFg/U+rkZLQICmLZyJhO6ZiU7mcTSEDEuVqCa/Wfs0vegCZtt
g5Z5WsOeXsNGOJP+19UbK+G3Yxlz+pijBG83cQzrTBvo/nUjeNpfsqNsUaPU1+l9Ij8BY8hbrECl
m6sL8maRzbuCY+b1AaHlmT0fiWfzqydvLtpjn2eymSdxjf9tz5iPQnF6BkPhn/N3mS/o044JG2zD
7IYw90x0A+yuhPDVIdb8bkdvh1t/I0meIVpICs2tU2gJ97kPHSR0UfuHduBszRCGe6k/DJpn5Whi
HbCywXRpFzDxLoELGxG68iZI0CXJGGDpDoPD2uD8aBrqqttVhLYCbwh6kIVvGiB+HQLkSlhy4aEE
lgMYD+JaB+jXn7LE31JMoJzFuhaiI1bHuc3VQnrJwoPNVkeMfH032pgWEyi/m4h2X6U1Eh8MS5nW
GY0b+OZ4tKjEWvlJO7PH6iWt/3jbOcWDRZu5gGdpQZ52Q9uKnBTWtrmCVLUgdvefcZVLi5PInqkM
+Du4pfS6FeaztHcCZTzBI7e8pQpJF7i2Xu9p83tXn6N16o8p0iUEnyYEdpWNpH8+sPFCwqmcQ11f
4J9b5U8/4lgyECaWyRgFgc0ONlMjdRB+/hjmIcFGSGQR+1JgCKBVRSJ+GXzktInxyIerkZKHFzyy
Xjvf67JBA1+94GopjTQgCvVJXLZC2JYbPFVlHqWO1fZJmsmMmCOPXrEwp3kPN8LxrZhFUgJ+kBtO
7Q1IWi8wvLLInFPOR83TPoaY20neYEiBJKsXtDoNv2/nP8WWTdkeymgowynvzzcedmKkfbuGCDxW
/npte6MFMpeA9iBdXLuWjvFSaVbcoPT+sduvIRTZdTfNHSj77sv0jKSz0HLn2wBlfB1Tj0a9FXcs
yDok6nKx004fwferQ6ruoDcR7MTRn2v+X+ns9Ov6X6N08CWcIKc0hSBaRe/HUya8STzqlbDQv8e3
+fD/JB5oY461mK3n3TSyCGf+0l0K6BslOPeoFX8z01ZnWXQ4d+gnNe3Z0oHbgZ+1wkL1kWQg6wzz
0iR6zANhH5L+9EZ0pZN4DLOQ0mtwDkh4wcKNfpJSzPWYVOqQ85kIEGf2mYx4t0sP02jqgtuGEkYg
C4xfeTqgsfvjbv27w1FPJg8nKpZiPknjBYaGUVOTrO/mGIlJZBH8bF1unG+vnB+SQ15n45/Rwjmi
kiNvYIZac5tQuROaJOMbIfyWeBeMiIYFKbHcU6BFuYd5dflyrqt3xy1qWVY7meOGWBy1zrwQ7Ahs
mt5csPmLO367ss+Eaj1jTgJsIsv22/Gg3EH+RIqk8XZfWLsR+vyP79LIqt/iB+qCOLxPfqIXXXy0
tInCYTMWPhrsgLuDiXyCjoQjM0oDutf/Wu0XpI5cw2UD/BBZvv1JTiyQPn9BRIU9tw/3RxLIuKEH
QKUO1OHV9SsLoJHw/eWa74GKOW7dcUtbrNzKVe0i20furzoL6Rv2AOPRU2/GfwBhaSH/x6lufKWe
cuA+mmrsM+wT6xmGoj8zvCfnZ5QQNmVo3u8NHqdIZnIGQJ8Z82VrF8GOWIk6em9xzRJhy0fT0FQ1
+kYdxeRcb9aWOBHc9OTFnLPlGUGVP879rrMqiVC+Qs3JIvtOuSweWWTJlLE0tLNxD1fMkNVwSUrC
7w/GXnQxvK9franESQIB1y2QlEeIb2B40EO/5lNB704k8MGsN4sy2I1C0GPiWnE29RdtAQfEWJxM
/+wbvj/gIPh7mNbzIs/OBhxZyX4FkoIeNXuidGa82iKNY2rjkpCObpSzEJ3iB68yXKwiYM9FFPTG
GcofSpg0ShHm+qECnLhJgmQq2EOu5lKaQffVtOy5u7+YRa34UM9tKfC3yjI1Jq++BqM49lothUET
RpPFtH7HspmrWrHIb5soN/UHUu1Qm9iZL3cqVBODXcqZe+SqNaQENfs4OZPsGI9QING6fpfQ+fxq
xhK/zKYVp5s4weOvyVR87wR5h+8MEUWFNGql6vzqxwV6oEAKVwUn3ukqw7oB+CIAhLYrettSU3Ei
VPspf+OQFtAqdTNQZUzHnEf//8qXSuLZjL+RE74yZxumHC4vHeLj+OAhWnm0T7zmG4oaPfUVUeA6
3MElnLa1TnYhVL7hgs6+9vHFdW3ylS2hiHD48HZRqD1W6hXC1JnLiKwRhvgm+CpnIffVl+EIYUyx
US8e0L7Cfp9J3oX4Wsr7mLfzmvz5sY1oxDB1Kz5396KUt4Lc9MgEUSayUODQJXtusIvf5lWk5uyn
xl0OodcfG6Y/IqKRkXu3wPhIRhSzzuG8FTPKu45Er2/+bYqzIphrN+amLNp9S+RFl7S2wfddfs8w
Vh0RBEgSzt9QGtmXUQl2Jf4+B0J1YGBk883HFLDoFPVO/WRRN9DayOa2r9RHbVNT5UwQvGnsX1NP
1+aANWEqm7Qj/poRA9K39x4nfxeEfjMOKgwZC5lfx1uCeMfQOsGft/JnvCSegxRYCdUGGvLNOy43
6yFYUPdfOO5lIb0G8TYDN1teH/ANEzbn0yUG3GzN69ypDrq/FgzSZrk1ETu/KDbGFOnKst5X8L6K
+d1/GJhJPX4oUcD3iL0KynCPSyvqR9i7UmZG8K1KZcZOEgPQiQWODOGKam5roxn/qwHEyxe5kaeH
IxwFSCvex5eTGfWqGGR5dy5Ba00zfY/jxcpztuDN2mCu9j5O5/+vmk6xvhDyFMyjWgT+8MCbJJuE
ShDzvJJy38abgNAN1Yc3JvwfGXNiA/L8j1WwQ0rkDlZC0xMspSZGlkD4tdDxjIg2UHomzP50xcJo
ukbJ/+CLQt1Ar9InxIlpUDv4ozy049dy12s6Gt8CRMDy0laaPaM6eU8EVIMJv2rz94rJ/u+osbzE
3Y03fwKWFcxD8sAEP+BxqWI3OV4VRXhNAKw6dGtBc6t2NgbnVQFFeRWywDZn5R+++TAMvbkRkebs
PBZ7lktEWUWF5ppSZz0gt7dVbXhTC/ElLNXXIoGFiJeoUbsrFwl16dNFFpStUSRa5iMDwvc5hPws
7l3H41ikuycc0vCi7TBqCoUTP1hoeP6eR706vqlJJVzI+B1Q1KGotKHCtqGiBSzHalAXm8f/AU90
EoGXGy9ith+AimC94bWs6lZlJfQMn+s4Uhhm7F7+oanXbvtn4FS7rGkBYDOWWbjB69GXaYP16pk1
rbUgnBn+IDhkTstA4C+Fxb4avw6k9DKwyI8wAJZTUtk+a2h1pU6NONMbJ56wp+YgsNhj3YaGf72P
NC3nreeyC1scToxUU6fP5ORZCOOFwreb9DgQI6PtHZdEW68TOwkkObop48zE1JUPmbBpr3j4B8DK
oRIbzQqwqXpIkpF4r1J7jPDh3c5UVcyR9S/hBHgGAPCcwGMQ61ea9WAfKWGsy3OkAykC9PBxJdlF
COHjs6QldNpMPUvxGJmvpYKSVutcluzOnhyxr5o9gNAyrM0bYbiyBN5Ye9DMVtKTez0byXK01q9S
UvAv+aU7Az0ARonP1GjMXJ0MMGfb+Due3a+juDlZ2WeTxYWVKWDbmjX4lFXOE0mIycJKUsAwZLP3
vx4cqmKrE9BhuVZ4AY8j6ypzJNsITAJfHAqu/o620J8HzNH7aYGFx3he+AytwMgTt+ZLUfjnvPAy
wDVWRIk2GARSk8Kc1TvaFxpKSPHr/EmWlJfJQ4E6Y+QQnaPNf/dQ07FD/0grD07dpp2b7vDSvzTO
zU9o7FjTGTtv/UgHNH/C4vlEmMveJSzdDiNKi943zb0xc2/PGLTC3iouNIHN7qTSsLCLOfz1L5A1
ZPTaKPQxiVUsJkS+cFenMVIgAzy8q0ENioUozGJYCqsYkmL2jrpFGA8eeRbhRCi6bn0nYyd0e3jC
4EBtD1bs6ca3XayKL5DRVgrgWY4GSMBdnZVhr20gbRTMYXcoZpsdzGTj2QknLO76nsLx+JhEW/VZ
EIfZgZjtcnmSMUUio4/XBGBYwNJ2fG0FbF/lukyqh/zsqL2DBWhd3LCwa12Jq2X8GU48jWxAfHZU
2d7okhg+IfrxarlLml+gAuYpIEI9R3qxud3yvFCcT2I6JrMF9v9xuzYgyKs19aG02hF6oi4LEKGv
eVGgZW11n2fz6uajKSAa/qqW75oH+oqv889wGZwEO8YIGSIKFtHFTG6oktYmfdMceG1fH1ZjQR5I
FD9bS4Z3lO2N4+v868p5ATqhsxrqnUy7AagBNb0jJKX7Qgh1SUVbsnVvetPBWpAs+n/T0UjNbux7
KWYe2EwM9P1X0v8v/+t78wkkCFk37+BZy2x/D8jx2jE+E70t469yF2cgynfiqQYNArd6AfyrEPDq
Cia2NcxZKksOh+ZoUdEA6lpZKO7PXQMJ8tbEeZwL/4WR6JVKk6C+jCntyQbePuW3ofJe5O9hXEEf
NGTB8ki5nMkABYpnUpxvmCl6ARGzM2ZFuRhVkkp5mTLcpAtaYGWfjoabvFki1oJEUh5PUa7pYNq8
ZpPhA9k9jCXlOFVJ/0qa0lc1JEEqbHOIRCIh7HPo/JLZYGbO9P9SxG6o3ETs663WTDqCwTCxTDEH
BGJjLSLPTbDq1cHtJlq7ERPfPCPC3H0u0MjR8x4uKa4h0eIoFox9DiYrGJ47zc9QH6X7qdPqkOUD
3TdUfAX29db/tkRiQXsEvst+fdCOWfsX1HojUC/2CCHwz3YAKyX/AnXk4AnWksdnYABHEtmrC1F3
1oC6YIDq0o0Ku6PKwuu8vQDCHIQtEIb4xLmqqEPJvD+AXYQfjbGa5mdhW7iTnLlHKTv7unNWoxIR
yF4aUArQ9ny4BGGWyTeaimxjAGUoHokuMib3ZYg/i5yDxEuNhPF4e7Z+7XBedmdC0unlgd8I2wYF
JFB09Owkls6WdZ/pYcLLGNjWPUcq9XSlFjO3A/FAX1ALoIzMwBR/qzpXC+4vCaRm1BMoquQLygfN
ey/vJppQdjVNd5a7pB/UKrHkw/t2JNAAby6EbibvdlK5xxJUsS9EIg8WsNbDvhJR2MGgrDk5ls9Q
y+V0YwEs8sAGFaNhRewu7G8xatfyxCcvgwxCNZT0Rb2qQ7S7IvieZpWgUcLAJI3rwVx1NCQdSdbK
3AyoNzRcurT+NtxDWWt16Xs1sBYU1o+qZ0jXj9CY449qPazg5sqfXg6a1q8fP+IoqWurp0hc7P4t
aMa8VgoBb1D3P91SFkK3Idno1u/5ywIQds4AimwpUxaNxlyfrYR1/elf5R6T0YdodPLtoXPoQ2rz
5Bgg69IIIn2itN90zzYZvDAybVkaJxp056ahwgWnf9w2YEj9mnVfBIUpYi9Ge+bVnVnBzi3Z6ZPN
xdKJcxvq8z59ToCwcT0fd/SlcEg+TjCX5jAtkuZaViXSTvUnO5yzexpJepGoecRV4qQype5/Q6QI
C8ObBk+2kyA7VghdyCMHNckxovGYe2HaNHY72ZyiE/ZtBUAN04mhNWU1RzKap5yvTYGVTkjM1DmN
QCJw+01ddvQoa/xk1rUvitQfcUIxkSgWnE/sUYsfHzY/4dY/LKKxUpKaU1Rkdw5T70avMRl/zcKz
eGt5qOuYTwi1PojmHZjya6I5KWGxoHKHlFdnFjm/IrRQW3iq73TnT7I/nGjR+CL+ObCD8svFrWJ9
nC7um9DEJijL/5yh5emhh2nZMzhMy7XcvM2pv687UULHKOihNRSU37CRYb7z0QyZGhc7hEeevEwB
/t5h6h7ScO6NcYRl8e8lUGy8oP9MJkdMyZ46j+3+xhCrQKKa7KXXp32QGxBBttV94dTxyvxTE079
IiJ4Z16mSEme0y6nohDQK5sYGIgJIJJlAWpjoFSodBwDZRGlyeMDkh6r7OXPoc3BkizSULQYjkkd
ySR8AWi+o5JlBBGDZEvuT7VvUnI1/fb5CzAb9wRmo3iaS6X0DVg9EYa2YD7528ijMOC/jZSxVe1m
Sf0/NMLSjO4arFZbf87vezxgnsoH6dnSg1jJFYujYQ5YmlSdb1JmYYmF94d7Acou4x5VzojdB0Ks
4+MSYZw/FDUhrcd3yCLtEK+1MqnIdy6BjgY9mfW1I0qKW/KHOY6Yh5ocG/Y+QTnAcDPBQJ8M3DQr
sPn3SEOT02P1fOnZEzhF3JgbANaIC90vvbHuSZfhuKjBbDxMopLAoUcuwxNtxbd7qNCLgtNLhTOD
SnpysgINFoJeZVk6rykrVdJZAoCVHERTw/QLGoK5YO4b6IcWGLhn1V4HiK2xWX7dweCmkopx7GHj
uAuzs/5xTBDd1gEH8J6SVBi8wyAUoCPJql4c4Gi3rGqJTeKPcEaq+tl9d8g2ReZZieNeJWK8dJyW
ogqQnSEBOoGsd7XBs7Ghqrq3MN3DYrkPV0gFWJybiLOauWohfEp7KFShCGrX4VQP8xVh2y/CJ9PQ
THnazNYDW/Gh5kK6djZyvTzIejfKF/rf2XT/G+CE72UhMMRPXLbvAufTKzpgaDTsZJKA1wk5W767
e3n1pr9EXxC6aYLjdSOtvJEPKeN6auOFgXws7/d8y0oS/sXGW4KDh9hJq6IjeBOFgvWRRJujw8Rd
u4zm5lD+RAOW2dQXGqhRnFj+T5gHz+bCEEW+swPupSh/KmZE4sXBauuo9KKuBhi8kYPMcsEpLRPU
I8BgcY8cJoZqz/QAcj1/VcVYYOQyDGHb30U4mo4K5SLK0xvAOrpkTcibeiCpaToxN2oOG+VxXm22
ckwnWIAMIkOfEJMcvwG686jpfLDDhevt8AHQRNVMKIjtASG2drq4TimJWm+2DRST0bLYREPey9CF
4IPjLCL0rl99uBQXcR91n2q6DvI5JfPP7HhuDA0N+aslGQVM8rUbdcUAHhLY2p8r+nSqypj3z73x
xK/Ir463yCWSoO0qwBbZQQwO99hZwhyALgH9VaSWoeypVtT2akfSuYcEZOM95wj3FMNdF+pkpYmN
rI8vZ3I8RNZO9E5koZNqjqUp+yDIviTgkgG0ytxPXx5a8zfXgXVXNjh1mSDUTWF2+ZgXB7qdynrc
QFZx1Jg1g0/XJeEs023+I3G4AMnM62Fj+Z4ctH0ymrtRkqg0TS+fifyVEH5zqTOwAHsOFFPnP8lr
AJ23ySOGjiad6Yt1s4ZohUskpkGerUUaOwsWcqHfw2+7veSxals3rJCK2J+PG9zHvhAs678iDcaU
+G0D4cpdJtSwhBhkzMzMfti4IAs4aJOr+eUzN6Q1LSIqZrQSG2QKdocjqjy0puxBlcJV7QzZnKEW
qUxXjTKnofm8Oohpb66RINqNe7+irV/GUR11y74NYl3TtNoo7S/zAQ2nF3UUQ0gQ4dmmOG9qv/Mt
okX2QWE2nrHEsBdrjsggqX7E7hogvwAUZaP1/vLVkp0nYjA74NDixSEgapP0B0cpTUZwOFpFexDc
lWKyrQPSDJIP6x1o+IrT9XlPuM9UQioCywAr/lv5AYcK9g4X+KKOB1Zk+e2FDElPNW8Z8Iy7Odp1
4rwj9D7uMKxqwva7b0HdwjfKDIrCJi3T9Fi44LEnFxXBvWQYqgjoAQiOIhnaIrs/IHBRFAdQcCfN
pkUmcz2zgBgYb614uofd3+3JuTRg66IqAF7SS90z+VrEyZgMt8W3bwfLfdacYepq5Q1lHq4lKo8f
tbKjjnCCeHAKCAelnC9ozcHX1dokszvME/jIJay2CxhwEtNonJUDK4z80iIsGUGUqmL+0XRI+Q3/
jzbgF5QjqNXzXE2Zlkj6a8RcyuyYteHL2L5k4txrWOM9QixVy22w+pWW5hjUPSw9TMWR6LGcdd3n
1UXG0k9LReC1T3arNWahsvZFok4TOV7v3k9VdYRs8621xpAKSQeHmK1xVv/zvRDtSdKcrM9x4OOK
ydGW2iod2KWb+jMNyXGK7CD7IEU4aK3uv+GCSj3zOWjAVJ1Hj/zBX0MNZYxuTMDOi7aPQHTIU9XT
zTyt06ZQ1lNIcBMfKhYb3x/15FGFvKIfC5Ic8dg7C+MP4hFTk566ZhfuIoMVgVJj9CyVhXjpkMK+
mSCI4e7SNxQnQ8MjReG4gVEg67Y82M79EgP00Qme7XBS7qBgU3/IYBmVIMv/xSMpzNkG63JRu01m
K8MAJN8HYSN3w2GJu956TpcdIrqUKhLc0pJ1C41cBbgbDh7mvgcSxHUH7DUNn59+EhvNDlOrU45Q
/zzdcAUR/A6BKAwyWMlZoCmOacqQ9ekhYi+eylkdK5HUzSHMSY9qwhinyg6MzURbUmMTyWqAURX+
psj5nn6HncWAVYO2XT0+U11dSjvxJBV6q9sv2TuItBRoM+xwLwWvPXqZ++ONvaApldgxS0KGocDs
3jEuXD/gqOelEz3/gWYQkM9aRZQsduzSKMQU8eIBcxuGvfpmPb27RrYNPtgZyWco0J0fPt44aKmd
5iQDbitu5tKnGuPkEtbk0BSVEPhfnsKHIyp/FromAUIh2KK+GvRh2OlilVsCtZ3XqRXV60da0GyJ
dDgNKDwpndrYH27ukmdjJGf+jOUg1NfPwkb42rIEtpF6pTFsJiMvyMfTbP9/9VC2CzeKlnb7kSmq
6ASoTqX7XAHNAPcgHjhc+Fus6k+T9jc0COAFbiKfxXlatAi8Arnj4Tzdfjr0tJ9lE/0gttn5l+f2
GpNvHwxYmQADVzRxDRpPTs+WHDZavghHycjlxBdMl9AuhIzyGgBcBYe5Hn72mTSWbspbANK4+U77
dTmI/MPUA990tJ/Avb8/9Jp8WSFIoNFvB2lrNqj5/u3K4Euc8RXyLT44HliU02M5+1Rr71Cxr5E2
E5QzRzIMV515hUKqnC8RZM+5yMqMURsjYxGwm3uUGH8Xyqr0mY4jxSw17Pz7PYZuUc/9gpna9NVG
DWAq4VyiO9D71qVmtevjNXYSkuMGeSfX0RW0y+rxwhg72UVM1ueIGPVn0ldgGViog6O5oO3aLA7L
tVKd+DjAKQ9qXIVrqf5lUR9AjV2tw1pH3aZwh6vLWNfEsi1+4pMclKzyuDzn4lOZhmt4LQg2c3hd
i3eBP5aXMIFSvFT8f9dH89fody8h/+tklrg34cGCTX0/OnEULdkUM7VEJZ8KRyp6rrpCZ+p/33hu
c95LKFNBV5RDqSsgsvHyK2+dSvtbfmkvsShH9+YdEOuCS7RNEe7n6k03UH9h1b7I9YDdWBIZweJI
+U450pWQ3r7S6ku/Khs1AqRu9+qw/knNVUDpIo+E9yamzKcYE4QxSnegK3D7dNZ8sbE11jaoinTD
ZMBenNIc4qkRgj34CLtpSnLPBrZKA1cHBvGhDDo2JL3NTaOCcsX9FSbWJTw7MOgRtI/kVMVdBaXD
0G98O6qLCXCtJEDEt+syeVPVHidoiKachUq4UZ4mXuLFem0bmXdEARLVwX3jqhjCRBnHHbmRmsma
1M056NycZrO+0qQeULhdogSyOh0BY91LYoV3jjwnqsJyPfKYUSFoDYnOYUPV/enfVynJmzu4cZ7l
mB5zWjYNAQWyd3ZCZnxHtc6xYM2iv/76gT7txZL8bfqOP8MXN8RbsQD6DjlVY/7qn7UgSZQMSrtb
oU76EXWfPWKeIu2YkC/Ea7qLXBifLcYtVqev9jEP8b+eT5KPE5tYbgBR25xSB9qSaO0Oi7DIcsv5
btMbOks8Ok1tQz6KEqGVyCrCps6QmhCQbxNvLSgXquUtjNio4EMmdJh71VF/6kzlR3+GKoWrAwtx
b33wpfsdZoMbOQyTv5g9FlHSDua4+OiGNSz2UNW4XJttzZJVtX9v2orMb+iGdnzBjnhfGVWafVh/
v/f2uroJRu3i17HHkNyljVxmUyAZb7pHfr5RFYPOqUTXACRuC+KYv9OTU0pcKXD3PwYgp6Ektupl
M9KBR9szaApod1z+6qDNqIwePxd6YNFdIrlcPPUT8dQkRAgraXxxvAp1ES2i3FPeQoYGfigthZQb
OImEY9MkRvgriPklaRwCmteZL6yKv58p/pMRgSnxvolCIEcF3NGRlWhXWdLbiX1RHyYhkdk5h4rJ
9iQbVBvDuegjNXJR30QdWcFTrUn9mXUiCdOWxormLSwZVkwi5fVG1TrPSyw+CCJ/Qkc4NYdauTcn
m0fG16c+hZbfesUrB091l9lSfftgwDdTMBAGRTajObXm+/I6OR+ePlbXLQZqLlDxPLHTsYzImMzh
29H0gc9LoGDANlXVuBREpMgeaLHG/tPvkIFLU5nViFBu+EARIZQZ/dXz3LAWmqBmTokSjQ+Ojr+/
SMM+KrGQrN/oU/ifoscRk0H3QK2BPfxuiLrEtyXoktXeSrUZlMhz+mkn9sCCj3Xu2nlznmHiXzv6
PWRvbhylpQQFluACvcOizvaKKESquY5izKHtAvWy9oCKonANbUb/udbunt06bjzSiKRIsTXq1BiM
BwHlX1cJj4J2rXhdUjDvcK69Aq6FwYEbemoO3cHkv44Rd/JJgVwmAoqP0H5UuojlbAbg3mfEGQSC
3F8t2JuOCmVvnlsy2Nyr3T565Dous6F+Hlf7cFJundEgHp7XF9l4aYxnzQo8n2dVfHANwxMFr/Lg
qkcGm1HDmxJ8Hy503WF43HmQopxmgMZbfhGQrOo1HbDH5WFbSjv3wR7YD/1Zi4IGzCYl/JeUgc2W
Zqch3/RKvEmVcMiqZb8ir0j+0qfrzd7Ggs5I2Tmy5VnZye0E4WoUt6NDuXIRebC6W05gxAAC1dL/
TZuFUudXYnHCPi9pI3qRKtxB56HzVzHB8drF/DFlTUdfMyRbQJ26FJogX01ceswvkgZUSAIzpc5V
Pus7hKjX5A0TPs+h5tNuhoJMwXNMbP71hunrxmm6cSs45dLfYBz2BNlEDqOb0xjxo5N0LN1m5iBm
dKyo29dDOF+w6Xze7iL9+CTyxtZ13SFuc0FQ5rCXGfsF3h0x8q8pjX1hHQLd0LQfV8JtzkYGpeMy
Nndt/9dnzn/dI2aLsEatQfMqyuPeZnpJAzAX/yNTk2zMvqxMlWY0jAFuzcHchJ+jWL+7Xudchulp
8tm8Vlf/FGWtjciu8/+2YzjgcQYO+Xvm0lmoIMT3wS9rnY9XNcmAcgnA3Cb2vPfogMTpPws5faNX
dar/2xpmgYUZV0eaIgMg6zdc4zu4SmsJ2BWC5Vk/G+1F73a+gpkF3pv9KdQT4JECl4r4tfCLWbUF
dspJfFfCfazE2dN0R7G7ZBGoDaX1fbL87EdTfNBLzPunPUWtbvCzqHaLcjYzdFQv32we3BdRgCST
tfmMGvZAaQiCFCJ1qc8CZTYPrNRRXLA3K7sweqtSp+jpKlvqCRYpHXIsLFAQm+9ZSt9RlSgtCpYh
LwamQkr4z3ErSzxWZVmlXYrKdtMrVzuBiWp3C+zZExWjQk4tBVMkFOTC02TkxL+z/kXRSplnaUXh
7jbZ3uz2G27Dm1I827bM7MYRSFVWGaREZ1zBgeJYmfyDF/XBo5+uO+NyMeSTe4yJr9f8mmZ8wZbl
6pkjCdfzjQuwAVYCnd6TlF4qduuKqfWp4k3UY2GmY/zo5q0gT7tip0w+JwY03f+XhZB1GRI/t9l4
3+Xi7MpaSvPihHYqvDWJIufwtRMtNWMUaikwcj5xsxdZADNqrDBNsH1P4/HmAHlQYNyQplrvFyMn
rwGH82IUfeTulgvYl3i6e8y9p0ez7W9gFS0Nu586ls2pL3moyJ1ShvwAnpuw9sG0zhHS8NFmfrty
5gMAgsSlGHW6NlcqYGw5RsmVBw2KQGwR13SeHHrfZRdFYhMPIXVNTw1CbPPKKVk1VoclQMjWQEhR
9p/xKnL1ClzGCS4hbCDCO5y/pJdbXbPNbVoOyBeNuzmkY0FDKu2OunXlEIg/m2xxQaIJWbdYAk+g
awKH1rySjmIvvQi0FMDElnXND9psNhjtUAYvl0LwrSxxyNEn1wSPE+gqnR/h5qgiAS10y0ppDbEw
0OEvwbu2s9ljKz8HllVzQGkMcsslTcwu81WslHoLOw0rI/z9+uDsnQd6Vlpa4yO/JEQ3hw5T4mBt
YCpxi8x4+fZyvruMnwwl+6VMK4ffg6tHMkClEug10GeejuKJQ76cRHyQlt8mXlvCP5sZWacEIncp
qkyANV16tWtAH4XYgyT0i51EzayvgB5JcJHLbHRi3OK1zQ3T/fyZ6jPRZgI2kEbpmnzqjWG+m4WS
oFMelyDSgW/sPH+BJl13mOkb7l6l3U9yh9ONjqHpOhLnvm9j4bFTkI+Aw3p7UHkE/bHTn/Dj+4O/
Drct6A0rQ6w/tPFkQsF//zvYlySQyg6H1joI1nQvCIJ8+1jiMJlmMyENhKyGXs/fzsLBc3bMcG5x
LK50deva9bg9NnGEagHA6jzIZHTbQb1I1lU7eswjOky17N+o2H7niowzX74Gfa+MvwZi2WJNKVcx
4NvGj4DjBA1zO0LNH+vlznQBecqB14A7Wvr+SsJ8TE/0w+CcQFZYpQ++PHuEJ5KDxIbrZIyVwqsU
8tMZDRIISXCQDjpE7XWbnOZ3RT11kwaX8BJ8Vdpak9V26fU1Q8sdz89oS+/XmhZ/WesiNYGhTRcY
uwn+fLUJcMm+sBNv2kTlmNu2fZCGx+9j8d5MPaDfFcn15rikXjY9etqGlsaIBicHwmW9cvlOYbB7
YXJBfX9PppbIDOiFYsJDoll5lSaCspOHGkTedxRKt8S1gdgNQSxF7/iosPCuEI2+lir45hvU5Poa
ZBOf/7TpB0v/xgOF+8OgIGuWSU4kZbAifC1REn5K1WdsSy5WAn7uQEpiTYWBQSPc2qPPBDnmBn/7
uG6G7egJR9oRK65V30zSaY37pe3Api5oBW3LrYDjGATBjoiSaNeOugEMqbRLxKs27TjDKaouCqZv
KA0txEKiDLOYwGtIlyiDK7h3OV1apPv/ktE8tzkHk9ooXzDM0vtuuZcoAj9M6AFiphl6sPlx3C/h
Ba64QaaNEn2egPpTzu+vYtW4aku90s0bu6x2o+0hcyw4A9B6f6rZ1QrGV7kXv/mPuBPAli0ulXCb
lML9DfevOt4gYJQMVo0drM7vIRLPiAMd+yTk5ia5vta5VgQ0iZ8PrkkC/epzBQGAxdjrYqevtHqJ
wIU+uyZjMpnCwuoPIr8XczZM/n43a5GnuXMubXEVvTv5/qHEOVbPkTIlur8YsAJvbZTpZRQWkwfb
b28HSQhwXTBdG28yT6mAReHq+0HIFJFDbkVPNJzCPXqN6EoDMGmpufo+K6cWirwk9hGN3kLZI4Kj
nE+iczZEAis5WBjDBL9xGLyTsqTgOgS2VcvslBAiE6g37WaZm7vqdIwbAOxkMRvnucGdGvMqe/sf
86hpHDolaHKoUJNGh1ziOs9PZ7cXeV6Zn6uOpWN/jGZsU00FNGKmHxIrUxnrjErgf8mm05TxMKBk
eCVc4jD/EOt9pK4KQwZXKFZTd+mawGyHGPr95u3MsRCZ8nzdIin5UjceFLULObUf79RFimcV8f4R
UslCKYsm77qcx5rBcRs8ac3JsGXTOeT/awOJQ3uyEmuIxDFXY0BeQooquGnoazKz0AtjVBVoVMHu
n16NCxSWXSLCE1V+pwTzT95cV5oXACsd3i0eDvp5XP7NACTrcyiNrxwy9RF15fsCUHqUeWfRka9I
w/LDlJA/DfkRlJC9tRuodCU3PEWtGOkNCXowvUT/HrxCRNuqvG1FVAaUSo+a0ZBn94NfZkA9Sfsy
17JXVfVox0zpbvC2O96qF5eKb1JgkzP+MzZ5SGVSrQrzWHEa3MusAiaLVjyHjLgXQ2lc4/STxikp
8wNT9MQSS7T5i7sTeaemarKsGGjmZkYUQh+tlz8WqT3TKKgT2s5pHo7eR3qd3f181pJ7Mx98Qz4Y
U2IKOJ7V8zLQr3NRs8nXI5SaM1syHu7ZLTALnCNTJNRuqdZ4+8oBgildNbZOJbx6sTZw+JqRves7
0sfGLBez2rrVbVpBvD0RLYl+djkcyTIF0A3zy/sqLczGVibqoNMNkss+k1OZR2RPrNqz1zlS79aJ
/1RUZzOonYxWVgsssraVwrh2X6sfmx521fln+QoSTLMf1CZ2wVrUaTXaYktaEnQbb//XZOdCPDgn
iN9bgRmemXmfpHMZQazwIGnLU0mevfRo2K9gvKFzfty2w6p7z//zkPINkDLICrDsFyE8Mkn6w7Y9
WPtKJffGjGL+lk1yjx3apfCrEGuww87CGCm5bC6C2g0LmKkY0SsFHNoAcczJ0jcQiqdfDyz2kV/Y
f9UuRssgErnMmmOMJMkGqIrJ+thMgvipuJCb+NVg+FACD8GlinG7glV1cyUsJUuAzGb1mdXVaFEW
ymMOeIrIMd7Z1OWsSqL/0r+L6S2qTRbWrAE+zikuXBTu+sa4fNxJnWbMbwyQHJepUCHmOPEOGfkn
DwQtJQw0g6bNUITHqcFMXVrBUV5vdcSuLh4GjR/q/81ShXCiIq4Ju9fUjhzJAgjeV7Tr/Rqg8DEj
KwG/9AFEQVjI2zvOwR26VQubOyuTdUvtBVFsEsbxsKpreYZAFrPP9BoYdh4k8mua5uPlYOIci0u0
qDAHqioyhQpSuS56S4UsWh8a4mZL9CXQM0xSXU+DZmzGjHobfbCJ6zDW7IfBcrQKzXmUvc1Ad3Ei
Nwv4Rp9+ZsNXTlXbWVCnFaUAY9O05UoMpMi/LfSDEab6ZX9oYR1n0V/JE8enSOeUlmk38QIZO2hx
gTz7q7QipBRZONMEGO1dmgd4OCoBtGw4j6Jtfy8/mO2nOeEs9ApJZ/+lUjPxEypBh0fdIGq/kM6w
jlSh8vwFD9p6VmjNN/BXu1WgI4pUgfAFZ7DG/xlEmJj/W4Hoz3AN8wlE0dElZ50PIhiecrxDd7lX
MwLs8IoRbWxj2cvpyVlgAM1tt2cTv5hvoAsEHF0memVYeqey6T7fjStWs+mPmEsTkVhUYmaFzkzY
51kO6v2qvsG6lbh/lChK2ZPEn+tPTXTBRdo2+GWZC9arnf0SId2wPT4iV8de+pD8XoU2HAhlsYq3
Mbov/OvclGriPhVpJROCW4hQDDfQba6FOjNci7PyE9Z7KzSUtKYh89TfXxAn0ZS/6KpWeZUgGUBU
v8/Q4MLIJVnPXFoCpySMAkv9Hc+Yj7+ae71FRPBljw+ljqa4QIRbs59mhqQiiLLY9uAb1iLzZYLI
MZrttKzmj/9O/N10nXh0EGfvdMP0GxOCQLuzJClBGmadWA7May3Mwt9xMbqlM1wN8yIcPK0hB6wa
mIs6zfklM9OVshN/da4hlCJ9Oz4wXZV/PiynWbtXeN1syWFAIpz3XI8FqmX6qCZsaijSS8KIMhzA
Rbf/FgFnbGGmgK6SqA184zSxah4zboq8WUPJ3q03QcX9VdmXeLCdo+yEFCfP+2+ON/m+2LgRsyMI
0xuWSuJv602fs2X8ee3BYiZSEZ3HHQ76lZi63NDTPAbytzvmx0RHw5ngDkMOq3XZpoLi8BwDnVUq
ttab6KBnCkx3TT2SMKhkABIZxu4B0ewCWE1r6Th50wJFA4pxOghcxc2DFzfmd207XPVFknnEm9vI
dUFjd35KQtYdEDGVkBXOro8ELIRqWWOlU38RtorzE7TSVb8S2X87MSFaOaNqiN93N4KKSfG2rfxy
mcYPpAxZifTlk2YaTFZoNjb02ZnkBLhiwFOEukGhstHPAFlM4g4rWW13RnWqe8OAQXHznTqYy0MC
qbifB0nw5ou9ou0RBLp46reCzzRpThxc/2SrQiZnyi9g1ZVF/+IbMpcFM9sazWMSgiMeDmnE/p2G
goKlYAM/5kAXoUcr59hDqus2BDZCx0ExXGVPA5/w2JX2QpKCmBg0xIU7kLg2h743D5KQcRSunL10
eJJNISAGExbcAuc3/uZCAvyAnDGZNPvW0mhuLK1vxjAL3y/0xGXGIs9CPpXtI61OqG/wLWKHe1Js
Xm+kRFU/Y3Mm+Ho2p56zG5DD5wEkKOxNE8LstWZxfpSX62XS7OEKQ/EgIqYZ7Hl9yrhpmYZklVUx
PqCSVv/mewRKlcqZPtKtlPff+Yg/EsztRPEV9+d/Dw+fHcqJdeDx5lDWnSM3bZZAmbDnzmYKPzBN
kZ+ssVDW/omYjfKRq6xx1fxvD1seaSEGLUuF6AS4VVGFS6tWFpBR4GqErgg6ngxzglyACMlmLH7E
maSQ5tJ0Q3XaEMQhIy3vl+Y/ryCf3GDrFQEMDd3GbeT2nGE/SwGrNQq00R3n2kDpfZTWO7bNO2HA
w4B1FnM6oCJqXpAqv6yITcUDthhkqDU70DwiQu7r/iYcNRm+qMSX9+A2mXurGwTdb2BzxSYxaSqF
uaSNc7yhxmNsXuxw/P6qevFV2R+AVVVHuV9SP+kW6rg/ZbOoO5ba340bGErB22qjiRrAinATb7qh
I2oy1S0mKC+1oHlR4ydZsMNVteWgXnyGPPFNFNtTaAb9PhH/an5plHtCbFwcULLryZUyyzl0322l
n+Aemgh51m+ftadtT+3Sd826hM0IKWRTlWT+i3JkeiJUEXpeaWdMXNCinUpU4z9cyAZg2IJxsevZ
zEAKi1uAhq3ndXb9/8gYBROZ9Qp8UfPBqbng/EVnDAEE0cTRFwsG7yJcWV9QzvX9Zn26DjkyRDGQ
p6hZEt54tD6wQ7KUEUdnZioFz/1DIp/3mlwgEBngVA4z/MRfPwM7/n/jMpyQrm4814T9tDCiZpcA
M/PBPpok0++/lnBHtCzxjAC2YVinBeaOfv/YGqHW5Msn1EHCyC7MofO7QBMU0t9GFvMzi1NEAunf
9/Wv41t972Bh4B0buap1PRNesgbXpsA+K1lQhCXri6aLBdznYiE2FNhVIWQUPedJi4DxgDbYk4eJ
x4uHulcxlo23rWpWmsqS1VQlSTYNO4ibZnxzx28PA6Fjocx8y0pKus58nsL8UT8iapDUgodIsz2/
UC9aEYIcne+kL1/xkyBrDEi7fjnXKCx6XEt6C8rk83WKBYxFyNyT+N18Gie+G/wN1iYauYxtp7xR
KVQ4qrSurmzW2Pn443jmGrCPTqWbAQvZm5JrGd3cpjz3Y1pcemUgNvMRFHmM6Lr6ArzKgsNcgQXs
l23p/RupThsoCD8BdifdVUEJi3pLwY5J6cmvoF5kmLmZPVXFanV/vHAu5t6Hgfd6qBEce/nP19uv
IAYSfmRRlbP1X5uUVI6R7/8qsNGYNOP7qNBieeeOXt+A1OA1EP2qMl6Shs6U7bwAs6Vdf31Y39ak
wmtVCU/Gkf2t4UWgG+vX095PqkBzzGzNnDQJPDai8qiegj/jvOjcgX8ADh6IMOwM/awu3w2nZ/Sk
RCr5SFJtrojwb5Kq8hKDkqfzqiKBMte5HGdosj61eKcAHGTnxlHGHDlyLrdEw/QiPJK6IB68CqN9
T+dBJLfc5BP6urla4ji8YZ8YlhKpe6KIe+JF3lpOGYuv0riGTS8U7TXR6QzOyU52fRGb69saVSRj
tXyOtejjQCVFJIEm3Xe+NiYsJdZGEjv8NeJY1nOLd3c1LkM9/Yu45DSNMGFuK+W1c3Y2jEvbHdAS
YXkp2KkwG/T0zR3FnG0F39FGaC/Pr9nxZGh5Y5TMgDmT3FedhEuglWycoA66f95fxCMH3jQFSQ81
u5Wen8ZnlDX4dhNmncXtMMi28HviTesjRBB3JoNNTlro4cpC/M+BTMCiNYmyvmZAFbXWS9zFnMG8
yRkq+vDMhUUSdhjjQTGPXBJR+YPo7RlnGZFLT+fBKq0wEm0MIZW/xcXl0TPTLz2lVidKp0ATGman
LcD4u56ZLXlZ2BuSo4DBQH3X5vS7hpTfaMcXTEtjNsNfvNSl1AEI4cibq+TSl0vkd4ckYNij/l+P
DS+ZToUTbkdAD41e2fjMgi4ThAZcPLEISj5BO+mwheofAI5cTurXWB1+KoyvqLoklrZnc79zuM7b
zR5eRkTo/EpO+7PK2uUG0vqE21aKnrNeHfYu/ioD8AKwNJy72MSWYkk3WLr1b2NfJ8LVHFKVo5yL
ESApa4ZCrgdlTwPkKUhEM7Gp3iUz5um7o/HW0RLL3MVDUZe/EAlaoGcAOX5n/8GjJoxA8IiDXaaI
FP6LzoqBPePj4faDV58c8M2I98iKy/llgyO3Q+g+J4TMlaLu6Wl6rGhOeB91JEcDG6E5xr+sh1fY
2ABY0lEZNSBwZ+cUScJ8WWY8TeHg3/PX5O9VsqQwIGBXelcIIMW40cVwM3lRAP/R6VGsjTqIJ/ub
P8HS8vWZTCbVZifI2VX+pyoAIWBcf1orEFfscmms0jwraKfH4OMZMpMkOTar1PuecXMhaEKchHkM
np/RBJNk6BwlMmtXbnhnHqzAMyKz3Tapx/IzDQHRItoDOXmHpb6kwbNLl+B1cO5qunP7sAuoWwCo
UAXANba5jJqGlR3hlJQuGs1W2UGly++2bOsy39UPwT86L0XkKZPX8iI//Wnz8Otfnw56wqs3Mnca
YuVb7ayVZ6qDEJom7OHEuS0gjyKD2lqsUUOBTIiETE9dS9SJF8qlLDLTkSUlpqmGxcEdi9cGmxib
L57r8uFuGN4kNWLtII0t8DzY+9WTtKhAK2U76Vr1ojqRyMVKgP4QxAMqH5tWigmes4DhfnGn4WG1
ngpQo5EX3qgEMxxMuiYdGjlYJ59N4xMinB6cGHCbqrPPM56OwLy2NvMa5uv80AcFCq71Xap/ZSbT
214YM70IeayUvea4WX9a4NM/UdCSCvu9M7RV5z1sFvKERvn7jarfdXYShkbt47cPs6TiW5h+9EWk
T0rWVU5Fmq/ERBxHc1eBhzjfOKPF6FecS6BsUXi+ZotkkGOo40JwQgLKrfE8iTKPDtIsAhxXmBKu
atshY5FgnpV8IPMLUdduU/h3rWKIig7W2D+/1vVEqja7KlSsMmUDHadqoK7T+QUhbg9X7J6LNIzu
zMUSyfTekIACn0sFZ24JEmPtYkFOcWw67ms+fJsSuqV5hsLxy0Hrjb2GmUg84fR4OYu11VGKyzQi
NNXoS5eoZ54/jLcEfbDqJD2vMdPHsWDcIh5dLyokMuwueQZ+CMvewnZVWKcsHGZvQznpMdlidYkE
GRtinDv0yEGKfs3gZjGFi/MU24iDgDt5mLRECJyW9U4eAoWB69gLqGn25j1TxV6e4i3BydPxn/uv
ZMb7gXo00d+pA9fX3JLVU8Xsk/zrun4/0Uw6DppqhABXpQj91PNgaLyiwy1pTPW9Zk1SHmPMdMUd
dcKlHEnrRsdYQtKC1OeZvEOA+fBO98PVY2yNkH8F0kj9WOsPB6KEL+D8lZWUNZzyv6NpDeLCZu4v
fOX7AVwFmt9Nej56MxZ5enoV1i5h/FpX+Z3DtjImQHlpBrCiYmQnp2AfxOjIvgJw0hfc2KKoksp7
9JGSvFeM5xC3l6qS0paSGNzHzNCWaVft3mk8e9aUuXwCGXs//TgWofkNXaLjR8H+6AWQuQXYTSy1
hqmm9Zxn6C+gNGq7wgv/R+LE9Ta42kFdYz49dgWwrvo5N1lGf57toHxLJRyPjlc5WPQsq6wVRVtM
MpY4JLTBjnwLKWXSjGZks6g++UmuX28AETFu1iGOyDLgvkoYF7s+bYX1e97vG5IHvrZw+x9E2Smq
xryi0/0MQLaU0AOniKM1VID9gHzGjXANDLYNoHxizAK36bZqZLnXBFS8BWS9kb0MWxqLyzmoxOAh
lKJn+mUHpcH9OqaY1iL73YaGIZpObyEQw9pY6rxoKgTvdlOQQBdSLrdN+HjneWnDjzAnAP6i1pb1
m1sq8a8PnsPg0XmkqNnQNr6AOfImwC8tB+3zmLkNPDSBsPnadWPOx0crfKk9jc5XPNP0z9PvOyLF
XQOQCYQ9ar2JW5uf/EIZTnvXGpCcAuM9BMkYDzk7oTiMMJPqwbPM8SmNBJvD+FlnTN0n9VxNvmwb
SGrdjy8Oozz2moJQzNYdo31WvM3QzwmJWKx4CBNuvmaJ++6+xhfwJJ22jA42i78bCfKrY/xR08ke
Of+vO+u/E3zF4l1ocQ9TN9/w6IlBHh55Lyvvuzc2ORd+AI77AA5jXXO/PpayCseMg7o3PgE8Rkyz
it3T1Qk2IQa+CLOY9zmt4oeolu/4tnrE36eQ2XHgvsdr9/NjWTKYejgInuYOZRHeyHjMNIfQCQeG
NBBF2+vBl+9wW8hkpcgNgMJnWCFMqefP6alseOKhkQDdfPZTvRO7UYWhIlLMqlCsnOaapVGcgbgk
9dcq5XRpxNBSW20qDroMzi8TUQ5hUDwP8yP9gXxDlMugn/DGKwBDb4y9hNhGffrYHjL6hLzICCCv
+oG2wMMhfbRpJaoDajEauhnHVVxDXchoEwo2os1u7vWeqL0ENLk5HGKPGcNfYcG+yTkiuR3B2R3X
9IW1JAicJQiEjNhQ/3yPD08d2tIBKOBvyeRjNWjA8Auf9E4xUW/bs53grQ4ws+HBSIAFknSCIDRH
kygsJG78vmgz00asSHnS1jGQFs4/BFfu/I+IQSTxHZlq79KaKJHkhEVKC+nqU20pKGjnR2M3fV9b
/tSSqGL8kJEUuKR9VWa+x9tcPCLk2VTWCHRoIoTCZ1XVqe2MQKBxJpdowGPMai3VtH8W0zaH0+S4
dxX2/J5i7To6CAoDf54r7fOMEVefqjzsAMP/3sVJtxHq/DtR785SUyBbhSg8xRHipc3KwWOy5KzF
I0bALluzQBtfWWLhNibnjnbqhnjZm+SlF9RuFL2p0yJeH9CLgk180Bqi2wlD3sB0TBLMCBgW1c8/
r33+rrxEC7hjaH0Ov55Y6NzqTb3G8wVVdE8GgAdT2H5gxZeS9W4PEHeaIlUGETH29x7SWiTft+1K
zVEvBTsptbCoHwxt2lidPfs+9uMfqP7KkOhLhhCQDOhARoGBcFhqgq2MLfV9y9YvgK55ZJDCJPjZ
UlZI6ag22xk9VYZIQ88iRoYoZrBrF5/reCHrFHtVLboZTPhoRpP5MjmHMCZn+g8bWBxZpKdTQlKd
EVEHEXFjt16YyFSKThTA8m2oAY9DKwhX60Q16c9hewbspFVmUuvkQKBjy91W5qX9BWQ8kTLYMBNF
i+SFvzYtYZwLAR+HtCZfgrZ9iiawIunrS0VFKKq7UdR31ReYEoAW1TPT27u0IWGbrXyH4OhfRUod
jQNDYG9PMJnVBewm/EfXcKTMCT3viG0kDw1prAlCUmgI4HMib1Mhbyms4G6vJOaVDgtMGzk4q6W8
rWfo/TdeEENhVWBG0bYTEWEM6uPf+99Zfc43ri/B26i1mWWrlLbX+ZOZBuyggMRwCmOdpaky/U4I
uQy77BhX0GvU8wmetXUyC4b2Rmu4PO6diyCiblMIEToBejfK36sMU5IhHj7+zy4OeokVqm73cNSc
ZzQ8O5SSO72Pzzs02C4tZC6RhD+xDH6I327B9F/QQoCIrpzVVWJpXGcGMV9Kl+W1F3MDIASOZ4pB
Ptz9c2F7JJv4q0G1nfbGA/AWiSLFJwbGoQ3lTuCtLZZtffTcYMKgAacsoRIOep7SsMy3psYoCyyi
9fPjH/DqAtsq7s9zSWqGHAf8vgKLFcib1uyMjz9/npARUpHpy7kSXB/EKiWEY1GA2AbvvAXHO328
ebK7+fpcWlGNCCR0OvJzDOmcqzqmlJ2KiYPp2WyZPXhVUOmJHwglbOipEdmnln1cWCf3i/+F0VWo
lg4ssU13YlEprCnxZLuSrCiOdXbtSprbl4HqPkeHdkkYnGcUZqA/KMJDGE4oMQ6bC7wAOehf4jx9
S6IPtLYNzqQaYmvFpkzXTN+hUusq0Jth2t6Mq+MaktOuQ4e+HWaRlIFsUFG/IGaINsH88d2K8tDJ
jdNvlvW0mhfwTH61crrYqfGcm4GDn9YwxTNjzIFEL45kxsSl96hMYjYvhu6Vq7LpJO+DI9q7RtEE
opPqIVhD+eBMEqRaGKbm17UFQOYgQ3xKQCva43hm1UUfiVt//KT2tCZjgo+DcgQ5bHpdrHceikw8
Qo8Ff+O/yuCUWhgnZn5QFpC7hucpfvIHmoD399w4nkw8CaA8rxLAOdnN/UpFWady5cPeYuMUeC+O
fhqEL86tpln4JiALSSC8OJ0lZPx9RG71twuSCWMvb/7cNwaAgKrqasBrbsXv0TfQbZ7YTcqOD1Yg
4UgZa1MrF9MoVqfWTgicf/WR9GblTagav8B8eKeaE+zCb8TJ4tXXMOxY2FkSDE4NoSy31yb3Vtb2
7yZBBjfDN+SnItqcyC6+fbJlLVfpOhyRBVCIrrOPHmI+v1dRaxJ8hkdwDsSv8Ho/yRMe/aXXiI68
/1TgjxhiUELocUe1U1U9u9IDC+HRDSkeOLZJiTPgR3KDKkH0wIkgCCPxCQ7sVLQCAFRKEq7A9Eso
6Ec6DLdzFpItN0xfSvj+gprxHKFSnd5yCmxgbHzN3NsNc5OsFWQ1icDGF4MnmoQMAHnc/Ca09QCz
LDoZbjq90MxAXAPXsmwVZgBkPeFO5URmfLFldjfD/8uI/5v1moSvcZ4CeB9JNo88912lDlIn0TkQ
B1waTgsb7z5P1pO4Br/rewgMqBLsiHK9EPjvCsTmYEYsNuCTaDOSB+HteLfgBetcQq3bCBs4wp0U
dhzdGdU2iC8s+69uCihs3Q6zmPwGou+Lb7bJdcsGkRuvWueGqwcBuWL71MPicYUDsCxXMgI41Vam
RbcqXNRQ0qGAmJ6phex6ev0tSjyxYV8p6aAbZXdkJ2hWGty5vkixm1sQAw+UFa6H15pThixtmDXh
kb/d9XydME/FROR51ibqLxzkNRopCaqVVKcvK+FfPEs4ePODJzEiZeVUcyJzyotT8t2VlSsCnwVA
CbFcpNPjcFZayfS6hMZhKZ2T19DD5QfW85yIMpIri+IJ+zXHLpmDfZGSMKmu7BEOSGVC+cM4m9PK
jpSbrl4MR9jhbMOhY6g0oxlcLR3lANPTDP+IG08KjGBWVN67b+S6833/zAciFVzOBm8ZF278NPQ8
j1C8LEiiVL12PwSoO0c51/TKzMTDxCB607isqBcZKLTZXaphULQz97ZtAZFVJY/3KEDIsnw4wWx/
4ed1CwwD9uGd8a6HbS8j10RGRl5joRE9bGtqb+FYlQshHVgsVE3ygR5mY7t/1L0A54TqlWyDJjyt
Y0MJq79yZ7MnXi+S3uRQ/tu/h/p2a3YjSAiOZcY+EgzprrArG4Fl8FwrXtgTUfR8fCaRgqmjJtQK
yu6crGqOjcPEmkIzYhDDpVciQAmdlGoOZYHAjv/+K4EQk2JslUTVg8SuDwWAf4M54IzTS9WU6GQb
gTEe9nMbElAhEYL3V7ylqwfcsluyGlPp9kMwkjtWehzTZNDAcWOd5KLKfw3zE91ApoKeLKyhYcO4
ZxcPeQga1xzLt25Pnqiu0ryc+MmGYHtbnXFq9rGhcFmNBAUwPfYbTicXb+/X3VKAF/+/tq6DT0Zs
KvFG+yQI1kjUVGExm2JbykmMBEFEu6u2zzi8KmWmt9MBnihzNsGSjD8gf7A1bkNxGD4qM30d7yMP
kq2OZOsPAumHIlq8P6oq5FxfU16FenfM/TiB7VM12mytqa9dZ0VoHViHvwA+5yUJjTp/JV2xGmfP
XGKxfTf7lhXPlmEfMaYJownUrtlHPZTPU8xWThL0hNYK7i3PolUAbdJzDaCdf/Elv9abNWgdpxKk
RP7Hqns0GXT0vR24bFYKHfjlbLgPRI6bQA5EpwYfDch3ZZ3mOwwTY22wKKYtlZBEB3rcyqQqOArs
vWxafBQSI0YTO7d2fIpjzhcBw1smfEK171Z2SR70F4ctcjrdtPVYdTfUffg+DYU+TJuHSY9PI2gw
NVUoli/cmTFZE5e5k+n0ZCSWl2HjrST6015tXSANyYm+BtCTmBJZ16k9xrVmovdypbqttsESt6su
j4S1LIeTYni6K5S6t2+sgWX9Xbr620Yfw6zhLQ8gw1c8hhQz8dmDPilGDwDKUhoufYIKvtWW/34N
SexwoGFzZP6fzv76pCvDZ1UHU1oncWrZacjlQxVKTZjyBaOitBRvGvm/plWab6ZcIVz0Eur7cz/w
4+Kl2mMK+xzn1nAvb2267oZTdD3Z6EqDJDP2mMI467dfVUi0w69uRTeE+Fjdup15YsGPyPtCaqB6
NZbRQYPsRND4IVM3DvoC4RGNFSxtHn2bNEb8mNhdMVUskzWZUKpZvEPYOTHawK8bP3icS4F8uZw4
ADHGR0Vm6ab1zHUxUifSXLxGV6eIEvWuLW8RCTxegteZkwUWg6srjzwewTbJ7+dhck77TYf4PmfE
NCg8C4ASnezCxXrNJzUfzKMc9kv3Bpt47PO6QjTnUuO8ChXw2nQ2X/qLNN9E9XW5QQNxUf9L1HEh
X1gTtMdYUAawkvoVxZIu7tqOIIkEE5Ujg9qZrb0/8Rdsq66PlTHQxvD9BTDj1gdXpO3qy1/3OvaP
8GYqbYFiBZCYG+7+bKP88DknTb2Y4Ll32NAHopLay7CB6kdhqFqk/OUeQinPN9BEEec5P4z7EqjH
NEdRXnMvb3c2w6cf71maQf4hz4Xh3MOgQh7uJV3Igv3498nukQVhOJidQwwKv91jUdVYTH5Hw6SM
oaKLfnEyjfBF6pj54dPN929ISpLZGTAfPUsQVl/PlHaR7iL55F0cBRDr7VggwD39tgQWUy3O5lVo
rAJc/PChwzdn0tacabeifVhzy0sQWHeBz/78mrXvgzAYSgQSPStvueOoxhoUAqESRjtgFiAGrsYh
pdr131xm7HJEjLHINC0+omap/yNQYaqk/sx3Rv2PljaZ3Wl3xPd9j9ri79VGfPK/UWQubEmo1VvD
OcoZYnvC8WIFwTqH7LXgPMNTv15aKZhOaOvtpddrGHu52X/1rsRwPF4hC/ub1lKRX8ZJSVKBmVDJ
qlTn6Wm6ITrK2AiddaElGeNGCeAAUNOXkI7mQccIwVBlSjf5k+JpAGHDFt5Mu+b67H16F1mn5NyW
F9vb+h/y7lWc7vanb0WSuU+Mxzpt+1DeSysqvTs0I+B4Ub6VbHYzwKNIAZdkGmN9GbsGUS82HuZG
WsP9mieoRHdI0B8I92yh50pjUk6GpNgtrqjZ6ESUu5NwFKv+AzW8lrFSdvomRNG3Wo7WP/Hsvrev
v11ZGj5Efuxishkz3OKUO4OizbEiKBFps74fJbypI8z8qZWPLRsiswH4KHf3sW+l9ybVpOzTf3Ag
0z/jtMrZoKheXuElnlbZWVwu513YkGe2xnmLJT1MFD71Vnb3tEIniOKHSC4ArQFtf+8wbAC77nDl
P0J2Ac7F+GsarhMLg/ouicK8qdlmi/TCbV+gVVF9+V1TbZ+Mrw1SvTTH7+zM0hmQY+NtI1e12IKz
fVdvnv3ne1QcLpoNNbby+fqsNX6qhfsvWv7sq228s1lfIU6DXA3PLUGqAj9GOSeHUOAfdsr2914J
UaC58O+j48YgL1EWoAvSg8oLAiE/LqpvljaV2kiEmwPaWM0KWpfRTyfkFpT5KTrFBDyyFgnkylQH
fb5VMUngmrkrOOChlXp6f9reltoARYnRuJjXEBUIicdG9RCR3d68AAaQeU3PWrDzzpVXNbVbkc1j
6ldBPznuYuBJnO+DpmmUAnRVHZguEv05ssFj7H5G9vtDV1L/wR+ZjYxV+xcFZ22j1r2uxjq7QnHt
5+zurNzFlLGelZzX/Iw/Ij3Dyb3NYg7ZB721GEN8nXfaMg/RZ4jNP5GHSLyeSAObcIfu3KdvFb+f
2qBU7XIceKGFVNKPCMEYnyW9pEhSbmJHwhTKN+9EMv6ERtDk/hsRRw5kzpAe6GBYgDHn9j/Xl0CE
C5qF1Jr8/jGwF7Y9JGPLzUa7FIGKykJdJHWUMvN7jsikTxJvAKPjxhLGVZEpQDTRAnqZkMuW0Rln
wMXXdbLhlYFLJFm3ij+h5rXKOauYYNcRfzeFacAMQKghJaZLXhFIUZFvc4POcXj0xm4JR6bJrcZ5
Syz4W3vcNGn6l2w7OOzKNbFAtBMmTvXOHvEzNIFv8EceSBjegUsrSZrpTTgCp3cveVI0HP5UYTFf
YSjtNUAYozDdMa2Xa6oZ7UjXa9h+yrIGZOXsekNE82U7MhUx5XEHykwdLB8kiB2EsHPyOffC6oWx
9PTTOfA1AWmWKnsO9mCLyeJxRJmI/waLheIvXab9vtOX6IB5FKR8elJqF+f5TyNYdwVCOflfqnp7
Ik/vTE4gw/yalct9goXt2XPARKzINf8gGPYHcQ3Bwkj+7qfI/GYCQTu65wJL1dcmbtwAz6kMnEcm
8J0Lg/wWVCPV/ep4d4MCu2YNlYxpUN3lqijxTSLkflOqhDwHNC60b3pMEYvbcqBTrvl3cIIDwGwq
x7/Ka3FGAoy3/BxfzDKdtMjH0ru8Ksy0dEEmGTjxBNOHAukxugPnZF+HGZ9oWwGUm4N5w8ljfore
x5lncOuTi9GuZgMHmZNbEGgyVNj2cRCRFAODdt87SMRNZ3H4CmfxoqT3/0FnPBOARLPWl6eoyBn+
Y+ika5Qg65e8k7AUheCAxA2xYsWkHaw993AYcQC2Y5et7CcaY1xTgVy+BsT77VKe4YoVSMrQIOGh
FVQqyTLIuLjeUS+23jU4pis8CTm4bh1MWCwquGfJooM7d8gu+Zg8l6xYz11vFVGbw9L+YqiquRwJ
z6Gbq6nR05UHJQW36UDJUgFqs4TnT5km1x5kYqO9buLUbGUbkXKwJD9gQzYht0bkoGsx8/zkxVCU
aMYVd/iJIOHq1YAdrfJZ990zEtfdhzKA91PIaSEOEKrWKMpX9OScVRnbAVLhB5uT/vcWMgQwsfzE
wLR8QWwevsgYEH1KaU6zcXM5p7lwAiFbRIK+boJU3Z/xWRlioh+HohpqBVz0NAEnHZCIE7BJVL0z
URJzrmyjWBx1P935A0EDJoLTH1Sl+RlV066OhDSs9rgOZ8L2EUT6oOrXJhTVLRfGyTZoBfVkSMzH
fR8gv+LcxxoHx7FoDvTCA8CqS2uT5R+NBS5VoYsB4yKUdGpZ9hn1aeCnDviVuRs87WaFe+K3T6kZ
QERDhyVOe9s4OS3O0TvopGZT7dttJCWgrHQaUxcvIcjzw5VlZMhun4RyJQrgdjmitwr/u9TZctz2
6e0v6w6wiM6AwqnFspqxDy2NeN/EVqqov7gZk+J689M/MoyHTcx7NNzTqQsy6tI33wbgFbAEsCf7
pzBTW5qQBwK8PSPFC1PpaLjMeHPpjvSTrlXmwtdmBp4I6hcJ0xmqj2toiwDabcEU3Cu4xAccgqVe
KLtl/wwV8KxGx2Ksfazfd5aZ9CsOrEpRKVog42Gocc9RT7XtCi/2IfmWvWcY/efATa1WTkvaXjQM
3luX6qwf8QSMlnSTHYVroEjys9GsU0HlInmrxafAw+Tx+8dHqt913LnKRo/cVsAg4VoP02Y2MQOn
VCl8qXhzFiV7Sj2FK3Ohu/vAbvXg44mNbSxmC2ndgKNplvG3IWX76GkeXN6XCyTQbTxVQjk6MdxV
C3ox3qKlcJM+PsILaLcQF9C+kqPU4ca3Iy1Hd+vtEFh3xhJwdgwEwJmzGMDsBc4gGzKQvuaJ/iRu
9C3/dvwFC/bq9aRy6Z02ZIy3eXJFBoGv5bRuDEqgYEFI5+xLVzkPOOndxSe1ivbw8merW9zeQ8rf
zy/peJDbubEmrg9Z6DFD2Z47gG6K9b1b6RlR+g+dpKIE/wvtkKiAZ7+BtuoT0RHTyt6rvoP32cRW
hXPDX1opsxJ1SbdF82TfWzfPrBdPMm/u5qUKJ0vzSnPD+yXS1izwDZbO5wuWPGcI0IQfx4W5UEOm
eDm7u5maxn8+RtWkTY4q6R7Yod/+nWZbML4hYWwO+toCE14sbOPmCJk6Svb8XwS7kWrKfQ44G7mH
IO9bEGf2b7V5e/0H1gTTh1g5Q66iZc9wGZSOv2dIonNxh4gY5TrOHFt06wITOjdVnrpIniGRjO+w
EYTUWxSFsT2A8+e+6uZAMjEm0eH3MnIQfCsS0/g+8jmOG+H2T9pHKkoCcSjUdn+p3Z+HMe31lNzP
NUE1i/D5Y7//W8g6N2+RYY9hdwF71h7Y3snz6JViFnteEyWYEqGBEs8lLo8LzJ3dB5DQaxoivm2Q
Kmi+L7zauA1xgedizMiSCSFms3si4AYZTsgpq8ylot7MnnU37q58Acz2tz4ZvRR6fYlTpQKj7olt
fKxqSxBIoTzQydjBonI1SsHRNvuKZSZrtPF4g9gHdyec8dIYnwdNS64a3Lj17J96Fg8Fn8sqo61/
r30/nWXBI3kTShxncOJOZL4qRUw+IDs2/qGe/2s747t6wLY+DdjL4oV4vmTILjUUiyt/aJ0Ube9I
mgChjrVmFALJpvbkby1JG8s6BEvY3AURVsfkCCt7Q877eIY0wCQ6kou7oOvzOW0nOhGWPZJoFeUT
DNZK0WDDJbptJCr+Gm5BZeJCimaME+gHqNDRCQaGwHFzqgcfe6J/i++ia16iafsJEGyBSwg8eAgv
gwTpkZOnbt4hJ8dnHLjxjc/UN28wI4b52GVo1eVe7Ac3bghT8GpclwzjFKKeGJPwgpoWvjDYFA+t
Cj1dlw1WpYQudCJ9F23DJhx5bffISbw+349IYqyNJ06U+4v0tud7gbMzIb3AXTHA2yFYFfJNjB8j
OAu4v49cIuiKrbAPo2K9MDUUcK5Dh9jL+Fn/wsoUMDc6TPC4cJS+b7yZTXMsB0akKgCaxvJwB3js
NHxIDd8aIeZizzKxgpw5q/VjPt6CV+nmTFU2qwAnykxbOZ0oHI2ulm993cMQrNdKhKszCdhLjIyK
fSevZGV9ndbj9DICgXxqJxi+AzeElz6N1qbSNbmhp9yzNGGtVpZBkqBqhEOojHxqDFaRcQec34X4
4ecj5QEjvMgKhv0s6XxYuSUQ3Qbajm3z7ECGRjAdRPjBuy0eOzTzgvgfQhSod2bJWbPbakKRbdJS
r8/U+0WqbUoho0sVGD8GhHcUwM9EB08iozBmc+p/fweWgO9WIFV4bGX8F6hG2ssvi6HsPVCn1JA9
/MM/peP9ur7jPSZUCOFGc7Vm8MsHl+UMfKxGLT0WVjOSAZNBLvkDkEti6JIcYpRMvB4+VSXDTx1d
gZOw4Bk2c/c6tmTDzMUC4Lq7/wR3r1/LHZwQk8C0ApVdyME6Fs58gO8acnI3Q1vwesCOST3o8l/w
pRZgUIGEFf1XIK7tNgCeyUkHiLo7O+g6kPOwrO5WYa4DUSYo5FyUQiGI8p4fCr3JfV7unNl5A2Bf
c8jdFlVEoxxHgT3jruAmJXwNpye2h6tmRIYPIjCiXT/Pyj4KlE33sLxW2Na759Q86WUIVr+bf610
MvT4GRVih/tNFEKQyr4B690rbhqGwUyVokUG1OZa0selKjTS4XwrqO1ENS67x3fucp+PPTvXWdY/
lmB5LOwUd6uFMsduBuPIkbhxafs58guq1TnOCu3EshdQxSJGbswbXgMskWcrIitm/ZhL5/reyTT3
baBpvg5VtDI3kt/Lwz2TNeMR0J8ZxXovvyXF0fZx8665stJTr164ghcR0xQxWVX4pRX3VX3Pm3Fm
+2oYLtenRgwsgZgEh4xUXBFxA2YjfcgLD+VbPlSYPsQM2uG3qzObPemtWlFcEEnRIxASAFlB7ENP
Yoy/sJ4B/AQPG8Ezgqgv6eUPhztRgdA6wEN1JuFMKBNoJnv39cuk1jFoaSNANA6yxesQGGFwx86t
643CEbRNR4UrKVdNIAS+lZ6SBHfiAEI6FMfR30/veSDlyjacdBz4LLpL+C3hTJLmO3q/0bO5Vv7+
NxqD+MQQ5a41Mbpb4e74N2St5HYOTQDqMdohLpINF0B13tBSNiFf+e6XXoPHuK7qECPujB0dRA4V
7jBwio1BZy/J7CCSWhuoeBAsDcIYqkodncj1DIi8nLSj9bcEtshzuaO1tlX3yxkETqCls3dueizB
slDhMgeZWfPBTaCY79BSDFtsTbSo8+TovFJIbVa9ClE/FyJMhUg/lgx4X9hDalfa/4EN/gykKuU/
hb8RZGAuk9LnDhAkAhf1ccIFpLrJe0Q9hwUQUF4PSvVHeGn64v8EJQICXbaNLcMH7UQePA2ACAtN
mdMX6tOi231OSGn2oGGWUsIUBzG8C+1GYKLHuTf4d0qd5+CZbBQ+nNW/BkCEkHd8E9j4K1JY6l/A
Z/Gh7UIlDQLcWVy6gS5uWNdi8k110xiPp6BFsqfhK1ZK0V0ahbLapa2gpD22ofDCWCDBJ3fEj1M4
oRAqcDS/Hw5rNHp5CwaupjKzRRCYyhFjyrbWtFWAwZcbW8oN0xsKp6c626JIV37CO5yw+BjuBgHt
3weDDvB8hL2Fw4Bh9EqAgMaEFUIFO6XLQSCNVRH9Oagiv6DsKRBpCL1nWkdD8v9RrNbWUesxNeld
AbyTBIT8hWW3NgTqtzmjzRq/81tTb2x5LK0HHxjvQb4i2OY70ygtNl5M/xmrpZwgAFMLctUmB8by
N5oPWR1t1x/EeHqtECYLfPjknC2s+12dm6VUhbR7v7LCOhP/DqZ/KVixDNK2sPGgy30QHtyVrK+T
vUtJkWKTal4npkSrhIvkxuj+cE/AkanwsH4SbFwGPp+XNRSt1fO+t2t1pnxfbItzEsbjr+5WRWYm
FgZHysb51vZ3CIQits/7ennm7KFduy8pcygdzW8mronivVLlMLKMswXRzGGLsWhbd0nuvTcyKIC6
/hav47DRhbadYkjOHqoJxzouj5VN8PrjiH2H0T1qOckZzmv8/f7G9yjx7rpa6I1ZCRH07P8QJj3a
rFDtoHqNDEomD6QVCShyvQrEuOLU+ZHpNcLj0q1Rs3o0viXNoWoI6EI6Ujh/lc2VLdqkPn0ESgdb
2B5YooMLSaPiQO9v2Emz8EF+2ssKOb/POCyExYiipZyLQHePPLqwB7+MH6Ss0EEf2h/oUq5DfovX
/TDyb/I+U75AMYGm/TUbkEBHoetJY+S8veJGhqgZHCv7x0P9OVRUdc0D/A24GfGu+KuG26ML0X6M
TsxUBWLVBMW511KsHpt0fjLFkdS1UaFO+BEYUwKNlC58/HVj0+RpMIygtYXnrpoDB5XK6lZV6yJt
467TDkNFsXOitFZlCFY7I6bG242jBVqdt7Ohmu2KkstjUKVJYzQ+O0moN91AsSTgIsKO7xxPmpRD
W+nuCWHnkopbyRzlQoKa4wkuRQTVC+lC0q3pDN35dTHwhE55/yGkj4akBm8pkAygyAYRCU0uu6ic
dCAfIoLKkAHZT59dNNbz8linPngzZRu71Bl9n7WJeFoVWlOJKDrEJ84t1MOEdy6pUsSKqLUrTPOC
lgFLcJ6Aq47edXLxjZrqwq6bJBCw0Ex6HIKOjhrEXHR852euh8ehbiOzE0bvAP9NBH8dNZ+v0E1a
ztil/s+qYeeghGxDs1yHHBKOnBIpiLd1Nb6OrbghitQEgIk2Lx0ABOkZ1ENkPTV6OpJfXy++uwhl
8vdkAzyjSeMDY7rT6enK9ZqLE2JwMYd+8d/bK9fcLr7oLs94T0qyvorD17t6cX3+kkZK7DiAyAdv
OJ3f5tzhL6aD/wEvOdx2on2qlx4EXs/5OAGA0mrQ3adcwcTjttA6ed64AsDXHUrH4zDQ6jUgCQtu
SPAeqOh/YEoN2iz66s8x04XjY1ky6IE0wjSpVwJYU763qv55cwyLIQ4XWpw3uaTrfShqaxTN9ia4
3uY9KxMIbR+fPkOag+R1MYMJZ8f95aff+uw+l4fKhesMAtJCsszVwxxPl5pItBDKDFq7L+hpGNH6
olu286ci5PAk48b4LVAsR46TxA93m68vFBWWsZf+PQ1GoZ8BEFjAygfI/pJCQIg4JQ3b31GtWb1g
VGoC/xMpYi7aM24AQdaSleVBfLwGnx1eRdv50frdt3vuHXTX1zeznPnYYr01CsPYmL/6/mfCFk6E
r4Oj9Fr0GoL9uufHRh/0iXndtR0Wms+R/nagornhNsTqquWWApjsbFOPS4OgKU3ufa7kRp/Rvfuu
Af1cw9rF31WMQho0xcxDb+ePEyPRRIPw2f95sZqfSgFWJT2kMcclqn9KTi4yDhsALdhFMzeTQnsR
6Px0bdw9XIHXS3KWtcJjya8A1Cx/cbgG2GFWJBNAUYqspAe0FUoVbD29uFheV3eu4a+OPgzOyWnS
OhcVL84O8axbCjpCao4IdFumI0OkPbPTTiMBpbTm+ExPs5gmxUNzvYXFB1yiEuStCOwsmRgrTzcy
q2VufIK4E7fbZc/ERW7Iq4sCawS3hSOqvLTWnYUKcM97k0e0UhG1+v7/sLsL4iOFF1at1AaJtqy0
KF1d4/4hlrbPqB3RLZbGaQPjzWgl8ppzPhwqBxTaceAaj04SBIl6zlp8l+xn/uzxuxs4+XNGOMC+
Y66HHasxe2cKnRkTK3vDOpPWyKzBZmrtqBLyQOsEi75Q0rhfd0NphuB0PkalF8c/Zq/cVzD67mhO
kv0sXHMzoV8eGMkJTFYe270fxhJD6O6TYz0p0u5Ee4JuMmML1FuKOi54xbbnuwNYa5fTGGWDvbdx
fIJCSqbSlZ1CKRKRLvX0oEdPAhnonSadFUGj4Tvz9ld1TrHMd/AStozrob8K/O5P8WqPXMEd6Ps5
t+vFRGv0boKZBs3ykgZ1B0u7Q5+NxFXRBoQeUc9Mnqy+UJUKoPnr/cDcsWxyVX20++gTM0q3qe1v
gLB0Q0A4RpkJMrQekHhKf0W8p947dyhEZBE8AvX45CQ7NtU7BbMJyUd5paBF4/z2moIw9BgQci1t
xukwhFrcbh3QMXNuMMJwJIW3PwyK9NI9u+kqw4fT/0hLD++ZlINWpbwNnF/oiUMz0N3hMrlt9MlP
rLFVQlq8aK1jBdrO3z5DQwA7gfQvjHypuvH2AIyANF9OpLB6h9n1WzTSbktUj0yeW1vbLOkg+NnT
GftsCqU1Orn0Sz6sYCdivVtfc1zGSX8n5Upsldc7iJ55W+r35iZydX3GhGBKog2lFvoU8RtW+++k
/tz55WxHfhvlqYipKzSV5BpUgGXWFZYc/W1zXK1h0UBIbH0PT0Jk3K/ojZV0nnXXVHypWfFDLPU4
zUgGa8AOdxiE3dteDlssiSlwS4gB3Kh4II6mgwWeeqTiGr9wf/D2HWGLPQwgoTs6+BO3YH691H/g
6ga18P5vWF+pA3LiALlORzgI9kt6ezEHniQEAuZg0ZnsCrgS41K3UAnUXXEaLMe+f7yhexePm624
xLcyA1zENU1kPtd/ReDw/nBZbmYMQQmOXmxFdr4Uum6QKqKx3Jz1zQEehjbND7rm6hF0EUnESv6p
GqYgu6zwB/Lo0G1nhXQ9d2JG6b7Ha4IU7lGybC/5JecOqkRrcZD2iVVWRDrign/BF0iQhYTpZjWK
dCiiZKwDqUvqqRp9Us6dd+kczjC6ohAnYon2aCj6JJF7goOZIF08uN2cjrwtu6XoRKVae6Q9MsIw
BMuijX3fsokgZ4+P6wGPtN37IzuNxhQ00mMlDJWtIpFrNx8ib6lLt/D7eqUeBecpxGWBL4+nii1f
zc7dISJ8PeK3pOrutFpoUzRLpIXKmWQXfgB2sVwZ5aW840+y18mLKPQ0W87tC+PvrOhtaDR902Ua
flne8kXUdPWp8/M0MQzOYsk8TN7lmI9DI9qj84KZV3NBUGJs+evOQR3ffQuBVfx1C13glgAX1LBH
6+26hh7gnL+lN/54I2XexESiTbnYg1vHuZVgvx9Ehh+G3tTrsxQ+3zM5KfouWIlji/YUGE6NO+Vl
4EMihK9ddt16tDUQTuuq8LNnzU7Rl01S9wQmzsGBWxEsgAZvReUe5fczqDPESiRfP/yxVHi9YzvD
/vgIJgK2Fjx/VXG96FKJx9gdQLfLUDDEzlHggCXiCEy2JON1KZFIuSmPAiSpo/bfu6Gy36IWTSGY
V66Mgq+/jRBo1GljpmG+ZlaHdCHcL7bWTvp3B4sOpgv85bN5ArRqQ9NAJdmtnlGEn1A7lP20/4Vj
YAdTg7MHkIGEksDKhLKlrcUFJAMhFrOT5TMWdfcDL/TaovqL1g3Q0CeSA+H7rYDZws7kZgbJfawZ
W2Bvbnh4gaKXSP8a10esqNcjVGDJL123FMDEGKd4Ecm1tGRwqXrYopcjtCUa1MsCADamhjLfOUDI
0zE7l1vcwKYR88uIJKECTOu2VAXZvUVLjb4CVju0iMCp/VdXP2b/rVF8VmtJIf9px65TWNv37NaJ
ZLAKqlc6PHSepv2CFGUjWUiEVMSnQ928CFcLQjqcub4JkhaEiX1DRQlCtYsupHslmEkc1WvgbWmC
4SX0ZF6laFta/6IoCLIVRWP7v0LXSCPT66tIu2jCyjVgcfdnPG9FUXSzWK+ffVH9Pd/3QLEyVkfa
MvAgnMnBJ6xEOL7LNGVIwLxMdLCqfwI2IECs0WlZEzQdXnIeeTysVVcYkJic49Z5m5iglKu7ESAQ
F3sybUpjMqBA3cZwOMT8Rv8U8NjQC3ofg7mqHMhegHrwbx1u9qKwh68M9jF9fuLOFlCL00QVYRam
5Zr9EX4KJOU7aw2av+byD0yvgUrBnulzL/3xjzbOyhmxHPJkSLORJCWlT9PRp9vE+Nas0J8oSkPo
TmCKuCWI1KQOD5QvfbJr/gW8qzf9cdEx0Ne1KJ+dYzR7sLlKjDzBOnNb1XBGnsbKPBEvstMmEZjz
hvXxJWrQxjqZEV6xP+E/CyRb4/ws3TTu75X6Jt1VmE2khof7wWJ7VJcZ4McbCnlOqd1qNq0+13jg
TmMG5MS0LRwPyVK8NpTgSEcU2kY0Ly07flk37PdgG5/oPHCtfBq+GWCUBMKeZNNMLsRrFZyPUBwQ
D9/R/WuefYssQR019XiOxAWjrChxb3ZbiTVDlEYItICwnDi+k8J4ClxhIU88D661cE0QuvBF2pAK
4BY6Q5vRi9ErxpC4iTFngFqB8A8reUwb/Q84J60SCJW6h/7o+4weYcnsDP2Eke2tfUez3tOKNalY
EIXyIJmdmEFNTH8cgTekcBtreeAAGWiF1qyXjLo2V+PLvUJoZ7LOSS8GW1pCL6SH3xutR9eX9PLr
hwGZi3H2dWwoTSTy8J5UiXLvM1K/KTWZ+OiII16x1sKBS5iBGsKdQH9W1yYgnKTBXfxuX44A7O+c
SlBIKZu0alkru9d8FNrQQ0s8eTYaDO/fPUMjipkk8OlB51m97L7vhQookr6PMyjUuOeSZ4umYy92
iB1MMXf6gKaC4I6cHmClJ8hEyMBW6wwVXqiCRZD4WZtWWFNXifVLzA4/1nHcDFW6zK44NeLewxHo
K7mIIcWthg2b/kW4zLMt9MoRaWwtpC3L5jGAfzV/s0SMQ67zb+rLAWOhsY2M+ehtiScBKCVa5HWj
6YH853mvh0ivaPVJ73z/XpHIncShF1WAloIgCeW95kcBVtUK1lvye3F5ACxWMLFSAsF2X29DIcA0
U4qL8be0el9yPAKQTgVhYu8C3lyCyg2nCVfx7n5yq9kTNWBUGeaNlVpq9HsLvrxyOKaUupees3gm
siuNNx5B08Uw/mrFCWoBJsLb4ISgZSWndxrTPE5vuCAiT8NWqvqg1ImCm8uV1MavU1f79tT6XRy9
IVuuTGsrBysAeuyTapNPiT8goko3d+4x+iRLv4wVMN+tMGTu41BFEmlNLnpUO6dVZ0eLA0I/iu1N
Hs1SqfodLhC0HFAJqoOW/V/ifcgFCmXST4293yWGvfcAPimy2PLN2cM2JKKLB2Ult1wldzFaCLq6
QBxxpRQUDseE077EYZ7Wl45IBbl+CwIdcBvKkbg+SZMo8heuyImcsW9cs40wD3UcuqquK7HaxLE1
xp9uOkzkc1qqLAdIewnDLgNY561b+grduw3wxTpGPvZExlrMKNvgEkWn98ucMXiVOC42lTsDWmyH
IKpQTzFKR6N8lnE4mnaICxxU2BduKjKzZqsxZ/8UWjwLIlvNDcUVtpn99cZ2ytrtaQ3kYbbJVEDE
vtRCC95SV3YRvX2F1wj0XLG69W4AWbtT1bQD2/dpc45Y7l+uQLDzyUXAq7Tpq8g7OVr6lcfAvfxy
4F2desqpn95Q2IXba53ir3NaYUiBFnrUkI9A4EaShkOEnjl3BVMD/uMsbBkIloxzrIqqtRRRaG9g
+UGLQocQ/oL4QJT+ipGciG62e3QgVIFMRiaAIkiHfNYaGYjnc/oIVrhYvQfqrIpFdJWLdcPDozpU
dugDpMf7gFv2VgIuy9w7f13gluwYElaSVlchxfTQFpYTMK5Wk4Ovd7osPD5B6AmqrxdSiVAJolYK
eUWw3x5VCI5RM75cXGKlXX3jG1S49Kn+tv8pcD4cpIbs4DfL0T8aWSldb2xS3fQtRf1zspe3Mi5U
fpPSvjVyNWyYmRqdnSJaUOlRCv5XqeGDMyRgmWAsqycMEQ9NSJWy4zNvNOHUuxSX8lFJ+PqAfJkd
/FUZftOQleDnZ6qXgIWYXArc1s7HjAyhZtwdd5+vpHHWETPYNocrLy+PqTj6D5Fv+8ZVCT0ANclu
AnyuKHA5uZTt0YcnjSZM8L0Jvlkg8ybumsFBz8AauMPJNi5EmFHciwTrHiPKlp577cRDTnp2RldT
YKbRYQSxzVFdaeJ94NKVnMIlss54EBSskjBQKXmOtvFP5tEcnk5x3UpKU5rEkS6y5rVqGKfg8ZR/
ob+WFAxcQao9pzIFMMjQi+Apt4HP1pijdcYUuqjpSv4O2yn+DJJEy4wukgKK0RdAqSR21SUuBAzg
66/jVn74NJmD5zCU5XxfuTL/pYjSzH+VvRr/KTaYuMeG8PzzOhcQu/EW4/rWfvmO3mjKvGYsWvQt
Ix1LTuuEt3NzXhzGLZt7JH8zN+np9PGNHjP44l4sn3S2Na90veZo/HiCjb2sP3QqGP3ycnYM/sg3
E3lBH2djNGK0FrI4dIrrX/1GEPxAWkZck6aDI2xJYVdHSSDFBlqWh32qqO1cDRm+fFqJ16OvT5iN
KcM6OOHdcXOexYZXHozHE4iJYTx0K2vzwogAWZP6Bj3WQwUhIq9yZYkV4RK6VpkwaIqMk3k88fZn
2Edu0KE1wxg7oiK6l9LSbtdB3hbbYdLyUMMQIic7KuVycLjqTwI2Uu6V9i2/gQH7+Y3JZOdiZ4Gw
1MPXf5+jQM+XmPx2GV/I9ZUEeQFkLhBnXl4oh1+nf5XFTDX625FzJBp03N0WfWUcbTU1M+MUdaWl
oX+apghOY1FG1+dj8f7BFtcET75m9l5wXy4aFVQJ2EVKfVK862hi4O0jhjBVmlHnmpLJZ6M6svRR
t+lT5LC1r4LpVyPynky2UENi3bLZGk4m/y8jBgcriDXdwJKBpgE9cSiTbCsvaaKZ1tKinjybIe/+
nlKGdx06jfq9cjg8wja0VriQAy1Gj1PG51yrhdDJ6AeQGpn35sil72YmZisOlgJ5qfvCnZXkAXaz
T0R+59dPXYakJCvJEY+XfntPqkCJBgj0d/IaPPl8EkVv/xWYtEsXn/7lohBMWewOZW+rEhIXfFu4
n6HUGBugxOT7yDGQ/sCTY9jxV9DdT5WvMl7WrZ2cNxN/nwKTPbQE76+Fkne4YN5IK/B9ACmiEB3a
hERNPGfR0/4Woob8sKskIr5r2uunaEVM21K9I+lrQArWmxjQqLZ8nHFmiVRyy5mCbMHalRdnGU5v
RY3v69srSThWd5Fl4J1qmNCD7Q19T/yHvYjbLbDwPPTSh1go5boaeAqW08GTY3mZGLMPG7nFdOCR
Qk9gwAvhoSfsDEcyvyR2PeJqx7GuPrHXbS14ZtrCNI9PMIzdIhX9v7OB5XMHWcl/q1VN/MSZtDlB
cKTv/Wb0b6h0FL/1+E7t7V1D9vnqFLc6BkCczu/+QFL7wHf6VZ5lV7Bbiy/bbGMh2BqT6Mjrtv6F
zjsSsmaHeYzsbMyW31pKbkn4SY7dUy9+2rj1B3UL4ZOgY5YqhwXkj9n+Lb+zkXl0IU5PD6pkWUjE
VMeN89F5SNfoGV97VBRYD748Q/r2ZUIFpimIRYwkAvs93mKPx2p8WznNj1NCu2V1c6iOjDBUEr2b
Opk+azh5N/nRHZNNk5aGYrQLfGVMnwKOlPzRYJ31FzhkbEjxSI1P+UQzrgLvaYTLTOhsXgBURcEL
KWBiH53/2fxiykpC1fHObrr6IK/ZRc5971DI+62sDBu47IwVvHtmtPsE6UoU463+wGyps/YtDQ/n
Zhr42P3X7BIep4rSyLYM13D4oqU5AyMQWSoJeQzYNcdghl/BK2rhRCqiU9O6pdzRICxrWcd1TnfI
l5ImqYoIoxVgyKFTkfZGdJzsttZalAeWnMc+vmcoffg3Q3iPQf7Ol2W8dSjbX3OXr1WjnJVHHBxv
2qh+U5xMY4qR2r5ymwACYtqk7sa8IJEBHx62s6BJJY0HRivFZ5va3tD0dT1xCRkuvRDBPww70kta
2TiOvePT6zbJtyaFPlriM3IU7Pw6hYksKHYzZF+yr79a4spfXHAjdqvDNrJDMx+ZkJgwS/0QEr5S
HaQPHWqb8iBO2eCv1drFKwC8rWRAbNftkU34LkJnO+IPfXqc8kdxiDIADEC5uMsMYtbbLMENoAba
00qg1+r6/rEXQd0+2vE/od7ooz4IVvI/8/t7N8Svt7FGa7RvaXCt337ClORgSDE9qIV5HEtQxIwO
SLos1XAcAWsn6UBZRs+/BESX005pfDTOM2w2KV4Apbw4mtSyGh8Mz8OoUhlVTLhjbWslEG8MMkdP
eplgJCsmz39u+h2RMpl3M0jTXBCT+ESLidk3bGt8jwuD+9XjLd0jNs39E+5zMQWqxYTc84B7Jax7
yLpj0t80yLRx3PIK/Qse68sjC5r2+PHjNRxlJHyiliKjXNwbjUZ6biLQPOXjIWdEc+HGyDgNChKw
7cyPTNfSujPMmEbEKzjLXtr2VxH6NOEMwSL9XRjIM8rCFtvyMbCeNbdlILxW1HDzo+u/wQm+N4v8
TNZfROdbwbIH9pZAIZObzhBFhHpWJGYIk5l/yB60JpKJSNe3Ub45Qb0uyeNi3Bj8eQ0FHFq8TF4m
DdAsJFaIldUW/U2aih+9uGOrlMkbNqs5egIoW3/cGWTrGI27tJkvaFzm2pxSqCR/WXwMl6hHZWAi
Siq8aLr+cgnOQ5OrnZcBj1Hy9GFzCh20htzaai3Njeuj6+lhEulHbOxGdseRZ/qb6amhqYmPgne9
7NZftmcX8zPUI/pY3UuJ32kXBzPAhsuQ2KhK+XJBhRUJQlyUuAFcJ04hr/T0dPz6a4GP7qyVUWy4
p5elUjedeK2qW+qFjDU/ZtUdUfJoD1Rj49tr1u8obNvfwMXKtxTfuKaoOr63UQI1XdV/NULVpTG/
OxNhYjqx0XA+mXspE4YP5oS3Udo82NL0P2xqeXEiq+QMJHyw7SphjocFd70/DZQEiyIcZWfg4jd/
KXZSUBR0sTf2HrQKe+Z+FVHaJ9Wg2iQoSUuBhj7MyepTrat1E3mkoAqRs6daxnz6wAX0gQHFQ5Ms
Uip+sbfHPL98HcPb7qv4VoC7byAc5vr3G3LQ0x3vPewXCPBRBIk+Fxl7U9ULg+x7ijsUFi6JWPnA
FnN9ikIUS1K8qbaWzi9xZ6K83JFL5hO+3WLW40HWIUvcoJx108cZMd3xXCXUEau96KXUrfuQlpEt
lkiA1/In2NNc7Z9fvukH3KTd8jRoFO4f8QWqiqfb3USp2fDPgJLXFIFhDpiwBo6OLrGvztJuYPaV
A6S3vCI0+rI6XMcssWSsCl9E1PzsDQBg9GtK28hFPfjIQYQcaYxc0xavMcbnfZWPrPrmPLan03ZS
YysXbiAkV3B5yb220s2SRmFjjck+EAXJmTIiMeQ8NY0VEp9fk9IP/7rWsXvPc/NQgE+OtVNM64y4
bOMhXbUrQflalky9v9o3caXAuW3mIPABLR+JcRfwTccMAzIvLC754krmrfChSnn1heuYw0tEJbzG
iXAzRjzwCBNanvAsdZyvDhbrMT88z6Uly0mnIhJHZmW5T384HR+OKeSd+g8YexLtnlJ9FG1RRaQy
W/VN3GymgZLw1T1tyHcywmrlTf+Mb4OWQ5SHlSXJu76F9Rj22soz21m3MH2+hLVmFItY8nz741/k
PSlY+m3pDvO/yjMSeXyN/cbES965q3KxWkk47gE6dgYiCJ2fIW5L2HvIAsZHMfKUUuGQSgmqcJTi
3u8jPGwG5t0g56SyHBOPTKMZ9KSaZrR4VkJeZySJfxvoD9fLKWn/88NstefWhS3RbM6QMw80pqq3
rpH0GGQ2AmKqmNlU3Wk8tp3SBQpcmZqdZ5Z+6oaGzqi5W6GSHeoe5IcZ3u6WDSaB/VkAhY16fwOL
eOHbwR/uB1FPkYQIJExodWNVWkOu78+PTs0mbwHUGM+emn0NCYozcD/Q4pcvTsvQUe3ZABn50mO+
H59Lk40o6uak9SQthIN/NGtnJ4ZdcWTVPI9uiSXUnEqqjy5/8//jtCx+Te/29DFzuZvm+7W9N6L7
z5WUaUfyguz/c04rFlKrlFRJfeLGRqzK9ZmIYOoWua+mnpHR/BS3eHnCY9ZHW5kl16Cs0hPd5Ufj
Q/SmBDSgAik896RvfzMgLtePLp/MymFQS2DDV8hDvS6SQe3CyK+w1IdXX8Z2pZOj8oMq3b3TQuhx
3b+8oqN9NG1ZKwZGQ+51+rwBVHDbbRYmeoSvvturRdDUQt3UbeG2Wb2t7G/FBkrb9Hx/g+edHZ7A
5A2guzKJt1moataSm+GeumVVTp9cjqHAoIWTAej0aWENpePJ91p7zi0AAiRoPqaRg1U/+lAJavlx
kG1DaV0nwLXJ3Dfwl6B+85q45LwRk3SsaNhfyL8L+ozVFmXfqapQwS+H+j5DvH8UQF6ouIts2S2r
bfykMwM1Ndtr0/Gg0uQ9FZGEF+JneKpqKQFoO2JxcdWhHsLnf449tnSwNpvsGZl5PtfPBg+/dDGB
TBIQRHkaEnzraWXoEDaJ9nh31rpH6B4Ydu5oVYGSNS0LUdMCimYGuDmlUv0JznSvBgTKLTaBtd/3
ikV4tyTu6kKWjRH2H4o+eoIvu1LIyZZA2NJJpxKb+klzsEt1Bw43FmqBpjJP+yifgeNx+gMalVGd
I2P/Fiv8WD/8YVe0E8ezWhIpEokDXiHZswtZx4utJ8g4KI/Bu2Qq9JF709vZE1RbC7hZUBsqqtKl
BWDK5PzDjjwbeSvkyicW5cLkI/6n26vGKaYi5PEidoLBUW8NZP9cqjH2rp8Y3t/i6QlPN2M6hlS1
XdrJ2lZTdYlRMORwOorIn8xSu+ciX2tOIeXdsRAuKNN3Hyos5+orviICig9LU2fLYT2h6NqDOLVT
BH5RKQavFqhtZ/5x2eozf4SaMNuvfgfRZdCdNXYbXuW5qQ+3te4vbJkuQ1pDqE53UGspgMRuUPHH
QeIBdaNy0DbjakPinxB28BGcxpQ7sVoe2tqmxO5fxptrFlvT13uVFVdmCV/iro5QbO68xxNOMC2Y
cP1WkbxZRTvHn/OJ0vGAFRXLjUWoBGCVqCoRzHXERKJZqpfUF32W5fTTYXSERwAhyNkbtdpXcvQy
ZmGXE2uFoanSXJTo7j/ZEQtoEXd7Bx/fT/JyJYwV6S6ohquSBqVQEaS2y/SfBMV9buEjCI6u0jvl
tMpGmkgEigV+q67coSHuTzE5KoevBMwwwcP075aOg8LL6ppwjvLTby82L3qfRk5k4xFoz0+Ctih+
6T9WcmMcXqpfrgTKSujeEUH7PP1j4/RvmTZVVIw/nKxq6lkvWhpP8w5WA1iOWlFFEK9V6z0TXyMQ
YUWL9RPkXRt2a3pu/Cieg5f5cU/gD7mHZCZnY/vhImvrYFk3Z9Al6HiGSK/50pJNT/1YfJJAexke
O48vg+V3cxDXR1FvE45rsMZlVBvygOU8/q+4a97wrXu5qvejwHbKudH+mlLyFToa/1t61SykjgiL
KF1H6VjeKTfySON1v099+IOAPd2jc4DsEcbJ2OYAFdlLhIx+xoTJAkFJlXDPN+yxYIhzMG6zsf5Z
GxHYvbmSsbXWdWKzF9huZLDAd8WLHgaFQqTUY0VQVvRb0ml+GG/UJPhHEUJhzU/5XXveHhrPCcQK
x4cetM87Yzbjvb9NawjOjJ1nk/F2vECvpj+HqMstkFlHmSmi5SL+AgqBpjjWr79BTBKWoBNGX1m8
1n4ZtPq0fleFgVTO5pCmHg6LeyxlXri46Qz53c0zUu9s2L65mJDRu0esE0v2rKrZ+zLJZcRDzyMC
g3/jdsr9CKh0wya9MAyGllAp/vnhqS4GizLk5kMnoyFM8q1cjE90FJ2q9QI1hvsGBuFYhbuD9aJa
X7VdTbwYOPFpYJdgZlz7c+ngQdMoUCsdfIuzqPyCChexPc11jNagnT5x7SVgUnfKvgC/XkHjqU6B
U4OYZGh751yrPxjnmVoCvhCj6lmrXu2bFqtw+J9Nt66FP0gDA3LbFMmmbF1JwhDXqj3jk+PPXtv6
q/3eNwQcM6orK357nhtkai0CQ8TdZ69s8/5gda+6LDeyTfsuS1PesrmkxWWpu9EprjV8amUNq7ng
dRl4vncuwfocTojxowrDpluHCkMJI1FYADqwqTKMt6HYaxKS6JPtGe4YDRsCy+Brvu5x3RLuOfoM
uOtoj6P1O3BSOrq9hB6Q0qNlUlEqUghet4u68Ih//VHqCJjrDWyTCuwdjr8nnStV8mMsN+RshFrd
56i7r6SgY5zOAnWjHXztfYbKfN8Yqo3XgOIIbSBKaMtp2PtIwyANKKIDTfzc5DDgQKKXQLsVSH7q
FETumxFIU2/DkcJve4MMCgFxVKDiSEnb4w1u94n5bZkmUO2TCU7XeoaItIGhJa9W6bkfpxXBqRy8
BxOiOkEgz4o03ck+ZQSQ7VgogL0pSr4sF8Y+v344KVFvspHhXi+9YRUKwX7fdYX+wldcv/l8puPR
VE73nsLqJoWOdgEDNlVaBCQZkYcNMCf4xMi92R9SsN2rwqbxd/NVdvu5h8WLksJO3aKXytIvWUar
8WetDOLYWD0Og0oxjWm/xqcluNlkmtFf1XjAxzLUELHUjadG/sIOd+YkOmaTMSIu6L6Za0D/M9jz
Sz6SBRLhJ0DKHVfjHafIQLp26d7hUp5ZQZn3Wo4w3K7r0XTJ3ZbSSbb79EozQ4DnkqARPDza9d5v
3VBCGPl0xd3yTPVfA6mZAqtdcdrJZ0up2XUu0yv6h6q9RdGQUnkxy/09QtHlQyEcufvb034ffK5x
7zcj9hUrGo9HyaXyHMgWsxlq8TqxrBgm76nZIss1u+esViafTcsco8vpdfsjlqvQRCpmAyWUrkI6
qbtJoZUV3Xsjayp8AcPm0ANlb4FuM63Tzji62ZFWV10UBmBiwLNzeeG+jN++80JXq3denAM1nR14
sY0clby7psqWEees0+D/L1ncmB9UG5vNzS/pwHOXiNdYm6lo+jB25Y8KxLgS8TIc0hCtlosKj0IA
EFIh5zD6VzuL3VwPLyXyHmGicyLY3ckPUFps0gBYdMYFXknDY3tx1zUxKhtA28rSUQ3o7Ibwlc6q
Jeq7DREwDkvo3f6OQHVAjIZrPXoruBduI8+Vck07I40ug+XzeqyyzZzE9Z4u8JikrI3/rzJznObW
grukL+powDIYkJtRh9+lkQCYCjK1rhpMcltLuBqkMTlmvSC3bXnV1NK2ZPFxe42BNa5YSMSj+Hbn
CDcFzis103MGD/awM4C08DGVmwxYn2NhOMwRXBSoAHuCIw1nmWoNIJPqCodwQ23ATAZ27tM+0sKT
sM5x1q/QYEhRWnNl6YGdv0OaBbG1/RRjkewHK1xsWJ3baGAKo5Z/AAF3ckkMSKifDCK2Mzl9UqRu
WYWjjSwON/DOaETZ6hvgCh+2Umqk2YChs9Uqc6B/SXpEY26CIZrhkqxEpFDcv294kyGq3+Xg9zor
Ex37hMEuKDjQcOr8tWUMCZcPL5sAz355VqoMMRv58K1FiAn86VrCAU3KyFYglrPGUcAG16vmbPqb
ZaDIV2gji3QwIFVU+IkLCNMV1jN98ZbejyjKf4MaDd4hkP5bTP+IlaWYCYJk6kTBwtaofQMx/vzh
dQ4llQEiG75a6xTGC/sN8yMFZBa1QyYhYze+IIsNDqxOcw4PGQdevV9uUZ0yEJ4FyrY6cDuLKzBw
XNspLk/2tYwXqkUWAURc+58HJtVr/ISlzkVM3RuvnnoV6xsSU3t3w8Iokt8pWnzXcuezaIL3aZH+
Ap1R9eJ9e0qxPc7OS8sgpLEebHShnCaoRNL9VLiiiBE7XUvGOnMcmssD1Vy1u+QQefoRG74kz8QZ
WTq7N3n6N0FqczMdf/Oqh6tGagDp0w6M1Nm5pJf7e1y8GjW/IhpVmWTMeY5JuBj1v7w36mbOkvef
eIFolJV0oe4oemdpftD0enRPvS1KimSmo+1N3MDDa20SUtB9aSW/gYmvL/casGf6oVly6+7emM7/
GcNoGD8LOrg06Bao/dLNJe8lkOqaw8kLMdP7C2jOIcPT3rx1wxY+HVdKWZDwpUZaA7LiiMJScHYK
DrDHB32CaOJPa2ar/NK0xgEp7shqvl+e9DR9DTJEYSXKlaI25GnfygX/NCyB1Fow8fKm2CcqQ/FA
GKwTr5L84tEPCICU1kZCLtJ1tCtNPX/YCvvSwf0NR13wo4ay4Xa/WkmJiNdSprqHv+QcpAdOeZDN
OFcOPZeAn3gAuq57SsxSXGXLFVhsBRhblaycZ8cCCH2aQSy58DZX8tIDfx4dUU3borYEVdg3UQH6
2V9oIFI8ag26vRqpnseGCwyiFa9yDdCKb31R6hnSKEYNhgrXY5yJKnDh61/cV0bIeT4xQlJRc8/H
aABypNV6eW8yyrt28QK8UoN2aqNK9Ylf3I+tk8MyfvHdIbdejoLS7O71pFwcg/SpADycIOWiBVh1
sIDy+l9vwwqsY9LWbuHbAjvoZnO8+DAzYnK7+aTrggY5DddNVyqWQJKmQOHOep80wcuqKaHOHkzz
s1gzgHv4NnL9jUR8mIKV9L5KoG75b9gYxi0jmB5IEsnAz6vHixVGDLL9T2rs3j11HfmscL34d7hJ
cBZTASlrHlrY3rJtJWFziglQv9AUoYZKqLDZLSnsRZn4JVFof/OyoNkwZ033b9jx0T9qVxdC/q2m
EPdUu9MH9aYVp8QQD/nyjO68G1LN8oFy3Cl115kELJcdVoBFZ1gn34TDe49jpxx9OxD52YktKaRI
enQpRZB0cbVSumgUoVFmZ1tV0VlTEpS5qvwmvlf+si36HXlayH4cEIKXeBKQtJIxGZWFyavjbTvM
iw8FxGrVozobCqLGO0q176QfYwcGpNs/VbpcJehT+xN4YXGCHHhBlKUhB9XANwYN+VeM/JANdxaE
t7PS8w1br0MIj/6SK4onkydMb4YFX0elmDqIDdJxgSDe9Svl5u83GOEK22nvATRLTLI876WyLwyL
xoaKPPqDFH8Nzf2pzP1YkqV18Klipz0cnJijbEIOkUR3a/1PS0o7HwKmGoZYFjV0sefyrGjZcuCY
wqdNbNuyVaL+crHuaQN4keUzAATaeYwrXdfyzR4rd6eKwxE6WiGPV7ypzWRJ69vcnC7/JHfbkAIA
epvLg7dx+OuwMeIW+SEznoeItkrH4UVHn9w9spCeI4HHDAxg0l9iJOm25J2ZNqLYPte6v1Z/3IY5
HlCIWcH2yGm6qN15wXGMpZfr0Qf7P/zX0LOsAMJuFF4JWxbFMNKAqrmN/DlL61snoDyyCp0hMzzy
+/oqKw+VpSJMLkv6V4ZR0KZfb2ruyf/uTkB6Ghk7yeE9c/uiHlwJhaeGmJN2eZvC7uFwHJvj7dMh
v4wDvaOvcYIkss7Wsg6ad56pic2hbssAm/pXJE2oS6VKDyqFjbMxXPgRDiKIPFh0V5P8CIOL82mo
cJ2VZCDrvKnoAtgtfYVeG/3J+qSe3Mx6w+PvN06W3mSwpjTLan8h5Jo7Tgkx8nnMgb3t8wwUWnID
W6r81vtONp3C8JWW3eeUD+Pj91qxvUwTw2JMcyKaKVMxeaKRh3EFOKXUKeXlyY4lkGDrTvDxg5f6
XNBjoVNVHGnh/nBKF56Iiy2hvZIkLiNzm757pdVfJigyen5AYdAnqIfGfl6cmyfrjXcFvVBmMrbr
TVb1rSn0z4J0DcNZbEFMka34uwo0RCtuqszNX7eFjgx6b0EBHPieYyMulTclO76YxGxoQD9bbr/D
LBlr1bDT81lZnO5bzz4S3OeATWsXb6/3jbunVFN02KDKXreV6i9tF76a8Ax3TgCIRcFCMaMZt7Pk
/EZlinpL2nscKHVZPiYqB681tRopS7GFjZ8tKzwIvBNeeTaiUXp9ALIcJNvyBEWt20ybJzLJtB9z
m+qGgdtXCtqV9LqFPFvziQhG00LWNdCbluIXgrtzP69e6SVMxATjkuSeooAdU0T119Ko6IJ79yPC
mE2Sp3LRv9GV8Fl6T+WgYxCdeMP/g+sYOYaaKcqvdDWb/UQtkfXSHJTJ+K2JYooz0e4pfvDDTM8M
1GQvap1EokaIFe0oeuh7OetoYAtxo1qcg6EBhES78f5NWsKRYTzU8W/uZ6hqUUSPnlujysrDXYZ3
Lkc0K65lBBfLcPGerg/ioZ+PyuOycdVqWs3a8xURKO4ooz8H8ODNGm7homxCZoWjZWJ6Acq6BIop
jrB/hklXUrrFHbvpwL+bxMu91Fs+C049ScB64AZp6hYFEHcG2268yVnyWXfBw50Xf1h6gd3LLVGK
MWNMDM2YWrt9SvvBUtn9NHIvk5bFtkw9m/QO4pybLunSAdZ0OlVwyK0TQGH+OE6HgjvvwK74QWUx
On3aZTUn+jCbBJJ0ejpJZVWHcQtH/jPgvPasFyBMoJMJutOxFvgyIqUFx3V9TUXNucLpfeMNdwHo
PYsYgpg6+kAoVLnPin4Gp/GD4QspN1Ol8XWtNUZEuODYWWw9QrCUZQ0HriFK4WZydnipKbNodYkj
zeduvQ9WTXmwLN5jlPmstCat8+75oumQTkUNjaMYuaBkd+VBJMeP7hg2xToR1tlnhave5GwSjDU6
8tbeXpw/Pwt7yiDlusK4+RLul0rAWeCvgt7YtySy/slBy2LDzS7KYqtJ4F4R/Uc5AF9DBbcZdWz+
OyChgR9Gr2tom6gtBrLrrbKGNjrjrU6zcRJNWeLjNggdn5+HGi30ZdiJLXwvaFvMRRWGLd76lzPG
FWkzmPDdXdN8hHKmTFjcH0pmVVk24BmaU+nPKTC3Y4+Bpb8cg1gmexE0ena0Z3oQewEKE5Jzc2CS
dBrG8GeukcikXbjoVmzUurSgzSAFWLyHd4PaydTRsa5KdguJY3TfUQOFK7DXdWImBDS2S0K40bvj
CUW1tNMTVifTtso/4bsonedDyxBLsPCYcm2pX5qpRBdNrYx8wEUB2GzYirKTRUpEhDgy5cfXpg1B
FSJSh2TpT4CCrXU6Lk/lErrCfIOkQQyo78+zIF+/8hNW6skl8ls3KVQgIMk5y+DHfhoDECrprT+V
yvoZ3UfSbKD7ujNVcDCFuzMhEbKxlWjOorQY9XnHmbnuCe71G4K1mm/5+Ht3pOVGyVZe2Eterf4G
G7HbgxMki91s+Q/nkezQLPqb7jZV6vJN2/UaeZWFWbhyc4MjgbCDt/oD3JO3OcQSKjosL/rbpId+
0kjSMlO2smgNdeMoFBpHSFPk5sn7KuqXmbLMvm8ZfYWVZ9awRXNRcrAYpAabz2AYsGtcCiAP08Be
9KsIse1lpnviGIMHer7W+IPkotvuT/Ra1jCevJWQw+oarhzD98n20+TNvQbYCqTl2wgy1zAwdjwq
2vPybVsB8Tl15cXtRnXFY/KyKPFwNxpHQn+kRLV1jqOxrlpkahHRzoCz61aJhG1Orpz/fcQq2gfS
CMLuqzDm4WE2uhu2u34xESu50FHVsYoGmwwYX5OLDuYafsAhWE1wQW3hQdofUUevSGsTaULuGosR
micdQXY4OP+qV3ZbP36+rvkp0/VIAV/uzpuFQeT2Tp1HkHJUNMPmpyYsKjkwWMYUb//mwVa1oPFH
pZDloIfeqKU3n3/5YKcVbQk0mavXuVDszHQhWt3XVjHdcy3jqbqWrYNP6g33GIv1bnFqBLQsOWCO
cSs5qPptiZx8WNG5Mf0RCsuKyZJVJlDtjXmpeWP6H/98bu8LeDhKZZsxW0AbWgouzOFzM4uiBKNO
LFyQq8tP86+xA16frGyb6bvllVdjUoPWIYh9cQNKWzHcRHz4dK7fqvuDDxU74iDXRnAPXFRIp8BF
MWSzSuDuZgUn/CfYPMcKYu8DRL9eyYdOqos+UAzLlvsT1PXgjqjR0DsZGUbp2h/n5b2TfV171ML1
qy1bGdUfl4nR9uOsrxKaU0JZwywe+am8akwFxDa6tAcPWldlKHFTEblf8uiBNJEbePGtnIFUaLlO
RyzK8wPuKckAWXkbA9h1gabMxYqKD3PsDj9bDzDGNH+RZItXPKAOq9MYUyovGxMBJA6BtTuAMYD4
Q0MKETzFkMIW41XOatfSGobIMz+HeRWOKyqU758vM+PdZ9CEkK2PJFkccMXRhS+4RLq+0nTPZ8nl
Asa9Np2psPN8UYPYoBAcFbkNMWPNoVd9wRErc3J5oWT9Ja1npODqPvFKpelgwk1U302I2EwJ15xT
zEopNhLBP16Jafvs2UhB3FBvwYOgC+h19Z3b6P2QuMeQ8A1o6HTtphcCj5zBjBWO6l6Col9PU6mF
EFmFMOLpG3TVkjeJODK6syEma/kfbsCDhwTLCmxJdTMt8MMTItiWEP6TsL1NnWvmHlZX/WRwqkNA
biyw6ChM6MvE2ycWiriltpbUHn+UtDSBzXTYPcyIXSgV+Tga3/265HAQaBkcrt70v8jSPCccbnEK
WMMWRsvxIA5h+la6DRVyAZLSJIDYJ+KWozjYSI1lro6AyY17QommshtQxirzNtTAj43tpNtEdQx7
iKeD0un5by5v74N/x18wTYKHnfHjURsIeMC8eTRpcEpM/Ptk/vp7fX9xdbhcDRS76FQtqSgokx4C
K7CBEakg8qqO9wktfvBLSDyhrucGFohkIcX/qPT5L4KHl/FLWK6NIS69gMEeVWOVU01PRoce7pQb
/Bob8kvy5PiYvmATc+u21RNn+HkYjMjSajPh9sEOiNcigMsrSQWEqn7Ur2evvMz3OFL+w18vHToc
RQHWkdVU5fYtMZKSoVDvlA/vTsC9Cj8pImDc6aSJPZL3OT8WSzE8bGN2ZpfuD8gLNwBoJo0mM8e5
yVZPDivxE/EMsel5GSYlrKTl6EJ2SEuD+liZbAJ3JslGwHP36aUEBY7jeGwqrNGSDsm5kHktnLwd
kht8J4e2obS+gh6b5TJPB0cr+evdsIHdJbBzvqTwMc9nANT5zuMGkE3cRxQApnz8sJe8x/Kx7fpJ
xJYYtBvAsK85aeL1cc8z96ywunm8s7VAXUl11+XregulvlcxVREoeGnGIophQMmb2DXgNSAUUbsS
xi133NNeScEEi3UWf7bS1hpr9bvLvY+5utOPVj8d+y6TomXgfS5kYt3HkwwAZ4uXRxwyuzzdnpj6
JHgVIzPrBHEwGuS2pw2aTTMqnrUfe2RiFvLXeu3n5LMRtdz/BsoUgkvSefdF0aSQBYqBATfFzVcl
MW6sJuSxI7I79z77bPJCBmwei4xxI5hzdzEIQOk7Motzs+kj4LeyxrlbbodBm+WIkzGJ/H35hEUu
gXIN/8JeolBpjnc/tV2jeonq5YYjQp9QpO8X1/L4SR2Yrp7RAaHzGdhRCHCG198whc2tskxBRBMA
A1I04IAvAdMBuvMnxbl9Rm9FAsfyo5aKxxJcirJT8nwpBS3dM/7/VdG+4uzzv+Ng+xxFziHjiDtN
gsQMNcc8+dtMNZ3961dEv7aircXenU+cfaxSHOKTsboqxlNzK0p+lMmGvR68T6OvVBIXP1T+Yxhc
bHr8LMES9HEqjNMA1M8pLIP0LK/JDcz2XaJXy0uRHGO2XZisLR8v/iJcnTrb5C2LYmbjryg9tNOH
s3kxdUgZmAuCngAUxm+6Erho7dbEzDCvM8Wf2+OL5ssl4bure+7v+QlelOl0x//BHaVXOFjylqr7
kndOcAvIBcwKHoMFUSPhniwwzLPCe9DcdWu27sTsgSpSczrMXaMW4Q4oUhIZPZmXjdyZzC50fOG4
yQj0NVgeIlbEpfKPnx6bwDIXI3qMzWegc7RDiwuMGJLa1vdnr5u0rqgA3sVpwIY3KTUEEMIY/W8O
RcJcqDUm//XjRHkdNlNAtBGT+g9xUbRjO1IIgQPpDc8Z4bwehABWCBmPwAPBlcAJ8XB4yddH2Gnw
p7C11fpDOwKbRBa2tZuMXL6i32ScBwBrtn+gggi8DS0nGsRb/98VokKrtgIJYqlgSve8fdNalFgu
XqhuyZ1e/J9BGgwt+FLT+/9Z8j/G/bOnOBBcalLBTKZUwiodtqmncXEzw5GyXA3Gb++wWG9/Mv9P
oSrYWfEAbLGANIw1OoZqYCqXV25T89vp6xXAGhL+iB3CuiRkwqRXj5kpItDtHqTVsg0yas7BrZkR
BC2HJ3pzXNnAGwEQN/m53BUWfajB7esGiPkLpe7MkCsIqQW2Rt3qZFDEa/WsvGfhhbFHZdU/nKkm
9BmdlwLd1+F3SuXWz1XB7V55/Wbf6G6gLyPF+eodRYkf4JogCSM5ZVBdW+6Dfi7K2EONmAkwlPqq
orR4k7XLw9UHQ2m1CGccve9GfjNwC8Yy2cChfQS41Cn22wMauHBiHLLarCu+oSJUSag3Q/dmPCbE
7VtqaFSDNiglB+YHY12319LI0hErphnp79fum7e26JmkgvDCNwyMYBZrJO1W+X3+iaQavapH6iRo
ACGkdjp4/85OmYJ+rAcUI4DeMKc1Xkj5QPpcnZeFpJGFgiG9WmurEoML8GOLngQromT45/Pa7aFq
b+M6hBr/Jw+rgv4/0NyZoRxIRds28pyLFrY5mVKF7U2ALN3W9KKF2Jzf+i87xA/6StsEhGbp8hyI
lmHQkIhTiXCBoDELOc79pFASKIFfareXppQLioJfWhx0kExpYNWZelaCAJnIat+kL9jmDEC4vIsn
VWBW38dwGJglFlEvdTS63Te/jnLfe0aoblBtpitipmhe/ZARPNq+62paJlzvABas7kwmtPdosjEW
pBZagkp9pOoWs7I7IXflKNX2yKX2b6X1s19eCXU3G+notx407Ow+NmzLe1q75A3Y5lq/O1Z5Jip9
N+budMvL5IIHKNmbfBxxX7M9KQTDTQwNrrm1GsdmbQT8OYiCoQkyBVZbtg7Tgus5MY0hGHJS00rx
RS57jtDJuRO/xiYt9NjO+MQ3OMi+xMAbJwTy4U1jX23mE15wwfmH8Dnr3G8Wv51SVXzqeRuUU9aL
JYq8bqgcfCli7KdgRonUpIe9k675db01imLYO2ZViDFf4ZPuoQ5aFtqTuAJxxwDAg18ZY06PKRTW
y/lylK9Vnpf9D3tdvzeyqaWW2OIRXCOHGtUXfZLwppXRhKpZFzW+VavqNaFdEkA4l8mP7YYzxFzK
IDd+/I4VSSq6lSjfBO+YvSrrdJQSF5pmgnq4Za5s7cf9jUAqqKb9BVux19DFlcZ0SmM1kumeiJ9P
X2FEHkOQ5el9r/RR0azuLV3k4p1Vzjfi2DlUYmpG01vwU1MgQucZeCHF0IbHOPdk10cZL2MZFE7m
CM1NORKAgHErdGE0K18+EQBrsGRdNlTfY5KIKvvmn90vJQTgewgfqMpZExiVgt/5tDm4c0YhcjCU
tlWDcknWBr84QzrFv2rgM//SROibBX7KC4MSHeSm/4ivAmViPE+gjRigxL8TW8axd6IU7FZtyHyd
Gr852m3A3j6FBgNL7gSGjQy/hPcpd/fp2fKUaYY7lJ7A9QiX5CHCCGz+7qp+7HcDNuxXQETX0oBl
HGRQw5Sew84M/IONPoG2nbDviwoxLXt8O8PqXEMnapx2hgE02UpzF1s2K27I3gE9opNRwuLoGCLX
4SgFE0LzNkg2gkThQcwnNQvCWsJM+JepH/6psp7cQ67dU4ctP7frbqAomBHnK97A9HM4zHQ3YG1w
BpnSvZrg3RNNZcZ4rF+fzeNAq3lEb6Fg1xfwxl+zLv3mVbzSfbSWAA9O88Gg3wyYUOlNf4ntP3E/
6wvh+2j2cYZAHx7sl31ZagTzoM1FlFVMjJFZZYuKgjk+KV/5rQ52KazYJ21QuiezYLybKClz2Txd
NKTpn+riEeYoORo8pZVZLmi11MehMiNk4c047luSam6iFPPpW+VgXkEwGlj7/wLuzBzpOONSA1fu
+Aa7lUKnMeNAKCmxA7e/H0tUdQVIf4zCbfwqUlTBhS6DePKKj3l3cu0Bi9n+B17r8lvKN2LczYL9
wt2ssMuHGoRaNkVFkJtmym6m5x7efpHX19i2ZcczrGqSsVBWXGOx7HyCpVbIPvQJoPkb5wZtJzMM
8qOtzd9fqlwwimUCYyhC4U0OTRD8o2Ix9UpXr2pDnTuFbejJlCu+2ZGpdFSfnWVsuciG7j7XQmzw
qaxzYi+20k2xiuIk4gWXh3yZiXgEOznNbiZI4jhTRL+Zr7ySnjdDwcUFDfPMAFUu2Rgbyd/E0UA0
p/mDnOKK+BgxBxW3AbhVNcDa7Ehzf3GuaFuq4eqY3fgavwpMxf161f0gM6g0lZYA5sVZDd3BZ0pf
vZEE334RYC2NdNhDs3J7Fnt7kKTFKs49T2DxFrHpkvWr6PQYVKuOsyNJ7oDen3AD5izuNbAkkS+3
Maolm9MKlvZFjFYBv0lZcbS6RcdfLa0CR3+/I0LFt2bRFzB27DXCrZ7VuCpklfcOprX2+7hBup1B
vF3fXDj3q8NFsNETBYCW9WTMuR2x4tUjw/Z+77xDU567+XdtKR4O6ZMeTsjJN2IpLVYrbX/cXeUB
pvuN2ZtDeVgzCqzT9RA8kLr48Vii1GKz8wo2Z9hB5ttlcWhowT3lLhp8oGTSfFpAkilRwSfZiLi9
qZ6uYxl2ONr+cvMhphJXJM0hFprFB4vp6Alp+3Ismm6PCGJdS1tIpiDPsu1tKKIv1R071Nb9Ov++
g7yacbxDFTKDLO2vaflaAdUWCQoV9Lr0yUsarVGnfCKsa1DuAz2Rv0knn32jzTDOSv4i3r9UT1wA
QtgwklivXDzx2VVH9KTT5pIFdlO7M0ZqyiFyqiYAxcEd+QFokUi5QovfK7CyxOLbbKTIBQ/wXl87
ATP2shE+FXbD0eH0o4f16gseKlz1bK3aNfumGZane9zp2BQHKqlOTWc8jDkwJyItMeY1mBm6/oHx
Z7FKYI8db+B0MNPMsqjnNLK1n9wP/FLD0KSdu0EuQUCAuJzhl1OoJpkyyXEncR7Ck/1zosV6mNQC
hZzeCT6RhGAFEylIes5HeYORpya/VATffxgpnJiyL7JEPkRz9FKSOzHQxnoT9ngM1ghhcmzVZ0kT
Yr6p8rpc/GDJWPiS5bYb3TPJVZi7vNw7uHEnBqAzOgB5S3FRUtoNxFcqwje20KB2a+r5ciqO9FGK
fBxTYkQ78caEs7z7Cocrdar7UcUvFDie2PGWmkOQl9mfkAcfdI/yokzlSYBq0dAHQIti6TQG3hSP
Ogs61prUMyGxByOCk8WWKrGWiBtAnLYFYkSOd83qqda1LKfl7JDwIiNF1v661MPDn2mWHT6ijh10
Zbgcd5HEH90aoD8yag5dnItrWFstPuBHZy4TpG4bqimUIn6si6HmpbnF2GnUjpco5DGndmXwqVFt
6cP8Li2zKwaJ9zoHrnB5bmNPe0U8pDJKf9NXGoMa13fPdLHEbRnviV8A40jVbUN2ub1Yqeut90bz
Qzc7/33nTHPWNvpACqiatmBDifgn6Mq5eSu/Fw7qkJC8FERDiq8UDrB8CH/Do7mopqeN9c00vT3W
B3OubegFsYk9FniOxZFnT7s8RcjiiPz3W2GQ3UP6/Zp3eC5s5SLnNiuzi5DyK+hZvDF+vi+sWbmU
HpK9+e4OWZOOQOOpwxjYHMd/0SMs4LjqzdvRU1DwFV3TL8NFfSJmP1+yj0o+T4eMwwjCvR3WCZjr
fiftZQr4KdP+Yq3hE+TNd9RNTeHo5+DUJ+EzJZXlmpC4zDdj0KRO9jJUS9xe8og0ZpzXTA/4qL9V
cYPCKkQUQl9I9DTAHkmJRd9J59u/8vyCUlRH+Y1dZHZp0FyUMKf2tOA6RETh1DVPWfg1WHfVIttQ
TvUjT3N7M4N9UtMJLpoVGwBdX+JgT2tdaCv0nP2YzRmVJUYUZDLJ1vAXcRXdqW7/mW57aX9ZfmDJ
5zsFBdzRYplF0fEqVBqbwMnQWQOo1PsCvCU7wQuI0CITd0XtZCyf1vsy7Drndqi/Ai59+hxqgr49
FyN+cayBwcnTh34BNDv6E+D606w3CV5VueQAQa8UHO3bbl7BfvXjseSAGDfmgTLiCHecAQpln6ak
w7+oXEvESPuxQsfD6GHWARPAtEJO/tq40iTk8H3M6SCDMBH8f2nX/Rc82839M9+xhg6jtT+recW+
+KwMgkfim8UhSzpuUbGO3ZFX83YcDHIogCiIjEe3EVkmMBrYPzKh+6Ofi2g5dqnrfsGt/w69BCrB
iGWejr1j99XgHY/B08fL8PQ38l9nSB1zF9tGR1ofL5dT2uua9823+9DLynIMP4KwDq23INA+RqjQ
08JD+Z5ckUJpInSbCp4sjxqaJvKsO0WD8FriIEGikRcPjQ+jF8OEBFli07pwADoWRZCfADM1eCIW
BYYt8tchPRVEbB1MRc1LrbBWdWtudPGVbm6hBoIHknDX89iKBVoOy7qvpg68txKZn7FylCUDj2KL
qLfki3xfbgLJ6ePIJNnhdSUpCgq6QamI2B584bmXSwP9mf+qK9Pde+yWf2hZv1pedzFFtl+bCY2q
4QlBWcdLs0evSByXAcVcPoa7t0POErNhWE2I8ZXPp3wPNkiQ5iLuPc5D0A7qE2vjMkxtEWqNoAQt
V0cDYRmOvcl7NfJHen3tDxN9yOuPRcw04prZuOEBCCqEMZUvbAijp0d1dmyLRngjG5dOavyTx4JP
VcFE85hQTUlcDDiICMo2C/Y6uPIuhKcBpUfptQdocbO++7a2F3k026Lr21maZJ33dFzhwTqBKwih
n/72YUwkLhssDZkrsWr+SG+F5E5oaL59SdVj3J2lQ+c0CiFlqR7vYjlqfI/3Yt8AhvVMldSG9LqD
L2OqUHg53ITOBp1IMppIjAGoP3gD8SXIVl8zbqeKyv//UA9ot2z36zBkLrYjgDNfZYQlBY/P48NZ
DBArkmhE6cb/CAGFWnB7dsj6tVHGMPHJuZe8ljr9ydgm8FQ+Tp3Z+hovF2Vbx9Un2ductNxyQGes
8zSemVE3Kfm0pv4qD0Ght8My3TKi2L6CFisSyxVrb0q97MzNFXa1G4f91/Vi1seQfcfBZbPuWPoG
1t3rgVil/L9wOYZ0+6cbVfCc/ndI6s/PRHWHjefRctxCNo9gsq/rj/Ccy0p6URH/HiSUlQm6Oorn
/e4qYhGY8VofrpSzDuqSjxIUTm/JV7c3P20PcArioeTLWbYh0vZJPWtZVxLZ+99LKPZOTRwpuI/K
jSvq24+LXQXAZ3E1/An3EYmrE80r52jzLr7i2b40GIC2UdiH4WnjC3prHRfCVCvNnROlS68pQo14
lNdj2lsxt4KEl83819qNIcWax0evefssyR3i5jVQSY8VbygTqCHTF+EAbnmjILGDPzCtdJ5/2QCT
V3S+vqbdb+ks7XgFbhy8v1bhRW1qL+5XjNMaC8vyA1JDl0a2Pyy+MGRFEbTPGT0Ghu+Hp+9iOeYl
PWe9TV0DrFvRCp52JM2ioioaGH+hvbHiunDTiPNGq4Y5pdUmibAGRKFNttluDokE7SlwtgnppiM5
wHMOoqXOoyc+P/VDk4iD8cX24gMX/WQMtlbrT7S331oK8QZj6Jd5Xu+ej0m/FbdanNbV+ntl1ep3
hW2LQI5rRU4LGrqDif/5msYAgGV/aJXEx4LvvkFk3sX/EHueYkJnNRTiT/LmW4/aa28tcMTNVIO2
XZG1ljZQgxlB5Ia+UTbXycw7b3BVTQxx4/Kbk3N9gljWS3PSZ3NsEfOrY1uhjIvKr5N4r+KhEdHA
nx5WZFXkkZkk8NSj/Y4VyGW7C/jZ+Ry0vqr821fydtx1GLfgUExeyJZXE4UHFlpImSG5hc8tW3HR
W1JgPme6w5hqk3kQCjerOVWZfFLvjd5iU0XouD1Ad2JFW0sicBp/o+yW8/J98eogZvByYL/ybwBI
Rt+WwDx4q1z/dpP0MHZwvIke3jtLsTfbJoWsn6Bgrntt/fNJDj26l/605tmN1hgcIWzq5hbQY9ln
7lq8Ka94KNHD1r4L3seTjvCFlivPbAK3n18TKpMuH7LPl4ELymP6/iJnURkzF3u3RjWGrqjBLfjZ
wSOorCSvmaikXZUT69q4mqKvcQewgPyGITe7zc8rUDFbUNo06k+v8uA6K9rHYxk/YP1b1efXqQNA
qRyOPckFYyqevYaFb/VehQuNuIl0FcNU5IiqOa6IDqsMjNzS+ZT42v6cOP/2y71C7we2Ji0lSB/D
RI4vg9mxThFy+1Xbudv02UV2wImfa+ImcK7me36IWEs/3IQYhZBd+XLG5sG3kIfVMhAreg8toTxF
BwnZs28uJAOsbXWbOWRasvfio4R68EdJTNDsjzBlZ/V1v2/LwZpk43HvF30GPidf1MCbpSYF16/m
STiAe/QPqd3MePpRyomqcAVCW4haIsXJg0vA6vgHG8BiT5Iua8fR1HOTJ8NhPW6bHaBa4c+G7y+G
KnsO1BmkzI/+xmXYSb7V3j5E93uLraWMsGNoTmTMGHb6ktdd3TX8iAe7YCGG2bLlQ5Xjh9FVs2LK
FcPdsR3KCDcLHpE9vRolidoQ6N8KSK1oAsTz/V5x3QC4AYoQ2jnkCnrNzsGMWia/Wy7L7W6xKqHB
cM1RjdZkxrmBPR4KbydNUsgEOdIYMkR964H077OVZO16KqhcnODu3K62eThjRA0G5d3MYS45LE1H
IYWd4eeqt3Ep3SVqrhZR9D9FasapGwF1Nqelexodp9a151KUyc19+k2snW+xtRA5a3+g4ECGAx0L
zObPpn51WQPe/3hpfxoLqn7c/RxI6blHgxPHuA0s9jhA/f7Y6yhzQ0Y9DyWZxf35bBPGRKxvIQBb
/kbRTcsLPSnnV9cpb2TMC9wklBd64iYJE7y1nP/dlnqFHj6d7tSTxBmdY/u5JvXX9teOPCiiFxCQ
+Wp82/Le2Ulo6witAZalz4PRWM9/oA8CI8mWE9a8mLIdtT9enuDIQ95qUctlrllyAwkq/KgevfZl
+l8cxVuAPj5tNDMNmbjliG8MOzyrQnMWCa98ObtbzkKc35nP36E9fy0GCdBW6y85dead4PJwI2su
RPf10s3vh7FpEJwuqw7iARXQtpVOXFwr3ggXldislRfS4B+uEeZyQ6SPtrWLMGbsmYkjkfxtwE5S
mybUnDASN3+vFSMCvarZcLSqD8DXiXSxXaE/A76h8RYs8DYWT0cYNhh5LoTgZyz8U83ksmZF5/dm
bF/ssCCK9c8Q/Hlbz0FSag17LFXsWvvv5YIWZ0uivirokoo7fjxGlEzTZPH6o8Kez4B7G8aWZ822
/Ym7/fglRpBikhiJ6pAdZ0M6x9ZBOQafVAGLuupNkaLauMgHaCOw96grF2o5lnKSuvbrXRIU3tj1
xn181jffwe359a4Oo4XXj+5nnJzQT9ZIWmL2OUaAAtHZFci/TNZwoaGLp3/cgGeOH/YW3Wdo72FE
8H3RBVxtx+Fmf6NPpnpIF+onETAqitffMgQPTWnubaDd98i+VtkFpHiAxMAdPfk2saT3n8d1Mr/p
GwBpjx7uoKrsdBVRNdiCrCtOAN93xONPZNyH3CenJW1oBGLERyeu8XCLlA9du6MZpf3qwe7t6p5b
WLNaa4XTpc4P7OBdBJf3hlQQ8iFR1orYBEEvhJ1JV2AWFt0L9pGNFghaTQKPy6XTnzdMk4JTdVXg
1hqDat6/wnJJTiMsFCEfYobANmtjmNXSA1LAw1cGbypXWMmGxV5qyukEbbL2fiCs9F/cKPgkfFL1
eVgkNX4+4ptrTThOh653DP8gFr4F0BCHbwSoivS6cnggs+f3znypS/j4ggK8Iem2cM3qxrgDKAt4
m9s2sVOCsGw2GbhB+WQIMEWEMnZVUqqm3nsUZ0BBAYQSCx9iL9Mt2IT3eqTG9YzYK0EkEaWP/L9F
I3t31262WBwtN9SMp+6vwN9zKeY3vkQmUTxs860YVqTQC99IsbxIElu0fBeGzwHJr0vmCO2PABgF
XW3YlW1BhRlrPAZU86gP9Q8XYvKgMc3iqzqnvF6o7Ei5+/NiMTEYHwzL4dqshdwn7n39k5nK9OU2
C/cXNHm3UrDJNUMt5OnkVN3m/KWPUm81+Qe4qxrbbrrSSdEiJSqBpYSlp62quSkPQTkxumbF4aLE
62rRy0tvMledFbwK5/cKEVp+tnh2UMpSeJw7eJkn6w+xxn2wTQqJxBPJadfhmzjvJN+TqDWyYW1S
ABIkCQVKNhIMjhf5G8NS0wZ//Q58Fm7J/M8q0m6vaFi35OQpXo1XpTBDLic68isCj85j75+Pq9gr
XKoXvM+fLRWoAjd7xGSe87oXMjYNzjAOlc0n0KcG6NxpwggbJVJh3s4AueE8KF4PAYN6aWO6TiIz
jMm3k7a3TZzcj5IVyhpaVnnsG7N+cqETIX9QMYZGsg7/Zg3S0smLwIcZFlRXA0txRXvZ2NRXfE2t
IiAHkfNa/wSmip7LcCRBTevgcd8nA/zRF+h6NuBvmFwLdMPqzJxhS2RnGjWz4m/E5rdoI1bv8fyK
FXL/gtmgD9pj+zqNr8M5rrdLvYRDQU8Y/9kFDMb8sP9ynZ8dhaiaIQXehIFc+akQT4RpstQwccKB
aRTL9PvIJgk9kqfZV1jeg5t6hkaxZKKhmdJb7HZEGORZ5JiE8HAkADO2WD0OJQnnXwsfulwrNxfL
OczDbd6oyOTbJcvFbj8Kxst7fegqVKJRoMv+WOvVQHjR9/2dG1FaUl2vkgwYOkqPCCpOb3qXZr0j
SCteXo/ItIcFpX3ZaqGww8yIgomaM8VB6owHKIN5BuEko5EhIWaoWPVn9+PA5Y/lrOiKW5ob8ayo
FjjqJkaWdI9QHKeleqkPjLHfgqSzP1+hKTKUVw5JrtA48W+dbRklW1TWLp4dKNOJcdAcUfF2b7kG
Nce39Y2/KPCNuCBsdY0X96D6S7Tl+CLUdrIQOImBVnl607oXUjlk5BkynLd+y8xSPs3OO5lozoW1
/Cjw+4ZcEaGyBOv0iqu0BOf3bTmnxHNcaVP4tt6nrmLbGLM1uj8xr4S1E2TuQWfjeeFBwlKgSszy
4vweimgJrrtZixHKnnH6TnZvwlqLknMePLW3LFJnpgVBQKXGWI+/vwyroQymQNVH44mQFyycX15k
jXfXWCfyl9fdOcnwIfQEQPlnnuTwazNBYHoCoAAQy/+Cn76DB9KVd9gBar2Ve91wGKiu0CY87QCE
DKP0Kni3ylwFiueM2dn0f1ncG1soYMEnPYzN5y3EqV7X+maEeK21KZjYoKIbxMO/znWtio8GYTtn
XU4WuEfnYjor2eF4PrJuMo8+KHhu2XAMRcoZBbGgv+/fIylL89GqPF1ePTPE/03UaHF3/n5YhjoM
1Jp4w5RT4avHwIEOfN7MfXliz3tncnolVlJoVDf2CNHCsPdOUFIE56WlHHDgsGywTwXNO0InL9dJ
34R2hzLS2Z4lgzJY3TlI4oTrM3Y9BZEGawvQ632PnLMRFRKnd/pQjeJzoy/PtoCAVBmCzC0zOU52
z97DmWtbogVho9IOc+J9NmAU9nq0iht+pvYiACBHHczPS7aUkTMaQZlSkDTUh1ZwQARPhHySmySG
vkDhnuDkTpVgcsfQkJNXJjcdaf+BndDmJ3bM3fXXGhJtqHdf4vmQT3M7iaNDfXH6G490AQhxY1fB
A+sGzt/kgvtMujE+7+rOn7YLh2n0MBF2UNwRgPRevnQCBgBk6JO68QPwp+14NjDRWiRkMwVUtBn8
T0ee1lZZoiLWbz3oFptlEJUaYBTxIfJTidJQE4wVekIz9HA17Yn3vpillubt+3QEAwnMr2fcwgzX
SFnJr+yC98IBlDqmcCnAuL/2ba2ZEqwwez/JOD8Ycu5ZvctTktRf4paHNgveQasNIkk1IhmrROxI
Nwoa8ey1QG0qFXuoFUdw1Kh9TI1Aj9hQppdFvLtLCpYo//pwqmF/q9GO363bB4/gU9dvaJBUy7Bd
f7dfINEw0P3+dTRekaZO8OZvDC/5OUdBiHbGtJ+LRO6incuO1dFNg1jBWSBtp5O+ywvUBSfech9Z
3/C9xVR7SKQYxnIZP2er/QCSWY9I1xDlXEO7Cfx7+YtctSz9116Kg4iefQ+GxFV6qSxKsNZlgSAG
SWgx6BeHSNXT/WCa5ohMZwiTEHdrdHDVlAaUmHUN5Z8hZ5EtPqNMsaBPCmkqmFaKGBMshD4GKKa9
FOfYe6J+Y8GOo/7XZR/87/0rSXDRaRawAjP5BBhdEWBww3R7whDdvtNBETmoblmtYDZfthIGMe9K
GyGjIhmGFGxx5uuw62gWqK1W5za4fVpOvZ3OACYFCPhgHrJF5Sycbabe9AYYey6req4AWH7MX8Ry
ImhgzqXx14MR2umxvoW6noqD6rM9conM7v0uwLnY4sOHhlGb4CC7Bw+XC23oVTTR+zeKUOMQ/JTl
uSvpxdgFI0X+Qvivp7yoxuYanaBpyVsBtxCV2HD48u4VNWNpZVu9ObOj63MHYScyOBwK17+gwy65
MZjgmEDk3kAsFHElO6ddKNeT9gxo4S6W8eEPOvfaabwbHQU8Zr3YaBaMBGICwSiQJ2RvH5zk+m4p
JIOY6t6LjdwcXiZbX7GQzfMuVfIM1Qmhj3X01IImVQuG83+b1XSWcgWuqBCJt/wq2RmbfHFqVjyv
EwhvxiowdYsMUQxpKCWOAK313mgO+xO/UkVCXDCT2GVakfqc+KWJlRKDluow7mBVoAf5LcTfcfDk
TCl6JzQbbxUGmNhWYVSgq7OJQvaROMUvmL63JP5KI0hzEhQcFX2JhaBuFSw+xymvkNgqZDbGLelG
yK4LTT2Yf4i436Xlk+9RWrs3WCCo8fLXfGyLJt00Vcgmd3BYo5PQ5XZHqLvibm5497ny2naayuf7
gOgWn3SeI/4zPagAgSTtGfqME8RR9UpXv7egeYRIqssnlxnO8dJzLpmBxdO63LKQZkSfABa5mNCA
NCzXLZs1fT0Nt3JcUtXhD6oTSnJVsH5G2pKGFX9/QGCItKHdBD8vqLPhO6kSVmD/hh6LELw4c6ib
VgrRiznTC/pNVIUDjWHCmdthMJDefWiu8zzX3wVTjtQ/wcfhlIsZddbISJkZDpYvjwDuFdy2KbYE
VPR7vesGnmt/jxihPb9oFa5yWh1Sh3yeS3AYXzZWgeqr5SoE8PdbHZ675igJ1dOlZKl+RFkU+pl/
eZzKlubGt1/sZdMmPJX71w0f8wrloY0oj8Vk+15MpyfPF6Rqfd/ZcSDRrKTVuwE/wW4Q8G11PQGY
HFcrKulQEmG/ep9eIL9ClHCQB3JV2osIyr/MDxKnSDzYPph3mvLTKyPS4iJosL3tcaeZ6zzXja/n
qjrGubAJEkx2ISwhut6mQCc6NsGVsmZbceWjlBvBBbt0SR5DxAcHEej0GhT4krUY2CSWXQpC5FNa
dvAC9S4Jn7j4waYeQfd3/wTTJAMh49a2vXxcblrsFX+3mo4URVHf+XhVgy5TG9TIltaU183ioc1h
f/OXAOVc/q9zoNasBVY+6F86M35Ctblna5oM/VoXgVkv3ODy9t9koj6JXt/EABRgYHFd140eN7Mc
hvKOopXpILxJG1mp0WsxhKNZhz2pukkeLieitD9NftT59rf2cc8PlLW1W+GAZMKhx2TU9vQCN0XZ
fa/tAmbpfnXKZRqT7SadbSXN+lHVknI8dbnnD9vgf4TTdILJ/VHcKpnWupsIWfDHG0aP750JkWY1
hNpnqVAt5uvKuAXuiJsGPpur6Ts83t+A1NsieG+Xc4DU+AV+98pTq7xSanbZuYU0kLuVxqoPnqiy
esTGyhCj8pQlwDMQAtLO4e0ZaYf52sNsET/IFkY+RICaphRtOlEFF4KbzaI8XHj2aJlCMJMGHS1c
3FPedcOHLcazq4ORVl6mCVrhMklCkOddFe8XVLAVmJrSU1PyW0bCwIgiMfPwjR+uxKFWkQExd+7E
TTlOYV18wACH9+Vb8zi7aPmQy1kpJCl9ByTD0OSlHPUU9pDK3AVimDZIdJE+Gh852kkNO9bvyXmq
GhNl/98s9H4ecJDMpmbiqKfjRKK20BGrADBDzkvrWZLOC7aPdHP2v+I/yosjNRkvsqPmTXGU0cY2
EAiWbKFUagEB2grMZbq1QQJBiF0dWv447BX0tx0JY7tiGX/PtqcJrPdkeGDcOiBtFTXdv+e8/lQe
C+r23JYFpNqUlHSPy3NjV9jMDJwEmNH/nSTn1hGQ5M1hgQUPcM3VZbI5SOJh0gXN9Vv6SNJ0pCPL
gL1XXNTq1atCLOarxiZqvJ69jz6ayQJRFmiywTv+OPRLcz/cNN7lSyuE6JfNZ6cbzcpFEWATld7d
crrPLsIiJLMPNFwXP0jd6vhi4XucvCSDThE+qCx4ULeYBB31iW9fY4sGPxRnS15A6ijY/SGTQbfC
bKIUPdJ4lHOGYceYQXGgAgMRjjzM1+ytcbYAH/trNNsfXzXbJtY1UUZ49BOsC2sta5ATu5oVJ9bS
MJ7A5PaF7gQDH6X1UBedIgd3004Bm8XSZgWTuozRCnAPWZFndTuNivWYGZzDRrSsLePtqWhyYsF1
RzRJ56xy8hkdeJZPofzT5cCac1KFCyXbeIOX9XH1edBgWt1Zah/JNFi0OiD4HAY9IjR67HVWJycs
6m2sdV16ccukfdzAw/xgT4oMphlWZuBmqoo9+Hm+2rNIJee6ZA6w6cPCRHQEUrODMIC3yDkyRHWk
2xgV6KIN34pdEIqkA30oyEftiNPXjkLQhRJJgR/9tC0kCG4x/jSrOHw4sgKjSomGM/eCBXWUXCIQ
W9fMGDxFWVk6ABum2AZDCMoCokbffe50tjXAnvZH4udw8OIKRKdm3itXmxcItw8uTV5w31mNbfrS
NzDZTfWwwOp3QW/5z/iBjXweOm8EFxvjMiAxhKwU99H9t98WgCL9TD1qv6ne+K9V/oRC6kCI2gZ3
ygqBYD+HxvACv8n9JKe4e8vjuRa8KH4j/uU9kQ/fjZyUdSxZEKtio/wylwUySzv92NH0llTXoxYj
YRSZ1ei4xmCjLA6JUyAiC9/M6YSaMUNVP0yCdylVPZB2GwBJ39NExX2+SnSJS3MzCNDB3N8t6nK5
Ts/bGqaYcAxcFREAo0LaxxK41v/BxJzkefl/VzzrXaPIT2TRLn8/TH4v/uu2k0lLstli3H1X1KZH
1wu+5qSkNefQkhv2nXqIhgY5VeO8dtLRKQz2EFgSGOkU7SN8yJhDrQD22qwzY5EpP0ixwqmAd+bQ
vyppZVyI8D+YHn8UeVQ127bWSpEdt1aV/k4fq1rM312gyah8Sk8ULJL3H+4EhnaAwsU0s7eAtw9s
bL1WHsIgehTWiulv7a9SGO+25QTnEJ3T/iyFlCFsBPeIv7WMnuV3cy8U/nz/BHdYF+OVFzXepkxR
qGtpKFSwFYjsB6WoT8s9DVbPABv7xbmU7yPrZKkeIXlAhMZblhghgZJNZIa5o1Qp1OYAECO/frb2
bzgYS00iaV+6310ZvV4CfRByW7RSKDk+H8SIZ/SQ06L/hwJb14424ErU7DruX1t/LwOhcpE+1hyV
mGqc9BtTewbnNXCJNGn0RHBwp1AN758cLjQYrXcVpawkUPYisI3EZnUuc95nJgltN+8i/J1Hs2Sm
eQsSp8VkjKjpSKw8Lf9/YCaO+dQvtQebF3dwzeBKsUu7E0HzG7dSBX+pI83FzSbOszLbJnmNyZw7
93pHfnaAYREzoN4C/2w/Z4RooKY8p0oqEfUWxekHKW5dqVhW4BsJA3wp+inYeJ24BJHpRY+4/lZ6
VknGumGcQiAAqgQu2xlrphDfVKllovyfc02oHOaClgWIfEvY8s02FMMUllFE/tOY85zav4/zbm7o
WsJF+hnJKUfR2o1ANbfrBpGE8uGH8xmI5dbK/Clgh+DCtzHZHiquUQJYiwzGzgW6AMd4XVyn/ahB
nnES/1gFiW++fupjDaZIh/wV/TlQi9M3eVhxeO6tiLpZ8nED616J1tHTaDun9xZE8l1jIZF/GIE1
Geh7Y26z1juxRX0FykZW+2UHwZJkZu42GVsPMMj2p9dUcRtBduRjwN+6DYz382/McL7pOMXoeHB0
e703LA8lV1qK88gpT3JvSL47qv5tNQi1XqxxXwEnbPGBpafQF3cvtcoawkz09XdsnIQhhvhyJHOS
jJi0qAsdA+yN98qPAKc93UVRPZyDMu5AlZK9ByptjgBTFDHHPqvTHGJdzJ2Tjqf/097LJs1INjvU
1mcpY+MQAyaVSKK+wd3EEIj+ITJapL/mEas4w7J6VOLQHjF7wvMjjmBJNkeHHZeFjbO7vqIYhkDq
MoHF1Zy066bCH4jHrAlOS+808u3KwpLkarndBKLPMBK5eotXOp29lU1UszOIIMUTi2+UrLO5OjIT
FpBueI7buqjgVWzbCNVRNF6Tn+UDQF2Vh0oPUeWxvuokSOuLtEt9WpWjrF1rXDvUf1VFTos8n2Sg
lM1J7yga/bOBmKB0ozDCKXQa2YYRYCUt9hN0Xp5WqJLqm/bpSTYg8hm1w9ZQFaKovppaaRuhLhIH
FeBNaPD5OGn5+656Hpq47XmJi/X8nNmqRPjeGiXr8lL2qhJcaKfL199OuqcvXys6LOUSecku3+TT
dnpGTyaRF2cFVkJiLYosGqVM8HMWQ34fkiRWYTjL04y35bKZwTaIIIKYxVViGKLODS0hZmTTj3B8
FOHU5Ua5lUzOf5ZP7Qp0FigxcX2oDU4pqzqSlaEM4EwOUWBaVXW3cLJz93eblbG/i5CX/x4dfUnc
7LK6eXLfQyVLobdBHNn/0mAdqsyMuozB2KC3k+aeQiWm1AFLsg10fjWRQUnOD8OFO/DsPRQTUplb
gj67lJAhaEexWlZ4UxRubn2ZsewYx/D6AmkRjW5msWKqIIHOq4VQS8mqF7bOjJ2Ur9VFiBWry1XI
dKdBp0x3NxJBwEAth6FZ4MITzC3V7tSa2l1lZplQ7AAFmJxksBYGq498yk2l73S+DawO6xfYB9dA
CJLINjTt4+lZtAo0Ledjr2crFYtHFZ9zAJv4P2CjzxpkfzTtzKW75Y+HgrzVp2rloWZaFadWKB8U
DVYModdfYS8EvsYRdkMP1mld0uxiSsMksLV3Bu6lNN5ZDmNaO2nV0UCBYscq74w4+N330xiDb54V
CI6rSL4U0kF1g4CxWbe9Ig15gLjvL9j4jMpcMfISylYb/nEE359Rr2XnBIiZRIM9QGiQ5wrrpcId
UHdWpt7IQW6KQ8Y6dFZArIKOVt6fBDs2n7CoWgSZqJhko7/Jr7xkxgEOdXyIcojSLQL+YTzKBFok
OdNXX6nCiaCGpUjDiuflkB7ngypi1aukvLaAshUjMbIwMLiME303d6x/Z4ScnMreuo4RrRRkE1W8
81GWE3TXsLro5OZTP3pOU4nNeDQKgQlveMNF18GYSdeQbWE7TGALyB5sAS2HSDhWv2dLVHb93UFJ
li5zE0jJuWKk498+eCL23cT2OWCgMbW2+8DezV2Wwjp/+07L7iFCRF8Stmev6FZBj/cW+GJ/A4Io
6XYteeA7rxx8O639T2wsARsAOKJKq8UxRjgTyXJByNvjP7ekYd6do/UJWQ6hyIZdR8ILahLL2qxv
XYevzXXoLBimVk/drE8K3E776aDhlbhSaFfRzNaQhw3r1J+EzuvS9INh9XQPbhlF6ODF0dTMOftl
tSntIv6iBwKIqtYdOkjrsT92wMCW7w77ccESovJV6aTYOguYOwoTV859+T1JbY3JtOTmJKpQkKja
nuY7YxtH85VH+teGyVEGYhOXsvfi4Q62BE7YISieq3chjNdqzaMCnVnQis/MMM8JBhPJYpKghJnD
eU64/inHjX2i5kBHtJnW4g9Of+Cpc/NN1X7CZhtRiUCi73a1pW4NgHjc1J0U/fzkyLRvMVUJMh5/
NXPXMFJM1+PbaL9Z4SU5Lsy3VnVzRqyB2HHjmgiPR51ze5b3RHjALxclPpb0kVOQj6k5k3HVTeHn
e/379MTy8WbZXEouSlKBOiLFv53TNFaM82QuWWG1P+wTq40UXzvhrY0+NjmaQZ6PG+Y1Tb2e43oa
trO8Tfu59BJExBA+70vjjT4uTyMv4mwhFZxLfyGpoFSZBxU88zrsl1Jnzy4CpgDXPTJQo9FMTYfX
osh4XiGrzNnVkMyn0lEAOBfW6YzK/UGKV1XjxNa3rBIjZ9zhyoN9BUlzGhmk4STnIf9enQnkvIg+
puZAfb3T6jeSZM+dbjkcIIE4OdM0Y2FjtcbxjrLUJ/TDKGbIetRWCZNz2W+sJNqmK+WyDYPe8oDF
fNqI5kVTOLQ0PmgvUc1O8juW7pZwkqUT6VB9pSsKEMPZ+/mOYwIMRiunzZm3Zt0tKLUMv2i1g9y8
zxMSWB/UG/UbgxdcWlp42OyS9w7Laz9rYVXbcx9eJyaACZ8ZFBNb9YcEQiEB2qGB9m9QWdJITtN5
puufncBopIPFt4TA+1BmoTP6GNtft3F42OoeR89VbCoktnWBacTQybPUrymGnIY5oziR4TFXYZHe
nald8/1rFFK4CjabK3HM/fwyeM9LICG5RnIPu+Wu+WgD7vczVsJGZzq+au2EI+hNnJsUi+4AKQw/
8JpBKT6zcT0B80moRwvc3rVoKXItOIUsaTO5m3Xb+1HEXRxjEamOFHc5tviO23vMmVsBz7F1J8rK
7edsGbYqWhcw5TY22WPe8TcwwpOUVAJxBkhnXP7V4KiYI51NaR2MSIY60DTxgq2PxnHr/m+hzyWT
Ukct/uPh+96qCl4gGcSPtcYWRnK+X76yn+ZJH4RaSShllqtQ5BMfa87OOouLxg+bWSjGxp/HXKnY
3N/rsDK2LEEr6blmouTeDEpVr/63daAEwihJiO8OAGa6gZx3VCI1qBC5IjR40rgqw8MSND07pdyi
G3DuWXqPXUJ+MtTddDoBIiBf+6ZxX7FAWYomtvcdMEA3z2zxTpnMAPh5HGnHoep5x7WjdW0PeCwj
mqgpCY/VB4smM++YKeiBkoa3HS+5ExulkEvnhTJSK90wrp/s1RPh45yycHcSTIxg5h1pTgVY0+uT
fid4ys59XKeVR64s5mGoaIOqoRG5OIhAS/tBnXt8jK2txbf8rphvQsigxw1+9rK5VuGVPyXz38YD
cKxdfFAuAheb/kpNmLxNXk8TwSKWFoQKdtj4bAiqZNsJWb+Nk6r/XuNI8pOCNpIqzDpF3+VI7G5Z
r0vicweyUWaYgWoZ+0tncNjqwvM4lGP3on/vwqsP6DTXOv1WQg/Fhpwnxuuu0e4IicrXsu92Q4i8
IzCitprPai14NPBN+5xJH5AEczsT6WLUdcMYxVg0D+K2wwoKe6AuGg9ZKG1cZBaWrY3UJ8D54R9/
hd0wjxaAxYqBnFeYHAVgoHT5G7WGh3cbDPgNd+TeG534ofm5OXJNbEM985F0YOpdX3HqAS+N/dvY
ZJq/z6AULrDQ+9TkU96NFJxaUG7HxKjubfkg42OyrW3UDl4OH1cBoABUVYJYxouZKKGgCoIFIO0W
3oF54sPnoLZOHv/LMQ61tgil48kLI55liHb4NOrdFh3SIfdSqAJB4ZDNKWvzIXvGdRncSuVXcGQQ
4+o+S9HX9Sz79cznkpVMMXGLp9usLmY1wEELSii/OIilWhHS/pqK011Js0BmTMLt0PX2l8cLaCDM
AO5+BWzo5BjNhMwUdC8F9oVQdR3xkiGxDmGPAsXja63AEWRlu1N987oDmPcJw/nBesoJXejcNg+r
AIr0iuZpyC+6Dbruy0wLlhVo+p73QKrnvDnj+bOgAGHU179ta0IMl4DUaCW7sdxL2w2ShOmTCrim
4zyaYMZ7UDGdNs4G6iD9CwK1OSVSGJq7LfwAjU3eTJiiOjGRSwcpN/hTy7vA6V3+P94UeURgT5bc
rk9HXZ6V28cnyl76wfa6g5qiMAsw9jN5kwQBfOQhqiWnxdaY//LrZxnymc8dYgOakRMmdr83dioB
TSgv3sIu6B7qS/bRkkPwtu0RziRvg0en0SIQlIbu2Z8v78pC/GTYVf3AIK0drbKidg6e6TeBg6cu
j+pd1EVnLdoy0dGHVHXPvsXyDBjidI0SpT1wcZQmG5yCv+TzzWgt6bJbKZn1zr4c7raLfi2kMxCy
q0b4TavsWN1O3wsjeCVNpZkHycCB2Ct8/27sxtNxviUVUgnLfrWFXKC3wi7v36eSgQiSe0dop+ZT
23GSdRWWfOjqZpUfw/SJdC75QNIWPTGTlHm7+a9gW77/1cEF/Lt0R6Nz8xfBCDMZROA6FsiQ9hvW
7ocfmZcF7cekpeSadDM1BHtbFhaWvyeeKFqybj8zkGWd4XvHsvQ5Vr+ceY5LtpvYytKGTiy5/caI
ivknN8btmIF/KSMB9HIsGS4NNFlCSuMwnLZTUPl0joqym0J5GIIfnG/CQwwJFg/HWkMPf4sBZ+rr
SCiXofI6IO50ekC5j1FLhpMCLMxIHGRoSunNIqK+uqSJ20OCemZ3E1QaaiLfkjr2/U2PRbmIB22h
V2yAKg6swEgTOpF59m7Ji2dgxwp8+C5vtGdntn+kE5Q3O1M1sdW3bl9+W2T0AnPDeUTNglBqGGG2
GpTiJ2pkydFP9CDEs25vk4vpP/QcQI6kMo7eeIMJovZQQyYqyhu46TRPVdH+qa+NMy5NcAu+CzdI
cp/U9jH6UyIJxDml9Yfr85zNRVAgRN5okLb8Pzfx4HfG6v5JWKoDj5zsZTXGpPxX+wXFWYYo1Xd2
xlNWEEWY8lZYVMQB77V0HW1VCK/rbtuWqlEp6JawOLHr/QzxQ6mXl+dfrJA9E50MG/VwXoFyFnHF
I6YewysR/ka2pp0E7AurZnZDpnlbFzY1O+fZbRaYsYCUamzBANvPP/fHEnjBSp3+bLaHOGilWZVL
eBo9Uh+ISbXzrH75pZbAJNcifv1aEawjJh4+ChFRHo2CoIhVp0jTQBf5HTS4jjSOoZPuI7fMoSf0
rWavUHp9PXx8WefDXk1O/ps/RYIc5TEIwjXm/ZbnYX6zba+M1k4bxCvJQExLK5jXstAohoQZIPjM
zbmIV9DAzrLjegrP5FLocaxH9nn/SS++gBDqouBcxD4Uvnfk1geIboB8LhWzxsizZQg6fC3V5hiX
OAyKRqdxT1+uN1hlvTrVuhdDQpeOEJLH6/Jox5lVfoAgTU9PMbbeG1conuApTR0gWAcEZpJw4be/
KciDiO4kYUYf+oqvsAykmvP6taUXEhYiEFLWVsa0VAxfNGsHr0zOvSqDtaEmKuBZyDsOQqsatWmE
578AjBwL1yAA1KDhjOdpxfjWN3SxW00HcIkSFIbCZ90vShyrcuAtKyhBZmWx5ppOXd7O4iH59wh7
WM1icS3JIbXgJTlY04Il0xIWD8OsmhCvyf2Q1ktAtjdVH2u8MG/MidO+XJisK04oEDL6z0KhQS8Y
BiSbzvRktVsE2XgFSzgegNTZXyN7w4UB5BrWoxs6g+RHpABMJMg7E4P9JiMBVNgdRr/CtlhC5HQh
XzCP8AbMi+AgtPDUhNbvrtBjfZtRALFGy6tIl4mfJD07rMjFnD9k/wfv6xW6+NtzKkwF43tM9rxL
Q9w9rrWpibPlHrN/UXFRgizxt47AknBQ/56QxZJ8hsjQPw1yGkKkI/YVpdE26akbba0qqAddA2rs
Kl2UYNyNBlcjEm1l6+2oAhPkUnsHZOQ6m2Ssa7pipwVaM1AU9IcnQ7Frx1F0U5ej+HD54Hi1phFQ
7WNzG3/sTL/W9QX3rIKMri0XYMFj8fwWRVA/qkqyzHwe0ij4uI3KtqiZpiv4/pmJ0uXn/FImv5yD
Audt6COMW8TpkdzO0ldwyLTzYJM+FXzPrZXccwPJC+ZMXrImly091kN+3L2mgEDUi9YvZR7x+QMc
5PGca64Bf1aS2I5H23a4WIiS5F/ukbN81JlZ6wO36NeJDRanezH6oW0p188EpwMpjN2YbA8fhHeD
x8T/5L45ZgcSygvoawD82TaQpwWlJxrZEXkDzmNXJ3DelJFfCf5MyqkZIpvaBNh/TOa3lasor+SG
FM6oVWPs6Yhql5Lp4LKJXWGjL2KIo+VvnTfQ+VVaPGWJHwH6hdfzJDDrhgDOMN2N2iov8+I/xXZc
iWoYKJfPUTV+NLTRTsSd/ozhQDd4ulfgIQOvIrwFqa+8RB8gMyHsNC7CCTRXeoO6/dVDJHiyNkes
9OACB8YnARH3H1TixwFeqwhDVpFdNZceTbERPAx1ABlpublQ1TM3oNhOJj3VJ4TB4FN6X48DY2qP
rF8js++25lS2eETTM550s+yYVaCrPWLSxd2B/ufnxR3lNp2hzT3LoWG2s2tbOMXoJxtIofaoPb+T
5piEy2RGgGbuwcMmBe/L/sOLhDeiG86l/FqB5LnfGCALoKag7TM6wyVNxR4uq2ynjoMn3G0j0hTh
o4R2F+gccIP0A5BUqpxJ4ibIKcB9+n2yMT3D5Sszmxwo/LMTfo2VlYF2kMOTU95C4G61ANdI8veu
NYs9ijbEMM8cUDLLZHpv3i9tziDY7suJ5l/SZAqwTq3xwpQDjLRscZK6sDuHZWUsJJa8cX0JKizT
+lvROPUoZHqsXqT1gABKc4RT+7wZzbrUfh5qwMKtoNQJIDkpPO+tYf+7gEZ3V5VqASqWCbtx4MFv
u1UhlQtrofqMNgxrX3xSGIr0ke6BqAVqaNmNDpyKGMbJSBCm232V0Vk6IxkF1nILiMvWulPwyGew
FWOaZxR74fdTwIHfOCEJmgPxcq3VN7NJ0l9JfGoe6PnYcjQFbjaQPHFbOl6VNkRSMZjaEl9imvGr
METalLnnd7AAodnX+NlySSTm+ybGsMzSG3nUbxhKOkFHhCWr067qYCfzKpMpr+cilRTwsQArTWVP
9DL3A0MbtXl0bisPeONBzdzdYfq4FDIGpv6UpC7zSRgrqj8U/42+Swx4eANyTesZ6jftJ0tIIy6f
f/+aLCwXojgvR//BHLxfBkxD0fCeoMkcb+ItxVDTAnAAd8/0jedBuBU6XLCXmF2B/2QpnE/uirDM
ZqudS41Tq0b/q2M9tUqIr88lVDIihAM9JD/nUcperDPj+nBKP6OtwzxT8Igh16AHH0yyMYGygpPV
jmXrbfxNXzR93Wq5UlbHjveW/1arBitNNblIEDMxa4z6Gs0EaMM0YC16uDeQiqGrHRiP8awp9MO7
Fvz5ZRcTHiTk6EAQxH3Ph49jzsNGWLS7IDvp0XEaw9DSvkDkBXgQhaXfDPvf6Z/hL3BJOfeMyoYH
xkblvuuNJ88Qc+k+2fsxzBHybLgtpGKm2hvxCt0Um4JNXeSB7yLecOZG+u3r0mSq3ANKWCbB/c8E
WJCSp4Sjob8SaXBIBaDjrlzeotiWOnxpd1bOeXeyDoDvrQEFOJXlFTENYybjZXgJD7EsvmvNj+l4
ow7D0GffmxiaJl9h63d4AHWKV2vGOhyG1F+k02GWOePXAdO5F0Q06sF5xfJg6Zi774mmPXsy5VY9
xGVYmuZYsIMOVSy92+kUF8qwrLjLjXEatjjxj5ggfvGBYpk+QCW1Vm3ZWV6v4WIyOt7M6GgQV8eG
VA//gRzGS7gfca+dIXvpBCSIqo2jsmEbnIEaFlNseHUaY7ae21Fbw36xWYyUbosUL0mRw9korcRr
TMd3FCAqAIq/KEDhzorEw6JJJAyTGXLhFuBiElcXm2lxYC0QYl6XTiGAPkuIVAcoWdh7GNKXpjCU
rggUHnIuehASz9wBVQBtmfp1S09N6egqzmi4J9XD5CoLvGvWogEBC897sdmQqHUVbeigXBWjCJVB
S1J4rvv6Kmf89pumsD2/BxI7EbX3NXc9FNV0NhG+c3OlEiF15rabkPkSNDC2T64aQdRjuf6PGJDz
EB8nliaZZImNKsLOsg9WBMS6GU6XwoGkx0HIJNBUk9N0q76CqhV91QvJ3I8T1YG52tPG4ytG5zCf
r3EsV5HqtI44m1YHJfYW/MU2iwxxRwMXNQQBP7zcxJ5weetBl3a2x3+s5dU8Gxz1QIWLZH2NBoUq
ex8zxFdSTDjork47g+g19YiL1hsxf2qyeCHZkRVUTKQF/pMT2rg6auSSR+nGag1KY9xKi/q+pMk3
PNSs0bErD7qGLHRwMfCPkpP/SiX+TrpnCLW8zvpuCHHxEnOMz2E4XP3tZKQMZnDvYw0Y3q7ejLRL
M1QXSkDal2E+KEGeDYO5SEKEVcQs36N92J02YM9YkiFD1f8HO0bfJOFk4KINFOCU4NI+87cNPZCv
7Ls3bZJaDF24iYKOt3JdwHQ6Y1I2cqpl6ULDBp0h0S6VTn8bXTLd58QBP6/t8K41oBBMEtxGvzUv
rK0O+Mz/CkRcPxiZa5HRnlDKB41D1l5uoHlCXiRyqtwLtk79tHGOms6yvTwT+bPPAfRLKSei6EL+
FZuQPMj7e6hl+lD6bPtGfFqetn79WlgTfb1brku22Tsrw0RPNT3pH++Wp/fqBbjyXS9BZxQ8zWmI
p0yoUo59T6v9jX3yCgw3oNJoA91bLj2NeZrXoC9psmXkR4JFsioXNbDndHokQFEOT1VPUxdGrJgZ
NLVkT1dXnM2Uqv9EHUQL/sbE7ToozxXys/8GL3dEgr799laB2KydhcT+8epBugZbd55N3y2+3/4H
oHLdGtAR/6o+3mXS7MTKeun/myFVeaarc9XqtKvDlWMGvpzeoS+xcIQvmBdEZRdLFpKTUSdaKQ0A
rTBu2q48AuOfEg24JmkZEcMfIMxM+2FJ0fn6ie5WI4H1FFLE7L5ZaIPmsd76Kd8jf8q6IMhPaaZa
lm4hcnqUOoJDYhlHZvQ68AjFtQhDaQgOsu3D0Rp2zfRjk7qBQa94saSgXAlfPgvHSHokpzvM2+am
enzo7oiARGG21GFL5jI5t7nZSKF6Vk+eJdYXEsPtlG5megLQalDbEckwLhjIpCLV6QcMmU2SDX+1
yMnJG5ADnNJRYBZ9LE9uDHYYK1PUrlxUnZiU+VUcrPp1T/hP0zF3cyYdlPmBSKCwM2zb1tA5HU14
Nzxy1kkaLxhNI4EnwLjY0dd6MBbfjIFbyHzBDlJJmPloySp45XmkOSFiCOH6DlrpIe+6GIH7iWGY
NKTvyjr2/BMCcAfT94iWYPB0WBgLZADxbin5Id9rZGUQOh8iH055YqYpMvD2Hb4TqHjrV3OGm+Mm
znpOoM0X7vf5LTVWn1p61MCg2270jGu5GBpBul17mIkVh1gfBHD8YjZZU4BEmPLUqNac7zaogJV5
OccTsne7FUqBqB7ok0rBM5v/fgkxV9vLW1JjWDcFItv+S3Zb3rJuYtF89PmOeImwG8njR7DbE5im
ljvkSgUP5i2i3zYGl6JgciE23ZWfrsDPgwex1Z37uHA4IpYf95uZpHNfLDUBISEKSp8/PChQQcDL
8/2UT/WfxLnhmKrSPG9JWtxCWymg8P9BjDmaYJeVnutLc+19fVrlQVKURKC/QGA+8vGUxhyylNox
dc6tsnn6o66uqm/UC+2glS+ypK/UpvjAeRgYH9Ejaa30gliSDLXYj/o9uV036CAiNoyHmrc/uetm
LYUArFlCm02Jbrss70S9nr6QUTvdAMsI/WkkfGlBx0VJizDQuQH3gH2EVlgij5Yt/GSVCW62t7Qj
/O/YlHtp10EHMMawnCYrlDnc+mF0hZxrxlNKIgjZKJ8qDgWKhMArVDA5QIQJCb3B4++6e45saQ4g
aqcVDB3/2sXM8thYC9ts5G7+2wYne7Cd7h0X0eNYo5iLU90YCG5f5sS+RW1pdZjfjcvbaLfhtI9J
88daEFizoBgQ+xoeTChUEVMHf+Tu5F/yup11x506Nz9HupOgRB89jt4XE0I3OqDSze/x6SvYIdX6
DsEEsrpc/XKyZFZ4Hz1qcgrM/KR4UODEyHbHMhMPsFYHog+t7X3waxK07eoluJ5EpFRPLeHx4xcr
bpEgo44msM6HNOA7Y50sz2LHxM4Xl6rI4EgwwvZcwckewBq3if5wGPEnKATrgI96PvlgSHn4Hw6y
fZLL6Sb0nzdfYyBTFW/NX5ZMXcDjBu/BYNXcbFWHCsvfU+GJILhf5eG5UOdSSbCw5pJPGDxxVsSZ
lirONhoEtMMFqdIb8zjFL22HE3mb2HzzkN6SgD9sGj1hcSqPCnPbHQ61hWq3a07q3GZwAmexB207
ZaZbOTOCXX0bxsIr+tm+Dgz2cODJNV58an5BJ8P/V6tQSXA/L7423HZ5wvYMP4cXoui5kPUkdCcd
g0+PPCBV7WJTzCJPSj0qdqOazI5b8ZKLXB9zlMWP1tpCr8rE6gVWZzQwidSsJNVPrV/aWhGCgi8v
DhjvAtrve/seHlghl5J5wRRpfLFe6wbqgvGcYZr5YBl7MEfRGpyfp9meEtrTNT+KAd/uFdPywQ/U
N4uLzzF6/P+nTMbR5VVArxE1bou22dTX5EPg1qkiUjNMKRFkLv+KOJvjuacI0k02oDfHprC4rD9A
5RJ6IODziUv8T7/k3Cq9alwJrPuDoDYnFkYETHnijMb2BABmFah0EsfaB70PU6hF52L7FT37JMjt
FBULf0g1g843pIw5kRrZN+aVgNPl2YDkTiA56937W665x0oV1QRLhy4Wtx3vCjocYv/7RQjwEGkT
qaREpluxFi2lH9kZ/9uMqACwKVdHi7wpa4fD4PgpyOs851vF8JwZme7TFc1Ae8NAhPdB8SnrkzXd
L0F1XEZN8mamCU3uRm/b+DlJM/IuYi/+HTddeRQtZ4a+5P6az+a+grtTOfHTav2lBofAp7In4kle
++bgDXN3aLFdRUEVgTGRhdywMCUsCkmj1KqIMQnsNttp9r0BI91RMY47sLDnaCU6ucjD0+ISWct/
wGeHHdQKTTJojYlXF9yvxQ4Dv8ByR8p2WETn/5uY86Umw4QKEgRBc3zmFb1w5Em8HPb6dItj204o
G2UzdIWcG+wmISICZ7j3yGegl/v1r5c5aCX8fKOonzl7vk1hZJkVMAgf5MP9+YuXcTTRuQxzLQGa
sYTM1EYBHFxCrbTQ4OUWMWF+2UXZgPRGf/fxCrJDcVNdTum4tesJUy4kaubB7WyU13dJ0DPrYuEW
4AUwiSMzlmxn5Glo3WbJdpbrKtJGmB0LhdizrJj3HXbq6hIIznbze1h4jg7zFSFHKO1Zqt77hMx5
ziJMjhioYrDIx7J7lvwo9LO0C4VZmInhLfGpkk7xSpobt7VjrAeL5MZgN6E30zGx4C9sjdNBsbbC
0sifN0lr8JmGVXA/d6RBFK3IrF169qx3O4dS99Mxo7KgTiYj7yKVtzJzQnuEFfjZ7iZtIm5FDh+W
QlNFcd3aRlx11VZUOn1TxhtOhLOjvxB3QLdDCNvf0y89qlkBMqXqrYtkGkqVp55d7mCWidw+9jOk
3w+22BBHCcZYFoJFXSBv5b2+ZpFyBhoyPbtXnDIZgDl4HGQ2mq6eXEGTBfHPmuq+9fc3jMdv0jB9
+N6pZESBRNDBidugiEktfYQP0Ybm+VS49uAu8FUDHztUWCZwUQ75BjvR3pYuEhcP3ViuvDeYXHIE
CGmSt4MyBpT+fOVSRPJWVBRK+6iH6ueGdFfNpmG8HokaO+nfqEvc+U44eB36NlY9Bit7bWCvjFSv
Kv1OjbVQkkGMit1OGCPj23Ef9lFgwGqPbLNJnbX0Yfjj/7OdWn7rHa3F78y1ycF/XIfHnFOOkbe7
6hQ7c3mLuYaegy8KTGxJfqOZ6Qx8uiu7NPXopkmzTeR59/1h5+D6Cy8ehg1gT27uXdFDOFRFBE2N
F2xluIc7xJ+p7+VqbJkRvZHeR/epMo7Cfca057m6HzThk+BSz2z6ZNFRIivaaOc3arhWmbJ4hzbn
XFaJf1Ht9ahBHmiVrLYA5XNnOQeT6LNsPprKpRREsd+bQ9LOkYyB32gx+9UvvNopEeJqD26PfBSm
STy8TjlGAlIzPqLIm1R7hi4Uaz4N/Wp77zbUY0QxalO+crLnKDW8uUv2fUvaM23qqqr9IhzDeBEM
HsNfDUkXzSr+b/27tYFa0VMkWw51NASCL5O77unUrldwna6adU0p6VtLhoO/yi3dT5XMN5aDbPT2
U/rw1FopXPLnka1fn5DUTMenP2GfTBzZ1W3rIcXVMzTEhZ3Y2OIAkuU+zbcDgSv7GSKI5rZJfh3C
Ufejro/0KFITlQFKIW6uInpiTdgLRYNtXjVmspue0uXvroDNGVwTEQaWlB6L+hs6VZTj40Y4tiyb
alLwI3xWAVZofY4no81B6i0ijWqEig1W1qcvouv4FDrYlgzmFMW3kCx77kIjtFw2zphjdLLnT5Py
0ke1aHjl89kCOKuygzVFaT0miADRLq58iXYYNkZQdAuesA8c5GIYr1jzHaTsxFcc2H7LUJMiHEXM
YSTG0q8x0lB727AVBXxNvTqnZyaN1nmWsT/ntwEibiScvmqm9SmEAd1khdLeWWpl487c9JWYTuPj
g0K96pO9n8YRS4MaBFa8/wx/fhinSep8ZVawLkiCCGrIC18KPH7epSyg6SbXPl+4ZslL8tOerW5/
ipweeXyMnNLUc8vihcTSUrszIOA5BQshHOMgjCl4c3NU07DoaSir/GjEJj+rk/gSBRKYsCjSI23+
2ayHBaIrCmWvi46S0O6ynKdBFey7Nf3rj4zT5xoQCetApIa1PdXegYvwX0ktsU/1KW5BaLNkOsod
T2u4xNE2slQcJaPTC6ZI3+MmrFSp+bIm7G86UWg0WK8SAhhzoyvJSKHvme36/od2gcdXE2SJ2rbo
Wwe1Lj+kH6ix902BdasIHUPeEME2VWwDyjKDEuaSH9QoElVD9X2jsq/mRNefM6IM4Vqx7hx3pYpF
7935+0ntqBENuc0ekxiybfbspPsG0qpuI29tCgEbY+xu+aFBLPVUjkacm/D2t9URacoNVwSIPA28
mmhTLKtZ4JzU66zCWOl//YkqO0Vpts+Ar6cAyxHz12vM5MTOo552auzsJPixOtGRrb4R/I9QzCCc
VVMdTu2AT1F62ytlwulSc/ZS1E3HOF/vdZAgDvjYzFmAm7na2c7HCLN3In8fdI/M14pun397Oru4
SNlhYeA/mYk8S+YRv9Yv68/j2QnDjU3SuXVcCz+WG6b+C3aV/YdpKfJ65oLfJtsu3uoHMq1g+DPx
73ulNrRCBMVOD9ODGwMbmbwyzlhlF/o4rkFb88de44jF3s+cXOrak4L+LsijkSXQGfFMxCOznVMm
4PJy1Y8ju4M3U6JYXk3pKaPF8CNkE9jVPPhSEz73cLh9l6gcMaZNbyb18I9JMpJe4u1+dUCWhuPX
o/S4gtFwp2JM3FOw7vMpHVoiqL1xj6bwtXhS6DfHR+SKIMEk5M7BthrxD2S69fIx34syp8IYrDgK
8+hUucdX0jpsvpruhkuPXuZzfjHGecDQ6CqxOkARvTpAJKuLUlYIu3YVh/p/32aYbOoxdrh2Xbvl
G2qeyDNHV5HuaOW1oVi1Tbp2moQpEU2VU4+VD9ry9JVShu3rJ52h8Jwa7fTcugGAmN8nM6rPtqcH
tHmqgWnQPIfa+bSBOgr2v/mtNx5x8rY3xdTdpx++MQHzlzHQTv/r5gSZEeIvHo0hPlCfv6Sr89OF
upko+NIcleHcgWOQTJhFq2i/b/gOhj4LiEDCDWVLD8oBui/Ue3wxrjv3QFZ/vMdu3KRGyRc0Cfhg
lVcmmKjC0hB0bumJOAntVK6lnOa7mBldWpMPARL7uj6umwfLAt0Gdjt5irxL8/VSW+l1LaCQNBzy
XJi/kkYO5RuKsTZw2oHg5O2+Sz07GQZEaOrBvYHEZ04UfyST+QZsElBCJDHZfmXk8zxM62gtV2zd
Wp/cGFdGYUmpV9iVl93g6zBeTFm3I90huYw0b+B8K2ihr6AFWx4oxLSmG0k238dy5vihLyeSy/HO
d7m9/uQ6beuGnSePdJVGkmIYB6R2ryiI1E9T09AcPwLmXpUg4uoT6N4UXsoKdzdwWD4bc5ich4I+
2eRFvx3/pODzxfo7+vpVZt1FkzVRjB/9vQnV8ku7R2mIOq0mGr+xRvj4H1E+teFSIWb7LT1ALW+E
fJbc460AVP9jPnVKcimB3PIzPmMHz1HkaMx0LAB2hfEqASj84JrxnY0W93G2q3mcK1Ts2ETO697h
m+mnNMf3QIgbvVlk2Z69bdg4anBbefeXj8pqxCIw+EG5KP8JgCSDuR5f8b1boDBMCMPedLKGDea4
Rp/PI4/3tKnuIejiQpOXetR4GJyJ6tm3m202Mvf3WFkRjxzsqp7/6Us0iHVtfZwO1HfY+SFhNBTB
z05XLUE3gN9e6rg0HaNoEJ+K6tJoDz3V12PBMuIdaSkUpQl03aInAIW5PbQ8FWzLUz2qskHL371f
tguOlfWeA5o7BdJ8UqMkPsVPH3ER3BtHeYAYc5ZAZ1IuEIHCt6aaqy6pbfsl/+jk6YL5YKA65BHG
dgZy/uYEIRdZo8k8rM2PwIhP/hljPCPcDpywYWe8ieZoPmldmA/GKPmSX9YtyXw+eO5VObTgzeKg
lP/d/maZXxPekewKaRN2/1iuZlmbRfJ4OZ6Moawx1ActeKMRcC8dAAVXYeOkxhvjNMnyrhSfsHlu
wYiZfj9J4grStkQe0TfCySEwv1az94XaJ++bRfqbZayBq3hZQwImM0MdYuASKKqpCFJYJpVVd/d7
Ms5i7p51MzBhxX/J5kjJ0JWmpl2b+aS+w5B7i3hEzvbb0A+Z6kbr8O6Nf3bnw/zvEPY9RDmaeTx4
QXsNgcXMFtcyp6t95g4xApbjwqMETmbi/s11NbVUoU2uX4z6GeONRKyckKGblnc3CVzXNk/lo2jl
SJS4aRr2wDZGrT9H1G9QiL0I7jVXKVsg9LDDJ8l2kjKBg7jovjRHY8qceQeO2F8EYQuu0kRmAEN8
gX99qPJelplmBle7RH4YoKHZ9hKYDoZQOE8rqf8NnObZuUpPT2iMiukTZMFZmF0AMh1N4z04f9zg
GSROKpAmxGYonwVz/n97A1TLK9yiumgYZkOihtxtiMvLZpNiEt5D82UEfusCcH5+Aw4ahSe60SLt
Ie6V961qCKvGVv1xlWNlemv15NsomPkxCgrP2EI2/XrRx2QXQFhaY11VoTX8y7HBjRgHL4AHuYPE
roWGPi9US0hF2nD28B/n6JOsTo3pB55Mhs540RQMzXq24QyRis+YHx70jCXyRmeqXdrRPGfG8p1f
441wtlsAiigOUiwbxMXS0HpcX1fSNh6tcVAWxrLqDcyGULl6ltCFGWyieDyLoodQc1NHTzo2wS0S
w2D86+37qjGWVFBdQuvhYh46e9474l5Y6E2r18mSgb1iYpbpkG/eC+ggHknH6tWNRT7apuvPz+69
kIcNWqOsR8+RfXq/5ipFh4bSrLzlheyxgcbVU5MMRHW81F+1yb1ekJUTsMO6fHv9E3rrsRkMYFQn
KiRRc1xgZCCdZ0VnNRQn+hW/F1tPsmeMKDPpl4SwZMLEUXiysG8vngYJjfvKNxp4R2AHoed9NmTp
f4HKXz7PcaYt4dQ/F3xVVM5qsFSZbJVxUSQGwBxWQBOIDOlMC0HBpOpoJDI4t6RlJaAT1EECps+P
+McbnLdfYiw+FxAh7IZHVy7JZ7oMiwHe+Mx455jLYpkN5nPkxyh/3DlDSSk/BJr9+/h16/SVXR4t
XWyrD7F/eyF/JzU0eo8ZCiClcPxqtAlUGUw1WLnIDGoRGjyEvDK9iClnz4n9nfLsyVvS9iARIo+I
HGYt6WmySpYVeqC1g5vu4zWyaRZrRoLoMzA271V26FeciXwgTFTctTY/zRbr5LY3XY6XxKiEKm3v
kTO8si0y5IGxvMvMwFSQK/zHzrtnFGKouJ5Z+L3LZ462DfWEg9MjuCVgcok2I2ZtuTCy5IN/fI7L
npEEp2wH9lVsPLsP6rPmAw+Zk4gx27P7t+LZgNzDXL1YxH77pMTq+Bu9hyMHxKLBfBiBNYRZlclG
ILsBmqZxDA6aVKkGLylYS/gjCff/yprkkNqJMl66a2S+OaUkFdIXDZh5fx2Uvx1/IAnYzi9qYxxr
ChZYDoY2XpkDCAqouibF26Hdbdohmllm0PjEu2rBxdJOS6Q85yQK9NOX5FZj9C1PQin1/Trfptzr
r1a7UDcGjcqIHxsI+y0ySAEfsVk7OPykUxTefaqVC89o1GpZf9pKgUvl7FciFVD3PmVIud7G7wmF
d+DbBEK38oUFw2g1Z/Fi0LsA7wU0dcSvmnPdtmxyazY+/oRYVQ5f7ONlWdAFy5zlbr46OupE8jqZ
bQf3uhY+pdH5HB+gITfxeU94Idiw0Vqquxw6f49SNbbH8V1W6zl+UwWtl9KCoHWNF5wxzl9IyX/G
TViKWFJWAbUDow7roGlsq+3BhtoCMShvS7AX0mYVlJI38ZY2BqGCNB9FpSyGu+/Kko5jyrpUF13r
dJkqN+DSiVRE5Gv2wMFSPJS0NcYrxgwJKhiV92/OIrWUI3e0TidjoDoq5qNJkFvIrsliKP44gg7S
38O6N7BCQKBAeGrZQ8BHVHxrrXPEiUCMvvUWWODlcS9/KJvsCVIqxUkPvObyv+dTVmSkZuExRLGM
JZwhJ7Z2vsigZmL0Jqqp0LkKf2AtQxuyHHvKJvMhbuWOGcf1PyWI7gHdswWzbOerA/aWerO6Ok+k
r/VoLbT7s42uSEBQ2VkTF8L6YHP7Z0Gb7KHAuNSmo1XqqlNIQrsyNCEtWmhr+9LX87PIb5k1H5WK
yHvp0Tleum4x80XKkz3StxZSzTDdUWoa5Ox71bdRzJ1WJU5oHS3fxcefA+W15c3FhP8ocBOJax1g
WXMex7lykNs5BdIuvpnA2+jiyHT6XZ6Cnx4IfDAM/ou8atm3hDlr9obd0CvFDaQi1MO5T/UF6XRl
+ktLJiIjHj/iJQdnNnjU0/Cdvntrcud/UN+KoBlkMS8UClgWOR1dSZplvoEXQt8EnaiU1BdihCUy
RvUlJttlgX1L/ZHwwsvigwSwB0kAbjnWj7h2cwAZYtGS0HErYq0LjiLQpkCWdjIgZwdgXqcC+5XE
xu6pksUckpdwLfIiCtkd1sUKnerJLl7skzTdXjtc0/A3IU8XLUM5m/MPQ+R0XRKcI9RTzpiMqCBO
HKa2uRZwmM/yYJiWCoczIios3QRNKI61yGWyczQOrkEH9jr/e5/xHd2WyxpPzmvOjWAdzTogCbsz
3DgJCFgMNtq+MwJaOaHvBM+GkQbNv+CwdxLV6Lw02R65nSA7jIuX1weSQ0KfX/FrVvjdAqLshF+r
TlE5R2+7MiVJ/lSaMZxwgZelNs04QRLhWug1XLxBPRX/3txEZBQiRUYvMrO/deZuqDTcW3bI8BoV
qTTr23olxFRuq4kUPqvswpvxFRH9xcobuzbzFKZeUWO/xMLav7hGfz4g9TfgLo+nXMoWBqVPu+TI
q+CkdDYsBQ3oiX1PVEiD9U1oyOj+kyaQSL9JJE4Lh9jDBu1j8DHK0bwTjjHtXtIDVI3BV6avYJnP
qduaEhx8DZlNEpWNw3qpif0exGuWLIaQO8z4/LmbpMJenf89nIchFNVVFxJHRFTGTKYB2qFahRBo
5hY2furEzI40sU9KxVeVad8u4J+5NZJl4XxieVY2wW/lPlXyQLNh1QLTd9abQ+cKx44mWL4X5uEb
EtiOCbBqZfqqsB51ENsASqWVCUy0Sgdr+DBd95bAY3wGG+jSQdCFk10r7nSKFMnJJOH2/DcEnRdC
UBX7sxbgfoKR7IcvxW1+/2ZWucM94IZm4CR3zjL1mngtsCyQb8Dtb0fC1L1gcUzOQ6gEI4xwU97y
2d2wTiKnM0bMcw/+wZy8Sa2hQeChzYlLtgCXX0M/rk6c+RJ/we7NwPenrpY7ul9MO1XYThfI5rNN
y9o6YRxSyz9OIFKoS1al+v5y1qAqno0cd6bTTaqgKOl/gb0t3m/OEa17IGGxpPCjX3TNP6qUNd1X
COalz5a4BOCl4VMWQtw1vkrs37Met74RxLdobkkmz5C2vyQHbBQmoR5YjjeKKe6wJoTxx1WNzp3d
y1yhByQJbYgPJAis7LuI+GClD6K+1s8dMUNbZR/U5of64NEWMazSpG1J3Huq3o6emr+vp3ukGMpw
ygKRoMtrnFJZX18WvWx/vc4TDyZ5RxbDpPAKASZkJp4+qg3ZWOXFWCgN4GzYPX4hlwjL6PK4E+5C
6sygI3Od7WJ2+fayLgo9DzVC9/bxkQz3OEMENM0FjwR7P9l4SaRFRSTNyn86tNlg6d73htH4XUit
ks5lRpshlKhuXWFOVnAzgMUxV8G/posC74Hsan7LlKqW8KRoqEbvottUwrl8MI5DVvwBvQiN6q/a
nAiE0DYP6ipypRlLFnthM+1X5+0oNPWzQA7bJh2qwj1TCq7YxJix7iaDiqoj1kITWCbUgSDPVYRE
iiiJfXeYwwhBe4EV4RkrRNLgsj6PRr+NZWLvbvlYCNXj7XVB4RfgOo0IvtoBoTffRyFcXM/Pb/nu
ixTeokL3iqJbj6GwtyOZgKWEK8811o8LasOzdFKU6ZnzQQhsG61eB+KrnGi8HWtXB1Da+AqK8rUP
S2Y5yhsKd1GC1JqebkQEw5XSV6qakXA7kbPXxzSnfKWZvBLRBAlS2/MAJrt7b3ePXbffu2XCr6AK
YodvS+5vzbSmau/eWicqUrEk5b1v24zuJ2k8472pVrSCssNqgl9u+7A9y48A/mSb1OCvMs5HMs8X
ScZFwShIzHqwGTWy9ZSD49S3KsxfhWxCODtJY2dNq/3ZMGWaUAzFywqiErVdxTT49xEI86sSQEmS
pmNeGid/vXKyhRVOvTgP8K8ZlkWImvQAjwJqspJVQ34ZBcjDL+LYqB6E8VLTGoQhsIh28HLuCoGj
iwDeX3u2aEjn2X0F3IFfpFDk4Tv+GG0bmWuLarbbBCcygf7d4bWvu5ZyK6Cpzh2HoPd1ZVODyZ0e
mJ2BDYLYyl2TFLMuB5gFyC2pITXqTv4fIabgmKzPKZwIIFVEzFo6oZ1+t/fL5uNepkDvi8Sh7LTl
7qN+oEJfpBm6ecjhhzGm30wyMx2814ubO5HQcVppxFhHDZvEHWbIWbfEwheCvQW0KCikA/sc8Am2
78jXIp+VHmPZACJN//9aCHqGudZ14pbEKeqyh2WhTUoybx+IU/M3wwVlRBvbtYWUd95Dup9rhQr+
QPi5yYnpEa9aCQWRVuWzQy42WpJXkL//ab/hbyVZaqXC9u2J227+xT0majDkD5btvFCCqNSv8Tpc
OHWrcBpvMj3NFQv8UAoamIH57HTD8IefLEiShF6af4NOmyda71vFmsAq6RMZQyWgGlEcd1r54or4
Srg6RZHWrkSxZ+f8rQFgxtOmQgEvJnRaMYfTOM9bjx//F7WQ+vvqx8Z5ybdttCTKxioMfXOFETAK
plJIGYy3Ca+xl24kRMiqxg58S3lw5ma2NngDtBUJlz3PX6vmNM0gvw2lT7u/RWV7VoaAGOS8kHZp
kHsbq3131jnmL/Y0Iw6KOs5utWOW6fVuuG5KeyACDPKEEDrA5wNIDB2yJItFuUbAg6x8czQxVmfi
zhV5mVuU8p6GxzIde3bDyZSCKr6/pdtOu3rhsMKskRpnFGG3XqkpRh7M+aXn24mQPuyUWvJJnlsD
YzeaUSopbGk4NqgKa4vFidEIEeQGVBaSb46hXq5p8KLTBO8P9xtQJDpauPeMAkJHWjJvPUOcWvDJ
H2n2JKFrrxbczuBbWddtOJUREaambvFPTmb//7/vIB8yBYJM+zGGag8cj3mHwBxGPrT1XincqEQA
uHS+CgXhdCLzIVTjwX6iOf6i9sfeczUBmnM9amLEywHDxD+IUS+ry7Qcr73VLJbEJ1f1gjwSzmP3
7FCaaVQ3kDdurypXARxuBecq0PLTFzYs576Hd29fAjQymepwt7A9wh0FPIthUf8i6OB0Yd585+sF
IgSADOjkr7oYMM+I7yA4cQdUT2TTK9Jya9VFgA2W2WEQ4jh8JQpnuUCYSZiqtYXXHR7v4X9aGhZN
OLXqDHoPb7qyCrQjO9vA9dWejvMc52eno1t+P/Nkdy99sGas827gB5aG2Fy7kU3de+9yuiPB+EE8
d5U5M9IbDQOd8Vue9IYSERJaih06KYbV/A9mxwhnaWtIMT5zFU4vG0B43PVHXwXf+DuX7zAjp0yQ
9Qs/HRa6+jb/5WMiZC0+iNVIDDT0RdffPud4KVIaW6jHw3UseXp0MNiexasbRN04RFsdKtyQ0LpP
KQz38W8NzBuvxI8KIFxoa7Nst7r4r2b1uxOvouFT5yKQgT4r6OugmdByI3PE1T5nrqNiw6Sq9u0X
7QqaqlcrejlX8PSoMe96NIaNL6I6P2JxylTG3cfmZdWHGW8z6PuJjqTjvrdA8Ub4GOC/6ZVeK6wr
qPPwJT3Sb19RAUrihhnhXS1lCEHuUwWm0KUq+MxNRqqXOQxxCHrVLGQkAX3CKKjcTjxGhC01XBB3
czzoN/zTmVnF2j4V7ndObnpyytoWJKMN5tDBr77plX+15iswtBH7lmJqXj4aauP5943IB4J3aiCg
s8pUPRf82FY2uUGFQtdZcJfGhKUb9DTJeCS4P+nJtOjL+URenwyAHAB9ab9PzpGj33c4knPCGj8W
Y2hvTH3kuukoAxkeTdaFqxf1z6UzgBwEdH013HCGeKvzXbd/5zqZpjgANwzRBPPIP/vP9wgUQjgn
oywDKKdVlJjKXYME/wzJD3OycEv1UHBZt/fmpK1l1j0JfD71xYYywp1ZzFcmGeeZQ9kGUd7kxPZ5
wbzSA7SZS8MVISVfZENW4y4pRJhKWkKzGmYEDnCRh6imLhf39n4Ma/nFltcYOp4nUyxhkAiUyPnn
aGqpvdjUwrlLTDIXJAVb912+7nSyZLhjrENUTDVxH1zeHxXmysSgxTkBPhQbiFMPeVSxPbDaL0NU
fx5nGUAnVjQpo7E4tvo6P3g77ZCEoaFiFyAJlaH6Hw4VpMU2+ncve2ou1xrugGdC+5qsK2rxAYQn
hhXGQaNtjHmS1AqBmlpEqUR/XdbWjEwoJImB0kcycn4ebqGZUAA6OUsn7SxUdX6KgaNOP3424Jln
McyvChiu90gcc6zwqfV2i5uSby7YkXr25MWLyBlRvgsFJ11HS0aCARlbkyuaMYywRB8MOZKOG3p8
Ec0qJ713I3fNedbaS7FiSeQ2cB7JjDN5wt0mgGcraF+aVza30Vbogw/XStNZT0PxKz32/EDVila2
oWi2OYk2iHlOeICfrnyps3NcF+oXxMlyxezte1Flf5CKp7RmAgxuvM3rChUj2gxT3dkwG7Zsr0Za
J8OIGNMjA95hQlnqXnaYpaYwOhdEXX+FlaOZ0mq8U4KdsKpnSsBJdrBAFn7vzFOfZkC26F31ZQIG
YJR9oLrWl0g/pTux8HFhZ31/icYflOOD83xeS+Ip21IsIwXGeH1uMqLMY3qbTWoC39P6gm0a/sXn
NGPHD6LOgq88LJ+sZkHNjhsY/G+fVZDgW2wn1C08pM8vB3Xaf3vN+7KdgSKhhrP2OEbSphmgXXPd
qqYqsdjsf0V4Ke1xjxlkHuF67xchtaU8d5dA69BS1CVvE6MC+6EPCUo1WQ2kTpFnsRh1qITDXTmN
NjuVA1mj+h3VQgTv4OzZHP96V+g13pzH+tBX6JwBg+aV9NU9PDM/jKJGQr5l8h52M9Uw4e/U4FUX
BCoEYoprt7wYRdt3JTouytLixXbVbJf5dYC6+0EkBTJjWAD5gH93W+VFmO2N6Xxlyz2rP68IxXWK
vjJnms9Fv0jvpuKe8GZ7BEO/J2VtJu6gzcLXn0jJafQ8+7puxMV3OHlzvrvA3ftVstfq1GouZgcy
wlzPazbzQyXSu67JVsOAdPEmQQzy6Ijeys5hrkqBsCaJse3o5HHcWPBhkHqsetQEGcl1PFqU9nhD
KuUTmKZAPbsy18V7PQIq6Kb4HjgNPXhsOLTpQ7ecHj4ViPAFJbkEhgDxTDbnU2t04SNWJqPtxrWl
DiiC8xvojrMAAeveZnMC9U5Bfbun+tRST7e2r/xa9+LB0Ekz6GTpn9HfrGhrogr6Z0Bj7RCuStUq
G5MICJyHgBXzaViRWbJ062hKMJsHHzrJaM2Km1diosYL5BKNtfiSipbXvKg3FG/EHdvcxxAzfv4E
v+qctLgwDQYqVVaM9T3qCAm+LI83Jt8nb9nGcciRdcpWgqfuXq37EzLjlnFN79tFGfeExACw5lut
0uHpTOdjgsIlww8/PSLNm1MEIP6VtkeAk2D0aMwXaRhy5LlHm40RtlC0Rd3r6e4jLgBR1r/bD4sh
sdTYTAOges8KljppWon18JDGdXX4W/olg9uvN0q+z/PNF0fxbPyui0fRnBJMqiSn/lH5wr/8EnJf
4XJZmfghb2+ViJRxA8AN1GezwUqeN1IbB+6auC5sBZ65hUgQQd5FzG0G++/QsbXX1HK/uFeyVBD2
6G87FN5zMWmwePk7PljtQG/yWP2jmZFILKr/igCIx2hAWnSimOg81JlGu6OyAeteCmgJdMmmKsbv
7bW1FT+JWGf5lmuvPQP7DEvuLV+pn9JijBKrlpG2gdCZSYdt+HNaFWOlSCIQokrg0bswr0CXecf3
W9a01cAWt0U2LIb1DXlhJ0DBsYvuhVue3kaS8HGzJgH5dLldpTem/oIaC9UG+yYremT3VzcCcnR5
SZp1DUnokwvGaKCjKj6+dkNbn+t/riPrJSBNrK3Qm2K7K8mXK4FWGP4ZvLxLCB25/zxhIFPKXg2y
BhLEqwY0SpfZG6EttYqDETNXfcGSKbabC4zC8irzsphvI0guxHrKk1jePxJewqux3vFHW9ZCQ3jf
FJalnjgU83MB6GYas02lgDuS+af7kfs1jhbp11tt/eXWfyTqkncqMVZ01QlMcx0asUBl3SxTlMM8
DB9WlEk2rW367wXWN04EQD+RJHn1lDdvtUmqaErmc0No/Ry70n32hee+1pNSPVM2ZKUWkHuZMwLw
Arentw4aTR3kPIaw4KlWBdWcimd7cogLlFmS/CALk/33oFGuls45UOR+w4oFdeU/CNsIuQG9Rnsy
G5n6wkEiB3pX+a6nR3YGjH342GJIGl44R8l3Ob/yVLlVX20MGu6H48yMqZxxO8UCUcIH8NFWxsZd
7YUgJ72hI6vWDMk2TR7lEVYoBWiXKN9WNxZLoA/D6UKgIt36O2YE9TH6AKyFrbtIAx6S/k25pgHN
0OFSTjcTeHt/tVP+8DQ+JOW20Wf8lHwgwM2/G6qTZEXb+qqdhpITMS83DFJQp8WjEBr2NoF8ZZCq
u43jky8gqNPMnlTJNleSqW09Jy3An0L3dDArc9CqKuSviyOwAd9I5vrhdb+UEHhKBwqTIK3/mnqk
SlJPXGmDZZFdjnouh2ou+TEUq3nTVqNrrsXXw+kAvkwrzgkYdOsbi6tIQtoo8irP33gwiFsoMpQB
vM0h70UG/+DtmAqf3U53DIG9nBM6pbdulKAhmLnuak/zXHuuKXswyH4Tqrbz1boXtCM4o+S2UAuF
GmzYfQ2/MENl6eJ/eBuTzgtwBtvgk9mDSvzQ+lPGbdCymkjMS5E7PVUqrOVU2DJxvVbcsEAueRuN
zGHsY1VCkY5ktpSvrzGZ26XuLd/maEdwv+bgiTqsVdNnGJC+60dStViLWxtkkYTIV5dExnyLppem
mUWuKliP3uk2fRu9CWVwrSWm9CFEh+MNlKCnLRkJcsp5az7CMpqB0oqFFJ+MgDhMXgrmfjzHtbYB
UtukYbCf91U4AgBskFNwHePd8CBVk8lMbkJYPP/yAFmN6T++T36iBKTVaYIi8ebpGo8sZd4PYijW
h7C/l7QOPNzwrTR8iEnx4pCPhoPhUaEsbvEezSYFbjJK5ecdfbTW/J0Mbg2Qg0c145t3gkOSBFpr
T2UHwk/gmHh4Vi9ARQbeQ6O/s/Y4W3I/n9Ud+4fHpDjxBgI0vNEpZt1Ib94csvCUCamDD/WbJrI7
CdGkO2bkXGN7hBgQ4WVj3/TVM8Fn0YO6jEzKZ2QPuGlkY3Sjq+b5LeQLSzlkWCTGUTo2MOXrZoNS
kXLM2/hWSbdsLDEYG8uIIH613PCV7em5lk5iwQ+Bjrr1u8eAkJAfGGwoapSbHLoGnWZnu1YqPVD5
8zzSyIbt4PbwSZJ+mGFE5oCNi+zdh+3t91TuGr97RzBpA4mDsgL9KRcbN/xWVAFxSKP5MhY42yRF
ARDY+7YGZRWrGGYlH+GgWLohtMeMSj6ngB0AJeVjgnlaka4ag0tViD+tCc8dtxlJjYzhhGkuvfoB
yn2aMIbKXKhlbqNifhgbPUe6tRQNaVKI3pHC2MnXro6Q1RixUyavsvjonzCBVjdcBicH56AR6rmZ
sSkqXsNcQaUMjR3MKktCCYHgqU+RU9XAY6EuHfhuJYZQZIbOqdoOOjE+ZmFxgAFkYmjfjANLH4gM
tMQ79xnflxRZ9dEwPVeumcCYjKbze+J/fxo7Haz+dbXwoBUeQh+r2tpBYR9YeWz/2mdrb+QEXH20
hzG8vom+50JSUbzFLdgOIQyVLJ0wlobPXsyWZICpPQRUfFtv19tqfqldrAw6xrp7snrTuzLZTC6A
uTQA4W0Dl2KaTJ0tWTmTKxOH8Fo43zVRhjwBgCGhrPManzItPI8nTqWneJ+/1wRDRq7DquJAJVaL
I0w9S+MKzgIhGKpZ+QuHxHqDqxAbfPjSdH7lXpn/ZgVVFP3xK1ORv0mrmiem61ddfqPF24bRRLSh
tUtGIYytpk8IDI+VS0Lgqfb+e06DiaGRtWyNHG3Bp1rgKNzLEz0wotgsrX201ZKxSeAio8EgaqN3
xN6S6xJlqM0lu7rq4uOAsZERATIwWyi5FWC97zUaRNlb64FukOPDz0hLE2H2oSKafLVfK5UUV38M
6cY9C3FSfdiXklsKxoHHXkXVrmZT5QDZj6CjAR65+kWg++mzJLDYUBszoBlXNrTO5mkx4oxKQ1ZW
OSWt69MCm3vbWr6PiVJxFyMppodlAjCjEIBzGjhPk0cy/hCRJotK7uaWR219iPsOp60/s75sXUwl
i5HgT80+Ainmsy7eXTRb8+qyFitNGM6TgCp5rMke8JzgdHYGk2GLo2E5USKoM6lBwFdVBstdJihc
3GE1i+gFDc4HpO25Jt2x+3SaicCk34wBjjnHkqyna7vdEOJCBiLkH3rlf+uqtZQysHEfDCMLG8ro
H7JgzkUG3V1Sx8etR4My07TAvW0FIl+XnAVIkqbRHXN3W+g27jeAv4mA9luu+kcFsKkdpZdYm/uY
lSDN3DFOQCiPx2DlXdo4+0zHW9s0Zvrn4LDujV1cngkmrS0B3Tyg1onTCk2syqzwD7aCM4PV7E8/
PGojASW7aP/sg72HCDx6y67uh+RRlmA6WpuyxxRv5PHwVZDfxl08ANfXUIhCDjsxQiW78BIJgWCU
i19J0v8AZ+q6fBkhFaAgTpv0mZJ0hQluLWQvPA6njE8p/Dz3RdhqYSBYQYQmyA7j8hkxbWgfAL38
h+pJ2C6It1AaDb49B+WTmjp/UnVdD5FFZf6RBh1WslKN90BImGYfEOmWlH/wVMT1xkBDnZ08TOGI
lVPCjsLgrlRiByKSJZwuvfDsIkWxsJdcDdtc9lPhYVVDbrfkr3p/D98eVXnktBOX+WghSfNV/mH2
sSiJPEwnJZKFiPTnem0e7JhrBmuvIVNxYxL2809JK7cxniXpbZ0NEhKeIWzr/QdXbNiB+1PM011C
2lDmAy3U7Lz8eJuGvT0ctW8uN4mljhPWZOt66/n/FN99mAW8U8KWHPIN+uAF955sVYGphHgnBmeG
/W00uuQgmlRmQxzuHuiL+3afdZvaDHJSTo/UqR/JncXAazX2P3oWZ3JFV2K+C9aHfFw7sNJTYC1Q
jhEy85qwGy/PNJEJJDcMdtQRcVwelRp/qcAemdrX5Kz+BG/i+d5DmWhN6LyDAd5a1xgIVQ0T9uue
TGLDz46bPStUxStFB76mIv5iK6Kugj9SzGSjb/oXgeZXaWfxqVT8L9gafD0Y/AGpiW8RjwGz7g8Q
R7hqegUja2OTGKVuvOZj7SLcGuwz5+BEhYRej+FPzMOee3+pwJ8aRe+adHibrrai9dn8aavwNIRi
IS4xZVOGXRwQcajVII0eXLkWfesWZNMiB/gREdiuV+Pnuj9H9Ek9EVrES+QT5KFnBcBBKKzIUwe/
r+Xas08MUwlqeTW0ULdKGLLpm0BgW7c1wGKt7b7of0Wqx5mrpyqUoVSvhwCBO7Vay6iEqO9t+eYS
nfFFSu2f6wH6eWHgSvBxWy3EXUxjGOzxgTZJ4P5Eyo+XceDqgjHa0dwtL3ERhycEtowGWtU2pGe7
EHEJoa/5X8DIDLkFq5e+uBy1KNhC0zD0QpuR1GHv25+J+WZa3k61JQjKFmQx5+yu6ZpyRIL/md5o
IDbhxnFMaF8D230GI8V8LkDo4hx+ftZn9htlYjwAYlAtyI7hrfr5zo8DhwXdmDrZdRPVMuOw4wCl
k7BfWyVQSqerkNInPB8BtvYcg1RGpxK544kdkkVsYu+BrXjp9ZqFx8dlej07SYk15SQ5IMP9e163
dEaOh1zc9eOvBLgp3ga9r5O/2VSiwK8BNm1qxiajfaomSge3GSnc9GWE/Jz18+x0ZJfgMFryNezZ
uUWjOyqxpel7iyB0nLRYtWIqOQ7hlMCWltBFmjclg6KnWe5XukuoyvfSN1ut8Te02h+iMpZdPGTn
qYJWCL2vZ28C+DCsNebNMcfei+BxKd3t62I80K/DaVhPej5Trpi/BwHfLVr6Ka+FzNtJIBBak6Od
E+G3+naznT+hmEvQE6CfZ8uum7MpaN8WbLIUQDK3cS5GyhCBEarlBMekGU7G2p+uSpM5KHJmy/Ez
vGo8ju4Mc6Ut/OHQxjq5M9L2xOtsgpNLc3+mOTkJqwce9Od2s0fiYjvmduqUZmREcFfND2/5lhtT
mATo90dtKdpGQmABeNmMQsh7FZbHaM3vOYrlyRSIUtTxXD6iQod4+FfCx6tC2QcstPQY2iWDAAeG
hBTs5FwexuTw0lO7U4OttxnTUQtWSlsupdvk1H+muYawWu1JdOpZ7h/g1dCVX7t00lWGjZ45/xay
IYd5clJHZuR0887XwPu0MA0yHMaXDwUuNADW+opJ3E1Z1YO57QENRxexBAIV8m6DKJUkXt6H3D35
iHg5CcI09HEhMomiZZ3aY+6pvKYbGfa+ROAO77OOd6jd+yi7kxBi+Cqd61AmZzUfK8senZBuaivB
SwSn84KsyuUOCt3roG0GcBAfOpk4y9eVN5nQFG0iiC/tia0E6cc3O8vX1pOsD+QTHQSU7O9X8aq0
6+g7AHjhGTOCGqXVVlDqzTU3/Vu7gIYFGGTTg6arZKB8MqHvr8hOYqVNOCN6ZzgtsrhIl8Wnfib2
wSDbLtUuqbW4AL4OWK9OlUOLESXCiHhesstVEIBIbNSV76WObTY9JT96TV7yVFFwUfd25Q+WIVbL
bD2bJT3iKJ8UCvh1wLQEJzWMx00P1WyNCC/L724iJkPX6uLDEgjFHMuMToUJSYAgDzaCTzq2GOa2
iJGmpTvzblp08R+eDuN19OsB+EBJ5+TTtIdljRKsW2nuNkMA3ZtRrkHl/HTNv9W/VsG1zLuSkyFg
8vTZqhi660vXqeyU6cZ0vl47vYaKRQNu6iSCS/cQNLh2nZ3U2XA1Lr6Ngm8xVjFRlKqOPA2/W8mZ
fk700gRl4c+NuYJMqG+QJOdjL3fzmg8r9UJlVwSb0frhSneFAQtGl38rIalmlfWQ+tcqKjEgOaq0
VoxwYMiDyi+KPZlUwIhUaIOhK8QVAOcdtECKBBGUwUj5jxWzt70X+l/v+E4G75vtBbeswvdp5UPm
UijUDbSURLGvg0XXW0dz40oRet4TvYMoWxvFP8Nbww9HP33BDJ5zrTLeYd+RY5Tyu/vrTdEHGCzi
IPVTlfT9v8E8GZxbYEboYTkljq1ayCFn7ftlhZDKUahl+X4R4fYyDx1IDksAUkZ8DEEFIyZzTNn8
dp3tK2YAe8zJ8zMpj7Il/BmqrLd3vWmD0WS5iA4rRLjvryCRBIw3UU90UzCFnfPRlhviwdiPEgd2
P3XJ2H5z9tbRREUXH8M6/Rpv5Fe+eXn52YDCDJHRxHPvyf9B0rzgnLrBZteH1dU0wrGvDMzgjZdv
Pe9tm9BGpni+vvQYt+A1WzQ2T/YP50DFtosJ73cjYa1dq8UdotJR95STxBfcCwo6vxdtk8UI4nfr
A3tjCCYc1nzGKik2hsLrcBdX17jZNCoQU5BZW/JNOC6lNOcXQD2nitNlgwKEVwxWXehP5P7I2GbU
8cdivw+7qEnGCfHeGZUNOUYYsHAgdLG2j1bcVYjPcjTngvYpJK8PnGffwPObw8MsLGlfZBIa1fm3
u1nZrJNTY8G8RkeItX8IbWP5e+XnXeEtQA5MjZJSar0K9uhf6eQGiVK80OxU//yy4VtUhTDn9bo3
lZ0CQW4wJ9LTDZ+n4+rNGnj4gsRiimJvZ8RHfyXVAdwhl+meV86ZvqaHDukihYt7+XI6LVH8f/7S
fkvpZMUfPviAWUi6eXayx6Xbnc5WZhMknjyTdfnjSCZTG8QDXCbOrqcUXqNkc3TetNVFT8u0T6oz
br5ZVlfsO+Dh1YQeEzx3lsp2NV13DaUCv/MliIVVYB+kEQx0eQIqrLCgT4wmQdNlH6mqeZgaTP6i
1+HcS5g2JluHLjRN8cn6oRnG3hcjjKOuMqgpuXGsEAHymm4XRiW5Ew7p1NcgWQfZ8hQRNEAKZFI5
yb8LXLC/QEr5v6dyH248fqB4cgE2fDGC0dU2jc9fEwp5REKQG6ycI7WNLq4KcxVxQg/Mz0c/nesW
xBi4llLxBqBXODB2euzhFb5evzrVA80iLAX3dLRAkKqESwM1zB3QBPoGRhaXlNQeEMOrt6kBKIIl
oIOYJWlp90SGoY2DZPpvXt4nDtv/cYo2343bHtoNFlwChTanVH2l08z+GdR8IKGXhJTQMrst0sGi
dZEJS2XPIqfZGax6DUjNki3Ba9rJ8qxk8pJG/8N/Ap4D8poVuENl3HrzUayRFrZO5hLWPM/fD7+8
WTmJ8ouc76uCHgy20Il2f049mMDZVMrBT/5XRWfPHbgZi5cVQ77ef6eCiF1v24cqTn4WQgR2xMMM
EoPT7TSuERJ6WHrmvOU6N/MkUrH/xc0BqzobMItOy8nexcS+6qtBuMtVrbgq4UFqVNWT+2d+bCdK
L++sp5mnpaRCnufHVeUom6kBTOfpSPw6TvoBaA1cCPsvQpRYUfoknmmKG3yMwNN4mKYNI92RgCHm
vmw/4T79d6ZHxVipdVMR1bepfmJmKU8VZoOGbBLxuL4Q+5WoGds7DjHzaHRa/Jf1mFlUyWWVcHDr
QmMC0pfEz6FCBPskXPomqSpYEJNUEctu9j0BWLxSxcpvrwMm6WUxs9lQR4F8K5Qjsz81sGojGmH0
V9o7MBaOjBoQFOfgw9C4RpDENp0jvd2TMUN5fReWIvF+huiHpBgXQxFsgF5unLnIG2iyYT3HOFsS
dL4AvcVsvINlg62fXBEHDomVGSWytW9G4IdEn0SLhL67EfnwD1TaXKY0X0Gv2Nvh0P/VBLRMY9J5
x0o8o/B4yXy/peQ6ZuAy/LNC+H9ZwzzxQAsvFdEtj1nyYpi6ekjYra7VzrQzYvwtniq9qZKAZnQx
Z/6SW1gI3Dfu2n25MLhttBJQEPjfC85BaLLj5Y15Z6yhBgF9IctHAUVkvBm6qCshJIyjx4N0Ei5V
NRYzaWISn9RfTK1/S9uFYne9I70bGvgYMpYyIvznwssa3t97toApK0uYyRjc8VItz21beoy8exsJ
6vxwqPtuE/b0wqRxrnTdsHY44rz95jaq+zH2H7JcAHNMD/JqwOIdW9JGl5vahMDhZhPnkqYIUVDe
IFGDuT6z1nl2bmHsnlQhET4/nuKuCF7J6bmVN9mnVH8KVYGltYqvNZeAdtKFqDGao9pRAsLloEj7
+OWl/lU4jr4mPzEPvI4eBUcMAI1rcNkdUyNU6y4XJ/reIp+zkvIiSZIk5e4BKr+YNZ7HmBK/2uD/
4V1n7qr/tVA8ZE1scbcb9J5qjcMlAYuJifRAeuLLUgSJM4qeZc6Mz9PMOkh560g8OX931AjZg1tJ
mlnrX3/FOTvYz+csJO5wC0pu5gzjwOl/PRdcLoN61IhNm8/stdlUC1lzPT0TId9y6EpHiI87CE5s
zZbx6jLWLfGArAJHDkfRbJay3J0iuiWhzwhdXDX8vNpGoHwy/ez+PkDI/nrG7Z0eELZiZNs2OwO9
3hDwZ3kOqMV87OGJnn2SPxOBUGJrJdd6F5DaRB6VEiXdu1i4cQV+iTmsIZc7LsUmJcyRvk2BQoND
60WTWvyWzFNqiFzqA1LmveXt0uoAXi2QeDg9R7rwmfc4IWq2qQH50fGOXZ3Neku4P51KP8cxObsC
ghumXeaBkbfKE+j9bEQ0PJREiHYlKAhOOYxNOmrEveVeqde3kQDCkl4b9l0gZ5jCs3vTBIXu9ZK/
P0S+Qo8EpOooJ2R2wmptiNM9E/ysAP518CMIXwMFPTvqBwUeqiC6SBGMIQXWvwzqL65MxM/phJvH
c1EqDm0OgIVQm4lQty2p5Gb9Sul7T27VkID8xFGs/1mWS0TbI5TdVz48CBOpfbMhVcvtdgEtcIgg
RYQehXQAskLWf6l53hdDEgJ68kZxiCoU67tJdgxEeW8RRemAclY5NJgSw1ArB1zA4bWMxb2EccBg
q3a3ZFEnjiakTWEo9RMGSzHsUbR2TuiQ7jtZGJZ2i7rRWaAc93r77ug3Mf02dgmyyxi1x2BUTFM9
lx8/Jaf0a7Q3/Qc98NYrn5xhuYXmmrSmgIdFhRZMIvvLsrxZqCg/A+ctNEJNqtkgNSQ3Ec0dxaXx
w7hJLtIluzQveamjAUwAeGRM/5UUH7/iZtgYvY/3gLKFgB2ZfQrrkUYQa3MeBZwBvYZmlXK4C1kb
rE3L4t0lVNH2gCNaL0q5zPJTckjcr9EuGn/647CZ+5Q28GFCefWtmyTCneDqywkUooViHCvFuaps
t+jo8iUll4ycbzeikV3Alh2GGQ4Q73o0thX+JfCdDDpiRKPQEwI861FXV6P+Ax5aURoSLNyKVUaQ
Mz9iMaQERLFo8kUi9C/qt1WIlGi1rPo6qtYGWOjYZ2V7HXa1BpUtHd9oHe9zLQfoOJeqjjpYTMPJ
ctEJSzLlOeXmdkQtVEnNsGo/YwZ2Ev596IUK5Q/zBFPZ85SnL2gfzsocAWw/Y+/Ku2O6LblNb5Zr
9ugzySy9HatWUhhCT9UPI3YNIu7u83N3qAvBkfLWcrYdzVmoUN/UY9e2pA5wQns/diQ+RdRtvArt
x6e4X/0kKKGIj91/0Y5YJQHj6wk9MXffji4BMCcSxV9K3mKKKEZud4JDrdmWKIdwdQjENXgf/wyW
0ep8Y03tHUA/b2HpTEorswp7XMEkv2na/AzonP9znDzA7FNI9KUAvDMfqEx2tr0FuLt543NkHHzl
/PnOMTfaZdUFvNNS8ioyXM2LEw2E9UHAz5LiSq3ZePEKohv9GZt67M2JHRuB1mo6peK282qpnJtv
R0FSdc56zfJz9WtFwLGC54WYEev8oJQf221/OC1a4A9/mESL5NjstIkWzllk4qV56HMokDbt9Rat
PgpexFWeFlV1kg9qdM2J6cD9ZTRjmquMnhvJPTbpjo8Zd09PrfbskN3Sr5aoWm/WLPinjqhnqVdd
oKwBisP7deiuEwRCZCdQFEPaYF+24TKdh3B+oNTjJk/AcBLagx5gVV1hTiWolS1fBng91CYb6Ptg
rpprNQfeS7+8COfaxnGcFMZ2YfIvp4qoh2uObyPyBHqeptcT0YvvJhvWy4ITsw8CWhGRN9dUTI3b
kllguotI033KLvGd/XJ1b8eaC36wHPalJjIE/mRNSCtjp+2zDoBam2nfjNERx/BgQzzX+yW3X12i
mjdoQrEd+e9BU/CIW8ym/PPgD90ayhdrgKZ8RKqUQIR00OjlFb/aOuhTzije6BAlTm7/2d92nRIa
t97IBb6AS4XTeZnMjvJBp65N95QNMGUDToNh99q2gVKzsItRiwmqOTAV76r6t4v8fE4qJdiDWplN
SRVF3L4AjlFUiPd+xcXz9wvSt30pRr/LhlDJ91XeoupTh3mcnBcSxkWfcIhsb+xFYbqiqS4YsO28
tVYmkZvRgtmuGDKCXFC+w2tbcpRDtqxA0HH/F2f8Y2CtoAg3URV48uQ74dStF5KJ/9m+Ua/9vCfO
ZhRjri8may0TfM7ySgRlbFpmr1M8+VXyRh2stJtscV4l4Pez5NbsJaNWybH/eJmcTO41z/mMYAoN
HP9Ytv0elsYFd+UZH5zb0CyaszRC/cxhghiHNMYeeEzu8GTYGdqACM2uJ9TmfSZMePPJkdPVaY9e
PYBeNdY6JN4/Q6mXh3VJlDgep4hs443m7WxfIdkPgTjU2SPo//ywsQFnAI8Qy6rNre/+Wx0zhyQO
+4BtJxK7IJyTqVgMcyEsac0bM7RlP+c+Ety06uOGUab8jFdOBYj0WCrZCVQ58AupHcYUlbDdj7j/
hQDNKJwuuK+cJarfBSbXxNzGR9Hx91+a/Cmj09vm9ihMAuQyKPfVOZUbNs+FchHG6A+gm1bfVwfR
ZAMEsiTFL5lo7an/HYXJIpQwWydS4jeZLX8un6SWSlydYc1sondTro6VQ26QxUB+V5Lz2zFer32x
YBeGzjkdu4kbE22PkM402j/Rr/ElyItRGgmJFLUe1Qst3LhkIVzsXvkWpw5pPpxWcLaqx/EF8cIT
aWhpC1pz21/sohyxqGLVTNsdAvNTRve8li/bIWwrpU+oX9ZxT/3CIPSit58eQT9pDZe/WaLFHcHb
g+8cqwriiEi5i1b677Yy9LyFxV3OAmvW2qfMcYoEMHRuEQs99bySR8xevrFDtibwNZD2qehxv1RH
5NOjKmnr9vJYfZU8skfjBwjMm/A0kCL4aGJNiIfdi3YfGYtXVQBaROxKCTkPF/PtR7CAcdsRx2cy
D/WR28G1XQX61gqT5yTHNBF/iXKvx0QNKJxfUxGthCH9RTJqCcr0ZoZw26LktCqlWQa3dVbSMy6n
Vgt0DDS+NPBouPiqEcHeeg30YH3PczyFi/pgeUpCpePl2EYZYbDJyfQz3nIoZ8KIU0wLM0IdS1yZ
IqSTMHM9jd7Efety9HGykyxc+VXJh6PIay37x/hRxWOpV89NxrdNpFoKTyFd5fe48oS0CymGdUXp
9J6MDfY/d6zwie8M2cGA3EUOcmupOreNc9PTNvjfNc+RvdmbFISNyc77Gg8NQfIFfwjDzqD8idLf
5Bm7STRGex/vMbuVuiRCEA2c0FDACUHD0xYMJoSxug/oeGtGa0hAj9V4EcIuwpY9HrLulkpDgnaJ
8tDPSdmLcOZNXoSvH8xtL2C29xF+1FgMMpnhC2sXSzPwt8mF6noqDwuT83VIZDrsO/SG7drgAHBU
oWeFjgDjwg3UzWyVPVYb5GZH7iVIyJ6/FF++y7LQ4B2IVNrrUwnZGr2M0yOSoCETG7nTn5M9LAj8
TfqR9b2t4kTv9I+6vcgY/A5kdFOUk+4PdOsf4LGZBnfaeE8x0sRZOrR0EHTTwTRa+g9Syem4Ind2
PaVcsjnupo4PZ2wy4wscQ6U9nZVIq8DStLwy6nvebuYngqgQCa7vxea6D+XgOcAVkQRUwq1IiLvY
ZUzd2knx803MdxL3EJZXD6UKJZDkljb8MkC5MiyWp9lE0khLBg8GpoMSJpVTIZkUmOdjOF3hv034
WYmu4bPAfEFW29OEAiJhkNeVLOzrGefTaPPIfDXfnMtFlbmPTMOBcRPIqIKPLPQ2maGG9HuQu+18
P/miQkXpSFg81gJZ3EnpGQMWwta8KVr+x/HlpjMNEsuEcSLd4rycRE1D9wZTe8keyMCcV0TEIJW/
2Bhvt9hkRGDoDKsA9wl/W3LbbrtY0ueljtAXsdehivLlSGlTVWVcNahDxOncNJwOZbnoKmZA0nEh
nhxRf5OHEsIqSnR90BwDcnwrhoKkMvvIzPzMWXt9vK465POwTcW+sHXBOKyjw0GtxxRrFjFZ0YeV
C2jyxnCqGAfJDH+eq+qBx1RGOIFdIg1GSFeSDZIVgwR7lpJ9knu2VWva/Ega6uasn/GgPNIciXMn
JYLXqy1I6H6w30ildq2sLamBTh/lUnFc5nKlvslP/q3h4HSHzPrngTNP9RRs+rK9O6gJkiWDs5CB
bes1be1U9sphwLmoRg9kyWkdM9NpJ4F4hI1YRZtnTle2nhyOk6783n5dAmUhMgtcilw73dnb/0AR
RPThEKR3JZm8L6+HmFJjWOcjnI1HwkeINJ/yxEHmwhGMpkw6CemMHYLbyCKLRLQ8zX0ZV+Tx0tS2
ELMEHHf5a6gco7Am6I/e05G2MK6cu4Pb8dP755/R5thwcmyzigf52xiNlI6bu9qSPW48R6nVPJDg
3V2Mcmok0zvdfvvVuia3xiDULUDdLjAk3rA78OwJ4+5ch9ysuDFLnQykcnTZG2uGxMnzjCYOcsij
JUBabPO91tkax+tbTnG7q3VDCX3bWZpJ98yRkFDxWxTeT5dspL8ywsq7bezyv1xgkFE6IM3UdChz
9tLa9SkU7Qhl9k4etHPx0LkVvvuv8DU+eTuSkahq01A1cY36Laq6UkS+nMJRxurWSKOagHsEx19D
Mq79a4TBN3q6hgUpDVjFTOPDx/uqzPPdJE8kYb1rT4ML9EdZydmk3X8QbTX12uL/rCVyJSqQtrlx
aGdTKqzyVd8ZSDB1Lu4kTfJW+oJuTDqmI3+HgYsq/EsA3fxjOU+zHwTCUGkkY99GctXjRpzoBcCS
N/8tLbvmcfO9/hG5F90uOq7qogw/oA9Ioe6M8/sSzpWgVLP3qKI2zzJVvUn823mpDjK5p8qKD5/e
YeuAid7ZLMVnVyLYxbfqruQHwxHFGo9GxZChNlkdTciRHEVHKdRy7ufcHU5T/09T/MMW6mU/5wxr
5kTSAyDIxoSIcAQbFATKDU6nwxWTfhK6fgym4icpXBXkUr8vrH4Bb6fQADnnKxCokRCuSVLS2ZCd
28CEtm+0b/Kq/nCluf5ylU3UkzdIBxwwinWSc1yEARldKQ+wSCqeEYXCy/tUG9dVgjUdmSTfxLi5
U9Nipi8Rj4o/4bhWydT7azNSiIaU3f1UYKQv+jHaAj4XAm9T3h/beR+dYuk/1E1IBFsjzdcYqee2
i+8+A0S640U1vA90IfaW4qoY+e1s+JDDvL8uOv42XNaaYU+I20pgZW4/GIWcLTpyxS1pOZUJXrDg
UTsdAl7+vpQ74Is1cuFAEqwCqChBzsd2gSkpOGC98wK7oon3NqE2Xaq/yGH17/2bzOheCyQwzlnn
red5ZXlN3C9gPQiFOrcpZsG+NUf5+mtKy0kAkG6UR2AbVb3mB8d7eUdIe5iQEt4xNlnM+JtV2m71
87Lm2yIG98sFCAYy9B+0GHuLQ8XOSLJE/rP/U3bZ75IioQc4EHW52qH2IAmO6m1sHDQSNN0b1XHv
jSJRw+dlyKINhDA2lHepTN6J+vyqNNBEgDajbgpsRD/KRf6KSGVw+cv4QeBcyHyCWOqPP/7+b91g
bUGq4iMH8gYncZCV/CbeiRJMH+UcwB+DHO2NOWXwalq8KGjEaXZu5U8zkNcsjUPuZqGKfxmVljJW
2pkAviEeLqtbPhXxZS0i7Np2LOX7VS/rod381NyOP8xDh+ZdLqeY1qxOVI1CXmmhIVzMy30gvB0r
q8QLruLvhJNMt7kLGam16ZbEX//YrFl2cNp2O5/lbhXGtosCjQ9/T9yH6pqdoHoaSbrVGK21FYdV
c9GFYHYxKigz3uFGw4pbo0df0Z3TD3pkk9Xcklm1pNYCd3qG6Ji4/Ou0MvkFS5dAsmFr3haAyhm7
Rj8zucYL5cH3QBCKa/o967+QJOL+PV0PGm+MLYL0VUM78ElSsxOwYvnOIkvRNtlq31LZxEJsy0aC
+oXlhUSVLYqy/P6c/WVsX1vh9ymqRKF5yT+BWz63RuuGss1iCWt7Dwf9dsVOI36XAm0emIgXwCAH
/wyvGoNeAOvpXFFT5hRme24BotNQAhR/xesv4KYfCU9lqlD9WHA5+GT6G3TqjQfvvjZ6ZGv3/Dxo
3MWvKHd0zxDOZVKj+S9NSUYU+ABIv0hWJUGdfA1NBuG4lkSNt26xiZHTvx5dX7qvWToiBX6RYL6w
+osZV8sGqcQJRR5Ds9YJfykc57Hg/8v9cbw3z1upAJPP77U38JvEzK3OLCK5c6co+SqSXgMUWpLd
VZSJmFsV+apeaUwSf5NYGHica6fzJV0pnwHznNcA6S6yMZd+i8afZtKWj3IavEZxf4Kbp2COBU/M
aqhdJDgXOeHXW8wN7VZMD2o+7fbP0SrNslJngsUUdKpdIccwS1Y0SDHXtgtgvPPnfEI62C1fLTJI
3/EIGsx6HZrMiGnH/F4vYwMk6xjN2BCPFouAlIp5meIon7TwNvDqJC8yzeVja2CbumLzDcL+dvtR
cb/oAXr8E1/qswqKHyJu0O2zF/bhSEKnEZyvdkq4LBzaAh13OqR5lXQGumIbV8+sXtP2mW4R7nw+
xvdiVe2B1cKUqiKbxlGFzBkl0lX/NTzV2KsfaGxEvgCJ8VQfOIacPpBBNGa74Rgjby79bY0cZWq4
waEyhEYqHIbjIRSFSuoy3M5ZLNQIyitlPXExkn8plRcTQYfkpY47k8mestlKwmvN8rl60ZhzGgNw
igBZJBIm7n9VcERzcHhJh82140Nfq5tXJPE5x/ZILU0WS5whW+ZcGBtvMLfInIdoFXQF58wP9Jmr
NFGhalJ1//4R7Kba2W8H3n5cn3Iqj4BECZvOD4EQOMic2nc3amgOgK6jscvQq/8nKQkfNCC+5qsT
CNUCkmFXu2SBXp/vElrX/hJWPmo1TpiDjOI4laFAQ1lV6px5laacl8mOJOaWlwDxRoEC6DLkVV+/
RaWmgA5LT53aoKeXqtjRWMSPmpnGPDYM7Gnbv9DRy6BFSoiddlVrimki3UBwDCTuXQxiMPBG8VtA
d7TnfyTEM3hBKVU8cHqpLYrgyJ+nU3Eu8y/Zqx1A93gvA0GFi+8NRkyVNN37uge2adYdgZ/+qcax
QABZ6bV5jJz7vIVGmzx8MX/uTzR7n5jre+Jn4ihOJK8bXrqQ4GSMZWkBwbNZLmyMlW6yOejSPg55
oQlva9c1LnNqY/jp92zppToJQ+N4qrMvHljqP4OKhySUBbdC2CRn0lCCKGvQ7eGWtm8sd3ijeXTy
5suIsqEXECWWLZYOSL74Sk2bVrCzYnBvTojMYrMEzUwRhCCjYvxH8dZkopg/w/wWsqueuARZXpnV
ZYIR6NLU3APUqbOiSGNvvemaRbbbEi7SfQIy80ffpsvMd20GEtABJgbHUfu6ps+hVAoy2L1OEaPy
W+PFjZJHA5TwWafB5iYkLoEZXaCAHS6l7tDonT4Z1Z7FFalZzJV8oRFQHZsTUsW0ymKsPO/BJLoh
IiEg2pQLECG6dJrT30W+L8UHsIQJHLXetZ3JkTmrU5m+pMwuD0ho/D7Tn59gw8SXujZRbNXK+3F+
T3K70EogzN6U1anKBdD26LmArS3sgKb+rGVX3LQqt6aWsePsnYKn+mBAaRSsUX0EVv4Yx7WDM1hV
9a07hoavpShQKiw1rKo2IWPwdJq9GjimoP+xI71EmxB/8JJMsTsUFRSBQo85AQT9ebsiaG2J18IH
2h7Jz8IkRZ4Dh2mpBs8EeJE8ZuNEe1r3zGyrdvV/K9s0LEX01cAjUdisOXYYs355Td1wRnrBkoqj
mawZgnZgZWc5jJg4Jy3tF5XHognHz1vJEFIxqfMS9FzMNoQ1u2ql3dpTpA8C0i5PDBdH06ksu/BX
mcA33Nq2iB7P7dCbD/WiE/mEbeVIDKmdM1PcqhjMSnCLX8HmvSuyK7d/ey4UFyrMnh/SbMFxpKY2
RGGkG/FXdC1VlkoAonF/MRzxQbIbqlolVwt8HH8+7ha1feCskDkR3XSZRZjG8MUujlAX07jjI0fe
W2Sdq0GolzzeMgFpxmbDQZzLBa2Qa9EbnTlhAbxfMZBSxz8e/xCm5TWaNsAL//aaYJCquRSvR9TI
NAEIqPgJwc9ziFeS8D+HO+bRaUjvG3BIMPZ1Ua3LiSLnEz0dNDkZ2ypjmF+nPBXe/5uPbU2Z9JEu
vmV3Wd0+ujjfxZYUm4RNhTeuOhFjv+POcinFOxXHdu5v1Zf4BIqEiAyJEAaE3Ky1KlmRhUBjGaLL
shFh2djhU+36lYzo4OjypvL4C8iKFZTPEde9Z0CFOt7Dpes9Ca5trPSDwcAmVLa11L43c7jlf2NM
Ofq6ikaGjt2xsjWOlNNVr5gjXgSKbOLlT3pk1wvp3fbOH4HUJlr75Q0vdP0cXdGSAWL3wUZt2CAW
VxU1gqzcoMQ03gzz9yyy14IJloGjWsK7KmaroD4kbz6Nqr1zRR72IpeYJiaHa+IEy2AoKz3AwwVX
IPNXfwesNGiGF6gnVfUXJ4oFmwka0NTt/kPinbWMZJEFJWg4/phHQ5QfygqVrRzGMC3dnYZfAHKn
aPnyyzhTg0WRw4iArPUv6YWSZh5iZpmzFfUId53BAEnIzqyaTe0mMfyf48RFQJwzjDFObYl9UTLT
OBhCDHmFd36O1klYz0lIScLlm3/EDFznpEnJeYy4T3KBicUUnht6jSooUGNqo+Q1zlV9jE679bZM
XOPnpyFMFFYVYHWyZOmnqB/9j8FjfvgnNg1jbPxlR8qntQTpHH1bmcVHrf9r8edywf5dWrr1LkaG
tPf5yxoF3n9Amey4+SFMUVvg7v9YWDQyQslkQIXQfOSZCw9HoPNl6UjVszvuU7ZdtxRh6qPC20F9
WkdUl2itfAqvSSRrtXsgdw1pMIY/c/Rb3DP5TMrWQkheHIi60oMaWXsoJ9ku6wbjOmOAgQ2n3f7p
PyaIXthdvSvZeUZPJqudLdXZ5cJAtTQlwOM2w6Wljj7SoXWlh/sIY3kmvsyUVy2ulmCzxKP0M8I0
nSf5qWK1sdItSNzdMBJr6Gln6fcaTMZwE8tiL1lYRjM99NOUXJCit/t6I7AHcIJP5+MSGxv6rgTJ
AXbnQwiDL3+nAokB88gkODn5zP8tryyk8HbMHJYcg4+WQm+AhldUEkHV7qG5lQkvf56zETM491LM
pkQhLUqHUAEFATkcXKwmeybYV0Xh8TVlTZdTDwbKZnliwR3fdJWu8MrXz7tHEjgLhZYaaci6a8p4
OYaQL20/m9uIxSeM41W4E3VA0qeM1HcrEREnXED8/vS2/yKUsdCigHFPbWpEwoaagAl6dPMum2nU
t3c1djW3/hrUGvf7GSZQ9gE/MeazBY4fzXcqJH2FTvYyt6Ultc2otT5wonZvMslaWqJUwxvWsajl
3CcIFVPh/20OAZZlhLncUps8Jse6moD4MXyu6sx6gQkGo5THg4VFab1g+ny6/7frfXwjdnz1XARl
cK2wvbscqNATxFb5DttXSsQ8VhcE0J9GaAAnVRqt5kgR1y2waYNVD6gQt2WiWaQ4Jgo4ycIEeCrF
CnuYWkHizqVGMZu+a//8v/4kXOk7ugzmBqJz6iYba61HfayLCF0W/A6BkP72ThFkWdO7xHrz8NwA
bP/+hvLHVXJEvSUq6J4Mmg3SGUKeJ2ejju6i89Pp7xOTk6LYT2UBhMeil5bEvNNnK6aXIWoqjoOT
UJWluBDxlrWTHTlPdnEOf1E32kcGHzeIzuEFtXOGW9iMUB4HfhOwl7KJsmtuCOEY98CKP6Fa1uYO
4LktloGyX9tiSeQp/qF3/LkO+Dyk4xpy/YxHKs73QtBEZyyhVZyGA0uw1QYabcYf4SIlU8XpMU1c
rbUXTIPoaxe2wj2bP2BDna3lYEUha0QIhcFkTmFoyVniKFqH1LyZAyixBurjNoOgke9qx7HmWAIE
MEafobhNhNLnnsERsolBJ1UFpvZNvONLiCpF/C8CycNzHTw9YY3piX+HaC8PVNhv3iSUR6Tc0uRB
YuVcpF0WJ1ePGa2xlcoo12GqXR+taxokugIAVJH+7Dy6uyCQgrxtehS53zZJFLPZAdEPQPWvP9vC
N9QWEYNQg3qVObc8xddncK4GCQHP2xTvxfaf8VcaC0wuY9Wc0s8uX7vPPqkZ/Jf+OZ82oZ4IQl0j
x67iecnKpfvxA9qMaq+wUHlLEYW3IrnxWBUxYIzvIznCEDGtBJvF1kGiY6hyzF2uxHhilmqBmMmO
QSeWJ88y5vR9mURmTGV+GKOHHpUBwJwg7oXG3Un2p6EubRZWPya2zFJUjEJaJpy6TW84J9zx/NJO
zWiYq9riIJhMWnwp4AdzyKdwPOg+Ryctrlo090mVTu3f/3SQO0FUQ/xgJ9emZhdfWBUcjP1q5MDB
knimd2DkM3XWzgCIW6Nn92vHq/wLboox828Rhe05OpThjekROLz+XAWIST950adCgq6Fxy1Yf27X
kzvjvD+wSgfToJ1JZ5E5CACfJNkgcxKU0cHZdDCz7UQ1tsbJo5YrDPs/kVZeWhUigzFI+z3f8phm
KGD2POnmOT3ySvH1XYlrSdoEDzIepMGcND5O8u4FzkTyvCJydRRLWz3UyT46KmvEfkQ9zqJs/2/Z
bEMXmcFHHjRVjcxq86QvQIiVp1QaDziHgmwbOFInLonlRYXhyAw+DvkrmReqfDXofN027xnbaeuT
VuXgZSDkNRYQZZleJoHzMK1h0/G0YFGFg2fn5gy0CbCLwauDujfkbwJ+7lL0NcJtSykFse8KxNMD
sZuY1b0WhGXxVZHQAXXG4/WwUNM3p5GSrr6RfPuRnj4GeHANIlPceHPEI/H8JGCEUHC3LhCIVM7e
joegqFgtyiPrif0sShbc5TpyRjFjBsTmwhsYVc/xaZsZkewQ/wJ6kiKrAWqx9UU0X2rYFY4gdIXr
3RtnunkENPhuVRzOKLQa9oNc8lncfoFhVYsPYIRj/TwYVK1i3AeV9jaJnv8RWYnkHvhYAxvC/TOL
6ArS14+LmDUy4I95STXSlvIv3mHt5WiT+7hIW0da1ukg8EoEAuXXj+nTKbp7ty8VqT9l7eiEjDAL
kNP6rpmV8cUqWhMlHCL4pI3fgMu6uFbTD9sBeyiP9FfeDSOi+4wdkimHVEKYGS9FL69gaosapfKW
vfqh0HI+obpxSL9ph4WNhQCB9RJzjiwds+Bspy79tmgeel0F++eneaxZr5jm5e2Ca1PNOpUz8U98
agWS+gpvg1nBS6EWglkVMtsTSO8a/lanFH/vjEOpDbLY4fW4UX1gBSCvFW4bFyMmEz4aJhlhMPPj
5e2ODpoJoHzUZ9hFv0cKX5ULyl8rAvmqQo1qnSAEl+xeL+qxLdxXPJ39U5XmBhw19cktRd6OGF9e
4/o9hh9bxcGD5z4IaQGj1J7CIzf69A+vQZF4wF9Jr/9nkSTPXew+yyG0gEFjlsanNFCotUBRLbS9
FEn17nLSaqx365W+EAimBpdzv1AJbY0yc53AXE5B1wOjcRQbbHfO7uZwPhiicnWeQPGXN4qngJy5
9Ssz0cPh8G2gpTd9PogV5QgLz4xmpRnDwZingFCIISQe6cw6GUurHq0H+Av9Vqrc8VUoK2FyNzrj
owpuuXVJ+7KCseUO7qojq2wSj6RFcLCC3BAKRcR8pz9c4brjj+2EJ634ce1rRumQl8L22YdqJFwe
pYc9qRtPu/FLRmwfGWMD9LN+z1SbrH0YoJ1oGKGiTSIM27BskZMqkaVR8KIFZWOeSi9hjCnAkmXv
w2RP0DK+DORpa8xqdAj199sQhwIem4GWLzd6uM1VAU2H1Ij+oTZaz2XS8DFMMuzT6/bpvSwXafs+
UPlQQzwCNbpl1vYP0bTlUzXSmYAkmPvugKSe2EalhYbTu3F06sM6vxg7cJ2lbQ4HCSs2O2TOwdIw
zs7RmE0u1BtcXKxLzEggB/FOCS7XLChG7bfFS9HBUj5xAwhKZ09BD351/fHVl1eOGKPpske57Blq
DeuPBHGeciRLE2vouI1X6w32BY4GRtFJjRszQ5zsx0ClJfdX7HwRmlL/gOUglx5nwYdDnhuQINyS
BoizUarnHuijVg+Ahk76Z4zqqKxryFMsq1JO3EFAnK9BAazhYkyoijPlNcr3JcqgyE4hRoQ6MX48
oMptsjsYQpeV79axmSfyVnaczMenwPeWLMIT2ZrrYPQlbPOB0ao5QXa38rsEXlglrwOE45wNNIKh
C7tpM3iMwgCLNVNzigkzx0+anWVxPPaQI1qGpMMoGOunoVeYueYxu1bSUn3nOcAM7jFv7D3up2o5
xF2xfwffnwiKU9rEbyXIb53O8yhxTkN/7u7mRuzevdrLriPNjeoaBlB+tYTBV/L927aEbDd/FQIR
KtIo8KptuwM+cX5hs30/ODo7kuEm/tkdsqsYf0ynzAll2Tk1w4y5UymMbWX9H8ghHcgurnUB3qKY
LVhhbXDvQqCR8rvmesmj7fzDmcnB+GjHLEAdK73uVOtPZGSdCQdInjXhRatWjkT6lulChIozDfxc
R7BFf+NOVi3umjLooFwMhgm6nxmB0uozFGGlWCD5yr/3OoAvbfZfiD6GSRriYMaQ0jLHv2p1j3dp
bupyV3cU7JfaMtghJlrO6dF4FvA4GRBrSDaafvX4v21pQ27nbM8/DIW91D6kpz1lmPNeS0wE0H9L
qxk22HTDWU0NEe3uxL7GIj5Pl5doqu7g+4n6QyXbH2zTukvxePUQZePF5pihtH0D5ewjGB1WqT6W
v+Pl4498u5DWqOW1MgzMJglInOrBtS6T7cRK6r+mq0pr0VIU2GdJ0YOISo0x4RxXH8OcYKFk1iM3
Kgg7zTTlYSC8vN3Lkw9GVt00X+TOQzb2hu0zbOfeaFwstK07HPZKMMALntjyp2XKvfLyLCRaIrgq
5HdeBxVt1ofXz461bMe6ogouAfnsQv5DzljRtnxdon8XJxZrbG2jvQ0IVZyyjFfa0Shiwx0HJcYm
olVdsce+sdGFchvr692im/XpV7QyKVyeT58AAPxcjyKvJqP6PLCDpiQJnrx9MfFKOPNszZ8DMwjb
Ta7KG15PPTJ/6AbLZKwza7I9t+PFOnOV+fVCZqdZwkdrIE0kxVVrZqu8D6efUIacZd3oZhmHgj/2
bWiKwke3QKM8DkbStxSnygsI1gCvQ5Mghou1wqXx/hnPGi4j+VFTzO8KgVsreSpHx2gh/KV5Ajn/
dUppXiwEl446HjDpPYq8wCJfZMeHPMAoKkxdqo4Tt670s2nGDeaj9OBSMUlbndFmIqoPLgUp0FnC
bXqQTyagxNoWqHeQiNFwn02Ztm4R4X/joF2ErNbbV8foggYbVvDQUygZm/KtiH3v8QAbXnY+iv2z
FSZ8CrhbDvbQoYLAGMIs2v+J1pPrsdejz6BMwlbZfLSiEG+5/jUCiIYcU8E9WzdI4GStmVqpzUBZ
VnRONk8wpmvt6zc9tLYFWCC7i+PUd6NEKQ1VsB4R6Sdmx4qxSS3h0LuXGBEewZPk47/mTDtvKvz/
nRBdi81D1tXJh71EUo3NRt8hSYDNb0DzAOMwrfXneTSCDVshTWte5pHMSfhRHjFKCnhYvwgbhuD9
leqE12+jY9MSs/i8mQcaDWl1S4FlxjymKTG3LIfDSqFoG2xgSKcbrDDjFEp9ImRfECgxfkmOJT+N
2nTct3JStl2uMsPalcfbRek7n/+3HH3exGMNsbS5x40bVSAc+Oru9KpD6LZqWWJEzTu6tX/0zjhF
cF1G0+gtkeor6Jp2vs9M0+ASa2eofMusM10X4VXoqW6ZAy8iaIRPNkh0N6gcIY/HFTDePA3L2f7v
a5Bq8z4O41lmyMZoWtANZucx/cGivtpuE3ofE7I7cmmo3q15JteFe9FCclGC3Idoa2XRUc273O/Y
DhibGv4CPvwh37lcnqNHhiHBSudCf6vGRRhXCc8Z+Wjp8835YQqhAYQhoK8J3KKLva710bC8aPXe
all5GKqaCuMUGL2XUZjydDHLuMv3Jg6w/ep7wknh9Qi6D3zg8bI/Tsvot/aOGoHRufuXgbTp4mPO
+SIManYIwuKmdxP4IAmJGgxOOT5TK5k8U+chfDiTSTH9GshiIXFnbUg2GtjRGMiZ4L2+4YOA9ox8
ljBjKz4/b9SNAL94IP9sG1NFDl7v3irsOrVJMfQcDDq7PrgwLXNkTgNR6hTanEO+yui/sbbp3aAb
xLW08WYKz41vCvrLd36W1XGC4ku6qrnCldkFj9j6/EdcBxnjAVmm/HE4ZbUp4ZTdxQqB7XY+lPrV
I8OouT9XBVcs59NTZALCpCgo/IqlmRDRMQ0y0e42veNE8F3HIHYzQQYfRqahhmycwbfk7sETBwAr
dEK9RBPzthPZDGMRJfj6MVob25BI6GYmBjnOMm8rzPiPxL89jJC4VBRvcVlfmyAv884eYUn+BBNb
NdleVzdXb9CKSsqA1T5PCXC+ok383cDJtnBl7Y79u2bS8ShGhSkkcnUfVjlMIPM7zwUox4FhuGKQ
BVKdyar/sz0bGcJocvJe2ev6/0TjB3E9PKQNo7mihuQPVpBdaOcrCiuK/nax0D2z6O7eCaYmk+vq
JwoJEAOiG8Pj4Eh26e+hycvyxMqLj9O19SiCFCycEx+QFQAvZEInMWdjo/XTAT2Kp/BjGNhwzIAj
6Yc1EIzIACs1ChQqvAZWIduHmDLW7Td9DKxIlr32/99YcghYyzL6FhNRzn2Zno96N2vIWZDvhgd9
eQHT04IHRzf5A29B1XgEG0n0xJa/dfpiQClGplLta0IPVDT52E1efIkHH7TTdUH7VX1h4BBkSUTY
Qy5LfCJzeBpo3XgPwfw2n5WkwWXbGkaI3JWLynct8DpwHSN4wyZ92dUQileWKn+4lbFf8JJ/0y8K
Ac0EEqyA3SoHFJoeq3qwbG0WYX7Bmp98c3epqrkiZREBplW8Xgw1me3k5NzQ+hcBAzdjGv5lFA57
trUuQWETBnwIWQQfazzpPLr+Zp6SXSmi/Vhh8FENVyXNc26P8NVx7S2QWCYMStqfooaj71CSX5Rw
SMKRN0WkxufPQ4LaHxVE/w2Zy/+At0G+TMv9OHXVVpqviFwtAVBF8Egl5+h7AQu6prctnASSKgr5
9PkcfTotYe1ACpAnaOwU+HoM4/fG5+m/21KbCt2Qude3K6bUBfXF2heWtsmlJxpGvPhmoW5fTdXo
awvB+bqmG686k1FuHOp1c6lT6udnKGZgYS9SB70IYvFv4Kfj5FZ5UI8EaI/WXmBEPAMXbuMlF///
CL4xZt03Eb0iad0j81zRG3m5fc1xIfkEe2dGeAJ/yLVrfC4ajF84GKST7HpOZuGIopnKHDcky+9m
c80POq6X803YEcvS/0k7+EF6NVP+DPZfbcbfpSv7gZcudylGSVapt7TQu48K2h6eStflEuSnsk0U
CNzaLj3LgHlHKk5zB4+E6uK7hsAYSU7Y6V797HHXvD9hxuF/fp/sNH0Y3ESOhh1EdUDiC32IDW3Z
4Wr4i+JYhIU+3ik+LFdDfoX9RK/Bg2cSmLZjPYHFRbviscv+cIlyHy8PBlQoI5K2mtBMwwFOCzmz
rF5HSYNVM3FGKSNnWYDyGQIY2s1xserZ6DChmp5tsHeT1bWnjudGdPjPeJa7DC4Q6DPm2RFuW9EK
aOkXM0M+X8veua2/lmU0zoQVCnl3Cb9z585cPVxLirQCwwCkgWWtiDHG9U/0p+LvJvuifinbSZQK
ADIsSCyVfsb7nqId1t4MhKAoy6Ug3S4iidBR+T1OKQNveTVK9qkEum2SwG4nV/LcPPsdE2A6hyUd
vlVGixUcbIrtxcd58mckC178M4bUFr+KnT0UnzPPxaLJHtS1Fucy2rlYelJbuzAq5+5Xxg2sj3t5
n805mMFHt3VbGveTp4o8ltyzUq9Eobh04lXe1/f6UGhN4CkX4IVLNWmKVZO0xDZcrDoV9+sC4FM9
7b6rF+6k1xUTgp3ZWQEU0GBy7e2Vxg+rlsreilUpaGTB6lycFC61oiHXeFPJnEkGKWditfkJCU1d
4JFCIwF7//fQuFF6xVDf2LdX4hHaMdUqjj3b5nUbJkBcJCnLD0mN8mbWieuzvz0r+1z4XpH9jW+Z
BX5c9rz6wFmXSW5ydRQbRC7PT9ii7aT4Bwz4opFnzOXvtu290LwFYeBPrXqzb6wFt1eaZ7OgGD6Q
8bLQatvdaDCOe7YCSN4RXD7eN3BchDMOIT8JmmDq6H61AgzVHtxUKsU7jaI0SdvpXQNSg4JarniP
Y3g6jT7ZfWWKAdQyz+Mrp93SPpYBp96i4IHCW37kFloFC2KNzemhVirA8Wh2jYWoMWLlEgR4XxrP
1nGmdif3O8LEAjSSoLIh1+ERTngO2sef2CmisqYkv01U39EF3qQFvee34Ki7//ndZF754B3OEyfG
sxfagztIPhUaV9jxgzEVHlYUsiWHCO5SKcZfXWMx2bKJX9+IaVvr3guVyzvrlQIjr2MLd/3S3r6g
7cO6iGPswLlTosq8Bw7UQu7YDspv2Y4zFFxAGXXgCwEAfJAaiSo3JZtrbvVDUJ4f4vBP6qMuTi4Z
8SB0i3I+Yv4d+lmxCaan/USQ26Di9bTrpMXwPFtkNDSH2YIw8MrLRR/IGqSU1WM0SaBMgZPvLim5
EsiBZ7nlQzjsLlwwKNmnVKweOYDPC+kDMRmdVZgdt/K7Emqg2QPIln1NqayA8eDnYRzK78UVYh4L
HAbdiH5Q1bqkV3LzdLC/9nTTg8l8tNT+enHixrIRn7RaRYrTqf8gzYvNrp0RIAZ/SYFcjBFr7M8e
9Mw6eSfm/ZCenTChbjNKMySaREs9cmwqya/59mRSkIY9RPmkLNffoB75DvqcYyWjpvA5nSFBrtEG
18CuqoANTXO6fnj/Us9Lvy+0Mv596U1Y3BzKPSSY/6NHWEcuKpZkWoHeN/A/rEiXcN3G7J0GZEGC
2cvaFbfr1pRP1fQdt1BNPg4Js6GGgTN75I/e/ltRRRtzXMKwJieoWHb4OJp89xIinn/wuI2arLTs
R+TGo7laNbmYnBftmkz+uZPl/lw7HzSYU3limLQ5NgTfTZLxHwHvyLf0/yu+F3FYIw/tLbmcF8aF
9x8gic60Ri6SZgTxvjFhOrVaOfWPWYNO7vSlYPUXluebd7qqPm3YhMWfzS4/M1wF+chEcXkmzxTV
bEQUrMBFYeNJvQW3jmKoxNRrkLPBuytFkoWWH4ruUekPS0nX2ZyI9mMfLLoljmvnjtWKWxhjr609
V9idJ/hnmTWTrL0baYSon/X7oOfuCKwuT3gqBbjMCEHlLNfyn9g+M+KyDfZmkBuY3WMl1Gb/fmPc
i0i9tBteHaEWDgC3/yEgQl/JnENRpxvoiBwlLcQVB155PJTtzOzl0AsSQhQai5Uf4Ak2H/2tvazU
K14dF4BVlV6+FDOIrzk0LI2hQGPQ8/hU/3QM+RZopLHH1SJEBRwNTzsgcGXw7lK/ToNpYuEqT9xc
W2UbLSD9Mw9PatST8ploHrML7jLqLFWrGSeWdV9KULSugvUTI7GvEf4ASPs7KZyncTKGGVLnSTlc
XxFhSaw8sT2C+vrq18sfCZGFP6l1Iuj8YEdF5xd8WHe5KCm1XNBFE+gG2zTAh8wrRNoF2Eevv/xt
GaJZf2vW9zLO3NPCYM7hE7yly+zECR9+g7c6nqfDE0Ct0qvJHLTkvJnjQZfwj8LQ7sf2EjJChnDC
L3mtNJkd0NJb+bguxiaecaZ4Q2Eewt1hfrf5zACY2pmabeOw4hxqoQ7lv2c50sRiinIzkIIZEiPy
YZhsL5rg7MbggqaCAjLhbFDOQxH9WX84l4/w3nzy6TPjQxdF+Z82npRkNs/NXlUswusstXyoUOrS
T6qxlRxkwS2KupkwM3aouua7mqo8ip4jAie4ePuE8fO+ocQg+hkCxIX13EZJcF1CNhByLPNcWeRf
ytU+mBE5Y2SR3xiqIhClbLvl+plN9ClRZjKw3TxFqUGstR6ZhXswdvIXBGZwcuSdDjk5DmJIAPL5
/+/tCwi2/Xd6AX3NP72wfpT4Ro0GdzaMTkeAqd/y4tiKjHZxcaXvkKFka4t9TsR2mrOFiDr7nkIa
GEomQGIsXqjDUvFPQFFsU4izKWVI7T8X5oc7cY6CjUbR6WbJKKKEY53AS7qcpBovHoFdlv7JEro8
6LsJHeCwdkjqOhNuUUA8Rc/5GKnUfMGtkTWi5z2Om0c8Euft6XEg1mAq+yOyzzx2zrYUaPDq24sr
/viLSdXRk/mRCBdfCWBJJzVDFjkUYoodadonLLziU7vYV+c5AnQldWtqNu/ShZvMXVqfcX9SwFU4
8hfKEL8MpfLlk0bijqZT/qSNfusMAT+/dca/zI5UcSAWqR379/AS9p6ezMHn7/jaD3r9/9aVuefn
tO6jiCj3nDVPpB3J0KCWvLj/8R7ThGAl7M0EmccaNTcV7cb/dupbBG+mvscUK//hgkwPXrqVIsTP
LUrRhY9sC8XV98Y7OHV8EHG6CvWi6yl2Dt2prrPWmKboYvFIzUNhnN496UYJYLL5M/csr4PL317x
XNu3lmqsyL3iN9qzbeSlbEVbNLCLofGcUFN0qUU8ODh1cXiUZEvMfMC+2YupLIbN9d+SOwPmH2tC
+1pmaV7YPEZTLiXaye6EL8jr+PPcYZhVG3QMM4l8StyIBiLUALLTMTr3i0YbkwK+YQobmYXo8e7m
vLA1mpL42qIOOI+LRhYm7uk5oMgPybGC8Sfj0OxoPqeaW74fJeb6NnDPjC7Obvy5vYynW2+yj5+g
BYp8uAi3kVMiVlmcso4cTs+51L6cpQWmTfYgTsUN8qwjF2mWgypO8oZsi3zRT/ubY32rbOWF7jiE
kqC21U3F3r/YDdo2CvOVxYJOFXxtdHPsz3VljILH3AIbsjjHFyKmr7u0DpJ0LZEZnYhCDTRtEV6S
Ic87zy7PmqIynvXs/guv3Q9Il5ZQYAFtN/dancWqgNDrW57cX/zdXNprktSU6/sgk1NyPDyQg4gI
8uA1P6xv3/tPu0P1PWkrAQshlabxdOrK4po4hkvBE1tR2Dg8QtZEdhNfMxTkTXtk2B4Q9Ts2Xn9o
bMFywlMamIeHRlM+S66HMDu6K/P7m29cGA0+ShYuJ5RJYC/Pk/rICQmtw1mGIFYvncHpJl3HmWRX
bw+zup4IGd0OpDt3xo2ZVE4NzlQ/UGTTVndFH1/b5sJrNvPo+CfZAnAxHnfkB23OHfqUzLUi/chM
RE9vzeb56230c2DE8GhJV8dMdF2t7yoOVXqyGvzyDqek6XMu5Vvf+7z5yRIkpq6MhpkIXwGnLy1w
vg24SGk5S6a6KfbmGqnzeBVJz6uoyLI+tMVyE5ajDpQ1qM+AIRB3Tm7YP0SfX6TC2dDTDKoyCY4o
z3TBImymtX1P/s3CfLos9eWeObTXqmf96yEIrxWVce1wDlVFN8MkmQJ+m6FgqxI+41HfLyNvsAkU
z48PhUhZaYQSke+gzOik9xLlyzOb6vBwfWgXFKr6aSZWgKNFTUhpXO+5gKt/cxoMtFoFen4H2vDs
ZnDpLJHheOUaGA7DAcoATuBp9IDCfvVPeGwiJrnRZPTzY9BWUtMF2yr9eAs1O8/kIZG57ZGm6hhQ
D7EtfDQ33vlMIGbnkxHLRSH1UKFKYIIb9HLRXTvu+iiSkDUut2VdTQX+Z41ly4KrnGrzpbzVAITY
ZxhqDa1duL1wi+MGSoxMPlVNukRQD9k7CEkJYfCIBu2bIEeVWDygtiCO4Hh7cKkTDdGBI0IhgWQJ
jafseu1QELpb8CRzJNuFFGBLIAaM4ZHeZG7UZzMaPxHsfRJhfGyz5cK/+wk41GdkT45tbFIu1AAa
QraD+58dBLC382w2/hQsvH3Lfac4muaDCoqyBfNQbG1D67v/ULJlikNeIAOfvgXzep3IX8x8k7ck
cyYTEhneSO44NvBrABKZNF6986qzIHufrPBss8EUmwDrMSLCZbXP2WXEGhMThM2WYtLeoMGxa7r0
Oaq+W++AMECgqaq6FEWJz/AUeEBWW3/y5LWxBNt26IV91evbnUb0L2QccBpaedey1e5Dg4ZC359f
zcijE7sITI2Ijo1Xn8Gnuj4Tun6thtsnKNoOQT6kBNcijEHKhhh73cKyPSIgdFeJL2N5oqGT0KJn
IlhYtOqkS8zcC8SQQu+Dv3nq5QDfYg3znzT57ViHdY7Ty2FBAVO42Iq9Kpx6XiFP0SqFdAZAL/yf
Yu0Trt5fQbgG9+pS5KBvwHryX0osDIFDOBacADLWuWRo/nHuQrtm320UiouLgHIrMR6wqadupgQP
rQyVf8p1URIgGlyoaWjz/s5J2De9ZBYvUOQ8FsKxyGI6FpDUGa24a/fMeDsl8CeLGV6wrwyqCP97
11fIFeLPpWxzZkmhWemCp1i7dDkgeBRElRmPsgcct08K/tNpW1x2UAywtzAJLAa5JDo3P/5Dt4Pr
bdQm44Lqo0Vv4bQaiVGPZILm3199vpK9Bf5X2rVtkygWYjHWF0/SNpl6l4bqT8NzW1AlaYLrtIXB
8+EB48FXjxzHZhMwy/jTbbQYkryNftVRm+crymHKI/TlJv9P6hfEA/kVO6blvd8UDOgcTvWuo1oH
PDkOtEuQlZq50WHpYivgeEDiOqLGrSJbqfrJknzSElxrDrpegvTehPFstytch1FeJNjlOHcdxitD
UfS+58/7XdYKs5gJfkQ3y9Uw+eVtgKLMbsfyQj93nBEqseM480ZTbgjlQN5zVJGBS7OFEbmw+xHD
ab/vjDKnyCuhEgFJG+or34fw+hiy6jK2JqPNSyAp0Mn1d7FNA6SmDXy6BPu6k2AUOwE60265Xy6A
FQxLIquhBnI2udBkuY44SrrROrFsD9SU30xL9FhH6LeRBgJKI1imDcieJrEDQBhErBMtM8uXS6gz
448eJmNijiLPLdkVOqHeTBz53RYSWpycpSuLWvsk+/qEOMnIu5hvL6y/GBZCCQTCeW4MvddJWRqA
spqDvW40LRrDl1ewZbdzhz0eYBUxPWCkcgKtK3K41M1wTI/AqMhbt8oqYJNkO7cS5QwkIon299Vt
k/jkYp1ampC9sFsG68+rF9DA7FZ6HWEsyWJw8pcqHO5chyWdjbXQsy3Iguei6H/UYFbnLZORjxvw
LosBqAyLn9twW+K7jQwSWHGozOzBXQcgTV03ZTVA+RsPi43hJg+C7KO8IKyDDuRD6H1KfcHOBO+p
MA9lxAcJ7nMVhngXIh9lwjVnarn/JNeUslvy4m3IoDarzPlqm9IxqO84RjVFg7joEg5U8f+3bw1v
UXN8dRdQLG9+waVm9n+MIqx5TjR3gWGt1PyWGc3QObNcaQnVKhzKoLKPfkq1BSAiajnjT8iydoKq
vePpyJx0FYA4/Qf7yGhQdiFT14A6uCV7ivG+Ga4Kn++uR6XMWtexwmvUETwuutBdbpkXY5Jvuk3C
i3GA2NJ/l6w6RKKaNn7Z1fWp5uauQNSymsHAsXt549pw9h0fsRGYbJIzzhU8D0BHLunV+54NMsRd
UBTIQob9RinYsSE11S1vnpmrCKOziJCN7j+8QGfF0rtSwXH0dT2+VONMtAsjxCYqTB6CdrEV4G8/
pKHSH0gf9GvhNe8e6bCMcNp/B3mM4SW4fhGZeCOdyj/58/lLzVXvR9K7BSbbYKJogvyBUK/0Q8IY
xSEsIW0xjWyrVtEhikdeD5raT/aak6GkZfSs1cOCz+9Fi5yoVlAc+cZHULbvAUdiZ12qAVBTmgJ3
67ftkcwA7sqL3hdRa+z4rw2KD7Ii7naLmkaf3JMFYeKd7kkgfSBJw9GNAmncA7edVayre29I+7UW
Slc4/WplaSizArfUsJlYubFcXR+mK7AwYwQHfy6Ri4jjWmVOW43+RBUkVpq831/Pg5q/veI45qUs
TfSGaBaQo5XC87qs5kz+OeQEFRIB6KPnsiM04nMfk4YuXaQdUD8715rDLJh1R4BX3dvWJjwxJW3a
knajUmvtlVKCiCRIId5+Bqg09h95Hu/uLLU/c0e/keUO0OZtuSuExf4EA/iwlbVC4huINKDJ11rP
y5l6Ss96lOtvzZVoB4V4dsR9MN8AbCkMVB7cvzX+y1Xu/Wc4plbfR7CMTD63pjgFQymD6X9zM3U3
UBuRPJZy4LjZbZ1bfXmLVwXu/3U4wkrKdij5uzyW+8m4qNtf8FrQ0IwonVEznGd/YMinxMJoitA4
MxWWwdSXIao7irDG1hN26lllO4UUR1GyysspftVBRcHWW4t7sHOk1bbU4BfHSqxCpiYNJUryaZvB
osTxbC9OIknOmbFDbn0txnuqaqMFX3oNPpwN4JbFNYzgKJcJYVOhHHv2wUEcBFbKpw1rDmAMVYha
DUVDzk29GDsYWlFLlPYanjqqOKPaOWo479tO5/wXmQKokBijQgJZDpFeFSr8hvp6NXm8KNe8lA3Q
zRRKdyyLcWzV5tkU3Eni6N7Rmf2e94yBrJ16DbsZj9urVDNMTsU7NolrodyGhk/cXMYsEIRrTZM+
4qWb8hNRJMMLiXC7UPS1E3ML91PTd/EJAiViUzm30g1QB7zwhLLI3TSeGsUvBjL18GmYVy68c79U
oM/3Ho6OIo0arc9xl1Pyefb3vySjX1GBjKTERr9ZVlU77o+kDNqXhYwas0owTw2fp70xqkrTiE9X
Yk74F/Gt20qSL5nzQETASWS9oRYWq2j1ZDTgumRr26I4XbE7yU6Sg52ufKPU7Stp82tjytWoakm2
wv8t+Gsw+rz5DzeMle6IqC8T254Ikat4T+1px2svtB0qyNOe3TNCG4vk9LpKxhHuBPCBV82kQmRM
Ejb7uUeAD8PhJMUZ2Q5DNfWSAn1Vv7DR8VEqNKIPrqFtiGiDV13XqQUVPAyCgJIgPf9EcRvLpWcy
qmo2TNOoMYxFDXICJ+30dGuvzTIrgcKh39XRcI2QnDY9hdHhafo02406qD8/tp9R5qjY36BDewnL
5VDl2yGI9yOh1EdS4yRxhY0LyWK6LZObfVsjOE8vgx+Bo0xAPrM9dt5WWLirtQnncZDF2zwDr3hE
WgLIlLPlruAyFdPHCRhpyFnsTREz2R9Zy2bq9chqtagufTWsOIdiQMK6Uk/ibEOkord0av7z5Bvr
5+omKQTHfycHH0JVCcUm1nwt4OZYZIVhqVo38CZkCpHGf/vXQu1xTdi0vm7ufY1TkPbHIyXlFv2/
LD1cK1P9r1teI2Af7sV+PDWUNEsHs/Wg7DpHAUqsTYS2HLLOBvfHjvm4ezFisIGLe/kLuqao/Isw
2w8tJhZReXUkruHpX8/WXOCHKIRKSpKN5LzqCK8CSxd1ZGcOvYqa0LwPBAOO7gRlicCg4m7X0gCe
1OccjtkNg1JC4goqSFyM5SM9S0O0QngefD7YQYKSwBqJ/2UP/nA/5Lrl8UnGMqL+V7qQFYZPr21s
Enj+6LMOqD4LyCTJd8ZHLm15dQMEC3gaJNJMQQcbBDX19Lou2l/nu4RkgdsctH49I2xCvXRr5z4+
tggIS/Ih597WsqYmLdXTXPLUslE/WgMw7RQHp4vtJIyRTAegjB7cB7PSqaJFzFd7SaVC0nxgAMTG
IfkXkvVindC02zs2oyuauS7lgMwWfE1Y1gb8RVXIIBYIqJnmZR/6dQysX2n54VmoN15W26rRhE3Q
E11mMyeq7p0z1dRY3saWFCflXhGcWm7O2dQQ0ZtKtcJT4eH7DEMZD6RRoTAkpFrQb51udk3DIC19
nVG25MAuaLoMggwMy+XReXNaAAXRr9ukHPx5yzTr7amq8bGLmblozrWZbGK1n7mU50TViCKxtFv0
1aU1SNPqlgurW5AGip1P/uDqjIUKEaOOhJaadzr2RpcPzwbAeOMXvQH5hsxmFjW91kQIujkj3HNM
+rOC+fWOv+B/ImtBkCZZnpX7KGMbxuVRLs1ZrEwDXPJjXA9XJsuacWEO31vy2V+mGw8pGDu90BMw
STHwSbCjGZQZzQ3ZjULEnTpVbTw6nPZDMdbPxwhg+24W643m5kkWuZPXC9cR4296D0bVKt2t+oZi
nf9neBMQeMT5o7WrLK5jkPeilwhRZqw+k/W2dR+ItR26XrqNkNBDQvvMqjkshWEeKEto/zLf274Y
O2OujoEl2PY/EHA02gwKq0AXCOXVkYm5vmphRU7719vpippi8KlDwXd8ok9/5hguVRCGpkZGc1Hh
83dolBjsYCgC7p5h9OQHoSx3HNr2+qQ2UaqGR8q9y5OJTBiHKKfBv7w+qmKveiNz4+ckTcd3WD66
djb1W2KpNnfxyEaVQrkN0GfZmQXxx3Y6F3Un7jEcWxJHslGxY3aidXxjNEWRBi1KZW0A7ESodtXT
oOpWNW/yIyQQtnwwZOWXrR8PqMsUidX3dQIdBnKzDopsbJrCIKOo4aJE4xVpkoK68L7vPaI4d8w4
UjCZGVRGyoF/l9uFTPJIq2DgdKfB3RbuEhRudue5rQ/Gp/idppWmqnUx7d7mpoFgyGOP6r6RbKN7
0xfYYMLE1uNBEAGvpoG7gwTx8X2ubQdfTvfpnepcDfE6C4VhLVTKGeknYFhEgxsSjXG4m+7tVil1
LCcSeJqzYbgN4mR/vURfhvMfA8mQVUzjJWwUyOVXxWi6+oaIVW2I93EQI5aPvvpJeNUphThKTyGb
2QvZm8ZYhAs6VZpyVS2e1JCzeaYtGMoxzdo/XVYAHs1KgJmj6EUNEDPF8vV5UY1Hx7mzqOgJdK/V
+6qVKJMqs02AMHZ7Z38fexYJuWcJSv4fUd8VEuX9JVk+Z5J8VQwhUOXXgBmvetXD/0XEBDIl9TQJ
uvqi9o/zfsXcEwpK9RgmAw1/3pqcwmiVxC7hLk2uWiOrL+oOm42mZlloDU47hewVvGt7+17oZ0Ng
mW0NNoyVWaGKyMhFcpEAyC6ewIEMh9pm02LdXc1ud3v6f16me6wmRFKRnxcrNgHHL2n/7iKbyhdE
L70EgOzd2UyzpsAybFEEb/UOy4cQDYVcE9gHqCKoXS/OBwpPZbOrO533NvwbzTkCIfyJjeihSCBQ
dH9ISAbWQwdr2UqKkdv3fqB530kvtjJKRVWJ1LmjgFe/82N7w7NF5CHNI6mIwKn3lVt9HjxKgTYp
llhzjXNqyxAlOFiSjdlknFUkjSFiSwjpt9Oi6PubIWHlHKtWsB/4htj2ADNUCaLJi07Czq4eFgin
4yvjSndWx5fTacJZaYIREN7JE7mi/l9SJzRkmv55+ooThzPEfZmPshWiyzhoC83LozLFR+QfvjM1
X0R3oxf9zm0B5XK2XghLZOQS7lvA4lvt1APx2MjhKoS2nzwbN4JnkYF479JunZMHuQ/TF9fcLwjv
uFIL0ZEGYLH+eIAKH8Waopp2mJlU79A9fWnrIfKklprrN0PaC+LhB9PP1Q72TTqgX6bvEopU8R+u
9GIwnOMLuqPQ6pZzTXPTMtCa5mFipfOTTNaEskkho45jMnxXZCZMaStZfnxjtPs0qcqWthF6ex+Y
aG782pUarU5i+jxMQMfus4GZzg8x+JsfLGotF2knOsexKH7Ecjxu/8NSYQ9cV8/16DQw8nN8ypER
lwns4JlZj/FcF5DAXf1hLCL3gStt26ErKgeL/QsSGdMV8DwPN9t41YtJGhgcLXNoeY7xirKxfyCn
DY+/QhinAQqzitKAHwUqDNiLWEdMpPzm/nJQc+jIMYfTZ04MFzAX5/H+dd4ETT/eKDXB+SX+8bAo
lJjtsi5o0KuDc+KSVzwZJuQLXMXUSx1XmUKvAMUmaYRyA6k1Jori9VaJG2kW/OiS8j8u8S6BZk8c
f2ruk01ZKE5870Vn9iC+eDmYBphAnhlNPGItQAylhOBhnZsGZVBHGmWcV5Ikt+WpBLRsTvasHGhe
ulkQqeQL14s0+ZIxVimRSKqQapY8DG7bktX8a/m4+Nqf40E7kjaq/9ZsmZXagKpDvxF3IcexPssE
gDcjYAzsQ1bZlAmanr1Tq2g+Lng8HyU4UibA1gVUer2MUG5PpaPP6hXHHROBEb4kl4rBZb72mWnd
kS+hRfHLtlfJJAvvEkQlHyJuX5k4kiDzsEB/Qw12PIfTTwLrKItB9ar0cAsQKtMIpxLiz6EFjNYu
jSMA/Ygr+aq8/QivWM9LCKU2kZuZom4ejAfSxK8VVA5av7FyG/FbQWCjYhO5eETeva7SBGmJVGvF
/oJgbvpy8rU1i9hfiOkZj83KEzee99Qfa/W9V7Y5yXw1zEgI7wfuAVSOoE5cCE3HSJGqmv9X5MDP
QyTf9QN/l5ZzWxxaTODwdC++kaiexvDq2/fZs1pah0i/0OF5Vhty1/PA0THSGbbnfpOslMuyV+Il
Vtsqf+gtn7eiLpB9XXQl+f/JHyRWD8XZHmcU4TAI1+WChr3LNG8Nb94Cuq0dvGKYGGR+xBU1XL9T
4gbg3PkW7XgDtCFbpFCmstnYtmYbff3GsQAN0t5tcQ+sXuoXRjtf9DpGvt7HoNq4cyETvJ+W4Eyv
pF8I/QBZha6P8ClkkmAjffJHbYRyaQV738vxm4jFXPfn4vfeGdApjlxj0CCnegpy8XgGElmgEkIJ
Q/wqMr6paiArdG33W98nntV/1Fe3TlXxD6+GYT71OU7lywEXZYcV5nNwuT2fh9z61A0tlIdYXjNL
yKmWIdYmN+eY9VisBpoMK4OFLqcxJcBvHohA4clkELQrBq8ctQNzg2wIjMv1m/FCIMrzG2Au7X/F
d6mWEVVd1TZhEcbQ7THHQObfs9Ld1Bpx8iiNq/YpAw3mzEtvYa2VLX1aoJCpO2RIxDu2AzTSH3D2
8Knc0CypGo4FQDTvS81Uye+T5wvY2lzyZR2nR9R//jXRLlfY3/z8wnnl0isL7ObujfxsyAvM24iD
u/xnhkfsvBp6D05vRhyhZ1Qn6965rSSDWwsR2FRvStg0OMi4zdJZU59c8v3DAbVZFZg03YDo8C/6
RG2DjO4E5LRET5WyHfi5BKlHBkTCuZa4YuBQfH51K5kT7OeXAIB7gwNyhV9Jie9FTGRKTilPkiaV
E1ZJUtPES+INmifqTyPPNrqWj6p8FBPJDUo58xX0TX7E/uPnlDFk4FbhOvEtC2LzztS1O9MZ6US7
7ESZQkGb3mSthw+YFLoBejg38/L5bD03ZC1v+GlvZzjf4SJpU00tjw5aG+TSn8JC9oFWqSj8y9vi
+IStws23jZ4x563adTXjN74LXnYDtPW3EP6JfMihMW++gL0mfbQnzMfxoRjiMFXPJNUP+Z6OcjmT
IynMFb7HDCUsIAUoljLIKLM8v6zq6UjwXYFi/1KGPBq2QN8BpeFF5mtfb+u3QJzVKoYcs3btM/Ny
oP/W7T8mvl+0zEtcRHyeYpnzMzGciUYjMlULr015AUkkm6CnvPsp2H5MVxAgu8fmLZpuzxb4poyx
H8SEB65Gdrk1KgAObcTTEBAh5wyMEUKxwZemVJL3xDoX9Iml6hg/q4Qj3PAxi44JH8zDwlRgyQJQ
jQtwgaHGVl6cMIKxhQc2zxamxicK+Spv6p+TYKSaMDRMJSfSAnAqgOaJp8h9R8XCvJhK11Wg6O1m
Y8E/U1XXWBvFiYHCWgswYl5T+vDuzofMVCLJMNJ2AgWaDKqC0rnnLLwgZmQFxB9qt0JnmndGpnAM
XZpjvZOyQi2W36QkNM0u6vrUL9Zbts8cYF9YaC1+l3Jrk41EpU7v1DTcEjNsS2O11bM60xc9tNbT
POidQ02lw6UmWDVerqrmRKPLOJNmE2wOTj5m7RmuAWJBytUkeot9H8m62jPds+0kdTH4d1Jm+wBV
72dzbX77IYuA+Y+XtVN8UqzFHDfiZBI5zx3/M+dhNdfSkw+6dhggM5aEI+6As/NUKGoaF4djGSP9
dvYdNPLM6fcrZDgyYH+V0jSvffWsEdZ5h0aLEjWTqAhKyF8kbaTMMXmPOzepaF7AwwLXpdTejMjv
ldwle0TCh3QG18H1209INfgHvuaH1JgEjDdNQiAUU8lwbX1kyJ7HnyPQDKNIy2UoBCv9a/QZ9LH6
Yc7t3A5zz/Az2y1L5kSUtqGfDjSpEPFkWHyq3JiVzLyumAVvq/VkIjjNPg4DzKNiKSfimzjN6oaw
xY2cQDsH7wcfNpPJhm0N+H4cSNgeqEp3HsP4oiCNJKOPpqvAcPT1qbx1QYaKLzx2wNcvf0w5exdA
kesH2djG4xWfqPcHBkW2CQhEyCCbbFMJl/EbODL19omGgYADPxRDTB02INnr1+RAo0nVbHicgDtU
AlemL1akxoQyeRcEtsUotSMsBzzkyvHPHjUdA6znTGNhlVCR/pQoLL9rhbTS8/M1DVUcSzQxiVUQ
sNBNYqLT0Z5pbPiMwZovmWesHdNuXSVud6IiEmlHeLRmVyPMVw1E596NaY/KglHWW7CKaKcWQoOn
c+ABHDwkxqPmnA4c38z7pG4vmU8e7Xw1njaprwE3gpYb3TWjBDfKbTlOAGCORNcGuNbtyv0yTZ+q
32d2aiTukVanCUtso8gO9yOPvS8wY0K4e9WSxew30KsajJ66TY941oMl55QCV0P04g+ObPE/xmaJ
6oM5KOZHArgwqDbUC4/ojMNUhD4msigOOvvO9UQdfhbzOGj8t1RWYR8sKPx/gtoJLtsfgwh9U3cx
ODWHZnpLL693m8d+pgweC6DVGQVX8oXNIdCihkXFV0vY6KiFRwQ3yaT5x24uSufWkWafvDlrnAn2
bJnDli6eh6lytGiQxRVBcrx8TiykL5VU3qGfTL5sAR4Iq7J41S5gz54SsXdOraXvPnhRL/sxMyyO
ABfnYh6KMjb5ytk5SUSh1i87Scg+ACF3gckHdrmKLIyQ361CKvf6LFVespA+vj8ndgCzFi4uhxJa
hn5lNOMHd4ZYNvohx/tjEEsXG64uRJY6N+U0Lf1XodwCzWm6ODfa+wR24BOxFsi4qwA+hvTfY6gp
tNrCuVNYVokdjoIMAYeEOp1j20Un/YeKnZ02vFvK0xZhAKEMvfo/3UPpdWbknXKrsY58hHmLXckr
61ZXWzPw4q3qNUf/goJMK0/Q3dxaUJwGk7b9G/s8JPcswHgoeo4WU13cefYL7wrXsEU+xmD7gCtV
r6cbyVNyqoG5Xux6X/710bW1BuAWwrveHJKr2KA+P6HkkjChDzfyfaCIH01cg1U19PCZOIJEcG8Y
gnpRrwzN9GAzWvlqxQlo+GXbpQEDVVHpwnqqKw9cn8frI2vHoI7+a6FkpgOPsMibL4DMdwGsUbly
Y2hNGlgjZQ3jUT764fZ3on2xNkxVAIaibHteMw4Cw4Ph0lWT39O9fZmWgGS1y4Wir/bubvvp7e46
Djd0RkR0tSjybdhXTvJiSqauW6YcdX9Nf9g6GF31OmoBilmvvwkn1QKO+ymfSePtEw6yxM6r7msm
TKLV8bkQW25sIG9ych2FZkQHKHCcF/lwn7z+rkXzZSeSYMsV/2E4qCoQHZ8Dljr66yaQ9IXuEeMu
nsEFmA4iKU3lnlUYZ9UXViVJRAXCz4aw9KRy20t3XAqwSJAdAUDeN2D4eckf3J9eaMhtZNzBY2m3
Qq2zAvepDK/MASj/QOp5Skx9TuoGcXRt+KaPVcL7FJyEVm3fiT8cN5otsaayrnBvbpirvPtD57Kc
FWK7R5ObzwLl6qrKPggKuCu9zkHUE4DHg4GKu5pEoYtFclTcTefe+P7wE1MzLy3az3jlq1uPpV/7
ozclBsImKHkQsJruveY0dRwYArecX9x6Tj+tFJ73mtmtdUQ3goi1xM3i51HzrPxtuXmdgyd9r7rU
08hOi4j3ELtg96nOKR4et7HNPgtnADc4+RFKNeBx/fNaW717TF2IT4/BC7VJNw/T1um7cvtCcGIB
6ENZBP+zQPy+pu3jQgcVVua8ozZaWeNZ5/1QfRWNFTksNcDmhu7YVYnepaH9jCpuFSkXmIjUNL6q
aRTNRg9D38leIU/dVjItp+g+Vannol4oZVCIzqgN0/ih1YayLkcn78dfcGQnYmQAdMvADTDbGFIY
SCNQNoPmeyyfnI0bxBMv+tvqF7fzSP07v4UWO1pytJrFXhg67q2A8wvZaPIz8Ey5GJRoVyxEb4ZC
LX0aMtHds5SD+gJYd+Jm9XQCLRYjua3BkSppAusto1LK7F6utVKqFrg2Uivz6aXKUBXOz2GQai2I
21W3gZfFQoWqrPrp07ARxknwAobEBpl3aDNknxpoEIpxqRtsyVfv6Epllqu7S8A+ouQkoSxwG2PX
3tFOV3Z1yowxn21p5u62xak+bGMcYQ8VVUJCwK3OjqPHYN4XY03/VlFZzZ4rw1IDTeZMmoe3lq8D
EpmrWP+nU80jtXDbPjVbQ9Av3JOLv+YZqnxzItzUeTi77txStv7h/sLERNdVKGwN3xR1Kuj4ILvv
zp9SU5fxNCVTTwp7PnrNZEl+bVNlkhxtxSWMqc63elANPcOVjthmkyHoGvkHf5xIwYaF4VYcPtdN
IgJsTcyU6380PfP5ntOJxbvBgbrQj269cJ8LEq091MUsiO5ncjt4D9/NOfFQT2GUKHf4MFyyiLHB
Y5ZU9gYWwzjxM1DV6yN5HQzH0tjhY1CjFjHUEiWxSAlzYzdK852bCgPnNYjsaKPw7KmV6NAFf3+V
py9eWSnnS691ZxYtubUs8PL3iLTd5cNRNa0tmLfZyxJX22sO1wmVjkFPuEGO7bN5Fs4VipDmmKkq
bZKZCKT2rtR+BEA9yU5yyY7x+zdN6NVSNC7BadmuDJ36CL0AO+TvqIzQTGxP/7qqHCEj2YPVq2Rb
Mf+cQHrDZbjsowHOljFK5MEpKji2Pa7YKYyMk7uP6W8Ug4wt5x5mu8AHM05Y0n74zCeO93OXeEry
5OUqnrFujzPM/d95LEI6Op6zp90VKXMDx/AJufDLMogftrVhedtZoyliaDjp4uVAO6wa1BgtLKAo
upumEtyax7UHOAwX0U8XUMEAWMkAPxPQkUBDFQOya6dTTKa6AHURw6yQIjFdXjp3cInUdH8noK+f
rDrQvxUasMAuhgqE6VLi181+zpcihGYf+ollhY0l7EPz6S+5WfyLeepbNKl6+qIlvlVW3HFMW4hl
oN1Vr5LA5n4Hrr4s/fKKmvJmRKVhBjHt2JKH78fv9ZDF8dtUr8/FHBbUTWlCRePVz1GEenUYaapd
EzbJaLVA5BaFcZlZebb8VQf00UWD4Sh0TWLG2sWQv5nIaVao9eemwlQVY7oJHpdK5KAmALM3qG74
uFY7GODFLyyPIRIg/LuBDx1P3LAPBy7ECQAIPytuYwKhFWQ3OOgmeiiZL6mMHjO/7yvMZlqEoKWC
yJPHa1Euo/YNxINQZuMPk4xcx1Nk0aYjiubJ8d1AHefi0MQgade1F3GtT+/Ab2dYC2oED7HPD1Ai
dVMShyEpPlBUotadnYu93zNtTybGPxCE2vYt8QpJ2wTusTIEI0lD7S8UVXF7MY37sF0RTWG7TcGc
uagJNCxXnptxWPi0voSb6P0YRy29VVEz7+xlmRluHBdC/6ZQS+pH9G758elQVXMtatKIZyP8FNuR
j+6mU/oSjYypXdTWgEZTpj7+aUweV2xjURCeB4itRaZSS6oZX+vBkplo9q5B7WH69HarZeWgZaYs
GfxAwS7r5HDk1v0Z5S1QmzeJ3DPjQURqdMQaPl62u/ZMWYYz2k9Gie9lABs5pMve8KsPeZSH6qOO
DfrqbaH+UI9vc1bTrd8MAe/ZhksZF6FNG075aombSymp14/Z3XwgV6RYlMeVC33YFa/7Y4ga1uIh
3JXhoHzot65+eQYm2/v2IrWi+scJjdR3l+1SEi2oC5V1YSg7IfDu/lvj01aDubAxP+QSwG1z23Fv
fxEiAQ/qW8xOO2isnHQRF6S/xVbotkC0xKoWuMuOwW5bgWyl0rYyKqRbSQbwdZHaJazpnThVkdO6
vxwZWqynOxzk6zyzCTsZ9Fzi/hOV1IWcSChSCXv4Ch0Dx2u8HLwfO6ayD9lW/ByNoBew1H101BQ+
N7HuLVfLofAhCFS1FG5LSHErVKtz/ZwBrVnNdodv3EtE3S1FSxvsdaEJvqgORAbzej3gHm7RRUgS
RT2flL2wHIyTTFkktlLQyV8c+OUrBRqcVjJKcNenyYgzxNGPg9Jy8SHnzE5P70NXtj7M2wKwj/QQ
49BprE+V+CwLn+x6aRLVsGlJ/dzCLKRjAKODZiwz9OoFeT1R3UO2LDyZnNERxqsFyNEu8DpQKz+y
aOFYJOqwMJ/ZoB7COfweyMYtX1XJtGuhd0c8zJz+8w2Ze71Rb7aBhE7j06TKWXHbw9XETzNVK3zm
73aB3Z748sSqvgRJ42akntWPr6TTKbgiEod9C+C5mH6ga19VPBLPMtJ3ET+DPOh8lBwrUzPG3sA3
4/mWhhjfzTtC/bTzzkBmGa8j7vgEWbEuzA9RnXK2lnNdKVoDi2i2jgAYHgwNGNNi2sbJ/18TYWr/
7GEyNQ6RHP0uISQ+igoSNcBHYi73El7IE3LjjaWXzAOnXjx90BTi8hy/sszti1nsxkLjqMgJqmen
AAbgObb/Z2xv/SNkQptmfCp9hwYqqscoe0L5W8qJZRLBPP3LykO6WrvvUhUYY+K83WoLpE+YXGWc
w/lBk/HXaGRVvb8vaY203iYKicGaMZJ+ix2lTE6XU/R58xyAnfoW3kTmjCdIa90reTC0ECpiNx7X
GbYiCrv0nC+4+xOBIg02aMTiQ1o//YnS03K+YqC/4UBPtniDw1zorpWZLN5k1SE+oTxPWotU9QRe
EyTB0De3AHjj3jwZj4D5fTBad6G3MBL7toEG8XPDM/CCVprdfzyWUcWEw+QDEG0B5uzlRl2PVXgH
1freeElmw7zmN4or1pFBfqY4XLS9bZYfOrmdhN3SHP8naDBoLHbcecEpzTwLg9GTflq+Rw4fiD1g
NFdCQtEsm4aL5l8W2XzX9dOV+qJG5ixFOPCUE+or/s0OvTXNRYN4hP6uBV4nPclbAEtC/WQfdi6W
zeadI4EKXLgWZbWYBJohFRqgQrA73Hs5Ta4fxyPr4qkiB4gYJWVQjVSbkRA3d39hPZC9Fnz2d5qs
bUxsPDGZ8FcJF4+gDC7x9Cwd/Rn22MPiyorGmo7rliEqx8GZ1eBC+83HJlQzkUt+U4HjC0I6u261
Tg4ulR94LBf0WT5xs0/hCfCETwFxCi0qWZM3fp5/hpHjvQCx8aDncgMff2ZBAois5Yr9WKIIhEJm
Cdji0HHtQ9P+4msgMhqpYdtPrC0qKcICNtq9iZncyJJGyJEBvmG5AAYZigBMecHAeDx77IUqhfMK
OS1jr9poFJWimwyGeGaE+CroBPPNeguSWCGYDYdYP03zEauqp+wnQu//gC4xux2UlTSBONAdSaLf
Asy7RgtFHbiD5/HctRzjxcmi/jK/pu1Jyh3q2VNqxN164tC+FLv631WdxJKZVQ7yRNAnPg3mE+0W
2hLk7cex1+me8ElV4UsOUvlVcJ+wrPnbb3IKpgo9/ejXOHwNWuvucRzyoXUCQMHOZ5ghQ1WyQrhs
1SPR4nOz63CJeOqHt9FwkCjUcxzpU7EKfLBRoROFBy/aTd3vm33Rz4kYjzVhLWkhU29nbrMGFkRQ
MmQHaoxMDx4RdKZHv8PSAJrJXU9fURq4XYTGgk5EUGEHoTm34vyyt3cUN8HakrmV3K70rSqjW36/
oothcBFNCI8JLENmnUT+ruch3a9AJ8OnQGe1E/IoBx6exJ81/lLJJxJZVewQCZmKO42QU4PrPJHA
I0dP25maqmTJaFwbPDMna2j9olk53tYvENJ5X+9B4Vc0EAqChA1ZBlrj2LTcZXCi28KSmG9mEeCK
1uaDZ/HK6zNXh494nMwq8i8vOVxlrWeETWDfFxpgvODAKa1833k5lmjL4Pwj5Zho8qmwpQVFT/d7
040Dg/SMEX7hQjYKxNnVtqtKCwdkNY0AMwVQGvHmBjVzb2qa2rRQyAfZiyKY6iGLqSX1lho21tLQ
fUyBnE+2R4Y2GytGCdCdiATTCEJu9PlWwRi2F/UpQO6/jRXA5zB7wq2aft+AGUxpF4GiTNJI1UXO
pmqn1e863YamA/GriH4aJLKCgQl/PB+2VJJITIQXrPLg2asQIq0j+SHAebEFneUXgoRcJ7efJPpp
PNz2oxEexNm8QxOC7BsQ5VKYieWiYFvc1QZyD5O9h+9is3SpecG0Rg7tdUByqFGk/y3vtzKpnsZ/
nfUqgWxDrl4GYAO5tijrq1oz6K7PuWYd/XZY6vp070ubXsrw+XzF/Zl8wwtlcecrR9KOFE2Vznxo
dkw/IRJdvwYN5qh9lU1NtwttD2gLaQRMzpFpfkHafgUKsgQVHTTSUqjntOsf6QquEfJX+23T9/yE
91UijtgN2W6Tna/QhB8Lh7CF2zcEFb9fcmO3Rv5A0+ASFDJsGVnIFdKDJIpqIPsT3XWN+D851U5R
LOZh4gnOqroWg2Pg3EAQAP/tB3LtEsf9P/Tt7WkB2HQ7AfO2zckBgc6ps3lV3wlIi7G/orPgIfKc
bV1ByxrXVN0kkSjeHNUAbG5rZzZiWjZBfKUm9P1hVgsQO9i+evumLuYDDB0fHhN4QWPcy0d0lAXm
gN1oB6y9xQJNY2Dmf4AenY0qecQocbSL19RyorFfQ5qFs6u3ZQAGBPZEUNGQ0bImIxKf9QkDm6uo
j+jC8C0VMVqCu1C99zYvfHwZF6G2WuASjtSMY6NW+AQ1SIjHAKx+GXpovOBPuOfc8GJvGfEkFeLY
x/jJcIEKdIoXKthSTbYKNjszAsuTVUjo7bUPzbZgi7BDSiendWRo6PjtwyaJ0AykzNvmVAEPdLyV
CedR9vRLbvt0egzB3YPYLGX0qls4yozH+Olgq6ojFjZMSd2uiKEBdoSIPAvUmtyAd/YkN4FTlnMT
1DhMmS77HTGCP2+kLvE71XFU/C1EmY0DE+piMFGkktAZ9H7eHZAAciUtmlZah1vek+Ps1Hpa+b6l
li0nSOs4Hvx7RosRQxDbZaShFBRJPwlnA+c5+dScxZpCnESjp7MbnPK6yfBUPVK1yrjXx/gs/i7L
VRO+FGeREwfLePN1wj1/ahyJ6up1WvS15l0ShPxksMcjbzi9hMxoIhrxi/O9DREBMuQzA7cgfHrS
KxSnfTIFmQNWpK6H7AKd3Sjnp3aWoX+eNVqR+zv01t0twPyeONWdHapBd6BD9SSGVAcGOvyJTQvc
OXi/yidQwwWQcEGNeq9Kx2Qg9lhurz8MUUNoo6hH+FypI8vDEkZ60dOKi9CEiWgr/P/3rt9o5sen
qQ7lmnVSJmEITWvCOIvVPPuxvWrewib7sc3K5SuhSHKaiMdMFjTTRhIrMSaBRV2abthtQ3W633v2
AH3JgDHJmTAzpllA4KAuWGVh6Gy3O6eAaCAscMeOsaGLqgW/ctkWQcG446z5X2X++fxaHthZJnr/
gYJl4PFiyXFzH/bl7PQwBp9GC/wNg0fEzF/OZrc53CGMp8JSnjw3zfiyqCmtxCXTCJITo3tKY53p
RRp7xtOyG0E4zPuzYAMHuM9mssSqB+Gj20VdKVMLsBuJlJyvgVdh7oSdD20uu79T6nECiEzLIdyh
LOzqgnPMcPlNF7btUvTV4bCDe6xy9UUEin72Y7PeZdPZzy3fPxgctlMyx23tatyrM5P214iWP6bu
SR2aWvq8ABE87mkgyEKsViRrz77fd4GlPOgZqO6BtwoXDi1bRNOLMO9oOPC7RAfXzhhLwC2JDnOM
xzglVJy33P6r00zOGv3piuH45vVYWs8CysKnjKlGMiSNtfX+fq2ZezPc38ch1ozeRQA3oD/ZRBaz
QfYG44RoQQsUHMlRlaeKnYYx7eoxP0KMyWHaLJ1Cd8TRx6cV8bm/VcFUOanO/jmHUwvKhGMn+6ZF
IsV42JNf7vQlqCborIPL4SnVNNB/Jpw0m7iHiT7zze3WhvRQPYVc0CCwtxytKm2xU3hvdHt2VWV4
KA0Xu55ATYSU9clJrNWp9qswfxcKiR00wUs+PMUT9yS+MFmU8RQ+6VAdXAa6UJUWyXNJ0fCRjNDf
1C2OcgRaY+mvnlM/NUbeixFK4zZj1k70aWOZBeDW7Zj515lA/F+PVkjr/3SZ/lz6Q4RmNHXKmJOy
5btXbTnLWzvOT4D0uBTAdGe0/Qdj8fEzPwixsKAlTX1YAXtz3kwbg6BmyKw2e02Qw9eTzhmquL1E
O/6qjJXxBQ+50XhAeF30DZ3+neOGYEP3mtRHCNVfnIxMK8ixbrgTtTS0kWkkBlZwMNsr+TLqhJBx
K1dnS8u/XTRgvfsYZEuwu0WkbpEYRFcMUqj1U7xdaYgcb8hZPjpZ3F+YBnZQHuVuJroddLqwjWKC
fIag1QAwP+JjDMO1/vBdR3b+UYgclSBXhgqDZLKKERM/s4X2i1bVZvX6irq1mGEb+n/nH30UU85C
krmS+39p3yCFdZduaZDwwmj2j6R49XJleIVfmt/VX0cTVp6/sD3viP2eNRrh7AUA+6E+85ZKAA6f
7qJj6YQyYUrpvReg/lmZg4XqS7+R7jdMV8CGRxMQrNnlwCozgMQSLuzVDKs19NjbT3stXGUpAZIR
ZopnnxkJhscQ4CF9kJGGPesw73rqYfGDd01u+qMJrsr3YffGQgcEejJRkum/coh4NAQpatosRAwF
1vfjYsYjQh+LwUcfBy37AVSmzA7dXhxMLGj3g+cZtiU2MnWOAheYRWQK6I7corcHt8SGEKaCPqrj
XowzHCGln6HWTX4UlMUY0I9rLPZ2lqGwWrA8peN5uboWSuy6i2rvDE30pIGeUhOfdC0grGxImPlD
Ui7FQpU246KmdHK7nc3etZt+sFLORqsTlapQij+JU8p3NEq/2DfBRJ9VfPLycjzBf9IZWLXbuuJ0
ONbjcrAJd+MPOD/wVq4qiGtIPkRF4o3Wncp90KDKZSg4v/Kfmd7fzN0g9wCj2Px32tCfUqwLW20R
6i5/mbtc4ZkrHbW5cpFcxvnIa8hIEo8oLlkc9q1gdbRtXnzqsBrPDnpKBQgEqXAwhsP/fVvX5xDH
dum9V1RL1NYFUzL+8L2urZ44JCB9Wx4yBZ5h1/52CGFUM6b9jXDkPZ98bBVxQ4D4a5qHADJtPBQy
aDqQCVag5m5mtkzlV6Nnr3Qov833joyeFUtHXaOO+yQDZ93rtS79Xb65RqK2mpzWYOgP0jC47TKZ
8+DvZJ1fzRONDi5dovCJL312rLndTPnkOwxid+Hb/7WeV8f7oaVoePO/50+Fj4tlckiucVoU3u+j
h08YTplWxBkEfdIqaT9VE0oDnjY4/TeMFqdqEGcRhHZVX02U4yLdCoEYAjz9R3p7i5mPRv6pRQ2x
wJYMrWOjErNSczRYaPeXP+OR/ZdBnaAKYYdCac+T75tM+IKLQam/DaZ9Du/RGQ//RN6c+Y7YnsSW
xm8bZW7Ab9eEjkFOMu8psO0+abqXpZ2KR9BjGdZZx2HKvVwGDiVGrQdg8iOASv14XWlTaGj4IylZ
S/PSJovo1Fsg8H2BTYt9EPydYIgR9w70H9l8jlSJkUrYsSZtaI0R0D09hPNStjqh44uBZvtPPimR
p4syFDfCtoqkx7TQrjqp3v9LRr3KseWjNujDBp3yqJ4lPO2klLd2WL57uAhfa7+FocKQxZJzD4kL
hGg/1opklO63CaPv7x8+9YGvhBzi0YAgzkCEQQ6UwW7efj/S+o9y/9Gfu1LJdkO9Hik1DcWFiKw1
cTx2FxQ7B93Eu/6cKa72S7KfrjapxKvM1anzgauaaoo5l3JfYKtb7idEQqBGifQYIZ8dE9v/+3db
rzrY73jYba+RCWbS9hQXI+ExMpcX08ef1WNqCP+FuYbJqY/2nr3T3q0XC1MR31+3EyPG0yMG09h1
7MwLdURPxsuh/adENOiAJA+LzL/SrcgiCVekZV66BmVXaHo2YfEpoQxPA7YYC0sbDlJnZ/YVj0TN
pTZAldgkjx5qwlW+FhwsfSs3soqsH3AjrJU7THRGkA3k4rBbw5wl6sEXUkVUyBYgIEmo7NcbnS0T
GuWwPT2aLJLtufWddQy1YgigUucX23bwouUZdBMp5v2CvxaoahUFE/RZXSdHos+yFiKg8N5JjVLk
Mai3KcUNHvBp5B97uwF3FQzn0McWxH5YAE4U7J2sYqjV4Fhdud0j+z1BTBecmD9mSUIL9WjVch9U
kz1ZqOpi3luvaecCtPU2MacwmjfVN9fO2oCoau2W/Uyo9BIgXklCkV7ZVnbefSs4Y1mNOIbIRRh9
hnl3p33E/04HjymPcfuxxz2jJ71jkTvvYV9GkXCRdE3JbxvMMOQXHNTUZdimknYvekv+Jg/H+t7s
s+aO9NHBGvm+alQUbNV/d7vfprCvOf/fBtzDt2l+DNEGAQCr2Ixw8vaJgeRgbesw+vVmvxPSXTLt
WHCydgK8vrKufHOlPei4h83SMyEyiBi1xv02sGTRLrMde8GyQIMgW5MSpJx6Osn/1i5UgTR+3WRC
e/SQKivPgbIwLNtWcdauTF4HgimJNeovCJ1KY4rKVqI5f/1eq1GYXEMNKDbZoRNZ1URDAFWTY2rM
qqWSEUXgQ1BRfw7g9rKgTYb6mxIvER+9rBe9rZalCL6m7twxpH0eTGdOh3r4830SLVUPqwMH2cU5
xRhSrK8BJz0tJcvypK+of+ALWr1wy4nJxkKNVxvX1G+pfZRyxzRi49InTcSQNc+1KEYJqfTbtN/l
04rGPCOpf3GE2m7c9g9UgKfN6OzM7siJ0UWDtn9GMZAOfWZKLWgwX5HdzMTcBGXLUZ3Ar52T8hrV
Vn2qh+iQw6ff5Bexq+6G5xjPY94UqP7bNQ8Lf1qLheWjzCeC/hV2J4oixatgJC0zBXqPeMGHjwOh
eqUp6oPmeTciJ+hRGMxQf0B0tTVXkz6T6RVEyAqWi6BZ8ObsaBM9IXiPJpbnmuY5mUL03s3qeykd
emV2E/DStVAAwTmWj4hdODz9O6O1/eExuOgMrk78qeGVONPt8FbiWDUybqyvkqKDckUWgbUT8oMm
Sg2rZLorXa3Udoi6dQPBfAAZsygkPBkOJsTEBFE9jhT/30qAx0xX7J/2PXHz2dEKQFuMD2VfviI6
/M499hkGvNPohAUiuEv7uyTID7mM3GtB+wHUfoBi2WGOINkTWoLVzR6WOnIFAkNfSk2zEpIJj4Xi
JMu1D0lXPGPSQUe68+Vf6MNBEr2mvfDjMuwwr2QYhwpimEkGWtLSP5t+4kmBpFMe8yjwYT+dwnTy
LhDsjzU2LuLOEiQnfSzyMa1kXz3MGYEsIbbtRK/SIahK+cFzT8Pjf63sxSG1i1wLZnWwVBwEA4uC
9TMlQNX90X22GPSULZxO3oS2TNE2hoBn+gE4yTyhPT/MSrEWAvgCViSSykukbeb5ELOb6W88GYfw
FBgJ7ZWHdul9W7/w2GdNmw0vkt768CtgGyVlu6kTnD7Xkm+qMuKcOu/C3len/oVw1IwX+QWWQ/45
CN4oZGKa/75z7LceQXRYdnTPj1dDJCXpwgyAAU87v82lbv+ukkQVDcJYA9LWB9PwIBClcD9Wbeqf
ZeyTw+MPvy4dB4dfEoBggR1Nn2v4qWcogmU3mUQq0G1JX0iLLuX9J0eSaE3auAT/a0hbTQeE4CLH
RxTZlHzMDhbL43nbfm5wYEIiGg9NZmhKNrO4VcgpeKLaw22itDoc2lKvkTJWvwnPGCIBGP8Q4JAS
yYhox7nHoU0gLXfBHFHBUlABv1BScPX8TXrjHG0O+Y3+uTlu36Vc0sWBinFHBWJaOh9Lsif6F6TD
o9YL0G4f04DPJI/Cg9zpT4cCs9Ub4O8LOYAv8GXtXCh9mitOeBg1LbyngqxMkMyhOCWJYgNSK/pF
0s3OtfvqTQQeIYqo9SQk5r5SZCpG61Q69mAgqrJiT89oBvZ40FSEbtGZptZPjYpL0/g9pE1qbP6Y
4+a4YOhaFVisX5F9DxbnR9pRngeJJCpneY2ApVa4xDEbfDN+g7TqpTEAHPc1N+pG/eS0euC6iaYU
kamPErn5h9U6+O4WYKNUD3wc+jWqumyxN7L4Rx/QK4s/ZspnPL9yXgwRVV33qwZYtuGCsCvjPma7
X6inU9FrO3Ke/v3XwTdo8WR8XTpsDqBEMiyAWRkd2KNIUaNsSsY6JcA3I1W35iWQzpmsZ//zMKjs
vDty6o426gRAiGAZFoD8kTN8fbtlM6UOGGN2Svwbi4374F6FcxPWwpYpz/AwvXKCINgdKLG+v5is
pAWbkaRz2U7zYoFiV74lHRXZUKnzSTA1t6YNy7AdPIMh6GlhnsXBA17+XobLRpgR3Ky1ZFgDk1CQ
m9MNf+XcyrTiHgVVKced2ajSlJ4LhZFK8WuN++cdCvNbTj5nDd94dy2ytk7eaoCFyS/QOjrWIoJI
vHPo6qAQNw+nraZ+DLe99ELEOfW+ncORp9GEzzWJT1lmmUVdj/DBlBSc+D1sgvE5lLXmcCl1xNqd
DDueQjHgJdWhuodK2g+52eJ6IASfl8kAjhEd5qxETjjIP0BHSoperJZwJvhwrLtCkEODY9Sv4ycz
ibfUXx4BVDfcasJnBrq59z/BCwFOy2l5lGhujJ+kOUYxmVtBmV0IXjjUuQvcXtmJ1xAJ6CC+JNQz
n/5LeU98jg3mGSeh2w4Kzq4wnBVxi7ve0KPuT0qgLPNd/SuOsOm16+o1J/Ba7tdxkumJrBDfICkL
YhjxmSo3i4JGeXZ455JvekejWR4LhaPWRCgJjjRcLzUfOsFIkMToLxNRowcDXEuTYwM05lqr7W1x
itjsbZtafx+kRxi1x4d36royptCAR9AXUjXOA4Ta83xKdN6UEYmGgUWlQ+pAnt4/TF+NBiO08cne
KNGrSTvWZFZ7yk3wcwm3aVaYHG8T6gmyXO4XJuXWw2hpQPnieQY2hd0TBJF6NyAHjO9EvNk6WsVM
PdUtpLF/cy8j4eB6H8Zw0nyDlwlvwv1p1SEUqMM6KVEzSpNwdBQjg1AUqVSMoiwKw7pClfRD54tT
mH6kXeYe8HIWl7o+giTXRCGJd1ufXIeOepuQ2puycvlAlSjVqlviVW0d5ommoQfT9IsL7Lq/3LLS
WSobuAGtzlA5kdSb0ON5KmWoXr8JxOcCe5357OQb00Il6E2SbJX2OhfyeaHXhD9JEfsoBiOcyJM6
VAmvcclc7CSGNeFXWv+SnvqyeUK+mtTVmc8ZvSat/5NVqIhWM6wNyikbQevUpiMZm8kVbTieG6LE
9DBeHeK4ns9fYUrOfc0Bo0abZPx9CnWisPtRE0Tmas4YKSxTjXNu1h6Nw8hwy9NXkEXZrqO9CIog
7c6g0C0zsFbbA4NYpDktVzL3pDil6T9mKEHM2T1OMPL1Uzl4Yc+CL0F3qPcNsc27MfzgWj3HxorE
b7XW+LKzsppHq+eMVNjb0hZQMfRSWMDZgQUXAPghZMG2Bz7PovpZYXCQ+MzNUzblQBiuqQGxv7aI
PtRSZK3PuTiuHAVCTv4mXeZhNm4cDhSJ2P+hdnCeX8LWjRS2A/Vg5OEqrSg4N/5h3T2PE8uai8WH
HdfBl8XVnqgxv5YdO17sufUr+aQJAQIy4WdFZwdqPtFyP9hTqL5hsplHvaZcOQ0QlBAvy8+7Ga8X
ddKZdBBEzK0Y3eUH2vKZsZyW2dfdTskPqSJQDUXKBTLk0DB0f4j7YUPtItN+NH8gIFyQd32/6aYb
dB7bWXHu0SJ6eZD2dDCZf1/pM9rQfUr7trR8k6Ln7KMNe8+AtytmJhQbLU6Ki80a5QQC4f+kLIQp
azMBF9xv79CyLtZjlPmE3JiOuQmQujo4USn71cOJZFtGysozgDb6e5QeX7bdCyzOHiKHSihUqrnp
e6TpZZmtrUnq4sOniDUkNVEW4bHnkcBF/Kg+sAq49oqvjO3mc/xoLsSrf1WpnJo9B12CHcIdRZKz
ieowaZwPHgMKhJaJIPQDHSmvTBb95VxnA0+dSWTuf20VBPIrwdaCiQrOtXaec6dyJ1QcVfs8s4f8
lolNr1GkN/917uwRRXEHRfrEO3vkG/cUNlIkaDJEU0rU8qS7qeksX7OQC9c4OObPEbd6vPtASHqZ
r+4ShQH7QwEkNccpl4dkeBngVHM2chbKyxCFJAbIC888J0/Bi3Xp3yzs8AKjtN+T4F8RE4L/IYjc
xkwOTri67SY5uZB/+3NiEJpdcSF07Lxx7FFyVrS797b009rZRbZPvT62nYGx0XFqRIRI7UYuJx/q
fwq7RmsmLeR55JVbXZmGHYL0O7SahJ3LnIQcVzI5cSYoyxc6j4Y7AID9KN6IkFgDKT25zkjXTUgV
yOoBrB2vv/wvzaUtlktRNRY/5U/gbMLxDgyjDWqbLqyrmUqdFGOB8FfwEBeFEWStesuZ+MjXW5ra
88Lpu8tEk2xNa98lqDkKbOfiQyLtCUwNDE1QcqOwvY90O4StuGOfQKMfom5hRbNYR4BuJh/k6oxS
d9Q5664hH5rIDYV9zP7pciVG9CHrwe+ZKew4O+FQ9SsdDGAYoUvzUma9cUvA95eJsxQ+7HmIFzQy
/xnMVlMW6Csoc/y1ZlbOaoO2+lch7TosFdn4ZbmwQ9wj1DJti4uBZ0MshgV9qjgUFR0ylm0jpx4F
BxpebQgVXTo3GCLdBYf96XHBHs303yT2qardv1utC7JnOJfFe2qzliTyPCNGBeWn/rZH90m9A1Rg
TjPKj2hKHQE/H87N6ywAXkHx9xeqQRv+GzzSKnfspWa5ehaOFaYsHahaRd7K1LTepXPsUx9edCNb
LT7jjYQd3Jyz0pLJnCaP5epsw6165VyQKzGgKZdNM/eB5lLFNilLZo0a/cRM0Gs96xOG7xXVAJ9X
1eZFMibme52FxRJDqoM7XVbV4X6Mt48rOx/guNLNtDyhkw9dLVQk1TIJsyRNaWYLH8uKz0qVGAkP
o8aE+AHLWgv9ranPz4JV/7FB8bSD/7YZzVg9S0WNrv6q5eaWWFiUk02ZwR/zkEvs2QulHsEQuhee
vqAIXdHp9MGW8TUFG9lDaAFiSaxBRt/bIPPdWMCOhfT8UdWq6AVJLO3IpeeiT1RWkozZNZipJUW8
WmqhngY2iMHPF4yhftgjISQG7xrCoXrJTkKB3rD2IWIWAXJbtnBlGSCxt/YCSNvBO+K918ZHY9k6
9vDUvY9OSjwBjtxqLp6dr0BlB2O2U6Hv25uAWdGldbAytPRyDjwxzo/iwWJUPNt5IuDkqT6H2P28
KMikGAxkRk52SVnbjR0veWBkBySOhg1YQlEzpppOcBRmrITFr473cblQuvQiP1+XyIFKj/CHncb8
PnSst9c6xbmkE/MVEzlFzOb6kiy51ZdDzQJDNSxgeRGyS3rXZD8jtq++fw5riWZRmB8ydvh+Zn/t
6cI8N1OV3LWgb1CY+ub4U5Z+F/AEN2Sw1HBzc79+jIUtsedkvUlRl06FLrU4g/HH97r9oybnEev6
61yyBT+OWVCizjQxWWLXwQ6AuzwpmWsGoN4nudQqq4OVUThHFk8pKuEoZuOEWhRXnItvr6YVh0VQ
7l4nRCf2E7W8Shw8RLnA0qJrKjhLerwx/KX/ILMLSwP0eGbO1UxVsenGQlYyxbMK+rrZ++mLPsFG
sDMAmtmMgXQ0Dpvzs/SseBVYnBIwg+VV7J3ANqrgP7tOxb72lnXz8XH3+YvkRE3uhW/fe1QXAE3i
TeuPl7MNgV2I2vy5amgVl0Y8SK55BJuf8DX/dREkIROhx49XjmuV4baJUmH0gsR7GSTAqKMPetaP
pCru3RBWC3Drxj6LmkVxYYPFMjabonIXbyP3S561A/6kJEzDOmSFxG0lD3Yn2QHZbksDzoZajP0C
kwgxPQylLy9NC+1PpmN6XwP+A6dj5cqZNw1gdEzntpbhsNq20E68ByqzIPy1hRsoWHgvc0gAZ73k
2swEC3Sj2n8kBvlqVUOlwhNr05N7cLvjFK/LheltjNtdWYyoSoe9e5k4OBittskkLU/tGd1C+e00
Aa5x/Q+CTfInaLUnwjNJeuwm6ELVnZ2gHPXMF7AoEX+KnCif1nSqcn2jb5YELehNqrJk1Mds9Ew/
WZpWQS2K3kPcNQzJexvlYmeHe+3TE+LJSP4ne0t/uDgq9na9PIlRsZau95wBJAEUDRj20qQ4EfM8
xYrWNZPFExfyT6Bt0xhR9GPYnDKAaGcymJbJ4cO+aNwiDOZq+ItUyMs6K0Vi/fQl3S17q6aURiLT
73/yaqMwMcva06d2K0juETqemw0crGVovkXITLLbPxSJk0njbzbGoqaN40CPjZCVPRXTjYZPhFhT
IZdQVGMw9oQAnhmiu4Vxb4gOCaJV7jlF8RpLYLsVrBhr+oXwPv0tPmAEwn39TGkmCb+ZfH9h2CII
+XqS8Il20y8HugsEQvA0HYAGYPPKSJ/NsTCL5eypVvzoMz66jb0D5qFBcOimFYzFWW8BVIoD5AgK
VuIFyRGbswwkxbKCC6KK2qTUeP/7R4/ICr1pE62cLr/xyRaCU6B3amKpfiPCjaqbpQOgwra/9Bjl
/n5xp63QLTltVMWjV/RrIEkE61rbANmJ6gCp59xPTFL4aTeYs4dQ9R7upXo6ivKY7mUotUFOMJkB
qP4ddSMOPa2ACQQYG/P/Or4UGyVC2UidP/nso1x/i6hxaDBTlWzVbx5AkmaWdCcLQ5r0Lvn4C9uE
B4ojcPpOMh2lyxfSJbfpXDF7ZDmMprj3cruDHlVqLnpC3iTs4/P3eB4599vT5Wq4T9088x3LtQEn
+CGOt/wbGO77vEW+FvYOqpM8AbikvKARzGgXVoJ8eImoM1ns0Ly+rXdytmUrMn6fiJ0kAnGtyqyJ
5CHKv59k34ChRE8OFzHXgoqWj6tBJOA8rwCbP41GuDFoJqWBbF66jXDEvebpLamB5F3BgK1H2XZN
qZq4UO2Vjx3VIze+vCQWcpPiPFGzLZWnz6pEGmEGPVNnAzjuo/KfD2rNBR9yCaNb/u3o9NxurSBr
oRbO8dpV9SNcBtECob/hTG4YuIfzjT5GjMLbVRkwK6Y99jkG2L/gbXGIhtjFNeGFCQzaFsJdBoGM
h5F5jxzLccCbNt36mWrNidhGxhyKdH4P4WhQdonAmfVJoIGxg/fmL8jP041vBDT3RTK18vlZQvFo
4qLJ0QphVRq11hksXfD2ul/83TBAcrBTUQsT14MVLzfvNWWlMeVUHj5w0DoJXp5fy+dD1UfbHwom
AGGM0yuzfnBgBT7UVQEb/XCpKXky5MexTOPmBDQWUxdxEtXrnbqJUJ6nWRB7EYtnsaZxGHvUopp4
+V5OMGZ3s1DvcvK0Q6psA1tA6qLDWPP44OXxOvhttnqKZTuP81zOU6BEAs6YwXRAnGSNtPsfM9aL
S0DV+skbmeb0RGTPINoVeaAWsvTaI//wh27/nUhnEPRLpkicewAlGiwG2xvkG9pRuwP8VstEknhU
VZQSRaogr7btYk/Q6Yt+qzrW7ljbu63gB4ZHQG2XqKWFXkIEEan8u8Ml0UKleAvN6RXgzLLDEXVx
3eFypdcC739uZyimriTuB7CGbS6xe5YMhQNc5+1unUDJVynQDXXW5l6DUAR6oRWakG0vsFGIrqvo
SkjgbAUq/egDb8NY9trH8QhhUnJ6HiUQCWrOOTp5m6JJ46VHrQb5CvIivsnBg3sdgimNOxZDB2An
FLeDASF9TG0L1ysGJrfHgjk3RhR68omlXQ952VMJTpEOvLNeGNBvZHTl3sauiatkSnA9GNHxDhJj
RE3nlukoa0gbxgDuwUOwHTXnH12BB8SKZUujkHhAx4tt4h5Oeiwg3TIBHWsz7Cz6NWfnWMZzLLnv
YVDacNtqYJFiZ5MJONfkKpNixByldjaFjJVEkh1vsilZ3sDQK5BOXylMDCfHu+hM1uK1unKW4BMV
pPoiIhABOVF5N3RBvfxtDLLAl/CAearXm0rGv+huckMXIinGP29whl6fHbkSg0R+LRkatbpWDfgZ
X98Gc64jeID2TkcK3wHyUJkIjw1foyby6Kp/+Squxs5JPGjKC19g+e2DNJzZRykbkpfQddkhkQHP
6OTPaxWKMqd4k70kyYjbB4FM6nx9anfwi85TbEFk4sIQ74fCVR547uX17k2GqXFtkbq1TpTVHbzG
D1EbuPBwXxn1mNttNxudFXlSfcQaZNSPXLGFWus1fATBP5RCWkVEEvn3hO/jOOv//DFi/Ec9IzhO
t+XsLvwyb8wBlhYkHfd75IleYIXdR/kErsHG8Y5o4XBVyF0i1n6baFoWMSlJigFso5wqHTCN/o6x
f6KzkZZ3il4/9Gh4JFTfmuAGz1wpZ39DKAvZGM+V5GOesgVe2scDPmOt5tH5gizSnTNyeU0ySbmt
WXxu9oCqrfshi+mIDuMGRPqeM/mmuSjuprpgQ6svfwIS6YNIax4ZU+uNuj/AnZ9/b9gIFbtd9GDA
c5JRXeWJNapqjD9b9wldC3a0jVBf3jYLKO3Zp3QPyMeM2na1lEI+HuQIer+JRG1rYB+s4tTaXcLk
UZex/N3aWQw6L7pAfxmgihlZsLcamCIOZ/CcgyL1srM4jyzO3yTTFy9Yvz03y+sTmXM5YDqKcLqs
TkL3YRjbhf4lXltkApt2Szl4AI+X99WP3a781SXNANVBazcXjELROQuXQ+3iHuaUoCPf5ZoiKYjJ
kVvImo2m8c+M2ILqJfsyE96mWoWWGF5SE1+LoynSF1yVy+FY57CI6Ah9uPn7wKW2Sh7XdMUaO+SP
N2g4dIC5hjPjTUh56JOa3b1NPf+/jXO4WSxh4eOJksn50K4HYVwgttov261fHAA7DwoC48lF1S0T
UIteYK9TpHXKLZDlPKnoJbLyTEGNCtXwwGRZ75lKKneiWLkv1BhNi7/0GMctXOII6OfIvbyQnqne
ctdB39mtERAlizK0j95HT8bVCFk0OYty+pT+fUt7Wfw3yaHW2hG/iVl6HwB2KbX5pmuDajuxZUuV
KX7V49fNvkevFmm4knkwcUph13uTVmkbEwR4S/vl7WQe80M1NgoSC6hz7YExuE2Ige4i8xJWxDSK
w3RsD86L6eXAU+ylm2apaL3fKohQuK7KF6NNpnyUQYxrdTcV2Im/2MBbDltdcB7hst6jc2eYCtF/
iGX2jB2TDqXq6DP8uM7OblUSSBrJBLggvLXayyBAMeS3ZtgAkXnxAc5QtDDhvZouqRV3wJgL+zeF
LPqs0f2M8hRVC3jA1nBlI1jwnWWYa4B0JFdfB/9B5dJwMV9odKO7OS1mQ3hvOFGSazuUKE5szeSX
9eSWtEB7n0ZRh4ejunAg5/9vn0Z0bk72KZtRrud6iqI1TnaTu1DVNJ/ap2yOPfcaY016UkLm93S6
+5oSz4xFX3hbI8UMpu8WicxYyQIRFHJ+89vl4Wy6J5rz0a9xWfoXyYolSuvC09isZ8sX4AWhpdQq
HSsDjCiFEgWMxWX5Ejvir7efJyLQPDiVQJ4OkOgsXyCYKZKb8FU5zFJ6ArV+jsBjg9PPrb432nQy
h9zTmLviptFs37bqLcGQa1kLjL7Cnkg9tG0AvCpUnZ5gzKUtBw9JJXQ5+7ga2/cO+r+/oAtria7T
freBoK7/gaaKvyzxuF4+Q4OEI8nmsS3lnNAQ0vJ2OjSbNyzaLQ1xqAFg8RMMUzNIQpAjy5ZEmkDr
hoKJ0Yd7/RiAnbpQLoc1BPFrd3HdXsevxXsd98F+xrm9fGnY37hpI9H7u94zfFH3zQoTBkp4ERBS
1rDrHR+NMNUykPp3yGMbIaI47NiMg7Un8Q319k2m+or9vP5azpLjqhGhqLIutsKAwQMLuzl9d1iW
b977fkWeXJjvw95g8GYtTScOehhaXIEo9nFoyYPQWGQ8iL3QdjqEEy72KQI0k6agnYQl1aJPdKke
kcTI/xSSC2PZUy/2BgG0svzmry+FRyajcVSRYTOw/een087SSp0LSuVJGouwxaVdzsszOi4p6YJl
wuH9fldwDbOnaKpJ2MUkRrFCGJO9NhOT2vW/hvggPKVrMdEjet3zF/uI5La8k72VKmXmYBpEcfnF
oK4nDdDT0uFsekp3DqGKEY+H16Vq1zUif/GnTobAKVazf+wcP5ucmZa2tBLnwS346bqtkDipKx/s
zxCQ4+SAnOBQyzIBVyC7TFl+4/X526s2sr2imMMHC5CS8TW9d8Om3eNEIpTizJwZqMaJ9jzHRcpT
8Aa1cJHkVpMDXSw+dIGF7iZ+WklIkre7CG37jxCNKZZUhdWkQ8ipYVpkZ6SWareXCmrsS7R9bR3w
DvH2ycRRpPIoSp5QO42/VpQPIJrXcpF0lNpk/yL6tkqOxUvrMTuATQo6uGF2LlEOVl3cpC3ktyIt
fjkaGKM5nm0gEwUh2xzbql6j3u5IBlOOBXhI2XSUqJPcUbvLAOh68sIhxZRKc/iNsUVqi6EtAdi4
ODai5VOT05Okzz9tsuYfsBz8YXXJKPUiqn0GioQ550PhNSZV12BbkBNth6HxVAEaSQ2ionzQXBiF
PSi4hD8d/pillEqYaReVkKIIddsuf4ZIRI+3D5p4HGWZNquodlgD5Jm1agOsHHOTGz08U07W5Ntc
BPVNQKjH2PdZ4VkqvVyHNKr00murDSxn07I58Ega3hYbQWzC9KHkxV1aIUVlR7VJzeQU3YB6xQRA
3xc9sOiegReLdgAXbxZKWUeZbC/w002rhqLUYmAfV4tNgAcAaiRpPtCsy0t/d+1ZTyk6m7Yu2aPw
P7lLkkln7loH2+15KPSiPwowztq+JsgNIeryNws91fbyriOG37y/SQhjjGGxiq2hpLc32niZ9U6u
ezeN6x1uuoJaTK7+urN66UiEjoIJJVLn0kc4pM+jI1eVsLrbeG/92pQ3HuUJXjuLllHlSOgAP+1K
YgmJruz4Uq6TWBM05bddjpMwCtfPVT+LC5sM9QVVmw+pn11YK3Tw3jbpKVN3n5o7exfVZK9mDgHT
FIBjZflIt4CEWqCr4yzMIYe9h425WuN7Iz5/t1K2yywQsMDvOD2Jb8rCOA+Lgi8UzoulL4y3aesM
d2nRHKmcgqMDorYzvtSGKKrmCmO3sy3fWErzv8awLf2AehS7WskDAC129BZoFBOmhCCtYFPXuW2X
Z0/kFbngn5VuhoAcJCODN0EnBHdEGGu9+LNobyYWwZDDfiCoVdEpqhElk96fJ24GU4A0ZcgBxMMs
ARBAaGYUT/Fh6SEmFr5t14moLw+v6OJmQDYnhv02D+MNyCD85cXtKoT5S5Jq+c9PjWQXwXKKyf7F
c1k0Ph8hIoFr4SNO6lwa3lfYa/EtvX5Lv7kvkIHONq3LlpeyBom2FJYtnmhCYIJ48/AqOpZ9vaFq
4WLgjAYolB1MLddTPlmTYc0iYYAesc3u1DAHMnJfHrKWJ8hC2e/gf6Yxk25KkZST+0lkQjKCf33+
oCa4HyRGfs54au+w8V/MGrgL5+yz9T4OitSOXnURRJlVwJTdWJ/wOZimNf9hwaHyCCJ/aiz6m5CD
Jc/QvDLI+l5jhByOSNheQ0FBMgLz/7KRvA7v2xNOaUVmEtAoLeg5PZ+9hOVKe15j0rJUa4nZFQUL
EcXSLq8+RIjH8W2/pN3zsSdB+l2TX8RbZEQ0SKoyKFeAUNcOSY3r+DP0Sx9nHsC6i3WhtvsMdtH8
iywlRWlsqULCy88BySTVIwmZne+rVvXlceggtjbGUq+nVF7ng7NJLkgaTH1NUjXQF/4Ut1dYpK+T
dZC1igQ0NhGdw/3Qg0zAwtyJkdtVTihygVO0slL9kZQpGeDamw/y/x8nujcj2yE2FuI/pUk3kZyh
6Y4AYrihXLbateTKLodRJFn7iWYj+4PdO8qxKfZBkq+oFcoiEUISTI7Rm2gjMiQVSqHXEV/gKuXs
pt1RnMdv39tW39rQc7ViwoOYJ8FsuQrKz4xfF288WT3YSi1t+fCr435hA/I9usg+z4aI9hhu7Ohg
s1ky/qzfqi4czW4DvqxmmqKRvHMAH+tGx5I/5wx1/aUQF+A1s3m+my31tHWPjGxApvV4f054VZpP
I8lKZSLc09Yq/lGAhiC7YqfxsWAgEdJ2qlONQq+Cn/DPYEIBXqPUNIWkX7ShsRV5CwWeKertkt++
0Z5yg8D57EfiGxUaPOvpCuFFbZc2AioLNf2uaTTxmS7/E63tCkfRp17wSpdnFKkQejkW0e18bjES
0gfs6A/OveArnr2S9HMvGKST6ZVMagKXSZsPslnrSHMh59O4jL8szwVRyHRKH5K6CzyQJYuOBMQZ
oRWkbQj49ye/0paiGZHHamqxBa19ijnHGHqE3k3xKzpGxgxgwH+XAfZD7vuFiRQGZVy6CFbrDo5y
WPoobA+jQqZxBONcwaz7Rvdg51K7/kTfID99SZHwhsVgGsPtyiTyW2gK7PTxvz3NYaGPbdq3hUN6
KOj2DkA9sIPOnls5O/c41HclW4Kgpu+XlXrf824DkAQ7HU55eqh9aBRCtVoq3YdGXfhygceJ6f9l
6da2e2poKbxsT6/dOKK2XafAKjrRuk8NxtOD8GwJ90rwv76gV/aeBkrMpcEMLyT0bG0pY9gcRdc+
FNOcvQICoU14MOyuTySkekPKqBA/Q9IhsxSmbht7nOkbZcYKStaTbs0wIseX1CCBebOmzdJHko8t
rLK8VYyBwhAdDKZ5tnHB0G8RLAqc4JL44c93XRoDR/Oqq44xgjvPnevRGyWjuk0O+/EZaLxJ7f3g
1GWOzL01VNpatJHvzHJlExpUFuhOflW/CYEuxBUBQE9RSMY81kndSz01kFyEm5PrIIlmvRWnpccT
EggpA0SDViqhjXOC7uFJ6dV48q/dQv3Iu8HjyhnBiinDrftF7C9ifgdmM6Etc/SfuHOBvd6AnMKd
5WLyUtqUTIjtPtRV3LVAsRI150xmAXkH7hSjTxeUa19vB7Tnvo7UrTnt31NA7rXNrGcKK4piT9Gc
LyojwGGORdXNBB6jG4x9qsOy9nhEIfczse/ExxK8Ef2dY21bxiRQ2FXmzeFb8k0inemyv0VRU+KW
wm2K+f0UKa0AUtFhNitCKqlYuKwfwjPmAqUjWH2t9+A704HisWwEA0YxuZ5Br2CN43Hw6kNzHtIO
V3/HDhrFWYPl+Lb6z0K9cBE4WpgufH99ysr6lGvBjtoIe154ATfv7rhMXhgR//tpzpdCC7lSWbEB
CEITPhqE8g3ekg1RAr8jSAIR9L7dM8Pjq9DqHmIMDI2DhFEZ6rjQLRwiGa4W1nUvmmkE+86vaNtZ
pIsR04MGpPkTuAy2GnnuUxoLFdyq/5rto+hwC62Q/TYR5rlmwlJfPfgLbfXbuAuceACwvgFnfQ96
hVHglqGDL8Jbva+PBfZnmRwaBtHP+GKBdVxznz8bXPd+8U4fwbuyLMXuGQdoFEzh48zHe+N15w13
iE9F/W7JKEvn5gfvQyAFeDaTXduwcBzPSauiUUr8SNLq8f1LnBdfR5nZ5igpfRI2trUDoHsMeuj+
P4slV3NKVxyqMm38qI+eOUwXSok2jTVyw3mVZaoRqcJ8bXpQaEjhIOy3TZFDhqXuges+ohWh0bot
b+W3EGTSEzOpVpN7ZJYQBzTz08LUxeIQ6dCqBQRqpk5Y/+sYqKjYVvb30gRLUXdT29JQ4AUjaUkR
FW7FDyDGyJ3SSq6YxIUxZ2XzjgS+qmz438ORfJUcr+Q7Xp08y1QxPJ9HCGpPWN2TOmUVOnfF1Ph5
CPBGIeIQwIKZcTO9Gvd2Sh9NvUGXoEiGN4YO6eLuLQMAf+Q1iKrZfWNlFOD08W2mnxeszu9oAF8c
4ESUU6TSA39+X8u1P5svaRi/gJ+AkggRvGwNq1XiMCLm37KbsZzVanssCWbaQ9WeVnzohg874dCt
7NgbvZqQkn603dDHJZnmNf9E/k8iTs/0NEXgyhWEklLfWl9NpCBhfva8892ugjOcCpOrcTgxWbBN
xDaPDiQtfUb+Th2pnteNJUCAK8LmQHc8j+kY+sS2OPCUuLq8viWAIFZ/f5ZxLfNTV449ph2soGxc
ypiw4XPvjfpqwt7CvQVIvwctvaLBIIrw/6IdWnnaVsfhdU4tA0imU4k83p2ZL5icpADpYCktOuwK
xHqe2mcJB7KQ+BFl3/q5QazQl+t23qCnzk3054YGVKzDD739eVNZ74MUlMd9xy5Z6ip8ZEEDkELQ
pbXdZR83mdbXmq0lIEAWVqzSxU63iMaxN97hJFjQlUTq6CC2wJpNgolcgg8ykJm/BPATcv3jLDF7
Xn7NeNAFUJqe3kd1CBMO4I0SwQPX911mntux/EWEudtj4QamOKFC96K6+qB8dFRhwLWjZCDqBNzS
3F/cKBTptaFhOj36hLMEn5EPozj4B60fA+EYR3YFWHYxkN0SXWhN3Ylo+Gjbsye7lasLA3Me67Ku
6O8tol6VEniBAzIvpQRTpdONCKk5tQG20nfZhEJ1DXuiaKAIqviFbP0lDG1LCdsCY2rquBav5qIy
N269Hv2mcoD/qlNC3cTLickv0KZvqryla6zX8jJHhzpOTkt30xHA1fRg2IVCzwEw8+Ow+5ENf2c+
VsQN+Sc5WK/7v2LztppkvaOuqr2RcjJF66BWZ4b66qRye6X6MTAQNKbGXLDtswj2NrBuOKZ3lp4f
f6S7QCOtkppS2GmBEQr/Xt88siax5tcP4SQeIBdjG+YyAy5ze48Jws2/yX4pWep4333G1uH+iJZl
vUYN7puVzn4tuEv93AyEg1gXz1IewWOe11iYuO7PUJUVIx3wn94Nc99BhX/YydQ9aIoYYiuXsjdk
NpWiCA9szvvUS5PCCtFBto7BXbn8EZvK9jQkITj5YiHcx9NotXfvCaWJmcbbDVgHTurcsjfivA/E
lpwxkCv3GQ5zqvdkGz8WxMs/AI4JHo2QVrYK1tOjcHrg0cWyfoe/y0YZdpgBqaNdOos8tl/h+qeP
QI02AH1j5L6D5TKoqwovpbiHlcu4leTphKlRJxcnn9CKXHPixLpw6+RRR7GG+T8rwh2bynoWDGqb
Y5/+mFCcd+qVTGvMsbDADvlD5lY93RrUX56w4tiYIToRM5aDpp/+1Wf/NJ2WJfUhCIVTSDJcsnFp
gEqCuRlv9GY0x1XvB6GWPQtHZAtrVDCqZEKgOYjI84exK9/HsfVixeLibIoCdnQ46yEJ+SzC0kzj
i/WrlnJngRwwLu417xH1OK3eE6SCKrfbXTfJhJF6KHZtEceWkuoDORkNv/mEf1ZmAyPjeEJxup4a
hURsOQpWK1xR6KaoLQgceIpsnHpzihMYCDL3iJtQBQY8P9FLG4vwHKidXriaPrkQzuYCIk/AMJ9A
HX2dVa6W5mTmETQR9YpyA76BaoO2Nl92ai/lszpV2uGD1tvnHWLZ8nNEkjbbQ4Na0vMyuI0OM9bW
RC1iqy5/d7Ux9Y70hoxThuHBncXP57pWsCum62OBcHZgceW7mbxdp+wkCtF/z/XEFB+o/H0bh95H
dMufJso9cLf4nIonQPnRBRwriLNXr+hRGQKDHrkCIj4odvi+y1WXNUBmMHSeEM2Bf3B5cFo6HQsb
Q+G/BmVdrOn4AIKPRiu2KPEThm0ywmDXGjEVpbx4/IxGB/8H8XnSw+cFnGap9R2DVeo9GekEDNlg
5dFfMO5gxopu9tGT397znnUVydWoFeXa/hNU/Z13hi5BqEwJ+GZyWk6xJshoA5XFyvltxrgG4IAZ
vdvpkP/hUIXJUwjAdj5G3e0Lxem3YaI/g16hUeB+8+86OGp1BpfQfugI+E76VGkVMn+a5Y11jPch
XArEgnW5XQvYkdf/frxHhWqys+5NAH++PCxTXXcPPTLwYS3DA8OTCDH6RNdbzliqkN0GO5ad2UY2
yMpDtqEpEmQP2FlY2AzFRB6h6wRhjrZlOIBsXTVZdfJbvrdS6aBoxQEz+VnaWgjktr73FjyaxeJ9
qYmlIdAoF9LOFfQbB30r/qubXInbKmw2di3at9lCUr46kqN2Mo2UFAkNXenHrOJA8LDzFclV32q4
ogbtzKIrexvmQXi9MZkHbxyVz1AetTA/AqlRUaMQ15NcmCjZqcwrvvR553NXe5m1ZY8B6EJBxyMd
AJ+OI/5asmmkyJzgppLxIw1nf7hiHpvcJOlxait5vehcjqh4X27tuq+hntHcrCY1BIeOEqoWN/Xf
nsE4fVQ/dL1Q4qmCgo4n+erExeRrO8mWPzpG9rvFDg5ijFQHvQ2KyxgESZ0hIsg+KpXmXCcppNwW
B6us9D8xyLT7k8wTUf0YiW7etoEQNFrES2EhNY+VCxj8Ef+XdxYObLIysX9dLey1aPp417QbrgMk
JMNUUwpvIt+/MuOmbrlEjFqtPcrxmGr1512zjB+IVGeRuo2rl9tctBvN6inK1aXUvcrCy8K3e92P
NCYOboS5pVpRFPDVze1DaL2SavSxQBfVA6fyJ8FyAag6FowIOsSG0psuP1JrIHLuxNziOFa4dtEH
4So7bvvVgOE9x7FSLHtlO7uk3OqtIIe6GLxdE0gdjDb/phoAgZMksqeOqmc2z9i3LzdQgrCWJ05Y
m3h7Jx9K0Ya8fphH4Ywg69anGKeZaEMNAJtuZc5ItLByQfZcoKqkvijSN/colNr5CQkiL0Oh7JWC
2iPQc+3rF5h23qnA2HLMIX35uJHZm9zrjL7O1+vYHwX5YOu6/cooHVEQiIK8Z/Me7cT//zfgLyqY
7e8483PfIhQt47K/nORp9JDzKtQb4tum4RDD2dCdzVn+vDEOD+xQMCdFgq4+LoYCJO79WcDB9FAN
1zy86av++r5cvPJHi835uYoyoCDxNdZn0D2Zow1pXvy2ljVv28WTFhyBVPKHhp2qSzLUcUrXOyb9
Q2L/ZsxdFa6by2i8BKIGCwjm6uQ2EGutCrAIjcr4CD0ACLBIpiyMVADMsiAfYosVK5MESG+qhL/u
YN9sKAUXfzGmxMrEC0Ba/QDI5VrHXlSvsNgpNJgdrQFIkU+uEFkxkOAh1Ki5VQcfEzaCXjcpklVx
W2BbS2FzLUwfXPgqahQhIYGukJPjwHEJsYTJqpvRDhozqCepaTiEflX5rdzdg1hLem7XtmQrvyXz
RogQTDZjni2OGzT5l6chmMHvoM9/em08PwDYZ2HM8p3uq2dZH1uGsR7g6OEQHUvLHGilVmMxeRL6
HYfWRzInpu1zAcSXLXRFcSsPqhNC2RIRE/1Q7fNEbPjaURXWQnOGl+ZKm2XR0K+72/2jyhH7Z5Dg
5UeXZRpIYO2wfacHEFhQH7h6/sHEt8YSCTzEeTErxRIdKsszncK1P/RZcjIUdzIzEBA95pQlNH5K
Rdm37UZx1q6OmGHLFa6U7usMX/WpUDimIuqxaIXNTm8qPYQMSaQUDvH9GvsDZR+HdJ2P0HZyGfHi
sSyg0EpKwidSJRWE9EFopnMegDfGfshXouWNl6ffej5fVCu7jmsU27l8Ji7h/V7SnECUs6/L/x7t
DMa+yo0EkEhMhWjV/Fys68CZmkv3E8JB1wmGFNYqFuW29ZJJarBYiZScXzmEzY2n8pjat9HN2sM6
OAhBU0vCrOK9fsTk3oG0KHmmk6mbSEKyPAq2ZL4aUnmXnSlpaGW9YhAGZfi9KgUfnWb9E203jzRk
YPrthR2znf6fhfibgHx/+JSN164jFppZj7gT0yES1Q98n3XbN/n4Eyqmx6xPWGHxFfni81xsQYPd
tq9C9qZ8hrScw7iV7beg24c8AdyB3CuU8AL7qZZaIpX6niveJsMaushtL2G2rMGs5QMmbYaDqCl8
Yxn4Gd2K7txYG/zenIXSBrAGIqrdaANTjkkUG94zlspxsH+U3jAYzuHCEpi6RttuX0TCcKyBPUnK
Of8ZKfVvphuN2649Gg+6jZ969ha1/ndweKB62ErmZusHZjc0qDALN+RIwSNDVRyuPi2BCIoOV5c/
K0HL3rOyqHamOYnQVenSQjFTMqWmO0INH4nomj+0ieLD98UDplZVtNKfp9MlNkPfnLoB4f1tnSa3
6ecQZGrgpp+ifncP27aRiqt/tCTtEjtU13/P95Mlb1shze3hdt2Fb1wNEA2jO8JqqFgq4jSTCJlL
08OPuB9zO9kOib1DdxQ1adswpl77wuHbKpuh0pePcJOzkfJWf1lvGVlmbKVsOMUYgyCRF60hIbpS
Ld94Sum3GbUAfJgLPApigXZ6BOKtAWXfXSlHSQO0CoQOxST90jHg2hzYtL5ciyvnUvK4lK9YjJ4S
KuxflxT2IGjXDn6XaOnbv9KMJ8VzT5jksJVcJbiKwxVIO0NCLcQ1AzVtb285/PZJK+TlmIz/FH5y
ahd5ZRETIMJjWXoKRVCekJDyjk5zED8Y/PuAEnnbEiSslJvC6xtVCHf+OyfBw1Y15/dtrsmJV3fr
9w5LwaKxfJOVqsw/aY982Zcy4X3IaWgOnu0kvYQGXdXFpw9797Y1Qs3sojqhaabDsE5bEXd7P/aa
Lkb4dB3oD2PTNKSrblJYMyyXm+bEPQb/qcafVnzhjQfZc7IVc+T3BZtGiSUPIjqRUHkWE7mea4z1
yFDy9VQDSk1A6+MDZ7ksfN65I8uAIhpztWlCBe9M6vd4TsXqFbcEeZfvOqoWQJdHiEtW3WFILNpC
wxasrbAt/JmQpson9kkjHVm6j/+qjnBA6Ui1mNPJG3c8Eu+o34SpFhEHlqJGkVCwlEH7r50m3m0J
8stzDYrFuYSTKGolv9HlVs14kZHigQ0JwVrUMfWsN832ewn5ou7kMPRdsYddSazn/tzqWHk6PSAl
bVYcLUT9RPCISnD0X9ZFOBHBwOdibNh+1tiEGLGYhg7jXnbSMZR1Z5uCE4W3iA9ayK+awJuZE9pr
WSE4Ev9VXKEV2HhpJHcsNlh2uMT8Y4I+j++E9lrniLDoYw45ZF5sibY4lsl24dyqMaWiL7e8OhuY
BXX4Q7sHSMtRwLGw0zuYoetkDGvQPlYybU0f7p2im5qh2FLt0Tih1Dnb96qO901zn5QOLDBlTzdc
Gp9QNtTSuUO0HlZyMeWWWYMZKjyxTRCZgoTVFt07dQgVAv8TWprP1IQaw+U84XltdyggA/tmRS92
u2rdRw0Zsd3M0tXBHeyEjlC0FZ0Wq8Agz75v9nRX84J+cqxocdML9MMDEQBpqIsB77arG/xF/07e
9/m+ILXPZHl+krqAakbjcGHEcuFcSKXIFb6lbNl5SdMbE4SwNUGjrW7dR1sUFE7whPurkaFyKhAq
F2ST8wNdV6PV9AqTlTJTdbqIPfswWkYv+cnF1mxzlDfew3537ThwrWvU+U4S8ZHf9ErnaRN0roho
W+1mxauSlKJrnEIthK3QWJOczv57vcM/MhoFIrKxJYI7P2YF3a6+IBa/8UifFYBhnDLBXMTwaCew
GXDDYtQxZu4KhXOWzwSyEeRJ8x1Nbu3pQolj+TL55kFXCeochd9PUitXkekQuLeX/zx+z/qkYW/G
1jidZRjLRlvjNpfizhhpKqcjKyHG+ZKX+e1FIK4ULlgmO1XZMLLUvKd5mWCjb8/pZYot+f01rFKr
X64pEprHAKUfquY1AQRWkkNyMStaiG1ZHAV9U3nP3pGpEtgzkx9VjwxYVGJeapqmUbRVCmKGTxO1
aCXn6QwoqwCgA/rrmrlHhOIN3A5k/pQO4bFKxM4D+/85BBKROq8AwzqI6fRGyv1ohcXlWr1iQGvm
fDGaWgauorFMX+Rfjt8YcHYUa8CFajmXZd8f5bLZH5ZYU3NU2IkUtlFkCqeviEWuvtX/7cNHpPHJ
oW8gzw4llvixzdvvGGU7kzjmdA/r/HDpvKtO9YtiLHIDPeuC8oJPELndiX8k7VJ4udSiE7Y0erCR
BD34iOBx9gFzYGsQOiz+J+Vm1UVBSkT2XmyVOHm0hv+JF4Q578sBgsa2Vne8gR0MO3I5+ua6m+AO
pcCgHX0y4kRRrxhpRTbIO8//dbbEW1CYAOCMpzKviBbo85g7Bw2p9cIVGpnxsWkuwXUEfnwULDOk
H2nvbByw8mtIK8Rto7CLTZfbRLCoN1jcQKd+LANfMCZp2WRwpSNtYohso8IqpgM5NQVcC3UxrHSy
SkARyGJnyP2d6siDxtfUPa9tJCnnIwISrmxXu4N0o8U0DwqmFsMz6cOJ1wTsO/HTx1JojaEVqqq1
/U/aAaJcDgkG6+RdV6/OjC01XkPTvUdmXxWetl5/Ptr5OOu8cFVfmRgTmPeV1Y74K61uKy9F8jIN
dwuRNtE2GGM7blzpFV00ARRzdVhTAuGMtsfPrFMXWU654pjUmIqnUiFtWbB/ZkRAEQj0qp5z3uPv
r6/2h/81z99WrqJ/yql9jZLAPK+dTqYdItIKk5v80UC1LC2vhEzpkwbrJfedoPmuopMTiNogkVFC
oxd9gHI3WV17mZc+4Vi+75qDsf9995wZHlFn5trA2A5nuZhzmByfjSOT8SlHrXzV/WEQ55rOoFCP
d+b9QDLnMC+1hipQ/3Fm4L9+SEhPzOhSsV6NsXKC0aJ44OcDwS9Qo81W0qRqJmUlNlJ69IFCr9J/
lfZh4LpAe1gLQp7i3V1lkrV1mtwq+ZwSQjU1S41O7ONMHYzUVENhVRQM78vLS6aLbSr2oAE0tDXb
HfA3cEXIFWLvREs8u88zbJcYXO7vIC2MCynddmLSjWfC4j3+Qu3HHZgMan26LK8laT6EwPFIYqlL
O+L7Yl31HbaNLNE8EK8dOVNcNx1bAlwOu0Xfq98Aib+/1cqQroep3BvNry/AcSpoM0EiLpxAdV8z
ueri+wv9TNsLfqUPVX9lXL0Mkln7/nmkhrV8PRejDz+anI/G7J5Ky85XT3upzTDY0/Ez8KpyVJm/
l36a4ni5MeJgOgJ5QYrSomhVLTXG+TJhiwZMPjgEBugIz/5st2pExbIMXsRdlXHS6guamka0P9HU
pKI/GK8BxkCyOepRlPjwHsEmiViSPJhctq47jIVCfZYfktAQwc0yNcTmSDNYy49TGn/WQEzybgwN
wyvUN9SrOZDODaS0jNslhqASQBkO3PFkKERtngqOOanbcW+MJmep3E8iBsG5cMouRpHXB63gIWq6
6YG7eXuIAVONz1uyTWaA+AXrmw9O9WCjmppYSeU5jP0seRTTWB7pzMjEdovw8g3yj0p3PpaQxOv+
l68GRe4BjR3kq+WJ1MYyMXkJQEjLrXRuPvugHMaXMBFpe6sZAK4rrKtAhSnS5FmuhsCQCm5u1CsJ
S2pqechdtENtdqL8REBPOoM+f5StU/TafhtMYwXiFUGzE9/F0BJIq8HVG4BHySlCmp3YuF+HYsOD
DNRNSjoghoySgOBmSA51ulA9h1Lm3mAS69+r32PKUOfgg4Guglbk3KRzDJuIV1vtFd4DL1KlDcE9
JqtvlUIQ8qCo8oRWmDnRXPOjSHshus1NYjRui5vu/Zti0ir35Sl0RUl+UMMRIhLLc0sw/Rr/MVZA
m6Bh8VpmMdX0w4e5d2tJ1NeyXXjhdkvfJkBmO72B671rPo0URLV0mVGYu5MGn1sO2Q+bAjCrG5U5
7qHortPetls7qKg/G9VSMPy7TabzxovfQAKCnNS5pLyh5F7A5SQeidmNOGSdAH6vS8IxR/2Aqzpz
XJaoDNlmtGt7xOyAFh9QPeQzioZ3gV/w9GoSvuixoXafRrhMeP8UblRfxV4ReHd5IHI9MnDNDEYP
yIDsXbFVJpqDCsg7RuW7SIsndKxqE1/RkduW27ESPKH1HGuh/2GGATwa5RXCWi8M9ZWcb1MvL6Yo
YzhOxRLq9G4RgEe8mn8UOMr1BqKICGJms6Iy8/2Wj4r1X45r/LifGQzxEmGHHs3oaRsSQu/q1DxZ
Yf5q8b482OZ04pkQ576cdiF601LNWVK5b0bvF2MFgIjD7IbcrBbfWBGleXXz2Mo1Ep5C6YdZk7tZ
U6uBQ73iFY4o94aUnMm/mte96v9eW+ufWtPqosoSEsl6xv4xtoEWVoHuzzXlhE3rhDoBFfVP44qa
5hk6vOI73o//78/MEyK+RIHJAfmdSWPkHngiO8cBrWDu6oQ8jp1K201voASKVcn8m3by9nD4UO+7
q1gdOQdCWrzBh2MxaGOCSdwu4+3FZDhDoiEoVuu6f+Bcf5e1bONetij2fTQMejnJT7eg7j6yjTuR
jw4Ooh5cP79bJQmbcEbpswpvHd8PdRa8o/y4jA/LoZnjJHXXXwJV7MajMOhDLnaW/c8UjITHT1hz
UZhu4hUFoOqVTEqtFsO8MhlQdjj+fJMuvV94ajyz+iWmIC3aI5LfNGfa9evvaYJ9q0o5FELjfHye
quwbaxQe1aXqKp+oBOLwuz9kk75cBYfkofdoyvjjODCDiHjDZWMTjgpUsE1/f0zuPqi9dgBrRncW
Bxg169kWGHneAoB+r8zYu+cDjW97oP3DWgwgaT4SL3L9FjuaibollGiguRaYhyHM6HEESLvq+OY7
lkoeUceNemivpopzmUYLXdZ3ZtA0E8oZ6U10TraokF4QXkbl26uJYEoXiha8cYUAzEzoQP6hNjQk
d+2S7eS/DmGBFNP3B4MZtr3vB1f4Kpcwmyi0ReLIxpxxiFsYXL6n4YSyuI4I7n6zii17OF/AFjr8
iJJ+Qq839cUl1fFt7XrWRUOOebhnMP/GD5CwGNQHIDODQq2hhtvnB6SYofMSOAI2RT5ybPOP/VPx
9goS+3QHYDDivnD3PZWajLIjfPBh2VqbsJk0uyDLN3LBcOMSOpIvaJAwu1P0+7amnL3Sc0kiuGFk
XPKdXr0kvD0fevX3ZpjEvU2u0+rUWhqVeMc913OdBw8cFk4y9UEnceG7OQxRbtOR+rz9rlJP8WC9
YvO6Be2Vg0qO70I+JmJQTm5XcjmMFlIcgSNhglvbOfYPglcykGhHy90P5uvSwKbuy/SYSOmO9ehc
5R6yhCgFvhqqCNyv2KTC9sne2qZ/DQtTDCwSIP1RaJtSPR8UMfoAFzvu00zEwSz++Fm/TD2203Ew
579JCL3oMd8urDJVVVSY6n7MicTP8YKGInp+qKhYhKYUQfOtzeMQO/WcM54PD5TMK8bmzP/ljQ6h
B3JMOZFU/z0jLB6sX7xMaM6iyHI/jba38Pp9ddEUc76LtAcHLQF7PudoG1kV75GP1ZugpevCCXyM
4ks0dlN9ufUZe1c5TacZ5C25aB9ISSIhNS3xpuwgUspO+yx5ZlroHzU3uE1hLRD3XmRCw+wOrjMQ
C6Gmv9WQODeuHCfjbIPLap4jgYSppjZ73UKXrizKiJrqOWYy9JMdnu3Y8l5qFAWMCEmxW3aQHBQ2
C2eUwhz6upf5jH63K0sXxHnWrp5R07i8erhFG+NW8IegWuNRFWaULezYBShSaQdLwLC1mMww9WbF
N+uKyVTM0/T5GFXDdD9rmO/ehaaeY1JFgO3EA7iKJoDxKESdlj7l/v+OZcRO4RneRIy5780s0Jdd
BplC1dKO5eD8xJnm+dQXRhhkuCCffHE/ReXMhIW7dJYs2n3Mf8gzTsyPfiT027teLI9bvDNtXz4N
J1Hhy9JFWNUTW/pBElHctLAKeGTCDgCe89WMR6Sc4AynQnSJ/NzdMRaBAE1zTXDVH2l7GG8unfX0
wNOVTHXWPkK3VCCwLqCNPPJoOYqGbZ2hw94Z9rBxIyeGhNkHiUYktCHBRkDsq7AWWLVsmZ1gc3XY
WCQkTe54LLzKM6j15FJUlchutG+kveoKng8gzCBURO4auLDhU2gUhXzAoRGuNMZLxwmJh/T0zyk1
T0jKLLD+lH6gVeZ0nCWVWIWWCw9zI6ByeKrvtI6zGyxQBqeW0UDPFPw9EegVDkVuAtNldzOOPO4x
UmPZj5Xp6m2WOglYkxCeTZqKOm4DvHHzUqkGNMyLn99hRuCXtGI3yU+IAdylecXTsTFi2fbHfmA3
bWs7RiR99J81v+eqVO7BZ/Dx3HyMpg+IOdj1fqORtqxsHHXzg0feJ3EOm1ooYMKOdylaHtBjNkTi
qjPCdmn4rUpbGcqt45BqzpMsO36+bJHbpOluK5klvbbbgQdNPpz86ug9xnJo1cSfRu96fNEcVPKx
/khVqS4cqW3UAPpPX6OUqnMUfa0Y1StLB9jEClSuqFHiQbO9vabqYetiXl+idI0/2gY70zO1Atcj
XAQBnsd2LGskexJArtNajSc4tVk5GY4AmKmSdPq+XbAoovyAwIQKlW1wft04/O3Q1rqR8NPm2Mkk
C8AFlidvVkkWNppxzNvKypCWWh0JiTcNctmHkoTFMg5s0PA//vKDE1CnmSxt8zeoxSUkBiz4oQwz
tgpNJXkmc+0I/3a3d73RJMLGVwLuiJAD8k7wmS5N4spYvX+xEjrklQfuGNgOASsIvwEsN03hiDzO
eVbkueD+4sTdppa+wqYGQsiat8bnzJ+/Jwg9U3n2WJgLBcgbHZDnKesF7bH71W6cBwspju7WdaQe
q/BmxpY0XhzMFF7KGMcirhBskq01WUViPCadPzK4pCgZ2GzPtUMgm2TwFbR+EnxBk6EuwpxmPKgS
HHovKlCgAitMR04Jb23OpTJYvAne8eGjZOciIJ7WDD+ifE3WMd5g7Jb0+3xJpSBPjcJvsqpsItBK
CuI8atwAzTAhEM2MFhWWicIA/6zjQsewDCjqftK3qGa8W4WVfe9KL/2CWkGgRm4JsY74kgC5aZIn
p/I2NNuh3SqXh59IGDn9hPZfTduDd62v3s4b0xNEOqf1sHnhT6Jvv5EDn1ZVF4TcwkzR9rFqmTZ8
2o2S0my6t32uDjcF696107C9JOv+VL7x4xjWG3b4CgIPBDdFDXw/NWcpU1gerWPV5ml+58HraA+X
0AifKkFuUjc/FfJY84QIMGnKHIdISXPw2thtZ+8QHjEbe9JxY4gDjDgGPN/aHYE8K1h7gWkD8tXa
nrdYUz33BN0Qlx8zJfUf3HkNR1Yiy6v4kNdcQIWruHC6xNXkcVHyxHr0HE1homagzGVDR8J0xgdb
z61snsHY4RDs53Me3jb7/P6VDUMqnZf3BstQyjcpmxDmqpUNgfXwLZWWQiIKuOAGhY9BCaQxrEtw
Qm4k8+8kwsglmT40SOUEGQ+IMYKCtK1k5cTSedFWDRhqYChMgDoRf/kRS92BBDeODMt5HdRcZgcV
RkHfC3nFRO4noG0YH9/mm8U9DJcy8yiXlVZ37gvkD6Xtwgr7HgmyfgWaSEes8FeOrITvxSj5zywB
/3A9VVrlbYyN/vgVnbOhpTiFQr1uXlY3fbeYqq8TB+UrL9xJbYtMocyPaxiR7zk1VxRLFb8Eef//
jYKspMQIb3zz1vG0m4LuoOOLx4EbGIpEeqWAdyH06U9xLVRafC5Ol7fqTn8GafUbSqzihCTKAOV1
7ITmwpWjCm5b47Yv5gJKiRBPv7ueqn6qxVUeLZ9J2BZ5yna+iKibMk9dMSLcShjX0JlVgtRmuw1Q
DsJcxrKQvJYEKzPyjm5cnqP8fZRStArqByCs376q10IpHsKNoB1JWNL6vFf1mDWGwgdNYh0EahYa
vv5lhjVzKTgdqIVZeGCQCj/0vvt2M1xfOKfgKusRAFec7pvCqYYloe+txA3ZKOSeHAizf6rOsoe3
yZ5xkoCAFBjcHcQ6LgX4ocFmHON3gVzV+G1MRgEiiBzGWOxgrhd5jCbWzCYslZX3WHnSJHfkC6LT
XIuoo7gEXaHg6qXM9IqyWmesPRPf6np9a4Xsxqv2wF2GuwP5ssZQPRc1qIOx9YCoCOW5s7/xHTiP
skk7o78O2L888bbQF6xEuk6MBG4xSfnMIsexHrDf8gTGTEXboNJZPoJzUF0kcTZkMvCFjsflxmIE
VXjiUKT/KhDQAqo7Kvzw7mnCo63db6Ky7NBo9htYZTsJ3M3iGYD1WNfpKfMVED6+lDjALBIK8z9M
n9dB6y/u+0mhsgCtkwejez5WtY1oMvz6rzCxY1Z0sLgg+vl4NHq1flCAQ2OWfFD6xi2l5nsZMo7P
OUJeKTNGb4Copu9y/cfwc0Xk2hFWRS8Dc3nQV1Ln2gw07l1ZdWgjEeFCabKbE8vieWtYoE0M/XuL
NwRPB3FjVZ/qpjoVI6GAToFa56zAQT7vwno9NkeupOXyoRTPfCGaLBTib1T6ir0L9rGBB+My2ENa
cFaS4C/Bp5dYSuWce81q/w6VtODXngHc0+YAavgJblZw1YwVShm1kyNAR/jdKzHqEm8ZWpoVi7px
HHGVKm32fBE/0AwGJVSjSRyrJp33yRZFxejUFJHchyhShynt2tQuplLff+3nlsndXjXzc8h0gk3g
VjfG6ttJ7WEGeYIH9zygJAlWUtbsPa/GTzdnvhAsTe3e5Y4DjRzFfH/IChzQScQASpF9AR/1cxIP
uJcwRY1g0wVgSkqoT5VrjgEGJmE4rcSDcWXmUW+Z0iLHiNscl0FUz6Sj+0PX2JKW9jnjS7PqDXEp
ufaoSg0aImULv+a6l4T3I8xu+ve5PnEkQ9fPDLCTJ1u/LAappdvwO9Ndaw0dsNw1b1J2GovJ6vpL
EB7Ce84ZqA4c1x+QxkRFQYyBr6b2Kro4N5wpS05MFGjoQ4aQM0M+4fjomuOqE1zjHEe8NQSkoVWO
1onbxJIcpZ9YYKmNNAZaYiA8abTw8fIeka0hDc18l1SYhELElGjk3HrUqOgiq0l11JJmBifTg2Zm
Fstv6fUwqwOVMrJpHdaBkbUwN28aXTqbheDBSJZvnvLZlnh5yr+p5f9cC9ChR0XVSdQn4qDB4ZGT
sxi+T7EXBEftcN5RkKsC/7sfW0NS5JeRWlRdrLNsmmjFTJUg/WTsGUL3jAzm1QCLGxOGvsjMt/UB
/zlAYnzTNvTr4Z9HE3myFjW/Vd5RPiZtSZFxSJg5mW+fN1BTsU4sqLIgtEz7uKJFzvdxzoMnhZHE
oMXjmrusNLqo6Wv3IGnbD/HmAzHPMT9e5G+dwB54fclUhdDtLcdAPYQjEdoikKHvZfhrd1dfCzFQ
eMLN7uIRlSgSTt2aykh+BsXGr1FVOPHW9MUxDRsXaj/wkuYiM9fsEy8WZKpkKZ+ElOfr/YGDjRiZ
lFkKj3h69g/NihyemApBRNI4hLuQEpX2nkVTCKxERLDwMqRla4IP7AuTZSA2GFOutbc/FpeS1W0Y
BeD9u6cNNTxroDVnmqtWzlrrxThx82g07TXQNu42Wb+um3g4+4QxnkcvhVxJqh+Ia2jOOQHX3XDh
c31zzfofh8QWqN/sAxtZOsUxLsGgDDSj0krJZhYvb+HZa2CT4HPewCmsB+y4URO4JbxP4bBLHgw/
AvcTSeD164RxQSeQDa7jqNWsLnqEesfK3ppMom4UcWqcSmWaOaZJIIIsvhbeTfvkl1VQ/jRyXiwr
QglytNnVxY4Le8HqCbtb9h51JyG9MmfxD8tghCii1J/yLqO59EeZj4hA8XUYzHnlUdKlSUOo4PNH
qVB6xPoiiJWSqLWEAotCE/EZR7iJWy3PpyQOYmsexHuGRdEcN9P5cTpntoTQTrlAOGZbT/7P3T7A
movVv+lHqphbJPcGIYBOEjpbpHK9U3iEJi2c5jb7UznXEkR+i9wO4t+i9Coirmys/PCh8v0w5VQm
+dSq0Uqh+alWuUP1FbPZT3WhWjy9PFWwaoz0H/dUuqOa2ESAr4obagxlLlgEQ2MQQx0gKRIyALYG
AH/SSqWVHslHHE7sz94wga12ABxb4Obe419MpHkFWA/3FYFr03yELbmq7pD4YIMqD11LgB3eG8GY
28L2iUVnznjtyPW/fW0PeGmHt7GOwML5DFYmeuof9DrPhfjkiTK5uIxmQmxApgk6MWhsS6cacxKw
7ZFtnKzRVYLXlvmsZEZQAV9tT1BpeOjfm9suj1b1X5xOoYMIr5aYEt8/fqMsXyFV1tBuW+StqwJQ
Kxko8idzPc36A4Di4X2RbEPIUb1Y8PLqQ0ZDHfyEzcVvTa42jiRp+0K/v0YxIjgTfIGzNxwzCFiC
IxcHCShTLLxvkPAn7EbLRCHL1J7K8f6WkG77piC+oXkFhVc21CIcNC+a5rTzTTy7GxUmKn2fMAxf
cOlHqM9YNGADEHb//vZrY2GF1xb6fPfNxL83THD2XVc5xJsqxdMJGtDXvFpRj+3lj3lU+cKHXeQF
tv4t8+OXoEjW/OK9IxwKFSxkao20otNfks359LgPifoKdwadH7pxQIZOGtaz+xfLzd8cJ7BVszwl
Vd3j4fPJCFrWmwjveR1mwEYx0IZzcwx6jtFwxf2SZTbrnnXobmY9tUUhOe+gn+QjcM4cRGW0W5gg
ThsA5sIwxhbqzRYetjSgxBvgbHD3creqCa4pD1qzgDab1WniadMQDL5uv2hpH86uwO2UgLy6rrJV
ryEb2zPFt3Fbu59poGb7CC0g0UxyrK3L9jjO9DM+2YkoEZKizmmGt9+dtdvo7Ce3G3RW2+6OE7nx
G1aOOw4Tyl2FCAoYoLMQl73Kc1qIH6Uga0nZJiP04533SC9nLxHAuiZJCmSyVFCX3z/dcmh8IHYM
NdQkOXxgeM3IwinGnHiUeIfr/kfAyQS0jebL1bIuD3ogAdt7OKw9vPQizy2aC1pUjOBnrHFGkcGR
852QN0eCJBG7TclnhHRY6niOeE5MFNlhPqVkSFd3ssABBHBzUjnXD3lpDZyS027KqAGcrhjeobRC
vpNGmIYI63WfQzmBVpgytdHk+GcoyKIt8aFazeRAUZAG+adWHgqNJUNPEDb92BhmS3x959UoF3v7
P3iik735bCjw6aT+4NH6e8fNGmXThB1vjD4Up+IASrjr3VvkBQnx0Tg2KW4nAnnqywJ0C4vLRT6N
1X7/IaGE4SI/DSyNpOsMI5u+3Xvbhb20o0xWiwcQOCmA8qww0IksSvxgAN1UdFNntJP1D8GA/zgU
WNHGLffSHKoZt8snkbd/g35/Twv2rDEa8rZdsJl0kZLEqaEbSTIFduKZ5ee/za9/QdNbwKP5WX7U
LDQMKU/ldv49WaHJ18yOdUosvbtprEsogNgxDwE6aZ2ol0FA3RLtlcPbz0yIyNiFUSXQ0TGmQ94I
GE444RHOV89/0RcFj2n/KlaZve7Nl7NutmdBWThnv+aU9FSckHa30XOSYPXUYnSvW0NDXDm1grH/
0SQyDabemPYNZvsUgF+V4/3E1cZcKnEaE+5omdlNYPD/z6ZzMRbNrHTyvlECGkaQxPhJhAuPCWCu
CIcrNLQrkFrzhyJ/T6N4vGLn1L/ZG8u+nxGHct9NWrCYm5D49s0PHFGyuJeP1GUDYT32epPtcjNy
+I+h7KdVBDt9t5lDOVryvvnRerKCeQQZL9uz8RAId3s4PiHlHdjTq7R7NwaUqV5NFyJSMbY8N5s8
WwUGKBRywa3mn/OG4bxPP5W6x0ZpvRqNFx3yq+HgyqGpZdfP/4oxsEnMnvVrqYq7uKfGA4j6dVI6
TJv3BW/INpO0uBmySfk74Iu7RIhcEhEreP/nvXsK5ALUHkBFeOHDp7sWXcs1defLQXmbkRwHlbMH
7d0xNgjICqqNyFS6U0/jjzQTA+OPwIDOfdioGbyPERzINV5eQQWpKQyTpafUApepYEoEcM9CSAw6
u2mJFb+tQmSyBb4O8OOif+2WwQXLdodKwBky8hqm8eyBDiEqMxvLIeDsqGzPdUM/6oWSOClJyecU
kewPhd0yld2Fsy7+0+vl9qjBfHdd1ZIVmXEhq5pW/bDmYQnQLN1bpVTNqPYLUQqjj8mwfEKCNcVQ
DtyqAIvmG1pVlZwxzxmpgpEsd7Etz44PAEUTkp2yZ/AjIFrdjpZg1OkrbcXP3MqR1AhH7ndxzqMo
cwtCVp0w+6e63hwoE7ggn+g/w4TDBUawkeDNqPaThc7CmWxS1Afn7t4hJqnJyjNFLZG3G8rWEuGN
9e9iQn+cf80dFfUUEYGoKjD6ferTu+UDV6I2EJ+XaUqt5RG2Y/knZeBBKsE3FO27y99cVyRldvNl
Dq6oZtyTdkZax0utjZIUXNICYPLSDlXq6DTf4SpeNTbIOpdLOIKLzDTgldXxHVHVC4t4Jz7nYdyi
SOQZwnCFkdwUdME7GcjoxoiyoxJBwLsjqlV4BI/BJZSUokyyVnIttBhySkg6EOFfoKoYKqfZw1x2
ze6bboM21ci7M+9bgG9H2NjyL8ZZdXChZR0Q3Cbospdpu34sQ4QUCjUSyuP6RsYrSb3ilGmpZpt+
XB5AiM9nhW4vzSGTttNCAff1aDgKfJg5ZV18Xck6jbhAC/NfVhcZ8SH9W/ljbZ5RbytTkcMlV0Un
TpLGnIGMr6MEVrcQ7cIWYnIFsbax3cC1jkPG6aBfVpOocfLossTAY2wimvUfaXtggN4zScCFbVi7
QFLg/SWX7qYm6CKKC6WwvHudYrKr0nMDgi2WNhwR+n7CF9j++Sh8ENgh08QJt7Tyf378NR5qNDoV
elthZYoFGxLCv0NRFIRy0pmFsqZHzXIxxYDta/DBucVZaTkGm4Yms7r8ckLaZWhp31gnIjyz1SnG
YWEf6qiAQ3veiltvOqtSQM5LlBD4uLuOnTcgXy6GMSH60cQdXWd4R36pYF6ySJQIambFCnJSA+XS
CDFAhnFlLWSAEkmPeeiAG30Og0LwAfFkcBfWJq+FXl0UcsRKmg9KSSLCVLYoNq8eKqu3IyPNMFUL
VPSDJY2ynMyBpIoEbkRRrJTb9/KgEKrCLMXOBZEIR1IHxOmbSX7Xa6gg72CJzwGHVoPq9Sve4zlt
IW0RHka+YHbISRVgURUKCGNQYCPWLRXybHIu1MeGx0s1TDX7k1qa44kY4ZzVQ7d4sI6kH/CIkmXg
cXk8FAHd7cyVALJxOm2L7+tIUXTiMeIMapLxOnYOQZ0z1X1qz9xX794EdwDJ6c0FeoG/oywdW/U/
SAi0P4TTyZZf+NlgGqg5Fv6VWTe78SCHCNeHLC2NKN+i1AHdMu5m/zvts9z9T05BuFDHlsm+sKCm
qXGHFMDjTCufDS8cv2s80ugjVPMPf60lXyJVayfNByXfF7N8WtLqvODpJsW70ZGG/Px0GvZKZx4Y
RBDvJ9rNgBvB+Vsqz1yGtAMmhP+XkpEb8Pz7IULgRkupd6uFDDfayAYEU1TCmT7rzsFCLMH1AYx4
YBMFN5XOtnJ3wbFMXCHKd7aI8zv7Ev7OK9LnuIDh4/GSB+71dja8RXEtNdfYJzoFBBw8Cl9FtRBc
tVUvM/hBNIRgzgTvewENrORPLx2RaDXOkQrP//LRwdwJaIaJuNzFIlyAXNm1FIC8kGodiXfhbIZY
WOWNV7eu7+raE5sVxGlo27jvFMD2MvFQp4W8Cv3SeyvAB7G+z2vg4gDjVA8LuQzlILhsI4JZon/6
9a+gPUxi+dgNOtP3Vr9uENCZpGIG/8mhMruEnKXDdjKDe3dQMcH7L7PIfIZOot8VyxlV13/lPpGM
Uh/af+t36hYxM1KAmnCMprsI4rFnqAezeeLGlLYhlVBRv5BVdmTgg5NST6luxOXKDhX4m28dTY2c
9ywXEMgu+7dKJH6vwZViYdB+uVValZdiCfHPbXKjQXGWYJzSCLYSOLdVrlsjHIb9AmMdBaHvh/Fw
I0k3O6wqFb00uWNeyqOea2T9vTxHNkDqqNWNJRWrgeMqqRyrAP0yIO+WbyK9P4rijmjVlkvu29j3
MRHNrbgDsq8XcPJLH/Hu3s3Srwu4aZwZoozV0r3/TR51DxN1ewD36RjIqO44zWs9Y0qhxrbfBKqv
weRKfLsjU0iKIkjfyrqodhhv0puIpj8AEQoGDukZiimCQ0vpdu8zPvar65ZiWDainrBPlqqC/wl5
IeSwZ5sVxTnYZnysBGx1/UZh/bOIyhAybyUb4ZWhPRTUDptllJPcdd7Y8w/RGmIE+AeW+YEucNk1
rG5cJJOgd9RoI0biHY68aeHS1nyP4ljpZlWS/mDhFeA76X64KKvGZ8nF1tJaWJndiUA4tgvIJaxx
P4bLh7mx9R9gyogJNTEzaegfJULd8uJPQFF1UZD7iImroaqkuglf1SG9/zmGYduz9jmxZleeHYyU
ZDS1FgP1QtCM9cLg9rM/QTEiJajdiJA8ZJymQiblKPiLdqkDoWAhEazEoKHNA6sVjGbSH8TnjPDn
Rgnn49K57QTFhsqZ3BFXo1B61HoN8j5AbIMj9C7v/xgYG8JwWxsQG8ImQtr2ijO5P+Hj7MXgXHlk
2Bq+t/lVDt+i5/aODp4aVUZu4zpEBvcI8Eh3dhT4DGjVQPLlnzfnKiTsAw7pEx+6GZt1kIcBzsjr
WBfxx0vR+iDrANWrYg3ivHY/n7MUAj2sE5QYJwYwTjQSwMhHqtQl1z0VRpd+A9mbwzx3grAH8q/8
73FAfSziS7VtkCzSEJVEYYUoNhwmErLH+/wO43ckuMMCADnWISLdjoMJJalfp/yxXCH0/h+sq3YJ
MkGaRuM6coiqCBjc9/4fTJsCIRmSqyipMLo0raiLRq6oMJoPnWUi54X3wG6vH8TJXAHRFG3M3UDk
DYpyz/PJr0SDIN/PRlfgSCSk9Cd9I2mT5Cre2q1SwDq0vtB7W7c0HvFdtrJbXoloYW+Qfte0WGv4
4ZECAMswgo2OeJds9GZ9Fjy5Gd1DdncpdZ5v8/9/LfA6BumgVrbD5Lae62hRo0T8qImDTkN3bD7C
FvtTqHk9H3G8srcGuBGI/GpepE9ZbNarwFhuTR+tk7tqaCp3ZO0x3fVI5Pk0I4yTGNpslBG/YM2y
3GJxavp9WMVofDjCb9eUPVEgN97GKs3O3tY4IbmJuj6kF9V9xqng3mkYAfK2TkD4/1mKSkLa3EPp
whFfehLoO+dzkJwFXLa8OYU+Gp9WR7I993lDESV4yt6hvMQWb0RKpTrL5tfF15BbJyM3yEmbW6FD
LbQ0Jx9fLn60arDdlUHEtp7zSpk5dyPPZxK7494gaC+gNOPdWQ+T9AU+BKWL46DrFVOVdSFD1R/T
1yeHizeQr/JBDvMVdHRqrBElkv+HE8rnusmeZXOcM6tgr8bRHP7HIIlaBZmpt5wj79X4wj5F43jU
1NmMyzptk+r/0IooMyxQS4p5cs98QcskW2wKC0muo3ejfi3p5OofD5L2FPoam0g2dwY0lCBtVjz4
/ThiPnDelynE3PQRyOUSHoz548nEA/72XTD0GkV2D6WUincd+t9nFBkFrIlzil3+vJDk1alD3num
tjq+lbsjmRpiVSHAYepg3jdBbyQuSmZi7u7dnX9Bc9QpLw6x40JxpTw9bLJWmBoJXeqlYgo5/0QO
JWUbQubIvw1uVpAjLoV399DaGH00csedyYY0I/VaeOLLZNcXtoAuFoTwyfC4fztD9nbpETY4gB4u
aYyG+2byPkdZoVXMWLqhvxOM6vE/f14RbE76aYSJgPHWL1j6kaDOp+2dOmERq5gJc5T08svFjTZc
X0SeCmojGP4SbAjnGvIrsWa1Gdc3oB4CWPuaS91WSjgl7coZiyD0U7u7jM+vjc7R2ofJd7uToqyS
Q1ibkFd3K9JF3QQJ0EN3spqNQUeVLVxIEsFvAYBZvwPIvp1zwQbbn+VBkGrtbhZKtxptipAia5bZ
rs2n6rPmxjbuRS9DBw9WqO9ayTVUa7Mf2EcJ3Miu8mEsEj36g67tqjOxfIT6Zn1nqr8D1qBZtDgU
mEc1H02QcqH5auDgcPaxUOmjVHlpMRBSagziiF+Lq7ywLxi7I2kPEYPS/0J+ktG7mhAXnxcPsknU
pW1f7zO7HvK4n5xqh/c49K5KWiqzFpnbh+5YUW/m0F1NawbIF2gXxxPWixJzzkX7LgMGcmdAIe2x
YyBgOuXAjc9M86NOfrZxOhIJIIcDSf+Z74GLVyjoEm4pF5uPmqy4LYQPyc0PDv6RoxEVXER/XyGa
A4caKWifXahPJhZHr1Y+ARc5azE9WbFWYugq5jx01puYEpV0iPsXarek+IZkQpKPL7j+WIpockp0
yZ5FSvpA+vUxLtYIAoHm21NyW4L3QR3H5w2/5SnWbQkZnEVrBHskKL5gAKvhf08eA04+jFXYzrOQ
72fjKCh745oTY+eyzaF5NTzQnkwv9k7Rkw/WjFgrc4BpiNA4tiFdITT2+WqOrW/fw6idsJsuIQvJ
2t6yGwObUv5qBZ+3tTRHSUCqHz4ZT1G6pfsRW0URpjdNH7KrdPIGPWDuSZaGzIfcwMYpFORyZApc
fgChW11c47LjCHl9ooJvcirzgRA0719TgnyUs18+Yx3aqs4ULGB8xQZPaHDitHZU2gjhKqFAH1cb
vk3cbLNartTbF0ft43w6nWsYAeR/x/j69siYpzyxQwZ/UZraDuzCpJZZi6pYFdT975NBwY5z900C
QzoODv4ebmCQZscG+oAPQx9WEQKtUoyu07xwTohuX/k+T0Gq7xuyHs7jPXxg++Mz+uzRGt5p2Aas
VG92CnBqgtOarUkNea5ywwA7LwgczRdWnSca0qsxKQVzfRFIgH7HDAERqeLFkMQIky/E5nsxJtO1
q8ybEelsATSFTKsRR1+lfDkUH3kPlxgll06nOgoCo2LomRv7ahnE9100lqBhB68Nm1Hm5sY1wNXX
WJN6/tsbkGClxx6EmVHslSSpQCDun4Q/md1q8XlgBJy2qmBMOM07s+ml6S5hm+/h1sS5tvuFbMTp
7W5d+2Q/NtyM4Sf7u1PvG2XqKy7h2xO+h1P6+utZbPheafVHR58fC/pI9DMXUxePLdM2riKqnGbr
yrqTNDjue+rfV+dHWjTTw0qyFBhffo6Y758Qih2zM0eFZ2o4UmEKgeXCPqRKuCFV49dGfdAkpTyf
N6+nvMjxOFsI8rgYWcNK/W/YjorwX7rmRKXJ1M5y6I4gq5o0dJusOdx6mvkkBF3/jTQWTjv7fq7f
Jc/qekI03/htmIbi0BEArqZk2C81LpW/1rHRcnBDRwf4B0ApSLYLUlw/92RRTjug5Vjjc32njZOW
+DwWXorVhCiBN56uauFqGDke1ezmY/jWIV6Q/ZuPVzALH3wsCDAFftMQNDjnhQ9AKbnJNxkKvFFh
PMQnICOGoC31NXi6ehRghmDAVkl3LeSuO376T0tvgWyuXySZoDIu1bwOWcCNydhucL8nE8E/H1Fk
aCQOaHaEkPhDP6OwB+f1nlB2kGWrImtuv1pEZYrIAh65ibnO/l6YwGNSjEJuVzVcbVQboK8eeOIQ
+/5LsD2k7HgHxrf4eJHZbLb08iz6Z8ec3QZTLWSDJy+It71A7y9ZxbW1TjQVkw42GnxYwnI0gMh/
EFFedq7uonDVAXqZqKhdn6wLfnC4oBm7bLmE/tZPdSTCaDD9/42n544qEAO1bRStq5y26FmtE988
TDAJ2v7myW0uMJHu6emva5x9wvoGLbfTtZPEJnqyxn/sE7PU7iPt2oOGClnUhV7WpHFwRv/Eq5L9
9vHN0fzBPaNMIoS9m7vSRsqme0c0F8LeboQVtXt+m/XZ1uknfNBUbWsTyMR5zA7PiU2IyeBaOW0E
h1dVXO8ESG1Ot/T1X1R1ieymaws0F1lN0BDWEvLNE0cmiXPB0jCyIhJWvbyqYOYyQGtxHfUdWMBQ
ogYePtGNORPBPSxI1iGtAF4Xn/m0A7jACcQX1SB1E0/XWp5Od0MR7OV1bMBvVSXQ/fy77zEZe2RE
cHQjHIysirv84XQrntXiQFrJAIH0ylY8Cnz+bRb8BewHXy4bBrFaYTAnKxN1/5PlL508qqQNjFr7
czZDsINWnFNcRC/N5MdfHwSmh6f3eTMU+iZRrO/yt3Q4jqx5dyQ4+aniBgDI4jlfUdpPx0JcvXfK
R+DYfrk4FbNrrD3j/RDdm8/VTkP0rj5H4FcBjTKteNO4LFfobizdH8mU0Lxhl9OoSTCLFJESQ7xh
tzMMNYd3BKf+ZZabbv70+ICGgcc4ob+LskOZ4+uKdf6xFqSZhuFB/dbjakVscUgdzKHRZPBTGKzn
Eu/v4+Oz6018BTSDgjyDfYwEozqh9gp1DKqhcLIEqVZ1EXTcgvyO+D8dJA7TPSIJJkBUdDrA/Ggn
i3PHjJba68i/lw8lGROpaSHAeWQHTjw4T68SQo4OfS6UWRgKHohlCVRnN2iohWXGIZ2fpffzyyeu
o76+AQv8cFe3awJarTOaNfI3+L1hjl1kVfqVneY+6e6vv5NihptXhn+I1FHoNqKf38OP1njM9/Wy
9n6KthKnzpIqKJiPC32q46tNdcnaCfge11rzhFKH2rYbhDewHXQj5lpfPFoetZsMV2rU1SMIS8o4
Y+ZgL7JKLOhWg7fh9aq43fqmHZ1boqqVOT3vVRcf47r+VC/N3ljjcLy9VwCAohqXGXuZwvHR/aYE
TtvL4WnS8YIoYWHmqSR5iR5Wg3Nym1AMvRdzUnrW2oQ4JR1vvFuWTCuK51EzFSOLBECAjm49euP1
BfwSKjxjIqjShTaJyN72geScL8JkzfyoiMSNQJRbO3McAVWxmaspk8cJ3dV0isZn+GKxpunYfj79
EW0BpaEQtLG+UXhSB3N7h0fJ4OdWminR4QxMxKxGh4XcH/SzOKN8dNG0A5nVIhbZ5E/jKMsVTy7G
vr1l6465QjR8qX6++UVXpd8KtfJUzwjR1URv731Ie/qBJmU+2k80NEnOUSyzGwQZJgckkF9uwzXd
9xYp/k9qI3OP2QavTzrL8aAofP/DKXF9MsKdhS8ahIOdH8w0+6s5MUN513+HR+ehedGRgLi+1k3J
PVhn+p3H3ODcoviiAjD3rG63c3mrmB8tOK7Xg2KjqcZPkQ+NgMERC2RMMzusWLja+xDQrZzi6U8g
syiYU36dvRwtY9ZUpGwplWGjvqg09rZSxQYDnBtZ8leiQb4EYCRQ/9LQEv1M060TsrnwYSHFK5RG
EF7sj630PJ8knhoy2spsrt0p7BbmwjDZHRwLlOLA9wy2JPzQcbnEC9e2Q6lNehaN3gBrVNF+OXv0
KFmZKk76s9NMO3FpUYkyYp+KNUlBjuBs1I3J7VH7U/kj7Nfz1Dhwin95atV8SolusVVJhfiWSx19
NHyv3yk7ddsQmZawDXNJ/mNG5OqLUxo+JLMz3kpwzO28NnuOK/LhmFh0srW7ICLuVG2/DHJgECLp
r5Wd8lA6uJu0K6FGQep/m1Nwvk/I6gB1utZ6A0Rx/2Ab3cD+v5ORlftiBZddfwLtL84Oe3wpM++S
IQWKQNKi6GzKGxyI99Dm0Cde5GhBsWvoBi8iYt6ptmu0WafuE08ct5BIw8WzB3MTGQe8q5J0Zptt
O3S7dxx/ZIhBvTzDkCZb9LdBiJe4o31rYcfXg1vLsW2SomL0U5xQlfEjefyFP7NMYwWgnDFAzQRs
+yb3Jg5KPHhWSqAmNYN2U2wuBHYpwcBwZdnMZQ2moAr51l4J83UySbtt65UgLeWQTvFT7WDOKfMV
49UPu4BtSq2ZVg0t8LUrmaQLcElCdHOhll1f+yOJNfkaxjN63AJu116kLC42o05mQSTdw5Vw8fde
ORcUyEr4ywNSqo1KjjCJobvcSclx3igVyYW8v80uDu1t1FtRi/lhTdFo83dWgxhSCfsib7crmLNZ
pQW0sNmkw7ZjEgaN3fBPHzFd2eBQ2IzbsqWGc3TGV7KOOoUH2QnmTovsJdQxYEsv3bhpHebDyw/7
15wWGRPeN9wgAwCf4bTZq/J23Dr4sgSqsGpDX/OWt46E91nxowSSZpyUI99glSN8uSFGhG5bL4gD
JPU+Hp6od/TZM+9CoXZxpfNQlS8pH5rH0pqOJqrJmSGUPms/CnW4qpvtw7COaopDasUCvigWa2Di
CNGsQ7ie4rK96VaAA9I5Dltw0Fmsv2uEVXZ6lPvVUxQpOV1BxJ4qrb1+RVLBPFSHbt7y/oVN0aK3
0tJ+PbLURFu5HfGCchglleHD3CVBXTxT95wy02sTLLFv81lxl0WO11irZ9TVXMe4tVBrXYGrCjj0
8FVYr/qFLZCupEI9glfb6WMW1k9cy4JtFm+twJ5leDOXJE8Ra9GgiPlpV9IIOLAnOGrtrqTK7e75
NiU98dorZh38N7daqKtNHdLFijSPYheg9HMiIqQe6+qG0s0MPF0Fw5XkuG9Wl8Xble3Bsv3KBdbv
VOa8jOHNq55fFekTDFfZJXL4tEL2Hvr7SsbpsIBihc27/48l39OcvyYHPlXiAWeb6CQaRUmqTTVG
vOY5VHhGzueCty0p39MIXurLPQlmdYRQd1jIMi+Innrjk7D/ecTPuX9G1aOiPTXvWWsjfRuFo6Co
TJCUITtedRdzlm2qS3GJjUc02fhIBgXjMR0IMvDXabcGiDXl9PJIYK1zmbJs4cFafnLJf9KwoEOx
KbQW6uu9SjBvkTiiLtvHHvWDbBvgi0vHZD5kt+otMnTs9YoC1nOjbtj3JgcCyNW6WHw95fmUj9Ns
F9HLjog97t1hSE9U05EDYwTzXmd8p1Z45p39q8byFneALMLhUkiwgvApz77o3N9ksSgupyS9JMRW
RGqmbE7FofsQYnAjgCk6miI/uj1/o5sgHpZZb8OTRk2902O7CM6EonggzhFrPLxUuXFHqK0Nl88g
69qXBCgsgXxeLbiS5VdUP/GepClLgnKef88FfOJnArwjdsQtISL8sfCiLVkIzrt/OS8w5bdiTUH6
aqfjZL9RCMnEJiWAyDBVjvr7kktMArgRIBf+KLbUGADKu8EaPSjoYoxxAmLWDOfcn4+JmGfFzHRC
QqQQ5xg7KhhqdgS7y7KWImjsVMIovbhZeYfh62QsGdeCQVK5A9eJH0Jkzu2RmaV4uBeJHMnAO/eX
cjqPoa9GGrxy3nFbIXwaH8AZWabak2G0amKLERBtlsOxGmnusha8P22k+QOwIDjPHI1rvjKwJVhq
QDFceISYMhl+wq3WxS5WZn+xEvIwNEea4gCc5futadBoOdqgrCovlxsDSV9IEcDirtpAeDF3b4nM
fN5sMCgQwRgLx8gtMJLt+f8TH6kdQcZumcONg9GMN58wWFQdHhYVxKauGASu/ZWfgPwspCb2VnyV
iSyRrriQ4M0EUp8oJfqqpxHZW/HXYwk+j7+404OkPkgt44lVLGUbIvCDy1P+KWtgPGspluP55YwA
9lF8LCic50ZWvq9k247xYWcfttJfSDKgxdGxP7S/CWSndxNBFnoPA45KBEvBThdjbyhUt+8p7jAp
ruknNO6/jKWlR96jYWmveu08z84h88WazX21XbJTt+/s1iGTz36ZsToE/CsEBJfh4JcJu/Ro/+GT
Azeor2hGNcfG8vjIsxAVN32lYvzd/ff7bdTGAPnEz4JWi4/4WDA+jbYq9OhXZ30TYn3S4gsT1tgV
rntpsmxPl4SkUqIxDZZn/UjDMS4Ffwwd6qP5UiiyG+5YSgsrao+ibvcyk/zaIUTDoFojMtiLuJhj
AcNqO01XBY2cfWfTvQC8FTNf9ciNDctEue5DvY94oPkgXxMgxz+qnvHv24q/QMpGlLl5v/+mg0bX
9fpYMBUAD4i9hN68Who5IZ8kuEvzwH39D0isG6QiFnNbL6QGjkSEUkgpiJLsK5qIuK/oVZ2wiI0W
qb3Dly4jyMLs2s44ZkHztpCqswfkQD2HBeHYh4EiKy6bpFHvyBGNNYQxXmFepW7FKwdPe9Q9z4hJ
Yj6lmxH+/k7IPxQMf9QIGYIDZvaAvAmEdMGGzoVOJP8+8xN4bQ0WqI90XiyK0TN/iJwSeO/zLeAV
Q/L80fGnvKU6jnf8HWViKmXZSG5bMMTJ4IQcn/GTA5cbVDYNf3U2lsvFkXWwVgKDm9w8Kup2JLLO
PfZVYewlrF6zJvvbP2V76UERpCARULoe/GqS57T7uv5vpgdTML9oq13MWw4V1rDtPspOKIGNqQ4I
Mux4KgirshRY865eoXEMZb0+L29eBNfhyDmJ2MzprIxxE+2+GdYNXHqc8EV0ziFhJVUEdaiU4DPs
0bH+s70VnDT1eqa7iiIDSakyr/XFazCGdTSgC1/THb/ZkYEuhfnXd0oeNl3R4OgYFgFL9G5tPYoL
fEus+fqA5ZHDw1gNuCz60ZkXtJcihCAF3eKluY1a//Tyg3Fzyk6/nztP/QlpTTIDFRxsewOEKTR5
kHigq8U6V6o3xBrQQmPTtZK8Ov8+3VWwjPO5Nxv88sCenIjrdNL+wsfhsgEfDNtfRLyQoZ1qOT0y
FaYSiFhgVMjDbKw3E+juVue5XLabPV2Bx2ji0dC+YT+qFmozjO3pjzQm3ouk++dKctn0uvQKcTW7
3O9zCnostN+AfohzsoSkCNCrTbdfOJRSqLD7obpfHwB0vCr9GURIAE/FuIt7ZXJWNF2dXowl0h3e
1an86pHCDImg1X/jDO7Xo6DFL7rmP0TsJVQ1xSL1Tm0mN9sGqhhbFTOew+Q0JDMM505HoPqn8ejG
rq1uNo3SM0kzokX8mfoxn9N7ddCcNVdITRhCv1R3+5z8qkHa8hHzqoNqSsgRmYs8wHYwn1WFjcGs
EOMhLW/3lxdJ6wFeLqdUDubIVH2Y2iCtM6ovtLIrPggZnYCfysL2/wPaSIaMcb4ravyZroSV+2B+
hu8lcpJR2XSzESpU1isGlNU5DYzPaTf2fMDqmh4BV1tEP3zuiFukY0ybBIwQan4s2V7c/KfYQxtb
52ZAn48i+M6uDsAMl5rkMYjGJc8Jf8OzCvvhH3jVGoE7GFXfItLEg5Y+szKJZbeypZ+BHzCTgQB9
FZVTrRPnPRnuxhphE3FeusoZ1OCBfexCyfkAZ0DeO8k8cFEGGs8lfpHZT5fqrsht5rUX28D28VYh
t1GG7ui6UwScGIhKAGlmA+UduooFc99bip4zUH8ZRr7b3dVADcc7azOC46t2yvJeMdfxJYaywkcE
2fA9uG6efvx9L4sSZ11tjkHC5q4bgLYsYTxPn19PO6XdnyPQAV/swUuNxtGt8Axn7xxw2plPifui
10BpOp6yFbp8U1wjPnisu6IQz3+xKJ2w7TuYfw5dWXLNwN+SH0f5srMY9+TfwdabhoWWX4NSS0Rd
+2/Qqt2ZwSexcddTg9jawS7gHTszzjs3wRpXo5ZCftMGW/T3vVeHGG7xajG0UD2Nxb2y9fsUlP/b
NBcmJWrdEQvMwJEBIfmoqsTdCwYyoJeVR2t+P2hVACfuOBtG1sopyRnFW92ELOhND+mBBuhLI/Mf
DeXfDUOOlfjYzxlwZgBx0fKpd9sk+JXRtqOUoRxDzR+K6AnunSP3YtYwpwt9ZCr7AkD4CLlClpvO
wZmnCkG/+9qFGXE9rRB+Yp1rvPzYfr3oxrvrCkReRFlnAHdS1iG8FJpqfAIucAeK4WU9ogY06pp3
k+E/Lms2LUoBMdWTfVMtjW+VvHlzHNHtagzGnP+HrIKPXT8Ba7IRw0hRwkrjFuDbmMo+SiZ0glZU
NUPOumrxwEjFFFVgl81hLRkcKeW+4FPYJCo8zl0X+ZUcBlPuppQfIeOXdq9CHi3+UgXJxS/oetQX
XmB2Rs97l7XiNvWjfkVX6BYsgsWKmaTF0m5gdPdgu7wvZ6ijVAtPkc8jnjTZYWSBKP70T0fB9oQq
2fCjTxgyX+k2BuOJyKL3xm07Pj6PLoqQKAvswNAW2lDTDDA3i1EPVotQLKClssSAw4RZN7sVIcpi
ORnkFv/j0/GZ7lu+ffa3tW7MpqwIbhDGjAPesLOxr6Uha94uAu6GQ+LXUJsVV7GTuNqhC1ubwSZo
/dM997y2yJrCn/Kcezxpa6adEaXlDRo5ZgBgoilW8CmLxb63sudIC2wu9IgOEHxGcz7hp93Kuxxy
qYaQLCaB8aN97WVIkPGzwj+RnbYzuThcMB436JFsruAFLl91iVeBdcLrrhLnjRzlw5SZYTuNlPF1
EacNdi/nlF2FPKNB7duSx8uDoewARbpKo5GtG0atf8k7kbald3C5cxnUFv9VDNEQEzJCEi1TZgA4
5udhtByRN5/dQaZwa+HziY/eU2sxp58+rW9gkmtHbrMer/hsyzu3gn0h6uGNZScXwzbsj7JYWTJi
ke8y9wlIvVpbyhEObCobAzqCvma+LtzNI9aRRq2TtOD4vFTRU07jNABMsZMnuwpzovK81ywnJNTr
XdakuugUM8ULE/pVY/tD27d6Tyhf8BjFKllxUC43bfJdSGT25vLZkbyWxDaDCi9RddBvB1L60vBW
sTm+5JiI4mUFxIxiurLbEqRC4NC4WA/J3Ali08x5h+18s/pC15E8s0ymPAufGqwHrPjzUhT1i7Ld
qzaZtPeCwyD/xRbgwkmPZn9zT7m+3GKitUY22+OkVah+wVDelQ9zjpLHxk2bjVumoWN2W355Q1Qb
80YVo5iq3WAuIPVlYSUnZZOezRqHA00KHsjf+tztUvgRhte+oDsZyWZSAn/xkMEOT7PBLIVwLoWa
ZtjXcd4CCZSMxnlgQSCHbGnDwA+NmX27/1N2Hwbyo1rtTds6HdEsPIc3gZS/FLWE+xyDTEI/qev1
6R+JAyCpaiUeRFklUOT8qmDmzIUvS79iN/SXZuFi6uKD10eO3HWP0fAcm2UXM6QQCqEq9EDAe+tF
blFdtov06lkRzaCgH89jeaShFVcuqMZHB/4CIUzgSGSjDqkoV5m66k0jUP2x4OZThdRVQ6L2bDgh
pwSdta22txMtYVZ4wMlkoICWJstYekhyOB4wnepXgLGZNdQpKxrm+gPl6RZXC5Bh2ZvYAoAuji+2
PlLPQ322BKZJvKmxyO2EB89gPMkjQQ3jM9zqkeRsUtq7QJaBIZjg0RQvG7GLyO+8YZQ/g35Ew3TX
1KZE5qYE6TvgpwdGMKVXfVHxqZwtPgKkbqAjDGZUX3E7qAdbiyrQzXcwTrpArZsXcl96tDVJPxBr
/0ZmCF/7GVbSsQwHRNT05BTQKjBvk5Ja1u1hiDsbXR4wnbDI0xL7Q3DOfzI48/jAx/lk10f7K7/M
M2lN342rDDerPa9e2o7Mw5ySdEwk3KrVQoIMwVURmIRebzJgQhMQSIs0mAL4i1GJv12uuhv3gRMv
FxEs5B7d49BW+FUcJ+Pz0debGen2njCL1WrQKQ9vtTpxJ1fTf68JTt9JG8cxCBRhCwVBDURjB5Rb
SsvEZSlAkyrYwAOHtGPN3QCs1uxgcBJngYpa9LGefJmeuNtgQ0B7NWQji5pM2kvBlhQLt38HHfNb
Brz8yo0A0zGf08unbwQl7p4tsbQiH6+NyXOYQnmwpv5818yRqZ4RmtMvKHTPVxykIYXcLpruOOwa
t+HF0ZQfgxLaeTPnVfgeKJsHPN53xzIfwW8EhJwgd47TycbpV7u8850vk3ng+2oI2rxmPanG1c0w
FFSa4q2BvvTE1PB8NYHwqZcgq3/YTkYiUoRIZAZvc06ZRpoDYoKvSNeCIYTJ+47c75k/pivq7pD9
JYqB6Jd2k7fFncLKVkYh12vlV1FqKF3/+mJ4BpWi8RAODVNBvZh2DNSprlzvUcaB9rASLFEnNZ7S
EDb3cu255wDjIrJfjocu9nmdZ9OAXHGqj5okzo1dHWd3abQJmRCmuf88vM+0MOVuQvR7xetvwCoL
MTqH9rdqcPUHkEEoxJfda4RUXQRgu0eB8dQGRecORQQFa/O9xJJG2PYJOpAPiuyva/euEKoRTzJB
96HIhmSJjqEPCBd5Rw7FYvSU3nf1Bjn24Sg4w6NtwLFyNE0qmN/UGxTuvxW3PaqiFqRRPFU1CVu/
w+wSHPcBi+KalA/86NRPTIjphuH/cwMXuMS2aGy7E7BGuw9CRriA+lJSewT+3HUuj7JiBBbrYN7i
2Z4zML1FyZBigqhfeYKHZFJuTtLgbTJwPbg9tirYJig8wgg/1FhG1hJH1G83If5jOIR1OJGUcT10
SH7fDBO/r7oGT2+tgBSmMZ7o21gj2lGAGFpUMqSsRVT95tmFv1/P4scIHRdC0mTCI/C8zThc7OR0
1eWOcXAezA3PkfBtXrmIbvtjuLKIo3ah1En3+k/nwY2F0D5D3j4IIK+jj8rMguB29WiamjCpYotV
joQmgGjo2i2taCltUkkkFQavx9sCakVTG/SuNE8Nv8EPRTYxhg3+xaRsgKpNc7Pw2GjVCWPGwm09
M8jh8CXqOoECvsSIvRg8QwK8nA6bekIdefH48suOXmNzNudYR4eGL3YoaiRN8rrTVKQ1maW8AADS
XcbXioSymy3U32K/aBpAqgOQYWf80xOTKdUPRKpuobKT9eTBnpuvxPK3Dx1NpK9WGEfo+h1emSU0
tduTCL3bVEJqhUD5Z1kEFEoJxBjEzcQ8I8wHCiVK0Hq6gQe65s3e+xrtueqOLT1UX599CjROKQQB
1BTNGmBYKQMOa+MdH+7ZG/rTEpqWlAqzwElELZ/HzO0iff6nDQjc7x6TqrncTHWAnLGZnZqWUJ1Q
cps0Zyk6KlqfXTQNUUH78ZBBqrUnYmANI3cA9pWpVXF/fav/KZF+8UiWX5Ucm0TIbSWogAPH/U1j
YX63kVUFMQXpcPhkduJ/NDOd28iTrfVaIII8kgSqxvrcUbAzCe9IUqrWkogV9lHaoqT5wFZqfjfK
2IDAFdzQrQpEG1nUcMSl9XV4cNnUk/OL3crtgfyw+KBgV+YbPlP0nA84EyoGEdnwOIt6irvjeigT
3mhwDVnQ2OBXx3oDuEFvVD9Z0/DKKydtYqt0Ml2l1+PU3IeJ2p+cBRspO7XLb8XnK6rixiJ2TAiH
Gyf2j2MFGfKYOlFu/3KlbGAc2jb8SxNOx8M/yqFtUTjGEBEbXfaBOPAeC/23B81WRewwGADDufqY
hdQQ40RClNtUV86V83WTLlvsOPLlRw475efawVN5OaBjkSXq5VF22On6HH9iKiZuPLhmcbcd1vSV
+opud03uEzYdtd3W1eAK96ZmHRuzBIDCLhoMQVD0xoD5+XLrZDEwCurTkS8a3znBscyKunraUfhN
pba+igkmEMw8RdqrvMFX8aWy8sRhVblIOIEgxtfv9oP3zZ8+GgdC/KI6L5UQaqw9X5rcBk4b8X6O
jDF+9DRcWyb2lmWaWDYx6dVAPKppoROpDDVezcZ0XUlfDaTCx7flEvzu8NTMZIlefRtrTumPK+e7
l3U2FRZbaBu4atKyPEMFnfWnb1T/yoqOrplDRdnu7F/4cdBt4zi6U9DN6kJBBUYQAAmVtXLzQM+M
9bEJHnPKPsYkzGTMkUBoLtoRrOdKrAbU/VUnqQMvG+A8ky8qnOAGCQXRhcutlXDvnB+C0Y7pObmE
muaLeoUQgPnDJgeGXJq6F1ETcp1YSlWLI3g+O+j4AJvX621zStP5P2TqKc2g7AyXfqlZBkPx5U9S
Ouv4iAiP5pQGjohLY70bV0sMOjA5GFA3/acIq+tFY2Kxr/G1J++x0L+/5KuZT4RFm+i37CkwBcEP
Ghn0UEe4uKAhiTyCztbha1f/UHnqbIUx7clVPe11XFDlHQ00jdB81YNc6aTQLVO1hCgwFH3bAs2W
CNSGR73zN+CQfXB5A9q2Sy23jeTrJIB5aUYWc+mcp36p/CKHqTpjrD/ctaX8cUxtOC/4t1RUD4tD
lRmnRK3mUKU35TbxPdPHaGGhDPB96BcIeHaOfySyvifWs4ouEr965GSgpA7Z1PRan9sooUnbW/ke
fSofHH4W8k1jP2iMsK8IpK0hPopdbpOs3Ls03xwEIlOblc42PCploT6crTeMAfJc5byadYKCqNtr
L9Ucy0/jQvJyQntUemb1GL7c4S/UqdW+NVHmC/GQR4DBwdjajlJwcZ8c2Y3+QgaQnPM36Sx/Mp8O
K1F66xcKyjyXWQIrsdb94u+ULARPpcPhlF/ISJxnGpnRL0TEh24dASGvSawHJe7DBpLZYJKlOfm8
IA++uLni7aEjs0CaedMbirwQbk0Qx8a2oOSAUeocKI6HpoangRJMxQR1U+Wls9Pl637/XnE3FLMe
H0oYWlzwhtvKT5AeaNcEN4HswhI2RgghEAXhJ6w8SSu8RhYrQdDNybuca9DXLhfXoS/9GsYDMU62
ZIkFL/9/iHPrwfr1oIAsls8ddDU7C81a/L+uFQ6MwyjyA/bl0WSCiYih/F3lRBpoDh/MIYtW5sIm
71Rl5WE5ZOayyhQV/5f1od5Nn+Xn7A8XqYIt+WgiFgYl0gYZ/NVVL0hMr7Ox+ps3Uv4ujxy5XouQ
MxyPObstNETvpBPXUxOOZm01U3ArwZTFLVjaQKRbVeMkki1PI9FRCWFSFWowkg8bniquKuz15GVD
Vk7dJgmPy5mbNP6jeH4Um2OdOVJ8Mws3D0gdcLHvY3k6z4M7flg+imjqSBayHSAdsL8FhfLIhtql
zphbZalDsLdUTIjzTlJ8g8KBsnlYebctOoFcD89CjGUdmyM0hV7sLlSEGBlicyARRb0QUShkXA14
k88aW8C3YptzG6v+DxItBaiSFvuZG3SP5Un9UF45vaCq+cb8cN+uznRWcqCkm4UWux0R+GKCiVHG
zcweU0g32vnEes5lM5iI1dMoANkQ7edGX7QGvbLXcu1231vzsyLBVVXkwyf7WQXfw+04iVjaDcVt
Cj/foIFjhVMx8oYYQf/l7J6TRmDtUA7GgICPOubPRaOa/mgAJjgTRKbWV9uQwpWytVs0hKYTihHD
R3AGMxLXa7uLOwcIPY4VsfkcKvk9CNCzPD/wlOp2voDeAxBCjZ9r4kciljCkJxo9rrgzn2NMea6c
aR0cYUBe3ju2oi4pS8PYCayIoiGf14y8OjXUuoWadqF3W8zFDgppv3iqD7cXBhv6nTzfRyRGGCqp
LBQAEzwK9XQ6jnxaILdkDKppI4sQ7GpCxzvZmP5KIJf1F4ROYpQng9wf7ONZP9A//mqNunRLdk/1
Hw2iDL3Vs/J+uWaSCgS8xYoZILqBDNv8aI2YmMNDR4nEtVtQ2qlK3CA9Xr6zMrsUKr0HChhszsep
TJoa1SkpscVpFYuDNVecNwxs3+Xv3Q79t6TGjXtM0Empijf3Rz7s3ZVjkIaiEIEFZs9Y++sEjm7r
ZU6kMMQAmHYi+e2miOHR3lj784R9yIQ7+5NhHT0F/Htrqm1LlsdzUjfP70ESQR8xB6LgXlIHsl2W
2g2FjOj8D04JakmWGJaX6hMqddi2//FOCFnda2S5APOzDfu6haW7yt7rwBbX1Yx1JeUU79RpbAxg
JHLlwtjvsy0nqHs1kuHHML3GtNaWhrw/QBG9clV7kAQg5zn3+1vryIm1SBUq3hLl99bqnt1tTrv8
mlPmCEQRvsserPD7qxWmew6iUH7AKyBz7fefdPS3CCzcy6Ewfd9tLIAE2OZsOEM3UDZ/A9nkg81h
HIot+Lvk920EcewEPhkXEsabzoX7JusK6sJTC9Ka5BGeexRYgbg5V0vAoS8ck+X2u6JSmgbmRJJc
Vs9QjkMl+91IGhoO77aIsRWmz/Gb2qW/pvohzuvsVlTQU6UJkLiXe/TN5mgKIuHXGLLIPItv3vc8
vVl5zpIaPFmJmt2DBFLnaRf86UC8rr2h3zXxH2WxjGeeg5IUAJvqSP3PkKPBYRpixCKbQtgpudoV
sYU59E5ejPTYotkRRm/G0mKbSRz8kNXPBWVDqD7SG4Aon0zbyjKuO6p9uNQjnB20atmuGg9dfbnu
SDKqrNUSps2fA5MchqF5Snz1zxBydGQz38oggP7GRYXBHj4LI3kjQlWSkJ8i8aT6yRofRNZ3SzN3
y1Sk0/sVWi3fozbGRGU3Qyv+c/aySstaPmZnv4qYZhoUnOhjwHfh2UIS9OBZ/nO5z9JBoQ6egCvZ
HFGvady9rgQAhlRytuq7YoW1X7PLFaSLrx+IsNYl0ipRXU5DCRg1tD6rAVhIewZbhsEdon2RhXhg
SryTsK4J2BigsVbdClbIiq85dKINchaZeiIU3RJvpUET9n67t61Gz14YS9eS0DFQUy/H65asPsDu
te9z2xrUZ/ywxvyIC+q8VIXEYe5BHlQRVWtLK8O7aPfqGSXH/KHpEHCq7F1AZsBWZ96m3mvElByC
7uC83++erQL+ojSSOreVt+pc/Vh2mZ50WOI64AYcqGYHD3KgjUaaVnRddn07cH5nfP4h2YjWYUpM
mFTfypC5MTb8YpGRhNw81H8+7GYUd/YTJR5ngka+zjObc0v4Qd6JfKMZn82nFuEdMpWWU5S29M0K
AuHsnj2ExrXqxR8OWRgMPJ3YZKDE0G4DqW/z7j8SySL8g1vFC7gg8ivvVTTk6f7so61nIClnvSlH
L4X5twsHqX0M9b1P6Vhz94FicOqMQV2qn3VSn+UARIIppLtaaWyo61KzUb6TtKBVWse7Dpm0Z1lV
IRq/7lE33QhgDeXMHzjQuWVpDMkap3ZCa+WaF+X/pFdIeL7qjwO/ZCQ5biWXoeHSvMd6AUdhtZ23
Lr8ePQG3tFfTP02w3H0PNU1Rn+D9+as/IB82Qqc1jfY0oDGf6Oe2mMWp/ZeNzTesRlNEoJEbcPBd
HQwIGXMGTNhl6djM+EiNgjPZe7kPGEafr3GX7sPvmVbgQrM5tT2wiRiSzGI8H9bAZgvSYwSqP5iV
tUChmmKrs1fGlowAbkjL6/8WKbjJ38i+/hP47595pW07DMVpnZ6IsVzkzltzO/yD/CcvV4hGwcO2
/LoTSUzIR8HYGvJoIZuDd4GRJgnVWPNP29q9zG+Y9gWWKmp7k+CgLkedHgGzm/NJ5mm0PeKgy/SJ
c1hJgmHB3ES+4yMBDguS5K3YA/SSFK4kZWLegucfhFdi9+bHEOkQklT0I36ewdQ7vQ1tf++EwNIB
voPHDcJ5jReiosN1QPASYmOiHRTM4w0V9lM0Emkat1cVv+2EzCErI9W5ptvzug8AYszn9NAHgJmx
iEbZzI/gpjM2WcO7a3KpTPrpveSjJ/y3ME6o5W3lfgLIrk95vFQenGeqMedP5Q78O/Dn4aNdYyLY
xicPC8g7EehJ8/VPtA9KLEu17tKPETpO+83u7zzFOft+KHT8GeJIRodlFf35O4W/7B3A20wyudZ9
Zbn910a3IzJqQpq70RxTk7x6CnwSyaqebvw0v523DIg1aNvubCn0zwW17Qyfvg52R815gRbngH5s
a8OgAFQxKADnfrcGOpfi9Ghf2qWPMJpKB9Y+Oo4snBBj5XRxJgrk0KuGLwlN2uspGRyrgFRG9AQs
MbtjFnbghJX/su1IgpsJuGZxTdLvEVp6q5S+BbEer7Bp9lcy2D+5VPZqcbxfDasRGz9nITHIRIrz
Bw7391yHCkZvpIW17KOYhOe9+xH0BTOh6dBaXChiP7Y0Z3tDIhcCDJYZn8KEIGAwcNsGOpI7w9ZD
TPLGf/mvY831Fe2c/jWWMu2yZPsTJDMKXC6TeZNxqDb5KPATy8ax/6TQRMMYlXFiFYUF3YxcSHpW
hreKRF0PjdrPHdFRe5hLrygam1fKXW1xnpDzodZvNtxoVEZG+KoaVcwVyVcugXA/BdElJlZZtVvm
wkyYgOlvMmLxXustHSCt4EBe9ZdJDufkrkh5XifhNzl348QshroIlk6kTJpZE4M45iwbq5r6oz74
lgPYHDLl6F9dS4umoURTxVOgZ7fcgANphtq2EvJygDERi7QNXII4lab8PeF/ZqOzNOiC/RiRleIv
zKpqm2HzD9hBHqbUvWZYYuZuYEne+TsNTH5+ATiTgTyY7Y/kzgm2WP3LKV7O0Llq1ZEqWwMEeKsi
TyYB7t9TpcrgPrj2Q11KLZEqZ5P8RzbwUqJAYYARLs1Nrzbg5DroGjs+NvTQqXLzcOTGt056jRuJ
qsvxKOSEjN+I9TTpp5W4bnjgLcmj3POOA42Y5N9rY7dwVq21ER/hgI/XHyWQt66y1SpZX13i8Ep0
FEf53KsR9eqeWPxOiglgdZJmhOFkNa0ANZoYKnDehI0op+fjgkZTZS0/MKaGAPXhXBOxyTN7nacU
jaoDZcEdmM92wf3wPF932tQfE5TCMv3TG72DZz/gq+xk7n8B9qY0MIsfLUn5hX95aq+MJc8Gk/Th
LiHf7BrGd2kDLGiRdVhakqvoAfs630DCO6zZoIQpkgrpsDaRWX1HKMPzNbK5VfCE8rE0h5oOQtI4
zK+5Rc3stkDDcTw5/Tj8b1n/75u0sCw0GkSsEOrONqU4R4LT9FehjIhY8BJgVH83+5G190qlepek
9y34FJw97Iz/FrV2Z8e08PGv4fBvQTgQVMXJj/y7KVU8i5LTNnbiSgWwYLr5c5qpSgxpIyorlP+N
7wMdUb+INze71ixCfH/rR+HQngNK1Kb3DGrCO05BhK6vbNyvMmV6AuRKVtRSSK6eE8aTKk2dR3aV
Zz0x+hHzuWPXwb1ey1+rcUpsTm7VGBol+XI/3vTGRd9wW+G1hR3PpPug9GtvH/r4R6F9sXsV1DH2
AwY2SqGUqjB2qkXm+ib6wIf5dO3A2stjpap8fhkYLX9FozeQNUsP27Xxq8BypW+MYtH4cvhevle9
f7WgEAt0aIVdFeIKgKR4Nr8mT84+kZLGGelJkg7uzrxG6ixlSQb+rTV1P/FlmWhbg1zxf0ralgRR
xmOhhSQfhL2WgeWC37DabLwHoT5MSOButUf0J4B1F56oGDjHnauTLFcwZq4Wv0ggprQ7wc64Edo8
uMv9my5/4U2lDltUwHa+am0OdykLp9U7pBWHqctTTfWQdreVFIiAkaTxm4/6UyyZBz3JrnjaWdl7
wg2+D7xtBrRLqVu1/qmQ0VvDUpSpPE0AJUGPoIwUCxa36SziS/1uqsR+kmCOpIf8nfXd8KGYamtt
mf1hYz/IIAWLS5Zt+kqvFj7CS+bkKA6Kp1LuDJM9EW+QfIj5H5x3WC+XXVhQgbR8BWr5uJhqa/gJ
nokJbV0FFBXl03rsXHZlagQ52H4i5zf3RZBCGCBT3pLV0tH/8rWmd3IVmJ2Q24Eggsf9l0N/WNRn
OKNfbwCaCAIZfW4DumqYKPkWnreieT6SUogFopbISaEt8uGKUm/lBOyS3xyrpx7m+qysDlwOBJ3O
taJURUKoICPdGlg7llPwnztxA/jhGo9IY4pN/xVyBWYaEaFL+xmP53qo6CrHDPOiTY+B4lPybEZ1
Bw1dX8/61Jfb8NuwavhTcAjxmTRV+DKkn9akJvur4iv/X63bugCk19Ro0V7UUlZnzyTKi2JzACQJ
u+4jtEh3ITKUDMZikCYV0F+txARkD+vMDXVf7LBUYJ1/vMvRdNaG6AJabPgUicPBQGPEfp1lAu5x
emJfWpc/9O2U+mq0llSGdb6Pkt9AdoS3BMSiOqC+kEfVPci3aldNlFdTE0k9PskEoDc0F1A5pNr1
mKF4B+PNDRT1H+W+tCcKMgVOd3UY/PDbnUIa2wm1Qb+bOwcHPWEJIIrKkOIBG2OXbrGLovH5I2SF
f1Ps7lJOCFTP056ycrWDkijoD2WwmS9R3gG8dqE8NJwxeO6nI/3d0n8IAZ7QlB7EarDmac4+1F6A
hkjVgdXLSJ3CCyJiG0DniszmVC1KjEkiIjHlPacxPOrvs22/sAgbkYXPmZ3MJAMNeTYDYxUiKeOB
VyyKys92261NxPzezwQUlMGHc779xtCfsJY8g5E71eWsnou0823zajP4j6x2RIjE7jSg3b+6OyWj
+A6UzfFSYdpvsku6CSbWQuPVxcqNEQcCMvVWQhRlYwxQbmkEsQPGZBrKqlPJPkCROly2crYPX0Q8
Z4vZx6TqK7oVwQMbyI8QTacugyApB9B49cLXfJHmKfC41ndmqqA9LicjBM+uw8Sv/wgbFUWARjnL
BjvsXonku3wdwDPgewORU7X74Y4L4XS1rF8zADftGh5cz32iI3S7YScbCSdqw7abZcTTWoD9o3sR
3kAbjq0rDp2hmqGGYs5/dO00a43BDKjMS8OxPjkoH2t8dz8OvCBJwgaKDNWoAfIJ65aRQj1iBsi8
C5wHdGV+hW7CuzEkSEgAy23D9h1wRgG6MS7PnQz1Hbc9OqKfhzWFiG74Hqp1GEifiv4BiJASpT5X
QfrnCa1HK+fKv+7PiDj1c1/h84lq41zqb3Sr1g+S5nNUCvFXXbRaY1CyYFMVncGv06+fgHesBs4q
iYKHE3SjtywuoTmO4Hid7hGbK3sbFf6zE24+eM08uKfw6ngjdkxKNK7UlFICSE5r5F7y8+8vVprP
hCrMygqbai9Lu9f4gCaAjMBg3Pme/dXLpFm/KBzmE21Wu2SKTJDcBxpU965P+nxgcxEWpBFp+Nyq
tx13p3ORPE6esYZt/3z9cJij274T7f5+lYJjqiElhNs7s16ivCQe1mw0BDgN8R2lCcu8l2kX+kVg
V4jV81xdB+EuWXC35Vwu2WLRgl7dhxYPi3FPIA6wKkNRJ4sm3m/2FmXQpXT8XmM4tcBgKKy3F9UM
Rim1Ny5SFYc9pgvEJjx1UKh2XJ0jGcQqMYrgapRHXEEDU8PJmwF/HevIPb74FujRorC5L4IiF3KE
yc0/XFXzMT03QBzP5lbmhV/Z6pI+iQrrnWSBPvIi4Z2wM05M7yqHacFDKzD3P509rHQLK5W0GFDq
v5O4OsV5Hhlhb1X8GHpiSzTrp4MARZ1YykVS2VlrWzfhQbJgllo6PCKUE6Lr4ON3P0j/WVJBYqPN
zAV+O6nH/TCVe8Mz7V0lNa50ZB8IfYr6POhDKE0p4nKE2oyL7Dsw1GuAZV7N1IEY1svqLQyt0rD4
VuierhIddYnM8eZ/sC/0LUt7u5Y5c4zGIH3Mg6BEOUP/J6fVUKFdwxbuFrGSuXg/4exUvHJOjtsX
Yl9q1FiSuAfbnlbY+ntRzDykWml06LXz9fxfb198UQfSYzehFjhk/sjuw6vZ84hfQ3ZsJgxLH/xm
NppxSGZCnH+nYxpsgf2MmDiYJJmuC2KNcEAQTBUkHtRwDh2KrUH7gnllA//ppkGx+3vmh0cTWwWN
qsqyQUoo4HabNwuw4LfrIy8TexyaCBLr1q4mHTJ7hVOL/B0p1ahx5PC6mMTu8960z5ZMjnQ57UXH
iHHG7bbWsvRy/yoI6LaME0i/os5S2awhhEtv4eHrgzVGSeU/bhWo8PwSa8wSKpZT2kwRlQp6JFoX
U9EUTlLOt+w4xBlBvytO4Xm3APT62LE3rbJXPIJ0VhtMolhl81t98GTl/qz3t45DMsFqG7k3KspR
o4xmKo3zET2J6ObMOQ8Ue4J55iFiAAsLspiqYf1zpqJqq1xKFX/DCXpHd3VlsrCBLSaux+tu+4TQ
pg8LnPI3XaapqY6znBWFUG9IZ2ZqFkjVx3PwNiHUj0R0u9bcoH0cBQelLndiDSZX1tlqZ3uhzWiz
qyWEJGrDkUJ/FWP86OGVtO4q1nDOHXT8nx4hr7LXSaP4sMT/8YVyWFIcUMu6TQZYX2m4i28hltMi
lDGgx8LO4FmqHJ0eZMDh2YytFsV8YjiCvxpAzqiExXcgDiB2edygTTog2Cg2bga2c0BwMauYBegf
7eBEsFZ/IP3eXCWWlog+AV6d+/TalNDgeKvkZGbjUIi+OcF8c7C4eP1GNaXZwhvfPXMFMN9qusCv
rs7joT2Ik6P1idOoYDuVDqTTbMZ9lyxFte4sRingdLg3z3Fa1DMaT1CFwVl+4YA9ABFfpJAGfbMz
5PaaaZq+61P20OcxzAJEku3qd8F9c38dikNdauG+aPKFwROdsf01OZqJ2AaRX9qHr4KnsRUlKpSc
RKkPsEAODHGRNNARAveTWaL9u60SwIXq5M+Wg2jLk2How8S1D4OypCrrRDCtp2cAJiuU+kBb0BS4
wNntzaSiO7aTsuqfBJbJnHFd+6QVCc1ZbD2X/V/pAGyRerIU9EiFNDvQ3kfcLA1DDqQORR4V9vyk
QVfyqUbggqgmqb5/6+M+5egNlquVJ1b0ktm0E5fH+I2xeFzosEZRHapcdRbtn5x5/cX067LAgh4k
cC59j4z77ta9Pqa1QCk2USbx+N7uSmJzQJzjIB93KpGIfxO38D0C96LWGO127d1Bf3kTLa25i1hc
LCAuE7Fp0AqdAE8+Zv0WASfYEI0DhYKuAptgJLWygqoPERNO7e8EJOucYidbTLBtV0eAozvNM+Y2
nzQijPEpFIx58cxv5UpeVxNP0IcaPfalMXNRODCtb8S/VWXqQkxCWBh3ZT3ptj3nC+w9yDdKdaQo
99qk/s3eMsGxoHDAyawUK6kbAG9P/nRbDhQyfvgMeCpGs4wgqwRbIHzl60UxHioruQp31XMmN3N5
rShJACNj9BITwPEU2/LDI7cLnfkdQeGEFDYUvFu18I9bDaOiKOPRvagkO86iOf5hWtSJIB0aVqTk
b5jEEos0d7seJEv7gMMhqL/6TaYKBQjwqHP7YXyXpqQbllpmxfs2UBP+8Ux4JjsuEG12DalPDO0s
V+FXwtyD/Fk+i06+0WNSlcy0KfYNgmHwP6xEZTMZsrtN6kPHKmdbm40qDyO+DEI5CG7tmYqX9edw
fyIPGTrLJ+uoaAnofEiLrQLS79QgJmBiTaJQMAPFZffWHEu2+eMM9xuyZMCfaRKyG8/hxxk9qRMt
6YL93Q63Sag3ixkn4o2IEClkuVyMeMybGIR4UmxIYJv+VkNli4Ec1Q/woXRqwOdA8EGRxfMH5kwC
ZIFdFStfXoi5voYjP/anoA8j7DleVBCKcTak3fVRUdOneKQhkqtgQGkbtMKOBHdlifyQsDvm/ohO
D/5rrRU66g7MbNt+grsaqhN2N8GmRS1uYabjsAbVJgH8gB8Ebd9aKnsvYx44IISerVAJgOu2L972
WTqIajPVPdQZiF/aQrX4FTsbQ8C69pGdIlYjebM87hsaVPZByt6mujZEBwHI/TinNy/tsm9WZMxE
X+2IhEigycyGW4V4P++SYmVbYU7EEugdtAxY9mNGFIHbY78z7pThWmsw+DMmY5CC5e0ONR+Wjq8k
W+8eUxUDF+WnCBmech29A2SHsHXQFJh3hV0xFWIYohkApjMzJPa9qmVXhAdKutTAcTwrv8oRfq4i
/HVQjOqfYnva+cXrjWW/IGrWAnBPuMKTTk2zD3wSXMOVsKSda/FL8VQ3FjM3a1wX5a81+dN2Tgtg
LvIO59pNBIrDVYl8xqXCe33wW9G3ffXt4MYqa6VGlodN1HlS1r1753B8n9B5VHeRwSa9LhxdmK8U
jWnbZiz3+GdBy4Jxya7QswUxcOaq3rfBIlF8HE1lp9gw5iHMAqh+x4rySh6F0P8b3r8H5vLXKAAO
TdR1kKRCaNDtmfBNEIdMC+rqwU7tp5GbxN3AZ7er++wJqPw2M6eApOzS4V/1/n9fvRFMYEEMNPcN
Goix2U8WDKAdFjde7ulY6sHeo41KJd22iodww0sAMoSshArZXt+bYuNRk4l7c0/MDK+bwFFbueOz
7FZUDR5V2Q7js5TGiupjdbZB8jxIRWqmqJhb0y9ngwR8cfnWk28lgPrNZWtmWo+/5tAfxRCf/TJW
wnGtDWxxK3RsDR4XHiB6wSmHssL5AP4ivlwO38iyi7RMcgE5q9csLiQonf+jR7Ro6WIam4QKVRm6
avGWNkNe7aiK4TePkVxPRyAdGLwTbZCRIyPnw6buRPqVOAVaTbrUiAtRIEDqpnBW8V850zocx/zX
9jNMbjmWvOf4TcOaFOz6F5F5QnMhwbPqDn0vHkE4cW/4VGzzj38FsajQIiJDe2A+FK/tMmfWwKEq
IyK+ZQk14nQDWKNqqh2d1dx7Z5ZRb9gKsr/QnsLU34L7d35cVkPkJodCA6OHpN4UNevc8d7Om5lW
ky0LDob9dESJmIodypQuvuWV9UnTfTlVxSIK+nUcLaxn/ufegbcjZBdlBbG5dvnGAgdNMOszJOug
toL1EzdXE6Ddh5ZOpMyNaX4L8cYITUxZPPgOVqijr5jrwuq2N2ICerjs4FHczyxNQHue1Oiq1bWu
idUDzonL/jSmxKJu1U8E7Q6OrP8H1l/Dz2xcgpuManzkvDjlAET2+xkObfhZ9seJwxSgavm01nr4
AIIXKQ3CtZIlpkN+sAarFYaU4irtO8NA2A+Cm+gdUAdumqwI0SjYI45TgOPmuSR3UWHym4fLqYQU
E7hJMO+UYA6hJW59Vz3kNMTJIGWDt9FHrKsG3eTT8QZQLDNJy3O9sCl4QdcYy3LRTZ8rd1stMVp/
6BYTUe0qdXiKpE+m2f7/WI2fhQ4xcSqKAv5y32U/JbgIr+tvRFFz4jAdZ6ByZqT/8TvdwL7unb3K
41UYXIuSBikYw5m2oUzj/o9adausUbGpJDuTglSD4t5FZJpZugkfd1qyuSXcTVTkSq7LKC/x6Y3q
1q4tQi350VrkaSthZwPD5vQc6IoAOeEzwZh+fUNDcwPOabkK8OwTkaP1+rDUPrYSOP8WmvIIb7oV
oqlSoyYdZaA32N+mZVBwgZH+DZgzvilqKtpB7kwVhRPYzTWVOC6FWucinSsDA11jnqggzLL60jEM
6RJ+ktPnju9iuCr+rNKnRe6CCaEcXv5ZM8ysqKPeizFVNzag18GjV3AZHNE/2mLC4gZdty7Qs4l6
j0sTrZxZXSxTR/lhEodYBqHlhjo1GDrzCtj8k7Pu0eJOg3Fyp3tEL7UnXr93ODYVFvcAeCLUDPnu
BIEUAlVL/mo9ZsN+fiusYoym54oExFmBJYBxp8CskzSnqp6TMoxAkYrvny3T/Y0IMs0xZhkWyj62
a04cSltI8ce7lS6INfEGbxA5SUqEOaWo2ouRaiDpMn5vC3eq0WED8so0Ws6cmPB6t/2H1kkhcqdg
EbXZjIcpCHO0UA4D1DACMldckMzgkGYYeTI1qeZmiJgjl8FnUOL2I7C0BP5e5LwOTJaLuTaEqWtZ
764WQ1SRfrZXm2dN0PuOP0ySPCwRwi1oA/IWcNbGwuMmKNaBtKVtSWE8HejKDCciNcLv3fTLbN4W
xsavSwVTTf9LKoYZY3GTyQ6DuXCIcAXEAWo+p+Sq/1i4A7WYbPpKJuWoixMWsIe1eEYySgif7344
EXSBz3Lzx0WqNMD0rpY7c0Ha3AWgGLCcewzjhANGPK1tcfwsttmFwcNC07KYGNlXu7JxPm6PP7lZ
d7ycApBA37RBngfC/uLTq8Kg/Va4Y2r4qb9FCIb9ZL6Fa8Lwy/WiYuVrijGgNcny66iPqagxeX2K
iI+ZO813TVYzEbIu77RzVr0o0wIfpHNKoEUOeRPqqyyWWMoGgdX013umGPUib8b8vmYhmPjzn6Ok
s9qSdOexyWS/CLqLKtSGCIm1cqQRp12LZPW0wwZQOtscmb1rE5Jw9aoinh67+4c3gVO8xS8C6l4W
1DlKaTliBJz8b5MjSQyN8P8LF3deAqV9uqSa2d1XKNk6yUr/lU1X3MB8ljkM5Z/eEt8ff7axYCai
/NodcYi+P835MXUPo4KXf7yTYR6vBK4eGIPDr61cvAYxG1qT/34YwFKLJ2r3niIgNh7ZtIrNPfje
Q5h28I5Wx5SXArz4TdrOwP7y4ib/soNRzOGrDqJmQcLpnUC1IhEOqjnBFYejmeJunfpzcqWCyGv4
9B2KHytVIKFLszyP88+sqHPf+m2h8g8rcYc4yzku2+rwpFc/hJ/InyZdX8539va1VyyBlLgZClcI
0meBzQmh7Fw7cAvA+g//sqotzoXmqcKlV89h0TbqIvGKRKJuIYQ4HWzuspDAeLCCM8GPEHk8iX9K
4SSOjxKVc/e0GKFB2wBa7Y65NPqo6SaiML+OALVDborBER/0gKwhh27kLvDK+vXjqu+IYJv3KTp3
/1Y5e4o+nZanBCXZZKe+eYwuBFAueLBMPgFrwTUqvspov/VVbeeI+5c0cdczdcdJMwedcCxqlP/S
O1RMifgEuhWfCWfaTP3bNiv3xijp7rTREl8VXwF6lJtkhHg20gYkvkoc+G9jrCpdwNy2lI+DIP32
oG5Mt5lldNzN4EinYFZEJmnxSOB+fGKL4F5bmpdsL6T3pB3hooOtIgwUcdbfSlC6OQYsAMJs/EVd
3GvhyY6wclzfCvgml99CBeU60aVDiVofMWQ9QXDdC2Xq9w/6bZKMM9gFl/qdQtzHAwupYNho35+J
/eN55YGVUmGaMQssAovhFd9QuoEc/tX7KuJ2Q21+CU+v16UsKvLNufXmB9x1nhXE1jyyp0Il2xsF
CkmpxWIcDdpATEAC/VopUxmMHbKHKdLxJ6+rJtU8jUaYeWA1dWEjKbSDNPUeTVlQIUW0OMorVwbj
lxPmpRlBgyQmXwM5VI+zqOEwnTo5Z9PynmmvTk6JuVQ42gt3ls4J6cnXTpdHhjf97EQLvKqQw7xj
RfYW79e22afS4W1z6X3rtvfp63pYolLrF0SD+VUoVxWw26j0B4/TlHezGqWDjFNJDVEW2E1NkpEb
WHLA0s3aHglNJTVdfE10+Iq1G3wm5fucwuaiNVtT+pu23IlUDnrMSv6jdO8lqCJxD9Eqp/u077WJ
mwm4YFfBEKt2RxOWYGuhC2qRDcnfba8tZHZHve08kKAQz0TGh7N69t3nLfSvCan0RXScg8dtw4pw
0fU/1mSlZlu9ihJ6BbayQgtkKl54Mwk2tFvdWb7TxDIVJFB6waw5jxGlXNTfvGCujsKIYxR9zdrx
z+G4EcDcOT3ZKc7549yFFAzTIIs3Nw9CsvI4hDb2sCKlBKs2DQ+ygbp1EBrTLtYFsZVoMGyuNOmL
x6oXhYDLKWOj+AfekcoSp06JQXZI7AeGCJ87NbgMk32qwoEzZHULFp1sKE43nNcV+Enuy4dzjFQY
rQdy680UPXanD5biMIYKc6yJVj0O/1oB5y5Kj0Sh/qVrjgDVD6Ntp677wAirnVsTNs/C54MSMf7f
lhlsOYFRjn/zslBFFeg1KTQnWS0rHzDrhBqXCX/Ko0lr++u1gresVEAUrHyLoAFf08eBJ/TtgH5l
+FvRQAx0lJ2LCsgvQGETfusTeOyb4JXPgxgdnQipsPuFfTDck1fgCaobqqdsv7JYJagmWvWn+M3F
M0ou+BctltXRMMdpDQEv+uLSMNkUn9Lh4dDvEzwnC+zND79v2BMoBrqRkS9P2WQTYuhUGy6fOINa
08a2HmUxtNkApI0nZqieM4D6qBh/rR+wiSffa10SYHh2FYuKAqA+l4olv5JKsftVvVzyp5MPQWsp
Jh5YWp7vJleC0q4EQCY40JRA4lskfn7pfjjHJhuSfqSMcaz8wXwKllU21Mux2jqOiGHiEA9QK5ro
zhBAOCXM7pu/NstmrJFMGLzKz9T+Ks6SLyq9ex/h1MfBubrA/KSEBQ/kX6cqIsU33WctmWO1WF9p
1c6dhsH2dD1GxvckuH+6izF55k5/IOMTaAMZmidJcFrItjska1qL3X012RHotY5OiUPVI9okwyWX
g4nDdhdF1NTW893MC8octLfJVXtlRtR3+aHOtoa1txwwNlJdrwazAJozPamrGoeaDLOo35CdPCqY
OMybuJHBWWxpXOeKLSsjSZuQO/TFSo/n/tUkaS85QlCWRH5kYgqKoyDdDKbAop+TD4CbIoY/fYpq
owYPQ/GbH5FVFEZjaSU3G6AQEz1LlXWSucQjiQCiZSpb4z2sY3kMoJMe/maHBEtj+bHElLleRocK
wpgSS3D3iTeYuaZ4H+4q8ctCToIooz0qs31uOLLWDJGF/cQ2m7QgfD83OFIojiQiqZ/taYwdxaQ3
VxuHzQwfpBVUJ8OQgxwBUTd8SC17o1R7ipfMWRl8AXWfoVXitc9BLySb5dJv4MfrGNQ4mahrMtTz
n5VPpKDfP4I410vLus2mlU6m1fYwfp66zilDdXRlcDXmWubayuSU5Rba/qkH2HPyXVx7fxUslj5o
Rzvw9L365DS92z0D8NwSEg68w7ME5l8Zakb/tUm1K9hUlKmpUbF5qkhxY2DYdx5cJ93e91+WPKBv
JBn7fV3HEbs5KytyIc/8k/sRz7Ekpqh/uXEVKp01YZtdP2LWjoFdiLn3uTjN1zpUD1rfZ0lR78Ly
wtyQUxLW0iAj+MtHhOCeIQ07XWpBZN1isAtJODUGO+RESFIAdniUTBlpYgrhl/s5/ELSCPCSlEbj
uGE2xR1crrAqjU/Pn6IyA0bqYzSPxvzytQbTZzH1Kjc62QcJuz9PlXJrI1ERT1cfOoxHU2O6+Dpj
svTOQFp3Kn9ZqG1F9imMqqHJTQP5a1Jx5yu6a3FoW3hsDYzvQ0Ni4penwwRlVGAI0LsB8s0v1fQs
dru3W6M3YIN1biAs5fT3GkwLzuRmcYT4v5e60lKYgzwtRYnIzU/ta131XkEJd8GnWtkMurvPhImk
5xc29IexKD+0YXytpvZbcKFG95mWtrMmKfNHkamFeUjmqSna3A4/jLLX+yqabPLTtNDqaNiPMqQ5
vpGHkDUqR3Nzic69lnhWqmyGZFb9dvYOEmr7EkHrDlwNri3+UN6IL1swGmN6i7dMFFxfq4CVZPIP
DEPGjI4qgvwahIp43B2JGd0JsK7m0iaZcydsYoy1Kj1eYAYvIg6fzUCeV8+UXeO/Fl/RHQnKXJS9
cp29cqaxOK7LceVtvqwx4FDc2cWr2R4gTRuMsIljRjRmCzcsFESOSYpfyAlbSKXtj0HxdASAH9L4
DMRFsjQMaDBVfXQX0DOUbo5BAJ7mxC6sCPiYEdrftrrKK/PlggboygG4ut81kzVPPVQr/mS6zK3g
j3PL+V9HlRz7km+ob8SfQEo0uERSoy+kM1lJ2h5PQXGYDHahreAFZMxCjk2LlMF1onuXTjB4SC0Q
3LY6WAPwwNRsKxLvnqvm0gN72vZKlOW+VhNnIpzhrVC6v8XYsQB61d9NHiBlrtEyY1uCjOplVs2k
JCZX649hGbY2tKAyh6LY5Oj2nMzF0UkfNnIAyKE6Hek2WuSrdTTemJT45TZA2yTEOvaVKkAUpW8c
bVI/HfBJqM3gePWmy6iVzchiyYWVvcAi2NZodmy4ohhqnIVlge4pWucPRAnDrUhKXaHQgKUe915D
SwTSbdk6pSUJAzqxMnCf6dDU92v6l4zG5maHc7pY4zkCW+P2l4zk75TVV39Z82fEE3an+RBGv3vX
SuxAt4G85qy8mIvkpsnOwA+sw4vRkePw1d3Epv05bjG+SkTjK4kDpxDHXOFk7zSSJ+IDYzeLZGIQ
afUJ0ECqNC0IQOlzzSR6p1AdnkmpV9l7YIQjes4RclXvuNjLNR9Xo180jnIoaqEPfHd8p9CXuIUk
ZlhTQIjkJsh7lmbMTn19TzqlEMkmPrK+uRcN8UJCqLDf1jZ5f+8C0hQ7uYoohpUtoO7CGEqURClL
TpDW795ck22TEZwacm5GAtSv7xDtS6NwnS7QnZ/DK1K3UUwxLq/1kWBPhQ4shvcJVYSFnW5p7Ih5
YiT9Ev3y4pa8wrpf62eiiQxRyn+f/5co1dPXJ7yzZ7aj9eEvBrUDntu7fYa7vnQG0x5rgZ8gI1ol
g5IwpipAGaqvqU9pnTcDZTpkaVYmVpmEcOfNkZIaaM+kXrBkjl/3pQkRRGJ+4M2hr+azrTmQRzNN
2hOw3w+Ulat4+iY7dOoigoMrfaTiqg0nctfhgOUR/Y7UgCVuFtKuvoMIx57wAk6v2Rc+pVUs4f6q
486bOfBSQhAOY1e3MveYivta9JvAunNFY05zA1y/2LFRWWiy40ebQOUvrHRCgg6PNwQaFOkJDxyn
TiQU48FROTaKgYaBLK0BIR3yLxEwMwabkeK5EadzhL7nmjQYYu03vGEa7GMmoWt2MNUaiEE9uzzT
g5SQBNoi7EBeabSMm888G6a2gVQP2HwVjHLw/XG0jL9p1fYtIxD6ML2zqG9Uz2kE2SQCkGJpgNq5
wY5D6+A8BLONKl8maBrGpDwFJALcwiXZ4/L+phR8r7qBYU+XNjmH7THWKVsEPqYlMNhSHHrf1wcd
UtG7qhOsRMO7djRmvIlp+l9UDc1eY8JtCmHbwayYFcCEmmsT6F+gUH0uA41Nxqokl9Q94u9WTUYm
qIykMHnQgp0oZd+YTJ1tZZ9nKWxuTT2grCGmNq9O+8T8xBf3lGicp8H1FelGuX/7i/6Ly9N0GtET
0EeTAaul3rZneo9EFJFv0TiTjHosCa9K3bRVqWeq1AFxdyWnVUTeobgAB4oLx5inRU02h0ISjqSj
WkxCuCH6+tvrX7FzJUSeB9vWrKH2XfcnPJ+PaX4/FSKUeSzJj+mDHtthTtgYy8CTFMK0bMy2xksP
ddLtf9NPX74k73BipO+MFykEowbtdGy1Idj9RJ9Gti6PiByvaeAvG8TspYfmI8H8Y8xqiv8DvjXX
nxmevR9mnOFSFAKi2fbjHgFexlWbFxnWHLgsPw8As8NHuKWrYl0FlIONg6hJAMRSGpyHDTWI3cE+
Yq75yNuCstqhJiXREKifrfanep3AbiJyTezzl0mfi8nvQCsoCmu9LHWujVYOmYRgxZWdVcUjKW93
HnbHqsYXi5amD4WKjGI8O/lZd2ImjYj7ZnXk6IBgxq7wdSCER6doa5hIPboLi/2bxGZ7Yr1hedbi
YIfRn0FRZR+gTUE3nHyyaXFpbeE9EvF9RWjtTmgJalaj7pE8/sXYc6RvxaxKJj+kVbjdztklOSxR
kj23dnty9UF7rnxMen9OIrEbFSgVpkJxU4rAjjB1XRzeLpORmZX0rwvaV//F6OAr/0D9dGuKV0Zq
s/2um9xOY3eWRqP8qPEp370evU7Mr+4RoX5+8nIWySgs8tiGCyiDWa2UQuomCLOLjW49+aSBTx3j
Byo4x05x7n87VBPzDn3sNd13ow0OQBwjUNkSAHJ0UPhoLg58mgUU37xyXvtegvdXUirpmpMNayxo
xzlhP/qoSAWTC9FuF1KvgFfVfibvOEnGHBeLUVzWAekdgs3F7Cg/46abrEqfw1uYjAazG1yd7f1d
4l70gV3Hk6iNA4yvATLZuB31e+HxHxMEHeLMAAZcZ7PA+oAfZQeBzybbK6hXokZJQCr3k81IrL+Q
71drsAQX8/dB1bB8GRmrekWetO+11UQo8PvllTLvQV2cpHzY4crK/oPRHeMffTItt0J82VVXIv9r
1srFokAYO0J61ryYKH/DmS8ZkKPrHySRX+GdBfqd7SO0orFkRuLS+cSz8nYrbj50wyEu5V0bCZQR
Q3F77FM+UOejq3emvUBHjPnCUjBVw3srRFV+aHTsiVB7xSs9Wu1p90V3Jn0GQqRW9eEta9FwWMlW
yDjbfxXdvykB4Ud6jOQtB6JZJP31mI+8BiNIOX/Z209A2MRnRlIp+rJ/4LjI1kPITBAzy/frjlfa
b8SgvJdd/p1oWXbqPj05BwHxmctxMJQ3aksvSdzY3xZFTgHWe/CWne+9j0mS8da7e9HuXdqpr4RV
4q+w4fpmL2Wm7VUUwjg48Z0JG53hTjYyett9OcjKjCCAYOVDwCQNhQb1HdEC0Vibd+KCN851yATX
tf3weyaz/mNy00H9L/5+NLErjHFtvBc5E/YzB7UMntycauLzHvK8iYGXBeP5rWYLl7A1KnDgPsCt
aOwSgT2WzHRMOB9LMnuvK66UfwHrOilxepCubyt9OBIxxZSB5nUGcfdEtqxCk0JblH1Ej2nqykt6
LcRo0WW4tRQL/TwihlumjtsCxny8Wc/gCepKfs/8q0hs13jKtA3wHB3PvMGTQNpclIs/flZEw9ty
uH3mjI80pHYyE78i9cMybwMUVDWUH8sWx0I5N/f45DAqrVb9389rELy7srslfD4Xd1bKzGojl1B2
zHQfBkoEZMS2S4Gw3G8Nh7LBJj/LCglkVWZRN4Hp8uummPYBT3mOx3DktDXk+CRYdxbdTyhBolg/
0canTSQsbNtITqZmxHdjp4rkrx3ithczhvspF+CJTnw5RbnFgeya9SRRlO0FVUKGvsu68cD/0TCW
Oledceq8oMsjAyNd95PuVBJP5tRes3gqyuNGVOCGTZ/vrhym2iBOSND28/qvmUt8kF52wz0ffrfz
EdLDPkbCjzsYhkZt6AWqTCK2jbDjS2tK+Mot0zeUNxHG+JNgor21W7alFQryT5MSeMHeEvu+3u7+
JLAQqaEZda4iMBmd4+0U0n8RABvdetw7qF88oZRxhUX6yvXEkZBOlvVgLAWWSAF/V78FnBU6lAwM
FaOZEZZPxRGBIHrCunz7Yi1598ZmdoEveX31S9Moo53cTZFA8pi5ydYPyx4PjZ2Z8XwobC6LQKox
5vsZiCSfYFqoTnoZ3xRPS017Qy3j1TeYuMrVYtJTMQERyP22Qof61OxJ+DkNt7dhYSzACRW4VWJ+
6zS+daCxJjJJ16pu2z2PKkAjF48rL46QTtolsOyL/uLB8HhDSjdUKvyO+GycOsSBAcjVJh7HDqI6
r+RS2UpydNX9gLLS/90Ad/mPQpJJ4F22YkdsWIQCl4rsLLg708Q3oN7KFaSmqP47aWC6qrRK4vm+
/YVsr/2JNTzCAhPdE75U/vGpII8bCHewxNCmg96No/4bhIMOEMbJl0YMtpLQ1+VK3rcs72VmBR4d
7CDNdtJIebeo9inlaz/qPWlBglbzVCyHanYQYK+aVYS78BtXTj/j2NUeOkxc9mqsLt806+DXH0Ox
1p0mc7o6m1/Ll5dJb7epoLtSwM/rKuKnHSM4h+qAW2UaJusr+InYGk58+g9OAYQGOwkooy4zAn6B
Q6evlbI75UiTJ89J12rwajrM7EQrCx+NU7WwZLWI6jHg5bJhOlGMLfcGoO2eljoC5+sfROg/ULAb
jYqvnCeP7+m+MqajK6/tksBgecAz7MH21IusUYIOYjpGPyI/lnnnOhwk5zZ/JLS9yCUmKXPslPAU
NkrC/WD/s78/6UzTszu81dTJ3uG+7cT6vqVbN/Jxf1/Z6z2dWor9prQ1v/J8K4qtUXlB+pA8IRQo
AxEN/X4wI9PFQgn5oYs2OkhCXDiJPZi9fZr1xufe1iV6/aOLgptl1uR9w2OTBw9d4UsfbqVZypZc
EGrTcrmkUC1qqjqtIEfBpvsKLcjSBzJa+idRdJ41b6lvts8gLzoVQZvdoM/i0RktnOpJJ0Dk2inI
LTQKVHZvv0ZnMiUU+dY4ViJv0mIBarGnvx7sY1ii6b7qm3UtLEaEO5PA4MUIo/U7jNuvU6v5Oc42
0PQ+kl1A2Yeg2W3ssNA5u05cSEUIWnP5xt1k3myo8obRPTnIgFQFJXvG6HiEnIF+J7I5RwtTLWqR
H2iHlc526WFbrx4YMUG/mKny5UgwLjLx4jpCVMhW9TGXeX2HIOzhmUs8siEDRw29ibqsDuImmWYA
sOs+dpoe0z6OmnAi4o4uL7uK2dVKWiAejkTS54G0KDMTjfWqYhoxDQwnGEfqlUhO1Cp1rlGoW8MS
PgFknu7R4PUQSfGnCTRt+VByOD02OmSCax/cjLr0SQL34DYETJKLEjI/0zUqJHuEfPlzSw7ypmYR
+GpfEwyEaHPv659EUp88lxYE/R6z5rn2fRsf2T+dsOAOocCEY9SPu+t1EHQ7vcT4Q+vHbDVAjuxA
EFGEJEEDb1Ri4hfdhUs600r9bY8HVQHDH6eHp7/mfMrO6abzXHq6SAtU98rAm7QE+MVv5nmuvIxo
y3L+f0Ba7YOYKFPe6z22K7EvC0aU3oMlitJEietadZecwW0PqxQ+GfBtZNoVqicY1TjaeXwOvaVt
+MBAzJrRJhKYtSAfJQzYHDGMMXtPnbCu/wr6iV3oM5KUeGk7RqfuIGCbbb9gwrn6wZBBmnAqA3kn
eyaMARI9JUQeY2//zL+2/pz21eHjM10dgDrn+6GeHzgitbfHuIaR2u/duX9uNwnk8wAHUEDmN/2U
kQOax/SafcpwupgPfrTLsTPJLS365WB24l5aoYPLMObExe9mBqOToFGc6ityMtoqlRAlmie2XjYE
zfStj9uIb7TVgU83z6GHCaNNgSShoGvQY0O4awVY1kTO8Wptbn7UpAm2w9XKOrA40D6BONTmBnLz
G1X/6Rt9BOmoJJBvRUHbwZZPr5ES5UMPYux4ZvdcTa/ogsi5iXFVjdToHKs7UeoAkT0EfEIVTFVJ
zN0l3Kf8rMphVaor82mtq8dKnVgnH4hEpEbWjtL+ly+S6nuXH8uj3FUpe8L4eCQUpipY0tTsRBk/
wbOLvN22DpRBmDhN6TKXldZmpGOZ7YLkgB7PeXmHJGc7A9TIA/TrULwINd+6v9H7JhaQxMXppbS+
zV+i3WSTzuax8cjXbfYJeEgsBJLPqL8HHeZy9ODp1wKztX1onAsEhjiF3Ll8KXO0f43yC5Ev9ZRR
yMljKsAQVYlkm87MJzDSPzj4EQXsQgpP7GIOqxRHlV+RXTE55iLf7upapFHdCc3+dok5FjC+lrWX
zKwNFcS4ZPgvSHzhl7BmKjrTAeSO2nbC94cADJNtUD8gMl7f576hPT9HhS8ngnnINZhL1cmrVePM
9ndfAz6iCJfj/oAigZg5F7v1nygjcKYHgMesVTXNfcmN3IKnip27EPrSquQow8BQVJ2BVQFLU2Qq
vVXQI6fzTgP2ygMLK3i5bnPWhA0Yz37RUTK2vUh5o+W1mQYPz9FdUnwGrKkTa2l1FHFVr0W2Xn1L
0PWDC4sCjPJR0pUiZq2CdRhl+EDDsVNeefFVwl655J02d7wYZEpoppq9wCm7bsKBEomi9gYJt+0S
C0vwnrdW5z3n5tlYAkYPAaR6WqZDB9ZNdXEV0arsM9NlsXGxWpCThyCQHA1gnpMPv9XcLUcRaIZp
knMqVPJsYfbdrZJhmro+KYg1bVduPMNZNKHfylWmk+S5XxfsdSx64BV7fbD0KWqWjp5F7kIT2+3Y
/krsukF3XNHGNJSRvHzkRYh33hnwXhsTdszwxCs7psMoMkl0/h6bIkW1aoSNW/FiHb+zTD7lyIkC
te8eIOrsLdWFSxwTgcwOJ9skK10yKt8Ixy3+aA41mlHLmFfj1NzY8xr5NA78HDYC6sgXhaAaZx9x
2MGe8dJQqotfMGEW9N6OCJtr+WfDLNXuGbI4T7xJ6NPridNrJuyjvE4v/ig1QEKQxniPg1ue56wd
L84icPIdcnFnsSLgEmN4Utx6Eieh/5Xy1eVhlacklxuMu87IHTTNVm6+mqHO5SsPCZdh7ZLiiBrR
U1J4F3CRa2M+bpWj2g6Xrf5bPB72T0SL97we1FNHl13WVt9apYnqSxMYc8pJqCBWdvecBIKWSQdE
MsqmCi9fWzxNCWiRD4ZKQhvilr/oXVivbw8g5UjVKkyZaJlaaI7Ju6+qW3EcPScy35OCs/eShB7X
/XQaUFwbZP8RMa8l0rDDdvWhyKBEVtuT+TbKzXR2Aze8a8G5+GPAi74pI/fFxezhSm6ZNHpl863O
FOwEllqTByaaic3yDFTKrBadrxzaAkOwvzUQov6Yv9Cujs/jp4wmY1o3zQLgyhlYEuhco0Q2r4mV
h9sGfh2oOS+tiByN84uBfDLWIKL3F+nThVwDwW0unBOOGfDyU4AgriP75k8R61pQfYMzQ4hSqDTa
5zpExjO2W2I/N3bZlAhFXbouOMGxIC5DprJxGQUeOHwE6G6sOCwq2z6sN2f1c+fhrlUJKq4bc8bI
q9N/toEumoWCfLG2KaHvJOV4/ksUGV65ZnFX7FJHQuJwGE/cU70pPCGb6ysfqSZh7I6wFMysh276
jjdZOWOa4iapKpeJ65WrTGY4vPnBOarOVAfWH7dKusgt13f3kJkfcuYZPXHEsbJtoUcKkNmAsQ6Z
s8BO65so52XsWDsTx64DlijEyl1OS0l/aYtRbfIejWzbc5+KluXJnAlGP313UoTv0uiO2jamVMdL
M5B3lDlawxS8YKNghOQA4a+calvL3hXjrZYLAFOAW10DeDQEhqoPiM9rschpRCI8YvxNPHhH2PkV
ggScnDp+solxVR0i+XxPfuBOBkX/SZXm53JDDcPYP+6ohnkvhjzUVPpTdmRJbXdQpbKRZl68AM+u
jtw7yI34CK9ioYCNtNl0WAboUJPVZM53CnDrewj/FDCPz59XocyQSYvVb4owEpH+OInxNXuIaoDM
FzXh+myEdjE1jqNF7N9AgDUly70PoKD0anLrqmaxFwIyeyUNrt9K3g2FxncpYL1XO4MIQqQmRnt+
E+X133WOdryoxug9ugFwTpF8UTR28fGf2oBExJ9adWjCjSHkCDJmlm3DhaQMenksNMDLEjCVk1nf
dJJy5MU49QPeTyVCHlLcKPYQJjGIyRj4l5yMOBUiBAQl+oltdApL+cPQdqMPR0C7YaWJcf/r9EBe
761MkYbmZxHfcD3S6s/K1ZYHWYHs7hXijzwp+7FY5Yobpdi3DOE+gUz//U7ZwBGX7tuITOGYxgCJ
hWhJeMgSCu/KVgiBqDBrZP5di55ISxiiyCT6xWyxqp49FjRBVsnFrTpx0hTycqEZZuNEg089tAm9
dxBegvL6dwLfQWx4LsDIw+ANIqqhFGX/qadfr0n8YYhBvoGdXR1zwcBeHg7oJB1fuccGFEuatbsL
BmhDi4uYKVwgM09hDPXF0PEL5oR6H15XRTTK5mRIvV2aVFiW0oNeG/O8b6gsAuyakqeUU9z63ZH6
5bVu45gLuSucSx6It3EsQTAfPuh0PZUIysi1/O1rGhylgEXnUeIp5lK8J8WMIilBaswnl1M8ZZlR
GOY4u7mZSJImf9gquntgYZ8556VtVifgY3CDBxmcCmjTY49joskc44kAKIqcCdQJHBgsvya2yWxw
rYVYl4vZarCialNKmlg8gEDlCfRUgcMzRjdeCHc/P4z+h/BePvaC1FrzzhTFnCL6kZPvccfFZ4Jo
bvieXAThrem981thPEuv4nmPBTjjLeVAm44+ZzWLbK2jcf6/ok4eOr5lHeIGEZtOdlvHk6ZxheMu
DRO+J+dAnSzo75qwuedPGPXoX4UrgJR5Qic+ZNqs0abaWLu5Vn9nZTcT9jGzsWsvn5hP20gbaL9Z
DqJClDpzpLNGZuB5yJDZyIhz51l5aYd4JbOAWZp+lcNgKwYRDZEOdp4MDTuO0LyElpCtq+hO6eek
8LwnJj5EPiEdYGVUuiGd7bWyEtQWgIFFFpvhipdUFLfGHLl/UptJx0c9g/N7w2vOulNfxZzfyLNd
L4e631zkZDeqPaJDoQDemH93XvfNgrh40SvUtaZVvSmpMsvMk8Pgt2NqDO8ZerNW2E+UiUfSR4PM
NVPlhxfYsx078a7136JoOQalPKFgY1ZLWmzP1ZB1vWpGFFJe3IrC2FB64WN9TA963+jfQx2ixpf0
8MqrYdhfw9pPqoLwwqcPF10rYXftBZGWepXOqhCmo7W04W6VSx4TTciYDAdBKWbEfn2hnvLqLSxZ
Ku+BPdoxlCIbOhK+UE2XTcFLOvcojI3mF/lIBHTYveTUOTpHnMk2Xt1xooxxNwOrvX2CqRdsnLUJ
VQSe76IRsy+IuUlpENClSJbTvO1hZyL/noIbwqLL9QLjVBS3bhzvm0ztguTzG+8wEqUIDiyKYkYK
xzHNKx5mYYuGkKIvhyl/lOGoDjdLc9oDlD2Im3ZiCVU/s8qPsVfkbSum/IHLMsAstPH87WAK/jZP
Y4kc2Y045JQh2LZ2XN0X8q4JHo7oKZIwnPZovUXdmtNu4yIXQS5acTUWGDGxqYoMTWUq+IidCCfU
sJ0s5a1XnBprdgcZDaY6CBZDoQavP5Phf2eRR8JEZhr1HOjcAjEhBJb3BnEEqvqaVMcRxSHhAV45
BfdZDD5ILEk5G5sBpzH2ESk8++vIQNolTkOuIPguHeZSualZohLBBamg4EUHFwSEZnBaB0arjJsM
U9d+OJul/6m41IvO1L3CnTLRVktY7N09COSq41jS94hYgFFlnnAq9v6L6w+MZ7fCVGqY4/NfnMrD
7m66UwUi98BNtGecHevNeJB1JYp3NeYbLYdHTMc3WgLZxmmOrvGwkBF5wYzIVPxb51vXgRvUseHK
floongghqM2LbnKY0RdFLdjXO7rXxVLpnKTze5oplTWRBQAV6rlEp8Y+5d1B4IBv4yKUjNSLBwoJ
YUWGr/TbknzzaF5rMHqRGKkLGff88UhMMpxuac7f/gyyFySvAsmX+KtUJcFo0xxx6oKKKN6qptcM
mrmcDPDH3VLCVuR3vQgxwDCMBP0Rys46RuZUbseYjJ3mLePe0AsYYOFvCCw4xGydqPJH4cJIlY/v
2UDeUuXBaV5qvjF3Le0jcTVBdiOpM7FKF+kPhQGBwB9KF9tKkClMbDwfTf91Q86sOkxc1yInS/1y
z4/3hIjie2IYhqXJCwHDTLx4JRUksS+ycFuY1+s4v77hlTapSB97kaN/y0N6DllgQNVJKxadeXwL
A7Iyh/d2CuNTk8NPN17nyJ0eP4r0l0ggAKD5xmtNPb5q1KCQI2bXL+ubZ1w45bEMrP0AzsGIxtxf
5WJgXb4Relnn6BERD6EySMgSls+5ewtfJyQAR6Vk2HfdQIWw+brBGBeSrDnR3jbfsnV+Tft6aaUH
4vXDoB2qAFVmLdaVN6+1s+KynlGr12bDwtE1bqCLbl7o1awRyXaow8US56hHFyhEh1KeSuv7+YzF
S/CZ10KBX5K/qNX/zxK73ZKZWSalEVgpc3FpUbYG+CM2HPpGaSiXshRarvCBQ13DwDFIwtqHAJCQ
b1qziz79xhsArNMyNkW3KtgDXl1U5opETtWVT7NFe+6uwD3xoLEGswy2gV8pMn55jFcsceCVblwR
CrqV6TBnuMJcRlS661d9JxMp6bkwxwuCVQ/GQK4uWYe1yvS5LQvW3aexdUtAe1LHz06HINSOFiN4
vNyLLHCMMsGXZeNWuGs6wzmavsKKK2ZUxFjdC7K5cH47AabGBy6BbPDJvAN8NbjNtorQvA6ZbVZ/
Pmsch3OD58iqpeIe7C56qBaKjHG3HFqERAfDo8CxRNsVJu0UIdMJDoFmLWWLxR4/RB/nZOneGd1f
syw4r/VA/eVsdOSDox403G8riLlOtapobXf2g6UHA5qrDIq0NFYDD0XqA/Cp+w8j2jHsI8c0LVew
z9nE91fo122z9R3JXNmoWfP0ReXLZC1F4plDC7y9IMQR6+X5uK3V7dL9REu3N1TYxOwp3+WK4jf0
gYoFUzsCP/xxC0C7+Qso+uzCbdUcaHAFjjbG4VliPBYSNEzqpk9sii1AaWuIoJFD4WsIW17Gugst
BU5CI+0IY92Vw/P2gJdoGLWhiOl+bnICnEXUJQfr2s/6MWYbtgr5X9wWo8PTGwYvUbcyCEob2CCs
727KfiTMxNB8IQHqgDoGktrkNm5ab4mikRxlq/z9BbXyECjynGVH/z6H7sMyCr/RaBP7cUrEtG4k
KyS6gdGxOAHWCVRoXmCNPnuYzEPTobmiUiC3mkOKUc/VUR/hUkQhZCcC9ijgGgaAmHAO5BaQmFwP
V71kv3YHMJcikc9KIH3pdu4GkniLvVrx7oL78WL4yX2ZFHduqsNaDjh2reZZbKuzVQ5v11ULwVXA
YTnDvFyD7RQVkCWt3EAh3iIHC06Y9Q+rJ1tJAVKi+FSrMoAVDiKb6mM8YOet177+VslXuZkYw9FT
INEetye0VUnQJ4Cnsi7CxXgHGdn64GirlgOJe+yHCH+cFBZXiHn7FCWsGJqeP4eRVVVz96lBSp08
6Y77Zt6HteXx16KzBSyzlXv96yPilBdGMJT2jwbV0Lwgp4apnmcuRPIoJjlrw07d+zTVP0t2APeB
wCHqpDUbfBbUa/VPzmxSEX8dPmke41PTmS3YoZ/qUMXBFgT+2U/xcvePb2vWaITL5TfiU1ydVD0P
VZ1NQyeoG/NdymW+LiV+YeZd9dYFeADbyNjLS0EzWf+jNB/s6CCIo10lGnpZpCdJokPaa2hAx0FM
iff/5wiSTZJwfp64UNJBpgcALYYAWCcmg57PQtdmiuLQi/8llocirZY79hMIdL7pKduycNbHVKob
oqpnho8IAvHzLEo3vBh34x7LNj07B/XRbsBW6nu2uypIrYUwQJvyFym1dZ0CFEhna0tj1esHmP0T
5lYmzCnSwWmjwnXFWj2F5c2CUvKIiviDctV+JHGdOG0T0GGgbFVf4ioXoHv+pVGZDahiXS32GEW5
gxx3L0vjK90+t6emJfyN2hzHoMKCqd23jTUU1OReSgdEc1bgrqf7mWKuuZ0xSxa+R7isM1SSE0Gb
ZHBSFfN/uW0cQEjGJc6SfghldxDKGfxZPKD+I1ked7I4m17KZHcD8bhIDaaU2FYfNuPf8lhgFqUp
g8hYcrMBzs4KLAy6ATBFpP9WLG3W7i96ucW6EzMox8O2eX5/bPTTJGEjLxPJ5YM7m+/BoO081Brd
uijDb3aMwmvdGlbSnimbniCS6o4NeeVjl3mHETC9Djl9uht3mLwUnm+AmyJDbt3BH0Ouf/poBzZq
RcMrZfMI84navWrgCYa8QVkJkM57kcDC5JLPQ1yD4Yw0Zh/TsYsbHhLWk1wnyUoObmDkmpzalfC7
R3UjIjg+2/7/hk89mVCWAt9hSVhLI/o8E10OeLKSxnKrNQArZOPJonmR0FwpiQU6GRhlHmL/zD3y
iDtfgUOvt0se9Onn391ppf//5aMXiDz5T56nKLXY6ntPXTm1mkwqxkxFY6ijBk3Ftpxjy5OpMQsu
YRSsRURk4gex04yefKCoGFq4wFnpsDuLdEyFFlBXGsYw25cs4kjUYwgzGudJhg3FYIQ+JV//BDpR
57q7mA9Ke/ZSdTduj7AGVNl26fTTufUFRQTY8F616Hlp9wGLE1tsuda9Nh02pSCPCo2HZUNM15PR
DMadQIZIE023ZbXfV7rAOO1P5fhY9rOnIR+JFmLTNmURJq8cQDlSpQcyEoZiyYj8BshodlA8SR9P
ass/N67UYt/CLMAOrRwySdpYW9m+/R7zHMqH5/SaBrAWdqen4avBNKJ3OA+yDuf6uQ0OupNDsWQE
1cqqdJZ6ypZsZQ0nO/lzdsivuPhla4EplYYLOSQQ6ltkVmO0/ecn8QVmvIBiSw+d0p3AFWsrLwzL
NQpWt/QzfKtXE577tpgYVWiBOZ5wyistwcfQBt44GVbyTb3C4AeFTFu/Rr8pg7HJl9PIldco/FQ5
jf/M3YPg0luU8e9WXS6Dh+lAPVpuK7fUl3d/xoNOc1ovxPMvX2tsa26tBefxYQ+yvf57vuD8xwYp
ly1UI6z0G7VxqoFLeaPeJj5e6oGgwCcGMBJe3kAFln/lZYULsECOkWobjE7c+QCHvLXJZgjSnYi0
omkgdCwMm17sg38FSDLgTMusX6WZbt4vjBtIB2CQA9qAP2f7prjE7Z3Hlm2W11JrpkaSG/PKChnF
TviMrKEQe6OaZQkQMqdcJGfmhN0IQ7W13iVwNYW+mn973FuMoI7P/HI7/NlsGpgAKfdO7n8bU1Sx
/s3FcaLHFqPZ9INtI8Tjwy0P0ooG1F/iaIUPBYnI8+P8+726rZKQxZnnf17tKz2hm0jBg/lThEY5
F6qhDn7FlPIvsW4RjC6QDTx0R9OZFRUubZk19lslwZPLYJaFTwWXjhGDjb5vzX14a8VuJFZpQutl
AHCMA00VC55HlK1i2oC1JQB1ShUWl89WEsiPjcKt5g0Ogg4//xRpqKEgkqcjV/96xAo8iooDuq8W
kP2iSnuo1zGxP3XOafkQYZBwa3r+/9d/2jSdYa2iknCHS1si4jhFLXuUl+sSwDk3vvg/2W4DCjWH
85gIbCiiUAK2oKnepWg9ogEl4v0Q2mIKChIAz2eN/fxK4RRi+rT75HaJyXnkmeJ2o4SiFyFpeZt7
+B0qvu4RP6+bRu5Kq1SuKSaMRNUQ3neNZogQilOFo6vf58U6xWLrCk2j2JaLzaB4BwyS6F0/v4yB
Z3B/K3ylqvAsCLwzAYS3DfFJHXWoTR+3bbh5NtoH2QCVscP3gZ6t+TZsFOfrTYvpCza0Lv709FHy
TVvSGG80TBsru1SNbp0eMjYd4qPEDNbpKdR++KkU230YSEPW+tVGz2OWVs+uIU2c1dJfSSZFjN3m
wHM2xDRPLYkwU8guVc20fS1sq8bsI/DyNI5VmW8Tvcn6Lo/7R4VBemKv5MLDKYgWpbvJohY0Utji
KoqxNq/lImU37HJPLn8emSaRiyrggQeHBfghqCUBc6iioEiX2jTeGcMYj+F+vDPoZBES/sE78fx8
887nILr766KjCUomLaVmc0QIaoazZPWbPbDOgWL0gdNsVVR5vK1HvMIcDAK6LmO0sXjzLeA0Yl7U
7e2aiRJdwu3oiZNiIK748DzoS+Vjg2Zgoefj5EPnpAGV7mtzcCp8Ux7IiQw15563WkoLFedallg1
Vt9flpNbc/zehKYJHbjjNpnLpSRTMtnxDZx7OW1nqkPz5vTwXbUL2sqr1NaZvK7L9x2xq7TFi5lu
dvoRpFlC1EO6JIbUuBXts+2RdFMM3rLzH/eLHa9M38LLaH6dfix4TNWZyzYz16vGCArmismG3JQX
B99x5mkkbuAvSV52snzAhx5TS7EJNFxvuf+WgTvV379RmibWSthtI/rf7ah259mV/4OFO+DGI1fr
LXWbQVqiNd71+Q8HI2G3M727/8q6jlCEBuIt5BIOI+sV9ij7UCrad2oDVDfpBksFVJixAEPABsuz
wzYKJLmk6G5OLwBOD0u7O1gV4HwyhJjjM3bG7VYll/tg4cK6ZEDTY4f/2DQHMpDQo/l77fnzw2lG
m1wrmYc/a4s8jZDy19hNCjWEtpAWrlVQgOm0vpobO18+GKoqdEZF00biN78VTy0VF5LiKOTB3j0O
UNj2uS1ag+9hMTzxbW0RDzQwBu0stxo6X/SRDkG1xPBD7Xl6k30O8qKYRnKJDDsA5yHM+qyH3N4w
aekzW2TQOPQRUz9zBWMOOq8va2ndfNpmcUpugCIcFp7GSogNpE3Q+08e5ozmpdY49Oxj4iIbL4Qs
blh+IFmxbHUcbx099mx6WrXePlgkUcyPxuEF6XFK1+owSre8zcsQsbQYhBFCiLGmwZ5d4n5mXU5f
5Y8dq567jXOnojj+MFWo7UWb+QxkgAhANnXkLXRPAK59y1gCS3zwd34O1BrGJ8HjAimUtvfoEU7E
O1McsMMS/rBuI24WxWTtyoRYrZfreSu2IVMvm4n5ymLAuqR3G4jZNKNwxjhBbtqFX+FHF33G57xT
EHUpshBjoe8HNc7avolDXo7QGddfCSTdHu6KC7EaJ9B34Lkcm0uXQZ4iTFTdfPrSW9N5SM42IzF8
bu17IwyQZslykv2LDS8zaUAqxU9tkckMOc8b3VzJp0UvU96ozu2q6UrTPeOSgM5xJrXhL7Ns8Gbb
43434fwO9YWQsM8Aj8mUjQVxKJ/BEw8S1Ew9Qb6eMAktS/PXu0Cv3lTyiFydJEfzxv6Grk7naX2Z
yjQmtkXzyuUB+5EqL7VmRKYAKA7A/YDhX1Z1o6TqcvpdeB3/EhTxrx0lkADS7TiZ47hpTXkJDlSL
OSvQdodgAXeXAerxkC96kEZymMzGRkPImdjmNftcXiVeeKx9aGLfxN25mxNP2lq/jxzQphGTDLIP
HCgVvbiI+N4WnI/enC+PMJL9ZGNNPC8h0l+rq+h8vwe3crEkDTEL9AocHu8ZUM2LMa38TJTx9di+
ZmuTQvjCtQyW6Vi13SOazcD8ah2rrzReM5Jcbk/cPAIyS2i5zTLjWfKLwPGOAIJipMwouiJ3AlNq
OKeq5NuHTnJLxiBqbYqu3TrOIseQXDKSCC6Y9Ud3qNs/5H2Wx03YSsEf/y7BXJIdUDiS/wg5yI6V
z4qqsIBKkOWwqjlrFca9/jCx8rOKYIjn6ozFMH5Xcz3UXXkSHWgeJiU6hmOLxeE46d+q/2e9IfN9
efEOIA7feeHGuPWBnm2UGsDds+PfXtfUmBurU/zaIbxSv6BfcIGIy1c39DSvejkiRyXBb6kuYy8Q
QhHY8px4g+EEmnro7mFyrfCr79Jy1ptWmC6S6sTidUvxJTAK8T6En+xLLq2FQGYVkc6JuyWJ1doy
GW/HdumYUKkgMWa6+J7TFrG1UjCRM4h+Z6soLAXPE7FZYJYmnXgi/hhwKUJsZIDWfkt9A19f/pBI
KwrnE6pRvZCIqlgyv7aXRRhkaRhlbgxdEbqaE0P/UohtQ64JqMAmrcDp7NZG8Xj6lxwFv0kxJOsT
HbCBng/KpWkuOfvlfN8/b7whDOQwXYn4IFxRnqe1aSq14ZJtoriFniKaCBQG1QsoXarK6yrlRuh2
c0jTykCy15v0R2ILljclbIkGaGRDx3CmjBsmfbsv6Nz6YHbGx1ugBr5onkrPYFtkAO2yUXsWOClF
2O2ZlgXZSZRGeOPBK8M38v/tAN3tK6VwmFeX6lFTnTApu9qfIawLQlQWwtEE3XQ9pXcGbJ9Um5rf
h/zHQPEkK9CHN8xWQtAJ/LmW63yxA2QsVBJpc2JhScWNIh2GwY+6lkibgjZc4yiB4ZEodLtjzkwT
8OQE8qsWu82FqEecLN1EtGNkhrM44t9J+drOazgmw0NauR1IMKbGbOEudiVrfkogT71t6X+PbtYe
NHIFfqmmCA2ZtmxxTcqz4rwTqjJw+T62NhWZyOKmP+9xXTAaZwmD1CMjF/cyNj4zAHTS2x2QsoPK
z6JdJCR/Fw0xqKk4BybKg0vc95Rlv9FBiam4aQgDzlD2WAAeEEmdqtI4b+E/6IEJVd1OJ3C0FRln
xUBNX12DWofx3ikN800YN3SmYi43P6O/CknFtPcZ4h5iqa0nROm5W0IYfuMvB633hOjoR2uufM37
jonDzXEjKkYiF+DBzPOX7Ekd23mogAZ9NPcfpAUiLTONPTShBZzRVftiYkPK6lCJzQSa2HuP6ipm
fR8BoVRv51CMpAtFGjezogmGAKcTc6HHqt+jLaL3xN0Bhge6C04jVmj1W37d99iP+PgtOWbQQsZg
gJ2TcEvJ/ZqBgCEZGJMtPWdJrnjDbzI3j00Yq28VHrhkyoAx25YUA9xXK343tmM4+bv0k9feXDOJ
N5f9LZPr6kOhfz4bHJ4MRLTjzVLzRx1f0jkRmoT78/zpB532ZjIZGiaElO8zpt2VTGHWje17H46w
EivHbGi1N/tENpEOrjHhiJtYn95N3CJj0lpFZdZwpqamx7Iz1kLhnUdS0DJ+kAGdHKkDLxLXO5eD
MrBep7JQV4q5Gj+yqsQLpVVzC1Zw8J6efUOtD3QBf9yDIZhJS+Dgw58QB5k1le3BGkGa/7sHPkhP
uh/2DDrJt6iTSJSmzDkI5XY7yqC+3vCEpZ5nCUpiqCSyf8U//YqJUEGm7MWpY6kujHrgT6wDLG0b
suqIFlTv4kYWnTAuTHch3cRxKnP1GrTWLAeUKed9EXlzV2/ZE/fTvtwcHac6H57bpyzmqSFLQkYh
ewjQd7DZk06ar70sq5Udd/OtVyBXoP82aAm3zY1LwTeCq7HgsTkSMNqaFi0D+YRBXK6xEpGde5rc
MnPrg+z/suR2h/4uSVWiRExvsDRu9RVU0kjAoYbxKTtkzdR182dA4ZyIulz3yKqiQLI/4ate2SyJ
sAzfDVBCCAjMPtLAMGJRNSIrMF8TARiHBGHCi3BaG7RgT/IAz4qC+I3RHQ7WuJgziukpxUl0fsq2
LjeS+HmTscXPUgZWGNsUMXKoYDyR0WTjUlS6zKwoeZ+Qo0RqWBgre/XON8ktgB/z365RQ5u4LceD
K1DhL93RtCiw5UHir42vB5fV24eoXzYfgtE5tYyWCRnjJLkzvokLRiNTpY1JyoBXQg5P5bvLmrKS
vfsX84pbdmkyYqIUTLwJsOPnesyITsUz1/TkvTJ7Kc3OrTGttvsTZsJ0/XB2Cy8nqytb7f3O6cVc
+1gwz6gntn9UwsrLRRaLagWTiTRKD+q8BVf6Id8/YnXwdld/x8uBjFAxDy9yy9vYyeg7Rq6RzisH
BlrUr9bI/x4ykqZW2tXa5C0PLkFFCIhWro+MvF7dN083ydu/IgN7BkWc9bAxAalzLujU9v87GZYa
TUiK7wWMw31XqM38fBS9t+by+fmeWreGxYWbBIfwl0bwXjMEHdJ0YFH1XcrmB7hoRSYlOfCcxaCn
7KgU9B45mOaG5BQIpFldAjTprJCxxEo8yYRBJetvijIzeUTk/aCoVYstgq4EMCCKPULZ4bM6cXXS
FpawPjWDWDp6SI5e4LuA19DQsLxY3dNJOfFbuZBMRPtJfr50v5wtFw+N601CJ7CYFxBQIxy1sny9
VR8h/PuHzWhCEA/sdEYpeP6B9tp9xzfjDtCgrmEKCwhMRNaRjJrICBIC0mCH6vV8So3KA+6O3Nsf
zWk+mtYw2vGWl6aZTckogCDS3zkRMt54d61jh/aEdmzl3rEZ2096NfMSdvBBpjbdVE3lnMYn3y3k
GPzYRhSeK1HHeDpGD1Yfq9Dm8w6WPAA6cTzZQeOTMH46X5u6C5Ty30T0/FMGDmgfNkDUqaqSIfSb
44nKh7ftRchyZTx95F/DS573/X0jprA0AFumPWqvia49buBeC/6c3+7ruT8cQHED/leNg82Z63Xd
wsEzOZdOd4BnEQ021MKTp30XOJuRAE2L8tVV3wF1HpznnL/dHYYFCaxDpVpNhk7KqDCDBWte/8xF
9b+P5YtjC0/oDREtITF/Ny5aW88MwLTOTfX4fIgUZDzHJcPjNz9CcaHb/z9nhFFP3IH20E6wim7X
VsaB5X8/NMzUGlEW7dKLZkJmEdDpkWFU6y+8eLz4kCeoNZFBn04Aheat15ABsxRNQubHuv4hN4xP
0kx8YjSVRy+Oz+giJmdg+nSU4BUIb887QCgqnauU3mdDPGG0EKfyljXQYd0bUKfrFfpE+gC1C7DO
1cg8h5kePf4dRrz729Wi7QCdP2LPNwM0XBH4xgdZNRgUO0WnS+hzIGJU4k6JBLmArQhMH/EmljP6
8o9acvvFzpGWSMmkYsNABFL7B6UwMmqnmkS/Tfn3TMfTSFXc5nuRnTy/JCIVXadQsPb+J9tglxwR
qx9xQtOs6/G84dlA+c2TryKuB/x7AKvXeZPHFDD2GVFCr4paaWpuP1PKrJdAgDcG+R58b0yBImOw
lBUUX7Qszwwo7gGeW7hlPVK2RjIGd4e9BdOiDabPzKA8PtS9AkcDYGcrpLKHIx3gxADi1cHaqeRR
B9c+462G6E7YfZGmjOTK7xAiyRueOWGc1bBegVu0y58Xcqp6sqCjUGh/GgkinQC0kEyGHmBGG8rr
c+cxWIDm3bxbllDylCktP5PfihXkCchUpqiD+r5EUrreFstAUSAwP9oRWbaHZCTgQBCtHnmzengm
edjl+xjMe/CITQHQRrK3FoHLzNu1GfAMG7fHfATVfwahFwtDeA6OBjzNllW5C8W9/1JUQijAZ4cn
tBn6LL1GyyaWLPG9NT/IxY8PDeNJJRsQN+V75ykB8qRGj8iDvMkRF5LpJtjDksqYE3FRdWhrnowp
hFXzMO8Nm8mb3M2+iW9moVcYE7T9LGQyGBht9x/OWDBwf5v6JkdrUXYoy7EFSVBxqSaaMadjWyBs
uRv7wpThcYwyKrDLEezNEX5n+P4dokFc5iq3QPgIwrCxBLWuXiCBrGAJeKIwORTtNnIeWED0C6IR
Y1b6XFC0wag13u0peQMc3FujZphHJZE0roT+VE218w7VoOLp2ZyXYt6Mh0gygSHeJkh5KD3OBiD9
ZQ77+nzJEhoqGeolSL+lUwvRYCoKtEgasKubLYBTFUU0rK+6r2PQFDspF6j3Po6lxV/U6fCTR1as
xEyN2MlZp1A3OZYbDqJ9CUrtysiA74k2JQaYuvP3vCPGiQ9iE9rkLmCnWmkX4UpiUFxwJdWYSvDK
GHrMROQUoX8bJR4NLh4NSvGHktfx0gm3Zai2UweexZBOcAPKevt/vmZR+qAMoqhSC2DZnycOfx8A
Ev1JgcrJucc8yyoxrxtXnnDrZpG4QNxwCQ0LpniOD082WZ5IuBhhPPaAT09Uxl/NGZ5jkPPk20UF
oZgl4TA4pxJbZHWyvxKtRGIqQjpVNkOUjOjVKn08jOB3A+SiOAO6FdiqwbzGX03yR9LkAxGPDiLr
SEIf1zVlgDxtiYwfAUeppzfPRQL+KoIqVvX7Dc+7O754G8ztXr6CP9JXletiXoDE5hISGBVGx0Cv
xKh6zBblyLQz2QkIG8Ry5chuXdWyNMYqYrnkMx8mZjngIKQChwVPken3TRMET1OeOwTWPJ5W3+m9
Affz0j+jrRgwXfm7W3gn4/eelckBWmz5QjuFrJ4XlFb0szfN/ciSu4fkJZKGyK3ABrNvk8VevFMH
unN0bCanfa7DWW7BrSkkh1GXLHfpqeaCw589zekAK9W4VlrfTqYbarPLMFEXvDwGg0V9oerwsTDu
Jvce1w3AcdZ7IlLIwG2ddxtALX2fJAOyGXK7XpnO9duvST8hGDfdEL7cEpRU2duSlNbE72Iooza5
+lM2TghKZDw9Gygu/ZTyf59qihJIppuWCykKLJbitbB22UHq6iFZJgHbGELNhqEPu6FS9x3HSAgY
dccWaN0Y7X/cm27Vkzi3U8uIa5ionAvHLEqfeCOrcp7cYC4iWHIkBxeoP1/MSPOxS+CT+d8F60LT
JszgOIaUSoaONhK6Daan7NRf9r7/TutQZ8QT0WXSR4bdExDBVbm8G+jGKQVvkJ372mn6oYB30eTP
OMVoqVqUS75Rmz432I/nuyw0zxIoxC5Ism27mjvXICqow4F3LH0e1RIVrt44cL2cD3qvO0nsSkOX
yue0IRaNA4leKtUzcmDNsUTWMUOVZt2gszXKp4pWBMmYwnEUfj3ResQ1C9JkypipE6WAJIp568Mo
PiZqPu3NnfFVo7BEf0WWfnel5sJz2MQrACM4i6VlIig+3w/paXYPv61UvmmDd6Dqmgis/qZNyxpG
yN4OZz9RTDvfxiY1g4EooyfYFvU7AhtyMc22E7MUeKJj4kqvzLB5utgiXYzkbbVBMQRwVXaLUQyp
m4ZBA2f3NnsyEXXiA4C19NV7LHTY2J+4ViiE0OaJBBM2FS1qMdDHgLDJ1YqA8l+IsTGGJ7fMl405
ELjL1FcT0+h7MeaTOkvgcf1ODshy4I1uwHIIXi/I8kL4HFtcgsH/hfWDcKxCE0WnGTSGkiJHAtR4
u+c3kuF3YsD9UNCtikimQ70ph6bC+ZaofGHSOPh5/tbytQd3njw2Jeke6YtlCK9who0G1yOaPmqs
kGd7Zaxm2qRYq4u/OKDIdDPS0/zM+CdpH/B4EPdbY964bVe/uMZrrx/czWuparP+ZWSNSTzcLvzw
btSy6I1aknxMqFd8vU+P6QmTV7GJ2tM1S1L1MeVh1C5A+pPDBO1Y31exLc0CwWNE/VvquPmaAthN
opkRxdQTD/vYhBQtz9EzgDgieVWCn2DdyQjHHKs/ob31LCNskXEY6cmO8YWzc+JKgo5o6NSSl9Do
o8t9ZL+Duo9jVUCEHabLXuB3F5hxmbtl35/rLZz0H02w1CYeYrcRVXaQeS6bxi2Sdf8IhaDqgcfz
RVz8nO8ZV8CiR+P/kYQ65udUfaauZY8xc93BjFyxEjrv4Tqxbw7Em0puhz0CmrU+gaJX5zzMjkxe
fKxJaYFbDLjJKiIdXB2ydRi8KNlH4Z7nx6c1vhHzKvxK3pwm7Cjc2zbRfpz5x5qht8b8Tw/PxOSh
Ya4PqC7UXugI/Oie2Z/KsbXJQXU9zEvoiE/36JRDuRtHCXeeLaQVYkZtBVdZOQyJFCnM0a8fI2+o
RJ0QkOFHruwi36FlEJOwqQj2EMDNyB4QbIHnPPuEekB6WNSS6Vu7lP5DSNPMVT/3P2dST0NAMO4P
76OffcJhGfSz0eVAwUauvzQy5gAZ2Nts1sJ0sFu7Iqct/dWdVhPHCtgzPj+yNYcJrkxxCSmrm/GH
ZevF+e27q0ThuC4XO+tbLUNu2j1tE1jvmYNTAveUQNMBHqN2mGHLp2z1yE2CKmkVBkLfBAgvU5VG
8DSmMhlPP5JrcS/lp7/hRhPWAJVTMh2/BJ/StlNzKK6r91G0vV6B9gtv5bFmR6rvuA5W7FzWLWKQ
DNNgVs1WKTNm4256XE+u0DkP3cSds2F7HcOD0AGLuUapeiSOPDOEmCKZzorkORhUwrQhDoadrI4r
BSXtQ4EHJ7Zmx3TYw/L8XJ+9x9CB+OKFPNZ0dr9ylEQql4L7/cb6B6P9S7AYm0PkRZud8HYZylt0
mhB/CdGBWBVYHik3dRUFnKlQaspvzFY6Qt0Yjq8mO/jGbgbFWNTLqOwW/s2iipygYXlxk5wrzLCR
xNWKE5bB+2ptTqRxc6vE/OIzx0O4fqkD+pgz/5qot9cb55dubMfl0m+PxBXwwL+RFp7P55kmSHub
0dt+hi4o3Ve9RbOv10AES0INa5z9WrSVmsedyA4CTreRIjbXHbFKL1G+MyFpqUQC9Vh5cBQqDI4O
WGn35cdHWIxMbpN34x/J/yJMUYJX9bdFhrLIfM7WtUTWNQ8lJNkWKozzsbFVOJ6VdDDtHiXkcpu2
053fkAu/c++oui9zHmMr6nzUK0cJbbw2VwhUY+b70GIyh1if68bjtkXLK+mJlHeJZtuLcJQYjru9
CDDn3oBeiJotsco5q8egvVF3npGiHCVCWkqNoqymUSe5yH7O88khO0pyxsu8eS1J8Xko3bE7IJ4M
DrQrm1bY42etPMGETiKFnfS4jM+bfWaGxEBc2R+HXTedCQeWPYoM95+rzQ+csdZPFHYWfUlihT/3
9bLvktUuxGGxTHEcb34xHLXeckyKDgQ+v0T0yv9lKdYUmI9c0y3ehiKLJBHsryhVIrYu7YVLeOrR
Qp0VOZHnXF6Cd+mzXR95tuIozS+GWTzLmSvR7PdjgI2aZJTJc21ruOEE49YcQrekXsZghba/eb3Z
cJSyZ+l1WlzOzH2Ihv9hfW6Ifl/9uVTl0a40aG+kKwg3qRDFwkvAq9fbIGDYaW2dNV7Rf2TiGvm4
xJx5Tk2JjplQU7oQeMWp0WGpzPZdAcVtZ/y1IzSiuL7SP2S8pHYpIEp6xgfaXrr8dHeNnwKoLpDC
oGmt9gGGo8nbokQ4KlkXBssMhZDfp+jaWzXMIovMSqdW98k9W/9qyxrSrZRoYoj1x1008eP8o2tR
Vd9ZhmmFqFucEgJD8f+s9zgQzvqdMBY6Qhp/kQZ8shGaphoA4QvXEJ01CI0oQhL5flsHZuiI8Grr
GOJQeTvC2V1LCOysRi2xM9oyonMKTvkLfni4NzGfTVwPQSheA1AnSO4hFrJjj0TVRZJgyCVIo6MU
WvA8qhZZYXv+jCT8WI9VXqfvUGz9y5jGyu/5/BE8zbWT+k/o1Eql5ICnsmSfCr0PS3OxK3OQA7u3
gUrfQhSahDVcU26zcUgrs6xI+IjrzvD7Qe4yBxwmpmayYuMvXPlJ8xHK7IhJm0Rbabnawucn2Jyw
YOCEDoPwWXIaxC/kycgGAQFN0ZPnzAbvtJDiHRlpdmwpORdaHPLgDN39vYpQmttPOXO66DEOGAxb
tjaTRlFNbsBxKvMIHPWp/YAyL2Vs4+tLxwxi025bY3p4wS+xF2vTBwgx8YRLqMWbls5mPrhfCGP6
aopC+Ok7Xvt3NpGkGxQm/OKqJxfhZCTvt6QLcVLGXjRDT7m9J8subCJXvSWTaSwQho/spUvdLWC0
yeFO1V5Bc/XDeGOIkaPYwosqAHGC9ty0cqhD67MSJTa45CLxpm53jVH4WJlHiFqChl/aH9d3V7+n
iDWG7cVXh2KyK5CctTa/W4WNh2e0wR5d0tPJfQC6agiDOTMtIuyZ9Oji9+Ox+1glONinDeHoWk7V
ptrGbd/V0tzvLuUNeRj4jGtGcTX0P8RXXLQEjLub4eE/ZBCGt4Zi4QY3WQgQ0exlzSt0QKexa+JK
u6Sa8b39Dt9jzSJ+onJOBuQzXQgcjnx6cvMcl6peT2RRxQcfcgBoDTiuX8v64dsoL+7+Wnr53QTv
zOqQuVrf7hDUNv8Z9z4ld1tNHu0lnmOd8skatSvo8ZoDW9wzYYEz1aa6cGtX3nY8MIbrXAZMGYnG
lI/l8KAyws3orsya2pCqOCTTn/530m9/twdJ75c6Z4H0aPx43bvOuhU8WYUHnkYkytjs+wNySIsG
7lDB6VsiWQ1qc+q2YJ41p+vFXOqzdOpm1y5FNyGeucHmdxP7QNSzppDJLk9xcp6LAq4SX3RBXpR2
W9waij7qY0Vx+hAp/wYHxIgW1kSaSdFvhvtRPuDdJqS+xEqtbQ7BULSDPH7gt881HSp/MDw8aqDo
HjjcekV9IJ9ThWOdcjhtQo4ROn9NF1VCYfWBBnTbdyW9XmLAihyQYCVI4QL+AOg/MApjrBR6MaMc
Gbs41o7jnW/QYBNmTYZI8U4xz9BeiB+JshnmeJyeFSekHlDo6PMTywyFou9FF85WnVqgH9BecaoH
hKOOjFFDeus9PcyMLHnAKtuNz3Ijwr6dATBz0mZvHuQDrpgWVtjfgDss+P9aLHhzAEH3l1k27hfI
MoK6v/sBWgMADEFdqumiYWcCuNjHrWdvIjT3Ch61yP3oKf15dAt8zCyDn7cJMf89Y6FvrVDILIjv
+INPPMRjcwZpFVlabenGLQ2pZdwXMXXY6RU+b+SOs1ModQCyM94Onw+kqFXCjNWnhiEPVMcJtduU
B37H2cxNcnI+XNSoEZtTLNAr3gsJ/HurV1pM3eQneSnIhd/JN8KabR3MKUMZKSMk1aJZfrqV2D4t
lKlf3/mil5VwIkhR5SkeF6AifzyuXZ7JZ+ISI1O3L2cj81PoL6+Wpyhn0q5Uh92ZSoL1hyoTD3RC
zb3WP1PEDbfENho9fw7nZA4J/S7ef1W9HPrCDGJj0al8ESSJeRvOcKJdLoLZXrrCm81mvAfBHj8k
T9WHyW25CvF94/iUATuEZpsUrLFxLqcWbOAP8hp8Zrro+tIzZFIUpEJGiJuPQ40vJuumlD03U+Nd
ym+GF3m57qyhWGHO2W1dLlqbIozfidyMKkLm/H1Qj2TSs33JkJ6Gh1Aj266+d+VBxAFaECMmH6Ah
u5NJeHdtjcDIiIO7pht1Yba8LtluaOKi5HMK3LS58jmSqbIW/KtZcqJCEUMVMGitKLJDvjCZC6AM
j2SVXDeW0ZyrVshCq+IirP+b1GBgAlOlCuLK7xbzrCfiVgqbTX38R9uo4DfQZ5A63bA2q18BxASS
w9pjUVe+1NXEsFylkxUcWCrHMF32Z5jqIo3lcLEjgYYUQkUs3uwqvUwICg56nfVoyxkInGvBBBzh
GFwb1zDc9ANN0imcQUKAFi+aCmNSZ/IYKfxqZI8/UkaYUGIqVsPfpndegAUbonOoNz/7ZLS9ZSYH
WwFXT14Lk98FE5Ymvo506QPS5OgSDUfyOg71UV8qHKY1yYpGcdXlz6bPvZlBYAg6//A8GKSfo0/W
+zxXr/meOmz/yvFlaJML50M/4Uq28cJy6bw7dxuhoWuvLrgxTiKC96Fwb7jFaPTWknK115azu8SF
Z6OM5D4wbtSlFxOHE6Saiv7rUXbExbm6OqlRkqbSrhZK03xNapXUr97YsxYp+K4MrX67EdJKq3vD
IdRhYKpPdlf0jDqP0r0e2t5vK9J/1r4kqOXZx07ys+f0MtXv1U8SApheXxPynxzOOtGpS+qD7jke
bT7VKuZVT9e8snXdJEiKcZwjPyWk+gzMwJRH3rHfofG8C7zL0kLgZ5qAhXrQ4Yi+LMfXcTGmb8vx
enxg7E1Mq75DJagIU9Evc6N8OuZGBaazXFb2DSDh7byC7Hsk68sCmuq/m0fB/4XE4ButdIpVFDVT
IKT/L6KixQ0WfI3AIThXH7Q5z0jbhgfoXFp9dD5C25/gCOpuZ0MC7US+PDtDqMcSzc7abYLLsOqx
oV5zflnF+XTry/nULonQmeI3mYcXSZAO5Nu8axXnv4AdQIL5tlqa6th4cn8UMVXZarUe4STpMMES
n+EpEDBdTrrVHBsbAhaIriJaJVQwLg9jmGp1z+tD0MWV+XtyYx72jPOSyBNZFsbMg0xk4TnShDOH
84sP6C0OB2PeXZbno2hyZSp3hrGF5iUk2VQETKtBWYb4szxUWBNq8B0xIMhPOJn4d6BPoPO9y00N
EIPCZEvxY0Xul7RpWFzqZYxJWNb2EJ36LKvR7uKvyBthxFDZu/Fvp2rwQvP+rwdW5kTFSsHdsZVg
gQ5yiTlLxNQ1Y6t1O6JVV0tG9Ct183d7b0IP89uQZpszUIHZ6J8FgAoKMR1KC8lMk4dTg3OkPVXu
zpIbQuNCDDyqcrjT+bDweMbGv1GUP6x64ZBZgJHW+dpS/cy8E+d0A0eEQfsNAI/6EkVvTxCw9CcD
QzohVj9KO5cNLBPtBn3blR5uTZCj72LJjk8GNKFX4+Etx+F5FRbODkozROj0bkGgQrcU7YfZknF8
m5Bvj1vHKZs3ZEK/9V0bpDwTPuW+tXp7+tz7+F9DaSDH0t8ozeb+7PBCsTxch4fJ9zC2NAo/lRsu
QE3jNhJVDPCbwccJwfwVLDtM3ztgBeFeXSbAR2Xuy+NH8eR1icfBTHsQTazRYUFacB9RNx6cRXoJ
H7wL948rEwEkxdROlX6PpnJ2DpA1XK+RsdBIjrISCamAX2/n2rXXh1vl98TOG/FkwpzPunrbN/2Q
ocR0Y9qacWwMMIi4jneoz92fvUe2yLlDpHIdr5mZtiVT5+Ay/XErrfAvdXnnFOLz6YnbJEEgOLeh
fDUMVNoMcn6rY3htq+X93u22G8s8e8322ZQEL6iGwtEfDp8/m45WxNGPGe6se4zX/J0BS0DnI6rb
OVmRcMPtEDYaL4x/rGrXCLgugEKxFaSdqLsjCVH1AdvpLybV44rwO525MnjdhxrWavfGLuegykLd
cC9pju+psxFQ6LaAP9HMKARWKyapzrdYdYgVTvvsaDON3fAA5BR4994lPagDH7tJW1iv2M2VjKLi
CtYdw7dRojXDwws4qOYBSDQiOBt0zNirP5pWCZnCa9iLihev3DGjJIY9COxtree9j3+wiZaQrg6o
QROjZoAscgLsjqoqB04lEljvjB2ob9JK9W+yPclRSXltqZHSMWTaZWdxDsg1gKGmcLDqYM0n1J5F
2RX+o9xa0h1jaTzTSAOVBdvQmeYRdqbIGeJIWIG5DGbYtbfWaxTVpoy8QOd2fUvolNFXTWypZRcY
OuNzA0jjK+LF5kslZbHCpe8zQ+HX7ltSF8Hq8gjiMU6SJxS2sGgA0coCb7m4cxiQSNqmo9fWMeGY
Mc2si/0ImExszTnEtHV07ps8JxatpCZmmt7wB4BNcroiEFVIz30RtNrF6MkwuwPynSBGaTUvWWAy
p9mlq98AJMJEM0rbcvgX+gWVP8iKTcROfaW2kdnF94zqjYhoKSg6mNz/LiPiFtVWDyw9dURLZU73
AAu1C2pcpdOv7OgQrT0QDPQ9M4AaZCWushSJ8A/N8tyrWKn6za0rM+lLMuHQ4lhFo6PjFjMHhvOQ
0LFIaCCTtf+TVSgGQ/4D7CFUJ+aSe+dLfxyB27dSGRpXLWz6QKvEEOqq7TgMPodYwGz7m22ogKYv
ULFSeTQ4Sldo94s0AKOlKnDpcDXp1RWRGg4KV2HeJ4wOBh8bMqyIOH5nihJ6dhkJ/QPNXM4Jc4F5
/eTR1vi+UzmpmCN2fVzdfR3wChHpv8WtZuGZFGUCg3HnI058ClU8baOqELOTbGPiT3VcnLMGrBHb
t9rFH0l3iX/TKFogiHnvMUTEDr8192LMmcy+qVKVvsRxG6eZNeGlnDVVojS0fXqMVORcr4ZHkEG9
R9tR0d+USTw+tDD9jLhBfB+frmgYNuEVHF3AjKZrCrsYFb00+nyeWetVRAP9yND5Tji9nx6IV3g0
9lYOUjDD04ha6jqmgm+DtR5CSrR5gUAT2FvhMHD0Us3LWTkuXDzfcW4CHrsgp9tPZk9i1ONTqvri
IueP+4hFLbhGz91WctDnK2v09NA9SwjB3H1AJZrYieHSqud7D8N7BfwGKqFtiZZoNXLh4azTcq2S
2/5VW2eRggTbC4HhrjPV8irs6CTEjBsuWiuiijto8ZYPzyPG4lyGHWjg7T7qVssHYKmB6s6bfK48
/GtQbAc6DLnDgSrEnpWCHT1gIYYCF+YKTAENDvnK239yno2PNCAyvTgY8xyE/xJwvCrcWcr9CKzc
0VWzlIQ8GAR6FOcylfpzD5W90V+qFwOFDdVlriWMte9zelA7AZTAHd98SWGwTwrOWfRZ+HmUuQlm
uo5ssEKtR2VLohk5z1G2H1EMgBfMyIsSB3Boe4KnX458A2lEUOzLNt69YQzmR7tTGOISq4RVg8Vi
fVV2jJGMvlkUVC4vioIPkBQdAqsvQInsNUeBIJBQdjEQW283qJZ6tPUwuLWZtOC4eTGxMd9o4ScF
aklTPde+6twi3g3zB3ZwkXBMw7FFm7//uvSWtqiGYINCOfIHGtzT2rRMx5AHQGwwO8BosKrIG0vE
RD9nQfeSgKLTrKR0R+pmRI6XFDvaPvIsuCBnCNlkE6YS5qG+u/Px2M1RzZYdYWLRg5v2Fn7vx36c
bj5CCLFvmDDQq2jMBtT15c3+4BxUWl/z5vHhqDC6QNY4bi+7hpQhIzVmDreLhp9U98yy2xBDwVaA
6DT9pgXt6A3RlJ5Z529H/KapYkioVHRDewT4qYJi6QGXQ70h/krDJmjuFlTb2TxrXyrSRXXF4Vhi
RsH5cj8b9XD6fL/orwWS80WGvUTr1CtfNYzlpR7TCIw6MRm1tND8rblfEbAudYGcflMOJ42r28kW
WB5B1ZJXeG/Sz5CLSk6zhVvN9PA8MaBDm6Pks9RgyOZQMM0uB9G5wZb4DDeYtH5cpLvDWXRCm5VA
jrUmzMuyX4BPOSauh5reNsBBrWz995CfjDW4axEQ3dbw2lDaUf4H8zdjjZBan4tEbOymh+Rn6iow
TnOE/LEFXsuWKmCBiVKTmprjDp4jH8uG5w090e1XQzmBoFtvqlUnf3A6+kbQzCWfywLDnuy1Fgw5
HiujxtqAJxGCNiib0gfq1TnIc/f+xQKabPaNj17hpIyiEp9wDXi3w/7xIte9sXzIT/5j9PvWF7gk
Yht3du9N4W7NHly9/nhcv0pjmKM0LzTn1AiZm+UN06ZZ0eyp3mNOx4o0Ix6UYwvMz2G1shvJyG1l
n9434cHryo0oP6fyv8YYG5egsTt2XpPKhdzwwTRK4hNhcwjoJ5hpZDcnOy3zLuVQRszD/PpVAOLj
te+AShhHe5zFaunGsCp8PUNprt2taftbt+JvpsCWEDj3ndvpSeA62XE7WbRe2gtEfg63cDRcNZd8
MFy9kD9x1+LZUczyolMQsg7V+ibJR5frTQpzBIfUR8yvJwlSqyio63C9EdLP+ge8CSU+8LNhqOy5
vbCO9pPz8eBsUk9PwZYtoAPWoVMjY3/bwc1KWvq3jbfVQpBTZ3ByBsnaD6TOIVIECta3lX2oZAcg
vbFrjOXqRH83UEb4DeK9MHQ4iSdvaYCb29E7UDR9/CvGfSQsqyWnyyn5n8JJCAvYKHCxiF5y2lxh
KC/45TEn07Tl1418q3eVXAF9ygKmYw99p+aOc9c/Dmv0gOdh/wAes3ULNqOZmpVzfrclFlaehqS7
kr89YrC7mQjfjkFrY88wEkcgpNcfNStRQHYnc4m4V4BHxSg1tgi0P8L3TKXOgUWqW5W67Al12Icl
3Z7UhcZ1rzZBF2bvtEVHVNRsAGz9UeVRZxagU74gzaXQSMkRHUdqBW3oRd523B77rAVXmB9wlBVI
cJr1SdZu9R00F9mcbMSyKHqzwb67ojKRAojkca7WuJof5Pz3ZlmQH3hMgEgBimJP9vPBSkAZLu5/
VCoNUWfk9lCM3AxU6k1AasxdVKvKLyZ0qaevK1QUrHWytphdXTQIGI4uY88JAqbvDE8yzyyJwtIO
rKmubXAb5R8rsi57cG1N2mJ7sNKBhWzObYjWgNTwRABu5CFLmdseH4+qSETC9911x5WFGU8yqJIp
NcBp9UO38H1iqqyi0EIF8Q+fPK7yZ3xIut/FaGaH7CchMxmxD7Mhpaw30WblW6jKi+Bz0LYHnSNb
Bs4ZIQA43nVMFOOzFsNDy0aU4WN3dmawLweC22DxOpYxcVgiASqOzn9gQ8EezD/Y+Y2mBXr8upws
f534tW5CjAHow5jHwf/ZCZBDisWUHVNDA5AutEmk40CEee4LCSUSnolQfQQffSwpf8wEE91EaSgf
nfZ60mhSglUXmwbV57LkFitwSnkl4U5nuWPteL0t0ihNWUSmnJo2CV9KRrq3WRUMYI5vDBB+Vl5P
J1ISBf8RlxbjBg/0tihP68iJWmLC4NKAbc+SJPZb8oa5TIg7oQKofl3OPG9zh8CrrdnULfSaGfkD
4i1gmTUo7vXwww4EA8Skb0K3qJGUpxOKW3HJBNc/6lTUHeKrdJhpC7jajMkA6l/HhKHtrvgxo6JP
e/r3aHmg94BRt9N7C5gWyHMhjcUP4P4NuJTpA5FsQZG6xZ8fQKBRQI/vorV7Gig7s+mbN4jCYtMz
quaUeBQjSnLYU61YGGuU/vDbTFUMcoaObYAaug7vIi/xCHHZ5WuUPLt5/pQ6eEACsg9umcvIh77e
yA4ZxIEaGqAz9jS6XkEJGox0bEE4LZ4LR5q3SrHu2XSll6L4y1BMffrdAKQAKCaqgWDwQBW1LejP
ilnkm2kGnG4Z2Of+KDnaqoQOqoDusgrWJ7GZEOhxzSH0Q0zyMU15V1NMMfRexZoQ1YCCQCnZYhgz
+i5I3x8Vl1v03aXP8UHb085yNVxUxBwl4iE7wC07dYPlmCZNaSqVFtOtnEjvgQnN0naXzrscFYR6
IrcFzqGl/WsNsoqfZM0R0NjvbqvlsBskWxP/03Af8LCsg6UoQaEYq8tHvKuKmdBQfVMNukJGUs9i
0oOiAm9yNL5YDhMLumipryn3Ua4k/YSOJffToQ28rd7FF1/c8bmUwp4uYKWWxtJhmCQ4QpwBczxY
QHUogk+pkOqhu6All6Xsn4vUWB9UPTVYIgLRlg6Ga5+MYGXVyCXm6GcNnCuF22Hbp7TNzSDD0Gmw
vndQ2et+9YJGPGmTTFl3hA1xN2Zg0m8SfgzIL5JRiJ7fx8+lhQ4nc4vlsWrYIBBRsUGfIePxoFDT
jnIE16PvQVmUi6LIPvBMT+8lecvBmxch1J5jcMqUuNJz16BHP5f7HwKMoltmQG/eWufzlpEVZ/iT
qpbJoBB3FtXCQXjn7acKbPs71pvz7KHrN24lPEA09NDc1ZQC/BmSgFkVbGIfpn4sQditDhtoO5H0
S5TT3jou5OvU8Ew4A0kFK4ErmKonfNdqu5YwoHAs+eRlUWDwAtclNVQlS3MWoaePWK9JGvZVpc4W
SufPuMTSxjf6TBDej7JNNhtntLOQI645aDKZFbmHWvvp3Y2S+HCMEIbq16C8YwS2GmERlSUSH4qj
STms1t8rRZlCtlAGVaUJOsmH+JDSVbWrXef2EIjbJwe8XoyKqvb/fDZSTGBTYLvzIh+AlDsgcRhW
fjWt5t3fZo/1bQ+4pBlmi8jyzg0GK6dxTeo2XwXMhKB6AVLx2BtH/WQcoT+YC8vpLyK8hcTegMHQ
BpsjxkH77TSZqGIUxS/u73EsWwg1xQOFH6XdngQ7H7gRkRYGvbuOXKgWfi9nIE+cUg+gQLlQ1VOw
+m4QaLbmknv2IXdQAxKDdkpVazgjEADtC0G3Rd0UTbEg7Zvg3jVoZR1clhr2uvS72pNZ6braKekG
DmLFcVhwfzMhgDrYL/ibcf3WJ+tNn0YPBHlWXhJbw6LRvu0fKjCyjWVVfhNatdFrqn9zLRrU1e/o
7WgytzfdPyDaQL4lW0ZvuiC1kFjz6Y5o6+c9Z1lY49s+C+PMOmKpV2Uc64NlCV8lxHoN2r0LmTuS
KhQVROUjIvKR8xSBiVom0pC8o+iC2867Nhs8thrQe9vYmIy85lsMzdBtZdHvbrQGWpdFQ+NiKHTs
2VdcLDCsItF4bblGvXXMztm29QS7ZiXC85dV94m4KBs8r7Lms/guu/iUFk3W203ksLpm/qYHGzBm
BiSqh+VAsEDjq+NgkbEd/lcrWQ+5Od+YsmGRUbpAcB0Gdosh4wY55aZRZbjjBjT6LLJVZOEIRhTQ
l3RWXxO979S+oVj3y67skVz8fkRuEdSgyFUy4toaLXZZZNJAYm0X72cZT8HmbZp1H/wZwmg9lPJq
UoiZRdqaL1LRhk3B8LFIFLyXxEq236kFlDT57BGO+AQ9ur8BOSdy3EcktsWrADKve4/eNHD1KSrp
Yx+OxGBEAOhCAweyGCaKXIl0RGju9fEx7arJFeViTgOxwiKBthZse+RKTRgASvzo6WFSf2UZMlYw
yWRL8fz4fkEKaAa4XuH3+B0+4yxvgA4Hr354nc91QxJonkPOgyK2jyY31iQf1gUEsOSAywnddhou
J+ZFIe88pO4/bpkyL3pYAh4O+PQ5mlfb28oMMQ7tnpDN5sNXXdXiFHwIdDBgcROcNoS0NbwZ0j5J
lASXdpvasDbSI12QiBOVKMU/DdB4Ddg0ez9aMP3Olc1aL+H+iFGafo/t9x6Y6kRKt5TTChbT6Pih
1qDAozX94hL39DJ5lO4+p2dxlxpXDOz2foP65w6V7SmUSMMgWUmloFsavjZYJATW41WmJt8O65rl
PXAzFKsYvJe9EhkCaFKZRVCwRazp28n48d5No8dBszYXIpXLkae/UE5rpV6jJsQTWQbwVIRPHySv
gRyoCmx9HckGWDnoydmFo4imkWeJ2WWhqRQyY7/X29/FZmEdqG7N2I6myO8i5cioQvdN2X2FasEg
NGnSe++VC01MUZWyU0g9k+hKlOihHzKdhJd5/j+uOSlhrVx5U7thiIuPtudQFtAvW4yD0OmfFF3W
5CeHxYj0YogaaCd7hlhW79pP0kab0lI81NohNucj2H6wYMpbH6icKkeWXXDQ3y2KFk0chVxP4nv3
sKAGIElT3gYQfr4GU30EmMTRvYgOPM/UQLBI9H0yp79c1s8OvnJWnWWWyAgX8BrI12006BTIk52y
1uTLUcMboYQwENY2FmPZ7nBcNKnjPBCGXc+umwCy7/G3BjKhPJ7+5/c8JDBtgg8b2lZZHABle7it
NkRl6qAjkHtfHrFQ/dRPIhLc/7icDwlkdngv5SsQSkVPURTR48YBfFR0tZJDF93A3wcIBR78wr7/
XzHYotzSACNxordj1Owg3D7UvHGQWDn7DL00j4Cnrv5gum8URvOhpaY+wTAtwl4PLwdyn2cik1dB
ZVTGBFu3Wemrh4UKVBD+VX1GzeYAFi4F1T16qkR8Pw38hsQkC4pPBGZHRwVqICzbNtO7UFRWLs/H
n1wke2nY7nOIsluD+f1hFF3nBiJY2ThhCDCyjhREjkuau52hhF8FyGezPrmR1eRINNB+r2o0YE0C
zmadqpK8syuQSi0jilLueMjG4rW5kKGLE3nbgISSWHQpsFfo8U0mn3fe06payHKaQabokyq0hHxj
fDT+RPirhMhGeeuVB3wxDAWLI2+bLk8/jkPour3kBmYRTW41/TXaJXJcyDoU7y65IVY3HFI4Sbdv
q8TyRuwRddxyQUW4yAGARxDO0TyOxyff0/J232oQbzUvjPaefn1DkbkOduV+kKSSjeixjDeKIN1f
BLdnOz2fc6OllKdYAMPNlTzF+V11PML+1HnyjGxLOMeAQryri8Jbf6Hc0pkk2xWYO5o6bSkKkldg
ncJwLX7dINcLvkc8EjhF2hwQ/PWupaYJQqs0HzfMxvM6mmo7NQBcQxObeFydhqDOGWS4k21Mliaj
Vv2iBwom6u7Xs4ZUH8GoOv6byQb9keM4PGI9tvQ/4ySdnT6EdadWbRPMcOhN/6IW0e/XvAzy2orj
QRop+jwXd8DdPww9N8WOVhMsoYO3OiEnfW++sIX9+KPy4TwStcqoJkjDk7rjREVc8Qx2u27uFt5T
lRIf3qwHjN5LYeeUaUOsiDol+pfvGq1J8JOxFcbA1BZSXwW3shQv/oOXXMOUTjKEuQq6nqAILUOF
l5yDY7fs3xRAy0UZzypgbmbcNz40LSoah4vnSzEyY96ARHQdVYyzY/fCFiIujI4RyyW9b2lKmlvn
WAlXN6Kn8fpDbEj0MU4EzNRSYWbOv5HblNI6VHYKSsMNk42KwbDFOSlcDs54/ERrXcwfyWHYWC6n
qDx6AHbfv2rl43Zl4NJWN3ws00b3OLEQmZ1COz5VutIESNXaLit/pGGHWgBn/NwYRjQ6GQ46RM/G
hIB/iIQXn9McipyBHw5bKKqWHhKEf8579Bzp3I7vRhxkS47XbPGIPCUK6JR+BWU8sHxAmBe7EwIQ
GSF29SzLs+cY6nDSVZlzvhoPQM0iBnzAfWysNPqkX0cxF6LLxqdAiKtc9CeKsWwLoGC0I4xsDD8v
iYI6/MPebAB6JUqaCZAtD1Nal2Qo+INPogh4lSy9e37og9AA0R6fsdaLpgQgQWs8/Y6lv4cj2nFf
AJs7MisKZjWXrkbK/S8m3B0+vE+qXrmben3jcefcs7Y50chyZV5jnJ/XUu7EiQ8mTZ5joNhujIrF
ZPQ7hw37WWv/B2o1jmQPG1bSiI+tASqclT22luohsif0zRS/arIc8pbi2diHeWo7R92aFIoN4IZr
frr5m2GBMQqhenfnbKmvMD/JUmft9j6HlNlJtObLDt2Re9UKDmhFaa7oUnQeVk4x69pzR1+VN426
byZ+LG7WOCuOKPzgRB6OBNUiSgFTSqMsqXG/zV9sdOHHTrC8gde4FS2NFQpJAw2U+jt4ijbnyA9v
WirAo5zJ/lEFl1JGphiRnFagRQML8K7478ogIrJcNj4tdPUi8YP/mfzhiujmDd/j5x4SGLDJ/WUr
xhXU/qZkDmr97jLSmGH54TpcFCmKqfBbIlWkuLTdRA0/BilVqHGEG0/Gl/zfY3wmtF/P6+OYNKeo
2T0QIsIoaHKKgLmCnKIp9tjn3x0hajnujMUj7UvNlyvB6ex/tBDBGmsDdys7iIfqAAy06imf/ffp
tcsj2SOk5ZEOFaXwmJB3RKyzBGOqETe4XAyxKH0lQHyP7yAXXeYlnIl6ic4WsEYmudcx90OYMlPt
OB3pD49aoAKv5sbiHlVJP49d+x14KyKyxTWWMuK9DVZ2T8OHCEngFT2yNqen6r2lIXYmvMNM4sAb
wZ+4kSFL5S9Gj/tm8YHHSEaWU2IByfrtjdNaokDzCpyJvVso/yfRy3fLvAzG2jcWikExmsOItocZ
LygvPhUx0vm7ozYSRWoWRC1QR/Aqc1uXoRAQ4snUigqgFBDT7b63Wp2VTuJpsfqf1yRwYAEhu2YK
2orPkVIa/6M3/p0UJgPIoBxJvGLojgl8D1kU8r4D2KTMHQp2N91NvdvqTdBYmWnhGNxnTzAulY6Z
QZ03usVHEnCvsbAUFvj6MMug0K/L2V2g0HaWVQyeO9YyINltYgs4k2pNLpMs3Rg1LdiLHqJa74JT
yjnyIJ96nFdJt4CpxgixvLygM8FhgKyeDIzL6KxVoeqfLOutVpDju6N8+UfSweDmgE/ycbZQs3PE
PevIAtM3+QB780pbjWr/Cju7L1Vz2G5qAIjzQsU0l9PO5xwZw5QCWoSR6tGsa9TtRXxS0u2DFniw
nSN+ih2jrygSN+DcYhXBbEbnfc+pMhLR+75hF2bnEoFjdPSLc7RjeMlp2I1J4LHBfDiiIVISszte
APcNW+8TNyWkvpx408vmpblz6tdYidJ1xbgzeFJSbmICuXPHOoSD6y5lLfK8VyGdR+AeeqPXM2YF
0YLM/JJ/R48GO9j9x+x4dQTV7ZMSr+IsvvsOPqZ/92DpeNGum4mA9neXaebanStFNoLr3EiZJ3GG
Mot5JxpSPdLhl3eD69+tu5yvzSHWi6ofmFS3beHEOeA/iHHNCt3O2q7tDEnLsxq+AtIwzzxvnfLi
Rj1v4Eyk7faWQJyzRI3AsQFnvNDuR3g+Sp/NPzVgiKC48PgL4ZISLl49v7dqMULQMwk6FHj80UkC
zDC/M0vSp6lB6tVIUMfUgcMiCV4DQYX2fogMothdMbQLnJh+ugJ2xhg5co6dAuHm+nmEF+rzsMqx
UAJXMiWgNmkUUY4SewYnUfinneNEeJM2bW2NbPQwOo7FdOv6Ga5i1uK+mSYqnKLB9h95oUm5ImK+
dFd/iO3jel7jaVTO9GoiS2u3zYovp6Vj3tqzSaJ7H09Tv/33aXlggKhjwOZK7+dZIJRHNlQ9VEzk
dqY2afDqXdpiDHK3aqiA0igbBGtLCQH9caoR2MZ2B7jsaKe1fE3BMMRIj6jorhxgm3MZ8xoen1UR
Bsb8EWYuDqRYWRP8CXqH1TAVaQ4sv24hKIrntPHsyylCVJMKOyKx7bo/MAT0mUIstxEOE8uS/pIO
MARNrX0N6oRvVBKBBjBOHsMs1glINm28peizNWtbLwfjMgE0ZIAt1nicYtUzh0yHprDmd8iue/4C
cEDT1k6YkQ9qowEzVGIwzS1vUUlFmFf3MRSIAploIIGc07jwMse/F+AvB0Ogc7uLd1vy1JINSQ1Z
f566fEWQb8cIfC0boY9+mZEGvz51c0jrS4H2a4gtw2VCQf8yNM5hhPUELEWV53LMgHcgnY3c4Wxf
FBRteIkxDDU1nzpEJevmfKqUej1Q/6Vket+wEXnL7EewXkfDFtUVtLr4PgYfwsw3fPX19hE09Xt3
qwgrbT0HPxCXyCnP57tE7Wer1mn1yhpHPXDCdD3r9ENb+tlQEvtOPbr6flspuc24UnZLX4uCykJG
W4v+l8VN4xbSMyj0GmbQplyugQiT8bS/WLLYAjW6iYZhurRoRBLvq+2qHO5kyPCisoL3R48ia7MZ
9RMgD9qepM5lIqSNdvB3sxw2ItnupqZhj+IZ+aukDZOsMpB4A35I6QA07QiBC5/zdKsxCIiDwASg
bevLHWgUdLECyhCeseFtdiBZxUU3V0bvDbcGnEOlkKwPiwQPuQK2lJN83zBFLdb49bNT/orKHuft
+OYJzVfae2TT/PAITZidr3wDnBKCY3vXZg9HF6Rp+lpDDMVVm3xTchuI/mv0wuxoBmJVKE74Q+CZ
iFOzkPsG83gZ7jIUEOvoXSm1SlTaeObqt+iESUvBRzFYoLi3HF4FS4TCbJjesmkX79wALPjxdN5m
tUUt2qpUKcUXeneFYOpd0SPyOqsp7bTMTbiQwjoOCQK4fyytk7wLA0JsZtIPIKGsiS75uCGtb9Zp
22ntY2JTaUsvRUB/yZUpryo+3MU9FABme/WTcXOIEpReJuHIJH+TTDcHky4fknEKwZ/e+22ZrVRj
wOsKebEftJNjPloXa5nHjlUTYXyXFWJ3+onMoEuD57GdKdUEesDtpOkc+DU41wUbPnFMrBvaecCP
iB+ymQN0P/u7APwwihT0Oy/apPApJfjdGXUiWH4fUb5IhI6IWeDbHwhfYKnF+p+tkYGseJ7YJM4Q
PDFYRpG++QFPYp7fjh9F9Bb+Ecb2M+RucSCtDKRtIBAyDSLTkMF9d+N7akO/T4skOPepPPf/ZaL9
+JCD0Heh2VkZ//pCsDnoonofGpELN6TiglJg2qeFWOjbWfnJA9869+G4bUEgKARN/QcOxX+GqGU7
64cdxaN7kpqPGlwCEwa1yJHWaBZ3rQgvl6iKQF3FsAfH877//dJgdV+84zMzCY/ftkZQr4dZBxlx
/Ambdlho1aENbN2IbPFgBrjC+2gbR/HSPiT+uCn4WfCrKYU08g9/9xvZwgMvRNdiaMfkpQ91npLD
SlAFkHN+yWAeVZ04o3DADzxHdWzCUdgwywubmxkFkFXxM1DCnmdlnnDMKacHPbu7KzEyAne+T7Q2
+Ga7AUgWNJqqFWfnZpc8uwRhZZpOKO5zSRUNEaQrooXaGkaDZGfQumBB2wPh0RP70C0xrNES2VtZ
3qMYcp3W8Lkhaon3h4JMslYzFpB5KZfVloRd1URmLUZ6DpC9YZSNBoy7O+VJ2m8bcyJ7DO18Wqs0
yZTnpWAUSOGZgO43KreIuwWddGaHiSNP41mhbQ7GGej+NSKhkK6wt2i8SVPBjf7vZElUY/QvnA2P
QgBiKHyhqxCdkbDbetaiCjCY7smmBbbxUGijD5TUeF/MoP9breOWsIVY3jt1lDj8QLjAbrjUF6jg
Py1/tzqrwBpg+7m5l32+trtS0pf4ugMASW1WE9irrCaAx1AecMDG+3yHPoJH4HA+wVbzEVQMBpFf
lUUsWbQqiNGYZiQQrmEhWWrBeopdmkQsD8BO/K2R7cH9XT7IbOHjTyhejwWhpOYqcrckn3BFd10/
xp4GPrBUaT2rPD4/2wHcLPUAOpKPV4gp8rx4IlVWxPFxVedVzOejAUzQ9UTYvSRbDk+iNZjTovHz
QoNWcR/r7cjUnbOGRUUclLYlrVFZ9uRwl7t5L04pU0WXO+AMz/H5fo7jTyFml3RoR/F3X0jUPB0D
I/etKWt6h4sslbwAcbJgZP82AlwQ0Sb3ScN6qw/SKg11jeXlcj+z//FL/OWofRGegXaeFRzBElTz
ee2VGv60PRmAzerVUeqeIXaKHtD8ThpvJJjqNDHMucZ9iOo14C9dZ4eGw3fSTVcH0vZMgwjEZOQx
hGrHrTKR5Hra06ABX+unCEuecHk2Tcg0uynJwhQUbyiLNYDVW4TCdzeJOcO/es0VLH59A15mp8GH
0Ea//UmWQu/PsGuXzWXWLJYwQyBjZIly0hVrwRz8duXdwGCQgrMYdRWkQPTsEua9OSO11whr9c3Q
UmKI/tjyRNFRz7YB7iPgnFHIUGAwN926Cdl5AvY8af4XlnmLeU5Juq/ZrPy28xJS2UJfM1iq9Ewh
k3Z4g/tuDsJ6VFMbnDYdpSewMFkeXKjD4haZRk4w2gZ1qJBYkInqNoFW4xPn6pS1rq7NeIBzM0zT
zHA/E/IHiG4CbV49KtwqVjYUkIMgjtKiZSVL56dbuYNwTp5PSqtYNZgVJqzyjKdSzPfPMecb66FG
jJ/ZeMY8HlPl4d3ImsziQ4Y5H+6J+EUCt6AjCvyZs4ilE3NRA5gn5L7S79WaxoWJoaTlmTTZZowd
bgRlDauEPJ3USPIj+TZ98ztNTTOyu8oDqv5dzWUMZemeKHz15NZIvjLOhFZPkBeQdUu3lPvCiI1m
AXpElm1qlz8b5t/T8L8ZPTAPp+1RAirUTECouwjhngPJahGianYo0nX+ell2+YZvhVLsVKJtQLJC
Dt6COj7+S/egfJ8ba4q6HSDs+h0ot3mVADdr8tXBHNWjVOjtPreP8fIvjpTlV5GM3dAIVXzwTmSX
2EvTBLxvrrjthFKPOo8Kv0+CzrQPv2AMYTnpZPQ1tCYOkO7Q4lL9m7qH02VA1NXaGRenYP4H7eAY
h8ilzT2jyeg/Bbz1D04YuARWLELN3yJtT6MS0nbBcmX4W6jmnla8xzHM/jEM5aFOXSkW8orGhqWw
rWI9HIrB6YHnRua8Emzyr/n3PqOXeRYGfjgfqjC0ea/FDUB+w5FbCI1+GqVxI/TSuqZ3BG9V+OtL
RREBKTWwF+W+UHFabu30q4JFrBRO0g8SraJPknjV42gaaG4LD4803GSG9BFu/E8xFq/JGq0Hm4HD
o2ypLaraV1csZg/LRdQt+M1EpnabjhcMj2IaK2IbM3j6cKgmjV5ESaVptPcXbz0yxWWtEWSV/7jz
sEV0RLFJpB/iP+2QOt0wYGhKxt8iTBVQxK08wnwKY4htDIXPccsYgORnzoEIlMDa08Nhl+5FbiHm
A+1L6ucn7C/qV3ABbGkZCWIaq9NVLqfpl9d3tqf5AcB8pKa/c9xYzV0LKppvmoyJ4fylIMZcDdXM
KKeIvwXQZRvWzOSFYDyVS05/zzZJwC/z/rT0LtlalQcIo2DBiauQKPdJ8stGXd+rsy0xqEspGDuH
vJtWsdsblTzTjXb/6OMIirhBEVDYtRFxSidGGW78ds/K+Ncd6lb8hPjIEmIvDUCuXBtZt1ZM3P0d
EZLAh2A+fL3n4MJY99+0snLfI3BQjM9owsqJJidnW2Iu65m0B3j4wjqTtA87XggJ/ABbVMVEQbk7
9+blbuvRRYVkVVMgYjAmrA6HYQpM6wV/wc+RI9xesCF5A3UGGYT7av+pvEKNAuvFuAMXZYiFkI8Y
3GEHaOeSjc9a4xGD95V8L17NkP04gPYMX7S5T4Rin3PFZQ8ddn/Fk3oL5QqLwtGslHdV7kqASzj7
NXpN5g90o22ao6H7IuA7b532W6JYdJnXWT09H+3A18vEmEZM7UMjBYCSgoPgF01zuSomJM+dk7wF
SOAA4Mzi6o3v0IycitR+1yE/Zm0BND8cBmwq7LwmKcwNlUnkc/0ZC8fuusivZG2AP2xVKvZn3qg4
EeL7zKQrJyhlR24oHGg2nz6VTGmHOxpuMu4AQmXvQjlQ8e3m0jBt4swU8WQAc45cg+Djm3/W9pk0
BrfR8WNS849voSQ7nwl+oI2kYNXZE6Yzo8HKyGD7wdbCBWlfdjg+K2y76z+q104x6HoNZ6zCB5Hz
CQJzrhGfDt5NawE0zg+3+8aj30ULPMD72KfMNL5M76msVjuYk205zRvYQ1Z+/QDIyoKdoua5lL7m
WhD364vMPYFeL17lg+UNWn87DUUhdCTR7rqOX3HAIydYpCy/0gd3K+pYtZeECv7KcidoOAVwAlrv
+bRwjV7TZIiJXqpqd0Nevn/angFqka9DaXF+3nJMJFHT7mnU+uHELtq8zjlmar3e+VDdVes21iXz
tECvJlFQrpBnqeZrfAwnKyr6F+S3YQIsPhWLr4Y11uII0CsxYGCZI3LTSAALm9KEagDM5+axbMM/
kb2yVfmOdSTgNoiCfW+BWfd3Dr5GniA3o8xjMBrq8BGbF0gDCnOXj0FpZlDUgEESCTaDD7brvFBd
XOv4Hak0XTpq4QNqnDvFU1krCzmWK4SJj6Sk/6/DhGOH1Jk8ESKu8XBCtPRBrK50NTiZd/YmlyAo
9ulHjTUICkMt33um9qIKVB61JplAn2QauUoAU0hxLTL89pI1inYc/rCSydPmAtUm22wYZpcMztJM
L4VXxyfm0WvKOqixiu4zsijAMP8Jd8645Q8NcFDvamUoD1fJF3EYQv+WNC9NNcVC+lmazQ4zSzun
JkilsNs2biEgYDaMerMZAujnlGT8MPnQABo/XllCnEUaiNEwLDD1tbJDGCavqmFX1d1j0F0FSBWK
4zLTZdzJ9hNbWCVYoMPJvYEj8LVu07ED35VvIXYdgDD5n+cgpkv3055txDwRHPV688oTyLxxFw7r
s3rH/pc+8hn3Z2G2K3zbz9pm1qXfFyNor0BwOHkflwmNwLYGpAQ3kzNrbIN0zQfSeKmA4ciX8JtV
bwT8VHJaHyGpFtd/HHPY5UuTUZTQ4/beS4QYl3vgdGEJDukAKDIr1YpiLyKVUfrmpy0Z88P3gQjg
g28CiqVpumWRIsFVhARDK0qgoOiI021f4KBApQAgkWjwVoc2hqtzlK3H9ocD3BCOW14IaLZYRniC
p2h72aCYDHFLDZM2XV0xFGXSFcJd4cS7wFUhyQ+5LxqGH/VRsGKcMHr67lkwRRSrbXUij/5Hv5kt
9WPFPMimHBkgF/EW8KatzOK8NHddhtMB8UNOeUFwxdfjc3/UzhXedrPct4e9MxkgfaeVWvgBehZ+
vSO2bCX+K8BN2HD+xpfDTlkAIb91/80kXsZSKSn4ehGLH+DCoMTvePYur+MFOweCsghTaSsDfZMN
rdPi7zR8yHhlLw9dMpuqADiH1uqqyKtkc6KLJEe94YD0MAK+cAPZQgqe9apPp0P6d7X5mIDsHq5g
zKInlTxeLIfeyupC2E6Vi4rmexuw4DTjiEFtf6b36zdQpdFChDI2Ut8Lm3MAlBjN7BYJZF2H6O3k
fingebEBqRo1LEN5MXwP2hJAvzbY3M5HBcC20X9DeF+bt5NT3qfwYPTH6Itmg4oy58WByfpkqs8N
QhljqWAB5cbVl5eQM+5rDh5eVww0e05TD3sCZr//LpZ2BMvqrVB45uwT27feVNyomiBZP1oh9tc5
ti9DnntcvuFxc/K+7RcukNyywRTTGhMReNXCCcdwwAV9NcpTP7zWlEZUf0c/yUlPK2kobfOC+R2S
cOVZUKUCHk7BkTqNmNsVrX7wKcDzHaNoQLMI74wjjbHDipzw6KKsMe/onJKRNrcXc65MICGcbwVm
Xg3mK8gZ8x4zH5yJfR/ncUdy9V0Qh9ljHQlKCIIBeJWrTuT+gImwxuXudpHP7qr+sKqbsK+GNd9H
UiGRP1V6XNXZo6AxHqlany1Oj8uine42brOlhdHXkm4wL1+GMj6dv6KrhUMuoN/JKj4cmxCP4Ne/
MM8TBVj+ipLwyxREqhIGTLYDzqFYv7jKmITDxaHCBBe9f5WPTJqvTmfydjDdYaY9gU0FeT/okwBx
p8XexbRdOnHU5aoYt7+DirB/NpBu2l/CDIIWW0Ga8tpEYPJ//cyINjgYeH7iavzoavTlgY+gvsC5
BNDJwyNMeYcxR+mPR8rgdV9qd1Qi0JvZDqR0eWMyfxU+mekHQIneB7BVFQNrFZXI4HjE4qhDNWzg
9HORwpDiCKgSBM/eWX36cMVLQYbZgozGIslT8SYA4gjxcwkkwP2Oh7h3wpykJueK/Qb3fQkIQ/do
iDrWA+hkLDi5myNSknSiHgROg8A8liA8WXYKMeT04WkPvxnmXPh+TlHd+/JDKVJ/HnSf0l4+zQFO
ZqStSw/q1jUmfYi7U1+PKHAeZ4RszS9PaziSS0umq0YAkuEVs1QKHM6TTd0P6BGh31qpL2cw9GCr
PtZS/xbKLWR4Eb4zPJuE0yM78WiOI384p72fSEpXCxJdi7ea+MhG8cQg6574T2vQfohJ8XqAarXK
Sf9tcD4R8WN459Ti7bAdL8lcxH/16YGE6ZDJaC5xRzbvMtkuHEC+nBdnpeKRHWcYI4IGzjlU6v1o
e3YbV9Yrv7N98+5cakWNMoYLgqXhHspxH0o5AjwIAwycULxu8rVb+ddTdikVcP5+U1LyjG4xmitj
J7nHeZymGBiC+RZEtJvRziWMkXPhGHcPmbHFvOL/8T+9HYpGdEmEivywdsCHKFpis7oq6FmdthXH
cIYZApVWxi/f1lmUkJuD1oZ489DnLPYyZfvqye8XwG+wuPFitg4ifDC+5/qWHv0irApgHW+G7IM1
977CMnEckXiWbjegxCdDz8oupMy8+8XzI16+zvLAEHISwacRVwie2tt8fzO2lgKtVALzTZb2o8a3
O8yFXrZjnTtSJYum0/nQ1wM3EHzokzBcnLDpMuUVRJKMusNblvUaBHbv9ZyBserh2+tzSVH91v/o
+VwoSDqtDPXm5tvKqxdh/6m2oGybW+VK9FGiZr7uxI/PM2Dl5y++/p17nOpr7R3I4PcYKZGzb4eA
FpMXnHaY+glL3eZpr75QOUsP6wTDjTWu+SbtLbyqeCBO7EC9NQnqc54JKxzo2uQ/4cK4TYdedPDE
Rur6pxtkI4c3lOApJ+GBVJPQz9HGAlCxyKo0fENvxAChrTVxo1PxjcTkirTGZAmtm8yhc9E7PB65
BwkZ7aoj71S2REjTie4SXSuFJ1HbW/PS49K3GHFXDfYStVLdjPSDbhUIEf6elDJAuodXJFxmqwlI
TvETI2VQ5yi8tnM1uX+h+D1sn/jHdQZCYdp5kwKuz7L4jcuPL8M9Ml/y28HOe/tlzBGW+XdKJNtu
uLx4S5WBxh1oYsGzc2u2qt7bwj8VO7nW1iUusRUG5ECXFoCWxRFN4fggXXMKbx2qf+9j1a0MPS/C
HFpf6cemuzFQvNmtyUV9dmKEpWXJ6e5i/TTkiJSdY/zeujMGsQDbpusVexnn6UYMSCv4XGGw09A2
mCDFJSxShWQ5958Z1qI2DdsWDbl86TlwVfpp+hhPwpnIpS4cnn3zPsTMV08rdjuY6Lare4FVtB6D
GALwEuhu6GLf2sWhIZEu1ubK1v3VEys+1ZkbCMqxyiIKl1EY7xqts38osWCgInJxTPQfIM9QMZR/
7X0JWF0yyE+0JDdrv2aagTxwbp1gpOpR8YpBqOne7lTvsIUxLqoVfeEeWvbQNXxaPmzW9zkhwp/p
+9Ut27OBO0N3o4dnV+1FFKq9jls3Lqo6agYUhxPK6WFE740fQKqAh7/fW8uQlY9zadzJSXGZVgJA
4AfmoXvx/rXv82vxZQiMLecDkqrCSPBxo9QD6c31RiVihjsP7md4ZDdgTLID1RdmZiv+ph/ulY5o
vGVEyK7OYgZdIuHmR/Y6/DBZtwskMhaaGk+aHwEnkHNK5Z071Tsefu/13k9q3RchWe97lW5nhZGF
y3wzRgJNB+gwp3+qAmpDKZqAhHIUoYCGEhWPEhidoxDhgdRclnIGqEZPkWCGC4doNDyL5FFHtU3+
yYoekAXRcyC1TJAbUawQvbjY/HXEON0ZbvePi2BxOn18xaWR6614SSDOMDuq4sKQge5cHlaRfQ1B
/lSoJqUbyhS1Zu8mC4AShexLzk2xj940sXhEWBZ9JfmjiNtGzA0aVgoVlS6CeT1iheTDJpCx7xQu
zN8PhrBCdoL/mIARY8yvjQTjGrLYLt4ZN0Ru0RzDUQKcjRU24dPz3jv0w8PsKTpMgpgAaVDimTwg
pQj5AXqzVrP5QOp/dJWxVd8Mc0u29SXmN4qsH6WqXHeVS+VgTQKgPaB6m0PAu/YxRRL3oie6OKYC
r0ui3M7u0PaG6w0ROtFNySHzR3flU+O5bmgFgOM/W4aUuXggK7s9ctS895CAfotke6C4KaZVB+F2
cioGMMje7mzIXfJfL+5l5ZUvEergrex06Hm8Yau2hNCf5qeJ205q5p1EJ66vnAIXDaUR6QdNdH6Q
sagsT//gqKhYO0ITNmP5Z1lOOYCeCNK+tgeHxT76FzmcjMYnZfG7wZc12OTQVA8IhHNc00Kh7Rut
Yhx633PFTeVjyQrX+ej5rNUP1g3JgKR6mbjXvfxgb7fRLudc0SHEiMbbrXWn2ypuSzg1ARROoPct
SKxO5yZEKwDW5Khl2E91VIIECA6WDpfB8ASBnCyfHl7r4soB32BBY2aeXXRy5V8sn920HPyVrOKi
EL4pb4BX+vCHYu2McjUaQpqhaJyWQEhhaPdX/ZDwm7RGhXYs2a0tq26JFTMCF5Zkb2IcwRfRofdi
CmnH41CaMl01h3nq4Wf7A4aCTSIu7KeJ0o9rylw0Q7ePQw+tuwfDAK26NfjWUdhXBRDteZRQYfFd
IDrdHQlWp+bADaa+KKrWHON2AUMBDljHAaOIGEyJ5RkuhzHxvhmMn0HFQ1GVkF4BFZtCYuGEHxwl
BKuZH+dEGwHYgHzaHf3Q8WjzM5FlfCTwti+PvIkKe1HAstnO38+wUJ3uFXZ4KBegOeoOqnd74sX7
legRIi7KoQg0OYFFk/0UCv1G3YtzTk0QCUqARDkgP/x6KQmyM+qdjtj0hb7cFgJb84Ct7iYQ5ljB
qe3//O7b8x8SgXjUHHZCTGAyvKbNAZbYD9yID92aN9iGTm3h+by7Blnj6f63mI8rgkikEdl9ctMt
2pvZIoa+Z99nQBKNBXhwph8G6sg0moEfVHsvNKODAcmhmJLocY1z0vODWxSbWmPRTuKGdfSUxdgk
E5UYZ/XZlkFBZsV5z9LIc0mXE8j3hDjqpRk7vbjLsuv5TGrlfF/qkGZueWd/5+pbmxHkxSMY19Jx
6JA0Sase9vChJT8FXfarrV/Dc+V13qSXTabu00JV9njrqNpKcF+SXYl4ZhTWiNoC/HGGYtds12+p
swqIHHwQbThYLJNAWkmgN2rVh+yWl6X5oO/jDazxoRYq3f2N6cCojqDVAZlD1uitV30KTAB2bmjI
cfJprNgHsrxCX76JBIgfr4uEyfa5closCs+oCayVY5WjuGcdmR/SDMLpGofV1EXdNHJGWWvThcmw
i53lcFuFVHRBQH+5/LrIMcXfT09pPWtGT7czIF00CIUq4zlEXy8LGodjJKp7c/uvtLI66TQ1V5AJ
yei1YiP/UtWIpC7demMsHEKtP3q4TO/8BHOUQ46kkO5nQ54fIkBNE0r+FhNNUAUaQFjWaso9ocMc
ljTrTXTD5UllD+LDhP0oTvmsFZTqCewCao598OmckX5pjlv9ZG1AGE+FJm3NEFuIPpCl/Riq7TxR
KaiX9cncRt8c52v0SdpFDfv+dkIOZy8k77ln9SsHc4gKTnbMUuAft5o92cBlysqE+KGDCp5rJANi
AoM2+P9Xm97IJLbXot35TQ4k0CxJM6RWpieki3CYHeYJcHbj7+QJH854hPj94tQ6dNReu7G48qwI
s37lOY85+qfIR5MG7IsCeCK4V6cY4QeHnIo3VL1oiuRQOHc9NeeOoiFpDe0gdx7KpxMQ4bxSugUe
tw1+YgyiloDxExUX9itiL2blkViaxo0QcGuSqt9cCATL8rHuZ1QR/Tbs8A8oLM0iBRFEST7vY16/
LJLPuPInITZu0y/JbslNm/wYbwm1PgH172DCJGzxeZYu+nNev+M8jN6h9ISXC+o+xfPURJ5/crHO
xraizE6eqJe0yd8NSQyRscG1nd6anLmPL0oRuT8+7vEj2GRnYvqTV26jk1+e3zE/vF4P0sqvsn1o
nD+j8A/7tc1KyAGrLC09tMW6ja0oF3QGCg2VVhEhfLZ+4wx9q7Ud3Oup2xJF1hJ7FPF5chTRHC9f
I/w20lg1mB84CPAiyDrc2BqaoBXClS2gfKelIDuScvUKyTu0qbIoaD5g2+203+jSEH0v2JMl139S
77e8y3WazFLRxGLKlXlq8otsSZD/M/uYv0VehLldQzG0qSb2t9rL+MPJeK+JCVk6rEZ4M//ifN5S
7oziu6Hf5kFnT1wtonVWcVN4yay1Zq/tfq/u/l7DgqgyfFni4qRrt6Jvl5/Srvy/xTc+r4dR5YQV
tIa18Yql9CzdsD3Lm94CM1DesWke6rkS06Hljkhb2AWPOY8V9VnxTmUVNBeZrhx5s2scW8lnQTAN
Bd7P6VJK5DnO2TQ/60Pqws/A7t90NPIXCGBLv1Q6XKlKV4ZpbiK1eWj8gTAjjueIJRPV5ndAdeL+
A/+CFdvtPvo8JkKgjzJNXT2Pyadx115MNsLyT7Jtksl7A4XZwa1iUTS1JEf4rYs3r+yRzvSXqWIn
pAcN2uLluE9PSryrfxoMGZZQNZEXZg3Ue1Q8rDI0q8KguandJGdfIibeYtM3yH3yAVEsoIB2JV/W
3+KOF0OGr96wkvgU9eRm2jBPXg9alphvKKO3kUxdE89DsBG6GZfJ76BXjZeNuOseJn5D9yedGkHJ
uepLfn8JV+arMg0FeNtvTDZIeHtji6mwQqrHKs1A50vteU0MY6H7sPsVTro67/ruQYVPYwxOx7LP
DGQjug17r31yIf/U6McCynThK5LjCRHScomKwvpQpIw3frNCMR5kVCgu5JU0z4NM/ndblX7bvhJ3
SDte+gOh2DbwTyCYtDmCQGXsfiYwqaIxuaM0PQ3O0Z22iyFFj+8Pe8fjU+58y7NEd89O/9Dry5gv
luZZE/gV5KAlMCMV7f5dizDRTmIT1Iaf4QM0NEgip5eeR1vkrSKkJNFlPevf3ggzuvoii6xV2Cxi
5fFHABpVIEaRfLC1zFvYgLKdPlA2e3N/UL3TnXREw4yPNhjETKM2EB//dEK/uGLSpZkcG5guzpv1
lkvDFuW/UJeoR6KQjktZvLj+gsGIArCbV6//BYhm19R1FYGHArJG3bR24XEOTqXJUIWXrX8uIx+H
4uoN18wXPAU2SyR1wNFHPttGRaXLHPGJntftbBcVbqO5vmtFE1xSUDG1WZ4+uyhOhv8WmwFn5WVA
HD7OaKjnjqCP9hGlYGMB26vj4lDsDgJREVxRCwio//UOCYkmvH4xUPpMo08LUu+d9BYzte6oKd5Q
ckB0dj6SZW+QV/G/TQOt50ADvEOQ1TkjuHM8WTqxF4pX6GTltM7hlfD6eE/WyMYN8JnzyPD+fa20
iVQcM6GKhntzsozECXbmKwVR1GzpTO15wtLndOhy9QuU1t+Rq4P2SI7UW115yUUFKu+ntzH5Ob1+
NYZgRYPYs3g5KX9anU9NZ4XnoSRmXOvgjWQ5KL07F5009Vmlr7E0U6nzoRPlL/ZGLmSCZG7F5tzS
SxfFT7OKRUJ29BR1RJcu/1KmR6ELhbNdW3LS2dOFiRftUeSNrTRAet/et6uZ7BWMjRQF/iTYg5IF
aGLLVlq+zYOE+wFUx/8h5PCVvMDtTSHWVCeYkWs6x0TsmJQoBxVFMV/ozXuPXap2SeT7MQLCmxRH
9FVJgU7KWLEk78lGQGm6FwTmNLQpBgnTyYKoKMwRLppYLniyQ8rWHlBGZ4BGnuwdb1aEXFWPOOeQ
Bj9/JcLjbATGhmpxx3MDrdvZpCN5TJ4EiL8ACKth1B87L+LFkRvmhRe5LpJa41R6nedP74CQB3rg
+6almuHwhlUddjQFilqviFlGyOBChlBpg/+Auy0Jxi7cGgf020SfLrg1acpx2nN3/PA4wsvM95An
fFmZQQn1hadGknkV2wXxGbZ0VHaswXmL1ou78Py4FkXWCBTgoIJnWlbHg/UsQ/pWTIvM7+NPh3zT
AIWTunoR64+walMA/HgTeDyYaR+ait1rylVgZfoYp91oUA6iCZ3yIqMbwNLJ0iPzIAcA1IudkjnQ
XJgvE5VeJSYagINbGVAEOKGEuYu3BhGK1fnP0UoKikM0yXse8e0Q23JiRqb4k3VwFAPm5BUAEAL/
WmbVxp+U6vSHxMkBNFZMhbCvKRB8p0kKLiYIapy/m/K01GvYuIoutdTitoEYn4wV9a1JFGyUe3ne
hnnXGZBMI5WDLIsTlPwBq3517etAT3rGqUkRR2uNSJcAqS34CuAepR/IEyyI2zWfOXVHyVl0S2ij
b8R68EeUA+74uBMq9khAoWFS3ixfa9qECxkG4T+AxKiYElQ7AMnHNMvpFa2Pq/sqY7ZbJUWgWlho
l3tzNLNw/YtY7+GKBOxd3IBBfqGuNMwFvek6iIEXeckKHVRAkdZLR0Qb0q6kO77wehp37uO+yr34
lgC8CkQS0NiyIq6N30GOhnBhjDv/hRSpXdP6cng2R3uFGihnYLiM6bAYOem/nFjiTaHxj6fhn+NF
Mk1iV0/ucS97Lf1eOSTuaH8ar7B8hTkqcw6Jbn+9eaxJYeR98pF8M2aws9ZA+YZe2tjn5/jguVZW
S5Kt9puoWG8kxVIpQ4FmO8MFqSZmFN6kMH+gq4rYaLNWVeKM5hijfCDOXI4EcR5WypcBQtzo1Ydc
FZyn+m4Re17yieHEhbsmHVEt/XocGH2XvFDxIfqu3MyUM0eBRqR0QM9X5EyogTve4X5Dy9waZo+K
oUEyRW1z1/r9nN//nXP/GRWGuLjupvIM6lAkoq6KmvSQKvx8RKixwo1tnQANEGT60lvk8zyuR46R
Ks0quOmM689jRBDZ7G/n1/waeYn9stuC0G9cmlApeDLTmqNd0DjOpzTTCgtkMpAlIxhfXQn8p+2G
uBs1gIdoyCHeWH+q6GRYrbfQ36dxSSN9/3HNeg2u9yF/gLRh/H0H+HOBldpSlyP83xtqxWzNHfO3
vskk1p/tSOFEfbOZS2oxaE2OEd3qU7eXGoX8oh+N/t8nl1yZ1500F/ZhTLPTx989r6HbNs843u4x
pK8hwmdv8YcK4fDq1splZS4KvzMZS+mY2WLnN7JLx+LhABD7sS36T7ER2HIrFdQ7TkoFH6NCB6oj
rnLcvYNrDI3rbWxy+d2HtPKC0N921ST98xv+uNfaXOevN4Tz1wedFhv0NEFwsNG86hjM72E94Edm
Tj+1tDWgnC5q0mj9qzim2czcOoOQmifGYJmbjalNAs8bRFJ+83RDDf3Y4GC9Ul7+mt6ghyP7i2Se
KvU9MVuzEeM4na7BuHUs2UBOxxCQ1lyBnBZqGEU0jlI0Dnjv4bDHtyP9LG6y6F3hwzh3+MebRxZw
Ax1aEA1kD8PipOp58HB7pl6JowVUPC+WnrZzIvP5Phv5J9m8IAz9beQUZ/VnQ9Z4lhTRzh4yVHr7
f1bXWNEe0Gbiwih72yOwpOyT7+D33MGemr50We20Pai60glv1M2/aDgyqE1aVwjvrN3GSjD92PyG
6RkV2vjPhd7VU6OXVkr/m9DNYeYFKgTm4+rIMJIdES8Qu7JVQuSRodJ8e+VMzAXguHF5guMJ2kFf
YLnylnSdPDYB4mjTuV7a5dMxw2EcnDh1LJuANXzE9uWrwzxmsaV/fAvNYEL8TE7V5wBoKf4+xRPd
wjv4DT54+7VmHGTqNbTdpL60anfP+i1w5WXWqkViwOaZFquVz8ZYs3UwFqvEi2wGoBX8AL1Y7Qf8
X+kiSkJORxegaiiJLmwAtd7D7GT/GHmBfDSXlg/mYjx2NAJS8DgFdjLxfYqaeKnrw683kHAOZQRl
ja8Izt7quhPhg8KkEAF6y8h9Yfb+yyA51aUFM6QTG18lavKBof0CAEO7DmoR+8bOOmk1RXYdeClQ
K9DDmGGZO2M/LDvZN+Y2kLflybLCFiwuRE0s8f1GXqNblI4Ih/I56vuJNsVVnjbd/tZxDSKTlLr2
18P2Xy9H4M6Yedv57+JS+sdqavKEGcTzYzXOrpwi/fCrFcAI9tF0oINcjTEwSSLKotju61VfWGB+
AKv7Egn/OkJ7jd//jW8G7zZpv0Jnje6O6oL6oEj+2RBbYqgxJb363fiu5Jp3T6sRxEoQqCUl5/W0
4kOaFgiT/rGCpKKE0Rhlr5ZIuEZ1I8WywqSHCyHvIQGHE0o+V1cXlCeEoAUCfxf6NlQL7P4FZRRO
WO4/h6oPQJsNSLVKpTQtGURVT0tJBFEPN6afJMQjtAYm20phbpipuanfb80aj3dv/KV/SfIz9twr
5B/bfGsVn1Huq89mXE1Dinvx0HCU1HcYGewVZh7unRfMG2QDIPNojlEewSiet9XsQv4Nup9I+kms
lQtNrFmxuDUM/g3YE5eMZ3//3ShI2h1z7EzeDeykK6iJpEMDW1E0kaD4nYGlCzQOSlCwZ3sl3Dv0
qa+ARqfIKWKRWT9Y9EZ/XLknbBpmTYemW28wqz+DcpSA5cauOt1iXD7kQhvhjOapQbZqOiSGWQdH
W8s2GrE8kjR4ZqFIKUlXvgNeh6KhcjUscNAn8MFOtpV2wo4IoC/1qDE6HAy1F4EPado35zaz1GcV
pfYZLChZ2rQQPMhWAbp0P5kzgE5+CvSXFVZJX0Py2hGToyls0tsVCZUTDMcXSAc6itUpiF4bp2NO
SjNhhCp+/0PcQRKQAk9yo35VnkbHgqzTMpxTGUKdjYl6Mez/FDcF4+eDULq5Y9x4iaj5XhA8PLiJ
8fa1Uk1+Dt9yxCO8D0xi0lf50V63gnjgz+0fU1hBBKE4GEcDYjYU30IzbSb9EcF3Rx2GVHgMME9R
JskSTGx8AUIACbbA/JUzdNXvXGdNAeZdD6Cyn0JnU7FnVAHG5rl4itI+KjFWM1h094eWVrIH9t3+
sf3fdflyDca2trBSVZC9cnWqIqmkmdspKiDF+Pu/JR8za7lZ+moKQ6q48jubqSixwEyKZ6q5odFa
FUVsj3QGq20XTPVBJPjavvPACE86zdgTFVuFAKOVOWsZurEkI5M3epcuuyl8TZk6TJs6x1ofejid
eJlEspxJQJgSq4Z/yU4aYVaA02gg6zpQ7sfAqA/SVERrngUA11raWThdMlVyt393H5hE4WwHYPdS
9EDRYE1ttoDyEwNl1NKgqjxOHc8N3yemDhUlXhznuNaHGIk2+Q0c4znz4Km194B5P0XwL1KiMGli
lUM9UkXf3XDW6FhPn9ZTc52B8jIZttLlXeGa6BetZP1t1VptrgGQreeZJHKfK4haYmFyYBCUYJGK
ZqSxUb4r4eSuum9HhZy1Ycc0jbrC3sO8sBK4KN/4RHfxTWLE48tCczxnrT2wtJK09rVTl3Xkh9L2
ce60CkCliqPL7x1MT/19ejUeGh9UmZzTAPYG5/XaYBukPXu8Ms13PMZnTOzhADOlUzHe1N2SJXQF
Gbnm3xs9UIfFTW4iBK7QjKMrAWO10rAdPI7ayaemc+mkGq48jeo0csw68Nj4u8uzjlD1p8WMYun6
TP3anrqbsaaWMInVJ7XVVbr87Wc6ISgc7NaD3d9MeucOVfcN3CRxHmk77agxscbvPxM5qGxiQ18g
0sncDyr/AlByh74UcghsltNapWphWNpjLeGex4+B6YAYo2IWZneG8ztZwX8KMtpElnlUkS4KpU/V
SibtZ8lVvXYrov9mvvd1ROhCE67wMNIirM3fxCFDxWhgewHyO55BrS05ukPpW78cIVDX0MHxjs/F
/UwgQHlcyHOxU19K+h6mZd70Yd5YgGEVNpxH6wcXNo/Bq7VFL6evlpSAXhoI75WsnNIw0imhWdeT
U1HNDAI8Bv67gIZRO6a1EYOXTqa2r1nseUR0dV978uDewqqxxX80hUxg/OwDWtuOIGzPzO0Y4+O7
9oilZdUkcGoR6gyZQ3RaDKVOIUBRbXA6rpfHx1otz091n8C/4+nPz8/HqoV/UcxDpueLsJSd51Uf
VOZdJFKs/OwmFD9yVH6xOOWrsO6nEF/K5aaSXmk11+U5E+AIyQCdcACZwFeYxbzV4uf+vwyklj4q
ghb//b2byet3BqaTgMF+XkvWj0j3W+JcSE5V8FKEddKD9ZJIaFDYHSPGskPHHbEbQZlMTtRGbgWt
ax+YVNk9juanhujGD/ytd/VpUFHla7VIG6RnkOkxkRp+fLbtA5AygVam57mTs4wP6LI+Uyoqh2bD
ouTVVZKcuBfsiw4NAUHJ1TjPmSwaEeLNvZXI9U17CdMRdCR4fkDPwxO4WPMDqVwiAH0HyjbIzrOH
NnsnYqKgVO38HjfFiRmepXrwj2GVeVXzSADfWY/6eQOTpL6VWBJBtmkSlWKnkw52t7yS15LXS135
oDQITzVGpMxXcAKy0FZ9asJbX0Sg3CYHs2h6loNtUq/48WcwNT+vzBQ4Owj3eInTyxo2I8y6slO7
vFNijJODBaZTJX3Qy5BUVZSeV6y6x9mcFIj7oDdP4g0scrzNZrepSOXueXr8A3TozUkzNfHsHqr1
cEWYCwJ7WL6nY7dzkeMaBuzh2x9EXgBroAzZvHMgc0j3b/z8ANVBDRVP2TIyr23p5yRMrNIbzWNn
I+7WQvU9k03nx42TSBd2PF/eFbkMKbfqYMRpcIDQ5hIlHHmKRkCYnSY6eFLmXT/k4fTjNBHwOlEL
ybBWS+7BBbSHgPG/Gs7v8EAbjmLvdeVXamVLT+TIyW0dsY7HjXlQl1z+Jb+e6LgDblxsH4KnuIPE
1GUkiuns1/qOWphFGfeEED6euN1MiHUF2YfX/6RCmmEGDVHnfYUZbXnY9CynyrLd3s38KkXsFWuK
OAjuE1TvRmNc6G6zDefhXN2OKCqw6DSYDnuumQLn8srRLpei/iYeLZM4uFfcRwlgpf7C0LBl7n9D
ECiDtyJwW35Mv7LycvkFD+9w4hth7DqI/mQt8SSYZaM973PsJUUbgO0Io8MO4ARALQkiejGmYr7x
THOIO/uznqNmpyRVAcGAczWQkzJYpKSPlekajk4HufA9Dtsitgx/IMlghY1Nm5uDs/k3+FxPptDc
hz6FWdkOPD+L0n615SXb5sz2JmaJBcHYTrzOWaWHQQ8AxgD0OX4cZ7LMmBs+6bMLwgDq6Yru4B6y
eUaksz3Uc9gIuRBsS7KtP7+CeoUrknVx4qiPKR63Ssdzt5IrvaRl67o+VB/AP51JBg7sHqEICap9
UZlhdmOwNDJI0uHe7cXJEcB1Ggi+IQn+CS3b1ap3dqdmD+7DSUHI7vorGUlv4D6a3A8o7IHWKQW7
M2xz5zUiFrS1mQDC3GvPrtb6es1dYdSC2nPpAKA2pD6ZsUmvSaPUNTpKdmeKf5cYDhc7TaFRdb5y
fPXs9lWK6218QrvLQm/hRZ5edeWCHA2Vz9YqqXZoQxvObUP74p3TRbAx0AGuOrhuY4iBToN0WMQx
PO4mMUc9l3rmJOC2yEm3/wUgaJGjU7k2F+Y+xUM9cgSG0i5bODAwGwv/5EPZ5/z15DfB/Q8NA9SI
MnyC38XaShcTb5a0nkuAyiwZ0wvRGQn4fWSCtr2Hl3VqZJhpuhQIdx949oYiE1XKIacVuEtHWwYB
sfSU51/5ga+jhJ9MBYbxsFhmSmzahUwWfdsBHZ1b5FVIqslTwwFrFFE9C3Nu5oy9WQ8rbLbGLS0p
tloFU9slPYf2gD5u4paqkkrr6hrevGCm8/32RuzGknA/Q4C1lm6pMI7ABPb5kDkIHT93pzeklD18
UWveXMyUKXtyZzsUqjfWZEKOB2pzujUoUs+I7gEd3MJPkBkdQET5ly8SxzTZh00AGSRcj4sYSOje
QtRYyNroqZlxLIjYM96B8kqVqeFz+iJwo0jXfKJZ2zUhZ0Xeci9aYj0+C3rJfFSc1T+JI20UhMl5
TfYWTieFWmmELCfoHMAM3gWHOHKweU8U9bHuZuSWL7BiIv7wYSEzN60LrrFQbcxMzAq2jRayKp9a
9P47ihlZTWO42ypp6vS7qUvmoqz/hxXWdU0l3tlwM7paPciA/ROtdgZIurgtrxi3gNx514avRtXF
F0yI32hNa+rExVaWRDMtB4UdxlwcrOekyqU9NqcbmQ9aTrKdSsLtS1RHVQKLvx4ZnEHk8EjTFtdt
jhoCIjAp39NQAEQ1NzQjDAKdjh7IGHdKFqo6N8hB3zEFd9eeQCpV6GaBAoGye0yfaZip0ln7QfAD
FoDwlVMiKxpU6MjFm6+6zD6kBZdeYKYnK0IQi/JHoh4yWDgHZa3F97xrev52Mw1q6kGRJvf3BlUX
6iQoBLtdu8MfiYIvBkjj/OExu2QDeUC3KmtyoYaiHzTfxxD4N3usUS0Nbl9+BccT1KXGsuNTeJZc
NmywVYbNsiYwTH/B3p0BtlIJmjufs5ZFzfTbtURylqDYkqxJ9Mq2SoBFRgYtg9e+T6eFE92u/tXF
QbGHN6UEJnO6d+OKesqAnXwIc3knapXECPCeHcfxAQsuqFwSDJJBA31U2BzwgOCMYqRu/vmSQm0q
RKR4BNstZJr3pfqAoWhZEduxBTvdWdREsRw8ekUUzi+ilOh/GgNLiy1CvtMduUFwzJ5gwH2W2mNA
7JFtFltDMeECHgSjbnc7sdL4kBx21OvklibrxcseIpL+whE1+SXqxxLic01Pz9MIqg2y/EK/lMXc
UXTKIAVnbuZ94SGr2l795U3RUC0bpWaafunXUX79oR7ywc4A0XPNPUjgMF2RbnpLSGeVqbhqeZEp
cDInzCKhsS16+TOKSX9a6R4vqvKKWd3gr32sCRvj26VYNRzqt1celxO0SKwXt/+PP41Ji6JUNvZd
YLGu/BUoeIDDrYGHWM92mN+rKlsRnyN/kXeIrrwmq/2H6w4PcZHgfpBxwphs+yAi7InQwllJfM3h
uRcWAABuOXbDxTN8ZJm0B4y7kB2BU2A/1P+u4xlQ0x2/DqeUhZaQe0SfxN3DBUcXEPuJv+oY7L9g
ZvNvXS4F54C6opeQ+Ow297+0iSbAsjONbh31iJU8Yo0SlesUufmDfzu3SY6o5/6lNENwlpBtyQ8l
RPRn0pdaOSD8mghxD6kjax8/kbsm36NmuRcCtpCRbdYbiElXEQgyMCDv+kbV3QF21Aqb1Y+iPXVY
+XUSH2wa6IjyqMbId/oByNecESA7ZCSDEVMwnJJEoNIlp/BmtC/mdighTEEfBN2l+GAwJ5s3sWn0
pKnT6YNrMSzDd2oidUH/e7iVVoAM7j189K5uSqA/9S6tWVeMpQPQI6N3sBefoYGTvIU5KaGz3sG3
MOpUUx04Ryvo4n1KGD26vYMHgYcY7yDuIp/lVdwfejKmDDDLE/59O9prCqu3tG/W9tWAI0M/YP+p
rIlT5qOKDICmrmi9Y7/LuE4RWQajiyQkwNRT1bNOILY42fz9vStgISVOxRmq5HN6me57V7rjQrxe
Zz1GNGx/3NIOWSkC7uavrtM22Jolf2IFsTNu5VxUiTqJWa05PIEsynR77bIqHqLh+UFFgmfrk8io
TwToH8+jlafK0MOMdlECn3H64zRxTutP65FVSc40PwTUm6Bpno83kJR5clicGgyEPDJDSTQ4Icxn
TMWh8GNyMylXYBxf5GDmNU4Lw6ZcMadCr3ep6waJhuSS+fvMqOo3ywmm0cn0TRY4Puxsu+wdLJQn
9ircQvCbODpxuYwkDRGcmw1P2+NEBh5gWRe5j8EXBy8UaTnOCt6HLJN22Kp8tN0eml0l3rNvi4XW
9QnxsmGW2at8pVTrBkjv0THhxtkbGT4sdv4Fvv3S4+afXsALhE0IbVOHa7YluRSk/jUOJr62CbhD
Lp2kHodjWMwUtl/1EX+WdD5QwHuXuZZ7HnZTR+CzsIZAnhMX6NpfxU2X7Lm5BfCMoaG2ROruAoxC
KQaOR/w5Dx4DYCabjBoeSnMbXfn4ZpuvKP3WSfQhpIHkZI4Lcu2aRIKWOzzBqY/0d5asR/HmmaWe
krcBnaU4sRE66NnRI51SsE23dUJGeszpfPPs4UacjDclglDaoOYITLi2Ge6p6roEmZY5YT4sIA+R
MH+eUVJvvH12QM0erOa32/hh3KiSqowtWfo5xZoLuz75wmB5EFuF5viHBdTcJKKs24yqmhyDp8TE
hyh94cenJOXskUdsgBfjPz67xa2Q0f3EV1jKbkPcDwAoBWuxXnw0+WwohG2S7y/n5hTZGqFtNRwa
+z+697GgHCgQSuGkdXjz5Jor8ImqLwuIrBYMpMkaM29fpYC/vkwcWaQhhJ+QpDZyTvkACaV65nUs
1YXPeyOf8daxnwA2wHjWC4DreUQVqMIsCBZb1hoDEsjO7H/oZkIepLpro0Vse4zZqncCsenrZNHM
coVwBzTft+sVognmuneKkVB5eSMoJXMWe7w084oFwBVp7ztCeGUXKkq+IP276f5Up6CvgKVvkprd
zw9mLTbVxVoZrJn1Zr7/7F3AlxgrCHgNU/AoOMD/L2hBXQHxK+I1dr3F5dUXbd+L4Q0Ss8MTzC4Z
PU1QvPZ/JY0P2stZexaC/aenLEMz6MXh/AQh280Ah5CDQcog0JwUyGhHyDkTrzPMiXMNO7BOUths
oXig21kEdQtuCu6+3PI/2HWDrrkyc14cBrhkY5dx8cffKFCqmSywjVUXRz8MCgKeIqOO9jjU0KZN
34ZsV728yra4n4+mv7Rlpphs3NQd0djHBj/nX9uC2/raSqQd9gNCVEqhDM0FmX2KDEQTbgbtpR7d
BSYNuvg9s1xSaiBtt8UJkAqcIZjrcythHXdY2Se1233utrS7G4srxxL0/A35H8VSdKQBOFk/CNnY
gLY0zPmGVva9tZ9D9mm+qMaMKDAoNARYg9IM6icToj3F0B2Q81U6j9C/wgEk8QAbp6DDG3Yh1ZrE
s6ken5Xg3oL4cquBrFWvohkIH4eD9MErXG2FWmIMkpvGlbq9oGPlvNa1rma3L54aIhsTbm/u/Q8Z
cafJlsXLCIzntHFCwpw6D/y0PyacbuF/yHMgbgjhkRaz+Tbg7gzD68N1HZOPJn0cJGaESiHGGSUP
HYFPVXRwDcyGLRYvd+VGpQFyPBtKRKV0wgdGq6zTFIDIzUqxzFWZ2mOOJ6mUrgQU3DS4+lwMxhfO
4jp3HFux/wot5l9hV3LtHFqt1KXg3LJsZsami1RS3D9JjULinUvtS/2oZxTkrMSYDzju77oM3ML2
rsVFLAaLB41rLHQRicJcDypYiZslX3c2jzv14trxDgWuaoplU0XOM1RrjW7Ut3lbxczGRof/7SqA
63El5k0Uc6NbTxp7iOXiOHzpcP9gtjlhfAM8tyAziK0IPVJO4HonX4OtAvcE7JoLbLnAiqxEyyHq
DrFmDuKgAj+euy+MSAHVikJseRje04PBqGIk9TGXKN6qYV/CcG1mkI4jKwp0ZbFhkqc5qb03qu0Y
mFlOIYdPyteHr6kmcOrYs3yTzpKNgbHvjNyvTjJcaF+IrDwqgOcwkhcV04y7lDzwSJ/J1Q0Wi1hh
nc52ZFIuZNphwc+fZq70UuMV8ZzwtcG0GUkZm6EnnKixZyjDU2aoCAhyxsmlo5Dqb6q3pEd5vEG+
11yBLlnGUwwlUNU5Rv/GWFlwM8cD5e25xNTrm51sMej+he0/w5Z76sbrMXxY77+STn6UGn6eeJ8I
i63BsSTPA7Ohv5FdzieSvxvg9N/uacK1tlMmDQMzm5+OFWXnHhTlDQabJQ6JsNn1pmuiush+LXVZ
5WQowU1s7wGPmpbPeD9mGMHcBNY99Kzt9RbY/Si5M7FZLkubCCKQuo9CZKmfjy5RSX9LHnZbJs9B
uGkcPUt8HkLzFXb3M5TncODlGpoUWxwCLu/MxIJuUskJfcNPbWQ7aB8MPlWMBJeDzafu45Tlzifx
7Y3Mcc2GBC+H4M6fbcAN29xsX7GV5LTEi6JbLRJTNBtMvInh9i1XtdZN5+Leg9tQs3fxcWzeGrAU
Gh1TA29StOVcN8K6d1WWsDVEX9wydci2ZeVkTcTdLAl+UAR+fdKrl2jNFqN8IHOu8WthDDK9zqHK
FjOdANjR0wDO6bHsRc37ohzVWOJQjtBKJjkKDNWUwR58CO74+AU9IhLi3gYRKkZinRFMdjNgasir
S0IQKkW34U7H9ycV4MZMNJyXtUzTN9LkHAbCU3odLpHb4F7zR7tDwz1S8jacvyylWUhfQFZ5Y1xX
Q0A5ekkDhQv7IUr+y5mnGqbOcS0UChQ/jgnL93Eq9/4/j/VbzjDPc51q3OQyj+98fvsKv7ZA+Oy3
bLgMqEjuPrTlQDqe2pKreDyrQ3Yei42UeoL98ojzXLf6UKICQbKMCF+oTd6fP9yR3tOYSYjHfPeN
kJBVXIUgQDEiFVQU8OVQGJTLsVxJ0TVZbJY8Wxxs3aflFhnC9+zG53dz6uzgqeVbxq6lL/DekRCK
FN71HHB6Zjddv6UVdlkPWkr3n5tgfCX33ar2/pRWF9LQkBvl8yEbPAuLyyZ1+BeuJG7bnPnaB2ma
9PxrwBT/5SnNR/X5kFcVPvml2B/8P7B7XI7/Bu98bGRNK+dhw8Q/AVN+bDBKNL7oR2hqPku5Tmq3
cpcPlWBZPxlCJTKmvr7eSHEGZoHc1r1NNnSxJ/SHmovwJG+8BImRE6WxxWH3AuB2bo1oif7ECl2C
BfjZRla8y8NxTcCs3GKcMpf1/15GmfERikmIidj4E8azOQH82UmUaTPtS8UqK4kUTMIZVRaWJGVf
08IIhaieHIBO+0I6rZZu3W/NSvtNm0AYynbVXKaMf+mrpBVhLnQWOErNpn/Zs2QRjt5Ic+VGqjeG
VgncmMevY5g0oT2vzESpvSs7MH0zvMdQT8XjPMOjtzm3XJl3rn8CwdrabU8GOyTtuev/r5Hv6z1U
UBv3s7D3A9C7Jky4dBKGj8Zjq/CDZ0x81wXk7DNsVlbJDWGgg+yceAjw/wealPaSUqwZ5FAjZZ/T
eX4KN343b0PMX+b/bJLyOQlVFAa6kOjOz+aVpsvzYFb9zB3pEUVMrfjAAcFcTwXPnRYYZ0u7EpxZ
nZO43iXAS/nn+yg5A5ewwOy5zB732jmqQmKO7PfokOde8TRguU2+EvtnhlHQvOhd6jLCJpTI/KEd
ejA5nHOImAEGttTshcJOkiH4gYrmScD3X5fXrVTEJPR0PsTYaCuY9Y6Qr6SO9NJC1TFqz9mlD5j4
XTc8abcMw6AyShBaCz3BewLlBjWcVALGe5C0AzmMxLdoH8gu3cYZnaJJEE7Z/p7+rbT8OjRQD5tC
mRUqNtVQWQBt44EJV1kl6wZQT2KlVyg74dmNN1DOriC6xsI4iyoRhgsLxZQN//Cd+sYf2KDa2Wc1
fbC3q5Jh6+Zwy8cgAKb7kzr6cis0+rKTJ948GSVaOE4HlOE1kCIKpZNZQXWRNg5m28KkTLuLzWol
WMoWQqZs3qEXEVhtTtyMOu295bmnt+didr+Xql5Y8SrXjWfPcs9MIB995YLdPpKYmFPtGeLNviiD
nFv+yU53fvFuHWuhUEPCI8MNojS88JAAPJW5L2Cb2j1lHADC5X9luvw8RsZlFgKjM2F8qEjICn5v
1bJLa04GdFxRtoTl3ph7U9Nk2riP4YofXP53EIyPAXY14TxcMJNR+chSPP06FCAqyl1Gz9jfinfG
uKauuKT8xd6vekBQY5nD+0ToSlTT0hfNf+5LWDsH907A7BqPaDF3xNFWQWfNG2YJemjRbxCUUKLB
DByXcAUR7SG8c0PpHDgssPSBWgCoOOMa2YkgnOI2l0VoLTsxyU4eHJEtfgE6DVchOMscohHE/I17
Wh0WW/cn1f7WNL2h0lUkhSsINJ2fIj3xAud/zsLv5HQy7M9y/0rhhNdVS4b6imuLnCXpxHsWwSh2
hxMBbca71MXO5bNNgcwIHQexMsMXZqwqUzbjDLt+qCFrhroWczkni1xajKHOsbP0pKWt/oh7aTfY
yQEJ71yTToUFg/cqeriSbSY6AppF31Iw8fxVYwsOU7bOvivnp3pMNABScCAcg82MB87GgTXOcQxL
C4elPOLW+KgTB5V17H5hErlVVBpHAdswq+x4InZoI9ddCdi5m5HKUj7USMkrBjm61GavHcBgNGnh
pbC6SUE7eEKr5jr5rzfxIh6u0QXFV162mQRpH212/bWS+xS3jKmUq4a2Te7fCuGU7TbrLVlVva7k
+aQoA8aZeaD7L4HuuDSvmLUVXppqxrdXp5bGyg142/KtGQbT2AMHJCP0gm5gl4gBI8tEqd2Z8JZ3
sBTMRr7+jSIsHF8AsYB1aUSCH32y0Xo4q/g7llWxszbshAFrDGoVsRfW2Npu4hii+rOds6mjVdOQ
Grnc6l6mbbQfX2/iqkTN9mcbPDQrpn+pHxUSAx9f+eJVmjBkxps3dZ5vgXcIw6J6bhiWn7eICnjK
sArDrK2jIc67QN/TIogRN9EKMUfNgr+FGnzm5Hzx42/RGRbWzOfqjkoqzb17Omx2T/RlqNSHDqHJ
9KWXEgaXThmD1lfdzbTWimZGQHzlQDRYUaTLxwoRMY1Sh31EosG5HXdkAFZPA9TBY3CfANCQR+m7
17q9U4T0Ju+DOKVacZ3FjfbV7Fx5PCRT008uJSn0aOadsgxfSysI3SP0BhY7YPWekd88MrUtWM4j
WlrCVXEAjXTuQDDdWjplsDs/+qxuA+Np/AyXkkgZDv3O/wjqx8rI6kE0GYO6dfPhv2bEme3SDD2u
S79D+VbSJlrwDdiFPjTW8FEYr6n79H8oYhJ4nSnUkR+TG4dVZ7q4yTM4+aMrcKb2wUd1fOIr+yQi
Riqp2qwigyfShqUwHxKQstBhj9frx0mgoeyqyuH6iX3mWF79TjXQsbKsoNNO9nzF+rDBaWVdu+Hv
ArYCVEkJzxQdJFxOhj1uSagFkszYxTP/PdE5yoXfsvRvE6IXAanMoupJLVWscR5J8QDRKo7SVkTu
Z4I801GBbt8ZFCHJ/SvUySgNih6B+yR1+lQ+zR/59de4kTbgJ2iLUhC31Qmqi+Nx9KPwhCUEUPCe
xmZ/cN7QB3r9w8oAnfzRMPzY1HbLyfA8VxDLzD0Pf7wyc7oUmG0FM+r4TPK9WEHR/Fl3ks9lsHW7
f429t7yqzhCkunrXQGyxFKXEfgSNgEhegFWOrUaRaH0p2h6MbRy6RL78lfmT0F9CaCNq/N5lOpuo
p7v8OgHd3s3EDrqD2QHZYIXXRiMz4HRSSZKW8VoQXt4es/+R3U2ASNIqokXy+NOBU///G3FeUuRN
1ER7QF2Qbe9vj0FqzdupkxBQ/zb+TCWEvmUH3dER22fFgM3HaVdZOuMON4CUZMG1ZSXEkPaRpBeg
JUBMut6cvtHhKQOZWzB4gtlPCUd2c1E3a/y0qo1OJppdUwO0+VBZ7dYNJA8juEIYyGdZDvxZcWbA
cvTgdgmHhMJprWQYjzzpPbzMki9LqFCPKeiGP0nLI3cSzDw2ehbK7+a4se1S2j61hFp8AVRa8j96
40sF8vBsMD7/vrXz5oltzqFPga2RxgACkVOaTwbYctirmWKAL0oOuQYh608/Z60Z4RkVaKCc35At
DvAlrUUAl2EVR/gNgWrdL3Pps5FxsXadkL37Vuyz2kWCpvYbDGnqV3DAXwK2LNfjP1DbR7aFNWaM
TrOA8lrVNCgTZshduQUIpvGdxekr2OtiKoYPkvYqRKLewGy4lJJnKopYPrDc760DmhdYvxZAhvu1
u2SJnnsu7ZGYpxHO/m1IzRyq3m+zclkZ300bV2JXzH3Zfry2q7slPYDsxoByG+KdNMTJizX18ajp
dOn9WeAkwRMYNp6jpyNmgSRII0EBwxQtQFCRWXqhH2D5IqFEN3oEF0FsWRPIPNsRE/A2mqDMbhNx
g5HRZUZUImqhQZ9mLbVMHxhY/XCJThwmJoMIrSJOLQAKhDmn5yFROg71drdj5Rfc3zYU9dCIyZ10
DoQi95/je4yPBo5RXMmNAGo+J0nlDf5zjtmErJfUuQ2vXFp+Qzocm6C0+KkKE4fpb9R9ZeGEfxj0
0ZT3EkZtsZ4Zb5fnuYcbysB0sPmjxa/cid6wLn6Eaps09eR8OfzqXz3sF7yTPRcaYXX62JVsAoxt
CtHkvrIJOpVhv/RQbporYTLugIfLN3NMxoke6spicsgurWhq2GLYpfnUwz3FRDqFOa4/nDQqv8ad
vN3DSBo/UEk/7vKEo1Nt3AdezF6WWpmdCqzPFPEL14sNCnF81MugMt4lrB16lz0Dv0TIDdPAtauS
4WZBAO4FVQtrs1ePEef5F2YyF6SqxiRPngQSM525PDe28wuJ2mewVIG7262Gi7Uh3+80JnBfsDgZ
pRbNaDY9uI7ePtfyl+4X2zm8bHpQKT74qmYwb4fRsSIVeAB2Igtn+dnx6CwKhTR7qCm/IDr0FRd4
3ZI/XNUHaTpHt1SZEpbwJg1kIztJ5QSp/1UDJZ3XWu20sPCbatYwqnmdEr+lGy+nYJTkKcSecSS5
MwtZe7XYP0so/iwWHAv4H5OUBK/GVw/S4tIr9XWUkTntncYRS5WEdpk9Fh+DTNH6tXrRtG3YagWd
mJ7kpABgWwH+qgYU7hU/OCv4f1R2ThDdsGqsg/+7OG2BLIf73nzDvt3yVxVr1tXqR4iA8hsZjEfG
3tvb1yO+cQHzIMTUd78zmod45c4s9gNp7owHKG1g1fIWjsN/YPZ0lYmf9PL0bN7442Xr8bso++PJ
h9aDMVoJuOw8SP6UOLcjw8wamgVVo+LltlzCf1S0xDT9DyuEJWfi1ldf/+RyukzC3syVlTLUGeNm
MBGnYNiQNGW2SIiTK45gBGFWgFkFFnvuExNmJ5CUc+N1qxIz5AddXDiVSq08LVA8MkUlhYp7C1W+
tB5p0nIRzyvqvJ/3JXsRs29MHdaxOVzoiNegIrargnJ7sciVMmq7xf5IGFIUK72nQF/1cWXR5tzE
tG944kZJYVDWt3wKCNVbfc1XXYzUM1l9if348R0jPs27/y7yyZyZ1mRE3dlJnLppIRKK2+PrI1yz
DUj4tDIbiEo/fvqgvEjdpooJeVGvGvwqW4poEm+kspcMd3HsmreMBzV1VsfQlqAF6HdnwWgzTa6/
6FVs0fLSozooH+EUFG5blInyFFBO0Irmj9bJfk/PzgMjdVGe+AJUmpQcZpguo8Mhf54FC3yuY21B
222z+P22GJAm2j2w9/JTv3cFQWRoDRxZ/2xsrfZJtXD0GSDFOne4C9KLYfT9Qa9VvtUu7p5WLNG/
huuRmWRWg2UGnAWQHQXaSkz1+8vLraFXXmgy5PXx/7alICNwHZV7rg8aID2GYLqbmAx/fHWklCsV
OX6kK5/gTM/bqJ/ODDTJkzRj/KnU9qg6d0dRSnm17T4pMt06c3VpL/N+DKYhK7YATsdTiZpQVWcj
5Nt57ov+lAntCE8siYf+s2X1NOOHayRQ5Nv/Db41FZy1me5ZrGYvUr0IFuspcXBm11SB5Nz1nUIm
PKVfHLQSQbyumwFqOfElz+J6/LtHgLdUSDnpoh7rlp2/ERgq/AiNeTmZ8Ew86dsfcU0tQ9yTYeNq
+CDpJPP/FG8xS2Y/IgeTyko7BG/2NBauMSbSbjIzdkkDnm4qUOyROnZ119Ecc6ENp2CeH/pwcu6Y
AF33z2i47QE1sXz/kT4kbpuUc3RI4VSVaZTcRRsT+NHwmw5J631pj0JoUt9le+Wn5E/XDKpsQbXG
6iEVChaXsO3aT+JNVQkLQVE1hA7DdKWgftUpwMXunVjw64p2d727f5ALbJqHbLgA6mZlYoacshZp
7qpo3ZJ5pDP3MljiqlMhBUqlzTnFvFe0D1zZKzh1f/nPeRIhw2mEC28hG27n/62WRN2dTpiprxFb
EpVaebJV2AaS7nCv4VMPO50jsI+lpngCuqkF2hSZtudBUmQm28Hm9hZltjOohBlk3tC+nWb6teXQ
V7GXN+B9UUW9UOO1dsTdWgSKdkEJmsAsEj0XbPWPcdW5EIe4PqOq6QJSeyfZHaxn2HtUX0JT2/gQ
8db5VDV62PscbYz7E+w+OTo7ktNsnHYxUIufoMsAMOCetvvFfcCrVQO885ela21LUSHEzs9HyF/J
KCx618U0Qk3RUq73CHmK/otcU8PQvWyt+NDHePnYO9MFUUlKoghEfbCmustof6QiymH87X7U4PDz
y4nq+oOwwC84demnyvLZ8gglJtv8CoGb1IzcLBXSnv3GYzXnA0mbcohtiOM7ErbTzCT+hUN6MVev
Pce3eGXDG+umOiz3cLrdGe6jUqdpX5+Tnny5fdwh+7NHJGipd9e+5XTwYgDc84rL+K4GUiJBCxVj
DP6hbGO5gPu9q/mprYRAEHA6HRLCiqz1Fl6yJNwWM62ebBVMppzuWq4APPr7sWs8PzHtCv3kfoJ3
22diHMfJBc08qVwEep0sP80HCppipI/VJydrb0z28/F3AY+sJHAKrbXdmYUr88aKuf/t60j+dr06
AQPDID/jH6tlEXpkxqj7sDhwUo0ykaDGLaE3dtVlX8aXXeAjkr9QMxuz0yFeCXiYMM82PG4RDUfF
em59UFYGkUaFilDJAGOVRxwfVpn1n0m5wZRqlFKQc7f8x+d36gPU1KJjgJZJmnN/lrS5wBdn07k6
+5n4jPYaV2UzOViy7Z4A7RffHrtLie+93M+qkiMu2S0Csx7y+Kj7+0sgtgP0ezoYxep6u2JBFH5n
yW61VI44TQUBcMJRNTqrtvTSk4hLRbfyKM5TrdnYN7aew6yWVRcowpI6yBKoN+R0AtEqo48hy6UM
KyWhFqXtgYd6Uwjv486iFMa4A4zYVhKKzi6rGoH0H2H98+dL1QxwN7insTTpP0TkgDZ+0Aa/Hljh
eVC7Mz1yfcF85t8VH0JWTq8LDZMXL1gf4UV3h59kKvtI5cjxYjx0lLMnwoeZwzstRniL1d5iRiXI
SBSpNx2PutBb+OL+Lq+qph12wwQjKU9uNoeBxx3w4u9u8tNdzqAzFqAZCW2K5RaRgGCi6TZXVu2m
E/DSJ+PCG9A674RdcQkvi1+P2UFhzR5/h3OHg6XEP2ikLdxo8tXFOd9Dg+T/JuHb34z1SoPIQV8U
u1vBPk/rPIti35UGDjbG7xpcqbv0U2XIPa1XU/UgQ+hx//jT36g37zG8sRIWT3xq6E3A7TCrBNbU
AdynPCRMnT2QGMr9Sd9qkton8kbeXYFVOvCGuKDTnDHTr7tLzryQD3RxLyJatiDIV0raMxTnLUo0
Azu2s6WUbAe4OF/f+A/o368n5K7gtumhZyqYg8HA/TTy/tpKk4WvBp5epnVtw/dsB/Xr1+hMlgOj
IMCmCsOtOL2tst3PBPZ5matHLYoRCczrDGqe0VnObamzi48fx1FLsPMq3/AgrS6QPCqJWIsFdItd
e6CJsZSKUpzqM7lX9/84tMXlJNvc21WIjwwnUy46jKAb3fPnnwRd3FOfthBAPHCQKfWqP6wHEy62
SBhArRPjcfBtVxiQLBP0oMqTSpGAnsxfTTslLVUKqJ7+Jw2KtBjpS5XB2D7Mfb45xQvfs6ETUYGU
xEYF8uyB3mw+eNYja2JdSlbaPVjLGuHFpMLefVJ2YmRlFlsLnFxxzPohm265jqG7Bx6J0DRDZF6R
M+J+rQWBiaPheUkKfv9eFWB1qnBWnMxJUtC3giNuhCILmy7YeWIyNCWJuThMoW/SmLBQj1367OSv
PWe9lJdWasJBXx1usthWkp4u5OXCvB9df5IMeYbHvEDzp2UntWJAcgHauydxIX5q7ppAph6o3FKX
05rR13/LGZVzPCMg4dy4aXh+EfxwtrpYjWB/+znb+fr49sgfC/BynbRnZIpWyLZ4hzO4Li0MTRdX
88DRu49bvci+c9neryuIqxLaBZkCSNM+8Y5IzjGmzmar9lodXxkgzgYZlumVz2My3aV9lhxHi7Pj
7u9z0bBOXufWylaXOp+O0zWrBiLHemgCxZpD8T5pri+3FsFziepMAfM/ew39EfZRMw95WduZi46h
ickyRMEFlOdj1KJ2D1Z7ifgELtteT2a9IoRmAAt3G5W/DxRKU7It3eLrgu3PrO8yef5PelZmUFBd
LInrik87cSTaWsmpirV8FXsVhIVJtg1WHGAipZXBgLGZi9TzuabriD+1ODSBczXZu6QBALnPPnlt
0IaS4KZlNV2ykpS4iHotT6u2kJsZ9dB8g+KQc3pi7I/U6cdPKQntHZeJn+3s7K0sgz0LCjs0/HsW
KQV206DWI0mQgboagJpUHH1SmWnc61HfKQpresWHMS1SsumO3+asNebvFT9TdoJiV63FqOyxzTC4
WNrbtYqx8TbomOHN0CHMNCdDvTGB0x7MY5ZsdDZNoQvMkyHvA3yGv1VvArNFmJ+XJ124LtMpTLjK
tc9sfoCIKPW9b1XO5vTMCKs+9wh+5m95Uugewq8clRL6ROg99aHutlr4TLzKMmzw1nIOHfBtkVLM
ODShZQsVumdayxwiL7ML2c+RAgeO2YD6+woIxd4xHBa9jV921U5Lvi/Wtf9O4FNHqEGcTf6P915+
TmemRIWVTZTnZWokSJw2PTJ1hXWXT7e4wmzOCVwRIM+gm7v2WhiquU2G9C3ybbZ7K+lCtOyLd8lI
urz2U+qnHwqF86nHqdjh8YTFuQpUoRTagHCGI2d+RBDgfL9IcOXdytwc3iHYlxXL65vYwt8n05K5
p2Svs2cr2DdhnV2Mc55Jt5pYsN3jwCilHjUBh/K5myF+W+WbWSar45l2FICEFjTShFF+pnC219A6
3kVnTzlfbIOpRsR1LvsBc3vHpf/GPobCZjbr5QCIYyB25j53RttM6PZZB/3tPsuO1H1ED/guE2gB
dCdeasJzBJAgpYd/p6FHMir1kQdtnKpIn+ZehCMgJMSPvYdj5z4CORm/3VDEHv4cXuyzGCW0L8/Z
DdB7jJO0VYlvFbTBULovo7kgM/BuQaX3q4+Lu62MOujXys6BEDzD49aCTfTJf2z0f/XlUNuj8iVe
3bQE5VQCN1OVhpjZjQOBeFcF21iRmAR/g/toLwqjSu6aP47OWN7xvKFxIoRzv8rGO1r+R4EcW/d5
s+10aYn+vVNFRNFdMrSMW/jFTS7i4sfm6bDisNI2RWrp0sM1hMHtsbbj6afvosdNXL9jJtb9vCji
kMKxwZ/V1wuE9HgTkJtK7uyMzY1oxZ5LsGXgDzKDO4aM2jEFD+Tq1KX7KYieoRDzQnYzYZreyP5x
WkKcjcepwtJjiCx2bYvaRqC8BDsqv4NPC3kLthtnafwgPH83PkXSt3jGj/kgXpTj95aa1XejQzb+
Fw1QrbyvNtQzNoOq8WcmVPxYt69oEd6Y/5Rp1trAE6SNBLd1UcUIVBYz32iZLHONuhwyW6PBv+k0
BsN6MJuZELm24Lq/oGMbnzNHaZMni23nhwAxxFwX4RJMJ3YXEtx03bxfnAAsdWGYwLqUk2OxOvkc
rghpVZCc/And+uOyWs3f9gpM/+KG1yPKKBgnNCjTQdY9Q5lSOKtwtfVq9w1xDwdZqBg/nkms1lO5
3ju3/WstEXD255aLon2Yo5eETpMEh97s//0hbEmNNS+8ZmJ5w7C2kHbp2Q/jFFRb9Ok+WTZ7wxdG
SDbNiPDzEoI331zK+D/+cEvXWJFpl3AfgGOEZ44A3vVlvLkE1H804RiIuDFKa5aNQblLxnJCVfQz
zktA8xy/+osLAyJnavrdGyfPtSXvSAEI6R67MFM0lBQ1g4UMBZ2pIh8eVcRvJAAiXxCC+yuEWgzl
CqJfW51MqKygjDoay4X05+m9dgMa8tVrfz6YFJON0zQQzZKu0CcBC+59ZvGTBqlh9ZcmBSY4QKge
nXF0rI/a3zlioiVSV8cxCTDu/x9iR5LnHccKZB6PIngZaG0zoGNrtz2zqjBy7u3rbpMoL8TjA/cb
A21wTQCEwfV1IhSEmsOECHndZDtccmlpNO5vOPSzzdt1V1kFKg2AZg2Th2jYwDePFdh0ViiEzMLE
mNwver6nhTfG6saNZRqshIIdsTQUnKKUJmqmtaluVOGWOtxmIl8OUEs0NbCb0go4Ijgt18rSndHb
FrhOg7x3hobpW6edxRoLrDtEr6qncRCpZq5l0qGbSsBYtqq30Mu3wlu2ar/3uRxiwjf04XZ5rLI8
slLk4FCN7ephfgOOyzlUJW0Ji1ffOocD1SjwQy44ApfyzOiVsw6dBTZyDFmHLipa0zneG9RTgsoL
JFevxFAJlFrWQsom6KCupqp2UrUMg+cABq/cCXLy8JZR83LgiCgGdcxt+RBiEFZUWwfSnStMTSd/
50GxEXBtloHWz9/fRXn5WawqitX9sg//nCWmViRGTJstRefDsZ0O8B9ZCYaP09G5xibVUiALjuOb
rwrYU6APJs84n+y/ADYx/Ya2o38MGponkXAC+64MKaK3QE6UDwLwaq7A6RDpZxdmc0ox+tZ4xqXj
vGCzZQViQ/EvInJP/yQNy0SBkPjYO6i0RJ/0YpV8Cg8r20PP3acfuNTSkWaxCC7fOxnDd99SRhn3
M+Iz/BmNv1mJdZ42wl292zhttYtNxxP9smv+rIh0zQ1lQ9hvT6PRsnkqcE6HXwwHUvQ6nQLIHA+x
TdQqRRFtGAYaGMwhQ6ufQJHgOHsyjDfmH0XfhevbSZo40aTYq/Le57Dfau/sI+n33H2t8n1eJln3
o4BKzPeneFHZniL1CuIaQBj+aVdJiIuL3xNwhKWOWebsa+80mh5dNsHCb5oxQ6c8nEsnaEPPBD6d
BAdNFE40HYWSl8fTY4UP1x9iEgI40WbbTkx4D5HnHmNwkwRnbci9HTByeSHWSUkt2G7W06mAxbz+
6Srkw1NRJw/vKerLkuaQ1/tKjDzO+I0dwuvoMzqLVmLhdSqfD6aHI9Ofn3uy0Ry6OT9e5LRQyCXM
Tv9NO5GDETWvOLOQMjT6wIdN7koyalR2eS6vm3Hmt5f51TmmAk4+oUTiiOPYiGLWdLwyVwJELwLN
sTch/JzHCEkoeiq6caQ6YCmSRhjE7ESI8Z2iVpWSUcZ+4qe5hAY9e5tMV5xuih9Ki7dsp/4vtXRE
Xy1Qx3CwY9hIaJ6Ql+LQ2UURl7uvkRx7r6bcEDGUr9b9KqT+k+erclz1BoY+6fUvPC8+dV0/l7mF
n4GqXrr51O6jaxem4BTQenBYQpT6vgn2jVktFV7u0S+R5EiKuuuwvIyo20ulq5heJ9qqqM93J/Ks
hCm6pRZ7OzzB7GJJWP2Vt/IqcvBGCYJ+dfk79MqUKqIF+fSPRZhjvgNh0hFp/ZcLhoy4ZIPlLGNm
NyWJvtNLflhliNUjdPSO7TC4aiPwbUmYj3Vod0SZGyFnph2OEEelkah8HdhgoxFjDQHxosbyM1t1
pRbKavWg2n3dpTNTEMO54kFx2pG3bynI9CIf1zf4OggWyMOur26HfNzDXywKr60BI0rJ74fsOenU
efPJcQI4xt3+2Jb16MLDZJIYdPwyQrIRzwE8eoT3M45Evx8TgPCeBOFAC+/bdN2m+m1h72viwSSR
UVbosIUWaT7yvEzsWugZ40AZ1JUFiQDsLCbBc6p8et8sq0z9k7yoR+E9fuWysbXIsjspeH2ssjgc
RHcNn3Q+8f85coo49ZMrg1F6jr0klB7vS6VbROXuKhyGthK7XbPgC4xWjMSjj28VJjkd/z56MiBd
9NUKSeaYeW2aZDZ/7bjZ09ygOcVF3Pzx4BIQMfvuUJ8y7i4xowzDtFiJRpyk3aIrq/BuiDIQ9RHZ
l7zNBL3r8s2PZZAMHEuHI7k8Kyp2MJZ+Y0FBL26SH9mOeeFYLqkMlHupZy6wC79Xr8Slljbn86bt
oUzNY90/w11lJhulyB4nZPlNLnMqSpQgibFBWMZviHQK7TArFUYKPT4jBSB9hMncX+GWUUrGRClK
d/epHT5nNMMbsbgQ+isBYuv6bc/ye0cmO82+z7PIqUiE9tGg6ArDDJdOgeCYe3fV6Kmt7BAO+Yjg
2Fl3bSSNNZHDt7ZtVArOsDDJ+ERnDp0hQadoPuN71GmnWLKiDbn0RZ1tKbHChEhMEb0WGJtP07Pu
7524X7CzWTI6Ajz517cZV8CUfPDj9hLGYF18pvulRS6kmnCtgIVV137DTszFmLEq0crkCwZw/h52
+BjQpfuQUDqvhsWTis+9zEJmEdRZo4Pq9DmWeaWU2sMmBVpzvwzvEWsZO8a1EfTY0cYPJRdKRJTj
j7y2w0iCPlSAILFS6I7CkxF06NsQ7CufpAkbStcddrPCej2D4URTB1qZJz1BbQm6QwU9h4wUj+6d
BtukhMJmdBPwr7f9TFrFlbiNGB+n9kJHJ6zXC839QSSoiXFlqVskK88vjvCTdfANWNKWcJNvrT2i
Mr1K7Sydn1g6bWB1RXqCWAXzvmV/pf9f+OY0gq+NEuMvg3Zl0Zvsh6PUIjaOJI5ZbiLKFvyvZzbi
0mICgmmusuZcsoq1d5/a45hOLd3I06bYRjUGmhYfqlHqMLaJGNNiqTDZXLGZ/m6ZRGSIZBFiT4yQ
HHlfo5pJkxdJW95KpJHygpPbGuEZwqc6OfPB5jgygNvuQHnjfziWOUMupg8TGOIczc2LxQTjHNQG
c9PCoCMq0mrc1mMbLporeyXc3l1m2Kz+8JrKHa4ojhqz4Xs6rzZIhxoX9CTmFK2/szChwXiFhCc5
9ZhZflr7lcYO3AbOYm8NoWHjT/7KhViJeXb2o+PxHuziFldmASxxUsAOOFe3goI4jtN6Jo2WvaZ4
CuzqsKGFqqJo173Udf9dE9facMuqwJiacZV3KeWVWQuJQDf9/1A6hYOIi/d4fx2MtGsY5oSbfyUk
V/Y6v1LD30rI3KLZAEgi8ivjaSzFqbJK7yjyWbBfPFA5kquci7s6Gtw8g6ecDw8MJhokNyT2QYBA
Zo5z5+tdI7PG5vxhATp9VuzeFyB4rWMDeO/eeLl2rSxNoyMkzzd/6wxcbLOBNtt1k3duwYOzDISB
bJZXxhIOrFe+gJ3v1l4Dwz2AO9DUYL5RlSClqUu06dg9k4I3MRxPgX4Cxt4rnWsessdYzbyduQq8
k4nTheXnRkpwaiPkkyynYd94JgFIJXFGQhU9mgwCnPibmrtdPzw8tcT21nj2bXl4sgrqpCVsCIiJ
24/IebNvnrIKA90rBm0PfJaELAolIGhjW0LrRUXtuyq+quFk5AUzgbEs5h4jrDtybb1MK3a1PQjn
POWxcj085dAO5+H/DB2X08VQNagi7xK3U0hwPbRatm4FCmTepPihtJAlC+TU1PdsFaBzFiqWL3Yu
Oy8+U6naqgtuMcNmBCr7sNBPVDaVfkkDCjoYUI7o1/wUF322LDR53Hq/+GV+HWECXc1S+icVI+PZ
AhdYkdPTlgT7tFl7SLG0vwS0vOjMj28JeMy8Iwyy8ZGs4Dsbmb6a0S0KNLDanwiyEU7oJElUcV3h
bnqRoXDseffLGvmhy2NUgk6+j7AZL9YOVh9mNVRxQaAwXtz2/UtcPmjCywlc6gFlwr+XKsMx5n6/
7S3E9xiprpebjyXmb/b3kLhndg41E/RU6gYi3Lfhgb0IMsvZzUasJVtGczBTol6lyqaMAMTHCU63
DeTYUaJZbf/zMMGs0r4jcNjLANsrd2O7keXihkGU0wudmgQp93WQQTP6YSc9U9ER6EJd3QM5aaIU
v9PpskoSuuPAgqtnKU5x1cMFwH6QVAz7H9I7GD5PsgrFc979pqQ17iq5Hu0YcBqn6U9DfuRgspo0
rxy8VeB1tJVCG5+Mjcbj+EOncNyRKIoe2fxxWnYeLwcwdIcrtRe2Emg6LwLYz23vRMjEwR93UbOA
pYX+uCA+nISatEa5xczJz+X5uLcD34ItS1Ebl8utCSdxbfTUZRqW8XD7L3bBElftaqQKPaVENwFz
qAYWpMf2OntLSkj/eWwCVIbhqtOAT+djYIyCfAvO7NxXOQgX3mVqwQUb+rFUGUOqoIGGX8nLC3IZ
WJHHfPl2g9AeuGfkTwUmlzx/5Qgnhx3LWTtDvZUJyCWr4El9UJVMlz1vzZqrg4FGMxeqMPrtdEXR
etAyKk7vUec+F86gdBiNB/5S5w5jTeH7EVJqgS5eCLrBASkQpohYc7+KdSY4p2kunhHG/N+BDdjv
8agwyHY5ubSZW4gC0cLhNWicZd5fog+qlGS7qOsH36XPS/IxaFtsBELTRnF/Z00HYiYd9GDFKjHV
h5eNtylxqg/JMuCgU3nvlxOnAtJj3blbVveVE7R5TQ1Vi+ZDsIRvvue9uYeCpZFa2KRA9vGPyvdH
MnbxqSasjmqO4RyoVCqGFyPHF6NsuCgrZz1II5q5qwvk8ZnYKY9QRYJHkEOit33GhrLMbl865QW8
yP8hgOPSgcIjBg7zihuuW2WEWhiyIEm45/o0qoARmDx6pZl/XQnHDkzOIP8br4StC7eQNjDlykGd
XWEbZi9XF289SXJnUSsOLDZ6Mwij2wQiOiJuqgrm0UFTwFzcsnjlAXqtyqmorATsiCNjtjaZYRSX
47+8Fg439CsN3TCQlqlSkCLmtvDxAjC60JEvPnrrwSEqIdwGAFAMMgEwjr4cyxQhhPX7XXlFY4XT
Nc0fdrgyQf4njslUcUMUvx2QP4a7zB4JCASrKCCriFSLJdaq9td6AOamYL6vh7FMT4bEGLhPl1kQ
EvlN55ThMQAw98yKiwIhrlwuRLgBhFioMnHC+r7dKXhUErf27zzYll6bN3uoaoQ6yb5T/wBpo589
9+aDZn5dpAENK6E/nfzh+HKoVzpcYhuU5pomhsP/juLrBp/jj9ncbKR6o+JOA1g03M0cdCwGF2kZ
gJMQB9OoQcP3w80RgbHpp8TrhqtW3j/e5Q8Hb66AW4G5MZB89DslIqse8AGgFZ2I/I2+6vLPb9aO
/hyATJAohHePIq0A/LeyvE69PVu+k5LExrOxg2kQ/EkJaYJYH838+NBFzdIwSb4xy371CJ4bguvP
q6Do0wDDAwSqbec/NqDf/mZklCrBz6OXOQkhlX5OLDWXPcPSpxF36eMYcTFit+b7nxhy9cwcpI/x
ZOOfQ1WaxufiH/9xP0nZDH0QoMOQCqMr6Tch4TBF+6APiCvRBI/0dMIp3f+orgTIBLF3WHDMDG+B
MuhhOGIDDSnO/gOrlLpQW3jgTL9roPVc++ynGclkvQL7K0V3v0iwDzb9lKIiY4M3jM1bpPUC4YYZ
m/SODMaLTDsYnHA2IlZ8sKJhZ7js/lEgZoy8M9OPktE/hTz/Km3QlGkl2awDAqXQvbSfvcQVfpm5
mQCGkWkLVsmyfuAiXtP8pe3yg8izOFgTpSa3jGeQ0L/L4VGyrF1HaZaQBF7ABgvIFqzNj5hsp9jN
wmy2Y9oirUwKjILqJYVMcfFxYyRDiyZOM60Xjif5PM5dOk8z8C4EMu4n3ydNH1cybyrMrB5o54gX
d/OovlaoSFqymE9nPvX9wcq7alsqSYVSkT9UiUSwfYDlA7XeiYWBEyqVuVpD1KVtRHNiuU4yaP4u
roshoBxGpjWUoaF6vLVdERtGMoCgwm2uMnATnBrsTSgcniU1RHIX36RBMJSqqe6C3oGrPa6kPQBm
l/+DJljL6kt29m62M6DvOmwWY8ZQEjc6DIiHEYX8soMzJO1pKTeIit5DwdZ9MiLIAwD2fn77ONIw
yql4+Ch/b/oZmY8HtUCadSBxY+EV7Au/iI5ai0v5iRMU7/ZrRPaKZviN7xqtAiVbQiShgMqq1HEz
oRsDiRNVeSARr6b0GQmnnKHc6+TslBx2pyLUTtLpl8JGG5RyUuCSkMDLHL9rUN88BZH0X9UDMjk3
VKie713KshL3zcZEhh9wzOQaix9zeYRJhw5JeBkG7hS9LCEoG6VttNvnKnoCCtzFeAvBXxQcNZ8p
++oUgm7pS7XMYRPRiZrysfkWYz4mOanom3iECUFkbd4RxeBN4ifX494JB/h2GRR3ru5efvp/NFoJ
wX5a4QSH5SvCa8BYbo9gIaHs1Y3khigqGQ7lv3319FAxe4ycKSum0fIY0LFeEgUN62ZCdAXwamgf
eSJ6iitm9X9knaNNQrcL38wz0jnJSXL9pSZ8jIkYhlOdWaTJdGASbIMGmedQcI1y+Ux6vV22/Q3K
odQdHJ+rzxKoadCkN3OA0zXgvQhWGKJBvZClf18mtIVRFLVV/lSl7+q1K6lfKjFvhvpn8cIkGx0V
qQhv+oip1wdTAROGVcC0QBlOHQ0LOl2PVTxfDfwPtA7PEsjkugWUD9VSt81Wn86eAyfY/beYkh2T
vytIy7Yl2yFvzwYSAj2PH9evVjzKNuCDOQbFPB3snIy9NKoJLcNrp8TrJ8YrKyZ90xem8IzsaC3f
Zknl2s4iOisqrcTr7ctYQU1YyGsywM4ywiluSBwOOK4hr0wm6EOLse0ApgxNkrRmOK9ZLody9+Dg
w7G8RlwqlCS6BA/5U/MBZQMLtnwLV6E0oPc7MmXy+oHn1gm2/IwwtpWEovrG/8LfaqgR4BnPnHmT
f+xX69fP1clHuxicHWd0qfMz7VeyI7nXc6hBFhst2fbLYXexEycf5MjbEVGrDMpUa0BrAReAu64Y
rfxx2sxdYcrfFLww/TsmkG565TqsyV/CUMD/7rQJq6VHoJ80wn8+gH4i4Yq2q/SsfI2yaqyzd3OI
ynrEjPN2ShJEUzRX4NMHaBoEpJmhTbu6qo7oKlEj+QnfX3ZELXGOEULCqs+yzmh4xPegKmMf+DiJ
KaLdNmfJsENgqXosJ7WQeAMBP2XmerjJBKjN1KgWnCGyt4MljzavEwhrczs38MCECqTo4txHHPjr
OibuPXCaYTk6cKybMJwZtQBTqws/6IPWA8wPKeR4DuET+EbQd7azGWcyThaSrD/yIsgl2wFLnFeO
23coanFUoBSZEoD8goUL0CKu7m9DgaWgZDrlyM2+qQU39NODJC4NHG616Nf7A9QmBlov2jiNa3+s
1anGiCUL5MOFSeUFGowtehzrWPciN6Sghnma40PqpOxIehUqYcjpJii3GXmZD2YvPy+1y+szrv3M
F8m0obs60A+JM3Tp539chCLx9mzN3Y/MSfe9kQKkth8mQmaLM3YK4TlhPPMLCWTQzA/diY8vYb4U
NbackX37EM3oqrcw4n+WE4GMZbxK23V27hgNXZC75nLeWAzNlus4aLzR66NIDKUOkYmPB0CFSAb+
rPMh2J/qgfX0dTKALs7A/MA6ZojNthtugukpB2q/zT47Qw9P9PrGkScIZ0NawFykKwaRAVy/G/+n
b7EWX0gywD85uHGxULmJPVKqx0ii7US7n7xAIhbX4xzpPAzi9Nv0wHT66cDz1g9li5nRKDVi4T8X
fOkUEyuSx3ayySBomGCzM8whwdS6TNjZTVOS7ZYKaN2bY3QtEhXf3uop82vmrYMaQkKKxbTxGmJG
kKCWFcd9NenDAY+gE+s+XKeyyo5dtu4oozRPpAfPgmfHiugTj5JdScs6AWdZKXRIErUFA571DlQ5
Pc4C6hU7XwiNipGjQ0nhK3zfCyD7jaIp15dF/Oa/hgkzZ4jzlOqUz+ZGcUajqBY0P5lBvZGa2juP
Y2RT6XsQzm93kIz0mN8FeZirrIUfDyatZRmF2WV7ByGVBFlBHXqeztYeP9W18THA0Oag5Nt6+EBE
UntuAaKYRzBBNi6guFPSeoE2QOhbyRWMYtscANRSIEEqePa+B8lkIxYLVurgyI7Tlv31rgDfzrH2
NIiOqR5dR4dfVatFARBXWy12rzgnj8T5O86bZOnq74G0+0s0FYCt7pcQNTmNsNi38WXS7D+IFekU
09FQ7CHyHOO5oSsR8eDbLTv8JNVlFJeIPPjHJRvprfBtaFHEJVJE27vQ3NTTH523ayyGpUTXNrR8
/VIWYWG3vd31T3qUTN4gQ+05ZevYY8gVmTZrhFXrR4HV5c5pzjCH1gJ/EUFF/Wor/xPdkPFtcCiz
9kPGLk7HwX9Aw/OsAsylhrWd7JnZQdWru1ZsdV/MAq2usqLog8rUlddEZwR1w0dzz7At+CiCUcF2
LYVAoT+UFvPisbRjuGefQwNPWuBLbVp0t6EXGk5StMzGIgQffDZT9unJ2/B2Kp6iwm4sMYBS7wNk
zcJaj+NnetuGLg1yoFjo6PWx34QOr4DDB9WCXl7ZNGC61sCvUi+zcE/qt7yEjvjido5t0/VPFURc
FfocVDp4QpkZQr9fERy8RRLpwRyki+lfcIWIX6P32KwrpQp5a4wYSo3KmYE5GMx5ikkON94BosOo
01EZ3JJNKpci88ESl1grfw/qfff1v6VlOcdptYGDRpzAv9F9scJezI9zSnQ8aaprgGDwaA663lNZ
nSRyzD2dhqSAAsL6Ovwgp+IYG8bSa+oEiOzEONGmBwIUhN/B3kMANdITkM60CeJtIb1NV2Zjeo0u
gfCzjb+rgpwcgBlb+lfkWnYGCYbsLAzQcMrN6qWZhItWEi2uHq+UIHvigHl9sHsmZ0OiIDwJwGA0
MhOrXiPCdykrQLv+lINxtdFtWYxNMHTD4cjDBv9G3I3+vHKazm1HWZqw6HoAdmbsNZhJ0q4e8EwH
FjxFpoDqO5m63Js9RexRAiUHwa/cp6hDhj/mPBhCb26R6gIuLnQdVcRVMO5i2GxR/ajvsylQWoMu
FhVQVTqPNuVqt10bOim4sncE4jfzIVWfwq8F5d4OcmNIBfpe6tB2yfys/bdiSlp1+kFW/bfsEi6x
OWVfWtVyxmE2+jPkfA6feeQkxIM5e4H2ETk5lC+J/FqPWwYasMOv4BWzTbsDO3Hhxpgqx8m687/h
54CxkEROqzPPkHiR28mwjq4EWBjI8XU0A7GQOLk86iy92bF0Q5GiNthMIdHrGKOYTl8WzMVbl1Oo
ZFmZnpCcA0wjWqiJF4tTFCHzyPXdNMVZEBGxZpwRofxjHU7acWy1o4aPzEek2J1sjl2FWP7PYCfl
hfvKx/R2NVXEKMU7OjTXnkwBpy7bf2ULTxGHlElX3wRCEjsBSbyZpJvX+HqvHJ7yC7NF3xg9p05E
M/nsdPAE0NrW/fX1N/EgmW+5G3kwSwe1PpJIORCYlHT7Y16PdvDlLc5o5g747ZFtn9+poaH008aO
6+4tnvGoyEuN/SiyTvwbQwrYxsRtUS6UVvT1fN7a+ejtDRF+hdLbDJ1CoTVQogs9ReXxh5HEZhID
e3Uv2VfDHUpsVG56XTrSkqWqN6Wer9ATFqNKaeLYS2RXe8UyxpT4zyiwa4/tFNiR2aWTGVFno/3A
WEOWuTaNcU9IG0vrkiLOBL3fNRWh9GXuMkW92iFmtMpl0nJbkbwN/2nYf9jxJ5QKG252QNlzi9qE
2pMtX0jRUm7/4mPAbOLyv1XUD8rAfQo0sGeKoEcJgWcyycsNr+SUC1K1SXVGcw/WHbOkGvUPdVWx
Rxc5tZ0CGi4OYlwB8TmTookuF06+xkK12WPcmqs9MUYfZ95CuCr5Wr9Afdne/jWB9StOcrzqwPUO
z9gVVtQpp2oRQTQmEYMDCwKo7CxIdjfoUR1deWwjuHWHFZLZAguLaLwY0L4OS63WNI5psFQLQJ/k
GFcsry1yXUqXA/Piqnl7onsYm2TKZ+1fv8JLdKGtEePteC/j+aqd3++LRN3r0m7rKyu9g6vj0wh2
egsobNNHAlRTwPMD3qvfF8Myfwxpqj9PgyrxsuSg77LFkEl9cyWO5lfVexTZTZEr8zeE+RCW7DUn
9/VSm4KDgeuQXs7Rw4STvcyIvQIMmXNhFcwUnKfsAi7NHyb1uTJ2PAd4j9bqOqc5O34PhyOsaijG
0QL5msycKc3q0NqinaEQS5q+rT6FBmqZCS7/wzd8trt8kDx6S2Atj7zj1SAIhh2snrBYLcvaz/t8
1AzY3gvPL2I9zJi203cXAesUpF5kVjaS/NZminBAwCi4nLc3sUPHdvW1VJj1HPQKdc0QI0xnA2C5
CMc7VAIJN0KkS+rvJcvyAzsiz6fNy0Eu6dCvWOoUX+vaNdfyTdXelMf5WbRdDL+R3y83xLZnedrO
mJWo5X/EEZl5gxq9nedKprkOzf0A5ps7Yo1RDK7FJtGK3hVQ6onl3lVh5/S89WBePXTxLWR9kT21
DSYoHxuEzMzR2l6h3BJABC+GHSMNrbYUPb8FDejh4780jJDYXHZpn47UzGFWucN8jt8dG4cAqnEj
jFzGl36S2KE56oue28jXAckS576J+lMgzyGrDI8E+xiQ8hKmBo6yFbNP2TW0rTF11MuRInpzhWSk
86p4DcSmjvovwve+askvQO+694GhrhTDrNCBiA160JriPoqAhOgDYvPuxEUlUhCDZVTqD/BYU/M9
+KaazOcpLU0Ha0y5zkEGsrqr6svnPy+fRYbhr1w7cRz9U8xrG8lxBH+qrMQZ4OnHMsPADaNCIp8+
eJujKoUJOAqHbmngzvg5JplbtNUyXaAUYqEyKHUxRTLB8SOHQVwZjEOiWqxCY9qgpx7UU+81HvkL
MISZcLG579Gcr9rXGT68MUz5A2dtkZhWozS2t/lQLHqSHhxa5pGILYdf0qvwYgAMuuse2U6wNTLe
l1jSlpr6sDCFo/+9yu/+sKOpT+HLumbdT/3AZCsizeQTsD3Y+drRv72nokR4/QhDTGyaXnvTFc2v
3j+6SmE12567NS9AtR8y9KRJQqD/Y03A1n5EXEGJBGcoGO0E8MzIp+W3nm54NoHdEmm9wvmhbO5Q
ndCBvAv4xPncfHBv0B2oaLPXCdgGVEZSPbDn9iD5QjxWVToz4N8uJTBSLp4b85D3PSuqfZajCJXr
imfrYD6ceLQkTyoRTLpsoIeNuqJc3J9nkMNAh568seDXDfuKXLw+uv3cqPA1lzEiZmCGtEHhTctz
eTGwxNt/fjiqH/HMiwlOvIVpuSEKAaUKjJZAsWzCsq8lWnf+QfOX3IT+WI6gMbwvdGNCjTuM9Ym5
dHtKP+UKd5Wg/AeN0jeSz8CBRcIzfocvQQuT5Pw4KaFMU5KRN1hr0UFfwIfF4lEbPHmDXNZTdusK
BAeWsda/ijR58XH8qwZNig4rV+Px/YT/PvMmK1XxPatQBr1UG1dD0TiVBeqWC+DP9ixQg3lKj+F/
YfC2YvRlxQPPCbZAior+Eo1wgb5JFKvRRA/hlDQ5hSCzNBeFDiWdyQNDMbtoTyi+tuQNYzC2DkXA
iYvSf8yuEAg3WNpFnuTYQxX9PakpMVzrCRrhctCjOOWRsiQy+rCSErQa4VJRGfTiuUcSadqYn02h
+YX27YYBcskJYK834KdlK1m5giifqHV2jPsILkdS/gwt4ifkEpduMkAUS8AizrhMj7z8+oYWXYb4
Tp65DE/Ta+Bv4BlmpPErDt616JTwQxVnzVLFa/tPZmrNXhD1+aWE5keIPJF1j8P9caDl/h57edul
vUHE+Vs/MotqASTrSt3AuULeKmPNLKNibNJOktAYNcIsDs+nJQaPOi6FJ0NTP+Y6AImcSmfymWlb
QK55/xEmx7eGV246GQsKeAsUeMNkfinwmFtVJz6us8jymNajwPus/Ie0cEWMVoYaSkY1FOd8BXnQ
YnjAWtlrgXZf27Egxz1gi7jdi3JIGtGkpDVukmtCmiR1cFGSGutLIypBKSIN6RGNG6Kr8Ifo4NNt
u3XrTlWgEynqrw+1YbkDLrHDapbrMqZpTglCTzrCjrgRuhLWQQsyDMkDezjevT8dggzwdkx9qV47
WWBu3IJG7vO5i0ohWjfoYOspFdXQDoJjrwX7meXBEo41sqBONDPSRzk1rdGRSqj/xdsBZqrmQ9nv
fPQseELEhkDw/tOaFnbt0UXNFSozEVsfAjEgx8DTE05iMJDncxTqGdzmOFFi4MdSwtMoD9uWiDlA
dhPKLjqQ3KqnHJ7AluugvSQcKz1b849avLlspoiUtu5XpHTmKqDnr+p2mh7sxe1Ctibttz/0XXK7
rcjiOB70AoMJpfsoYvuNS1e/jg1bx04NRuPOj5wLksda0w1PYO9W+GCSx0Zv4MH4DXrkU2eiIybn
SBelbuE6ZoPlTZ/5O+z8s1O+uBUpzWyco69fZGkC83jgwpHVmm8v0M/LMLwkd5qJ/gYvZeEg7tWY
EMdp/vJMbNopAaxWHBvvUGd1wCH4yOnmFrLoXhPS1hdZ9OyhIO3kh0QLJm9UE988aUfwfkMY1wnG
Ttt/65r3av/Ih9guH04E1r2c/cueuXcon4hmljnOS1JiRGWAbOjcx7ZiyAE4wGUN/gIAgUcv2HbR
n7xQoyyTRKCX7lj/4fJIp1TSbEBP+JYub0kMXTQq9xhOHv11w1iOxO+sK23vdi5KXqUggFcS2q04
s7vXz2/Ph2EHLETWioO7KESrc47+DNMDqSLf4fcJTwpk+AzzGJsvaJdKeO1h12jABaZONNbHbpkX
0Tfs1bFTk1ZY54cpVCNT5r0pHx9UeBTXIrUL04ipdXYzFG191up0nrYXfpt7ntfMB6gXFy1MydfS
gKQ0hVM76YpypCJO2rEgNIDVn7L+UvriUZdSQOwu6DSKJzVA3eFYQYz9dw8uyDf2DV+b+JuPHaFu
e9UurHaIIDzvNBTJ4Ul8+C76r0o3OB2M/5G89JNlEeBIMZiTWrkC8CRT24BQwVFcW7UO+nrMVoGJ
mGFKJ0+dOeBI7pBAMwePO71Smk5IJpDfq5ykUkupqH07jBry2ECwAn29bVhNpdHQIg8kxf/PJiQ1
9xJ1PaPpeG5VwYR+59LlFUtB8jWp50Je934dGIjDvosNOhkFmwn6REUltC0GiPMPn3DTMNYM+6b2
5qsATp6qwgM8kyWZJHzSsF9+G7lZpR4N8nY2D0UjO7xb5UrD/IfH8pzTXaFiTF59sb8B1rYpaqfT
aZPVQyxC3nxvvLouGOCfUy0yGUSctOhlLvQEo2XI7XlYNwcIye4U2rdrV8XRPHI6Kbn53xPVb9r7
tSQx65Qt8Vd/pMdxrtdihHYy1nonSJ+MAoIpYVttF1vmbAWCPQS/E2AcRjPnbxs1kf4ojNLxBI7Y
cGXjvzKW+HFvrszqFucWAxgFluFS3jehMFa/zDUMG/p3DH6r7TXZbdsM8ktCorWCUc2XqMhYqbj/
07Mr4lQy/h5jIETe/GxXvvtsyUMlusB3AIIukIzMqLHD6rx94CBM9EiiSUkfxmeScHyBdxgkf8pQ
ZYIRkLGysXCUz0cNuKdo615NSI8RLa+Z/A057UmqsVQ/F5B6MAsyLXp3xyIhhR43SJQV4TsJs+Gq
D0utO+8KwNoKHg9P76Ye+tWDVQoyXkeASQPuxNvc6aR8UOc2RtOlxcmkJKtt1MkT1bXQdnVfsyCQ
1kC/vOVi5NNyIAel1HFzOQqg2+f9jtR97xUzjaLriZ6R13x35n+5Oh/ejTx+CZDhToOF0/7QTY0x
tfrN1Xs7jJ4ukHISu0c6VnJOsw6uF4JiSyPLBbPv91fRRGUYAl71Nractr+UhOyRC3d4EWv88PvU
UJvP453rsM11GRDDjrM+qxGtPTI7bX27DiQVnML4khan7Dq06/WdYAE/FDNPMhySZEpWpaO0LUN3
P4S5ta+4GaYWbFk6g618+nJIXvBnfeHOuCWx6U37MBq5aaP7wo4PQCA8KMX6CRS4KA5/cEYAwdl2
vXGgeudT9jbBg7n0KnxXF6k/nq5zTKuJ3TCXNecQxcO7cxMWwVZfY1RcF93yFOclKx+7jh0BKAd0
uuIdUq0ipVtf1Rt39MfHfSWKiu61/mEcJhWe0L6RKAVD7uY+6CzuEZ5ZH6dlAzjOJebseYLOWDKo
1gWO3twm1Y/p37lIZ1avX7yKiTsslg7ucfEWs5NFSZkxmJ6CySPoHKwKRVZD4DAU5wShIxZJOItd
It7faXj/rGf08hNqHTwEdA2koWvnYI3TNx76Pxw3Vh2bNBDo3LR6EEcj/SYyZnEh6A4fwAOdvyuu
XuIQvnjRdv7AhYV7PNHo6sq9Dz9p57LybkpkO2ocKg8fXeIoHxp+meZRXMoLcAnSlYYdnHEsAfJA
3D5gDHOKwgZI2A11um5Te/FSlZe8eL5TXJuBPLugr8whyngVawStaKtxYuvB7Rgs6MJfInWgBsl4
yMnhqvb+uVQBXFECVYfD+PzLqkBEUPeF6k9Al+QyuCZOJlAJl0UozttysiJLmUX+lYvSpPKPlOR4
KIoBh7FWKSfEp+lppwbc6Qr70Kz4NBKpRa1TiuHzBMGxpJhvwwfOwgkfMFFoOWxUs4YcEEklpbxG
/9gQnHhsxHiZwt4k6Zb1gSrFRnpuMdzsJDddHomgP6vfl8DT9gV1avqq18+L75sz3fVh/lHZXxN8
OBdVKwsfvujPMxNSi/rhyb8jzPBjhkJaH1c9zGHmYJaOXBAFxOu+qZctxnnrV2bMsopvqyPy8TvL
KojErFrrOPapADXdceT/66KXkLMS0lJONVEwYIigUBTF+5XIfuKSRZxEVR3G0S7gg8X0dsjpR3O6
FxNopgkee6aCLGLqvo6TPJej+437D6nNR0+BykVBaXyAW7c8LeV81Nuff9UWFRX3W/H6UpELbrHP
+liDNszJZcsp8zyWKYOpO2XWgUvGifrYTPjwSxP+t/UXyJvvnrd0Ikmm85iP0LWGxTKlSx8cGI4/
N2KFhXs7Iz7pr0WebCf7eTXF85mjFVRlsmNWjubswvCE7TWIqgoePrPhX6NCUEHPj7YHOWN8GqmO
UGxMRH3kigZyIAa1I2G1JwKyfyphp77zXRBr4KW+O1HY1c+EB575lAP34NGEbZckesppzewZVOpQ
fdCcXWav2Z2MYvn6IeNRQ9LhMRX8PkwiC1ijjpDxfNRY74ibQHLBhw3w4g68ImGMoOvq/to5eXK+
tM/xXHr8ElKDwplnMlMMJ3rOkt0T6V3j/U2rHhvIyRMUBiYo/P21pUZsdQKbUc44aCsrm+S5LPRs
OJ22mOxBXTD9IyomCLc9PVPKD4P7M59282I+ik8IoAAWkP34OcqmVF+QLPtJKG+xmlX68l8M9hKH
cqBDHQA3pGAhHZttyIa9BLng3eydvh9pTNMd7a7AzRUZufz/I3r9yK9XTHnGY6h61tEu0ufJ11Ri
x5+2G1J9eA6wCtzFobn0MtTzlhTmmuK0zmUO4Pn775Aslp3pOayLsIS8+RKxwS097mEraPOJjKcz
i3hPU+xTAMZtCGyrd30uADrq3KhnOrZsDVAJITLk8GW+hE0iGvRWCi3GMXsa+jFH0lslF7biE4YO
WRTRSM6uiJ7uHJdkPPR3EkBl/eq3wczQU5sSXoH6wbx3YfI6PMHe0IDHxU8XfYdiJrKdDwulHbAI
DBIAFQzb9OPi9kmU+B+7HdME6EyEgEUR7XloswImLAOVLw5j7IfcGlSvH91YEX0zoLoPcLAQq/Lm
P7yuvJcVSgSBDhyTHhCil6AzGAs238IjusVnHzifciPJwlb8to3I0zmirxlcB3upCKQa71rRU3kn
K0Jw/E/M/ewxJPswoaYvN+GjQFFuRYkl1uKmmYKLogQoq8w0NV97Kg8RXL3glEN18SeJxIAy5/HW
AEDykvmFmmSuTrCGNqXPILBmjBBHMxwnjnwWzEoyyCj3EdewAt5AI5mMo/8d+OB0S09/Fna/lH/6
CA17ednzoLy0Y7SYANO9wTTqEV50F6Psjk+YHPa5fxk4bCJr1P5M35Ewg3U31XBTQhGRdaqK6LpJ
9k8xVrGMXJy9q5F5RtRJuRvuwiePjKnoTyVCgFU692lTjDEaMp3Aidsnu78scyut2MZe4WjB6b/I
bkxRizV+UMvxI/cuPl1eie9uysJ0w5yyTpkAgVhan+knSWMrVwQhTaoVl1mI0owSg0NyzsynXvEi
I7ZKPjosNO3UFv4I8kGSjELPx42hwC7hd6FykFnoymOExd7ySYSC6T0eAS8oomjknMfYvqbwgJVC
53dRB6sSWdXmuX+EGq+cJZ/06jCfGVx3YPsseT+VKKhkxszXGwgzKe4cbt8w60zumxkM+o5oBg4J
Nw1kp33bzLYa2VgJIxwUy1aPy/tf/BDZkz+R4m4D/C1ddBiO+sh721ooHqTbQTMp5ehtDZe6xjei
16k91HrpsAKBa5oz+xBQulfF0oP90vHR8kgtDhZ/Z4oqXUZzJrxQ/yFV3tXNa0QnjTmwXr804J1Q
QM7Tk9+CS+WhNNRSyfh2SSLjaw2DlMv+qHhQ7hforp0zCMOe5Ps9Yzk+f/DWOIF/+gE7FQFdIzjw
ZXV622CL1iAHtsR74Pv7udEBM4is3/zVCcgAVd0hvNMrknQL2EO60zmcxUe7tc5oq59PGWnNwucF
miuS3CYeEnjtTwlZw0VC74AxhcZfuQ+zkd2LCLPqXfnYjrwmjC+ktEwvln75E4uHk0Qwh06IodZJ
+r4TLPcWXExi0egE2PIXyHxUTb5HCW1ilFjEzQ6Ss9WVMCGOpzJ2iZN+IfHCJRuy3FSHmoh5Tcae
0mDJlOOS4dDenuj5gPkhkL9rL95srRnu5Uf4zXDUPt0NDCP94r94sMj9iiNk+1zdRQmysbwifmIp
6JXz9kcMJGhOB2WcHWDYyCbBWt6RbE5Q53g5lbXS8f+cuK0mo7jEvm/H4WVoDMa+X9p8HCRGEOfU
nbUfY3Q6GeLSszDUmF5JfHKqUTzTtstN5Lg4QJGAKwUOicapXSXOQa1vploqaOj5Gpf4YfVMLrSa
2oZu93oqjqpaYsAouOXM/ApcLl3oCxvXWYbEK43QeBl7vHox+kH2jtg2GsdMWoKASiTQWYme9G1B
aG5vdTyWOx+opB+LR6e1Ey4aCjSmYkpAPrc467ZFFzZTniZbu5J60CFkfQ1NKefC31q7HoM8A1Wk
GaNbmk4KRWp22yKcYk71UeHCHTn9SV2/hKpikMILW++Ww0DWWLxEzDOYrp2SLJkvlz5tcAhqKlVu
MKfl5TTxfkFvX6J/ejMCMaJklTRaCxURk3JFKpkIu80Zj0QsW9C9A0CdEhVz1UGa2lW6arZuWZC4
JFeUlGbXmcdlzufZGPKF93qhz7g+ZSSd+pvz4ZoHqsNAl0yRG4MNUyp5pukw7T9hbT7rZLL46u6P
uhOdgXlhZQSyFgmTFXtFKr6DjI/8fEPuO3rYH/dKfuEP8gqQ0hBMjtI9sVYJ6GZzuXWIYOk24D/b
EOhic132+5Vr5qva0ixw2e+WnZrEAdeRCCGFvbrTlIH3SFUwIj79m05OlHFKNaE3DGT1hxaQqPIu
s0HP8bE4fMHDhWTXDg1s14RXvOJVUG7uPkP1Op+mOJAjh8nNXSkU0pGNO6NlhnI8MulxdgDp06lT
V6cRrhzUct+ms/QGnaBFlwCqtXBK0cCB3hsOrrEoYHmUxlc8rMCKhRifA1sOF2+ALYR6iUXy4D8h
oWBsXlNqhZFO3VgLFEi7nxTvIB3Mh8+7aIak9Ux+xjUuGl7L3e5mYHAFsbgzpx7QTQCyDZ5saiQO
sv1Jh4jYiPsJq92k24VyelpBQQOclm+qE28wnqSBIqf8MIJbObW+hGppnLsh5WNnlJ9YhAQ42hSD
2eGey2FNqUoVxq+ficwTmeXIgythn860bH/4IZReC1S1CbkI7c8R2A8EWSGchAWgq4hnZqBEtN54
nRa/L5Mj2dzOSCFxwgeOIzunWT62EInAvJ2OGtDjGgeoY+wHnwvXDsUX6p/CKxHlrk5+TPNGELHc
bylmHup5HhOBanE7LlDzjLQHJulBuYr/SBQpzLjEpj7Zjm2BjGHb/dH8WXZ7zzaEvum6RIOFDPog
8Vchq/UpfAbDQqLDAj19lr0Uem3O+flyxHGaoW2boKkuN8EsXLtFFtIXoNgKQqDZe33S3twud3vO
tqobxWhCjnhFQ4X2SCiL+eQ7oX3CYcPTVRTBgLtvkwfTis1romlJ5pLePeskw0sk8uUzMLYSibO9
l/OprFqzZULwod12hRrooNxtj5e1uVj/qoWKGcjNI93Rzd+cnjs2RvAiIDNH2eimt5L1s1gxo7xf
jVnV1fkCReDWJSR9mu0i5qhq8cQOLJAV48Nx/CBdBOl2UnR/tMrlltytIv5AAj2u0xB2RS5jd/Vo
/75/9lwokM5fbS/Eke+sRjpMvR9YiZPF+uYMyuXr+gYM8jH2O7vM0lnglrAgXMYZ5/6jLdqpJ7rB
+McjsRNeLucC0sH+orB7AFuxApPqjBpE1p5qPRgxqJIh952JRPto3hmwuvlSk0e/GhsMAsJ+cNDz
daLOd8QeRSXbHy5uwZPNI+zcwYFUAtKvlxKritnU/dtlg85CuaZTTLSvPyrljwRJPDXTd1Pz7hhu
y82Lvx7W3AmJPCnTEwnRlHVIrE3HcHbPPV0fxOUgJLc1PZWppOjdeQ6FXH2vwsjOGWQ4hM5+Cchi
wpVDuaJvwPXauBJQjdU98UFf+u0oKg7M1Ml6/DeaErljx1JUKY27e8KPuVADfd9EBHueF5DEmgQy
cbC4ssJZFCdG0+GR7hbqMOTFZkmq7PwlWJcri2JQeyqfoV/q3i80/S+QDy7uaDn2uTUmZ4FicBZq
Y/eXzHFGg3jH9k+n+/fYMlSakLUg/RBOTyJ3ryQXmfIs/836NHgyYMUG88qDJHzwDvjpikVbX14b
WhZQTF5iqi4PjevoVEtmkPAQbBMeX8fzUNLr8J1QrucEdopoYDwVSZeHZ60uhrwZ8CLSb8j05W4c
H7mKcwjEBXEKGAQKl8Bs9RagFixJJDRgIzhGNT8c4vnjL0Nyr6sRHnAlqOJB7bPeDgPeXu2oj3vz
mOqGty0cuIUgYRlX4hnX+pBmtRn1LWWJiFXcXs+ynIkMJurBodVQH/C+CiCpeG1v/WihDZyZV9YC
VXwzYj5qPpYqvJ7iqb6aVFiNo7cGlha2Z6cUVVMXZsvwf00fhxGfWCzshE+R/a8fd0oQLwVfb0Zv
ok/f0r2sMpKipkkFxfUfnw9Wn3AWGZrPq0WNqgS7VolKEunz9roEd5l2pX0t0b2LRp+zWHeK5g1W
DFhUalLAnSTWBoFJud6U+JFztqrTymTqsssPA5blQVSLxwwgqMxGkSgIaVknL+tg0GFXywHi33zT
F7VFDLkvaailYr7wVT70dzIQ8DMGzTT6Vsag193FTZCz/ND0a1N845mlebEAUI9CjKsFW/l2qvVc
mYQn9yj90mA8btin8BxRYWoVbf9BxIL7nSTwP6Q9Onyl40tJMu/+S2Csncy2/b4xlxtKaHOj/sAU
JjJih9gmPu3WKnYwoRSjV6wtM7o5AAwwkECMsXBXsMibBzT2vjGzZ0xsaxD8xihVAeJtixqbHHbQ
YNgmTjSavvX7sgp3Du6LvHZkYtF5R7cuxD7IYCsMT8+xu94iim0HQzN3pkaWDWlYdXACA3apv/hP
wfTOmSVXREdxfAOyAylGyT/NpOR3eTSUQzt62BPQJV2c6zzbNz8ZXWBBs8MABFMhXP5GAla3JZ/p
0GJ9L2Vvpb8ZaPiA/IQGObzMPcSZg/pyvPGjVBUE5Zcr0rgxzT5x7/1eJ1sxGhxjrHc6Q883Fl/s
QHswyx1KZ3hm7Ro2IF/xHvEfOLAMWHCciyDeof2z46HxMNbKFBxPAYdoyswFvB5rTZ/3Q7BSgGTl
KFoRiKGTzD822vGUMNDpsN/Z27DpURECYv7BVhWriO882EqMZzANxHgLkoSTVDnLKOiTEQ65esup
IShz2E+Iww1VLBSjcM4msRQqTgN35JtmPjUqV2GbCnU0J0HPdpyp9KMukJh5ABc1fcnYHa+vLf2k
w9anwVgBN65xUjntcCy4nk6nO3A4zH852dbJoJsqydj3iU2YcN8UwquGMCEOzauIhLIty/iNcTcQ
X8+kDagMH+DT5zIJn3NXdf/gqvW9FgjZeWSCsJGvw4JQsgEbQiVgwIh9FBB0WxFA9BRGm+F1si0W
DBR/2Yyvhab9cws4Xn2VkF0alSvf8Skk0GqtWpyyCrW/PF1xgAC7JPlyZRwhJ0IHQYWQaW/+p2Wz
A/+iKUImw7+js3cmjrgjZbrcLVEMqjthpaLrPlbUdbA75sZ38kJi2D7S1yEC+EkpidHhDWJpGaWC
Z60itpw1vjN8Rv/hUOPRhRxXCslhh3AAIRvalo+XthLaGIrRHIXBBF6HD0+X/ob2J2vH52wX/tBd
3sPSnk9v912fqj99SMzq2vdDjUUcC/ivve27V2g02edcBWPdi//f4oJOd0ouAj04aPDxpmIxayLd
bgjBhwqB9jQ08H28uCQDU7OWSRijFzNCwF4kFV8UHAG2VXVDkQFCxxLA1GR9wlWO1RBrg10YAkeM
kRxBgUHOOmM+eJKoVHwAvWu/hwLuUzeA82IMtVtwaGhnZ1jreYWGTpDCq9+umyK+dwpdM+NEfV8W
eBZdXdD26Y/agkYSTIMf/QgzmodYOLuyeS9XAGRSLyfx972J4oc/BtGGRG/bEnyDw4O4wZBXhQO+
s1iWO3DJ+rF/irEaqu2lRPToruD78v3bMXMccSBEmTaOQQtMBVyReFbdIOKyuVpQyjqCSZfxBe0F
IsEnZedFrtBbAzpPb3K9vG9jAoltcfzZgxP8lIb+nrufiC9nVWNk7E50SAbBQNm16vm5SyQAR0DE
VDAJZUILRo6pg9Rblh967tx4nJqow4yGT7xO7kcYm5P7NjIi0ApM5L+cukWetEk1NDdjj/HOJRR8
nabUEIT+oCb4A8sP5RVlQxTYKDiSKvwAIqpPOvms29VtKaxdO9fmcyF3203QbGiMJWYHkm6Jqd2W
gXuVIXvQZcf17JRQ3WLfwZF81vWECTK7/DNAqS9ZZoITjtnPVxBtzWrKRAlil7/mINjETEq9W2D5
g32H9AArY/6Tq2yGaEuZQ43E1bNNVZzzRvk4zZht2pxBFHvWdJ7MvBpoazLEh1CmqIBjM6gjAYlX
nfsCPc4pf1iAQGlVPVFeGh7BKgNrc7EBiRsPiqLPGmCDM6MQB+pDiO4b+f/4tyrxEkvHxDgoJWk9
SChETtx/bBk3pMC0i26uYI93QyvUHo+yjO2pS3xR4HoTS3ctMZDjET+O9JWtl3ONdbSzbDskB+aR
HN5zdhvorIUlC2m9FMelZAtgyRb4/vp9PggYSh4eWM4vz72riXD3m2PKA+J65AnP1cENGZLdqLVI
K+EbWuY0lyzIpmVjMVZbdGd2wFkqs0qLwSZqD88JBLH9R6NMcqJajtp1hFutcczqij8KYJ0cRMnS
Wdco0F7I/x5F63217uoyk2xR2xZFBTusD9NxE5oVoiDjsMh7D0t+joZGcog7k8acE9MrPQn0tQoG
7gCy4WlT3Kr8HeMLehqMskvf7dE7ep0B6EwkKfJqeYMImdp9M4kF0YbP5BwSpufMm408Dl3IWg61
amSU0ZGonEXZ/riZX0GDdRyzT48XgBbwRudkd7z4xExJSpQ8r0Hy+ywgcOWMYp3+0DQ75pu85Q/J
nwv8bWdAcNe+XcyyJpnHVPgI/AlOrt66dOCQq6eYbiMySpunY6u7A5nq1IJKBfNYdWdvJS6z5PVR
l9tqVfz3cC170+fwh4LM2PWmAOeQRq1zhkkBulsXGiArpB+9jmGzd+4WT3pqIcOXFEp5AMQBgxl6
ATNWKx+DLon3nQ/F6PMtfbYfTRE874uHSrgkGJoYPOlQNqvJ4JXiRL/CJfiGl9cA7IRqyfKgdSvP
7oTuYtVpvdQ/wv7SiHPON4il++9zaNl18u+Km4NRV3nF/2GbfkeUZtV+Kg6ckQKzQ7oH8Hmvl1FS
dGY6R5dh14RPVIcIEdkoM2AA0QlCVIBQrjaWsDBCfSUx2v5kf8qnmPrB705m1EQ4WkdmNZEqXFiC
OoTNPh5rSIgAgY2ASHVxdxDm7zKJM5aEef78j+9qhfDkTvr6mhovGwdKejU8NU7Kma8JENDeICrm
qu5zFcTYwo1wLjPZwoK4iNTRS2dCEeHfOSUDPLOZnvTQviq+JETwyvmakqDUI5742EASaYxvPn+t
7cpZNmRB6ZvR/g8xCNroYePS6G2FlsRVqZ46pRZ2oaYZeaTZdDSuF0SLkG0jDEuukoh28M8FARdX
MGksYjWVG3E2C5LMMUCZdJ0WlBneUFHHwgbiGtwpmIhqes9Jv43H/H1YKBtU9F/8MWL5KJHv34VL
d94VOBmWNuawEj9PXWIUoEhZz3wO7vbP9YPT6O6aVsajX85/Z5CBfTKGArNr55EPoDHQp9oebFUV
AailW+bP7z8kAYWRgaT+YTfWdNd2kaigg1mPyJpmjGbzQOknmiksvhxh+cNuSX+WJXiH+O2w7KVM
oIfVnGffVXbCxMFsZ0cm9V20zfaZRhROmdWT5TNU7z3H0SumcYwubbcpCPWKM59czq9U1CfSlj91
5S2PtiwJNJO941beyZ6Buue5SsaTFTml599m4zbOdcTQo08MLNKnpC6AOgNeNnyh0y8Vvo8ErOcF
J17vnIB3EZcAgxHTt/OkvdyVcA5g5zhP3WqdDlD8qUL/vl89LyuledjkWNznJVRqnHaAtEmVOxq4
xiSiBCdlfp/QkXXTEkoUSd1PI2rlwaRTLWofF0l5TqHcOiqPCoV4PVpeAtd6x2uN+vGcVL7KB0Sg
lJIZNekk0SanUR3jWhwEpzqmGmdDsuprbOIU7D8Rtrn/0bg9cLOkUJ34gnCDhK8PG4r4+g+Xj3lt
YP81LJJGXZPn3ja8/wBNQgIV4q/a4FAvsY5/lXy+Vh7n8j8k6Nh07X8G7OrCy1h11tLbXkiS40U/
62Yta6/I78a/2wyLhXN2axj3if/ul30Pk7t/Sp+YMkN5EVe6hSmrcjTWS67/9mwPVTz1kBTRaFAB
5XpEPxNyoUrZaeR+ogTQSlUeggHsnLzT0vxY1SYOk8CJowRU/stdNt3+HJ2Fnc8V/0fL0FwbLd/j
6S5T8R/gBVpZrUvEyfTC/isOMtmvuQzdKsIqgEV/5Vr+mYkZRYEO0M28a/+4VQGT7xy8isovci9C
sPBwMRdEJ1XdsGczy99bQ1Q+EbjOwHvjw6ulkYAmYru/LrNX9BbK3POYGlFC++vkZyeXsFdkwkVf
bZ2KSvjhjzFLjr/TnLAYVXlx968S2soQvWyHQQElBK3Wc75WgddkuICst9zbNnMOXAlRVjJag0ss
epjUJyeMvJR0ZF0aq8tNg4Y3ZUA4YE/jWodVDg+tN6W08gFdalQX/2lHk9Ox9Q/mAeYKLHlM/aOm
GXI0qnS6ywt2yQigN7atE4lcwLa1HunjJA/C317gTCacKSF5ll9sTv2ZFKIXrJ0CbVHKgTGAQfpe
rL1gDhqYyEDZJu9XVS6aFn6rjPQcqmkgcASS7iXf0hb0EwKKTAYs9kYPQjuM2PcdLZKM2uBfOnA+
QASTlaHiuFsEYUfZff1Bf78Gq/Ti7WLNQpcoVrts9YGyVpoGuRYrQan3ElimloA1oATGzlb84K9l
X8JZ9UpienaOGWivm8NkgLjPnygS4DoiVRb8rLF1ilgRWkL+GPuDwwr1aNi/e05qr/5rWkJ7N9gd
JN0au0/Eeb22O2E0L2esG5MI7LK09vEVsHpaXVpQ0fddgGDN13jH3w2P00oLzMYdI89L72zmPLKc
3kaHNnalt0IjeYZdNTaMVrZnumTQb8RDa+Pb7dFXyru+w4e9CnkwcCL/j/uQOBVQNVtICjlxY3Kj
u9DurGYFpkSZ2a4eTOagjsT61eH+aLKjtDcNPr/gzuNOc9XJdEBw1yRWo2Du5xAZl/+HWPD03JsY
xliV13rw/ev/5vbCJuRW9e0JxzYfET+umH4l5WN4Qj4x+9YrCifdG5VcvFlb4yudcBG0JY9ZXcsp
xuKuTcdhsgC0O1/j8qP507L3J4vpOju3x0sTvBjPCAWqHI9Oynle43jT/8N2FSwQdsN36lp+31QV
m0NqdpXpUNP0TRLL0FSthjTpXaMhTFO2zOyyaLXFPpL/ThkZ3NHb1VvXfuVjtrGpKdZTFX434rI2
RKtozAnms/n5l25CT9yj2tp4eG3yFt0BLW6UNLLlC7DxuAAx7peu+2jBp4aMWl4ZP99lPwM/ZSWl
zwnR+6DjSMRzMYw6fi9i5C2LJoWeUUftaOZ4N9W/49MFQCGAOfJwjqp+dDwaYnyZWqwbHACdXBrx
4N1zLAT7kNbD9c5Gvuqu1xW6u6llXuMaK3ZelByzX9T/JlPjsR+1Tocg8CyDkRinM27qKEoYLbAk
rtffaqd4CwSuVgUhQ4fKdrQ6D0ISYknwUOE53Bxa5Je6v9/nKZRmE1/BlCSs0IJb4LDJw6EPwLWQ
o/CMnsDy/bteIyy1Zj/5fiKgz3VgglY3qYPDt0vA2GadA5jxETTVoPPhMuDdEjgdzxP8CcnyhCNf
DgBESidn130EAEYNBpiRsSmUIgYynk8rvQzJqk/QNQiwPc4mxNGzFk6JwLzyLKoL3LcguUi1gnql
+Wrx7b9aKFG3DO0IEBJGB518m1PHCQxh5QY6KwN3of8NcL9TTLD2lbUey4jcm3EFUh2cs3hrXxBO
XlKm9a1iU9s3StMYDTwKowdh2ZsgXmYBffmPEQXKM+eWriO/PrHhj+eX+J8fA6mt+ldaS4Xq4tBj
uWkvyb6tJvpaJrqVD4AjHUsLrNdh8S9VhgaOzufmBGF4YiJ0defz+bty0PBxSmaX3L594i1/O78e
CYc+mC7l7PLloOMIEtoJV6cdgZEP3rS3RkrIU/H72EcwWAYblM+mMTrdXdxpugUHoQECaz4HH1Im
XbViYsuxuVQWKQPynkZ2L3zDfG7VhCwxfBN/y1d/ebqxlVn5I0eaLmZ8zJbI81WU2K4iuhrWOiWw
imnMl8Bl7/KYIckK7frwf0ox7/X2M9Q1xYWRwImbJU3wUKqmNNJCpNgMQ0NpYkvdDvLBRe5C4edJ
XUCLufRPJRTbenT2cRzBmy8gq8sa6IN3fb1Q2f6N1IOKaMC6W90StWczB+7tHJk3Yitvhvy/bXr6
TrOF59AbDGohBvNQ6Rli/0cSZGk8vQnS/CLyl7/QY0Md6i+RNN0mPCxnhkt5NFyW7cpiWMpZbzg7
G7huXs9PSvSlDYHHJhHvoQmgEB9nn8b0JdCAaYdBW4w1WL1bLoUO6gYERWqu7qzRoBgPs1954hO2
eqF98/uNZQmbIrMH7MExlbymLjls+f/ITu3w8B2yTwaRm8H5e1Y5tNR9roVYPrnxoyk7bvusXSBo
JeiubPTQLtr1gGmQ9Hma8eIhYGaI1Oyqb6Ra/YTxh3CgMjv7lmZ4kFmmNzLhADAP2rh3tlX7vqF8
b7KoOXYHyxsJME5c8qe9zr1eAv56X9uGrrp4sD1cztp34eoV7umriQhlRBeMYz/Z8zGJ2/5JPwqR
lxyjiXFoJo6Blq43Ur4FNj2CKu5uILg0yHKGZNq3Wb5UnHqzeCHetCgWtI+UElHCykh5KBbSciB2
UZq2Ku4zn4crrSnQKMv2pHxiscKD0JMSyFoJfmdKpTuq5/2/tc4IvIxwSTbmJwPyBzo/6pxxalBc
12OPZIqKSjnHwGma/qnDUFmITk+m7LL/KS9H+o1DjyNLNWM5w+MK/tF5A0USr+/aG3MivauZDV3f
dWTC+i6hGPx8qkVkDwTz8reUdKrhSwF80IOf9blKJu5nJogzRjC6MVO8xjhZIuGflbSX+3MV1lOf
V+dzigq9BGayZlTmQrtqZmBYaoe8L46RsrBXFcCpfJdb6YPodp7xiVSU/9iDc3Glemm/MQbOwLkA
hRpEU/ljxvkfA9L2JbtcfKr5V4KuJqt63Lyx6TJYJmCMpIWO06BWbAPkHKWv4jsDfOffuuDR2t/q
u+CJN+8FbksiLijPm+SM2D1WNdyxZHGZIJQ1c8lH7G9ebFfaHahjBh+bfhWAV3+FKYDGcv6oFk/U
VJz3m4dcXWK8ilS/M3mn+7emCvSECPVaIgWNfipV5tt4FxJrZARxOiA3CB+kO0Xi0qmvCZgiCP7j
qo6P7YxYFuqIEj1mHIh6x8Fz5yxdJViCggt4jorSqLzER/BplyoaPff/g1lv1wGziwXMmR0tTbA9
7QtJFZDCpUcQeK8p7YS/ZYLZCJelgvVUtRuekB7ANPteOPirUfN9lDwpmG2QXQGn1SatxZyKjhcV
XiRG7tpN9o1E5d18OM5NZ05e2P6sdGDW/AAnXjV1UzmpV8Wfq2fPKzTOaTypqUnUvAbSGY337uNk
U2Voy33nRo0YjgFRONrGWlUu8rUaJi5Ulux3Oqh/XSlG3QYlX8Uuwyfo4CCUDMQoqtD7mmTF2Y4L
SlAtNN0EodTV4nMvjOm8UxdynzbHj8Zs1EOMeW8PtqXzkOHDtdfkuW+xWU7uHVow3XuQesm7ThKz
1xyEkL1ztNK3kUJGlc2GkjYIXmq/fM+A2aU/QPf+6zvJtTBXSl0KQwbvsqa6kdHjtmaDubID2O9j
7nnl39+gcmviRufOhklHtmqBqcATLaHiVJkzIwIH8q3rwlhXxCguBkYA4bTA1S4brdwQcvLoq9/t
TgD/QnXpPralOrxpX4NzOhWM66LgbbHCxBfMs2wjYgH/qpoa7QU3AFOVhvxqfsEFg1Pho8FXb2fJ
Yo6D5KjpL3EA6EQAlmW58UK2nNwuTPTcB9lgqF3zMZhD45X9sGvO60jeYgLmUMxXPG+8laBmjIdn
J0drx9Cj8A633NhEf1fEreYA24R0KqwmQgFnXH06UygIC7TOSwsIuSE7rH0r3JwsvLLXQz64javD
ZM25iP2MWIuz1mW1Rtvfn/HoPCLG/9Svm7R6VQMDaEhY5xio3Gq6vlXiknDdPH2hAiPVS8mIZ9x2
K2RlSzi9TKrIxmYK5XM9PM26iQauYZHFA6eQOb7PQx4sCtml+8xbNzSfbYf1qHJguwc1jZFqAmMQ
JrOpP3yF5vF0JbHb5pWwsuHYrl7d3yxKmGVZKrUh+wcOovQnECEyZuWUPEmcFyrEH3pQuT6Aa6Xe
++POGdUlD7gSsTWnJ6fKVzckCDd4TV2g/9gVqrVSC5HrMVeLnwy2+L36/9KuKcnNLQVt6QV7WidQ
uWpB1Jdz8vYmWZ2C0TExpmibxBHZqP7Qctl9ePtUoYqW3MpjzCgULmjYZpyUAot6W+7kB/Ag1IXO
iXoWDSS55lEBEfjd3ZC7ZVcaky8rjlidXcY/vIJEuaLMSuWidz0zsJEK1ZuKSozSUx2bCEzsAeke
+QoLNgHk79C6SvWy059us60bv+wADvitLXR83L4IMccFTPvcoEWRaF0vYgbdeImfCqFb+C9EK0Vm
+2qtpPgb5kOH6EO0SrLWQz3Wmql7IU7EOmYDE6nq3J7oPHcPyyg/6zSdQiuRcWvOWN+VVMxR9KsF
Ew+Ji9yonwsmH8fpb5CXIbk0UxKef72bvQvKrgce6IS+w5/zSTDved4+ZP0N40rXoEXr0ioN4Y8j
B9u+HD+ZPJjTDZ64Mp0qM9M0L+hfyYwFD0BZWDHMtGg1+WZIvY/wpOC16uCi5Hedl+UoIQJrhrBz
K6c4kK8QwAbgYYv7s6Kp67NSzt44ArmP2xQl+4PzLCiI7F68EDI4ihPWljG/67EaGTtrhVZJig64
BD7F7hxS/6qwmYhjz2l+jxJwhORtTPqb2f5EHWp9oSjk3kADPa4p0VP23AEhjLINjT1zg0K2a6Mx
8WRBz1BB8ctndifjW+lcYq2RLbhcaHwmtSSH8LatexB74zS8sddYtBSMl3++5Fbn1zToVPYZ7oP3
UP9KgpI7luAbVkI79AQtaQDz5C8LZ5wOYP+wih6oaxn+Ce0fkfTwoPJPWoQVTloANIuxlKfoHW5d
sME5s8qr4TGnX/GDss0XhLZOM/4n6Ik7+gtMLvMq14gUFYRwhu1qcg2ue5DDRFv/omhQomVwv9QX
FBcJ+jHIYJLo7gi4gvmj1Ui5hgwrqXqAlVPmMvV4JX+MuhJ+oQZ1xtvLxabRazB3iqQjjH6LliS+
2ZvRY1L8Xu0bTH/TRGKh+ZYMGTOXoLpWqB6TsHbePdMRnj8FwmX9+IErFb6293VOafxp9AzAughz
9/BR4mFpOH8SV4JS06vNukKW3TAZ3BvUwxL5yfspVBAFNbvK1qJ63rFf8Zr1SQ+5sRg0go7n1a7v
yxqL9rkHE8ULfazWyaWsJE/MeJLR/NqSZg+ZldBn176aLDRXE/ptDIF5MFQ3QrZ6JsZqfcFO6YZs
C8sDVNPBYdW5gCxZ/q9NmyoVef3fX5ZM33pevWOgfoJiVA3RDRBHea+GvT/XQG4YVK3CvsOyVfIG
S7aMKGZUyxZ7hZwV5+asv8N+6FDB91GuLjIjqnxuRI184PdTu0FhoX7GqQP9A38VHH8ECDGX57uy
p/ARbrDTg7bhyCuvG6rt+CyAaIavSfyNM7QmTKLUsHihEMVDBaWedxPuMLVaMMACXRbKdSwk2ReM
C6ISDtgUaOzRE5uIjMRNOzozDi7qtLYi3EC++LTnJCMMnyd8LcoSYL5wXzfI5V3cm/gIUeO6w2WW
h/1Y8WCzXsR7JDhgTt8QvYk627CH+x0WsEpRm2dsE4P33RmInprOLHe50z/xGRPU1Tzec+G9KSCZ
47714vFat8FSY6pqNNohdTqLqG0XqHueuvL3n5MhN7wmGbl81HH3rLXZ2Ly7fraOItW4FmoS4TL5
3kAXE/1UDaG+EO6suuTV+hIdodc+1xJFu51ZoBIFZsmwatKBR6W0JpY+kPCvbvJnkjH+/ik9/TON
oIXciD3sMsQZq5PwvNNFxHtJkCG0cEQ+z8bi7bRWr/EP11z7Bs/lM8XHCXLJFjrA+eGOznfMGXRR
V12wUMzj7G1eQFVfxELyAE1fqpogl4PTKP/JDB85ja1tTaQhsQuAmDbTCNKhJ/joDl6kk7CXzrNr
CKPDn+vjG7+znqGZRSA/qgz3X8c5yPiiNpMTr0uLPIDXHnEiBvBg552t/RH3qr5+btJ24PTPSMOH
CMqwO6kmCwgC6s8pq+t9B+wNRBcWNrJT7BNTp9Lpe+RcwSEdB40rhebCeEYG1i6Kw8rs509jeY7W
c3J/N4+pdeI2HJDNRjc4MQWZGDcahXipyWhKmrDAbVXXEutfz9DOxrO2i5zhnEWGSRgB0jqLuk3V
8pNvG5XkWrGKJpMMdlbbKc6hNjwia67Qu8V5Ye2yb18kdbEFHDURtmT/5F1t2whc2q7+KrfPiSJM
G+IPWaHOn7Jf8vArYQRUxUAtJd5WJkbr3sSnSCaFHI2QQe0CHZ051HZcKEqms71r3ZYzK2y9PBB6
HAIRTyfw7Ms0HyWNEHOLVUk4FfH+D9b1RYlk1FUblChixOYwSCOJT6f8IxMFGPH/WqjuxWZwioL3
2k5Bg3BNKOlExrQS0ZfsEwuQgWRNdlxk7IWzOxdCIswuFNh5quVFotueEXHuOybKy/nG0pPYjTVr
vkB35hJ7kYB4nDWJVEEpWW1o0kTb/FhdiFEoS8OrjfBrR0an4SqLptXvQW4PDDYluKpqUQOfp+ZC
8P/NKHIgHYB0UQ5R2ZUj+ZavjqGLFCfjchEpvhEAPaEGLvCAae+qz5esEHRHqy6ndz3LnufPmav6
pm8iVM5INr7YawndRigzy7GmKW1wkp9Ixnq7RctAY7dvBWt4OgxdLn6UK0hix6tix0vY6SUrbU0P
aVdPyHSXzIYj6xN21q2Vdue5hQ+g0f+UlIN9hBRxe7bArBvjd0PClpeC0I3wEIXJ72kl7+yBKLxt
XPeajV064sLShGtYxxHJwjd3e6QepWatPQmmGXITT0K6OfDQqxi75KWyGjTTnxwGO43QngNZYTyu
fXHrZN2MDN3/U36Ri0XdGtCcbhJ2I2RWldLumM/aRk+mEE1QB4Ge9IiQZMC81OuaT7ABXExLEVax
4iw1+P32yh0wEmb9nBNoPlJ3D8oINulIwzUAlXTy3DRxaQ3zKtT2xx0jkZnXp3XZmccmkfJHe5Az
O+KuBMrY3x06YSejq/Up1VxAxwUbZSkBng7tO3EYe/fWerhFCt3mZ2YjzrXSIiEmZvzYdZE1VrgI
7tZn0jRIJfKp4cbfZujP33xtcV0ak7u07rEAuPVPOjjExwwgKsvTUwtOdueov3qmzzLaBI/RuqWX
wK/RyqdYa39jNQYXgrYAv65nwSM0JGu0YRcpThzeOn9RhV/OmAsORSHsYGvJYyO+3PkBGQh8GDHB
ywljHNIbI7kcGH8s5lm/I7jAgq+jWO5Knko1kpBw516JIXBm04QaowRWOWDi1T3yzAiFPt2NnwIe
jCRSmLj4mWCWheEZEVdUByb9Zp7EBvyTsi1RVPH2AQ0u3BQfDE4JxrBchi0uVyZLnAKSQeYExD71
CqklLkfHf7c/1rdp8s2Kp9mLOtsc6u/zKgBLoT7gEFZYpMRwlLy5b6AR5ZP9SvBmtago/PAAifgk
beTJHwvMQvZd3kw2zta2ecvtn0nkbt7XEmppM9Sx22YjLSjbYsy8DdK1/uL1A/mKTakDuBNvge7y
7Oka97wS6/Bkc3X2xaJwCAbw0vNYh2WF39vCd9hqfeahsqxkwxq7eIouX5wMTbW+hgEN/DAQI7iZ
5L2gCL3NmJaDkgNDBzzN5gEWmOg8MnyHeBhNFhLzJsKHVsdehl7Gca3jzAYI38G2dFsc1CPfkNgN
elAIEQe1TN2j00k3XOZz6XO8eExX0mD4ATTQR6cACXM26e72zZjIZZi1AX48uUobSVlDR8FvWZN+
+OWeh/p76evBxb0fz1Nda63Y8UYOoVqZu3tiq9Z+ZYnKOgtIErdCMXGvxni5EZ/KS8CcB2Mx6HKI
zdj63QzR4zaEoPSv67GuR91HmQR+qxDJBzb7kFV+Q58RSyRyDftjFV44ER2uOmwd0JJOxWkUTS6L
3utLvejlUifxDd3E0WeyMS6McVDg3FWNIDRHaWyv/M0/Kj+8HmB2xzNvgi29UYLqEHzMJt7huHRF
1JQvEGcZuZqSKHqo6/cu433C1pYGDOyRm8sN5P/P5Ch/Yzm41Cp96nTs6ck1ZuDzVmiye+QStibW
wdn1auOf3bldLq7r5vDOnNYG9OFxc4vCWuDdwWLOfhUnTn+5pPM1ZzxxPs5NOCFBG1W40LaDpxul
zWtBJgxB5DznGlWc4Yyt+UywwR/5xYtxrfOAVvSdmJK5Gk5ygOq7/6gIJ1wTLzcVZxOuU/SsDRAa
Q2VzlBhx2wXiwVmPHTBXp9XgWlThJROFF7zgAh4UgHlUYyMd94prLRnkY34bvpDP5h9qRU89eFBk
6xAcscfDGBuhmF3rAO7ILXOPHm0aJmm/mvvO/0B3Ap7R3gRqmeuowlODH2bb0OhvYVjZdITMsALb
D5VUE7776sSd0idHMpRULffOYCvmGmgSeRjEuVwnJ6kb6/ejIQw+OnLjsj0AcoS0sc+g9VL8bbPo
hssnycW/FkQZ2l343zD9qjtdVUAE+Qg8SrHSjwn8drk9OkLvS7JSL26/mCO5fMNi7T236SqCJoSL
8zMJ7zDcd1HDdbFWjjwxLczZ+1SkIRwhLpwKCniKuM1ixa5BRxXBOI944cngrDUDN7Qh4+fEt/iX
oW6bcjtwRPeYpwRN8n99KnqTFTdnOWDBkhXxPmMs45Y90u8582swfCWkLTTv9hZeHiBIUpRgl7e5
UFfQ+vOcuFc9bMRGXWImyfDAyGwvkvFS+wxH/Yp6iUqDauFod/WPnM7p8T/9x/8TUkSxnJwyxRtz
7PqppsBwlKl7Wwt8jJYSt8zbgdkCgvh7mkm2uzbk6ZYFfffOzlZcjflWnaOm/ZpFfxReoAA/Crzg
o7PUuqOmm8TE0bJVrNX0eCM2IN17+Tc2RghzhzxawhTdYIN8U2tjMU5CLVLg0wWkrUUyjRGjjkvq
9Hm0YoPA5D0Gy0IRoV/GrEHzZbftkRDof/muYlvT3peq4qWIYi+pFe44njwyzlfp6P3xuMxZ5ykH
g4EUVSbHFlFfKyct1BFrWImZ4fPeJ6WLtsAT5REaap8iRND61nLviQkYdKfeDuFNO5lyYU5Sg2sV
yBduF0jkRYwoixI7DOpSI+3JkVr+230t9W8Dh9daEbB30T8SHSL0DeDmEBDtdnnuLRx1L9k9HDRc
k/xs/W1ntHxvsVq9aL8MdaZ+eQCLAwZcx5PbQSDU/xOdouCJ05EGprt6qRno/OY+pshgVAulhcTp
iP4+D2k0ZLr3nYERuP2y/Re4FxzqAeuJZyVzC3HoNJCCuQd8NodUcWzdzwe8qTBut887k6k4dXDb
EhfZfjiVeLZahQr9AEN8rYrrX6MHVXn+8AZU6F9ahlt5wvoFyc9xh8GYxFRWAt9PszOHwSTYXupy
oRu/qj6KuI+UBtNX+mUfOn37qNjfYRiz1tVXtk5VAxVATZhoEftBRWJm+DfC2zvE87bbst3JjGmA
bcm3b/JgweGXBIrWia+eFpL23U5FF2K9ofXm55q6fQIp9nqlS+yv4gyDK9CUDDyEBv4d2UBYGYpD
ZL4YaA1v75UKRkl+ePbB/DRgX20FUfMV71lP/I86U6wrE0GXmDGJS0r2nWEx/qxUElAwH/2d2wGt
7C+kHlvEngHnAbBaJw+UHNJJaOQPZHn+Uh5lCeOiQTAkDd6CkEOEFdNjR/mMX7qfChBTRP2A23qp
6A2nCXbMiS5EbE/3rNRgWqnIjgKFoU5RrCJ9e2sNcxIgmvmOD8RndWttRnQKco19AiF2V7gQs5Fh
iphVoHU8IQJZXCD5/Fd6NlnYMUEG+THiq5KW1gtxfPzKyPQ29mZ/2P9ietCrFm/9uDx7TAVSjAin
AkaT5V1eUPFY9mHPGTTiMvsZHVo0jFcHhU0eXpwuEFMMdRR+dApPlJ8U/0KXrzhItiyJ0i52bAab
TbnJgCHJVOjuowQz70CDa/b8dgacznswpXhW6+YyuitIN3xATa+9+pv87XTANtPoMj7xfgN6135g
9ElbP0gAQ2vuQYrAn7gUkDNj6on6IPkEbAMGR1bu4Cg6MRMfh/gLDGqrj5rhhHzQSFiXDtr9v4hr
Q9KiXzpfwL2dbRbnRiI8fn8lzyxv8TJN+tQ36P1tws0dkgKCZCuSSMrK0prK7KZdxKOoK2qBZvVJ
b0U8WPADNV0i/vosGNcjPD4eDgSF4JMIYur8CdsQ/Hx/ulfDe47MBNM26+DKj0AVsCQtNftmXBZc
VNjZv8Bm2aKjfOmqYpbimTbHhf6jYtfLmhHq+72mCmrsT+8e9r9WAQDKozawjoofcUrZ5TsOFy/G
zVJiNJLxpQ7Xec//sPko1w6UFmWd+IvhkBdV3KhA4Q0vcang+FjcxNB+0jLgPUvM5I1mgLqVr98k
R9sHD2qjVT3k9+LLBQ/i4Zua8SzKQTBW33IOJpZxILh3IudObZ4mr0zLtV7SAyQVkTBKwyZzHprA
HQBYD5zuo9vx+XBRX45PuIBR+NbaX9BjENgDCarw3XXNzMTDp6ikaGkHsQvMLlTqwbLVM1lAa511
4UEUtxIED6N/1WjDYROwAJPkWSPG3w9i4vfyq7AGevlUOAHtOKsbDXPtufaZP+ur9j2evgppk+VF
pRLsd8OXnocXYfO07Q2FCbcExvPCC2VrNIGf/1CwVOWiQCvMQp8Lk8tiEA0AOpNDS/pBxXOzYNYv
/NwhW/urF4rfDJXqvlI8xicgw0cTd1NIPJilHIcGBfOVp6BpE2cn6LRIg74rwcfqOQPT3Nzni5/B
6Adrjk7U+WqGOwYBx2IU0u+BFwkI3ctdtytCn2G/O7XcaKoPk2Nov5yc+FM6wPF6FZPXxNMpQ78C
ZjmlbCM5excxkmy8ibyCCeNAuu/dJ0tJMfvLBrEgoTe+KwV9VnwHhRn6n3sj+hhndd/NFUoZa3Y9
l65eE6CupMILiz/4N9l6a+9Ft4tNYjeDSswTVm/KMfQpwvajgLyzNYTDaFaSI9zsVuEgC6MMfY0B
hEQQXhq7yN0+PvL49ZdfS6GZLAlVHTsRGGvpJATOWSbY4E46Gf8Sb+syPaJcNNLVcMPE2SZpL66U
3Uw9bLCspJ9lrE485PR9FmpFGlGHFjxg9PAF1v5LMbXnRQ1kF7ADi71dkGh262bxQbyddV4DOWzV
vpTgeNBjLUlhvBGAI26zeseUO8wrtXVswc1hPCRdL5BVG0xTHIwI+VLyAo9LRAFeVEM8GLrkzVRV
3p/OcOY7xMacYt+HwjWzjlzGuLB1UNmbMxFvcHLDSd8l484tqZDHJyvjNZH+qc2b72V6gOrRXC8I
FqAZAfmXW9hmeU/QFC1FO5E3bwDJUaJP+uZd3Sdro4hRoxG51hfmBrVIxnBm71oHBJEfWqJ5Vz8C
SjNM/O1QiFcrkSeJpHDkPFk6swOJjbv9sL/AMOw6UCCsvKWlfJ0OCE0CrYyVtPiZnIZsKOjl4U8h
CMI92ln47OYtk+SVI+KJ40pAMAFthi4ztN+iTpzGEPp1gg82Pi9ApdFcbUm9XNGUex2PUEkGfhjI
uleOEOGS+OzrKrU6s6rxuLgIzyFQ/PbNab6PfDJHSByB07vsnMy3JAHnSstLJxY6rJ2/GVbCkRhj
i4TXZAJtwULcOtyRKkZmkmkthahkNwCfVnCmo8ExBZsBUoFTCPCoz8RluVoF2fM49TJ6dtK3Gu88
0guvoXT8YPTlw9UKLb1yMHquKhVUp/OH9S5FRJNSMbxYR/OTWhGIpBTVE4FvI2GpFlougmQV+9gK
/qoHrjtWre5lBWoVZPkfd1MSkHczJlARAGDVSUzP2sVQUAc4415mZewaUJvnsTiUkGakIy+BNjTO
swJyEE6KoJedBnIl06QvgaCd98JzKok56d6LjcSCDIXTua0u5kkj+pSHRGyFZPpteGfWBmIr84JS
aFqgEWBDfQaapQIh7oP/LAMroseBiLLwN1Iyn7s/kn9jwJN0wJEDfm2TS1DYAMSJsCzN3VKFnAU9
8eGiLxzE8G7MDwNF3IcNBymR7ApA7oDVFW5cGBbpJIJAUzYEP7rZJEG18KznINfZhjvqW0iklYOO
8lqxa1CqsokQFFuhgMfaa7G1yCIiPSph433x8Ef++66SlYU7r5U9PQg7M176aeaKICSPL85YFIvL
GNLdzOznvVQcpaS5RtYHedXOadWRMD1v3K4Ir2tmg2rPMaosEwTa3fhl1jx15inGVqrQBwy18FVs
WiVBGsOfgtwVprdnJnztZywVI1ux1GOBp8MvTZ7tLlSPWLU9nr4qlk/rSQTLr6AXRxZEeTgaslAg
hPSJiF2hqtjkI/bNTjLaE3b9UzBT+V2ZvF4ujwt6m4I1BtrYxNFmDcYk+QGFPg7p3CUulFWE9Qfu
xeo9UglwIUg1MllEblymSRSCOE5gZRXMPRlA33OkPnxWOKffJ/6ZOaC16L2rua7EfiX8mUzgfsJr
1ZqVER62J5hm4FSGKYljoTGlYfemAxhZk3gKtPLYstShADxdLXFPjrsj+zMw3EEhlP0bdIjSP38b
O1NKjBceYUj3qESy43Sej7FAyAoUYFiV7sZHtQ5cOTEI6tknoOM41uRwAWJ6ag2eTHcPig/gwY2a
mASVdHi1un8U80fuchz2XBEtwIJql5mcJiBhoj3GJJm9kHcXg9VG5ikfs0V35rc9r25xt62c6U5b
yKd+S/JYa5FvTKmeBoIR7NwPUgCJSpM0Lwa8UXcfKS1DiQtKfIgB6AaVpUEfwIf2R05UatoBvV8o
wGgrh/xF/4P2Tkr9N9S3QshjzsNRVrShe3ADbwXyhb+EOgBkb0klCk1Bnxll4ULFjJn/gc3VSOmV
riNSbk5+LASUbYM1NM3hpt57RgqBu+V3UY4C6Kg81xYdPFsVRHCCg7nQIxZDUXZhIL1KGPi0q71S
Z4D6WWZFbFPc1wxuDk8g9Zz+XPyaol+LV+rWQlxe7myn3FT7vBEOx/FYyNy2ITWuwqXZGFZ5s3R+
1DWs4pmusIXVZQjxTE4e8R8CuLGjWMZfBTTi5eX969tYB7+K276o0xxD+B/4KRsQv+M1LuJ2W5us
Gz3Bj8lQ01pMeiNSAcmGnr5+r4ccStL1EXY5qEfIm1rYKV6ghAub6edXI0+RjQoamPx5A1xK1h60
S1tzwJ45jv32X1SacWElk55og/2mDkn0isKRfkWpEDzKiABhCD8boOAaqZPvDZHtotPBKGHdNSPe
8hARv4Cidm7ON276SE2IC6MpxzhmwkihYmDWPFw9Mp/octvQ/8m1VAEjxaawsPXyG7JO9X35VEF4
df4IHGjLsMXObMeTNPJUIwsmvQCCIoxycbgC/msb1iN2YnP6uASx0IGy8lYNQgwVQhrWojt0iJUa
w/3Kya8FnOHuFa0Q/s3VZTcwC5lQU6OCEQfIKDHl/hEvgnv9cvFGr9l304eRZoM3rrCIBCWuIElV
ZMQQoraRt8FDSQWj/3fprmj61pfQZQuPqthpA4tIfyusI9H9HWtyJos2fbK+10YdqgBLzDWVPugb
hLTX7QK0F78wTvoUZifnXZNATDe+49CK8clkZP8pk5aDOiL4zZRexE4pKKekrA6/+nC6GvZ9BVpr
D3oSLVNW4VUyAjJpjopr5UyA3fYtacN7jvXO66xZWl7UuZWACCd2GEt1DVU9vAor9Sds8mbTl5El
xonn2ak29tYB09/5Kv30TuMKnJB0NfeLSMxRK26V5G/gv5lIg0n04i5SOw+HCzrAYrtOChLjnOhW
NllJjKcf6gkT2y1SQofllUcTgZlLchej7YaZgURWXq+IuApRZo+0KhGACeXT3K0HhIyhQ2pJp0+d
3kP4SqAuOf9cT6C14zIk2+mBkgEx+SvEWUtRX1JdE1oCXRj98kyVZLElge/rnp8gKgqlquB/jwZA
UKSS8OwBdqlg9P7rOk5OT3Eyxryz+vHHmRhIvFv3Na0cC8pyq4lShYG5RhH/J1VJ1VwYqGY+hjgI
HcFp5ASvSngjCw2Q6BdsinvFBAnuDQamHGFoRmqcHO/Wmrfoec9eMcwWJFnRuweIMEEl6GldTu4a
s553LvnlRbOZ4yQYhvNKJYzynHLiCkh4A/Yl7EHP5jt8usI8DRUGyTrJPWVYeIr852T7W8l+Pcpw
57QjRQ0FsNwdvicRYURnn+11CKg9Ra3B2xsPrKCLCz9Qj07yvxJmCbI4wyjtLD5jEHf8kj8kX36o
sFIAY5e0iZjMSduXcyWlgAEhtNlLaWYHFa24Eq9STQ3kc4TG37xe6pUOsCykT0vANLqYkALaceYf
xqf5sjYT1LhVqKkwB7MEAkVYMKirigth8TN860zfA68cnCksYaYTiyjzF/VV8op5fDMIcfn9LI7Z
z3qVb5L1DQDbIhTDKvU8Rg5CkLQ9XXEG+p4gvsKxSfI7FPT4Aiw9Sa3TbSujGdUcv8DQ3klTd2Dx
zvjPDieiJ9zsoTR5gFYyrkCvI8E+djmG1//s7qTO1GYWi8/+njDMEk97IsNh9GWOajLMYVxZkS9z
sHfPhIDiYp92A/ksmvcQpZVOgFYH3KBJZYRlbn6M1FW/LK2+eh7xIS9y8WxIoVmDAI5Yz8tUl1WE
VfQiLjmv75wOSLGvr2V8lGfMsDsmtiTbs6C5tZWPZjSAlvOr5uYOJ9AvO8o3murJ1WYiMjHaY0/N
t3O4BBbXfKU9ECBRcmdgD1Erq50UrV2aG1cLut15rvFKHMR+byWquOpDewLs4QoEKjpPfq0Rd4Gw
FQKfl/igqD59sSfUzD6+4lQ3KVoE+HjXu3E7urRY04ow0HbRBMy5oPI+Pir6Twd3kHX7hwdLQX49
sJMriA4O0lvwEtE1LiRc0qH9vlGhlQMAGwFVG7FX/+l8DAaxROOSSlrLykQWEWSW+IGclR7QXCrK
uuKinO8CM1VsESRDhWQRRUUR5Y7U5CuH+oAu9H4qX2xgnZH/iphjNlzw92iqTEBvdVkojjDs1wL6
x+KNMGGe0y2TE+1DQ14VJrHw9l8xX6nVC/FDfV3YFgS1vIfCi+mFQ6nIhYN7Q63ecBEemGWckD5N
K0X9KOW6qQZqLujQvBw+404ghS+JG6bAwKHYPvDSJFeLRlGLRAUPIWHQaFaCq6DmzoIm8dDAcTo/
QLYbCYMmsq/OWpOep9rBHO2XvXRZPfbxQWmD0F/YzEsD2DYYke+PIFla6Hn4v85BPTuvbbxzKtMC
z5SCDCU2qmAHkLy6WTPvZICu2oe0N0jycu7dWWV8BweJ3lDYUefE34D+3ZC2d39pO+iFM+VfMZ8e
Gxp99yySCh2Tt9yTA+9mXTHT8ABow76ODEgIGAVMN6nmsoiaV311J5EE0OUfnLDZYv/AgfwpU71n
h93xSkYHVoM4buMv8iXFgQ1CMoVfEe72aNqcyku5zuaHxdb3VvQbWVYUlBkKFnmjN0rlBv/fl7KY
MHqTzEosSYZ5wYf8A57lRyfRmOTwIGvLMHWfDb7RsTvPj3IZqz/rdoqSrBurF+2Cev4lqNx3cAPh
/xXQ3gtIzHO8OXZSLQgNbnllBaeBcyMIt3x6U6GNExKUM0N9CPc+HYNLQbGQvM9p5C9hqbu+q/O+
dUJ3BP3It/Vo2p9ApBh44V1OHMRTI23XHkxsWKUaNNdmov0s+DtJpdnTIa8YCe9QV16vB9ktWtFW
zNiFy0kj7uC4dBsZON9eEtaQ//HzUOSECch9X/ylDqc1lyW4kGdiYDrjiB3ygw4aC2Yt0IAlY3gE
nnkKpqXhd3qUHLt4sAfCG4tATA+bXgL97SWshASsZAKWDN/Qu3bHQ1eGJOP/1wS/UNdP+HLBFk0r
xS/e0ZzRdgPXveniltZymGN/ca9lpoYCyZ+VkduMMO0vGOnvIlW04Yx9kKoa8Ee02suP4y0YCfFX
Nt2JrsqI8mrt2W4OUPViAmnCLwvElnaLLPUJ1aaPyO8EQjG3NCdA1eiM+EiTcgAVFNKxh0mUVB66
fOSFf30iISX8IPEYduLR+MPbb3Q/qlIXSmVe8pd44mwDr6xNvJz4bWLdGUUtXSMpuwrLAN/jW/ly
bth7wQtXjC4vMod0esWBIR7K9QnI3Gun+aamriqmPR+vAE5d0eSl42KlraJnzQ8qq3s4A9caVSof
WZBW57TSXrHTa7+B3Lh8BeNh+d4hW5N57yuMY2ufQnr1QsqIDDnZvXrpoTeX0jGYtZVXC8nSynbd
3ALtnY14glP0h4Nv5KNIl25rS9zs4JBV/yWEkklP4IC0Ush3SDvWlPRtd4RGe0lAil+wr92OduHq
+OLfJJ15pPyQnn21vC4FSIrXczuU4yL5etujEodxyIoRyZDklycuChcmEfcxYP13CsKLeO8pr6ZY
AwGaWbbenMbnCflwvsYeNYuNewcpILE4XRTXheW/z8EoN0/g/sDPbMWlIP/XN6k1R/W7WXTGo+aq
zjkNKnkF2YXxMX9gJe5FKKEBAmM5Y3QGM55cwoVBwe3RPJVPNBTjqMQLK6mKURorWo9jA0+7gfPW
kwRdFNG6SFWsp+a5HJwACtXOlcCUn1IEo3U/CYzPfJnvg+bnRsSIw/4h7KcWoTc1UW+n7SqaY+qA
CO4E/O00VKwM+XSXe1VCRNYivTDFsM36GEfk0RfStUfQv8iyCcirhns+FkGczuHHWawT4rKybRwD
1qYCC5fi7hatFLs6uhd8DMjbvxjpF8ywbu4y39FvmCXYQg0Qgil+OTAXijQETJvjTiklL78mjoTC
RRjo60EXy45BwUNpBaBAs+9ZFtQ+b3fUPRqd4t6ShiOC3gxSvV4eGFfKR4DjGtGAvU9ioST+f6i1
dNNg0poeN3sezM6uqg6Fa2dYQhZrH+A0uhEskLXmQG/3ioDIZNLHTnZFZnlGDeVfPxLjd+zKyfIq
e5VpFkW8SefYWjJH+QrYtuXjv6NsB+AA1i7IaRCUcOTNctIeg2dzWiKL2MpGD+suoZ0hpzNwkIfu
yQFN66Uvai8rtlVWSuU34ysCwkgD93ot6WqiSGQtxnDiUiRxU68S3TujNQ2EWgPIR3WyCl5nR5x1
cjceiPz+cgzDokP9YxJbkC+mD46/Ob7nTxbUWpdh/uy5wsQ5EFdsbWTGtQnHBSX2+FKWjE+9Ulr5
UruCWJkEdmRBbFFPd2D0zNqimzsSINXOOX93kBB/swvYas9UK9pbmhjVjdzptE4beyStLdpsf+C/
bD1lYZYcax/R0BMVHTIdpaes7lB4ZlBxVdCHGyUx+ZqzFDubGSDZ20ANSEA38gSGLpuKuGLkI0dn
s4/zMBK6MMNIfMrdSEjyJC7xiWk3Y0xDY5kdwnHjUq2QhzG2gFEi9ISbDfmOeWoavcNl01ME2niu
fip1qvSRkGUm+Y5CroWiMmFNaMs5B3xHSuzbcil7e+L3YNe1dll1cuvzKy2uSTf/KT+L+TDdEfNq
QUVSHVtpiGL4/8wBOfJiH16kdMP+FBGZ2Xhu+S9CIdog1X81/RkSZmbYQwSCLsGkWq+YSK0okRdX
ZRBADHnbkXivEtwZTB8HZpoqrwOttgiioromXpX+E6REJiTZqkETm9hNzwJQamAIlB2EbhEYhMLn
eb1snZchvC2hau4ayVQY4v6hcYcctoT2Ly8k2kEvJ3DCBhZ53MrM0f7maN3ltzib6j+RsQ/XS8hW
rXWR6u9O1+7MYkz6HjAgSXZdIL7MCebq3eYpDXM3QDcAgxL3CJpOijIFppyR8vQFdkWgg2kcNnEb
6+SolN8JP/nCzcq8a3EPKQ4xkRxgw0T8EWuncEyWs1JwXksv8dM1qv4UkCGcvuhJP6uFiU1tmTtf
UY6Yni1HGRWsFMzWFm3Yr4XHUPJ9t1vuglFfDYlOF7q6VopIWRyfMv5gDOhoIO+z+M+Zc9X+tgce
zRzQNXcrNjuNbb57iAIAQhK3nDAS5tyNizRDQSpHXCoWDB849fmhMrL0OdpoyYuRsJdqMwOTZ5/e
TztCQL6NnElU2fKupbWRSe/zB4SN8UECFSmoOug5iY9QcFIb+43MOLMnajGy7RVSn/wyHSbjlzKC
9eYU8uqvkHFNloA4nljbLqMl1fJ/LOX0Bp0WTpIyyo3wnggiMrgi9+rnVTOmaTVxbo3dsRZJo/KZ
RSkXnbNUV8rpQSvtemsQ9Lcz/gC20+Tc8r33M7+e/l26+JmvAt60FR7bWexNNQyIsneVRfmx6BKE
Lcq9PG4gIV7Kjxx0eQd5GEAeG8elEUwKWxQ/8CR/T6WtDz3kQg9TGKLPG/3kTbLXHAuPttEPY8Nk
D+HGwUS2VgNeNNCipp47iO4KZ85uR3WT9lbU6jC86DO4l9Ih5em6rSpU0ka5F+vntdEny+oTMrtm
RMkJZv9BY/Zl3woxHTdqo4OAG1WPnlgW0e+QUE1AI4obfHrDsG3uflVoXtKHLDDwMsCuV9UjY4uE
zDB8AtKe+rl+Pe3+7vn9K367nI+Kw98V3/d0YU5lWsPKduOSVlGw8OO0YXXi0XKCy62RvKs8hv7r
vMSadvsGmM+qPGIAfQxEPfjpq5gzQt2HdAXeM+fWlF2TC6hPJVq927yi3zUKl/koAbwk37PHQOzj
BdRQwYT4TupCTQb8hWYwXHZZCMicZefXX5Hotkc2B4UtGPd5xGLV2YuTY/ruXNRRDbtKDPDKKx3g
wjcCx5S2skhZw8Dw4m/F/cVt/+nw4OYT4TyId3KlBURs4bdrdR1525JvC1hbf7m3BgdNXFCt+v9w
ANsNGEJvQm+SNgvMOdB/LCK8dJPOe9SAbdzRTcsrqbK8n/SPTagiFAw7QRTw+21UdApeMllenyol
9pLWf43B17bbKOZPGrdXhOQeYQ+RT2GSJXgI1wtL7wW0Xo/5it7YF5Rrwzmee0io9VMHVM3tdBJU
HRGZ2c/pg1VFemmsfToE5xgcjVBbhdwMOpLrJKhtVYvHy8vkPyvE6mKaz3NTvQf3CLSIwIxZ4X0v
UWNCmbvNx/+dXz6u6JG3WhnD8LkECif9JMMGie+l+f5523G6HoI7D3qSbfsIlrxeieb1/XwVOcIw
9DHLKfZ94VQxViqx79mOM4rMm3PMZPz7Zdz0nOGTkUp1cHxQ2tto7is5rLk2DOGyVi1j91Xh6T02
J55McPLNotz+DTP/+MVGcmBW5EIAfokpcu96OiXlbpqaJKs4QV1HWjmIQ8qK+2qihd8/bFs6yT29
tE40ZBrIwG1OT+UV318vPq9GTEPEA7jyc4dqkWm26Sx8rUaj2Mkn/+u905hoDEkvoos94jnJAWp4
C3T+iUzKOqnCgL/7PYZJwmMmIYGTqMLAL+MVZwdMMBReY8JkTfgHl2f9wPBwpfByA7lDjvMUslg1
2AIJKwhsQLmg+Dx+s2du1lMV6fJbs/b3jqJtmmgXa6xcMrAiTDCDYb1tne8wAXg3Mr6sovYFP7dA
/JVTtYl4p2FPLnG1Ka1IheMfJGfTvjNKH/APNCkfuoR3Ko3ONPvhldz0mGedpIabwoGrW5o6Tymi
V5eOLF0sa1asFZKlSN9ltD5C2+sDjZIPNfYqWOzHQqyWCzkdb4xoETfvSHEomv2OshWsbEFLHAR6
xcXYu4KzQeVxTUoik1I4/0a/QqOrcmPvTC1cPJjvaW54Z1pg9TKrdE9wSSdMjRE23JaRZmk5Acpl
FX7IFPLik8WuofTuoWkXYwtQWocdCv2H5ig6RuFo2BYkilRZ8pX5cjEx+mTu2kiJ2vuWlyUYYacG
C+Sj+lydoc6W+IHfgZO/E5wXfNtN882MP9xJYxPdZQHXuuI0uu9RIR/yMkfdOl9pvweVjsc/058Q
nUIdnyxosSBSHYUzGV4+Zit2p7xhG4tIi7JBxixBfvfeezpBylkgUBWvTxyGJ4lXsHwPjE8XX7Ig
ea61XFcKuBa2OGqE6+/19jqlhoutf1vYoca+hac0vu9ndFlJ0ynwu4JmT9SfAU7q126Xnr8XYoIg
ze0L162gk0qqY6VgrN8L5VbSksQsf+aOse09UmmAjxp8woL6hUGOBd88wpWr3YeKjINn2J01MoxH
AIKwL8AzYKuQrRIu/bhZhbI018FPum2Ga7dsaXZVm2BydEPMaLoLB3udgxVHWck3MkoEmklxpOlx
OS7zHWWYax7fJdBSdBPAEEGDZd7/Tl56fhtSTd9cadcusOdOCqq3/Kpvxy9xWtCbhq3B7liGewD8
G30HWVsW2/dRdhjGY+vzVwn14iSVZ25qzxI7hlq4PcHNI4B2ALLPqgKgTARmGYlkX5UcgpjoSyac
4O0ZvAGny2ysfa6axm5BHvzdnGCZslQXjjbHcx5pObK5kgZrLICVlbZxkkZYDAwFm+D/DMRvyPLq
D2OSSp3ZJoOlKZqBWRtZMLnmuHJTsDtWeEFAB7AoT+E0pgoNdZLVPEHruN4ajaR4Byxgr3ujD/uR
kdY/J8r5VqIlibOASG3l8H7tDzbFyey4uwFy9GLFqhy+BLYtgS5fpff9WCae5C9AAwrTjaB+oFZm
omsdXIwZdA1apiW6s+hQXuljwLLRXtoZ0ssdD9Oc0OMQEObYhJUAqBAUqmqBT2olZhK8qC0vTsXx
+RtA+xpm2b1VXk+G0XGl45DRZodAD7y63mIckwTG/uE5QQDZ7Ra9LxqIGxyLOFmKaTuVwPbKCR0u
AdC0xx4Ays9NZn/O0zCv57c323JUlAHQfh7C4tU4jqdLdBIiAvYOXuhEjJapybLRjX57MXCDyreJ
re37fOkfQuEXX5H6d0nK7BZK1WgJ6rHTjnIbD7pqFm2aow5D/gK2AFMaQt/OCz5ZIIIUJeP55cd5
mg/BUr57mRhzviWmNIjEK/VA7TcXgliUSwL6Bkq67Uk5Bsep3bRvX0n+rdn8a+Ui7PH5Kepg1gan
r3mMu1MyME2tjsm9jkzRxr2u7DUXNEqmtH3jFPZFS2jlVpXq6vyAJz01HRkZNs5yDIlau/WtcO+e
fiU4ICSUGpC2ItivYrulNtiqTBvD3iAEBKW/KU4aKT3Hm42rLsx2nCixKTpGh4hOAixwRHmsvvEA
5S9/lB+ev0wV3+LZ3P9J630OWerFhirk2T68iBOQz07W4TDsL1JjzwTxbZN3CY1rCcHErd48PKkd
rpBIPqIs0TfZC/xgVFB3QXVYDAlzuxYqCgSN7Vzo+BLzSY5fi6moJS9F7Dp49AY+ZEbMwSZM+4Z0
W00Hls4EsQLP59Qtw/+fxKjEpTN9Pan70JW0YPbIsaYkk4TS1+2d23ZGjipYlrj39QwEpSn7NUTj
rd04lDseJUZlzp2Y60/4o8Ac+z/vVj2G3poTiSZooWVLSTuZW+4c4RNGUTyo1/mqgPWzOnaeYcw7
4SPl28hGhAuLWi0EMctBndVlrAtGrrdNQZlmtMp2whPCIPoXTcMB7E4HVnLZ6+u189Yyoz3p4eIu
2zMZ0pcQCT9CXS88G3wPJKIeiQVsuSE66+aK2qoVGCt3aGOXui/J+kVJ2WchaPFG404DxYE8lr+X
5JyvDBtCTnlYxgAnou8MVhRTn7BvYg6Pf7k6ua2oIGniYiA2lQLMynxHfbyV/5U2uH1zlA4iyKZc
CdhCPeYaHx6BnwFOVYnddHYZKC9w7h67JYSpoDJFUOdoYRobowV3SPQJvy9GIjPdaIWml4Sl2RIc
yxlE4G/8mpEaAIMZnjkthBffQyOujTn6cyrgm3raBDYt4MIpvtR2P+f5VVQGyXl16PczaHMzcQuH
E1J9qu22siseu+jQ84hEAs/bv0cSUKqkQMBVmEcuRlAIVixO4XEmpxjbudXotKQCaXv+Fjyh3387
I5uE2Vf2b+NlLmlwkntki9wPSI4GA1C5AqWfVIfJfas8viBBkMn2x1APLZwh/VTLhbV6KZJ/UYgD
rYQFjh0QiufWU8NP638pGAoas5s1Lk2fjokkSyX/3u9rAxWHv4tk5NJ945WAOEvJhZzmcFK6qW6E
ToNMjpjiX+gj4LWldf7eiMnLTuLphZJ6JyDoSnGEtheuMECkRXsYSSfN1rLow1R/fu74KFmH8U9S
LQ43+aO5P/2a/o1p7rIzmUrWiw8yy3ZYUcALoV+0nT7KsdnGpjJBW4uxqFd/bsbxhYJ9sllrzxog
qXxOZxj4lFFDpYtqxjiQvC5wKpKO0u1yCts637I2WNsrKvbjZRE6zkkttVe3gHCisysYuREQb4Ha
T0kLHjNVEGgq/UhMCg3jAmllUHMOs3VBZ6gxqMhAT0TR4W+tI/Q0rBRVssuuKFQTXnUqbJhyKb5i
FGMLxXZ+rXuldA8omuKhMdvoxnzdKm33O2mU3kmEXQMPI4f9s/Xp+8pojbTBiQ2swYCpdkCMIKvV
GVoeK4TcMzDBLTm6k6NLnRgJB5YGR2kzz6rp7yvqpXY7lEPtJszdPyq8NA31T+T5p0q2KNH4jQEd
75fPd5DJD/Up3rZDYiwRaUcKPQ8YnUsJvfkqmnanDzEMMwdz0sHgAMA2C6yuOUxVOlJ+kITTe9/c
76OAker4XhUer7rV1DJUC7pgzFFX9YG7yY3HesvAPf/SUE4im+gJIX4DFXGhxtD7QllLpl2ZnawD
DKFS94IrvkkqFraPD9j1Gqwg15YwnrF7lP6NPAlEp7/K4jVbRSm6yJbWYlvdEuiRiGujJtLZLY/u
4r2PxbmQsxmMsFKQIFYcwoi/LflRgucghepma+QrrhoFppxvfBw9UXK608AmQG4MQarYQLQyMvda
djdYx9xhVl0JVRa7YBqUoRuypxxhQ4sdWnVcTqholwc6E9SHcms0rSbHQg6BXOfyaCwB7DiAC2Zx
F/kJjrA4TugLJUqUSH4UeigC2/ruI1icx6jR0A7SvHvuupve841/prurdo2m66ufz1hTMP/CKkeX
XBWLiCwzTyyHCwtk5rjeXLY4UH41ABjis85/4t1nwkp50ohl/EnAD6LLjU6RRduqas2eaoaN0LTz
OMkQI16lQYkjOn09504ez5BvhI4bd/0XMnAC1o0tWOf5te+WjEIYq03yVyRklXIno84fTY0y255L
2jnEonS6yjwajZFpL3zbbs8m6+qzQFZzyCKeuieeK6ZQoNhXefEQF987O0nrsphou2aLmoF6k1JU
aYs/y//RU0/w8tXjZ54QH2RfzdZibArfy8z6h00EiaAQ8CYPhV7y94an7Inr+McNMBWoKlV8ZSNY
L8UbPKt9PcSN/F4oThsb+MeflLsOK7nyWWhnmqLs61Gl4+sBIR7NgIJLl+Anhc2eKmFnq4AYe/b1
D7IPQ4BXcqABIkxfcwIGqkA8SzUEOgIstdZa5b4C3rWHV3zqtYqu+jAGPidccwv6KwVwVsJfhCyT
01byfYGPWIccm2nrUz2xrEOJ7TrCGFoK1e10cKltN3PxUGTfkRve0DUHg8MsNgi8FWy1hKwMIcnd
5glc/IqHogeq9kei6RNA7+zBSu/lmfgXsXktJrZ/p1gi2VUDttnG9odVlO1Ohsh56dti7/OXdOEQ
LGNfkEbgKiAqQvfl0IOt3W/yULnLSDOUp2R3888D6Wq5NGnUgYsNNKJJRTiawAUpU0IzLk+KnJ5l
g/GtevXN/crV25yUeiychnT+CV1vJ+UaI/iwBJdoiR9E2ld+lwHm0vge4EA0WbgwrxYY6paHTMQd
NpO2VKt/PdRb+SeH3KfI0us6OFpkceVRF9somJqcfyetRxdl4SyUnxbAYtlj438d4dCmLUULN7YN
pnQw3npihVjl2WSRxdxqx54F8pvHoaoNYTaZbO5rTLqDWIUcJ7kVtSjaAVB9n3HQyqD276e88F/3
OcGYzG+a9wUAcXje8cLASR6Wm409qyisC5Bbu/eOjDQXvK2ESvYchENTtZ7v/v4F/RGhpgNUvttF
L/09sCwUVJGcVDNHFanajL7HDLxopq19SbolXcxMwtQLhOok9hsd9CeCoHkRVePWvbd6UsSD5LH7
mf3iJzU4X5wSNKiWWuU77kBG4q1wRrXn6EnZlgQvdKh0BhpSfHWsttbLJKmVypmYBJmwVD1sDGvq
mtfbypE0zw+HYw3TPHBv8RkHFeVkL+1uXiX30FPpKRHUfPpB8+ZXJ/+s1i6N5o5ayNZJkbLnlWs5
DfLHd1M2MYV/Y1L5v/kSKWhTOBPeikPwupwbL48hrznZtd1Esf1KtNlOBVtDaXC43dmrYScmqX4W
OYqJ0uMmCYR3P+mZiYl4sJ83PJdYN9Ju1bnkDuRZvgq+rXDqXd5DjfxkyLka9NznFi6FwLlO/Z5+
Z2AxC2O8oKVwAENHpogT9fydw+XNrM7wdpz8hFrj57FrMEnEhLohMffQlnitTiobScn0HMkIIQ5U
bOiMMizSnMYNnf3w43hVtjE6axnfSaEVn2RxoQo/frO886pQsIf417ET4/6XzaodHjMeBV87lg0/
doKp97Qq0rJUFPi7Qi2VMwICRb/mF2hTrPb0lP4DrGht2vj1NiT+ztSQTLei5nI5jWa8B0uweOx9
r/uR9lfXJ4SiC8r330S7imn1o408Ci2glnAlR65LpF+FDAInltxKNhccg91NRHPT9jLNlzVVEROn
Cq0LK7VlGc9IWNx7rhX4wkRHcaYV7ez2RbirUFlRd/ceTUPwkLoj3YmhNLl8q1RN9wd7qRF3IZcP
k3ngIlKKWesJnGRpWnUqiLKDscTqs4UI5Zi1kVS6YVBE45ZBz/rRgXZhjkvtsJmYBTLLCLwPtoEF
XhUVrh85gPrSW/649Xmm1brb/0Y5nNuwcoBmu5y1aQF1NB5vtJu+nYvMZanXrBqHZw8ASZTl95/e
q2bgLFvE/vbv5TAAy/U3jPwaA7ys7rsrji/jun/Lob1xSxEKnaGp8j97bZaM1OYkyGQzjYRVtrOp
kyLIxtTLF431YQEvIlSorWZHckfCSPpMgkalWAkEIEy00E3eIHIK7cWm2HyUafzQv2SCe9NCmHCr
pPIjyoXmenIx7hp9EB8tjfgW8Mst44fg9D8abmU78WwQfnMlphq+0HL1gRBAHRO4likYeTmYl3OC
R1XoZcF5lXLse5NrynK5/iDwwETjVM5nDJhBliPOsPOVMU+nxMNDkpcI3X2G9jaSjjxj20qq5BhP
Nd8Czv7ywneF+Ozr8R67aWz5o0FXW9bCfn9tMqA+UEXU1YmJmFaJNHf/dj0/ZLc0g9GKFy0dJnDf
a9arI6U1AtaK66+FGtK2y4FnwFZFCHuhZoFPNBRJVft/HvD2GEcT4ylIwqjrh0mRIti/7sIos7/j
6SHFXlqgNUch0VGMLy+pv7PMF60vexhY2yZkQgMh/aJsfhszKb4iNfi0fiaUil+aDDWecncoyYtG
t6I+vxhXWpptMzrMPsWH9NUfcXMeaYEVWRINZoyAEb77cdKXkExg7hcDuok5gWfrW9Ta6VU5o8Ln
m5aY3cpwyD5dvdi3Xy1kP1SFc/lWMUpnQaGLUeazRCjtz5e5v3Vjr6Wb285+EshdFwxsBmFmeTAJ
CXBSKyReluwxsHJl9xQs6WDHTdIll1lVsLHcrGX4KFEywD1SxXB6pDPV2kRDRhYArqfXAdLdOoKq
kWP51zHQ9nye9zbP2W/CswPaTdra1C9bdEgypXm0sxwVfsR0QIuB22nxT96dZJBS4aU2w168fl63
OFLUVOecyy5ooqyAwmN1P3jcHlAqrioA2OJ+U/55JCJCjFQ3ktg+o4xs8cYLj/xqU9HqI6eGSg3X
2vs4IDLWOuASqzwMJcdfs+tzDtox7qWT+E/nopUXOx39/eU0n4CsRUyOr8GziiDzmZv7DT3lniCO
jJcJ+2ArL3jBIBGpgloJ01k9q4xG/iz5y0kWlddqO6BMXGk8RVEspZsxTIIW7yZE852LJ4C7lroP
OG/PVPQg+EK37mBDCHIa84sVWi2MWu7ZHac0zev/ChVEVoGNJMR1MVQKAWBG+/mosrxJBCLzmEiL
N1A8lIBUgXp5qz7v414F1tHX+QuqnD72/XEvUne8/YsKKy0UkeigHpEw968Qjq1uXM1H0n7V0Dd+
Yyo4F5UmRpc1Vw+QWMZbDfRu+7ehk/vnB9ZC8GxfCsEeNmKUyMlaj14v8F9g8h0PlrEww8hl+zJS
EBByibR6dYf6OQPd2YFtmWr9E9/tf69thLBRHJ6Y5QqkQaf6BpB4S8hAeXqkqyQmqSSYV1SPcNW/
Sr8wLGGmoKEgj+dT/aToyzLh12oif/kjVIuSuCu0yXfFuEbsNtTqD4cZ+nkk+QZ+Hf7xcZ/EaADL
3knXi7BmRIjw6R7Pg/A9TOfh+Aw/YhwHM1IVB+Cb7PySV6WxY2Vw7JiR9twJQPetzE3X3NejPWL9
0Mqjo7LCJhZwsBjuLYEKnr97F/lofarMDgowX73FdD9JvVUYm+lbeHZ5GGn9+BLk8cRsByn9BAaC
7dfL7CKozAZDGed3NktOOwVfWQKzKi2xIDdnu/BLlYdh07s1VBzcczxlIfXLcJsvjCjM3TDmcxbo
432uaX+o2bVWoT66qMowQu74WlnHs6Kb8KKewNpGDr6KP7veZH/3i1K+1np7arr9HOJwyQ+WRflO
ZTJ9xDOGAbxClkk7PUljkfAlxNIrokHYYdwpBl1G7FcXtq6eAWlQ4dy3KRFW4rwkWYEvQFMQ0fnx
HV4q83j2iqMJKLW7CzQn5hf5nMvCT7U5MLRNxxi3Ps6AGwdgeEvFC60yEXRjv2oKGzz1ZGEW27HK
YwskGMswxL1Up8WVs4/Vi7axeuiKAZnuIyCKT8L69oWSze0VQ7G7JciAn3C0AR1Wi6HuSyzsI2DJ
q49c7mrHCa4lJzfu+Uyoe1wZkUYg+k8VJW5UFFDWNdiCOvwcvC9Qy1L/cHCBAVNp8AdSIGeIziKs
XiI4VqWZWOoHuS6/M1uSB2C9pBlKlVZeSrQrxkqAsvHQbsziII+xCcCoFp4++SEUI5X2WEUeKDI3
Dpks/Dk3cgY+FX2MH2XwiuhWiJ7L9gJyS7pwck8iSI9Fv8pKNV2i7QztmQ/HXhOn6p/Is4eoTPbQ
KiRPIkKy80nI1Mzckbyik6anTQG2kBsuL9P4IBzewlO160f23G3FM8FGJeJi3o64jhCvFNXxixgG
C/Y1Q2lGtp6rKOkJiGP3+RbXSwh9huNSLTYcS/UqIsErOhGhgUuxadCO9pJxHgPjWM6FM8w4kv63
L8+IEoAqUiQYaAAWEVyjj3UXtZFZG0XJcxpyRie3Ymw6ghxysnZ4Q+NPTJD1ZKS2XlHhqU/qzPll
LuwrmDSJ6KPumJMR6dRFf134/XPnxy80ES96T4bdFdFnncxvjPx4EDIRQttRw78uXh8+gLaXGCEi
9RZE5lIdWpn1YKzjIPcottEV9XlAn5xyXmNnc6Qp/Km/zPa2eq2FWbolxI0vV+/tkjHmArQyadsX
3dfapfgxZd1DZoInfxhzfutT1lglANubfwQAG7ylQmGhPGtsHLt3vwCm+Eydcnur36DFB/PoOta0
8sKdFSeqd4JG2Bq8IW+9PbgGP8bF+GUMiN1JtILK/3Qyo7aSAezehE7AsIHMvnP1FvBKiUM5OTC5
SDqbLsozWM8wijq5+DCix72ZKsqZggap0JK+DGYOO0HNP4aU7Pq2OLe2R4BYY6nNWLFuF9ZRB7WG
8KQfOP/9eRGUMwlGK+ePxz+5YCcEQ/KmFaopU5wVK34yPo5EfKR+x4nDe6UEojA71dB2t2648wI3
FMoyCYOYjAxkhK3dPMW9JEZ1DEFo4fOUg4jVJdM79eXr5nlNkAH2lpSr3XIZPcgao+Kpn53e3MU0
Hp/CjbPXTr15NbwtjtLuLY5d4ABuhYMhVgqEa2gQeu/BZWOyrT8ysH/esMxHQnmdTtkixAyKclw1
WxbwHouq8JJjXNqewSyGd8LZIyunU5UMICKXJxoOa/nBfZaR95eZNYX93FJ6FzehJNNGILqo/48s
gGo227wfeast6z1t+3YneYgHtz6mTDxix7QpMMK5ggCFnrMG51hCt5t59GeGZ6WhT2wjq4ep4WUe
1h/Hi5pEkBisYAk5kAwaa4BzZI6+IcdqrrXE30BTPkzGZqsOmtgPm4mzGfxBy62OAz9wp62/77xc
oEqAJN1ncsFp2h83TGodvyrwXYCFbS9tXhi7HWZO7rQNXa5PslHxldINPVpf7AkBtPAFZLB3HRwB
Q6zuQIBxCQTDGI2fCvHZ6JHjdqnMCgk+Eg/KUClwSJsjGvh8BhJvBa5+cASyNRHGZDApr0cva3nG
qj9DrdWtP4pXEL7WPWcKnirJML7QPoxKxfqyHpR82mAQXEZPN/zw7x708Oe82LZhqGPe3XTi9uVk
+VUz9FvFJGhRX0TdiODvD/1YgIPs08EbHE3wye0Rynxyu9eFYIRFeM6QPsSma3IRwbRG0tXUuoYk
fRvnHLt1VKVLWZPac1VUehLBghDdl9cjZ85BQ6Wk+EnVRaDxf+htogk8P5pG5zPlhiFKgTTRd3Sl
0KYKOICBg+n+1Ekf52BqVhOvwSrONkLWrCLZB2Deh6ND27TzNlrWpNE53AgfZf4v7IH+7D7qBVLG
XuJpB/NqMIbiSWpaGMIDKc+19+sHQpUX1Xa9epsDG3hrJNO0jQGmWAJLIaJgR8YHEK4hcmAGGKQI
Zk0qSEVieLJB/du9ezBSR+Kp0ZZT2zdhci6OY2Qltke221uaQCM3116D5aGljZA153gzw9ADVdK9
4DziDn6zxYkR64QMl15YTR0YSZRD6qJSduwCjSuIip49kzu7obKzJdmAdu4XMVx20OZ2lf2bF1Ya
S2LDmkiyFeQk8dtPzmLKMuJfxPnlSQBJHEpgdtMzO4+6BcmQdHL09va74hNH5TzqvrB11RuC46DN
+5xglTjjZ0LhaVjdxApKdlQR+NJFwwYijDviZDA2iDPYyopeP42gM+++vl7s8PwYaQ4EEWrBBq76
itg4esf3RElkHkGmxN+r7E4y62h5H71c3esvlaRCVn3UfbpCtjufCCizZWucqQLN9jxIxDOldRGz
GIAnpwfBANrGg62mGV1tGHm4uatQqExvc3JV5C5bt8yGb35dvN5UE198kZlGJgQEszNb4mngmAtB
hvRMWeK0/0okOrCvJcRs6nGIrhQM8j6jCubsfl5rg2WiypmyoE+dIF7Ud4wlCnc/AYLNWjKH6KWQ
mVq9pTadv6fk7vGvHMkJCghDHD+E/46P8mdW0NB4bu8Ff1nQH7dXMgNttxtNcxZGuYmKQDQliuAN
Td47h1WC0ltVeA9I3RBFKIlI3eEMBBwKeY6KAVoKRbiRnYZeBeSXGEzLrZUgUQYzy0zGYCKSs9EV
SX38voXYDrbaGIKa0MPGbtxWZAE+KJ+laEGxwyxbZhi/4oVr1Xr7JgNlW3pX5V/TyAgO3MiITRXi
LFPQwz5sv04GWgzyznW2WubDPy9Vwolb0rC4WAhUyGLMFejhT26/SmqrcgOr+I2c6DP0UXaAeMgi
DKSwgO7f2g2e78vtxAt8VsxZcJtHNTIw2ErnkGL575WOGHxOamjAjNUNdBDfqNm49Ncqtikzvufg
9YSUFJY0vXsf6gMXYYRV2SEY3W5G2DAj8EhvV8GhBlD2PNm/4SZgIC9hRe6CrZgXFjuYfl+wBkQk
qkkcloQJyKgZDjSydK/mZsAoDeotkyhrsZjnQfqz0EQ4NaZjw+FfZZfu5kSODs57a4RTWqTG0Yjl
WnUAsBxJDrTT3iNMLu2vryWXuQRYy+CcdH8PQpIdyDwh5dRd0f8tlGHkMvmUMZaVVelRl2OZ4S/i
XPEUi2KjrzxthH/Y4Iohq6JC4DZslZF6AzyMq/WoMo7ibhAjDh2Dz4UE9uRqOd3LRbhMKXEWlael
BajuMfGk+8qsW7iE9OVkhI76wbqTGHJ7RggawqRBAf3nboyky8HGkynevb32tvpfTV0JCB3Spxuy
p+SispdiK2XIntIQ/zzg7mX9KAo/kLGvINAavhGLsLH4+GHsBildPQqsjiNx8hA9roQcZcZUgb9R
a6GO/tHHFA206uHV+FhkXFbb9beTdikeuLzE2/3gF4YC6hCFatX9AuaVLUbQ/5fMxMZkhPvC33zy
nY1uujHsz+4lvJTDlR9eKYIjvmR33133BwWzQiDHLDUwxoPoUugpLZr5iNIaa9G0AqFuk11AowJY
IoRI6zBkvlJLhF3oMrnlKOe4q82qLmzYubDZR4oqoRFVcUQFM6HG9lU47oKDSzcu/MlRlDGtvKdN
JIYPB9RUL9yCv57BjFbduz4oflUtVEVGGHJlD2xFlwrDhHB70pf210PybdVqdDB7kP77LlsCVg6W
CgPL9jGAuQxfuxCDryyvWJhQYPB46lAah3UXsqxYil8sOeSgvydVe1IXWBRxnh/XpjO8ugel9lkR
jMPsilDBjtSWoTETVgsafJC0TDoN8vB9F/ml5adD91Kbjwtpbee1gMCh/NX3+3tgLSBcH1Kp7ppX
andvrS74hKz2BPHTZwWbFun4vRe9KTrXI21ThtN3H8xEVsa8E5Sp/+jiD3JduBLw0wSOZSx4twlh
ohQN4xqoQ8Ye/R3slqUouZcZSLGBoCQz7HVgwsjnIUgsK6k7rf/3pSRrW1SadSJMIzJ7C3kW4Z3Q
FTj8myCGMHkb5HHH3oyEBiH/iZJ7a3ByYbgoM1KLmRh4UfTOREea+EfcT109rHLzMdh2LvS1DWdl
kTmZAOrc6HwlspMM5qrqcm+lrrUsadFkC6wF5Xi/pwe20Er8a0RGmany0ei6ZcE83JrEopHBnlHV
8cPNYX4DABhOX9d2DiCDaeVIdeq8IQaqSvTCp1AICX1kAGdZAvvAfkAhpk4vnYLv9oChq0F9zWhM
hw8lyjrofYTFaNCLPiKJ1sMiYzW1lROYcOHvsaUc14kBNKpBvc9gEGyK9H79sjBli/BqIiUG94+O
mA0VKBn0zsWxKOwwC065CGYaQ5ojeJD6/bMq1uk1eAakuFXaa4cKkVXXHIBM+RzELntGny+r5UoC
iAdA8vpbc8zaaSzlG5l6SHMxJ+vYXHNM0bYgabgFtnVNzUt6DxEJhKDMGX26F6jkysRMZ5N+O+UK
0b7zJMNJ7TZtocCrCV1ndwHsLEoizsKmeKQjmaZ2wKR0ABvJl0rOUatf8m6m/Mvf+QhIZcd7ApD8
Ic6NNaiOgUTcnzu+97O4jW8lMLb+LoUhBJzqHHkUYZhdJFSfNjSdpLigzgiWbWjvebPlcwvqVUEI
/Y82cUcs/tvk4ZBvNmS1dBaIVxn64U8j9fboQOp3bE8oJUqSDE+VaizJZZ0TdnhgnTF5nPm76SGF
VgKVnuusNDMRJucHR5ROwdu+Y6xxcvaUIO/T9N2CrVLiFzLh+F+dpXjGoFXcrKwEioQnDXEI5aSv
VLo+u4Dm0oX01VFCGv2MAfjzWWRJekhUCahotthHBNek3y7YbUiKSXVia9d0hzuNGqpaN+npi7Ns
IDa6oMX9WaIRpRc/noHU/9Dh1ctJz7hgvp82Q8mSGWqE6OEEuntCcoaA6VHHIgf9Rt6+lk4TT5y2
Boy2+g+DTl8xtFZimQCMvwCBssKEQEc40Ro6linszz0XvSmd3gsL7jHhlwz0tcdBgynHD9YNfSG+
3X5tHTerltzcT/MnZFcztW+JIZEkLgEMc01YhITnBuLx1YUG5FpIeUkbY9NHw2tpeahPB9dEy7GX
B7I/mNO7CI1LUtzZyxXwFiXHa4jvGhMLraDHGUCsOtEJeHADEBwkUzrvyjdaVWEzm25KG10e1CHy
XCgVX8FxqNVZrAclZXnNwPLCEw7T7cwVY0VBLul4BSTiegJX9gvPCk9HaPXGVvpJNHJTSWUqo1nx
ykXwZjS6c8H6q+Kk0Efi+W2zKKWUdpX4bCBwKYJTm0Di/9AYHQhIYi94ZNuyEmUOjg2xG4UFQrul
zLIXrLlidW/9iKslwmX2BhFWkFKH/ZedOIMXmEbVWv2H0nbWrIe24+LHYDjwjwPNjD89ziZkgaA2
O7sZuaJAVu3JDuhltl9j2bmSiE5cuFgReeHU8rENh1Xa2KBkO6S32DOu8ZDkoQQ0brdzg2qGF8iH
AlVaMsPIo9aQjaTtcV6AI5PrHNeENJ/pLqeActCTMuDe1lP26m+yUtfgr9bfg5Tz+MzqaqabSlkC
hZoZj1ouqoLKM/Rim30Axuavr4PiEMyOCBTw6hrB7f5FVG9jMqSOVkatBu2bkKQWIUGcKoO716R7
3pP7POIM/b+kdr5YrSeTFitkS85GrDs8s8ZVOJRySP9SwlRaAWYL4cTYV+F+iMeQxJ6/RUYRB/Fn
8dKwdAmiBmJfLjQ9EAkCcTAIZHSJ3FdrW/KcsMuXIoeQ8yBJEPOlJqYiORlk3IHonlFPtoQDfF1o
lPcRzudU6Z1GAoeE8VvlNgBmSKmmC8keMRKx6pLGxC2gJuc8lkdl6wrfPefKwSHoBLvNVVUcz3BR
qaaxcxCu1bcdxr8nu+vaBQVlMhfxtJWwMjDszrAXkYoXvA5md/XsoMIMSEGw/D1TGpYdMnapYiOP
dtEhbhgUJ2VOfgUq+I040vkmC5r/sUpCZ2TcX4BFPJEiv36olFJY2KoG29bzzYwolmTjiQXsxscm
4x8d9KbHfeC9MD6JGxam4lFZx1CeZ0w5yMFOK6+Kny3eTk8GENSndcSf3Wdt7QOnR9dRy93BtwsZ
SLAE9QsdUKVcD49DU6dlXwo6syXSI7/B8ldE+i1MCOkcqIbdGOMt6lzXDY962XQ74ZDzVAXV20K8
vHpF69DDtF2WX/IiDVuUxWEhre2+hrGgkHgrKbZUP9xYTpaADv6qoB1y7cEasYud6MP85rMThq6V
yQPfdi5eZwyYXGofXgGxg/lXIB9Kgz9lKAjRE8kxfmXH80iVky1MKpUUEWCT2myQz8GKJFwsmPcd
V8itWht9bCrUGjdLmqeY8v4xAsOZcS2oysgEnH2SOXu55kkmsksboa3g+kRqu+rNCuplN02ntmdu
kRVTDe/s82+YDZn+4Qnxa6rxxTwjlGKm9v1gTHX8DXYVqc/uRYhwCpi0gjq6MVDjVnq9Dh0FK/oI
CskoQoz1MewAeoWIStbAASNfy6g2zRT3qqc4CEkRZ4yA+mBR4kE5UgUWXwlpJRZ8Encrrw3Gsk7g
eTMmkeBKQ65JQupD30cr4fFDXgnvFNF5nATD++VjjoSP3p1Y+IiHwHgCz9E/LoMu+E3lhYfiruu0
Kdzv07sx+e7UOc/89Tm8SEVbYQRHKG8ii5I3DSPRfBK0/u9zIIT8RQXPdXG1WQFRvgDZAFuyC8IU
rR1eRjLH3Zs5NAGQDMm5YxquvThjqDdcPkcpM7UbiFL2j7PJL45PhKFInvbpNwJp9SUg8qjJzqjm
M9ffOwSIZ9PYIQCIhXupIu8ZwYaBAUPmG5fmabjHTqKZrNGEsoBy0icyrUItdCmJsii9oB4Ql3u/
wUj2SJYukty3SNPAb8w+sTTBSusB1wqHPUUEeT14mv/gzsnjzwpp2CJd3HdOGevRXYo75yXswF3A
SuWpDQTeaB8941mcgeLOkbgIaUEy95/IfF44BcB8VbTAvNaKnk/4yo2UaVou0dfkimDVtX9/CqRs
ATB85rkI1EQOAzyrYKMCSzikja+GVZhUB+nCeF0VtIPGVkmfs0PPHbOx8NvWXY9YtIfUl2lCtLkE
Z62WgRPpDZcMEtBZ7pCQHxG2dmeIBD7FifbJzRNZjg7lNkvbTWwRpk6MH1iTcM82PtgbenAWX/jY
rnObq25DtyQIOupeGLi74iea5rOj1hm7jthDf5gCiUtlrYAKvIdlpVAxk8Z/jhTY9+PuVoUwbCQ2
iw/5ZLjEfufC6ccJAdSW1zpWLaKy+9UNjb9jb9UEJd6qz1gnVV1TLgV53FQaGV4bS3Du8A0I0h7i
4DHSfLT7HLjtR6jj2JZLcfubwHRCmZS4SdkQ63Og3p0mNq3vDu8fYv6VWU+4jODu1L8X5QIILND7
H0J9ShaBy9o90FKVFB4bGEhMM+wnh7DzUXFuEKjfFeiPINtzpYMfam78iL64sKrTdpLe4foBTw+U
ggi8jYLc5NcSMp3Q/pAJrE/kK2w3fDRLYfH7cYQGvgrUrzrn8RjMNXWQ+F1b2E9I09/pmm06kqdB
w4zB84O3FnC7NNKXOK1rc0cuyDTVBH4KJnJnCXObsk3NAVej0qmUJFkhDZXQGbR/HJOQtvSlPp4t
G6T9tgvaxqQBxad5L1HOueSgGt/k/fYhutIn0ymq6oXjUQHvxJ3sW9JxsfOAOj51TxCshYjT4UDx
Tapc6GIRPsjm4m3Kr2Rw4YpHgyT1KrGtFz49XpVK7thYHDz0LeBxc5bsCS3jbJVNquYfdRr012mQ
hWMMd7GSlrUigmZ4EbvmJS3zbCkKA1xGjwFBFel7f+heYzMg2NolphARZaXuDzVGL/8ywdHAeol9
P3qGypeFARlOzQV8f+GThnOmE/GtDVcpIAAQvtCwhgSWbywNpzkOHDT8edtDJ0a5slVaB7RvsNwS
QGeePSVaxJwZv7FQ1aY3VCk1NAeYthCqLO0juvGGw9036RB9nOLlEfmzkiDkmXiZZX/DZ3A0hoF9
wRKW6UjIrBgJm7qe9tYnNIyMnRf4NIBB476+u2D7DS1pUYbSoBzHgxMXU79SyF9F1VP4E99IRnWY
sQBLzrG/8moDKpl03HjRwm80zttCyIQp1uo9pPgeQOJswNpIm3nYmqQbwkoNfAMfHiiFLyaQyHC1
LpocKPz/gwZ8XkRaaaBtPsNOJ7lwZe+fONRHt3/0cDQOd29LZrUv+NELl1B5cVKD9Bg+J4YEf5zA
VXm5DjyLFdc8d6Oll7DmMsS8KowPtH7IU7bO8SXgpVZqk7ZHKJSm31V8jDdmCIIg7zJQR+be+h64
RkoNCIb6XPlnDInf3/KEs87mPy369clhqLNMTt4TKz9lv5iau0WlThcD97gjRld6DBNkyvDd/Uh1
ebVfu3aZqmRsAwXDzcwDu5XKQyTAJeU4VIxZf0aVwD+s89ZKOFifvO4UkhslPvtDIio88fI6NhRd
S87osWx7OjnnqfayqSNXEtsddy+n/TkE5hkdaQyZKwKRfAVhW0q1IP3AzlK07rBz9PeYMEgD0+wc
68KwaB0qwXdnBdOp4PRWxsbkdzoPIBYKaFo3Fz4u/vLt1rDROjucblYTlMQSihXFtC18GuMjmShL
uvGuT7510l0rTXrPDgpXMZjsnqHXJNkznISjaT+ATRvT5Wpl5TUxTnz2Gbv3xyIFPEMvpHdMrpdp
edtLjadIjXKV/DGRvroRISuupiiqb1GifqUutUPnaaN06HAmGdZF2nZ5eV7zDmBk9M8KB7e2oBOI
wgeu2EVILdlf7+/PP7v1FQSPfAluwQt5nUj0IUV3kZ/Tkdp4ii76cnptqqbecgRmZYHyESRSaWzJ
VC0rXv3DVmd5qM0SKsWmPsZOJ1sW7m9Of3Y2eWQkUXIjsapCcX5Z2/1AQDnqf/ZGe3Izvc/13+oE
jH7DSV/mSVRpspuXK5MwxUHCOvjQbij9rAjPGW3y432ktIzNJYOCgD5BwXqt4g9ARuSGoc51umSd
1h8XKD9CfZpXlo3BZummDeh4vi0EuR75eJjM/0YmV5odkwY6qmJY61oh0HVa+AN/GMS9+BGQ4Qf3
OuWX9c83h2mis9yXpU5oKcm4vWfqKb3pihKv46wcFkWxbcpwMM3SE9MwqJjUKVuWGL0Y6kLfB8oB
NAoTKpB7GqxfkvHDheU90HNyhaz28JXo8C8f4mkJXos+b5Ov9G7xwWmG9im3uHwGthGj1mESSOiS
3FcqmSrSJ/ZskqNOSCvH3kbC/S4eBscjalZrQAop6HsugvbKjXsRIoBpngphYxxlDsY15ewXF+gS
lRAjC0Iu37bCtMp5Y93TrXwAPJB7X1FhaujHZZZHzot86/OpJvsbuu9LKbC1LWXj4TqEkcyn0SDA
zIho9DX1bBAQB9go+5Z+hmd5+CElew5NYx+Ve3wfylXVTpInlBHZf+7zMtEomyD3pnDRtqs4xBhM
Xs8/Kg51PlCVKmguS5vHn1Z9AQT/xohuc7cwmXrcZb3sP0zkP8wbhqkRu9auoov5YvDVAGlYU+l1
Cft5m8FN/wULdWo5G1D0dA11cCv0/Wm9u0LSKgtah1XIPs9l9xgI8hDvx5asp7GNTtdsBRofdTxe
+Qsul+/fdk7+g6vECOZVyYs2ED01KXXt+42Qyn8OWtzvjRC21LPNcyR91c2ucXR35CjG1kT+5xuQ
JzHlmjc6IuYyf418bIzBSpSBdeK35pw7Dbggal0Qd7V/X+awuzBa9GRH94fAW/50ZrV9ippZgBia
EMJeSD4nyG6eOoQGO2YEFXuBpJgoBzdX3bl0/uNVE2gLMy0+rBW9PUsMExHUl9pq5PqXh00UtxYG
xzu3UVETnbAnGK/G3eKHSkLLauktsKwWf6SUNahoQCUX8sXN9iOzFLLB+Xbs8QxH2KS3+B9GZ8/Q
FG98u/vYYdX5AX9BBejLmDa0qxud/Fpxula0nbe0nrTOrhjdjH9SHkXgLv/Yb0emCRZ0LoS5kFcz
V5/Y3xumpzAnLEtNKl2QAFE0P2XeJjYaDlC+kI2iUB7Qpg70ASD1ze4BO14Ju/H8Jy3Sb1gG/6F0
yKrh1yQ8nCNoDoTObzH+iI7QARWKiAFEG7InYrKufEoLJM6wIuvE6f7DQqrpSpnx5Wwb15QKEUdZ
0V1n46+VhXgwdf2W0ESciLLXTl10IsYYCbB3SiRgVZLWz8ems3n3chD37EbwsvlXgWjwbsjpSegv
f6Wn8OH01z9SsSa14HgdAiwSbkPmkFfISvejU5aGjQl3aU7hrrHqMJ5+dxiISZG/2zZkFBAmWOe+
zBJCdiVgsyhoW8qFEC091nRitbiwB4z29pYBWGhlyjUinPUwLBYI5LC+p8ixPYPAl4WyKtctWhKh
EX86IbDdG4kvyVHnYgBEnlR9kuB1TZoX6PgSmHXGXOHdpxHQbbO/LdGtX2dOQCnMOVTUBELRvso/
NJ+2mAPH1/jNKhxKlFLba8FC4Heli6tPgSycZXN8fa5uToal6LWW5O7B8MoV9qqNI+n1UdkrF5qY
aYbS5/CFfGBofGc+PjYLerqDN3Jr7w8krvPHASmWI9pGEpy1/31qxnPBnI3BMwidHSqYL7+BahoH
a0/xR5I6kXwWzcUZUMGPAclZJhT2JDvLrAjWQOT/sKlRJffwzi/lO/uENt5G+R91MovDVBe1N2zK
2nTH+bffkiD/y+CM+lCsJ0sM4EltVf4XKy09gdKkE22D7QuzelSAOeCwBAJ2+GLVrfXhOZkayWhB
u/94rd/wCINTShavApfO+5+KSq+RJ/TDKJwBevEy4LcjCjAPeoitY28ePSEriwdRs/dYXJuwodQ7
7bxwa7/qT6li+89QgHljF+ddluhShIjPNBoT/vHFPOqC1UQIlrXvcPG4qkMqTtkaFXJScvgtHVDF
D1Ff4ZoZods5oXNOzlw7SiEZdUw3eGc0sef9ADEolA3J1Xzta6R2EYbH/IqDz8giBpR/EOTcpvdh
fMWcTdchsp1pRNy9TkOwDXndDbhIOEljJ1mi1Si10xa5r1oLyw+8+3rwZ2ezXTUay0Rw4oFxl/7S
Rqpf08rZtpib+3sN1opOLwg7QCLsscHZvS6zrZcHYHVhSEhMgT9zrVO/aXBOAygrKTZJeCchHO7Z
SKOay5AsNsvtPoRrsVglGVyQjcwflV8quP9GnRnqLd4H9E7l8KQdZEu01CzWiS1fckwCuHpHmprp
Gq7UcJJq8yQZvx3gaAg2KF9enKpDcYZO66W9rQfynR3s/n9tvMRRyU+AzbQbom+0PctlBVZEJh/N
9Mz3/K+3a/cKXsmld/Q5n9uNRdO4cG3071BLZ8CeNpqxVpDVtH25jttJYkXZwXgVKPfzCzDgUCsY
wwnJFKQEp8v1oRSdIH0vBJh1KHelf+tZ0IS/cAc/TC5ymRElyI2iuZHmT4YXvMy/d1Ki8gLrgVuv
BsOePt0hKp+jspSkdDgNI2iL2jtMvoC4aBkpSHoxiKy9A2y91hQHv9qTf4gJ45aZIu+k9sqy85z0
I1cGvfDg+nMRdZ1xErV32LzfH1R9/Ms2+srDujVpDtlg7jmfVzzVwya0UMfZ8GdWt3Yy1IKEiBzB
SKPiKhr61PwQZ2YI3/cL/S0sOFrDRLyy3vB+U5VGYiDvfkvTuYuzHWJsqn45BEvXVyPcjVDkAy+Q
Zvd0qXEs1lWnOmF+3U42kT+EHtcNxB2IaBClO3Fmu1GBBlxO6/dBmREt3SDCBkgb6qYIERuR04oB
V9FtYeK/t52DS+YBToQ3L3kyu4Zn0X2cV7qNxlHZ2ztXm0cynhFtxvj3yYnj7dy77/YZLeQ7Iiw9
QcMcKkXhrnPpfzjIB8+jdEGB9ZrAaRUFRN2HDDFVwfUTkAsb2P48okVzXg3kVDnpZwBRrL3sZS8O
Z0D0bh0G5Rbp/Eu8OOPuBjW9Iv/RU9/ZgehwlFZvB6enKQwQ1Dh/IHMh43kPaU6ujsiBZqgMPZuE
jVRP8XDd2JkHdF+58jQ4EyanZiHw5HYn1gHJO00Q5bcwlLGrCXxl4xPUE/RevOaK0t7bAj4myGzo
gZYdXRvTEOvuBxtzLNIDEJa9Ebt6bzYrSkXHZ42FTN2YmAz/HqyGdCIPocPyBxnXfj6q3pPS4Fqg
OsAIosRMtpGNXZMfoXCKWocWkS5fDbzAHV9uJNZPJuXnPrv7ohggZU2hrRuikWHXzU03ctaqRpkj
nEZ/BC8wtZFqXmW6tdhuvxcZ1UNfgssiY/9+BzvhztBahBya2GJVLjOk9uGdidGH0d8ih55YZh+d
+AudVLEAZMASQA8KA2ulcKSomXvcRPZdiP5ffYk8UB7hGSzS2+4+GN49p9ReFuy7H0Evm8HHSiv4
oizeH+nqX3ibh9onsc3ERhys+yFehTbRR4W4Py6iUZv/uTsD1mw8k9DurtKtvgvgb3z35n6HNrrU
XiB2n7OBt2z74jz/x0aKgPWiNk4Q4cc6h7K2BHnjR+Jj/bEsg+4HWkZG8Jkr2TGvOt/s5vx1M7gM
8fpkFhbpEm4+bfAFTQM+yDcL4/P7fOYH+5y2/030iJRcZ1FSXawi6HklAzVIXZgXOIkzugyxLR5S
7wRx1m5+4CMc2ycPBGA74FtCkVaRkUahGIKDlh7EEJY+fYLEk28Cb2PqtkGy7qE3ccQrzSWdNIeM
nTX5JPqb8rER4FJ9vToA0N8QRW9AP9qXkr2nMg4hpPJyL1FfaMFLGFUWunimy2DXGYXl5DKeA+dp
jHblUg1VmhdErHkpNh2Vw8M0pFaRk3wPk7h7NTYB8CLkE02ThFv7Ed+KNtL+HH8XF8wDWBYNqKCS
L+Th9cveeE1X7t3v+T6q80UbF6/4VrgcghHlvti1ZgQtzc7zjKVWhnat1mI0Thwio3BcLmiZSoTo
pNow1f0iM1ro8iEnmLYpwuHDGc5DgdsLVpEMLf+zXKQT9WKZDZRX5+ITSqcrTXv6pghqSNnmA5Mc
RcJtH4Gjv+3Nz9QajPUzLzMMNB66vLxl3jSR9/cyGQlBwOhqpQB1JIAcoLbRSoX4pOXPWCmhr93s
rYHZcpu+Wd68pepQcZMccLq+0w9oaSyrcA03maC34k5P+IGiNjn9WtumWC+WNy07c31nEQcL25kp
0radLmcwbXplBniZvE7jSS4FQPLewMHcbwVZlL0OWbaWKIlUgoXAGzi+YOE6YXxwzZrujhFqVBCg
f9prZMXhy66ZGDqCIdQ5mE/tfTwJ3iGR4T8LXtkV8kPGN82taLMprvVw3NVX0qGHWOgP5s0JGLFs
GUcGJGZFFXv6zZaqhiY+XnNk0UJ55K82vOHNx+xmTdh9FZ6dKpI+Ib6J1ROri1VPkK+w5jOXz+UV
XfS9YerS/2D7vWoKcoxGd+DasN+A+GfOMmdkSbUzIsWKu51JgkaA6jCdkd9qPUDkwSAEkMx2+11/
Jmdz6q00A/SJqk4uSKceO1SYQ6kkoMjnBBnu/u02cmVT7LELCOKRRWngR9Qsqb8cCkrv1Bh7HaVG
KZrWArkpLOYnKDNcgUL0L1scpzUUdnSnNVTkwXcGi7pKLRhBsg17Zq/X16Q3AWkWgom2PlY72UlA
tEdLr27i9Wyg6Jk01tckBctXHEQF4+rtxXWwI80j+nrT1yoGhJMVT7OdXFxo3IlzrcfThtdhS/ds
1aIhjvZnZnI8QJo1HZkODNotclPgCu1pG/71Q5GAAF8KvwnKR7T68YuCTJQ6lay+2FIXqoSjK91K
zo1znHOfx5TruEU4dCk67+IMVYP0Vs3zjY2PVom5p1YAG+5d801fhDYx6O29QBp+ifUoS8MwAw1D
nat8wf4VZrDuNw8fDpgvrG5/fWS+YZ4Ek7qkFeKhT7rk+UamFBU9bAuzhYEEum/1oBB5ps5IcraV
XIkT1ytGYg+w0tay0d4KrBgyVbrxVGmO9o4LBFCsU+5kJ5jpEtBiMlqx8rT3jW2XwPABHkepxyoN
uYEoqxWP/K2T7CExnRK18pbNRHbZZxdHRWwNHs5yTm6e9CowMc+X1SoYElOneSgTrYN2B+Am6qly
JzdyOoE4Z2ivyt5v/JTZIS5CjLWDCwJFLO0TO4QTAzyYN12sd2qw5MOL4lFLjyiuGuK6jXwpBDpc
5lbdCKr84mCD6meSPPmWezLf67l+P0bG5jh1sciav48IWC5L0Qm8PFzmqcyVeaQkEN9DW7drtRhs
mreDs1qZwKmMJk5y09kewm34Zxq8FEbIP8Yqd+H94S0qob7063LjBb8zJsxwMO2KnuNn/pcYMmF1
wIkf1fjKo0nVwTwAqfBngeqKsWUdv2pdoU2CFS7w5dKR3TyZrX60F5rQ6FiVykZjCPu0cPs9eIas
AnKdqzGTlAGmykRtY7EHZbJ/Ohk7evS8sw0TxOd/c0MTOonGKmRlLlba/xUJm/am4b9OUnKEImF0
s5liC8DooEQ2jaefZNowNps6oEEwMaXEZfwDCz/IuL09zgtsRu/n6CTglR8ZjXAE6JW01Hl3pZeP
xF7JsQI/N8X48FCjeFpiJT9hxKpJlwEJmqy9PyPFCto7snAO8wMjh9Z/EjOKS6Zz9F+oM/wGTLf6
zkZjurv93lYT/nQu4xL7SE1WxcSTTk6fwr9s0u3unK6hW+qgY2dpAGjYmdaftVHDQh0GBW5LQQO6
5w9ftOnx7i0OwZJJOjV8K2qlFF1WzX1oRmKtWQ0dEHgZbzJVRFVDG4hjR0QfTv2MwIDfOpO0tqYD
OIceEr0nVm3wkL6+j5M6KyWe06HcFc8Jzt3dSnkWOWfC7a6o4DMHoZjaAcW/OohtrZkIBda6l4yN
VEjcGb1V1RoBmuGFDwpk47wMiqz0Nr9FNjYK4eTZ6zlMdGOu5m4Z/dA7vJzvnoDo2kfz41dZbtT/
2Bm1Qy09YlzO1f5F7eTds5oM3S61j6bsFngKsrYUKb09eFie+0Z1tm6dypN1zYmrIKKYQuokSQot
fuCw/D4jWiv9W/1GPJx7C3D8ztxYOsuePsks6UMqcowGmD1EZN9CMsYQbdcGmGLN500BJ+i8C1ve
Mj/BwCGaO2I0jAPNUtubUGuh4hHQsf6cII28b/V5A7s8BUrzX2sCWMC2a6XfD3oFZkQRftEsSIti
CBKRCtZ/JqWVTBTt+7eLEUZYZQ46EiSb6HjAnKHUdnRlXkUQitXmEXlWNRlQe03PeaCqFQUt+Uik
Ur5V8+kPBl+vRgCG6bsu0Gj24o+n35cNTPJykOA3YJX5x2eDaiext1+UycOOj9J1ib7vSHRmZqMD
rzHDg/skNazP9yEtvVq6VG9cigiZrqm+/IiQZyvQ2HZdVg3hq168mV+NX+9+CmCpwMEOGj6nwyMr
NBpexZUxEEZv4p9v5pvwzny/vJUrXDJji2ArlsaTh5QzyVJOfXIA7juQOaBIJP7xGoi9iT0543wn
5Z+9Vi7YUVxVSITWUSA0JJ2z1C/Hw2WCl2kGHpkw6GKwMbeFP9Cx2o9+IIP0IUeih2MqEIKUe9js
O8UGm8ng4XU21FNYcOb2xgjKW6UCAMtLXCruSqHx0WvPgBuTwysiDt1mHOikPZqmIVBRbs5VVf7e
4oC5V4+Q1zXdjLiuXlF3y3DmsVKhjyC7MHROaa/0i2cDsxlhyTv/a89BhBtBqlf9IrDU/H7zbfuT
6Y+pmG08BAl8zXQoWAkQ9dvy9ovPQMDPZPHbV0Io42kFRXeAAm+JxLd1QaQBRH6x7Azk7wlTYPB9
nyal1+4i8XZMiAl3Cps1aJCtm0tS/Y5ULWoGRiepl/0sb1taSL00r4qtlo3BC3eLRWRCDWGjnORI
feNeUOVVdPGfR8quX2tQrJzSXBF18r84sMVReGXvEgy/DN5YKhiyqpPg9P67JwTXyc0vICAuwv2J
A4dqhvSw07vW+VNQp+4/Dpz4hCQluaIAO77sF0nMu7EoHAuOLZvDhSv4Ivm0Zp/GKmO3P6EbVf7w
QG62j/VGNMZMVVWphBFEx1YSxI1+iawkmMHCRATHMchIb/8KfgRWboll6p++3VBVj2jC0nEHhOPq
0sp7kRg/EfSpmsCEbWasSz4tf5BpSD7KrhyC7uAICc0knFCVGa8rqGNb0r3jPGvnUmQTczEgknx4
ocDPZM10dvavy0EtMoc9icY5aefTyUSx1aH5rb3ho3234mqmiMu9KmSZDIls8p2/YLGbusroN2By
anslEUhVH3aZeh5K9E4o3bxhXPclhKUbp7EnALjzJxfLMUHGil2VqGVGqv0gR6qrPJPxnXUoPbgy
HeZFIAyELlF2V6IfMD0dmo9cFn66HgTX0zc8iwBtJUT3cYj7TAq3t0d8NTLgh+PyreAds4Hhw1DO
cGspwwi+V4tAhJAQM6psOEu18CJ/vuK4lTHXzEFR4rACgtdnUTE7aE08kdw+yesWt/AC+qpJ6fRD
j65DyBhfWiq1c7FKfdqK52m892YTai7fgWF1o7K5ZOyYZXMCAAUwTS626K1HQ7W8xpQv91RdhB20
b3E6YSk8sSXV/m/LuXCPbnx/K2u1HXOMOnJ+iSVq6zPaQytEfXxaETT1lMZdbFPJJT4yaTt04qbt
hTDEM8vb11+tLiPc/FPySxtRX6muobF91/Eq+Rqo3jlBy57ZR8FHORY2BpyqxcBBOlbVlFZHt/v7
+qBeyqyCAD3H6ADNbMZkBgzo3NC9s9o3beY9UFVTwVqorJ3IrToz0t+K4WXGc+dyUGBpzCp0jspt
7MeTtE08zlpsGcX+19iDcXUN2Pt+KLkIO2TiT5VrdCTFzV6aWRxcCqLEC815NSwD3+MDHNn9tPBn
riGKq1Mz8EyOnOUpffhjT9sOeseWqFrqTvCX5RlTG2dLhK0om4ZSSBEXVb8GIGQryWN8f9I6ryre
D5hFEaOlojkALmslBLCAMtItj4dJfMn0vYxZPl+gPlEUH3QjAJuVFRKh9cPf8yPMz98YRSHJlyu1
BiJlgntCjUqLg6difgoiBq+G0mj8oGrqi2iwAehkwuo7s6fwaUZi2N/yy5dxZsg3aWcUGdwQOkXI
rT0wjA8UhaAQjxaauPnggjpEbEqyrmWErK1QhvqU7VA4Ejnyul3BgBakU8A21qkr3AyA0Ns2IVl/
roenWAe7tz3TIKx2b/NWGAPfLc0tUbSyIQLgxumxgbnWs27l07iTRAyIymPDJvTtRpaRAOwAax0C
Bj4HsZb71sEEFL26NpLh44eq/hnlK6GWw8wTZqSGEv7FJR0ajKRV0OyaMMOb4TEAXnDLbllc9/NE
nRgHoJnYYgutxU0lPCX3it6qPZtPGmnaF173UWnxF7BQ7U/JPeB1V/Z0cOa9viUImMjwVlUyOa0v
Zj+LwN0x1SDE0xhrgE+1zg9SawzUCpOBuWsCFgl9/IWAJn1gCgN2dCCpqFUHm7IMempQC/V1PBS1
J/juV7w5hKddNe5POUkTEDjDIfFNIUqzjYgEn+53ZdNuxH2GonQ2fY12XyWQQix373v1lXugTmrI
3tt3KoEy3V98I+JrTY/eBsU8oXiC/IRIRjq30zprONmddeLdBMvXlX0/TozLoVVN7Z+QTeZunqiu
fVIIsiliMo32Li5LfIkT47/Z4F6elAfIDyK4M+GsMeI2tTzGs9tIDJMYgVVBQMZLjKhjDcunf0S2
KXT4FuW8hTiopN4arv1/F3mrNtdrw77Gy9TO6NCK2WWppTeAQtjLa79YEj/lHNmvv5QvcBjRMc+d
1Pg8zymvwbq71BTMXDWKUDv5vArZY/FXqIRvdXt8c+XXhEm6bnWo43UV4LS3p9mkxC78jNK5D3E/
wRai+WKkTKJ7euWNdA6e/6tIlYonbibzR92Z+jV28SNpIYNU50flsf4b/TDOw4gPV+jJkETGzovJ
qsXdpmJ0ORzPBa5wNoUhxVMSdzdpBOAOtl5fIc+RH1LZ/jAjG9kR4AT5TQ+oreLL0NY+UlhbXgRV
vF1tbjzmLpz3O+v5dja7UQMvkC/1VTN90SUXLj7r7LrJf9wl1RTlIfXFV5hQ0AyTqLIK+Py0s8hR
0O6l6sa+4BRP8LutIhcCXAq851ovdpjY6COB3RmWAdYHVSJMboPl+J97LhGF23pYc4IZfFMpRgWj
1+i2U3UMyRfpSwrE2Tlb+ZeKltTX3jRqNtLmgQZghDRU6U7BgH2olO2rU7uqYvzews30vzj10yQs
QmDfVZemwkKLkgFfNdFUxuT69K+yehOErGwVPFvQ1JPHZKVDVCdNw4H2X2dwhpzTcP/aduymOePv
PB0kACKe+N+rwMrsGnaeLhuFY4F90Edckto14kOqJsZcxCh5OowjEvcIJgbqmrJvo0bC7yDTSact
nhjkb0YvoctbP2CT149mPgeS57WNgEpOtMBpYM+GRE8PG84nBTaEBhaZ1zfVpPSqN6ecbJVSB4my
yroUbp8pDHw6DeN/qtLwIah0WMDPtMNB/zrH+NJQy3/tjDEKqvGmoTNA2/Yyb/RQWKOeVXfpKWJD
/Ce/1hYt5amxqJRpG3pVJlnZQVuqAp3F93Xd+MjkAtIylaFj2OuFbX60v0ZyllVD9A+0/ZBfvmiH
CTHyB2ugwldzpXktzJMGUuzwPdlYiHMsL7IQs/nTlQlu/HHNOY0yZwK8/cM986rRl8iScczlWNxn
26ZO7t5QVpAs17E+I1TnKw3L/cikiMmcTmmNY9kABPLf+2R4AfYP2HMUUrYoLbXnqASjVfkvJROl
UiEXNbLYySwiJ03zrRxe5hbSkuUeVDw/2rdT86as7Ok4cQF3qOZnJLuif4eTgLr6LoZ/Wxj4HsIC
cT86TOmktjxrAOyPz22/0AL8reBypxrp1HcgMGLa/JwEBrudxfV8yBN6OMUDZzaLYfX3TloQZdPI
VYZEJ5Mtq4Kea2bKKAsd6sgZXDx1P26WE/IdPQJDDi6pFxT0qJF6Z8em9I79BWBMkL3iJGguP2vG
qBuBmnCos6RL+W4/zgvSCHcwSFIRKhBoffjOyW+AuV5RaWTqPo7zlFf1iNhIV8NE+Hypg0uSab0m
yZYXBDX9wQ5FLxaJyYIZAPdAChv3xZ1OhMX+de+8HeymxmtZXDlt0JE3RT7mCbZDIKpdP3EyCr8E
IHNEt/McIDRA+RQ/L5zshkuWeS8C4zQZm6XC+a/7j2AXGVg3zBHOZvMg7oLiX8Co+IF3xYlN9PMs
hJSUT1Z4onnEYc5xzcMm1pIJp8B1nGhkvcIcSzNMvkRbPHi/OtUWtTqI90yRBYKBrtqN6btBweBk
koBetRQqrWXKF3kGLLj6BHKK3petFr0Iukr2TGOwB+1fQhod8JBWzjx2FFPbTm8ToufV7vGvkINl
LdMSFgVOe4n1geSKhVlcf1rxANKPYa2nIDjfppxJn4ksq3oeBrAjyDEupJndwKhYwUkFa7IpxdRP
a0BdNkH+Ae0d3z75XRzAVToEEzLrNhgrPi9px6WHwr5VW/SQ85NYJWW413tolWLL/3qZqD1nuIHn
zCQTqeZVGDAsIg/NqBJbMmG4xsql0hRmtPk59CoDoK9SCRPS7g+vjwAYyLvXAFfMtfyLa/2nNCYW
Gi154IJyrQxBie9gcIEn7t1zYWgbkNQTHPCQokiDf98DrJqkh4bHaW1H+oU79x5tockL3SmHVIPo
tLp79bv9BDdTI5ZSac/JPD+cWtUJ+LlD5IAL1B5svaZR+gu+uzqewat8/Csl4qUhOum/cc8vMUCy
Kxv/xmIqzu++a5iASVGMxq16V3vjW9428xhQRhMFB/+kq9RbRSN4Cob9aXyNLBdpu8tnEGcAyG9J
+uMCqSVROb33dbdQ/QG71vkM/q4GaTgtnQzJzJ9d33vmksyqdGs5oWAZ9zQSZ1sPflq3wUA3MSLA
83NHvU5U/J+zzaxdEigGFLMTuk+Wp23MYRCDgBMMgdUrJ3CpSfifrqaz6hpyw7CqL7IBor4C85/J
I3P4CCpY05MuS/j2PiOADRjNbAce/5xLxfWR5/KCw2xQauqkJCMytYABSCt2B2VdE2C5jkiarmAG
YYEKBP2N/cMG0drOOO/N9p8H1idm5A+FvW7EILFzbfVKI2JP6ko6HoUeZBJsk17Tehw38Gi7edyf
T7dHAC+9Da436uW8xmgXapTqnaVe89x23UftpITa9abLhmtAMj1DYMiezlj3DWjDRf5MoJ6H9rUa
taE4LanRaT5xbkR5AaQQt1aWbjYXIlYVZSTuWmzOJiwQaGoHanGSPd6vAI72ISGTIksZ9P90T6sm
CuQMRqI2abil+GRnt80z4+NpC5ilwwQkF+KPJuLhe3YZZyuJU2Rbav4ej5ofdcNMH31YGjewgXCa
8h0vQ62z/mXmdHQsWiOpTv6K+V56NHj+gkud7ZQhVkjgtM+oNiLqUYZUNAwz3R29ILWZPM5akn2H
bWldfmzIY2rYFIygBJH4J3F1M+YwZL+NC5ROj7v5zhMguPTn3J7rNijNB2F0GoPgBS1iqih0CQ32
xBbgiaiFbj3Q7Ar2gqsI1ZQdixYEFdtXwPLsP3mla+CEb/tFN7AP//Mi0IKR0zHXPj7RLcMu6sAy
h4d6kKAlv0lTCVndD9mXO0ETk5ZdimmKaLzp3hd8qfa1n/eR9mev9KsypIE98EG9YznPFw899v5x
jbpV0P0jcJ4MhMNFVMunA51GzU/9yQgUzin8jcCm7qWn8fhJX5jz23cZt5eEwITFerza5cXVvzsg
eYOqo0PcklAlG15I7E+icHSoWXf2RB5F47z+sbsrZRVpEYFwhbQdCDJtfPTBua44ITiBhhH9ILT0
NS2Rbwn+9Eo5HjPuKvqp1Oy1/GpkktVg9EZVhRP3NuoaBGWzVW4MB99nSVAw2hVKjdNjBZsnCtQa
uXayR7KU6yDgq8m0ZRtPMC8HTUY9WB1EpiGT2jbh4S6S9DjZCFqaBi81PVVD/WTuvHiBixiucDnN
Ci2snEJ2w3tfm+bjyW7U4sxU6BwIfUUbq+mJ30Wqg9fUPWD8U0rWbRqGKFlpx5OSbJlXpZ6fwd9p
M79fJ2L7wMgn/aTa+0ZRpp5zC5BQ3Bxez+akgohpze7iIVVteLG5WT27kuL/FNcl4KWrFqt4boWb
FVmoi2zUo3WkTaEscXZdoioPWzz1qUAxWJuZS5oo+hMLL5Mf8JPIFQFhBP7G0qmeNtHUUhnOXcDc
8fRyevP8H65Q8Jc8dxd0RARRA/NSiegunhaPf9Wn8FepPccPAQOToG/vdbaiLwcOzruF346VsMGi
zxDNEmrrOJSAoYk59YQMgjhhmmquG7prqff+pO+2oYVGYiqmKhyKaHlFmmyCVPigpF05VOHlZXk4
UYpZeOrFsGwjuaO2YvZGHcXZx3EPfsykIZWRJJewz1LO9J6cDY7xGg+dUU0Q2jLO2rh404CqH0h/
SHb/Glf/hTz/vfIheMoyJZAPYVPWncBvoPw9UNBz2HAqf37goUsnuDi3//weoyeAE5ctcNQtoTkS
CUUmxvTRTKddyeY2J57FJ7sAMg1hmm9kq29KbBHJt8gglWnvtYd3NWMDwBfwVWBplKs0TpLlXOPN
NKEio4LWKLcNgxyDt4h5zNeOXVsCx6mV43rV5JF3/aRS9DtjleO1fmn6TsXYyiK2CKYmpzBHaiZX
x60/pdWNSn2squgWE53Rk8ONKMmqPebrUKJA70l0GviPhGt4NwEjuSIsY30U1VD4iTFA2MkfqEJV
hu4h23kFwLtocOo8BEmBtrmTHW5Mpl09tV+mJ/dkr9DcpKtKI71Ys3EaHBTSGo/YF/f8+hDtj6S9
+1rhUZNydJka8F90uHuAS2PCRYwqGGlyRCo/39WEiOAGRmrRZQb2ca/GfRjcaZ2boZJyWtvMFuzy
Tf60G88asn1jtGJWNtyJB1ieMVfDsSDLWEOob+LVsIevxaXObJKYYcZZ/G5JxnNyayCFBo+gSwxH
wn9fWo6mFHRTiuq+qymyxUAnD6OSJs1ZnbsgklVWP+0kaUVwfWbFu757hk5jTCAvhV5GB6lowhO5
DsXXjQ1vAU904vT0CIysdJycdcZtawouFVEIZWnJ6ObB0gWGWefNWWwK6isScGn3zSW1KLSK08qS
9YlrazxyLH1gNPzAJ+aOM+UZ5Hc350ah2CPYaJGC3Wf4zD4WESiHUAFvcG04X3rOI7jEE0STceZZ
QZmTTmO9iRSr2Bdw771E73clud+odiWonUY7pIk5GcVXOK0f6BXpMNHHPcMPzD5WcsuqVfc4K1q6
3SAz9VuMV0SiU7cGMdBwdFBnC5at+JbkLGVdhf/iqqJusPUq7gWnFRQ8pokVTqHl1HerOBm4ZotX
hqg0rkkirDXKaxoEHClhmE36x8LF87A0YY7cPFF8d260vfrr71xR7D9TvNam/u6ffR+5DvH+x8s1
nHpw4cZ0OXbbfdojWEyZUBTraeXoVgK0qEe5ZWO6MRnNJBsrNBWRWnm7vn2LSQH5zbypTPYrWfYR
6iSHxFgdXfT63a0zJMGElG4zo3QkdRXn5jDivJNl4ffooQsA30nvcDxHNCYlnS+AT2IaFBv8KsU8
MjeOqLRF0pQybvTwT5lh3hjhEg653A6vA6N5E2tmMqtFx3ywssQ38g53FMKlixBccbAPJjFJ7UQn
HZPOJnLBJL+q72ykIwqB6WurHy0v/7OCmGjE/uT6oCglgR1QKXDlNPaL4tmBKKPsXfZJutf0hbHL
7Pl56LdrWjzJe7cMow/YY2zhxXmQclakG1ixipjcekfc1q8JH71HQ2Zi/BAMD93jKxcG0TuETiYy
Dwd8yDwM+gMxhbwa1JHlXssVKwaYPIxtVqGD4zqIF2dldjuWdFe1G8lSfBFgyDDVV/tL/VwCpgKg
pOsmSaUlmbzDCusCtvE5L4DwRqsLv5L9u5T5SbWqWOaeyXTSvgR1Wcfwl/p0in3A7dEYLHYraNN5
C2tx2MWnYYkWqwUp/SVXVtiBuxhJ2P1j+6anmvIMa/JM19Go+lQQsZT+uX2VPM2FOvAEaP5Y6RdZ
+iQtB/b1G4T26JCNSZGA5ySBYcdrMdAduk2vImvplFSuiF7gXmeN7x16v4fE+qmAtrAXgV+3SIHm
PIBzSqCFO2g5xtUHzwYMjRVFwNBf3H3yXFwQSlXAxpGIAjcfPrWG0OFBm9buy7go6hGN6xAA4VWu
cHjhQ8Oc3uaGpqDK9z26i1rozbEb/bAVVFmsw5+pmSnr/pEt2HDs92GSiPhEdn1kjWVcoYJrN1v4
bI/yNZOPu+tmnxYS7q2X7pShKdw2JwUujIadj9Dchn4F0vgfdt3yVa2uyv3uiZam4pbgQIFCHhec
dBkUf7uzKw2wvhH50TjFeFMbLzzOFAtFisoSgRdQgCW4idtbj9m5+4LS84Tc5KIS5srnBXYWwF74
+8NFY8Bk8MKc3oXuZb63gGcNSH+6eEZnyE6I4og/oZxegddAUojYVIESqaoykY8KI8B19U/2xhij
8BgwVGCSdYOi6ZWRNyC0V/ZpXzgL9FJhNW98Wbo+ZRlqzOLo3S414u4lUyXBPxifEZAe/bvoeyUX
J20SO8XSgxgH1dz7h8CjgemNLO7OAuhXeshFtNJFHtb83jMdgCdDzYqiMQGLZ8+jE3mTaU1TrRdH
Y6v4734gJGBTEOhoyzGd1Kgnm5nUj+NUxN4QvlxOzEogIO0Z1BBmBzku6TD8ZkarrOHbGjW8W/eV
ETPWhyRXdsJTuPamvfA8Pn6liBlGxJIHUwcJ5DN0WetaoX6BtLlOvb1s4GKhMxP7mODTVIMLW5ak
UqCAjJ8ufTOwY53a58qlqT7BK9GuF4BRTIceFhJwfIpjtHypxhC713nsmRI1b6STfpFRniCy3X1l
50sF3eLPz5J62X7L/enNJI/ExcReswmWGWKji8ZVbdmvCpd6j+o7cN/l4MH3L2mk7vccp+8Dh9Ts
6nVqCIpn06Aa0buUoPhMJ+zNaeekQ921asC0knt0vPXdPvgXTphWz0TInKZ7IGo2t496BbGEWDKU
+c3sOvjszntKkM1GxGc+pOyIT7LfUOUJNlcguusryS0HHsjHZQIf+4q1Uf3kI7yQanZYMy1ayKGn
A5X8PXx6EIk0/Pd35VZjOfd9hvFN6R7gFtf0ji1Ru4VrA2Dp3lfIau5IM3EUB5PdTfBjfNOk4rRe
uPpeb+6qMzS6373Rd3oz7RWOJH1/nMgM2TXAQfGptWYxVzS42xW5nEBYZicUoyvva/F29adavNK3
3vNt9nvWqrdS13poyTrsjqEyxkDzG+/fiWEpNAV7jWJv5OrJen8Lkl+0dk/zbdmgY8rIvVdFgMmE
PV/VueCaAVXb4ZYiRZech4JEL61kQr0xo403uBHKDrXMxRW4Jve5vWvYHYzJrKKPIYS27O0apmUm
qAONYpXllc06DyB1FLwpcdtyJvuH/QPeRFZupS5sCrHOneIV4erXSqSSLTgXwg6yUd3oSWoP3+9E
UMW0bmrrbjsH8iKCZa8Xqd4tDCrjUjdV7awmBK3d0GbKwzR9pnz6M4MQOegGQ6L959RE3dxzHf3o
OHukPzwNHnPHC7RLMwWR7IaJLEhaQxkgGpm1orQbXNqYKsKzvp3CmI3lMpcJzpIvBpgaOORQATft
XIj1AIJGKM2MasALcWCaJbO2t7R3bNEKjvw+SJNWlKhWlpolN2e2sD8ZI9ndOq4vChjFScFPmkV5
wmownrQIkH+88dPYkUPSKkh8+zMlgBKIC2perImql7qQL0DXFUUo7L8m2m3HkzW2RCjFI8GuJTH5
yDrmEojqba2VV7fdQ1RfFNX2F+cY6xoTGon5cfRm9WKlZj1D5lJX26Ve4wbNqQdL9D5TfzgEiL0O
k4ikAlPjcRUttOIhfsFIEntFjgOjtgJMpgkv6emUKW26VsYpEcwS4Btd6VhgWA3f6x8BKeRzUJ1b
3uTu+r1Bwtysr9BbZF85k5S4ut6k/Pnr9wtiryWb2D5Hssh7UX41WM8mmV984mXlXFqkt6k4wPT/
eTiBmgWyp9wsqYUa1XJPPE84mfk8EBs4VkN+HCNNgBbvwBgkC39yZJ1H4y2rGH4KHacrKL6ey4ED
wtUXpxFwN7JLXrtvfZiiZMmhi7pS3hNXKun2v268Jw6UTR5MAowVyKY5qyjqvSPiYQL8E3TDFcC5
c/16SsVMys3YCW9RjUXYYJPAPHbfWrM9DVbCpl9TgGw8RA5kUoTdYkMOwZ7enLrB143yfylUg2VO
ssHniPaxH+AuwqyPDusw0Xg+vzhwVWIy5TS9OaPb/MUdKdLgkqTuWcIhd+9fKNiUiIzY+hCow16R
kqdY1qBSlc8FWr8tSQm/rVQAt0Yd4zryLsi67PU9QyPVGT4zg8A4/C9fqTV3amxwX/5mhsEo9Vi7
feBLmBiTEMaFckUMFD09Tsbl3/+O7gBJSrfslKbkfZ5ZeLVXPzsj3nGrTeKBFrGnhnbWMo8AACqP
9HXEzfqoDV63uLmHN/RRqx9PpenN9wsTYRQ2XFJ6xgOJOAxLbUCqxyw29/ReD8IIvAC7rtJ3/Ze4
sY4l/ctN9B2kqrktHf70OdZtDpijnLOy2x5r4eS5j/MPsipyhXznNWlX48oRbZI7d+parF5TEpJm
L0YVt6SP1Is+LcYTBztxCMglvcl92wRJy9athD9Z73c3nydS4HZzy/kQm+I3SWrEZDp23R3H/c/F
pgsfLsI4iZY91bfVF4pDAhE3W5IektS3xF5GT+VEOlutYQlGQvHf5Nrp7qNejTVYAV7f/YVUff63
c+QXOdleipyVAb4ibs2IV54c6npRS8tDx4FprfjjdKwL7ZREM4X99k2HqnxkI3qjUXm9/6oVkuMI
+EXWNFtiUds7EdCQkFUdWVBxz3Iy1YXh07K6kWxQz6ltbQ5OaXiGsT1yjfEwi6lorBxT2/VnJaay
GZq6vQiWSuoc1PyT94fDB5wUWOzRGUwvX1cQfLIPO3E+HBYxofsrxkmMU9BQMKprSElKPSx8Q0Dd
YSN+4BlF5EeDry1CL1aLaGOv+rDRjtpoMccBiTuJvREOTMChcN2NbcSI06t/Hvx8EpyCuTmH6Cgs
eE6r6mVaZ/GnjXoF37jOMu3DB/pEG/UrU+5oA+mtxVJ6zlamHooPWY9GGgxSWI+mAYnRwL91zcVu
l3aCJq6KDE6VWGhy1DEK6j3o9/rhOGCtbQc3YO3McBH4jOMz/AvkJsaho8x4KeCg/m8A+uTpTE7v
xXtw++V1qu1HNGFGy7NGFXaQV/TLVbZi033nBloY2jbiZRaNm6ElF5/bXRun51aLN8KqT22gpmKI
VPl/enDUvQdH3amG7gu0d3JvjcakGBkX4um1piMnZ0qP41awHT4SBf0g01z4JJ7bdERzNRFMMjiQ
4U7spSdyjLd5IopPni9elt3U7vxUCDDP2UwgERYoH9jd/lVFjV3dLCdkb8B5KLfx86G3bXd0Po1l
X4Uvvz4Sj2uuXQqQ2JjS3YbVBSJoPKkNrULUJvH6OjScYYSZTmHaOE9toFiwfF/btnZEw3Cr95hV
SLyzxxFVm7tsLZFS+w4Ic0K1Tq2wsWV+ZkV3DH3WMbCEPD2gqp6c9erbpABT0MHYDDywrM7Tkkt7
m3S/hrrVG6eL8CmdbDxbHRZjvcsHg586BelTOajpvAPyXKq9+rhw+T99CtSMGlonIC4mLnWR6XQk
ltKlRh1B2KP0YcTip+VmXP3RzCEbf81xGDEzBL+/Pau/lw5nujGoj7VA1JhLhlk7W4UaRYDzO3nN
cO8xMBGhOhJOm8mVykIdzdipqXts6+8Rt5xnnJ2oN7f54xgUhX1OJjfringBKJc03UGnMGbEPoPw
puizbVIvDW4e/xGAjoaFRXBT3TGeAOYRZtulKZfX5rOYP91/MWCBGU2b8hSq5emsPWiNd190xzP7
Za9wR+AIxFnZDAUbu/hvzS5CkdftAt5heBXqcvkxqGTSreU+P4c81B2jW77A/9Ekf4ILgnU6oKCC
nv2n8hn544nikW1p9C+cJQtloAd3jLFNSBYy7X3txljaACUwFmfTydztNujbIXeCHTgJCpfHOLSp
olMy/kjWL0xQ4BtJPBoWGqWT9f7VTcHOTnElzvFVdTv+sj20QfxTk5NI5GPDrNZmKiKaTYWD5bjA
agSDJ3ERJ5t/Z7Ln+957IPvvn290+LRcla20q4EfH6503vTRxtfjpZDJDkLrimvOYt3LQpa+WPYp
4np2MCdF3W7+jgyzQ4UTGgfbZKeCX2stEWdWhFO8xBywAcN//F8kYgkDq5wC4cG057k8ErQ41Qhr
oI0/Y8MgZizZrTOdhpQOdcuiXBF0DSPuRldN7B84lpq6YtsmxAob5jxYGQ5BT6fP/JbvHZ+YF/pD
GGtNJ2URYt6iN8oKx5GoxwL+3s97vUHaR0ziUCmLOEYBEk8DUe2cckTIeWoLhgHtwRrZkdQtF9yp
nYdLcbrja44HfX+QRZq2BIO1bPE6JVqahLUrYBVrGZoTi8ODGMlQopRiHEKB6tuy2HjuqqoGRGT4
7riIf+ufDVir3FbxoV59wuIt/IhVz0D+cxKpJ6fkpklwjIyn5rhUcE9w3V8wULkIK+7JPQc+IJms
HA/bUYDppJBZVt4SMpoF+vGTrTDFXOeB3/j3XMHgGVwYIHd+GbnMElEw+opzmp2AJm6NjG53c+3U
NJUzUkNTXdnPinVUUsArqY4L5SfyJrUpsbW9j6YsFLdVh96JrZCry2a46qpVP+Di0qOiB8SVsC81
J2lGwtb7UI5uYA4qOq0ZHFzTOEXt6Q5OX2rAHkxR/NppSp63yI0ot/+CbxqGZL2disl00H/IIu+U
pvhuKTC2cKsqqahbh5ZaAF9aEvf5FYxPS/oWQ13pYqjL21ffiMWI6hwlBW6F4hfFoHyKbAZDOYyn
8F2YOxSU4en0lTtAco/1cxV0V1hWP4E239ymuyk1uusX6Rg/TA/06KNKaLdgM7Mo7JbifVT3T/VW
oGfSO2YYkKPlu25/oOP9N76kxlc32WF/q/hOQboJpHxj2kd+AwPP5zizW6KsWxnhqKngfY4RuqRt
Ls2OnI+OpfXBXhS25jO7J303gGx90ZZLIz7m/9TfGoFeWTmpV42TL+0xvT2NJjUzWVdHO0zdpfyt
lqoCJPbnEK82lhmVgWrI0PTbPOt2x31rphGWiFdv/7hHOiT8tYdv4NqWiZk1HbJcz1aUbxdT7vu2
L6jbCDPBQEWxd7rnWiDzF6d5TIEdEeVAoUY4JE/GC0aloH8g6V7HvL0bf0rwGFRSmrKJIkvl3vzW
XOCOYnday3CGtDs54ysqfOCjmqw6v7CxUu1MT6lB/nPpl0kcC/AhBlPUQOA5L1TpbqIIo5GBK4hw
1k/x3YiWHbFBJPI3UClwf3wOFrgOEWI3wUGRpgn3XfQQ6Nus6IS3k5TE/CcWSfinLCXVbfEQ7sCj
PThAbj+Jj1W8n3zxQWfom69V/oLfAhpaonj50/Pu+ZFoFiPNSMk5ZGoXNEkVqzSD2jaNKkxw20zU
7hyT5zzQ1kNsJx23vcvCx0Iv29iZ0cckf+NbUwSZ8zoVn2od4EfXciignpw+INwmvRkJyOIPKjtH
SjGFyoVBI9jExqW7mptFt22uZeB+bckLvuRRko/nmEqlHiEUmuDee8NxI4PWNYBc0IS1zeCapf39
ldzdY1npcN895wOqj0RhDYJVIMzip9c3offGe58lGlsqTsFL5uV3EYdKuAH2ecxV++71kzBSqbWB
l5qydSvZ135Qm4lZJTtiTPyMQFA1nX/YL05nG8MCFMy66dilp8lLe3MmGqPOjHtNt4WDqC2fwPFt
uBdoQMEgqpWQUSWE7z2Hh9QyA4yEwN8VB+tT8fk4q9bo+D0eKFmdLciyjnWBiJ5ySbHyz6tjtTVk
1+7ntxRnC+BhNmxpygdMmD0dtJebe7ojxc4rJXg43Ijxsh1jVCOB7qjRJfH4lIFDDwaPMxslb8md
uz1ovog2Eijdk5rFPM8BBuni57QBF22tcZJAWrXokpYukVuKrxTQ7QV8DqQll0IbSL0I/Vo/51+v
E9THICl7fp2anTMSEJSjAUxRfSAlXdMMkKWLkrzk/eaiNZ71xxAtaI9zZx9MJu1ZUs8PTWEbWDsK
s7A/s0OXEXfqZyeCVAMm7lCM/x41OHwSRosuKm7zOod6wUNfq51bVuH+EhiAIxhmZNu5Wr08ochF
e48P5TStTAuzUS58szWN3rc+wDdPnlDLIPtMVSemRrSsyv9NT6fv+f3Sd2FsahWdjLOSy7v/HTsl
Lj+W1GWrdS4QtHIrWCaZN1mqxy6BQ8X4GZD80YWq2FtIN7imcO1Fjh1asom1nJcXSa81/RfEW16s
nc3CP1Ub47BDj5pxRcw9VvhbHTlF1Ez9rzQgf+AZD360bub7tJ3+fIVD+V3o7eT8O/rymEkFKjIf
quAy00AIXRW4xc6jnB/KokCV3IdWgij50rFEAx7gqlpq6W0O9zDsBZaFQXMebk7PFRrP2z3rQA5c
I6l+oxAXlt/i5bdyai7RouMVrxNyiOcwKWbQNC+6Y/FZxyATv1H7uG84GVEPUYPy56uSdb5R5KWc
0cII9MyXcEpOySRAG6sOXE0uxLTAsG7uUtQEMCn70kmcP/ctwHr3gKjwxvkTQBc0+QmjnnNrCd5i
9KnpvWFDFMfEp+SBH4T3AhejE/SpXQuPAqstDgCeGuhplS9t830QXUehfl/UknR6gCLmX7RjOF6P
01dDp3wfDC2Wb9PYveN7QfgxEWMEuiBcD+L2xMjJNNFsHwPVXwHrlycgSq8Hzcgh8x6hjM/x6+WB
pX4NJ8VMSmhe/ff7wp/lx3kGp7pwJfMQ3DN0CFP8gi8KQvS7qeTHrpqwlhT2lUUHaJG2iUE/KtPY
RX5d9HhWT0ZXSTe8HR4TDzthqpXhjCQ6Q7594IAEt/je2csu1upvd0eJ4CgUCicrbu1GSk6LJ+qz
pD2VFPUQrO9AEn5ASdQyTjpJNZji/ClTr/WqnKA4vSjtiaVyN89FX6qh+2TbEz3/PDNlHzFdsb+K
nDiDGd/CjLzzIMKxgF3Dr4WXwtKsdW9vC6jG5GIRw9lvJDaPjShvOZA5IhIPiO5VYsjkgZRZdpwB
IlfZqSg+TMaqHavmUDx5PJoxOIJ7cCUKGli4x5bD/avcLhciHG0+7mi3T8IMaU/DkM/EOd+HU58L
Zz67nPRlca63U7YIHiZQ8b536lyMzvf2/XJwoysWLOH4RFw0EkFKZzsa3GhHZgo23M7zznWNGHav
/An+60/K4RfxmXdKhot8+qC2oswHlOZdXCckEfyYxD9RH75T+Qe7kif4vTEGkHnRZ5F+6s0H8uXX
TnTiFa5YOGpVWo1BwBToC+rIk3RXy3Sjm4X0BglmopF0HoZ3dN9uEs+ho5pf46f+fMPVwW0mtY5U
B4sahduWCm9Ojac1upnv5aqz20cK5zU9iVwHIlp8kNZJbAds+vCi6SLlFNiD/3wZgJblSJpqJA8g
4CUo7W5ldP1zIqnG+hlhf/30Ev2o1QTvNz+8daD8kDRW14TliIcBocjb+y9XD32fkqIAii4pKSbE
DOsZ3lJVB3tomMrSpVtEKSw4CVqcPaKrt9xnNGE16aEM2jGKsW0MMmBrET24M/FIx3DSOG9MqNi6
yWevs6giM9yePQVMbTMEaTu3HXFjahCwTYPeeTgIe8bvpGAQGGuLfK8RlPsGFzk1/15u59O+Ri/Z
fje+LIU091wOUB5DF8aXIywp6chdZKPCNKfulGai3cpcJAgS9K3ocXaYWhe9s0hipe2sKOwkgCUE
A5KoGlV0VXzinpfX2SizQBqCyioJCDcKVpe5AgfJGN9r9taOHa3lrPxBSgaRlmV/c59wp94DbsqU
DiKVcWsVmyLLUya6hsYyygngFemqQADGmRnhbKchJ2WDTb40xi/jj5w21letB3BKm51k1rMk7yz1
x/AplCKLFnxPJtOQjdXRRB5E7cMfefQLUT2KiOvj/Ln1JG5cAm2SuXoFaMIonEUnhS2p8h+7h9Bv
usUmq0Ij4SokBxNo83nnU5GQQWiGdO6nIVKwJ+wG9EsP+LbgnwQ+iAne10UiYBPMgeLgBp4RGsWt
YTpuCYNxyFeeqkRd60lwHYhl2sDje1txFnVQ+CyWAx0BHkcIXw0cB2Prd/P/GMGBsVvQG3b9brX5
/D+YvJjq4ph43ptEh12MLgm8gbXr37sAv/sIpxT7UiEi4uOrH1+SctTA+2E2h4BApbeqJ0DiNIL3
HLx40tWHs2NpXLoBh3KFJLfgN5QY/nGa12HGabqZ7Otkk5ObX7ILssWViOqqrghIyGP+qLmLJL67
bMfhs0ItGJjkhjo4tECrvQYkLvZCYLVJ1rcc12yKWyxPGzE5Piy7MNHwA2HaubEccrJwgmPtbh+Q
ZVims5dyI95kMo/GJ6rsfH4Ah/EFnse5oB8rcPJP6ylrOpLwjD9CCcWZjI5qJRTnjVLXB+56Pj7l
vlOQJMl0c6hsouIGloMqM+S2d07a5iDmfnYi6SSRVCTbiRQ+iIIE4BmD46JxA2Q8SAe8nYFUK2SW
vFpqh//PyeXcTjwYppaZijMAUtpjX2clli+MVwXbVkid+nUh6DPQ2d4fHbxXUbxkEJdSyjyFE+nq
GdfgqJOF9M4ibcKev+3qks8hrx1bjNsR1jXRc7MjTBBC9LR+IK8rvsGiOlJU+eMO0FPK1sA09Sw/
BZ7xUfoUJq+l0McasxyMmYIpmzBk15R3z1Q8K0LVQZKlZaoJEbeQnkNgrds/Ny+MwrXhxU/vTIv/
LFLr16bSe7JM8d5QSgjDPj6ZlAqUKZ1AlFB41/2AI2J8c3H3vDbZ7kIxEif3aOFosMTGB+Qkaehy
lvUedFPQQLXuWQhTUqFqPQXrjh9kV33h0KtFlQLSOvDzCANS+yPzL3msjrSoLoRVovZU+tL1o2k4
pprFZPu9PVWgJtzIFkrCEdBBYpUnsoczPgHLS3eVe9kLH02asAvvggaV/I88TNeEePo/SoxHtGLy
i+mvPMQ1rxegEs60ocsbTu3rLJcHNymrbTGAUXiRM2GtFn5Y4i4MYUST5yCOhC4/pGejDivhi4IT
wdhpGDlLge/bihsybg20hDENK8CbLIEJYBlrHhUyhlQME2kk1h9F9Ya0UXMk3uFSoiCO+Yfz2Pvo
m7s9muCPMRmQx3qH5XwtAcSAzuU8flc+OsHUAz4/biXOhV9m9AYQ3vNcxJl3hWq+rJz9KX5Ckgap
WbgXjKerZ/E834zQ8LW0J7jMuvNZbpJREmwJ2/kMCbLGJHXvkBuI82vW3mdUvrF8IxDcNRwNZVZK
05KbxR711RoBkr+PdWtIbp464axoLx6mo92Psy63hH2+2hgihGpQS7TBsZ9t7WHS8EtxRqaC9TOg
5z0F9y8uXn4wfJvJ2iMyvvtkDXasWv/GE7WhWexcrPpVGVxTP3LeCjRYwknuRTYeonuZO0Y1Ptu7
LeGoBH/7wTbpvJRN56EIYTonzakL1lsm9wVSYxatacWQjG361lnufCzNVkrXHXVfSJ9i8Zo2Tv3a
qbCESt/6hcE0eeoOIEr12Otl6QswSPwmATU5eftM3jbDbZy0YQf4969cz47vYGtg8OIX2cUTjygj
g2Ekk27o4npCCYZ4KM51YBK3hsInBh3fyqluDOe/j7x0rL2trdM4IyH1dmEW+LObfDTb7GUy8lBU
/jC2rkbBZTG2+6BBKXPEl/D9SXt2tN9TctKvXBGCN1t59zsyL0URnEd1z5kSYqTAwzRx2NyrQGU2
LBZyHZ4+UN/SGhFWQNpmQKbKsktsoK7ckKO/X5myyp0RP6wUWOJHXiYzFMpyjLRhA89fbPhAjJjL
9Q0+AAK8uyCXd29UbVbUJ6wDqTYvZFA5CfNOOSVz2SIzEyy13bWiJxR+pgaFzImXVsFIEeRliXVi
MEjWV+On9S3XtueRT8WYMAmXr4lLmmMgHz/YwgnJx8uZVeB23sn6gvhl0etNFOvoRfDP9QOApzse
LC/B0NqTckJhiN+mjEgFQw0BR85soJxriGvN8rXBpKwg6L/cA7l0qhhCmu8tagyYwLTfoK5qt9Re
VcTxXWTtLnh49ACCPcFKBnx+bgDjL/gkXO4sYJbnZ4SN4O5mvP+90EllVnlV4buaokuOBj2k3G2V
Bq4D1cjuQTJaLfJnW3frZMZSzNT9fYyTcTv9pa83YHsbik0fDKTTaxnEYy8I12sIm1vp/1NB3CZh
BiAJZZ/ceLo6zhX4bSNth9IYX2U6HrnDrShRgFa+P66ACjAD88pHz8z5eKXtbGY9ilJseZWPfGQF
aRUOduZ8YyLYQ9SbikzevSMl//VWxl8Fm+sZzzLXeJnQVKkBXY5dvQzWt9txcgLCkKVeUbUkGp9f
CfOUrFusN/dckfHlxpmya/hLwBXW/bChPXbxbXHgWfkdEyUVN4B1YQtVfjBWSkP8rjk5mLJ27hxV
EmrnxUFCHHzMN1iERk42KO6aXJPWFYH3XTmqpZNd1jMJ7S4n6tx6naNI8SF/LUldn/sJXX6wIkzq
A4LepACrrM423VxSZSaREjZ20g1vC79rMDKz3nW0CCzaZXCigWNt/QFJhdgX/Q7Bu1ocagBd2RyN
z7RWZJtGMBtmFkR2w0P0gj3or7aMDmlVf0r6t7yUsSYfA5yvinHgHOdUtaDa/gHW7XmdxvrB3VNA
BiZuyDj41ApKtWAaWYtICarj1/wGfXb4iDjWr+6nij7S6eWzw3rrWm56R9B0eQwbGPfPze86sHYx
iUki/2frgr+Z6qwgdG9mko0382NPZMVBf+/s1xH/9SDynxXgLxC3LzrgJIVGwGBoe4BTpUyspOZO
p1lP/eBR7NXixrfaf6AYB+EvyM/P60f0hMcoSs10WaB0p8ZBZmN+0jtbFueoC5+FepA4+m1kPYQL
E81NR/R6yUQLonh5wdrKHxoE36P77uE18B3rSG9DDJCFtf40/hiPyDbOQyxW6znhDwhOkYSxtcfP
bl2S58enULT05arw2fuZBvRWXpN1j3HjeJ1Umv/SitONPwQsQEANvwaUhCTAPO4qJFJx3tDPupyX
afqcI5C3nOzRGFA0FWyyoDv46C7hDt50KLer+cBi3JJLrY0IiZdh7bLw6pG5Rb9u05qTzA7zbWgl
sSDolCXhHwTIe1XjxJ5yZ6JBr2S9naApG1qEdOw9T8hpvk3Fd6pWCRJHsBAWgDbTx8M1pXsuL5g8
EkyvPNGat0BLkj2QOYkUO444krg541B/MpCbasYpoW0NZIoPd1Ewo8b6ElHvhvzTnnGjCLnz5QaJ
O1EXzqK809AKET2St2HNKCitI2NFoTSPP1Rynf5IfbFGvUchE03zBzNf9TxDVp90o0heVaTk7sxJ
Mz9XjQd/N2wRh4JVfPhagkhmQ6g9VbDlaSXIP56MhQdiUXsn5zAyXAg0ojPuQhVt98Gl7M7ycgHe
DyGE2heDJ4lT6KqC+rhXxvAjnmGlW0udBa2wKiQ/bdhmNig7ESwk2EuKCuFgXm5vdTCij5hqPQws
CafSC0wFy0okZ1KV+e/GEHUmv7it0r91bTb8dfiSNwAjHnFc5GHIj6HoyLopYM/uZteRvNYmEpRI
8QGAptKk5nBZ8P+YXq2o7UQ9Pl/+lSxuLzLbANHqwotyZGAET0FQJrQ5ONCYL8k4pZFBYtlhvMFb
vBjqXux5+l0nEmLQq0y5CPOQFRql3dr29zdJhuER0nDDwyV0uRaFMczFPdM779BP2NqtTivlnFmd
YwsjJYPyTgo6nLQJYZRoth4fzgBerxnDYREIa6Z4+Udjs6TiFeQ95JlTJtvwsBGJpVuu6qo+Qo5j
o9m5qGcxGCsfEZ/G4ZGUj5PNXajFrVEXWxFZIrh7h3dI5bwyT1fskMoM+KtKVIKdtlY3sukhM9fq
WyH6FWWSM6wuyfvW7y6xmTlNFOl4B7uONTNjeRFcUmInH4qfizzTDT3EWZMkeJoFoENbFj/kFgaV
eZfwzlSxWovi0bOnX+OHP282HJNEBJzXPDtC8w0gYuw14XV8crL3RqNu5ulAyq2onOnuOr7ex8I9
8kokU1kpaGBGP+P47mQH1gcDdFtxNGt9Gd3WBnK6fbmp/xu8MEzIsDooI8DbD9GNFUACzE9UQJdQ
XCNoWTpQ5cXP2q68AA0W9BxTcoWKks562nF/mLLvj6IJHniiHIo9QKEuzR1Z1hgd0s3BdBT8OMSe
rSjWrNE/4wXpRlp8nnoWkCg49YNhA+N2b741R8XdkjuoT+P4WQlrWkR0o6o+Qrqu1MhkgXDZ7L1B
6OOematc9sU7usI8tY3YjE/Reu+1tKZgBFk/gqhi1mJK63crURCEZoVBTJ+9QxBvB6gtrzicfbmZ
QeXSX4TRzxDzLyJiEY7HOxFhpBXzUZkFDHQjI2/Dtt8Lvx+7NN6Nn2bXFawdo7TFqcfTozWh1oZO
YPuegm2yDpGEGu/sKlvcPcCEfI/eZAisWx+PG88qm9mrTwd5vggDLQR0IyXtR0AAMt6JXdpDjMjg
pGcDOnCYC7e9/tO/bGuJucBJLonGd7FJii0wJjxNfb9AM0ImDilczbqzISNhDnDJVZSebq4/VrEY
5b5ABsHWefb1EomOAU9Xablajrvf1Bohkqg0j68/YgVRh05sLXADyizXARUy7TP2kHS7pMTbP4dD
OgPDtoJfLV+zuQEV5mWF8FOgq6v8cEmuuc8/teiQVVc07EpQi6VZKazK9Vso3UmetLhW0Lh4k3+F
DBISSc3kaRyr80DmpV14OS391KuTLQsAZZlxJM9nDUXRFaC1HH8lmDlVfIA++tUy9tzCwyEsVgAp
pc42MqLtz+Gr7lPrxGtf1jsTZbZ50eB0LK2cPSFuP4Sz9Km/8wG7tnnhzT72QunCUix+NOij5ua0
LUdryh/KNmHN70Hj7irSIya/fTRf4jiTi8t2iH1EYS3aMYJw9gJqa6ud0VgYOXOeUNFAQ1GeMxq5
GZvPgApjF9RevU1/AZbZN+TGWpU+IK5LayVQLoMWKQBNvL60vey+x5EJXsTqByFgwX/j53bVW+IN
vrQhA9OpQmZpx+QcvC5Cro51p0WqeGFnew2kYEuEVcqdb41KBwq3WVfjjEqLkL8Szhr5o5aPoQyO
Bku9e9zKg0Gqgwbu9994wGDh1scNb9EL/4Fr8cfs1xeF2VWokwWcBORjHbAlCfI1DjsgTTaq32X9
CKuTuPGn96KJ0/6mJ/1BZ4fhDOnyiDoe2Jf2v4bT/OOOULwgtF08fcvLI8pIi6cbmensQl3mKLhi
4eC57/+lmYmsIWl0kOY5xzgRqEy94+W/CFfgNOYgaWUL6Zp2RpQYzQJsG/g1qzkYIG4Gs6KS7Bkp
Ue+ZrzzZ3zArub9C4TWbwqVohdVsCaZ5llxyNDjpxCCc/2Sa7mnpYa843dDPmm71XS4j28HWcOIr
YeOXm5IOcW5AZV2OvZoYhlpk0ZbelIyr6c3YfS3ZKAbe75xfsM0Ypzv/9wERGK2atQf6IEuEsjjZ
hOl4ZXPIXyz9hOx152DogdiPP7HdJQiBCcsZ60JCKWt0z11wIV1hPcf6FQ0mT/eyyfxaPWzGbgb2
Gds1o+A94QGnUfosW9lB1X/UgG7Whs9LXyi9ge71mduMUIFLvVL31Xvskcu1cVox3RVW6YOap/6a
HonWZQlIh16chZY1gNDpJErfATq1gQE18fFtBiEUNXJF0xo7/MIbXrjyTB40mrdMnxsizq6h9k2X
E8sA8NCoPcJZw6O9XltlA/Xfq8V59lgyEmdQUFVCjdmZ0+wIuTnGNh2KkeWK3sPmoLfck8F5PtVO
gU+d9X+ghKLOqKFTFkYDH5XB4OKZz4+m/cqkpO4WpYS6E+2VBTf+m24Vk3EjI7BAU/AdwGa8oFZe
K22iWKxytocB/h9MRpY1Rfwk+mOIvnWSTcDMClQMmAgn7WE6i4Fs/5L5KiwU901ZdfS0OnDouaws
cEbPMtN/hbNwotoF277FXQH+6zFIgOSjSSDGCHtq7s4R5bFl4FCjwL+06jSHLYz3lU12PwfBUMD8
vEHH+Hfm3mgY19kciCHcBqGyRiGoHdsyKuyf2tt9plYnxZIRrOybEk+ygfltJI1wJKD2H0J5OIeh
iCZSbMQUHraPsiVF+lk7K6K+vAInBwo7ufqEmQypaF5VyN+dtX/v8PKTQDc1ZogtWozPMj0VTUlk
4i+Ju/jKdIAgsUO4Igv9l1QdfK73udNQgZtz+gdTwLtTpDT84/iVdRs7gnJ7ceNp5cX4sr2iMfUw
D/Xg7WRFAfvFg34OQvTikIcW2tv6eXWcQYnMfTLwpuXJGZBQX1GVoSb2K2eicwxSOn5E9BDtwDY4
VxBAaIJ8Yye4NA5Nvnqq9G1YfKFxRmlITvnO8oHJb5vkZYf3MeMv+srR0Gmln02iw+qrecoJO8ND
0Iyu8KBpy8UD8nwXndYHWBu6uzmgUxFx/lgm2XvBn8HXbjmFhvoxVnSQ6cRgchfBq+XgmlS6lwbl
5UbM3LKCn0gKYps7jjnRGQ7uw5h7mpxYf8BJCe9fx9ycJyRnAwCxMi23WY0F3okb3Q/PNQGm7LCk
LEKHXvbOn09uoYwxuWXV6z/7OCyRgg7SAbpaUWNR6bjAj4sskTyAkR9rAP/aX6OjN+4FnMSOiKHr
y9lx6bYP9E01VFwHcRHgLjsP6k+gcI9Pngs40heBHzPr5McN14MwJkAiiJPoDEX/6RV81+RsDfgF
+14PeS2Kb5da6uvlqXg53pgIRRQylXR2C+QHb01FklkhOkPaKQr6K4VMr8SkOgRleGx0cwJ+E51m
cggQucenJlwbBanNMPGfWmUcjhBROd5ARIvqRrjEhjoO83aus/N1QbO7eH+lYC+rrlnr0Zcg4J9u
56geodLQhhcV/P8KOuH7yrYjewCmNPDiaSXqk6ulcBYhPnU5pLAOwrWtR/HX6WuhG7gF62HzSUcY
zBgB6AaphdWg88dwcjLcRNgzfUvxEt0kxPOFaa+IKqfRucFlRuptV2Shy5DkDo84BUjOsHGfhyY4
33zm9Igvr1UyF8NtlO2OY2mI3D/lwxPABIQ/DmkecpGj1sAfFLaXXKHWJr9gucXw6ItIHZTnIRFT
f1/3Wu6gndYmnMw3pgvyzxo/V/tiPzPGsqVDOr7TtdfqYeSbpX8hXMOkjRBMLnCB9bG9qPTf5A7T
xgX+RPwuNNyOW81HgmhXRcrYRKoVKtdvouJUR/AVH2nPoBoFKZqJj9qq3njE/rkUW7gVLkh0DjNP
IYZcCu4eczvTfYlBJpljNzT0tTfebe5VXWIIyE/koDm1lK57kFp0jjM7xyCzd7ghoxmNVynYEmq/
erVWYd8c5bu6BtsU5aTq5Zc1xEEclv4HhN3PRjI+lGFXpCoLGfk+J5TGxvK0JHYo6NmUtmtVwjWz
T1hxehR6VlYTRD9gHqh4SjBIDB9HQF2QOeWfVqlcOCggJ4LGWXDpCmelCT5/YmVhaR2YI9n0oabt
EsosNF2mA0MYqXhn+lxLO4mqrZyv+jAU1QG5hm4hmihrRMA1FBHrt8wN88v3JXtE3bnqv3EingIC
5JKyG0ycjx9nuUP+aTot5vYd/QwqHRU9f1o+k5LhYXqcT6Nyf1gqq/ESRL1GBSkXGugzp+IUgArx
MB6r94GjvJPXfr0gE8H6dhXgJNFdz26ucw12ElZ8v+p584scRo1IvE4cx7toZJi1TzfopBKedFxT
GQv1OfjxGs+pGggrNwVJVsukDI9MAZQgzXnr+v4OmDO9MhQl30xNpgzQTAlaNFq1E9+TpkKmr4E/
GflAYyqzlLWhGicDcAP1WfIdtOI2m3PraUuGoHT8Frrpt7YTfkdv7rp0pFbeh1KuTlcWDUYaiwWr
ZVEpj296nwtRRadt1HEpeSYgx9zCRjr4m8osF4vuzVY9SbCDIW9+kapBJRai9Q8BfckbdwNNGryR
l1h+RgjsQ5vd7pQlpPiua8Bb9rfHtDydWCmZiJdzWD3w+ZXb+iIW6LsNkE54eKJbgJ0HMmh7xQ5R
+9TNS7lVFUJ2p5wyawXYzePK3Ssoy3dgZyZFRCW1JFfKVCvWpQsq4hnfQBOWayaQVIL4MF852D6o
cUGA8GLzBuOlXT5lokRvexmGxodlah/gp1LhPAh0g0UzL0V84th0uR5KGHuG57P7hHv1mG7AUnhX
UTHGfzTeYbcZByrFVumAibPcj9aVrTmWaXozZpm535KT9tAFaLh5J3YeARJi3Up2tVmj5XYYc4iO
mpk3zxa7e0d2DYdfkHIxeHThk14brwx9gWOdJbVdKtmNzFJVyfkcoEooNtHyD+Do6MmzACT+Hl2C
7aTTAIbI9Fefny3R8Ra7758HHQ07lWF/3apzi0Q1p+fbyCnQZuPLQpwmOAdq7URTXpxzqISxL3i7
sifFhKSNBkT+IteIJ7W5VOh29BgHL2v6duGdbpwc6kRj31FOkCGam0tA4GVCtnEOQdby/84lCKhn
Kc2jLpIXzxzcyfELS1WSZbbnf79jSh3+xvryYiaq2eFpHzpY7eckAWjcyuATwGAaUfocxgOZYT6X
cY8iDeVUm38GD6xwd9kzu0Q1zOvdPWnk0zXYTkD4asXRkVZT+4E+zLW5Yd/NcoU9zzvIDJt0Qm9n
fBDDr0fdA7iQSfz4cQZNY7n7EDX2B0DHalP4IVFrFJoeGEZFUMkBfWkO8kkcF8fy1wgMTOHHH6U+
GhSxk5EnB20HlJfrEaBCITgOIdZcjGtAkNZ05lFysVMOj1b3b3oF6z6aPL1bq6JZKW5YAWKctpkA
LW+nG304Z0J6Lb5AMwtdSa7cUI33Xs7ghM6werylNL4jVc4K/rTYNGRkto/CJJ/+O/ZFNwZcbz32
p9gqiKP+JZBkcmsGoPs/rI37FyXWY65N+puC0XbVglW00lz3D5OdWKe0ODSy7uSTd0XJhzL6QbuO
w3X+a3ZO2vsYZt74EvdVwb+lsWAWIMaho3BUfyfom7rQGQ+nekgbJPzqZAs2Eho2LmY0pBIpNu5N
1DF7n0IbDYDyk3NmN1YMjCO0slaj9o0sLfCJibJaI7CifgJ9eB9onbl6H5XpCwe2XRGMydgKFc02
lD1DBgNDOZ+daBODbjhvxTIJJbXLwiXwYvYjYoLSEeKGyTJbZR62SG7MDpvtoxZpdm0V0c7Py94q
BFv2gupsSK6ywzp7JVxlQfehDL7oTCIrvBWoElJKmLO4ql5h2/WdF64WY6iacBFgcm+Vv65FOesa
0FTlOVRNUFPFxyy6LVzNTNfolPwCvcRDNGy23y1+8qia5/16JMAp6sUKkwt+0Z1BYyRq5g3V5P/n
J9FTusmBPAuIZrBxPt+sMZcQInb7X/wIkAIHrDIHvmh00u5ddIQhXo94jNzeOimODU57SYtK9OJi
EhvrfPF9EtYt95XcsuxP8bq/axbwjXtGD506hNU3U2e2dJ33GrlSTYfW4s2lYxOrp+NmjuL4VO8r
Q+FcguzID7IiiBUxpKS23MCWqndoFH/6htqnTAaK76Anvonv7seol/rCYkiH13YYokOxGFPKEJj6
E1F79PDXd9m/nJ/ot6kOJ4JeHTgmWwWSJAANlN9vClNoxNbTcU0ZUy/ua7VfMxBniGdndutIJTcr
e/VomJcEB2S3NHi94RwxbYtxy+0xrQYbBtrfg2gazd+2hH3tl0TmYNTlP2OcU8wZHfx64DeWPwGP
BfFAj9rJYT+rWbTgwRSbXAdEswQ441exqxvmoMaoo/pSeSYxiRXCmspbKsuHH7bKqIR1R7lvlP1I
52wDyg9JtkHRnpf1RvJ9jJL2zVuhm0tIPh8Wqd1IT4m/oTBfRK87wkYg+zsLR2DHE68eHRuq7RDo
vcpzDXuYhBwQ99LbFxAoZIJqy7zgfr2BxgnyLKhhzF7tu03nmHEHf65pd2ne7KJXZXoIrx9w9/Oq
618iww6/1HksxOP1Y/R0ChcpUm0qG7bJj+TrmXY/LuSLIb+y+brERF8fDf2R14HFTnv8qtFuaDxR
Z79SaXTmfTuDdxa7EqehNTDlzI1qI8w0GY8I/kYOECeToOmIMxYVbDpU9z5qCWXEXYTEq9TdGC2u
AmOk8pnidKdZf9xZgqZQDxG65aAZavqYwa3joSGby7EvlF0TrOVXaxQ8sjEoFOY9l644knX/NP/E
2mtZVq1lSFKn4H0RmgNbw3XDLsyCH+CQS9z06bU6IFJ3xrk7+rJWCDIhpr+rqeJQYMyEwujcvnsi
jnA+xyFvbZhdE1aCs5p7zjnysL1FLDy5jVnYZIfNAZ9D1rZDeQ9gOhiCq4++OiZXvg9a900AGx2g
qFKenRjIURiDtyXE/1vpYItZoXIiRj2h8u477uMgkH5LbxaNFjs7ZzCwn2b+ZvAniVwNqRoB798A
aHiaAbTcxx7ewO4HPWVnU1VTfzv07gvT0soJjtrBm/ickCyiXtJ28P6JXVr69/eSbP144kRyCPEU
IiR3k/HLPM3666/hJphFrkLthLYsp/iWWBwz32YAske62gne22tuQTX/EQ0qUUMWqBrYD2MRHQKP
DQMpW5XVNmFvOHZnz/1kSu2cEem8itCnkttFT+Uoyn+gs8m1QYNnkEXQ1X93xv+WtMopNPyo9TwN
udaUE+iI9w7m6uVF2hxYKeR6lvUQigbRWaFH1XGmn7toH3rCagB0ORX9oWl3iABDG+BDEW20NOdP
iQjxQC3/r3Dh7jIeREltAkOulh3zYMDQIY40tBmMcs9Z/vjZB0trZcvwin4tuKYn44jJ+G9D5P4G
hHBR1HFbiUVfQ1cHTaHpJ5vur6crhuBbQm3ea7Rgiua6nbp2fZ83uNhiHqLV4n9wneXwMqZQ8xvS
k4EwlLXesA2kqTgQsCvbzIZqigtd0VcU2+agQ+P8/7zM2lE2YhJffHU4OBIeAhnhKpjWl0A2sRE1
YnCb5fW1C87nz6cxAkINBKRo8b8seEZ/A2c8ShJKY1mElDWvPy0S9/tz7ln8XiMTRRFTHwgAIuKx
0lDVPsYVMpNcgbYEIRxfZmfQNamngC1IMe3gHSNBJ5qkOdPOUcjBV7q2zkdsTZArM8YOZnB24hbZ
Wt/ohTFPYBGY6a05/xplvpqodF4ttTFwI9k5gynXBXlCQXmYPJq6UIy4LVnWqNq911Pyh/SAM67v
0Kaa6vASpHLozPSkNRUV8vbYiqZKu7DzlDLXhRrJgRz6Tl36+NY9HYSTODsr8cHIfHakrlcEzeDS
7vybbWoGwYx9UYCUcBbKy7ElS0oYpGast/fVkToy3b+2/wX6k7+QLmAIEdIeGffsm6goUBQ5A8gC
ju56NUONdYJBKLtSDRTe7Nj8/kUlOCWDle3T1eLtAdhYQvaqevX5+8g89VRvBYMfxptnazqrvLfp
5fN+i0otVuS82r7dwsUGmbBwiKq32uBvHQOVFajCSHFjV7owEoXqOexl95+xLv6enYUMsyxhsNsG
Y2nzfHtl4aNDf6nsFWAIdmoOxyDv7EURMWgE8bpQmy8j4DWtJOThoWITj5sVMzix3rd/lZA+BEnB
uG+4AJbi5T4KOymnOLrcrp+tTL412h9V7VuLygbcBNFBlg8KOaKe0W2gUknqQztPBPLkZsa+4bgF
P2fCkG6eIZBgqWxl22veghpAJNGZDScsZ+0vgNwzvL1ih4Rpr219FCw3iWcfG9Mf8WJob9wcBF6c
7IqlxchZ5nFFul/QWZigpi0BMPJ36a0Qn3kSkI7eaGg0Epjn5nxCmq08wzbXRAwYY/fDd5xDKOEO
nPgrlAXhAUyFUKJmT6GJW1zYVWaMPoVS6niTf3EndumlhSZK+fdn599zGu7e4fcOUzur5RNjSY6t
I6UQzWU/BPhLJwJKRbcEKfPpngDscYjkRusEfPiIuAbvX1n87QbfWlAFczd+C8mD+tKeaE1Rx4V6
Qv3wzEnTVShT2n5AkGrJsvuD4TozSoh+mvdDKFY36a4QW/qRt/de8gb0Zl1mcb97Ncu/O+S5jHMT
jYHXMNBj4XXZNnydVEChl4Hjig+Q56PjhW5sDh1ieBQoYM8EKj9n79cyASSFuxd85yfC5a5MEpmH
02V54Zhl5qywFSNrsr9B0HSx6fqpEC4CiZgiX7yfNirCWhJFeYfoR7L+9XjWbu3O1PD8mkyLN71t
4GMxPvYxT86MOPQIucJZrBO5ukstL1zr0mI2DlKZL7vFVktI2zxj50YJqulimWJDE6V5HPTX082g
e4be6ocAF6dXC17Ed3SPcVySeXS/+kt+aqa3gPdAk9fZO0b0tu7sXso0R4Zdv9p1LqtL+ECSQzeS
Rb8t9cGu3S8MdlN/DduJROrQ/SdGMm2JhwM6OtC9pcFZriLBslPHkjK2YM+a2Ug9glMWFvaAVMFf
+yfjXuGuMWkwTq/riJYo16D0fJfCu1Nao5rJkCcZDHXS/jTPudq15JmPd2kKOJm48eJidG6qvktJ
tmmkJgK5w3CDKBks0D9xMzHAImYS0rkAW114QYiR37CRmuIyaojKNhvCp07fnCu9xdG1Yom+MbbR
yLDCzXg6eNb6fFynhp4ZanxpJdA8ePSAZBjMggZ+G9Uz79AvQwOUvPJXX6SGELcAHVDBqHGrKUpM
Sx6DdtdY+OoLM7R0/lbZR2ZsKK0wfNoyDqrb2ZjbS27lN2sB5g83BvzXdlXVu4xzo1P/AU76hduN
KWZbqyK7nSQWYqlS0EuFtkXxeJzXMeXPEqwBEfRTvhZcvgGJyV2jhcsOdwP+f+1woMpvKcM0hJ6A
h0Yhy8Mja50l2Dsm6kgA24asjtC3bfqH4vmwtX8TvcINmbMH6FsvzTVNCuoMB3xHB7rqs+Rbc7Ua
w/w8ON7ffxYQhmAEIptCWb1ZrdPixbtYIV/v0+phyT2jDPxxpql7xkwWFNKoR5PbAK07R+cwNpam
KsfbJAMU2nF4+ERNUWCTBA5NfMRKTNVFGhrUPyAGoC0tYF5WQJNYronI5QPPgIr78PoYD7imKjye
eJflvnv3MxKLNWTB3fMC4UpEQpZmyohKQydmEJmhscBVzD0MsljHvNlYmp/U438qXnWu/IcIVodK
2JvlwJpkBU1vFa6ODAR/5NFGX8zMJxrHEeRRNF3gG+tZ2FGbCv6pvYAOBy28nkgOHQ6/aRedHrqI
P6RLCNXTp9rGhG1GLYKu81Qqn3Y2tVMu6SuPS2My+HfYsmOmhwA6W3rZoQuFLzQdIylux30ysuo/
v9nuKbRCIEu147Easw65vzvvZYDEfHZVtyYj/+WzTXCFGUwzStkIlhhaudcNJKTshL64biAwodAy
5nALsKeBwYhp3zlFCglEgQn2wJWEK04nTjkHkOmnt1mot+Yjz0781FCJpHhcRq8AI7LVIpwu4q2C
TiE4RD7mdJzn/xXtnEBmitHHaFUrYT0y57eyzTwVLF9taaDkKEqstTusTFMmsg2lMWRomojsBNqA
//6HK1ytS18zI+ExHc6qHmXRdES4zZzAxGFW+J5jHSIF/SgGh8ZDyG0+KASdSCQlWRQriBZJLDxB
3ODR1ZAw4gzff3mTV/CzAIIaYcTVxgvNNYfcoBDqbPQe61yOOU45Ws62wzQq5nBaSniCiC20BuJq
SDM0WfiziWCEDg/99/KuaPLPHuEOXFeEbUc6mE9LQuZUtm7EhowK+gjzbYceO6RSVLfx8vXEPiFE
K8PIEpkfqUH/5wgFw9OpVd0pPmTXHp89m9dwtRHzUgYAK7sOerFiGzylPL5ixgYoJjuqhbnsoy0n
5bZLT/5Wrpy2aVS5yalTxlhOXRob/Lf51WfsSiPQH9IwAh4YZaNk1e/gXGnueoAjF7++eTgGJ0Rs
SR4HWdd7OkRgFhVu1kCnms/9k5yM+R+cF0dJE1RvbQ0O8V6EiJel3mJycCJlam4i1khNZBh1fotP
3S3Qo70k9BIg4OEO9q6H99Inzr7ApA27sN0JuEmvq/xfkF5R0SSlzuyBd2lVOSI/XJj74zOwNDsx
JaZTNd9+Scf/Xg/X+/04DSZ0QwZZwEdl44l4pJE+V9d0kPJHF+ZOx4sKYfWa39hQ3Y/qnYHpQYiC
3NGzP2HeyQuUWVl1V5HRl570CUeuTQ78K2fMkfnBE8N1hrlLKmMRBAWb1b/mbpC26IRoapHIegf9
mdRmwtHl1S3u3BKLk7o//EdXjKgyyuL5np+PCx5WoyEQkgRXvGIsDrsk5dMQnbYW6xhUQyqI4QKI
PgH0wegcK3iYQKEStQjHvCqjn4zdhpqEOpbEJSh63aOQJHzRlYuK6lOudOnAEFNOZ16rZi+hsUyV
RgSKXs7Nlvi4KUFBJkxwecx3kTyKfC2ZTd2B9IkpKTVob50nZctwSgYSGCGrcFS71/xFuWEXQqxJ
gmvR6aHYuMkwaDFvEl++wKBHYI35GFBt6IW98q/GUzgkj+nT7cECKdT4GraOMlS4m+oZadlPx8Ex
Fz58qg5u0hE1TLXoeOP3SiQGdZOje77oW178frTHJEUU462yRAxQa7Oza9509MNk7hl3N7X5hPv4
RxsF34EKNcfcxh6QUE31nhibYVUXknu5J9IIm6Qqa6zWTeZSh/xXxC19r68RloI4r555TBpuFkJt
Z5+FOW0M/9W6sYyirPj2lFqVh3nDRyznm334wUrAh5n1iDiF4PVptzBJHkcYkDmvsOlDhN48eJQi
1JBgcu6WG4RwTxQEmizzKPuvARxcWOCV3zUL+hqKVR9F1aVf+W11HrBziK3LyrTF3toBvP2i4oVH
KGjOvhEJrluanVTR2tDbzIDyJrXHz1s8+yNCp9qVszvkW8yFom2XEm6kSM+MrGORvZ8BxqiYxaSk
7c18UyoR8Efi7Uj2QzZKGToK+hTdCo1lK+cwDrOMBrQm1Y/I0BbSoE0wtg512LKF+/W65w4Xtoj+
c3uA1nnP/6hOqTLw8iMHkxbX6t7+7Sot6DY1G8oihK+Nt9gTgxnfSbeNr+OrSsf22ItTRU0EQyUg
O4fZuN43lf5Xo4FIxAEVk2M38E7Si5nIIs97+NaLOdo2w1KoU48oR9LXIkCu7eE2Fi2JvxbbtBAp
QmkrdUVzsMPRUckyVU5LtKzsP5I0yK4qy4g47lbgUP2bepWNXt0hy19NaS4wLF9LJCI3Zgb1vLvF
S32N4DJKl3fhMhpHyo/f8+rQmEfrc6u3UEzkT2wEc6OVpMe4vGp5MTT4sVF25jDp/Dex55vc3uno
qtUFZXY40S+0HazBw6NTUpxq5RY0Jlr3G59f5q10F3MalOeBW5xOu5YYPL+OCBTXk+wzC2oR8It2
EJkJoXpEd5rKJL6FHA+LFVhb8NKI7xSVRXT9ZW03fqrSfTPIc4PFOdYWrdQX/aOJj7WlAsB1fXs1
MtUTUQxs1/2HFIz0essDdrHfWHSD7A3IG3mYu/oPgOVjvy+7X1XiChVoN/5YsxTvQuLDWPRbrVq7
haLW2Uh+Hd1Hm72JNoAUzQCgV61aloIKqeqD171MFDzFlzvVAOMsfsG84fOLATXQ1OpQ7UBjWyLP
KMkNIgsiA/B5p/zbsPDzFbmmYPXpgCEJXLRYkEdYoVwDWm+HZkPu0RMjl5rWMK/ZuoPqTJXNPvzc
D1Cn4Vi7+Vyfbpwbfm0ldnQ0Toyi0bhy/5gMCNbGiGwgIUXpR/gp2y2qUtLLchccg4smSwcmxE56
Y0AiXL0k9qGJsUIQO4K5SdVuHSdxzna2cvNEXksRPhe0+89siJRccnOtVMvkNUl8fNC0bB0wq9Oj
wh0xL7AAKVaolBG0OG6VOvgq3hVdt23mhNSskmX+Vl16Adz3AlUzZEVVtu05tMHpla44UYcVe7pS
DfIlLpHqhMD6+Qf8zNAPwaCWmEQMBy8crJ5BDzjsUjYrkqcFud/kwMgkr4+3pvQ2lyHNTlS1nagf
JfCL+TDRq5z5AosUWBig9IVp4lpZFxSNS42c7ynYRgEL781VavVBE/Q1wR19TIkFaLC5Xn6L4BjA
b+0FmDrwvDdX+5qsAsTUJWpX2Fh6bPf+lNt10X3XdLEWzhax5FHxeHODIx9JsLIGqqi5j4/IBuXy
QLeZRrVwQvk/6kRDcGAYrpKJDqlYr5X6sh5kcuvjcc0MJNx/PKAbHQIfBQG3wZ8M6Caco+THRWvB
n/WlsMnFL1Vm7ubRTPinMNnTyU2A03N9+lgtkmq9ZlOlpVllxKsb05RT8y1f4EG9Hi2ecHOKLoGx
d9n9nbGza7tcj9C8PDVnR6r+m100128uIWmMbdbxGfhv6rjYeXpkob/qYSBqGG9FLmeJ1jogF0uX
DZ+2IlmwT9Wb/+vmK4FwTDKQLjlcpdU5PRsiH3bu1/kQzcG2P0mY9pA/3J5aZPslx61wK45QXZYt
xEy7SLmkezIugJTPZhZ8oRYXwLE5YHlSqfAUdkcxpeTsX0Rqa2BOqARIU5dpY9Ug8svpgZHiInrD
vdFUaKnrHAvaZO7olO1KGPp9367itklVsT9VplRwQm8d70qpxgx3nlfKvrsrIfqxDm0+I2Xwv1hI
dvWITrxd1vtFroqpl6Wi+HGlsDCKIkc/xBf2ScagmN2MJt22gH1YMLwBOaRFr+XCjv39CO9ragh6
q6kJL+d9ffaHDTtFwkpYOkiPg4HBYYNagZkMrJz75tk0kCJA7OaoDlQ/bq15rQna9eKXdt7Kedm3
H20qoRnQzuEyp1lN20IwGrxFcsR9uneG72r8iIHUHL8DZchrjBOFN9WqVbhgHh68SOZNq9Cq00hM
BDny2+azAa6JgVkiutVK0r83D5FbovJNmGX3AmMbEcK0mw7dpjVZLCVItt/0a7IE/KO0VNEhhWaq
EgYE3FDC+g03KpIE7sniSBZCQ6VZitftMGrsih5GUOFpVVNKSfSxzUcRnhLRwKaDAuV+y5BUA2x2
bqb5gAtsdFEGEYwRoyDNfIMlr4cf5Ra8toXeEE9/N6nV+FbkWon+ACbUZMumqq/lj63z//tv+ypY
o1XE4/UTS5UHesd78PTD1dYtOZf/3UJ6oQIOZhKpYY9q0LQkb4XA+h5TOK8nAWn1WioeogDz7K46
64EbrLVsTE162ck5qAWdW8fp4kTVEcAFtcogbh26LQmzHrMnKxcRBKc9zQbOu/CetLIaRYm7YdDE
pqGPKiT9tv6ynYn7QkrKmpgXZN3PsNM9gBdlxxo49/bkplgK/2Vj/eolFW9sNLMTaNZNDpOEn/gt
aA4+tWXmix/hrPQ0eECmtvJ8Ezjna8/dRr27IBPD40pUdPmGEcW4+C9nCucFpa0EzQtApIl1ueFJ
miPeoVHHJU2RwkYu3yMgng1dnmGgsESngkS7epGbYvzySybD3hWtwUsbbHItNESuF0CnAyAa7C6X
9zo0tlV7r6uBpLe+g0928ZbLo0VoncPskbYjxAaT/bQpwMVjLPMfTCZWBHro/WGNDQsuHu5h51Ug
eG712eZ/mjYZ1H+9k+iYo5YiUc/k/lDU0XM70AACAwI/XLro6uKsj0waE6DWTrXMiy+0u+Yl6hYi
CAoNmZGacTdfwL1X9iXF7/7siNQo93kPDh9BTS8sJE23Tewd0g0qiXnG4BCxnbXYYV+l4itGWBGU
OwGN7KYDdgDjQrtBQL+CELgPpskj6EJlqwHR8SHrvzYGbQusPPFgZ6LQwPwivVCQy7ghPvMOdx5T
1BoO8O2j7cJ/HJJGgwyPBfd+4zJDdfbkr6XQWK39yt/Nxoa+fiBpftbZO0GrvQ9XRTPujwVxE8HW
k5Vb9ks7eBd2heUJHrCg8DjjpzPZlFZAiXIJ+z1eaxYq7SON/XHguMc2nUxtPg2vnDsA4REtNyu0
bLFBQkEUgtv2GRazIxf3aLDZJdzHO5G5c3H1gsitFwBbUNsBteCzywaQWjBuVrXZ0yRH1IfEEC+6
NLGmByYDjQQmdddL+9xmp5YU+aJqaQ16XNuJXPi92cfaxiTwsuQCTyni315lD6mui3NkubyzMkWi
wyyMFUcif7tXay6K/kGonPmr8z6b7t/ga+Y8uaJvf/6jTHBI3UOSdFevdUkWjDPvSR2dVT7yfuJX
xzKYz7MeLOlxa/J/InC+KedZINqiFYngt+x546FgdR+P/HWLP3zSeD3T8il17QNcmCz4Ay82oJaz
KNgDVVq6oXldkdA19hKJ6wLzbeTNafU+03ldaNyQNGrN+DssneyylalhM0g6hQnE7AGzKaOaAfvK
YGv8C2K7pkYNG3ZeKYzeyO4NLus12BSNmiuuAAuMCAkss0vU369oic2YwSjMBvbzHmbGYtIUX6co
J21YdIc7LfLprSJRNsrrLQcf+2e8k9u9qvoGHoZtVYs3pz23M9sFAPaxQIdYFJ8vHIvrzZfFh1Sv
vLgipSJXj7FG62MDC6m9IT/zRwOe3wTPnaz0lhwwIhz56NGfpTfIg5Fr9wBCGGcFfOczJeWK8dJv
pYB1soGhyDkT5eitYeLz/TGhqAQM/7r/yBKLI6XtNVGk84AroI1B7EiHlD4h4oWRDXclRPRuNpn5
WaUnci1xeaLVcLCoRkJPX1PcJ+1dSo4Ee0pKYoozLKvsWKaeq+Izm3mARWz7e2TZmmH2RpCtwfc8
NWYVFsGCraqAKk86bee8TbeyXGX+hJZ1A2/P/vh74vbecOhVZp7usq/zZgQntOqAMop9b5eQvtbh
DeRHoMxnvmLpFQY9PkGFTwX79n9RnDOJRvBZ7B+484bQCTg6u8m+GCItHyFGGsYSbSLMhiXiysgs
hsfyDuyZOAUSLC3dhfELiAVKOrbPORBhRXjHT2/AV3VqkcrNms5+P44Qs3spz0XMh3aOHytlwfEH
3ZKEFJB7XyCTlPZB3Uvdlz+z2zZe6TGSGSrFLPhlj6eAYo86JFd3JvS1F2XGLtrdtr2XQDU0Iydl
3XodhFVGnF/j8EHH2AYOhj4CRpcN+lU4kcnL+bnuZmuCM6ntx7lgRESFLOVGk73Yy3JfwYkehn9W
CWYXslU9hyr7NzSa1WrptiTUGd6K6d6j6UfeBhGG9kNXGMb8y4RBez7TBRjmBtKSxctsF/8MCLw3
kILOBpjHgKYHjogGDrmtxfkKFix2DQJa5oNBp+gXe9z8xN5+4cPxrNc/WxjWTiHJranBFM74OB8B
xLUnZQ2iuQ420a4kUTO37ui5Ad4O/E2V1T5k9ZMRQ9EoavmG2LSkS6nvdOeu2NhC1EyPl3GOKYHB
90+LVN2Zhzen/Df3gIA1k3XR+HY/+TrCS5YzO3H6Y2CWORxF2Vm7nUTAo43jDOtIRw/JaOIU8aA8
XEwb4Lprnfg18nEMYE7rOYYgK0yntTo31v8KYEMS6/73tS6IcEhM0RUqp6W8Y0SwgsdG0ObwGgTE
LIM9F/rUEY1RoOtHGSdL8CWPDWfHD8+N+ZHhAvRks+oRoMNoYClMmL0ghWuGcjkoVDfTZ6NMXwSy
EUzpnBin6Irj+leThLpV5sEzyYTdFzkg+O/II4d2RkylGFjlYJTV9UhmRefQB5LFvF/jMaM5DJkp
ogfyWD0Jr6crJ2JGKWw9w6orG2KO9RMblbuIZ3vz8sMpyYWqztXbIQnjrWQ6FgM6REcVO0QUwUts
yz/umAMZ4XWHeyqLLBoc2qXrAg0Mek80tcp+5z0+yuZdZYHGtdt29JGpbeLZbvqA9u8hhndYyQDg
sl+oZYepz2ONq+nd+uN7TK/JHAxW9D36R+UCi7xBIkJKCyI3k+1ambXy5MpPo+q3PGvEFFzeH2MB
pCbsVlRoiOcGRbDYxHBYou8+ZHlJ8wM2H5u8HFrvFXwpD8nYXFxhEXZzuS4Ucd8sNz+YPLGko2IH
yd+vtfFh7DpMmrJzqJNqZ+EWZQyjHpyY+ZpsQb1E/tpParimtdTnPEvxgoJpW4uFLP86QMu9cKI7
i3hc+VN+XGrFsQj7lJ8sumvfmrfI5wDIq6+3l3LFJt6GoMG75DOgALQz+V1Ivw48UVAk89xCdqF+
JSeBrZmQ5IyHTPARgeoBvbJeALD8d0lYNIYgYCEjoDweRkYh3nz02ewLQsARUsS87AGGeHjk0pHA
gYxYXw27tUiLRkWDO7Gn+R9ScMexzAHl+3mKiDw0CK4fswj+9QFzoyfcQTAYPKSwk1Vlhr92ohI+
NqI5+TeKfNvSpa5P4l6W3gGbX2iUjHQsvXJHdqGNyz7nvFjEjrpfWsG+nJbrAlhuf2k8/ybZ9yQs
Id7kkZlKYVzO/kOX5yj6qotWbM3vXV4y7hRjyI/A6cEUkHMB5Y0XurzNt/OC0LT6RHVAo++X2Zdw
7kTLRpBsDtxqkwK9Mbi+b7XToLysRRAkI3Mc9lDCW8u872qYyAfIJdONpXrBaltNreNMypYIJmOd
cp+NTv6kwoGMYOk4izxAeQUtQW7ZmauNugA69QJfG8KnabMZ/oD0RM0lXpvOEUYP3M+bKNbQMmLD
tfVHFKU2IbHDGau+d8nvp5h8/Tw1YPc6si2cwez1Yn5PnLO1R77y2/fDu0vE0X2lbUEaZWpFmDeM
vNvQZD/A9o3uiosnqGHUXNaFY2ZWTjgs7jaue/Cckjg1ilndRo+XoJ8Z9+frl9qAqZ0/n9x0cgQC
knoJ6uJiDgunim1Rb1Zm0CNOxIM/ss6bqEjBXLJMCS0ZRObVx6zwGhqElmfi8W1BkkgGWBJE8Knu
br2Eo1t+qMUGHrp28OOaZbaGWHuFChzeNvDWcj0mDNkzIB3X0dq8+1dKJRVkczng5eBWmsgYjueL
81tbufH79/bYEhzorT0NuSLYjdHdY4l03/VqO16boNjuj1/+u6AvH7qJhVXsJuIp1wC4aVmmx4Dn
dM+vkkY13N3qXczLT203HWqeGT5t4VbKYxcfhGSMkG4od399eHZeV9fUGLAXDZla/v1z96hqxx/3
ZetPDiNfE8wGrXvUFjRS3a5YoR9bJOo8GshinJdSsPRfveuBXlXjXZxHy8DCojFdQbzEx3ZQRNQH
Ig4e9bGRmLXbcY1Qa5HUmxQH+Zb4k+Q4VsVkQ9FpojX+L4HIfojOFb0B4pkTj9XpaYbj2NZz3gCB
tE4blGQGzeCDFjixGenEf2blgCEkMCA4hp6Qrqz9MG8FEIXI4dlK4iLdTvuUHxucrObvE+CLnjwC
pwbxuz4Oa6Kx5JXEssN6Mt7i6z65Z3SXcRYi0OaRWUwWkHO9b0V8TD2nIUpwe1DPvhsB3L8Gq4+a
0AVSlS9QJ6fm67WB2gT2xgDajtVEktI+/QJ/oNryyder6WwSXfnq09QhyU3ss7xl9PTnjFPkHZsm
LUjsUqLRHGl15Uo0OZ38l3/jG9d4NPf0rfevsIDzTBWpX7IOTwwt+j/NjVEAniaBq749BgWR2oZD
Y3bJv6YOxOa3TIcjiIYeteLbJjgLXV3hbe10P+/0Pp9LPGWSOOWgUUN8vlUlgg5yDAEBsBfDXNKr
xG30ZZQsgAuL7dSEKOmzwYoJkMuMPdvqaJmnMs8LOhBfyHAaczk9+81fnMcmN/apWTt6mpzIfeZ8
cly896kEoqfIU9yKzucwldozPg6sj1hMc2u87Hg4WVhW2+XJf3liIvpTTjJcrGSjfs/BSwbIIKE9
+1YVqRcQtITQKthHzQDkhRhkUXa13cMMcnpj8PhyYt0hQPcxajwWUAsT6CjVWdfAOLChxEVGTaaD
tohA5OVpqqpQWWIoaxWV/Fitqr7x1me+aM9/2w9CV/SjqxrxZnV1AH+bhnrtfDuTEVsMvF1p9eZx
yv4YqDhdQCC3XhROjRM6PPEWiNQlu6CaaV/IJ4AEyQszFmCSHTAnOdjHtaw0daF9cApecwtuuXdZ
bD+Ro3dycAjTXi3A79dZrPYYqsAEjvKPcgGrimID2Y/bwzWitdb1rR6jfK4fdCD7IVT12DCPql/E
pMVYEloi6SIlvffdrEZ94+z986Ckv937O63Wpe1qM9l5XRh9bbUA8/AeYdbcOZlb1Iwvn9sirI1g
USeVRfbdaSrJtTp22s+PKAgpuxqWoZBpTh7FVey1bZxsS0uR+8pOZV1lEWXD88F6sBOzfJ0ds8R7
nC5LBzKpZ+GTmM2Wxa6ivucp8zpWNLheMYji1/bw69wNMjWZa28nauz8cSHt/i5TdrFWiVPvV7B6
Qf9/RnKgnFSImeE3YMg0Yta6Q+/Ifrqu5Wk1BF+KZXRBIAe51zreQTYsjPZhBn0m8Z5ZzQznmrjs
HIlxVdYr7qIQ3tHyTaoUwbOK4ZyTrVBayDSobWhCO0uNlVTBWfqileooZo27aSSIkQy6GVKVSlab
0gCI4yHXARDm9OWmaBLS0f8CrpNc37lrvs3z01XK7cfrZZWvCqxNnjYnYxr7VDPRqvS1G60ypQt1
gvBNyBWSKDSU+cDOO8lhZ2/ylAtrOuinPfI0oxKm2yD+ZNeAd5JgRsjauTfIzvFbadyVo5DwIzk1
iFXf+4zSa5E56iYjZWU3/9c9okxM1AOkfhqwBqlxp4rJ965PLYWVQHmaJWbHqy8ySn9z20ZTD90L
n6SXHv6c3yFWJTZY/IpNtxbMjvBKMP098vO91tNnl9gLntatwVrKve0/szJST/SCVA2XQzMyWeOn
iklCY2iiWuNz3aDQHhEHJjrPiL6C8kkvYCHoWbPIy7mzMiUkcwpxkR910Rnm8Txjx9BvsKZEGHUb
aC4TTPGHhFUS+DdlPf3wGZz4NkBRGwoLF8R9LGQCqAKyY37WOjp/QhRut6Lg1kn81f2LRkzqydjo
28Y7isBrz+CUGZMGvvC2ybOU2F0t025ISuWauEbvR5leQGAIeIe33juZkk87P2eV9s7SK5XqqR8t
UgycRNJsChebBa1UZRSCF9dy/mAGUL9hKmhc99Ij7EIQacE6zj1vTgaDwai71jKGy2ljT1i14YIw
IU6FZir71LrSele9l4GxojjhEoVVTfAwTaAO5i+yhQ911N+xWwqFy67JIYQgwfD1xWF204JbICnk
vhYtE644d5TsiAkY7YuDvA6UfrYIbAbpmJ/CGGnQ4sLcJSvoLJsX0gDvg1HxvhKLREmDV5gJnRyo
3KSiSAPZLldQeN9TCZ/J8qOtIqCBwlPW8FKZ9e0MXDrcAtustEl1ZZX727DlQSYtE+QHYyI6ZSj2
Q7lrpNF0ygR+HOi6w9lVmygNetamlLStnFpM2gbIyOvOa1xoHjRcbsN5FMCaWA/0Bd8JzA1DbK2y
m2V7tH/3rNeYs+HP0aFmvxyfKs9NnhFWVYaqnZcrOiTELA4Yl/B/X63Ng6eB/zbbeC/0F8jzpjuV
XwhTSvlS14HQQQDnNZMtcJJ/J07iAT822cwazI4RJgLRxui7k1iUDBkqVXUXvLEt4FojWkv36Rkv
PTQYzLBAq4D6yQhrUmazfFjwN9axEWfMPU38YLRZfkOTUjHT48EjZP8wvtp0mvpJIw0yY6lMzmT7
uDdbGtX9KJYOni34bnjM62Oq8LMDHjLIAPA+0zMXhnSM6KTNQoU1CiZnNgnQpC5/Qh1yHBJDiB0/
yheRg00N6lTjpcKH2JjArj1tooxcwvZANri9psdP6pUrgO7ObQsq6RG1p6xXYLJIempM5BmVpiQZ
D6DMkMbr7IHP0PeMkcKrL+OuIUzEM1t1pDORan7nk75vjy0C0siYaYp+sWDWrpa1XbfHD0gpd65O
Igqj2FcZLTlZnUH0TpRiOKOYcDQM758ckhjD8uQbTfSg/eGsujgcpEReDzwqfNrvhFAWU1XQJk4W
5o3+N32UL0MKelKRJQJXOzkj96ZyBGOwd6rX5ViWTRxuqQvt3b/x3+cUal/bGFO/Q2ZLy8d0wWcS
G4YIk3wuxylMQ/hhHWKWrAgcUgHMKab77Y+37RxQ6I5hKk79xhfqMAVutbtINwyNOwjuHGtfzC4Z
hWIsQpYdxQey7c91X3/LVatwww5GJGJInV/PuPAGrtcO6DKi0wrEMbtpgkySFBAoakOy1prWngLG
sTFt11wlHx+WNYk/aIg5WV7EujivcZNP+HPUQMZ14xV2q04PyKEg0zPQVPC5JZN7dKedJaLeY2AG
Z6iF4a6jvw5rrcmrRoIYeccX0oe7XtL6k15ahhglDOJK1wEKgbqQ+p9awI/FV2Sz6LeGE1DyNxK9
APokhadDZSJn6D8SmovVZFOl15V8g2A/2/SF4qwmIibmTS5TaDBv4U+YYOL61INCihlp4b48WPtf
W0hVo3pnkW/FA7rnB/apALptRiQEdOULCZO2G4+AzfgxwDl7DLAsXd/cZZwYQNxJR9ttwV9E/YKU
JaOT0bts1+CsljEzq2+/bsf/gbni95dMjX0G0cEVjS7F2h8RJ6c87USoo6ILeaY7h6VqgeE4Rbpg
ly638HDeBLV+PcaBHrBmZfYkJLYiB6DP3OrvDIia2Yqg35Aj60qQsUjfFz9YXnWF/u+h3Uf6X5uk
7XaNlOFBIBLuXmH/QSGJsRgmf0iYaWeWOYGewu8MOiN0eL6w4db87wl6JaebQXuSz7G85x24BhQC
vGuPnaq8Z6gI8NYc0IJtldbveS1IeVWsyHq7JuR/Vv0SE7/cWxbbOpgGNHMzRljEBO4Xf6k/DhAt
MFek3ko5zBUMxrPqfTDPiinm4Je+NfgaCqZ6MqRY59OfXZcSbhQJ2tc1/CJGakyHoUeVRWdZFaYB
7LU/A0gTdp7f7wg+Q5kCp6mooOe0RADuwIXsWCV74N3fZpxzmFvKpLWQF12Tbs8lOrLxX1WtTX3s
8ZA0EgZx4R9wHA2LduC2wT7QeKNRIqOCu57Kp5JaDEa+kz0QnfxyHhRMgXmEVQ1ulx6eIrBWJurk
bjMH1WKKgYowLjuwMahgWitvQWLUj/GDf9WwpYXt4ZqetYA5UOAMJwSIJco8hy00xrdy1SBbs7+F
8BmNXaxaKXlPhv5VhXJ66sKuXmQ9Z/7ClqPg6TomrxBxE5helzW4Y7k992pNLG27ZBcnLDYILHh/
FGYhDiHBOAbDp1NFHlwX8/lYaI+yX6MOwrm2ZmNACG08dRmeS3N4VtFF+FKViIU/FzOeaV+OaWGA
2+jlUyUYuK6bMaiV7viS5XcMxhYbACM1NhJy0hpgHRP8bv3pAsXEyV3uuEaEPGR6hVKs4c6HBdVg
+RkXiSv/XLgmPpo17l8gIM5tLSCeX1QTH4jrr4csT5VDBHEFj9+SaUK3GrYAVPtNxJknegZK5TKg
jbtnoLv/39YiSBSmwWRSR+2V6TykWX0M6lnZ3kall2bp7Gi3ZEkgraYlcBWy7RqcJsFVHP1O+Pvx
/1U8cr72aadSN8txmmBmGVkDDAzt05k8HNmGDL1hTYmSXmYjLMZOlXXQ2u5JpMFzokxKH+O+r9pM
M9HwN2GKom+cphmKac4AXzfa6Lrub1zpTnQFWLR/ZAr1oUjTfRs/0K0OZA5tJUlLHxhL6GquofOu
Dr5wSebhEIeIDPT4OeB+eDAcmp2kRD1mjGOphw5cprnoWeFL87/Fwg+Fmv0tpDKmc7yDlqsOuwLx
FegBQMIJOp3jUrCZYuDGJ5h6ULSwsu8sTBsU1oCj/PR2JU/+VHgPNcRkIDvcSIjmoMa1vD5ednZW
NGMVEojsHoFVFWo3bP7sgOSgbCrNetnBjA0cUCztPDr07vVKDYmCqqKCPFD7Iw5ZBxKZ5uN4y5qY
cK5ZiFhBFdL8NcAegFwuD5BlGfMKKLjrie9W7p5vttWgx5myqhz9tuYVGIbP0/EG2E4UoUiAJ2HU
Sqk69r9TCMdsEGvZgMoH/S7d1XsyZ8PzhZYksBSaXEGYTZHopqDA4ZWIDMeUeC19ASp7mZmEhTQ3
eXUjexTZ4EMCRrokYpjpkHxGuxHqAX4kRaXk+7RZBKT+QnfXxkl0QEIDdXoaGswRKfTCnqfv7Dyq
v5xjA5/BXP5Ni2BtoC2hBZMb/jC2YINna5sjaK3BV/ACl5AJnDwL4FuhMm2QvsFPjoWhS8AyY264
5C8zjPOsnPQXN/wjKxBxNf/Z8LrGc5XN9hMACbOqM25BFoNxCL2X4Z1EyuAqPkNtdEGqFC27MF74
geVG/lztRmIyjuIrpHnUAlOsrN+rn9QhTd7U8TQ1szWXSwdnH+NAm95V3kmiJmSbY84OwJnbn8SA
v6nCYlg3p8ZZe5cNzhB22Bh2Y1gy9MDEfsPk+tmeTTPpP/9V6x++YifzBgkjVPbhdGPc/XRX4SaI
YDEwfmJYFMgaXO3UrnJ65FuNlGQLYTsAmXufEsGa8SoVkXPO3TwcJLRn8WMAT2TwTiw+U+a8qHyr
0nLAespBcRNKv5G9lk6sVNsOMqz8url/RjFfs2H0QkypwMLEUmkkdb1hGfQcFzME9xikxy1x7736
/wg+BO58eN1ZWjkNk6Ug0lBCIWfpWmKu09DUQ+ksms3IakdYuZhu0E9r5QTVmoP5Ep2IgrhUMHGI
VOorRkaYxUx9giPkD0H2jITgqiKn/TamzAHfoUFjbLbtg+9VwJltNuYXpyyedI9ZMXB50Y2IILoj
IriFyKA+xgE0e0xqKMwNIHtqePCUdLK7XCIAZMAjunG1c+LMleey6upaJaLrKRvhc+uiDbB/SIUm
bfWSYW5VMpwVMxdsKczwL6plbsnoXjkeuYCoHkfA62vWsR/pNn2D0OvM6n5wHFiDSANIcyviZyJ2
G2Pgtcz9qrriagFI6Vo6BQh7omSEllhj7zHFXXPZQLgfh+d1Vi3o9cq0TQ0tvdJbqvwok6a9X1jh
9wpOq7eb3zVOrYx0hk1l9ea/rO0YlgakGrr2ZNb01UdCeUp28mjQmcvSCmu1uOKmNnUw8KZoRIp8
ObTuixzaPRoYXH5oMs5k6EAjGQwtHbJ8D11DIX/WtDX8agBVUrXYrjINH7CWbiPmL560bwAJVwM5
iKnYtuJsc8uyjhXmIOAlmK0gr/Rapg+dMjyxoYMKc7xhuBBEErPoK+73by4UE/IhJKscoL3DWKB2
w+6l5gkfQohhb/1SLxEhCrQOOTUhcjT6ViRH7iTM8BvlDMqTaS+Jf5RtjygcAqRpwIBLPqjkkgwp
GXB+oG2ZNgdGeB6O3XVRu0VNV9NUXYl23RGNqVsLKXYXuEII9BElOaOMoz1v/6lsXVJ3FrHidR2M
sMyQuuUDftf98oeJbIy87RUnoEn4Hq/BgMmJx4/DJUvnbAT36Gw74dDM2MS2NAt/W79bATSZuN3J
6249ygtIhQNnT4T9cpU2qo2riLULXbXRUgDBs/FCPEeV6uXRhTddhlWizYW7LSVir91D3+o9Q5v8
sZ660HG36W8T6fFUSBOoVDqO8V/v9qfkQH3f6YwZB5h4a3iEIbQcqPtNgF84es+4uMzYDc4xryHe
d9kjSo0ce1zhFjpkuBLVB4fxrZ3U+CXTg1Yca+BIysqyjdpyWlk/rYePgztO6QqtyPqJl9DpxZut
+YUhDFnOY4llbAgvmOlR19V8PzSYUIBODnCaKRmMntXPOzqPo2ImxrWzSa4jR5EF6oj8jn7Il5V2
67eapoh8gUo9ynBMQdn23t52TBAxAiMEJqAAuWuuvqPWNkGl0GwHXNYnKzBbcyB7WfJbzKsDKJ23
xmaXTtt3OdYrWcFkHvR0zb9xvulr4YPZTRmgmBB9637mO2fDVB3VFRCAEn/gSKwlSVoEfOo9tbJw
Zdu7Q1azTM33MtvEGJuGq4ValNYPUb3bTycFm4t4hicvx29RJ2asIAuRZsrpP14SIrJoLKXBVU8v
ETcDPhil7zYmmqrq4SXpR7yd+mh/H36gyjcU0kN1gF/1sNF8/0yPxC6uUzBNCkwaewx9ZYg5JjBE
xtVpVSq5SUSbLJAL6b7fxcsJWOuuEqWfpevRwRHCZZrxe052xqkn9eu6BWxs9QSjlBHdbkZ+PSVD
tmK/JlTWw9F1C6vaEqcrmAlQQgYnwqMirLB01sEy5XJzlf5vE7xvFoE0R+la3x9vNCfEvOFVRGj2
mnJ+LfcMDOA/3kQAKrd3x3ithK3hpoSUUt3dDCKxd8thnUhsNg7L1uP8J221LXp+AGCf+hJjW9Za
SPDPsYwnuJOc8WARL+aQdXNfuRyqk5TTzdo8bso9GhVa9qPJo+8NmSLaERB3q9J4PlqPrX/CYn+O
obMzVPcu4NynTkJY4SewXi/kHpVEv9Y23ZLwkdtC9bAHCIMlMhWdgS5Cva/MMTkNCk0VyJfA5QA2
XcxUvjxIbt21an4seV5zrHwNMBl4ZXBdn8RuMgTXkYaI+8Xamwe7mwKfta2s3uUlzTZ/3DMzCJzm
JJUIE6zudeFt1M7i+ngnGo2P21c+2qiWBT6XCV+cD5dmCR9y9mMzEt/GxKQ5yRSiHk7V+eW4coXm
HcgIcvJ+AMR0rPYymb7CcLU9qZ8qaKqVxjnm6OgFRlB9R/s3AUCbS4zDAaH01UJ4MBIiQnWV+3xk
2TufpbCXfmRP1+6TlvW2TJev+KzhEMaWP9RieOsg14xV/JHc128PCVVeHCErsqeEliBKdb+GlQsb
ACKoSF1k5sPgObMq8Tzfe+9iiZVkMB+kjz0SOgB7xZwM+ttJ4k7vihRg77ciLkBzSkyK5PkSuoge
qujoUzqIa6J+2wCBuIriqV9AKfOrW7Ne3EKRUCPfM7ep05oUZJQRusVouLVKhshOduUrp+WPvc+z
KURSQiU/XGfPZhr0texytzQrXzrGmS288VYHOPz/NZZnK0/sovLfpMg4gYYsYEowdkcpww7dTZGl
wOePR8RZId7drbdAUrFyWOuhkYZh8YZ8AsBSzcCS2pwG1r2LGe0i9q8S8Rs0pSPMgMshx1wbnUUl
DCSo6aTHqnbX8BTH4eXJXJol48nlpi95mxIB59BMKkbdBKgtuvsLcs1WTTqM2QwvX8FmjAtL24ww
kieV76wKEO6mR3zG2n77viw8A4aMKpi2gHeQXO52VgqUftWeOvpMfXkkUjORE5XscaHEkRjCSoNj
7/Zmx2Fc7ftHK+7BdBGKR+1d4JZkVUQ4JWIFTS1Y0UAdzuDl0HbFUUux4vU4V/6fz2mzsTL823nJ
uKiGVr5uJQVMmWxNPBv/9C+MY4srG3O39fQV2lALYvzY2eDMbuwjEj+VKv652x8WhBNeRZxSIXPw
0ZY0ZxikJ1EW9bD5HZr/7Y+uqeCEiDfh3A8zMV8pbgRkjIZgj97eER/Unk75SAlWagyJHgDFLO6R
9+OSS0RONJk12NEGNEuON+WWmQg/MYfmw78W/fxpGM/zmaysZhKdRWz5LzslYx/08G2yGMDoqUrc
/LkPpoQQRPbYxE/L5FNWGuDJRITKGcJSbv6Oo+BUnHRIjY/2w3drwnbkkJ1wzIXVy0G1qigwZ0yk
sUJP9i+umco8stsH29K+SlU5pqaQgl2VDxaWn6hbxwKtp1feNaJ6kTHGkKOdtWnjvFGuGB4pnCSg
SU98aKpGwWg0LRUhmlZSH1vsMvRc+Z0zDpy7PlTa22kNlRVjYQg2aBZZlgp+mfl27sicnkJS1F7k
e5oImpvB3j1127YpgrnwdqVy034dIxLsX4iST1fsLowNrRQMvtAXrD9d8y8cHCNv/h3A7kbzsMI1
wBZ6GGX0rDVVc6kooNN7v1RDbtIMEL8JQC2gwAojgoCo7gN+A2DjRZ9w2JY1YGdUQMUjoIVGwEhq
XmqBV8cG3wjPNeWbYaxZ4FcFIhX8olvKTmD+2HIMvzAr6u/NdvSbTu83r6xuSC+qBSsqDLDN2wlI
BdiEVWKZeqbIC8YYr3DnBn0PTq2A1QurYbJzrhKNl/7okvK3z+u2cMqtqneWe8meQH01UubvwDkQ
UPdZP1vKZwjOfkqPB3isxli5dD+cBaqrRcJ1xPLuFOPDCvfrKaPyrVUEGdAtA/YwqVXekhnMcNh7
CW5+WWLvi/xL88UB+ISgaxRwiDV18IGxuihw8egH5clxFCsw+cJ+IAaGMioeRf7zJssBmQvnm3lQ
ebkxJ8mK+hOuRqPrq5ZFppOatKUEB97P073KuoMjTlgMoRQ273BUc4e3QF0w6sGb29o1GS5UnQ8e
F9H556L6IwuL5QM83s3VQHzls5Q7Twbxa9qa0oSO6ziiYMfYAFcDc2CEkOvMrTeVPjQSVq5NsgGY
mb4hfC7kd6u301LiSwXoVSGB/bV9ySuwtsZh5+SdCrJ983E6V8bafo/awZ6eK7Ebc4y3HEfI+qu/
WUYrxF75BtqPW53PmyMccmAq1o+BJcBqJQxFMDX3872BZOLIWeGUuSlu1MwTn3pUnDTaQfTWAnNY
5n1HKN3Qc74VXl0eSob2FsSELNtTY/YwOfRn5RG9D/5Q/771+ID4dUKedfzSD3Wp3nnoU7HmHrZT
Y4LOYwmGIHOc8s5wU/RaplKff4i9DhrMeYxxMAOTvQXA+bH2tkojSmLFW2beLdVY+rsaXfhPpKvv
LCOrEDjildvWbWfcBRf4zscrrTmduzLEGoVO0mrcNs3xQfNF/5Z3Px2DDYZljQ9SeqFiHEPnlx/Y
UKGZvvVuDaQIOXyc2ow0TbxWQlA0ihl7euJrQplktOTULtT5Fe++gtFuapZG9EUAjQFYTQqq9Qg2
oh+ZWYne40eD1DgTzyX7ClMJClebXV+PSIz4+N50UGRAedUZo38t6f5zSuKs47FA4t9ErA5YjYeq
hw3gyv3Banr5K78SFVekuIm4Mq+6Ykol7miK9InbRtGF2WHQ1z3ezLO04j8bZOZwcooS1LscFl4E
2tgBHOLnD1f8vZHZRGe3LnKQ77Wo/k0/+Lut2oNDrvi21fB+D6Ndr5/YP0H4QkVhh7ruGa85VVPU
YxwALAXWwsZIw5nGfXnu2o7Xs8mJ1uCauhJN3WDgrk0f1/nyCFG0pBuPcPs0D12RQTLjSIjPq9ji
rbV/A82Lb9BmmOBJ7EVGu7RlS7E0jcsUN9H3k4aaGD4j3THX7c6jhnVy5oGHYfFPf/EoNCGAFNSd
3UAxhwiwd+E55KKgTJ5w6DZL43iK+/jQuFzV0X1qbLwyvyLyzJzV6aYhQsTu8EXQesu757V+qDmj
nQ7k6CGk11AQpmNaAkWhPUqcMI6ZT6/vEqTfgwVwWRbn77QFgAF4s8W0gM4tHTJLPtrW1rN3TCoo
VsSt6DceBhC/JO+2O2HDaPfqqIqhvfEiff+eFNyTs0EfFM849uSkdCl/kjU6Oo+idY2P2QcV0wLM
VPnYKPyEmV9mGQDY5plooybxQITo4+GL0GYdl2E1R2QhxlFWNgBnIX63EsIoyulsBDXsEb/8uPcj
tvXI42FSvcf6jdg21DkIQ2dQqnFvDpmpyTVNZ16Hlwl1E0/3iCEKDVKKlx+H73CsH3+Sbu/0ZC+v
TiK4bQN1Wq3n6NE5//2wX2FbbJ0RmXHLMOhOA43jPehk6CCW6254otiMdnK6wgV1LXCpBoNDsNi4
InvF+esTozZhLW7zxjzwtHIMoh8/Epzf5vxeY/TWJogexErieO34ZyOja5mGedDA3l0yAsEcJv9+
0rLvyIOan8MLSuITV93lr/BJFialZm+n4BGdpmu9iGFckZ/059VSwuPl12tGRrf22rQ+DUflejOY
E7n/k9Naiw+q3Igz/LzC3+9mtSltpJDwJdmCKbfur9VpTEPwSVOyo5ipIojC7R8N0pYc3D/F/c33
AGKW98XxBops4nOB/nrp9Bk1XJ5pVSKE724CQOfk07dzCHb4DyEgX5iomqKvOrGuYaGpVEO19+g/
o0H+gDsBg90beAik2u6U89zA9Oi1Ffz6GpUusMRsP7MFBdEG7LLkjvgpmNTePCjeA+B6iQR82mAl
L3ywtosqC6gxI988ky1wWauiDcqvOkrm12VfxfPfAfHNSb4QiAvGwJZUpvrH6++C7BQIyN/YkKG5
MsECVxBuuxND6v5wO6pk/8vzIJe4OkcKCZQoN1WZUofL0fKVZtW5a/yf7Rn2bJt/vXzy0b6BJOar
QR3ztyQwHNBvNyeQsOSRVT6fvGryqS5Es3tKbyyJn+MIsUnQBxq+UWoNY0hi3LGls61FLj7XH6iv
e/sStn4vXZmItfNMomtVwfespHTpP5YAVUFIfrqE7z5RrpmvlCgCrhWYjXMjtYFM9AcVIEUitHS0
R9I1IML8nDjmGQSIu7G/TMHsaStvqiYfTjJ5AR4JQj1uj1CMaRMQkTGpBd+Ksc7YcLmI8JDI7UT+
ni3fPuWTbTcJLxrpNqpQNKzdet/HmY/HocIZC3xshenycldvX0oHVfQ0jkw26Gt3tO0BD6wj8FYn
amCSTn5xjvbTdgQ1kOAiYFyyI4Hq+4bCWz5VOOSA6miCk1j1EUMxufWL3XLn6y2YgIkEsYdBz5CG
GLdL41BXKjipBTMbwEQRlEtpIVYRZhhF0j+OYpJ/lDIaLjrcdB5gIC3y2hj5voStb3QZZHfCDuJU
4xJVGVna8l47l5FRYlwcTagcfcpYcFrpa1LLGLS6WL2wBjnzAR7MPHiAh/uyXe8LpjEKYUWWqm56
KnM5xMQMzEfnIITIPoMJsQ/2YNGRVH1oxH/CLHCAV1YxWBTSGw/HAACmZ3jtR6lRjqQGbSOD9M/m
jblig9OIokCOLxVl94TnyfBkjgL2wQBz0RdjS4fsU9vFTtl36cy/9lSx0IoFPq3ZSVeLykRzhp9n
MZSXY4F12MukfCGIESxOUFn5CSegNhnBVNrJpm+LD+deWKEtPxcU68XBkyMhDblmajpTFS3Pxzip
/0d8u89pDYVUW7BsfU+aT197SzERm7s/kD4e6Acn2C9O5Fdf8IVQj36cW075urd9BvUNoaTsyUqp
3EK82i2slE1oAIUmg+hT79X9rE4YpLsFqghQbqpMph4KFhieCLEivOcmmvIObIQFJoUHLCBgzcA0
U4KZv4AYgckBnuUd0/aPt2phKPGGbii68EhK7iDzjEdaJLgJN66JYWQCLOILaBpg3Ij1/tLGHDOz
2T0/nGHVBGCg+Km63b6GaJKiLNy3HN5RZW4lSpr3Hg5HR5qvbPMC8dfvs3B3kRiTbvQvOp3sn91o
7TzC+RvAGvXw/Wc8hryyxbvePdP/G9Hj8FLmZszJnuoVxIdHfiux/HWg5+Z6QftBSeSyT0pVNcYo
EGI0WCa8rtHJEvmcoZh9l7S4EBKKZtII2CSeYdaZlnPkmzCxdf8M+q5Dv5Zd+pS92yL66HOQ1b1B
WU9tUXL5+1gG0Mh/6TXuslkvZN8fErrnG2ZDs6Dl/N/UnbOMQYUrgryBvpE+UFl7BxAebKLSnpED
BmUiyoe+GMhbeWfXhB+RryzCsJ6btl+Kbo4j0j9pHHEo/OQocULEKFGUHigarDo2avSpgVzeNkpw
yPDJeQr7liCrBFtBlTiP2IEE/ZlzEd9QiP4t+qSeuarn7yhjoOkA2hp2IsKrFISDSf5j4eSVRM3N
zFzKiaHoodORs9Ga37QIw4aFLezU+q/uGO5YrSBG6r7mxTQjAtnKsIgBWxChOw7aSGg9dLaO0iqM
w89SBUZjQQuUJsp2SuAPIsFrtFQZ71EEA6GOAd8JLm5GvkfgYmVFSLIVAM6vhhDPrK/BJH4UICF5
hJN2s3+QzcnBDXQ1VnlagtsbI3IjRcu69yk2vJ/qmGM1tkoUYF9eikf70Rn6OBFSkKL4THunP1b/
P+vDXPvJFS7U9yUSs5bdd5/yT1Ug7b66T5aNuc+LVbKaLiRu98CA4eFw72DbFh+LyjLqj5cSk/rU
2uJvy854FlWfpXIjobjU0kgkgoKTLx8vKO9AQMrp1JmBjDdZq9/YoZSJ/icI/1i+7R0HiuRJRaLH
6S72VUSfZ7wGkXqsHaMO3KFPVZMvc8RiGPTffDFbcc2mg9Z11KndA14CXNFam9x1sv/dr0KlWTYl
jXJeNM8L86a4wN2oWyg5g1v+JGhakq5v5yt5Efy0tCS1cMDT0PE0Tbh8v1tr1nuFGN6oPhK6ItBc
bABqQ+WrgmJCrjA8bQYZZ8EHg6+Ca5OeQkbv0smhmJ04ht+8f2B56edhUtwtqigLWACgjIHJ1SR8
u0SPbFOPDZMeoZ65TUDNmCV982g+uGecVi5KcA0KyawBCYYp0ApZNvtsZdmL888W1oMDNcQpE8Th
sfFrbpFNHSwc5GEAQdm/eVl+tGXQLwarNJbdWkw3K88iQAQgkDdl3Y4AC7OviPf1zUI5ZJTNnipG
+ZbKZ0fgK1gyiVMWUY8o+CopVbzXdUuqyuFmZxQiUyMVyAnLfS5EkyVSjjnZ5/oQx1y4o6xuehsv
nSVLnFfwHLH0/E6jqvmKY0W7cuESaSYBVhnDEWjRrsTQvFvk2uyzLcpJblRMYJA9aQpei37EmF0p
Acqc/g+Xzr7SJtyZTQDZYKjACYsBsDqqRRjEoBPG/TzPHIRMSrTqGjzP/SsDbKh0GotcXcleXEV5
9LSNr4S/pXGcQKqSXl4I5JEh4LwT0NlFMWFKmuH+18vM9QSZ8nBJ1BRc4m7eG7JvtXUYIbwOZ0cD
6SPcTIawoIbCDEQWClJ7iZ9hNQUpJydtjI28e1Q+3iOQx9Sw/OrglkO5BGC2yGRI+qSj3n/s/zmN
Qxqb8soHoG6Pnrqk43F6dxY7PKwGzDHw6DLGfBUqto7tMIB+5/qiQ7xjjzdVd+DuGoKOENYazQeh
AofOej+CdzaMa5DEs550w5CyWoDGXoLYqiDPc5Dm1BfMgdmohd0+GIUoswh8drOq2QPNCZnE+Y1W
to2ZGgcDxQLuFjIEYt/fYkXuVOtBvKlT5pbhe+a104sSBcRq12Q46Slw/0TQmqjn7M7n1z+04TSw
AICf8i47xoduVm7+rtoQhpntqKXUtb5wJg4Tl5oPCRLxJdmb9duKR5/ZsKc9R7HZ4YDjKcDjx0LE
ZnL+irV03pAg2lWPIkk7u4z+Msiq+uZOy5S5h6vmffB0ijQvOaJEQk7l13b1Buq3PBhRf7OqBgOw
tyIQcImSRE09J8/Q5Di34OedtpHrF/Du/4VGWcc7CuWz/iJxjipZ66VqVBfDA/AH6Xwu76rrHgwN
Z3/a9t4Vb1mc/gNUgVkjIS/YkUexCxVzl2SyMr6gRIHpcpC4u8xd1zuB3OJrDm+SQ6yeqaTOrmlK
J6gu2454U19mgG3YWSc8aY7/zMd1bGeRnJpokqqpsclr36b57wUAeFoh/nNi1T+TbhFZcjeFkqI/
6dMMtCyd55QLZgakGa5XDRAGAruiWAiodx4dkWvi3/3oEPq/ayerBsP+0AjzPoOpblYzrfmYL7yA
uXNtldAnK7f2RKPHb3EzZkzOx3XQ7QOFPIrCH8xH4NN/96qhSaz9v++qaoQ20NRugcRijhZ3Gr/B
g0y84dhdnvlLPML/m53PdSHBNJ075RgOc3urv/e5gm02obCgoyzRsDyDARqfjkSWE7g0zLIt5Uva
nwRMLof8N+1PZwfQlwD0Fh6Gy4gHxeNP93Ili2tfU+gw9VbGBfKCaPEc7ffj2mAfZhaWccjIKDbF
656rTn92R7Zn1dx+I0Bm8XDv85QpPvIiTcen5g58z/xpWhVD1mjDatnp4Y6ShsO52LMfOxvfGvBr
SXOh8wfquFvXCEw+zHD5aF8e2Xr5wmQTeF67f+vIfXt582oYnDdll1gf2ApD+6Sq1Nknksq4OfFX
sm8UPCv5zYfLIa4zvHB1ZiGfcnyUxYhuoXVBg9VPFW0muZXMHoAhE0+T4Uh9g7mt1oX629JK5fnM
KnRATjHoC43OmPcuS7poKtubL+cNnSWwS1SEUjqT/Qy3BcWagybu5MU6heyyxo1AHAg3oMEu7xUW
exutWHLEmLuF7/bd7GJeJKHeznFeSJ1HWT+sOlROnjIBWIjj6Pnn2WAb9n3j3Qklt/hRN87k2yOE
htr5HxKNMAdzxRcmZMIXLlm/NMiiMzMHn3MIADgc4vN+kCECXx5aCapv4QncQg6iRx6/2T9NtOr7
iqxhPq/3m53UXZ69/nSzOPT2cyBCmZM9thm/K3p6NSm33T5FvF+qL0SSaZD4h2QYvq+0gorBmmbk
rgBW5TdscXf+MAPYqJDAGMxPXo153AnK6y1BQGfwhV9j+n5QO3z/SOaclLN6Wcq3S8+9fl8vZ6KA
rraX9lO0jKC+lBKGBvIA5RBa14A+4Tm+rYpJa+rr/K0Q+ThOgoxWgGzXGyt8N19ZStvFFbaNNagC
ONiWvRDMgUHwY88RNAM5AE3q6j/kWrdOwbxseS3AKMAql4geCxA+msvd9IcpV9jH/o3nYqMqPFX0
iSuh/wFxAnuQkU+pwsSh5KpmQylqQYthwqLeew9uvG5O7IGzYMVVNbq35dY6CrsiyP5uJ/ECZsCD
q1RT0JUasg/D5TNTQIplrJZcv5wIeJ7OKhTdD32sFfvz1dsVV1xLrLd62An6oheZlEYgSsfdVuyu
oG9+SCxqulHpM775oZB+4qEJPyQnM5SXXuLb6lIYlNuyEdPs9l2jmRhPFtpue2+IvqQRys+rUCiP
lVizo7Mj3iSMchrfA4MP5X8r+jL9GjhTa7TYOQ4Dg4BqWEV8Jw5AYSgGG0WAks3w7eHV3gwexAoq
jo/yrqm+YdnCPADJ9P1rmuA9Mhu5YYrQdse3kNfJqV9e1+7v6mKUrWwJN0TyI36L0sB/Ap/LBruJ
kr/T/EZcnp+kn4tQrQOYoKagaRA4WzFTBiMom6lcGljEC0T4M8wG9N0Am9aFLWlP/1xR9R2K3iBr
OAooQTnozBrlFVWBo5Cxq3QIuJE1IkHaSJNt/XOgrnqX59Sp3xy547msHjNtRlK8/QFNX+WoI/By
5uSrOnWWnI1VbpTpGcCb8yDgIVrP1EhdeJY0Bm01hMO/nwr4vgPmRLrrrO6scKIBldmQZawUKDg/
YNXQx6jbUnTLgQt2BfShUTxIrq2BQ4dtuBPO05YtjP5HU3rMZagtg3tgHTO0cD/kijkd4FDc3EM8
Q5LwdeRNgu0eJ7L67DcaMTs1ugAOXlDs1hgEu9+h6kmaJqBSKLrdNh4H+HXn/BzLLhKND/wWjRfb
x6p0ErNjumyAl67cXJoPmUhMrv5O5PaiVJ/xiI4AzSz0JdK45zpF1p2P7dGP2FVi7Was9T0L3+y8
gPpLZb9w/9qojv4CINnTW0/4LOARin+um9MEe3JawzktLPDcQicz/soM+hip+GAMia2Dp21miqXi
Yoe3mP6iKuoswH5RUP3HZJB/xgQgK0fGwVGcUTN56yRvuq/eMNF8tmRbaRcetjW9fHA3222mRRNt
ZAw/xy+lecZotR+blG/tWjrnuvnSdANjFVuujhBBsrT6eESOt1Q1u/oIp6xNloh09iHcyp6XrSI6
fwKCQlp562cJ5zzkTfcEtIOf6L2sgJpqg2uhGCXuePte+E/sHeu59hx2Os5AyU4wG4LQLZeH3MGv
7leqFoBr848e2TVlY84EWc3z55kOiNpi1fIezE7Z0mYnVmzZu6YaPgnOH1LOlyoV2XXRX2m7g357
CWNmNcfAaAa+z94Fw/tA6Gdtkzu78ztC7ikybys8fT8rnEzk62oCbhwMIRDFEHBHLwJWsxUn0LYP
nYh1z2ZSnn1ijZ2oq7bowY7AYt4Y02tIZ8M5Gtd4PtgZ0zTcIxDQxzHmKr9jTxUbl8pXxIO5l5Kz
9AV6UP97N5VkAZLQ8oyewKLoeYWAss6IMkm8UGRiugNGGWKEycHhEDYmMNWVjpStmUwVgmjo/ngK
Tovukl0Fi8X+tSAkbYkXSqe9mNEi3DCDsvfbVmx9JdAId4Xm54lXwkHnR6wv3dGTWhSbUVmGzJdJ
AdsAFJKLa3KqkNp0hZdquNLWR2Y+pqtHu1dGQwyQPW6ykh8q19eeKn5K5h3ANCHJQWmHsCg7vb1u
sDnHKTxhbHdJx2Y6lE6yjvW9HVHDe/EAhgq4po33DyUkEfBBZILNnrO6RLR1LyjqfqVJsDbN2gEc
ONtJ8FM3jHx+3Ubvo2fTRxzSzCGM7SjNEoLgIcbpi7yl6Pg1+VkxTAoYIjXP4EpEevYGCQSTp3Ba
vRm+u/LLSCrIQ8yEQCUMM7D/03p90bCtd4TEVZ97FkoWD1O2RvFSq5JwOmR7Wqet9+aclgL0s9lD
xtv0N3QpOeIl4vAqtalmobuX5WF5hxeobqv5zIaki/tHgGppWz1BRk72NJsBff0cI1/p02Yxzm/B
UEqUmomNnifZTX7zIWyUJXJpAcXXwHbSrt9n7aF487ILXvwFP2AuxkZbcL4GwZABbZO9TUBKz1OE
WShL94Rr28XbUxLdvOeMP1WE12RqUvgkTrK7PTw2oLTFPeDCI9eAUkmORTx4WRtE3jJhpb9YULFV
+kOgCyE/zNH9GjRs1NsiUidyqLOtS4lHlbWv9oEw3gh4HfV9BS3+nxrQolE32wI6pilFToERHUZ0
v25OQDdPb2A2oBJ6fO98j2tKaEV16W66wGhQ8Y9C3jjXHlQWalf6o/dnsJu/qVxU97yiYAGZC8kZ
6nKlkjFBfhWAxJ/HQBOpwLLPEpHf1xdDfvwrS9wCnKZgDaJEf+BdPDM4THzY6diD50SjnmzBWNhK
7pAsubqtrsR2sp/39lk/xQ2zjFGQesJGlm7jmRgXFd5PZ0t8UdpWPdBV+TPXqQI1A/oeIn7/EGAs
GwBcNCG6fdpNwvhxH7BYlE8PoDScdSVsD742Ds1u2K4XD7jCfoUxcYaMTvCGKYrd7ea5pAPk+nQG
zpYhCo/eQHhqFQUEN/m7QXpEJ0f8ZKUidglTje2l/zw6VpKBGRIYDuFksv9BK79ouesuugFvNKoC
a6iq5jll2jkuuke/21TJ40m6LRObjQ5crbhyMCulxgLQwsb1NCruN2wPpJjgWTDt2zvbvytM31OH
in4byFf/ni0CrdsZUFC/49z5U0Xg7lK9xVMhHZWdbz5v7Xoe6MS1nhIVpqEVR4ybnPhTf2eLA92c
ntZddbcU5ynxmmRvyYIC6tKWJTPOGIfJN6t7iy1g6vNBy+HRh7uCTkdEpQIcwYW8pwaqGLgKq4Qf
LrG1E/RR293CBfbqAmtcgnQStwLuuXmzFpiLvHohjainZ27PRLpXR9klFiAf+pesA0NKDpY9BOtA
G4wkM8c/ineJj5HaEdeyBLLyLWoFeHHN5GzcaTTlMUplRKS7LzJhqlk4oQpXs1xQrIybCdo33llB
gDaF+xuEL8ka56Tvcoa1RP13BtdunF8Ok8S91KAtUXA6PJ4pxIt6wC2CN8ymIK/stu97zFOSTUvT
TR0wE0+ixQ7UkfAX2peDGcJnA9Rf6A2JlcJEm1o9Kajq8xGzOC7C6csPBLpOT98TP9/hZZj6jLsr
s1WUcXGNri2CTz6RT09K3O6Y9HHJhfHIG0VadxoTX7kmbRwYOxKCwMD+TKRFTPVWWx8XR9oBYd5/
J9du7fQ83Y7uipFgmHrny9dDtws5LUxGII2BZawwNHovXavhQ4RbFVg1qcyoEgXPg18UM//8JNSt
ApwZ+I7rumtjTs0ZsvcpKSCME/w5uuX7h5bfNqF5LV6L5fk+kfecU+KzOPibOi5kO2SU4Jjra2dN
n/PT9iAkBLU+ctZwIGDcwycrOrN+74qle59gaEIXqNhgBsHpWfgrztLD8lLVTQSNU0YIqVWxyDP6
8BLCoVwyBqbDm2WbhrGzSzADiHBOXZD/Co6pLoTJsCHU4MPVUIbYzETCqg5Xaw3OuDs3/E8QkiW9
+gdaSI81zpHtbjLEV05v1TsAREIuImRRlUoNja6vq2LMH0ugS2w6yl2pBT/2CvrY+PDyPfE7kvcw
qoqt/u5ujQJ1qVeLnRBquex3eTELsXvIRXw6hjlpGs3J7pbXjzwhqjxmPh+HW26RILbHNt8lra5f
hx9WoeZhgRonm6x6wOdhZaHzfVKu4qeVm77227PQb9jtXsaVDYtRl8ALp+aGnBAhQ0002NLASfQU
TcErP2uKHGqynf4eTvfwERPxDn7OgRgHaOtkVO6fOhPv9CUnJwix39E2QixUIFcmTuTj5ecBOHAw
cV2wS/NVzkZmFNly98FIfgpXSsNLQIaLbLVjTFWQh95rb4dkRk3/hd3GUnZsO+3KloxpdFHS3xFC
Dc2HSnhTdFc0QpN+SbmvUtbT5+bAiZ0zsPEsR5go0FviEnqu0Kj7E7nbpzbNESLDl0JNJyyZtysS
Fck4vtSLvlwqCqiE7w2GQdeu831FoHxgPQsUErLI0MGzA7p8Nh+zqLsvXIFEwo0zuKMR9+uwfOts
uXyCjCrGlg9PoEpJ7rkowAlk7yCDX3XxpzsXn+m7fMYrDIATevWTL0OcVbsf7LpIQqq2/Qk164cu
SNZEH9GqASK4UDgNZGms70XrCNyNhxKypwmJMpgLow5q5OJL85dltJD99hYzHR1FLXrQp7xPLsps
cuV89TmiJWr1q1hU594Wr57M3Zff8TgJe3BXDM/H5NZGpR3B4hJZ3WNEHLCRQ3TN+6iaX+VuVLkm
x9796otEzACIhjU8DDvuVFkgBkiTIWBMhD3MEuDOnOJRfVL1IwuKKjICfpXYHMGDGSPdJEDj4pYb
SSE2EsbVybjv8iTKWwkgRPHsgHap4yeB1bzVTQeQQ5HUCMW0AGXdiSNLUOiSKb9CLbzAYi04xHVu
dFTmniVqMmmMg9U3u09OWgeyx57SgaZikYFgXfLLT/4ofjkuB9KzYoB47eM7WlvuLBmS6ZaoJnEG
Ob/p5liiWj+WBVxBEgY49pYMs9KaZeH4lrFiXEXJQAlomUybrAsnWoC31l7T2787vCvGhUeKRo9G
OU/QAAgG6sOE0sErAJAoHygOO0z2eWSa9grwRtSr4SwaE+4+HDl0p70TXaj6nYIZIoCO0WCD2op+
MjAg8jI9NREQCs+qqwf8Dn/7SXiXxHx63GzY6MgXZris2lL2LAoWHmrOfFUVAfslyT+Hm3SpOufg
CeqzAJOo/OOtCONEe/UQDvbpeCGlmLSj5BztgxNtNzLuONqTwQs7i3LnMY7fvET/5N5WdiIDVKH1
WWS9tRaHd27IXa9nXdI7r91ZdcFgPC7FR0dYoKJUZ7GTqxq0vbXiBKrVOrWRDXJaA3rKk7Wb91SZ
yPfGyhpHzIGOyulG5QwC9reH3VJs3wDidDeMeK73N1QdYFSjvqxpungZLNnZxCL0KN1X1b7fg0O/
/tyQ/KSiywcokxTwjCRpbBapiTnAFCSxfbMvMgpNT4xea4Upw4xogAWOj39ZLbDGD4j8hRP5cSRJ
EfojBP44BIpVEZbYMGZr2gBGfWcB1Of0QACOcEf2M0FPuTO5fE5ukD41Ugsq9SMOncnLTO6wqjP8
7NE7ZZoi8PD5WCMYLKh5R4bcyVdHap0nJpvmj2qPetSk0re2AzZjMNHS6hKnzYnR5n1RLGnQEebC
dxlzhtRXZ65X75CSKBJ/QR6dKidz0DBUDgVtn471/CEmYnF4XVFZNUqynG3TRuypJuCkeFGV3pzv
CjjnJCMJzlisbjHI5knkwp6RBm5DTxeqmN+3qC+e/VKa4PBWrZruUEoxSkNeGKMIv6YY0REv581J
coen9ozP7FaM3FSv7hw15r3WZqnYacw9sF1xOxwt331CpQpB8GRS6DnulkfYbkycMkyn6llv9JZQ
plaU0kkZj3vePS3RGYypsTzTvqmlaGVH0TJIj5tIoiSxIh4Qk29nQqHHdFJvgPcvJP1cjq2lYt/n
F0biGr9vrJf81N4IS7wX6zW8pdEVj0lFsgr1X+wfyEneG7FVB9C1yzrFveLab00O8pde1RhXp7Ze
xa4LKby3e7J/pPCo/N4BjLMGnT/bfiDuGFxnyyoApbQRQlC5oORJOQDxHjNXeyaEWqEBy283UbPI
ycu8Rt/7yyoInA/xJmiaCAatJV1x+vQlD+5j3BJxblZ7YH0A/VXpYZIO6F/hLfiV/LLwkCea9jbr
Q6owpUhwtn+M6d284meq/OBBjwzk8bvEagExRwZ/dDl7n0DNplfkDyiiS+GYQoc1VP3jBLT+fe6i
LF++SDW21ft4725KqNdWIqSvhTLdhz786r/5Xb1tGqqPdl9Tg6R54wuGyROrBpmi2X6Sd2cK6yjW
g2qO/UqpLECE3sXW6Ug3Og/MJSMRKfoYz/lcPkB9pHpKFKgG0tKDMMwYvxqdEydoyvOPnW6tw0lH
ScZ1VSTntIy7zliWuE/hYqIusifFoNfnXaoiZ4landfu2yDq79xoL3z3+eUJpMjFjMVu80HPpSIc
KiRUmImURBnUaNYqpVH8icieHMICCsWxySoIfPmSrrEmvjNZzpgU0ZidJLasjVZX4raTtvxAybPc
tRI8Xxu2TfilZjSsu+96cCxN7EiOAJjuCR/FLB0A4FkWUwUvEfkM3qwbxgOABUTY+NsEpCrtMphX
vDJivzA1cWo/NyjwMat5pL19U83IRR2yQG9gZOJYD12rg0VmH4SGV2H+iMc2eGM9BM3GL24swDl7
yRcbctC5O9qwq7CHfloqmcj40uh8v97z9eOi6jdmZqDljKQXQcTfGUqq79ODvUgByNIDmZcOMrPG
tY3b14/Mk0khxoT6VEJCadHwC/SV9VU1bK7pIdpx9VB8vi+hSpNou727LQ51YnIhKZrltMPpe3xE
VFWwXlWl/OTvl/M76iDPoETFXZkh53r92a7z6A7Rh+5D0lCq8UZFKYeoMocVNTjTdXi9EZpUD8gw
mr++E/vO937RgO1MKaoTKk+vDMxwLk8PBQ0qZWJ8VcDmdEE87VeT1k/xL5ZTOd8n+T3vRQxZtszz
FHUaws40EQ8N02O7b67c/YosdryDMCmRmAYf5iaJlV6x/1BnXn4FKmSKGFjUPUe64nHXppOG3l8j
P5Uy9zjsKQG5fiflCsr6Yaa6RLpc5sWV8+caNfvSts+x8WrCQk9wy7qg8ShRJudpwjd/kgGgw8TX
D3V2xsZiM8nVP2U7R7M3jIoO3QEnV7d9OYIZosk6A2Q7LjC7HBVpXYNbSLGGMOGZpR1HpyxT4RbX
SQVd9DEY5ddm95nw8+gdx1LNbuOn8NbX0u5Bd6Tg68gqZNfWbrEt7GlRpp+4DalWmWPIe0cgiyCM
UZlVAzsrVF4VX4Vr/IcaHOn6IoaN7aYZzb4y0ycp30osCSNJM+dBXa8IJgh8Xoihw75ZJI4pyNfg
9ASMcdXXvh0BqmpiJhptcIFZ2s2Qo0XFqBaXk9bKDVl2g243jBJ3Peh9yxiRrtUKL2VXcEcGDNJb
iwMnJ7g4IvdyKtGzPXT9O0hIxSzRyqJlH4+SgU3wur8d7qTg12Qe7PgiugI/ZvdLOlyUqzrPd06z
UuAtH1UaxHrEi50DnsQmyDQBCM3EwI4A+OCkW29lUM8rynQmexAkK09gGLndNTSckj712fNa80eO
K/NDPoUwX/GMArsFceM17ROhf9nP77d1NcFNI7q6YHpwt9NdmZDhWY30MbW4eTu9JIDPaUgPnmAA
lTo29W4fH0g24ipspuLDisvzkjBOm0to3S/XP7BTHnASBJ3HOHD/izSm3y+RKBj6T7Ncvx04JWTe
yrVE5JYrtwFI173grF34x1MeJoJrfv+9740BDlatgwQzA3FuQN5vBEQiAI6f/FWiGAPEkXl9/ld9
cm/0NssZmV7HW0f1+WSFtEezcBQeYDeSZOqXbRXS4gfM0Mp6X5AyAbNNm8nn6HAsE74m4kkhuPfX
4n922bcEf8NUGmYckJV1JfV9Wibk3cAyxRZoygnO5ustMCcvHUF6d8GbNkx6Wi7Y/iDF5BCRIA8N
OyPbmvodojN0NP9OxzItdDwpp63FLZg1FbNriBxpU2X23VJdLSC8xO+vZ32NRbFyYCfQ8I5qd6SB
ypYizznDNAVKWb7576o+qETSaKZeFvZ/wEcv72doq9sjLmZy1gxbBeTTUzU5P8Tq47XbtsXf4H8C
9XBFFkItfpteI2VIQvva12t3cZZXDPn5sMJYI5Jcgb+n98MV8fVnpIJbfvZd4lK4vm6IO1uamrgy
6r9ZbX/yh22+UbjifaUVJ2TqQzLX+q9CFdxViI9WZw0N7N+rQTBjMIiUqAbp2M0V4ZxutkQvw2NW
cDjDcFp7zLa+gqsUEollFTTNVGRRLZN/hCdHFEFf/RsBVU/L9YzT+NK17NXsNnLfFa+MRH81TCVa
Rg3Z1Lz5ZI6iusFsuFoDtYRL7hRC5CVUznEudukpIvX+10psZfDg7W/GijtUA+hbMe5jKbVED3VF
K06PeK/xubBRRMK66+OYmSBXW5clbH2Afrp3M8myZtkuPSe2QGUN5u1tOsMDPTE3FsIZWhlLnITQ
2GndkDaxZGWZzsK05YpG2U4Sepgj+DMXuQPGO1D1wDdaCjS2TNbztrb/DQxiWDWLAOQGYmEkUX4D
uqReGG/Brb2y2bBiIYlbiZ5P7YqdqrDEw6KALO9fPYNS0Q7LTD+Tqo6R+KE9320/No/iG1pUDsGL
5B9ABEHN8CvXIU4N24pCw9fbGVtqfYyvgzo4I/YpEOT7f61D/ULLBBghqmC5W5OVN9qbTeJNXOI5
08Va9edfOyRs4NEU9eH8ZgulxQL3QQl7WfCRPz6v91nhyBJX4DOcpmhwCFeR/UlOdn19YQ8aR81k
SyIqqALEByYzJpRj0PyAGd2zO8bAI1s9kzDJ2DevxIZlk7O0DyAiN/jrIYC5hJxncsB6HaAFMqL6
IwoTi/W1JXAoBr6LBhGlV4dUXg3Y2RxxGUkLAE2IV0JVcPGf/1tpp+O3E+viYC2g/VFP7KJPe7Jv
TW28ekiq9x0BBd6In3VUtUt09a8R+EqA2JmhX+IEpubnXdc0UCJ/8dzKlhpELwQ7yN9k6yZ3M26G
zXZFp4Pjs7adwWUQ/ooOBpJEpumpax6F4sblAXueoF88ZFm+0DwkkQ4rSrdvrJKUQiY/eUZ2pcrP
HhdM7xhEhcDnzSoF36L9XBz25Fvs0AVV3gUPXgHt6N90aXeRKEPjDGTzFL2UTiR6j7MiHr+CnyGE
cqFJHluUYHByc4zxOB7mFRRjjseKnV/IbuTNTgoQAxH6/ZnyPC2gqjDDCSAe8Krl55JU2EAooFR+
k3wNRQtJM9Err9+Pz6+cS8lc4aZjt5k9a5+4YtxJsvwFpgIqdHC8ASyVYzWwiqfcVwqmix1faewK
lSAy+PzHxkPlXIeoaLqZPDFp5ymVItpIynIaD9CLHfg7fBfDcx8yHVEqEi08PJ300WSQPOoo+waE
ShnQHvJiyn31GIW1AnfCg4aT4f5z4H7idY/VYZcFohDqITko/rEk6DznOev7azzFx/SyVkkn2Qc7
LwEyrENBLypZ4R1PBk0xXzsOH9ccmCiR2lLs6gqEugtu9Eb7vFqSHqFN62jdIC8Xvqxly7hLzQDE
mRKYWLmYWITzuCpYXckDJFHVD2A1PhWN2UwNattV8rVHCXZXxeh5vDuGwMB/aMO947aSi1Hcm/4/
VQIO0Zx7+JGDUVjRTkIxs/HpAOi8t79aBvhsAs3XadIUMP57pl1fOuIwJo4bHhstK0WDhyuc+wvH
t3N0wYnobkeo+X95lfC2/6iG5jiB9enmtQ55tan/F+dONc5PgoBcGXUqlIVDWLv/FV8TMgL/GjIA
SKpKQh2JUISAlCIL126eKrw6uqnjvL0Xtfcr1qOECgUq7mL8dHE4JxyGAKF1CeYeSuXhOfFI/YUu
OZTdXZRqbokkkNypNUfxAdASuCrvKEBD4rPJPEhaGKRYcZ/+/1xjyvhlLFy1TvTJsNhvUjpVyV+j
svKby16W7w5QVO+73gtc93XtflBtoa39nTiqsaMB3hp3nrgRjYwjkH6sjUHVBh3KrL7aQB5fO7kx
Wrg3fxDSxtlcqjH/Gb/zWjaaVBGCvN8Q7mPG3KChQ+gT17KHLnWj/XS9JVkHZoDRCEbJGeJWd0Aq
rUs+cfdzekV8mKtUjmPp2pS8A3iifyWQFn0364rCIHAPvDxcDIE83eq3+Kzmz6+l311uYNOn+Awp
oxYnq5VmQMsCL3aA61lLPrrU+o1QW2YKEGgWaViKCYKQ/NG1mYk8Wr0+1bopU5R4gWRbIE0fCxRq
pNpJd3mRhRviJ+WpfdZpp8pHajX31s1y/kNDDASuWfZEz0D/oEazWqkqNTpJJ43o7KNOnwgk9+0p
/OrVI8P7S4z+M8RZdI5QyygCAh/rb671sRv+lMLyys/OO/0Asd+UM0sELy4H9FYI/+aRa2UDkzJ/
cs5OYBlBiSbK8hNypgKvrYuLO9CQPvjromueHMXkt6yweQZ7y3A/oiFpqu4ys1R3bG1fS194Ey7D
9GV4SvSAaUhj5RTejzHAMOKCtF9x7ytg50WBfkGNv09JqinwrkxF+PaHwhou8x88iyb53ttksiMZ
/6ML9AarqtBf9AzKR3jSgnG0vD6RlVRfVe/eyWSzLDZFOGtWWzXpJ7e6Tw4UjN28UQpRKuc+Q1qt
KrURjCThitVvfk3K/nBvzajnAtwjqYPIRVDFcHYWv7QLJykvzWcIU4uonnHLLODaFQ+cJZMr/JAU
eniHABj9uDM69Hhwy095lKY96fCRYhRban9Hjw+JedVHfOuLv2LpL13b47F5oUxViGkTWG6w3Fv4
NOF03iN/D3Wx/ubo+5dR8TmsK/tGuAS8uzzFjG+yNbfdu1rwGJM4SH5oRnZHNhONOB4y17zibNhE
VI3qkcl9m0Hjc3+E+VXNU6yGC8vM8gxZ6T0jlv5GfCp9vQ7sTos5ghC3rxUHy2WhgKQ/10GY3xCa
vea9LJN9eqALyaqTI5ZdZdBsrjlrqeBpQU878i2wKM4hpA3K0BmxZpwW1utHRpPvjKzkCZS9NBXL
NVRa6sKQozAcMW4eDfLdJGxXsXKevK9U4ncw6SDigiQVVkQ9JufS7P4eCLU2KTOTK9iyHkUcu4TY
wuBjDs5RmXMTZcmDnvjdGUsgcYwk99A3G2t6zHb4wDOqDIYvJY3cZYyGjMthroPntR86TerDivPI
9zm1S4wWip6B3HAZdDB95fe7ZImMeF84TYZkGKeBCGCmtyUPxrjn+5Zn3uJn+lzdDzNBEqWRt1e+
tZKGYR+ZSsOAbVZuLcjMoq52OwOB4iNNJX1u2ppt7ROV2tt/+IVb4KZg6udihMV2xI+Gwjtl6oMS
aG/2AHZVDr4P9XgOfxAI4qFeJbxatejE1CRJMlydMM8MctZKHwbBnodHn2psFp/F2sKbySJ4P/Mc
kmpPulg8bK6OIGoKtUMuLLRDBIGc3P4tIvK05uorWILLGg5FFpTXAOtYOsqIDsixfY9MIbgDwlMl
Um2rjgCcbvyYibynzq9IdflS3AqQoK6/CyUuMLFRHjwEwfhkSWwLnmbN8PQn8YhC4T70rCj3HUIr
nurJGBMqMSRnr4O8jvOIQtmZkzVkc0+je1nOdpBTqHNlI8fAq6b8Y4dbIvtMJhnAN6rjNcbEQu8C
mMXiwQ2dYSpcSYSz953OOnWuiP8Ve3+1CcMeFQde2vfCqCEaqBj8d9pjjU1CNbURwWZ2/4rXW3Xt
8SRXXtAGZquZ62izbhrfT2PTj6mE8f1vbTS+dDKq4hAs+CBJdcFIc/QnUucqBv+v1YiXWmK5ZPrl
gazqZyZ+1VNHhYNFLwQX0jodj1pbmaMsMjZhZQ102E6PqSjjfzlXxcI+Qvs7eaF3NqCzALo1xUUY
Qw+V/iewTyTNWwz3e7EmgMSBfkABYj8W1RWtd7I+aReHp0mp1xeU4h1hYYIQgitKa7alPrcpv0P0
ukZ+Zl3/mB9XgysjnBO2uLF4SsUw3VL8g0Ir07H0pVEF2671NSJaLRbA/UQx21zonxW9iLEyVfCQ
mVZErgD8dpUiZhbus6OTf2soFymos4Xuvcq8HkIMwV+aaHRGKP3Tg48VpTsx9Mklg9V5zZEy7eD1
5DVLeSFo9WMZYUWEyzY+8ArzcWQUeu8jHQ0sXwNf1d+U/INC9woXwUzYvsLmlQwATVBEXzCW4vAw
Yz/RWc0cnKZIXgvF0nmctMTL/eC0O/Yy2vRdW17XOlh2AP8DPYNTttUWMSQnUPkLyRRwQ3AjYA/R
nWUsbM59KEAmdJO0Zf/i1/fh4nhpT1vKQPsdGjKsLmgs3zEozbki7rrG1HuyY/ohqb/uwwgUSOGD
Oy+4naLlrZ5Q+GQuJ4coeV2i9XFxT5NTPzzV9UVhAviGC2Gk62BMtzHoCoYjLOzKutxF8OkbncSA
DGhnKW1APCQUx0exAm0dGw382JvVFrZH8LSGAl+6pi4Rdx8lHmAk0uZAhjY/Ljw0q3H/FFpz09k7
drfU7haofmJGdHFhYzScgxzRJXm7XOm8y0WQc1BwCht9171CgLtaWPn3a87CxKKCBV6R5t0p8YUv
xgKxrcsRl3LFkX1Kah6s2CxRjfuRFuwgBq1OB8Z88GsLVMXP2XDmubGKKx+NRYGH1+eI+NweL3Xv
mntXuIrdLSLaW7WhJESzG27RzqU7v5RJWKotPqioxN1yvB+Y+V/IBe13tKEfzpl4/4Pwkck+pRjP
u3KpmYeTM5gtU+JmW2a1BVwKv/UOMv7VXi6obbIDrJFKJTZHxwkF+VCyvwVJvSWFCoQv6tJPjs8t
khXYhLfsbpMBx4uP2cagPhNEulXJ0X3x8I7xk0Hdtg14ixBNNHQL6PAjIlPtV8KDRkpUDags/Ysg
sW0rJCjucUm1Djyx2142P/NaBdCydbU3PiPxPSJWPPRT6OBKKt3fObFCyBS6km/XQ98VrGhDyJs8
XDO54YoPbWpYTNC05pzudHaNCNL/NjFO2V2BJoRQwLY6dBX96dxEuJvnRBOVamZb4NexgQYN/yyS
Fo+RNxts15v92lsg3xM+LZBAPmVy2MZUrzcmoxmohtiTXg+gHteI75exMnaAa1QkRa68T8BxVrDk
hXzb94Mc3DUXNhYsLMJ5o4osF1RPKd980MgjSN1P4Pn/3aWU1MlVeWbU8B/YZWxGT6Fch+ASTLmt
mSKx8byajY0LmL0aWGG/JWmuqFyL2NVp153+xME9xvfzU9nhutAVCJuJBsNxfV0tGOLWIVtrZKgz
RGPe0JM09Lm2oYMtVmIyHGdTy4RfvnfT7XigCNuIQdVomF7VEoeZBKXeJgXybHA0roW+erKsdUPh
y5Rxqa/EaNQIHiC7CjGwBxwrFybruZZW7N+dlej7w/NJ6zT3tIKVNBDwHc2Lytn2IIVioGyTdmaC
DCWxsNDTLiTOXZVw7BHtL2VRxA2XHGlGRedN7HXpFD5Mv4NzyT9IlDGoOFN0N46x+6xt0JwDe7NB
f80L+OmvLExzivhki10x9WxY3yBtXvFhnqkuM0nlJzySkzO4iG9Ch0xkGguIdioXCiJRmax8KvVE
eTktGpnAbtNuyL3y6BivPD0qK4UTNSqqacO99Km6eI4Dnx9HS7jDPGruegsp1Aju8pSXiRlsvzSK
UGRTcXrsJzTUFQ5WjSaubPEaHbfA0c7VcsISXBB70bcfHglpYUDnJQCLsj1PnOuKcDOG02zOFAqn
f5vgVRyd777F891NLTfiIeEqfnF2MwWW/XVNha/PCdn/ViVUpRUJzTWigY57ykW/jy8EDshbS58j
029FikUdZJHq2QWMUC5f7IJksMpP4CJm8ZBDwSHx8dEEz3yvsk9kmR9n+SJ5dVGOlwmlPgV3UoyP
q3PUCy2ElcslBaiVptA0L4XfIz/BpiWjzjQX/qZOFSUcI9wfk2bRtQ9NUDQXe904WafoBSjWz4iG
N0gZtLm6YqU0Hc5S03MrOfxA4xXxSgagEKdS1V/UOU/D+/S9d1wb+uo0isQW35b1osuIB/jXoIFX
uWUaD3zoA+ie+YJOccGq8xDUpEpuCJclYdFt0taef4W+ThwLH8nxfXtODcHYh4h3xt0OHXNSZb6f
RPD0m/NXEFFrbfXbJHBX0bU8bpQceLAQj54ZsOYHLnAp00ESgKqdLWCRktvuHR7SXM2AfHZY4Iwf
gR9Jdj9qAkvE/91kzwOuOXXbU36+e2vO9YvJQR8rGbFhYP21AJDKS8eyXbtYmNCzBQf714RTrljj
/jKz29ak0MpiT/+KZqrMctsr0RaRPFzYg3jLIHPsOxR5LDd7qKjjWYjBCM6m+5WPw892aP2eM0E9
eSfDpQupZM2aTJCzIrV3239i8m7jvsMD0dbutESxJM/eO2yKXsTnClyWpXlcx75FtDgwuqViwzSY
jRmAmboPbGCr4sSmdke6/5ECS2ZexVQ/JBEDqERojISluqb0voHjeKw2m4Pu/b56PNqD8QG/bbC9
jfTsVyR/mMGLBeT4dgxThtPlgbONzH+e19BIbuIlCRx2nnf8lfSDr7MsuOTurLf3988rqcvDz3A9
j935RpZ6T4NLus6YmegMDjpHS+/SGvhiONMMogfQrcRFYOOoiDzyX41ofGmA3sMU7sdeQ2AHUbPX
X5O5vPIAL1byjEf4qkkfGDQFjOBT6tkJt3gcITZssnx6zRUMZtoWAZCcMnQ0sN2epXs493bTQ/dM
0xNFUp/y+zduh+1EbEod+MLIC7a1T6SlHm5YfcOV3yWMJVfcszC6I9pZZd1IH/qQbPD6ZDL/1Ap/
C0/GjGiaAEpe0RNmD9xqCW5RDD4HrEC4dhpmBbpe3/XlzBHnZ+d77cOExf2glAb4QJuiLrutVfpg
xr2G/v4AUJilC+UudbBX9rghfKDO38neFU67CBQSd9+6FYhHF9Ozuqh1tG44/dpi1s0/fAj1vi8n
OpqeMTQnbuoPFs1q36hA1taZtsr+Z+URkGtpis657paU8UEGIjK9y6n6TXoLb1AYyeHZW2ulMfWC
haabk9SH51YyCzZ5739cZXjPK+4fiRJroxlmncqiCBGuZ2qdufBuuukdCNdLQKePlZEFB0lDxfCS
fSgTEB752EjE9SLB4PNXpWjpxRASOEz8s7i1DsBISHsAztn3w+1HiRmzgYpVfKRiXe+gmM66fjk9
5eSuGhOI55nkPpQYLet600BfmSsA5fLjEKdIgTkCptOd2PI/ZiflQK/V1ICNSWjHL8jUVPhKu0Td
LwDoiY62iuKLEhyPQMaU0RTJV5oUwu0OpPQznpQsN+rm79+buHdBLhQm3ZZrYT1G12B29Nt5A/Ta
dQo+EAzwAzwCsi1ZcKHMiSkUUlga6Xmz3/Mc6QvEp0stYd9MvOnESK/Hokoia4Zf3eDVueB1aQ5u
q/fGp/J+fnP5oUAsJOfCITh8RMe4ztiVmxILnSV8pei3Qz5gNKr1b1rA6lLELpHJDzC0E9/c3n0V
DBkwTpY6DQ92aOcwfAYg2MXNrLZOqrAXQ2CCoblbq1APSgiUKc0aR1dIZN+bHf8vkcYerg3OzHNr
oiFjwZJVY+fF08YP8uHmYjy8Z0Ex7fqe8BRD2nZ2K97v5ZMfHUA3gi40w77udLXXVHjysuLhK9MV
MQJrN3wcho7Xb+peydPOpdCE5pJIQhfBjIRjM3N9h9pII04VSJHOjoyVdfexYhTcMiytRPKqs4sr
NhwLtamOCF/6RipRTRlaJ8nrMqC2JkCMr9+pb84U03XcZZUpQ/CFj1P5XtBSBQQM3pXPwiNWrEHJ
DWv75SkXWFQob6OjTxC9IPRg2C/wSxGMl+GMI7MrA03Ltdo3dngH1jOj3oo6nJWi28pLwZcRkqvV
B28Tbq8WuEiaSWsFYbepLJMvJ5LWYVtssPHJa5iBm/JvINFlDrm254cpeNCGs6Z43qP0JcxbmdX0
oSkusGCiYBbAcojBoZEQb00tCSTPI8/TPQFYkK3LXc8/S87zXJBRSW/CgRIFM4QCjG40dd9VbIND
qwl0v88VEqrSgSgw7p2oqY4NKLKPxpSG9N4PhvqWiXtC0ZNu4L30vJhI4IeNdCPMsqGYNtyQsSyz
JfirWFmP5qjEyozt8kGvZiEoZaUN3J3f7xsIn2e3twWrVoJmfZFMDBsqlTklVEkqDDezYTzvTV+7
G65RlfsPnNkeBaSW5xy9Mg/0medzGnY9m8hSejAH+1XrE5O9Vswrb+WijUHCnrGw9Pj5wzT3exVh
R8vydcqZ89b2RG9SFYxR4oSQmYGv689mdjIgXNARkqjEM7Bdblt59kADi2Lj/obEaaq7bf/cvtt7
dZz26DuebOH3WO6Z5E0GOy6/ISMlQ0FK9T26ixSabBzgR8kCDJXf92LjZzpDbZwvIWNWAkSecZtE
lC5ys9COeTM3euW15FVtnULhcjABYS9003zLLzypIt5xdzqgvQHHVpswGyHdZxI7nP2x8QTRVgPa
NC34fsAxt7rT+amtlYph08Ep/J6h/yh92WlV2vCbgZpzpYJkxfYwRvHshyKzF2XCewaOYzkE2/bT
BXAqIzYdr+kwFpz+gaBA85CvG2880lfv3w1hugVK7p/8AoPj3BG9aVZgjv4niaqN+3RCiS7oWtEi
b01eRHdlA8+2p+BUtXWOsWWKLkpWlVvkbNOTsRkyUTml4NO07d+LO+2bRF6eYdkDYPXNvMMN7BUe
bxHNG4i104vuo8Tvi/abS6qNssCSPL+8LEhNVt4vGxK7ipvopRmScil8HgsmcblY3E8v1HC2+zf1
fcPHKeehjlBDDkWTIRM5ZNxhoQOqFi/jNTLDwZuSWIJnStPMUD3Aa+QXpJ0aITw851tuKXXUBfV4
aPbtLECnvZTqAg17Ltoub2q01mVJh1V/N2cuXHLUuxysdpbrdU1r/jb5nX6+zdZKuwXs58AU4w+2
Ov41xvwQv5xJ5ly8P/8txuvUUn5bIAZsE90wospCrhBU88c4elf2JMebEbQLQq2zbnitQ57GQyR6
5uH+1cdezAul8FfAC02pSIqjtwVmpJVQEmWt3P2aaEOi7jJ/b7W3QwlVbVH2TswS+Wnv6fiAeoSs
FqmN9RRIzd7vvEcMzfRYPa2Rf7xFOZrHhlaQqll0f5v0z47q8XMd4yVcOojHnIjkuZCcDNeO7sKg
+ScLDTFsZCBPXDcF+hpZpkffxDZl8YwUfOHlLgSUc7TLQPId3+RYfCb38xl20U9CqqO1+URmpi54
fdWW5wAv4tJcFKylWsfpjbRCvtuPw636U1wfVv8U4L9M7yeO2x2m/BhqFjbugphKuEidgCXv7eDz
Q3lHO8WJCQiUkI3bYK2ciTT/PSrjiYN/VmV06Y6l5nsmFaMysBRhuXcNcDZCpW1/lUOOfT8/HIGm
f32rC13Y14MLxlI627TOWD1UA/fXsOhthSBbEhsHX+UNhDKPicGXcItT4cqy0nHTCa6xbu1enoTg
t5LSOVObSWmYGzEjTHiltnBZxpXVQac9OPhKlOBmkgozhJARAYb8OJL6IIfPCwvriAmuzASCrx5f
oH78FvHXpe43m66WoQ8mJBPkKAiItHBBwLuoXU+hVwGroUXTvrFaN7M2P6RaYD5BMidsPQo4X7FU
RulpHmH52wJAgim/tCjihkXP/SGPWdDL1pfEbLhyyvzElhf7a4k+fTSbTSC+26klyoxCi3TufwcE
uEK1NYi86JtZW8C6VF/noU8uMV+YMUdCKV4GuQRZb5r+w1hmTnwtH5Tnfg5J5vj4Yj37eFpWIYxG
8ak+/IDd/f+03vlPOpbmqGirZRCZzc5jTN+qYS5xc/x2nqDyD4qy4z13Pr/6lWSvHIGblifYFZ/0
6iKSt6tGWix9PfTBkaABIAzaIUpwGpamSkCHA4Rnq395QD+FsF7JCMGMZrhUdaT/0Zaqkmjdlprt
I2PKDgHDYTt9wYdypNWDB1Rv88PMeef1D8aq/5ASuUV8enK39vxaub1l3nl4i8iAUppFrUztuYRR
O6tf/c7ePhN/1QbsFqJAlbKwSANrm4gmgoSvu6izvkgC1lPK3k1IUMIFE0P5pHpu3v0G8ENPoevP
BR/G8YA2tkcyGHUyhcyv876jV/Nlw4z7WWCqQXP87lrfZOAGN2lkNburEGDMwXYp1ioMoKT7fr87
69RZmzBRPLgQK12oRe9bGNHV7yVtg14DnhaWQH81BRMZYGc1Zq/6fd48p8m1UNX69VbYfd0EM8CG
QuY19opfJb/h5iKwZpmV7Ah5mGrPB+JFEnWyEpe97D1WGCSPCZRReXGVQAOabjGdcywqQUm6iIYI
PnP1LlSWQ9iK/VTVKeI6Xpo4fGuGZJH/dE9E8atji0OgbehUvdeapid3fR40TJPkOXarFJdWOzFv
eAJV8HEU1kTDmdK0LNK7yWwCH8RKKZYB/js1jRAfLKD9I4LrYm1/u7vWrClvEZCeXw55ZVqj+teO
m2BMjan+yW10Q16lqlyF00BJ2vSnPeyZHAVxZ1PVfNhjowZoHn/Ay9rkD408M+wmx7kDMRf/gQ21
lwoc5SqaG29g966Z6RTCmp9ZT6el1emhcjwj45VRBTA3l7ySqYfhx46wnokCHJCMhrS+nFEBxf/a
FnkREJofFmsx9XTaPugLUfpP8YJeivu86JtDf+ZvidzN6s7v5VnlXD/o1E1pl0T7y1XygZUXImk1
c6LYXj1RC+X87aNBSmQBBq7kHw9JNHIVcRfSO6iGbyicBFf2e4HAch7M+0oqIISrY7sm8jWrZ78/
WUkNfmdbnJ8igybPq2rElHpvhdJfmI3d4k+++zxyq6GWLuo0Inp9Lr/5MX6Sy5O3K00ff9c5/u45
tgFGVIvHSqeXrHOgq1Ixs4QKDDvul0eeo60OPpdTtBQhlIkm71fIkuOz6Rr9O8PB8ge9ho2oYnHw
qn8RevXR/uHZn/CaUnSGDm2pOoNodLM5aFyl1c8itmdngKdPyjDGJht5zZDukY6IVIlh8jpPaeks
uggE8IqNtdfrmU3hFlAnNOmnUh3FOf+o4hhFcoAn54cMiUVyO8Vfz4xfI48/fYE22bxmaP6A5ZPF
RrOMsO+vTTM+3lI425JbZCL+qFPj3eM0XsNSjwROt447zx6qwtDN1j3O0IIzUSWN0epWa+/NnPuZ
Y5P3G2heD3Bb/TaOcB92c5WCHA+6AxHz2OaSdPGbhcDDEG+kV0CpuwvHgJzX+yW0W5uWy2Xltkdp
h2Ap3xP6u3g0LFTXjERDv+r8p4o6+YlZByhuNAjjPaAxLIHZ+X2py+GTz1cNTOIhKBfP6fdkDfeE
tzhPieuTjGIoSBS9SijXDaUzFZXD1PmaJtZpwwoKKZA/R72x2XYtPf2bqO4yMBxo7LUaH/Kgs5N3
lF264tEdzW0gA+UOfm/+zyzNXttH7w4I0bdPL20gGs+7YADo6/pdHoF67xJTLfxrcXnwzAH9/ZB3
T6xo6450Z4o4Pq5Aih5m1NrjObzPQPbf0Yw8q1ll1vVccZDGrNgRuLBq3Xf4rVIjoaLI6dv3Zrae
wHSSBAop6zu2f99Ya7YR3nU2HsD4SKzeFZtXOMxYGt0eXkNsTHdYHwJi9TtHOB8nh9JS9wWzFzyj
RvpAvLpS4RPdMn6wx88uVd68RjYfIigE+c7O+wR/V5+GWEpmlpibP4t5n3TxkGVYxXusqniXUSx7
IlVSPCEOhaIx4aambd9GGlY05bTt0ysaW+G+ouUxhC6wgjosqehSum9vf5ySDqiDgk5Z1xbaYNnm
Pt4IWIdARznf+XdouBklh5wUOEBgQ9ptYY8SPk1FMYkk7kJLh9KaShVEoKLQHV+KawtE3gWI4bzj
1Dav66qUVjsRu2Z8bHZvtoux3mmdAC2eMWnOSYuPIF0XXD8JATDyVVGzINp0/AMX8INQe53gs/vy
Lk+cD0zO2T85sF2wFNi0AjzGywZsOOKk0dDpJTwmbQaTflXWm7Urr8dUg5KLbcqCm16HjLhpEnk3
ZrO8d5cSAyJ86L7jOxhvK9i5+rLyfpRBZiInPDrWrGpKWI2t9jBeOTOHI3Hxfhn2chPWB8p8faJ6
H4ErusJ721uXdhSnQf5hjijTh0w1W2jLGGEzxEu9w0C1CfWa2RD6a7odin8cD5BT6p4nUdDxc/Uo
4IMCUfzbvpfoW1FxLWysEwJiWhZ2tsLsLsMcIL21Cva2TmWUkGuUHbUCRtCFW10cKXfdj1HzT4+d
lCI2IevTdy6/DeRMJ6uNC8kHUjGiFRimOOxS3U7onB2tWN5XEZR3OJ92/LZpX4ZbcXRH8nA0JCFw
zLc8Sq2DsJqtQjtOEWMEdP96CrvL2sELf2SyoBJzZCj18LCFmztNMlqzvZiqlKiiytbBboUInB4f
/UtuchXhdPcTAL+iienFFqV7yDfo1XT7a84XOb1Rpu7iowwA7kSsVxvT65k/LOVkGp6dx0/y/Qbd
ir6kuTrc3egfEUuFZcfyung8bj2GieZkE5hOgj6yuCirRbRyQWANY515xjfTGPdwPBrt7HgeP31O
BDIPkaqoj1V2awKjyjAZfy0aFgLeF9+MsE593p4xw//rNEoTOijV/oZvYfotAaxkODMOYNOIcddd
C/8KOjprrhXBcn+BpXmIX3IRmoVthJwQLxbfQGwjIxLuFzlK6TCOctgRUZPSEWBoeNelWeYhnxDD
VjHXTgm7HW6N2aK6wedflTphyw4CAPKcBbt8/sESLj21Nfkb+G7r8aXjO3XWhzfUkfcjZF5dzFNO
pROENLvVKx/okSLBtskqLRJLGGxotWkuCPV5kAuxi/fLhuTcZdY8iwVmrAuptg7QP+46HZKp5Ghs
lVEzeGrFjWkTSUOb0bxbGQ3y6Yasd5ts4G8lxXtiq/HjzuvbkGOQ0+zd8w1qKhs/N43jAlkHpVKg
RJglE+GD/1kpBzcIFkMa5azOIblaq9M8nTuKx7daAoYDc4UN+Evqm6WgvjkJRSdDC+xJtvUjBeNn
xPZ1yjfkdbIRIAR++F8UictL3hVvP1EAN2oJv7pY2qqhZd8Xi1wIa8nHTeYmdy49MbPt9BbsWFB0
mDRj1swLgbETTcT79T2kBWy/YHv2Jb5DyzNqekuVph9xb7oNie+98FjBDQZnWnProcxE5EG/WR0K
SlMuVti56fkPHxJUj/w5JIXg/08f/x0KGNi6sYf8XfKN7VqqMaEZ4qIh/w1xUk3vyOonEodnfQMQ
XFC5Cak3qN4KjxE12wNb7nPNmD6YcxVKFqIo5hq2bZ0piYSAEqdxXdDqWI3HATrjs+lp019P9I2V
8wNY0yEAd3Cp9/agTTZsNPEuA3nGz7U8Kd6aaiBqJedddXFKzVwhHq3E6VODNXkisZmz3Cbqn/T+
zm/I4gURtP1n5Eg4LAlFLtFHs6WUw3WrhEExlcDLHp+z0nVmO2DoYrtIbHEwBHbSgkZLPNj+prcf
9KxjPP1m7+cHH5hMPqVGvlwrgfWXPE9lVSU4oq4pp/0uwhojxhNKiuQVo2kP19ggmXaDqaN3Qn66
4oqV2Tf/YIeX+9OYjlqc+wddkAzvHTDBkNKVQSP8u6LzkMoCR/TADiEhIv1Od6FFjvNmDLR/hUE6
Kttw0WQw5fxuxvyfIIL95Zu6XEaMJhDhbCIqmTwJv+yA7sKp2l+dJaOHr9nSQv0RDpgFHRW9SBtX
oyCTne5Km7bzEm8OQB7LqaFb3dlLUmViMs/TT2ACDXqU2dvTAXcP7mqaOuAbIFI5ZYTqwV7m2Xjt
BZol9TcntK7oWAUsY/xRmLd9lQXSFc9/sRzKR+q4Ayh2h4hZZlK9mMC7YmZOb+V96Z7lMsKTcSzT
GgrsZzQecvVZrJJUVgcFq42zntjuegYx0oR4a3v4DFtG/xKwvzhvU5DiytpV1mPi/jIRL6bNGXej
Qno4OznMVmI1LvpNUV3x4cIJPD+fOq6duUwDOQ3/UaUese57AmpH80+hYnr/DGWxY5CZPIqrZ5Hl
z3XwswssYLY7rFNTKumjZ+OXTRgLcxfKs3KEXD41f79FEiND18M3+082ClNe97gbpuAybKtomoL6
KfrZ7jizKT2xAWcXBZoJHdczHwGUQIvVB7zaQH/EMy5hVfElIx7ag5Mqxr6EZeQmToSpJgMf6yLd
PqZCWNVPhSg4/3fWhVwL5UVc9r0jOopxUqpZ1DUTDLuCTXaWwlG3C8pGF8hoiqCXhWnOiELzc3sF
SQqb5IQS6hV4duyDSWdmKPYhvCG7IUM4XjSvkRTOh1rHmfoVaT0gQq/DMEOCZ97oqDlzAxng1qeg
nSeEyKLMk0YGdOJqcYJ2IhrhoADxEmh09Yz5mleHddTAQ7eSwO4vaXv2mUZa9Hoh1DLymZ/8boby
gxbrTdZm2ut7AoZAgssTmuAnXv3fVfTMoI4pMe3al153W0LLZa1txTKZqHExolCF5m5KMxuhJciI
yS87Ics42GNNgr9hyYk/NxrDrSVSYOwebaxq9sEep2fFjilYyfvgro8m8f0ivkTq0+9XLPb2vSgj
FIHJqvkyuCNwJvaRebOos9qEEy93BjkluhL8W8zXLOqFp9PzX8+D2mKVZKGs36/R3Uc8AdM/nTvN
GZ4Jl7QfOqLM5gQWCnYWT+2O18FTmAKqhTSwLK3zorWvusmuGxR852OaO5ilzYgQqa6JcAu6jlyY
aolbb2cqU28SaPr0BqTMKAjPOM9vHQ7tycVBSP0xL2J+4q7JQcDwcmrvFtm8/aT5PrbX5PkSEglq
7RqZquq2Kmyks7qNRAM2K+a/Ts+EGI/fs158zBAg3omOL5Dr5Ij/myyBfqExpAakQIVSp2t2LacE
xt250KUhPOk0LsGjoR0gjejnWthKntqSKeWsLFC8uIB5rNl5O78EbzG2Su60p3Yq/pQ2GEfz0HbF
7XzH0dPKLJn3yJqwru8LiXNjyVARonIomMhlXgcuuAL+egAcjTNrr75a1M7/uIy28bKE0nS93k1c
zGy36hPRcd2ZtaoM0ZLRkaMiTF0J/SHel6g4E2he3hLkd1qB/g7nhQuN2fn2SpU7K238qsFkmZwK
HlWF7RdrwFofTPBQa3NTfqo2R+1i8kWIsyHSGc33RehMvYRviPgT2DkZBDSHPZh76CjtIHb3H7zF
g+Tm0Om17PK0miuWjKyrEZbK9lDiI8CL96SrJYDbbTikdxwrRH6tCXqy0ie8zTrknNMRXgI5SjgX
jxSS0pgxniGedu+wHxT8hRyavGGYNMGTpHTXa8e0yn3vp1nHANtYOOEq1oib/cIhBJ6fZrL/LbxP
/RwZ1eJ1bR/Bw5EKyDDIjBYfzfcKD94gTwVMB4jWcUvK+LD6ZcR7BGeQORgS0Q3jIgpaWfypzAyY
wAahoy2DHpwbtdl1L0jjodbVxZRt1qvlf1yAHyk8dPzon5KsbAvXXG7HkaY1AxcHqNmNkV72tEig
MkUMIYSUTFnK7RCvbUaCPcxNWzWyhswLRnCCFNdmfdsaHQqmpyenrfwakd0p+scuW3qoZ8e6ojMt
eBFEbL22uvi3YzMEdj71a08aR8wdASEgPsHBYKlBgpQ7IMXxqDhp47iWfFv91AgGRLIosGWmCDvk
Q3NQ/yx/0Rbx17uU2/2Ci3BnggwYC7nGfzU3AizW7+tCX6EKVZE6H7JNLRJufFBtUN3vCeP45zVK
E2yrEYNx90fCYnO4s04tbgQfcJlofrkG7Ty4oPKs1Hg1nBJcUKuTqeg2bxgV/UpVjjATYZvCRGbG
6C8GcLByGQWy67dMT/2IERjhAZ0P7D1prGASwFFyiHpn2KoqeVl+ewNFW9O2OVam/vowIT/9tppX
OjcznGl1o2QHVrKihDagzsF7g0AlqgGDO65weAgFFEi8ITj6mvDbk4/YNLg1Qdh5SnqqiMMv/y30
3i84JApmmN3S59rd7LMyil9wTvhWhRa34QiFbqFjo6iBuOJIk/w2FvvEZWvZyKiX4KnndksTx2/H
sAJxCNE8tar9nLWYcib5e1OAeRvroUj4g+v1OxfhbCd3e3E1xUnX9GJxIXhEDt/jjeDw7LHBmPzb
XbcUshb3X6To5YuOT+erRHnY18xWj++UhJ1kKCWRkUGmurrR8tY4wtNO+yX0D+PFIj6n7soldYIv
/ErGJEmiRXLnsr7+02dfDUosPtHc6zfbb8sxMerVYmX0JIcOsXzOJDRfv6nfegQr7ds3XdQ6Oobu
jCojyGAlICI9bbhrnRbBSbr5BmzkCRICgGZ/0cWlph7eWxaR2PPOdnQTLluYTwFicT6AGGXjKz5j
MrCOBgWqB46CA4ITFDFzeHNuwiNzXiyF9qB/t1gVAuRoM79fwNxPxWoxRP6D2NmdFk4eYb26eU/J
NS8jCcARr73m+lpxeGRgwFV4psWfRK9WDWR7oB/Xm+2IlfLIgPqAaPVs7l0L+kIbdv2oZ/ri/MbK
8BYO+8+n6qQMtkQNPGF9JboQV1CaInp/+La/fescA8PhoWFsVoNRpp0/ebNIIVJYOKRbovbJ3P4g
c7dcWjr18RF0UIIcg9/GErcZ8LW7R2theyvtoUibg+GcU6SoRkcf5Ngm5g3i1KWf5lpHARk1b6wG
s02uvjJ1kYA9oJBkA8zmfNAjiZPoKN4DKTKpoSfVqzVr+a8+db0rHr1SkJ6aafJT5Iw5/i0p4EMN
DVmheefqDB7pr7yQRHH7t9A82saZwaI1EK0jvlF+XVExx1N39b//HuwLbQs6GSaCQ+25p/F/DX3u
6jQOQnnt8oyT1/57ukbQJvkcHqNs/PHk7PlZmGOp2MaK70x1S5qydsB132CEb4ZEt7arkpkeqVEI
f4kWS2sIQglukWe8HrNnRvBgK7pN5OJWPbm0dq/b5tUjXTU/4EZIebdeFxnQJInn+7oYB/E31CYE
S9lrxi8Mpl+blE6l+R6sAr/+wBHFCto0NsIYQd/2J8k8M9A8t9PerNgoELElBB98losiD5iihDnv
yObX/zizagyWq+8hjU4s3W6tNn/mrlRJNO0O/WuUNWsV1kBem04bM9P8wtxeU283j8kiI0GcbmYq
jW19dVcUzicedyImjjeVWNvQWtfkEDuROIKzTeTiCDme1OKNVWHIGJ4ZCpnqi5SCY7M6CMv+8KAB
NM3PMrqHEitNMPF77tnAZ8u6wxBLnN6VeB3y6P9I+slOjvc6ohvv/u2RJnkR7hd1ojujGzz760X2
Azk/kA+aGOO9b1DcS2vSChK8sNPscRFw/vbiHhOK2CXggXrmoQijkl28/V4lUe/tCuUtyLyl4UWJ
AVYQ3YLjHiI0lBrTnt05fKZ7DLpFKTz+W2vBIOjx7QNRIOWspTla1dLz3divJc4P52k053g+Sgkz
AYYcCpYbpHqP1WPXoaTlaDfLvxBWLgCCbeW5omayoCFw4Ob+y1YoPSDLMBNHwcm3K6mQ1dx1U8Nk
ew8DI5slOdJL4lq3T5hvt5heRl6Mx9Jmv+sFLv14+g86sanb83v7m+9rfhzKRN52Sj0M58W5AESZ
dXJDZ5LMUfR+eDKQRlOHolWCh+VL4z7vzv3lRWEyT7YOegAbgW6sWaxpnssGJXAczZnl61hWByrH
vDGMKRCMg5vfZAlvUQV9I71ZfbWzgBX84RtaJfjtuqlvHKPnjKEekbfc37J3Ge0c3GjDFeDhegJO
7bXs7Q8Z3w4IHAnt+1HzGdZHgMF8lCsJ+PyLE86y8MWAyAAnjTQdfJ8axFxMu+yJ6nsxBJrZf8wU
6lsuPZvNnEleWql4/y8iXKYSqAQoEj0Vh6tHnXgMbJ5QkOcFU7uYlFs+GSlfgU8799l4jBPTJ9EP
vuzx2hoCUjE3P3uDUovlcHtk6R5M9Uf3aMS6OKBs+If+qD7UCwCtPE1mqLwpVDYwmatbHeO6qNU6
oXd/+CgbR9kjYAdbtXSAP7GYI9/luhur38xAq+Qzf9yoKRtBYmfDQRF2jZ76KgPnYy/1lsBUF/Ke
IaKu6+LsJ/UkAkCmIbkBx2FrOJyi4rRla2txJyvW8TAF7uz8cEWI4O3Go3Iw2zlyyp46c+NLm1gQ
7enuYY5ui2m1be/fjwHLIE2kWbeNNTXvqXTEenB1+6o2Nkn8Z9tLajwOIN6Ra4cgKDgUowJjAMbm
hNEb3bXWP2a2ExDdPqcT3t9Sl7RzKe1r6RMGYxkR4IOL6Ox90JxbZu5BrnsqySDpu4B6Yq2rXFZK
eG5Ld0pT4vMExGjk4KLeQ9OwwC4WkuTbiZ1ZHFTc0yo6nPfGeNrsISJTsBsjJZByzBfiEwCBkLbD
VDILg+IfimCxgU9yLBW1nMKKMns/pgL34l3oaYfghNTdCTm2vNVsFB5uucG+9+AVl1IqRfcuXcqV
aSdetFtrKm+EPRFg4oHEieKX8UyYyuh1wNtNyPEJ0vzMpBrF5cYcRkhacwpsSs+qRbRD/dh/QiCr
WrqNQvsmWg5f320klgjzage+SZRJehgSOVra6GuwgheMOk1DiKHzRPOlsLPNKqDS05eA52ESXVtg
yoNUw3vV24NXMQxKkGZw2Q9/V7QPyCOGuzhc9++oWSLAPrtl6jej/yidpRISx/kspLUWq3G3wN7L
5QvQMcMzRGayWVwTVjVpJIDSS8rsSoESbuWkY5aHrCKjvimMCXL1bvtJlf+bRahARANMn4T903J0
KD2G9C6ijggm4PsjpA0I/enPdhFVsOsmoUqSYuAWurLb/kMzuvhQQUFkkttAzYRO3tSUDa+drjhn
tu79QGAYj55ILVWpE64RLBnQPgbPIVWDk7SAuusk1KevhbFNj+IwIAB+yHjS2cO9iPGLpkERnyqf
d61jSoi7p+AoNOJUccS7ZMQUHkFVoh5+QZNtR9rooj7FE72jHK06PwprhWFypATyqeBkppbANzzz
4RQqlw2XthXcgColjmUmctjyAEvEdb3Rlq++xVuCUjtCMnk1kUUW+uzOM6cLPR492AttqYRq2Z3a
IDBe/xvc4ZQIeHSju4wHoowudKIfbTqCU+Rec2L38/49rjKPes4gUcMJ4Y4fGRXK88i3FnYVX7aC
QxU9aOAIcsadwttjDr3cOkhwq62Wv2bL8AUgBVMCBE+hyW7JxxB8Df0Q8vsY7dE2DryL+4oFMdqo
i3SVHCm5i7gSyRG0B4An/yjO4BTkN5+j79ROsB4PuyQgw7h5B00hWnT4fT34d0CvWL0w4UVkzRDd
w7XyxjTXnNe6+RD94tuIsKiHN+rgzDI22kNEpPhbNxDEGxKv1KXYLLS/eBJHE6fBet/F4v8BiuLD
iBOf55IrLHLWEdfVa1kx87MB78Rs4Df3hxj9SHI0NwCNPbyCqDLSEMTGXZ55uvY8HcdXJFBkfzQW
12Vtzki+gh+UgvnKGz8dzt2z7taLkNGC/GXrg5puJr5FC2JHGYDyDQBtROo/peQC79xRHk572TeG
ClEAsiZdPnCdu6uaecVybn2KzUgWor8J6ZArjkGpWIqPEgUyL+E0yAVJQ8n7nqLwWXd3B3N3zTml
zmuN6JUknK1/h1/0eT+BxlEytJd0NLC1eMMkWW5Fj690X3o5FLi0vS+C2Q+optm1F+Q6Atl04Ns1
FySe7Z9d+raJWyRn1X1Zi9WZHdNfcSmxrv7VCR10jty9/vH31fBoCu77e9dX/X5D+waLI3XnGiQ5
mm4wQHMC4bYwMdM1DKS4Oe25IEsFTkzYJTWpF6yQzDUD5Z048malZrOjQ3ZwrM83b0jrvuFEpUEK
cXW2OlRR48Lk96lqAzeCNuspmhBnQlvxhtfN4wpZcfMjNYgyGeF5rBnVFHh1xBGDDh6gjgXAv7y0
yB3VxvJdAbRQBXwyGGcfwx75z0jJdKcnZqcvEkmgYx0PKq/vt/rkbW+exdfhzT2jnzuzWTKivRG9
22v/StEvWARPv8Hic2rsTy9aZwrIkU9eueVaeYUhrMT7a22WC4VUJBVd+mNExLXhiY+9eGgoAr9H
yQih900D1riKExcQsRfqrNX1Dh6yA+0Nphb3fRHWv0MWRWGiUADu4mxcIdStMxeeel0YDHqTBxPd
LOXvKl2L9+jf3TdiIHNyt6bvJpaMJhtqS97flujCo+8W0EZcSPNAeoBBwWtd59Mjl7OH4yxjJjkX
a7DHIxWRmJS5k4oc3KM//vxgbpEzXFFEwpFrXkh7fklO/0Nr3Ng5g53ha22y2xN2EGxihd3hjey5
yqzVgtrrQP1QzkzcU0l/3W+emwqH2TH6PfNS5bLBKwU85PZKDhri2StY+BqJ6z3ouVMVuDCMHDYK
brxbv+d8luspzyzr4kUlVI+O+Isas31bRpVjFa28V0FOjRSynJSXhTnJii9pOzGRPKdwnivEOYRi
+Bm+AbxOxLm3QdU5ERjVEykzm7kqC6xRcLY7fHNSCLE8zxIh+8v4GYQgKd7Tx6vYiH8gbh52vzFB
DnihMWw+XAZGQGr0Sc8TqToZXP/Jj1g/6XlM3rr2xQf9+aTmZfcyX1BnRWlf3M1yMhuKzBjFDIUi
cBYnrEaJAD/hLJK0NIAmfRSmbUB7Ij/rOStafecpsUti0u59tw+9qIDFu42PTwqI1ckKnQrllLG2
Hkzt4Pp1QNXX2uONqil2SVU9rh7mr8B4EzzJ8Mxzpskg98gm5xMWpp1VWUDv9G3JVy/y6jV1nY0P
X7c/Bjd25KVsXb5yEobNEry8PN4NvGhv1vY3GIbQYThPu6guOVohSUQNYKn0ZYTteu2FsetiSkzW
Iqz4bfXcFdsznb4bqp+UYAZNhB83GkqqEzNtPYXZT/ygyEeFZd4cN8BJ95wxseBlI9jaRDtIe6Qm
SKiXUgYTVvTPKwNsvezSAaJUDkZFxej1RQghF5XA8tYI+CIILOov5dVq1oyEkK/Ur5xVyhKQbYFP
ncyMxRgWmHqySHlG0/3hGUwbeaHOJcnMfBI/1+CGpFZy5ODhiruzJNtvHxPs+FstDrKJ3lFHVNO4
qtn30S9x10/r+7z7dEonybgbMQBq4rCLc7i0gM8y5oshLwebCM822GYKaLya6CZ6bsZXKTGIZ2vn
oNYjE2LNfYhl9Hvf+LQOvnsiBcKz+KpM2Ce5r3CuszLSMLbSTNsmV9Z+3ooXoOeEvlEN0HUTovhH
Tyqwsy/hrV/HJEKIOk6jxU1mCI2deoAdtSPXPE9kZZrQGchndE8S+8QhLICY4htBiS+ffdjZbswI
a71IO3zQPlvJ94exMo+QJ1kDsJA6fShW11iBPziO/Fhe4AKAOeruJ7xqESCqsytzv80rxyxP564+
4MYo5vClbbiwcw727OYYRJ3JgtgZRrB5shYlYh7AyI4qS1WJasDjYOuMwBT0cBxRpg26pb+i2OV1
DqYSh6DvgE3IrbiraM2xqjOXvasOJEHTiF61eocfvPkEIGmdrvLOVxyc90dunAbREuuX8gbRdFps
AzZw8ntvXawCDCDsHwJ59hLuoDGDv+mQi2sI3x37RUr75ktZHdF6sxxh4iC0wN9GhQ/yt5ewzJvT
8jkagXdPLu3FwCAVyWFoutZs0jClm2OcDRwCWPzSMtTcD50+W+xD2mykPeOdZr4GHSdtqD8fTO+v
jKUXzl72029vxEU8fciQobN0qZQL2QPleSpudYsdh8lPJQIAjGCZXRzYhVusjq0MT542gXHo8iqp
8zcwusGIJAP85PLnb1cDEK4B23md5LQQHFHHtP17XS8DDsHwS/Y3DOW+gcfI/Xxd/e9NoCtCGDrK
4CBR/p36XLO3mb5F4deVDbb50EedNKHHIFlazT2ZVGlPrC4xIx+BnU4hPkKQgOS7bNhVNMsDUZlc
x+QVLxp8/sESZNRKlUn1Zx1LAVLVU89j0NlezWPJAWbLscODvqCwdeioaI5/KMg6fS9VCzb27OIc
HPp5lwaRyHutR4YANqVbEoxmLuHJj+q2ddJt2/myl/OKmFhySvUQR2cA0qwmEgnCLn4ph8/GFBBl
5zQH5ia76qhBjPFpgGxia9jzb8aVyPCoE4wxJhnFf9UAxlZfdiQ9ivBcUgcrjxRJtDalzgSCJ9wh
w4co/RDaGjDYniga8JN6JoE2NFC0mnzn5UrkpwIEC6sgrt4vhlHN6PkqqhNEXJxwqne+AP9fYuzC
vjrpZ+2G6hbX0b6u0+r27SdexNoeptEPd4f110yKYCmn6QqFJ9+7sVrudLUgGLKBsfXWlc0kbCRV
dT1FuJyzIEV56sCy41DY/Jdb39J3oUs7oPb3ZRd649MRRrERvthL8h9kI+LAOVPYsYUf6h+dHu/f
a3GxrIvbeTDvu+VvIjVZCRlSOwGlWUFpS1fr2XNV3jMCVq+76lHlk+Er5a4WXunmbdfhN8Tt+WxO
LouV3yQh6z+MRTSFx7hQFOwHPb6PHCrGqJNSNUhfXqJcZ1Izkv0XXOIapXVBwkE8BOoH2yfZmZAP
IG7YemxKR7iCl8agdSrb1Efcy5dx9FX3fwkcIVrEyhhISMQtsPqpiDE0iwCFbn990LiX+YUhllHS
RC0bRCkzTlBm9MHA+J7qy9FnXyz3jGsegPHvj8uDdLCZSw8EupnecUYf5YuJ9gA4+O26XsSUpP0z
9BQMZZ/nGBJoMMz22egyiBMAtvubImq5IrwjpmqbgWdofyRj2G6nEkJlVtalH/yT5tAJ3/t8NaXM
lEioOjc1A3KYEcfFngKoxi+WsFWUvGlig78IIWVsnbvvJwW8Oz5r0lpBsCNcBnw+Ya+LwFa/GXPZ
Y0Df5rAm3EhCM1WE3EO0tbFJmK5X2utb6zv9hZXYNKKqB5jfXjuhMk7HpcgL2xCNJLvwoLt3Pqqc
/QrLXHqN3ZEbQth1agMlzof33vpofEy5nViVOkesGWJn9DQK0Nvg0ud89Zb1+vMnAvPCF5FRibyG
iQ+sTsHdbEjFHVI4nWNI+OoqRPhHLjcah8jpTVE17/WNvWJt0cQjS6aU0i4aL4isZ9zo0/GlK7MZ
ycHmR8Yp+1nUgAA2KTLZYoodqjizfzzKOaFtZZakHoOgzZEBkbbUMiJGf0NnDgOOdFkY3Ra7J25V
4f4LNzoeonvQOm9pBXDH56r3rudXaQMb+H7fp2msIRNtgLHI+iusIKmnnkQ37prhpJWIYOu6SxUJ
JFJ4yBRytsm/elRAlBe8uUqzK+O8V7cS+pLmx7ZPcGzD1N8tAEorbDw/iccfwD/xh1day8d6aEb4
b3t6P14sWtvhz1h/Ui+IpbyEDJ3+IVxXS8Ixypu1S7xZhC7K9hdOU01RE/oolbtM3PEBOwNgo+4L
6FcLw7CC3lQNGhyHnI0ZSWeiZ9vHpeBntgw0Xg7McwO1IiSbIjg25yW1dtzR6U0oqr5BwzIXcDFx
EfXjW8NX+mX+Pj/LEV2QiXyKmmGR1c7rh0LXGQjdkVjtAC/H+ZHPBa4VBIaZD+KFPkeQ5EatuO6M
meAnZysSYMtvKidFH7wilVEg1rhW8QMafM7gl9Y6ILs2bfAAniivPZ/80QxJJkr6N6AzGru/LzsO
8bLWxeCreQPvIGmrEvkY73Y8mntz65mzswj6odUNsrCMcGBtm/7JjkPFIpbvFA5YuTcoCLSuxibv
/+vxVujOlnz5W0o4432T3tlaCDpHuWAwT6i5Z2fK37TOen5VIijvOdVJ3+qsOJtNPjAv49qkZolc
6k4DFSwA7OdCW1HwlaW8LSLvBoQS0GbcRpV45OsVnJc66W+Cg+IZhgm2k8J5qIwNqkwYXcwYORVd
QdsGReasBwE+7TKAv2qQRPpz+pL4X8IW2N2RCA085IzDufduDuccgRE9pDEfmLlkYo/fIZz6ZZZ8
YvujpFRCYFabk/HJYn9PJNolkpRbC4OTBckWfcoJAmFev4NvLqlOHKxBiYQb7ZWKbDs4zNyzcnLV
H9bQtDL4BLwHMkTsB+CSyY1mSjs3ykkzr48BuCIMiQ3/vBrsX9ZrDd+bp8s1hP58b+zPuRR8MOR9
GkktE5K/1O+CqYI8lTZxu4A66Ysv0+ClyN28MbMv7C9334PPwwwMdputn1lu2uUoEHPDm41V1hP6
hWpkQW1C1jjHO4Jg7fJELPuro0f16LRoayJYFawuCKJjjdxSQ2QohAY7H4sHHrS6bIpFgGva4hvT
i8mexejw8X4Ib5WcyB1NS+vSO6wmqUEfm+la6oGegnDfBl/ArlBrvjm/fn70YjbRbxwBkh/zY58w
bdlkeh6FpBLqptPNu16VwKvhifWKXeHlmwNStyUR/2MPdp6jVuxCC2WD9UzJkD07asKA0YkrE63v
PZ/qOMLbVD1zdBD38auA0iWU42H9Er8VuP+mfRU1F7u1JRUSIgvMCtDcbC8t+557yhcVcll9C4AU
c9nmC+5n+ECzJ1ZpUOC7mOqvC4UQ2Lfk92WxHDxNe7a6HmbZe7MZM93F0EZppbpsWGeYbNs+cpU+
MMC2rcjuoAAS3EwiGvsfIIUlHY5ogmBct5gIPcGlYw2NTmzItF12r6yUU9rCv+QGAXlKf3pvSn9S
N7/zvstfUKhuFiVrfMzReNrsS7RscN6zhrhqYCfsTB6L3J9GTSColPbkbOjL0nXmD4khjkFoTZ0w
L63efubtknnPXvsEnAf3aZCmc4GvTKY+jmlA77QYDSa9DEe0C42iF+YyR9Hr8ECEAqTVPVKNXxz5
D34/NxoBW/EVknaOmpIww5ooAh099iQ1RsFc8Gd2Wz3P5VlONs48MTjwgGU5SYpvX+9HDoyZzVYS
DxqILWJQpbIFMjqdIf+KdRxTQIMcyvE7O4wfxOTE+8UcXaYuh7/TBWlizo8t8KZ4QcGXrkAmNwf+
DTQNZ1NS1/qv8WHIbzkWqBmq7Q8tC3AXf+A8hAvqBFVWcVpWjYGVNgfXu83W8vaBy2fNNUW8qFfB
WcDEoshgsWvYL4wgWpgsk4SUSU9pOjFCwaB+UoGXBKHQIuV7qSxVNUI3OVPklL9BHcWK6qy0NJZZ
wXzZckfKhjMefj1i0u7I79MO85tgIKAQkHHATXoRbGz5kFGHd7dr3yd0iSf54p14iF1Y0bL9aXpl
t426zIr255zjZ4D48x6QpoFvS/m+7iXHOlwk3i1/UNlu3hSf6Pkz7nKAau45RrJyQCfYnTqapea2
rhv8lphYOvjJ403roMeZ9Ky0UYlPhPK/FFM2051bIeTReI6QyiW3vQXaSj9In7S2XPefb0aHTRKr
U7KYBIOFrXf7okgP/tdnanVxjBVk70Z+TJyi3THNoWoBJolJ2M7Y9oYEilewMN+d8rAEIHBPTcof
OuT4jTdwAChBtQ9EOBQvmccg79k0GhT3GrifC+I4Hg5gNqUM0xccKnzUdVEnQyOmBVTLx6OtK1ns
R1SCiRO9e2JrIpd2cHtdJznlYwyjdo4cotXl3+IcJp2COuNKRYsk2+W2WrM91qIX2pvqCX3ztOFX
cqlvpnf3BWdzW1iXQuOQPOIgLbnLdTmtnBgiqRDIQj8/IGRk4cfuT3rxf1oMHRb4PihsxU4yVKO+
5+OcCAeEgK774GmcIfnwTKW8b2DE/SRETl8xItpfPOedmkqB20CmrG53T0YpZJHmwo2p+FPWtaFP
eNJRgy9Yts9VDb0N9Te/TQDGoKtLSlgiG2JI+5fpVUnpUJF5gkxCfaJxkITOa8AK5DJ8XBmthtUa
6G88T72/b89nGK/cS/XNWRfA/Fb3BPfSkV0/O3jyHZsUD6zcsqz/ELbf8Puy6/tWXo8NLc3WoKi3
/wI9pFpBIhnbZmRia6C8vJ3qzoKsJDmM2JuqBMPskkW7CRMb9CfYiFikMpN60LNTcnAxM/qb2X2V
Z+1wp7s8WR/t9GTZ7xzo7vB6VOuy41Oqcq7oljBxozaSOs/1/rYfmpvGD/s5zK+0C63ZpW4FxbOu
on64+UM6YbLMuE2Q072c+Ohf5NFQDjE6t0M7aBluy6ra9apX8ZcAN3E59sJroVP+SEj1VxXQOHw9
2VzeKs1xEiXSINlvWdZg8DPYA95pue6A43QLcLl+K+NItrCyNyTmkXq6syHo/Igm5I9hSA6QCVhL
YvxhnYtcGnjal6RA9y1wvIjOUyxBIgT9bRUiG8ZOh4Az5xOOLATUMjltDfwKk9l4e/NX740zos7L
ADizR97ZvBKErC7bSf7h717kcQEpmfPdnK6++WV9PTB/iW6ZFYaRVn4LnwJ0jyYpJWeUKD5gInYC
DEYewb+16COe1Ph2CJXtkhmVTZL67o1G8VoVRgYDDUrFB6reGRSJWyDTV4yJeJo2zf4CspMy7hHQ
Sw1G2xFJRdBUvkccBemxJ7mkPYt8VY3Q/xxGOXJRauwoDiPympmCuc329y0YUjYJx0kKqLiNLgJj
itMp+YEDiPEM0jH/9bUt7Z1kew9s2+Av86mGE1n9O3fVQEUNuXWYQnULCCEvsaCTYNeJPsAJ/bNA
MafZ8RZ6gDQApetB0nnbgabJnlmIiUvxpMRDuqFysT2M//v3/cVsOzvObnJpYDqslqc+oSaW7+3N
jUu5SKZPjFkMC6oFUrF/ohOi+WSw8RIdvfH/vB1gFEvWOzzLSSnhOT5khcgVSZrGhfwPpBeXeUJV
Wufl8jG5ixooG2PkI9CUour8cA73oZ16qiyBV2enVR56JIhOsAZ8sVDz8nus7nKTHKO10DUnpaE/
J22iwnfKtTKqMvuqEM/0Pch8FmgqAQPXqJrBmkhlTJFgB+Ura1swZbnvrgWUyFTYlcqt3CdCAhkq
25WSoUhcd32i+MWy6IXFY9KAb+2c2LzhADy9sDcHshsanQP5nsNPR8dIj+WKZT7+3E0ySLuTjhEK
KE/D9XWKBLcO1zSTiI0z1JbcaeOFCaeLx1O4cMVbk8ICGNu6hCaNZBfk5T8BeopdUqnWtORz1mTr
NkJHz5CZYqDNsWOwctBa/NiPTNN89XzD7hSrcFoR0qLe12u3RX35Pf6QgsNnVU4/5JvuUXm3SvWl
GM6kGd0ULDSGJ/Y7IjhAe4hIgqEW92BMjm2/MXgYFbP4C4zG6BBozHyNqhI+aIpl4LFLxMXkDqZz
+sTbNVSEVjMIFjmGUm3RI6mnwJe37A80Sq3+Fwd/nvyaa9niwUgJKo89QApAjw/opxzhJSLHV507
b+Gorjq1lFpbpkIhcO2PdIBPApTYx+cL4Gk8JrQX3i8UX240ArAjwaJNVYYEuQ7FaT63BNK5sdeP
+3nnzyuexQrmZb5npF1zth7YRsW+kwn0LDKI/thZ8zTtDc7E44ps/YRB0x0Kgre2f4sbsQ7ZLTC/
1WUimdAh5LfA9X+X0Etw1BWNAjJUuYsUv8Q/AVG4cmCW6oBZGaq8V2QmDikrB0TRkCUuP0bZTQ6w
OuIPwdS7QZNo2TVP0x7hQ7/N3xUvYhcYSHmfAj5knUk8ttTrdkxIiTAs5gl1doiAKB7Ba30aO79N
yZ3J9SCwe+GqGOIJVpFVMkOb0paufYQ8g5cC/z1NsFBI1pHzI5mb3hzuqlpGIh5P82U89CZM6YaN
7xEgyfBevytJCTIaxVXExgOmkrx28bgaS/AfO3913H25sdHxXZhHhe+tZT6dB/EdVRuE3GIlnTT4
QZMiV5ki9tNTx3qZbEbyFzzsxICwqaT+F+k7J7gHbx0CftdymBiZcth3TI5CkwFEaFN8060NnuTT
Hq8UzXT3TF7CxQ00zThAhHDJ47NssUhc9gwcfsftfYDf+thXBQnyE1ZAFmpAz/3M1YoKC2yDjCTx
ahYuVecLARgmKZmjnZZPA6IH6nBwEbNFJugH/qKW2G/YF/vicX6U7jQiu0fxhYlnejWooucGq82l
MWmTinj94emepV4HGrKyMzV/yM9afnjHMQ+XRDvHWXre4LUWIQlFjq3r7XVT6mQl4GZEjd1qPXmS
eEvPSAHVlhZieEr+LlmkGstSgP1um5+5S1WIvw1pPGETfpjsh5uc+dbUoNumLuY7HBhmg4lZE8Fd
2npbh1hJp3Py1OHj7pCAIYkNBVMcykSCEJYGkmEgeioGi6it9rvDnVx8Em+ctXvx5LYtpxKXgiYI
nUMcobaItAJIy/uKbUnLhgs8qD4OPRh3w1vBabyKJq6eTwzJeqr0pmhs0Y/TJ7huSuE02lQF7bZ5
pPCJNC+6x1SiFExb+dqBNuLXzD5UKFkiP6eHrTNBuUWGukaJYbm0fxkD7Va6Rmz+eunn7qVT2WVX
TvGQu12/3OeOCQQRbbLwqQfuZbI7vghkEuqfVYleXWgQsqghErOekQum2H+1WyyR5twRzQ9sfbvY
OWS3fwf66Q4C89xOmBc4foYVrb19J1HggkXdlmCZmXogumLwkuOc9aM41ZUHI9ElapMPoc5/fbCc
qEdGquQszq1G9y5yW9HpFUxutG33wF3Nru7tdaxQ6d7ttEXrfD+CFRi/3ObLi8ZWmdaoykOk669V
GyGKMzyXvkzUBKqI5FT3+aq/U5rnyn8mz8ri8lGxaeI+ehXlee0NZEIoRo5/4QHRd/Zzz/Z6e4zQ
K52myOLF77HVRHrc14P5JGb5HqDM2adTot9RmoHHQckjp5jMcn2n5mWAezX7lWuhZTJW045p8TWs
3qJv73v4xcUlY97OjH50ruaSjBGL0k8ACunhHfpq4l1K7JUm8Knto25l1XSkeXXUMMYqcsx1iANC
CM1fEhH5OLFK1HHcnU+YGxmxNLdV0H5GhMERe2s+ghEuMesqt/fKe76PHAGi+xwTHvAzTgRWthoZ
2ho511xrF5QXAj9TvE9km582WmFAKiHkQnp28iC8mJZomF4ZKrO6RVvaGrqsTwSiJDncbXnrxF0a
2gZDckBnucIJyrZDO7OHHQ/riHAqNM9PLKg630KYka8jRPvFW9Qt6BybwoQ719K9cFqfaRPoW0dr
1jy0tL3DygKsSbbIeoU97vhnumUosYqD8WLdooW/J5F6UXJ8ZuIZS3c2Szj+U+Blp4H9AeYljw7u
dBo41GBeAxIHnVtZF5q6infrLP48U8yLfupa7X1ZvMDP6bhAzt63E5vRSqx6IrDmuMOrCB1/Y4US
mwHuU+yiAlMe8x6RSewDckTZKVPzC99o0KgIxwebIeAaMZliL636FKoX0X0WzRc/yFNQy1noAJZ/
T2BBM8EUstYdOm6rkYcy1C+7jqLDZsdeUzqBjjKhPEY9KxBMkj1yKC0s0SikXwa5sOEz2Aqayi6e
xfO4wa22mJ7vRy/E+WXYR1jZBy9t1VE+yS0WDLGF2yi5Wiz6+0kwNbGVTZ14YVLHoNX4C+GdD2NF
NCv8pC6aNmpqPjpTd4teugFnPozl9b4SW0I5hy5fsLC6Nil9KUnUeeZvI0PqiJYm3irH75ybpf7m
ggbEfnIo7UsaiJGd72ggBf/FUbVoKpVp+XkLsbIhqxiphDCf8hzU4e5sZgFpy4PqLjrdni4m9sQA
HpD/IfqowKOGRrr8sl8gL9mx1/TF93jgzxV3tXVjcGHV3Ujv0CxQhq1MjqFPg0uGSkRKwnGPaE6C
xMJfC4LYKYAQzjngfl1wwSrslqaJRJ0JD0nHtZ7p8KS1aoQEJTbVthxpAikrMaAJqt/jX+o976Te
XcLC/e0OMLQHCcbK2NYEPuPUwz/8Wz08Do+uW9kJyNqqKgcQ1iIJzuNp7+FbUIY8b3Rrq92nX66Y
t+kyNIJVbTUm9e3npbbeSzVtS0h6zKJcHLTw8DnduVOYF4J82r3361tFbIDQ3isROF6lJwrPTLJ5
ESwOz5kwtkZXpD6Nm+PVeiJlwDhkGwuQBLVOIIO2610fzW+YIFxcSMC5kiVzwvo37EXJzo8CYgLu
a6GDSgZvDK/3s5RcbvFWtBZ0yJBaHV23JUr62xQOC5pNYGtplQcFSJl3iIQSaHgZ1E8oovSBxHUf
PMhAdtzAtHXLHKaRLxMzXBtH0dDla1wegXr/LSRV5wXbcB8bToGHIjgQlNINYNtxHBVW9pUzgYOG
Q3ncyorYPEqeIqlIo/T73FnIuq+CKgr4MSVveoyvAvIwCqkirQR9ifhwrsSOCA75PAfA7/foTrap
qTfZMzdjNqG2qbq56NJMukGuIPm27EH5j6KtNnUJpBpUHz1oCeWCYjZKjvOTeo1bPMA6hcxRKoH/
Ugdb71KyZ2W2Y0XHIJAj4vpMakdZjDh9WFZju69O1GmaxZFN6PS7x6BAqwcaCwjCgAHj3r9xqlWa
w1pDfiJUBQkfKV3dky1zVS/OtEK75GAMnQ2iAF2cIqx0CqPa1XXELMwaA8lY2sT2wmpheKtqrrQe
uI5puwqhh8KytIceuTzAjlcXjEMFiBkiAtDxjWnWeXGnZL6QxnQ5hLu/aZj98j3kKgzWRcc/qZwQ
rd5xGeaKR8cTb6eE4UzrkPvQPpW/JwZ1xwBQbvVlLja4WidTiLpoiSjE6dp6ZCZp6vWHuWquFhe2
/7mGW5fHaf2iktUsPCo+GZGlQLC2ZNmAeZXnMKGHK0hI1cdO+pvTlqcHn91h15jmPIFDulzfbuZ5
i6rsoItkQ1B33ks/s4XbZTzHmg/Kxx/iG2J+CJJU3KJId5BEsZS6GWTAlUiSFG7jsbKsw8RWwzjs
rYTAjsNd2VviZEwLSHqfhCuXNo9UPKWDMDPHFlTmkjFkBI9ZL7pXEx/Ks0KteWBdOALxE/Mb1bQQ
NPe7Et3t2GYwkIR7kYrUCf1pVm/p49YSV325xCNLwWGygvzXTbtDwArZ8aN5dXQ8j7osNjKeP80J
1Km5FH44AP4VsoU1IwgHK5mkVdmW1q/5TRQSMc+c22kLLPtZVXbFZU8bGdEkcj4+t0bdj+kIe4xx
BOwTh8HrSPQcUKVico0eN/al8wX208hp4u1RwZwKsd2g4C2nq5XKONLbxy+REnnC6E1Bd4BwzLVL
gR/Od804aYG/rctebhyOZktmos9Lx2A1FtOYmzSvgek7w9q5qNhED9p8nf9cFAFPcReErC1rbdMy
K+HQORjPshHV2FeExfegox3ohsKKkJPWXslxwYZrU/W6+X7T8asDHqIahEZk18XbuTvhs5PgJj1d
AwcvnGurLXEGcpY/QMIBmnW6Brx0B4mJQSyszJgqTH+2aVxEJFGBunMgg7QNtzWE6HGo3d8Z83BG
SnOEa4NxzCsYRjGpwXIeJjQ99nJJlYnKnWQ4kcFvargZL4ED0HLH1PFDXjXv/zTsitkbWiuR3lr2
yA3fRdWJ2JIpcsr3+NWBJ6K1GlgOpfddVrPIYoMhB3CDvGjM1lL6g96PogQBpKllA/SNnkv0eCb0
x2t2SFEkiqEfKzmp60pZw3QGcEyNFX3KBEVHGj5kIKj7GA0Vir5UHObp++egjY95uteTqnar/Upl
iZMkTnstJSOJ6H1qKezWQ8RWemo/FloV0TupG2ABcSWTMdExm11N0q/mPxNexuYxCXq+b5w9nf6t
3wE+1D8b0XjSmGhMLMFXvBHMtFQsLkCF9n4y74z+cqCl35fepcmNW6eRtEm3AV0rJPdKILCpFYPS
k8z+ff/UyruryCnmZc1GjyuAv+NN7LsQSeFSEds0Khjm3Io66Wz3Cr9gJWwLO2E27Y6p8WuLvkzA
bK7x3J0tRScBjN69aoSSXDh4N4WsTlHI3GIIaEGS1Sm827SEUhwOuIoniY+spPm9Mrvco9VIjJ4D
ppkdfbtKmK9GiktXz/NYtWcFDYUStr0n4oomC22ivW08JojI1Rw2I2fCQYrwLNdUdlWoZUz28nMV
BW7u4OeQpw3sJy8yBf1M5yrKUFniOnQh8ly/5to43j9O8tXgbnDBNeMwVcmgr97g8Mpgdf/LcDt8
ub0jMIgRgLOj7gCI3hCr9ZrQLfInzqIx5Xx3uGDbw5ydFfeAiFo5Ab6yZ3a7kVBd82Wq90NS7BGg
XO/qFm79INCD/m/ra0dfbRURKIht6wsyh/jyYK+7V7gZ10/A6aT2hRh55fMk85CWDci4WtVCYETi
o1dl1yXwHz0juFwtJX7+aIYDBnMrheqE9op6epdCe9dqXkC35LmB5mEWkRnOs9HQS9MtlgSMmHUa
xtOsD/EHd9rxP4xZcWQdgVr9qXAMlWx2jIMxkFYhxc1JXXRZitB+iObyD2icCApTHxtKR/dmGp4Q
1GdpUelS8ldUvtDorEuDArY1/AKz5jtT/16KTA12csQJplbNYrenSoiV8EwXsXykxBoNla1y36wt
uKeKQsGfIYdP+XqPRwlGyWbBRMZgMY9KICHTwvmyPrsktGK9m4zPy7rcuaSdgkmFz6baiHq5G8A3
K9d92sXXu7LiU6N3KjlGAUC3oB7RsX2JTqrsijLSgF2w4jgZPgFRtpncNJ500xvrYhNJf6EELpSm
zqY15/LOWECfhFq80utszXn/O35PzahJ4k0Pk2nmpFT/jC2NzLrOSRoUTvcwBz1/NiuegoNWh0WY
5ZTtsHQ+yLGZPAAcD7onl33thPiCVC6Dky9KlNO+TZsl3hzFCyR7n20vuglWxbb91TjAjLU+pD8h
Z79/PnOBE51Bamb8dAadAqBoP98Awx+aYxm5aTvml/t0CEQ4H8ux7ENFfMCWC+IrP2wa0CNu1lZq
QGVwdnEKYN5CiyqJT6XRgAijR1cU75cDXq6/aqggpA1hbJx0ZXJA5EG7C+vgVEX/KVTIGtGIpOSf
3Rx26+GnxOcn8rZoX9+Uh0r5AlTmrGzE1bIQREncrOcDjxJQdws5wP+gkD2dtyS/LK5Lzeh1P/0I
yNAaWXfY7zSb4IAi/iq3XToj14Dn6wMgxfru9vBZ7coytIZY7b64Tbtoqu9QTroC+ZUf6Dc7lp8T
VpiBrZPsC3EzwLnSZ3/D+18z3RNFKbBRorA81DRD8lSz1z4K7Gzrr2dM+8abSvDArGEHthCkm/8y
cS4EF6qkviJOEZhkk0OuBUmjdsvsM1qrAGtw1xTsG38zuW1n7kq1y6hpg1iitauab4nhcG0pNX+H
IK9YIsPNdvTOGukZ0UFbziVHquUhxtR0BpyYCZXBWorsSTAsm+pm9XZ5jU6detlVpP6SP8nbESco
tf4/JAAQDuhuK1u7WNhW3jKsZx6f4kzgE0Uwc2LhcfD/fwMUGWMfO55Qgjo+FYq1OcKHgCEqYEwA
sywdifN2SJPGSgC/erNijFvjWs5OIYlPpllFyzwUhLrje+OrrYq+Kd3kVcMjLDGZrtE8ELzvoTg8
3RGkzMLfescjmctro2I3FXrWfRNcs5+hI0o/UjmbHN9uLEt2rjfmHVUATJuH6qql0g7KynDn0T0H
l/rdtii4vcCIqcLotTAIUcA3OHryWFONIoVO6KsbPgMFmcrm4gVKwCdDl5GDiHMlYsTeFUo1cdCG
o98Ur9mUuxN6tRp333qYoertKo2imA+mg0oa43Tmq8R2fCfxIjcQ6yd+PoNf1tnuflmePQKIvwD5
GXZPnDbEVkc8EYADiSL9qZ1Jay30nrM7rFCNWmdzsgJo7+hodQPhiWT/XioB4aGKk8TG8ee3UY1e
PNpOzAsLYLgSGk6Pv/Y6JXyijtM5s8tfrRR2nSWMUFIjWpDO1mxPlFikSuUQh1BHCZJhShhKuAOd
7AI6Ci/+JfEj9nLqCqAo49p+yL6Vq+9mhKn/VEm+Unr41sQK7wrNvegq9lCadLFN0gYrdlUxOtBb
Z06ANGxAa/IB26XDdgkqkYcVf/1gGEBfDma39/Q6kDqk82rWFTXfFpThX4cwTN3L3bk1at8tkwsJ
eoeJqrFWd/y3tpnmsk7YC+U5bFMKscWhFutG07w8zaqjYagna6X1BWyPw1SPkKDq2DwcOqenCs26
MMcrJZSu8jOSxUoKjjtOp6RE7zytNivmnDcLTG1tTMhasgymXitDY/nRrliSIk0AsUxQCUkPhI9p
EMyUSiSUe6nYn4GkA826f8cQkYvzag5g+f0em474Ae0e/q8oVb/pUSiqvgk3evfhAgh6SAQ1WpS/
HSK6nR4aOIvE8GBid9264nZLEgVNduUjudr+voo2zl6tdj2L2Jl+G25kMM7v0YR1ER3LajkRE4JB
LpafxoEr0yor36T2I9rAERjDaYpdUO6Ih2mvup21mWuF/TTo7qscS3qFQVKgxMjcBxvpg4rGo1hg
fcGBNdNURKpZP8QotabSTLbhYfg1oBBEA1SR2vku0qBHKPQvgsdrgkK6zINqJKjQlXP/CBeOq4RY
Fj/hDQEVZhjRE1im0e7WgnYBhiepyB+89/VvaTmyrDcfmoScw4A9eVZEGr6G+XOXfe+XGrQcp9yk
nai4FctRoE2gfaEEeDbXY+SgdlwEzanEId6qqE67RS20WTHp6gpHc6Dyrg0Dudf9gV76VOeZdD+M
LcOavR0TmgY4IIEjNrKfyqEbBsaxR40a1b0ijZUw/XvqQySFcGhCb+NXIyYJndalaZGDfUm5qimT
jtHc/5xP0eLkyogMVvwcl6iMmhihxiKqXylZdFtzRuGVU9/mSM3hvX5cjcl/CUhHU9NBd54ek9Kl
NSwBbJASFCYn8eRNKrQ5HzuPrIaCH2b7U8EfuSfWiP8BGTJmBOpeZtjSkyQ/VwdEIke4QUgwuxSJ
2SUaDVhupAQ00284eyHWoOIhr02PzY56RPhE5BdbzOZAspZoycXVebykQrwI230R6Ut5C3Uom2d2
9RhVZqFK6x2dB9P0dX8xiDMqJt4ZdBUsLDt1ekGqCKBRf0IQFqrLb7NOstYsT9Z64e4DJBRfRV8j
KK3/JR9eumYUCo2MteuW5xml7LkfWUC3laRtunrEMKYcLh7OlP51AGQgd58aSXG0URg7VfodgHmg
fus485G8vaMnubLpVPQsGdVlpuV5gF7cztVcEP9JW7tTpTNxnc+LgQOfrAO5rIK7IZGaOsg2s191
4BpMDA9l2GHZRapM4Ab40jIF5ctOsnv9vCll6R40U/PP7DCUQ43VXGc1i+h6c8Ra/kJ8Z7B57syy
pCkluS7NYqHuj+AN/axwFR1xrVYkOVHmyK/j4Db17v+wZEMJcn1+mKL1UdGM+zegHJctfhBREaR0
GqZ+S8YmHNz3KAOhbtPpNjPDgRXYTN+W89GoR+wp67hdUKwpQFe4JFXq8M8+KTmK9+ASPMMZcG/1
++XBqmANBzcXEuStpQB6THW4Pr/zABqtFvWsKisltk9AVWbAai6GOpZXGjpVkuXmtUDawuaIM6GZ
Eil/hEa3Xy47ozewKkqU2sRr5t7pgCIJFf4UAVJeyD4IFKeiQLWzjE29Vs+UvZN67edXWXvA8Mgh
jiqqfBhn1BmI46mw8gbwgqgbN/Yz+UtCUC0S16KUoYglOUW0Js8ZaryGiKSDht78bjFVlGacfEnb
fjIJbn6SybXTKZaTqattgW3OeVla4AiDct0KF1ZZh7DLrJE+dryFfcQPHGusabAhkHBv7WJC0IoW
Ejt1+ieFqj7UmJb1wiWTkrurxo9mC378aqZf9JGZPGbLMEb8w7YG3d7N2iOJ2S2ICJQefqcz1ana
tvVZswfI1XjDk8ontK1M3bixD7oolREg4DU9ixvqCa7FH10aqKwjLjdwWcj2iMr7CQvgMf1NmxPs
RwKFtEEWEWn1ZyKxQrEqzY8A5dO8XLeIpCaqQfz5EXo5/ALIdn8j/YSEPKCJDOLb7mo0GZ4rs5jU
GzxaVtR5qT1VeIKOpC+wrUZYSuocRZXVX59SnosxsnVmKRb0NEJhD9rCX9Q/nIU8kWy3aRa81/07
xq1wK7026OMz1x9SQ/gbDWtyseiwNel0pmLykQY8p+SGpB1tSZl3i81PYeznj6Z+jWp2vgxjiZZx
7/dTvMJGJ9am892OVqDaQIs/sIN0dzflqBqsyLSN674Ul90rqqGh/UByJr4GNN27iXpV4vQ/zHiY
S8dtIVMD4bgpDjrsseC1su8R9wESpOB28KJX1hGwpHiVHPLPafXeM7D6CH7f8o1GuCHbQMS2SKBm
KZECCBAfGedsCSL0RD5Tka+GWDcsKyfh/d0Q3A4uVlzeT5AQf7YKKhmZMtt+cn79wczMHW6iWTzK
lfp0uPzcB02dbEfETd4OifrVyuQLghoCaCfIgmUprf7MC54W2+fbcl9QuGwFfU4eD/RAnzX6ReRZ
2gMv+LLidq2vuTC/n4PL9+08YmbOopFwsgewL5YcOV51w5oxCl/La26AH6UVp7qUdCa/H/1FaHhV
NKnzDzk/auUbicUQSiKMiiDF5v8WaHiSWVR5r4gRqXiOLkVnI6JYJPR3EazBi8SfEUIlL8s1/dmf
nNcD/kOKE9aeyeL3WGC9BJts5gzjPbP80fqyNwle5A/QOjqDGG8SlzO1yXRe5aAkSTOBsZddC7R6
2AbGGwbSWG+IeolTmLndoTGC7iJhK0l5Tr2fAy4KXEavn8L+lSAVsvu637t3jztNtCSVTaRT+/qM
5nD/MZ7LqfJVCeNsLDdIZc9y5qCtiDt0QIDn5B8O/CpLXAbwDtAUFmWt/ihwHD7tA6n3z/zXziJs
xGwY22arnKyOSpMlemvkeDazpXT0UoKQj2y/BG24/ZbWa6IRY1kQyaNOwf1BJb+BL4tPnhqcgf/P
E00Xhj9RSxKHaqYbwVIASgENBivRpz/s5rywgoRy4IuSZgcIJVKUsxx900x1WYCix16P4Z5MGayX
MBlpw65/yOfh26pnxeJJcwbQCCr2IadXqkdUdXEItCu1jAHsIvwuoHPe6znnN+RZ3LNftO1vgF2R
mcxkvpXscirdUo44rIQdbyP6ERphwrbwOhDP48P0gGimc5vDCCgm+HIhLiUp3zXcTcVUMrE2LO/9
UXQOIDmxbgKWt1cEv1AgQ2i/0zaR1/nV/KfkSRj7ubjUILashEh8XBk1unkzOgMRYuQOPl7i76BO
BF8Bz2KHljKzIvqv1rPvuhbSekeygLQgl2PrgSR5DCAQFeKXAH5XDFqluB+FEVcfqWCuYhwwrMXO
OlUVBDKLermOYI8pgWyPZfrAQpxSTnnt4CPWrruUsD8Jp8Sy6FoQx1Sw/4NicGHwOTIX38wYkO55
Qbc9z1qPsf6HfOUa0bHmgleVhIWCUkAFKsZ1bxqCuRYqOxdxuQGMGvYZEx7H2V4MYLaEby67nBdH
jdupPg89Z2Zy9G17nzgCTlS9bRyX64wiWkD/1ASrBiHazeD/0dhSQdJvGckp1ey33t7aQCNDCBGu
ml4cHiqbJDycN4FdU7c7ELJGj6RPQDDjbWXPd7ecTXsw7m4MmLdoUA+Rciw1iH+MKaCxwm6cYPl1
1G85SQqjTNHNLuToLfszgxmtfDMKbbr2YTe55MrhWF1ny6H1L9UI1fuRjGTNTEI1rEv3tQPrKNaD
1b+DYbNEC/kouVhPVBDtCREbpz4JE8jidQJgaJNvSySCZAakmFFxROPHJhvXW5eDEaxadr191v/X
xk2J/M+zYcSKHt+RiWeCgmD7UeMbL9egidnzr+9SwF4Xx3b1V6DyGEuDv0IsLshvmy7BAUuCIZXw
1aeBte63UNlHK3BJhXtEdZNpYGmofkM3MA3/Tz6jSrgECEl9BxKiFJTeiy5v8O7mBz+3Kabxn7cj
oXzEqLJXkAgOJDrZhDUSACyUSUe1dhhYB6PPnq2DlxCSYkhBetLe3G6hHXPLjaPHnvQKRhk1LOjQ
W1Hsnb3bA/Igkx6IiQIownEseo9hmccM4rcFAFbLaO47V3skHYgBlms2AA28qcDVZ/KOR2K3eFg7
tbAmYemxTttY68lyfFTYVqN9EIgfsKvhNS6lrSSqeMwC3TrmOqvC6oF8+f8VG3WwlPMkCQTWY+Sg
yllmURcV+wm35f6+AdsXhSkgd7AFVBKoqjFyo2NQ/zs8nHgbjiRtbT9Sv+240b1/6Qh62zOAxfzo
TfCkDBOr95OHghwEef3w+JXH523EtIo6B8yk6e4Mn9FOrwulfl96avbfxdULe2UAMUMb364NbNSw
/yLmMc3MGCz5VFcizIMi4ML+zpD4wwCMb/1xkI87VJhUSoAJwXKOLaNBMXQ7tAPdbYVHB98UIAdb
3qthNCBtT2qjeMuILgaJBHsF6tTUGlh+ib6LYtzZuZVYMeSdYtG1g8xEiP4XrT0X4lGngXp00ejC
fjUXZwsVoH0FMKQOG94GP7tTEdnBkp0uR+fjW470QUEsbja5ivw8J4v1sZM5+1RyqLy8UQzkfr3r
GspqRNKvZQOpx2F6x0XdhsYDAxA2bKK4ZWT76gZ1uKIehf5DqUb+IT6rLUVy+YYr94XGp6tOWDXa
pg+w2sEIPIEqChNL7SFA+b/Eto97Zv4J7JVVvcCEuzbYjtUV+Izr5fwhKaS1q6LidLUrq8qBDLLk
+hiGpgdhoVTjP2thNroDbwW8azVm0rGWfx1rPM5kBRdIoaL2HmJrFYZvkB+XJc9H7KpT4FPiQ9rP
AWkeVZE/WataZOaip09jZp7zgBYMvLbVrGEW87KlxHidbXikIft4NQYNswCxnWuwNi14dQdItxti
8V0laFyHqXEMiBXhaQGLEP2rgNSLQAOzMoPljOkg3MAloWZLOLInQLRrg98VPTgzZw/adGnRJAmk
TNWtJLVDe703kACnWCwbqTerjybQXk5WvA0CWhFEo2IsO+AgtSmmqSsNFgA3dyrkEgk4LVG/aTX2
dZxjDUy0XBRrpLkyA2c+iRW2AvPSS5n0wzlMB8q8b2ZiSxYETBI1zhabz5ncMBUwGoU+1GEe9PDW
w0V4vidB+fk7SGFsn2HTfdRFA2WNA+z1oYdwdJbUpLM4jD9A5IqjhYAl5t97H1a/gG0gECu75Xo4
1id4ArbdL5pgjSRu9Lej+ru82dHN1GzQX9VNL3cnWHD0lSWjhZTVk90hn0lUGwciPPffY1jWbLkM
hgJHE1OLygayNeMHgev6wwGsK3DSl+hrhQSe+L5BZpRdoesvJ3RJqOQb+b8IqpAocmnGdhMDhYym
FAL9u4qE7RtmjmFjCXs/L0EaKVGXjngPhLwU6tnuX3vTZqTYzzqacQOD9llKZblhyWGMAEoUDV0g
+4c8QceMfUsBPbVmiseZXfCu/iPuK6do85d50hmyv2xVsko3JTEe/pArRZ2TV2q43thXwvZzAcwz
8dNHJCP0SVgAfn+r5gudwvFnDeQAd19NP8Ka9ZRTnkQnjUtO4S3vyjM1iYG+v3mesOn3Ajzjvpwd
5JQeURq3xE/3uPI3wfwxLDv3F0/NYzp+VbiNHgarcIbjaDG1BwfRLhsc5Chc/l+dkSOH9TT9A/QX
QEjD7Gc5mj+h2Bq4ri85Y/ITdCN2zhGtXOwhjT/6beO2xugL5CoDN0uzwL8MJ+VfIcKTebMjTNxM
NBGjJQMZ/RySHOyr0P5CCAvJhI2rX2uMFJS7apbcFG7DeeqBAeFiTlIKPW8d5h/moZkSdXr+E9Qk
DkYcakhLVPESQJOmVFDWvpipndOoQ6GLUlb3+MSYlx39dBHa42bX1kFOsV8J0RwYb9qcSJfWnaVj
FibjV4lnuiZS9MnCuAasbi/o5Xf50xG5epoYBoUESzRA3Zuu+BudUPKVjBTqgZA+Y5mnBuM6lhtt
fRAFbN1t7QJ4fVhbhTSMjW/xlk9GMNETeZPdEq82jd5IeZ7q57GNBj/G2Yalrjunp3DsgbawujgF
KqWqOdnPTfaLfnLoDxW/R/aPtvnWnKYlX80Qg9YuXqCLlHvJDvt2JZyqsKQmtxXfnCJarzaMBEad
m6zrXFHKErhRMaoBHBYy4quABSAmnb4wW8xwpwYinHCaaB5y1A1CakfzSTR3xZTq8qapjfMnIAaq
+Ao7B8PyT8dBZGQfsy0AQ8ZN5FjAsn729dvVG3qb4r7v80VmYQOHqgY6k8yzgMyf5W/5U2UF6EIL
EJkdJx8ivw1BfXSHhr4C49XcZ7HlsNw4wSHRrvMqCUFCj9lh3IV+MWwgyftw1u+P7ecZ8F516oJf
GG46pmESpuK+MNC1PLrna8iP4H1PgQT4LktdPnk57s+VEaXX8FettZ8fOF6wfEPBQ9TOipqFiAqL
nJsapxadh7+5j1I1oe5om5wvSSrWqz+wTQ3CEnaiHNIY3/2tnBOI4Nzz7JntlSveLAEh0dopee6k
80qMqa/mVBcOq0NbKS+wor6OZXSeQQFZnPjKe8MtQrS4yVhnvef8vwJ0OHuZkNXH88W9Jmvt5qKF
Xnzh5KsA2/3n3aPdwhiIq83LYBb5E37kuukxgdpEu+CGSbr1GzMwEYtP1enQiCG3oxE1U30g8yBj
OGydDM74gewReCwwhF6drc8Me4DotIwICjI4L4lqB4k14hij990EYvbnC9YcYQ2rLBehNLd0k6eQ
aEANk1v5fqiyYw8ENWJ1C7hAGkedO0kjRyg6raRuz8bZQkANgX85VExKjBePEC10FG5WDupiqVPW
mj6plJ4irFWCnTt35FZu9DEGQIUrvPu6IWW5NJ1Kr08Ow81osqVYMVQw7mT0obRXgJzU7pSwivtA
0zILWujKX49SNdTeoWw7mhoVYBaVTcuQDx0emZVOd9KyFwa7AxZ2kW+qpkliJYkh6R0zF2IkHewv
EVBcJ4SRmuzpvYoGF2SxSD91Z7ttvUIadf8IT/G0r53lMlsOLJebALMg3q5jy7TA9VowZpC1f0PD
hR2FS5SjTttl1SrsUdWHDXHsaulAERAMV3NmQeT4xZa8N0j5n5MZrdizVR87VNjWVfSb+5YGimB3
V8jsATzTFfueb+0XX9WSdTkG2vO2sRFzFlwbgShoJ8gJpeP44Tblv1aFUz4F8xlQYU2bvKQWMkVq
sKsKXxdHA0O9JeIIrGgW/AFIroFWh2hwJPSIxBAfipshKexX0avxDCIp8IPQi4ARxEWfUP8gAg+p
syywwgtU06pEFtqEC21N6kwWE3oZleM9Rt+qpqom2HqH6WCDrrw5y8G8tD8Al05HdAmQNiBWswIR
0hHlG2073cnf7XSwkLBL1O5ZBFLm3iK0U8qZgBO7ryWOqIXSwxCj511E7r17mRGzrMybsEVsmW/T
Vcl7ix3WG4dYnZ3o7mLfDBvbPgjugb+QNMDe2GQbLY0/5+UIrDyb5jSnYc4fv4CWvvLwgYCUMujQ
dOCgokX2j7D363FR2N2EGjPY6hl2Luf69vvscqRgE7n4ByWdCkpjWgLjLFRJkSA1BLEo/gt84cAp
tLWWokyY4B8Jfo3tue5KNd5Q0athOdZeMYNGDBzvToAtKjYX3dIM8CTHrFh4ND9s/Q/rmH/rcSfK
IvBKg3LHBzbxz8hdldzCV7EJfNadTI6R80ns3iwksj9C+ayfMlUBjnCvDP9Rb+OCt6/nJ9SY+oJi
A0ukuR6GlXUmOfdFJriJTICFwu704EItWBJ6DcKWBixfONkkmr7GO9EI9JKQ2PRkpPW6bhoghS8s
pbdMgvQstlOHaZSmPeH2+4dFwpyNW4eP/Lav9WJCpr04lfDl4Nurd8w0kBRoNXYkqRHwDo9oGFrx
fUy+KJmC9TmPvbNi8YQ8InHEjQ7V9G4ofA4dIG4k8hji7JPXoPbuX6ittizf0C2PoFVFiIX70z6a
iMYV1Zj8F0azAvXuTscM7LDjWR8POiUCTYHCwE+Qwy2TqYD11C0HVwUyABn/I4Lu46gTGp2eOdbF
+7dbkhZgeyJt/J2uu9dSpOKr/DAeVkGrKJHREQa1r2cHTfSw1MyYzdclsQ/MDeDKpjHOrrRe0jrn
85LbuKaGdwgLyO3cK445wnFvgUMTj6rSewH1TjwL+DHQep4RCEAyMTA6/zjLcLAUVMUMNj9wp382
f2kPiAA+6PAoroa6jcc796tWcBZtVuaY0BKAxSBBRuyUa5w3m8vm6sYFyU3UvKKFmQPTEHxeAJx3
9Dt4/vjmCEbjQsSIPzYr+okO+VS8hvR9cSCHpv7sa3hLi8wl2noBJeFdJC7bJWKAyHqty7x7GfLp
RiI6UEIdOSNeCzOuC8V3TVUhyPv0osL5Dn1YCz1UsO6A1/vaSgYx9kMIqYQwk1Oy2CzP3qPPT82V
SUyO2yxae8GKMKCP1v7U4yfOKjevyX7Qh5smDU4muG4Ni8xJxz9VBzuaQnQc59W54azu8JtgVdWN
WGyfC3cLy3IVYBqSUbCGRVl/tduSYXpjI4hqLIh15tCnP//oTIY3UtXZSvodxkJmpg+DDw9nBuig
q356tDZJRvchjfQn820YBDKe9Z324DpFNCnysGE7+JksPgFwlXAuoJxdupKTacr1UKhrdmy0qZ9F
OfWHoVd1TmPuVHmOr2LWmnIdgxF36ZhX36fKpGqhekG9haPQFwzXKNzZ6b4CaPvW48pEs3jng0TN
o3BsM5TAhce+lB3vqwww8ugBe1eOjpHV7McMwiBmFBc1u9bIPewVfvuOQTsrTBCzQi5YyulD/cOr
uZMuWp6bESzDQcTypvT0yapy5wNFlkG8qqNZ1wgHkGep8vHoanh+yQLMS4lYNX9QvvB1qx03cAVc
SbevUfTPkbiSGJpA7vrUHFNv913HMtDLF4gQ46cloRiq75L8bYlmmLmh2aKBaEH8iV0QALH78KEK
lNUPo6gC78OY+aeVoJtcBNZo6QCtzFqaN2jvIl3q2sMXO3fVC1gvfMHHVPd7Jvbf7IgUomwc8RIT
FxOZS4sHy/mEK6vn2aWFLJhP7cTeZvIVLwtyzIWOCG/Kh5iveYGUKjP7GJLfgk+3MdUCZ9HfI31P
j7OrbTm/HcUnht2O7ktrez/dD90xNfuYOK3JpLmFX1s0LZyEowmBmociBpB7sEQIO6Yr8epPY0Gd
B2aWiC+bObsPg1TuZJLSYT6mHXkzxYo9m8uGuN6EJhQOCqQ1pPThShueZpbi7DeTXYXB1HZCukWe
n5C1Kd4FIzmVuJH5ib51VeylJJ8aAGEFR0q8wkBbTRSKb4u4Kx/Kw9trVLn3bWUcvOoGKNtPIIkv
wXliOknhXOdrZesBF9uEZ6GzLlrsNdIwwPY7w6tJc8Hn3/YI/bigsQ0xVYf6uejWQueyfM2q/EJH
3rzTnSyUInfZyJJ6CzqNiROLJ0MWCeu3RP7XMwKvyshNTF+jv5J+jkFITaexxD7cj/VnB6qbzVj7
rNu5ma+Bu8McjdKatUpDTdlbVJpQ9ouyMj/AHvcm6JrxllDavguq9vuSQezWhrjCzy7LGk/iyqSq
MeSSjY3KAAoegXywZ0buO1z8KUnBW2CUJvXg1jEQlr8J9LfLdGaN8JGr+uL1LKEe8afljmbivNUQ
s19djyxaLDy5GzNiwxw9hPQioUJNPIXT9wH1AyBwpTY7ewWvONsYriGPJSZWHrYBo1JoQFuPcBUn
GorIlMXBSem2fwOEJxoMXX6FPaykzMddwnfn3IUL/XpXgw1Ymz1ITbJe+pIjck7K3ZmylhVRuz26
c6/w1nE3EL8gsvCWw8x3gt47CiJpbSIFOkYCptrhB4A7dTh6Z96JL1NPJESZH+hsR7B97uKNi80I
E2pDQTk+Mb/DQhBh+c3Y2i4b7TNeTM2H5c44nzX+Z6Lv6feLg2mq0zlF1O0YHzp7JKvUgGTY9+1g
RDpt/jC8OAJ6xs58+MjkSMrOSsg0jnE0Pcbpm+RIV0XLx8001pMbwEhI/BtVKdzLlSqSs4/vOE4G
QGGOzlyYDRwdLL5Uak2USOCCRklLXeFuon+ZkOHZTTN9D4WXyRr5glh9FmcF0bXU07qhXZOy2/od
1/4ExZ/vqlciGodlFn4ICgDIVcFR3GZGpO8b8Db7VOhrMVYeiB5qFhWGJ1tv+Omdv9CIaj0WNGn1
Vt1SwiAk02OO/wcypTiqMNMmlNTuQtZ06VEGqt0hb23qo3UqEAWdlHkMnUjQMCkG7F0i1GoFp1M2
O7XsT6Fs1u6/PtLjLsXZYNM7/Rxu2S4kauifyEN525GiWNqOP/JKMwJWZmfafXye2c2p2w5jcjvi
T0hIS/zAtaiVwE1jbLAOfDXHmKc5TvX+K0XQNtRuSoeAVoorBK5Z2x2Br89knL+2jQ25ceREs8yR
mfCECbPD9viY+fkIPE32HrwxarlpW0Pb9cCYhzOgG+jQfWXhshbgbxMEk9vtJzjSjNaaOsYHZgUO
wk7VDaHZ5mr4u72wCKjwXSACTAZ4qdmfAM4wdNiSIK/2j3fSisRVpFfTLBVtS4VJnQExtm2qGkhj
RiyiKnadeHlEwfB0myxy9i0Hv1OTUrlZWoRZJ372qeb+WyzAz7tJrxt2TDeqYC4SeBf+Ng0qwE4n
mr2rBNLkyYTt0FZVknKBYA6OeGkeSOrSv9GTLAF+lZf2f0bbbGzXpXm3xhkkvJcbNvJLwwGs6sw2
viJQGcNz/NtTndpJMx0PVDzruPiafc1vmXLqQKrzgP13df/cJKkt/1z2L3NcksG310PLSg8E75Vx
mUOdzmHQzEaJ7i7UcHaHJa/euuGmji8ciWf/qrETI3SnQXfXXEwyBl56cU9Igt7cl71iNC43Wyd6
ZxyHxfiOXyhWpkM3i/TGnqPnSp8wsdE2ZGYHMYO35uehTkQymBR4a++qLgP0VAfRsuWYuJb6ZsGe
NfYmgJ8345LFSOjLJEVxk9n8qBAq3X0h5P0jX7FBBeuVNMURhT26CqMsVs5ONg4vXfYtRLHht7d2
0tIwdjligTJ2y1mfjSwUuJRMDN2YJljbf2M5vtdRuqHSOtOGB9JmB8abuZ3MABIncpWlSt2Mx42c
Z9BkReXByjMhPorlJ4+WgOfK99kWFoOCs3Gmti13EInRGgZw1PRWKn0xm++lfnnLxpk5Hg18aEm2
5PFTbfYAM7HBpiGmRrwljMpBtOD5ilRXlwPQUl/nh7fbVU3k+OU9IoyTGoJWwWXY6nIEYMsNrzY6
HvtklbKLEZCTG8jPM+NawnxYiOTBvJIBU6QK9twTdqKPDEjmudVogZrD8mTqtd5KX1y6NTnS5KzM
MwmZfww8zgo804jHNdRPIp+At3acS7mqicvZ1WGI1WTvuWoez/iC2WdfxNeR8m0F5NmaH7WnTrTE
r5pwzEth1jnhcXeyU8/itcB91hB/cRtI8umfs01R9X26EtiwS14SxMAaBIpwKlahb0QSNru2DIHw
oZsbOFagLfamUFYJvhXJAQ7cb2bpP5lkQ1F2q9Laf+NjdfDuT7Q/+otuaZew38+em2xGrhQWAQv1
BW0G8mxFRgBiI7J07oBkjpFTiT+g+RWSlR6Jor01ZBRlBllFkcWA+YI8eZJFzYYwwKI3b+SqaZ2o
jrsrHGnkzsFvS0iQWlRS6T0xRnP6bGNmdImV+aYVuKO/F1b8hiPBm1P2aCApbMbbSMyA9HWAaXnA
Ec2zajtEZ8OGov9zlWYEWb/bbKNBXbPBxoI0ddtLl04i87FCnLViaME1zx93rE8V1i3Ci1nodD+Y
yHRso2QNI3cNyuvqxuEwXfU/F0UEyXCf9It4dinp451NEofbtXfY62rTwFXR+Ru+N3gi/x17bv0A
yT0Qt82hFl4kBqZ6qUunVt8XEl7JsATa0KOssoX3Qi5NfNxNr+KNNiE0xMPXL+/gE16bZ+tlYhQy
YpInb6oJxek00t369o853LfFu1lJ3Rac4gYIWw9aSirsOpyAhqJlrDL3VhVFriRsBRoEutG63NA1
hMnc5yuEoJTaZ64Xl6qhYrhpww3Ee2TgF8olbM4ZkyPkcypKBbPMCZGxelgeXRxjaDtWEZH+kgZl
IFcKsdVU43EAjipezR3Bp1zWwNjeAGwJSjTybzs0tWOKGDkFdlnMoRFLpnfHANVo9oqSEe4HJURP
g5UgENmkRhIbOP1UFQG6PvAAZQjvEC2VCm1gz03EWDOdJ57uiBQB84almONDq2EfbDBQmRNQevL1
NvejDJi8tTxMTLcRbdS6FH90lmi1kZxNzTdiuY8ZekwbE/1xcWR1Pn8yWLhw+S0LDDsHXMh/l7PB
+ziaGq+dOB8OG5Wo15gapHyP7JvYdnmIVX5hpkpee6GKXGoLtw2qXClz31Rz4dEPJe482vxiNx5h
X0mLp3XQ/OAfUA7W7hskGvwQl1tIZCsTLxPHCYw63Q4JbNa38ztG/d512ox1NfnuEqFhlguepahv
nL/oAYWe+iDG7TaGQgzkBvDFGhPcYKYqHdIpoZRT5+cIV2KkrM93aodNe+ered6nNB/DZ04rqaPC
WZXivpFSIgcodF2XpERuH8SOS8M+E7JN2bGxSSoNadRV9jdfMnrcQsU5PqyGvLVwuS9czGGcK2C/
bpIU+SjSw7w6Jq3+022LjkbUwNTbcxvfZ+EJC7uDfRFfg9CuoyJ+XZvF1TBVScApco3RiC9EhCgO
sibjKO39dr/tphI41B/mzzIjYxmpvka58i+yQhL0/+pHYIdRRYKrHe+vCeRwNDoecQ1awOffQ3DC
ndkL7ZamHiNdPxCy5kgAFKWFTWvxV65sdus5hPN6Y4WiDN8cGlUhCyz5u4agoEPBtV7sM63RLjJT
pgz26ZCVX/DgoICbsXsr8+UC3DI9tHxjKyyYnYiY1nU6/fUrruEpckfskW4j44w036ft7Epvvk9X
/2ZPD/HFwSk8/FZpF5ub5q43vwSnhQjU1HGtBfN3UBlc2EcFG9qnaXR2GJ0tM3OWFKo9ajdVwKe8
SuI4hSc+dVz4yxoQFSPhWzi93u52xePuJECxLaGRGobVF4OeWXGC9C3zO6iyh2L4ZvOctvDgyUBY
DGLbS/5Rw470oTEAiRCFSrahbnigmlKqB2Vpul24UT6nHczRw5iZC9vHmJqnXy8cWh3vaXabvoq7
QGwIqL4wejTwFq4cT1Vqytgn22tqBY6qiUC5jvS38kwm6Cr05nk2BjE2w2vYwQf6v0ZKDS6/0IOl
2VnLoMD4H/NpA/X1Jb31Yr/qM4bdqEdLWhsGduJ4RTFL74PxP/KMQK2fZX817TOF2boLWIoAkTUR
2LFsJzW6GQWZ4YZZ7KYbs1HVRmd50gFXV45/NHticPOlFc/0VK0FpPtrfF7+S1/QbzH7DrtsNZTe
UVQiOU5Qg99zrGUTYwE9nECuKxrfv7W6d1dIFafKGdgUc4RjD//Ql+nAmzhdVYBxY0Sdm+/jM5nB
GwVdD3LUS5wm7KWsmay2ArH71GSf72YyQh0WmYiG+A4g9Tz8+4XfgCKztPWj0d6bGKzPWJnfqPNY
vQf+jBZFPin9hzHMthxGSzh1f0MYwgUZL4DH3mOkDb5H/DYVCOMsEEi+BZL+sRr/rscjJvInaU6a
ELmSWsmBd8NEtNpweZwOA6rYaho9+oT40aMLAumMYre9LK6kjd0s++hX3lmrFupJklaOsjjEegD2
WUTBfo+H94bMoCvJUU0d7VwD5eraF2vesjPMpAa0kU/Bl2S7xLxNm7JhWjar5cRi+4BjkHSm8DYk
/MDtYj15+6As9Vs4zsASnyb+2FvHRDe09seIAMN8gfhJD8I0W50bCQDpBJ+cQwig5IaoDXdEgaSe
wAeYzhNAV1eGNDRmR95Ew8EKZt/tTs+3gAS5RhdwGOyDe7Uk9jyTqW56/SiV2sQHh3hjweJMHYQd
1YK8RJylV4qk72qtC58bxxi5naf/2+HGO7rQbXql9AD5Cri2czc2d1Zt9Kg7FZDPmx/6eyhHVu6v
IMJpsvnDuYe5k5ajVcEUPic9JX6iEeUiAsaskFSewOVTROdjQErbXb5b+r8PKdfKVYVyTvmV5scl
kszJkIv3C6jkzZr5uW5vie4C5h0dxd3Izqb9se2qwe9FC3e4g7TbgjzB55Ae/8/3QleuQKs7u5a9
/erqthz8aRUvb236aXy7406OxK99d4vhIWS34Aw1Wroifn8mbEwrSDjr73o+NN/OBBPLyxT+HiBC
lb9dJH9dW+qxdbQG9AZtahEXhNQ0t1tWhSjjR1SM5q/+M1+3kWAnwzkNH5AxM772rXYrWmejk5PP
1fxnpL8tWFs97BEqwyGQDStos/mWQ5VbewPEq1gceqMyUz/vLKS+wC7XVVi7ciCInbf05Ey/g1/o
hP9iLmoChMoRxgm7c6WvekXjptcq7MTQkqbB0ys+NHoL/FGkHOxaCdWLMqKjYuwq3p63DPCe7Msq
0MDtdr6Sl5RbuYC2rYF7ZbiKExVtVXRF3Is5c+u4dGDWPYefSDdrvJeWsSm5Wuq6cpSGToLKZD/z
CMS6aRNtZcRGB+5VBzu1jIgxvRxBkr4AhwHzc7dKRJOQ//szuXcs3vUUIIm+FY/nL1VEC5XJOVbm
XASpdafL3I6R9cShe8U9uUPSl6+u2YbZgnVCHHYTtEAWI2WkvGJtyk/G6W7/CSAa5m6wwX5D2eXm
jv9esoW2XPGt2ANJ8AVMcN55ztoxbyhahNkAWEzA1tkfJEbE9eG8wIO+eZfLWIEoH8lwlVFH/0mb
Vn2GVTlsvHfEzyROarUTt4ynV9GghQaON0S4fwRevGNtiAVtJP9nN8bfFtM1V3mgXZcepNBsbTGi
EyOSLRZzGFFYCB/j808xIlU4jXV5QHlP7DoXuxUN+/wmec5E/HMeeOjqgAS0NYs6GpVbKCVNLxno
igXWs/MHhFcWBeok8LyF+tHtwn9B43uFm2gl9Ct0ufz7xK4M18mrvh2f5cFvxt4k2VRH0v1hosEB
K3LCtXKOviiIxdpbTc0cTXnT+x5uQGFEjJnPl8Uyu4pNaYjhvS4KneIsb4NLJtQoJkm0kVEwgebo
eG0w8jGxVVVdVqLZf+1CYA+ca9X+HGsSP0d4bNlWRtJz3gR/WhUpZ2MTghOyOV3RNkPC7C1k2lPR
FmWVnkg+iixrOf5iIPBkLzy7nK9WeTiEs9LSgb7Dzm5MtYE7ZHea2jDcHf6SGBQs9giBhdwaZpE3
VGxKjGBj5RLok6xWVk2+B5Z9Mv6GO/F0E/kzxUkUoxxriJ9eqOVAv52jB/bqzQSZzCcp6I0IW3pa
9waaX3sQmbZ+LH7ErQWkdf2yNKhYxzyoEYQaehj6NuwA+irfMwKEQgpf3ru8jaB19R81Jl+u4892
3s0oMw7R6Yb2ZJjQXhGjV9hK/09ugKEoqWMmCRx5VYkdldo+8RNR0lz2oVSjHQDraN9K841142E8
lRhniKFqg6ah+hIQ5SY/N/Y3Joj1fwXWfxbhoRig3z+Fgu1nH+UC5Hhzjuhq8fM16NefMcfIeaJI
OMnF9F1xrHq4Sohp0GO7L440HCP0SnzuCuxEPdWndUfo5segJxp+4GrKhQzdEn25P/gtRtGERY2X
OCGacplW2to+xC35gwWgPA4fWXj0C4XkLl8ZhZsijQRb63mMrsCJNjrB3FIYEtjPPuAdtow7GDal
ku6QsMHMsTnhyiEpbbSFc4c/CE1iJegOIS/Ffk8FD73g/KSPOQOmP3yUyGe8MWAnlNEkscMTryNb
+UnT0IrKrxJ96B30pkjm3RftIFoBToyfY2OAsvbZUFVjlkKoPsmxbJPMMM2ydFvWRuNRCeg2czrO
Ob4S22zeoP6s2vnx2M7Blj0BaSPSeJOWuEw2ipAlMikHRmrLAb/86C4HHtfadLBDHj+XsaWAIr6/
l6lEtLGoa7XxhvXoKYaRVai9c5MPao+xm+cyEOeBwwf1o7G0s9+x/+tE7nS0ncdSitfC3/Y4g0EG
1Dox+Gzcuq4aKUx0u04Nxfae2mZogLrDp2ffWt6+N3i9cNkEkFTAseCYvIb4dybzgBWQwDKXVvh1
TkP2qCrnQg80TnL94GmB3zPf6oFgIAcwtmAPFrznTfCagZBJIJ0u24+vo43dMXA8CZWK8mDk25AI
aRIN0gLapGPOsdMvhijAaSc8i0PJc7TRNcQGlkM96Sicq14hfKwCX0QhkCWPg4kAeQ66rODf4oso
3aUU7wuz152gyy60WHwQXBVln+NCO7+Tc3mEenU07a4bq5/3CQdA+JyK3MEfKx7Uude7CV/pn4ll
2VQNzJFZV5TDjAhEiEhfK+kQdZPbxA075bVR3uCIx9weVlCFsR7hsrA5/00rCmr7Oix6V6H0xt4L
Rw8/rGD173XqL07oJVI5M/OIPF7fdJmKHT8sPhY1TSMpxnZ7bOvaMGBGxzZ+LsGR5msWptTEM/wX
I9T7Ek1MzRlA24q4VryerVKgMg07JtWFoz7xyOyjdNwwWbfSN7fd1hP3K/qz2WiUc2e1Lcqzg/vI
eWbvP/ZrNcchHmSLmPI0No1bcP1VYzr52KyA/+opW/t6yz9gDbtLXDOulTDs1v71kH5JL67Tl5MV
8FQw1ypqtGds60eF2HQEOhzJ582zaLxHccB/TiPTlpSK9rKGxZLNJNLcJiHClcMNFKTqM4HXES7+
okRRMEmy8pd0UbzUxeg+X5gW9rrfaIk4+VRxOFzF+AjxVudOiUUSDQNaF9HBmwo980tbdr5YowxQ
EiWvujuDZQplfNY4gZx0sFyX/OG5vvxSOfBcbTk0LDMs9fBHxyM272VX8lvt2GCJK3QzDVZ48FI4
qiXgH7VSApOm5XOSxqF5oycWNNXCa1cuW0gLJFyV0YTCYmWpfJA2hEgJnmFJ7cI6d2zeARor4PgW
/YyF9T2zNUQIx6BKNdcQvIWPqsdphEc752IQtT77GdGn+AEu9GBAr46/nZh/7OKvJczcsXoJ5RSi
bIiEiZKMrFli8CSeLke7xt7SoxiNEfDQWsnXAYC9+Hur+JwamBiv3YmI9Z2iN49ELW3848EggZCx
HF4tVSb5toIFiD7EGDYMjtwJy2mT1RNluqVPxKqvQnbIn5FiwslgOoYZE2wZrbfZlUZxhYhX0+mi
guu91eT89W6eh7UXGHJTJu01CMC4g7nfTgGkxxxhA8yB7eDQz6Oa1ORIrkTQDy0qxj4bZq2fWU3K
BZuSqgWX0jrWRnk9QAI/1E8XnHfOxANT9eMQzMV916aO4V/EYiC5QRHHR/NK8nlfqQDaCTsN4uR0
84vlDgGQ9pLrIgZtYigMl9+8qTmfuph4uh0Xp0n6d+ZnFR2mZcg1ZW8NVypqLTHn7i3IushpDTvk
XUEPvAsJzix253Lm62n48kiYn2w8BfWY0Wd0ILF/2QbgUm0SJdUFl1F6Rju/SsMxNyTlyItRT9VI
0GxNNV5ouXgZxtanDrXIJ41CGoAs6GEERByCY2Mj3zXo8StQIlzFG/Imdubyvyu0heJJ9Q9LkKkI
DW5gykaKm4OmjVLvPUCk3rwCLRC2KB5Wi0yde8GKorhQbkh1OU8hOwCPQQ/3UL4CEi8otsiUQFOI
Q3XTGPw8pfSnXgaryOGSTAx4VQJ7ATJWXQ06w8hImRGC8jxxRO2eUWC17ezPZB9xu+mjeZ7XeohV
mTchanzN9VmwCLI1yU+dOU7imfD6/0X5w3zbEHUTF14iumkRt/16B8cM2LYn/QWCIyq8N+FbZV1Y
Xe8OppwRgR2F07Nv4HP69jOP+wDhCR/OKHOW64asYZXbYUX/SQqwdqIO+1kQdy8o1c+Wo6JsYmgQ
RbBoLy/OiCA/cEtdEk/94IjqOqcp5YMfPtHYq8RopsowwtLN1NfCHWNNJk7GfG+Rtg/UmvPWliYz
EmbvtMmewN8PG36FNJr3lA8T2mOfXi3vlky/IEzzROtF0IyL9p+Su4UW25SuYjR6IPirvThpvPqS
DuGsRn2ieRB6Dy9CuXK7l40qtuJzbnh5cbDwCcv0mkCIOf4WfzHuu8osJ53AcNeLfUqLTdUvtSDh
FeK9FeNNV+y3ev423neU5R/bbZrt82dGTUdlyW/XGN54p46pX51IDaHOJRnd6677IGaY6SBa/b6e
WG++5PI1RYCCIOD3+rWJcOSGD7GTwMxyi1AsndztGb4Z0YYIIdqaELzstM3nMfsXmmvAGb+mQuTn
MJzWutmTh70zmRhL9LqdmhLYZNw3ZSDSM8n+RxH/mkcLPPXqKM/Q9QBiS4K5Ot5nLG8zpKg94/x+
aa7D47Pxzt16eXRQA4f9iecu8xpiPN+xw4oZdxIXapVqsbfKweTFuYxSDotHxFdfdEN+JlulETOx
Hb4Q9ftv7nkU+ShHr4AshZ9mUxr6TEr2Y0mQzts1Zw8N453xvePDXI4yq+I1/rpNTHM6pZC3F+PM
G3yZJmrdt5HecwBsGqpNcScq3saWRYnhWsugzJaqJ+p02kNoAdCxjqQcveus1e6F5S9SCwgnLRrs
0XMcj+PwWh1aHfOitp3xzEn9KCDnFRPUXSFAccsKyQY4ISgBY4GJyALtCS4n2GPO27sHxAX3TL2M
joBRKpVOwkSaOugceONWjhS8Ce9vYbMS4LhjwRXbEsCx0HWZzcBpZOwRvRuACZRZJejKBJZKmE12
TnGjH53w68iJPDFFtQuB0gMF5JEjaIMBdSzkEt5VZm6n6aHmhm6gQUFkEtTc5KL20leJNb3GbYYk
sbYDJlRUbofIkraijZweZBpj7bzr1cuOBXMUo5Jfnd6Yqw81o5VNKRXVg1+xDeMDqylJ1xStmqK+
UOJkWMd032krEg56waTVSelVE5mfLKghfpQQfSDWkzovls8iRvfOdug+YKsi78tcXWDmtO9cTRjo
GVcNLAnPIxjkAC4JUgVa097k4nPVTp9xStPfxZIhdzDfN01OMt6zFeh5blELId9JS9CabAkSdSWb
ROP+UtFq8UYsfPHbGvkmOhF3fvh9vbIQ3rk9kJMLqqxHKYwdtK5klV8TTcjNRCWO50K8rV0G4qBE
uwuJRABG2/l8Spgo0dSQIqPhADe2ycGChbZeOGiKgzvkVOZtLdtB2BTaD3Nd2oTiSKrFgZ/qHYBt
F3fqnuIe0CrU311ftD/QwJcSIUhzjK0Lp7j7hUIr6Usnn8XloPXcDQmwqht1O5WHu4c2sboMupCu
4gU7pVDD5EzdYnGAS3VjT3fydysX7z0tp8e5oLpU+ID/R1nXNy1COmhzNrB0U2mIQhlbgi51TW0J
rziD/E/WX3EBGp/+ptreap/j/S03PO+KVkNn+BSEb4YNsw0WMMQ4N6b0J0kjK+R1qHRevqF9n5DQ
5M4uZVbJktG7aGYKASSr1m0e4nA5p0UzkNTPFGUDtUUO0ENx+uVhjdj3JSNnkK5jprN8j+ORj2tM
fhoyVTBuHQa0y5jI9GLWsezPv2bpUjSsYy0614NR5ZXLlK2sYLAwWHZhJtUmlqJg22B5miMGoH0u
3mFQjoZh226nOflmQUO1cWMaqeXXbZzxj+gAGNc4hdUwPABVSEwHIsiU3l2GrNwVA5VLseGT4a6C
L96unWup68Cduj+d4FAMn+OUyJ4KN3j11lDI8CxCX11ehIZrU1e60saD4Zyvrr1KlrV2nQXLXJSJ
YYf8oQeVF5/VmISWtoawS6mzcIFVN3ja0+7fJ3XmwIqA3h9hpgaV5BSEY53vhhIDfrzavOntO6Bu
pak8bMKdxY2X3qzuMfgZpS7UZUS14YTwuj+jjBI3qgu/7YvGPDqr55ee+HcaMkLQUG0f5Ige2hdk
ALQEhxSFJM3Kem2LSLLoNDspn6ie3EVyvYnpz547XI/fYJgBdAgqEUP8S+TdewJbwBRalc/s+Xcx
RW9RrEoYmW94O3J+O9q/9l2SIXwNe8W8NUK62Uy+o8SBFrH/PSNRf8c8ky061N00vSA9PBGDkrLx
rgdENJdo4nxSdBk8h86fkKuKEBZ/aoC4mVv5G6KWeoEMlSt4000XGiBMFU3mNfeSO8SMUq8WK1er
XOjoaz8A92tPql20KX5sscVUIufYqlMBJQzdsg6gv9zsP7upVBI/bnRoq8v3ipziejbPlxBkTZB7
I2ht1se+9dK3ura0yY8QHGa4AoLxxmsERIXBtcRIdV0UTjN5RkbgRI20tOyujQNfvQPLYQQvO4OT
zkw3edpPzGyQFqPREJ8tS9QJHY77e5Cr1tRpJ66XsiHN2IoCgdfBuNOPzeN9sZ4cxuPicDxQor6F
4c+fFtuEP5GErridbAmjOZnQ38kSGjy9510bWeBb3Zhyuy9SEHAxzVOiGMViwC1KkZ7fqQd62PDp
p8KDgoUUXZUG1y0gME124iMDVs/9Z4Mefkjr/s6wFSaoKI6VHnlV23IlU6IPlRcQbXd+qeyPm1kl
s1oX3AmrhuESXQXXw621wG16vhsFE3aVGucflZhNM6UdAYdlsgaCSJPn9Omogd3EmwJVIioC4cxa
OdYdni93RSGkG4Lu4hKfePWbe3b3WZ9VF4pYCX0L/Dk84n2kZ+31d5iEvf6FtzwAd8gxsGTKFmMa
XQJI8b3hIS0pbD7/SPmWuOKZ/4Vpp1VfTGQG0JcXZq6u/amZFFR37L5FyNau7umDK0mKyasBUurk
3ohpLpvlGQj5MPWJMo3LMpexqgI/nL39jmGXmjw8FUQnXrZFN8PdZXBZZnNa1Rlw2dNC2maB6JIy
YSeB3Y/Zv9UIitD3n6ERPE6wP5jotXEW3GAvf7n959OtLicBanUcm/buwiU9oOPSVpELmPaHoZ0T
nomuvrHHTMRmfdYypkk69Tf+WBXwAQpNvPkGfNzFPWSHLSwwhB0q3xwF14U48SpWJQyNYiba/F9H
ZdvdGcMegXB+JfYoG4yWGeL5KBNQ8N9rbR9EmTQBCXn8IuPWpUgV0iZwLd7otdL0OnQ4UGdu5mDg
tr2PuFf6QUCAqSYyBxETgKUtKh1IqKWPqc7LIx776ckKo9FeN1k4tKzlnCg6T2uVN6IhMwBM6Qqk
mq+h8iU8+Ax7Nwwdl88R/ckV2Q7f1WumP7RkbYew+tGO8Izz/9CYe3+wgwBgAYObbp44CLkd9jmw
rvcV9c0S7B70OUisAHXHzmwaPMmCVTx48DuH6JfVISUk+beojCLCKnfzqKlRLSZvS+dZY/vnnVd9
9bIByI2sDND/LRSx1xhOgH/UIPs7xUYWiyAN4a9Sam6Z85vDH1z7RYlE053HVoFwss6uLOwIj7TM
h3bBvJ67Ht4xbgTj/emxftUAlKzkK3mYgrY9xBkTensaQ9vpLiee5HbspdupHffDz2BLoftJBrvw
bZL5Yz1QJwCW5I26Y/3igIAySFN254aNc9UYYVv42R0BwdVLVuNHj4sQzzuW3Qoo7wls/E0Sg5K1
zR1gwUeYFvulc8ahsBkMmqdQfTyaAuHRYWWMjzoniinlD5v5Z21qo0GHlUc7BVNqMgm1q7Gh1ZvN
75mekzT18FsF8B86KbPwf0q+uxSSDfR9E2tbSye03H2g/YPu2QQ4dPGkzcO4q9VmxrlkVtUkkAKv
4b6HBndkSlvavHsaIFGMjoG7Uimaexo9wyNi0DqLBwzxWJhAdNzVAKfElaiBfXoRqY8oOAXThXAi
wPq+S2IXaIPg/uwBPehcsfiHWee6iobPQSFkpPFp7fsXbdurGya9KKIauw5N2qqpvQygEsigdnk/
Ld1g11fLzNAvLZGLDdtlyRolAwkUqgBrMUwpH3dXXo1sQ/HzeJGM4B/A5b4ci8sjVdlb4w/ZEavB
Hwdv9dENcT9M9+wsqS2qbE324UouulvItl4fmxGK5XlaikGF3ENBcFO1S2hujz2lYMhR23+g8Fnj
Xl7POIvi7HHFog1U6IeXf86txHlJ9NasUxR4JYH+Y8jL/PqXBn4PWc9hcLwIXvzKh0W/ki4mGpq/
NCC1Cb/kRfYuXm+CaRYrLv3AACR47ptIsLu8r6pWx6wry8DUOc/Y2sF2+13PhyBpC9SInNp5ip9d
Si3NSmD89kGrlgivADPT47zNX+cLv3eatUQlzLgZZ7UfAoMyzcW0zCXR+e/r7/f7q9gY4Q8uRmlF
UCr8RJ26RG9oncoTCazGLsxHoQfEkSFIEyFDsQaj9n+hq5Sf1Bh5hyhqS2CgOQ8O5w3ELDPfnD8M
c8DA9mAw6rbqt6xoltjuRGe1XEIo+F/lRg1TDQePsrKqJb1WvpZDsrmWc9fz4YlaMt63vLgdZZSB
sx7ZfdP0fHgY/a2+RnGaeXDsKHo5F/IuLHRdUL8Tlcv5rv61eKqowRrasDIU6828Pfu+aKXtBIfk
Ur/NqGhIjhDIukUZgf97UFK68ljgzt/SP1WEWCHA9lsedIdHEaf6rt1m4UHE4cCWSf5FgktTC5PZ
oBFFNrX6gONZBnkQV884/AMI/RVKJb1QMmv3thCU+zHfzTcwZgvdfhoUr8VtUe5HTfOAdSgEmyaC
4fOtmj3F2aZL2gLrtRWByrQ/3R20Ufhczs77Lu0d78M0KIJSfJmo9FwHCfsrhPDaaZxeC2EZK13Q
4dxnU/5iX85MZHg6LW+qJXQ1q4NY/RZQFcW4LyCs5lK4/t811onEmKlIQqk3PAKlil71P4xYXOpo
NLq9z6Hogfrwmi/c1gJDl4hCWB4QUlzkWlOcOxPbvzHT0Ndk5cOqZ3SgDFAmTR0ZJKbj4+gUI4d3
AggmDalgQh385Cp1XJqIK+s7RpwGN53htP0FqFZKvhyHqB3b/nrmYF+SC5MSS1b6TIaQHSELIx01
JZF6Xkl11DM6w6tM7ysVkGk/irzdyNKpD31BKj0qmtxpuXt88/ZeakKcGBQGgeBpYp989TJbCir0
bedvcPV0NGFHQm6lH5GBGGSOy7ix+OyIa20ncVz7BC277vj8cKM7x/YvotmfAuNWDieXYaMZ96/O
lzsG0j5b+pWA6+WHQvKO9U6I8EgWCwtuGgD7gAxKgTzjpJdejMCmMKbgHBq0A+7buuq6iQeSw5jy
trNUrLRLlsOeLdq3fYuGFWm5tMsbl5jOKs4v4HE3fhiLSDCEeYuLxeB5TEg+6s++S8+Zfyj5ywSX
Ktn9ikmjHyaufRWnAKZA7uxfXsuTKwySmVHqNlwCL2A3tvl664cM7O+X/xr96Heasyi9H3Ea6vlc
ylHnkj3DceoJmCQN3tdJwLM4vklM7v46AqVM/bxahdf9sdIBVJimqONbKqIscNrh+HrEJzXO8fco
+FjPGnYbZH2WFocVDvHkn+315ACR+k/QOBL7id1edq/676Ha31R/5kZf07YKV0pyLu1H/FnM2TKr
mXwykppnwKTNeKpp1LEpBDVdaWesJQtUGzR+/Jkw66ZMVJa9VTn7KOsXz6gW8hNQhhIsFqEC3HKj
tMLCm/TDvvVa/7o59DhlJIyX22zNrXp4YnOH2ftmyUodYaVReyN2RV7RHNgTFjBRuCdEUyvwdYL8
PWaS44q4skApD/Lth5bNathOLfLjcoMUY1Fa90uOUShvIA1oYOLEGdwiwdmBzCjQtZZJALZ7/Hi0
iom3iAfq9JGuJgMIuH1FGUmsjLECHkUqmIO1uhGb1rPq53b1zovbyBeaef3gmAfC9Edxe3+6tOjU
6SM7vLgN4182lYi8wT99UGjXIB3+j8mQpbls1pGBfeRU5RHXlhCZfhpxS0eCQXOOIE2RPIwxCkfl
AebASnIUNZFk1OvNDH2zEpAryxmbJamo9iEfnxvCSwLXVmjR8wI1Ti9ycARp/BbvhKB5+mW+QYpU
I9KqctjxYUy0LwEJZxcu8iBnVx7bjPkp8afY27v+zaBJRgLUQpw3Z1WwpexzN/eg6iZUraQ2SDSB
AjQrzrygsg7LLV/ISykj9c1+1nCNdmA3WtnZkBgZz7NU0VtCSZJB0Pbg4frSAjb+ukGH4EcSAb3O
VYLYPZ0p9qeqp8/7fJkZgsMtZZpmxylQ5kiw6AnqFVZD24fhNT4pdOYRVD0XGk5n9WIan7zNHaKA
LbSo388TV9yDhprIDCbiNfG+YcA253KnPxEVkNy1dq6qINFwWhEs8pgNAq8wl1S4kaC2ZFKWzJTW
onQbMIr9rsRYaYhWuMsg2fiymrQG+abpKT3hocThDIQU76A/k5NHUdhAt8zztP5zuVw/xDPTuehp
K5664O1X0rGdMqfW0x64mwhTzFamRm8tWORpLxACnXoanQzZIjKGrsOaZGEkNkZzvTS7ZAxicXDP
aWsYHH7nHlziJCBDw6dLOqhNhsWdxh8OTl/rnBOnE200YukPqb2yDoF1x7jDNQYB+d0g9Oqft3Av
x0kMl0rDKfGR6vsVTNFR0VUeC9PD/4mdBX08mS2XOFGRIYrGHYMZ7mIOmGy+90epuS13RDkq+zys
GeM2bG8QwPCanL5vIDMbevWkQoTYI2DIMS9++yjJ8gXyUVD3KwVisn8x7joChn2NBtVit5fqkGPh
hyt0GHtF4IlB3v+EoJLsm/IsbU8Ntbl56XxPvcZkxeiGIj0Ucqim8f36EdRr0fYbPY6TEJVqR0I8
0fuYaYHEGQeQf7tr16N8q6yxXR7YYF23a3EuCk63dl/JUtALAMVnfDKj46WZAdEWDDHBcRTZ8URl
kd9SDaL89FbmnRKQY0OJSAKjqtadkUVDmILuDtl6H+ndvXKGE2Nj9DcC+TGNCHRyJejFYtBmUtXN
5ujLFSoG1zsE+DW06Ff0cBvk0VNHCAhZ0OAcfyTd9NvjlzOQZbJF81qxfXO1lJWJN+hfQJ9ClW4A
DJp935rpntLpbmk4uh5tyyq2r3z9QMfrsHeOhfUUxhUGLDs1+dRcV28vgewQFTbu5q/tIHaFk+kY
aLXyJqRp/j4oZ+UXifU1nhMtSA/xqKENeMpwE34I81/SaHy1bkW+0M9vf80ASagNTyy5Ch4vbojY
yAPFAIV5CLXhJtrNOEew2PEU3JXbIcAR2nDglKSoU0JLhRX+CF8SgNwCDH11D3GF2jsN1Z5jK89U
wlDoVwWpZtwQqPb/wEaKA284bWB0jaROGWo+s8LR3zNFeazq6iSoXysSJ8t6R4vWXqN/3zOOY9B9
usyrKoSFbng9IsK1U2CQlNW5EksyFdJD+c9yo6xlYweCFx6qqwzHsd7iJzQjSOeP8BKzwjU/GFU5
FiRDS2fELWymKvMzD+OeI5QW2ssi0jMMNKz7PSqFEWx+BYfwakGx6QCeTBneuGs7rs2y2M54TAC6
GEspTimXoKuo7kSSurRB47sHjlVdyrwAT5sbdqtveJaJeek+8OP73tRwPOudAWsgTHGs6wAoCWhp
ENIIm/rT8MV7iaUVj1i9Z6/U5Rtx6HPcrC48gbe6Wp/3ML+XsNa6XFVJmwLK6oqnOm7WWHCk8rwD
QUgLeB9fcbpEQzwVxOt8VuNvyiWti6/CZP+eWpl/PyIuKl7Icsysnpqlj61cKTS6EBxNSQW/d6Q9
JpWEQti+VYix6kE5eKA8o7h2u92yN2Mqnt1YhCjfqRBWaRhR9UJ0anuthadC7lpJXquCy1nu5m2Z
cWe6++ESC4LxGxphC2Wqk902fG/n6B4Ks+A25i5BilCTOYTGuHeiPWYtJHLcf7uP+o32oxwToRD6
710koqa/r76kbYJRF0pnoR5w7CJkU3TFH8dJzFXKkt+sd/T/pQXBVEjlEUcOBKcondR8bl6539we
rTCwwGBjW5KesiKVvAySBeHKGrasw8+2DTQnRJCZw/qU4yxMKEqNjRskD/qkVqg5Cxm/wOeQNhXw
bc5WcxVL7GPE+bwanS+EJ4F8v9t3hiRnRXZgB864DMBwgVKx7CPVL1lFWP/TC6m8BGMC7zfxJy86
nUiiRyT2DTNN05BBO+BepcqTmQLGo9Gih3SatxFS/paF7gc7b5o7sYzgr7MRNSF/yT3ktZIipfbd
j4H8SV0+zbaTf6a0NpGWzwDofI+FqyLnz0fL66HS0D+fo+cpsU1c9cvGIKzpjRB6h/COff3edfN6
YdXd1riHYQcavSk8UgErTshAPKR3vTTAW5kO7w0XRpxEMJ3DUSLlQERN6eVg/1TvEIpH/5IgUR2M
2fuqjwVwAmiErz1Pv5TclrDnYE8kHz5kjdIbDszi7OF5WA/efDn41t+J0o/eL4mPhIybFsno36Jx
ptt9t884IwQaZd+M7VEPauWUHKWAzefHibE4d/JIpC804MJaauGkmDoKVcEru4ESdrg9gQZplri6
rofBCkhU41NUhVIpmU/gM0QSSi9z+6RWTouStQeNe18+qph2VqPMCdwApqAoG7m6OEv7cOnqBUCs
BCGQm8A491fljkfEixPbeAltR6cwGnj1JBJyIi4c58ecc2y/vKoM3XnidciRhzaicMyu9l75k2n+
3+a+r4OjOqI6iiDuTV4SSR/WRfm2k19y2XZQVPXIEEtG9a/FRlpBAZU4ZS3ms8QuNwf+8vYEuf+u
3p9nw5EWdVqpkwYpNk78d0nofWzTh4/v6G54cnOK7sZzTaPM83dxuKQH2i2vxXacAsly2HRdfzGo
89SfBj17tUn6Dn1BtkqysxYDv2OAkIhmCWxfbIryZh2YFRg+QDlxdXAUIx1drmACyAfI+4CrK/Jf
DLxRnoNlSJqOZF7sA1zT+AFPHO0HGsY7tULzGCXsi+a7dLNQJ7a6rZ86/9rd3TbvzQWmTFvOuwD5
TllBfZYJ3IPpJSOvDx+ldZmLUrdwqliem3HTlpK7aELW70x6b3v8bwkUEoihPB3gh2rx9CDNbErp
RqF9PRWz1omTrmjmu10V5AagNxqsLuHcXsHOqL/lJhdR3CaoFU5wcG3YjYNqJKv0r+pcuGFBvxRx
1EwAuud3vSmBPfgRg4E3phtQDRuqO0CNQ3/m9hmY9AV7Ub6BLdqdz1qdt/Ml5x0T80InhFtqT0lw
RkfMZjPNfbGmy1f7zdIRgqB5VKtaWtygkA69mpfH2DZvBypWOzHu1j7GdaQItb3LtjFhOjiQ/7NJ
6ZWxtkvdCr8juUVddM1AtESyZRlweFD1IvmcOc6XmDST5QMJzCltoOmq+s4X3zFNKvLTDFA3+uOs
r1Kg2rwcT0BrJiRjNWNxG//VIxHDNXUAMywtTIfRQkU3smhC3goYNqSJy8pd0AyP+n1blaBmjfTD
3jG9HDDUScJL+9ZJNgngLJI4q1wVS8XvDw8kPlrx+eKWRdbTzXClKJv1Q4HhbWZPrLjjSaMbDf/I
DoguxjmWjdF3j6d6kklGnZeVx6WyCGk3XNmKHpplypXiQM3bnTlsc1FNt963YAIqFd1krIogZ41Z
KguyR2TKOJxU39WCo/9coklFVGGMXIWESZ22OsISDYuSl6+4G2cvs6GLjXp+rhWJWODPoeyo/7jK
SfyRViHq+8TQOzoXETYDF0Hl/ciY4P9efC0yO0aYn0JoLlK82TVNybqvNC680pDZCP5dt/tgHiZT
fhr6T3omdlRV1nGXYwAGw5jCbyvezbPNO0epx04LydPg1E5QD5JkeaSN3Zr0QOFaJRFPILz/9Ta8
5/d1LyhJc6MqnEez/y6Q5oJL0H8eDgPiW67yJjxzfI1H9nIsAuAnKfx41ypxesnEnuVCnxfMv94z
1JFyEDgDrOucDZlxpWaieLF7gCd8E7njAdQN4jS9WAPCP7yxaHfoq4F64JhDPhqxWw9cilI2Xod6
SlBzv4F+N1D0Qm8rUM9kKZJT2iS46m/8Ly2vAIaaPZFnx7kdG86MWlx/xNqbhOw8/xxQPLXy2WcQ
XfIfSvqk6QrkVrMLIVQ+8he6pD3+Kdmz9x3fp6Ye2TEsGvjX2fz3rZuFuVsM3f48rJt3+lmMZRcH
nd9Thu+Bxf/B2d1pntK95nW/t2v9eOI3G6QfxUtsnD5kgZWZ0IxdD6HTC4ST1x6atE6hDgcG75zD
OJpY0YQCZbJ69IBRCA+ZgxpB6LSlsbBeBKbsHSSwFzw2gGgkdkZQIHap2vcJhbDHoci8ruxz1uHv
9bYDyjeryD/MYH9Af9k9qpQXZWj6cGFeCwtA56EqR+BEwN1ukpjx2U1ht3lOHfRn9aktooarFUES
WPVxmPm0XZ6M1PgHNUCSSn4zqhNwbqhQgKzVMZXVpbmqpbphR2k/xMGvOV6IfXBE5hdDoNdvv1Ug
nzX0tlcLsTwcwHoEJkXql9c+P3dEsiL8LzLNivQZmq0cCUEQPZ+HlmEKMPCiEgzy69OM3Wu285jG
RF7QGpqB3T2jYwhhJz5UlGKZXbjX0wkFe418ybM5ZvZMWbjroUxgByTbajEtc4dn4y9ZmNcKOXSf
9JU99HHSe0uL+xlkFwdAXk2rLkKyEsgMOqymNcjjN7Qix+aOs77aqDfHFtiDb/9hr5S9j5bC2rX9
qTQ2vqhRsz+Gq9K68Z7rK4hUaEa3TOmqD1WNUPXcUTwhJZknHJFn7g+qQK/2IFm+0g+/VR0c6ygE
fjvd50t+0+Rc7e3b1Esg0j76nLoOSYXC9QbgaYMiqcy0cH6dOEeVKWhPjnI1On8uSWwTkz1wslLY
Si6pMQ1/CEmKpLACpxge/QNaOKk/3YDYc78JsJS/hHT195XkD41RwFEEEp6Bt5D/K9O8UswzfbO+
A1rn0jaItNG6btb7nD3WfSrPaHpoNcxhYaOBnJlbCd/OUst6VzSMbBmKqGQEXQwN/8xW5TLwRuWI
xs+DU8IYtnxbQmMoTHGccLhuYKu5r5U49vC1g3w4XTIaq+NuShpPb3u7KFAZ80nYcIXY9m+YXYHr
ZMcy5tRpj8VVe5bE5P4jzdRlcs8u+EOIhScNz1bWt2BIypyDPyanH3iE05Wj96yAfvBbezlLlFbB
MqYzkCqglQ0Vudtdq+cmhbzflMaA4E0PC2lsM5vZ1q/6DXnTK6b7RcbhHrD3KtYndYcHr+Z7k4+E
DhCk5E05Nh7JYGQre+x/XhyipDumthZ/gSWw7HEREDkQ6yN/Qn+dV8gqWoNCPeruUIuUbgcjOK3V
7UNE5SlV8fidzP/ZEdHLrlEHXCyVtcM6i7pyCnABWot2RAo3+ILGBm35Ti4VJwiNnr4GY4HICGVo
qDMa00EEKCm1eQFefhFKwNqLYgMhuaiszw+YOGkz+UjAxwB8H7pjHfaegkv7xukzDZoSA4w8wm2t
UY34hJZ5MLh8DD+uEnnswAef53fBTf3eBMNoLd4Of8pnlDnxwvyBS6LGyN3fbVUq1ZmOur2mBYR3
Bq2EQJYnlHhngZLaXoOIylko2E1mRr0t8K2KiTbJam5cWxdafa0jEK6oo7ho/6DvHRMk0ag3hxtH
bRHHcvqi/Tkmf3/uYe8adlx91DXRSmxkeW2AnJJkfcRMwF7ksZO3BRFn3UYnUVO9FzkjYOHLUnry
oTORiy160XKcZMFpOMCMoWnEvDMD2co2emWBJQCk70YK++dXqDeuEnlGqzew0ezCEzhpc2SnnL7J
kHbES/rcITLzwZYZ54cvMM+x2oA5BRt/czrIdIQraw2ERJ+JofjJ2km5jrbYclgFCI7JtgpAedZC
h5ZC0PnXrEFd2+xaFu/FyaTcCmjXGsg1Y6oNyTpHJ1seATFMKfulLO3b/ft5Sg+F2fJKZrfxU5wj
QHDpS3ixtF+SjOED4Byzld56dxu3VvWzOrH2NkUA55Dhrutew+D6Epr/Zl0M8523/32+AfcvR/xr
1J/KY1HrMfbMRVZ+vKNssWFIxsOTD9y0CgBvxwmIP3PVvof1nvF0FooEXO5X15OrIRerM+IWBXR1
ZgvovFYc1RrtPo2bm06JlKV6f6bvv7segxAFb9RErGVCnp8m7YQ8hK3KjONyEw1eyTvtmqF4z9mi
RZa1g3y/jjCJAtNzCWzcKeFz6Omwl63YoUPb5eU1qLM1jN/tGgtdsQYF65lPeTxxTJ5l6tqc5B4A
qsvXCsS8kgaKE8ZI5kT86rGAuS9Dj7EfWRiodKfBq4qCqzDGDDEH2CYMU5SkWvkPQ9odazDXQTFX
aEaUFXh7ql336Io4i2rfqmBKZyoyZ3zENMUPg2mfdI1FeMGzJz3BYwyRjX24lEfXArncGfiDgV3m
x2v3wewUQQE41XePqJe+PKlxZliXT/P5OD8Wm3IUWeC2/3RcGulw3DR0KIXKWsX1v5ox4RM5k54G
PnoxzilUfXljkano8UV4cCuaVxXvS5bAC03w9B7fLvrwCrBd5hL0IIA1X9wNFHN4UlEOGlP9Jz7g
gijSrm9jn3b+rWm5q+V42KDYYo3UoSXgvP58q5WRMTGVUPIhT05MHWMyRq9ip8OifHvKVKqmzCNo
tLAp6xwdB/ZfUxNfcbzvWe6hSx0YqBkx95LDMeX6NpLZbuOmEYVQYFiFLIQIr5SbEKJqCYzTSNNt
o8lEJ5/8lrthpy7e5oAtuMCO6YTM8iCDwsdVigaW2sd3D3YdXODuwH2rRUQhHSEZDdGPxzNicofN
atcMtMkHhVLqb1g0yJvuf9A7/HBAQiGIu2IoodJCRiAf+dIjvqQz80W7EEmSSyMap0D5loo/l4K9
Lso5eVI3BrR/6rL00E43MY9M+W0x5s3xuD2ABR26jgVXW/xoXLKOWkKLd9mwDmLWqXkiY7Xy9pqj
X0buo70o42ZbWNbJqcJFRF7sGTfF6Gos1J8u8jO0yZiptbK8T9CNsjA89tA55l/ZstM7tnlMPGqa
3dc8iiGMo5VWRpaDH+XNQWlh6ySoOAyj3ZdGNAJJ6CxbfPb5Fz8OknYKh70sjCNopEKedBkaLTJ4
KJIklLVNBCuOJPeFccr6KXpoM0aMNHGGPWmTsblPtudt7MfJzAGCdnTp7vjrYkNpmeL/rzkiq9gK
VV/k0PK6hYoHvdg3oJZ98SZl+p44NfP1kjgdr8A62pux06+jhPGDnJFy+r93X+t2R63MZRYbceu/
48rRNCcm817HoCLVSzm+3TAk29G4oUI9lKcFnvOiobakK3aVRsgZbhyIXrz8RrDT/w87Vz4e4qwT
jgQoZuCqIEoeAoJ4ZB081A9oFKsW+EEPMwxeQMy0xeR7BaAd+j4nkxJKVMZO83AOLXp/UP4WL1zw
gXPtbg/RKzG93C00cKS1t7ut7u2046+jnsAOtgxuLP7eK6WIUkuldx2aCqPkN84Dw8IkhwCWz6AC
AJAAkNfxIU0bM8EWJ+DYCO22sOuz+qRyOW8UTvrXPNC2NZUWvlx4BClnDfcK+ugktt1QPwMuqi4A
5OIQZx+iGiGp+s4wjL8c/15OOL5j/kARVqNos7T8YGJU7p/sTOxOrPrbobyeCLehbJmxqDD2/5mM
tiPbEYsOuTHzeq8U3mHuIS+Tcb7d7/JWaoUr2hfuSQVW4Z4rElgc2zBe6A2EzNd5nPY+mXlNvOEM
jumRxv+yhyhwItADh0ermkgZs6cNYXPMt3LWa3Du8eor3ywoJP7CWKnzHXfDVxn9ypSsVSmz02sf
KYZLsSqK4EVh4+G6Oic347eRUX92WYCev9xifJZj0CpB3eh94F5YEM/KrFe4huJE8La6+AeEd6Ui
YJuWE8If9R3UXbxOVKGOPIQGlna01nde+1o6C967h6ogosBDyZAVCqHGmILCvX/U0z37SDYIVcsM
yZyC+9u9NzXLVUDHLdIh34Vqg6k0cpBlJw5eyy5NDS9UM2MLD+JGQMFpn8w+JydtZcNIt9D7DWod
zoCwvP7eyqcscGQqxEm9+wbVaaaxMF8Eh6bWbZjefgdTzROshbRFWXkqLIp2CcAikUU7rLKeaxNG
xBmeqvBL4ufOU1MImF53tb3CckoBkRlFO7pkivXIrkn+lT/cWwFmfH9lBi6mtHvrenQXhD9JAEHm
Y8WVmoW5Fphd1FYxAvbZmuMXjZMoSfyBVxCn+Ch2t/380UrR28Kvw5DZzjWP5NJx9Q5GiPxro/9B
Kj6EO/onKsKaRgJmVxrJVv8g2qxID6qkf/FxHbl8HahTvu/VvppK3bfGg0ZG8oQD5Y74BWc9wo6M
yDNgKymDQB5ARQgPJEQuciUATKfbMt6JplhsfMO2LmZo4wfB6FkYJFB68+cQbdze8KLC11p5ZvlW
6p2jG1Hmg/0nT7xt/D7kMtmS1zWCJ2MyePRWLwKiX5L8CXK9HSgmnNowxFil7w92pSQ+qE/RxjZT
NfyYpjOtlWuGXfgul7Vk8BgS75BLNVqgaw9SdTaoODI8KO3tEPJbdCuJh2BKtk7IcrtMrp/i5qh5
RbA4NJ2TNrXPLSwrfzA0nw1xytpa7vwFztoKJD6Jxz81miHf81eFP4JkHdaqtobTsd/eMpJ0XQv2
iaK5HqHIvPnsd4b8hwghGw37fUjm2PFQucVYVNYrORjOY5c8HfAcpq88W65usqnmWjRGjvawjUg2
7t9QmWa7RKkFHkSWxRC3jpTPQms9kOSdmACBSjKSDyMQZsztp5tCu1Fj0GnOGjeM9Gzw+hbrcYXl
kfuYfP7Y0FD/Al3T+n2QtVnxDJ+4I5zoe+ohTrbFZRc59qa+ns9KMvFD8C+8AYp12Z8N5swqB00t
kxkZV41jWfv6TMihn/6mjcO4eCNzH+eywQkc9c/cUVFU0CoseAWH+DFqL+FkF4PozeUlxJPboyWv
pkunXu/OoF0LXgk7YBO+FaW/rNflyDPTb6FiB7f+DkmO+IZXeNdkx17pAsIQldhS832KcMFqdoD8
VmpUGeTWyktkl5XWpmPIqrbx9elQHWtUfqOgY/7RV2PINBZlJvUvVo/wFDOlh6CdggiOlM1TsXxY
HS2vvkR/c/VUEbH/P5GRLZTv6Ugs4PK9wlGcLbDts4f7XRs6ujEZpvPAJYUpNkgjNfOygQ4CVu4D
UK8bhR9zjjBLZywBQTGxUGJcMM1x9wO9LNlXk9Tk+vCw/HFIVxqIPwEbo70bXJ4/oKVVq24zwgcL
ppSX7b21+jsV5/D3+B8C09D8giOW/NR/MHyrZZHxVPM/FYdzkGxWEKmfy3w8Vettje1s6ipQ4FLw
4R5jXMOq1SJ34JUSwt2jg/4YVfCWHWzg1bZ4EjXs3C8B95WLM1t1WRFTkCFZ5NWVIwE5sIJ+KhAG
wFTGCAEWvzaKP5UMoCjWfZG2DpxDORfKRIx7G4304In6M302OXLyh7206O+0UrWjE3g/Rpb6AaFV
IZnxLe48Zriw+jYrSupjn2q49goV2ymzE6Nzh0i9KF54un4Mq8UgUJs8Fib4lLXtcCiiJ0/gSdjj
/wOCfAHIHQdkD4DHx+AOSCd8MLEPJQtGPs60CCFEOfQnC+DbOrTDs4lvmrjWJvaC9u2XLCOQ9k6W
LVlGLQF1ve5tyUHbEJSJlfIEbEiFbU9dHckV1pooMcrxQD8vD1+JEmc4u01/mDKyY4NWqtHCJhla
jcF8UrjwDVxLICA857x7bguUFqmBgRrebaBCCMtslHR/5bPYsiG90XIf35BebvGXOmsf7PW7HTtj
bWT3iGNu7la7yANSLOR8iAoHuKomsE6iWe5iAtDhyPgql0gOGFlYBfQNtw6sx8EUJf2i3OYoFQN9
qBnCxrMeWnIEMe8qUZ1CsBMeWHpxLGa/MMZSDP1DtFhzVtatY0CRi4pN+/vP+AKsmp99rwoBRVBN
DL8oAKB0di4RJlDVM+ElYPA2OlLlq1h+Y5kREXnfxLWviItG5cFaDJIyqe1nJ0vCxEPDzqC14cZS
A3weD5V/vK5MHXPyUPY0nbPcQvSlPjji9RHf/X+zgsdNCmwN4jn+RmDDErvIwUEA5/eqvXW+QmuB
F83GmgMznXlWucL/FXhlRqP6XkT24KhfNpk8KpZ1TFK//SNlq5EVs+ox8dXWIxIVXQfgsTq7oJ62
K+wXiTuom7HmN28tSIdNwpG0K3R7GxnfAJCCP4tCd7sCws6K0Am+s0yAU0Ovo8SZWnyGQyFw/wE3
nt1vc7pJzvuGo2dceop+hZISMvx0aZ881DwElTlRiA+RWTsWjvuvmz0RVI3IObp5v3nV8sIRx5ad
TYom4KYqx8f7MqwopTQ2Gm4DELhmFqYnvGg+fgfDEkAhIjE2qTUJTj66hgLAOo6LBHwtp2LinM+n
B2zzoV9NBJgeMBkLguKV0QMBEwmH5qx/p+mTqGRQL6aYbi2hdUmDlN3ldVf1PwYTQw7hHypwtF0J
V9I/dovXKMOyBsjwnc79+veFEu5qDRKnsICKnIvQg5rmRs9Iq7OQ0tn+QZOuTTjGkkkp4OIw72sY
E4m81EnzvWQlerQjc3Hugg3k6YFz7I8nDkCuctebfO/iXw+noG6efWuyRDNwSCxsTMai2z+AHWHG
Idz5GdGIZhWjfx5+AOHPlAq01C68it+u/RggEJSwozvXhRHzT71DOgH6ZYoIOdCvKWc2p8BjS0Ky
/rw2h9AFCNebEmjYSnyL1Qm5kyWrO1ZpUZ94y93RUCuScOnIEGFRtsy0YBVJ2DrXOSR2Pp73r3OJ
pzUL2Lc8G6nYjoL8f5PPQtBdqhJ71zBEzcJ0MyLL6u726VaE8ZKhYZk8vL+yfs7i+/W3MVMXJLhs
H+khk6BakvjU2aoIXEm/1lWrv0kiU/7QhNfw8M9B3YCwkDhfwUw6Ey+4f/mnq7us03mGWNR2rIX7
9VP9jAIgjbmL+H6zY/HvfhiTREHq5Oel+mnZr8FzzaF1l3C6BMQz7jIL+JVBEa3afemEcsxFB8hR
6IJ+ronMsN2kqiEkFDmZ5dXDEE2pH9cts/Zx/VRUkryf7Iqz5fk4QDlHe0Ym0UCFPfr2KK+5Ywz2
yO3WZ3BitQViNsHSLKQTppDCUR97rZ4El0GyquM9B7jW1PHyQ5/ZyyBxVW2h3x3EaKzISVlmP+Te
lgCd36tHNq8rmLp23W1JfzD+hp+hz8PewIiI+F5Lp0FM212Hk2kTeTfPNu6clXuMDeeN/WRQ2ibW
RCKrFWRfnK5KDP4cchxSRsI7aput3hxFz2F6LBT/e1l5cyznqq0kWKQoWkk9seI7UTVuVZVaYQKW
00ETwuz/LoYbsI2KJWHGSeGMPDy14JdGTGrpNrbgKxxWrGDRHg+T3rDdtYqAbdJNFS0oaGDER5+Y
5lD1QZcKafeuZHOjUKtSR7r9MVu+gZw8tOYwqSMDpqVC6aVytBEwDhwp+A2WmFVcN/wugBtpIadH
kCYtkxTzdt6CGdrAjT163AxU59nhkGBqf2KOmQ5XUxmR4iqrcsONiRZHAyVE/2uFkyAgTQ+WPogF
WjU4m0Zg+9IDFkxfG1a1jZhj30ar9HU0acPzQ+aRb3nlM/jSPLWL2BlZyvwWCUIwRGqR/DW1odlW
v9VnL4LiId95CwT8s2soBUU4egGZ526fFjLmYXpBXfRDbCHbgMSuj898vdaSa7SCnam6vn2acqM1
82gwD4G/t0c50iA2xwRwVrzbSik0tX79dVw4ENXDewPWzetxu4y6Tytz18WcAIPfwhO+bc4ch+Dl
ZpnXDIQOKGUa5MlXQa1FDxCKiX/sSby3clczI74//TCsKMVJIc+mjuLRPuntr65DKgAa7+DpHMBA
PBjrzw77mitbw0LaJbycskw92iA5HOgLPoJsqYIr1p2gvBohxUeAnvrKtPzZEowQ7qwLyguE8g3z
k0VorQ4zUkgfOZJ5nsUBMdDkmNjLuCxj0qg9LxLP67mUz42FRrBJdyxC2Cys4kHsQZfagkCbpXAO
p8p1mMXiwWmH99U4oMsVM6Oug03l/IIIVeZqInzvDmrPMiDr/muCtof3WStywd0ds6rkQXf181Fj
/PKbftF3Gt4n/jTJH4QCSsyIxu29riPrO12xjIg/j28bO+ppcX4fAEbz7zrvFlV7tkokI2qYd/Bb
jSTdixvx1e1NziGk29+bkd+SaGcMHvpjzbQh1SewshZf0sfIN1wWsDpgjgYCOCkUVGRJ7jYprf00
Lnxfx77czqbJ9jZ9UB+CvHjjcK1TcpCFqvLF63E3ZBddI/AysLkdVI8cOC91KRqW8QGS2mjf0eg5
2vjc9d86Fq3in8IxIDmUsyYtXwCznHppHdmdoti8RmK1fQw/eUJPz/WCQK83qDlw9lw42zqcnzrf
Ox820LVtmtr8BYkmIlugq5b/HX0n4Vvoxijpjq7BbU/wYiAgwKV2uTbPF2cBlkkOWrHQaYZ2aS45
0IVXHyPN9+UQ5Vg77zdkhs1KX1itQfQyG/nLTV81RdhdRJ4SON74mvlXsFX81A8nVh4VvsRBxxjT
4SYHlrbjeLxFAI2XLLADSvDwjtd1p6Mr2F6g4gqMHLAO4ma46awQvcXHLaR/DW/KCH5sGkZ6BUII
M7tkfI6V4tPvede7Rxp0BnHUHw02aJiV6w+zavpt4h2g9UNNW2msMmxew+pMMQ5gBtwGhpHdRw5K
N+cHG4c4MFzYeLr4/soY0ubXSuSevKQgQVUxW1Wxx/eHikCatflL+DaIlDn8p8/fh/ELGOXo0RHK
mYa/YXaarEMuvGWEE2DuDC/Xwle2a2xv6QXc5zbVDgKH81/ZhFVb0XN0Uvr6+nlg8iKNESkHF5bh
jwFB4V2+NphyJq4rj6knFu/Rqa+tdeGuDrFo50xumQSzlNM3jgsWmD6VmF/L1yOp3i5iVxnR6pcD
efn6ZZEyzKL0f4E4hm2l961CClaZ7B75me86P/FFWmT7zHc8UHGjKV9gpFze5m0+O5z0JAE2HP1B
f/cAFX5+iC88VZ1x/pacikfBBTts0WVGnndrZYRb859fX3chMIUIet7GrEQra4u6PXF+JSK5rNE0
x8GaDMPm3dudqqcKpEyHQTqbkH8bIPwq0/7wQ8YFvyQcHNaBs//8MbQhM+pwCeMsWywRPoHk9b+g
XfWgOtsaeN4qjK2aq+Bq4f9NvDQBfmPaPfX4EdurjW1761vziRkrFd0zXUm1Cd5qvWj94U0LBSAp
zwOUByl3O7Sijhan0cGMUZIXV2vBo3x2F5qFteHn3MIMBARy6fd2w+S7nn4r8yp1J0b64HBxIJ8w
teFVuBUbmSAOBF1VWfTNSzKTxB9diN25JmrO8VH6vmJWPDeaX+FE2qlVPij6d0fMSngZMpIP+ko1
u1vSRWJO7/TycTLG1ovPWACSXQAftj4SPQ4fb8+bkMCJ7b6cWO9HElXcQyL7+cdrzBORmM6wfyrO
rxiU4azEgYDMSdmtn6FDKIaXOFTcdoY8TFedFy+W1kbR32GOys+6RU3xU7GlXwAjf6BH7U5f/9Lj
EqwaSiJCxJm7DucI80S+Znl2P8jEYfD0gO4u3GhwJXpdLvIwPm5B1MSP2RVa6Ky56zXgy9a96aOd
bqiJI71D4W82C7c0dmGDEBKhQSSyb3WYfuUKM2kKsrWqZPPMtRuqKVztxsmxnBcOZ9vOhuJAOqT3
86lT2h0JYg1+CQe4bartUNB1S5JY8MtMJixRn4voYmzjLTRcAWEYiZr7Yyt9SI7Dbf/elGwN8zYW
thtA05XsSKFAP0UyXH1suyFX51Iny8Ki6qwtxfzAMMKHXyKEDsw0rp2Z9nnfQrxXEKX9M2hvTrrZ
IEePlnUvoyi476xmrpBj3M+2jGSOCn4gSuGfGVBCVi6MNYa25Cz8toYcnQazwB5Gw14yEowYKyei
l53XP7Ubus7lIcrV5EJhqoUpI7sRlW7nOpTvlmaVsuZbGEQoztHZ0jXdG50bQ9FXagF4qvUsgbUr
SxmQNOMp8EAbc4pcUcNPPIs857vG7WjyPrcv6Nnd+BX8wMzTdetzUASfYZ5vNT+Ez8wigbHk80dv
/eCTL/jerkleRn01Yb7tWNfMHxqU20AvDV0vp/AcCizYdZqPjZ6evEuxJcku8ZtQ+g97ibQXkU+f
ijJTrrkDu50p5g+H1zjhi1ny+R5L4zUEfKAfet670+abpD8ftOY+Ap8uXnX0ztvFgaDwbZtA9xvG
7EvV1iJNpNrKhVly6t2gnaH+zpkAkbytVD8om26zJINgwYWtri4CgRyu5DvLfSQkLAL9fc2MrwEa
yYRgMOvcM7myd8BUaEJ4yVCAP5yWSwMsfybEa7mCK1PM+OXLQdahlCI0MH4cZzO3CFFfGGw9toA+
QtoWgiveYeUe1kTdiOvZ5kCo7/T7J/e0wbdxLLpStqn+HeuXRwBC6RL/NjKEr4KzuMlMKVgZgYxo
X6vKXEGMj9RueOd4uYqZ1QFIAtyjLdhPM5xs9rjFZBUTOyyBZgA8fXqEuaea/+uXNwsQFyXecBRl
zk5JHv9b6k85lhZQOsZ+EVAWFJJHE+twhg7o+8Fu3742pxFR+qT23+Z7eXg2xzi3iZDRuk/KCGZo
V6xwbBlhIJO/mPIKxLV5DZxSlgBrq17ffU5CLxl7+QUe1VjhUrgaxieFsb8/lIOsDrmwDohDiYQX
x0ovAsEZBqE7Rzgbe67YpEVBrG6bK69X8Fzs7OkqWX7DE6YOonX3TpW8bS5gulmWrGQzVLVN63be
isBPh2QzLgHfCNgqS0cGVegxZPwcLWb20suR0Ns4okvINw30TIsoXn5uOYBlc60IZKSdcGXhgHUk
AE8eJId14xh93D94+WIifUsIw3kuEABenAw3DwxPv7J/WPUlEtlGpa0UT46DrBswwo76rC2+tZRg
zn3QdGx8Z8FQ6uAnAt3EeoM2cEud5Xi8MVG4JxP5SGuV6+tSf+3iiHaNwmsEZgS0ENYKPNqyp0TS
9xlugwA15EWb/l80DuUvk/ONToZIz0pIv2L64qoP9mL9/vOvf+EYiAMA0uKOo1Jzxd6nayi7TVLY
AK9R2lSfbkg/nTGqoLeJUrvFRIDFaDJIOXRodFCvavd1QCs04EABaZHIq0IoouVvQasCqaq+H2SQ
4YtD2IhpLS/1x3s1//ZYxeC5IF+rRVLAPS1Qk2PdNnpsJfNPwvJLLJZfB0evw2YSGzzddr4SZ2yq
MlW3dwBf9UkvYPDrq/UPcwB8JtHgmBljHydWrIJ3AdQcTlYHVdb/o0+6Y+8rLRcTknuulT5PikrB
2g01JZW4oZ2Pxz6TYHGdw04hyI6k04X5pud37eHh61hu0VcWTItVjOoksIUln7u4QfdNxW5ceGYL
EDIWzW9vF86eQdIKpiCsrVqrPjePwdClzVZsPasOsl2k05EPn+imL09gN9iVrp5v+Q5jNlcVG2XY
WAly5t8uvQye7ZZDofFk2jW1lzCpf6dp/E8UNwujlOa4wPl06uR0G1ZzUN3wj6Jtgm4ytnAqZ3f/
MqE+mYxzlCU52zywXC2yGetA5tnoSV5JGwFce/Vf0En2yF3vW1QeiYWu1biu0Hl2dGCQGWQrHobc
+jFeCTqwKkawQOuy9N8gCLPpiP5yRoqnh/Zab15ibjz2RgFAUcTy9aOkX6mIBRxpUH34bQ+twQhx
Nq2YqrLkCjAq2g9etqF4UpXyBm0lw8WJCDbagiuUhPeVyVKWKzMAMzIZz0GRdZ0TAm19fYmbH8BP
lGAKedsT7HlAETYubTAoN4uO9oHdIYNOunAQRQ8HqNxWTFjpdzSodf06Jm0jmTlD4sRJmTwGhBcR
L1JTMovq/l1UH9L3U+U7FyWIv9/5iHyJyGZdQsnIoN/vAheyfCfZRFgfuab94mSZgv3LxWI65YUO
5hsrTwh51+wQ/8U+DZPJzvPtJXO+hQwLtr1DIae3mIzQUGzcwzRzrzyRMkvx8hICMgor4SzSuBPv
t3YWnsJD6sBpHccYUAk3wwlRcraHLI2evuu4PZgq9RlyYCZ11Fa2cn9jzE0oqIDVAxXdXZ1UnQTQ
C2kbgeayQXbsnwcdO6ck3OIKwv1wD4VYeV715ecRg61Wl4kn+o5IliTG8GV8Z5vuAAjMphKIwJgl
AbxQ+BPSRExAHsy6XNf9pGtk+6LFL74d1wODZNYD0nbIqC599l3pcLN7pkCe++x6ZaMcj44plHFA
d4JyYa8Zs+vS+mBD+SvrwCV9YCSSKOtcQnTurjmc1sIMkBcv+iwer4hldFiGyoTnRoTiHdqOJ0Rj
0uTFTIqQpND/n1IH1wQMIMFdMUqEAXMleb7i5K8S4h8JyNxfbFMm5fuebgurli09Qsu+zT99cDPr
Du7JDWTxWOZDdOGOd2rE1mknjLyorQU5dZxoVZauAQwITYDOjB763T9Ca3wwi51o6E64reCIKY9w
88ceh5srWS3wYeBLQOiMcXdOd8Q1MGKjSj3CiVnRRXuhiggLQ1uHOZ6NpNXjlf6dUH1nF1Tixivp
Cq12Afe6vdbCO/M4LD2oy09O0vW6yTXDWeS8wMYaYUpWWZTJnchc81nF+L8tUM1s22Um7vbV/Sus
UIMt9pFBfGkmUV12WuPgGYyIwfVEvXrQ/2zfDGnw465G1hFRVrCXHpZSlE/vNQIcGg4J4d0/Z/uf
Edtwa3PnB4f72EIrI9qY6l0KPfO++Ov6SYn4kjGUTEy4quMr+rm8UYjIV+l9Mc8XVojrvkJilvNi
y8O4id6V20hSh7EDX3pzXY1rYwDqqBdFX2qltFNJXTodA4kql+3BrIAabJvH0VQE02gMkPnbxAhV
BptKnEIa0d1zjyialnU7JC9853ULRmpGYgcD9RvUfPSsdEX7pw3XbSADO7X49s8paVpCGe2QQlZ6
aFbL8Z+qFNnC5xcJBaeabSlOqtHiiea9WkBzdMFcW/6SR3i+Fa2pcPO+VPHYICbj/PSG7E1F9Er6
iPse2+piR0Z7N0UlVnwRQwRzEVQms3uXe6OEg8i9mRUVVP3ajxnjTu0zmq8O7QuoUgaTFM2gwEqG
amiq/f1BNUwOwuzOc4MPD8riq54IIlqk/w7ImZYWtmTnAVMtUFiYjf/y58G8di/lF45qGCS36Wqu
64mhicq4OPLGtJ25QDFwZmxB1fAiYr0AVuRXO0DlUI6uQznW3+LrZCdUO2aDZh8t3kR9OBXyK/4s
KJ3HhiTuxTIEchAdxIK04U1Mz+navoIXmTFfVP5MdNR6aKO7bHrtyXiB+jDirMqkXD1Q6yYm6pZ4
ulyiv4gL5FEs1p7jh13loOs5RwE+isUfCKEEx98upCQcus0KE6XgTe/UrsnJxxQKEunanbG5KcUZ
MhQ3JmqZH8HnMUwM25u+qPJMf9IDDBJcl4Hat7oq+woyqDWGjAiLTtvfhNZGghAu8EJE5JOL6Dr5
1yhmmYNQUhj+b4gBGfbWk40dwiiBoAco91e2qJz8VePw9Pd6qy6LEDRgvnyhSRgyjXTr3Zy1AQm3
JrO7ZfRXUeKwjQYDAlKNToS/R+PDkvok7u0GauT1SlB2nZ0S456R/m/CmhTE9rUvtdHuWPYuXPrs
0L3dYkqTlDhoF6v2Qf2Q+79DfQGmt5WUo6oG+g9nkwoAEWk+W+xyyg8bZiQ1Hlf/vHfFpD3VNu0u
GZhT0eQxqnxHfe9iEVtUMSoBpkcK8o20NgmuM0wIyk/edpdeucA3DIO4nqZDSfixrl8wyL5P0SBo
nIg5Ufm4MkE7U+O3cdJWyArBiYXuXS4wVjO0R43qPV+r8SXOHsvF1g3ePlKTCUqPCgbwyj0ebiiH
/xiEqitatxfl/tnb+zu7iLqgbThp4mKF4dKhwjG5Nkt9q2/T6D+XbDVd8AYv/1I00OKOUFMvksjK
+IvQZxL1K97HS/m8pQ1t/Knc3akGnPJYo1/ermJQkWnwIUPpYDo9FwEXNP6ZKTshjZs8k9jGBIGS
01KeTPhmSrK4/I56onsrOajHPGQTnysQO75KWSbqUHwFNR5PSVh1rQBHTienGZXHNf5zke7Iub/U
c8YMdDqdRGfC7qyyPlzTta7bw+BaDFjSEAcYzUDwJmcyEnwVaPCAbOu4ZpRmDUAUSKqepUwC8PEw
bAlxGgGcr/M0hv6cE0al1sfr40AWT/F7o7YuT0N2wOaZcj5llA7G+iGsNdsqFIM7JpVhoBnz0iLO
KPaFtaoy6k8YRV+NP25T9X3QvUPLLM62ki8EfsXEZbvYsnyz7g8G1YprPP2sDFWI8w6FxtBZ71Iu
0wltPlh3h8FCeZaxmztBzjmE9T1MNDHdhEcLtQTwJIZTCrHVWLQpJLClDOymnK9re/OJ5Ghvm3qS
tXZbZA4r39iTsVw+amiupqS3/WANGxwRfRugKfIO5w9ejHdYpYoLzxCfHNALKb7D7ii6IqdNa39t
84tf9X5bU0IoEg0C7J0I2sNACvTPisERjTsEbsuw/10ov69jT+fmR/gR9nhjS96KxkxOtdUmgK8/
vK/U72+SWGadkmkNvfowQAaFc2fP1O2R6jV+rpYDPBPUqNMDmunVtG/ybBDbHJKrT2lzUtoefCIp
hTy/4VFooh2DZMnOKYM22yqd0Ko82x6hGOLNa03d1tZxqviYTbTK7pWMtDI7+jfjRwmb6BMBh97x
HBOLOJdY+dmxE7srgSuIalj9yf2PDhg+k4kcPQmnuq5DTi2zTOMncnhjTYdeewc/fEsbGzYRmF2D
i8YlkGNhbzIJtb7RXRTn+64OU75yTEH3DBn6r7azhy6zhPlf25qhi5rv8doUEQQKjjfxIYsG8OVl
JdUITyTVacttF++Gjt8kVUpyAUANUMvWrqrtdixIA1BgxrhZGWomKaokkLVDEVmDjuFf4Wt21eY4
13ZCzP0QSH3YbZLwW5WabRUR2B9iN+PyLRF5u2MR10XzQPspD6w/NuK143wn4Tl/y+MSr3sJsRqy
2hzkN/fNIzxRJCs68i4qDcRYPHz0vvt+3RcUQTAuaqjLGNu/tYbXFQihrhnIDgNd5lleS84yhKbL
YeXEoNfrk79cTdPQlEs5ycPllBbpg2OQhgIkpcX7OrWbJR2RelgHpmkz7NOZ5MJlGNymEoqvGmzt
FukO50Psd2wqGY0m3OkH99rdgkvx5npaUqxkle+HGRbisIppFd+T66Cixk7vprf8oKXIFVz1/n3n
0jykLfHdaFUe6tDnNKpTZSo3bhQQdkODcauI8O13bLHz/DM9cPz/pqpYjqu0dmI2heJ2NRFzvmbl
RzJyXN2a98uufWz8IYFrXAvOmU/xd3fTUyo9M/ESbj79GO4zPJW4qnAg8gCfmuHd1S3DiynwrkN5
KJSxFVsWnhzw7kIbK7fQIL7f8CjZNU4BU2AHRr+9UEZ/Ik67C8GyRDK5znSRxWnnn/ZPYS6zdjRt
AlwAkrVDUQE3XvVzvh6l0vvRGUADNlKp6D19EBLmbB7bdN3j4yZcSSl5L4NY6J3v74dsQoZoFb/0
CmxU4h7Q6hcdBdojSUyPMwe+rEGTkBnBbgEOAyC746TK+fpUV2u5h0nlyyaVaidpcjVVMmDM+Agx
uqmQqaXGaczip0pWHiUJk6z0xPnwkEYdtPbfViTbyFZRr/sJLsN77Ia+Czdiia8EgahGroaL8vYr
8NyyYs+es9m0w7WnvfA33i1yE9FGfoGqlLIxGhan6w2ZcDEb1YIORXcohEzuCXOQr7r5hSGH+yUG
PdbNbJSQSM5+inj7wkx678IRehEpgmJB6D0zBcGRYmyd0CR5taleFHpinmYMej0lvlCfrHGOyFJO
NRgxyDWJ3NQHjJ/bI1duxi00zvANOTsdwZK6GxwmXWnJ3DNtJpScUSgoYtd0wiTpTG0wQpXPaPnI
1sK05iVhB0Ld373DDzV23H4X/BPuDglIESYKudlUldlqsWryFzU2AYcQQ03ECwoHRiUrZ3xvIlFq
7CRa1GiEvWJGLd9NVnfMG+yF8uzZhA1xbYCop75siCs6g0hxqe84HZwBx2/rI9q9yNabSXlMmNjl
omN3rrMHkhJHg4hXbiAaKvjYOTMTPDA0X2TIHZiE/bcAGLmyNcCCWfNQtkw3vGhgtTR8NIAEr96I
niNOSAOUZKNWDU5roFpFs0DuaI658NqN1VOVwxuggNGlZWo58keZtl94gu4fdUst1HG81EfleHFf
JxoO8sqpL16ODfKbxcKrcworpXdzgIy0WVu7LKHP/01gzbcXbGG5CcCU1ZMOhPYv69A15Esmjw9p
QHjzWwUhcfHjIJv5gkZAGWNSX71kUmB11rkZWxanWc5rTX1e/lVWJI3CnaRjt0wP91frJ41P303b
yi1h1wCMf34kTOca6G+Vc/EHi953IP65un0qmolnqZ95w2UFyYaGp+RiGK0tCRF8jVZL/pfeKiPj
DK14mljLH6u2Y65/8a4oN+7whfORpGJ41OIXeLMap7iv1ZMZe5/JurOVRK1QX1gxppFYeMs/G0pz
/3d9Dptr0x+yrtjsc6LLK8zjIrw9QukXKQnD/P0es3eI/qOSGwsvOq4/+ZhBEb5kD8ua/l09TRxJ
hdhJUcKx9ADgV1gy8uehmQQqyewh21kPECXCLHFwN97cE17dy5DvcHqvAvvTaPsKkTYEH8jhPztJ
i7Avffs2HunKNzwSQC6LiuKtwToDQNXS9FKdDhWnAfWRb2AL+9ajCvaM2hLN/imrfVgzpywqMisK
RELYm2qQQEPnivLCfnkSacbuU80L1QNZE/rcSondUHGDX9xKKKdrILphlDrNqt+wJ6iJcWytw06/
AJ6TyA2491Dvy2jA1Ww7kvt1BWQhYKFpjtopS1hzyp0MttUTQorr3tLHDwsWg+YenZ4trA/MFGzM
Hk74YB3BH336gOLgxFSmUlfZUNEEzDwsKRjNPoSEqHxvKbLb8EAXNLlVZsGmktgX8tlcdcIr+79k
6dvjfifMSs7QMMViZgJCq8U2/2YsBfxn7TSYQf1q9p70O1QQuL54C8XGeDYk58ESE9L42uTs9sEb
tDWXHsn/aWSPkthhSX3w0LQW9SEs5ekakjYMhZPIabOb836QnL+o8cTj/8qAXJx1SDHtdKwvcx44
KMtVLfAZ4bErq3N8Mb6k6Of4zLa9T3oHJFisteA2VddHav5OHqriNrmRQQ6F/P+01mIwoK4GLKe8
4FfljIwb3uRx/x/m2+M+MMAQLNuWofhOUNs6F59x+k4DMPn4Pf/fyZFtAw9YlfoeG+O/sMGiHric
yVzMkAQMlAFh4e0wGJGGMdKxlrr813wt2TCagyuVrRUgUfKUuGdJa9TuZcFFip8QXfZxddDAIdpM
fOgshCjT+7WkGO5820jmwsAYodUVu6G/8Z6pdFdK2OZOh2rjBuio52Jt/5+CM00XgcvAck2zEZ0j
SeP1ReVJLYRg/ysjbZaowIwYkcfpkJ60BC8h7CfgUW/xLEdSJfGgnVgvyfU43Vzb0m+5H7Lo9tIw
Zzs6P89SxIeWM/1ot5WzJbzuFhMOgiB07l96tKLjA2VrZYSw6Xe7hQZHjV8cDBxr5QP1R7nyocm1
17JwERerLZedFJZiX3csJo5EE1VjJDDo8RRayGZYiDubIpHZWQ5ZxVBpG+yOGSV5L/qqumr7n3zu
p/j5a5R3TMiVqAtuEFZvAgLIM2aQQj5YIc+PAVqmGPD6eIYcYSYKME18mSijYbyU0njlgir6AC64
GJLdejPRu6209RFV6T+b+bV+txtf32gWJGOi2qFbeEizuOXoeTMp6DABAVIjrpo70uqTp4P8Y4n7
XkH8fQ3mJjQ7UYns0KrJS10cp+w6CYFg2mmRfBisbhjKZhTXo0Vo+F2ognW9J5nFRWlkqbaGnrHo
yy6Oim+/++sBvACa1yYGArlCLTZLHBRhpaIH67WSsj+sN4ItHbDyU3Y0oc0ZVXoDOhYlkALWDKnS
DmHbmhHO1EalFf5pbXM9BlFtmX1jbR3ahyW2D+VF/xqA4HYcK9Rf4LNHpF+SBR6byb4RbkI9N8Tr
5heUB188JppXoQkuLpGBjrrylOa+XYOEI5EBTSF9iMtRGuPQgDLwuk1gpgzlTMOX9avZco0t1I2g
pWzgcUmbbk227anzQESy0EYYRVRRDF/8+6+tGKmkJBgvPt6AgmiSwql6HpX8lAjUPlR0hWxhBwCw
nkUltHXoUk6u3JCLE3z41U90yZgwfihNVpK2M/XIPE8oTDAX28ez+BJ8zQEIe2ch380yG0kh7lzD
y6Aqt79F3UOQN+wmKA9DmDFisBBsOeb3HqCwRz3ylNPbCZ+1/FV1KJTOEnkOsiUq0Y+mZ1FhcXBa
8zV2+ioNXI0Hka8qKcZUQfwj98b2NDnoosA/Bn5pVrZX+6FSuqw8Py6Dw4J0LzauHCCRPaES12p3
FzW17vehQZr3tuIYhBlf5ETzgo6y+Eob6CfRQKOVpmK2MpkxnfA2OQqDmAtYRjKoq17G197Sq/2C
HDtQp8FFqf21amCS4oU/N818TWDAz4ZgUsrcwqwLOIAEBApdvpcr897vvNRChQzd/ht5pnPSxSyO
QXv1Q7WRnQGD/buWJfFooCz0tL3HzSunR0QWO4aNNJBFoemy7EVjHvvNGYVBcs8FYDjoBGZFX+zX
KNrwmlyqZQk7XDwtT3CKinfPNLboMvD/HAGKzgxR89+OriCVI6uN8M41//XdNbWssKGZHDtZ5UDk
eOU7Kxd1RdRUgwO1+fSZKHq/n8T339tAy2HJOJG04KN3aIn/0psVOUIIZbS8fMF1SHaUmaRq8UJf
EiyQtqV4s3h9l7gY9GWj2Z4zLMtLlJV83wlyflqk9tlQzAFmgRXSmvWE3Hn4ZNMLWlVnbXeSunrR
f9BXft+XldROGLK8WcpOUtP9GHH2IurrFmftMzD2T72xeqKdAxA8kiI6HzO1L9iM3epXRCC56Uk8
dK+kW6Rrehk3R81R03Cu0nLZt2ACAh2TOTHl8nNLHVgtVC7l532uZuTkdIZ2+HMepTjGyjuLZcO7
KN6gTXbhmJjSjtpU1Z2KVASiCIfjbZEeF1+nabYAdCGAmDrpqM0pN55auinWyLom9rV/BRVgKFon
iKIOHO1YP5EedWCps3hrt+59WssselSuJ6aVBBYilBr0Q+w3/EL+d0miYgqJdJU5ga3U4BdJTkUD
HZ85Jtmp5HBOuaAQjBKjhhpoNKxHBtzZkjYe74SKg+9Ud51HBlFS1MA0BZ2umpDzWBZ+IC11ZHQx
q1Lxjh8IxsqvR1eiQR67vJqdpj34bfW1ldzKIx0KV/mZjgCngO5u4VOHinNLvRNKyHNo79ynQQV0
/K/ectuojz9sz9lz9agkMgQjlAEj85rj7L7aZzFnVyZu8mpCzE0NgV89FshpalAuoCvyuLKG/xi7
n6PW0MbQi44W1pN6jn9w5g1J62VmrWShwtTzA9XFa9C/ZR1gh4JJXI+b2q1AXEWS4UMzAGiqrwRK
t8QQ6I/cJbN0UZntRKfkT7g6Prvq9T8FA/BZJWIB5tnjo4E2QNoCvvNi2KmtYChuzeWuZFuujRKQ
faqNhDeTG0CgfbtFihyf49+rMS3DPdbJxB1Ohm1DwkJH+R4Af0R6g4BB3NHYw5UmEbTY4E2nN+a5
WH2RKPMMPPrU4yQm80PxtiCM61UCbdQF5Vvlz1IwXm4NhgJbgu+ZNZXfbeSS6a53w1xdRSJ7q0x/
hEUWA3+fuVTGms6K1mA3AzfxgStcGZgFuy9HMHe34enrOl02ejxeReZ2x8yhu0f5GAiMy1X1xykT
5OdldDfqd4FEkfnnBdUPQd4ILBE9GrX2F8RF4no5PrJ12yTwyOo5EaE2KCwox8SJobfY7RanyC+B
TZLxzQWI2s5Ua1PAsioqh+mLAvj/NvgcaYFjzL4qSl/hE8SnJu0zmKK9Uy6AwKCtRsw+yXM3A8YI
GY0odUXCbhviYceLNfcqs4+WJByi3/rBa6nysYN8YFUCSxjUq3ZnVAutRfUous3yjm1vKjdZB9Y2
Gv6M6IBqbQou5UKlR+ElyQe++zFm5kDirLPaKPwxvr0988O92ggd/UT3JyVCKsbQD4sHeYMTsfsW
ls+FFWSYFAKOIqdASoNfPBlX/EL4AdgC0p7xSyzkcufUe41jJsPafbjXRQMjOQlvgEcn4G8JXtdx
AEzObX3MfJK8OdT8eFDLLlWD65hCiXsp7A4gulcA65ple7Bzs8uZHEOnrVvs9zEdMJXfPalVgTHY
Qj6edqO74WqWltqpyVWq9usgoXjRUfUg0JGB7X+rmJbix8stQ3S8aj93PmgJtV/vQZ6EKArW6LJB
d/Msq/u70qDqi5zWCdmd/l3/qiC6EIIM/fYvBZ8OEf8jFkcvT+r17S5+qRy2VlOH/Jrm3letlwFr
cQ+onaIPHKd8ZLhcOvcP+dqgcpXDkc+Mc5QoH74aA6bRo2wyJFPjbTHhOFYZ33k6eZf5j4YpyZfn
/T9S1O23NcGTK3B2Pn6a4us6dg/p1RkS9/El+G9a3iM8zr1OL+UuMGBdKT9QgDfX6AmC52EGfc1s
D/JctKZxJi/eIuvyEOAzDZRRy5+Hk02nNlZETfRvs4pKZeTQlgXkcWh7UeeWgQaq0gkSSQau3jjE
skM2jCu3d8Jy7tl3SaFd4bO01ADj3tBKQ9r7rjVu/7mT4eGbnzAQaAkGDDY/XyORSzDB5kSNXo/+
yYgV8GGv8Q2pMVBjzGZgAmaprJ1t2hQbTZYNOAsGTnOZDy2AddsdQp0buxN/rPjMBKkyE2crCHBO
twJYOFlg6jaY5fn1mL7ilYXJ59VrzJLZGJ4QUDe7PlEP0wUlc2xKnd4wY2qTmI4GEKr8RomNFBV6
cmDffNz2ocHqH4ZtTeEIyt1z2plWHfIFObXXE8p/xivpmkZ68VqumsLWD2MyxWnHr2MOxHnizpMV
aWnracCDDs9QdFt2pd/Oggv400Nv0IC1jZHbmM/Se9lE7xnDmjy+stLuR6yHFM6E0lc/6jEOGD4Y
MpoE2tHyTLTwOwLM2TFd8lWrt4NfTnu6FTdS6/PkwciZPSj3h8OkYuv3jUk76IQtaae1Iu3Udnwt
sups0up/Zmeb5sErFiNYSQUe+ZhFew1NHBxQyjnha12hDiK81L/MK7E3BcoYNM65x2cByZQ0e6KY
Oml0NQ+D7IYX5BlEVGHmf3Nz18NyQvGlMP60IyPySuMICe4ZLb2H8VQvRSVFuWqKz8oyO8NEh0c6
tPYpZzHjh1NZ5LG/uFP6hXfLbLxeNjxAV5VQOmNaMgtc5oCCLhTxfOh8h8nQJZ/h9Hi4bd3JAZzC
gXj5iiWNvbkwAJJKNARMmgg5ji+O5xv2/5AAUL4g0bZVq+Msir39MxUaPQyU6DaKaw4H+WIpz7FK
lJZEN8hGCvvFL0BH3s2ptKdVH4PjOoJsbnC4n3RMmF5JIzty73sByzW0GsUJUqoys3W1YdUYkymT
utrh1jCwqsEzpQHpe7BtU0N0M1l59Od794zcooRZQ19GEfW2NQk9YsHvYIzPxhMAuN0tVA+iWVe0
39aSgJf1Er2dPQmShPBPneoZaFvasLbSA/7z/g5oEHou1JZESXgrKB4dtMMhb71ZpKCxSZx/cLuK
rI64i1vwqS9foXC0j5tbq/qflgBsYS7BAQxwJpqQBeE+SsyaGh8vBrP5uMG74zIRKvZ1HARZOuCJ
JvlD714wc2rqCMF56ZeiQmJ7fqj3LCUcrc0EIrKiLnY2ynL92Xtt7P1OFkiAT5ySl4nF1vdibGEI
Q563aG0lL7LzuhV9vBMNz2eRoQP3tCk0Rl4XsUYrk46WKtR8r2Byebc5dL4owijj64RECZb3kB2Y
ANVpUrkLxTIW8OrkMV5X1P28c8pdyxRLaIRZ11UNxCNhYZi2hyFnmtGYSAoHVQVyfr5rGsbYqG7C
uQEv3cLj+7uoT91HuolcA8q92E36r9OfNpCk35v+8stWIHw6+udoOaIG8jMKLw5JctntoMIIIMi6
eoqHu69hXJ+cVBGwsKsS3TnbZt5xGDQNcQM5+q0Y9WN8HYig9At0454FoUSaZ8MOKHrcki0YVxhd
i3oZZQDEX3vhCo5HnSEeOTHIPkxNd4OAkaNmOXuv9h2RpmVKTqiB0pwQsFukMKaRrHfrgkk4SwWf
i9ZIRPTh5TbQU2zIXPGMNCqnPOuXgEjd6s5zjaK2ORMZm7oy2Ms9YHtSM7/8NlUqs87LryzBK8sU
YQy6rFnvR36oTrQnL/N3ubSmc3RRlRxk2bMToXXq5rn0uNvSKsu3D/Wg8udn0LYxs/qiBXlt5Rs2
jEXEJ09oY+67tUM80zjQE4pzOSfLx9uhb0ItUmXOU9xFpfztZo48Fo1Uw+Hf9rJ+O7nWfFt81Cr+
dIseFaPt5pWtedtSAta+HkvIFk92EINnu9EE1LHcVoNGlSS9DkqA6fvZR1bY4GCzJCYSOyiPOi47
6FkhC//S2gM37C/aPP6lmG4JLwwWcgsFf2MHpy4YRrAczB8NjDpMTXADXh9nyTRZyBJgnC4JwS2U
pJ+7qoNhcMhEjPxLo88Wzzbix0tVUnT+uv1jfhcF0YhSshUmSu9z62FlPv317HyP38t/q3FnovYY
Zm9F5prNaMIvdUg76fq6WPsJvD7ZAPE2Ff0NNt9pLf9u1EFG+GmRu31TCE+Ok3dSd2bOxI6g33Ud
Tw3uZbtmQOvbQfXYpaHUU2G0eqos7LlRv5fURw3znMBVRMWY5kWpZ8dv3QqFUbB3M5DsuroV8VQf
5egyjziL+oUOypEZVDFeEHi1XAHITjWAWkqq2HfJ58I/GtJ3LoiaecHssxQOdFx3G979fsPqVCEH
1smsxXJW1168/6bMvBQG8EkzKqSerwKplkULjxW7bm768IjeO/gfJYEZG1qxX6dJENybIOqpROnC
Tn/TQgRC0Csecm/yHsXdtQVphB9SYLEnUdgF8byZN0pzjIk499gg3ey215Qo0fIPrn0oAa1DcN2W
oMrk5SnWv2OiYnaKpvX/BrkpIHKCsx30cD3HzNtCYIHXWxCRPSWYMqP5QKNBvzaWSzTYCaixATnQ
Yq1ICVTaWcxYrBPbzTD9pdtRF/PhSQ7k4ACbpSVrsxAGdN9HSvAa1RT3HV2o8hPt+ZBbU/Zz6TYm
btHyjSuI+L6jrEAdWiZ51aslFydehsNxvNgVmYN9+qW7hf9rLeOEr0Jbb92JR2H3fPKlybBM1QuA
Ul/8FUeaVC4dPrjHGBXSdIDO9UkaaKkfWDJTCIMqE+QEKX2MlV58clkCEAvyngAXzvOX1N0l+o3Q
rgNqmZoYi/B5NcC6MNOpf7tgVFCSUjLL3HXX8hpU7h1MinR8rZTRbCgmQh1y5tFKoui9SLB49nVf
lRXseuVK73TsIN4GpehZzbYiQLcpKeL7k4TdQdzfxKa9YFpl0n+zvRlXYkscVw+2Fix9rivYu/VC
5uYvHLAqjd4+F/yPMC1Hsh5ZINCXzxNy0ABYAWuymndStXBUzPV4ODdiUh3+vAC4Y9EGP7RPPKN6
gp8KKllyTjzL0s80e+kQm/RnAGudjXbA7kFtACAOugbB8fhF9xzFYbYEHecGiHs5+/+/951IpavG
a98z58EZXOyY2TAh3L0J3a2ylTKBvkTVPPKc8ngQu5xJeDqjMRT712QAFwfXpwGfnuGo60NviR6N
r/TnnLFksjdm6uql5wv8MOPAIviav76b6drRahgnJVjeeuVpU7OiRQr8aP2achGGHcsBMD8XIkp5
dbXbFYmNgSDAnHw0sOeXi11CZvbRTxyPxLdRfMk266MO2gClBOklkllyNm5QbvjajY1rJ4liKNuB
udu+rBuJNvKOqbT0MPFj1nHUtwS/fd+pJywYr2nzaQ6TiCpj/OqAKo0aA/L6Dm23SnMflD/2+mKF
7hs65a0E3SAwDlMZw8a4JcZrt9RO6DHg6PDLvG6Mls9SJ3C5fIRguOmt5ax7gxn8ulkWC0HTZ8Hy
XufqjM9KTr+u8KLmaaRHn1bm8ptIzZzAVVqBeJBA1FmHFtakE4/B9ewikPLhLSLjo5cakAUqxwwC
ub543vV8h01yKjElpst6MAfBaHmCF92UOxtOM2uDrLt5d+mn8zc38f3KnK6K0FFJWtaMvzT2seSS
/5rd2pBHYdAkNhi0uFA7BxtbaXEDwL4P7bpdqE6+w1bwsUH4dWGt39t6im54zgmNiGFkpDjYRbGa
oNXacRwmpK04B/nkVC3g4IbhpTqoAZ8QvWuMuFKevt8199Rb4mCozKiH8U+KAVLq8oEre2mT9+G/
IFu/q2tTnLL0dtA+gh1l8WdT6mhvQ25mNh5T78TNBob6UNfW1MgHeCIyCeQpXq4MXmklFowCSAFE
cZ20vC8N0lmv4e0FsPiDAL/ZM8TQjKVhXuslCoH2LS25tovfW/7GJSJ+BvPxEUieUeizKCXdAj9/
pABBFAVWNo205jlI/DcgRXbzSAS5Tc6PFZjwLN+Ox8BzuRZkCJFEgJe8iYeKS5745ZIPi9O94542
OUiKCywvL8s3e57tHtceH5JvLOYxTciPej3ppU1lhwDvQVQGUO0mfDLQqO4/J1RFzCgjuhEzY5cr
WktRAS1bxTXVVUY3OqdYrF6bLxbdbEuOIDAcdgWxT1z7nYBTj1nEU9FkUSD2HuqfRoe3unXRlm/p
fYGUTFOYgvPyPmRTqmDpWTx5xGPsnC5fabnUuW/1ZM5kCb7ridcfCbX/lfqWuktmMxnt+u3tRjdy
m9grjhtiVhZiVmcIj8a9yTf+zyK18nATRLlJZjdY5f++sqI5ROsKQJ2ITk+uAWi173g8tCas8UQl
pJAxgNCQ5GY6sSCRnIED/9SQZrzGQo8Ek08LdeB98GgkTddTFGLVgAWHFlyQi5DBPtFkBf1whcD3
8UnLMUtzheBP+/1lYXxFEVfjUNpwdsYxvCIKz1URw3xyeunax+dBq2V2MvHM5iKX8yDmg0BMB1xl
A/FZb2yBPmfrdhzTioeJQsV0IuPw4FLCh5t4gAqVhDyJjTPXBQPwyBAJS9lbYWXb5vtLvfF8rXzH
qn+sqrpvBAweFc86D2tgJv085K1ub2z7rhnIjR1zMaVBLKlWMaGCHxBpqCtOIiKVA3LxpqVU2iwV
O0Y+3qe405gHubMlFwnnrTOTt/iYhzrNAzklUilg4/4jk3kjcvYHAeAOA+qJB3GZ8/FYfEpoeY0W
F6dlXCqDyQ+vOvz3MTLncqN4JAAkswjFSZbO9QvlxUOfzwtRoV9bj4+8a2L2H4utt0IRAKaryyJ0
geQJ05vRVPlYNVaDgIER8K6KVraw8ScTFqgMwJWG3JqPT3smkGWEwkGMMdUBuvtQVa6xVZt2B5/l
zgAGPfAHVapVWbOhAcLsK89U8C2ApMMCV7ySO/dEZH7KH1Fu8WktnnieCf67/J+P7wfHY80wP9c6
b9igkWsGS1PV5DEiG3FowS0NotChB+/2RPP3im8CSoQIib/cxxsaUGPA8COqmkMQymkGq8WUM4fk
5H0ZEkIjDVpArCHdXspCDALopy0f51zb+8422zKoT5MtBjS2Q4WCrbMw3WYCna9/zBkSFgbwYZEw
aou/xjOttc+EiJ+0yI3aSlVGcDah2s/59Z+gW0mNOWEhJhj3IcZ11Q+8Fh5MqUShGN8p/doKfQdx
49fIigSRXj7VTBb9b4c9FGwX1G+bqwQ2c5CSCYTkR+8oZ26hTYhDEuzrc1Z+GVQhaAfS/i07eIX7
EFygBcojktYLqOc8a26zoE/K47qtfYEuv5P7+gvr0OyX1cTl08+Ixpbo+Y3/ppGQidfOWUjriPPK
HJ1CieKAD5xDQd/U9ZM2eqbRp9KoWmqtkdtQxrXbD0evsQ1UzfIqsqprLplyk9Oj28EtFPAC6Ur3
w55q9iR9xAyVYBu99zFKb71NI/AJCuUvvhNzLnsh1vWJgYAv0M91FEq8SVmQDhyBAK2QSMkfHkeg
LcO+LFunRkDVE1tGzfOYn6/qat9zkdF0krvokZDYrB7GW4O204VC0IXHCH+kVUxw7WDVUXPH6oED
p3//ZAo5ThGrfIXaakAHfpBVGpfeGZwVfEGhr4D9JwkUp2ERZsMDDb/YSSk3AmzQlzyWhzfvpMRH
/GP0TZ8A0krdguxRfFmQNGMIy2HikQPbSGv3pTPhIcG9UQT+pNdz28pAb2mTacSz3oXZWRKE4gfl
nClQETf0dMR2a/GwZMOI+8qm2bWpd66HDQx56YfSkBwh6FjGv8Qxo6Y1pnU3X9oLKNptDnhMjZjW
cHvoJ/JBMGaS6BdxSa/PaMVHPvQUl11A9SBa4fezQdmPfyn7n9y0AvwFO0c2o8m/W4dWD1V+08+b
KKcz5Wal5LDa2IgOo/X1yFi7XK/yv7rIH18fuepS99uNwSHQiaHotjntP3KOSO9fiavwddekc8jp
e9dWIwyxEHt2Oh4yFwXrx0EQA+MXAlNvY2rTMBK7S4wIiRt0SiiRD9qJczaMb9UyOwG+SLJZ+/2V
WknzZz2Niu0K4guKZaO7Xi3IzvQNR11rHiDR4j5u0kpedIVG8dF+NCBfcI+nI68QV9s13mMQQ3cF
BJPgBZH9iwbcVPMGhKKrIGQXRi/nsJgfpDyTfxWjEXzD079b7TrB9b1otpgGCDHW8YA4oUHqXAwS
0wy3kiD8COIQswp5WYO99bNzULOwM81QpBjqchr92wQJm3LTyHm1MdmBdj7Axx1CVoRJP6cbbE++
gfBPRU5MJmG2RICLOhIoGfAwWlXAa4e0hyGVlOTscGekCwqWeAQUUroCZzM+9Ew+VVWuGjQ+xTJE
VW8PNYqUbhdosh3GdAYY37mXsdny7PMC9GWr1dHA2gBjOtSpJyj6kcGyBJELKpmlZpfaLZdPFoeJ
WXQ8wFR0LgWcYJ2lCog1zm7x16YomLpK+T8T//R2nrYM1k2aqicTNh7nIirozRtpOwBZZPdWGpHz
Nblup2XTLIoBcryYrA5qzRezz04xvT1pLbdGOo5r6JKDjj78qG5K1Y9PSdUhs8su9s/35Xl8cX/R
8G2pX8Tlz6yyLAmFo3vHsv/mmwhrk4sMSD+YAaNxr92yySAAb9YuEq+o8c3EKL2IGJggTlN3eX+z
aQKiDY4UMUJ39bkFJ1WSV2K+GkU3jXEXMeIbsrmJfW3WXVHCD01vAeKzuuR+dLbnVlDukS15evTN
JbWxBsbRlEdQobf2pEPifcBDUtfNAquerntFqVw4XeFxWHPSzJPcfh0BMiUXPGpR3ApBmVvenBJZ
2KkceHV7+WwgdOMW/os9upjMnbz3HmQKGQ85XKZsJHfJ+kfXljNzMKzbPQd00nTKooqyou/6qrCq
8vSBseWplFTWhn0RwBTRbBvG70jZnVUuwAY2U5LRRrwftBjqKEfqLTeN2yOvWythbK+u9ixenv5y
GqiY6KN60x4noQrGREwVMUa4iO5ZtBAlxa9ZeD8yRbA2dJmVVsW3NZvOl9uDeUNqnzbyrS/1Xqti
UykOuU0ll9VYSeizECNSaqI3CovbqiQ7lVRm29UZnH2N3+xfjlygAJi21XsdC5V1QumLS6zaEXl0
kbd7drERTRU6zBGamczW+Nc7ska5ycSHe9HL4WPbGmSSJrefNLta7K7ReMB42xJHx2ERapAIQOcl
yQsN0kFaRbBUChxWtpRkAgvgv5wcQ3erDsyPaCoA7nngf8n9G4ug45PiVOFaF4hP6Bu/IrJgrYk2
4sLmDRVnkB/YCKMpy2Dgiz6pgkDTFe4srwGbPKpYAdS5My6jKdphJPw0TQbHX9n66ODVM6YDk16s
vbnh0bU+qNK23QighrN997EIvfWoyA5XFFASsx4iWHOw7kAlFoempqX53YZac6nTiT6O96lK+Mxm
yMjBd85HxHT++I3biOtdZOTGd1yuIMmyOlg9Xx8ltneR99w/HGEa6CNjxTCXpGcSBg77hmu5iZFL
/fcQAOFfWZaSPBPd09wGJSv/mTZGSyPixr6IHd5cd8Mc4F1iNHPelo8YAyrzJh7o0H326ZQ9F35Y
a6WwP6GEq/qCcDL+cCqyJHnuMTEUYfZj6A/87CmvIXBLihxBykl+ynkhHRimmR01rc9K/uCsrlI0
JM5y/MfIMbXxpZwCRANtl1zTkXrK/zOCEmBDUGgqsKWPJCbMsVETmKZuOEDaMONGF8NLpTX6rGlp
nb98WO7HcC3BM8S8aBRS+6hTGTMSwNKVBTgfbQJkE9JvzK5vjurqQ3h04mMmpN0gSXawKxooemOA
3BZkiFygwhx51i8HXGbw4wEVzTdDZoMJN4EpFOovd59Kx/uTHvU0lOJPttUh2pmSGjhtL0tpIziD
QplWGPE6pX9N4k2fUO0rR6jRirlW2PQ/7pXI3OVsm5Ne/J3bEW6B7nzdKcUGEnCR/YNHa0gLtDFJ
PrczTuiMc/pusa2LOxUTBCHrRcWgO5yhMXs28l8dz6VakAwmao0j+RoR1OrpeVEmc08Fb06YykRX
I9YAlQvZUaZ/vq2C5WeCgqaM+c5L4SmGc02MJ+9dS1L63tk2buWszuakQZqR7EAhsDTMUbYk6RDi
h3j/P7xOH8gFsHMdBsHAL2l1duTA3L4x4yefVQh9XZkPCIn8B6eNtKHFe40mvC49QYzdzDfRgth9
kIz3Br5vzgi/mJJrnPtn4nNmxf14JBfAqzrWx/HQKeK16LFhtoTUjnFRpXOf+zaHs3aIjasVDhm4
JIInRTIqQPVN03W5H50k+OUEhya7UHg01Ppyfpexn37pGBOxWB1x9tMFBhlb0nta4qou+AN9t1LY
5jdnfokXWRJLyvwJMGnfZDDC/Mrtz35iP21ZtIRqpyZ+LyVmvUMtr/RPsbbrCyhnEGp+jeMsP5lq
yHFb/5pA7xkmsn07CfMAGXWT+YrPfKbnSv0RZsiUwDiJ+33zvylDWuwatOnsaoBEk43i0ancSSgv
R+uNKpo1SIDixpk/G/nWTfxCYhvhKakccUvLAPKKHfmaP6y6Cu8CGBTRp/XCBLtN78O6qzBsdbYl
pkvnsyd+kOAVR+UoOHdSsEKkl+348QGEQmNrXa1pQA+J6Fhx0l9G9ZOcHWhvH6EFC+2ofBRgrSet
jqvjmuVbME4Qv7LdLubuFRizVxicmJZoW+ULbeyBnQwogPL6gbgLJtksovhImVar553ktn59J0LE
UqeKdlKDDxqGxRsdgEkGMr3v28jjdAhUhJoD1lMWpDD8HJytylWVpjutlAQj/+pqbbSgqFAiHlYp
jfegbqE+sbibOR2r6Im6sUH3Na0EuAVLh+GRL4xEHu5vJImDnW7AK3NVwF02Xhd+aEA6bUnv/cS5
KTWAffaoMRmYrpi0R9DCionLpJzvHX08Y/HsTFsWl3OuppvHjAMbPnp7jSmj3jp+jt2vHrtan/z0
vDVUH6A5USiJ/jz2pCUNCvbQzQlL76sSlMoT0bQOMNO4SV/NyLGo/yWYb4Ke8auYC/IcOwtR7FA8
vJS74V48gwJmO/sNqKMDBsIgteC1iNuDChylvWzktHHsTg3957P5Z3x2EGkNavH8coJ5+Gse/52R
DgE7Exllv2QZR1zyjXUfl8t/YpOwMgFTAbzu4e6jJI5ia+A4F37DI1JCqJeONcjfrM4jqWm9cWnO
7Rsz02AkPtjMpH3t1Og95FBgTLQdtu5yXSvOWKCPpd3HiGh71bjNxf317qxS0z5lp3uNl1Eq/pDF
95s4qlQr4whVNfkyJ5ctsu87oavY6acJTqHTwnIUTASo2GzWJ0JDjCmNEEKjwESb44daanS3ujIB
CaVQOcSTybBbFLQKfvEVAFka17P0wwFksbyXL80sSCIrFMvtUvlgdOWbUD96DDDRR2yLxvXRlCrZ
EpeKgyRdYZXpYxqKvlYMhe+TQEi0h4FP3+dzCh8R8c+z5w66+BubgxhgI4xY6gWigzlkyoOqsO+7
yzRw55E56YxUkVDIGfv6xC9ePzFRQRqDw9Amq7Q4gwcwJibvwklPmIcPgenU/W7Ogd4nQBCbM1+r
ySsJ0mW80u5SXfXnkgn4/4cfhDCJH6QZKqcgGI4W3YDHCBJbN5Loq49Y5QR9aWdP4hOltpAoHzUm
oqgfIiFCWXJIw3nMU9wDf4b7x8cjiQWlSHSTCQE8by7J2soqfHaHpWHrnq85Dtngl0We0hdfnGdm
iQ5qjTKgCqmFvvFyZGXEooMeRqcQNR7XOUjuXl/KAwO+XWhDWYxOtzeP50JCEHrL7k1iRVJCt0gu
ffPruY0m0lo+hfD7UA5vJ1DgwqqMyGeClXWUd2Hal8Fo97VOlOOFvxUetAkuS0AfWdP3jHmtE9e9
1kYRl8F1VBC70iC4W6rXU2UIbjilKytCm1RRWEcWFPnmdOAqzFz5EaYDht9HMo9A0GIrO6LvzVP7
tLjWEObQofV6duZZ1ZCWWmiI/K90s90muqK/LC5kkOHKnB9/KMN41QX+Cfw8XfS7QGntb2XGPpP9
ukf39y0aJv+rrwWmHqj1viEh3Ik5rg3SKyIjhedBMMBsWFQCOIQiLgxZW3VReZ2Zaydh57RijlBu
smiFXk5v77MkbiT8DQHzvcrSvriLFzdquSvvUJxGk20XFZradE5b5fQY4CPTlKONx/a11WRAWS7l
70Wd1T/eVq1ui2ETj9QLdjRyTBn83AeWA4k1XFvIKD2rKycojM5ZUVoaoHUqvc2dgkI3jsqInBYt
/p+KccdclbEW3DU7q8ytrMbM6pZyz3dqr7nszi6GfmXMIZA5ZsW1l7EEsQiq+ZsKFEEMVzRbdl/s
rhzelxW9jG/wa2Z8dmUxGUNQF6UGQNxaVYvWXFZ5UNoGLo2sJ5W+XpUI82sKICfMFsToDez5i9ea
sKafxKpCNHATNpVLHHQFN82Cz0gNNWrEvSR9em8+Fu30i5Nuw+hUWf3Ar5TIiaaDvTtKld/p7iu0
V72zwvUCzU9VUL9DL2C2BdNW/7GjpEYh2i4pHosWeTn6Bs6+wr5pDdxOrT2wD+3ZwMBxeLGBYaLE
zR233acJ3RXZRscXyTZ1jFmiT5ckXGso3gA1oSTEozrGuSWUq5aJrOIVwenqcDGjE4kR/2ZRXSSs
uiwliAtC0fgBnmuH/SR+mDJhelXc/ymf2KlQMLoxq34EAGH1dGM0KbCoKUzdPZCxoeDj7tSNhuhW
Nhld2suKF4ppPNldtstHczUFpXM/lsif+6ewE+uysiBq6QC9jCJmbuv5Odu26rj1EUcKlg5afp9G
EiXzJCIDOuk+qJIQN4SePUmeR0yx2kx/NLl8pSk8l/DhGF+3763SWlP9yRdFaxhyS0OePTnfZ5Hh
/EEb+0VBt08maPY2ulBcw73OZRdtw0ymyQ08zcJW/gLDHQe8NxFlhiN5LnjxQOvCfyYCliwY8b80
Eem2X2b4EfHCxpR8dgl4P3kXoudO0uC6YURbOHWh6PSFdoHxyNdxFaMEX8I4QNJJ2YGPYO1BW4xC
T8EvROXlNJDf7rx/pcof0kUqDjUpjF7M1hgVksloYFHRH3wkKmEDv19Fj8JApVjkanTtEX6oPCTs
4tLACPPpKEPd1H8bP8RrF+KXl/mQIbONPEd3QUIK8Zv08Sq3pUW32B+onq1K8h7T3gMmpcCSSlTQ
sg49keuSt56kssbBdlBHbDvB6d9wPgRJ5RdvS4qhLEQyBtpTGV03aFeGbj7KCOxOOccpmzzb0fry
ALB2U4qTWmnRvsqxlgHFMYAiPIfNRAUijUsAiPrbTKcIGlIs/ULEIkkocURq+Ps9WCL5X8hRsrbx
ZC4AKZaxkIG0IiTfhL+A0HOuw0XUFXPiN0Bh2mGSkc2EaKDJVmMPyn7F17YmGLJWjw7l/7BNw1gw
jyIPvH6mh61yLSkUbAjf6GcRHq9qSbtmgLQfxBpozM6CsV1MgqMtrGdXCbdF593VkipdaxCl73Gd
5Cb4FB3a1uS+/Gkg3fbnDVW9Gf+BBpscY4gfLF1QTr/P3hYqK+P+SMm9Z6VnkEmN8EfOtV2fMpt7
jbK6OFklzDLlxDq+ks+fG5vedakqjvccjNOPUmq5d4NqTbstUj/R6zUr0yFIVCf1VOcF5RlFnYw3
L8O41B2WvJnf8xigLkH9KTAnbRiCx5HRlz2ZDArdy4LLDaQ2t7vsxTktMSCDQJRYC7DVSnH7aRiA
qdQMmUJxeJfkSVCTTf3IwOAZ/5wiFCAUzDrYcN86K0f1Fk/PA0oquGtA6lWiCIJQDmfr7pbABvp4
96gFbEI5NZegUpKEkCGZZ5jSJHO0a5f07dBDdAMw/sjYQq9DMBL9XjedbG2r2l9veJtzT4o2A/lE
CXm5g4P25KWQtwGI01mOgtvI8qLxgsewckZ1g4xXn5eXXopSC0gAcbsCxtbnO8QaiaPQQaXhDDm+
C2pRO7QBtbVNMsvBC71juyGEBZsHF347bt5WpFJOh7IypQXL7DleES1dl55GeBp/bDPBP9HOzPVn
fm0Kgr7l7dG9mDp1dDaIYt3+bQjWxTiAhkvY24jOttJzPPsOLfNUpD/plOBgvb4eE0DKSm5E3sDa
EyFVd/lVrbLbyUwPtTMeD/DdPkVqTcRPCX2qtfcFa5CGKuZ03ysSzoQMC7F6QgHHaDy2M3zaVKsD
A3ZrzLI1qBCzKDSGeYOjDNDMa3bhrhAkHn5OPmBJlDrNevGC9F11AhelVRe0eCTcBNxY/tWXhcds
t4p005rzuQr3dnoEay6T2ITpCjHIIc6dIrSVocCJwUqdiuUMVaLyvEAynDS8Q7CE/A8F/zuI+EzU
zsAHyErvgzYO3rrnBl2DetuDmFcr6zCynW+jlUH6f+le8LetXBGnub70BvA4Rmwp/2WZEsXiJ4Xh
Flj8poz6OiE24E+dAsqTdRSSGR6GTq5X2lRaEy/zewMUol27tzanEKpDWn1E0i57kkv9vvcwIVVB
zoszBqniZ/zgVYwh1lOclT/bb798tpfxzvIDkSF0Ib93mNEX3eX8+lu6xiouyAsBy6x62Q6uDEb6
EZnDBwZKCJTN4ZfTWBW2jM9sNSc0bFj+29Uf8RBEEYJJwOhZ2U5qVa+LElAwSkmEQnC5O3pgpXbR
YF7D+O6pm/bXaytg0wfqUk9dSf3o6Q41obxIO+64ZRaxoD9hIhtMZQ9lNN0bsai2YT282MU7yHaY
XJ/ptwcfraxc8/xTRDGmXiywB2EFnbmMLv4GImNbHkhL1a44cWLYdZEaNW9mtR973/p7uQGK4ouI
7BKpPmUdT0FZYm+Z9w9m+XB0qte7KKBMdSUVJ53zlb7B6ZatfzUpsHAkpcU/9WGW1XZWFURp6cMy
061ZHNza0C4rasViL8j27dnFIvZ8mg3U7tkiWbmOblSufTgXbkiU4HK6gLfameAHxI9t6QwhKdVX
E18yqiMpRFrsk+O3S0Wy/BlFwOUrXTwMLyG/vGoTtoMdVI6XDhT4E8ZcX0xaPRQVaE+q3KkNjB49
PwA1Ndirn3ZDueCWzy2NPjEpvCbNZ8grFLqZ/6ElEPtd4dIjQiV/ccRCt8vEEzZc08tYiCvxeE0f
5swvvfwg75fc/JAmej4s74gWF3SKEKBh5eWOZNp37kq9KC1ohsd2270B+Ypab8pzdPQrsiaeI+K9
PC5QPeRupYkfqKDCxYtP8Wh6CPAgE9rtEXnmsBOy1/y9jp5jQmnKBw0A04CFJ/92NxwZSF5bieIW
OW4/Ox8TPzcJq1YkVd4Fb9kf2B8dPGG+mwA1GhU9uZNRkN7TynMBnacnY7RIr8FiLSyyUUZQATkI
qt4UM0rwmkVPUAd2+xzlcT/QlHpRb3bO5EzDqnK4dqlFYcS+Jq0kDThFkHZkc6DdYd2cSVQOncS/
JIveniy7oIVEtuM8sTN3iDXiEOwbbDLUfn7HyZgxBYDki6umgs8QGlAchBJo/m/LYt6IwRT2Ail3
B+ka6mIlpZneKlLhxR6cAtIvzK0gEjaMo7LEJBAjRjMG4T5BQuwa3ckMhJMK9K9A2U92SjjLDHzo
RLlxzIraPxlt26rLkcZV8e2rRyhO9ZLUSXUwWJq16KAbR5DNZfbmPh/Ynj2tHDBiUTAJid/Ihwec
jkb3vj16lSfsXHl3dVkYAo9EsghL+1QjNLs12Gh2C0zuoyW3lZA2YUp2wOs6ewAeKrWkHqx9H9qO
5jvW/0aEpMJD8R5cuZq91dbK9UBFrUpWwwyM+UyAVipE7OGmxerNuSaPoVyyrG4vti1rVcO3f8HV
TiuOjVrsflECm5o/XX2+dzbRP4cEf4WUdADnzQ6qm3koVskw0sW7KKIwYZg/e3CyeSv5Phb87luU
uMaCkmX7+tTQKeGhUAZryz64qRCdKJqsFSFp8nx8f3DKyf7MtQYwMkZSvyxbW0FM1W37LZYCSV6x
rgl/otvaHEWOoSxWpwHlWBehWm6pGg05q19LPDHnsYcc4+6lAdDxRnqOEk66zcIAZJWyIQ2XNr9X
t9SG+RiLn9MNtBz3XkzU/6WJsQaAfAzZZFCq5CN83RcXViwKv2vg5i0Bv2/DP/D6UrJrZuzRd4YH
G5gBxkUDdaPt9LeaRV0ApDgI4HeF4F857yxli+Mk5x0m9tY2P1ZSOuPmaNwotqnOcbXvlg1B0aW5
r35+ruZXaFU8EsPLkAKYMs41WvQeGW4m/MP2lwof5NTx1QBjBEjmVrT6PAAad23iNcFjkkc/Xjbv
A9IVe7hnXInoB/MLr4qsKAZjLFaalJF6SAfLxPP6liqIyftmlgLA/63TW2xyFzig9dQ+gEshqR3G
kz7CgM/uCLw+FlC4BN8uTWlFWTTmCjzdT5m2B7n1ojyXKdiU6phTXj/9XESMMejbYydgYhi9YPrJ
6TfmynwjEEnn89wis6pUexwNqD1eReRqI0E/H0irANxZaDECqZm2xXSmu36WMS9L0Dz01TMFY/vO
kVk3xBW0NSDV1/NX1G77+6555bxv41SbWJsOoimmVGJG8xjRLrxqWks8ipisR3H6USOrrhyQYdbr
+Kx2MvHs/FW/xRvjNS0NB4HGhFWwcFq0jCsNWVhnokkzWDaS49ZMtnlRPrLVydBxcN0FIRs9rBYC
ocHh8xugWWF+0Nn5QGXDl1KB2ElqTTKt2o/2o6gzRCNIEzu5BNz9txsKnOStYC/D96ZtmT0arIp4
Nr4/kMyW7D5dPMB3adFAy0ZiEZ8XlO0xJ1kMfSieflnJx7q6Cenzb+1jHkrnqVJSivTYMmz2+vL+
ljldrPIY4mcDXZUzBDC2L4jBkpZ56PJJhBuxPzYGTVVSg0ZkCrm33DAbg5Txsd3jK2UOXSYTZrM8
liLfc3xrTXdCac+cXKhvWPPxtXAajf7Cr/S7sR791ghxqkgD6tUWm2E+0t+HzOP0bHvOLXx3kBTL
0/rSKC6KGvCGq4j31akQF94Zyuygk9YgS9oAi1pTZLNDB92/Gc08D9MhiML9Uj+Kl/TdFhUhM9/d
i7/tbjd8FCu9PsyZoCGWH12rJNmm8+ZXVb+kNpkKVKg/N9SapUuJpix0D/PXN+lU90s5tqqTrgPS
xNQ5ALlVb70w+zpVGkWZmJAlCFuHs5U/fcHIxPOmBDbBAUKH+BInJtS8vf9xTiyfvCC+tV+bKp5A
ssJ5h2imTzIq3/Op8x+NcWzzmjB2rSyHP4UnfbFuLG0A9RjmD1Pncd+Fhn7v71TbEo+7L8Lm6MQL
WvQpVOxIAadvXXJBYtG1eVFxxOeLDGRxbsloSfc9bM8h61NG3mYXsy+2l0ze7KLQIl8+0Ag3mzYJ
WkitKAvLKyemYNBdO8xVFz+ednJit06ZpMkBE7NjA65ObEAbjNsUhEFsUxF44nUG2ipRuKKztgJo
VznJ8xqQwneHN3v1CBNyyoma6OIDzd9BMmR/T2psCVfQUbwouXat50eIeaAGg+JO5wFMEzr3fyda
UIWSPQaIKELHXcZKaKE3cJamVwrD8WeEnSoRVGbCVgF/NqODXetWz4zKuqUyBpifB1tk7WWbFHz1
YAP2+WFXKrfGVyfVrzIllthiNQIA87CLCeh8of5JaaW/nd763bTgNCuiW+tDz0JVREyk31HS1xnd
cPT4GtMILEGZDqme7fWAs3oQqB/uyLHVqY1GTrTnU0ZEbhVkSdg0xeWxwjofUFsoy1+cFP3ki3P5
JWHR6zzL8CAmxqAROWKGZIBUjKlKvOdEXXz1NvOSUzXD18VmKexMNg6PTGEsh+44L+hzgACknEgS
robzKoE67wKQq2emh5OYkI0mv/zok+TrriTB15z2Ct1fb9hh5e9eEV9y9DZnLdj/MADRrZu7z1bI
uzS0e+X+G4RbhAVgEf9OVOnY3rv8eU31wcYA/dfRNnwGzQnou8mNDj0hq0YAuILGkKE/mIapwD1w
z0e3eRS5YrnX2YPXw5rKmXUsYbFqHPvz6VTG0TNpkSbCupQunxM4cdPqGs2VtYC11GQol1LOT0Te
HTWoHKWimXPC5jwu+MArVvWxayHNCmE3Kci46HIet9ucDxG2Cob6DmJcVCeIFLLrIssR2KCSgAxW
v/X87smObwXp89OWom7i0eLfNeTST5mmgC3RPwFQ9EtBYn2rTRLQOtzkhteOOkJutaUJuNfLs8QK
l9OToocZ6DNSz7eJ2il5Fjzck4lXNBAEh/H2eX+ApM5zN7ImIbMczI65GvEiuqEksQcvwrB37JQV
PVkOHnvnNE1FMnHD90Z9Meur08cq1Rqix/1yMuYkycw7WHppR/Mmzx3yhfyQrdNMiTAopyIEW8OE
6QOVSEkS8M5aj+JA93r3BN6dEY6ez5LZ+KTNfy/wfb0tEyH9zqGDsS8crd5QtQnXbCj5aeSewhaS
7z3BlRg4QROE/nOkmhZGRB65rj7cpsRlT52qNbL8SKO0yEYUxYQW2IKQ7880AmjD1I2O5/auGp8Y
kLXsFviPCWaWwZ2s4ayF9ln04pRmEWBrMexyMuvnEkaIjiliIs10tANmQgMbvorQdl/lnrS6XlE1
ANLM5tniKRAZ+6nuyhHDieUyDgYQDd+pZ9+MEdSau5U5+e0aYYWcljqQBfULYr0ydZT9MyqQpjO+
aIW3ZeAtLpTOE5+PX7knPQpqIZMBc6CxCIiN4OlUf/9dz7xUW/JKqwad3d1mbCr1jXB5c4VpLCxU
BBejZoKSQee0e9x+oO2eKegG03zHAjYa7ATZaKtmTFUnziFfu7MjHAKg6l0RrW60bGNnCWL/wUh6
MCxEoLbJAqAH6+PEHoOUseCRHXRV6mzbIu2znVXNfKg2PAw5vpLDowryERimbz4LEXaeA0PkIsXi
9UdOqcXLn3CFByxi0P7V/mhUOqZj3Qy+uNS39CspKOu4gGOntxzxx6N8E3/fI/PAm5Pi+xqpzcgt
vCn3kRu37ukTgd2XSTa7JKXKoW4VDroTfUaUT3NT4gtao5oxMnZjcd3RTHHzcUxJ0rwXdydue60W
dCf4nbxsceJms4HX5VuSk+j9eg5ifBasSMyr7bq5cks4KN6TFvVRox8UffEFius5+zjKDPlXkILT
j/nEi1wNbtt91HvLqRy0TSG4oiJWSIpg+T6GiOnWeBmYq0LHAzA4xWEDjsvdIVzFkTa4koFM2rzn
wI13GPUAiDGChUrL9q/3wUtqVYFPOzjB7c1hKLcf5SH23LtU5MKpoXtBGpdpcccgzE7uiIVfhSQG
oDL7QSLNwO/bHKIe+2QnIPUuqygM76vZRSnlTU44sW7kIbCwTAGfaMSHPsNw/1KF2xM1FckxgQ1N
rl2tKJ6kcjRJ8ilWL2oftega/y2Kuw24lpYAO8bKWpw3fGSb1/zmoIW3c3WxZx1mWVh2bmOM3u+h
ZqOh4udvvcgMosp24fxOBVO6bqEYBq2IHB5vnKNSzzryrfA0WBaQMTsJuGP7Dv09w9yJe7CPl22L
mr2jQeG5ag2R670igSbHE8upCNT2UgFyefcTBaKT+B+KyVQBUrJ+t9FM+jKFxQ29VLrQmhgrttVl
lm9uls36sNIE8OC/Jjl/Neaeg7KLvUT86QYFZ2d7j98bvweklCAz7TINa8yeYwko6iCEIRYMn7Wg
q0TjCaai3U2vCN7gdWNRMIXWPcdbUHXyQ3AonZWf/EfkMc91l0umN+FsqzkBVzgRTBjJSXttKjTR
tjBcBcp50MNXChow0bvLWikJEL5iiXhUyxrBaMLwN8R/vve7CijX9Zn3hXleu7e11/SUcD1sbk17
dos5+x2izv5KGDMJK+XIQsoS4BZ6BxbRoHOiSGFvXc3nzh1FensFa8O5mRY7hXIHSc/oatuTfYk5
wEGmtqNyDWFP+VTwi+TmE3+T7g73aVYr26Bnj6B0wDgqPseFjL3oncggxxewOm+Ff8++wUaukyBn
/BiwaPTpO+W1mWERpAr0c+hsGasf0zoO8KOHwT6moCrOu3XwAZENVCZuX+pEKmrtkP2z4aH0aAYp
lRM+YeP49M1Q7EGnCKM5DJdTjgpZBFj5wPqqdYy1eSigxdGxImV9Ynklft9YMP+PpWswmK1l5zKO
WUQhGySyeDCvC/a0g7ksarqWjfnEzgGvJGIa3fsUj/b3A3hanpQ8oo/EHaeERfOUGD4nNaXWWwzw
eG6Mm/71dG0EBp1MWooRnoDYnkjTy19c0IZIOk1veegqbwWYF1uSpHYsjHa+QWTe7m7/dxUX/dV7
9k+9DJu5RAh4rsXIR4F/0md8H+kxjntzFFdNbJrW+w3uWAPSt4wouw5UT4Ze1a5UU4LP8ez6KYlt
3pRLyLmD06XiRhOATHrHXBbzseWijTvIp5FiXVh51tPlqNXLURkvbOxsFpbDsTnnAmhHIfehTZAY
H9EEmSEATLa45dKDykDOeXKWxNwQTgUAVsN3bDWWhfPQm6eQHEbLzsZiFaOZEEQGAx9S0vKsckSA
a2aeXneDu4IqGYokyUGJhPPMKIa7KKHxlQ4nOhQPeWVDNIy06FZ6KynNCDFIOwhdBZC9fN1tWzXe
VkHUspuvz77kGygY9fqVNUZnYDR9Z0R4WGvez2pRxkBgNFfjmaWYvV9pdwLhZehbiyYxwXt1WK4u
Tskv2U0M6MEV5HBAavaTtdeQPNbPToqpa6QwHzMr10tquTrfn/nuXl8jyAo5T7d11tOV01EL8Ja3
F2O61FAK0HsvcldoWqlyDKHf9eVlBIV8qlYkfr1d7Lnii2RV7I2YGA+VFiCgxHMN3ycro1t9xEAL
f9Y346DfWHNFyUdMB9K9BAI/+AXr1AxgDBm8FK0K6xx6EIBywHzUxR442pDt1KqqEFM01cOxCTMD
8z/kS4/9qQzJ8I3st0IrwCuumNt8e2efvDV4h0mp1MdSUJ7Wlm8VC7qrsMJNl/rIcu9P+rXrqyUB
Gs5f6ZqQUm6jbyjwXdyATlL12lck+PwBKxjIJ+KUErY3IZ+FnEFm4w3xiLBcto4PTrbr2J7VNXhe
+tpyL0F4S4BbxpyroxW46ZJJqrxonHlIrGQ8C4u/w8FROrf9+yKfQ3cd2am6I4N//zIijfycHCm6
pHyYs/eWDs0M3TUoqQ/4E93OWVudPuWexZgdY/Aua8OhwnPlVCGAlk50kRVP4WahXsc7plAqDta7
ujPxt+UbGb3U6BFSLdd5XRzHZbN4PddW3+YOO7dAyFb6kwSSg73DXDBzx1xRXpUVaJxXpTYff6k4
wEdJTNVcb1jyFWQExT3Cjxf1kPqE4DjXojw1n6fa3CVi0MHlwWkCYB1vqlMjYuCD8IRyhZqRdbHA
cIkjgSfZgGyawsAZSgYgQWBm2D6MEDIiqtdhW1K7KlWmERJzno9gT7PNCVBHolrDQJ5OjwcBQvS4
MyyFE73n58Nd/WaWAtqruKKPj+8Jg9uh8sZvF17WLiXKZ9puaR0CJwdB18V2psZGh+j9n+AS7Lsu
oWbl4gmIxtVX4szUwTIjO0v5CQSxpq/TBpWGbr+Ji7YiZlQgdI4RWbC47mfszZrqz9fIkqjvioQL
zem+Q56oqtRzdQIkpI7EuXAHomb5768oKljn+6jf6NSm8wkNoB3kcOk4k2tVKi5hZSunr6b/40EC
1ZmdESL72g9JLkwkylOVnP//4fA9251E4dqsZVF8mSFj1kpdCkluoO/hn92hykxbrOodA2WyoQd2
l09hls0aG/wbob4MzucUXhSk8FF/gx/+RJd72qLZeEAipwg2W3Yep516BQ/M6VZ3SzchlCQxp1ma
Ee54QN4kGpvbwfemdsVTk9gdgEFremK8Nx4K3hJ66/HUKuYwmOPFu4X8h+z/cCB3c6sidqxTWfB8
a3MeDFCcZgbEd+TDnJ+TSPBQEsA0SD2OF0tdTR9U7XcWRFGsQwIJFwyPXvB3bd9cYBLJi/+nRaS8
ItKIh9Jb/qQkYOQth1TsHGqQWZXhr/oUb19pqNHvPUBxXRQjOCeG3QxW/6YorlwG22UqTl4wIiK+
mvQajGjbq7f84GWpS+Pk/C+RryrFva2yuGJ6/lkJP4zUts2WxzpQAYr4Mpz6A4ifxIpfNKFT8JOU
70x5X6T5b+zOJodBTf9bZDU0vT/4KEBSVnQBFWQeGre4W1BrenfUP80gyRIsw3tHfgdfDMCTG78X
D+DFD/wbZxVFG3GqR4yT9gszhZSnrKAvTvuh40FsqoRvjzTGyKbPO9jkrJ/vSMqKZe1T44TZ+1i/
afEqqBV8ZwGqG8aW9D5tBirMX3aXmn5Nnf3RL4ViOx8XS3YEudGFGL5b60CRdWKqsDX/rdDcQQqf
RBpXaHFPBmqbIpmCSElK07e4MyEnPjnOGDJZGqFXNE8KIXjzR8oxGwZQL8UyZcmavpsY/kRnVnaA
tP/S4hOdvBSUKmSMLBFG1q202Lnob3fzCr4biEbgeHwzg4UlW41OmH/4m2/RUNqqHRMqtMq7pPQ2
AtgG60GB4kD+VD4XJD0ACFvbdme7r55VHpkKwEZnaVNb9mBSQgyaRaVavdHzp/PfTgnduIKEJnG2
CVE0ZIxy2CqcITmak6dOqXhN1hdSdyHcE37wGxyDD9oFs/VO8GZt+8SUJC+ER/TqAU7irJuTjFRG
jTjIrBVauUBhldHoMcjf/cc1h1veX+MBibfd5H7AfzH41yxYljFFsOHPvGO8UpaS3po0EGblvShk
bZfPvImSNISsl5Pd5trkavIjr7k12zDu7adJ9sdewhi7StS23sLAXXOmOfl36M3a0ncmT5a9w45k
+w1Q4Q36yyWGTFux/48q6JZEQPWpn9TzpQBBy77P4Ms3d/I6NiPU+GiYeIOqgBBY2DUsQHz4PH9G
5SkrLRgRtSv/uyB4JJ9MgeoQEUH6ApmlxUmGC4o8b3gq7ZuNPm5OoWF1XWCejF24ch3Lbq8ri9Sb
gn6dEYGtY64FT6i/T1QLEmeQj6ZGm6jwWifJiO+DebLSz+74h3gspBIZG3PUgRwR2FDa2UATmiPh
CgbLx5BoOS4ca1AwX1C7w/yHSfeh+QsYWecUCqpd4dXrw72g7QXMh6WqbVIDmQGePYtfE32ujfNh
HzATqI5jWzS7BZeJ0TER59FXj4hkMThhkpqmnS9VP8oH1Cfa2e2amasarVQazGf2b5Kc4PxiGNEG
QUaVIIks7f71bLYFwyKs4PWlEwl78QkX+GwSJlTQab5X2IB/bbhTak5+Q+1NeKWmyIr7gtesJTAR
U9Qcw/Tpm8kAbHJ79d7OVJMUkD468BTahx2h9snVAZ+VVEOHTV5ImNFNrduchsn2gOIjA+HVl/+l
n6I913iTZr6vsOu5A6t4HuqBAHiw0ETmZqEi2JhgXg1RFSfA2oEDY6wqZEx56DG2y0n0a9HOslYP
Ua7dxk2vBvoaPXLgEdNM++YKwEcNsnyM9Cvkvx7KArbG+UcFQcJ/DUJA9fi+nNp8wflt5Ag3lYU/
W706LvKxGHsJTcMkPkkIjtemy2167mRQ4DSAgNG0W07aEN6RaRjAX2J76NlF70HarGdrQM9JiJu5
oSezuh+yKifw0DLpPJvDEtWitSPld+MxxT83bCLSCg7RKye52g7Fh/LQ1vzGD02wwFyRc0mkXbqe
j9SDlzVcHQflrRlf49y+hnZVT8mbqVmqLh9FQ0tkf269JU7dIW2pTMFx8x3daomrMwxcBHur1Bb6
yThthomXEPGzzVT8LcZsoG5ceT+1VV8NnKAr/hMw0n0nq8kw3UU5fiKmF8/Gxm0hmP8+0kuD6ubX
p0QFqDrZvaxk8WNGowgfwtk/q2CigHQ9h/FeTt2dMchvLVVAuCWon1dwsxCBt+UNxqbChCV8uEpM
rKOi7oPDjo4p6y6VL3Knf9i6kEnSiNntv6/+yddx62tOyc+m1ThVYLGhx9Yj7uNoWLX0O/sfLuzi
Z9v3/cXDQHUk3uuGvi5t1Ij+oBE8TJTbD/PUpEEBu9vlCFGpSoA8PCh9KvmX8LiBbJlLqwhGNTx3
WYw7yYseJMQO+T/fX9hwIdtctYmpEq2iGJJISgDSmNLRPlmk1fbtQEAxQNqo+AkgYDL2AbA2ezer
FWHnqS+6xyRs+lt2hBkHHUs6R1R3feDq1m+LPg/tc0SLsIcQaHOzU7ihrOFPsa+hxqdYuJUP9HyZ
yu6kIVa0LT/JuCG01D0FA8TebKI3kys8u2IluzYbNqEh1Yld/pXa4zKELf+NSST9eWkWanjVw5LX
/xK6maYuK1AJCFRzVp7PaunH1IX0GsWgXklAJQgRemvdTfV5HQwduEgdGSYaaCAy7qDksPL+QKFU
9UvFeBj+dO6t39kKLnnBY32iZ9Io5kULBO9ubf66I6aD3p/ETehDDpks0d3tXu2bZm2NAQwkBfsh
uoWBqm8/Ek+w+wa0QIdvC+mTQgxUZei187I8PFynoJxasYnaSbPno+Vs3SG93dUo0r+i74ro1lHo
/b3qCKD8/pTI1SAGaJmp8TXrJBn0d9zyVNXwAV7ETg1UqKZaMewsfYmmJ6mKS94S4OncmMT0k5sb
RJvVUMGF+9i482mUqbfgVpBhK1QxiUspUUqmpq3ih4vKopMrhkAKheBnSM/bDW4rjH9chzBrFDqa
YkjnhSG2COTWZV6dBL/ju0+jKOCrlBBT9p2PuHSa14qEXAf8LVsxsFb2zypYni4z7Eb31nw2WHqp
db+up3A/EQFG7JKybxbsGiOr7UyOjym98phxdMiY5wkgiJskTQnmEqyMbEif9niazIGEBRO3AgdF
+wEr/VQoAzEtGdO3RJGq4az69hTxMb9o1fJPH9uU1Ln0MFxuiWWUZHAOtrQNdmyEBmz+47AjkUvG
BbRY1ZQZUDu9fDWIiSUTJmAkmPCkQ9gfkIpgLWHjy5BD3XDYcyQeAxPfM6ae3JS1BJD+TfusvO73
Vj0rXV1Ej7ofleKiwGQ3xnwPIJT7Pq1Bsgp9w0/0fpZJ6Xz9Dqjr+2+vaj/yTB48gCM/moJK7Kae
2gEZSKAS+fgfZWQETpagzQbPrGjfgDOAwjf5Po3pnZq1e5AND0FgcgsByPEUwLQRtEam/FdljGsu
IxeUAwJVD34ldo1YeUOVnI3si7f5B1njtJ1bgP0SU5hPRgi91eKJpmdAyy8DDMoZjyFj/34Uv/Mn
FrfCCNg1Op6LHQPRf1ZXTgzHARD4Zn4hVQG0Yj2rowfjTUKElY0ANJKQgLChcHFukkJVcV1uXMlV
MAXUo/Cxl87JipTtnbxqHVKnuSLg6DUeH/Kk6TI40qCIC3PHe1STYR38Hlpr0JoZE0OKeI+2/62U
HlyP+OfbzvSLzs9T5tYGySwZeO7tslPFRf9flarftJhZtexCm0tbrK46bDIibY1cqjQon3HqvWfj
+ack8AeAYxlSnha4uDfHUhV2QCfkz4ohOYwTN80q2xv88ACUPSbVNDKZX9IrLGKWp2j+ETivTAv+
8xQ2WXLU6mJOIjEz93fz+78g5jUTAzeJy/7T8Wn2qUI3GNtMRjQHaXwej26cdf4MARvfF+7dIo9/
LcB4ewyUiPpmHGWru4K83pURfMzFXJDEDsgoXdTXzvCoMVcd+g7+eM8rE6e0p+ny7ka3RWf6FO6c
XHr6Eunla2xbHA1fT12P55pB3tNKDcxo4jMj+hEN2vJrJwvvjeGk3w2WT4kE3w8dzErEQgcnt2bt
5jAfl6jxzkEh4XkNrSdoVCCCXyuT2Gqd6fUd3v4Npud8fnlP7fDBpf1106zxt60gFIPpsleZTU2K
bYZljsBIVjRq0n9/TWA3EbmJZOMnyxEAzVSU5Ou3phF2P2Ri1OwZ0fuF+bgmNco6+0CsAF6DvS5F
r4hdAVb3HKNJ/0rsAxqym5BA6Z8nHS3hP0Mkg6dW4GN0KysgzZBQ5G2AVJiFzPdB+56IFr2hyInm
J3ZauLm4D9kqVvorBzQ8x3L0dREbZfEKpQfihfzPqVIvvDx9qhy/kHphVgCfySo57XPfY8qdjutw
KXKsefRajaMs4cBevupAO6LrZpC4iTGAXT12dva7veF8kEG2teohqDUEQTsUwFxMXxvq1S4dDFBS
G4Kai4vYACmUZxebCBGqq35dJZqfDWazz2wFyVgm1eYgGjfTtVbQOZkYfXf1+VOjzmoVoXi0yoGK
qxqxbPyuMT8RZr34xw1A8UTMUbsE09XkYcAf9/NWu5tQ97z364HuWIWUkFUViHUeorKNlJ5IdZa7
rQQO7Aa1L4Dxs0wn9gBOJGiGRDGuoliZ3Qc9zFeCXe84y7mM1tGlO8rloYLOU6Lanm/6z75nLAuA
Tqijue6uMcTvip2iivRotjOVjpqCThrJFFaFQxr0UUGFYrWpqgD0oMNYisDm/1P2tHX9pVUKGrPW
lOSKMs7IZl32fHJZo5++SH+8ViRQVUkflRDJmcmpodaKCEphn1hcDST7ecgsJdUSY14qhNTK4slK
iT35T8G3qqQLlQX7l49S/4xVhf/DALFRN2x/2cvRNOe8UwUnZWSZcrlpzXT4d6ZzQHftOwRrLUsX
7nKS3IeSUHuphBj2QfY+SCtENC8fLdebV9v6VjVAPkeGeA1o9io+AM4g4v9jPD4MLW3LI9KoE2HZ
KEq497uOLRc0N2qEqeuGRL1KTNhqGg28JE0ITi2P4dKuFFXQuifeM8Py8wQLZnqYWy2L8q/lo8YS
tAF4BpbfTy2HqAynfVB40kmoezSE+9UAWnoBwWWFUKz0b7+HWNFsugRJJKb3xH+tDcGALTz8ih9Q
0UR8rlorINQcc6vgL1ISjqxQUVlxTsuqE4vIvpx5vsB5WEsW3lCzAqka+ywAi4qdQvgkk1abH0Bx
BTopWcrM003pJeR1qiKJ+LmOoJrJoO7GnB9URHmHCBjOTQtqfrPbyIyzjyod9nm8ImVJ+vYvFXw9
f4vsdFqTe7lQOQ3qyBdGsH0XwPXXXXejviRjBD/61m9uR55xXawSm2NBUVqDWCum08EQe/08kCcw
QTPle7fyZ9l/qRwpyQddH5hmNhc6MSYJPPehaFr0b1IxBXBdehp+JjjtIiPP9T6kQMFJkKGRzchX
L8MsXmOGHfYG3rB7x/c6uXfHwP7NaW3KIwoO6ppkV0xIoKC4uSPgKgzgySCyy8XcyPiQ9NqJ0x33
Lcq50Ir9fYE5dT12gz3dXEuzQOJzMsdv74nnyIs3nNjh3NqydVpnUdM/sOG+UqcmRtx10ul2VK5+
t7OCBeaGHh1QuB6+8H0xZ3ZsiljWEvekvLZK1bvIjwos1djwRMOIF7fnPPfgXu2teHaBugDihoxw
JWzlodRfsNAsToMAlxVFT6cGk9fZ4CSBThEKKLrK5v2eyvO8TwpKeezlrZ3Oxx35VOm920O/57sS
e/HrWCYKPERq2OJFUDYzrX3blllH7z3Q1IVZm7Dt3xnZJhv5/bJDGBP9lH7baS3/7GLgDbqgAemD
19gO9Srlbv81Nr5L0ulyX0uMS/rhQNzO86xeYMhI6VpLaA4oPY2nrKjY/jZeSSaOyQwW21LtCSel
AflHse0yJo06qKiLD209Y/1qSkz7IuvHct26zO93JMa5ReMaJSPpw0s1ZNmFqOigUCjeXPp+wbdM
OZXQQQiO1R17diFCS1bJmR8sOfMmHXwTZxCmhT+P2aA0EB6z9ttOKRU7DRLZHZazAN7jHg11suCK
zfFk6yram3X6lio4eA1p2Kxt5rvw6pwig7Mw7yMvOZq9CCKMQKD2E8DSLFO4x3sdy+RkFZTfT5AU
Qm6P+rIBdt5Z43c5v7r83wto9ga++0Lnny1eMaewMsPO3gWWPPCyT1Z70EX2qAElZDkEAEmaRxLy
xrjT9inKNHsrENvxoCEN0+Fb7v4v55HWgWVGkv19waWumoDLIi9jE1iDkLEPB9BH0UGXCvXpAtXx
/yHx4h0nlJUUmRdhS83c0WxgAd33HiXOHUDFwbDd/yOVJtPg3CVxiKrHzXoKK/7Cz8votdmv0roZ
VIkBDDBWCLjosAIpZNXhjM+FpgJyAgfFor0+f/7F+7LegpaXs+K+0DlcoXgPgWtq9mmgK5Gv3rZg
OXYHbkGK8zBPGd2KZt9mdgMDRGOf1BAjOhcyC67yoDEZLBEZZp54G1uCcqxEVqjqtvzQhhk4WorY
cvjoyK50PXBVTMLKGzirU/eJNuXjsaWhqbT5ZRSVj910GuJSRPhvizaCr49Yjk2qJ74fTCP3l1NK
E7nxZLIDC3yGTzOci6ezgWJGUEaKVXG2uaruAy5sS49yONaXhykaO16HlKRP4K42o7MTueEdBi9W
gKbC8zVR3ifgnKiuC81496KGoO8rdpy2gP+YDTBcmOHf2ImX1BgzDrJ7NqiKMkra+wH/fP17vbWP
LiV+NI3tFD4xRXMwKESM2FaNXrY52ps45nBlfAYBk8cqmg+JPdjOucYG7uOuCJlkc0c2ezdJUcP4
SQgb3sZAmaV1qvKWSgLpMi0uFPw/g/528G4QVLZuyldM6jaoJ+SDL+36dcCEbatHsjgqSnlZBL69
poCJAFhz5eYv9msZqnsPVW01Zq4/Er4PveIvoqFLyPlqf+SXe3D8W0HTcu7fPPMKJ0b6lteqHd1Z
Cvy2dG91648y7Paamqzym29o/ePlrco8aMLoK0q9JEIusXsQWxIf9S1UhepGYNwGX5BpkxY1GqMz
3+zsbH6/EKjga/MZi+JtZeA0ltjIwbNjnKoLBCTBB/90L4BcORHqXJ2OqWh5OUdl77uCyHCTBww9
k7puB8l/8jP4nv6kSEHQOznhpzmthDMamhqRU/mWbU9iyC8J1l63w0t9OvbMiNK+ODddN1OHH9Px
dfyTfSxPRDQ33s/WfDBaY+JFm1wvrXkKDX5tVFvdv7YZGNnFkDCFzhg+0sy+wMlmDa83SwqlwU+E
bTvoJMEBUpiGwp6aZSqo2+KG3g+mzz2M9V0FWnYMIfeVwcq5I/DdwfJNcJRNqRuCCuZwpDKBzhIB
M3NwbVCRNdBuGzd2FWrTJRUsE4w/o7rc+H01lG4KTZlT3J5sMjufO7piZ6gIWR8F/RfuwYL/N/l2
YwtJm6DyemQC53o+A0Rd7JWFSz9es7XEbVNPv7bXEImJCddBEz2gOAiJLNfM7tPP+qbH0bmmIumL
R9Rfa3z9pveT720qvcULVjiDvLDxdroslnYFPkMe+eHddl/eDl1JBX2Ho9aOapqb/z7ESuS5VrSc
TbbzqZhJCxI6C6HHo2U8xuCtsS5CfpFtfDc1Mte1cwobGoA72EdiRItYwSse8+RywV0eYHF61VOE
IVvZhx6JYi373K44538dMIyJn1APJGr4IC6Lw86vf+IOp2siYF06C8ne/wn5DAwlrTSaQRBMMFDO
vDWGjTJ81CIEPBQlQ+jMcdFfkg6wu0oLlZP35jw/D+KgChGYt2VBO6lP8krRnb14zah9hmzMDsYN
+rwQ1eObyjNhp4blzbFENm7vGHX8HE3PFjteTmr8s4vOawPfMkaaZAJ9nzYKHiFh/DryBRVhnaO9
Es5rW3O8Sedd54ibJCWzXMh8cVxYigK+RvYYqBeVf7HxDqz/Guz5+P8h3GOfEY1jESaD+K3htN1N
kvSJQ11PGFNSNmKrm1W6TZx9INcvjOX6xbP5dJwM0aS8k9nlOr+HacmNPTEPwfLAJmvDnAKVDwJs
KyF00l89AR9pif/w070Z9Igmc6rVFvnz8wauV/xyvqVvI3+DdxnKyqa6CuYBoLHbH33kio0mSsM9
0ytWYf34I1NqQsN+xOhg8Uz/IY5S86es47mASEMZzXMACKzGUdAiK1HMGVNjVBL3Pv5qPez0UL+u
sGwQa6BKS+HQQVUMmXnJHk0pQaRqAHhB74gV4TNDdMZ3QsbYKH62SUDFVryWReMHBdKFBRC+RTm4
XoRCg13Oh3sltXLo9PyMNgft2csm6X5oc24OlUKKFRIofU9Z6D+jbmqlF5Ck28ZD/3WOx7IPMZYU
EMxB0uMg9UXZjZ8RFZHPE9d+dRD2OONAolMi7DyGKkH1ZSiJXyPYINalCTH+v/igvRkoG3Wodu7L
+KzSakudk90yW3qirfq6UB2PJ4TZQWYd7ya8Qnl4Y34G+VgPld6m7SlOWgz9vIulacX15z5+1acN
urknB8qZL2ma+mDQlOwN/rlipys6dmZuZjI4N69qvOEKbj0QgIjH5TLtqHBtfirz0eRBAhmC6Vc+
HxxM2uNtBZSDWzNGklGckbjfo7kA391c6/onhDcouAQBlmdGwNgYQHHSMP4NtcXb9+idikirC4vN
XEsI/AjWFKMFMQx7FLDTsjtLYO91fpAxihfiCR2LL5Y5HaH9soHW/aAAGQXcF3KzI3xG7oHEw3w9
6mNw2Drkv8xseoO9e6WozD1BHX8Oy1JZ537FsdS1nAJ28wErujR8nY2UpzyRJHmc9dxtnYq6NNLb
3OhuB1mtPxuPxfwZ9BPTIzNJchrGCfJq/Okbmm1c/k1xcW2TwLvgaf+iJ7JF/J6pkgqTQUaxfsIP
YbMfLF9MMd6zvzdEMTD3FVuG7Y0uwmlBJlVOCliv4Jc2bERHhGywZClQvulZF/Hv2W2JKFZHsk9w
v4XuJcE1Fr0rje0wNbSgD537JS1HP3lAgwif5vpOhsKmC4fVp/a23F+yMvrG63G7yJ2d+Mx1FOdF
v1a4GSV7RbRuuG6u+arCMu+Gexq6fp8pvvyH45Dn818G+si5iaF2DrF3zsQq7VxIWNd6fcegPyI8
LCCzYV5F6VlgUt2eGe4xMuBdWUdtptM9ODT335AVPWSvZucpdl+KEK7ami+dRZLAwVspCDM7lElH
gaWNkHTa6A7ZbeaHSn0HAdOmaS36iyiEKZasz1URdYro/P1DrpZXHI/ySW0yHUONMyCSSERbmkwk
8mUc3DEeMS6iIqvSf02dTc9JyZfoppbTBBYX1MiDAH0lZR0Q8AtASF1jwxZwosWuOgCZNKTefn4M
4rb9urOljqaif0JA4mmApp/TVL8iXdnTZu3LJrhZPET/B/Pm7gskhgFRGA+xEseweTwnMXMlMKC2
GZCSffw1b92h6fSnZQirJMuKh/VsX5p4Lrh+4phMu7hJ+97+RV+W5i4jVT6+oeB2oRJX/HLCYnyn
qrjcHsWhOP1mkj0zh0+yVhSms/5B6zXb6lf3OCN1xurixE+M+yKnkqWMGqmAXJSsnIfHbpc82GmS
0aaa/gKxEP7bm4NfG9k+Eb1HS4QE0CYH00DI5jTorgst2PHaJBw3ncOekVj3nzUcL5WJmq9SFxEr
su3HL9mYeuweW/q6su03UwxWZcj1opnQBSCMWE8rxTUhjIj6I/TStSCwC5nodQPEilMVlpL52pZ5
YTA8Ga653eMJ66iXeU+PC4FRdJ/01cnS9IQ/lFb5NBulKiWq6Rh2cfgjkyChhNDxrUktnU2t/eYt
1t18pDW3IAhFvC02f1QTmDclm0Y+gQ/0xbpNBkqUxYBg9cvZeiOAU5mWVq618cZjNlLzdjjCPJ5c
CmUsyBeM5DJpZH7ygPUAHhk66zLZYAL/qxoh1sNUKz8Fw0h62Nohm0sr9snvnozFTHLXzNA1hXQa
+nY7RorwPsZZ9cBk+CcZj7VBIBc/3dX9dEFoTJos2eNTseY944wQGhdJ0HxQN3LTlsvtX1KB8S5w
+ge6T4zhFmsRRbLTTY6Qyq2RjaMTpBwr/tDLGTHyVHfzx+3T71sov8itjyq6NraMJc5vch9Aqo4P
sgO3aFZTEdW/u5L2Zxs/wDT3YdAWfeHdg5pM2s5tvfr5CHZNfNsC8nmHZx2j2HjiRE9YCl9W0h5M
Id82ZkAf4Dk7l0PqGX0TdqcWsDU0r9QuBmAf7BkWoqn62U+cIVGvCLq2ToZjWK2k3TZ1mA10Zgqy
HAHsXezYVQyCV6o5tartFmwEvZA7CQwqF4mXf1kwxhfGq/kEaIFzvEVxco8dHCE3cO+iNwtMErzk
oYaMqebiDKvPM/pmsjGrwlv9w24xoTdfuRB7hV2TxyPUY8MG/Ro/BCABhA6S+8EPqxTdYURMXvzI
TFyd3cZDqG6jl6avjL4l4yIQhm4hTwOsN/VLhnFrlPggqKH2EkAWovQbik7tKoSfpSAo4Gz5WcWh
pN83rWUQog0UcqIJOL55ScsT6OaInMP25Qska2Dyl8+dl+nOWx0cjqGp4zwiC6dcSNtBiRqW655f
/hi67G6lqGEGDnMXATQm+w1LXZDfRz9Yqjwl5XwIptYfp8ZCEk9jhka+6Iyt6WI3nOpuLRTyL6Jn
AneCCcwj3FdCTvhDfXMr2Pb0f9joW3oFFR+6JXHzrk0oM5+I3/18cmTHRE0paJB52iG4NBf6maWq
FpsyXdTwMhoovbzll9Wy0V6e1r/adPIMzkRxVKJhbs+0GwrCd4+toRofepiv/8iNaEe7kzdZu7vW
7Z/zdMgi4H0FODXTV4TmNYhRf4YXiOwfecR6Tq+HwiI5Uz3Gx/LEOf+l3WykCLukUvskOSvuLI3t
XujQtM0PFsu6M19fBINhIQjwiV1IR3CFG5kdK/TtNhlzsbyspetteVy4VAGXfBsbZ3wJRUf86n2y
S8+1e/xLAzuNP0hboIycjdVYPMx4nLqRa9EOHbUlXwAKClrAXl3wlI5bapbm7dqflyVVXEMJRw6u
TRsYwfmmKBF/6zTTsJo0UdUNuBhkACLPkCZ+XKP+GfpO1JoSVVBTitaVSiRe7vBd816LVms78/ZU
cZabGNOhRy6RZGhu3KGtGx+vYtAe2dJE1ic8XRbOb+EiDixA0uMDIFi0YC9Ca0mG0aktebOZ9cdH
Z/pUe5hr/v5GlMadJNAAqj0Vr+r034gcMd8XX1O8eI5aYVNb7V/IWNstZj7jP8NMIQzCgG+2GASm
I6n1lsnVXejlORJ8UlneG0mhkGLuGIg4VlIi5scnipYT0wEtFl6Y/h0tMaIhdzVjEAwzcPBsX2gR
NYjuS3FcTbPhSty96NFddVd1miujghEVSNN2jnWLqG6u6sV8R8x7tBIMQz416GMufq8oBMSXi+sc
q2TYe9OTvSZ/8am5isLkTc/V3teG6zi5NEZJ3DN2Axppqs3zVB5qTyIO6F2eio8b8tn1Ulc0+NXZ
J0gCfHotsQRwLyRMyM8iHgS5O62LqmBZbR/h/eRBbrZPYtXs7lgOl2DHk38fvzkD1RhTe+pwrGzu
8s9NTt5TeA7J/dmruAQX3t8E8RAP3VXo7EyJzKMhdTyXQa1QJZNtVErtiRHqRYMvo+6E1otnkxhQ
5E9/BDG7zvtHsF4VmuY332qHndZyT2Lb59vP1pv2pHgyrNM1JS3ZQnbG3Nl1WYcercCowTF2is6P
BCGU/yq5pFkyrZNVpuEyhShgbtNfna4qTgyuIaVypA1JL6fo67LQq+sbfjecRthJshgoGqIRXfVP
NIhXSHwmnC1fiRgLpA4o4UlFN42+CHRRWRHcKSKZP6lIfBOege6MNOyZOJCsd11veN9OgMNsCu4/
Oir1XmD+do/CLLPK1kJoltj8l0v7gKuAzy/YztGuuu9qIdSl9O45V4kri4gsdgtiwxbs7/IUc/WO
5NF6j6/2o9WYdSOCE4lHqsb8t3tliggDJX5JYMzTLTjvGkmCEeU4rufO/qMFCJ1LHeNlG/zryeEW
Z29zE3M8prPVYRRBf6LTfoRj8yCyIclowtyzlGwdoh0G1aeL8Fs0l62SpGo6d2Rj0H7MXHvbr1M5
m3Kaiojf6M/+CwCjUZsNMqXW5LAazHsAA3W3RPmX9FvWuQiOwR7pn/VI4OhPSXG0aQJPv4rBaR0O
xlG3LpHhcTsbQDW5rXDHcDdkJOKUxwEPo8UWjQehAtJOFjbTt7kuwMF6Ww8EXyo+wxeasG/9UawA
Enh9h6HnBVo+Yv1M38GHBl1B0WtSw37WalNyhOvh6UT/8AA/IVCoeKBhACHeCBkBmY5DP3HuurLr
QBpgoB65V0B7q7zEaygeSPF44Qj7pK0efZHv2jPMBmuLcP1m8RLaFn+nLtI6+qTT7iCYu9O8zSQP
B1mgvScC6TnB5TtbFT5tDSXRz0T/ac/2P0MnmWyyT8cj7GtSKn3GpRjgR647RtAnc8hk3TtI+6B3
MhN5j0ttj3e3cv2WXtW9Rxr6ZwnWXtQjpU08saAxaolCXVYJnQZUMXGtS4u/1/APMpv/F6Z2TG/X
8/hskoW5Yx8AlpSIJE1rPr0TPYXM4ugQv4G/A0b6oP1LTZQfjbJXjo6j0YULXWl2b4r15nO4CIXk
iJL09X8dVkbc4nzrJk/ajnwVlBdqpoymysL5znFWEHaa0g6WIwTLU3VrYaci58Xzn+EDzgvBTHnA
ZUj4L+yU/n1EzkfEgy8x9/0XlLzRTFrOVNOG7VQxcX+7p5nri+Y/qfACICFA8x2HitG20u2J69Gm
HC5/AM5UW4pHoaZWSrngloB3QpEY1e35TAPJvYfzpHWxENw4nn8KZa6xs3GN5Yxd1ggtcYQi1qOa
45tt9XK/uioBP8OyLEAyt6VUwgzlkuh2975LTvr/PJW+AgImE9FWDGmVWgvEToZE9YCfBNzUmx9d
rCwl5C3VjmaEHf/LxZtrqNV7SqWc4w2hdDV5r8/pCpwa2A/vM64CYKavNJV81d+glocT2C7enf8l
AeHyfxtWPmdGslzNcvHdJlpFlKdZooGxEpXxoRitLoGWcypdc/u5U+fb257a6CviKC0703+cNxMm
TkyY4mcFnmSa+FFQo3jsckif30g2PbNAs7zGfX1cYiKLWexsGt+n0t5yhGuBhzjPIRqGmYzSc7LW
81dKymwj7YtlI+Kf481upxIeszb+gFasQQLg3yqlYpUp6WPBFyBomSbnveKTL2+LAIpitLADWHcp
rUQUXwfxbliGpmAsYGehahL+c54wRv9/Pzyt7m6z3P5fwujQJS17H3VMZudB8qK53cQT4y/+78RD
VWNeMl672OUWpGVY+/xgDqY0kOFVYXjh/ey8JIprKe9mKIGncu8XMuY2awUVNF9UNa7tDlZuu4XR
HAOrK44alG3MYzTblAWmPRQXbby4is4CjbMddovqSFv1/vN9C+mBxZuBUzXAmFBpx7IT2ODZzxRh
5CV3lZ12I/n6KwxWRmCv2lz8ksBwqaGAuGPz8ATtszWPUrbPYgrdo/Cj3dNXG0FaKaf0Su/B97jt
CPIR03Tm6lkm6k/z52R7tEOHu1MTSDQ3t1PjfvLoyhPqOH+qo0/yyQOMl5iIEsRpPmJrMAONvM7F
WuoH2pGJNH+t5dNyKtvjhYj+dikKGvlR5TQPso8lXq60sOA2wN9P5+jiheH99EngiLqFtnAq5iSG
e2tQTn40bRP7qRtFTZbfgf+E0v5Q/WC5gZ3hGRWp8fva4IpPbJ5bD+OLCY7DGfBpC/8UT3J/k9/4
cL8kw9+zIHLdnLogyIeFEEVxmEhdx/Q6cja5JCPx1OaehsKUQt1W9t9XXb0kIX1HiVO0MXnQl2sp
6YOq04O1WRxigam3V5CgD48gyrBjkW/cx/h2PgI/dvvq/ShYEh/zJGMmQXdAoYHf2PxuLlPPjBQB
QUp6oLG72sH34XKhu4W/FLnZmFcef7+NgCQOCSiBlP1E55qFSUxiVBt6V53+6e4jwR8LcJeqHxjr
JZrQbvb/luuqCWBZ9W+qoo0ORDe19zpzZzTQagb7qO7GnTtLIYB7+6kC7wbtVDtqQI65TEHLvFpj
hYyxO/JN2NAcarmqspaTWL7TizZA8afI43A0TOjHKGnuG6Th9TfGgdxjFnfthjtDAsNDI6r/KsHF
5saZbPI72hRKGSiATB55pkziAgrLxACP9lSx/lgYe9itRJkzj8izH2pyisDMqoMvMQ9NqbT2XZyT
QqGq6+LlbuwVT1XGk1x6p4McF8D7UM55Kb6VesPewj6Z7cQmIqcQETzqF4mshYXVCsS7rnndyFYl
F/hgHcyQv2wAIgEl0BWQIXjigNO/kiYgzIPFgd+QnYrtH8CTcdgdcZs+M+xdiR9osFQH0P9vKiNT
nQOgmCgv6edrcs9qxIEB2kcEM3TgsYUuT2WD+bS7vuUSP3ikmyIrGLZGim78Zk5TBuFrcJ38+D9m
nhZa3m7Enx63Gk2aYqsRFxsZ0kGIAm0O/2VCDW/jb9Df3W3tPqIvJvfLQ9ccsVW/izWGojQYcpDZ
DGhdqRstjhGyHFAxDkDfV92KMuxipP5a6SFRJ0lnUZGKzcRyNmb9lmtsmVCN7k5HCVyxDOaL+rt+
gCa4aiak9z6voJUKkcdhAD4cglpkqCWX1ELvOWMqTSpYh0hg9qdXJ2XFWbcnVn1dSOcvbtgIvRwK
HCXqP2kh5uQIg7+h8NhACyMviVsd5C2ztZY+JBc0GDt9x0xW0CHMqLE4Qv07qr0s7e19zYpA/hEO
BNtYfop8z+MdtCJgbhuBs0BN/RaeubabaF5O+FZ+cV53U2oCPZUq6wNe1Fz3KLtExsQ8Rm9NJm55
eiQiS1ZTq8Q3iUEqXenyEaSIk1vKXujIXK9r42GO17Cb10D271ENwTnlTNW9DhWKv039UVLG+YUu
d2flZIt2bssGYUevHmUj+7DvBKSwUAQDBJKxkJglXpyE4IyxMoKSNKGGxMK5l11QAKQK30K7Mm7E
eU2WMN5oslZvbDDquZD98tOjbQ8t72hONCr+iwD1WPQ4zEXqxa2KjDuUtFVUtTXaM/BsdhrsJcgz
K0A2cG7IQNvGDBKzsGQKmSNSnIKZzvBQLg6OwJ7O8Sq2E8Iqu2FqKn7AgdOnsc82RAU7QMZDbAue
NmSR79mTZJz5MplR+tldjtHT7MzMSbkQXrMIS35YCsUW5bpcq01ABKTBA8lJOZdGvs4HtwbM+qzz
xIe845j7N6iTz6iufIyU3ZCKfTTwZTq/YgIjmP2mOXA7XceR9UBjED4Ws8fPaWIdANb1AIDsyHgp
PgXVL7SvECwJFMiExFUIlfrYpPexVaGHAkLKvaACThEAkABY6O0EDWkfizCljwadkBELluQjaJ02
HN2ABolQi12bbGOVXPTkiC6zbJe+q9vlu8G60e5pbAXBGFhAReMK7mz/l7E420qiJAC/Y6zkIxEM
ZXEovZpMBcYOgyKsNkft5jg/IQi022v5lnCQUmwymAhnYRFbwRgWdbS7KPRRfZnWg+buUacoQNEk
38qVCZ56RxtlGZyo/fqKULWGzqjig96YWMFpEryz9olcv3HOSDZIeBopmJUFBxLq4BeDJ2mSGCid
GbQcqZNLTNQP9SQ+ME9bfvv9wdM156I++IHNXXHDkVr6HOdCpon3WQIK3vFjdHIhIfDxIgRovbSF
90H1Tkai05fyCSz/vkjlRYuuv5V3S0W9Ka2U60j5kmM+yzEF8Z3lZxsbeX/ZYqv+YDZJk/IN9HKp
0VxOwko+2jVdWaR/ufYbVIK9ESC0z942N99C5uL06ysRQMi340Z+guwTLRAheWy9lzsb0iW4BVij
yV4IxMr+Qs6lYechNEhNtj9rPgP2g6IE+vSswXJD8odNoCQRCP/0nmfNEZgerA5lplfcgfkmYMYB
5a+tsNx4XDEC0PHxV7qR76jbKHDHvWqL1sT/uoLLPJ2cADSNd6+jjA8Qu79Qv3f/FiuppwVvz4dn
TTBAwyDr7WkgBTN9vI1kuJnsloitTq7RAN8Ift4PEe51Oqg5ienC+DWYwOhJoL0h2tsNMjrfBLm1
gFbLojm425DKAVrP7gzznqMk5JyzJLVESZYdhZNqmuxz0s6vVp+vcXmzIcXz5Nz0Ax7mqaMS7zB0
cMcStoCisJ/4cCOk8bHAFThrxPQL0UcZ5JVbBdde4ysWIFLjvO2H0h10XTvyCu4kftQkPrMhqD3E
HDuHKmQsRIh3rsNp/434LBaTRio2QNwuHVOn1lla0DdywwTIQJd6g4/eVGKJ3rbpL0DZgKevo2iA
5a0oI0bwl5IRK3qUCrUe1IWOKyHZiEIpJjacNSHQtFboOrmTtpxKrn5tsROrlIqLKx1BruXJtzVs
ZaFcvJV9SQIjUk2RfTLeiK5wTh1cMisAVhRjI/z6HsD69AiG5CFBN63N6CMUbWtwaejKT1G+K5kr
l55yZyVSDiuh5/ImErO6g36tFuVCl8vbDCtWCmgx4bMI394VF847P9yfUyRmwGVsUgMi3iap5Lbp
DQuCMrfdeZmUXxZG2U1so6OU7croUXys0nhokg+gbEBbrKv/FHchV/zeldwjUyeu1RAIleFCh9em
C4m5FUSgDtRHH0UJvJhEgvsNU5ExFGt9mINTeaY9jkSLYVZQ/fFqdydHhGSi4F2remJGda9kNpcH
O02IObwJQG27cPt3cjrZSZ9lvBBx2r6U3Ub5+8GvB0c972MzcaXy64QN4GPl4nlHaAkMcGMxDF//
0MzH7RfXnr5PbRs7oNMNp0rCfvAAjKNri8tQ94fz73EEnokro0Kp3bP2q8AMAXuYItho5Rk6kJvD
vHQ15ceKFFAc9PrV7kWI0e2PF1se60BBAR2VEWnQwnICzQ9StpXmWWVjdy3UjwBhViW4hVaALG3c
D1FPsZFNwDhQrfuJLGRJQgjC1fx2SRWQL03u6g+wFZQpfNbSNHEbVFRYmgQMpn7NanscsPZ0oQLG
ESYkZwWkHKKkIjQZeHg5cmlo37pfGZqzpI1K27HbUmbTOmDo3KZ7bMkiI2LZRCzpFz43h4m6mI90
kydJxUaQFVh8+M+i4v5IV9wMV5SvGUE64+Jki1kROQQsETLqxT5atiTum2USHZPliR6z2A9GcYiE
Y/7lFy7MHWSrrqqhJ/vYhK8n7U4uCmz2nTB8T4eV5PW9X91Ii09yDrDcj317uCuwTKakb9Ulwgme
PozW13HYXXdof3WY1wtGBjGFCq/lBFzVl3xbbSkj1rMp4NJruhXHhGVh+wnZTXaS0PpLjt8w7fl1
SVV5PlU6OZqZaQz/RcveCYgDbj4s8fUNfzFB232+V0yR2ELNKvBSVFgAUJ6OEn8h9FVsEsBUv1B3
jBOZpkt1NRA1aQTtjflcEcgNFv0qnHA2Anuvk5+lT28rt1yTGB0kGN7Q463ApP/I6deSJ5J6ZA5a
aaLoGa2DaTaMxtglUDOxOK+/lsujkrEEUgXdS5/hZhh1DkCSfg+8gg/oLYHZ4QlysxJfKNOujOR0
d8cxE0UmwlzQsE1tW34UfQ+oNJ1qDZBs8UaXZzM0MRY+flXppiXsxgTakkf2dJoM8JPtYuRCU5Ir
kkznr5lbRlVEbTo514N17s6KhL2kE+DMv7nc5rBXRW0m3KC0TDGB5aZHdZKG70EqA+7v/0h+4TIy
f5WlGuC4gZbfpat5Qdw6dNTKAF9nSCzFVuQnj1uEEY/w5k+6QodgjbIuvcUsoJJjpX/brP1irxYq
iudHvalxkdvypRkQNxv1LBgG+RNuJ49DeAPObfIrA+5zaDbWM6dt0xwGnm6vlS45QZhuZOnWNVcD
WXg5APP/viwFjaQhNfbrfpsdqFehSRzNqV2KV41zOa9/8joRonbtAPM3+d5XMRbtpD+ggh3zASBy
5x2N1TAOMUAv1EZxh+XJIWUlIBoRK9RX1oyBpclclB1yDFYh/oLPzpd+vhm1PK6FSOboGx428uHP
NgtkQiBaoJ7YsvlB1+r1qXPuXVElDelEgxxFUGMVsOdDiDaL1JKU9zG7d4aZengmLFL5dvYVBW+L
e52DF9DLCsgrrCnFFFEx0Mv5Q2qj7H7Ls99gD7lvw+uaS7EHpGctzvIIPVF4ujk9A5MAspSN3Mqr
ihdkIjR8R+0hb1fmAN/dpAoGh3o9iewKaCUg+yt9BWeV7FYY3Z5s0869SUtj6+BueM/2QVBGhOae
Fo946/35XH66mfZRQBSiqlY+SawPUvRXpjuIu6oJFlawsAIEmKzDhTXuRM1bu4YzdqocQGysmpiE
+8dTnyBWNwsar/V6bVLtC4JbfKy+9qKDCL1lPxEuRXdDVmzrXUqe9JOLMHSgeCRnZAgMxhZMTEG7
AQw2P3CEBmtNuXWKNbxLEaN4CnTiGTLLYxebfCegUU08tZ659w4HPJg8cLv0WmL0Qw8w7bU3kMgK
8DvXakOSylWuaSl8vbLyYH9P35P4kT4Msa/27693z9TbWZqrSedeGo3tbQAznb2R85Iil8pm8ibU
I98Ys9flvV/jF/4qlgVYt9RpcFdCMHeaikODs2yY5aCuORekaaJF0SuZamCfw5lRaUhK0OfHD5RV
Cl99QxHyFzSsJS6l96OnmF9ej6Cpax3d+oK1fZQbWM3UXQLYk/vtUX8dswGt5+pF1Pw+J91rppU2
JU7XV1yMRcoZEtLCsK+Ynck4fm6MKJS7WckAraYagZcXzTFjKyFzVum7jFCanT+I8vXSG+CSO4of
X7Wo3N5UIUZjs/ZY0UJQOb08gow/MsZXG8D/hetyvcP5Wa6SKxyrPCsxDzmvY8a9RG4Mhfq3JH8F
I+XYP87IenlI3EGk5vqQhU8C648EERJ3GBxaue4kaPYH6+SPxe9ulLvxtfvvIp5Q7357bWFpYoR7
czDo9n9GdG3rk4Ouogo0tgnhytOFd7Xgo29Jj0WWqD9S0uCakHJCyTGEKhuydvW6ll57npOzMyY1
qOLb8BPxJ9oVs3EP6FHSHDZ5O98McSE6xEJVP7NJKPbH9cz8Da0FwtRR+J4j49zA1NE+ewWqyYlX
jH0em+Rboj6MOfL+5Yt5WYtL46/4FQhtCM+BCTwhpBrpjaCteZHCuIB6ZcUCBR99QjFpavhQspQn
70FuXPlPMch8ge+EoxQDgX8BLMSpEw1p3+MZxpWexEftag1sOd+yi1TNw2KxjrWuB5XPBk/Mdnga
8GBqNrrS6skdja801PEh3DOk+UKIf79MPTgBW3IQWQ0Q5fQvXt/FaW3Sa3hhfp3THf5vyNp7dyec
ToNyI13gy0OquBSh/TzcP79xbd22zncA4fHXbwyrV9MagqXJ/iGCGUJa3UVpMtk/zy+lwHC8wiAE
B/nPKWY+ak6oIukp0jekKcD05DCaCx1/zwR0aYrK5DSEnlapFLOTfWJRi3jTP/y+5q6hi3PGEjjz
Erptpb1mSeU3TV/t4PDgTTcXDZZMgIrWeStVuVPruCb6ggnfH56QigTqS3cJaG5FX5iVWUbqrtfP
2D32HykeGl6KCKoALHVB9Xyv/Nm8KnPZXiKZHmVdo+14JyVL2wjJcfCDpGeGU+axR28pcVbDr6WS
oGPJyAWL+vqzQ18BwJql1EhdUSt0maBvpjpf5EcCLIieffhXr6nTFDz1hx1TkAMSgoaLmG3Avs8n
vJKimYS66A0v0nLYLj72Lqyvm+mLXe8VBiE5tUuy+VR+KF0UE6eO9s4u+LSz+oz+TUkIUyRYiiqp
PAbR+JLTGXidnAJiMNB8XAx7WAisITm6kSl3cREITpJnDHwRxFdOAta6ADme7av8vFtJB4huHKfy
UHjILlF/2CigQ0XqRY33wolj9P7NrYV5TjtU/2B1cMsL9DyaCk4naR1fzt1CfF/6Fre0CY9788Ra
zgcY/eHSCZTuiZg7Py+lBHnhTny33T0eR+63xIpenfNlRq5oIZUEUM9io8aKl531IJRNpaKZa9XT
AM3FwUBDmiOGatTsbfDeImouVaEzvNc2KfseH7OISE6pge6GPkP14YqcYAHtzdWWDgHLTVAvBOVt
uvTCzot4gXw108o4cTtbJ+8KUmVICGrHvzN6z0x2X1SpNV74ZGrFCb6EVgu+Y2zFNFl9xpTro0yL
6WwfwuNjFtofrfWK97TQhgvmUVkNublkX5nQ0KhukEBHHMjxmgabTkZDk06ZUL1ZehA1NBoT4mJY
GrlQP7kLaTDLbrLT9abvljo3PN/GxPxbHBW4UhEJ5LxR6+r5WsrlCvCkdZesIXc0k15pPQy7gKEk
QfwfO132EKHOZ6qo7aXGMnT7pdugXNseGVPTc6+kHwzu041pCqn7oNsqsuFfDeEIc/ej7jxah4W6
3lMjIKQKc+2IbKCZEXutKr+FMy3u6QA3XN5SJOZg50ts6771a1Vc3w6hsqQDHTGyCtOzFxsf0JJA
Flc/SDyRn1mKaZl4+fB4xldDAEjgNjKLHLhlz+yy+gngp0RaklZv+cQzaaD8XGz89KPavp1WJ0j7
rdpptROI+DucsUTB1ktNyvjOFa/lSEO3GaHKNzOD31pY9FgY/gY09eNWn0Fr+PFZfDvPoYAE7QvO
DYObj5FRoSfr8iN2KLiZKknLoZwBA4dwUr2slZSXPVHC1iu3gRlH0YBVVX0HSwTeU5mFHfdj9bZo
X9Lr/TMB51wt6cTUvGTyFVlboDc1YDMrEFy7ILVg+JbkC72zEM5TQOLkekqBu9P0Z3gdbTm5JpQj
RaveYuoK+oSq04+sQqT7beSCsOBASp70KGyr1rCnpG3Pcy7kyH00OX9/Jn0WBTXIJtyaUm0NuZ30
EfnO3KEIvD0BuN6WqFvmoCmGbXl+cmj8vD/D3FF+5wxYxnLDRCR3HEKcZhBfRnXB196O/RKxo2kf
CuTuO9+cuO2qkeZZWwHfPFSTYCBAaN+UYGRmYjVUZGV6FPgqQhiybTUgkZihU3EzzyfnkABYPzdg
C/E/+e+puyVzR/WCIPISTKtBj27Em53L2PnJAzdshyWbXjIwdE+WHVUuQ8TDWRberrmS/ThyZrWe
NxCMUwohm/aGWgyW6oySRUEvQpaQoZOM0+Ihy8pUsPR841YCTLsqcP2dze692CK5TzAR5y68Kw9w
kqvCwyTjmeRCkvgGRZs/gsxD8JkQ09dH6jsdrXCmRMnRo5JZM+brey5QZxB7fmiGuKDmlS8N+ngm
OYGG0RrwvSG2uhwpCJMO4PA9WnrZIEFghc7J0W7msatKkmi+2JrCw6s3WNdkn7p2eSmg+KWwSs+9
M02MQ+WKlYs6juUzfd6WTMSPvbm1VZQS3OG33ixUktW3TXf6BuEgQaW3uQ2ueqy0QhCfJ6zrglZr
8o0hPEeOnHTnIGzDkxi+DCid9rJjKuA6QX/IviSslX1qB2ZRCFmgao//fZjbsoZDsYVeetOZYWE1
R3E/MOa1GGolldl121BQdz5R0fnywpKCdimrcqP3dt/fHBautx5DB5qC/S8jxUAnEJimPEc0BmBU
gV4bE8SdbVz8lfL0EUeHgJQqjcGHpBLu1IGw6hyva8IXnAjHPbWb0OfmS2wbzZyzwkri82ZfJV9t
/f9qkbcCicaml/EYBt7c0hh0GLCPJ8rr4UfZ1JjCV7cq/FlJscoEpdoi16tnyOpb7Ef+l3M/aXFR
aqSp4PsX0PMnB5gHf37bxOx3ov9opAKymZ/gtn7nGFpe4zD7mgEBp4cQPEi/stU8BGXssz3ufffF
/kPXBazIsk6zz+nCW0xR/C9AQBx97W9yR/V6A49sVKKPgkoXQb9A7NrXmCLqnlPdUeFwqzCGjugr
zTUiEZMb+Y1jcQfcEiAf9ZcPqDcC0xNwjzv+yZRVwlEu+JdjqBbvmD7pAACUM1o1zQ1t+bTDGZBP
D4qRq+69CiCCUzss8CHH4+ZfVW4tF61Oa1vInNGdFPSrjlrA73dKTpnR3YQ27zLo0fIyaN5E5J7I
YXVFfOJ0U+uG4gEOk4P2wbgVOwgPPU38IdHSzAAyMtAFC7zKiSIfldgS3TGNcBX8eB3T/wH5ajjg
AjjUTM7hnUYu5k8Sel6sFB4v1Z+3WXfNfi3ufmuHNyv8hT55NVeXHV60wQ9R5ZkAnBeFtDc4RzfJ
hFfTb5ZirmYAOvwfh1zN1mlVxRi8WDyZy8emT2PsFPaq0ThsTj4ide2QzGbc6D44+a02OxAaWK3P
I1c6KHI8FIOE36NoBVt2rZVLDaeRKAkywga4BAFsUkGouFiGeorL3jXzUNB7P1OG+/DaxfvdfHnX
6oiC7EokUv+IxmmBd0IKL9DU3uFfT7sc2jtwKEg1WJsE1Blhr6Wl8PrLarXg3CE6u4aizjQ8QLM9
2JbXZkNKM+VFucXWcge5+yXI2tO5f0hViBwk/uV1DNv+Rq6aw28VJHCNQaMBFFOAGRokKwvhsV65
NOm7/Xv73j5X8qPZC/0IKYdQNpt82S44jLin7a/IuzCJkhoYWq8IXl26uUT5RMwo1/q3p/FOxtFI
NbV6taGbvaNKaf6Is/SNKoINb2gejOMEVbCV+w0aL+XdCVfyGZzHwePLSBi9W0JU3JMlMgu9ARiI
mJYZIrh5fA2ut5/9VUUs6Q+eb3mRVFVzh7OmsuD9Gx83iBNQwh8KT5Q1QFfv2QOOdm0CGlwcPM9S
n/2Ptd30fzTfR1hL3m1gOSmbSzmgr/9j78alk2/QmAtMh333mrZunEoxrJdl4vVYLCw9j61M3272
tIDAxLuex8WhkZ5YqllEuwEw5yMq0i90MeMV0H0fy5ikg3Lx+A4djWvKg5UHPxNyafiYgpVEgf0u
S7FiYeYGMzOdEiC2VGW0LevIyFE8BkOV+uoG46cu+WhORMLEbDh4AWAI7OaiX8KMOn0EicdbtYuF
nDDKivBJOq7DTLe3rfMPFh++ae+Nfv9vc1IkY2ytoRr48e0Jh38EIsnZNvyeljRdWA3mlU9n6CPl
g+aW3TDszpEozJ46V0zICIErbT+yC2XrmyEkmiszUi08V2O4DvitBjOtx91v78mHRmxRwaKMQyNw
lRTIQuRnPsSXJ+7Te4TKfluXOHlO0q6EGtXSqfXB6nN4i90WkphQcqqAi/Z+0kn7R7B8lXSSvg5F
uFmOGAeuyMGfI/xwrhzuLz8ofr7cQDRNau77L2dYPNcPnHlmBB0ldGfhO7M9yc/PMXyiP8OntxH/
moNwpOn6BEy8vTJGChZa3jfu654Xc13wBN8p5/vFcRG32xqKcC/PCJrC4g9mEjYXvuck/nOZwNVZ
6LK6zpgN8A99j5TOf8ZZ0nPRI37ptkV6jqpRMJCsnAtqWb61RDf8ii90ROf1La9piAYdeMZ5f5oE
XQai9NMBLO6/uV79uhh9VNu0T7JyqaK292eTscWFF7H1wSuSpeYTlHavy4WdqReCMbpj9JT5UY1c
SSXvW93zM6z+NcDhOJB9TY6qOaMfLEwxT6/km3JyEpCXcyxJcdLQZKQmrduDJ9keFAp0COKZP/lb
PGzPbJ0RnT7+Qufb+Q6s4fNWCnsS3bvQL3jnzhC5b+S/ohhcdM91qs7KL7nnqfWMGBiuTLZauqLY
NRiZuUpGr0GIxDprFu9PT/uAtweliFkSKrQU9OQRz3len0YozlGqDQES61YlXT77cXV4naYYkjh5
XquPVIPihOdGahJz9Lqg+31MTBxZs1QhtAq+i3vYTX10LuHV2Dzexgch+/Lq+79FIEQSNCNGKrNO
52yicWGY46MlwA3jzeQ33Wzw9mKuxgPBUSY7bS+zYOs6E2g2d1JAg1zNJUtjNNk9EoKY1Ds3mBuV
5r1pOzpurpxW/o8eKoqgr8d2dCT0Q31yQM7ifEJvG+4G9zn4uE6oB1Epw8xKnTd0SHe/0lt6IxjD
bl9/tIMzkVZ2ti0nGl/dfgTBP+r+2vl0cyeMlffGndXml0M8zYfxxtkqhKDhaLABDdxk3agJJsKI
kGKe/omieYoHMHRVUAB411s7s9IzzTYTZHi7wEuPSQynik/5055/DRj7vEhJ4YMxWd6+QOmk0mzn
zgWG+x5ji88ZyyHTdIUFEpBVNNdr7yVC2t0qtg1+KmvPP8ZkZUy5wru7Wd1p9g5yhAjVj17TzkfM
zjwKw8pJaRujvc7VOHN3OZR7ikI/5gPx/DXtJMihG6xzgB+ADmYcYFn6MgfVx/Ki0DqD5UBKML+y
F13RIpFb61GhM+MWwG5iaOnTZmd+8kfob1jiuq0CSWvnCZJMkvrGMISVwJcaaA4IaSshx2RaazZ4
kSezQ7u4RraiAAfNJ6Ouq5mqZ6ZrtTVwxlKEbXNUeuzSvcQsZju7Xyxm9b4VSa2cxtDXBAFxwS2S
JChXxxFQmOnV8EvnLoMtZMmBBvpP13ygl0XRp8tA39uVUZmkY9Y9qUmU+PbIaWWNUJyqZ0UINe95
pErKT4wDWVvFuDyy7fHsKNZkNJ7q+MSC8iN04El8LlbUrqHAY4JqKE4NpStjVHqY+tRYSJdiDEEE
B+64LQROyBSoq4mk3jzMyNIJ0XC4hOdNcMg6PsUF1jzE2iBRxR41IQTm3zTgzpw36YChE+qBXWyF
ILsTGm+Irkz/WY/FSQ7GwUYEAIqnjjvKyJzFhdut2MrcQoWSHW8+R97lz+MUIxffUcx9vHwpy5U9
lJQcvBdUl2ZPx3QPtt6W75eMrYbUpQUViSldMI0sSdAdLgDP7pw+tfEI8d8rIuEcka8UDf/tyWgW
ZIM8QwZ/q4TYssOntXNVemhZMDS3UX2OPWsVg5zwP2rGVIorIdWXuMyuBkBaRFtrKSIUq1EMqPmF
ogtf77k8bXryFYYhvEBYyG2zUIe6C7Dr7N7C2kQkXBFdk/njITsLpd2aXbit3Z+Xnbapx8aXdshQ
z052NzkmRuIpLI37bG7VWyj4m07NDDpsCibgLTm80XI1qRHl/HmyH8HFZp9MslkrTDZ5kDLPaNYS
E0SGbTPimRB39NAUplP5IeJZw5Ee0wrm6+NYqHEleBwHG9Z/SuCABxegO10GHxfUasMlMEWO9hAV
15cBm92+Ptr9Cf9YGOy8L6YFN/4OR95XyRVZ8ph2u7Ow2nIxdOwbdKBI/AjmuU9J6yS+ONpB1JtJ
18g58uvJ78qaSAk/kUUfBGKDJG26afsxd6lRo+LUeqMwIT3dzmeRZsMbKwPhcgiISxLNDDYyfk7z
Gi4daS8kEDRL8kcMMRoURs9lAYRJtDasL5gnzcJ0/gWwXfogFqrnwtOQlnHIem1IHqNAR7169km6
RrHuND1XwUm9PyK//xbSaJ6sndllDCcIwPKXQQuuL0qoeCXia6Dp4VMNyppy/tI+VgkbEsQAyw+2
6aM9gK7KYhKavFkSlfhBvMPV/o0dz6J6E3ggrnEmQiswdGuVZ3FgS6p5abSVW4HBMDPuugSzCdZq
Kpn/u2zwrqJGVDQKkELxkit1Hq18Dch5LsSKbtdVZ3R6TJ4ETPm35UrP2O2pOHTAN7nas1igHo3J
Gfz5WR8ycVCte5KEpHRNrw4jTYxxnx7yIMIuOuKQ7x04D7VWJzS0nj/I0MUdRrf8dBPouJvhjjfg
Q3RHM4yJ1oP9bpOXlfSgDNFWLOfQVaCzdkWRh0D/9ZLSYc/If1X43vH2dJTlSyYsFALCFAdMXUfn
d4B1Ew/UqUwztbqX2En7LP64CyiY+DcFmsf66VkvVFzYIurcygzPL6Ts/HvqKNmGcHrdWzZFEhFV
Ayxh559kSpFkny55EgcHSnTEPUhc+4obG5qCXKcJMNZAvb/INlaCgeRrUxYo+P6VaDUaNZEjKsW0
bqVy64VQUvoy561x0HNcH6snaJPCQUG+6/7JL6rKXKuqSjCivD2xrMIjVeEMW+70ugTuvD8rHVzO
MLt4z9uZaiQ/daFj8TKe53F/x+mhu0XsayngDSAbZPuPWSnTN+ojulp+makeiO+SPziEnF4NwoYS
Q/Fs9agZNCrbS+PuPIMUakylk7UJxsJ25tRxJNkaOaozXgxMuE2Jd29zla9Q3uJ8l+Q5+tjn6z2f
SUE/gJDxZe9eEwWoCb3WGG2vkxReDaxOxxYPyQGuontgASpRHB5KeGogNtGE9+3dttlZpek/dgw/
Bvd3/TPuib66ZhhD5qRLOnrvAAy39JhU1a1rKTeChcGTd8Z+ioxXgkb66T0eqHTbjIQ+L+TspfR7
flp0uP0geiqL6lK6PxTIrEcsSlUS+Hj94mClhFxEIt3UPKQ+jzC1q8wiedL/LslVRNGdfK2WmR8X
Pl/ddxbrQCOY1wLDQJoJKFpfz4jrmH6Ue6JlE0FX7kTkVj6byvQs2LhgnDvXozceBKBN2CtTHtXu
eDiwD9CjmIb9UqDQYj1oQE6XFtRS9D4QtT4r2p45n3vyTI4hsG7vcJDoPR7xsUjbC5vUgM1J8B3M
Ng5qmkWvXT0Cl9PbYxe3kzGn2BJO4c0YQ2NOtf9eE4mCqT/bTN/hchoD/piMlM5Z1kJriA1/igl1
IrQOQOvc4EoDy19DRIxrboYLwKBOq8T7BZ9uOhaNIpVAfLvutYBhcuMMIciAgjgH2Ub0b6KISQgp
RmZLv5Kw7NfXXDp+v1SxgNzmy4oORlI44he9cxGp8RsO37WjQeAp3dlsI6xIF/pQO/xYG5GdcRHK
lqnMnEYNiA4fd+Rxd4lwnRVHFZ5zt8xf5yYMvr2esDtsAyLjvmWKPUXymFMY1zrOkUcPnSFL9hma
6dVtOoutINFEAEXvXAmRFTpQk04zz54fA2+Yq0lEduRC9kQ9ClYEB2KdFV7S5bgdv4wzv0ucMyhP
+hR8sevtJcNhuhXbOW/KPQNi8kHluNuLQ8vm631xWLIdZd16JSnfR1OEK96ptRWTIB2TUf2bIABz
Ge6kHLuesG1lsw3Mvor5l4JiqTxcWAT9weWctgSEna74DO6OFPhQxLiNSpC/uw0AJEXdJkTSzS5a
5Z3f4MjrhnYX5aNElZYuBUzMPQs3QmYx9i3d/Vv6lU8vl6Yy81be4wwKv50HZzTtzjSr6tbq/Est
hwHqNjUz1VAwQ7Eh4YmB3YusMcoCiZdhKKev703Wu9zVgEjg8AIC7hg4rwc8nwagfoNt3juOWVC+
02rVpBLFxgPOqsnEKYv16iy08jst0OGyIxJJX9XziuwPleFIWawP0tt6x/qPMIY8s8wrsBThpgNF
LLb8GoBPOVwFBfMYbygLYi56ZSDSSbrH17+Uz3u7HcyNVdpqiKF4ccxnCdH0NV2KgrTE3UTckd3X
vyyENqRPgPurqoztLZ3buMXCSnL/efEBAFHarmPFm/9FL7M/3Jx/CN8+3rfFVCHtAJaT9DmYgE2R
PwwXiIfWltdHcPI2XscGF7vtoGgWFcdm/CjXkQpTl9Urhz4qE1vbPKdqwH8r+f9SDfxLQT3j0ly1
BZ2rX3zhnKEBpz+fCb9J7gR8GYVcGvKONzvdSmV0u4se3pD+R9EP+gTlVukZLt2MSziZm195Hu1X
kA9tJlZm27FGA0vIw+yGh0MHHUfqDGiIEsMnANxqqXB6XALqb2nyDjGfoL2wSHZ7GbinTl0K5DhT
n/TyzckYAQwP67I6b0f5/d0VjnE65JT99yJcefRHXRxO23AQ5uZp0P7SfpvljX/7Q3TwtazFyccH
SiuGrxx3b4D4Nm/naRTHYVhIvKeQeHZM74mLrzvlgmTPRTJJ8+5Bmnn3YVRBWQNO4IA6WxsZIxfS
GPWa5lu3W2aq0weI2lElSr0aP27tJFzfoeeWBTBP99qDSAB6EwjuFCjutKo2ag2UcUsIj4vNyRy2
HcSxnkl4+IG+vKstpUZP+P2Xyx2F5oG7t8eR+Qe+dwd28XiQeOMVZYr5xV6oBJy3pFpR2RugC6o2
JzPDXf90cKcMeUCFpT5THBoduWQv0hbvkEs2YXpEGX6gZjm+iQxcycihO6zROgawCZMCnnrk7FKq
9Zg6qJRCOndUZ4cxQGobqR41Pxsxqg5BbveuuI+bAb9N1EmJhMMuNpQt+kcc6bmL16RcDfy2Purw
kXgKVkLc6vtujIlqblT1MaQpDEx+t1zrxhhJN8srGaLM2nWFB779Bn2/pbhChs1X0kpLyAqHEfgU
r0Ah2ODsjhp3DXeDr1mSZdLs4baqhEmyjyqD6lsjblhvmkeeJ7uLZd9/p8108ByI2EEavGhvEcR9
E5hB9zW2aZVWbp5pjYRY4GhuGzEwSq+jyU2W/SfkTbgQh5tqKQrg64t1evn//N3/cXBS4dO0gjbd
hNG+hmqR3qiPXBsWC678Agt327M8opDZpRUyWzRMExrY6XbIPhDTsd/nAOzQ2bRa4NdAJBY8Yjen
b2xixX/qZw8YG8PmaXozYFQcppTLoan6nafdjHc4eCLaVXeyJ66M5EicYNsalQb7JUNZyGkjuDPm
Ddhv2ZVVs9JgWKapo4LVGZ7UkouB9qwI6/KAb1k+I5Re/cPC3v8Slc3f1Dr225LqMSYPA5hwQ6IL
+xfCQUJisbZdBnDEwEYXTGdm5pmSv3Oqu6g+/DmfPQO4Nj2PPjssmm9lvHd29JDq/raNMKnTzeOB
mAwJsMQIooqE9NVFIZxvRoPDX0sdSam5IOlBjZQ+Ad0v0kM2eklFIC9zCeHUgApYq+QAIzbZtW/u
7/oh1vQYPFD50nnK8hJAZdSLMBc3gkYGwR8sEniyvSQrsZlgy1nkLMsc6VE/zmNyE9LmgieSXSwW
ciO1zWzT7JnbLX1pj1ZN5F4UK9ywVrnuMe7XFsdGpxhk3qaoEfXyS/zIq7NIGyuFIQliwO46itdK
IKe95terwKA8S80ZwRG3QP42H4zeqX34S8jMUhXpNTv3yEZUrhdTXzw9prrQDlie5FZyW8C+PHXs
xIIz965uFubqYywgN0HGVwrVuRpAzIxDSvvNoS5Ykw1Tunq9ljmTtjZMkaIzgRVW6LC/TSHZojK2
o6gik+cIGk0h0aCBKUoykpXEwFFD87MaO+mPBgEhjnq1D2n3wway4B2OMbi0s4ozl5rl1D6hoDSZ
6hFwiH8x/HZnhXYlUv4F/X0mLXsfQ5ih7PAfxRINbDveqm3tJrjYNw80P7mEcaQpaK2kPuFreJ7u
uUcXjMEtJzSXZkieT68cSnDHPPO9QGfiofRI+ZYHkxGp+SJbf8OYEOwZASh0D+nv5kxgbA2gwT9M
sqKBP0/H3VJR6UUQGKy/QaCwcj170+6TgS6nbWlEsgLgTLnGDotZls+OZY42eobGhJ5X1AZcM/I6
hjF2Ns7/+Gketq8lG1cbykpSldgQa8jGZCbf43wBZDXoSBgXTbswqWxwXlFiXjNUIG/XVjHw8Yg0
W9DKPN3QsNS0KiID2LWfF/FNFfIrw60aPg5icrM5epfikoT8iENWuVfKgRDhjJmXhZtVhcnCrBIp
pcgrO2ZzrgV+/FfwP1/lr1XNbDzRSt8u+QaJi0sd0FWF/R+ZwRSn7fGpJsJpYzd+fmNbsgD21DS9
wXCNzDXIKrJUPvB/EEy+ID9K2ZEbksgPL7OBJD5GOkAJzzR5wb03sol1GOfjKIHvCRtsvSKfgfEc
BcygNeN/xrgUuM0U0YC3gnzdZjDeyg8u4YYLZYylXY7nhQm8gZGgC/B7AVGJjxsJFIcGSwMPPNBx
JcLJdzhywj5jDMc2D6ZY1b9FXz58p4ksmFHlqBmIb9xHOweJ2ybfPWCcC4a6TCcDjPqsjZ99+RCs
ksow8Jxlca1T7rG36pa/kdr47KDOzEQzjFYUsn7GEIRj9k4C0ABvwkz7qFykoLBmqLvA+FAg/mob
bYMCwKnCN0x6IJk85xzQDTJUZ3VMvhBPIPz24Yqe+arVQqukY9trxzgy91XW5bj36j02613butAl
OnwkhhWPsi253lGUNBN5ypJmrhu0/bjU6kX0slwD3y0LxZhBUjIpbNSnk3ocvdA+aNhS9RWZ0sUS
yGgE+97G3/LKWLwjbS62gH8MMZsJASB/jAeln2tEpbeU6K86vBRBPE0gnvDxN3SRngrw3qiP190Y
wbY/eY1q9GPq0+BjguxG1hqb/qkIo+bxhhu2scguQOWohAhyizkrsyi7rvxsMpMutKJNfJL4DWey
qbEwKQp304QzEUVmrDN1DWtdfjuG2vpq7w9l3OkiIoJFpVInfBHtWiaTlBsVP1yD6kpf/axnr/9Z
I6fd87FLnunwearLdNhCU12vvh5Lsd93q459tYvuCP0GDL/DI44mogtx/TPtgq6sA4+yiG0gjcvS
DnIpVP3uNKA+4humil0pxyYeN/B/TBhKCLKXtv6264Rrvs3qWRJVWdTIegXKxtxENu8AJA+goUww
AlZOh974fSEWElhhtGjpAMYJAuyuOexf/1rvUH3EImnpLvWFX0aDs6/GoxzL8kF8IQw6LhFzyLNi
LlL4h6UxXVuZ+6JeAMzCdQroHEIRZCL21BrRXyqehBQMf1FoyhmgqC4iGQFC117hte+xrQwlngws
zh3sSCu67OtI9KAlj6MXzk7EiBVhhQTjJvEhOUqkSzwRha0vvecr9dcBsfLowbWC5wZc9Bru/tuN
5ELCx/RgdZQiTueXLxzPkhJzf7Bcywy6lihIzlz4LnP3hotSkGycIF0ETNGCDJNVfmA5NNp0w4pf
KqTfCSXlhC4oedekyADhwf8i6ONjnvQmagIk314kJv82t6jdrSYuTO8Z+qkF3G+W8MN/HeZ2WXZX
m4zuv9cYj0k90uMMJJD4CUhcpr9z1UhrqTVXnAs3QA7fPqK5823SZ652uHRBLmHtGIRxXdejze3x
KNk77AebNVE7NwA39Fl3SByd4iyHpdyf6pXKMYpPLJ/nxu8ZUlYk6HCWc7+Elnq2pVNqDIczsvW7
WpHZnU/ZkNskQfVfWcoGX/JelTACjHzJXjNOKyJkia4eH1r3ffGQDaJhG5EqVnKYNpZYm0eHGpdI
hjXccyv0FiXrmSRod9h+leAJ4V8yjM3E6Jsw7WPoEmM0oz8J1Dy7Tk5eFjN+sI6/rYKRTKedW1DE
sUlYng+LpwLc/10HdXRaSfXh9f6pRig/ucWuvsIoIf0MNG15n427mubjvybJbB7wpMTOMO0N6YBT
d1uIuPSKQY/bTy/EGamcKZgMr3DTElXHOCw/WkWhVTRB5TsTCgg2B221gWshjLwC3T7aTwuu4vDJ
gK0OAfScfZS1xO0UWQJMjYUb48DO76ooxna1BoDLsUFfHjietxGgIAikETfnDNla+xPvLxl0UVD2
syxJaqbltYnSZxy9YTk4R8It1wXbn4htkjMMYP4tk1ssYq/KsWAdKQNLx+9tkCZ41taFKZAfVTGR
p3f5IvURi4xsDFlLXnr1ZRvpyLyxbcc8XKSa+ZjKuHK+bdEBU7rSVlDEBmmw/jIk4SLMSGglvVRl
kkH39SdTgc7I5IL6vfFexwVBfOvFupW/KyM9Vj3hzPnHP8VEhi/gSVRXVh4/255EkzS55jAvlkew
apaNi8BCJ9NE9MUvYMYyC0RpvMMnp2BD67cfTen2FhR+tFCNujXLVVhTVNy485Z2w9EDkl8EDW/U
i+IOm+CPFd3U1QFNomLsyaqIuQ4bBtN1UQZW/kbk7vsgi8OXke/r2u1aNVFe91L3Fj+g2tekf4if
Ltsrcr8Qvrl/jFJFSxDYUO87bbFidgS9v3IMojX+/EcLdVPzR/kWgjY4YWMhN3rZ+t5Ehif5Eep7
KFdzt46pfMrRbIM/Pwb7yKGmdrvmxV/KogJo/fi3gbXxEDmw5Dud0vnU4SXt94jTYdf1eawsdolF
4N0qcd3TSkqhiclEsSfMRs+HcBDRZz4nDgbmTr3zbmCQBoTfed4RtdjRYUPuaa440966r1SSMnM7
kdooi85Gf9OAUZjqfXKWFUq/O87W3s1oSZlIyR4gmMRgMVwjjukwbGW+7OJxxjk+0/Y+65KYe5s/
AH7Yg69TkMnZTbh46yiq31lSb6+lzfFsdSeVXXJkZq1jX9ykKLsyLUPj9RRsQSjP9mTcsD0yNV5b
z38oqbwyC5eksvyStITz04SVoF90qOD69XhczZ53Wlih4EYj17gygGtwH4+ls6rq8Rai8NYRvekp
JATIbVv9lHGizg5b9yHpJZZYHSdufEu+/hgd4EULCdCNaDBH+q4OIMqq7vn7KesTDmcCV9Ys8Ihi
wPRq8ZJhZ2ndAvCwm4BVNkZfR1cw6ZnTkOqcDiuGTQG1SCTmtQkb64twbd8SCyNCO5inNBEWE0Eh
OLahRIEVrSz0kI014q56PyxXJWZI3Dz7FN//ch3d3FB5m9ahAQCxejD9/lnunU8rusZt8buNbl22
5wJyWwjxaws93tcrHrWmaauNBn6du/6RV6IBhV9f0tBmOWlaW7tv7+ovnZNRrMqCdjfwpgxRX0j2
WW4kyfTM+OLlGMIMXWWTBh6vOHKNfbLwo+ETq7aTe0JNKOC1s/YsCvno5a2eO2QSPV8ZZHDqpeGb
jlcuQdWmE0lxU/bJwIm+EcOto2NXgweTDNwVb7pmAhQ7EYzvvjH42GeFeqHuBrucUOEX1R1Qq7ex
VPziFKpCV3gM4nb5zSjPyEjDKeNe8EmKDMjIoHXHmsbdjOGFYCau2YsImY2iIrj+RHQhHpaAmS73
iwprwmt3II7W3wATKK1W+3usJe+HJv/SYI2O2W27kHGUZvBCRB9V+Lf1/Jvc9MIajSsLPFKfKeBT
ppjxku44KYbi+CIf9SEtYgUR3JlUVp1MziTXM8gjqHKQRnSF7fSbo9qOMtxmnUTNMFcWy1vjC8vt
HCrqJuTI6NHd4oFkn1xrOQeuFNiw1KRILlI/ECpoQ/co1hx0F6rSrGN2FeiOZDyDgWVxjSc3+zHO
G/m02BbkSmmeNGmb1df5cYpKfbg5vCNoVzbpijueiPCMpDFjA7qkFHkkcQ1OqqmZwhaO5ER/GWr/
4qCFiQGXFCUYxN97ivR36T4WpyapHU2VAGpgMpvbSSE+Wbd3JLJ9Bp5Xm5w6hgMKJIOWW/WaBaR7
Ms3KjVdlVt8f/fkEUk1AfA7Djl+pZTTJENantkAULr2JNhu9JdSLOzhhfbe8v1To4jtANYTmTUvM
QHqkLTKBn50QHIsVkWcpH1mqlEEGeAy+MHSYPgK9EiYh+zZE1/wGgkLjYb9QuqyR+UW8LNknayyB
+f0nHrfIHs8taTgG2sLDuGR8vvSDDv768z8oONZHT+Xx4dpBgdBbfnIHFhzgI14dw23LcRe0BT8Z
V8GSOq9yV63iDQ6XkJ2TYbKAHAlZIE3n54+WRJYPLfN7vDy9B8v/KGWt/WlE4I0mTO8iBceyAPjJ
gqM6znw+7/1jTPI90JgEaEQJeSFNDMiWmGZ/cIcwBO4BEStDQZXhO34BxjNDZh90cWptCj3wrncO
OEGSx+Dhw03tPawmiJq/f9HcphJHnh6qRMleLlEXOoKJaEFpKS0LPKHjTLiJz9HeRKeByDlVJntE
BKedMKZBkqffiOfKFsHENdEm6xH0YGmibLVFvwdM2cIZ6E4vY17+MGW3QhmBJuQQ9q/X3GSadydv
JiWZivIu9ywWUBfEBHWvmlTS7JY3WEIYS98kp9NS9bwnJ08yqC7So1IBgxna7FrkF2AhiXRKwOd4
1DRLyQNaSaNXCdd3s9TlkbejhMAK8E6cwDw1XX8G/QW1wX6/yrM0lyGeXOphyh79nzWO5h326PqN
IImOorxAzmQXVcHonBf6c0DSHi0eB+YWWuty8+NYWJ2gUkBV3j7ORcmolc3+EQk+sg+Qtb+nC11G
ZuWNSAoFq8o7SlK3WXM/83FCwRQwKnZFXEtGhvNq9wXQ2uBDtxCSffK8y3j32iMwHTm7wnP9M1m6
ReT37qRPwIJ5tyHAV9jMO4wurxcH4VSurtpTiFRkIAmE0zU2oAuGIjJPXPsjIeHDp6IKIHzLtxzn
IFCac/ZWueNJJuSTcx/jIF4xeoDrlctUe/NDcTnhfp94qbjSquwCcscWutAckc26KcFR079AmJE4
xiKYphxCOVRexqSqnExsf6L/xaobrCHZx0QErGGoheqe//gRzIcT5FpVdKjQQetiBxluGoJN7STy
uAGsYCRnLX5H1JUuNTlE0TdO1SmXEi0pa5Yyff1tjkfhlwgmeDwTj4CNOcN1kRdVatcZa32Ll62K
XMMnH2+c/upp4Vp3NKPjujKZxRs7egqoJU+Z4Ab+Hy0rEb70XjiPajNTRyPYuOeFB20OmqUirneb
ZdXa6jvBI4e1En8Y1EaHYBJ10ikUZOcdgWJb3lLeW8ywru0QClDGzxMDER54xbsE3i7AW6x3P2Fm
kafAZmyxVSVc7YHhGo/oebH2E/SHUbRfQ0PyJVTcj9pULa8Kd5mykYNimPW5cvaF2sR869PDWnng
yLWzbkw1/DC6wyfXs8jx+Jl/WQSAl7TXk95KPMFr2tCYZxl9lGfknoni7yfIVs3WdojK2oaNtgd1
p+1DJnWABo7xnoE77Rpwri68/F9GEKV7VEqk68HCgCtkv77WR0ohEbLvBZPhPAgoJCKVmv3O7hwd
BLu4GG9Y12lWmD+OzIA4LGqYhuZ3CcR1RBKr4nVmzk/JOh1r/TzTDS1VN1ig25eYPrcdtf/IzqOa
g/fALdrVGmxsudaS2Lp6neQG5VarRtmFPEX/6n6UXz5LdmgkD2GcaCr3gXj97RErgt87N+gktMOE
yDu663a77Nq0dahHZlnS2A9ZX7ksfs+/R6rUlLZ78aausS06QNI+gvwHZmHl3zvOekh64tdl/fRu
XiZDFh3YffPXZW2xuGyUk1szReQkBFCtpIaa6nc2XOsC3zAH7mdWwLMx29CbymyL3vVFPCvycg4J
1fdlOAG8/QdaFKbnttLltHx0Sf6QecN8/JCyN584nXtTyWkQRM8ejQZfP0O6n2dvmFdPsPHLUTbi
flYJWrt3n0YmgYX0X1mdfPUWVgikXKWMPEBLpsKASY/2Mjrhio1cqk+Ds+dEcXIxibVBg9bmRHAU
H24SjysO2mosz/3uIzEHZOnjwTm3zIEeUtl56yeJKczvku2lIGHhji2zrcIRKrTzAiOfVvSa+rGf
E4+J/S1zO5DSdksQrmz7XWf3HFt01fpDTl2JhPcXNMUri6Qo78mycMfdf/SVckdcVg0VR4qd3Ygm
tswhqZM+ed8BSB7RYq5GTYbosCR5px2uxy7jcOhaZ5ZiXzd7UHI8V047z/TmAnsjLTrvbM1x5H7J
1lIbhsfnwDIKVlWEmSUTuAGuDysW8+M+x1nUXX2lEmrrOidJ2/lZ2+fzSb+vUa7nw1BvnCNNC3W9
cQ8L1KJdtKZrtp8eGGsHbrkORMOyf7nB4+RIVesr95+kWuy+A/7o/8hmHyZFriG5X0qk53OPKtqV
4jioaHbgbo1r6isPDQXxwpVPL+th5TCBApw4KYeGQGJIttbW7/VkHpzV2zkIk2+zy9wj+C+9DQhQ
BQ1fD0/o2lc6CpjwRgbcNExZ0hbOpIqSmBPaupccNVJ2I0v4oNdw68MTkHKnNhIvCxeHLy6Ydm6U
tshgd450bq38s3gpWy9kSNYKeKOk4+69iV/0Tshh4gEw5YS5R3TcqGtVCAy7VJc19LVyYeC1vf4c
U1csiwgmaZj5ceovVNhieknR1xjs/A09fNJDXgDhFmeOQK/BdCpYWu490C+Jyo7n2Sij7wYE4v1D
MHSmYgZtOUZIV9LEGu6i2QUHpZXHFZxzBhZCxdp0G+J6m4/kdSfbsqVJ7v3qbAjn6Z0R3UMNL19c
urLOagatTuzTHuo77qZBVOkni4PeosC/tTMdw6LLkPJV48emJw+fpnfhXWxdqWKlOdIFGEPi+dXT
HqemXjJhcRFggxpQzQm71/9R1QhkiiW8RE4vPTzNSpzH64T32SxhPEk05oRKKWYMFq9Wsp9ASBi3
G7d+JMtfKLJhPzvN5sgyZI2jhxxNZ5e23hZ8s86rlsteeCh+loQ7R1wIZkwUZO+wFG6hooc805aP
/Tq4qm1GU8JS8Isvfz8CYiCf0OD/Q3bVyrPyAi+cXptVEROJCn2uwPiN0eX8xxbnN1TXrHWXs3pJ
LINZi8LJ4iUkUXyWcy+ZzuOOymGFvkyeVqjvyosLJFlCNEHu/aKrdE0TmlvRzkilmEq4jMQztc/n
7ilnzIR8V8kKHSIkgm40d4UjcIHrSwK2+cWoZ21HVcwhh8ua7SdE97f3ZWsylEj55lkUkPbRBE/b
bHLYRJR0Mob6uVfMICKVSeD2Db1TyzeBp7683A1bEOy7TCPLzB9fCjU5+UIEnl7/6XLIwGNvoAhn
Jpl19xS13qNu3p3KM9gibqi7cr0PDaW/RQQXUriOhV/MRFnszQ6th16BuziQvgsz7aNddStn/X7w
mYMX9Edft5Acr20PsbdRVSb/YFZkLd3HNE0NvS7POhzEqKHDJ9VYUkCOaVEPZlrECwk6EAlnZxVz
U7ANW9k2HCMQkH7b7wqT3KUrZj23c3P2KhmMby7kvGa8zK7UQxi8N4xBDjTVwO1c1Uvx6DxiGXIU
dupJ/rsoNmV742gdANxzG5kP5Qcnv5tC1SA9oimmb7gGSGIi9JrMD5aq4FGatNrXkZaXEoEaGh6Q
csMChmmFNPIDWySV3eop+BdDwiAwTLpXVUe7c0p0PRGfVCGlczFw3ctOn5wGVtVtUdnm+iheXiGY
9KFRExPNfhDnbZEdUwqW+/e1oVLM5jh0qi9zm2n7AVXiPFUxbuJMO98cIOvsyFcV74+uYeye0l9G
cN1oeFc9Zb/HxuDPIc3fzSpCwyPs6vOV63iwHxIF5SIPSePEP3I+cP5pWQbmu0EAeEcXFkzE9XQH
4DNjYU0FtgY5H6Bwi7SK+MF44pBg1Yn6XuFE/LqaMrURAC7+x9KdWoXWxhdxFlheHFqMIf3N5Oe8
GyEYGtIvbOq3v+bJArWFgieNqZzQ0EdmCvIxrCSNDec8piZwTJZFK5BRajq4vj2IwHbFksNvJ69h
1OVfS9VbYHuOMREACOM8u0t0Yr+SvoIu9b1BoZJTrAc2IjId7vhYB6xT9hYIrogX7njM5gVn5fB/
6wZjHw8kzFNnJnBZt1/birlrEEmu0yA87daBhhGD7G5jSl4voh69OPcly0VJnHDp1KdbQkUVc/ud
Ov0yTXKn/rvKRW9rPf9NCQS7ssCKCSe+0BTOpStq72fL90vy0ans6fD4kJ+z3isJpnbWPrK+U2lO
I/vcJ6FXVrN7IOK07G1A2od4EVkLgLzgKYUZu1AhvyF1Zs3MZtgymtP58bc2sge31BxReCvPtqwJ
cE1n51vRdKghu4omfU04CPhkU7jFvyneF/zOmUOleejvNqeF8DYuWUr+v6gGAmMtrhK1J/HaC+fc
CuQfLPp7uIs4Sjj6SUWQIFu5ANINNgoyi1KICGThHxPkh8L03cqlsqVtMgZbANd9EKm9iLs/J4e8
54e9VONLs7Pi3YcvWjkLJGGGZiJk7v6lMOpnOeZW+irS6UvveAyBNDTXP7NdIQos8Llhq6xD+rO3
161VUqgDxjzD4A/5MBhA54UbnWtQp+557S3aWB8qPDRWeC+Q+MnhOQseS9mteN087hVbERLxoxyJ
K16/lkAJjvMBSRvyeubgRpgAjye4JiP6F7hAS1REDdsrECh+pjcZDlM1DAzxQ5SgP0GxlbAgmTJo
ZmJXjRmLQ00ZoW1BpDdIzd3TNA9DskEDs+OsWL4gxdWnFEImFHEua85oT8iZKTxPerDqqR6gfSpr
YxRFCKCJxiYgHYWAgLkfPS8fRAqAT1ZJ2YSRCagg4XmJA9JbJq222MRRZitFcBxLMVimhCldfQpQ
alKV3E3BtUYQDrKdD29EpS0PgMx6ArpaRLZwMO29MeZy9cHdkq7RNLJO00l90g3WWMIMn1Ak1pSq
G5r0mJFSpYNkKgtXWK5Qg/80rhUGGGgfgLqmGFcq3f693YxJ/ZcbPdqRTCvSbKgqBFpPNK2+p/sv
QYujHnOhohDeF/mkkZqDktAouXS7ShlMYeNlANfjRQDK9GRx27i3xeQKD7Eqi3d6BABJPAK5qcS8
XzxybI/q8ilAa95HMBzNZrC2zlbVn9TP2EmqmeIEYtYiZSvanoh6XpgWQo4raZa9gabbh2kQzShP
S5fYZkmUhCHGIMrYca8HYUgEsAo4L+eSc5iGlk73Vx/O2BjBemt5VIVXG8mrbIRq0ZxNjORq6493
YdSodlJz7Z9gtrfmm62zyCNN8tAnl00vNQwS6nyOUiOFtqo6nn7Ivh86kg3+R2sUiACwhu3EwYBQ
enl3egRfH6L+W5LqEHDHiwF0kdLVU2FRY9jIp/nqx6hzqFcYlp9v0wKDZqnwsOhIkd3VhiAnwHIi
kccVNgAgxQOOXsCdBkzqMyIXkbHUZqJMNoLOZgWEj+sdgCZHW6nIRUhLmLVLHKioge7aaqnJEIJ4
9C9RL/b3QCVVdtQZbaeMG0IBORnyyTf3mAuOtYASPkIRXbjaM4a4XqKkOehnnpJ7ZpqJuK+K8nAn
4cdxesDqlhbzoptdl9el8vXoMN8Nte4VHA5sYbx78uauCiIb27kLWtKfySlr3v2P9cgb4eNT5gXP
bkbvdnnZqsABTe3UIo+3XBBCMNBh2xTbFbdOH9H1ihMxORrofIIMhA04jA/Pod2lzYc3etVt0hne
HsGmdWzRAfGifUJvyugEy31e5y1eFV3jbw/xzYUFfUgXFciYij9LBhZ2OOyyKjLEFQssFIM7J1a6
oanv5JBTdSSnN0VElK4UZ/U3G66mcB94HA8waLxdAFVdcZraECypTJZDONYeoIOSe0bmPCooOmxb
qmfo3xpEQoMsk7SehRVtY6PUQObStigXT6A4piAQWGc4k4d/cWwcaOMjECFx//b1m1kC+yH3fA0y
us67Qh/cZItd2iyyhPWk3D15v+6C5vYHmehX919osGZ+FRcJKVY4S2r3umQw6q4RWnTci9PyMcp1
ekuTEl/h72WlfK1hANnS9n7kr4JgsKyFH7sYL3UQsg7Wk625tN2wRjIhwgoDJleXenBS95aQ6eFz
qH+BPT/GATY1/Tu00eriLikUhZrLdhpcjS43/6/6z9e4+/LnTxFSXzhhnnQfae56sLwL2qR677Ju
HTua+nevt5mkhsi2GhGOzQMrLc2b+cl2nXrpR+qcOeAral7CJe2tD2RyduZcnnir9i47boZ4q3d4
ZE66rDk8ltfeO5ORovTKG+mUeQ8vSN+8D4/78aUxYWj12HNKIHpYi6lqHIdBkreGqWTCl4tWt8HI
o1y5GG4apVxSktOldlu2KQ5OpEGj96yJMOvMS9rQiDzlUBAPIMv8ThHLOjvqjT/VZOrlLglBCtA4
26zS07cOgSKPFdmVCoi0/8J6ta5MEXCuIpdAmUjeegPoxDeCKR2cPsFTmYmPOgXmrUt4+beSVequ
kn/RuYmNOL5G2mv50Xh0HmkVBj/pC1sGYuZmb25O/UrwylE/1ngLl5Qs0PtU/Q66XC8kqAFdeHxL
CogVt4a9nOrupvm1kfTzqj4XXiYdHj8nEBF3VeOiDmblQ2I+cLWyj07Rd2pYYPtX9NZZtfcxiHOD
o0W9RMxGUzUs7/1bS6Mwd8PxFGkBEjLiSlBAnQI6NfO+L38Gklgme6OPB+KZLdPxoeGIVOoQdonX
G4sOdksbfizRHQwQNdW24VfocE4InbGoF1M8a7FvIoDmbSMk0S+Qu5TTlwL40CpZIXbcifByQusY
cS98I0sKQzsbM5bsTvVL9kIvm1cuO3ZJF2N1Bt6GcQg8X3q41YqrCM8TB0F1yZ1XYO+R1RaoqAOq
SWDqG229PSmliZwizLgoKyVKYZHObAOLzFlj3vbDTKWCF7ITub6o1jS3NjhRgXbYBUBoC17lfTA5
U7WTYMM2xI6D6xlafNzam0LaxJDnIRxZAKYBO0pqH9/BqC4noEN9izKRA0VT80NLSmTDfHCmhbEJ
EWhM6krJG/a6gIPgIi3/LP/BXkwPL4p4OChBtTIuMJ4FPXEFRoSruKNnv7aHDCIMpIHkjQWIwx89
UGEuOxHC9p7wn/6Isf3lKrKBxciC0G9wbkeohIOy5XdFROZx9NgBTLCHF6wxTTPF50BpFcIAK+f8
+FWZd0rNUCiw1buRxc6IveiJicym+ByGGXBXyR12qlN35FTxz00XrUnfkcmTxYyo6eAwT5+D+Kxs
JrrSWjpvI06lDvk5gggqnPc87+qlxxGQy8fH9T/mYlm6sbp3T+5Oo4GibWclIP2IxDvd48Vp5o4Z
gTUf5aoi/zjAfIsW7Fly9lDsdVJHubDhPt+gAoXTKqlIX9cDjlltV4aJmRSTILiIqvNbYgfVzqY+
6L6dLfWG5bkb0dkLFUhMYC0aUHi07rA2PTUTRGxtR1zIuj4EWRSa/B8AkrjbGgfotgAsy9aZFtdf
1tZXUUQis8Xzj5T86yJA7ImrphF1jUsClJmP+bqkopQ3VElj7uJioLsfhQnCH4GhiLRuCvaejm5l
VSlMft+TxrQgo5fEVbIvzFdc8pqxXZ+eCroOooISSDWlhP3fhCB0x58oZ1trroLER7hS7yBbn4p9
WR4/sCzHOclzjWxWCF5c2M//SD/DIZMmWhg0p8MO75WJu4e3ujv5y0FiMAj14GboqIJ0/XgzOqC/
N576lkHqvkDc+76ngaLZGNM+v8AUu3sfiqlUgcxYHQwLzne558OhaU8W/V+AsBtqAtPx/O4oFoT+
I9sbVQJjOaQozcXVIkpnOob8hYWKYngUMSjkLzSd1wws3DTiJGS3Bpc2/cs14lQkGpx9WDehkp+5
gdQOQMTjYDA+6YXFXrVGfLeM59jWR4HFcW5DnlAqynO0ZyGLay4eVf3JJ6ImE4+z9wm1zZrYpy8Z
xSXJDm+0rbpy87wQi7SJMEs+Q5kE1OqUcogJUR1ZygUV8qS+vSVxNgvntctyyPmBnW5KUprddHh1
M1pRxNsF3EwBMLowNeeQvi89atLJOOPZ/Bo+UTdxNwCdXxWVRfYeJDC/3qB4h3ZTDZbO/xjrId7m
Zu0O5eImMp/tfG8MH2fvxBQPATmuF0dA4ubwp8GNj8s7LshClHYmX640gC7qdAV7iX76yeGzxcg8
p4ZfBY2DJteMNVHHuZIrS56Hv8usUVgKB97zKIPxGsFov0NawX9p+QiutA6BX2Yhv249oe1tr30O
iK4Ubtqy4EwiPw1VvhkaTp49YadYtdot1OJ+wvYJlmEQZhLBbNjtTfka1frWGfCywJCG1NlcU+t9
lXd4yzkiaQeX4KKn1QQPxj38ajiHZN3DcHHvwzUFipWx6TwYrYvtdo0R2jiaU9aRrhREZmVgHMpJ
iL8XhAZHbuPjYYDLtY6fDCh5GvESdQqusBdbyrlp0OJhbv8QGlASuZmgief2vkCNg0ph8jTieOUb
kwpTpDSVkulO6VZfSyUc5SdJaJBfzVFZqn6hukQPwqV49ZgzTGHL/aKkR8PzW+WeR6c34w+Be55U
7npu3/cstUVJvng8b+TljPI1dKN2AycigePsuiE2BbEBgJaZknMOL83Xczg8TbQjxmsVTc/JEcoF
9Xx0tuLkKp6YMfs/VZkO1bWRPKXR/DYjVHzn1aRMcpGTi7LaYzUSRgIC9tNw1hkDqtGPTCuiKcDs
cVpaKMLW5YiaZp+nvqt6AZLqfiAMziEHyqElUfS2dYohVAWFGelQbOaSuzIaSpknsLaG/prXhh8Y
tqmt3bNKNpmLn1ZQ36T4vA/TjHexnwf4Knnu/QNqvi/PMhd+eCmJqiHlPMw5Oo55DpMDy4dMoAim
vMIhUcrNRbTGGr8OUI7I0PjOrrRKouyT+7BZK1GE8I898TwGhTaQYMcWCHup5aKQuQ3IPGtTxc63
GWUkWHZKezf3MLHsJd75rM+BASO4qwmty1L30S1pATfciYrlxpP1y8/RBGiLKPwoL/zAOUuCeWMg
j5GK0SPe0alhpuY+gEhDA5pCm3v7MOlBl6RkU4u031oMzOk3eteS0k0fGOpLQvAn2zGzsygT0qye
T5RiI196NwP4mWPQeNYyXO89QHobHbWGB+YJxOCs+exiksK1TmS39+GiGk+R253IUUEl0mJZYNPq
/9D0sa4hC6t3p5u1Bz9AFypoUuT1VLBUcTTC0/bkp0MVv9E+t9m28aQUHPwOAQBVBESlOEAs3r8A
6ZYsHCyrjbkygK++9OvsLqEOg2dPjbZdJhlPitNR3OzNX/nWddOxjfzA2m5QTQC4m1jTlIwWb33r
RRvI2RlNXrmOImwSKhC/vu86sVvsrkc2KP8x/rJoN0Kki25YBgZxtzEuOFIOn+8WL7FzTotRQTqh
7Q7TF1PF+dGBP1v3aU3m2xgmW/vF4pwJumKF3gsO8HmK1Wm8umWP+nHeSbc+Tb19bjoBL0slMYfc
ZMUeb7oPDdiETY/GrU6vsbqApPploSQU/8ci8IEz9e4RXl3fabdfZjx0ls6vsP1uQQObzgLY8Kf/
I11bClj8clXtCP8DJ6AeeCXRnWJOFFwOIsf3Ixnq9JhLNaqy0IkE6qbJdymt8fg0FK2S5jWnmIjt
8PiMQ6jOc0telOcJcIWCJYSV36/bRE9TjzWbYBczf5VXrXMacqU3JvGaR+IYtg3CLAEtsZ1H/UPl
7jy4ZoJBCliD3YuSPR0VCc5/Rdquxtlb3KEl4HCfZWCqt45bjLhg78bZAJ0A0jB35jC5NBXcdBC9
PonWXykUAM664V6PhEO6Drk2wH80b6Dpxt5+0JpTdOEvhYJ6e7ciLtADXkdwuQhMlvdaPXbtRBlN
0gmiGB8uKlgBFw3eBi9VlHkdq56kqsuJ59IOkyczfRorNa30R7vTmXY5Nc9b3o4t25kI2N14j8hd
hIJSc/2SzPS+sieJQMNkgCZDIIN8NTn99FcWm1eM6BZTDW5sgSUt0EgbIOXbMr7R29RCQq7DCzpU
B0B05/hixmEwtDPZqibyFWWR1rjeK+sbPY8EQGJ1I/ZFd+zVI8a9UAZPqvolfaGyqWTf9jnALwzS
URuD6wTpg5oX53oBJCexvWyiU2S9XZv6i2yU7UGat1WfgGqMy2C2/mNJwQITQ7ziFejyNu9AW7oe
L3WOGX/8YLVZYWc33gDfuI100QWbmfeT80T72OlLYMQP3sQTvHDcNbWdfLz4vD/z4nx/9JhS5Iub
DPxLa5I1wAR4Ojj9fpFy/iU0dKCQI6+3Ya1hrkAyACX2nO47w1GKDvBpTH4PcXnP5f51RjGDbGsg
dcyc/SJy4h/lvef+6KMaClejomfa7Wavmg9KkdIzUqQRNJV4pZebe8/BSDGadxMMB0LIy9+RPwOB
yLan6RxnlSKZ0zRZVhPPe8FVbrBTDW4AdJSG3onzZPBOv/asw9K5gKGORqC6nYw894I/OOoJ848f
PO+lXo8f+wI2KZphmvJc7MSVA2+1JIotBdlmaJK+fkzHAFuumIrP+5JCo8sEFbEYNGuJMBNeaxbj
3/UWX0kZhMND39aFvKnXhhE/qgIAdw5bOVERVDuL/+oeYZf70fXAbeGbuHSOwNCQAjjC1O/b/LOG
G6b2QozzdgYng7GujgWJuNou/INwAa/QwFJ3QyggqW3oN1+Cx5CiTs/1N1JQ1QGd+/PGQScmyENG
rEjwR3W4Ywwd5XprVKbXWBjHQ+7AJArJncSN3ZQnPuM5trVncyQqw2KxibQtlED+6bpT/Nz1IyiS
rDk/9LCA0oZ12snnHL+k4jKTESzDPt2ijpB+AqabYIvel32p1dUbK2chUGaVfGGkWsMDXd1ENClS
HW5jO4RkEvPwgKtknlr1Y5jlurBRM+SOXPriIhuIfjif7cfg+8atMliARN7VITiCHhaAhnwd8wY/
OXzz5yd+j3t/C2g5WxJrAAj8X/j8vZm3F5L8NAsKhi/l1O9pcLZTfYMPj0LO0TP/rHGO1DSxuwfc
PC25cSIYIseR44Gnjql3sYho4X8dxPHTnaSRxHvVnpHgQUd9bwTr52Z4HtuA9oxdtfsWxkNVmyyU
TCMrbhKf/2r/z0o2NuGgZgX0wx89EEfat2XR3WqcGioHMY78q332EzPBoxCe68ui+sd714FCtcew
ER0LqYsFslz2sbgpxmPUsApWZtqYsSPD+r+jgQXGyZyNOuNJg2N/VwjOmSi41pzovvc+9rAx4Q6R
I9Uv19+i6BuWwjPVZSxpkKZYdDuDRsGbqKLC/UKmde1d1SPa3Ia0HH28uf33rYPgyDrfbbPOsyGI
GRXlHdJYO7Tp+hDF97GtWjWFj+K+a6tJ26tTgLbTbF9KxSxl5IVF0uhE3MYR5kKrl6sXnhwA9Bph
vF5jXFrOEY1RhjPmJ7HS6WC02B5J0yNVqiy2RlnX/HV4hLAK8T+53VAEsyTPLYNiWdfGfSS+h0gr
M8ByhUSagWvwpzKCvCc74zXUbiWUdaA21VDWEz91loG2mtoZ/JiSpE5czDL3ChEwxoJu5bt35isA
Q+lIrWuRuH3NM+bGGt5oR+7QKgU8SFspCYgRvZo6Kk8g6RN8Iq+RxMHywTDF0bqRj6RHmZQvDSuu
uLViVU9Xr5W83VDDWa0GR+Zc3MOTMt65Y6odTK4LGZ4hIK96xdmpxJFmIozVUpM0DXOCqX38TA8x
RJQeT24c3JyvJPI3kQJixNbVC7jUnXVzG9RcQRpnosqs6KM/2ViXMfcfsy3MPpCodNidmaZ7R765
nofIEHZPPEGChcFiW+PNipEicqOrOAI3xjcY+qrAO/YmxoMlg3bBWaMtn6dWjJ9OJh+WIGTfs9I8
6ebPsBDh2lP4SQlDLBTxudz+4iw3JWdioySjb9U4nWe1gGaeQco4LjCQfw0a/WT2LugFsnQ1gfsV
1bc4Gks6EeRrdQZnhPfJVZF2VLs+52pCwStiYxef5pTnBDKpIpqVS/cSsQn79p8LDRndduyF/d65
LwH7Xf/58xIKAk5DbaJ0+a1RBEhybGyt4TQwG1P0J1Im0j5WOffgr9Q2bTahIcyI992FKwxss/Tb
CdtAzFofPEpVZEgV3nDHGsWf4cZzweJrWaC5hPe4V2BdOdNY+82kd7Md3orGZW3qyA8tPaWh8br5
s0NBqDiVv7h7BYlYsUe94s9W7GqDO/4gEa0uNRC5NVbC+mNXX9kqITfY9vizdJHcQfNr88rj+lV6
Gn9BDTJxhJTkq/zCF4EGd3npmRpm/0Yhc7TB+nB+PBOB7qIJungR2oMaxqiXFRFcsx+HbasNt1IZ
IdOkmxhaQEA7lkaYxJlPPZqKdPnn6VYwCRpSzqcGC+8HQhaPZvYYWbtQLdMKQ+vae1QAcftxYVgj
tz/vSRhqZlfqOVn6Tt7YdbEvaLDwAc6wdzE1XbXULkRntL5gNRleLxCFiTngDlpXvedj9aUJ1Jjo
vjRQNi4+KzpSLtlYlsuTF5nVFVDXjwuKZRw9q7X5KV5Tln3DjDKGcTc439ycG98ya3d74dpzQyaH
iHgJrLpirNQrUeu6yJXeMpz+klYK0GqR1+w2tMOWDd6NveFnE6bKFqQGcOnmKoZcTOkForBP90qF
mHju7oWauxEGizKRh2yhbWrCuyY/12/xIP6Ii0YflaY9XYYaNp8nPhkOR5N2mM0SrtkGX1oG6rHk
LKp4TGQx603PKpuWsr+4h1SiG3jDJTabhjRbKeQWtwtVmwnY5rGaPhmku5kiunXFNMvwnbYNdJCz
ALZg+wCia+lwOBj52C58wuQGIyTbb49Pz+++vwRKdQqrbJSTbmfYtyh0rwBiJUs7Ah4wfFBW+RXX
5psb154lN5vsOFUMe7UKutckC11px1qZ6DXezywKoO9C30m0Qw/nbFrHwT/GKLP6mxcj86k9vLLu
ix2l4p2ZB9C5pqGYYy/LsoCpKfrEch1Ci6mrlCMSNAjsLA09ThOGJmcuWVUtwVw6W2mI0DzO9d/Y
ml7OumA7opiiJxwSf4mTQYNqyT2N2Wv5wJBmO4WSPzXK4p51kJTUjrxL373jsvQD6mIdOZkFs6r4
bN5hzimsXYZ+UKbyzxLeZH5dWTA3CQHwh3QZg1dPOzWGUGOMQXp1fFkcY0BK8Eelrk34oCiFAl7I
CI95LmFnYNvCBs9LgZB3sOaV+ivQywjgKHY2sGxzAHk+PYOTHgQs4weACFo5w5ejJGhhTtQJKNct
f4oRUgGjD6XRoxmK177MbyEi0pdlQQORoMedIkdLNTFPF08lbs/rlqXMaiUMkqM1YQQsy4XDaLgv
qXeDMgJ2nWPQuv063N6vjLJJqOIw78ZOA+b6P6yqAdZd8WGk5LnUGsbvvpaFbHLQTNE7wuT4GDlU
zGKbw+h5/9bPGkfBb8DhAHKKolPmW3AaiIJccW1VPfs4mdKl70x8LHBmxe/pvG6pmaeQRNW60HOT
3NjRA3ZCKa0lwGodMj2albn1JP/TKf8qnJR0MM0h1wNZV1KxchDgWP7IPpjvGS4ACNq5+7dIKi8C
JnFeMJumOCo81VtY/Nez8xscylnH/F2aja0E6Y7obbWowMH25uDTeUbAA5OCaaZnOYHNsRwkvxXP
O4LOhPykD4PyKQckgHKPyVH24Gry4DOx8frbxmemqXm2gIeqsvvMQiYWpMFt8mzvi/8s5AwlML8b
7E4o6hgbKFG0S2TQBsTQ3TgjnGa8OWbNb4EWkfzPcpmQ9swVD6D4IOHPZJHEwrpZrcDQN5GfxE2Y
zIueo6+v5gqk4KzMMEXTl6/1Sg8rScFYccHU79NCKVC0NZ9eoJpgfFP3UO0wPqpLAE0lnbQAIKTK
Aeaz+b22+r0SuCG/OPsIzKucvHBiX3upZKgkct5CSToZssRKlozOgliYuTNwKe6jRH9wq9FbbdJ+
a0oA/wRL4Y+wsJLs0dcivelZh4dDuirwmFUu1j7sO4D9YMyLy0BKctdLsdn8hy2qNv8L1mwK7BWB
nTmWnIe1DgPlGZ0rpNvgnutyvCVHaNhT5uNAQLQGJ0hFp/auzwvhTyd2tNKQbyTKtZiL55rGcB5G
XaAN6U/oa5uBrtP2qwaFd3g9+286+LP1MSzSUfFwB4amBfPQstFtY56PihsIiNWFIHC22txq+hYs
ibMoF1etomffIu7ZjiOG+tqYnjiHY82NPbR9Bt/XACX58AD0ZwbPR+ARBe3KQFGhbMup95j7ohuO
fB7zPELtaoEGrKz+pJdu7wriXveazb4UYBvbPqDyUPwi+xpRsOmJBKSTmk0lSjp1CHhftDU+lFtn
2yt/FAPTDNrBosiJnFWfrNfB1QwTyjXLJSsBenpIqA5y2L1r6ud47+6hRDWK1niaBj9d33AYUI/1
nKGC5ShUxDTwlAbvqNLMJSTxuEYwo/cVXchhj2PE2xvoCdVXij8ZPFmKBVQFSDPfEOpnjnE9zSMd
30fGiyZMazfrYbhyQBNF08CY+tFFztXc0EQF3bDwDRx/igpXvOhPHJBWgQihpkblDSbBXEppOYgn
bh19TqRQ7vgISp25WYDUJ20tXVTzZdsArCQGYka1CjWLAPAg9K7cWPwDEOZqTxvxlqW3FHG5AQg2
h9IL4N/39+I4uNW/EfkmstDCAe8pX8Oc+3OdBwjbWLv9nYpuFplWuqworsMfdNGDW208/iTM46mI
K21Gh2aT+7nHvTYYLvHtsccls2qqHvrC04PjhsNTd0QF/N+HOb0/w5aF09opFrYKYUWjjDo/me6j
WAO6xObySIfRmaVlf6I+e21T2G8FBspmlOgcLglW+tX/OfebocqatoBQ+061tfN7MQspRkwul1Dr
hPk+JJe+eZwpbowVcldSE8CDjS52I/Bhznvv0dJP2MY4ybLVQdXEMBgxxTh3deeVubDHEROTmz4l
IXne7l83guQWRK/Va9UkbfLwSjnm4/31rjjYAU1Sbw2iNYM/vpmkIA1CP7kGGS73mTLT6cNnJ60M
QwkIwTv9of9m1zD2dvwS1oojmC5yLH/cpf6S4FN2IkTrcfZ0o2MSTIdWWT786ET0wKy2UY4l+RQH
M02v0eTJ09U0t9ROfWMrPMUSIFRW327cFz7Xlt3LC87WtvIh+xLDOT5YcKMkKZH2s7d+17TejNdS
rWe7MEWLSnFvH7X9hUIy5h6oq5S/L5DtfEbA2iknc6QIsoTZPyMSlMHBdWhuWZUF/wrJC4i/U7xb
LKWYwPLIusJ3AJ7fLpl+Y6KjIaUxgCym0BDE+x9gin4c+KU74v+MhQtgKggdG9RFemrsG1mN0DMt
QLa7/x9VhLC+baXiKRS/8odJkjtIwMDAYFReI/7hQcmx51tWay98Rj9ZVHJ8hd4/qWW+LWQhuUFt
Nf5sQV8uW40qC6Pulud7EIei+q9g01yBT2ih/tHFTmvuJegrpQecyJb+wkRKrNiBAf8u4lUCHYE1
a0A6LW7aKGlTyQ5lpx38gmA/D3Vu7LwNuPyo4qLokfFwQMpx8DBL9tSwhOBABHGx67bcw4zm5tm+
bGGM8Yg2T96LO7vsJ+O0tEhk81PKsQf8xcAbZrDgqQJqZGbf6HEfwod5dJ4OfJUQe5Cv9qTLYs32
+Qg3WTHU+AKdJpyTN3P3T6/sCZgQbD/7OH8COEPm/mc7I36bbHNOhhgGJYr4Z4vYucdpX2bwh8zY
kiaKnndY7MuW3cUIQntgk7Y2ZRZ18IIV1+7xIdenIzeuu3Ng5awI+ViFCrhyFbwkqkCNudtNZ6MK
oCs9I5972pI7kWBvhnheWCNdS/FrZ/n+90pF0l4JuDPSTxUDlsPEteCr82PJwdAKpoCna9CE3xAs
JSWGqt7EbW1Yb5JztkEZ1jasYLfBtctlCG3Kxa/OUCnWMd0kidr5lAayWzCtPSh6KH+ZA517COhc
gJfGzNOKqK4Kg9TAsgMDiKbN/pJnGW+XcuoqjWxjIWHjOm3INItQGWU8ePLaUK5IoAKwEZ041M1K
2IWtwkVbvl/4dZpSBPKnc9Zr24NWjJNh+eB0AcTeyeV+Cb9GxkuL86ZLhd3w+eh+gkNvIdQkiDpD
iGUxnIe3Ry/eZLFg4/BZBz9obuvSiktfOjTRpQU6LgZnlSWaSTLQeqqcMDvoT/vbddIX8fbC6hOX
si6H8Jj3h2banEDVhFPvBinqagqJvgjjqGVv7xSL2kJjQLbpydVlVBpZHqms5fQ93v2EzamRPVqt
xkAioJ7NazaKjDFgSsiArnTNVJqmifiR9z0JhogACQa+/kTXB61yg6NEE9C5UsHeLx1LLQTW5et4
qVCgq6WuW0wSXV9EAjJ2inUrp0Dg1mcEMcPX7a2FT7ZHYi7ifzZ5u1f06I1sjioSBadr/9BvSFXq
OSlvHs6nGNLdYCVfhm7LY2eyN4LYjRRF16UM37kBghWf1AWyfRtDDfZcCBcYuo9j+LcEJKRx7+0g
QaWsn0avRoIib2qxMUkVOFWhkhLXPAlY6j84f91oDVnpNnO5DfY2zbh1natI+radAU+Uw00xxX3P
d/KoxKLv36/P8h1Nup2eBOkDDnQzBk7CexEsu9Ed8RyUHbFH8tBmYSHY9jIAqlqbQymrYxajbLkg
IrcY3W/3rm62oigNbWhHMIRrP0brciVVcQyD6tkkWAAkUxu+9b9LMmOLFCf2ILc69SRA8lk+XOq4
yZuaQMOkTDvyBoAfy1PkMjgS7cGcQH8e9Qud/+v95OvbZbKv1YwTozmcGTcpepFjiPq6+HHGJ5qP
a3GH6P7wPliLZktVH933jo2JmXHHKHeogKSV+04Ij6HUshE+hyqqbVTPJ5F2weTLvfvbYYdp1tA4
ITgpoxOtFi3EuYH3OeSjdGrA87DqrHXWJdAVBpVHo3hl2i0Tn52ERpxaxW4usvtb7S3kJday02XB
QxWoeKd3w/ipjCrWHGBcYsEJypChu/iK7yEMyuneEmojWNuDXdlMcESZ2qFewwibP8NOyTwXyeWm
T4Fc6tM13HNmvP9kNXvH6OZoZHFbPoVOd8YMfPHyZpPndnRMHeprCGsSUFK1AXSJInWmKZZpCnhg
Y00LEKwt+3UdYWjE07Hgy6exGQ4l4r+z8CN0BM44pr3LGIxX+GJbwXyCr3UWYO2Jj0FaiIvwLeDX
ovirTfXzEDpQbAkIUBk5clnlj+Ry86sJ2XyjbmxXN3m7m2FN/UIFYEndnmdHU1fRf9cAKjICeIUG
r3gLP3VcPAcgchoAB4HPEoNiU/9ymJqJgrfpkYAO3nFuwxAIMZhZ0A9du3DdK/H3QcgV2Frvi6P1
7eei71AYfJqAYZ7U6TEyyBgUJUUSYpA74oan4JT+bVYE+seYhoCZFHtY7auKZHsFQQhsX3/vJWxL
2Ie61Rd+q7zkk3QR4Bm40T8E3fdAx+kARyHuhzUyNt7NcepRu/MJWQieoiRwezayWffTgOy2xKpS
YJrmQViD42Rl5epzr5poattp5R5IqwZtJYcLFenBsw9HZq6i0aN4Zuel7Ax1X6E8FDSTPBeryCR3
VowW9BzdrdlkUorh9BtqJsz7BihZPrEUjZTb9dL6BYVFNavB+1a+YewtCL5ScHoVujvTX6JuDncR
LygMCNg01I/lCf/gfAJIAeDfWaCwpQBA+vi7Ki/NOP8jFiGTR79DfzaGNrLKlt2NgVStocu/I7Y1
Z+jwdtwZ7TFwZY51AZaAlz1HtXwQlF5v4GcZF/gOFAbegLzgBTnrvhkZZIQD6U332/yc9tCQfJHx
SEo9aUdbCP1uXDmh9AtWAG1nrYrAEXbU1ljGlGiKrdS2O2X8HGGihmrwrxMz+RDSdoWG7HsA1N7f
iDTC/q00V2t24M7HBZUjEC7HXLD7q95TImyGGTy8E0iN5iZpc+3zes8JeBvgmgvxf577LfuCeb71
xk1fq1EnJ8UMWWojp1+wyv2GmeRbppDC6oJLBHcCs508wPON2bm4W3icvOPIuuhIc/1IqvQ3M+oo
TRrZIiuAQyWqqgCm3uDruONnkZLpA1KI4/60brM1GWhdxsOSBnEndL4vxbdXnBP0nA4mkLd8vC9V
5VH8tif7d5aoGr3pe0JDPxNTyUsAJ9TiiNzOFC/5btKzzBmYlylqBQrg1/UYRxzjmqQJigZEK7qL
KLUOxzurD0UsQr9IGFYJjN3mjm15loFinmlpAxvsG3Rdu0VxbjZDcSx8sdxhYNBuODCOZPVENZQ1
5kXzK7Jlvqks8AKnz/CkgELtX/fWQcbLh99Jxrcpf3C6k56x/6OyEylz8nB/RjHZCDPPGY2yGWrG
zmJ4B9T0d8ZybaSoVuw5bX+ZHTa8tvdvhb96spGjpJMc/YGxh79CvkgfRCZrGRv3JI3nX5KpYO9F
ok5nDT9JBLaXEFLcJ9ax1cWAG2q44jI0NYON2AJ9epPtrBPtF3kDvIn3JPc9fTrHvo3U8cWsHOR+
Dov6qsjazdEFvwcqG99PtJ9VyoxK3uN0g8+rmyCqy3avIqHAl1ZmfCvC9sWtzLgz1ClCX5GeNhYH
bmKTzkIjpumZa26sq2lspSGFwTFV5qooUk14R29iNMzpUn99KbmmlP1dewaHVWCIGHUaXZw1u61h
eIW9kYpD3EdHLfNb3LcIHrexOrazDM/uo4ILMkWD1l+/4yQ2O2MtUgriOiiAaIwaVftDtUXdzCec
G0U4RBrcLhE13nhDJZtyIkJg94FSYtfGblrJcCiN/rD0qj2Ft1AyV24EC45Wj8/gbXsze/umN3ST
ptUTWMkJHIdHGA4JxHQEKw8F50zGAzS6DkE7f4v21OIs97/2l9hQFqQ7yYbWED/ohtWhqtzcCPem
9aEtd2Goh6AJy0003yOaHSiHkTIIx23o7jNFop3y/+1f1aXv3vfNKvQ1PZavUSCGRd5udpOgYj/w
iNcH/obQj0FKpudgdo+zk+D5h6wssUqqfx78jaQhCziPkwVp7UksiOMpJGkGuscbUkzAfV51SFx3
jsD7q3Sek8sIvhm6Qey3yC/nLYRZ7iSgmUdopSosqFHTmGmkF0oVzqanQXX5rjwvRxisJEaDDMo+
5RMWGB/hRr3QHTTXHC0w+AiddCZ+NK0eaPRjdkkndM5pJC/5lR9x9druYPmnq1M0uQIYMVuMrwy/
f+xB+1NsN9UpshnTv9wpf2UwvMt2D2vZdlLfviMUjC1D00plVjQ4mjjvLqv5ydCBSnt3zyEKWA7c
ukOv6MqCPsQSNgpDy6Dm/uD2BUj165km2bLKb87G5TVlUkv0yWUwL656x7RKKl1mt1Mq35uZDc8g
zdBd4ZGTmBYWxwune80Bp4VhkoZIAGvdRiv5c6kde/s85C07Dm+dbVSPvsg6I59EkcMPAwMyJAf9
wZfqD5W42f9AUK4i5nSz9ZOxsBflM42x8wFx12NMJ4APvGMvcDOilEJ75pxs/NAqDQsFh1OHIBH2
s2wTmouSjMcWRm2I0BekKcOoZK5hWnYfWWFiqVDXqCfzky9xPdxdcqIqGx0Z9XXC2z5/xSZ6w2D9
zVe0NIy2t/K3S0Gb2bZnSkyAeKqMZ1K/RpiJh/LsMmzNCFWNMnRLdbpeDF6pjvpY6uHwBjrkgVvR
ozKyL54KjRPy7/W06bGNb/nIIvolFBqxIeOn/svTS8ED/niOTDsS0eiWHQeCH5bDO4nBzb70gZi/
rUpZ7NmDF7OopUCDQPcHgSC4qciKxD8VThuOczyPO6R6DipAV9kGJhNnYztLHym1DH9+tbKupeLg
ukzbGDS8UqT7cFL0kgekr44ePQ5fX/DRYTP5JePCFnfBwoNC8Wpeuh6fwTdVdU4NOkreffb+zg6i
opag3c+BvSYY4+G529UWRgdaUSAIL6z4wc2kYtoKOFFqRB4ZHUxsacBPDj7D2uB+XvtKexrZqNcl
tDUmNqlRsK1fIQ6ClcrPQQs8EqhltZp17Sv8D5KrPH1oK9B1WCHSA6uPU+s5TwtSWkKLNrJS2gyj
tgJKGirGLOPmj5r9SwZOQBqi9c3wYGdS8I1KIAj0MPr2GLWOxxsZRUh5vUDQhRr+AWp8m+wPPCDg
dhWumitF5KEeVUFWoJSjopGhFn/rktydXx6bkXGCaqysFFuqK0GeaWzinAog3D4QrKHy8isHQ/K2
qnMDI2uNLyPLBLEqXq6SmhjFNPP0yW1EpwxlQ4OfdMCbz7V+WinKqjS19SgYeqUdWnhR5O1aykwn
nUwyuGXmh7Sbtkl9BRfIHKOjdFYsS+P1LRE1CPDXhcSbBgEwPh52BHfAwWh0TFh4uA5nBxK0fqBX
oRWKkkTt9D24etNT12GBVUQPQ/9Ntis57qo5J+HDUvHh5Zy8ygwPJ3e7dQz9Jo8/NUjUCdqj/Sz8
nZmsdaqH4kJf2rbkNGpm0SVJ3BBUrWcxVgctbCoruqCDCSr27OKGZVIV+fkSAhoE25JS3o4MX4PT
PBQEcyPf8nOIwIJi+TV8qSBBEulIaTqZgJcN8u28zvWGtMJ49ErU4uXMp2tSgtt1o3j2DjNj10Pj
rZk0aLBUigX4HPWhF13MODAb1e3Gf9FZiKPq3/ZR0qPSyNwih6MJinoo8+ULb+pj21wMLe63vYKc
Pz+fx3ZzPutcD1H+Y3h9Dv7FI/ACigEW20Ov9htjqO3fu1BSoFryAjrIT96dhal7TvBIu5UrXAaU
Ru3zK2LS9+om9pcThitLjKWbd1EghXt9ft+oloT4H+nSc8R30c0WvjDWhtahnHdV8EaYBBfTksIN
o6wRsFrf0eF3NpgKWd3WvTHjoDYuiMTQK+4XxCcS4DyAKIktXbOKmCWts/wTKQbriIsE5+EWsFap
C5dVv2OS2dFshQ1tz+HlsqxtftjZ6tpnSwXW8cPw81oJTrBJYpo0hrb/H4Pfw9NtH4mqtKS5a7yt
6xTubZMs9Jh54Gyx6viuWRMHEkVH8R1kZ0IQHRCgDURUuT03s+o/imai7MjauZynxxu2MpRn4tp7
YGdaT/kjYIqHWo9+E5V2YOhSz9CCOqO/CEkZu+eJ3SAdTZYlGbVshnGy2lLNS19xjdtF5goPZard
R1lyTQXohAsbtdVj25mNuTsmd2HB4AZUtk53ZjRbD839LgPSoEESow29TztPIJ+tZBtAS7dNKfXZ
7F7+oF0grxkrHIjSrFM7rLhtqTEUQAgaBWHcbvu1vv2kXy/6XE0sDN8UF5mXbH/EG3TtllV2VN3S
r3al2CzYKcTfv+wCiIr1N2vo5pErY9wn0mfcwSNHXO48poo1k4ok23vTCp8nM0YYryHS83bh08Vz
saCaM98fSjG4PH1PRrdP62chvK8GGL8Ihptl0R4qsrJDMrlYhWPoQhmrlEp1RxaITaaO9DnRSsd/
qcieJa9dsT/AtdH9sk7UFqRkY3wNYf63Uu261vjzfc59s4DV7UFI+HqH5ZXqd0LhXMOJsFWS4eRD
sCd/azyvXjNOKUj9yKR3g2CovGhD0ym/5npnptXPA48c5N4Hsx+ThIJ3oE96AkeAlp93TibPTP40
w/kE55EYQ8fM85GMZ5XI87EDjj5jfELD058TbKb3SKX0W1gJwU/I5582lUw5ub1pwqmfNte9hILr
D8MwfB+3UvpOGcPYc/6iNEv2lifPAh5iwJT/9xF7ojaOIFtrhxQVusUhhXq3eclrXJK279+o9JaC
wzVIMCYixAI8LPG/ZEILOQzTYn6poyl2KYmQoIXjqN1MSmUrNqMNX5GpT2KznArv9Oh7QFxeslAV
7I5tKR6QHynvl09AAzSlgutPMmSJXkqdweK10PA5X3UDfk8JWcxhIUXLQyXce4hLYXf5yV5+wPzs
QEX8dJF4cJUlzvvuL9kh8EycGh+W6sTiXJCo0HmtZiNq8tJb8aBup1OMG2LBIvmaRD/R99sAjujt
u8AIHQb3Cv6OmNE8oq7N6YS/Yj/cconx9+ZMgu3GTtRZ8yDu6cuSxXScha/WUcubP/OBhC6+c0dn
VEDWI+PedYg9LEbQwziELAJ2sQFGzb1WWKD3f5iJmHD1ZksI3QeNKJ3W3YBkJXGMnga+wix9poGa
MuhDOID78IU4CNeeYW+HDxnHJLMegkP4O7M0I8LcOhk7aa2nUlUBuhLZFqb+DXH+VqAfIkYStjIe
lplSqylH9LMkGR4bHnQVjZgxRwlmWkuK+3WzFnss0LAqOP1JwbXebZbaUV0LV/XC/nHJUNwLDVGo
EUGPgfafCFqt5niFupJvF4G8AoDiccuymVCadChJSDSm3RA21p1cmi1gajePMwWQ6cVnhl15p0QI
LvoelwGVstRr/PLGWRRKQOBTm6/lJwFy7VMK6OLtjYkTr4DwUWVHDjv66baKTnoIQMhu7H4LUQR0
TOL4WpVu3FarlGtqNOP5uo0VtWo2rGTcEWJhGpWpq9LFJbySjO7pTIK91fA/62aTmvwkjWrvHtj4
trj2AeN0bb+as3DBX2SQvub89bcwTBwrV9cSasHaA44O3U5J205LS+b61hK/wfX/qMbvAQqql6ZH
5RDHX+bPGK9VdIvQSh9Dp3UtRb/k+iolP0cl7wWb78XCXknMYrLUIJAkRYNQRPUd4Q54bSwfVPaG
4vWjxM3m5mpcNF0rKWJKuoCwB+tvG3jhKfOvGvnqfXanj94l+W7W8gkkLzJ1DrvvCMhZa2KmBXvI
bKfCzyLyam100N0c7qweArBREBq3n/gpj+sk48CrGi3kgrg/cNu1LBGus2FwZGZ+e9fNpYTf+Vi0
YUatRRFcX7+IVkt/9M+dvTvjpvwc764LSwQeLJx5VmmIJiAa0taVZYRDHEB7lTpeaayzCLOCbmz3
6NzqJoNLhgv37YJV4RSfV+p3h5nTkLKUVHK5Co5CrMFcHtvK87v54zmzpM+Tue+jqdyK9t7M1csu
5y3oBMs7c/57ZIWNc8KSM+Q0lm/HcPg0xf86ixY43Jr5Ntf14hTz37VSGwdeJqbtugXrlIXNMA5m
byNNHdNxnOLlIjSReMj1xdHw1Pxog8tp4CnrQLUykWy8kLSSosEBT6okORbCbnm3YALTbTq7kdKv
eAGC8Xfvj9ZwsnFAZWh2TKN2/UH9n84PWKmv85lIDdCPhonzFLXCA+5y+Td5EXbpDqagRugcf6CV
DpfxkRmw15WKN5vB9a1f7lfxwPjSsKyBNgH8mrjlhmxG+ZErawrQuMj2YT/LYcJ7IhwbhA8xjT7S
cZ+KI/D1d6LP2AMk30HJuIOJ7cUaXVHSXf+bU8OB3Q4sMAffvb4O4KGR//m/57DA6HXHb+lSj7VU
tC4GkdZlFnkLmhIC0drMA5ViFLiVXURXyWtEMuqqKsFWYsXHf3OqdxFv8qR6Z7gey61ibvQ1rHzi
slt/lOqWzUjc1g2+OdYJzHHhtPLOzQB39wt4TUNZHZFeFtcRnRt49NdAoYYt9v3NzQdASRhYUPrI
4b6+n1BNkv76mPOUkeVi2B+LIZmagEU84bJa68FrdxkshRmv8ntqtA4CDl180g2r4Kwbodh+3pIK
yDqQEKPkEGxWFC5CEeiWPYqwnjudWQ/Bj7HG2avkChAI/4CH4euZYWyqQDDZWngrRdgNhG6VEFtN
S9HS3Le3VXIZGHC8MYq/uNRoriUqQENHRa1vib1LfSaIAnuSxNmyNOeoHVgDnWKOMAJBwc78l0n8
sZqzRvG/JIahoXHHlZml3LV+MnHcadaFBVI55s01tOZ/q52sqBgiPP6GstfeI8X1e2ZHxcL+tm37
DuUGVRjbfKuWBAhVlu7VJ2Mh3jklic0X657CjS72PHqLiq3ADvMRzXIEXhlEIVr9DNePYhJnuf6E
1ykm5F6HBBqZ8VgG+IcHPG30nnoZsFxaKGAQcqJD2+bGR9Ysoaobb+P8InGDKV/iruX6uXmIlrcB
Ape+Uz+8wvN/i/ckwlCvzWkvR7SotVR7Om41hTveMXVDiDHbjdjc3OESbZKtFEzzyG26vTQHEC/W
JOTVOYvtWTYs7VWFbMEagA8glUFVSkCYPr3PQUv4GKrOajrCHqHVa4LOEYmzWoqoNoHHch1KtoHE
/0mZq4Q9Rtjxgwury8B1V7ioe+JX/PJxrkM2CJlXxx+vlVZF4Izd13JYylM96zaSymJipP80PnmQ
ixK/Z1RPsTZIRnFHZiFfcdHjxHOhShcSnJMcfrAmFyk2hz2LmQPj7IAZVH7ohHjGXWiPasK2GIbE
6l+f2izDLNi1ZgngP9eOZGbphkBBOgi9xu8Z6oryU0mrWFma4P3F+RLFTA4/xF3A06envAixgsUY
Fg6psAbqeZeUrHzW2QSuFpawO8T1+r+h9lZeIBQQ3Ed/4DuyQrYB4BxuHJaj4vNQ5p+Kuawykx1P
f/ECeO/LnYEaaXXXyVrUpyXuG71CjzLEl4pHKw16DOn1JkgQv9PGrYG8nNgiDHF/8DDROB1hPjc8
arpgyQso4ru/wbc3501Rs3vPz2ySpc4NWgVzBjRv4Cs9cpqgtfqY9gX5N/T0OURLBZfnuHCx7yH2
TuoXmr98A2VNa+mXx1HTY6cRel+8BlNzTb60O06nPnqT0flDuj5292Rf3r4BpXpY9RbdtSLD6xaG
MmVLmuDjQQjSsBdXm/AmAWWa1QRtWMXgJeQguANl6EFcpJ4760GCttPn4cY6YYtRgXGrhiC0t/QH
AuLNX/3lnlwutwA7p9UXbTY6QY2LttO5VpMgTFSdySDhx/GDgDSTD+bb4k+J0dKtboGHBMvrwxkj
2kioRUAyD7hMPhysiHm/ALIh0HxUq2Drp3uNMOPeXKH9R2lmZTvOFabmGXQA1MLftRQE8qi4NAwK
7iEDMw6th2I/QHniO9fRb8rpvbvWutDopWEUcO5yTnuxPuiswVOJ+Zt8PllMlm41UzBv+ww0pXw7
r8SB7fEvlCE9i1FTSrTruHgJrmAbywkdHLR6ptdKd+WISESl5CiS6i9i/x3VbFUkRkhvTZFUd36X
wuAg+hem+O+wEDmxwl/CZxnO63Nd/gQURvtfPCPZqTwYw2YE9JOMoFxhwMq61HMUH6NsNdcGJpXq
BTuABpq91Kzw6vNMbQkzvevWooJHLUQY3ecTarNGSgtohEXtCoPF8HvhuuWZz0kcLcpvSj+y02AK
EuJA8kQLDuNB6Fo2/t9Rg+JP4FuNw9hFXmAwfm6vELfTf5oBvkLLgLH0CR8PF18bQLarB00w/RWN
+thKTZMGPC30UkTztvnUuzdrdjCZDwLUv6lZgYIxVagCopeQb3nSbh99dUzSrlxtWm6rkHnkKWHG
WdxxPss+NURCD/SkqQW81FAPNvXZYoUPSPwwPB5UsW5drklemJRXuZb31KpessTuf90i8qdazQEC
GYalu3vT9+/vIUNOmdXguZ8R2Wi8XZaASBFq8ILa1MefV4fzH6xB11mV1aF+UyO3ZnLNBaFBRwTG
oxFhi7L3v00E0FpZo6it5bmPzV19Exhy/0p0QEra8QhgxC+Ses93d7O6hIkX51r/E4D8HXKBI5/B
ILqmuf9ruzMvsuVXpLA7cR4r1loKXAJktO6xXaIQrXmZvP9rAUZmQBR4/wBbGy7eyBdAmm1sXRZm
f4SDos2TMfHcNEFLIghrkPOphzI0hDhtyF3p2gjM3z/x8onXVYICGhUYWj+pmLtYgYAf+mkjdw6Q
ktTB0bPmo10VNPnTreX0ZFwWmN5/fCHKaRfSsAnX8sawSzkPJ9InC+D/T4EgGjZ5GeQPwj5u+Eux
pp1Up41BMUOSjJEGkiA3F79B8cUt6TJ5ueGhXytHskkuMNNNfsuJvL0GAwBe8Lin9Ja06RoSK9Ux
AA4zGTnUvYHoBAzKiIaRV4ysnXBbDFrloE6EgiHTmkI22/zLKZlTAKuyyx7SN6YUOT5AkgGLrjG3
anYLzLBnq5+XnVSqqpDvOTa3ZBKk+g2fLCuPAg68Z3qHD7IagJSs5z6VQFLp0qGwGTdZumiOKAqy
YFk3p0ZSpY0vbxMJXgCIN7wahKqSi8hmcFamsc1KxTc26CDvJo0PXWg5vYjAosrsMuY4bP0epWR1
ALrBJC5E85tUyqRxG7+eFehTSJIww/CDDA1lQAbSTbNki1OP0DuZratL8ivfqzcc2wS8+BH3HdsW
Tsfqnzy4byYs4qz4unpPqn6BaPUKQGdhmK7jGzdiTAwDc664yaGtqBoosXCG4KVKYeINNDe2JZt9
m3wzq8gFwuFVdBcHXrw3B7F0ZbnB1oy3Yc8NvknFttgFGV7X88XvecwF+KCHUxIL0mS2EM0xcwHE
9mE5mgSgcGhZwj0+amRsv9AU1IE6g1qSRUjQGplqjSMREQmrMAiAuljdn9JaMFi87OxCF9QimSX7
2HDYGAtLRqlNv0GeIUCrDeFspdGo0Rr1910X+PfRdlv7vGTojijxBk1Q0EYFMXZBOSP04UAqNySR
2B69PcnV29GtuZP03v9c31uSuGxDaFQ4gtkj4mU9Bg/TdOa7QXXsPJC/4bfJC9VV/XMsb2K/c9iD
WTrBRhK11KjzEjO9d991reqMeu1+1xSwXxphnqMu96QrPOzy7JHCdtlUTw+dXmu78sgKGcRqEc6I
nqZNraY1cVtn+DH+9LEYXaq6cmCUxlNK0TcDL1q3hOI/MTJ+kAqW/AVHMk7m+eygZLs2jr+rxO6W
X7dig/6MrRyqnME/gGve4Fo4ue8Pd0g0xsRnlh6exo6UHyhGBR66haeMj6n7EryGZvSA4GbqU2s8
gPiSrKL0oZP61N2RjtMdxip53eK+teBQ+EwHqXh4R5gtiOHad6BoqmjeYc/TbXVA4RjggAC+TrXt
F2uZYH95fEGiER2BC6DR/ZoJnhdokOsut3EdFo0vVvz5DiQQMNwroQxZW54tlCjh9Z7EPb/Bvktd
OPbX1cK1mS5bQCb/ywBfBkCVU5WOxzAT/SyJa+5v1ZHiELD4If5y0aZmb3gt+AGwoi+Ei8RtneTL
snxrUEL7o2OFnKras2OrTc9Uw5NKpCPiy6ineD5PGUlyPKP6rgnA51780ntASseDuHrI+kmbxVZe
xbt5c/WhjSR9r9VjUJym2jEg+hdS9k6rUFyMXYVCz2U1qn8BXE2w9C/uITjIutXjiX/aTc9ytaGF
xfjgfq27vcLUPfXKMLtGV9yA8KpDg9RUWHDfZOog7qf6qEbKCNJ0B09Fv/XIpquVt2gbdhp1wO+o
T+wyXHtALpbBS2dKNixzwZY4c4qqLHDuvZ6f1LaVw+rRzMapWDZUS+U2VgvByCoVp9A9NJOgupNe
d1wgBfx5MslyTW8Kqhy16C4Jta5MUpgsqu6fZY6Ui1TKCu6uJu6NGBsQzEVSXGh277GivqyoXkTY
7zpjnoZTBpf0tlcEYHpJ7PIf4IVhoc8SHp7ZT0cwPDphrrUsSsXFdlBpO3H3uUorlfKnlqfXB3YV
ybxkiTaJvcCrPvjv2rfa+Lc/twwvegjudqSD4xZl9tsp/AC8rF3nSecXvrLJO7jYI+YvD6ha4tlD
18IKSH5rK2E9vFZ1EeImq39pUmiujkbwjUahV4I9JFDq9UGWRXPtLwVFkuaa3ySo4Rv/y9CclM8b
L0fJoXKnBr/2pSs9ZXUOaMUGLSmM5YOsfvHll3KH1fgiwU8Htc4oQkwp1tRZawazNIgN3PFysjPd
UXdzzxXghlOdSE3TCNucUOQnbOR5LAR5OeeWp0a+KxafvUrtyVibAWuwa0FXiMtMrICwaX8lCS7O
dHrErl609b77uyipycsC7z+StLp43HmTFZMfBZsH0SPXruL98R2iH6rWh2fHF1UYBcClclwK2S8A
mSQgXWqPY/7b0xxGlAT74DIlHNCMxg6yEoY65+UUbI9CNGLhJg/pNERieK4Iemfi7ZuZbqr20vCM
3C9i32kxAdEFj16I6yAZu0nRhm2KseSGcO1oCBSeTITYp1RPQqnEOChMMBjzbyz/6fyPiV6VW9Dm
Z1I4KJC8mRygBGUEEeS+w7PvmIPiUVm1K/6/m4LyYUhDXyH7c0w2LQVlTqM5J3QEmYuGGsASEZd3
7zfreFN0+OVSVlLKrOvTwvGB/D7NMn9gkvtsM3VSQP7iI9xRxe6qrkVbfMkSJNHJ9fDfqyMg9hZ8
1kxtiN5ywlbeVhsv39X1ib9ddaGpEjGxks8Vf+Jv4ghajVRZglweCv16vw7QbvGppniUfxQdtRlp
HwZsrNlaKkaG4f0cDa/NRd4KgaQxcqzI5SEVbREoO8aB/t8hEWpMuY6KVogGR4r3tYtOCrFQvuVm
1Q4guJay/zzejhaQIXlx/lZBu92CjW6mej1G6kljO15IMFnAPm5qPl0cbl9fpHc2NihERINA1Cyu
dVSUHpMuFjO3781uTWfbBZ6rHA/05Dk29kkr2io46GQgP1nncIBHc9OJ5jhbsnTzzlzHYcf8mla4
rp/+BYUpmEDZosLQ2WYwEjbjLJ65MP0ajEIxSg5og7osPUaOUnFz9dNgUOqwJxagZO5gMX0upW/t
FKl5lohTJVWkJD1NWJkzkloBUo07Xo3ZGYvY0YWzJFwjZd+5kgR5q2GF/MgEgaaLVYsjDOnCDEQd
E5DVfOZKmwcl7wcrAAv9zZPPR0iKzduVnlK1B6juTK1NhTRrfaWqFYNx83cRtck/gXeXpj1vDujn
BVLj/j/Uk9uBWtpPoH/DJAnT0yvd1ufzx095A+jfLH9FgkQp3S5+EFDmbweJicKsBLiNsYKWtRoB
YwihIQS8uURBD7TlHRYR75odkgXCpbguQUt/+EzRB5moefJ31po1dXdR159wMLZ1lFNgBHHj6BJa
k+/SN+ww2zMAn12XrnXhLmsef7CaSbJ0zAE+BCWIIrjWt7BXq4Wh2I0DWJuTMmG+v/tk3ZtYf/yn
lpp//yiZjjlbnI/BoXbeFEBqUHRqlTjPP99Pe4eISUSkB9ZRm4aj3liXLkl6oOdwj5mO4MwtG+O8
z+fc2M7YtREAn2J6GTSrLdCRGobTpg7In3VrvIwCENjMM+kw4KRJkEo2ZsvJmXlp1jcf3094ZAvH
Or27rg90WKXJdg1ldZ2RNpBhUlG+X96e7BxTEuw+TnLqoTFBU0Um34WvP/w99WPCe+ItOowQcE3/
1Wu0dg1GbtY+QaAj24k8F+Z7edbPjHaQ0/ezYlpGZt4FL6qvJvRBQGw/srjTnj5AtjiLFtqUYSJm
QjV8zv67RFt25sNHBNsFn1IAA2hUn5IN5IG5smcCoQyx/uwr297AUEYIE8nCvTL5DvJrW9lagfRp
Q+QHYb2S15/idl4WkOQJFT5jENQlM7gFrJXgwrIyLZPbEFfBJ8JHNEWOna8SV2hw5g5UOJ/P5/jL
GFVxFm/0RwFeEMrBO8Gw5DXDEgqm7K7o7+z/ymvhy8HXlai7UG05qt97QLTQcO2ktirYK/ROhNbX
3AFsdJ9DSJUskIK958mJ5WLZ0LiKdDDZwYwQ8o/ljWIet4CwzmPWi7KajVfPdtRkV3pntCB81Ta6
1FLeLhwWqdx66KExxHfwJ6fl6kqAtiEStLhzbeuMBD2dt+j7CjAqCmrJ+bj50f5YI2RQCTS7z643
Th57PY/KvkFcw4tOH7k8muOfqdK3HywPEswHRR966ya3lFA5S/XszUqVoDNDiV5dfTjGjJSt6AHy
w5w87GCYykNVnoeURgN/A9DbWHCsIe7itViUiF57MRqvogpTaU9Sx/DxKFyXxCb+NQEa/xTpBeNk
0/0LiB75x1R09uiYhwk7V356X4YbemPv6qHF9KDIBbOG+ZRDR2NvfdwZ5vL9xuWYQGY/CUEiHlnP
a2mas4j6U9ryvX69JwSK98EWuvBVWjzOR7ymNgglWJXmmhLw+BA+KFWmvFMhmpetuAqqQcZJyy1S
TyUDw4vWoUEqX/vHfzujF3QtDpAssZUR+fMMocjk1tiQMwrvNuWWrQC/pv6jQ7w0XChXL6cBP/4l
4LubBbkdPbZIFjo47vrjDprciyaOdVx+eGKdvGAuuHhWTX1jQyxPe2fZDWst6btzEYHk+ABIK8Vg
dMcxQkg+kb5axYB15sub0JTtpdjg2f1woAPatYrdwbkKFQob2MipzabgjcPAUr229HLmlCS6mvcN
cMBMzykvYQCe3YWMIL6ZQIzfC6BK1rOuciB0Qx7+uJsZgeG+6qy8D8qW0ZbHCZDiigBFaLvMQynl
psvHqq0yOk7FE6dq9+iUckIdASa4TxAal9yRO7lSZinwk8KjziaxLkPiX+EyOOFuabHdBUHvdmTn
kJAMxGNiEI2h/Yi6zqlZbY3WIbfZ3pXintWmYWA451r/kmr9vmSt2IyQKsPXwHfcHql8XMrr44zb
Acb8is43fmgz7xyYdxA2DlfVNWcNCvFF5CXcG/z0iPqCwyEEmKfN8JOF07e9OPVgUtmPXMlyDlVJ
OPDEqKgv/1cYZT2vDcIQro6ibWAHBsioF+PHBKBfk5AFQzOYzIriHg794mn5+NrZRyHsamNp1tqE
bCQnRJGdAr2z/mgQ0H5hB1e+7D0NzqbvqMsglhDnO96gbTUyLgtVdAilAgnLxP0NAf23/I+pdDFy
7nIkZc/7YoLtIR6clzeqvh0IAEq+o9Po/shfdW2ged+5V7oH9CxG+gdc3HUTELypTmtAG+mir97I
Y4zs1EfjNusr0JEcp8AEMbVtC06mqsH2I4X/+c7wyTUZEo5PDofM7U6rt4/086cNMbo3KxwIHR5X
fnZkJXiQxmh4df1Ar9mHQpOOvRsIWcjYlU3vNle+H5tiHxDMwptEHDPPFjHgVDLs6xeqy58Lf5yi
JJpZCREfV1kkOa24OeiagYY3vq6C2NeY5O80ZnMquCCH7fUk24/Hwa4fAiqQrp9yQQQuSZ6uPgI4
5ekHYQ88wAKEFjVkoNDHklvr4ziYn7jvR04iDtxy0qffrKEaZWicI2UPdWEWsdwwZKt26iFKMd5L
lTdwbEokpQz27RgFC1EYjLWsdZ0ay9MAcMPLw79EWtshE+v0Myv5GerNCNajgzgStRewXfq0nLqo
CSc3FuCndrkKXuWODRrZkGykkHfi6AwHzNdxaj/zAswPKqQGgSXBztFnzBp9Iu0ixEMi/L+U5Uwe
ihHV+m4UnC3Wo0BIaVjIE5wp/uGesRdLA2We+gNjyt7rBP0a8gLicG7qU0Qh28+VBPCkEUIKVTbg
JshnDnkBX3XUQQyJtVxXCCOHv7SrguntZUbh3HgzbOCKHGVve2c+KavuBvXAXsGhR9Xbq7VgrLxC
DO8iOKblmGO3j1+Yhq0sweNBmx/ZD3jWWWDmPq2nHkwwVq0hl1I8UAr2F+M41bY17TmwTetLqpzk
NqWaN5fhq0nJAlP68G8XdHxIEhmsTxQGj2kQkwttsOrbg346CCr4kRe0HJ0r79bep4V8si4x8mX6
vceE3ib9qCUi1JUqlQWc96CxxsoHHQUWbGbLeeLUlj4+czlh9+M5fLxCIKEceHQQbNLlBLF8YREZ
FSs5qPt1aBOk1bctyhAhdZxPejdJjVbfXdsBj7EJGZHryCxmuOkfbnh0XwiEAOoSbktLh5qoXHsW
+92MJjQi30Jg7IElcSsb2i0cM8kqw70HrammjOolni2G25giYm6HyptVhm3Pa3TlbiCnOk94YL+Y
ogccQZg9A2i6ArTGhmjzrH17g6s7PL9ujylYxCjHkQEWHM7XO16tpThI+cgRgctFH9pl1HhzrU/H
2TIpHzH+nXifUJ7i02p49tceypk2ujjnTU24gOAOUObrK05RHheYkRZZJB5xm3ghQ084uBq8RYi/
DVR/oeWzhWrAs7MIa8rjDi6dOo2dWLnfjxCQsxj82qYaHTuZuYJHGBxVZSS784tx8KNz/keeiB39
ebmrkxD4qHfZZ7HoM91Rt6eqk6UIaB5jmXFXyOC2QU9H3T+tSGLmfO5SCe8kYYo3cPwW5RTEYNDx
MI/+kd5o1SJtVMRNln/WKSVvPh6esVm84JaZ/27W+3pScrlfEpB/oHShMGERJ2lb0XZ1DLefNkRv
hG178n/FcrKl/B4CY4Vfi+jmImhkCoNoZr3Rca+l617nOGBwdkUMJgYWCPOY25CT4pGeKtqHNrfo
O2M7yPR+KPZa8yrGjNrUtprpr4TfbFArLyMz1Kval5xtOQVW0Mtcc/ZmT9d2bdqPZlEFy85Tc/6U
es//Vk/wV5OmFilFWKDw9VFG5fBktsAIdoj/Iyv4r3JAr3qzLul4nknZwslD4freBUXtZtRMXtT8
+1RcdJx3CvRPUefbJIiF/OZFbDqjtuEsVU5tV2TJ0FNhg2D2LkL8GBLNDuFjmsR1w2MTOZDs4KZI
TRSMdm8/IW7eD0zN6kNwCAOg1gKIIB9xv0n9iS/0Ja66wQEpcealtWC+RiKyki+rlxEgDwcFkHaB
0YC9onid1H0RHsFIOQ3v9Br66AqNoTRMmrKzZLca1RfFNZiOeFpC2UKUcCl1HCR+PFHcBTa6yVEb
RFdcDo2PLeR2EY4w4t3YqAS+84sdqPK41z/P7ZiiH6xQDpMMcPKeq0G1cEhUHVHOgA9NdeJ5l0GQ
EQbCkiSKNptOPcPvsc7WG+pgGX6Y91eRkQsqiqEltpPUKuGKzcMUz1SkS3EfuMhA+9O7xSQ6citx
8I2cOPykT2fWHG+jo/PjIItBh55fP/IUyQrA4FRhSJj1JJogqCdm7QSB7qGZgumRPv6bAXfVI9l5
dp+a0c9GefPwmfuXj6lscRSgBj4tCwdKQD1hpTgnJhU7NNs6UBsWW6hhzjdcfByPZn1ZoRkctvq/
tGWfvdZQHnqSSE2nLFtYQbV302e8S8ffSPGbdv1XVhO67WSFcCrlz0UvA14FTm0IcQw25EFnbPct
U5HiiLPEFsLZiiCMV1eq1Fp9ab5VdnhWAyy1r46jkT3PbULX25fuGmV6AMy2idifxORm9ekqBfZQ
B82AoswauXwoaj5TQ+FLJc9cAO6EeNKIXWe6aEIMBu2jPJ3ziDxDUJj7gHXBqyJwCkw1PW0H6iiG
lExqXSywwIWAJwE9HPrNT+Pew8c6SiC+T5Wp8WMpf89g4GBqHIIcR6dwI802ycqYL7dKjj79R7bn
3z2NMpwB6BGbxhoATeK6+nkrUiwBy+1kNWsycAzx3Zwf0sr/u9zx1wsTsIvLfMapiQK0fhbro/MB
9acylOGEBVydqKOTSEWu81nz2/j3wICchL1Opc8qUfcxYm8Fg7CBbA5saDsc3lAonUIfc+XPYUm0
bWB7N5Bfjyhjzndk0vGkCbU4Sm56s1teJ2zhSXc0N+0ddu81iTwboh5y34wnyrwW4tEEW2CQ35w5
ytT0mmB9jOFtkXBSOU9h02dwzS6fJOdufmc06eFHHIfkHRBbkLSVjssH2Rbx+lq2citSUcp5rbdu
9b4+JCLbF329NE9I6X7LvTgrsAHqeOQLvpiS9AOOGcTJWoXvJWRjhxsi931dzt19pRnix6hiaOrZ
jmfiRPXYIiFBVJC6KsbCDNarUVwyccx1wF8ghLaQkhsS54qRBFDmZSu1T9S/k3hrGx775Evh5Xi7
4O90vVT7Cl/9bN5LfU9AMSQ9UHRApgHiZ8lP5m/tR1dMqMPvylWQsGq6HhqPp7jrZ2cXPwOy7wCZ
g2RUgwPnOZxf6YsRBKO8lHuYv2ha5yhvB9HRI+Rt0/6oC+mTtoq1F46H/Xjp29wpucTrxnT2PclU
i6ICvaSqhcJOFnjwm2qZuFApEc4kYbgmsVN9j+4ej0Gr6Z4dWzGFRuylCsy9xXDVzjEc9Ia45w03
BQGd/Uawu6Uz+dlsnrtA8vzH1zLlUCHDSYLYyP3uqUQAI182A9taFXycid49XcF08OfxiuUTDpgf
gnqzuxPOMpz7hvXrzRouTXnMkId8zkovRWGoTsWMLf8FPNWVee90TTx/JfsD78Lv/ujs8jrZSwNY
TzgfCmx59WCkFK+sOHDWwYjmLlMlWNbAGX8sJrcShu1WAo0paXcYSp3Li1J9gZwqXk+VXRE81NwK
MBoMl+vzVGScV4qgTLKwa6Jjc2T4/awiqvUc4/YAW8cjTAa6C+3/GccCxCUqA7nwI6uFiURl+s++
tkg6pFBI2wRrjBUfhwq7QToo9bePAOxv8Y2ioOdmY5Ukayh2r3UDExpgUHbOV/AgbJ3+VL9UMHHl
LLe+sB+rF/ixxIPe7TssbbyiF2g/cg1+HlB7BRTDzbCqaGoaq4+TNXr4dxlFjhbfNa+iIiAw3Yi/
lkNGlmXTNalWs6jExYMI0YGROngxhEGIAhW6jzzu0HdkxGcDzzR+tLRKCwecCmtMiBt05EopHf8T
nCEjqzq3XqHU84G7lVPYe7BXqvKEGraxBlHIBAIG5/U+8WKehgBNs72KyZW74Ah7C17/CVsmCOw7
zhOzhjo3rfPYmPnH7X4O+jXc8iRX9SEKt8tEPsabvB2ye4tQq8KoNRzun48eOXaccB7Ux2eLqCX2
c2Fn5Vq1aqgZBCTcQfn8TAuuQlinsOF4krv7xoNY54erBUBhw51Mv4cUd0s1du9Lzj0pI0c68JIz
w9dWbaIaqEISz5ZyN2m+5nUWcCaN4WtANoP5SZTLQleQmruU59h6XhZt4AjCd3beTkQfgd5p/r8A
uoz2q58MQstjDfGcpayV1BCZD7C8OuEtKbHPm8ESm+Q1OWjgt/wrcAWSQRKIgw9xYos94z/4Aaa5
JyFQpA/4yxe0y9v3TsWFZQydmVIdJuXH7sNAjOVO68wvuEqXQT+rXV+OaacLGThB6yD3YazcYCFR
61qwXe0ZItYZpOxhNG+50uNKZB+P5YXmicSdwrmGL3gAWFrIiGpmJwyIxyhHvC2/FlZ2KsjSE4J4
lsfS/fUPoiZEq616mldeIaQeJ2UiIr6vLgCwKZtC7x9sTCeEy/xGKEZathzxBocRsmRUCpedYbKn
EjLaRwzln3xz3o6NwPK2JwvE1R/2AvN8TnXR+H1iABFNbxTV24zo29jzAJ+QVKy6kwJuIvvDtyov
wDjy/LLkJ8rS2PtQU/V5Zj/HoCVvDVu8syZOgSn1wrLbFwa/KDPsH5gpq5h5CvtqCJNPpNJLCBPO
gBtGMXQVGDQnUaXa2YEwc2w6lsW1IMjYf79C8AT7jXmE3/DPABAR6q1zEm8lkAM1wOP7N+tH5v/I
rqdGlOK3Qlj/DLR+pFrz7OD1t0wUcAoDqEebRCdl7tIAW2uexw/3AYcWekZsTuMXbVG17TypONH/
IezLqwD8JySJqTnq5YW9I8cHoc81ELhzW1+/JBUMctdXvDawkVwtWZqEcJcdNrHoqNcEFpDDzoN+
P7bG1Hc/Qg4uHO2smHzU6GHpf+kbPzpwd5UIdR44/WquOjkPTWdK0GI5EbHw/oDRUv+NeNq2Yq/U
5J0fstLsPWbsCF6vxaCPvehfwSQw5tDf8Gf2oYxCaql316CLKFDmj6zDTvJcDvtAcdq4LGHROy3b
7id1dUog44MDExo/pLvCq0WMXuR5LcMB3HXjdMzsI9dXlPI1GTHx/G+uOvtsVA1LktXderftTM7v
vgmuq678Kpeh2k7UiLVqQIs228jVRJTuXlr4XKEvzavma/q1InRxdAZTiX3rFcKL/oRRHPlZN8J+
TPi8G6By+N/yUu+IvdRaGwmpCtGdsdzdEha0TeAj68fOmM2y/XTlBqMS+cktqJIk73wh1K9P032v
XcxSlWSfOF0+cUrtC3OSsRagSvlbT5EMLp4GKvSLegE+kPo/+Y6HNOxvswly9OfICp+U3gTtYQC/
CAgGxlZuHCEAjUrBwNtV7b6THgEVYvBd1qdfBcG2ReP0b75MUnIL19S1Qd96tUch9iRsm31TqbpO
7eeHtOel8chvQ1LeZhb3Q54jO7pHobCjhvc7DGIQGU0Le1mQgpjiyiJBpAMgJgP9DpwOtqdPdI9S
degiInSlT1tRW/9Ti79GneT6kgeQAoIRYhOWSDWHkwwGDkgD9HPL4ahOZVC4lKsI9vCqT/qdWvGb
pTLI7XwVSwSsKbjhKyMNFUFa7mhd2EiF8oPEsBWQYhFFXajHTxhDDze/h8pFg7cw4N+b3hpGqdPZ
R2wnuFTwhJ7AI2xslR8u9WjicoRICz6kdKh1NTaG7xxQ6B29iePSjiUkCA3n9EZ3mazqsSqhA/+g
PL8WRWZIw6Uh4Ffexchg/GtNLUV3H8SpWGTVSuKxRrHEUSH5VX5VVTF2OUD7eFgX+O216jRFpe5/
0Lfo5mmH6qXM7dGRJPQiMvnPHjfBvJ4rcJQ7wKj4zhHTmPRB0JLx9xMgcAH+W7eRv84thEU8+M/K
iqH/+v3w/GjgAmWv4jfR+Yb2T32cjh94Nmog4bQsTqQwTlOxyM4iKnHY0ZW0IZLgZjIR8a9U8SOp
I+kt5HkxW39REao0tJ8h3ypxDrJAdVNlH0eSW77rUhgAqWb16sRXqC+XN/4cbL1kn4m66AUyBqJZ
ZFMvGjgWoRWNI1GqvFiafr9TTcGJTlZZkfNCApGB8PLbj4W4YVIdY20es8MvX3OwZJXLsqT6asz+
XlV1nTW0zjsNMX8MOZmbakIJXl1pFd7c/rtwsigzJbqTrj15n61Ac7zf8ZORnLVli/99W2A08SVA
iHzb41HgOXK0MPlJ9KIq43V+IsCNY8tCGlzPnBFjxw/2eaYGpvSQd6tSgD6KpssLbyUSH+jOwzF4
Lz36+V2LOp8c4hJASUROGy+HQ7mF+PjbupqB5QXnz9j09LlXHZ0c/ffzQljbtWI9FlWjGdJ6lztD
inGa43C14tBXhlKDoNNM4N1Wy5Oo7EAjpnXFDBKdiBuVhE01fhFO5ikp+kfsbW2oYTIhlxcwsUsv
9GjRm3xuGH68MKXqOO+N5cwf9J56qFA1ZliuqWqW7mYmVCkoWDOnz1EJoZofnH0dghh1AlrCKl/4
vXmcLEx4FBnX6vUYMBD0G6FKsW6GTGU77+XRqiYt7JfOdFF+KuTrw6+wWgB4mJqsnAQ6i87WoKDb
4p2PKY9htUb9gECYcGYCPujl7KGzy5F3LFO/l1Xl3DxHQfqurFOODu/zC2BMa/UdJ33qXchms1eh
wltIO/tw578XdQiSbj5O0hSQT637/RzvuSo5bc5ONIZyIODA8HoMdIBDP+udXAphORe+C5ZRMJzm
v7Uizu2DgCoFf6cIgyt72boRS2HA2ydTRKfhEMt9mc+B7DwV8LExtHpCpjVPYFCKGO4ZfSAMYG7O
Cvu2iWLHrArHldlknwUVN1GQRY19S1+xguXuz9BM3OKZ12mOeUatOWSaUnXFy0CfTLeS+WyHDpkz
mtFt0At2smCNmDR4E3Nyb1Yp3v5PQ0B5IN9faerPWkoOB5xMYnJZFUiNdwhsQRJifmYPcWf2JyjK
OyWLJC1zPHFdFLDUT+u/UK8LMUyZEzzEM/9qarxmEopRy5LfcZXxEpZpmey8C6xY4p0YZcyB6C56
x0ou+NMDgrY65l6kPAtXEeJBnKBcR/GcUpb7j9+uXdTdTZ4cgCcdLiN2bH0pVkLYu/FUM9iqo1ft
2CM478Ez+ScFTss+lqSWM7Kqac0JAMImQAIvDrZbJqB8mIIT3BJZ6rymNpYvcULQPvPDwwdQOUxc
CoF516C2ryE9urGkfLI1gIjZqmDjbEB8L5MTIp8gvEz+0akpH/WTZzOqYFWJ6nI6db+vrtZCfSNq
EcxiSrSKofyPhAscJAnbXGt3ey9jpt6uxzLja7RYybI+H+rUebfL743kY9CuQfMD0jz5Kv9n6jqM
22rKhKjOkORRsodLeUVRf5cSf18MkuhJYp5dORqTmmUuePD+jqlHioVjGATFhwxDwWNKyvgV/cZB
dQU7GcOGThOILOrqn2zqovhdlyJ4qcV+cUeW/RR0Tfq7kNAPWTUJ+OC4ppHlShGeOHrJJy4+hHmf
UWrs3mHcwbtRS+AxoVM5Kg1d6/9pono2bavhiEeEmzYue6WWDTbz4AZgpTAE9EVHrvcaXqiX5EDT
GB8d/uOi6JArne8h/7rQmxCZ0RrZYYsnTY65ElVPwt3IjOQY2EijURBdZy/ghze0ivmD6ssIeQcg
eWVNz8i+sOm/QNSACyyV0yAKTH+MaB0q9aMKfEunIAV4nE+3IsDUYO1sLNu8Np1HjJk4PCqgpqfQ
gXytoVCXZiMoVd9I//jpdrUhuC3xQWrc//1FY1PyFFK7bhHn5whor5bhTHHvGQ0CADsN3UkPrSTz
5cC/4hj0yfo9c8ZEzz3md5HkHzLWUx0KxgQ0VN5pzQAjHC4wRjqy4HNbnNWoFcO6LNlAiaB9CbmS
gjL33JWBdWHTfKpTvr6mZTC9GClWIU74hhOPmXcYoMnsbjQjnfCYhVh6u8uvrAd0ra5hdK0gf1bp
TeWVYO1jhr5/45OvcSiA8GKbEddzjURiOmN0wgVCEHkg0OsCjJWsiaoSe4pDJvKvSCvwXw+x8I7/
xjtlI7QuRVzPCNzIapdX+NBQ8FVSru7A/obbTc2KN5Cc3Fbqi3YYmCxhu+hNBe6oWmCpHodCZ4kS
f/CqYrPPFKpRz2r4qHiHbxYPK8CPYFrXXyOHn4EXkPQjt3WSBf+ipfSscDOoy6ujIHkm+quqqcW0
Msz85mNpT9trfFb0WDCKIrXCD9nDluxJIISHRnwqTTQeitYPrNFcUZVrlGYwVbzUSfLbyngM/10i
96vGFKhRlpVOIx0EMoA5ozpG+CjopU7uU3kwSf0J7jyUiIn1a1xm4S+67u/35kRZFw/QVue3nBFd
9Lg+33YwWGq1hij3lAc33+Ehmoj5Dhqrep3egmjxpU8WyVOnQQLVFIc24T1CB3TvSArh3FiJHj2m
rhqjYR3afB7YjrFOJVr9yHQ7Ua7XSRLdRaFhPkmLDmP2z2m54N9ESyUEupyJPsTLvXftmPTcecqg
ToEregF7PH7fZJ5blYur0oIH9RrhWqQmOo33xCl4MkxDcCROFQitX1DP9r86s6AIKA33mZBKwAMa
9fMlVNDlAhxcOfJ0gavRqNQZfZdlw+nlBxt0U4K+6fS/9I7s1uNfinkh9zIXMpZVPUGUgPTLJ6kL
ke6AfMJCUaGsK62QYGV72xDKgA/2a3cRi3yMGQ6SxG9RbaEFbFh09tmFlsSUsfDWhu6EkO421LNq
tF6xgbcXYriWk8WtUqtf57USg8kM80igq0xhliyYs5TuR4Lm7cysYpYmPvQxPgwzdrduXfsUxe+/
cxLjhjl3Bx5yHsS/2swgq7ZfQAvmQ02jYItmGBHWznScRde+4F8zlnYOfwsUmMCpXxX5usZpaSpq
W3aTMcZxu+slHxkLXoCCKhJp94hPWlDbgdzaq5EgkAw58gVHiAGpzo0ogNZLLii0BVbRHuqD5FC2
w65GqHO9TshRrv51ycDdWBL3eXdblLTwVNcbPbQgYpM4sXZwiZYkFTfpxfqL3qgobZ7B6fnvQr0d
/H+zxswyPcWx5ovYS3NdbZMzJx9pZxzCbM+zoBvH4eszbSCrnjadJWHEOfi8zJsvanIgdRZ3Cd23
cqWLuwK572/d1lY3NZ1mu/pwT3L+MBQAaLr3pcuripLVP7OJkEbbviKNitrGQ5JIqb3YWlfCkK5M
T7a7T0zkHM4hoSwgG5u8ucZXkBKba1z4bF3MwJqjG50GiQXQy+lzNwXN+fMTOA6o6P/5zT0B4LQl
Tk/1KQe7sFzWWxEprvKun9JMj07ng9iT9tkrwvTuLrp31ovosJAzs8qJI1gqcAoSmKc56qRs3//5
BG8hHeLIFhjhdY8CkFHKcOr8qW0dL1nt7e62l22bzGicVZht92KlxYOGL3ygh1JexQCnYWYbwTN9
TdSHS1s41wKVpi2W6b1jOD/FyUEU6XyiTxu19We7iQybtU3OLPQyu9xBiahd46wsfByY7aLh8VNQ
kEHvZA7RytZD0vMNa5M7tZ45PH/IME7bpIER0T9bUTX7n2oL4ZUHWDjR/EQyte0YZL3iEgiMQvw6
9l2lUuqn3U0VRM8f4tFttYDA/Aoid2i7m3LcptULy0wvBDqAekUGC4Hfy8U8Z0Dfj1348vGtmp3U
2t3QUOmeTIONXVBB+QLNnJwYbG477XQxHKDdsBpzvugh0tJG0gRrfIZGGq9erfwlIjRAqdpe/dcC
1au5xVu42sIgSnhTcO4nPTd0mAmrhMDsv+WbWOwvOub2r6xZ4q/DiA7dHmTBW5BfE9WMZ/DgGIqu
UxG0WChA8+Xdnpa4/bgTRjmYTKnT4rLk56CpBaihz4JsSqTHnbB8EuW9GakBMlH0RpieGbWZX/gi
yOXepKSNzhr7Nlum/s6WCaX4986DcPUikgpLZJiR8iQ7DdDU/N4ovjEPJ3BXX6Xjr21//6tol0XT
tUkYaXpB+4VWhCIvpgr/6SeIH3URkyWBR+yzn3gf6THjfkcgaK60T5U0Le2izZnoaZ4DZZAaZSaM
cwGILi3yZXoP+fmQIT9KUTHdb8wHWwERr8iZeLuALTP7ogOE8trG024UYQmOh65CeQn7dntgWnO2
Fgw68s9f2kvN05DAUx40X/FHFapXhldEhkZbQT2T+tQVr2s34X+5zx8wyCgw+waZl4BLZuzNk4cn
jWgsHB376lXGFbC4R0LKYDpV42YkDoHwvxmlNqMx40qgzcmxxlesbZw1U6epvOPnBTv2/CXVHlh9
NZ8A3HolXBxoht2LOACmQ6othy9zJKWnB6/ZWFZsKrGvfS2axUBppoAXa58IzIUovT+PfLGiCmY7
rMfRdY08dViO0c9s0IbGVJshSKjiH3jRCZOL2OhsT11gEGaMVL5p77y4RCCmW5bFzVQh9N3hEa/F
gqI6ycVYD2Y8CT3xWUpsVvvK0NijOwenlHoUnSHxarI5y0ZbwhfmzT8Rd4VfsC5DBPdbySayeEQE
+Zd7kI+Svveem0Rc+pF611svjJ7YbeFnA5YeuPHk/ZrrrhprLqyIUqXTkhOhUsBmauszBrI4w29T
P9vSOcQ0wk6ax2i9CQbc2RWi1bhvJnE+ott+dYHpi/3MzScNgiVDyjMBW+ldkcVSGX6bvzoT2uP9
DhxKBwu8I+tM+27wmDEKGODvE2pfJfs9LKGLOaY3s+8pqQdTDZU8RknmJhlhvlaw2Lq9ZW/wE37w
Owo4j6UVDDKa4PLPY+gi1PdzqklSd53AmLGK5EEXMmXZjRfefYnu9Mn0aTEkZsSuA75WXJC9J0He
u0xnBeDn1xBxJZXaAS6uKB4bBxBy597sBMBVqj/w6cay2HNUZiOP0yeAuKo+NGHiNnq0U54Dc2cv
Si0h5QSpAZojxeiuPevqJ97X+Gsxglq8qi1zgZYZ94UgVkxshwWk8IaP74xfvNt4vH/dS+6sIhuV
nZDBuXiWLqNC7kxLycaJ1YwlSJjnYzLvNytqEu61Bm6NmW6NiPzl26qzsU/yxsgLofLyJYuzf2Sp
/b7S7zUILKYTM6m32+UemmUaUps8yVGJfzJToz07qhLy3kqyW7bLpTZn7HR+QisLqcmYL9dNmHHX
0xcyKOlG8eMSqcIDySd3rzU+PMWnLEpY96yfSfBmwxYZWmycssFvk5kTZORtx5RGWg4Lo7BAKga1
en5GJpYshrbiYdIp3V4/W7Vo70M/TO8mgYbb1abxkY9oRj3DEASzYSuGId8IUjVf3tXffZYTt2v7
UlkPBrXI7yghj2EhLG1zrHAxjfinXg5D6N5++kjzQ8c/rRLBs/MVAQR3uWoXbIfCnc51ceo4B5LQ
/MSwvGgkrPVmeBsiIkiGXwHRWO6ntybRFBsFbm+Up49bL0JSmQpVUH3b+++YaC7O2xMbBImXyJU7
VmLwPoDNkwXf/qAUtp5a1it/6hQdL7HvoGuCTxIwFuA8ORu+XFp8+VoeP39XGwEr7A0OnafDljXd
FA3np1QG3riksDrJHlXTq+nLg3P0GrS1Xu2zALsZy1abPefgG4OViDjl8WQMDUcDGRcqqLAb3Nhv
4faW4DwD1bfSK+psGtrbDbw+Se+J9efdHytlipPLyN+Xc1mJlUdzE3tCpwYfCXiiBHiRQ5iQQcKE
aDCEAR6Imz6qJpmtNZXlyG+0gr/ZkaxdpEMPCZpzrgJ/cPcpZYech0JvbS+Cwccbuq5GOLBOK95F
8uYDCavPxNkEY9oaV2DPc0VyqItFqGy/KxGB6XwA4XvT4PpYAJzQd8HZRv6IDcizIDW3aWqzz9cJ
TIu75DgiymGZ/VLHPqnzvjzS4wH/tTOMqiz384ghiD/xS+dKi5T3kFgw+weZMyWD0GNb4+cM90HP
LVnkCZGhOln53T+ziStcNdP1ZHCAULDT1YXZi5tJQPsyAH1CX9Ac4Vv/KKs+THgFV3yRzLDdIt0b
xSbW/oP35ZFwpcPTqKy53pOHPj3eYlw7yZ2q0D5LGHAzJJK4xFC/M42HE+01ya2OffAK78t0j5EX
uso7fAo9cimyD4IgJwtY0im/5xqmtXVXVEASrR/c2sduZRAI2AybbPd1wsYgTHQTVUr+pgXvCxk4
6M81x6iOKH+AY6ICU8GWQKOtaK47FLnxpqZHCDiTpG1uhUl3TrJmWS30COrXk4ibR4VypzNjpWFN
d73UOX6jJyE8r8xzDiE3OqSViKQRmPGq2mOxnBBeFgzkcFzrOtGOfW1xrIsW5rfUDTC+KH+/p91p
z+CrZnmw0PJsuVpnvsljWtsazkKj1I6ega+IuQEamYKDsR4943j/Z4v4kVWweLPIdK2FW/a71zhL
lngCigqAJR8Opn9/DcArtPMnCNCd78K4p+gL1g+QOnB7VX9F0m2XpC+JOzL/9SGSEeqy984gTRQW
7tY4Obc1H+uO9GROz26QdPh2jha/K2JEsJAIY4/UdQEEzPJ8zqf0zhHhXGIqHriYt+8zWZCB1CMz
TPOWxwqk0ljSoSqK5v/jlhFhliYabD67Zfjqc+Y37M5KzwLlPK3fGSSJEnwDrMbp98ddQGVhrpGL
dH4QGmjFISRcdpNj5eIUKQ27yk/CcGM6wz3UV6f3UUwZPyjp8Nb7Pn4TToyXeliRZBV7rEld/j+5
NczMtBlT5d85OBuFoKQE8JtRbB0efyXgcczoklBlPbCNFVVgqb6+HrynOoYgwTX/HUVV2pC20geR
ZjoQWp0QM11qbtsQT5Gi+WyDTpcO1oBgjTDxyIkyBRKYsIi7Gu3REITOcAD7TQrye3XvHPzZ7hEY
cPk8IJvVY7OAZeL/wCnb23jW/Vqu+EEK1XBwj/lgkhcvRHOgMQjDIPhL/63neNlswREc3HbTz4t2
R93K0eE0X5aljc93NQYnGjWBpjtJ9ZqihLtnOwHf6kgqIkYsVydLz5PjB+FYEdgB/b/mgFS6Qu49
iYkkpVJMw2bRXz8RecsUhZ/kAwP/DZb7LZPaEb053ZhA61sVmJ8+HLLLwdFZojkSsC4fWp9jxg8C
umMH4eoHww8ErFGNNt2MzapHuQiJu9At67W9DXuZA4TH78uKnd3uneDn/JOnvtLHXjXwp6/ZF+uZ
eceYV73PjKPgvgfWYWsw57D43Olxy0wdchWZREN0qvbrc3aA1j8S/sWA5oYG53zZfUllBClha72G
TiS3I3ooPndZP5W8BrIDR2QaadjexuMniv+Enbuc74iLNxTHCFnfDGeOxOXku9Zj3xM8zmoplyZP
3aLGS0XGVojTuMF0QPeMOMsOkY36lR/G39/GvDt2ou3Rk9y2xHzTO10yB67RzabBJzuaCwbEKnHA
DE39lcJmb9yIFzExe9LdoOh/0rpRTY9L4OUdZUkw10MnMA6F4FXULzR75Ucp9ZnizKrC3x86Df/N
oPTAM+cCFc/XWu5QpG2cuBlygVsjG0lbPPcLLP+9EoEniDSyK/JMiuNARyhQ4BIkE6Blq6MDWBb8
N6rvp/8XNkx53wNyjP+ypqv9Wru/q+ATzPVQog5LIaFRNI/qqlRkWLDvICt1a0wLAay73vB7cdAR
5nOyL2XGQV74TR7IDHOFFD2hCBTaol6WJ4B8w2YYNbsTELygdAJ2YN2IxNYE6oBNm+TQJk8WJS9B
gBsOf2+JTWLOgiYytKY0GAKLSoyb8dTM5hQMTpdOB9nR3dH5MM+nMFGgcGzNk/wajhvQ1Juc+1M6
eBFFjU7sJZZ+ePR/+UQmTnO8PwArFSKn/6wMgE8JGNl5+Hcx1JalnBTE6DqI4GKOMrXcsHspX2uJ
gBVKw/NXRfbvwkGXi3I2VuHpOXjzH3qYfioei8Tz5jbbehMYH3y51FS2AydXoFKMOEG3c9Chro29
ACz1TODQSeJdHPEk6JsoXFncXlXbb8/K9SqWuzKbSNnVtbJ31x8ZsxbSl7Yf5r9GuLeQ7e6t3CZE
3sQIl0VyQTDSUU2GTyqqD7HrzoSGuEV0Ywe2INJk5O8j0Llhazs1fVEx7KN57ooX6R1f/ADPKAFb
8QxkdTkHAmmoeOSOHZqCcZ5yM3bKKEPePZr80CZYyUGLKmfLtbzVhttLjdm8aPmYWwkM/XagY4Id
wbz9OcnihILHLdI4HdbU6eGM96YZRsdXSxCI8Cy9I0AY7EGrnWVoca7DL6CXtPu+R9W2lWhSN48c
44OSj604SWCuLurV7sobWDxB2ywW8YUAJaqCe+9sINYQKlsaeuZJNl7w8P8VTsfFFL4pDoHzZ3iq
Tpc1d/E++CNdTYUz5K6cQTEJC3OTnuU8UXRUpruej0DGCDsDfgY3w0FSzp6/JtMJAEkKQc6GVBcv
wGUddXclN+TP1ZymA8qYU+2ZbDg2v4IwPZeC8rq+yu1MTjYdwWMZTEJ1ch6iQKwREekIy5ruT3sd
u1MmiZKI9ie/BTJ9JU32RYMcunuHZDsCw8J5+pA4QCFs2BfZmXUBtiqtSVFmMsnwfppIQyLY2I6x
Iny5M2vaT+yAaHu51jXZGSyc/HYbBkjDC4Vr/6OIM2dxVkN5Myszmxx95foq2jlfaFC0KR4o+XVl
sZYnL3q7I3M+GaS7Hqhg7+bIoB85/F5vfK/MTxshD427qPzC+O2fwin1+kt7fYu+3BbknKKl0EPl
2zP6n6i1Gzt5VD4g+x8u9dNchd3eiBHuAsdBcILprO+anPkXlR3aGPH7mhwRN6TELf436g8f8JXR
QaxnrOYMBP2cLsjSlMqi0GuZ5CJWUI0NhN5WS4jV9U+NSkNzewXVQaKhdZAuQgiDFE/A90hwcbgu
kXp0/rMb4QeI7EuW3HwDAVMWCZPjU3s0WgqpPmCow+fLvzTjKm6aEt0OEzYBMmMGnz7doMq9qI4u
B1XQthngdf5LYCjYjjrHFLSVdYayE2BF6i+apoGL4qgCs+W508rdsXazz8DAkI9XdyP9Kz7rIb/c
MmkT4Vrx0MLuhfRUlj2olgaKCqOUUD/PPHRBKY0KRhFV6k3zj6YhinTs3OS9Sv3qziZIAchCPPl3
/o3/QONFAZ/JWNEVS3QeUeqUtMRxl52398bJEJz4eNAk3nMnWgoeT6U0npkysT5sChuapQEMiimI
UdmcGjhoSfDLSx71VWvJ0Xv7QhSFUZsNzOzdb7WW7vPboVeeCVMPL9Xi+DlbQAN/mavctmIlWPXd
SVY3GIRbFH7W8mtXFCcuemsbgmwPtB/n/fbUwyTgn5HHDkBnAcEuOF4bgZJC4grAp7+iPv2kYZiR
6WGv2Rm0uUi+SQ/Z0raMtJIBgAKYJXtivS8cCTXOjPUwx1tMp6Uqx87M4usOsex31ulEBb3ZesnB
yYUK9G6xUKgav2eSNDbNNqBrfboE/AQKSbRmGjg3ozAFfAubX3OF0GiZhEkFTj8gTPDxpYo8B00d
kawnZa5gJfDxOKmzfpQjhmwvIdHp+2LESnlrGd5ea75ifumXRRTgVZ5u+CCF1HsVNpFpdQ5qS54y
TmuLNIjHDSOvq7IiHOS7YDWk8VC42IWDqjPQe8oZUwmHa3PubKqbxaMtRh6n2bOcG0UJCpQtzi0c
p9XiP46QqKzLKgM46vQ/AzxiwMw5XEJ8a4Emx1kIgUbReZJ63AyR7U0vnrnFjZgE5CijDyLQ/zYz
ARj6Ux9lZCLOff48MJh4p1Geo7dDyyy3zAsJSN/0W+RQVdZoQiMQjjcMjXWnk2S8L7B6vwRWZ07S
QAomJDZlf1yupiaE52Y8/VLJr9f3XH2FgxPljlvLQRQn5AF31NXFi+1lgE5hjDXK1W2fkHVW3kHk
1aU9RMQHvGeWPIxrE51ivOgRC80eU3kcdjzhdukW3SggIp8TrA29dQeN2hvNPGYVyhI8qhZMKA/f
XfRTPG36Z/T/NZL3makN1bPCIK54DAIEoYgcZPLtMjLPPXLcgV6A1bgadMgxjzD/GJQg/yzSwhxC
rjxeo6EW1cAX6BZfI8f71gLnfb0Q4JRPoKccSm1zunl0H+gTMvM0lgpKnE0Uor3UT27EsC+KoWes
DGqKxuzyY9HoQYntfMXZYmfyrTnDK8LifYPzkQWEhZm3KBnPccLl1RAm3zvU3NPuNHuiuJAMNyXw
yqFdXy62mrhFp03cEXvuW2o3cC1glf+o5UefODPbeT0G9Pi17Al4vn3UlTP/9l/9pSc3Dmq/sNfJ
9k/Yj0AUfcJmXffqcZGpR3G7lAzGkX2xS8oXdaMd64v6wikVEh9Qn6fpr1J2apWN2qpS2h/eR4U0
pCaiWQilaCH4eT/V9PaCVn0UplQjQmWqDqHxjX/K1Ucpf1gNnA6Mnv6JqH09X4pXWx2YpmtDmN1U
4jNjut3TW1tOye6+I/SCRwVRveBsZIk87iuDPvo7UFv/F46GFZyw25PoHMPkFH9MCXlirelYIjbN
dvcKrx692uJMfG/mKMUN4A/FRUmfsR1KQ71sMN5xAohXQ8BNlSNqQsbJjJLZTOnImYa3GcYG8f50
yfetKLOhYz4bxHHFZHy5qFwSSC1I82KNGa82DGU+bI+k3ZXmyyD0GE7Q6OTugRLBbeWwKSifJraY
Uz9lzz4AbIF+0JuBYcOLeg49uMQzhCk+0ajoHMAy3dYtdanZg9zhSvmmHc6elOvvNZkrH5jtr5W1
jhhc18z70uYXpCX28vCnkiD/kzO4es558QyJndp5p4egq3rOck9b9nYCnPGfWNlIds3W6mUG+42z
HBOX17rsR06SQU7tBua14WOL0hb2LZTYxtPlO9XQjFWrKNIAJ2pH9jHaCL6gUlUlZK/mUiPgcGeo
b6eYBeL0Y54wFATCHKauxmtOAf6RbSorzddkxG9SE8f0yWsEpLgJ7JOCkAW8YZ7NXpBC2pOJvcbd
dOjUloM3JPJ0p1wLjH9GA5ASd0kxDql1wMjVj3E1nY9w0RGoksjOAJLhLsWxeZrykYYMX+XQISMc
1uShq91MYb8EyI4yzcsfwwg6RsH6Ce58EzWG5WEPsJtHVK3cUM1ASJMl/eBw466ms1cq1ipXwEMp
suMYr9bIccYs8tFFg9m+9VZQMZ/rxQXZj8Q0iYmQVxqjH7xlKxVT0Z2LIDsuE/M1CqqtKSiBVGqz
XkD1ba4eBmZDOExuULsiwyqo0BvMvuFCEwKI+TEASG6SNpxbitpH2tnhbPPFQTcaTj0jej8y6rs0
XLGjLFhO/KMmp8eAS/L8L7buYoC+6RTiXKUqzlfwEZFrCp/np05Exb/IOC5KFw/BvTxPBtb6N6mY
rRsJCFM1ZLET8pyaJBxstRMKxfxLKKtPIzw/u0r8JZuihKt5Jt8fQMgyCxH3nhd249oDAkwT23w8
96CcOyG7DiWy6WsPrI0s2RR7My7TDUVuz+yGrHXJPQdGE+2DAGfOH75//P8j4t5+RPnlOLAOq5ju
HaFTRvAadvNz5gd4WQx4PqjoUV0qBhasRrf6yQKnvoq5w8X/MdF6RPCinhsS7V1ysUCrZzyC/ICt
YznpQvWuEcrF4H3hRwNqfU8SlFD5/lDa0hrzZlh3fyBD8eaLbIOc7cNKlYYROmTTlpdymauaXpUz
UlsmjU5lS+Tq5N4n6NITHFLqUoFU8i0PfGzGp0l3XyT3LzH9coPX9kW3kZui0130Wn4jeDJbB3RK
kzW5Xe2/z/jUW3g7H2PGD3hmFM0wvxzAJiyc0wbU5B3TXVZfDfzPacOsjD/Q6Q6S46E3NvdXXkWO
HfZdgFmvCPSEJ+xInOuweI4Xw904+RfGJtWaNNZHaFDbVux0gEMu1kz5cgyvKN6j2xHhngJp/WcT
aZ6gJLpDsQ2HvxGqXhnMowMceAbAsqSmUjSXyq5Op2GId6Umao9toaJrUj1WEoTE4UskwXFXfOvE
GbSQjE1QaV4RrKv5fH3gJERNPl9+p2qPwxwlWkcsioh5gIY8R3R8YP9HOlowjY7mFf9nv99+VlnX
qgQ+SJZDwI8jZ3OJ9Zotdg2EuT1p74ofS0vu423j3BzbII4//4xgbpkZhGO24B5kNgYRVmwTalMo
a6sn7qcSu1NPsV9DiA3MWR8bWIaPOGcnOXHTpBvvYiLN2SzomOJG8LeWP+LEGBtaYvoZaQIUXAn4
44NEEKSAy7b83eXdbh99onpVyzeTjutq3or2SRvA8IhRfsi887Q3OT0l9naBVw1zXZDsEN9ViJPb
XXd24Kd10w5EAAYIAUzKnxYkPcxIO1drhUJfftLKbNamuYf24NJnmnybv0+18fIeNu/+SuID/WCs
bUaWYDO/jrjcfVu/YSlxDAwA69kv/4FWvoQ1BT0YR6Asx5MKMJndylsEoWyAHQvR7II9s3WKm4M+
k/SLM+1NvV7EM9CzNBsYBct+4Te2NaANMqeYmw5CzUA0XCNrNBY+Qqtdi5el3Xc+eN1hF5mkTLuh
p56fzv/Kyo3k5nSlYQfKe5qBapceTfOOvPAd7uiQuHogDJRP0eyO7N0krbobUU/rbF137KRyKPGJ
5hmwTPk4pUL0u8sYG8e5BCP0s6+uZJO6YY64amVwTKImXBH19i1Tc3ETCd5su9xH3pNZpm1P4J7c
evZ55bCMeGXRII4IuaSLE6YzIoVn54vBfmV6kjPmQd5wXbFlNZe4RCE9WhHbTasWUQXWgJrqZyYE
Sf90KtJqshkJmcWAkELVKsnOc6DNFH4D+6i5tFokEWIV8Zznk5ttIi1j4/96x0TF/6Iw56kT/zAO
sMtxDL1uS3spvd13MtilaB990oiXqbOdbEyQZYe/k26KchszH1ch5R9dT7qNwFaQM846qaTvYRq4
3kRGA4sy9V4jF3MQTnXp5Pvm1O3jpXzGVTVrEDZgCt1rjp0hmvpSNiVQQt5vKYAQEJNSr+E8ofRu
8HOE1CQrrb7zWxVLP+Bjl3D0BmABgUi27Xy7BOI8/hUcsEXqRkO+A6HUoj7hfn/0A1LcRF7Ul07F
XonRAkDbGVL2GkuNTcekHV7N9mLL9wZPFQDuEeGOgTuvpjBUgxuo0AtybXq9kbs8EwUFZdeG9ac6
ixWYxFUURN7KYO2Nrkw4+4MpI4RpQ2bAeFvKd1M3+NW+Qj1k6/BuugeJG8XmNUy/kvuGGW5SHPKp
HkuJuNCG7BsZxeKbRCNlca3YjGrDyRKx5Ipssb/TguIj3oc7IZj/fuKUp18Uyx6JTJc7Vw50NNkC
a7KLVjMFNqgJXT6w+Y2+m4AooXdRcJO48J+W2SQZC7RpyGzgnLyxwAzS8cg63NR0v1xb6Mqf8ET5
twkvW62vL046fsBiNNNJixg2jk2y9AiVRNbGC3DaOVjjaOoEis0yE5xBh435/qcbPdzhkVjCR+yJ
nWV7p8cPyAaS2JdMxmzw2WBZ6hQAZDy9ocY91KbPJVvIGchZRWltAGAR+iYke9N7OZNSoRnZWDpV
7YizMxeXxnBUlDr6ocZX4ZxDim1BXjZQg6hja8rcJEDAKb2hDiCIoEXr7HOcNf/HC6s0wLY6rOVa
a0sFoVSupv0lNUYsvFgdR6zeXYr8Oe2r26lY/dpdy9LlQX5rZuqfvc4XK5qLkc9tZt6lIJtofCap
UkVb2PPximAIyVs0WD55O5dvjWCFClZdfPhsT/qeWwmr94bOiq8Cvx2Q15oLM7Uuo3maJ1cauSQu
Rzv0CE6cGQYb3zLM5ng1CF4CrK+sHbKxZ0CS/cnvm8QrCitAE1DpPgmLtJa9Cn/irrS0mDQklAFz
Co6PijFizzQZmlwVB+xmtsiNFyroRqM840tdBXNZcCY3pP1qzL7Rhas2lg33QqFiMaeWYZBQetx4
Hr1IBhQgDcyyx3LdD19KIhrYNOiQhZjEJMHmf/ntomgfYRXq9kxMW+3Fkq6GM/OEpV0F/gXSAnNh
Jiw8KhSwf3s29catjTm76cBWOMlYMSlGhTKbSD1jULQqaHpjwtYSApETjoDPqLs1K2sUjEgEnugg
eqie6qo4j0Z2nDJKgEG3ATVZ3fPX2ZFrD2EWVHjsOfMlHIfYblxtJevR+fhi7tDUKeDKXGhnsC2l
3CMhGMJdtNssPpMBfrzTm8v3S8v0uTHvXgyvYInED3xTe3YL+U4iJ8dEvyk5AfpanxVQkmITwMiy
1s5Dpc3AytakqNIns/ZSzgBGxnL7mS8AF4jtiTz1FRV3mlETXI5exB2VQXY60Bi62nPcw4FpD9N7
kIQEQi+JeslPryQSRvU9mGZ/IRYyWxqPcoxbAAtPOZM80+khUkuylNqCRhlNKUOFh7nPmoKKVS73
LLYa0JldkyTK+14Vho/ZVfkDJndyiRmorw4615bvnVAukgYkAuWo62hR7/wMFC1/N43Pn8D8Zop/
PfrpjR8lhAL+RUbcYql4QtJx9kYIGF1JJOpDAiZhYoZZasdRuF1g/QCVP5n9Od3MOtuVUx4B7P5K
34wvtDM5ogrusDqEy5+bjBdAAgB4tWCvtQPgWj1xm0q7s6TC1d9+xahk+xHN3oJkHi9qt9CHCnVs
9EbEfews2cLWAjCwSUmXYfOvdrCRv2p38WD3Jd9H2ydgPka/s20CKosDFvRYzso+g5LZW7Di3NOH
l0nSEp0H4viCf0gk1lzwrJadtC2bmIX9lmgC232bfhdfmW3rGe5OGysNiWSxLiocCe5sI04KlyOe
PjZRmd1z9+ODWNFj7KVQu/yxXAadiYfmcZdRkQtYdMc7cyt1jkHhQwqpG4rzYH+ceqH6jpVcVcLI
oVsQD1xOuCPGfkNsK7VA2YTojsNJtwHwd/8uhnRRCR3sVZYLmPJ7lZK6Gc1sEer1Pt9UQ19RlnJG
0ycxMGH/MGRER+ImKnJCr0M83KeEmaUSq6ssswIkr6z0qn/crLazKF1UvZRW/QR/MJVEIVyNfhEp
HxDVw6/wB1vP64bSTRWQvKuxdMeW/vXR+9RPP0LCE+VtfZnSgswPofEtxidJeaxsSrTA7ECwoD2u
n+C5k4X4+DGeEHoTYY1MsqbD6sZ+HLu2YU+vaBmbhr3ZimLWd3wr58N/2498GIen/JDxOFz1A5te
nnjvRFiJiYjZbXCUEQrDJs/hW6y2fqa+h48QLQKEZ6/Mlp0Dgn4SJTAvwL10Y9PuS8tEIWBa7NUP
NaG/5GkO01cnzvLgCDVh6lTmzSpmyz3/gKNF16nwGVSd+hdNgCaE5IH+MCURjJthbp2sXwvP+dRW
6LNG6tFDxMoXOmAaccNTckAM1XGYnL+Zi6zp3CvMrcUKiDbNQvoL1wqrFwfoOU8nFvbWV25V3xvt
9dDoxvmsRZ1zCI7k2cyaiR84wQEh9jicxWrakKEfvtsj6/QXXvtIKhWg6Tje0NTBl59lsl7b5AYx
gWtYBtg+EH2/WtOC+Od0Uzcn/pulgpXArb7bCkkaouMpaMGVN8FVWZU5Anv31eOAYP+flTa2LXGW
LkFIKBeOAkmF9NzSNkC8urKKvsBPZf3buR0AwRVVc26A0XYLChz5JEBNjwCyDYd3k9H92zGuPWrp
GM7g7O2Nj+WtUpTHDsYSwumhDAW/iPX7Vj+loJdH7KYDdWQfTsDJjViLa1w3HcTzs7DtsFAdIOpT
2znMI3AaSoM77x3etdmF312zg9qN6gOxVJgZi7eP3SybASVibE5JOt4dHE+4m2S7INb2nXYUyWwo
x6X337Qrub/qMn/ZJEqPnsNnoyMEQH7PmmF4PYYt90qSORg0yE8C1ztPC0IaP1bRKdu+ptLXDIsh
IXF8x9/58v5IGKMzkV6bkfSvWL2aI/2m1g7+fox75NCPBWH8GB736+cDz1tKiWJJ+up0LvK+spcP
uKFFUGVXrUu1PgFIh3f8iEx+lG4IrakPq7tZ5AW3D1IXrgnvqNwJfVPLAcspGbk12PbzSoTQVw4l
DRv2Qgq/vmTUzA4xkoceD3sKaAup1hw47JTAlovaeGCq9epf7TRHe1Ihmt96XX7km9QLKyYwU6nN
J5EKm1hIaYo/BimOHHaR/tm/riJC2wvjjBTV0oX5gnMxl0UTQ94IoV3SmZycimGpGC4H/A6q8FEZ
Ej0o0ml2TsAgZUYCkbZ1FFmI+AjRgjxoF1r7ifcDgtjvYHfIU4SgdbLJWeXIN7l39lDls5ejSL+Q
vKTapplMOwn7bWAMajBgcMCQfRW73bnXapYJ/vQhFn8O6SI3wlcQSBtv2uodb0XFdcLYXG/glCw8
uzZN8mMA3TJLUw1BvpG/YEJvxxfYfxnIqTgSYamKphBe50/N+VZ9cVtAmd6hKcwvR1pM2yK8I6qj
wQe0/oDPUy4R5CunHNwWDOK7STsRgoQ5ecrpU+LxJ8tHrIS0UFstKbTHu0s20j8gWrkYsnxrObFR
OGJZery0WYIhKGno6YdnHCwVrOr1+lzXTK0i8l+BppMcjHl62oOHUGXkSuLRphY8k163BRC14uYP
oKtinPWIrDXs9XLBzhHAJvfJoVeOQZpO+YjGboMWKZ5jeh3QpT1VEzPB4dtOYTmWFBPHTaIbuQha
g6Z/01hq9ydnZnt9jxwzgJHxY6fpKxzIvsMZzjZUIgi2jLL/VZL8K/RDrb7fp68vJA5q13IKoO5o
nvZ8A5h+uCrG750yx9zK83rIPnwHhf33eQfoyDgIP+LGoxS8Bv18JNDyI88xKYKMdAKuIOy6CyP5
kMfw99FtP5E2+FbnHLGRwETgXp7P2T9t5bIPLM5UQG1etoyhQlLePeSD1Dokflkf4ZylDbmVus37
wvRe4nMv0OpnnnwA0oqh3Q8sVXFLhcqt7seRa5AlKhNO9MsEgjEaejJ60J4zfXv1qFbdxasysunz
0BZjtNiZl4d55NhxM0RVsn+n0nykE5ufcug4X/DsEfYhZa0mKS6Qo9AxnECX6zi9Ar5zuPYCSZUc
JwYIQ4s7WVxLzig7HsQ0PimvcKkUwDKRHqdwQekBfN5k9T5XBgyAXIPbWa9taePootn8dZYiDhKY
0k8mjXkxSio1MMjgRSEFeS7pxlQFW1baG5UWdYd/9IlkdqebX4XeY2lZShhgBUDQ/Y1YYoU4ALgj
VBt6xmBf4VGR7zDLPUAEk5ZX6wSIfxk/8DiFuMTvOLjhBwua29EGI7IeSQEIo8SYMxrsI4Fx0DW2
0qZlq1n/ENJjelQDYfckvC3TByvaiFFEixVGkS5sMgfaLpG6gXms8w/XzaKTkOgKnKXJp7sNvDV3
P/JQ+gfLUaqc+eI92TFrAkwjnQ1KmxtVP8Lu3Kz6q+qw9W5RtQn2GYtIm1hprJYewC4B++BOk4BD
mYIY1kRfFdkEkAfXUWiSqp5UKD+M4DkM+qdxpcTZjp9hy97q9mERyDPiEuEpRyhDd20YxfmlwUA6
VJaajR7yiKH0Qh17hDbBvI/Lon+AsXmseizDdl+3hthaEcog8uftp+b6r1EiwVWh4MIg5UL97nfh
7WydNC3rj0jkoMjhFQaCOTbP5a9PvdjpMz8+bqdnN2fNKeO551/fThYUjvqxx7FHCS3Fn8PHjicP
49ZMjdF3r+mHT9qkhJwk5GTyOGQQnAxW8UAKkJxEhZLm3b5yH4nHKWs+paMXcD8wiEX7BKWLUFTX
1UN4k0gp26icvt/8txJi8d+VjY9jGYfIqlwBV5fJ9r1bBlCqeKN2XwIKGrtqDnDgyM8c9PbU76Cp
asDKYbcurPNM/N7l9kudpgappBhznkh7RldE8GpbPc+MN+2Dv1Viz4xpdjxesnqgyBX8rDxfwTzD
2HMi/fkhHi43NGOix1q4+A1dIVqjGyuPWXsG27ilc2wxomhIigGUs3XksnIZHgKThFkkEp4BaVZ9
RoqkPpUU37hDoZojgyiAASUKzhu1204lL925PSoaxNDjQlv0IXjv+MQ7n9JXbIZ99NUMvMsP/GWx
CG8tA/gtS7HPVLY5iaLjVzqtUyMSwPMyFj0yhNtVTro/TxITo83epsJGVjgo07ubIGraYBLTRI4b
vGbNeMexxBOzoD5bpdy4/qGOmpQnyxsLb4JczPwzm86BG+YEqZfuYMPh6IlsMBKFB5L+Y7CrF6GU
fKByEEClW5PSqYRQPc09vMrrhicfzA82CIBraZtUx7K66WEQ3E5brRpHdw9LP/p0s74rHUFRTMlw
JOnERshRP3iZ2ArSQsSOZgE+Uw5NBmsn1CVg7FVDxN3CLd7gORZoKnXbxaCqVC2uIX0jjTY3b+v4
jH2+MtNhFtwGjrd6eTVl9YCbvLizT7F9oetaUA3Zj3hPIZ/wUqrx926+iudCXH0qPBEd0cZfuRkM
oVd8twRyyo1b0dCVl2nELDvJl0VM5D8ra4M68HTP5CPeoB9rHd5bxqa6bDV1/FKG5PHx3XiDamuM
M2dzZfQS/bAANNGWFdoRe7cqZNnCCztkdLHnzCpTH0/4SajPpa7dScYcg0hi3j4wR6yDqpyhEGyw
4BkdC4woGL8fXrRzX9HAogNlrQF/B+vwUHPcnYtA7VNANbzzcXPDKM8OUOBv59/fnc2KsowRDK/E
ne1HT/niLs7RushFqT2UueHlXgaEvxEu/zmSd8+qALUApFVOeMOSSqHyw8VbRwHMMURDSGyBN79m
RkqgToL6+Sk1THi37HRvosHZLul8nAVCuwMx8ftILPAoiric7Q93VcjQBWk1mlrU5XJ2URId57QC
IHPKS8SYrxJqveF82oxXySQabnPqBLWqHHENP+ok/tR8miTB91g/WhqLAzbZqSdahgW5x1KrxpaQ
tXm1xJs6LwYqqpnGipQNgbykB+IkvnP2vzkqjbX3wU6Ip7HwD+CiwOz8cZIAXqdUxjw+dQp/g8l4
8HA/JltQ36S076X8Oa/MMKZeE8X2p3FrAdBfRCboAN1yPMwiT9lGLAxzjOHAPJ0IDQSVX0+BQvyM
sS3Tx+DRNzs2LcE4RmTrFrjz7U6/OLJ66z41I3CRLUGdQnnfGVqo8sLvAhgO1//sZOllu6OMXufI
OQSfSnwY5b61GFEE9kpUzLqf6+AaKS2DsqOsOsOsCfz+EiYesN6lcNKvd9boD6wajbQTc65z6x5t
aQRxKQ2pCGNwbpIgq5ewcFcGebjy/0ClMWGYQXsm4KMfc0Ayqv6ZbvoJCp06BJfyWLK2mTh8DNHB
Wn09ADOu9JN4udCKPXBgU45BuIMBLQhJ7x1q9naznnufZvY2xEKkUiaPNwe+Z6hRupE2eA24J3A1
KoSjGzQGBkRGWolKjUjxPQXmdALW6WEXbEhxLxS2c6+ZObsMyhoU6lzjc67CbEyD3i9uxeDlrlFg
CRrF6P7LBfkRKUDiP4RlflxWO5Z1zNpjd71i27GyiClLo9pFtKKBZ7avEVtFtoM5Yktru+sU0Rxx
N/ngST9QLpIrIMfE2WvgcAUNPrEtbqh+eu4scsnJisvxwN1dfIfEwMsHSWjMOrEHmJIVqMsT8xn5
puVL1DV0cIV0Ro2iamtudKWUMkrWito0ncMJRNWhoK5Ba9Q/P2v1O6hdZ822Es450zvxGkVt2pSu
86iDawUJdOxUX32GfN6H5iti7Zj1RKAwdlG6tRGvlmd5t1cNa8lDLwG8zCA8f46EWFwcmZtSsKaL
fz04s9TLBBddUXJG1D0qXs95jkgTuJGgINoLu6VZtgKv3L3fJOZqZ3quoZFRth/rrLZ6GINaZZjO
FPzqx0/uW9kGSM4a+36bnd53z7k+t+DNitC8i7ijZH8Z12nzqKWLCwDPR08cwVJVSKuZKmraQMMK
c7DuOv0tq8dDXMBpULIJBvcg09EaKgroL/jeWgedlINwVAPWHBP38TTqrq3GzBRj2petbmGyXoUP
SGpi4+uuZg5EawQlsmDJjlMOviAm1BfrohzTzQV91JCE7fVS1dJ4r11BYvLz4m9NF1wjbaTaM+yr
J+vC1KjD12EkYVhIROxmFwPtspvPHHgkBRBENGQKHv3BESi4sRaGfWI00xIJ6tgO6epTrs40APbe
ESGN0bV2JECPu8lqmi9nh65gRcJ5iZg0MaYT6uo18+BX/0k9+sxiAcTS/kMrc6weEdCG7oT5hBH+
Sc74ArROwlvONLxk7hmdgsAwVxDUowDPhH9hVIIy+0JIaQLI38OT6fvemUQd4rc4P4mPITYAEzq+
MDfhYwg7neso1VhEFmxxwqiwIQXraWVcicQUnCntKt1A1MPmXzLMfqd+sUOk7Ejl6w8r7xqnwwfD
XArtiOjBrcmthBvy9kI47888E+pTEmXB32NXwk+/uUgEZzMB993eSyLJMU4eGSQzuuEEizDKEbXS
3W2gUeoN4I2BA3yBVM3rHoeteOhLHDxr0z9CHmfufHDyaEKX7WnQBzFx0Wd7RLY+EgxF7W8B9E3N
Hdk8IHcxxEd7bSz1tc8N38GDhialiXvlJEmeHm40jG/Zfu8t6XVzukOEZelnme8vEdeZ6st2BG8q
J5OYj5k5o4UzqOLVKn6gEjJ4vr9WZRXlBM7na8gVFxkwjUhkvho3pAaP5wyCSDwlQ9WXaG333Uu+
tynenD2ON/luznOZxLgKW2+aOI8BKYNMULfO/KnDwYnOg2cJ6uhCFzspu52U0d32D94YEdhcjgOz
cBnTYgTWi5wFqXdzGqgPD65WY0G+UCITqMCgyH3jjTosom0izI4h/IHb2u79GuWPA7txsNKqdc3n
1EvJ5uFgHEu6MkjqthDoGu6YSiI2Qy5aXcMMbWVW/ECu4kks5kZcdLgoGBVjJPne6Kl4yxFBsqmg
TrWQwbwQM8ZBV2zzsVzbQBzXKTzXqIo0y2rvkSi4KbmYG8Qu38zTaN7fo9BnQl6d4ugW3Bla3qlx
PEnogfsMSdZINWSwRAI9SRZCRbaaPvKty6doPjfUTCG9VT+454667rda9mGhWzyOvbtfulxy8q1r
uIX1vrTR68P94gd1tAaFWMrZ/p/QoaX8oKVSOHq3LNHfN06rNmEwb9SlmXr5Kp1qsAEv8mShVgo8
E779xMCLEuoV/8KZxpJAlcDnOLb6YoVZJkqlBM+rngIvrBckYb2dN0J2dXE1nZTDPMaHb75xZPW+
q+opi/UKw0lMiKCioGJjIYDGUjnoGBEa4nYozjZyXUppl5Suep3bOTSf/rvi7s5PWHIQ+HmQTTMA
QLHqeR+j6BS8vKAn8UgUD8GgujnPqK7AZxIASzqNpxU6hYZHqGZQ+Ipj74+zQNDw35LUrnSaqw8J
8N5it+x1DXPySjWAesA/GKBT/qu7H4hDaosRFu0T1vBlGtO2bBla+hfu4ji1FM7fEvOBl8EtR6Ts
2REpYprkCy/K8FTG/RUuOCQYimAO20FhK7iiPpkwqV2ASGT+mN7gVc0xwj9UmAmRkWYpANOJw73e
h4L296UHyIyh4wmv70E4WiNH+J9DLsvUeMVxUpxBgAwlBEoW2hUqJC2WozXFnKhIpSm2WEhT8iSt
0yixugu/Z/S7keYZPn6SbA9R3tZIPKqyB8+C30qqiZvIEg/ITFlrjEPA3RoprEL4j6vVTLZFclx5
fMmzIlTxx2pZ/7ciVbIK3YDdk11RMwXnQ/1E4xkmAWDtU/YhJpllBBrL19QAzFPJUGMQPkBqvCQC
jrPJm0/3MtOhapXspFf2GFZDigF0FIXOPNq0LohaQGlG/xuci8tz3tb1YV9qDCpbXZK0kSLDS3we
Bfho11oCELLl9IWsPkUZ2iht1En9zTGHluAg31IDQrMqtc42V7DM4+PBG2KHKeVon3Y46bwOlaf1
wF3um35lH8Vp7n6iR0zUFOKHnCfa4vIaqcNCjvleJhY3MUuyv9VDhFgH0P8kHxSxtGyr/67IyO0H
LXCZ9BHWrVGxWgS/Z26e8XjALXOv/BLx9AgK3NXm+by+Cff3+GHZHADUelIDVJNibo7MYwmUWsR9
BcVHjhaP1poF813xbeDu/7vxoIMyBwJO96NK1mQCh8e4GHtks80lPtxYcJHUDUc4RyjWEEjxxje7
38lB1Pcrz9ZSNuG6pY0tb+AwxA6zxUGtDeONig9RqCq8/3Yc9h9ogyW9shrgI3wSENdG7+5xdTNf
e+0vxbZdH7hHK3nky+X+XtwCgWxMHYedWpRuxUt+cjLsdGt9mERtVVYFZewjH8Hl8wJQu7nQ3yWw
kmW/IzmrL3QfefpjQkQ9yjf2PF3PMmLNKyBS2j6AqPHowvpFiaK03DY24LFa7aG4QOGY9K3b1nP8
7dlpsvZfLaIsufN53cZ2Y3t9Xq3yERqBUK1X1Q/mrya+IrpfFmisCrKLZ6QECwv2wTnSkw5abBzA
ZHxvpP+Qvw45w5BymyB7hEyALxOJbKmDgWMG9m2AKoXKIJ37XAXdX1WtZF5s3bQEVhXEbsNCPoK8
3SbcF2CUc7YFSeE6Eja5cCNp5nHjBpr4ls6Z/eETHyaHjt4RAgiEkYghgR13evakTwvqXKXPrtoT
a+KxgR+ArBfI9b0O1CCEQQQ+eXN9U5S4a6TxXJvFkNcW7pR6Elw8JjiAdhGN+WvH1uSEMttxQBYf
3Tye/gV9SJT7zW1JIzdbRGZvEjDJPoPA2gVkfP7wyYjYEZwYQiNxE+xgzE1XU7jI6pTB0T+LEn7f
7kgijk5nXOoB6K+3MxnaU4CNCW5I1urHuyhL9BmngP29AFiYxRfMkDfVdi6yjYiQ75hCo8DtuCgq
qjcZlX3F8DfaaH/lR1C01JajXHRf1acIolu82OwmRUNm3draPJYq7LcnKY9vCVTfk4xQn/z8dkNV
xIWWOYxRF4EOnszaITRf2hCV5wUwyCsTJqT7ODvho0gbTCUiNV4/awfhmclooFD9CGbc4FHVX7nz
D4NPYqBoyOiF3dZspG5aBMzMbQjJ1cppHwXDKw9PiI4JB9V/spDVzz8uoaFPyqREsu3bCQpxRPiP
GD7SPHXivGX9XyRBSw2lGvIlMJ59AcqIkQbGMA4rJ5PPbluIe+AbciwW6ahd+aYIUoBM9jTg6TlE
TyBcAVWVGIRD1imXfutQ9lb7P1lP2C+HOh4p7eMqjALdnjfPdGA2rzMnTaSqGMdfrMZoLgk4TVfb
06DLHYjt+rNDtAk6ualn/F3dhvF6Rn6IXYEn0cmkIm8+sclQXICSHv7YnsmqxtzFpck2c3pYLgeG
gA3wHIyLLW3bCrHY8aKjNdb0JgpDyb0bWkLOPpuFbBERpXjGK7odg6DlV94D0ND6dFtQDwdmR7Qd
hERnBlUq+jKk1W+oC+kEjhOO5FItWARiij0rYDWY/Wt2gm8cdai1tXLf6p9Zk2/m+gIc7RnL83Im
NqfHTqb182Gd+afDhQoiMwcDlbjaDckkNPjytrkreeGzQIG9Ugx1XCHXd7ABX7Q/LHsD0QfBolVw
NH8yqAUdddI6SpQaE6fHxJqYUnvE+xSh05RKiDFZa4q1Sz/LQ6bwCSfFnZwzc5ECQ04gF7ophlPf
hJdaZSprCuUnogH/m2sOIrLXeh5/ndWI8+hpnBLuLq/bqZ0N4318RsZLumAd+FXX/Sn2WGOoq7SY
dfszSiJUyQD90n345zWuCOcDvZQy2NcEu1iLvbMPjSyGuNJrLas2zv1U4Vx1i/neRYmZMP/OwNe4
dtZFZrLc2qlxMIBUJMIpiGccFn09CvqLEZvaEs+U7hUZEz8aWMNWdY6Ym1wrMn32DDw8LI+I7Zyw
0G1qttz7yKLHsGV7i5a8KVaOu78Cu70hquWZRGkAlOXMJJkpBwHE2Tsi/dPDTTAC8Y5f4cIMXT44
DwR4lk1X8/UH+wbneAkFYbjKApKbPPFOjmmbPnG2WZXY1zIDlxwUOHu83GAFluKWLUS83pj7//9j
inRElFbaKLo72gleYYf+0JJn29D9H1eD+Ok728A7WFnp3F0i3f1XZK4zJG2kEWvT+QR6uToj+3Tu
GnnEO3ZPp7CdaVgYNhxLN2N+GpFzj24tS1E6pI5zR8esEy+pDxIKNSYFT0ls5mDHfaUt7O45559x
kZijR1qGRnde5snZs6hdC+3wACV0PdrqupRvbVm/ulCXfRMUXg4EFzz17TAIfssSYDA8sgYmaH96
omw/0wmjoS75lEnzSTrYTelAt4YYovaFv/9oHbcFdnnB+EKUggY2yVdScjb5rgR7SVEFMGQqPl5a
2lhxonVAC48B231i7RABex44aDpDiLb6bmOezLAY2vdNLlWpbKXbZsEyx20ZaKiSozch5FItE5zJ
9iK0I9oTpPnWTGWC5G/hE/fRGscILJ7M1/L5FiO5315r+zsT/fFWKfZOFjXM106tH4ag4QWlrY02
SADhr76e5p1LoxenPruomZ3UzhviB9KlhZOOByl9tfHFW+LVOImt+zwDiJpciMIcgaTLPUpQ6u+c
dqw+oqbrqcRbqSxvYWFKbUkT40bOkM6cxN+hT15mqd8RijASTtVj5qXbBmxGaAa0R7zIgFV9Ek5T
IQ4QBdYKYQo9pwqGMy86rd64Rmgm949XomLWijfysly4y/v3KYfbyFcbVl7o6ge83DDeWkJ2NDrD
01RDGRymWWIL1aJ7U8KwukGhXD5bET0YVUYlHEuhxFizmf/WcjxaaevpP2gAixqgcHosyPulvSDN
IcsoEbAmqutYtwXSENsyqMjFJ4ZfozqQOTidcHaP94uzYlANa6VzxFHcrDz8ydKQOLIoKaEMT0Gc
PrV+EVcLscypHQW1dd9mQY7+t6T4zfSiAI5Yp1rS0qfhAZtsotZF4daGdQaxOIoAJEEp6D4TwGvp
FKhirZJmFbQ8+wVhiqSyIM3/Wt/ZsLHv8o8E4L9YMiPKKDgsAmM6u42II8KS9DEOQVw9s3sepXfD
JMmfb4IsnQ9psm61583XZ5A1DDQB6limdl5PbzST0iKLO2+k1vYnUi2EEW3xsjPqiAgNfKrO5af+
uFBQy96EFKO1jf+bfCtvbiomGPuh3cqK1b8GKnVJtXZ2GebElTYgaUEPw/VkNlhLhljWCW2Habqk
6LZTX83qbs7E4G5u87U9gVG+v5/19tTqBQ2dAah32cwVX7Le1cQyvZ9QN/LGJWWjdqvYc4KuZh/f
I4svevptTSxcSBwQVy/RX4R+KbLx+TvH4fu2p154Muxe23LThbAfCPPBh3OoG2IMnY2tuE3NUmOZ
mFh5FiXfkemc7BqXYlnAGGLFj/iJ5fwbgcwgN0XNP9LBj/ogFBPpfKtJqEumEiuJxQUnHU4wrik9
9/QiqlUk+wQpxs2oN45g3cFrWKSPC0aF/wWqmR8LAKMxbvrToPEB4mAsjFcFIO+VQUdYeh65MgU9
ZqvWrXd9rzY0zb1W5szTn8+gPN57cS2NNrFmvz3ItDNqE/POFD/MDQQdLR8S1q8ixgZxQXOVq3Zx
boDnpb3C6mpTlv/sU/0Wv90TirDlu5n/lkpSTpMfT4eOy/lOaRtHDM5whX5RTPyOcOYWlrjXWcRy
IaHkj/++K3qmG1aZO7673sAV2U67pHRG+rrfxWpHmrkmfwoDBS+MBEXPolnri+Pr81vl+9hMnGEh
2MAYR3K2Fl3qG5HO7Ri5i8l/aGS1PomcTr6lLrs6T+DbQCS0h2x406yZMyyNmydHIpO6lCMmBmBE
oTZgphyDpq6RcijgafseH17GrMvUNw9nIgcRsPjPCY9qhi9VUOVMJiJ8jd7fUbY6xdys1mBwzN0S
RvHajzTfUhbJiH0HS3V54AX0GzaptzdciPWddgK/CBjLD4rQ+u1Ehjf8mKtnMVtgEVARRIzEpWN5
n0lzN1KrfGdvExJ7m0F5UhWQNjs27pXuDg1thOMTKY0NWN3UnxvhCfRRHivgCqQnBag/Ml+H4vrU
1g7WOL16c0FXzJyniYF/AOgVEwwq8eycW2OWREa8DShBQ/Y01BUR+piBc+isBkcRvwqW0uff7OwT
XADKwzu/e93uOpHpv/cZU1fAS2WtkCL+bTY2exx8wVwkOzgZR/1d3WXPIhQ/C8IR7GjeCREAvQTD
SCSbmzqJng+o0XG0X3wc/wK5bRXsdIdxoKum9Q+aSxgEqAaQsE0wnuEPRDuECkmaxjuEmO/gFxFY
0bLk78UNamgn8kEbTN3h+BNQMWeRqO3dwLZwrGq6f9PKE8+39BXsx2KGqOlNQP6+BLfzcO45fSZv
9mhn1XhudL2eaJ8xO+0uaK8fGVDJSeAMzYzLscqAwQtgX+/3h7JqGTu97Sba+WiMk/3pBqntpXNR
9zhWBrO8yHMh+jLVxPk4eQjoxeV+cQMoM86198zWSksgIDASBwho0Ga6pVvXipapt1E2XlXs4OjZ
+VKA6i0mQBFRNTn00QHDXNiShyubAE7c3bC0zZB09e3R/S9qm0XdaI1CyLjJtfhJuKuin3vWCyE+
fVW38ExDPqv6L/dA4pGXXMjDTtzkOGRHd5ggPAwifhyqfebd77zvo4ZU4skZBWOqs0Ls4XJiX+Fu
EbWifwAdt+uFQ54Q/g3gBpnPog19azQ+5URLEb3thak2AYsEpp4R6RsAqwR67tvWKZ+oRjvWm7MY
ii82xf3r2RjEDmgGdYZmfkNUCHpZl1142+c9wmxHw2K0tVqC5rC+ag+tNKGUy8mV5f2AlWhIKvo9
Gg/uf9suIUs9jPaTH0ZPzqu5AX/Hu/N4fH9Fvcy/sn83ZwI6B+kfKUl3LoQu/NYdF9q6DV5KjXDy
oxi2hiFW8UL9CPxbmgl+eHl/bONgqf6ehfEhJwgIT857z63TbYmmSczmvOxpjcFoVkhMhod+t6Wy
tx1mkgFAXCYuc4flcIbkJCSOfxSPC0dAblVQ942jS7ri0NusqSju729V02agisXbjXkCTb7qMn25
0oOuRa9Lk3ZUGbKmIbtXF1V8dYX3R4Xd32l6ZAL3ACemMT3YA+68vjJcYf+0f3lAb/vgUiF0P4Am
CBRBpNuoePeEPHzFGesIaivxNeDBN4sasmIZkpGFXm1sEdIi5vmjmIehnBvUVQTs+Tj5a2ZFY8yi
rQOOs1tQrkxCn88TFL+EAqVTQderE6Ye/IntigW5zo45cPLh2RYRxuCjMqnDBxawCFTpaPA0MMrM
DF/KmlBfQJvDyzPzWBG4YV6RtAZZYe4uY0vz0zVfrIPDuPtSYgu1Rp5mYudZFKbrMsM1re/jNWyI
INQjn8IgtoAnbGkyipBmfFPfOmDH6bc5FKENlg9bFY8Q+qgom5aaS5kNfw61D3AgyxZnmoWrlWah
e1+Yb8IWwwyWTJ8YdwQO3M6S6MP9RN2Nqf9d+h+xlxcWUi0fWaOzwYr8K1+nckVlkg5IcGXBM1pZ
4Ao6ho7I4YRib8iOXVl8/NSb+2wJg16AeoQAx4kCvyafrzJusm6E1EMWNdyOh1ZoiIL79H4NONA9
GJLDgz8Q/kc4t1Z48lg7d4h3CVB8hgYbRghLLe/tGRLzPi9UzLwrWSt5Di1z3RZCAYKMUwWLCzGD
FL72j/xh/kSEpPetEg5ItXiMcXFYeh8M0thsXAHlWDMERZncuTSslebzKMhoCudWL7aA4wfI5byV
0jX+9rvie8F8phsu+3ge+rNRp78tGSlN04taEpEu+2BT6l18RP0NipPF10R1FBXQm643dIuNlOjl
wvXSj6WO3EY4H9PvdbVCDMAP7Ly62pEUrrdmoYaKi8F9r6ZkbGTR4cg9D2Z6U7oSS5HF5k3WCKGp
KuQ7hk1YHOit2Z/cRFYCeaqABX1FXlwrGf7DpXR2AJC4cdjVTWEHQhKTiZ5jDR/SQd3HCXtcXysQ
kQpEljOQcZUuQ4glDTp4boke8svNYanxd5SSftXwG/tZiR3AMb+TVyBZWfXEA6QDDQNcf/HHwEGy
3cypNIaAfFXVPfpk7cL+vh773TJHGM7VRhADIJaScVJZ7sf9XQ00BzucxAGswSGUS7YGoExMCHP9
7PAmY7gyH8JuEnyc2RoMCfiKAi+xSe/QQ8+Re3vA1UybBnJUlet8rYpHTQvW6KtqiHKjQpX5GdBn
mS3jN/LExwivAq/3UYTO+RuW3KNMj74VewLkqI78ppbO3Cb18EHz+q1PY8c7YAS4ctA8UQpgUNph
49aGNGSnN5EBQNz6AA7cxI1xVxsUuFYNZV05v3Sjht9sU1Y79e7YhUnz8qT2qahYvENvSXHdbDWS
bvDNMKJFMOk453RzzIcdyFXHmjnsL3h4gtoj+R29/G2P2KqJvjq2NKbixTSNlSDkZElgJq4M7bcg
vnkh8dDIeKGbw3OtQhnC4R0zHlLiBIDqfrP7HkmK/afvWdxeBBJZHn5DlAOv3qhClmNyM3GxFsU8
fooi80aotUUixPt/SnSMmvsGSYNhnzLyWnhoimura/pHT00KAzkDxvVazd46d7Wi4MOwOyzBfgJP
xRde0QoVB+qwW1moST+k9Qi6DtpfdiPeqXDw1aatH+fMY9E1H1N+PwL2R+7fHLQYBYKtXIYlYHvR
fFHoGN9pukjJ0DvZGGwtlSDSPbPiriPXcpvryvQDGdFzNQZX5zM1vl5CBScGcnKbTLNgVyU4LoVP
CyhFLU12h/HggiWRG+Mv28YF6RTIVOtXoyh9P6wXniC4pPeJIhqJ6WIIFTkEb6agPNpOmUvGOmU3
ZfDxycYsVmDpmF0hJVGUOapjHgxOZsXbrWH97MWIqWwrC0Xq60qFtLKjSdH7pdOhjQSRo+dlcPiP
pLvb0cLshYVwp6/H4ns584coFd4n132rrhemwwsVcjKmUQooTvK8qsasMcXFxbdLQNVF4FSSjMA3
IPpGf7A0DXfhjM5Cn1sr8hMUGnzYupz+okDtPw0bAN3GwMxUgUyq88I40jIG0gsAlryMOp3cUgQV
id6DqcuSqsJ/eLRYVJe0mZxMlnLB6LE8HAvCHc3Tn+E2PyEe+8rOn98KWwLpZMnZVUBmDvZRxWJI
25Bl3GvSwr7QeseMNm2HRuROcHWAV5SunA2n+xIH8ypsaq4xH8xGkNergLtdWpT9MDJ+JMUfys8h
EmSr6Jmv0Lp4HBAERHo/9EKM1aiuyNaI8idlNAQExYQEgMzaV5AWsPqKwHG24RAkGhnuXiT0hnhq
7NxjSwYAT1SGAHPKJ273yWuK3jmFMPCa1f7EYY+fYeO/Ku4dAfFMr3VAygUh5PoIZ9NH/6Zfe/Hq
iq4avvLVT2UNfbN/A5Q2BrK3WiEnQKGWCSQsiG8Zk6honRwJNPrIHBYxRFF780NA8PVB/Qk8+wg0
G4qU8GtYrTJPlK+Nrfkh9i+GIl/cyJ11sfzf08Qf/XU7j9qBWzkl3z5+fiKUUfNi2TYYEuVO843Y
OjY5f35Ha58+8NwAM4MgfqfR74k6Jjcw2R+YlOYLauTbYAD/CSJKaq62yc6PYvVPBEsJL4XJyG7S
4ZB1naF/FVJ8U66SnbLnv+rd54v9Guz++zIIctNY6wJC4/zf8uN1RA3rAw1FnT50k/bGgQFw9vLT
jeMMcaF4mU329ngxQOgChiBlNMaFgSwG3LFBIwCVbQ8IUYLUZ317awKXdUmX2GTGe+GyZQRqkr6V
5XL9gEvPc+tM9DwbLHJjEZjD5FnaDKciHfQaoVZJCMF/d/J0OWM76ozMvCwGIMohLq+CSoPHZN/g
TVYYGsyPMUoE6hq0XqFeYdeVnWOKf2JR70Fk90Y3gnrxak0GYXoAnkFe+/48DBjhdHVGz25348et
1AZyj3bKWRMLeW4tCY8U/H9wp8okwVKF60YNMgFFUJSpy3pinUuQAlebMVUltEfDPDlC5eapm47N
h84oCFOG2WOiz9x5q+5EIU3cPcpb4SD3Sq22/uNp39YUyjS9oRfelT6QC0yXBZjDtx5Li0oo5UXQ
dMPKmfsJeWiXRY3aaP4hDVnuyXsp5DGL27/tZLIOjQsGikq3wVUFF6MeSGBluvyMH0VyxgurJIaX
t2jW/iHRUZILRGJBeswnQQ+XSyik4cbpMYkOmUIOdLWtlBMRYyO1xoqunJoTXYdpONa6i+Rga12p
mfaPPL4vxUCQbRcb0I66MjtidUSevFu1/4LVDu0CTJpxgBS69xPjzXNyhVDUHl0mg2OqX+46xJIl
a7FyyRYQN+pyRohLTy5IaVjT3FOZ+VA5ku3nYob+zavMhkF3oPJQAbac+Lq1SnzXt49V5NMl1oFe
OOXkYXoRJqZfVn8uZ9zs/F5X/BSQxOqRCZR+RxByyLH12/Kw8D+FczQIR2zid4xEqTMD3/dUKoMJ
ULitFkI95wtscYOwDGM53MIACX/KH6uFSexLU4fTKzUIYVI6Wz2pADI1i7jeqTq7wdXy1OG73HX9
s1QaEcJsaGY/6E4g1mQWQEfQWguszqNeQE/WXUxFlg/6bpJKABckPZqLz5ZFhPLwBDcKwx8Mk7W3
gzMj4LD3jnKxVmfPmsX8HVMiS+iyCxCxgFl2HbdTvx0txO0gCbd8zzIa4H5dpe5T63P3g8irHtyF
pZDi+M1zGfLwLahTWgjSWv26t0FrFLujKrnIoN1A3Vpv9MbUL04FseVPLM5pGWMecP7v/1RmM0pq
jiGOiKsSdw2UFckp8mj/V5YedWTMWDAZPCWwOXcdQnHRJ2jTFpxI+zsO9y8mJHoENxH/GOmAOvNX
zRjsApAwGPAv3XqayE/KN1IwDGMSjEW5ynkKV1zmafYomt/LUCjIInM4o9z6c9CsfOydQpNDF909
xzx2eYYWlupaEtAdr6+HbmpuoW7imRyHl2fZwIP9kwATfHbXZ+bwdITtwL9CYyhSOouRI7kvm7zt
n/PdWiW8wZ3RwT6hRHTWdg2RiI6v7WsLvLJCFtOjLn5S0Eu74wlZ03LSvIwje0CHO5IrjE3Tb1qm
NCdFH7+zZ6lvK0VeHtmvyarPOwNVYwq6cDzevivKRBacHotQ0/06598JsnPphFwEfWh2p+MIYYVZ
UTuCnsO3j4hbRloN1OhKeHYjytKnGd/zxRu+oJUgUDdwgoAFI7hUtSL5hl0z3uBEALv085HDe6w2
o5VpuO9QkZYAr8zTpz5wnVqF4PsfxRYqkUkpL121/5L152FFi++bA+Hvd80Sf7iI11ofYOtQjXeZ
BMztliqFZx2M+1ie8fuzUIc53nJ5fU+kALMShUpW4FbpphLn3O7AyMTCRwyZE2sP99S1McfFz811
B37Dy9NxjyCBLVC0w4tryXU+EbJTi3riJ8CUsm0SeRSKLJXDYc+IiNdDmwyls3z86rG9UFtquOZb
WOQ6jSpNLkNqhLXk5fIlzX2HRLCBt61fyX83kj/27jl5dnM8o92JNaPMqVybXjbOR8LW5LLU6Nuz
wmcYsyipwfxpDuQewW7ytixNJrd9hhB+88TrffQcAF8S8pOFHeOyRMkZlQZVOFl2JubPVYQ+LHBJ
etNVTLLZbNk5FC/86xU0DSIKtpzpYMbj9uEc8J9zeKF2B8SqgZgrBQK+B2acTczbIghstP3x0cD+
X8kf7YTcc9x85VbDIdVzwdWp0LWsrZtuaU9XzlsCfT0nIj9azIk8vUmtiNRAqfNaV8aBRxsSsCo3
Hh73tKwlyIcGalIYQvmTvASYEVNvS6ZT4dHyYCRShkuLHVuD4tDK9QHDFVHi0Vl8qBnXequn0mDr
FgfElYS3ILsvUt0ZcT2CSQNKtgKPPfDWeR3tEw6z5mTl7OdrlCapCIDtO+WtPL78K+BdwNzrPs+r
kfYBXLwWHoJ1zN5UzQEvo7EggEVzWvgsEN3lE7QxmbAL2xFolCbziwMe5Ei3vBpYTIcVu1C18FoB
hVQk8lccDChJF++z3cOm935TXjApP82pPmqSQ4j+oggBkIEyViP6w+1snCUI8aHzx3lebgKoHWiI
qKU8AEGQS5Bp/Yzeo5wu1L0jCNxzgaZPanzpWpfxBgxxgmuliozNfsc3RCR3T5qCCmQOhmdG3NIo
K1P5daYe7oRQvrGERXsApVtQ2wXvOQqpJrKXAy5vtWFuhmvExYkYYxMvKr3OMLPsZvT9wLsucJVu
hux1VTRg9ocuYu034lWrWKndiJRzcHnnmB9n3u91i216Dx/roFzIDN74qcTmCAwpz3YVIzI+PUk2
7teJ2GVV+HrHX9TFG6vqckH3Ot8pXZ7pWrW6RXR9hjuNEid6cW+zyXRM++hISLHMnartO8W0SplQ
K4AoFZVVgFSLUKJIoICH+hdWIvi5CxPmEyKTtz/04z1jWJGPv2HkZMuT+jCn5/aZJPe03fdMPxDS
vYUFO8oA72XRKRStOyO3pRPUtXpP+hFDCxAsYa6LjR1R/Qxf4eQZ0C4+t1iTR4Uaxujy85seWvXy
/N2pl/qZtbpKMpcb94hI3kpNZwa9SjNCxZhCjClDS8UpteXJtVDDLKd3MwGfSLgGSsOcwtCfJcJZ
mwcyRU/DqC69FkUPVNyEJ4rhTE+3aTFR8jTHRS2klSpC7BlqmoNdKmpHRBmmVMJbCfgO3wpV7m70
QjqkZdcF4iH7yJl6yvETt8CuggBULZxNpV+IjYUpq4Ns82FXn6RljgVz3+F+taF+LGV+iD0JmTnu
UW2ISFdkZDtHWwkBwwMggwFuK0FbO6Gzc7TiOO5a31EjI79hWzkhZOtPB09eMH2WSllWhRBjpe+6
X6nvsI5vxR5qB7ADd3V68awqMA5D32BJikpupLoHBKQQA+dLWYNgmmAqvhk5HAS/sXXd4tsltvM2
qiaSNTf0Kv7aWs8iYPeNDfOgWs37W4uCkC6GuYYXYkBOSRnFM/fwEYAGgoBoCj4CBinKz+u6/JMP
YVUNwmxNZGxEm4Cgan/5upw4Di/AF50f+mGLkr8LHTT6dlz9SB4qaajiceysC+6fsypXoOsE3b2B
iL/2hAH2ZmZq6Uaspazs5LpynOBfCFXuZHWdv94mXiq4vBACHteMEqi4BIgq7mZdNjGPgnErjguN
iOyZMbkwjbkR3iYLyf4AJEx5u2bhIBxNjSJLnUldOcsDFUsAR85dccJhZuKoOIT3hmEabsPf8nBs
02btdhJnWZbLzrj05+HsbhphHnAh2+Sm856htLqhGlrTGxXdG1eTk7iiydK3L5WwBk9hFvUdApd9
y1t89UoNKinhYJhW2NeckzBAoZtPJDqksocctKjV+/F5i0kgi841SX+DraoENOhYIlcWJhR7vFHy
WmW6mQzqKvIYF6GSKmabvRdjoiXVMHey0CA6EE5LtEqgevewlbfOc9DBlpnfuL4QjOjr57bhHXSj
2ooZy7+87Mz59zprm5DELeo2bagczck7m45zph7bDhqrT2fCzyWPNcnoXMTaP3thp0GWJjjhRvuy
5oAR8bW+L0hzXYevRkKKKFbceHZd/hg9F5ho6a3hFGjGhZ7ePeta7DfcY5Dcevv7GrJHWFAlk87i
sI7M3O1bY6yaB7eoFf0W6ngI2IxkIC2JStKnr+OJIIHln2vHXLzel8DGtv9NbcF0bxXsat+uxuE0
uKvPppzWTW5PdYPybpXWJwXBvB6NwhphpFqah25Np99BvDoBPYQZmC15+6/4CYq0wUVhWeyQlvH/
Fu0wont2Ik4uuofvNe86+iIsbrUp7gxbtLK9OQWlKkJ1iTaTuQRAWScC1VzHry7zxfZaoSnNNsLV
cbPKmJd8GDRpb6YFg6hVeGYqwAn4BCXrkmtHnbOsUCMdR8+CyrJMxvztI8idPaz943kcy2CUtCbw
x5Mg2LG27t4Dgi4rF2gfuWAS2wwJWKS6sv37h4lkDvIJNJ0fvIXYMnPhAKHS+yB5syEc9qnaa47l
xqJgGrO5B6+0CiSHH+zhn//RtYnMhdCcL8pPAOx2b3iitthOzUr4ErBWLx0Q0QNIIYLR5i4MhCjE
mKMh8R00TsGPCI5JpOxCANlN4Ax4lOeH7tNgs0OOD4ZJqeRIQo3w3gWecqPpSCKzPpuHy235h+bT
O+fkeoPvJJ1CbOQ+IBhNcw3/zYPILCJiCefSuRgsvrERi82ZcxiAA9y/ACX4bm0googqOT9bYzOi
FkqTj3qxvRjtVln//F4lTcdgAO8o6MUAFCLtQTC02FMv8oNNkAcVHOFj01Y2T1eHJwatT6L4tWP0
U6aJ7oNdwrpG0sEmBtj3kehNIIsdMGKWTd//fU4hs3kvOjx6u1QVWVNRz/BOtMJxhXLFp1b0/zow
ID40lTrpb6SLEgGojOVgafZejR+B8WWul+KPzwZbqkMCAhV/1ByU4+MXgMkc4xIzdMERJtIXwqU8
IWRGKOfN6h0xLUKlUVP+FaCy6ZLMdzoB+TDf73uKVdPJacpE2CWom6bcm67O23qIUY+53F8BjKGc
pizfcywavuC4IwcQ9nKYV9SgXNUECpDALrK4P0Op2PHdCdyDbXYSzqmHHCrPrvcs3ByapiNh7a1C
/evElA+1QeV1BmlizNRkf79VruKUZNtuCvblGMUM01dbxwTXYTb97nIiRln3FwcSO9ZAdBRGXAqA
vJBYdYmtZwUke9i6ulksxkH+0N+h4GEIr1wkh1+af++7IGlG2QeEFi8GefD/izprbRi2BJizv8fq
aAqs2xib6VHGa1NKRSC38vJJRYuooeBYLSMXV+AFnKDj5v/bV1nZx/AREU3Zbz0feMs9mk1GEjJq
0LM5Up8OmCgwN/hl2IJh5d3YBCq/kwiQa81WuX/q5nFE/W2Ia+NbsRy/Tu78Ex0cpS0jarTK40MO
3SHkdwFucgsaDHXUrDIC2Uzrhqde7fuD+B/vmOoJzOrIVOjpQ/jBHC+hmhI709S2TCdK6M2oWWrV
NPgZcPRFLHLLkTEs5D8rpyuwmfuDWoUsDewrZ8hLyKfuIWD9oV+uFn5oW37H+IJOzFOB33YPpo8T
Ddk9iqe2FFFTz6A18CrwJxK81AY5wmKvudpLyLakmvzC0PxYGRs93jr2c3gnyLVo018rw62uPJdp
hh+0I32WsZZXr8iIxrFReDvq3jcSQdr53SJXBEnYrXT+CyXD77ifO7EWVbpHFLpPNxzwsnguiF9m
M9lkbP30b56pMjB9LkN5R8nq8ObszWUTxZX0/y+mUGv1V3jqsfU1JK9yWUNFts+mWRl44KKk3vYx
Ieah0UYQmCp4fr0iKO4DFcXwWYrb8UjdN9ZCnJum8cS/nSyeyugHaexfXHx8ymNQj/xlKlEOBIOq
MTqXd00hz3A7n74UvjaIr2fzp3/7JoYd0Mq41Jo6GvBCuG7IVFnwzZHxFU3CMqMDd7dmOBDXM9WE
KJuyIvwy59IqU3tA2w8Kf+NFkZ+G/YmpuxmKoH2ewJXGHww0hEbvPeOjDbVr03+JVOaGf45D9q+y
HkrvrHJF1ztz6h7oIZ1QpD0uA3rKN+sp1Go+xlQ1pa1Xxtgv3Ye58KgMRtrIpfQaHAauFW0aZyhX
cD/MZA5nSeQetcgjzIKHKDGxhO4Oggp8hpD/4uLQ5LY75DLlmx8vOAOyOCtsWv6nCf9YU7B8P93L
Lg6zSg5jmSOsveIF1e/HZreB586Rl/8dvd4MC6GaZpkmau8WzY0BecuO1RdN8GaylneLEfLErAVB
I0gfc0PcS2+NAK6NVucPORg0vI4uPv4HlYsQBsk70sXRI0R2YGXtKUKl5bYGdZAO2XB2zQRMxFXr
DTrmWOXqp0e2hZkwkp/KuG00Q6lGUqWzhkIGbR7TDqJ1DxS4EQQxnzk7MwxKFqgAgCH0thFzxplv
t8LtrXSqeWiH7se+vxJqD4R2WURxhbAU7OHBgLKggXL0cMjsaVe38Ptdc2YGcpFy3vCzbZrqOQmc
lDb3eC84RK1HZ26aya4LEnErysvcPVSwpDA74BXjUT/r8c+DNvTJ6IfnfNaEi7R6OuYJBny0+793
0EJ8QysCd4Wx+BH2Cxad/CfYHyKe79Zg/33gvZ7o9/PTJ8+JS2QsgAB1ZfeuC5HPNz3DauseH/0o
vOA4tkh3jcdkJey5Vd9RM9ScnMlhTraRvzc82IzGENQ+XmeVAdXEPOJ88ZAUvcSnU17kQk6WAgRo
cvstY7CrJFc9mBk2fKr2X9/G97UUZ7bwKGgTGiRU47c97jH/b6FnCiwu8pp1TIQMeEc87oM1chf/
uhJWCwsTDdsYmMWEkpSeHDdiwcDI84jbmeX+iVIW/8WdeaRk8j2l3wKL0Var9jH08H2XWy5sIVlf
cz9R9eN9HFlWsTN+SqfZ6ekMk0prZNhGRZEbgPlUpjJu1GJ4vV6V9GRzNmLQlqsiRxNwICHQvC6s
JwJmGloEjQprA1sLNa6KIOq0XUXtK5Mpe95cG8hRhGHchpvtdumJSzmYZVJeTgFkv0IZHwRO1Bgx
jEzVtp0LWlQ1ODnI9YQlw3TPJiXxD5l30N72LJuLMdWjwAQXsqTccj2WfOuukd8juGOorEKy9eF8
OMbafD9Ioh2rLylWcpt+HwP1grbv1iR98copKHMHIsifStcTfreQz4QOJ/i12eilJj6S8JOBeGzx
bv7KNKVWze52d22hgiBYtLoJQMLRe7FN8xvtRdeUHCjkljLfGtG+lRynd8caqN++uXNbGpXpoOAV
E7O72BIgaXMC6vjo4rpYkBhsJ9LSpnUe7TUpoTlR4j4hDDJ8J8Am60mBruIAZzJy7xI1YpxdqOGi
kRQXFACHatNls7khCVNAUsFkIQY65AVIPLv+4/jsZhtR3GKuZRA5m8XadJj7lTyMQmF5KWU7SO1D
29GysEN9/ZU/GV8V/2+XwMk3Sf5HAAMi8jcXbSuTEcQ7ioAGhnlrCn5aoeLpgJapLiv7N+LrSVQ0
glQTeCtp0gY3K1APrg/j6LYxhRbUdUr0ImoBEo0zZu90tAPlbjdubMmAMDhbbXo4zokjwxH2A+4z
QBHf1GxpcscSltubQ8w4jFs5ib8ybu1T75HC+2drBHaxsljQPKk64P+wTYbxk6vj/Adsku3cK3xC
3o/tc6h0jbCC+xy1mUJwOQk0GLCkPW0qSs9hpu1oKRqTDSrzeHcMRl4LjGg9I6BueDi7EK3ititB
H8jWQ3NdYX14wmUxbPKhok1Hflcw7VqshIlX2URWiPWpW5VFyy+TiCQCu5DxUPCIwDV46Wn5y8nx
Ynv7smi0zg+1vLcXfp30oTgB7DajBUKoce6kd+xu5isI6J1EtUHyclhgeGbpSRcxkRuG1i+r9uY8
juTZc+P/fq5caLCEIQGWby2ImVBishH7xnfUxWyiN4iOkUnaEIIUJiCEbrDsKvsJUWZgoZnzHbfu
szHba2HGEJc+xMuA4QZuJNNAJvsMEoCW8vwA0OLVSpzn8HlIE+qR0/ETTy3cY1kCUzM5ZDObWaF+
kDUzQ8kVayGmtrCjTfGkcjEs83Ak7OfmP5vyeB7PzdlqMQHgRdBXhAqDw2OLGvhhDS1SrATbC0hY
9T196GX+asRO3X69EIfr83PbkLRZqMy070kUh8QId4Kw7Os2zHsNlXJy0ZE1b+WD/Et38j4pTps2
N2D/hT+MZ/1aoTimnr6cAsBktNbQMXRhsmhZGYGelyj7unFeBn165O4HPnMHXmT0tsD4l+dXUWU9
K37aXqbJFe3iC3HSqlgtFWCzZAcmr+XFQ36iQRjLcJ6ls3goC9JBdqItq15+juK6qdM2a125lCd7
b7FQ5T2tXmOiX3PZJ3+n5d/uKqVReXI3uDId/voECrOMaF2tTJjmUS6xMRkxezCR+XIXDkrVCCh6
TOGd3mLSY6bg/sIb8tbenD7oMlm3P+CCZRbgbR2ItFxbbOvXIBFPm+sDFYoG3IwJMt81inZfRxE9
nYrDO7qB++USrC1uxdYtq5ATg3C2axDH/UK2sGDOnWleYP+uOnbRhBhZIvz+5CoS43j3/CbPfCN6
2OXmmNIELqSfhaCkpc90dDi72ujyH+xSQdVr/+CHXv07hSa32yaDjQ8TjwrJqKIc1RYSUyT0E0hG
Flz5Y8e6tNTp8BSX8xglVpYmT2xrk4t+rbb52BayGuBQcnA462NJDv3OtTVluFevkqzJ3h6K+YSX
pgCRy48TE76i7YHUX27/H/WXUpAZmZqS4S7cBFzMqnEi8+ZpwRvIuoJ7x6QMaA26psJaJzKFYRwK
1R06aj8Fh9mGb65zfHnsPEcsF43A8AlOdpV+slnfoTJCGPLlIims6Irht+DwjbN3jp90Yzk6mY32
Sppu7ddm/LWnnTjrrzsjTUIOHbLS6oSJEUoob76xy0cdi4Tgb0qUobnslUEKM77QNLTwHhAp55tY
F9rTHoCP+7l8elZyMiSEkXpTwK4f0UGItystpIFAZ2+kiuFUyjpyU2/1mowfwnvGxt1+XBDrGjjw
VY6tFJ2YFPBGzxWYTOGA2L4V44FLVUH0Gies5NJ5kdsEon/wz+3sM0Ongk9fZJ7cXBMWDliH9pw7
ewhw+qczdb6aA4SnfXyWcW8pWdzK4GlYSeumswRYj+sgCaB1RSF1I9691yKkVFXGKsOb8kJnsO1h
BeSXSpc8OKKj1wjmvbanc0tCQY+mBWKGHhZuyeKQJQv8f25p44WVPv+puIllHBmGnyjVSlsM842s
FsBmVzGE45puXMLsJhUlbJxw1353bBiI3eykcpTowTJGBRkHBV28a6ZfJFqlGJfLiq7H5AaYzE2o
ePDAGTHZkKdi884hiXgkhbQ+5ngt/wGenpg89nNBm/pkcAlvRqczyEHG8ruT2ol9FgoOrHyJFylZ
uCv8DTikmoB0g1+lNkPztV928PP32HrSlMNEtpONBLrmHXFf4EjOhYQBFaf/MaM0E6hQ+r+Jln7s
GyDfVgsY2hNU2k7rl3rRaPVQco5vJ+22K04jahKjQALZqIOzCedffGhkzVGtvQb11wpW7F7W4HLW
IYwAVyRmh9pT5d/gxPhjntUI+KQiTmm78dYUaYvZwYV3DU/sQ6wxx9u07PoNfVOb3WjCHHbxqqp8
EnIY8z40BtgkbjgTDJujmzBUPmQorWbPXbyMrT466XRRSJ2DxrIUro7USU6UJQ23cbCMWmxfwqtx
j3G2lPZK6Ox0lFHyVk7PEGfRyjq5Ra2YOC8o1kXaapNYb2TqItjdrU/KBJZehkodwdtEajvWMfZD
i1zPYCkuetblHMSxrf2P3FCe/RJiXhj+I9sYCzNLRAn2fVNPobpuYdTsLrbUse9ppFZJz14KEoZv
FRzBeuIJOpbwBcBNW4KgvsOnpH+DW/aWWYa83YKljUVT+Xjzdi9HKrc7U9WtfYffdqvIrI/sPUym
JP4//cOYFxEFR0Tv7thlRRhcSDTOioqWdGlt0bKV76oQFP3wbvqs3EYCjFvdqpUZv032wePhGarx
UZtvl9OgWiWP1GOXJNI0SHT1cNmbNsIBaw3U0SyCkay91S3xuprxrYl7I/9EgXgBYkBE7Aobu1el
Tfm0/hiE6xdOmkUvqe7Z2hJDa9H1zbOHFKw8I8t9kiKJvpY7g1PhC3E9eEr4cQclfFx8GhH0sFRm
814Pj0/Qo7NI+g/okoNpDxF1QydyYIVxhgGvGrA+TC7xJ39dAeUWc/KwJwxX9Zq5DbeBv17Tl2E7
5nnq9y9rt2oJRfZRSRn2rViYV/TYnW7/qjPlopMu7vzqhgQthWbWYnoNmwApXD9vicdu6RqyNNz+
TJMiUZ/mq/k96Ve4gh5zKNuy+rdggRNMUURCJLMVEgA79YrLjCmtcARU2rutQCjzftB4gDAge8i+
irGv0XW9T8mgpH7HJ2u7DpaZVGKxazgoTO62H5Dv9WixcE+btfCI0+XhketqxBObXXosFWp5aqJS
uHWf1NqZmO5Kgdb7qaFxu2vrHsLCczChCsQnnDxxmvmqcxVdIr+4HGl+5VBHPD4fM2YLp1pKL8RU
L2cGol+06dNhfMyuPTr7ABG0d4T/6Hkv2FNB54IX1fn+DPxq5rOACfi86weTY4wHkgFA5AFsmCRA
/Mfo7Gk8rmUfFAbZoQC8wPPpwiFdlrJGrQ+A51NCk1jUdM/b2MxNAEXfNfy2/21hi7rrJtMLAoy/
swTu98snKgVR1pFPJL2lBhlGo3Tcs1h9lZXSDYK5ktjLiwldX+23lRwtnNC9KGDtWzDhdFpqyIaV
iNfFFle30NnKsnjATSA64Mn0f92PKpcafHLBeMWDIOtj3cXtgIGfLDC0+3pKv03ajhAiTO6hDSz4
QQxd/d37vgk0BB0fZAhf9Cu2zLYv41LxXetiDzWfnuwJdA6lQhLHJ4LvbcU1yB63mF5uOzLgrhIi
ZsWIj4toahNnzxHhq7fhx8S81ifjoxfaIrx0XmwePD4UjUd4mZwTdpY2n5XOZifD1z2OoG39d9pg
qtN5VhxCHGOlWhLGxhMiYUidPtkTBBBrPBUVr+3n1o9U2rx3BSD200HhVeJXvFc1vmNLX8kaplvy
FiAIoCIJvaVF+x/wMSHRMgaw2hVWtT9nkqL3hDRNapdCPmo5XG4RJeRfH5BIFBvS3p8U3Jp1U2P7
NVVxEb5TQM304JdS+wLXLPC/aKKQuyE0RbajNKvZzPNBMsNJCsQc1mI7TzjTukqpjpG7Z3HjWLN8
k5wuXWF+kmkudHTCYk+jXJprFvZcZ+Ner2cXv7nEHl3itXj2cW7lMMlsXwdDIrZuvXOdjdw4tPFm
q/lR4t1wFR6XIR7dNwDlccOnpEg2b1JKDV0Qv2n7QUUgbtNi9jiveBdzNvMBIXF9pC8Tb86+wKCc
9WBk7MkRFVd6d0+2a049CfmlAkd3fGIneANBVP2urVHWPaxwuBTZBFVo2szdZgdFeiXQ19Uk8VFH
2coES5MNeVF9fDQPzDeHeFD4grM4AF7rN+IRZh1ihah3MGXpN5V+kdOgNPN+R3T23JUfbVB1zoRN
CQ+IPkld02NXeTUI5xGAX9namhFi/ncSd7HInbqT8gZSvXGbPTmUsQELaPibAHeSZu1XwPomFyqI
1UwAgt7tgokKGUIv1yTxayy1ldiuPeq2Xr7acAi87mUV3RqOUWd+Wxs4QXmbxK9iBBZ4zNgZ7GBz
XRL/Z8wLAlUHZqnW8fwvyx2kNcpWDLmMrJK3qr2O6eB3z/sBgoP0nrPzRMQV1NKIFSilbW3gns4g
AdeajAbBqw4UOFC4eusk+l0dLzl1o+85H9ptjW8QcohQhWRQl9ux14WFqnPEzj48UdrtnPJai6ux
rR6nF7J7j2jzfXoAaByEUSe6z6UWiiooU5gcoldyhUC8JzQyWsGsM/Y9qSylCtbUE1ynSVtazl2X
BO15mJnIoLZR47mFYVtzPs4AqsL/n+uWulXRBrXXAWjtMrMK7mNtg3Dm/lqmiYd93L7H4tqd2oAr
BIwI6xvvfnZVwajFth7RJPx9sBN30AjlFy8DtXUBX4k5iuiA2YKHDhDuAvNZxP6yBSMLowKP/51a
klTOgrOsC9LQmD0cU/UZbZeCb7YRknfDSYEPCvcYdteRuXSpb8VKkMVX8mdlcOlH8+pr+gVmX173
avABhm4Xm6Kp1RQP949nRGBndqINjBF1SdZBETVs91TlDRQpuggWcR+4ElKChIO7GZQ5RkFhBrUW
rstD77LHLevgSAIXlHi5JL37ze896IACuf7WZYI/ZvSHK/2kKTwl/yuV4+XK8Mh2JEnE9c1XbFt7
Xl70ORyeu6KN+35aiFsO2q5URauZK5Gv1dw2+HxoftZHVvFpdMAPBgAPZoB9lt+dO1NUPQ7l1i7T
EZ+xfu0nOagOULk40FmbdM1aTUqmBo71xEOMngSFHdg48r5hxsOs2EE3gsEXVenk0y0rpBtuq36l
4hvmFrlAR+ihLamo7zgCLO3INNOEJ/3WjZm3h6jATrLAah5Fdk894kbNC6IfxmbWF1rUkRvlgoGr
iYYYwK/6yk7UXtfQOLabX0Y7h9Za4IFYGR+qMdB8CZzkmLzdqTvXc2ph/b7kNbS6p1422qnRDWV+
N4o4DUj1vI6OhGz2Q8FmaaClZZU5y/36MIzkDimKaqU6ikWFQkapBLtJ1SSJkJLulLVvWXb7291f
16bd0QaPstYkDuvaZNleQhO3YGKUfLCKFlc/Zb1BO0q4Cw48cmxnKH4bweWsAg0u8zLoXWRZ3pID
gTAyhFzx/zQXbyyFMMVUwy3qzVMhsYXUR4Z02dU1Sai6a4rkUzrRrQHtkXNGdh01WsF88X8VH+ys
geQ6+h/BXpu1HQCVbLmn74b4EF0LM8+QTGLiQYDk2M+1PB767zoceod1Tfn67Czt42Ksgi1Cl2U9
VnCfqqODYjwxdoxc8wkInZfUnQmvfj+Rf3z8a3CruvV1ksw7GgL8w3NQvdf1zW7jl0l/45XvC28L
hXoVs5NTrFpDJjhBLzO2AbwonvpxtgBc82+gn8CLZxCmcqY8nj27q0l2Fxl2nbGujXEFp5z2QODx
w3EVF1xZcCC6yO3JyTdCR0NqLXsw2br3QI6E8Y72Xlib+AK0VFx8Y54i8XGik0sIfm8V/9Gnonoz
fF7vF00bGDycQUTqioetJY7wJMVswCEbOkKca0/y7rRpSme6dED7zr0IRaQ5/sak1u10HqbcVEJb
TB3GUqUJzosrnuz9su5NUs+0RqQgdnksGPJGRSgPtu5sxXgkvg5X5IuraxCQ50jqF3qeTe4u+2Hx
yKbROf6WlxG+eo8olR/Gz0CWqXXuZ9gciMC/5bMFyUBXLow3pUo8eN8S4G0TH9PVUkJrc57VvP6c
+7+3XBgv7b76qNw8Mhfknj0tUkP0CZsmSYMz2+mt2KVfTDdnDsDHXCYe+Feri7tUxXXbc8C1Slq3
ndpW/CnwVIlZaa+AFLmLhLsilCK/C9pFbnZg1SLyvlMs5c/CkfzRChsYPQGC6UaR8slygLbMJ3Uw
Vj3eVKQBauvvAW7MC9/r6pjDlzOke3/K/ArbPoYf2cW3BVEYxhx5fjhB2wKZGPQE6kIwEF3JEEmS
koEj6FkQU5AvdPjczCvuelcl9CdDOTmEL1LASCkz6ZrqajgYtwcBXeu+Qv1LkfYKgpcdzMeUeqUD
3pv2YnASPTIXON6o0hdlYCuI53CLepmJtmIvQ8BD1qdk9uCILK1lfVRwmu5fEdHWLxrTX5TF7mRl
ZKAwi9AaV0DX6cpN/fJdLACR2kJhfrfWci+0TPWNdomDj6W9TcGW7ypxfsUv8jGaBuUsuVLgo4A6
2DXfR23emRY2K/01FbgZeVsZhnQZbWCOlENHrTdXikFt1v0qcvxFoBj9irG2tWO77al8X3x7u9RJ
Rvjxz8FxrFjHVAzmNe91rTpi/hKD8Jz3ts+HcBqamKB6+fiLRvqwZocLbHijbt+jfJCVXuTrRCII
moymBYsWFOB+X2XSdOwDgswNeg6aKZ3ELo9QakAs/XUYnDx0MS7FamcLgQuWf9GW7awx4Qg5RDRQ
x6lbi2IAivyxmQvaxfxil8FUoNUbV3r58egYKdMrIgVuS1XFBJWND5y5byll2UAVyKDSzw4jcJ7N
ryP4DBI0EMoqgP0RcymBQLBUvV4o4KCm5lOZLOe5kTTO8j0auJdfiwpYN+CJiWpiBMc4ciWvBEPB
8jFZ5d9dy2wt534jfZH409oxWZvmKvfevyBHCWWQybZf0PN+05RzL4NON/NDDu28oy4NjrVzbBdw
HJPoueV8qmAa3HTWSesv+13mH5blDj4IEHpeBPXU594gVjvCNTLGxZQL7lndi2YAvAIIdIkoF2Yo
9rtgMQ9N3PdoIg/wnA5/zZsxyUJlVBv5CUwu/OdAXyW46esgzBvd/ZnYTTlTNsOUSPT+vACE0rJh
6iPknNdGEuRnhuZMw+vaRN8OfdOk2zf1RlEzC9Ak1T3LGLhbdnaYsEg0OIM3njACetL9b9Q/JUbE
+yokuGcSBUgnGq67p4AdVEs8JeztMsE4wZ7xyHrc9hcnqOs16PE6GGqLxnTIkn5ktu1q3C8PTjcA
c96lT1o5KkhrsigBRi3H0OqmyuGCVdK4dvOHGrtbsqZznD2BemH53By/dbpglV/tCfA6X7Z29t5o
8/tXiF69/fkehHG7jTa07S0b9nvjHey5hvjc9Y+hsl7WOeZNGO7ILmsksHAT+MLIZQ6NmMmLz3vM
vVN57tarh4NRNy/K9eKvrcMDCE2JgIR5SgIh7JzkhU3jMG7Utr5GTVN1pbq0eYMrdwF6ejU0okSy
+2rl7+amIxq+8IdK0GG6HtQBpC8tOmpDFiVKeLhNhxWwDox5c370MPfEn0pBP1KYS5URpd53pMG/
JekaQJcJMTI1h2Uc36uqP+eNuE20wWQlDyCSQWX7+uZgKxvTwYUZ5vTl3kQmfp2wVPVH9pQOfqgC
0aWP+pTGhL91O2USqM6sloWD7TwJEB3gwhG3+i7cP+I2DNb1aQIGhzEnhd1rhrtgH+ul1lhmmEb5
WFfMu7NMck5wonFzkB0Su0BWbWpUKAjDlcrtLdhMACPRsgBLPFazxaCXlPxn03isp28zYEcD42px
CSUjX1HJziR8uLVwW4g2CAZ0ZBqRYiipDxj72Ie7IyLy6Dd5gKAWZktZAE+TzO56oA+FApCf9Vz8
v+2QG5gHnXLPgWetytZa95mO+jCZGW1Ha62OkdICfP9JXT1/48b42KL6mcQ/RAAW0Rhi3UWL6kKf
5f6opLKtZJFLCGk6eblcmixaP3YQW7VCVi4tJUkvJRxaRII70DaZ9kemWCDfQejQZu1zjGSzT8Vg
La5REYeqa/1ZH1JG/GxhUJmscx2OZKPLutOovuqc6EmkUi9niiDSlIfhsNTFjQh5CT2CuNYDGjGH
AmnWgvhT5NkYyBcqGwt/2Rg/FCTCo+/3/3pi07y3oJYVaqmfL4iNZJVlc3xm9lEw4MmK3/DFMHKH
cHAAVS+CpRdVPdJr/eUoeSWGuN+bBhV3xnpDD7GGc3prcqmWGgkqaUpQP8OjApO/BCWNHeChcCSH
hdo11FlgWfDRhvnKqU5fqpar5oI9zSakTScf1lk/ZJRYRRBbXqE0b5wibwCPjLlrNKZaDpxFJN0b
DQRg+5oWWGT+WHNckt1I1itY4YpQFCLHdRDom+rpfwFFoDtbMcl9AImlYam4vrZWtoB47j11RWbW
1HRJ6e26obiwZfiRA9DXbFdVfrQw3o+ix6PeHpI7T/oljOYMn8zQzNHnASW0sRkZR0VwzLXLH9cr
byO2S24ddaWgLC1Emfwsh1Bze2kzlTgALmYO0z0Wh10+FWa7eDdkekRR53GcgXbVLQjoWE80q1ZF
hCOMFyvVuX25CkRcJ9XOxtQBALPz/jQOb30cHBedyWjz2apP6RtS/wIt0+U0/TeKosvj5r/tP0nU
GXmV1FgzXwmaNk/+qITlMxQQyRyJ6MfeH4IxVHlH9C8MoYKYrJ6P49CrXL0nat5p3wys4o4DdiRw
fKXaWFzZrciBw8ZY47np0BocPJ6cxdC7lmJvC6CEKW8XflS4Hik0ZZD/P2ySIVj5uWupQk9Yqbvh
TxVUic9/kcLF3oBg0JCQYdt1Tck60Qm9BwUEKsTEFAz39KoU5/NdAt0SgLY6yW8jfdgVknje/fu1
5C6dHIfJrRUxHWY29f9x+o0BJWpRrf//3D/IciKOmigxeMFRi5Ubn+RzJmMwguT3wUBUbd0GaVkl
pTPumQ2oFTZ1Hjcpxad9S+9t1Ii3lkIS60tCJjsj2v5rqRtmomqwUHrbvXu+MRLMSJfZ5nhi5QG4
aQ/v8FvrPs2VMq0nohyerc0qg78jWMQT+Lp+hsBPUOD7dm+EcHF/z3eHN/2KBdT+LV6RFPp6dAx+
WyEdsJzA5gHfcwM3EutObzphEtu82x8Owh/IXvxHah/jsJTeAMrBI4CgVPxfROsc5mrvPLl+H4pF
STsP1CWplq0/BrwSI1adjLrUR6ud07Rjaesoz8Iw4vcDTt0DMJC5dxXL3PV9DKQWkKqCFReCTE6Z
sumg4dH4aUH48fxBuwBvJS3TNLrzduPlVlMt8+WRfczzvdr7YZi1Gd4EQSVUWGv+ms6BssKPqGbT
Ikt86hgJXc83sPMasgbdD46q61d/R6tHOYllw6G2nKWhboUNYqcWbjC+6/MajG8YHLVv+7lOelto
HBkxbiJsivl2Udt7DstiQWiLziY7RLG1n0e12KhiRS1WtOAfqgxeX+uN1x5Os/7jheJV3fYN3htZ
4HlvWM0FXrLy2aMm5GihLK1320DwhIdGePZVhe3/x9aZET5AtL+x32nKK/UOb4uuKjcCj08aHXuj
kuBC0gxIrcIJQfj00QLN7kGb8KBLPpaWeQftLpqmFJlcpyZtQAVQ6gB1V1CEgGs3tdYaGln4uy5m
pNFZiwb1s8Tk0pxblNI/Mj/BaPC32Q1NfKwENWoykgRX7Lgaa87e1QksnbhADlqCTRDBmMlLo+vJ
JoU9v/SGMbSF1FH72l8Kwlowo8Y5ZHM28NaA8CQ51NgvHoVeowdZm0AKYpUVVDQwvtCBfQBLX1ZD
Rx8BLG6Pdx/b4h2PVpxPFVYhIeqjUGYEgy3dnE1yrkMvftw1K+mxVf9ZCZZtLoAN1kMSxDgn+w6c
zbMbsbTTV2Bn25ci9uNo67iI8NPFbnuXHomOJW97u0sPKTrbbte8L1ZlSPjWY6SDHoJsRbk9AVzc
VcvytmXSrOZoxXQVSKYJVdn7VuHlh7H+ThuKe8Slaf9me5VsHRDMnKiY7Nj/CGNnF+dwhuhSY2kx
Co+k/sqJ3Vkan0iQK4oM4xJsfY6z6/oSGXTpJ5+p/12TLG+aK0Gz9iSyn8qFAlLNelsCBwrawsHy
yE+aDzf3wY4hhAuHXdixb7OQpr3zV3ZIcCt+RDQXDB99NiPp8dq37np98yaqGyroRKyYD8x1zQvd
43ODedtb7JsfTukZYq2RI86/DEY90fexxgjNS7Kf7eouG0mVOz6buywDNn6A0mrQGJo3ucpoKo3Q
au1SZxps3AgmH5d0gqYKnWGeNds5h5/hIppz6N08zBNXtNlYbX+GRG22m+3FR2ah4B0eml1Vhmnm
mjY9VwKYjlExg4HhPDa4mXBWjAm4RrxhO/57nyEmrgU9s6iai85CJ0qyt5WyZMGUf7nMXvs2AOrF
w3LWZq1JG+H2s+/ZrfDcT3ZaMNxKSWUMpidG8hPkZxEbOgbO2MfdA6JdZ4mYoNMWo0SABOiq7dYf
p8zu9M9umj2xXdYhv8whzL5H59b3yZpz1UYp8Yp4oRmHz4bGPnODfHtybCjYtchwIBAVBpiR3amP
0gIEPyWZIM4BdX//NMgDWWiFtbI1+KIbNR3sT8Ee17Usznf+qFpIXG1HS+yv7D7lZy7QByuA4XSD
ZssHqpR/8Y7GF5AU9wfFvaI+UYJBR1ncJHIpj+MfOgILPAnOECQteZ+aE5vr65mz1fzCF4dD5ZNU
1azdyslrQZNrAmS7lfMzplUtFSpsFQOyHCdFh+mc94V/G8vOqusOLMrRaNcUDuNmFop6H0y5fjbr
ffoR8rL6jNgXYcmTarF+H/Q6su8+fTevQjv9WfFjH5uqUy/tUOqT7TTNJrogtVBqH/vbFI0LVc9Z
mIVvADJqabx6z7XwyOqzPqHDplnlOSIKbt1YvNp6t+oZ/y3zkx1cSmNpTZog6tiuVjkarpmRgHvH
MhQA2R94wusmynQz1Bb2/Jn8RYC4YagjTXsMB/3Fqu4J3wHVkSAEhIxm2darTuWMZdsDp2zdjZWt
i/6tZQk4atDrWxhpiWnhiCpfjh0FPNayynld0CWXqorISwyTUVH/miYIz/U+Ibf5ppopz0ulGX8i
pG9loYFI7rkpIGpLGEELcbKiX6BXlAje6tKN1sNEP4zDsHaSpvGMxbdjphsGn0i1eHXSTovzwQHQ
ASx52zTZYidZz0CI+84I4Zn6e4fS0eHFWa2nYpkJJCqutLFqOrMUtSE9WBmrmiCX2zkgFSnLju4z
niRFP0pqKE5t0vIks4Fw30B18+59/fstUCSIO/QE6kLWzV0GgHF/YLTsDlw/8PvIxCFQ3m/zLOff
Yr0fJHRKVBiPNfbpSSuFugNIUmCsVw5m+KAPjPacDuk1uHYrKtODeVa7rAzZoftUI+y6ZM0Hzwpu
mnonaDk30b72kE8/wpKDHvM7R3fkYLXjQmzaqJKF6Se4w+JJkkRWD28QXvGZGnJvIXwQJ/0JhhHb
vFMkvAcJxbTo8e7wijaBMiQo6p/3hZIdLDnRMviNYSm8f4OJJmZMweFqmHGOmibiEx3TUexoqxyr
8zV+B/XOeXdODma/nNJekMXFO6CVMoaNpp0oM/q14LD19TxJivFqPxbRdHwK0kHi/sl6PTdmV1bg
+Zaw9ta3EJJrBSQ9bevxOVKwcg+xzS/Hc8jzLcVIliOaQJmI/PNhnQGWnKTQYY3dxe3LeeTQaS1+
KJyYEM1dc1XkLp7c1ptE5iDuskcRkxYrJ4S4YiCtKrBFRwpDr30A3qJRVSwiXHIYflyCSN5Wdwgt
aOA2hxZOnKOg1VuGdwGRC4W2Yb2A3Ala2aOZ7lCliKUAJv1YAPWtfKMi6tkJ0pB/cRZ6LWcK+x9Z
wdveiG1QXtxE6KTrKmqBug1MqXA8WVK+EjVnWBjYPq47uQzegfuaKF5jLrR6zuHATenATYCcGvQd
mMWdNmhqPM1SZauGICXmrGtp63dE420FlpPh0osvu6yXjCQA3ls+ZYFqcRSdB6MaCxu5J0zMxa/y
c5+UMqUHNM/jZKbyuJpCCVbgpPQRc0SJjr2dtLqjVL5S554N68cSF2QhQuhibCEdbMTtwfwHixNJ
runkgSjkcHRqSvhHhYRsXRtEVswhv7Uaj6EOSTaHWCXVLkxe1brLgD8GkplGmCwI3Ftum45BGrKw
seM92/XJJOtFkLXzZ1HE9suq/dP9c2Z+ogY5xYUaweJ8mg2qaEWQ1yhz1hTkb9GtuiqXQEN2+VcP
6ZeZutjWQ/LT8Lyf0g3DA9WG/XZUDUKAu7kni5eOB53vpnLmFrL6e5Y0kC4c4k0o4gEOUwuXkAJl
64y6jzA4PYZpJGX6FLB8FdG0DNDtlSGy9EKgEj1vmfgiLCyRPB4nP5NX3uz2dEnc0s817plN1+wU
uiriUMVE11Cpu3GxHdc3GILidsN21beIIelGIiYJ1f+wM8txgBJIRLnxDtkwVLJLUbvJkfUwzgrv
LkvSiuBC5Uf0qSddfqgYTGRcL3ovckknhx7nEMpW0lzbTgwb946H8+h5DklsimpmxlZ9tIjPqF6/
33tSmBWftnkOeQSFOuG0Q28NAKL2Oa/bxo3euTY/H6TYKW4FlSNZ0zDTXTIpbiCsRQ6MhqrC/GXk
sU/Khabs69PKlLzor0+JCUtEo4k8z0yr0g6Gi/qdKUwPkSROMLfy4VVZQSeTBBOGN6pMTQFxE9h4
gCTbkDYFQxjMkcQKvZ0hHKp7XGcEYg4d6/tuf1rY15WYOUOiXCtB7gIOuOpMc/bt/2lyLuHPkPHw
DSG3F2epfwcZz/a1nlzduf7li2P68PH6tHudN57DvZas+IKp4I6QZK2H78m+SpTc0G/TNGU4OdIX
LgOihna/RO3IwM3erbvaYhaJqLcgGml6KUtu5Criv3CRHxnRb0Vk80LLa0vPBFZRYfPZm1/8jadQ
EnVvC+OY3OJPINu1KF6447pYaEcz7Uu8eoUEq6BJnTYMt0Z+0Gp+rLeljIea7sMHo6oiKBqCq2LG
qxd/w2kBalhEg4lnDjzclev1L4vZ4jiH5FGnfer0dK4k6Pzlguu72LZZjOsZ+3dDzCaU7v2SlynZ
0XmZxvJJj0yxaeEoSWXWIw4zzsCK5s+thGd0XI2biRjwUTZ6ZtT4wugEXYObuGdY5hBILITLao1O
pexcOl8mev0OqPlCni/rRCpnnzsM32iLb+deL6uIze4R4ODdh2AOQ/sSlyvKBkHHg//4BSqQEbhz
cjGy9ubxCA8QXYHBWRBh3ITKAjIz0W4dlBn+FnctM9l6kpEZVlAJLKsN01u19NRCY/nt/64OrmJ0
lbSn54P2NjoI1EiVg2XJLAT6cCbtdg84R3Z0m+4GXfDFAnatKo1lZ1JYkHcCaFWgjrYzw07R86EU
itWPF28jJZVCFfNVzkvGofczEqskMr31shRtQYA/PzQfc8MNv6IxgHZ+/bMlDdOtwwMjmg19K/z8
RypLAc3cT7EWy6gL8tN0uond6Cp+JYlylE9v2/o1oDFlhMsgqUmXR5Bb56V+4SPi0fgIcifv0nL2
Zpn4LGF4LjXfKkO316+B/Y/NCHWBmoKPLTh6aNZJf8yrTogSP1dhXK/qdDjD+n8RHfK2F92FHHfZ
z9CosQQ+zDsmH7whLsEh5AYqlWyaYmAVGqGLOYgl1+jvhM72/VmxRRlJ1SCGgeAYqQaC3AoH/ZrB
qT4Hp9A7UdplvSiyWXO0BtgJkaNAVIp9Ja9sOY69s1nHfehMUU0AwQSEszjiTT/u92fDtsRCOdUQ
FjdFtU+iphRXxILGJS0pJBqkUY4nvE0GzwfteEJgW0nURgPb6q3jkG3sLSwAUnxYHCMtQEG1twas
jOyYRVQ4wfSmK8BLA8f5ZeLSU17XN93jn+/yQsus6qwhk4kDrHNZJnxBFpEzi5EHmCT8qV003b62
qTicXc55XQCjZFg9ID8IzZDIRhZWBt+mwiu6kb2ZauXqPCCtdidHGTgVWBI3qkoDjajJ8paFDA7E
ml7PRVcOUvCuAT/Pzx4cuAYuWDah7pIJCh/VxX4qCdeXZr6pGXnILIbqC4EcAQiQKpSWShsWmCT6
7mKLTHzSkEo4sDhvrCx4ozS+4Q4q2VXH2wdFKx4QH0AZr5gW5FMTBrWfZsUwsFk338pHua0NQGs+
t40PLyBr7wG2hp6DolMe6v/DWDnZE816pJ1cyVrtgemTRGgoei7GokaJ3tL46wbAFLKZa2v//gm4
0GlurDQ5WgMzL+TP0hNy9AZdMPodwDNTMEHXUVxhOGV+CJ6DE9QpafsWcVMtpAlkpPxNFCqGTjpW
Ck9LiWeiFNK27YPKiIFEHg0htf0BSu0gpBq88CpVV+VV1Byncq/VW/iQB+qQHuwk69Z5xpkwGPmd
cLyx+XGttv7YvFNEUUVjtBUFO0249jIt6DZQb+VbMrwuelUuO2Vy5QluBQynzzzTxi33yu+D/vxr
BOVXDG83tI89d/MSVB0+co+YWTly4DP73WrJxNueQ72iUHOYSIpPVOIBsEa78BBIc8HKJ1rz4nCH
mITFTTEBx3h0Z6DSqjp0/MxW8f1u5MxrLKoKyWlD3nDntRDfvLTo/boeEWlwTQVIsLB+a3NBj4Fb
dhLrBmfH77tCO4CWCKCyPKDopQgEh5zwxTbT19NGyhnGIpN/qpk/+Z8ppycZuHISp/ha5GHlI4d6
KuD11eaqjWOffY/gUivXDo7SHu6f6BqIh9UsTdPH6zgdDRmDX6tk0LZqFS1voDtxGGC+gGr70lxO
XsYODI3CkvPuLyszElmoOkJLix1rul1Kqmy3WjnxzWmO1AQ3LFOTDVYPqsgRWFJ0QY11UEtVAuoD
Jz43EaBWbgTXJBZx7+jDhB6IdIqg0eOhOcOHFDv154pSvWr8LsM2cPRy02xasxUNEaUaK//zb07b
rU7b741WfLI9PYB6K4zXjXTiYzywYHm5lmBmIkrGS7qsQ5uz2AA6NNpjcJVRikOuLGyfYqrxUWH4
XBchIF55vdqoGpx9qJrcvKR6c06vilMqt5GMEkX3zknol90vbeSsoi2n+IPXwIVTbQ3EdYga5UkV
G0aAltLsbOjJN0m/mxxOoa/wfZwRpLqkXxkHryV55nsOjVnGNxhNciDY3kR0JVXoyf7nJ7NMahvE
Y30igtIZT91WcuvE7PaKtSST2FHoisFPr1jHIP/CYwuaJhcqEYEPpJqkLSOKuReLhTfuYFN56MH+
r2bxqdQTMGgBfYrFmgwkljrKymuhFLvggu7KJ0aqWHmttHnGebL2XGCjNmkAj0KrX0ppAhSTUOGw
v9556V70ThCg7oxRGN4UFN0VqqvodzEiTZetgGQJeOJ0emiCyFmCg6ZK1phm9JBPwkLa7/9FqGc/
TrXEjg/ONuMZP6lrqfzneg72cfu7aO454Q7Lt5GKmYcHvjvNgDolDyh/hRiWMrhW0JUKbwkArHVK
u5HcVMZh2i+eTCQBU5GNBnBlvxMO6+ASqtRqXQ9ypi8vzQBC+4dORXmJpYnK5ecOPGD8BWF2fACm
ntQh1Xxl4MnH6CxF+CSX/hKVIVHJsE30bX8+Hn/KD+Vy5edOi6muYtZTOmi0XNau9MaMbBdVHmhd
mhLMBGIOBaAR6iwTiVONQ3GD0eUpq9klfFm+qwVu/KCpAx8utayqNSdP8SX5u+h+CKjYDBgXhsLy
k+jXXP0uUolM3nkLvccQea9IfNt7rhwD+3AY9/IOeIPnYOK3p73UBUYpYDSJJjvuvW5qdEEywceO
tctYlvQiaTP2yi+dSkbus/ECpN/oP/HtFqvvt3v32mLgyVcHhn1PiVnOVqeaCk3i5He7O2uxRkYZ
phCONRrHwdRlOZ6rogulV6Kdwt7j5Egqy8GwM8YDdWBgAZQFKyUMh/rQqroTGuMZSsRKIxappR/i
CDt+dQ++rEd35paBeCfi1XxNG65dBWMoMrsjU8WH9p8KN3/SfdkjEnF54AF5xphhnNspXHb+DZ8H
W0jXv3h2zGjgud9wRnbUwlbW2kMWb33VFVOMFcHpm613CF6BgPrqcFejDEVoeKnYuoBijOJYXS/0
K+sNRUtGFpmt85cnereOJbUSgt/g1yAAWeOPGR6BY5eJ0TLezLweEe5eMpbKSqoiN0nI+at+VZQf
LW9fhzTDvtqCbKvP0QSFsAPFANUm5K664eUXrGQUILvLyo9tb4+TR+H1B0iUTld7SGJB6R39hq+D
u2Ji+MTPF1O6ouUzOEtGmn8p3uhftoWVbCulFTY1pcLk0jiRVREr7NDCB1a3qniisiGb3qNSf+DJ
zE4xW71zGbvQx9ElBQEaWG0BNV7IYvV6qKBL2GZimmYZ9/xhR4PLZ//cko6N7ykq1yUuGjM+bPYU
4QGbkmPgaADXTodTrgdVyuA0+Hs0n+0M8T/zve6hy0ZdF5p/oLbju4qsa/TFBH2ALXsKFBC+CHb7
LGGgudh6alJVi8ZlhVQEi4D/2qzf7J74WHHyJPNHV/z/tXpIi6wizcAHB5iIKyeQEC1Z5ObERGbS
C+ho8AS0muShSv02CW15bH78/HPx6Fn1cqSQ/D99IqiWJla+qFTcx6JbSCzrWOsz7PtbHYJH86cn
5z/kR5ZI6NY0/nZkbizKvauTBajbBVGBqFiIiaBtsYFxeKfytIPzuoxG5BDIgrVFtyvYzx9mHE0K
SVWT0pVm4gIt+b1a8+YLxvtrIW9631FsLAETl+br7ko9iF4dIu0xjElPFkjjSXnFSWljwOOzpzgl
KkvAx7xWgSnPguEm80Nfq0ul8FTm7QT1TG5OjQWYN/jFk5v8INaUtqmVM+CkKTZAhztPH5lnvJA4
EY/ukOMIWxgER/+YYpzAWEndnLUE8C0FUUyV9NtgyaYUCZ4PMBOXZX345CeK/rVwZPegwQyupTls
CrLIdMHurqJ1Zpi685OVv3PPYRtG/CICmWXwQ3vIZfcmiVj0zh+Q6cgbVkbaPP4spm7AisjT9Wqi
AuTL0Ndi3t2HK4Ia9vxX43mRQFeZtucid4Cxz8ygno4aeaJ8qp9vXQtnTXedL8YJ4zS63OS7hGrO
kg9vlU537T06Ie0R6EZ+P/1usJTSN/i+nSO1rxtAU6i+QR1FzK6uCe6D9dytDT7dKopEoUEjtAan
wyEUBlPuMkf52azMb+U66pBdquMFyJXIyDraR56OI0N91Ae0O9A38cNpIg5evIpOL2rjNYD+VWMZ
brGp5cBC0CRfhN1/fwJ+jQh5RneCWscwfYvmoosVxBxwZG1n1QZrRICLNQwfluiy0pYeHgTosSLB
Feq+rYt2PgqnLkdtUAnyzmHi/yOrXhuKSIO7WqxlKNMIknXGMqhtXx+WK8yyYM7s/ruBBDIym/F9
Xg+Diev2Zb23Xt58fkTTnsBxt4adUFuAx6PmKGSFn5e7vIESHjsKnko/m4u5sfVX2ZLsxs9I6DC9
q+yInIHhqC1p5tQVDppTMTRUqEyiQPfDWjdBuvWeE/LALYc4tP39isdq+WwRpg9YWtX1r0gsb1dU
0DklvpnS4w+NRpGsAzXAaX8EOL5d5orNOyNWe+/7XVkRP6o5NGCjnLvD7rHUQg6tuN3ZUP15Wl7H
PK+KYDigEP8qrxpM7nycIfTyiBRmDRdIcRIejhGTL35v21ne4szJfO56ucIBuK5oMr+hBocVM60V
s5Ae5C2GO2lKATDc9uQEDMrBdpFlQp0z+hVMwt1mM87JVRLQLI0DVWXqTvYiAC7wxKeJA4k6wXFm
+iDxAnVqKYkDfCRCNDd0SXeMFa9bPSltgb6ZHkAV9697iIWlkaak0YJF61N1AEOVPHdFY0iKEtzb
t8pXU3vB/0JcsR5sYKpgcHtTqxCSnmZHBYACCMVNG197u8VGzfIjN7XSIaej1Efy9pdjIT7S+jPZ
mzRsnuqGfAUwYYb/Ays189xfieMHg/yIDuE5Ul1ycoMbFTb09d1QVQtuSvknO2QGw6ZVL4EmzzuW
lTsOISNc09/aqqwItKHT4OV/LpQzQbMQowdyBVe4ybEDxaI6lXCzmrak6Xr0scdBWzc9lK61n8PJ
yw0iEJQXiHDYBZdhSaDJHslaoysaltUMq1AUACdQ9qmkb85I7MPN8iVebRCe4zC4hMYl/BeuMRu9
izqCdBNj/97ejfSvUBYFl8k8Ln2R4T4UynV0i2QXlHzKFkF7Cp+PfQZJ1hH+lrB1sKn42Ax8H2ir
M5gBHmp4iMOs6LHD84rg/rM7A2pjYxSl/7frxboPsuqG/FRkVBhsDV8d+/VlLSGZdkSBg1v8zL8b
YVIw78QTHpO5nvAEcyy7QLUWBqSBbnimJVvLIZyxtVIU8Q67kVEUVhuX9LTXMw1Y2Hi8ckK2BQNs
19RF2pZqB64vlvVFxpmWR8zXjEcIs6mHYAlAACh1TGkf9qAZ27TO0yoZxCNX+BrHo9zYGlEnSNZG
9VILx8ZZPW3yvTn4+QavobvrcA4a+oz4Ogr2rogBxWyjo2Oems7KAibZq6OovKCjNfOV7hjuSTA3
8uY3Y/oKgviWboEwh2uuk+dhlNhU/HRKZrvfFOFsiykP2zIyOJ1h+q0v1s3KSyFRJTLwq46Ln2X1
FqDoge3Tlgg5EcUJwkUkIwTUWq0xu4ZnLGQWvPtPWtgTarKQ6CDbrSvUwUTchV2MSc6ud72p/wIq
Bwc6WDCmQzRobuL2/6uzi8OiQ5URq7docnjE/t9OoN+l7IypgjfBRfNUXNCo31SaZabBxHWVYloK
W9BIEpkMi7Bmr5nRKwcGqKlTTsU2WD5Z3HgTjbbUHwuDL+NxDBsI+MV4h4T4FQ48R/Oh48/b8ws5
QqzfjrrNjySF+jmEhdNsC2PfiYh01jLAXwLEyZihkdcbAOQQyKhCBFEZ9CK/+AtyDla9bdzxWuBD
SQ9z5kbcKLymVCDX/o8wbdv0UGdll2inkK+L1nP83oQABiywh/il+MrJhNO5YX7IUBz10YbfXCb8
rWdaNgg3hAZPmrCTTIMqEDplVNTcHISXSw2m0cL8TkdC7B5gvJCQv92jZe0gaXGu9AK/XR/uGQkg
tI1Gz8FWrcFwzFs4QgZnLX2nPmWTfrwWn67Pop8Jem6BTu/fz5nFb9Be53XTwRYAZEKlM+ErYCV2
8DPp292wavY/uWf93IJyUpqKa14mMGlgKPn21m3YlSAvkCdtg1D01xmnoKAPj6WTEkD7qZX/GnWA
VvtxHV/KLvA5+C6KSA+0HtudNXbufCojlutirbYg18PaEHoAmwYa7JHCap6AYYDG96sMBTPMFLTF
n/13lC/eLIOSK1monaruA1BJpvDuShGdHBahtOxzgvUYCJ14MWcIc0X0ZwT1JVX/NVzProFdaZhp
UuJ4iP12PwaCI033zSytUWeO88OLRyxfxGneAZXcER2gf7fZst4qjpKAf9EF2aadHQFWKsR6BsJb
Q70JM3FpajVeOWNuBq0h7t6vp8aZqZht772wlGSd0iYwcQSvKRSzE32u3XJfYpg4HRfQRbWL0umA
y2y/REVNcQLye26jdoj7Pftb8qURThv/ak3qYd0JwKswJHQS15QMWnfpOnv1I5bGKpGFbQ9DL89m
4SHnLVG1OBGpQcovJJ3e09TXrnkTCteIiOHngoG1zIqVUyD9wdyFcKDNZ7rBfEAFUqVR1iyOF1zK
OxDm/X1E9qCLMd0Eg/x/itT4PENmcyjMFq91wRd7KvO4BCFXEwNY1qXIQSRsSnHjnmMNy6lUkXrm
JmTN0aBMCzm31MsKh27yxhGcH5h6b1kMgnteugRO8jat9Cxsnew0cvZcaxuL3i77mI2GsjO2sOl+
nk9YBABq5qeq5JJFzC2GEASVsQCgnGSkM1bS+O+AhnzT4cYbJpNP32JVTK5Smb0bmJKzmAq0cf0l
NfetPlhzI6voMCluZP4nY2YQffrMUAMAfP9vCF/zuNR5uwItdVXmxru87etBZtxyO1kv7k3GLEL8
V7eOKOXL0WihjYb7XD0FPznyyRPqPgtNxznuqN77fWZ9DAlEhuTWow80gD5tg+zeauGWmEhh4STT
qOMCIaNG7bUZVZcobM+U6KDc3MysGF+TygA+KxpmzjYkCb+voUm7x8Cf3V0hPBAeAh1n3c/bZhRd
bpkrxmbr49d+BuXsR+HRoqW9HZ2yA8NQ2ncriSMINo1ZFshnyTCQBOThNF34ETl9d5v0l+odrIvr
X2VreEI+BhAotOG5XUww29KR9dWBWWq+lnJ7cF33KTCmtoyadJVwH18lrUiY6CZLz20/FKB/YDff
5QkzV1ubbj+YAnIpG+tqoGiccg9g/oKsrSzGaYfUArOJXo428QPiKEAcxZMWrO7yblxB2IRjbRw1
tu0z00/MB24aZ/F+VjYO39Bqmb1tgYOBYjLVTjbG+fFORYQSkwhV2ZukFnF1U5gga916WbQFTb6z
GEZTCtbnkDySE4Rl3kFBEGVsIHfCgSjdqX2pUj4iKMISCevgShQoX7ywG09mDf7xjZOLSP1WdcTj
ibTqSWikN9fUH0SZ6i4lBmuEjr4+3vRAxLgFJngjcj7SZofVaVde8zcsrlJ+pYjhgbGI+mDCU2lu
aEYoDrYbeuA36oqVwQtmSKgDJJVIdvPTRV1XbRiQEuPpmFw/BtCxZOKP+MlKcHHMv//PhMYZzkpK
oWqikGtXw62k2U9BJ+h/WDoJUG4KKNIgGdtXCDtyzhM4CyRrI/ap7pF1sfjPUmK0Rjsxgb36cRd8
tCl2a/8HEJdJAV9w/rccQ3E/CAisAYhLe9k5RrC0qOjv8BIlkz7Zc6JzsWFG0CbpCwCjUVphSG95
bYwphIW6IO1EVA+JWlLsMIPIylpWcByZC920yIUVyB25f/IygzaiJMklU1cgzxC/i0i/dwd6vz2Z
pVNozASkybCw0/qR4nPRptAudU9anUbirf6CE5GhjvPuBUIdAtwtczcmR214ll9H5V98NQWV6FNV
0EsqMKe8g6qo3ebb7iJjDkU6VCQpHYWaPCszUFCGrvrGVWbQD3p3G1jdw0z4xkKCg2Q7YW0BHg0t
57O4UjqHnw1K1cBqJrvWwnyPF7hoNjCKi4E5jCIUvkWw2FvZM1Rd5ovaqCZMqKXt64i4tyhZR9+0
AAx6xDDSjZzBrSx9Adq7qs07v0f964Hl6TzGAUQ6Loo9wnXj8pldmeVpeymKkyWoLZ4sDoinhcye
bNKpXh7qahBG/NRzMybV1UcEP1IsEmI1ckOMl2cxuv2bMAgFPiMeXLbj3525spC9Sf9T092GQhQ6
1a58A1+SEoVLPWYwzuur7HvsJWEhOQT8+mA1LyRLQNRpQrjziEvaBql+POcISvl0okqdR25C6D7O
hQw11f5pD+BfpDPE7kF4GFq/QVMRL031V+kH/nGageyFHx/nSt+7BGrrgYjvd6DEX8UO31YRQVIS
MFCqhycBzjBue2EbC4afk+plnewIrGXGsRRPGsjYv7gmctY+1d5rEIXeK2HXub7FyBhk2mraTxGb
jQ9SprAEpyLyQ5cC/A30IE5/2bJeQ6j4Aj1HK7O6F5t6U84qE0S5/civNIbWOJx34sDJTVvcVx9W
y5YN86vId8NU6AHSf0eFB0WIqHG1OyQJxcs+57kuhOuIBSnwPoRGGORXZd74C8MLrN/aCFMUkF7y
q30j8wdzikubFCd6AfWG/qvMTh+fYB//TLJKhMVUIaFGTBUor9Gbe+YlM/4hZIOxGGPdxMy765NB
dwHpvME9wckrmJ3CTapQo0/u6RWKcxxcoICRC/L4k/I2xo0GsUnadDSiBfYlSmTYzCvXHylm8kgJ
2UThVEi2Y72pMRZURCQesEycmHHyRYppew6Xzh+mo84fHj34DS6XAzdSv0LvnJurBuWmOLtTolCM
g7SVpCmXDic70JZOMK4GhyHF2jX2RjxdQIKakXerz1rvPwoCwvaJTILerdbCgnoXpidQZvWo+GY2
pe+cAmWR7y5nGFDh0mb2RlKRh7yuysS+5MaBvThzX7KxvejwUiH9KF6AbChs55yzBanLk2ePQKHQ
2rhel2lUS/b6ngg0Q56u7rsjf98agqVUWFlepe0N3RcUqMC9HvO105jkSZOnl97pHWr/OmvcRxv2
Ji5QnKe+tdcKLvrVcaRcb2lWoiy5J69uUo6rLN/GkzKezzle1OI2TqEXRzdm2DS1WdZQnF5gyOZV
KD09Yur/q7NRZ1otY3pkWnWk7tyFJuir0HL5S1BVIna7tK7SPhJNzMmHmtPKxmVl0Xmscuj19+fZ
mbdQs2I6VIx9isqeD1W2fv9vFamgWCoR4gSPGp4ZyxiR5+0s3yIRP7JBEaCPbegH+MPZ8hWadEq1
r68mvdg9t8DD7FkOwT0yhHz1Liz27js1MTxuc60usmd6fgCpCvPAbTyD3ti5mMXHbhTKM1DHwgYA
nEEAv0K4PHyc9BPlGmDAeT0bglxyV79Se6rosOOr67pttVHi5K2QfTne1N047rxabZvr1ut9AUbx
1Etxj5uTkwMSqh6JiiR/ZeSNlGdK9/96gKiM2mLy/ADyzFmSV01pIXoQ9z7IWFgz76uOY0l5pGnb
GQ7WHL+P1cWIyKfEb9Fmu2HgQsDlNFUlvW/YdKzhGGVPmrmLAinplF2mA9T3flR323FQsbMNZFf8
4RiXPW1rx9o2mPNEB7aoaxU5xbbj06b4TuUM8Snr46usB1qSUPPFyu7P9196YqE9NzE9vpljvf6K
Vk1wha6GbFF04ysayUkko9t3a1MTCcG+F1pt0y2kUxDuhYx0BVVieDO3+I6IOFKPLrPCDYJG5q/C
oeaKSdsbBLU91sBYtSybEzxc2zu7hYuB75m9z41N9L8+CO85AqU6B8UtpG7hgcZejcNUibq8Ejm5
SVNWLeal6RUaJa3w9LfPydTQ/YFAfL+XNdgl+HZWr+QJvC5Eo0Pc6qISjIbfwIGhsJTRGJbzg225
WnIWkUkTaTfk5GNYMk/LrR+yFEhTqQR3BqsJ1ECxk0KUHXthsFJSESYNaT1kDauJt7/0bjc7hwZk
exbIzU/yawdnG9dkvMTITOfZaQfO6woyEM553nHdeKUQN3ysHaihRR92Azp/MQodcsplCIUffFKt
vXDDtRcsvlh74FIB8zHJi4X8mJIVQhdpWGeck9i/hPPcNO4wDZ2JQsVmSE94f6SbkQ7oomY/1aYm
kvNQanDLwLjnjvD4x49b34E3Xs7idTT7l/eeTXvAIYTnTudlnfcm0pQjOcXL/G3CnQNnTYRTiWQw
UWwo00ch0l/eTX3Bkib3ebBFe0hbm5t6GYlZGrdirzIHvbe27qZwzSumoprysOvDzAFcocSrtVrJ
Tc9m9CCWxTsjhnvnFDbJ3LKn2AtNdzLTTkS7JB1acUjGmyRHzMF2d+ke72vlw9OOZniXjliJwz9G
UU1X5oA5aESLhNWDol7dZ3SDaCHYe4T7wiRELMsY9ho2xv0/xPXw38W0cTGMz57JUsTzMYV1/0sp
Mv4ptYC4e22vH6b099/RyzGfxCnGCZ//6yls1AoDswlFEHmJi/ipWQAFBeDerOklHRziQVeQa1T/
Jb/R7GXbEAkdnyEWFIitPWeVKqH04Y0B4qBp06HG7zmYzqB3KhvcVt8JfB+u+zaCPdojtxQP49N5
iyA3Bybm8ddsXAnf1d14BYh2eiJlw+cwoiec4KwwSb6OuUWdZsM8D+jFV902ApdPlbcGocfip5Oa
X/+szZWAav67huHOp1rFyl/2OMoniQRKqyvHBVDd2bBPwGJ+kZtoyUWtpBl38979t4OzDj6g5WqC
gwzzZfRfyQkdewfrocq1RO7kEXCdb9RJBKQZccSxKL9uQVHFMPSAh5MNTY3slztFraHSR/nZ99Az
RcTworOwZSQvBc2TY6xb3DBzDpAweuldo6a8U/30eJyfl2UeT3sA+EWVhmU6RzQxuM9LFUTkXyHG
UkE8TtuHGpPSMzXrdqoAJU+1N8KBOMYdZmCx03VyyZL/arl6i+VQ+K+Jub2FcuwPTF7Aj7jJTjBe
mTcv4v2hA6fSi3Y9c/YIAv3O2toG66xmkdixUc5/H85D/bJZCe3uZy4UDuhz4DlB+FeBts67utVI
RSDoAr4Iotnx59a5qZxqk3ONBptN7Itl4MJufrBl51Nboyo4Yf7lALRNI78tpWH685aR3x9nMwC9
mzRDqzSfKMNS7ZsgQD5VKgzSiazeuMAzWJVZch7ilvlIX8uPv1PcFpaQGZeTwiWyjL/meyK11KuC
33dwWaUkdLpBusISZrSv3oNDvS32u8UHuW4vFvAKDJ3RBilONi+l6Bt7H92ELP8a35oFOut15Eog
+HfGvie1Cx6c29VWscsS1BTyFyiv+NMhPYlPiLX2tkBD65kfWQlFe0Lh+/IQIvAFeg6lDnDJWAO1
jtWSMHTEEoazEIFCcKeOBjpKAvZzZcm5R2W61oq+OYGsGZaEAcJyH2Br/MGiufimr1Tw7NzZ+V87
yGOQmEcH897aFUuDNjtBqBlKoDQqfJjkKFUS1sKQWdwGYt3XC1VCB7guZraeWwbm2ZXpzr3YBKv2
N40mrkEovqo1UVHoepQYOsVD2A8v0anPsT7byVDfYwEVFYtSebrdf/g/I/Go2tGEhASl75cEwUsG
zFZlcmSKZq4syFNHhsw179OEtCgZ44wxeQVhsYXYyiAAI4B+r26zmU2dTkK/ASMSGljZJiu3KWZM
qw14LdrQxJVuvJpD8GwDDuhFNXn6tVQd3q/c/bCK38m8aZWAn4UOzfSOKlKC22PLbTNIbeuhEbgy
AugLxoHllV4s5uTxbQEnHjFX/QRWBjG/oumY9I6n8Cf6bOMLHz3X0X/bb8+DjMtTKwSHTSZ/h0jK
FXHxXb1TKXeopZeToE8n2BblpUGlq2ycs4xO1rANV/hb1VHl5XlwYc/+w6/Bo546PCS4h4qhM52m
P2SXOqhSixD5zhEo/nMDLU6KATE+Z2VgSodha8zN0gfuXq9jTQjuJmrUkQii15m42B98fSdt/8LM
6p+/wNsAQFjRYgOxo/ePewZ6b43hC+5oR3zp4b87pDQEBFwU4TU71vfkVZZKwCf0ToIQQE1MAfkH
F2kJqL1lBi4y8BpPN9CkldqlwHsFtEPN/BxOvgHsUkzzcAMYV+iI4p5p56uvEl0h+9D9PNCIXAHp
hRJf+U08k5rTyexEK7g/FncSbFtxNlri3SLn9xax7AwiLWq5+8AY3n0HEXvvdfEolwCODx1vjOu/
ciTLPZc6zvv6IX/v5H6Fs2fOrWwArMXuLQyxFNY3HCAiQ7OKD/veRfe6o8UOwcq0z7kOo1IHa68s
Y71uQEEmxfneoegSiwvCTQgeAnUsLb1Hpa8KFEVVX4L5IX/OBeUA8zp2qC0Kvcsq9Zm9mxkDqTiB
vjFhU2M4UYYKYLLHZ2/jzbd+4hH13NcDXlzHbI9lYKDgfDRaZYLqfBi1P+dzeuNrv4nYAiQoVt28
NvGDFcUksUUi602Cv+EoCYLUEd4P1QRZSZAk2OX4uaPNWmJ/55aG2dvCLbxV0lMjWDESkzrXCwkG
BzA5g3zkIElFK8gGi8Vs8JFd4GZ0yrT4Fa3wxm+1QrrVYn6VfR10IOmtR4OgCzQK/8SggtoMNJsD
qBxA+qYBNj8GtVvIfoaglx6rvKC2wA4lgiu8cNbLtG+GLUoudK2wJcWsoY/i0Q6bUr437wGAaiud
f3h0bVqJhMwqtpnFJY/8dZleuEtqwZ8Fh07nShOMSq/mXa8SskTSxZigY56Mf+/cjcjtCJ5VHN7a
qdU/PXuy6gQt/JzUOahAAiE6Uet7QxWOcpICPq2SZFkKk04YxFOgxKXFHiYkH45NRsRcxCgZWFvm
OwT/sd/OArRDFpbKjX42DpqTo2UQjxtbjO61PV0lsv+pWI/+Wqm3h3QshM4IiDSNJbxjidAsg7sK
av53SHalIHKsapm8Gg9L/zqHJylQtK5omSEgukO53/+9Brf0XdjNfTRdDhIOHZ7PFEGcvq+eoDfw
9UvZz+Wysmt1qFVufzDQZAIiPMBvP/kvdcoX4qex0Z4M2AMSAuWCdpyxfvYHIPoigMXDJABMumNb
NrfRER3rTQROM8Yj2NL867ryg92T6qUB7WZLouz/BNdxvgGPdZ9oMbMFs0APjiCg/sYNWmIqQg/q
UKygM4C+dou5yJPZ2FFT4zYUPOBVCzkGQ56PXwOqqYdarWDoc4ZEJBws08WXHzFY1pELIKL8o4O4
5Ro42mvWCk+5QhWiPpjH6JIkh+rGJVZ1WGxpacEUD6Oo/rQDKSKRF79soXnd3i8LBR4m5z21cYlL
8e0duLTfA5nPmh7mptvvfWYMW4rtFtP4TvtB2zeeuZfhpwfqlTT6cEXSddM+3mQjlYoj7w3QTDnW
9QCKmj1+XcCX+lZOOtXTkEmdjqHNMd4RcbLutmSa37cjdqNAQ/ous8nmvZgRbmZlg5b0s0Im/OYT
6EOEQlz5rBzPZP/sVcd6kAMfJ+2cl6WOpusr1JEspifqNAhvQuzssDbkJvUnyN0xlfBRLXoatPu5
e9Zjl7X9K0lC1UpiQYnYG+zOAl7+mjr+fE6YrHKzC3sYRQbw/swT7uQqcRPnIVWETdUwj2T+hLMk
IcxUEZ4kAMVgdHav9mzcQsMvgPlqBN4MpUaKwAaO/k18yQn/PKLiKVZKOzIYKHzB8SJH2gjQpD1h
vak49Lfax56EAnZs8GrP6OaqOd8hJhDMbhGe9mi/z8iLWsvqzjcQsTXaxAT4hIMs1BRDmGPYLeNb
ITgedup1A20EpgEmVVGcs+89BmxCD7o4ZkMjnQO7xQkwanYkG74zKUqbYPwtsHfCQ7Kpo44rk5FB
jfPoo5bBtHdsm15N2GzwaCntjDsZhwNA94CXHPPsQDnINwFPQxsJEa1BRtlMxU9UQnIOcgdae8PQ
3LPNgcfuK3eiu+aZ3hoX2ccVXgKAASbZagZF8FVHYwU4oXiGlHj2vX28zy+RkMYce+Ev0l9W7kQf
EKkN5BwCnL03gJaNlvTZEFrTsxqjftZNLHrWkzhvQhjn53u/2cuA/V2Vj8G28PsKNsG0bIpi1WAT
Vcczw+XxjtOI70D+5ZFKTFcOBbOBE7S4WWOfEG50w/oIxVuFbEt4afBL9tgUHsUmt31aDg6dYi/K
dNNFYNhw9WN0wtUhu1dDcyZqnOOeksmggDRpWWC5kvmADRHEmT8mVI6azEcFeLg11pQpwZa/f/i6
QN9nabNQn1l+LHB7xKmzqFRFML5l+sx3Pt2hGyaeIo037aHwS+Pbw9Vu938HDAobGErMapMBdxP8
9elQiFpmAzjAOVir8Bk7bKKagb1wiQkqyMsfuOiQHz8UbVVnsSSymmVpFYhLIVAXD83vXIwhdz0p
2OK2ljCnQBtjh07EeiRinB2VvqoEWPmoGSmWzRopyFkWswQ5hhkrEibVaAwtW3+wBr9FEwqR7/oh
2F0LnnwAxaMwEml/1I9ihW5qT5V3wEcpa+gXNAixmNr/yUCpSFGGt6yTjhaYQrsgxaq0zyQmq+zS
3hT/0IxvuwDJD9oFfjY0DXUEqGoIjtrRW2z/OwvsqguZykKEH7+SBae+nF4cFFepC/eDz8fqfQV/
Cn5cTwmHK5UNG737q6yLZe6J6gJE3HyRkeHe9tCwCUPUqz4DIvnOd9G3QEWXPrAj+Z5co7GQvvvf
17Y+PWh/UYRWx0axaQ73wfJOfonnjge0rR+diAgU9wQ7ZIjtRD0feyabpkhYC77em7t41BI7UwyB
jswYHgaetgIg1qvSDfGJcrKPVRlpi4f5OTAmchx2WBg8MZmYi8kI3R1WFTXcKMGWFBlPF36xBQZe
fjtxlZt6D4VaVkpOtIcHYiLIdTP+I2lwN3xVJec9RCCj54OBNiV/ZFpotiIy4PhIZklwIZq41BJU
8H+mL/LBdpAh0ABaQvTCBDH4LYFT3MUcwEbcOcDW8oG3mcsOEImqVMx/+GXw9TJNlOmYrg0K6CVH
blSFZ0CAeTcObY/wICfJteQvqov1Pp2R4jHKuZikDudBl+zxBRF45QBjk4XVZ0+HAMDguxJWmsq+
hOkA2sm5JbDasVwXr+3iYZzlz2jsmIgfNqZft384Snwfoa88ID302X6o2/uRKFKOzSyTXwBiw7ic
KJcQfxo3yPn+tM4RjXzUsYo2H5jKm35po5FVepb9gc4YchcCSZPNxlIt6oQfLr1L4toQE13ibZ5y
cWBqc1Y0MfT6GCVF5ycYJhFA5hAdL5tYKVFW8/jdpdKKwnLJ+i9bw+b/ohhwQZaeGPbw9IGQecCJ
yT0XYtUHUpHFd9kv6c8wvC7vbA6aSsE4SCPMmZfrQo3/SXikPvZmWPtfvZ/+xyIPixvUNzcs5cBd
wVibUmhc8ee+Uc+i/5VHPha943E/1ZgdWC4FjlPDqYStRL6zrdFFAl3+yvc+87dRjwq+weWQQ1Rd
x6zPXk6IYZs6vhnofykTakziFZFMpLYK6nlQIoIp9e6k6qQ7mmpygI+URBMZvcCxMoYmOkgj2tVo
k6jRfv6gUbIDQnWT/auKtr1W/u8NVGxJ7sOmcdBEhU8QUj3ZzipafVSSDQa7qQq1puh4/Mr2nWTW
SKHuhdhpTApmWkY0THxavJRw6aHyWtPn+k9K0aa0I0UsXQNGMl3tfxbycsHq3wuSmIXyLiNGyvsH
I7ZSbjiX4l25j1nEmWfzRmXrjuW8KcLBsVZYokzjss/zMH2nf0ohDSY6u0sBFrI3LGRZePYVRoSt
Sv1+9JS3UdxKG0tpe0hU4aCLFWebRKJazCRbzjzoiHfzCS6OS/yyeF4OmWHXaTD6pFkEg0EI90j6
DWjIfWGXKjOStuDMTnJefLeCq4XwhLBSQyOQkG1BD1B8GZvVuJT+LvB4c4PX/kdW3cYtfTnVehT8
e1BugmxlNjeTYdPCnfMF953s7d3hmuT2U1AqsATJzGaAdBGlw4ubJ7Deu/PLoC70eW6U6ugGu6td
aEzZwQpbihpx+1Ah0f/EmLcEx2JZGyvM4YimX5uZN19a9CKkpAmqoPPp4RSAC3lwa1/0qm1Z0lk2
WdMukJdsamlBbLPIeiCQK4U21BcTZ1FbRExD7piIsnTquES2d0FCaAlEdp49tCXSGGcbDaA4Vxra
2eHDeiTyIQSqbHQ6KYlF/lnRTCol8Pmc1QlDs2yXltHKtxVlUGkCsLgENMzY1zwzoIuNl4KYl/Ya
SK8IQC9PMn2+1Fj7jSEHAwqil1GrLETq2tCgmt7O2nUgVLl0633lLNPbV2SvZNGXoT3o4TYkCQLe
OOpU7VnmPbAFtAUCjzLXubl7oR0MljVQXYgjuwaxa0+f/m61+/WI/+R1W4MygBK7Ptm8i4M4yCA2
74pcwSiwZ0YXHWCtuRRkjB1luu6F41RdIP4vKXv4HXoTU/8sKa4S7n3ZefYmTiEDNKqVJY2Y673v
7PIOp2AqG/7o7P+7c+xQoVD8mkbx1+m8E+JxfYelyeQFP9Hkv/3zlEdQPydgIfLMB049etllcXnY
eJXZhuCrV0wJCuDVEtYoMy60gmRPoXcJKh14UPaDOdwhSF8hJGhgL7XQZdVBkc2XQZCZeVuk+P5Q
96X5/J8xy51qxcGB9jvmOlJgQZLcKMNzlImn2Td2+rAx9cv8I/+j1BPHm+wFyG1CQrP97ue/+pcB
tBBcGj+xvTLobJaBe1Azof19YNlq6UTwEwxsFCMfNxAdbt5qBSyU4OCrhPBlGbxsE7lrvLchL540
SULWYi2COP0wcA+U7NaTapr3NcqJaf4n4OO0EXuRSC7wpElU38XQxxysi5cdxmpVbfduH+ywZyNb
dbozbJBqLLbAQt5WO+r8wgKC2wQII+kMYEIQMNco4N2IPjd++VQyYA6HqmC9Zju0T8730W1WpJmi
n8o+h68Ce3W5KMHtvj8RzmSGa88jbwSBsvztLWLT6sfuyl3BSUhqhMnyFqjbdqdfS+BWpA5uy6qz
UpalZv10CBzbrV9p9rUrnerilg5xMGVSbxIcFnG7/wqMVifg3N5VdcTL/67LKC9/x9TKj0kAJ9lO
WGBJiJlNs5sP8yL4E1nkh8WR8Mf2x+KpSlykALGOwKXJDYXPzRkhRm1pHaw+PMhfydgetvDuy/+F
CncvOpp7qNyJMKDU/AqTaNYKSWWIAf3naHdjazAZo6ysAKfyhr+g7g3NejqYCUsLzolobAyQR4q0
V7Sw80yDEsLQ8zMweDM1FRxZO2s00GbTPMEQmix8JYpV2Kar7wYOz/sPNoOvnDpG0JkqEmsKdt/e
Eff6ZbZWF5ZdXYQtNWC/9whkQ7Spbo9MKU9LEERZN++Sg4Q+vf/yXh6rAK4Ysb7F0qqq1iRxqUKW
GbddKGgSgGvwMpTBQDsd6GDQSXeSNIwUq3bGnrmb6oRaSXiLU0pBChKZBeHBXGM0P1Uw70BL1AxW
UCcN/OyGUKe2TY2GsVVUY3KsDS4b+CLNC0gvFD3a0XNokPiYnS9bNH9w0vzDjJjYh9hiL6Qvl4PJ
PQPW1iagRVpyJGRl3htxXg7t5UnUApYsC1qN75wIAyGfIPY1TupmXfsFDQ0zoc7VLsGUb8EwMAzX
R5YVBXMaAj9PMRv3uu0R9TWIgn0S290Ap9uvA+4hci4H2+bjRecDzFsPT40NbjmM+ZO1D+McxRiJ
jf3CT7WSorutgSpl69WNjXfbs9yHy6k8iyHrmIpy/uGwd0kSjpEWa9LSb1Mj2NDSby9+75jfcA1c
cmrDoPwNLZkTgG56phMQKB1cCSBLO1czCAuYTynvJdCySyJgA038G7SqL98E2avx6naKB7YXKdWs
jnomLAE+wdvNjXCB+aH+HSzUyVe/OMaJTZUNzB+yBJuz41BoHVmV0y5b6IG5xOPfVeSd06ohU3Dd
lumjCk0KTw7FWQkcbu2Wx5lal7l02oNmmwzNkewqplwJrlYb0BcK8xKi8GF1zAqdgKEqszRaiTJa
2a8+2pp5D88AcHX1e4RMFGV9O48SfO5v0Ii03DHwQEWW3VbNu23CiR3vv2GrZyIXQ9Pzn89vxjNB
I3Qf06MH/m8QpNptvKANvg91CuAdbInj4iYo4lHcmRXfSSrMyc4Y7j4g5BKU1Kds1U9yUY6hMgnD
gT2+ZakEfEP0+NcivxocPXGqK0tMXMimJGc3uYVguh/OXGXFOG693EYWwXdCRBxEAlyAkLrl7qDc
X+iG7qaHwSOOdmxKAQbb/lGc8ZIIVvEG66aCAd++qWIZyjYXcgZaKNXcjZSyUsxEp7HvbvI5TrsU
7e40vGdtu62swxJ+EFDo+dlGnWL+YPbPOHHCRx9E8+VpBmVpSvFdkfkA+kyqtvJVcdLlj3KBXyDM
KXZ4a+Yl20gaVb4AhFDiNK5jrB2emA6beLJEY7GWbIBPQdSd8hM54Hdp5ScsGNyIfKuzeXc3Wk46
04YR7WInnRbrf91Fd6Uhst50r8wxZ/jv4VJJW7U69Z8EUvtMUkojTjZTruKyWc2OSAZEiyPq4paG
GwJkFu+xNpr2aFaYElI38OKBksbVtgTDho1yEpEkAIEgeN3vezHYxAnrbVEjlMiBeHeN2nluKtBj
KQAsQ44eTt3l39pEpn/KXhD2bfRzbQWdeMPgw5Q655nFgk+oIrFj/cycQkK7QWXHzuw4H5Qrk19H
XxesRDs1NzBFKY3wOrWQHXf7yBwflh6M643fdk8f94mitOyTVBp5GBmGaWadbye10SjVcrqtijLw
ldu6NrbQFTmll3IFmsUcQH4/HTOZK2m9oh0Gt7WjYBuMICIG8r+XmiL1wIkvwg0tA5RDQ5iBYan3
95rDGp0bYrG4TcxCkKRWWd+SAeqag/JJdaeECGbehvcvpoiikEElUarJ4nUm9sI9VGG/RtGF391K
dbQcs7d9I5NpL1HcoZXvJkRvYUpw0pbjR31r1LEFg2icQvPsIkKpgJPyTt0cCdrKQT+px8Vmo3xG
9m2VohnwI0nfaBD2fY3FcHbYDDgnV2PemzoyA7ffuT080jo67/5DAONKvHX++spwIkE8TnMfd1O0
F870LVqX9T+OkeQfEYpHqui77EXMXQNdyxRhJpdeW0JxID4bq0bEzdDIjULPLTNcJhJjxVP4qdj/
1cEq+wdMvfnRBJ2baZ00YrzEDr5umTbyahJDxnovKJcoxwOfnPVJ+Uw/mFxKGftqjWYtQFKvrKXK
8AWLUWoJLsOp0hzPNA64CILxTCbAefdQYDDGl8K0RZqNLChxzeuf9416v61zJDizu+LlMAmx53c+
GWfTQA3qipOeSiq/2+KmwBkRTtsdZBCIl/kr3uN0qnFpQYEDYYiojFzkb0PGp8AggWTyRwv0puAy
7mqzOImMCFkKe89tVFlemHFYbZ9MCjl23qebYrjvinNm62D9IRb/y6W2WOHRGn4liZqu3yHyBF//
f0KEoDtnGMIsuWKm2t2LD6EtXvchwXRBlCJrdufq53iBTkRbLZGMEOKSNSKXQnDimzs80usQ2YHk
oqrClKgsPjyI4wvnts7hJULY8AOIPT7rdWiSFSCYVM8Tp3O2jQbSLx+x4MfRWoSncxfn3YO3CwB8
fe9CyH40LvfX7R2E7Las2oI+2l1MGxOZF1/S/nN7HGzBCgTJqSC/fRQhYtKikx+eeaoS1xkn6lbf
eNhkPz3tL7Mq1jAWmMjSnBEutCX+ABmh3CxWG+HMQK0pVY88yCIC75VAgdi7FZgzo8ppbsnx6+Ge
OMweSwR1ij1DMXqD/geuSV5VXBNQSFj9m9e7vVuMzNca2ewpg+pp+BvARdF+4pSJvGBSBqZqdxUP
1NC9qu+GNbt4oOLH9IM+EgpULGTIjSLF+SAiep7nXC4i8rYVw0e/FbXcAJ2DSOyKJcXZHtdKWJit
RjovPAAAY9jtsjKszGseWPRZ8bZ5WW7bo+3QK50aEN2rXecoaY3F3m9ii8JbLDlp/lR8IPXGh1qB
T7X/y5A2GULzD88/xPLCxk8FA5MChN3cFFU65dLNATBWqiPLlpFiF5hI5AjRpy3Jl9I2ZLoIEOG6
Rpt+D+hOn6VhjqB1YDkWHqaAAfe5i4m4bt/4chbwsrDPAUk2aIiwuXW4V5Xu9IULECf+xSJQpomd
vClKtdJyo5ZgL5JR6HnhQxnK3ZTckiFDNBxFtG68YY5+nZPNRHTdfGRNwPwBqkn1nKbKTRna7d6M
pLsSd9oil7xj8/6SlVA4YJz6aib1WRYLleux3CEcDhGlXL4K6bN1pRKUhB7GE10XOuxZemRc5ljA
q+475U3a1yNoBNUQAeE/hX96GcGzJdR6YjBbfNpqDAWwFdaDONhm7w9rT4o6EN68FNzMIz/eC5WH
TyS2pMVcWzu1cL3/AO6sVCyLYZQhkvwdekAcWz0GVRqViiKYSk4R1tscj6MBPXArlAdaJWpoOQru
GsZrli+qLvMo+Fc0sN+CXLIy6Fkp5StZPO1L0e8QIEmNL2Knc8IGTgsVRk5mDa0l78MZke8XenUp
UkUsR+AJ0ZA8VjKvwiol2xbCt9ZenfXp4MZHqRSVOC4M6XM8VZCvZcSGJ82dMdW2nq0PuOKoUqXz
+NaZHuUOgxu1bcUuTInEfMCFCyt1CQPJnWQFGMoRyy1IZWKPxHBiv0OgQdxnvJtZTmqpfiZRki4p
p3QeyGzHXGAj5jW3h402rzt6QQDiVi2MwEhgguOAbtmc0dJsZHpNFqp+VRUH7U9xdnoD0XXJLnNy
1i3VdaulRe30l7iEfqCMuUU4u4juSjbKsfU/TqXcgNo19S5pCUaRLsS6ZcfEMmW0rW03klNDCMD4
O6Y6B7+++7Yi0y04IR2Lcog8PFeiVkZnlAU5nbxyVWX67pOO71X6lkvJtpZZ3g8muigYT3CFODtz
2OpODnH/00Of4+8OeyVQxxprLpEILSdqMbDVAD6zuK/QXxbXN0j5I7sDFfQTRR3XpPJ/JbI6UzqT
d5azYTqcMFxmXfqt+2jTTxDJDmGW2Qqa92lBD2E2obVXYpp+ESK4mLN/9v1kYJjsGAFRLP9GC5Sl
UrrS7LpXyn/v7fXYvNZxrrSjdDehFvf56NN+3cEshTV1GO7Lvi5xHP9VLMOAW7/eVfascsrZaZzl
pnoUmlQGKZ1yQeW9fxHBxWk2fdO1gdyfW3ayNmiSi/bmEFxFtf1/ITi/whjzyJBN8/lrqbulb+zh
UZg4QJsn3IiQIfVPP1764MoL2Y91DLbt6ekvcbJDNve6SDHkTdxEu7r5seAYMYguOjDlFE1IAg17
QzE2cqaDIw6GRj0STdzH3g7cn52LQPLDkIqMKDdBD1of8S3+SwjcLBIv8PNszqJ9fEUBH73y+5rM
jaTWCEYrjT76/DH2f+t0Svd3lhjJET77teJno2H/2P8x+xKXB1qpMYmq6ZPXM//aVhwDJ6tnwRZ8
RLhHV7K8c2dJfEaGvueKw3GJQBL1QWZBf5f9PiIaxKTWOumfjioRHCXtfhTqTT/X3xGJsrV9VE9E
olD7tIVIdADI2Ll4fzvYFlB9nHTN24wyTFntvVf5E8GXx7Qzs4DgdvGrjLGTYFq1AAY52rgZOucZ
g+4cBRFGGWmwgDuVHO64csXGG9lsjW9CLPpTc1SO9pl3IRLy7ADpFkfMDEfyXq/gOCp74Chql5Yt
1ZU3so+bURIMARnq+Hc1l1QLuXgp2IXAsF5wnHf0uYi4PeJOWGC/oOfCBZo3SjaUa9adUFPfB5aI
q29+44TJy01YPGYj3Of1KbtqkNMvsq4dZtDkdWe/tSHR5Fysyw5XlGmOv0W9FM2gMx9JKNGIXXWp
se1fWrbAwpnw591p7KOHvfHzswaxiasZiaVnVXfskdj30lhjBFiTcL/AMgHMTV8rUCHOmEokDpga
C8p8iHoqEH1DLOJKHKYLNSMIBywHv7hC1xYGMEW1o23JDKb/0n3SbsYAHu9hSjUKs3DASmCjjR48
xYJPRKZUJfUrdmDlqmXdj9MLcfFNxU9sB5AN8HuTf1tVB4op295ayFshv8PEmrv0FDu7RIFZ8hoe
VqULEJoT07pOmmyAjGKni5bs3XRsYl7jyI6E6U4oJDmh30NRD84AzePA0z22dgPkNU24gitBjING
J/3ebjzMWHYskQo5riWYx9fVqVJhcQu1pHgfXIF3NwVG9ETD0zD5JgFJ8ARqOOmMwyxDRhYN3In+
77H+56HkLs3dMaYPcGQuA3GCXfjH4w+glxFuLs25sVg+6uHaZGRE3wvBYqwGckpMWTJbagCsxrLA
EQgy137jEu0hOmVkz74rQPv8xe5Fe39OAexDzPJQUiO+yWgXtHylv34HHI7BxZ5HlEPuoWr6E8xx
lCEpHiRoudd2NSzsV7FfFdMOR8mt+h3+7w/8d0dGHL4qDeooSTThG+0RpsJMZI1r5xtq4FACtIuu
T95ZhkrApmx/b84cN98ORgxTU6eLD/mkEB2m1frT+zoD5da9fIrQBKQReez3H2TZDKwrztREInQr
IE3mcVR9B5qBPgElKmENswipfnoolIp9oTUxlxjwM5nNn6CcVwtWVRME3TWTSY4FOEXszUUoOsQS
9DDIPBi+LTVC0rgbHFyzon86zacXpe0IRWY+aXRMmd+iZGuAcZFBzME0Cl7Wk/nQI/r84sPplrZQ
5rq7c5GQh02LEd9pnnfN5F3F5q8+I/99kbiSuqMDx4gVOvT5EdeN9S2zk1pIh0MzpyWDE5sDZEUI
mpXlA1vlwYlEL/yo7bwJXR+NIY2BLUomIQbfszFw/6coSGCAJ+ByAjtS/XcjRRy3FQF7QbdJ+8iE
tkb+NTLD6+kiw6Ms9oSgcN7qQtnXEXp9VjG8uir9T9JH21TT3KXQzKqzzfPq6HU86rgpFmfrSriu
nxYTjK0tc2GMGEjccBmCXo1CF8LtLvu6hbnA8M3Wi/BJoSlLcCND4bwXyiJ4s4SzYOgEl/8xQRYs
BiG/8FSG5innTtD3RaZUhLDxDB4lmeWWWrtlNoQppNIT2iG+WwWxoWx+NujsDqepNyUL+78JGQ6e
UXXeEPeXPs1InR0/h+OWaksxiaBOcIaLB4zvEOnw3YViBazIR+DKXiSVynu/nvLyZlPmM8s9kXmG
dbyNkwH4K0KXdiYE76i6ag5HGISOmgaoSjX4/RMZY4gDs0mIp/sZ5bLAp4t7WRhyxVJXeiJf7Ff5
E63GicnZ7Rp5tQXv7RAClos0tBU9yZkkdHZcEFRRhgZG5dBeKWRr5i3SNy65FeIBWMxViqTOz943
3bjp5t/nlaV+UUBVJBTIYcG3GGkKeopj4a+fETzBr+WjfbX6ZSooAjSEYvp30gG6iDt4CDEU/rTw
uAq4Z9OZaHn/Ue6+j+pmU8gSRShX6Yo66RdhEpuhQ5QYQF514e0DOoghfIdUKpC5MgBYjiXhVBlL
RriLHD4wZRN6ktOUyFgKkipvm12wdFkL97yO8VedtATrLDUMoy47ycOV6UHEkxIUhDM1/IjaVgiM
nBPb8Sf7U9/TRMwcVUUqDDi6vFu156h2J8ZfnR9gd1fZBq2xUuFGktSw8VHcvgiiy4uPi1WSHw7F
DXO6eAMVGSOcpSpplvxuNL7rAtgnnyZRl4Em+oXB2eWmCseeKBAUrvd+nTAW6EB7bLGpdBqsHv+3
g9rn0R7sCUYwlN9Evqljqqtw9pyZ6co+VGt8pSqYOhRgNucHr1yK+lwnoHoR1/yn5e8IR9vKP+o+
rzpT7nMM2bfmm6seLfv6sXl5hdo2TVfPP6PYVX+sjFURgKvtI//NraV2+qgAgW2pzqUPQVG8hdln
K/071MKfWFyqdh+/UHqHlluqhQO85x2VCP8/6+dovA5OZCaIz4VTkW384Y5bAfGVfq7nyZtwI+7j
ePmcAz6aK42xnpEKdGevJSWyztMXLTNcyEGjObI28wT8sGYtpXO0S4XFwo9R7ZTc/cVVZST6BKTr
xYrJzMcOz6US5RI2ReD2T9rluan4y2YI4+cXTANCd+f9zf8yDHITsJINDDbqXwckq4Os3rUu4Ybk
LfRsZNxUOby2VB2dUOqhOBXCiAEqNgxPwKPJDoj7sE4S6hJOG5wwxkKRiRwDsp1vAHlo+QJdMpPE
vexaxZrVgwcAGNhMVhAb/W+NczpoucwUn3il1RSz94eJ6RuWVv8PFnWETd15ZRev/vB9iRtBxz2x
NiA4PQ7rzhy6FFOQxXchbGa7ukBEvlYEQ/sGCbaWDI90G6fIGyN558anCQPnWA4cu8y0475fgaV/
IF0BnifIwb1FU+QLGH3R7bE/lJyh+sYBOMCk3TN5lSQP46hEDlz+WIngZJJy+kvfG/QumlMxFSLX
hP1CPY1LIzFL6qh/Naqy9v7p39lf/V4UNNSgrUeTvjZc8Olo6jOCnCSNrta/ICjTxSkQ9JNfxprW
mcwYIBk0qt0m4/0rvpivmRjarOlGPBsJcL7IFc3umt3EUshiXt8ZnPWq2zTGv9Lku1mEwc48ciaO
opRUmZS7zfAPLk7igkNqGCa/XLJjZqNwrJr16kESdc45OR2/XfjPHdRwF+e3U05+WwP7/T4/jBpD
I/ajyHjflzvA/nVhcMoUjGE4h1PzjwEvmWW3LABQ5kHh/DiF3ny2SBp9Akb9Atf3WClpkpSchkPV
Iyg9SX0yQywnXnLrQ1DKvFZx5L/IVmK+t/2JlP2YWFpj5XErErAg/I5rQhiQqB8QC7dZWc4WrZQT
ExyEllHcaoWlSaBA8FvbbTc2fHX5J9AYkS/Njq9sUeLat28D528dpSaZmmjhZFvcJ+AYUYG40rZx
40wo48+c7PaE+PNdR9CWEUOYmgNUroVCf6A8L0eElReGnOrm1p3gP6qbDzPmVKrSqyNEDOyVR0My
5pN57yS9CTJjRNx3Ty5qwKCcI5AgoqpZxInwKTaN0H/Xr1qx7RE3hnYQpeYCxb8kcu3ZcxmrLMbk
9CPozaWeMK/Fn9vkdTgzS9KyzFBNmCmkNsnI0AD9UpPuNVp6klF5lu4rMk7mdzZq3tJZOY8NavuQ
qTJH1RHSO2xP+4qkzXw4nzi2++bEu70docjOUmK17pGEZRYqKmuE9hk7DerJc1GCwTXIpZrEYTfe
YcW29RwJquZBzwVcuMWOBQ7eBtMMJleQEZ3JTk7wXPu2O4Pr1wfDXJ6mSBTb+mtrjzQyXmfUV5cJ
gERByCmrLW7QyK2qfsLIg7mb4kffrnFkDrzD28BIGI+8KJ/ROiof0n7X/+NHrjOdUkvaxTEqm6Wn
Ox2SpVF5Y85JE0XlWDYR6Q8nRmg+Y58LQeBDV4AgHuLTrVbbsnKlnoB2Dmfjwyls7vJZLi43x0Rf
Chg/Of5RIjYD5dtFnCmqeSOexjq3xWJ/mlbUk4W0wZs2Eo1PEgHFE+rSu2APOsBXdXVGT6Z1ib+z
RIv9/tFRk5ymOm7tlvqn/j9RW7frbWHa6X8UTnVFj+0tjlEqDOeFURFXZDg4XS+aAr6yLgOm9zas
Qc2Hdm4UG+WRdh0RQuVs7arGByGRJ4V9sZHaLZIriiRYZoHUCPf6w24w6d4sjB6+lObwUzFplK8U
b+HXEZdkbKBJ9y5GVSxZMJUMvF7IA+zTYU0GDTpXY4jGXLPBBnQruNjDBzNeN/9zSPg5FIZN1AXy
g6xXWoeCToJlU3JCWNjL9N4PY79KtYdt9ww8H+iC+H1SESZjv43dvGd6o+om99pZToYNlPEgqVUH
kNtpvYPtHxt86oX/aHLqDWbqD6FsskM9wFjD8s9Dzd4BO2fWNO71CEgP/D66dO/Smb5+jKTwTrOv
88KYHLDiN/OMUPTGsd88F7zj7hR7A0af9fNKdPuNDX6P5qEG7Y11PkgPO4IzuDkSXLGSWGpssjW7
sk3OPCNBjyKBOWOAHgGA5skesWxo9T7VsvZnpqEzoEPwlzi3/gasW5/kcoLfwMDWWAgNOfSF9q9L
gG/vy9kHbH/66VXhvwzzNSuFBL6VfMnzBmieVgmGKJZaYVj1DfW8iRiy4qiOOZIDzb6XpmBs6u28
FERNhqsszlFEGdB50+ssQlqcFwbjUmg7b9tB+9ID1I+4L5fXcP8qTwmloNGwIEWoJE9mz0PzNdXl
CyhhIfFtCnQX+s/gZBgEow/vmnud2+JJrpZa17AoOGNnkMhzc7G8vn74xOsQNHIRI4DMFtNLoxFO
Vy42YP0cBG3VmVCY/k6AqmjjZXtdEOMO5ko5PwBel7ReHf1Rd6I9E+o268QaTOXmYIV4M2H/Bw1W
n3WJa5eSDd8aVrWKRkln3X+xkh17/yoo3cHv/bLj3MmZRdH8yO1b4wvihpfGFmg2gB9WlwmB1Ozd
JZyDBk6xHarIQY0h0NbagyGtSR2SmIVQ6gO6+gKSaabCVLU2WTH/iWMGNR2CaGA8ZP0ZOz7A0efo
WbjvpX2XrwhAHr2rppi0bmwg9lKAgXLEHODdL+Oq0nEXKQ++FnHJGTudNSV+JliGSBI/ybRt9L/Y
We4glFHJ5WexMtp4Gtm5hLLfmTvR2KoD+wMyGBaaiNMggVKMnetMItXnDeCCKOsGvOJCI1IB8a41
dPd3quqQQ7KiDH8PwGOVBuawL/wnAJbBD6zdYdsncCDgvAwaUpKZf97Bjwgp/oQaIO02ZyFYW0+8
5Ub2XUO1eV7Gr53eiOKP/YX/0UH4NmeBE+WmNHn4rStBWmhZmJ2aDwrnFgFN7/O5yK2yEw9GHyGR
Y5FMtkET4BBzccBrp/VdmQt+Y9vclBbHv9o/Aozi8xNeZvpenOlYoIKbnzwAkh4edR/87BF5l5Bc
NJERMsWZ14q7OyR3ekPaZpGLIlpoPrhju6OIGuZ3mQYDqjceKOYcDNgiExEgTT7FPnXW0g4BtFN/
xmRVkh1FDe8gEil+qKFl7L1/E0K613vOHN2LM3r1X0c2KH2Z5BrpW6zn7mlWD4iWlRycScGoHi7W
3OX2EdGYBMOv9jlMF6Vtuw2vY3MAgIGacbV1yox8FLHIlUPclhhDIiIo1xDYF0xJPBv3bHz4/X/7
B+E45dZVg7+As9MO1ikWFNRwjxDAy5xW8eCz3RXGWLDx7pYW1OnZ3clhlnQ3avlxV1gOqCucUb4C
cQcORF3TmFO7N+aBNhSK4/PcPzB2vfRW/EwOpaA6hTspD03grgCwmkcRWQH9VxW/tNDr1XISxjZH
ObjQD2o9QZCiG6rbd7J8bGbZxoDI049988BKF8zrZcp9HEhCtenPumLf5kf/2aXPotkxp3HUUrML
y6MBo54tSX558QtcHP4rqHsBUaZAY2Cg79BxFcSmAw2jvGj0y/Gj8fYt2Opo4p5yarKCf62d28fC
55yvOmOk72DkSzzPQTusPCUnEQO11l78jciOnNW3HXbebbs36ZDk74LBDS92cESGgpg73eYq9NV/
wQ2WNiPX28PacY4vPco1jRTJ0c87JNuI2jFpEf7d6YsILVW1b5/witmixzzHkJu1xPvBf20PeJwR
uNr/ETZdyxJKitWg3tRncsKC5oy2Y6UZFsXCfawzHCBcoGCjN3OQao4qr65/ykYPGMSC7Ei5rw6s
YzmXbsIXBAQt76LC/ZBx6UbuXhfejAEsHAJNIA3AKxlREBOmB0NrijMtd6qatjFyImNe2njDwaJh
7+UbNaMNhCKyn+RAb8j1Y9Lypf+LlFY0WVUjBworbqwvZUjJ8TlI7Tt+UdY0r3M8xV1xcKZmO5ph
lRpq2zCipiPaZy+kbQ4rnXsoVokztcXCaIpBT83pax9UMAY7MdKTIErguD7Emk0p4TtDoU8r2fzW
ezwk5nDcrcS+sYE8uhE3oAN0fH11ADssPACyB357Q0d4MdzLc6tQ7tKMua8K2VOenP0ixk5oWERL
doos6+ny88Kcnp728Dtj9Ti3DSHZ4LN6jhBtXkWi64QLii8QxxQbhAFTl1uq1aeLR4ZkIPCx31xd
VBW1to0FGWj8gT3jNx6rwC6jHz31qA7rqu6KQ7tJwPA1lfbMThVIKdcunGJpTFqnf912+4SUt/cd
QKcWoZj07IbNxkWzlOJgVaqTEpVtaT9w0TFCrDBmHU4Yx6SPwmvxrf/ThNVfOWKas+VbRH5Ap+C8
z+DA/PtQGoJdbWHHA+0qLsylWT/QKdx4cdaL01OPEYz037d36ypcqIaMnnO3AFpPe2tcz+c/Dtsr
pDzcGAx3rz33Q9RyK4gjaa3LFXFeEdlk2lATLl4F29j/Rno203obT5oh/2f5Mf3Cf5uwNypTunY1
LYojkvOqqEUdjeX4a5j8d5yXXyZbYW/kIjXCUyKlEVqgHFP34VLXzvvVlB+gL/uEw3IaMdbk0nCv
pgkP0+DHRTk22FWXQ/2A//7CCQCgLtgvN4Klt3YmshOYrq33nl/8kuxErRv/fFFiwRqAy7xIMoSD
+68HvQTQ6VISP2nPpBmc5rck8oDlzggivdOaPmdlLGu2PbCWAHXjU88yPZ86MZx+z53yMjYiGGxG
RgAqYRlqx7eH207ZZeA76OPT/pgPeC+uulKBQnPNftuZpYnmFQQIX7Df50TvWNmchi4MvvUF7bRM
zplNvbZn7NzqpikDzPvOiyT66qIYy1kYNc1Na/ZFaAlBa27fBr4gleEFKa+gqwX8lwl7Ick/t/BI
gaxaztUiirmNLb6m77r7tw9+GOGg3fd62qqU8mRBM5RmUNPVnI0gGdjWWXzTOGBdZo97NRZj3dXi
ZDOefSI/0a5H8WSCRm8VXlYE9KkQ0P/kgUoFoclDLMJJPZMTfPplSAlvG6WK+Isk9x3sd7RFGiZS
iUQ8Y54b3ZC1Fxcmmz+BZCbmyBqZym3GvXdEBtI4Z8LhVSItD9tdUZRyXynJWcJ0lDb5B1z2JJau
E3V/p6HQWSi8Qot5TYh81uenjdyzdbr0DMStoyvLNxG6ZoL22RRY10/xxZ4iAAg5afnObnkGsxO4
KyH1oxCBB6eRQTsbl72Y0e3/6lkNFDdUuqZMqmq8reBBcluLkKHv56zr/02alo4edWeTFGn8jloU
CCBNaTJRSAbubKmpE0hMjpaKf3cvlnFESUiN/yh0EaXMWIM/QI6gCZ5mLzrOAVgAjtb0bOc/jigc
b8GPJGTjonnUXxp06uhSHB+eFgg7DL/LpvJQ6ulj/TgpxXnL7s+z/ctgjVZAFC0v6n2do6Lsylv6
Jv9WuphGU39DALWYmvUDGZLKMyEfmzeMUiuisQqlYRm9BwJEyM2kjE1oaxIcIchvGLsqoaZQs5Gr
Z/ohodaxR+RtsmmXO7C39+xNE3Rf4OiVA4sP/mfVfPN9uXtm/EwmyRQTFYR5BFX/qIjsS58EEKfg
FjqmDmOKtYSlo8JyPg49CfJTYpP3ET0GZrrd/+Rg/gOtopFzq0gIvc4QlE3FMSsPSlK/8ELpY7kt
TDwfuiHMIqd/h7g1aichyPwEZC4mWZGeGAHt7/6hh8Qu21JHAY+lHnpIhnNdtTZVUijPrxITuA03
fs+fO5eauT0KrFaamTEvxCik0qm4SY2FHSeEIYdkMG0MNqqP+l22mlv5TuUnnoTDOKBVSkXQeMfy
/XZNif7JST2zmk0jcmqhzU+CS3Jqx/Iorklw0t/1TimEqhIzY6TSgaFY9zppPn/PGF9Eom4OHrrg
xWfWqamP2PAgnLfaE1XnGnUlSxyXLbvfJMKYj/ceMfoxMd6o6IxJ8O7W+Op1SAMHoy4mtnt9PLJw
h+sNCKv2TfGFvNLZ/HUHz6oUoZpdNiPYaESyvv6a5rD50jQdUU7MUUCpMYaugid43DgLTLO/BpW+
mkTAZLrb0TaubDuyMXGs0ew0IoAGygbyd6szYPvO8+l9W76Fs5sYRZ4tMYyHzZDP/CdiL1G8dbnc
TNoK8Qdqq11KdoTWTGXWoOKzsIEPb0YaequacerzylJHCWXizcOgqXX/cm22fd82uC4aj/uqe36g
CVLbNZlLKhMr6LN09Mx/OswoRQuewqG99dz6NKU39pzeA5xygF/Hm+t2BKh9f06O8nLhp4WeTISp
v6LxcbDD/5tu21toO3Fnd8By3lht3YiVyyr3IMYq8/0FxutZEM0mgzYtHvp+2xJe3jGu6m5uF8kX
lueCBKCvRSgouwjVVPuLa+/JUQsRAqRO9dJo+VZiLwVL3dUdBwQUy7t3HH9qoKp+eUOfAwWHLXpc
SQYvovJdORHV9NOyujbaWciUcGK7KZBB/u4kJD+HRrFkSOikBD0T3FxkhgcqkivHVAn7DjiNaAQL
5OpCg6OtIUSNzXyYv9BwxPghDa+8WxiEQeinTF4MTgjaTNo/XJxd+wdRpwAUgoWdyKQzi41WtGqk
Hous5jMRHg3o9Tdc+yoFxeCpgq8lHNGJTQGuPJcaFqj0jFvIWm+/ew/6WgAWHirteErSnuoZB0jS
m16Iujfxf3FO8tHj7xOEJ65DKhM9tkSTV8eF4lhzxV3rR3zBycZ7eKfAraFHEdATE7adzlte/CKJ
EpUj4vUNVUZmYBeyX+q7veMBb8muQV1BRfsFe6YZqMqGOFZGYYfqJlxMj8Zx9oV8KAlpgGAbAYZO
DlrQdZC7ypEW0Z4c3YBPLQ11PObMZNIZQ1VXTV1rA8hwEWm62uc1Xmydkhbdoy1zbbt0oqJ+vmUW
XIAt9x0irjGUd5uR5uX8mKiBkkcMGZ//U9zq3pcwJ61hgMgvvpjei7U8YA5SV0Srtt595ZPZRw+A
ysVzcTuo8SqMdpUkMKndd/WKsGvyOIzpgZLzk4VDzMm0d1pAtYl8RLg6d8xN3T4+1B4ELvlowI5b
VO1Bd72q0McVPDBvPt3zX7AcwKI9yBVKRPAqgesq148XD0hksd3NPh1HrsW9k8E8bWzP3NxlIY+R
EZfnnXm6ZIPTlIBogEZxycoOs30xgXcsvgIcbUD6c6hxAVfJhwiPl/S+u35Cw5hqZrmoIKMlIOqy
8umvd9e6m2Ad8+hQTWPax0+M+S5bxkklKli/sVCN3JgnAa43PSsjfg79TWcZE3bYbvNkuewpiyz0
Dk143JcjzyYQIcHVPDSzKgeXc6LHJ9tv7zoXXiAG+qlFVfaxd8khLSRjtEGw8+l3UjadquvlwvIs
hxKZIR07ny9tdoC4/J732QIERyWb48ehciTi22hrNRlH35RGEtIiPt0ORIULMYQi7EPCFifijHGW
3LOQCeoGJAN4GFqeO3bB5R2X+A8s053uMksCP41T69R8uvcp6U9Pf4xJvD/So9CZ3bLTBMuupF3h
ZqHjwH0aBcCnOXwkC2FZPn4UBFN44UkajOOoWcBZVWAkyRuGknvpCtkuH8hxtbYwBdMKlvNK7pFV
iYzzxJYwHDFO/GQYdRq5k9pWSMQQvxL83EY0qhBCU6esKnE+zZecaSGXSR5dWQkNKPnkmCmduNDg
VM71kcAlVFQeKApSr3g10t6sNY8qndRfssM7bYrEWOn/ptox5Cyc4gCEe4gOmOmY00HH6VrdAA9Z
vCQ4U4nXN6fov2hhKv99m2arksc3sNLDAx1XP/L+0er+tcaovGZR/VctCwZDOmtRNbAZmiVjWVsd
Wl1oWTGyXhCxL08D++debxaS2gw/CuFgqfyjccxMXXF/ydowuTwMLbX3r1VcIW8d+uIkAecqRAWS
5nipm9eVAHslBVocQhKtRbfUV8vm1XfXGoEc8M7itd2qqViH8wA9Y5ALD4IdHDtTQTAgr4QP4/ox
mUWS7AMp9oFGvjOfSxXPPS3ZKrtYCkN7kmsz9Yr+Ob3IrCQOti+YL2Hmro+PhNQJwTvp5o4PKpbe
AFSDgd00Xr6QdEoFw+3E39STi07iBGzwgM6tebfYQvm++GY4eyLP9LoZyMeiF9b0uZ2zdC1TOIQI
cOfrzHp/NgNg0LNNaNZeKQTD4/HhGaQLKTUgMIGFD2Qz82ZFA1hs2xOQ4uRQYYauf/cUmf0RTa7v
Ivmyd94TQmr5gK7Ui4mr1lms8YXJs1FuPmYsJTchLeesMuWWNeUkBY27cm1lZYLL3OrEQamqi7zq
N2xsDkUzKBXzVlW1lYZlnXgya7ZrwMWNoGZG3qfztMgkdfacwf376Y77VLdjyIYAw7kA1a7IofrG
97RmJAfbjLwb5q5C9EGTx2e00CvjcUiyee8dNq4t7EKnfGmyAAmJrEsqUQFi6TLRrZGHXfWle+Vq
zfQuL+DX866OID6x/4E5Ywfm/Dmo66XGncKhJ2rsT3dzHkslILiuUcYI9JcOBDFWNu67Q7BIijlF
a2z4Vy3BzSWUBCvebYxVL/rODoRq9krxBi2En0TAkS/cRyw3RsTF6r9KyiHJA36aXnHnDLKs8oj7
AdHAhY+aO4A6pYpsAVL0IUi4LTezDrM7pz3c8jHqvP0wlsLcGmddUYDypUh+DjQ/mXd8LscX5g5I
dGEP77NvTNNqvl5VOpI5CvbDPwlb+2sgWjVZ7lyrE1KXpQSXw+4LWGYE9bcLYcrjMMcSG/1A59eS
RODd8Omx/3NSwLlmFTDTOajtUbp2PXbe2OQla+iZA6RLQ2JeWjDndVVvjBI8ZgAJdcgx3CTrgtZn
Lnwre3/Ssq8fFPmj1laWnUjBONvcdOigx5VXxohvldbfsSPvHHEytPPCe70RGuGgIIYJPQoEvFm0
k95qrRk9oNJbglcukYHTNRJZcDgHymzj6VHDOJxs1r03FrBba+PtUb2ac5wdPBqd9XlLlybYmfU5
MyFRKI0NGeez9kvO9UGUIK+vhRAtQEI8FtWk5N+5aBGg5LQUDaluy1UVm1IX4J8qwNQDfy+cXyfJ
6lvLfYhVSHAEQONAywiVVJ2rXzZz48GKikltpL61ANmk3FSNNjjnFjHm/c2S75qvYrxPXj6CrHJP
5Bc2c89CD3hBMgmW6zuLWpXx8G0/1uMOdUNcwO1APOb1Q6xSquwo8BFNW/cxCXvnPtgLYiktP4Na
s/J8Sqipzo33Wtihu4Px+YLcWsUoxK8xuozORIAJ9EtQMmcWrApIzTsvQgK6rR45JeLXBJ13wCTL
ld2PoyoDLt81l/bxnM58Q78RcaiEXAilBuYCzc+Eky7OlVC3kGwdnMltEpglS2ZUdpQjQAQ4GN5E
287DrqSk5fvrWUUfl6Kgq69AzcFthaLvEzGihnS2AA05PusZ9fvHUBZH/Ub8siHggcEDau+mqOa3
GnbU82d4Z7jlhO+A/l1llBSuQ97M289wzB8Kf6Rs5KgYNFdCOVRvFlx2F5QXxBoikBaU1q5tqV7a
KxlBgW/AFeS1YiX6lUPh/KDK+JEihzyGLKQl87VYqxd3gLkgzCziS816gPFpI8qO/6hcmD6avnDQ
D67Rg4Z3Dm4vGdEyHHbpUQwr239eXmH1iVuwc8dTcjGORwDAfOUUa1+qmkspnTBRGE8bxR51jmKQ
SExsU9frUzmfYGiZ9DP7tv5G8T1cNz3RcXkgxLUt2C3QQ8f8qEaqyucKsjWLWOBePBhk2wXFBB7A
paku50WU0sljpFyaklZHt+xpLQKtbdPE8gVYH76iR52IOJ7BpCocVDPsdjrp+XxqNItH/qScuWC2
c17pMvVAXc6goM3MsdFIRxFSpry7DrZwEhdZ32qqpYHR5AZBdYOE4RTeNbJkn0UXTwuqXBV/pDQq
ESj7sXWhhyATABbewygEbtmgtX9rs0t3Zm6phWnKT8Tbi191FHIq17RBdKtcLy7NIMVXfNrWdCub
97j+gxQaU83E4r3Uy+diOTaxr/qPn2I1/aoOj9OiJXXktx4ZYpvokkjNTyMCvc2b4oPT6LV4iqjF
56O/HeYO+oW5lA5idsGXvB5zCyydX9tpZHtLm3SdrRtEOKpW35GU+fU1Hoe52VJhRP1SCjbCJJjg
WhMm2KqkF+jzCS3AazUSErmpIcEf5GqSWOq/Bj/rg4BupmobSjqWHSdbRjLf4raHmTIyO3k93JqQ
eus8E284pmGwoHR1QcCIsQZcVQdf1wTSxEFaSiEDI3+zoSwriMGPMWRtel9O3AtD9jJR4etFxj1W
0mJs+5WfGfgYAbbUygitERHcEK5uqk1WhezehBzSOIRzFP3yn0KTdASMTkgwBIbfrQYpnH1I7kyu
7Tzn+88rS9XWB3HYXsx3MvOAWO5FxYVLBqplRqyPiHskkwrXZ5deW9GdD09EU+ltfMMPIBrGO4N7
XnsfG7SQLQOte5jj1wh8H9EmcFZ+hq5+UI2Y5PiUlie9mS1Rp3p+wKnsxEckiuzZvk+rB2Vd21Y1
BuRx0Ja1bc+0yKp5Qg1SKl7TyOMYazf8yC9p6QF6xoTnEzvgq3k6hKZgF0swQtnjL1aPMkbeh1Js
FOcaddJtMJaa1ObQfJbvf8718CSsUg3TgNfru1C7uoeYLxPTPDd5dxxSWTUxnccqwAgPtbYur5pB
+ACvCCIBMsqBzLMu8/ORka8Z7fxyzb8f2plZQNbV3vatSGCHU67dlW/LpAInN/jwlwXIgl/jNcNf
axKkv8E8OgxXuY7gggBt0ssIB6i7SUpffAeub92iZvl/bK7eI+Cv30vTsFyg92vhoSAc1m8PtpOW
0T/hCB587/ikBQfsVCNJUNk8jyhVny/EOfSuo1dISyGe+1v8kEMz6MkG8GqnIQuSnxqfPLOQE3MZ
yAk18rPM1O66fNuOOJ8YniRv5pQgn186LJbBfXx4CkD8GZbXHcKYcFuY5ylf6J3TEwC6Ij3zAZBr
vMSdu88Df87HWTKugNE1szoERmf3Y6LAszE8nnPyzTdEaK2F2o11unHI6ep3fEd/dp4DDGayfkqV
HXiLEBvhSrqlyAibLNZ/kW/I115sx5epvQzjVC99EqUjV2kHB26nb5qAPWFfeNebOQjN6CCHJTcG
ZSPdObF1nYbfmclUHyFu7HTfcs0EclQMKDq4Is21iPHyMmMibIg54xADgn5Wfai6O/c8HEgEWc1d
Waqnr7UY5hCPCAVlhtxf/s3Km5MSBJcnJSRfxu0Dn3zFbWInvzGyEgEuXO7UUGjsuUBcs7MaOn+8
3wP9Uk+ifA122m2MnveF4lxSMzEgMupU7mEgLl+pXVPbWNEa1bF/WT0PzKA+1JBWBWPmt4h9NTBi
v0iNk7N9kURi1UdepbzxVsIzvg16tstD5ItFuPJDTjqze7PRMvNqz97/4G9a4GqVZTia6XvXvPvZ
j2St80V69DZEz5NDBooSHGS/9lx846wpw+2aggiX8oMdr9kr39N0mX7ESVznyux3hmygoiwFw0v5
CnNpKN+cPS00OcB6o2bB/SqFG+somOTDjFnjsB9gE42n9Hb5P4BUBoxxDaVkP+n6XC4CNOXD2DlZ
K3SsfS2sr+O85DAqT8/lIwrYe/oPVebd0w3gd1okxil4ZoDweqJ86cWrp5omenJdjzA164xR2DQX
APPMZ1ZWowb/t6/ScFhWFxwnG4elUDlnpC9GBJgmz06mIKzmp6JUJpysEaJt+l8LPaJoTsFGsp6j
aEj2kGwQbuUTsaNUy9TLZYr3G/ZyGIKEBk5aanPSDs+weijsSbPuq+SYe9jn2sVaLgKNlAxjMYxG
g2jAash+Mvna8giygfL32LDsDUZJ0MbFOcK6qu9fDTPFlqEjHht4U88uO/Xna/inE4/42BPrIgmh
dRMkSV4WCfCWY0//FxnZZt4+7+YZZ3Lbh9CJOhjWWCpVmdkfHjKhRVcobCd2rX1ZY4Mex+Mo/yB0
jrr/xi23OlL2FxavIDMTpUGBBvKpmgdtfMTv1YQ9nACGG/ThR599xVYn5xo3QafQTfzeOELbXCbx
+6A9UfdI897SDVnSF5VclbTSt9PMLze0XJE521VHnWUUipOeTe7TFEGIi7x8B7gUxL2dDXHeaFOF
xvml6a16bJNJdtr90poxE++HfQ/kLrweppy47aXdSMapLLKfsL5EI55BPyeTXlEoutGYR0aI2EiT
KudHEWbCTbF+rbVdbBYSYOJYIg5bCy8yyxso9eJCbMKIjt+rixXG6YRZstm5qhpifp+vQQhT8cUa
S9GQFC6oDgWPlhi9xiIW0IynlcgVN1L2rm7ceVSye6YYmHWukMgzIttbtDkRhAE2r3j3K8Ay4oVY
uLPiiE9T4aibZEsSo8wVYpG49bYfWhxhdIE9czB4QPQEjQ+SB2Y7withOjAzE9nE+XFNNk1nf89W
iX6aO/I2jj0SXeBtjiqliVNhWI5K0m5/xe5ug+8CnBFHZqpudua/qfi9nTubzIsh65m2cu4JRfQW
B0+8vAfmkbz/5GYA6F99ODawjBYc1KaQRxmgrPQTeZoL5PmWA9dp43NKHv3lZp2m+1mY51Y7AAgN
Xvkupb1tg2HXdsZRvckBUR1c/oVoQrCj/BYM5lOD29QutxThQZtQ2+IiD2A7T0YHlfEI/Hkw2Bhf
SAt5ZuXMCu/DwsqqghUGrdgNi/c/rVzVVjmD6B1kr/OAaFNGi4uuzGNlK/SUJn+yQpAdsVeuJBGN
yBJPf0kWBcoWcgvv1dKz0XipL8in+CdMqMZSGSuItZrANWtPV9xwIw79E5pV2uPwByNsnQz/PLWs
MBkxS4JnS6bMTc2+aestB564VBsxvj3Lk1UX4N6VkVgveFItVamNEyob8N2wr5npQxthKaT9fIxz
naqmZZ5fMDrgoTu7/QK0SkPdWG+GrndHbAHaSmledh3mFc3EGnZJebVTMiWyZCm4dBFnF4UXvpl2
b4LHaldsAoyUP1yk2w0iGW3YuuxFYobNeZ4srA5jNma8o99JPDzaBDSdXwr+zQIxwJP5BhDx1Xaz
k/VYiah7j2UD1YmWb1OzoBYW6+Z8ZAnpjwU0r/z2XvcLJfoNKm6lkPU6rdOKAYqPhebUnUfMoMAB
5Eml5+3TmBMhDOEb43o7tpcvQO819nss7T9pR5LdpAkuj2ciyKFc93BpQlciNUyaoZdYfBi/5Igo
mrxdo9m/rE2E79hgh1qYLz1yvHRYM7KRFnurp/SDAR896Q6RXcnzx04KtmJgwidsJjlLh3bAKUTR
BxAp0IBYE2VQ6kEiZJqDWQYRg+pSa4QKXB8fytfTQxMcYcB6r/Js94vgKAU+Qu7GhqzfjNZMS90u
Aj5QIA7LWYh08gsDR/N//tGuBskAtL6v9YJ9G9vkhG0TyiMgOTIXHXgauC6usVIsIK56I1gXty96
xTOVJsOfippj+ZibdbEnqnQNTLokKC2/muy10TWuvVDOJNetxLQLaHrTM87AsKMOXWRzrwKTyKz2
eRibVhmFU9soo/NbE0lIATA3dUO2HvLf9i2iv5coZkS+p7R68BYoGnTLv+kZvj9xJXOCRQ7aqJ+2
TyPeUqMnVNaL8rYflTQLJmpMoqhQp1CWEel7C30cUaqNXuERVoKJQJo13h1+oY+ezlGHFfRZyu+c
SSC74PkCctHCmHZNMpdtb95um+IrX0zb/5NGCyifh4tuA6nUy4vuuR4gu1gVNlLHcKBUh2C1IG9u
R0HwrdaQOJurPMM5rIBDjLeMT3t60/mx3m2QdA61X/hIYSGfHkuNnlAR/jqCUwJxWVyTKU44kkN2
OTHPnfnhy0pdIZQFXOgiU2GNyt8ile55tinqe6Om05/CaSk2yc/jCW378pq/xT4fHpSi6fyRZjZw
XYYgCV3oY9J4RGG3oAxY6db9NzFKvu7nHxrhIGlgHM1Dz41cl1ACQgONZSQATI0v4nTa4v8FDpPF
EJMeeDDBVYvmztsdgIO3VPLPsuOI+cGMG/R+Re1oXZ87I3D5p6Zp7/1/JEeHxlFeLfamZrGjsSU1
BLYggw/s38QyJQBzUQMiqSf51p8muq7ahgfD17ciXpiRvV2I2SPHVMIxyd2H3/3dbWuB+yuyzP2g
urgF44zYfUPltU+TsSL3pIVv5pB/MBOb+/cNOkACU8GdYTztTJQie5ICOsppP2dILzXUWWD34z5V
jYUg/plH6w6btZT/MuTtIyDxd1pQaByYt2IcjOX1Ih+NravWmEAP9uLKajGchhCaPII4qs7wf75j
sLTBVA3f68Hc/lJNfdovBq0xZr1JripL4Xn9bD87AjdfTEchZy1CwtB3ihJiJQ2iDn9QmQsFhhCX
WT6Wn4V9jqW9iYSndEfp2/WSkXt8/kTJln21+LwGTTzsSpiKM1T61MkIoaYqfeS2hGQfhBKR+7XH
1IAm7I4z1jaHlbOb3aMPBg6lPg26iHcQoqs7AA8Vqm4IglI9xcDBxQrid0N5amJApeigogKeooSx
PDF32F+FWWcL7GOJXtqPbAoSEW/aRvKm0SaxrO1Pa2dBYf6nvlavxEI9mZNmv808kiizwm7OiyC+
8JkfvUBos4sxSgBcVcWotHo8XLyltkz2RjezoNmpW+8NpGquqa8h2r6/kA9Q8PZkbf2v9ExBGvkW
SRkzPqpIYjptOhOILCXLtVoRzlTWhm/OAFUmXePh/g20598BGqDE7rnFD9FobRUZj+EOfJwLvLlx
ghBcH+0u27YPC294DpDTZGvPObcGhUgACO3TwuBWUEAegX1q+wXKQjub6/39KxD/yXPRdFd7QSON
fbevy05zXnOknyKzi+8n35vytYLA0w3P3nJ5hTzV1walLjgmqOYKsGRe4Nj3Bt/K7ErslhoauQgq
2C3e+u3cplaDbt2mReBE6hfW9AOFbmXGDVNqeGIN7j5OL/kkEzzsuIOoF94w33CtDIjYr7HSPJ4n
1B2fwIyUYrNCDihDtaf/qyLJQshInvbVT2c/6kcbI/K0PwWlga2UVes/Ru2pGV9U9jwZ+VgH9mul
y+2cRd7i7kzTjBbMpsaE7F/h25LWQqyyUMx90j4KAZ/CTUhe/xgq4IgJiCtuMmIDpuB5uk9rCWOf
5ePNX2CjdPC6OAHOYJP6Fuay3NZOQeL8indImcKdv1WCI9FIxZLm93yxHMK0iVZEUMdpndDowXry
omjrtW5AKHV2+51hcWJzVDfnX68NIyD2ONJwSv/f9oPlgHe68ZMWupAM4ORPUtAyIPFQELYmdZdu
Z8XQ75EmjUR4ITdv9oA7buakNmOYpi0zJ2atPwFiB/UDXsgvJN19X+VTL/YJSXe/mGOvRL1cdB0a
TI1jQpOzYmtS8qtni0lMcCzf6OzVdYNpVjrm5nyutIuByPpeUggRtquLU/hTMxnYp8hlt2VZrl6y
2O1TD2ejZu2kTPmVN419Q4ugygMbcXx9ykXfY3RYlyDXdjwQ7MK4Ohem5B3ssEpMlXZ4837LG5Co
xb6hT2eMOaBxdA7lDFjgMAHWPSb/5QlOh1U264YIR5gVpDqBG6swFy4KYtefXbVcKTxYOYdO9RlJ
FG48Y1/6aoYaPl/6mGyciFueduk5pbfCQgNFxtSRKZWxBih8lYSKJMKU58BDZrNkB8yoJKW2V2ZJ
37PvzdQ+tkwFXa5gBbcoeU98W8d0iWacXVu8/pVVrkRoF9epfobIHJCdnIu8VNQ38pg0yQfs3QWp
xH72FbuQbBM8PqepVJxLhxPeFgDRtrpiPU+EL9HA3rtWuj1kotzQKRBZCIhY0wTTpA6zDCA1Gq/J
7v7po6zTZNgRpXn6E4pO73A+NnDka/GcM7HxDd5rBvkRnSrKBJeWQ2cJ7CmMhxOkbMPlQ6+sUVoX
tpt8KrBIAv83V+pjkIUrQvQLyq8RnKe1UcOnLMXVLFtozwxKMUYMpBmINgBxcfSEdLcxKS7nkMFy
A0JNLff+vb6hhh9VN7hjHLiIUkUhu36wcQ8Na9MkHgMXLp42idP0r399IpjWA27qJNta+KKrafTB
g3ikt7HVB16qa7vS1ktPjm4Xu16u15ObQODAGUeQj+kstCE+iWali1EZqrU56RsTrPg5x+t5AOM7
KUlYawWeve6N8ikLPWSEp48CXCwJCA/TsCIJPwQz3m2sy3mFfE0DPuzBnUUvAvQSw1LhtiTlHfOd
PCUWCetzgNwtEgK449PvtPnrxSXSqrmVI/PfxL5Y27of+pW+FgkbV1gMHIa3SgUh37HKdk84ZD1b
AHpe331MgCMjEt8uh49capLrbhhqGyns9fEtQWo08sZthM51AxmDRnPwK1jVrrWzXvkc3jVJPsDD
4D4Oov/H7g9eVtGThvpeLKSbQHNumr6Kg2nN4jpw1Un0CzCql2GctTAXcn4yDlpdSaDQVG8JAqH1
RRhoJ5V+qm/+P3edApIM+0X0AOLi5fEQE1KiZQ6NHtA1PaWPXHs54GZIMksKsindZA2iGjZApvKj
92oY2dFGhm/JGXP5Y0yATJu3wVlkXtnFQ2PIguceR1qTcDJiroY6Qqt0bZRo2sSUAe32eyQdvFx2
Bsq+nXZxA0Rc2zXux0vILwZXPerf98mSwtowiyXeeuqB08tRvUCOLcwPeAWRB0zGwrhLjmjKalGY
ZnZwem6cQlKoMEaQksq5dDPHjBQAJl8ajQ6qvedpE9UexrmrpTGF30MlLEZzs+67XXq9GDVfirZD
ZzbobZjxmI+iCgUm+XdSLZT01DuQCGS1Lfn3/XVPCGf+plQXVTmmOdkbV/tMuPcBPnz+67+wqCzf
Eczj2IwwfWwNa2z//qAjEnVUqXhfXzDmh0+gvBBckoiNUhXH4jsA31hV3TySdkFYFwyzhfm6yxk8
0aiE2iJ2Ac+yEosLpxWWmPf13NnkHIcE9tbYj5LTU4endSc8qBBH2MX+6TqPhnmZXcGCRYF2NRxN
gz9gGLpH0KMPbjPhys1pCN35HTTxzaN6zTcDcRD2PekGzyGCuKABM+nx+ZQNqRQlniufy8rPEtY/
upBJeOl5+AQSRIVwTHlDGITYVYXTarsh7ANkfFS1Px/cr8eazzBy1K9JrdADZVr79OHSERhz70w9
h2+pvs3+NVjMAHUgYl4zu0PGPWEm6GQYv5uy/BHdq/QMWKKXkpF0oyz97TfrvAoeWA5Olx9AvH6k
3k0zVMmvC0GBrLvudcy8zNOYwStk5I9oV6Qc2v6NgBcslifd+3RW0FCWl0nBHe6TdPyup3Nw2Hn5
P27cwQZ7EHHnH6HXz856V6Ofuc8yGKox7nI39+u6q2Guuw8pfIyjPuHSQ5psl3MMzshrJ/DTSTYP
FIgzfIXK6mo2NJk+PgAZyJVAV7fmJDUaIREIDOCFRkJbRGNOK2A5BINnzomjoE5gDuEKW083jcfN
U5qfeT38SPZNFc61ojvplM7bWj8phFwBS2Mp+L3JzvX4ZJFPU61PdOq+K1vIM2mTvrTN80JqrkAs
KNzdzfAejTEYSATaJgo5yeG3UwVNdz4PoIP5GYPYWU9z3XB4b8pNo7ut1sVeqABCigHANd9REILJ
Dk58SZ/GIcr4hi3B//ioK4O50gPSC+x/qSTjDebFLnoDRwH3LhjktEQ+KV+3lmFY4xm6/fNFOenT
nDp5p+kowjFaifA7IHnW1rpQVWHdEOkToEZMRqlr0cnN/DE1q3jtDUmhfxm6IIe6LQ0tu3dYbhjX
P8RJ2xNa1plNaZQR9iWJFI+xEOhVmHcP4mPKP+jZW4MJFtGPXCfI0/J1Qs9CETFpGZ5N9iShnWu1
mhjh0G6VG5NQsNIWZfFZs3BYZYMsYH/SmXo7U2mbOc7L/2kD0gGCVlql5tgezgKvpHdf+418K5nK
zav2Q/Qg4elz27LtUe7L6nZloRqgN5b4Y0wdPJdgNrCDAy0E1ryUSCAz5iGE/iyKuQcPgmnrNsWV
3H3L8nEohXPOIb42r/VaIq3XaRiKqk17rSfJSRoc/JVp75HOvzviyGjyK7JS/fiKMXLcEnY7xXdK
OlWtDhHTrx5v+5hArTvDs5yUTbDUbO6d6aOwbwE+T0UO6G3H9MQhJFSCJC9sc2jjXqAFQQK9AF8S
KOlkK1QTVjSLNo1lla4GUXnoaM04oJHs5Xm5ZbT7e9Uhyez5HxifhAeA/NC5RAXPtOvAYgPgNIGo
6Xsdgv4iUIQNOwI3j0AexmedDd9Ei/GebAtzWauQvRfpW+wu4IRQ4rFrI2zN9Z783CKWB6PBIfF7
gryRn9rQvgZVfpBWl4nvtbJP62LIvEMCuT2KHyNWFWnd8TErsOMKvsx4+tAfjri/1HXpAp26Hk6G
LvtH7FW4YhDDKr/sTe9saWu/PK3A2TlFKhgNjVsHuY3uJ40/fcRZ9s1gxhUAGacPxSYlcBnLm/Az
+QC8LZRwGXP97FZHYWXH7Y/dQLCHepxVK+lpSMYBqlBi6IKRvN0mMje/F36tHW/NGvfwpEoYw7E4
4hyJ2wMaE8FOQCkDHz+iEBjMWCje1Aw1MagvfeQtQieQsXwgsTyaECnWizg3dkb8jBmDU6BGy5Q5
PvfbLjtgU8+QBKDJ7L7oQW9YbhWB7tR0BjmRccfyGFByIhEYK8AbILKDgOQRuJV9YfJ9I7Gcus1p
zTt/yTuDdbjUIwc7awrUKtVJO2SIOrUOkDg57ScnA0MN/JdXM1t/+VNLHYgmMQRyGg0w3RNf7NL9
nLk6P/+cXSS0pmGSQrPnhrRzVZn/gjUANYyKwAgF+77noOyi/qRZm3xrUhWdBa0lb2y4Bvn4TF6t
B54kse2qjW6ZWGweD2rmdo+7d/ett2o5rTZixhoM97mKOMONTIo2Cp6ssWZ9tlrRD6tpGPrvc9Ar
3OrB3NC7PZZ9s/mMKat3SiA/JzgXoIk5zWOSME0W1dbnkFAw8uS1vQE+UGAVF8EryJ48X8uNBYRP
zcKENjB68JFFjmZmTPuFSWQdKYZTbKNrEuxFJgOs/R9Yb4eiUMOmNu3W04gsOLcpy2Pzr4LK2TSW
/q64jlgU5/SYRK/fKubJn0yEt/kWMqguMLbA+q8jmQZraBAL1HtyalXYFEd8oJRgS9Tvjx6EsNz8
LE8HetU/r9mzusQldIoT1+uNrGIErk9dCkm29U+no5aRRhbZZ763MjBwxhUM0WVkN6+glAsVnzyT
suLKZZDPSrnzpKSTNPbtTD13TG5vFxpVpypGlE1JeutcJEG21P4Af53D6Sm9uzw3N95QGe9lCnCK
BdNby0kVgagvAOfNaujyu7EV0LQVbvE7wQMzJDdZqvJPjWGNEjmlYmFx8UbIXhO+gD7yegAPIpLa
sfT46PSPyxg3cdnN2ujDmO5Hg3AtdqtnyscXJbHpjKbCYNK5oTSPDuPr9s0xI779bu0es8cKGyVU
FgETdENqyPEwpBOpphua1SuYIG6QbKF7WADrEUOfYmeZcux1DsfD8eY6gNfRsA4e9T3ng1ZZCNcb
uaYuBUH4yoIRHDbrAEA56VJ/CCnulRBFe67JwAm0AGaj6sw/9HTRkJzJu3jBcZihA4YvemkoVcq1
PY/60T5ETv75FRDiHdc2mwuKG9whrXB57louX1mGWT28qBqdx6NUFNhwgSkwlmQix9tg29YqKd3F
hZsZPOYdmxkVOYtr3U4jPf0abZpQS/AEITRxovkC171NnuPpzbWpFywiJ6JzkAFDsdYMPUqa+5cN
tiscVfFXqmP/Mpqv2klJomZANX6W8R4FiEoDqUkbaJIb3S+6l1ax1baBP7hsP8LcK6xkx4lMpEFx
kamzBzI6J0UxHzSvXexTuZSW/KqvV7R5ki7tRMRBtGjhk+A6toNN1AWvgHqgxfQ+UoMorg9sG2Ps
3i4t0+1CfRpCA2Rbo5nThq49xT+XU9euRNuJjrZBaC6Zqpggrka8oGlWNaYjgG5E+sPSqFSQb4Cx
od60FUzqjanIo3V7aITWOBg+UjOQ6C3VwjOSYUf5hUa+PsmhbST//Mp7xX7fRMP/mba0SYOGYgqG
6cakB1GDpCFOKF7jT/tch6GfyAY3ZdidhsXrFMWSwqCbZ58t4aq2NQWLadQs2Df4b4Ez+fq8ZdQE
eO6GcmCsG4Y2SwYMLxVb23MkHqVAUi4v3m9vt/kmDQ7P3E4MY/DRMGknTvP0bgb2AMuvbWOZwCrC
5q2DYLIZXvayN7Wk634lkND39zOT6Zk+q8NnAEF4H3G5JHJp0caak1LD/1ox5qRNdq0DcsvfrXtS
+st1UGYL1dvU6L1kuy3FrCCjf0zKKqrcCYA4KyqJ0DDt7m46nKQeIcVCrzo8vQGavqNrWi1pTTap
VFVZIOEyqGBxv2u7kDPeXB7Vn6pDVgiYLsK+CtvZ13gRMMrdA8kAYJi57WBc5x5sLhuKWdkYVaYe
sP12+TSNRWzI3MnfrdpjxNPdIfxFy5S1zdoNGOWRF+YRDL2NIMEftEj0LIIBtNVbd2VE1M07uczZ
j99Ucbkj+GXEJMEfzWywlVnuDIJwnSx5UqIKVJoZEscbJz40+L75n0mRLrrGffJRnnNzm2UWvJbe
69vo5eQe3VqgQuy7EIrwTUF/NnBuL4TIL6SqoIb+PmNFGqtBTuCThk7j7L3tgZQygnFXynn3knsx
n1rwHF1YGB6n8HqGBUwapiyub1rKi0cmEOt3xMkloKhOEFUwisvDGsfuMUfTxTqyCN+tgkUBsB7/
1dy+AZ4aNzYt0qLtnswTQlfUgBFlSOiwt5Lw0J6Wu7PExyXgVMfywHlFry02GtjeHv1mponXQAPT
/ea0zPSbgtrD9zpAFOu+y0UkdlKbRHoC24saIOlgxGPardzqVkP21lS0kl6l3m2eJL2OBjLClAZl
9BmG/jSRgwA9ZqkHLGvoCRJKTH61drQNW9EALQqKml+u0voghOG9lHIuXRLf7dZQm8Doo7kvsUCw
kDAJ+JON6PYkVMCFTz1/m6XLuSGFeFdvp4j86wD4GjBt5vyByODMoEne8/xsUqt6GIWSTCcCAFgB
R8tagiT40QX/AjSLPvS2OQCGbyhxongAFEo+LpLeifT8DCTMFT58ZxTISDn/1Eoimnw0ubP9DK4e
H7G4LvmuVHYI8jMKEjH58YxB3SRjvgeT1r+fcLatLs2ILRVDlR29r9BVL6MkP235+/uKicxplgV7
WbYMwFk35oi34crOxhxFrMIHY0ZBZ9giVc62cv6h7HZnHwiWQZrApBFVltBzB4Ajh2ylMWKgQkqf
T6bQ/erhFMoJRIBpgc1Re/dIsnO6rn7qcnM7ApPQAwqmGpp11EeeePqHv4cpEsrWcsKRa4LoZq/T
P/PlewI9FPmfEYV7AH+MU2eGHySuhVR0gZFhIDy6d2QrR5UG2oSz5TfcF/s6I+keWtyKATUQ3rOi
u7ydpTkOyx4z8CDpKOGOo+sWDWW51rxXv0+wxabC3q0JalXKz0ZtLr4PDT96HC1MeZu/5gHhks03
LHA/ckATVYArUgZI0uECNgDOspTo7rdEOuWDHLT5QVaYRJK31K/8wUXYlF66FlsIlEAxd5q9Chmi
Ymp3blrKNhN2aAYDzs0JqtmDdFJ8n5JpTwn05upqzBPXpH8FKG4+OgFkI/NDtfokQ2kcNsLCLMrm
TxerGX0L10l0/qP+h2j9++iMvY7qre5/I34kinViFczNyABpjkIMRZn3hNJBL+TlIJZrLP52tGbh
73ESAfZOi+QO0V4mwsXY3KeleCOvvEQZCFU4wvqZQ4SW0+kLmAnjpkMpsEe0SFDn6F6zs/fvLOLF
BHfaBYFIu3Ey3+dIegh7JHLtjBdNZpGSjNVW5f61wlRnHSHH6odVX2gs0eQV23QvAlfwXj9d6xjR
k8bOdDtxLeUTYGjScr8+OsKs24oH/8tolEq0e0DebWnGy9qgt4KiWZx+AdE7BujaB58iWLkca0fv
HoHSEowPdWTNPHgcAcgj5NVZzHrqjKxn1ccVzDwgtCATNUl9IZ94tgQYn5d94dpLPnCRlKpwjoji
9nVRqu18FbpxiQ95/CqEhvMEASWpRs4WNQyYGd3H4fnstBvyQkkASQHtNtmYg6WIJuHMv1fTMKbE
vI/war3CfPvjHtijJDGwHchF5zrUxgn6GrTQUhRKjx0X8EKipwIZRCY8VTauT3aEAwnZc2LI7tg5
Huzdfcvss7n9thEa1QTTElOR3mZfdvQf5xmB27+fSf7MRLt1+8Bke5McZiuVm9HTTUA0Mnz7astu
IGjHpk7/n/yBb1tMRsvGEXkGnLTKlVEOC4z5MH/fyS/u8BFZPxBO7ORl+kUcpOEiD31CiUUdbNdz
eVohaqUGEcsbvA6I3OLXReNI71Am6gZ4iRzWsjeGoyq66Sklb3pJdLusCKE0xT8NlZwQTvDl02yH
zWI2oKZ6So1HCmvX20Vq2Oiphy3nEMscSTuuOnKiHp5RGsJr/Mu0K/SejU9BkxsNrhPQBBYV1V5K
exhs0zER+dCN+a6B1V5KGO2WRXlkvQn1f+Yy5EJgjvJH2gojE0dwMInfplUg1G/I3OuE6Ndb7Hey
sxDIK3YsVgkd61GH9vCvjxsK0+l3rNalUY6RohCRdEIwN9Hj4OMAjQhv06k2ITC6DK++HliiBlYz
KNxpetZPL00Xs26aMSN29zhFQbjeQhckJT0hIvMAJzVGx7qImKY+BXrCKlBKnfuFYL9Qfqq+iSDt
JgnyPox0svmfPRQ1+Aa+lwEbarAljgZU+aaP1p8/9vaZ0GW+IIBTZI0q8rV8zG+0NtSMNtCmwqmJ
WDS3VMI0ipA9qO0iSNVrPL2QUdAlD5jtcbov8E3QEqgXJqSywJE5O5oUq6G9w+2V/LfRaFhNF2Q9
yTmEAXZEeYBHZqJv5bkHV2jXxrSB8fOql7GXMxy0Azmwxn1G0Er7EoMW5eqQOmifgZ1Pu6PSKFuH
kVCIMhiWayK1i6h5FIJFpVSwGRtiafYZi2N8NFE+7PJGS9L/Kos1ylwWnpr9K4EgZW38ZyNEgqpJ
sRF/zn3Jz3WIsR0SgHaBvI06N9R3vBM4S9iGedVAPOhk/6Wsf2hstKcnBe9hhL2NSN2+IfnhaWtk
6Lxmx2lc/5a5HImAW5WiJ1l53iUE0yFu/U6dXzIb7GK6rYk5zAtzpJZ/7WprrmANFe+bS0XSgl5k
eCx+uEe9Zl6bBPUkpXZelA/wDeNONnbcTVNNsbXmOoULXzKdFDHEnOoxjNvICs5cghI2qqcwAXhj
PRbl0ci2KVm/MpuTTPoXy7nalQrYGi1YvYrIH/DuCC06fekz4NHzNGQAe/9wj7QR+LQXUleoWihL
D4TXjhg11Xla6XgeNBNf+Aia+CuRQy7iAwQAVuKvc7nuwTT4o7VDvgjdGPqN6qYb09JUhQYKHwqw
7y82uuwh8Fa+wlw8tNWHibpbEt3nHLt5SU6Xx7uHuPt/IHOCBm33rLniocsicBYKeRs2QvI0acep
TtmE5Vy69wEe4kdunkx0eGUD/0BzchXtR9xV+OWZtL4CeKw5ywgdLEp9T82ji+avuMhk75cf+Mtu
5IDKk8e82DQLHemrmgPhlj0v9ckSH2bHAANlGqPB/dn5el+2D4BsxZi1At2gjz2EE0p2MEYh6c3g
Ypv7wMZgnR18DYbskjzvrzCRkRzj/bVNEnh2+FgsLi7QHp+qlW8Jr1qNl9pEJLnuHEHpmLZZ5GcY
SlJv6xFwTmdhnZYGIFN75moGIL+HnPnIJJ/ko1nZ2Xde6E0LV15uP0EJp2fgEfGTX/mHdMIrwHGC
E/hHVn4SnG93dZKbGtp9Ru9YPb/cC6pSqE+lXtsQa86LlwmcCwxiZOnfvofJ2cjXveZq3THv0JA+
0YiVz/e7pojeXbjeqRcRJepwr5ZMzrYVlBoXSe/GtMzkQs7Ju6r3tihElsDNI02Ilp2XzrUHbOrU
Lb1IATxZAYxX79ex5yWcshtaQgxgm6yawXnr7xFMUZlxbklE8xz0UTPFRnNQzjhzpYPIFAfNv7M5
jq11XecatXXp/wqEqNX/MGPVXvNMyhVwJ117izvJk0qYMrfyWNYXirZj7JLoHysXSkoS2jWQ2PEA
rMVSIkedaPrEYrzHdBwWHZp3sGJMwASzuhr1l1AfmDWuM1oP9tjnurzt/Yu/H8HY94KwY45EQ62Y
Dn3Ca4wfOdvbRbRW5UVZ4F91+htYKeVJdrA5wSzktba66s3t5IiDwNObDcL4DQLwY6NIbx1A9tCr
DFDrkRe07bEK8VG9y+jGLNpXLCjITJV2ICrnkk975FaLr31TyFR1fZg2tM7HK3l2O5cCTJAdD9SK
s7pcDTYXYf/KiWVXAa46m7Lzcsdn40HYX13jViHe8vZoIqwNivOomaj129+jCDrmkQQOlYZ4DBcC
H/iYjIKeh7UsC5jSHcD+cLZ67kQ7t5xfDYLwXlxZGTBkdpf11AU26ItNe9j5kjmu8YKGok3XZKXO
XgzGaeuIqWsDknNNCvAbp2kaJKZtd8AnviekU1e5/SbhsOSc7Hc9VDQHWoLiaVjxiNRcV77oK4bD
tUSyNp42MIYAplgypBK/O9chhIUdkWTCf5nqkpduathDOekcPHU54ucxBe3ud7hfcLWM6n6+qTl+
B4ztOrfGFRWqPFIg+andSYLOlI/sewp+V+ud+HpXqOfB5cT0/7UyzDv8vEk69CUTNVUl+s+tTqiu
ztFftHn38DZUrAj5TD7AiZM9NTpYWUDs2fzFJ5dP7SktLKfWlpj3BhlOuo7JF70ra8/3WWZkF2uV
OV56lYQolEWUquutPckQahOB7tWzz9RxFjPKws5z0+iomdhNCOeuG80RS7IJsYkzjJYG5//QwN/g
FKEbRV8KQFQbrtOJbsupAZGyC8jMGjFgmqh2B0ehWV2DBvhsMDwVd/Di5fC+mRY85J+hJfziROA3
PNhlIaY27nPLGPi1tAh6D7HCSnv7OIp7IbWJXvNWLr+0Z5YQ07ykGBhpjpov6SjyHoWWvvhLFAAG
yd89ANL8auhR1wwq7iLt5T93QK93NSR0yNxJlX+FXJnTrDYBRuvqz60qjpYlGlSZpHq7oiCda0W8
9CVqyjIVsOXhnX0VrYddRTvVdzebrCb6eGULC2ngzG+MN+jsJPr2QGjIHKKbKT00f/I2LnZpKkrZ
cR4sGTB4S47eJCqrwQpMiXzaLryuccWPwBC/6PceZlb297Vw0MvJtCGEquqanenRIS07kD0R1xWm
hX2T1XSfqXUNHvSt+i8SFW798Mjfd1UzNn4SJwPIhbb7d1h/itHOWYI0AQiohFaobnLk3VRsKqjE
9RllMK7ee4fM0ErSkaegtXrYHg3fWoHMzlPrx2QDWFgkBn19hylr3rl6SvUiUHJYP4klL2v8RrM5
Ca+tMGBrK/V9tMfOTSToDSsU9wVi9MelurHNiTEIHUUtNDYU/ibfCO9GoSMgqNODnWQmBImygRrZ
lct4keYJp06+eL/rMZcpy2BoGxJE8iGdBWI8MED9bLVq4H1wKphY14M9iHqkjJ1zLLSx67R/kV85
TwjQ5Kbta311mWK6Totpfx7PNxH1rIG/masXAiFnZmt/M3cMNxw7bobDz9qfqDGoIeFUuR0dU0AH
w3Wvps2qk+MhvEGTGKON11wec7teEahJBIq6FrKpYZIr555O1DMY0D3b2/tT+yuM+GjcsgQqUuLK
Yp5zVnLcXqdfv7ALSxjYqEGMgfrAyW9/galillH3QITuHLjSJN2OURV+Zv+7rXSA4ifO8f1ueWTt
dusQtMdsLXuDGMv4RjhZOt6oK+5KneVwmBWWab6V1oLc6JTwvK1Ww/s1OPkp6LQkHGqzfDQsHST/
Id19ql9Yu+njw/JvboLls8YSc/iAlLof31sxCUulE77vhaEagXF+HK5+ZWuB1Qv5XRup+2x9QT9l
+Whg7tonZHkl6/8qqNiRfc4tjDFD+4SRfg0hQP4lfSnVuWIycpKAo884p9JGt1Jjq9izKQpPNnbD
GY+7DNolpmhntgqcqjmyolvmDJs4Op33LUp3zebSLJ49LCnNLRs/PrrfF3cPEha47jl9j/yccmL7
TUA/QIN+Aq3gKpirHt8kIoVjKt7lad+/K/uV05Z87vQynqJMwOp9Ucyih2jObomCPe5mE/6B94Ol
NKd1t8zkIb5Dm6hD0dpUtytfHc2iRPl37hdTA35Se4NnBlHsd7WpJQbDCykbUBY89dT5em5BydsL
jk2aUrGykeyhfc9hf2RHDFsg6RxVhzJIzLfHuLdHG5gjr/hTkj4B4yPb/6sGTwJRPp7KqL/8cXS4
GSpbVGTQr41kox26OCGrs4Twg5wH4Pp+IqHN6eRhfuBy2T80Gquetc0Ex4XtmrZaMwu8ncr+JSEE
RtgMmZTAJJ8AivF0WQcqoXe04BjVPC3NyMIjy8K9Pb25vDIvAq7XFAyASGa6DB7G/aPADqD/xnSE
WYcrurnyKL6X0/0OWgSUe9ltJfNx7ogx6J8GSACWNmXV//G/Ok2QS3qvy+laV2fVN0iXSMsbaWbI
EXVzvYZ9t3Pu0NY1bFInPplx+j6GU1ubrbd9d3KM5QBpbOR2p7Y0l6gFFKz8Uc4xtbBnkpUwD7MP
pQGKKgf6iQXcjIiX1Lz6a5ei0nlpN2vxfFaP1JbDmFnoZYGnFuUKzkzGU/5KWwhRtfmhMrPO6z7U
QJrCqyBSi8CUCssCGvfRgONU9XO4/xOmGVeJFbrM2Fsr9IG2zpmoruZ84WW8QxlBhxLF52LTwKIV
58j7DiAJk50U8s6bjox85lgv3x8N4OhzVhsmLbqddozwQ51DqJwCNwfvTdm5CVbZ91iyHCEO5hAR
b2AvQ8uM0XuldVKVhTYVRJaTtr75cBy54NFE+OyMFCY5hmtF0PCxJpc8AdL2MUFogWlIohiwkFw7
ihhDxJfmZPM0x91G8d0ZPyqzO7LG4y0SF9EazdSg0+Hbgn4b6b6zWuRut5NIgH/dVGKdO2tSIBv6
R5PtL5cMaNVbSGVyH1qaC7VXD4VgSw2OCE3TGr6Ro4vnl7jaXhNaykdXCGPbENwU8YPD1VUeNUFq
dPQVg9nRQj3rsqSDylG7nZtMwEy1K0VuCqEl2XNRyqyMi+Lf4fGxE0DRtX0t4/HsgvRiSWl9qJE2
5FdXWWGbpTYMRudH/1XcX+Ixv6toKR1ZsYjuqK9fmBMILBiZraGeGwvUwFKTD3IdDfZngA+2l0lb
wvtx3gDCB0xSdpOp84ai9bougHGf5eM8W/15PQAZb+4KXfYmF5Ktcf3OxJxnGH0ZpQy90q8iRSzv
Y/bYmcbBW+Xcy1kvUHBdae8eQzDB9L4DYnEkJnMsp1GdpO7BT4DQNhYE9j2rRNlBJXXPez8B/u/T
g820ZBddS2I8+NARLh+9V1TptnRjrIak7QBjGSqT+KOqXydS6hsqFhhW/Gk2opoj998ajUjRyox4
Y0f2us3KRla80GlRDM8DHIRVX5QBt/s++UiNse3vsZGtArlVfPDf/gUmWeH8ZYqRPJP1T3nJMlHE
tD+Pv6brJyXi8SW+UlqrZIH8PflvzPGRjrpfhwxZF1XEhYCtxvWrM8FfAKqyrr/8Erpo5u+GDb2o
Cfl92Y78G1r6c9ku3x1Ta5azMA7o8p0z6MucA/s0J0SpQrN5DuMn3LX9F0t2LNV8TYSwR+6qD0qi
949qLFRatXRu7u9JkPusMkZmJR8ofD4bcwiflXtxY2/vQrZQMFAycZf3alQ7hvDWWiVgTyx4azG4
bGnwmDyIN1q3UPNYD5g6vAxaI7WptEpwXkX5pV30M2AWNabUg76Hlj0yUQNZsuVxHqHl9rVNocFu
KHHxCA3NxiI5cxg09GhwefuNeT5pWTUZyWOlBjXedA69d8SYk85zR00EpEGYcczJUcJVmWAZzfzP
O9F9iJ/nmNGo7IO1q8aC+Ps4HkRPJgaY6RVicUYL2ItHvEwWdGB+aAq7oEbZ/fyPueVeZzX6NyYi
H+FmwbK2f//Js3dGEud1BBHSUCO55UJJmJd/IePXTlF664ZBkjcVFuHwGNk6FedtVWqvCeMqsiSa
0d2C6WGWjy75s/uXCzlMYcPIA7+8KuwQhfTW4ATH0AYrw9+03T1CfPqlkgq2VioWYQEn2VVJWiMb
PrklR8S3pi6waE9YddRpuwr5QChvflUKEDweMOisUpW/EKz9P2H0b8hOhhJtJLtEVbn0QjWEJv1C
VhMCt8PJm2vsrY4I0msvgFYWtDGQRDrGlxW+p90owyuyDTpqLXvjTFpRTLg600s9LBAhniDMFOeN
+wojgc3ILsMFxRozGiNgvaaVakNEz8qoMumL0u4ONMG9CO2Hry/YczfTmQQygSPgwmjaupCdvNK5
TEkVNdXKzO/1PP5u6ml/8nbnJQ5Nr136BAco/YWPD76L++M8GD7g2zuXEy+9TkR3xKkjGRus9vK8
sPctTMHfCODeylXguI/PUe8qOFTDYIgVPKr0ZK/tCHUuYceMr8fLKXmUm+uMWQCnYh1x8wBRbo4n
h703L/DRr+5hIXHP1qMUPHYThRCkYqpOWX3ayDWHCFMKufKfG4QxVx56nYOCdfJ1ms57Jl+lTCZU
WJf1ph0/gEAsHRmXlP0CCL6q6MPjMdgkiYrAKvcQqD6eBN7oGN0M4AXkQ+SmrWyjy4EefqYJr3zB
WSJMdSUD6V2STFW9Ma7vnHjKjM8xv4nSZEjMxbJXj2x7P6ms3IDrpu35WLRYu52W+UzdgruqTJlb
sCPFOVDpN7PFV3Ska8Y5Ujhd3fCuqKhLpWXFEXU+inDZeEGMDCozOx3NqHP1e5JMgdapxg3ALW9y
LmXFaXk/0kH9GfktaxO3OH6b4ph9Y7B8f2Q6Zs20dUvsfL68geyXA0iTRGc7fymlF4STZosDRKt3
qyNxJyOonSrq9QrxVcoFHYszCuyRaZrASTvhXirrwjTEbZV/Lc+0+TiVbkSb0Cb4TNhpLdVYA8g1
Ag2DinJXZSnu8+tOARJkd0XArRKcMVx/yh46dQqs+piF87g1g4/d/K7zG/XoOxl/nx1KoaGvhsQ5
cyOgF5oZBBHW48MvgkmtOSa6L7WJBW132PuDNOO/5QSPopV6AInLLgfTeD4CRJ6IIX57RvyWGa9K
rPO7FwLIKry0H+aVHCJKmJ4jlRtJAhJvlQk0/US/AqHuj7T5MoCHKwtsqsPqgB0lvoUhtvKiHIx7
Qp+VHDBOEDAipn2jehCx5rQSWQ/nEgWZpdqiYOUe/FOLY1k+teGJHYmGQH0F756UtFU0re/SHWg8
PI/mwkp5s2SA4Ajh6ioziz4h1dazDVGBNBj8UxGoK8gOSGfHpISDJfd4lCSc62aOwB4+Wv+zbcAw
ld+P4yvUB4ChH+gkt9XMnVxdZw3jvlpN7VzfsO9oiCSeUXImjJb4ee4fl5CDHBXcs/VTs0guIYMA
ZFx0HXe+50nf+z3sHAcBnsppoNipnH5QVkTGz+9iTRHXGYgU00pzfq9n/qx+2EpqZxDFyoscueT4
lU660aHwt2SsaB870c1qBC4W2jSuteib3+yKHE3LdZ4aiuszl53FUcu4AvdvBpyIA63lKYN55Boe
lim3FEzEXBcervMsu7ilQjZUMZ3wkNjU+Wp2ihS8eYrz7rrN4YOFbcNpEevfMmWFiEkb4NglbqRi
TU+jYYAS37GtGLAG89E07e/gzXwzDpL9c7RiQ5ZDx6Dimt52GezxjSXrSqP/a8Y6BMiRHnZ1T23Q
9aSshNke3HTq/JCsljqf8YVw0mB2/9/PssgIKHB1fzzPvEnfHhRbcXAvYdQIeNa8O/ZC9QTzdMj4
BKhP7JNsFVA2RxRZeVO8F08O5LALkhDfo6z7jtE0MA8egunNDYLQBnHj4JdMHuLExpYEyHJiubtk
EyJQJ70zNhFBysfWXmKbQPUE+/DdRyFndeU9ohMZE+7vLmUs1bCEJufhTfY8s5DjWBsZrkeF0ige
w1n6CiDWcjUP9JbssQv9eBdypI4liSPnBSEeysCZYJ0rqweH6XRUF8hcMqkKf3zLg6ejKRC2Zd9S
X2u5xfkgk+xnAlBfHxMfjEHZ3SfjE3EZHxLo7DJiDFBKNzCHo/uXeeoNTlXLMh1J43N+98fIsm08
Zur3g1b31PKuO/1vQeLTGNVZgqujLKjUzc/O7GtPZpEA8ZfaKo1KRvsX58X32iyHgN7wy4M7VUTJ
jJyheXtpPCI8WcUx7voFP4xbqXXGgcxTEAUwveZr5vfe0AgxlNQVa+gn1cg2U3FY9Y9hY5SGUGPR
QoxQwqU/DV4HbPYGDXVifYwMdXgdFznIw2LOQ0O8qbDXRUfKEqXnkV9gLk3bOx//hQFezK2JPQyq
7Hrdt+8mHRVvw1NbJKY8SLxHEk34PbVGZm2Q8+ORDhp2rAHQapoAlwFB5iQpX1m0u582SoBjcPRy
IlfUQh9sZh/YCvKATrgoXhut6202mo0vozDo26GCkCa1/G3u0xnnQV5Y7umBP7pF0GTw2I8UMHQR
CZYDkTc0NxHQVR2raIBNyhBO1e1Xtm2qTnpe7ojsKMo5pFcRaY47AIgHaF1sKXvSpALHi0j6Enax
qPoW6Y3gT856s8wbG5TTjIpE6KxrgzGPa0OUShjcSoYG0wYm5Z6D1XcCX9m/VVc80ka81Wl1E0HL
SR7ytDP/SO8xO69yFqqf5O4BjlXjTvxy6kfBbZnifnp2pRMaVWf2o8aUV3cjEUFpRD9eD01OKGtB
6ntYPL6oRkfOwR7L25nHTj9/+MCR1Lo7MBZKAWBFYsopTFkqzcbogPP/V6+vi+mSMVAospbLrtwu
JkPzV2aoyyy8v5RfsDjcSXpgeSw7yKHnqpsVn7O2V1JkTG+x/hj1xtniOpG8KGYvKnJOCUMO84jZ
09Lw79Jv8viriGXwKJJhU8woZru45SaeJVZswbuf/fJAQIE3Q4Fh7Jt4zqMpUgsouL5wSvlCY8b1
G2zJi7NQKK6+QllZXjDJe76QwrG7eVR8cxs2xgOxXmlRcYZs46917Mebo41G1qUBJb8by+WV67yF
XmcvvAd8EFFaQrV/3vtI2g79napY3z3864M6XOytsln9UzMcUe0LCHuFJnYd4BvJTEJnnLWsqu+e
2jvLPkc5FgApI9EE7aEKSkfHUXTrVh54Pw3o9I7v+KGf7Dw004QwX1vDexnryxfNR69m7EYJpWaR
7Lmy5qm2HGF1SBI+JKO9uMV4TRwxS/BvdGY5P6O++Q8igUkocHIFqzsY3NIH2Z41vwqGsxKB7T74
P4mKpZONyRokzoYXs2xhvbAI9ICPTg+1cfUylI87TkGFLAp5UJr3qw+PkyO9i5SNod0zDJRxYX7h
epZpts5mtCVjyVRLbn5pSubeU/wY0M+iBEmQGF7MOjC1qzdE834XfjOtg0tP4a0gt56ViQW8rb2T
iUgILaqdCF+S2Uo2PpXp8ZbAADZNsgA8AHd5AKETj5RMiYMk4p/ZdkBthvq55FshM16+Zt/VT3Ov
aT1c0VmmXr0cmPiPq234rPh4QomUwGUhUrRaVftdkVIQINQSzq6bylfbvS+jewL8XtFDRON83fF+
g41JowIFHKshEWNO81FkaZJDI2baWEgqLC99Bhn6BWCK6Nj4gmnR1Jbs6D5+mfxX99PHWaRppJd3
SwFrt1htitskvz7M+jif7tfdBgb1R3dpGvrv3Jc0o+12xceC5EgGtRiHI6swCyLObgpcPvl/+89V
lqJswS1ZpL/QrEF7szPaTB5zq6u/94JeBNY6ikIJ9S3SP+t7Z3rIffimyBe/7vWFJSevkO+a7vUL
oa/KevUWNJlzI3mH/ySdqasJtVU9VD1EVgY1dLlT7Da7Krx9lo/e9Nzd4Ie5T63wc6ih/xtCl+C0
N8eW+WmruefGHF0ecakgkqwWoAyjMNXzt4wanXfB2cYZRV36cQ1bDaji++tz/kNQQMDKa8/x6vf0
4h2WPINnTTX3sqW6qJpkpMXQt7GiCwTgHChLpfMcZdcCIa6t05g+vj4qK51Cm3lblWnDHmLTfn0m
mvv2wEJEltswS4oqBKHJR71yM/BDtZbQbqnheDyEWI1pdOmInhju4tjcVeca69jRC4NhhbRlsSrk
Tt2mWLDSPZh3uVoH2dnqIRpUoAGTP4Ciolfvznmx2GuG305HOYcbo1aeHOelUTsszu6iDQe5ivUC
c2wIeWgJhmMyTg3uRhnWzlYcXqCVeJwhJJpTe1nkrrygDujxn5bUk7iLtcJJc4FBzpmhhpEPVBcO
Hhp+cF/w3trgJbEm+bpPFmWFBJSWnt7PfueGB4EA3Nuvi83aVkwn+wgx3PFOcdfRABpQhDQ9toMB
tGJghkwkoHePeHFVBrnDWPbbSBUbebnGbapMoI5QYNy6jYaBT3yKd5I0Nmu4VYoY6JfsebhInLU9
JuqdazxZscy9NxDTXH4hSiJsC3V9o48ITHFoXN5BTGxMuZ/ZlqVwl/ypsg7VZ5TSfvAWkHH1Iji0
CmRPOQUCcrMUR9PsjNQ2+bMdZMsdyPrVJr0+oBN8OfTgmZwnVoIANVJY3KK51FCRHZJmGRXq1xsT
w6z3N7ZbRxgA93BDT34cv+D9HwNMcihZjE9fe2cyQugttCW4h+0QtQPFXvdgYnxK7jFZFniRZ2vb
6WYyTzpfGE6QCi7L1XFeCNxU1evc3qHSPX8JwBiyopOHE9MeAtswIjfAxTrF80WSS85tgZIih2tq
/6ETj5zrZ5YzKz1GJvWjmL3/7X2LOLsEPmh0izh7RSxP0n7aVJnnCI1W+Yyt2XTyJ28R6Hy+wvco
edzUT11PFtCV4qdkqsYqR5J88LJ6Re6+pnR/w41+urP2QxQuZlSfI2Y561X+D72/gT+F/yXblH62
nW7lutoqV22Js3A6qXHSn6AX+pgitGv6oacSgpjL0NDP54Kaf08JGph657x/K2D7Ls5hQX7vCxnP
ivrTBt1zTAUHQ+6szoUGN5Y/KF1nS+Gt/SenRvDXAQoxafWPaGzjPmFtXrCKr6PBCva/Nw1E1rvu
Xfm87y/s679GC3mCITDlWmcIlPgE89BUs0bwE6kkTfdnL+MRCDkFbbppUnEhSNq1y/6XGW3zWfH5
/RMcSewd84/dsk21cxpNnP4qTu2kgEAQPLhUWzKzp+KeKdXt5X+I0nv+Nruw/REJpSvOy4JLVVoj
rCLASdMFBnsZnpxbgjA0NK6jVPPPQ4gpgdKwBd33eVNpS4XuaT3o4bqz9tdSKgz2tyPNPCyz6XTq
8OsZ70Pzp+qpyYcqepHk3ysZAbvKeLcL+2juIO6pGkZK+XrE7fSujYENt88+0f8CqLUN00gbBkN+
4ft6CPS0gRtLaDVYei6g1w2g0DG2teVU8tM8GoRY38ZWqOpwUpE84FwIakwbks8ZBW8jNRuCeD5j
R2+9gIu6rCupCCNd/Vu+oOREHTiSXBf0wTJP7KMzqlngCDORXNkJtu1Pb9SqFfidNDdKumhyLjEg
CWkT1g/R/tmxo3IHsjcsb1pD8sWsIaVju2mkwDzznyu7wRp7vtu7T9pl/aasML1VyyTfU/1RwfEq
fD3CzraegpL6CpOwMOckbUrwpK1pHVwNnvNU1TLk11QzudPbEVkGu7/JAivdsJuBPCuI1yPXabUo
ePnfRo5H9m4FzhZKrqz6sRunW3GXtTiiLIWgUTxBDYGfg3tdCrjrZOYE8u64qWdl5fTNDWgyA9zu
/8iKBV6XHtDorsO9dVkv7193fBufqB60QwD2eS8ccMUh1jyungGfFR/A/Gli9AlXahTROLCGw4MG
4P5zIEXJniJkUvbJ2gG3wDLx+W6deXSvO3n3X7wFa/09DNBFW/Y1ZA7oTZCto6IFBbUBEvIXCig3
jxKMTljhCDES9k3ztIC5Z6Ve3dxdHVn1YrGUjd5Dog/oupsCU916TujdUOHzSzSbDZfogQrJdfAh
OoxwzVrs/ODo1hI1D2lgrpCLbi7nJVCKk3YIHZaVjN2zm6eONM5pTtRhoVWbmLmrMuOTv2sqfZx7
+gh8H7+NLTXir5ZrX+iCEDcblB/g3dmDAa1aBOKy0M4YQZk0HarVjxdSTFa3UxlJDKL9y8ckN/XL
m9QmotIMMhXDXo4hoUulAn2hleJrH5jk5ksBFBOuFjHc72nNa/8AtZfQDbCeTXAFxsVp5e8RV2tS
15KeGf2smp3Q+F4VVw3GU9qEU9HA3B0YQ6ReYgPGZw4q7wScncok4WLmW7z9wn+VOVM7GcUlcAsg
oURo7FrLCdRaAwZl41NtySpAyUb0DYSeTrJs54Wm7iqbtDpwd696/5oFQA25RvSaXfkgxmHTqcjI
npZVSs8or33vXOzCOTB1/JSUXjfHuEOKWZ+QXPkrKgh2P0AI6IOlnzH97DWfmbyCL1mZMAWAbhCR
7L6PubjJSGVfbB/8qCAWuStcQvnhFJSuvWs5NmT+WX+J9IGplO6Ppd9pH+Xat4P3g6wovqrcbW+z
rZsVMhct4dUol9gPQqTrLInLAS3yXYGE5+keUY2l3JI7xVApjt3yS2jqqMgPiSP1M6BH+QzJF04p
wwvXpj2PWJArUz0Z/VD0mxZEptgV6bC5IgFgE66iXKsguFG7EPCIsPb07ahGPH/zMPCLqmu1Sl+f
bNO/vVQNOxXgkrov9zSprVeLVMYzJWbK9HTVMaySYpwLtNFUQFWUKXT+Hgemm/PnSK3chJeCs+P+
cXdIvhg4cGDmCgvuYchz174jsufYkWwUA/ZM6ihaxm2VT+A1chyW96UrwPLEseU9UoETjD8lxtfO
7wOU0tZZuNUa75DfV9O/KdnT2hqqQlQO2FjAW8oMn4gDnFb4RRO9oabwG4CDc4Ys64H1JDmcZUKV
+DobA7S1pgm0wFyfkjXJPPX8tQY/kZzQuJC/5fu38pYr8J5nUwOnkgCyeA842K/kLmjugjvFiZsK
/VVf0/FsWvw2pzoP5xbFZhtLaY+JoIReDkcMc0nCBkaSNoQDgk3PAY8XfZF/7qLqpJNzQ2V+xwoN
PPInvLCQZJogLXo6QXQQVbCzoonbNZ1npHjKm4ryLcTznv/nAZqnGugJd+ws6tWpDY+6NbMrJ+ny
FO/yX6cb30343VtISNU51181nZSeshNrsWlqr8gXTmv2bBnyCAv9SdqpwyfDWWRqZ4Rd/rsZUsI+
PZLYPwb4Nf6J9cejp9vSCC4JhF8NcnWnutpYQlFdY+d5GkqcgvPGvXVfwR6sUEJqxXLl5/TFiRKW
yj1W7HTkLc1PlPuiYQodX4h1NvlQxTsj0fV2gN2czkoWyXNeB6PUeRPgzkKu0N7bSL7ifhww76n1
XH+fJgU2u0VMB2O4bNbvnltRMSqu0sEco8t1/8/eXl1Nml6Z3Z8QEiYRi+NcuUAVBF8sO19VAVJA
aqDwucldV9M7qN508vspIOU6Q5e4tJ4gRQjAl3Oid9Mo6b97e8R60sA/06XWUPb87hQxemvEu/fo
kjkzxuADTOPf+Tz8+1Y5WM+3wWlGrBeOhNJGynqwtltIdh80nvRbKC2/itsE55Sm2xkTEMZfrpgW
XkbaL+D68xdflsu9IjTvpQt5YRF5eEK40niys7W4xwfKK445dYZqJwzBnMO1PYkQtM7BPAclJWXi
MeKEeJ+gDOw6hsH7D4a9Ua1oBxSYbwxQZbUweDWSFA3uWwPmI/lxuw8pXSiT+jI0OTjB7x8rjuyy
87C4vwRqNPpPO0q6m+kG/Nbrc4O/C+FU/xffjK0QF/8gYtzMvy8FYboC0MjmrtB/IaDCOmcKtaiI
yqRQsSCcZ80p9WTOqZ2ncmDpPiOMooiQe82C6JAdlN+oSnEut9mooPT/5x9BA8d+zs7UsKFGNTnK
ASgXAVmJhXHzne0obi/dkBA90yVY4aRKSVkkzpskn05aWj1u+KUsY7WvNlEPzXxSy3OG2Yvm4/EU
MNLdFWUoIo338xbCwDUT7RvlRRQdOA8TglDkvpQ8jbcs8EgXVBEc7riTm8xsdsec/tfSnO7BCFSn
et3Ah7HizKB9odYJA/QVU6dVuv3/HWpw2xep/iKUBI5F5hEFvfp73Q81FGUlODXgM/Ld3MIGnpeo
EtEpCEv6b5NJzIdxMisl+JQ1Nz4atltwyyo5RM9gg5uCq57R9pfSI6iqUN5ZWKr/LZ8fVujWvvsM
mR/5yfqtIzHFljeDSDM9+Gpo5XRDULocG0XGKSqz3/yD8ttXtjXdhGbvEROxMn7Wlg3woeSPnPXR
dYQEh9E/ZcEL87nHaKtEVLFqiZ0DuKxJftWzAHuzEcDHoYWGXDvvHt6B5/y3ms6RjW7J+HaEalj+
ztNz7rLFF0r8g/9DmaVEWcxkPj0QjWhLZtqlnxFUTAzkPnbPjc+1fS4A4xf8ozrWMs10yDYXDmIE
lnlaXfNjhqAvBn7KZA7+CoiHLQgoVFKoCmMdBMUI5GQCTZminX4EJLtOpJ2LEQdXCXTzEHxQdmSR
kxuauf7D/QjgLZUJpiTRD3R7LyghRf23IR335GnvYC2tHBkVsDlJSkDmC3vvgU7AiSFb5SrE3iMX
ptPNOjjHZF97FkEW0DFUSlQPyum/2z07DoLBzjm3pXepDjtuCKxbYvXlSz3v3TSADGn/tJOSn+Yt
ObKv9KgxINnodj3a8ednV/selifniDLuVM0RW8XY0R+NzYzD6eKWyhcrJBh0AnfwAOZ7bDui3kxs
wA/OWGsZuc2VJyh/kWb0ctkXwvg6uNZMheGS3DauarpyQ7jShxnWYYR26+/9flMw0V5mO8rH5GPa
Z82ClZ2LtyFzRvz8avycXmJxq/69WZ5nL+XBtsW1JP3zeQSioyP3HwZGfy/EcCdWTsg4hdY9ATGH
G1zy+NQBRCQ3NIfOooB2r4QyOtsRSnHv1moQ3dTnsWc5IxzZA9fraJ2OFGJxER9LiM7p2/qWQ6pX
/dQVRDlmrlWeowx2gm3vgdI+/mivUPtu1gjrDI9+XBvz6JO6YvHecGcZsRxHdWSsXSsX7P1qgC8p
hSboceCEujrAbmnKjU1+/3UI7fqJ0Yildsty3CFSqAI/mk7hXV5hvaesT9bw/eoEweP+oGaB85P+
xfHhDcQ81OS5PmS0iOBpzjr/Cri8+UPySpWAC2MiaJiXdNkf/z7x6J90borEzWeirXtIkMbS+s2f
/krEznWPUc73auEJgPl7Z2mLm5JWIo/mjlPDPW0WAzfVUiK2zzHrtZGt0D5/8wdy3co/Q0vwMKh9
2QBCgBIXtE/PXS7IjtvviJe0yAs8J4nTJ0vrVuQQPbwtym62sP0jiwTrXEXvbVsMA2LlyNZTh0oL
Sk9u3S+i5DAxR+3/T4aypVq0iKLO8BWTbMkUQjQqXc+qEmJGbRVB3DIxtJ0aI904OLe0bMej4feo
QQ0P5LTvI1e8/bf1qnTMZUIiJHyj1bhzHNs2c4bY5B7ztgphyS8AVNzGun11uyCyDkac3MTZB15W
02MEbrqnN2XrvyL3J8Ux8r/JAyZWCCJAFGBdReM2UTFOSTxa2VOjErXLzigTJv108tXqP15QMFXl
HlCbJy5UCHMfsgDf0LFkeA5f2e4asmRhX5bBPD2zUsKEQ1pO5QN16UPicwh84ZP4+hmU+aZrdF0Q
zCm5ZwDpCpfvhmLZgaaxD4hcjK6ZVlt6eFRwL0R8Z67B8/Ct1zQ5Dy6SS1jwe9aVCo5cy9NtVfQa
nZYmTj5QLRFAGQCk48Gweyec3jjQY0EOFtWsm8yVysc7rMZEt+4Zm6Oa8AfMIbqVZOevz8SngjiA
zj9bbyKUD/SD3B3/6s1bYoFW5YxX+EG8oFYmqcj0XjYU0JS70PpBUloAe361QiNLe0nZxzIYN2QS
BEr3OU5GEGr3i/IFOvu6xIJfkR87ClRhMB015ghbBOqM9UT4QX6Gxmuzkn+AqX2KRVOxu+lrcgog
tvZxDV3p6q25pHw9uF4qhaXFSk3nA3khVKxN2DnCH3U7+At/9+p0CTVuLfPOit/ZeL1QYhwy6sVr
L1sUkbGWMfDXigqcQfZUbsbglOZAU/JHLlUnEJsahLLyOkE/DK4cPmZKab589mLxuqKjdGhYsJZL
I98l2gLeZ2f6zwQKJi8oHF6Cvd/904PHu9iKme6buE7AZXDAzcgwDaWidZFvjI3xT6c3w9tfwmgZ
T3b03vSu1UgEXOkCNx2UHmixcCgIdjPoIXpO6nbK/YdnQ4/bQMc3jWXiNxzR7xswAybPraUmvE4F
pDdPj94MATTqboqEro5Ya13Gtgnj+i91vyuZgcTBWxUag+E+rN+TT+F69LnsDnOB116MSFl+QISU
0pgx86lpeeZmOwxlAf6MYG7Yn8k7PsBpeY61yP7W0zXBa9yTQMskz4XJXx+Pp8j5NOq2G16n+NSy
Bjb3UBJRYo55fVZFCLBVCJVnaZ599gLjVafNDyjy6H0Qxlsnzx85ARM8DTV6tLtaLjwmnPg40D/T
pKXY66ffOzVzGHqQDSh6S5LOVgBeVzCbeQZNeCk3QaS1wC0H/C3C2CfNqKEqDLiK+1MZCpKsrbKm
wKvGulEIcKwTBAkcpjDE34ueYEv0+i7UVIiGcoHXP0SrFcZK5ToUr8PUcwQB3lN2XG762EU+UUWg
mNqhKLrBbdZ5SOMiv5jwuRQlu/PQpAIjG4VdECgPFZ4KbG7XNqdIwbkwjetPXRsct4yTSZv2MUSD
QSNDYZr5ixZSsJKQ9T/ej2lQCuATDUpp1gPtRaPzVKogrP48lmXytsjkeDCcwTEza9i4bcOExdnI
ZGXmlTEbwm0+cb209zr8ncPrZecBJwRfq9AREmcg4NrP7wkuiSg1b0E+DTPFXviGMvsizy5zaEmH
4Zc91rYq1YQU7PWILD1UjfjyzbSPXIvNGNH6KnnQlYVaG7Xv3Ye9GzwRmWkhqmekS9E8UyXjkPss
7FSyDZhDp0S1VOKXbkjx1Jfeo2LuF3lZYLzUKleaJGnc0UUlfdt5sLw0s+wsM+ymPuWsKvn1l7A/
dxc0pnhqt0wDieyqNJnjRf5ncKcWzTVehVpj4efWEBrEvfzL7ny22pwKJqlbRGe9Z1VI62VGq/rg
rXiGIsbuBYyfn1adq53qxFnNDe7LhuwJ8wj/8zP60n9R8hvMc/MPHpavf6uDgiFU/Tr82YNkZXdg
StuffjOdwyI4DLKmLGFfAd839WJewJjAf+zO+/kFzMFYrBsAqbUKFxKyOJl6T/87FFeMjtCsZ8F4
c2fZ4/pPGjdcLROX/FzFNQ0OMeNQZ2vak5C4G5eeIeoSTdsIFuviAO0mikVcUaN25NyeFaaxI3AS
L2jbeAKLt0hphVXIRs+AnZMMLfZhTLp8FesBbeAmFqLhbAzYIt/jhsXpHWlCVHZIGs0WO455UPSp
vQ5QcJl1ZH8R7g+Si3YXc6i1hHl6/SOXDz8D2rpeFB1FBBdeZ4oomf4xFBtNTko0faLzQyWv0Esj
Js1a0FQFoWsNpE2zuHVpZedUhKHe25I+EJIE+YeiFTtd01jZBziqNlDy2hSJOfEZ0HHmFgd0JMpZ
BJPhee2+sRB8gSSXe2Dbi1YhOvL3BNZTQ6ravIp1CVwixIHLfYBX2Wg0ImnXqa+N3AJ5EKEocFBY
pd78xJLhQJmTKT8cY2tueDLHIYVqV5+Vtb5U9VZeOzaTG4d4cbupWJ9oVWO1TEaSF3Eswx4uXHDf
Dv6sP72+0/BHnc0L5KsD/E9N0D4RKxduXuAjJi501IA4IL/CGTg5/myMpH17wi2Tm1GQbW6H9JUN
l/ttB3+P4hYwZ+nd5S2+DfrWqhUHvA3V9F1zc7f2deizuzBdtJXGtTNKwx8zy2BB9zA8dIeNm051
xhtbLxSgBau4YrvQeHodla+j4V8Sl89L8vKzXn+NzXnKkWExINwDnb5hQiiuzztp7qGMNvTdr8Bt
ucjIKMqAmK1dTDQsKvgegiiyXE/RXpzjz+JDcohdaRzNakGOel2Pp6DG2yn7gI2YN3wTbDpOEns7
sikyZILeHmh1AKKvO9LarP3wDLByWt2CPNLOEawtoszgpCiODnq2Oussf5t4nU3fmxRoK9IhwWi+
ZtZ9qb8j2kmaPetLS8j8M6uSwwK+osYETtazsQW6/rEjFabkvcSKCH7MVglCEFD2AAEBO0d0vCQ6
WKzRv8o5u/sumiNDGw4XU45Ng6JTIAbbmNhkTfmsur89nVY0O30xLP4///556gM/KLxdVvkxxbpb
D37MBZY+5wLWc3nM/bl7lEqyKfq/x/TUF8usnOts2JZScmvAXpwzYitzhVZx/qn91i5yED1z1JAu
504YbXGDXjFt7lgaDkVAQTUac6d63waVXjU286SCcNPjzOu/Nyb3TbE7lFyJaWmjZg6yMYRUdDqq
hLYl39QOw3a5OKUwWdfp6McApGmdSDG1HWdSk9avFtBBFgIf5I52wToy90D+kxQMjptfUl2BF+8m
X2WUiXLTSl2Bnz51VV2mTsmt6siOToT0Onr0O1eDTt1je5zJnQDrx8F7AiHpvA1utwu13fm46+WW
0p5M/0TwYk5Yjsh+MuMjg0NVq8fd8KyHm620MU1o6exFZvX/WjMwS/x1NimqMonO8vaDrGkjO/C8
xp0WQaCd2E7u6bfL9SdOObGowAfKT1TKGErseDlFQEidVB06vRx3Jyxia4YK5CbF/bc63OwV8P2H
UAVoBDp0hBFcUWyUQf15toiYqw7xyS7SAWRatCqcD4up0jNb3WLIPa6WgO6jX96GmLA9/s5UXNuN
W4AedMMh8stSfUKRnBvSDHax5qySBic0arLmtd1NHO2iuELMCQ/FKxUqFa+IvBbrIFDfiDsOz2So
ayEeGsPl5biCGs+MW+LhifcFTDKpwFOsOZaFrLk20qmuCSb7lUhKZyvgxJ2EQ09jBmsi9cj4HHgM
KNy5N2cEiFzHqKMPQ4Wjyl1ZHjIYk4n6KInWJcrFqb8CTEduLGNeN8dP8dTDyzbLeR6/ToyZEYcD
hm12OjocamNbd1o8ntSht/o2zG6a92nZqfH1dDyOhoALB/hIxOFaxrdsYE0tl7HkaVxjjXKEVMoU
HJGrzLCaJUOiWCByngxgyWqibteaxmhKphpBCsvmdDtQvDVqjfdAf+t8eh+lhyWYpzLpO2HknfXM
GNdmWb40hB6+tJz+gyIoYZyu4moUreqjCH+mynDrUVcoGOFXee47SqFGoM8guZvS0E+I12tXijXY
XJ6I1ZFC3U4Mrfmzbobf2CfQ1V9YFLoZsj3RWZHUTvzB4RHI9jNuSx5c/feMgVhpRYZzqYeqKGX0
FSp2LQjToyc5pclJnjDOlPWNJHx2pCoexRIrilCuJ/bS5OHzxve3jCKcgWcdchl9AW+dqliklXae
IFo3MD4enFPI/56USoDBqHkbotJLuuOa8E3P56Ecb6N3VOsJdHUrEE/A+jzepKn2kGl8dqP+ozjU
+mtMBp+Qc7iVzEmtpoO4DsENHYiIhqVvNI+S2/1I1DClZd1ECt4JTZ9r4KyRhuZkH7oNRgzagPAI
ubT0TsxLIT5Q5nqdVufgV6prW1rZKNF+g5afN8A2fz74wJXMeiW/p+nZo2dK2MhhDkqNsQHuuuSq
lRYMvIDUP7LsaRjrOM+SOM20wMnCToUKrcID4f7/22MuHRGY9og/4oenLq0pOFFF377/scAr6VMB
RZJ14weTYMaq8J3hffewE5lajt4x5u6lk6fgmnJMpteEYCJNrVkBfgyz74+UDRN6fztxIp/pSU3a
z0Agbp8YkQGcZDkkAXuqxfnGEJ3JK0kz6AWRAw6eKaT3UGnFJVbk7Kg84HWrGbkowAJvQoo5bCFj
B9eILdR28a21PYAvQoMXkk4A3MvwBQwRRMQMWqygo4bur/+zzj42HETMH7yd1Pb18L5qPEJ18QZo
eQtt/2T6Pi+ExHkLVTqihuhYydEcdpM1fZeh8QqvD9GlKYiYJV3gfJn3rgb6w64ne7q4+vcfOjb/
kWDW9pZzhsKKfEZeFpMBI9v+itXjT52Lrax9h9AAsizmxGwoKPUHO+oGisUMx6Pr0m72RrXCZas/
/xrZ7qk+i0JSoH/E+uEV8K0EodQKYoIBI1vf6oChmLW7kiO6UaFQUjCqbwgmFQ+Tk7W2pPJegbh9
HWDhKbNon/AbF5+OaB4t7UUvDH+FzCf+bFJXBLhoudl8eSHJsnQeDBt2GCfARa/lwRg63YKQTKRX
dzTzQcTHYUpNT9RvQC6rbnHpKStijh/cCEmYQZJVVhn+h8OxbI75zyNg/0KQBX+hfPH/1bcQsBTZ
yA4k7DXy2kr6iRUy8/HgHzc1mSyXsFN+H1KBOZaIQuy9K+CFFms+FoBBTu6Nf0PsTAz6aRMdBRjw
w3HamvfA7sK8e189AhWRvUBUrCeH96vfUArS/RkKN7oMjL3QVa95k8Xw4LZwCDVaIsgide42ebFv
jPDPTSMT2pBkZ5vA5SRFQGgx0riGp7LK7IiddY6cZdE6t+EQm1oqW7AH26Ak1zVV8vrKpd5/mIM0
oMAH6uynsR1spFIyEShU1giNRoyX3DXyDMmY6vHFyZzkxipRbWr/+wgwoUvUbYtJJ0Mnabuo3Hlb
iyXH0fMZU9cU7V6sE2yVhY5PRUKMmVULyJ2NpppzgefOoZBWFfMouBlcYKn+8H4jDXyWUMboszx5
dVrBrjiEQzoSaQ15uTD6pjgQH6eoNg0DozCrvRbHUC87XSVCudIXr61yoTCzD+BmHsWOxB1NSpUk
75N/i3VdQOBat+Y5m3eiQt/C1JLAPpPxoUOVShoW1fpgn9nNGiKzg+8qqWvemZts0l2Y6VnblWqH
LGjOtctWRSw+xCs1QwoJV2qkuYL9SP2XpkVbvKj2hkfLnXPjz2Kor6RPuGnGxAHiM0xveFaFElM6
z/SjVk1yp5sCa5NDqq86DVeQL9pcGbt7/cgnI536FEZ62xGjR80TO5TIhrlU+4hSy/YQBKlEf1VY
XY4PTOBFZXTT+9aWK9fx4ofE8Aa84A4HlLLiRXeFoVyQ+lN1POwN17psLLPaG9a3gECdW3MAffwh
yiZcbNg3EvgH/LpIKCWnHK/1Qx5hVlPf4BgXdMjvZX1I+IO/obq7mLY5XtReXF+jXFkekwHMaNKR
bF2OBOeTO6eOOx9guUkFNhZM7ivK8fwEV5KO8BViIFmSQeINHwdJfNmJbOo6i79vUziekL+81uov
Lg3YprKgbmYfYKQZ7YvxFkwADYTC0fHeLQpv04zpm7KSWY4epLD83RiLob+fPfdnyMaKVXmx7VJH
4QH8L/DnEOc0dp/p/gCmFEudfGMu2Ko6ezuZR+d1LtC80YRP96Ynu0q9dlONBpYSafdf3aIJ0/G5
gfo02It2yx68epl2jnuL2NaJoB6gXy1Vq6TPulQ/MR0zcjfdvS7TjEFgzaujgYTjTCdInjguXGyN
3bvg6OU9CFQ7+TM9ybuh0bI61QbswonleGn8jsAGFO6N5UnQgZ1Xhq4GJSa8Wya12Efh9eHVRtMq
TpGiWwRpHs3Ct8ZIp8Ii70uy/2R96qJKimrgdcZgC3iA00/kxmrGgiH/LZbDDyAE2js4WPwMhCyC
KGrhngX9qJVqI3q0mOs1aT3OqRYvWSb31pre1d7GMW7DMRLxzKuky8eSggXkXLrTpZ1P794UA3ls
xB/yZ+V5RJNas5KNB0SI6kleXZveu6plknfSqy2bzxXnh8dUP/FZqa6dWc0GhfwF7NLLE6jfmBqX
IUfjc5Uh4+7kkZCLwazW5bFR4EH87nVGJ+1Vx0QzQpKG0cFKBfxdjtKO5UzOVZs58h0O7j1sPQz9
r4fDjVM3bRLeo1Ol9Z5hZatBRXmSa7R5Gw+RUeIag2lEGw8YUWA2qnDKFM8h9kZrGKnS43/ZN92f
BI4a8Ofc5uB6THLUKywRrGcR3tzsv48XSGN0FFiOJxW92rHQk3aaxsH5QgZzcfF8LG24141dL5+m
6V5n6pIe2I9v5kLwc7tCXTCWTib/X8g2xVQqKl1rGM9vEqNgQdssPBF6g3GVd41IiPRztmo7cp5z
tmS5wn2A4iTn86VKHEwRzFEeVqKZ2J4ZFsm3oEFh/bXM8BrAHnA32aBzENQIWQhh+QWzOXJCBZ7z
rLpESzAYVq2/qdsxER8uMVLSTfGXrQ3rFz4LBfhfYUgf7tJ/MXzNXNpagjSjygWab2FGGs5JF1h/
GzqsQDbhw3FTEOhQ7wgsRuJBNZctzSG5Pma3WRSQ3QRvV6b6JWoscJsffk4t0IUq4UwqdUK/5xsI
Z8dfJMjavhOhwvyTB5PqMi5vT5f3mmgU9Ct8/A8sTdV2Q3AcrSaIygKJAOti/CswduggP8cIDFIr
3ilpBW6txquKHQnGXX8XHJORzeuXuPprmWG5QCWoDEXE8w0xHHeeNqq+QLwRdRvRmRe8oN1KBhrh
ZtiDyNRUrM0gfgQb+qvx29Q1W3cOkWDQfmVvuy2vUHowX4nR1QYgoIPE2KB9pK2fdc+HSm6gObSH
Y5fY1YoZom+J+L8WqQP1I6TQT5X7j9QEVIt3utDdHD33GsUd/Q76b3nylu9+VST+9rMWh3EX0F1D
ENeZQep+iGWKnA5ve6nRvtOZ1+nj7Jy0WwAWiFyTcqc53JSlGiwgUQwa11FaSR/pO9kdrwg4V/W0
UBBIQaQSd74nSPIOAj5z1aNC00Dz/O2MmuDvndincb5ZAxfpt5pUQJs7FjgFKmrN5coVes8MTERB
mFhjiH4Gg4Xi/knPThxkyVs2ZQJq6rLHjKusd3SE4oFIJsOgH7Wr32p94T+fnJTYAf7c4jUHMxd5
KozzJDP7/jxYySyOc05BnjPMqqk4W9kZOSyMgibT70KFY2h0asxleSC9EDsERCp8LxLz34n7AbwC
6trJIGYqNN26LYJcenhcv77Zi/bkmZbSrgwHOpKPAUtRZQifLw+uR3YT7xvAg0w4JgqCmUfjr/HK
gdmNGFRKstLr0ECM+TvzEV1v2NSCJP3oli4TQFafCaR1TqeETSkLhonB0zE5gHgSmkmKDVyX80XS
0EgXVR6BxBhTjuuUpS3iH0qblkpb7+ZM0LAm0DO684WYdhdVrDcKHt9SiTNpYmH4cCo6s8ONz0/0
HMSFcg7bleDFiveJkRTgB4xE09WusM1VVVZnn9CnF5JnixEhqPauWXxRfL55Ax60WP6cptAEXvWL
vy9b05iOVlNu3OYIcXbARt/xStv2167bFMXL5d8yIyxF20JkxWNwLar4H318ULjbaKBWZ1Uh2QFy
ZdyKapeZOeGu17f6KH+5Et9XLSivqeAEQC4/R961g6KPdaX2UxK9NCclizd9shWA/Tq/fTNhxrnM
v/nwslQyPrtZURwZ37KksJQkNvEEH6CWrYQVWVSlfR4ijW6zcAJpCLchj2r0TZKC5HhbqWUj1+gZ
mGcCB1CZz/JzimKv+x5fRpy9jWFTr9gZEZcPVaNIKIzQBnNps7YJGIfJPsujyekmQjoOdt9cXRgF
NyopDgTj6sGN5tQA1/JkiCWApYTlig4uq0ZjUC5XlVEEp3K8FMo1P8/Md0o+GacgaeMRgw61pY0U
i83CmHEi30mJMW0NhRajU9sXUFgrFrrrhDistdDtUdn1iifiXF1ot/5ntIEJTpM/QK6FzVoAOnlV
YHzle2FQFAOBcMU9DUULWMtNDBkKPqOjKtYKSSftxEHGKy0Smu1qn7dgyzDRag4hbiW7++8E9Rff
bDC8aGOt4oe6RTGr5RuCcJcWpVK1rxqIrq0bcDoUuXztv3v6EYJSggdj8E8BtFgN7VF63U7TqYOO
ySEmWcFWx6rrlHJfS6qIDspdhsiDRCR1n/0jmScfRfWNh/yMddtbLmsTIhjYMVSBXBWyKUMV8oRs
nDMPJZ8G7fJwYUxHLCoghK3mxxF0qL49IKOv48EcRpT0Qi7zbPjhJra9O24rinonDK3JewTlIAh+
Z24xGKuIHC0+ygpZMagJqBJqDVyPjn4Vqyx/IaDOuxE9Oi1amW52JcnDeqbBP6M1767CxMN1pngL
saCVffW4/xMWLOvgahy9DDqA2kVhSIxArvWROKgLkElIQlCuzbviVI/Tm31i58tm0LlbdV5tDKm6
lMRg50p9wptqE6aYBukILsAhWMAK66yIY8fKA+2a/mOagu5zvAjeazVWx2KcZfSkoPBoa0ouxhXM
6/fJ8phNpma0H5fi/jolOEI3HZSrg4th6mdioHgWKdZi3hqOuaS+C7rizsnUPwnxMrR+GOLe0HG9
rnjP18zV2782HiojvC2aC/Ftu2zXimcmRVohZTe/XDxEad3kI+sxmSuQ+AdvJrI6ZmPZ65WS/Huj
UcJYEhSegDXumKQNz+Sd18P4z/1XJlhpSWeZvpeyOfh0O9zH5pkcjf/27x8YonDi3S0LLLh92v9P
ee3kMgmMRFbXoaHdOSrDhMl8ze1/IE/JDMcYzZeg+Pn11imlSRf5qdGnbzugyUkVbX4kmMmdDOJD
4wruoRHlxwNfTQHVGJWjkw3j/ShwCFjk5YHmC9iyGPci+9ppSLNfEWZ7xZeiKlYcDowvUdAkxk7m
AqBYPs0ZJfEZzfdoaWF+g4LY3kbKebhm63rQkr5EAzdyYSY7F3loJ5tMJIcM11AIQA82QKsMQTyc
DHGSUhz38FdGUaoG5IJlnoUf4FOr1cgNG+FCiG2+fF5tHzweYs6BZuItmMBW5DgdWd4NbwDOQ4ye
2k34B8y+T+i2vTdsWCJrMRgkm1LnsGX1W/8xDIo/Ym8BhkIblguyYXjokdgaUuhpUhIwTe2N8oqm
DEClsL5QtAZSetywjChHgVfja3T25dsWdL+J2Ye7y9N+1sCHrE1yF4dNp7ICDoZHnzSE6FPv5owe
glbIqC3SxNcXkn6kXDfCdqxY9XXiteubtz3UsejjZ67wM6xaxc+qqDuuPzFksyF2yAaya8w5U1xm
r+wd9h0MA8/tlJCBoYxAimGIjB29iA0V/G8/oysxwwpSuj6sNm78gXtCztNRh6xKCtEGs6Syu6yO
9dx+X5gmsP+7++7AA29c8b557zmBkZ3wKxCjf5JIBoiDFXJnW3drl6rG+j8VOttgmktjLVvLivHz
ieY/BXDxOOz9MP2D1zVGooPJfMsz0+OtCHSDQcZ0GcykVQcHEOl32GRa2VvehIyW6Hv70MOiKCt1
OyqmYfcNBs+CzqBalmGcBwJZSFrWrCbkqI6LfP7283YqB09DrhDoHKewGfUClwodCyy4zWdHzf3Q
kglRnoOhfOxEilCo/UrqKDrX8tVH+IdkZjFxwFwVE3eFPLyE0mty+P3wdP1yMIdrNlWUkk0d7PpL
j+xc8kpVwBgHl7wUaeAJ5EWlW8/c2zUaCZ+0QpD9qYx7XePfHLMbPTVKMJO1H74RVxNxSUS25g8X
8FXSIi5tnfNuCBBCp42Vvy9FCgHyXeMeW1LGnn/aX5VvILsZkRU7i8ymhtDNjdTs7224tUYMVoFy
0ysTF+pE1ZrVV30hLA3cV6ip3fArBDC73fRhbI+spRNtDYZBGBOi8lgNXEgavGMbjv9/KZsd59gc
4Dgz38d/qMb9fGHoORsxhNTJBv78NwE/SzmJDaVN8dJj14RgbL9MxnpWvdZuh915EpclSYOSFHM1
qxNbeZ5dUDxMMZYSJCeSA3ywR5yoJcUNjfzpXgDfq48sBFx1CDUpkGLJHlBBp2r8AV6DT+X3XLaP
bdUysWKe4sbhZFDPgSPWiUYApD/lp3GXUMen0QF0UbBPJbUdwqsTgkm4BMgyb3/nbQUlhAJMFdBQ
IO6T4YBMHL7djgKOqOcOLugCi59ubUTt21ar4ymNYl7gxGGwRVtdxGe8cGYXPfFYmkeQvsxw5cpM
mPDm7IQlPJALSEBS54sG3z2xfIcUiYuq7Zs42k8riFbbSVDQlf6I/W/OCe4vS5oAlqKEcxvINSqI
4MC7OfnzRv2X7UFww2zGpzynbXAM3r4+PuWOE1DSwX0qJGo55FM4mhPO8+XFPIiKkiY+/IgqSEmk
7BQNN+QO2mcWJ/RBxJSn0p3e1BIsDcQ4XVTO4ukt6o4f5J+oiWYHalgthv+0SetuBIUxwRsidcIf
PcjcsZiMToIOtxYZyiUFp4DCVwKCKMPRaPRzRY0X7IDVkHEZ9slWHSvbUfX/ywrL2MG6yvxw4EyV
IVJJBB/2dS9IdgTSi4vXPbRJxoRceWqtD9DkHY724HWVocGICOIDtQ65Gn0knIc4pq8+V1LHIzQD
P2AXAGZGy3+RsIhdM04hvQowyySevQ/R0BB28l3XCy0BEptjquSkMPaJ0zuFYWtvgvVRWB+fAeRb
R7/of73W5koVcwRIum9elv3hjEpy0eg1zf7jFdct18K+K8Zzkd5Rv/Veig3VUhDcHIa9XvKD1Jec
prfnPL3qCEyb/X6Or9Y1eHtmwhZSBhPqrKaOWB5u++XgnDzazc7D4S6vh26p32MOxDwFVzpe2Rqd
Hf2fe2HuVLE2yd73mfinogMViGIewSfMhZNZRbpjGrIPYCvaJvArq0p6p883QEZYCTPXAEFHYUFQ
1dgPdWcuewV4v3YVDGCfOAnniOO6Gn+4CEtqxxb0AiUWsnbITMsE0bYcntzDTEt3YpqNsVLEqfqi
2k98sJWftK5vXXdltmiKqsc7GaT/HSPiBT/3p3Rz61KgJgC4opzgV96vJ86Zcrzrot8RUrz+bNan
8YZO0nZbuYN3NTUfJYEMCQMASlM0p2Kf+PLMWUv++YAiOl6eEj4xJRxTP0s5NB7+9C65J1zjfmUV
y8kwuccKVQ61V5BcBPPkuQr+Md1Djf/IUEI21S7fQzJolmP033S5ouMFPP8yoFVALVOF/nwBvup1
VOyxW0aUoeXtptXjNYZlCcvz0/TwwNzPXrak/QybPLhF57dL3klxFbZGh0/zh3dDXdlBJRco28Ov
54I4Xo9EeXKKIQED3yF9DNKmk6mGLzCdZlZkNplA0eMSR9NTcn3MPn9/YckUKsQZzM5ep4eOuGgD
Lz/FarcyoMaZWVIZIrn6RNjCyPUkApscKGtWizdWJm+3tKgnEL3O7g1G/rz4K9jtiJMpJsWKiMgj
BK4xDHdT8B7jrDuoJbqOmQepd/Se09HRc6Ugmy2blHi2+mVgnFPqbjEXN1PnQbM4ag0f2Yn27s8+
izZspwmarSi38Ggu3YiDX5Sa7MDxZVv5lG7tBHhKymPEPNQU1j4OnkAWoPW7GP4ynKcbBQSKRzxD
Jl5vBJ9poNn1mtsdZCPBH6RhZtMNZI7t2gdJE53sUDdPQP5k8k+aSL8b2hdJJdcEItm5aCAtfO6/
JiW1EQyZIxviMaLkfjpcTEBieLhLjn4w12r839r8YfQ6g3U2flvMOCjW9X4rHOfpiDCKTjrw8mAZ
5wuUvxSydzrw8VhP6d3pFXzsOAmGSApAimN7bpWBRGYPuKrOkQJwVDqCqpuUA0CkT8VRL8fM3fw+
zlo7IZPIZ4DTFCKdB/HV/h5zQ2ynFWbwVOh1/WzYpXhT/2GulOi3aZnlnVXl//dkVdKRPZBNcZZh
WlGzEM2XiUokyYQU9Oc0AHFylvfev/jAlqUuBPid1NQWw/IRWXPd/5l/85gTY6pB94b1eZJbQMMK
Xi8UotgMUwsV1F1TuWK3RaLL21dFJbfogmh2thwD8XoYGCu0G4jM3OF4gmSXJYklZdP7TMlM0Xwb
auXrd1m3SQdI3zwOyOBCRqOneOFybUILnb/ydanWfMNtmfohg3sVy2Obd4pwcI7T1fFC7xEDyeXA
lJMCVqE0jXGBHsuNK3ztjUxm+Pksc6rn6tPNyCA2qRhbtij4iCO3Ji2aKMoMRL3D7tUv9Mx2xwhu
YtHPPXllgb7XyqYdOHV2tL3zOq4EeVjVQycvT1NLt1DEU283QTJ4SGGLe6cAAZLQjhS2DqRkDbfq
M1XXCH08H8O56I/S2pBRXL73zDV49MMFO2HoPlWNFDwqPTeuiq0RyZkHAKT0i8h1FU9FkPpElrGw
Rq32wLg9/iO764kteuYPwzUCU9WclsFWxMnFnWffMHNaZBKrefqoVSrM3XTSKH6eWKE0dJ+hDphW
pgzI21TR5o+p+WJxAthB860vKD7YJQbkjA9OLwgsXta76MewbozRmOcqnOXAAPJQsIhWApB9tk+l
PDHwYoUevNcB69MjR/2pkPl0K5NwhsUoHfRDn+6mCdAz7W/hmFJDbSoeTf1+TsxMfkT2CJSOhvZz
vb12gtZeEv4puQwvrY9hvncLq1Tqev/oCbrZChCWtoOKQikp8tFByTAQhaROFkTfnavEZpR0092K
t/Anal7obPn8rOFpZqY/CcGo/Ht3B8RWVmIqxonaC7ad53JceQftanlMiqf4r3u78FXBsgTsS3go
jCCLbK9IHEArpd3iFbzPxsZ5L6BrpFiu+8bDijxl22Lrnl6L473JhGspIhXyYsb5R3G7tIt5UyPr
TRDbvqZA0gY1/umkL0TBjD6oJO1yOCHk3LjvO4hRO/TwmbMrAzYXz3WN9wWS8n4yqLlw0euci849
51iGkAdcjGkXN3nyq7dcd/mZI2fg7H3iFNRRSV425U9Dz/P8OgpWuYvJJaM0NguS2htQZwrTVAqG
tL5sKByshbmupVCoF75j35l5BjmTmosoEZO4AP0R3cBIcgBg7QEnL2TGL/JiopA6Kqx553rwVZJR
bExQOk/rpVfNdVQZgdP+9lBv+1yC91O0BjLvUHMpbPgFIe8mRImTLDrjmBlA31IdTl2tOGA1Waw8
1AxcYIa+uojRmHMggGw8ohHPYBJqSVSSQSWZAjJT45SYQBebGMj2f+14S/HxpkUowHZmc9UgaGry
J1w68wL9j1Psom4JvVMwtxIPBoVKLhOlFWmjGZM4Xo2+BfqhW0J7S90ALjB6cbRuVr28yBXIfxce
K2wuEcZk0XyZy0SAzClhMOvVMurZzutIIfrX3jD9VeYsM584Iv8sa2TDcT7qcvt5rA3QolTk8snH
qxPwCPuk9bHKlDi6vjB4R5eIELX/IzEFJYfixrFWierYwhvy/6mECCbaBqIi5NGKneB4lwzo5n0S
jak2c/9uyYV5M/Wtil/sqn797FNgsqjCi+SFxXGFcn8avPrMYsHors/AgprMpKgnFovbs45BOpvi
0RC/iaJ3FuFKpiFXqnybfxC6OnNR+UQck5x+vhbM0qDWFnVJUgL96J8bq3eU5E4vmy7U0dNvVWZx
4H+LnKW72dXASLNS1yHIbMK1HjXohznlR7F9WmvkrHN/xHmPDuzWjtc2dnLA7S+iL1ZRf0l0ge3i
Vc/vvxfJGQLYKB/na7GP/ue8byQJxKB3T9sWPcxomwj11WeB7lshHm4kDOiIyPkHu34MXOGRYpDB
u7GHWVOqIbFtmnmQw+EOXtpSKTcEIWpb0/Zdv/vq2XcBDqGnJt38N6f0LdoUquXqG+p0K3Yff9DV
C+5ycOay1Wj6pLj83MhC9Ef8RGxFQF8sEsEADwlp7CKOc7Y9yZ63DDSeRx5YpRlLUOnwfcrSw0BJ
EEQk8/yrf7NFwK6UhogOvV/oyW5zuub1P8aMZuWc7HkD7MC/rEd7B3KCL4XE0sWEa8k96Y83XOnM
ruCbY1M3UmJgAZ0D48kOUnD5Rgfr5pxKwY9TlJjrZawtf+PRAFCjbzZj6WsIwqqjfmAZEhQjLgeS
yMclhB0wK3NEYk0JJB+Oa1bS7D9UK5tjzA9PLRCQ8ZBAlohNkmvcrSA2OslYhJpjooEeIwnsMiyF
GluMnKSRqgl7o2peaIJce7/COpwcSOpEREbXwEnikhNl3XHm5/VDqFmlIhi09Dglr6mMfrb4v07E
vwVkzdTxVFdYuQjQBKAhTSfFI7wVDoJV1YASGeLaT0cdQr7f4jAHR858SrwSUHYELy4xFHg0gBK1
mM0X+qRw6APmNC0m80eBEc3b0f2dppMgzibdOk7CBE+T+8m0L51pwxwBN1hhiPD4gpsVMbWxATdM
cSDdYKA5WTVsd5429rJOqIUwkN2/dz0kuWHeCg19B+a16d2SYgZsEGg3nua/15+l9P/6I0lsUyqq
/7hDuo+TFwLYPKxsZwJSxYv3KKtfM8R5KQO0VnxzqlGUnxbb4KjFTCGrbMnl0279iRWQ9CTScquk
QSdns6greZFKlyAw2O0FTmcAWP+NK5OqtAYPW205TdDYK0/6ge8D74yoJm8aLE/uo6xAVD0RXiyI
YTJ8OoLY7mvtFT8WApmy2at0YESGKAP672W5wkx4EIK5np6TLBWajZS9YjUGqaONXuAFLU/UoSR7
XUVTOiKFaE/oSv5yE48XseqsGTVNrFwD8fNz2gEiPDd7n5pu9AHtaezMq6zmKfKgttZBV7XZz77M
yjNiiS6/U0TH5IUst6lC97OjH3UKnIsjGXshFfNC3UzZUF1BJ//6J8/2UEIa0V6EzRN/uxAnpFJK
OvARX4kVdaGAqjNytECVhySs51Hf73iQClP6PhJ4VZwp8RnvDYuqA+emP7iobmloWPqrDmwcXXXd
Lyqli38b6Ouf1L6jjybtKfCyn++3djEgcvROQ3aVxcVRE/WwTQ7ytE9ManSQhA5f68IeId0UvbUD
asyNRzPF+kx4YnWb4126Mi2A64oZCh+e70X0fX8XajmT9HGzNzzEMYl0uguRAgpUYGSi81mKA+UP
jrehifho7EYuJWCjGtcUuLbjfRBl8Do6GIVeWbtlRcMzAHm9LJYGdoeKxwlLOeheyQJdztrYSxYn
FmnxI3zvGxBx4mmnmmq3c3ZY8/s6Mxugk8+Z5USZD0ePqgxsBBAl8d/U3i3XMVmBEW5te7neOZFQ
W/xnUyqQ1Xxk/dZe+u6V/FrwJci0czLFYZcQ+2+DIM6IQhkCFgKEyoxAW1ZbHVAIGxov4BfCanih
jjwrjgsi4vyyO9aaR8Fm1z2qtRUimCzd8tdNQlOxizmteudBQYAz7qxtVn7Y11lUAqzd/at3eNOV
sWI+TfhRhQo9W/UEGJMyiwMvmai29CQFdDY/jI8cniEzMrNbgvd7Ipxwi4oNSKXxV6gLhUU0TbSz
Vdm2coIg/m4CcfUMmK4tm1pSidH6ccJpMwJpqFz8yxSsrLcKAt00qj3f8jyM6+IjGadGiWy2DJwG
mvk9NTw3jHVDS2ERskBwTAv5j66AuL03pEMDb7cdKjymOldkxkw5LN9AFso/EreOREErYhkWSQbx
hIy4QXbJ5zEtSsAPi/3zPr1Z76+eaZEpzjs7Kmfc7PzkZLWh7eD4fBZgsI3VQ1s2tyuJTmoc4+KA
i9GXc9KbuhUC8w7kSSoW/jW17/KbyQcIq46qji/9OaCN/guEXWXv0h4TW+VE+yt36EnMQR6H8xnZ
jjNI3ypga8w6DPa+k2b1BJWRhmu/ROag5//1SSKoncvFUc3Gsgd5WgTBa7b/yMOuEBRJR1oW9jlM
jVFyZmGTqFOrZC5VcHhvNsugYxsvjnk3nRqUvfXp6+Aa2m6e6HbO+mHEbdXMLEmwhZXCC3Gykdh3
wth34YpSJO1Sf9QLeS2scaZweDP+YxV/v4l3Xag0l8KQCaxZcPyjvfVfuYRVrvfAKdYR0u7GviSq
7YXU3nAA4uHkSly6aLFj3tv3RuapDVezK0Ux4Z1LvjjKxEnqS+fNl/CeygGR991jmaX8Jv7yQZLy
xFfPR78bDKCk1fGCGWFDBwb7cCRiEmf6i2+bJPA6p8kTH6u6iB4kRZpAuXYeFe86jFjAFg1cBdMU
kpim7Tm7tDaCuSTqzuA68/e6dsV254pxfCfz3TQsoLgcjAJv/b/JW6x7ghKR1Zown1wl3vAisY95
3UxUcHXtD08cJG7rqrwb50vaW1P4FjwwrWTN0LUXt03CDvo7BhKFHs+FZum8GPXAOfP5McJ9kI8f
daLqn2MEOXSiXAxHjxZ6jCrwBlXGRPQ8CKarDGJbH37Qyyz6kbYREJ8GVp1G9mxCapglSN8MKiTN
os61L+uXspuQUAP4IZNlDn1BrBSLNseFXjyM2ZXPVZVpwdonfskEUEFYZWVd5DYgyuYJZnaNAEI3
qH8jAAnH0sjy6PkqbeUShIweIhlTYvjAayXqLbUB3qmc5P0lNX205NXLukSg8KvMl6WbKIPaLT7a
71Tp+2yThjjpmtRTQp166Sr4WK6hP6HUpPmf4A8rfavKo1+Vl7lL+JRflDkCmwEPAS/j+6vNwq00
Rs5fkeCH1j+Su3Rfg350jOVZYc125s2aEHOtjZXrtvPvXCYStUaNQ9mda+W+HRZ5Alk5AxrtDvxQ
KCpOEKNIR6bbUEs/TEmPfgOFXN4jcItvYBXcKVIBABZw9t7Gcm0EXX1JWNcadUGEovD0pSS2XSBO
vLzfeehYnBChrnTQF1Fr9FI1VkXrzTVAxfby+JODbnxOZZbpv8X4UiBPjoLjnozhA5dE1mcxCe/S
NHkXqM3W0Ul/GfRvldGHziNeDQSRAUaqjQGCZhIVhb35zoGBkq2aqw2eSHyH6X4bdjl2+d/dxWnQ
NeR7s3yfbS/PS7o3m8WuCwm0x4ZA3mQH0NzubAZpSDATjimWFe77B2v9r5QfIM8yG5Rmx9Zaj8XK
JtZq45blHZCFwbBmVgqgnMf35jErmMndlGFlQhJvGod+CACUMnGiIb981p5jxx6TY40WujeissBV
Lyusp24mZG6OI2grc1ucA4Q3xs1oqWPF/Ljciry52JFsD4zmF+KG+xFsY2nHtaBaEchMMI8HLMen
Hgt/I7OchclZhiyMqWK8KSVOADbv6jibTKxHRga6Z4wKXmpPd1GOLjpvOqXAzgCqpuTu5PdjABh4
9cZUc8sMBUp0oXcY5mPeVFbj//6g6R3ThAHSrdimLd4XuQ/SXwyu26/WE5FFddVjKFW/MnuTxFP3
JabrQgPZD8bUL0oG8fteKFt+gcEXxwaCpDL+ULU/UFg44LPUT16wtIoL90H1lBq7zv3NB+VpsZ8U
yISbx+ov//tHczWunyzdnL/uxQm3O8vOWI6SpmDHivNwowcClkORa8PaDLgUs4d6xdTN0cYsAHv7
SNXigzIps+6NcgSPGlx+ICsFQkwWxwiCamuMNr03OfTKAdQ9aooSg8idx0kSOFBWwvrok6M+wOJc
QzqV6mkghOC6sGRYIw6NGb/9J8rKjO4YrPExBM9Pu1whHZ9R6c4q+uC9j9GNDrSosnsL+tAVJd45
kIuBwFPAv9qOipoyhWXk95OmXbRUuKYmy7ZljnCKvxNskpDvn7J5cgINAJ8mTkqQpSJ8u+YfL24b
CcKSXUpwgriRxQlwtxcuosCEMUHQRxvKU3aTcj2NfxtXkLCd37+qTX2O6Dwm/D7hVRHl5Rnv1lhh
rUXKaUcWnuBn8eMsghLwIu5VxAlwTLoaItxIdaEqR96ah0Tk3KQq2BfO4GaF9BXZZzqWmAovXi7c
cAo58pqdJ2tNfyTbS4v6UQx8Bd5gbV9nVksUiLCSsQ8lWleXJsSXj9foHC5D8ELaiOx9VeKYGDiU
xF91ammtCClz9Ng+D14bXNNhP3QKoYjlBt7ZxkAvlg14nbhn/7Fy5XMRIl1O5pXpM9znutDOL8ro
l3HrQV8YHbM5iAP27mZFlxLIee3KpdUk3y5chpmKZuZrkpE1R3kER1NHHttklB+zHJen2HBWES3w
XXd8+wv703DlvilxGMU2olPEIKcxvD3/UYxVfaNqD4m5mxKi37Kn5tAVx6eXgk7Jwp/HPDxbXDrM
YefmYcePelc8gMd71lbCulztBpoXG1sxgYp5LvKKPdzuOvBXJhl14T0Z2fL3tcn3Mg/bCg+QHc6p
uszDJOQs5udpsux6jyOlyc3RAVqpGGyAecPxfuzf4jFTv1lpy1s/sJHpu3FCZIqrM1fvXWyE6yGS
trfi1R+MFr0UMNvfn0Ped3CVzpqalIvsMOwIGALPAadxnsheSyXaMG4c9gO6j5ClAYevUNRMYo+k
9n/U/TgZphvBLMyF3RTW6AJOnndTCgGucPsDOdnYUfeIaKvs1YIHLVieVfV6b31SGcMgTAs+EXVv
Wn3HCCnPy+07dvq6hYUZ2yOnX0TDqfTgAzKXb2zrwpEQhiozzaOGz1LB9SIBASUD1K9z7HvLDjXg
gqV5tz5i9HSs7L4HuAPKPojE8MTbXw1AxZ5eqe+QDytnKU7KuI7sY0//bU/QkZHPcJ8WaKnne3BE
aZ3ePFRrvlNpa7nIN6PA2l3LlJnzof/2C9IXsKCCjJELSw6O1HaEb3Gz32NK66e+74dQv/66y6LU
fJiPcYD/UnlljNO+OwJLF9O16yy9rmI1qKkTi58os+Kt/D5FKAC+6kyjM1a6YfFtbrK6wADXCurx
nSYqGc6DVB9AzQvcC/S8m/IZqrQeMt0i6DLvyQTyErYt2mFJE3MSW934LYDu4VEMKJ9DKlHFjCty
VjVCv6g8FsJYguQk9SVVLXAhn8YngDG7irf3YVRFji69BEKi8qPvR26xjKP+2E1Ypw9v2pSIc93t
zkxYHbyq9SnPL4ORiVNKbmHZRXYVK9TZQT3xy7qcyjTUn7cepiPqvPqeqFOa9WykrKdBv/tGhj6h
dmgt7HnmjRYKwrMlLp8d3gcWtiTybTgeAC8eIDGTfPn1Mc1B9ELmKbCdfxZfLT+kuKObC5FQYq4z
Zk2XmYy845hgNd6Eica5N7i6fbllhC3o3okOhp0VHmmE2wdrYsv9aPQB4n70vnUQsBIdiRo/VOxe
astWcInwYVgVtO2/D32jgUPuUs2BMVBVdTk7eKFnLRqMBRYJlmoOEbmyeB8Y/j2cXcB1qUQdPc+e
xm/6gMmJ684cjMu9sktmoVODxh7a6pEG4/BhgHkAImw3nHRoBP1jMZE3PuvSfr0SltCVB6jLpENz
Z6q9eQfzF32UnUf5GLPWzk0j7aZzzjU5WFgzCCraG1IS6d41/JZ3k9MEW9Hcrq74L1vg//fzs/a2
GeybcqgrBc6+bLnw7au5Bq6Hc/j0HoaB6pC3gSVamF2HtDrOEOYGw018iB0QD8ne6C9b+RKEktBd
x37b5X4zX5wNQjkF3h2+eAKI9qF+l448i5se2YJQvLljjTicIJjgLQzkNKObf/CDTga24T9s1+1K
DP3VYe3HQ5uIMFbNHdLRL31WFIiTWo5BrG0XnSVWesL9d78YuED1MFr23OT1aXVXmAvAgnjS09Pl
gI8MkA+OvvhTR89z2TiJUPjPh9I8++4CvVdZdFVXMrII2/lu1h8r50Q/DeDUwUoLr6jGQrgHGvRv
nmKxGcAzAD9BWZhtE+hxHY1eEmFNITsOeASrpBatTLdm9FTdCvs5dFuH8OA6zAPWnATxxcQarQ0A
mwV8Q/LVX9BKcyXb+R8oL9zpcWppA3IT4Fwk/tGY/cAi4mUCuSGkjIxuE6nYzGm9gA+bFssP7aYK
890jrEQ0ItpdbGq5ovHqZAKg/ZejA2pMiSXc9IIp06znLpZ8YUMExTweXj18RIDMKfIS1DYMnv7u
+vZzAEPWYDDKm7Oj1bx3WNsAq5yXC854oBuel3FfLmFaVwPdSpG5sJUkrAqouocFxNk9mh0iNpaU
vO4UW5SrevbzggjMJ3usSMf3jWk8limqLmWOnmrOgITdmmVl3vFiAVgkgCpKKr8yRovFOVIofvqF
hVLXRXIQjXajMrBpJF3f5Gxrju2CTi7fdmjdYx1Ph5YeFX/HWh++IDkUZY83UlasZqEHTZt72Lz2
xZ0fa6INysLD+gkTo7fnPAOJhJHsy0TUzxXTKVpuQ+6liuMLu57N5IEWiytXpyhoaBLp64HhFgHG
NgDEX3u1QzNkJsxReww+acHjgB13XpI4I1K9+TT547UscLmizA+C4oJaDwDgvC0YFl/jNhT6Mdxo
1n095FDt335iMwaLuW5ZWakdisr4Ledm6gTiahqAeZq1OEZ0g63dA5VNPv8DJuiP9hFD/4xoSxXd
d2GMNZV0sAAVDR632WVYJUGVjEQaJmcdDVx6WlxR5wp8sUx8jc2OiNq8NfqOsGKRUK2LN4BKtPyH
nQJNo4WOdykqY+RmohsvqTARb2LndhwQYivtZ3K8wQD0/Ygv6C94bnKC8tMJmKm6dzg06PYZFsJ+
uGHOf75BV6Dkx0bODg4SYyyLz7RgMh831Lqf6r4joCWERD8YhbpHFKMfoBvoVxhDeS9+GPR/YEtV
qYaARoJembNJAbBguhdbW83dazarzO7OxDpgc5B+jqUHPD+GqqaZXN3C9TwqgtenVnJh1/uq9z9Q
eFN5uDI6WECpPM3ptOALeYwvZLEkyh/Dw6uN8mFtJ/AbGfqsntB9pbxzBsvhmucITYFSvv/11EGC
EBN6MSJqbLsve94HWYiNdp/DNkjzAMt9Yhb1Hy6ncTP/YOuxCGiQeDYyX1Xrkf3gk7ixBgrznojl
5h/ZP6VRyZqU8/1E1XrOPKMY2oqOJ1Gx8Nl70/vzcDG5YSEGtmCHdpW6BfxysVsnPhnKka/5nHSQ
YdKxRYdGJJroglsHhOPIv2nXX/FwaT+0XficVOkh0P9z4Ru5qVgUAjXBCpjpdPUEsHUKBHFoQIS/
h7rtDKxzjN0WwrIiO+WHgZtzlUTDNh55M3v9uVj5+h2Q1v49drJJMqEGYmBNrowqEPULtlKuT4NC
rXhVHISCD4ApUabGxmvLnhfVub5Yzn9m50UcvLmC9cLULFW9ttEGcLWq4d6UEr3nHq+1Bo7Y9LLg
CF/c1tNkY9ef1QpEKW65gysKhwAfViIK8/qjRrWylGaH29SdT7HWf6Oq/4SiYvN6ddtAFP1hBbWz
57uPUFpOOhpuS6jvKjl0mkPGW4QlYPrwzGWZefDbo21R61zwAGIoxTVFJMO5HDp3hRokYcYpU4T1
bSdATT12teaY95XFkbLF3I02ggjpNAVtLYyP9hiAHT/kw61lR2Sdve/bE01kwU6Cwg7FRkREzovk
QWQ2xOcqVo/JOKwsLDrnVbkF5Kkq3fMXz2y8VzmrtqAKhvERzcltA0qScJm46TlEGwLFncSsZLfL
bpte9P0KZSSHuBkcBnhXlI4rQUIiTuu2oQ47fFmduYDtPLgwVlL6Eich7bikW1RgT4CNgaVqDpia
CzhDkJUcmjDo/0xHo5Fu3RZWq+cv2OG71HTD1NMEOEecJckWJ8fKi5nq4dUZ0pJJHhwpPL/dMmon
LNXL1RaRNmRAJGjUQNH8cNURV8Xi5wrxI9++aoMBuw81ex/psoIgp59ZQzhxZ1g80DPYhKOTiHgM
Rr6OGrh1EplvTk5kpDvr2wxDcEvBQfCtVmG6nahZs3uRcoFEKYbRaAApCapgMC6nl+8a1JAM5VrX
l2uwgMQ8YkAatkS4tSgs27DXGVoWuXVmiLQmuXrlRqgLr3dTRRyCLcvvQNndEYXr5+9e1kR1jCNy
4JVtAfeA5yc9PT+5bEsfMBs2SfP1pF70R+/RfOl6aermgWdrcyBwmxArjeKMiTEapYGNqNsObhU6
GqgeosQeUDycfA7VSLWvhalkGIbNIlTXaTTiyikZQa/n2KpksJ6sNiLm7iUXWTw/6l8Lyjf6P5HT
qkCvN6xNwJmgrCQHxYqmUtk71P+FKpq68eVWYn05MIc+6svklBP9n1XvNtG6NhEaEGqfxYLGeJ7Q
Ax88NolXgvNsF37UhsR4EuiHHYMtcweoi4IKPDye3ffEY5DwSx6esnyfsmZH08ZKSeumstIffTZH
NO9zIAXV9Wy++xgTybnnV/zXcB/lcQksxCq5zelxtaRU+jdPtyhNefhoV01/eP7S7OeJHIdmG+zM
WIOQnNNnprhmBvFR7eF6Lnf+QgQW1mivSn/dsl4VkQ0ytyNkJc9AzixU5EJsmY85wKrgdxSBt1/N
l7D75ch7lvLk3S4/VsGPAej1HZL7JBa04dekE6xUdS2mqDHBdsyEKv9nWL0oLhdHMqX6XmhxnzQ+
TvcPBsOS+4q69Yu9Zm1m8DC4624yQ2kRCF45gAtFUImGGoET3zkLLLqzPYB/HC+9vazICc+Qv9oy
/il8F6YhaIXxSkZ1TfXQqfjewf/S4zLd5itwOz0dZ0TQiCH1sGIS4EBsnM6jsvbZ1nOJtqoo5SQE
pI2YThJ4HHkb/PUOX+yxxzYgRl/cVXoE69hI8NgWZ9e2nkmVr0xY+JH2aC5CmR7uKyAjROdtJrVP
necv29sYeIFNMJt7vnjkh55G9KFbeOm6IAuw7iOn1QdeTtsXs8unCDs8QddgsKO+KxF476kBKz11
ZHAIO2LxpCAYZsSfXyfpm2hRHE7FD0uIAaJoJi2NSR+AjlD5NXCtLu1xWA+KcfEcZvg73+U1lcDT
FBfpRBNklAQdpvRT/mIh8pQb9PYFJK64HA55MZx+UxKC+XftRc6hpam7xl3gvuB8us8To/aDU3ED
y+50fR27/ZtGFgN8Yjju2TqCq5LPVE7Vp9JwKKstGsB2br0gPhN+QBElypwR/5N58vnW21fePBdH
1d99HLH6SNICs5rU85yrv8q8CXzXlXD0tyE8N7EXCDvsIcb2g8Xu/wui73KAgpj/K9QUVLHRnMR+
2xDt7t6KWt4DJE3IxaJaxP6bUD/JhurLf/MCu3gh7Uot1gfXrYP2GIZn2csx8166/Gxp7mNDGCcS
LqV9sqaOFznd06uqLI1h9XdMSIOn9GWqej4gAoZOVdmhjOh+PJoyMP2qrY3AG1jjtPBBs5Cb8Qrm
ftSYms+eejpQNCbvW/krb1JgxRUga91N9b1qGSR0o74BiDJt7Br10NDPrAsT93b7yAxk94k2wc0/
W3Rzjsmp0cTIjjwPHOFlaEy/nGcQiCzppw85VVbxZcGgbSNY29tTCwCOLodpJyax4gfKoj/wAK0l
HlYS7DzDB0NonIpAIb2QLv9q24SDhejFr7gIRw//KKCYPQETp0PuxpPrOJt9OnBAjjJOwR8a0pFK
CejflhCDgG0hGyaiCLigWrxH90J7OY9sWkGTVouJxXNvVq9MeGul1j2WMbL7B/qYaNs+YYRlTE5Q
zR8qRy7WLQYQ95niTZtAto5fmB0vVey4rcvKHvzL4XjbFicUWSlxMI9tW+a/RaMvF0Z3WjYixyPy
FFv66y5ytTN6rt3AWFZ/yMt8b3g3TNYLjoqpm+AaE8IU96QUyPTq1NWFgdr10CIFkl8Xnmxbmn70
/Ir+61SS/8rLaYfJi5oj0SoSAY+457KzQt2FCeC6IlAK0SVme5cHuaS3NR09iO2ARlAJuXtZjmmw
bYir6n9lfh2zkEsWdH/8K48BxD3KGBOQHCttc2N9fdIenxxVdZ/TzTmMRE+aXNv3bK1e+Dj5Ukxx
0h6aKlp0JcyRrhphqdIzm5p7Lfhpxcu5aJCAeHDIbfy87gx1y3KOQYBkZ28GqTzqzZjtnXxk55M7
rFXnpEaXfwwyo1u87EynoIZ4MQA4GuuvNxy4i5jad+UwCboAqFJtsLDQm3Jm9LSsnSEUHJ7geKrj
El0/v6l0wVmHXzuL2DjDk+ivryyPNb71C4k/ki4cuAkyzdvW4YZB2Ym+QDpX2f1fZMiEhS7Wn24K
8fi+4Jljv4LbRxI1aAchVMnEd9EWYBNsepCTJIKCo8bbaTBB7GuBnGDXkXsi4wFmB1xLXXxtutys
axfolzFKYOLfi9EiUiM/Uq/03TJ2n/YrhGU259DbNRD6OBCzRosUtXIfRSeUzvpJt21YXuHOB51P
qTEJhhuRIwxOOrH7MpGRNPMUnl4QLcBeATF6o7UPRPNeyBOv76TBXSn+z/bbw3hXqYE6c7akdlgV
rz2PzUXeGkGLvkexvYmUcAG6VS3RB2AMC1PiVS0Lkv4eohUF/ZA+qpMKWTDFbtlzIexXCWesq9XV
nwm/Fz7/Dw6a9h/W1nROIYc3rN4ISzAGpydWu8u6EClVTebC+LKGyKiCj9YXq3Zc7xDZLpFUfaT7
9+teMLbHpao9laNL+Ch88QeaSsD80kJ9ljJqgW/NmSVQ4AiTaRoCaRuA8SJx4+VzTjr8o6Bpby2H
XwbTPUdCQQ2fusdOOGeFFMWR3yRt9OoTabso/1IgVvVSFyeIvEFRJLEu5wTNiDeXQs6IgU+tGaaN
+4LLIl3Ud/OTFMPKrzFoTCOhjPuHJeTucauj7YadcPbMoBe6pmEhfbgNMHuxsA8EHBzF7pLULVmh
Ng3b3ymuu6viVUV17fmsYKpH830MJsdKrJB9+Vkd4+JDlSP/xMLPR1zLB+fMse2tQkSDTRN4//VF
H9yiXJCocPDfwdM6TEGLgy+awRbXjtAD2Vo7lf2tFz4G5xKDLgx6geH91WWnYuhbR2Z5JGdc6cy2
Di9S7eLo0w1LYY5N7IOI/L07ulkhUS+hC/Hl08l+PNCO8tFq7/1mEdVPESX7S/f3L55wYie7bK6I
P2xVpiJHrzDPBSDfe1ysrAwS+zGm+WDAYbeB1f41gKOkvpfzIdSUpFvIvdj3ZdBQFhK+hqs+3CvC
0VcaQmb1UrZt2GsHL8Jf/Z9zGsjOITJJvh89P2V8LlcyeK9cNOD3HOyauNWpgF7ZBbSVpvw0cKkK
ib2MWUMbBnFR1sRKXrDSIGXzjZLWmD4Ozlfx390pssHOaQElUxr1IvqKYoeZfACe8Z7Y/lrptzMf
8onYtBRTVGqKTxRm6vUM4+JeSyFaWXhL3J/v3tjrXhcxr1UOXnT8bGU1hHxT3pcL4H+mH8ufJjCu
IqgTBxpf4YoWtOBUffWCr6S49CtwYuMKGxR6sxS5F3EdkRVB9TCPvdC3/zVqI2h40dKhQxRmdfEV
VISQahW9+rhJQaBe/na1dP4HZQZzQrNvEsGbIHbXCkTJ2azcuWtpdLEZdqWGwql+SDERVIOse1JA
qgks2peYYmY8q/POtJpui31VlRnARjwBhaJ0fA0sdqXuL+DHHgABWqMxAGD4h1ptkOtj7Ut/3/7k
mBU35KMpCNUN3Lr2M/wFNS8v5xeW4PQgI3PvqomR3QNFD0S3xJ0K7w2HJLO/EnUHNRw/XYW0FuKA
36Ju9H7sI7+6sihFmZWdKwS4kGxTY+M5gY4LUXzTfcClZZlRZVDOhO9QxXzGhfM3/5lg8h5E50mA
AkLaPdlQCd1i5fMD1MQl1rbqNbZyFptzJSWSzVxB4oRy0ze662WYOXH3yl0NiKzpIStxlJw3Qu54
PYZ/b3xQ24QnSXUAdp/YwhTfwPPgiDFS5kaHjJvSojQTapRO9Ss3PJy9eUDIzG2QlIubzAkXvYM0
oH97wR+hDMLoctHnwUIRIw89cRJFDl9dzEVueciuVXhXunixtZo2ulKSMwksaAEWDGF6l48Rw46a
iKaW+RTnqQLOzqPR0OdEkjm1ctmn0dUYrrpzF1M5LnnWkINLSbA/9ecFP7pAW+lpbeWgB7Xisbpb
0v7ALJbFy382EbQ0uROJJQuMj7cl67OIzaGsL7eJi8e2RpdgTvNYqWtLJD2ALATUaSjGM+M463h/
V4fEZB9Yiqk6X/1sfMh6LorMR1L8u2kWFFaBSnNCVap2PxcqllRIEK5k02tBqg+uk5Yuec0M4P6S
Rl31NbYZFHilAnga6mcUw5RcItUdQz9Hn7aML3W8dZmvHZOGqyu7+6n3AQ/Mm1iTRBdq5nSMvIq6
zDiZ6vwctRCA2LceA3UdzNs+KS9pFakQMx0dIRGm37QCEOZ69gUxWsQMHWz8YGC+7IwFhWEQWVRq
gd8ZMI4QbIQCWNW3ZcSiuIi4j3DE1eODbPtYKm0CXXbMheWQbRt8qTwNHvlgV2s9ZDvljobpb1OI
OJhM/sqyynyoQVosHOIdnRe1v4YEEuBOqI87sxvxDCZJ0o2IyosH8OOjR99oA3xZzHPZXDJt4phv
F2dpdFDIisOta5yj7s7pk3KhVNY6B5vp/TkmR2VipQCUOPEw+9rLKbpGR3HeWd3HR0jIAxlMWKvQ
2XTaVsWslpvp5nP9TV9MwNEJZFd/DEt7v+j3eo9UvQUymwcTZYBnAT7KbmSNo8AgDlDY2Ql5TvRx
C88M0sWnn3Ejacr536BqjctRxfiPxNwYng4ocCR1wue2WOPvWsTD3lw02p6+QVMVxQyglAayN5ju
xSG/6THgZaAX0uLNINhb3gB0V1xPZl9FHgOTdLMWqX8hClXj6Cp8s2CAYLIR7wR2JsFhcTP8Y2ku
UnSnVBSoKwJMEGFwN5poAwe68PJU01g6AQ7l+E3fXqAA6YyrtIc3MXeRjcJki88YQretT6ZXg/SO
oRi1nNTiDsgs3Dv53mL/SvKvbDnHL024OsgsUKj/GRY5op/SHbRaUd2RHrbGjIsxJpyg0N6n9zpR
Yfd94FiNARRyv/RJUg6fu363aABxbcyNQfdjbTSwVXiis1clKpfvTCLkAnD8SyEs0QNAqddND5rp
EJjat6+pQy+vB1ef9zIbNS3pINdKrsgOvoz9IX05NdwfaH7fb11B+X54JMKfVN12WHURSrEl5ypn
v8pk2hWGs73UGEr6q0bjOcfnQ6CJYY04HQ+WDD96XqOL99TH4u/jkRpBswzlkHGLJKZ5M4nmInEV
ZVT3lV6KZjXHSYMjY3a21dWGGPD6tp7f2Ro1pmYLXD+hUy42kEGYj/+DGDCFhX0etnoQiX89butw
ikVbjPjIv5YWlOaPu96naLTRpd1/2KU0En5QxRIRIts6oEcmwWwM0wSkrQiqG15LfCyQl5Hs/psR
kLsOYhf/ZrDC0Iqdq/QMA8NTpI8siR1mZFj73gS4LpQOOHqVN0rxrbh4HtmDdP8cymc5yc2XgQfy
SyJfNShmqzUIw3QTrcIF4JVHUgsbm4wrUwIST6l1BrBblokUnM5HCCZ3s/8d2s5myiBgRTC1UWR0
mny2ufUSX0VMsFxHySHO9NoT9MXsTXalLJfUrpavvFEI4LpOww3+yKr5Fs3MmFn9foeQXRukwpAz
rrRmC05A+e2BW7ZGNQNqNi1wNKsW5+AwV84imk+f26tZPnaEad+NImeM+lKhHn0Fr1hPU7zBgxiP
KlmQR8kWl1gnL+FY6tQ4PyeHxZpjvPK0XMvawcEi1ABNGUTQLgP08V5Mboyd8lhBlSDhZNSEHS9O
Xbz6g8mgWJsAHEXdPWg4tJx06RSrSpV5KoWbjFyjF6E+IfC1M1LspLWho97i6IJ3KGFM0/ocmfoD
nZO9LuzQ44xZZY9LpPftdjYuigirSC2Oh8YOTVdhmhEOcI6yw5u9ngohoZ+ewOVsndQdm4rdWV5M
3vIJAatUO/SbJTiWth4VM4lZEuYNWaS0clAKfY2ilmIUo74YjWax0DM4yOX70h/g9hDrtQZDzW5O
ksy+uU5m7/75EZzti2kgcr41hmVztbptX/bOKN2G9e22m9wqEQD9Dh9fRpIGcnCshUAhGh7UROec
NJO1WV0pe3c2mofLko8+T9cgvT1a4NodXy0YbPD3Y/ifMhg4A8Cl+4nPQRcwW0t6gklpuCPYLzWF
XwnmV3aZsseqsGitnLfyk5ztRfIuW02S5qOTprR4puMM4s5WiiU+sP7+8QBiIZ/vKsxZwZNnmvUC
onqWR/lw41f5c0VSXs+QZdbgHi0TfFVNZe5k35iIrta5DY5fPjljpPiOnyytmyYSVceRahrnN5ou
b7I+4izdI2H2xK5p7mE8rvP6IrjCtWWDJ1k9ObHbcXgfP2rQpzobCShp69lZOJFyXviK9zhPtVi0
gaZirEgDiyvDjO+ZksPyNWKoEb7PzRR2KyOaeUPILN691fK+jgpMW6GCseSOHq4xdMVSrpOTkgTe
MZ43oTWXxXRHTokq9JI6/Xp/m4Rg6HpMGbNrnlkuxfUsSAlNEzuGVdF7l4zO5m8Q2hvbvh+Faosa
J/06/uCj7ly+Y0U1/UDArRRuwcOOJWD151i+tya707517sgwEQh0IdDYBjraBMv4quCUw0VBMv7q
etbtm39iVMVK8Khk7wQdct8DbqzwfX/LNpv/02yNcD6W3FTIobqE+TL5hl0Y3J6JcKp19Az3JaK2
h9N6pm0tZ85rECY92axhsypCpwC+nzAAjrffZbAl8sw/6Mo8w5mtJBD3UEYRbRUyhLQILmhnPqXn
vjEH0NAHj2DSsWg0JlnjeqeTFnWlwbh15QoLXKMfcoH8kj7pLMgU5Np6chbsITsEcGMU/82VHzOD
Arff9WRzsEle2MlvF3V5aCgQhANWwymM8dqvwn3eqiULM7p2dcb+NxYpu6lvc1NwI4Lk1yDuf4N0
3dp5kTuJyWaST4UKJR3OskK8mJTvMZNGrEuoYR0vqzru/sjoMUDg1VA0m+UsjkE9oWjCizwR0jTM
6jcH73vpMKZ5+6awYgGCTQKoiifjvHj2sQrB5abbfzK8jMvoK/UQtK9EUaQZ52wxyZqWyFkCuXw2
3OF6bdjVeaCMTjVDrEs9XC9MRxL0Aj03axeMJ2lE4rKWoHkVVZm/n388OKMrqAEAbb1y+VmSiltQ
Hvr3geRNjMFg++QEboKreVBiyVMFBPMCKXNjF7t8XOjpoVBAtllSMly3hgWR7OmEjAIRbtioJmW7
uWFPfBVPF7JzLCuSK+u0Ciptg3uijl1nfILpKmj+4vWxtc0tqWZ2iCrfaVa8DPstMit8DEPUZwpg
Px0zSCKXTM+TDb1j+2ZXIsfqJKoahSWHBGdoBl2y5hR4p79euRDPcUGMwkFn08iaPRY/9VyXC412
HkEMOKk/SLY2JQA/zxUksb4vT2AW4SluixivjrGEGJGgn1RQzbKhEDSBuY+k7IhmOf/pmD0lb73N
w/jXs7ioFkrTLgzrnaIv/y20b7XgA9dHEsz6eyQpMgwRjVsvQc1yh3w61lkyaMgFgh1fnm5kUbxf
EwqJSp6s3aIDqforp7+tAfx/4+AIz2nfLwueyHPnYKGKmv5ZO4FycSfY5iYI4zX/2ifgiYAZqEMI
JkcJ2ZgFoYIUSCKrV1WQhXKtiTiufztux3zJ8IaRuTB/s5kPhahz5kan1jiPdAuCjLuLo3jh/mSn
tONy0/QDUh2y/Vb0mjiOv7hjcMq23xT6qsI4JMrUejfoWr3G8jzh8gFpdK7W3PTFTxAY+ic8yRbc
cH08kql40tKWi6L3tj5OikpS2JWQYpnYfPy9gI+2N22m2G1DSUeIDrYQRB49RBZWR4tuznD38l4Q
x3Ja/+HYfyyBr7+ZI5ZkHgibZZ7WHbNNqc6lhbiS2DiHxwPU7w0b9G7vc3DlG6QaiclbWq4Iqz9f
ZWbqvjnUKOzKjnewnaxrc6vP0uBPBqukSFZAbYayNSTdTZBJUz6KFOuaf21epxU4OVjIbZmJyuLh
p4TZjJmmYHgFU16kIRf/GutrYhQyW25jFGB0OHX6bEcVhX11KUxM43umde/6ZWil69GvsXJvGcu0
vDEIXl0igQsEv8YKqZJiHKZv+aUSdjpDmp7/Tz51Ks9TDtibee8ehdxsm9YxdieThC3OPbu9QcUe
QLkjZt50YsTQQn3P8xa5fXFqHzIOZN7k6EMUzICtG8nj++BPQDKWQUCtWmwwzpa3sq+DlubebbKI
7UnISpq2r6OeUR4r4aWMCArdtHHwJ/W5fPig8jeZsvdVuHAGA30Rwbbu0d56PFPGba++LB1MKS1k
eaPVyNKO4680CtYTZoucXMN1MCrTcJ+Bb5HgGeurUppTaZ5MSx3gxYA0HCFk6W4NRdUi7OwNTE7o
Sk3E4g/V7GX3BD3INfu5vAAAz/HQ90WBOL5TIfuel6bxlQanNpmmRJ+pgSNzAlLJWDbH4qmlV/sa
LHh1ARODxTAWPJJ/L69/zaYbdklgHNRAhvil5BWzIAUVMKEMGCUq5jJTU4uaNL7r3cEVq1tQ1rcF
AWmt18NMnaZ6yxLMY1fwbWjBZaizBHM/Ebkv5m5JFVqw0Qt+bDx0ncoaFDSvbuyt7ia/7fAFIdIy
ueooSJ6VYFML/JMvaB2/n1Mi8ScLUKHC/ksKQd4z0YER+BDUrt27+dmx2oVeCvDRV4Y9HZ6OdV5/
QBOAMMNoW+buWWWAsHVnZAUFICKr8tXHcTFJVNkC9cGM0lW6+nKvJVBXlnqcuS8i9X7rvcFxkMOH
WujS3NIA6+abJIIZwr7pUpgyM5BXXrf+BDLemUYeexQ3zvaevfC6rRG4JK0OWE+TcwisxE5cPKr/
CowlJCIOZBzUd0Yi9PSL8L7pmOhyqSFe9uRaOTgb1ko5hM3HFDwZSlEijv1jjF5SsMZ5G0C9lGbW
NI9VWtt+CJ4qUQGbbIDx+X55B4FydJ9BbyTSoKMHfLPvlTjqxuV5PmN9P2Jy8MKV0UKQXL9XzajT
pnkguHseiIZdN6Hh/P8/3SlPWyiHQWV0Mt1S+ckskWJzU28YmqHGMSoOHjuY9zLekOycpaMm8S7D
dh4NmFQonY22UindiqFIpzPxZjx8q+7YU4qD6m+bFSp4kFQoYuTkYCNCosPPfJInBukC30UagQen
G+DAZuSrdMhGIfsbIqrOYxqlOh0pz1LG17k2PfmafT2GULrMG7lpnZ7Y93sxoCiQqzreU5YhKch0
cxHttK2E19UdTrAohYRBegVjPU95TjkAArg1y5FwJbNAMrS57bhExTfpj2OaTSIlXxkHqx50Tl0B
2H8FJF9iAbPt2I4Spd2abQ/RurWOfNBaaCIwua94fzRejzB5VJ0sW4yg9mPqj9fBYfFNcyYdvkM3
NChZ1bAWhTCDpAXv4OQpuiajvIdaEgfi7qrKJoSk4kqVJYjGFOqQ073DtMcQcy66bUjvVny43OLz
AYtTQUl7tFcd33skTuk/cNevl1kgvN0G/2Z7c0WmIu9tSemZ2AxRvby5DunZmkqV6E5sTN7YWXNo
FfvuMijwGyOwasyZswMcvIeJlflZ1LuodIZWri3ykVWAjsxRbfhqlKFe3ZuDGj7WZJeglFSzxfrt
GFlfj/U9K/lK7yYnZoTGAq86fqnCjsCbFOKXWGNTirDe1yxAT2VDAPHfVJfTQoyTA4hVlAitC+f9
aRAp7DOk8rIZuyZPrWub6WARncEvSy90WfnIVenS8m5L2mChGkCCW9QYtp2EJNw08Q5qjPKhDnmi
ISuOpRYm8+Bw/hQg833aQ1QezMe4HjZc04GJHGifT3W9ePVG1TmvOgSO/swdbH7vK8GXCObyjGd6
q9WWtdKer8POXYtJfH2pLg8nfiR2blUsIwvd2n6u+IFCmNwhYR1nsSK/hucxe+djErR23yjw2S96
m20wnP5tn8w1Z5ropc1CQgwP7BBTQJ5D096o9rTHpXo3go1bdQo8FNBTSRzcpCytAx18vjHvd+fD
ICM0S5c2QLRG1Amzrbvd4qnJI6mmYr1EQ9BXrv8a+u9GxrtsKDsTJToz5dn6BHZfTMcQDmVX6KDj
ZL8HvWWhG73anTrwLwt4ATTED8ilG5+uPS/K5pe39IGyMwYsGyJkyqXU61KzXvX61K8dwqtn9QaI
FZT8JRcvKspc8GJLqREkn6wJ09LlYp+ml5soRwesAvnwNFxaeK++p1bgxedUipHwkzX6qubz8Iif
nSCiltvVNNSxY++BKvpMIfQJsNlDmhLakNIyZMojffayp1EkIRSUpScwkLGs0ZNkXYtWYJIui/8b
QH5zgXJYkG8gAYzs5zfl7nRJWruyxLEloTjSRKb0lYh5qHzCi2tcIo5f29E5ZbB+92TAO35UlGJz
lRxKqkedV4/YJKEH8vDnEfLLxVuuFCysJlkebsbZaBk3FDgIdnxMdNiCN9nIyZ06wBRyiQcfMyz6
YwdxLjESYFyCOTX2lZ22vu6IOMz/w+yuNfNn47RZETM4fAm8+G3bejvzcX7NQ9zrfh0iYiymfaTF
yeGIRIgn6GK6tAFGRncQvXNkOuvUVujf7zSPNI+XSsQPL6FqpBfSn3dPjyIz7bcKbCfmS9qUIX9Q
1p+eakxoANMsjfIIELORVUOVquG2x5joOdJD9CTv4bNLvYRKwZ/luAIHEWPQ6Qsy/1llHFAO2hj5
lIDqSuI69oeW6Haz9JwQj4WzRsdwiF7oU9TtGke3SGATb7ahCLfYWcr7e1kQbkyY9AsGV+NLj0sy
cEQaSoTCxqzDNDy+ArEnu0QkEc4q0OO/BYe9x7QQARHP8ounA16BpGQ8tSuPfiZSILHgIbwX7jNv
5MoHtsn0Id8P/ii3g+VM40l6BVu+7feEYFxP8JaQqfOmFW7hZ0QFOzeyRQbDb7KcDWoO2QiBxKJP
Lb5UNZYIyr+Adom1VHM41LhIWiqVk4MZdCkvFwUXCYV/xlKV3MNz9hDvGX0MYzmDeBNs59U87Eip
qovjevYQ3qCmYWbkAvmH+Jqwh2aW5xc2+j6h+MfGwEq0NOcAHndIN6r4+SqHnv57fWZp8+wo1lzO
Kj37pdXXHOcSCthh/b25gEv5EdoFe5zgFTnZRvHLnyNvKaZusucFTPklQ0wLhq5dI90ZKifBrBTV
zqi9Ic3ye39nbaC5gw0QxXULTU0zh8LtJWuYqR4M67/ufWBExjp7mf+S5+V0K1A437v+dD01sZU9
s8MnUD5eOqrMFgxg6EkAF4QgmKTJNOf6q53TvSE6rBkpnOBbCLgkX3dKglQSV+P5xT8JZ0XrWWsK
fT4LUDpVZp2oWINKT6cJ6eNbyX6e0LLUrnxXe4aom3509X0//eYGgde2VDqLO2k7/gIqcoXlQSSP
QtoxRnGAyjbxIfAIhRy+TZ/P+LT+kOZ09oDtzju533yV3hjE7Tg1Bt4GnfuQj7p9kMg31VsQyfgf
nNJG56bCb0vhAKHSRFA940wI2KP9V3hyiIA9ooZU+/IXfORLdBTFUCjmmIyeAnM/fLWkJc1yQW9z
x60KLbQtpQyerSuNUWz9x5OYTb/PvOm7vhLLJqdO52cggoAn00PIeEsFs2RdoQizpsGPiGKZWPRP
960MCf50JDyjPzumqnxQXTThuEQkJGzVYzRqpidjNCqWq0HnO5o+IliArqpACHSV/Fc2jN6vBupo
lSHPwZNUvc9gpdB3gL/RojlZMzGzFagYO38VApks/nHPtfQNFB5nsclQJnZe2Rc0D0icTqMX8K7n
cswqwgfDAUYd4LI35O1lj2JeC3ij5aw0BTzMOhpnEx+AVzzIWDN3anVSVQGQ+etnplPH4HAR6OQS
3espQThdtox+CEks8rjBBaZJbbKtKZXYSnEYJQnNedDCw5Df9suwi17UHkTKJZ3Kk67NHDv47cz9
r1DGJb+ySbVn2N/kG22XSr4Uwu55DOPBU2VEpdU8n4bpflx0kakMYCPFHyhgVLl3HOxXwXwL86UP
7U3izw946xg5eRXgSTa7qEuVK1pczEePyOg0mRzciEWvsq3w09Cg7tiBIQDrDdXlXD7T+AZi3jLu
lGXXz+/Dhpq1tK9GYyRFvHKviVRKurrN76443SDQLGMtRVIV+C7w3Pzt/zqHTcTLwZdm5LUEo87d
Qf8qwjXey7lu+8RleCEXhTw8AdoqvgxHAU2z9e+AaPkIAoTxgXyLmnD0tsg5ixfGQhH2rJNM1prT
2JdXruR/wVIe3hxV2CGQPT9MEVCWJrRy4LfGSmHiEpTLQfioTYrJ42CLFcWYw+PPFi8x1VvTyDkL
CNQwNR2MV7qR5Hunwuk5Kek5bCMKnFmLqWGs4HlMrG5ZLfwJkV/Dx9Xq4C8COteJkU/oTBtfPVSi
bWP4YLJ4IdSV1THi5PB6CKGQtILk7Z/Cf2iSwK8Wiw501C4Gzhv9mcnlaDHvF2Y9Nr6HsKubkiUd
CneRzYeDYinfXwHandUBRO6eswq2tokvDyi9S1KBPcRQv3cjwcBLHFlJ/kXw059YzfcGMMXvg2Z1
DJl294eNUghgSJe60VcZ0M3GjOT89QTIe40KnsgAAUAHeIYX+tTKP5RZFg/E7L9K4dg3/z2H58g9
nYOuFCQBTEVsF0WV8gYSBUrUhHpIPCSxtIj9cWE5AcfM9GISwOUIyw6rzywWfUE1JbUlRo75pKVT
FWifm4ZYctN0X6wGk5VBSx27rZlmWKc+Mz4IHr4Y1nSHGyTYi0pBbdMp4dx1EubH4AGqrXlEPE3c
oiapKDWwXNK7SW6f3OyqjOSCoNANAunAagID2Ed1ZbYl4PO1/VjeYWSkjjQzcsMQ+gqyUbuKBSNi
Mgvont7euvAXNQavmwyJSE7fQe45C9Hkf64korEWFaRRlePgQDpQ9sL0eyyIz0wJRfOdIZBwhMXk
F1ZIzAhcMMVNukX7TTQ6GESdH3YQewTAlFwtxmNPWsCBWGTAymJvldLQR82TQcFJdiS+3dQVS0NW
Gn3B80xC/dCn8HNrHgDtetxh2D/l5J7rEq2QoOivTudZrrZktvAimQ9UA87yx0z7ajwhPA4G6Klv
zaYLIxlJjQuEdMQTtgWau0vJgvtVcKVhRz6Y6cBnToX1u/8+g74zp3KZduegfCWe5Dfgrq1Iokiu
YBYqdSF2veySPSMrU9D+BiftrmSrNxghJZFIEgqUsr2apVYb0zkueocqOLZg1oP6bSsrjir4i9xE
/z5mILVcUjh5UAT14rx8pNcgByIcAGBPT4zxiwjslskXoy23BgppTylUfM3YqRSNw+EgyCWWLnez
YYvUw4kW7z8oMl5+qoR6hlXIILtzzKJZbfkSC9EdCj6l87nng0V/yUR2ODMRhpfvz91RMSAjxqaF
hFsMkgWsKaGkpU7+Zj+CcX6RTD+cxzeMrlza/PNVp8bKHaYTlg79veI1dyj8FhNYLn/Z4KGCizgC
Np2b65m7e6r9i+B9+t8EK7l4v03jhXd4Z68DzzRweBNKGFnRCS8HiLG9aaMgECiPKU9nFrmq3kl/
Yh9RHFqBWeWEXnWn9sihRjThST0V3jHV5KCXz8TcatzwgT7yKgKVNzrtAqRU5OChH8omD/qHCoNl
Tqn4soW3knKTIeDO1pN3ne/R3j3MA4rLn7lHXP0D/Z1yEE63LMMhV28w28YdOc6oITnaauxvmhlF
+dPo8DQaNRkQ7hWXyTND2WkTWuDRMMYD1ZaKVVk2x0BZ67UNUJWyMU87xtjkGaTqQiTieV9NIRC+
a9h71bzHk8i+/Z+yh3ZSvU3Bla3o1h1pjI6IIJhJn6PmbjsV19A2HjeVpAKGHyoBGgITzDBLzPJA
bv7KewRouw9z7P9t1AlSmHFqGgnQOPdlgq8aN6DLZBLdEB8B182rJfLm5linzsr0xqC9zidMIHku
oPevpn8boWs1iiRhuITlSCEq/otHkRA438/cFdi1/AewEbLNh3ACHRM/zoMrMa33jnhasAaqoz8q
zaC2rpPIvf59IYSW09rv9WJ9MwMcYZ9l+n7RGQ6MbKGnPraYHLk3kOPixEntbAPXKCQtoFMvfBFP
uAKuGT7y96utnL2wgsNPZ9qBxu7Xn1lyJtbnBxiatcEj2ZmOsv0gwUXYHOvkkZzEhPMH+mSeY816
Q6rwnf+rva6UN2I0JUHzpRtArAzSYn22MlApPXfqK0FReNhrMoaLp3+oHbJ40WE8OTbF1A7FJ09y
qlJebWZ6BvJFiK/VUYlXjatB0MEbnB/+oRhotVWDu5gIw+ClRfMVbghDcifuJPMwn0xz335Mtzx1
JjJxHr21Q+RJDmnxOv0AXE/A6lq4nxKPhY9NEFNMjsAD0oW8ehyIPvbucciQKNvLaUUEULqO6YBZ
GaObEJPg9vSA/12LVYqWzLY4Nr03tym/Wm1rV7madUVg7IdxkNcOkABt7egqzE4F8vpNvyn5lNnw
t9eXE1NmfNuqYRvJxYE7qwx44keTSretpIM8rdfOLmejREYG42wh1P8IxOEMFcjnMMF5KAyo6EvW
k/VC3fLlX+nwITAxkII8aZxxKZSsR12GDrfxnTOsYWJdeFy8XdlETY9tJvXJRuiwC4e6Q312In3B
5uBqfpYxkn8KCatWJ+Wcw2wFiv3s6EAJRnfF8DKhcoIdgNNcQ+Ukur8OZsKjJMdcYsPSxiGOAnxS
S/iZFrDCI1mjQJXww+zb9dMMmVN5A7ScN7fkCIVTgtDuAaydwIEaZcWGZ/plMsZ8byRLSh5Ds867
54nO7LchVxhiGSTYwaum0ZS8cO/DlYkY+mgJ3EYayJFfRy8nw7gHMLg7afXH6VUG9z+X4CJxHy7G
2PaQ/+3sd6VgPWZxhDQJZcsa0YJBC9GOOxLmRC2htaFijjStUeX9XVMFTKsEVWB+t1xlFWx4ZXIE
k7Ux3cXR8KyvvmYlr7wK/BQ+jvlr/rXnAzRvDqsojh9j3uUnf6fAp5cO/w6tHo0Nn5uvLDRaK53s
XnKTxeSHNqvtXssFTImgBEBSPi/+GYq6aGUBtW7NmY3P0m0tL+4QnXP4KxFV4glWOhLA5KsCgk+C
CiQyc20ibvb5T4KkG3pWwddJvB9NnUc9x6YVAlZM/QLs2Uh2pjJ2JbFh86M0mVySpaOYZHW91FM1
bCKa2fHrybnZ7AzqIAEk9KIlsCcg33Lxj+9MeX5+KbjvR7GU5mtij1zFljXgj89M1eK+Pm8ep4y3
0e4QvjndtITSeBKKunuGIBJGKUwwCVv6eUlIqPkwdkSvJGrhcU8npeuJO/2wGZMdvmCo+gnMzMvK
46EFnGHdfW2xv33Rc+orjyiRFF8ZTG/EhLNkJHXnUP+/R7sSFwfd38ChQbiC0fIXkTlZP42v51xv
4BOKfK3/3p40l5uEc6FyZZAAQdRP+JQvaC4nxNrmg8zmCZ4AriWvX6N+0c0PsMAyWiylDI8P0un/
7xCjobg+t1MdfIFrZGnc3oMSreFRqlMx5s8JUOXjurwDKAdxTqL5eOqEC+qy5v2AS35wQwzDhSpK
0V6gOl8YOPusBUpIFA4f2pZRZ4H212Ux9c9ZTMFD5RR8kVLvxjK4GR1+o8vUXi9Ky9UxAhlmLCOi
/H4nTsyijrScnUwmmYElyx4mHrEBQlVVPNWtd9dRG3tXbqyAY7zrTgEYSvORz6pMlX18F75zPZhk
LVJ5t7N4F2dbOIsEihWm8hEJPKhT8vhc/3g+C8QHaw7meV+7dWpNV6Z1J1ind6DuX+hgW3xfeDqc
rTphFwIn8oIEzNl5QVHWL71ATc/DwzWaI7e0En2fvbQNMESYIxs3rCA1zRTBwfmRie65QgP0epjR
iCuTOwuJkPcUFv+mSwAmUv5VJQ88WFaPNtxNYRI7ere5nbVxiKcXDI0fcIT/qHtEhcZwO6N39zlE
QKnSQQ7qYaTSRqBtdc7qFuTgieKzEMGap7OWIw/180uEjnr0y0KNg7ez8HTF0TZtYtkRi6QfCCwk
yxO9JOjwDIsXKXZt97jB38dZ3vCsgol3Vb8FHl2VLf6V5gN9DaIQgZTAVJm5eFihAGRNw/vPsasH
JMtJeIv6WGKl4UxEkbQ+v+lF4LhJc/lNveL+qijNGq2YO53WUbH/sNPbUltegk1RXBGf3ACNTyFG
DrFiAHeD63meElVUBslbNSGHE18tHmMlHiRFJYSBKGCR7tI9Y3eOcZHWewXZ1HWMa4tQl8bUIpnP
CSUclrz8dpWpcs6P5ddifgkDDiiBOLtHj9tU85eGucAGzZ+Ck0Ii0c27vUwNr8AKnM6sHAsSEayA
d0iV74vHlYoPdnAEih2x3+VmH2/hCmrnrl1OAXhJallofwDiI4W1+geXEtL3S+/OqkhKU4D46EvK
UarZNO7IrCNWMM/cs+2ZjrgAeBpjx90LCE5Vosb9DM9AteAKY3T9KL5ok6q4+J1xnGKvBI76T8A9
aPJx/rg515sLPm8QSxIJzMkTrfU2dYTEKmxRL2LzFM7pEgzsXbR+D1IFsv83OE+gerG8YGCuKSIB
jl8ldBodDH6pfo+e2vtdvHtImRO42MRxUU88pagogh5eb/ubtNOPZBPn/6ZIrIboDbpqVfhYQxb/
ojuCreJI7Az1w4qNbhLFgCml+ns66k29OOAH+qr+ETkz2L+hNoIBn+qPYA4CvrXgh2baODOhtFTK
K1KodZlfOz6e2pdsEV2GmpC2Cbd+nL9122RIK13ZTBBVjp6SZnt/WKILZ/gWuiDL1R8aMTA3x85Z
e3kzKBX6p5P87n9FbCef4KT3bHs9L4FIBqp8ahDKRmKga64BK46wvRbc0lEJ8IzQbDbIbCu3Ze5w
splRIFh08qBur3hnhDrsDXiNT1xANNlv3eStNTyJK7qvBZxzymYMlxkBnPHJIvfLcZ7B3JhedFH0
CsSyec4MYYdRzER5g4monljciTieuaAUDTJmUNmCXTdpISg0WiyEtnO7jkWlLFmgXFNfGy+Wi3IF
B6Reks/SqdzoCximf+A0emM/MIXxtZqrHQoNG3v3BdEuTSBXP1UQ2g2CpRXWRvKbKTiUYqWQH8XZ
WqarOp+VREstWLbgF2zHU1koiLLDlVFQepjxljLCLmPEuhW/v28lFJ0tYYdyxycUvHQQvxkxAUXE
u8pypKH4pp41MVZu9vjPCPeVqiR5c3BHARhrQmi2k9wjP0bzWws/u21Uw8WPyNq8cz8Pab/F1DQ+
uSz5E/F+6d5sl/reKocorle/CYTu1XvYqaWX9CLL7OLBorwTdAD+LKBIc1QO8qZ5drZcPzUvsdvK
TZt6brdcQq7dOrzXnwSHgeVdLR9+Ug6tDimsEge5+ktR3j06i8EdZ2HStgGQncMlAUwc/GCj0EZ8
PWTP8qpDwtlMgfXZz9/hH5zFuygpRTlWHJ9+KpGUj8eIK5290uKKnKSyoxWUjuNxBkvDCUys3IoU
xWL/nq/9BBRwLzO7C+pBDokazLM8ku21HcvqEY/dWuEhNn0URJEpQk0/W0btGNOuHR6OP9RpbmcE
Mnjq8ipEYhxkURyYpMJibaATnFguw7QUU33W+K0vC9hn9NTUqDRXmraF5gyLiunQQJWLEq/Nei/T
YAylqi++t/YO81P4FVF4Db/x8QGQueXGshZHZzjfG6n7GfCGPl6FM1KkG57U9euUni7TVoxzJ6IC
cAYM9YQzFFjKDbi+zNFom14ONCmgVxtiE8HVsKIbcNwOj0+Ep6SAKLo+afIfeGxk7u36CDBnUe5I
G+kqqgDvjdp4AU27zPOpm/T0R1xOe8KqCkC1m/9zzVcrzAVPLxU4ba+zqe9sXbBIbrCyp03V0XQs
nfXMpSID/EByGKapP3ltn7HNq6QccPAUZf8YAD+5OFO9zYEGcgiq0SwUo4Z+r95jMlHz7BLo43nV
Vm8q1bINJyKuSCmn+yPSmkVIXfh55Yt0ioL+yFcdTz+faeFf9xlfuV2z9HUXkW/q9gwAzZfiwi6L
8W2b+PDw15vtTgImI4QGgRlYOIc0MWORobOXp8AKHez9cqqDUIpNfeDYt503Rr+w2ZiHcvUqGE3a
p49Ka/uOMXzgaNK7b00/Z61brAoGg2zfETvRawXqO6p6JjL4FvEA3oMvPBIWsCizS6yAC9a3m0Uc
h/VgKoeBD/oTCvwWvLJrEsrw0N1d/rYzS2eOdt5ut1R4irEEbZ8rL8wWwgHCoJXdS2XJuzGg5d60
H+QB4QC+t1/Ed/DwkNezt9JH4ANylBVBxZM/CVIjWFSsNq1+OWlJ04rcRS5PjWXQMkux+0TYIr0r
si6nNij5gq/hJQEQJkS23zWWqiI0fkLLBJ8ZcqafxagIAd2y1bTU4qiKVZ8Gvv55zBkTrBERQUkt
tXoCNrEEuFINvDkrI8ApugjWgYKIBDG7GHYFdDUVbSqUIC1coa+4zCjP49YJQWKqt0D2JZbhjTtg
xkIoaaRpnaur019R/LLLHG7a/o1wij0NXzXiiywoZv4Q1kPgyLGpQVYHlG4lP75t1+uuJJs7cvN1
v3hbo8lk3VxnQadlUuT8PsC5f6Q92YqKgTkUhL2fJYww3vsAiGXUz/ErkRSZJB/wbnT89HRaOAJz
0tIjkjCDDoxNkE4SD/kohsHgV147OGYL2hS5A835ACWqyVzOnjh4yhD3zNQfH/vdFNcjSUHfz0XU
Tn+L95+pCgeJ8h7eS7tbCRGu6XM9lGrBbSvhjnN1ArBDYMzE7zyspcHieINVqUhJiTfJKhuS2s5b
8hOOXr8wA9TqvVADJ2mR7mVQsOEQs5Qu9dtaHuZVTb1HC48eosXqwE8PMF8/IAU/BHpSvDHnare+
9y/MhmmxEp+EqBkHfAKxgRpaWOwm5xS662G3ruCgj56vgK18KBeh4jMvJUOcJKBNh7OoI4dK3Gx2
PLL0tlMjuTCWaGK2KHLX/k9lwptle6jn7jeo4BFM0jLyIX2eSWwSWdNW0X32wNsHDp0p6e4m2nmQ
5EIDDVS1UM6wLdrl6+EDVcAILTxe52eNIr1zo5KYE4AuTcemPcEzsorm/dTKoujr/sk8hdaZXVeN
op/SrHVuSle0TmwGmI71D3UAYfRK5EL1mIa9PSxCXho59qdoqaYA8BEpCd/LdA0oESbqixY5oSX7
Bsyv5a5HZ10VH8vkgoiILC7xh384VQhlKlBv6J6rzIJ8O77PLdVuklHLZVNi2CRa1tMWLBVX757S
xJsBXOwE6sV4lujmImas9JZDbR+CPUYy8UfYWSnxbVgwEROQPCplSgsXCFE+2dB0u+Rnw+HgaZO8
QzUwl25IR/Ye3hbb2gWormeIG5qW2oDpazh17Lfy87jEkpPBbl9ckF7mhS/eEZX6tbvfzbztM/W5
w41DKtEQ9wmcuQmC2q5VyQX4P/pPC/m6MIhaHxtrJ5Ci6cJTqBBMAcIhg7hmxMfGfycMN2yF68Bl
cdJzoEqqJcNX2r8SkAIgMGSGgcf6UAu4v5tHaiDAG7lLq4rMUC15CvQWWqVzdJb/LTbHMRg/NaQo
RWLGSjflbYByBJ+XX9IuNNbu0huQJCSo7BV3T1SC/6L78AXA9tN9Q0DQRndaPKA04PEpkfm9OVyR
SFwWO1grYSHLHGkj0jUL1PbmWVhXGVPb97ygeMfnh9YD/TTF1GOqU4ystq1e7mw9SgTm2nsfcBLR
yrcw5qPNl/ogjBSjFS2tstk6ya59fUhEfYKDcPOQedsys4kk2EjwnnRCHlFDmFswLjSZVFPNNeLb
1REJQ95U9ic428TJOoPVvAkTL2udemeMf0T/W/bjsM4rQTkz5WQUg+pF+dMzgs1gVOHP16g+uht0
MD3Oe9vZ3+ocuLRGo5z1WrbMQieWwJVbng7N8KCB+mLW80GK9JRnoibuaIUjq46K1bgetj22Kkfk
5EAO4e4OkZgShW3r/se9YpzlXZTZzWKOotlwo1STB07c1BsceFZ/KBIuomuBfu8MRH33LlUmepNf
Yo+zlDgmRUJ6MO3n0mJ4qD6CLUvI4h2pBEdsCrKLkSwd5WB3POs72taiEQ47nr0fux0oBH30LIcl
O7Yc5TDJy15wkpRfSGDIJUOx3YROxoSVdMDyd0m/cDgFLiPmp3arfu5T1ueFfwizp0N14t5rYzbZ
NDcwRSAdMsjKb0pP/E5YwQkfX+q2D1VjjHjVvSh3JXlXewYEvFiO9hoh4YqH3FLe0pDKwOQw/fYd
DNZdpYEiXlwAxfQMAy7AtP/9tZkaRO3phaUYU0YduGq2D17VxLuWp1A7YgqGSDjtDq3wAMwdJyQC
yfAEA4MBi7NxHaRAdN33ivfMSp8FT0KORbHd8ExMk0ebH9Q8HyzraC0q6g+er75ybZ68O0FNVj/Y
LhWWl7Ilx6oAtxmeg8EB5G4Z98CgGV5JaoRDKjDGFS61HzAaaJJ+gmcZmcI2ftT7kqCzyA+G+UD0
wrpHpGbuXZU+DibyWk6chpd7KQ38/MmP/PYcqiqws/Xh/fUKiLNbElmvdckZ/yu+BkAXyKYNnQ9m
Tpo/g1XMedkkznm3taLGn00FVD897usf/cyNUCqtEHSOw2wz3DOxjYMafZJkotDdzqj5bdvg8YYY
MRlxie0TzyRZRxSPgrV19xIRS4RkoBZVFukSXRqhvacraJ9p2D6+5d1D38MBX81O3+vsHadzotJx
KkGa+C9tLXNW/5iwuzl2tXi/JerY5B6XbxJb7MiTb3wdID9whIi82Z8pq9afpYFagkbfaNbHp384
GuKBFyXVnXQFQc7N6Bg+t7OhRfillTRfGVbY70bxkI4pFfsV/2CIw5erXFCGkFczDE2xcUlJ/dyf
7LRKuX5BNVqayQc1fvcccd4OCEvMOdCFtNjpIsngznnR46Bk2TJjr4kIAjxeXcAWmd7ZmrXfM87T
itewehtueeprDuOxRL8R6qTfJ0xBkc9yNzxGjmzZXrVBWh5MmBZ14nLCPGbi14aS8LXPcMZ3eg+0
buAlXE1h7aUOTPSqgQvOoPKnDMQZucI1sefD3sOriXsJvc0e1kqUJv09/4Hp+sk+X1lTp5hj34CC
R6smfBvFVOEM+JeIgbIAIuOEKXMowZG5VMWzgYw1maMZm3F8M2pahoB9RZuxMjfbXPoyFYOwDULo
pfG/mbQ7chsd8rGz4kzg5lsxMViJt2w+pj9Od6ZPD6HieRuzX+IGgI2pBEdz4tCYXrWKbPpHZoj7
NwoOQ5k06u1SZ3FrLtxKi9IGWmdtIHmHqHXR2AVMADrxtwX4macv5Znj8uT2p3Gbtdnpj6W3Jf0k
fY24Zizus5jtnQGnF+RMP+t7+L9BvfczJiemscaHcW6N50EO9nw6zgvqUN/eY4jN7F9PfJ7hf/Wf
V+C3rkfIy7RZe3TlmWuaqAggREOKzysDA331T0YFBYLZjL2MWYsR0X8qzy05d+F+8sFJu76/DrTv
lxzxW0tjqeK1ogSj1YvpCCRoWgOJZwkyUpcsG5XpJuaX24QoUjlTN24gclDWUF9mqYLrjRQDPJ6N
lkT8DeN5o3mMXaSBsrd/Xe10j7CAKpIACU4LWYBIiU5t7msa8psQ3mTZ5PS3EVPqsU6Q8huDq7kt
ggML7AwVySOLiFXbDANbqdDM/I4olgaoWj82wA3HeFPNfihKy94ZmmjhhCw7vBBmtxJEZmQmZ0Gj
Ul52G01D7tSgs8F+A2qfa6s/In6KdkGSXRJryYQpy7DT7o/Wu5wBRXEBm8qfMu26L3ht7pHzNcOF
cMZ4FRh5Y3p+HhoNWsiKT6ILNv4F7cEQp79Qxf1G9q3vdKvvdhEd0U1bMgPZxXzthwIoHeAdxUAo
Wlh2b8Ga0IYs6rwDrUzQ/AL+zYdSFfaCxwVkyiBr5aWOizcZYVT16x+mWT7/uCv+mUJqAPtblLCr
9/Qq7fOVagwcSsXSGZuLSgHCKvK/tGJZKpXU1onufpJ9UZ3fWdSU9UGAfGD1+tYU7quYEtnhrN1z
W/Dv0lZ41G6zcEjgshrMx78vLnLzxMzXJ+0vH/d9yCfZ5WR19d1vSmkEYmnVStjll6R1tI4dybct
xWc2Gmj8PuTnJFIJnSEexPxx1XX2fqNEOjCB6sHKAnhNRsvqSRxBmAAY+PFbJjvGLVhaDLNXTw6x
Gli4fUFXjyiozHQ2bBgrKVM0tF9kVRS+czi/H5rR8HsnrwNsTsKC1Y+yiU92kpUrkFsaO8IAWXZ4
Ze9m+RA4qJg+sZPL6NME2LfRjRPuQ1rDeYOQ2FbZaSKdMkfQlAwjm3XSX/F0ZmcOz0/L/CwK4+Rn
Vs3K9My/LVbTA5Ov6pyxz1LlM+Nt917gWeoGrryft5d+eUNDosqZEn6VTFIVJK/ZdWYpjL9E9UNs
QqwtE87QdH/GrXSuzaPPiGHt02ZV4PMVWe23qRUHIFhxUjvwlRzORPG9MAJEQ00gacDM35Z9xrHO
dFdN0TBzzS/3KbWZYoPWSR93JdK3+YOOZu3STZL+yAUHZ76mi/ABZOBZL3vzeOhPp5nWknTxOLpr
8pwDlSo9rkNXPJ5VBrTfNNUWB/ZUMGw9OAupMVLuBv0pwnIkac6Mzlfrg5zQDl6hDzAgn1IDm0Ny
X8UvshVql+piFlW0S70Lb9EMgJvt8Ze/p/5SOLwvRdwipW/FGZmYIoXuyV7PNhFqoHaqAd/qunYf
/2s+ru6hobnaHWaET2G21HHh3bIbNcv+SQUxEg7c+m7Kji2kzYdZ2ZWI7BomSH+/Zyd9clhmLpva
Pxj37ClpzR5rHqNmS1WJ8c0QwXEwDXbiMzbJ6mLImRbu6BTF37LG5nUUaerJ8bKU1qWnwIhEWcps
o+27ob0cXlQ8YSsndhoIevFho/63Rz8TIT//5vLW0ZYKPt0UILe4COfMEkLesg35f/WvCo3fXFfu
Ew903N/gINiUVHbQiMFqXcn5EcLpjNsd4d+tftU3TjzZKY2k85sb5Wc5LvLGhtZCbWjwMcDKF+AO
kY1Nlr1Ek7/lrP6pc9Egi5XUtbNyz7/FpQHJvH11rIJmB5pWjL2+MjqzGzHVShEgWNzdAASSIz1D
H5C8WyaM1jS5HOw2DukT9MX7BhJ6CAZa09QCcuGQNGGaj00v+R/dt1A482Dd/eALlJ7dv843/Uu8
m5k/3UhcmyHL/b/+vB9lMUuWu4nXsTwa431cGgmNcR5Fop6VV1qZ/eCVWfPxJ+ZfnUaU3BlfMfx7
Cq77GT5AisoE01zPXTxR2xBMK35n1+q7ZTHAfP9rPFsuFJMuwABTVZA+raCDnlkPcnRC4aNRyXvf
vg1KIsIatVeWvHKMjhv5K19od0Wu/fY8WPv5dK/uo7RQJZyQx9Rt0ieE0YDqgZBKq/8wVMJhRNFN
ytm9J2yRyZDO00RWwpCziiaCgljGHqIad5NXEVyfkPCJEdfKOmhHlViKiZ0C5klCMDWCUsbzWlgy
AE+VFoAe3tQycwPR8+BsCMsu5glzw79pXGeYmu0huedGJM8RJytFbsoO1J63clWppIfmxldQGvPw
/qUsMdy86SXAQjdVNjiI9xSwEIJgxvSyeoYkzJcn8K2pv+n1L3vgVNjWCOGajiQpa2793f19y+yk
aiE2FUZfBo2xPieez9fClw/A5VYSE8+gvMngqMrAq8DBxzvNOvHqKWAC2JOefgM3UeWmF6MMeO8m
Jf4k6PvJ1BerT/pJ1m/SxjN9w2fPFe+7IZ6rSBA79NfDRqXbTQO/gimSm+Gos6h0GZvexS3hmK3F
vK+PAlxcGd4Dn9t0S2Wj/v0z9CSaaarqTY1gIZkKQ8E3c/jkaDsM4sjfBE7IzhT0FWPsi5C+2rlU
AYZ3UbdTypeHLRRLrbUaHvASywxsFknBPbRxygd4R41twnZ7fLeAX1UTIrRcBcR1SUL/hW+Vylep
Do3+Xnj4pSTqjF067peJnzUhBF3Cd82md31G42uxXYJjV6a+VkqgSu1B3cmWfKj7vCJwL2+BqKAF
fvolhbv4nZj8L5wfDLPE9Szfb894RmHebdWN2WGXM9Nj8F8lDEJSg4EYEatbkB+eaAJA0mvJBt6L
XON6MTRNXQ9c1AjDILvhGTCPElvSG0Y/+j41suQuHt3us/1MYkpw9eaYYj2lFy8IrM0m/35uS+Ph
sI6SpHI/k5jSV4kAEeb6T1M/FIl8HOrxX/LOE6tBnyEgYxIKw0LSYs96vdOkTM83+EJHxtk9a7Nf
X66kv0wmiTEuEj10xYh76CwjrCBAvYfts8wG8S9vpDiStwLJhq47+z3LgjB8C6vejQmhLhaFmK9G
jzZpPxYSq1EbRWJDlTT1blpfEyl5UHH+KoX7UbotQm6ZdcBYbYjF1YFFaFu6PE19TAmOuKVphgsx
AiiUMh0ZQ61kdd/AMGDnT3Ucs1AiBsxGoBL6hU386UvX/QnZ67JqL8afjyOTOJoaY8h9THo8qrfR
KzE7BQb+U7nGcTH3BbcNIaJJgZslzNMCW9Msd/XGfmbQupUQqBocu/C7KUA/ktWWYVUy1cDyMCGN
6UCHq0cM4cKNi7OkcoZAx2zaI13mzyE5CCNpeg65PuncfBBakKUZbSEI+FhjFMMs300SHDh2Jtpb
+6CzsdUjj3sUDjmsGQ2YCzG/XIYLkdJrVkXx+Z6Ojk6l5ywxaawacO5AlGikp+NTL8gj4pZSYsDL
TrCiexrxDcyoXgb20eXeQdGdN1Rt4YK0SuaMVUeV0DSMCDRyeVHlngLWD1cDpoyQSoLDeeTbSKug
fRELcNfi0oER5QUOmpnO8ESD8Clzv1p4odhYrJlHxfa0BZVKPbj9vWelAAETBaAnxxUIQGrqDGdT
B7PNFxH+ATPy4R3/V4gnsQaMDfSnJYQp2JhVfPaTfAnkeN9HB37hHLDHt1IW8Y6GifaS04vRExaV
yKkrgfmpILFZ+OGEMZXt1vCXXqGFke1ShZkrT5p9eqG5v4Bnbq+KhJB5PmOvBuy/5EhgNfdWA34i
ocqHf3yn7q99ncn16BOoAgL/v8aX9JY8PyCB6rDpqJYWXiK0owx0HdZnjf9ZXTKU13zGCHsy8+nv
OC5yBejohmJPzHUOp8zceUCHkVbEwPVT+92N/1j8O2AtfS3obxolTtuVUfAK7WV1l5PFMrc6BZNR
/fMeIn/iOsMCA/t5CGq/1x4w92dP9CO677lWCj+E51wParCBYnncOmiAxs90CcPRDo+P5CQY5oZW
66amwMokppBV5mCvLwUhgBzMx4wXkSZLAgfLwF2bJS85THJqeCz8rUnC3RLCEmvzswELd/THKtaw
u92CTUyU09v1BHJZvsIZ2FQDxOEms5QKwGjICMrmt4s8Y9qbHXRA+xJi0zTKcXQR5ZRnRCMKnhoz
iHvlUMZ7+PJGwm9q8gglJGHEoi/7Mszcw/jtXnn/zJCnrxMl70EP6Q2rEBpBSuhLXg7NCK0qAwrb
eot62+QtU3FYx7UiDKQi3hADUHUc2xG0UaWbAHdDOnb6KjFgYWMpysXO0Hgl6smBreAnLyiVEjX2
Ks+r4J8jYh9+b4k0mnTEiW0r0Au03zimI4AKhiOx5jEHSyL3Tkw+k0NWcj2Q/bEbBKCaHVjKMoup
RMAB1dfQ6omIV5D485obgwtklQNsrh76MGNxz7yauMFa4dcdasdHkUNLKL5X3XKPkNphMJxZNLUf
t+nAyR2C35ZPZF+17W3TRgjSUWFj8O2kWbdXPmddhQjIl1qPgYI63SfDQIjyDKTKaIFVMTFn1Pag
cmhRe+aaAOwIjbklI2CRmgc+OitvVVByuHl/PUMaLQSEuBtGSzgeUGXQA72b1VQVs56i8HqEbt7k
ShSYRKoKTStVsYy0Q/klKNji7HFk2GnYohJeVr/Nj3DVelbEtz+NHB/O8bFy8pUcWacbeVdRfvbG
uzXdcsDS9D5Lx2m7x3cQagxjQTye4eNcyWT+kj4ZBPHP0XJnwazSBCOUMKXs8UIOFFmUR5eLt9Au
04OKsig8T3PWDRkqzmg1A+UHORr1gQENbtFLgHUdHC53LN/Zf08iK5sNrrR4j64HocDKLfmvwoDm
q5DEnkXgoXHQgFHpfGC4ncxEYUo4JBsTr/MyhrFptV5cWPI//xGw0kcm8PUcyultOQ4kdD6GKeRb
wNRsMUBYSF3rZTloux+4MmDp4iEaXBO196Clkfdk+fMqJWsuhx9rN5onmFaW0Mp/u5uUtlIPbFrA
1fdZQX2sVwtZiTsfL+wVnMz0HoAdeWTGsh36S8oxn8/afVvibN7/PEbeYGQfWWpAPGC/8C5U6q6V
9w0XhNTpcAzVlknCGSMeKJtY3TrT/iOpSYCJGS1K05c95Rw6S09z2LYIuiqXBcR2vOW0rnO9NYc/
UhBiex7BMYN2wMcvrRgNNV9FNcN847xAhCNpfzV16dtYuZtjjjjCp5npGXkij647lJCAm6JdaTvg
JfIQi9bdQaLsYQyqjASZGGWL+PO/NidBYit3l9xH0OuvLoY4lRI71eXQyAFvL9vNtwrKuvAgiJUW
srfrE2fQIxcQLatpB/B3thJaKOG/PVRpyyfOevu+ArPeOLSh1VkJKer+g/qz9dvWFmC5LWWSsNc5
8Aw+7URVSd2EaKWQ4NYBHtTZBeyyyuwT1T1HUeOmEcZYh1W+KxHlRt5q0bWXLKi0+isSDBEne7Il
QtK9MGqVX0/e1+g8aVyfp/SSleCk1l4SeWbnRN7g9GITFpka2Mvi99Ip/GiDaZxx9BwRsApYncsG
bxqQR7DzBA8IFphymUGko7+fbJisqSisg1sZDVW4tGo6jto3ZmhCmACk6Trf8ULgSxJVOPkmPaDC
5o+g/UjYREF+XIn9wxKPFk7mHaJGjUHUidNBH5TFpNS9DLwDWrfmYGzlWRC1sw7GTPMxU3Xl6zNx
Z+9wjRd2yF+s4NKcgMeA3qpLCBMI32q0so4fl3/19cMCVK9WZ9h2GSCPjh2/u+bCE/qdmwsmAmcW
4FSrcdGwnDO0zBJYxprg3VLnE1NvX2m5fqIAkM89o9OBM+1CjPH6rO8uQVGfxMhx24bnma2Ydmrg
oWH12+P2F/K2VOK5qlKmVGY57BzUKAcSfOfgfc1yhVNaQ0LUylgZmnbJ/UJcSRilm+kk1FadEn4m
+AvLYA/hXZS/sA4aUnmAk9qwM9NbwRijlBAjiWV51ynq2CZW+Bydt3VKengdX8whKwrgaQjsrGEk
5CiSkIrLPaZSEgnm5olKzXymiWv6xc1Pe4pbbWb1CpqUXTXjNQuSdVfHOmUkymijneoIAitO5Oli
ku4vAiJ6ScGRTyf4oRtQNxWByFkv4hdDX0VW5waEZrLWf2FJA8FG3HlW4pZZKysafn6H7NjuCRSC
M+fE6Yt7wnsxJVUbwLmxfzRp5ztYurNOkJT9pj8zPxL4d1Z+TxkHB30jdxY4n9vxLpqmst5JUBH9
gx86PtwiW7rcV80hQF+f2N8OwGC5gcoiU5AVGwazUj0s0cEllMJlGD2bZtLmM41S4Ed4Km+F+Nzv
lFOVFXlMh9+TBqTHoknPa/gErG+zmx3LYAwbArRgOvHdK7hVplWM9UmkGv6IFaRzON5WzjUq7HTb
+3SNzg547Cf8UWV/5+kSh5+AJPws+Fyb2HSPzY1dke0cQxZcZk9z1i6vbr1v7fCSsiBnWpwBwZon
tFUcJKgb/Qb8dlVNJtAzMzC8zCn/F8M78B0E1nU17TOLbAeORzpv0ddD9Ic+E7K5X+HmmJrz5Iv6
UDIkgl5IHknYN1J6HyLK1NehZXXUMwNsLnkoQVoUPG9k7qtdgAL+5ZDoQ0WsoyNTFHQqo+WLfQXU
P1QH+BK/01r5c8g5k+Z2K9AHWD8i27/6fqs/gFKH2IZ/hH+nOv55Pk9uherW87Zy5IFpkFA6wwuz
EZHqFza6e4VVN/Ahu8hWTjYZ6yuGYv7BNuuG8gMVoJUDHX0lNVmaLZGQJHzL9Km2Q04S+bx96xji
AxcyJiW4LeYftU9HKDl6uIb8vaMq6b/qgyNSkGm20WrCRguIQjebxR10Dyu55rvE1v/YpWMzKoYo
2WtSKpM3nExcEqYQYUzdax0g0Mpv3WBtkCmk2ev+iIFH7f3beTft21HJQFlzmCMY36pjvv68jklp
I8d0Jrc1Ipj7sk7IuifMZNTuQuyJO2f/J3KSFsE8pbHBwyEkrMn178ZrVFZwNALiP640ilbtTGu8
bjkSeg3dwoQHyWl866VK/ntQSixcCT6WwgIghLAh69xff2yoALaJimb0RgpvkSLYIjkr6yEp+fjs
TC/2HhO6Lx9vrQcTANF7zCyNpPomAHRMxfd6GCy26YFKzOJCg6c1HlZsBf7om6nO5nE7wTqCkeAi
cvAyvXR+TE9z/OW0YPanU2I1RnPfKlttDiElVChp6uODppIw5oycQTajj8y19mc7pGxaMCPgjP0K
OQTd0Eck2VoAEAl+kNob1MCFc/gmgkTTfJ5yw62k4M70PvCTjE1wgPD+3p+janay3JBVcX3KrTxi
VA9tzBE6z+fZnYqBRS0nez19C5SyluCd6dIYmaABQL6ceUgS+kbl6H0UnhyyvPanmzCSdf1xR68v
PQoF7Z5lA9kNQ1MOCOd3WA4p6sLqYzT09MOBxeLYvxvWuJCJYhCCeqwT//iSfWTVF4pK/OIfWrp9
1fEH4r5XUGhokIar4pWWcxNMK8UXJO2QN1HOemygOs2D5NA471JJHTh8fPocyL9MLiDPB2dUqDlX
v6UMdMVqeEuTu7o2uS0jdv5nKw/zwwqx1tICjtKJuUZTOaXjeSc368Yzzhb2/G1cLvv89YtiNaci
o1HqkJXuIQEsCFiAPHbmFcLyT6iFszdkBzG6SwDBygGNjMsXsMkeJ9dDxm2s06SnqVJLf0lT4NKH
Z4aYJ48CRKFNcjI9XzAQexgyyp0TpqpxxY369FXJBpavs09E5ddDvvseQtGZO1uKCuuFqIZdz0lc
F+eC+3tyUFHVlWxcVHd9ByCr288QmSkE/HDTfAV/Rg1axL9oKCGF9O2n9GJtzAImn9MA2oejn/JK
wci6GVNrGYZ9V/nHd+7fTCg2iZLhNDXXStt+ZUGRx6LkDMVvyAB2PvA8sx3gbNybcyhXqP8VmGDt
7Lie5rgtWiZCdJ6XA90AOU1EGPzcfjpkb4rhLX6DnlbdSRhOlmHnSuXH9m+iS39uswACFq0OVp3R
lcQpphRLVPbtxaZMfsApsQFFSnSgxmAYRIYWER9B2ml25fcVlop07EO4Heq61rHkPVQqASJhya0r
9ZmFUp3kFPQn1tTbE3ju7xvEoRXDZuryG5eDO886dbRp54Ng5L0OcIbre9uQXJYdzQqiZcwnicNA
RxwiyveLmHgPXrji+asbWa2V1dXBXt+znPXqZip3DLVs46E0UGoHJtN81c0hxGyAfj5P2nfnw6oU
k7VNf4idDTp/l55QbWlm87c8jdTDgFnIbe1hpIeuPKwbRcQZIQSUtytUTF9oDyhihd80SXgAgutK
UPtXeHWqHG6C0RnTlNSIrB1T5FtIIPCen0MXDgyimxtRe82tg8/dvLcrWEcjPwsMdVa1Oi6yIsPz
jd294dS9LXBuLVjUk0iIx7qrmaK4SBiNzI6BSNS0FjADhTdPyNF1gh+jkEkDYvwvOw+CILiIByqG
+p5yfaI7vlfEgr7kOtIb8pdbIlo+jo9/RZR3O6dyGpQ+7uKwWmrz+jL1VnozVCGjYnf35WLWrg/7
npGslea9X7uY4Aipk78Vi3o8NzCk7DXDhZP68OH3jjLM+P4QWLRSkBhnRXUjSyiarmR2znQSMNo8
GdG1dTSJJbXNRPWdE5UAA7nDgrh/8XvIhooIHtQOzHadaVMXVIE7ccZgafxa8sgW/pHnFgSegzGZ
EusNxVlMU8UqwvwcJQd3lI7fW7esgKl4GrFNR4SSLAEsRzn68LEOmStatbjToH598MLPb0LHWwC6
Am1aiON2HFgcsZLdUdxgHUrLnu0Uu9gvqS8ohHqOYq5CLn8IRx0tNpJjlvf0/Pp2in6vgsM0Tk7v
mVPBdNkmCNuARO4uasO3YDA2lnOaTu65W7t9SRBQNw7O+Rs1kXobVrHdsegUqZ5fWcaZTMnWikeJ
VU6tV1d1SHf7+jlrr1/Rir0At6GqBWBS8+wbFBiCnmDgooDBr8SmPWKg5BhEiHeppQK+c15SMcUe
gufgbQMR0Cwkk5u4zKKfSPjcTzK5J0TOIfjcJCBOUa5pX6Yw2oaeYykIx6IWyAEiPlMxinGrT2RA
c5PUMtemHn+dV/rgW7u0cSjszUSZI1ndU2Dm0KByDK5x+qqGwCD4xl9v63mLOIx675oeu/OIg5iw
JLSaX+O9uoXSez7+UpCTYQJmEfPKNrRiFUXiUoMFREiwTp0n9o/oJlY0xPtLkNEBUsof1zsr+B66
7f28eMBLIx3K0UEDYoRSfmHMmdXi88gA7Sp+ntHqXtwtXQL8iVBPGbZPgcRmhOJFE6TwB+R59RXQ
h1HRdMLkNy/GVixY2VfU43zXLYhIdNuDTCthkRi/zAYdT/FjfzGoz2mrs+sKMSqtMrLnsNOG+MvE
qoRaHyTvqG/f7GWX6TXVzoKzrjIGA2S4yShefKv7i5A7l+daBl91LbUj+PYRraFY85dNkK7GqjoI
Wi7c5izIRfLJYsbZuMSk7u9Gof6CrlvBcB6e1Pr09YiRczsBKOr4Yi63Ys7ASSfulWk9zBGNy1mp
HP2IJYLyjqBVRhDhgdZEF585Mayn4zaEN78GXi0rPCK3KO7+fLJ1/acKMe+Mma/ogUV0zYrGJ3iN
FtXTKtsCZFRj39BouB3qT3bV2LIfffSLpaRP6ZFZi4FBUAHtUT/BFCx6B5Ypi4pZdImLQ4ACLKL4
Ca58VuE3uB6egPJxgaIm4osTQQlrtqrgaYXilb8lpllsRMpfSy09BDbLD7BZa60TNw4IjmK3PhYm
unPAyWk0Iwq45gkx0mxna+/6i+LCqqH3Sgz1ItmLIvdJ8wTE/zj3NrgNmY5M8ZW9aX9H27TlX2pn
MOFAVFPB0fiN3S3Va+y3TbdT5NrAz0HjYFlMDUG1u132p6X0EYeS6OtEVSvtFwvGf+ZWJoCvA4XX
ucyFNkD3YAe8f9LfocWmVW55D1LMC4Q9wB7ybDbco8ulIHXy/bvfcT6DlW6a6LInVZik6WoIl8wL
empeh0MjVAt4MVDqK11A67jnpfBXDUZfoHLT712wB9XErAeMciEEaTir6Cglld3VVfeBx9yY6Goj
1O9Y0Amd9vbJ2FdnYc0pBgxVsYUe/L64PHqJm40uP5F1aVeR8dMUCX7TyNTjTa/eWgl3rRvByDBA
DmIne6piATkTEfTjAmBlz1VLrU/4reEXz9dPNEMNMBXXVKB3exUlsXlMcQUm663nCf1HGhy8z+qq
n9YV6+6nHZ1atdh4JG8oEcX3dcf6zyHWLoGynBLjlnec8a2y+dT0Rh2X/Xu9RuuahdHeQiEOnJZk
BZRVOCx06s5B4o4FrF/WWDU/J3TDTsmxPaQZ7t2/rtgg1cwV2hM8XcnSQyhHWPE+m5qtzTcCQlyi
wtQLAgzaZfYvTK5fq4eFzOy578dAZaO9d44JnuN5OXgs7+xG2ie40wu73YlKEp5se3F3J+t7TJcR
gHEZWjuOATOSJyhcQ015Jxxplq/8/PlMFBMLRhu2IXEWkb5A97WeDfbY98kpTTh6GXT00u+h/Y+e
SiBydTspvoB0A/yeGEkzgzCio4VVIZor0CpCP6cQz7fCRmvff9DNsObpb6GqRQkaDTA2V2TVLBXB
xAVneKRreYNVH/OJ+OZWUSAvDQ6CG66YV93Asr6wns3GREIrRWOrEhVD6CYPxEi7p6ohnpJ0dHSs
hr1PNRCYrUzSlgAtp0BFTbHXJqmn8Osb9xbMch+HfkXYdMK1Gz/CEFzQ0VRKtQ+KhDh4o6GlclMr
XWvw56mcRGevFvvIHFj7Jocadp8OghcTBreEKVTl8we+dZXejIoN2IRGrf6IdD14vDYOZuWv67Ez
nqv8EUYzXWDoZHNTR4i04627VC5afCfK+/tSgTMC2RAsIDlPWbIIz57x4tfyYJWfWkCmWD/KTFq+
9QezjDKK3htrNlHpPtfHPRLSPjaVYsEBB9ZwXPBIBNgZLlQRpqXVyuRmJ0H6PJTo+l5MXQ5ja047
hdB6g4ivCC1Uu2PxFwfuWO3+Qa8H5swY+nkPeo0NBhATuisSNxLI1fdcKuTufIw3gelpIq1NbRa8
sWEZIUBcEHvw4LNJ2FO9px8sJfWV6cM/VTf8nAhOp9GAWdSgungmMWzDpkLR2GVcm31CZwuLdg4E
Oj4KjF2W1tVQ5xO3y0RgKLkOrr4bJOlCXemJfEpK79siUU20D+FCzBc7kh3nLJAXNFsPHLhwU3V0
0rA62N+CF5QG00ASlzejaJC+ylpzWLIRc/SSEJckBveN+N/XGnHLhCR8baJXLdcjyo4eNEN7dN9h
cbE+JsGuB0Skrh9pplmPQjzlk7eRCmd1uZcJjba6N2CXHTD8MjWZ6gYCOcjfx/INbfH5C4QPL+Ha
hJNUkNZ219TboPf4H7yuGsEUx4o1xzX5iE57uKtBAPmnpY2RbFIvaHsmN6ennek9MgUxuze5Q6i1
oRVaRp7eLdF0YasYvSb3FieYgUXmEifsldk02pDMGywjfntDs/XtRHC3sWxppyI8NYUnkI5BWo0T
o4ckn6QcFDmw4F+1YBfWlcCGJK1UZl+Qp/KDtC78y0+QrWXt+RRbSVPg1Lwdfir2SwchRZq+L0Yh
818JW1bYJmSxloLN1L6kiGxAS6fEQoBERcHd/Fw11Vxx52TOYXWme8YQAuw08rf3Dzu4yb73g4b8
LKTwbP9CahBYdAaXPXiZU11cceeTG9A2sm8XcUUH4j3YELxRplGxo8NDCp8ErCRw7iF/Wb9o4R3p
fbZ/TK8qhGSAIO/ClTZba9VYntUfR1MCligUxSL0opPteTOWxpZgEbkQROzgKPOvU58Jpnm5PeC1
WcvvUePNO1Jf1Lo2eJ4O2EyaO3xUiDYpzRl/XHQWWuF1qfZq9INqwUsVVNGRmHeFVwrHc8a69t6t
nT/1iGsuIg633yTACol0lMVKwhyuABdinMiAeddRuUezW+bhmbCyTcEj8p08F7T50vdbIvVn1ixM
Ik1haap5+kt1jASwa0fxAxry3OhyQRQd6zArFh8KWQJPmmme3QEyh1aGJ9Ut4ew4LvCYBXuXZmfb
S/d6bxVQ7OKqrZv8toqNsciz+YHDyHAtwq+0Cfp47Ahvyr1MnQFjRDSmfQxqD2AVphTu6ketnajZ
/bLgQxA1blNsetKRJRlfZAMAVcghNgc8GhrnUFUN8mUUDyzAhVAzOiiPyG02jtFX6sTIBjxm2MOD
ZS8dfs12rOZb/NSYOXTDggwxgfV9WdZ5Zoe3BV/9moYWXLdwypC+Aj1C+VWXdPeDYB2AMdbnW5AG
i+KDtrN7wefz6Tr2QXEexsuhwjNdx8vJviBtPeEE/1QS0rhoTLhudBZDMBKYGGxJ6doEWsy4SImT
nzM73TnVnQGWjjnZUHoPFLL7uw+46p0mjIR0pZx84gHNmPP96/Wp80nJE56aTWrAkr7REOyL9yd4
7yhNV9OhmUC0rihtx9hYaoE5wSHVvHPlTq1IlG3pZtfoIqUxzBBW+YPNcvmCy4IOQYH8JqMqQE3q
LqsHTiS8xAXZNG31fyMTCc3dH9R1fbS2zjny7MMmOk9uIxZxYsoETpzoqsDZyjdxwKJKiolY8boM
qjg8qc55Vhv6Ir2mf5eDvriKlk8nPrmW0yNHtpAofACfED3jTxtW33v8LbLCdKygK/j+H4PbWjbi
SgDg8fW/rjstonr45fDQXgybOUFZ/0z2GYtc/+UMNnY0Hqr1gbwG3A/3eAj+wQP6M+HbyPvCHnf9
uryt5E3SFpag4smp4i5h75nALSTdMLCHNfaSQ+a4st1eUq2FdqneLoSp1AFpmN97K7qNUmhphwab
QoiJgwhSgFaKVFXZXAIILbibG45/rKFMWD1n+eSxtFf1oI+i78HZ0Z6RtvAoDPRJwJTct05XXrXL
hSmcdwlW6IP70+zV4GbhbxKn4SaD3a7xX9vItqZLTP03+NbT5Y0WBykxgTdyv2JaXwbCrjrbaDVp
25mBTaPO1+i3vrR6HRiaDJ3p/M6H+NEFLDxcUkctrxtwtgYBX5cs+LpTUHajHY8D+dMYf8q3ni4L
rgQkPn6nTZ6vrD+AD8GduyxH0O3aVRY3+iXyro7DeMmFu9OFEihzqh7abTx4yqPAnnTPiedGuc5a
XYsU/2ozyckm8cXV3OI79s+E5AuRanCAZ3V3KwWQmiNb2B/IktoMs+F+V1yhFS6kOuiz2zrCnRxx
Dqt/cE/NXgou65FU9N9FROyTRoVOeXcvUmL1ATBkjXcOlraZMxmFa/kK0ojCJuxoQXtDe20Qle1F
cpV+SnnTaxq17fSIm0lDBPYHRq9+1dYDqlpOGbO8bRqqYnWcbdgjv37Z9cv9fCFive/VAU8i0kjs
6dGCWZ7bc3xtFyXTf5PfAR7mdmXYrTc5WCgbJKJ5cAVvn+crwb9fVaz9tmxkxdsnNRuZubOyecyS
Jm4f9B34HGFBZjuYP/AginTXnaTiCnZoMRL3iiILOLDToqCki5xoRFRk/icu9a49/1xmlKex9YN8
X2MsGfw5jgvtzyHMxuv+pL2jZ+Oztz7l9E5Ur8hMCbbC1VtZ+mBj4ngH9Fa6DzpjVPfo6L1E4WD9
RxcNDel9OhHOphvNNqpP3DAnHU1fQpgLdTe9b37ZdHuJMTA0DxD8EB6cFHFlc9r7pNAMYpeRiJFg
xK55j+XDH5n+qb5Qf0txR7S4YkvFZG0SG26i5SdCmeSN1OL1gwxNJtjxn6p+rEJ7gUsPn5tobVc1
y6MoQvn9+IG/oC6MmQJX8mHWdtwmArljQbC1lYM5bOrQ64BAIds3/QwbQJa09rfpggwYlr2oMDwk
E3qMwSsJMGpzpQURO13xXaDdmWSq1euE8J4hYYAwJ3tvhAu+kXqZabUVlX0x+3onRExAqN/x/1kL
aqtM+tDpKSW06jD7Pn2teZfXR3yXFvvrSGHMzf0F5qesHdeLM1FzcFYLVV0Rit0kzIFWOnrTSdlh
H+8vlD73fBdww7m8HBX6353mpVUeu02g0DwIug5jdWqFDZ2a520FiY8q8sugEUcYX+xC6WZ+EQw7
Rx/nIDbJrVdPpTm3S7D02zLKnZHM67G1vx3t9nax9/jLH6Rm0RCd7n3T7MA6NjE3J49Ht272K5Ly
+63hYZU5sEOlLEp1Y1IcrvhBL480nruBLQzGYZNgcyywHQB1OZpvvxtwMqIuKtoXQOwatLm7kDYw
g+iY5V+LhS4XlJV+6Ez7fzxow9V+IbqGqMOt0vc8/zNrV1/7P3sIT+0h2W/R3IqPuRgMcVt1JqJ7
hGapPOINEzUsl6UtfL/tsfFso/B2541Z0zbVN7woicw++z89OsgqRl0qqQrdwjCWxWC+SaVNoWFv
J+Hnd1ZC41oq5LFarcUZXU327pIE6Iqif8bqsI+QSeHBZSLCw4AVtTPubsbqVFrWsL82HtzwSqTg
uOOfOSem7ON61aJ5Plx3aYRmBnrQG624QHt1z6BXpFtX1QSnpJ4xLIF07hY6gnS33wrNJ+o8cbtT
3P1b7mxCP06Cu8mOPH2rUA2KowIW+bUOlH1H0buvUCbXZ2rB3FssoJWHwjGRnEMz+IuquHccgGJG
AuQHcwmr82yna9SxcrWa6pOo0arXdMICX/Qu9GBqTJADJAwmD/gRyVz5Bm4tgU+TvW6SNZ2nTTsq
acjk6VtKcZN/nHgj8l5evcxe/W3SLTYf91sjTk7qf9+HZedlXX5YkCdCENWC46pl+z4N2yWyPN+7
BY3qmuG32maaXHMp1Iw7AO8zl8k8dx0BuKER56zGdcy/V9+Ew10uLCR3AobSV0H3hBaTJkOuasIm
l6JbSbniTXSyO72PxBR72VrbJuN/Y6ElfFWhGdZ6PJXef9m1h9p4oZ6pSYAJssSSmPdvm843QYbe
AldolBhjrC7n+ZGVweTEUWlacHIN3ANrLKn1cvRpBRGCzJSWlBKBa4niP0Rv5ONbbxYbbhqJ8T1L
7SjVmHnBdJ1xAcmaESyRtIictcyYasPivrIqK8miuw9rdAzBGfkCL3bSDTfs4+JuocbpA5b+vs3P
RxSJUtyA4Bp+tj09/Iwkp7kJ1JEQnh4OK871CFz8TfzH2nNKygZYE9xpIsqhm1EcmGmD5cQpZeKQ
2Ot8RpCyRxRGI7VojIkblSBtSSHszoBl0h/php9j6kFdiV4H9KzEZixFRBDFJ5QSP/Glr8XVnp8y
efsO6gJOWoJFjouetWbvzJ3luAvFNL2oaHvYXL3Y+0vqEhiZXQoDGJzzEN6kZV/aHyCPWc7kl7Y1
pOn2dgH+xlRRL40txa2QMRjlLdrJv0/FFPopIFern3DCjPvHjSvc5N0UtmVmus/8A68SbQdmurNq
RoGuZBWBv5MJmlchC/rCJLww75RcIIPPwNoI89KAskliT9qrfqP+L1lu9TKk+2DUd8nVEzww+OOu
A44kCrl2J9J0l8AmWxQBy64vWTbMcZGdpFSi343coio1P88uXauLLL86wxj71P/Sb2wxIYNM4jz0
Qc3O9nTWpw774AwhLtChllhPmowGD+yzBkkm2a04PBU7bUHXz7YwjEDxjhSTwtLO0Ba2UyTkXdSq
fUggjYNBiI0zobxEwE9qtZPft16PQpR1hDwrKPdaaxkgqdzjlEfr1SfCmfnGU/iEv36yenFn3iYL
WZ0wuXWkwEz8HOqf/eNs58qzakCrQ8PqhWcsAo+iN0G3Qu8GhD8iaogrFxAh0t16l2vAsFNSCAkg
Rpyobf1+1kAxMSDzKwud8WOpeIo/cW9yCi6JK449o2wrUtqCgLGM9CariEyH3v7eQYAPAkaGqQ5N
6v2tkVt23i4vPGGHbYB141eN+HBSfVXTSKK+hsgEul56HW3DXCEimrk7VRFR2ws3L08UwgIDaWHa
xRrIfmNTU7/OdXQLureBfYq4/y5N7mSYTehBiCSvUWcG4BtJRFN0sH6au3bwrGwJ3AgoNoI/cN5F
t6QOHwq02GaVbdPfQQ1JnPgGAGCjP0NHAWutYLg1LyalpBgaKbc5NiCRmzaTaM5lnUfRZ68CRBs1
l78I+bgM7Fbf2p/V3TDXrvvbHNlF23OwMZ6kyNAX+Y9UHPF2aCcYgJluiMdJWHNwlAai5jnBfWZ+
eQxFqRb6Fuu81+tiRq0DMlcx52HycmuZRBHH6adDskI6LcOUE/bZECBuOwJOTIo9ORlfjKbj3ouX
K3FNBWZh35eR10vsCCnCJaGetAYAOaMqtJtbTTsFlC25gGAQYZPkxlL0k9ccsJbxCuWJLdWiLuBW
V1vFTG7Z4PcWZMvOpMFBPHz4RJUgMayS0F57j1lE62peBVngMS8lO7Qv+bT0lH16S3foXf1NXoaD
vhK1K7RkcM5guJC/Cm1CKQ184WNPUsCRF9LZV/iYnQ0OMxgDeTyCMHPxgv/ipmps/rmqVV/Q5bB4
O89ygHCx1Z64FaBP6b/Qb5snS3eLoxYaVoA9bqp+28E/uWlHTgbjbLafxuyKxaX+z6tADniblCGi
QeCQkmTdRE2nqg2M40KQJeebitBSGjvprgoSP5JbLXKTXiC8ZjVleHzsF5IGZHX4toiBd/BQLgM4
jFqBx4MXVboiqPRvkdC3sZ+vliarH9WDvZYypE535P22zqqdxtZgw1zUlskh7RQ393q96iJ/7MGB
P7M6n1oxxnU4XgXgnKCTGCXVlQrAWVPXn0nsekxKZMDGT9R2fpUYSy7t9JNSKwF+o1XKHWe/Y4PW
e+B5O4Kpqk5gjbhI8l4gEKGKw+foimKHDWJPmFYy1ZiU2aXM/YooDmoK1Fr4kl3Bves+NXZ2wboN
p8kfO6jaqxpze5W3vI2yVJJYNpIcMVMU0CXmjnW2loNkFud+F5qjryVdVliZv7myZxz0jF1cP5mP
3naQ9qqVeqOlSpIc6ZdHy8mGALrzQaWPXIppLuTAzr4UFLeeptUvIARRxHgIUbKzBxmJ0FkCFs68
zMOFDpBxvcW4kw1Ib/OrdQgorHlgw7uxYCAF8dBMp9KvnJmLJh2qkEIipJBPciW+Ut5MUpDPGaJY
tJW5w9xGLKzgMR6u31JTx0kFB8ElJOh6vYcHsmz1XrwsB0Qmqbzn8nfwLeZzg2+Nlgt4cH64S7hh
M35DQUHzrAg428CoqxymzNCuBgfurOiPzzlAnOu49KRng+QApZywThm2f6rzgdSR6vPCjQElhX1G
a8Y2Pw2zdknfERvb2vWWPU8Bbd6rJRxhLvJPlkW6CvYWUI6upDoy72qblwx9t7DrZSR3YEBUzvI0
RyNX4GxzqlSjfSk062VYZn7X1nV+NpaAB2juje6WeHijpKhWp4QEmpgqybQr8x5zu0ZrWXH0YlfX
242S7uT+W9HEd1PObQlM4oXMRls2IerVqCPltkD75fvKdEM14PqdUe+5hFrXa6j1U96+U0Gp6+GF
PVPvKXl3EW5OZgKq0ZRfqhyDK/wSEpZebbHg1RshFyNQiWjY6jz6NhGoXRHGDzrz6sS/KQP8grzu
9sfOkPeHzwhk/0dk5+qI8N6QZnplW7yTDKBPC+YFLW8KexbAyrTpdm6YFBVMJ93dQwNoNbBspr5u
kgjEvirBWdUcPgYZ/suoFU4fIDd7IHOd7cTRCqaq/5ThenUk1J+o0tGR+QoaH01NVpd7/mlTr1Ki
xxL0J4oEbUU3VYkKdeAWS/2BWFm1B7Nc6iAVcHgpB51RKn2XZ8hBy5fiSwUpTYOWtw4TkS4TcHaL
SX23UNG+AgJFViUp16PXfliQvenK7YA+8YZJO1wzGh4jm2efqQh6Cr2DQ2ZHjSrVuHa5n5XnwR0c
kPl57a7QcNp+TlLo7xDo0zPv/QJNEpFBboJcyJ2lOFqjtmikXniv0lLT+cdKKbyoARtV8abfMyYS
u6kpY7Gl8qNMCGFYnYq+xdbT+iiQ0U1S/ZRqeZmRhZM6PDMp6nomPDoSoDALrY3QOWkS06LvdYJw
fGIhkNk/m8f0QJyuezmcqiZVbbrNzUWxc9vJwTDfCANVBXSP43mejHa9KR2lYegDzp19wdY8Ycx3
VGS2oPgM+teAyL6WKRDwXIdEhzhRTrEaWmKcLnaOxNeOgP6QU2Ew+gJNPm2sj+QaH/ztPMgVxjR/
O+arJCqcFWNc5NnEy/wks/ZrsFshlNMG70Xb/PU1evDVwjsAOHv2qeHOeY98R/XYwGifg3mqfaYQ
Ig2UeRyjXR2yudIGf2hQUFsPojBcAi7pxTi357qCp/w3oGJjC3ZuYyFEi7pr3nbrLEekq+hyCfMZ
4OCX8tX7xNinqq6HQuB0iqLGE09a0ATF+H4JeXeFc4a2e6FBlj8w9jQvghMWOe84sjZ4SK0BywQW
biEojER0YNFCFJpxjMzR2ppUNuqC2IY+dYLMXhvC1/GmZLnSU0FMRI9Va3EZBC+o+z76pAON9C8R
fwT0eBe46jJCXnWrhp/0rhg1tWwMVUQTk5FlD72NJsKskAQ9FsYQKzXWu3LjsLKz1THxxDOHS7AG
JkmUTAhITzUU166j01hyWiKOnohGHd83Rfd+Yw4OqHGq0JoFo8QaOFVUX/fjSbVlFh/afUZUav+k
+gyKZsKG9k6qao4IWkrWntqL4gt0VizR3VQ1Qg+hFXHWDhGZ9XJ3IuWCWYCZiULCPXlP6l/JPNmE
xqqX35SP/+odoYCt9lhR3sRuhKTMrXYXciLi/xkse8ezFOMbqpnIC/HyEyrWE+28j+wP458vO+X3
Gpb/3Af9FYEtEaC3t3GP4l4x5qpfWwn7SMXJrgtP+iz5AJ2aRgaZQe7CQUy8SXgGWJUPTN8SAxGk
uqti66uO4hYA6B/+qv9Y/D2r7XVaKw452jM4058hUKbF4d28wX/x3s/sCYNAEOuAsFkDFLxhdJSV
Ub4VGMs012nn4bpRXUIjNMd9hvkBJDAxqTBmm9Cx1c8C9/447CE6A5YiX4c2KRQOepYnTrJAMQnD
9HU5t/+JjMmmwmbVYb5a6TvfVayTMc9OvNve8rpzfdTCoRId0yYtPC2dYCvwN5pdBRrraLmIUFn5
HiV7qeKBtXmYoK6vMbeXHFOjuvb1TWMuPdwBRZqZThIvX6jKqC2kWTf2Ry1Q1S7eyKR22a/4PfWW
FZUejrDBb2Ex7KxErnGja7qxSm5DNvuWwzajCn18bh9K1Pn8lLUo9qF0RJ+2gxu1j6WSkcrgKy+J
vtCOKdQ/JwHTwKZQfaQBtvRr5Cw/xjLFNmVaLioC1suBpxHZkTTzemmMyC7mZ2V54IME+410O5jL
uahL6NOTuCFd39wRyoN02D3UdzToz9gCr7gCcEsnFXrGJm+CbmtcFHC4srYPLqk0a8bDoWvIrxAw
FkwxvE8ABvhg6GnED9AbKJ3esmj00YSJ3CUthmzVCGoto408Fju4wGAsimlWAjioh9m52tuQuBe1
yKftnVJqsS2VylKn6SaMjttdsg30ARThMUUedgxdvJxCUNn/7ITuZHNN5sJ4A2qj7tsV1gCy28Xu
B9/mMTLicRxqg8AV2l6oFmwHZnw6Gyn0lk5V2vb0wTuJgULWaWBOaflnHi8PFuysQgvHoMe8J6+9
uniGlBUrLi+FSVJOzUlK55Moj2pT3Ba+mN63fdsHq9aUOVTr8BTuyS4h7pUps2emb9vPzapaIdd4
d0exb+TScB5SwlTv5uzFxZrG5a4YR8bobR5bvBRCaE3iceyboWB+uo6edecAwgzPOk1r39H3a7wo
LPSz8mjlQZ74KdG+vmvmdPCNRNJqeIA1aoKNWRyCDbnXn/b/UsxhCmqrAs5+G6GMrkwRyhLCdWqm
1ynno3ZRZIjwRDYe1pCs5dab9zNPPo3RevKW1B6PYWmsGAxGPHsdnQhzVsXfNPnkq6PuVCpysOG0
G1DeZKYS2l45TzvJP5ijEQWeSVvW4TPg4/0nLr9ake9ceDpm4nWBYLWanKN9c/XkDf2JiXcras+K
FLg9RDhIrDDWx84Brxd2utsWeDMP0MLM7pbxFtjAm+J59D+EYCDIWSd18eCQDB9NuoullVsxJIZy
AViIQ2YAahNloAiaLR7kvIcQga9U9RUb9ycTx3iZEJl7GskkBtzW2Jy8vDvn8jxIhrrQlFn3hW5S
Z8KAOViUl+mAQUpx/ZIhULpvWl1HGfbL1PAQeLTi2ZkZNluA16lUnshBh5EdG9yO4JJDQF1hfmCD
uAtv8UHKvSsRrGJYeHTF1NtUPl9L0Va3XkzjjEAqc6Yg1qIGBKO+MPIVavg1ZspLACjW1Q6lFRc1
lHvqy+QXL1vrqS7R+5Twu5nw5YANEmFttLzXpSNEYun5Tj8QDtfCwEyOgEGeT5E7AKnQiCNUR7OX
F4E6+RqiK7ti4mJgmA4gT5q0HFv4ELLeD6IuGtoBUjSe3JHictBHb4iILYE21joMxbecx/qVR5ii
vea3xzZofbFRpXog4ND0vHhMW7AkrCNUVXJ0SbygoQafR3yk5O+XPa3IFegE56gaAmzBi0oVR/O2
oNVzu9C0qX3SaYDmh3yx7RvsLqXYK7cCV4d2y5ZLC7PLvBROnh/07Obg/zsJGl/sTunprJQIBXHd
Zn0pgJ+K+i4ulc4l8cPfwr24fAruKwaTGWv5lzWMOviOTKvvm6tdQxXp+fau+tTDjJLkDD4toKA+
J7/ZTj1ee98hCwHxyRjoES8MHClwcDqIIAN5hEvsfeJWkVIGp3d/eme7nkNCFQpy2Si2+AChEYvZ
VfCCJyAKwfqZDf7VWPBRwTpKjiT/OIcyBU51yulFy+jHQXgSnGaep5EwEPyZsXyHuru+z0t5Yqe4
cQcBCeXlgRsQ29Pt1qCO7654p4Woyf1xLcp9xBR3crEMMurUcMweTrshFJn0NnNJouJG1hCLnNfQ
SoOOOWD6h7OS32xI7HyPl6+4cpcAP/jRZBlFnMUKhhJ1PrZLvBSgdkgBg84aSeOql7OT3MXM80hC
yyJ1pBvDfhOK+lGUvyVsn1I4ge3l7YlEs/g7oKNhqHCOOoqxzMFS+5d2YhrsCny/8wF8zm0ajHIT
caoua6HIcofrmr3fudHsLkZn3yZJrUoYqsxMhtuShl2a00VVL5prBzUVxMEg32vWI2XmlUSLHx1x
9k7EUkO8pQ24W7rtYOGSG2MbAakTGB7vtoVN2l8KeVH9wZ5Y5k1vpFnjbHiwgwpwzx4lN3yCdCIO
ZNO69qhpiwJAi+Qejdxcjz4GJwypYPPT/VsM/r2jOjZdk6h9kJKx0NcKKXHrIFssasZcpwc7qLKl
gfO++QDAY+ADXdChyWBR1B2aClIXgDX5ShnQ7ouZDlbXApv1uoRlaR3lGOrmBgDfT7U9eColT0Ff
yS6R169Sa0MA9nhrMCTlEqhT2uZ1VLumbwx0UWsdFZFnFQqUqe3aoRsxKVLyNrzNLWoJYOTYDtsh
S6AIiAvWO8TLFnBVe+f780Zm9sEy/VNZ6A8mR/E5lZ1dIoTE3+9FAkyQxTXKMjl4Pw9aEPLmTTsK
O+kvCzCPjsnda7QytoH5zPYsrP6v5bKST/swcDbfJiM1pY5v5WBQmlivRI+l9VWDXLhJjvbCQ9yS
96W4vdxl2Ow/vhAhWpWyxYEq4WNb8BrMvumbBjy+CFV88ZW3xB04Eq85lwRmXQBOWxvE797e7MxL
FrK+U+5dSfG8Kq99sMRz6SiP0g8HEPOkH13rlTteI08Wp6FpofktDcv+BWHdzkmLbCe1YVZgNMJs
cCr5shkMvE8zYpGU3KjmZU4OE6D08bJWdB4lC3CV+QtQWnkytF6HwJ+fKQcDN+ponB/vJ3BWDbhH
yNW5fHH/hulrGSjE+0vsDrFkVlwVjqtuFfn8lmZIIvE/pdNILngYfFKDZVwIMBlwCgn6QTLit23U
/sp530QMlYx8E2Zffnbm3icN2sIQmyA1YXrO5FgsKmttTfuC7r6ndNJnirfr7uoTDmeDqUuUOCP5
VEYqOeNRDaSV2QcBfZKczltDILUP6gj/V5La3ii0UPE621HjkoZwCOLi2Ub+YnjMvWkjG44Y8Z8X
D9XfZ0p2VWvJDsqqHB1Eu65qY5J0R1WK6xvjNkd38yu926z/IG81xHEevCgy+v4HweiFazFQQuIQ
W2XxtUeNqj8MDM6wV5Btzk4YXPHz4Ta8h8Dgq96ZgsmZX91q/vEN37cLVTiPcu/JUYl0IksVRRzm
fCO/AT/ygDHAP5K6keJEb5VOBSZs56OBEJmH0XKp6snuxnnX8byL9D7Y9xtcQjhGnKbklBg3z/q6
Gfd//hsWJ1kr0CvCljYfO6/oYIMFpWn468WbbUMlRPNY1WYcJ6Tj9rt+X2OXJxYfo8C07nRB2H4Z
c/mkFE2AWSQsa4tbz6vBi/yIGb1ODHnwCWWyMP2z3ASDYAnLdCwouEd0+93liPgOeoCTGzHxfzh9
/i7BAnhntiQCtSyNkViBYdwYOq1Jx3M6WwPgPbCgsqoNQyB3ubVIpp4Yzu+o3CX4/8RbdlMoSaZs
bUkGdlw3JPMsiVVs0tvNkiU9Yk6FrOIT6QacrHVrFD/dRDTncu+jRe4QFT0EHpaiPR7J5+m2uck9
cJROvOwhn/EF5LUehSd8jAMgvAAYtYq2t5kU89YrT9bbOJIPbwapN2XuGeAX8CZ0DC4D2fJODAL4
Do+aNvYfqKUSNmi+Z0avBlIz499wjFm9oMsEl0ULtlzVu06Tb0PdNL018dsUX6mCtU31HluoJNQs
fEkU3c1KTp8FTPdk12msGWm7dwMEEqNO4E5Ha7UMSyNIvpOiy625M7eQXc2BhayfiV663s9x4EQw
Lv+9zUdhVetaGdSWuNKmgzy0C9zI2WkiSUs88+DjLZ354joZLTLz/iFHw55PlkSufl69rIcnyqrE
0dAdyR8azW7fz9A3StP7JWunBmC5EVycsUUX4NOZxIfFzb3tD8Ye36DjKTa1lCj6BcWlGpN+TAJN
XNs8LqFg0x57OHs6hDTf041xbW9dc9e8HtKaRwzNWS707ZWI+R4hOQgYsJAoHB8H1NOgOGh6mooh
byLW+AlkfOw4GbobF1moUP9ykZYHwx9UEuYReyXegwRMHC56slBYHp1OF4Alvt8fZSRQ7rnEf5jq
COAYIlzCvWJx0phan1J/XvXfIsx4exIdqbpbwoxbaRr9vffJ7B6ng0pjGyMLA+tUG2HQuUu3vgJb
ovifFezOO5dq7uMSR4EW0vTLvztBmg/3RFXUMiJ/4y8Qz5v7S64Ly7wlc8vC00zsTCb1VueCaJ0d
ffwTqJWtcVIO4wCbYknzm9RCqVmx6fokmpKM+e/yQTVOQtlaR/0z8d+e8+FQ0WxEp3mqLx3emu9/
jmyVPCQahs9DyLzoMCPqsa65EVL5FpmenFiNsENRc772DeUlVzJ5oFrw5et8dzB8RVWg+W61erQd
19EeAu+J284Ygp8SoPMgTS+51oAqaHW7XFuNtFKl28UEoxVmjav0J8ezXJ8DG1W2EsrUsERBrWlq
k9Gno7TB94pSYyIiMW17ZRPCZsk9WxWiavNGx5V+3yC0yGWRoafQ1CmXkPKEKzWVW6AqhTU+a9aW
5UITDZOG7m278JvTv2w37H/rf4HBEOP1Fb74fKIbRWAGHC4mck+ECN7ZS61yhvkrZ8oQ/EwNZG+L
gE4+joflma5RHhvDafQvcS0ytmFFl1Kmj64S7F8mpbuuYgVmo2khfavcI7gRcXfVZKPs7gTn2Q0w
FfR8JtappzbqgsBQmFtLeEJ/3Unt7cR8xsOM41RZDAtLUSfTkOXrixvQCil+JScsiJIVG7dHZe5t
fAgJhkJooDRRwHKtcOkgBJ4inSAJOBc6CHYyr5zznHa7fZp7GcD628o+lfnaYs6V+c/PiGsvlvjn
6gHZ3YqCMjP2ApgSH66vtiO1dlSzmfjjiQJ8IrK3tVDpfttkWtp2uDDYpe3aZ65KuGxXi+b0nqIQ
ssT/WQd6KTPqHwNQFIgIPBojJ4Mfj+mZVn2Y9KdqjAYrCLyhxrfir1c/HWMdmiO+iphE+sgCQcMD
pWB8RaSalcg3FK229tDEFYxHYOOERTL3I3r/QT2bVfjFtNETZmd9ahA/qEyxZzpqeC6R3+GWMyV3
m8cym75YdQ8RiTLqlfH+VtXVb8rkv/XBv4FaIulJC0UkXWLdmssQDtgIcy0d+p9rGcZHtfBY+bdt
NJ4iC+7cQ/Xw3UAtz+DUYV/pl0vafSJM+Cd9iMfSreWCAso4ChYOCaEvcZbz+QtkIhOf8dRrLg65
QmaN4dHEmxmPQ1omu+Dsgu+ZRQ2aWKyXe0RWHCUBZg6BjUTlhOaD0MpDaoKj6MQT+jgM/AsarTVu
QIcefyIet4NOXRrJorNZuJe4xeK0+BMIwUd4dx47zfcfrb6LbBOwRtBTsRJHgp7rWx9oBO65cYdZ
lQNANfgJn1iFdj9oBDbwaIHBsKrUM8zVAHhbl+WZwSPiCn3X3ZHjBVF4DMckTvSHbYXXzQcW1bKW
2Ev6nkDY3swTh9ilXaOBOgXEX+nIzQCcR9s8boYJtvSRT94p3mISl3lJRQPF+FyK0BI1e0wt2S/S
zlhqfaT0EMv3SBGPedKI+h7kLtKmNXCRcl+42HRxMyQaGvJAzjfdAIRlKdxQIVcFpYpyGCSUK+Bu
5xSHy6nu2IExu3M8VjBpJ0Q9cpjIBSpJV8+MRiUlxVxmZrHMjGKqhcGiA5vw/ys5SGDcKYCb7DGs
llden4gl1c/NmxvCVYWXj6L6ad786RnmHyCyWCnMERIfinDQlPBDqrS7QhWSP19BgvhVwdF924J1
cRMX8UbvmpIskiaDgywxZBfjdjaHskWTLh50fkAzAxBa3Uz0v0N5Ezeotd2ju9fKG0Tjjv1Ajir4
0ViLGfyw8T6UcU3vKjqqAaTWM81x+kKEjb0Tr3ro7+ZsCoPvUMJ+G1wl8MsvHDbsXNIk4jmo9F/E
dyNwEH7l91tJoxqehwk68tjdxIPsZ9/MQeprN+sXwpp++QO+Js0bT/APZKAzCjQ6KvCrwU0dTKID
RgWwZ6NAz96qUTsAaEi4aZGu+430BbJyKzBCeqpNwEaHKJFv/Mbxk9YXuamTiJD5HDCVY44iYAoz
Iu2KEuF8BECc5gHEyGR5Eu8iJKuQ+ToUAFBxyY0MP/vFzNnxEOUj84cE1pT81VShP1D4RvFiLqqf
Iq7eipAu4C5CAKLCSmOGx4Lf4xNECQ5yY99LqawnnCE9qZqo9pRo0K+nlVRuiVdIZYF1TrmSn1wd
bJ239kPPoXTiCNtRKeXsmZTMv3EbgwG4T8lbdcDB01uoj1DS3e2cJ6LbS32qtexjwHY2gE1vDW7+
PHus22hXfuaPsUL71QNGFXICJDV1vx72y/ORtiSICCXJnqcmLPsZGAsP5VRLn+a/xlgB+i4A2nsH
v4KmVrAl2N/chj0drqJFd/VLpfGdwqcZDUswAiMmY5Jtjm2ZUlAAdltGkWI50/JEaBV/X4jzmTyF
IVEbZJzDcvu2zXdMPAB4j0dg8OQAYTQM1d//+AydezV5P39jm+ZrqmREp8TO938EXFI+MCHyek3G
RzyZMoqqsZaJCHvbKFUbTf1D/X7N8m/MEwvOJSPKptlRzoGFsJoVOWfRAFussD5vXJJRB9oCdkow
umVLHkO96tUCfpcOEOxtIMVuODLoCQshgWFoAjgTfKnZZg6W/u4wjeH1qs3/BrPs7aplUVBLMkPK
UDK1HCz1BGr3j0YABTnLAiRE5fmFbCHF0nA3yQIbHjJ41tGY5IPYbBwSNQKJFa9CLxKKysqjNMUU
Gxjxjalyzujaz/YXQZrIfENHid2I3kctIx9APWOR47HVHQudRJU8mS9RH7jyE9K0Jd5zoq+flgGJ
HTNZpZPgBgoQcRp6IylT802sdq3qaYtSmjLpS7J2ygR9t2PRcyFlx383Jpg9zo9MZSXxMol6amDG
19ElHm5IWjjLi02UNcYfZxwAqZAI7bo6ucQRUiD5rEavhk0BqNXzoxadnXsQkkr+wtShUfza9GJW
TiHpvCINnyx6pLQ1yBX3YMkoB3ruLdsX6uY4TdSFSs/OMrVNtMMLImA910bOVtGSxXydWMhc5p8S
1oZu+m5uprWhgecjaOGEDzN6gsMSdMXW33EtlbazX9gE9mFQ61sPw+X4OSU450FVDqVCvKlyXhD3
9QorPV+zSnolY1hC3JikPkXfXwqKzi3jZUECa5DC2JFerKWUh7a/l5oWqCvZulv50ZryeMmlL1oK
xna8YqjA6NepgIq0BJnSqpahWRgY47mV03K+zlXmx+becTs8ivr6rBeCgo+dNFLxBqg+wVH7dT1X
RAYet4Py559OecUCWf4W7A/fSc2BBSYemNP3j/tb6LNpgHbjVtwoE5EJKhmp0jvnEhrpDUOfY55c
nF7JUXLWlCXB5lsuXOO4o4YL7gRx7ivo/nBNtl2dTAhunolQe4O6U/tCUkHRKIPdRORmEz97OOIJ
O4Xfm57yAillMQ8dEotb63lKMOwdyjBpmrjeMiTcSZzNwrVmvBigY0yjnU2rDke1lFXBsubZ0A4I
FgbskLDncHF2ev9QSxsV2LX5IMpMsr7BZOdDap8Z7Dmm8KO9DCXl9gjO99OkJvmvp/NOq0yp5WHr
HSzt3Pcfmec1uq5HCErNv7gEOc2bHI7LrXCSYI86+JjO2Y9Lconoardqhk6t4EdqvTaV1kswajFB
v4s3S9HuvdLpueOohCIxWLhYWAv/JSU+BRP8PwnrFQYa5aMKsQWfbzIo4n9Zofsb7nMTY6UyVfkU
JNHYQVfttlpmFxFrMDMbWhS5Vby9cPzO67rY1Bob+EdX2NdKsHBR+xhtBQ24Pg4VGXB9neL9AcsR
DtyD9I4LbPpUuOTHkK7c586e0sNDt/B+EpsoUFKjhD3P3YmBQ8ofHNPxhLCNQ8vWdX0NCG21w4/i
u1YxZlLum2Db3WQT1Jiu6q5sIecczfj3nKcsl9PRO7zl4JL9/FwhZgAUfZM2DUESfGxLN26TrLoA
4LxMBxs0D8LhELmtIdde9FfnZjHnrnET7BJnpyQFVfydPgSMjKfuWrhR8nTSLRleu6xJAnM27Nmh
ypx3UURzG5O10gfP3VVc+bLIhIhPVLFyPUYVTL1t4g3eHnZOK4Yonk6S9OX/77yoXxLprqf042pi
Lb/vjKcRxoOmtvtgiOIEW90GoNZ4MPLb7wK8jihg+5xTh99pUo180bd5zFlsk/LLhzNJ0knUqpDT
SCfaiT/UHqIZsazxdznntIuAy4SUCuWzw4SLbK8232+cLZha7TDeKCX300xkWTYX7bNt8wmEweUV
HzLS1vp+sC7gI0vvxWI+0QYGp3aJXUR7/2qX/yHoTxB+2Jff46JnKLvvjN/CfBLnaV3aXq+1rfde
5INYUeQv0x+wWo+Pduw8/aIyMuUSRX2kBz5QFYGpgA/+TeVOVl9va4VTMdbTOriAVSeJp5KduBVt
s8tltVlApl0AD12J7Fo0UJO/qP0/kNz9EpBr55xUqD2ysu+t5D9N9SwRsOUDyKzSb2kQklUAChdN
8jZM3b1QLmdQY2ViYAe0Nv67PkYJQ7eFuYVL4/uap7EoMuDaUcecOvtPlFcFuELsgHVRTCOW4kql
Ydb1nS4PCJLW+h8vKxmA4kNUWu8+q4+me6khFOCu5/SHm9xtQQGcxLMy8tSKSNSZm8vX2hpW8Hr3
cBUt2TQnYap8sVyQWaFhWjIOM9Gt9sH86MIwfteX582gM5dJDIoKaUy9N/dySuFMdTTzCM587d1q
onPTVoG+JiOciMSyhAkYkfwffd4FIAzZhYi+f67MC9t+9icx1z2XSEFSvyXW6EUNIzGfsWhPOdca
DWv1DL8HFCfHrCKg5sdwARb+ec8nYPu89syB1CriFml+pNSJCUOUHQ8KGagh0h0YhsSY0c7xuxD3
e203Gko2zAK5p1b5kpdtEUZT45rihoe3semeWwD0v7EH5ga8nlPS4LpGwlWwn028abmEG99KZnX2
XWzIw77+fkHrF3Uap20VtNM0TVB2Ly/lFjU8C1mDL/g5vaJ0eIWibEMIZT9mncIGhw19SLL7Mroa
lxKVOgcCg8cFxunENIN+49G9fb9iva517N+jnHx/+yDhYsHPP0BHPKSUnC9wMhcUoe7wv5fwgCQD
28QHyNAT+83i1U0ulhWR4Z/4tlWD1p/kmZeWnvgtV4RR7tYl8Bo9tmLTovGj3OR+9IjCXusqUsun
raex+0Jw2mS84dmnoKAfzLQfIY1+15ANDbe0MgaZ7iaADCqgDiyYp2gT4s31Ui2gFkXXIstFUVxS
byUgKzNmGJPgh+5C7RPqZMW15uiPyO7+tQ/C1HSsleRFXc9Z5VR83Z8/zCRJ2rlhCJCT9LmxFDpK
LL58G1bVuCRG4JCc6Y6+6kgxDeGNMt9n4z2QlR0kCT0xX1AR0QVs1fmWoQ7FT0K0+PV4xftpPgIC
Vhjfv5PCsn8O/DNIqB2NPXJYFGSck8dL8EyeFQkkn3rEXAVknaFGLjqgbGhx0TE5IB8rwu/Goo7t
NsYKgF3mZp88rjcMzP7RRXD9Rtt0Ftf7Bz1LsmiqVN8wOSew01FNyZcXBQfZlkmnFqgnArIoLCXE
+KdrhWfuhuCN7jcXFr7tzFpR+vBDG75IF0KsP8SeiwlY2MQrMJwRHYe4uZZW45BMxOy8mxvSK7N8
Qv+rWiyVJ2Dzn/4Ueyj/AcikMuNEVPZWQ4KRbZeoKO9bdWoCaQoSvOIC3lVyu1yzDysBWNV0wbk5
sCYd0orC+YlCgOKW68a2lCspA5QKg6mxDPQsAsb7Xgh1Fjx2bef02+DHkthq1UqZoJc7L351w1qS
liW/X+3nKgEUxaz2YH9KC4Dw9iqp36pZnh2Bmxi/r0Amf9nvN8WTTqpbqQHxe18D9yQgvHhtb7XR
vcr6R1orHyuASQeUlZ3BMepIh8W+rJ+v0rqwSRqxZ8309TQ4EVu2mL0+PcVbAkkdODRe0uF4JeVT
z3CqPSxipc6DUzRjmmWzZGe4nWlcObvoPxIidxGgG51D2Mp+t4UzgbJSlr6bZcFiMh9x+qAholkD
14JvD9EACAgpr0CKWeaAQXCl3z5dmGC45wgHnJU/rE8CNYcwUAACw/yO2VZUtc4XCXvHOtHFJA+/
VqPgHlnaZn5hj4L/fDJ+bhmKJSPXYLdiNwxvbboYZ+OTXqZqY/zP9MyadNN5naWItJYhVv1m5pkX
7ueIfMVWr4HQ0fgSnS6q76Mc/k/Lkwx+wfqwqZR2b7miSpKUg/QlduD/R7a+lgKMhc2Iv9jkZzRO
U65NFifPFlaejHC8pqTYhI4jY9AWIuYH8ETDqRClL/7P1RBvE00MeCpLUkAqZ0COLqJKGYI7eUV5
9LAray9sz7e9Qphz0JwjWiVg5Z0PyrVH/GQKvcNX5MqmFRLPaKzKf5wtOqGCm5snMtoBqhYj9ppb
vgyoADSZPPtNQBfkx0zgKS0Uynf2POwu49FcyHt7hOWp5myOEMQrwVQi8btuNg3sYZFKe5h8bY6F
0ePmH7vYqbWVXpHXORCjslhZtUxIJ0njE2gDzGsfDonm+OkcvV7Pte8JZLASc273Qs3zFZmMldih
2vM1661RVuz01VAOoPfxL4GkXf99p3te3O2MzzN6vylQJBy8XtmL8kmnTHrHZN1sbFLQGL0DBBO4
MFk4/1WGC2pEqJSdOQiSD4ZtCFiewbS/ySoPRV/jbZ4yR2XpOj5a0wPHTOFkloDwXV0YJPJjviQc
ONzWr8+6PGp0FToX7oJwS6v4fxE/FS/beZCwRSyLlzfkDfA97nHv9/GVMRCpUASxGxCuhjFLvSTv
SS8r8uVpeZ73rkgaHXNj2Vg+aAnnqLKk0PQOEgJPFOPpptLBe2qRgisOfMWfnVIFihDBfDQMiDdz
oNP4WobEOOkQ7e3AqRW8YfkFJ+04lix47Mjyf5U62iCw2XTufDdzNQo4ZBPkhxgc9Jn6t3xl4HIY
vmY9kA+k9x9ZxDm6arRinY7XCqsiKEVHhGM/cvrnuhvokxzyiB1ULHDGlc2el+XE90s2n93/fWCN
eoezawOj3N8gL/GYK4NFnboHRa1qLgrKiF5+AYJi4DkFcNlcgsEMUYfxyh+2TsHdepxzPamHSVN6
iQVC0BeA2g/ZWA85LU5wY1YlxJj2F59TK/MAZclAs6QOEieKahuNZLR3Pda2kd8lnw76AgTp2/B3
alHVS5lHCPejOYRvRh4QkldlOjD3AyoffNWonfLo8/VFsEoi2B22QUNattQOJCN2XWtlQxvAdr5z
0uptHTSdELOQyfODzZuKo7O5B6r+f9+b2XQHyXtIGedXdjbE8Nr129D7Hhq7ptOJtifJ/lWMMMA0
2RbzuOevFSkKsLQHEXHC0zFPmsETFvP2wnFpIhqbx9cem2tKMUYVsDmZsQVpiwDwSOU4jvv/Mbod
TA4SeSQNcUx3brSH9buwGFK/+I/H0I9Sz1RrD2MCqQEJaTF0yhx/IFWD9WKfNYxDL2bvl1tM0SOn
9XNrvPNiXG7rbWJXWH+hFL3yqwf5mez59q9LPnTmmA/uWK1SfWT0Hm6FalNp1LeRhJDT8E8Lm3BA
LTU/piB2rBIDJDF594h1Ocj31N4iPLiFO21jeStaw+BM+TUWpQaVcN14LeOZ2L95QAXlkATbObx7
077yKQ3mrSFOyD6/Ql+Gyq6Iz/qvcv0C1TTSb+CIdvOWocy8enHAL1Qoev6D+WRrYD/0iC+bhL0u
8kNOe1jkx2O9b6LVpq7ShSYgqksYaQSblkUbiq6pM1+yISIFUZ1ZrLLhsOpGACJt/+IZdJd6K1Tm
7cLrw1Q6WISgFMvWHc0aLsdlHoIJDW8G6ZH1AtQDCXSfEVG0+KyDtqY5anavVFLVy4/YBStqVRiY
am9zxXKpvd2Vw95epLGozd5ghDpw3G6q9gs4nB6U/2Jns4nbGzpx+BwSZiB6DXJR/Bi82SV+BIir
tPsfWLcHc6FJOQNGFVY1QJXUF2Ply6k/dn16qFbR/EmS8fP1fCRqzoWI905M96cKgJ1DTa3awXJt
lQqg1R6Avf4TF1v1jO4ky+IYqUYoEaiub//BR4rPmFrHcx2Plh7q7xKhMoPJeji4RUjqTGp5VA/T
kqw8oOMjkhi3i7s8sMPLNpDWvLjtEUZEBsGH3cMCeyLz34+O5ulfSqThzFy/aKBr9yxQw6s59hgy
iny1yS2sO3wHoUjMo0KN/Y8J5DJPlnXxSV7hcZCGk05DeUjyHxOp9XJGJuyHEc2EhB/dSFgPMPoY
mPfZhVuEnXAL6RDjahJ3AWYjamJzCFdxk+wnNav1gkY8qxlpFhPajtYqNzRUmd4e1pVHjU3nEMa0
8+AipICPjYHcNqjmz69CnWYRBoOPM5L3ipyfWrorjAhSJ27QGbDq/b0qxEuFMr8EN9iVVFKQY52z
5H1q5ySIURBdcg3Vc3cHa5Yc7ietoVxLANyXqJRmG5GE3Cu0yyC6IOoKNb94NMSzkrWkjuCFeSyC
S13rV+PEDcknDzWDqJe/H3pyz46gBfk0LZLsn12BQ8abhDVVl/kbdBX0dAzhefMQAHAiJdqPJZ4d
+8f62ohwqnLSwBOAHxjvwNCgztPX3Lc5svNLgQ4DRQAMbyupp2DBgmTSThlsxk2QBah0WBs6Y7r8
PX1IzrRukz/Jy7TeuOWHeWzprOruPxhV1GIxFfSDxXRk94r5NyQ0czUrO3No6owPIgPHeYsvbn0p
AfeQvUlJNmvqRrIo+4VcqHK9BdA4M9eNfRaLiZYQz6avshTobBHG5JgqIRX/SCu0UcGiHJOizlJh
crpXGKWH6V6V9dJPISw6ZdwmDnrCZ57/5fMc1kUifpB9L5ov3Xas9a7L0oM1Z+soZgeMBOO7k7iH
tNLj8mvLW9XexTW6xwWqv0KhxYnQYw3gjl5x58n7kTHYeZ3MVRdWnUaIQD68UExjti+nUhAlCFnL
abb6PcnsIrJZvbVVVW1Tdq31oMagGElgmvCiA4YTVDov6pjerk6WjyAuh7NftFm9D3Kn86MxhkHp
AfkgCfPapVvmC9H+J3SlmC3oNHd9Uhjm9IHNhjaqN6e3/nHBx4cOPaldJlxT0OLZc3yITCDx6WIz
uGH1XDWUki9+XewVFNtpCCseRtGuPvEDXv/M4jz420mwFgxF4XCblHm1ikEOhy4zT83cheJVQtEO
NPMKw4NjOfNvprDo7k/lWI1BFXi43NQYppNuL2MEXQLUwt6CBUfBKy8zSXIKGcV0dtTfD8e9skgm
jy4IEE9DnMQvC9seoxN3+0ePmano4aJ2W09M9HTGMx0VJLiDusNQiWV71YB/JK65rW9DyapVQAeU
W0XARppJ9fi0JLTMvebsc6Ff68cYnCHRg0Tmk3NcvrC43kxDDkkbe5R3Y3I3tqIR2JGsedkkJLLw
+OQFCCmkhBXXR2AWSctWhZp5W4xFXYe1fvKBac9x7UPyO6LZ+QmO7pHKKPHGXubrwbVRvVz2r0Y5
jFDZJv4lYVSiltq7NN0uINv3Zg2In5zoKqJv9joxLK2Sn+49Dqk+G/h11i0kfJ+E5bzhSmsZF5/S
EEYw/Fa5jsjPPkcIQLweJXtpq/W3epseceqqMX+HqnL2mOVCbOahNmilZ3GoQHy0Pg+WgZyHwW1A
C2GpHujKkMhhI2SZHygX2ylnazeT8qbHElwIMpVVexOMO4aKG9B+xDrYSN8ya+5clCgv3M2FNsYA
2edmqLL00nnlv7yBlpkEn83n9ydSN8J+XrYtEsMtOg3T8yt3musF/ayDXW7sCK0XpAdy6YqKOmyD
z/p69ysLNnPOvtFzeZF6lHn3HVffj+wCIP2Nus1J2Drz/NQ51NCL0Z3HGrkbW5HmlXRY/6reDOGR
PKQzVPo/JmEQWfaKwd3YWgIN6s0tD73LKygbB97PapzkwscrLAk6bAzPtjtuzbjRUDHiYovWul3k
XqJ5tPIdv4Ef+wGSDShLFgf/RUFvRqXoMbCI/9vzyscos5jIkmCOcVuCZ8aGXxdxiPFv4sByiVdY
4R7B1XguKnmSbm6Mut5Tl53xnPnxMccVVzi4HpAfb27AyLfdiPDQd8XZH5xCoTiZN+VYisyJbF37
5OwCynN4JU0U3Ur93R2OcXZaZI8+DUHqdtWE+opYxmKvqZlr63yCjyQi6cinz/TRyDYrZT1l59xL
Lbhn/zNUW+XUgXBaSniGRCqNdWTs3/SAcs0H+/QYuTNXVRsaDW+kf8F5eYWg/VR8EnBap3U3lgeQ
PxdyNv0KjVMuOqkuZb5evMs2JoulYe7iHw/bMTrUlqC6KTMueuPImsikMHa3xRqS/1YNhRJoTR1k
DAEHzgrzymKfFN9/iWfMQBud/2GUT5tjd0ZK1YjqhSuHUU3knsa4o5wE/ojRbMhqviaVZjgvkQFO
PypBRtvDQ/gRvjZQzqkh6mOxtazxbouOP5ia7/ZlwU2MOXZUyPS5CdOMVHHeNBYDGzlUXZMVHBtN
7fTBoHwpcxqAzTQkwVEReUZC83uT3IRdm+qAeUhyZ2jxpscVgcgf9Srxv6R9dnroTDXPNKExssdF
WnNNbchgsLU3FO7zu3df9y24tFmTXcO2A8iqxA4sJHT6j8QMpX39OPBYqi/VabKRIbKCGbNPCNGT
TThb7tGsKuC8PxwZctQ/aDYB44uMVrs36lMyZ9p0RZ2f8OLI4Kjd7rbO3tb5z+vuTdGr0AiqdAUC
ObQijyOMNWEHXD0IMjwmst1wrogBlqPBuzbke/iLG8MNokOfcaugGencsAUTf9hjnqAZJ8mh69cy
YUdE1tW7vpt+S2LKQKBXfzTNrJIWbbwJf9MJcDBJ8r7Yn/cdxWYdCBoqYWJwJfBOihlWzIr5j5uG
lXs8BV+0NrBVwInl+9rve9X7GHWaK8kfqnX8XWK8ildVRfFmMVhtZ8i9GUVK7UjYt8u0Ry4PoilL
gU0MYOF3pc94BfHZzW/BvtHSZPz2+88WYA1KsDS8lJ7Izh3UsHvwuJRZYt2pnnmceSSvoenUaEsz
zGJb7HozQi+Wb3wydOLeKbNeRZDATc+rgkuhCl/6v0uxjQmId66TVBKf+ncJgszWFRijSSDQQVpx
z95VLLam6EG30vcQ9APTd595dhbZh5Q86qdi4eHgns6LN+Nf5VE3X2hsxOw0NK3llS23tQbmOw4r
v2Jx0Z9DOKdVDMSSTpYXGV9ShPP2okRpEaOtal/fBIQbH61lmGvtP43HMsuKSjhNcMzmJ/gz7qaK
kCpsFbgxcLa4SSuKQmDUeKBvmTh9qE5mhmYg4qK78C0xAlmDhWiLKxSG+SpWw3tpkUMGNECQ8FYK
kpjdL1XxwVK7s/k9JLqJPTpslFo/LeRtnFsWXZ1nLbr46JgrmwVy0W8pgvf4VTcUvjOfpB3Q8GBX
pQGPXT91Iehjb64BkoRrRPwo04SYnOTzWutFlsybbEc4ns3IkeC+PddTOW6LzccPbyNOBqvlhZr7
Zve8QG86wfYOKCi6FX5wv7zSglTNUR0ToBBlwSdshK9tQClnsuSDwx4844uadsP7jG7Belo8XAWA
fI9E6gKrC4owfpzk3OYEXEwhftCouaajInMxveh/tk5OTeTySlh5QEzg2wS3dy/6PrTNqBJt3rvn
cJwtlLRROEML96w6nDeGieIy+SVAw+zU/E8xdqR5eTarP5LiPC9piNmNTiFZhUqtim9PLfc8EWQ/
ewl5Iiek9Y5k3EbVrc4deP0+KzvhRsDCtT9TVAypMK5tEAC/gpHmD+Jyw6hRRVAhKdAvVPrIr659
OaCUET1X+54O0K1wN4XEw+Z7+59Ipuh+Zjn1MgKphwsAihqIXHhuM7M6jdDh234VSTFMH0TAnBGg
l7oARBVGrXHYhjkZgm5ICu73+3KVm6LkFQUPIuNKyI8wG75jD0ljXNsh6uiTKPQ864g2rgpov1Vg
QQinUtKKoTvEP1/uAwuK++jm3DU9w4MxBZUVI8JKlY3Tp0hUFEDcaJ/Nrdcu37UwKY/INmOkKZD0
eFCFi7L1lzQZWtTOgOPUMvhNPKxN10ABL9/PVvz458H3PFJSonsPXDZadQokqsSscYY8CZlUugzG
W0wPs3J8gthVu6GE27r6N0Hk0Azhpr0qm7xyAyP0dYJKvD8d37kzjOPJG756aGfBbT19bYY9BGVe
LaoQARKJ8clenMj3g3iT/CMy35a9oMx/1kkZLPsHTLW2K4GCTIlPHOB5wu3nhGoMFOcp/IVWvHI7
l1sN2om/eq69leNwRA0Y03bG97IRY+tfzzQJnBdNSQLy54HF7Ypg20skAHwbDNDz/vyPeVPWqgGe
dvA5N7HRtYyq3kAdtMqA76F1qnSiU+7aAQqGDM+kn6BSenhNR2bRVWOr6VMy4+X8j2XjVVt7deyS
RHqbX2zVrN3kUJNt/H0X6vtqHd92eLn5l7d0K7B8tppL/b7smou5Gd+ljkezOzmDj8GUoGnXIVyu
0hTiJUuD7nvDXjnn64W+hrIMm5jMr3p1FFmdJSTP8riK8O2JTbNZ9ZunkUhXeBoUczp/J3n6O7ww
CuB6bHyuWnEKvf4Xx0u/DBUWReBIjD+Bb781dYgH055QwduMsPWiXYozp2UAE0PKW3NTkgmfgcVv
sDAdgyZUeZFEw3bWi441yln/U7spvFpxRBj4/9nchIq0dLiMbxbU9NeUjUGZYVNsTnsF8d/NPNze
G3ZIe6P+7/xiLRS74o2FckgtN6lPrpFyME9YrA+7S4QSEIK7jvYBmBya71lp7lFQvEfyeHbX87Ir
wEtvpLtb+gS6CRqMqaV9H2GXpuRvOgXleuU9iqv91y3JQskduJTuP10QKqhx8B6EBJMZyaP6/0MN
btmc/n7dpkRQzpOcDXji6ieD1FRozA6AjGr2RPET50yUK8I5HwhXRLD4aomDtTyE6D1AmlBfXCFr
it1L+KnwRPXwji0VFbYlxDZ7tL8BqmsUgykrQ7yRFxuzlk5DYpmxySAkQsUraxBhiQ74clU33/FS
u3j+1wEIjIK63Gk1o/PZyIaooIAnnMvmn48RPTfwfJxoYQTwAGViAuTO05JLfiiukRY0XlY3lbg/
HlTjN8ut9WIWfe/LINfZsISeEHRcg1gccMjU7fvJO9wbOrnmWUFoIAPermMrIj/gLknUDUw6C6XL
hyMWgt4RQlnVzoZp1RN110bhljB9G14NSCCmyhK3XxBn86QdKOSXIfnNQaGxqvNCUjeKrav7g4V9
zNJ9wngBwt9+h7FA83G5R5oqa0YqO376J3KAzgrDN+7y2bs+jn7c9Wm/eMNYr7SHhprTjEvKIGx7
WQUfpn7NsWaClok1/euQHHY+40HxORV2D1LixyQ8RChtCrpKN+4WADa/11ABAtzs8tfQQQhmRIJb
fRh5vlEBkbywVplyvMZgi2qC+4wNPb6xNk4478g3Vc6F3osRtjh0HU5Z5DYEOnXFQG20No/kGqns
IZ5/H0dqiK0YWbivMDVzwYR8uDSS9wiAMyF/rNYlz0Rq3B0vHi6wREefzU0BoGIV+tjJJMugPlBm
zOnzMaB7CMgeguIU02V/DdpvWjvKgNqQXd8z3R19Pdfpr/Ycvv6LmSyOJvxVqHAlF2mS8K84fn61
4qX7YV9OyauWZ6REvpgsDuHVzUZfUOzpZ0wFsVu3MVT839fzM5VLJCmfJuqfqKU3KgCCNvuiMxJU
+yxsr+W/uijbQ1EbdG2BmSOf9eKgcWAOrG7j93h35OtU9iFAbU8VxGExNZwAzxEDKjCgNUiH9ywI
IbsvZEty24KxWASmEOuff7E/TkiI/e6wBOhhziVKfEazDfxskaSH97RXw6pedua/IF+SwDU5OSyR
zdeK2s4tP1eNbLB90auz9MA9iYbChvS6C/254bu4oEsM574af4OvI577LtUdWizuio3wQLMSFNhy
Rq1ZtiYb+8UkbaxbLPGeGIDdKYcwnpHcWcSkdN4leNy0HOhshvNrxb4F9ByXFWAuID17HJLtLtcC
pVF0RWo93EwmxoRHLi7mL6r2f2MQviUVz0rC5YfAe0D257BTHCKGYWXV61xLqSw5hI+L6O/W3Dwh
GaYLCljTFTU2JJ/J/6hGJ1WTuIUeEGhkD4/pcVl0HFLeD4PyBgX/1AZpt22Hy+DA9w8+kpMZo20F
nJyhlH1ySFnTKHcSPVDS56m7llyYbFvjP1m1wJbAiT3I67gqLfuiOVf6G+6QJkPeiuZz/ItioYhE
6xixMlddyO/9E3L1jZdEoS3oaSPzC/GHZSAlaheUA+lpfJ135P7msU61G879hrNYeyB7fHwIVZQB
4ExHzTHmmx6/T+IeRKA+f7PfIXLEJp8I4b48Uf7H9ZBjUevmVcqY57fD1DOPSWYb0PVtOI0jVDog
u7P2OjTZ91/LBTIXb56Gri91gzsr1iLU+8fEA3iSEd3asfFHiMAHP2w0Z3ikLvjuZ4yLvIczbaSV
os5OJ+5wqsgjuxfxNaIPbVNL+nvrIbzkgKKLHLWYFQXY8fTYz6wsMME8Upy7BvPUs24OXEZXeq7h
nNnsa+xI68tUU6RNOhdTNLYoLb+sk6OVTk1gGXW6nJ/e09PuOzgX7x1T8hWHMj9mek6bbsegSiPO
cD7C+oBBfayrqkc/pnuTShoIGd1HbS1nzNDhsxs78ZVYcUS7+EImtNSiA1G8BDjNZO6gy1dKZKIx
l61dZ0hVBsRjOQNzTbZberHC0R7tMF9tJw/6BW1UczEyAwzF64odiNcholtAfABtcTyQf6+iyMQW
4NGv2rV36QdCvfmKwF9KEMeO5FsrukudUo46jslohLvSzDDqAyT6kCFmBhEVuMePKztthTBqU3ba
yMjzsYwq6lYN6GK09EJz3CbBiu2C384vUIjohlrgobetnnSnb36Pdoa7zos1HdgJP/0Dk7lIR3oY
UFQE4rtWiJpFTT+DU/jzPygK5bApOpdutepTzvSJHOS+U98xBpjUEOyZg74kJtw3VEyZobzvJuoo
SFXRzFdjtLOM741KRWnna8WTopsLeOnryP5XkOj+rsbe0d9FzTJumUEClaOIKTtZ6s5liu9xmph/
zD60xpXOiE04T+olCX+3Fe5PIrkbihM24qe+Rdw336/b1S55PkJifkNp+A8t9VHY+Fb5+gTGm1dN
J7hDI3/QgYL8OpDpwrJ7uQ20gEGg+JQIeoOnjUi+QU2uC8DlAecGfeW7t9t5nuPPKlUMr3/NibDb
A63T0roDxxQHxjw13+/5XcpTdG2JWngsCAp8zvi4LCcg9angcMjzNyGZkGVhtUClNF2/wNFZKsrO
P5hRIZ7qANnEOOlz4vTy255DVaAlJlTg0SoiXBjLbycttCSCscSI/n89FY+J+g5JcZCqAxBVBY6M
R8Vezns+D3aF9nTc5eXod/mPplxXBkS+EjPrut4Y7ZojTUT6mhp/1dfOgPDGYOajmfiCRwncw+Se
zsA+lcVf5VH98Xn0HDlfl4jnzmJSFz8QU5n/B8Q5zKuL9l722HHvqXZhw7baJID7lvgilbxKskun
22LlaAbcuiXUZR1fDk+Drz4Cu/Kn3STjmomr6rU8HPy2wVxEsYqtBaC8KxGCr6kQMG6X5wOeuxH1
sCHl+Sxb7LNG27KAaGaKnzAgj83QnHohczcwMPQ5xweYvta5pJ41yVJPkluGD7iOcNJHInm/10ib
Iik26+3sp6kCYjIresKIbLSjQa6p9pRWZ++pNFFDTkGNRDELGB5Bei3j9Zr+lTTBN8CEKsIXZomx
uZLp+VjqaBMmjS21vHchAnaX+bh9Qkcn/nczF1VoJWhmLhkP6a8kDqK1zK+FAcc0bNK+AZbG9gZT
YKiGzYR7Rc/JQBVdZjwxWw4Hx6p7LWND1JqTBljLWLY3/G0M6trX32rjqCHS/H6NyaSvQ//n+EQA
Cui7WbkYa+spDsfu2HUl0lZCK17EjFEbW2UVh7WjwfHBGwMOnHe+hiDlCH9zIjchKjNPFX9+UE7A
j20lkyTx2Rg4I+7UrLJVs5IjAZVf/4V+0FMNmisUnCQ4TXvIRhzD8PHISDQBXKnYpmRylkSLca+D
6fjMcdKLh6hKUZ+nsWBLJMHLZu7MsmlYHablHt6xVUMr2snryM5lEwnIMAMCksiS65YgHPwah+ih
ZZIcbwwFIBUH9uTjDxHs/UE3gcJpbVRDMTquSyaKyHOD4wa/0OD26LwLq7u3XPkMe2Corq6701Eb
swl/SHVIyB3HpejtSt/2AY8rUhUOhNc5AppEf+WfXIWtqF5CajgSN9fMbWHW9pHIwYQDlaHU61og
juNo6XuKRNbqGLVznrTfVz5wpmjGNERLFP7U0cI0VMP1tI3kY+arj96h+JC7DJWgoSohRZJDQ0TM
n44YX0kzJv67czoW5HSHClW+xQ25qaVL+v0jOPpfiiMr4S52Hjm146XS2NEeIWYsHoHEN5rtOm/s
z2isuf6eEGIdjlHYF8tbBGr/VIXT8m6HsYT+UYZgqZJyRsU55kffOLHwHEAt8dfwL7bjYWWX3qGZ
ypZ0ZMnbNTsziKmVe/zw9+u+b0Gq3ihEhOQi7+tZ1fG1fn9q6hNsK7OKz5ffGvHELDBfGFBm2Chs
EQhQoOpagfGstbHbR6lavm2ooKlh3oxPPmO4/w6vjErIE8jpj8WTotAQ61yoLXkakvLeKSwjfd1x
oOCfAiPL5Lx3J+lfXtp1cHdh24oz3RUVpm26gHGhZInM+Ig396GIFle5HdmYiEq8kEcddk0o1Vja
xSr/482jEt0fUubS0MhVvXCzciwH2ufjaBrMi390VrpxgnQoeeSgLHTRdTo0O4mdi9aguVXaaorC
agmQWAd6WgVE/ZbM48q5jEzLTMAVVtwBWaX1CL3jMWhHTMfT+jhKFo34PcwMfUJ5u93AcmpZmvWb
bPIeaiCo8q31iCTTjYexZ/Bx65+9YSYpXDEeg4xk9wV8RvjwzNiNM1d9q/fdtYmX8noG2t311lYm
4MI3aSpGya4vPowFfp+yqZ1KGG/CAiiU+D2uSfDalf5Vqg6bSVRgTm/R+nfrqzzKPPIGVPYNBCKp
Ti0QuHO32u4+Wx7fPUbXIBm6p7jkgHswdHRLGPEpo4wY7t9KqPgR/nVn8OGBNQ75Y6IhQ83Lq2Hx
zFIf8su5DsgwUv/jZqp03y1WscHheZS358qtR03AdwGXhZptF+Pb7ruHEJ2sFv26qwySdhWYF/EB
tF5IPchmwedcOGvppBsTEtytg/7qX46fQIfMSkFt1gsdBE+LPm0kjLhpVzcAB6SxTCS/2KVAgR/J
P2Y3EbURx3ZVwibG1VVK0rfSoD/f3WjiBWAJ1LQ9CBH3IuYuvD589a1LEKJu82p7zh8YmgV2s9DX
Q9m7bKr/XhQhgH05pTfYVM3y7x5uANORNJJjom0THkzdMZrXHcu4zToXrZaO10iNTDE5QlWr/KQh
fnT1ABHeixe0MmXiY7Rhu3vY8h0u7fHjRbPU84huzobcJLOm/hiTpmBxD2GciSWtKkNaa8OrWaqk
tmAwCDF/a/L6IccjbS0a7f3k6cQ0O1zSBzOQcJ+pqsNEC8Vr3LWa7+XUmhKonDtQZ+7SgIpXAjCZ
fpsSpnH1U1vyUZ1wa39fADGw1Lz/W7Std5R2lt4S7N1gwP+bQmM54E5b9GD5cYNtk/Hq9m33AbCQ
+PUzgi8MyQmRaJc3q5p4U1aMjd9wKFKmEE652JPUGO74QuU66/leYeso+ZlrCmjMQbbsWCTfX5hm
56ET053Dh7/hQ3meHHBP85JOoG2GtfL7SgMyYbj98Mw9EtNmpWD85RMM4tFWU1PGdcV5T/uVLtfr
njGNfm9h4+X+aIR2qB/UxCdjbV/Fo2iK3jFNmJwMu21h0DTJw6O7taPdOiNHmcJ/CSeIiyoukitk
w5+PDCFQF6/t95gBKiuZTF1Yeg3hX6Q8HawKw5HHS/2NWleYljOuuBn9BaFxHOossOjP4S5wVKAC
aBkuAiJNKgKhIIcXq/WNt8TRx7SzQVHVwip7m8nzJTEhFYsMiIoWIQibQGdxwT1PcBOUqwF9qprf
KEcN06i7Ry5aSX3pspQrSgUGDXbO4UmmREcDoxS9XswdzPNrAFNk9C4Y7WBTRJCKEVcE210yDXZk
4wCdzANeOAfTynjnKXAE9z8/5llyu+P+jc924odjYP3frwH+/tll/RFyuz7N+Ke8ngTjtKmd72hW
jfUqDzo/WOXjtwgTHFkF1HVIib5aR/w93VLOu8OJzSzgbja3Vk5w0b0iFymHkx4NwolXSxVDWIIW
OXsgKq9Cg2+Hqpo+VbKXCFOQmbmbqwt5JyTVEAalFwP+fPDPKLnaDVaM2dCRdUxVFFXwij0Q3T3z
CjXYUpEBfVJjXjKbyCUKt+jwclOy5HyVNk57n9Hu3taq2lbFVF3VtxIaJlTUle6vcCjAL5IbtkBl
fnWgHfcT4blwm4Ayum36YOdXmR4NSZD4AdVIHxR9WWIQIyIq63sLwuRGjpkGcd93miNyFeumKR7k
d99jzVXZWnGBC8WBZGeQWmJ+fqYZD1PmLKTD4GYr+RH3jyT95NA7xUp76uA8eYNbvsAAs6/7tFY/
L/D29dn/Gvai3Bg1YUbO76l2NMD+0nIMq8JqOq6hiHUfHcfu9YwpVRaz5uOqBj0GBGg1LFPOxDgq
T78+ffzY5pCpRrqzTfzfoXeVJkjlOwyrFo7OUHzv6nTYg36QMRiwpTqBb97LewpaJhdaL7nPNA+L
VA9m5syaFDMErbmNXZ1/ENjSmaF6VibTAoTCX4ticCytwBSmfYSgyK38DmstyW+7eoLmLOl9BMJa
5je7M682zlHzqv4fgEUE55uNHghyYJZ5hwxUXOR9cApGAXHmxPVqF7HeqZQwisN2yeArp2+T9fJU
xX6BDOgp9zO+rTJxIeFJ2gmo2WDfjMfk1VbG8bmeZqtu+Yrw4WAABUZwt5MYFeBVVki8ta9U20uG
7X6rNIvfczNcy88+9LojcG8jNheqRC3RL+Ft/dbFL2XD3oWZW99OGT7qzdDiCz5zhC4w5ez2GTYu
sTMc88VFUdcnrU++nfvmKp1KjxAvQTYMybXBpR5V4lwk2KgXm0XMMrJSdsyxT7A7tpEPnDCejVeK
2l9gwQd3xwpsbF+Lno7/5UveAayT8YDEd408FmNnhSk1qCkXjuVaF1NBxOrLGvu1pH5z5MoIt4b+
GgrlU7fl1IZnVG0NWPVhZ/aH5v+TlWPEvCwfEgIjBo89NhxTFeIEg6t+Gxcsla+uGi4LqsUSC+LG
5wsU7xIg59rkaZZwzZ/Exrb6YXaw1Vku39kzTmuZ2AxjE6tWtQ9YIs74amrSwwHRO2EO6cq75TW0
fXFvU6Na23fkL2CJAkhhYDu33Uf9ep2Ni1WrEi5a9UQK4GqSN8TzmcsNwbaJGcRpr7BFWE++ulqr
wyhiEDgvll1idf4XXpilv43HJTMKG8On4zR0ZXIbQ+jbp8xt7E0Of8xk5JFlss6rC2BfQBVHcaKD
J3Bh70q2SQlh/nEgfvzsS7pLfSHOQWsYBjqYiUbhsxK1A0Srq2q5Bq8nw7On9hHkdv6EQU5BdMNB
OmnpY9Ih6UzcyEBH8utnJAT3TiqT1GQxgPrye3u/nxvhCCtR/nE+rI514d9PTY0mcDQvp+x5VklQ
ilnwO3tg52uslhna3WDmeVujK2hzryoB0wEIgp8UEvhTpOV1BH+rgkdK6fTFPGUZn5Gd6hJagwHo
YksS/C24LNpw2doKBv5D0kTHqmONcqtjqdUGMlCemeTqSCzcmU8e55r1D/zSnb05w3vYgrzSN+Xo
LzcwtdHjJMKgeDuechfr193nSOzJiay6+QqJirebBwgazZv79bW4hXKUl3+KvEgKdkORUlO6n3m7
b33yMOn6UY9glJ4XkBKC0N5ffkjfFXMOQZglEY9mW96RObv0lCFuahLCLgwFNT0e3fWLZ0nRcwhN
TIiZhLQ+L1BQciJ3Krm2c3k6TRLdAiTwIe2yDXNdZ+u88kFx3Y+1yQDQKLpeOzKBwzOH528QVVn1
OvZEcx7tk+8Tb+Jz0nxLfcnyI9eoxeC2hJLlqpU/hj/40qZO+DpODWb7iRd2oAmK5XbqWTQ6T7Pg
dyzaO5jHgNjQN1qCdBX4IsQBQLFJOaZe9bDME+gobn2F0szuLVNUR3XzcV13z6HNTfn+07iP6OKB
KAr95Q1x/bNhYDxyv8nW0iw0NX30mwySco1Ofywk8fvuq234VHpM+SLyU+X2LDGOv6/a502+IhM1
RbDmdMJR5PPAilSvm3aqCtY6tKenVIJgmJON9V3ObIh860yY+o3yvCtSxebUo3z0zr9yh294gz38
//0b7bTGXBGIb0VkwAzF2FvaAvr6iyKkOVhPRU8NZPOTmTP0zXVQcrPjvYXQzvFHTzKxtAi7BKrZ
R5TArT0zpOHgJQRWllIIMTWlh4MnaOtxXe1lviRlft3WaeBDa4K5xZlMvT3zjc9LH3QAhX0PAQVM
ti+gf4AE4uQNSkLrVqqbWvb6N34Rk86uxQZ4pghoNvsIIEOSdawp5zuGVgV+9+1/9nMDj1GtRDTG
hDY9G+ZspUWFHbqTBCPx4wIMu2aQsPFL+LyXxsemRC5UlSbiyO2hVDa2Kh6lSONgpTigyuXC9rgk
vnsKKH7b5yBldhfdevA/pfzk/vHmA7VyB/aaJ1Q5uFG9bxytwdXDwlPpdakDAzvNtuG36sCpgct8
UhOn6c3z8ustaDSsOcOtJfnrPRMDXLTw6UjAuoJeTjG5t7nfivLON6qZiDLyhSAd3pCp6JGlnsFr
LJ5NN3OxYBitSU45tBpdXY6yGVZWBSlClaRm2Pel8VXNF+kvjECiottDCAAM4Xt8A4ksc4/2r1rl
jXu3XNUz6VoHUU0J47uCUffkdj/kNKjlWPfflQ9GoILxTlJsr1ixCGd/kL2YS85PThWxb/GSl8Um
TtP4QmsTPwd9W96UvHCuSqcQSiGtHftvY3kq9nyNrDXKwfKOOO3wGWeS1Ybh3rjKM3moGGQAe44V
LB0rEFQIbQZxs6rivWMX2A/yXq1hVqS0aAEV2rNlCyIsePT8EF6pzUcPg9iK/wqlD7e7Aekj6uwU
jRM1KKvmmCLqc8dPqRzOuB6bATBf2OXXFdmjLK0HQXFl+DF8EdS8ERtcc/AkbvHKQTMq1xPH6DIQ
7ThDV9VsNzm/fEdWJAEwkF5jW3kqI61w52ic4FkB0nW+CCP7zqwnr24Js5acGYJLmn1qsHi2yQUM
5TrGw2nl59LHv4GNfXKl8IWV1qiKIlvATDdPR6lE7y/hr5sYMWlmidU4uA20IEwZzG3uXFm7XOyJ
rmgBnGm3vwk1wZXB1/U4h8Iq4LucPB8wQPivq7lGsk2c6/CvQWtUEVvct+cWwuMNNDtIj9IdxKgZ
hHvqieIkpNVTRMsct5lU6ln02WYzHVAcoj108H91flAafLGnvGh9M/BqkSFGHEChPVUy74X+SYAF
Cff53AgHqVSrnXwvkajI8sLCddVyCHeO9p6e1fmO6Xwrh0vzoGGKSleK+S1IyfCK4NBMThhTHw76
OSMbttzIVvID0pt2KYEq+JHPK/p9ZN12IjSSpgSKkH9E5cBx7jsRkf3Y394YzoT5V1waBtl/rKSC
MhhzZ1n4YstTWS5gdlLv8hlIMUhjE0C1heENowKnhZXB5lS1m0S5UwfL1qnJQ4o00No/XxgjYkeL
Msi0oOrZvCfFxCk5/1JeytGo3uO7p4pGj6X0DmZ7NRwiVed4MfOI++vTdWD+u5MbYL1KKJyG6FAw
HIYmMzavaRiIsfmiG7dq+D4b6YY9RfpZsAz+3QTkECYCBWsxVInG0ra9q/RXHX1wz+zYnGMc1Qhn
rHEnrrF6RIBB91Mheto/3JK095cYyqWAldqcmnsXnNcO6dTbx4csF52nD637xTU+eKJ7kTpHwUHR
gkSA1op4EpvZBpAYe9iGeGkZ5AHR9QfFrOX7IYWbW1qHWVSuFZ2Li7zMJrk9CzLqb4DxPe3eZIXC
C6k+vCdkw+1L4T4JACnZ/ydySZZDfhkxNkOMLOhTEY+kP0s0D5CTU9RPpDW98m/zz9MEmXaOlg95
amWR0CtRieyFr22PeOeZxNvopBQutqCkX60u7Np3AIO/vnaE1WFWNO0KJTsNYAtDp6PZeDtwQFvr
VE2FXbIODZgvaebJSG30t77MxV+e9OhDPYMgywmC26fviLrmi6p6A7YddiWpqF0aBODltJtUTLQh
FB+DwM5Xgxch3vCM+vPBzmKMXts6K7qtZXF8On5y3nFiYJytOzXaQwj4QEnzlI965aqvFqLjoNVr
H3+NuRf2xdFRMYiBS5Xypjsivgn1soU7TiLHs7Dm+zcyRSiLQk9ISXPALJilSFeo6EHRfTm+RrdW
0mcK62/Nf6cfrOnIAmplMeT+10gLtJw8suF4eHh9qZW5kkNa5dP7uqufIeMUJp3IafTZCdyz4Gkq
Uxzyx+2Jz8Gza7jvy9rFEQW9UaCIeTfxf8ksGTeqZqestXRBFudDwnm4LH/qwFudIsVyGuFZ/tSZ
fq3racpLWl5dh4YFAywhHT5FHGuerhF3b5GRgnrAkXLwWBRY8oA1b9RsD/+Gpx4L48UKLXqBIn5s
Gj2DRsiYfxJq3/uda+bOofO34qu43y3fyDqsi40Alh9QN4A0UAeluZ+7zhiexlwZ4RG2uMooGBkE
IwFZ5H+0OtRFxyCQxifyuTimwdqL1qBt89cbIE8fVeXdkDhXJc95J5U4ZiQPgp3z6sosCwc048xQ
r0Y7/ldJDyCsr2KAA6wJDyAY4NgmGa935Paf4nEfE/oESH6NbWJiLOYsg1SqJUm31X26pUNFNRAr
URLVftSMIHNaeM70Rs8Ex8JheIS33jTLH2q8CH++o3GKuY3vGvnPcZeRg6RWh/T9pkAKVA9+SYRt
i10PHalY1O/kxtyBjecUXG0YTo4zzPnkmSGkv5VXaVZT3upTg3dvT8LOSU1+1PIyvikHSvl68F7y
MJIamEKazkw6+QzUnMbcM3W59aPkxcUFZB0VWQI8g8FPgcEBVTtnnPu1f3jvMxkJwB8BXCXfk2aL
3D22u3jx8s+itCViDcdUfJq9OuSM3HFtO4dJt6NfyqkvBG1k2sg9AsDB+vjUZy2JRPUMitxrQLe4
7c0jPzs1wDqMv0YKVcJUUqR7zOgKC+n9q2ozWJklLlM1MAAaiht+98lVpRdZtTqLZpk25U/GWi5f
JhNWsP8cbVxRUZ0iEJdjVJO4F+KDioTeUVomEtOZSNoSPJUejtcB3vhpJMn++KbwtmAETn3i8YqU
k2ovHt5cavdaYYhByIwRwDMh5JbgKWuPsmx8VLnCqh0Tds8Bmwk3HHIGFug1PtlYuvg7HKxYiWeK
RyI3IVVP+84NHebEMNQ0HPspvYDAmz+WcCwbPSYHxAa2hMpsD36Z9EvWTFZFSCXIsRNHnYgH4Jk4
vnkRYimRrXMf4rXgdZGpOHlbMZD1G6V7Q/d9AaSCClpNjLlHa/avnalsfklRt73kdPjiPol2Fua4
PQjR6+kiwHeCO1Ny1zcmSdA5rgu0rfFHgkY1k35nhG//1Ds76ZczkKMQCcwaqi4DJcRvJ3FHbLYu
tLbjqCfykwE8ShNxsc84iz9sOF5Xo9EwSyncIXZMOIBCnuUv0y+5L78uoCdA0aHU/tz0hzxR6kWl
1h03PqNzsNPsuzAXOD3emsD7mSqoBaeXNn0orcIgoXZR7sEdp94AlyqNLZOz8UkuYWONALhvc9rQ
bkzu10az4BQijZpSX6Tgw+tOfc79XIPgwqknxHNG6eGAj8dVhQxEGkqR25EUAxHYbr9Db7PjCYjY
e7zFqpv3PNe6zCeiDM1xmYDi1UIgguzia3ze+3XvLSg8TXxE/iZnbGQ2kqqHPrHtHvfh2Em5yu4R
iJet5+sWfXYYsb+liJcD1OHZx7VJwsyTogu0TfDvT0lVorloccQNRewQSx7hHu/CHIhGOahSrh7k
mlc2vBlIsW+lMc3AjtEXrXnASrj87ng36B9FRJNyK7X2YK28NxJLTZ4eSFz2soBtGnshlYgSkFAb
uJfq87UdV48vmMOiPAv8SAKCEKD4GtH/ZyquhjbHlmp89zDmxaR/JQPCChis4CSEsFaD1rbpjliP
I8oeiZRboqkThnuKfLPjlbbUGAmKV7JXkurc1C5WcBOdu0NHpvc1TGHPFt1KC46zaNmE+L61yKmx
ueiaC9jLgHcDV7CnH5HMivDBtRudcScSDcdbNL0EdwLALxUv/aIVw+icgENkgc8m1AgtOZn7DuFY
AlHPm7H2DBfs8OALnrLtCZFubgh0l3Wfi/h6f/IRBzWK/LPaj93OP8qQCRP5knsYrP2jYantC3Eb
Y0OI8B7HuqiCKT6Mpn8Xw/8pKiTCgbvpTZawYTPnaFNmf8X/roK74UKNbZwzzxuy+MMmlgnyJ/pw
VmevBRoBlFzoraNhAcXnuItJQwfLz/YE+3N5HAkJg8Op22kpEes6DKeuVPKWo5GtV4A3CV3C3QTn
mDGM6w89XzHMdtC6ZoiQ+UNQt5wgb0WoRjZ/8IWQCitmJOnAH+vYA4d4OpBAEdbvZeHaf1eVZeZx
4/53nR5YkEgNP7wiWmyCugzWbaeoAqru/3d3NAMQC8GlZo/6LzAhuXpuxSx0w9iHk0VVTVxcAh71
+X0JPOTpWB+FvOqnlafethsDInnVoGZXn75HrlslCoWPPVTRQeWvuPW0nRAyhP/4O0QzvE14Rp/p
SjCfMP4oNtiII+mxenX04W6d0ir1zX4zRDNgBH7xnhftnHFp8rAys6Bzob9Ent8I5eGYtagISBVS
Ctxck/OtURw6I7cvQM/vCZIEoa/KiSEWZggjymxefrX4JEOiQDSDz2goxMaARqwozDzFLB8Te1/r
9u151p3EEinWg3dmffz6NhONb8lE0+hVUlhPLK7pCv4KKqzFuNm7etnJiquYjVVOZCFeGzU8XcrD
wJsK4GlpWPcE8YmOXNHPKBzdx+UuBfBggNXi3SsGgCdGXHWfi+UyXoO4X+Za6yUJmBr6Q5fdeF7I
b+0rHu5S8uoUddTkAPtb7fm4u3T1qp9HI+n1kIkAoEulEAhwTbYWliH2sTua183RVusUAFPfjXzg
d8ELDCF0YUobNKX2saPoprRWgOoGcO6/jkGHUG5/RLRlOMS6w/swkq72uT9Agw1n11n+6t0Tp/oq
NiZzdzFXpiw00TaszeU5YPrvxO8H2PzuQK5yW3ggr6I7whShDZZ8N88bCX3FpkT7tisD3xeKip+s
S3oaW8zOpMfqJ2C3AGHogZv92eXuYE7Si+8WXxok9RKdSFTC5McMLfORrhad5YCuEvLIUn67E+9a
08JBMJvfgZ7l61tE5uYYcQLpvaOJ0L9pJeQzEjlN4ronb8/AaxGEoWOHSUpovC9Uu8dCRlzPA4xB
8y0i9XGRXQfkg7660pHrN/9/T1sQ513nLDp3uOmjYZWIIMkwt1lVobrkiCEepBgAARTY3L3e1B+c
OAKdk4jQRkLqYnTqAcLj/paoC7w/D6blNMVcUTZFN7UUcMKbQKjHSpxKbf69fUITzGgeaoP3HGrY
Jj4SdgRn+F2qxUk/6rr76TPZz9v7Gk7h+KgXOwHArDLONh1i1alrdlJANoeexTRwdbMCe01XZqzZ
EjvG4BX5MEojLD4tI1acKsGT6ZfMxdsg7T9Seij/ImrtU5o9a/OOWnX5nMGspUQ7+laLD1pcsKt1
xZ82jG+fMW5N7VF8dbB3LT6WUbbYCaRoIbFBb/BEa7gYqXDa+eGZmwMrPLTV+4t/B41w01BnlwHU
ADa6EZIrFosOwzs/F4+VB/szwXgSLZNP0M2J2S5T0uM4hLpedW5KowSNZ9FJUV9vZJ9iVm/DYkbq
eRkjT/Q4VRqiWGmLW3C2/n9tk8AJwq0SartIk4U7gpjWtzM6V98A9n4rcBGYZQSzPsztMRyvuMVu
qZBBXxLBh5z7AoIn8k67tt8T0H7NpgTmvh/grLSnjwFWHJNAiscqdTEDawrehTdAQFv6FQxHOGbt
lXAkpg1uQMNvidaD+avBhZ58156yBs1SuUQliBGHSoWbW8Br/Uwxh+Rh0zzlJ3QgsMe2ZMJ2RkFq
wGivp9uDoqkdyavSylXy2FD/8m5LaNA+27oVvhmKhbzMy2XPrlxxaObXYING+X+IR16HpnpB/5CY
H2jKwiPmB/R0WhMmehRlEpS3bSJv10lfh8rgn2kAKkTIbhEMKMA7inhy4NGpAsWkdrDh2YsoDf7X
qwivoT8Ql8CeMkYfJa9C78tBUGcnG2rTSlJalhrv+5ljBUqP+b7zOxAj0TLEH/fpTtO2v6I4PE3H
GiPcxWoUjQmmrOI2PA8hTDpuBeldX1Ye+NoE/c7c2giU2/SbtS8TnfOB129tqqh6Pcpx1nT7zTwt
ScIbaUKfAns0gv1K2TCw7pW3OrK2pMEpFnGtXxrivV8byumD7CKXesf7nI3BPWCMsYROf+uNE7JO
yY9N0YcaG0heOzZlWWBx9afxrlN8ppXb0Uq6/2kMb3mULUylFd0sD5WkmvIcZ2fchIwfhxksOIRr
oDHWle9L4WrKM26Fqg56HPxCmXbuwb6ZN1GTt8ntlSV53qqWvoQw8OzdgfuTrUiFiSFFcTdpV0ph
paRmzcxthvI7/vxdw98TQjN7rRLLP2H4s08hXiLjAALBEtvsVnFmSxwL/KfA6LCMWGGmcn0Rlz20
ET9VTRYiHCH4O51GgR5x06bHcIDMtq+/ntKUQxOrnPIfo1PRlIqfCMZTK7wP3rdNO+idYTjYxUTV
3oJ1iK0RpFpWdSxfRCHZIhrh6CjJ5GZtbPNaJNp01FdEOnl9iQGSSmhJFlWvPCcHLB92NXOaaojc
CXjnUQXqU2OKK3I4qC5bAz4lquhGl31bCDuhDE+wb/Jse8Dy7eh/a9KoRmDu47ki/JIXut83CHgf
m8Z5GZ4IhnLSKu4DQrFmb9W58ur8Z65LzBr1AITgPTLLEuzJdarDYcYwmejU7tBvHFDvbfY2Fz6Y
cZdliK450fkXF1UE0MZUllhXR7ndDS5u5Yj8R9E3DsKXye7D8NRtsxavtIQlPwF1XLP2nyOmxdfP
JoMHM02qg39K40P5xvR+CLC4j77tKnlRcebKO2KVJ5733Mxr5GQUTicVrFdDZJyb9gxz49D8a2Hs
DFOQClIuDHs9MZn04bdF7BvENJvvqRotUF0bYeHqHYeuT59NCwopXXEDY8Plju6kgm6YJQHw2UGq
u8Vy1I3/4sZ0c9hGUDkAoQGl5TVwc5Z/camHN11wFMdIDIDZizKyfrGa8nVuk6oWOzl4l6G0d7j1
4UwfyGTllVPCf8RfrK/3aBxTHqHXBAxTJ3oAvdkyKLskT5HaPB2mUGWxpQfocwJM2j6PBYk97RC5
Z5RD8Z15HR2vwCA8I4s9fG8hwWm8Izpo9U+KYS7CRTWqd6N3yj5JmMD6UmbkpWyck9pfQL+jNJkT
9CpNvOf87jDZT1tZgloCsbHerwPL90CsFtfWaK+Ypsz4qORhMYG4Vlq+kiZ/qqrnSrIJqhOvWBVK
kkFpFFDIJCmcMUU5sug61z4q4x5/LDxaUTx9ofyjIxBUQOe0hSu+x3cvpCUYBOlTa4FfP8EaIV0g
TJ6gIXgRGUp0Gz0n1QJsqvWk8I9b31gc40pFj/U5+fYDQ5YFdny7ACVtvmH5yH1RINMEVxp01zFZ
v7WnoWwX/So5k9j7CHmsKqo+Jbtq7A3/bPnEIC0+PMow3sSQidiwn9Z5q4SVFjzgNZTxxI7AIL/B
zmVFZiaVlyuBw5+24zPJw1fgl2r3QeL6mBpUz7F1yi7k45jj3JyGp7FFmBloUzTpdQFI6OSS+i3D
fkKAWgoXnxKIObSOFyMWm/xf5iYcGSWb7QSMB2GSR7u1UV1jQwK/0w4KdzouJhGGNr17xYCxUiuz
uqQBjBJd/wVbjabfs+J0hOjGMBwrX4yr8tQVbih6nW76T51BUjN4Q9ILNIZRFn1VDsmvnYloCUhf
6Or5agt8SDjTJeuPUNjryoDjoslr3Q9DOWFbCpqTn7UoXBKzKUOEZJWpyp3HNeUQifdnzp66xNT8
kTM7pxoy7WiwbzCxDDFoPDOaPrtWLlh6pMwNiGJbh5SNnciITMJaUwbUFs5QouMM94rEXPSPfkb7
LH1qrwwaOapyrIAfGw8WkcJckeK/3/WU97k3LBknuBNeOzjtEstp1bfHg/9vqO40x0vVRJ/lySMF
zKObhK3L31PEd8T8YGJEaTdf2IZd7i5VegiLT2yJLdR4Nhul14OZxJLQGu1RHBeYJRJE10aRrmJC
Q6u8IN4Ih4mbX9Ix9/xAYFWRHLzehvbP+PtEUCDjL3swmq4HmZ0+6Y4GgQyyR0IlqDQ8szdclhbN
SDOOcz/kNOzzOkCfRHZFMmm6w01LIXX2+Zxbv8jM+t1DsxkC2qnmbPnQ2EV3pV27PWKB1Yq0cQv7
gq9TYJR0O4igMdsygD3ogyxBrkX+VD1/oHxK2qKswuWWG72BFkuRIyCMtGU/hwV51NmoiyHDfpWz
ge15L7EIpziYLgUGLY0ZqXSJS1AL6RnZUmEX1DPdr/dV2SKJuVslpENtAM4qIdNZ1b4EXu3LTZRE
gaD3DKGxZLedC7Y4V/o9OXT9IzZv3t6lmOn1PshbGS0YH7NOPMnz2qJIvojAZT3TGEtPMLW4PwJu
wL8XjofCRycRsx6FCpu0qSn1EJQl3MeZayTBKQoYN+n7Oxe4jLCX2Eg/ZNe32v6LE7iBDFsPrbny
E27wotC+ssx9OSm2+O7MFIUrINF48jOsvNZPl7ARxjVxd7DReRl+05P0nPFmkHXpqSuKi01zo0D8
yKRNBZexxZcbt+g9U5MY0iAuSJThhujX+MMMLnu2go3D7McygVv6sL0ErHXK61OHolrx15KM2Pz6
JDq3AlUMWxCnSPI4SXg6MSWImrGgaTGm6qVscqlTzcbJ4EuTv5rqoJE/GSfMkoad9OH8mR/55W0L
xcU8uUjyxcZFJXWiHaYV2QkVhSwtfknTdfqmAM6CsN3YrdnP/vP20tIvtV1lNA3/hjiOGufGgJrm
Ju0m9L6I0epE3Hm88FyUxyPtELtR0iVsM+qUF3K83dpKhH70/qQ/5TmOVlwVRsHXHVsBO8m85FxG
bwgwFsNLau3cYDj7bk1QwYu9g5OrSb1Wd+ZP6EYPAu0cWIe1gaRBNH13P6YQLVGNpar0eT0bgOrc
qhz+uDWVdq70/x1SWndcKDFmIWMqTnlgGI+P8It+EZdFZHrNMtew+YOFDJG5Hi3K+AcXRJEou3WX
nV0MOGxrEpe279Qlxb6ok3lvkXL6EMjp6kseMqxP6fI90AXyQa3BRK7hMJa5UwB866T2H2TBQy2G
gXQyr9ennRYzMe/eF8+vpaAEwFgEHJHxIfzMuhikHfYzAQ6aBV+caUaxc9L1u2OUwLQV1b2h7Y5/
qyOCc5hc1blxJG66J1NfYrLbLI7LBCIll0ho9P+NJCFAh9vauOhXBnVIJuQpLSGghBZWT6VUq1xx
Hbtaw4ewl3a34Vyy/aFKqUbcy3+xw9RsjVz8i7ZhnuF+kjtvygQerHo+neyd9uWCvg3vM4t6hY1k
Hz4zMj5U7PeLoCSnuNnBT4oNnnzoyzOrvikmDsKNrYvyYjtywg20NkDpKTo7YC92cCzCAek214nW
ZgQZiEsc7n7gYCEAKSQQJQx7Wik9vZ/vO+cLJ0pge6SQmfrmvJT6LfPlSzQkWhUNcg8bdn+jbiJl
02UCoiFAxsssDeYTX2MUS/nOIronriAAcm0ceavxgjp64TrB/21v9j3pX7qQ/QJEjzBd1M5DuPGW
xLQ1B4uKos4C7KtcYFpSm7B8+Jtl8BhGfBIWbhmXlfzfvcx3S6GQJqroZs/lBJDBB390iQ/iO3G0
kTDPxhAQ54H4QbjZ4h8cy2fuJiyUzsTQfwn/8fbT9X/OPaIFZSP2s1GbhJKqR1+suXzrjVGH8NDy
rhu4goT0YJ/RmbUliEGqJ7gDG2QUBukAGrHiSqEmsOkG11C2Gk7ffgLeH/IHzfYEK0teehOnVt5F
1L39eDwFSz8RZ4xjmvLgZ0iWyLkuj1z+VuWtHLESrAs0W23iPBTSm0bp3D2NBnvns3IyukvERsLb
Z81Som9iM9Z70kKkErueCwEmnOHZH8sdyOtSe81R7p/OuMnFIv6BToCoFmaL+3t+OLwhcz8Xci9x
6RnXyU7eeusUX4kuUqrA2CDUclrjP4d5I7Bps+xwdNC/aeieiiGHGjWajLJgRBz25EFF6LI9psXI
g4BzYjl9eKN0V4nAUlq60d9KjeZ8ah12IjOa6cEjPmYgpFajV+bCp+7GNfTCG5vpMuRr0f2+8Sh0
nn2/8xweTTMEELE5nAt28PRakbXl7zBX+v7G7j0neEni2a+nmA7CZZxyq+sMLQMug+yadSU2HDjZ
xMYM5pSmFirsom1gvqkzH0cnCZFrEmhwQ5gX1zYcjgFa89glZydnDS3RPc27Xyb9jXPE6JAMePMU
daofsA+kWHToAuUv3mxq+vPYNjg9SwaHrAfuVieIVk66UxsjVIg2CJoG+zI9GqKz4w+mYMr2zqZo
GZxblo/EcyjL2r0pot+9QjjoAhd8AY1C7GnsivgXLqL8TwTOSDa6DlmSNv3UOVeIMduCebjcC4sn
XwAxDzcNV6xkLGY3nAFbBRPuzuzXKcRIIgNVWZbg5OFO+pC1GC0xgt8EzPHAkLZAUFg7cd9Thi92
wGQNvl4HRstP2+Nn75WLqtkNTuQCdFyVLlgKi0yjgglweYOwEtpMpvUwQ98AOGk8sX/Ee17S6F3g
WO7J8VSRlj6tIhAByRjQixvypTdIK76r91lcxmfzzgsYi/oXVyfB2pe5BO/8xGIq3/pGSMPn35zk
T1sR4k5VXxND8zBR4z6H4pVqwEfRWkCucXi0ucTAoLQQI1pJduJ6R+9r1CrgSV9pZg3QtUp0HmW9
uHnjjUhg7IMu4sLdihXopkz7fcEJplSD1o8wpLfa0zKAJ4qdZqbwW6CX2jfgeU9udXRVZ7FwUDnj
yl0qcchpyVDlNkUrBA0Y5ediIyii/6xA938kUf6hdk5MvjKj28LPDy0S0SNpyZ/42A7ZgBDZ1BqX
xE6oGR8WR3TTvAcUFbTxwSyrzQO7k80wNhj5YdHYtZDv8zbf6unXjc9YVyQBL9WQWiBNIOQf88JP
Aj+IFIjDm7GHcKV62HA5DKWzXITyUCJrhw8uPHwnvT6WPojIwuAwZTwOc2M+qtwjw5zzN4J6337v
Lop4EmKEC9Oe7HWOJb9aTNbsefyGK/oG9x85RKncEdE5sTDqWLfQBXq8WBckEZm44cNJPDWI0IFn
KMhAJdINlLcfHPVHA9170Lw1bOMTCtK/tRsBVfiAxE1hwbx0mDPxPspdtVzGYrLRcRkZWUpnbtQ+
OeoweLQu3odf+lTbe/3OeDfj4u4nhbQlqpS5zounqon6Nlv+nd45u1hnrwB0zxy/1ON8KTzGWPUa
KqrMT0cccPZBBxZx3/3NCZriNjvktVbD1Tm55P4bnZOOsrS9pXLfV79UPQ+bUvAN8afvK1w85tO/
4YbBmX3j4Jow9QQtNPdLoiybOKqPR6ayoT5pKgQ84w6nBn59sGrMRt9lFatWEL88IgvgC/DHmShd
QLcuNCy+pGJ7agHBURm8P8vJGjalS/HLU/wBTlyNEBEddhsCn+ikFPG1kuQ16JBqG2IIm2rKXJ/y
yq8I92F7PKiPXJtnpl9m/3VqAubuASSRw9OVLAHPvNOGXJ36X38wfHPjI7SXKl/wLk+bu4ElvCsr
ww4+40kK2a40sxmFypJ4pcWpYgqDGonLVOvC1+NPMDkLQ1tRcY8Bl58FZF6JT2Sa6PB0cmZxzFUV
dAm0/vsjzSFCH8muJH9RpYhvuD4Fb9baZmsL8n8Q790pJv/4LjhYM7gvzRk9tclaoxP0Rp5lmgDw
/6vJhn7tJPOdwRSHteeMJRTP9cz1zxgYgZxZZ1iW+veU4UcUZSmsqu71dWK4tS5+f6cQGZSToQ+k
koi+GE7X3Bg2qYYNbH3oy80ixZC/OvniJxQOczADXp0/ECdBoC82Vrs+I7ptRvykM6hVfYZoe6yh
/Opqjg2oBvnwLBou6j3KtqYIzQe7mT0ld8UOxLwsNzdm4H+uZrsFbEp+aSVhGG08gWRJJTku9MzQ
kfBzQmdpxn87OkvqQgFyoBoa2VfoMygi2j1d1XYkMVLbnmyFTS4bLb9iudZKO4RdPs8HCOEIKoso
msdvI6nhMr5U/hvVb82ZfisKxnuV5hznw19bf32BLiNr1UbiJw206dmhGBEWqBrqWomfp1p7CEEM
AsTXJ08PAdrvvs3E2eMls5BeipFshgMttGh+uvEsqWACaFMmgNiASpQS/AbNxrahKQbUtnlOiwON
axsq//sECeO7fcA5nPploqna8zzqpEMDdQO4JJZoNbe1kiCoUqOwTwwmk5xKr6I9tIuwcxEoSpAN
1h9cwclXBhRu07whLa9RGhy6jC5CabMBIAuA9kB0b8nrIx8eIGYJp331mX7XUT3aPlfYfc6hlq2L
+6jEuE5OZD98rOlMwkv9RHi8Nx/f5SsMZbsCvIZzpaEEoKBq9GQCgd8paenSPbrj8ZwkZ1Yh8/rn
xcyDEpfEywL6O3sT4G2HgysQP1JI6p+8yZI1HM83pqDedJyPYfhTIAsTdThPDb3Fm+t1QglLwYmT
bbYkWwj3U00kxIJueKUJqkCQxRg+KEGACQLSTgmB1oH7fqDtjXqG6sfKWtWkxR6+NPC4aSNTTV8+
xoGv9JZD+uD2vKfBAghV3DEWvsYkFbkjr2WUbTzdIFeQ5S1zOZ6z955vGUUI94aBD3ZbbomxVe7N
wuE9KjczniZw/hl9oEgBtWg7vTb6YcrdmZNVuOIZm+77dVqKXNYXha3iht0d3GLCyySB9UVOU+1V
JkLNL6hDEAdmTA5OCb9vsfnvYLNIbklpKNhBwYrBBw+v5phDkvNwh0UmQ43e+WaJBlul9WYIDf/3
VsrH9fku6N6/IwVOpa6og6t/a083CbHyb1SMDu3vwDJZxVIdZv1IvCyacDCNEhiaZJPR/8t6v+WO
uVlyaHQuoli0rEa/vAtg+JpAWQ7NdabuW7lh1bfO6kCgIoZLo26DDtPBkmMh99P05lElDwlMClVN
kAh0V8S/bj7kgbfg1An4UQk5gyPysjKyvllnEJHvmr606ctQukUeBM1z/NeY38UmaaIrY/WcBu9+
YOpfhVrAdtD9Y8jBQo+9m2fcFHxTi0up2uBZiWE4LA3ppxjrqrqfeBOby4u0pa6Tw3YDDqw9g+sa
SKdLkiDkGnF8+DTT+nInL1ehEpJjvYuLngS9lvVpVO2EWJH5EDOZCLHPeXJmZdqbE9u+u/V/qqNg
J2hMCY9uRsSyLxSBymy4MgrXrQP4Z0KMXOnOCZaa9ZDliZuJqlH4BiClO/EQQWxBO+7n6XeJ5Lje
od96mVNa9fLhZApX8USHUkcA9b5Bm/RZ9Axl88eKE3LWjwPIAYWU9i/S4t9X5VcERkPYlGCulw9m
WHoLO0jDru1zh47Cc8+2/NvJRycW1E0rmgMwDDinG2Fu1Vy1dq/Z13eaDBYnRuS5acqOKThQ09u8
kp9SQO2pOpxtHrE6bUfiOJfEI4dFGkKlAzuJoqzIYh+nu9kSU7KL/vEfy+ntbMfuT/qHHifEYsBP
cL2zPnpWcj9STiS/cA5TNY1TDJxt5o46J99A3wAXxRVYNduO4aX2QRyTf/TyJY5MC/WoQMbQvNj6
rA2KIieQIDjmc+nrHLAJaCit/tXTUjDsEB4ljrIRFcbQcjVMI90sLKd8xPXvTxQCQ/ZrYH4o0jmV
StPWTfmHf0u43rGSAsyfOVPyNikjrS5FNN2KMemkWl2iA2x/eiI3gkicUzBWnB9o8MhC9khAAHQR
kBQ7+3QRtVYqH12JDUZ40LKTfIv2xsnKBm3LbQROgUvgCNk0mU5Rp4EIpXRMxRRnMQacCW2mQOEg
MgoJOS2F+U+y38NgIEMvX8pNbedRF2Ge+yA12tIVWCvmnf/PGkNfdBa5t7/1TwDr0o8QX8sYv/GF
ZBjBGirhrJT0Nbid2rWNxI11ISVpivbafC+IXvg2uF1BpBn3u3r5/RxkIfw5RPkVFLBpfzBlbyGl
fzd24jzozctNoG1ZtU9TPjbqjJxMFYUjRH1XBeXwe3Ud0F77jPlGstu608hiMsR/G1Tcx3DZ4suu
yEwgCNfU+TTYRkcniOiji9kRB1G5Px6KA4RIf0IRyfDsRnBvNUAHdyZTwYXKbqMXgZ12WfhlnMdh
6sL7mxUycu94fF7V9OJOaUUcQ7uvfn/FlblCz2aB6fsGUHSK9s0wAKbXh1QQM6SGinkT0GUxvSn5
WEowWRAwAelQuFSLvYo7Zfy6YAOusWCrP2oCg0gKPYHf+l0FeCOlMlK0+m+I2wSAP6wRo/Riak7S
zWRlZful1KXP34pwTxJyJqvaPJrmUuo69DcLe6TYoJtWMuu1p7tr2ZgYyU05o0ezVIpEHqaUbI1p
FBsSG3YpDZiyVIPliYsDntn5H15pmqXwGP4pM6ML0eoDIP6djNAZcRmj2bwkNAlXOjXFys+ruhks
qc/1MzBagtJSjU4SnPFK679pL6tEWMncW9B40pk5GcbWksKvoOZ4G485HPgWYDyZGh0GjQphAEqs
j5FtpdNOp9/du4O67fH0RNZCSEtgC4gxqa+/SLLQ6yaRSvTY+k9JMKPuFN7aoFxz9C5S7zLq0DfW
O3UmKrvXCXfQC88vqkw/DdAFUHcKWsdhYgvpj1WhN1gQv8ifF0I3hugDkgtkYOHKBiX03O/D6i96
x6RY6WhPfdiwSThrglnBqf3GzbNhvbpH6vUAqUXSdq14GSsV4H7Ex/4lxpf2RDk+aRau2l0a9RJt
rpadcu2q83uobH0PqTrFyqfsffwkaFs+ykPqwVe5YS97Xu4prS3FkNM+5udfHnfIWi2Ba41AyxoD
D932jL+V1CYdT0rDHm/Rcw9oJOxuODD0iZlAlVziS+24mJbBMePWoiafxs7p6vW+Rg2XphFAJAm6
JtX5Na3+GVowTfOS9dNju0vX/W+oQM48d7v3aI6VUkjo2eTcZpKGEAY7/2RTuPaSmUORdn4SJPIQ
ywLJU3csKZgBYZjoR6GlzrhqKrvIjctmNP2HSC83FvplPx7DELRvi+5+apPOsIqxotlzt/wpJIPT
vIlrw0Cj97hqesr7hLMjgCAoglCKwu6moixy0a+PSA3WQ94ceY6OLNsM6pZh7aiut7ZvKg21QI/y
S+/i24O5Gye0aclyinPhZ74ZfyPWZJYl/dwQNudgvlBwGdoRy8Dtzl4vvRFyTnq5KCAwG3NY9tLR
mVeGXXHyAkKz9bvJJD5sheWcDqYqQZXm+z3QyPx+ntFgpK+kqt+kebBZk/wBfGpuIFe6BRE0DaE6
NIYBBY7Wy37chS4GPXdaT4IIPKx1/f11f4ge+E/pjgD1ejYT9V93NSHXQwJmCqNFNNrCjQhayOYT
Ih1Uksvb3dblU+SsDiM5iwJGhRMuZR3K9O9IcxgoMhqfl2csag8QIoL5+PH4FUSK6iZ5PctH6i/1
x6zSb1oX/y3FQwBvDeAzUyhf4vJ7ijlyPHtFrXFdlhm1bCfqvmmuMPns1L0cPf9meXHPoOsawa7b
n1nS0ZcytGIiKcMog9ZA0WMLxTKQRw5/lkuKcyaj0GtxSsOEOHiujrT3I2uaAfoImrCtaaFN2Jtr
E8k1Ih9jgw6KZxLSlRBEe30EJave0CIv/tuQ4AfH1cb5OxcgOg7tiPQz2jDaxpomNFURZUgp0VpV
jWzYNIJwgL9e0daesvRk0lQBEtruB8/iP1LxB4lrU5Y75u1cFM4oDvfDfv9mu5wxhJEFrrC/yq/7
gzQALjBQIjmKL014ouOIgQVjPSN32OSoB5RPW9rJLgSowEMbjJ+sMtMlQ1Leu6WLbJbwWKchvGDq
i1+GQgBHLMndBgEPRku0+QXrYCA3r2CvtytKo8B1krIYQBAi/49sm4ZZ/n/wEa3XvPQ8gdp2U5VZ
FPXxthlf4xr0eIb9nvrmmZWnxhk+jqGM5Ij0pZcnyMGwEpnylKVCU6isizk13XZCd9LBc2lZnrPz
COo+yUMTob35antPeiFiQrRWw4Fq1SnhvS52Z+cKcTt1pvI2E53J2XiBnL8lpkUxls/1nIlXGvMa
qxl9BJcAzoiDpT2PtU2bTIoetJnfH1Cvb5vwZOimzaoILkgDwt/v3ylo+XBREKv/WQVPxo3b1y/x
9J36TzsdhoI1e9z5UROzm/GVDz0qcLfdUktzQC9X9nbW/4dENUrLw0nr9YnHueZevpLMXiIfdNKQ
0mrcvRNRUNxSQmWFKVBm/xRpCUlTM43uo+SqH2FDsZrzSgJ4SDR+mJiikZaDkFlre+qvnVEZyTpO
e6BIsSD6qLbC3kEsFGzNBKNnrwEa3GsXZVBvaiQKDKmRuoQliWbmP4rmEE7OF4NJemFJ2olboYbb
weiEmsYhvJqR2ZlZnTVXf2GMq3JrWHOdEGKbwFuwdF87I76wUMBL2pKJGX0Pz/VL4l0c5gamukd0
R4nUkcaEjZ6DxXj8xiX2kzCJcEheP04ubXpzg/r4sTL2mx66dsfJvZUAJqOU5hGhom18eH61QvQB
x6mwcye87N4Kvxchi2DLXspqWGNTbmtB/Xh4gdNbs2TwWU/V4pnyq2grhh8nHr6mvOCvq5+7JEUj
LZpyIZU9SJhtrU7y3CS0bmDeYtZgjtCB7Zk2tcPakbH86xJ5e5ibXDoRj728PGj9pRQ9rUQNyxmQ
PxpUHtAGK1cX6A4/sf4cN8j4mv7aAab0HNukS+5i0qrfBfeq+UQLBKn2M4Hh8LVb3vjhfblyqfN6
zRxIR4+/cr4ggmOHSObicmgGslx/+L7gB5+qTZN2dR9YfURZs0kw3424BsTRLfJyq1gHnf45LkIa
X7uiQgb0fvg0JfjTbXRPPCCdoXoi4ITJ9L0GYupeYLAp7UcbyF/Qr9ojE5XQd7LRzw9PJqkP3VHY
tflUA/JamZCdXO1RRvNUwlPuJEkvtUnVtPKMbzhdjiyKy2TF9EJ2a5k0fi1q2IBzf3TPsMne2G5x
i718OCI7nS8mOs5pzbU7S/Gq7FQWwJ68Gqa6o5vt7kwWRnqhPHoTdESEIVLa6JI0NWzkOzYF4wKh
7tn0e2nj2+tQiTqMUSdVIoxkPmJwHm5dNHeq7Nv0A04Rr3R9WGlalA3M3inShKZO0ETk+72mSLzb
UU/h1y9G1s6hxVu+QCR+I/i3F8nTYt+4IfbfKBtm7l84c/aBCgt3Rbr+p5GokepNgcMf5HEeHX9W
y5NGqTYUh5BPpKhdIf+uyHIRxL0sEG+i1tIHQ0opip6gGov89ogJkvM7YDMw6zyaN48tcp685CIJ
r4EZAlcFo+i0NR4/XF9BQqYvy1X9KoEILjWwSkuysODywVyvBgG/gPMfOyLqFzQAWMrOppnmyTVv
X4aUbI2lo/Yjqwhu4UYvXDHaBhKJl5RrQamTUNIW0HAjXfsRu0Y0a3i4HPITVgF/QQieBbs4/4RE
MKof2QC2U5PO4Ztu4zr1FJa/v/oz1gEB5ZS5r3FD1PieS7r1YRQHCqZkkFsY+UpAhgbsHElUtXj1
vehnxUiTh3ZIRCc9x1/8LG4f/bZ9XurvkTm9Eb3ytcetlvsRJNFOgD+6NqusQeKitzpsHZVnjJZ/
dJVRIajC0R7Cp2yEqDfBf8X8C/6wJ/zb6SWEqzqhtkcGMU4hPrDchrgcgxUXkp3pUqFINhb22+sL
HjToS/zPX8EA0CJNYPaR595bS1aprsSH2pKg7B5doRiBXwLzumcDRZHJShGU8YrFf+cZDn9uV3BT
8arZLPqEQ/jLzQu0fvyKFc+JNKqu34KK6g7r5ox3ltKRSxtk/Zg+/jr6rfOQ9jaBsqMY3+ds9Jmg
9voZogm7CExxVTOHdt25vxBdFa3HQz72YJLl9WnEAwHnWz1SRuYEGCkO8ELjVcHsvZXDGpv8BWUW
y45ZTLdH4Pii3HTj221loxMUcDzyk66dyaBKy323r4Imj+i49ATsPXB9M+oCfs15YlCHlOYKXB3P
shlN85/3O2zXhQ571oAH1pOeuAB+fN/zaJnlF7dg5Qvb5ohZBgV56D+4Hk7jiuLWrl96FW//XBsn
SoidECZY8ZpayeN/17/KRBiXYO4htUIPCbARg7hx4TAu4V3MkOHWlBMa6lpCOajnFtBIntkQhxqW
OKrupKK5C5AECoxujokxOyVBdDpuiHEmvsLJsUk83lSwzYniSe9RsHNiu0ZUEPD/vag0kVyodum8
KAT5XyM5J3y5bcxxfVHNFp+IbNPvjE+SwsdIUumOCBMnQJdQXfqXids2yDC1/IMOF5VZBhQyxfpR
Q4TUKpjJnP6Eup50Pd4QQ/AP4cekgFc2aywggmgh6+rNcVsGAsBXwZ7jUrHvUP9g2cabytyf3ylV
q1qGTrALWWbyeVSItcWakpkQsVzv1omxCyw1gs5Y4du9mBRGFPo1YGZ3Be7D8AFNJhbmrP8mgGyV
sWvkWze68k/o/bDJHaK/SfCUcF0ALStAGEdVM40UlrEhcTjuZ93kZSOC9ASX6US6Z0uk2QOpLk+S
RqJ1TcvQ61ASiNp/caOnTv/2c0WUlvu8qK/jmD0mjYU3LqMLDweQUzCHCxbO7DrzWsSs90q+qhjR
7+ifxng8WB69Bho+61CcJQUgKQaWnZDi6InlRr57VbCLFYCbMI8//Xhqnaxl06LjPr/hD8PBkrzc
SnYN9UnAkhwPFZNiZ1xdw9ESenZHK40yOnGpGr1lQsjO1YENklpCZWi6tv6Our6i39mUZ4m5PmMu
pDdUZcLLxi0lqfWVXYzbu9VDbgJeUMvke37+LFz13HJHwwUxes0Y3qzla5W7XSZMJe0VktcRNlvQ
2YHIHQOoa97zhv8m0MPU5Rojg3Qslgq9A0tWjmh6sI7+15nCO8rpFeFWr9lxsvXsaTQQM1sV0s0h
LHpYjAyscQo4XAk1fUUtxrULlIN+tsl7jkPJY17k1K6w63x3vdFkoODXaIHnAbG2rVD+tf2hXd3x
Jh/Hzgjz+5JFy5ger9Z5qg6HLZp4IRGvMJ31aILnoorAcglqrZJ6NaaEtiRN6p+5oD44VJCeK7Jl
/Mn563knQfJ/UBeWj0siGTqbvhLURHI7vlyAFU/2X+YhYq3pP3DroLiKdMmKqTZJ58JY1EhVIGH1
0VIxA09j/FKQ7ECMPMHupUzwyWJaqU0FI67H9Vsz5x/IUIjWRuYktiZgFe5wOEaoOqcmNwi9UdQh
4i190TusCfcwKWJ/EVOy3II7iM0nXfUpQ3HGWzzGmpvBmYVvwA5XdqjASA1sKXEPwVDGw1vn7Fl4
48euasmRUARAeJvE8OE3PvrWl1VHc1bBUX4nBYMlZX2cvqUmarB7GeNAwcbOnQWfM/nCgrgYOcd4
wdBYwriF8Mom8MuMZEmJ0aNwAHMuQ2fCyopG/pwji9bB2i0GFnFtPq939+GGkYkfgLDaP5y3HMVZ
yM/pTZ+bA+YE2S2bTPpX6tVxnwPZXA88hHK9PnNxEgLVhdY/+D/b3f/bH3RameLOfPCKAhmEoMs3
aZJC5XBFCcBP3V7jvoW+aAbOT9vll2M4kI/CxfGAkFZqfYFwm+HSOD/Yj728MJnRPY9mv2T721l2
80h36ncoLkskg8MeHvSIlZ09TZizq199ZVr7t8F6gKiQh4YOniTw+m/3hEdnT7D7gLvNkO+o1acJ
cEEx/1uCXhvSfHN4AM86ZggTryY+BYDyoYPnbcdaYLm2HWLmqUc2NjH5Iq5BkyToWaFomBtXINMr
FSv9aJj9lQjfsBBog2fhs1Zo0XideWrYq8JB9Uq9d7E/SoumttUCZkNpbI7CCAsQYNs8Ldas8xp2
sCyDnC1iUfZUH/a64NYeTf4WkJgvVZHZWURKiaS81iF9Sf1HcorxurcSKsXgkcIr7T7KB3A5vr13
KQ9jpFGn9WemZUjN2weJgDl6KB5u5JVebIlFNEbljkZP8IsxsOSfiMFMit7JK2CcvTN1RlhhVpXn
GP2NsuzBqSGq5IHVL42NV4l3PcqNsSRiGWHTCe0buitij16Obxsxcm0SZA4KYoI8sUL75676SCEs
bz4wa5pYf9WJZlGnZ8ylJrTi6eIe28i1H6tm+RCwzwenCkP1e0C4ohVFaPIBnlnr3I+mJF2AUF5S
Od1DSuuYgzew+N+m1finwjRwtgpezBbauGATvXrQFPNwVwXwe1OB0IoVgvXERTy3zELwHTSO/zzE
irreX53Z/oU9dwjLrvb0/zbFhqYO3n/AqXICkulzsa93eg9hDOfWoebDGp6ARa+QyFWsQHdgPevl
TmZ6KF6FeNz7Z1CvCKLWmFvszsGKvDPI6VRvaVb65KXfGQeZOovs6vU6//Mx6/KWPYuQtF1VMqWX
RUkt38mE4Syi4Dfro2KxO4kd1NMqc+aS9YbTFe2Svx7UQ+SCOSHsmVElLa9NgK+xN6mZYOKqLVHy
T3oS9IJDnregfTjaulbld4rgk5Um7Rg/1S2R2L048AZtN2KjiLsexXpAbqjLRKFB3dMrMtGt2kIj
usnFzZXM884gOj9uVBy3nlqJFgij7vmeSeS2JUg1WCVc62Bc86+R3MpWT8KTmn7fWRl0+R0Tzl8g
xN8vka+9LW1yRKfcFTvh9nLF2f2rgdxIiSu7YTnpHQhsOCMma6DoZacxQSnKtpt/3vVNy1eRZ5Jj
eemr+gw4yJlEjzo+bddHd9j8V/w8XRcOJjmyU3bhwDhH++DzUvPjHql2vmbs90BLVhZ8R/GOqp6f
Twi/GTANvFtYcnYB+TupZYzX2mvsO982uuKQ6MLL4yrYMWg9ccoKC8HICSFulCuI4Ak0IJ0eo7Q8
Uu1vaX1N6ZQzzoSil6ez7OyMiwI/36gFC+c2aI4h94BJnTg/iaoD5wooPmg0Vz+QkAv1LK09rw7L
vqjZhIea84TYHLTjZrrfoXNu/ylXlWyWdDmyBsD/PUXJK5mtez0dNLf3c2PxLqk2AK6ls+eEy2SB
9+6x7B5GFUAWRfZYY3UTVZ4RxbXPbzAdMC7w2NtZawoVse+BC4tSiN0smoWAzl6qZvn0uXuCVa/0
TNeUWC+Q5CK2JqWeTbmLrdP0vGyDd1W1PlU2sMID2/QBh+kB80cej6c4MdFVbcvGNOn1xQ5BEPrV
aR1lsRxhtvdq5ogxIFIDA2pA//UErzmu7HtOSNvY37XXL8faW6ME31vGj1UlmwXpJcizwaxpjrUG
qBSIRM47OJuYlxgSiQ8vsP24k4hoG+8X11TjMZG6x6v89hk7jhSH1CsjJmLqp4nEl3unP3rTFcLp
O7ECIwLk6PLR0BHdrevk4wUFNRSJmQQGS9APqq+sobel0VbgPxjtz7km34SuLnMoLK2rq9e5gLEd
gR645kRXqVtXV8Kp+U5flF2r3wQHJ3gXsK/HeTy8/qVj+CGYfg6y9JNfuV7aI+5/zQx1Qdt/80Nv
aJkGhNRWfo3P/7byNc18CbZ99jGjy7qbIrQzrAXunFXIXaOhUUFllyC7ur+WN/1lBwMwny0iKYyI
DpZ6eq2N/cPRSSin5oEy1KeT1//QQy8EI2+EDGAYFxBv6xNv2JaP0SGy3FCCx01iaDm+LRZVpwz1
T4airOfTOXO2a87Q529pF//sF4YBB2DyAN81SSCriFrAxn0kSH/9FaI3lmE5u2RU42NiLxmd9Du2
O5SwZk76AQj0/S6tCEt4SnIVNwVAK/KdgmMQls4gqd6V8fKZ/1h1aKcyeNykkgy7vqm51S9SxaJ/
jqrSSnPqwp0ucsgqs0zR6qjF9lSi+F55XzJqCkPS/ae4sWsDCfekm6qUmUrtckvVOem4SODfeeQK
AZznit2rR446hdlAZTTnefxrghIVdPo+JVqJntx4/efnpSg9uQFAgaUFze0iJwTaBg5diw/EQhJl
++JJBwiw+iSqIFZj03XfcStvwOP57tRwlwh8ijb+CEptaha2JO7B6Mfz+MEBFu7bwvD+YSPJRT52
XoPBLJES4jyRjzVlWCORN7bFpoRcpS9ZFoFg23IYItDlhThgeQbkdwd0VxXhPDYRXbGJDk4PSpRM
Bcx9q8y1fqC6LfL23l17O9XK0OoMgqf9X6/jxn1SkQ5CcQrcjtZgML0JmkU5TQX/42Pz4nQX20JR
zsyPuMjMsDVlGBrIWgdc+dWAYTMYtqZoEv9GT03LU6pLXu9LvC5Zu3L7OsQUkpfuE9P7TOsPfP16
dt0h8aEWHNBcvWa2T+QrACApmGpbi+xaJ1GwbnSlzcewrNye+a86LqftjOqsjNXvodmJhI2FfyOJ
dDa5L9de09oAwBmHf7kdsqChChdYj/0OIl5OZGqMFje5G2WmsWg3R9tR05wNBXl9BVoWK+6rByk0
ZDcKjsukYtO6pcUXwU7sEQPJ3xn9rtFyS200Az6mqrnSzEAv3ugGTO8uQzLvI0F60b9Fozi7eorl
2+L2sNC/COubjJiFqRN8ArC+27XId4A1+xY3Q+AQ+s5/1UXR+08G+U/uAMtsSAfHEJPGMQfngUDS
9YDKWHGtCaBr8hLtaDI1m9e85N0GSldsvdZJWSIa0TYgiYyKyWE29yO8sO9nmTq2K1Ic/uUqnffp
FWvZMogdrjqh/q6qBJ4o2N7Hzk9slPTiBkp0OTJuxw4ng3BUUUyZf2zjIo9PHh84emZBFO8UlGSy
UnMddEBZt2wU8nx8rcdSvuZqHrr1kwQB6G5S2Z0n5RClTnc+yNL9j1jtif8lY/E4UtOfQZBrp5E7
4XStrAOlIEMdD+7suXNPPxsTOL+XOitAwIfe+lJQs7W1AShG67OUzHJ4m/5JcG56qIeDeCA75NAz
wRBaqtHBHj0iJBdkGPmoG2lnOGoIqp9xiKDrC2VLq2bvedHDDNZjmIo6WpVmvxdllnIcejUSpJCC
K2e34DkheEjmhiUDIpoAHv3XLn6N3GGU0a+Y7p0G57QqWEc+YdG3pkNOVOjNitxxuj+eEQb4zFVd
ES+R43D1ctX1p7pjhXd7LzaoIoe6oyBZomCiB3ZQ10pmv2e7TAy8NICm8AYbB+Q5WNArqAQ1Tniv
d3GwBr37YVjX0aSZbi34t7yShNEgwLEH0O+a+JFNoiyBsW3J/I87cx3EYNb020SpZ1Ksv0fMoCV0
QVml5Ja7VkObEh2SVxDp/1uTdNOK7Dot5YNS/97c8lv/jt+eY2uzOqiVPoxJjMJFDS7tssnaOFXs
Wv7/DcEz9hFL8GzxJU1BdZ1xq/b/+PQjsRyorNK7oVDPD1yyMyve/Y5fKj2cGO+pLbyRCgxTrq4h
PhvTlT62nPQtQBdA1yj+p2HarTKPr6zkk6y4tK2x+wLoOsZwG6ylV0gh4sBc7W7PcqVPiOW2Jcyu
6qF6ACyneHjsOwkTPRXcoNwfB3DWzLJZ7YWApiuiOt+7RCK4PBw9VZqQILPNwM4KSJDiJAfF87hT
0kyvCcLZPZ4K/bJNhzXwOb9GOd+p2ivA/f48jtR3tctbbvL4Pws7/LikVYjTCTus/zRcBOBthxPF
x3/LVIay5KhyuzupoZF9nGbY7agss+XuFyb97NzJVnJ8rQn4YjAbNnl5Kucv4cSb7SDOG4fY5mW/
9xBEeg3qapNF7rUZ1k4X3yCai8tZhE3yGDKwjXkAP17cGxvwJj70tL+buMLrFiS1R57WMB7NEERb
lF50loWYoslAlN6whIKq06ve1NIkDdodbMCm6PsBZHt82pnc7g1YnQNS8eaVHEr67UOZV8SVBgBP
1grHZfDPyctMYdhSi+OpwWiMn0s80egvFXbFDCoNVhwN8e+PZdnnDIXELroGhoUgCOZXQGs3yQ3E
ZiE2clzN5Mr3gh6YhxwWdMCNAV3vBi1NAW881VwpZSnNuiR5QhKJC23MTZS8VWPwZtxaVRogN+uQ
ddrLJ1r/936BwICAxrshB+Uu1ec0dffa3u4s/BP+ciupqVJ972gwdEePsFP3Dyx5YRg+8QG0bpYj
VVkDH4Xd5JJmC7j0lvEmIPIxASXiCvay8i1u25xF/0scPv9BRJANY2IDJWMKb7lG3R3FHvV8TpAg
JTVKTh9y9ZxM9iFeEpC0Lk/RYgUd57lF7MQykkkSaxvKaNj3D1Qcax1W3bjGENuIu1KAbSLP1SrN
arSA2UhM0me6qs8wUSk36JkP/FuS2+CMhBMG0ypWjVOb+NG4v+ZoOmJWGZ9gBI47eeUiv4uO8dcp
M0no77SRioZDbHFV1Tn5/hcG0R2l4ybJ6SMsFdmDIbsnW5ltxqTr/dzj5+LqNlx7erZLs/3xoha4
UrS1EK54d3KqOQeHe60m2ANfunaLpCutSHpWecTSzB8RpBOx6aTnWJADFSlBBZN2xIDanPoxBQUr
JteOGS/O1cTgk4nAI60i+++wh+aKtWUbqoIwvucz74uEouOYOHklM8Q9hL4Jr7f2v6n3YRW+6vOW
GG2tgX09iB430h5vS+f/nBvC2CNqefAsgPIO5mJ/H7GDEO4AVMTdPMh6a/edKgcpMpCP8PNnu3l5
tT3BRlDH8+mOq41sBty0oovwzoYg3MetMKpi8P7zSEDsYL7ZXjBnEk9H2I7lce7P+Z7ajJeKxodX
Pz5udzWcgOV8ULArMO7WWlZAigLk+98rCDodFK5oCj2P7WqLkOvr42OnVH6/maegYlkKWhqpImgu
7kzyTGCuFuTXFtiEzN7jyjwmWBDizut5VdySslUXzkD/r0NjWpA8KbD+Y9iMbJVU88nCBFrkMNF9
t3xyaJB6AmG8HFgl3p6KzGmvgsTnsrHum5f8bMQ1ztI6iRsBNQuO5ir5QaiMNOvB8sLNpnW19tpN
YJ5LKo5+MW1RUP3MvOm2lROYcvVUPtF3jDCVOxxDsxyaBezbsYdrpTrCjmaj/fbM07nnPeNuxZW6
6Vvb2z35z7ZeZY7zVVy6gbpQsjkw/HuwIpsArXRhu1rUGiMyvf06mzFTNq/LaQQysarD88dph4QA
/lralpaHIP9kv30UZIZ2/tKIfwN0ySobYUNTzzhOzUVBCrxN0O10bGD12CPIEbw7CFWa+EgsgSTy
Hv34SvWdD+DZ1cNSUh1JtN9CNyjTYK+tgzeVMv/0UIQOw81qCbcTZEtkrKPaWJGdRbr3ZegshXWS
ReKS+KM072eX/o64FBpL/V0Ljgo0IglSn0eZm9KzUhiPBP2GOFEfo7uT2MqdrCbfDYD6N/0t2UvW
3IsYJPnbnBgNCN4wyBLSFXiabOLsemNc5Fy07AGS3LhzahVWSpCxMHKIu/imOe1xiWRhwV1BPRKF
Rjml7+VLSRTaEilWLvR52Z5nqif5bAt0Ix7hlwUzxoCWLpKvIwnDejmir5J4dc0ypsrBHmDVi9Bv
i9c8afnCUNmXNgr4EZj5+puYNSld2jirIFlYtY56rH9xytJkhwxjZYDvExnI82LLA1BN5B2/BtCq
qS2t7axX9XshMmYDXxBR8s2+lhbb/0gu0IDLYOnN9TsL7iAqNljwDW8/hA65RYkt97F8OKp+3BMP
R//ivDmqc3MrVrVcuy7OaxTVn08lvRX1c80hdcFgWaeP4aOdCY2Y5+d0Zq1TWE/hvajO6ku3RQyg
6GwVfst4e2uVoqMzFDMxnQyMj1/xhj50xedQ10I+49HzXnr/mfECegPQJ77gUVCPOSw7lsvemkT8
e/qoQOIiFMKN4j3ai73b7UDm3E4swoDUu0BiHOIBvZT/cWCpdwgeSGYzd8/kFvUHg0D/+biqHp0u
bi2giK/E7+cdW//1aOHsus8Prex/uIBsPg27fpJBqlM9qnzNOxFWN/w/oUMgHgWy/STriFJsNuG2
ZlLoHfJtfVKU1am0GOpOqZe9Dz5btJx+aguHHbjqc5ShhdI00f8jGeSAScp+v5c72Z2htz8t9cl0
5MKgyjLnwbRSMcP7xlrKwv07yRxjBlhu1wvO8JeXOyOjmNTYmvFFIK0FPWpUTVf1gbVLs4/Ag2Hm
Tcgsp02FA5SKeC2UN0PiGjqb2mn5q9DGWq5MzG7qHhif612WnRYv0S5UsMvwt/lX39RM4VLmNqCo
TrBpajVh3wRB34S0p7Cghpqyj4/CNVzNv4Q3gvo9rb0elTjnQqV0tUdBx+Yg574i5DVavRpEYVSc
DTIvyp8ev9nglo6n0NW5dNtDg+MEKV8Wy61RCOLqtKKyUBScaUiAsp9QX1Ug/eGy8jhZu3YVqmvV
wNGqbPXQXm7KpzxNyTuax/nTf1K/ZOQdpk/CXi+rTd/un7hXr3op0U5hb0d1NYtIBqrAVEz6xtHY
s5aSevHmVx4LbIPn3lS+gh55T25qslEmgXhN0LOKNCiAGcWHFfXBcQTgA+8lEW2zVqRvXKL0Hiey
OZAi8xdpsrQrsHwcuTqhPhakx9ehZeXcHMCd+MjVzkuX+Uakp6KOERa9bt7UDj2MYXpbsYyYJGRK
DcoF6xEAISUFFL4G+PjOh4Q3aEudWWmTnE1q/8FvudAiuUWbRksylN6//zzC0brdloUD1zHF9waE
eszCDdh2lkOfwcE1lKuMCMPzXNip7WnOY0sQqAHjIyDYLVJT9/QHpZiIrpS4dIyOXVZ72GGf4ZwO
yxcfcKHelrYD+cPPpF9Oqx7ARvKj24vV4Z4kvY8TqK5M1IEhRrvifFBoRY3cHcs42+vPkcZ/ljhm
RLGRrp6TniAn7bkk2K7mZrm7C0AXGxSV1P09n9C8yYnqMn+SzU97Q6X9ty488npSXizhB0DZAT2a
G9fzsulDxp6cbP4teTF8b3UVygajRAiKyp1+270LsuUVs++eP9iqfZiMsC4+wtnytFc3BGCGsS0z
LCj/toWGMEmtUfP+SwHnQ5Rig+5WPFyfj+cc5HyIv33v49t2Mj6KhAqBSA6RzFBUYV93azolv++r
DxxhNA5KNzE1ZuWiXuqZQ/owbrmNfISwj9P1yiqnj7K/TlV1bNFF92ASkhNKoP69qgSsB6mUbPWj
CjfhXJ2FEEMk9jQ+tZUw0uNl5StIeYMi9YGOlMOHJ/QwxQKzOSIzz83qL3YwrNKUEXGkXFzR9aul
r/VrbzsNS3wTi8oR0+c+D52eTuqMniPy0U2uELbgeAhL6SzLPrAx1/BtaTxOYnsT+1lbt/sP319w
RVubDcvAiciB4UxPnMB0UL9fLR2qjEC+9oaJ+d0abXTI/fOn/e26HqfKvnWbH/9G3LG+TQu1T9/h
/wEGBdMAv/t6h/6zjBJ1oTsq9hHLKZQd++9syw3ueOVW9mOYDpLKH/JDA4J/AfZpRwfZnUtN7SUY
WgmvRs/+KlwmgMJU6rklkL4eov+G16slqu1x7w+ZVZF1tw2PkttoQn8K/ldYMhqE328gI5UmHed3
cYHHpHjHhNr+jniAW2XgHjvRRhmz78VRfLr7haje2QA4H+AD6xsBXDIph4RLjQoBrfqtLBf9HllB
vcz57EKTT5mR4HptiEBKCUq1GFdRgyFc8C5f1u3/jjpsuZbAZE6wOlPoPy23cBc25/q6wIobjDrM
Z/4e72+xNjJ9Y2NruP7rUe0adlsBCLPaLpxmk5mDzR0jsMbpy66DIlxGK9poxKJwtKIAkWlC/bbD
jW+N45en8oO0fy/YzFKKeOAt9O7QkqbOqBYDv5C9hPT38/qrPL0EsviqZMnUp5WAAhGQH9kexXTN
LQH5qC8XMeSVy4GjamcWp8vIKSjQQbLVuIWrUtwMmfRdhbcWVhe64Sr1GPzhsToih46CnqXfnsJK
G2OjfFBmvTMGbv2EvKlDE0x2inZiCm6jMRPIyKQodZvJw/HxgdY75QtcIQgJGxOhon19d4L3Lf4d
UrvCg4/EiQRnGay4ti+OWlwn7qZ1GvwzLTCzThx8MoQs1Q7H57rcLW+6/FeVquBRBrVyfgUg0UeX
0g90J8z/vYJhgDD6v0F4rnz+wUIsRyDOYqiXbK3n7VtfK0kxcYIBh1mHdPiLkJvHjrT/G/k/94wu
ZXR2tlk2uX/5hq1mVUegwXKmqlwcGY5ABBhVd2e+ydT/kkoLPIgTpEoiUrAKPMkJYQ2MUSwGAk9L
0nFb40TZlHIkDS3Q0Am2N/67p1VxPpYFYdJeNcdlFE014W5XD+eSrnJPyA8HpFdqrR1TWmHp1fdP
3faCRYCUgAmNyff5UCW3j4jS35fG5hNUVlg9MGgw69o/Tswq+JXGApsXsen8JYm809keQuGW/gX9
StUTB8OvS+lFhERUm8fV+e2p9SeBM3r9Cg+eawuY+axW7x5d7/zBoUOjnxjxdAXMuKUP5sZ+vNXu
8IWlBv5Se9lK3UgXDN9R7yZS1oSHhCiDpNikD2uGBCBqA/JCUjl3vXPOgkHl6U35mG8rvT35BNOs
ouNM31ydbnfIBI6JbrGtFegdScZdtr7e1pmt1G6Em21bXWCohKNhIJ9JnQ90yQMITapQV1Zg/Dug
ynL8Ja50dP7vtHNNj+eIJvhezCyqMaW0JP4yAu1JT6Hvcypmwqn460L1XgkNtpx89Fhr62qmsIqh
kMTFgILXiknR8cEz+3W0bRGU8s/gSX1mrAHrR64BZFWOBQLsFAcHsq2zDcYcYw2K8fUG78Wyg6iS
cAvvl4XOWuxOalyEjJiioD6ZbKSk0zieiD900RtKvwTZT3ksFPvqn47nftrT16nsLI5zTtxRNyFe
iDFqyIrmDGJzjN4svmw7QrLYfy1aOKSCt/p3Y4o6OF2UgYlOb2sCADKb3YjadGKPy8R5QVX6JaR/
kCgJfye2oNXKIr+v6RW5EQMg/q3UBdI/aJTOyhR23BSf+eqOhLBQAAYIpy648kYujBk5kCTOHbP1
wpMtndPZv8Xza327l+gJvd2NBghl/iBGG4tRkwhxo7o7E8iEN2d59oZw4HyDjCCPfb2VdjgYemhD
G+Ev8DK+EFeZv5F51xaGtWxtTKbhAg23CRqkQqxvysk0ZuZ96ZTM71Q4Wzh+gUfWyiA9QldIcQtg
Lhen6E71jwcXZ8ns1xlLyGBCtYynSwwtJdo9Oq0UvNSkyuAhuS4RLJmqKzhpeoRpmsQeo0qeb9cH
bdJbZCtQZaYQPUpbGHf3cegFvIVyHHioR4/tonSaaB+A3vAk2HLEScc2ieWCX65Zh20gJl+5DmFY
YhTKLY7txHYfXHbP9NugeFtyowvcAQWxuVNck7u9p1xmuP7j8KOBeEeAuKCTS8QM4QKQOkgRXO3p
dqnVZxVVg4AbW6knqH33TanxvJlc6Me4vfu6dmAZUhm7ZPI6jnbONdoJs2SkrgtKLjvbc84ipDbU
sFHtACeKeuOF0JNbZQkg4TCA2lUMMb56c8r2/Q+NOwUY6Y3rm+TO/EHstJO/P9t8rxUU7+R8XG58
hHEjJPM7YHLE4kt4cLEBGw4ChHYlsYU+lzO4G5cAsKz3c374KjJKvcTqxog9So5vx1ICr0O6BGz1
TMfTv0VNUpjSWxPj9fWAqvL4W6OHHzyUZZN3VTHhMG3VTan/OFSwxWo8c6wg5Tz3XKUBisIVYp/5
bY8QMxF1NbT80JRD7svd/w6J2LVwPVl8bR5xvc5NsBokz2TCb8LUfxOS3WtwSuY25jDjjJme9bLE
5zxulyKtg1J+oy6smn2W+PpOIjLKUk+Om4utJRbpoeNQPMMCZYHTZ+aJs3BRjYFPnWlgb8YZkrBy
X7xhPzMnQaojITzcxFoHIYij6LCfGA+mf0m8rDnFOQBR2oes1FpherEKKWknKsPm134tuXEm1Y/z
qBiyz9SbAswFtjiqWlU+XPf9MvyN55y2M9jmWNbFIRpjMOHLqj5U0zAtPA8JbAb5GGFga1QOdY3/
ucUbPWF7uj5bHVmqnMlnQ/pt25fnL8f8pRMt+o50R3rzKkSVJ4C4FtxiBNHPUV5/7+USQ+EYgc4N
089IIHgmWXIqtE9tzur+/x1g9vZHAXKtrV2NdBJVd+x1/dLJSOrmCiKR49z80wpm72O01fk3qAv9
5uKta9PwiTvlSZOyoyMdcRv/tn0HoVYMa9FArrdLFvcrhzHYYwWWi7F4IwXQcSvLuXgLGXkrLTxL
12vVExV1kZDR/7Q3dP0DHWB20pRYQMCNuH8YhxpXIjHofVO4Pbn9d1RC8wrcHsTY8/5pmUfH31Y/
yNPpZSVbwLnZVdE3JicqqTMHPNe6qlxdUyJut1pvdRqDMWLEWasPgP8Lczgrw8hTh+TJ9LZJzdrp
aCBunKnHzM0PXklTEMXCW6t7OD8WmIPexvZbrVsqi68WM5t/OyWk3gJvDvF4tyvxl64RYsxfFGpo
Fs2UeyG0zlkcDzxgWVS4JAQY18S9TTXVJLYQbeVJQ+ABwgKTZJNdCWWU/0aL7/8K36fdA1m2SpDv
ZJ5d/TRZNCw+S2zG3QPDXJBlFh/67PcVftnUB4rdHurB4HaSNwhwF+9N1y1BJ6MrgeMY2Iw1Uvu8
1kT+rPUSiO91cewNX8dWdcJKx4fLw06fgdHY+0SfFH2AIaCz9pLoG1YYpfw/+kE92O7gUBkJSF+V
4/WsZ0jS+TU4blSNs7miO4PRwkroZqreDJhd3xYAfMjxp2H3fSV6TKeo2U6t8Hfry9IK+n+CkVYb
5t5e1HRFZoMYC2jrxP+wclPO5peV4O0zubshN6P/TyPxrtj4J547RTIETSW0pBJrcIWEUSKiPYUH
GOpHvXtS+9YzWARyTNyE232EULDnBbydTFmu+sM4sU+/cf/PS7O5opdECa1LL0gIpypvOqW501tO
HOpM5ul+1xc4WM20iyhhomsUUXFUC8Az+rqZFktwnprox0AmvzDeSPHY99+xDZo9k4z8N+78ooYX
ICDmsW8g2p1DQqM/x2YTphe6zYZ2I2CNlqiG/VqZ0hhv0a0UmVstnTwE3lh7rP76505Dk5k7p7CA
ZzgSRo44/fdtja/LkmuW4hP04DR2mp3O9KcDtsLBEkzr2dH0VLfKTKYev5e8WyWqgy9V8klrURDj
42U3GR94OHArOGHGYz4PuDRvMTb5t/i/xetvoWe9pyp8ieHiPUbXES4UHVVnjqopCJ5t6+inHdpo
1SsWPTfG7qc6JZNIBdbB8e9G+5P7hs62jBd8FfP9FojmXqbfRbntnXnOmKxZgb806Fnh2z/WBogT
ZWa4U1qRe1HB0mzoZifZFHMN+g1Q4oH3yTn2xAO3ESBHr9ECTHcMsFI9ypOqnbJRPKE0/LYDBqVh
xVS3Fldw24VkHoj4dbUfHPfSL565zPUK7ogX9SzvBgH4gNkQmyPqRx2+haT2mgj+2qZmTTxsXfX3
iDfzqdsbt5f2YZmcOom3M1hpiV/U5JrcDrn/FcE1IwN4ghQxU7l6fLfy+fB6MZ6Rzm70NVyLIAm8
p5HnjkDsWGwl3vSVzkQsTs9dR+xXmVeOqRwIhLrw/brUnCuP235lZoHk+LVRpR4Z7S49gbMJIqIX
a7sCd/Vy1j2+qEbPqNRg4FjcG9c/J0j/Qvgw2OjilOQCkTsMSq6njoUcxAElCDxwLFvv9O5p0S4l
u5AsxML6F6p2rPBeJG307BOifj3W0Y0AHkx5f80lVmNKFkwe2LZMSOQezM5oc+c2qRCxba6iE8jk
eoaTkb1hKFKz25nqSCU//AKuMKdrAzYsiZbPOmUt0Bs276pAstiFVhLKBnnP/OKnRC/2S8BZqQL3
fUXnmBi/rtkOcXNwZHRM6h3CWXwkS7o3ueVT0HQJdyi5Dq2m8P3D9/vK1q0t5bu7N1v1CYNYMwRl
3Z2R+BpJ9zuk1w/scySFkP4A2yAFol35GCKUB0XSuLtwLsCC4/ZLYMxJfwGpmBNy9rH36DMpUUr0
9+I4JhjYERX6yVwHXOzQqzD6arp/gwWmvLTx+2yjXGmCoCcd83/JbDaNCyI+6WKdbha17MocALC/
QCJxPh66AQL3Rsy2KAGS+/jobcrC3qHKjnqwyt6Y5/7bDc402+FkKNWJh3K/OpPJ7Qi75cPTVgLL
BieZQ64dQGq29xGN7ef+793RGHPSUQnip3md8vmG0Fbn0Fq0DeOv9GoJySLzh8MRsaJEytZcbpLl
HH6XtaiSfoqj0V40ylw2zPYjOR6o69at69OrilP1cEaO9pTfLcu3jgEEYXJyLKydiFfC5J3bXjU7
AqkNtSt/pOgaCM3vba9jRYf37x1ylNG1SDXJzgEP+o+lJ49ezdLpz8g3sPMNp0XIfAJwb2G58Ex6
02VpK6AJaG63XaQFHfr4DDNoAB/wzZ0cl99N2EEykYuEkZSKfY2gXX3nCj1Fqi5Aa2jo9tBorsbn
8wLUxWFyiOIjNydDicGzxrVq+fbI1tiY1KbpwbUIwjiZniq0spWHe/pST2/xx892IqWBEBDOqK+P
LBJYQ33CC++qABJ/yPt9Y8wc3FFWg1Lr+UiIpPW5b3fZ9ui/Qmiuqjoxug4TVO3hwHLPc1Bh/NpT
KASmAfa5unkHaCrEnttap/YK2QYuxpb0TUApkzR9IENDeiBEzxyLDfxFaiy2CjDGv+6oyutSTWHJ
068rTZp+JPOANb6eJd5qszmDVwEKBO1Dh8/YYI3xqYkWLIviJwpVENrn7w4UtIqDHjnmGPvHoPlZ
i+UBIFD84mFP5wKXyFMMvmV31TR8S0l/G4GrPNTc6W1XgXTLxR9ghqAuiPyltbcUaLmIb+vrERds
wZFDGAa/s1IefKrHeGigROijOyHhnslqZoW9pnzWq4iBesNEoUYGn/wwhErB1sarIZRqek+yfHnD
URmAYsNXzj+p1X5Eq2bsQLHZoE+WrbkZ4/zsib7enW0wgaweNbMPuCXexSElWgrdU0nHEuUatMIS
IHhfrcbytBtxh6ndZYUKcoe1Li9ADe74AunV7vyDyUMvpDIBR/RgLTr0jzP/9Rk5WN3tXFfzyd+k
g8L7WJQ13PtcjDFyz9G2aQnRruC79cAaB3jUrSLnvEEIoj6BTeecl1MbBANpw1oS+WAEiKEX8LxC
Li4EqkbNDO5T38XCRzVCS7VBjGghk1UWLKPzsL7i9bfdbCK7bMZyEmsj4qsA8zl73LTb7r9+wpun
fO0T6iZsI8Ftjp9L2lAmIFGbpkrRsZpAu8z6IMkDGpNDZP0iF2SpP6gH4S1RJjxw23CDv3Pa8Phi
QFG1YtKcQv030Qxgm5F44/yctLWCBsmv/ReegtXvQ4vLiDWI6xO1+i2fKoib0eAwFNkpXJmJG8En
lC8PUuPNkRhrtp0UiFlFSPI64mL1QB83RFbjhhwmtt9D2E0+lHa953O23nS063Qqh5c6q1bTHTp3
/g1gYp3+pilUULDADsfLPeOcEF9LT+Pgp+4cZGADxFMoYzyD/1X3yXTKsc7+gXqdW/ywL+rr7Gj5
ailRkkeb7qb0hcQ+eqFU8hIuVsKEnuQ7CD6TnaJJoWJTuS5dKmJ2lV177Lp9Z7CnUBahgy0FrDZW
qUhjbR4rCp9P1dp0sj7qSG9r9VYcwo19mS7/wDLq6CuqMYpSvs7/PbfISuAImBhPhlah4LtuLhS+
48NLi8n27hANGLDQMDB9DSuOYimS6QPQQmIgRskuw7ZCMI/tlQQ2+Y1g3FZrVNdDanL33PvC9ate
i+V4+Zh4rvHBPirZzlA+00fY90HsyxoKNz50F6LTxyGlLflXODKBByRSZuYRcwbCEpvUuF21PYrN
sZeMkvjZdPt43FWmdZLa/7GVvv7Wah7QeCk9BgXZw3X0yRTBdW5CRWDO68ZHqFEz8JVRWNdYo7r7
xRvT0ivkURS8OwkZvK5D09HIapWV92KtWrp8PhSbFRCqFwpwbZ9ZmzTHGktAhj0s6yip7iloeIee
YnIxcR/Iix2idR+yrHJb9PANjEnJoEVuFgMdg56aYCcL0c4MaX8TvcaFZd3C6c1a29UaEXa0kVYD
iQPIy6x1InQTHTOhf5Ff7Iaitz/gMz4mVXqWq1jTsgjwR1rueH5mEgeg9RkkwKwAFcPwSH2CGzA7
oBmPqOfGkipDCiQnOcy4WZeFi74xrck9sO+hONHqZ27A/hk7bB6LoBZvV9Q0D91kuioyoq4FhrsZ
RXTaTm75CZzw4MtQRogjhmtGLiB5ySw7J+nda4BfpbZy+xxjsbB7GjP4zP9yd4azDgP05WCyE7VA
UaqPWFSrXJc5JlVkIPqiNhBJCufT8eTm8Ft5KSzMD8W+/Gi4sOQKIQ4LZyKvJnf9eS+4mJqRqVyp
xDM4Qx9EF3VU/cjDTsQhdTm5us5ABk6FwmpzMEhu54uxpQIRPWURtF3TOhsIjL+nMSvASMkUn3ba
pIRYIwDEpaei21IhFx/mcJkJXhql20XvaVIIV+kEdeKHWAGSqCnl/h2u5VzcU0CzNKyWJAIO5I12
OYVXUV/j+M6XHMsOXX4BrL+2hYMO+PoJKZDY3KvRzCCyhzKUppDJd71v7EoXcxG5KK7Ky4dfvsd1
GsuBEWAKUHz4S8tfmLIumgPMV5dfOfE4t+DGgfCrq/wLY0qHgIeQppX4oObGKpJbeKnH10IJWvfU
KyCr6nee3HadNdR31ZRZoFlYD9jRk9dd4FTRlqh+cLWC3dXqmQt2y2leFumyL8GL7TedmH99vRmR
ALhQ7X+t3nHgwkT3s8GagU3tf1yCxOWuwpXRykEz+1r3GaLixaXxJCmJMwXm87iJzRKezT7QUUzF
69SNy/XFwdZV+CiHGG5SpYwpVaxS5q0Uyh6pMS2gjD/eT/yx5gpoiLZ1kT34AJxCLn87geykLhvJ
yBFUQ2ZtlEw6R9B+PK2lEghvbzVLh+nE6wZmCkGmW1t2MTTo3UOIcborH6O+qhvbeYGBTFP4lABM
Sc+FhmYqG/H9K9421GEPSWGG+11zCgYAufpO5YZuhf62O56Fu23hn724KMG8CAp5qnMU0X3fFWl0
H3iY0g3RGhN8c+tUGTnqsEsJbKwCbT/HZIoqVIqdGF3DwKPF6hqXFho0uOAD4ULFqPajlCOsK4si
Bk0eI5Aenn8+AEI0o+dZY471GusQWMapBnA7Hcb9WGKxvFkfG9HAjWcSaRo3KBxwleDzgE72LXVq
VNUutoYej93/nhL+6ScoOcSK/+olvvEYQYtki5BgUoc2+PuuF41DDOOaO7UGgZn+1DMm/so2SxJV
ztbh5b0gyXbrYdoHeGkLDD6iKS2kPpiQIoQ9OXJK8yOw2NVN5UTQGtBIBnXexVRipmG9S/Y7jIyL
YyCR41w8MafaQ83uf3pm+y4pjEKlqfLv6zF1ZGvplbRNCL/uYRYg+7/APXyEd6wFEtD9lgy0Hsg8
9ojQUIabQPEKevgXu7k5AfknEedbhtUyk622d2/DobGl4K6kK1/9nCApiVZunDL4YxIM5vwBgdOB
54Bs6NZcHGINeU9TacUunyHNdQWS9ucNWFp6xNQy4y9Z1voClW2Atp9BsNnCl+FzCYleLnwhZShq
WWAqfQpx237VM7uaoQv5iSLGgvk5dABHKlhTXWbSBncNmU9VX3saDAsKqiuQOgCys5vrnHMDUEL9
xCmjznNlxSrSBa6f4pRVUIMYbYiGqog1HlNBEsDHyVV9aZQSPj+qhR9cOKhAbemgKwSi/nNgiTkj
GWBAFn1k3Euq2TvOqyCWRgBvaynVnm3UeMbFSzUjWDzSD0XdkXN14TxgGphF5mE8r2VJ22Lrjmn8
pXgLryitlzOASl6xl7OTideD4QH0gWkQAKcmLkJvF+vkjWx1U6j9kwPP7Pkk7fJ+YmuonhEy/IU+
Qj1WsRkKPKbJL/bl9QO010jlWEi7e9yjMXWTBLUNo+LL2jnJhqz7WB5JilbejBpuKUOU6WSEZhlK
fFVdN7YICx3XvfVgMPHz6tLOTu5wANq+YZYZevABS97bpwWzBKyod0Jx4bjkbmbAl87ONYg4W4iS
CH40vCkXV26ZFvKmbBDTo2uBLNjYlfqeqQf/jgJ+EvjT3Bd9j5SAN0HR/g9UgvQ+ZlpGFmWQqJfK
U0BMnCKup6G5SVnoCAeUV5hKP115ySHROsJopmBac0i7I1iGk9Etis3iwjDmMz6oDI4up0TDairP
HLb0jS42XY9F9F2UejgAXeah5XbiERzdYkPzxwcAoHYVIJywHke1boZEj8/sBV7Cpzy3tCTDH+Vi
zE2bPKz+1i0hl6KHo8Xjtb9PS473Nnf7aoA+C+2Zd7B4q98Hp/VgBg0Ip9a9jmS5x0kCfCqEAEJj
1MYwN+10HJmiKfQwUhu0QGSmkSMRNvt/k8bCmlUGojoTuNEN3mmWhg72hXf0zupYZYVNLh+vv8JV
swbGoYKWLRDykflHe6Udum1pKvzLyn9vqTYFY7CjLe/DXs9I/RMVLWAcYwInyWNdACOMXBulrqIB
keFRQrZFQdGVIxTjnk8jFjXSwYdOevmrgYW6nhfCHwXz/ujnSs8ApZQzPU58PhN3kHavqkyTiBPV
XR+jXRNqxElfkIRk2ngJN5S3KH7bIYtDQ27tN5k3bgEL1W+mMkrzTAPBhRBp6JNZIClc1Wk1Dg8X
t28rLoDOU/KesFPkZ/jFvzawBsj3FMKt7jdJ5eo4fZCbIFq0Ciec3DfnwxptAb3oxzHxHLms8FVU
t/RfvbaoPLwkt/Ao+y8OpqDW7uvyljksyUPI+NQr5ah6S4OGfLerJURizVtHlRpHh6oazJIsWECM
CSvi7dEpQyIXdSmJlXXEc7l2C4aRzpPEkAJZs9E5oH0gSPPYsJFmCek7i+PPbAJqt/XiJrnQ8ieE
UxnfvDs+5sFH6ZebNwCDAFruz2S5InTNsjVw/CalflUnMQIFJLPxoHKWP/j6TGNaoT+rP+oWVt6Q
ewcj1r7UypfFemesvu1+mnbbkPgSmXI27ERa/z3HHRSE+4B+5adCfhlOKZBplzkVwKzl0xTi3qaQ
LUy2GoEPhnDneGKNykLZYXkxjPcuKnM0/oSNFzTWCF666x56Bis2v9zjy13Kp3H9S2Ac4ijDKoqA
AV7HFwW7qOvb6+ixApf7qArruyUSHmX5wgma3wbuGLjPjI1PQayw91xn8CtECH0qtJjQ2V/SVZft
PtfI0NPuUg4Tqmv+D6ZWNmHkmr2ZcxPq+4nAa16CNDQSSYh2hJKi89599ri32VmmG+4olguKX/+Z
uLJFNtSS65zh8iKMouK4nd29TrVYvj4/RxUZ2PMLobCvvC8tMsC5FzLHUM546WyMpwwC9b8/V8B5
RumapKnaA1NkHSF7r0AemUrgUFo7P9+RxtKiuSeMCSImMqNckqNl5bljF3wq7aRUSstemxXSvSQD
wQBTg2P1IMLONDMOpn46f+5SO2HM/Bhq/4KCJC2e8b8K55DM2pGYw5m8mAgdNuW0mcpYY7V9S/UZ
qJhsOyPrHdsOKPmpUa5aoB4373DgWvYTvaS6WOBDgoohWTXIc9Owmiv/XMTSsV2STkCeXDNGnuCr
XNE8D93Ff/QK/DwPovd2tbP3CC+Ij9dL5D3ZwT4sUjSBtyfmshX4i2nxDnnS2ufmucQ7DbvaewKg
u3xmt10FxxbOKXrDzDW4FtCBf7YP+Q3FopiY5sQQZBTtQpXsUzVV/XDFIf9a9zKAVQg3Vuzt+2Rs
vXSewUTmVATmqPAgnIrcWgU6yaMLaZ0WfZaiNhsr/wDVf6HMOFRhb9O+kbZb6Mn+uS0XE8o8TYyf
+uosjoPSC7e2F5gdeZxZad7yNkGewNQWM2H8lj/YnsyAEshn1CskixLYpgvOK3n9YvuCJdznBf0f
vURKHVL9Rlvpwdf7FU/fVf9R59+rzI9tPHXEuLEqDHIv7I5/8NRtZjSveU1eZ97sQCaxywCxCUiY
zD62LH8Uc8vho+I9lMtJbvPrmNMVLRchqj3Y73Dl7BdYznREzZmidW4mzM9kA7wSMZL4ArqCc2yd
Ie10mAEbQDDi1CyXtsF0wZ4R8Ei8PxDcWealMFLleH+Hc2yt3tmdrLjaASEEkjC6HBPo9egFjgF0
uFU0fb2CtqiY3FQ59uHBapvUZ/5maPlL8L6nbvHfJtCYbUPumqTFvWuVU+6e5HmsaROYQNIshC3R
HuVRyFFQRnOXg+41scMQNtFDz4hRs8SktYMHl3eemHbeElf4UXj95NO9v7Vf1GUsMB7SZQ2Z0YO6
zoyIcRIjP6XSKSxCvZKu7d4rogH4CHrJh2GNf10bWvfjQaZg2+xJP5kokScZK0oMf4osENh+qgt5
F1vZFenh20g0DBDHl3Cm9Mr+iQi0EEW0pL9YZ9xsyR510Sspa4PRrid4jez+UiCOoUykvJuZYnKu
8rNtdLfIX1NhJrGT0FtGlP+72U4KUGGI4LB8oZ4VKZmklnwaTRyFxfaxwj0wALDSsDbYlmErqDJj
EmZZUKTz8ked9FWvCX24ZH4i+s7CtPD6E74L1qPyIIWK95z6UG56Tx1dc0ruaoDmbz7UHp62uw1B
ptUIgcGv+D8aiifIOY0JgMH3PBB52S0vKi3HmlF/LlW6ldZCPRu10/COVZa7x8lWvaxaP9Wlzjyx
NNmY2xYaYTt4+S4Yg+Xz4dlmd3NjscEjpHjougQ18OSOWpPlwIwgbDLRqnv7KKG9GIRCMfs13nNj
q9enTLuRpVENuFLkt4rNm0e8NewnHPQjbaUiVr4BX43kF5XmrE9SBgfZ9w8EHhlsoPaqHApKLni8
89a33lWIbqQVxS0oHLeCBUQwc6rJZg0f3rTZ0Ka1n6qfK987Jv5GMgQwM6vs7aM+XuxnozDiavmg
OH5mSGw34qK0qiUeEqAMUJIPpPyYiXG/afUSXpH3j3+nmLG59UasmEonCBJ7Phh4gHs17SimaG6W
4spDNc8qAK52kbb6mF917hCIo3L30wtO7HfI7LAeQh60Jc1AsDMfaBZ67Eq2Ers7nlvqjfjdSd/8
gd+cvTgaxhvgGdW3XL+zvNUYO5AzS8H+DrmFRFqs+3KfhxgYSEVrS6InUpl2vZhmED7VQB6BE9ql
Udmlf+H1mh3z7J7il1tqatPR15CmsxHpJrgRqnk9N6iLldkzSWYXkspDLk1k8tc3fudKe1n+40Bf
pNLJdLl4M7/9EAgkJ45qeM+Nbiyhyjd9C99M/55jZ6M3hSvesbbfzBn4K/HRS/UwjtLAYuZc7OZE
eL31NZkrvfsQch/YRXcGN2Jg4gQuVLfKMpk9DgouHy2zeDwC47C5ExjlHDP6XdM0fs6ijCXV2YUI
wnfxzg3jQOhNP8kVfteFBG2il6wgcf3bxbW7/o299oQQxE35wloYg3yRCRafBAw4qwSAZW5YSacS
YpfXXzR4IgOYjdOsPp79ftWTW82HvYbMOupYNhFeasxJjTQCQrFJUZX7LXu0V4vSD4xV3xO8nXAx
6yTBNJcHIuNLZvAnMzweGZrnLu78ELVlNU7TrD72Ga0vCoCI2euhhG4eL8B4fzhB4Kq7EiZBb2/s
DIozmADi1X/IYsFk8Ps2QUfPuvfSRwol1oyFxwwKBVXpvK2xiNcdTlKe9e8TbJUOFJbnsu7ovf+T
iUNpbUWfsecuupmaya7g7K1pZUQcSz2k7aNsP0iMB2JPV7vU2v6WPTw2Oo8Xf1fvZI7VxOGyxzFP
jaHx9NbgojHlxC1ezWPQ2m765JV4hdlsYzfN5UNxBeulK7aABgGq9OsG6cbG2dMc3M1mfB8JtaB/
/cr/9Cxy1XVWQG4yiLEpBpy7k/WoTXj4ChicG2Gsi/Di+6wDGMnbCDPNAG7y07K1RqDa8GJAzfvI
HKaBFBtWaODXhD6vsg3WwfnXCEhijMtxrUpxz3pMvtoxPwHWFMvIALp+ZSvmcEvrk0eZN88XWhch
wMEUjpkW9xJOA5xSE//scWnBDZAZ0rFYfqUcX0pIUZXQ/LEqF7WqwCowdZpKFel0MsGRmF+3HbCP
+Ln52nJbZtxrKe8q3la8Xi0/nGj/GifEiCHpm77XhN94L6kXjAzGpeJbi4jE5WSR1PaWT4zoUqoW
PGIRO8j2Jol0s6HhhvAVjfB02f/eNA5NzoORs9VZGf9nvKsZvzDo+yZ0REnR36B+KAs8z6k+zre9
gzi+EWJKpPUAQ4tF7sDohdweJSjgNFM5RmJXpSJ+xhHVsRQE5eUB7zRB9eDZeMj14e97ubcHfsn0
rnGQnNT4t4FmUxlwN7MmbiSVAYkY5qQTBLlTFQseql15BN7poETmEM/yzq2wM0K6x0jlRDTQnxGG
jsf0MOtENgCexxDkP41WSR+OJoWxjAfHeVlKxKcDSzXscfpkblelEYTleS2MgroUy3/d1ajEWBbR
jnK2+XLInYyx1OwXIiUEttgYHVoPniktSmx4jjmw37LjdW50lMEDLTFmtaf02BhD8teBH0Tdppbd
dOtRLXCZWARLx+KIAaT3mIN0/Rm6ZaIJqSf3XY0tf/7OCrgRA8wSd2elhJ7p23kijmd0ycZZu3bh
66b478WqgVb4FU8k+LS4rcFo7z4Q4htNjX/PDNlIwsDlf3+NI+UFk0rqtJUTfwN38QM5YEI4ras8
g/iFYreD96oxS08BFmLhtQVxnSMV5lxfsVlya2CYwT7W0SZRrIf2ypEf/RGZYmAdy+pgkuL+avLm
wTXPgJnZvCgiqtjPthG+Dk4VZSNH2a+HGdg53TklVEZ8XCJeFZ1OcP75yKwyh+e5oaNkDUPL+isY
IE0+trjauMHYjlwAtkvV8uPxvfnnOz1xeWL/fL2a1fgB8lZoaA4gWd7ZqCRmqwqG6tWvtXC/rI2s
9eNeHfcB7OVRBeX3HzHXUFZ0jBBbhN+QQeShdlgFMhzcC2rAzPNNTI/RClfGMDgtyQaPpNyK/YUR
ipm+bl/WgkVdaadN6C7j5aKvXSf3Ewcx8Qm4+wwo9gxVGp1HWEZjx4+bgQlalTJx2zW+dNgA6FXC
YKIWmOCPWW4R7JcXfJn/wI+/AymkqxRw98tLoZqGOO24ykf5f7x+VS85NfDLF81Dvuocw5d5j1cb
iI6g9S6wt5Ce0sPJuB+rh++bx81OlbL4QrvNi9rmq5VVRMOXjxGtUmSJFgfNNzb9GCbe6BaWiO2h
l4u7mfRATU7INsBO76oX7QNzBBFjp1nOHUhgQ6wbXJoXywZs6rjV+B2AiJr7nv+WIW5nsyFuqBCK
OrazmQ9qln5H68HAXzUURt+W46Rc99gk+NNIlCa8guRxn9FCZzUd3ZR5w16xPwn6vRLUIDlCWwRP
Q83lqAGoENaINsWwODQdy/vXngGU65NVifxHXRWfCsdrftHX81zoCNrg5JapLvimbfL6RC8f6dzC
+I6EZJtcnexcsdvxq0V/jjBkxyCjrxKFLaQCJeXbG/INwheuMIAi4vOSzR9mZMzgauBSCBMrAYcG
IDKqw7y9szmjXTnWDkv7oxkzdhdFyz8NKx3LYtgEQMsg5R52q3H+fqb4jZAwKtBkzkrLeDtzreg3
xd4oG+C3QDZHqDFvqRqzJ5Gxen22WgKOmfCzFMyaoWVqkTtBTq37AOWfoOP1HmqruNg3nQgih4BY
viL9r+kEFcXcdF8iSN7syR1NKeso6o6cIuhgikifwliZwQijtGVPtStwVvDp5ZiKB92zPDiAtRsN
r9WJE5d5kW2QDiVawfxGrR4mnC94MR6J9nLa8pV0BkBi4QcR3QftXXRYR0kowhX6DM5TN0fZ0ntz
SHjPQEsVZk9sucpg1x1hHtsfzSeVA31I6hCGdU44WSndeMuRPzSlG7QX1BfWTTdgXZ2SwCE6pxfB
ykOmiw3gWsFh+C8lBKoGKUKOsTDvuPTXRBzS9eUWRqymnCzKYhTjFOPcASBv+aEfNR50G7PHx29p
Cir8rCdU4YSgykqnYJNeNtS0DjCFl5JXiw+879bEthHanehqtsl78De7j+H1TGCYo3/tzDm9eZO3
I6M39T2mfpwEZrYop4J5wVPzqqfa6yW+ACdaIllQkxDx/NP+sGH92kvnwzIXlZ+gP7HCaWtqB9a2
inBUhJf2QOD/n0SFbi/5HFwMJcDCI6tUdktwh/QsnFk32G/gFo5YCarCwKKlaurKecyDVV1nowrd
8FmAAjO8n1N2Gu/fs/fWxG4yEfE7gT1iyNCij5guHndvuqx/NAZE/l0nMchQg+9A2zDO1ol2jIym
bAro3m9u+TePm7csBl1htIXNAp/mNyUfmTYarpJeu2QclOuDeNaHGNWau3qD1z2uAAmGoXvv0YQJ
lKCgVhslEA9jtSITftjrWfQpKaS/ZXF/QCL3IwR1xeoOtdPQabNGjg3suRNT8lmsfQO5zps/SIYY
Yczqemde6+SrczNVGW6RmexJOA5eXoh81/GCgH5vfcEVjfhDtPCYa/clTcMjG3Nj2EilaRul6uIY
dylfP5IXJCfGHy4DbPncjVqImBmBqVnDWNccDVjtBO+nl4Km9BpZWEokLDR8bEu6EI7O2G2G6cmM
lj8O7GWnnoYl/DdwoMhAdN3cL5EwRaky4twN4cTOZVElSbLQiAhLQG/LZPvkRBbLVuAgApmKZGtA
6PJVYlrb7soOcvGdk3+wX4ei11ZdX1kzq4qZihGCQOxQHOMjwHcK4xaTfCthQ9dAw9v01xxrR3mU
TOlkV9FrAGiL3BOA+eCss0NsL80IIRc3Xvi1gwqjD6KFVM6C8ps+K022pg2fVwIpvb93UlO7kl21
BsdQStfWHRkYO9tbZCzVFJXtYVnrYd6jeXg21P5UAyMsysN3ACBeyBBuNuww8m4DiOcZh9BoTx7V
Uy7gicNs3cIdqpHZwajZoPbJT6bJsqsaCefquBrJbxis98NTuK3GOfGTsIH+gPxvWTZ39+Xv8aXb
pYPS9hW9rQYNZCfNNO3juCrzQ1JbH34TVi2MocmhEwDzQBRaObq0eJmsY+uZpHSPmFeKv9aXfXrc
CDKTm1k5cDWYPtx5kBvCQm0TqByI1bLUYeF1LcW7n6tq53iJ6s6RNLw/mbTPXsQcmKmh2OXTUp/M
t8LrS276t6jjohfsH1cjAI61PaS1TyyKHWxt9oCxObnxcrlVhM4pxIOYfNVtryAPJ2NRk5yBtje0
GMJ7pBVV3t7wGXXl1qqaFQIA3OoqEq6cVHil5flhO/SRri8nW7iwtakYySrwdgZuKaVio0r9suAC
e9TSqy8gP2JClq7nHjp2L4pPmpJnMsrLakg9cMqDxyrT8ipNEfi+dv8VMi17V1uwUR0yD8DHZloi
1Z+etqXl1jLERUUbfC99U+koyVIyof4Tnd5Wy0ylB+bBdgE18aJisIfI0nBojty+yJTz8XADhBlx
FJ27vVj3fy304nLl/GRwmQ9dPo9vNsINkfxKu1G5o8hJBJO4qSyEXSkTZX7pfC7AXq/e8uxjmjpH
wkkZIfifr2B6M5KHxWfMfSN+NrDL0FzqMKMRgZGzNUsy8y2xGTxdo9BkXrKjOMkPbyF0jip9JdZV
JsdiYes/86I8y8HXewo0upgkSZ2FI8ZUHoinspDq9n3rDgn74GWrJIkzvj6H+IZn1ggDW7KmlcF+
V7rRNFIWLBqQuigdfjucpH9kRO5WEmfuAKFTFy99ZizMMLBb1/5YDMqgXxdS5uOMA9qhe/IyC1TU
JISajGqubC/l4jTY86qsJpNZxLK/v76p8OX/FS/Hf3QUycdixM9m66U0jd5scNm3K1u+OcBcJo9/
q1mw3C1i839w613vaU4vZscxH1sVzMMO0V4uzQPd+EcBQ4yoVd8vGvtmd4fUjSFOA4fdmeI+C94Z
mxKtEql2VWxbvnPRVItOi1MsTNzw+8oW0iV1nypFs+aHuZ0iAawwOsNOB7j7qrxANSP7DQRXkTrE
+ApXgobNxr9OrxLlqpFUA8r/MVpko5wRqTAd1WivacdUzYZAW8bFndwslu1QtTDQ38dotsr7f/p2
PwMScz4QCprj8KOt8jpZLbwpPEU90vjYIE4yCHevAC/IxpRvEeZTb3YvAVpFHwJynhI2QuSg/PBW
9j7vODxEcyxZDBKGi2S/bdAZShfEfD1MugRlMB3ke87vZyejmT7vA1xFk17ZDEqi9NNjsXqJpziC
lOloGhZAWrQoXlKWP4WJRIRiHNanFAobUl8jZYAZBs+XsP6VH7Lf9hD20augFz53fb0r3q/ln8nh
dG+Tqjtbm0c7sjjkdrcu10/OwKZzXWrPNKwPfnfXKG7EYvWBCYzn/SeeIZvSW8Uozk9P8KSYM8gQ
imNYDLU6w8zldGxzCEqX7y5wGWH2ImFDdLSholnAotnTssdS+SXcSnBQ642jlNHXyB16zovFgs/1
beCsru2axlFjoqCKKOeKRtmLUsK6CazKOObQqfYki0poDZ8zoinzHL/j508HfrfRPqTeqs1pfXmj
14ukkIC5HiWRZF9wdXFvST79PJiZaBkDFJo2vvpFn3Jgi6sT+oTqgXufKELtEj6fQTGkSDoTtaXS
D7MLhbMnMjl4kOI0U4GczGNNylZ2FiO/McbEJhKQIMkpZECm//U/axBUbv9+tIHGeddMUMK5Cgxt
+75frl3AaNP8Yla5EAH/8h2qZjo6TKeDpDoQUVeOi+o+VLD0eTv7bp2r4gVeJGSsLq56Nwmk5gwv
SLufibEDap22dil0ajQzF2GKu5Gguvz7MjJ06gQyBdpkB9qj3CPFzJVRNcxcMuX1yqdCd9xNy5Bg
zMDVNE1ZBOQuSbaVwwFLUCbOg8O6EDRqlQtp8Rz1pOq3NfJX03kDjvhJHypJ2c7LBuD6XK7I8OQZ
1xU/LdwVrU1aeZOj+KenVnjTs9wwca1aBRLVi2ZHfV1mrbNx/HEhYQb34tdtz06L2S7nP5lsjhJc
65IHuQu+t9DsA3SSP/2pxyMXDAR7i8mWR1zwf8a4w45mzGeZBjxCM/uZhk+s3Mz6Y6rKGWXCAXcm
T+JK7qjxhaQFq6XtPJIqYtfExwQfGdMOLDJGtH9y7PK0SKyVjV4ff14NUjec4UG908xxzRreGqWc
DqV5QyuoCVxPbFk7sXXR2rL4a9qo2WLJ5menSnw/tphSHkskZe8o8r0lv3qTu53RxNS4sa6c+5O8
lRhZc5IFZDCCyJIMH4KErOc898qIet0dia8cfWVjbcc16E1HVLihjos10tdV5L+EQ9qWQq32Lw+j
bsFYJm67kdSPQ9wTbNfrC4J9p1MAIbhPne9NXm7oPn3P3TDKiDM7pX1wmoMTUzGC5ijevTArzjv+
oRYNYILGooT+al84C1F3Hf7BhLAg4Sri/1p4DRad9ZjLzaLqA+bfjZZGd+ue4RdI4IleYLj9AzGw
ihM6KKJ/FqtLn9JIewEO9eG4XHYr8KQFeSMkyNM37U7hOOlXdixxsOaf520F8L04wLsW/IR7MIPm
pimQs0T2OKA/C2U7hb6GJTNjJQz7tjWelMlV7Wcc14dEOeVbrADqKA/vYm7n2XlfZc0w6Ft4ficy
k0Wi1YM/cOBnciTd98yNrZ67cjbpkW6SNUS6a0U1MHU0ESKgCoFZrqgoau7GAY/Twc18TXuLxnP6
9M6dDCIsblMK5AZzjR5hc58xlrB9021B5PUYmqfH5pOhXb9jbP+HfKc4TWQl5HTVK+1zL9YcoHqV
NRgtf7hlR11ZwaQiaMhX+n/USduyKHprwgaLgTPYYVFzu0R94qyVrVBFQBVBc2929PY1vhDk2Rzi
JYFUQAsr7I85l/byJsC+NghXjqPHWxbwnfEl+rNswh4taEO86U4QKxai2dI+uTIQMYckBmTdxbHU
YCPJdpwSqRBSIZKAbRR8v5QIrGS8i7UdaTyEWXtcvbAHeud+ButBsHNfRdoSxHXaEt0g75z4f7VG
WiruRrA6T/aGBlba+3Zk91GdvTFaPwuQTlZc9RsC6jLC7qSoa+J1Wca4S2yhZglfJ+L8r8ri0xp1
WOtQIaAcZOOuuq+t6pgH2aTE9TEjKB4+veiwQa+Ky4QN0qc39h3yZ9k5NImP4nhoHHjkzuUZV+n7
lUiOkvtn9p3BIgxrV74ddafehBCCMntahPWvefwAPLQw5N+PlPhwDt/sjGBRVtvHj6/JFVnkUnya
ztWVtPdfew/M4M/z+m/IpHVOFyGOeXxZ+YzvuuxhiyYWyk6w4lQayhsbk2qkg8RYWT8GUYvOJ6Fw
Muxeoek6uCSp2J1yVJYpXCRj4BEYg9AT0S3p+zUMhZvq5lPasIkq4Bo3i+byy/00KRnv0dZwKEME
PV13Sq+/UoJwZc5dGRXqrRX7SPOGXXoUfHxaEqKtVyvZqRR4srjpYGVrkO9yzFOzG34eOXSzFyul
DauC136J2lVl6s7tnEyXVgPuz1b0u2Qj1fqMHcTTx5xJskNX6yfEYCq+eNmslqYukM3hgEtwTC4i
s+csGA7z+jiwJTOyCo8EEUtxQap2yrhuskfkdGGGMA+mqy+4xqm9hebIZ7w81EeqcRa5/wAuKwVb
PtGfhvFHXAxC1gx7V8/FlrzThryw4Pk6CyD5UmC9xXzd4UEDt5Gg8a12GDGZlu6bU9z9fED3yTHA
nTDeZhqT+EviKZOpxJReAq5AZjHZwjY0DJeMgJkST012GcQVU2e9dL/sk5DRRxCnbmKbIRS59isF
VTiDOxuRN6OoE2Z0Kpc8xGAT4WX/1/vreqoYD/Fu0nqCtJozENcgxjhemiUiGGGLvxauFvo258qI
KnOyMH3Q83kOxi62dWzpFj+OZeOO72vWy/gufxeWDGOjtA0E2eVgA5tPwwJPXcs3Q7ovSeepT3C9
OXqvvcpYH/dTHeVBIsGe4XpXvmMVijA4rDfbKIElQYrCapEbhVnXE88rYmHmOgH+Jlm+EneB6fdx
CEU4aZoDAzHHxQS4pl1fb4s3dgrryKDShMjs9gbE6Oq4f9AVBUj9Ab9fXzSOUAKck1ifw7yxb2eU
Du9VGcq11LcRBvyT3GKcdOwiNHnNAN9tulfGXhHom76Dm3Xl15WpqQjwKP3hxme00xINHY4S1ygx
WIgMZqT7JRc9u9KWdFe6v44JClYDbiM4grKIjClDHgyQIiyJdNxgyy6fdzR6esH+JHrKLFAUOFjE
7QPlVeF0MDEkZY6km3hwwGV7meWBh+F2xmqzGb1FJI3646Czan2pzYDTGLFnf2d8aFSBK+CCYuF/
Xo28fSwBz3i+8HYYC9XViNyEZxGa0HLvpfmxm2b2P1cd3o3iqChF5kxUEtd/oclgbZeha/dyjCpv
GcoD1js1H/l1boXGYHC74BHzHPwbl4rwOGNXTr6nzkJ0VAVJAyeD5tdVb8CoMzvKwm5Ueep/rGF8
a+O+BgSjNbFFMZXxGDA6carX45S+ehscHFpUdhhIFpl876E17ERV3A4EfJQzc8hK4tMAQahFc2HI
Ngi/c6LYQBTpzTD/8wQCvOEdBaVcXXBpO3HFGsV89uVyNl2MnCoev+bl2UlU/TxraHlyOXAAGPlF
ajPxIZ4whSJeKR2xJj7eXQmmJXueBwOnqcm2xBXGInLQ0J8HoUuUwA08Wq7z0LDOe8+eAXAvtavb
D0Fr5aix8nStcj6kHGimjRB+pMo79EDK4mMyj3z8LopkR6aJgI2ISGok1KfXM4Ux3tqXw9BDoQ03
6+pyJBCO8SHRtnUr16URcarTNodu6x/A3FcMhfo0azesnXKqg9LVNKLmX6G8LxBRqgEcy/o+jxfS
amGsOs6PBYalOVSVK5n8bmyTqWUCfvXE3I3Oc5MofGc1i3DykHDn4Vk8w4luZ4Iq8Xl73eTVrOJ6
7m7sqYO1i/hOBFID07U6iYRiQ0jN9Y+393EUhjmlA0h1mJjUh6/w8Jk9RDrh60tvD1jh00aqCBhk
EVeEJVAC3CboGeysIccjlLfLKpucfabc3b7vL5HFXzAGSuAJPgC2lJyrFBlYxKSe+xVVVeg8VkWD
Kah0MIfZwBxlw8mO2bNgh/TEp4/CMmVYhRNTmSrZdkPXy8KXbslxdCfxV5whT6RZIeQgpg+G5vLp
hWi11Y/ukzeYbxt55sH4slyPYp91yQUHKk8F+kmwepcUF868nyjG1Jsi6Ep9hRp528GmuDEV00Zo
FrfpSdZG0+n5H2s3Eqnx40J0mSxNSd3QiDfxHWZt7opkuCarLGpMg9eG4uITFMcy9SqbQCt5kH6d
SzclIKkrp3ptPPeCK4WsNy8Y3ixbyrX/6+jOv8kallDr3+Z9hlsI5vWROHBuZXS6OErbYt6LWISy
xYvwXnfd8TqUsBonXMXQm2LWoGaz12JSJ+RvkZxW5JVM+jkuuJA2zc7XWSU+nlk5jwrc2mVWR9hU
fkPgN8vYXXA3NxMyMDTUACTWm6+C+qiUfDsvFst5Igdsb1NkIPIsCQ/9XClTeJa/awoC0OQbjN6k
Kvfw43vVzgcX5HVgJ5e1Xs3UaQmZzvtbFQbLHXUEIFGfWa3yClCdZ8O3c6oeDqrtnnaQBpJk6CUy
zqS4VeLgAvCdGlnMw857Qr+A88tNZ3T5KPJdvkKiaSW+AbJvcwmEnhIxR5s16TBeX7WnTgzWw+Fb
TEo/OI+mlog74OGFYUxAL3W9+AVfCRvnfc+xMl9gS7lecbszdt0zGR1u5CzoQijSrdTTW2F/KKnt
xLysqEy+XOjLXJe/bncT7JMGB+MKnxSWCjSxfkCI3USe9fWQ+GAhmPYHQyvViqCMG7ZthtMeXyW1
HI3iXGra8WjVnUcl/AHORZoqUuOH4vtScLDBOvkZPwcWxfD/NSo0CvWrtsx9c9+/+WvHalbFa69/
Mz1w1g+f/uyUMkEDnk+8c1SJaAC4GFcif0+G4Hnqo9nQ1jjZJjJIiovwpk1t5wYEwNuKeyJVGd/T
8JpvsAOgIOJ5ehqsFVc8oBpZmEQ7u/wpFfO1Zl7iYyMue209amcL3mxCeBYIr7sEtvuEDoQeHkaV
OIYjqK4+w3ypR41v8sj68NNblRSJuq7DrmEYCefF1cIkP97wnMx37j/TSA+LNX2s1f5xW8aW+ZzW
NGSm36pA1NZrI1mtfjDUekhfXw3pfCQlGmzqNW/W5ttkkpqfut38TPyn29z1suhyuvazItUTG7C5
dtchuKfAhnIcvr/X5HTbMsQeo0jVxbUAfXIF2Wu1YXlJa8saCubfnj3/i3tnfjGW4+fZD42/23Ur
iKqYMcG5PMgf9mqfNOqE/xjK6/N057o3KSHUdKt+iW6lqoVdx7C5tIV0gZCSC/+wdBdDOSiiI7jx
0wigVNka+VFufAold1ht9Az8y86dOslhMKdJolbzrBXQN1i72UqDM9HAhsq6GKY332M/3FIagHnB
03ahJ2uViwyuaHmEXbT4KhuldxMvXl/jKwDtZkbS8agxbOGTOsLNfsvgJ8SAnjvX6hUAGnCdcWIx
8qcekzRHFulcqkilwXVCPf7f63+7ifk7ixGj/pkRyHJvUxoD9GL2AnHg8exC9M6IHNBHc8KmrxKP
wWv6L2yzeqLWSeVgC3AMHJng4oDxjd23dm68uq2cNQFRWdSkQhbFlmed/PEiq2TdVCSoAGgTJ6So
cUYmp2dD6H7ug3A+ePPTphz/+MOkdsGNUlFIiG/Z0L4cW2LqEXbkbr0tQsulKKlh2bPphzKUnczD
HGzdzXrgJ6U9T/evN5NMXxS7UyEXGgu0OwKu84TJIRerYsq9W8vmZJnwapD+x+x5LHfTfnLGKyDo
msm6p7035cLM80JKbZQ+NAxjeKbl+L/y7ujMaXJL/XwpwXYk3a9OhqhMTtcnHLJgfoF1nuAc6r/e
OTv52ImV4Tu+o1rRVgV9VAoph6UOcFazOepHkSQuh/AUXubwPDadDTf90M8VTZTD9Mt22TenW7dw
xR7Ru7/2lhCA1zxpIX1RxKSZzd2QUQu5OMKetJYTLoCtggdj7vaM2oBdP/423NfgkYgwItmkx96Q
/p6vcaDR4/fTSsA9m3CoSyc6EKicsWpawV+4HDYWsWsxEA6no1idfkCKhm/00xyeXAm0NdLzQQD9
VGzlmx5rm4jaIbG3EC66Tl8Qp2orF14CqqDCH6feKKNPcJKCW0NVcFG82AwXyT+KiYRh0/rwxWJ2
tYQBgUsTeKNmQGv7ERJBLNHAdMW2ZAIS2AfH2ANh2UuIhcuOV28KUDavVsPTVd69eAFEs7SoXLTg
qzoeThAVOOZKin1xzwxixrFUNuR6x0LODFOcYeoYI6oxYhib1iRJcIw3pgAyCJjvsb9fZPtkCC2k
LxYi+jhLmcnxOPi2rrxOzmGQzcsKKRpfbiOlcEUNHXM6HS5+ftiDeZKAlsfV6Jm3Bpp1FGQMuUc8
f7aSCyJCVNOmio0THqMJSoXq71IIy7qguhtTDBDhY3E/Lam/1oiArkaZ2GvdcK12Zbl/LRXtFC/T
fw77ZawxzjxWlXJ1RI4CbudBqnHkYOQXVOpY3Jg9EaSgHBlwvlWeF4Gr88kFJbvNHIj8keiMokR5
07iA8kLSNHtM31H6uKB+HtT4qq813DmqmWRXoo35IpHKrInXiF5iU67iJLOYHIbHCqpVKwYrlhfM
L/lnuqrAAVuhu9vOe06pjwiMvZ38/kn0tL8TPEE2GJReHLfZe6N3+vHo7tUpBWj0wA+ydzrehZ7K
XHTnKU0WryVMZdG1aZh3tk0ivxS71sAwagAtdw3ZpnygrPdwHHESMkMRmofN+WBPAPaUrlZeSKqB
hzcyLSyCdmU4/wN82ATkpVXW9IqLFnjWbi1aVp2nFMj2dUgscu0SKKquNkFV9s9oyI4/a4AVfOQ2
q+2i54S6zWoHw4CTN5YUEwz9ys/VfXTlb7WJNSWoImIjGAuL1PipgAe/+dV1LILWpMDBZDJaEJzP
vVaq7JXdHHEEHMAMhF86YT6xMek6rdTEGNU7UZJSA449sNw93mrmc3l/PqehIZGM1xpGU+AmA7JG
jypW9DUzRt0TR8cT3/h37jxrS7MNhT7bSJWbkMJEVF5nSsvrRxLLRj1dWU6q+U+Ge8zq6yjpjjuR
VhFVQaLm1ZboB1ogVdGjZjrDCJGcVtAlr/2U56SNgUI/JcH/nMMldo7F9SOkaX9rBO5GQRhzsVHn
smhM6B1gjxOxYBP2BZI6Upc9cB6f0c/6CoQ12ksRl5AteSW1lODXfqQ/W4P8hSX9RKN8qZVGTTyu
G2PU7F6NLI4xIdxWXjK5kglvfPBAfAMQeO8N+nyeXde9XHvYKcGYtDFH8V53MPcwJKr2ShCV0VmE
YlWOEoEK1+nfkeizyTeEuYBY6bGfckXuAgMX/lyCUYGF0ALIrOa8DCeQ3Pwfe1nsIISPk212q/B6
YbRXYBDuOX4R5LGa4zK2D7NZ51N3lf9ZCWlbjlOPIjxft2SA1OHq9/S4gpxFR9HtBa5IlYHv3t29
aeAjQuUd0Wvk/yZ1Baoh546ZMHkH3bPyPX/Y5q+7fO/ny/VhLR5+we46hOhLTCLxbeNa4E0v+8wR
ikM6RRP3HDpaKFJ51xnMnN3vFRJgjiw1NBpPZmaXqXx1YVhuHA66OlYXEAH60SrEAoO/oBjTOmfk
xUCUBtAEna+ejzUQm39UDnEnbW+1FzKyA/Hhub+mk5fVpzxlf2rgqwqHzqKfE/lALfROLzbPe1vT
RW3YEZEGJZnc4TvbDygv+E0MPlSY5r42E20g0UO1UOo9aMB5msnDMBh+nTUf7eh83zmAndv9SHMG
nrQM1NUz5iqQ8fgi69EzTF0V0B2C73bxYiB3ivJggGnP1lYsE5sZ/HbC4GvZYARu+53mm2U57G5h
odrRcce2/gdaWUJcladFYcsKIRQI77skzA7FZK76ttMWbwkLM3e3wvStIhcGjo3CcC3B50TkFYZT
RqIiAuFtHy+bWm7lFi6QS+7IptB5D43SCu0PaiMD2CR66qSDkbhyhGIhFz8PeprsWaKZbNfCqbeS
2zjsrBBrU7+NDRvwmzTDsZMOQgRo8jLlW2jtCtokcjGYLcEENru8O6EPSA92/5EyNGXRkuMaqRWJ
QKvx2v9/y9YO55wiBnkmi+jCg8ENwTkOBGmZiXFscvqUmkGk3P7b/lFXtdABFJEk4cLJzhZCLiav
PsRBdj154s0YCcp4uddH0kt8gd2q/3m+QvzFJBex0wdW+HlbwGHeqUBg7xipYiUC4yT56ItZs9LT
Q6am9T5s9L3M3HUvrKZKzswjaISXoPxLRMwOGksf8PA184dtzUUA0E53PJZN09Ea3NsKwN9kaxVd
ZSujDsFoG6EmPuoPdnY/gsUX8kRmpBQwmILqXdgEy+hFbM+v7L8C0vqiPy8uSYIFxTjaK2l1TbSy
ojUn3f4jInS6krlMgjha9aSpJwLs8Sd3uddJAZsmRhbtuZLF5+1B3K5U6KxCKjw+jL7WKoqBE97+
zvK8YGRMUQ54Q4qWMnc625K47nmp5zM19OhVr8C9rRRgtzMFlycrUGYf4vZIt0D1WVElglTmbzWC
6lIOfpaKqP6NIJjdxPCTcKsWb1LPhAA3X0EbrQkNBG5X+SbTp8DiircssaXarHNtyYA6YLdCRU8M
X5IPstyYXgL5+IorLVMuLqo7EBlzQs74j00KAlfZO29mJD+r90Paad+HaNpI/Wgldx0BVNqL+V27
FpRLoer5+liRu2RAxgIjTV8bt2vQoKuUBC0Ux/TGyAn2vT4cvFulVv9x/mjdCCQwRYkACCuBL+JV
VZ00AMRUZVWEcvD/mVnGuyddF+W8t7j1Sxjad1KErHdZ3m/yrZpqWylSTIj0LBWxQi3lZ2G1G4PC
aeq5sHKZ7zHi7BEECS3G48IpqXkUjKTlHEmnV1Xh0/szNQN1s5orDoIN73nGuMKuj6QZ7700+PDZ
neIblGX5djOb7Ey0NhUvveZInWCTMTza3ElGrkvO9j39MaNj/+IyPus5oCJ6xhd5R/IpEgnVSp4O
g/+I6aJY9Tr6VRB8XdNQDkC6xhsciFK8YcQnKktMuND6kWPVk/XfjDJip3p6Xx/1kaBQFNsszMRO
608Fmx5jPNtnR7V0IjntA7QeV8ZMehmZE+dPa2KkDhKDWwFAjqwDq5zKHmbI9hNJIJ5MNZjgUKdt
FpE9kBqOVGoZW8c8VG+YKb5eaLNWsSIVUCIjT8aBSUp4ZZ9qxrCmWPEZrYH+Uorqll+pvMSMp4Qw
+h68fRjs26Txz9bYsgN4m95ENxYOeDj3HyDqfTGtE8oB8Z0apdOtYlIa7ZRcPPHMrPsGv3guWldg
+Q/O4uv7Ap+y4MHL9Vekm29hhoEsBWdbAwvHGMbdM4o8MCoHoNngS3HpM6nP9jaI71nZXPSBR8Xr
Vh8U1JFAcWBZL3WXFIzbZRfFQt18dQF7XZ13nGgg6KCn+iLF/OdkLDv/tjyummsJKU19uuE5ZH6O
O3WL2fquGcctMWnWvvW+0lCr8s8uxdyj3AXSr3T29C7WVnS0Q9HazVfaGnXO13wfgVHnIZJ/VFH5
MWetQY3cre5jI5/gN8hL4ngbs8d5u51lpuZAZUM75M1Bh95C67++1XI9Lu7cnXL8G6VBIIFug6EV
YuZiC3kHn7ymIRTW3DwghJCcURLgL6gqXxZxRUk2aktaV3jgW4lhDymXE75MmlSjk7PAKpgk7nJq
qixJ9cR7yW8OeMvtG7Ra1jCaTfcMw5rAOTk4UY9VKmSBYuS/nz0+fs1Z/gxkxnAzfGtLNSlUCwLY
UYchAuV75J4wZbWkMm862nQZe7ZTiHWIztSXsDJ2wd56CQKZEs66iD51N+78oghnsbYXQu/wE1+3
zPaaRdOWEUSesnXtbPRIrNiuCwN2NHbBahimCTQwRNg5Xecb4cspSAiCVY2F17kj/7H5G2GpmgKP
yCszqUzFEk5DtRjvQDzl3LNbw8bhL2QEoySP7jUC6eCjN/Or5QTDnx9POsbSOOwp/YbVeILnqoce
iJfhpG2iTUkeF6yPYYm4FBShWm4eqibM3lmpIQ0WwhUQo0wS4UuwD03FORUkNwON+65JTIfxNZ6x
oGfPxQyE0KrVQRgTSAaVCyfyF2VZtgoh6iPVsUzo84gQAnrStiGcIhUI4y5eLOMJsOegyWygrPZa
VYCilXflIMVi7BfT0Nj0qszjV1khFS05cCXTrt3HbaoiuA5SX5T1+wD97DxeoJAXpZUJvThLuQ3i
wpmBB1tp3hWIVGln0wAVipzHcRQ9FSUq9UujtJ44se5Ht/WOufPyxfRdJii/BMkMRfpEPPzg8C8L
c3gHW0W6YodvWmj3MHHNuD0L8CwsykMcvIUals/WpuHZU5/EEX5leBy++hKrqSVFbvDOicgP6doy
/h83rmymIdriUFvoM+5trxVBQCVn8hwOrgtRW6Z4uyN5OsYMic2au6Hax+zPcFCiHF8MspLLLAKE
qUmQZr95u+lJ+XppB7u5/JkoRVtXLccEThNPaMiCuDei4TKPHuRYAc9/9lBTuNAARF5qekcRwtuU
v8zfB97AcwJc2kutG1zl+TuzuXtGb81xZ/8JEMRg6ZwuZFeDpc3M8J8SIej0o6gIDA8GrgwPpteH
GKBOFHBpyFwmScazO6C+z3ZG0BP7/z+T1sjS6AjZNay4WT+jFIFTWEoYrbwdSgXMe1DNK/ACYgPZ
VC9D3NGvNCWOZbQOXLF1Y3ZgybJp1Mg9QffxGZfMQSBFst1u3DQj3qYvw7JyAxQ8+MIDZH36QzcZ
tbvNXRWttP34CPVFTiZL2TtSUcMXPK0RRfGuwc6bY+BxxFVRCE/eCxOVKHtqWBvt20d0ifrd64qd
Mj1BaOwtW5adygQnDEwzovy40JDJTkeglHGsz0wGEttqfD7N6Y13G6UrxfDd2KTM5NSfDjjfr6U5
B34Awks6S3pjlWoCQlXG06FJm3l36AEYHiDxHoiEOkDXiHjfZWk0UkK1pAvPRZ49htzMLV/+8xIB
Qp/j9k5APWfE8SAlYe2keyyPrjKOlU2JPNtHKdMEaD4UA2tjNcMf0oE1zFJrGSPsknMcRtZx/3iE
ch+NZf1fpNfeNrqOrLr+nTJdgw6V37T4Lv5Ia4U/GEbdQu4PWx7Nlw5VbokvPo1voP9qQdQFs3wK
H/f2fVF8aV8a9Zd7PD3kCwXznY5y8egO4M2NDQXSPpb1hUyLVCMLTaJZxg85nC8u/+krJuNgEnWc
HYU62qDXyY88HmEEyLpIftdzKDitr+rWSF9hlRf/jtkp4MzTjh+lvAaIHPy2aeVv3QPyvaWnEkuu
zNJZu9x4qDfqttUIP+WLO6aUHPWwJsp5dolpLZKWd/OKbOFfDq6CnBybl0EISe+MFDwrH7fbDzpU
AxQYKMozyf5cYbRMbBJR+VcsWsQ2uGgSwVDM9bK0ZA3QAseUi1uaoa/0Ezwq7lmMum1V1Z9ikajw
ekOaZVSvGyc40Fp0awxjfFv1BUDSq3dqh2Ac0AzQolMR5otnNOAjzg7QeEP78Nr3dUEy0FNU+Skm
DRyvVSTrvhE642+rTXp0mlkl9RlLEN6i4cFLuILfQHX+gxJrQRy8Zl15c/EGDkuIRZHP9DSKPhhm
5IFCVSi/+Cyy+iUYL2Ai9na4zLQvucmYk1e80U9a8s1cTuHTwqQ0jVJKDsjKWk973wyVcWxIbz2t
sx/yxZHDW/NwtW4d6tn4qX/MHMcd7d9SH6vxgOe695dPwJYepQbC0nMx3NtrgqUEnC5+KDTrUJ6u
kON+aGSh/slwl8hJpBmcRE1zU5IrKr/DB8cISQyYZeaabfbP3S7hpgb+dgEm2uIFh25TpKnF0bTu
gZlJ+zzsvA6vOFms0bGLCW7rin/+JDpIeg64DCaKKxIzup7x+M2eZFULBRL/h5MPkSp9jLhxPtcI
/6vFvWSx+zqQ9yXLcjJh+6ba7U8vefS2BVTiRMWhiXuDcimRXdREoPzL+jhGPLS9CrfIgXkHu4X+
o8g2vzIUEjmSRZQr2rPzhutFQ3yqfRmpRIq7hmb/m2XxdqiGn64r1FBIdQprRZV4+vzDD9vm841v
cCSkZkxmcz8VLQvfBW1BettxULY5vzJljpbtpS1bl4S0muIVEl1/6eBuZR4TQzS6dIsjWB2d21rF
Y3c6jrfW/RJfcVZwdLUFe0f37OQcn2Xcn4Dyc/JKvDhlFo6kqEE31Q6jLoP8fxuOUknt030NZ+6Q
W3X+PxKByqf8/fMhw33jKNtJYVqkhmGle4HVjXxhsUWA2VdnBaKKu3gA+EeiwHmkpgVXbtYO2McM
6qDMMEqxBEat+RTjyjq6MejeB+QF4yV0cLBxix7KeDRZYiu1BZiNkIEC83eYDyxnkh0p/Mr4uz4f
1UfbLaSDxaq7LEMJ4FEzYJSGZ9oYlxXfKEzkazrIgsAvVMgtLlk94mqty0oajdnL75Ld+r+lmiaX
mPbG1wk5k/XE/B1mT/9n9qDN3jMFi9F9zFPqzSByFx3Bvs+1TVAmrOdE2iDUwZeEH5H8Xbhsa0Yj
umGmH/W7G6EBmZp53YfO6AAV8b8OUyCDoxZ6OGJ/1m36fhGQhHzfT0TIJlbFDpPnuEmIxynvoaRR
IaZ6tUp9OoGMhPCcvNNOqu+XNnwpB94kGMxoeae+W1a804lasGe01Vvww42KCp9jkMtuu5oCrcKx
dk0g3yZum6VYbptzzu7NmrIsDqLPFiYJW1Q3iWNepad14j+45nZa2nmPSHY8PdLFoSN7D4QxYfqA
h4cbHX0xMNzF+/MoMxwUK+HulrF4iWux81Jjy5o2wnkP/DMp7Jd3Vw7Q/IIJKXi73j0t59ZTuvao
JIHHLQ9Rn0xmLEIjd1Hrf7rQDqpji2odHzRJEH7KSuNMFZujcO399UMsC/bNnWMQiRuEyrWmLZ23
oyS3j/DYwUkRC0oNETnygxps0Yu269pmy24mbc1kmx61HPf9PNuFNCBN4vo22qkMM7STldh6YKaf
t5XlU7qz1nJEx8x+Z3xpDgmWSvOXOjzdwP928Kgj+farjso796LLLcfiQZlymRVCqTyIljyzdNb8
TgGJckRd5TCtZNoyi2t3Zw4g/+Plo9aFDt2DFjnrJRZCD+julhJiqvD/YNLhkuVHMiJOlVmHEnhK
saUUqEzrlYeFdRfipX46oNUAglL12MG0Rucae52y/nYVoVIl6/CpxEdeMSvInBulj5/Osskxw306
jdup1O9bOFsthDUfTnRO1Ko/nYDY2S8aPVH8oZWXohRZOLb+wnsywUpZ2Ug/xWrdAQEoKI+LdoVQ
F01WzdSVkWls5sNC9qnjkPnVQKNp/CzAGHTikXKyXG+rEh/HtQsKw8NxVKqyZTeodU4Lbma3H6tM
20nB9tUyFbno1nf5pkMjxppzlZYL8vs94NmKk9Bd9WBAV6yLS1tzjv9bboZq4bD+sID3U5SFpmwq
M6PeQmBc3wQyTM5P3JuyLThQp7n+ru7THmGgGXk2Rpr34i/5orvokDf+2YZsosGF5hy+t/0LYhzD
NxTfnVUrcTG7TbqcRc1RRCzoh83g7cHGb9+YvbbhQ5/hmlObNmhwt+UsXaJC+UU1maM5goD5hfKF
GskuHA2beoDwmNRUEXsEWUnEKD2d7hcUuuk9OhY5Y4IhxIq+dOL7tdZalWAXOepnhRRCUPk69+RL
Tp44nq3k/Dmndc2BL1y4rQQQHzlftN54lnqwt6ZJZA0I1B+0oSrmvFeN1ZhVHksfg6d39UsXqYSD
ILS13XsWNIf93zvof2FTnPHmQgoptpHiDD5b64tzCKXRX7r4Od86m7zMYVh/CH5zFEVbfH0/oN14
IYGImXT8BT7Cv1Sr1HdiEgp86QFWxRTrV2Yxk0gTCeXFUxfFAx4Calh4njTpmH9yURpAP6Ddr+lX
3WZWeFVIu9mbkGmkA64tPYrVS8E573GoJsghl5jMfTeEEncmFjxtl0s+purL4sSUUw6KhyOnUCej
qJl8whhyjQOLU/9s5Oy1nHYTCMElceXtnrpxm/+M7XuUrQRySnIcGOVhVUC9wffjkjvwkoFrgsFr
JERViWkBTjk6JxWi+cGfcDOsorxDHESum5OxZmRe9OyxrpIeRbuSUYH7jCl1vp1bt8X8jv7xoLoB
2Vo43EHIbeHnKdqbztL41GtnbGtC2v2xrXpIyKzEltg24jrA4KWeJxUCrvgo45/Ony5wTr+SRbuN
OeTbddKqAQqzaoRbD7pFb0Mf51Z0n6IiqCEbjiIRPRU0qSYDtFELCTW0T53JBybSz9SzzeWXio+9
c5/yklKCLhYcWtr/ZtyaIfxKCjvog9Qg6S53iq7Z/spP3MO4hTZGDocW5QRtjPXyS1Q/oyFcOsO/
5X7vMo7qc4HZl3Djt4cUdUM5a6qlT6iBqWW9tzMzlcSCN3IEs/JhGIV6GdpBRCMAun+vflon337l
mAkEDqpNup5ZNLIAnnH38WhqeuEayraFVU+QnShCtodGNcHTdK5LEY0BLdWj9Dbh0WJSAo6GbCH5
cEuM3ssUzpegVzMciYsOrEtB9YN6NwiUaA45DNHgOlu6JR8bfSAg3ZFX+kP3Z4zzGmtYRfRYO2YV
uh5dYcIHW6BjlWL4rOTzB4DXmmYxDmjZnsp4lKnqGF+qCUALBMmznTndrRuKAsYeK4ynVd4ZSl4a
2aS/jy/KAlRW6qaux347RXIWKZ2Em9mzWz7kJP5LJld2t8p0oXyMfGEtXWUWuLoogqfQhDuOXZVC
7x/kV0AbHeERZZ0EHYfHUlNDJCgy9skB0/yPzcGmMWmRHN7le2d4cn0QeFcQLscIDUu8bnSfMAZU
L0rmbxXDAwuTGLk06w2TEZy7yS2aoRHTrlO0TtBKEpNpPFKE3vqDPoRxILh2yFRA4/3e1/qL2hmJ
YeGVQWoebVQuPRtT1/Ap8efx4E89MXXIwSbREz6bUDQbHFAk3dvsYXwqR9+FntgF4cPcBoOYuAcK
YhYsq5btKxGqTL270ISsl3FeUwF9WAkjH5eVV6U0RDVGIRe9PnxTGvZbshqIoTI16qQ8q9aTBRuv
mE4XSJrTuD5m8rGodfCYxMmPD6HqgpT9KNwJq6HSm2BfXcOMr2yM/FeBd1VvEfmhgot62s1qtMhP
1kZT6sPUpQQHrkGDZHeZNioHm+96oVjxs+76BTLQ6AweP/pBDIn5Nhxm21AViapg1p3j+0jhVQg0
Ac7P+1Yd1TVWaGrI+0XfFKIMIozK/ot8GBZa0s4qYDTZ3D5R7KHxREihs6Vs4RKkl3IrdmKepiKQ
4xuvm6pMocZcOL0oKVdyA4tRML+odhP3r9grd2VSvD2655uetiDCm+0+tg8QYclKy/pU3BGFdsIO
CUHLno7rO9mxrYx2NILsufnTFz0+Rq0jL6LV/6OOvvSNUc8qdQ+9mvzXTmGCUpZaQVfXs5IsHVLg
AhTREXibUBzJMBxmLloMqy6EHHvo/HPOFq+tG2pZakEwOTF4hUszk5H+dofwPxZFzFKUL9qKzN7f
cUbRNfXdryUu/+8sUmkPz3wDMYTAsJfZ73dvZ2d6o9C/wnnxm9wPTF9NA6AR/bvezyz5UCi/rvq7
kiZjNJdSKQugDDnmvyFq/2lknwtbV+oQK5OWEvYv5PdsXW5q61/eWWBgzDj3iNfOS/+jEbLqCl8/
VLk+uGegxCzAJYzj2VWvMBHTNOlXz0VjUhYOOYEgyorWmHxzmBXupAkscWx6IoxqFdR31K/UxUEK
gGcIh6W0DH+XJkChavmW3nH/WKRYA8QYKFxTVMVAVgI9ZHORzlJtgYwHzJUa9ZehNyy3Wi1//+nd
Vx38JIAIuOv2nyWKs/jLy2L6+BdVjPgZGWPqIhpxMS88qbDjADdt+ySzi2XpolvI81SYQVct1pxb
n96zL5OYsVIfE7jT1qPvM2U7JigPlyVms5baqqevq/kC5WfS/6g71Ww+Fg6EyTl0PK4UH6nysvk3
FQAr8nNfIYJBAVDYDveN28mA+2d/VRfUgOdrbzoHDFa+uJ7R4+BHyXN8al0GlaMK6w0pku/L9Puf
j4JZ/C827t7WlUNBU2zYpZj1B2XPTkn4RHU1IgKJChd0jPxUv/SoZC1Ih5Ru0bgX+nUesf2xDkZ7
uxtZXR4Qf2u30kuMkx+Scog1YbGsFnqdf+uGd6LUBZunESAua2FHu5R5L4ZEYkna2fR6d7azjtyI
meaeuznUTcfgU+uU5ze8XcSpPzOQrsF6hszrkteK2vKsGMjWrHPELKkoNteErK8EWYQTPvygf+Da
MUQbNEAhM8rpXLI+Bdtjbg8cM9CdZw2LMFiqXGYvkJX3dD69IQ3NoxCTG18GbGcYS30KRi5Wr/xx
aIgtkAjlcOEYMb0nMgyV1h7rs1lCkG9mnbKo6m1mIHZ8cUgzqTqU/iZ/G6LPXtROa3ggQN8Zpoe7
mELq7RpFGRiWgR2olLj2LoAn5SRgmilTNbzkiB6qOAiSL7030rLdxSUlHATX2zmK9rRbW7NcV7Gu
8f32ybtTteXF5MAYsaqXqZpjHu1Cq0qiG6/unl77N5mql7wA1MpXtcLhD6ENqIHUX6eOQfYlHVVI
s92S3WTe5GVwPi18s+2HSXI5TDgYGzIh0BtqzLvg3OmffvZW+RSV6b1IkYWFCAtZt1gL1woWYtIw
qQgkJ2vRqvwlMXrq1GJM5lgqbcs3aciEt2qBMfcCh9faT3IebrNjaQOa0TsxY+b8PkUTskD/JRrn
1xqqwEm7FZIzdVtjukmHBG9mBvQ1BuzABzzX1BJf8Y6w5omlLtFDz/4699dNHaZ2WvbKTBvN9rcR
l1XsX060CfWV6x2vV33gGLEDG5Fftlo1nnXVpN0n8iuwfthzwkmT7RAndMgVtrOVHBO61W5/Zn7P
PTZr1yU83e9/PSuvp2Ba0VX9Hu0mEpDuT27wusiiyAdkTwc7rClaFLqlkgPgk98yIk9530BcCqaw
7Onhi09zbxJTfS82LKRkEol1JVhQ5BiWQupZSUA54RhxpUQ3qAMQP1MO1BGQZBeomZJH4eB5z9vQ
DahTiFeXnSkep+/9RLFBYxRp6hvvp+TNeETYGhyDCYG4CicK5KdKDiJOn3KVdOFjwsL/HmBHdbfY
Jodo8M9L9wyXdEoclzlYg48xDGQgKqYUTncqGhmfi2IC7mCVAP5veZT6MNPY6xfGzdWhJXL76s0b
3Kq/Q2JK0MoKj5Jx8252Beudkk8E6BlKj2BPx+9nIg15xOxfk7CAXHUyaoiiB5IqBiAVOm/L5EZ1
xw3vx+myNTD96JUjZUASIohgE6rMQQwQ5txIlKJG3WmEVCbQ+tFG6U4txnbXn4YzGheORUahSN2r
hqlVRtZNd/gNkZ/K+Nd+Mx/eXv0Mp5Mif4ZMWQboDoG5PLqaiTJYKnmmZlyol1G3eh6gW6k+dI3p
58x+d+3UJOyw7EZ/N1AkMa9Rc7Rj30RsYX0RYPTL5g3CKWfTqbSS80zJVGInkl8Mr2BDjObG58cf
buDISK4W1oifPvOLQnW4h66U8hwBb1KEjr8XVRbLbinkpiK3yRTT8chj86gOR4NbqKzoobRsQ7tX
v5dHsNTPicbslPKgIvIFeqYRYW53hqtgWqRsJHnJVfozSU/wFsQNrZCTkgeQEeiQfM6Q4e8TEOHl
o4Qc+8ve3NwYjL2A0jhVcOEi1sT9FTWc87AebtmwgK0+nv+FzXVR+XowsiH5rTn05jitotmpm2EQ
VIiRqEeRM5xOA85gsEmZqCwpIZ6lfgpFZawwD4NEe0/K1/3kRTOLFhqWoOvzKZHcuQSHcUBgMGc2
aHCM8XisUIee4K31J98iQT+Ja3Ykt1OqvthU90SpN1uY9nReH9BmWLl+OC0w7ShnCI/shZkBVcc3
9sfbxMgG5S9G0rJrB5e+tVi1wlICmW0gCTMjCL9YqRm2CPHruDWP28+IVIrrNU3V+kIZO/1WoH+I
fBS+CkB3cr/xJbiRhbG4qEr5Nq/T1r9PkNu3SypQNqqLMM0PcJvnt+CWhvMeyxqT1DcTUtyZk+N6
dtveiaJ7sfZbV5c+rJHJeVGnP7YKfH106UTbgixjBDaE3rG/C8c+GR6j/gh95RV2WdLbM1WlGHw3
0iPsDiR8Yz94JjoXacodDmHxvdLqFL3XWfTrdrufAZaYdg8sIxrdWUe00bhZzTCVzn9unQAfVAN6
LxaqnV1OPvYuu5Z5w/T1a5D/jb2bnBjPZSIwdnHKY10nL5dQ88tq01ErW/IAAnJsYOtaLdTfib2Y
4qRj24kCL8YrjHcs1aQYKi9zObKqxdvzy37VgkDNpFSQhGaxMVB8q+SyYnZrXRPE6NMzMMALL9hr
C4nVnBCenUt2khbPKwTxzRh31Zuj+QJG/BdWztGIZe8hC3CPdKNy85TPm/zTOtBiRwhrMsHoofio
Xa0rdstjjgiq0Vc2f7Lvq9WftT6MSnSFI7u9r/afcZjrnQXrY1wQswF7Rryoq7PPLObeQKVnr4AT
bVGvI7QCJJsBXA+BbrAfg8joeLspPKKA3WKh6sbgET4EPGq7RgTzc/MiAPxE4QpApmjLWrnyj7zH
3xEEUSOpgFlKHJoOgGwCQmwFW7bD6NUhtGgByJwdJVsrFse5xb6NfqixJuZDw3PTwb2kgC+fVwky
FTAccz2G3SsGVarDraZS7TUZUMjC4BUgSreHmJolUG0tTAftGoVuyNHi3SlGTzaqh/ZpRZbio28q
6VgcoWNDvlV0aJFPslNxVrv1/esZTyJXlBoYk247yRcIFXWp9WKYb1oA8AiiaZpFm2bEm044TAlx
V/I5ugXjL5FGsKgobPhF+vw4ENk0gXl6n/PsMgV6iwVRppn5yLSFsRk/zXHu8cbL7VPAypJ8cl1F
jHP4SlMNHCj1t90I8bYdHRqDTHs/bEAln5dZuw6RdkVoJ+RCjTzecs2XIhqSZulxI5ODDCKvHxBs
p1ODdxqvXqsjNCu2ec07EZV4mb1nushzgVq3yk7nFV2y0Ul/LEhmQvvMQ3dTSmH2NcGo6oa/WSWS
3cDSszNrAnc+gQkH7pKd3QXJphGsfZPOkwU3x6yrF3tEsamswArGWoIuW5cXLgYaddeP8u0gHXrr
Mlra5Gsmx65s43njN9Rcsgl6ZwSWYYvqb9kwoW5JFP+9/apeViadLXlvhC80spj5/qYP1rmXQMnS
R5zu59uYfubiQE7jkox7TBkIKNGB9wA4J6/lFx9HzlJ4zlTifaiAKSFUFJZwG+Vs0yXgCGLGyIpA
P3pd+NdcBq/DNf32khAsbB5+OZAWAXjo4s4JTsm5pO8HSP1JDZ0bm8R/MB9abH1sc5IuhXj1dEBr
MHa//7dh3TlbkDC9OhQ/j73KdgVv6c3G7+F4QGLBB39ozyFMShHuQcQgSWM4kVSSlI81MqvmBhe1
A/995fgHYHq1rnqDTvgmsxHQEVyQY7VKk5qrNO0KzFaAu3oUSoNO7y1FTKPwCUq7IEGaGGhHaR9B
EiVUfw+nUltOyDBhpr4udSZYcvoW2oBmxWNCgOQLKEDgk/XPVDmi71g47IK+C2J7jSsdf0qswZBr
VPyIqIXb6FW5VfDc6IxLbluL2lYBVwkvfyfZVy6twr3s2ylltVorkbY6iM7XlYpyNlVlExa9TE8j
yJFINqffeVBOQqIMIyk+el2F/Ah0jE0fKhWHxiR4XqBWDMpYFaVbZa6QLCissGxRec2hmzm3Th9A
6nbx1Qut6epHGKc5flDg6m/pPgRmBHTcAfHdvQdq0pdcTqjMwN+JtTxS1UqprSm8Gw1KQ1xW5pl9
RSFGB/3eVxCakpb2NgnL8b1cJ1EyMLq9GN0DJ+4CqU+eg6s2pcQWJGUF2NwlHMto5o/0uFXoGMfl
kpTGEBSoe5jM8Cc51KuQyWJCyUG0ijJ3jGHYxb7TYUqG9RDKbigbhTzoShiEZKobDDgpCz57gWFT
ttW2O+xYE2HpqrHNTgfG+T/xeP6R2PghjugNxcN8k/Yk1ZKjNM3f3mNPBxRV2kIQudvjXClPM0v5
SXf/u/95cZob69OIndMrESxcwGj5+DblyAgKvAru60+n4HlSDoAGVPtkH3iHrVqGb6xSY0eY4zV/
dsAhpMWMTRulzQp2i+uKwLKOojU9os+jWUR4Fea7qwlMWDNuVar9/SVVDzq+W0W3n4SiSIfvdBj7
JNS+zRYf8atTTGhq/wXApNsnlj9i6RrUU8r3fZBx5R6kSOCSuYfsqG9ylvuBMkpZl8Tzc4q7H53X
7Kaswwf7CY0daIhaxfuWUM6sWlBZsktIQx01dHswRN/o/V0UJru7dMINGXOg7kbiy7VCNUYlbIAQ
O5DfMbTo9/yC6H+yfd3vDZ1Hs+GcBd6qDElvDDtUewylDTz6L9ha4LAy9BjBNXmONLUNlknODUVE
7dICMcZkHczMRz5kRq1NuBXTH5ej0eaJN93qsCT8s24zK5jjik0HcAlI3VCA/CNC+c3XuS4Mh3KU
EfEGxx3JZbcbWsT9D/oJeF8GQGRUiRpCYBbasXM5icHkKQbPsOoFrZV86uWRO3B0NHQxKDiQlxTS
W/3PWgZapY1fAMHQjCP6CGnTsHU00Bi20lMaP0cs+yY3JVfOBCyLbUiplBQoAyEcQRhBjJdjcTYC
jQtk1L3fESmBLurTgM1CaFEpmqgv3oltYfDz058hUGrYsCvYvmQZfUOst4JRtSpLKBCkF27d8Xl0
OV2FG22i9tyBsNB4xilbw4Ihl2zALJTA8qqfAWD6gtCGU2qUGVnUE0W9bcZdftKPVaTzvLD1hcWU
+HIIKhYN82kbzxOnZ+xyrjeF+4ZLZj6gg9WgFVDtZ4KZZYwbq2x1hX+j61RyAjY+N33bwf8bAc83
vSh6ICqm95afbx2k6T286CLHPD0hHv+r4ytdhW7ekV46P2fybnlPppAAVgPlfbsVpXXDzOR6TJ2M
1LPUdsnXQGf02zHw+kavZt1D/BCCOcUjdmsUvd/zj2ujtL0OgtX9DiXi5K38k4ovU8NC1g8R9qgn
OzA7ZrDqM03RFKSWjw+LhX4jlKIsETmPMTvIzoFner2x6JtXirR4BgdAoqhwc/J8vJNMVJp84MWg
kY/vPwYGKNp1R+fbVaVRzCdJ+Wpz1d9oMIgKKMxz9GFDvDS5hTLI8zeSkOiTjzkQ+USi+y4a/S0v
yMhi39KGS/lsU6UOHePn0LEi2gNkAY5PHJErrBFyNi1yKyE9rWKjELLdH6K8tCmlBejOVAGyn/tK
jr6QBMkeDhwSXNNpnyP/OYVrLRAK4+x13uFd2ko053B1peJW3qDmeD5Q4kNXv0SrfNOeUrFmH57d
PrIFi0QWJ7prydnHvkjjrqUaHsWlMco1ncc2bRm7Pn1pa6TWfe+JPZcUyvYIek6lQtsGqwkzuuI+
p7IoKSGgw0X4fXo5iEII4P9hsT84TT+t9KaFKP0FIoSZglR+liiGnBTXU7jDu9lC1Npoy1hshFE3
izGMXTq3H9o7T9fJxdlvX1g54lYDNwWw1guHAlahPxWW6kufDyfLXnMI8lU9LNxjG1cUCQYbOrDf
/qft+Mm8Q4bdLfreoh1OkGhaJOk8CFfoH134DFfSXR+TmkvXV0SD1gH0Gw71ufbbVOSpAwZPef7q
C5gR05puQ52tliL5V4vaZPnVbMZsEuaBZiBKQZOrhCYUHZla4SszK98jpecM+wqWJZOpUmchekuM
mBD6YUxiGM0/pAd04q7dD+ihhKmkkUUNvvwXE72NG1T/FJBXUZ0BIooJTp0c4IAK1xsP/haE7cub
K7LSl1XH957BRB0S5VXMI+p+pQkREpCtzYZakUqxXMAaarI3T7eMGJbYwyn21dOHjZmO8WZ85g/F
MOm/RiuTRW5AdsoZHMEWp+2S4AIa+M5ox1cUWGxUjuoDLxLStPNJ+P9ujIai9nthi20lNRCcapSn
Rj8ZPuoYO739U/7nwxUrJfq2nH/kUW7mSvJunY2oHarkBq5beV6/E3dgQWQPemZzc0Hc2gLf+cLj
ZQkVL5m/AmNEG9W2EErYL+SDQHnWQx6kqYHojkXJj3D5K/c9ttndmAhXqF0ciAlZNEwF/bKtJvUS
i4Jm6X8W0wKI10HubAfbLXcr7DD5wZYx5pGCGPxuWwz1zEkiVB518H89SLVi2xNyOdW94sNPiLRv
EEnqBZb/xlVeMvga4sdHCnDvqwsWl/zGabRdFslFulwrXi4YwvN/POKsDLUc6HEDk6iDpwL+DYrB
Yw/meqLDKT3AT5zNkAlniwplgQriwczjBJy6P79NS3VwSZO1DbtAUoR1ja08c0k6VjLU4/CUycYr
bQyKL8lBpdMK8GFXRQ0hRVaJHLvWhHj1hk/TDSGcFr3RqNRldj/jn728K53jaRi1F5VhO5SzuxcV
6oNQjTbi0Pp1FE08b4NLZ+OnK19BejfpySGlhZmpKorsbjB54Liz8ve56wK90WVQs/bZQoawTgWX
qMR6jRBLXXFoHEoosLGbYtrGwx/j0Nf88EObL9MfJhAiOO7n7K59y8C8mKu4uD4BqWrnHxLaZQFQ
NZd58j+4gRCn+yxwacMBMgVvcC+wuYuQGoU7OLNpF06EIEKvyO/gWa/VCLUlVfihLWb9I/2MVatY
TvTDPaSNhrNYz6ZsADqbdwsc2oDpUArfncX0qkoAuGu/HXgwE8DW0bR0G/hqIHKGrtaHGpUiNCOY
Usy2lYcXGIbM5AvI5oY61Sc//A2CvCjczu75Y8UJH5xAzOLNoGeMYmOn7hiYU6t18PtE+5AQhSrl
UQKx8SzkV3GNNL2lei335pgYO5gmEyKThNcWeH3qN2ezidZN8f/+y+bhqc6i9VNpiD2CCUHRQBok
WG/kVBlN9CMaOLxpX0Fu6oM2cm0Y+VgRJr63X/2pkJuD+vrdlFyibvS2yyMJPg/Bx8UiRLZm66Ct
TTr5fD9mUVdGJTa1hm5gA4872/GEPud+Hx8ZgFDwBfW6Ei+/fKrGmSbgahW0pEtpkM5pWvLUeV/M
5S14QrAt422NaAkmydGjO62FA7cotaUuO6fwHrc68jVvl2DiPc9K7t3dFxIHf/fncG18zZIeqdBT
5LmMhzpN2MqqllrDTYaBzwKEZoWE9Y6ZXtQihoh+TAOx8Z0ixbECF3QpXZh1kM1OOvnDSvKBomcX
STkqTz9naZQ92H2xToQw7KLuy5926KM/4wdcD1qMLQbceGak3B7nNeirYjLzZDq2Z61Mjr/eJLYa
z0QrAzmAw9IfDF/Aa2loHKSGcZO16OiJl6VI6+h6WmZI9m6tBysT7IJkZw5geM4CBYN8lzgzbfgw
n8ymZy+1u3/a46dqdn6m4XukkKCiRp5TJRURX+z4HqKU9+gBrhLUxGDhIcKLUEaZXKdPIXJSh/dT
1elM+oFWiO+LRhFQFfRP/eQWPxIuX8VZInGAmw/Jx7WtsjgVTqxzKLZLUu5jmbeEitSWWmHQJK7Y
/QjZ6xKIYA5jdkyyfSf2Co+gqsj+UOv2Ku8dJeBkoP3rlA68tqNDhJ6jyZ2IjAozfEzLwqYYYFTo
GNFsBVYBsYqDbynTdcNiE9GKTHjSsZqrWJFdX4cUf7UP2QdVNis4TatLvwLWOTpoCiSCQUAXu1Y3
hdP6FFW50vI7p66qRzzeQvqj2VywHlLGY8fke5Fdxl+ytLubcHXsAihoiy7BmRGeV4gtYbdivcET
vr43+5w/S6Ai0RPZNPf0YhlTwSWm1aBZaoRHgdMzzuge3uCW5rFAFd6WTy1jjDwRq25qF/ldGdxy
nPYroSD12XUy9Ts06Kyjc0dpDpNiw+NbhbIE3u4EgxAdT6+/u2hruXCR4U7THrCf2yL1rnGUlQp/
g0awpC/WrUN/b4BvAdusVKzEHFu+rKDxnGeb2j8pFympGZDKITaityFp7WWlcgklL9w2rxQSCM3R
eXNnIEP7vEe+tVm16+TPQX7zeeyRwshLitia8/2GjK4tdKyHstpGx+qvKcuJ6KIL0UV+azUereSi
gjzBqEyjQmGZkzuDFHAyeDwtm4vlpK+5L6jxmwYiBkdode518nrR3S//iiKssEptlvIDWpUMxuDZ
GIWPYaPGw2Frw0rPpdkft8xdWy89CF/tU6qqlkKzr4BcesLTPoyMzPP/FDXhfusqnWrBkT98fD85
Guyu4fcSycT17ucPXYRyg3XZiJe/ZK+jsQPM6sSsCNMieJmD38HS3vHAJhQTuS8/EZXaD8AWZVcX
QoKVz/zzHxrVvWwKw84HxZqrG2MVebC5DcCuYJsV2V15luWRmXFWW2PQrPamUY7JShI2JFXNWXWA
vx1TJ/m7PCzp3ZU4pA2mT96owp+HwbGM8ScOGmb2vzagOJ9dVbPl5Ba9RneKpNx0gREotMAvhWiI
LWHVENf/vqJ7Q7vI8N9iBo8Q5jpH5JErIV3Gaol9weXEfKTVAoVDnlGKpBtE1pv1mchFnf5nwqGA
pAJOc3k6IfJVIy0bTvS4KFnKECcYkglbAdbeybfOfqsgXMmM85aSyEeItkIoygS5ZT2nm3D9+yvP
ljgqQ9eiflsUW2bxbGMqTGPaaWbZq85P1ocDhI9gcK4VlYgWyLVK79riWwHpjWIZkCJ+cDkRyRJO
mOi6i97i0CagqySSc5t2tD6dbYIP12WsGlXrg/hdLJM/EQ9wjJWI+MQ+B+59NC55/pdpuG/alXyj
Y9in+MUjQkPNM/otA5spvQXQd2ZPxYUFT9uxhMJzYXE5uJFrjtsLvU2CNdwMu2+9EQKP7zz3Uzmp
kDXdlHu9B9rVqjIplIaZxh4QjJWURn6SxLAPlQIDA4eAjbx3M1e5MyErmnAjpJKZI78THw16+uDs
qh+ETBoLX9KmXri6aDZY1TCvoOlr8nRxUBhghFHBAjsXPXYMUnBbI2JMKk8z+Tmkd33CTr0nzs6W
pW+eafDci+wUGrnWN8gz0Q7NOwVA3zWwZ37HclJZClqU4TbwF1ZQvWXyE5LWBeckaG+BhtAWYgxp
Zuj2N9B76Sapy9stQ7LdcbGIixj1/UuT7m7+RWid7IU43Q3KDxaiSwKN+pUKf21+kDQiHzfT9Hk0
SeGpX2FqSZ9bvxjajc99vaC8ZFSpicxqmjEWNaq25l1K9Ni17cAOzKXed9lpMCTeTI464huJo0Rs
K7NcvzY7YqjA207rGTr6gE6OqGcFjPQlvwajJpxJp0EFhWKv548MZqo+nSRcmLCHIt00daiJ4dat
DrHAsW5p4s1KnEeRhe+JFFq08WQ4IRsMTnJVWpvbU/GHEUs8mUxFx/Mpa+I3H/RS7B9vPCznMPtM
10u+HxxJqYBB0zcwvlNiRdBDaBQpGYvyJFtBtAdPWCtzDX07IXHFB0+C34I1V+q6s+dUsx6TB+n8
INqPVLceKnUGlMdWNcsKEZgqO52c3t++p9lqwV1j203bytdysf903oSktuG7yYoVNYoqFhFd1+hv
Ux4rYGF+8i5QUjVBzvohUW3yZtVoCd6bUbj/BocvCQdt9lj+Eru/N8pmtM3CsK/6RWrMReqFWkJ2
gcWWpKnOf2329CfnPpsXoaSLsCwx8yXwxq8lOPOtct0bQFobIrtc0VREp20vBzp2+4vXWnzmrpBZ
jBt6JIdOqnYL7e7HbClZfZ0PNr2SEpAWBjmFF64ffvU5jC4Y7IyiBzQw8ObvGmfSHSLKwuiIYJO5
K//AnZVNS1Msj28q+G7LPz8tT43hzj8Od6Cnjdf1/+kNlrCVw9OpISavvcYMu617fGjg3gLvw5JC
uImgqU6QkcMA5DJ/Xe/oq/lmdmah5YSw2BGDCx+tnAdaezD4u5vqqr1l/OHqBdlYtscmrHvU7WKn
ZjWsje1lqyKHSIr72bNlf45vjqoVTkPAQh9BEMlsVSbc4VPugilvaBVMaVlvVWMTL8OdoS2o4zIP
EgkKfcqU/UmGfwvzke8K4zOJsfK7tGHoTubi8eESiUvYdf9K57HyVE9lC3/GoQLqQ46ZDu+diU+n
/NzpcyXI7zkscMMFRdOre4AvDLmLChLLjDn0Iu3exrcoXNM2DaHXk5EJc9UVqgo2d17akDwbSEuU
EN0PoSWHMI4gRb0ZCyS7y+6B9eefsW9ToOr+b4SBgv3lEAHE6q6UFBt45/4uJU3LZvx7L3ZlEYu+
GHwjONEiFl28Mbl7PXCQ3QgK6ZDIjDtECPtbjNhcv+iajRp2S+xCQSmU0STlTGbrX+JOtsqGjjCK
MNMIjsna0mIsPm0SaZaMUrWHbBBX0JFizZk4rgbbGXpAAv0GI/ir1Xpl+pm096/NynOhIj3uSVm5
KEg2PHjr7q3lA4mBkQrOHKONH9E1l0OkI0ib1aO3MjVXEUBaupH3B6BoJ1Cl2AyIjYyMCHw3XkjN
5M9RZ8S/vrF4zgGLez4hMC03krwLVRwsPMsxmJIvOAaNiBdkNse2rzzFXZe/K3OUTwYhktg7AL6p
3bw6pE4K21hZpcjRRUPyDQm1sgRRRBNk0OkfiOG3XFUyVEU1N6dM9bkxI6oD8odUW9FFs7B0cgcn
dB052OIp0i/EwnTcRpSikMuBEGSn+YD7Rnnd/db1X5F1UfHnN4ljIQUXq0hnWdxTYPQOP9xsotzr
b1GxVboIcMvhXKapxpmRxJp3CvQm+5p4ZwwlzmhRd3Lrh+IOtNrpPnCI3E94VzxOafJzzKAul+n/
IwnfwTC49gjkL7ElPzvJLpJb33QHTt6fpNnwxqJxZAze7txbHVKMFa0MlQysgmla2f7cvslWN+Ck
qm02jDNQGB2by5JkSKmM5tX+d6z65KkHt7FhDx6INKHnQe/mnA9oII1IFn2crY8DWN7LWqt+6zMz
iRTl24l4wslqwvOgThDkXk/yh5OWBxTJdq9cYWCEn22AO5DqIUtHIwjI1ZysV5z3o7z5yZ3K3a3n
mkDisr92s6VKGxVC7hgO1107qXzENGtC1AH9QpJREH8R07HzTImAd7edXEM1V8+tP9nKKpjofVhl
ZG5Vz1flKP4POrsusGYNCmcev8JAXjoO7+DWTzjtKRHb2zCjqNiH1sudNfr8/ea0XvHIcjwV10/s
9JH3boTV3zNog+tUk7zND3ufBX1H7rkk4ENlDG2MVbDdrJikvdXzdGLs1gsaNQ76cOJtpJBow83T
pC+u+dlDg7iw+49fibuFk6EPeV+rFC5ynmQc07wb/CyazUKISO9jmK4WPAQYpENT4mFBdDiL/MiI
86AS2z1Ts++KB7R83B+I0jjJsUFEtrpbsC+OUll99y0WyJKC7JDy3BAEGj5a2c2u1mYiQppDqm4k
N8OlaX/Pi5VHHd4VYpennXwtGulSz/U/aENHxBvnXccd5+gIJyBIUA81LVkIK2fWueXN8mLQaDW0
OxkSvxLPaMm/+iA9LV9HTboqCtInjmSPHVGP2N1KfrSS+mr+0c4AbVJQ0cVzaU71kUauKLBiNSsd
DtkPdnNg4otuDX/SOn/Y0Ual2MQgcxC8xk5Mw+qb2nceRFQbPbX2TNckyrq0GqBLihFpaXqZKUgJ
aUR1E2WUdIXCToFD4Yrsz7RyBmmBtNR+/m3XCSniSiwATY0PzSyEJyYUHLBXdmmG/upmW7PSqyYN
UF5RBoQw1KH2DFWmYCAsfeyYIOv6+95UoCEf5dlZ+vwSGlciz6emr39EjGfwaK4dkp6kosqQ+ztz
OE0vxL+XP9e6+xk9Ljpa2x5QoieOi/NrSYJY+OPKu4ItcfE6zv2Jl0t7fnwH7kzcMJZIIm5Lhbq7
aboitWucRUZu/XCDx9YjKusNgkW9P+v4pdQuHZgQ+BYP/8dcrv08hVMkBWP5yFtB9oHGQeDZQEKr
U4gzOtP1tRP5Zf1AeRZHqM4kqr9D5I1N0G3oLMHwxlud004VxAjRlGMFIMnF1F+c84U2BiuyEQB6
V5CG974LNTDphIE6MkxfOvj+w7O850JcFe+JKfsjH9lkC4OSoJCV2+3rXYSo5ITnRBEgT9VYmETj
J4HB9zxFyDbOZGDANKEKkJD8p9gAFWAPLdJBvsMkmIM1THdRsqdz1HxPBrnz/U/GVYAf7clORM/0
sARvvlxyDYFuvk6fvrHDVLS1uzwtp1og/UjIVGzl4NB4ePCwvFO6vMlwdrRDwzjOiwBxUV2Yhntu
H2Kkk0ZAfa9fWG7sDHVGY1P1raql9mwB8yedy5RCGY2/w3ky/xTXVpntqQrRuwxw8+/f7q4ACEwB
ebCBBmFMDqJzzTOLzL2ahYYHn3RRwe0ccAFTkp6bAxrMxso4wtFnwH9y9VJSrEEK9D5g3HhWR329
SBwTROhWoULjcr99vBdLtVccBBOycopMaLztFpG6mqi5HRFu/x3oxyEev6tuYDZIKJnAnoFi6WY/
RtcFV4UGg9FJJB2Kqv2lclph+IIvthBl63+kY37gJC4VW5j594Xw85c9lhBLaRUe6oMltlDpAmMv
ALb+OdHCxc+BhD8H2KdyWUWhU+ZeBMFs2Nr/z2uH6Iq5y8OnIRDNm+0U6w09yoV/Y3StEK5GwEOj
HdXjwGI6sn+hCozMqjupM1QI0GrPiFeD4MHyzxkTw3WqDsKBa+wnzGCn/gkBi1HTjQIPNc2Qgoup
1tPYq5JJ8d0TH287tkOu+G3eKcqRGPLcWMh6jqvxKeACpN715mq4ce2C1aANuQx2blmH0bDBBVGZ
obAEjaZRpqHu8S/cQub+vPoBj1MH1jFBbFsT4TNQEWt96Ac+2iA+H9qieWTDt4VgOEozgT4BDlMt
EalAPLH+cRz/OWU2YttatOIpkh88HSKMNp6U2l1VbeOMyU3awDyDrfrljvk5rU7Auz6yH9VdxVvA
aq59+fZOrYmYOvzf0ROZYPAHd+5yTvFaGbmSjbdb4UJ7bcos/fJ+9ge8IocPjeVUyDMXG4vkcyS7
UrsXqknPzBczbppZhF6tw5EuGE189/b1sINpVjr6yapKkWDAt1AaipzZtLUEedWRWn2RgwUUd4ik
bYQE/1ECUwUsOZPtUNv+E2pnYatYkuTUnsAmUKvS1LcmDENEz4pQlfzSArrcNW+K8m4exdXqeM+z
m55SoWLAAcdSD1Fcc9bUNvAhpkn9LxTwqIDVLiD57ETjccjdSFt3QYSLTkDnIUFsA0VgdTGnCGt1
H8Yswm5ZfiXe1/UYNKQTAgWvIq8Eo4Pfht2wucaTDB9VThp/Nzl0vmgTLmN88zojKv7n9nuQZxc8
OEh84rXSbyxXmfjBgZWYDhYhSE0NtjAgIlFrjzATffzRZeSZ5AfDrG/ZCXN3s5Y/vde+LXJ3EZ9c
AedDtPs2d6H06QIamiF1vBvhnqyO1z2Wm4Hx8T57LJbIJpqueQJ4NQhDr/PCrHo/g5v42Ayq0rY1
VnXBK2drQx7MwD3oy+EYdQxw48I2JJF3RvrTQaapyY3FbSC5uIx9dWsD1EQVJ4D0Ygt3PwddwI7V
xxIqbaaJSHdDQY7j8R+MlPpx7Plrg6nqALJLilfbjPyz8cn8/n7NspreyUe6tkUmCK/+42K1o7ti
kkCBFQy9KmzFfitVtbjzkWvcK+2CRlvFXagMzLP+28wpFqnhnKXQozJvAK5thu1Mn7b5vxSFwgID
Xv0SM1dYYjRrPSUgrzyWjTkH++qRv03p7pa/NyfWtqTs4ndpoE/Okc+NzuyQ/CvOUTYKy0jfXQOn
8SGqLLMbcqTY8Ep+p1TTb0H1mupmPogK/r8lU+wi3V33PDdsoX09PNBB3e+xiZr6j0gpluDtOuhN
8SVFPQhx/Lh8pTxFx71AL6sTYD+iMWbPvYifFtipnxUSkmCVh1tBsJRKS+uYjRImD/5MOK2aXUkG
6EhL8R7vUfvO6eb8SV169rTsRGw1TGdX+ACxLxhegTtk3m2sJ708LyKTK0UzD0V0AePfQrljCyq7
T8/zJMY2VHiCRhZS5rlK+vaZj+eh4w0OotDXyxpy96NMNteuhsX35UzSGpZDv5HOrk+nBIgZA2C0
vT4oCVD0VTqkfd/Y0/M2z8OXEyu9fWunBW8gL0gulrHHHkcTKC5ElM+Wj1cOcX7GyLlOYGB922q/
g58r7BpIyFpdy6gDIZtfgO9KhJN6cUVhbCUFRXR1n9Z3K68KVuGJcmggUmkEsF+z910rSktJVrg8
feXZoqQyhxX/2/3FA9Fe49H7L3kNWtMHtCCUKhwJ1cn4t7wxOa4F4Xk5myTWgrAWUlDmm1yEHKNG
SK8ipj4UZ55a0vateUrlAFHVk92lJXrekqz1oRisk9LHzBBQ3memStwTZ1c7KfTRM6QjVyo2wHTA
atZELpYQj6NeNEdsBnF1asPkpy2Nm2Jyqc/8hgfAfj5IjCJdeWTSHgeu7qqxuhyZxjkGZ9gmGpyr
+r0t30jc1S6GixROiCiBxbailTgrhnIgQf0ijlood4wfrbQUwZM6nhc+LcDcMfhhWIV1DM6sffQO
yJr3Bwk72juptpmTP9UU60uuqsoXqHJhbcTdhjOnInVBzXHRGWbRXXAjXvK+Jmj/e9BNh3IIkrLN
XIeafYBWBkTAGYhiTtUh3BrcHc5FwgU8ooEBL5Y+AqW4o1cf6NdS4J0y4zwAC5JwsSUPgUpGaiym
5r1IM+xd8H09h0Ddtw5dKtfRmsC+ZxgFbKjlXM4k/fMmEzdjsRWthVdoCz47sko+fDxQ1KVNbbtA
/nlEmT+nt3oqSVmLDXgZdlidcfmEUSFfrdkio3gwF197bX2/JFmMARWagfHLpR/f60KmrFTxNTj6
jj4UPqK+XKH+lur+DGRS9iy8YSAyrRMe4wYshV4RWbu/IKMEfE09/gkUNtoJK8CCals7jqdh4A5v
IvFYPvaldrfVh+2tj0sclgaGs24BvUH1u+asAFXRDLVnryxc2Xm/tCoCiLMSwmP+QeMkq1d/rcd5
0LV8fgNFKkTrZhlMO6RR7pZ/sdpFwb3bpOFJ+uP2k+9AJicCUSIStD596nD96f9iHOgguUR4F2S6
KvemOXcIRboMDY88Dw38odXMyYcrIxekb3WbIgDEgUi7ICIK/t3A9oZH+EnKCUC9JjQkNw9gsFAr
hUpC9pihkI21rfR8XYaOnnWhPjhN11b+3uXzEK78N8dcaPJmoJIR04Mwv03uICQFlYDILTE+zBOw
UfPKg3phsr2q0tnItlUDMHNAfTJ6KzvZo+0qCoDCgtO5xTB7QX652/axGtEk8KQJZoOp6B0SV6kl
knEkJvIMZEHcq6l2qOnVX2vpowvXvPivkehhi9pbWyrXEnx7769CQ5QnWENB9MH4NDgOvMySSkCX
vaS87eHzN3IOGpt24Yo3dFN9qE/wkTbEX9VNgWU2er469wpf4pHbacXLgb2dkVaLLv+N9zozbBz8
DptrkefzlEMt7pSk5leeN5AKJzvSapXDUfMfvvTokbhqMDLE6F8uhyRNLEQ2R6lw0Yz+Ebx1p9fp
LYQZza1d2BRyxCUKThyAYgbNjfOgpKOG9X8/UYStza/354E9SDfWmHd7n/StvEENlv/naJdE8jOb
Nf0pbc2Inss1uEz2WlSO35MtLqDUOJAkE5V+B0/3xaqL+AbSHG2jLkWwizC2hcKxSewoS83I0GOs
cEXSBrJtyI1k3xMCeEO6nz0ar+40k8bL9gcClMt4rrDGCOA5/IaEgJyyVX1xuyjoacKV2+OZTAna
va74/PEtXqiF5BI559v9rubDCwLrVUSYB50BCrDAjXUa/1qV3ht+j/7YfQbz6Eu9jEWlTqLp28Dk
v7MNupKxMuwT09IJk/x956bAb6Jks4FcsiHfcPNyo47MNl/tQzrl7GVsxPAArmtU+QLitCcQsQvL
I+CPzRX4+O3m7XUoKv6NEbPp9BD01T3UY8LXdcW9dmZKMV/W0g46OHRFGQGumJ/eX3WGUc5euAZO
jWsHWATBuJtH7d8ItrfLe3S4eakitTCtSDlPKl3sjdI09HiALcsvVuQP/fb/BgOcdf1cUG0VeOQp
rqESKh74EMpfxWM9u0cikssYQ1LsokNrgMl4fu++AH8RvfkWPjZuFX4yGvKJS1/fta12e47/gdaO
7nBoimrOmqj+DSS08COTSHbbRIE7YhqTSTavjpBmhRGRgddbD28UYzjXKx4suSoA/AJJ1BuJrc/a
WvKeKhshFUtu3FFPTQIqywFfOKd8gd7k9CaH3YnYROy5H09VhNZu200LK4ZKf2S28asi+oPW+GIV
QvxYiPUhBrpxrawEueT8EGr6PAzlFTKiDUsYCN9ZrJxy4/cQAkXrhsjerviBeeT9eBrXqh1oBNjV
thZKaIbOOcKEWDd3VxoABmBD2zad9kj5N5ZQVsKArzsAcAhkgakiu1R+3Q7B5m5poqPpzOFeS/VT
xqwA0q0KVURTjULqyWu9kRzIn+EHohNHkPnZ5C2tL1JlyOymMV2H3pEqnU7cip/+NNyTbQ1LzNE4
ZNiwDN6QoPnqS0mCWDvOuYMYm6PfrZoh2lv6bBqXb8Snb6sA183HPPRaUeJvEraQWJK/O0hmdJMH
Z/U685edgiRLhoj6wWlvalMhmu3ufEc6uEEyXFI09pbpVigwkLMHvW1JNjdcVRRAkK7yEN9+TpqR
ce0SW5E+GM0oxKvZj5pqAglYBNl60y93dKuHXqC3NVVzjj93W7KJ3ExHP0JL5N9dlP3KqYplOCYV
jDl+GUzib+UBctio2f7fF9WfFRkuvYIuJbG3UT8dm7VMb+PwaF8laZhoXRiyueJaJ1CUn4AD26oz
xI8ScpAzhD+GQAji+4iQvlf81w5ydT2pFAZu1AEygfwS0S0GJIG5Y1bASxy2oAvywgL4B2kaiDGS
mSb/6zaK+QfG4VCiIstGqu9n/4viT+7lRCI673z5kGjmgegVcHbEjLLaURSmkYvS5ztl3xvQIs77
HNuU37VeMvq++1HKZJ98qNXeLAB3MKFUfZHi3MotWp+/SV5VLiA2IhE0xQPylDEUykTHjeOT35/s
MqQACHIeONXtBrz5PsYFZVWiByosa7rftIGtYQGgziIQAd2if7S5S74WSQNFviV5FOs2I2Eellnr
H1uIu/8JctIPXe8AHRcS3wFwEggdGZqp7yKKKX7UJpAyquMhCL0rbRA28kDfKgKYFQfVvJ3klzfq
8v1sCPMuvB32G5mbZg5Q5wnyNhYoOaJYPHTp6V7t4RT8WHmvhQ7WzQebrbnAvGREqwPFHZoimL7B
oJv5Qzl+cgAz1NXzTbGqnic5w6kltv1XcrRS0ppO0Gh5tzyWaoO4GPaE1hJAi24Cc6H71/XCjCl0
N+oy8Ti81iPfhEcwJJ2s6jh9u0OWme+GtZ5xPxZTKaDMMeXr85gVB0IXpYeQ7SnDDPbu9Mj+k1k9
4wi3zKstsUUTYgmehjBJdOdukEBxU42OuhxPRBnrF8xsuJfV3RnhtKGCS/0Tg4ib4t2o8eixeUtV
6pXgKw05Aegi8FdnQrgMsqX55rc15KC/zrjgzOiifqcYdBd54roddBdA0VCMS1vss7AAQc2qEYfx
dKxLaXo3S5rb0sGHy/aV5kqB/PA9XUp+Rl3mgF56xXcXMCTfzFb88z14J2WekBultJHJww570afg
9CY7R21Ab0KPDIhlgMJY9h3Q4Gnl456Of9dd4si33EOuLFAOTxJRSU+j8SQ08V2mU7Am0Tv6ItFH
RahtOKudEFcMFJKjdMKH2NPPz1Jm65GTn0Kk1rg1fXL3zbppGj3w1N03YxWdD0dCsYxpu6RI5Ion
llPMC0sE5tBpXIFXBqoad10u2y5OeHxvv1XfRmcohe5oVU34oUp0nNocDM1abYHXNS3LrBFt6+P6
SSL0Ku2MlAe5Du3KgA4jUVTP+KO8O+MGvZBIG+SJkxzIrDO1ruPvnVASXfxk+64kFFamZp3/rN5W
sGMa/gujTloL8kCym5Km0iiagodqEH/aYPKAKtRZZaM2RW2abbv9AKwbGcJfXdheSXNZrq3+ntqe
JW6x7ixWiECkpz8NegtUcll/piejqVcCX6kX+dXJYgj2OwsI87nE1K0j+k8fyJEGbCtp/T1f2crV
WYe5C+SVIIyIKaV5OIKmd/Es9jXLZUnYFtN3tL/k8VP1APG4fZG8kXZwjD+i5WOwJpT6KBfTPP/o
H4dXigrfJpLHGiD6kYfnQ/q1lpEp0PJKZtMKo8oJQT6vZk2krs2Ioaqsw/96hq5C7OU8rAyVDTI1
FOPIbQ4bq+/KaL6xblXA0zvsUuJ6xPzGvg1igdZSAC17bjvQgHZYSX1nafDs06JQqB/y6fU0ibKj
yRP8omeSvnhilQgDyq4xN/CJvrjPj50JpieX/O6GT5BacWsP1SRsMI++hTKwrkFFoefFBXc7Wjj0
MYVFu1l2hdPDS2YwGdUsjZ0A2Sim081dSmrAP93NZUMnFtKsX4EOLndNMKnH/YPKhzn5n6YUJD1P
LeSIFbLjh8/ckW3a7uYh0gS6FaKZ+U3ay5rbA1Gme1w8EAXFObtkMdYtYppDxDk4AvJ3A+qNa8kx
z9gozVxBvDkI0/dgq9yxvNqwHIZMrK7OTrfAArOGsYxR70CpbTDkOR1JCVrlSE9tWn5BGhLqyO7z
o+F7AEqrJZHpP7eLkCuCfDIqpZ9QWEFPi9uNKA9BzPYvNTRYlV0iJGb+FaE2EHCF0O1tmyxV5gJ0
89p6kGcJRaoy0qU6Dl8r6k9zprx+x8QlJuNiS/5gNXqIzJmS9svKZu2p50M5z+gKuzu5ozqUXKkt
cPI2T61EMoy7qymJw4uFyAPlNAo956opApGFU7x8Yd589VLW/KOIuS8DG+zs0XJyFDau/wE9JP2Y
fbMGpFupD0h+QeJ3xpPbb0kGd7YotaTeIl2A/KfV0b53zswv7AcO8VTR4sqKeXRMUsbtuNhXNsuF
x1dSmtCnelzPid+43HK+QivRlIBlFwCGFu1T/+1j7E9oFDADg/Rggy5zfZG2KLBrmGbjn/zAt/ui
TBxnS6MUcfjrX0X1xiA5FNP7aZDSTBcMvgQNE+owUgJkuiqtCjIKXV1rdcXruLjXHEm3gzNzbswD
k7OHFQtmRIUKvY82OYwirr7oNGyllpKAgS+JrYSjjfs2KScOHYpKR33YOyZUSFwxEK6MTWKt5t9M
AEcL13CgXgmELtkDILFFnlDcEomQuxnvF9zTgpsVbb7YRVD7B6UbSY8rpwijnoSiDkXNdCw62Qhf
RAFFaZXGLI79jSwGbp/x/GLVIIZQ4Tt4fO9+ynj1bxMWWDoKBgFGPzZi8J0Dib8dydATG+tuu5n+
2vkKTEpGlqGGtD198TT84k8PQ6gz15L+3hIfyrTDizWXxL/qmHZxsRkz7DvHoxxhvIpHxPuIgDFr
vtkZZ9vxXhnG8k9G/uZfYfeTwSH+9RycBXDmDfE0CaIIna7lieTMu7QhATfbBXvoQiBc2UsmVGK6
7QkfXLBLtswX3vDaL8hLCm1JlkqnzzMGOO5c5yHMFa9bwqYSCeX06XQZp8MvMSWdMDl25A4cC7M8
Tv+h8hepPsmTYHpcNCvHICjxCHQw7iml3JXJUglKnKjLYEi0wxP2EfGJ93DzOCihl1C6/AF12tCJ
b5ewoWfXGdxnMkuvF0tQqjXXYKCMgt405bvEGAM3WIstUPAV2Vda3o5azjwxdJA0ZgP1crM+Gjov
RgHEbonmljxo+zjxn/eArGxV5+RVTDdnGhiyUd3HC8iihwzmpZH5KLZ9p0/W343iPBak+3KYLOdx
PYl5ykpe+mbvkl7xU06O0X8eKEn8Yff03rGjRHWbtdEoKMTnIDQcPIHCkp6eNRT0bxdWebWy2A71
dFK9cMPFAHZ4iLj62u8hthshMUHVpWbzx1++GL+SGxvhnQjfWIAlfikPAiqtE9KlMSj+4t0TqbAa
HV+OuBbPdHRWOiCkOjBNpnQeFXDRt62XHy+wJDV+nZJjdhE4W+Qwg2LFj0k2sQy9+WM6+3uxfXiA
tRZvFL9xekwET+H6G4HNW79yf1oFc2lHVxWD2yqTbV/fByh5ASIotZ+0oJU4pPhuH1oAeg9A2bF/
Z3gqC4Xgv9GC2Re/W0scscuFIlxIbPQc45KqrD8BieJ8f3I2fykwg58HSlA2Mwm0xbBi0/5aySpD
1MemGdH+Ia4ZxvshVS1ltMEzbxnMMDnybFRdpo9XTN1eSiQDiy7YjAJdknJ9zi98nqmVY9Do+h+H
HE6RgXPkR/yAE9/w4QOdyVzq9RtcK6sF7954UpXBXxIrHEHfm0jDE5CYtdJDnhMNFUkSaxI7JGWg
+vI0ir77c2SA6rh82tlW+s7YFzVr4JLrxnbqB6L4OHdAgrlcCf/1c87/mEszHEP2XRwu/N7EY7d6
3+WW2AhGKAFbWgqQeHVqJkWpT2krEw5sBZ3NKXjHuC+FBGgY6zYmqR01jHMiQdnknPrL1cLy7fq3
i0ME3eMgCwBRBQkO11Re/KSwbqpIm+3Y2qPe7gpfvfw08mARQ+xA5KNS3gqg20SdZTQVYOex6R/u
vD1J84lHpjAjjMGlTEkILjs2LCa2Fg/malT4BtuZrU52eyzvC0I0/t1uzemcFLzZOzEMY8UMQDMj
Q6aM2BHrNm8NEaZ3JNMX2hK+8HrIDJp/EOlwePQaxtXknaQTkt0eyeUmsxzLMk1ncezV+WsinDlJ
Neqh+yvYw1DKFniuJshh5371lPB9BV6xF7AUWvYkYS5B1Hy0Oh6qEEC0dzq56nHFpftjtmLztFna
Jmuk1UbdtwIg/Y6BYzA/vQHa8ke4SPiVX5/N/VKnklO7WMbvyFP9RTmoLWpw+O74s4B1W3Hi7Gdw
nVM8Kqoimses8e00Js2qm1JsngQZEzCzeUvWuazgYbx2rYnFOCSZ7+opl51hjqyXqC52knjf/S4Q
cvAT2/7FLXRNqFuFks6U2aGv/SqeRSuglkett8iV20UrVhkcvvhHh+KnHv6j6zoJXj9VkRw4ykKB
U0nhyVL7+Zj4GjGekSYr4y+E48otdAiY8YQCjYTxDLozBtTcyEdtIOXFBRPmIIE/+ktjl5Em5auf
J5ODiB0wZf2UXSzIzbn8lOmKGYTmkxyEMxpZD4mv5nW377Ib5RmNBDgIDRTvhyZva53zOQjjUO39
BapOjyloszSfzaEwzLD2ooblAsnCtKGDOV8TxHcZ5OCuXO+VqE9vpdRgS/2IHt52icnFGSU+AMk2
P7lW/YTFxbMRTyYaPghos2OHDanIAh93hy36mXDQzVT7eEzApqM6O8EJn2L7mkMwZuefpxyycWL9
AKb7UnVgGjWs5oBeAMdjzonc8XPgUUSe+u2RZMJLqNvT1LW9Tr+JEOWflcEclL/r/yoY0pagzXs3
UFl3BAK3kmN+rDvX4AHbBVW1WqxXY8JHIAJEir4fIMlf5xuSVf1uuIrUH/N6cPQ8x/wGpV2yAZKm
yB9PvzCiVy+YDjv70sWq+kWQfc6qeeyYDTDOtr9L/Wj6MCvwWDfwKMoh7t+w2tIOGiiwYEMI51Xa
wWdxcTMA8I1f/0KuyXNOLSau9s/1KsAK4mnR1Ip6m7mwn8HAe0NewP55gIoVKsKpfLdoaK30/3Dl
bQieBQr2Syqaq6picQ3guI9gnaMMDtm032DglZS4ai2FGoBCWWLI+3h+fz5z2crWMCAh4Bug7U+f
vJmJ8e+VUWQV4T7hUP6SNGR8lRM6Y1wxvfjjiCxPvW+JNn6Yx5vNxJTmYj1BUt+OJSAGHrlzTkfX
q7sdortiWPcMU6QRyI/A6ZtqzgvZ+n4/0tt1pVeKH25qBTDetf5R1B5lApvUO8+yh6zHEKndCmSB
dyUHKn1crUQ62gOgbDxBG5rBDId+ban3+X8R5ptgqa9S4mYTk5f/Aqu2owoHMfp7cgogh5q6Aw9i
9ydZfKAle1SSJAx6Gz7g2wiAlElkdFvFtjl+jKncrPSpMpW4ZMDQORfKCfTDFC82tcjdyKylREcO
1kSmbFS8rMQadjmwuHovKQRSrfYAmfgMb6ibmv3ybpXFSnyUxDNhyV8S0lda6CEQIcTVs187A7vz
0EiMkc3AA2nrqRcHynIa5TyVHJK2rG7FV8uNz/JEh+EQPzHy0xju5l0nvqb14VjdTCNW9N6raAz0
cjAujUtD+KKBEpudd49Y12xWWKB79pb5E85sJaXbDxvB0ZwVGn1P9fU5QJklJp2nZ4g6dW+Rsi+T
mTrjQkFFeDaZ2GGV0Q4mzGKEHHjZAU6/gTaIEdF6TY0nCIEmu4FeFyMSoC2xHXGUY85WdAomzxkO
OhciVN328P1MQiRclWOPYyD7oP5DnOrj75AQL4hs6itxDOdF3BMbUgwB+CI1zTj7lU91PESTMSau
JnuDxPcSsYBHaDOG0LmN0qv0y2nHxRoST+6w/HRcAhdIjhyWtJ+bnbjYmTe3KTYv5pDcqAb92g08
kV2peGpakDhaAgoF4zFQVPVi0BHkL2JfVIbNjEZ4dbZZDZCVoDGEeP5QkBomeFcfZEHRMKnSDfJ9
xpRNcjpcYRUJnZK8GUq9PYWN5t+UKb3AB0kYjQ6sPSaCwn5ztPRQ8Jdd0TFnzKtzhrehmeXJ3c9P
HTNWxEvouEuNAFmKJPqeHRq2Qu5Dt+u/KBy9XrS6doxa2HG4ZH3i2wrACrihlaPy8T8jU8cbLf8H
NY8TtNX6wL+zigUV8ZbfKo5BoqpKmI5YDxZJMUqZ9Nk1GmXBzUWPt7XbHxMxFD3+RrQoe+5nrtZk
+0Iuxy3LMTuN0oQvFOdK4fqdwj0BfQs3AHp4/rCEWM7AGc7UFRDuS+OWhoA/+l4XJra/hU4Db1bb
e86XX5AGr8QHx7SbKExegI8DJ1xVHN7SI/Chb1GidtgyWIF18y3vqytONFumcGccDul2b9/JjN85
IVU0cTpM0ONzSuNGU6Iqy5VteYmRfLGWwfS6i2/14OxJz9DNodS1CfpW6B5EA8fsHAy+EY2awSnA
/J0lDCu+XFrXtUrSLXmjDGl7xAehc3ZUh3O88uY8EBlmfwnSzq83CBkwhOZb6MpqyK5rTlZWrGg5
ae8fiSSJJNw/biyFWqds56WDlu/o0PkRCyO0hUDQGnz/txOsbyCFzETX3fYMAK5myCEkmZejqjC5
l0RUXqVo4rdqJRdvxLc4b47xopnOB+boWCu4wmbCgXhN5qqHUMPYZYsvVUV+CooQbutPob7ABvH4
lQDM4p62dvD2Hb2WNH6Zv2HS/ZCJ2kdFb8vtnk4K9h7qhfnQPc6DZSAtqbiPgeUCDu7qY3y3lFgZ
XKJZd6BeXIgTfnjYWHs0wDvV6nyxZOfV/LL6ic704EwnbIS4RVDNQgfYZiYJ1vNum1NMTaQ5C+VT
ImsoqYExM1a0DVhLLM0E0zr04kVCGjCsJ3js4hnEd3extbMSlQvBJ18M23dSWIhT/1tHw1bDPTqi
4OZi0+oeyUyhKwAbmjjEu7sJJpWtTF3gNWpzKn4hGV1vNLek12MDqBEw8DL52utSGyI4aDnUK/d2
F8P7cmvv8Rylid0Ncg0fd+XG86Y41P9FJAIXf22HQlvS0zmY8Rs//1IWvDmnWS9vik7cX8bki8h8
uWIOxx58RPk1VID6ATUbd7a+UyGs3EvE+bJCt+KHHVVu3bm3lupdPRzcaqowdT/Gv0s+GUq6rffR
Pk4VkhQB42ZsVjsyWCZkum8N2SGbyTy34Ud4Dr2x/8xn98Ca+xcvy/1+enN/DvXfFHP5t5eDA199
F6Uxp7f83QPNPgLl8U8o6irBDNeXBmeLXO0S7drceKUkCe2evY5yOWR2sIV/K3Z5abew4NE6GH5r
Ibtd5nCb+DAh7QAU+ViRGik7caKBpyOkmDjOGGb8M88W3zoE+E7r/C5F+JjolM++nqTHcGRfBGau
0QDY34YpkpVD9lsDImmll8X20nxayR4vW9frTKtD7T7evpEMHeT6vZ2XuHvy9DUcBdgjZ08+wXK1
s41kRjJfCXeP3vqzL7CndLZ5hhd3OZpVNzMb2OzrJaRGmheZ/wTGq+14wiwUYAih5kYGCSDgTmkV
5rQRCx0X92ifXMNoOHa+jb/589FaDa16omKAYKv5vhZPWPUdKVAeN+zYKHfYXwwh+0/W9/pf2Bpi
wakHGbDlNmWz3FZJ31W25/VAPvbxw82jbHlFq1wi4XQgMH3EI8opCSPlBOK9+T0VxqAbpMYtmWtg
U3AM0AM0i4CIu5pkouWhe0YaWxppJeaoLFio1/2k4dRtOKlITs/2zGQwyWwYWXhRc1VmDpdds1R+
digl3lPErAPEQLVO+wVN2fmN1Z2ZEZsxL2vvn5lTBsYto4iuxM5c3V0NuEfCZcNM+KI2L9Wyg6Lp
xJMaEMIZ11TW3p9ORX0SeWYrmuBH24Kfkb+VLGdPGoYQzf0N1fIE0vB7rUuKZvQN9BLyEXxlgW4H
qJc3a3EVKOHkmtu92S8AZyuEt6AzfW9cbLYEkS4fnbgH5dnY7s1G6l85aPtwALoWd+jpcYoXYden
Ve0Qo/ZaqtiqEP36GN9a+euM4YbLF57M9Y7vRkwR19EE4iuk2TCsD04Mj2N108Q/9D1y9JS5ZGLJ
8hxXrS55g+oQ6uSJOBCRN0lojZMLvNCerkIJAJH9BgDY8PRJKT1aMwu2whU0bV215sbrTrDpISwu
tfxfUFxgIwrOFogw0cLFfvMGuBmRSP6llYbyWVuH9bkPoH24bqbwFKvDdij7ibcT3nRXkqSHz0nx
jKvFWFb7mCf2Rb9xTgFPbS2lO3aswgOX9T3GmXGQCHv5CLgfB91DM1OlDOFE9OcEInh3okXInYlr
kfKALqlbKuoXIoR+auJWMC61ZjGNPBaONLZvENOeppN0nqWAzMgxFyY0sQefr7+cLm6AWKui1scA
D1MOF7nZUmKgZFZkmG5vFkwjomTuI3ajVeMnlYy8hg6iOruVMw25Ml442Ban3/LsnmhN76GuGKoi
lIa8JWwpd+fYJHPaK87Jfz0gAtDMyf76MCLtbZ3vsaN5wrUHQnhUogwqLj32H6/lDNT58EWkc+Jq
EG7/ODSnmHwLgkXxzoZRgExjL2RSOzQioVlllW2wESIch/lGkEE/1StwPCZM8P5wh52rh54y5BkD
VyUnxcIJ3KujF7t2tLgSGZkLWuVXQnQa8cByZ1HRT9zgA5+H5waSoBe7AAoID6xOusJptSyZ1EY2
NiNc5zehd/20i0aRd/MFwgMcrCgkYpQ8debbn/9zdnyiLsSwtNxRAFcKh8Ef0rsR98sVE1tn3ukS
fPMO4tXHRsiRXw5iJze7KPE/brMQy0rQV6ix9I0XlHuRKhRiMxtLYH+8P96qC9mjU0eDGggTSRKu
aocGacnGYfzHAAMAsMy8XSlkSFCpqYyJw6huFKEG3mlpkmwWwjxfHAo8exGcu9Z0TmbCe0QJovyw
LZ6+sacV/CT/xJjnNdaWCaSn+dehisZwWLOKxdgeJzwtgjcacyPr6DSAZBUIVgHVOD/RDydPoRrl
Z75vnJEQ4hK/KVYI+fK3axn0fBFuaT3DXz+UMNEvD+51SQ8VZq9gP3ZOilTly8PaJ4KUg9dpjH6t
GQkUGZUUZjd+Wi4xZ32AFluoyaQEZEp+utY5n9C2Nr0dQg9mrELvV6oReZ7z8o93Vf/mWvAwhnza
yf0E+o0XZ1c+rGP9U376mgLJDE65I4ILntxRoIdMbZnDDe2Vn2h1fkCuXVWNT2YQqbNfPMAnZ8JR
E07SEOfINtiW3+J1UveuF5pyIhbmqa3XQY24poY1+byBCi2+xMJV01gVwUOtB0XtxtLSkWMK3u6o
3YipESChOcLRRuSzh7L9J+I9bzeW6yQpq/+sifo8h73zl4AD1FbAEE9fvtnhlnvFdWZvwAGZKgSn
QHgqiwHa4k+rQyFVXRUXT8ChFWvfZ1E0y9Ujl+omLZ3sKbbuo9cH2ka8iI8dVbn/xjjehmcfLwxE
mRGfjxYdRREIVkDH5CQQqW0GzEQlWNLUcsKfByatIN+R5ZoYaOY60kgOXRCa99WsHY3H0cslB3zH
LtuCe658YWCtU9w/b9aTW6z6JZmtot8Gs+sDBer+aXkeYodSnrcBHIoXHfqP6HZG5PL0/xGpdQYI
FelMWotP0Dks8xEJg5xb0G9EPDAbHKqrMsIqIj56H/37aJjX9hRJ+RmBArRMV8yy0msbSVRmaCoz
JTcN7u/WMNHxxS2oQTC5Nq43ksYXrJfBOSvDZlKMywwshWfuLH6T/Vqj0OtWEBHFZQFWdWptl9sp
swB8TkylsVl2cngkA45ZsjcuQwX1Ba23Z6iM1I/h/ExBH0nJ+Vfy69SYcM6nN+3Xfbwk2lwMGvFU
t3iqTKzPZoMDHMDFp1V0QoJ+ek8rKO5LJKKpJKL4EkCSlHKyRYbl8/V2+DVg1gN9QSakCHMHs7GU
aEpbr39MWHbWSaifKtt5rfcUucBF5ZYTyLkVj+HR0cYQtgsKOcE2JN+tBiOjp5tDpmlTRwrFcTc/
29Nz4bj8XI1oXLx8r4v10kc/wYw2Y9fZ0L+i4owTh4ACpONy+6R85NLxyMVVKkeCugoabRGdzxz6
CePJ8cTomjkZRX9CxBjha96eOmBddUOwUwO1nSGHaT/m+TjSpZtEZcvj4IwQlfOTCODhqpz9IxWa
QgU4A9sSQ4uXHzJO+4D4DBfxv/+6KIYAzr6S8X1BxqPOqzlOJmXX1NZe+zULIFbWrxidCAOKfChs
yDQc9b+PTEgNuKMEmkEYibx2jTFRTPx8svd+N2fYVQ6Hk0lDLHOS6BRsxwCoPA+z2LH1qAF68H3T
zawDihLuHObkSjb+CZ09RDovHRS2uFW9uvjKbg1VGoWmZYRuWJtoWbTlNqrTupQvuaOo27T8/kfD
gP+MNKysw1vrNUZaE8Rs4N59hJsc8Ko2yeoojT901l2U2iIn1IJ5xNvGsxnBkYrdll4rTaew0GsB
hjsanXrtG5DXWQQ7kkNVDxWOoO3xvHUAfvTdtHOFKpvl9H1rPYnOSVCDyy11+Rp9cGN7NsBT6kHP
LzMtlPGo+x+A/0UUN7LaZJhk8sWBylnCo+6XQLw+4yZP2mzRD4nl29TPNZy3j5lIHP5bm1/Va1To
Pqa6CVcAo9cvbR5OKzORPQl54qLvugKsRCYOEABktZ7mpv1F7II2k0FLStrZNmLGWZ25E0za8zpR
+gOSV6TOPy+HjjcRCO5/Z9EELySz998tfKhxEad+iVG+3LoRGxOPhmpmMzIRd20wY5YM7Z1LC8hy
UUXMyaFDN8p9hZccsLZqaHgBVAHUKgTutojtIbAG+1jkNh4jB6mKTik+/UidVmgSgu1BsBhhossL
OxBzNNva4Vgcsg4s7rITCH4R3iHJSA4th0WrMtEuNUpUMQzujGbuXcrd1rkH1SifEMWfIudjabdE
tzw571U+VFrkVuFa2MCLwmeVS0Jw1JlzxoRW68p0YSnjgzyt+TDFZ5SK3GCkKEAAAHLKUbKdNaqL
8KEiIk8WfvfnEC3Qgdk1ACZlKq0vHkc4f8T4GIAm0f43/uYP97lWlV9zzZr8sG5PAY4qNbCo/cYA
mv2AVT3L74r/zZDF0XWy3sF7AV6usAnomwTAHo+5jVP1BXrcpcxkEZK+3twvGpprFAyh5Vhd0mlM
4OQLvJ3d7r7BygSwySeMsSZIl6jzDsk2pObUdtI1fdZ2TseS6Fwvt/Uk8PFrwp1ovI0IXeMDmf9X
Ey5cwKKTYA4SSQ4+C0ynEa2pgEyrg6aU5b4IOPveDWwvQhihy4EEmCRcCUAqpmR87850z39Mx5pJ
NbahKKfab6mXAJbi+v3CdAW1UPkMeoDkczzobLnetW84zdab2pINySa3ooYLNNj3wEZH05Q20hqi
S/pVIdfxsMk3qxDI7DV3F1IZ+YZkVbfN2wvSBWgDOpo8Zb8UmL/4h3Db9RkKFOot012sLSnjN2Fx
PpZTMnfUB4rWCQEs5V1WDdBN5aP4sPXUZJWFI+lUI+jTSqPjzTiK/UylW4jHYmIoscseGLpZZl6v
FnE7RWuABWFt6hclQ2h1UJ6ULzR6gJbPtE34pmdMHtFQ4+9vFxuXS1ojYlwKdd3qy8JMbb44Xxx3
1uZtNvBaRun8Di3Vt/j5HsRYBP1aiJI5RECnKIb1UjlhFzhDMlOHiErMQidk8qAEGhXnZrXQaLxS
SdMjYFzXmr42QlIio85j7aNuynjdw0+y7GVv5VT/tl0VNYtrO73i7fCqJiKhQ1l1vyh+q+ieHFQf
1Lx6sQ1vWFk0/OzktOdg4sej6h8FZ6poLGUkYhiftu0lizMvpz2jOorooUKFcmwlOwE/VREVWme8
hM0v6vm2+gTZ8uk8AghwkV1gs5lGqVlRwf9evTTmZ3SyQXQtz0FTdIJ2N4XpzZg2b9WoNnaktXZG
hejIJEEGQOxDPpcEas9tQUupPPjYPqDWjUyPT3I2/mTQwNI/a/lSA7Z3b79B3CGN8Mjq9igNdqdH
+c4byj1Kyot8pGhyHu6sKJyCrJVX9G9RpACT5hWt1iktz0sq1bMdsQe6zO1vTztoIsE83nGtWpMF
rrmbx/wSX/0yjmJLhuKyygxzlkQgIwF5qSKn9OxlMZZx7GFSO3dGZl1eshCu+b7a9RVnLRXsV9Le
GiHP8AjcPys9fb/ebUwutuzv89D26JQ9iSkNFax9sBovYUDcA2u3CxQuhXLJNw07wj1Vx5BpCfML
zuEFo6RSVoYxC3QfO0NYpzO/H8S4VqMPswliqIjmdFNSEGDf/UDCPEh83wkg6R5TdQ5o+GAndUIN
78ggH36Q8eUxiBtVxMCIzauOGRgcWgMDzXTH8VtmWnn9NsjOefnjnEhWad+ncaDCFj9+5/nR1w7M
RQDCSzbNryZjTAHlSV9V8/ZQASc6/DBAcgs67aed7Hx/Lp1O/WDUZMhRcVKn2u09iP2dWS+KGuXI
WrhdwAsQEk447Fc35GJiXakrE6/oaw4ApV+4oXqO+Iv+dNzMNtwifr7Q6B8FIWgRoBmz9O5WjUP+
Ve0UjnL4BdALVgfFZ5YRsccaq13FBhhq6ZeoXnt6V0gNs9aZlMwaqI9NfQR6H+MKBdBEvNaveLPQ
8/nx2f1AjA2xPN97clc39jqed98Isi+Xg8ZJ3VGKr6qAFULHT4qRhMsWXDVMAaA728zaHRdF0K4Z
rnlhsWiX67zeRTL+GrXNOh9E4drAPBX6gyPX42vp2ScEQdLQOnicVa9uei14zZFA/8usplfUL6m8
a37IAnNowsBivP9RP+O2qebaQWBl7If+3A2Gpw1pQkYmWTRe7+8iIWwMQp9ctZlC3lB1jX1ps0ko
Y2NX6QJuyWvWiFc0zon9Z4TKgtplY8Jg75TfQZfC+cc0ZR/STos0I2MCUWwv3pXuVwSecIuWNHCb
tyaZSjYQqOgK5xRAey5iHoyIKRcd/KObYOzLHYfPQbm2qKkb7cZD2kMPjMn7cBkPRzYjVWeaNNJC
GLa12l2MG7mG2S9dhETsdLEC2YaSgdvTpEs+rmIaAaFs5AL0UyLAQi5WXW79G7GzJM/4/McUZhYU
eSLWCt397tsoI9RAeITDodPA4cqDU8/7EBW46DYIUAJIayeWNWkw2XVzEm3b4FwwFxVO2Lxhoo/4
tWA4dofdYez0hnhk0qms+m8O9Su9u5Fbs6wNFbkZOe9obrGz88OZ2iSgAUc0Qi0jfLV0bWOVdGnZ
vCIg73W+pw9QUGzEgzHvqpqL3IspgobZDMmbXpBngt6mxUQTiEuGkqPnESXUl9uIngwPwn6diwHw
NnbLjQSyir9XKRX2mTaY84gV80EPPgMF2rEy7QCBWjNGXFrbhOfEx7/32bzIm/4BlGRQwtaXid6l
RXjxkhXzP29My+xv+nEF0r4w8U+tekxDSjJ6MOALq4g1Kqq+XyD2HZwMsWZhl/F7VONKAFU7MbsR
0YwTacqrNOT70MnvBXXC/ZVkiuWektwKjtf1wdPIcD4kqYfp/AAFbSuXoAbw8/gNdXklkJTCbJ94
HWeqljtalSoL44eH/3o6kGo5Sj0QUuV3AKM2/r8fR0N5x+t6WRXlS3l5/ykN4p360kHGssBG0dXG
MpTnhaNc51OVA3QKf467i+ZlRWeNboobI6ImWDP7199wZnjWV2PcDYpmKA/lwFKjNCkhx2GpGKBj
yfYy4qUYQRh7NPFMlAkxazmxnUGptxt1npI/A6jqCBWhvX18KEMI7NET5eJcauEqLFFd+zWFzpwS
smT0T93G8Iz2QvpAQygk7X6hedTWKPfxTrrJzUlI62lkp0v9PlMEbPbekkxvlcROiSmYMIo+cXbP
BVeB1B1lCL+8vGEI1pjY9mh0NOdRoGQXtR9EKmNT5p/exmW2jYKmgA2ZY4WM6H03stpJb290sAUM
fU4N1vUh8gBRCemlvvI+EeRAPW1jE41WUhU8Zu9seIQkTrF1eHuntMnFplYz1l80E7j1MBvPezUw
N0P4NDJ3pxV0EIN/QBFTJyzeXOoro8iEbUQZUszSAo2YaWAUnkatXBHqY0AR0KWaZ8h/7JESTiq7
A1rwHB3ohWmazKkhURrREcape6fGododCpt5WqjhM3bF0lbel65EAGa6kHyTB4FkUy2Xw7J0XSCq
c13qYYeTC1lc6TCXU6rNW+Y3dgXACLhOvIEV1hAgAnEDIPEWBUyNm1I/wzYNPbzA2uf/D4+J1VL3
/7nmmnsi1QQmDiWQQY9IaEandDfb5XZbtf7txJCMJHxA6ssU1a3voEJLOvIaT8Bdo0QqVywNKoZX
zsBmtjchG5uUhSCowYA1ALkBoJAl+dQd+BWfW4QXK0LAMHMt/K6Jv15GNZvOVUI2EQluf+o/XWKN
/kF4/oi4+t8qP7/axvr/smRIbbpqwPHY3TyrdCOEKgCHv8XiBwTTZKLvtHJh59YtYYl5meSugpdE
OJpp5YbW/I/voCHhIi07dINRGl6sseiSALK2j+6qF9f+Z/kHeWPABtMhpe7Rt11PhwtPq90a27lP
JpSBYrM00Ff8q47iEU/bAAe7bfEugW+pmAjLghXmFo/4h/8QiHEiANJDa2B2/e1oV9ycARF+vTot
H3LZe8QEyHYtSXVH+GCPvHEGO8ux8Ro/deu04Wf5oTh12Jw9EFtsADHsnTACH7eb8IBszzlutUZ/
M85nGaq9gp4r56b+9Tmlq2FOGZdVa5eR4e+6+6VWC4qkCATXSnUcy4rmT6pgu9z1/DixxbBNcUOu
H4yZAjY+9y03mPARwc0+Un7AXSqGL8A91ZqPlu2bhzXhWO7oyluAYZCcvjDboCMXk54TAwzFJl+Z
bo03OysofOI1p4/lK2VQtN1f+C/B48Hy14wc8BZXvVP7GSKmAJA4pOZBnFWu+Yg/58KIuiRN8px8
IeoTuVVZHBQY4h7+h1+qggomeUSNIUPLU3UQZ0K6uUZ14KRrsLjI809kdV8LvLmF0ta6iaKZP1Eh
QWdJVNGKcJ0kH5cPbT5mRLIAoAeIvM+Sv6D4YBlqVk+9Sldy6d4L/o2ipqmuQ3PEcXMdnrS+RBvy
xD1jcfHLc1+EO9uAKE28UtLrdE7PC8ktRL7Gi3VQ4YRCD1u9uuTIhnzFQLByexKSmsmJydiKFEMN
nmEDp3R2ezU4YbbUBJiBUcxL9t3ObJ5KgEZeTYFMEc3RaU+4QAq5McheB+KM8zrW7Dl99pgcWbUf
VLSdLAG0BFdIgNXncFQJygeNh9QZlJCuvI66sxgYMKPpNe72yPcySrMQn90AVNzC58hxDQ/NmnAA
QjO7cfySNN8bMtRyH+/ZjGPdsX1sWYBZSJ84Cpk+kKtIHzAEZQ3GSKprdfiKQHlLDgLP0VD+EPc+
CKFn+ASa9kf01vUKVB+W+HTpt4qIwIvw/R0415s1+HkHM99XbI7px88mmSi+W4Fv6gqoX1yeKosU
bgKsFkx1GTwS1qgO1HQ5v0yfqypYF/ORlkqufyP+47Ma6+PVi+Nd2Pqjp+z2xdOrEiLx34icj6DW
fjW0VCfnYunDILEiKh5XstJxJ2fWWcoOyDvHDWkDgum+Iiiry4Y9O28laNl9peCrxHaYTiP/l0nn
mxK4ccEEQvxlPoMP7PbQlkiUk8468FfIARvEGeErzDrSaakDFaPeHcchS0wR4rT0BFBYVbGJvy/J
GtCGbngHmP7ZIWIcuzRKzHwSoCaXHKzc6b+eJpgOkJ1wwii9WI5fKIMbNL9nYyosTElxc+6GbHRU
/EhJjPyMP3KAC5UJHUyNQd3DU5V06BfesD1lkHvrp+d+5nu+GEB1CSFGHrWt0LWvxRfU2aBSWFIT
Sc8OS9mQvkx61yXKgjuK1483KSJBlV7l3XugfYqWe4nUOs8TLHRiZNV3gIYB/f4fxza23z04Fr9k
4QHS3qkAs8G46TTwZoLTWVtGkrUCEHqj98wLXDxXeHKOEe/NQyltgWPqOwiS4WR39wtIaSE5jSYX
ljNjOtggCCHhqS/O9DOqvPcwVLllALuDXSO1SxakXL7naNTFHzkaWaR5nWxU03LiTCoaCAOj8hS2
xRiwgk+f7M3rHO4QcO9BPUQe3rISirswMgSMB1Nf8Vb+W0pIjT5mQvRPBxJAJzVbmvH8n/Gi+IU6
toCi3WMBk1Mgq64DEQl5LGLYvly3R0TIcVxisi9uJI2Z3u+ecLeWQ3Ky8K7zRnVNsTtmkoIfI1Eh
nl0LAKhgSV57ktpnSrnfzWJwJsPRcxYM71H4z+xB1/YuoK+kA/yWGwOGRnxCpD8l7sd/TYiCF1qP
gwWY6cqLYnniwEp5mjcdhd4L1VqSC7zOr15lQeGXJwWLyZq0QScUTMaP0tsixyxye2psS9adpdCl
0+DEmAWm7T9Y8noONmszse1lep7y7AGHKSf2OhCd/DLUl1QbswXsgi63GUSthm8GGR8w2HzedSS3
JAKGx/2U0h4dlHum/eB03Ximm0aZJ3FUGI/EgAAkE1IRcOgXZG1RFv1u2d7ettg6ndFLhy2nHYD3
eiXaesSECGOhfyzr9AU0w2fmd9GPSNyoikc2mI6E9LHLBtTsvUPY/WBFjNoAgIkRayNxzH0t8Fev
D+nrsSWVKf2D0OPwe2/XrkbgrMjbCGUcRx5TFYd/BIaR44g0wuQsLScKs/VG6iS7xNHYSqVGxv9t
Az90p+r4+IQBxTDeEO1dOCNOdGaxThsYduts0kuIhKLETKvv//FgZjkbjip7lWROua15q8CQgIXx
RIci1LCF/bQIKenf4d3WXhkoZb6avxgtqb9odi2LGk5HqorXrcUsbbnUsMcvBfhz5zywVmrvvbEv
7f7ziYfADvSsDVOo21mc2f+Ryhd8NeK9/8EQ5oM7Hj4MUyGfL3VWnynF+Fh3JoHf/rK9wbdo4Dja
hy1t64t+vAIrz+9GVW8Y1Aqo7p6r0VE+QVIZAKnsnmMdSuX42Mul9kVuwxaF1ZZgGV2oLpPJk6aY
64kK1ojGxXmZaTapivFpa6dg/Bz5eKvCNT0DeZxUa5Qz6KUyDHMWdS00wCvUCdLVw1mkSlniO1HG
2Qtr/AavlC/lbe5e5YxbhIBjgNB6RkuWeytmRJrkQPgxHcRW8VEknRfEEfYVMpQkMjr+UKWHeyB2
YPG7/NpVXN1stJHFaEnlSx9mUlZ5cqzOdO0K5WCqbT9opUldCPvf1bMhBoLYBRv7kHFOt320jSF7
Jz5kf6OErBp+aqvjds2ETQS3+FOjAW30rpRPLIz2JOZovGKvXZupLNFvCNtebBjHY86QaAdmMVps
mnTx/U4FTYRinaHTwwJ7czNnRoF81ltw7q3sw/b923jqyOR7ZLqWqZOPtypLDR5O0Ig8stmjPIfN
louw2yS6U9orBol3bio5pAHwzSf4ofL/WsL7V8nps/zVsGbk9fGWUK/QWG/GZ2ZMcFvTcg7gmFLb
/7Lr8IUXH32eiVcYxMqs0UvksqsCOzOdV0hQjHA3XOzQKFNdxi10I739RnsN8anRFduwTqdZZrAQ
fMM46UR8l3IBr6I3o9bRMLcJ+zh4vErgPze/fovXcSb194inkUOzUKqPQUGbEKYRXZcLyh/gMe79
6FE+iCENrITm0JyFcIzvLzitYA+87t4M1oEkiqunXEbpSeUllnZQbnnRKcnLH8yJL8rV55/CnjEH
ta2M3t9bBh2KK6ngX6tTTDPnuFoKYm39escXJBsjwHfVYjW3wfOeGcFGoRBm/KhXyWkttMkA6UvC
t5ZaZROByKnVhPE/k3kyx7ZqvFzdiisFnTMo+uxAZCbWpuTSvpPO/+CVq8sSWKl8hn3n1ROz+08e
SgfH27McS6X/oH2l7jDaKQ/ngpdmeOsBkW+aPCJaA+cCL2rDO3PhOEmcTEIn3iC5Ql4dPNx4Q2eF
nFPKfyWEYHFBmLOyabZmWw/XQ+YqpAhLvGOTgraogPp+6VMX0MRX5UZMPi4XpZXdAVJ3CkXSW00L
KnPVbRP35uSeqrf71YsliIm4pb9KaQOfIGEiKgN1J5UJmLTuSTgh2JTSbIFRutwhaV8quWabsvpg
/eEP1yffXSDWuwYkbu8NzrSmSs8gtIzpTkV5PWlnq6Lu+PMCJCo+SboVo6vPUJpnwkt+wwlNZKb5
XH3RTYhkUxIra33rw6ZsKIJwL2zkZsiD+hkK5j9DNe6Va46OP1MzJKmbN/ysWggRi7sDkq35Gl+C
yZxPLwVLBaWLcdifGWyWCVg6rhqxy9G8tgF4T4F3yweoBPOz3Knk+PnMalpZ1sSjsDncYGyEpEmT
caZKLchr9Etrs59KYOGfWwYXbi9BPK+UzazOvMv/3BgNNmR9YIv52dYCIp/w1TTQXbayUxQpy8yT
dpO19KdV0ejcNLQHGGwU1cpKWAo08V1kYVVVrCBgQBon/GJ/pVVI1Ttpj7NxR6/9jHYx2BWuMiiM
Aj4NMcuOJAdgygBv9wfr1iqK+I6ss3W/Mjqctgat7ECPyhXN7RmhOJFur1B0pi07QrwS2dRsDnas
be3EySdJOmc37LzGqCm/zLm75757zMRA0XsoulxeRmFbCB/KmGTKfPNPo8ay9rJYy/s6uWuF5Fif
9vWPgzvLyEnY+D0hE+0bav+m+2IZYTOM87HxVaWCUnonAvHv4D2wraZlACNew+gBzEfzDDfZYr3K
oRzRnvBY2rSt55sZn+T7ALRQS8eDiY3fEmeoI9rHLZ1qx/oL7+c8/GnMp0wKgopy392PCiZNCjga
vkhuQIFdP+evp+6NMjmipPJZ58wq/eyObdcvC7uuzN/ksQhhlGB8Jx6cIRygdrAipuGcVib2r8eq
HhV9lvGHg4O1CaRXKXZJN4HW4n0qS5pkBINVYAO03j7TB8K11Jy4vKiOZdDSe1A3RmglT+znTJM+
pR3KSwf9ErIXAkFlDaqswAYU6zhQY4/YyDzRP0S8kpU0XNcL4mnIcfH+hD1wOs4oYhC5yoK+Ybf6
aCdiAEnt+SaJrG2Qx4/5VBMTKk1FqScekEHzeIJAz6MFUZYKGUpXTkT+ya02HC/kIHkNEgKOAr5f
Hecjg1je9s7trc+6nhCuFqVBpBUAJcJqlz+S4IcixGMUl/RIpYUtGey315hAsJPq6US7e6I7yq7g
xuVsRlJrR43rfnOHkeFwa/oLYDhmiLiGIZjzza7TH6/AsRYe1XHz8VtAmTlZkiRresvLFRDvH5is
u/T80Hmr91rwtKfx469npecuToL+J6o7LOWqW3ndMIIuUnhVTcOk2OmSatYVwaytU4Oq7xe1K8GA
vGTxCvQF/D3S1IEyKC/vpuu1Ehwa+S81Rd+63l8D0lfJUqGvPjkqdQBLeGXKcM0xg+hr/u/klmLd
MTrcF9ymIljF2zQWVbcNcz9yQdc3jFd8qUtxVlucoGKPXzrysRA+xrMwTCsIGvSa0dkRLWkzz1Qk
rGYhZw+Iw/bNnWEYKR5zDkrsGNG+66t5zBc4ViZicY2Pzzcf1mjks7DyyySXOEXc3xxdZaGPE3Yf
lj99dhh4tCtYjuSbZrqof5kimKE7KKVSsmOVmKA+6aG28hlAIfjuC5uyyZMIfqnOD7OtY408IaTZ
qBN0mKShNm7yFNqMpq4PnOTKj9Gp/Uq7Xb/x3QYOa6fuYz35631z+X7A4MAt3U53p775B+0cBamr
JYILHVA1ZrOpPsq8kUjv54iSZftB4mh6+bNA7H4uwy6Ylb04Tm25YRDMuGm1w+geaRVS9EMu5PJ6
gdMYS7MZ1/BKQkoRttBwEAvu2etA5HuYBnkD6O2GfQLjAglWMqo4HywCpzyHDAVvHje6KCFqHuLm
zioXrBZp6oi2uCdto1gkStjdrFCKkFXAllBycvERf7Cddj7cak4cFjxQXo5rpdAV0oMaaJAbVQnO
gSefsi52cgUgiESbFLT/Z2KpRn47dwtYddVafHiPKJ8MLbQiQQldtBXDkoJjH98OkO6tV56AqX4E
RZ07jG4liYCl8JAl87NKOkDnIDC3VpsiHky7AVLN5k5nhuBJ4KkxG245tti4tShGXzI7/C73FpAh
D7UXOXcnBsGXAp61+sbHHqw8L7Hnkjey+JaYgrwLo+qwgVqpEficUgdMu1cxhNhL/qqsDNqpDMHE
xADu3doDwp0gNuwL2cB3zUJjBlQh8fIRYI6PuYc90URIPPcNeG0pLSkhKWw+JfYTohtjtAot9oIu
Rx9eJNhQNWg1/sHhT9IcsgEv2meILWBMnLycM7p0WfbiErPpQLEFEesW0U5TcbEno1pXCUqfb6Rt
o05ozNaRKcxvdiP0uZh+YscyyHVHJSSNKVzg7P7KrH8jW85UFT0pKR10Af65I/1YmEllqSnw5ZaA
WfjV7DPomiMHQXZV3eXSteMF0gUJ8XkopbsvaxQY9JKdXKmALmKEX187YMZOXfrrFD18ZuGzz3GS
SDIcxccV7RiZRqF+3MIf/eqQ/R5g9jG9Dz9QWXZIaRZ4V5yrqm5MnB3akzsLF8LcV7Q3e+TU3hDU
ayqBF1Px33AlZvxhwIiEA7qdGs3wRV2hfPr/8LcKmj4+qsjOZkgSKLscLQrawZwlPkZDDsRBY0oP
3hFOkDehuQfSz5Yj6leUl7QqYmFiQsVHwwq8vJ+YE4rReIIpiTYwLIk4jyRvncogkyptWGoiUBKu
xWdyi2HwnWao5Y0ZPK6JJGQeMQxPguXy3ZPrexnQ43F69I8IS5z4z+JY7SMkXhsCRPTPvyIadSYN
CQM4gTSA0ucoRSvL7nYToRr+qmunHrp1qyl0hX40ZWBOfAuxd5u4tbHIg501lClrxhTtoKqGz4N1
RkO99MJoIlyLTn4pulLFbAADVcn56kns78C/YoeW2Jgkp27Xlgmpayhgct7JMJiZY4K91FaChmK5
iMG51ZHxnL7Ilu1l69bOhsrJOZSuW/IumHyegUfXFiEPDToXwHZmTumrjnRR9/y9yNX6L3TI3fIM
2Xh/3Av90V38IjUk4+2ZwjyABT+SPh3K70Ww2VhtBIA4Sw6yuh+b+VPVvnNBRWqhp0ny1JnwhZIp
EYfxbVFeg0f2PmYoPiMq+6mWpt8+7DOf/9EWojbtyGXDiMEyGXlTJOxOrlWLjvkjKvAgrAkO8XLs
tIeUnfhPyW+wfynWjz/b8y26iF3fSd5kptEZ61y5KW7VCovD8He5eBIwGjfmE7F9z0qBdJh2Zwb2
YgKoYNyXBeOQ5FkYSDLv7odKqJm1MTiIhIDQahABgUhEJtIT3UPCnBfmiGJpCeXORotFWkQYXo7B
LsHtUP23TjkgAHceO3/0rkI4gYqhDThSqgLitDt5fxZHEr+tv7yV4f5/PHfGKC6TowCtNfp/V8/1
NrdjOPjljbTlHV7Ky3ERtmjINbk6lpiFRI6f8oXVkE3oXQTM2lKLCm313IMsgw8zmpe+1ZGfwT1b
921kVapoJg1anjAexLv3M52+d5Jq2D86Ha1OalATyGUHnWHnbnlQljW8K255j+WQPWZ1fj7dBW9i
SYqxPX/9EldM+w+uwUoGwDb68jm/KZ51E8LgeqJMYnMFgZ9wbkO0RX6LsP+0+KDozTbaOJvNLgc+
k0+kuR+Us5Gye4lWBjOoJ3j8K80NVAuinHwUxgyAe7FRbAHGoPy/jjNTqT6BQeV5K1QW5NHw/bQy
IVWdnNaCut4QTZ+BWWC90nf06DLMHqMRq9bk4/bZ1iRTuqZk/MoCjJLAFQxi+i4X2hA4z1/vnnY+
D3kdRWTVHe0RYNlQHDcMk6jMb3439vKq+kRlY89mYcfPJliziA8rjoB/9nlXRX0pROmJw/sTD1+y
4JnF+xMty1gBHRxGKXpSckERqu5kNBaBGLuFXihXCo7aK9KVuCrBfGpaI2ywrVcxQYje81CBpX5s
XzAYTe54JmPxENssGTYgAr9Ems0VSWsTdbbdzhC6uuSzNTWuoURpE6x9yV+SHvNLsmmwu+SCJ0wR
mf7CooLESvUz/p1nOXcZ3s3eMp5CWGk53lpmFLM+2LUDx5zI3P98gh0gbXJWeqdwAE3ebHqVzOJE
McsEHSVpe7m+jgDQVtiO8MOY5gIp/oXEv3ggWa6jxF4gSwTfYzJC3Y/tf4nEn/a/R7/3v4abHlsW
pCBLaWgeUbkPHAmL2UqtC/te1BrkqlnLtaeFExhB4Om79Eg3pJcD5dIiPgpk5irensEv4R3LtZ4P
0Quyu6382/1XGMPa6vL7J06sT/EhVTRWtuOgdhwIakWeUX84HUW7IHqHpuNKEd+gsIKb0TTIr+pi
X2Vur1JqbXCuLmseLpMW7lgahi1tIgsriGChygxlTw5Jznw/uT36ae5zCx4HCW08EG6ZU4oPbE1q
B+7iOVpJmRbuk+ObBZsUm1hoPx9+dfcTa+VPK6K4m6UAWUHsNZ0KXcO7mOw4f700Csc9eLMa02ps
wUb5hxwWEh0eJPx0Q8Pl9aaJKdRuU2Aio1zqx6bHKCozucGa7PXU16hixmoJ3j+C60MHrgwW/Bc2
hipG51deXwxymo7wZLQ7z56PqgvtnqoVaKKl8oZl6J87iYb/OnCpNvqvNt1H+woUJhFaRCP6vj0G
ZCETGsHnvkZTyOQOiVK7W/xd4ex/rJdPJ9O1imESqd+Veh3r8CigNStv5A0QJBIH5xxzK7c78B9Q
ahohGLDYIfAk7hNo7gOWnIkZ3O5F+FpCNHI/KFt1I9EwZcFYHSXJXB1Aycqntmsy6yKtvP6HA91Z
i4YmxBXvU+1VypNfyEd4s795M8KXwBUXTmW/dLYEkjKevokMFJ9Dym8Y0EdWiEnoFbsLh57BiIwb
Th4aWwd22m3oIZGqUN26D9IJRt9P+ksb7vNvVipxAV1xQngdQHT9LR8pw9VXSds6KohU63LJUiis
UyjBen3UzirPxJLXTlTpsxmiSsZVh+rDBpgE843guipXb0m+FkuamUgIf2T24W9xTEF8sGPuy2Nc
XqTudTQyB8ocgr5xcxlA0sD4Zam3hsaUC5beaFE1J7AU8RMhd8Mbxshr3bu4huoZewmLnR6PoTFf
VmiOngtcgKaHzKwyy0cKZWiaqpPYMaN42dDYasFJopw3WYHKU3rXKO1MMBY2f+yZiowsuSiSMjMA
REVVB6biU4+954l+TbBRPqZNyHdAPujJIUE14ykZcoK5CNJmiRqVUrzIE+ZwUzAGU8DJab2311mf
5Qnim3HYAB58bHkc8WqKhJo/Hf16nypH+Mnnit3fTNUZfHKuQHtocEX9Hxte6luuhbsIjLeKdG2T
DtD5Zf3Pue3Eax7zOMC2oAVLhejEoTnBXXRL1xvnNSubwIReAHOL/x3zkVyjqQsgFrE1BlQgqKGS
3ZXjiI5lOZj8PtHd+zjcqHqXesiOp9TbXZg6rxUYROlZPtAmfscN7b2+/Qcm5yxPBx6aiVwQShkz
OPuRfXK+sKCahE5iFy+nhK+O5dJM4s/pld41hmJFkMAjvuGRxnsiSS90/mdW9g4FOClPEHkLrUFo
YXPPQPdfALCIYwLNU3zQkwPGrUJRInXwi45R1Qv/2TbN+/VWf35v+5YIbS5D9+DOR+FkgJ8gnUUi
30OltQ+X/mr/xCG3Ycw5wcAQdbRg0YJpZOaXefYxaMT7nfqZnZLZV4ABOMiUKYy3/rrUE9cWTU9P
B3V3+b9F98RHRPBcCfLVze0n5wZBpOKdF3/qOfJCzRVqRN/A+F1ZUxUNwIbFXEh04i6mpHj3CBWZ
D/RGCws1qwa+BPld/Hji869Mx8rXWIZC6tigj88kEmlY8fi2N8lw2mv6Q/GoahjYnVQHNAVcD9OB
6UykRhcrS4UtBmrStxvBnObAQvcI0Lg0wlXvfwDSxv6jm4kRX1CpFjnMTXSMGcyCrf47HAV2OEez
lr3qC1mmYSR/NE+k7U2poeIDmkW9t5n7XND24kwnTZkcTF0MRFlPq1oWaszHaYwfi0OKR2h73Shd
NebY0JQ0W16rLlbjxE3Y6QX/06nevMWHPxWeS2zSD8ndHkbm0W+ih/F/mQKAO1/KFgAtFl0zkDkC
pgfLlYCHFOM6jpfHQJzdaxUBjWGRIWa2D4SYpR6t437lxCrfAPofXlDF4U/PmI0MfmdXokmfJ5ZT
vI83rph9nxCXWU3R1PIiwcR8vLpnRnP1Ew2AlEtrET1UfWSrM58NaIKlJc6iU2tCWlVWgULgVMf8
lwPaaRNC2Qd4xR9UQzSkslb4OojaZCJDKSYgQbsfTDftuya/soajqcnQkVDP5QLd5KDcKXvu46b8
Ub8L3qrQrXQJewlNmMlAjIDrnbn8exexaqdwu9Zbq4lTInBbrGENOMWAK/I1ByH1ncVDcjWKGixs
LOMk21pqAyo0MWswG2bMpymwE5jVjpTsLsYiBAEUfF+RDoUTtCsT1DUrL1hxOZXm0udyKEDMAxNy
ASOZ5nnZH/+yvFRLEytycaDy33RntHUGILU0x0zsNeY5Zm1kSI2uu50VqVsfMh7ZZmSUlcofbKSN
FLYT19TAnDFXUc2DoysIHty1aAyN3dmbbYCOMyXsjGoOeKRZem7lsW3U9oiTDhNo92jWB4v2PHAt
b79BKrBKI18GkxImUDYtCQUdFENfGlv8o0K20UeNRuP38cqcUwKleAYcD/xc+TLI3sHcOYT4peul
qWji9aXJW8X9kY7v9XZjVMR0yJQZuiL5DXVvn1635xFcg/zYPb2cphBKa7H9joIzhjtkFHdIITNL
8Fnt/3G+BDPfdhr/rerzsYuj/pp6PUEyfeWcBBYiThQpqc1CAJfvg30CqmubRyddRVhP2ei5OclD
6sJFulaUprY3H38Ro6PJDOctnNIVjglJIYjdhoEwvsg2qzYIW5iDjAQNBd87Y9OJQVEwB0CLjac6
Fb+LOVq0XkX7hDBZAK2xHLI/kEWuDTk9EGF5HsX8/LMUlSx5Xfd2IDuyYhjPw/GJZCzTm9E0xCJB
7Kwm+FqrIpoA8Zac6yXsGGsYGZD6J37CMBOr+gkKKhA19nSBiui2l+DLqrNexKxRJAkbsLob3TWw
sXU+0vzn6qUCJlkhgwNrMlSPQw37sJ6f9E9xjYQyYX9SICHU5KxLT7Ev5MkpUO6iY5xUPrB6L/li
WQff+3Cnu/zCml7kab2pnH/T9WUCRwl48c1olD7znI+TTJXjpdT3PMuQukOUXZElaQ364k9wM+gp
YM/cLh9L3eKJf3kxSoOeC6sNO9kVKBPQ9s0ND1ddgJe0XOXNf6mr/cekrz2kCiuxZ9/WaXWOw1vN
x6sNASBYJq2rQrJoc361DrqIE9aicW1+ukdPFno668TwmPiw73Yk87aNKUqw3WkV6qhx8roqjzOE
iJvYdLzMEfdqp7jVdnYBX4BGF8KYmXXMb8AelCkRp2f2lEksrVAIhNPAG8gN2MQ340O9HHcYlCv9
Bit7eYpCsV5toilZnY9/8qZrQqnm3zElX8gLXTyNEmH1H6MkpNRxjoDvYtpBzPElOzp+C65IOAB5
0lNWxkxSnhFz18kriseI9seTGC8wY/3bJOsId3K0K2UNllAetspPpUeMyFI8VofPnVbZ0iaBx5F/
cCCmsK1EqVPOqJomr3Gnb9TJXd+sFifQIVQot7CcMqDUjWbMAIB+w1iSY8KI+hZKkB9yGXn3jE3+
6eCFAaAk6jc/7VFrYgxuvCtz/voZtibpQPdvmBSCtKe95SLKQK1RJ2vtH2a6B976JwaaL5i3Dncf
KK20fTJhmT0bubMpE8tBVl9kd+RnOo1cf6Qsn6Q9uofpByCIWlYjwnPVrovdq5equDyR0ffFoiWR
PMmdkrm63o32pE9sSNSVS1zx+eQbxOcu4vTNx4x31+yCnRQ3tqS4UohSpEEqCUOsjrUgE/AKJJLW
qewetDqXW2tPBp4/rhLJb617heDGwe6ZQAE1OUXQt7iQf1aqhTYIJAY8s7Qju+hPVOTOgb+OSBIr
6/SVnzraTSOMqQlXm2IN6yj9DbLaTHbXLsDBiLJ5dJ8fbWKudN/N5+OdvL8QTsqJADbIOBZRFBLw
w3TydKf4+Hhui/Mgxg3CSjKHFmZ8nLqq/XE0QRh9huG7xirf+jFAbNjobol9zC3h+KPZG5pCEB4c
O3XLrIYXHkbEWCzkY8TcQ/ULghtSjqr2JdbUJP2BMMFiR0spjLja6hKofjV0L+7K8kn4ODftB9O2
gmndjU6AvsskyZvcCPqBXSrPxxj6KMqjqyWlhLdHs4mnyZ74W/RubDoz/5Kf34FJS8BhzYWfFG4R
sPFgZ6mxgMtRQvmv31m4T1YY4ZQCwGrRsfOIVyKi/QCODWGDAwsRX4FbrYywF08z6CSIGPXNwEoO
wiAhJCEKLDOD+OGkQyWbs8sQKtZq87gCzDMLOkPPU+SyX5LIHkylNtWto4W6KpnYI1zEqpbhpSJY
N71v/+oHCopwMLZaS0UHrnKS6kxS5+Mshg9mTkYolCb9JaBI9QBDuf2Win4nRIvZxorIs1bZEJVs
p0lIYRtpSrktUah6DoawRaPfp8GJUqqrtVFvofQhv4bjTwO2m92kZ7s1FbiYu7qpri3A67UZPp3+
97xfEj3c3NFG4zeWVCnxlSsRAV6C2gRuy0CNrA5+TvyOny5XnBu5KtER2aF4/Ecml64KQosnXZf3
2RW6HuRpCjzu/4gLgQt7phuxhovuWRykx92SgzvPxVzAyDBgdHBrgM+c8jPtd/0q4PtoM8iJf8UG
7AZNQrXp+qagHg2xH4vAXeH/irVAUgMEbGV5SLQXngl6JPSbH7m3s5UKrzm3Mav+1cjrCYJDQaQT
yVfNZx95FmqfyktRjWlMKOezM8OgnTNsKq2ukiNhZuxCn9iczl7osrlCCjzoo74gv0M5Bs/b/tYh
D0rR6RwIf8YZy/SiXU4rJUpXiH1p1Dq3udXIRT4vforGEV1QPrqgN/eY11FhETbDglk2NjYA4+tU
k2XI1t9K0FyeUQlFeASt4N4B0iTYmIZPGCijFHgPOZe89Jg8Q56NiaGmsbDMln7dbSI+TxN89X5F
FPnGqCAywUISemFFAGyzt9fXu4b9TJpppIp2O0dPRWT+4Uf6snpiI69rB4sPu/y+NPB2yZQgrhen
02oNNMsj+uDzuSlAmhU6X9FKwbyj0oqelAA7VerOPOQymrJ1wtTLKQYATPVsq1emrqLiCVjnGSkb
bP7IE6BAOgMNgGzM6fa9SP85FqF4DqI/1DG7v7q1bXywSgcYSHvH3fl1KUp59MhefvTnq555g8A9
lzpEOPNrhGR8ZTilaF2j+oCx8phF0nYpowAppDwEj5PVdCKjVpvkc8iBAPxtjJ/PqqA31Fo7K2QE
3N53NWVGpY3vRoPInCOSF6JrafWds3YLiO1LDI8X10AGa/5ijAqpmtDNTW0mH+ltZTHLV6PK7wD8
SAWY7VghclNTQibSp6y9VXumMtnximh1D11FdJ4ZdAoyJshOffUOON7nYr9WdiwI2w4L0sw5em66
gJQ36FdLkgGjf8NjLJLjRb/P5k7Rp0TDQh0TZRBerCJSk2q2p+ZmJFzG+zAyVNAilGzpu3TaCDD0
UgLAH3oWpZLT4+nbWWK+2mUsf+EIfuRYc5G7fKteJXODp78I2SZBCxaRpgtl2//G6VHW27fXnUkc
7rMZwjtixQeb1CU7HIymf2cBCgzHIXS3iGodGw3xCgFXSF9IfWkrSs2TLnd65RfhjU6ugNFrxpo+
SRUrn9Pn9Lmvc4jK1W4ZkoUko0gq9nciyzfCyJUhHmjqAatWJkZkqHZ3+QQZiJSwL+8AclfzBYXJ
r/td+ZXfKNw11l/5h6CI3kETvS3p9HXpScZwCTxzYF/kbzo1iXUCMAzVqzRdaPdoEmOb8+PLCb1U
xpt2heig1+ibq1zad8NvDjvfhz2jlnJfUOykC43CePjRm3LHiXvRFb5k+Bo4KUa+T/ReRc2YT1s1
uZQWoloPLdsRslFQzH/faOeLDkCz7PAKIpaylL/xKpfb3hmnUDmvWJO+GWkddS0pL1SXqHw22TAJ
gnmao1NVQ1pQDB8FRw5bFeA/Xkc7N3TMswc0fUx8HRCc7dGyaDB9Ed6GUGj3uF+IXdR56elZ3omE
bmKVWxTkBbWNuFg/lMuVO5VCOKOs3BMQGwKRhlVMetUq5Hf8Bmd02fiPORqIn6mfdHgmEJjGT20+
lI5ZD4PJi1RIrCTpGpamK+nmfBWQ6U32oTjvmlP1oMKlspXCHEALVjrMf7Etw4nA83cExPvoOTBG
/KxIiTfLmfI9PjhLHnAurb23+oaATo+9ZLN1et+JZRSW1BWma6zyiznb3t6B5GxRPoVl0lkUeN6T
pyDXPixPsqFe6DkYkVbdEnhI7F+pX+/Mvcj0/8hzkqjrO26wLBcNRZLpr2XgAEvxym0d1HOhBkH7
quQV7K6lmKURT9eh0DbkvNdub1yeaV8MVIj3gpkiYYMPsCwsQEijjDwjPUwvX7PoGYv+RZxmfq0v
zez2c519PcLPakmT/Tby5HVHymlzUMT5O5CNC+Ez6/O7LFzFKLAHFyibCHuDMz7oka/7SBQz1goa
WCAFx7OaJ+r5yr+v5/JDdcql2vrsPSa6kCTBmRFJCaIGzdD5zR8q5G5jiaik3wPF3QYryNgFdppM
P6Z3snMqBdeQwCgzoH5g8vRRLf2xDU0dAjAB5YKajD9dTKil9V3R2RP2/uoT/t7elXrv1En/9hP4
czh/21/nX9AdWlxIfNeIBrcTRElc5Q+M4HjP6Gq9MAUnc8RtmIet23KLbLqJEIk3+JpbmakWMVQ2
OLxQXHF4wChejIgrIwSF0AiOvn2Fii1GW2wxhz9ZaQG9Yeo3SL+IQHckvvxWaWS7Q9gLfUL7Q4uS
ZCSfje9+TKy/6TlSQ67rE3b/ZiW93JVytWZBPZHdvWUWxDdaKANrr1qI6VtzwFMQqnDogmJIGGi5
FLA1+LA6YZ6yCaWPv4yhKlC/abD2Azc4mMUkPIBCdOh6M1lkMZfsgpHvqjVHlZUq41YO7DYAZGA1
nb29TGXlb8TtJl3ysdg0rnuK2SDaEA4UjcO5N+gsSuPgVUhkuahRRhisbPvMUxjMQ3b9WbnwQdTQ
X8prgwHNzLIo1jPpkwPIFhIXLfHkSHNItCHQtUQ4GikETr4g9S8qsZhnhrVRlzy4oZH3CA6qXoFd
iAVO7BDZyKN8wB0Js8UAASKT3xdU6y8v/t3r9cN2QiZX8gd2DOSNYVe1CugMsui9gnj0EXcZPHNM
18OtkCUceUzW6wkD+tNDYx4MvDujQdac45IOSaEHEGjW+sp/C2WIE82DTCgihx/XEZNzU8mFHQzz
jOwVBi9H2JePPv4FGKdBhovXhVwe56EzALZU1Cinfh9zfFngczD2hbCAX2DBJqVlG4wqy+H5iatN
K2q6pcoNFhhbf4fR0v6zbTw6+MNlp6aSiefhYr9Rhxzaq59DCDG2sXabOb1XGJKj9n023YKMRdLY
AB0Uk0Y/wUSvljNCNUZB36EKgEOSagK9fQZVTsK7qEYtuZ5rkd9H8NfD/752F+Ya6sAKQ595a9uG
ObmYDNTmgdCiTKURCSEaaSxckS8O4MUFTFOOrXlj+Xzl2tRsaKnkNY6VFIobd2+dMFtzNOTZPhtJ
NXt3UA892nfJZDl2eaUW7YDAc20RE0lCtU2nILWyebZgHtzDhUlJhDxzfqX40MIFKUoaBMdqzCJf
JrjRI6EPUrJqPT46p/uhBooYJFt5sQbgmxdQipfU4vWxnb8hgZqWKJpSYCwJYmHM/9Oj1RBgC13S
xu7oY/yHV2YbM9ykXvciSgx7afxlj7Uxfu7t9BIh8jJWo25oexScViNhMqEXIWpUQvVVHBTJW3ZF
gxg/c3TZKpgSM91AQvdF5MT8OogvKikqs2YJUPunZKTe0n0xZn2Ur2hIuiFYdl5bCHyqsdOpTgXu
y1O2AtH2tSQ7aozCTZr6sFfB4vvk7iWsc7gA/oWjjK5ys0ah9u/l/Bwvk2zwnrba3D32OE07Wfur
z9Ajf6j3gXBFip+ildlD/RpGjiUzDDd84KxQ/fkdLkFt5YJ3pFL2e3DK0ftFmVmJmeR7DWP0+Kdt
gyhTAZjXX2V+bWIfOXymDz7Sj7WJDJIgw39caQ5qln58Wp2YpYollt4MqcL5SWuqgIAkOPUpU7dU
T+Izw1cCyzvTXYBHG3nSUdZib2xGzRBoTpSOczmcMlKPciybRRqYzMhAGd+6Hn/fBdB0UehpspJ2
qIszqE3svbQclD+lXeuJ1vUME/3GYPQg+6MFMyVj5BfF5T6ugij8ZHexQeL/frYkaM0fHsxAd6bo
GbLFCfq21N6eclwGjF0D1/srVxXukn1o1XiZX/LkcrfEOs8Zm54dWbPXmwP8H6gfZIy2tDZ2nHcd
63sOJ+qywFi+nmfm4IlBslZUsRFr2YoCuVU8z0SudE+qQBr3mxnpLuZyt+BzrkULG6nxHmcbQsI+
UhP44a6a1mOy+Vo6EUpDLp0TH2UuKnZqa+H6WV2VBoFEBS0wrgho+GEZbdl7qJ27HSsOE1QWaxw/
psja1+favqWFz4NyM1JgBaDB12M/A5Fb/kPyQyOt9/wIlrLAtMR0AfECH6Sn1jzTxb7Bc7V7EiNi
D6eE8s4xHrqSjbY4HYQ6h8iNMdRwbRapPtae8cfLta660ZVrNZhKKwDbhumgga25koA3p5MQqBqG
26+448ZWrc/msa7pmifEYjcT4uWbm5FcQYr0hpaC0atpcZrxY0tIV+nMKqY6lYuLdKLXCtjXqGMg
nPUzMQMLH/Synkgubn4PVY4Eueh1HgojKUQeWrgcciVSPbuEj26I+BlZHcOh3ll9kgHHJzog7Onk
+BzA9TxOtOw0YhFoAL+cnOx7pN7/tIbgM1qROprVdKHSWe3qcS8vTub2it2Tc9KmEKUAUizp7FRY
KW8H19ZHtK2oemtl7x8uDTyVw2OZeBQdK1BjUJHGd9bnwbdP3uegNRzhXtfeYAMvzNyTFWqSScV7
vE1RGqzl/ceCZkiyGO56UPRzRXNA2dYlEqJRfPrS1r19KBXeO2yzut2jeAlgoZZbwppLtO9zWPdp
oYgDXGIkVpyoqJykpt46ebvLZpA8kEHv4Y/sWHh+SzucTcdewafOqgFvra/Bt0YZzeW1xwnYgCuh
8xa40yhR0xIHgxVE7FjyDqip5bQ4mBJHTRGCWYH/qtjVR501oTHKJWiNYE36jLs2J/3puv1IFB/O
KE39NieFZKdLQjqLzYi4RU2VVju1qBCyffyLV2RxeI5sRv6qRQS7s9MacZeYSi+7zZPCCYe0Xd1e
vCQbDwiYFcKE2QkBTehA9lkWrcnOL8huGPmBgIeeEnVLgko+drt7fAU7kAsntSUg+HeRVzIZKOCS
3Be7dxMRo1Sc70lz5SItUsr1PjhvmBKZWg2/sl2rXg/622Nk1n5U0N6yaUbrVD7xRj3/bb7aoSQS
75NTdqs9We5tP72aDnw1Fq2LNv6/z0/kj7EImnx6xfhBLbPpyy1qIqcCGu3RiTFuZ4uwm/rcGH8m
yAX+/jShoDHQlyfMTtE2qqqKAzdgrdGP7/njsi7Sv/Z4e8NLhpTRmrTWOjANS2QeBuY6gWygtBip
+wI5At8xIO6qyLzl0tO/AC1o7LQwSrJjkYNenoXluKXG1yVK+RRsIrgK4BpeMERuC/N5VdISeNbg
01BBW7LTP8aJTqU4DRLTDTU9LUJfWzP939hPfhR7wPl97ro4URe4N3MnASj+jtE/fr/TxaADfZmi
p9rjzhYLRrwXCmQ8B2IPgYcE3zEMadFlX8vmTYXX6JfdJzG1tOiL9w7TwYh0zuI2F6nUusWmW6yn
hsGBs4Xdaq3hk1LPfM5Rxz/5A1SHt6Cz7UNyz2tp/od8jogvoNHhBEALhCd7u+NrlB+gQePXOCbe
NlDhsytXR7YXmK2405YJ+3ITp/XUYOBpmhPyUh2DfqfFHaAyqCpOC8GMyYk0M7nNGhXV2WNWbzLp
9f1ec/0MA3h2JNnUN12KeR/3PWj6VD7EUZzjRmCMLN+KJojEKF+VCwCY+2uuwZ3R/om1WBxYJt2t
Lvj58iSjKlaDRFTlCqa7UvDtAkxNya8c5wFE9Gi5Xv7xdIQBaza+tZoZ2h03/EkfTQ3yjsBnuk95
0q9JA7G6Uxv7fIok5MhX3lw0LNE09G2o66+uW0YrVXJU+/3K68odXJUm7JFkt4fOj0/gu0VESeGU
D0rFcj9qtQWs9TSSSL3NwS5BAPDoy3I81pqJJgra3/0DcMJYgcf2B5VJrBBpGeG0I26STBRo7kbk
ChoQz2Ez73LCkSJiOO5lmR56tCb7giu3sgn/i2BPgzAFnrjsIPywddOWbRia1OZG+hVLXeTjk0Sn
WgeDGuDiJ11ejYU8U7HfUab+QNGO7M5Lu1v5RgCcPbPxrx6mPvHMzwulHQsvGU0vxcAPPvx3goA5
miu95mSmzydcAep8R5DpDDaw6tBWgTEtLL6sup9hEnQy2xh3r+aleoqFYhcxoIrwDD5MN+5ZnmaC
dSr1HsN2/CZx6r7R20FiO8uLIKqXMqsDasqsd9LunHvazHyha/8vRugXn5jFa01cK163GmnBOWrc
wqZfLsnKfXaJNVyQbBMOiRaPzTeR9F7lU3iLVy1499XM9wEENkPk1TTyOeJNoJ3Xb10jp5yyg0HW
OdeD52TpObAtCHvkM7Rwwv6bUf7HDxevJKqxkLNkI119GKTBZhAsaUp7Hm6Kp4D6mAsmjSxfxrty
KXCIDRGcPINKgQ3xG1MDofQqtgMyBiY73WYkzHqwkfZCq6+GXvTAbKQ7UzuVvbu3XK7rmNX7iBZn
cSAjLgsEAUaM+TzGu2jRc5Xm0vNLJ3i7uFL204NactUjALZQTxk7FeQ4bXxNv5/pKf84oQqXeqS9
qE+dREIcbAsbBwUV16a7H3p3sY/UUwMuG5RROBI5FcvP3gjOt8EeNwLoLL+s0jMzENdG7tTMjZup
bXsQ7nAGa9AdIC9iPILr8CIU8XIh0olOZk5WDAaWMJPUzAdQYuwSPdSB5jp+Lb0uk85rWZUHOEa3
xUXm1YY6VVq58OmmRgbHZ8AD3/Nr9XblIM//rsWQ3Qtj6XuUqSW+KQFQTivGVkVLK2e8+YzUFGHV
c7nkhu4jhreHv4p6ZqI8/QywBWcxLZZTDBHCruZg2tB8nfi9PZnhn6p5lals2NTfMDNrC9UPsU7E
gRfmOIr04w0UzDCt4/Bkdp+3/aFf0wnuxKdMhJad4n4iAntlC9wI2cdxImOXQx6WMHxWqNl97KF6
oTH08BMYNBdHIcYZMAeYOFCeNsSe98USBk7POLBw0dJB7+eAbr1m9ueon3Z69LkaWM2ImSAzkaMh
MIdNpv1nq0r7gOkE3H/mA7y5rbJMygcSk0Yh/skWIHOZRQticl93P+cB6MyqVYu3Lwa3j6fANmc7
+EWh0QPBXY77JoSF2WigOsFVmDVRIyZy6fPL1SGzPMP8C4nHeZbyGs4pd6whA2/ooTVkPz98UFas
IDYlqO2LZplIZ0+T4cxombub9LXCgC1OI8ztu3Qt1G8AxzJxzd6Wfhl/Fh1Ff5ruzlfI4wW4QWOy
+ndRQoFu0K6z0JxvUOCnwESQe4rum5LXcNtvHziaYmY4D3Lu7hUPda6yLhblH0WZjyKM6y0fTKt8
jvOjWqk3MQgMj9Nf5NdYjKqUXk6PHl9tjOoz39lSRAbRi6ldLmemAirEc/GWQmTG0PK0FSnLMRIy
+5Qnq4rEhIU6iCG/uwXkD/L95kT52r8iIYtZ4jecN7osBklRkapzn8TePobdxSZusGo0d20Czy8K
PwGh9JEv0lbxg10gMPPWFrNuLYc097gB+U6rkI4JybHwSIFtY5szlqxL2KYLZpq13LxGrTPhfsLe
vW/HNpE2x678JAA5F6HP/OgRM4y1GXk+mPserWvjQqTXYbcz8D9STqzmYYMIcH8XF7ru6kPeeZY4
FP0U0fR9Kdqbt7kOQWAPkK9Q/BkwAyvHIIKsk2PxEFARpSotnvwCR2bIVyCf2ElTgj/MTxw/xdVu
HBI5Strjila2QSQK9f37sog7a+PpjWjxYlPWBosw0G/jXt95PDvE2u/c9i4VVI8W2eIpg7Ahdap1
5HDHqTy94a+6mc6uEhBx8cBHBCAR69SOP1Zo+dQ/jySeRW5iQz0H/VA2vwRUR2Xbw4BEXKMzgCmm
lK31MpS31ichJ72kBQwpgSXlRNcjytuwfRvGwW76BTrM99pSgmtSq0SFajHlHDGTFhOYm665Un6Q
omK9DykE+0RNO9+u1/KbejV8wOg2+tYwTt64/IvFXzWSz7jgZj+SBYM1nQHrMU2V9qKmzJOlwHPT
KYv5BRY34FNB4FldGy1vigV5sRpFDAN280ap+cl8GAU1dShYOTKTscjWja0NC4bAH+u+yUVpmVNh
OhGYZX6itH9JnfU9/E4y7YFlBGupw1ruYuROqjpLaMzaJ3XjlWxrEX5ehiEBX28dk8pifYfYV7cq
omtM0fv6PStr5S6q27s6KcKUsIp6ShNzpgEkPIBCqE+3gjqL2KN/A5DGTJY74me/AraFqYySU8WT
inP+Dngutfad/A36MkO0UrBsaTF3vth+B2nOoWWX1uLD1TlnU1uflCkZKAcnuYpDinZY+LBMd5wl
/+eSr9cMhbpWoR/FxMqyH5Xg3TdFDtsjKaywsd3QiHlCys6L6qp/L/L1NS4U5M9LDCN1TQgEZ+y5
g6dphQOcbyRSlbdCoaaPiTKg7g28+I4emRkWWcp2J9Wt6a202Suvo2rlg8Pw7BjTj8MmgUjLMJtz
FO/vOy0D4CguOKoFZjBR/yOktE+gm2FAWf05Buhsmr28klndnmvnubcQUZoFua3hEXdZnoKan8GL
z0AyFdkG6/Si5rFasgze5KZG/3gj78TQxwlycN1R1WLv4QR2Rz6uWntDYimebuuUMhdU0RUeU0CR
uNpVPmg0k/gj4NsMbvcW15LjDnU9levuqbwFbrqSK46msPW5cw+YRwzBVs4Mo+LRH+xAnjvYAqf2
4CDNZapT8Wq4YRwndr3loX+7BIZvP2Z/aF4Ymk7u7554SIr6hbbdSWZVIScHGWLBxGenH1kAsXA0
m9dkD8h8Pk4ayoNEYEaKay8qEbFBVXQUB4sFiz5b8sfhpJA2P36DXYBvyDnvk0/HDvHDN4QJDXiD
wdIefgBdiWDsvK8PK1LJb+/Nbokin9JUElHJNoa7Izfj9J/5yJDE8IohYEBCABHLUQXmhhQLOqXx
IJM5FLgoi4WX06mNTYZ2lOp6/NFNCnxf9VeFetcVqWIWJdX3Hh2oaH120MqUE7VEm5xkNFl5BeXw
LAPa6kPIXm1RjuNVZnIL+313KWzAYgBqH5C6A7fSZSYePZZp23+wserxxVCsZMublQbHLF7t0AY2
edbPzVn2DhPUm14sKFbWy9E/PBw90RTU1yGYVKpqgws28iKnaaVieI/Za6aUlNMblYEWSE1u0825
jFCFRhPu/ybc9cRhnFB4f2hk6cJQkePRxdnfjiM0Vn+oQk4TVtl6b9RdmznH+E8w1S1tAPIcq/96
6/xB8kGqf1Ud+fHf95ky3zzz4hZ/uVL6urqIHBrATW8GJUUWNELMs5ZXH6ieD8pEdTFOs3wRf7Ho
WhvvXijAwcFdlzqP3G/e7pvsPye8mq6rId6NMTyLYf/+PUWoH0TbYNhi8n5I5X40UG78m8feIjtj
S1zjtFifiGfBxXU7p1/mFxeJyBII3Q1v/p6BO6Rl12Jt1qWjRT8xpkp/nGnkbU+tTPvRZqp+Bj7f
dQg9VKpAVEwRh3iXc8NP4ccMTFU/NUt4gzyn2ZkpkLtxRXW6p6pZvZS06Op48kv2C12wPLRXuJbP
EEtTbek1xco8d1cQ5c/JQ5qCP9v3EDisjxsP58/HM9aHwqOi9awe+pddCzttP50jgkio2Xpo7seH
E5OOd8qxsW1U/FqPn3QcGzUNcNzfhDNBvo5DzszBd46uMa16RSTw0I4+9JQJGsSv6Xw/vfrnBWLp
S7E9Rg9LSB2PcXc9WUDMjeg6+zjic2ci6EnselHUGEwz4UKBXdPGKKROx29YVq3tYTMXNomBSVFX
7YbSlBreqzc33JX68AIUgV02J5E3iqOTl8CeCYtNdYnx2J7JUZ+QlqEFjmg79tbIShR/eDOsz09n
yNo/9xksw1tDvzXFihSGkW7Mj23uceoQ7qO6wI6d2RS8sPk/5bqPVTwO30qCC09Q3mx6bUwt8EAj
dTd+arGiHsU64wCWVzP+zDqKWh5yIIxrc1qLCPixzXkhiHbwBzd49SBw76OkrlMRQhiNkj6i4y/9
oYZLN1k6v2i4By9PkzI30aLJVncjffYWEAabKK++l6X9K9xTCq4s/IwtGjvkW45kwds2k/ZE2fLS
yG3A4x1pDhsIn4UZCHK4L3DIIcFdn0udcWcFyGWv7S2RLkgZuEnUWc70vPnJpZxnK8sb7a7x+dAc
AqfF/UI8ZmmGh0kun32hDc7O2VSF4o3n2goaDQCBEbnbo3m2nx4eBkHkbYmTIfpWEwORbpO3BHOi
ne0FDij0ZkRBVXrS9aFSOMuxjoKKQWN8RASUymGdhif3k8CQ7d6hISpQNt7FdqswYhh7cIb2elPX
kyECQruyVbLx4UTTSxDp6cIY9eoOY4U/rq0u5t2xXZTSKZTP8THf9v55oeoNwOfJZpCv85nhaldS
zRADmdTxVFOYonnAw1PTrgWFlOX3hlrVVvY35OsTMdjNm48utnUc7K8/jJ8DWyN6smktyGZFmXS0
jHIfGf3ZN5sZQfDJ5RyhzykAgHQ/3GC6f+BLZuW7mZ15q2NHI4vze/x4Ahm3Jq8UtIkw51i1y+Yi
fmpVpDb92ueaVhtMuqAaxQFBtL1H+rd1hIJXiYA73tloMURv6ulPFMM26vuwXO9qJwj+1YU+aQ5L
s9V0otOeEgeiz82t0zimp4xX1mmGZ67FJd/wdoRJWeggPhBk2+9HkTEv62S6t5sLhaC5T/uUXVcY
33H7CrM9sEV2sFRfi2IaK8GJBSA8YdC15jqC33aslv3FdctxL2OS+mXB2EJYG0gletFZKaRS7VWi
VgKecIR2yc1keV/pHQMNbY0XxWwCkLVYpIP4TrKJd6059XzcKpJrjRjCKYq2S4QYvz4rfonW8+ZB
bWGj9PtKWvbQ+qN/DIZqlGCLnM0lMmJePUZ5j8WK4NfJnAShvF+yET9IWv9zSMWU4+/7TFQIYMMW
P2sfzULQLrjtvitKMWBQchga7BcLk3oW5PIcGERIWEKHUVblFMSpbKZE7ppkZ971by43c35658r+
6xWvBvpdUFWjC5aNYxel2HxH6UMG6c+kkRn/X/qrR8ai+MwK+7JBE3z43MvBcOif3IEnJYkgxMUR
N+FhpEDlI5CIXR+Yc61fcdMkPrkRrLDe5/cGIVa7faU7eUZiuc8AL/vr8DaewkDB6UwTgCAvGzgP
lpDe3QAaAD583HVrxu/A7cVsLnJQru6KyeAX+eAOvbgVCqdNT/P82h74d9uXcm8h1nruO3le/kOD
7z8DwiC1HjGCtygw23SAQkXfJ+ZSAzT4XyO0d2uBSZfka2UJKUUOr+86Qa4eAc3fqF0h2ixO7mfl
LK7H9/22gK5sPn7qPwnlLaBegqBAKQN4gIDLx8AcAEAS5wYz1BezNaZDUc5Hrb4W5YZiLYV7e2/v
Z2ikIL/9tkrf7O8fPVwgcYqBk4NBbIHWRbpJIgB1W31SBwNG2dIn/8MaY3fSUoqvd6LUiedr8ZH2
k+0XDQYQ3Dh6xP7KVWNDAO3KyUTYvs6Gxktjxbj5VnLh9VOAQdpTxfrG2Ay9x39M6l1dxP0Bt61U
tt+6rGj/fuSB5TUEFwdXs9IH1dCjIOu6ZDA8/xdxZjSD/3rdE1eG/3zF1u7d9ZrV+E6P63pXO2wU
NODUy6WeVs/csniWQgS5xQ9qU6A7VskWeX4kuZ7nR9mTfYDQoAaoG14WfHAIpMdbGCY7zHucm/hc
8xTPuqGy91NUWlpyeiaAVLxuJ5jpaX2OQvE9FFgxnIa2/iXUGZyot+8/rSs8g/lwSc6XFBRTvI2R
P5vTNZAnCMYbnbS7WJn3cxBirSPgUaN3ipphisiY5Cch3F416bQhU+biRwr+M3o1KccjakG5GRzi
uEm0CXKuUHmyGbiHKsNN0tGQuoK1mrs82rro4WQXpW6kP6bcjT54EXwWi+FPXoLRNH2Za/rf6nsx
ZzyuB/6qsGARjdNUr+G8ddoNX4OuA8WfSNCRG491oXr5IwA3P3H+ZXXBZ+w1FTWJNA6s5c5nUA4Z
BWXIN4xwll8GzqTyT4V75Gg+4osA8uRggfGsCcLevh1bNUEu82Bd/pjQgSIr803bkwZJxix2VvQQ
LhMRndPHrTEAWcShCIAWMUT97mNlfOdL+VFvl/KHq78wjK0REzdmGtaBJ2z8ydtp/Naelc1EQ2DQ
b6zZoMNGyF0uOQTizE8r6PBKopNuCvIVcuS+7lG+KdyNtdLTaUNUMYsQlj9jtsbtCUKtZYNvC6YO
DcH2R+/R665K9WNPbl6MTS7UgIxoSAEkyVIWTdgME6jhUekLXIzZve59VOidiJjGNatynGwdZGQ+
Ig6grvYdg8rze3PNpK/16Z9nXh3KmLunSiMGgHsGX2dtHhTFKdc2CJTv1hVKe13POVptG2b2D9Ia
aMBrqxIV2/RPIjM96cc8GpicNd64r7YpST9CGuHy14pEneGtg8D3Yqm9c+uEgCYmcjH4zwmJl78d
r4l28mZUobuU0q/0jBsC4Bnv8XEenkAF9XGg5MPuv+IHWpqPtFFU0LiUKA0uV18LnK2huVM5wQkM
Pv9I7C5Si/Q/ndfHkn+zd//2zGlnQrVdq/X8XbzOgdBStX+S71vGuf41aTYopvf1ZNhwLe36v100
+lIGrhdAQLxsp7j1+k7DXOUJhWa3pgQbGterd40x7nVLlCXCSOwuvfmigoQEKh+thJsUKpmcuNev
oK2I1JhU2YrVQ3BPNSpFe2KMTxs7CuDlJZEmHf/bzSOaM9aO+EC6+vAkK2DOoQjH2VHHeWVa8K2O
DXXHEXsrkKvWe2rHejAfeUQihGNGp23NjDDQ0VPnDP6f9UXF71c7c71iwgN/ubJMIpWVe2bMUw4n
XbHXJk1nt8C5Xy9m3honNxGty818Dsli+ARbN/JOnC+QnkaOgt4MsGIxj/57j6kPHEA2RIqYtnwb
9CdTuwZ5/QUUTxCdqn9SN4cB/xgWjzYyjTantBv+MTe/rWbKMT2W98jy6OqEjI8JMPpKcSevbZJG
u5+7sT6B0JABQBvyZoK76+Kr0LI/+qRqVN77EpG5BH2uY2xOtk/L4OxNP4whk4T1bqpGmL5u1oYv
CMrQasIKmC6a85Y+KY8QM9Ad80O1LC2SM8rxftyml3DDKeYZ6A6hojJ+E5mMUwvFboRj4u9QX2tu
0sIK+q747yu/Qb4p22pF9V7/2caR7wLF0NTs8MB457tmFeNO44Hycjsd92R6iUGFHAaESnsLSvyb
Zg8MlZoe0UskmH4FaFqlafclyoqQO+yd67aDtzsn++bzndmV8K/w1XRMeU7ZOR/QRMZpykutXpn0
swbqq653hDyOf7lp8V5pD/NbpgcRijI29bXkRFuZESa/K3PxHGnZ+KJGzdRoVlLVA8haoyU10ATy
Y7WvyzYXtC/vYA04mtjF44wxtSyaEovIKesHQmZQcvl17zAHiSRB0fKKt7KzLpMUjU2bCTqNy8Ix
z5v9LnBKZAVP9THBWk9hSYvzP1TPLy+I1acUXrrBvIb1p4l/ZZTgU3j69NoHeoImJ+Z/SyVM2yI2
LmKAYyhLm4s0o+JZt3oEWl9tIqnu6wep7Q8FeDUb1jZet2nEeYgmKZ89HaSESPXVHDXYai2nICUP
BIlf1m06uBQHCI/Yjh+xJ8Qy3la3lig2ABTjwM30RhIZn8KKfDE7sNfoLmlZGf7YT2AlZst0Qvpd
DnKR8fs2etLX5r3hN0oY1DabR7Su3NwRiTvXUlg6/wxUFt/u79cjCwyECLdoRrqY7ICKPkK3G59E
i4GwAMa3COHrfMgMygturKG7xn+eIT8abnpAInjHKCEZI48gPGGMXsnxM3RJrFyojwVQTAMpHJ1P
z7xEfPdBFTZPQVDmefLtSxNZCJAyzOqCVHPqZ4/9VIJllSEL1Skekm9cg8BBPksOJ0J0VDcqynmW
yh07hs4Nd6Cx1bqPgYu7/NIxDM3u3Msh94s2vuX/xrDIcjL4Hi90H8ptfAtxPyqxIhenKGXgGXWf
7/vwo1q0QHHYKAS+ot0Q5LOynyVs+dKeqffljMGG4Q+aL3lzb8MYuOKk4617XC1cvtiuZg1V23lz
EGKkMSVbd0yhvNj/jx8skb8EICxTJqb5tOYeN/3RmxINjhdTgkn31kiOg23Q7p+VW2OgVQrYq1tS
SqlI7NFCsdevYMbPqd6cnUrRevah2dxPW542DC6KT8EXvVzDlykn/7JcKC0xOT+1gjZP6Iz2JVtG
BcBL2pp8X7by1rNjTKqHRXiD90IW+JA18mDaKCHS/bGuWnth+cY01CmduUyiI2VfZuQozqlEUuJO
lQ0epobcSklSmWbTgGy9DHVmFthZklgW1PT8QGvqqp822PxQ89m3msU70GE2/Eq2eJL/jT39mJ9N
q2NSF8qWlnMaQff71VZDAxbHmAmK0uinDLtsTqveKDLPUjWWvdl9x3zf8ePP0fp4CVqrLHo8igeF
u6dG87u8+coS4kPaRUPiKQJ6vxWrw6yUHbt64TxiZUitZxhJ2Qycw1K117eqZbWtPYHPQPiFOBoJ
jur8/sFB71L/78ocu0PqlfV7upt9OqvgjRcEjNnyCIm8CkkuS7vFGWaK2VTIhuhbHokKSWKGNxJf
bTYXGiZ/Z9xeBSNI3DgW8yFop8C8Ek54fXN1c2fbpupnZCauuU2Vd79UOBjDw1oQYrWtoG1eIKt0
uOHi5ZnoAWyg5yOsIBNf+1aY/ZTKjN/yI+MlIL5Cr+HsGdgeTYXKZJJA3nhv2dpcIia6pIUhO1wo
h+AmSNE12KTHino1eBOqhly4GYeVcBm/kAyEECDDg2P1jer+sJe9MUgxzTxEoi0wmCqNaPgY1y2s
YxuSrcK4D6X4RYO6B21LTW6fjaZU5t7n5wnSuCrbnbBpn818E0eVwDce7l5QRZqw5ly8p/TniBmb
Is+SIpLeuMUOdsPZJUxR+OezD11PjL3PiadBhvUuHp45ossvcFBmvvrOcfYrWCM6xoi/+h2gol8K
jz2qgTbANASViGODqNFUtmyk2tv00zYEWV25zJRsdQy+z/bwWUMQnURMREDhPAUo7xSIKFX079jG
q1W0FgP93aJwczrH1J1LuzGEpHuk9iJtxOu60XAu9RVOB1a02Z/ULQylxwbrKgVOLDqAq4/wCors
qvtPZTK2uxJE3kj16A3vSH6lE41j/ekgCpMTuuLeD8Ez3ETEgKsEQ+WfYLDCWXH0Or5n773qLFXa
RWsIIzXOHJr0oVnEYiR9OT9D53bjn36G21zUBlvJ5eJtB0z5/1i3L9c0Dj7eT2G6rQ2fg6iBfTAY
4I2ksatRzwNHsrnKuFVlIzx+22ypsRs/nkXmkj3C8ja4YIMModi76A+2aTkdsV9ST8lYnCWgzoCh
X4Luh6XD4Q7iehTdWi0MS7+NDPYPT5Y9dGDhCFH2OyBuUZTisGE2vfSwJTeJh+9GPhjSZKrlGQed
VQAk+HdZAEkK5xptfHOpkb+6nueYCavf42q4Hxkl6PU77tp4/kV/it4r9Y9I5Ney2H5ReINn3sza
lG/J63PXl1NzSsLUxAY3oqNK7EqbJTjIR/oNBxe0PINcYT6Ax8Y+s0y2fVTdqCNFZypcj98wkidy
WH5TEQDmGFEF9V47XtFwF6vS6/a9y3uKR085XPXOq+Qz7RPQHxQbJidaAbhP5Y38VpTpeTTcrw0m
kddCDN8HU8T3UBJlAvUK6h/GmxlhBESPt9jxdvJtVO3/LTXqsJRITbyRJiDYnXH8/K6yROeZ0M42
xwIaEUo8k92j58vAvJXEt9IAAGAdVg0to9n2BbdzNlM25u10//9RRNCZEV6i33ze1ludwW9MGF/w
XX7ptyHOMxaHjxgZ3YPW0trJuHwY3bnZK24MrqJYIODxdJByMqQwBgCytmWXccZWGkFrt+fs94KI
o4V1KAwTijFGdSBkwP963mk9K4Mba65GuZbYZIH2WMOHI9nqwzEOLRewlhnUxesDdLEDh/anjEVD
X+vDY0if0FRuamOqknys3mxUafeaNOhToA2ChZDExY7sTpT1/pYCWLwmE+CcLAUdPuIZPvxJzigM
jcNLWXUq4VgItZbFOkXD7fZFFcYTVbTO4DIdDD7q/7p/hATANXLHgtbvBYs1hokg2w90xCVtfxaf
U7H7/ONTVUCEbIflfgfnSrDbDSWzh256gUS1lvd6LghWU47ZQqxbEsTlrw13H2gz9TyskJ3JliLA
30hid4/dKl7cGBX0Dbgz4tXYthW4X27gncAbynmjqPqDW19il7JMesudreCzc1yEeLRg3RXTdoVP
RWu2bGudfz5xgef9C3ZD5ujJCB53vC0Ov9boHwmVgNalDzj0A4gmUW1mwH8GkWrM/oaOKKN5xlYS
Z8k+nnruo6rlWFzAYYuLjVRpzqURUgZgIHhn9vaHsjYTYu9+kT+zfXYRbmNnuYQ0gfotyqNLk2Av
LZKiQ9XfCQqPqGiA9Ro9TYgQ8U7giCWMUqjcJ0C92C73BOM8C3fE60moottsYDF6ct/Xh1JwwK69
sUqL2spPV/vE0mMudZJwo5rjPm0yX0xq7b1/B61ZjArTXWQg9/xTT+RPQ3I6vKWq2DS3dBdACRVo
5IdQslRZIOKqrpeglBNlIRprULrqknqwlTwcjcg7rkjav2YCczkV3wW4jDXXyTqg1evLYJFIDhQw
7Nqf1gg1BsD3Av8c9Yp6XnQB/a6QtzMAYsbXQG//JKHHoZ2J2ibrMYevcu5BZoYLwNJSWsYI9hGz
CeK728eFETKtAmljxDZe68eRAtdvis+F+fkCNJHsd7Ii0cAufZ4Q2LELvXQ6uzxoZyLblifOuE3X
BJ0aixz5hIqeZihb7GPD0+XwQMPsAU9lJ+7DxWfVLyWlPEJ0KseO8KrbOoZ8CoB93tUBevJJeBvY
lCUoiffKRmDDXoF+k87Yqva0RXc5Lm1RUlWiaxY9DZfHyctNWoodEFzhYyK3ZK+6RIV+m2fIT4nr
zlMqJEEQkGR5W8N25bkCXz1Jy2+p49wR2FUZzjhp0p8CW7JDho58izI4GirXeCv8a0j44Xr0bzkU
ImyJfyybRXb26/XQL4WagJdLIj1bzqhFvRYoJJ/tE04GFHU31q5w5h2zSiSyiogvGct0CKc6Do0j
EGsuMxAwFRJIUFYTgukInqbNy6OccbArVaJqjekv2kAXUAZDNvCVOUhNdgNzwhOb9+LWpsrPzzK9
t+ovHck/9PQFIzVo3LEdG3oApBvNmXCdoQggu4XJbrA38tcAzSwoKLb4K9CtKEKrHKsVi7KvzHTM
36W0uBhDcCnlt+MdqYx6lpegSRCLRtuWLBOOuagoGgt37krcD7xiYG6C9pEIzDS6VQmpYOW54eQy
iA9YU2SqL0SJOLRFVs/SrRg5pqQhq556cqqBZFvsJ4POZtlUMzInXf3zpGcoPjKEwK6HXfekhejK
QWoBPj2ARhSUOVWGAuA9kqZFfKL0sCg+T+MkwFFNAclP8empYtHjHORr8tO6ZWm85NNSUR2YPjS+
nJH6bfleUJvE6xLFCdUyYJpJkM1gaVLJypPkWJMfImYa2q0ExduKkWbOTT9rl9suxP9CAxehamkx
gwqjso4N0IAZtITGUWHX+aNCue+VkWm8N4wgfaX5c8lRDUYl/kXV7seoIuapjMXtSBFFJa0q9ny8
V3trXVQOUQi8byNHHDFJJFt6cp+ym9gINRYwXcU9tXlXmBnMAfad/uJEpMTkVOLqHUNOAzUOO1QK
tyfbc1CSNa1+183ogId+QpBUdTbCvfuH7zYn2V9IBvhIYTf0m5lwRUK8VPeNffKJ7Om9OUnUSNyS
EWjDlaHhbiojQfrsoH0TF8WVRADm6sh0O4Ghh30xRFim3bC+5mHsvgZ9V2iWf1VhEQsFtvw/Ir9h
0ebqb9wFyFUiZYcOFk+cBoH8AoydWx2DLbrQ2084T/s0sJtaHRjOuBFZaVTHXUoH5BOjkhuSxJGs
VLuBLvYtR/VoE+VCUCUbTVBVKEmxJYNsRD/QA4jnnmbiFd/XLEblKnWiuOtIOPc+RqWPgFSEaXFu
/iFbgq/I1/PLcXqGJ7l0oRWOKNe2jY8wUV1L+PIwG6Rcmxt9Cdk92+R4LMvKoQl9RPYmK5rsl20M
FPVZB2nvqb/PDOM8EBB8zX2RgZ/2RaoXE7aPaVgIlROfVKwZthkCOfQu+ULeoiUiOZdr2JbgdZ5g
njXSTivEPIoI2zYZpUXRasa7aEmmRsvFQc4AHApqZIizGHtyFDZgLw5g3L59bUXnjtz+s65kBaAQ
8plO8ko8a2q8cKqAv1OiqQZ/isVpH/QCUbOY04oAOTudpcP5exKLwAIJw+Ea/WlRQP8/bTeUmpS7
vMFL9Iq0omM3Tq7Lhw2QI0UfzyGpbzPNGmlQwLKvG0Mb6+hQcT+mbYs19oUo0GG+Ol76GyJStG6E
WDsBMb9PuR0PwiJzVzvo8RnbzAlJ0XYWVGtiTL3u0esuOen+dtP06xzeB+jvz2mDQ13gcGMmDwPt
C6XatAjM+K+/beupOmF4jdZDPCf7U+gf8MGqOreVjVO7zV+u5iPDwEkreYfcod7c2cnUKOmVKF8L
/Yy64IZ1//unrOjq8QvIPa/NH3W7+Q7E/KZrAsn1qFa+qkgwqFqhIzdSW95EprRz5chZK73OzorM
BMWbYzdUw5F8qlHTl/8Hp/dYToUtZi6GQzBTIEvspw3M1L8pu7ewmKwA5iUda/kv474PXGNUEGfJ
bEkiab8PjmCbMlxdJ6UgSOuuyFRMtg9+CV1aaDIp7T1+mQYml98LYU7NQ1/H2v3HvoADzjOjLRb5
BTcW+hLix25CcuIVRl/Tx/17MX3cfyDsHcUxH42rnUhnvxU2EPv2FP08WRs0md5Sa+8sauAvfymP
bN5bkxgrgrRJtxTi3sVbG9z43nJ/JBp5NsK0kdIUaf93g7PTDxLzMVvjBVK7dv57dZl9bZVAZxor
tYFGFBAmQQOaLxz/48H/Prczxz2JMoG+Omvqp0iumfoB7/fyKppQzS/E5N39KfRwgotudmF/EsRQ
D5EG3/9iKGtPJA541IntmzlNUt5ti7KOVbCXs0rOP28UygNVzhFNhpqqP9swZsRg6tZvyBz8+ZPF
EYt6QSAr2y0sz2MLSlUfYramZFnbgUPjs3zDfnvHjZarXuqgSCrZe2Uemqc1hhTW6XT/XixUbo/X
gAg3TSwATMV2ajBb5eAjrzxmAAMy3R41lgC70WmaNYfxrc4JL2ojrvD9ZRi5YjUgtyNRNw3Oh3GL
khV9D4wFK9VhQ40X2eUyJGJ3uPRdsAkyDnuOs7RQW6kMKVm0fQEcBrXb2iXUwmMLjUXZtrRYOzhf
8bGO+sl2A+tEoeqsEHqWy8Gfsnw8QsmaKzeFT9d8KmTnxCQMF+h6RnQyXQ9adHGf0MDNBOYWmiiR
KFhnhDCDODjtt3N2qg28aKlm7/aJA9u7ZAZfJ3P9AXc0Vk0Kb2+FmwpBr3zwfaB3UCGaih6k5Rya
izX9ZyMO5F7pHmSLTOWmKvxyy1a8hRdBWFQUxOlJgL2eyUovH4AbpZ837w9AI1qht8VpX4x6bdQI
8TzgEfAM2uYkc2BczlQ+2ydDCTLqPtDT9RDQiIeoAK2mFAW/xLzFdXTHB1619U8EfJ5Svbtt4jSw
cnZ6I8JsIN8rsAjo/9XwaevG6kgV5KrbJQVQix3BdyNpoc90w8Fd+5vMsD10KWtczgpEnRwmjdpP
P8AsZLkirlh4I1HhYHmWu0Jk9AvCwP1GQk+a2pRVo5bhDXgEY6D/dbV0AyHdaxODp/tfIGA4xScH
MaG5C7kx++bbJezmtjD13P10Ufli0ETy4qYHZyXJrXP2pmciH+q+aD3uu10sLPr+yKR5PbnLeYPf
G41l+pfUtBjvTD4/CVUKgFW5qutB3ZR63N5PaHkIXBOPnknCpjBQvX0FoLRF3jKVP5/YhUCtGCSx
sPOeUFJLjWHkf0/NnPhcTka5H8UMHTGPjBZBlft1PhtK7yaErCTO+MnIlJZ/uhHWWPhCMx70TkLH
kRGdAvy5WWJx63r3nKmH17EewAqztmZTzNr9E8zC7/ARAFndmct9Pzl8GMaWUiIVlpBWyb1Ao7ZM
IUBXSsGjeZWh0X6VMwVHKdGehIGnGiKiXQuD4OqAuiL5IUuzqf3XC+/maT9Dzt+BQJl2SRkZG/wO
q0SvOSPe8bk+8PTMeEysr7CqwX/d7ubnBhIal20N9ClNZu1vAK+syRMuenhW6V00zZZwLBkGOnrP
uq+opzakcbCaTjTANSWW78YpmuFaoJE0iKmHjgglEDbnJ5dkK7qn1REVkrWLfSRinmxOLLC0DlM6
+igWZfzDRKCIhaj72wM5ZFR4Ad1Dt2SapqwWNT0FTgl2T5KoprXNeKCiliDhpvfp/s+ctTWzex4s
3zlXe80dxPiYUsFnFKVyKxjjK+zgXcWK8LUNEgVUtUj1OQOGxW3tSZMmueuXVYNsR1hWez0+YrOq
PyPPEW8FrJ/mC6sG3LE6mHyabJnAJ9eA+eKAxw+MTyIJSX+wTF3FeeVQ3dSYlAaxYtwpEmm66BDN
oISYAkWnVP87MvyslLAMX/j7m+id5QhpINvXTizEMC+wcJ1N8Jpk6W4I1wuPN1Zqe2X7bEqI4DEh
uZVopn3eODN6BnW6OrcjkYxjoqWH71LNJmeeJoRDr1e6Pw9voiL6UD9YTQeJ3WCOvtOcNftfKMpj
lOt0L9Vg3BiCiY4gNDwxRPR7yBJ5qaeFG0yNiYt521eOlDRRz4YqmKOfuu4bxO5H/wQYn993/cg8
gx2XtjrNQSLSGGNE/43yvSYFiICT3yfaP+BOcuUOSYADONMfFTs2gmcjYLEcJ1x4Hw+ayomgo/QJ
/EeJB694FycR7XVurdxISOpThsLE2s+Z4G09fQvNLTq40Khavo9IVdWTMWlhdH8ViyoUxq8Sg7V5
NIiEZ2vyoO8S85VEPB5o2hz7vMAMJPa2z0jU0+ojT0cH2iZbT1gIYtOYilIWjRYC1qWF77vK1ETU
aQXIxVg11iQU+jvMkwql0IUXNTScfCxKMhdkPfXbcKZub66B09SCqncvbxgRK8O/F68YoYMQqvpI
y8nvuIOdy7TQ0tD4K8LFOWoopxIjEan1HKAD0OSRbKBdb0o5hTTNRqWyz8t0Th6z37+3vkAIFEQ3
ZvJn/v0Xv3nv51aDvcvxnjyN1HNWk13+42trOa+KLTnrg7qgjmVtdEajZScrgBIWFiOOn3PRvRCK
BOXM6wKjIAhichX0PqtpU336TAvyFQROxoIJ9+VwxSgJappjGliVfLPDVpWWOcmrFm6Pefs6f+Hi
4ek/9ftJfp4Q9mTZHuM1IfprrHx0T9RvTNbDsH6SXql5sAr57tjnB53TafH17RLOTAxviXvuWxwr
K/tbzI0PsnpxFSt4GHDIOWVqkuYIl5ykjXiL2ze6bBo9Evnx6yXG+Sm/q9ZYq8/Tjq3ghvPeX/b3
9o1DmvMQZGIecwqOfcarP/bk2HkiigG9BCajVDXM01iI4US8vC0hssQYKk3Oic+Gsd0S63MjJSk0
6Iz87UeYIu1LZKueKC937LiAkY2wReB9q8uFHeGADNTLfUzZNxPC/abMth9sY2yrndNk8T1TA140
6S3nPMi6UT/lfsgEu9yhVnyt5LsHHIRX/Rz2NAG6w4HG4mWpaYakdqyFc2X776spAuSmq0CF5HWX
9a9g+o3V2yX4lIm8YXlgg17EkjH6rby6860xfHKVG0g63xB55id0Oxwc887P7pPadLgAK4vB8O5K
a3GasWGQ41Hhss4o5pROnGxRoAuZ4a+kdIoQiogWBXKIMU7Q0DR9wnwHduo3XjDt/hjaWjia4yqn
3aaWytqkakQ+Z6WrBgIpcOySeudvl+tEJsEX5U0Ew0+S1V5QXJfH+3gDvz+b+Ge6fOJ75o55qfyy
jCkupiiWPJZLS4QtNoYcKPo7w//B7wSWvRqHz8a+S5Mj3RO5y9O/LTskdgHeZrd4dOfz+pgUfjon
NUD1UZNG58tYKLc+Y15WAGwMeS/VHZWMYMt9sNqcQTm1MP1vvCBY1AWKnq2FwDh11NvasdfYwM3W
p8GY0Hz0olR98z7NI82y0HG0oJf9Zb+0kODiuseBvQiqLdrI0Icz2ri9XaFu8gvf0XZATjm55pk4
N5WCHmR1zAKGg7mKJrNLj2GQ843sQU54zYoNYU4olAk//NH/wQpqMWTeRJW/g8n6O0A17l3XxsB+
iCJWl02QcalX12pNwApp+8JNFfqfJ2WiD4vPjexXWRWil1gNg/rPWolHUYx9YSkkNtPSOgIHsO7F
u+WpkeeNYSknH1/2X4T/X+XGOmU/6KnWcUf8VdorFEwYBHtNbfyQMVxUmkIDHfE/E1w0YbtaPAyZ
ExXdJIitEBL7LUTTjUXt4T6yczQV0x52zVwryG/Y/3OR/ffzgngHshaOz0XvXNR3MniqpWlhKDL/
gBpL3qQiliX8UNfQEUMcRFsOKPyqrWf5N7xPClPY0mfgdMcMaauuPY49p3zqfBYtx0YezR7nE/JC
5MT2I8iRxiSpXHANU7c5j08wFGKUl1WvK1Hw5v2LjVA7qzSrv8XzcDH/iCJjUIexG0gSAMOQyQja
J2SY83EyBIa2x1TXC1Sg/Qz306m7E1FlZIoKV9tDjoATOjsYjcDRUP3By7/WKfRCF22/79s0pKIN
fqdmArzkxhAwfhb1TUPoDjOA4U3kWe3Gt/isck1s+Rnijv5ALAYu14mtUfcVr9ee2ptZhrM0RBKQ
nfwehIPQioJGqmUozcnMNCjPBSc+evmJkVIQ4vDk/HUsAb3iZVbDLPQNmIOPoNz7J/cDbfb6n38B
dpQBAonhgvt8vA/wkgLt2m/W4trhNUjaLOzGE0isbVll2y7yMYfhwWGVJFyye3uE14/rM9+5Bfo+
SpLBn/D/ETYTOOOIYqJ2GZMv2/QwFi6+2WiKbWDG7UPdozEgf9ZQO0570bqJJwApZgnC4FyMDnzq
AKtMG9ic1U/orwOWZLbaXcEGcOLpiRVgz864HLmSuqDpgZ0eSA9sgEyepxe6ZExq9TND2LM9p5FN
G3FvMQRj2hZAzLOXn83O2PO1Z7bh5mmDp9EXcEJz/AtDSrIn2wQHegorUxtBNyDbizFOswp/dDQi
QlkKVJMqQfYM/CnWZqTwEqrowf5U+DCTDwUXAFAn9kQLggPapyqU8yv+AN+5b8DXAg2tvYi6lIEA
yxH0doeFLjjjdV3CauhuJLZ1RNl0yx2T5cpoQMAVjJlLK394B13gkjQVRUagsdluU/5X7lV8qMZT
dCSXrk53N44UMXUYC45oUo01JT0Ms0OHbl0Fpl2BR2acrfbK3GLkBDKLcQqFf+JCCEcr4TSYWLK7
lkM3irniKf0GdoTmtMp5WZlmOpJJnAhRtM+34KDYaFQ2DwJCfjU8e91zfPRL7CDNfB4Fz5GEFHAz
ee1br5ifEDGa6kncLrYkTSWBKBwgG/4USydVk+FSY2Yik3iy5yQKmSpuvDtaeNBv6ZDibFtG7MHH
6iLOxxN8VF5pohe0KEuqYN58DSMVQtj8yOMLwc/4E0/KFElJcG6adopV6M0xxlhr56u2HOajld/X
AsaoJqTBGSnqt3eeZxSC04QFf7UjqvnpYxBXxOONu0LAlfg0H23ZWZS2WjUYjddwLptGR+bKB3zk
ZRUUZ80J/6Gq2wdH8NebDSdvU21FY9zWHQobKLBFHhnTVEA2DkdBmeNhZVVC/0M7uLe/X//62OZ7
pICJzhQNNrF3RW4C71ctS3Fm9mEBtPRq9Afvv/Wr0eiDI6FfHB8ZrRCRYYrWz4TK355QrfFM4i2l
GaKn+9gkanpxlumbq3OHzpy/FW1iuke8775Ttsm9DEfclUYSMMS1sPT5sNHi7ksbu/3YpQXqjUJA
UySlGx1ljMO+6kL0XpEC3HHjfqbhOb+RADhWxy/DUDAbEoKNARq5xXTWJfVOlJxI2EbDBSiJFIhB
iLT9jInkx00kWKUD1lFuCH+anSzerD2mjB70npX1YxVQRRNmybkWILckb2lP15lzQ79t31+Q9y6E
c8lUw3UtIGUmZ6mjqNIj4d89RuJAuHDIWFSgYkasF4mxi5Nv3xWj68RRJdj2wb87AMF8JXLDgi75
4iCw7iQ6XJ8ed5Obup3tner/C7F9ttc7MKpTVJLJ3ZUpzxQh7acRgzcHWM2LBIacFsuOhEkIZJAS
kKzDti23FlLlfP3upBrFuGZCd8XNk5f78ZgyUOAcobSrB53N6XtU9X3EthxizP1TKlfVNRAcQtAV
zJSXMnHIoaXZnj0zQgOuaJ9esVSq/zdtVWGt4V0FAJkr32gKs0vwaumwFnELKqKyFpu2cxaoPV8C
Ei0At0yg+7BVGdfyYG4/mjxa/r7s+uBg89RU3Pp+IpVEN1rXXewIgy42/77N6GOG1UryrSXZ34ns
vxULTUj0PiJjj6KhLz8HHr3oyNDpCKTj1/9hnj+aRfqmTyaUHFdkCv9E9YheQKd50xbABrr41Tb1
qLgkbTgQ1VKQXkfKWsyBLOXnwdWIgw87Vi2Hq5G/UOsdP9fdphMCz9Xu1ZyMJMT9Crk1CSEec80u
DdajwYpHEWjjBiUa4bXxpqhbSHnweCKgo3doLCsdkbAraHJIFAqtIEa7Tb1C5l+Q2jSJyA4FSDiA
zSpLRZFgHbiidwkOEkGiSZvM1QfapqP+CUwOx3OqPB8gFejJO3a+sVtSv09qvjvksH9dtWMVrTqI
r/ctVtogQIW/Uw/GRx6Lij5MOCMk0IuVzQuJgaGJX1FAVMSsKLnfToua2CfApsP53aPkq8cclAjJ
N8VupfdOlt2DryqaNt1Zo9UK3Xsg3aHvXmdNgr6cWaj2IwOD5G0fZY3fGO4xU9kmISXVJlbt+b3D
CNyOF3rJUq1TL0g3kNJza5WmM9t6GcUU+XtLNlMT41YkYPTyLELNxrUbo6/Huq1c0xl/6KQlqvsx
jPbmT2ts/1ygemyOrYySehIlRN7UyZZEqrAMFYCR3+tPbJeKy6cM0D6/uYM3GRkeIVZ0tsiVifQf
2vID48g9Unmf/bOMpAy0BOb8skJcFB8hYIHW/o00EFGPt6fMfja8zOwQd6XCBzasNZ87752O8Xdq
PnUZZiwJT6PlU2aP3cGq6SzH51QwFGded0kQ1UtnKTTe68qoUATuCpfvy9NM34aoV4Osf27jdOy/
VdMy+zM5qiEx9pNucpIIqVLIkM9tpjJQSdEyGQcL7W59kYxHTR8ddpIwVtPWSS+q77w95gaR8R7D
uQVbSzBQsya3wt3TKjbNrtrvwguvHq2Xbf7MlMd8Ql0DMu4ELXY22w9K/Y17B0bB8efB3NomeVTN
LH4jz9TLHEBBhZqtq5nzNSmalluCknZc+J6aIeBk5AL/wgr8iM7yG9sOLId+3RvFp3HNWflnSgo3
XumlGm/BANbLX/9PoQgBe6brSqgdXE7WuPjxauv4kz6lW6i/8SAIZQBNpRKCv8nCL4sqkQxppFDZ
mtC+TExPyuPrbeYmLu7tYGYjick99mQnkEwj68m0e8ABkWvZzcg7qrfNbRuXKa0t6GzyY5rQnof6
MCQLLiROiPsuEfL8/foNvPROKETwDdTgL+p87O2aIfjWj+c9avtOBhkqvV/v1eYzToRooQLaXHFY
MSZgg7EljVwJFZg2O9rKhGPuDkVK8tRH97eLy7VqZaXfGkbqVVmXD9+vzxh7ymfubMuTnCAHaCbh
WH88s+OHFk/4yoWQyKcT5tnNwEiN83LC7/dRb4VkBTAg5MfOTQdp5CjjRmSGjm3hL2v8aUyzq6UD
G+CKVZ/OjWAKNrsPjP4E+ALiJSPtoeB07nnVTTiaDrTFJMHfIOZAlz1NdPplphEvJbGNKSufok4C
N7ATQgfrnKzljAmBm0ySLnRkqUnvtuItEQ3ZTFoh2nBNsOk3WgHp87y5mlM50pO+LcrFkp+Woum+
5a/PoxedjNq4PIACFaLDH/mzD+C5JMa8mv9AjsC3+wU3+pfcXWFHi1SCZmlgOKpu4xBa72XqKxZL
gs0vl9dz2H/we+H2DBC2Frmg4lFpyQmkOIubb/bJiZ7O04NTnZefFySCelcKZbZyPJ7MMJtHPjdy
c96dcTgI/4oQmygoRFkF0TD1mQ6eA7p2DZeaMIfW6L+jrOKSXTKeAs9Qu5naWFmm//tu2OGIfPk4
9ewA4vhougBolAWi9p9SLCuy9fs+hFG3GlMZx19AJa4zxxacEMzKMTrzCWDGFJnZWzutunU+mzMu
WbmVKHFek+nLY5oLcqzkSMbif8fGZMcZxedWzs2XoUQV9jlLgfr7G8oi6NRzZVO/Et4n3xk3kMoQ
faHYQb6/D4Bm0f1Xgv04ZTUT/lk5Ng0XA0aEh41kgZuW7/cAGGhNam31jtdPfsMZqboToQIJL2u+
q9kCoSS+UtVQbhdl9d9Rm+uoqq9TUqUwuCn6FCVANQcvkkKeWenv3/JW6Z6zC0JZyRQbqzEzSP+5
rneVk8VoMKRp1xJmOyHj2UwkKqsa0vmGvnri1c98xXY59728n5D9OL1yBSFdtr2P86RwNMBmA+pW
yBdU6vLHrtl19ioLnTuXbTwqOMYNMf7181lR3Qkm5h+YetShFFIee6/ptFQ1ZKHlCpeLqAZo3u7/
wDiuo2i+wNQCzUG7bZqHG/Ww9CcfrR4mSIQpamE5UMveSRvnnTmKefDkaXr3q56uUJaJG2JAfZ5z
gKBgZOe/CzAb+Flqb9z8sJ68687p49kOMXWVVAllH0DJsWjQVkqMTrmsN5V/wubE8Ie/cgA5EReE
s4iSqlaW76osh4BSrVWqY7HKibYfBpfBuPCoy2SQlL73SP5TwLywZyvAVN1XiVxqsBHrUaVTJRPY
c3Q/i8m69KxWkClARhvv3Idz+xBrljn2zrbBXkynUkOExXuzYM/+4hBG/yCCYJ/k48q/qURNAKB3
fh2FK0cjCYhosvwGmfFNId/gwRCzG1lt2MHXqinuk0lpG/eWwZFF7+91LfbE0/xMYgniXHjn9orr
QYO/XzjHStrFLZ+5wTaXkXX/fqzl6gLIp1yvZ+t6wQNoZuxkMqUVFcnAC39SJKlqjoeraXr5wEO4
4BSWZecQP3P/48KfmGP99o7X09aSr7/7XamYkLqdksTA7P9/7Q+ZVMempwDjhYLucvZW8/92vhV1
Rvxa18KtIqwhKzC1yvb6PuesbVR54Uc/ZiUbn7SO+QLMFXaaPHGDiD5QeAiTUo40XOjjzn7cezaX
ElVm0LMC8G7/lkYJAgRIs3AI4spsjkiiNiPI4oW4zAwWYD3nWUht5CLzu2FqL2rPUKPCsWuWzqSo
TTfPIv61LFjRS0bdqBIWTCm2jdspx3tKD9R24rol3olNzUYbmnI5mvajXbJs2k47oVeQOYUxKzBt
20u1auc3KdLlugJ7PetGXvwJcpuDwuNtt4IY50Qxw1xHFnh4nJ+H3NdSIxQRBMN+4T/H7B6EyNDj
U++JU6ZQQWgaF22pIHeoPjDrXMu73O3z3yo5y8zOHDcQ1kIY1YpjGhQq0albbXuYFvDRi7jmS9/j
QylcazVhgns1tcDlBRJdlFpRvi1pDmxKmNkydy+W1IGQxpK/hvj+cGoJe2OQbzLSK7D8z/+3WrdF
8GjO3S1ktjpVFGtJAQQR4ok8f6HZAP370bAsyTfZZwHbNd+ZWzaPoWgu4G1B5waLUu8HX3y/dkzo
iT/Zzyz1lqTapZZF31oKJMSlSREUW2I5Hrg3AcFvQHG24qMz333sJpqMCDLY15J5H18YxF+LDW4p
tIsVWMDZKxMqcBLBMFiPDqgGooJWJBDSvN8dSoBhfjqJqiXyT5XYedep5AFEPTkzYMt7qCz7TtVI
cXqdlMdsFxzf0PfeOiocw6gBWuq/aF7nnrt1s3OHLeSDI0i7jlMfM+3MUSSa0Yq1xRclViI5a+qp
E+DOuX1eEDifYs19Ky4lETG50GwnBBAyUbdvQIVDjQEJtSMa34LiUW4Ox/tEDDWeP8h/bde/sV/h
NKJpJ77kHcw23qzAGSdh3VRn5ygDHNagHRTVjKiOryMzDrCoAwwh1UVYH6w8uDeMe31lrY/RkHQ2
Za0tIqtd6DpNkbco0u5AQMW9mNRLRbq8KrXVYBEaLYM1HUvdeW6m87z5+kzH1ZHEyaK2f0c430xw
fLEGPqRuOrKga7Z6Sk+F6TANqr/9eBjhnlEOKYiWKngVVCjunb03tB1juDhKTFo/OIEDvHHMnqU2
VnLWRuVX4DkPTr4ckkdrdP2kWQHs066rm9182+r6AfdPo3CrGfAVmXE+EFoPStm8wYelGAGwdcYs
qSN1fhAptZ1dl+kj6Lhgxkgttebt4ym78/bQHIeUKLgaGfa1TVq9LENesIgAPYaw9YlAwkgAFSs9
wQlW2muQwdgncqUZ7MS2f6QJDTQHKXHOMjahgdmwYx8XckTDq/6rZL+U7Pg2gz+w4HFOjJ8p3yfd
GWOhcK+4lg3UKzs7tT+wss0etY1X4FF1qhuY3Grwv2/9cshkIf1awOvlARt71SIptMa2nPeoMJ0p
Rh6FVmjNhODqluWEA6QVIX3OYg7I8FcabBYbVpczSzRETo/8juu74TMyGCcQKsinqbZn7bbbeRKG
TkUdtUFQamjvuolP/VVs5RqvLKl9PZZwZ26qIvaHwko2atHRhDwnAyW3e8ZmH0nRkdOZM4nREXeD
fLIPc6L+q39XrlRHDHbiGuXBssuNZnZNXUgQrWQzfm1ZoRBC+1ltvxrd9yGrRkaCM/AXVmse7YaQ
2D/SZs0DnSiC5OmbkAmItpf5P7qBq6A4jeX6PjnfaJU9MbvHOxvbgeOXYVJt0+ck7Zv1BHoy8bM5
MzjfERP7RM+37M7FbA79G25fIbFy1sc4+54sNol7FOqk+UUMoDzXmcsB+lhvi2XoHtFCEmmuY89x
M105TSYIt4hIVnLEF8zqel7Wj5jrKDuuh2Ba6uF85YEmwHfAq9BOvsFqEMUahIvDUEwtqI5oFgWJ
Svr3GIKnHyBhHxomm4a9SwyYKUE/Bhb7NtOA/3qY7OICJI7kjTVTU5K1iN2/frCUlpyG8fnNOWvx
FtfHnD8a4D1OBxw+rcLvFyu4/Fd0ongfKw96/CiCTg81QRw+1fL1Yc4Wpf2azN0dabPlL3n4YrL4
6swsMXfvxsnYV4juEUVMf78utkSX6hmB3ZyulgDKa2z1PjEI4NrB3wzLU63gkC8LdDs1ZzkOAklc
yY3NXiZAQa7/rbPH53v/QNGrIXn4TgqtO7vAAE1c36pwVaXJg1brdDb1rfCoWjTpqFxrp1XHUw91
2TU3tV1SpHEuR2iOfwHwx+xyvGY9m8yX2eIxK9GUn/vuvFkTVR+0UyT5+4bS/ezL8HTT3ZzvxBQN
xzdVSfK0vAxBr6SXfIrreoCEE7U3jVE9sUWadyI2SXKS62urtl1fHxY2FcFvZ1wD3txPCg30WTgJ
Ryw7ncGn90uiGkASdY5ZN4JX70Yk8GTVwahcZHL1nYa7//bFQTY24oha0KD1uMezNZHL8CO8M4Mi
96WYOrPsn2iqf8d1f5Lp4yZtMQapAz2fb9JSCOazR7l7I50vczdDdWeQdIEEz6VrdB2XnfECjN6D
LOucf8PPXswXfalQY1i7tamDsA249wGda68b0IXaC6084kGeVkDzRyL5M0RgpGg8/UFVYv8EvE43
MZG4nsTGdFiV/tVxWh3gJTtc4ndWMsEYtrKlESX57TjmppFMittU9jzn9dujLcC41ofbB5SbjvQK
irt+dakos5etJwzoVc3XpctY45ImGZVCAN5ZX9Y8qEm+dwfJRN/H6ZYCXMYGqcnzDpwBw28wo9DZ
+7ePUQwBCdcsx2aE7VissTY8YaLJijACKSotyKRbAGH7+421eXVQZSQvoAl+J5OKJ0C4YpFWoRjW
3Fo8hUDyrTLYsBsPm5l2HgGp8atqXx8sA2UrSyMWy3nbpdkfl1NPVA2mDdGFrrAGPFfT6qC1UOZ/
TsV2sIJJoT3tgk6KsHh/o7fyQAKrsvz7q01XXpMAlSz/1y8Rno+4NepbAPfD/+sQywtj9kcRxLu3
tjRu68wq/14ztp0nWW1/Jv9SKSGDXBqL4Qx5TqYDwfiTLOBHC84DDNHKGmjjmFL0aJnj7PeXRYa8
O/4h6UuMHNRlXcoV3xqxEOOnbFrgRP3zbf1JmRRH0xLefa26vrKbnojBQcq7OvtKXEB7gjRSYivB
GRx/zxtAQKtlHp3hb3624yi8GLlSKmNq8avwwZPw85seqEGmd7qsYcxf5AbBhoHhzy4QTewzcvR1
UFcOs5midMJik1c8A900kKvigYoMw7eHPkJ8cQLqsJlS0R42Du68f015E+FPqR481MjIr6+vUHUu
ctLw2lyHjUsymHuwPBUVbXXXBDrRT7b6PHglG8mq1aTAaEIAwhqWohdPOienNUcLsyi1A5CA8hCG
4B28Jsl+C/KebIqjLOc/tAS8tfhb4zLGYDM+Pvantmiom05D5OlZGAnoD0HBSSjO8Z0Kz/7rTGik
+ChIkHanSxA4KW1SuV4j572kyz98cRja0b8Q4O4Y6ZE93lU2flB2VAODSOe5J1OXDH1wtmawi3ik
EmriZCXvKWfHhT9fTpOLxXOwv1HxkxuB53NNegqfFBPdOAWDEYEQjG03VN05UEjI4sqYVAUjo2UN
NP0FweLgKJ1zbubYZNk6Ri1gGNy+JjThPXhRaEwwdbwNT50jTXS52XiowGV9QJXgbmcdWEWY5YFU
JKbqcH/4YTHapBAWZfuOSMaZJmEQGbwgcTdwBLSxbFggWZ5HI77jrfnPS1QT8EnbgWFVj1zkSlSo
189MhbNByCk5OJfpKtxaz//cQhtYLk+Vx+D33gXspQin/uiCOuZJKpub0xIR/bxz62JKKMe/uMWE
su22VhvN6l1J/vLgW6NOY25UIATDn2iZQR/bJpA8qvUa8XZL3cwU0M18zWXM6hdT7CkV6fxZRnGm
xu5f2rbtd3RwlfIGRjCZbsajT819NE/l+bX5x9ZcACw7noCu4UtpyDWGqWnmjtkD7BmMnDSzFGi7
f91NAZqLAc2sjp4vKXim0xghJPn8MDRoAKM049KoivS6VqeKIvrtYg1R3iyazW73LA4xA3jh3Gpe
jLGRC0dJIX8twjX5t3EpNtNagELdt5615m7N8VehfVXvnYfBHW5G8vfvIdBEGKVfVTxiwWZsRIQg
8V/2fgCuiQPcFJSc60V1HQElCgKxOhpX5cMo/p+gIbOXhY9GSFjIKtPGwFGJFR8JBWD3lzDcLEHs
o/qswkFs5k/Ce48HewtMkxQEr2/tIet910yNhvGBkLqJ2WuzEguPl/rREOZoQsax4zpWTVPHHZsU
MXqHHQywRd6E2aXzsnHx2R40TfmAjx8U/Bl/+BU/B+4pLruAWSFT/GW2MbbcfX3taKwykQFQm9RC
noXo0kFL/h/+fTV4OEqwUikeGm/LuUyH4YuLdjhSDzI9c0ldk3G3UVycLYWCIkoi1lMLwYXRu+9F
F+c45mMCRrF63RlZhymUlaxEv4vheKpD/RLdNy1QLmvbtQHi+VyC0CPgfHqXmAYrCeW6cByc/JyT
i4rtAIhgfrQreTtFthoRfE1FCtpD2M5Fj04BBGAv3nW90Xv4wzL0P9vcIWxL867mTYAA9sgdohqL
M2RuKzpxbgrwkgoS4q4agR+DAWPB3iHSSHt7fWKxGXno9YYJzxD3wdQOIgH2XrgCqmVIaffnyVr+
KXUK8QxlfOkW6gweDSUdP9yDm1Lh1l376kjHoqwYJEh6m6lH6zp2smOLAJF8XzIaknpS1/9N6mqo
KO65zI/bS3xE1GUkN6RRLoj0ro/U0zYPtd465mJDsfgazfkYEXdo0gLGj/ECvpWWM3dgNp68ksQY
kuk5KLMo8DeqVBLjpKGemi56rN/TMccV7pvGzsSqLTD+Z4jR8HTQVlmSw9V2qP9CCnATGyK1XaFC
Y+JcJdnR0NUR4c8Lcl2wRhlfCQZ7akatAnFIwv5TG6qE2T8uMq8auJnR3E7OQC3GF/UvTK6TFe/Z
o2/kv9bjF+w3XgWmHnTnv98nSHdw9gcC32V2LoWpV7lefzJCsBWu0eOVBM6A4JzwF9lxhp3W3EyT
JglnXyFtndvCeqdNHSR4tEimNLO0ijqYXzmSmASsm3/Q7TbvNH/W3Kt6MgTArWF6RZWQEUxff26S
lAD7VxdLwfssU6ht94tgTS+dYa8uSQrbZHh17W9EpEaodrU5kind0A+qkuH9+1+SRjwnch7POYXl
BoxMdPeajtXfy+s5cRcaeibFWl1Qffrd7lIaURMUuJgJrygjU/LwbQQpTl8cLvu1VkIZnJpgB0nD
Sl8O/lJBDtSSHHTRXeCUKwkmBkr2F7azVMS4og+mm2ACXxm0FeXjaeBwWGIQ3srcr18OnY0HPPRy
fs17fZMfnGbuMR17psi1FrdsYDMD5J6KW6JZk/VG5e/pdq5D+QtpvdwUIWt8GBz61U1BjXCyMiJa
uWt0b0o3gKYeCDJZL+T4jkGMX1wGtpmC9LQtnSfP9qFRG8mOx4CKQm5nFWEAAsfdW1ZXkWVsf+7l
g8R6NdYtlbI/tScQW6H3m/S9E/bjnt2m2VTovXU+CW4VEXkYvYo5SmYQccXT4gLlTNCqEXZAFReW
fIIO2mBlb2bctWdmYY0WQeIEqrskZekBxeVTvS8Vz1Lxu63qQDEhKbEkI0/NlV0fuJpSSUo4kspo
rCILJHpviBIdCkPCvC7PKrsIWQJKOfQudXe2RQHUWn8p+BU4PAkzEw7IXJkBUvOEhgcVXpL2ectH
WBUtky7y1iJccJioUH+6r2A0FgFEfRp7YJZKM6ZrH0kzjhD/MAiGqwy0XNQRrSjfL/6Ecu9ZjFsb
mc27bV3vj/HYeUCiaMLM/Q+czfiT4srKuJqSpnAHLWs4Z9vsTyjIL2bTRC11/zK845uAUEGyEZpr
AfgWkJba0i/pr/HvCfuuiqZ2cF0h2VAxgOWqH/MkC0wMqyarOh8Zkr3FCX9P/2VmBqr0jnSDLu1V
1LgO9H5/sVUN8ghPXs8F4ZpsvAWgKSwXwmNO0/D3LvSwvzdJonkaL8SqQ8ecBIdomQt1aFafE+Sn
WPZJEMP8jTEUKuPHZot1V9KM4ecu8TbGMqZfet8knm1LjbHxGx7VD0BhRIdu07E0bSf4fzye2XJ8
2c8Yibz8r7HnGi2FGqdqlmwTlAWEkFZqSU6wU4mzcsQBmOCCWO3yUubiuwTuGK2rfrTeXVgI/Q7B
7FAVUa/bG6RcBK9rHmMtt1FTJgMgtHjTtMM2us0T98StU4yFN7HKv/1uwpsjxOuNY6qk6AP69WbB
Hnbm/kA72eEmedZdomBaU+9fx9rzrfR6/beUVMxk3Re9eyKHqEFfyU/Bx03vhd3+fN8lF58/1qSK
WApQlIxGyyfwmBIDxZ9eMQGqF6EtCYSzy3MCQ/mCfDohP3ax4yhybJGF2NfFDDQJ87HvPYQUblhA
cwE4VScoo0cVk3hFRp4Nu6Oxpo5lr9aoWaXY/kqUEVX4iQrMb/nz2WOqTTPY8DzL883NgixTYVCs
MVjJHJ0u48HaX21Bx8g7NwKQgMCbbIQarHYC++MAfcWBOGjks8Qcveq1Aigamu53UrH07d1e6Jge
6UdnbLj/5zQjRGRIJJUIg58HdOrBL1B/Ej+gEZfOfXcjh5W2F+Xzazd21eDtWJBU0dXJxP83TTOZ
z/BB6ksglv7qzYWGf4tKwaexsCV6GawmVll0W2Lv8pQM1qJpmEZDrKEgUi1CeNh7Qp/NiNO7PyS3
Zq2N1268KBbIMO/n2sIUlv+fF3WlOjz+9fiNHasW7gwOsBtOMWZ3eT6DfpynPaIibHmjzW6k8Nlt
lKabDnKHSQCvF+p4lQzTmT77lqkpLCbDIWLNtAUrhH8bxjcNf1kYkSwpBGHwPdlA9mt++wqoKdsn
Vfk5XiUp32x0vfOC/jcZtYjX3R8lnFfE8b1jIg24nuMv21J7wkEVUDhxsvXECJJB8i1AUrGmh925
Zpy98Zw1wjaXaebYJv+PLhvyvqiZ+T04y+uw5lKPJU1Oyvdob9s8rxY9Dy/0wHfA+Mz0sq0iAyTN
xXaT1WKMgY1dyMvN7oCoVe6bpRaWLGlzA67AiQt0sjA9ouI+DEvdqKj0BZVBm/55UMSXIczEasJS
FzR9m5Y3OkCWT42ymM3r4bceNLcIx0yOt93BnJckYJmEuvU85CUPgq94z2i6EmK0EHUM9pCaOix6
fKWajhaQrXAuZ1QnUxKfR9cvtUqgnMGlfO7icSQSvvkjeRuG/M4IsmFBgZdWUqJo/5XiXdKs+Nbe
WM2LD2LxkWMawQPbwOAfSqQIhlQJTmfJAgPu0ooJg4fSeZ1zy40KpTk8svHneTwewqNRZ89NXp+z
LFMeV0xR/WJOVCoAgYYrf3S7gGnLpNB4OTsQciN4gHFeRFoh7CiY3iGbV8aTjzThOwsDrhiT4Pyk
UxROcBweoVMoXWP3HQ36VWy1q/JJURTFAXB5mQULhVuHbpcAGKiU9Cj5goz3yJuem9+CEEFvqzu+
0OMIGeGM9Jaa3kLsDEzIt8cY3sAoKMF+iKUAx5rPRe2qGYXZ636p80X74TAtDDxgjEG8p/3ztDw9
DqICoCQLRC9iGxn1E5y5ImmE4D1Jgkn+PYJr0YJQRcfcFppL4HRUWKL07XwpF9DWwUNvbJsjJuZu
pNEvvJ+oConoz46kC75S3EjTT1A6AbYqFeUupqpFzzQ3nPqVGDkBdiNs/xm1+q+gWUCzpxnqq+d2
XzzlhW4vcD6Gz6F1H2HRX2RLoS3Ot2DRz2n8Mh/+SOPNFyxLWyvGaVnMysT1/KqB23umC+05dqKS
prAaWrBCMNVLb8y0aWta3wKPRRxWWhdAIbLo/Zr1iBhrpgVB7foDkNteCeIK6zrQapbrXcC5Aj1f
YBwaZu4WbfUzhxvVesARJNe0DYjT1Q0IRCchPPJUeJkHMGRgVDuQM4MmxjqUR1zVWPwxvlJTTzmv
nZCvi8C5ATlH5aZCOSUm0oIzVnQSDbKtcCtWxkFe5WYooxBES/iHbOKZLxnXvIgMwdrXf3lb/0dM
5HkUPCrCqkE1zXDv5jXW5ae8wg0r6jA26M5KcICJmLPBJN2RH3wKo1ueZHlPvwQKBvQY6Vgi+0WM
dV9U9ZEox2XcPiMGEcTSwFJRbc7Ed2TY34xYjF0IjPnj+tYv+xJVrYILh8yJeQGsBf34YKtC3tBX
uDpxC6yRrro2I+pHTajy1SmoKBnJww0IEDdC8rxlOErDW+T3j1qHEd4C4yWKkf59i7bXh8t+jF5R
88f0AuzsagzG/HE80WUKjL92ZxWIeTg/3TdJm81YbrRwh8MRdtQRYnMG7nL0m4JEx2s6uUdAx++E
aY9gFuWc6xIxR9Yy08G3KsEhDP25wOFeV/ZDH9Ow4gKmFMb6qPW/BqY1QcEqDfVDMkirU2qprW5s
pUFYMhHXVOyIwVWLmYnDymo/CQUG03uQzzLzWU5Wybs4kfwIeBbpI/vQU4kGzmU1pgzZ9xg3XxBM
2s3uwUeyeb4VvYorxhaqXKGUp5Me6oqa6tYf75Qvi8b0j6Lj+Llr6Z44QsFq00G3fA/wWTloyr8S
Lr/pghOckSqQcH+F88V3DM74IhifmYZ/0+6PYQ2PYb20YlNIHIK0y2YN4dBN+D99iSV+/Tc8dv5M
BRR0TxPD6aEHFoi6xd/Uib1rEPG4Pxh3Dewki8gZThh7qpwhZWAoegZXLfFM4Z9wBcJUj1gjHGgJ
Gzx7vbNI9wwEOl8O0WWnq48L8cxFLOZHSCBPwPF6mIoGWaE7xd+WSXSxQe7gHB8qYGc3IafuwpPl
0UGXhVJBbvj3xFxRaJf5yNZEWlqH84/eUvdIH2syU7Pt3iQmNhajHnpeoNRUCJ/bJ33dHWYajaXh
pBTyOTnx6bggH2E4fFNsz7O9IrxRRFEPUpYFc9XGzccIDaGKd2qIyNxiGuoniA5U34wfcMul+AG6
o0qOq+QXT+2NTrXgx0bhxiX0eodP63HKn6V4R2U3S9kaUp0rPIZurIGOLwQKWTodK0BfJAqUVmFv
W5ZYEaGg710F0hAF4OmzRgYY1U5vLqbqlcyNGyOhX+U3u1QkhWDHolBV6rTlaoPhu0vJt0aB9cdL
CWGSYuxL17BaYbCvWuGQ8iFmObuGBY8LZhV6C014yNmOngsetqEFla7aYjbSGqVtqdjQ5Mz9OeCd
wuSVmVOhzPdpKUU8YuGEt80l5XWxkoUYyNsNjFtg1KLlDY3RlQg/R4tKtMxIew1WBh6QCtOo3nsY
zFrUvsbVU01ndlUPSyLS3JcLCxooizyQ7p+OqohHzlVSPaG7yuXYQOwfBfiNJWr/F/T5nhjygtry
BPgBcrTvkvuboqZsxfUO02abSJbFHyT9UcZGwh45JAhRJgKGmldHjU00D87wn/EBbO05r/kihLNf
+PrkzL4LxBNcfCSrqikXh4+LKbDn6NnaDIuigzJs0novo9ipLWmMLUQGJX4o9GAo5qMMQEYmJZjh
qtBSI9od5b354K3s1+CfPVCJ04mcNkQgW1eht5uDW0TbwfNyH75nBJA6krcbh00GW3d+ysBS7kN8
ruFo046e1NRAIJNNYnaqPPiZFwPZXGXo3uNC62PjZ04LODWVwW3NlpcLjaah967A4I+VGDgUw4Zb
VB1MbW+SBtAsCS5bCz95PDYBiVbg7hkH6KHwlA2Xyv5QAicQn4ARpqePSnj5UU8eb0tQI+db0XsT
9VHdIfsG2EWeXAGGuaXbd9/3bFNqE+1+oqmeiU8XG6ZiedP+ChcgDzJtEBDvaU6XUuPv+g8SuPlT
wgZ0IiXd3bf2JnQ2hnHvG4wU3oBrXHIZnX0m7w8PXvYTDSXB+CAAGuxhm/BsgVKqhIHNvsY3slDm
YBRfPwZjDC+Hm7nSn/vlBTkBf3JF7hYy7Lui7ZJq/eF+YDEvXBlc4d9CV89bPSv06CuMs6yEceSY
b9GcHFeg0fBvzK/KukspN8vUdGdvG4pCZ1M9nyHvW6WYxz9aV40WE3KFqgbXgacJ5E9PunGfcV1T
FXkK+4BHSuIW0i0VCE6peaxMuWAE9vVwQN5MZd0kYAE1Pe12nVk1GvmztuSYIsksCyTyty/8fKZW
txmRpUktYfGOib8/eXDTic+RhpmUwr8Ta5McUHYvlUOpv4Ut0A8P+RlIQNnkTlGfDviUbNF1isaX
cohn0f7E6kscz5GGJPLl9A5SrzyNc1hJQWJUYwQ8qaQIZfbLrXnixBs8DCAXjM8gNuU5cq8eYT3W
lFfZ8mofoZMNV5n70y/0oTmDXgMtb33OSctuOwPGTyN7LzHy4Do1EyC18WdbxjJZAzeanDEJulzF
12pH/VkEFs5BGxll4buuE7Ip8nmBtbgOfy73Ce7JEL+snT5VxKS/lCmLkGpnjeLmBpii2J21awn6
axqhsddfu1/TVhynpBTxTgS/Fy6uIHzs15iXZkTsETUjCAWEtcUnTMu67BMArhCpecYXcC0CL85w
aGCQfKvm8uWucN/bdNhl+iMcvFFgJyIgIfrxlYyrpbNNRvpTGuitTl1zS9NDb972Dv+m0JvEfWCW
iCi+r9jswxXpzgdbZfG1ZMpamSQyiOqMzckvu9o74up0pWsWL4nFgY87xDlxlvJficlXmaCvRmwl
E3j2Ne6B8k6dFyQsLRZzgIhm+5hM1lCCQH0jFWoIspmKaCVG0AuSZQoJEpwGB0nBfgNaPAkcqlsx
SJ5sFmhauzqrJHVNuCXO6qwRWOzg8euJmOkSBLS8nSyLfJDQsEr9Rq+SAKZEiSGRGB0J2rMtYO9S
lV2Qbd3RfVa21HbpfG7qC5uL9XFUPuiidI1bUSldzjUSzJrFu/Y1DhONV553fJODneU/+B1yf9aC
24325uhQqjqoQfYABBnQZNEdSYGoJ0T4U60EcValmVNCoNK3Wys6RuHhY17GGHw2PCEfiZjeaS/v
h8WvLYuaZcSTvgkwb2/yTBA+bECc3yJB5mK+IR+p9035NJL2uogBsGvgNq/ZHzDaHAubqS9Kv8Ln
sHzbdiBZQt2SIi/T66jTZpwW48ZP8wM30bwggYh8Q+J2d1p17ACrNDzprlsHoaGmWWkVNfetKMyu
LbTX0BVwJao6fNWSYLQqGVBo2dwrAy5wViVObWbr1xgISnDJjzu1xmdmKE0w2g/0VeWIgAqBOjS9
ogOyrrCl32upFCxHkOTgIfQ+kN1A6c009kGJcq3bp0ZUGL4vwjDbaFM5FaPtYy4Hswzp+SYKPQR0
pamhKJw6iaiQ5UxxogXph9tzVbh6zg5dwxzUscl1gfihsCrZjGPqUUJfwWunQo1VGpk/FnTpSqhQ
z/LgWL/HcGrruKkFeIu8Vi1pSqkRpEBM1gcr9rHA5InF25VoyO57prwuJxksbjzH/r6xDXI/MmKk
aWHnu1hhrWz0+Wqf2kDIbP2bsRIfX1Hdg7IZYr7f/sFjpy/iQ8g4DwSTQEdIlnpDnQwrDIy9LMxT
bTXBkBviAVccGrkFqaXp49jbgkfLo8ZNeOCPQG102d3kgALNq4S9PVFeHEFXJDuD8Wu+RTCd/eQg
duTwtCd8Y44vbctgzj9G63rCWTrLvA+yur0xieBJIGhsotW6Kc9QiEd4pn1Ra6IPruPUVI2jL94G
UxrlJN1LvP7YJ1lWta6EqtAG7SZxri7JbhbN1SXmlV8CpKWr80eSSPtniVcNfHvsPPUAL1QPmE2j
u/0riVYcia3FK8q3ofvwsrp074LYqi9CeI9jNw1zofSBlVL28Fl2kykCdg0JS/jMHQLb56y35KLs
Vq1+wwUHLVHvDz+FT3rJqt5EGSdFZ0OeW03lG8a7+V88WhvWtEVdKmgVfXPfMs2VHY6cVIde5Cxn
LIC9NF3NluDNxQnmZYvgPhIscTL+Kl+inHbnmY1PdJ6jSeDrhJrkuHIlBaQLNR3C30HQZy9iOSup
ndo+PxXq2KI1/sOKM/vi+6Yi3x7H42SZc/mEG2s3WdzXMDzvjhIY6EnTs3MFkvsWyRmOESDFYR9s
MuRG8dHRMVYbEJqnZMoKXpFkvEFao65804pac0hkxT2kwdz3eHohKHsNcI6vLKMaEcpmyzKbHoxU
AH8YQsJfxfDHblKdExqRYHA7Ktn1f8CwhKme6BU1yW4XGNEgTsUOTLzWnoSB2JXVKac6V4AFu8Rn
uqdK2b3qK7REqvtXNLCtIdRfx/1kA1rlxNxAY4WqsqdThDTZKO2rng95ZpiArUv/puCjjzo1gxE2
eOMpuPKr7cJnENW2i3agkcC/aiaXjj5++ye1ZBeb8BSFW2OtFSTfYBdq7GQ8UJFd+98mpDoJ2mO9
ML+/OQQRy3NPf2l6L0iI2L0FdMwv1uwEaDu4flUpJ37Tak0aSYMoZo6mnteTrSZM75IzKrOYMH7+
gESaGStL9MXzwoR8w/Pht+S2+o7xR/FXq2QnY2NSQZH0ltmcP73vLMWjV5uDpgeLub28xKIGkJyD
mcltv7uk0IgBtpg1gHcIotHMBPNkGX4yGtHIHcXTJABJqJ4MJa8Czk5sMACWoFvhZQeMSEPVBZv+
fhGJwaQ6IyMmr6dd5TLcwW7gCZqZioAFqlwMP7X0IC6rRSOP75dyZNU7A/drTBl3FTZG5IJ6DeIf
KQeXjUB/ory597BrPW8DbIHKjY0lBJbfd5mNqLGJEAHw5wMXMP6mFujgFphvRT7P7PNIaWgJdHXP
dhRqKQIauToa9hxKaWY7svPUzPRYZlSiJQY3qXZYCyIpsigkERSdy/+zrABzLJQQbmnOlBNyPyHO
RU6xgElGfAyfi3WDMnP68NsqH6HMT6y2vVeJomLE1l/A8kvoem540ZAPuxwOGgx6gIROl8c68iiF
TCiMIXWbNt32Yr2bgoWEqGaybuxjGW5o1GPtyfz3sGCHS6SrdksN/NL9M0f7wGeSLsw3RmKYx4V3
W12aNY/WtUPpJ3kBWTBb6BeNBoWF6GvNA7RoOv69rqAMoW48GIos6kWjnUFEUmgr7a0OIz95o4FE
sq2UlqaPjb9Pwe0JiGGWFtfgyToMBnzitZwajqHhnLmSGETO9NM2gc9VCIlG86FEU7zoZqnYv+si
VOGkNMQ1rrF7F66Fwsv0fAHTsv1+8pa4a7gLef/8j4R8OXrN6f/It1XKfH6nYLNrZv680lHbeS7D
cDS0WHPJINQenUJmyQGqUBhAm+IGfGIJ2RZn63L9vDC3YlloZ9ik7tCAH15wVuYNIqeXYGgpPvE/
P+hVJ7/bKsRsdHhK3OS4OVq4M7gWNRl+Cc77fLcPaz6AXeVFvyA5em6KfcWDfEOSx4Bfyyb/QzAE
wX9W+GWigY+H7dpPr7+FEVGGjjDRBwBmy3OK/Ttuno8//N9hmlEQMkrLIGv5SQ49mDjnDc6l6PQt
w/z+6sBl77j69D46gB9mOzxTKuykR2jHDcqxtko+vMwN9gWtfEXvQluLk5eAoZTqiwhtig4lArk3
/NYNcpylUl6h//FefB9myYtj7gkGEYWzvGanb8KiGsp8bAdc9Tlz0UYol0pZawz1NHobMb7sbUUD
DpaY0n8yo/MBYDOygSi5oAF9Tr+IyJqPNdAllJqhMtOOBbhEGD0MjcX1heGHLM6EGxQMhSmN8kjf
dY8ZGZ7/Ec3pFVUYsMpnEVeyyTVLBilST9RD9xK9oq/tbOGBHLHZB5Ij4UVUwfDf0kNRAGsZQdvz
wvbohZG9m0SvBmu5ocZhf7dg1c8g94AGueblacQ8tivCgRSQ9veHUfRvddrJMkBPy+jYAFttCzg2
uF55AyXbZrDakxcrd0aAB/GpbcHiwEClBTdVAuVV96HC/aCC19F+jI+btKJBwfkACJaJMfQ14sfa
pk+c3MNJfAz1VbuJTa/HJvVorpDjBohkT2yYLPvQu1qK1VtaXeVjA6rgwL/nX5YzrAVU+kX261zG
SJCxIe5eFut+HS5FEUJoBQm0m4F/1k3lcVqh+mVjTIR5CIHFDKjllyMFOmQWSW3etxGoWAN6Ejw2
E2XMxUPrOZ5/Wpj8XR7NnA1Q5Ps3f+ckUkyffDUg82MED/2DggyoSJhFO42QNg/2xYzlJHPfdfkz
QxJDLEV11BT8oV32LxsarJZOhKhEYMREsZKVYAK7ahm/YVj0zfbQ/1GgziYHqC9bTVMbp8OsiDt6
VY9sdlkrDQwZGFIT84bgDQjdCim5yX4mvzDBz7py0ur3bYhqf/+qtkQ4+1SobB6NVlgpZ5JONoil
e3c+XlkOcy1rTOS/oOrKYmdXviGH+gAiq10hCMkIWSbCogQu5yOtqJo7MIl+Hg8DaFcz04CNOAGH
iO70wOUzKaEreOMn11hCdia+hyjDG/zK7J/WdosLu8CsJytWyJzn93YP1Uekk+47dWIudCgMt57E
YSIbZ+gtc/hOcjZqEHru5K8Q5LEMkGTnGiQa7y/u/B864viRxNK6Vy49oEu+vEc4qFlaVw0ddP/c
3uBAPnpI5SVXYUyhpipK6W6fGkmSBH5uJ8FxucDDimkxQdjtjbHuyvSkzDbFbz3xMLQC23u51m6X
BWxDhDYSqHMW8GRGBY7gZgeCW5bqSwMO+FM6JXYPYB+bwGhgj8KgcR9+2RECHxjlutboo2+6bmFN
dD6RwogPLtWoMrIAHyMCntAmqPQin5/lK+iCgOkctA6jHtQji4olHytnvuCI0huWWEJv59N7MCD3
yhG65dNOJXXdBcm4LPHwi996bE4ORxDUfaY9oLm8spBzrchClWdJrltJkXOlhJke8sqR6DBDhKeH
xurdLLRaJFOe2wdUZPyeDQLu8ztxf9BReiaYhtFkLJoATgGC/1z0DKF9GZAEZ3dtyQKjYzvqx5Dy
asrm6dUL/jBOyd7iXUsZWGRtRRCPs4afCGSLLzMEFaVZ9o5G2j0pEuPlqAJaLms03hiCxCze+EJu
A9Ks6O3KskjFv2qfCRCy1lUeGw6l3Z9DDDZ2MWLrdPRevyBJKA/MGDaUtrHmGH4RG/q9Me7361bn
SFngQXZo2SqNleAkaVhJ3UokKB7dSH5RtD/qOyd6mizdyAb/Uo4x21+VV7ZH5ebb+ogc/bQsmIP2
D5fxW+J/gwMa/dPqYyS7hfA+WOSFQ33LNHqY90ModOuxZB9dOgCalrxmIsMCTXtYXeuwjXy4C6V0
kne0J9KB6YU5/RCy+yS4d3vUQ9EtfWr5eHCN8KmVcWDg0HBAHxOboI2S1aCsEwMQ4aP48BO1Lsra
4MLSH/Ld/f8KD5eMaHcNwM67cU3wrW0x+7ikaDIkkkPjM10nI/nxbPWsjJzwiZQcrHTbIDq5WOgV
IvvngxZ1EH6TPbkrmBl3Ca2AALbdysoRssAaCAauBgDo7nt+muuMaSW3/fyU5nsaX+ZNZAqgEsZQ
EmSLI2/z4SF8GzU+G0KKkbusDCgZskKBspFW2nKW9STx7TJHwDSecEPhFfTZXhyyYoSZhqGlstJI
YVfY3ORpiD2Mgc13QX8SRbq+4bQjNUAJuIWZ8DXHqzupNYol6cRjFg9CJ9bXZA6ZsYoJ4yORs3be
Fbb0ZDAud7/5NT+h2JvSf7H9xjnTK8cd8Q4UxgdDri3zTWwPjKASxclheRgGNSXReDZxuJrmqkQX
K7aIKESe2IkPjofQtrF7b9QSqOS1YyMTgC/UtMdchfegQSv4pyvD4NQEWQsIoYLmTxiAaqVegrde
UqSDLuP1YiJtjWlDB9SLkfhBFgKp+iJCpT8z2QIlAekrjTuIPaXQbNYtuZ+l9DvuQ+A0AUXuz2Il
jfVjI3xJc49Y+0PMH9wRarZILBgbVlZGc51YRnwgvVnwf1+poT8tYsDi6YN7BZ9Eakyczql1FRA7
l+U1zMXgOI4qkdjQPuvvh9sX3K9AqpYbTO9D3fIl67EZiarQ6hOSaHLaTSs+oSVdmBv2KOtaxSEC
YwwuVfSEvAvOw1kOpIsQlyhxKgiNtp+1rDwf+dX1vKQHsGObWxge45nO+Cd2xct/TWGoqCQuQed2
hm7BQ9ka+M0t0lQ2N2R/q7LR3uF/BGS+DeFHQDo+HFjhu/0jkAReos2cBxoDM/KqnDBrozfXCxKb
qjqSHfiMi+aEBqwyKQvKiSMlz/1Z6PhpzJL3QDO6+CHE3ewGlJtODwNIi8/VPbXpeQjwIAlAuutv
5cnXvL8zXl2uKM8cygy6tkld/jUXXM5KlQnQa1qUcmu56Yut90Dtrko0n6muruUvzgU8xhulNcDB
xKOb+AEaNWVjLMLKVhxIKYhbCw1jYp9h091edXmn0zxiDwI954nE7TPcDJPp2IgCPhrDp2rAu41f
sJDhOn2EnXigQLDMibPlOUT4qrZKyJtEAhltRaxhz2DWZdZ8q/CUsW+CMN2sM9VgmvC7K7s4H4PR
gI7kocVwFGl4Y/JxnxfQoyx/IEYJqbghBzV6VjADrrU20Rl3NGg11ZrL9WjwQSYXQVVHGbeBaOPu
9d/K2ggqwlo+35Cm50upnFuOajP77i4Iz2lZ6RWz0OjEqIJzxEwzj2/zCLT5Nq1rGhkLKPxBK+JG
qT/PK4Lpgpb5vv6h7nXuk+D6I+BqbYVivjgCXBHcX1VDeuAY8S1/jrcwI2F2zItat1f2fHRErh2U
2YHoz0bxGmK8mkjgkRrEJF7wbABOtNpEXejvGVJuUvzSBYlBBG0XHFvFQ4uWTe1/8f+XScsmtnoL
ZDC28Bt+aOnh4wA/WdoqCX6ov31Jo3xWLtOTGnhcQap90+eymX7HUY51PCBfDEfLpsRYq6nuFFqB
NcXE8Xx6sr4o8r+cY5oxBXKguLqQu/k/h3KCN9hYi/ew0/ftlPzpKSzIbCJfcTRrvSP0xOF7DAL5
1dHfM4uFvmhMgIqwjS5lKI8x9qtcqTC/NhBg35zssL4JMsmFMH6GTJGtKWSscd4wl2knzj26ko14
DTPdmvH7M+QKlJCZtK3fa13dQYtAzt3GgDObt/DebB1+FILpgChN63kpG73WXEMCLBVV19SSUPKF
4jKoUiws6LN+/3FigKYplQH0/u4rxJ9yBIaacbqg7qE7911NsrV3ioaBW9RfBiNh5lvi65bjM67B
0lJDfULPBVItgDdzymaKQQj809I+vIs2lGMJUAV4gibFXsi99zMapDc3rlg8m8lT7Kxr5HkJqOK9
gb4hOYTJZ2Axn7Ta8iVG+neUknuBRphxKX6O4wp0PK+hiBIIM6wq6UapRdN2BLTgSt7+rB8iMbPa
El+2Wl8HiaSdqAOiHUzj7BXOI03GvNUAN8rVUFn4eOiUSxtvBbZzCaWTSEh9jOqwe6qLghdqzQ1q
7D2a2FDfqPnDPp6RrdltGfLkxHP+Zuuq2gbF21c/ZY7RLVmttf8j1dUuRY6oaLQ+wWw31Y98HVqR
ecSEH4xDa0MQcm/fkY67Z5kB/vFyjZWUbERpPgPDhf3nQeUXJJ0zTR6f119SVhi/tT0zzAjTQu79
PTiiPhB+gl+SGwLIji9ItmF719K8b2wQOvwou1TLRrFBoRKb0XrE+UZrYMmHFw7fweevIGfbhDTa
CWvpK4vC7rF1PJ+JL025u+QTBjt5wyfB7JolDiBeAZyuzaBmuYpWQV/dh87TSoAb3HdwU6C4rqQG
xWI9vn3y7jYFM+Ct/n3vSNgCmVcPaVNhe/sZDLsMzwEPgL1ngX/N+cBxLF3hdHZeciQJJ4eep81A
iRVHUEjOJwNmTg/TUK4Xg+WSQIz5nY+KHoM6bYI1Nov0ACnP/FHam1glNTmWW++ik7Fvsu0F6Hel
GL4EO1y0W/hxPgxWBtmqNyF3J8FURzwuepkkBTe2N/vZJ4zmkTur+X7LsyYiq32RuQzHMjM4kM0G
92PjITETyL5DlFjkfI27KkY7EPjSa3uESP+lJfKHwEn4+WnWRDd9lX3oxSfcb3KrXQYsE1cskM99
wE1YNhqlC4RdE2T/nnlEgq/ZxTiUcUfbDABBlGchILuzSIk4KEswFQQl6IHL5bwzyXqGvOlfZQpi
yRHLW63TUZCjkqdA2vwJSRUKfkhXFV3/Ji21+ziKjpm4gtkFArjFGhBTxIF3uKgn7ZVg/4oc5z8B
JBf83yxMVzGc1USyoIPX8nEI9bxC81oEhbS3w2PPu2ZqtSeGMakQdfMuO3L353KHI0TlmIKxFI2F
DE6DmPOBvq0+05af6Ip//txOVsscnsKhCtxr4Ix8prrIhUbwkUxTPn4ZoUkLt0NMjy37J2163NgB
RVmkMi0U0VI2cOqK149HGU2MCxIFkt0k2gqcXn3/GfuXb8L0c1d+zqJKJOYHvRkRhzvSNjnGPtEu
O3j1utmH/OLloMaITZ4E7ky2gJLqLBj6iiY+n8ItO+y5muqUMx32BoM2wjalrqA9Nud6tTahyQP4
9mkoZGRZMf/AYxkF71+98G5ctbR5zHG0CUr3shdX6g/fNvE7B2gihfc2j9ydsPcZJ2NNbafjUQzw
nxhe3aNKNy+yGimLRM/FAgzyj1B42z+Fj9anmV9KhHyrxFFVQqVq6zsMKw3UxnvpXTynWyTj+BgS
XjG4wav5cFwQh9+gKfXllIteKrorVitYR3S+JXB/rQm2BlGjv3UCckmESIjgss6+8NvwLkwqIMAN
5sMNClZ4T4kuZL7sNIQHbZyRwhuMA/u8by6PfLRZMnN6ibwaBF7mwYpIb3Jgj4k6PZQs4pCNq/Vn
JadMp44xRdnYhh8BFkYGvgoMJ6+JHj7khMXqyU0uksqQG1z0DbNovo6uUMtgNakQCGWZvzQWZbz6
e+z3Zofb7bqsKN19fB4X3z0l7KKqE505euEGabTF6JLjSI7egDAZwNK1HKT7NAJH6S47j4dMQiDi
RS7JDTvXE/05gJ4a9hA62fuiBH+HxZIMvSGlTf6jhAIYKCeSY7hV5O9d9sxtD0DPpzNln8MXuxlC
XfhyrOVYCjJV9TsskTdBIv67vR0L2/HV6E/wXbNKCQsccVtAQ2bmifw+bjyNcvfVRWdXdbZJwKVA
8w4sDEFbz7YgrlWKhwQw3PJw44JZ6qeOcCzI/T51AR5u87j5yQtwXvzz5hCtFJgJoSjK+iv61QTI
5P4Qo+AOa/+Dw7irrvWfvmJaEPpVLEquhB1KxJBah7nYaEn+r6onGaniRAToXmXiJvm9tYZrh2Xz
W9PFdLxklSvlneteJ2BTHaRXCIjipsKjTm0OGkz7VJYxTxfhxvgdDRGr84IBw/YzmJlVpdpW3oGC
E2h6i7idCsKKL5GtD4TdSF3LRSPHOomTcvl/dolL+Z/XQeEZEUnQ5qaVqQq0k50JKLJ2KjUc5dp5
jy+IY5xXDgHzDomNk0Poe+Xe92CGDuus/w12ClmolCKddybS31sI75BgRWY7GYVzgwMAqNBSvh94
jk+rgY6OyQds5Nd56cBvLQdpBTHQWKiKvOCpFwFYyTLkGGHstbnXPCRCK6HG6VXzOg8U7tcMirJ9
QqBdHGs46USlUK3SuV0h2uadrbBWDUDo0k5ufAsRx0j7jvXjf4njv1xXW+IDXapKMbcpJuyDTwrI
xkofLNif3vpquPYJMImIHSFVK2H/G88UcijT2FaiDs6OrxqDJxnswdvmwOa3A2+SttKtS7c0yS5J
tFVcXQoNCQw9dlF6rxRxsf9v+zRzrXZ4uqmblTr1HYudrh1hYgzJJK5sHnWhRYrDYQj9v/w8j2vy
DynEjdyIMlHSxdoyYMTwx7gvY6v41l0DU6HCci2RefiAEsRy1y/OW3EPOp3LJFFXTj5Vd/G8jK7C
Vmgef4etWIufBNEUS+JrQE23/rDLxEtJKZMCIubSOK+op6J4395J2leMO/Xfs+9Qq96JYcs3tIBl
wpm3AAKK9L0OOwG65/u4i41UFAdLRhHemISzLrKobeKMEO8Ui8GleTF0u8S6Y+AGSEQvBL61rZ9x
U0bRw7bVT3+e3NR3IG9Hh+JKpEYkmOuGCzeEB8BnawZw8IPawefI54SEx89aClYcq6Crrm3T4jyo
k+GVWncgF7lWEe10fh/CKnmhL2T/6r2I1+PiHpnFxsdIQPMDtWmK7q9KIvTFHaaW5xqLpT06t8ij
YIPMyI7qc1y39kVHXOslAPobxhrED2JLvTnw05DTTJDgn1f9G8aYSpzb/ML+dqVr/7Ip2ek5Ge2y
gnsWKluYku4m0Ik0UtQnXgs3taRkw1Inb1Vhi5vv/S8FSlRn4q51P3N4OLa/FRPRkdE2WdReKgGP
JrIrvwwE2sjSnABed/AOo70cQQcah0LkO/Tt4N8WV+bPewZ96wxlRi2moEQJo8X8xDDG72BMHt9F
JFSf/KpezxKyK7Ay58RiIN+WIVLyfTMhuWDIyvdZEcX5CEw9nYCtFSTaJA6IKn0oWlkZ/CtkqiXf
n9kpjedvyhj1XvoLGAbdIKlx/6mi7db06n2PaECufMti1AhnhEquXVfDWYMh7FeUS9X+Ii5Hj+Cq
rSjWTbwUT3XTWc3LwP37sziUBIHKyR0SfBDz+v6JOvf0Bpk1ntrKAQiZpiaxPXF0o0HCPGySI469
3kOfrje4znvITCqyIa+DRSG7G8g7okzS8LWDsUjTg0dWN65A/9qty19hC5l4AaNuNLSucXd0MTFu
KN/NMokll3w6Ubu5tYeasZYDlS3d3o3aN6grgbrkGk4JzGncyO7oOiNOO5pALcIdujt3s9JkGo+d
whfDw23s2T/9BQY9aCSgdWdTX0dzK/M/kCMtFYHkMlq6S/SOLqj4c6wl2u56c51vDiAzVQP9u85x
+cWMZxMPIQWkuMCQfurLehXWs9oMyCc/Xdvm4IHL3XSD4xNAIrxp39xpVffK10qUnkJCU/RWDmpQ
J0eMGNFFRkDGnVWHdHH0trhZT4KKBmiCk8Z1wVlep1vwRlgvGKuTf0xdP1jaMxMKL8MMJMgKIX7a
BmkAfug6YCe+kLChzjg8qtHX1mC3Yy4MRtlOGv28Z9dT14x7wetbUXFMUZQaKbj1SCow5z6MpDus
vWmmaBxSImxAiCrq9QWkcFD01Ha602HUaj/gDkZC16b9oqcsopLTKo8UPVSleFv+PGLxyjx77Gqp
mOxKxL3Ly01Gx8B7+fJraVNjhtw51KLSHJPDCq9mFOBbkW7gJCl8y1TmDuQu2lNWFZRDV3VDRhD3
zbIORSjc3/px+My9CDkC3QlAToRtAl2MrgJXRo2ACHrgDSe+/61O3bRaSQnwKX6Ypwd8/5Q35U+v
NE6BrReMGkBG25bCdxxv6+xhNHxNIZLlwqSwE2XgCbFYtXrBQWKEFkteLbDrB84hC8SjWkatPbPC
3iyZPkbBzCirGgYS1yi/AeIZMa8q3PG7sELArXdYyA7oC2Q++ESa6VtwaRwzxPEhnc8uRWdskRhf
tZacA3hECf3revG0b8fQhJOQ/tUG8BMmq6vFYfjQ0Es8sthyUWVBEn8loWIWzoepviIzr1yl7JUe
TFzICpy/lGyba+nv7il/H01kNtE/ScNytAennchrIXDu4Yd0MBMcdXCrggf0RZuyaLuxqARxVQ96
wP9eYxkLsJ5AhX13W0JFf/1QxtWCH+R4YjH1syrz+JS/o/qvoQy03jqjuhbGi8uF3Gg9eP2K1LVd
mTFrtl5sVCQhI2m9vpoXbDidRR/0buTlIvLsykPcuzdHg5ssAdhBA8TsWulqVyW9Ihkevlprb+o2
FJCU9fJxEv0qBvtHH6B0AWxkgXBqV+/balEWfc5oaYNrVYKyRL/G9w1VYk5HYwk8swIh4KE99woT
xaF4lYDKp3Qqq0ZI+VmJKkWEf8YyR8xr9ZoU9uA0TtjsLr8g04uUDKA6SLCdlhg+IisYKRfyL72q
2qS2/KlD8pz7Pn9m/Lq/rB0qzAms+b/KdFZ5e+NXiJiPOGAGzRsD8F4WrmBjxOowKQ5BG0BWugrO
27mtOopURxGg3Fc3AXKmgPOR08zfsBA7r0KdIwjagtdUDh3qPZWKkWVFmEglvwYK61FAy0Oz8lJK
yhgoDPnFNplIgEwEyV/SIrxgzcPBaD+dyrmjLJjiTiffCje+51QRZrqhItW8hNToLG66zGkSga0k
pdCGXFyqwZ1kmuuMzn5gi/Lk8GX/esXUBjkgFT3hx3uy5cH7JHcSE+YIytUgcoSxzhUUQyI30tSj
0zJXUKcK8rPbBou8c2nn93RXMp4XXhJ1yuluQmHgt+RXmuIY9QXktx2mGzmr42iH6Nc7KHrMS2Rg
yZ6uPnlpH+9RrIpSG2GyNOyRvaGvu4+J4ZHyKo1VI60WrjUa4j3n2cbB4KQqw9VB8Q6XA/OY0l8E
QJYZJWSmzmlagTu/Uvxf73QCQy01VbPcEoXE/bRDCcH6d2J9NwhquQupHqGJnFyWztfHHwKH3wWb
1/B0V5whVsjzqxsEDXbVF41mP71297UZKX67szfGVUTYH2CsftGpukKaKNTYYj05nnVGT+1vOTx4
Wwn/ozzxrx7mndTivFbpvkg05+yIy0ZvBFtxYzQZuULQh9KbUSy/p5M/6SqWtASh3nKFLbkuh1zO
6cana/RR+Oj6qK6etTbVEH5PkKc9ZlkMAmqfGFSbF18Yn4YvQkxRZTEXOa4EeaanpNFSqPFlurE9
xxf5OkO+EdA7ZV/+P0ITec6Qa4s8pg7RqokrwjEKMAdSH9hqDmWo7Te8FywwKASj1Kx4vBbi7n6L
H4Duhl35H4J/F0+ggPFqKah64t2zhDLLJlJv/qQkC5N9Pds6OcQj25shyhNcEVfJsZ2MD/hSm9Ir
s3ttp/CI9d880JgtHcYbhL6CFD0FiCRTZ4YjFG0ePiENVHvgwi0QMDRPuTDC/YLPURMeupREiJXN
tTMdpcQBhNvCEsBCdIyksfgwt/hjhENUPwJ7oxQlszJZJU6DKyxB7pMti2VMLzz3WNdHjWJgug7H
7IRKy3arTcEpG33zQtLEIYTzJT5wdxE02yMDB1lh88duxN9atC7cdE+fu1W6mYiwOc1bt+DzMUPF
EnqGE9qTsR/tdF65tmSwndj6HJtNAy6XfoFTzT/33hAvCeDOHCSsNn2GIugaG6Lz9q/oDnRB9FDi
Yqz9jsbLy8KBQvT5PjD/KP1JOpIzIxikHLwHQI5fR5/MWG/z6Iop89PzAn8/Ycy5dgqFS7UdZVrJ
5snQ/5Q+rP8fJfeO4+UGy+mvkG6vAXnITPKOcvWZBd6/stPse6Kxv/Z/9b/iTt8Ijy3XgZhIZ4qS
hIE50hBubJflSsqJkXh3AIwH7DTd0GnFNCAcvUdBQf3jdK2khu5cJxzUV/eWVWTlYvCLQJpfG7Lv
A7VnSXN+rqQejeWP/TUOKb0PJnVtfm+yWKnmhfuJDsuq11apTe8+MxkSJjuZIsyC1XodUwQMf5tl
17x817f6lw9AYRz93HKi+yh7qIBxC1o2G0n+6cm9+GEX2ox/fAUrxSI9Gf8ctd4oJ4RkHDl0QqBS
FHPEZ8x75JnrKJS447XS72X2ZdLgcfikH8XtsXBQufZBR1C7EMDbcqH2IKri5CEbVh1ngS080PjN
oB4p5ZFUly5muX79TXU35YRp7CMPNrccsxr6+d0dj/8A50em18+Qdr9S6tem/cGiEtR1dR0YmuCk
d/B2XVZPR+/TJ9CsCC/8C9hPQ5hhaTDZXbvj1GI+8KEqLUSPhYob25qw9MyuJafRfBEz8g6keykp
SPPwnmOmopNSe+CxCPXTjZpFqUk/WjUNuUir/WeaZ97nAhiKXZCvnACknbpo7sb3Idf706YEYjAa
FXOWY7Jemmhr83dWC0+9odhS0JllI6s+yRK4EMA0kZLCXfDAAZPwLLrwZRMAE2pZjuRHgMucIDSS
YVzfAr2RUsMWBjZJqG6cFBEjvchH4+25hj2WA178xsQH+sswgJXpBE9PikMUiqMLBPDA2IkAMMXV
l26rOYHaXbPQNSj7uN1v00YWviUCS3H7XouoQpU/Cx6/j9vbasGR1zNvnN9B6REKez2lAs36vsWi
B8Ho4aWxur69kQ1i9bwyH1AL641wPLei2OYQbP/UbJ9cpVD53s5xI5BQLxCbT8vzqTGvDRclc00F
k4JyLubkhX56gadNCbBGrimcxDh3YP2MOHKbHMVYpTXxumCQUFq3xzempeDWSz/glhimms8ygjGa
5M0LeKzVy95Y5Eo7uzAtwYJ1gQ5GibtmqKNSyKJogd2NgoRbCxtbizzWaZgW2AdOt8ofNJyqrpTI
ETKM6SGhy6D18DmnOLVO/HtaXTM4cnXDk5wFbTka2uk3i3AIc7JMAe2P2T7qiNgAdRIFsG8yfXFS
UCFbVIGx10aLdEsKgYZ30Vq+vRvL6x9wbfj+ZkUBMRP2mozcpzKBELhZsFZeyWdZiyVVgjXj7UnZ
dEDuf4oWYiyoXcuMdA2z3vYpHXLjo4PRSq+nz+r50Z8k5MNwJjcO+OEGowDVkEVpduwjDHSbFsg/
CVyYWFcsRP/8u0tvFUXTcHxasq9zjI9fI/cw1jbzdZljMTtPiswBsl0lbEVNjcwxPGwg35EmIsLg
vQfVbfqJsJ3tJBp+Uu8Jt9z03l8cXS7H8Z18032DcCw1mgDKnxKP8NHsI4iwZudDhVy6mVBxksZO
aBZSsNCfH4+OnirwPYnujU1LSlQjOfqQl5lS5IrSKlWxandu7t6iW/LOt1XtqYHm4IcxkXHvLush
SDWGcUhughOstKmkP8KSahi7kMsTGHWs4FfedT3uEsl92HgDNLMIUjeEr1sojdxfMszA9fMR8q6s
6f6DwrcjuPuC74KyTFTgaG51lmxj1VkCKPdC2T2EP7DGWmI9C7lFol1cZViuZ4mjVLrL59xPoIVL
jE3OKWHUF/DgulT3xAED+VDf5HJxIQDZ4Vm7LpQDKH2iVDAu5M6/w4ceT+VVZPACIMMf7rin7JrH
xC6OzmvW69uFjFWt9rBWPbbfYybT/0bijXHXbIEL/VigjuQUOAArzYHn6YU58dipa1B996H4HbbS
rJRN868PQtlCSAW5ZRv9OtuYrO47tkcJy2lgyDVZUDc4zD8bXzNC94cargdz+iIphwyAJYlySuUk
DCOG6EaU/E5lGgm5owowxYmPoQHeskkn4TE+ArNtkPWfvamzx340OxhyDLIu2NGXrgtzcS/fZjjc
YX0JA699lDCuZB4JufywLdTSAEcoPPkKYPD5HeSQAenNMJH5xsqxRiW88LC9MLaZLjabFJHzcmi9
iAdBHCyLHfQJcZcwxgSXZncEreLL0d2qCUPSN9iamgvBLeMOmIgx/kXn2VrgOdvy2g+6iU33RQ6C
MDlMjl1zIxMdO+5uo/nX+mnJYuzhVb66auGNIlAa3dDQ8Ua1iajRHz9Af42AApkO0ycI7qKq8ulI
WGtRJ5HwjOeGkkP4K/zzYqjJfNQ74KgltSjJpPCi7KC8dkRFBijGRe9aMkOS4PZLtm4FEXaWEB1C
SkO1ovsKa09k0mo4hvPzgbajeYvIYXG/30vfkjvW/Ppx6gcWOkX1pksa5GyqylRRZBhaoTwO8MYu
3xFuTF0cne1s22by2Eb9Po8yBnLQkcZ5LWWH+8c9z7iN+K+uhtMAyIRehKVEuuS384bg/XavuKw3
Wi64eZnYTjdBD0NW1ss0Z3B8cEKGjKIBD65FuCci2PUXpHYdl2QjZXJq89xtz4ahkjFy8Frhy0ix
FJZ2yqDgd6S/10Ce5/sFy0Z0oQGLiXGuJILjW0Eox/TUc/9Z7nKsgAT6fAvH8J0AdOR1ZsK6vHdy
kb01+pmJ8Iks1KtmiNouK6XSuzNWzTx2+TRORnG/DYpAuety5G1tymhTF+FSqSvMIDA2sL4MC/Xl
ibD/kMrKKV0b5yNXBgw5w/GhuuUze+QUxvoYfAJCt2JLfhFTtKjsOqQApQHz9NLRoKM7X5GLzRJP
L8eOOHQ2T5+zFoLgpgOIh1HgUafMidfqPqbGrgzSmBDp0e57NqZ0DbRtMHAfLCvZ6qe4jOkH/2ro
g1dNOQMXhWV8Buw+BpiP31g48k6ePyT+j6tDbCPlpXb2MEtZKQf2yLAZ1cv6FX4gR5bpTw0mSxPQ
9Sg/ON8Q7JzMOFgpS1RK9cySnB1pm6IVVQdk8zdSfX2KfLkiPfT1CoDqD7y28dyvJB4D2FPeQUUT
OY86Vs8UB2f+ZhKIMJeGRrP+yy52+FksEkYCWXhhi5yWQ46wqfnr+nm58bTTz4lVylYjVHvcA7KO
TL++ibIPwl+QJwaC3fYN3V/iuj5M0wDadicyskp0/2A20MdYU4o4+BKbBb2uh37GWh1XKI+aHQ9a
p9pGAqMx85s2DvBnatyVaP9YRWkHPQ7/6cHVZdJn3ox5LtwN6M8UGfvPMIHhOS/aXuU14NMXOoul
j+j0Cp0yxD2h5rjhXdfg7kHfRF7NsqtxztAiNBLrrr839Xsgt1LE6PFfF9kwbRVKKBhqDoh0PQdE
jEXNNiH4AACwjjBCBvOM8p1TThBB28NH5gtyodAnyaBKBM1K7k/iiO1EBq/QdziZ3op1amAhcIuP
WjO+zBPiahg0Dt9A3C3UQrDRYSPgUdAgQFEaZiuuZknY1tk3Y4rV+ixM0MbLHwg+n298p/kr8fxp
I3HlmKmL3cODiJbBCfLQkoTKVWx//ARoQe6C6TbMEiSOnvKt0QmQT+ZHjO8VMe0c/hOxULGVG8x4
bLTymSXYB+iMZ28fVGY1auKVkbMQP2rn0bISaQRq7nmHUhEOfBFxJ6yL4JFa4ZwM+m4jjg5Wqijd
mZUoG8AyCgrNzY+KHuZ0w3kYlpL45pElfSupQT+rgOgQ9AQI6HC60FJPsb5lKfCsUYerMQ/Rxk7j
A7sJsKvwq+nPQbwPFMbhhXBaodFo3vE1SVrAGpWVd4MAry8XK03sFaX6tvpMUgQRx3eqLm6tIpSN
Yeeanme5aIGzRVQcP8ziFnCkcKq+oWP9OWNdv8G+kByt4HAssjesKWSOW1X6WH3ppN0GPA8RMyYi
1L3woCtaQeRSAi599jVQr+GJEDdB2MJxYIZ+LZaT+UORXFkpKD47Tp72ztZ6pSS274vHodGH75dP
0+X7/ykZwwuTO9vFV73HXcBOG3zWQH33JdKb2sGjy3xxpxt1Pl4PzP3aoG2tQcWlBl7vUlNzpiao
Q+RiFuqEGTP9gH87yExR08rXAEADxVt49VPiLhHGRulHVIW1T0TvlUhiVlm8WP8FF4GdLlLumIs5
ySUyw2UFxlfUFHcd0wW/r1MP2hpcQyQd0qPvPAcwB2FlRXimY73Wl2HLRNCiVLu6JqdechABAqNV
a1j/HtrtzGNReGALdWpP+u+8rXUd7Bqo7j7xk7TRNTI0kAksWYfGTv8GKWAEW/9sYkZ5YbrflROe
ytWOlkECCuCiNvblN4pVSRqp/PdjcB7w3j+8B7DCPXdMNqUxtD+kGt7+Htg9cyiD7XFpfAJL0wq2
eBBgHKrj7vFbic1dYphIxu8qRfP/V/e7gTYA9C/B1t4mz69QAX+lJtXsI7f3IbdUiwni5i+K9eDU
u5UeCOy+bDb3KpJ8gJL8fhYeWLpe5dPBAg8tunMqgVJ2R+b4OepF7PTrkvxH4rECtmZt6r5aaPpJ
GWZvsU5T0pFWr/QNZz266AT55EO4Eild+YkCA/xHM3NLs9kNLHmNs2D+8Zp7B4OiM0gufEu2PuP/
/vcv5yommjkO331URBF25XIasJaptSgemQkJnhU2iPfeyyQIYvWBMM0thohn39c2+7ifTaSITEH4
mN450dzRr8YoI7yeeWTHRES4o/tUrmkK3rMngZMYSrhlLeIitD6Jg+5ebTSlB3W2fjBOB81QKsL8
hwmqHE6FXt47+q4uLZ59WYkazirZHBDTsrDhnpegPTWm0KH/XePAj+MQ/OXk4AIXCpCt30xeMn9h
xwx1nrr0EFG4AL12y1hQSWm81vzdysy4Ukpu2s2ZZsL3pVDf1EwyvoR9Hnvf5YJtNfsOHsqQhhxd
+KRFRQ0IbyExTcwAq4ortClZGaMf9imooNJtuAzsVRVlmVAsS+4XscvYSGn06poAuasiPgj52al5
YYHfrOYNq861RFU1HpSSSdceELNO0DDdxNXc+mvPspJv7I6838s91AlUfmGPqDxblaM2g/J2XL0K
W5ip5TV+Pl/nRWoPTkCjxkoOI/XuqzL/KYuFICnoc39Hl0K1l1gHxz2mmd+zCrXVGvo9oxCoNpht
1lht2aOW0KPJXUVXtpmHyiPY1pjLA3wisD6ZhakcYbOAeLg8e8w8iAqOmbdj2OoH52s1x64IQqYv
BI4v9vmmOSsz+AxCeoHgrAqwqEHIHQzVIAUdlN1bY/Wh30UMZ366s/UvR93EhkjP8+xBz32etP9S
R4Xq455tuvPsOLT2gYfGHDickedJ0R4xj/KJaTjQsL3fUui3lACVGYiIz7PRwD7vkx+Zz2jVoFu7
V8OUa914JgU1ycZ6D/jpCsL6X0xwAvGC/x8AeYYb0p3aB1xp2n7vCsvbfUM2vOGr194Y15iPWBPq
myG/RY8LI4YtGRKpCegH2ocRurLCALog46Ln50yyY1tyHS/aS4ozHSDosQ8PruO6EhgM9RV3Eabz
z+ci+/9IZpsDwHqQlQjdAk8oy7VGLSiueXhgQWUrxZTgTR/vhiZN9PNcwlWBPsk21b9rHs68kn6T
ZL/OrFk3wb6eotjQXQLLUw6Dx+abALgYzV/Di7tGSqgThHWZrPmFolHQVB21ZpLhT/+OxKEuI0IV
f478MHuEvkJy1nDZW6y48k71qhdExZNWuFp7+/clyiFQrirZmKUahUlNUsBs3j60NVhRVQNz7j3u
j7W1z+0zLRYSxwpoN0DCTzQHmtDrdnsEnT05MSM7ZokUMN68pBI/wIAEIYNibK2d4cAotlklE4Bo
IqlBEcuPH+VUvbFzIlYsFqWMe/pf1SbXkWcFn+RvXhA2KT1vmofyNiSG1EpznjkBp+HBf1F9nSWq
7Wvspzl+XZ5uHrD0vQmdVe1jyQ4ggqP5VsNVScQePQVgKim83rVI439fqQ8MNR4BO2eFxUyqg7fB
9n2qMoAoYdOaCP6FjP3RLe/yyDdSuif2DqzMR+2X84TEEYZMo54heOMHDuCccDtxLSok6+Sm/s3V
loAQP5DKThLS1lSRfuWt9+Oa0E8f4gQ1AiQ8u0dRgUMzUGnwqEuhEFdBcXNCxz7XhDm5e5z4PvQh
b32/zCJE8gU4AcXJfR4z2LCMOcx5xkgN62YvMNLMiF/IcXGN59XWw+s6zTgij2O3mjm3RZpdPGNN
T6CGsY8LJFzH+PWutQcKiHqweJIBt+2/KjJeDvxBJePyHtYXcIUII9bw+/E6Tnehx4paKmgOb4Qk
jddAkqRlJJE/slXp0ngp9gWmO1mpTafR0O2I4Wy9RnRkzX+WD6oUUXvm/mFe9u/Si26MZVvO443l
6BtV3uoGIMt8c4zM95j6FW1HltQmJdSt4Qt4wMrynjtFYN6SB4CIzOEOegWrIpHwdEGRQ8tC70zM
0mvPUKGqjuK1nL+Gn8eP8Fn8L6CeKMEKlBCiowKE4q31pA6bCijvkoBq3kGjo5dxkeC4SasSR3WE
YjVoA5ib/6coc9YkpxMmBXLxGYG7jG4C9zOYmNv7b5QiAut8npz1WibDlyuNCOfRTckQGVVRqu6X
XU3XsHyuAsq2Rt8KJ3H7e5fifX0mCmXnS1nRqwtvY55dabblsTlcpGqJuMlWZ9nfrvhi/Jh0E2jr
GnsoFjfxMwT+Et1w5uNeB+DHVnF/dWyvIdlpSeg7xj7PW0QqnXkMKgjM/5PvdXFd0xKcNV/Zn+HE
dXX+p8helUfDvOAGgcPibj+BA2GWkyPi5wx3zoQ/XI5o9f63nM+0U8uStAIFiYv1gXkF63VwiyLJ
lcLt1gH5la3ytTD00oMVH8/ORe1XgM8m6kz4U4zW6YyOVTf7pE7I62KN3S+JFkU5w1o4qlnwU5uj
0ZQpCuxjYuaA6/0v/uocRM4Q6/FZobKqvV4l/tf0Fngo+cQNGxnQV8qcSiHgdBWcW82/ZaXL3SCf
EAYln5FcHoYH8OhZY13LsAC58/aMLprGravi9sCdjVuc5y5vWnvuwXbUfvLCwfYmp3WSwcEDoJ9P
h2l3D9su8GkqNF1AFOqPFGsmSTnSQSABA4JEpGa+gwpwevlmLanVS1MYzUXRN2s3KOSt81xyk32D
2WQgznqqMuF37BU+Eq8i/j1v2kHac00zUzlq4fdywCvDFvNYr0XOSmW0JY5qcQCeBN4ePmldztvo
4BC1+NhW23yR/8fypCf+ij60D/5/onpXGLr7D0vE18aB4IbNmK4xVezFR71drfVoWTrZg67QNihD
aoKvI4pEevqSYGM0jp+F+THwvskgle7y2+eEqr99o3+Aym0AHAQsF+UQfBinW5MjVuwD41MW8gtx
PaBsYQ/rHCn7BwxntgiJPVwFr7fL8MIJtaYaIA2yACWN+nPrr6zaLRzmdVETXV9Tb5C5Mbu7BvZV
zGOkZPNCeAZsICEL3sQwRQ5EwtciBPE7hXmwLm12kw4CqPPyU+e+fcViqouLn+dRiSVTUyNbg7TN
LGech4mMla7PFv2QG+73BT1slMYkNZnWrBGw/eU3ava9GJ4xIHqd880YQ5f4KantX4CO8tIM9qam
Gh0zTuaI3sTjNU0li1EyjGFG7oGyqGgKoBLMPuhZo107yWm4nvXVerJC38MHcWQJ+hR5N+LBtDSd
UdAE5Wff+asflx6woi/F4UNFZqekmI/JP7DSo3bDwrWN4ARsouytBp0v+6XmxyCWYCNqOfPSPoEN
J76+LvGQISB1miKwuzNYAlUBt9i8MERQlBywOmymrJ8JT04P5mWk7iNTWLeWsVspmTZaffdah0f5
CkHhFpgRfukzEfb9J7KUh7SsviNMAjWmdPB1gA54ZJRDusjx7cSz+DpwqT33VEamhtbLGoikXIDl
+oM+oHrW2D82prtH7L72D5IrdUMnDhL+EDOwA/iom/RVpB3Z84DUj3UFoUrvZ6AMmyd2ux9/khvB
LIjYKkSAI39Ks5AqUnv03r/EsEaCqdil44fk0dnALwBTMTVcNmzm8GGkzYnkmNNFSvtR2U9ekwIA
yzSYOH2j+951ZhHty4hhAF2pgj3UvOu0TmcWdR0D9HEhaGD2DPXz62CRcFHvKkuUfKkXrYGuYQAH
/EnjlaN+zkD1RTuwUmq6zxIrV6H4XCBSNlGxN0O7NeQNZWxZLn0mSpoS0JQziFUAz7dka5FmqbLZ
UBM31cUVT4cHpXZpU8GcNyFlWuPkzFEaHDHOzrYDCVSg7rKIny5fhi4xPksowOc7pngqJ+kjBnfP
F8p3Q5tmlwEXs3nfAzEzJTxB47b3JhKhArv/dbJVLunqTOunm4QddCzDSdmyy6f9XFsx4fFj4qC2
ef5P+6G7A32zT5wNobQUgI9JlUmAlFovJ7XXePzdblh+lejb4/JFgW2FqaKuM5CrCGncO26xQQvy
kznyoI6FlJcIF7XSM2vQjpmWfIdIlZSrTpUF4ejMPSrzBbaLytrYc8fXtvSLSdn+vvWdk6tuAZWT
iOJbEhvJDM9UPhKzuAJ/04pBl4wW0+IstQcOVFRUChOI2uJHpWG7CnP9noqKd8wNEpZ6bv/Mt3vD
onMiew==

`protect end_protected

