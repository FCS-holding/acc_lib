------------------------------------------------------------------------
----
---- This file has been generated the 2020/07/30 - 18:15:51.
---- This file can be used with modelsim tools.
---- This file is not synthesizable and does not target any FPGAs.
---- DRM HDK VERSION 4.2.1.0.
---- DRM VERSION 4.2.1.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=128)
`protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`protect key_block
f5Qen6UuzITB3MkaJadfTg1r5H1dLZUCaxllYoduzADNljJAbrGx2fhqgI1/D8KIh7/CT6YFL0A1
FZa0jTjsBjPtnWeltxVuiirD69wCeaezVwCC0dIp/3q0ufWEPMJcRf/lJLcpFxVnxlJmaOoO++hy
++VpQ/MbbFxypmJenLE=

`protect encoding=(enctype="base64", line_length=76, bytes=884816)
`protect data_method="aes128-cbc"
`protect data_block
5dn6A9JRoEyZlMtD/ZT4m394D+7B0tKkcREc7OUDMLgyhHj/zGrkbvg+WGcGL8Wsg1lQgGIRNyLD
kEYFfi1/UjQof3Hhb+KB7lJoOqoC3X/+Y2UcDYFovLDKXZqkvj+Wt9Oxyith7t4PB251o1YC57AY
3steAZwS8IE6OuqoGFrK7s1lbGoMW7uFUcgbiVQRI1t64zlyoeE/ZJ6eCoIvOsC3UkTTTb3JqvMb
+SMlEZlN1SjsvWDDUrF7rpqRtFM/80YlCXBpH/R3O7wq8w07FUWH0EiVvrMG//zba+WEqz6C5wlr
0PfmOcNGCxpdbGPl/yA27S1bJhfjP74CAFfLidCEIe4oRWQjToF++70Fl5xzR81rE+eVyLruuEFs
8Y4+/5NTH081q+bdFKP3m22ALatgg2yqbIDlIf5f2KOCNOkNDHREhotv2T4mLNQ9OBkpXJ0j6Ncb
DZa+wzj8+k5l6SKh3InpTcRr6vrPfnQ8FqT+ke83LwT0PpF0Yk6y+vUJ6I/uZBwUUTGXmCSaDznY
B0AMb6yTKBD/FycdJryaimS9hmtie9K5jYXTkfC0kquM5yEgtIHfavjNNfBdPqiDQZraUd4mqdxo
+QOPtXFmoOnT9/3ulI67Im8KxRbQNUSLYP9v7GXjCLZTjklW1f3K147Rffj9aoAvN5TNVaP+Ly6X
akIFQ7LqownponJcBoXXtsm/Z1Fmn5miKEMyDkN3NOyvLqvPSNn4p/pCbY7mJWKdr+gq313K+Saf
Ri/ZAm8U64hR6HMn+gsn9HvwA7SWRiqLE+AhLXRLVabCKQF6jFeYDosp990oRyUWxPS/44MKFtsg
ksb4gOqgpZXxo1yytbv2ly+PJmVciBNGEzfYP548o06XFCCnFvxTTmNWojXfFm8uXFDI0Bt8NDCd
qBYsqeHQ7Ce7mZrp65cQMgEGApERYLv/lTTbTdRlLYu9A/IcmTyR4BdAt507Fd5X8R1iW4QyLdUp
1e4CuTR0ZMFXpua6XxL2/AqasXvubJ8obK3JJCy+Q/9wtSFtZUf/216pJZ8/hvqR1aoRfWl4eN+C
+OmDkdeuOKQNl7DgLHIFAddIPEimo+wvfs0RyV+/lsZTe0h/eQ1AVdRzCg+PCK/DKOWD4GlZuqfy
C9tdmNjeRzMFIVsS/ZTDorxkqTqDO2IjBVamNkQGOmzGr32jphh+Bnoq4kKpCIf01Yb6wJ0Z8IJf
7Gh0mE+d94TuAVKtPUhIu9fmU9E45U3hWxF+emUakvxy0yAe+Eti3BNdWWsj4OO39Lyl3viupeMW
K7iF+7ncybCphG/TdEJWvsNfdcTeQCng3UJcItuLyJZAqJK3zGJDKa+JllPPUAPdeahWN9I13UeP
IQVs46HCfUtd/I3fs4Q7DTzG0Yn7ab+EkhaWBeLw/3CP0OszTCojWo5fn8+Q2n4doiaiI1vYBH4v
uF6tP4OkPqTCfs1nIm6pOAlyevIJh7mXC4gyBJI10pEeFOXpA3doZs+W+WWTCW7WiLMdhO64h5Q5
O8tSsJaZCzSI6ZjR2cAOGj0m6lU7xCBDhghY/DY6Z20n7DtXh5b9eavyt6uPCw9RMs3jbt/lEm7C
8DTO4YK4MPIJbJXN4yT38jfZKs1FbkX8HUtK+gWgpo2dq3ji7+TGhTHrEN57Fa9a3qGd2YnnWkJG
onIr+lwNhLWgriFY6UG1M6OtC14/O8MirHbxoV1KJDVKD3Arv3D+wbiOaR1dupPEVu2LHG9aGfMn
ARNbzxx9cBBJmTco+NqxSsaj4DkoAwP80Reu8DoKKuiQVWguwiJNiQor7NPKkRbZuI2d2Z1AUlNp
MWn2VulKD+CaBMEgjk53VEg7nw5LFzJNym7pJP4QJsZjwsoeLFOH03s+gqV6+eR9oPHhNjroPO+5
crJSAREsUeWl2YQpzH/neisBtmixkZYecrzoTM5JFJUFfGwxfQR35sSEVbKFk5Ce+SDw+B0icWWI
OxgFb0+9rYWXIM3faGvRHxCsx52CG2pKV8yyJS8rploWoNovj6cow92GMSi+JweOMZtdYR9yGAoS
LoHa49QSbGRKyJu93p44YveeKNSczVXyVJc2Dzim2C8W8WCmfDJY7WCgGha7WYETF9hJ9KtFztqs
0yyQAGy2U8cQGJqPYUFTrUCQ8MufJ85iSCCmkcQRFcDubuUv+v0+eoc0FrMMv2RQ/8PbzEr65V7r
vqtw2ElHFiNjR5jRqw7nFMImDeqTFromOwYsPjpPX/5agVck2p+AGr+zffItsRekr6srtQEeIGGs
HND2A1NXURdd/8yrtz8ijhg9d0RHB0GI9zuT+GNfj4HOcDO/xmyNhm3l83ax4x8/gI1UluffxC17
yKwE8PzCrD3s9F8O77Mx4qI8/65NVhBCroXzcq6HCSutDnU/tAQHHYnBnWy3LBWiI7zjNadcWtOV
TmpPTHSgc9eQ3HOmiIligUSw05wvJF9jhMbMaG1BCRWYNUN9T94b87Y5buRpbk6MiMOkPztMo+4c
FfF9W3POsDpXEdoRtLz+vCAI421d76tUO78LWuO0gBspZjITZZSMYOL+TtNCdl1ERxEje/dZ8uu7
tMsLqP/805Utw4ZeZ+1B6/Awdj+wi7A91JKdoSWlfLKZMfrVErY+/QnHmHjvedisTcqpqw+viRYH
O0A+H4afRrltl5Az6eALTS6DkMS3IgmFVKTkdjnemzXoKUZSmRhJFF3Jnxz02dBB17Y2T7irc9vt
V9wktDjy1ki3kw6AEMH9NhDBSN6tYB6sps/i8EpSUFmh7SVo419+BBiRW8w3DupX3h45VhOx+p33
abB5l6NFWuTx/PIadt4u9LsJo4ERK2D7Z0f2qbV0JbDfGeSk8ZMtKOet8koE3XDQEEReOEUPaJo4
k8DVxBH+kAr8XSkB6WSXS3Z/+MisoKZv9vk+DtO6nonkR1uZ8M/bXepD3wI6p7E27d0NJIanqJWg
Y4F+/J7eMNiQ1Tq0V3o/TaUYfYcS74w84EXBY2NG1uC807Of4li6yORJ0KTVbn8hUy7FSGa4eOW5
+IHGZ97R/K2LVeDWsd/WztkWwZ2uyIXCC33CpgGjZvIyXg7XiFYLdrd6UQaZyYZ0yVA9f9r3kAO6
cZSAG85ksTAh5wBbXi/0QfAF9nVKmhWmy1MxqLn2RxQD5yCISrzuyZwdTlltQWjMELTQwTNoeNSH
pVu6eiVFZG5gVeiFjFnEngInJleXaPyQH38yY3AC3FOmdG2lMHKJLjwgjbikvlIdnUPApPSqFh+a
gSfl5VFRdHoNO7iIEQZBfShUN1Juo4212fv1kArqhLGKlLAailPmXDEZcoLfoXCGUXVH0n9SdnIW
0GUD+9g8Pfg37vY5ic9C1O/YOw0jDrxy54IG6+ahOi6O0UUTsYqJEsvp2g/Hux+2eaU6x/fHJIVv
upMdIgYNlu98bRX7cLBYgNRG+VaVLXendyqxhS9jqBxnJbAvO96BUf1V+aIDPyCurxaLkm2+A0/p
0KkO51QQJtycN+sRGJqPo73/bjOAldlvkA/QekLWhr6G2FaKjXP/SmJ4E1fONOs/jCTBpfm1/8j7
HN7rjDhrXumo5igKjh+7bLwk6XhaGxvPPoYSN/thjKWZ+I+zqO+x6ytQO7Psfh2a2rZWR1wn7y6P
JB+fqDrSeNFzXCftqmSCu49kIxjsDSDQUrQQJknfVcdG7tfvb+nus7XF3P6RhRvETKYwGENAt1xv
yjS1EgfVL/jLSQWsue70G1cNWJNhseicFAhUes90i1MOxLimnmxFj04Idub849reuW3VHWsR0mxR
bHgLctXigUaCvqok6voqe07S2isQxQ7rsei6p8MOGG8cGU6oVfQFtgckrd/nMdTaQhkEZKueVu47
+gi/fClqTX88dH2KBKzE+9NGe9aihZ77g1oaiFjAig9MNz6UcfUx3gCUjifoxIc0GAPu7R1ijpC2
tH66H9lkH9Wg4R3rIdSosPrJ3uNVO8XENZ4xLRV8gSzQ83nxKBIgkxkLwDKJzsNYXVgDvdlL1sGg
Q8+ZFoOjuLNdzXpU7Ff03dAA09aiSGMGG3+58R6Dc4auta78GtnKsmlHuzoJDOQRn3/Mpbm29RRt
hLEmxpbNvNlV6wCwUeB20m9JOZV8dub66eRYyX6ri+RGTbPJadp5tKkK5dDC5K5rc1uUMzVTxYS1
jdM5IJ2LLc9y1mhPTdQDmJJR9eAyFKVOCizSojzcfOStO2ngMkC9Ce3F5s945ZiuLIkcrobzU0Ar
gE1mHZQx8I9NKPNtWQXVx3LPy7EQ5GW+LWW5Wam1LIWlcAVoV4n3e7GiYQR0E/+RFV8iEDnyFoy0
ddRVZo3T7E978WStLjcDc2KAzFSXwD5rRRAxyvt8fSkgZREk8gakkpH3SpZJ+spfXdUP5dwI4jg2
CZ6DlY0N25gooGtc8Hco/LWHLmBRIL0Vv7WTzfDkycBBT+jjZdHOYJK9jEUi2Kx6E2uouO2z1yVA
X/zUwvcncCWkMPSgIZrNhn0h24jDNm8NMUzRrfQfOgVzOfZP3SjMPLhoabyjmi+RKNPOUl+PuYmJ
59xmi70B3tg1npAdcYcXGWQ+dKax1ihk4aF0cxVGDrDfeBhzlNr1W5/tr0aZRYw+o5DxNzg293YB
oxQNLuKxjaeEC2M/iEgT5WgG92oHnSmyNTDZ9pgnSvjdDFP7DYsEMHwl+jZ7QTQHdH1zUcbf6FlI
wJcINwW39Pcj+kyJpXzaXNWMUFG7seftx3ngpMN4VA+RYBnNEyxvW1LGMPelhdIi7Eio8cBAVi6I
R97FEsye4z0n7r0Gs/17W9NNQBLo3HlU7zQt40GBhwE+8aybN7bssIFybDTQ0I0osjdgTe57CrfB
pdTxFItEMsylGkqAXlkgfNN4MAwUCpy2vSiicNz+BiX86q91RAqXYQwBAwlRH46Oq7Seu3c1BqLJ
FKAVrwWAUgoRw+1Mj3yX0UBZq2EgYKrVorjWWE3rpmDgV7BSAmw4MGPDtwG4HGHah6EfzAkM+dtT
BOPZi46AhTOp+PAVasAkO7XAIVHpYMbRhi+r0fFno+wxx88LMmO7nNspt0MokGomNhvD3eu/dFKq
e5Qb1innIfif7a1SdYhWswGkJIaQCAloVXiQU6ab+zmJHteKZgmkpTBcq/1fdYn6mp6BSplLVr5M
EizgAGH228rHgJbrsT3MU/Nv1P0LKA3nsiL/hAydr41w8zyaDkX/T88w9XAlDVoVyhgK3oRuBTNd
Cpyk9YDLDdM81ryFhgfom3WklOzoS1hH/uiw+CBHAWzbulZlyu3I+19lHmfJIXJTujP5oW9eplcZ
RK/uWG+Z6dbvdQaBBTo81YP1gh3DL9hqI3H4wFX8XlkXADSs25o0Vpkx2ctNGhMxVyKcOaBHdaLF
HIrxj9GdBAVuzD6muxo+65s8FMU/4gED4t9iiR7iDiIH48rxcsg5rtGBbAsMQpCY5ECur9iCfLSQ
ayPr6ZuTBIIqGI4MaHJf+4a893PLL9pnqNUtwLXGzEXVoGUVkxbhJM0XZ6TrfZ7XhaGGUO9H/qoN
91MFff8qHJwqJJF0lYR6GGk86jQY+12dmuxYe0Y04zU9emOLcCWqNPeA/rFJsHc38FbzUELtinDu
LwaSbZiJCO23kH9v0p6zyLExNHYSpio5v56z8+HPusV0WSyC3DsYzbB0PNypHpYbfDUSsSK3Ift5
21hzQi7iHyTQmKCF6NLVXB6yIeg92VgKBWxbpkvlaREpbJFxcrEfA+8noz9MAH6HmrWgVGHy7rEY
L6+dV7C7GUdsHOEtm2wWRNbumcWPZFb2OTxloyeKL8CnKeVNzmuv/9wMsUzj5YGYDu7guNyS+PSQ
rLuC8uOOsKzXPyDRv4ldB/2zVQC2ArxoY8U+Ng1rCdEKi2maB4dvUV4Gbkn1oiYO3zA+8q9CMOHr
2YWaiCqqiRrVOrtHbgEnzmRjNvn4G9w4WQTG9u8bRdRQiR5ZlB4NqC1LuXT41gUx7JyTElSewKRd
TKDZAn6MlXL2o2cQizwsdcSqkX19Se1viT84N9bK7oWbWTGQ48S1dLjrjpATGv2GF5Zqe56irxoF
q0ZvBjEW8Sy6tU0FOIz+AIopVI3AyFQWlqTPgeMIHs2gTcBrp0+nKhrZy0XLZrtthZe1ZRyKzrtR
+lNbwzmx9XA0+GUN3GT2aLYj/3mS26wfrWm5Zp9YcO3sm4bxQhddp5DCCNvmSURgwcEQ64F1m0sW
IHJzzKs5MnyAN21RveW1OUYQDQ+TmV4O/tboPAJ6ZwYlxiXKfh1dzQaBB1R8f6EdbdWbIGCfSGdn
g30szyU54Ny8uSlQYpNU1HliXdMn15nT7oLd8FHd/CBcAccLVykKbU6HPyF5bEl2yKhTI6UICsnl
InlIDp6xTF5b6ypoHiYr1b5vFNUlgBvlWHHgd2tNDdLDi1SPItfhxdHWdgAeEviIHrZJhaeB3eZf
SitiBOSazcxj7tOqUqwuYKUHUZMeDyvmbbscSkGywPp6pi3uR9tAg2xHYKS07bx57bw9rQ+D1rhS
MYiqyNblkBG4V4fs92jYxC2kSO2iTicjTbg5RernQQLDXjlJPPyg/B9DIxC7MpdNYRO/mQS880ao
x91RrrmXMeZuurN5SGVt2NqbF+4wSkKP8fac08bQTmCBhoFhVQqJ64R4301TxavhNHHLsfHT1lCi
PbIyPxYY2i308ois8vOVINF2BwaOPkvccFazMcPFfcDI/FeeD+EtD0DqHjJnEtxfPdI7j5QEwp0O
jg5R3sYbh0F/SRAog/AFAp+am4uAx0KZ1mdEgHGnNGwGdHPSgVyjbmi55igCQfREBkufPLk1CvH/
jUFvKVOniv8VY8sQgbvgVsRY2ZlpuFTML4VKtHl9nYLsQf+WSCjAV9QoEghSg0A6vsSCl5zwJp9C
va/tjGj+fGU1Yhrv+vsQ2AAkq3GPu/s7zDXljKwNqv351UKaqotwFUr3IJzLh8TzbpeZ+T0lzuWB
UOjODyjr+MT67F1FGI2Yjt6i3tOr0lXV0q/R68P+XxNEK0fddPwTnQBh17aDaHedz024j+BSeZDK
YkyCjA6GJBTzrDfB2Cy1MpcTsDygmcsZnIrjaWT3ABsrHMuGZ+ikUZ2i46FbfaLIU+SzG8DmE8uv
MMkcxIigB/3qEwrPJfq3bAMVmGOoZ8ogifPOMzEmQdCt9v7hD3ja9msnPbrV/BHrAVLCkXFRkuDw
QzJ+hLvBrGN2MestH0eHahGpvCtejOpJqYXh57p5YvePRlyLgSuPOlm8CUxyLEwid6SLBr9d9Jtu
KcRoSUvLSoptoht50QNkE+n4QxjelHy1y60d1XyZqYWuEX4JWquLaVOseaB4z+50MYGvbKlx/6dQ
4mje9F2RcubeUZR/O3CC1bFSdG6TRp3NVXCgQM3vXixjLPZ9lUry+Kz+Ssk4PccWqxkIWDL6NFXk
+ov7wL4FtynyudEIRtUK1DDBWXOOD5/G+BPx7AQ1sDVMtG/H0bAJ/2xAAl4Qzv7O3XZ+kkkdreq2
t3clcicCBsvto6XpeE/cbH66OMmM1gh/IbJfhEQ1n4RMX9oZr58MUEHy2onIbQugpVlcStv0ygow
10nQNISFdMY0YYXwRFfP02vjSXB/bPYnYiecPXbEQ6NIYVGCR9eHup/zDArDQDbIL0AUyHM6F3hB
Xj4JIp2VzvAUhu7OCCxMjAWbzrkHnn1EgVVp/kZxX4Pk9a5CMgyaLygXhJ89kh+g+UhOE55DQfOR
Zim65uOp9Jau3nhqdlxs+W3DFCuxTMUOdygbq93D/e4TkxkaF1eD52cKTyKP5tS2CEJ8+YjLSat6
5flZScyjUYUNN4V/UE8+c17VNHoWf5wwOj7/Bp1P2EERP1Pw3y+hxtr7OgzvCqFhPIohCnRj4kNg
Dfs8+FS4HEX+shDRwIdus6nqy0tGu8B+J6QlT1ugP9rK4yA3WlZQA0WrDh5oGtJb7eWnLjihY2Hm
AQ3mHhjfKMqi0oHVCxluR4j1xcxKooEcZ90aJmMir0Q84oef3DCF6Vi/UlAuCU2kK9ly1bQ5PwPC
WGk8iyXuNu6qlbeG/sbecEWoYJkaaQ8907nj4t8CAZzlKl+frQlb8wU6Gprzmt+vxHlTFcdndqgJ
/8W7dAr32aNEG+rgiETGqSOfCUnUVXKR1QZj7elowvMiVKyB0h5d4LvGGe7khRGzP9CEB7AEGbI8
yRUaVuR+QtIc1fuVWPfeROBD3S9HDqYlRIVa6a4q0patAGDEUp/1WB1L9fsw0EptDk0z0BiryXCh
Ku5lJUyodhTinAViPWXfpxGWaN5vm9qTz7gtYKiMieTHm6LpbHPBbQJxzh5VfRQrbijPB1EtzaLW
el5TRwVNfsurax9G1tWY7A3FzXgXs7NC7Xv6NkNZJmEvfhmtlCXrEL2ncGBOtQwUb6A2XniBUyTm
2zPT19XDqF/xFB6wHWJ2poPmM2C6MqcDf7q0KnJSD+98OHOGd5TaAvnpAtu71FzrOeQKHSkt8r4B
Pq8r0pDzYkoYkwVt2jPYPhkzBg9UX4plxkmvVkn9IUgT6UJ0nZ3YktLyATL5zJfguC5Oa52HndHa
gdaQh4FYCp3SZgCk1NhBrXKGjQE7exQ1Ks6g09/j98HR3cuQsw82QwnbsFDth/4dtVB0sD5r6827
QSmg6yFG+KoT722BL3FYoP6OLY0rRG9qmU/QkVuZYPA3Wzd3d4U8QuVWUbb3W8/axUPaQwSml1kR
PHlzmw6iCfNAIxSM4Dr/9AImvBhoWZGLoPeuEAxC6DrfTscvU6pEobtSUFN67yOkPj7I17hYL6IX
GfogWbTYJ2D/gV3RJVmZvScBqKejZyy0uWg8De5ZKgLTWdHb+DD/xzknfWwnstMoG1Oyr1Fb2+Q/
/mddQ9ndKcHY0qbpux12OhlCts/1iLKydWgWQmeSI8Ww4tneQNFVSlzrFmYfhlWonDdcOP2P+IAg
1+51c+k/aYTzbPwB6KPGhF9cExtEXRC2HVpGNdsxRFWW0XyMctFIbA6+UxnKejWdai3iKpTnUYaD
sfWvbQtC02kJZ0tg62NZ5uY7HQWnPgEDhYCgwj0znuTVPTMJronlZ9aRYFvmTXhQUW3GUdR9Hq+R
THqETomkZWIHQ4SvGNoFpcDKBXZIQfnMvA+E5gw1xIIjpk75mCSECJhD74tuRped7dIp5cQBF6+o
OhxKl1oCnTySUWN3Xz+gKWm0+Wk8wAYEGsrhEbUShm1dgoCqJk22F+79rb08uIDZ6vd3QPUPFaxm
IU8kkn2P8k/Xg/11EV4v4fAnmXZC77CzNkNhgt60xqLBmTJHfKYdiXQ9/ZXe2W4bOj4UOjIrwcPR
Q3beBjvWQ4dM4hhRVWH1b4Z6D8Djlml2zICCgPULdI+XddVVMSG4vDs3XkUki5mu2soyc9XuFSZd
Uaak9xATXDexZR0rHGi9TynwI5PdqwOSttjZiWrc1wY98zNSH/iZ6F61dbSiTNbKe97sppNtrIsO
LHatSK5RSK4aV3iTQvjkN7caYbuvK1PeGIcKmR3+4+XvBw6eb6g9wJqoDGJW0DkeobdxYkEVwR6F
zynXEZdLAlaycfLF9SZxmCRtBknyx92eCl9405Gx85K64yJ3Iw+JsjdszfDyI64awyi8UevJn4RH
qGc0fDWvXLb4D4uZ8NaM5dkot3Euce3IbzCfmlHExRuvV3t011p7MlLMDiud1Sv1ZYdcv1sx9KMh
Pd7T6sBs9tIdf2mohZb1k31VR38daR5B8HiW0aPxoLn7wQsnMbTZC/6tTwlR//a2+TX3xEW/FzsY
sZo/Mlhpd2U9622XfzO73rbYz71YZgJw1LYKO6u3OqmRTZFIPNyrRnTwdcD681ncHstJgpoM1Zu3
TPUYeMOWjCtLnRzcQZfnAbChCb6l+iXJyDdYA93n9+JMOUrqtgLrT8WbJf1E8Utic1sXQT10OAMu
KVP+Zh+LT7Q8Qm22xUl1KDxkqfBT8AYOBIluPF4imkjeXY1OAxqpjocxkd7rZ+HuzZSBqR8yfIgq
LVlPLX15aHbDQ0Bn+xeoI3VIcBl4n7o5TlRaLTPH0ki205eH1B5s4u2f0xRz/OMnO+ZM05r4to01
mt/G88x2SfCenlnUT0WWbrkGrs6KEp6TXruXVlZHHNpY+G46YSh3I74Q/DsJIUdWrr5w/bkzx6CU
OZnmQ870zpT2cfnzGSAVMqyn4M9f4SkvQPpU9IR6msmhNmoBtkD9MAbgtXQiRqQXkWPEnHB2PKQc
rAZtCjeCb4qV30pZTxYOS+0Kj8PuSBoWf6rcRQHFXhhyS1nhecrvcWPTFADrcmd6PJ4o+OOJnzQ8
aRMSNGVMfHrV8JooHHlKNkkWtSJ1R+Q6tRrES6AcgGZl4z6dtHIClglU4r17s5qQic6gHhJbAFGk
jqiI4tLqM8+3pbeLxLYS1EFjsjGv/zOC1Rw9SWz9DYpSpz2BBtcdfe9SvDKfLMYhaFGncqXCtrb2
78+/g3g7qoFyq8RPmHboCHKu0ljWNP7QTBt+KdE+wPVh8H59qjXycQX3VF+GRl3xLtiTpmjFnI6p
VwEbAn4Tk9ZFFDZp0d10zF81YeWOFq2SveBMrnHbxtJhoyMD3ToWqCUAx7Da1OMaFlk8RDQK4iF0
x/4KruCye/zTqWoVDOZv5TmM7YRrZL8nGtJEqwoMdmeAStA8VbbgmdSmw0efOgTyRTeNKW5d1+/8
VBXiCATOaZKbOfx+Db58r4NlAgdTmnEqbDPcFX8QQP3qi8Y1yToOxcIy3pmfP96sPweUe825+aTp
BVFc4XgbAJq67AXCzOEgEZ3dHhMrbAW2mBgwyqmgjmZRzOekrKzsMB6S7f54Dhz/xun3079zDP0C
5mLxmr0ocuu9KjDGl2eywKziGUZd6jizH+iuq0Y2LgwiZ9gwGR+GjWWxLL55xomIx+vbGqbH3giB
vDLwXKPzbtel3dZnp1GUt9UANqoS37HX+WPcWDVjoBBlb5Bl0XEXvV45LaeEyF4hB1iUAcSVWel2
lTbViUUVaIXpJwYCIxmf5zesbCEJq1B+HbgavlNQbycAHK4AMOi6CNfDW5BxELsRc+yl0NYkNhKA
PXq5vFan7AWZ0Uj4Qu/gFwJaDs/WSlzbhkRCh4baXgBJIIsjAaNnd2NRJPsFx7MUEq/UA8j0Ufp6
MNgOsHh/nGH4uzQ5ZoP4MaRkE4OAv6gK0VQ3mEOQw9huyYXE+i6ZTv//bs+UzlG9Gbs12Vcvf5I1
tKJzS8VGZr9PTpEkRZT92/BfgFtF9zyB+bZIzYlPUjcceUPOF6PHXpisfquOJspvW2jIcRS+Co4B
tmV0kORwKMkChThyRhBxAoQOlLkQylw1FmwMF0CXyZq/tkagija1D+rmYIX7/HHjacPXKPUViIcn
9S98nQmyqpFkimJbz9E4pe24zAHr2z/nGhmFDEXDgnW0x9RacMC2YXDNUIzQO2YZatJzX9GIK8j4
EaFZ+GrRIiMs9StB2EseEVc2/JlGr7hXQuGiV0TJtRfbAon1uBFD7GNWVtcf2RaLz6uv7VSbnlur
C86+oIJwgkWt0DnUzjpnmYDwIBmRdQvUTFkXAn9QK8VqDcjZJCIwkf8FBfCdEnR1AdTCvN87DVCi
oAKG9m3C0WMwyiKtaNnBvwyL2qI1awIaF1Z1gHR4J4PKudbd9S4NkFTDxCF3gD+6g99GvejiSd6k
MYe6RPJuOq2hS+HCsNyG7f+snJLwJZZzZd7E1iM8os7i4BsVOffjE64hXxE1Ny0Zqx+rO+DDHbvr
iDiJchnR2Z3sdOb5IpmWFCBPe9MNQdoUuB1zbFRI2pUGP5WMF7uaIVD64DW9cEqLQPeV3wCctqGW
dkNMs6GJsndWEcM8c7QwHZFWhN+yE1xiO7gi9Rine5LLeigj6sNhyHrDJ2/5ooZ81lHFel3im8/v
7WfmJpuxWVEBFfvk7Box+Wf4/J43GuzbMaz3Hckhd8HC/E6QnmKN6t8UX4E01mNGmM+neADa7Yq9
mJz1VsKXRkkLTJEceos3NK6YHtZY8Z2ZfEsP4B1Mzc+oRlol1DB2QccnW3tCEO93Zk13xXEBatrm
IvTRIJBjr8BIAtbd3cKhetiYLE62kk+KGOLizTacw1bQeVNq52/Ga/kI4cOExvn3hW4KYknIICzf
cW6MIOFOvqsrGmdxN3tUp/6HOyQ43/1c98pRG+2lcsXCMTo76niwXgzByys2fLBtK6qAnxG/t+/9
IpL9v3euNfBOLzlvgi6kSEYCYYlpt6BfehKEqd0/yNE5kur+d8fy8WHN4I3Ev4tjYM9E+P5MpU4S
SHfamvn5M57uoJ8UzHuzPEZfBaSPWKw7XnzjFz3RKOP46K3wnCBNGv4qdGwPHKlWXkjL+h6uISca
YuR90yTJzy+PaYU5Q/QOtHxFuiG/qZFfvKI+k5ocIeztcOhALDD0Shf2JaSE2W/hRxVVhdH18wgf
R088W0m+obNJpK1kypv3iLDRfrNwoYwxfYpVmL2EGi8XJvu+kO3WTho2RLayqR6UeI8473U0NPdZ
6TskCWwo+9/jA12lljU24Y6bO2trCpuVkQquOr3B5Fs3w8WTDQcnPpU44FP7Su3JYKtnzIOhAh5Y
An1Tmu1Msei9ZYnzr7uApdazpxeGh8+xZ9qi2MC2Mo5TFE6Vy7VDaUyVYt1elCWBvLg1OIaoFfWH
fnuUCoWOVILseLm5uP3fOyy3EEE76JSRTN0X4+iIFZBG+Cbp11V8/JS7y2pQ/kJ+gVgBZlt2YWpq
078vHDnG9E2ZJxZtsWu7LXB6Q0UAMllUfK+FvYpJt1jJBf7qN/Xg6Lb4XElRAK9uoP3qoX4OtaxW
WLue8fCNWQLgC96ab1vw5cqjDCVoApQt5MM09aXYV2111rdysebUfpJZlaB9w8KdvWwHDEKNoclb
3DWjSxbwBxsvei6lrPe8q6VVPB4H86W8qwpL5oJNpoxDeSOwHezPjrGKqxvrkNgvxEDQg7CVMQx5
RvbTHDNYO1VB6n/v2u1up7BUXloeMq0RDkd4cJYdxbBmhZisOfMqFR5olgLjIy1K7HQUaA0Wxv2x
WjYUfcCxZEv6olW/d4ar6qu0o1e05A/p8PuPfqrbMLCPeQ7vv7f3p+7/RcMWiUhsFzSito/nfbyv
52N05+pGuGsWZ/m6dSr9JRCAYpgaVCkWZBtR3F/cuDqEzEqydKITUCzEExiRBf2i6A6i7x62tvS3
VVCKkxbCsnfOGDUA2M36FbTkTpd2vglc8C39ag3DY6IeDfQo35/GUgtaYXSWx0I/kbL//gHCnkiZ
tinnWwhJfside2yQv9ohXPDmSh680HA/0aKzzd82CkGvGmB/ezPLEoDx7kCiHWG5/FnkU4+xsKg/
3g3GCLTMfEn0zsAOsP5WKf30MJXT2PRJ20nqiN8gDe30Pcx3Rf3DjJdxgA2YH7zBz6XVI7HjeVKG
rAK9UAcKe7vVIeDNV1tWaj+akVR8G9fCrr8GPI39WPmtOWBV7wYNlqKMBdndqipIVC2JbE5TMzML
agKH5EM16lRDCg+BJQN4lMBy7U3hr2rNM0QRIdBDezDdY4xwQ3N63Otc7QmbcZz2ZeWF7dOVK3n9
fv86xn6pcMC03U2meNOzEb/LYW3dNGrTBSxBw845FTahnlpuxuMdRIeGeytnzVLtdHrD1H3Zw9EB
pf12EnNNIpiG8WocahpimQsQU3USnsm7H4gSiZFIgoLRjpn+fIOfk+hKhYTahnTJMy0W3UtiA1B0
21F0hgGIGYLloa3dg+O8gPI57AjRsi3+nK3eCPQc/tEPgxmRDKUFLkr9ci5i5LWwwkaQ9hCHGZOZ
Oq8gTVVjOaqJFdxEIcVMCOtAvVHk1SJRH6CoOT27mFlzOiCXEqw86ITi6fynKHBWoVBwuHrceC5F
cEJNAlQLniUfXHjf0vMS5DrYpW7obveknq0/ApLFiUbfl/Q1JcF31l5azGScSlMn03Mkv5nM0wKO
kp0crDZ+ZeHdsSCU+gZUYlr5qiofpT/i9UKqAsN9EVZ1s4Z62PeO92FeQHTT4TPYAnw1l+cXccmL
gRZdofMa9bQtH8V+Gg5ViLIBhwGXG4nRDCENdWM53Ty8JKkJE9jBRADjH61eqMqzKTwwplVoYDDb
QYrHrVm/r7JkPqxK6qGroV5E+yZGypbX0jp/fgL6bz1yid7Jby3VoMbYdNSq9/kAOFDPh4EuHjVK
+CEFSo01+HTOyD/gWP2ik+Eeu4qAZ2F3s9VZ/Grrd1FibRC0XVFKdEv18hU8+bPqtk1Du/K9XRYY
/uN1YWeVm+aJOd3o245nc9PIutQ8p4sE9OC+FbcdX/zo3Ec23Bd0DL0Kgdw/x/BvfcvET3Bib0/W
Tsn6TnviZCZ+VX9YrayZlTjvN47UYnwBzs0nxYGZQ5RVvhbaQ4Tdjq8M2CxyAahAyG9XpTtJF9fx
G4/X+X3U4oH1MW2kXiQDDDG4AGaIrAoR9M7IgPRhsoDui782EXmdpx6DqKByAVCYXEXX3+TW+maT
RP2FNp2DdW2DjTIR8tJkPsjnzX4qKydLdtGx2IIW1TT7P5cALw2L8zktb3vRqWjOkg7xi/+ePBeI
aiFtZsFEXzN/jtaQlSAmGW1t1jEg1f7ynmYhqrYjp7cdzkUUUaW6gICk7Sn1F1aBx/9+6PCVHgd9
Y67aFd1VNLC51QoFRPfyuzwaSM3XLSohLoy41DoLdXpN8jZoQnBuoel8YcoXDFNcvN/022N9EnM7
ixFZiK+4EnoMhORZ0D/0DUMd5QlbqI/HHKQfsoiVXCyGeAddjT4n6hD4/OEOv0rSzTlrtWjD9P4/
ZJY13Wf4LACB/DqoUmJu81wWt7DerlVNwmk2j90O5moWC8QhBwYW7o3Ls4nXGK2YO4UtaiCKsmhg
T9dc0tjcTJ7N1AibC9tckx8B+myUOk0rDNhr9hroG+BxUo1fFzCfvpLjHEGtCHOmXYWMa9BxAuEf
XzWBvfzsEuJeRbcnBPmCFe9jGvbvV+gJZ+9TUiHaMJFuB/yXFHjS7TpFu3juaujmfebfhT6FGuLa
g7m8gNCxywfQkh+ssX4BNwy3qCZZ6YfpMvPlpa7bWEw9oxSgVF14jgvJiXCRT77AFE6NGniDfgDA
9smlsuP8RQJ45PF0tot8P3Q97II9xAUQjAjymbryYEAwmDzAiSRhQZSM8TnVkkogMeDMUOqbQ1hN
nWoN+mAABCxBBl86y85dcEgyo5mjQHDYSdpXwi36ZJPopgU6rzZ8x4k3q4PylM62gSzJZznPGsu4
7XYc9iuatppxBNbKA7Qeg1eHAxs+8Nwbtrpgb5wLrqI2RBLmq3Dff9p74WCeh+l+csWDJmDXubyK
pcTL4I9COUAfj+5Y9RYTQ8Tp4b7WvXgnNKizfJqpiS/honChEFCTZ5UAYCRtt+pV4xNCWTI+q/bM
v1u117kppxCUrHOUHH5gfvZEb/Co2DGwur8cPILNPMKA8R+z0MZkMnJojrE0sDJfujCXgwlqZNkw
VlpXooCdPfIwYVTjq86+sL86p7t0TPPmFw5i2QauXHcn9dyRuxq5noyJdfyYwsP9r/C5iTsaebI3
AElGN0TuOSHdZu+pA3J10aNd5k1HRgzDLpMmlhjrICGNf0Eglzh0pBIN4MOLvekvh1nf/Cbp0sjF
OBANG9ZRbXjpxGgF5x7uz+jqROx27WjtnoY+IVDqKuWqVMQxCnCWmeeMmOM1uM/4AFuhMy8tq1+7
6Ioe/gnQAK368ki7LCdOaVMi+3qVTeQvfSmeLJP0vc70MI9OG5KK8CAA00gPzKuq2whn7kiuCrg+
hIu5o5HOWpKcRfy3nybL3M5tVkn0E8Q2i4nxm2KioGEIdNdOPKHYfd84uqYQjyW9k6kUTx+BdIE0
1nBTbTavMvkQaZc6GFZqpb7F3lGNcVhvNUycddkwCmYq0ZmPt2fjSB3I4ENQxOEeIEXdK4fembL3
31GRQuKwsnNCkR8bL2LdiDHh/MxZE8uW7O4fgpan0mNzOEQ+4yZgAiiZqq6N86g4lFJ2dz7TJDLl
BW9o0rvpDw4SXKXqcY9pUgaWABlMmNXvblfM6A/YrCOzpPk8X4f0yXEgdAQE63gGwHAd5u32f/n3
/g43NEfOMp2Uu52beM/TJ1zDrtQNGA4BkKSD1S1YByoTwZjAfFkJ0a7fiKNTcsjiv3iRx4j+JG8N
6hQRw2sy2Kw+qfkcfxDKhvqHA2pFFHg/LjoudnROkwKM2EzoUtfwCR2TDR9qPaG2oO3mJ83F4FmV
g3+XwzZssHD1vsro5lDtwphV2gkqiyLwSsj5jC+JnTn8pDcuMTpuuBh9yZT/S0IOgMuqU21rc2t/
ngjiKJbgRoIdBaOJS7R4/VGetPxjOgH/Me49E0V8/fT16CseIJlpckn3t7rNwf7/RCDNpDwm0zNc
NpzBtaPOAC3G1wS1539Z37+4NOKqzxr8gS1gUQ9gt52hYsMmHGV5MbERL5dU6LlHxv3pdzP9QA/E
e81GGUuGrH+VbdLD3tPnFWisUlV871pQ0jRu52J9DdkUbjke2SwYhQ31zwsAqdmOtbH2gOzYDx6L
OwnIIAkgTnHroijwMwhL533X+4tHtyYsNnZaYGW4JYdYK+jrInQdHh2TlYTt4jE2hTEZnMM/iOlB
bIJzFO7nsK+lzAbCs2VYRnu+8Eoa3OhNkFC6oFYrrucS3PrNPtOS45GfxjJ2gImSWCbX87BYoErI
Z4shSDPq6/FUC58k0kWhAzYTZFWgdsz8nUjrHolt68cd8yRcieyquEEsAUG8Wp5R8G/5aitzOsBM
AwOkZvWTOOIIASttFw5LZ0r5ELuaO3dtac9RKs1Ep1vpmnS6Gb0zB4FQwdEm2hiVYxpxAxYeSA5I
KCJDcoAmOUejrFfQRUSEbHqKvo8iYO+EZO9wRrcrvO7URbEUnw1zdKcpHq4DVFlU42jHjiEjOWZw
uZc6qo+IGbbJ9y6zQUlMzj+bYNaXCHr0jLL7p3fcX0de3Hx6I2650iLbe2A18J73W0Fjv3WGuqnV
yOUNYOeFkUi/wRKXJAvahhELHf5TzEiT16nAObZpJgDcG43e/V4Apkzo+TM17gn7PAfEFn/Zjpfs
Kvs+ElRSjk52ZOGLs8Li6DCxrwWc+09bIGcMybBFTAQc3tu4+qrwYJAuiwlB2zSg1ouyaO2clhhn
ku3u0plSGAjrgsbdN2L6r4RsWVh/6/3uDVziMviA+CCGnnQsqzxTA9RezTKq3RAnc2MdD4DOCNK8
8FPzikudsHZPFrCYEz22wodc99bGxPy+6HS+eJNlH744NQodd75hhL2Bj9k2xtDibT0JEtSxqgkM
PrLIELh/4/UYRQ+TXQOnqn+5KM5K6iVAxeC1Vrl+Qe4RNGVyjuKrvJ2x9U5C3jvNzYCMwz1nN9fh
1nm7Ufy6c8iWpNYSA09OxuIOjkf2L9YkUbiLwdQCRL+dR8S3/+JeZmCSrQP+mq1HAsZreNjd8skO
VT0c9QyBA9rndB40ODegbtG3OiPMa4pUWzkmfQBXy626+UM4s7MvXIZ8wh73hJ/vErtLOt7uVVM0
3Up3jGI8lqL6WoaKJXFlIOrLEv5VAaAVEidcTVu8jGwFt5mDYpPt91uOMzGlTLMz40XCSV380Fl2
W186dghLIcfnhp0hhAmHKntNNRR7sQiFKeP3tnL3n/aShg97jM4JS8p0yObWkZIQw3Pdvgv541yy
PAyuZ/7OIpqgoPGG/GpknPWMJPDf+4qQic87dGSZ7Ez/mwIcCAlWjKEHOC4TBtf9Ha9XsSWHk2Hv
Qn2yKzs0O9cPN6arx9+ydZWrZN868qodQkKH0IFd13pTQKavkYBzrLB401BVOO/FgboWdRNNczd2
+7UKugvzgtj1VvGO7s7TyPLBIplJUe2EsVeR8HAb+Zmd+5em/u2fVA/N9389gqo+sQjufnxrQSpe
+JSdKM2vGqhKIBphR3O2GUBaFj5XCSrAgoSeyUiWiipebS8r/uLrLa8Ai/yGQsj5GsBdw09vL/jK
HQPCw2qLlGuFL91cOgWDpCr2RQfkEeZ3rV2tfY+WXRP841nBx2wZPzBCkiUSO5UZgpnfX7LK0ZEC
0voiZF1f01NQJMZ95QpPI7vxcrQ1aEQ+2uf0G9i+NA9fDaTjh0Pn8KcLnGV6sf0FmXoXKKtP8Tgb
p6DlPsUH9xuKLUq9+OcK0ZatUvsQXRuQtxzcxg2c9zk1MEaMCYOFHntQiBDWR9ANjIx5m1jv0nE1
czcvbDFe9jPW/XZNXFMKXFMJV7VUCrDiGcM6zfJwi04MogRRl9DHV0IBrue7Nl1cFLKFSisQWNr2
LS5DW8wF0/Siy8bbQijdZlJQUIDOOwJbHk7UZFgJA3FHZITZTnrJznBVU5OGo3Aq84fnzu6TFjf9
Flg7jjG5ND6yXLooxI392EtFw05DZbkAbhlW+y1/zKj1a0wY5UOno9xNJsm7+/QLBpKsdhUVZ/mb
ngsyME6A5mXbBMT9dVSSf/8ZhK538fXhya7c+y6v3ZkvIZ7Tq57BITv9+aChC7FmHmLCAhngizTe
Nwp2XDUYNKUW49xzU/LWnR6qaJ/9SLk2GEazbd0dRe0kqNiL4I6EV6B1ZfYWzTAQ1vKCjKyL7mwA
SecGLjYjj09h2SObVQ+iWXgbuL6SkK9QZucMhuiYQne8+pXNXUXKv90h0myJN5y04WftgIAjhmzz
PA3pHkvgV69zd5ICkP7tgZ1AqW6iS420G2Ly7biHB5kGo4NlOykycQG96SZkiue5hDoPWtqSsOFJ
41niic/Sho4+0eQf7Y/4X7AJXhNBIAzSsWX1k0YpDWEgyY1VzYqWAmPi6N7m+6RqbV2giVQXbNI3
LaaEVHoCyk5ocPiDUZK4xS4S3SxMJxgKdE8HWhqwzvvYgtcLbPE3tL1UkNDHyQyLZW6d3/GZB4Lm
68T7TPlsHNSrN7xN9s5t01L+Tk5mO7ULPMnWP8X2MKaxga2O1OTsNixSc1zwG+R/OsYd/MwI9vaK
rvfFFVezq/0uR0E72v2b5AzRk24hE+WMl+MZMdqBDfjQPAFts2K/CL2PJm9yvGVsN8oY9F+V7TZ8
FYHdR3612/K5pjHN07Hg8hSEQDJQPIUvyJ1ouVG2ySpRYFzXoRHUXnrdDXlHkGgtg5JixzoqwfoB
z7It6CPPuxiegVewGP5f6AWkeAv2wQX4hkceOew/ry+ZUz4DvHYvYrAwd0b6OtfKbLcViqEiv5+u
wu1+UcGRYN8EubaO6OlwspdSglL12pm8I37sGhiXoOhvPp1QOm+SDrf+ZP3zT7LiuPcnlP5itfZh
GEkzf7FJSbg9663x9b+R6hDIXxhIvaO0NUM8FI9qfeqFDrnA4g7E+bVA1tP7BNwG5jBfvlj2mPqx
kW3CrKvFf3XNpXdVzFGwt2NCQM/54kCl5kAbQb/R8nohKbDPZfZXjPjLf0IuGfFTWgFDG3wmAQLh
N/fI7ZCUGhtFZmg4BeKGh3jJCdbrAUKiiH6USP3d/xIYg56mmbDEdoiak8GWvokddeFkXCMLg2e5
3LtKrkCqiNxM7oy2ZYZkoRIAoVLD4JTubI6RmG+bkFyzFT/aoWU+6Lmvsw/iBXHNsL88pdA2g79O
tW3A3NqI/4a97DL2u2l4Fxq8OYDOtX/rU2l/C4UR+2QMgkP4zpsEL2G7PFSONxeJTcsST3QwvhG0
cFlnkvSzcvSFNNHpg9wTJ7zQq+lASYPtYPfINU0Inc7Z+4WVpEugX/lQqiJNhj1sIxj7LSNkpfnw
stjSaJLmxEoBGABVXWpYSA4t8prfUXRXFA1NHwnmYm/Y3Q6a5xCCFhjbSgXEkPE/32/WSmXD+IMf
mFe5apPpRlx8fnR7V5LUKiZaiNNnXIgr5NkvWta2QO8ZKxdxmXs+oed/1ybatG7RAz01iNG7heib
HhKV4YuJRb+B74erGkCTQNeJ36Rd6uyX+teiXx9b9DkWRXVqvN/n1GaRBGYudRyECcmC+sKeCpbf
gyoBRkCgKbOWaNk0udmsvdn0KCVSrJjRpnOG3zsEjW1C0+FAzVGRdrIwv/mmS694MKYeOd4jUl+N
Tm8T39G3uI0BRzxGJSEQVX0nMhV9wcrIMeH1CaBJH/7Fu5/VgfXPn/sYSIXQuBF300tswoetnqrQ
i/arxxZv8Q1z8DHCkwzUmazs6n1r19Rv+TFkA80O0ok0VKmmOgc8n42QGeSAoVXWVWrseBfcaX2r
XpD3nwVycHUBV00qcL7zFkAnpflUtqjuypL5Qt8FNuo1SSUuEjaA5k1FhZAGZhDLHep9ax7J2Hqy
gI7iLJWs5NOp3fG1QCBE/iQIKVYxJaepUmnbTGyvuxDu/UzXj7X3LlukoGf7ffXdTuSjmjVSwqP0
bVZ5C7RLYS7df/3d6qbwAHTDD2jX+8xyGkInysv+vyN0tkC/MJblnwi2kA44dRhLu1FwVzYEuJoQ
bFhhIlFJ5+8xNPD0zwaDNnjVkFJlE4ZHYTiqQRVjLFuasTXidb6BC2Phbao4OntPCL+vX+LY3dsb
8SNhqw/C6UOYRJwmEiy7wT3Na/83oaWhpDwZA8Mob37pQF0tg2V14p/a3uiP79cdMp4QqB6vXmPj
ZMDjpgZsGaKcWfU4qHhI3E7gYtjzeLlU16cPSs1V68TBB6Efv+ezJE31itl6ptFNlOvA8BRYTA+I
P4iNGOgXh7BO53OeTBFXoqBodMocU/cDT95o0a663rMuC5/EWeMfGDOnXnvBNDonxZvPLeT7rrD1
ioyzw2Q0I90nSo18O+9nT8DD/Iis4/Rn+G1itK7tAgLoqmlpi862BZ56tG0jfDmPMbU3v9yBICL4
SYVtvlKmWokKEwrdRL4ydxXxoO1JfOweM09ZwAdkzHNISZiPTkHeIf62VUvpF/tSVi1wNZ178sY6
hrJ+fygSk2nYLmm+9eZtOdFFcuSparFPtDC4fvakt5r/whkrwlBQ/z5AWUw+wrWNSKbOc+PCTUWR
hWN0qClma3+5VBHrndF4sGDkdbMuA5dN03RagX/CgGttZ7Ux4KLtxwnbDnPeiIKVbS+EXdEAF7Vu
Uwk0GO/xydaOpYH2bVTnAftrmfv4kUoB4VmTlaO310NaP5HogW0fSP1Khhg1z/yzbiCDDsHfO6PV
0yi60VYjRvJrEDPSqNOtzxtCnvrKMR/Lnan6rApuZJCiFPedMRJW92SCkYTH5w0UFf3hKVUII+ER
p5i5AeBEPeRJ4DhDUtybVsCUuV7LzCkBSsTg8ZgJ5nWhDwyY9woA7WhgA3AvlH55+MZvUQcFUYbi
OtZ8Y+WDUaxlfDfMe0OCAdRUMAYG/YCa3xkKQmAB4zPwKYDyP13GCu+WBnjTKl33NnA8QaNJBAlJ
HQyceNXg/lU2GX6ie1FwmloxXIzRNrh2HX245XmJDfM+EF6+ePfkUpTP337SREWfl0quUcILB/U1
Nvd8iKrylen6kkh4jW180/QD0IE6B7okbjb2xwPW8t6zmwmU4BxcNoMnw307u8gXg8PxOJ462u/b
tRiGvekU0mYhP9B6naS8xuwtxqtb6MK6nIqB6bZbf6QMMzC2vfewy7lGuat4e3Vr98paNCCkP2lx
xxcTAfTZrzdVYp9Ugm09w4mpYI1o5iaVWaf0neKB/h35WYtdNYYNey3ITD1srjJbukgrzgPPJErD
EgmqfdLczse9kBOGyrybI1zaB7N8odlszLftj9EgHei4j0AOx/dWAxNKGwB8R/JuCeXdRQNCn+it
8ESlxFLJXeiXkl/1hAbblV8iZc5vL/zDZ6pwkXaZm+ByC7AHagvPa5IPYJ+ZXXdxo1ppqbQ+/68o
y/1DMtRueQgmQBHttOZD9Xpgz7sXP8FCh4f+0/jYDLgH8imJRR5rgmaGmMhdeBbGyTPS4IfrIjAU
ZYZeHoTCsEGmjOU9yB6dxGAX7oIfGr5Zr/CePv03s8gDuUdyUbk8K94HAdZmlUC2yotsBjLqY7CK
+qTYsBuEE24sMY9M3ueOqlNId0OdWPUWpPjmwNmsda2TdH3+E0vbIBJxinoiLcZ5/TlTuR1xJiRp
qjE+l0yBed/FEOA7xsSuFWPHEZ+3rWov9HdvX3CAIvMUxqK96Q7FdQeRIg4fYDpgXNDdwS7+7JGy
PonPLWcBx5vde/YGqwlnU/Ml+WWyup524zIqSVNA8sfvDiwEDDofDUjnBSY3Niyb52okP20zbUG3
iZdyB6mdFJ75f59FaB5Q1OABr6Rjoq/Rr9LgXZCZwL7qaX0MTprjLXBjXAu4NsrBv0prj967tcuz
JaDpnMBtMJgIOIzxaa3gYnsHRxRtL+Yr9j7g67LY7LRRxRUsZBwjxqhuU47N05xIdbp/8xfapCcs
gEHXXQ2LkcHKhuNamki/7eIu2GN55IbD1974trmDuBMYwPcVdRvtaTUGSQQuXY7LZGmTc+Rb2gvn
nR+tlKb6cxagdZrMM2GJfve58BrvlbogN9xuGCIJH5h8Gz88+apAwrgCUvY1t12PDKi3Od4oLrp1
MpsueHbZMWPRttipAo0wqYIQ+BpOpy/PGEuwFICsUHpMt2aW4+QsTRl7x44r4D8qXDuRyCkbw/d5
6CkvqkIbBkfNLITOVGI5nHFvT1Xa+5rfcKgRS/IimqEkT1FG2uxpKKFOTf5YPbV1qr2UMBaWzFbc
ZW3SU1Ba6Bfvy1c/TeiCGMsHlAcwAb8RCWHRxtV7OAwFzEaAo+wCUpPXus6X7zHYlZlIoN5BQoGa
acBisVtbWZVt8HktXXLBrE87gUsQqsfKzy8oxMTWgGh2s5ImalOrJn1bG6AOQJDciSTBn72OdNBD
KuWewfOid7dVP5PRfhype+xB9DuBK3Ea26h/aQyYgEqrFdr8kp/NiawKu23dr7q+2NDOrsfpEcWH
MXv3TRlNNdPBIPhzKAeGMyHoDXrb/UvzY/OzwpqG6DVp16+mpEeNWPBbz5RLsCzazoShwpztLfYY
+2IE+2ys/xLlK92AoIPtq8Fzbsd9Bk1qzYqWhJv8utkkiHD7eacoVMf/bx7mbblfVP/FX0dHLQoP
+Dc8kepJVOXPLm+wDtq7V8mCr9bEdShZfgk/VBJhhBSyRSYgpPVTjeY5jT1GSFuECeb7lWtblqD+
/rZeShCwZOCZMXOZDumWu0sGHmtx6/UYAchfNMrEPf4gxhIjk6C2yE9t7Goe5LULFKxZp26Ja8Ge
EujXiJvpYDpPC0pK9hzV8cOu5JCA5yrHVDiAlEY/cwl/pa37T7Bi0a0si3n3rS6Gpchp8ksaoH3p
CD8/HAKYVzEkuln5vrE0oCXGygBaliP7dz9nVOZlbAqNEM0H8tBSVdhHfWLjE7B7Rb+L24FWTj7l
T+jl6U19+HTOAya+0zIjAs6G1wM40Wn6ovw//GIkLoTeZOXDnFNJJ6G93J4Bfz+8J9A7vwzSQgPr
DAkLOCf1MGPs/FQXC/dHk622e2YQUp51lCKuSwgW17hjBPnpgpUCgt/yDaOqHEP46Ewbo0tKxJKi
hbQGcPElcm+pVlYlY7krvQKSirjtYKF+6N5A7RLViq+uHrDv3VO+M0l+DqUHjZVNgAwHzPsmI0+k
IMmL3FfncmlM+tKVVgwHNUPQ1tR9RkaNj7mjzbfRVDd/oju/l0i0usMkGz1mU/kos5pIx1m/pVdT
WPTewBLtvFnK17K637GylaDQ4ZrtU91nACSNvQTlOlsMpmqOcnnR6tKNj2eNkUxt9bDFeqQuIJX7
ep9PrkiV4JvccxkT9TlxIARtvVBvbbNM7TjblwR1ol0fnIKP1WS+ZL6J0B5d8kf5tMqMui0bfMFP
7bcFipv8d/0X4ZOp3S6zaHDOn3KSExsmLCM874lijZAs+8HzpC00O7XN8hNtxO65tiZ/BZjTy3xz
tDuyzEbqwy/cozT3hnj8kThtxhpmlM6wTRItcN+CxSN8diohTxza9CKNSnh13hpVwD3Hcy978VPm
fwLEh8uDwQpuaZrnt0F5fBV4xdnQoZF8YpQA7GUdK42NSrwDFyU++53F872b2WfHRutCiGELv9nM
/Qn9ZUVftJAdJRdDn00bsAO5lqFrD/dhVRu11T7Emk9pzbmVCwI/fd0HGfgqfvM7uz1s11dBbmqH
4wTckleB881EqEeNZcZ7OFPBGouIoZuLzsm1xavzDuMveBykbS9nmHeM/6/xgWypan4Vg5rgxFy8
F3n4h2oOE2IidtmAwWMSWMsZwFHnS2/NZiljZBEsB62cb/NlTsQXN0EkJ2jHJW4oqfSZqmaDz/+9
AWYqyGqfKobgx5ZypakK8ljMOiCLMcMDd1ntmT8nzrGwGccos7eArbIZrxSWhVjSWaD5lr2EWihF
4oVie3NHF17qwDVT5x8LMvWXs+zYbnXislWmXDgVKLWk8xgAyXHFTiLNnWYjAD1zZ3hmxQ7eTJhZ
x4nNuG1FTrGmrRa0R98e+Rq/r6hnanUvFWk8GC4VcjFLWDsNsqDrvenVrp5f4N9S3emk5SPfidqW
7xTLJcxNicc38AOlVDG0539oKjBKsWpq9qb/7JgB1mrDXb9CXfpC0jgYTcpvXG2bDsT+wn0t6Bec
VZS/Fe+c3V87vRWS6pWep/Zeix7fWPTnwCTsQHJahaL9yTqMuCidmGgLCY2KE8wXeoaz+a3RLoqo
lIS/fj2Lh3gBe+qvTSPOSkz3fUPlvrvIg02igYyN1UjTvTBjOnX0PbvKRJbtKJwt3n6TKULjIPdh
cfZv7cyPSwQVALft6Afrvx/GqfAKn2v0rvzXdO+CR8yqj/niIqwxYhx2sYUDkgsVo/9j4RKhR8n2
S0xSiSbNkgxAu/1vBH178uXplsGmX+c7nuNGtznxFraRJGllEOXJuY2jC23asz2JQvFD9MSxahum
VVh/9xAUJEJKYfbKxFvokd1MiC3w5PJj5VOzHFoCsgO8c7kEVruyvktQGdzOkCYX8APl0qnarkZk
hOlW2bKiCttlkiwF3dS8oVtWZRULVBwqocW44D1tU1zzEzM2/4CvSSWZWyXMOT15YYdAbbsd2Ofi
HZNB05b8cc32ChxXLWCqKZuJZ1D88Vv3OWSMuARXYSpUQpRJ8AR9sDraEwHIALzZylfVriJZtRwD
K+WM+wWVllsNZnJMD6W1S0OZx1ARCBjvx2j94gnIAR0P+FxFBuB3OL4ISXFdzMnzYRW5DLJDEFV5
68n5Fwns80a5K/VNkVLZ1/Xi5MRmxWJSPMLhF7DCaS5QAW3mW60oIvQfXWH4nozROia+fai2QK3o
y6jy87EbV36t139o6ljtc6oln0yJcaKQvQW7iriDeYGMpFATw/7ijp7y9gdjTiwfbVoe9b036veK
6ztaBnC7LbJE1mmgQngl0ERsqW2OLwbhibMcK46kh2QVTLk/nHWEUgr9PNXI76Lu+ybsck0DSz8p
CcdweUMzgb8QFrO7n2D5+PBM18R+uUyXz0uE6SNGhNZoKWRs8pE3PRpggfKOYaASa/t6Dqta4/sr
a+63HNBE4MiQWZvWgx8u5nw/A3xMnEsCeQQEFboAVZxFqQp8/IUMym17AHlPT3KcNRXlmxVd/NQb
MU4PNmXnDy2J/WVWwXSmtEVHEoa4gufCbNnLEEvC3aA+6QZraWcACf0FUinezvCE1HxnmpAu0f57
2WAPX2qEYqikAiZPtCIhx60m72aGZs/D7pAP4i861+M1cqAyW5yF2+ZVpaxsx1Bj8k0PElWCIoxP
TNwgx0980Pqs7Qx1Biap/84STyufPABkXtQXsFv7XZCOE/C9CMLMwRPWlG9PDP7x5QtNPT2uvVf6
AmxFrMf5PPUyl1bswMRZ9vRU14gcf42R/p96EyfnGx6D5SWuV1NlQ/Ji97H6vdBip/yrtBLk1Ij0
ELnZdubvdZgFWpMG1CBFR0GWilPDHPI9Z58qG/yGJ7TLYBMJpsBezJ1TmrwFQlTxTKjHpBqHRowJ
hhpW0d5+d1/LbF9zgieSOH6l24Dkwi9Q3EXLveCJsusJWRAdw5bJb03PdBIeJgqBjMvgVwsCTUun
PAdcyMYWwHDVx134xpe1p4yKFSkxEvGvr626c2542Dzox38Twr+n9t5f4JNjbsO8TX/1DiZ3cyBV
/DqBTsszO8op3sTADsSRIS2jmw+wXgcpckKimlLtfIHDIDAgKAYY6hkb/TrevL8mozkIFNjesl2X
syPw9uiQONlBIG93xV84X6VIvEQ1w+939b5juEw24szrfqy3XZQu1tR/Zha5W7cwAE+/OnfkU+4h
bkDzFduwxXoQwUh/UcgY/Qk/nvA/cNo8QjQMJm7xxFPPxQGbeQn7inSugNp0GZ5xJMAAozZZDLMi
OZtvn1d5AQ0oKjow13+Ek1SSIwE12RalkS3guq90XNUodhTtNppfoV1eLF5D5+RE3Ze4wh3ccxDy
JYnsZjOGgdNMOQEB86MonTPaEkcOUc0ud/UQ6xJGxgw32W6N04rUIJEjHBSZ/KU9hjeEgmbo7LOj
HgVaogvpGSerjwgO4wNaogiELHiU2YOVNVMsFaoqRx9VUzqr/+108qWuZz/jerJI26ZAQ7QzJDKp
Zf3jezYpLnXJ05DPDXcAfO284Cwaaes1/gZ3e0Xo3ua93Mo9Ck30k1V731OCJe4EvJKc10wayiLr
I9HxvhSturq+RM8WmQs9x5u2G/pPa8BuUVGnMW1wIFYndIx5N9bSrjZdg/MAWFTcZOYiT8NWmjCE
10swdvquJO5Yx2RzA4T0EWVaZKf3Tl/Z7zZxdcg7xPBieyfmSjfco4m+3R5sSty2qogqEeclIlXP
rQivF4i4H9YBYtsaJ5IJn//Wfe7kylaoE8iRABdnXF2JVY3DFinidxpEY3bG/hEe67irDLL3/cZM
fwrg8+jQiIZ3zxFrH0xgSSnBQegVSvnm/04tZbcvfVM7u4Os+7prxwl5tZz2/xzj8l4GVMP2aZu1
Eb8KSWr7O0ooPJ0PKPdDWabS31WC9vDqXlYqlu49JNY0KnZR3yZnaJNRjup0qCTY1TFm1+AVAwcg
hzGgsbS7OY6tYd8tU98jV9Lpzgfy1W7vGcGIzfx7oZlIBstiOVwl+vbazeA/jgIUtcgUjV4PIV6e
KkfQ6murpDkOD5E8mJLaguysjCs2ZInB5nSQy+1qPWSiEuxHZv2ek5VEZ3k5od7vyl6xWGMy69DS
9yrHVOUgAIz00GIon7gvUzInt5re747XwX3i2bZ6p0vwNLlc4cexEco0Ab7W67AklmfG5zvuU67K
wSeE/vvt1r3U2XP4wTXaDseVhouXlochabvbn9Ijksh9MXkS+AFnf24x+dYClrbOjeJC8bOTN8lI
jSZweX/Y/lIDzElEJy0ULfs+ZX+3qcuotBFrTPX+KBdZBibFAdwa9qvmZ5sev84ptnb+C9co889E
clPhvJ2yDWWCQbsq9tjDRPJwS2NOoJ8forSqgs10sOzGHr0990y3P9WnV/SE6M9F2BOxnRXGsogo
OIwgVYIGYd/S9myT63zthmgajd0N+dXYxkG/p+R0WfswMJ8/KSkgA+N3sbAOdkxX03s3sWcciQFD
kAjh0keCGyfWLb+Hw3OdVp6SgEWCpnW/olpxhq3WV6fpVJkykZTTq/Txl9PrwFGJP1G1HnH4gaSa
ri5q0x2wLalsFU6r1NeozSwVobx2GmuFevb2/DZOvAci3My/zoP2Crrccb1fLaxInZV9meBoHeWy
pt/o8tpK/ZOLv8qBgmneV7WiskQSyKSYXTc23dhEwrrgGS490/53DEjceUyIYoR66HoQ4l4UpnLH
EpC87GnTFIMzTZFaKT9behRruVkUxqJQNhpctreaZuAPaO9Gbz9yF8Ipd6SM1tMqpiR8jhC6wc7/
nJA0ddhjLzrRKpgNMXHU0ZgUAzsrTFGZHrOlbC4Xx3K6EuR+QFgNgBqAdvtGdfkRxQHhrXq3dijL
yuBYlPXD4PRzX+svOBePT/tncmJbgzyM6wJVSZgrY4dYg6x4Sg+W3cUePI7lvtXPzJCW748EeQuw
x0xkmBTFlf8VaCnWz/XnlnlomN4VdMSI4e8BzrqPHNPi/J0llAVK9zNu4or46nAgqTyVZ6o3sqwQ
Eg9qIfvAGXRA7orXqOFhZSO8XLl2WvJkImKSzXTaXiu6dWYymDMuB6dt68M71SJtRihUgbaHI0u4
VGhLOAchX3jZJp/K0c7PriCxX8xjquWRWiDKe5E/5mPhzMnPHo1KdkUvdJ2vf6dJj97iaqqQN8mu
q5xpYCITPMJ7lzyZ3+kqhqJ72pVV05IVR/OGLo9j0oDCsAqZ0OYpZwVJ3S4m6kLuUU4tSaTuwx/P
MIESTXz/Qes8k0VGhsfIVrb0WHKMbNjndAd0rdXKX3y6hrFJlrHBNEUBcCUBNa37V84qqpe9bF3F
yI1dakJLmD+KE05Sn3Rjk4yL6Qs5b6KonPI+3Mlzw9xH59fN2VtyaSEZUaS19euYh7oGua6LnWyk
q/xjntyYUrcdaQxOkVDnGCs8gaT7lHA6e2rcB2EGoBy6f+rpeU/dEQ8Dblq7a4fKC+kJfgzjMAN+
kUVCfApk0MzHrO6Bui8CkHNk1e/M6pLnEMCYnvSHfrbrkdprOhQw8+0NdTGZ7YHJqWYUw0PJQH9d
uMAC+ZAequNAGaiPCM+Wb1vF/zHB4WjyEEvxgxXkX8Tl3/m2LXrFXugwp2h1dPTzUmYmwHhKcglZ
0O4PXEP8lN65BucVGw6IzFT/BSNVOeXvuZmF6qj5M8jJ6pQ+U4EyT9FZyEdWqqwM9/EYGuiGAKwx
14PynfqWJJuxvRmouoo4Bvmno6+G9W8N28wQCbSle8+r/KldD8+XYjxHBN4ytTHdtEqSw8cAo9uv
W2bakJo9GOxrd62RI0w4Vpandq+E+MXZEej31Uuv28zCmu8o+kxL1BESyqbaf3iBs1DyF/eitsMd
hQ9AxRSvYBqGoYtfEyf6tJyoN+nRZF2BK4L7RVtHVTfu3rMJksvJM1RUYUC2EZ0pS7riqqWiAYYI
BZ0KzdA6g2fy1Ju0prJt2tlldQ61zMKl390B9xc697yAX9BEFzAYpXlsa7hgQovexI9lZNFKEumo
8yhJfMJEHC3bTIuXZQoWl8Tqwm1V8cHOJVgsbaXOt2YAO/14Dd27NA9VFea6OyKkCpJcf+oihSqk
vLZEahijFu7XbC1jdChHt6aqMtX2yCi6rmtVbsOC8N3X9Jmx24Addz9SsbgC1Q922ZwRHGa3Kdhk
z2jTTjTDXN2ZUYTX4zxIFAsude4dwYWMCLU76oYmuDaRtyFoJN1BjS3NRWBUKIbaZ+nTLUqqd8Ms
MLXve6BIwd2X3AxiGgGblcbePke5laePPiio20HORftkpsaa82ZRhBab3RNFEnIGsyp/GxDywcnH
viifuSJErTQThURIo7VQEyzSySyYGfQjcVakzC0fsNLbc+sXLNoqWzknuUhuELnaH5dNuT/eS0DK
YQNzi+eotOtOO5y7a/TP9oanLtwwKVhPi5/ZZZqt6ex4bG4QSyTyhGZ4dYY7hQyiVRfkSTFZBAar
1QUZdIq12Y8LGutd8hdzdO/QpJ5nXCfVcMysFvQ2bYUx2lKLgq99bxYeP8SKuH6ue8MWZD2a5Lx+
OuXX9hCFVY1ThZz4ADFxcm1+MeDsLOvA1R5PS2hpyH0QI/MFwq2YCr6+AWFnZukYhZk/qO4uLG0/
q5rBhferRyKvm7L4w7DXtz/HKn+tk2m7ovL6yPUPRLPV7KTsMUY3bydSpowxfJONkaXS4ZIn7HK2
NjSrItdR6KS7eOpHeboeoHxk8kDYFP4As2OK5zqEzo2RP214HYGetMhgT9VpnqrKLXB2M0ECV3ol
IkRwIoJtvbwJCddx5SkKWGB9hB1eJFwxb+fI/GXl4/12C7aHeHywRPnxWodzsITxx65cHiItX9j6
OwvCkpSDSRnv58fEg7/YbdJcJAf75B2LfFBQkNFnMJr/C0nxs1zcJ+ZAR90fahYt0tn9CvwszA2+
SbR9AnMEqozd3OOicyPeIacxKwSTzmuVObLJsLgUdFAUkKoZjip+xAGx0WEc6YsFYxg4T9uWot/z
JmSxgLMKZC7uNHIPCg2+ULqRuqfK1im8w6Z7TbtbtpnStBqEgkH2j5BrjxLMuefow4xm+Qwxz7dx
1TKb6WfWWzI+y1PJ32iwiSsPlVm9a09IVhmEgQJx3uackvAmvJT7YVcciIEGeYWHh4A9yDXXwdUk
h94RV4lh+nVqicvD0GWINXp7fY1FwheWdBmSidmfSk/Y8D/jUgczKXhCXAQ7PxXslqbylNbuL2Ag
X9BjI3216EziU1oqpSzqh+XY20rOHTOAkJVKasy5RpT/0/STAgnwzne6qaA/AMvJV6kk0PnfqZte
+Q8109tZOT576g9Z+Ml3OD/iqY9h7d5cAI0GR2biijVGmc7/hZ6K7lsBxOys66HPORtz8E/jfuKi
gw9LMjIzWziOqFjANzgey2M24j6M8fBveKHQpbdraUBbNO21Kx2A4cazw4+pIxKt59CFDVfDPomY
WFEVmce/dU2U1RJEFcWA+cSp8KonqM0txX7LfoQKcSZPa0fJQBIr8c+AeHPHruycJRYLa/a3Wxh/
aXaV8uOehlkyBKEJSG+GOgX/YUFRThT70k07LySzHKuiS6KgGcnS2z1sZBElzhc1lNH1m3PA0fNa
c9GltZCsyj218b7STBx3m9HmLiGmDl7M4s+XqteSbgrG/jUTayyKS8SKvfKXyNTVsLUtvnVTOxTq
DRgkssBbcQBB1BkqPkJLASmESnKvr29lfICL6jwPTwNKN9UmK3IIa8+Yr0rLy768wkcsZ8p/A6Wt
UYMMUGS8KiZXxSIpMfhCAnsoLH68bpjkLao7kzhxCHnoR5rwcrqveXc9+UTjGEoaYmTNrBAf/cuU
I5H6tpaqOQgea8KhRlGxEdf2gjXzCAlsYWhyEL/ZlXpmAtnRvMKO/Er6iazQEZro6NqaYKH7O0s1
THsktRWlJVw960xKG4T8lceM7/UOZ6dB/k0iopCBW+8VnyR7sUIAnDzrABqB5QLwZsMCjPSAQNvN
4Qc03gz2BwVSrGm8QHPndYatOvH4y2BTfUncZzKYgZee0qN3T1SPVquxS9pm3OZ6478G+g2bwj0Q
THpe2Wa/BN8BbkiQzSjp1cL+NZjU1DeLTy74TUVxsEqe2PqfPK9iclZRahibvFRJ8TX0p9IyWE39
zvXPxG/6+eNQkyrO2YL9uASU17gDZg4NYr82iMk+7pR3CWTfaSK2ShFOT5Ci7Fx6hEbXWL0Rplf2
ylIvyJ702dFqhCRHWswNoRmEnzHiIlkNAeRuwqHrYkGd3P9oxk5pNJTOOrQ1U3TWj2LhVnYyguaG
CQEm/y5e3Cg3QPdySs+R544BsUJAOzmty5URGaqLesMiodDwoePBrxHQiNOBKsdsgF8qH0LCtg5V
smRHunr2pBF2sarcNL9sFS4WcebTRnbG9KPGHLid6eLYYNMR3+jm5FjPvjUfQLe8l938Ig8TkVuN
L7eT2hOXpFEZqLQQzTtQS98qrg6vk//Gzz2lqOdXPZp9oEwCimEOC1Y0fsbQb/kKEPyvk2sxuLn4
Hw1IUMax0kw/utN7dP5Lulk16Fw8q2rF6SsJJPV3sQbcpNbqXpQLJ9Xavt1zO+mQdv9cKO9TIkSG
tpsebqwbTMtO4TD61C4rdiZlcoHGQ8XkTMNALhJXY/4n7bjmgBOLr1hfZTjYc3qMiFOC67NGPI11
7PZeHUZ2lmANBi3dCKp9UbfzT2zWPMPQWmLAuD3jW7T6MjwDS8tUQZHrYSKti9dRehwWMnPVuzB4
Ac00GX3q65hb1R+tO7kPfAG3p+AzVrV0xbmcETeImLP/ofnxSRYsy/Mq+80IKjPHP7wXoimNmXd/
uf97bEaka1ji6Q3+9ffIRDEIewMt6/J4uj9to1qdwHy8cRwc4dh+cOlCKio/YPv7Wzps1z6DWh6h
MHAOgN/JHcKeS9Btb3ffi9Q3404yyzT0ivsyQ0Qa3Bl4xxfe4jvcz5/eWiVI48gapmZAgkkqXqzZ
rp9f7Hv2X1qr+oEvbMnfXGzV3WDR1nmsdO9NBufLN8oHAUVXj3Wc2FI6WYdvP6mU+25dFJsEdTCN
NSs5p/cFCg/HVDKEb7t5AL0RI0BjRnn6DnSy23hUpp4cw1NSkQkOTNW5oi50DirVx8vesK1t2/gX
0AHelnHhYy0uIBWtAcgJCnkn1IdyQR4tpRxjXN3qLL0WTTe/bXbQAd0KNgl5AcnxtvBBcNPGup+H
KVm1GTlh6Be3hNcTjPcb8p5L3lcTaupuEeEEDIwr6je+QK5yElqk6ayBkzoc47MJwPkUt8bqOlYH
472EYSrcl+WzD2lDTdpL9DGVSt+w/E8Hvs/g/jiI3KIvufPk0rX9VN5+0CBXzfIDcqhDrVXnsrAU
R4HVq2BBYKCkOKWpVXXqhd3AZ1QgfKrNvxVn8garneuZ9E+x7f7NG6iFJm8JaeToftk/BJeJWSiw
vA9azqm5/c6YgiCTZorckPO75m/m0wrXuuVM9bWAIEPUzmGAa3EC9TcfZfMEEoUJnqek7U1nd7UA
L/jMnFWaXxoLlUU/88iWAc5s80dVuIDfrdG3BNSlE23LsZmO4f/SvqKnr85yV0Fda+P3CZsogUUP
jlUe+l/8qTF/29gu3tER7MIDmUs6L1YeFg6OhU1a0EE+WhTie6mFar/ugW7tezVxMWwNutmldw6B
eLb7MDvN/b4+sEOH5ZSGw23I0VciqgyM4Doc/cobRiwAGpUQ4VlgRBreXXcFa1JqLdvOY5s1P3uw
X8z250NR5NxOOSMnu2aS/zP9nEcanUGaqL6zgJhBSW0mj8AQ7PQhIatl0B73zly2051NmKgRsjpr
7dbhFQzGooUyrjhnk7of/yZpTLrsOHK40E84FmDnbANSABQ8352EcHvRTH3z2ug+5nrEirSDOXDl
nrg3ANT3AwOAu3ifX/62Znr3WXiNyqwWZJ9K2YaKidWEhEXm8G7zEi5QEb5cpbf9lm8MIMpEVf6i
tEK3rCo+ywm1ol74Hk7RYBGDC3aY1dxOsg/zK4H5Pcrl/GUeILOreBknOUeTcBMztDRf/mpviint
s8pYBok8KIibLazMqThLMPNeVzpU9rM5M5FQz64S1ZJOEPH2CPCCfMSOURjCiYh6R+e2QFiapE/I
kb48/NmJ+XTX/xcbZ3Lw8aCPxX5B2A7wsdqeKeyW7SzDPLLQ59WTdipc6InrKmlLZCZb6Qgmshne
W3t18gsq7/W9Jmsa8pBh7mpjolWpexHUMcrwWpkNtVfPPe5aqspvweFj0AAS7yYWeTRQ8Y7sRPjE
rwAt6XHJIMVk7O7OMgoI8Zkg3FEzM3RlMZXW2a52wKAvGlwGJ/OHSuIJDWruYrL6CrDPDSO4/q3h
hG4JLRS9Lw3EiXRkup2FJnsZC4bDyq74QiCt3TMWknRhzCQNEmB1Endwa0QQInXPkFGbHVYvQyOG
1a0sKJPKo6StUmjZl1ilS+JoLRxvJifgcRjBC/azSponzKNXVqVhvaSQxI/ymuh+0LvApbjCAE9v
u5QSL+r635b+xmQwctAh5bWVa9IR0K/c6fE3xtn8qtIUuKysR4cvh3pihWMltBfqq2geqy25jFOC
knjYYMd3TKP9gnY90akyc3t8P6imJswvXL9hw1uZVdCrOk501jYU15LAKK+SNjAEEUVBA80TJcI9
0lUwBD2FEWSqSHiVbfQYhi1hFWIsW1GJpozRaFWxs0h469WbVf1HSMIFo8GyALO9Af8CySPQ1y7S
0NyXPSQNL5fL7LrqTMDOco0nJwOlIj/tRn63jKxdePTefyXJqMJZ+u8DOen6NguwTZ9M868rbuJQ
+SvqndvmQTzuwjhEPegCRVGBNLh2IuuO8qfWrLe+lX6NZg+bI+WAmuQhjfbjlwh1d/pGHMSjSE1q
IBMX9lmBNwKYYqFKVlaRPiD8IOo3DqezOOWE460M/vObfx8YflFPh8Ul9CvWQ/IXIcUVUDq+uqRt
2e5bCaTIfgvb/PSjjIkLcvGy8XI4rbm0GnhnzuJmOJ/vV2N0sKmytK01iE7mc/cVOybNrU1Z4e0C
qBIlkim2CFiLZ8r2yhcqNL7D+88Sw7a/gjsdohDhUel+xQjZ7mLh+xS1hMsrX2OpggkxKkG9coc5
Rtp6b0/9s0iPQNgyhOg8gAtH4PhEReeEBmJgBCdfeqTvxMSLOY6PxlNY3UbwaX6EDuzJ31u+jgMt
qRxCP2CNobM4YPDJIwUKjHXt/W7W+IG8ZVWL0IadlTsJRPkTSK/Bo1utbnPieMpP7qPuDHuwWh3k
CEONqAfz4n78EQTvs4MLKou+jlcVqwXcZciD0DNjtaYZh3WXg37Nh+Q9WmtPgA5ZxOVXwkMoAWKi
N230fSsp0oYCotg908AhkZo/zotfYrOxJKrQJfFj2TSIn0ASg0mXHWPBZxDEb+solCMiC3ZcnrLU
oKOcgGj76t20DmkL1jgrFYARibyAhafTwBO4+HAM2HbNxkzU23Wpsqj6TwcD1f/UX/3BcsrlQ/li
keB3U3UFk2kwI8941x8szsT8FMT7d6pW+RnAbsUo7ru/yL/G7QpkKN6rWIQLv+TTSh434JGPYhSk
j7zcmkBpU8EipkiCSQdnXBuYpB/I0IxANFRn28de+TuFwICmufyqMcRcwTWayUzEO8GAMkxc2ZoD
WqNE1kDnutdY4fkIs3m9lvKdph1rw43dR+O1tapO1Ba89HEiRl1iorDWIO65Uoo5SWI7v/B/neWM
3x3BtoUoEDZDQlMmiLhXjSl6Cg+MUOl0l/CrE65syIaUjBRbJ5NT/8R44+OXqXuh0t/OBgTArn5Y
t/cuMtI+/lMmNFLgUpogDakF7KtLHKEvDbNn5oJT/yCLiSfo8TFS9gnEAhDh4zIH1+1HVHRxTmuU
92ahzgE4OHk3mOPA96DCmossM0io+N+AAIiAQfszlGZgGndKV1o4/yNnOgBW0TyJ//sDZU2Ix9Z6
XevY2U6wzxDXm0mNzh0dYHZ5Jv3mHfpuXdEueCEwdiAdOMgSjfziQQpeLVLng6tl/4TjhpT7XT2n
0EZeaDPcIy1yjad9qQk8EoMWmz9jfMOUbdwahTGJD0qAEkF74xZg4Jhmr5fJygtxNYtYPBc1AanS
iHc/QR+EL7+oaWqmj8GhYFNeC5goYUae4UkHC94T5hkVBqot7VkKq/zoxu/XI+ALyFnArjkMPTSV
9Ut5hlz8JRVli8Zr9MZ+aPXH4SOBIHkwJHs4bGKsKUOP8bLGREP/gB63AdkS9iDmyr4HJIV9V2Y7
XXzlI2dGzpihT0xmRn4SxNuZP4xlpYdYtoUDElJnhWxT/6VP1HVONVKEohkblUX30/03pBZhwDdR
AtLaCpWVm6/uKo9PgGR1kHNtCcUAPRVUXrCai1bwevY2VnudFoUBC5u9lVuRcS+XprkNZodQt8bZ
cbOm/j6GsWiB/kmHbV6tN18b1CIQEnymy5ZXBr0d3kDSNQagjc26fUgJvybAZEsm64vXB0aLNieo
0tUmMGZOjvt3TdFN7/5YKFSzmnGV5mPPpvcFdKdC8jZbvWwXzVV6i/L5LjJJ5NqKSVJm5zg6j/YA
G7RdC7635TbO1b3nPUNUJAl3yjeVyRPJubdku5uMddrYu3wvWlAqRsti2Bd9pfMdflOw/uXc95zQ
4hwDZnSdEZ6QkQbTXWZLKRtYjdUfqVfhEIaMAqjfnYbzrfevISDzpM2+QclGlBjGPfn11SBt1hd6
7japJw4KiIpeHwN+3UsK2lziycYwKuRCy5GPwFEkVTYL4qqmCsSz2JpxlC1JYlD2/O4pBDnQP+0i
I0uRFUhZ45GkaXXHUvSprhDZM8HCRgIkSDv2OkjLZrefWEa7wg3CJGUOhiJ/CM7q/vRWUb3thr0Y
JEcPobi7+uSlKBmAs+qCOxFQO93ydGCYnHUM91z/L5UiwW6tLoecqnudNlvn1TxgLjiHrngVv/Hz
3dT8KvwoaafuXdHXg/xdLoNzd9LqXgyyOaxCmp4siZDfXJI5kzOqCHatG0NqE4X3D64Bec0fVwiE
Np2lPaWcR0sC3/9tXx3XDkSzkBWhdsG6sOhx4BGmy7Z6yD8Cl6VDmxj8U83VpA68vGngqTmT+V8w
MJO8W5/YjLwF3ccrAd/AxFVd3OoP2+jibgPMQeO+VPR48CPCHVGyUsXFejXv6WVIP+Nf52bVlWO4
xQV0mPoAmc7oiohXYyU7hUmOxzBjM8f2+O3Je8wqw3s5MH0I6o5cA103SkIlEM5c9uf5PXoicnZe
NQgoR+yFqGCY7Z349maLm797Om6wUmEZ1H6rAFhwMJU7jIfAuM85RZR++YfwnOOQuFj+PwphqFUx
HfHfl5csvg/N/rJ9vt+ZvA9pdGMmnYAqCSCWyd2KCT2zyIBkJVV3GNh+o0TssdUB64wXTOfkgOCL
/fItdoVnWOCQFUqCCSRAJV544qgZrGayfjRe/SUgGzb9KDYgZ2j9gGMWSvY74K85WurPF4ZIMszt
GyaRGhQeVlnptQ/0utHKugKd8FF9Aixtiu0Lm1ws55Ruh3QIf8igzLycjjIt4QjpxMOeaOAW0c2K
GL9btUvULsHBkQSy8UqFPNparOpB+75SddN0ShnpXYoWR4TdXVNLGecsK83r3N2wiqfKbXjqbUUP
XpyQ4LZGX8OR7NWEC4+N4Q3rgDtkh1BVJPvWgQrQKOVAvMekRZLcdh1/9dYiy2C8EU4OpdKeGBxm
4s5pYe0y9uTViYCiHBp/7YOKT2Tb9loXrAdBen0VBONEE1AIFayLnZ1asjApV3iIz2fty2lWmz+l
J0iQ8SZVFOLfcZGJrcqDeouzxA4tRk3vQWoMJp95bBYzZ8SuJyTTTOJdXhGH08F860/P9rLrZIag
K41EylP09wxQ75/vX4OjiBYdfVt1B94nsIU3DfTY2l6lD6iavFyEhJlkYSudVs7CBBPbBHflz6vF
L6gXsgcPnhC9qGXJWEuLTx0BmkEXroR9fEzS4g4Gi9vYrO+lt3K5OJYtoz5PEvz3uZ/0xNisT/jB
uU9AMd5A545AlSLWtRJ/51DESMjWXdvpMwBhq/bcqV6N3ugMQO3N7HyzT0AkUYpy7vvtLllJkAg0
g+H2zdLW/AkQwVILx/8gnCAGk/aL+Ic0zyJ+WnMBLwAVjQPBK7e3tKodPlLTLbdrajbmuX/Z6QCJ
Wukp4uVea45Bwp3nbvnLTsKzT5jG0Lrkkt3bEsdrqFQeQScgF2fISXF8rj5SIKJHR4QMfBkpxL5v
6lnfHc3Kr8kqk96rS6Vq/LRlRj0+2oZiqwek5e8uKb+rlTSBtWT4G0iOHlsiGSx8XiOPEa73x97d
4PU+oYstkI1lI+XusjEYn18gSsyLLClAbrPQXD7SNe5LojAj+iz6g3U0uue80ecB4mFjzjFyDUC5
P8jgpn/N7uS31e3+PJs07+hgJkowYQNuRKM1C1rENWcaYiuBlMNIoeJtDtf+N7IksRl0pbm5qtyo
lgkTK52mj8jsfbKB8tmpBXQdm4C96whGcfRXwMwp8ptEghTDk9lcA8phxOucWbPycXqI150DrMN+
vw5B/HXoxpH0i3eiMv3G9IEPPuvhgEMQunNPod/zzj4FpxkYdmdbJhcLUqCC5/71uMbd+lSeyoDH
nUv+eYPoq3FI3ZboCsu70KqmQ9mzL3Sus5Z50bX71QpFnByav72gAQDl7KZDuEfnXKURxEoGDwTv
ckaqha0T5rb3Qe2DDYK32IjF/smZCxMUD9STJ/8HQN9Pofjx6DpISm32q/Tw13ftAmrc35Meac/h
7KY2ijUDRaEIIvEDqu08EmWmkyqnk6R/uLZW5csfYtFA4y3yzBQVUYonF6wgiu2dCBfvUbNOzUh4
OGAfjZLFILyYjza5vblRL/CLMS4EUtOxFesekqvaz/ohYNPJ6F6Krz8KKTh0yfYEVezh+rLHal5n
xpZMk7ahfUGcTTUWrqOotIcW+pa4zaomdmqjtI7VgHmvWVpkGVClMlI5htYliPamrGPPtlpF6z+M
oXOJEyAGdhpb29ZlGdb1RFXAHPxaeA0nzfBTuC5O9pJzWvl20IsnRbcIz4VYgABQdRPI+o622fhu
6QXnWixjaKNCGZOAJBzxhk/Ikf4+l4hcVD41+LtceZV0owRIzXetbLrAOKucwH18lzdhQ+bLQWN4
KrvxtMZWrPNx9rZhvuYlf85E7+/Rk6EcZE5JpezJhOh+Ev5yJFvlwZYDit8sZ4qxj+ABs1w61UyH
T6gFcoTveBrPB+ZiuXtqv8fCrlUpRbvWz6O6/Alu/LstG/DTkhvPQWi9Z4Qj3y45qLNnh41w2VJ/
/TE73AA0PGRKGHnSZAsDzXJnm9bSUavisqb991XRWNQZ9Pi20ZWVtOXzej21u39q4tkSbagpFPd5
8ztJCSnI+Tr99qFo4bJr4L83Q/AgXfQ2zx2IhBuFzpxSxmVZiQOgrc3yh2MRCr6JGIiHW5IE7BGv
kkGv7B4P9MqHpcOqCKCI9dmeCvF0dL9MUmBuTfdeHwDQ4c6qGak56xr94OJ8iFZhMrx7L7LOQky5
Aw+u38wLDc9QCH6olf+5pw9aRl7LvZMjy3Y+/gX5kKL8zTlALcnh/EPz8ZQIBJt+iWUtgtx3X7M1
gzTVRfKVrmuzQX1y1kl2IDQuEkSelH8feyXttP+Mnpuyhuuc05Pew7fEJgDKBn3qKBtthWi6PX0n
RAZhtUbaSLgpMrKHPasplTqwcsTjP/HYPETubft+M27CJKmM8wVgNqDIb73GJJMv0JcP8O6aUUaU
5aGtOZljBx6U29YDtQk0Z7V/7bDxRXoqhbEzzw6nRO75Vqc9FfkHLxBaID+Bv85kp9LJM0fF3/u6
rNXUXeMWBwso/ulvkhHL2SNuWmstItIg4WhxRSbzFHpMvsk+iHxEP6r1Iscl1/Q+XcXP+itxkVEq
bkEcBV3KQfgx1X4AZ7G2wWy4/1BqhnDdiCxf8WbGl9VJiEv6xkR4EqnN4VMkKphOwmfYAQi4kKH4
jo5KxW53UIMrEaops5C/cZiQy5ZtIodTa2I2I2BsedAlKcBxJ7EVehwlvneo4Nev42DgE3GsulK/
640YPm3jho6BunuU1+2pIC6xTDywyUHzRjRlZfCBqxSyKAtIoP+paIxhap2mTZzgUvNg0kUMibGT
wvescKC59Gi76cUJLJaeTw5UWaqA5kRg+67bAffJwG0XqjnjOeTrxiAWWNHPvDIx6kWCy4xmscjk
SaW9k7GO1sgPNhC46mBDvDSmq65FuqxxHRzEyTJlkDzbDfPd76kNXnLfrIcBKhmPpLzkGrb+vzzb
1zdx2wvLpp4BIa6w9Soq5t+haEVekBA9THUsBO4dacic/owCstvvYSs/oUL+UZL17c/9bMpwyIxh
ccHEpp6PTsTsu6IO4bX0b6YTCI5tswbQ07t9hepdFVSqH9mBIiXG21OdC3vAe+aqfFt4cZmYZZTB
Vbzlp8wdBS2m7Oel6XyAwZRoWfSdPo73FSQNqheTiyk1kpEQLN8bGtxXGD5R/2QFEnynoZEnW/+6
wIjrWSQUjUi+ZTSC3hbhq88XapKGj84zYTL5db+T/CcBL0q96vvLydVE5GOxTd98eAUX7tBGRlHA
D+MyQTJiraxO/1jRsaVmn7y88YSqmQc/7x2jlLQSb/SJSdxJgdgIrbg7sMy4BhHAe5BTVSaLMBAV
X5Tc6LfojxIJ42JY6dRG4QrUfzzH9scBYuwOp1Zhvnq1eX6/V41LeV4OMDGhwUigf/hEB4EQ8Nu1
B3LQSoVMuxzhJVBtpaqxyp3Rc+XHY+0QJX449DecGXYWHiuY1UtgDd4HcUEPOLeFRxU8yhEYjNJy
OGiooX2fHZEu5FgrlINqYFAoeSoJP41MFl3+Acr9zjh+dJEDjLNqasNI5Da5HA4L0xRkzVxARUmi
YKJE7faPI3sdhgleOIloE3UptHEpkVZM/HQjM5Fndr8yKx7IiHj/3ZuP0HgjLYPfsWkly5+irkyo
Qm2lldFMP/PdnpDryE+OpgWG7llV9KnmnWXQebW44U5/0G+h0fzRo+PwBRwqPleF7tq+KhVwWkXW
Jz6CuPgYTKjpAxwRhMbj/4l25uAJNHr5wEKqpq9y+t9EjcKiUdKqTrFfSeZ+ZLWzLHkdalPWQX9r
kndFqBH5N+YAm5EynXB6qE+MIJjdLf3W6RteTJ/DGjaoUEDjA0Tn8umSYUORaZkHb+FmIvQjM3tw
y3ohE/IOtjVKOd/O9X83ThdXWCPvMX7DW8l0AJafp2S0ZDHE9mkBGLP5hIZn3MI+Sj6MnP6fJxLP
r+cTpHAZhyPP0ZSg6nJGuBvQHyKyvJzFOqKhLfKwZxF4T1tMt2s8toNIlispVyH9mH6pHRtE6pNd
2pJFyZfaHMapc0NCMuKUDqw+XMRmDydWsJNNxgjZUYDUund7srKBRJLNrH4bb4pIaS9zUYhy6BYn
djXEbs2Oo7sbnUFNBqXf/ONPOPhlyWp9ujk+xkROnFl/HL81XypmQ79S4PY6641w+wec3IHt/evG
r7kbjnps9aOBW4RK4Kr0sBTpfixerZRj9awM48ULealOPprhY6ai5ktfp6HapsLe44ENvhdk3pXV
8YNo4W8Gg1wnCb7y8CskUVNGTE1Hq43oUC3zJ9c1OgZnANZvd6/l6h8fvpN/B87fnd6mth9LyKLP
4C1DlrKpy8NG4lyAOErpK1PSE0pQDsmltjFHh10fi6M7Ww10ARCBFQXE9Snj5xQu03Bo6xZqH/S8
Pv5BIk4qyBcX+Tc2VXsoHDzLxCJilDTf7tB3zpEk0wdYp3IqTEibrtJTU+WipR6DvpDa4Ga2hraZ
BWZ4O8XcqZjS5fW8LDUjXtbiSMUGmyAgMO+hxcsZE/b0yiGBMDNaBiYsHcZ3/1ZKalCIcsz7c6My
uKAA7rh6z7yPmRBYySpVp19mTltAuqjpL31OVgkNmjvp+Dsg31CqDkbscZKMZhkso/DeOXAHtQW6
VdUwyDCVu/PgpxKHW+L4ffuTu2Kyl/z0Ip3nva8H3R0sea6aN/dBCxM6sMxGx5AmJYBS+zCvTT3E
0uJaAOsc7/6S1kAwlc1H+fQCXKBY9C091aakJcuagVIjdNmu3h9gWp/hZiHRwkzA+PDNtSTjg3LY
g0Ioes44LNV0sBNKMB5KmD657HqmC0eAa+DAqhCFknYmYd3ikt0KUr3GnCC2Vd+QiheHcAQ4QOe5
pbPJvlExpe/dKFBEsfN8fk44S72YG50duzDSwC6wPLcRIIBX3kc4GpCJ182A2hLYt2TMneVhltWb
dYdA/1kJiGK55hmLkTIYXMbnHbCjPCKXhDTY32VVufJtutncjl+errn+wnq66ejPVbUfXgzxP7fM
GP53NOCzPc0XG6RWAeimE+2NLk+bqcNZwVsV2EqtfVe+Yaa9kNPwBis6aFK+VTLAa3DxhglctKc5
IBMNYLgyxMowoDXIZyo9OveCq0rVcEimqJVBHXrB/7Kqu1cu34HFJ+rrdozsvvpCr2U06evAk2Er
AlBB5Xxwbr7pUevjMzhXVjHr8OYoYiDl9aDDEqMqhHZlpDaPivy8xlmZDA59+PhXhBa49jbfJj0t
20B7hscsaPRklwK7m0Vbp6MoQ4H+Y97xc+RmIBTqjqCpIvdRIKOAyv65ZrN2Oqf3gdWks/2XtgMn
9C9HXbLIhsfNIBo+U2Ys4+kVJ4DzPdgdCcJx9qkiFV/K0qF3/oIrMwlscLf9KOFG+dDIAnldsJgJ
LMO7qub3zU5gjw53hYheh7Z5yAfuahx6t5gU4AmVZaKI9KmUziC7Zu7cprKbOWJ1bxl0HgWJFy2P
/zOE0KGhSPg4NjajhAkaTareYnvrFmygcyFaDdd7hlfHrZN0hTs3IzPdn3PSy2bY0tACVtY95FOQ
+1ygbQrtV7UlSlcwtDGP6x/3CA/TIjH8Yqk7khOcWsOuNvk7eHcyFl33Cr2+K8/EO5HCDrHpwSAl
i3R07U8lie34L4Y30NXSrUSXmM3gLnujNw7Or2AENjxkvWpaXQsJzNa5Er6Jz822nJg2MkZgaT+e
A41w4QCQAWsZROCEA5gHrHOlu0anxZOqTvNkipvdSqSFEQFgdaxgqATgLBI9q8vjbI1bpMEtVWkR
13iUSd13cYNP40ajzPGdLfX0Yqt9sg/Sa9ovd759TNaYSfsaGqFR1t2FLSqrG8tUcmVuj9xiJmX2
mh/bHnSg9homSY9EnyBzrFU4dReC3hsGeAv1lpqdURjHGm1vUQSRQ1m52HT30CGocYXGOMO/m3y7
aycbInA4EHNsAzBFI4mSgZszUnOr3wFe8SU6CPIznm4S3e1aUaJC39v9S+/7UY+CjuNKA4/hItjs
wR1ZMWerMchyRIDcNJZtvBScAFp+1/HUXcwc4QxkEEJt2WgvMjWnTqwATJa6WOMNUY0ThNxMgeWQ
aaJCA4k0BVC8MUBUA9ved5YAr+cx2wzJeSc48omoMbTDdllm1qDEj9B1JfQLG41o/K88ANYPwuAs
Ln9MRZCSPKp6pWqWPsXP4xJiHJspmb4MF9Vc8CBEAAgMBPGS1uyxns2c3dEj+sinnpASTL2tDLKB
AzD/z0yE/epdBNpBoRno3r8wc3fToz8z9t6fEb2DR5BHU8D12xjyHofNP6ZHjBKkUcagXLyulcmf
aRV1zteW2Wn15VNpyLyUkJGBDmfe+vazz4uxyGIv7zoQ03ynNkmAU6w7DRSHBJqnkFTp1+327G5h
18j8oXSNzP/mO7PUmG3IysiS9wBi0RTnONOIAJTzvsSrM9mUmYvaznsHdN/JuPHl3zIftfvrzueK
+AHypYxIaa+lOAS+YQgb69IlkFtEbDobBqwkmCsYlOG31X4ccpvAZZiJYehFTp98CcfF+VtbCOjx
xTM1K8fP4XfufA/qXvrZp1z3R0u1PPzBusRL7kEBjMii0dUQgPdZJdsayTZwvvJRikydr5hM8TF1
3A+cjHUaBZZdxHqH3XnJSp+vpai004VrTzgrRr0nl/nANgKeMC2D3ziyoXpQF/ozX86LcaTrvLAx
z1syApakYFv07TWACy1mzRMfKd8q5uW/Duzt3tzxgpZdPMuqtn3LXlrOP17FNzGW6ZQtItuxXxee
tNoI3b31V3hztG28u6DRklwRlFhIdrFSPhgewwNFCGyLY21zYYnBObFDPtgoFCr0t+bSBTHlBeka
kJeVtrE50vlk536mCzuqx9nvFC+jWNBlSXGlJKWvo3AtAPv20yayS2zblaOBhue+p1FFpMtIp+et
zpxO7HiOJfPBuwz8pE7pXSzaeng4lKbV6J+QeEhkoglGpf4AeByAzWdI+aDudT4UnbgYjOm5iiYU
DebBR77GX6eg1BONnN+a8Tu3nrcPvyFAmeTNEyFWBYERzNKCUL/wRK8G42ZUfCJNdEnywi1kRX1Z
7/3nriclXm+iNyDwFlzB92qHv53+GS/oPnV4/O2armI2uKFogx+PKkIzks75w/MQuRzUr+afihLZ
9vShXQ8jqquY9Fw27rwfKF0lxCelqE8arnbjl/7vDPyji+zd+iSg9Ab6LW6c1Y2vGxtuW2B7jP5m
a14E/SaP98XIXssOTjdX8vcI0fzn4qtRzlB6QRDsGZOfj81UjRvV2LpJpEZ1mmT1HGmSRBAaqgrn
W7NvQftaQyqJ5HWtrVHL7OoPGOuJ4RjMbv0YY7r2uCBTTsFE0DCrDU+5fznc0LQ9auWrupY7BihQ
OcYen91URD9CxYmOrmFinad034IbS6WeWFyHmE6HH615HX4M5aqIOT3aam+oYwcKTqPmkFVdYy9Z
kO/KY6jwUqHrjOnm0vm/OA1Op23uGHayeGOQs2zND8iZpBiLu+oBtH7jgqC1CO41bYZ0YvNj+JFi
9lurcblN8CiDxgO7txXE2bq11cWx/U7AJgpx0/cMnpKqsBPfVL/Ti4sdMJtYG+L1u0UE7XRLI3Ix
qBvllMYysT8rQcjhkNKCnX4aCTLAA+WwxSlkOZC6xf45aaq8bx9ML0KHO8/tlnWvHteNWohFeauF
LIQsStHVIW9udth434QQoLFtUgDxrv6HCTAwrTLy+00FwBzm1S18ZZe3TEb1im7bumyMADaS4V+7
uO8pIuCqkpQpxxk+V97GTiFLUhK0+aBZRR3twc3bT1m6o/C29x+vl6fP9h74L/aT5RegSobPoiOR
5W3ETDNd768fUP2ZjmPKriEMQxemt5mjAHfrY4vvhltX7kRcocDAUfVL3kOlLZy7WupCD/RPOnG5
v8WRRQa/p0BvKwBQBQc/0sFlI9twGm/zUYHPlc71vLMiJGx+IcyB7BPYdBCnrF/TvM8sNQwqalTB
h7VgzVrENybHnG1tBsueKLi5FWIsJV09doDQbaNTtrbNQCHHvCfiGYejWAGYaWVeE+vSR0hq7e2F
z09lSTDEeUl55P0nDhsMep9Vyy0ysXcpExuacsW6O24Ti1nHMexBt+D8NrC7VMxaNiuF78/ThKwV
0+Y4ZbmaLS3wpoSYVIGlnCRFjyEsY+jw11g7Pf1WrbcwUrIBB6SgSEGfU8RCSGR/LHi2E1nWb1kF
XQDLbgUndy98n02TXctoEHP3hVlFeigRV9kKePlTCJ/AHtNJUxpd9DxvR338WsAT4ow1XKE3Akig
4W8nOeaW56wskGrWoZ7MTRE+sfrGKD17z6fKWNr/XswcrFy3Mxfrft75yYFgtPYvza89IhnZ5fZN
6eimhwZA3jIBHc487hrigHs/nbHAvqCBrwY/Z5ZVlZJjPL4X115topAVIo1aiFxcRFUAcdxicVWt
mOIhEGsYnX6wwo1tA6zXtNLqvHlsxb1/45oKym0FFbBZBSfbOQ8zr142pkqhKHpanRHCd+oiVb0I
xRmipXPnGAk5OVN97QJVVkZ5V6L2kWz/CVOaKfCiXHsttPICIQ615RPapmVgifMZ7MfZ06gYnbSc
xJ7b+K56T5HBezC9hyPBq64Y53YIzvea2oVFU5dDU8sVH54y63dgpaYI9qU6ak/nRuALPxQ5St5e
uWqQSevGcryUVIhML8g4v5YbDOKb4r6UK/nvPpsFmDLfJcDew4nTWfiiQBytgzUOHiUyRoawis+h
qGbvSNXM63V61jQ7acdtZ8nCcmMinUebMha9o+aSd2wlLJ5s3jpZmYFQEjNGRbKpE24vOGCen8VE
Yb7QKvMDNijTibXI4vvOtCagNphf9OQXJNyhCr3wbHZVOGRIn2Xp/NjNMMQfRZtSpI1pUoyVGBxM
iw/zTb+jzkUbNNPMRjdxN508aWWBx7hHcqzVe1bMYnuPJRX5NYBGrIUGp6Xwh6QzhXiT5g3vAWs8
BsvCkpmQ1pbtyJTTpZzuoMy+yAXQCkZxPtjrkEfY6Vb7RJ15qAizBmvcH46tvkCHVQdiERYahDvk
d+iyw+Mek9jbEpkt8YHF+cBFnwxt1rjhA5ftppsAsD0qAnkYK26axuGeY9ikax4+rky5Mpx251dB
sR/biSUTKU9NhKZ2kaUxc8stkTEb/Ue4G2/26w512oEdsnC5ygYrdj73o4gOVZ9dLpqZ3VOKhz7r
D9y96cMTer1kNe6ocq2yEzLgFjX/cGYaAE+KcVuvd1GgoBZMnOs+SV5Dvaf79bfymVPYOdVfZOAV
R1jOkYgY4D/L53lGhviBWjdksYaKDrt5EdWHC0XKM8tqi3sFrmCz1ufe+45Ampkfi4VbMu20UiZf
Q5ATlK3z8Nal/oDQ+edRNEBndXiXzNBfgh1DvpEy93p0QTwHpC2iUZKphDV4NLcMq8fbR6ih6xTo
IzZUg0E35y8e99bJ99Iv9zKASMod7sLb1Vg/bG8Q4ZAXgr4c4dRDfHv5LVMuQMXlJLNp2VmdoChj
tUuZEsZHe+/EIZ/4XRg8JYQpIpg/KHPksLS6zOa2MzaDqa9iPc831v2SwvJQwluA3zjZYMrmXkrJ
RvFft14qGVsQjZfW6lzKOhFJM468jDVGkZhRngYwFhLXvRN+yN9L8jcPbMO0gnF6u2zSrXAJEVys
a2aKCNylR2rr4TQe8l95MX+EPJYV8HQ53+Cs3Ls69IwGJtYsLhD+NWR107UIgbYjjbbLAfjDkY9O
7otatkpj9DS53HtdyxtGgy5P/YplAavBv8DO5946Isrj3UvFTjE/wio55xvqZFoT2RfEpM4XJvcN
H1RShrcMcjKXb0TFe+ogkW00CxvntNrfPOZXHDuqAVihXxL3zypdOWl4VMBVnonZbgQI22xnsgDk
V7bPwha2IXQQdEUAEyXOKnkR6lF4i1Ur+wZLwM3IuX5NgwNxEJpRGGec8TEfDRHPe8blPBZiCFiz
L81NOPZtb35aa3FgCZ1lNSM90rTlNwngRl0/0X844pz96ahZ+096l6RuFEMrlSMyz1KVOkEQX2+e
8Q8WVWgrelW/977oqgTxUsQFqez4ZxVDPK1fq96O81NC0MW0uU3NEw1+fQXSxUWp//hCsp9j0KHW
6tTycJ55z/1jEjrTdBIFT7G93FnYROF/Xc7kkccOT/LHY6sKCo3lOgA1GTBdlbXSX4W/UuJ78sro
gFK9hrMDgdOO8sBN2VygYnrzjzq3GdIcHGCVHOE73ZXdmurx1ecL15mmSO/XVauc32jQAkNy+N6o
cM5lCpJidt/lLwjXHUkw/86yXJOIV7tR/b1MFpeOYIzDUShjqovIcJ+kzibYGHWdpSKCTiNszOgH
0dGu40YCfB6GFGi726YpKwtXN20XafxHV/MOwdnXkBfdNEVUz/P8luLByCd6pKhe8LMsgNuZ+pps
+uUcgDzRpRL0nfthiCd/uGGrgBja+auaB6VUIoUk1zyqI8KFgPTmKI6krIbRIOo76cyl9pHFL4VV
0t1QocWO5k3J+1igCWZdDNZR1EXiQtz0ieTUisg3sZQCo6KrNstR5KIpM0Nh286p+REKNZQ90VN/
wxpxp2u6s/MdmGGbKnQQn+v2uXt4E5hs142eEE9n6yEPXO24gtsz31rgYAOx1v0uoG+BTVx8qpV7
ackimfURsBHwjoA24IiTZRKCTvH9h0Mo/zkHGhxQfXFfWlZl5yIp9AmYPeV4gdWNEwviHPm/9X/8
lzKpWVbmoEPdZTiVINWASftPapsHwdjySOT+gI0erImYMw9m7Qr7qPEWF8JdAH1cpcelGM18N1zu
0P+j3HWWHpGGmFYpzH2gFFIn0Tfp+cjM1a+15g2GA4DiWYlDKHfqOQ1ZoAii643nE8J49IJ753hF
bRa1CXhCYRAnEAxPpSl5LQWDauxXZz5RfVCinJrmeJX/TLn/DYx/Fp9p4EqEL6xHPI6DOfO5ipKJ
ZVfX46xAHPNXdL0IMt/uQy7X1aVeLWaiE+MQICol8WAb0AqCFYW+g7clK8FhvF4smly38h+7cV4g
Ba+INutOfJOs9FCEp/n0QVRoZzzlqT/SIThyeM2Q0LmXTZb0dqvBzLLO23vtcNJ/GZrI3e8qRVNA
aEyEVR/Hr/gUQGiujyDRXu0Ze0PJQ6XG8r0TWnnaWLxBRByAVKBpDJWEKtzZCnWs6Qq2OpMftZxO
/Xk6Kk8zjU9OZSIWHMrbp4cIk44IqZ6rwKU1ISBe5ksrvrM3SVpk9EdJh901DlkHwchfhdTjnnky
T5FlfVHy97Xf/GLFUPLdmDJQZkCQHuN3aSx06QWyNOuJQK9BZ7b18uSYh48LvlWPg9Newpv2/PLg
ffdapGqNHoBlnAIB+ZOKizUemt/ujUZA41meBuoup6ANpI83ptzQx/SvrgvjWti6BOTGRWzO2296
B//OPLwFXa3wYRg/D4Gj2V+2I/gQFDwS4UJJYK3+KebWRet6+cBcQY2BOPFmvTTQjSY3zVcGq9V4
IaYrtjhtd551b1PE6ibLHY8KwzVrEpUzrI7+7MsBmjmChvoh0Xdcao3MS6pyCbBbKjDCsfQbp2tV
1oCyH3ihbklOHVbzn0viLF0kEdRSb8J+OG0+aX/x0fpvNGpCmSCkW/3XSr2PHboJBwlTtOxWXLqN
IzICuGIKAspA1mZzuLVnJ16L3W2kX3wMSM1o32xiXz7wkzgsrImuVLfS4CvC+IEJtktf1Rzl11gW
I8DInwQzlTVh2uquTgF5NPHx0FErFw3mzdliaZYfqsFZY6bH28K35K4zjMrsYbGcF+ZdUzQJyrgM
aGIhIxylu+TUdfCyNNlLgQtmNkPmjmKMOpaGmbyclzurbbg45VZ6l3IBTJT9Y4DYqBMMoMAZ/UDl
iy7U3Ww2Zla1kNZj7xYMfOIr9Zm1Peg7U8//mL2kQ34ZDI5XWq2F0aRq8WsYri1161eilnIZwfBa
68v+natNGM+fZrmESwNAOO9dXiWYD8oycJYR/48r9nOuMSmh0G0EU+AVYJfY75uIMUYhLZ2Od2Fx
K37DDvnN5VnR18ZOdK47h/1LlvV3nPIQA3KTZ1ipgFvQUP5KrSCdygswV8ZKFwxAu1Xwa1UaxSYt
PsAkFS1vtWb2vHmFDjB4JrWA9JW8ZklnAkVjElcLI+SltaiPYJi1UM0txRl9tTMEHEiUR3gWs2PL
RnGvoWyU8ZtmOgA4aecaUna+dAv6LRT6ZZ/WZyl4GzqjAbvwcUjgDbopzDq0EtnBlruaUdYoafAq
DdosNFVtr2sjQiYwXzQFmbqxjAGiGG1SasIulk9/JqsIr3WJPZrNp0bY07wvGV2xgJKWjGuK7LVv
P9pYnL2tFvVirktNjt6zxo6F294OX9ksS/qh5w/nuhjwql2JJxKgYruepiYi5tX9skwZYtva6RKc
QPQpuFPUunDeCWZcGdXzDP9oSkXAgp1YXdduZ/OziHjTmmjTX2ir4QRNX36b5PVoIoDOdgnSbxbX
7DbM4C9g+KkBI6RdTTP18M83pPfC6IKqSGl+gmsK+F2lpNjPqAe2amY0fikJrfN6uEfWxjsTeroO
3TvgiVkagGo9Vi9NyOEuZBHMbeHb+Qan6UQOKUsNzqUD25hUVR5bflEaNvXHbpdnJEkgLlHXt0JP
aVUOlveWN7TNrTG3hBahInvzNleV0ND8cUFpypk7yVfn39Kt2StUiBE3HbK9FT1Xmw4iir3Qk4qU
tBdpD8mEw5fDgLmYTSC6hLnuI2DNSRbH0OdGBgUdiomANU1+W61bpGWJ+RfPLLPgDCV6vzGhUEWS
xazh/1EOw8Y42gPIo0X3qkKKwYpKKmdy5Vd3+ZtksWIXBmntb9nUENuevHbzIRpPE72ws7Qm0xcj
QH17WqowDbdImsvbeJUl7JgbgtNrftAhQbMdb77qy9/BRDhqYgW8fDllXuOSDSIfBVNjt4LY/f61
uqjXQ8krapOcHq67mnVmhhzHQzY+uutCrjlzRVEUjdmEbmBxtn6phQF/wCAyH2XwfEmyiITSUqrk
bjgqwwROml+iOA2riunI1QfjLEtbnno4E8e6Jfaq1XHWYjFHJ/G4SQ5bU5tlkGcUd7YQprFj9CuT
Q5ZxvSHJv+hogLTgOnQRbFaDlGmXVK4x5X5CE4GU4pTTjHaU83Y+m0DnvsLKB3GJxgDfTQmSeLfw
vmRD6mOGuXzWyUGfm1wDuY7vpxyjtldOmlZSxgK36Kt07dsRC+UNyGrWUW2iD8HCcIHiwtjTFwmm
Uur3QGYT1S0ycMekX9mdVl4n/+NkBlHadr3I1O0GG2M5rBq9fWq6pMswytaO/Gz8in6vJ8IC7yrd
C7+V8g/EOhskioY9l3wUrwnWpLBth7v3Tts65omLNjNJ0OZzuZ1capEv4Fif7MKZusGNDbaOKgqO
EzUPopX/jcpM2pDi6lyVkZ3v8iie3fvZOeu8mLjujnFo/6zJCJ1H9v0B0aGqTg8McstW3GClo/7S
n8atqT/UTapkfn05r2Iy6qNThEdL/SssQ7HCgjxuQn9WbGzTxfdqPlU4+ogXvWE5yb1rL5x8FCiJ
MeIkaokWtdfREcR0o5/cQEFog6seH7CcZgHZypikQAVTdUnkL49aobEkBVbLlii5oYgqeMXBKM6i
Y9RmuGjviHae4NyxV6ZrvwJnVm+AmaKM32o+dUp9/upfc9zgsgOui7Rt2QsgXVvssS67FT3Nscep
jxHM0DBpLLchNCA5eMGqz9/nvImjNlm0Pzw6AiR1aXG9rusrKQpcH2lbmkMzvKFhidmncC93g3sg
k6Kkv5cY7ZKGqkiHtqK4TYR6WlVo5vV0avvPFBGFSIpOufRUlfyao+cLvwGTKLQxdFe7BfxW6bvH
h+thXVIQnoiKnYmxZ2s0O2SZdrlk08ZTuZ/fTdbhVwunnU/1vFwR4riWgVOAbodnYJaS/GGFgjdd
Et9DdlRfPGSSzm1g7E/1+bdKZBl10+qKepyvC2w5TObvtiNSv1HhAZM528Iel0UXaomGa5qDuXR2
wVrtNGeTfEqQqj2NEru8zPBKwClvJ8oRWiNOCo/KuZe3KsAfmOIq0WlHIFG6ugMNMeSy7EfoMPmQ
qDxOJLyDStHz/201CXLGk3T/cDyE1Buvs0QplwkHEO2fNL9rbN8SGUcyKXpQdKg4UeC/seM/i3Ju
oz0WhBfyZhW+U8hNYtqQbsROfFwC8fZJ2xfAMy6M5swkRTrfKCf/t9WO6Ncgg5Dkwn1ZJj/f/+fn
jquaMOpJa6MurMnlGIrFlJliE/Px/uOmKP0u+x3nrd5f8Mrexf5de2oZUzl7aAQkSRjNbL68nX45
ikZEawy6r1XVCgOt9rcTha8nGwzEoDXugjsQkDlxabqn96JOs+UOZjsBKhgNBx93b7ltNvAlzUnr
nKZiBl4cSBwkoqsSiGLVZNk3BMXCctHqplt8OnOzOK0oeVga0DI4od7BCA9vn6J+3x84DQHSa1+V
rnVcJRqbGIa1PDAilPMT87K084AKR1ksWnQ+y9toOupy/BUR2gKFXfknbOLL9MbuFIDqfXRtvo5P
5xdpOJNm9zcnhP9sKEl5LhScWF7TuQtrLJ8HEueOtXqnuomXagZNT4n296q//T/RjHaqb0ShzbsY
ESK+2wleSyOovAu9l9q90k1Tt8K+Xu7k+7/DFCi8Dub1Y7yUW/72fAWQybLXZLwqivpIrbrF11Bk
f+z3wCVtn91I8/oOSLf8it71rHoQKFjacIwhGYQhmjewO3QuPOqpbCyUgHvEgNxNPXeR6suda8fK
kNK6e3IwqTJFO2RPpIq70Z/d/YzOITK10C0KsMbJ9kTz3bqmvi/B9Izvq5F6KgF/2ei6z5211q04
qSBPUqfdvECRTQ0rrSsMVC430TPd+S6lK9UdVUl34Z2H7ViveGa+udTZOxRgN1B6yg/TY5zKOzpU
HSqoY5+lZfU4ASCpMgZ/hXUIK1we/MskkUayvmFR/Sua4y6sUejJsltevOYFYnkg/HJfk/nn/+4w
te7PwxN+EQ9NvZqYaubW52KYLokJl8BNZhabm6zQN5EVlygvIirTxOECspMhUgtPWLi1ehc5favb
UEM4+8ffoSPYInVm1EqKmxZ0dQJDAibv2YSAr+W0HR7aQH4ZENWizJ7VhuUvEDhb0fer6fY1CmMf
vL+nkDEfFZkTnfut5CIyp6wMBXwdHGZTttXURaXGFkrpqqIT1+CFekTRJuqqdmY37Vy/dwSe+0qc
2tYIJca9scT99igRhuHuU/zoqfnYlCgaQDkwJtfVDgkxyLHrplU/WBacqpLtpU5tbee0ELSQA9cq
pjfu3T6xewOrdDmPXSSgRD3zPghbWgLm/RwlgwbMOxkx/Bd1kmbc+Y6uz4i1+Zy/JftNXbOFucnq
RXCaDVmiAt6gFcORktpvG6bu391o3K/hJ79LV6jfkI6G025SHOamhb8L+VRGC3NXmnwRxaizm6su
EWL6NZseW/p4RaDZVUsyrLxz6LWtEyd7QQfs58X5d065GPGnU9TlCyjlTGISGraYjlgN368bd34e
S8jB3jR7R+JJKkzJEQqOxXQ8r1FKl9ZnxRbQmlJ4LuVES7pEwCG7mOP2VerUf30pM8gNl+5qVI0/
9wO6xd/+YMfOzcCfPv7dGD9+5mX3OfcbgvbrWR/5V2kr0cjO1z3OYTNCsxZxjkJM7ZRKdMJMZ048
XejnlDtwtH9N7c+EKx12B7EBX4mlWXviYmAk07bdFw232b5dvvSQwbsr72N62NjgyOcnHLmAoiT0
nVBHohFxpjUPyxnWm8x8GHFKK3ICY9dE0DJm+ZidkCGcE7vCzwBOuwRZTAWUuSvSew1sLfHyziAP
V3ljAn6kdJbu9Ze+2E9MibOu0k3/+Z+kPHVUTX93YwTE+8XlaqybPuwxQVP/wOVdnxX/7ZcbKvmF
dWd2EMvxdp8qaeDMpSRZn8QbHpjYux+WdxrS9vgdz8AUg0XqUXy7vv5yrcvK/Mp4bYp9GRlYn9lg
bvet1VPuiMk8JAr1Fr2PD+th2LsZRDBIF8llPtIOpebhppeZzAnKgeU5urwSbKc1+usukcc144jL
U73HCnn9r88K9uaPBQTYm39WhHgCugX5byz0uePLi7mImo7q+kyQSXSuOWUEgyC9uBbtjcOGC6ne
UyWQSYjCJt/U8LXdG62hv6ZdXSv5xvX1hdDeXAr1xJ2+RqZ4sTCiU25Pmleo2QhTzia8sW8usIc4
ABusQPD4QXxZNgvg5ebG3h8P1QDTQ11W8g+o0mri+quE0Vt3g2nWjYpKBku9cm6J6Ho/3B9jFMfr
MrPgqFJxdBHE0+B3nhKSUm3rUm+Fgl/GWfumcrmGvwpeXw6gwHItlOSLVf/HbBq38BHOyyZN4JVz
KAPG0PboVVrQjQEjE/BapNHeg3pSDHgjaCmB8LeN3GqLIFWQKCwDQawf9nCwSV8VNXDoriLlaDP6
EyNdzueEP9wopZHGxSqUMvbBhYU6K1yzqmAzcSytD3j02YET6ZS/RA7l/0sytr8Zrr2La5wiXOGO
vaxL5joI2TBglgnv77Xa7tZ972Guc+AedgAa+PsXpFNMO1YwLkpWXKpm1ZA+IrQwIW8kK2QIQnMT
+WfinyJUWkNJFvJMd+LlKRkC9TS7xEEaxoL+u6ae/LGMq0885sIK+Pcav6TeZeeGgoXm24GTAL7N
saOIba4S6OgKunzXoaJcTx3iD/LdsSJ3AfP/HNsbgAl7uchR7fMZwtlXhMPM+EbxWJ5BfpGDWrkd
JD15C7PhQQRY/s6N48GoiCbc1arMaXJcALn+o9ERjVxM4UDxu/DQgB2SCgALusvvCOUrFRsstM1j
+JIYDfJFx/vpl0P4ZEQ85/HhQ011W5EWBDdVuqxyZbNvexEFQ4okkKceXzdFfo1Adtn383BUzBuD
/FUImor5v5Rfvf4O2aJOvpKe65h8ljc3wLc2ZyjTvryYwEsgVtnYBHM2zlVpI9i21mxGuFJZUxYX
Zhj2JpqG7ErdpTV6MjqU1j1N0wp+gnlnYAQYvNnJfQQZmToRXSKsEEJ9oyNXebwqdKHYbL+hq311
TChdYTO4f5c5zeE5hHMnsoaHk3p31SZvutBAraNWixfocu4Sqa6pzJ2fTonHnDqtFq9FGEQ7LdoA
VwV2tGq1yPcpK2dZGaQrHzfgn1LGHCszc7sXUUN4/llVjbBZo1S3y/KkeyEoS0yNVhTccfdti2Al
gJNDuMx7NI7tp1GtjlrU2D05GVVmjOoOlD7/W0bTaHb/G/zDjMZF5UTeaUHjLknwMFG763PKt7Ky
+5ZJVDQ3opUFxqi01KydMg/Tj/hHkq++E9T1bSEx9Nz0fuYpmB01EccUtusULMyaUZMhFpEBpw7a
EIvW3DeWE6CDgXBHmy995mVNiwE+2HqTurxwuu4r6Ls5isgoczWQ7C3ZWv2F7658sIzv21mqi3Az
MneW8kbiNruVi3nrgUTH5FB/+jAq+3WlqRuEB438JlYLYbELGr/CTIAVfmnbFkQJPqvzHZN8+56L
YLZmGXFcYp4EqFoj1P4He3vDTIcf6USFU7uyTZGiKfHQNS8NqDIZqVA+asDiS/3sdgKw315vCgH9
pSm9q2nRnK/Yohbn3NUO7/XjqjR3Zh3t1rTBeEZX3BaXJu3OSanNh+FEdFteNb6T11KSSvBDK3h3
9oxv+b4ydrN97IbkV/JlWQT9Vxs0GMjzYzO02+DFWOkoYvxux2x4BdJv8HVMZy+6pDgiZSWBQEyj
46ajztc/iMrQeQAXLM2I6xQoiaU6ZStuAM+KrS2ux5o5sM1tk1JTNuVW+YZ8Ouf1JT7I8m63bc06
55VxUvQulboAwNmDhotPk4jGDnHJTwaW8wKlqTdLGhVWnd2gEDZPq2l+4ZEgWaH3Oq0txqhy2IpJ
UxdTEwCovPB1t9ePrlkblPELoQAa76Wd5CgeofP5tlY39IkneMRY4gcyekaeKVhxf8peIIPXeeYt
LzPk5HREHAxxk2GqY6YYNPm69JsKcO9FYjHDhd/yZgj4iQGbZAxlmah40vNPRjbBXcuYEbINfRVP
Awvmk/0ZDrRrdH6U0EP2NzD5JDJnWUeVCgJGZrF/JNNaVpFLasglxCPSwYtx//882t4CvfD0Jtp6
ncWzRkIPWxQDkgKAtguUyR6ITok2ZcQGd56iaKW+DVJ9pjZsmDsXya+dLObXgnDarvcFcgvCGZSH
JE/x3WwjtkrhNys1QoivWAwKxHpbHX/3+jZ01Sj9GTTHSIuTDjI/6M2gQWqyEwtrw2VmF9hr1YzF
bFqvNV7oXXssLGk1y8XOZFBkn20eNRTWDre5FNB5HFwUlPjL/cSgKPbacGw01rejNuPWGOaUR7Pf
jnSlkgiZY5Dt6NfeLj8J+wj/TfHt6akbPcWLz0CMKxJeXurQ4ivSjfII/XLpTBJMGbU86qavZVwI
HIOD7L8rW7VhAs1AYbFqnVB+3TbyLrU/XM8ZrU9Z3k3LO4dplYc/pLEYYAVrMJb28pUA06zQjPZZ
OiVs6ltMG/CQmZIUo8jROGQWUs9T4NnBS/X0TKCzhHeFQ4P8l7IeDkR3qT6rHM2Q/ZKPYAmOuaHK
Iao4o/Z/WsQMEOs4ErpJOgoj744p2hXyjARKVD3wwDC7x/Zbr1rtnDrr4l8SFHwRYpyITUpueoZL
9Xg1DLSj5zcfHW/IfEGGdTako4dZoxdRiAeGZGeyDb7UahosqNphuXDQnh9m+RaEcPSCjj+kAwNY
fV1QAdZsNbwTXyHPBc9WIvgbCxfMTg1f95a+jmrQlGKkWWmyECG9KUfCCPnk5n5+v8xgY+hxp5B5
GGmriIVM6tz/VK5MFqKKr2kon4CJcniH30PkCU4CAMWUZDzJRkqNnB82ppe9+Wjid67EuPHzSz+t
MS+TX6Ua000c3BJXI4yrXhoGMgQY2MTGDMKXl4CAtdZbyhISiG0W9lreRt06tKHa5+QyxlVsBtQV
jnXQTTJBpFQcSmJjCx+gpS+O3IlIsiNp39SC+9sgzHRbEDYJZ6snQpqvA5Fvp1/0IyUQIeiqlXyj
o1RsyZTZvmeF7HGWHFe6vhTixcykz7TXdNWjFaUay/dTGxTIlyKw2BGNzbg5PpEDa11mJ2XYSxNH
kWJf+W1+12rqe6TiKRBN0IF3Pu+bYf24aBLloIFLh6GoAslE4f6GzRbCzTX/Rq9709wbhKS5zjJm
CueB4jFQacIETk5qROP7d57/1IK3x4BwxhzrJu/7iw2T0CzCC4HUa4gXitfdty5yj2W9J9/TGcJo
aAtaxk6bnJfPi+xf9vDDlbtkoQKNXsQVKEh549VIhIk174GFZiYgqEtOVVQCutgpNgcrhU+wmXjQ
7WhdlvZRmVigA+LTGBEtR2z4O+sQRUaYna+ZS7XVyWh5CSlIIpgWxqBLLHO1TK0DHQbekQEqBwS3
h5YLVKMQiSZWzAEhxpO3ugMeuCYga5BLUtmYXoyPKYA1yHig05y4hwIHiNisbkKXt8OPVxXbzsWR
Z7Dzxc2bgjDvJG3phIQUxsiHRlt/gBpZgvfyZTKKhQyGSdzMoChUHdistGcCngT7+pLIoqxwYzxL
7wbKSrvPnIS+tJIJlmWqLErKQeSvp9huui/R5gvA3ZxUYb48wEPT+70Rs+9DesmVySA5u8JIdDKC
QC1cm6R78mFC0q4hAmZXusGtzWBBeCuKTEGGkCa0unvuaTzxofmGSpMMF9bkJV8PUN3P98ECc/ZF
+kgMm6ugtVzt2HJo8kxrcFvFBV3ITGrma1OYD0bfr2MlqlUTD+n8tQYjDNzHi4A1RuCohNBm4Si2
2T77t4FJeuLLmj8NVotJkZI2DzM2Fr1TTy38WGu2D+fmVSCAEuN2yFvE3vdkJ2EP17X99c/VRStQ
MPPh8w0UkOA55wXvlTr5n30khB+6M/egOnOWuuoK8bTjJi7KBBcQ1jKthQQj1KL6/Wb4HGjREqbc
b3qjiFK2QwxmSHs1Asp8XVCVCbRhipz61ZsG++Mg9IVrXdyPq1kgC1LdkX1FfpHFIB3WJx18+YOr
LlFXYsfZR/pOWcCgJM9lLKQipPL6M5MzOEdsLYjhqXI37xX4i4iBN5c1cc4BEl7kLqCofvbypvhM
Bg+pidtzs9CP632ewuITZJt4pxcVV/oFmREavkUqUAkEPNq3Y+oj+Whpu3EF0axpq75v2U42EEeT
w75r1/wztQeQ/sb9hfSjJyBi3CBJa2OzCKGMrGbdGXNofXdWXpwL2qEno771Fxxz2oyq/Sh7T2+A
FExJcPCqZn126pm8S78bjAkKZ34jOtZdGO5owgOnpZ+m73eSMsGJpqte0LjToVkoZocGXgCQA6Gv
OtjP12PcwvtZYpJDrVSoH4nTOUV5jBGdG4Lsjk9RgZKjQPaGI3cCYGm9c3fBoKDliBQXlaXzJXHS
tzlFpOvoDNrF2y++XAvqbE9wooF3LBNkNXHxwpCA0dgqqfP4VClMhgJtwPRHH88gZN2JDkwULWyF
COEVR568furzBbmVs9lBmlJK9OLXLAk71qDcnNLH8JW225UOEJMuA38yyEURkyJJZcKSWOf/FjIh
JeNswKdA99frbthxplIrLVnZ4q21s9SK+1uBdHiIqiw04HaBBsLFGXSxlve6veGN13bPeDSZz7Cu
XGUyk9GhsUGXIC+fIBEgeGALZ8/0WYCFwqL9ik+x2iPQnD7TP7lqrgMJcqiZKRAJggakva15eQ69
vymH5Cc66ohXr3TjHtxCr01w88IDPVK3ugeZsR7LZQrROfpakjjQ6aKjOx4hZlEO0w4dRmEd9FTH
r7FBb2Q8xhdLdzIuZYZTziIRZPOaERr/dEjYBqRnlMKBiKIgwfgwHAL4EdN4tr8elmieZzzg25FG
IE57uLuotB/CDrY+f3n0DtfqdpS8Jw7+zVo89N8wwzae3iW2wM2Fk9aiqrbDYgKBDSChC5Iqz1bs
4pkaHlgW0o3PFh/3Uou29/mn4AufWyJ7rrI4sN6XTBxvfXg3xswMeWtXCWUuQN8257zYUABZh+h2
0nGRpW3c2JsZqf0/dluR4nCD02tz/aI3QNIFk3XrNA+5wIGuXC6RUGhCP30mlda8Lh3nEUFWcl4g
CnRlRIVblrw9TY17JbycQ3ol9RRfBLKFl+SUm+C6YuW1IvBm/6jLQwZLhtlb+vhsQ7qVsn6/Pstw
zx4109bgUwE+sh9CwjqgnUzb/eMpqBW589GAg3EZpFzOCbMN3Z1gIlJnUhI2J1yf1Qj/M9pZNaX1
2mFPmkZNVUFXZacQ0p8zloU7h5xX53RnVJ9pKGHbU3v7lpkNtK/QckbLeO6vBdUi8OVYUyd27sif
JB/BA95Frt49+ISP0VKXDYz824DKxV1KBJLVWSU1K2q0gc07PcW85iZdyjsKk7aaSIKN5RLv/y5I
1o2RrKqmU5a31vsniJQlwVv4RqXUL338CbICPbYFco4ZbTvZCnoQZpiS6+3bHoOPWtMei6bCcT5n
HnHqvUnYUa1j/HK4/+wJw8dof2uzSBqWsEXlG6PPw+OSK7n78MZm3tvf6zmytej/GzGTDj7U+Xpa
L+uBjg9N12ayvkrJYhgmFE5nYR7vMzJOYrgLnl3JY2hLOfEFDNZxPZsMwrIosX2lQmGKfWx2qkju
SylDuZmTYI9Dh1zq3rJTjitt4tf4aefhRZRbmYkkSw9YOpDCXBN6JBKoxCDT1YIQzqy7hgbSqucG
kg7ORVwhqdhBjMnA4xNljJ5Ypwpu/Kxpr9Hw+QYIynHDFIBqbkhXUfsL5DCAAGoQVICLDA0RGC4V
wbUUYbZOURWTM/XOnrz7jCS8lTD09g1NNK90DRPjphnjVBgrdqSGQpVwU5bhlZey9Jbj0RUjTnjf
aMx3V7JmEJPNiepeNB7+w8DEHEKQwtwxZGuewJXGdV93cbc++DErUgiwDw2ka85AmMM0P56cVN8c
kw+Wctngko5h7rr9lnJWIyjN2zCWOq43/udQFae5vkRUU77R5QuNME6PtIjVEEv+w9FSsWi4ewDw
Q7QObmWmylpC2tTpLgc7j4Nd5O4RdJtx32sK/pxPCWKC291ctdh9EbsBCiWJhR2DABBU0NfmJtuM
QhB6LYpjf7op9Bxv5Rko8X9Y+5Q8Zm41lraGpGymFCrkjtAwmwcfntEW9DptL2uxNkzEH6e6jROd
SFlH4ZSsQ8rFx8ZczpUAlXGYFAqCNnOQVwMKBItUcpGqN2bEIsPdTPtk/nfrZFN8Mi+f01XL4Tf7
NzhshIW7cfsBvrBM4u5JQyUTqmuDovkYMOmHqUe2P8197IZrtfioxDedrTgq+sNfHGbSifWG6kMh
J9KGrvUB0Hg819yxISgmBKoFSRjZEwh4BQCw5itB4FvZd7nkh7zvvCjYDKRgV5ziae3/FQVdCW2V
xuH9a33k7R6dLrEg5rNF7wBBtMo37rw+YkIZ3vDIMNJsjhQgBKycp9YBBEv/JmHdgxFwqXY1zV+N
jGX99F5zWO8g0soEKZ1pQEopxitIjIX69EU8IQev21Wg1iMZix0KTDQeT5vZk3yfvYSpCrd/ktLE
uS88A/sefSn1SO4phNDU9YHZeNeBl9X8Zzlx5zzJvJ3uu0nSLyTVBtxm9+ba2nQ/qxy7yDDd0JDK
aYug7FjgypUFsTCBsZWSb4duNtPuiMS7+X53iRPoSkn3UnIMp/Eb+b6JNnG18qke4+yXpqS/XrVD
SDxPGxgc4k9WF4DitVv7gtRSKhmv7xaqcJesEFa883wumRfxodcJTU1DTZrsEaUrZ35FgYjkKJLf
7fyU0pnNL7SerQrWEIMGKA4FMHO2XOFaOw0UxqyHpqZhZKpfvdoKzFzW/dL8YXfl2P1MQLdnEcPT
2pqeIY6KQKz6o/OFg3ifoca1uagbQlUMdM4/GdwQLGRrTwTxTOdF8iZeD5ZLeanQOJJ3OnyTI96f
zjuvrY/A5KSJWVXAXpbAGudfwlq2reST2rAOI7JODLNVrOSWc+0dzPD5Qcr2/SG5ra3c0YXvnk/I
HPQhvN8+EUyxf8D7yxbwM6Aht9ptxiekHZf9JU4J6jopJc2L9It+AEImp46c2OCM2+AkTwEDpMn/
zHRAnCqgR1O8Zb2GyL5ZJAwWo+yfMIzbYr5LjZxD/qJNCJECUkGt++Luy2Anl3YfrIxA8ulAhHFG
xrcVNuSigvCfY3DsJTYb3sq7O2mTCymxt0jGkXaHvVocYsAC51qEKzzzsp1+BaF2ZZG88ZkS9kJk
h/w3R5eNQM/2IgCg8wj8YjG6/jRQ4He20/llvm1pAh3mWCG3AG+feh/Qvuwq1rvzo7x/MCGqwCYI
HDWoR1GgK30g3LBNT8WmG9C+5GTARHj9o2PSFXTZXC/POEnUhbscPwSkFdn7Nyh7NYsTvU2Oiqf+
kFG7V3ri7fQYLEenw9Ycko6Zv78SzzbKKXop4x6KLJWRsGbVREIbCMkP3iL1TVDDnvbMuGExwNEq
/5Z2GcA4MNxqE6QQIqYFIsuOtKfLwgM4yqrETJJ5ikhm2ylkBiTbsSNUQ5dgd8a3MGvv7nQPqmo/
JACWLhYPIDTgAjnSJ/CqJzto/IgtfCZcmR6l98LL/6Ae06yXNK3mkcIgksmL1tYRJhq7iBofmRv1
fHxUgyIx0nNjSwZa9HAqafXZpFNq7NJH9jjFOHEUyTmwnh1eOQsGiLWiCKpR7NXnvqd+pQmzkJ4L
KaU6Rs0XzK4CYAoGMiakbHQd0X9E3M17qBpp+BUr4KNM+Jpc1u6pQMAFkCaQgqG1Sa16Wk5S5ksl
ZAPwiLibX25B08rISHXzkoZ5RhzQtBYDhTi15vEF78aVTDBEVtYuwSutqteRSbK2eKrrH9jUU1gV
3rhfR4OO5nEA4N8wK1E0Yp6wb1S1sq9s/7PGco0lkS+8Zn+Xj495KD0hy/pQu/apHdqS/01irmY6
MtzkJKtmNqvI3zbiSU7Ma5IIoGjuGvWyd5FgmVfVMJeLJw8l6yqHpHeAaIcoTn5NarHZwchBkL8o
kOMSvHNTUFbXJtu9KdjB8PtV0PnloOfPRLkjlwvsCsU54pCANVfhWbtSlWj7MLRcEg3WEwcWCqAi
qWKuIqaWhHpQcpE9amAQo5u6ESBgnyES0F7WwqzZ30+Og63ZWHLgRUkzEKjYzdzn2b8Fx/83NHky
DTZkmODj2fzWIf01vzLBK4Vq6VkRN801+QMiMKuICm0nulGp9cVo/ieyUeXHlmrwep2EWR3xJQDN
Zfu/SSTk3/PVA/YCjCHCqbfukipcJj/C4HKOcGJgJtqtg7r+zX7xdK3xtNhWVWosVMt9dX1TLB4W
281v98hkE8axHseTBUFlpQNa4AybP0rSbI5cchqaqXvOOZs4ghpKWH8ujvcEiFimxBefpY/pnKEu
LYYlwFRWc/1ycq1ImJsQRbz6hED82KHZdu5Vxz0bvHD4FFr/RcRvJ0CgmEfyykEg3IhxSXs6rTFa
Y4Rf6NefbWsZ6c4GzZPkGADaJMsrtK5rpIjthfmHcq27IleM9S0QhTT+TlxY07moMzVzhtJ4nDeh
OBGnh6K6sFTETWpivphRAVsovZu0jgLnvLLIKScGeMfbeDlheFXdRdmWZPm4gX6zShgM4y3UOwKj
Mt3FU3r+q89Cl6YdzDvl4WIY+VDTZm8NwUt+13XLvw/f9e/zSrVBh4bLg21GyAkM33CITzP0JpTL
ZtUHsDZmEekNGrmbGLDQC64QcL61s55rck3ICTRqtL5RJ98GmlPT71zTtOH28Biv0zY6RTmyt7w7
GADjb5rb0I1oT8CesqhEhFVtQqbd/BNB9XkkurooM9OPOdXNtbZUJzHiK+lrbYUmIjgAjVOaVsTs
ZGXbA3MvwrAXRE/IVBKDEWlU54uV7aiwntHQQ5la0cADv47gpFEfQIgoFhjKe8tjTjdA/Qp7nGja
2RfGwAjSximnZGJQM6oZ5ZAt91TOziaQUhfeCWDxJTNwOFOiq2TieIHk0CsOGW5sh0IKE2PPpbXx
dcdT0luz1TMJrFMSi84FRtRNixyfyW6flr3VU9MD78JkX9I9HaHAdeN/+mrzPzjh6jJZIcNNIYC0
AVHVcNLlu+VIuaoqgGZygdHM+WztnMIp4J8mHjanqTQVlI7FE5E77VMww1I6WlWkzeS7L/cPf6TD
Ngv5eNecUOBqcMdXJ8wrlgqnU3HRIlEPrvkD2XwTv2Dmn9xjbcpR89UjLbLZBoE+nN2MRh9TEgyE
TV6z9bSWO97VjOG7PGJ5MpDSMbLU2sjVobheph79L655VQGKhcMQ19pOOwxBO3L8CAvHl7PZMURg
4H2dOqHS+smNZvKQfVcq2i7H8Mcpw8xAg1lp4U+jAlwFgbSo4f5BrHc6p288FSwUf9385uyj/wpD
CSu9sSKG8k+hVUceLcNwHH8OnLbL+Q6wyWY3cZCxrn1GtlbgEISyG2HHJI6co3cdFgs0dWmB9Oa/
3p/d4RW94ilzDHtEkw3UARuDOMjraCENzhEcLTzM51CckpkMmLGfKI/0QyEmLP8Nj8NhBt/cqmrA
GUA6O3tqoCS6LpYpj1IjHtVZUz/+ZrrDYwBTyphus8fbmkAvkmYpTg0/qsE6jLnVYxc8pvd/MRsC
IWq8j3oceiMzOdNIDpQRHAR3lOPOrobRM1JO/KdeBEn1pf6IgTYHCNqyj15Sn99sk0ItqjJ4SKg4
sbRb9gekWSZwnNqX6qjjj8vfo3QHYKlQeK6rPExlBAfftbsqSglx3C7mYrFhftE62OW0PNIu4W7X
r108+wKXHiQ1+LycKADq8rUZL39GDcO508xZWM5OQXMf9lU2LR1BbHN3MKxFGed0+4FTFPDvdhq1
c7VwCRYsx1T4Fk5ZjmfQjDkSyg42MhfJ9QXqWBSPmrXvt5uwS62ZvAbxijbkH/40uEPFGYXy37Bf
eykp9/kI0HMMjsohwoEB3CSSHriwf1okuQOxaMi8yWbTtj003XmYiuKyzjqYmpwDitsROxK5rAhu
n4h8BHPPHxwjLE2kuF2BxKuHplF6G3F3Jsl/66GQ8o+7ShgPiPrLtiLPfqnbzDlGUklvdByFwFtg
wtbFvLAOVVXSgsi0TnbkZnfJJTbBZ1+JI1uCQHKl98f2hPRwBWiokm7ovflhJyKLVW5EO8O0jmtr
3oVsvLXsjWAZQuHnVPt/+QihbZFsyAsZmZOn+BsXt39QrlkQEZKbmEy+VJCB9LiBy7vT2ySVwJbt
ofafX+8fd26NpOhX5SW2DKPfP4KMIv1uD1ZvWdwROwIUyAUSpe05X/oJcNls9V7UwDYZqpz/QSqM
5eEVdBx0vSPGVcbaX0J4vd/gqo9+w1HiebnFz/NXlZeWUPqxGXjWGw06j5352ePpiOSKFlGb90I1
edJTwQUsxlguwsGnyGAKuWYS5+nVyspXPuz0zkxJ6f3McKaQOtSinE5S000mLCkm+hIn55lsSDq9
mcqe0kcGhd4xv0xZaZPmix/BUI+ymIvkRWXjnwUQD8gKsHvuYWmpRAgnOc/xMQ9r5LfNQSNP7ccu
/0wucCRO9CQTpBI8nvpb7XliuQAbww26oTdJZi8M6oCKMRVJzdxNPRzaLMqbaq6d58+ZBfa4f3tu
frPZ5cf6UFjZBPdABMnMAXsowqM3pXHHiR5NWXjLzCcLOvjTinp3+Fo2lmiCNgPZTymefXYF3yMB
eAUws2GmxTHI6Q+2QWDw+w12Fr1N9rywZQZ70jM34dxij+3y6I7wjtjtYDxZ5pl3yUv3XoKg20uV
X8D4YI4x+TsK/tWgufAUojwdUsLdoPuqYhUrXSWGI7CIIEzOlckLhkIiqAC7AqVFGI7kK9MCGzMc
cokOIrMBt3ZwoEr5uieWzrwxOvJDsA6LZB9GO4mjRifhHgCM5CbjrPiGcY1H6geIj02FoDGatJDZ
E+Xcwh9PTY9UmVgwlU47PHNDUXSyVR79xcVCrfI8akDzuQQLVFA43EC4FLJZ7pcYuPW5aOk6DAMd
2F/cN1rCSxNewH75XRpP22eYh01qtuCZd3zMLB9xW7HbwzaiOL5d/ETSDEGsEc0Mj4vl7/xizNcZ
FDhcEUdmq6MczZfH6C4XsCjG/mUG4NtdEtSaCVEv2X0WM8jdzeWUyBTZYHruSsHz6t10S5oRtwqF
lg7DtnLujiAIt403iUqee+8hyb0N/bD4nPHFYq/6bv7dgDprqSw6D/tfE4JXNgdhp1vVnowZiYFZ
I3OKOyKh05fBccNjKRpa1vgMblKsurd5sxBNPiXz94vu+FifjTPBKNBfvObeUXpyhSlFNNGJMvFd
ejAOjwtPr4PqfQ2Tg+ILGtVKjERB0ib0c93896EEX4/2pMO34A18YAN8j2wIFCdeYNjHu1URgp7G
U9uEhxL2amOIiCGLqPnGtKSBjqKq8NZAbYQiIm9SiF//3QNdZDJ4wUWkaQKPr11E9jkH1jq+P+m1
rTCAobzB/bjNDrhAhHvcBem+stoH7hgN2eXyoE0MTI2VEk0FEXbl/S4bBXUMcUa+acylyOMcPiW7
yHkj5WbTwDCVTm/GAIMNpFqaM4CYG7F5aU7x36PTqe/v+4koSROLVPIXwIBeuWhoBAqb6B5k28/G
tHaL+o8DLElt8PlBdC/a0G1bNXVPZ0Ypl9N5TE/Ppu04tsXI9xOzbHlrmETSxojC9Gw+0dQvS8Fu
60BTP3maRyFc1i/mKt+5X5m5XrNV/YzJbbYX5QkdgL7STDaxuIyAACi/NVr9ta/6cn64L4JqhXiV
km6nkzUwDM4cexc/NW8Ugp2cfyL60giY5tTUpOWr08oj1K9wzLbVbxvti1mggMHNPOr2rXg9qYHN
C2Spmx8+mP5bhfp43f9Nr1ga7qtnQPf283RQFsnYsVmRA7Wt/aZaru8QnvQgLvA87yUeO1gdo86D
XL9IiafcNAH4caqSr2YoxIhVmlMbXufaW0mOGR/jcqNLhu5aFwpxDxWBTHfS3eiX/CxPrj0rL3f8
cstJ2dgcHEDJQ3GfSgLNM9xRTGtnx73N5dZT9MhuXjULg6l0pxpe1T1YQ2eeDkOWYFK/Vq7GYGIE
uzUuKeuqNd4c0wt0pBLE0iV0GcULAdKS0iEwhXhk9i+2CMUByvOz4oYKpUh1xPaW3+FnOZgLfm2A
A5CaMqApYVrOtkuCcHhKNfvTkI/leT0tJttGTF8NLqcGPofFQVTLkcYQccQGuMEJzo4LvbbyXL2w
wZlRTYvjPgwKsIwCZb4zGvCTfRHOuCYaPRzYtcfmPqrp+E7e5Gs5GpBTaKqXkCAN5FaxhNx48659
afEuqIL5gCFU7pDFrj/HPLKtz51kqo71tOBB8eM1fCr4n3nIBe6mSWNv7lrrAFHjdD0Qv2AThnn7
+AgHa/kMpvtXeZucnH1WPzXd7aqeF/M/5BHVZ/Qqx3Y6Wi7ktOn+z+8V6rf67aDG+GFNWX+L2SzU
+ub5OcCdKnreyAXvlZ4gNVoRCo1xhdYy3GVEiK91E3CF8MLPg+rEotzejU9nw2+qCduQ/y/NeWE2
18MEzm4Hff8J97AXTS8j/7JnmMIc0jlPcPsmF9KvedfBiQyFUEb71tqzyyD8ZZ8RAXr8Ejs9+D5Y
5djcQYbQczO9lzWQsbx2/wyGwMe3/8rv1lP1BJeRJy5zUhRQYwdbw5bCuseUnGbMMc8Khw4VaW3V
hau0zVwdig1ueLWmiPA7oC1hlg9IpFkSIdfxd3FssL4XTPbepqPyO7LU3wRcd45AyRJD986pr2c6
i3JGRcdi+P3zaIpbB09KayZLapf/UdAoyJtPZqAwjise9mcasLHr5An0AV83y1BAS+VMeBrwzNgk
z2ECdVsn3HGlc3vEHW75S0iEKmG33brSZJNDPJJgolu6ckNt/wyaC4ovPi1sDuukvEbs54LkUHel
BFNOdafII4TNxRnsK1wOKZCOtWT3/hV8ObIds5fP1YPE9Pbi03lPnYz0YMBfa/XTeNIGm0Jd1fHC
Id9BTbsHGaunwW+Qt6xx991oHra8oXZjZI5vrpGw5+AKaJRyR4SdWe5dDBw//H55KOD4rAfBYbVl
QkyLP+v2aF8r8sZNW1iccIb/wgNAJPdtmqVaEeuAnI0VWaLhzVWT1mOC3Y4WYrdFiVIwzQk60cHm
PKomwArpskXTJEsMxzO5Jfvx+ou1sYMIArKJzrfSK6CXlwalZM4rOnS1b3E/5hNdBfkIqjjlaJuQ
GgJNvkr9cGqtbddaVyL/UKjnljDH3u0/2zf6zyhZOEauBxQn/xixrkKa0NA5fG+21umXGirDdi1p
LUobPrOC11GUiTKStLX9tJTQO7QPdCq3z3DN00EXmo55TVWiThnzYQ16AZZxPtQVqs2EeslaNQaV
6ZqWJpkFNDVGnDL9O3PoD2sQapIJDmugU4RsP6fk0PXxaXcFXubvdnXfGyoDhrQyUGc9K4J3NlS4
5pAkxxTWadKIa9aO+pRediqiH+mCdWBYTMkeSfg0xAm1oeJFoyNBIqZSyOJhSxznKcylPDenKzDX
zYrk3dYWGnw5y3SV/6C9BXxTyHP+xhKcwHsDNR6u0ms16qMBrjAxf8rxwwJ44eeG/+YiIuJtTMOV
LIzB+soPnFHNGs/MQRoxf8ZnIdQf6KDzcKvu1zwfV/+YFGxxNsYibD8NF6cjZOXlQ3H1VKLlV/8g
UQjV2LVnnuMZeyu3jx4ki/Z4jPgBxi/M44U2+ErkIlvk5WjAirbO2aPbHm0783sIVuao3pVCow9b
F3Tug5JJO/3TlXXk/e8r/L6razX6/yOBQIm+tTrS+5WQP1xUqH/RWJanB/K69m+Tpb3rOTclsWXx
sxXxUinz7TT0l9fC9zvljcXzsFG0DCqS1tsUdOpZSKf564pKJ7LwvkIOHDu9r5g3lVXKV0Rluc6Z
RjA72mepa4ZBC7tlPHAuoeHi/MfYY1HInNOBwGaBI+HNaYxlVEF7DOrVzICzsPmmOfv/vZpaCkhx
ikNgWAtpAzIwTegsesOUjZUUOcY3iC7mAWGFTQDvOr38YttwcaZMjRMAsfDxkP+HLuwpJGTSSs/B
M8+xsPTIfDwXQSA2S++0iXTjsrAvExKyANRrQWIa+Vs6x2iLANgovkLhJq0FZHDkqCPVbRuAVQgc
gJdoSLc8bgxoBUSTSr93uoybAJGMgiZAY8auhhDgvMfyjUTYBznniXNlkPPZ19B/QZt6X5xQDOOw
mKmPSuH+0xTSgIZUdZDlJ7SpfVTUkagts+QGbP/ZT6xDDbAzoUyx7TeuM+WINJHyXAgonYUY1Okn
0VQ352tjwWgNMqSNAmfFwy6bkUnPhHaAPv7l2KGXrx03kl0n/D8k6RJooMFBengdO2BS7F4psXzg
fLFd4HYHHMB3uHF/xswzyJSg5kRHBuU52hpMWJAjhBDchlqKXK0kSCqnh4Om06y9nk1+BHEqIcJp
JC/EvRglRcJvo3DECRtGOfPWDGMQwLHsSOa79sJrmYFUfE8LaHR0PqxdPR56dR5qF2pJPJ7D//9F
1716v4599cvi6ygjbmd7ymS6Y36ImrEfxkIaI/0BWjYXTL68aXR+Bxqwt+WU+w9LnfIQUU97lOdn
6tSqtFCAUCiBny+UcWCNHpOBzjzMYr1Qxf5YeL8zxaWA9F4tVNiBKacOFmYLpzVTIXsYdl1HqeBH
jnjFkekCq9JFY9ulh3CaPcMjEulb+2PefPIBGR2/dMUEyhBfVc1gm844iqnEnutFKQ4Y6yjIEbWp
VoPXdw2wYjRHnb1bPWWLuj4BtaEJA4Hs/BoZPCMP5i4IYqKa14mpc+IwpD6YUpPPE3Sjm2B6Z19y
A8sU81lwpM3TkDSmECUGDGarsiA8nikkGMlCqmQ8Av5FQfVBOWANgJLrr6oMRFp+cYoJ6tbVituA
CufYcJq/5RrJ/8qZO/ipCGlmtw/pi1tG/vb0wtWHWSbzkqPhS4BOb1JWkkYU5GFbKRL94ZVqJ2MD
Aw1Q6+GLhyQS3jVL/do+KnUQcxAljYd8TptfLQ6irqOmbxJuWbUTB7RvL3BJ0VCTuHImcdqZyU7s
LsuBdALqqtSnr73mfOBK6BM1iijGvf25nSJG/LVBrpSuC03f+sVXOLRXMDZrJGhv4MwKDv8H0l8u
mJj0SOUTFsLmM87D78gh8SlINoiRri8dUuYIVUh0XCs8+QBhn70CWwJrG3unXfrw6avdS1ry+ZJh
Fl2nSX+SmDnkuV7+jiqeL4/a6q+F5Skj0mLa8NbULqZcDxqgBeZakZvLz7lwENy+rn30dtL6oNKF
Mvrzt/3uXEw4CxIez9OV2jNNByJm5LfIUscSXe1xZcwE4+A8BgsTrrdPEx9tDdd7RzlD4LYRQ0dr
/NAbHL+Eh4p66pHmkOmA1Ntq92ClZByR85WVibJgv7xlFh6ZbxBd9U8dJs0bpc67ErekLZe1y+KA
eDzYCO1kZYPeDl/qRkZq6dXlBJHQlszZyS53qJQxJAmm6kswZYXt3HbXjdBLNdSTlnyFvCbwHsev
3FiDVP6qpQbHYR4bkZ6Was7kDk1WHecgREp5KApDaTb80sqY/Bg7uVOhrAeoWoe97TiwIl4SeBnO
5q/j4msBk2iQOCjQL/s3+zC78LlidM4f7UIg9Blb2Yg9e3qc3Ne9zt7CD2gQ0yLtEDJsk72ttAAX
pWCjIhFPHf083rhppvdIhUKW4Mij+eGJp2pKaVeyYZ7uzq8/FlMR3HX191/IxApucAp6qRWk3cLA
hkXHma29nrJEOPcvx3+1W5QYCdmtt5m7C8jSwC0CCfNTDsKUlcaHU6IwI4BsjEEEIMLy3wNqsKck
yna4sSsb2t1fYqjfHfjGPbkcCHQYM+mG4oZxlqOe9gFiCiONYYFDyIUh4k17hyEQQ/PWfz5XrqVc
AfPz7DPJ8ugx1laoF4hX3FGT73lz0iv4L3+0SXdCDOcnSZrMENSx05jYMqEz2ciEp8O0ZUZzINo9
Y10P22y+AGy9UASJYcz6Zvx9ife831GNYkfPP3s6PxTk7XExyP6j3QuXEoCXBtEPCmnXhZTE7u7B
ZJPh04OFF8WTGc+6q/AUpIWYE3OUdMZDajWrlz52/JhyB4oJvJ2VKK6zh/HfvrgaTDuxz9hHztXJ
u2ZhTvc5qh9Ji5Z6g4CiQohwyhB5FiV9lRd3kGtwkAMQGVJXcvhqwxczg2X+vEhT3x3K921+MSbN
/+RqbuC1BtI4rwgaZrRzhCcOSfn1rLOpWnMw7QFf1xhUomH5QgPDR3IBPQ8pjNuHGuGtTe9A1BoX
F8W7JwWLOUvzvzOIrwkRAN9uAdpXmcc3iw9MsCEB7oZhu6/PkPW8WXqH6wJN1EeFAl5WLoA84suD
WIHBM823LqhOIojkc0pTVWGqTGHkxUduXFPh7PFhUamRR6SAr+dZo3/ygLxV2Zl3p9RQCOlrUKVi
DjiKbv4DSKerbB8b8JmY7qo6sWa24A6CAQTZVl9CHVNoc+gCOAeBjaSOIisjuNqbeZ0ZOMRzZ63s
0nCjL35N+zq+SbDIm3kwgebVyC39T+FRaK6dEsQHPie391FvwKqUqjf/RuqSAjPjU4EFDkyPeyXC
rywn2jxREMczGtg9XW1D7qwb4hQToSAvx5DnCqg5mWcwCp3Z/gpRl7+ElyHFRtOAlRigE5Ku3t1H
D47yc3hyi1SXU3Wupz/W+N2h9NmketLSsSbBMRG/9wGPSnpeVdzbyoRYaYE2ZvvPhaNQGMMbf7jO
w6osk5uuzUUIcu5SyyNczAWmCi9+ImP+MnTiuwk3Sx/CNPv7VbnrAmIuSw6+SKGO1Dl1lCFZuFPG
DO6Y0vL5SBS4O5Smll4U3iWfITl9zDY+b6P6x9fkQ7cR+k45qbJnK5nXuwzNt0K2Tm5L0P0ls+9v
N8GNk0QgDuIIowsJGdEQCxKLAnB1oNtVith7fRv7AjsT+ttmkrx70A2xZVLYUujcs+pI3AFRvWyH
pGun4okNatm+T66S4cSoNiWdKy1esmW4aFkemqyRkIOWau1M49ktkAjORwEBnyZ5+H3plebnm8S+
5+OLjOlwy16qslVhQa4GnnQVwRQ39yOLtFtYe4rLkS+rkQ8dZEkS5ReMZ5FvUWf/4MP2LsN0LmqX
UizLKEZNU8O6UD8avy5G/QAECLnEEy3UBr7nHl3mlMy84xiJelI1nC+EtdfqxkGBBE4juGlOIe8b
Q9yCL87JmOXa6UNJxCzOPJgFVKDb7VWeduN+ykelXiDmq8jZyJ8U7wuXeaIAH/ncyYQ/Jhl+jI9V
oXCsRx+gtWdX8CwnmHH0ITDbMmfTLF97qffBZbjo3Zw82Xwn7J2D3kfXORRaHHLjn4nl9saCkFAl
GEQMzE4ffuQiPgbX1KCJO9arEQtcxGAQNcyjaDWk8b8mVHpSU2a710GiW3YeYeE3zGqEZhW1z8Ez
8QV95qNy9WvWwPwQeOz5JucdizsuyGyu1HAs++AuCUTSNWcnWoU5mE8dJZnjvEqgxfaEX8TVaqcD
4RoaZpSYWDT/CvfvjgbYWwXBvo43AnDLxV1We9GB5D3inDt1QVRSf1ZbXM2AG5w9mAvCccY9u1jn
Y+d/5nRo2mDSAVp9hL+lCzKjLITkyQGkPliY6Vycos+2M734F5ogNx6wi/zpyZ6xwO8zUDtIMMk1
zjRoSwKgi/6sCpSd7ju/+fKY+ulr9tN4latfNAQ1RVlCHB8AUPjppdWNG19X8Ce3wuX2B1FqllWx
RuUQD7itDt0XDerYz30jPQxHrcYYveV3azpHwIp016J5dhugf6FC132fvhH6ZPaiFnd6PDluU+BS
JVQZ/7lJpk4da8APqf+UnQ1pAOGOKEVnokqJ2X9AX0x6HVtQ3KcOn6et1rn2JweDYqvqQgIJC3DV
vFyGrnmidsAoL27ffDvs8hSDXlDJhhe5t+4WQ2AYDduWwfdWsYh36F+gl3veOsFZkkFosQ5VSwTX
0R7BtRqFNkWfRtZTTxlqAqi7IvD0r9pX5UKHdrjrIDhZRX3dqbVSXrROg1Epp6gIvtj+LVwb04FA
7+y/8vDZ7LbeukPV7CpcPuc1CJxS79cAdm403N/hhTd2gy4P31UXmsY7zaj7w3X88GL8PE4S5Ua6
D/MNGkYH6IyaolnQyXTKKvxApLbONlm/cncWSuFBDvoRSLqM0AbpRqXYbTpNZ8LrGrCPnk8JJ1/y
xrG6p7MkIgpwzs9DjKa7RZ3C0Oir36w9F7zAnzc+hEnENIcRImZzlimlGyPHM1egF6SNire+O8mK
Z3wabqVQq3FycF4ZlYJntPKKOsUR0IVTA6Gk2xTUtC/zCdc7BWFPBzJ+TFuPfmlImO0SsKAJ+1Ja
gYJ2kHD+rxw9QCtT5iyirouxIhr0SG0mSJHUmRIFO3cgzE1hxnmO5QAUD6op5mh0JWtPqNPjnNKv
g+7yqLNWIxKGlNip3k3VwggZNC24vxKQquhZfKmtu+rNfVQ87iNMFkBV1pWgTwiWdaiRa8i5Ph55
0QYmr0w5DrhDruconwBei9LYdeWClmKs6enqW7qgooF34jRRY6v/tJeNbMy751H9CL3ZJpYlzGS7
3AZT/D1CtCoJAMiJ9c3HFJE2W7pcMt8Boz4+RA2jJIB1J9fSHdjnJACRAbeTGoUcDW5yUu8YieCB
gZubk6+PoDC5Mx3NHRXtAtsFoB+C0FtD3Ht2E6AqXO+TlV3c1fGb2eiu5Y65XZ3ruBKar5RU8VEp
zmCU+T7lJBmLeP5vtk0FYcpovuflAJ0rixXAkifefm7D2g4yIM9rm5siTxqaHjhjwasp/uTFtc0g
KGpqirsk2usDvqmffSEO1zXZiMuELrwcrinQ7vqRRC3PRbhOKGp+8b+AEzLzdpjuhz3Y7M/yHj9O
2m86adON3Qg3fZ0a2EmYTDEWCdwtg4f754IKdQxAbFnEu1tHe4C0gW/oA6v3wSY7s8wlGH6d35kV
sVmEluK5qsEGd7t9QblAKJ17vLAzNtPQFPCcTSziQZyfW5x0aLhKvL+oJpbLE0Lz6GjLoL/SkzFo
bjmHzNZzlsRvSnv7QYOeurx7E5f58v6gc0nrTWC5hVHxPL2pOCpsQnMSmTS2AxzTjOQX/hdnCCpI
wha9p91W4n0ao3cjT/W0/C+P2yJ8lJZ+QcbHqbS/FsdA0jt4GVNtEySNHsBYtl1YBUt4G+TaxPDJ
5NdeymCHYYId5iRZujgiDDN77jFvSZfY6qKaYxenhCwigod6GYBbeRQ4BsZ+z9FaMSOSPpMmcKO1
PkYk5rFRvR4OAUg2tTNS5aTZYaJBxvWbyG8cGx7+O9AzKtS1FkGkWvb5t3Ql/0AZC1R/KtfxKXzL
wWnrF7rpyO/zFMvvDSPWJinbEP3z8tZQhhAd6pxWFxpo9F38sQ8wJqMqQsdee+vYPMij3v0MD4d+
nwBH6Gwh2uEadItpgmj2/obI/Fy1JSXVJhNwcloJhiz1bh/V+fUiSm6JvenWLv8Aef6OSsY/nAcm
Dkc5+QsMcDUrNbwQG0ATNHFfljL71sHlWFFKF6Eop4Hhjv/Z4QnOLq0muz2KEyvJi/jCtKxSBYPb
jtjibQbjRmZRn7LdLYhnEbOP03yguASLEqVzzUfce5DunFfptulvJd6m9DviiPCUS4Jo4Hguq0yo
EdH1apUnaSP4W+I/kcOvLuuuJEYW/degQoQA6kGWMEaLtb5zaWgVNYdvuvjaADw+7ZcqoI6mEa7F
ts4Gwy1g0DX/u1q8wwuEINHMFNhR/G2bfKhVJlrSukgURfe2pw3Hvh4drKr8c2YgiPzo5rlLlKWg
ZUal8HNWYSwrV3cJqAe/7umxMqkhgURW9g+qXc2n8xikOzbMiCJ+X+wZHi4JHdlEx1sd6pZ+p+L/
Tgxx/2yEcjELz5PIsU07lhPPNI13HkgOHWXn2EvRx6rjfazIrgY8MIATTXT4ZHTEoPmfQtS0k9FW
kclYWHIKocqURYMenL4JqcNqW5OjRMc+rLEuCz+KGaqGDtD3WyeRFd/ayFUFDkyv8E1lYue0wJ/H
VK0FxlCIyyjMxTzcsu8EamPtn0KFYGfIVmhe+w5tVjta7Ocu/Uy6e9hOVn84Q8Pwd7w4vBDfnYgk
MzSeGcX0AgJbGo4VlEp34S2mXsAZhtVHLtXOj4bwnRbUsAicyuLqHaONWOgi8UswBvp/fxI6ArZS
zBKLh1dNRV6UTmuAAO+b1L3pzJlAshRD19PPMgFpBAAletdvHX3sehGWrSkDvrFgxLy3sOBITEvD
7dZk10CgaHY/wtozAj5twPbDmUc1c6ot4EuJ09diegHGF+4AdCVp4Wb0sSF8o9XREXpq0Mg76Wno
acoeKLcz40OKxSmr9gsWgR6f2a6bqTf59mYzVPQopfSC0LiDLkmyDEfMU5ea3OCszaBgHVZU2zoj
AveeIdUzwXMkaQoFx+aqEY8FycHfV08ACtkF0tgx+kHze3cBvbPrOsIlPdyorx4f4AW3vmlG71BH
yaXsIsRzzygYcK/eVJuwDo48p3qyfByjIXxC4YgtxGRyQ5d0XlrQ707+2+YDMqQaN+DJ6BQSwu8+
tD3pJ9qItWDXm6eo22BrSFPDFYH9ZbLOQr0b66KEJT13PaNQLMSKHRPz52BPy7JIoURCGcbYWucA
FG0vqXBljpvw59BrOOB0pDYPJmmSxc94+0mslaMwc63YkA86+2+uDtzz5uUQEtD1SCuoogDpTAIq
wH5zQASIrG29tt0OB/qGPJfntkhol0N7/cW9QgWSbpXZMILcqc7RjMk8p7wer/DFRV7DUs5Pvlml
4HKc2o/wo9k72JUogGAw2a2m6+eTezE1rU0+1fNkVevJyhR5RfWZQd/16HNGB6drp1LVLd+BJUPa
JX/H10TjFCupD2EcFEWmj31IaNhjRKDJrVuj1jNKOmiHJWmmsmLvbS0EY4fYwfavipb6SNZrdAuT
xtzr0KHq7CEBmU0yTBnyXDgzLvYRR8YsuhxNRC8m2d4gjmcKplbPU8mDMaLqB75dt2TQJBXyhF2I
8xuNjT7Acni/nx2C0x4798bXpLZN03+z+7LvwRcl3iRoK5HZugKauKQyeCugMFsg+GMwzde5RsWm
Pm6PQr9UDtiL9cbxehlIajexVw+OqZYsE37erw3kHqs8dWgujA5bxGCBEPF+9H21l+Jjoz5Xx4X/
JndLWrnIXh/I1Yzz80yO5owyqfzQt9JuuNsV0uRiVhxOWY/2VNE3fIW6rg0lyjTuCY7NOuWlk90J
Q4OYymrRmPbJTgPjbFnmBaCmNtZoCVshtH23Wi3EYGodQ1BnS4Bd1ELpP0UEK1H9SUWoLokludiY
lutSs0aG0lzSxLfCz2Wm2CmGvRifpWKA8bom52/2Frd9cWeBQ3EpLjINgcdSZbZYYlwTGcxhckVu
6pge0dCyUJqwpHhK4uFQH5dGaVRQowOs+3utEcEUbs26Z2ri/ixOHnnSVy0oeNlZh8jNHWnD2h9B
flJ06VnDlWSvz0LgP9fRJWW+OjZqqpkSPamwiVajWbe7ZUE1lHLnPTo/LLe00AXfMPFTtFJE7J9i
ZflBoif09fxKA6KpwqkaZ33HaF/GFH52oLlPRuvbkqfiQJHeiSL5AXDOtRD8V6dlLYgybyX0+nDS
k8zBsdO/o+L1pWMMb+8UcjzzMtep/iTB86IBAmg+WV/BD9Xm70yyELO4Hp6AgGxN7OkV4iYSinPM
U4K3UB+L9bH2qyVNQlW2LWrK5SbPCPx+Pi+3FC1Ph6W5bM5uOQJQBlqOkoI670zIoe0EAxrwFrzH
zVq67Mxtp+Em991NW2jE/B7oFCM5Iw2guBm8/JYmwmkThdOjB2BmopcOovlXVU3tDLzd92nDUITh
OEveu7WOiMSW+ZJTMHaxpOmHMRLuDI7//03XSaUKYO4VsFEjDKeEfsFjC8g6Qge7DjxmnHS1bGdQ
NV9EtwI9hu+sdiAPMtRgEiaKXC0ZfbnkANZ1mig9aylhJ5JSE2sZf0CMqUZ2NPodNBwxt8lBbj4g
sGES/ErqpYQnDvJx2ms/Bub+ia+Lyafi0hKFL4ZZDKkPHdpTM4TLNzG54QNmY1/rWP9Vbdlr/zvS
GhQp+SaneFUc02Z4Gt8Q2NYYC42PMpk6rrqJ4OGg3yWtS5msepiBeUDCOL+IK+4ebUBWho+Wyhmf
UXfAg0pKbNbw4pRZkHhWGblxfMcQL3OfTzdngSLV9QEzqxgTk+wZ9KCW3y1DCAAWN/BiahYh0iz6
YxXcKLKnd1jEUTQq4HBweUu8un7VHvVxSzO4WLfc8dJT22Ce1y0OutRs+mTj4VR5/lcjDjYTDGcl
HL2Gzt7e3KzybS1IE4QeTYZoYaSaYG5aNgP4xEe8hKtCLmSgteAGLg4xg00BeMZItQNr2b2erYTm
NAv2wIpr2GG3BR7G6tLQM0+X9N64/jZGpuA9JvHDXxK4LQHFtK7QFOK6PqHtYV879Hda1n1shQyW
mGCV2X7/pV5E4UMlQ+mxvSnKAv3DYkSohGuNcp4WoDkYb9ZLL/SGU3Pfl5HbgkDYMramBpIeS9FN
yh4T9dxGdHsWMludvF/P010/hXPahC7LOUh+u1G6sYJ+wiTzwzA+a496n7MLqpZyFI5112ULgX87
1Y2UKNwarryu1052bGBX+29gAwiJ6IeBzwqZKR36mUgw0tonWDRi1C68Jzhv+NzOIW0J+Xj2uUm/
mSl1/3uWs0OjtcguTndEhO0S0YIc8yyxdbQ4PkYJ0HE7LIrn/RnM9BhDfS2M0Q2ydRRMlvgMR/Au
W9J+/UXGsdRyI2HFfhOsanhyq1vBP/DE0+fevi3GBozAyJ5oCtITgvNT0tVRx4Yr6ECfrBhZMTR2
4fX6u6pj8p6f32sbu6b029TR8l6zUKMGJLtMWOGJ8nUrOBlNPjOx6lmAKDDN9EVJ/+w+3K/A/p0u
U5RCp8Yh4S9njljsSXjIhgpHk29uiP5y9G9GL5YIx5jauqmQ2xBccUNDC2jOi1JOMJFm97h8hwxP
IuKyornQivJwGuBlGb4fyACSYX4oZJOk8VuBo6vX1nrap6f8H2tmdRxe2QFVb7IITeBUpsUxz/ek
PwxVGWD+Sd2XbPpHRcsQSksn5T1BN3c1DMUyzepn3sAlLP55LIBUD2mwSsCUJ6tzVOyKJJ4UWfna
HpLHTk7BKn9nHTepuNRvzd5OPZ5MW10j9ZMuF2higwPLvtdKF8fTaejMNo+9WYUwenwSgX+S/siG
iTelSxfWG8btOs6ZmSgT1DK3pYx+7/P2yPaI2hc4e/TFuheo32Dz7ViYGUqBbSZpdUJ4auzXESb6
ZygYXe+0Cjio910p6Ekc92C3BApHwh2HkBR5PMJm6rOFnJZDqB0gQqCfKkjmGFBSvQvhUIzgJqWl
FzfwfSABqjl6GcA3ugI61nJK8EUVpYfiOovVXUxkEPCgzRLwxBWV2k6mLxlMeiH6+FTYkf8HWZ6p
GtGRVSRHOsWFPU7jOAJZKoxtvrR4QNOHepWsW9sJly9gMTiOXybXoeCXzMiDDMO0UHFqQEba6vZE
Xp62lpyH1ENpC4M51DsoJUgoBVdaKq91VVH7UWe/fKgJVdwZbcvHJTGrlfgFRxZ4yFZk+rGz5+aW
dyj51hU6KGLcqkQZ3kH19fsiWkxgLE9gXRJ0QyAVtm+ZWcOyGiyl6O+CtzPD1eaqC0QmSAYVtdES
y8aMlqwliY2OpgYhJjKW2xigasHAokeJjqLFOfgQxv/Mb3/MxSGo+IvW0r2NP8fgIoq0H7Jd/QQv
Q030Q0xCZIXJzGC3mSkao+VtnAnPFnLYetqx6UTcIHfEBbWPWsqD4QCbYC/tz41ifgzkCrzqHo3d
pmEeY/2gjKx8ltXLmDLId5u1+wNRgTMyOhIsmejGbenNH+1USvdmgoAotmfehfWY9b2uXbscwfJ4
gvbWI73ouMrkTh020QlQBcRPsV1N4+9Xn73eGM7yH7kmgcGp8N19xKo8+d9rK9qnDw1NG3XKwplx
goEXEZSL/kk6BCviB2qDnZg7MhXQSzu93VT31gZCGyS5Z6hmidXW4O0E3ePXacwJAYBbbFMYx6fZ
76K5tbsPveuLnKs+3JeWYiuVoz93JMR2jISSIMIO1vlJUo58B99kgWuVvEVbju+kEDpx49hUPqvJ
vESkP+cTc5UO93foQa2ZsfKCmhFFKGBfQEchHU26jCmN73cXe1w8Nc9PIFPKxCIvPPjD9DOPo1qb
L9m7RTRg+67gEEkD5Ak3AC/c7sQz48MKxlsutnzi9QMro7DyaxRIoPbZrqzmLp+KeDa2LO1gTRlU
SCDqHV8QOFYwlR+PC9LiBTIdWnk38+x1eVEvilkK4T/jtWvH7JthlG0rv0HuzVBOxoccRePQX8xw
wUY+6NSHBAiSP1R9aL5UO0mtIfjV3s0TmVJ279pppZxkpSJAVEFoi3AIX2w27ea+dwJWLFVCAbNj
MV2CFOxJsO1Km76b4d6LvQWbdBYCPMw5mLbO1jLRbNdYqgFIDSe/ossrp2VBVzm8M+swthmbldtY
PBPnnVUO8TZ1clLjGa0/L61aegQVHviRotaYbHWA8oFJQDqj5XD1t62EknqdqEGerOJY3/waFsAs
CvidBgFGK+MfsfTVuHU+P9yN4mfsLrBQpkp9TwDcfq0mBdYE4BPcdGJb8UF+lx+t8bkno7fnTsE3
MuuvxXZr86Aqqi+nYisnSfy13gp714MivKFuIajsXfrWie3MUo3uvJ7+W3IPKBZFdX4Lb5/DgPv6
KiQNnh4cXfvS4u6AbHfDt3PINL1YE2MKtgFU5iPToHJUQWkZsiAAaZy6oAv2iknBAolIhPas5Gag
N87DnroVD/0VP41U8Tkii25YQi8OoBJKWSg7EeQU9NmGw6SoI0E6p/vV4kq3onx1t3wM3ZfdJMJr
7anumjiYI0iMDH1CkXpxGXukL4QqxOEraq2aJdUOgtnOHcqg8vsrbU9ikUfL4+wpkxDg/4ednfEu
U38C4PKrvN7bEZ98MyBx+cvcVwLBKwYxQIafGsEpy9pl8N4caP7LrCqqMX40sn47ya97MYl/QiAm
Oyn6AVRaSKR2bil9AKD1WAGxwaEug3x3byA8+rSqTq+zGXD4CRaA/pbrC9M3ngvhaBDRwYLF+R49
imdCRVjo/Cma2BUJDFtDSs7dafopICGRo3Ug0QQxBkyvFd+zHFEpKVXWwQ0o4BlKx4ezciOJZpym
br4Zf1m58c2nWLanR1ZJkJcy8WL7o0wci8voGBxy4SbC/MwnQmKGY90dodjxXN1gH99wO470pmL5
Pri27Rl2/L/0++q09Qv4zFq+uAeJRM+ZjdqVEIcv9AQ81X+6yZYuJTvgl9iOgD86iBSF7Fy/P4u0
hNvwCiUS5U6OVZUIOZ2jpxRyD8ZX4nhuwOMK7kv3j5e+BFoslReTqW3ox4FSDfUh6g1/7kTDLU9n
ZJ3VXHUoueqLN3sBLloqlgmV2NXAY51PRdHBYe53PePOoZe/01WmctLdbf9+6x/LkX8iE77q0HVB
JNJVpl2zp10FHEDnJZBQNpwZmNrwcTdneoMBTSnaAYbpmVqxh9qB+iCaupFw73K1CFxm6bpMu3uy
/32QsIqRgit0IeP79RyNZSgcQRUVZUdwoUAUa1G6i+waBbZISBz1bgX5KslrVyDHecifPthgACqC
Gv0Hz0DEBlg6sgLcmy/bcVz8WOfoYFtBTqWOpaxduokmHuagsvxSckhiVuC/zGLyVNQFTRsj7izZ
5xxAHqcGXKHJfK6GOuO3tuC6CaOY/NuUS6wdtKcy1HithZ6Fwl23ozQHdMD/9lsZOxqcoBTaGdkB
7rPjz86Pr8AcvJ0lEjD6B3LxMClD5l2MvaImvrJA+QIClBN7mwq+n1EQ0Wli+sSOdsdzFbnsDamT
URK8XG8Sk2yg2SYql6VCac43C53FaJqdjmkJTxDKhfuliAdwpRMuoo3TYjbzLBB9vckUo6KRWzG9
yzzG7jdJ4nwJ8ANcUWjju52+nCB39OVeAcszQybsLIuCKSlBCR6DFfwO3ASMCvMk+Q7NE+lFdieS
2cFvszE00Fih/QVtDV6Kyd2zzh+kiVrI8tKGqkY1n27zFWNuS3rPGCm1lGEhtMDMNo9DZrXtzokm
a+Z+g8O4QktTtL93DR3xqwMvHrE/9L5gdkLfYr3ajVlmriwJdkBIPrvhCBhLzRzaWTWt4T47OO/d
lZjZD709lSMLW58C3eesjNZz8XzmcAovQtz/Y/qkp+CJxAoXsF/iwk8pPkYg5amSxUrtkzX+FoQ3
qXpdxk8hmMDn6ezkdYMTWaGE3kcleCQaN+YDj6GpX98B3KUhS4sZk5eINMs/ItZOKAgGDgD/OHXT
RQjTjwaePusvtumI1fO0+/KqZWig2WRPq+Eep5Ce6naiBB7R2N52aFa4+19kQRmKu/o2XIlcHKOD
mxKDvI7DwsbjYpqF/hhGvDqq0ugRmt5RVA4rk4FNxxZlymrFez8ZxTzPLLP2vSSE9eabDtq4FGv8
mmtQHMH/WHKK7r+iJ+hH0Hs8aWjJjZV4SNtjeHgxWEUzSf/JswDD8OTQVa6NDjyZL7wguwc5amaI
p7AA6LxC67ikJOmnY3teRSr7a2SUG72/Lbnf2hPVGJX8lpmRhtlo9e+B/69i6PVYFWYfcgsW5sXC
DF6220b++Ueymvi26hP3u9MGjE54G93r7WDG+Qv6Hv5UxSu9NJKz/8AmaMbadwrren3Ehq1WZA0O
y6X8xtBZeTWrAeagE0fQw/Plk7ZbQqcJ5fekQQj/1XBxn/rIIPv7bougWGREWoSclRkrIysoKYsV
DzTWtPZwh+8f4kI+1GvSwC77/JOz1Qy9qa9digJnOP9jjsfNiycADX1n2+fA0Z9PJ/FnDoH2BP8u
mHbJpeU1byFwHtMkEpeyeZQ34Dv7jcUTu80tNCgiX0umWL83llid8SL3lIyTR57teHDbGkqgc7GC
M07pDsrvXfx/+oh5dnWDzQgPBCw+fvR0RfV+gmWruKZACNcVMZwvih7wkHwEzGqwH9t5BEK9LTh5
Gs+JuAI+qIZtTyvrjyx3pmrFa2WtwOt6HX9H9IYkDSai9+iTO/Lbzpor/WByQKw0OdkHPHT6t/q5
07GHEyfEusqkFrLr6zjQGKCqhQaQuoZbVmSP/lQvf8jOjvfiYfG1klL6nNywA8TBFWZXkE+RQcLz
qz4C5ZoozJctiNqJcqVmYciFeySI1trS2naZ3dHoYMXlu8iE286JIqyIhYxflG/wRS9hiBxD+Qqh
pnaOjI231/5NdQiyXkTN12W9gK3HRF6GF9/NNfS2a95/h9eJt5krTQUSHNk2MWCwG8f8y+j8o8BA
NeWhNY8/hUG8yG0GACC8QT2e/wDMD5H/XOPNckDJu+/5GN/75UF+z0eIUPBMO+0EojNxMZ8hRV6S
oGPclnH+FSCrMmq2HJXbsJ3GMZWIgUXtn9TcLItk5QRFGeiyT+4ooElzkExR+3L0Yl0IWfU25/TD
wXXpgJEc/WjgQNJ+2+UbnrhCVOnZqIenonwwUGkKaXuIHokU7TQrp4WeMJsyHhoXZcZ5I2yI1fwb
MluIddvNFMRGq0BZ2gw9uGnXADHHBLcn+5XHtfwHWwY+fFWEoP9wrCDsu4ZrxkJxUR6qe0n7PtMe
v9gZceonvyZZk5pZd04nhnqVcMo66eN3sKACT8/GTflzkfcrR/dWEn+ixNy/fk4SYsTIT/AKXCc3
rWJy6pSjxATf2n/GH6L2YJ+pERL+Plu1eJsrkMHoBqsa5714kPW5QgKICvmLKvIK1huOy8/HYM23
D81CkOMcmSKlAZMjyfC9ZwqQq4dULXQgSAxLsNpqEarbs2jljifa851cs4D0lmHbk6TZJdWlYA87
5q5CXrdyn3cT21t8Ocs1lLbeJeysBEpVMdXzn8/lkrGcYyXbz2usZ8jqWLCPeiSVRUhSvQkvYVeQ
j+UO/1Xi/arrTO9nSxFfU1qinE0o0pRNO3Xwndq2hKMk71g8sioK/bYasLfM4EFUF37EAFlnFCG1
cv/sNsAn57ANFd4U96I6NGRSNOZF8mrzqF/KfPlb5t5BTd9JAzHuuagbc1gdIF4krHsK3Rgtx9QH
E70mC6/FMidFUYQdQq1qXIBxEXtE8cNzO5vqnVcBfmpH6tHAIIQ12RFWi0oYadiVI1P5XoXv5aHD
QvqaJKCqs1o1tx4ElNC+CGYddY4bJMoJnpTczOB/FtBD51s5xqldgc24D9zMFq/HO6wdQ81XnJ2f
kvVVkJgTsqA/GgEm6+1uThEReTgczb9IkTUFlGaQEjpPfClmgIC/uU0iUgXwOZPWQUopVIYz0Vk7
TKCpEEGfQYoMWTsJa0jRVaf1qhOneygv8I1PBDXHoub7C94+8e+g6M2R4OEdILCe+gjyt0/QJPnv
IvAfKx5DQW7ERzivXdTZq/5wrTD5n5yniePnBgRi3cLVQTUyiFuIf0U4f3vGMPTrzoEgWsR+uO5P
p6DLg/GX80z63nPjSPGcTooVltUi0QkTeIevzr9XP2Ess3NdUH+7EeP/SAvLQAK8U5tuCulNoa5k
kQqXlfniNByS2eYA8Pg1Kw1CEeYu24MDK4fW055/ERn0YnajvV1r1g+VunJKDO8urYKRAK4Al+21
Z+SgpQ1O0Szr3sYF1GC+egFOaUfYuL/GMp1sSIJrSaFVh83Sndoe868CpOM50vWyp/WhWEtZa460
e2/ti9DjfnTX8yLZDyIQYgWFPsEh5tIWGa41A6IMXRMOVNV/I8mG666Duc90w/EYN53WKv+ZXdJ+
mAwJHIN5tmlbb6GEFoRdscANySGsDgKfwm4Fingn6kg3yRP8Rq5yxU0pZ4vPI6iYMjw3fkihfN8G
xAmlKviEAiG+HqmHVLe15zKiI1lpaOAw479ur/31AzRa24+xkz9zmkHhwRrLmYF0bElMwRZamq/7
coq6FmQGYia9wOIVDyl5l79if+WD5ZVczQMYeQGs2O/eDzIWKSxQXLTwry2DGSaD5gLMeoxCZbPg
6JmFI+9PUJqkDDXklTfZrLLn4jXwkiUoQzW7V3l37eRB/SW87C97ovUiFoO80eZhtmyGxpI+pXx4
BvPa7UxRkJ3t9/mtIJ5KrvvdnChOdxyAluaMIqSnljiLz0NiWsFJIuRx8SPb6xle38VHddXnrX/7
ZaI+6Nj7crvpylV05h/Q0m+Pj5XR6rCy9seITw9gRY3Byr4/VC3prSLbDzHjCWGLAnPjEpnhnh7O
JGt4myQjmQg6qx5PyRM8GojQ937wM44hgSThp/Blg2QEqYvsTaVJXEZ5Tp6PdemG2laIabj7mi50
//b4H/83jFwUrvOVPGHPkLNtwBXCwvtgY+8wNeXkFyIWxZzyzyU6pzaMCi3JzikC5yBBuAT9irjs
JPNBmeEasAulN+E1gRvwK8+YDJxmRaiRgddIl9tq0gQB/RxyT/inTbMMHX7LkY9CIXwUljxa97pu
6Exh1uFYlE9/iP5A2S4opZJZQOth8EErgO04XM4srUy8psu0Pkvmx5Di33rP8inbX0Hp7IyfLsXX
f7dbvgRNSvv6Te2Y14YEGC1s50YO0uuKj93v98mRyFloNtXwoTX5NY75mWrI788bQ7MpUfaCLHNE
6Neo8XhMFby0ZI/yfeVZ6or/wZyh4701gfVZynTgkJ90IIAllE1LJS7WxyIQHjtAgK2mqkyTGGDa
NcqPYSZbvMxtbBagMO+T16zBLhPVQo5q1qVTnUNNGFY1J3fs+P4sHkkdRVac1sfJyudFwDsXaoa0
QOgSriRfJNkBXxQn2XXk/hw0A++G69ZpCcaclHmNlHcuObwR4MAZ/iGQpiaj6KY+W8Et8tq3iWd0
jTVXxx660Xo6Bg9WR985/QTfpmTDQx1WdWQ7RXkt9zC96bYKQ9q4GMPqyfFnMjvmDvLKGd5pHhI3
ucZs0XbUuwimGewG67cWuGsU+cm6HxPoQhXFnnl+C9wHaeG+dwTiLxc/ah3vdNa1TvtArD2t0uQM
xDInqNjn+9wWZCvEdwdK33R8Nhj5oC9UoVyA4/BCYuYRc/VI/mjNQiS5Vl6Ft9lTIJaBOJ+pQTyP
uhG6SLduAq+rmFMIKtxnPXtrkEbBs9h+Q6yC3mvP9awX7nQo8+2mJuCdzAWUosZX7aLUucH7x9b1
o7fcwMaTUPwkE7W7WN7/4aHvdi6YYK0iN9l5AR5e3DPzjmWPqvKNXnDYN2CFzeMLvKsA5VwY3GlA
wdI0okwItjW7VhnCM1eP/x0c/f3NRXVX9/4YdCh+Gi7K8uqqifnsRxY18ciBZyrM8L3W/lFpwgmH
HFkXBNbh//VNMYsRisgjhPMRZZ79Xs0IedqzqFcLr5XbPvfGHkpIPOTlh7mySoigBg7uqzzANjuC
52zFasnhIXQs1ikaDUQHNYmWexonCkV/7zP1xT5zs94d85241IfChzNqSOjwgpr7DZ4H/iWJIXOb
q3ra8AZ5yzyLvZSIx/5lgE5iVAeIK1l6oZd11Zxxsb5DNulnTvAne0aiMd74Qm9td4fGtLYjCyq5
rTg19/QroK4+sl5H2ZdAcO9fZnch+MAxhKRq67XZjyAUPfkjYuaMTDmOP3djsols6WRysHZ0rxZO
o3YyAK1k+rpPrDYhsfv1nxG+JZzfoS7czZC2UYoZ7ShIgUlAzBJ0qfjJCIfj6xSwYd3Ap0cUUr3v
8ugyyRwlX6WTgZsXyHEBPvZV7Xc2yhar0Co+qpY6CWFs5rmnWKa9DxgLJLAv9S26ViBs5OPdMQtC
HVfds9V6LZ65pGhxDEV/b4nthYIbeJ5sADSfBoiBvbh3ffpr6sAJq4Emr6i1bYejCuzUvNjF7pdi
gz3C6MVe6Gw0bQUiFui+OCDPiizbI2RzLHFA9meyWg0Gze9xuhfwvUBF5RnYtovYtQj9PfUYiP67
9phOv4eyhgJs1KmQgzeEK/+cH6LbXAxMIx9KRqngO2txKi+i1S2P+HAvo7E2Ds0Iz335CbVUpKi5
V3iLbnEsoDtk2zXOvWQbmQwOdxJY8/wtcCeqEYUFLE8SDuYU1E+1pPUVSComW6jKCcIwMOgFdwMk
K5gCBUOGcyAgfCHtH8qbBlZ/cySwP3QAT4+wE4UcxqzJLfsdT2xC2nmmvspktTBX9n4senBGRfzY
rza7SehYGZYbL+4KIYsDSq80CX0PPDvvKoFHwTTxQPu6BTliegYguUfGEDjPMHyOQAu87/jByOZA
vp20KrIGZ3BiHcdrcPWOr0B1G9ekd/i+91wr2RScGHQh+sSSDuFLjW+mDdqNS9ofbawU8YHLekng
sfMBj9rRmgGJIGZkLybf4bQUYqALOFfNr9SX93hpZZJ3EM+fOctNEIfRMteJaR9NoUHvbe2c//Ld
GJW97Z5esIzmLLUoy6UZ8COgUNNyPHeSS0pZK0Ce58bsSgb3zk0fEAz94MVp7Dgi62zutwYHLWU8
eBseoX2D0TmhG7UU77NSKiPnA0B4sgpv/87DDK8eUTTNL5UnJoPMiZtJ2su4xGtdxbI94CXCVuUS
aWSG14o48bXeWLvl7t7Mu+3bjc4vjeKeJ7uVMRVBOnYOF0ESDUpds86gYio+9uYz2yne+0gx8UsO
AY8A4GsF0PESLmgCgQKXcKd0o1XGbIMrWwl6yWq71rbzutf/lfhP8dw7zAzgG195v+jGp/jKnG9M
uhb6WYA9IjHJMebMu4wu3D2wLPJJLcpfjuDYrFMjCSsBJpXfkXD4Cbw5DBv+SdBjzfOKvHDe34r1
2lYLM6hWzroZ9CtJ1Ez9pcA7X38Wu7zCXpj6AwwkLVK+r9TLq+KKa1C1dsIGOps3RLTVAxfaTOzh
uFl7TRQKpu/vsmT2jBqjFM62VbU3ozjEwElqR/gaNgHZ2MXx/sL0DTYSAnu8iXE20xtilyQ0XHYN
gYItcYx+1007IIGMoFP7vSSN5BxB1ZAxRiK+A7opcxRG5IHqXcQ4l+r4T343mrr2wYCUG+qV8V20
OWjMkJMkOAz87F4TJJRuTLETvyp0j16Fsqnv5HuU2jtbNou24C6wDVL2vd6dQd6krOSOOSBzGKPD
/OB6PyAAjo8J6lqMzonWefVskqXWrMupmJCZ25I3AJnuI2KrITVSx6tZ/JHu2CF5UC3PLDOxhDgF
7FPLM4pzDHwSTc6FZwh5tzQM1KzMHEd7yUlNblSrpt3Pg+hk0m+JxH1FaLtAJR6V3HrTdoOJ8As4
3slM2wdG3aHiBwbbMU+y4q6CUX5/twyl+tf7F3NjjjPr2lTYM2GhKwM+3u6FZV6B1IvqUAQyNHIW
FsnjI1PRT1EhIRAr9uozMqLXfOagQAO/clrfmvC/FvdTGpWCQ3tgejzj/GdbF3b8HCa0ljRj5Wmg
z9DvXNc/jwjQNnTEACt3q8+a+Swjy20uVVyE7f/LwdiQtnTFV+NGXhYfHgNbESSBqC0F6xH0Wa81
ER/woFmhIepADrjwHuhIGHP8oRHdQCWEIZx/WHwm+zIQgQ9Vqjh8/hZ5LZhWzryhgOezb8WUBj0d
7lhRdE8hQDK0xE/dSXVApMr1JpPjCUPiEsf0I9E5o1SoLzlRGJelT9QmtHQb8G65Dk13rHEkjrsZ
RJNyGUk3CC7BJ7LqXOT27RO+nnLlQgoWqWujusv4GUtSVZ+tSI4xI1eCzmyXrp+BsocGadoQMkI3
zM16Qud/doFz/35qi8TaCoq1w6VfesgPF9kvZDGIODrsni6EcUAgv7Ls8JrsqCteWWF2J9eEp6st
Ra3euVfrJwUUfQJU7xmByjiyzHQ/lz/Zm4CZc3NLFfsRlFoRWPRmPL+A2nczvAIWi19EjmNe19C7
v1lDmvxMMdg9cuaeJneZjikdC0wEDGGCoYXQyrJuC+n+NJIoUPxPuCWsHD4UJEnM3rWig31rgYzf
fbyEkUO6zJdxXCK5adZlDELFRR+Z/XZFE6ozE1jvVnHsSiIpItcEp/dJ59d+hBES0BIvz9XjqdnF
bHCMK4rokRVWwc85F4wD2XUjQcb2pFy8HVjDZxc9MxKBKp5yB+WZNeFRl99O/uMegMOX2KxbBExq
BSZ626TRuHaH4ve9GnXvdeOWqIsXaLhsmAkWPzPiMdao4JbTyWPcxoqtDoYELEOwIxdz4cwO0RUG
SAHtz6vc9XizGfu9ZE1mpSeXt1iM//eqrYXOFe4q0ruyGxulzVZrwv8L+QrrmnZ/ekPD4h5fbrYz
Qgovzxq9RaxiU4cPeiQwRIblJQzUrPYM7fCsSkw7zrfFtjZBqt94jPznt3UEl446Utt1wktIUWlG
3NNJlUH91eZtMFz6MkHo+NrPCaqp4tmGmPRX891J3Esyu/hibiC/Q6nq6jA5GvSrXuIi0Quh7Zwa
k3eMXkdYgzkd2kW/XOTUmeVEJWKYTN/F51PxsF+TEzMBmu1jJIHNq4RXmFWUfoHXIEYFzFW0EHGn
To2QVYp5/ZrKY3IGq0xpqebwqjBuoEnteig97Fu68P6fHtiir6akksMfSW7Q6ALXhh5h+wrwodeu
r+tX9pMCGNa6vmaKsXU8TYBRcV+6k6zofqFnebflD2vyz81Rru8W6A/mZSNf9nB9TYvCka7W/tsE
F0fddiUPfREp5sWhJl1tPdsXthvGOVUA82KikGX+kdrtiNxficTe7jPlUfgmbp8a1Kj8UTPRc/1m
ZZyE5Lq/CKfW5tN85NRBLtyJpQvi8e2pV0V7JQHI4deQQt+fr6HWY3trg6+w/Xc96eT62gDyJgiz
LrINKtJpnluHUZbO89BAk46W0JDbliI5OT1hq+uVwPN4yiIYymwLmqrcZNbh1Z36tj6E2mOdvKO1
NiV//vTxjrAAMQxXwRtBUMKZpmobQJ/6qS21vMYjY+mAtFvE0jvAva0cWcGVqv9uTcObViU8S1Ud
Cyag1Ua0I2hUIZoJG/OOTNJZaJx7Cl4Fh+tFjuC+w663sWPv2VPvlPOs/PZDfo0TclzALtT4S6h9
dnZLBILWOqTX6Xi+j/oT3BxIxTruwKawtUV9sfP05AR3oB9popyYCQLPnvTLFo4ttvChZexAPGMD
B9BqrolgfMHjqJEgOyPzZWQAf7TIZbxc0xstZfigGrvv3Jv7TF4wfioleJNNmrhgqBRWfZqQAw64
TEenur1iKCRflqizGPNaYFTz8piuoQbtgBmFT2lYJtQ81uIupNqZFmMMBKyrXOG0tri8AYvRpyFU
lwBlmeVNCo6bd58KwHX5z4eBK8f9+xjnM9AoaghIaKhWdE3DhyEZppAZ+YlpnNYaxONT+XcwmkV3
u+pFzs83mFSbcJn3nT5AWOl/WEJlPzn7Ug4uKCMXpRsqnwlUREu8Agq5JH7rtXaISZ1Y9Mqwo4bT
PTT3B8rPEPfMsNBCLqhkW3Vx2qI2V5gfoy+fzzDrtFM6GvgATZ/e2zVjOZFSfsBBAgrZXvNKw5RJ
d0HdX+ijOM5GxtxvBff30NJq0wTLDxWqAObY5WxhJYKISotf31t/ZPAJY0HvgBw8qVcBjxjOo7o+
x5KDJE/LMlCKiLG1ZmgdWxPQxVhQMtMcYbMAM5Y5Dlz9tpI89bIVRGxLpkpi66U39YccddXhJDuH
3/8z0pneQX8NptFwAvpbrZto+oVqHRHTzPv80FzQQLyfMvJM74NeODcgBtoP1Sg6jIWPk4caWRno
PAJIPZqwWsStaxtgMHLmyAjHL7bFZaJ6PeHu4ZBM83Jl/Pzeyq/b/LUfQa89zPd5V5HqygC224YE
Ruppl8+/f7Eh6Lb452LD9Y7MWkxB0+2mxVdQozqaRGd19U9lcvE7OmKVURWifkAU/TEyRgZ7gzyj
iHiz5+TyflGEcy6Jqot9IUqCxN3U7LZOBAeoOruPGUe2N82/018L/Xzr53wyFaHME/E/4fG9Ulk7
KhBLeA39KF+Eltb1ZeSgtRluX5lSXb+Q5m0Gs4YI62FErVCjOUWrer2t1WLrH4yuItGra3cGDciN
/VLSbx19vCiwuon0vLz9M+W9xFBec4Xj659MsuHCHLrm0cdv5UcNcyNCxK5GX9zJVPIgosQ+9jnB
xi7DMFMfNEPy+tHYnKaGQSyph97hR1Qt8n7gyRn+dP4aCJMoFgQKlJGqgzooetqkF4dGDjJORyxO
APZCenMEdPMUDdbia470y0/PIUgzZ4hrwr0VYwYQC5Suo2tC36LJ/x20CvNtiCx2HJnYS9iIJCDE
BV9N5/GXf/3Y30CxmBWuH0jTzzLzB0SN3lW1HAsS5BZ/lkZX6vVLZLcUK0g1LWKLP51T0rFnEhGN
bhiKQtr10uVhgjQluP3xTblxFf/+ZD0lsuA1pNsNXhLoug5p47VHNT/m0PXWeOCSoVnZNXm+l/rI
0RISU4dw220kzzGv3gvG4ph1R0U7qPwyxGgXZQuY19yKIcglaZKFTA+TiHhYczWcqzH0Nk1B2Mq0
jYYzviCk+j4u4OgCXcThVdwLLD2oyvziFx7eG8RXMM4BzfzUZwMjo6A/h9p7kyhxOCOycd0GsH+6
17FaTwjfKuvJL2TvJ9phPFIvsAfvQKg2gIZWaq16ZpjlI8/FcG7NTVDS7IxTHQj9dJtxo+2g1zh3
7i6Xebt2Cb2mxEvOTNkPA9xIBcm6ecqQhEC8Rv602trNhCP/1ihDTQ1Ew/+kTnln/0NkGOXf3bt6
J2TrqINE2KsZncGRNh+Rzb8ofOZ9wr1LLV4dtFhzXxBttTxuAl4Ut2A6MbxR6+ncmanQ2snceSmv
Jwg2fdvmnu6hL5x4+lF1rZdqQylBiV2UOoH8rU/0XlgNN2PQXhhg3S8tPk3Wgjak3drFyv5RHV0x
amvXoS3MXhyzvKJXB+2xUJ8b0wp/EPdgjyqW9o8KNx3lQ+jAAHJQ0x6vIsto2uNHMABbfvfM3h9E
Cez1mn11uw9wjCa5CPp/Di6sa2vaW4iQV3EN/Wrg0sKwMlquVXwZ02uvaS+UdHwRQl0F6/tiaMO+
4hx0KdiJpP5Ahg0FT0E2i9uf+MAv1AJkgC161ZiLW9oXfJ6jMN7O8UBR4Fb3ljMRpOGREnCcZH2Z
uBUuOFc9px9FlEGLw/ho7sWihbAYaIcfGrpLD/IsESC9pbQYmxzq534a7At+yfW8V6zqo4mjGikq
F4FWVmP64AHdNUe8Lh73lgNi556D/42TNKRr5eB+lX68uHpjgJm6tfHXAXG6wc6RlEB1QPs65CfQ
m1/Skp7eqw4TisaoKAPgfXnsdfDYtSdcnQ05tktVd3MNXckn+If5F6EQZB1/D/wCkZl7YXKDmv5B
I86hBIVAVe3/B9di/UevSo9gkqa7id5zwxd/5kFCAcH+HLB+Z9mS2+2cX5gtFBcz8hjzaG7eYk5E
yFIbDi7VJd7ylAsb1tqhUMxgJmAQSicjJfSs9ptkq3kJir5vrIDKNHxTPz9FDrhzzSyxjQvuUzuw
TXYRM/BIzinQ0vOJ+ZtYDiwtTQTnn4vraPyvfM4Vov1AowyRbbeCtXnHCuZPInJs/v48zwqkKV30
oh7u9RVQmhWXKfp0hvS6CvtS15h8XdiUIIqu/e+3wyWEjKlHNhhRmRRfttMbMFnFXHIVTO/bNsIB
wh1CcDJhv77kU8P/GbnZTxTUZj082hbM6wxvWux0Y664Nln3Ujoiu7qOgECARVuCCs071VJGcDhm
VgwhfMsYHwt/YqWkBPWfrz3ySqzL/aJsi4LJ5D0fUNpHYEGANlFfKjK/QAoYhOKxy9Q2/xU+Dupi
4SWgNumJyA921Mr387GG8x6KnfuMCuCg1Ic6l8nGGh0UpW3A0Ybc31rF+9JhbLkY2p0ibphF9mIW
EYYzI7O64TJJsVzuHadnWxeFD7Du2X4HCjVsHbzEMM/54M4aJJ+0nRhAj4ogcpafyaSnh7/Yfx4l
CWcoTxFkqANRxspgt7FFAJWmGuOeDeEYOCidAY390YivKwXOnh8HurFbKSWBUKU+vIlncEuBs4xz
H6G5t5vLxWJ3xDe7fxHIhLKsvpim45mcs/zQogfhOrhnDTl+ay38yuspq5hkhgWW5pZ+Ii7n5133
R+VmjNhSSOGe7bzgLmBOkDXihWGdTogbtKn9npGxanWk1JMKd4XPtkrq2Z3TFLfI56TmlMAmtp2N
6VNRniT9giRESmhvK2EcWDzotDL9yjdt9zNdBwpEQU+M0Lf34ftBwjAQp/uj6LU/LNJaIIs8lxnu
sEBys2WU6mOUUf5+DKmPAwBDBqH+z8YzKeb7YB9cb3sDQh43AJqe5ejxl81qfMn4dvzozcA1QOa7
kZEiRdyQ4UBC7KhiRTMsFSGFPU6w5mmLYSXXPm++23NeLWCUEYbglJuA6PYmH2vy/1xZFP+TKoC8
A9sYjvdpbFTCdVpYO55VXtncr/+mbYx0MfvJJTvHN007ACJsVFNMTi1CPHSswdEO2n5Sa/Jx/fR3
czX89oidTydUuNzCIIZaF2NazlBODBDqjX7VCehgSXxMmUfUVzlwIiKrWMEfu8EnVVVyU7S7Ge/a
G5YVmjHyMNd6qmB6h+ZSbxpVyE43WLanWM9x9Xl2IajqylttBKgQ0MHWYmuxPzO6fpBQdQOi3zDP
ywhfi44MSorXTxkw/U9aH16nzR9ciu8j7jGBe/EQKS+ZQ1GqQXveK7spL25ccobRjKWCNxw5Tj9q
5wozti03c5Tm+cmd4zf7kH6NpH//RHUIzupubqI9fDkxbX0oRxrXCGH54mhxJ/mAjxuq97ARDaEd
+Erw20LBY42HkOItwK6EWd6qdRoJ6JpUZxT0e8W3QtBRjoTtjzVphTtIamxwJ+e8loXKgSp6aMZY
o6vumJQa6o5RrkdME/5Vuujfhib/umhK3Hd20VOIxoQZLwnw0pMsdq1xy0OnR7azaIBSO1mG0n/T
sNgBYWIxO+Ch1uogSgcDMmE0ub8ekO7hEFZ0MB5iixASCljoEa+4RZis6viSF4jbmy2FtU1lDEQF
FchuTl1K3PZB0nYYDZBocMIckS8y32DZwY57soHDnS/bXF2I9kt7UJ6boUyV3tTtS2e19IaHj3jj
vV8qXsYBsP2emc0aEEtHVLTO/uNHHmIAqozWa351S8Yuyva2zisFGfFuKIQyKNVqA31KQdSwh3cS
+/PQa4kIBh685CmeMiqhRSqKGhrSscPbTzsiwWpD1Z2mEYE4npoJXEc34LeuwatGI4gQb8oyAl+e
/0U1wpALZxZfeJM4CTpwF31jIa0lKa6YGimhzGNAA4NlCuDZEXg9MOs9Z6sz2zSoXQ2GrPnYAU12
AJn8riGlhn9+7juF4J9C5On+bhAsMcvDBo4e6lTi2qtAlnTiSSipsIyW9qjKLbaa1wT85AIn2sA6
6taXQg9WfJy2RRbpVblBBfC4dkHt91egiX3AXqMZIFko62/HlnxzFvKRFrvlkJ6eGgUP7hjNgdAs
XVlcPEEkhVJr39c9Vh1dekC+AHFgWB1ZUCWrsIIxQ4hgkw8ANsS5i0QfrXErcYgRs1IS9fFw7vu2
D6WNvufJ/qE8/EJJ/eb1+PmoMTxjWZQ8tdtAvLSMsYLUQtyBpil6xY27+rLvyt3uZFtBD82D2he9
6nLjkOsTT4bnuQXv8hRBoUTsSmxAsRtZWnJA8bKPTHSi+BuAhmkxcXxRMsY/9Pn1ahitgd0gktIZ
QLyj9r741AjnwV5NyKf7G8Gdp4isu7AoFROHOxcxZv+bDtKyJemFK7RLnQRt6CEFTuzC+5h9X2c4
KjrVctxJ6J8Lnh2BesAWbEoT4Mr553wD8mzuOUwY4Z1S2GPsdHmZShKyzRTpOxRyDNS450MnqTE8
4TMEYwc/4JbazkCUPvWLF9rKUXIE05SkfipNnDNmJurray6XRvOyxz4xl7vTot3uzdYuLCZAK4jA
abF0fIupq3qHTFxjHbv+9+46o38MOUYY9tK+AgUEa3cO21imT53CwSnOb3pjUeDL7ydu+LxIA5DH
hDMKAmKgXtcr/84A+72vYVVRAhHqacgXSQ2vmR1sZIW+gSAI5eInEEhXAzlY3VQNBh1HAhnzMd5O
Y4UOZmE7JHUPRBBxR1nH2lo1KlUm40l5bdYq1fiaZfDSBXcRHA3tRptiZD7nbpE3ko6YHyJWeO2h
KOBwDhwj5H290bw6unKbbf0f7iVdfHXbqVA0/ESauccqchRbe+e0RqLlMf2kTV+QUdG8HZAh9Z8s
WICMtzSOT3Qx0BrTQgTpGOijJilm7M86CIG0Eu6AMOykSfRusbwQ+UZx0lncsv/QB2tf2w+2h9dG
hQ7+Gt6NP++Z7lzmD1IxJmGJ3Wflfe+XQSS0qhJktL5hJcaRqB4C0wR/m67eptYHatReR+uSn27e
PWFck163q8hKsHcJNboMZUFsbt3dbaZCfKiH09UxTvxK0yE9Y+IalJokvFEpHzfFk3FjCn5tkB84
SqWCEF5vJtog4CFPoOZarBMFJL5I8kLCMgKLGrZ9GTY6jQMFUgZQ75815hkeG2KqYqgxz/F4jUCb
W1YJmF6JRtIMtbfapJcJopI6I5GWccYe76/1X4sVJFiXK3hgmjk54zEnnNAMIm8MIA1QdHK5pWOA
1DeDJt5D/EtiX+HsshI1HLfKV0/DKViN/zXNS5J0kKPQKJrw9khRUPH6BF+Bwdm8ODIWV0rQWSFD
XpmFz+9i0w2xd3saReb46aF4zwIHfY2MKLWhiDhGQpq72E94X6QMxv6/Az02oG4X6j93HnYDQH5U
leIX7z818ZR16Le2aQAx6+u50DEI6PfBlCebfa6gNmeSOjCXubpdYvwb3c99qWoqJC6QciR5chrD
mpfBS3cEsngt0UpUKeuhbsSgRbIbFdqegUU8G361sSYP4oN6FWAcPWQjcrGkvJyC81jOae/OdLse
BgKEDuujPlXQiJdbWqwMLWwVyRy7F370byGGd1LWbajXSXC+V+YRptlKoiEfxiA2Tru6wGPP01e6
DNSesOOy2YIIOh3PGygPkRu7D6mODMbr3R+b4vPlVHxehD1bkStNvkvrk5y4/hfw+rqMfI9XwVcP
SSp2CkJwKsWW4sC6jP8oXFHzVa8sYzwxt44vomUY092PBbZuIojyvzyupBm4rkIgfMvFUrGjsJfz
PHtNK4+qbmnliq/Jfq7N9IXYfDUezUy3jIYaAuBE9isgPXIxZBmJQSCMAvVt6w/Hd37rGRM42PwD
4lbSPDyLHEIUvgat8kpfL+l+x43ZEN3Lgkc+H1v388NyFdKL8DimDBLteNqpAQeGjnnVNfvQOHWA
HIrm5bc89WGym+pcQb8KURMh2AZ2zAKrVpxkD5+b0V0VhFiioj0lM9hDW17t//t5BcskRzK87Zeq
yynsGF3WAjbMsObEgNIxxxahN79McvuS0TsJ7OPJF4W0QDHvQl9xoHvR0sWdDwQwCTDhl5qRckcQ
0OW379Cq7NE9kGdk43nlaQw7T2aE+M+2Bn6kGrqnok2wz3wKjh+StBSF2woL3WCazOedrCseoCoY
RKdoeus4ZPpbrmvHCCjfSeMpYhLtRk4pncH2Np3YshH+JHQOCR6P47HKqqicWLi4zLSvZH0UQQK9
cSbaltXTjY/6LKdtt2Ua9HI4wcdTkuE2WbqMBFhKBflNOLLn6qemA65EHnqfcbOoaTVjS79qKGg1
QAFYGuYyZNXK/oZy0FtjceSyTsrC/1qqOM22KX0u/6P3QZs9PgGadVfSqTifUv3jFV8NDKYE9ZPN
gJIs6KomQlMothQmsuap0kzsBJaXufJHS2TqfwfLncP7niUEA8HrQx+BexjA+/V04hM2hLsUeAXP
iY0tQTq3FQoP/dBEc7fnGlQJIklVtPNS606JlAPECCEcpBrnIPKDXCp3C65H0ISwFr3xiWL51YtB
l9GQ6wsiD5gqPx9WsFe6V+wCcxUM/oGq+ygEu6yeqJ9u6kPKwQxQU0+A3jmviOHOswPzqQrTnG8d
WOZyxacmDeHNrF9+wAU1GvnHSYug5UYC7WZAAKzvUXTlwF3RZ4jzdF+7TtkA2aNwYwoRkammBLxh
ZRrFre1ih40pDW5hKyeR+GkvvSsxUCjfFA5LMCB6bvuh0s9O9V9jUJzVPsKh1nc7kzOzyJtNxVKe
tWckiqwLAqym61aoY9iGBBSd9FxwGA6ggPWvswggrGVkOAcHAQkJipwahnUM5N9Dlu5qUGtPg+3K
uktYg94nrPSymWY5KBim6GSflRpdI3MYmX5MatfhTW0JTeMcylH+3VnS9waraGKGMUUhvWI9ZEFl
TCNQcTnGl4iCVAmdlCON6ZJggaqEfzYszNX2WvgzinMWvWCAaXtYn/8Vd/S2gorY+dh8x8J9i4HD
yOP9WjeyLCRc+qbVjYKNOT9zX0pZ7eHJwcXgwPxBiMR28T2uq/wDgCcaV0RL7lTBrl0UFDcLh4Ed
QI+5uOj7SvgT0iflp8VHbrNfcgE7SfLjVNzg087moHpaLo6MDuETfoduG5SUn9OtMflUCiZ04NUz
hDnatHLJ8RpsmjVFIq3OYSs5SYoSaKufxAFw/OjaPG7LQ21h0AOoPrXQpbd5/gXceTRRCY8oLIZS
WYcxxxSJNDBTSPTrriBwl0LGJ3+R0TWmKzksb4XmIAg63Sg5BcB7EwSvoSyDLr2wKS3ZY7Wap8Ry
0LZzZkrqj1Nj36tWnuCyQGQOLcdsYTG84PrXYlilLb8TCklqQkhN3vLMezuDIQIS6/ST0bF6TDFk
tVoAGhDIhgLxYwaP7ORMu6gj4Y+5jgWtMio+988l0Ec1NoPcMj1zU3la4qvJe5+FI/e05go7/NHI
v8B4OXypG7LmHymeMeXEr4ZvL5I3I2QUGfYYEXO9C/Aq1mWIqWK5dY2/R87qGBmH70Qec7TGaisN
BMJp+JSszLyEsx17AmX2djgUQU3dSTm008XJlq+tiuY/j26ev8E1UykEhMqliktAam2zvZVXdl25
uA9qTJgZvE0PxTvoaRWBaes9VawiAzauWSP9x4ORE2CckbD4WTmSLKgHEizvLFoajrJcYZpMK0u3
pGiCPKsZaiqMGwD3jjk0Pfd4yS5aPBXzhc/bKJhn2OK//ef0caz8Y28vWvfWXrg7baCKPxBawXEZ
wiJHM3BFYLYWo5UOcdf1/sCss9XyvKtFtSixTLM4dO3cx+qJ13sPVxP13EFw8bmlfu1D7sVbfuM+
GFLd7SNspvPKwgZgrSPX8G266aRs9mbWeAFHgWkzeP7ZXes4YnHjuYQR3Y8ujY8QlcJ7dJxIknUS
wbJhfq4mU83FoMXZz7ShDvpetrCojPLSZzyW75OD6ai8uSsqcVsiu1GO7eIdILrDw7WoL5F+VCAp
U7QIgkHqFwkXgHX+xH2qtHECoBvIvRH2OXbF3HzL5vomQgFG6YhtEL9IT/Dd8b2d1Rle6L4QC/rb
MiT+K4snWS/Tc+nM1/zn/cDWxzFCitRygybkOVJstizaQ7AHtl7bgm60sJdOlQHkvivZWmFCFSAV
ZJQtndSDJY/vKnDT1zTcjeereh2pCXBfH6RTRPdO4weK/IvHCTqg94oUhC8OmW0ISprTy407Mb+e
gg0f8Tsu3v5bu1Vr/1vNbeG0MS2boE6A/i4Ik4PpPQ8uzc1NVCs2IVNEywzlZdrsaMUIoUuS8cLw
TJ6GUJLUtNpLlW6mbhwOSNcDk5Fwq95cmG3NFZSGd2NW/4x7/oGH/3Frafm0RZZ0hYVujpLP+omR
XCDSG8HA2JiwOpukMGXgkiT2zOo6FgWJsc6ni2Dl0V6x7l5DT0IIyohQ3/I3YWjamfGgF8nJOCtf
NWfu2dV/fN+84ut5c59kmz9RrKDgUbpO0+QkoRnhcg0QewBamtEot3GpDpEniiNsw4KOpnpc/u7t
9JRHjnM4sMx1G1kJufHn80JFJiye3k5Rg31zBtxCgA71Bt9A5m36vc/VlPYjPufOL0KpbJ3/JxEd
fUIbu+fXjrnsglXF6Eb/h5Y19Hhng3Nhy9Fgi9Enmhj/bV+ZNo0lcapnES/UFDnbjutVanz36p4J
qYR9TqLvltLzClOCFtmlJEAfJgOOnAzg442R1vPerz+ifnGGRb++Mv3uYrv3P24wVCpxWe/Nic5L
yrDue+29UPLz3EK4m6+ZDFv3ttvDkThtksx12dL3Vl0fVFeENUbYSxXFChB9z3YzAabcC+Brb8Cc
1OWAi+lKojWc98JWjDY5lD5yw/w2x43Q1s5ILLkeUdHMxyu8rMo6SfYpNvMfg2dOl7ZGYb+2fc3j
cUrmEWrR5lK89iqeaybmG7LEvsSKKPiRHv9RgEhtfh5nZFpmX0T0LmKP+NK7nGNuNngaTOeh7Ym7
nl8Jni6c6yJ/4MwcRv9cgb7BhzVciwzuHvmqZB1J9SiVR+Kkgebqf25YH/Q0yc8kDCdFylrQP+WV
s0emliAGochkjlFn8h98BsnNbiKWMr+2JoFg2u0qshzoUy22y4O0qtafOB6q9RLjI1wrq1AmzjuS
xIlvNXurqJWeHTW5RZTupApazlE120ou6o3B2W86oUoX4rgFDb8CMn4CgJQ4oaoWHrYm9lrY7RYI
z+cBdylOSqr873YjvOWfhduoHukHj/AmZb8DiYn/lpkc7FHKSmSFcV9kBvWdFl39AqQTrHFy6QVu
zI6SytlsQgT0gTBAOsInyuXPhzYJ5qc139w809pxIXiWdA5ZyxI6EEON37QBxoOlOEfZD5gBAKtN
YoLDQxxSAfa+C22dHHvkBJkmV25mN47E5NHd4p71Lq/c9iwGwh8HscaJBz3Fw4Ve+W2oWrKehe6C
WoDF33sP55r+8obx+cqXs3ryc1m/yclXXcU826YSuCrOcVT7w/fqzWi0sXxhE56yZ5UEdsk31Cl5
soO+hX5jh3zapFcwyf3lWq3meQwS5xryROkrfc3/8jhWXx9wWt9RKBieU7VDU+7UXS2sydLF9NAr
+lQTndzPbpviH6b5JqIUWHAPJYACyOKtlsCZt8LUB/q/FIOWZ/ZV511/Ia8O6yug3Zibjm2y5cOE
lrQ9klr9QfyORK70N33kyEeWZG5jcM6fO91buoo2gfSmDo8UXvnxdi5z2P9qTeKZx0yf9jOrnDjj
wqCx04Hdf5iMHPTKS2v1mm4miafEYaFik3ETdbaut+RVMes5vjheB7xAIRR5ADdgOwKwObEguHOo
L8RAKIw9WHO/tU65qAU58rJpqKOzSqMEoz2Ar/sDt97CqnDn1Y4VOX9o53QOvop7UbMCgWwDaXr7
ilthqQtujUpctI9f4CiWmBWa565LmGxIl8u2QZ43ZRE6naY4zeO6JHbI6BY1a4CqTORLbUvvAPBU
pkYnt8QKLENHjbAShKR07KQc3ZGlgfFTh5LZSiPxs3JdumqdEYM1sL/id4+loQQwbbI2JRm/V1fd
+8Y3xpTZQiUYRDycUMx9D8KRP3FNZq5Xg1L5h9uda5Jnleo5CVJBnwzK+d50a4C26TjqssGi+JH1
4qOvCEOwi/FtZ3KkPR35p49rBllPVomEqb03D6sZAo2+1CO/OzKmYcEzxZz/W+LID2/KvnY83BbY
B7ezS26dfyj4OYLG9u609eqEaZOw3hYhYdMPsnSg9cRix3zz/u/cYF7DqNSY8qUBFKVU3ZLnpMYr
DW+p0qJ9X7CTa0kG8iwjRs007iVy3Fgqzb28EHISYd0vcZL5N1N+I78dpb4Ymqc9/K+bUoER5BL/
48oCVbYoxz1R39MHMSA0ZwsUMGbz6iLldm21kE7zl967yBJPenLJiuRj20by1IdArNPZALpXpIFT
VB2l7rvW8CJME84K5Xi1Pa3Cq2b9aN81axI5Nb+++e4ghyOjOEtfc7UU8B+BXiDjIzlvE9EyKaSS
ivMWvJLEdhS5YFZNa2n1vciAht0EI0xpqomkzTVy18l0DkSmRHLWC7CJlGJ+dVgSXZV3f9Z0l5Zv
nIfmpXJM4Ea5Vy+XcOHdHfotiY0oV/Xv/lz8PL/rNr/jbA2r39Kwkcmc12T/feDOF/ywBC2Etq2+
2HK+b0xQNo9BgkvR2vMi/Zu/WS+E7Wj4vAKnTNwMgnIKT84dJ+QPK0mB4fZ5elavxkUQSYhH8LJE
/DJAOftTbEgr3WHXqgSh+nw26cTkIK8pankpJXMzJo2aui8f2v1JCsGgYS1FsDWqy/9/ax9Kg5xd
k7GaZQcQVcV5t3RnvElntF0HI4pZQWZ7L9fq96NA30VOrY43HNqoUXA0MCoyoxkM519iInkEyPK1
hQ8/4V5LTKda0Pd3leEaT0MQKOZwQxAcsWNQNuSZXJsI95tX74booe4rSDiZZ+sHtH070le1JVkQ
LTyKmJT30t3+AjtYti2qXyKwQJPNT7P1ijVDK3j3Huk7hUcMRlJmy14bPvmydin0iCEcYHeKMleo
gkNRkBRkKr2JU3jRAR/6Ta62CAjdKjNJ70rAoG+Y9Xj3RX5atsiUXbZmoAvQHQa6UBa2VxnYrR2H
9lZqqA1QHNHiSwxAMm/4/BcjHwtLDzQRqWbi9/3UAiFGRCZE1TD18OMeyDNKg0tsioZRPfGHWuX2
r1QfSkydqttE3fxwJtS6DdG3JIgGex3FmxqdyiPR++5ebF0TPFXAJXhDD2OzP2nkwZOw/H9Dtpsw
cy9zYpwojoKL6Ob3tPFU2Q734OJdnM6SS734US/6ztm140zRa0EIWd0Pukq+K6o1yKHvXludWBKJ
Iu/jsFW6D3Mm+bkFsHi4SpQCiIHbXKUGPsqKaU7yueBLVBCc59jcMQFEg5XWkLxTtJt0Py5kPKRP
i0EuAn3FoIsATZegvEqOqEJTRCZw9ncr7FcSB91VWWrVbwPT34hC/dOsgmZ6PlcpRHrhRyx6mP61
jzC6EnALL7GntomQyx4ODx8b2E35CaCkr/boHA3Hg2xwbPVvsoTeEA30T1AB/CvRmudhblwqDZdc
DoYvrJzmUbT4CX5Jxq+rct7ccMucG6h3XZOPaGMEweUpoHqMCBiHKpmy/CTYhe1p0i7CdGKKFvKv
IlAvXb9yUAIY+eygNFbIYF4zlfMHGiRFwmBv0GUE/Cc1PCxS5CtJL9HMPGiQ2TRo/unOCB19TSOG
BYLA07ka9hkXxB0oCDK1g1w+2WxDxHAZnS4X0CKrVmlyUR49dTgLPZbqnhezXhwi5JBE0qqETECO
xYj1laqkB4/mwT7+Uq+kd60c8fNc+XgVo0p5EGifBJvhT5cAgYSzPoTi+r+k4gOWaZBtrNs/Tj6z
WTiKHBQbwYA5wUn5aina/nPDSVoqNeLRScirfkHj2syxmic5ErKxgGj8EUsVSrcxfsbDm3LHkYOW
ImK3ouNaLfG0Nv4+UKfWuwhaFMqNBIW+dY42gWN3xTXGGx5iLbOmMdNCJf+ecj3dIDYpvBgmo/8J
AFT+aZ++ubznL64JSl5oLgRjgMUvlIbEfBPTTb/T3NRLA+RNRgDF1hjmdy0k6UjK4eXON7+Q/Pb3
P1INsgOEqy7onJlG+VGCcdqdgMdm8g7bEqhy8G2tgcYC1hQOaxLg0E/jHNbzrryDaXcYAVAkjYuV
Cy19VHMkSm1UF+opuCN3ioxcBBbvOOcSIa+YppqG1NKPQ3tsDUUSPBLeRn3VWeQcUuirJOC2HsCd
Fwo342GZlfdGQ0OYvzzkUdw/3QrIGPglAWzmPby7BVokobBCZ2HzodDuImVVG844J7p6glZWX9WQ
uIhHEhqFcNDslANW3GLezQZUUMv2MspJSE114MEY1u8XVPt9TYIkPpORv3UV525frMNC5HtYr6EV
8Odc5pDaritlzCXHtQqgDPptTmWUt4L9eVMDWsuRVVRQsM8E9jfzYsPN4WDPNnTVqBM1dSubRXMy
Foh2ygO2uIGhKsLus2XSzFvUjmCUOqJC0hZHHR8x/aDNjysbMEOjdGgRXJGdqjXgfpzGo0zT4m6Z
pK6+tRRICOQu8vQMlWVsZCR1uF3bpyHT8d+dvnzW6Dn1bZ6PRoYetb4ueckiHXk54AtzwlTeYlh2
N5QkjkyFQfSXfeOlEf8yFWYNrskDM9o8DX4GCdkBYydWTW81LW3RRekQeDYZIx5eK+T/PIRxgkKx
0pdt9Zzl6hPbn7XXqbvhi4Q8vDMCQLKawETWi+RajmknKHR1YbmItmX6o8kZXqISq9Eo8nMvqvCn
3utcvnpIacuLDeMNPkZ0fgu07wZQITUN6ziFfMsVb/38RmTEvfv9Gceno5IqAsog+9AErUDzP/RH
77IC8yjpRULXkP9l7gs/0Zbw7mci1vpTXve59ysEPvtIDRXldjWdyDlSjHxr8hwEo7/Mz9I28/AV
UT0lPga5r7k61GFd9EcJn/Xfqzn4C7mL7TNJ9y46+mt3219lIoE25ETQf23SAQW33BCZXxSR9wae
S9lm2471OPnsVWB0rsklUNMCld0mneFfJWORlGIQeTNgd42vaMLVLzHC+nirA9RN9twc0FBLSKxI
JFQiQIotzi/Afygy73OHFSHpwawglnYQ3BB0MX1jeUgfgk+t55WSg05GbYbHA8zDCHpz51Gyh6NT
jxB8e7H/ig6jbCFWR5YWFHQtcER4UKj6eL1DZ6ag4QGkmg+Vp0SpCkQ01nct9n9GrM1ZCX7RQp8B
aqzuQEwDbqrqrOwMnzE5VylzUANIMGeus/3/6ZD95XtIpliNM2GnugEZN066h3RiTjeV/0MUCLWv
QbSG1PCzFH+c86m0E3sdg8zjkLFEnGvdufenykBZU84yaMs+8zrc3xS5VzZCbZPtSth3nTuP7rBp
rLmaw4MuNaUbXzKoN3CHmRjNb5WNIkAgg1hCnU9uB4/bfuIV2ZXrQOB33OaNQmQiAWt80ssyVpDR
Yl5C7NqWLQ2C2y0/QW7JwZh43ATzFx/isF8+/i3gXjITWCIxNPTcst+KuONJK1aUmBiHs2rIG1v9
/QjhZ22OwBidbtl8x5HHZjhTivXQmeD5BQrVi/e3cMHPMu3+zGDkQY5jdHv5lB+poF1qZu1B55hS
/zusQXf3p51cRoAT/k53cFvKVdJC0LI0TzfEV3O3kX1QguBy+on9rbdhyxsqwAosVrli184rO+ZB
4TnVX+Gb0mG2TeTdMMfeWGvrOo/K51sALIx4dGCdN+mE+kMlQodhz609zUkoYwURx0tCP7CIHLCm
YsUjCarwevElxkxkIAOaRQ2KcsYrkFCSEstckSB8PVxcRtQdQW2PKrm0vyACLHUHspmoNsNLdSPn
hIA1wR2QHDfhJlp4UYWqAqbp91NL7scLiak/8JAlioGYtDNPnV3Jh3ye8c+ImqS/CKPujHe5Jih3
1GIfKo4IL2WuXC6sdQVhzvNND2AvKXwbX9ZngvtLwucAltYyI11T9BJH1HBB0IvdupntnxaWt4Fo
7Bq4YvkYfsLvXd68vaybptYxtx+VB1IPMrvAO+mvdKRhZtEXodPi2dk8BerVFTbwrcOSJXsVA8cV
vABKNCcTYXPAxli7K4zkP5COYH2lgxgmKOIvXKBKgiiksPT/V+8/EpCjkKMBRjc6P3DmK4zCUiBc
bwbKMW96e771E+kB5FjLIOio7AV/wuEPMy7mBOyaEyN/a8P6e4lv6AiEpN+dI+plfY7qokpUVDCx
bT3JFNy4HEAkk8mjWwf4sZNRAnDv36h6SHY0Kr9VixNbaZ+9cK3+F0GecjsGgImWjmbYdnnf9ezs
+DIhEVZW3i4AOCmnPkE/xZUqQLA3JwSHrvZ25dHBzZ8T+g72Bg+zFJ/hD6m2DD5w63/BPsWs4/um
9xLDTQUXxQMqNc73fpXmdI0Caa5b9TD69XRqRayhzhotAqHSHfL35anI/Ti4sa70f8/rIbm66k2m
Q+vvrummwl/SpJMci72bKI3hMgPZTWkIBJvTKY5r27AM2quEG3u8hckUnarkC+39yS1q+V7HA17D
/AAlopdqMS9lU4yeUXqdjmUZa6h3/J++JQt8iIXEJfIwpqvU0DrwmNvHvDQy8642zdeF4qAbFrLv
8mLoYCJghnPtGnjACr8PKqjA0GBsNKpwkgatqs40Y1wfceSzN3bU4uK+vuHVWNzLOAAP/v3rRtc3
ghDtIswhBjIgCWLKT0esVrmNbD3Ay84rI/YjRyXcDLcggoLszlXQlwa0G76DZ0DuFmueG3RzsKmB
nflSOsiyDXQPavb7ubOAsX2ze6b+CGaEuU2tiDLSJCbARXonW4ZkRu1jGzaNC1vyKIWNzrG7cT88
2/3h9Ae7kBlmo4CsKLq61zaMGWvgi5GkaxIj7hUN+3bLvBxPVJiQBX6KrJlgrUdbIwwm/Bu57heI
1gDR5kjw8Z7llcegCG/jihmVsE310QynHrfqqJ4leFPi57PImt2M7M35/9VJ1LZMfoGuWPm1uqoG
dt58HAIA9UzMCexPDQPfLluAUAPPHPDcuIuw2+TUaDBpsloNbir8dFOu+jBxD2LsUAMBvayv4CXb
GaeeNNs4Op7n8VVOuYxKLW5B4753+7CUvo0SBbvaAN0WRL31d/t/w4RdBy1gElNnNevxO9GpOGhA
hasbzD9YGrVurjxeoWkKX9zqJJkcUAyevm+o0ia7SHOgGXPZjH15txV3iBNSfELlaKWB5kkB82Yr
5mPDs2Ah5/yzCU5DhW9l4zNywn7kOhf+PF3JVEqkPJwAly8SQkNYneGnX1+1s393OiqgthxJ9byE
/G8clWW11SuzwYnwNOeKl8umKOtNRUF3QB9AMCnViWJ6Fj7BfWyNGDxMkr7XyGi1I6PheKvZB1m6
foHMGY+cKc98Db15jiiLH4n2CKcN0U+FYbAcGAGB33EXOM1H+ztXmC+PFWx/s6hAh0Ym0yHdKmnZ
gHpPhLKz7cMTeF7ISUFPcvud01CBBR02m3AYNhdh23AWngvG1Sit0V/EtNQ09Vg1kNe7Y5CTmxo+
iDnNO0/cGeDtZIMw2/7sb+m8rWA24TX88xESBd2MzoRdE5wWlAUCrxJw/28hlbf1czsOMRFNxT+N
NwjPiPyCiXeLfLuKzbj6rxZW4VplidQtslRI2NRJjGlF/xmIw75TXlX9FPisS0tgP0zYg9DR2TZQ
kXaGSUYu2Hb44ssnvCa1KDYUYJco8bI2CaRjkVho1sTXg3Nohn32uR3Da6Nm99R52D+6Wt918WxS
wsjVeVSVewz8cJfDO9Z075CTE7VlHT54zbSAWu1xcwZthFCT+jo8+20LKcUS112D18ar99xDEnn9
TMV7ZpZKuAuwFbwKghWpcp1Kr17+GoQMK1JUt2CWBt0Zg8GdbAILfToYPyHA1kMD1xlq9isYz74Q
F1amZR9jbAwC2Py/jbfAjYjaEumZK51fuDFQMdVUuBtYatwGYfIDj3Jsxx0yR3MorSV+26bb92tG
NWR55iSM1KuvI6pnHjdPVRK6QMeiWJQGavM/eFi1v1ZZ8OjLLDLr+BmMktcaAMI3lKbB7iyLnfwE
iRWT2YwEX849zxX+V/zy/QLLSaGXoF0O5QuumD88qXeeEL0iMi0UoMJ1PqLx83Ton76iIFBMvjOM
WjlCNJ3Jk51ncWIK0aVSaCCIl4DvwrdM1cwrT5J44/Z+SYTsc80mNFYdiXC+3qi9F0RoWil3XEh8
kamMjLnpaCvj6Bg6R5eNVLDjAfu2a2Xwm41HXS0FweFORGM8DG40lb6uFjIMVCqbCwT+qT8ZfVNz
joyDd60GHezk3EY78JMbN8UOsaR0L9J8wggpARl4FR5LRXF78QUpIzBTZR0u6XsJ4CD+P1JKWAlB
2p8XsIgoebX8AP1RZ1aUXkZ60/eiSp+aGjhsdDUrwRDDP8TUi6EmvDURJhwLf05XlZd0ND9TxG86
B4uwfNd6e4vMBKQ/uWWo2iWtmBUuYCU8xQfvnGwsrSRNYSIn3crF23UP/OPq11Vjqu6BmHzHhog8
z5J5V9p/x6PSxpWYXNrEwN7r4kMMbrFDvihWKgbUE+xagxPPZ3MWFxZn1te28TRhwcsB+dV2kAHx
odisNO/rwOvTvnWQ5QQYT3X8tIpXyU5KwAqoblgnyXWSV4JcgHFu631BRk0s+Ye+TtZ1p8FaZfKV
a4kE8Mnj0ZoWlzsR87DH6yP6FUYYSmi5ZJLrbAZgAOex/y2TbW697Rr7hsktPjqr69oUQgQ3mprV
fLfyshpiDwIzjeUK8XC2uGR6BxMjaMue6BRLLQyEHN2CxXi0w7g5rapIe+9ZEhAyxUlpSpZlcOj+
6TNFrbe13mFHMDxtaJKKjHupdQqZMshNxpSwoBPDd4kpitEhSaZebjQivAlpWZi2eTSGfLYThHFc
B7ugVHqHIeNdt8XL6M6Vkx6BwL/zQ6uujG0ksx7qQfpwa2nitgawuUYhlzZ0FzlUM1V0r5h4VwdK
RT4I8rsfjb5Lx2+z9Vw9jYR3plrVZm6lw0ZfiwmD0v30JkGcQb0bMKb8PnZVcnPMoc8nmdGrCw63
SzNjdq4Aks16t2krsosBLVRtWnE6LJwy7o1k02+/VVlz/o9lu/EbX/W2TdlPt+dWmy+r7DDNDImA
HML0xdOGdey3Gx2HZ+INNOVFA+KrGP+UYqIQBEqe8n9PrqVk2/fPofklIDKoocmF4kGmYecbJndY
MsKr2yQaSgUdmZ0Vvha+yFEz9TecoZOusj26jQ3XN8Gk0GAalJwlIZlmClR2Apb2g9s/UYZOdcSL
+7GIju2EwH3rkvmH1Ro1LaMxMswMcm+9oWnpbbQx/9SDlXuJYVjXdfQcimT1JaAeOaq4IyulSd+C
KjJEjUuOrfueS4V3sBniZTA+cFIrnzVBQ6LPTTy9fZkRMGQ3x6DcSExnn1sv08qHFyBn+CvRZG9i
3fUxoJm4ZQbJxZPC1i5MmZD8pYUgGu/NesL750NZESqiFh6HY+6EBD9NWVbHrKvQIFk0QKBl7wdS
JBGo70sXdCbzFOAV/R8Z9R8nmEbQjO9af8OClvr8K6eqeI9a+O++zOMPB3rUmdXErWckZDeXCEPK
9Ebqhuw8yVayk7MIDK/uX07WrkB+J1XSduUK9YKgSh5kVwe/Fwr4733uv4DuKDnGhrBIeODHQug0
6irh/6KQPhVJhj3m2tciqGef8Lz9WsUMGDa8gbQ7rmQLcrdIPzpRFuXu4wv7ny3fYpeV6YlOTNas
Amb6+6yp2pPpdNrJtGSCPqmUXLdXpmG3X54EUbyDxj5mwQuR8BzLvBdFux2EEodZ52hUfeI53PA0
KllxnnRbewI6D9hGjMhec12hFPXJ3aH03V1H/X/JEbUuD345VC0+BTo1DlNjgJ5pCkzkL1vGECdH
Jg8J/Co8iae93+JY9jmYCWd0gzK8TRHg08CZTv5qk0QyHKQJJLcYsmg7T28HP3cNS0zdY5baSSnt
hlPkiYnsGwlrFQQDhZ8HOO3lRwKMSTWbaH/oozkCLNSB2dWrB1yrWwQkmuZUAmXFQ0LT3BTwgKPI
8/7exa3l+5WjhPzIbk4EGzYLwOF+mmc+XSyCRra4K+E8HA6IoUcON9lRHAdbreOHf3MDDP6J8bdY
jbhecK1e6xrfX6+NBw+GgOQUlP33bFiF8vt81Jd9hBz6KMl1tkGw14yT8XWSWafuweZZQWAPJb5T
ecsWWm92VGPwkAzJpOEEEs3BXlwMStIC4hU9VyMTPh/m8nm6PjouTqnbp5g1RJpspu/APtIlkbdM
9M0O4miimBclgXIqJb6WP3KZLKvzHr6DGQp2q5ySmtiQDsJNyEBxX6IdBPdmPRhvSkwzZ4rtnlgl
uqLys4/KAM7X3mZS9Yoy7OEuXYHpxsllxXNgqYzDJsWwINyt0dIjpkkkPRwIxPLnOZUaHnIeOK8R
H69WH68HCVw3JnJIMq9CY5Beh+fAHPLx2B9t4gnJfQcdGK/GbZGr1Gp2bOmzsFaPE+Tj50ETidPE
udzrP3vheV9W9T4x7OAfaz9sFTN9paZTa26qIIgRjpQXU+Gib6ZqJFLJ+VSa9pI3aK689O9rRTDZ
et3ko0xvR9WBOSCoZ1Ru1DVPW1N8Bi2Y62X3VeOaJ1DfH4lxO2dn3R3eaTFcWcRnvFmhG7ZOWE05
Hk6JQ1RUm/NQcnGYqMGN/T9CvjAL5gldbp1sugYkfWis7YG2Z4V35w3dDQ+mRs/yZ78i6m5Pxihn
kynkyYFVo0xKX2bUMbOTLTBbT3bvjSBkQPc691G/IxQxZ7cg+H7AyhS7FxYhx0R3cAPNU1NlLbfu
4czYVLKWzeoMDh454obmt5gNes2PZuv+lW5ujOMmRUDXwZHM3ZCMAWjXUYlKix4HL5J15OPnXhrq
5RBnzPGEWTLfopKi63Cva7r6zSI1blb3VTaaiV8dZIzCU54zAnUqUElLPSBOY7fjNdXZcYiGW6AL
JvCC17VgO92qGe796rFsE4hX5FUqPhsSwYoWYZnET394BLAllQilCD43w/xGE3DvnGbu1rwiodCE
1i1Ipzg/0UCxRGDtEAcH+OErToUPD2rXmD5XfIX8SeiFFbhg9Tz6K1HgN9RpgwOo77ZYTr4BqPsP
tV+Jll5LQ+VlZWqsQR5Dv46Z0P5tHIJeyQRzSA4s36ezMPMn/q92Vr+uZWdCKBUzwyP37wOmjY2d
0ogjWL4OllpdgEi1GKSWM4ZGMhJcg7P4gCNeypvd3PUzYowB/v3DAp89VefsAkHDr8aKI/G7p88e
cJnHKF2mYZMc0uNUOwSe0+NmPRD+7fJ4ZeBuZvlD3xNsI1RAkDI5RZfpZFZsVS7OldCbom08xh28
/kEwvh7rAzCXTVtnqbBtkBAm816tfaR8Jl/IfKtctpXjUjX3cXfQO2JaRueAVf7/Av9f3Lw7Yum+
rpTTCI4OJB/Nz293YufWzSf3dXLIn692sCHNhAlGo8Z0TEx8jjSGUGwvlth9ln+iyiw4vpxF+P3c
2I01LsO033jbMYi9J7YGo7VozVqpozwu+ocmgI3QDFzZYBKo50CBsTaH6Xe+eEAUywCVzr6/eI34
+nprKea4Tn4eCH0djNbrmnghILADExOj5HtXcJcPbe4mVu35QHXigmDdmblbFxcdWumb46rCz8bK
GK5RwVhSmFAvfsEkTveav46yOwomQGkCMUgYpIaci04rToM/Ek8GTjZhAI1oQ+LDo2dF+7xc6YfG
bNNdhPX6t95YxvHZP77P43uHY13k5M9AMHLUSWXi/lYU5ko7KpntnqlFmAGCWKa9Lx92kKnZQ5dK
21jLyiD9f2O6hJe+CO99PhP7IhmP7gmO40k04pxOF7ivgbCcEluYgnkCly23AfxayGbsCy4INwxf
e5jnsX0j7GgKwfjSYb/VaXth8gYjoWlixC4zX4W9EvGKuMpVKIF/f3o1PitTFPasr1fzQ0cr0VGP
UpxsTaa90nW/+xVu9y+jTdPNGuCq7c8qcM1R3dPMFgYz8Eekm75rsbKsMB/YQlpAtqoLnyDXFmuC
qClI8SRhRJplYVz3RizvX/XXIRglAS+wGX4mictDdteCe7YC0/PNEp58L6VCVL95U2ZlCgdS7WF+
PAG3FKUdbzQ8StrU/C3dhWAMf95VWlVCTSk/7qwn3r41B5DR6h88qH6Fk8yz5xt+5pzXaxuLL36y
CXCWN0KUD5RdW6jvMl47i/9bLZm6HMcXq1nfrkqONiQpJYAdvKAsQDf/g5eNVxqNHapmequXe1Pv
zL0lm+Ug569oo36klxW0XBCBVpVjX1byukZJSCL5PEz1qO8dJkaXNM+Z7mNUQx7Q2PvmJOIB4THN
VW8bbU2O3ntk7/Ab4GCnn9wgFQr7T/M3sNpBQSVqP/f6pFhcrnNvMn/Mi8Z4gPJzdjkLxc0kHnOc
mww2cKs9Sbj2sqEKEJ/zTP1RPDyGOhiqDl3aB/FtgUKAX1QBHswKDyVdv8RfsTgXxXvYYmENFjRm
sb9OsHq6mmFmy3CCSByPa30Xqeg/xf3lzHz6Ul9ovfphuk6VfFEkfdieMx4NR+/F7V5xApRVL03X
p0kQj4zTuKriD2Qt/Ut+Gr1dBa6AxlZ3js0lTATIhUXk5MfFifhsP6vazhWSGugIbjpqu8+3oN3r
/hFERgnPJfNPTx9DHUa/TvyuFG3qtxk2ncwQK0OQCZAogS4LFY/kSLGits1nDNlDnh0sBfMnDFRz
YNu2ImRyzVlrS/zBWAovOW91OAP5mxIbpeYM2wWMaJ5h62Xa0/PAJCGtofe0mwFqCwOIMmstfy6/
PDs99CDurr8lqvBOcDakDRi4IalEp8jc1xmRLxcaYt4OJe6MYOQmdqzHSF0UdwZGge+ws9OJ2jrU
muKPHzORqruHo6iBAMMp7AB2DpWoDPkbFPB3M9upIaPqHLXAyV1qIQ3hGa4MU1LrhnO4O9LnrnMW
L4R+5sAWWdaCHfS7HZkPIh15MPhgZzqDUlEwMlKsG5K4RI0zwgRtq31N3APyFY/8+dXHtppDKMdv
v3GTYYfHxkDh88kEOaEMNi3joBFBogn9ZzgPvSkJ2yYHeKJN6NZp+I8GSlPDfpFT96QkLN26uk4j
saGzfpd2Ex+bVeUBUi95WHEXQ+UGjOnnk9qTFYYftsRfMYvzpkvkEheq4e0NaBlZ1ZjIPwc3k4KH
kI/eff7A3uWbSnXSuJSM8ovRyNzmE0zZvyVbExB9L4E4Ao/YbJXgZCiW28WoxbuRRK5baJRLXulH
UhWq9jLDPewcGxL0dlLMx9Yay4CncLSo9dI+1jYdid92z9nSvT9tC1euRIfyat1ZiMylxvPjiJUo
zC9vP0S0efVfxqMMQlU2dczTwrdM1SFvaxeFqV5X9JwNHp+Q5nf9Qa1JsoKqcyhmU9M+FqlGfm3P
fL1iHNVIlBeJYBKuafRw/skHLHTUY/3HnnIQ2kyzU0NfEMFbim6jR+/y+kqv3Ek4hviaZ9LyZ6D9
GfPVfc2fbAWRZYeDu0jgoK1uhb7eT799pztYMhQXgZgDIBwmxy4c7eyQBk96XA/YfampkB7MECwR
D/cXOpr9Wo5865wEPIwM0YFm0TV2wZRtSB0FHYmKxvP+Jhfzv7YGspkGPZe09X7KDctr1zz/Yz8U
FXEGL6QDwiquy+ErkOj7M19E+RxYZYJOlw8KBHhYrWvuWuubtHeVFEbM563WTo4WMsMX/owh0z3E
FJYiYZuFm83bQZ3bePLvZfmgB8M/7pskjyuW94rL2v9/ibp/nOOmkaxKVKeJDqFFD+x4BSIIdjFo
pg5T/a1eP6Swp9o4BTfdUA+hVOLO4xDp6Zx6Ftwrv/NvrdQec/Rs+BUr0yXtGCWWW95qVbQ0GxKJ
hQ6i34AL6u9iamCXB8u0+fG1r7MsyJR2mGwmGlMMYK5/J9xLD3OPPqXbJBZbDxCwYTrVVaQ4B1OR
89n1FwBmeTe7frlLibBQPYx+wjeJUhrjpZTTXDnKFxZ07646vfg6d07+ytNKbH0oRQofrK0UpMmY
OydSV8u+YLYe0NOsiFdWVX8GvJ4FqQc3W3EOlzwYeuO2OWYYYUtAy65LN8FHXU5BOe2hfbM7j/kI
ysgp9Aa/EDF2dYBoZDkH2XqzxEBZr+ibhmcXzfMp23pPRP1DWA8HJSIqaXLu6n73MuAmQ2HCbWpR
D/KD36HtxjB41/31cfstsoeZzADt59O/ltmBk2unZMAJuwbKULUTSo6Nwqdy/rhAlmwDFoIkQrDb
8tPfjqoC6pV2PCyQ7vfcJPel3aBXc9lDWb55v41bWeBU76h3htXe4U21Z+GxGpabTa70YgqporlE
ZP3++k+gYfM6hrKyPysWp7igv0rkxVtz1gJuyviFLcfqlA8WbKsOPiqfSYizucBx0IpLqBClpg70
QnAMFTprdvsk70f1s0wHcF7Ndl+ZxIYclaHOlBMNGROYy60NAfxRiQ8Pgkm3JJnTAvavX9lQTyiR
GR+WTMjq+h2yJYl2N4p90W3aJwO91RSCb0MVOaGaIQxXtXf6SaSt6wGLABOcF5x6rZxwl3I5YfuE
F1eg0MVtWLISJCNCSRSNbIp4xC9JTDNVkqw/9IYHKl/PDP5jE7s6gbLTiV0ttvzZlid4rtBodWsH
We1ANtzCRMuqMdkeAC7Z/yc1N0efA701G9jekjNMBJS+18493EVqhdrOgR/JTAAbmTuZntoWM2vm
W3U57MRJf6MkJG8dsdp7aXvvHv6FfrgSchl4cQCsU1KeggkhsGXT4JjtYLFiiiWbG1Eo5//Xrv0C
jZAXI8MEBAd/Y8PLgtgm3N0D6SHnzSNE7UFZiGXlk51uZTf+L8vgOCupSecPOf5J3iJMdMbEUs5i
1oSkmCcGK655f1ruj9sFoI2/Bmxb8vW06Vui/NB7fn/pfvidktdQ454JBhIo2GYfENxzo9YnrViv
55SA6OfwC3CcG2XDD/2kQD/Jlx3C4RSvC/Wm3wPDl9KFzKwIqTx59gsbQV/2mCWlruEpdAkaqnqD
U/A2yOwO26RCXk23hOZBABxHAT7nUAixrCgv1T+1H9VczxVJF6nYAQAfTDSDvcddedGXbiOLBVtG
MloshR4OFlsfDMdga6GRPJj9a1vLToCctWcIR0NkyY+/4o2MuOkLWdB6pB5+0yPNtrubTfE+tKg7
Xytgfxu1ojAi7SIUEAqRUrZOPSkfuFp4ME3vewGk0hx7BkFcZux7sLgGn0ba+ReX1NFyo/nyGruH
dSqWmMWEbModk3kVSocGplHX0tl+ZxU53DNOTsibPdcsj/3bk5z58UTmhAQmdJtvxXNL8L29XPhv
hirGjnywyYkxFxfteMzdPTIc3cRzjyFO+RxKFUyaCWCglV0tdLo1O3sckkHX6gqk4FpwlKdKlDMg
hDdUIrdvSv4FWz77k4FJNoru8coh9FGMd0eNBxSR9PhA47r4x0Q2nysJKVGwtSeIx6etzgXNkR09
ck6TNFcpNMTj+FADAwHNhIfERyUGFxvnWSRmKYIcM7n8Gw4s9kEoIaWBDmsjFlViRKgBPfeWZ9Ej
UGF+ALRlMIVKL8h5iDDEnl89KnCWR/o2U8jIWTCd6k5IVXuVJ695Yonfc82wY5dxSyKrRmlJ39G2
wdY/nJcNw0mQwGdAZKq/Lf/AEjHHSAxXwc6Acu56F/eqpDbE1nyQqnnqZJZbk9LFMmjY85X0iOuM
FHs+bZFMmU/7QyVSYG1dvT/mx/WGp8D4X4Wcc10gR14juopetrYBQtV30OiNOYxXp9DTlK7WVz69
GQ/IuUX5SjoKFzSEs2yTinSa90zvamQRj9ks13f8A7bSP4/9t/T6wGrsFeux/FTGQvJIbVoSXzpJ
G02S7ihdqwe38tyG1eGG1gGjv9XlmsJ7YAU7PsxSzrOkcP1YNeQOv8g9y619wWQPN17z5qJ9prPM
TeDYCj/2al1lL7V+ZvpadtbL7B9JBMks5rNZElVCgnEtTiJF0S3GuoEzlqtJ6NXhthak9DvQT/F5
DDDcFyl8Cfqgl1GE916T7xc07JT9+ov/8TSYtlDrZ55firYFxmUmyV1ae3eFweWFXAl+gCGCx/5Q
M8gcv04klxDt8URvhrBDJNrvX9gKQh0zeclcN8OEdNVSA/pF38qJPSoJNRBRiP2N7wzJ/27unzog
VqW3Je77oW6b6ktt0UEV9aEo5FVY/RtuOStKhcZd/eBK6H/zDVO2wNcOwGdA88qf7lyH3rO/zow1
TwvsE3OUqkJcab1a44x7VvNaTOCEig87zzJywCdDYm3Ky7Gf0eFUocfaeIQR/XYNPOojUOQEXn18
bdYlQFam8RpzS5yg8dTGZ9plVgBsMbP0quuMCuEBwCnbLSNGXFEchk874NqQPDS1H+7P9CTkeOHo
JtLLQ1FHV2HVYn1PlG38T84cn8v/ISY8hJynYHzQnLLT1DfK5KIb4GZwaR66BZWPCMQOTXClJSwF
NOQR/5kIpj58ekLZe07rZTAZggS0G7lQNjb7l4wwkW6kz/BTeH9/5pPdzyehshQX010z8P5Lbt+1
vbmqp3rKqx+u+cAVPAqAvED5wSVMRL/0mX6owxV1P+QZ6kBgQyWlPJ7OysG/jC1DBwhErV/NkhN9
Am0FQxI2+DsINnRH4CGOG+TtHxSa/rahrRNd/bBINpv3G2gYyVlpmHQBYPTHzo7/fY44S3wh/yC8
Ho5y//PMsyd9cEtoeFdAOjat2e7+bUYvg7CvyNT7Kr2DSw9jTN9ydmwXdr6+V1uwHBNQ78bQKCMp
5Aok56VAD94+rS2iyNxGL0tArNEtl3xzZoTef0dtHc8IVex8VDMx+xUyBK6ZoMhrIZ+Ew9JgZvgP
bnYqOPd4CnenzwU+KCs3QfCZZM8sIgiy+lF8YnLzY9+ll/+VZ4zfu1NS6sFbMVTcGdAwpA5cY684
rCcybIpdanr4wtGQUuwdm/F1b+gF1pYdGzc+lFgx4hiisMy74I58NWourWcN8e6Hi8MLZpcnpCCX
hXlU5ftA7O8yMlLxGsWKwI1DHQhrou2Ch9OdUdlY/O/+mjhqaOg3TeQRgRBRR6z6VjqQ2ofslpDT
s3xzeZQP79K7i7/qiMiqitWC/YvzWrdZH2JOeB4xxWOSr5le5OAuoNXgt1BogNMKVE/AGK6xhPXq
qRbxx8QwSqxLB+nLtE1CqL1YgGN7QVGw5g25odtBU1u9AdYjieeuwK6pzsM6SRMZzjKtI1nrXEp0
cqhRsfIzafyVGf+6BlDCnluqfQl3B5rXGk4zouv5c+m5/vbvKBEEnDc4BiCARM5xH+33YYT7Zhpy
t25mM+w4EIgs8KNaaxPcxRGbDFAiV1bvw6rJ3PMwsVzIz5AFJcKX17tZ74FbTRsNQyLPZ2J68WyW
IKcNzJit3PlcVlAcDaDG0T4ltWV69Asc/SvI3OH8yi/U53iEtCl1X2yVHOQULQ6BsF6RdlI2uF8n
T7fk13LxaOpK8yPQGd4lXKHPDlsattQFWMayjTeD06Rsd14GI8rgTxObohC/uK4yY2nZW9jfhdZE
cRiCVwfDky1onq3laWe4wFxdfIBSRgUfPcAyHxshEHOCzHNgsQd+aFnJlgV7A/m48bTCxT3W8H93
N6PMz3kgTGtbO4uiOoBNpl7arVcpkDFJ4nsfFilayuIPfB0+6zP+JprmKVLNIsmh/qeH1Hfu3C6H
mRey23WYphKWn8ptOp1DwvABCgHCRfTxoiRdYQc7ylRpm9AyUnUEy93wVuqKYSBL80mBYCDTLLu3
u7eKSCniXFIOZ7dei5gWrwX0Sh0CEK+ipHjg8jtsO1m+U6hk+TeYRHEtykbLjUhhm9QxOqwisOkA
orLrz8z50if0yzB4df2whRwOz15ZG8CvT42N8V2gePKHCo6QTy3WhMd/B13GaKdxacDoLd0NjQbl
VB5EQ2R41hfHCKSQHiy/1WxV5THRi2gboyjVwJL2jesUqpNko4/vIn4Qo0m8FqPebaH8d8JKaU4M
4fYjAsGHr6XjpCOEWOj0i7H1fQ3iSQE2YP7O88zIqMKDWtNB/kr2YZAF0+P1aATcLZ5es7vOxP+k
AMKsBrxj0RgEmsXsQwUreOF8XAHCwgDrGr5j+kVWRJZbka3TmV7UFLt2erYMUiP9rVHh5Ut48IP5
/DTgYMr04AST9cODeYVOw1Ck/cO6WAFbzVaL4sC+RmUg6XY7n0XOUsePP5IOTnIZzGiQYc+8BwiS
ETZE7r3hY1D9KQ5NMPv8flDHWwqMRW3BEEuZjQMFOYo2DO11sT3CTEwbpR5Fs67NjSwBOSBnHJOJ
9p7Z2V4kU1cVpyVoXvruiDGAE5ADlVEJEMR73vP1y+biubtEp1a0tqVQEGNSbgB0gefXySWTCWIp
qZF3k+YGb8iSvI3Yx9DdJtnPdp1sdr2DVJhzOB2oEcmpnuulBap1NLYVc2nbSQMCwE1T/E92EpOp
oSjgLPg0eTec+8CImxKhD8JDp0Buj3HpDgjGpWqXDRbLoM90e9QWNJQzEJMTN5VxICmIcSFD6iJx
tjqUL7Y/eHB/pepLXR2OSU4iuT/Ihl2AN8pRGJmmGbJYXzvmtKWFXeXceHDp1Gr8kkXFzF+q/rDX
hVkiX1ruChzh3vziTlztTL/pQHzW0ToZh79IQl987NAEtOCeGQ3/6RUUvKX6U/TPbAk3axdYHTHF
KrKI6ktozON+VVqzFsKRF9ldgwciVRd4ZfCL6+IniE0y1envah3yNzzdMCOW+iBLzHvMpdQ+P/uA
A2iWVi+ftrvkfKrnNBFY7gP5kS/mg43NHStqXycW82rHCdDSyQpengtv5EjQiAMELo6sb0ns+/BG
2HbxsomdHkLORjpCbHvXZILfZuAa8rokwkx3JXoRnKdpf6mkS6I2OWDrfpAJ7u69vV/AMbBpWCpz
ZSfgQx1K9FdwNIrwKnl1HPh4gnDGePxI4yz7CZj7nbRjhTgQo/Kpj5bekOgtz/wi7Qyl1Tcuon8q
EdP6wc54lPEVwThyiRidfqSgIInRdmaIh3b/QYw0YCfO3s3VH/7qHI+nDiuzdBEjyuYvT6pVA3fV
CqqxG2feBsCmy4Hl2x525Z2khwvvyNCEcnyRRl9HJ1UNUgWILNqtPcodLph2zNx1nI41i9IQPSzG
xFbPr1BvXE9pN0yZTXHMlamwfCYBS614+0WnPbQSqVG3XMjRk5zymQDx6akfbt0IcbPigpV3NJdY
gUrknEfwfZOWoAxdHfQ3nT6rd3vZRLs82cs9oi6ESqM49zdRqwqWia9ypQAda/0v0b08SuGV97M7
Xq3DZY4zoqLUUiKErQr5Ubn+G/lGyITJE8X/I+6630Puoal3+TOzP0dtHvzM9+3q65a8XfBLw/ol
XpBHUY8UFhVu+vfJx+gNmpvGOtWkjB/mAD9qWSDBAL2+AvsEK8zIfU5cavGKpwW+xz8xHYKXsNaN
9teNuNHgWbTjtwjD4N1ZAa3Hr7AWAfruseVsHuF/aEQ4pIzSFUdeZcWHRTzkuaoB4dq+DF4VSdiC
7NDB8LEREicQccZwPYiyXWOqeoJEAqWqClUGdRrcX0v81pTEWiOajaOGAf+MldL12vou/3MmhOPD
FB1Uk2W6QQ5dyvistcNbbeddbwE3JEtnSSUAqTrbUwBd7revY/z+uWOnqhgN2Cmiy6L2RBiVdVff
Io8bPoIM1khJXaOth1gOuaF8OgSyZ4XvTg1LfmPgrAn2t4P2tJJRLjWdSFm0pq3MM5m8I5QxwcGk
yy4iz0K5JOMyScddgz08C1OMGJ4eIChqzpR9yk5AtqSdpuu6G/TZx7ZsCa0GbqF/BarKy60WndhR
qHzOQoRwk1gUfc/LkOIa9ilo8bBJHHVwAsMr7z68SrllPDk73bJUMwaRp+kdswUkksQNMjzUOJDY
2H5rRiKZOKSH/+rZ0mtwU6sOsp2B1TYV7ep8SLRTEgZP6+JDeBcOCLjSCj2c7uNITn15gKYCbVji
+jhQDegBexPT+fs4iLKY2ruJwhDvWrF4G3RqiB52DSxvIwen3yY30P9eEXWm7j2RX4jfWoczx3EI
Fo45FEmYsjq7l9ajD7FB2KTbEByJYB//fKMrg+xlOfJxaBG5kHOUmKA638d1Ts0uxkl1EZegw/qk
vX/nd/qdtgTg/wUB0t94B8egX+DQmYpZm2m5PDpRrFLEpBdyPPcvG2cZyCIFS0CJEComAfXzQ0hQ
EF9Yzjx3+J0yEpt/V6iR2b8b9VoqXIBK6o0KNhoMUfCSVsJN09HuK/4lf0UkIUove1maboit6Ej/
nUOVDRywIxigtwzylgipsDcoit4rhpByHo6AlwBGOL6qAlADRqf5nwHRzLa3wNctljGNYT752d18
PoxkT1A9pmu/SJnqE+Ch7RSO7nNQLU10N05IDUK5/e8PX61jFV+kjQVdEq5kG2SwnMXTn1HIlyOH
ERwYRW3yx5YWfIjTCB9H9wvBuUI/Um9nIOiKRjJGsueYdBxkV0a/gD+yqSzSqwVRMFjUBoo6Hp09
F1fX8HWNpa+0AZTm5Br1zcr1VzqU3rlFygH+xCemXEwgnSZXTcyPDkyu4TWTi1PS/QYYgo9uzQVT
15MXxYtTWjGb7/7D3DQI7Gq5kKsPAFW0BYlZ25NA8s9gwo/9lSnixJvQGc/TngJ17OlML/J0zLMR
DLEre+vvDF/KYpA925YiylcC0EurJ3bquQJ1o6QaHPYhiuhQqxwBI7O73Qa8Qh8C09ialL4mduvm
7UH5q71b7F+9xv7EF2j7SbQ1nR1Emu+gygOGNCY3I05gGs00tFfFPjcijhzbOASbcIyUPSMCnerr
DMSTHAkr+RS6ZvvpNJas7TRUDN1r0DwVQfEmRwtWAPUGZqqszijTTMRUEmt5y8brpxoKKk6wwYGH
kaE4ew1uj/BYAs2Sp+elS42MPQitgJZvydGUbRkKjPAQpPXoqxOYvdpofbE2t48tm4Tp4LXn7XF4
KIIqeKBd+WfKsjVSFOEsHtSLVuYPIpphzqvJZ/mDvMHkd+f/FmLHbrVySudU3JYXs3IMwTGoG7d3
brFsur/bSYGI6PnWq+KvLy5cQd/3+Iv7jMd5j6r9Lx1tFtFXZdRg+eyqKlnSjmzAP/J/0+qlspfr
cY4xL94d1v/vePHMvhd9IrtdQf+gE4aoisYYu/dx60JCyjVYwtWgvMlB8IFrqjhbZJhZuK1giDvq
f7FcPfNDkL0bMser0wyFfXqVmjD5t0Wh2Vbm6dHiFC0sDplBxTThgJxrBG/9KYJFp2cZUkwlwXmJ
tHb2sde1cSQuMJqY7s89VkIu8egXp9eRH0dfKe2oKLX7uP56VA1WabtJ0rRp2C2gBnWWrE8pqKfF
rSEd1yHrArtdSZ6yDGA+pa5bQg/x7C/LKdnLEbLPYh90bm3CxJdv99Wkm5/0vN9nk0fsjbgGydQZ
wjJ6YcBEWxar9epmXCvRdr8xgmJONWoftKBAB/iAHEjD9AhoYJtQK/4/6GZ4ppabY+VamwwI8cg8
HZITEnPr3t/K3h9DlNCGz3yvyQXdV/LTAlxM5JDvh897VVEo33MRjgW5gw5ALLzyW7akPDeKga1i
xe1xPf4TYqtxRW/c13tYszMdr/4MxjhK5M9GZwmPPSjuyAv8fik6GMWqwpXql4Hi6+HYz2Atx140
THtLixsTPShaCef8Pdk5yINCwD6cOoXGFDPPrmpJDukJ3bdEfeJildE+rWMxvL1Mys1kQ0FI9RGN
qmuWb/EhQAqtSsxUU/4dTWmHnQyYA7bu8bQNJNL5uKlNvlNnuDTs3bPD524DZR1F2y0SHTWfU3Zt
+rmzYE0Gd1VEvKZxUjJL2kqrC1FFNUV3vGeWMAOMPdzlSr6OWznYJKBv5PgkZz8EPUkRAxKrj8BS
8d6gR4omxsXjrBu/ojwKD5dgMGHaEeiGBA+souhAK3dUlAEL+8KiHa6VVySl7dstS2N5220wPy/Z
EOglGTmCXNOSUMCWCEo180wWklERmuWGJIcQuf3KnWiDLto7Nq9oEMqLwwTnnfXxlshYe6t5s6JG
Bxwh25ZIb+NTHvS3An0+5jnWS1XaXpAVFPbM7ke7a7eyss9hlufQklMVSiL+MKL4e0M5UGSOBV5O
Rw/AkfK88PKFeLXXkHmb6atesGfg9NLO8xnJJ6yaA+Id8iyc8QOqfR60823ZPhc57EK81e2TwFv4
8SegPhrfoQ+RJRFNu+8JPun3X0kNVSSsbDH9NMGJYoLzJCPlGPbzNhvYSndK19wyCiA2tzSvxALo
zOPKFya26qpGBjze0JNocipr44NBRuCqBMvCysDIfnsJobZXQXek7nHlLR0al5iUMgP04L9Q0k7P
lAaBpogAkTwp6ySE3T4z2mcDdQkHUACLfmcqPr3EZFa4NyhEQ+0oOvnPW/cdol4MvuF4WYFKv2Ku
z2GX4cKrpVOnwnBYTlVGVwkyw75NulmlO+xIT01b5IVcr9RPYstjr3wltt+S2E4IKWj1hOAzFPc2
oDHfvTSYye2Ng2yy3hwCS7NpcdkEA1Ck/AedwRuPgyAkICN1hHNaWeZ4hJId8KujpFmLwoYJAVl1
tUGnz+4mBovuygMqJUjuaFus5/wtMPFQSRLNayw9BUz+TNDbRLUkGwNKoLaUPGZwxGyCSXcsH4wt
31NRrZ93KrLkT8RiXXERjZYgbJXQmZkKLsl0PTcls9A/E4Wla6bmkq/+0JNQFJi8wvj/CyBwkR8u
i2zv9Pm05C1T/fJ/0jWTjM4U5sF8bOney9TSM/D6UIr5lJZWlQso1O5EpihtNeexk+QjZBBMvf0g
0iMflVrx4MbvNd7kOeh5S/6DcMUqhoOEo4vLuRJHqTGvb85oLY4c2dyfNIjRgwjd76LlbJSxMBaH
VzLmZGUW3Me2nEi1psQLmHXWlfhasuugt8HHbto9q7QPIxupBdABMXyZzsZKsqHEufdJVbI/jriR
SrVLhDZ1qeN23v6LXV9V+KSEg+zKv3E9vrwWWybTPFa3eNegeWWb+TgSAAG9d4X2AN36c+/x7iz8
305vrECaaJzgxZ1fqj45SBH8gsRuK2+seY2r2qMjYi4o7ON+ncVxPCcdvk87b3zVORfshzDpAXkj
m0ngBWhsfYReJW4TUJnxd3CgTJrI3a2nHqVjJA4vLmMDD94/HvLgkJ85HVUBxDXqXbgC0lLDmJvM
akd4xiItVZ4c8izrZ6EQJ3KWE1/Vmp9EtIn99/Yl4UWT/xPncs08dExCgz5WdtFTcOmNGiQ1XwGw
Rf5se8eDxngbXR5oQCGlGshIs5fxfEVp6vcJXMM0jyOMRpD7R/6gc3WtK1st1lciANvmlLa81NvB
rncLTop7GtIslAEQSgA6BqxWex5AV7SCjpmS8E9l95hWl5pxWmTZ3XkpKfBsAX7ZGenxnFlsE3TV
RKRXDEo3bJgO12Ibxlz5jS5Dt8Q0XIVyIAJB9DEN2BkUeWcqXq9cCnbO7GKCZOhCHIJzR4vt+T3X
+y2lYuXNA7kn/VSOjHzJOo+TcozjkE4wJ7iyxWI/clQyukbVlQt3CVyp7lQDMn8bDN1ZxEP8HKmf
I5TeH8ZrV5gHT225omWgWzRlowQgd5wMcxpbzckyQSXo5GIVkRvSjSrsCgmz6QKbBXkpzokI5OgL
yoMMDAg9gjWvF9AmJyCfwca/gXfSkbtYGVGdcZl699EbviGTSe116FAjETRPDyL1H4SHfpMBI84K
ljwwKzSgstOKr+FRZSreEdCskIIzUdRb9BhG0PZpyuGgL82gTgJCWYwGXQkLjsu0016xRa/bpmcZ
OIrYHKpR6fYzcEtVkT6dA7aWT2VUmsmtRKOMXTnlynGHFsgca4E63YXqnTXqfK+P8EwN4l+40+rN
IOz4fO7qWkdTnncBhGsKJd94IVNKSUdiI0FIsy0qKJozpimMvf2qkglTvVA0LE3m8rzNgH7pF/u/
z1HCtB/Iw+JlOfUSgXRXChPD7IMEBmSaVgaSuNtUopf1uFHhNWKUKFvUsdziP6eYupH4EjiPatAL
kH8Lm7FBcsWGCUuQ56lfG5RZ/foQfuSYzo3x0FE33Tz5bW2gMFLgF+OTzjVRA7T0d1a/iPHTykAM
V8MIsTtKe7n/31Qc030R7csuTmNvu4tm3XM2xK6bsmSI9Uu3Fb4BpVy7JRahaJHsasUO6eJAJ43f
y7UeC/S54HBZV2zT8hrk2X90oHFNNa78CagM4hbvdt78ifAIbZ3HtvT8XoWJT5Z/z+H36GCtdZ3A
uRSRG5VhbzeFOEPb3GA9PofKJoFudajqSXIPi/TxTIne9iViM4vSrZeyeas78DOPfvsoBLJULxLH
sHCOMOafmNLCX1B5Jh3/wdNraLH2s1djB/spkIwzxf1rJPSHMJP0Of0I9fxmm3jEBgnlFwVph3LB
f1AfjXqYapallq+FmOF6myeButW5GxpdFguXFbzZhRiH8Fk2H+WHkf8M3B6AX2y9fvf5h54261jm
7eC8rDHYlV467hjxLCw4ChmyrUgHPB7MQLsPkwKgUiSMvMhSBL64cRRy7HYeMn730CYDE1EfVR3l
i1bBFYoMJBCKuNF7QhgLFPDzYr7bJjufVZZkFrZ43Qg6TO7h3y6a2XpF6MqiYCdmivwKkxvGDJsm
i0Fjq68pL0N9Zlj8BtELeHVTok6355TyKXzFzbxq+YT+/o0tzdTf3bhmirss9elWUzNilh3LyfPL
xULeh6llytWPSzbrAk/Y85GAK6Xh2M4wvDm3tAFwCa7Fou0tvEqpvw+DiVRynlsC7SbsuVm1qHCt
zn4NkGGRUnk6K9RdJdEevYvoFaok34Qs34MO7hwIQv0SvCGK6cHq4ZmQFEln1EMP4mpb38x9yhp9
RumqVpv7urkOKGN3BALoUp6VxbZagDZxO6vV+74JUmSNL+WzrBV/G4MQr2ikn20c0PMkue2thI5t
cIeaIXa7v2Hjj+wOmq8DOi/sN8mFwMn/hoPUlm3yhYtOBoxWvbgfKlWudAWzoiUkdd3cgrAVgySe
AE6+JdE0/JIZIQLjpX7PSw9chkx4RqFxSY3xoK0GTw5TL8ScrgvSP1igs/6LFCKHIvIGQu1Rtjp4
fXDoMnzKaYeKUKVEgACmI7t1LDWqAgDGhYo6pIOYM3Xv6lAKDlqoJvyBclUz4QBxiAtejy1Z8Ubp
HZ8zWgH21noNMCyA6CIwvZvTwX570sAUpzjRNHTIe40/0iHm5Z0kqeODujusnNJaw6OrhKmlENwC
8ORS68H8GDK6oJS+nekFCnhiBSGhvM18On8FQJWc9ZYaUWBnrw2H/8z/RRJdrDHCJ+H1JU0OXWpq
K5ffM2RrHGXsJW7uUj6KFPtxzI2+W6uFitHUafbgHqlf/D9gb+0iN4RhqS3Hoebg84CqzF2Lv1xp
tvImkpZI1wk2SzgQGJJFsRJhyL7DPEN/9qkybv5T9NG6C2TK6f8sVlR3ky5XJfnGAbjPsM2e5I4B
WCXY+KWCIZGd8NSI1Kwar5vfr2dOaCpAmpECVohi5dxid2CxkpRb1lGVKroc2MNpI7qDn2DZo4ZO
3Oo11D5+j7bIpIUzm2YCSjnBlxVivR9iBUKA58Ul3jgHhBlLBe5yuOrTasCl3fTfodb9rLFQtATX
mz2gX+svRh4WSIOoHMbVBpDYYNXZ1/ziUM4ZMcgD3mbyHn5hIo/z4TX8H3yuB5ZoNnjN8uTj+aBV
iiF8EtE6DiHYCLnZiFXyVKzlm2oHhzZdNvBZGiUFqqlo/W20TF6B1zBV9Y4xrjJqNr/gCyJW9M8J
BgHMgAuOAtWGQz4RRJmuuOL4/IKGEowa8SPQMDIBqtsss3BVLvG5T+V74bDikFozoo5unQc/Q62W
hirzb40aCNH+tovnD3/cKfnuWRNw0oIRsAOQSJYSYycS7h4ZJvYr7NnsXgzp/BHl692Bg73n5nVg
e5OL5NLDntKDlx1ePijTiTqRk6HgIIUjh03IVno3rG98L0IfpSiEmNc1lyLTQSkhLX+EI2umKlVb
RxZK3gtOlC6R/tzsG0AkXnJzi4LdIOeJor8G0zafu0qSwJjTq7TjBjGwAXYIxtMytYsHnz4O/gY4
TpOOwQ+p1qgB8AYnULaexBR+OlnmOSXSM9quhj9udLzyFAA1b/KPBqGTpW5EasQ79oIMsG7EJa4y
rrq5wCZpKNkb3BW3OxczwNIbFMIObfK/0IdRVhVUP76IT5gWuQJW8Gh2+MVYnZQIKkOWhLBF+HkQ
O5qjdJkJDYQ808zNH1pMQXFuLQF8q5yxb2gpVCNAsTq9b8m8pRyqp8JnYAbs3v1sKLU+i7AAzGcq
1X/DB/fYbd4UxbbG6c8oDvGz5WKi+giw5M3Dhm5nBVRetaA6Hqyxk8qBbiKL5aIFlg1zCzBzuh9Z
RmGDTZB29qFJhRW865lWaUdNg87tpl+sTmc7j08Muz5erqSrmPtBq6E8tQHyksvnZ5A0GoqouHPZ
EHTdREYYI2dW9oM7W1lzwQHGf0QNb5chDlUbJTRRkpPf/Vy5xFEGL87ZKeIdUOLa8x8hJNky1HDW
o6W/wkLslLnWDutFK+OdRIYYBjscHeiYFVaUSHjmyhgFLLoBs57d3Tn8jK0KGn8cha44XM/55Pgu
Pb5KAs9Vt2GyvY/GOhqtwxRDJ3F8wRxu/Jo5o3EU9Tx4o7DzxcEjO/cLBIUjAYmrC8vLw/DLMK81
C+v6REWE8YsydC8wB5FU5GD0R27EcVzzG3v3/+N61GmopRCoJAsgD0UhUtoGeeUsklocOWqn+Nlq
f+1hZrduZpPanpJerMRiEmA6dTA3H3j6ztgiIXZXbZy+eybIExOBXSRDtdfZhXbEoIOua4VJz9J3
y/DJy1rJRmT2tCTtpJGtbfseso1AhyQCZTt0TbrB36DNY9Ba8f2rreLsApUT0WSNTINdk0yCKo86
con3V/paVa3UtRCRcHwPGhmpWnQ7EyrKWZR35m7gCmylAkDlJDmZah2VAl+v0pzGVpu3KR3tqviU
IsclwMuk5lbmdosoRqHODQo2IrKBixHiGf4AYaXgSKzK7CQW0Eo7X28ZHicICnc0gNGJpDEwLUxg
TGrT0CVinI5tvbRSVzOzZ9ppeZTWOxAAiRZVLJpIeCZYQ87cnoZqu7CzTP4Hi1NLHXHhavQZ2TAT
PFwSdzELwOJszC94jK3S3zc7uRczKDe2ZKBSGueefgUwddJlDRdefSGLdrsBO34cce1yjAIZjwDV
VnLmnhDN4UlfkQ6Kr8B1wjhM7BrelpHW8QtkBrEAW5Nqm7Rpp/AohSA+jTWjuS7shF+2X8iCgnVs
s8Um4p4wAHb06iMq/pzCrJ08CNk9yc7MTOis5I7kNN5+NkhQEOcZlAPh2LNn/8+9BGa4a9V308Uu
Fi1QQZ4z9iF72qijfQwwseUZODp81oM2AUmlbqL5Fzt9WsLwZ1cHWTj8eAMrtBe1g7YErAp9rNSg
z7fW00I0e8+xfTvq2R02y3HyLA0ZGUZNY6EAcFHMlfOi6RvCuY7nKxKZ7zeNsmy7FacsGcUiZmHb
n8dUPXfeq6Fx7fhSsIexfWPP6JjAsmt14SheErml15Pp1kLjNay9T4C4CgjFrG7hY4UH89iTyQpx
5iDe5LtCGcS54OeW9mRq1IFxga1WW4avWhuVriptf9LdMdAPnjMF9GKJUBwbQLi9p2WlGsnh04Ap
uEvP6cMGa8nEQ9CzODgQA2yJ7kj5EUbgRwJ1L6Zs7JyWwhwpdCE4V9ocH0Hd39gnZmvgpCrGF2El
kqK0r51gKtJGQ0EkUBEIfleqFlNtaRtKc1Rl4zqf0/zaYi5FxNwVXgLZpGzGtKRbQJy22RWFiyQ5
g5uXqfzuw36QjxOGtVmOq5mU1wtEmOXFUGzLfKwGZGf4NETjDhQtkzUEFliu6VGQl7VNYbQKxQC0
hhaa+v1O8xif3CVaW3/aTNslMG4SdY7SwwXe9Imoow2/Y59FXnF47oZQ5Kw4tsf5Y8j0gBqqKSDk
CF/Qu/iFxzcuuooIww3l9kYTei4mR3pft1Bq8ctRpDtHtLo2SrXsCgZWtzxJF0UY/jwkTNDmTuMH
ASPcTSxtXi05FHUNo+voev9/M6MFPp2U76hwLOmU5HlD5HeI5PjqW5HUzSjHjXTLy4vNuCM8BviX
XJllnOc8DASJa/ggb7+8qQquTm1htqT08PqHNJZ9AQGf0PTD3T/Ealr2xA3p8Tt6KE9w4v4OgXbN
JOGhnLUm6DVvM4omptteb9/z1NOUn/3yx4D3lQNPnik9RJsrEzNQdCdF+T8mTcHaPSc92hYPpCs4
Dv9bh42BbCvS9W0TUHBCiGCvodn1cld/bZ/IOxh0CQT+lFChCjn4dBgde9goJCypGPoDB3aCdnE/
l93SbpFrcU5qTnaxcmMoc2p+l4+xKjCOgcEYM7jACYV1FLwMx+b1I4ItpLJNiRS+9IcnJElukkTy
DsJEPjqJsUpn9WinjPxxVJDyOXrGni4w/cvjeAv9Ah7iRCdmP4jXUQatm/tNfo2vbe7mDA8ik7Zc
fSpwkrxSiWM4MZjdpssIUxbKT8XDt6P8fdWGR3q34LHvmwpsrixShFrPoqitXZPtfceHfJZW31D+
I+wIvHwQ3TjwdYkoUNBN517gvx28vI4mX8auyigDepMudbSUA4TROrpvYMh0gkJbjCZYeS2DPGkF
GG4pv5zccO3lJXQ69HNxQLz+O4axk8d6ad48aI/IpowsTI/efpsIBM7aSGuvGwhJWH6Xp+UWK7pF
wdWbu1R2zrD1S3blED9uvLEA1d1a8Cthutvx03cs/816VRS5x9hltVqUnOsxh4JEjPdYPnsQVMbR
iLvbkyHZ2/Dagm7ecLVGodjAGS4wOR0OIS9OVNlS0vHlyvZ4RCpViB0H7zPon/rrTd6vd0Y1nQuK
hrjn7Ltks+NbUfTnv4itZuRG51AIw9SDvvPmoN4cVdw6Mxev1SFABhJ9xYfDflkzy0gHpPddxrZd
eAhd0iVLesI1rAHZznpF9g3Y2AmyDFq5Aw1dfV7c4KDWimtiyNoiIFzzfQwNoE8oWmdXggha1cPR
VsZ14An0FFlznfKTtdXT5oCbkU6DuRIMXZ3BGd956azVvJOTMttRli7lD5+1Aog9aw/W3yjk714E
W42x7vq+7Ep+Sav8D/eBGqcY4smk/KxandFE3BmaQC6JAZhaRNxWOVQsKWbteHPVORSPh+UB+mm7
j3xBYq73lLCj9vvOeZE1cxv8oie4lIimgcD5C/RE2gBjJnxl0ZwJowK9QG/sxpsCNZkeQV+DYeKL
nFPNZpdLKqaeN9YQPqlsffEnTOTZcBE+DwB9KhHELecutwfnla27n1PdZ6bLkgY/v7/WfYYuwuS9
uDEJ6b91N9w/BxMXt17h2vpfTf/oAaNDpcqGjFzTj96n3DWasWJcRDruqVm92jiThwX4MvCIpSME
szPlPfFbEO+6QeXRGTuRcSzOYwzl0vVfMmYOmcdSrEnF6do5+MU12G2/fII45zEzNgpLCL0UXsEj
0uYYNow6KGd8viTgnXkuHutq6B3jqShfUUnQW3Pim6yNoZtdewfqYk1MalLamr4yn7hhgGJrueWh
M+/2JysgRObK0h4t90wT2ITpaozgQnEqW0IK3VeKJi6ZNq8TZZwDT674mLOn76mrfa4lIqa2q+fe
zSv+1Q6KgSaCYuOEvGZPkKgTZYTnP7SITektjD58GwhBBDBuEmloIGyonWCuxCb/JEJOcvoffjpZ
82CoMLpxGBLoFG/yfsY9CNkF55tywtUo/HrPtFXvftdzLznoci4ZBDx1MbFB5rk027xVxnESNG1p
GakrynwPueMP3DW/32AD8c37tvyjTtaAQckjEPk9N+TnjHPKJbrQnEnSHmi3PT0aYKEUnk15eBhg
MzxROhfcyQ+AbAiC91vlvBH5uvME6+1REwDd3OD4hsLqrIaB91houP/lXNuooLTSqiWi/xt2MQC7
MMkAF3CLbRAF39/rhkPH3qXeXKjfU0uEWmwerd6N8TZfi+FMHBi/hBDd6mbC08DGTdOnlua2I4Nm
dLot177EYuK5Ezag5KRJs5F9rjUbHihEMtXd36KhpZcR/jSwWfqJfwGh95YBQq6kTM9NFd05KlIW
BLrL9ZJK2qbywMHBkpztdDWrnulHdt4Kb82jAmSnpVIygx5UC1/Wsbjm18VVFtMDu0yUvCAZoBDq
A7amMM/xcZ1r5+001lf734Q4lW15gMtxdmj0RcefO5URtxyr4Ct/sU+dfJJOPrfvUZPPTmg064W6
ahFaZSbB7rm60aFzucFiBQO09tULv0mTym5PiPtqhtIgRdnsRY+tPgNhpWwtOmzK02wCp1690bU/
JMy4fIRZeJj5I+NJFwpIz3aWPtjZtH7Iif/RHqCgQWotI2vwO6AY21BaGLg3/sac2DjfR7uaC+/l
gKvFJZvnqepyfJI4K9Lg75IqMkj5lZ5NXxowlMYYSUMk63Wa6ssuvYE3Bd/Owuk3geOBisSJ+xu9
9zNZsPgoIfUJuOt9GDdpObjyucsG7foo0wDSsVJn6NeZmmHicpzg446pdYCV29Qq6Ab8wugd8/PZ
mKskDoUEqsT7jGyeClHGqIZFy1m5dOoO7UjoBuItKQ79AiQNkvlv5zkTZavCCi3ht+59nkjbOUeH
Xe5SrSCsHqTS9/XRAVeWqLtaTnDsrstNAznDM7lqTyK8vetiAoXqBBDCapXODTBJh/hldKY4NWcf
BWZHQmKcHeAFIpDwlPG03tDkLO3WFypAtQ6VbSZiwefhg2oaCEp6BU8ZmwYz9491w0I6dFIPomlI
1vsJn++Gd/7zao58NhnN490JOzlA8W/+Ks8hpAQBl//gE9NO5qgdYFW65JFLYfN2OnO73EubqVcv
fGHKZKfKZ9yI7+q3zNqf/IPsvjekT6RnlixUi8XcrIRll+VXW9g+0Zb98SDuKjZpMeuoExs3BzVt
feAKyGpHLypnr9HG20OoY5JtKfW+i7Lh8krFkSGuJm14CEU872y6LQnMLlErcqy8RyMrvVGanVGy
1h+OlHTCgNPgKXUzQB7dRrlbEl882ZqG6SEx0lP5dnQD2Dfayj52Db3PuQYKnDfsylt7FzVnpOZG
DffLnX83FpfHEuWeJNvMx4KNYM0XTe3mos/kzYzEs7wOScsSNKiUKakCueNZEwADK+3TsTmCMPFm
DADQpLVfhRc+rVZsJfN5c+KT+YVm5d5fhBK4x2/XRaxBYNVz7CktGqDEQiljx3qZ47eLueFgo9Ve
6oyWS6kzOkMu6+OSYW5cr9gUaaQn8ZzHuwB7+lqw8arBTABkr7Ga2BZwdjZYBze1sJsi2edj6T9C
UcsxdV1r19C8xRhoFQnOPvTpeLuSJaHsQwMNRhw05JMQ/5NJ7me3MSY9VlIVuJlHplCFu26SXOJU
eShlyc5IqmnkOoJv91+ddRR5ocsM7FqweVDCloj+mbbLl8sjbaqz36eiFIlh0ME+fp2jODA/zMVc
X/N4EYTKG6fPgeYHAR6I8EMdzgNsDn1RZUt8YWsaxUUR32BBLH3QZoGJHKIrkfxtJtkone0NbwOU
lX2dBLrSfmwDf8Bhetp8IvDDRGas5Htz7p0jMn6jcSJk9TKrKFMC3D0ImOl6YAb3whFZnuhMG5/6
y82s3mE2LarpARsZNuyeYiGehE+zREo9cNV7u7+u9c8Vo60wbg0I0BVygkxxlXpgxRoRgpZwjH31
KYDsTmReRHGE1jfKmbIUPHTP6tK9WkFinDcc3dINC2VedC/BV/hnusbuUg6Z5C7k6+41hIkrA9Xt
S0cCIpZWJak5u4SqoJhA4kkTHTkZqXp8NZMKe0s9J4sLTZqJf0A6wcmMW6X2B/YiyWFeejmKJHlL
q6XXVVj9VCaDK3oeKvJgyD8/xLusplgGt2N67gVhQxVVl1hzLxWYF6UblBjnzw+6o1AH7vPdBRkz
3kZ9VGIPQzD2SuhiDVbjiJs7p59Ai5aaG86Pd0C0aMBEOzsl/5G1stBpzFE5aiZ1jOJvmfGRC7B1
NHZJXiwAqrwqHvR+7W1VmS819bnkVEwpK0/Ihw/euClYy3L0uAMlqYpYWG15EalbSBwsWibFMQkD
tXQuaTtBzL/U9qnKjxEXF9XX0UriC3bQI1YA++R1jz+NgZhGETgRuk+1HngKi9nqq77BKVNyRWsE
zaG+MwXK79m+9e4xoFZT1yPPzHVWeyLJBSo+mtRiroDSw/j59x5AggrCjvzjYhyL4ucivHnZxHwd
crVBcp39ky0J8eaL8D/136D/3jPd9D8alnsLjz6ACQF4zLz/hRWj1+8z/ny7M/voUffSCmpLkbJj
4dqauPPiFRq4xBeQm89ihm5jOCCkptvU+U5KEg6vBluugIwiMc9BldWgXwGYh/Q46zXKVv4keAB7
JYQORWFtuixWYilqiWy8W98FSXAOToHej7qJAJBr4MeCMuNwBh9FDJrimFq66ZH/+qttfgCZI8ZU
tl4I2R30R5M8zVvWVqg70PtH8cfftentDqqrndWGQWKDfIfyTDeaBOGuvHZg+gqARIkI7rOGppuk
qTakZ0bi2l8B02yv166CrS6LFdaWYx3bzlaoDwno6J71PctLFpfyUdaE6ul2UB3QHl7u51A+eWe0
5LRfA/eeABB4NDyi1TPG6mNKsOBeksDgLFZSKGgwaI/cZ2/kZz/HJ09MW4wQhp5rOH1Cqqs2qwKD
omvm2zOV6S1/GPTr8zQUz8LYis2E4ZKzulTX0tGhIgWfRkOq6YDDSbW5RuQW9WCgaLPJRXmd59eh
vytXLJFYNeO09n9GkuhZy8ZPBDU1lM3ZtuRd/B5zNsA2Um2NsYFW9snUzyBQB6aWKTlh3body7CY
h1IIuEAd0L2wohReThO1GqMOUz4LsOCAgfJrby09RMQ7V8Gw3esi8RS2fyN5iO8dNckgOUXeHamn
enAG5HPRA0WLWvZnC7vBbi+Ck4X8hEvnIrUF23ehYkfGkI+uLuNGB66AIOMna2z8VEM5KKWQ/r0J
G4kmtvlna7thCz9AaKl7cTF4cFs5F1wv0VGcDQdrYiFgWx9C4IALWi+6wsMLkFpY/DEJe8Xy8s+o
VRyszxjhh8s8Au7Y/l6MKJzB43nMWfmssTH3GI662JDeC0I9wpAyYgTjXR2e4bEy1fL3QuiIOBRE
gvXpggDCH7RlCqLYjNnjR/N+gp02DsUjk57PsrE086vx5gVyWFCGVS3ts/VEphxhoqV2PaPbPEpt
Ww/XFN5QdlHwAwxAdK2BNzJTlImgyaMsaYfBbL4/UoHUfED5uT5Fh+DQ/UBR+FQURQ4eyFB3+tmK
Fgr4xixe2bwD+qwICc2UOkgrxgPPfaROllv0KgbeeywUJDBvHqDtab1tzxOEWo5Wp2J0hVhWCmkC
jkrLrPhEmcM1uKv600x9BIqvycOanSi6eMn87VfYrh1KWczybUnbKqYWxXmCFM+KRDSZj1XhY6D1
j0IovtEBhhtD4iwmsi6OKunsRciPMqwsZlwpsdutRwcRvYV1s8oikRQAPGf/67UHtQ35yTbiRPyl
UqNr00FEK0QWZljUE8TZQCRmHwS2GSJACcHbW67IDEhKLcCxtt2w5zvpJJg2ZsBQJcUhdUCsBp2I
X7NUOIBjeIxKn32x174chrfnhWKi+Cpmr9wqUPX4LtChVRnpMaFZCQojF93HfSfHcMFiPaTMWYJc
rNUyAO3nkdPu6xp+sij+WiSNhRmiwwXQb5IrH/PXoWzbTbCdKY58HZPegHESDlyGa+1ce1V1vWjR
v7THM9WwUbyjYo6+JemcJfTF0bgmB03sbw9jHK3MiG+Dhu9ol1afwum+szFf4CuYBaDK43XMVm99
40HYBpTMluGqCOJI/bypRx7nQOe+m4G2tQK6mFTP9rRz3FLcEFoE4PF0VKxoQnF5UPkVJEEgX5Dg
6wU/SDpaoGFKNHU8DJ7YiyKGMIHjIkioX3HQFmEFUjzcQi6HiYPVAAuCbV+FZfmjRAXc+bFxUpTV
UHO6KEYl9Qn3cjskWkaYlXGt8vuC3bojjJVku4Zo+bzLyNNVj7LwFpFcVp58ehEOs9tStXbd669/
SFOl6APrhCr5LBaqa2q/2YLjHpXiyXh11Ib7FhKPgHjFSZ8NdBb+QJzGs+WI0gIZHvMJpZ85V0BD
14DkPQtwfyhjrgmqAg0vaXpiZhgm3D32BKs19Wyl20Iw9C7D5B/GNh+Dq9zvXbKjgXHjJlyLiDYO
mJgg0TPAC7NRvuXHBZpaMW4qE4Cidp9DH52JoSr2GGO0ZSbSyAVp+tIajvD4KIhLeD1TvYnzxcv3
u+VxLCQ/uLLRbSTYKLjMKpcvSVsFoReDxrQSs6PPvx1zlRgWBQPEaLujM8G7IGBwPmmUrRlW2+lT
rD8Zr7ES6wcZsflM4DBvt//M9LriS27rq1PX5Px7tm1JGv0pkzQu5DisZ4ZK53xTvQaE4gPikDcx
prSdR3VJmhBGCfdqgrGnR1TwcZLAwl2GsH20MUodjBMUdL4PIzWKM4rnbxxqCYGK4Gmux+3VbG8U
RMbR+wg0fPvM3DrYp2eqYj4E40Wj4fW3vgjJjrU3hPFKg19o+NgNmOFRTAig8vBQjd5mdpzL0oRJ
KEO3ppE63mznBhkqgNRAQGA8TPL5B94Mzh1pVlMzEJu9NWATq3wilyABECWMKCuBPU2Dr6mvdBUc
6skgB+ufLwWEvZbeDHXAUNUzBjgd6aCr3G3sCTHajExA9X21sY/1zoBBe97rUPiRvsIKAAhaP7B+
Mjr5M2E078M5WXRTi6jPmA8OW7wamWbVcs8kUDtbVjd8CFwFX7R9ANNVAsE3BpyxceFwz8U0/z8S
LW6cSPARdMbNUIykk7iRyfwfnHt6aAisdz260Xt8UAUfbTfb4xY4Lb5wD0cpSHojVjAKiaUPxrx7
IzTP1/KW2cFSQ3eI/Kkyx2QD6RDyyRbX09w42hBpc3vYXnZNR2p3sRz7OnNcUon4qBj833zxGFt8
Z0MEY9n+StJT6aqew1uNa+Ll+Jt317wbsK1jrcHUZOBYLokeTo4FAVi4YCxjrb1s3AmpQXxdbNwt
jlU/Y4RkDIioqXgAsz0SrWfDQxn+38RVyp7MmA444FaEv3tAw1Sf7WHgIGfkgFAlgSLQf0VTBK9H
wNRe/ssnIdpSSs6iXpqpXM1xeHQED1IlLygJopLxKjBGKAR0sph27qBCkeThJlmC54UK4uroGuRE
1QrYPxXZYM1u/Z/kg8WJ3vMsMOGbz5n6wMDTvFxKDur4D3adsTqNzHfDAk8I//YAQwLusq0rIiPB
LyfOwpk+GCpS3psae4CzU4Lo2e4J5BjqDVw5MNkyYx6mkZUUp2mOE9rPMT5DDuXl7Cda81YaXrsP
MmExAL2uqt9OY2T8QPIIfmoNuctWFEiZFO3oEfDBEKlVPJOro2k38qis7tsqRmmJTv2GEmjkU/jw
EAILJt2JWKaD2orOxzYxMAB+pcgZ1DEz3kspFwiaSkSf/R14gJJr6bJIiiFxpK+ewsAmebW5w/FS
QHw0cqic1cpNneTM7VOyez1RHb3Sg+5N8i96E4i8FtQpIig8dSa/eSiNnY1S939AjSQAk3p2Jsk4
TAdD2LGzfXN4Wdh42QdBgIF/kWH7c5e+/VVfK5PEHul9mu6pqgzknM/2okK7Nq9BW66U67pUTZ6A
875sMvavS39STMD29Fm/1PFwu3rpBXuK8sWIkFy4a8gWWUabVzj5GijabL0+FXrkKgj1erbiGBj/
wB8NZDNGFm2vE/sluscAC7kX8zu6o6259OD1bnDQevLIM5gu1kIDrirN2tOZoCBphMTAjgnR4syn
1j6oAEqs13kXFYC7gLChnDOKk+GbeoSQ3WoNiGf41j7GqhQIDJYZfh01/znbP+o2uPxo2cyyjjII
+enRUCruu0E1RX+E3r0/VgpWuNu8tPCmZGiRZJeBcTA3aircalowaF5GnuN2R3JxJLt+Y0mED3Bm
ifn8+LA7yFJdcisUuXLRu9D/huGLX84SpZAk6qzXWkJ8wKhv9GHt85cgc4xCy1ju25DaaMwcEu06
sfYES+fTJOwx8+m9IlWppo395JiDRxM7CrY9ytgBd0A9ZpK1piWM9abMLfEbILHyfk1i3ZIPY1qq
Cq2qvMyEyATWPodvohXxXKM9DxrT7mBFqGHd1Dv8GiHhgLeV4CS8vrxZM5YcwcrTWxw9hDtViHZW
bQY0yrT1eWqYTzY9ljJV0cdiHoyOmhmQusoVVr4IgNDCrvNKxBhtT/2sEqwFGt/GHoHEVJndjr7n
gQF82EXC/spK2wX7S9FhrK4hCUIci5Ats7HAP0uUqAa99oFkt+T9rH0O5UOrpx/Rdv2HbpiZMp/K
ueI5do6i0gls3p0X26F6JISIACdHtn88SgCBLHpvUgPcHvK3XjFsnRtUxtH7EjpxO4zB368wnz/3
TYO4UxJIFoYdrdCL45wXVEObsqmdfxzlAue2FQKx4CjA2hMMuzjIkdf/49Bt7CcxQlqr25kqpats
An14Zjhglqi3Lm0I9MsHqzimeykk4u249hHYC2i2If6wVCzqQiYaVd/8iJNYkioBQeg+R29fJNcv
peHjC+t+r9t14PvQfLhmJL0Cxfz28pTRiHFVOY1ePYCosV3bwW92OQMJnjbRPAFDJp7nrxZBl2GK
1Li1gYNjFBx9YIWjV8Qg7yfH8VZ0zvw2jg1CcMIbkZJhLAdbt9qaXByDGmlrt5rfr3qyVVnZDyB8
+iiV1HyjkBUFE2Dm9vQznovSXZJU0tM0pQ7T4BHkf9UskgUJ9qDU3OG86xsVmmQ/AS3QenHGe2DC
v+DfL+dDi4eQhZJ0wcFlLEABeParVbZ25OzYqjbru/Kvz9EjantZnlKYrhbCoVpUJLU7Qqv2Yich
NhjqxEEgveHMQ8S8S004b9HSSOMOOCMsR2Ub3lKBwVjCHN/HAy3JbTBxoaIZ5xIAOmNQtW+aJ6cj
ZTqr0NzaQyF/cExzl/pixuXo4BUcCaElGsTOpDyttDw8y7Bg3IJWM51aJwNm2sLkrp+d3nWXSv8m
pjuBq7Psiet1c9q4BEhUWMHeFABQFJDlBBieGUBmrf7sF/dKM+Obkh/5j1FMuPq4uGpfPUgES4TW
ejBCFAe6Ax8krkNYGUiZJFl03IYRkmlTlEQK4ZhyL78aAcRfZXiuOtgqkCjC0Wwbx2pU7k+zBxev
XtUywx1Btqj3x4eJA998YTefE5ERWdm+zp/zIQw9M1VTb9uIXvsSxifBixayoObUn5iaYgjMwfx1
UWf6uahrJy4T4Z9hn+/qElevx3u46TbJFQ7YzUpUdZfBURGnqEKURKSbebS7hezUMVrMVfqzV8C0
HJYuXeBN8Tmcm2qCXczMiXxFHoYTeIyaz0ofXdLDXFTKiDY9m6PoKTX/UKEWzisU4aFTmu1IaU8Q
etKN3Sk5xAFF0MTdh6x8WtyiZWycfI1RqrAaRc2r3OVboS6CgZXorCeh1Wlk9kNeEy3TGcYgoHPd
W4KPyh8N3g/1dw59lqS+5ZrlG+6F/7WeHKDhNHwY7kvyxL+7pQHq+DsrqZn1eZhDSPBx4ZSzEZhK
INRjxV3OaXIhsKBoS7NBRqSw20F5kekPAiGohSpJLUPoVTbeOuxdnszPxBx4inohJcLKGFQe2rxR
80W6gWCapZ8LfmDN3EuecXRmImS5gs1odCOjfOiRpYjHRhdKn8oblsxN+20pu6tzc/fTP6WKbu5I
x7nQJEJ6EFk5Z9ytwgS/XGKbggkdQ57gKooT2UDy8zWu14pcDElGchHlLFikqdy45jd7aQRNUDgX
finy2KcZE6MBEXYjN0OGxS2gASpbwBwg2gB2Hpp86lYPmvGPcqv2dO2hzE5FEKPhmWCiqDdm/j8T
k8X2FvSYNK1cA58TKcyS1q4Zxm1NCWylh8p0Ci05An1GczQhKD0X3C59lIOkYCs/yGzbXqDDDdBZ
mT9NpQK47I7FczF5nlHhBU+d9tBqorZYZqGrOtHfDXQ2k55aK4FtHXTiT70MwHbv8aj9pkOhGIUn
iDcEwKYz4wcTEd7aU3Lfw8GtdnpVANzTFC7R/YWT5OsRS4eoFvsfBFFc9wza6ytLpXUZZZsm9bXN
kx0bb+RCHwwmRGUw58a46PJhCXm8JpHu8F32/n7xY9CdpJn6VH717/aH0uylkancrWvvl5Vz9DVT
i+2Y8DFUgsNgwBvc5dhUYgl5maqkHvidyn9rHga8mFzYUd9Lb/hP6YFnd/1mkIKO3fvffnJbCMCa
5b1DQ8OjGqE5mhxY7uzEZsnj02VttnYVFKLNaVCTw6CIOhags0ct+b9HYxJEYWLiNwrf7pymoRet
UyblXywVLX2Lpy7dCfs8HDJ+F8V81SXkwPgY9CrjWuSYPyqncQvWVeqeGv0B+0MdM7uaUzfesxBv
YJ05Y1PJfEyRdhHHjypuVDvhEgqX0AgV1BdppHV9BqupP8QIXjJ9tvy0idIuRgE8lDfcgkBwofiE
fUFuNgvsb7Sm2lCyjGrzYhoYaGYbbCwWgQATN2oflvdOMTh4XZzo/cqtnFqbaa6TEdWo6CwgvrVB
OZQv3j70iwcGExoIQ+yfAxF4GrO+9ADzpCysfbxKWi+2yGNq5vOKG6VyRmGacrCOtJbdJbHk0Gfh
gh0Sjd2rrdS8OxZCy3u6fr/uW+CF/70x/k6arGhDuVwBa5P2gVHjnsrhoMzsAypOeiU/Rg5EEROy
VQ4wACD2MuDya0pshQwymWmlVmlVfcCGvIWpMBowRuMi4ONxk0D6isznUL+GmGe76Ms4BlPbDhzI
LJoJRhOe0JuGyxreT0aIDgTLqm9rFKKlbIM5Rs0DznNZXSEYYO4amVQTIgwL5NP3LRu10bxgivsg
RjXewtz5Ynri2v5e+EToJ2lpatTZKT40ION+/JxmVI4gfsuoAigoO64t99vJNSmarLOCpWSKe4/2
O/zeEgI181XsCGpLQMR/riKau+wQRgmNg8EBLzYDTDT55cL9e4YC6t/rxP1kCaF7DzTt3gFJvVgz
kzoo4ojFRcGadx3JIGRdmfuO7uarla7gJkzn20GcypjrexjuuXMoXI8862k2HheXnKqfvoKr7H8P
O6PaBl3pbHVU4VMTRfT3d1XsZnP2Cf/7MfI99uk0+UOXRNHOkq5J1F73ZvoKU9GGI2SkpJ983YsA
YWhP/Ke1Nohu3owfkpWGsI2Q+cFG1/AJgEhG1p5MPtUIKrOp+jIVZTVOIvgSHNRJKpu6XohQghM+
TcBrrFyEWWa7p0rTyjb4cFbiqqjg8UpSos/kh+QIPhuPIRh9Ahhs4MOGhwlIHFEw7wSnawRzHhNj
/CbmTW7qwIMWckjLJTrxzh/LmjeAN59C+QunMWaJKes14UP9CvWp0WsWcDVpJf4BHg+x/Wqp3JsB
Qs4M8+OID9LhsX9X8fSUW2w9ppRbcoCGSQzJBx+OecjOmVq1DGUjhd2FK5qhE8Bu/A1/1Mce8dJt
byKH/dMbTTeDueT4ktPZsEtLA9TOBvU2oL7StZi4/vghNZucEG9QK6ze6qtgthOYSBeWjlRMIeky
n/mZud1TJXu0CWWugT8WffrEwDyYO9QTaLUJ3bRAuSHRQ2NM3tTdoh8Bg9Fi9IO4mp7nMVtLFXSd
tJHG7AwJIZmBRNZsiCqjVyvc//SjlAom7uj5LauGH4BjfL/atj6dzkMfHiyDyMaefgZndVuJjIHN
PN4xVhn0g8i1ICXAgp+fmupw3TXxewXP9kQhZWgo5DEEMaAjH1B17G9KoMUeYJfKyGLdeykeHYDI
NfIlxFu9yOvMSp6f6bKZn+aKNbtSbkmT7rumtEAUzEnCygJ7td8PN7+lGF9FhvdSADpTwDVLCsJk
MJa5kH1cS2cSSt1lfWD+2Br08QVeUM2/I8yxK0GjrVXnlncak9cC6INZDa+OHGpxqRpit3v0VFvY
28nw7xV3ex94aIlbZPkEa7pp+N/fidltjlf7q1btMuahQru/ua7XUsbEla38Xt2Xn0+iCG9tZcbO
sQJEKaRpaG9cTJflimzzO0Oda121tu/Rsvu0TrUSl5zmjUUX3Zl/GK7TZj4ixPsBlowdsdGaKVKm
BggrO9h6IkDVEnVhpoKdbgGvlVvW6WLRTmDK9QESDqSY59TPK72t1mccguV5PYW0o4hrYHLJsS+v
cOJvf4hwJehbH1yH8fQ3j7yhUPdF3vW1tLnEp8n7aigPlpuajGOsb5tnTGAjJNHxXdCuk/2UoXOF
fdnZJA67odMBJxulcC6nlezzoaJNtiGs4n82xbBfEjTSuok50MjbPtFKwCihb3AGCb1Q1SKWaar8
lPumyPQbtzbZ8D+F7H0Yn3t/1R24g7GfBYSYL20y/AwBdum4b0ujl2001gBKA77u0d4riJNh9kMy
2JczLZLPlzbPTaKOIsmiWCkBUJC+snbeSLkqhjzbyfkw2gSTPMfFDtC2uAksTHoV4JJPpL6PnOJ6
c70zIeksIsgFVLpTuaKXAA4DRtMLyGinTLsXh7RwIqf+dNpsKmi77xVkAYmoceKh+4Ufw+AFJ6mB
S8JUAbvom+DXteVPr78i9lowPF6bH2kvE4byb7MwFR3uLKZCZXPXTIFJ+YUnsH/1RzIS2kyXOeB5
ElQDh1rGwAkSo7QKCTjvLYjepRFqLUp9aj2gekZ8bSBOLdukr0ayv2ub0hHgFiBh9DUPtM7XE0ZN
/X3FWuAdMOMEVzOGAqDg11jEKaE1ft3eVhDbvzPvWqg9viMWM7w5ph5CIJKQrCvK/MTrIpX+wDTe
lQ8uRR7HtKfE8S7b8VbMHg9eEubxzgelutiACRdPgNPN7E+wdPRaaU+JZAsI3t7GBuBRewy0h8+f
Q/EGeo9UVnjikq+KC1Ez4erL3ax9sKd4dswfojgqEfUVpc7uj8HLk9h9+3wZtvScV34sgmQlcOmX
uxWRyvnpGmbe1xBDEN6vVWIR6M3sEtyLpaYkm0SAdmzWj92J9LBslf0FsgvY93TPR4LA0XMwRMsI
ftrTjjGSxn9R1b/V1z/9lvTMxJ2q/CiSOukkcvbWKbOzlxc4a0We5OYrL5EGnYkGBFYIr0hVrCSx
Tfs38y2wdZBxJ3Rh56m3IePcJOP9/NYiKZNtRDBP62Dm8DG2/+IsdWl8wIMgCh0KIJlcSSd4Y1OL
BP5oalIqw9y5rDEthg94hIMHZoYVurn5gd+NZrjNSvtlg7iE/7EswcAUACWYd7wM4HwviY+29wp9
+Fo1LQO6rc3BzsKekPewHNNy6yMz86FayvaQiOWA79Q1fjHVggOEc6fYn17F+TJS9D0wb5ibtlbo
k1o3PRJj2xf7VDm1oX8MUdiFFL1AffAkg5CwC6Z0hWu3QzvW3TauJ4liGSkR/GgFeLtAxSjTFd6o
sd7D9sp485VklNIXzjjlwCBZPRzMxntWd2GtBFKvhU9L5vhCX8o0MZXdUfI1R/51O91760XNphHI
MEwwGXjN+3Vx2WwHAPrZZTrk8COTpiD5PJVmnhcPMqOI25iViqyp2fcEjq81ckmJOhG2cL7rY8H8
9B1ZS+8muzDmdj/DKUlPcDy5YSiqzB/pc69tIJdwLaGXpyBF3vmMvmG05IQ1mjqMMlPM+7kFfaGF
NaKLBtsuqdcj9MDHub6lIXAd/zzHjdyG32b2jNvnyBpeq4CCo6Sq3u9xALVR1YQBfTbQgXM76hbZ
KgG3aw3mz/4qu9xf2XJt5blZGrHcYDp8V/potOlSSvU73PZiJgxnx4tOMbgOipsb/1y7Kwze2CcQ
+7NxYAYwrL15dg8dOfLAoaC67E1L84hYgqj9B9yHltADq6pZJDM31zXBaxsZSS1xwP6ahdVMZRtV
GgFRMbg0EDwkx+QZNB1ZRdwMo7VV9AQX7lVxiZU0WnuG/JeJzRha8Y+hWZ9DL9JSmF0CWgdC2Hd3
R73x5fK8jyyS7TWXXknWlLG6P+Zcr9zfda8YA08jaE3LIp2SM/v+pVJK8U0AkUAJPWkrEOH00DIY
hv2ZStBgKB0chUXYLtzYXHB/yesWyfRDob2wyOLuosjqzK313hHq4Zrc5B7Z63IsZwOExpXyNei5
kVQdF05hp4ztjK3SUV0TABhMqn2/CB7xqX+PZotEn9+MdQiyDZVvaJAkF1j8KvsJ3xDMeWJLciFV
PeZ3fmisUTK+VrrtAAoM0Juo3xDQDLiKQdzC4nJJ6JaByBYZdwYABGmMXPi9v5uc3h0WYxanJnoW
pL9mf+HBhFiDdYHAtdC6O2JUXdrJsMM8PrbVjdLWsOJx7EydqvS52gStiad0k3VCzaABCEwmp7/8
TJ2L/L13uER9Y0Wiq6lwUhXfbj0RcpScpCUCQX0LojIXbHr1/t39W9NEKt1Hg2zsmKJtECA+r6UH
ikIFLxSGmLpKHeaANuO4L1hy4Ej8jqOuEaIulb1vJqj5g+yP2++yiPa3Hq8exIkZ+4sAhHPxIdX2
BNR+Y6qU0ysoCLgBYZkoAjtofCkr9K+zkklF2A9rJdnHb2qKp2ht3PuTPyOHvqGCfz43KZBROC9X
ZlpWxd8WDBaxcztt6Ir9Kl/AFMDPgP7AuaT49xWFZy4MPTnwcwcY/FdEneB1bnKB8PAZSIRRO4Qw
68SjfpaSwNuaoDwZnbp2LhdjFVKnc7nVAc9aMTGHNYJNxWeaStSMADLYOIijM+belYT7dxbDnGAc
NidvoLCCoQLfZ0U66mGpgzRlzkyrKCfyXc407QNVBRUpoQtp4qJw915oOjo6efVlmWo1ksg7ItfC
eoE8nRK9pXVWSU3llriAApLpSk7wNqYgWv7Wkjqzw4xMQGoeZGWDskxAN4RbK6UitHLBlNiDE5sS
17Tj8mOtbjxiti5wQowqn3xC9HnqP9MWHRduh1XN98NL8nIIm9l55WXh8m/C5VYt0rB64PS3EF4e
BHMBi3tFC6TygyhO1l6N9IIQnxNHfdp25o4qXBQzJWunv5bbQMmglI9rR6dUUoCemqMyIWiT7NiD
YFY7HUNml0jK6p5kJnLI/Af0OIihH+K1HPQg3DKTCBxdFiRpqOxq1a3UN2N78QAWdjQbJpk2xX6p
9hgBaMOujzXW3ZSP5cmtdV4Cg0bLrLxb/nZQVNdvUlnqu+898lTwTgt6QICMHUkXYASa4rXNP3Np
9EfBPzx+/R1T76hs8DcsknFF+QaM+KuZldXbRRRyEFloseusDx0xnXrc6ZVQ1Ip0pRFP9O+TfKCY
W8vZW26Kq7+jiM4HDd/IbTAZfMllIfDrKD5NkELxjscIjtPIcqU9ICxpOnC4SxNZf03pyNt7BQxJ
h8MQxsWmmRGsHNJHOb9sbC+I1xu3mrnl31agRQeuyXchqxdtd0PGdexJTt8WIL7s8wjDFCcfRtdj
hfHSdpXetCX37V7rlAcXLw4hgy8M9ucJ7ngEQXeW6XkDx2mTxfpW/HNlryr0ThdsxtrRymHBD2FO
sIS2CUPy9J+JfAEMMkVqo4BWmGE61jyvdDHf6otV5SV30wj+cgfppkTK2wSC0we2+IiTMjm0pLUU
/QWkcJzwWBJ/rtolNgfVKBwCSmLQseBa1RgxwpzgLF9Irs6X+zx2VUxzHzoS/AMgZa/cT9KoZrDC
S4rVqOhBfjGPIe6TRrKqDOQyu6nhgHxJNBLirXZb4TuPXdEMDK2DF/Z+zsdjqwpjiBj/dmvzbF1/
kVFHxjHdlVRIg8yG/4J9iZ3ZB+BBuCO8aAAXVqo97HXfOpwP1bs6taYFCh0Z40lBnklRqrofmFUL
jAYrPS5aVBtquI+4sANaU9Yh3hVlAlVsl3Tgwg8nlJ4XPdTTlRVlDyXeX8PKVG9gAdHXINncKvGr
ElwrGrME+cywGerICiqnmHCyABw9Govf+pFg6vnq4RMdlNx1wfLa12oFcDHczs6zgpTI26KV6KjH
ojBeoCOzOpKqWwe33buOXUehbVMqMeLs7rKcIoZa4RJIalxNY0LC7wrFuDQxP7f6pHsFGjnUWAb4
zHJMUon+ZDhXbNsmlfDbi8N9IeKYdoF2w6+egiZ3ECHblnbD45dynDudTwPyVoODUJVa33QIuFHD
2YaFJlc0ve+FmOXR2WxH27VZkjAheiXUBQbcK9yL0vl8tM+uUg4qNMQZLDpLdgYs6GUdwV6x3Lai
x8aa5QcjGNUzLXa5xby1DXZDGHbDhtsQ24WnRIG+T6SG7sXnMTjXTqaobnM6xJ3SbupHg8s4tOkP
IcMFYi0MTN3TZRp/hhGbwwayTCQ9h7D8DlIGoPQA5Sr8MlozN4f21A/JdnJqmbO0jGx2pYEG7m7w
uCauJmaZaFSkrJ+gXqdlUOgpla49UYO6xJJG/VWcwh9qpPy79CvkRO2ygtfFmaUoZJ5zxhgz6+qN
JA+SsIYY5c1/4sTZcbvkZYZAPwThlqlFXcpzVgVT4bW6kaiflRouTHToeo0Gw3GMU4LMDW3WBGRs
XKaybogHaO2YAdA6Zb6uxQZSMhL4PtJnbc31XgFNsHHxZjR2PjTyV9MtOfT1To2l2/nHWU9JDiwT
f+wx94/eX0xNlS8opA7FqvYg2SCy0VydjV8niwpQp3CP9Gln6mztrSGqxg4Biwi/K29Gg/GgQpwm
msSQ268PW/039i5ZhLMJtHxPZLOKmUJpHWmeINj5UQPBNQMeh/952Qzr6lY3Fc2GdwjrLXQZst5F
p2UzAvaOVO9EKGvG/2dMpd7eVQJJ/xHhUBvtbw4G5pH7439Z+hEcj0rkPoa5/o0mKr3zx5rVgYDC
gdDqPh1X+YAk4kzWw7yKVnlrRAnSHTl+g2Du8KEsQuTFZvC3iR1PNrnbfp0rqBn0svmeX70cOgWO
GhsmUdIjFMqtfmNj/tlUWLbzSrQnwFsXl0ZMnRZ9Q8uRuWjWk0BgCjs/JGVNyIdYebsJqF/InU+8
jTV6L/5k5iyPX0X6/RmpwTz/FW/lSJ1s4foyxn1Sq4zY5nRCXWBUCLTNm2V/P9rMMy0VtmVpQn2f
WKvvrjIJnQ3ig25KzzmI3cjqZG1XYF009Qd9ncITIor4ufvTy4jhYO/EdmJS+UAFo5s3LA0CKql3
hZY3VMPFmEzugF1FgLQGkSxq9OMZn6AtHyo0TPKt+kk0a7VX2hJD1icJ5SQojyZM+kw2WaCl7OqC
tcvsgO/qqlh6c5Q/kIx4z+zFtuYHpfgb8DXkx3fJBw9FrD8dqe5fDxILEbXNOfak7OnH4+6/cDhd
9ypeqLbrxKXBOVEZg5Kz6kH5srMFWOqk06IWPHXQZ8KVYNdLhqq3meQN6HSXnPmdDkt652Xe6pLD
rrfZ+dRd0blopx4ibIf3QUz7GQ6zxiNySxm39Sbu2Wqp3a5+9icwZJrrJ9hQmrHOfmyFh8ekzpKH
TJkUqcKNrwUmwSwc8nhZAwCK2EGD6x22/VokeNzrBH2kPAUGcW5LlZQxz0ooAAtwLo88Gu6XFd2y
tDK4q6qKD3eUQ/cWNl/k5K3XnItyHDlCPbe1zl8BspQdzvbpIsPcwkMFFb1vwL0lC44p/4c5HdJT
5nV/UpHf0df6UMymeLRGlmyK4bPriDW3QZoCDvB5MgKoA44Kbb42mVzzMNEeNzwyGMvgBLtK1abe
0DbuiYI+wlN7VnCN6Z7Pn1/U8dY1s5lIOYCHcWVo7CpmjGNPCNWZbnhZ595xi5+XHOjFdyXoxozO
3jkTX++YC4EOX8/8ywS5J9HB8acRWcBT0zuH5z2WPq3egVtyMN83/EopptK1UbuT2zbQgDls1qMF
hNgunxniIqHpbH3QWXMbRW3mbXxsoajiCUtD8TSJqa1eX/zMzIGQh7K9ah/HGBc+APxZty3TJeIc
MM46dKx3kffo1IOcJWzNmEeFjEHneox6rqsOHBpW2e651mDXUaunfe8NZ19JIvNjoANxYqIfRKFh
DdAxcegVt4efEN9aMbqxuosq30gALzU7U7xXlhQLmPa3P1A2tb1Bi6it1zMvwQscqqKycrQNdAgI
BIFlmN0GNABKN0fmd6vmmztqHKZbalmKQkL+Lh6KqE5swvPfvGOAtKXVLx7r8eB1Z8fzA2iCmhUF
adcx71q5/t57e3RnDUNxNKbN6/LUcSTUzo9kaplq8feAXnetscuOj+4LIfjca3z/X4kpVQX++m6D
3iaCqmGat22R1QP9IITlJGPSas5Ta6DO9jtJHb95I99FxjGPsV+smCPftN2uU0K9GOmYA3vyOfkt
zkbfuO5XLoMD8PTB1GrVwlF1kYoAVV6eaQz2A/E0gkIdiQEcwos9GjNl0Jlc8Mctc+49I231yYTV
8PVaW5yv9m/DsG02HnXdnTdffgVYTjyhRJR5LxY3+CCFOr/IbzYVDAd8xbAc63iN5CqXa36Yu9du
XEOji8sOqrK+LXfgzsLBW/9IP/fGJOa2EZLfJ5unzdXZTfFRQnUYTctnFIZ/bNttOrCEcPWEnwlS
gJtxaJc2WPJ0clMeuqVumsQAdbK1Xe1wDXo/NMZ5/tEvz6/Q03Y4g1Xu7VwXwOGd+Z20p/rVjKjO
Y2/A/WKfjNIE+D9X5EOjb614a5knU43jCMPuCaHAyoGjgNlVUeMolVo8iWN7Vi/thOA/nBhfh62B
PHBGrTrnb5svDczVGPdmbbislYGN97ORX13hv3nwcsn/tMzmmk6rU3TN+/gOMu9mMqoYGrnDhGbX
/WhQ/ct9hWzKJgn3p/h4TZZVjC6e0owaNmUsbJEq4K/wA+irMquBbac3075e/BHn16YDSW2UH3/M
Hrzldl7zhEiC6HfmF44nZsC1Az2q/7XTSxnczEh86yXB0NpPs+Lajt6EAKapLBafvwik40YsPXcR
Xn4pKBj5J1MndnrOqnz3viAGBaWOf0lM1JqqbXpJn+a/rVTRal09PlELi/gufLh4FpypmPDF8FaH
3NDUSsy911gg50aktTDcCNJ8N9JbUgV9lKonzVd1LeMXuh3j9rI+eENFR1ucoJ2rxI9w5O68Q+/U
OihBT9e1y+BaHNpqGgkmLu8SgiBGmakzPKxOcYONX+z7lJ79E3rcGPh7IaAXpnyr+poI2/2jKmgt
8xlEv7J8BlKec4CPqgxJPnGyEBN7ntEVbfKL0NjX5TzjEHbeJmvmTgGO/sCJC2DwPxVEmplMvxNt
s0fTyWUna7+20aJN14L8H2lco7HznJC0eBTu9P0zfn5DnEOShMJ94sZVznu481FHMk2zmRQo6Aka
/7EGJm4ZNhzWqoNn91BUk7SsiIqMyDutMrQxCSA/YeRPKl+dEq4z9LZ+Dk1szx0gajrrhDUUXAu8
FmZN7DmrJwNxDvGxz1L33I037Th922TEBODG3k+kqEUc+On9uB/9y094Md2gcvTygZxFkNPn+z0+
B/7NSLAPbdAym9RtzaebecHB0yb+l77Myhu7Uq2FdAV4cyY5lF1gm6wJTsfxP779jwmIApCS4SYu
PW3Lw6eimQoJjdn+7cyQAqCkuu4IKONkCekUcgvHsPA/iPGn552pbqequrVz0WXQ/lXx9yAO/wdS
dlYI4nwAjlACEy7zQiEqvVqf8k9YyS1avGY2aZdU7Yv5pob02wUiFKT+FPmTkKGPdI0cY7pZEUZp
YjG5fGqq8iExnPk89Bw4vHAC4Q7T7AVLAlZOgb5RClompKoozKKFHUlYb+s3YwR8eljvcZhrpePz
v6toNfXMtQ+qNZcUzlmB+ZgXuOEkHn/TWiSHVG14pO+kFGz9rvcTsf2v5BrXPKOaOQP4zhcXfOvM
g/+79nXOkbzrX1TlvY0BaWc6jo7GNOcKTuHecMysXR0jHr6rvTYbT7i/0mfDRDEMs7tXEZQ22JFL
7B2F/5vcs4r3iZ9noPslmdMCX+BKE4A/eq7BQLeltCziAQFqiSuphSzIDCSW6lqyXAIa5yanv+Xq
pvC8aCA9YHr5tYjLk0+Rw8POqT8Ebhaixoz1EtUYopTn3roFvZVfAlGQTBJAMF38TuY9atNEEtV+
DHxD7My0I5xCNEtYrZz6nfGJhHr114zxcHNQ3pv3IWnXgz/Lghv2jXTALoRhQgwTa0gJOBEwXobR
vIB4WugpYkjid/8M3mDskaHo6uqyBrGftv0wKNiem5G7QJ4DmbH174GJV2goLBbXLvm44TZx8IOb
uHdD5CK31kbaf96otvQKP3oqcuaT5aFJFg7i98FxD/W7tloFPDKGHdbG0CpG+G4nGpU3xVresZFg
y8BufSa4s5OK6Jhm/6ld8Ifg+uTefHK1dUSGWdSjPvqlw9aKJLCjY7pe5WSIr6eZulqlhl+9gZX5
m3k9sWlnS2OEwA7fHz+kIIZ3BigRQqtSPad+V6hW/aMhftaoCkO9WqIl8iiR8F0M0B48gkW/dt80
+7bbDPzSDMULIWWT0tABoyz3qrizwAoXFCrWRypdTZNLpz8IWRikzXwjiL6awPqltWSztv9f37g9
p5oJg9LUXfpyYjQ1E7StquGOIxkxV1QiCOYb3j2GuSVQP7JE3Es919yEOetTzGot8S8b+OdpnLyO
5EivBuZBFT4Z7soveAj/GGeZCmXgqZWewTBEIyZjrZbMoDbHs966xB1apYSH8uPOrpUFN8HkE2RR
9qNcGoeyDTwX4IF9Rp7Rkemta9pN3amw166oDOJOmZxk1A3c6MdNAK1SZOMP6Lxd6s+DxAusNfDG
eoxWiAgFXYiZNYTEBJq+OtMbh8VYvGp0KtpTaobaB6Mi1wFQ5yGQjX2zM+XlFEhMvkfRb+DsTBTd
pGO0qrPyqiYnD10B2Wrxs6PZ5TocDSLX+JbqhURo75NOenCsElApip/PQ+glZMG8dApyTNJf7jjX
4+HMaJsGDYwPC5LDmMgjhkCqY51SJ3VnVQUEoAery6bVAvsdqnIB6zfpMxhv6yirXKmXc6LO2ywD
JHpXJD9vRkeKuvbIV3de7CVGFvs1D5YVzZm1WdzC7q5ZRR6g9XXEZbcDSSswV1gO654ynM3mP1wt
p+zk/q1sRKSqYnxMmUE+NIAJ5xF+rlBh7TNrMQiK8ddCzZVKYCM7mVHc82wrkSt5TpeLnAnWGChM
KMCammZr4uDwIlDWbMzPO9ixYdUeomn1adp3jXB/jdugyT9RCVGQ4HAZQQYNwYMWViTcUbiRJENL
ycZJYz3DrFv9hP30KVf1wnw8IhPvvR29xmuI9/EQ/rpwMllVPebzkEDHpj67WYk06UjYojV9N5lV
+x62UbBAWqMQE4hV+zzIOGUvwiQa6g60VJFgL7+HnL3+gi2tv91dbTDOqPznb7oN9QNKNZ4A/2hX
BFPD4YiaqTln2Fg9IPppVTcl8v2BF+fBsXqRa0Y6LRJNJ8RiIl8gNqxE10Cm9GQLG6AwEl1OIgye
NNZwyJSLZbal/AqzM6C6qm0Hi2y33q0rtaZloK02OVC0kmbyY8KB2LQd0Uo0GFCeRmLdwQpDXgZ3
pzTKbXJl+2OvJPOJbDbePP85zpRxG5QkGRFG55Bx9n8hhWF7vCziU/MiPg8Vm08BwKNpjH+FLxmT
u1vLQ9cYIINXM6bfC3YgHiijaQxn5PqsoK/8yR2wLDBlEyrLouiCV/pEgd4tYIkhEssw36VszljG
m5oWIX3NsqEvuZ3XWZvqcVZYEwFb034yXSIaH8lqlPv3fHUFVQPnYJ34AQUAV6jHwuQmNh7l3LBT
fYe1RtHKN87JId8h+WdQZUrZEzUK0w/QDnNU9kMsB/TAM74AOXuesDXQPK3sP9XkjREurmwe5ML+
5pWOtzKUUltOSQIYjyrADvMHyQ3B1DTHey5kbMc6eEbO1NST4MuvnJPv0XY9DtzrZb+HFy+WujtB
srU/7Am09H139G6+Dmd96sYYQY2AqIoKvTsfacZAxDYR/W1BE/s6be9N56OpzOuxibDJxAaJliA5
He+qzUxAt6w7f3M5a3Ugtv/uLjeUS+mtd6ruyQDRB/EUy83oC7OSxYttPar9E3d2lQbMEgm1a7wO
RYk96ff0RPTrSYFvdTmxLIzb63p63xZt4lK7w8918XVzOkpBW0g8xQwZ571pVfLGJoEzQNrFZ+Qw
rRwmH5Wba4q4DEssI944FnuUgfhOb168CCxAHpJkURQnKTDwMhNi3zTkucY4yUObUOnqbifE/noT
NGAquz2el6Xt8GGd+k12egJSl3G3PvSH+F+UMj/kNjZQ491Oz7oiZ79auV2rT5g6esZegF+djGdm
C+IOd9f0koOBvBMCKI4UkZPMsnHm1/MbGxjeCH0y4zBJL3NZfjfQgHePNhQsUNek9R/7RkIDt4gM
KcPVMdQLL22qQ/FzFLHj3ianDXpUv1MEboI5D1llUfCEmos+sYzCqT3uGYI02CAq4FqL1IBl+JtF
nV9BbjIhbkC3IQXTyP8P4+pc4n91seA1cUbO3xxx/bDp+hR8eUsmENTVVMqWwz+8Q5iFTEHNVqtd
5jyZZbAoizGAYoRWDaDnTfXitr5+iCleCcewUXRBwl5KyzCe3q+YjZxeEl0jMkJC6IvkbW6ZT8lf
q7lDcVBXecW6v+VFb5Vv+/JuD/aaJQZqIhdIbvOufZfSIh2Keo3J6Mam+emuDzrQ3vEJZNcbomBs
ppCEBwtaCw0KmGwZFnowFMQCpjsxfF64LjAhoM5Vdyc4bAYGYsxZCSe4BdtJC1yl6sf9lORg8D1Q
DugFTR3pLrVR+n4Vul7udtpnp0qswNuQ4cNSIQTt5zfoDyPo/fru+UFEtc0GCi7iIcNOCqFJ5G4x
xSqJDJ3sUsShhQkDJDXshaUrAvqHlf+amN6kG33/8qDY4Hj+t+9J/EYZ3tF9/iNLv5sMwqZCqbx3
FtkMQ3bi8lvVeGjKJNJf7vIomJQJQ2V71r9AlTvbOssxdZnX8qGxX1sMDt7eTuwNyYDxapBi35/x
wklLn7MR6iVJGf30NUt+3KKjOpjsYRJtUTBPaJbKYv0D0ihle8waf+SfzMIxRAuqC2IFzfgxgnvG
u/qtGPD02eJ76dT5FPQJW1hA1AZEfXnt0/UfmoC03+gzj0VKweEcu2/y+qchhfeSWlMRzp4JwOhN
sJWHQ/EzETEf8ZBAWnxLYXtmYYlgZDuZszlWDsg/yYIuZlrcGRQdK2rBd2ckX4lh+UwV8BDMciFC
CMuVUZkpiFW4q50Nz8pyz/+d4OC48aTNpyKBJRICnL0/IQU/VkcVBuWn8ZDDeeVu4773Zax3LkOE
4Ri5T3ZY7StLl4CQkPDbYU4UW2sQD+cFPenDV4HsVj7xarRh83OzDZkElKYwBdU8mhMcxETfD5W0
25SxDbYM/QMMguWFj8xkTOpnVFPiTIAH4WBhUy3ecE9neia5Lyx0SvQEOkxH/QJfs1FSHt1cJQZZ
OPyXFmNBMmoacyFKrRSN5IWsjCrDKE4aBiw8jHSyDjWx6YR//kL8uToFIxp/EBfH9X4I0Pg2lwfy
HYuq73l0B0YJBbFfsZftFiGmZL6xHveTwUrlF1jku6a5kj0H9iG/j2VXpSxP2aepZg/YJaGHqFMa
KTarxQ87dgFH8bHPcZz/PMcI9cQPpnvcwPEJpClkMAcirF+E7QnCgCqo9a+Ce9HjymnEv0WdSAUa
5Y3Ls3/RqisGMZAmAo3/YgXA6xJ+CPmVFeBj/KDCxEQNZOKtVoLcZkAKjpRueI9bTMhbJzZb6va0
0LvJy9KwYOD3oE7za/262XnvAqKOS8fSPU2+oPA22ygmcAQGlBgNv+0y5Y4qt1Sbda8csaOlQ5va
8rhIejoVFJRDEzD310fNhCzTkFveNmNCpJ6LWfIPgtaHQUHWHaexoNQXywG5PMDTYPO+cCR+Jz25
Q1C0PVOrxrsqu+87Uy6cuusg2lhnt2S1eFKjvKhdiE7j+/o1zJ7Cmr52VSGp7rz7ufd+cwrDsCm3
CnFE3NkG76xMriFstrE+iu75ohA9cXhZe0EZKolo/62GNp/ciu1z/rv9cwl3/dDeHz9hoTGetUZl
gPDCy1aqXM8V8JFc4wEjbr3ArpQ5YIsJw+Chg/GPaBL89KVVTLSREJWSbnViUFOCPRFsX7QoF3p2
IZT87BkR8Rf/JBiSB+KNsBgoqdp1Ufy6TDu0GpL/RYdSZirXi2veAh/vexVWWCBHhWszFcbJQMPF
N83fbqUXkh/uFWKLTQJeGOE923lbF9n+s2A2bcGt1/4q3Qh20/rzqL1g5eo8woOcvBZ/+eon4RkR
hZPiEjaFCbShxwydmgxmdxJFaPXLoJ/P8ZaldgI7rNJ7YI0NT4SDIEi6QnDEM7aStrGwvPoT5+xo
6PfmP9ydP6VKdp7M43HyNPFN9vTEcOHgWcy3LhGbNOgAL+lXX0ziWM8tN03L+mVPGs0QE0vigPYd
/fANcDKNo1AsFq4i2NF/GmrdwR04ua8IMc0j3X0bFe0VdKobqyAHvhR5Vb+XgvpcrDcc/AqV3ne7
EkLhnuIjo52Nr4X5k+Q6QR7id/y1gLq6rqRX0D/+Vwjzj+6qXwcGt/wVAqHCDq9W7RH12DcXCwTY
4UFciyMlkeC5TOhdg+dvcfSQHPoWb7YzUoxqAP95feuTDUhbcUuJGqn+lovdk2guya+dFQgHt2k9
DNYZZywNl0IbPhwgZj8U+g4FdzFLYBnn9rKbv8GoH5b757/vZMoF2TU090Eih/lqg6kKGyGtpZo7
q0dtgyjz37AD4TuRtprzwTomCwmPqlp1SVJON8IJB9yoNiFouRp9LjI22yscQQHfovYp6pPOW1l3
OVNFxuneiLGQpB8PIlcbhBqgLt3jfvIWZVJIgsMlZ2H0rrmyjwLGE5VT87QuNIfj1c4go/XNr+cE
0M1GK38MHBMVbpDMfkjMyiQalknfP/GIs30MOz+OqD1hKOkZ7wFoyoUn8poaE+iAV8w6ZPuKn3xp
GL4UxQXY5F7r2NNFqyvUyutzYgRbVWuTVntAzh+9HjcILAtxmJA6CDznDjBbBeOoggkNac3kcaev
YuS0prGIXI+2cJIUxWhD4CmK8gdawltFuW6zo8sKuGmZ+yxMTwGI/l6La8N84Z8TPA3OAFvFkLC2
R33PiL6+Tb1gvuxMaa2UrKUhSs9VDQr/SY5ILRQQOykrHcTgQMb5+TNfLZaUxC+z7AqB1GYq+gDv
zidnRTrojRqpjF2W/DTAeCgma/XU78GAXc3pXS++wcpCZeDTYzl3umQtGJtpDlGtosSvsqRLGhCb
uaiQkuHxAjb6Xu+qHedYiW4B9GM6sNmEQ2jrZZz2DaEj9v3GRmowXVsr6tXWbGDZbpQlB9kQkI1y
VQHV1h8lnYobGEpwRdP8phxhObG4UJfc0Ksvc23pB/fnp0oz2hpH7qAyU6HDio5Ukx6gOdgzrN/C
MRuTb0cr4MggQMZJRKXZtEKp86PKWCDe//ApwgfMQaKmIeTnSQK5yCOXSw2+Lh6R1PrkpcT4Gpig
2+5lrYJwEOqlk4JXWHHjbXUwbAjh67z3ysALZpBG8EAhLiButcteixzYxgPFaMS2+zQeBeyk9ytv
qMC0ZI8xUHp2b/f0Rhz1PTIHKLNDoS/TZ1h+KS2wUvfwDnoyX9tcrRluSpKt9++SvgTMFdrrHBMt
eoHOQFuOr85pDZIXdZwXM1T9xNUhd9MKvqCnpumArs8qDPufb+kFp9IZ6SP9zv2ZQRilChOZvy4s
XQ5+ujXoHZ5a42jN1apvwwG4HVlXNCbtU8AtAs79geuEuj+pVn3OeTYFQMJXOkATAHTcHCVokX8W
d3ORIwbQuyWgLC/swCgx48MRXYruCLqHs6OCNpjgGRkSZccFfMYmqNlEW2PCGQGedyZttTiRRYoI
5GbdtPJJ+smQ3A4bWd6t+BAJEKysYx5XnF6d08UEmal8df/WlZH/rwKEE1+AuNq1DGvmBePLCaf5
OJoK0D6fcRMp8/aKZ7h5cznLC4AQe0EbNKK4E1agOsxvZ5SK8LayQ5gUzjofYlK3Zxrmv/MJrQ7d
jf7vCrECUVXKXrsS52G4rPkTMy0MGab5n8QmyHl/NKXbiBNQA5ZxXOw4JtgxU0QGsXuUlgBiIDqp
wmdKCOMxR0z+tQgQWMVN0YKs0M2jLZU8y+EifYQfcYUvVRt76lY+dL0jDOE2kiC5jvPbpmr7jCLI
Ef0ezs/naahSIo+jDbw6AdbwYewbreyNIHw8kpp1GhAWhBefxx4vIrf4+2ODEDVkeVhhCRbn4zm6
Lh4iWud95KzxOeWOUfDynEBKKJjNqTj/+jjbSLxuOwwLJKpsXtzohhNPraBQgUW49WjgCLx9H8s3
TkensZ0sXx5k2VvocuPDJNuEPaa/kOgTP4jwdKGylrzbgWptykB7dRhYS30UvT8v8SMJYZUz3j8k
vgcSvkmAdC8JKj1yHfog/jxa9RyYrA3uiLtBSCBjHhm3Bva5Cn+BNuB3EH/X7vnidKfVQxblC20s
0OQ/qbw5U/01J+dNPKKc9b4tUTEA4MZAcWBTVOXq/wE3hOEclo+QcEYggba/G6H1yvm3/XB2mZKY
p+Zl0D76/uE9K3jPRz2DB146GSaV1bo3g5mbB3UKTdCImMkZT1cz08d3iiWmTOndseiGEMKzThmK
u6DvECiBkILiQ832A8GnPjwRz0LMXmwy5OnebR0knDDhu7MRv6RL+P1ffTO4twChTWmaUk3JSYeF
FWSsjcgMl3QtO6zPRyTWlIIXFbHEG7tGhUmFhLsVQEjJM9gAgsZd9HB/+NjYS41nih8eyB6ZAwHs
7YBuVbVB01Q7+3Fqnf4P2mNkaGhuvDWiD454bOQIxSCro0s9ZEivCBp2Yw1F4Ji5Qo+aCVao5XTR
u1lJHJD+zhpM1twP6rScLPdMvI4FMmZ5XqGjJx/ocSMLVb8SbkCGomjcQcwc0OWdxhbexFzIJmrq
owG6gOiDUuF9l8jnk5KqclNWU7otHWf12Fc2naiexFl21/vki2vohvoZ9dYE5y4hCRQAoQM8dfLK
atc9k3/s3cpB9ckiIjj7MqbuTnpzE1pdrRymL3NkhC/uQCvFE3GS/0YKpJ+KCWgKx9ohh7mBQakg
mCvQV50OUo8Am1vAkJUteVhHuGzV3wKaYKcDZ6te2RRmLvXERLyeTfeuBpYyIm6uIJNw8Zmghhuc
FbY5YMWtYVQcMPZVXswV1h+kbzwBCy67rDUnnsi2CqKoEpUectjPlb3oaUEK6maEPFcHkqFOVGE/
jLWWSMoMZVetXKrvd84NK4Wle4W/t4tSrxSm4uOggTf8bwZ6aXD2mIsERZ/0x4LD9CzF0o0/IU0a
IC+HVLTcjiWC3Ouchyi6ukasTvGy5LV35aULqrmh6AUdMpixZHAvsD0jp41XbmQleTSLAFHP33yO
jQuiO3lGl9C/G06FW6r8aeDd/7/YELlNClJCggQFcfWLFWG4IK7i8D01rBg4Kp4gDFEqdDIRLwV7
eBQrO8w60LOw73MZTKoxPe/ID03dGCyiWbT9VUR1gpljtScdcnRijiXpBhpB/8QDUWBt4ybVrBNR
e7IAhe0ebKXyNi3wrWMRMMMt1pVssPAAnW2JtFrL35v3KiGV4SuVislfw+ME8cPF3RUFWse7siW8
xh66EYcDW+tdRGpPSq0VwsoJiXlHmUar4Pt2Hd7u6Pxov4vIW3qFt5ZQd311qZVNiEQK6XggaeQt
ooV946wFTNbrLBqcLTINcnurC9wAoFp/gWReNYDQjCkHddgG7CsNgN/CviWS339ssVa5X9hyWZpJ
NvO8kE0yy1Mfm2S7D9MIZ0XW0RwBgxmgLUXarvzycOJB4PhhlYLCD8ylu5NOOh9XW+it83ofRVoG
tnCT8RuU+ym8DzZ3Lq00jAGQ4XeVidsFqs6U+zcRtLDQ3iVXN6tsfLKWP8XxmKbwJesB7lu8xcJ6
fBVmsDaGBymfidrgeB+R8uQBQZICuyn6JsWFa/ZOXpuZyj0t4Van8cfQHSoPRS/Jv0NzAL7VcB4U
t/dbWkYWl8pR4K9hfsifirV92kqU8goF8PpgrXpccCDrdNHTSN1RIi7MBpJMDwFkvxi8RpXgIN5p
wKX7Yk06qWu3WJsYCTku2k00nPmQ1v9nuMWafcKVaYB/EAzlVaSklvLRnngtPkOrYabGep39oVam
+krPJAjw9VIYD5fYg2abXF1kmKySgLKbRmt5pgZrSYp8LbFhlJrZuay3/8a3iwAzoxXJ8C4OwFB5
nKZZWB/aaADZ/oRpdrOBPSc894Y0gizmRR9n1fhbg6uJg2WIK/L2i7K1Wuqgz7AZehO/M5DAW4J7
5FQPkegkFCj2u7ikijHUAN1yLsnn9fbQBLBKgQIQbp720aIqPhlXg6TA/F+NsHPMCv2AOgX/LeKT
tY8Zm05kSEgrocGl37NSsfafjWlL/jDNVTRSlSkEarNvjG1FaYbrxyArt1BqapTI4V7/RTKc6a8S
nsAzkpuN1pM2rG6rpECJDTalv46x28GwPet1XC4xu+flIh0lSgV9T8fSCzjbJg+4cw/ubQ7+uVST
ahTYZewhAWjez42wV+9vLHER+KR4EnSiaU1jonW2we2/ZRapMzYyd+aK0Hf8+bipsGn+6YxaBOuT
Arr+pwJFbyD6BOhzPipWdfNQ+AE3DcCxIqALEJqSXUkG080eysTD9IiyKcSLetD8pR8fetcjQizE
GZqWp2acVTDNf6grtavUUazCSAKZxGmEeAJI+JdQmFb45ZO+SkZS/1Mo/H2vGUjipf7ItrPCIHdG
4qLt6A22bA/9TDtBU4CDJwcjdIlOZOlfJ60R3EH3NqoFM00VDOIqUIOBgZ4iKbGxImym5VwO+HnI
I5yQ46SmP6/SbGHj3FIGFyQ0GTLkTpyPptdj/ptSxkDlxAdpJTz5gcY81FwqljwnhAW7uAYDXnhi
KJ/CoPDdNRhIiIoX3VfZvDXTiIx2kwHvvzyxPlCKz89EFgm0tHq9+C1J/H5aG6FZP57oxagrILIj
ODXJ218HsoB/LuIOg+ypUoB+z4HBIhUkwAl0vG7dLVN7hrVP2dktHuld8QJoaBjSEoGvt9A+P5yh
3MK9nUphzOJWam3S8uOtlPe0HZWACUmMihBApsqG0ChD8ENLu2uknl8a187oZWnMSpuukZm3kLl1
9WjbPUO122ziwO1vjuCowhnxwYddrpD89mNR+JQrOnB7OQVbuDS4LXGWxZ9MUVEUt7TNuIWp/Vt8
spTgMT2ub+ZOMYwc1ss71OushnNLkXESiNIlU7jk5bagelLwqj1ASKpJLHdUXu228m6dk8MOkF0q
j42zS5WN0BURsM5se67HrSGpa/zqvcV+PF1oix3ns/lzYoAd6nUCWQXGorRre0Ox4Joupz2jgvBV
a0reuv70fvtExSTNJVR0SYm97TAIrK2TCtWo7A4cSPR+pl5xqdAWy/yLKC9epd9fL+RRmcllm3S4
Uygqycm1slZlwOkCStrNeOA2QCg4vpb1aj+92G/OWsyCX7eBB8e6rlIptAsxIC8L2Tld2TDdTfUV
pXRcq8T3JwYyEaNS9J3stl2BO1g+RbL5uyWWzITJpwb2UeOXNuGOkdDly5323fL3/CMLKgdqlRQB
+ajWozDzptVkV0MW54Jq/WqOYgyaryjw5JOqTEhXHmdOLInH66HU5GZr1vx2YoHnME3wPY5itEdx
6jXXZaepT80mPPEbkCdAhoFM8NPMiUklB2X0iCX2Tulhh+mPX1uOzl6a50HwVCAfcbwovxrhpP8a
UrvvSPrJeinR2EUwCAbHIAiv6VZ0uVI2tlozZhrLJy6GVYj5Wcit+rRMBS1BBWzeOgv51OnqtCnZ
8vuX/29yz4cpaTTdT+0y5zRf2sDkg0FOrTdpS5Lnb4lr/5Dpll/yN8aSHr9lXGQwuutywqs77uTd
PF6Ur6jdQw0scTRvtnHGEwk67w0RJM0L3PyKgFJ8gPPGxJvfqkT3kwdfr1MrL4cuZoBIgMjDV0Nt
r53+UQj0TaANPPztM3H9GWy5ej8Yy+i6QsM+wCcNLffCSnJTFJlqJCHGMZ4OujSI80UwQhmtUqPm
fvh7ZtGs0JkBpPQJ1LZBwvBvqbEo7YHB+NPJTHTXUCuOx/7HAnDIFqCNNna5f0UNQaiifRMuAbDT
Jm+wmiUU5ANrVGF/9RjHA4tlpKXEOfvmFiJEYvcCW4yY+owzHtrvrSnThQEShkTPGYYUYOR0qZxQ
ySLLJKg/4gRQgcYuou/oyLt3wKvOHQu7xEmZg9nLuwdfqsawu5fWbyZCVjrch6xT3fEM75yJQiXl
4Xgf/F3TXw49KxlYm8PbpNCNjLkWbeUpP6ORk90kJGkx+epIfOaK0V22/+SCVRmbySYiu83X8782
o0/m2syMb60cHcSOxNKUSAjFaRIe/d3HDRYCiDGAGH1uY9dtK4WWm1WFcJouQOTP7wXOcQw5XMXG
yDDeGNwTxKCRFBx8xzd6VMM4r35zCKNTgSth8icBwQJB46HY10lMWVoT5t8MNO/tYIv/QCL35dZM
GXBA+WExK2s6XK/iVQR57O3Z2wUoS+JqLol05IISpbpT3RuIg+Z8Q1KlVuIz9MpikszUeDEXpDC8
wLsRPaVvFfj7DKhkrICwf5qBJtB8keWf5/+4zqszCkzGpGJtTZ8f5/VKlXXPbtIyAI+JWnvoCXA4
r1A5CBq3uoIZKtl/V1JcxbwyDljynbeyJxbK9B7cLErbRPW+UaajluDMnLVxDM+0Qx7OT27e0Nmg
U5MG6jUopf/vmxU2tPIo+iPUyCTQI2z//sKCKSu4FY1JQdlOPN5kLobmJGsb2GFmlyQeles2MsAB
HiLZoNNB54/CPBe5X03/b3mMsfpqc+SNoFB2aeBhNyExtszZaEIJWSQRMiey9TWlWXrqWxcH50Wb
/+d0UIJIcaS6dmWkVRGKg2c0rsC+5Z07Ir7PFL7/qMfnUWDpIzv1gP7asogLiAsL4wdESvcAs/Dg
HEJdaZ18eHuvdVzYH1iQcS6sDCeRK28DKfOrAZxUHgHTImIVgugh/uXJTqqXs/zPJbAlL5tEq/GN
UDlzIQhnMYQgcKfg4brZvjejKrsxFTJdfIX6ZcIKipINCnLX6Ey+TWY6r1IFO6m7d4GCLhEKA+vs
m1Du7nV6HvqI/qa7695ebWQnDMqEQzeHD1zbGItS4hiaLK5852Wt6fvoIMW9+asTdDD5xZX0q4BV
ifnq9yAm2hsdknHXu/S9Oj+8IAGaAcMlFlXk/zWRIJ/SYMXPc6MlhcXYXxLnGk9lCHqOv+N96g/c
bFLtjaqMAhRTzL2OwU+qHaunzkTVC0hplatAaF3bIfhMpPoTZOtrWermZ7yfrF+P5Gx+ujDR8PQb
VjJ6dPo+mWMXQEzErhUBwesWDzaWf3ZWIXR0PyMNPjlS/zBva9YhShFsbKE8W7KNjdxrBrQsiJTN
DKUvoNLU6fHHQs/LvN0qck8swc1J8tjpvAnSpbvDsFmBUPIadywuMo1ITFeSVAUEJ1wbBqGgosue
wGc7po35/XObtscZHBUMG8BWJbfmI6G4Uu9dDPJdXlBlAnSI+ioH+w6ioB0z2Z0gzQRBUj+01x+X
NnaTinodbwkuWCwDGeR12QorRBuUJP+aUpAxnNXXtu5Lfif9dG89HmgByArm8Rr3qZB8HK8xXLGq
k6arudIy9VlEdcT77ceTKY2JDSHmAIMOkaHwTEPUx21P+o1CzHhEpWu00MlKCiedvDCtYJGMkxVz
sfS5Zs9XbHM/vEsnH8AZ0JSfoK2OCoSTh+YgFrpWgORQOVg8DRTh5lYblo18tnHmFbK2+OhB5Kzr
5Ed75zbfZH+BEIYek5/tU3QjaJewLmrJywSnfhJsdNeDCv2qdT4UtJqxlYgqlmy1Ggq+xtmv6L4i
Nk6+vJOTrTCLR5xmqUjbx4/a8TJwUv/2I7//aLVYjveF1iEbDizaRY4Pt+Y71vavl2YN7q//3/0Q
x4yonvQTitlf6xWhDxlveGPWTwUQbujWa3I6RuOeoRq37cKbXBn31VRkCTinF+cYXJUAi6gFu9P0
YnpEQXosUvoFLMKjTgdAmWQ82BlyJAfq8Uj3NvS55rRVZHLEjrfsZHdQVpnpZ2uMReMoTEuCEe0O
0S4OKArXFVHFX2GuzhB4xOLaiqiYrFhVRmFHyuwUlSjnSpl9kInfWpe126juFiaodu70mQLqQHe6
rOUvfqDXB5LG05S5ln3+olKcP074Y2sY3eUDTxiKoNuerlo4ym3XU93UZ7DpxK7HyO/fpm6EXPWN
W5mBjlEAK/+7KxRnSLvm6KpH9OVDDRTx5u3/mGI11FdEjPfRLNV2ncOBumCgs8hzTDdbExH9LCzy
RBzbb53ISGw//Ya+Sq6vSwu4oZDvq0z1i6lKe6q8tn4WrUrZkOi4lO1fBbCjRWVO8sZWO2MhE+tq
ah61+3pOuV8tl1BmO6EFgkxuShH0/BCnqpoBwTUAIkTdR7cycI03E3IMnBRbgJVydGi6QoOtwA2b
bHhhf56GuK7Fsk7wSj40AogbNDxoiXX+xAcYYHt9jwAyOxEGM//9f9HB7cQTtCqGFtX4xrPQEnHI
cygN+wz2tlifEaR7Mgv+EeiBbFetvdKDun/UpYZxlORajJPBGI9fZVwgYLmU6s0lUHxJJQXzEQkC
ToQR5UKrdtb6EdpHQxaBijDsY119iglvMMrNZi4su8BanUCvTvOaZ+LM1fnE+TsXPCqbWxGhxESt
2xOUswZWtDMbMRCTZ9xHKYAOg7FjPOOn/jZOHGTU+zKVkIemyhgwhR+9nCB8nTfNS/xTpNYBwM6u
ko0UtWLMbD1bgsXLuJg6vAKz5K8qS83pHRsOnKHOe01KSfSJDV9PoL6Hm1BQAJZMSTwJw+NLsvMW
AybA4pZMWp1pRDl6ABFRNiCKDP7mSqghpY8LTy9MFUr3lHMpgRMA51FkbOPreX/e8GG8OvBiB7G6
1cLtgZVboz/OmUNyuVCYIf2VIGjXNzO5quD0nXLSv/4CrxEjIbGFOb8UO1Tq3sTrM8x5DtYceswg
qNk1ym1XW1Romwo5eXRcGMX1cCv7svQBSWYk+V4vjH+ttxzoc3xfEkWAAknh/0z/riGo0H759KJV
3VUoXPEKOcFqY8TOLE08EOglw05WUO+vORApH8AX6rCnh530zhLFlPF7b5ettDv9yqD/Kpl63GkZ
sxrx0fV8jKcle9qPOn37QX2bkLy1oSlK50TPS0KrQxCtEmR/RzVkEdN8cvWIRgtxIqQmXBNCG2Gi
q0sy3JqiOhXx/IqwuzemDQpFXL01opZrkGyvisK1H3yEVx4RTqOidWYxdmw51zKjndzHwl/JRQx2
SCuO3EYPwa5BGwkRnGVLImRGmEMt0HA2rC3KMvLkCCTzOJVfcZrGI1MRXC73SKhFdgf61b7y7+Ct
cojYK3cWmim7EmH+yL7Pclz6T3LXzAyhRL9IBm7ZLLfD9omIHgWB3FQNTTgAkfR5nozq6uGDUgIT
mculit3sXVNv2ZET1GXEacOMwN8sAfsuTysohSBTrXqP4jFown1N2+5ljqYlXHN6aqDE+KT771dW
ewG+Au76IJb78DxElXFZ4d0mFTJoELjwnOosNIAeODksTk1HA05EUChQRZhqD+llalneG3zO86/m
Q+Mv+aVS3yJ9sOpW/sKIkltu/7BVoDKJWd7ovbngEJU7bE/wmkyzRBlRxdfrg6Wb92fYoWEgzOwr
ZCYrf9Rb4+63ywQ455HoMJPBCkaPpmptZL75olGSk9k0NZTZ7JH0Qvxv41UC28vWgJ7KoHysdr0J
O5LENDVybKrXtTohGZtEiZVpmd9WWKbVA2VLel5fkIE9e8DlVaSgrC0zNDez7T3iTqTDPjZE59CZ
GkXqcX+KP4biLaXPot07TZSOw++k2Au49VBXpK9Ha2VD3rs1fyzN+bhRoTuTSG+A8tyvqBgF2T9I
B1/H2B0PdBOuxFtz2ZQvaZNHaaCZK0DO1W0bxRZYHhgnd98FGJJi0hXmz/ef6nQKE92IwmNIEn9T
Xkn39OBEZoxl6zytumigBRlc2v2DRjupNkJeu48p2fFqyVR1I2Pez2b1MinuS0vH4TGizhXzfC7Y
rAQ9gERc1ujFH7aGLAB8V4bxAv4h6nv0dkFzB44aYfgSeV9SDzxjgQ0VapuiLA5hEocLh3JVRDJX
6htDx2I4Ob/WcJMn51rKBvR8G11s2ZsbZ90e0Z7ZkGTdWPvAA4RsHlUvXngIn94pmv93YrGxS6rq
erDd4s129Gf2gayxg8x3XZ7GXvE9obFHsF4KWHH4NDrqBZ8eJEA6ndiwy0xojXdLVmsTaczLi9WQ
RfCutcJKezgCDu5S3yueEwdrI4ZT25XOhLa404zqmcb7AWVKmEL/ncSoFqgzZlvBBeqvSXV66X2f
wi5Jc2AJBPPAl0kaBh+cifWVjLz9uTHg68sewgfRLbgNLoPrrNHKh9cxHqHFCa6+rJVEDKG3uYSI
pRSRAqpRSoIZy1Up/iIvu3FsptqyG9El6pJUaXTC/6fdPJNHSa8UnaGvLagmYa8nOJa1DrzUEhYy
XAJwavH9Ldu3ZL4Iv1lDHgTXk/CxbmupCRNFztJ1dGgjmnMFzl/zgL/3ALCWS4HLr9UACxZ7jqaz
+ifBEAZm8Upjddb2laZKYVsjgArBmz1KJVXg/RlDfnH9vIIVGadUSafNoQ62fkaqslgjwjY9IYEf
t3x167ojrhr7pVbBEeTOvYYXzpa6sVJ+k1h/vt5Qzn5/PFmWXnlGnc3sAcErkKIT0xP9l4kvzIt1
jx89+KpIHmgVnfH5kxVprKh4z4ZoM4IC8ItPxx0LGmSXQpG2oI0SyqCJSU/w2hE1+gPp18z5rQUN
atp0yzFw0GyyG6DI6BYfDrdRzt0L+HEowIQoE48G0W87MKm3Ux4AmilPJlbIs90urKR7x/kmHsX4
WcbkJbzUpQyWbL2MSNdhIdj8raU+OmNoUknqL1UJOw9fu6rLG9PnO3YJoIe4mG7+KxBfvwRe8v8+
qlj2g/kd203N14eL9mNAmen4n2cdinFjUWk5F8DqIoazOkOehM0zu4dsJuAwpGLDjledaBNX9aIL
6OAyYpf2QpZWeGov8KoZJDzjSVBrlVfzSQbVIceUmtDjlHvpwmc7C8CkZyoUjxT83yNJFI6HKPgb
uOJ66Qg2sYXsW6CR3s9gNeQ9SeryZHIj4Z6TNhSImL+YoB3H4wMCr4DIkPQc9avmoJAJK8T2GmUP
4ReRBDDI+AhR5W6iH3PWREc7kebJr8Gh3z67P9IJjXZE3xAelP4th/qyBtpJuYQ76uc92bf+YXZm
JSqpOVLuFO3wQbYSI4007QqxUMd+OL2z066aoDiU3Un8E3k/nRMSzvapoASNFh/ND6h9t7g3k1Aw
zF5wK9C1giYGhcRwxEOLhbTlCjN9fMOgxD/8DUAOivVeb5TzIlnJWLSpYfCxIgbbk+sGAOgi7jy+
0Iui4mCLT11rIyTg91F8fiy6yj5pY0rkr5/ZcYuBxNi865dU14+QJ9bNlhxbBbF8BMyA00ULfUlY
2P6wKTS+HXIdNeo/CtgOKLT3PwucKqMNQQ/0ayg13oLHtKhsrXkTVQ4OHt0vPiKJl0TIl2qkHRno
hWYrdIisxT3o683Z+jmF0upPt24UA0OnJY3lT7jM0VezS4cR6H/96EIZo921Duo9a/G/kNhMdZMv
63XEYPrJXjMaNi6xnzWa0e5nKd+kMFRCIP3Q07B+Jkk5XfPISOR0uNnjqAV7vsNPn21+2Jm7sVSJ
KBhtwNEGQ1TzkaMUvK+cA975G2qco7XnEsn/Mb8mrqINnUP9+vHKcpTScgi6uLvHh6pZW1CQS0Yw
cLUST5Z/1zHWYSgfF1NLP1hT/ALPj7K8pznahQBAVGuNqM4C7j7gjhqx6i79uV9TZwBvzxcGQzJ5
7B/IA++321k6FZ0MWh5yKj7+WrnKYRGv92ta6j0Ww/9GytCdk/4Lgl1RUBH5VRQZvSj9TtQb9rlN
Ze9cHQqdm7+uqTNYNAPB4LjXg5h2ncF35aZBcuBDm9eG25I5Mlfs+MPVVJ3LSPuSWtB/nLTGVvMw
2x7osbsDUwsm6drvexz8RGhvzriN4sm9IikfWltltSR/0JzyoMV8tE4eTw+MmhLo0bdbTeJuaeJB
l1n6xX1ivM7tC+wZDHcceyWCPjwYxWE4RT6u6zr/GOLw/wJR2UzIan2w73Ngs1JdIsIccCeOk3qr
vU/acvVq/UHZQ8X6VX9cVlqxYABNQiAjM7lKNImjAwn9JgCzapbxDH+4eZUfkbeyMdnwitEOVlCK
Fq8ZdQfOVWYpTL7spJsaXjNkRUUenvI1tMy36F5AmBfET7iHAdv5V4CNA2dSnFInXzZ7UwhV9LHV
O1wpOBu+jaVN5jUhxmqwjplImpx+NeMnSSbgN0UxhjGYpVbWV8w0lloE2EmNW3Q74zYkd0UebytD
Gexw1jQguqNipZ0Oby1CLH+7vZ4pH88mbb6GjKQjAHTnOtpjOfSL/7gl4OBK+YsJrJ0xoJHhjoPJ
McdtEN5vsuNrlLCsXXbV6xexj6lncw7nPzDRYPz8SSnCCCu2D0PnpLlJzW2S6+UoOQsL3fyzgbmC
m8URhq/i6euxblzSDKRtsrhzLiTrKg8BZ0uNPw3s0hhuSVdlsZs4vjqSreKzqgUDo+gj9bPWD/ee
3Y50uRTEwwcKqltvlxZSY/JEyZ1veF0xsOr6L4ABtlEKatidWQZ7hn91uFnr0CfYAnz8mc3n41+d
CBhDg1RVYU6rCvxBdVdEos7w9hxf4b8xi07IIdOlKW7TX0FQpk4Ha5RnzT51m6kpeoxLIIEHUU8g
+JR0xArhz665OxGq1LBmjKXoqF9P9Mrjy0tZgWXfBdfdfjg049IsKEl2nTrygZRbETwgLgPEltoP
9FH3XOvN4XFZlmEr/wJvhf4n+K5ptUqvaTa4zsCOjlafp6KPOzeJo26ZF436n9Ir2bHiPlPU59h4
0knxcl1r+dlKWV9Dzne0Dw90N31olm5LMRjEpAxMKPwQBfAvDK+wdbpoX+IoZPvIAyyPEIlq2aes
Z9VzXmmTjDDTkV9Vm4KRyk+kJTMPA1S/9ueHhWq+Vc/1cuT221SC6t30pHRfbrRs7oXAyfXs8gzf
s3j/AlVT0j7bmNomdVcsHCVoI4LIW+VKmdDOrEpVKswJ8v9TuggOcxzSt2PNvbmXLbrQdvRhm698
HF5ta1Qm5wxIBzrnEvrsfYKMGELbs+fEm86ug4hCzP014serxptfmKQHOjOmrGN13Fk/jeeGv8wK
Fni05D8nKfT5RWWyLIBYSUPg/ZHucRZ+Q+ysIV/7KeMwF1QKz3ePHS0RvKIGjEcoQRPKAKjOiygQ
nzlN9vnicXJG4kasGWLsWtA3X+N5OhSUA5o55B8xO6khlbwZUmRqGWOMi/JGWL8cqCAbW3z8TtYZ
QA3+YIiGfeS6BIIZyOL1ZTHJHvZ8UVJLpgYpYjdoXJuBxL1AuTpkPFHfAcDZ0mzow4SP0yf1czDq
SdM3INoAMpkr+Og4C8LyobkQgu0/F0yhxc+HEKsJ4vTxsr7wUfl6O1GdFobEhZP0tyvAYsArkf/+
hVkyx2YvkuaoJfvKG4HeJqzGkPNv5IVpep/gMfuofxsOnCg+AQ81Qhg6MQLyzWkxhJZK0IdP567v
SRciUyXmlij0B4O4MY/EM36bo3eLO0UxleXKKoS3AqSf4lYjrHYrbSWIt0JsXfh+cDrUHF8izfls
Ob7xVSmZy9vKAZ1nORcs9Dk4rxPJLh7eOOYk94nZcDadUrWIsT5zRUzh7fHOHQOfCjdm3I2F+UTd
/OEZroNEtmgKdRZsIhMWuf5W8TNt0dO/U+9j4UPVMJ3LXkFLE1ZbgoZxLvYlSrvMQfF/zZNjw++6
0xI2c0/VHhn/ghiKgCwqTQhx9+Ebkhq3CzhYLVj5osl8bGeqUMUP/y2Jj+UMBiRib5wUmXRjiA91
55aI47dfOI9ZeiOqOpGWga0sX39567T2E/JWJWi/ATr3WxfaqphCj1qmRXnZllH9XwSLQWqTI6CS
1vPV+e2uhxofqqgLwad8Kh7HBEHhSZqKqKG8kYMHpWJL44dXK7ahW72pZsbi9Y8xT5aiQbB8TDgw
QtVz0dZwn+y2bk/FBLWu7A1A3k/90V36grDa8cp9Hn+NHauDZftpGJA4kVgwWfp3V2dqeL4/XV9d
px2feVGnNlStfMVQbMfAPH7g5FNA9nnRJ0Ry5NdLRJ3mgHD3i5lnY+ciSqlogKUj2RmCDGquV9U3
yxjIjp7VFhM74seNN4ZIKGcMOhY/vFWhiEv6ktjOcLHR0ONVSfmSbcquwwYJmLA+4cESdY3Z9Ieb
Ty5HcdHRtRSMuHx+lHOgTmRS+JM0NLPTw+ggG/1JGBEzHfjdSA4fvWqvG7K+mEae3ZgullJahKon
hZmEC1J+F6noFeIVDl8G63/Vctp+ug+hyNwCSVvkSFQw2DC+vGICeUuKlCOc3PFJnQX4A/XDNB/N
hcys0WIQU4r4Eeu/I2uxOKS1ZMXi+Z2r8uNLXfSfvWXKOwAQygVJEHWT01umTqjWIUFOuTKYygtt
Q8kFmpSkL97fVQShB+QqcMBBb+15nrcIH5m/M9q8RQBSNDCDB6c/KflCCzuwn+Ze4UKIKlL6u9ly
3+rCVHzNW/R1xEjYYztX4URI+odmFMmRSeLeNrd04FnN5tv8P980LKhypyhDO+CCPtV8Ued9Cz3Z
+RYf1BeSI+5LkEfTAga9Iqe94Cd/kS+aOjk+gKBfG5JSrUUjPK0Fqv8f+2Kwq52IaFW57/mhaa7R
IBxUETcFY2L4FDTLfEvM7jeMa5+6ox6sbOix4HJB+VbsR3iBWb9piSsPq73wErwxedsgWG9psY3e
qBHhsczHNfUeQfBvFrHPzexsTfDTf5A6Ph4xcirbgCKSbBLpVBczSmY3FSJjsAlyTRE4sfVXOMD3
jmGAk5NSEON0/mOuQjJNMMLNm6Iv+VcMJUpQRYKTBoZJTKMFyIcieTkgarAAV9cTSgrjIWd0UO0c
0Yhykfkvb/IwnUQlYqGFj3FmBXkyZTOtJp3ADzUh3vUB9/JZbVd76cLSyM45qygR4NTsXOHWiEFP
v+DTrhlMY+5M4Jyjn4159FzPAsdjL7zzfWdrEh0nrBOn9WIN06sAJFdkixyvNsalHgWohL4dpUtr
6VEMxPBjlsWv+iblQTTWFAt9v1UumQsUjliwl/FJjGsLZbu73pFzqf8HzDatH9YfAjtrIZA2OgAk
qoOYP7/i9Hs89vvhokdWar/v7Jbgi6HRvsTuNCNYG6esauz6PZFS2Amfo8fHjXzx6H+oBgMH/1PF
Soyc5EPouNIdwWtd3b1vWefiG+AwjA2aRvQAN0C0tgD8kVP4lorDQEy7P/z7p2Td6MkA085/WT5G
6JJT0XVTXFXQZj0oI1uCj9+U5P+HYN7m0/UCJ0iLXEZdk13n87W3w6VktC+dhGLZIj77/GUeAwWu
ykn/vGP0ld/peg0rRK9QCx71JygOzbFNCmHp0h+JJ21qiBjtYm08hNEevkTkABAA6MV7cT4wErc2
3oGWCw6qRBOmSgn5UZlL8wH9KRTA3EXypm1MfEhmcgC8dnCvbBknNniro3onFOMlcLD0FZeq0TMc
dZq1KJtJv6fgkq3I3/txyqkE407c8FKbC3qk2mWRxoJ5GrpIpbU5ZiOxm8O0KTb5tQVYR+EFdluy
+2EPU2dSXV7nwe1NQxUrsnqn0zWGbJrP1IyW/6dwGUln6Qlza5ce/u7myJ/1CYC/LBSJ4EwjW1uc
P+4Bm+u8c7wVQLNFHAB+MQlqI3kPGxs+78d9pGVABS73y3tlSyWIJMTfmxwcvbQuvXn2BF1BNaeR
o5DHEFlPV4uYWhuf08bampX8JaaxlrUqf3iI3rTHYRDwrn9Ea4DCzpZUvaguMMsZDB6MG+34Ql7J
Nl/sKXCLloPF/rPMiIMP2QjNS+09TNRZc2UAvxJ8rx/kQbB/cfxKZ26XYGLKsGpCyRGNtv3S64s0
NKdaKsRo9iAhvYNst5/9hAJmw+2Vi9GnHO6CZOxWeXxpKSR+fWwokcfSmgPtT1z5+donA3P6bgFs
7aMfTgLoh1QwIYVikVwgPgFuiTkX5OBz0BiOGA1hhTcgxqPDpa5bEkLPKWbunjuUEaWj5DLRTsii
GvZKwzZKLWH31SmUTwVA71KnnlC7u4QExIq5Uw9jpFt6vj0DVWb8LyVmyyoAe27CgyM2+hi5EPWk
xjZMD399PRwdz1pAeRjrnhJZWKDMnFKGH45l6NDdi2TcYxFdOEnvnMgG5Z0HOiq5HQgbDdOqn1w1
RpLazZRhuH1bXa6TpfluB98a//DHT/j6ZH8OEtPJ+hkppIMGCvmaVTt8z9DnN1/bQyj2sXDGsEaQ
zt52I+ecSd+1eFG17t0gxVbB4/IZuINRtWVBbLpKsh1oiARpERc2+AO+Ltj5Awu1xkF4KaVfIj6t
bmpbR2bT77Enlf3Thtk+Aed5bjw+55iGrEvRIq2nPTbPdDkAMV30yW8Bd3inyFw7ZzQf3qr6YyKQ
MAg5XkUEkjAU/4ynxN6DMM253QmE42hyw3+Jji2FZw+8hQ6NipWWN2+lbSBg94CqozaZkGQLhfX+
YncPZrWL9J4Ccv8zcDSOJbz5KgKyZtlfzXHm+kKcLUwcjUbkiw4kXkeGhLrrDXqcmynJ5LCd9oV+
s3wexpVEbQ6yLSo0awZPRDqMSrHCUJA4HKiE4ZWEkYPzUjQShjhymsZiDUufWkaMOksrmMQjhs3Y
4Oz4G8fkmusOazBzsp927IgAsUIPCMe5OosnnSmgmaiQZD4gabpYFSOgx9k9TYr1IEOqKix+YbCJ
EsrhVDy0nhiveLmls7INuYmqpxTTDiLatvkfAszzMXN7Vazx3M5ikqoMYmA4QnIZeK0aE00+SQk3
GAooS2byKmprFpBaPqQy5aXXhhH5/nk4ZtQqtjzLEivarh0a8eiK9O50L91OixLqA+THotrnMc91
ZkgcfuedxVhVYFsZQp4MEUbNangFB/cfCI0+lAx0t2Z/i3zyjDzEVmPTeVzGdkKoHSJ6woMPtBf9
tUDwvKXjxDsKZA0fom7bkzJN5jBBwkI48PSWCdLpX8SijzFeKIuh/oruqR3oCXyuKEj0QSp773VC
M+RId9OmLDqs54bvU9hhfSljJGzqoR6qSOBaaU7HjaUsvdMQtHKpFyqO2XD7vS1yz5/wC+9u6DzW
+yc9vA7GtnW25AFLLjDQ11b6q4ez49qPGLUFCxB0oqCD0LgsMMKPowmtKs5kcVM0DE0uVF+C4hI9
JpI4df0rsPI9EdHms2dCXBHRs8hPOMDoOYrt5sg7ZxiejVHVtTr41x+m+nb12llObB8qNyUPzsz+
kfyO7qhl+MBFYTB0ULz7ysLqeGL05s5iwLCPH/zdPMy2O9rWDzjXX/XSF4zJdEOrgl+t6INsXVcx
YPtPjyZHsqD+BOZvisCvxJkMJ9L/2PjV26PODdzg4uAy1RtUamPpzQRTSJhOrcmXN6ln3ICYY5K0
VflxCHhQg2wHgNagyNjy2JV9ZjJnx6x/yc2YSNC/ddYztF1WD1OlUe/9KSoy6uAxyX5QQb8tDJLz
vuPdoVH+862aePnaxfQr9VG5GLMIcgHpS5WmXr/R7PY+CTBt9okTAsPdStasubPWEfoGL9rgT6um
Ux9HoXDFxxZu/bi0pMLVr3s8spffGey7qxeIeQczXNKgS3mqRDWUOIl8hdk1Mfu+6Rn/kcAGfR9a
KHlI1jtkegteP+PYKeKq3RAFUQcOkUMU5hnfM6ITiZ9iafE2n/1vJqPGWQTKQ3oMjomxAAOExE5R
vXrU5Cw2KBqCbx04/dZbvPUCKbhBBMlJfdba1ZFL1RwJnRQPlnP7Qy9LMFs0OwpT66Ok9hS1quPz
oBGPaXX6XEGzxlJMzHi1YR7DA+mRNhqM6dwjM2vVnrnaU9UL2WINih67abuOQxYP54c79iCpkWIY
wfJSnMkzvZLNVH8BPOUQjTBw85He1AqmqjcTJeBx/Y722wjSceU+vlnbKp7sntWnuONmsKxr7FzJ
cqeV25L83MyjRA1C0SIPU/e8fxMFrjt9Igxs20pqs7Ge50WiV5iwokULiC06R+miU7LYqJkmX628
srh4j25bWDZ71x0YN+8psVKBMTI6FOiJgzvTglrqRlLl4Fl5NUUzHgYqmdrSmBTM5K8/K0Yb9T4M
VtUNOOJlTsJLefV9bgKCo/LQPUuKh8XjdxOyoDJFQjA/hnogO0CYfOXT82QVbbcTaH3x1Mlz50Kj
KZhZnzLbQCUa3gf83VtkN03pj8J5w+3CyY2ACQxOl7dnNYVj7SDsmxsp7+3zGuCV4UUVGJAHV1Wp
NkEofNPNqQkFBYBdc9VtXwNf/uRc5tBpeAWwZlQty3FXkscurr1r97u/ddOM1r6wxc/1QmI0Jm9c
hJpbGpdqZqt/F8nktYx1ZrSshqvaizNWRDBvpuLCKX+b9QczVavK+I31Lnjcu9cJbWGQLBbeeD/C
t2wr9V8KOEK8FIU5yhLQa6CSdVbOk0QnxJ95BCOcQ33y2brIPnKq91d4H2REV0VjpHlMatcu9ziO
jaQAmlEGhoRUzStTAZcY8oW5IAn5gMjPdrUowfSCPrMT4PHeTgrvJohDYruwuOE01h76L74mhbBo
0MutDg2KqgSQNG0owy74+9mQo7psDQMioskdpA6Ek/3eaOd9Ic6g9S56uWAnPbeLFkHa8e0bp2y4
DoCfIS+vt2ga0+UtwiVwmz9tDkGwOfMt42Doan/aujwRroMu/dvMrqfoCfgFvYK1+dvjhNejCaXC
bQegtKMxz3mvjeaYrOPIvW6yqnwwG9PL/G2xWCIn4kTyOleEKYIJDE0T+dDNJlGa5CIuqx6ABVRQ
uXw5EAbBLrA2EaoDU6AS0oUBkbz35Nmx5qr60mskGOm8tNC4jxSX6EjoifxNIsSQg8e4lPUnbQYv
RwKZs8GorzGHkLMwWirblZLzLmzHKoy3Kem72LINFI5J77Fs+FO/tw6VXVj1lEqzxaNBLH1x+NpR
A49mbkR1eETaBx13ucwN57MKPWs8c9OEE11TwKxZS7CRWELSj0BN1PKbdwZ8ztWsfd+BIApPEDjC
kryt5CsXabrQSO8Nyzq1CY73XJPEuf1blalwsc7t3gCZnh5qZdOstK7SxcYt61Vh+bPIz0XavANV
6Eacq3QzKh09P95Wr7xETnHE4HdAohGQZk0ynXQ4P8220uIWRTOosm7O9hCWIFZ/mbXN5W66p7xe
hmDzn9kb0rA13DE3ZP7Rzp1QmnvUAQLymqWyEE+uI3XUUAeQ34zYTx7DoFT8Ey/UE5HZg+aJlWJ0
tw6B2WmFqxLgIjZ26Cwvt3tlBKrnEzCuH0zVpPxPO4dvvlTGjcx1Nr7Iy0DyU/+HG2lchSW5LGKX
gIvFCqNswsSA5O6xb212QGu3hG9YBBqkBhVBz1wYgFUFA/CF7gIqYmZM4Kn/lxbXGJDlJOkZdmzd
154m1gIwRPC6ckMXY4gSrYXS3+EQkHT6knvLl3uQ2jN4P7SVqSdwHvxRMSI4K6PnfLAczn+z8j/2
8LYsv2Xxyh/NKf/96G9lJsa3wsDUJBk6CWva+ZiEsUJC0lZOZ8ZljjsoQ1B2olRUZiuv7TvZJ7o6
7IG1DO2P4lAezX11LG+2GPm/2lShwi1QUT59r6d/dUb4ZmllOOzS2mgmhHq7tHVQWut1umStXZpz
6j65tDmR4ZiSF/2abZjtaWgL1TSuWPt3potayzyv2BcnObAd7EUkQFHzvBlIY8LPYltM10xbmg5w
6PgH8dSyvSh1QnDYMtgzgyOR6TYfX/LL9smCximwZJjfLyDWdknGGMMkEUCkxYZCJCjdQPfkZiP2
0qG8EcGnDNqG/DvioK8+yNjbtKDbIVTpg8xaEI5gC4NyexGJ+9j1M2AZ39NRIwXs3s+KTMjCci5M
hVdRNwODwJRtziaIE/ETG7cCfjtflw6E/uJp5zU6XpMVRvvt59k03FpNo0rjxYVHy5O5Hd5i2a57
yJVSuCjvJuNM1kumoONJ9F/vfsEi8bpWfwfWHk+wi9+MdwUqp//mcDBEJH8beqYTgyIECjIUCJ74
lX6O82X45ui4BIESBuokhsiEjCU3u229ywcrk71y8FMrbaYV6kZnBny9yS+XBI6/BsHcUSSDrxCO
hRsRJ60rzad9xjGcu7fxyTuYRkitRXV53h5ExDCoVTRgpUNVfmmf3ddjlC3OYjf+K2w9uz6RRdj9
9PWRF38ZxZI/BwMf9hJQ0ukDbKtKaAhBHS3naZSpXL+s72UvxwIZPLS46ajfr9KBTJ+oIdZSHB9D
8G+mFIQsgO6RYFaYLQsNl+EQq5DiaJatO0CBunx1W5BLlx3Q117K6k0bn3/PKx6vtXVIGHPYxEki
CzD/LgSJOMHAI9e8pJ9srYyHEo7A4n1SAt1d5CJ1Fbah2R4qnu+XWLacRauI97MJFYamCG8VsdXL
zrxsGTaThzuQzOuMUgfW8IvilWuUEin91dthAJtSd5QAckJA9ppvyiVW8Rl0ARotvt5s0oY870Sw
LE+jnZ+qoy/TWjc/EIA60Ca3oqjluNNu83CMPVo4/No6Yd1OILEhDew5tIfHyVMIpmc5YyLqZFyg
E9uDBoCWTf2jDJryVvI4WIiXbD9tsL2gZcUw1MfANAbYmtClwf3tQxIOQz20DkWZFtMMGiFGOhfL
UUgPV2P2p3LKT54hkotRvjevThyOlQDVuk0YkfLIitVu5yjORczqc5nlCIz6Siv4IAizJeThSaoM
hWqEPJJ45+jzUs4p+3hHj2EwyBpQdKBtYzGLkX+zN16es9Kr7BmJIWXY1A+5OO+lbtG+BsydD7Rr
yPSggUIDm4GvSO/TAnvWgp1b0ImSruLqLfYFxBKyo8Dzg4BTO+4Vr1iX3EDe8uytkU/r7M8pUikd
baopRn/cbMY0e6l1RbNQnAdAhbSTQHsh/wAPtmP4JsTgSHcNkw+mWQzbJUnB968kSyCeVfWXrL6R
Uf2Hw4iw0dd0tk+MBr3ck5HhctnVdC8/W3uHgWnVsTV7bWHNO14aKYt30hQAEBvpFDey8SIicpn9
7IsXngqdvZuFR7JeJz0n+6W1z3h/KXY1cWHWFiAT4/XIezfjq5KE09gilDxti1GGRcbaonqwjdxt
amfVYOsyslKUVO8zPHs/f6BoL9FadqWZjO9vrSH7NUxmWDf/vtAD9UZKNpVY65g1oAyc+27aOpmh
jexF5WRkza7FvXTlWfwFwZNdN3pCHYGF2XHLbqxbmyAVg/J+01x1rt8Lv4YISoLq5luPmT+ngnoE
qie97QSMpx4orpF2+hV7GPARrCsKStfrVOKKmfb+7jp/mZ4/x0bPYIW3+q5oXb7Qrl39zqCSxM8W
DUW+poZ47ITofEEdyF7uwczW4poHCFcOSYCN71yo525i1ulfNrMKDpOZlDY6O+YBZCiyjE2StaHd
z0RsnEAkCV1IYhm6ed3ARmKOcDxe2E3I1JEj7XQsBjRJEFSMn2m5NW32fB5JtGy/Aqy91MAVqAzt
b+RxaUrqfJzZ+cyvCKxBP1k8Zt9WmZp51IMykyep7PLOCfjBx+wmZWgE/SDYoU3TSrWdgbhBXvTd
DxB3L2KXJDmzxPLmuPiHJLtBW/Pd3xooJ+bmi5xqXpZOblHGPO0bmUtga1svsG+0uylmMnBbRM52
KX1Yj47Q6jkWWJlOR4Ji2YcsHEicFKlyKWCe7a+xnJhl7hR2dVduqQOOUnnLT6VhkWcZGQMOMVNW
WmTLtb3L0mLV/vnl+JZHNnHt0C6CY4zm/adWUYC86qjl3e0jxyRYwHH9LR7QTdB4z9y8Bpe7Xx3Z
5mkkRZvlBwh1jDAOV2J6ZufQrt7G91cxbMOP9m9FDHFAdDoAsm79LnZne6MpJLs/cgMnWd4hSteB
NyWadCilD0LE7D0cfkBwd6QbYsmB8QIjg4n3KrFcrjSoKEUpRxrKMJmKlGKYuBytxM3RIw+fKdzX
tK7lb7Uw2Xeto9XXZaoKx6coS6wyXpZlKv2PlibWPMU3kNWI6juNJ+yMHAs89fU2zWKjX+E88ka+
7VfpYYaTbgFR6Nn0PUB6fi+5To43ZvP76hf8A0vopiTkxEy9HSYcwTZr4nqnBcU/c2AN5gMJgZwa
xrRiwctFgvu/fB5vsZA3vKRGCQTa4CrnrUKuFnzKNhhocTN9JBwmyz3Jnz89eER/n8HwoxyN6h6Y
HGrFMRprEVDGBy6rJKAZ0Digqiy8ZAnnxxu2hB6bC+bqGnqlsPIe28H5pTZjf+93CChg115uSPCX
WsxSyAkMVYHdWjlDhWQU5ArenFLRO/Y/KS49nSWemzDaWgDn+w61DzdwAXTPQJal2O2R4+ziFizv
1NKruO3pQU+TjAo6GaruS2NkDhyNEoq+mQJfzq++4ZeVnIBH0g8UZR3ccewtZPSEiFurex0CVSQo
sNj3mgLmicVglLgZVqOXjVDwhlKO8q0LS9jsNXgRQCLKP7Q0c+zmts4sLEtW48bjJK9MGNEmsbaF
mv0Um/Qz4y8YFKDD1cBBsIZn8uthYiO2eInLJ17lwpiy3hCZOYfCBIwFpVHIJFOs5yRdXnGYuszX
rl3/sZUJ4gFU5C30o2nRkzlvhYXpH+X/su7zl9pxpRdXWyza6zinMNWvpAEEjub1iJi6ZAznEOFl
BzHMm5uwEbtmwyo3tDaqigz4DlJe0RASly9TBG5csY7lsfziEtSjqeu4LDIQ8K4Qk1ncprSMREIF
M9KKgWfubhXUd8GSIStoVJv0YH2pTjFJipmLoMbUbg+4atrpivViNSdJGTyd9zDDftolLk+EBeUH
uwDfKrw/DWSKgM27/S/32FmMwN0lF7hMZwdCFLllTtqu+zMnR6NhdevC8eDgZ16MLI1R7VWe0tQ8
xYQ0F5Hx75Ly6+AGrODp+PS8kYzE1bk0WYZT051snEj5mahvOcPtuX1NokRz06ICvpfyIfh4yIS9
rO4LU/pmJWHcfzZ5VE3OqEjdt7kcHNbOgiw8thUTK/no+4/4+zjWXeratIUpLbTnxcXBWMpUs23R
1qFRweBrqSQN5xIa4q6vfnU90Wodqq3K3OEAjz3wOQEd6USHIzhY9k0NZ5z9OEQwgMf+pE18NtvT
gRhaKvuG58YZjEj9clqP4aEsT4adhfsjgHwekmcuEB+ccWp7amQKTIbwDlbvMTpZtizyIUKWsz/T
gbmXjdOpxinpuUU87P4QiJxXeiBdljfySLpz3P5Oy9m1qRLjskCuAsI+Lp5yIb19qMRcPGuxmXQw
TuKX20caM5Hio9xpXoW9Hsbn2tco1M2RqcBmMpncmWmqHP7XeTXca2b1uXLIDh78OS1sUItbaMB3
6LEwNbrStzWpgNDtwSl+Ke5aFZMKbLIDw8Sat1qJn/XG662Uc2QLR9600OTWEHDJ/ltkUR9CJM7G
Vy/d0fofK/p5wazfD0ZfcyE1FBp0jGBGqNJijRLFq5R4ok/5VQ8vvUHUig1cZnrVgDaDQpgYEJSd
0T1F3+ECZNjb304cjM2Lk0cjTGuB8E5W2EekIcAdEhRfHYZY2/W+mHXd323+xT6PVNkDjPcOrLQc
G3LyqHgu6nRygiEsz0NlDdYz14DyV59BkUsCcDPCSLPxJ1jlz6arsg2W2qchIrh/CBTQC2mSMoxz
3BlziVerRaH8Or6M0Mv5Ap8OQlsb0r1W1IV8aykj713SRhAMXU7NvKimnpr+GqHaToGTWTZH+PfA
WyEY9Ovd71jpCrFIjxhHFk/eSs44zx5Yt8rnoV5VPHOa6mD5u7J6HxeebIoNlwL8lkXTxgCLA0kU
9eK4sF1hVZ5ve+3MwuWf+oSZEAau18DFv/tnm8mhO9NKGe2ijGkf1Nf58gNCO1bxOJrXrOAdasGQ
UjXssQsdBKITX82+gsYz2cL5yz4ZvjYez8l0zdU4ad1Xej57o4fIiQ0RQwOaPEzNcY/vLAbtArZ1
KdAkk1f42pNbWnkWp+OSsSKR0JF1rdHVnrwyinQeYsz8uuLyGTniXieKJO3O2UMoS4Ou66jMuMun
Wdw/gZnQ+U4xGWOuvmbwn+Nmuzqy81NuyKdLl1CtwRKK2mDqv1Ae4lhyE5MtLqyvheM/Gl3KYBaI
nyF1PRkKxR2xF1TLs1NF4mpEDxAKRk54GkBuu8peTf2sWkzVTKJEMnm++5WFLkKwVe63xq0jsqUP
S0hOAlA5kIhpEQNRce/Xp7xgzFHmx5DZnCbUckyfzDByJNAJ+EK3Vfljg0GDqw/z8eoTdBa1F9X7
1acdggtg3rYWQ6KaJISLre0A0jui0nppjPG0WV0kZh0E+Xlosz9HhKq8kxSr7wIAsn5Na34FItdy
/eBqRUwvJNx75tWoqf9Os/jcGuVhgzpebTCzVphOhm9h219S/9ahV4QxjkK6z/SFif/hjUa3LuCv
w/r16EmpPSUF4b4wRsLBXNvn2FO8zAiaUW8uCGR7H/MqObQhFglfEZK5GY1AhISobAAKHNwdO6r5
vuwgDqtI/G/i+XnKQrcsvtD+3zAjewVdOWacAoPUtc7LNlupJbkHpd5YaW7MVkaw5O3+qVgApiUW
r/AkvvXVrRPBDh4bMYhKXnS9ILwAEOwELcCS/NxWwHt7JqVvZW0GW+q3Kzu2pQ08c3KQOWdzujq8
gwDvCYlAl+swSSfBVH6KgaBezsS4APahWB8jFAZoUNlLeTMd244vfD7oIsZWirO2IyBg9QSBg9A8
5kcw2FEEXlM6bL07GTCZz+eGqQNbMm998d1AFWpC2rAnEQPAblCe2mcCQG1/OvbU/Z1y0k8qqdUv
VhDPjHqYg/uTypAxfOs6i0Gu9YegInupmI1Axo4E1/9i5Yq3UdsAK8ieD6enjhLaRmTeMZBxNmaK
824D7k8NWkZ7mXMhyaotiGB5jSjeVAj/fGT5kOHFLVx7saJb6oragYqpuJF6oQDOn4FrZO9Vmz77
dde4umGFnG4AZk9ROdUwX9qxNyljmnJpshfov1RMrfmzLs8CLRENrzIdU24ar7mP+KclRm8s3Thl
87BQQoXfXSXma8UVQeqvfu6m1lWkTcMZ6Ort9BG1KsgFpEA1Kdjm6HQF3BW00Hj5oKEqMRwn+GCp
JHJbBs0USLGayoQVvtdb0ZqP6DxHBIOtw2mLHoOvbSQGW5Vu6ENCLNgJVadiEOJeVd7+Ywqp1lGd
nGPbTe4J0vRu8vu+qrNXvEoJIvC7BSe5BORKjPoL0IcpfId54+tWWp/Hw5gedjV4NqbQPOm1L0C4
gruHBrDS1lp9VFikbfbn+fBUwd+DXDMoIzDHPYZVZM0eW7Wbjosr/7yMeS3anrxq+WJNdqI7LMr8
GE+k5Eiim8GhTZkyChmrCYjPSe61NJoYYWR6pCuBhcSwlW3KBdtgdyvQVocVeQCxUmfJtrcGSnKU
VG/w3u/aO7+6tA8uli4eHdKRAt4hl5XJLLnNaOqeNGyKb811Iqi1sMlytyZqfhfDygaE0uv7NGq1
QAkkclcZOYhHUIL3mzI+jItjK7dJUJAauPlIZj3FbWc4e3n8yVvySg8tYuhkrHf3Q46avk9PTBsV
pLIeFzSHdfzqwUaDc1iV+QOCi8Mizd7uFgC6C5jc9CIIjHlvQiA01HWMBpFL/eMSCitIfy4GchOT
j6Bd4dMRRSVb5eI7Tb6YoRiSMqWNXEWWk1jaBm1v1WRXvj3IML2R55hpVLKQeU9D5m07hyLKOCuT
Tp7hWKBq34jZgRJV6UkpRWQDk1RwI4UkO74UALKCc40X94z6lLClWDKuWOTbgf7ak1F2k13UXfV3
zAPW9O13U+b17KrcOo6xzW3S8S5xyhNAmXWcsERL8PDd5j82v+6wcra61jZY7DJFPKK0fVgwX8b2
eTBkY/UJpf1PAavmL7IUTuW4hgkxnojjCOw2lIPCoflCuHzUuXAz/bVH9gS5SHxAUa++rNpiSDPG
3ydkIjAcfqNgRWiKqp+On7CNNeblBwLCARDxTrv53w7kImdmUxBPIVVkHRGXJgJ956cmH70KSJyL
WfLYPYlY8Qe9KprLRiLtwnqW6dnlSq9YpFi5q8UeL4Ph+J0nTNwdW+dBlq7tr/DJReOMQJtzaplH
srpSeGsJjpgepWECzHi37AvJT0c+RiWqbS/Bw3cR9N+TugiNNMnvIUjCNPedlrSucczdEtkanuzp
isuZTioMil10o4jbdAeZJeI1pDT91sXrEAHFoCAp33M1eROS/0Kv7cwy5hCZxJqTyi7z/a/RIZAo
Wo9fh6Sn4GDSftKOGml/y6iLyLPtDRst9C8H/+AVgo0uo3opk9XAAN1MDsGHLRxDYiG4SNFbecUD
QpEhoYJaUYqsdprCc8YHpUfHsrURFAcAJu2LzxpHqYTiWCSPMtV/qb3P82dGw/3/L0tSaOnXrIuV
3moEkDk2nh3M2f3uXH+3UAOmac4/klYabOc95T3DVX4CkdWBH1THtjD1uojrjyDiLS3qSIJ5pD8z
6q4UQfknCCXCJhWSp+MThFHX0VnbuqhGCoEfYbFFpOZbhEC3x+hF6pAxbFbZ+xfP0NhiiUX4keqS
49D/M90ij2OamGYgd3/e2AvJJTH1VdHO6//Js33OomckGKlil2i5joFWd345IyDC38IWQYy2N8W7
NRVrJaQA5dhaLI7PVsr2ddgl8mvF3lk97NaGeuiAppxwGZLI1Hq2zBVNNuH6+/DXVqmfEyHalX6U
hZejBPP+pZ6TtvR2Iunpeq2Reuq5h385FefiX/fLd5MttJTH8uIH/l3r0S0tWiVIePdmbQafFYB2
f7BBaj4X/0BtqvAkR3Imp2QsveHut/0JsmMOCanhbprXl1uXuh4w4n5tzH9REApSW+Agbg089sIW
9copdNp3D8E7n08zQc7HE2TcInSjNSKXQWn+dI6QJ+W1xUu/XD+4/qh8M04OTB+uBmEc5e4Qu48x
JYtD65Rxpwu413L2RB3c51A0s01dlcjHCl/A2lberAW67FsjAo+pLu4Nz5Bg9OXXNu1prO8ZrZUT
CEppupivHbIGlvzAkz/Pj8sWHtUTVpXbATP0KMwjkGT/MDzJFX6atNVuiJDpItJQe8BBDEnpTwn7
uvvnxBBvQyhpI7DtOQ5Pbf0Pbz4qPPC2oGGChRLjTOYkQxHT17BI/W0625x1iSEIxnNrBwwoPm+n
U25QCL5RhTC+OIRhv1Ac5qx9Viibf2ENfP3nRB7b2VdQuIcwMzVepDyC7HGaFWyU90f1oAy3wZX/
oobBv/4svS4LUlDii7AeXdJM4W3qqQrva+O9QnLFQYQjmiWdxiQwZuYEl3kZU8jisFgOfP9qauMQ
Gsy13eaMLVo+3JunnLyApiPhO0yysP7P9+7SeGMf8/cWTPWdUgbvc8kkImT2Gh94LO8ac4Sno9ps
UTrfYPUXrBUKpRKswR6yGwrhs2XlfFoR/j0xnjtIMzwMIxJ9aCJ7OWPvYVYIU1KPktr/7AlTHXDY
qNPzgbPofLHaKIoGhP4ZYZ0NMeVZufKE2Yn0aRAA+sb4NkWXV0BdG3Ae4O2cMryuqMRClJzTkgEV
dzueiHS+WQAA/hGiQRx/JpVAuK+SDp/Bxqwds90PuJA+81k5fr78MQHQtCwr7w6EW4lhr2pJQy+l
WlTUHzAaRkV1hAV1Ehyo/eXXL4a/+DbytzYBUAaFwL3IWD7f7RKdeKcdaT+Jn7s03v0RIZRV0+Vv
bCocahgHU7eZIqLf3SpJ1hrKNXh4RwGViiwCdk0wZW0e+6dkqXRCMQV1wIkDHwxj2vnFKgtlrJHw
5g8PlX5uRQDna0AMZAwetAZmoWEYUt9x07oVC5HZnY20WzCTg06UVePldGV1+kkkXQ1zR9cndP7B
5pmdItol/7QS9Ff1Q100OI3WGGYOhUjr4VT6aNPaMK6IIGlcqp7wI+OMR0GYbd/G2YAyTpUNZVWl
3zE3a1J2zinPMgxzHK8iZ9agd3ngeeF77QahC0S3bOrNeDdsnZ/nzEOPchUxfAS69+4pgdZyRif4
wlZGjHY8gXUMTmHuspd6VTCw/+kleQxvAcx5hL69f91PlK0PwJSLY2mh66PZraV0vG5GDwaOUuEr
AdwKCL9VLsOF1vr+yKdz5toIEW7BBzTfWdhcjDckcbMq9q3rzvXYlNWQh23IuWsVrSqi+R3ESWU0
xDu+KPh2gZSRjYEUhrSk3+zmy2mcHaMG/Y3Wod7KwKseUKKp99vbHIAhupgHQS42939YAcXuFYzM
zcpBSzxcaThe3jAXpEmPsfIije9Szv+c2qe585pK7zQiV8BLNEnKhf+V+Pek43XZA4h2T8fK3LLV
ZN3RG+KRZ45c+t+NHHBlu0s9Y+a1k6lpXIjIm6mBWAfkpyzg5pspLXloU29wCITjfCZnN7wTGuCw
ggma1B5qO9JCzvEZJYkJzMAJXb2/8hlIrQSxbjk3civH8CU5wSVtsDjYYdw/3SgUfBotkcSDAfm+
mp5nbnvRvIqXpBbq2KZLkV4P1iBKYGYow0i1npIPNki0VkH8fNp3UkgMrXcyR+YeOgTv6zUekdui
DfXkXwhjQAwVRyfn/IIVH9SXvj0b984ot2TTSH+dM+33C/YTow5hOK3dXjPxNrS1FyXQnPp0tBJs
lNU7NGh5tZ7lq6CWzw5PXOAvIpZglFuaD+22dwQ0wPPN9fwBY+qkxQubSN0oNa6v98SNKkQ/jZra
qom4kdyXQTNIC7UxJuQ0rA8CR4i3RoQJhNcqK23bLbNmJ6I2Lo08GpdTpVDe3sioHJ/+I1K2wJ2N
2FKOCVhLR/YAgwH8wu0Z5TkmudUXe52IyVLUxk1NW1b0k46TzjWr5fWqiO0Wtv2BNQ807qgdtKgO
vomelaoPiQ7jOqturck8EADF0tqR5PCd6eHLNxkY3mpR8a/TcqS7pT4wUXsNZ8oiInY4XUFXlpnS
XmOEk0IZmvl/fLGXebRy3VLdkf1xufF8XVYhvL5NScLCzBdOn0rh0sDt9+FRtRFa4HfgRIQbIyvi
0e3TnfIm/dp+ydPMw5nrTaGit6x4iFhWRS7TXnP0M5ikS5x9ydOk+uKXAekfHBVidTyivTQxu0M1
k/OoMy1JMR9/aaKduak6YIuXM+9N4qjwG29U6SYrCcUMXqSVWm3UA74Rwt7ahPJkQcku1DB+9GsA
/FaP/DgkpAGwV2vSR6c0UE/U/zbfzWWwIyPhU6LscnES7UbLMCsJND9IRHZ9w7iNxdlLFlvUFp4A
fn1xahu7VTQlit9JeiCIGfkdcEGG6GD43DPDSNn7fT8dFtoI9Entvm94z7BuXfrjp8xhZ7AVW3XQ
YEYJ7tjQY/WbpC9HXEgaRJRPcxWFFMAUc19HDvuBvr9xXc4N0q0ITLyeEvpXWjAVBXXKowdgVx5T
mbDDxwP0MMrsq5fsDCphm4gWRATAz4vYv8I708j70PTBvSFd5+wJDZhFX5XPZlD0NElFs7EfqdkC
AvDgZJuz1BvU8yGiVI/GBdkFJGCee8Yo0BZ+j0hceFFQJzOXl8QVW09TxjgII/Z3+zckY3IgFJO2
1le72LbjutZ1nh5xa5DBOHJalxuxWHf+0B+rUMEc1g4ZLn1yg/PFOZpFnbCOH8AOW1pc4gBsteBh
xWxE8w2CgawaVmZSPLNEKJdzCFCA/0nRiVg9GEbAmfNtMZbB2VwxdjmytXWgOoH6gql2ulorHXXk
YAw94HLKoBqM5IUj1UZqjH2mpbGnOSDZ1x0BJFT5uvyZ7n2dufjpF3Vtx+5ojINSBM3i6dVo/nVP
61U4qRubqNtDYznvqBhzYx6km5tocgb3C90CQaDvxota0m7J2MDoNjq1wkFdrpL5BnLR/WqirdiB
yVEQCiSFkrLuQ263wUle0odBV9v7bqzNghHjotpsUIGVkuUcTbdU7crgBF/1Ld2u0mthP5RpML/z
spPGn/8ms7kQTFISN/g9M0YTp9Dqcwi/MyVcs+rCqgf1EeU2gv+JAblOFJINJN+yBa4aL56AqdI4
KRohj3tfJucK5rvKBt33jVoEXPiTNKL1KQ+2nzeJdY8xNZV1F2YT7hWla2Eq8/+HoJaiqhV8kKxV
DEy4tmRKkHLg8sSoagDL2ky1HN7ZC0nlfuhUSJXEV3HBkXFhyEug8wHgROJLjr04Sc6aYvD0NOdV
064yKZO41UThW2gIjrQcyc4oOuvX5jDm6uibfgeUuFj2r/GT5fjfrotNieikj6MdgmMYea2Zp84F
M+5/bdMv4s3n05n97GQszaA6wyyCRWMd//BmMWscpirN952j1tnQP682bZx4Un70iLWfYAuXxIsW
PLWrMp+KbXH8Bxh81L8MtLx5G63kTO9gmCAblZhA2i7VhSwqzAeD+/vwMY6MOXe5lQI0OkJ4d5xX
+l7vNcetnuZSR7fQXJvLntMO9dKSEsB/MOEXmjCIPo6R4hZRcPAf5ov7YyL6MqOZWyXkWgVjE0ep
y5Wi+4LKDK3K0yZtMzSL5rzH/Qm2RNsZ48Tt8ZXbpwLPq5m/MJhNzKdfPLHgldUnuyJqgtiru2bf
Uxysp5uEyXA8MkynOHEEz9XpWql5NPLDnJwPg19MFq06J8KP8a+k1qPOarLg4V1wDTfwsKoYYAeQ
qJ7EfA28ODdmKruvky83Lu2fOcAtJS8C0oJBteOaPoxqZ1lU/Ct+fBk/gRlkEN4hUhXLwt5UHHOu
LEaikj4US0/MiiSse0CmmMvHps/fXxgzNDlD5oGweKJMWcTRiUNO4uCtdn2cIGhUJLwZTrP2XWB7
ObXTZHuykA5a90Z+WqR12GpPqyyyeSRLuvq4znwL//T/J9FDX52wdiW3Ow7iWZsphHICpkuNkx4F
dbzxXl2/T9Sedgpb6Y3EowhHzEa/lVtFMnJ4tMTqgvsVJW2mFOpwJ3DlPIvZti+M4pGFuB4skhh7
xmxvnlhJQYiH2BQhF9v6wMGxefkVNEkXOXEb8dOG004W4Y+W2Cs+TVG+ITwgPDiZHYg1wcZW2SSS
61yusBaekWmv9Eog+kPgmtzZS1Cn4OHXO316rAmBuryFKXTidHSRkQhWhfmFZhzK28b/n/yx9zw8
L8IrZ4xEOtxyoXrIByuXC3M4TCjtSQbCkIzcznrqxECdmYyG4Kjc0Gzw+Ld46syTL5zWS1/NJKYn
YR//zI2alWaizctwrC3lq3HxHEmWDbtdr7Gt06HA4w3q6f7T2LUAp4J1AEkAHvLSSJ8GMl1+m1g8
o1lteh+4gSj2eLmjDUkjxNblAcJ/hv++jyZ2CRTSIvFKS+VXI7rKE15OUh/TytyD0nukMaqvDEAC
LfcnnwxjNGEIPcw993dQRUAY6jqu3y2ub37sjSmWHLObxYNhiGTSD4p+imIoNim82i1Pp+U3wyAe
Hk6rmxk3HgtCH74XpTKRxHoCp1FlSwmZLANkH4GEBpL/j9qVUMReXj+NzlzO3HyrxzaW4GKjfPhM
god9TrW03IfmMTCytNPd7R8Tpuh3x4Bo/P7rEdPX+8EhQWz8QAuEhAjW5N6FX8nyMJ0Mfr2J29fT
TWNGfbsbcfelkdJnDPLk7ni0jGcsg5JLrZUApR/P67uXsSJsTOQnkAboXedaaYlEckcjtTrHE3ET
V4qAgjqCcQwYr0xUTCUvOnfhYdmYH9p4jyE24z2L2nuV61h/JHenFR0qogl6VqPIKNTkZXIXzfPi
Vmh2ZP3kcJovHbH1WB8WQmTsXbnzQkNhXcxSRgsBgZZHHSr+2LcS6eSFl2scpBEghTsl3aTTK4Ri
5SQkN15u93QDyoZajDpUqSj4F/WQvw8WqI49fsKEabUA18Su1mqy3gaVFB9alNNcnw+L71JplCY1
s1ZdsxOUXFOzhFYguquwSOFkKePgrcjUH5gsUOT3q08AFDGpygIuIJ1eVjOrak7kenI7TQc2XwJj
uqVoInAlJwj3yp1Wo/0+sZAL2gG+zQ9p3V36+WZhxj/6TQy4QxZlQdrBADp3FPI+777xBCIMaLWZ
iWHAcHtyAFmmp3XhgA8CnW0Z982bg+ivMXEt0aslY1ozM4THCzYrPler9MQXrYFLTmkZbJNlsacR
vqIfyQtHN/11EDzYSSAU/gQY3NbTEZDiNPWwWld3ghks5euR7F2GVQ/m2T6b3ElddkfzmLztEuMi
D/kipMMaA+NP+2YjxN+peGwzMioUDzcKdX/88jaE7LnDi0k+pyyDzAgdbm7XH+fCD6b5klYhOylX
6R4ErIr4OADnMpJZU3QexLsHrOXGbqjnjvojIGJ18oIyPmFpkjBsRUaOgJretifmo7WyRLWkhqz9
zUJ15Gu4giutQbM9gYJDzoGPfnj3tjc4wAbN2qyOuC/P4/3BbY6bofqTGoNrYj5fUh3RPYViAtyE
5IbnTZh1xydg8xKlxwQh9QWBxWw2URI8HMBNmrCyJTUMG4R09L4Ukpq3FUBjAkJAMW2v5MyazwqQ
2qfC3XONAI4Ub/k4/B1xP9r2krBnH0A21IIIOF//Ak/+wYOGyyVcncWRJwkhljLoWJ/sqvCjpSPb
tBydONGRv3WzTjSSLcqnva0rwCj9yD0om0iAgUYSPig9A3GugnTi+SXfnbjufa0e+8/9JKp+Hm8u
1gcIJENbwfAuOINEZ/f9zrNAw2fuftGhYxa/oJdWS1y1ngd8OgHUdhRrj32xEsbMniu18BBQ/HbD
HF10OhNZypGU4f/0tR105UJ8pJA3wz6FgCQd8yRunk2xqLy3+qd2IA4bdGBd/uEAmYd289NUbWaF
+bPfiEcQLmSP3hj26kstaSe5P1j60kdk5HGGpqDdEA/gUeu1vguPgiRFfOWJPT4x4FbpD+6Tl+EH
f4rCul+cuosa/3iRcyRbYHx3lmB2wNP00oAd/fRsrDFRwPl229gfUkUhbGHM9z/XXYpy+Fd5jtPM
GSzASDHNLXM/S4pHU13nm5+hMtySGWAcKmubazY6EU4iZTeLuckvydYO2CGUXshDQSt5Ou/hqpc9
KtfA/hJ/CkVJ0gIZVY8fy+elhy1sv+5Nu8g5N44dRv08pjQ/AT3vLynH2P/JaHUcR+uV0Xy/3vH+
m3fBwSeC8UgWE9BGEjX4v1BLs0Yz81YLzvegOFgDxHE/DMgVoZxGzqc9OGtKg8XtiJSkJSnpbFVu
0aoJ7QhY4bGi1QYXkeXfARfk63/Zc2PIMoFsfYEj4v3KNNtp+FXFyM4QUFNUE3xbXW1mROW3PLYg
vlh4agHWNa6kktANvrtLQTD/CnLxUL1hB6h/Yt/AbboEyyjiX5EVLzGZL+md9n+2K73zvokTR7Px
fiWVjWF193+zBo+U4G9r2LqJmvteStvTkdWnrdPthBIqF7ebzlcItUaSRrMj2iSzv+puCtcSs8kv
C4kFe7hOUKJQGf4abjvH3JJo2sOcTNE4Q69Km+/QaJWIvA8hyiu/aXuUKEdumOsUw/Qu3ZOGIFOg
kgf3C0jYrAin6mshQX2ySswKcOLcDAv66ZU1s0CGqTuKtKvGzNxxDbn36Ua2kf4X5W2t3QsKRT+/
Zp9XUW4W71dR5CV6n0bIMQ2mz7GniVU5bQtCaNrdwdWmKPdu3gPDXjjE9uxk23Ryscu2X4TSc4Ma
ttaDyyZhhnvTP1lvFipz1qn7797KFH4pljiQxBJ5ILiynHoSkfzSdW12A6RmsUtsxvNGKyQ0DuwW
qdvUYbsI60nthPz9ULcfpCaF2PyD44bd6TzlwfcmhRVtPEcMWeVKPSX+ldSSHZO485kt6V4PVCpi
1HkhcaDkxIUxcbrp9BMREhUjDIlbZLcIuaY3lh231MYpbbZF9ZrBbkSvvnf5y/cR6BOpCyAmcTjp
o/R/2OO4e3OZFpkG0H5px9L1r+0A5DGOhvp5NVHVOaLYdJVTA3WMOVDapgXZi/8BQZ03p/mUA/un
rrJOaypXa093SOyTlLubHRsje1M6x/3lINf8FxHP+HLqTLJ4xyMPfOO7SgoRz9PPhzANa56yxKwI
nLGb1bCIblT8v5OGdDm+RUMqwz0s1CS6KmsHFx5fkdyyU0g3qnBitLGmVsYmogq+vBL2UOZRyGyL
lr6QIIDbrwpbGOySiyISwKMzvVWJimtHBLdVJA7rU7pvK+75kg/etj5rlMb8JaQb5uK3dNMtSip6
uM1H6Y0/DUwavsRWE+YNoIJjanto3kUWbdcgaC7/IddcwNB5N29sHxT4B0bmzcKRlqqzZRPaNPYo
cN5xQcVfaGeG6uHpsyIk6wk95CrOVLbIsKJlnFfZSyQ36Hm/8qtKIt3JILOBBmqXw709lBwHKnpk
AR/aPHdKSYPTRquFmJ66etwwC6UmXiyUJr+1ZFhY1Y1CM6+UJfV4F8I1XzkOTVjrYp6E02Zzup1M
yaqMmINvNQ8RO+dJx1PicU20L/UPofeiKSDyS8maxrwWlw6LzHZrkB62wuVbOfH1SSSCFgu58CrZ
5NREHha4ZbJvB7xKDjHS8oxkmKJtFWgrsI3Bo+ryUhsQTpS/nbkyZkmnpl2gA5r9lFvnVLApE5iL
VAdFRWauzCz7EaxdOCvmWn4ZRbW1egSrsVAov+h09pdw7AA1Q/t8ySLhU3BCOWoB0F/aIKeXwUVw
Z9eyszj0bNOUvXzZYmPeQ0AFNjR74mMkH0ZIdbCzsHzBllKnUFfEqV3QwwE9OQd+4f4ZX95ZdUME
7LN300CSpHrbenzOqqOYAwj0huggGoRigxPe3Vkivkzad1o/29+8m5SxR7iMtVnIucpitXFlS/Ku
mHZBg/Rz0a4xsCp9JGHdI7wV8vxbuAJrEYIhy4ywzSSf081yrUdupTLAUuTT4PjD2IPsCOifyN4q
cEFshUlCtymigfj1x8Ey6Va6PeRx7a5ckYdGpp6wQTMT1rb/LljtewLH4LCzw0xtdxjQLT4vwM7r
8IxfBetY84wgDFFqbgcDXIM1GXrXGU1iVfAJPXkpCSh89D26POoWkhdxjV7z+CvmP19Y1a64Dfvk
5Q7FynRBUZCS9uyofI6bsU7T2XtL/toxXDRxHayXlRno1iZrwU/0Fwq2+qAVcwLv55OxI5Talntf
9bT8fXXvR8SQm4+H5LIWs0t5UhmfnCspBIfzGJ50aOeT8nOVlQFgxaQ85D/mei82zKC+rrFz6Xxq
0n2CjsFndzXxmiZ87mdWT/K8jasNdg3HxXf4LNaLbsXx0NAGMIUt/02Bpsgl4zXXy/S1+DKNlXm8
7zLTtnX70oozBn+YHIeX2waat9dp28eRUm0p1hg81pbZ3PANCzxbWPktxvl3sTdVxP/xcPew/5yV
KNcoDFythHudVKgsBjWWaIK6KGzuqrUx96JfYkauFcCeK/TFbGfoXkjHtUr0Oci32yNfIOXhY0NA
+9FgDel1TE/anvksnL8tqDhPwqDkB9TnxtqBoGnv0XtwF3CAvxj66ZDsShQYIlm7uIhERpgZYQ0i
vaa0sSUmypmEnsXLTwKRSw+gzFe3FYZVVrpFk1N1Xdylox01LicmlnB3CZswuOc7ejAN5hT4/JKC
NOxE9FAOBAJOEjBJBwRkn6LCXIphb6vxB8SuLq3u0iSrfp4kQTYI/6DmQoHLc58IwRk1ulmjqAGl
4BqlcbgL+2t9ZOfLtygSVaCVXTyLLeC8DLPCIAuIxlMLoPzVke6R/WEwIkfGwW2eNOWEtug8yvts
VPmDGHt181BMKrIE6m/yx6wq6YxYipfPggGBZnKNnIwXJfgIOdVm9U6zZ1C4Erm5PH0JuzOSH8IT
ogeBmp6xkEGTKUjO73FsqJ6vLCHjgMaOE6KnovqaVkHolQmJ2LLj13u9AZEgzOsF6S2R+FxN6Xmn
M9HLwWK755Nn2a4WqgpepyRrgmn9KXOxuNBIfQhzeUMCrPH/ogi/tISSJBdn202AxJIYhOKxNJI2
UElX5n6yYTB6o9Rkr9YqS9IoDH3ZB3VUnJwzwPjVMq8yW+YDUj0MW9IT7nUhQH9CON0rRVsYl+59
AG2+zVSDNgbdahGzY807xNK7I7AXjRNthnLTk3uR9xMH/POiKdcv38CpdrcU4NnAqJG9P5zP8NNM
n6DE86xpQYVOqC1Gj4w8G1n6co7b/otx85hFJwnU24Dr6lhg/ALA1peBCpYnDQz7klU4tqJXWXeu
QF1cOSnGZHSjPIBqg74Gr7rBCHMTALRqdqIGgaSMWyjFMMPpZ4J/lsJvwzk7/9CDBvUyf4jmR3NF
qhYj3lqhMhNYWqtcjk8xaaK9Wwbi7ciEm6EI3EzETRD+M2fffWyFZHJLjCo7V3thwcv8zEt2EWCW
pGb4mN6WalpGXFpDZd5j48QNFoWoNYoKmZEpUuv+OX4cBN6NUZR/xe9gADC8jNh229JZ1H+T5+Wu
AbQc2+zXkcxScVtEF4Z1O0t424Jl9G162fb8agStWZD2ENnHexLXIyme0FveqDOE8BbNrDTqJ0s9
dPBVVb8y//YwMjEu2fPp0hgRDfsy0DoKJx7IwMZy5BDz/EGC8kIQIq+6AnmAYZFQlDQ/81xaW6Cx
UCKVgVTnY8Kb0qPy4cOeWEKf1jxnD9nz/Rkk43E0fWwbaUGhI5gJ7iKn0NLUeIlIaaYu95ITzPow
/o/NY+bfEcdJvsnC3urf7ccsLs/UgmmolgWwDCKSogdB2yHAfYawTLaE2ff79WFtynddzNiQ/Fl8
KMqIrp9qpDsfyI2eZEk7YLGxf/l6zrUlFTVPSeo6HzEgsb3q2kcAX0nTdbt/PdaKGf8UpxdBylY4
E9VfJCa8YqkXzKEg16NooeGU9uSkgnRCMA3c7esDV8NEUYDovOB0DiPOZb+9VFPN1wD1osqbOq9y
HFksBTBzFZQbkCNb/q1lxKrG2ia38bf2zSTtjqfifhB627v9xusIp80B/i/8ZCokGLHMcEl5gT5+
46GVvqcU5uLtnIssWgsRwtTncMKU0V2a9gCZIedR5jvhsmDyKVvhZ2yPPIbs5KIaY0NX89R3GQYn
+cWp/tpb4e+5hrruh4LpLmisfK8tE1/2MZiAGziYwDLYtxZ6bYhnFA1BymU8Ebx4aIZznhTzVDgJ
+65wXg2+uXJReC3Bq5EOrjaqu99kHD3I721v7KEt414LrsR3zKH8HQA+9UUYWdtCTUns7bI5Wm7C
h84v9nnqLiiTylPIkgnt4O2JbAVf138QalH/GpfnKi0JiaxafS/omTDh1mJxgyzCW59JbRNA9sB6
xJWwIPRkK7EylkZhprcqTLWLAitimFJ+jVbDIEUzvgmJ40DXw4q1xH5GG5Fitajpr1DrsAFIDaSi
l4IIAKgY9uE6xfAPOfD/r0SFLtoUpVonQA+oYlxMJjEnRyUUvsZR/9oWoCE4/spQKABfC183bC0K
0O0HOW272cflDSi/gLZQqElWX8ZmO49p+IkZEXWoJFogGWEEQFZx3ec8IhKNF/Zx8YwFh0ar+FSb
4I8MaN/a+iD9PioX1FGnihXczcvkWsUKaUKTAS6sHBIBgwwpRUUUWKLqqiZ9xrrO6xzA/kJpibEh
o9yRZ034qLFAxvrvwo5SDKeRmvij42co3XQxSgVW0Zip4qSZ9WJPYaWiNIMWiQpukOw09FkTfXPk
oeK7sRCRW9OwDPRZTTrluR1TcWAC9oz9Aa+XMj1l8ZoiNWUpHz/672d71lB0E2JrStCiti+WelLo
ZiGDvffhViq8RrqoNHnepnavCChueS6RVMevcVbSVhiJH1YBAInBqFqz3Q3kESysezZ6UjT9N75j
dq8GfBR8VOS1ks1gpCAEhTE8kMhF1yrcYMENfmOThZuheS8rUvB+lpkFjqOivWqr6YKOK8zqIm5d
qT3vS+CLbwIPB85IBuyXMMfnWzwZxM8hco+eTawvI6Pzgrw630rQZOpTw9mqRHwrAJDtHDzlsX8F
Xjy97yDnXlFJfG0Ehg8HlxkYr5WJmP7nYTsfz1CE2HPQVTX0whWoGtZ8ZWqJTzAdJ3qPw375gkAp
UyDMU06v/U/7nNjbVMbFGh7S5wQdMmkc95R0pQ++/6oRwKOQ+hFdfO4oJCGnfHpMqwYgeYGL7yxt
EACq5FKQnNQNg3uq+dnO8UaPwaWdL8V0OO/OjR48t8in7yP/GgBUZrpwXAjHIzUGtmH3+DkqXz16
m8j+p82LG2DOsZsshT+r/HNb4jjuqxViEFFxdZ4NanXd5LkzplQoDUxltQpN5qoKrAsOwM46z8VR
4Ko3ktVZPD79V2G5RG151gy2ofWs//B39MM93MLJKg1Pity0O+yrIq/O//yGUlNjDJfGNfINO0JG
B+9dCePLEkHOWs4w/BCqNK77kvM6UR6xR/WwuxW2lLw8DGClMeq81MGgKXdmhcshwgZAE5ixDKcE
CFSybbh/2+rA9fVFPLxzEVpkorbSU/Ds2yCPyqwCVHH4VW8GFeehbSNc67kQweotXRBKwG2Sho9y
0Z65XFd9OaKO9SZ4VJ+yrc7EkUAyTWe4Y64Cb9zV2cgWnMdO311RsF4tMhE2+OrpmAO0UHWi1ape
HBAf1PQJUCzs5Jc0QkGlkh6i3NtNhJsQJiGfGCZMPSEPnqbzejjdCa2zctsCR1TGTXjDdtqHAaWs
oHZWvTTCLWDQZpTqwKAs9sQw2pssF41y8wxqMFRl03fUDTDFIw/U0EuS8dtkqXimMTf366BDjPDa
iniT8F3g9OzyvpOWwKft+AShg12CmfEkbqyZPbchnTUbzrPM9dIED9tb61KJWRvdjvHcQ5Rd+APJ
BxU1xPH1EFpPF9y+4KH7IGK69Kbpg9MnwG1XtUUS9RfccEDSLaOfyTvkJx08jxEquryCkbtPlXKV
aj+FfRmQoey+pEfO5p0JxlmIgNfoCYjzGqfgpOCbRXtqEQYrdks6DXh/Yrb+3H3Ufm6of+KFfUOg
+1I92E6fDKCsvOmkttdbhmhhk+2xcC+GCle/MYEfgi8WWZKAwan5/J/IdLAc6dzvnlI3RZvMHxKb
41iSLACk6k2xpfbwN9WeSNfVTcES+21BLpWsWHOJua4r7wx5lLxPHJIrfmWK9LF7ihGPmeI2uzXs
S63es1+8QQU1GAnsBvLohRoy9j+u52yCjTLt6Ui0owaE2UAnF2gl2h0/NPpV3CLbvapU5xY9vHfL
mFu1TYJBYxpNf/kTTxqUNtJqg1AgRxvlRdf/SEydWKaKtpTg6G2EReo/xAAHxy408YZ9t4mdWhN9
g2AdMRQiV//IPIbGRlo0Z0ELFgUxSXVDA/Mu3HgR4yUOV/OLQRrCxxZxZfpx26jFeaBmFaLxu4xm
gKxdbgxopLPU6EONiFHI/y1YIFj+ZQ5tLmXvZigg5D/yb0SCOTlsVaZCKOESC5ai/4Ls6yIL3j5n
rfyzmq8m3mHQ4BW69N4jTzCeeQGnpf2VGLbkK9XshyMO9AJ3smcoGe6AxvRtKYVC4uOpVldWLpox
ZRBSqGgvyseR5AqceemlrccuG/rUaXy+itChJpALd+SlDIoPSaJXODqEG/8mOx3677C34AvU48CG
pORVweWQ+m/EhwcM/4SIPS/uaZTm2RYy0jyN4x+8/9v9a1sATjCXsjhSgFtTysgUrvJVURykkYEt
dHwVM+5/YBqLpZkKZC595uV4Purw2lv8UXtNxaJ3aVdm0tIkny7XosHScVBZHPgXcFQMS5VJnKz1
zAjePsd5IDt2IPS8tmk/0gW7GGBYemlD50KrCCUL8L3Uco1XigbNaPaTnM19O0iLB4nnb/RFnsGM
nzSb7H+/uJkBmw1SbNJLK8CVH5w3GG2itiO65YOveyzDaUaVEpToHvvHvEpA6PCeQx1VPMIyqg2H
FK112si4nXX2Oe0QyXHOx2qOsjFWfjCAxo9svjpnJZYNCV+ZPk4Am+r9vvk13T3uUhvNWcvANb0H
6aynFcFT8YaYzrYrEtV1YVWRMgBvCqvmXLuJ4hncYWYu/vYud1bzlcwvF+mqxxo9GEROqL1ZNaLi
wb80IvERQfuBqJ+chKj2+k7BCoriBMy0gmDBwS09Z0O/VIhVNHnMWY6fmj51ixfyFEpiImt4/AuN
DTQoJen00n73DbBojmIUkDgOCz0nODvOBgzWKm2JeZrQ6+r831Bpdv2kBZ6Jfad7UpMiqCJpDamC
DbRKWKm1dnpwIRXssBha1YlvKZaQPyzjH+F5xrmRzlSxnbvQ3xUdiabpfctcTD6G05zPNXgTKMol
NCMN56SYbdPG5RKjC2/E964xXoNQJ4ALEqjjzC2bNN8twbuEPZVCp3dmrAygHR4QsJtRoalmQLGJ
PpDEeVlRjlAddlU2hwicxnW1oc0YiblXOmHKP+l1Se/P/hqvGxR7x/rOpktQEAASTztOjLw4WaEo
TO5CJI6atZUEWl6EDkjqx93uYUGpPpbKFhfSLjwCQtlKt54if4wgFTmfaz3PY8NS+wvJFVNHdeP8
SRImn0oeUJXO1Sf7y5w5ucHY/sDSp+oPRDbRUV7wGHKoOaYScRZj+331+hyg3QBrdK7HhegEoTOc
czGiu9iGGRKPyLxFops7Z3lBRzFh75E81yfS6V+d+7DyCj9/DiMX29vM2M6UsywEy/RyIHLTucQ4
QTGUshVm19lb79GkbooTv3tAIZXwhbvDqRbkpaMa4bUa87J4oxAxD5ttgPoce4C3tH1vMuv/KglP
jJSEzeAQ9mBg+jV9ieoe8AHNDmp/4YuWIYzlp+SCp2e4SPWHZzs9z8umW8cEvo/tixVUIAL9OIDE
6EoDpJm098mooJGy7e5Obz5ehDW7Ouq+GJJ2OdI3UJXA2Fzx3WC1/GjoMFQorIvN1KI8N7WbhrGe
4rp/UL4QwT12YGZweqQ9O4ALq2YSkOD00Ghv8iFWsffkT7y2VXmzjptpbFjY13Ov3eBO+QGSqb7D
zlmBNogr/06zpPEUsySBJdgIWYFDlU0Ad1B15BKbWDn+oM6GTtPhZDdPE/1YSr/ux/6AC7kWVcik
n838+wn6unPlm3T7mjaShDB/jPKaKuSA4/8g0uzLl9Qo4Mpdj+VCFCJcfNlbSluwFSwn1RPRcVAb
ENJDpyFhnw1woZsTOfjU0U4NUt2CN/sNgKpZGhn1ewdJoY9NVbP6zqSNIDXtpy9Hi38vWfE7wjqW
7RZv14mLvcUeGLogO8pmR/DHWyxjhWPHdM2IKrkf6/X2wpGCbzRb+IADgNpKVuJKAzjZFuEqXhFh
geP1jSKOtAkYXginpfBQnDnGypzfsNA5LVx0Q+IPDdgYyjyRM1AWDP9/hLZonA0AeNXbKy6t7oNq
ZVbZ8z1JmLw09QIdvcLPiMOyURcQIQT/u/4HXCQmR6rGKIG+2JV5Dth2gQKdlNkJ13UR5CkV8nFu
dg0xErcK6uPwBohTNIY3byituPt8ePqUp00GTc3/VuRekqjlLCN4z3XqgFY287OEu9PuXEqLo5K8
J+WkR5TQbkT/b5TTL4v1wcR6ULPYlLiycFHL7X94+RPHrPCHNNS7PUg9rbmURuOgqbdzVnQAraPW
+YhzFwXfdYFemTJiGiO16iTVmGhEeL6kddZIz9Ris2FLViv0bVKe8SIuP7uNoU3deP2yiS0cw5fo
no2cMGSOIA/qM3JCIPznKYTFkolzfxxbTnWZx7Vja5afnrUxDr1SBJsji+oyrpnb3IURLB9bom0w
uXA3nBCYVnjfbV2AzQLAGMrzHBKQyILJXeX0fW3yqg8n1//Lq9J+bF4Da/DnRcAOF+4hMBkkdmzl
kSw/yIaeq8FSw6nI0xsKt+tiNOu2Jw5AXiO8M/cVuvzFxetqw53hfKzZdXGxzcAkSc9fl3jllM83
pv5sF8S3vh5ENua0B8E45m4oh37R+siIizIvmu9QdM4XSfyRG3bwd7kNhSSeRxvCCVUMy73OGx6k
8vkGTE+1ogji8GK5bMMBLfFrXLMumpXBmBiRvAlEHWORb8/q/2L67/uOfmxVYCyRlDgf3D4RriZA
ZsZmnmhQMMQ56Uh6uWMWQ+7XyERM1r+NmIfK6sj+mL1Nii0UEb/E6xVYfvgd7hRteqT1V7Bw4tAN
QQnUJ4gzkNaoMhwq8s+Ixdg2bYAFPvi98A2+kpVoZTYnlyYoyx4mn6Tu3U0DkjvhNYlkQOqokk93
gtF7BBx6nJQVoKdhp5Q3QPWrxBZc7hFh4XazD8gXvM1j3qcnXcRo2zH7/KgfieZ6jCty2R+MOaUa
WdM4rmCUfTWacClnhc9RyAtA15gzrxM5uxI9241zIHwgq396gxOq2jvwwGwXcXv0bhH8AKRecckw
p9yJeFTGwmI1FberKsaj9SER9Q7HPJpqSWpqZZmoxzMHEa0SMGMpgf/KuAFIXGBKT7AeOfUyCCXn
oWjgyLZY/3dmB2yjh+u9mu/7FLZ3OGynbidksazi0Stwj+C0mC7WV43ReeQWFk+2+mlW9abEaIrJ
63kPQQQ8LB+gU3zfnPPWMsXBPTLuNJhoTuo8x0Q7I4Z+AWFdtBJnnz2q2zhDDjaUBRzRh/VuUy+7
OqXIjiRmRpuGQRaFZOp3q5D5XfMyP8Dxu63NG4e9hFzYClr/H9UmcVvVQcumAYlENCUltuMox6tv
TUmSqMtRQ6nzfV6Gtjrt56HuA0Lv8Vms1JOpEDI1VqNwr3dM5EUq4qLJmcY0N8upDx1qNDVDIm3E
LKKUBod6JBMLto+FoQI/SH8LxxgmtbD/Krzj5kyIV/Jl3p3hk5S4vET9BqoNlqzT3tMXl//0aqKK
a4MMm8C0PHQIEDbx+aYJg/bQpVs2aTfghX+hzba6VBN0q53K1doZgBdsgEE4KmT3dIP3YTBsDEYs
eK4PlmN95Ofe6CW1em4a/OCqnMCNyEWZjnaAu+xi/9p1+TASGKKrX39cdO9wBkf8IFNkiFismZx8
mLDNcbELxjiAgt7gLd6EoGl8POgR41uhW8rOVBGdQzGKGfujihezHOznZbCT4uejFGt/LYZpIPpC
hWAtEzeBLR7Hagw4K2NB7EQvd2BoA4EPCv28PUmMo2yf9GwRJzH+Mo7uiWcGeTTjLEscuB2iXsJ9
YBS8qKpykqXoYOkYpKZfeESXwwnQcAGd94g7Hxx9vW/9ObQqXTG5kUsuE6HNPtzbKQhbeOVNZzO3
mIjdXEk7h42LGLbVpOhIkK7lk5w3R4Zn0uHXL9+Xb11m63m90NIAJ54eXK1N/k4/ylKHRAmrBpaY
TO3dUPMnpEI+PpKkugNstrdvU76pqbMVzR6cN41tektCuAZHdpgakAsR9jC+LL7rEPpa6pqgWdsV
Id0ZIm4k5ksN1aeMcYXhSfCnVOC4fiYzvPQjDXeloWUgNxx3W8+Rgwa/6WMVpYc332Gox4wkf7wF
JPlV3lEXFvbetGRjSdhoPFY/sPUhkeDtF1GGP8FCXnjyoTEX0Cw6C+y8OlCiCgrb+MY+JqayGjZZ
XnvSEezNhM7E4MRAvSNcj2O7mDZpXw05T/YN2eK4mIxkxVnvQ5TNCMh0OJ8Qx4qrx68ipidaUHSW
xAgKRdlfpYgVvA7nHpyk0BpvyJk6rYiuqRhTRBiyxM+f1rdRRlsi2UMjEs7eLrJrqHEGRepXxGgB
/TrWCxB2iApVW9LUr+JnRNyRltyDz1lkAhedHxDGAhphpyWXPFj5DVIlhnxucynsVoCk/W9QOcKr
jQviN/kenBHIrTNlhg7ET1qbcZNX4IfeNaKERT+dNeDy/711gWjZDH8GR6+NEZ5uRrjQ0d7XyJnk
WlDTCIyFOOTHqzcb5uzsV8HPdx0GkOF2QshdKE+VWecXMLG7FlfeUub1mB4FnCpZqFx8xBEoeG15
SNeLKDCf0OGNgjZnot1JSIzWIQzAyWwn27JEERI2l29eshxnPvrvLl9dgbcshvFUxWUba7Eil/u1
84zwTgKr0zWOoen8YKKXglmqnsw/ozfunRG/GKDfvd7+nKNxjUn72SIRzIeJJdTudIVKDGm3sVkS
EHjWjSWa2Q04AcUOnxfAFo6SI6RX5C/VXRivhimVBxmt23KEIUus2iD4P6RXxRlE/VCuJKjFFYe4
eT6ufK8TsMoExYRwMJ3/OAbEdKxD0QvwNMbO4QHY75Qxrw6MneG1uzebuWOhlO0juSFTmtZZEL4J
wCnl7xUvQOdwdh8JA1hmPsumq9MK9ATLP9eI0WQOOKwwRDur7mL9ze8X4LOhAnthpCCkSsES04yE
B0//KtWzvov23dxAd8rVDJb0mB/QsulB4RL9wYk51lMiq4P3KySwCVV7amOZiC44W6Av3tIlXNE3
rclIEgLBxWIXXstbdQIA/NSdeEnqns4COqla0E2P0bnj84aqUcs4dES1/gXNtAPJ0EZDRScnQn/Z
R625F1LIYr5/hcRPgQyDRbGah81WnYrxwMvOegW2VKXnj2tDEL/qWuNIi/tRZumqRLDS5ZEjgaV9
0gdjfxi93cyhIxdsqvfRU9B8EuETSBxwc+TZuWmGmD81kCzh7NPQ46eOQbXypWvQlfKQ4EHuFGYM
ncV6SKD9+0LPBtBem+YImy4UUb64uEupGoNZ7T+g/IBVT9erJSevCPSDMyfUZ+MwBrqjuvNXssxF
aQvpCwxqh+nFbO5c4zSIwVNTH1ku+IzRH43Vi7cIq3h48iycDLQunZcFc52AnlW/+aDLnrl3V02K
T/CfI846K/In0hcAYqgqypKZJAL2QaGDaEdtBXz6b7WJ/9rF+YqVzJQlOq5/8by9cBa6dzLAPLTD
LSLbKvIu+NDfApY9JeKKgeQecTLcW4+Sgjw0yK77SVWOKAXS33mZmRv6+UxACcLm+jHhDz45POzv
GBGbafytkI7tbLGszKbImD0BUlHHRpGAhfYviHOotKRiQojRbOVBP2PhfZdMVpDiz2PkALmVBEri
ltmXY2uaOKchMiGJ+j0syzV8+j9IEERzPXu/l4V4+zGLAMZl1wXY+duHXRPLF6l+Ks6VXLQ6gwzz
ASKSNIPp+8qxzxJrOmY6A9GxWKk6eVta0CcnDxg2ES8NWkcqnqFw/uF5N4gLdzwZuuwqDIm2fMwE
Oa8+V+RurALuwwdd0oL2F6a5ga8plef2BQLbTi9CJk2B0pWgnLqXuejQc8KumsajjNYjfukalt9+
EcgV2dBoL3fjV6n943Fz0Bbhv2czG+BOq/kJVCc93ySn/+xFjefOudmSnyvvU7jbvEfyCq8IedpC
t9IiUtZMNp4R81SRQjskO+w+sAJjc8aOWJFTuzlfeVbnCd7uTtqfQR9Li+K+yzMorZ4mohuScntH
mpLcZFPbjS6z+pmXvXYuhlF7OmcVVSWsZECDOty7roI/uXNz75Hv7ZnHNshViRyVljKQHGn1ns7y
Tdb5oghmuVYPAcf3OqAxEX+kVbs0MhnW/bBEJRH6r2cV5w/nmtnsAC9rqMy6lpWoVDM0C3EfMkNz
s4vklcTst4CbEp5tqcHap0Fhw7h6HG6rKW2u0OryQqwNt8ekp/PQulETz3M9E4yjJpuJ5NlgYHla
eK1RPDFuO0Fh2lc1TTI8l84S4md6Hc5tD4aWHQl639TvbWjCCjqpqACU4KiBBhbewbMar6hM0B4/
xtowuIyWhlUcfYvFVoHr6bf5eA2w9c0x0n+ndC3IV1dKzQTc5DDU1zH3UBbkHl+ybF6pOoTycoRO
RxdyGDkDTtzj00Wq3tvCkmOwE5E5IL6JePlFnjsnryz+9J/OZws7MIQSzPlQnNQgSVAGYgYYtOfx
8urdWPEdUAMBmweBDeY81u7J9yYoDjtFstrDjHYWVsstO7O4/9Kc2QWufAqzuPKHkJ2Hz41fK+Ej
ypzdhptvP85CP4uNpAk/Hj4vAlafCrHctssStmNNVCnB4qVRWtzs12/aAif7LOPhPO95SzLmPzB7
QdkaL78tSleZA7QdPvD4leHDLY/yUKkbsdinWM3bpwCJK/FLq2L4agmlHCZZZ90DsKNLCdL8pzip
rY4jXNP9BQkXlgQOlzMu+TeRTpKR6y5od72v8HaM7tjqE5NJDmucdnxYK4yQrE3ZZQx4zPSeJ7Ez
IbhB4Jn8r/BujW6zSWsAqTSkV3ZrN0FeCZDuKt6xH7VlORzaOim1+QTCZpgxCdSRA2yAJtowJTOi
Tf8mf0/dj+d4QpVc7Gjx+o8AAbF9wlbRWQi+1iOGKLuZlIUhx1kdzg3rLu9GLohM/BvoBJUcCjmm
9T7dfNirprSlMmyGeUOLLNO3v/ANhYm2NOOxYql9E+8ZfPNOP9zjM/JT+38nmYmywgRDkmtRQOEU
3iBffI56tGIQSThE7JWKv2FgZQ71dqopve5o6JeitjsRXs6qgLNBshEFXuriKh6PBxH/ePRo99/J
fffl+tpBbxB5yWP6ScdSbJxIFOJLF4yKavx/fuBpG4JXDKue18OKxfzRf6CMwi2R3/z/9Kp/BJtj
iZJ/aPnnvs9enSbvY8cu15cYibJNL8bYPGDW7XKP5+eufBMZGUaNK2zNedrYoD1EOtARnaxpFT6G
wN9nl24AfKQGkpkPm2B2fxFzlv12yOVm9f5yyYzv13B8naKMQoahlawdZ4zISyetqj6rMgH+90B1
s+66Lk1vGUWvIPOTcmOqak77G2zsIR+A/PhuHAWZZkHnZGtle4jBw8nCGksbXJhIT6cqTUZrgrXk
lUkcsyo1myw/YtjqsrI1NbkELYd0F+ps4uHoVFGerP/Ddh3IJ+UGCPthNDhOm5Lkpx3hGLj7ugQr
gGYg07+8b14A22mM0Hrj6o2EIIARDVeQbqO7L+N3TCv56peo7bGXili+CVPz1SnZTs4ungoHfPy7
rZSppB7LjU+Tkt8tACHnDchudjDeRGSxD6KTjW5cddclmSSHFk3CHG4qS0H0c1VDBBsOAWypW8+B
BNcB8nu7FO/vX3Tx/Pd2CbGb9x5ae31DzAo9aDOA9me18P6Sjg1KNzgxudf0kKI9hHlKRx1vL5kI
hwAVLYEo/cni+lxTVy12RGq8sIKpscD1nVXTOoU/vRpMBybl4ynjiikvPgZtOz4wbrM3zvFzeuww
775oHbYv3dQnmnMmw5728Gjm0Vncq6MixqnXGxdh//q8/U8GLRNLg+lXfi7l/5h80264X7h7JKia
ZSBwTqFg6C4vvJbHUFNmKa5UP2FYYa7nj8kHtUDvIoxo640OC11G+xklXccx0IpEve0T1oE4S2BE
yJhOjKrSkJLdeP/OOm1MYPc2GC5OLBioqm59rMXSI8CxL198KcqIEC2BNdsMHJ6ImGjdMpK7COs4
fBfmRI/cVMi2KUukBccdVeB/zJ5FNmWMpzQnJF+BOy2emk4LwyaOpJQ0qlFJ8gyn4QFQ8tjqT+gP
I6QkXCPFNMhiETLCDyo2GJYNvo+tuRMQzfCWwf/GIM4Ri8h3v6SL74PQBzUHldLsGZYCTNi9XjXy
GHhaECNqY5tlIxghuGaLZM2A2p1b4OhZ/RW3MrrIoc7JEkxghkk2DQfbSMrZd/zul5bWptSlznGm
6SNlhJcRCwQs9n5ExI0xuxMcKFskYG2qKdLb9+iuk5Xz8nqfkdHBmsqoC7HsjEQT7Df7V5omiqbb
xDYVafj6XUuShAHLvJCyuXXpvfhcw5Nk9U8O9EpyqcNIwFvBX63u1Za1jyZr+ZkLyIaSlCMv/Yyf
RlcjB54sc1KlKbZWDX3364FDzwIGM7NR50J6DKm/gyNO2w6VIMOlAAGwtEqIO4oIp3OL14NaSOau
hmXjhhOOoXH6midmOzl+Ih7e6ucjGAUWICA3sssaG0Wpzc1hqDi+Iwi7U7s+5cEYiKTtP2edmi4w
rhwjX+uEVyvHvdtK9GmmiPDeRt+SmjmGftZVbzlV4vn2JdLY9nzHIsC5M0X84pm7v+i40A2O7byB
lGv0+9mWHoHR40TIR1BdkvkE60UPTj/0O7R8EDqIwMdq8Q5GE5TFcb6jWut4kQ6sYLeqsqRQf8q4
pKAzuoVjSRRqiK/1fRuAvZ8e3JrPAPbPis5V6uAl5om5sGGY83VtvA6ESywUg6RSAv06hbHHJXwo
YPHY9smryEz8bltJzKChZcWWeLvbAAIieHWE7NA1ZAU2NVeoJjf/qqNSFLISMgd+GDbRazwtfLzv
MDoBv5XqrupNIPwjI9sG54cTS12AhFlVmAYngQxMivoiXiP/9oYKeDS7mdZz1W0KqpGRLe08643W
9yT6LzYUSL14njywBbHlnfyCfna5aRu2xSXnUik+/m9XZWGnLUU9mkyWxubwgUqUq2raeUB2Y9hz
4mShLWx1VbbVGkmXZuya4sqf8BVto8rd+JvkOrRT2XHzxnuqZDDEWFUV8/S4LaxJtZaMWcWjqex6
gr5C0brrhxnKM/6H0IumY3mBkxVhMnw8DmWcVnzRmxiRMDV4zcWe7NQUreIllFVbi9x0l+aSRtC2
5o6Jbimw9gGdBIbGRf8VFbDEf/h9nOINr5lXtFjrY5qIAgbN3zhVDjpDXu237QbfrpTQLDyaKOYc
kDwh0Tl9nwie4uo61e022W/ts7YnVUcUC7k6G35gx4arNlzSaI3+j/8q8fE5SGgr0YqKk/lPRF93
0SvvIxr45RsN85LxCC1bGfeQccquMwu91d8NmL98xWxY4NWlN9HpsfSHoMrJzCohoFIrvJHIVP0u
d0D9ZWW0vTRyqv7F8OGEYCQ9D6lCIikirqXUPfiClYGM+KdB5w3adxn/EFh1zOorrOAL3L/9b4HP
aJo3VgRe8q3/uanLDXsaQHoDLToT5SJttYqnXM8xkRg0bagDDyuoPX1qIEBAouJBoJhDsElyV2PE
YOJQWgK39IDRBVujZB9sA7ZV7DvLflLhrNaMKqfmfaCmCN611ZUjedo1WGmQRFfLdPS1yPi/ZyRG
SaIETop7xzzvIWxcWyFrFogYITIz8V9hDdgi1sPVDxlwoMA2itItPlXUPqbN32HneI4mxKCa1pG2
TOxZ6wd3W/UhklQ63tmOTUSCb9s6UmRGhxhpp0ok04+sJzaRvTCvmtzDgC06xD6kfxRoR05Rh0Za
sfNcxPkh+vEgbyQ5lUQylja54e7U2FkqV4YCjR6RQg+PuR4JP3u85brqtAzq2KeYCinSh+zUAbrp
oV1OlqUsa3tyNXgrN4JV32JydQrfRtbKWekimE0n5N6uWmh5RTOnQWe+I8EoXxrUS2WDrHuYU2l+
2ASEz7Nn7JVDzXameUYL4eCHsQYAc12LNR2e2bdNI+tUfjWQeXjvumsAVRH42y5QOBQIkUqZFkJ/
JH73NZQgvqoRxMJ5uvOoOhwwLXihN2DPR0DfOF3btHMSG08hpcyp4KFESaZ1gtg/90lUCun0P2cd
xX/xQ2A7TztLA+vsm2+jXo8dudTMCuD07aoOoc0EafK3chYJ//GhvT5PNXCsUvEyxOQPaFmDFGsX
ghQXfdA5bokz6e4CaQs4uyJrYaYGilI7hoFpIgX/kqRZJI5GAly0iKXUTNe5kDB2dFHV4d7K3IqE
8BAfBIbfxCkJGQ1+mV+DQGszGXlbgMhThCBiJ0meg9mf4l+3xG7l90CFAP7ZLLvoSj+TlhGh5lzj
fGp3sIIdFNgjDsNCz/PTDnphXEnijrMtKoNZSBtpreOvZpaCEcS4Rob4cxo39m47A5izAgFinCqc
eQFYqxE/JfaWgwFBDJfbA12c74vMcVhQFZIZWGoxjanXdSZgB6OlvNkeGNTeCwcv8DmGePIZmANc
MBWJRem/Xb88sBstmAfQ4oLBVP/WdGB2RSmPY7HhLcWIIFeYWB7iyjkNCFNIcTdeAWJzYTbV41TG
GHJYIRGGZzj8LHlHup8jGFoTAFCKnhpqCGMUJpURBZ+/+v0xlD2Vwr+Erf/t8bv/5xGenSlOtXwa
czo8i6CLCKuTebOF/bfAdWVgNJV1N6OnMXkJitOESH5ntz6/sujRPhGjMevh4yfeQSMJ4q13hMFP
570tSnUISmlORn4GbGwAntauZnYZoYF+kq6PpL1HtK2MSUFL0LvmnmadS569N//xFzzmdCbTKyJj
GfVIUlAyuNH67ZGa6fPZePMkrAX9b5etkgRb+rA4y6DRpcDZeQ43M3HG/dr6aLeLtH2Lv1b838AN
k9FDmIjLlcsKhsPEqi9DL2of2KfUrBOtvlHdYhzDsfxYCRwtHUHitD0Iwlq+pSbodWN8vPTm4G7Z
d4FkTDdVY1vdls/aZCLwOplaXpBW//QctxHTCtruM9g35tAP0SeWgPby/OD53OtvE0BLhe2wH/ng
wtkhvzIFGN/7Jx/5mf4UXskL8gx/PnWlC9J59KlLoEEHnljLVivJR1vRWqr7lHd/LlBtTZalw2a8
xxMAnhuPNJopOg3Tbwe6x1giqvCGHtCh+R04uKf8xqqhXGugaEJdwyONFpPFgJNQJU9+SsuXXr+n
yyfV+c/4d31MYbX4GHI5YieZXEMAcEv6/0+F9ABvpSoAMpzOy3vzQMky0oJFtoM2DHSoT/oJS+hY
wN+GqBcF8IWVfv4l+1vVq8Mto+Lb76qlFGPMdQlzUr2s2JjXzATnMuw3vxi7r4v+OYQ3eruR+YUl
9jFC+gvYwrt3CiVBE2IVZSqEORLzOawQ+ijzs770vRAGOf5V8oNvzyGZa8y3iEgffwISVow+OMu3
lU/Q53nwiG1Tnc89OGOWl+8jzTfkC7x5wiX29rlhUIngHC9z+2fTpFHQI0QAPeuCB7HKVOE0dF8k
yP1PEY/6mcNczqE/biJ/vugK72IYEHp+X9zGq0cpayNfUmPEsUc3StWlCB8CaoiHviH9Bny3ltPi
UJ+7Qq5zYNBaimgFy4eeX85L354tvlL3JRsVpz45Wp7p+eYiLPokoowGUuntO+Hu7xVChYdhGv6c
ImRfVwYhVZBuhzfR5rvLI+Nh/NSJPb+AUTWX4u3/6IaxNv1P73ylbxJDaYQx4AZR8CQA5fW7ynJD
rFUa55/KjY1Oenh0hArg+PcQOXIXNflynu3ltqKDJbEoD3imemLbTubw09CPCTjhOGiSRPKCIdA+
UpGvSXpfmeMHXjivwI64LCBT7pN5HmhAMw/T0cw2Z3HTuK0hfHCf2dtBu37nFuDCsaiBDlZknlDG
YYgTueucBz+0+SGpPL3maHJIBzZ+B8fRZBH9iGWUk6BqWpPcMUxJ4rfpzafm44pZZV6o6Uv/m/uj
mw33dUuLG0CKtmwCEICJRKLGLrpeoXrvbEbcEIwNxAMcv1In9f6Hjzw7sEQ4Lqdw58RIWRt3t7YZ
84LTj49JechVslO1HcVgeQ9o9Ns8YZ2q7gMT0ub8obGuATeSERJC8WuB96ePeDnWzrd+pH/6SLDb
HQ+R2Qx5zUHTiKTrMtFKx313/kfDyS1VMoflUINXJD/OBO1nKCFl2M8/I9SoBK4w/3EP4uFktE8n
fZjhDe+aGLjQBej8Vk3Rkr/bxB5pMaxbF59LGBuVgYIvNEULVTqGm6Ux52Xl5p8s+iArVHHyk2R1
7DdLCgslBK1MrxCUX+V4He96x5rvN50vHY3E/P+WDl6XvP6Cu5h+jVhVUolh/hcFhyLfJnt6pczl
PLkVdUe8nvJh4Wc9ZO6FDhJW9sXgLSgRJ9eWPRTLzUayrjarNuT0ztUM/iuXDv3hTyyFIjk2yo+d
9tS1Sn6fPhLXgjxikd9DggV+qCEMUl+detD7bA186nZcW6mNagZRfWt5bWB7zDyq5MwyHPa1ghk/
xd+GOE5XoF1JythUUtne9RQBagME9ivljBvjjMvEgm+xim1MZEhVkvh/4odDg2DkMqcCT6OUX+Y8
bBokd/Wa+y+GrEq6mg+pIA36Hv0ozn/0Sz1sy/Kl1hWxfo4ZP8CU/+Wqc8NUw44F0FuNbkWFfTwn
Hjz70MjzlcMv3ritmIapbNBiTH4ZUCoMrBjapw1faNVrGapti/uSwJ0wDvarAiGcQlql0DtcwFlM
33CHcdB4nynSO88uK688SOLjgQxyxWSxX4VMxN++CPV4ZqxWXrd5vnIkbwfHLX2t7WWv2B6icLaP
qjBZTBy8SODlOwhtiWtOUGXebysjzHIVtNqFoH1H+KA7QoQZwTnJk45xLxvgaDQSCBBtRRftjiEb
Us8auHb9czlcmroVZxW5adzXR//w8wLvUfwg6W4QysFDhDui/BhUvAiufBQVlR7XFr6aotsPJtyE
5enmihvKxmoniyKAV1iEhj3L5Ft2t9zgh6ml/aj3NXn3YCEcYohhe4wZMdIas7PWumgVmcGbbqYA
zkT8ZuJJFrTb0yanysm1fCcmJODIJFuEiNFBeu8oUBrRm/AjKdZbUnxBg/s+zSHn8ncyMfKD2CMi
vJMuzYZ3iKXSpeo85gumXlKl1E7tnWeFtAt4K7Y3/8dANI486+hzLuxMQDQOs7cvZ9wia+ARis+V
hFin28GIWbkpu1Bhi9BFgi8e/WEmol0aK0kUQqVDkLwnS47zio2noxhuY6V+MmcZQTJ5tfFSXubq
2l6lJInF7viMX5SHOBW7viemB90V6TJu6TCaj1D6Y4SJKLpCDSnx1S5InskL5ZVMoZZga7clYn8u
m9VU1m3AgqgN1kATxAd5QwSw2EC0TxD6M8XCefpfx36jL8uTttd570Gy3CLKhhXHUcctJ0udc6Bi
e3bU1aIUnff2lt9AXw29myBCmKJN5qbH58rsy+J0N3L6W7JYsX59dm9yZWMyZJO36zZBG88X+4KZ
wsbqHfDc+84SNuPJcTZ7GmtjEXGhWsH6r9GF5PN3fkKRYYC5RAncraIkveCSQlE/He5H3Ou8/bAW
yLJbxufCKL6kf/VnXk464OCqETTbRAyH7ClqzCHIwE8HmSeaNRD+SmacmcB+oLWquBkAcZziC92c
usZdqelq6tQhlyjQDze2XcBJlaA1ngQZuzrxv4mysEmK+F2qImveRpEFT/2sdhLJSLiR7oj4h3zl
903HhxdqZZo5Nh9iFXqKW8iFtu4i8fvALg/x4XvcXvg93sSmoojBO6zor/NZRgru0IVrmlnG25pW
GW7k7pFUAq6pMqPOVgYxp6GJLblB+hRZr3Yd2hiFrfSuafdhwpTe0bolQXP3QfLZgSK8bgPjG942
G02Oyz/q5gOq7mA5I6E3x3uVDAeOSNEe8qq8AJdDUMTGahQnYkMRvy3xlxPx34Pj5/CptLVsWHYI
369rkjsZVLw9V6Ub92W9w6a/owZ3YxkmsJNw95pF1vAFf4uiyEz05zQh0oGA25IVPgKp9rG7qDbB
xWSYKjQ1BK3xq5xkNjg2f/LFeKkR0uTwJK5Dku2do3Rn2Z5sFgpbRi+VuPk5GcCdvbeiqnpt5lyX
ryrC0YczEWujiLVdcnHuokYp2yI/b5Y5PGWWwIhXPoDRWaynpTlE+Zfr73kMtG+CdILD4XXSaMDF
fVxrtuEJcjRlbFR299ylbwXoUPDSyxRjudXX5UKP3J7R4ohGdtpfJTblbniJ0l8Gz/RDWF7nUEd3
D2Q82xEpQAmK24pYHJy9o+ie73WG5LWLbl0AY0J9QdU8OS/V8TJSeEuNwNT6U/0VVEBi04utJvD/
W8WxQ42fnueFP1I1L+t77HyZwAuZ+1/XvoyWnbzw/RvZzubBsbPWo9/VqplzbUhSPj2yAyE0sqNZ
s+MFkAo6galkIf4FyC0E54atcPVFvGWrZBOzMnN02gJ3nZCAMWI3+UrzvZAIBK2czIgDJlQQBDIN
sNu0rxBLsDVJ8mAT6bduGqJ3VT/bl39UhnMpyKVSKYcD77dddlGKv4UfKHC1fdVwx0XAQxsOMtX1
opgd0JgsQ6vxGcdPCkA7Q4KHcqWb0np4hP/Jy4uQM5Ff7D4sFYvSzXNjC7Vx2ApozfnfIw7YiAeJ
mA7sbEjHHxlwX71+oaeCridfDNcW0sTlrAcs6OozSDzFxl6zTTxjyQtf6huCczsLqMILrfSqkbtX
2k6chA2uco5YLZHnIbYjl/NcUKJxYMGh+qN7azRmpa8qmfb3ZdTDXDLSBcXSI8sXixXowZwik5mR
nlhwmmtDD3AqvfQit7qmioTqulWLSukbEr84Goc+Gkx2i8Bu+GgVrTEspiOl2YjRA2SRZwr2JUPI
/YTFj+H8i/mLxVweLnzbWeKsHCcf+woa6DVWP35sJqJwgEJD3zKTzVnrc7rAsBJrsGadSYzkzZpv
PrlQlkcm5P+4DfZ+Zc0iTmM8b/euTXZfUWWyMazdPOH4AFW7aVTKC1DYrJ7d/jnWasFS0Qnk/fGg
V6hEQQ546ZGz4ENvj2shNqA/r1TJS6yW25dN8bhdevbB7zzJarkd4HM/48ye0dfHHk6PSCcIdL0T
o4Sq586YqYxrlFzQuQJxtQypJJl8LGN0Z9reasOMORcOvasze/kWytcl65alg3yBzcQbVVzRFnp0
5t1guxqS0y1hrwgom1Yulsbcjak2Z2Dcc6MtuQzV5vjgcBoN2FJ1ohdfJFiH+qInoE0vLOBoxQbx
XS+26N43Y9kaSlhydDjaRM6fgNtd6R/wbLvv9iIh/mGbIdsPcXqzZJjuwh+mb+TqDWT3cB7Z0hCN
vehl8sKkreTqOYvLE9P7w7iYVm6ATszXpQf6LMbZ+/f7Qenbic2I+yGIYmVzntLiZgXjMmlUJarf
7Ynx20AZ4IgI2KxFpOFAU9P39vEp+IYaYSuw8Si/6qSe+qYad2N9SQMuHOV4u8SQ2vPbuMv4G0cj
LMbq/hWcnKlRpLCyCuWECuqzd7CR+PD/wCZKniRfzseaQ+wEVlYRqbXGNp8k5/q6ZK6Cr5FRa3aj
0ii6e+HIb1EUe71HDj75O2fXUNIeuXZARHMvrn9CeyPKgRfrKpUYn9rlxg08zb0wdfOUw2YvHosx
JcYmi1zt1V4r4j3fBnFGtYIUgMUhTQV/Q4hC/T6+ptZqZunCZxrad7zn6t1+CY4o8SJhTHMHEZzI
i+xDZGJ0V9UMaF/NEukbkii1vtwCB2Dmo4Ba9yxCTGyrHxKBApOgvJkX/JOc8k7wY8NpI8M2d4KY
sRAZACl+r65U59/7dvN11wYcEPnDB1vAPrj8xnfCUOdjejWZyu5HDITZEuSKvYQPALLUQB4RZHSY
9obWZntWlZ9fb9rR9MoTlynNjcqyFZyMeFFv2E0tgGn43CDJpZWLtPbY7mMnrJRQMhymTSkHE3NO
3lyv4S63vihAM0V4pXJjev7VLUNYj9uJskJDcw6u8ovmJg2Lm0U6ZW1iJnFnxTb3FLU7UNF+WxIp
XEzKNaf0PcAIM02q29bnm/hNeh+mxlHwbMn/LQhrvEj1y7Wo/P+H/RL2z63Ml2pZEZAWzE7ognWz
LhXUwQyzaLEbi5gYo68AMQx7aDpmjqAWTEZHYz+Op7A8ylGLBpAiNWfLbeZfxb+Uji+1F8u8r01X
I/lidaprI5AfHJUn0KzrhF9NP/6MvH+7XFMFTU7u/Dm/+PRXYwXACYlLU6ory9I8YF3OqOJqGC0z
yqtPk1seOPlaOJUdoKCdtKp+DExJCdpLeZSa1vt7oGc+iRbe1RlO1JrtqOplixS1AI8MmN01Lslz
QJKt5Pv4NathLME1Uqhlu8GLbj1U+TQCwgel3cU0a8E3a8VfjXJsnyGKhpXUN/2tSYPC/2moLoC7
QCgsipaGrrNaT8AU9scb04A9HG/JoA+Gs57ScYFaPvwBPFGFfBha5whWWKUIIswo5WI3A7laS5tF
BYoYkCFNh0p1jcjmUWlLfK9+CkDwP+i8ab3xmQ4eatKITVe3jgap6qKjVsR3mUl0AYprJYYpzCB+
eZ/ZPDLhqkw3y3v8zFaEMXE+YrOdfJuJAfyRiT8OquyEsrJQsiJujTOhjsbfngHcdSOA87aj/Bk0
1p52m3y13UgU9gANUKXffZy+s9HHncb7DM4lbiYwetwX+ZLUzEJfFMGtPHzPuooZax7GpB2Sh2mm
IV7O+yLDyBu6nH4bgyJ7ZoTaIHuIFOdyz58UcLxtf8vRnAUG+H5xmnBt5xKvODGgmAGM9+bF180u
jx4uWNWYWa6fMb00NAiiQwCtbAL7P8jbopg3JOXVmm9LVoZ+joBpDR3hWVq0aPi94NrwTcbJWbCc
vdv/BAMOuO6Tjaf4cXND3ya2KTZDwM5q0HcHIg1bHDs5i0SIWNlCA2z/FW74qjumTmxDeimWIKFg
sReXIfoJXj1gYbc6l7S7wP/fMyjpuyDu2QTFG08sGiBDw2WAy0JYQcgNoefYcoPRkI4LTAYcpC+5
Pb0zlG4+eqHhQOuWQmU7PHWZDZmOkn9pP95+4V9WQ6DHc4QNEeFfo3lbsIoVdZ69mvCGVkH6UbCS
CFTLDyfZQyQKeMTg/yE+ngkmzBj/qmYHIElttUFzlGAE/OXCM8JkATU+dSH9jXyT4eHnWCls6PGy
bbZ9YOs7rJLBEHcErlAmW/13Ys6pHstbnjy1ugaVIfOxg+TsvF+I+uh06zjzq7cKtWQQytPuO8Ju
sDD/UlPgzfyM8ZdYJWGd32gekNcyUi9/OAvffKqEtJA98ngUgO3xVYz2wqZdHFz0f+hffio6u3Rj
EoftRZMIn/10quBY8F1aY5HojQuRNEq0Ssvml39YDlN4W4igi5rmypuMhwqqvMRuxoShp/fh+kfe
PDDDOZbwLWfMbNYTyUrp8cAsiddqxPrIl2FPiJDk2KdHbk0Xny7ADQzZ9OcJJtRSoTCX0/IgzBQU
AqHTrAo/3hnneHGvFgs7e1JPRg+yni5fQ+S0Y0gztiMQnomMEtetiXOZdXmeWXNAwBMoPT82Vdw1
78c3lwn1YckJed8Z66nFuwPlGOW0cMDi98uUj0TEvPoHinuMrYH/G+A+hcabdMGF4wTIpAL3K+ik
VNspBCvsdbvLgCbi+voK4gL1LIlgKXwP/ffnlrnt4TnZYtYjD/T0mgdWhy9P5xqJdRiw/dLQ9YQv
VhbbRa0RYTteQxqD0gGnzwzRi6iuXv6t3aJGQpG9QYdr8Cv0O5TSuM3KbfquOz2bNKBmecRf9kbL
e7Lnr1SyquqaGrcpxzpoR3Rx/HPkqKeML4Qrocum7a1/WEav+gRhYcvObTZWsfgDLxo4zYZvmkzu
7vj1+LJ5Jhm4CHFT/R0+isc1wtVs/yjeS0gecloV+ruN3wEwV0vzr4DIfy4pr3wXHqZT5s4rbgWN
Fi2rFm++0K5/HpEUEKfFKmWIAtu9HimM8rr+Y3/nA3vPfTVlbMz1Egt6HDa2DV6fvAyoNou1eJET
dqIzAteEE7Uio+hu6t6Sm4kNU+n1z54alL74ERO/may6juHK5MiZDCGYfjpFgqvflUNS+NfpN6fn
kY1SAMIu6g3GyGKicAbwgG7hZmlfzqe/q5i/++HK8nJ399ptBQ62KAY/ISNR/QeODU84jSXZ3RTd
N1UkIxP7hhppZc9pQVVuVy+pxgkuNlWkhcx/3MvyUxvlgp/rwNMULgyu8S1MWz02CsIZrQ/WWkDC
1fnEZFmbSA3qFJPC+zx4edajrBF5PufNKeGyLFc1ONPCvtqLhleRBNSqJjp8CYtcdNtH0D462lQ/
lN0k/AO3V0LU7ZQnhfb7WYhMgbFkqGEBsFECBe2vkE2iVcN6B0wtfAwNUJJXTqOTuoquv8CVICh/
ceAfq19dWTwbpnKkm+2F8Sc7ms+SaemCH3QjdJsw12uRSxtCfLv+uJLQgekbAQdM94stdmnslxm4
V4iL/HFYh9PJNusCpHMJR20zAgY3zj6odRV9MJxEHBPl6q7k0LWsV42yMwTPNv0n3Tpgd/BImq9L
5I5r1aTLzn/bZO1lr89WLHI8Awwwh45ro/VhknxNUfriN3wq5OSS7W30tKS1rgxsCKxHsX5sarxq
1KrhpvoGk5ii0IsKaj1hjbJM/ykruACAuVQauermsShcs8TkPp5gJsqZL9LQExp1FrPBzIvi0J4v
xoW3g7qF5pr+dVDEGRzajmXRdITpw4U0fIDbuD/pTF3abNLIHrW4cA0a1DrGad7A/o+x6LU1Iimx
BKz61JtS6HCELAwl1icIBuRsdWw8jZrmt0P6KsISX0k4EVXUbeH1qc78jjmQg9BtO4m6aIcG7chh
a4aQdSVTbYmLNNAEf76gthso1Djzmp26eBCAX429ePs3bIAKXTFhcxfOQBq2ZezZ9+mxzbnjIUNG
OX6iNYw9yI1+T4h9ZyLABNmTrBxPOi6uEx5G83KLJjDqMAjFMR2qcyp4FO9u7VPPZi6Pqi64GDr9
qkt/mzKuowC8r0R2c7N2jDGz2Kc5t6nxD/6k/QfFSDV/I6QnwPpvvyDaHoYLCeXqp4H7+RieEpnh
CspR5mluMkKrxTywO5CFtTwdGhJJDmZnGpMoJuiCeAbTozurWdLjmBO2fZ8TgR+R19GHz2v21apU
Qkk7kMJnDaY5oFfwBdvg0xU35/4CjEtFFtsBIfC+f5kOCS90Qed3uBHx3mXxZV89Gfqx9zCC7BTw
vjLjfdFCEmxo7/R5VOD5PGRf3s8sE8qRHtb8BwWf87jKA5iu/lIw6pmKjQ8eVxTeLnxExuZGG5SJ
wNLnUSGHWjxKnSqVMwvqJoKc4uFYhQZrVA/yQI+t5AacO3k30nXTuhPJ2X++G+KueZAXo18Gja/b
av31ww2gTg530JCYF0/NaSS8TPXJKocf0XpQPcYTN7KgQk6YNQlDVDiKNlUnlxMciy1WXeoC0dRY
+MwT0+TKiaKQYSqonhJItayFbkh85AVM3uTuAXuI7a0qYQatcpLaGY/assZF57kW+L7xUPYu93wS
mrRky2Gxwe4KrdTeEblTVhvPH7Hhj5mY12iu1aPbUw6CvY5bY1CtaLB2m39zGX6wojQESUZEpdEu
AfHrTNRqj2f0sukbcUpZxZlJbUn46rYflS3T8BtofnseHhVAqm5/xmK7VNrrO2Sm+w1PBQCktC9B
CnOOIwLe/9By8SVeJocM/60ReQQ+1sVzqDod5voH7Pz4O7LBzBmpdi/A8ZeAylr9d+mvGkeeMgeY
8SRD2/R526IRl/O4x5AE6gfBhLBHr17Vscf3YeZKleeHukXwSW/t/r7U1QFtf2TOmX1JDnWk5XLA
wJTvoL25dfQ7pAuI8tS1FaVLBjwYKYzDtx8gC7M5V7RllX1GMUuRzyAWaM+guzMVH9GZrko6e9Hy
H8LOLJ9ZWh+qSPvCOlUaXupuVSd5XU4xn6alghDhbrfch6iswHNfeVTvL0h9IJI/62vNrQv6ahrh
YISZ0r8AUnpLdNi2K9sa2HXz0FQ0kYZo8uVavxNDkU2MSsjQIvQdhYgscFQdyBsV4F2FC1D5/477
6VJROgq35dEhfXCn38UGNbqC3jwUfKWZZWf97waJiuAcwKy4lZEy7yha68weh7NPGe4Ptz8zecBU
042WzmJaeMVnxjdgmVLYg1PXCW8kwYnfsZdtnwIgyTdsRJwzJt37SnMUw4eB+GnVwcVwSJhgzXXV
f6sMso+YBfeYHg/gLYhQ7SSbmcz8n+gRXb66U1truO3LIrTRI2IvUnlzGDQuXFXNdEEdKobR0/pM
L4uKF6pL8AYCc9+sFCPLR9MStM5nc8amEUJbtdpKv4SHSMKPxbSSMrb32lameJzoQHgG1jEpAu5y
RCIDLIjQxre/G2BZFZUrmlWLgNSuwnT1IVAyUukwdr2sGIe1FyTGlG+ARc1z0v+xGYQqT6x5uosa
r6MrctQTGNrZjXuGp/j+qzNgrsnWn8j2gCdrdQocugOVjKoazLB8s4eo0FYhZhzp3P1I7Z2gQh3F
pKqG5+E6BXTQEbRjyzBiM1nk79qqqZdAQkwmFdAaVmKwhhPOVfR4FiG5mioVxFEARi2DKZh0vf1K
Nc7XlyhcSR5i1DZcRZwrGaWu4x+2GFyXZDV4gx2L7BFnwJpmRxFmajpDgBGzFtYu5h+fzzWWaP5D
3tfAoSVN5UfJDNvpsoNrafmCUPsJe5JX0nOZ8VuJtpa+ZZlNNu1Q6IF9j6wCO+3qCX3kix1KX7wP
JAMDNpbBdtDQ5YGRU+IkWIa29PaWNOwzPTYp0OCfsiwdzlV6fV1FgXmLr89qaCpcMl/071CzcKEt
4NIKXVgCxTstcwHL5wmc5oBFSPUjpp8dUbz74QbgZrzqoWhwnYPtADArBktqPG1h42c1nVjf9qTQ
Ku+YtzeiDodR9NOP87MIs9eHlRc86PoGhYio5vluqpdOvUy40nGUznMdNYGqp4L+oaa+tpRW8/9e
IrP9jW4+2V6IpF87zBb2HxgRyc4GJe0LjrUwkukM2Oy7ql1+SWMhA1HoH8ENSV0gFKPKID3Pwfoi
TyFSGcg52KqsqeHSZS3U8Qv+KX+RgY2/dyAU3JOrooIvuRib9OMgScaKeFYUuuIcGmETFw4HEiZu
jsaoO6CyWPDL8cO7v7hatjfcemX6Q/9fa9NEBxgR2/qocnK60ey4mjWzPgW20HUeu7O5qpY145nP
iLoFgQVP0BlyUu7zdpBl3HrgZm1QdaR83Fx4ouSrA1huk6zCOafXqL06j3LuvurDKpyTNsRPWIVl
EGkp/gf3cCMreZNxqOzrKd4lUGXWaiYyhkurkiSPWOXK/e90dxznxGWwmNN2OGvVcZCCGnKJWS/p
xXG3FLciUdBLxvwPduQr3ae2rQYCgOpoZ9Xy8J/WWNHVavoihyRHRw48SGtBNeohgh2WSpp122mf
Iy/ugi3Qh7pgeKFRmcukqPbxzJk+TCPq03cC7wzhdZum4+f07a3cHxWX5qfk6QsCliQh7N7xcItK
fwr4rW4QpFsTCYh26qnFgrPvcU5utNolNiKZ6cSo+FNR3RF9CNIloQq1iT95OsZ2yP5zJt1EImRx
ugnN2L44Lje+wxuQZnCVQRn7fhoBUBUW19INyZY/2VPTIInqfxnaFgB7KDwS5T9fN3re4bHV7Q1v
sHbEJ/0panlYIOqSoxnvRLlU2MxxuIZ3ZhcP4GSIjJHnU9Sr4aFRuFrj+IM6Z8JTUdrEYpN1O0+Z
nvqPlGKixFvya3iR/5EE8RWUle8LoGvoU1fX1VtblrguDSD/CHjEhqtbtilDBUx1eV+KbM62ZbNW
xMOWvtPNhibqoA49eM9MklILV09YM63vG681/yhDMgKHaMnPMeyp0foYtg8aQy6ahGdVPuB4GL1d
DTFVGJL+AooZcZaPk3oWnQLc+c6vlUnhhPeZnGl8zwArYRcgKhg7sj41J3gwPYD04+Giv2L8o9hW
LxcnStwkKU/EeYcPqZdp51zG1lHbVh6KmNIWCF5hmk+xF24ryCI5P3BLNLgHbJsfMMsdN1+46xQG
okFafQW+7Dx4i74F8vaje5EzMSEnr8NRo+DcSeZzz7Ijt9JcZvH4mt/DjDsSMGefi0yBJtgHGdfW
2CFZHxpMXrEtLCqkgGFFHEQ4jQL+ZJbMATLZZ0GorH939W0n3JVSNBdUijT/5qqrWdx87Iu58hzh
lqz84D3aXlNnIQbilDUiQLUlYc6QLBt8wuhEtmEBcpFwRDDJrUFelctQI3DTl91Da0YTgB+HDuF0
agT56QRfJSvFqQGjnNZ5NDjR34mlSIwqBipYVbufK7XXBG6r7gDdGt7UXQWK3aUvJ0cgaYZbCAG1
FkrcX2Ki5hYpSZDLwgRoL8uDHu97fD5p6Sw1bm8p948aBMmeltgQzhQ+FqmtOzx1A0zCc4kryAKJ
uE+kfV6g6y2qzOyXXrdYWlT9Fv+4cxgRKTgVg/lzoKc17CU+zLJfX199gaOJozIhf0JH137Bqae0
YMg/bFwyUfbKSFynuS+0aBBSaT3BvHAluSC8BDGZ4FmrvE5fYW4gUwqiXpiUOJRRhjDmkXN/6K+b
h/infJtfgCazzD+dn+iAAHsbL7komzYjInTt+v4ItBUQvwoVl7xUwOkSSeSw3nRUOh3ACDq5VvJr
9NMhJoKsEJZxR8QMNy+FTfdI3d+fNz72p4ZgEKyXm9KPjk0tuScLSE4GHna3Urlljq8KZLUjGtK3
JWY1fssJriOgTlJU2Gu2K1kB80u8LvJ1CDarOt+KqzeDsMyY+bKzm8NCEohfmjUp0WYkpDMhN3gU
9s8UI3nVAMkyQyDn03LAX7WF5TF1qi0X7kakH9oPcTJsmgRhLEoPyiNa6rVfZOiGA2xHEKTs224g
mEVTBjg18l+YcASizMro3X1PlVL+Be6YO7edHdptW1GmjB1+1MXOqnulI0kRwgKcA83svxfT4tSn
H6tBWnuNGS1M/JPfvQ7iehvMQCY9LjVVVI4eE7H0p72ucLUL6YD3R77BchDlclbvDnS4E+LkEzhU
bv3svNEfRNdkwmBY3BpIMVHdMVe79zLAsGmvtRrpSxKL/WeTlEZOEYvG/JwJpujq0Jhi+PLU+/6e
JSyYhzN7OyBB+8PN+gizpUPtoUp8GdgwlvhF1iWP4Wd9L0XaxT7dKMNsS6yXdBk7jPP6UbabgJ6Q
YCJp5zadS05fG3DL/g9C/0P9MYlwDeJPotI2Teh32c+LO72Ts9fzRfrj+fpytSH8r+VknG7+24iB
PVPUe9X7JkFUxLgQE1YATn3BpsWhmURQqn/qzzFW52Ts4pTc65rvhVR2l369bLaYeoWLh8kcrxTi
vDU+KNh6NXJzWVJhLvcGJMguaEATqcRnonBiY3J1+C/LmXFB/IA+QhfsaDy20ABYcsX22toSsoXB
b3XU5EaKxGgkHgc1PrDkB2FmgYsvrprkJHFjR8O4zN8its98m8NUXjWOZFrbeApviY7g/te0NqmZ
qr4egH916xOG11o7/eIhzdKLn24/L3DLvHUsp3KGhO2z2Yjp2F/n5Fj/e9rxAxycEI7+6/G6EvZC
xfByvVTd5esH46BAZf9vFLrvJi02udTi7iRpHQoeVQB+4gATnmhCpZYE8GvKiSxn9giUaceUCNJf
HKhnpT6CKggEPdwZLBf/yH3cop3+vTiTmVvC4Qsv5oqMd6cYZUOb9mjSPvrK3Fxj1bT92cIylES9
0FoDi/qayNZ2/CkaFsA8C4W9uNZrx3LNY780U6BESxjj3hW/RbNkwoM9KacowWYqppmnaFtfqeh3
XWq3EZmkFC7IYxcTl3PoNQE181rPqLjc+SIYXF/TLmg/y3qtPeptwh5xcEugt1DUrcldf2ffives
X8XAikII1/Lg41Ay1colK6o/HTt7QLBx/qdNfgTgyAcjuAeAAH1ZkVs9W5C36oEUpZNHU0nZJ0n7
XmfKCzQwHFYA1yexk+Ek20JvcW6sappOpG8nNeHVJPSKVaH5J/roHGKVb9UHBD0OdP5KMtvZaSBK
kubkZjeoIqEAej2OnsZy0qqnfXlneJJgnXYHmM3mrUAdHJOKwNau4hBdYRNZkF41U8z7c1piDiVr
Ys5WLuwGbGV5i+1igl9zQtc8ANTkj59ltpaiwWsxpgSUfOihRfueClMAVm/ZAIo96GZLdIArbyU5
E+AUmrfJt55mNa19M9eBNBBgwUGNtC4LAq9ugSuyruT5btdF6hZ2I5GNq7Vq/WUAjRTGT6g9NUwk
9vej1OI4E0bPSr5klFGvZJacfdqwjbrFkaiVnhxmwO91kHXVcWV511qTtLyA0PMZ1KVMhe7wVTB6
FzPMSN7PvHNm+QnW4DQBCLYU8d5BiAfxJM111LC0o6MTP7BvvH4XuZoo2lJzDd88EX4H9QQS/W5O
Kd5ANRjn3IA+C495LqocUjPhLYAKaYeNWZe7KFTq2w5L6ZNzibvRNNznjpuWD7TVOK6XuxV1z9gk
k5P6sbWB47chEfRNN5nk3ER1wOvOCP9nH6iWUd8a6/yVgXUSZr46GnZjE4v2lISdJUKfEkXxxUid
Ryp4zyd5gAecpYsFmC8dqPvsVX+wPdsYvFaKJFC1otDx5mQqdGfVHFB4cvMpdMeSw0NPnLKON8aw
Vxv/f7cMbXQWcqDLzdCH7wlxZCsR3O3pIhlHC5iohXWj7SDlzvqu+PBNLh5TRzYWQe8iutdxmD3q
GqwZAByQwbavo38nJkOH1JVvvqI+yoo1Pfl0fKoPuHXQtGMmZtrT+3pVIGOe9hZQKCy5qE4zT9PN
mrxBJEh19uHXmOmtmlCiftDIcjpngHGXM0/4CDQgU78PsQQ7gMOJIYxZOJ66ejkF02A3CFFX4/JD
x8/vKY+oerqI8PQovKj/yeEZghSeZqc87O33JGz6DMzgGwdsuvqEn2PXJiYJzR1Nu6ieo3lFG8d8
EgR5/ZNtgouIk0JbaHrIaZeQdB1LUqMuj+7rPGU8G8wk2vOs1j6t2QTfI4YlzkToI8n1nwXiwKtq
0MZKHX6BbU/geFrthazUCVccjj2aSxCe/v80LeJ6ug9CF7EEtIQrUsEOD5DhWhvYogH/x9alF2aY
WsV4KYboeAyuCbgKZszE88rsdb+rE/bnsDFsavlj0/tMwf6L8eCMPFMx0JDs8/sMRKIaFO9RtsaP
uVFPgGRXpKNnt6rOvYeuR1X7UZ3OZfnQe2KE/DJufACl21XehEuEEHXeou2AOxpcIWEEeAwyvE3M
ctrV5fwp42cdor/V9gYEhyvVssFPH1j6BK2sNc2/6pFz+5mXi09boejd6GBhG64X/J+x3VuP08R0
h0don32R9we1uTTPDtkaODR/NWyRSySuB7P3cvzLXl29qNlc+6kix66fFu6rtOWIy8MlBagOt3rB
K8kNhyFCAe3DEMe4Ro8LIaXN+EWuB6qBmvWmNY6x5rakKkW50icaIZHacdnK2kQD/GQVytNsvmZu
s/IMk3KjoEWUs66UNe0gHszDsEANtglLNQxpgwTRbDTotiZN+NzocPBAaQQTdPQXjnZQ4L1v559G
hI74oecvZE1m2qBCn1TzVN7CR8MhBFH0bQmfPseYYmuDBm91/1OH3TBvTdrL9q93ahrCcv1wK8c5
FkWVJmyOpSltuCXO0mGcOsVsHU+WhEheVBmk2g446DCZK2igR7nSATOSA3SwqZtEVfQb76zFhS9H
FOs0mr1AWZ1tOcfS5daojcPRERi9ewJXKcD+MdPR0ZqoSAkYTNcyR6gItK4cYHeYaPfcCMURyeha
3GG6TBa3sV0rgWIWcsdpXu5i1xHIb9i/s2ki82FdqrQPjnt7LEPJvcwqUA17xc179YASncXSaNse
wx4lEWMrJQF+36eG0iLEXKX/oceYKB9gvrzHC2MLCiBILH4ct/iLw4YjKy9ERowGIqLsCTOu2wzh
NpeQENnO/ubye7OgE/+g/GiabqPjj+JQpCY5tX6JDP2r+f4Kmg+gEv34nb3IVNMb8aDARdAB+nst
L3JnwCzFE5Dwe58xKwP27SZCOlALMABihcq6XvNrweMaapgiOq/bE6n1D5fX3Ejni+nITUQEtwQt
1nSljR9swL1dBxCR0QNu5SkL3sh65ZhHYV0M2t+TMoXM8VvIbd4Ld/OSywLcXfrIAd1VFbZdglSf
m/1Eppk44RRf1+/Wf0YWTe/WE84qC9PAK5/rgFcCMC+EZbu6j6DA7kYfYJhz+bSV6fyrMBN227La
qB3wagzTpbwO492qDKXDy0jwHsJ/PRnllZAMwX3eiPP38rD4A7+HWvyDulAnS2vWxM8c0lAoXStC
MEy8i4giv1nKyg0u8GYRqLrYhJoUfRj14djiCZSjY0Kj7z0eVG9uIaTFSwdw6L250rprfz6Ee/LU
U0za3Txh1bOU9GocSIcUULLld+OA/aSc8+4BTMxCto9JHLA8APeibOaqDkJPL+x19CI/ZHrEyE8F
hjvxQOiTVE3wtXHM7Y4Bs0rXjgCW6NvyTparIys5U7tQ9qxqT//p/MUeXV2XNwD+0DTPK74Y9rqx
IpO3iLS/hcsydyegpfSvTt7EoTYdTMf/9Aj0dXAocFMZ4qRLVqiKsfm8tcWncCY6HKFwznKkX0gf
jeYlbGOCt96QJPt2cT0y7tzOj7w6HziMmZjOwN76l6xXdHuzvp3NWLjbJM8hvqxX5EV647Iq9Lil
HR25TPDTlVgE0OjrCaE9grZFtIUeYK0w8T11xiG34edxFWFvuXvFIj1P+02zTKtZ7LIDkaq21wme
9IAOll/3BBnG7pug4DLNi4+/Eo7Gt8QRX1OfZ8dO4Ar+6YjM6YElPWxkSrw9+tdzX9y2bj/5oYMy
5dBQQhbasvvTb4mu3a23gWXKyOw3kTX9SKD3UH/WR4ZM7NNeRbNsRFyaWCY8tjAk8thqXQVOxI6i
MnRmLl0Iw42ksn3TZb6E6mxp3DYQLbCSVwrU4/CmTt2Y2eJpVTMg81GGMLhQ6WjAgUREKVz45IDB
4KQ4wLUETbDRz+5+IancQ90nBYoCdsU4o2DOAJPAoFLJR/2Y3D85Tq5uHFJisxEfdeG5J7i3pdnq
/7UoeQC6UyFNbGPumGkiPkRyg1YsX8d6bY06CRUndL1NaeJgOOS7QUODH/4Z4vhLByeNQK4tT4ZH
AhMLJcfj1TND0nu4FqNQkkb3iQm96b5RN7NMMsJ+WtGZFthnSGQbvz222D0Zm6YmVNIQZQVwUyYW
85cXbPRsiDUh5pN9SmlKq96O9OE4QFGWLjNIviR+ZABJsmq279wJn6HzE2cBtRJiYHsxOtw9ml5O
9u9x+Glz0okdpm7u9aI9/HKB2yLkiSB9Ua8jsp+nthwS7Smyj8aaNqYmsrInmErnVXJuxHergGKf
7KvBBaueu5T2HGsBRcUnBP6CMZD/3DXfmke18ThFxpIzcNjhDHk2w1pDAYqpttJzaZWxXbpP03DS
dJmZ2BsXYSReLyZ3XnyjussvCIh9IZPX+9cUhjOKLch53xmyr6aHQ5ZBiw8sgd30T104WMjJFcZ7
JnhICJnAHL2OJZa5HgMedomZYQXCvUEuZy/fl6tg6ONTxJODduXleTKkwj2q+nPwLJb2L3HUTEGw
IRE0wAwohGtTk8Mp3tcxc+upIM5kwq+6I0L6bb9dyC3fSjvEOttzetGRhYBB9C6TFrPNQeHl5iWO
hGCzqKW39OC2Ip9XeZVOWGy9ZafIZGmyiPy7f8vyhM6phD4j2uEqMvbktT8hTUrm4fY35QI/zQ2P
RHVle/mgW+p7U/7YOTjZf1bdWOuRWfiAQdtCZMN5VNvy5xaDpz5iWqlPvIE8B0V/3QRwX0CO2/9a
Owm6T6wwN+dhAXGxt0Ws19K+fLQ9cANX/9Cz4HnNcwVENtuzHPrWsiUUCcNvd89OrsHHuLEd4+K8
ReztQgR5P+c1ZM+YbY3YnUHrRb8vT8SyFOpaw0owKMqjRT8v9lpYAW/vNDCzGSe1Tn9Q0jc1owkO
iK7YS4oQlcKKkOAiP2GSTAqZ9kdkBvMJOEzlKG2Kf7lNp7oO3dlbyJp2StWBXTs/gwI5aesLCLSI
mTzWbAPxJYTxXmVygx5F/goB2xjB+H2XVdf/QzPhH+YIFhDx4Cx9c6nXewOs9guC+l4RfbiLqnM3
j1NtjQtjghMEv/PRPj9Q7vhAzbJ5ezlZ9UkWe9e6zNDSSXN+6tYMPTZtYDv3kOOzChuOC40/RT+v
qxwFsmvxBpTc9k02HuI5CzAStYTa0EpR9N+kEFKHaV3cghBCVsIb8IeLZf7ZgBkQWMdiLA6z2734
Y5cPk+VyM8a+Zgnp/u4aQ4aQ79XEqJFhMV7bgpmdSnGz4rU+M2xb16hdXEGKluv8Suets5S3jNNc
LcVcc0LpK/SNfMnTamvtgdZSp6KUt5WBN1JycLC9xMUvt1Fwk9lhkthph4QgI79H/U0Q2KvdXK2v
5OP+tsQAUF9IltaVaug3GPDpynoZseo8c8E50cP7iLjJDtVRvA6uKpNC/pn30py39MYaW7PUVMNp
PlL0UdQNhwER+eEQ2eESYJ+Tim1nqSconbQVPBgHsIsFEZ/3DL++eB7b++qVfW8pSFY9Jn4ol19H
lkm6AiE8NFWfCFlI2aIbOFLaOWck6fn6KPFJUBJ6/8SQ7EPQOI6qEJyRfV45yiaE2Ye7MvzL4d09
k++l3cpXPx5rMVJ5f6eGZWpbiQCP+vE6dmWxpg/dmBUJVjK3In6pI0jTk/Z7Z8RKvraNFYRVmF44
dhP4NLb0qTMYRQFl4CDwvDpqMYDWKoMidj3x2OYVhYJF8Q+VZrLTg0ZpjypRGrzoJRrIK7R5y7Lo
ngSq3UQiRDUZQPFGWsFMB3TPukhprOaUoIsOEUzhvsVLNy58ViKLeiUVxsVDCE6cxNBGGZBeenSL
oTT7bk+dnTIsZVDDjpT7iqEPFdXgdutmJn22XO0uSh6Uf22Dh2uA1/NfEOno8cB3hNF5GP3/qw0E
jXw9dhjOKY+Ty8YcpKdH2ABjfdzQ692qbR5GspLPnPpMVVhEAT4woARl43yabbEY0M0ILcm2igfd
2jDyo9DcrwT5y5bOmdQalC2JSARBdItkwYZX/wHFdm9HIx+oF1/Suovuoxg1Z64sjekFYvZS063p
ElE2O2Pr1NdfMXR3IxsOyfFKrR9glNGpDVf6kFYXQzjpu4+du8gqn21NJM7c/JTvON9zTMuKk8GL
li3lEAxBwW286GAjUME0bEAtOJqLxyy/z9NdWHv+d37222fT7AwtKiWGytM1fEnsINfjTseg4eMZ
cIU2BtfUSB8bCQFwME6wCjjBCxw96MlIRolrVhz/CAlpzB9OiEfCMErp7hDHluRhnA/aDkY1bgJn
lHtfHTyMBbuQBmgvtMrphj7hZxui47rOTIgAKoVlsh0QSNO/+EtcOHLIkMFBJuXzljOo0HXV/KNt
IySoDVSnBcOeIOM9/sVuzcoWME/HGrA4nicopLoZGyRBoRmv3NnHK08uJlD2mPRr2MKljI+fPHSF
XS40SqOyDg2sch2jDS5oE9ntEBvJ9d2Otq0tiZVvLcypLR7skGPvILCkC9TZ8eX90dAJON2XNeHT
vZUONEeWYsEutg/3Ce0QmFWdS53L9pn/OD6dCfpKpJ/MJWiaL8cRMkkifpCowKVTOlLpkc2xyktR
N/sOWe127QBadzfwA50TpTQdeqPaVKI04EdSk6XKvPieOr6EKVCvMH4/Ato9wEjz6BNqBhMYogIP
JdEF2+dxUt6Fn4xg01o4XZuJIAt0mmU0VqoK7EblO4Fc7lNNeAjQitTNcMpUetQN/0KmRLBOw8Nm
wnYgxKE3TWNuJLFr6fLp9axXdE2VoFJ8E26Ev9aV/7ElYz2HIsClbU+mwHXM3lfLkAnDXEpD4UOG
Ojvl7sxsmlKfDOz4FFE2KDabJu8gsVU7hyu/M+OzERy1a21jwA8Qw0NmfnSHfQnX52S3LS5IEF9y
89g/CL7Jo4Kl/6lR03AtY3lsSOjyJnOqRxI0H64bfxIixqzTDCaAEwj6F94T8nTyl1z4SocL/tCf
1f+YcckaDDr7aDil2VHr9cmQAfEE8OnAzkLXfC7smFAm0atGVVBmGF64xxNyIqEPR6sLBc+tJYGD
spUjQT4pJq6wx0Ay+wYuhrZCDjlN7pFS3ih9nByE6HgSv0IfOdJ8Toy9jA+odBD63wE3m1i11rfI
dk2assUKa0B7XQZNREg0xnWC3wx8GLU+n6voBhzrvuaJFJLnhF+09xmI/6mO6H614e3/2If9si65
nxol7FGvnmT+MDaEMlK2pjO8CSDwviDta94E6RlhZhIBpsod02D4KBcfGBADj6lMapW48CQOQIR8
bTQbWe7K6yrmq59X1rfQ+A4m4kWGqay4cUMrCEmSgUZRuxwbkiVugH3ZzLFTzfqfoPc6tfVDKhmD
W1seJ1lvXsNVD9rZHcQzGnfoC/8kC8PdN9u8i+L2dXYixa0csqUM/PKtCrESBSF55M3hGLV8KqPS
YMUMjeFpS2jVOcHSlltyIaHm5Z2lPRiOvYCXbUH8OS7HvmEbBlXZOqPfVNmChZs8S6Z0T2fd30gM
i0w6TP+JJNIn4eD83UKqhVHkTL+XdRUkOghsbyxuUz3y5YRB/MvXSivE31xcRiZG91WnZ1/hCvns
HSSPIxGdVoV37GtvSy76GKSeloD2EliOaAajoL4sFMB6P8ADDfGEm9Cp3YfNgbNLTFxP56eUASeZ
4vpe6p+pls9oeoq0O18aFHcMx5idIQ4ktPKgi/y9o4LdqBRsMXR588RWoP1eZDzPDldwBVzp78Gk
z9oQn+AblLPHFqqL0/1E0ghW+zbf6KgYm0bcwwHeQkLuysE/FVSseUckE63APfqUfLJ6o5XqZM8o
J/h0BmEcTwF431l7oRQkygBr5C0Q099WVl81HFNEyugutvSLSGVhMWZcRX4IdLVS+E0h526CVTUy
0j7X7ARtUfCAI6Yaa78KvSiM28GskhMSAaWaTmDD3P0GIZ2wjfWHRoyYA7sFcYwF6MrczXhqjc8/
/Hing92w4ymOJ4dcr87zCRb1+R4xyVg2kcCI1pWqX0Oi8ro5c99CS/vOIBOrvSXiS2E+XIekZZdJ
FLlOmHa74PLbaAMsBMj6EoEJALqxgKvRaiD/E0aWS9XnmrRSDEjYTKcQTGI3MpokNZ4DoN4Olp1b
jeaMxiWELuKov84hCNmdqfsAwoY+YZ2tEoCXMk1XJq2LuKhZ1EVV+Ik5lRO9q0GuXzzw3oB+ZHmH
LBmLkQXFGxFqkMZV7kFwI1bF3ERamROBZi21ISGRB6wa64DRZ36U7knPEz7YUTr46i5Zaa+zFkJq
BK/9JG8ewlCEsFZmJGy4feTnBCl+RvQ1Y1mRGKzGN+0JtPdtiHXOTbeCb3QI6e1Mh3RVhT9l+FxI
9fg/CcRpaVRnFeJS5Gm+w/LyUGK+S81KkXgReOgz2UK2F/aRMYGl6wN3OyZPdYgrTPwIIWjX2iHZ
q37in1qwvf5TlJ1kuRbxvnMPUkSOw03wuwVAypO1uknILfOP/Sis4FOB4YLv2NlEN64S7/d8APwm
l9Ekclslgf5Y/7+jetItpSOSmfupoeDqcwBsosmXl/TL+y8NS/KslbNv4zy03qGtPUGbo/3obmAP
Zs616hcu8z/CHpN3b+ylsFJuR+x1qSzAghlQhjouOStbm5lnLxdFdo7H90CbfcOBjHBk60w8MCpA
4lqybbfATvaCKjGF/3X8T9PaJ1X8R6eMRduE0rmNyrEQaMwaBIG1/4sBXQJzhjYXUHqqrsINJTmm
t4qY9CQE4GdLqeVOjsesdXvz0W4g330e+eiP+K9I2yg63imZZtWK7f9FmL6vpIvJJvTQMu/FeVcB
aCWJKkrwsL+xb56rmR2rTE+5kh8GLgK6wC/bl07NfzpEEr7W+g2FFBIebgfORz3yOUfXgP8IcSQ7
x2s6qyGajoJbskwMAGAMcVl34YtVeb1KzIMD69fVkjrnTSGDfiYuBGbPyKevhj3DMND3XJbOw2d5
hcsoof3OqnmicscyAJWYVWM9SSV90zMYQH7scoD5+zU/NCJJngT0ArZPKEeFTvoCe2/LroRjTFtF
1tPh1ixzOMvGYTuLic/FEth7PXNKSzRSueJrH96ovUflIcUf1/Bbk4MC2niCllmVNA9tAUV/BL92
bYseS1GFAP+upItR5uLvdTjQVZ5Zy/gFpA6srRMLdPCxE5THDYfwlpa+Rt3RMTWmdvYwGG8CPP4B
qbhTjU4EI+pDDcbezEctiGqkB11kZE2o9uY+VV5DGjUnYFJDAs0ywI91A1Typm3J9xCHngqO9Vx0
xUE/hJIToxhup8sZ4DHa+KcKaqnamhthO3Q+RcCXQd7TtnuXoYCxWf7cav99xmA9RSOT7iN4vzO6
Xl4zve5gSIYKnzCFKleKHvm33uULGUsvWg26i1OgPNqXEG6Apz6jpeIjZiloGgIj6aXhplNFGrg3
YZz9B8XneMGAroJJAR3mrQjSOqCOoXkZ0ynnA2uLToblNdyvlBTrfCP7xU+8hOZMB7rfPEiYtmN0
FJjoRv5NBgqyBevqVyjX2s7GotYPeDDCQSWsrNa041mwVDehT8GlbpHQX3Zdz0ervUpKRdjKAezt
Wbu69zB+/+gOjDN8DySrFYxdTEu1sQfmGNMJWQpUNJUxq6PWgKC4Uq89q+euww4JMUc73xdGJ9S9
4mcJG3yowrsIfOX8OQ5oqWKMoNrOvtFgRUdxcy0GDnu4ev3Jq2PGvCK9JZH45KNylEGwX8c+xJsV
CAQTPLM14igT4WlidL+yURq0sQ2PSlZO/dWkzVosIFk3TxfLqXxkY29SyOxlTYAuKZCQnYBkBcbK
tXLigtM+7omo9iqZFCccye8qd9lYiN2ONGgpLAHr8UCfiPS3Ae95oZ2a4vHWtCPK/Za+a26cbeZn
KU4adt3YYR4lVZasVlwMqiv6R/buX9RlkFNCrtW9UQ804fPpUz7xlHR+XlnaqaOEKSYgq2oC3H5/
xoTgMzowgHNLJVPfmn87n7sp7MPkh5MWBSodB/IzUqcEGpaAVj/tXTPNeTVBiI4J4IQuoXACqAw6
YS7UavqPvHBtYw8OZmny3m5GxVzAUL+3cIHQUzbbQzTqa9Ic1cxPqgIIF85QpTPe6o+VB5Lqsr0M
uatyiKK87ZgWvmN3ysqVlX/9Gws4uoKkYd/Syk6vQp/xWy1yYsxQp+t9D967P+AMjYPyQw7Bj90g
vIvOKWduN1/sgHkDkoCXU3w36Ma9/I7LXwjSBVxmzrB4NWrZNRqJ/JVtnG3L5OSB6Sf45R6GlSwQ
uMQe4MUecitxFzFfGUTxW1jgCfG9IKUxmVDWq3d79ggLf5e2G8wjfO2J1KCIrFQt5hxMVlyZ69QO
X60SCtZvWDMRJxBCKANJrZmmZbGFsRikDRTkzFwHCGsgdFq0RQibUILMFQhfrClwoH4HAKJqHsQj
AlvxDke7sDBphpto77XegiOKnj1MULq3y3xK5kZAu1F2iiwbG7F9ugHdruPgoSM2nD/MuFXmuA6t
Y+fZf3EHKFHSoav0bab9j1EcMMb2kE7nD+6D7qzyDv2HGcP4C8Xlz8J7AM2DRu12gujlPkDLU/H2
AG8ePl/MYrrEQbFQ80eqGU2gw4XyNMAlzDKTqM44VatwMtMljwLktHkQ3ZnrqR0PpLjBWcGOm/TT
cg9Yd7H+6eQO2WFmCpJPNUuTODRmwDvzYNQOEsqTBzWBU2bfhwZ1IZ6pMp6bmEuE9zex7/s+Nh1/
YDcNgIrluPCgis/j8ejk0jJQuJ8t97e7b8t5dXVGntPiyICt029cBnUWdP90gJEnWF3FyEUYBZgx
4/wdZdPAxXoo8MXPbec4VsUU6DJJ2Us2rzJwX/cF69xeLbdqJ6MJxe3ozj/kcpv8mYWUvYW0fZzm
8tvFfQf1TBOhGe1JJ6j+rTGBk7dftxsUIgIFLPWIBWlqxCedyxfKTGq8cy0kXNzdgCwPUfctNOey
HwqqEIbvOEztXTNUIOj7xTehCpnP+scq8Mluo2HivhtATsvWPmJBXvot1KKqzOInTf9TUHiWWzb/
Vt2uFynImIxFrNZxKKmQ8X0WGBE6OjTn5xrguLXPW9LlTSVCe1nOJV+SPLh5z0DZzDK/pvQGHLu3
/AlnSzG97fFGhf3Pd3m/hk6OPaTtsa37cb1j9bcPxi3avXSi5cQXfeK9dcKdMdaMtQtZClAyctI7
YuV1sYlLnxvoRWZMPetwgxNv2zq89Xgo9LJJSCaKNNkKza/psE1YexUCShfZRwia/MgZxqu+c+rc
2FnT1yvaeuEjZdpT5CqLQfUt588yZO8Qz2PSM0zeil7y5ru0DKYt+MZsLfprKJnsjoDlWpTymbZG
iMKwDqpxMuuhUQmfCUVGKsIHt6yoc/cneJs/xpaYTt8M+TaP6GDwk8IwMZCaf6H8HZDbcD1Or5ts
dBQl80mEGTpwAa+rVqA+HPo46/6V5ptiqDJ/i2p/91eTdB+man2RVZtk4ZntcYnNhMfoDNRIX286
juCPcjrXCHEAkewfBS2tP+vZuKn4+LofnjWi9f8am1TomS1A1hGJahPNe6baxtEBwaxRdq2eI+H6
7ALb71aoRnK6fm6ABhzRpiOV51wEvD3fvWJY75zZTcCsRFMElDUo2aEh2lSXo/UiwoMcXM+8Ocop
Bld65TmLUFtWNo3JF14vNKH0VNAAfXEomU/ESm7O4U2tbYzjdHNstiiV3XevUwB4AzSkMnRiLgyJ
ecx9rqxroIlNAftlZ6N6w3J1uPYbnz4wBCYSOOB4S8Ygd1uq/8WqirxnlyYxr4lg0ax1sJ9XKXgZ
wDptBht4j6LkH3cStTDjuCwT9iQPfgzQt+olrNRJJm3I51m4PYhp7PWmzjZL5DHkObPte7pLgQuR
uzaQ7mmoX3WGk+Qf62h8OroQdZJql4dg/VyIvqh19qmkaIHHtoYayPJq/kMaCZ9ESaiFpHhc7Eut
8OI+rB3EN8W++G8ghHzZiWX9xa5wWjfkn/FephC3D0j5o6Zk+8eMauk2y/DDlElqayaejpH11MMb
UYX7rHtAO4QmNjJ19NsFvCA0c2p6VbcT/eFHU+w+M7yuidx3/WVSX6w6Ugc2dEHUxE97G07zOfY6
QYkffmOKJ1oW533GA+TE1D3WGQFSearHv0K9MRB32EYFw8lmJT5TwI2jBGLGQ3U9EFbhgShBqlqD
5jm+WQj3iN8DQ2Oyrnr4i5zAPnq0lKrusVBfQsf/H60Wuppa5E99svQck/obWhOljnlCq8xyKcPA
agZTj/9DOhUxNGgDF5HkKg7IEQbF+Gaz2n4oaa5RiS1p+Xc/aZD1LcGztJxc1VpOVvuvOu4sIEqz
QMe2UR2c0mG/uVgWfZ4umN979PKoq5iil47cFj/7g02I1a8SF4qU75pb17E330uNM0PnajVMmJPZ
dHUk6Lxfrl9YqI4qLDZX8Z7fmr/rN3//DzvZ3hTJobxdgrKXF3+l2/1IiF7P7wRKalYIKKPGWv4R
3t7jiO6JbSWg/ipaYx4o/AJKNJNjd5AlROH7AZOfAHtsXr7MIaLtH7waWvuUDynsGH7i7HrmAMMA
XKZd9UPrWMwjzYZ8baO2joN1iWHYBdTOxmlZUYFmVGBeCYLrCssz1KVrOsmikiOwX/Wd99gHSDoV
BqQ1ntmwJfLSYA7YW13aAlmr56pi2cBiU/B4LXruBZuFPzNwpm9BNxkFzRpAh1NUvESIoRwq51TN
vVbDeKoXBInlfPYWIa8RgdCCowAnTmFNk85x8aNaPKVyNqNv+s5/uT/YkSIZ6wYSh1aYfDNGzt07
Bn4tFAR4tjDI42qSiUfY2QMrhTs/XZ3izRF2bSyjcaHe7CiwDjiQU/BxMAIREQozkALMmca9gntp
d2M+wQxS+wgB/Y+/FeTRXJwERl/xh4+d5I+i6s2sD6A3A3rkuboWSbcVqD6RVhAhqyWlEOUcG9iF
ieO/WgVOSrWtx78uBYVu2fAHWQE2EqWnD0X6IXkdrubIqEpDHeiB/2kljSp+ZEXvChf+Qw+uO+UE
dxRBsSMkWPkILvx57IYOcogCbUMu4B/nS5jXx5z9he9O7mH7mJX9v58o5dzft6cmUwAEuvEqITVR
wJZ9qbHmwl49Bkqdh2bPtPVBh3nzoGsraLFN2ObfD2nTeKdL3up0g5iBvsq1NSsEHcXWJqUy4hph
m3LWVVFj0XUshOvN8OyOWRVDDdvCq97GpUvkY7Rl+llxVyHZydk0IzgDvmOU1F6s0wApVfsQNoU6
Ua8FVv4WJz3vV0tmeudm6Z81sDaAGRei6N15g+xpP/0gYZ+QwiC6fn2AJXJeX9DKGvc9XAgVEV4x
2/I2yS52uzjqKS7/hi+FOLCCpfTfs5sj/sfLd22eTXacFkoyFpJzcFbbfpx7JFwuRPv2JJMcx0z3
v86iy5zYq1DVAFE9fexTsxZDJUAMXhGwfnXTDy3hJa18yLJRkIj9YI4bi17W/hGo5aw/COB1xg8w
hQB3tPe0s3bpquPzVxI/S5zUo8PlXoG3hW18/fAasQzmGJcpcLuseA33TPi8kyBeVSMI7fMcM+OP
7yXY52kaGC1F3IVY5ZNDJswxZvfoLn0n0j3MS5TAQLv+YVUZcy4HwNYgOdUMbl8y0xVl3+2fORG+
6dBuCjS4OlkEut9Of3lBY+2kR0lnklAK6DAdqmyiK3eKZoUdUkJmdHiK9UPVS5nrFIPwQybUe9i8
qon/P8Is+XG8FzpM8H3PK96q/oH4pV1Tisxw4qzSYydBP+XErfueEjk2DDgYHLsXaLXQYy3hMKBD
GvJQPRnMe4VdcDlt5W5U+xblQLy4kzv2kcXgzJYLMhm7EH1zkYv0AdbmnxeBq278MHxwbMftIXex
7/LK0rP5D1RAiBKMCWcs+sH8+LaSzd1xShssnpvwOS8GFJmTjNIO98VYK/evDPIEVd/aoBTNAyZw
9w8S6dnwyHzn2c2GQmJfXbTcR0C1sMj2C04EPoOJ8L32PNn4dUCewRxnVZoYFW77sBZedlQRGG1B
5lRSmHSGNGR+2yW4cwu/KADPXJ4gH+cpdxn1lgqEsjfc6AiREAd6FyPCNw4La3aUxv2qDF2j4QZn
oy7mXJV/oE25RawRdOQP5BRDF4GK/2MnrHmnen9Amvmk34l8RGwLfoW4E7+9MKry3bzrGwciPsrI
1Ac6X7s8ItZ/y/pJCs8QWYL/VJAbVd4kt8TZQKPWEQc5JMFP/7+shykOz5xmy65ZE5MgugGQWr/3
oXyR7TD5Qpf20e+mdR5khqpE4+xtaCcOs1zqR2OLliIvdwgBJBu7qw3WTF3SSLCNRq2fvATAmwib
20K+KOh3MjSZx39A7MhusBUu/e9cy8rZBxFsjm65q//SoP/TetO7MRNnjQrecNii5MNSUVzH/3TF
7RUTNM3Iaf5vuH24mFck8ahbfhhAbUMUsyHRNnLP7pXAnjMsO+VtT+cI0nO3LQoqDFvTajDI+Ok4
aVLZ/ttfoV4/+bBy4V2Vkox+0qqyx8KKpWAvyUFJN3YCWCsxg1xt5vL+0IB9scpGWuKdBfGLsuSo
+kY7/B3Kbfi7HPT21/i986Yfilkapnke0SOh/zzKMLrQfXQ9OurMLXdbuUtphjcDyJfeKFTuKOQ/
wD0omvxej2z6Or/UntUscM3hhLuPFWbNed5bVUvSp8gnVaQKFW/2r5SZdbGXvnVUnP+JlP538aCD
Typd0k07gGUf/XEiZZr4x7gb3BR+70EC6u9f7FmH/2NSoADRMv3BWuKM2OVesQ/yqnJur0nFDqla
dd48ONXdaSaZhyagFz4g7teLB8mNTyT5mT7+4cGrql4wjN+kJKPyVjdml2h44yfqjrqMExoHj3a/
ePOcEGd8ga7yWYkKvhDuBV1Ugz/yNOxvcspEmdvK0nMV5a3WhTT/LW8Rtuja31WpZi1ax5ilMc18
cz+LWMyXRro1qkGnABbu1Waxv+Zcm6hQU1gB5+Cu0shKFdkH1QxveWXIZKufISrBTYrf1KnLzo1K
gWmEZdErDRV20W4qiLHwqqIPALoOohIYGLlbk3oURpdw99DEE64l77lQ4bcEyahR6ShiQBednK1o
QFXTmdyCQdYll2dJnjqbialNDrJZEGBx5VmbGdyr6C2q4F69+7MncQZ5uqRpEkMvMFO4vRgYUHak
EWgzGOODeayomJQ0llRtFF2WBi843y1o2nB7XfssIzE9DDNx6AmKEFLFVObU5zJebG6m/Hknpr/C
gxHw8V9KEl/EG7hAv7GFwFNQXPD3uUUwYB1txOuHqpvvTYnySSi5BaMa8bOfIL4VqJAUUp27IC8l
1rp83LXKpvw7f4K4pMhUoBHHcKybBSJB+6cEUM/eROhfU3zZpU1zRe0JgL98C9m+4ZMOiy+zFEJN
zObNZaGoXvc0FeNuYjHiVKH1yq9ie6PSTe9mIufUo852t/KJ1kogW5ORR8PoQm1B44VFUbFK0zLq
5069YP6Xa/J1dhEuuXjkuwEG8RbMVVplqD0ZB0I7c6nxQIwR+Caau2ZXyMN0qcRTO5a+S4b+vq+c
rDIAiggOBcB6q1lCmdcO/ozcUS+Xyyw8I49h2uYpkYbfWxTJcx9zHbTTAS83jap+phvztomALB5L
9Jt1wwrnbMpQ/ZzyVqBrUhKCdvZEtok4b06tOtw4xX1sBFG5YlwN/EzI1FKVv5pBufghBPZfJQCG
PBRxsnT3QltlPtpG4UNRYWpv0tN7LFq4rgC+rKsdkjrAFjmP8L8qW1EDrR7SGcX5dA24eHbwBXBP
7QcXIlKov0wTj5lPMExjDMeql/iY1TBQliqhSiwh5aMHYiMJ+5AVQHHH4usxx4hrgNu53VNByj8x
n9xHNGScXa34XdTfZ4Sxm7whAFB1ZQcBqyiKzj5EOIFBXtojBAF7clF9ikDgOY3qUonir3QXWZwH
0P9AGT6nGacdP4b75uoVQSb2geTVV8C4B833Ih1FlKrv0bQCAmvK80Y1Ou6WizwWgTp970FfcC5/
B0daIW90VCUSNbcnozbh14aMreaoP4aCYyKsmaS0X0K2v2V2wZCB5BhiU1t72g4ATrFw5j9BnF0a
tMvYWk8yh2Emlmo6IiFuTBleoQFtUsNEg2aA0tt4L1xZXB/RM0IqMR24YQ21RwSsD2yCEr1v69vC
3Wo+OqWXeBfRH91q1OBVU29DZH2s1mdCBzeeZTsCA7SuoeDaLsgEUbcwLIVumLaQMmClm/ZcTOnQ
Le3pFGwZ32kVuWR03O2diH0jUG+aL1Iwt55YxN9+W6xoZzRun+cIMT3raT+HWQp91iWbJpcgyLC1
/Ugqlx5Nl44WcTIv0d+WBeVxheYNhxtoExJJxw0G3JiZeMNFvOQEsT3JPIwjTlIJDuMI4laKlwEv
3sZ4aX5Cz72adQHmDVITmjMB5AxW8ILb9W0pvvnllpvRPS/ISMd9PqoAIBtXie7M4a/xE3uGy54I
9Hc/8I8b+opceRr2x1q+9O8LFo8pXSO4NDSH/+XPUP+VEp3qe+Moyz1PUmA3ETHp0FdZx0wQ8Jve
rZ9ZwZzDXUvH0Yw4Ko5EA9YDbLXYSzo2yCj5JyfNJSb/CdYlfCtrrjfI/OVUSZuZGaX8N4YRxDcJ
pSQKLfJBJ4ckx2fTBw5FUBybiTuro8tZq/5g+6M8KTdBWMEcrVmVp2AOr8dwE9AjNTexPs895/fU
1MX5CW8Z9qZv9mNGvZD6HMAJX9NC6gGZ1CyNG0sz2JzjVQhsz7vcBTdblTJWKrS0MC+1JHmVsIRt
x4NDUVE2ZSaS85Em3JJOu6zLCz8vmADC2Gf7oknoJgZk3OSb4iB2u2iaacCdO3s0/q0DgKjT0pmD
DiqKcze9QdU5GMIBbc6zn9MNecbhbaWnGuyXBxQ5BrVrZ4r8KkqWClAcsjz2dK6zAFt5zmHlhbgN
vTtNqzeqpc/mYlkQWym/grM6NP18BmayIV2RrcOkg5U8R2VoeyLouTd9N6L9HCoqV1X5jG8dCHAn
UaC0bmZE3D1iiB7krNZ/1Z2Gjg5XPKZN0czjkr6VfEpfIclhOyZT8OkZ3LjsMg9ZYIzYjt3sii1P
qi0HVmjoSOPlpAFGci04Rb0cBYPaRqWHWZ8ZXuh7HN+YPb3iaN1Y1kkg9g4HVloJF1gR6LXjNiOA
Te8au8QnoYdvjQJ6VrYXDItIGsm4LhlAqJLDonCnm9JiKW5o6ZhU7CtO5Y2l4FshysEijPR9RsVO
45moMzYZznes7d43id8mW1NsvP+8ecOQOl9qceji1uv7WctSuW0IEKFle1jRHmh2N8gfmvONh9Bk
5yH4QLmJ7AUOApTuFlBz8N3W35mioivxYu7BP5XprYQlwXkEx8hso0BoRSfkeFe0MOCiucaDsDDn
Q05/s5r85CjiUbm085Ln9/+MRNxf03JZiJ46EIzqgwhUjjm+AWwLWyCp1dJymQMGCJUEQieMB6v2
Cj+f5kKQCgNiAhwgUplcm2BM5yLQL+KX5M8G/X57vZglb+aCNQeL9lbLGJkQ0AztJCCPfYNZ1usF
yo+JAIPm/MZWy/d5tvy+hRBAeSTl8pWJ3yj6RkZQ8i5lIBB6b1Zc2xdsA+xVBV43SuMP/WPnpzci
CuPPUqSMOIuN9kN+R6Rmf0vB7eJHPBTX0Xq3OZG4k+dK/wKpm/v9Bqykl8UIOiZqGqiYtAoqNhDV
+x5y3ySanqcMDePeyjvgXEV1w/1GUzj7Aqw8PFBS6crwWK5iNS3WTtnrDczCfIccY7052UImV0w1
X7p5RFpffHRnzZYR3kzuGzVWZ2VVB4yxv7e3w7pjyU/xjevuzJrv/4ov1hYI/EQqpvCh5oKvPzWr
hfgwdvRiYkcICRHRPRDFxQlPnD43G5hIMj5xiokPDdNAalF9gI+7U2vDZj9wG6js7Bf0/pxKGgsL
xwK6pzR7tixKcyn3GqzgL8p7ype1+weH4futUfAJqOU5tSdToHHpUcXt7QtqiVKxgoExQZ/tBXei
d8QHp8UbnYRDbBXBHsc4tW9DKBwnGmC0Tz/iXDByBpbrj3fachG+mUISt1jRRnX5WVpX1DF+1GzO
UD6gr4DVMcnxP6Raa71QBN+3m1Zcf9ofolR2y2VaREc70MXZX2cpFqfOjEZ5ST0NqhY043iWyrJ1
SQGgumZOsoFJ3OHn3f5qjc3j4NXfcOjFQvoI0lbms0WjKqGnvja76AK2tC4upkB22CLidVMRFQYR
M1G31T8yR7fl0wXD58OJD9fkw87M6hG6u8ffhxxYIqRy9/motJxjzbtU9rG6uKIKM/KwnKUJxm5p
tKgKwiw3D5OWJkMNtC1+P0P5KEKlRccitNsYAHoqS1EaqIYiDZpx0gvUYX0UMLBrG9QfV3FmHq9s
W0BqlY06e25qqsMjfeD5dIPA60lN4uSj7G9p/eh84Qx9C7hZ7erV8t03qzZBjy18U5Uk8KstqtHP
+lJGKEtHXrWXQlOMJOIosOaGFWsnu/RMDStgkSlCvUhiebzvxsDTb7oUvHZadfRxwEukZCcwoN+F
J7jhlLBW42WxZoufXC5vonJEXqGQiJaJxq84jRlEtdS+RWlcvcjy3SHneQVKxUdUB/a4LcZHEfj+
mxEhrR0eFDr8SwIJ7nhIE0cv8HN3JiVPTi0/ADHiPcpmKHHIz+RokEQkawsWbbmVVN22IRFCk9Gk
+YLlsE4lX3qahMOCevb5zYKAbtQ4gEl+k5MepytIoZ2/Doha0ue9m31PLEWQK8TgyG/DWWkqRcR6
GIRSXkFMT6s24v64MUQJX4tpoulmDXEDQKdjNfJC2bmhMvs8tbOczajbpea9OdvZYlwJMIPAObor
Zn0xhHLoDXMzn1X5b+BV4vu6DgO6yCALXige9WGl1me3u0SeF8aUVUhs6u2ymUWqtugfIYdbA+op
WD3YR0+VdQuwZXXZXdWcYE4z+M9scIgmb0acp4NKladqu5fNzS3GDpoFyjFO38aFCgO3rpIAjA5s
a97Agspd8tjRGTVX5tzdRAM7TKl2XR2mxD9PbAc5hA2WYmewlH+lDq/XythLN7PXEjaIX6/AddVu
Mah8tme17/Gc6wTUTjHqTOC/KQdAij15HrsIKO8J0PrnM3PJE4gtb+cSyvC+C1XRbOmd1AsmfSIa
iODKnPP5q6jmORElsbJXRMYPXXZ/sOl6o2q1zMglGoHloJ9DNXrzaOMszQf6VN0FV2dRnA/St08+
RtBz85KaQ3SAje1MqPrdSLLGlfw7MTINMwU83BoJq9SIfKd6ajPJMTCGKtVJw1+4X8qAMRUIfneP
HJvFV8fZsqc+iMfLN0JwZewT8qb3pvsMqo1JxTzrSg+NrCFz41Vi8iNxBGOiTtdDcmjxk5Rmwg3p
ktmXRfREnXoJGlbaxdKWwdO7lOh3lyQJmZyORCwrzn4JspIpEQX2guNxLoKrnkh8mNvyl/jN2EoP
CHXkxZJbZXZNhPeMfCWaDdHTWxTB0SI9WUkXQt/nd3dj4w1iGNWC70vOOAFgZ4kCbPpmmkVPtTqN
BrYWj/2jLSitnJiT6yTKuzQduTl28Cci0CHy6H0b5XfN8q5b5PRFhQzj8nvwmG53fsbqqCPTGa3d
NrpGqLqmRWMywY4qwVj+6FJ8XkULsPUGPR5d+PEgdNwH+Imrdtdkcuit4zqBc7yr3EfhG28IXNaE
1XLQLqFBmyj7ON0ma+Xchax2xEEme7ICoQ1TO2GWaKp/QjseuHiwFqXBepMwBJ1/RanCqbZwmbxd
nHeB4h4xwefPK9H87gIwWceIj+ttqufn9W1J7hPecYOSY0wDJQ5OIaDxECIQCKFC85zsqcHIugPr
YKNqBZDqXPbjFNEnQ8QZw42vhtL1W653XT3sAim9bn16PPID2FHH08yDD8dZDOiedhXvdMNY2CG8
RBbTzzfMDVW+v7LXpriuAOndL4RLzBcLyQVePFqhssdpFjK/Nlf5DgQP86Mf/bQKyi7lktjDwEX9
0I59O0d76X9hJz8ZvqKTLZ6M1I6MWOm5Cpymji/dmvz6NRa7v4NosJ3eNfF6DRhinSWJWS032oNJ
Ycllf1uZrNFE11GWtbB3lLCM/XuzqKSINn8QwzvyW25I7gLoZwC/qNB3HHYaMjIeyUTGANBFf7QL
Jym2bJqMVxpEiI1w4yZ0UN5UPr47asWLV8wv+7ranPxJtPKDhuiszfqo7Beise/G6aWbcSStiPh/
tPe5tScGO6wWa1vnoYrgeHebBDPGPuPH+KtBqTTa1LlVY/rKe/jQ6ZQF1O3TmtWc0kpFRuXgojT0
dstR8MkH7vdGOeqvKg49KF9RI3bUiLEkZJD6UmyAVmzp1O+AbrEf+QChi9ocOsM+dwx25nVPctv6
R+wZQwK5EZUWcjxMTq/k8x3Eh/LpUMj2Kt0F7jhkngbuzXCx8nD+jlmRVJvTOjjo2f9i8lil+dmb
GpB6S2SGCgwOCDdRwt/7sstunnXWfaS+08XyxRTISpHHorm3R/8rrmhit5Z89XacjF05m6CwPzfe
a1FrQfROpvAy5qH6H8BBk3QXv0LENCtEZjzFuySrZvUjuloWGDTcbwlt05NXKoLXWvM7S1vLvMMJ
Rxwh1U2OrlxfT3/ZMn9wYRCfKXoypliRLScBvkkXV3k5R6ObW6BJ1Ux+C+AGRoRHynjN8afEa+iG
8UROptsjRCMQK80Pa8yW7TsoAOsM5rmgeoSE4tlOAqrg7o5If1Y+wQMPwphy33nH1344OkeZoUYt
+x5YLniTJvA3yBIFkwxeNkxEaMccQVQxIfHCuM3vBa9/jysMPfDbA1B8SIiuOxEmzBKvFks1cX2s
OppUzGL2Dfj54uxlgvea+8pmDbgnxcxq5JiUEoGwBingRmLp2QAtotRsA4hg9SNaYV9wgoKNtrLp
7AAZiBand2Pm+XR2HfNxKU4LOgemccUL/xpbkmT48J+fmwW31k6+sR9qCQTdMMl8d9M8b+FtWDWW
4+hqfKNVvYMwOI2TZzWtRMWV70mpY/bCnsVadtg0X0MJtATqZXriBCjRxgvtUQixwx7S5STRVol/
zAre2bb0iNVQS3hDv0hq52nMWTLQpO2r8t9Z5+XFYClPJ8UPtG8KZprNcRaH5gdIhZax1+x2UmC2
OYDSYqSP78jWBQXtZ8NfJKSL0hRKKMQ3dL3go9FPXygQCRvrgfZGux32GLEGfi1Xfb6HHd41xLuI
d+6DnwMwzdpvefjquJmQupsQy0h0kh56SGDa1zPTYv8MAeHfYS7A4p4c6UM/DGsazjrkGMHcY2OZ
OUhv2AQZt3JngmRO78iWqro1d7yR+PeH1eoSQef0cDzaiuFgyr/XMyBdQPNmHO3Q+1QOFhY5PnhN
D3/blFNEXJII8CA8yWn1Y2qBiEUADRZzsedIWvXurYFDVUEMRtit5xirXqZKK4/z8KZlKyL3Kigo
PIvr14ZbYozovA+2PU3ygZPv3loDb8s4z+pe9FFJrTOBBmaUb5azagbxrTV4TUEKMcDRJn8KwHzG
LcLVmrkCzClV/WkKXgce33yKzLOpN/t7imZpicTghiFdUkF/6bxo9Yjd/ldGtpxpa5lYWyWQb/AV
aZUQdQhRyXhvk825tUtDPgjtm1qo4QZjRoOzNOnUdMGkZs+6oB6uUSJUOOgp3Kz2GBGBRE6UDzEK
qkf/UYlcSnSSyWV2xplcBhzs3vqWpuB5wFg5ohEcKSvhri/IhUAp6I/vDn2kUnwCMU+rjrwd3E6w
PcJQrYZOM+AjBTB1xa3cpYoZYlf/ZP3yKHoLi+4A8VHEkTm9xPE8B9Qql0U88/uJF4ke+O9LsilW
GIAN3KWHFlE/NAlAZOhiS9CDtY36Whdwoz3SJ38C/SFckUNFOrhOIh1lYMjHlUrM31c6rIS3pWiN
VJnhbQZhf5JbiprrQnxqYVRdlxLfULWy0abiQJJSBskaTpl13fM39TG4QoSCGRh74r56sL3zO+Yg
dyXrEw1wmWPPIj1BilSXv5F4i14y0ozwT4TYpab4l3Ur/dcMz956NHke/N7RUHe/ZbJkCvrh8Cnn
QXLf5offeA18B+kNBX5R82IrvMs1I78+HstRWE5FW4LWVGEOmKuXjNITxyyKl1hcJwxkGbNw5fdl
dNZ6brt4hy/TrjH+VT2y58sq1pelPgGVr4JAAmp3EOhuKlBWbnjQxBD0++hE55xYbChxROGayVDm
WaoJJizqOEq4jvpsikp1QHPc0wXKrWdZ3XC38T0THBrRIt+4FTUwonBjzuLl+xKPVp3vViqNTcXH
t8dWmRDcD3VffRKpKAqNKL9pCY0JKBnLzvCEQu8bvJEZfy5nYhHtyN1WboLndCicpNsv2SFHyIUB
jYD/8dVJ1F+7aTpKVgG/I0KKRAmF1WHEwhlNy2Frd5aYlXVAjzjPQt0dM5TDTloyl87qn9iKef0J
UtcuNH+x4vWmTOz4AlDzGuWBCLPZHb7XXK/zVj2+Fj3Vm+S6RwVCIZbFyiPYUalhQ5yRrdDe0AjZ
01Yi76gEhkz9L3jWZKt3L0jMUOdYe+XQND9c62bE8tCpyILkNh/0dfJo+XDpriJw3xByol+c8X03
qhW9iDWE88CNp5Zslme1uqNVSJCOug+gpKIJpNSDu1xI/WbVMdxBwJvavo0fkATADG8x41D6fdQ3
GzMnVGR/lwUqGnEaQG9YlbM3Abb4Qei9UmxvsVRBQ3t4TrHWrSDxoI9TRWwQDlXCCv3h/AqestDu
4kjjfe2m6dGCtAKKuMBbqheEqXPCegr/PnlQNRIu/Fh50TaR6CkrN8YMS9tGcZVBr0+dl3AAzn1g
i5OhloerwCzv1iQSlKap82mpONyRsuIyhe5wlKKm/EZIa8oRpDO00zMlN7WuR6wApLbFFtjT+35n
zfVFv1pmCaaJ/2wZhe2+M5hpt0yPr1Ykl6ctbm2azIU/AkigZAXuM6Qme1i5XM6aaAhPZOz1+2CS
Zu39MmsjVHW2cNX5fshKJZN0dim/a639EK9xJwa4WsAENysrAuVZecmCW++VRbEgLlWlajfJ62Rc
6w2GSQzDNUBIMhRYBXQTgANjmBQFq8JnOOz7vjEBFCymnFU3S9WSFNAqS/2qccvMMXNrEC3bTdzJ
n3IcIp0AcquR2DwTMOeYuAjsJXax/VX5MQw9goA7Rqm6dZlItNFtXQhGjDrXbkanf4QLVHhRa5dj
LoimreNzfjkeBlAQbn470uTd58WHfos28qBDx2BT1KgYc4cytpJVoMnohOeIMoWB9rfCkS8qef3g
UR9MiYd7sS0emfT2Z2g5vZNAptLzUOiiYZCeltZygIgzUe7kuRDOBLbkLx6sL0mMU5vh+QokVK35
gKGnSnhYuxNQXgQdjEwbxKGrnoD4UdKoRlbd9khlC3ckv/9khoWgLvVygtkl4/HgLC5FAxB50aDO
ctbRerYc7qhhW6EcaqdTQWZx5/vDoG1EYmt9ftH3KAB7pZop652u8XtGm9/494jI7835RaKcUQJW
hhF1wm0RGlGIJ9Zrm0LbmHgolEPbP6zNXqaUbuWQ1WsIvQ92CSMaW+ieMssafC7XOvkkrP4nIXcV
M9gEmSbideYrFeT8QlctiGKgP/G38qjTH1v0N9gNNpR2C+LZS3eUfnLThQzojehv/UIyOX6djqR/
PG6rlSbQpYoUD5GUdUcYVKR6qqT5GCn9PJPK2vVQgwV88tsqjTBkcVTk+DFSxR9jYJ/oWLeX7I4n
OoYl1hh68M2DDg9a+z2dDwO4LIMa/tNSagFRLv7xFMw0T2X3clDC1fYhIdPp6TjuFvL2o/4KVJPj
8aQwFqtC+CnJF1jp4XR0NzpuwDaocVcZFJ2ZKtkSS/mX4KWPhBv0evrlULDxLxJ36qAUn9KaFUDI
ne+1wNKAXv1LDL0xeCuSlD0mMy+71OLY+rELiydgRXxLmD20MhhmRs/fJJ8w7vJxcmatdUEGX+8T
fUJTZz7Cm9NJNsxPug2SdZWXKBSdHFZVIovnCejcbVBrQO4yfPd9qZvEXIqKD8coE8upzhf5uFsX
V0nRuEQ88KGEm1M93qyu+ppzImqel6zdIB0wUL7rdY4jN2qAZhf/YEXONmIUZg2q2y686CntdrbG
fCC016/oiLN5jawG4f0/DNEogMbVcn8CVDO44fjQJ1SBt/weuHWzIF8DNjqioOkekbOPcXDg/zJ/
003K9pbtsm7M9Qfb/3FgupIYDtQ/ymS/Yznh9nNcHqPqwnOsbboX1JVTErYHRe/uXhj8QmKDeMko
odNfATDsJnJM9I5hQlfOFDPzUVizT2AzG46I/v7sNoBFpE10dPxMZBke4pe+YOdEjnV/WpH/NYqf
WK4HlG/MVE8+xFyueZy6ZI/eG+CQRCL69rsC9ufggoPbWbhN2k9fVwgSbZIJfeA9Fpkut9rqD21/
r/4tJYJnpfLhEUykzo2wwCKtYXqXGbdZFKucDPUOuMtP7bisOOMASWH+fqznBMIpETcQfFYAKItW
cGtbvo1AnJAzugWvVj2EX8IChxv+K2mLtOFqymPcnNxVKFovZNoPh8KoTE3+9nWk/h1PJUOSQ8TS
UiRd7REjvzV/Mij7Ra08YR3t7KbVLhbnM/YTGrGv5QfnpNmqGAIVHwy6f1YFsNwAn5sft2jyev7c
SLUS/Byuh7YHXnSlR24DbN0FYl+w7b0yM2SH3ELc0gtuEVJHhwyCdHWDTi5iLc0YSQTS8O38+Nnn
iMrMNZqPjpVaSAHUR66BsXn4FyBcvZdx0gXU9MSGdm+mP/se91RTjJsK+pAYfQizS8iWsA0FDEyK
wpt2q5OTksDZpi/uBWD9FD4klxhimY65tJMvrVSPaRxBg5veqYFDOQoWWI0BYLI+hloPBoeAFmeS
hWYPPre1K8gB24dRUEXzFVwQpQEllRBElSJDbX3w8d6eW0t7bXojWnOS/4PVUTuBoDQt0CWY5fr1
M6H0P0o9uwWrsFKkvy21pAy2jEQ7BdT1iC975CEtWoBvRrPOBYHO+LBBn/rkGEvsCfpYUz5kSWFB
tTHxYb2evaqWYyybD6075hgX/CJc3AZtyI6TiWINfPvF5ZIQ9MCWILoptY9ti+P0P8mHrvkzvtMk
g4jhrzIWtbzg19xVKeyaBndFux4VpNOSkmGzUq6WNekZB0PoWvi4s0HpMGSwUk7RYBht1ibeeqYA
o27lAra6/E5eS2iZBJU3mZBa9kEJvIwvzloj0mRQ3Zo1JoQwYh6GFYZHkPL0rt0vWDas8Die+9p+
tzfqEIqxKtCEqvo1npMvIVu5MmBhZlauPBOI3VYnWHQsJHbyZ4Ct6C/o0VuOkrrl89HQ6dwZ5N23
xcOaqw7H1QJG53aOiLnq/nrrUOXkw6qoXSmIPXDag0A9eVwqRlef5FCcGFFuA/bdxtYJTivz82dN
AZtK65CVDZ2b1xoUzrB4qaMTlin90WRfJ3nKj1ZYJ/bKQb+AiWjo4P1Zj94p+SMan+xxAPezyac0
MIKDOwr4vfCMD5ByScEHdDsc/6oOG6pb2IenPF9lEgubShAX84iWeaPKqEVAySOE5oEDiUUObNOy
MbQILjqp2IAZsp280CliIfN8yAq35V2XhAOBwUI9FQ/ksnPkW63eoJXznJWITsMjRENX0/bgc+4+
UFrWKjg1jh/ArnWr4eEve2IaonaQSwEuSa7uswCAN/ZnTJCc0TKfff2/lfdXAaVuJdawNiXU2xi4
azA40ygAytNqiX5j28K4drfy3Ph72MDX6/V4VqatR6mYtlKLmeFFPa1aFJoJ59uFdzl3UGrxRnls
j9XVPfYE/EPdUFwko6SG+gfcISeC6evkF4GFtmZD/4dWqYM2i6A6z4OcR4YMsOTp5r6JRGYQPatc
2PDRBbotWQ4INeVvOF7ZZ/fBQ6XaVhjS/Y3sGp2dcPvFJi1y1noseWFu9HUkQAEdftbR72VPXsUk
/wvxmE21654C0i9RVbWz+IcF9VDCrwXzoio7jtRl/tHtb5amX8SgbqaI1fDwdT0YSWJyy166dMK3
BCBeDul72LJIBHRHptGBnDoT07+rE0BalCqtJYDqEEL7jzoNJEB1pXfh2djekLSzC5Yauep+wHS6
ot0mFDkYmewAjKvHhjj6QtkfV2S0y82hD5wgWeu78VsICtGNySIXDTXTlOw3vSWSTpYgvh1M8TiC
rqDFzQtpWbvEJiJhm13JagPloq0VPKzhriXhhfGCloQpn5BqloVSkh/pq5ewEHZd99mVaGxN+K8k
qW29FodUGu77zbbohTEc+RsOLq0F9LxnMaaIlUPa2cpjz5xm/Koa1v4CsJKo/zkYh5ky0H0ON/Is
gmfDDyMur22B1oo25trSIoB5MCAbYqSnMyjxYyDCbjLWkCIh9N+YMYs3MiAHMCP1bSPpkxK7hXOV
7dqho9UGhazZ8gEeOurx10xR9ByKc108pt4Qj4aYcuqdyoI846l+NQbEtpXTU4+XFHujaS85pccu
one+9MnDzWMZwpbMG6dBvPt07zvfRBZbDxZ3yTlyHVPV6C2/7ett3S6Ohizv0lM4CdCcy8ikTlu5
R4BiCb19ivc/E142jQy4K1oVPV3rICBCz0a/zq5As8HcubNQEnApIYVZ+teHGIUhg4MQtKTHqXa1
gAH4As2zwGHCk7gX96zMdOFpTzLrGx8cQtGchMGDg2aV489cSqdMPklvVRepEP+8RJSBlYbOTQdf
4y1yq2dhKQlIerXgyy2yRwSAC5LCpxkOxHdV6AgX7Fsf78Zuz4REPwKZkdbTGNP2Pa/nZAyUkFMj
oc803+CeZolbaBZsFVCHwhsTNcudO2iz8t1rtncua3jb619D5hypNRlQX6hxGUmC6lvgJHiGf+YB
HD7B8JJj/Yd1pKwLSyeTDiYcTpXSbYK/IV0jOf6ItXcV0qcbx+3uQsww34NI/xtPLSdxgTaYbo2h
BG/tpKEhFjx/9hXPKrV0bmLw9r+Y0jfpXq+8jgPzy4sN0kCzvmJoNywwb8koB8rgV5uqnpGXWrvZ
wk8Kkcj1bFpOh3vta5CSA39KnvoBQacaLcy4xw8WTgXJyVeZlkDOXVxspt5WN6ot6cQGhYGhxk7G
X2hs5+kKoFn4shUlL/b+jT+wzN3g+fhM0m4ZjbNRP51rbKweKo2xqrfbCOgBuKHP2hvWSLQqQDqs
GaUjBjJY9xguH61PNWI0pZPJP6CAdxOTOIAJAQTjiXX2/QQCxvKxwrsBgH1sus46t4gKwuxAvQk0
rVnNE9wWZABLbLmNOZ2DdVZ3gUImYvk8C7wAExDnTrubEdGOzDnLAFZjiP6N3PYZPP246goM6wO1
RRDPQFsf14FYX1o2YcVvPl6IQJMiP4vguT8ROgKdXTvY2G2f2RklumZhJmtexon9Nea0FE0c1leZ
jVg3OD+ZRaCwJMHGfvM6FXLEWlLR7zBa7Btbatd6hpbFatKV5eZDFgqXf62do1Zii3P0SE5IS5rK
eXhRH05yy4VfqgaPRjq4GfNuivXI2qMLMxbFE+Fumc2bFOr5xKUp1Hw9mDzbHneB2ktDpnttSzQe
SggiiFy2jiSqyZ/FHLHju7XOJi55fIDPSfD4SLYKakO0+95aY7W+pMjIKSXiSZXnkGgIrHoFvQoh
woi2KAn3c0DmU2AgM5rnL99DTXLFq5VNHXxUcXTsEyq8MirpLs9B2L3QCEYS9e1uMo9SZV0QlRMZ
1Jtlo98mGyIRCSdEOd1l6LJAzZ1FV0E4RTAdLA/sqIxNFIDJsgizHi/0bdiPq/cyJn5Qh+zTbGdR
nfAyICa/2d4eDwckX483G4FE3AkcFUq9r6TUyjaQgZ72Z44TiWKtHxX7I3vvfgzDF00GvqlbRX+1
5wXReHdArrKDGqDRH5U/bf3wRJd+VfG4vkKgHtm/aV3sg4fnfpz8PCOtF8az/qIcZRk/L8IRZ+pa
193n9TywnYjKYSLlL2QqvmOPXubIQN+c3j9Zug1rq6BK9eS4DeQqWC12twbSAWEOIZsodc8xTbWB
jIp3VojJUoZz0mOibOeh55F6VwI5MWEP9UNh3ttVQwMq2cSrd1hbFRVuD0CsmUJ2+ue/IxZJV1sS
I7j6apjynWmPi0oLi+NKiqDOWoYpbyaFAGtygYtHgkHKXy7T0aMXW7kopei41EVWreBu0FsDAKXR
vH+g41Hg+hTOtT3vHBVMo0M2Kw9Z4iK43eRjblVieVpcRSPkdOto4hH3FQ3T8wtbimZ054HLXNTE
zpXmotQ6be6RpIWzNME7B+WCY6TV/6aFWvp5xSfvfuXvcwpFgeg89G60BsWiMOyhzxi175QLhIxL
xDx4/CSsV543bA8TG8DiBiKD18uZHZjObLE/Fp8w3712ZeY9Faw/eA6xQ+QY2RgXFPW8tfEFSeEA
doF7eDssHzygLXSZY2h0kOtrC6f404wRnQ/Qh1xUojgNhZWEdMTnNA/bq6U9qmcmPpHw7mcuq+Hg
ScJNU292rZ9jeZp8hSb/gsopq5cFUi7KXzvFvsDwuC8eVu0ra20lgc0y7ckkfmpd/XqA3YlFuLNI
2eqSui65D1cr4DJO6Q+Rk9F6LItlbH6j4KzeRHCWiR9wzQP+WbmbMNwXVRdpndtMeOn3oQtKQRmR
apMPBK6mhpJI2Chz+6NGg6kjL7U47E6oK7kcMYLr17WSNhXe4haRzb3KE0d3hj7SyI6phxwEe2C8
WiekQKv/p6hOufdT0F+rXUkynkSd9EcYzDj6Q+BzuQS2pCU6EzW4OzGGxdBp9oMmacDnWl9kivwi
iWoVZL1ZclTV01aKo4HbMudHeNB+zdrs77vP9agYx+UYkLzsEHzMPglpOs7YRYqWFTTi+RUndvlg
nHUSsKG65scvudRZZfQJoEGLsafcLiXSJMUtSlTQzyIablUYutBLrfTK2Vfd7keLNlLQk36jsthm
VEcHZt1QTijI03g0Kb9x/kLxH1jaLmUe33TZLgc10x/+pmqLuO8eFly3Da+issBIh8X5WKZWe+KG
wYo1uupod/QBuj24KvHFUiJKkWgRtPN3dnywOv+opVqjsp1KhGL9eS4UKM6BPpHXCZOQplJaQ7Nn
FpoSZlN488q8Td2QgMoH/L3c5eXDJxOT7Klr/RrMGcRVNeSVsMFLD9cgjwZ9aE8QsZfzhXv2zP5u
l+Ipzbiwa1bpUbutRvJnnq1hFFrcbq56icfpqJYqcJLrgIiEPZwWZvhY4Wjp0/KHXjNHW7SJdeRJ
SQiN/lGaRbXS5fSimVSJkXWTHSpYdHkHVgwXA637g1S7YcbvhfKFmEZyEkzWZQGohGIqeDcj2pyT
5MH4tk4hG3gCGSrAlukpGyJXCjNt1+cQHgMWr2ObbvgPkyzeC6H0fLnuArMdz/16q5Ku8B+jYTrb
hdW8gRiLq9LNSAH3uW8X+UnN+fp99YU8ZP5AXCCLp6tcIRszFI+nM7JX7rFmXzD4cvFc3UkIyF0w
x6mjKqPIw8D+MzsydtD0/DUxAgtaLh/0wmLujQUTyjzaGlHYhcjL06NZDvMltBLBfeCUFqn2GS2/
yS/toke//e2a4faa1D4OAtQIIOtCeoJBKumsHfyg2QWWY3hxd0LTTNYBCu5i8Jfac3BBHfdzuBw+
kA9WhSQqhAtfw0LuiAlrC8To8cLUz4N68NDnzzUO5L7qHwIQ25ciEDS+Os4ulsa59Q//Pdi+YVKw
PmaPVxPezo7Hbse8tqvJEM0kUyB75wHcq3SVDqnaF/Smml7/FmnbTooiCHzSw0H/v6ELsdRet1t9
S6/kzZNh4M3So04B0bTvS28Yud2oCLk8jt4fD/eWciam2fBUdY3+NvTNpGRh/qvO02Ho24WrkSJX
yg6OoGGmYXUW18H+Sc8skkRNxmRwI7WNWpM3m2auIEMx3c3hU8Y9hwSU2dp5fJ14lVAW17mvx/G6
0aetVgAu8kcQB3j4+hAMNWRtv62Ix0QeFsoaa5XgT//wzHqph5HEQQ+cXD/PkSz/v3DZ/OnyANNw
uYihLsYM7yfXHfeoAE6MMuhwbq8BCfcokPoDtZ+DJBUtsSB/NzpDSEZ4fPHRXR8KIDEXYRdFq9Zo
QjUEPb5/Kfpe6g13MaAFsQI4cqhaWDwd8hG3mMclH60ekaidMNbkWoaNCD4irPDvGWHcsxrQbaCa
YF4tKwtvHijgcfU1hqHdKbMDtLnQ6daW4BRGaEg/h8OsyMD7djQqxq43J22cndzauMELTkFH5HTc
NqPQj2825K1HgVsKlfBsfvl+6kwmcCGj7m4Tok8Q38fAgDnGU2Pr1quOMeag000nPc3elskGoK9T
3RgMk5Y2O0w0oKVds2lQMSyJbHH8+L+VBCCE8eJnbWzLy4pakXFVr4e56xAdeT0IFAvWz3jw4nGE
RafiU4bNaorPw4SmKlkQodwhgaUGVEeh7INWPTFAyAfA2R4ycQGz3qLzUZ5DdfzNX7zFScx2fM8b
XFylvIYhtHi3xOSTmlQ0NX9NphJJaFw70lJ15EHONjjJMuRLFxqYD9RVAbFCDdskC4jpYuA1lN+a
wiAuRkdlhlbV/9z6S9epy+uJCqevEkNSEuPjue0roCgRtGXfqfebPJAgmatAC5WuXfvazGlYQ2ww
Pt+g+e6RFio/e6o5YNDVUfqz2p461IMwkJZYaqxaQ1eaQ/poxC92NTlAOjYSKA+P2EOLZOLPTRbX
dJWvKDki1M3nksr0P3VmOiPxhX2bMl0oEFOTR7EMe+IVTfTTCgMdzQlsS78HW9hb7/fxGcmk6OZB
rz+AE+cI7A5kRDAlX8NisAMjnifmzIIVzrrE5tSgoVOdAIOqTkD5ud8X/btS/t87tls5OlJcZBo/
VUgb3i76dPzygcHYLlWZUYap0U2bCYOuxhA4ni4KRI8DJxpmkvurmtw1LvPx7p5jbxWLCtqgDnRD
DCYBU9ly6/ZlNdnvZLmJB/pZuj7Z/1cFM9VrzD4+tL3YywwQNbV5iJyr2ydasUKQEAClTy9N8/Ki
l7ngr6D36BNPIW3JCtIOPohOdpJjGLKEnLKa7cn14uK2Qw0VTyo1VjSLEQLp28KOYPcmRvJvYQp7
WzUap/QJYp1NM4SoJgsNENzKl9ob9/qerwFEZrBF3DOALAr/m99uumTHmomFMF0tJ+Wf7cRuEYXN
pxpHNqy5ZIkvVoV/Szq8JG1xYLjh2PFnqya8VIPOuyMH1rVSbh9eI7PJevuoR5GRMJrGPyq7kUfK
QLoDZaQXtlttoC3rnB0P0LHWOwgojJdFaqnKwvg3A+vk7yh1n8OSmoWS9R3uv+ZLhmEGAhUxgSZ3
yaSb4PXrbgNVlunuw7QITewVa1cOi/ar5/8csGwddk/TIH9Qyg5O5OLfnxDrmMzCmHLnFqyE4Wrt
4WY1PHAHnuPm4gk63FasFy6hLaAjLK+qjkEfoOEoAMYUy7cvNErUtjn6Duf4vGSrttfVth41rDSZ
MTMykWndzos8ZytwBItBYAz2XUBF9vkvPwXC7s4yZAOm4O+P31QmGGRsZLzXQa8t1vMmNbwIdXjS
Hf8mvRs8iuTFzf6m1Ww/2si65G+Zc/bcc3uqJluz6w9Ozyfs8OL9Lv9Nyn/4JmnG2DrcT0GJYwBr
MRembxCPG454P5TfQ8pFjEM1/Slp0giSQG0YQJpBIC4uULHAWXEBtO9QhtxiLx/HGWonpCxr+K8G
na5Ind5kRIuhIJzEeOXecCHTsHlZQJFoMZZwTL6sjFuSgKYAIpF7QKdZM1NYZR4cgugXCLmSArQ9
/ZvrHT9sKwNKCoiDTt1q6uFTi8uTussSYDLr2JE7x8OgipDwS0zdcjt+MszH0cdlnF79X1ikQv7k
73ySp6Hl4lXJw7Z1ViYE4VIdelSAV2z4klvNs0RqcAgebZvA7GvowRp7xjEdfFnKIV+5PTfC/viv
TUpx7SVd0FS5Wjo/v3MFZS2aRu2nGuMhr6qoUZ3uQNuHJphNyK/+uojvCrJDINsttx6pO1IOF3HM
nrM3U/bGcu7nNrIWbPz5t7dUSdg37eMvnZ8pHJ55JdyZ27HgzXikT9X0cGXxGZaSkCts3/Qbllxa
hMRU7Dj1F2XEYnaQ3GQMYM4S+nk5q5VouSyD51yheJIxy8S520HPpTlObvpUGit95X756VGXyyoE
VMyn3yUo1yrr8FKtuAFO+Ld+/5V0cOzf8/UnTV+8DgOorVZ+irrBY7PTEBFADfmRqFGpNcAdJI+x
67EJxhCeTCxunKJG3P7OdPVJfvB6CveHRf9nXvLpenojNOKJrR+7V9ok+6qQ28r2lGapvcuXl33u
cE/ca0AqY0+KcJqmVox/qlSw8kzBR5BfEHMHY3Q1yx9+9OQ4Liqe7RVMX0GFoNoqz538Gx97cX6s
V+W1Wy3DEGcExe9SCDmMohqXjJ6dAvTmD1J8GXqmJcM529wCoq4cQ5U4Cx95ZxYRgcxFvZgjBk1r
gIfF6r4HToiAdtnkoPpIqF/TpiY76TjSjaU2Ni/fPAs1aJ5+bsmSicoKCJ/0zd6LZq9kEoaCRGFs
0IXUVE2VVERGHm0UaB+Y9JMW994/Bw4oeFQipvTn+KBHZVIG8poDwcTa3WJmjt3PTV2OJFKbZ/2h
ote8wnOKe849T/9dzrb1FoP04QornOXsgzeU20RMy34e/+4eww0QAnla0o9BNLaG/Oxt/t6usl1S
7HjJc5vBec6TPysVKmc7ncXCxVEZUbMVrNzcivQgyjzw+1JbouifTlm+P7hOfbU2CYEPU7c1pOma
5ShttHHcKuZvc+vR2Dl6458XGgJUfA043CDmxbf9A3WSOQRDRMNFaSV8eOhQhx/iv6K2G5vu/wS4
XjbBX+JjYWX9RawcJAn8QDecxXuKcc6BloseH+Mw6Zv/fXcKZkyuDYobL5IsPOvBO27lUKA/SIoI
FbWPOZqP4BoTcI4YEq7/y4oRHPAU+UNyx0ckygrDiSheQIMehd33WizfRIL/LNmRphWVt19W+UtK
yWUU+ZMDovDiqCrlg1oYc4qciXMvxqR/KJ4/1LX3kaO5IemOCmWX5nvx1E/We01n/tIX0oqUakaY
HfEhQcJaWqG84GtmryF67zdhYmxPZ7p2EuvK5glOyCAOQ1ujs4vVI+Q/I6BBpoELSgfV60BdZ2L0
7zeo25IVHGWo+oPdx5IwHaW1NG58o07UIFmiIZsm/exbEdqCLXrXkbvykQLh29EepODNBSaCEMf2
RyKU3EYV02x+Q3NbwooQObhlrNhOb/n/EXT816FoQNrcc3OwEMnWYe37rQkDHx0CVxqLD+UqjjI2
VD6wHiCvm+1Odeogk+8UtidYmYcTxWTAlj6hW0SavKLQfjYh2wcfME3ii+VzfhaWIW9ISD9eNgZE
Navc+GHMsBEwhTuFuBVkpHTO87NE7DzC5JQ34TGyoWxUCZtU+RfO0Hty6WuOpT6ChKsd0tpyjulT
DcWMCHd1ZySYTEYIl/hSdm72nU8OEZua66xxREBvsaeZ3Fwz3in+JsBdT9THf9rUt911/YbEV/GD
xhEbGrE895sBbIAsK20DNWJxP8fdIXfihAMsdnX0h4LzhRWWCsbjRwu6nulR4aslF02LOGhomb0G
OYT0VuBfUqz6sohzzyQeFEFDhmh2hqZOnLrL5NfLi392u4ozo4CGB0VXrJYz8Sn+vLlSFNpNK1yN
pJaT8JdJY0dVQ45aD/O7rBTJdSwpRqzgzny+KWFYq7rbK+zHo60KHLvcldcjI+xTUrgwXTbimObN
gkJdOEuKCO2INsyclgpxqZPF+u1vwZvO4IoyfkvhsDIElx5e6QaKfPi5JfZfKjj1hCAFSO9Wq4a8
hxYvayuwerSd6mr6xjRBAY63mhVQGupzkyNjNSaDxbnFOiJSkFsMlAX67j8ue9pYW6rahIy/dfTm
FZTxd54seilE2+2QxzTFXtUTXZoMt8GT63c2wQcE7JBhjRd/PPjinBkBy07KHeWh6xRrLWIMYMwS
4p/GnnAVaSIRRFL4cq3TiUgjhoTFTI7aKVztAt2j5on3/kYBecQDsCKQ/T7TS4oUc7O/ZU81UKao
vNbfPKydnayAYBoNK4Gxqdmf4eL1lF2oZ3fLgVPuAHEH5k2LnKFDgPhfZ9m2Q6q1qrDXFlGsDp3y
hD4jIDCPNsQutnbCogneAMGd6IKkdQZgTtdNeTZoQdwwvr4jLygdKhj2SujK9EHfi+N1BzOv1Rtt
BDdvYQZHEHAI2KxJUDQ1Oh7GmPD5rn7x7esyN+uKirldz9ediSk9VJ9BlhQE7w1YZCm3VtKWB0Cp
16Req3so19Gn5x2oJQl7GhWePHo45Y/rJirwrqVE+8sxQxWtjoSYnYKmB20SZfahQUu5THIW6xxl
2IrFxCg3vvWbpuoHp3F1IkfvLPST27MDSmiIJWboS97P2BAqRjv+klNBMmtrJM7BO7WM+XNTlCwR
qz710ghvxKuXob6NCqp7Z++DMobze/jt338Ti1q/fOy6uWsIPUJz8I6ejdhnFNKKZH4zviu7jlKU
ScV4paUaqZgILsqVosZQeVrkx4keqDlsUmJwQMPUatLA7FIhsngXw+JwQyBtX01f0a1wPCsxPdE4
0H85jC1EaPPSSCyn4SWyd/xT9sdSbmGB88Bu6ZiJuHVJvHPugHIZHlXKiH3hQCcdtULax6Un5nHb
8elSfqYj0RHZHfsUhsfmhHJGJhhCFTWyOBJTvwFB5VZwzLzSqivAfKJ9igFKnDbFrOgZVLKGl8a4
f/7z03I9IWu8a2kA0gfoHgCqWwbyH42RDVIyQ4mEXTocyE398NUpiANUbJHsgyHrA7y758pDkg/F
AAEVsflJvHWucD92rycoolYIjmvVHKAbYq36Rqcn4DMnNdox1lZMyYXkfYp79/PLitelLY35URnF
U88qvnicEy24nE7+PA/4vBDL5FokfZQuvZffpPnDpRgSQl2cx8vUo0HWMvsVrAe8BtgPiD2VA3bg
7+dZs97Q3Ao6m23Q1Hc7gaJS9IOTBE9u2kUWsq6kFc1+tIi/S6p6uJQ5EBBvMJz0jwc/W1qSE0Lu
ryKYIjP6EmG+QaPBh7sR65PrZB8NfMBXsWaUIC2fZuc7uR+G4r4EnPZxSYs4BAQHmS6xrhCUj+oH
fhgdhG8K7PGn0DALJWvg+mG0fEwWqW8RBEnlrSYnPo7JiJoevrxmcaaheAAqonZzEFEfbPUuUdLN
02NAak4PEoLcDwAJugGt5WkTbK7mdb75GTK7oOwH2PV3GqCxjNvtGTwICD7z58OSnfAFkAraoR4d
aG0icxK0S69yzb/r3vs8F1OaXQ4gr8Cz0gdYa4/9x11o0BsLg5OENuM44VeXyUhDTbaItF/0k47s
3Tb5ljGjkLZm10dSsKVLQNQPA0wpiCo2AbD6FexlbupKgRRIqjgjufNPI9LEjBIJw2o5/9pgY0LK
DoGXZJWcSoi5Cw8wQhm4PsoZvsqoKc5hhjZkMYaszxuxJZpoVYiXytPxszec2xtWHvtRgravG86N
NWTxhrZ/m8CMzXE9e0gJ/7sU0ChU41rJipC5QLe84vn8OPf9zBCAIqobFCWggDkJXpt0GLzA3roH
Z9UfFAedRUEbvc/8g2xNTSPYXdnZf/NOu4f5Aaoqdd2Zj4AmFKBIrQiticFBJzu8nm18iJ+1NSTl
TkRRmOTvCaYhO2TAO1e2nkFgSx52A+241WFPVafTU/5SZeoLE81+pgum+TDdYVt8GVL6JQYk8+DZ
TGDHzkib2ug2jLiR9gAozbI6+4DgCA4Aq6kSbHj8AyLbRKDWTuu3NhRAJ8mtK70qc9Lyc2zpkKde
nsTvvSzRhNN0To32G7n/DvfSk4ExGdmVsg08FtXG22uXga72GNLsUxj+e6MrASMmW+UMvE4Uu8KH
4lsIzSH+5f/A/5VZzeavqCb8gQ/iMgKwOxhPZcaGkoZEDrYIFjQJVu0umd7i5XuUM5Qi3qSj4xoC
gIN2RiEWjFW4RbNkysm5as+RjwEZdvmLd+qr9kjaUfQ0GhYE1/d2Ait/FfCwQFjItsBPyNK5y85i
du8X2jngODnp0K6CgnyJVSuMsA+qFJfCW8FaUOgHd0SgyQtxcCsSH8Bnk1sHAGwjUCbGRkUilGzz
LePuywcdMO1XkqwNpVMwvG6aVhrO0oyIEcjk7xmAvoB/M7A4jdQFbbKIblEwGkFMjXjngeAHo61O
zUFGnJeWhaTUY0k2DSSs92fNBi5TFw/Mq3t7r0DCRHwvLajsSpo2rdhe7PAfK69+6sKiiMYKc5M3
cA68Vsv2odznMDirDsv505pP6mXQDgfa4PN9rarE9geKYUNsK8xSeGIUZBUxdanWAwSp7iNPJ+s+
X9SfCR68S8KZMAftfZ3T7AaZBbR3RNj1gvaD36tdg2/0fMuTTHZCoM+4YCKTEqFr0NMX7zwpHTiG
K+8Y6AnXyMkEC7FC+YSvEO29j0JbWFzxaUH3116dO6Zo9qhUWhplCF8rrHkYNl7qna5/Wg/sfJH7
Knx7wZCMC0XhX5nGt5ovO63xXPmB3MaH+q4SUhW+Fejf3pXU/TOH+wxh4GxW8kaVQGEnq/lBi5fz
lPvkSE9ij7zsBUEQ+qBwHCPpV0Z8FqlbPIfavgy5Rvanm+XfkLXDjS0PUVexjaYboxvCYbbFyvqZ
H6qSA5mBRKpeT26fkTJJXiDfudg6Uw8PjFjg85hUDL0yP5E3WvDAGOe/CGQQCZdVVlhxLRs5+uPW
GkCFS6rNiIK8DJaFhv1lnPZOM1XhU+9GlobdD9kApJar1n3clf3G1dwHHkOTOkhpKrQuwPN1yCfc
WD5B3nEX8iPh+/5sdGmB3fSo4wRUT/yBCi80EgZ7QYBWYe/R3WmqLvOTwa/M62HPz8CQsDXcxPEV
KpRl29SQNFrDp6MHARQ6SoULYLjhH7BTyvragdD4mZ3k/w3Q52y5fb7eZrlDm76WEYHTKbomhQcW
X4+x65NR760jzfdhU3nKXAOoSsFqhgwI8pCD1oI9KziVuCwyIHR4YcK0aDicdpL8zt5Mt4O3w7BO
4HcTlxzDaIeWV0Q7ZuT3zdmIlK/UoiDjtaD8/dqFnd9V2JOk73WsbVX5r8XLBlXwEq0acYbiEnd5
Q3EpSTEbU+DclZBLsTgWlTcHbQSs76H5O5D/Rk6PYz7ITEEMAFaHFWfw/wxqyRS+64nw5NWZCNNB
/Tdj/EsprO78NyxyHanyub38rY4FB7RIP61Bv4EYGMfO40eKPVcApZpQHSzQIFppmOTiL4P343ao
uJwn8j34HiclXsYg5D3wDSHwBfWmYRTpKqBGnqEau3i7ZVlbevILrtQFThdbTRZhhJliXVKU4Llv
jjzwaRGk4XUeXAbuXc4Q42E/0HrasVmQ61rTAX/uEU+/+vRHOqJAHHSZ7W2SeqJhw0wNXEavcFTq
3iofJgygnTrpB3OWSHeJGdCYqYLhvAA78z/5+orxr5fmxTNjT/t3MdhvYtnf+KJZ1+pTn6NBbJML
euCNcTOZQ6Ec5V+EtLmkiEc3NLGXJZh9fytsKvhAtjpJj3lQDtWebsxxJkquExJs4oHQtviOu0je
0bcx6ctNib711Mb8qJl81iwucjLFsjSwXPpazHnjjJPynIcABW3GllYhwKiydmL54xQjdX7ZWQmA
fvjxgmNJ76tlj0ljt9LEz5TeA+I9ZDpYFsDXjj4S/5Yyme8b2dWjym+3cb/2miuUn3nU42Ee/XLI
NUSNz/DA6772h/IPv4wr4KGVevKC0jFekRfRn7wcfMLR0Q4/dZv4F7wynNJeGzg1oMxkdkmczNh8
kTw8aw1KlTJ//fGhDFrpgIyDxyWqlUKAv3VygQiihINyDWv/QZeDJlN1WEbEJkgqQ3JfXPwW/c9J
31YHBqU8gW1o5faS1inWYPc/cdfsT4tT75DArpIypz8w2J1nopUdFFpWIF9peIrptMVaSZmk++Eg
Qe+wriyfKKSm+3aSjAtv9mouvcgzftHQHTDDzTJyNLlYPv2kAwLLRrqIjfXbdwbIyTdb/fD5wiiP
z9MVxRHU90gDjPPnxvCkv0Flcv0LpyImjGQPyKQMywn7YJblmWPLD7GtQLAt4NrCAUHD4Pid0UYP
/A1u3CzlRc/5dFeOa5xp2JsOKFYPmPeTxiActpCNrdhLhpez/yKk9tFiVCrR4VE1w0mL6Rh9ksrd
X/f2ygaXxRHF6LAizYttp03z4jhPl3Xj2l1DKhdD3rleAOOW0uUvUj5hvQosCnknRcrd2EJCwzui
tnVO77xJjPfY+HASl/LLC+JmP9Hh94ZsttYSke4cKXvuCD3hrphjW+2Nnt3YeYKPAkSZrjHzpCx8
SBBeluA4Mo5/nc5PQLbBe/0Z27Za8oT+Y37MlF8CWsWWxE9q0sQ9WDDpwXGx5ORdnhr/9ZNUtSvP
+Losj+eoi7OZ9LMdXXQowxwAaIAM0dzpAZHn1ySTkoqRwLPwAZZP/qeQFrnyUOe1uhoGGjdHkdPC
Zv2F3x8ZwkfUl3ET/HRZ3EPhOkh7Wlj9iefQL+HVYIbYDW8XZgrdRCszdZqQjQEFAkbi/cPRHLsh
qOEHUNHZH6h94uMo0vCJVo4TjyMqWpsxWSo20X7sz1o07u5eRSsR1/z0obWxNelO1R50G5uznC86
dxUMVI58oyYfi4aI7d5vbcUBoXaUJshyS6CYDktsl+0y2qVFL5ZkOwDmjiYGZJfhey6XHrfUnKGf
bKgiWKqLLqyy5Smbp4tX1AfHRGl016ZHC3ksh9NKfUdTkb8NdZF1Gp8cIMLyhRvMSN0XjNUheSly
L9NVi0J+jpM+hbIQc0z5UWjvIXa0kXoF2eNaJ53KYdCTc+23KDcNPr0Kvh2kCsBPRC4EutC3gEl3
lHnJ8ghBSlySirXKb0iE0vL3Ysnupsd/+LayWx90g+5abpPaKdRNzx+A8xOQT7bMtjnaT5oKB4VM
lNJu9ezfxvsLt99GkkJ0YXGbKGYRTyFhEdavN3URR+t/x/EhKL5x6eVdJXjhlHx4QrDgccjCweVk
+w8FJCXJ2Ms/LxT5yLE1u6GswVcFegvQqfUl/BIpraiEq1Tdmcdt0UNTxZXo96HyEn/biJnIoJBX
5nVh4DOTYxiJttXJZeTAfwZx/QTqZLzcGfuYM57uZuyBLTKxZCP9NyP2x7ejaB9I2DedBz51rNPD
pIozcIBcp0x3t5dHkvTh/G7jo+XBqvRIHHY2JJhSXWPHPFWKggJsSPKHbYE18gvBavwK/NfD7sIr
Zzn6Hxd9KNDF7MosYhHJ9MreEYSkkLfG41+0WUfU1WOYoaEf6lXVnmvhKCSqZF8YIQOlQe7Aubw6
6lsczugxbUvVvKPtshGR8rc1+hoHZMjlWTcnpBWlLiz8uK2dm4pkui0pqx2oUC7GThexkUNPGLms
XjaGkoK4Rp2zvcBclmzoRPdw5MMqpdmo7Lg++4q5mrlgr6N07b2/2rV3fi0xfEpK7m6qOr5jGOHI
JafQCKHBk2XFIAq/omdycggIs83VG6YXYH9qe4frs0g30Gjdt0r5TNr+fAs26d2QLxiCfSbbrCGX
k0pRZOGhZ9ITrnb3Coo3gg730lTxCmBhHk/O8tIgSaWMmAtUFBfdENNfAk92X1dG/wrybUUA0fb/
mijwCAnFRQ5QtnAHD6otICzwZaTdzzUyNXPYNp+Nc0PflxOP0Da289JgQ4edV1xlx3y4/qRNW6HS
gJhGLZCL0bekAy5kXlb4binKwqP9Ev5MY0TXqfdyeMW5LLlkovNOj5sqQReufB4/uH3+un9iVIY9
oJf0sUwG452BAfr/APuTMuY3IQhAtD77E6vOsZ+tEeRIwnqajB2+D7aKcM7qQ/hVmoySM9j+KnJk
jIF1N/uu40WjPEKbyXsnZinwVzZ1HYOFqdpAzgP67M8uMHBKm20dZdrFndx2mxhCYXvFJJPesjRV
dih19qzBHGcTJVzdkRYmk31xTRKW/HwkRAXA5M2326v+IllaGdiCsT80j1rdrBUQQpx6H17qlz/P
8vMsUAGxINylXRxDb5fkqEDxGgY2JzO45G2UKwURWhSA8oZhfKB9w/h8gwcd5B7xYJWm7iTNSE7i
xSCR/d0HD5eew/vM62qPVVz1zobURijVVIgGcbtlGtv2wjFbeWezCjMkZk0elQJpABMiAXISLV72
fDKtZ5wS++eUGOCZTB2k+gvbnLbXoA15WoYg798NED8o67m5fis6639oKrwIOaoYeD50FjyZs8Ki
p39uQjb0Jbf5PmKAsFx5OVeu7KwhhbkE52wizgSoZLRCYmAd7KAl+38XcoKVcxX+PV/4CyQf9d8t
rmdn5BaAe2l6Pi0tUaAUBNtXyLYJT1WfvO7xTYY++2xBMz+NXqBTV78VK64Y0lfhQvVUNFs+6A+x
lvcMHRgxHc6FiKjtxHVbERpEJSPvipRnhdmzhgddVk8cEpswAKVIVR6qPoScx0g9HYt3Ixcs0ZsS
y5b3wPzvlFYWgTSGTfmT6lYLiu/6GBX+rKkMsQKNdxyIYqKqZkX5AMDG7r7s8+HIbjHrVOZFWt4z
6FZ6Jn+K+EtfCyJ9j2JW4UrnXvoAj56RxmalAkGtfpgJpghrkvHlLHo5NJ9Mjb6UKhTjryL3rvgq
fi1hgSz3K1/Esm5LCACNmoecviAtmPplIpZ3FDOAE0kzX7w18MOC8DxqBEXcJpJn7wBcwKXJdxOL
0swK3leErmqR9dqJJS2W4GJVfDn4tB014fwh12Z3M5YZw3oBn4/o9k8/dqBLN4EkMRuH696RbwSM
SsYrfi0kZWQoYV+GeC5hQSPDN7C1+kwfH6V5zDZ2AUnCUjKjL/yN+VhvsCSeAHpbLvgZAWKYrvn/
pzSSGK2LRzSMGgiTt6mpqrYjqnD69Y2ewvqnRKtjad3UbWJroBRHaCZEYdzrC+vY4Lq85wm5g9nq
fVP5+11zsAeR3ei8WIG5OvG4l5wH+U7MaeZI9Q/sm0D6HHzP4xQZqROvCxq5RjPd11Yo0KbQ7nM3
2qQaeBp8nkt1h43w20/YCPByb7jRc/0fB91Zw5VdP5/eaf//jUq9PF8JUrIxSX4XlEtDhO8iS05o
IvTuM73OgsuLOOO0lF01p2Eb7GIsZf88+Gy9GxR4A0LfmbrQEKBs+cNRgSp+Zq0s6jqwg6zWbu81
30v030bD9zlLkJldjyrY5tTbPtT7Q64M7q5+0VSXDzgvpCVD1oBznFSSrDQaXlMa6iNB+HkSx9nt
ldUJ9jyLuweqmmGQ+Drfd2EaUHadUTurjSr2UBaWMeBzEDKIz2TczwnYsKeKYsx/Blu4EYw5ll2Y
TsO8R4zKmTAIvpJLOUjwzolOF7k9aXgKpM3PCELrToV6f+ALr0qEmLZyJg/0DMYa5Ur6VTrx/jfD
7pUXtm/5cZqxBWiLpL1cTgDnDnNvTUpSg32OJgT9ihJ+Ye6DX/891GwJA6F/DsDs7v2/G3m+jQV5
dZ2iyuRRx5Ul3x7zdSI7OG6yEF4KIdFIMqqAH/j2uDLegvnyYdF8dRUv/Nst43neldGr1yoJRKsH
A6jRPlyuU/mJHldwi2Jd++472iyFKdpUYTAWINcgEGIjfdFkNqJFozLQPa4DVMmEVNj4jKqR3Kch
kCfZf0tfliIjEdj3ILi6Fx+gtDPH7v1+bSwC85fF1viCqCqHtmVLI+cJDKKJWqjXXiyWBK9SVarJ
ZrgKGiqvRupKJDR0YelPi8py4n5tjzoq+UY2TvVp5UQ+QMCBrmEZpiLYqery/ZGupyO+aw4VzUG1
dKTDOWO5I7R2WbJoLHZOBcjYAqJvr7cNyCElsDSa7g2WFzs3LigyKozlH/fswhxIZVrhpbOMHH7k
NX5+nTm3T9nlwM4XhvHJpxq1vMoYqC7N8O3EeFuaa1/7LGvyUm6B10ynKgsIA+v/to1NoWFWKR10
KPJrNIS9BVIVZPHeQF06/IDDGCH27CFBV6habp5CHUomsvxcw2N6WNjuMbN5xIIvFthJyb8D12mJ
KTi1HguGEC0wXB2gGBKMpNjt1ubesypydrTNYUpaXz31U+GWS2oq3U3hJl7vxts/JNC7tI2Mwpho
inIVLjKwsfJ5IkCHsEmVRSP1dlQnSJbkv15j0XwzMYDwogCdc0brLRIj36ZkNGRoYqca/5lGbwea
CblrI9FkpCPNmJF/iaNn4eRNqrJJ2MbbpRO3nxPp8xQLdP1UH9HhbT+Z+JFDKEUkDVArYJG+UjYN
6OhboU7mX+2+t9YBF5inCkaCLo5/r27Z/bygzpEnEdqXHyCG2SHkKDUq3kTHkM82xhesYDaL7u2j
Bd6ZMy+yk1f3yfTK/4SdV6ZxMYIDYQ6N0/txn7aI0vGKFOZ1cJwa6Ocw53DvDLK09GLXc40+oARk
wsCRRbaUn09Bsw7DooN7eDB4ZYWd84MrrM9pM2jDgYDKamAMlAwzlx71GhpDfEWH2vKdWGuqRFiT
rhOZKBEQNIJNjDLGl/xxp4rUqzi/pXlVUdF0wiqx/KMdIEJLEQFSGJki+sAFdKkjoi4ZgTQtlTwl
V2M2JL/45QDDIbvT5Dhmnb7i0zSx/Jvk7YZi1URdhgiaX/FfO/nQ3GEsDH/3JF5Dp4NRysnRiNQe
F1/r+mJw5157K/RcP4XNjWvwI06lxnjqnIj8wwWS2uLh13NsyTy78SwZMMY48b+l1Kf2UCFAPyoQ
ZjuUCDHTT3NefuSEQnZjjYgxp6lnSe6nrvdBFDPn1JKxQe0dmbib2uAw//ke1vo0DK1XkcvtRw+j
5/lZtdIUiCqAPTEw0Bman5tpmjW9Dd+uUmtBnCvKRBMVQxWuHxgfnJ/EfP0KzaK4R4+EsjPmBCMz
iXU5Q0MB2cqrDSf+yvWOfldOLBHGyt7bRwV4D6QqtNT58H9OH+tkBe4+nhw+NIEkVkwRWCDT3Eik
poC2q25mBFDzAnayAqEESCrp6Pe9B9QX/vY5Lq+NfZlqZp1DoCcQ8q0PZMPAWSsx5DrIFXU4P7qq
iF7ek5iRmYA2BSm25xZWgue+pCNgeNMBW4f9IxBsFGQ1S/PxPw1DZwaCTmAOaJ0MCFAsuYpzteqF
OvpIlML6r/pdCLQk1DbS0oavfK2tNZldqR0o0vS/crOvROD+WoJqfPOf6XpYaB+Qvk9QPUKigLnb
JghVVXCBCIR2tCWXhF165GChEJuz976jyr550gq+4WZtTW4TF14WTW71Ianfyab75Um1JJ1ToOCy
KFt5hIN1JMoPcJkt5Y4BBJcXPUY2ak3JYPj8lt26owm5XW/SLHwPW5jwKSX/6XZvdRcRJMIELk+v
+cayIs6BIJVFFAhfJYOl2yEWV9j4UIlHmCAE/ZoBVaJ1cIU6VOqDPm8/2it9TxwH08BY0fySJxKk
zNalqfZWRB25iez7GqkODjhikh0WDD6FuShFVcFQUnnmrIquBDql2V1rgkEAdiXrx96bJZMirgGZ
yZ2b8fb47WEAnueQu2Rz+EmzX0+cygm9Oh1z+PFCOxWu+lQZzAakOCLxCFu9t0eX2o9pjmALIJok
O3JZ4IkbPC/bXbCzw1DEMH8k2glrUxcUlzgqSLcmAe5T2MIIGAAjvD084040xvgsBBrPW2sqfnaU
SOrcglxbs87byw5UeCpwkvnOGkMCVnpnFycLadX9mDXcr4bpADoKmf1IZWlTsIcIl07qly80+qRi
BhSrUWf0xTPYMB578fglQz0tB+7xBwvpU+p70D06YJ0UwoT2l9ZLEYe66bdWAU5QQg9yr8wl8fkV
FaDDPqhvmhZziSrSvBLCols+Kx8egYFgqH0yd9d/fNPtY9Ub/KDa0YxSXliSt1/aDnmhwqCHdBIt
0gA+V7Ssgx9D92gkjgqt79vjpbbaqu4ZyObPB3/gMGbfsS4PCdtB+l/dLNWs/1RrRPO9vkBn7Q9h
sxn1v1JQwJ/0I09Zjn1C44/2Q8nLdLwqTOGWl9YDU8nAfwYN8SfNkbt/0+HYLnU6ejLhdUtKq4Jc
71zmkfo+fRZjFswcvGx5EvKChEZWfbuAjWygYN13fnvjn2K7OY5Nc5gN37s7Qo01bA5gHeN9LU92
d2jhOGy0vmRVdqk239wWQWh3H8k9o3sbbIS2jAPj8dFIpfHZ96NGc6tQzcKsyc0uv5JvcexSHzJz
8CXOj7sEYsfhkrRWuMP4TZYuQYfxgq4Zt11eSRVvykdfL/kdqyVEywjjOeAOZGqRbZDYUKQ3d+0U
nUISMhDozcqdb9hnV/tTF+wxUo7SJUh0p0RPiT2YWSX3cKadKCrGyR/36R5Mt/W5telG+rOGWJ64
SA4q87eBUTuo5VTapXwlmF1W0LSKHhrnP1QXilaCfl5MHX/BVL92wCQcFOeNbtNTryE0Kn/KFW1V
2EBuIEV9cONjJtJjPPtRo0Lj55CrZpXe4va617PZZilHv4sDmmEbyDtUyzp5iDppYKtPgQuTFUDg
2IoGogmoMlVlWxFEZk9G+aDVo+eUDDAhKfxkAoNAeIwtwKh8uslS8fj8puICmLJ9OLj2wFsxgGSH
ciGY0zsWCpeXOo0g7OFIReV/Kk/+XItuSKjT7fw6cW1OnEOIlWmdNLxqdDzCd3iaikRphxyevGcz
Rxvhf9Uw3YM8rF5cR1jlSSnpZE32ckRKOSLid2j1S+sUWDf++eSn1ThMh/lTqI7P+huwhRb32V2D
55d4iZab9ZppiRNNnUZHqc8hkenJCi1KbCGgp1p0R6mUyleoSaGp66MCWBDazrASpytV8saeikR1
+n9oPg6AEvSQTseozZLRLGmsKkms6BCLjPNrtnB+Vdr3I/fHIfEzO5lWpELMh7E1We1HNR6CLHBt
1BGgcYTNNVJtf5nL2W0eJekc4EGQZBz+OIv5OPxqmWSxUclCXM/J+Hp4tCZFF3y8MWeSZyIGI+O7
EcptIhACi7fix1ThvOQi6g4iqVRIAJKZqpATi2TYk8vcjeqsGYZ/37Sp63YPxRourqDoN8tvkpwC
r1U6wXsKsV3Qrdyj3m/dN81j+DIzDE33KPLMUc2954zhaKg836r/p1s1xha21OUYVvXImW4P4sKo
LeM18bMKY79q1Ae6HVo/KX3L3afgvbXfT//5sNl1l+HUjMPz4Lr0wWI1KZ/Hw9vD7Te8SPJSZOPJ
P18fpR7vxNMLY5oi0A+GtIk7tAgkoLTzHnIg81Yq7Z2wRxr59N73GavXcJmn6lE2Be5bTk/u66eh
SHS2+PDWGVLjPHFvStzC6xFeZQjuxF0dZnaPxfw2abO0lbv08M4UAlVJdkh7+J5+rxXJDm7srugH
Yq33c5N3uFKPdY65CVADhrKVc2wmNjwPNx0Gtkw+HN2bt7qUKrGZ7Yy8AsrNN37U2T79YR4dU6NN
4brCHnMPp/AWdzrXZeTh8ayHs3EIp7CW+kGYOalZL6kGVneGt8UFoXAYLWP66rXFxJ9ZleTp2h+4
L+MxcPLidArMNIdjDN+tqdEl3O2t4GE0htfadMjC/ic88XSs5TamDvk3D2ebxXLGD9qK1Mxj4Qp9
ux5/nm4aSFKgoJJPcOAGxn8HAIQY06idJadUgurYlTIlZsulf8n056HooLAICg1t9sfJKHGFMxia
f7AUtU2KylnTu8aykuVJHZ0fx25fP5/cbYbZ4AsajK2ldpkY0dPy4HIIMIjdwWhpc8e7dFKO0bq8
/l/8fO4rsw+3h3SeRjwpArel4Tv1fj2dgdQbti0cMwA8ObXW/T5cibWw7spfhDT6iqGH21BfbBkd
TqV9wxsaS/VHNFEzC9EKVKZ5rji+yfZCO2oAXSSduu5mS4dGXRGZ3lvZ8m0a2lCQ0XjlFbdzRV+c
O4wQwKCreWmSNHTgA0low34ECCIbKkGhehpxEiqnkPh3jYTrNcj8kGbHM/3Jc5y5g71aaDrOr3cu
qEowmsNwoMlunQ6OIxPSrpa/8+h/BozQEy5l5JKo7TsfPzImwcJlrBwdwPfC2SiCXB/Nm4noYVdP
7GEF5GB0+p18ui3YkkhC2Nh1fUCU8B6gUaGarc+arv8k1IIp/i2NKvFbwkpvre9+4ssIaCb5b2uy
NDMCgxICsV7UnBXkJJQSJR3YbsbVzWzj5V9qkuFA01baookDj35644r+HH8Tir4dzNsj/evsYC29
Snh+CRfMyEAwDWk9jXMWVLj48EvnOFYLUw7ChDtSe/5j7hvYfccoKRJfytO5NRi+58lpmxejjUPQ
K1/qgulIm4NWujGomuAiRgKscxeeRgzvPY2A7wB8CdlGAqFj6gmOiLrJFHxoW+9h+xWtgFBlftas
Qpv7OnYrjjohb3/rxUNSiBPfmFYhU6heywPg/R8x0FzXYM9O6a7DOlfCtRAsStRP+x+FNAMfM6tD
5rorKwXuU6QKiUEQdNIoIqpzWkv2DEYxYeo+QYNgKJ0d4oNi9nIOr/UfVpcVTPX0URwxM+zqaraL
UhFugEqZwKND80m0l3Z1q8/qWuZBonYN0QDibmrtCBWQX5N9cVTgI5zD+h+OTWJ/+3gytnLTFWD/
X2XDoJb0eFXDZ1JETK0+HPMisHEej3Bbs8FCCWl0tYM4a+Vxmge/YFpSCSZs7XYOGCEU931rbGFg
sCclu3147mkl9Db7EvA9JaxftSLgpmRDWoCQnjfnLNVS7+4PXlRxMq603wucB5hw03tYbGmRZJg+
mi2qHqCqWlg/URuZGb71PORVux8imBBXaw5wqfU8UJBqzNU3yo+uSDUj8uL3MRvq5Wf6LM7txgco
wc7HYwtgLvFSV89zNrVKLcHSwCZ9d0oQfEODcZy9Xhx5R+Treys278bXqvkPGikpnZroNTirBClW
goDDnQ3k/jFXWyA0a0oh+5IrcvLYTM5i55d4Rirxc4PKFO6OU8Zt7eELgZCTsdTc4S9HQz8vD+/Y
uz+V04PulabArsnt9++u7fQ9WShw8HEUKKHMcc1Wg2EnNLmk7EICUai39ReWOPTZ+s+ClPpFWdWS
WNplES1crZqmdCcqlpUIXf2UeKqBaLEezjzDH/squ0yNQmP9Ysurd0cmV5ueV4Sc4AYnu/5/DWX7
yVJ+GO92uR1G6p76pFdo9aFJP2TbCbYGzJQ8fQcaK0d6X7WBMb7caUjZQPX1Y+R7+oM1cMZQNf+m
CQ7U+Xf5hXGA+qLY45z0cSHbW7EcdA8mV4owCm2WbhB8+yKcie55EMusyWF38wcmeV8aOnuSVyEd
yVlEnIOth+3C1cRSIFB91SCj5klj5hVBOTggdegNQsUX1rZyqsp+DZCdL9ojbFp+FgRi2mKNRHhT
mC/aFFkIUuPLGeA8+9V0zrRhEnQkbPfMXeof/qThZVAj9rOHF7p5mck2nGrhOg8HQ4d4q/MgYL7D
kXBk437iMefUNGns/xkA798APNKMQAoTd7VxUpw6GqII04qwJVz3ez8vTaQlah2PcoQbOzbQeDPv
LABZwdr/SSHGsUzbRK+Sl5JcgGG+il40p8ajsb13IxIp09/u+m0dLIzuhtRnZZO3WYjdDvghsROu
WDsKCFErd2CpNLyxrFOY4+hQV6UF9dmiXD2EJbRMXXWx01gyotW2pHl2LekxusphKzAWx+4pACwr
qXtLxmYGAchZznX5fOk13+7PTvOVIeRYJbK40rPc01ge9pXqd3yaS/3g+YI9mdjoDo2NpUIg81S4
bT87baEvLNB8WLJ4HLVW+dgABIkPWIzVXl7YD+FUjjL8oZlRHesUaLsvQ5qZ7GYFzROFcST0hIrl
2MKibm4M/L3mVZhn2yMeS/eRxUhqpnSdRaQ4NsoXtiXOtYNCN9q7yGVtfuv4f/SuJ65kd90UVsR6
YXHXntubUn3PzGcnfCdYWi3ZtAaMlTqAd2cAvM5rDLJve9HMnGgzCRuwQ+TlCSQKu4K42VyHAQGI
kvwZfC0ycG9Bm40zPLb2ZjK2va9GwNR+lkEu5xE/QBYpFgkXIVDaQ/Z8DWw2YLPYmbuhSBj98Z3G
SndeQxkHd2tmMn8KhMTjA8RJykJveFEGHG2sz/vEITmUmYbj/f3C463Dxmu9sPrJP2BipRQC7ZVO
d6uMfBGW80PCs9DrIFV1k9gwfR/82IOXSjTFYwaY4urT1xwo3wCDxaRFvjMXNidAJ9k7OMPB4i5o
EiLmHNyaJsQkrcQK2vaCxU4+iVbb9ez6EBAej+Vprdo/5ZLHc5DyMtRge0YGM85yNYUpWtZzlAeM
oMOeSIInYP9z4Ahc+eC/fyH0UZykTft8otm8Y1jX4LbPlZENdf7cQG5yn3cmkrb3wJyrvBt/qeag
FlXVXFqvIXMce167zSaHI/4qorw5zvCbHjb5vtjcTgj4VofT0wxwO++FuHZMJNAFID86UP4s5c3A
rt4Pf0l2o1FI7CJFh/hR3K8ffqDVPM0hmZVoO0bxScK63EMbIviAWVMgJwMk96Yj14IZY0IN+KP5
yjuEHf0ca0UEUPiPJhF7je57TRR6iTC2snVllMKWxbgCBYIZWvC/houtipxtvwJYtbHR4UmJx3Sn
xGvpo/Qtl+H2fDI6P1EGPVqC5S3jD23TzlgwVHPeW0nPnbQyafjsjxVI0VOkXy6cTctsv/tK3tAR
SpBD7IBND3qQUBdbvab5bdu3U4W3w1q3sU5AXU3x56Tzw/YNaA4axezchgIKJ1PaigVNRupVzEBI
mHca82c+RiUKjsNq2rB39oyB26gnwWIKTl/PI8ElqYSvYuZj6jPD9+CXLJYrfEvPV+etZ2IOq6uS
JXA/TYInuwQLLU9tPylQPPw11tNqTbp37VxD1BhIxWrv7cn9rcJ/NIUOvF+WTes7CBvy+q8lNXkw
72eFVDmqRMqlGcPa45ChbkTqi/8Si8oNGRFgRb9TpAy4RQWxjiXho94mXaC5x+b1zZDxRzV85QPQ
2PcHPIOacR8zwYUO0gS2KojFCMe2xL+N/rwQ249lwoNzMpGWUv0c0Z08IgUmXlOyAyTiGDJnPzWO
7UmF2UUFDlKR/NixagvInVtC4292HrB8OKdsb8lKdenRH3mXsfnOP2qr0xGtnc22qI1MjmtROJ5V
/y+NyZ/S3m2KAHy57dC1rLrjPGq1PrR2le7aJa+RPKQEiUURK4CXfbIzg3gYmY6QJ2TVKS4eUH9l
woWl0e7GA1s51thTbthgl2BJ9bsdNnzzWELPs+Zu6i+OYkvCGzog8mJYGaymgXw6hEL8tlrioY4b
EfYOiUA0sSzMV8A7CjkhYwi0/3pD8iEEQS0Ha94AKMhdtHtEZRnjDQsMIgktYlx0HiNaa+EoUqol
AeClDegnDWbACmhEolQnV6l3fYNyt3KuduDSGD6u7vrIRRr+e3Iu1/oxB+jMbKw7N/+VIk6pPEa4
CeV1qwNV1YOyVAmgtTWYAPlVXichoLvdHYzBQrSMcBVNLReNYqpaBgTjMQ9hlKAtkoe859rZI+4T
WHMG4odCvY7pafEDgQpI3GZcqUCB5cv/KcRNFAt+TelFBb4xvnw0ff2BBRuoe7rAEJA5A3e72J/x
psvs8m2DKTFGjz37cTWCQBWECLYaxiO18SBknjlegl+kNg3BLOqwM7Zc8HgbmqB5x6Wr+4wNSJCv
y294ofHrqkZGGhcA1vlE9ZH3L23yTZGnPU/AGkzhgqpNhuCLNJxTYsVxOf5graYXXlfT094DCypp
HSVjQPJ90mCd9rddyDAkGVeopBCWkRveEqROr7uC9PHm05MzfuN+Mu3+P692k4p/etU122dyReEd
r+RXlp23yH8lkKQ9S6lDukswc0vouf5BhYcl8RBv2MFItITV6lijqqkof2sdldgxs64ZXcy7GV9/
kWS1NkePXdhRQ9KcMHeoudp+0hPR3dNQa3I5RY1b3u686zElaEsq7Uv6rFyxioQ6zhCLI/qcTtTz
sCmX4MIDz3GYI4S+VDAYBr/eaSkPTSJC3HNsTyi7Y+hqShhj6Gfx1pSODTBhkDO6bGv+QYef0Wiq
3eyusOut9eri+izLYougXixTb6FYx6BzVeB4oU7g8V+xoYWQfzmy4G893fgvjzzioFSTNWZJdKu8
W0U3gbzZYRiQKNCc7Ok1Q+qT9Wi0tg8Rpi7FPS00r7VAcCVjx+bNyCAgkdsHhIrTWzMcAt2T7QI6
MQZwijzPO8Bi1VpvyYL0Bjx2UfvFPG8tS5bqlJNc8UvrJbq3i9RGnI0oXmqHeAhKjX7yO3YdhpAw
/h/Y7sYZ4bQENTZ/TB0Wp97tQFgf+dzX/rY3ruanwKZZWswylpdqiK0hhoY0vLk7Hah6QklqVgkP
BrCDmLVZPXkXJm+i3o6yFp9GmQmksmhzyFTY+yzxk7u/9B+iLt9v8CHaHd/WvsRCe5b4fgFWRK1d
v4Z8RJmpsDsqoluSWO9xt+tISf7vo2aN3vjk5kACHskJ07F005unhYCe2ccrjh1H3tParCYQDLhV
vV3A03YLwjdeu/S77/WTvZdIk8ui10d9dAPPcVGUqxAYNSH/enUePiGWcI4uMcN5yWe2ezE7xY41
J3E0isyk35VH05kqIHwLkEvJzQv0HWwXLcbsc3RjS9o2X78t8y5MZ6x1WYZoDdl2JUlCe6K3Xh3n
lLgV669JyNnkmQWX/yFGrVkRbSlEvNmVXEqb3tW0Nn7NsyncJJxLhCWqj1owUv9zD2PQbY9/ZB9S
FTapHuylIshFlgGx3+/QDE1Xt+Xt4gFQgfNeAPKhnCe5XagReaMdpFklU0OHY5+0W//UigDttdQ2
3t/A9w2hA06Cqbl3ClfoThO8y6a3LK1g+VOfgwhFl90vobe8d876eESDGTzxhA3TgjMXrkFJU+QG
7HUZ07pOdb9gqqsOdLoNxYjILSHeNAJoO7unZp8V4abH8U2RXcDrn8i42M2EdB60fgmR6x6bt++D
bgZwMLNKAwaoUDumm0a6lB3yH1UY4mpMZUwLFg4vRTsqTn5eHjlxosC/jMpr7xf2wPSQrLw3WKZ5
ZFYZVMpbVSAgBsKtTEzsmr2vtw6/r9SrlLaf5oMhBycyFbZ3EjxEQasCrp0SOBfSqqpz8I1mWipm
ZZTs7Tnrjb7a2sBfxf6pdw7YfNVz7YzTI9Z2C36ivtP6YrtxDKHwB7bYWdytefex0Z+DVvL8xmuu
ekq/eQT6d2CuET3eu+b0s0sI7nn2G0TQRHL+sWP/Jxglb9KlpxDEyZFozQRcPTCU/3YDazIfyBY1
YHU2Ivj+CmrfqH01fweNpW42ICwRvaHiQkdBFoY300WnJxzHC598a6XL8z1hvw/ujVqAdZufzQs5
blN83F77AqHnO5GuIIF6zaI0XvSPoPQMHg5SVqn08bh8l1kx34pj7xSRq8sHPdljPXVsffwXwYel
FIzzWB04PO/DPtB/FSTKxft+GfpcPFdJXv0Bm3u3PI+OMzrvwqrqA2iodLikTZa3O06C6B6+zUBD
2At3w94V1Mq8IOUeawERJ69Jsv30Q/nXkFn6oOjTLwEUoIZWlimAm7MQhmZ0TIidXvk/nLKRdkPx
ft9Nx51ntl8IoHNuh4mWWALLqQzq50SKz0NQwnwaZ045c8iRoFfegjTJVDjlvQf0R7L6FGK6H8HZ
GpZSstlNIqIjAat5/LeobPwSKMyWbR72CY5YserSem7BkTCYfClMAko4ca562Df7UBpCZV3be+4C
hdrXIgpb3OWoGWk4RMHD+gM1ZWlzdFpXByVGOvOGD26/9XqH/D/sS/qzMirZwkOdoXairVJUntpi
DZO98PjU+Da9SE9aAGMobIpFbzT8uzEEKX+luhvzacz76+Amm9QkrL60oNnUhiti2WcDNQ4yxnPh
4qeEnKM7zZtDNu5f69xeEbDPPnfuezu0KOj5BI1QXGLiX3dVC40ljGOsmOHM5Rcf+bXagqRex15H
2BI4GFs39i0bL0cJGsfPaIbn1gANUM93DyXx17Pft54wVBVK2N2/9y9VossdXoQ8olqEsOGF40f5
UcSjeGShFivU0Gr4CJVeQH5oYyNSdvxFi3FvjCOC3KbIdxGzc6yzNFQ73KFb/NHBUcLxX/hi/CUd
MdYRBgCNXJW4bWNK9kxulkJu0ul7ivfqME6u5teLVA5zY7wNb1L/XFHE1GYzToXsoCkcWtS3jo8J
p9Pp/gTsF8W+BRbaX3NT4+51yGpTB6LDp0Gtp9kSBlvMGOP9AcbMTHN6ef0ER8Grlp1HAf96Dt9A
wC9P4oyHrhAGZpCYZfq2uLHWPZ+S5/QN5Wm5TndHTEEYB9+Nk3OJ46ixi4wLDWhkA/qqOCwQi4KY
We6nqHWMjXiZFh/okqfWF4ODY2fyu/Kd0h7hI3AITD+CW/7VlvHLKfVOgUKaJfTmW3YFMyifBmAD
FbAiWpVWgf29vh5A+ej0I6kA3T3/ozqNrcYGznc4goopEZrRmiXDhkNZ8nHM+4hPe719n+wS+0lm
4M39jH9Pb0h4tfSMOvji9rqVZiv2zqKAknd4tJSLcjKCV22lXFVXEGl9H1VpDoYJuLbUzNTRccEe
jbBqSHdx6B6S8cmvccdOkmDe6NqmbOWfKx3YW2f1BdOax/ouOyYylGvkdM55o9/oGWBqY4L9raNn
Ej4m758k8BJNB13im/d8yksdh4leWqpfNdS81fTMJuW58bCwjBxjEPNOqZMrPRla+n0ro4PbxcpA
SDiwfNv0k/4goRPBJBsjc+sWUXp/Zmlvf0mQke3SixvWyHcCj6FTgFH1LQ8YJBooN7lo6ffe23Ip
tOCU9Vgsn/cUityGOIbOaSSBqwXOW0F29lbpOTNqsGf2JT2HbkBvYJa5QxLSgWYMLyaAZGJToKQ1
SxZ29moYp9y4qmHu3HnF+yeM/aOkHp1QO9wMx1Hnb4pbavRoFyn83CO6laamoRQreA66/uQFnTRp
3kDgYgpRuVr97FWPaf8ro3p9h2D+PBaf5xspig6vOEgy5/R9HRb8QZTleWl6fRw4/x7DjAMUCf42
TCh3XU7gVmE5MB8VZdu84BczFxneIRaNfXRc+HrkBj3+wEG0PWGN3yxoDs9rtmgofLPGZMpmP1Wq
nM+bx4WqOJVn605VPJ624GMMVRX/nOWguBPgYcTfBfG99IsEyeZwLVBM6YQhPvMtnLL3GI5Xj6dF
rLnUO8POMZxg8TVpejru4E6AACs8uQLFKrb2p7DYyritd1u5oV6+Lqpkb9dspFLL9VyCdxI+ke/B
LhRKh9JkWjrKjNpSHEEVHYCaQ6PFUMdO7Syw+w4f5G+FY2pe7i9C2Q2ZW++zlas9sd1T6NDZ8kiK
kazLrG0nm2DSSx2MirEIrO/sD2ZBx1+csEu2oQlG7rhwAq/0Vpe3PesNeIX66kPGcRThTmExlSrq
OXcrFUJkDaI5ugo/N2vCoC7TugxpF/vHOu2kNu1ZqMaRgssPoi1PZ+DDIFPJTeTVHWQbuPCGlCQC
vaVr20C0O0Lqfm9nGAFP3b+IaPOPWaBQXO6KDb3kEbIlgVo/TuwqtjZqJLQlJ+aM55NhBtdYwwjp
SndMUWxXsEoJ3uWA5RKMeKvweVwFiTgWV8O3dtw1agect/Jj0biTGIsIUHc880p9bCptdowjS1Of
sauzV8uyJ096qMArMX434bXIZ+v2CJkw4PMwjcuHQlryo76s0mpuv9ppr1pArKnDMmR+VAd4KnHd
odGzXng3JRt1OxyWYq4R6IdET1MNlGetZMUGge9hT1bnszaYAlczm+ohAwrG3ccLsCI2NTvWEW54
sHOI56RyeEYlvPJHKohmkpXJihzzbQTL0Ni/XAPO/Qh9NQCQaWKOImc5ONGd6h6/ypEeUA6jygaj
gId7iPPi3LTpKj+n0Wh9gfuLBorRviMi4flIj9zfHRKV5QUvoLo2fGuizmcchE/uPScqDTmxDtXV
x6ZVmQKVDw/G/uEK90BB8qfLIzcBiDZQofuH8buCKpkr/F9aBWrwfMeyU5iqtELBzA+LdpDMy8x5
K1ckNcvHlY/QEXY5Ja922qpbYPC1GOuC7hyXf3Qw99ybFA5ps66UKoNWsOT84L/tbygwwHqpu5sL
LCikIOiCQ7Lvx7kMq/P977X9bpMHhkIOusbGdm0eyjRWtDg68KPb7Yd7raxA8eQGvqsX/gVK1td6
cj9QzqKBA46tWt2VRJ4banTM0jukf5qjkudk6cNK39Yt1v7WWS9sfrQJm6CECWtynQg04INMVOSj
byt4G8EYNhv1zNnYDkw6On1yroIiEPTcWFn/ZmE+qJ6DkimWRdCnhprW+6+7X1A4Ka9OfW5gYOPY
KOG+P00OeIwIPsveO3u2tBwQ4Z/XIPMtcdZVax/brGTI3OLYYqyVNfKDqggPegWFHt7He5cm7tbE
Tgh1+3vChCH90bUs0mGIl2ZylCRqGPt4KnOsThyOlW6OpiJBx8uBxSFh4oGooawZ015f5gBkNBWn
RGl2/UwS4vMpgnpKgOqwmnXI8wIk5lYXQmPGA+pv+uI9RuoMver5zYR9s+Rtm8CSgEfuEHv5AKpI
JIjpDK0QdqFBxrk3sWhUcYBMqSSLWkJUQKxu1qaWMWb9pJZOnQoL+7J/yoh8U+BcIcbbXH/doEq5
fDXwwT/pf4HIn8Ehc9t8RhJBXxaPNmsR7MKEzbe152eJRkoDvRNoJ7SCmegIvOlvpwA1dPJyNQYX
HIBK1FQUj0eWbCYT9rzdGAhzcdhLIIiPI09h95PMyDZmVH3+A/zLj4Tnw8HPB5wBcmOyNC6QoEUs
NbR849JDxGmFZZIu6yR6OBlrUse9p7UcEu/I5X/fn033ChEORaGULyzmYlGpgWUD0UfJY/iE2mfe
z1nbQF7iJH54dtsDgPDg3+uYTEHuvY9ujkizBvmaLgnCydNdoN34xhXyEy5sNanscwgPGZhAxzsi
yvhquJeZbRYNOpD6qABbVxLp1LDKu5+SEMnqCSokYRvou8CWLZH/iY4uTTX/831uLtkK5fjYEByf
cXtZSqKE1WjIf79tmKceAQ9Ta7Ph74g9NF0mCCYYA9U/l533aDJ6GVX3l8Ry0aI2QkwJM6sBpUc4
BPIlzXoVK/rckKdbF0eV1VnxI7GAIrYppgu9OQDkmiqhmgEYcsQAFwl58T00aae0vRK+XEmi8+zD
BgdUI4Etckekpz0xL4NjCiumUs9KXXx0x4Zpsa2UFmbhF6SM4lsngg726t6R0p8bWZWpsAuO8HS5
Ljoh7ytxmRYouEfKbvpx6BnTfCBHx08j4mud6bpkjReYBhrPDKhVt5zUwPZuBmAU6MyZysQQBVa+
1Z+hKTkQ8ZSfYEmw7niebLTmCbCUtuLWS/HA2dZ7Aw9eWPKwJEvpvNBEZKqNP+/tLg7Fn3RvCfzi
ILbWZWfclqqvJEWrPOyrjj7H6thblg0eJfyESid2Y7cTS8Kx4RCKq50/ibIcHup2oK8OFg1X5Rwg
fRTlvK+ZOBqj/DIgN9XPL9HQHJ/klAofoHXO4VfPnwuQvN6wq8IxUb8H7UlEYahAPcrGWvVCZzpB
XlJYEI+exUOd6F6LipwPhhyU8p4CB+dZOeQDrbx3T83neSCVndbKkQc/6GWy3BA00+8DUcqh4Ja8
9t2QDTgV9S1I7cOPEx93F56ttwvGYlQXOyJTgIkVlWb8vV3QrHaX28JmtIDgLpY5uHjHo6K+rugv
xnkRWbMt4qhJiC8sNuTtTyNENOYtUKYNG4hmJn8wAHQ5YxQkVUdHDvN/gf4bipxIqqtfBmroy0zn
ZnlNXgxOJ+ydcfFaF5gOaFQg+iJQpvrCcMAsY38mRCIRlwjuDDmzwtrI0mYjbtll4KG0zFdnaRAS
86pR5dwpJKavz+21aXuegOU2iGkBS3dtwZNJ4qUMv/YHS8yXlTlJraPBxNqhmlQHEvsVlMjJMMsj
k6I/xAmuHYFRi/9VSGxZ5a2ej7HQ0iEJzxJ7zfgPDgNGtUTfBJe8iT1tyCPM76E+2vPP2qcgH8fL
OtiDdZoNLSJNYvw3VwG5AC76bq4K5Uv5miLzcdeFUPS1u7bz71G5vE2HvwA9CVtbOAI3I/YqdR7t
QxFoHMNe9TtJHFYlWaAwfdNhyJlAz7n9GXdR38CkJFwpcPCnkQbJXf9TNC4lpyYNxF7Z3uZigHyu
IrsvKyimbHJgRE9Ip16RD38nvJ+088ix6gkGBwhPEXRpdJQsxlPYXxiK0ImoUCpto4UsmbbUEXsk
z4MmsPXybLjvvoEVNMBmO4gsXVyBSXOZUI5VZyqA251agmByaXybxgdgX+qtsdQgoq42RQa4TO3j
hu3n58CvCYfXJe9SG5Hvl66Wdoy8EYAk2Bo9c12Q5WMeBgavyFr511eiWYXpg/QE9UkiYwqoPkBk
/LHlhA6ioiO5ouvvvWmATAkuNgCX8CgiQTQO7fOu8B+aQYVoC8EuSQ05NYzrrXcaapcEXHt6AMLr
jHG3VqGnNrbsF49eSVpzgoa4NNLa0kEdeeXanJC9kQK0dJtPjskYxXnHk835KKhbUFJJvKPhRriL
Ittb891g7t7M9+r9kgN/ti+W8zfnV9cKdVT0Y+OYc8F7Olyr0XVrjumgi0DaEOmL9Sh5R8BF6iX2
PTVma2xS5todrOwFux8vktqXNmiMafYjQvwqRgyW/XZgVsjWEJBQeDUQvDWZeTIQG5NqAn0l0TST
hPyOQWbvCxSQkWZWGrMwTfVQsCr9ma7FKK776dpMudMDCAG7cYqYB90f29bb+1O/zvpY8p5WASvL
bkliuyJ9cwvx1C8B+ejBGFlMkv9TFZEJf+LVHoETYcOh/sgWceYcbRhHsFP3brPlDsWJZ+shi/75
AZUSDXt1WNrvzBNq2W1eTP1TVSLQvK+sKP6nZ76it5EInufJDTInln/kOuHZbACMXdaiNjCyJbX5
oUmXV9iD1kslmfne2Bk/CcVvtswagOx7KtOYFSdF2WgC8LIiJ2qNYy+Ba5YT3qVeQtnckB7WteJm
K9PAp1VmYEizwev6BuMPvWRJdXmy8FBeOYNpwpNbqq+HoCty/CC9k8WLj1ltYNaSORTwbpweXhzC
kgqeXn1XnT8cxVhxCH3TTumno2M04zfNRpiUJqlot4CKMruqJ18kR2FlA9rG38ux+5CtAuQ5LTKG
h47YcBCbHmAvS9HKHgB1cYkCO/jKFFdbyib2QyMX/V5jbBMG0LayzeBKptsT5F4Hm7qSFNvQIKqI
gXoc3ZTVyS4YixWLNIvWF5v54xkhDdx8DqN2uzUBVkQaJezSnMfTcz7rCuAxU1h9KysGcRb17wYI
hgpgiY7IrvNdv1GJ/79D/azQHJquH34T63eK6mram5WHZh213RPcgxB2fiMxJbNrlEjbb2lU5ATl
NNj5+kntxr6Vk4psJUNJCpLijGp7zerd3RPj1apdRfuwVNVftlcXkgnA8mUtTnJVDETcyq5n/LGZ
M1W92X5H/qVmzTKvv/54hV3ynsrGfkKISc51vkk56SCnn/xrMuC0inF0M4L6YRhioubyFP+9lMm+
QgunJ5BNCjgF+B6MgBmoGh8vCdKRtcLLCdFAGl9F+7DGt1++c6QkV3ZgIneRP+Pnn5n4/gJzg+GT
zn66Z0aCWcJmdrEcmHClwafak7RFjL2MT1UafGPDAnrAHkIIvMTlOrUL0oe0+YMk2BB+8MeKL0DX
VbRII6tfTu1Ly61t5MGHbpeOfsVvZn+3iI5l/nROEDmfJQM/T5L42Xsb8liRUcpBRVriAR3X03u7
3KBFByIbhJJUPM8xHhOq1ig5gD2oAhr/DCOkC9QJfnHNBs8V0Gt/70VTIKUy7JDz/KM8LmbHyABz
0aHp+dX4pGrfeGjvmkfn0YdnXm7XBXMmkq/gisiUclVuElnO3DrQ/JmWrG60URlPL2OyoUbfJeI+
07jOvVn8W8Alep0YyxHQSpCNlfA+7ZqZBcrvRWGmuSwVOOUXw9np3zE/xc+v/S/CemnT8v7Bcfx9
gzdYOZDuSw2yPzrh5X295dcov78x1Bl6M7c5qwVj8zxE9zrljOSCqZ1pMVgebKglvajZ+r9ehdcP
S9JeArdPPeqXii8LhMpPRef2BkdJAAYIHBC50ljF/SP+ziOatR1vAAwK3EyfiDqqEoy65Qxkms3W
bvyuDkjoxQ5EuTj2aoOCqn6CjcRr9mJXMuBmL6pKC+9vMtZRrSbGBUUZUBhrZAZ1SHCilcJ+ys1i
8gI4KalbUU+HFmvH7AwT9mQu99PUXF/GKTheLlgfkA3yU7XvWTCFmJ1Rv2bzWuYf8EU6Ne9Qmetp
iyh+J6yyqAP36HowframmpcggryMWt2Hahlcxku/1fjKbgf9K4e/1u51tVxRBg2x3iX0IcV7ejw8
kecGK/oJ+MCsKSqr6rJ8qMVuuuTuwJNA+bad6VlHZ55BnVP4yT6aLegDR2bu0o7o7fvciF7tO/Su
3QuFFQan3EOs80E9tgyLRpcUtevqdM7G8Pi+hVlxYWdpJZpF4oqYcKldTr10nzBIg/2QD9IqRIxf
IKOGaW15rv83WpJJCxHz0mJ6Lyp0/gnNcp+EwrpckEXGoXDQN3PU1Rn+81f39a5fIljOll2F9Txb
SGBeyGL/zGu/fkMI6uN2BpkhQkm3htMDaypP/NXBO6/DY3zSpmfnhlr12j3/BSJVqmG110Zz9Eg0
9ZKCt0VtZJtgXkd/khERBvCQ506xXrYGmCPh1Es+Wz+8MrPgt+/WB5fCWjKjpsnWp8N69cib/4xt
K1BullzjG5O9x1sAHskGH89yx1RCzpYnMZuVryCZQhJXUIXm6obDqeCxpLmsSwPDC2wHA+AdJ5R2
ejmec8jIU4mB7Lp14py+yn2M8OhKlNJwKcb+KioML/jGf77VY3AsOnVaM0ZopjdjyBAESXzy/aBr
jyTA2MF8XAqh0w3RlvSu319EFiK1Vb+tAp0uzM50MWJ6dxLOFZAC1Y6BRQY0p9Yq8eNmQ33it5fW
VzIGnKjP7wujnogCkNbPGGTLNUMqVxG2EqQBO0on7lU1QM+QZCyRd0J7GNDGdOehshF9XNb/fi/X
jcRZwpIxfdLwWmeEM4pl0ZKH1vcWFrzv6930wXsfNySsXrpgpeu/B2QTw5Vt4ICZT3PFGz6rzZEf
q5EybxIEyUxEBTeGBMjtguo0ye2S5TjrhjyWNU+qtdcQtiANsP+U2gDZw3kezva7WNh0BP5Y4Rc0
LN7G5DnGCSDXZ//400ioM7zL3sJy42MLSk/B1cwOFm5bTz9DPVPfwmR5efRWiIarqi3y9/OixZeq
pY1IHb1zV7xI45o4ghd9pnB2aR3+8YLsQYHC4WeMPbDHBElyEa8xuIvjznkNdRvSRIlvWiEAcRAi
N4wQjhuCCMRF+lqdsfUs3x5AGig7PUPZPxFJQyT7U8ZxnwQJJkPdv1zeZMtSOQBv1cttTd70FIa9
KmJFWotps0VbhXzB/3+pJD119J8BxwB/9Wra9FXUEF08bQs9ZVegpXYJ6rqFFJyM2maCmKOoNF6f
QhQcXbvm8gx3SzfY19ScbjGvut1uaCbzXe9XdsqRvEZbUrgtKNZl7pPXjIMIDiZtRzWh+Pt783cl
I3fhs6QRa7wLqr3gM6gR2qsXMLX8yfjylF8S5Fu9BEcmQ4v8/Z20k23JBYXQbXoDRgGSRQNEM7Yx
HltwuCRSOWYvl5OQopM/LryLBjIjR21+fKZOxukj0LMNpOkgC23NFbeS4gcLtFHbcy7fmag0Tswm
U251ng8ApSLw+yIrBOTKEq05Ltfi0X6iX5gB9E4affRzebpORRNrD5643EB58R5itrBZaXlQM2z/
bt3KW+Ayl4j2mWUoZfsA9EhHa+nOMaku1gQV+9TWaFqRy3hm1oSHCosnv5ZrfW4cjjZXy6bUEyOG
HgCdpnGfA6QTlU1UIBuMKD0xYqy1p6WfiGVZHoC/U2+xYIRcsSr/JEojLjZ9TfBjSLEjdpySRDnW
J4pcVvKbs3yAtPIPWWKuQEHZbwn6gxq/EFiMiA3xoLeiDFwekKh1eGkDQr/wMk8mSgGkiBb7H/Q/
+GNlVfaXE7JFqs7uSQR/AZV5nbNwkfPbLVOEikqM57ZGeAvgYAaGaTiDGz4ew7PCCDblxBgGoF+l
lS0WLIi2TUJ2G3gR6nsY6ro352hTz1e3e2DywAAVOBZyQAyLkGAabop36Mv6Zo+1vAN6fyZsxQ86
zo0qREooHoVjC8kLPQXwUYCz24pl2MdwChXHjqIs5MuV167DRXnT7jr/L1VHaaoUl6HQ/rOM2vU9
1fxKDZTQjIgvbTfaUKdjlfxscmNo5Rvk5jY2hnU2zL4ZMJGIAZ3e3W9jeHRNEZH3MvXj5vzMA8sh
iCjNhfcw3AsrV919RaamHQDx4Ct0Rw2w30hrZoS7wzuZnzBVLDEtEvBp7h2M3qBTUCFyMKebv0Ib
zZxLniiwN20KELHwZoybsPlsOAXqUshwvZCZAO8+CAizvmAdQm90FeN4TNeFOAi0NpxLOfMG2cEQ
ZY9BoOCEAP3Nj1UGDplMlMkgqz05/3dFCR+tcBVjGvb+r7IEXMjZizIZ1Xj7hacVYGCzD8h8X96h
ktHbqpjqQk6jI7yb/D1M2Gf7LURUiXrQ8fILGY9N8lj60KkoKJvfYGz81jXDxrbPD+sBznxC3Dap
8TOkqNzcCXE2TicfvE5kgcPn4wln1WsMAPayvmjkNxMXjPcnfITCTDA2MMIbFnEuY9bXK9OW6nVs
ZgapKGFPWnQ4z/DWHjOZmaikSzUMNgdK3hIc2Jhzm5N/ekfnSTQZAxkIkEmcP6mqTaMi1FrVW5x7
mYN/Jz6aYXSoFnwul4L86+rGlUDORLGnnFDOqWXOC7/WYyNoR2+kMXuxM0AbfkP5isBRlYxcfhhG
YgEULafq6OnKkpGqcVQD/YSUp6RUVrCLSajyBwf2AgAQJqlHDaREMrGzDqNCMIqt5LWywE8TQKEL
Nsz1WmvcXXIlVK1GT/7zCdFpDssAGRjeGs8RsCWcq2XTcOTokYAK2ktf21IETWyQNQ5WrGjRgv6w
xPTaHeqC7ws9lMIqAXSXPYCsw5TPRsEilMnKpo1WFb863u3yq11spWcFLoZKvYheuOKH8aCNx6KB
c4xI3NNYII0V6vMcAcBexj96iIxmtvwOKyy99hH0XrhDuBTV8SBVDb3iyLSiUCJDZmEo+0CaxYIc
zT0QehOnXoild+DU1zln/A1k+PujglV/jruUH0/bxO9MshcMciA4zMDRGUo97IQ2pwv/17YjMqCM
e6zk384IQ2Yjdn+nYy5ZpRRDAtaPUcC5lzkW/dcHGNqd7yHNdEeTwUnv6owY7CPhsKr+185THbu0
FpK1YhdA4i1Xvr2MFuqWIb6XntvvC4RJOqUHhjnMuKW4cXPetXsA/NpBNxctrIi4XbgZ67jmHqt5
xtHr3GmpqDfaqXMLu8Mvckq6bhkYG7QrjAVR4toixlEu7A91uyj1ynE3lDIrnHEs5XzSmh24fVL7
FsTlBmPQAPZoC6xpF97aS1VWU+4JlWsLNsXFww/TPuLu/C/tVJYjnvdLKumiwnzeZLSJ3raiiC98
Islun25gXf8MksMnN9YlaPOcBa9HIfEhKj8KPC60gbwqO1r5sCYQeOlEjpi7VQXls4Q85ppgqaKG
ojLfkz4bfuu702Pffnw6WuNJ4I7+YwCE7d7z3he7YWAxr8qe1GtrEYU8NYMSH/CQP47i/R9IM0m9
xHDoPbyqdFtbDIW8Ob7ZwqX4nNpKvzeaB+es8ZhS1OWGgb4TEVEB4gvnSaPpHoNbzc6XGbIpSBya
OUs/pjLr3GLG1yJJb8EJPZZfTZzfTXIlTpVv09WxR6gFxjxIKlIz74WDffjC+6nHfkUV0DFNbXRq
JO/Vbof5M104ceLAXoP1L0D7O8s+NmUZSE4lDGcziMhq8KJRt1HfRCUKtNvbejD+j/aAeRMLM04I
geZBn0tzn0aRegndI9bxpB8Il2wKCYP85FQjHFHilEW8pheV2NO8ZhZPPa0L6dB+NQWIoo53hNLJ
QXNrgkDjsLEIWy6EANAOu5HpbgX4rfvO/JShnBtycxSZE7nMy4yMsyCPCCIWA4BS8sThWy8OXswC
sexJGpFDgb64smCFvWgxtFdF1wWlCYsgSGqnvvVZSXyRKrmBtCpdEn2mKWhW5MuzqyeZps7rtYnU
t6XfSNssDFJwW8a0iFeweK5yNd+GRjGxA17O/n2pmiTuEiSa0dEHbRhwSt5ylg/q8Kzda94HNsEU
4qBAMmGJ1JJwkUW6tbIa09C6TrQbi4XO8ea/X6tTEBxzC9i0cvJDivsyUL9YiReYbhefn5ylxaYi
ktbs7U3spOItjQsrOHDma4hjcMaloklpnyz/6tzjSB3R2yAXiqwsA6PAveUN+dFnits97jfie8Kx
KaS+8mrls3XVU6R2ykGSj0qihSSME4EEGlyzvXLrpBzunpR7AG2e0uJEaZI014JZoHLuFwMCjboR
PTz4UN8EKiLKLa7oGD/v9zFyF1FgWmC306Qqe/xhys7LwczNjFUvgsHCTSPcjaaOQOVSmR7lDmmi
Pq+oMOAuIu5x5NcG1fZv4GoGxuVyrKtwrLgFqVqRaM8a5b2oTapjeyrFLsmyXM4Z0Y/zmkz+p5cl
TE8nJfqhb3RYg6FhiIZNyOmRd94DpOyCEaWEHwg+k/sbCFzRPhvEtvaNbjW+HyTB6tdTBxzac0Fl
iJ/1uLdC+5BavgXscWxwq/A6FLBZ6Bnmi50eAnpIQ+8/GrwWikAfzJ5rJ8mHWFqB9RW0nI1J/c1d
8A+eP5oyp1TJcmvemzQO6gwlOOyHPNkLrxMpRQWPC1XLbsSJJh7J+u0kTey3++ydn4sSuhNwlbZk
IhHhRI1JgrXb/yjN9zaPYNzOj1VngHv7BjhwX1jXylXtrGZGV20uI3tUAIcLpyUU9YNxZxu9jteL
G0+KHeMrJ5JvxpsJLBI6jwxdtnOPMpKkKGYxwhQ1mgKHNgqxH4Mjr32cq2HSOywAO/7kXrtSnvqV
GWCthpGhwArJ5U94VdAm47GYGeg5sR3Utl2Q8aB3Xntjewn0d/Jg1z8I9Lkofc1IDZCSGh5E62Xh
LVh2gdgdEGGygAzw5eJ1d0MrGnQTfphfBb3gDMwf+hMGVM/t303h0PJy51CKbI9PzK1+BXYd8cuR
TJI5yj8FLKqvPlFRv5aNfq5DHC3rMGBu4rGO9dZ/Mj44UU1oD/6L9N11TogX2J1J8beUIt3vak3W
eTTlKafYqzf+nRhkEY/KRDV7aHOjZFjEQ8ImGtUrzG8t+13qRY2aCfwTVC8XE+UZhiv3Z5+x5P10
T84sK5BEcJU3midyobdaF0ZMNBBbJtMsl0uoGkangXAcPKdg4jFcJf8j3wucw7iTUq6x79ZruO4l
ycsAwbbR2Ic9uh8XnjJFxV0l3yJyxDUSjy3tSpermuCRpUWuZyZBGlkPRRVPL/bhWYwYg+xPIuGZ
Za9TSqD3eLxvLmatzad2nGzkKsWDgDhj7yHlgW9HLboBRgCtpckP/UCRmVvCUUgRVSHswpLnm1J1
avHTLhRdndaTt/W7CoE8XA0xZu0/8yKsTlZ3JMJeSjVy6cau4x694iIxs4OemK/3MprrnVOk0m2W
T7wFqFo/xyWZOL6IHZHwUI/ssjM9hx2Kg8rnMq6LpedQm6E/DQpG6DwkjhC+0W591Ij/zznuz8T3
rUyll5bT35RTBXS9PbZ+5w0UOMCNnvOdNScYknLF8eLcX8hSbwZq7V0ZzTOKX+UFAXsKNx9nYEmA
+s7WlrF8Pk8OjfuoYBm6kSgEjTsIW97Q7caW1BuSZ4KKn9uxE0s/oSTGO+G22nor1M3W/Wm2xBCx
MK0Xi+DVBXRgV9xGx1E06cRoIkfNrUx9VlCXZCcdpyDiSFdeFcCRK7ygrCU5muVib6BdzUPjnXjW
nayyo1jiCq0sElClL/XrXLKyOX6HbpQEoLkNtc7ars9XZcnbueaMRSy3y+F2rqQ0GXs5vKwuDRtD
lK6FW9pmmZ/H6A6DUdkpviahlbKdB1UoRX3A1EUiYjDCeIBRp4fuITWzh1sAPuk5XMu/2Ugr32vl
rNpoXC3gqjlxKkuRjgHa0h9v6HtM7xNBIWM8v9HV1s0qAeaUkp1eCwEpghILs7OgylOYghQuCzLx
fn8mS/uFYyklzU0PKCF5eWqRhklGqJ8zOU8ApvNjsnepYVLwUZQ0Za6y+NWz07cfEnYuyz4tPfwV
lumolouCxm+qSYCZ3dJzWmIG4XxjoW2h30r+QphQRhEq5HXlODY5opZ4IkVqlir+RYdNtxkQpcK6
nYoDl0i4aBn62Yj3jFz5gfmd7Vo1Qogg5YudN0mqq6U7tqyXCjLWPoIIWpxYrD5US9UUBVaBV+hT
uIUN9h3EJZZl1VZJe0ScyaWA9uJC08imesosrfxEez5EhAlUTpbrmoPkk6jVJEc6bzHLqggVrT0M
13++uiejxzidy9Qdwsh5KaQjz+5BgAji1aRFYuOecDEPmyd3WHy+hADN8xJ7k2ZdZOvfBq1u03II
P9O+QfIWec63kp7yTRXKYvQUbRB6eqaGlzsCdc9ta9qri12Kwps8yhM0WAqfdjs94IPCQsyyT3MS
xYJUfkeZT85LG1X05q9Y1QBWS31UkNn0gjFofAvB1zEybu6LFnCe7je/WdhZvhDgsf3jSyTg0HqI
vtAt8yM1uJ7LS33NqC0UOe67ebdKVOUNcTszKHsxnlayJgOSQbV9fCri01/5fdi2o9ZRceEUm9e9
ZvuOYKW5FOHzOfl3pXSprY6IFk8BXUfccZr8DyIbZQr7kwnesA3L4Q5rz1fOkfAMCytfKApHY+cG
QR5rS2J/Cr3M8wVb/m3hW5uwmENhtPEH0rV9zabTMq23KtcbXE3wfZVvx36cn5Ek2+ok0v6fRyk1
lomZryewIkkDZIqroD4jGQO8NL4KNEEOPVOHEsbwHLesLpIt/PaGuU+76zc35US4HzlvC8Q0SGyu
SGSWMnsdg56xhpSlhjl2c4LbY65wNivPClv+IhdQxmemFrt9M347wB5VsFS4g90vfD9GjxCdFVd9
T0xGWxmv/uW3qhPSl7tyq4Cd9riOuIakmCYniSsh3NnLxB9KbzROxZTPZngcE9VtVFc2EhQeM8u8
BMGDf9B5ugnfGQVwx+zx/YnCmSJ/56vJuXQbCe5v+vOa9XwsT0SMeJjlWcBSQmVxaF0xkd0Vo3Ci
zIx/1CQG80bfA4Vb2RicVyZ0Y3Hq133mFjG3RPmkcwHOS1fJUa85E9qdSdcwhf9gQYbqOdSLHrmw
pdnAn48Hhr8Cvh1o3bsuvtvPslJLlo3mUls2T3N1/BE7Cdp+naFGYD4kF28w20dE+W3ciQOpbUk+
T4UAJ/sEtW/gJjgPW8n3CAticNrh2MYlk/jAhfSRZXQwC1KmultA/FhoCAXMw8fONA88jSqQIlKf
zzaF1/sKFhK1v2NpjxkRqna8clmD1X+kkrOqNKws+PAQgEFvNbNiHa5iImVntqFO99dubbM2hdwN
7rtsty05Hw2ju4LMDVYmA932VdsWdgGKW2T7sYcUrkqRa3xIaE44yOSPhq+iy2frnTYvt5xK2Ops
2v64aJKntJAad0CRQk5LCplLjqtj79k7NeD8+eyGgGmpOYwiLPlVy0YFOnzlUIrhCWVRBwz3+FQO
opfP5u8TpeCBxbnFKConNVnpRcsZetwGgV5XCUJm0Qd4p7a1VGHUK+W/R7toiVlmwtmcuwuosIFn
f9UKz/KMmBT2HkcT/zgVfrL8N0BWFJfO+s2IilDN6MmMdTIWvXU98BJqUV5QwI8vxKdS1AM9OvVb
liT69nbTWlqiv2sVReYZLHZtHHjnGNF6kzg7zlatExYit7SZG7lZOXDJ9XZKTh8b1TlKZ/hcdF9x
bPRSyUdMUYcD4eQqUeDHVaryBQiAasabj1ha/DkGPVcf0xPDPThcEpWTM4t+5ZxLEoOuPngqLN3M
4+5vQKkFyNRVYVcXRoXhzHda9OI2RP7MQY5WqCEE49eeyJOtNPhNPXQTpVa5Xr/F8t7pZUuqgZI7
y6j8hWbMKWBv+I0K/2fr09w/KJvuWNfZpoAS1qAfVDL0LiR0bJRMcca7It5HSR4pUZrmov4CqRni
WDM3XopYpB5C2Ry9u0QoJGWcCfvm/8CkykwOnIEXHBCHavziQJdpHgHFTaKlUl1Qe/hTIV6sYfk8
IHYcZqGGCNjVUDCh7nQ1U3znbal19Yi92U+/ZZND/UIKe+F9PK2hIFr99DDxqGvkeZbAHX184CjI
8Ai0Fd62pXgSBTXO37OqwBXWOlNX5n0m5+2WKFiaiDYkefVZRL7hEvYC/kKOWAjbucQjZ436Ignz
Sro7YFj9Y58F7FU0Ue2Y9LyPBg5OlZJ5k3H+Xk1VWh8TJKmEQvwVMEIYKoQ/fdgvA6ib9j79DhCc
Q8Z7kS22xzp99YGrlII4ItFtwqLF4WWqMM9tV5ZNdmjSJRkDkVX7MiGGi3SgFwPHTDKMZ6lsGtjK
DWW5iWMpxp94Sks+DXbDuNlbbQ/hDPfVHyfHJU7Qm7gN/zMEjklHQ1BRVNxMfJUWD27IqUv+l72K
FyqvtKIFpYQEkjzHC2ce/H7uPmYREUOm2/bFqcePCp9Mfh4F4deSJg39LmWoGus3mzeZTQHZxo5+
Ax627T9u+oDXayr+CvUsFuCrCb5/8Mzc2QI1URN8FksweWKC64r5lbTV74cIdGKAxd3i/ZT+Gb2E
Lh14+XbcCHk8RKJRpadcDlXSRcW5+mCy9D86Fu9Vu3qLySuZeP+Oj3za/hWzAmaw/y5DL7rZM+vg
qr/8wRPZwLUJLzfoZFEcSt6BQWa06tb9s2zIW9ZVfC+TPfQY249s7DvuC8bpr8B1ZvEoVOcVsigI
iMRSz+UO+DYeF/C44Tf8WIpXj3qHLq7QF0hyCmLBx8CpXmZ8iE36FSiea1vE5qoZnZVOiZeg19eS
bMPLtUdXVJXLI3WFti0k180HgLqECtEQPrCeG+Zrkdvo1vTp/Ke18JMvDOg61zLUY607f/+M48TJ
bKr4sWoveCiKERua7tiXis1tFltUnmXwkoz4egL3GStUf6ampKtHToIVJ7HevsyhYB4JHpT+84S9
ZecIEH2E3OCDgQa0HfheF9K6VWXvtbPK30kG9eFThW4FexaC3XMUxp83dH5Ff2GA8NHpZZ/lcswc
THq7t8IajGsDTqmVdJlAHdNkMhAXH1brivqK8ed8EcukXtwnpaEDGEC2IIvhrZthnrzCTHXN7dT1
YmeSiDZmB5S+FjcCottIjlvYpN0eKMY5DLVDnIOliOGrp8eGQATYnFuLrv/5fX4B+bBttne8Fsx5
9i/SX8E1TkiN0PLh6hs0A3WXiHHKfPdbuq0qIouU8JxR/mjm1T6gqQcAYGOdE9iRQwF/IxwXGtH/
JmgWAizwl7IAf/UvnWg8z0DYXLPDXPzN1guzj+AFkLwG1sFvmbcp/bdTTuHfZgSSv1fgRjN8/ir8
wZz4pCFOBTSdI9zFI7yTtYScpuPLgZ/fJoH2/C2hMHeagVCIIIHDgUIMowQ89iRsnZibPXAXRHat
6Aexj7kaXBE980+UzsQIPSRhAyczirKGLhEScbzjNUytG3u+SdGI5RVp5fenUyqp8o40Jx4dj+JZ
LZ0manqF8MKFJyBoXvOUWHi2oOiYHzEhtShh+Ab6urzbWuDG21DGmnN00m7VcONG7b5iRiefSzdp
V5zhrVlEA6gRfuqCSLqZLTjPCFLyeYCVrz4+uMre9Ajf9EL+jc9kEOs0C8hMxyffCMIvP4cRKKtl
4oHsyugl3I46jmLvxA/ULvvGmL02NQmrGS62Rb7EulWihdpdvr7pb+ScOZBR5yQPswd6SoHBaGIi
+aMlBOisue14RgJ8xWdP6I7OIifAe7Zcxga06wPjwu0PQiN5hZBNe8V0hzGwAR28wUR/bmGTz40f
zTdlo5dMpmnAjyfFk4bGAItWB9ovGnPV580IYx3uDw6AHLACt2b+TH1BliCKaMevJqcClzZsR7EJ
bFPgCy8MyjEYE5DnU7wdVWHrAYOdAZz9c9l17LZQECLsznCnZOinLlDlafv7b6Auo6d+TGrlXNHa
Bsvkz1+1RR8H5cdZoKxLQja2Sx5puUcaTDoY/Mq8f9OOqtksurqfq8P0n/Ri1rGGJay9BIYBhiej
BLrvmc8cbAyJ0aKYFpr9d1WeVVETphpQhrlkdVn//JwEXkE/pFnlH6xaVMViVGZuSMPQfo0yf8vM
J4HcPjLgw/19aT2t7aiL7+7kPzy6n/Vr/pa0jzF/bZbZdWjUReBKfJNF3BfyaOiI/2/yh4/uX4vH
8Vjhopvov8Q12YEc3S00iBuxGauXlB0/XpwQ+miMRgRuInPpcnXNiYWUnNmNbP3Ezpqxn1p8wR3/
f7Cg5U75lI6d1O7sa6P+G66wWyPP8eBeuUBJTDMczxp4fQQWqrh9ePN8UNKuBsmPJgBmbO1LVmmH
syQBWizuMMoS2lRHGvKAl9CfD9sYc6nk/unIn2nQHnQi+5Go44+XJz5D3nnAMsAsGcSSKIFA7lBm
O1CACTCtuq8iZnKZ4O00SoOifAMcCMd77AvAirH5p5vA9t259PXEfeUMgPakO5cOq3aCEYErG9US
gnPxD4h84qN89WlSVTs8BB2fbfhvtWxNvjVYX1Arfut4h+qGKJ4jJSjxg13CR+P0J7FzYfs/wQYf
j/GmNC+OfToU1nR5Miei7nNXiY+3F8GdT22XkjjPI4KBgvCItXIPGk0F3Bco8kLFJYrhHkXmcmjH
hOiImaZG5ExJ5tKYoW/SeNM+Q16knXwb8RLashKRUVBAplaFyJUaJl8fp1XM7aof1pR+iCOpFAHU
ZSN911+3YSYeXrAy3C7to4l0Lfe113PoGJsI2pUSoBge0fddUO9dZQB0V2kqGtejWjHj/voj4hEU
EbpsxNUWjCGetQz+TSI0z778F8MF9ho0JlFdjy4i5fkSQZlc8QBkti7kXfQDQGRLreP1KrnqiT9A
GOkL+cLubsWSZRwWh0zZtPMNObbEh/fe4q+IaSGlWrxoFXAj7BxckWf8Qs2w3Krl0iMapfjnCF53
i5pozA/GdzORm8yROK724QzIYy2ovOp4zKeiuk8SUGAilx01h2jXlv0n8cDQ4EIKOyvdXoOIq/FX
mlazcKu8Rg+ZS7OjlWkuaMIgSrZGzgnjuvmDtW3u9k1nsZiL+urmrp8HtZQ9Eo5Kjhh4vB9AFcsf
KVtKZca2HwJqHft3XJjKP6rZe7E+O0iHPsv92iJC0mivjIrkJC30TmHW0LwVDSiZi11p8uAqBB+f
QlIGTNy5vtknwdlh1ze6Z1SapzPtRqQDlCIkp1YlDkqevenAzn6gfj1Cy85BOdd21YVL1pluGCgG
ZPPhOlpCMT1NbeDCGqnd14/ARPaZ24N/xePW7yLj54T4uL0SM1Q86t9DlKKcDR3tsmVelsl+luMu
Z4rBqc2XFXTeLV2KIcMfw/jTrXLBmYx7VFACd9z2nJAT25TAfNh9rJlYvNVO1xL3gdSpzQ6x1bgy
Wwu1h5h8c02RudUToInusQLhW65MOdAl8qxckMyOOr0plBFeoTRACK0bF9zYUaEmHbiXARfvQIWS
ReWDoY05DOmbb/1C2jV8pFUbOzNZRQqW3nlbEtBFNANtwZ/DnsqW1UcOkeClEshD3N1BAiurt3wG
hDYvmh5o4KoaZR0hZPThBR64PbGK+RXKSV6gPHck3KMl4xzoxoiGXFnM2qAxDwmjAOhTUjL59oou
pCneS6C7d2JJct2xjkM4XTxd4Or79y8JFOCi+JdzynALQBUUyiGy2LAhi6DG4HDoE5QMCHxGNPJl
FhGueV3YP/peZod4+ZiDDQ5RIZMSDqgVV6nF8xErfYE9ySscjn/lDccmOV1mjVnCwtVO2G6iMuwa
62IpuZYiKFPnSuCijC4bLPAzQaiLTBnOzHtEWBGJluSDV2JRvglrIg04lplNX1/ErfedusICl4pm
Y75HPhN9U0ZxL02HTQDsCc2lsDpCx2yZZiYmhLZx25gTFok0tx1jfnY0n8GQGYkuk5L7CdLQkrxV
5qqkzRQzZkASMPjJ031UMi7FQGkun12MLdlJ24YNfehRuAfCZyvbkQxPbl/QXBQdhamJORc1+BPr
ynYFFMplBj1QFOqRwIzlMg2OCcp4GbL35L1LazQtOOVOBBG6rWY7FfJFNfycLxXE0ByxZ0+nyPmR
moaSD/nCKPVCIv02deZdhX++nZlq+clmKHrox+gDcF4vEYw0uzcif8xy2xNDHwipwzTxukpHLkSH
Mmi28CLNneUH3ir18ljZwBrhyy6j2I3KU5ZJ/FgtKYS6R/kZGmd83AAVBOjGcC/wvRAOMgEYiAHI
i/Ap+KQnM9GIY6qJi7mxMk6F1xYvs17joJv5gJwiNNivoAj/OJG/GgTtcxUlNCLpxcY9EwmQ8ExX
saLjSCBI2juOXynt4PANPP+lqkPaMYPJwEQU5KsCVLHP+tqMbCwErkgXFRDgISDCx7niO/CUwxSA
8SRBBaXJjigSz+eV8OBwpHdyhQverGI2JOdmcNvd7siE83ofBPo8rfsLc+1SlxDjgSreiqoYn7Jz
4S5UcSByeOUF9rge0De4qyTcbAsoJ0P2TLjddd480IwS2ZJ0Qd7To9WLWvAcp8+a3/ULt06Aj7vL
ONKRQ6tCIaMbZ9vtRg1Jse1+F12ZEEPgAorVzJDq2h1haCR5T/yUK19oIK3owMRSRb8Cm8U0W3DO
EE4cluICottkKRvBO5BRTrC8v+6iPpLFUpB43wq9clZlPxLOVbP9G7f2y28IwN40tCSzafqNISEU
wOkb/gN8FlJYz3CXGbsM9p5EXFNfQ1PIuB1qiVzSVfbOwwKBAUDKx0jCDwUcyGSqrjdEQ3pm8GX6
HxJRmn84vFEhqqK10VSGZo1b0smZLNKYXrrImtq94lohJXjTxDI2GWo8rjoHQPR8guVHMXDGXOy+
odrerxrAhhzKDXnDDgzkRGhdAyJbVyJTBd8kPJR3qltViftZ4p7VOMSVID5n6nLHDLfCgBPqnQpI
EHOTYj6g5hDNE2v/+RwsOh6xRvQiR8cYg2L5omD0EFzgBSc9X/nOVr5WAGZQHRoKDi1bOCcGEUyG
llTcdWXGP/OgguVMZLh2tNMfCTXTPwTKCSmuhSuh+ztKXHrtM1YPFNdlFYJMKhNUY/t9UGK1cZAt
4M7wkl2fdLLMMLJS/8QExL7KhlnCs1Et/1WjjXayaAvmxGndMFkdORineKfrcGKelQkhUsioJUSA
iZIaliedseCt1uvGWGgGv37p6Quuk9GK06bZ6GBSw9hp3tJ7f/9CdzN/OIJGwF9hjfhI3uZFh7HS
vUwOYVCwFL6x50wRBnYMkZTN1eYP53qWYRdloAS0eCW9uJT/RMsQC6qI03uMaFDsLczKJvhZLa7U
GraiAQWq/Bhk+BT83BYltzVIrkeKgtoJ5qlEwPnMCjNjIOrOrYptzib9IwsrDsRCG5tNu5XzqHR0
UHC/mieqdsRjWAF/FylvG7h5OP9WxCpIvFadQmXOxT4IFrm329pF1+h9PC2iizLNHMCILf00VT2/
oyDq6Vs1aA1Z7TzvU/Rpsf1Yh5hp+n6r/Vyqy0eYsSWJQ5NDgKbuIn/kaRFec+FZ9a7SIK1Zow69
deSFoZGZS7ONqiS596A5dwEj8iI0NcHwLDGp1pDW11Ty54fvzxC5faUcUMxQmI8u54NSsn0C217x
mJNQIsHuYCUYc6A+BihFEYZhdRa772mEFZ7oESv18Bwg3pMyt7+FTb4DrjXLTzDje+RIZMeoPNff
Di/osJxWgAQfHoldz3iisZCnhn1BhSpRrPzc9Y84tLftPp65QrQS8XzH98YaixtKcWmVqj2Am8av
R5feS9kq1dRV1b/whEvTNrG7s9MGY6SDABhtW7ZG6vFhZV6enS51QRXQb1wemb9MJ+ikDtxog+IP
Vujl8JfbjswTLxv8clW3hLMvnb/Nv6KK6Rii9RXEVnlmAG70fcN1X/0vouQjEgw9vLF4TamLBxCe
++nxlaP79EsHDyYr95V8V3eUBFWSrry3/Dq1i+wRzO8BkI6npJGI3uF8vfAS3lHJCEXaFyF+eiIP
VW8kiBGq10/m6a+W2/4v/zbEspXxGO7GIlZN0yhzDUud5+u6IaZAQ/PoX3XsBYxX6dKmrSkM0Mt1
2wMQ0GZ1SXKYqsUdTivDMNCY+N8/XRS9JuEw0PcpWqrllEsZNsbFRyvrEsafe1bt+xaLDTMU1Ajx
ahO5qVOUTFkOT70xkl3YeVm+pbfBzujxON8CZ51x9BK1FgVTXoLorULGsgL6b7MxbVmnYlg1AwAz
FpJ5+54bHK2KBnv7bARtegTZFeblh1djBzzXy9Yb24Whctxyku4FR31zpJBN0wED4BheunBph5Xo
ebZEGC37Tw9RCSlOg3Nk4wZ8WJUvMBoQQtHWCQ3pmmChWmICh81GWtWCf/so5y91biQlPpT1fVqW
wzQq+pg1CJU07Bux3eployN7MMya4gwPe2m6Z7cEinJt5j/j1YNcAulVUjoXQYCtpfOlTcFD4oOM
Rx4pvBS890OX8ON6YvUiQyOI+JgH1SZwKzQUGXJBlVNNN0b1lgA32U9rOQIOJMjecBGTWSKUYwcC
OMt2p8DrthFqzADoBu14jadQ48+/7ggX25BBnLmiEFIuNxmFJ/Oyg/GjMaZq/AAJjxeGEU7FIaqy
5NZNBQzIvpnXedi5rdAS+4yPw4IKZqSt7ibvERchPxq6mQtv+8vQBYbDH3BPXIOjyJa1Imw72kr0
sUKAql9vOC8kEJYjRt2EnX7CGUwypfsFWOcXtyJcSTdNHcuwh+M4K9krON9oRks+eyE+egEGlSFD
XHmlpChMBOHv7k8LyrzwabwdVGFNJjUryctnmuBurgNGjaWlZ9TCNpyx5uFPd4MiXLZjH9ysLTsV
Rqi/1LvrH0oyj0wW3whH3GK1rhqA03uF4CrELTx4AiA+JhaL0xvf3yQTw5QQ6Jx6470cvmhCf9cv
UOlUxsAsvKuBCLWl2WMdjW3aExMxZITbzLjb7dJ28fNZUm1k2xV6OSGOLOjCWu4/eOTjbaN8hwYf
2Qhk335ovMkHy+wLGMAOr3ABWV6POHcpRGEwrsUaw5BehBvCSk+TpFwn2zlO9x+URC2k9QpF+L2i
Cm2hyy84LHPQuseP7wN7u048+C2vR+1/oQdljhzNPKPPm+FzQX1YEmaZfq3jHy/kUMIS7MzEDFPC
ABApbAfQ9j1Skxz8c0ZZKT+H0O0u13oTe1EhBNA1cx0J+oMhYq7C4kBDwxrQyZxo83zCtIfumJoY
hGG6XDBzlvHULYUzVsHsDXAbQVXrlNH1INaNpn4Qm3cwmP6wGPeW6g72yeX1B/E8lu0muaKx3uUW
9V/rGSvOX4jMnel8hBOOeUXo5Xkl3HtdbjUZehMxO7KJOAtY7CmY81nigaYkVCngQ3fCqckI7vRj
sE8RS2Je9EX+xVYWcppnZJ0WYHb5crxy+/bYxxR4JBvhVAK9qI3zHSQYc9GjZ7HzRiIecW1oCPoo
XlIoRgOTeuYwUbHSy8W2cppzlwDGR0joqQC7tYG3TXf7Qqep1btviXySVxlivhlabaMmFWsp+Q4p
nARBIZOTbtqyGlwvoMiJfrScO46Pb3CFeGz+kx+T3xefjzaCOG7wSQiHlqY6qxu70Xn0HIKgzm0U
iwou53WBWnzSFKiExd26PlQh0SexUraS78yHZWZKhg2N3S+0SKxlsVsb2GjZE98p6lcN7v9pAKN2
XCpGjkwciGDpLwVaQ2MknYyRu38ejbBWFSpPSHxTN5FEB68qfnifik2pi3U9LIksIysdt/p16Qu9
XWhbH2ZyWxr+tThRRX/lIcrZIBlRVqf9YwX5nqomFJ0I10oiyUjwzOSlJs2Y8mVREzNee130tOIc
LizP24Jpcu73OafqE7dBxzqBrLob1hK13kEzG+p4LHhce5qiaQ3SuT70J69+1+FYO8INsEUvvx8q
IcmDGAf9D9yaPtfLqhh5H+0mpgn0wBZFQCvD5ZT6+ulMlCfGeSypXjf+l7BozQ63QyIWYLYgNU8o
cFuHqiiwjxZe23zocyZpIbyOJCFsMMg6OOl0Le9HonG4iviq7a9mDHFj8bz6SzGeSThYhGpKKeMl
1a4yRCvyicZ8I5jPON2cZve2NVgqYq3FXmM1j9eot61SPHc9SATx8k/IYD3E2rWe5TETNIQyQLzf
k/X0/tGQOB35Dd34mn7+4ZYkxFPFOtW+2COLwQZ12nmJtC7hNLF1y2fmmWSFQZfEfAC8/KJQFTtd
UGFyXTTVZtz++BB8/mo8zgTzR0DLzJca0PeSHSqmO4JKZc4LA9VRLGZF0aeMiKlmmisA532DpnqU
KUI+sHTZHIAQNhxjgbHh66EFYGHNz/BIftCQQ4NneuMSBWVNQXNqadK+qxRXT2zfkvOfW1qo47CN
tXFmIAPqpnyatS0kU3gLXsChqm3CvlZ+AqtpqxrhHhQ+k/YaJyevY8CN6nU/h2u3atdwqnM2mZQf
pUDe+FvdzbxFuJoRlRjJdXWzbPVSFH6hwjIxTkxdCoxX5UdmVq/RnNMIFNagZCvffJ9N4wKM5qNa
opmfGKC2T+CexbSAkD5C2BpWcJ56eKYvlr0dCZZ2lcJiVGI5DULyvQ+VjAYJZyRrjDTHn0MvOW8P
9Kmk21odJrQC50d2fjlgd+z3apEF9TiIAsOYhdfYiKkAaEh6nHWwly7OhXOeoPWbgBOpzQcxK+BU
jV08ffRVURcgDR443AuLXHVAjpRXzS9NHse/ojE70t1kC1kV7nRiKCYSJE5lVr95FUkpl7GmtZ8y
9o7vKEq6nUFFAJXBwPsHrmtM3xiXqpdbQOxcj3B3ox7MX3mRMwE0df1ybe8SG/XEmaXS/OoeVUKU
hXmZcXNbhm7cihXzLX1ofON+vfiJN+uh5v/3zLwxtw7AZ+4QY+goGW+/4lIbRmWhw+Ahejk1W7E1
FWtStLoEZ0np5SpP74xFJjhAsD42697QbwQU4QuaYGlGfJIG3oFM0JX4xJqqrNu7fC3EvCf4tKTI
LF+XTo+bJbu6YcNPxZKEQtmnZFnljFPgT3TIqUaw10T1oE6V4Ol5J+Vr2y6HamKI5YPuD0kjVHiD
0nMEoVCTArFdnKT/tmnj+6yeBPz51c8ydC+xsFymrj93xq1UxsPzDrdYK7cMwr9v6GT4L+/mZRaq
9TqBziOisoR0TIzc5eESqTdP9yGh2lbIQ1PqnFrkVvAgF2QHjM1wSCSmdQGiNO0EV7L1Cjeziu+C
8BubTGmzqz2oL8Sz20EL9FdVR7PX28lo9pInodZy8J2lRv9H6xDx8igFvJ8qhIxmN4ZP6Zrgczly
mf5MTWgNsHB3EtMcUR+NV6Oya4oIQHHDvdL3haKoezw/rv4O6ilZpAZP/3Vwh7Mt6fxp0g1QUrw9
PVc3VvTAwH0qZJVqTeIMQ+hssPhAZLNlujbBDScFK5BcRQhn0IthvMi4wblXW60p9F+XmBuVE3LC
TrYOXMX0RIn2+15SQdWFcOKVMBsV795g4BXBjom3nh2vQC7fzDb0pJ+OgCXkGyIxBPWTvAyNxMh8
/X6U73Ltk/6gxGjFGO5Pcn/PI1rRzOEWh6rB1IjYWEIm5AH+B/zMxnfLNEVwLUEseJDu2guN1ZAA
WX6Mg9xZvanKZCyhBg6LYwwktTUMVvROcuVzOvxdsgAFehWQoiztvkD74XOBMfe/fgilVCc/yh5x
ugUGx1ADbKdL/Hfud7CzQ/JT8L6RADwDlltgpFO1omgEl9BbgWkOLYjZWwFlyYHRJPZZutwExra3
K+w0uk0z1Qx6IsB5BNUHJdMbeG5ifgEGGDID1zVcs/OkTpUfCyE2zGk5kjlKOUb306Ob+SGCfIbT
Nx1lZVLzovK2DS6XfCmzuVn63/zc5kac+MEEVlTVt5dahnFabQD7qFb7vjNv4vHBM9bM0HKvm6n1
hO78gj4zenJdx99hzMPj0bJz2Ld7keWWAqtjwX//pnpdTvjLe5nb0RZfQFcY79gtrkNc0YkBiTCY
xfRy+Z7GMxSTTzR795G2p9V0yQKCE6YlKLcPlPmThHfKhGBfbPfLCI7v+J0vXxpJKIfVaAYXT7Fu
i2AHpxsS4Hdr45hvY3h/qCpDaZt4TObFHdDFFQXZ5aH5OyomrFsMacn3N8yx5CLQAsMQibMOLaZL
XfpZpN5sg8RB09oOaHFSsHoULLu3WxW49cfRKyqmqCosI9cYr43BQpOEV5T3dXCibVFcjgQPtrBA
g/dqk02qYEMpXfMljSwS0zTJup9vfEWmixE36Dqv39kbUAtijiHlFlifwf8mDM23cVEIopUaRat6
w+xUpkdp9P7GaUVV3nQRF24c3YCxHmt5Hv/M/RU0bNJOur9VOXe3eT3LZAJGbbxGL4ZFHgQBI0LO
j4ksXDg6aB5yp4madRikxNTeqzuKpRzA6uw+2so6MLpN7PL6LxUJtU/7anO6DLD8UF3W1zFbo67g
G60TndIhHJMgvZo2vh9FZT8xiIXqtEKiMiQBid/XkGT1RxT/Wf7pzsX9NF99EpTO88BxCdwvPgqG
7FPMhXD7B+mCSCOivpw5OZ/0/LAyal5XQStwHJ6npWmpD1+WRyLbIm296uSbVsp1kY8jPKyqudDR
xyV1V19UgWsBkBDjN4Uld8nUk/+gDOax3ccDsjllZC1dmctqPP1dtYPX6IegVaBGWzvrTrF/Zpa0
AWwIiN/LGpzEtIOk5mXlOQ9/uq77vjLQuCFuXjHXQcdY4aCZ2mIsHBCiHLBwOrfZP2flqpbr9tyI
4GseCFpslFYhMbcMCT9iz+NI7oZgXdgMTdO6RZ8kO3X6jowvTtsSuMBt6BeluL34d9167VniNLkD
3Xpp+L93o3hyTIWkJyfdsmUgYYt9YDuYu00253jm4v78mR0a7emgaLxgCsEYDJpGHZ9B2L+jo/4G
NwB/49CmOnGql8j91Ll6dwGAYw1g/mvNyk7XYaQs0IKr/I4sI/L7mLqb+sLV56EBjtvxDa2k0ZKG
NAK9RwBT+0zPDnCpcHGKKmByo6mfUoet7qhl4UM7Mong+Cf6MFr+zfSq+6qC5gY4sfsXdmDTABw7
OkhOAaDK2iU1vKotpBwlq0q6uYvsn54s1SjWyRGz02slu6LJFlJkvwMO90OQ5Xiqw+aNUdmxkAXj
pi+UPo2kbHI/q51fe0G996nPxT4s34+XGEtBbanu8Kokhd8mWOKavZnt6o/clEeVe6a8AeUOh5Wt
VbqCkQWinaTi7ESyri1r/SDp1cWnwX52tFQcVj1s0DF8QOf188sX1nb1vDC4YWQhyqFxeQ5eOPxS
x3amCrZ5JJ2OlMOPqyf4ngXTx351tBSbRyVuJUclfxn3YiB3iqtSNclvFva78OlZJCwYaP6xWqM4
nqUxGCL89Pmc3Dgq/qhqdrHTE4W5/YzpZRqE8G8CAzRV2uI3ir7qvFr2KuGv+mtaYMnYkAXVBwzZ
mx9Ksl4DdaDWbealj1RZWKi9z0ObCUnRymBPbFbRO5gP4LHzsOlijpEsBWF5sBD6EHKwfhrgH7Ru
YPcCZn15rBJ1gaSt/SbItJA6uP3gHz5YzSmMbpL9lPEbVHLiSTbwXI2S335NlsLfofBdyrneObKg
RT/n/kuEc9eoJsUalLPyr9KP4k8aY1+8ACYARWPkxgCIqOgUC0yF/FrZ63RYTfeH3bwPRtZnf46M
efkdACEvS1EsdAImVwRrKa8vw0mpkEEed1I47sQts7j1YJWHhg4muJ0aXaibF9CJf4UAmMhBIfJn
aRamg2TLZzmOCycpE2jro6VHDGaTZBMfy6rStpEd3rTzHd8ypqamDlNyTldPgYw6xwCAn21FaKeT
OFE7ylRz7Fqbr79HiCCzAm5O7HBZjMEeRKVZXjdUblaLLxE1nxIU8YUxpCXTkYXXezgyNlDTpI5D
KG9HkXnA0TPWEOaW1VaZPgMieiTd6lTl84TEKFlcP8rq63EjOiHqGCoEyaiTqLOIDFubzBzBnLLW
YKw7hWBcHTEaLzOmtkNdDstk43/IU8tqCnzN2FqneVKPj1Mb+VeDc4FaFXiYchUaGvjNE0EQVOmD
IaqTL8gnAO4ZdSQAFjCaWZrUF3A4oPctHOF/jbwBr3BKXhNSXbxz9430zIwmmxJiszvBFCJj7bDz
L77FOd25gZ/jPg1wFuqbVUIChROIO8aOaQkpkUDNB49/wiM7JhuavMA+s1zzb9NPxKxUh3J+QWyG
Ozyf0q3T1te3Jr2CSUa5hCr+nHHCtOW6jRbQZGlu3faKPXyr8OBsaA2Tf3cXdUT2MecsYhFznqyM
73HSnHFt0+dwlFFYELrH8ni83vMz2DIdPSXxyoN65nRc0mj0+qBded8V90dAgi/8Qr53GGy8JeSJ
EZhJ+SKfER6qibAKKyuNwDh3wm0tGWJwOqkzb8fVMcjxq+GdnEebOztYpbRVa6I9UuxqhJxSmU3q
olKWfnAA+PEOYgwpabYGPDqkljSoviIrHVbi0qOZeY2JMb+m7yBrbViP9xwdYMyiyiCL7+Jb7OvX
wgIA4vewufVEWw1Jn7EmKQB9hSER0Qhbqw4Bh8UhcLCmW851+q6COYJR+F1+CqcQ6z4Qq4NjieHK
lwUJ6D68FYt/TktCPknt7R0BMll6IS7avmsQQ/GmHiwQ/e8nDFN0PajG2nAL6Iv2Bgyjs/YyJUXv
zK1iHSFV3cxtY5sF6YMjl8UuJqgji6QjivhCbCBCF2rPj9Fuqx75aZ/g243xh37lSc5xU5mvOHyp
RnlPTzRmIHgX2UEX/PfRuIKoKuFY7VbQfDkrNJYurs7/6fD0pUoIwuZxCUbQWb0G/itxc3MfttuW
2evJ7GwXp7AgMfDxIllHLDVceQr+iE0bpBxO+JwYPeUN6CZh7jyPrxXKsaTt4A5YmRI6lZdMhzGj
RPLeEVV7WuYEAjZFq7E7PFKpPE6SaR7P8KXYyT9AmXeArEEQxWsmU7IN/GboQ1r8jDJRpo72mWjY
Qxj3o6R0jXCqeI+P+7vUFflLbJEOveme5D3ML2S+c2efUI7EagATaa2PHrE6wHb99JNuaMllveuF
GmqnCMHtg+He1gspYZqwcFnLb7xuEiQyN2H0SQ41n+7XGAAH8nFIQfJD+ozYmy4y6zeMFCuspRN2
+Mxnh78a207yVGYUqtnCKUiLOLrC8A5R54N684Pp0WeuyMkpdB5jfzpeLSuslx4WNchKgQ2wI7Dl
Yrv9tmcW37ncfcHAB3W47P6sUc4yyTA+iPC+j/+wLNixOehuO3suNFa820RH6s4wzFvcYfynIBOB
xWqga5RphdNaO4Ns//Wihr/W2d/XxcPR9UNKcDwnxGHiDKLZfjyWo+etWbA2MQWFGJjqgqY8lu82
VI7d5JFlHqS+KXihVlHMN1WuIvLTr82AfaK98KA5VZhPPJ2ZjxaJgCApHvSAXCeBTwrxaGUk1IyA
oovXSGNIjkvgybRxR+7jc1cqpCnCxLByxrU4U9wQnkIWtbxSVo5cU/G/sLLBdwpmexrgHzoXfsq2
VGVC3Agc1o7S6n7YTkG8d063smrNJNCnmdzTQJvY/BtdW3W5eYNnKjWK7ApMbS2df3C9L3g/Ynmd
gFn44DeTnsxDQW9TWiGDtTOgVzFj+XgwhZvr+DD54a3oBaEQRDxMFIwJznYKn1q923qE9mfzURbJ
mRStvf81wqc7JaX5o1yIsipMwTyEsAAqR0WWp+UgeYOLbplnfQ2muhVz2FPDN0noGO//9mzSNy7R
G0wv8/DhvTgy7gomuih2xPB0+adbu++qEZzhFeWGR+MHF6y1s5RHfiFA8eNiU4ppDR5QY7vxi0sL
VLnxWMrGCKsoS88cD+GVZv3lU34prnWzF3n1+TWASXLk5i8KhlM95/QSYCAzNP6uGSWeOnCudGBF
X99KrdW5rzADtpWsC28Vh06pm4ui0RuKtiyj1AqCXTqZ4tM9CoEGk76TH/p0mcXAa541RdlADoUf
K6vDg0KOGgadIIEte0pUhDuoroSag9T9xdkhUVZn9aIncHGA+9DeR6NiGlEjVbJB6+JxtsOlSQwi
Xhh++6OwzRTdVNb0tb3TLgPC5WrdSxukzAJkOxYWok+U7XaIdzOPr/kiNT+DuzBocsQmKZlIFppi
k4LYxUmvEWwprvYR7E4CF8aQej/Z2oF0u9U/PJpEHUnhglnigdWHS4W2uHwijEdgdEHnouynKXTg
QpJCpjBKeclqcgkbKLTemXAtQe3GsoDy2GRXJow/eVPJlodJHg1Y/gdDJhd+Qx0gZ+Y+e3aILd03
FuwZ9slo56Z/pu1SEA8IlFV2G3YXalT66V4mxRseJFdLF2CK2qTQTr/l/ermcDPOUmrCpf99sjXS
r9CvyLRg5wC7GGsCAhC1cJ3CZyi758LMr6Tb7w6xgK9ynh7FJQxZDd9HrYz3wOx6Xo/+xCTpFfV+
1GUM1fegndaX1AqANSnZRg+XVNo79VzTlp/Jfh0tDew4M1AYFuXFrCh32wQYpn6A+QRL2B5ZWohw
KAimQ6YgjY7HtUR20fjySqniP0sDbtqOsPoQhuqwSK/5poDOe3ZIcZK4kT9cnDQ6l2gRbSmSjvux
oSsVVu23G43UKXEPm2MhXrdaFem5ha8GQLXs1pZbCyImB7wjYoZAvo4yVR9WBSO7P82SBDkfryJ1
u0bI5L8kHR3s5B1wPbChfKtJHopjE1uW+Y2f4Xr7afXGyk5KkHxLv0pCrl/C8mG5p9708AzbmOkc
smx7RqE9spzqzt3pDwLMrigJf0oSrAtTyGGW40vCh/dGEDrO/PlnbWNSE3wwjf+wXq2MBc1H7wzG
tKuzHZHqfWHFQ2Islw4IzH4WRI7njcjTTE3dpD02ZD7N5YRub5T7oBC0SBTK+bG0Bm2qRRcTl1Wn
IybRfbKbKsp5AZ+T/snqKAkSNnV1FKTXTXlIT+be/B168OVwUzHSXCiOjJNca28anzMnrptqPdt0
N/MLQvrZz7wyHGGluIzBfYAMCvyxIuiVD4lHxH4hGNSnP1+BfU70urWXC6UQFL4JR/UQKWTyxZHN
t40D5XdEJlzo6YkCKEBHmb7bB6K1A7BP3cRREn8sKGrhSG5goEJJFNtB8RAzzS5VVfEXFf1XeXj0
ChT8u4Sd7WQbm41EFHTvUa5up8aa5jPCyU+4GJSmppuh4HDNFHBTphGDiJ25jZKqa7jWO6DrGCwj
Aw3+iRjmPEijxq/iXFCfU2XgFwwvyPa0FUCOJ4PIA4602BdtC6iaJ50sPx9jRzau+hE3XMOvF4EA
HSb1qa1cBroDlGbEClw83IlVaG+Jdr9adUPQgW1fY1jC96TzxvVu/XvTVeP9/FnRD4uh187y6m5S
QbiYSMaVr505Opu/CnDhVdzQ6QSg0nbdCgGaE5xA+u6CH2/Ba7VRjeQEXDWNjEv7i+zbhIzXIlbU
8i50JteUyaGUB+6T8bIhjSUcySV7MZ0gC+cfkFI7tQpfnAICooHahQ4v/rL54N/bGTOzlMywywD4
FTp0fb4+pPn2GZBckz1RPu1WCSonk5EfXbWD4Bp7YNcDb6SnjGEnlARtAHKLXCC8CCR/DWr3sjhC
rp/Jlx4sU00qSb0bz1/VAAuq+njpysRc7eeTMbDacju8gCEogfsf63cVOGdarNlrDCAFJMm5ZTR5
UUCpY4Pr58sF5ngNNSiZDGHHRO4Hqa7w8DEevr6mbw/48aVBJllYU+tq7u5YIbqRJzm2H5iWkOrk
Tqn+nnyT5ee7Tms/UIXxm/Kbsi+2GWjtKGRdYjzeowK810s2iAsk79oQ2EOlcmsThSE5wzBQeQCt
Z++xogpxDG6JPvqkj8VHy+EaZ/8DvXUVI8BVWJeMkv7qpWT+bXznDvq32Ej12BMrw8hJ8WUsP/Rw
pZIhelOko413PMfrzp43bnIqZaGN4hdA4VlmzpH6aghIrha4fcRaxli9rmmj72Spq+2gPEUrQnEP
jZ/67ZQnxXioCdbbCffxpJwqKLfWklcPshH/INAtIJ61SJUPmlvqkay8zh/TB11eUQJA40BYSLZT
m6NhL6IsSvjux1LPRcXvrlCkVJyRloPUiL9/nFbVkFg4JCGoBdVchi2n2TVoyYbVGel/FeKuZo/t
rFfVMIMrGwadNdc6deXXXWSTJiQJKew7Yht49WbOFnLoRd93aKGarMxtdoNh6CbFCbFU2QOiseXl
lD+ftg3mZkQV7bP0dJ4E5yxMqekT2tEBAmvY9gV0qPnr2vRl+ScCrLZ/mKJ8NolNsz8hpq+Sumt5
GkY4P5IiU+gmDszM4PBXzS1idamMcETVD891IdGV7QRhWXarUE6k4TpqzmRiXqf5zh0E+DCUhGuM
vZRxuCKfrLkvdst3eJ8rtrUQxkO0OlKNdBCMQys5r0eM3YFy0Sfy2wiCYQer/9UwwHqloHYkmC4p
Wqr6LoMjsyTACYHbEt893YMH9TfhcFp+X6IyOWyr8svrj4vBv4D+yGdheu5ga0BeLQWfOdgR7HEy
w/m9xjGIFAQRDNWJnjlGPv/CVeUgCJZwspbPPKLD3pZcq/TMGd3xxioaLNKZVMtez2nf4AXO3z2o
iEdIVMEASBkpuk03wjtrS+7bpwTlHE+FgkXNjnF5rLNGD0zrFBl6gKcRyADUXRXIwAcBcTQOLtI0
jHs3yabSIs9TtpTlbjtibajTWHMoDYhhqrhn3Xng4CSWkLcH26hWSSx7PJKa8uIJnrhDfu9sCaVI
RxSAEM+eFKiPYtHe3u/+W78t5P4UzWH530NTNH8hoMjVSLdCgdXPQybKRmMMlFKogJczgJaEirDX
v2LX92SGmCaf0QqpuFatOPlXQwQq2UppbPCsyL70kPL2D2ej12282ZOfQKFlQOb0/JVYq/SpAtFW
ksXYBfPa/L9ZA9nUtFXdaOcugRovXkrtxclPmOtofpgI/y8+CYJwt47hF5Z5/6gpUK6P9juOHClK
5Z5c4L3S73yqWSWCTV/r0T+byfW1wvTvF3D4csRp+E5vYIN4QSn7Wt5Hu7tDbWr562Kr5AysYbec
n8gwop6TwT4LUOo9O7KV5S1GO5NU47OShPDMHk/vw3BQXCf7TPF526K/jgC0JlYfMFYvZTHFSsjE
FGM1bFhCqTEx9YYVnXo1sKsUpJ/zRvXXXFQJz2IOEoYvdPDYq/DK3SI+5W+z7U8fF1axZDRyEzah
Gk/0wxoo0VrSED4WvvDuF8jem57G5JMU/arvClXtYuma3nXwg+K5flHG6pT20iUCyWD+o+6FiUHi
wILOj5R7PGz7aEQbL5rVsCSk87Vwsg6pA7CWSa7h7gXCRPNzPps9Ofif+UT1+mZgCg4RztUIzbW1
FPq1tJwVjnILjcc5YHgmxdbTC8/YJOwF/SsOHY3DRqSVCV4UOPhnbK4fTWH9uovuHww/iDn1fJCh
JT+kLrTQ0qV5cNstFP/6tSFG5JLkC5Vzh0kvxpsiHg2j0Z8oRNbiRNrDORJmg+Xr70985kp/XED2
PX+FWWC4e6WGdGChC5qvrT3k9BF6LyDBd0yXAMqSl0py6ed05oX8eDtoGbN8UwmhGRPC+0DOkPod
Hin6TMDHnGDeMuExw3FCwTtxYBAqcP5vhvKlHr8CXxHL7aeg12Y8WrxpGE1JwoyZHaQIzI7iS3Fs
Dbz0ZcsxoalFhYkTvgurYD3aMFmC78sseL0dzaU57zum51/cJfZE2SC/Yi1d03gvbQthQYsof4ee
eycci/NouUedMY9vp1Li0+STczVu5SSnfQ4gb/W3rUoGlpsxxWEmMmZE3Gy/KEZ13hDS/AXnIh6F
S2CrB3W43LNPQzhnHih1Cp07tIT39V+9DIOKQSXGhTHn6dRhKUvNDesyfiYfKgIAjb8SFReadakb
4F790hluFTDXDtOoTgeihNaoH+vZe14+eaIX6TTMp3rAyWVfa/Ie6Dhc3owsRV4WEsNuJKXm7KVs
JErYAgqhHQEaqnein9oM3ROoAURF3J3jlyfrFhBx3OP5pjLLNKsbhiyXip/yWRpUcN8dDzB/Qks0
/1e2i/iKfsKMzeUQPg4XSFZCHmYr6mVjIGdyJioKbNJGlqYV+DPYA9IGaqYO+/2QHDHSv+xo+MnQ
jfwy+6XdXanxyOLt8l7BUF07Nr9vQCHu+ejK1kCdY1y2kxJShNwP5bFoMqKtnHOJOIzJfh7E3adR
/ceG7WTam8GMdp62CuYJ3ubr/Z/0+l0k+EHHuR1CT+DW9er1rCU1nOtGD9J1TCgpRkbTHb0Ng155
htxKJvBvf4LPWvZvkHG1tgBRJeU7DECRFkyyDzQBEI4wRujf64Fmbu5Nwf4imSWTZFXiGxqr+4vh
1w2klRyUmwSAoVrkIw6m27lzLydksjzDW+FrLxLvN3p5FzjU/+yFMgbrsyz8Gb2D/+7Q3W/ztK1J
uE2MGecp+WQxVP6e4E3ysyCqGHoAcfriBsl3pf7b/U6iUHNnMCyu17GRIT/vYwxpfBRjZ7M1XdkC
3ZMbVPsNdyecVA/xMNBZh7rUjuSqAndaIJ6gUuKL5HDiSVfoF8BVOhj2bS2cuJ+lyeTTVJpappj4
EMXoIuEfx0mT2rk9BQEEUZVj/X4q2rIUz/yQbXjx9GMJs9qw7N6LYhycOY7zZyNb2suM3PM4g0Er
zD3GqqE9ZPbNrhKgjvGUdTXEoKN2moRQ++9jSckboxD981p27AY8FRQ/uDNXLT1asRXzvddIa1ZH
jtUHB10Jd/LT6JDR0rj1G52yZfzI//6NUrSL9HRPWn9wlvc6C2CTQjAT0ZgM3f2Vxv3VKzN1ONWL
gOZxL5rQPPyXrccZHDjBBfs753B5EqYQRRWkDuVxPoZSPJOcqe5SOUj87081jQ0R4KWhJd5PstNM
MGbZ3fpmPsJ5Cs4nAgpCZPoeTfzXshCdQrhOWuyZHw7X6N4fUmOk1Gl1UOLaw/ZMpBTg0bA+vxb5
U+QqWTwh6Zn8hX0OKThKXowowavLHiKagW3G78pW7qSShQaadUSRNNEPjueSO6n0Y/b8BoGwZzS/
YzCR4tbC67pEchfj5dYxVa8TJj2xU/MKXJyHOWUb83AYS3Fi+eeZSlJyFtAT7woqQ70lcKeeh8Lo
/4jeOghvkUQgPbDlxMV9e7bWp2MAUt6pyCZvMVugKBfinZMWGYbMUX3Z32MFrLTyMn/JJ415AW5d
eP8sRMb9wDu6qOYK+3vYmVBGybOuF+YffvJkwWHouAsccVuvtlPvy2jPiiajfYwIiMCiB/RaI/uC
hX8Fqn5poLo4sIdwiQlqxl1wkqLajAI6Syu6cEy3zjuWmq4j00cjZ8+3pW/7JqV1RHPhFwQCI+/p
Dr0ym/QYzTc/gdtU9tt4ul2Z5YxHqTHFdgbmqj4G0ENYLRPzo8nIj6O/BS59+FXwwSsgmLYqQboU
S6IpiofTCpbC793oz9CehNwDsSUYbd3o+YbBOTd+c7E2hERnCOOj0Oh83YEK4yhFNrRE44cTDs7G
jWuQazdoel0IbwrsY65YcSEaF5g/Rsxyiak3gasQuG2bxLuHlg8QqG9wWtbRM4V/GOJBV2esXSG5
qvISol5cA42R7C3fI+mFKPCh932JBprq5iZhNVMKuNiAN05eEA/73mJPWmNAQbXyyo6xJYgAtBZr
NknArDR6QEoxoJEOf1xOTM+/lCi5L68kP8T7xgpXjorbM7/GFDuW7mI3GeFDTBPV5OjvL66iIEmN
iKdymlyj72Td/WzlXUAHvBE1eqZXO0mWUOKG0/QlXMiTcHMp+i7b2gNZkVt6oCdSwPiu1vkxih4q
EA4sWwsQZMW6DR2r/aUsEMiZXRsIZzgWXf6AE2dbI090A8XOzFgXYkVWdGkXWM81CnGzbHH/QurB
zs9Edoz5S91sa4wUJPI4UkzMUJNT3WFIEvB3aoWFHHLw14lxyV9GKYognnnmrA2jnpKtzmgg8nz8
D+4vK79hA+vwgUwA202lUEQzSg+z8SstaANySFVEvocyBPdCfJtxuhZ6KDiCuqmzYHmNIOfmP8K7
1Z1CK+TUnOZzGJYjsOgdb5y0D0Ofd3n8ZIOD0nDedAgn6He1C7HmHn2Wr6iVVxt74VbosQQwIBcg
wSkt2gHGu1JQx1lbXMModp5qqkaCZyS/US6B3LRpnyQ69K/uO9NOJ1Ngyd2znHyRbVlgyKrOmNau
L2Qs3dup5cQwtzhpZL4ku4d0CJ7nAofV4hdiJJBaHwHwwKVsBX7nUHF0XgLTB2GYZEiEtZm9cKJL
HFI8gGx8Iv6BVFhqnIR4/e4DdPPT0Knmvuj+OcUxDWMR7N7YcAZIiJPWPsmZbXKoM7zEaK13StMu
A8VYGkvoYd4CXeoRwZfX5jSOvj/5H4b7aRb3qsWD0+mKCbZ2geLtuhd4Y651qiISIYUuK7pTFtSH
MoX2FMzeoQgyxv5TzUNlbzmgIE0sCX+Zc93mhgjhRno2dItcauVmUCaQIOFMOE5PXkDwgmcyNw87
Bhh8KKIDnZrOr0Q1JJMPy5J/72VrRQBCzv/2QUuxiIzXaUGcQmdIsYXzNdSIpR5tVIcgdbm4bGey
yU+FUD4+FKCVl52WAhscWStPORB49ds5SRQkrKKDDqCkvgDWQcOKhOCzrn4cebuAVoRclrB9/DYv
tsj9l3LZwjs3gnAy9FdiXx/NtBjoQDeQ/w0evu2K9aBss6KgbuoGNJVZf/Nu2YaZ2whd93QMpbN8
CDHWjgLXHoT+the+Rk7d39SOxujlUmBAbjxVVhrhPMVHS4ArCR1D+jcHMp+1CCsVuXA+VgqZzdOK
g/Iu29gDr8kw407NyWt4c0ilciqFn8xhQu3FDuls2LoAi3l3FbMTgBHCJlNMA84edRdSRjxxq1XX
K667Quc/Q4BS6XsFnHJclYxJJWMq9zU+u9aXQc7al1jVykJPJ7ltEgWyHlSuaTd9SvolxR6jDrS9
9flBAXUKN0Ht/KVccS075y0vAm/bIt+x7CRo4CN8ITLo7pXlJMkAFbhJoRe+ufLQvx4ze2YcHcHv
tjsKjeJs1Mm9iDRU3S1le7AaqAYZnO6i4gVMExu4Q22OkF6tl/PMHfxlkuWNNqQO47gMLTQb+rfC
eCjFPwl/uwaESG1pC6XxQxHDjKsEwIRzw/4hF5KDjaEpqzjjSceosj5nSm3szNrFRkjqI4W4btWQ
cG3Snv1F/j7p9k/8Wma7Js/eH364Uv0QEnX5spn8eXReb6yZ8k0I/7l+DT/w+fxahkGR/sJyYIN4
dpFpoR/dOmuqrDOkIw9nnKaSMNAVulZEIlHAnpbuSQGrGlRlHpGokW6JCIacZJef7NN6WxtCGk1E
4u/2x3H9vAsrHCH5GkRzgr1r5IQz/78SkAgG6euPmdH+YTNP2dFDKhUWqJvCuCduNOvvhk5k4sdA
mKEvBxVhk8OBP7AXFc4aH+Q3f96kiRTgjOMgbZ4TImV/XwTBgLkfg14d7hk9G2+6PbZgufe/XoM9
wWPfwTtjKyHHPnByRn0onarQ2DlksdqXZj1Kk0Nae/pDNK3Y0uBWkKiPJ6Q4oMS3IUBVS3VTlijT
x9Tpi+ZltPJFvlI6wxyO/GUyQMWUjSi7B7khQ8VTZQB5dq4xqiBMmXSTTLH34WAnY++W/0Moe9Cm
ySM0G00We9GO4KwRyzYpnv08qYuqKf6i2t3lOve1j2/bObReFNicWf6KadkXPy58h9ulhKndih5T
d6ThR6ISbPrW73QnxBpWx/cpg1c7G4huATCmRkwoJlvB6l45UOQVJ5zxCoTpihU6XoUJUR9Vkejl
QIhfs3DBxj784PGS3EZRnHlhLVj1iMUU70+Pca8oUhj8iB+z4xKgSMaV8ca2G/1kFvXJDCgm5z+Y
Blk8r76ZmMBeYfwZiZKJt07rFfCosvBAw1fC48niJKtrSRHRsoAZ5VnklJcoGufY/lJ2yzqz3loA
IKUczeg4O+VsRRO/HvZqMJsm3+jV2z2IIg9gr3d+ssu+7bDiCh0wlt6vfy0vVDwJnjDpU5Gj3ZAY
g9v7YJozxVlnI2ttmJttmqk505Cri/itjI4TGqjUEoe1ytbRd8g1H2KyvR9150SNKpmAicRStSAx
udzX/MBzH84eAHtyP3cJDISjpvQ6QEiVkOCBZOCbva++Ef61mF0O2+vwWZToX0aAbt3WKYkR7UL+
4qBrj52Toi/A0z+IgZ0xNkCNY6g5M/T89j8JpWmBOzg8lnjCK/iJSIt0n2yiMHPubp5dTKazdkZA
yRb/svgmlOiwHKY1QpfcX40Id4gElgc8ZLojYEXd7HVxkQu9YjIvLMk+yvQSAKlJ+B+jOsPs6NaP
Ih7rC4pd14HWNYCvnQQwXdAMdE3xKNHRNCcOjZDxIBp170YW5TzZImaXww79xbzzbZc/YRKIC9Kt
qlcuf+JAdoWe4vbTma1XCp7EPw3m22ILIuuaMkFZss5ANw7TIEvUW/OxdVMxQ2PrQYCmBET4+ADT
TwkKZgm5d3vPy2xCY5zJIv+JKg7slz07IizHpwB+nocybC2PpqNL0T6Iw+dLAMpN93cLAI3Rmb8+
7nUBbj10c/tFACDhd1Dkfz8znvpZsYXqvaKOia3G0Nz4mk2nlMdYq+4VPKVNMYuivIYYZ2F4zt3h
XID91jjohm0qhw8pYMAB9coF6PNY1E2cGBpxlul1pAvmx11S18fsWabi4RDtwuLOI/LbMgnrOgu9
Rm+ar1D2dOQx52S+tz+UquPyz1OORtpCxGVhhTF8xGght+UbVheOQs0Ay6Q5CPZWIi7WvI3u8A+/
BTaSgr5186i6dvsfZl3SOnsDYQ5ZFNzbjtrDkVHUSIrxqZux41ATUwk/x5kiKuBgi+0gFSAox/T8
djZZM0qTAc4goIjN2MlZazLVdktcpVF+ydCaD2tM7jnQfSFkXc2Nr0e06zNc3gd/SVxeSQMNABvU
0CULGYyCof0ikwfcryyiGZLgbx5OFw66qlfzKrj3BJ/stqZPmXBtVyvwWO2xmUSGtjyaIa7zuDMI
qfLFxiQa8MB5jwpai/ynfGS9fDUC9Zb2J1xQVJLpwGG6DdX9b7X824H5h/UJM9ywlTbgoWOV7apc
KDVE9PYC1P9Z9oPC+g2LmBlOXx15gGbj1pllddr/n0CHGgC1d4h74mM/FJY2qoKy/coBBQv1Ffw+
Rd6+TPXCPVwlrJjwGih53MfcxrXwi9PXvRGCYAOxOGVPnf9tujK30hMGquECfZzMDJAdpV8rNDaG
dBbP/m2TAIQzopv30q4rhcMZ5nSKZMl3UQ8AEVWjKDzuPCvHVFO6q/JOv4itjpGDuWJ2EgCxYpk/
Ist/cw/x/AYdj6BVhOz3fvTCrngTpxg+ljC8dpx60DVt+n6ZWjeKyO4tGltiUUI5RSYs+lOLxGeQ
A9SJP37hXD7vNaNuMo9RAlzbk1nSIc6I6PEaYEPNE4b1CIwd0FtEO5GuNN6Z97FHN5axWEoXW7ix
lDol/+J24eMQ+4OFcP88ZNrRqq4Jk8NkjkizEzbSdpWiee0kqa287FeoHn40PNvihAq3qeN/qOhs
sNS86f2gLESngGwnxduE3gBCeUhYs14ydVaQ6MNWtqGrWxGU9uyUf8AZeeqdLgPjbXtDdcPLSuk+
SBC/jLNBhBrwixKeaL3RkcvCwEY+Ff/7P2WwLfkuR4ccwdJRkkGo4LGXBmzJxdenLUNbAthbilB0
Al70IcWWIwGRkgsV3e/BlI7XMwYSvYnfA/1SKEogQNEOv9w2oL28jZXxDBj0hggrzkRb6Z2+SXPV
cjh8qrCKafAZe7rKarPqd8971FThJvsf27Arr+Pi/xBHpsUeMYu9BNhsPfJkjhRjL5z5AN5bs8dy
MMYWBIoRlNk4A28OcxtY3L1DHm/1NBeCqiPaAor/Asq1IoY3quF898AW2acC9qllRyUkgIuVl389
gx8v7bSV0P/MM2ytucsgQz7o+5uqKTSYVtCecjuYAzJF7jJ8H5EIdUGBzgkmONiMTEhKbeFabik5
s0MXy8c+pzHBaL+So2ZDFxhAKpy6awXCR48UGZZMEp245LG2iKgIujYGidvSWltYnZIjI+XdhG9G
WEQfY4ia1y1Fse8P9uena3FJY4PAGsuPziww9or127rkIa9aHi7t30k/8vPaxkoUYe+mHMMOOHSP
o5si7usS7LUuS5tOU+TF5HsWL58Wi2fa8WJr7W/sM1aQrDmls35ZvzuebICA2kCVaI85gcRtEghb
aQKwRGYV9zmUv9mUneIHnJTiRHu57Vm0ZjULG2dNBvyYXoTwXOkW5kZUQ3yEuC1/g46OW/ldGCM8
iLPVyFP8NlculAGULwUEQE56jyB9HdolrBJHW1CvwhnjdQbQRcxIIupts3Ij05/ADxtc0jAyya4G
GcBHLt247qiMuW7aVz5BZeEGjNS35ui4O/leRZJK/2YhnIoD0mzmmog87WfgmkLdZbhXr/Mx8LHB
dhRz2sN5Xrg22TLsGN3rq/CPg7dKIxaHM6xUxH0SrlpABXj3AbFHN3erIfueHVraOTGPsK4ncQ0u
ZZ+H0V47efr9+w0rSegi0X3kZVtbELuuo+rzo3QrnGn0S8WbWXwDpAyBIyVcyRUAff/dYnrNSBws
fX5WHPnTu+JX3ti1NXFspfPNjSGKV3zFPIM4COsTdaPRASz0hREuoHAcmX7R18SXBA5RD6nUIgA8
/38BR1zqlf/qxS23CcUE+e4YeYVGdtv1m2YyCMfrDBSmnjn3TFaK9jhfY8Yw5jWTFZGHfi0+wtVx
/pbSuXN59ODlankPHCGQyWk+hHYo09RaQffOfUnyuZCSl6BnIEOv/cyv0UZHcpNpOtq+rALCOri6
ThopKqm0MRkEiu1H/CmvYuavK/bhq9dG32pWTXqt2ZrR0ehfiBLLWmJKMC3eMqIyRGqzSvurlbP6
/mDZ663jLpd6wzcptlhvXcAcDLtJkvOSS9njJJBfxl65E9l5DYNVam5KRJZtMvVMNIxn4RT2w+4C
N0+cgiXhUQ+sbhgtZqN41jTGkW6ztrVxy83EXQ6PjfPvMbMcjhike8dniPr2bWRDgFN1Lt/p/AaH
7uwZTRAFeY/YDHklaJj4ckYzhGyY/BMlWJJcF0F0lF0cfB5uFmf40n7OUb8zQlz//t1fI7Clb5Cq
Eb/0oisfsEzRCLy7B9d6fuMdtbNhaCz0AGpN5lwn++rjaCONmDJqIK1f9mDiUyCLR4ItC05xL4S5
J1Ww0hkze0N8/SnFPDmKXmDe38dB4Q8gfUvKSMglRu/lIiM2pNoLvHpWoCK85jlVVkWrNExdve3J
BqruZ+814CZARLGGr0fVkU1OFpyY03g1nPeIWjHuAcDIS8Okfm0KLYfNGkKc9yfTnCmOwMOb8LkM
SdClr/sIGj/jlrdr1ymBNYugvjq7iB7gANYyF4Uqztm2KRoZcNb8rFhksJUQIsJxCZckieqHViW+
mIPfRBjH3fAsVIgHbDnFjMvvHYE0lrsI+rLJ4OaKGVzV9bASxz8Jq67/CNwJGkhhn1aemDobRWVv
9NTJyuzx5ebCvTEaSG3VPEL4XrsGMuc4lG4cSfDaHDjZMgj8DC9ehTCGoWDMgNwNU79d2+doSpOr
dsxuNbfvEAgeAyNYmExXP2O+T8dEhe1bvw9Sn6pyhKIVyep4YU+09vHVl3N8hqyAwbzQZG+MRcCn
EiR7R6nvUAFTWiKmK/4kGntDWYVaiI5CqvLNatOPgXcyoL58CeoDvfjUWqBXqm6QIIBhH5ch9dlI
iHGMrkFXnI8AVJuhOiAuf/Z2p2npYy3HeYNwCF8/C4rtc0KnvRUb9dgB1JO6q0crenTgt4axoNkf
VR4+EAQvjThzYG4uzDv9qnTtyQo6Xz7zf2XbIqFVi3mQ/rv6CJz06pqFotFdVueGeBG+A234+5bf
mHVscrYYUT6+QJlVBZ6Y+ZEzVtmf+iYqLWvzTvvIitYfWLle3wTQ5Sv9lzSK3HvoCG7DSB+Gui9y
xxTWHangpgJN+mMhT9IC2LpuV+HCxIkk4NDKN39DUayypwmh2a0uZUOrBYCQo1Q5C/VIRWeyzW/5
ggx6R417C0J9E7S+zVk591W3lOLaIgXaH81ovFqKTyv+4j/HzyVK4Wg/pmn1kaR07AQcuUJUwJUm
P81S5xpa7Kq0cXBLXoA5frT2GOCKmQDoECPbPSyOBaypiB/ZcrzHk8bRCxRipEyz4807b1d0YZYY
t2rsZnYQA58KA9w7N6yKuiry1+iTxgcmKMU/VWoM5tAWYdB6//rMgs3wQdeDU38z7nAw2P4+fKIp
aGtb1IHOOdSw+jsM5+5bwcKJGrwIcZd2DJ4i7GPG69vD2UFZtxgPhx/hqGZ32U99LT3NqqjOKxxg
GYezWaiKwKaZhpKnq00FmJFrSWhiu17uHoHbkDEyIzgii+4wO9HzFWLjg6lwfJsJBnCsua9sTlEE
9fSehicIUC0ZCZrKf0RC8hY/Rg4tbfFGYBkUi02ZnE8xYaMHplgCBznPBQN2tNlCqopWa+f1cIK0
Xy9Agh5NiV5YOzCtn6yy2LSWHSZ+KC/EezqK0rQ0H11zKnarPxuhihmOJtMpjWpKnbfoFEvlOWuH
uWam68JsGkL68QCdZ7zbapAzzKAnE3EkL2LuufCGE6e7rsEq2lmYo/7uziHYdS5cI4z/rYWxhFr0
asAfAjh/+6lKroGt6trnfcUMIULYVS1tXUbLWt3heG32YEov0wb+eMnJOuQPKKN1b3l4AQAvVb73
/Y9m6MDk1hj6QAG2jUKoHHXI7QFlNF9oJ7iAJt9LY9gpE7/2rII6jea6E5ycTX3tgieSpILBPCX3
L4VReJ6pK2Sr1+pNW4OYEtxdJlYxD63/FnrXt1Fshu82JS/HqN2X/vD8C0WyuSALlvRbQ3GCrbqB
do5OS+4PHkcSEuNSOh0U9EgX0SwOEuEP3wdoaYsJHuoDDarrYjFoqITZ6VYsH1ZBS1n8CHSnk4Ci
1O95RFdVKilLFvVbSofY8WH/wJGBW8rHZj4B7sZ/0T6CrBb3TBlwpG8KQwJ7RF98YIbGZcBm6L5j
T9rfdHVpzVhewxBkvQu9E2ttARWoc/dAP0uazSoL+EnvsBf2wVGhN33lsl4qcJ1YH/e9If5QNceY
yGrWb5/yhOIRdV1Hz9EfMC1ZbVxFUCJHNQutfzsBs1FJGDVhwpNHKTqF92HjQ3+JMTQejmwxO719
CBLIUAXdKSVcgVc7KOsDBi0/p/IbGsG+CYFb8PjAz6wp9V8i/r5mdknpYJMVFZA4wEUNavyOZxv7
SoY59AE4xO0O2IauilAX2LXiFKSacrqG6Y8a1Nk+xCfGoCDbA5VNrrB3CfJXMZiguHah5EK5IgjK
sC/Y3W9jwawMrBwKSWwM8e07ZRdH3ZxZLzMrHMh+kkjvtnYnttU6ED7fsmGQ+gmR10/1qwUeopKj
lwb3zbYC6BqdwnFtXAylrVwj0GR7XBSlk9YSWGbK7OfPDBvCwIsgoaGV/293TelPtNOrs+HOxH0F
Pk8VZsSAgQto0YBx5mkaTd5t6OvizbydyfjDG4+SypKUM5AG62sKppCIk2jmC920IN9sXsFoCfx3
m7Gg/xq2CHq94PntGtsww9bTshg5dEX0o5GM6FS+LakinJiqyFJjko2UKqCr9oMMhRTymw72S/6p
p/lPcvPx6rUG5xEbfQ5t/92oPzZHS9OmQzjMtIC+TcC64n0jR1d0Q1sfbZRz2LWj5UCbgyLXI8kh
ZkHgA9cqSXj2PIy5YKQ+9m7qQcW1rRuGPqQbhpwN8DIesaZgMzuZr0wiRejTWwWqUxt8Dv/pesx0
VmltVJoT7yKyTyNQIs4BD/jXy2bHqk9OtvlKGw16Q8MvVQ+W4XqYB2EQCb00eOGj3P9GipulmONO
0yT8EFRn5QvQB9IitOtSFdhhfdhSgg/1YWDXF5OiGKd7+HZnmQmuUlZhVEOukPvqrw6luTDOskO1
5DD6R0jBa4wllS35A2zhJX7b11wKL5RQqWxlv+9hVxjA2OCa1arbZ24UpFOluCvxT5X5azDhx+1w
cZGiClFEV1fDVEJNm7R7bbC9K7/ny4nNx26Oe8qfG68PxBkMXYbc3fCtZD9FXr4mR/6Qm1qtRuMM
zZPiKGTjU1WyTG68hzgA5BT2ZGuoUjZnXm90SLaG6GUaXwfBP/8K5Zs/YhcU9b0z4LjavreVJ26Z
tnjrwokhUkQY+5F9XygTPk+xttmmO/G9YsGcbPJCmhkh99It0sqCrXSlFlADmjeMid+Rs+0Up4G0
a+wYlLtGUZGxF5m6YepF1x1METikYj/Vn2XrZo2m0oVMt13oZubSt14nLH1791Lc6QHsh9OTQ4aC
hA+gf/DWdV0QA6HG7daELpHhSPbcr4NzU/v5KQFlJx9CX6EknHNWr/nAGGhcJj0i9Vd5fz7KI+sI
+Igk+2i3trlLgkKyzK2pNNv1ZAG92LzcM7OAhCddUabvdj3dyEgnDrFq7Y91smhOKFn8rMlfb9GM
W/P5m29y/LzpN3dxb+WKI9wxzBh0YbqqQ7qYwFrjY0eHmiSg57kwKC8/QBSE8F9FIf7BjQ1d/J61
ZnJdypWUR7dv0qfgXll15UZtOJfA6aVrDm+eWN5E6FvPSC6G6GupHbCRq7Ko0lPCwPxSMKVJEUW1
QlW/N2/tiw3phXI6AhSQ7Tt+BBNUrmEtAPkyetuZ/ok6V7WPLoitMVzC3IQbFIenWmLyjpiqOa0m
lnoGOBIhJkjd+8aJXh+pqNk9S1le/PGXFhQMmniLnGngt4FkOvk41CEEFkZj+RkTiJQsNumz2k0o
qdKt1SVjL51EMclKQq7H/O/pwM0Hcm4RxV7HOGqel0iWqMlmun/lz/DfvYz6SiA8G3FnBPcJR6OR
Fw45UoCpqn74CiKtlz3B15/D1yZJKe9/6SPqJwlTg4CzLTNrpIMtDyQmpsw/Z3QcZbEicWS8LY83
gKG210J7G+e3OwKMuKLDBo/+GadUiCXGG2prWKtvMcb44OkkLzaQSjoUMaj9zCF0o4ipzwWtveAD
IEN6TDyv+2KqAMe+iaLdxMthPy1Su5wDeTuotpM4zKs5dpB+fwJWElPnVw54lUyOjONVKFbhAo2/
TfiDgIpIc9Yk119tz+H+eijc8xTyUaLEY04bXj7dov9JgNX+i7m/eZjSJdUOl8087LEXMqOvuEGp
vqU3j2IBCcHsBfjCF27scPpC7RG8vk2LIaN58veBx6YTbJw9n5TtiLfAB3T7kHUDfUv3XoV6wwst
50fyws7z49IKl2S7+K7CVtL4nKdYxrQqyVJXqcNXf9RQwXvlTrevPCtL0puMibussJXbhkNZJdqi
GnIp0apPuOTXowt9tsbZLRFIDW+L1kTVu7v5zatDI4pJ3g9JX6w8RgWp4Ob4p33Kj1dQLf9k2LjT
OFSJ/ADJi6HLORVQAl/ou0Mf90m+bJ6KPFci6LTyeKW7aptHoduUwP0GpZ5y/lDd6M7M9ahiarCN
ocViTIginc3DgTVK5EAcGpQuieKTOXS678WmoPBFqni2douTf5XGYRPLncMIAWY3vZ3wDAhJSplp
eFAjNZALhBDMKT1C0OauMXdqhaJBZJkTx+TpAJTxQK6YQPvoEDGpWZjVPL+AMHUtpmo8WlLajN8X
X4igYgVp1J2bDzdJcarXql0cX2Gz/xXi+9zl7ulM3tvjtU3np34O3IHrouKWvwjBN+QF5hbTYblc
OaKLtywE3SHnkYYAdicHORHDYjBEjrwmnVIzju1Xi8d1p8e9sHyhDjHWQuEzoz1NTg+QY1E/yIXc
qoFcEobif3YnCalzhJCoQU8omDGnqQ1NkJTYgUF51VPjwrZfABRNhw2dM89PUyB/gEwTNmLyrFEp
XejaN2U18ic12titdg0ugCTH4eEb2YA7FOq5j+KgCHZBxKuse1hegU4Fbu7/8I6fhuspd2fyEDrA
VjJUrh+CxcGd7AxeTxuFKX2qh+5lLG/21RgScC1J75cs7cUXdd/+/DndKBe7RvO7OSA2maQv+eWS
hiD1p+XJRD2kyqN3d5EPQ3HNdvEpWDYQH8w+S2SXQZORKALSl5+wHhUNbObXO9alULx02IUlDzYf
6iGprroLJEhNpDDLuHcYRZQIU5Nckw133VrUjRhGp5tjK8Y25vVsU3y0Hubu5w+H53fYOaj2VRiJ
iaxLiI407a2NlHLKnjZP6MvPA+yvcAQlaqrLddRTIFNdPvZXNSyHih/W67PW5D6mDk509dwpMbH4
s/b6FEM3fbwCxEqvO3AF6aglEj8Ia9Zl3Hq01UQherjIuy/4Llsaj2YFukWCDzFpwh5OKNkVWWd8
KCTQkRigIoPl4wMSmyBM544VU/5uPTsUl/pUuOFT+oIl4a7Xffku22tUs46N3lQE74Gz0SklRe5m
vAnSChg4wro85Ufbg/pv70p4RvLWD/hDf2xy7xbVgFpzi2mAfYMefxFTJq5f9/Mu3WIAkPbq+RMm
H3OXiVyLWdkioTOzXne/gfX83RnaYbooSLX2PxdT4gX8qsQShwAYLTMIEZCoqdLw7nEqkLaa5KfX
J6n2n5p1qSryn/DuMWVJRTG7P09qduEh9c4qbi141WnnYKOQoZJ+J5hK4uxCRoCidMcLKkwtwknV
2qpIOoeiqoRpcbPKId61UDoDk8OGnYqUznpddqWAHAEZm+/MKcw+U0t4OQytU1uWyFHwFDG/Aifn
yLFKHC1ZnP0JvV791voOY89q5o4BCBEz8z/gfW8AamFDY85zl43VlRmcZsMdzQY8MVPYcCaS/rND
hKs6PAEYlE59eAsmYLV/qW/ba8ZiwXyVHyjizCqbV4EORSUmJbR20IdmskoyaDjJerJ2YdKnUULL
wQCD8IPWZJl+jOQWBWoNPJKjFepUacaPCDNyV+IM5pVnvPqgAUUFX620swR1pC8EFj08Eya3RM1q
cnFJREZ2M16z20le4s6yJjE8z8TRve1Ln0b7DpqP+kvgTaF26hk89wruhk2KDaO9umU/FL5yjovd
QeQtCCPIVhSAxln1YzymyMO+oxwZtgdyTun6T9T+Vs8TgdzfvODTKIpygjfnRiWWffUELngpkKhG
BxnwCCs/Ng69++RbL8P0Amt72Tnoy1HSKk/Pre2izJCgKo4zci0NtBEFgAsbNnxFA0oS9jIHG0DJ
P2TSA8MRkzELW16NmIX3ZSDE/o9+s9gqSdBkRzgr6Hb1DBCGmIut8qk0Q6U5pX9nsfRwkfLAo+eA
bENxaRuJ/PYjMK8Tp8HFC0CNoA/ti4mzaqF7O0vb0HMZgL58blMGlSfwAqkvnLx7k3EFoJCkogHN
gFxAYt1/dHYhoYibetRDWkIVBT5UGlq5SpdzQxCrdHoVmZYW2GiCBjUks106p5gXAJkksNjS2I5a
nbyhemco4Am5aN8Tb1Cn50L8eRd/4gPrf89NDIml3MLpcMLUo7BNLtaR/n648OJFjVVhmyaf9tvQ
NNne1uEMpW02CNaUsxLNFoBoyioSFEbB5gMGAjV5egnjLvD3k59N+itlws63csKgrQWOBTQlnYh7
cdHoTqQc9dq0hM9hXixCrgE9ArCkd6waWM4IRHRPnhQOtT1GAaQs3qvAxAghOdf0ZYjLF/6CNSXF
SAhkEaXBKyKLI9Zziu+eiYUZ06gvksH/btZ0xpewBPmS7biqRA0DgOXwWWVBRK2EBAbZiypVzElo
utCE9lGzUY8WKTGOhfpWcvt1Al3CyLbSdJO+teDHe/KMgaUp+mB2uzCJyMffGXyDWJ0KsxVDBNjv
mLpYUEkjxPcRirRGmCLGLxIm0RUj86vOCMoLUSqeEo+eHmu6VZLGGdMa0gU4+NhaPeMalkRNBKS1
kjbdCJfxbglNjpboI86t5RXolS1ovfh6hmqSmBjDBNnE4UkCz8cB+zKWrTFyasHWQrz2p/ovuppn
OFglEu2FhJSNFXcEuLRhLJWBHWLs0wBzTzLaz7sFMNiLD4ATQW42T6H42/Ykhw23a3xk+nlVc+gT
kPGdCvK+MVtd4mlSfYmxVKaXvHrlkRbnDZnyeHrhc9pdW76cpnh+oTB2A1JBm7LWJJIHPqljzyvU
TNty13PrS4uvFfoXDsjtSD5zfBp1Rybw2+ipO3ZhYOIHjo5BH7LhTO9LIldAUtSgCm4xrAAi5z3E
8S+5Ykovzg0Ix2nBAdwXEcG0n66tMDBjSGDM5Vh+F+q6kvEPiTpOpvceak+HCYZ24OdVSPzd40gS
3/IPrN2iKH0DN/fApkQ/wM54imAWsl38iEn4f3a5Pfo1T37ad3MtQiPWxOBbUE6rRf1+qA30UyZd
iE/UwrdOQmhkeymcx4M/8cdiUWe8iPuOJS33tF5Wn7csefXv6eIcWowY0cWpKtjwzKh/cP3emUsx
7zmSTZVcEnvHpgbVZERpVjqquJ2MR8dEJ9l1g21sIqAo9AEL3Guze5ATz5L+pJYZ6uKPcKdsMTzj
HYeoEkk//7M6YoaddepTvxo0ost2PukX4877QAs8YtO/18CwLVewdTxjuOdJTIZReqI5JuZWVZEv
Sr/BML7kVlCvFHhBApI5uEdJiKESDmMJKyo8WqLLzvxOHpOq0Szt6DDPPcTZpmZnBWzeipW4oj8q
QHuU83XS5n9YnYYF1dEwvIRy1aTyYM+rO99Al9/KRZtClG8bfwwuRVJ4VhP1iRwtpxqCM6ymk9Gd
WpkAAyLOFGJBGlZDcaQHy3X6xew5kFzZm7DcRNbB0bljl9RTFlsbvTjfXexFVuqyOxk9d35OxsoH
7qFwiNmosWYxH//5A5sLPjRUmkMr8jdnwVb8m7R3WgnHtcL05mlikWJhQZtokIYzU5oRCfokNJY5
1nxmAVeSrVz8ieXCuJCxONTkoCUtz/DHht0FfhJkeWgR0OnhdxjhmPP6U0GN7WeyVtmqmcv3jQKD
FbCzZ1XxSd4Bn6mavoh9+Anvtx3GxOL5RtSoiFTajh54DwvG08wK6wwxg1M40C/amtwxzmJwoWDC
h8dQDWMBAGDdoocgA5o+9yLmRkYFZ1XmMQo9hJz2xP3OnF+W3m/bGaXg3yoAQomT2yHYBshnzX8f
lDbtXxMZl73EqBhxDmoRwJopbsIOY/JuJyIfF43T3b7R95C1IIh58zE2A/v2xsl47curK1UM/p8l
kXfymTY8JXeLexoJ4d/YakQGaIw1puhdjwbNbl8F256CiM97VSOKQMHPzyrtAe96ggXuCOIfVvxt
atClT3zwa0MpoLXkKEhq8HRCh1U20CYhkwzJIbGaQqZBGAm+4fYNlO8X/UL6h+p0q+flEHfO4BBI
s0GcEyyyd6LhCB+hKEGrbxz/fvRs+DtZ8dw3iLcrzG6wm4gYDzw8n97KCH7miJ+XDYwAGiO/yJD4
yCcofS1M/v7G15LR41tbyxm9vrUymUGE+eW+3S2TW3t+KmGxqpe8B3wl9PvCM2KWH7a5aGA/qNsP
tUhm+IzktUfF0m9UpOBt23Elu2zh6OTfoD8O+QhFz4OonAPNee/YTRiFOfSu0jph1BdQkLRDiEQX
aOBk5zfyrPcmgz5vzc6j8MNsOpGOY8R/5UTgGopotMZmheD5Lko2++lVAyYlIS3eR+ztfoPpSOdX
VlEZP9I/ceqR8s+3qsHmhdTYVQGEHXO5L8ZzSWDpXzWKO28TPdLDnbzKyFldfHaxPN2KcQz0WXzD
vQFPTFC0wqFcpGltQ8Y0znjwGXJLABCzvWFluLHFPdWEinIVmKxvQtCaL+k9xhpLByzXchgBKqDm
SvjIPiAr03gsZ6epmjRqnmoO1hItXHSy/0H04HPzMb7VYjj9eQ8z//uFw/i1S3/BnqeAnEEu1D86
wdrLsvIcUHzWQ+Eq+iJw3p6teYPYhfgQ/y1uJBl/x8qnHi453JrQMrRW7mU9mYSEyDlLrNMTrBWx
rGkVHxtBszuGMjg+XoCABxyQPa4BZvIHRcNi9410x2clQDruMJTDg6KU9nL3vP7ZIE69+d5JW4ZX
UjH9+qp75EOLqItCE2kjOtuswvYKoZBy6akrlXaRs8+apt2j/5u8yhtL3ShH092KuC7xrSQr8n0j
6wrF8tiHzJax/sbvM4loE0PnTIjCo+yu9fWRBOtJK/N+OBAdtD312RbvNfLKqB8UIJ0RNwe+aDUJ
iPWvsZoZp75y+nMUKbsBTWJFEJ8GU9FesMS2qL6t3+RDde8qEk0ZZuDZuNY/n28urLenjTz5Ju4D
PHy5feolyALsPGqlWDBUWpOl2wcapYl3f0QMBFvp0WqcWSMTt50H9SOUWaloMIvIhs2oBMgE+vPZ
GegaK6k1nRZBExKIzEQi8O4g1v6yx+V+XBiD5QodiaCxhRCBTE6HaTOU4513SH/dfeorvcYqQU+t
2e3N0FiaZ5eksaim7x0yBSzHH40T0mT9sp50zLj2RYAPc+3fGeKxZCzfzyNUY5ju3v7U+EZoy3CS
7MctoQpgSgan7BHhjoK4LXGfIfGnwfXMDq9tqaL1/1CuKFADrzTI76W677TkffeFconp0bAXv/yt
cHGT21quDpH8qRFexLLIzVXwb0agc47aa+8E3Xa1WcZeGZ87PBRcFQ9YuU0ZHRY9IOy4mVBgpFoQ
lGYsEttTvKYIVFNCn2BOCPTORq4nktOoL/cPjLRXQN+72YsFfYDtbjEAdFHPOn0/Vqa/LzJrnc0W
yImP5y1EfKu960LPSID/nolvds0eZ9Kh+CrURrxAesZ60LwaVfrr8WVe4Q7kQjnx8qz7E8GODKaN
XSeSnmnVaISmp1ZKS4/hBPYLpt1YARUKYM5jTBWNlckED3jbUjz0wj4wEHIplWIgM1RB/gMv52K5
yS7CCw7iX9jD6KYjs4czyFacM1ZCD4OcF8zK/azHFTJjTR9IqpsfPpMdsG49wg+OnDmVT7rlPBPK
xVWVY2sQaqMQpmLSLo6nqQLRdf6lJQIlHpb8y01AphH+001Zo5iB8C+VFEjEMA5GlaTBdvhhGzc1
v8KL9xrri6/m7UlW5RxuVKSqlyWSf6eVLqCRmBGZLjZbgq+MbegPcu6Iy50ICoOE0Cv8wLPVkR4j
XR3Ezjb9BkjCck9vEcuC3RS30ZdPlvq97Umf+dZ78qCk8YeN3affQ3UT1GUXnHNNJuBgjTcbgMUa
3Ql9Jok4li/18H33HKtAovm1ki+PXVbyKLQJTXMzs93dK7kZ553fFFzW1vRbtV57P2aZkYVONc1+
xYtQlT3GzTI+dHwupcUaiE0tqRAHIx6fcpUScZXJ1oFaSa/NGRawBHc5jAHSQ6STX6H5n9uYlrRY
T5PiPvyMQIaQuGtpZBSkC90oFm1x/ZLLu6gyGGck3fdQDknpA3DUkNPHCmOsUO4EQQpquehRlJu9
hnDwmnW0h1m9T/RtuWXen8lPWS/CXWYFkNMXSPHvzNS6jqn4EatApq7LjyuNUMRQJoo+AaRN1bfZ
aAZgv9EcYdrC4EpFtP8cR7lrMPrBRccYeSqZbJAKy0LYhHHeyJgPRiGlD4KQD2xCkrZ3RxXwiEj2
92ExVZVleAlVp+pV0ig62EtI+j2mpWRxXtxnOww0vZF/oi3NQsWUPXwNr+BSHXen7fDEdUrKulE9
IerQCIzemhKl6PGTW4DD3K2qSFqjF9r5Sx7d+16vPfCs/KL33YCdGicTjdUHD4nACUdDcn0OEbZl
LRTzGG1iJdlXY8GpNhXETafMpK340sYZhT9Nw31ytSNRIUijfNQ+6DySfnp5uec4ScYQzj4AAmvb
pWDWfJLQ+T0xNxeXBUi0xckvhnGO7Z/GKeaSu/xZmZjORU8pcLYjYB7ZqZk+ixHwyzQNA8oAfhGx
woGQ3SAcdHNfJ8vSb0GCxyPBr0CAGtMLI6rYzFUrhW+GkRhhZ6kO1AGy5xUTDmQmjOz8KqKTH2aD
KKWYb4l2vJlLHtvX3zU3d4ksB0L2SVO6/2gTfW4APo2pPp19fP3dVPV1x6OQwvWtBrbyoatfJfQS
43ZiUomC5bFW5u+o3fshtT6lRJZT+vqOIOQ+7OVGWYdolGP23OuOrZSzuq6yRmtG4boISlky8gIj
HWTgXxqYYeRIqUcHK1pZL8Zebvr3PhmcgGt38eKYb+Fd3EJUJpTkeTu2ReXbu5J9FobDq7qHIfkj
smBMd4+R1Kmjs2rBO0hfBHZT61h7pSSqauUGTkIePPMdjY6fKXehY2+CIEiXmO0UmWDb0AcMF6VY
u7mZnj/U67e8ioXmYRBxJTHIT+hDkY9HzLppYGHaxL8QsMadLbyD1krpngCz70c8pd8iYobTg0U/
ibNlvLWOW0XF1ej+Gdjai9E+2JH0ocvA1lC7Nt8VV/f1Y6kRTM7B83svjrxpxp55K2kryCYXe/zH
TxnAYZafj/LtbONddFyJ6Whh59vDjrKDigDkIswMVsFHI4RaC8hKk6Gr+5v1/HhG4IgoyJ+Ch1Wp
vyi0EA3F1jWPWayvgnvWyAVNJzcGD0an1UGwVEZGWMLhg9BpA0n6ovIwXOXDXwW5V4sdFBYeXtiu
1SK4sH2zOC1Xuq6Dv0sMcZJgPh7oAuH9TVEBsS4Vpr+NPpFczi3cZkmLfJ9B2cQknQAOCsMzr7M9
3uXx8Zad4kR2UVzWPWUO0QM6s91Ujhj9UIu7kC9pbaYw20t0dF3nVm/ixiwLlEPiULImlOzDzQhd
6KYkpI0ZoFLP+u+i8HU5mxx6CyKrEI5ojewwjhordS+k41QJIbXrBDEujbDhyi6jdEZhjv6dj2m2
47ZGaAUipTHQOAIN/jFMXo8VNV309plLVPLKoLz3Pg6vq+zAl4A9KdssZQ3HPen+HTUlxb737e3l
5JM3Yc/u6J8ORAMBwI2K8NfzwkG352XfARfbbrttt17ZyZEqlbyqRccZp4BaBo0GPYVbfIoKW2SK
cZWBk4G0KikQeEOlaKCUgGaBaI8WGWYFwNmJFY+vOefU34bZfm+WnTj/xtnak65LShxQQUr8Px9x
GZ3+8sIBiNuDvUezXH+OfQMyM9RsWjfJ+sPBD+hAz5iyB39ktOdWIQxolOWyvQKPX44d5TMP9VXu
CljPCZjuLcdtOVVmNk2a8vj51wxfdU9dt5Qo12bYIoH9ReFTwjRRcZR8XVnDDMh6qBlIT4YPJmBs
WZunmxyH2wB8gPR3JOA63LQg/YXVjGNkJzzn7YGenRt1dqLVssyCXY49MpIWgaAbHMtpXiWspeNY
E1/5IwmXn9YBMcyrv5FC7XNORnI51dIBY5UQHl7W6xTyV/RRLXt2MwFPMU+3WsacwmtuG2vIq6T+
92p13lVQjpBM6ls3W2UkcXLXZJV/5aKHiOM20Pnjmd4d3RS3sRJ9wUwrlEEf5hon5gsfqO2yEpDZ
QhWUQRkJA35MswaxwAgOrvczVCxm4iO8sle47GeiBhy5WWIPubH3AtyalOc7v+3xLq5Ty7yUKxEu
HDdgTDGFyc8LOXiVHKzkj4Fc5kPePCywQ30j6mUUxrGCaintKj/znUJFyLypnASpmGdWXhu2ggmN
2lMijp/R3bA/EgByq90D3/LQ6HLyWk81ZtXcNCNeeEIGdScPm3Ztixz6MK1mCaTumBgg/bLWNwXK
goGnUwORYnv/Y0CDCYa4ISwPl06Vi5eGmL7+Cvu0hAI/VhtotlFbb7f9cUpmsdhXPJYWBmr/2n0b
dz3KttaAcN71H6jLmy/rFXRFOha363GvaEszrQJMQVjqJd3AYDOTHu5CfrrS83ZlvdCR/sks9IyF
sJxgY/Z/ZmKX04ih5tuFBiv6/Ph84OYjsqz5gUN0dhK6XzDuNcnMndWbd0EqoUExdsPkWAHFGQIJ
vWqS4ugboS31Gm641upY3aJSNUhHOyRbWjscYguUY8Ra3eKLIdh+h1Km7P/cGwS2hCpMEo7pyWli
9Kj9snpo69T3WMOQUddPTMHcg25SaM2unHoJBwxouHoIEN42STQ/d2YMtt11uRhyCJ2AH/QpTjYB
c1p1L2m8A6v4l4Wj+IEIkmU1q1wmPgOZdJ7GCL/4cRdxBGoXqvo9eOzv1quVoKUnaCZqhzuy9QCC
jMoL7QiK5N6I7aqvrK8zPQ07EO5N0xT5uc6U9xYM3a1SSgV6D6b9sSDdIxvkZ59sCXVzDBqI/lAC
r7J0tLpLNBxaXuNxJJRf14ktODFXtFW5O/MacztLb+DmsaBVor5hQZ3jeHWWlJyqcA9N0XLm+rwb
0x0BZ+moU8CDESUwTrh/ENprCWrKEtO1+/WLP+KPzak1IuL8msEv0LocnnuxYNUUG4qr3SRJSyrc
u+cBUnRrLVGNPNGcEDpFVzKstPFalkovvNMHtIW1VXIpC3ljs2zh2o6/jD4CezcUecGIVIuQyZWJ
ecMzhuXkuDYnjJi4k7geTrA85nsqUm1NpLIq/eYROKdDAzbPfPYrlw9vWtR3usjfwSOx/dswcIlx
x07ssZEPbGzkdtODy0CrsEyzTecyQT148CFtYIk+1xi3bSeVp9Hm/euiucyCu5lTttDoz9VzJoX1
Cxo8UKhAihfh0U3iEDAfPQAyrvMFMg5LZYYJy5Y+OSK6H1/gN46+hPeUJIWqwEEXhrR4HPTsGy7n
E3r5YkFWL5uOhIG3hu725R16HM4dtGy8jVFSiK+K25oHMOxXPpAuQdyNPKI5CRhsmcUBATvKr22O
GQoXPeUtUZlgJ9h2aJQ6wFTr0yrGGxb3Wq4MrLxPYr22SELAyp9b4hGunrhcKYeHk31bpmm6hXXY
8Dq9skbHXgqfwN1uHffDqmyF8wu3ypn2Foqh3xHtSxu+SLdhkwBHDOFbrur6gK5ocgHk/gvageGm
VAYNltAA9obMBQfImvSAQVAq85u3qArTTTg73i8HTZ5nPBzz/VwEfM7f8dLXx2FK4rDsKwa5vPxi
my+X69pg2vMq1CImxg3TYAbORrIShSEWpokmsQeryzZd51e8ZFfMMJzE6Rb9Bga3FT0PQIOKfV3b
2I6WAkMZ3h+tr8MbdNhB5wwChydxTUyekPz7X4VhBGaW6F9/JN38yG26Iba4IJAwvZhWJUdexdq+
b2j+YSA31TgCMEiZaWqEj9ayGowTHkMoJZiE8VyGtjcPVnTS6RxRt7PnXYbHHaUv+YtNIuacP50Q
m78RQSFVtsOp1GObYyLxY1YpgAGgtHrp0+xLozUzLMY0VGpNaPQLpyPyj2DYIcaVw6u8WrrZmtjz
XhMTC1xp09RBc7GhnYc25VIR0ThncSO5pKVa8MYq440o81E0oSEWC99BH6IB4Gw87Cm36gfNScVB
sgfnAb0fKo8riuQBuRr8wGoAUu9BKvtxiLI12ej4sGYQ7Y4SHrujNLopnw/jIjN3jlVc4+jeBfI2
XP/MvRLhg3HQGt+7dEhUSFPvBaZptwjTbvMK7IHKDXiCWzX5AdqMUikHjdUfM8F7cyZIf9KBJX5q
6fO7kVi3qrBaoICOAjkJJDZRYFSuTLq5TyIhvO++4kaxN/me4ThGoXBS8ttk+TisT9sZIEihvu8T
eDjYQr5cGUritWEAq/mAJQS14KP6hWr3cg2+W5Qw/mE5cPyht7p588UOfpF+5XeEkIgyLrBKuk1K
44OQBWgpcJUVb+MLXBGBr3OY6Zi4H1yYpQsoB4hR+MzKsfHPf+zdC+7jKFjjSY0WmG55jzNupyr/
E5GdKTBkpi6QGJTeFTLyjjUYTuGM/fwl8/bvCH8oYs4dDO9SuZ5SGtY6o82c0st0NIkkScbf6wdx
CASQww4qIPoxqi/CwrzHUYlC+TU8znIUA2KjbToBz97NzdNJUo017zlhoN4nK5a3J45KrHMBGn9f
Agvx6zDx/l7HR6z3pzhx8gc8N3EKvYJL8GLSJ8v8jSqoukVYOF4WsgJVuYygMrCu7CKOZV+YpHuu
3BME4PNMqeCd7WpoAOIxHDnfpNHqCIh38dYJNFBxehuJVCgO5dgPqHAJkex0ylHotD89B2wZ5mzb
2JF1j4fJXh/KXFFHlHOrzDBaWeHJZH6+vhBQRxc9/QQiq8cuUP3hx+Kz2wGyKWChXW2/Om1gyAOy
JfP3TJEhc5EBZQXKY0myZfVSkh1LBjv1YpopgzlU1WLYfkAUNaeyNxNWzKwg1et5jO3mLUJD3gAH
kP7niXiyT75JbAwAehjWSvZIxr9UQ/VUnxOI6NqJh27WFJNY3ApGBpNOuX+TYi60KHtfNuCBZlE5
YL87qaR45bzKcyWdBd7RRO4Ne+83qLZ6Oc7MCzoVifB4paBxbjbnyVeAO4dZu5XonjXiMd6XGQT4
Y2g0yhNbVXSuZgfUJHzxkosPoLlpgZforHdDyEZ1cgKhZ7J5mbYfnWW+wlLPzRomgPVzxGWeJ/9j
Lmn6dVEV0B8NIMXKIp9ia/OzzSD65xCdHlpQKTdbdIt3cjbOh55YhEBHNuzxd10kCikzGwH9zZS5
lYscTGbdF3Bbc+C2tcdt8zOAuNfech96l3BdZZIzljVVdm+a7oinagsM3+XO27tnoHmIfsbqVlAB
3RQ5K4YpAKnSJa/a7J92GfW9yrOQmS72C3oDv9oTSRP0hkxfXqTm3LW7gw3gaKM+TP5DMkPWJnO5
5ViAqhJKQFl7Vf4ZJvnwlJLmFLqTtykozwQttBxtiFTVkOPw6MR4EPMoG/oBHHOtMOZm5vlQeaqS
VjyFR8IiV6GqoQhX5VyKDFqnUBtE5fGyz8bgh+95qc0F2B2b9U3bnXL+b3FvCNvyOfPQKL0J4Hvw
ua6o2wfVg89HdXzZzE1ABfZ9Q+wNoGWoYobiYgVb77mMlvH3J5LL9eMzWWGBNFNG3cFnXeZnpL8/
4kyNshLtYbIr2wln+nN7Zr98gziY7+MnwUR1bFaoxm7Ut32HkmR9jkS5VaKVEGeKCHZ9ZE3dd71F
m/b7G6/LGenFJ9CWKdIFv8cGm0HpzGymMDiOoPAT8SvwIjyzpY414ALDpGMcseC0qD83pG2ZWAXF
ugaW3cCKs5MCyJkp8pk3g4rVIKPMqhm/VEQ9LIzhU4REAujCfLiCpsaNyydQBTESzw3fso0lDswI
DCFlgENf2PukgyALomA7oelSaJFsyxAyxhaVbmXIFUHS259GhKsbweqiBAu/eab46T4G1QtcJ5aY
Qim1VZPj7tZQW11sNVFtkyRq6Vs/bkKmKiHAYn13nnIykwuKIPz2STkvst+LFZlbV/hzSguuSb5M
3+WzGF9eJDONqQrC1pfoh4VDivKI+YkUs6K/eIIxLTBtRdlyr1NAcyDIXHfN46A2QfbKqP91SJzy
Sy067QUltIs9PH6GlvetUNS9XY3IHz5aX41EttEVyjhYrIpi2SgefAY+BGiK7Asr/BrXipdfm09U
kza65Ma880oJNslYgWk/0PkclwkpYTC/gbsWW+xF6CUV1T5uiYTDm2jePVXRUd9uItFTk+tGM4oX
B+VHBoodqYBPOWZIG+X8lG5ia6ajpKDnigRVSNzdJcs/NmuTlv8MjoTDO77cRH6VxfvdS9vSOh6z
eU75NKb9527d8ZVpj+VWI+/UZYhxco0iJTbK6/i2cMZ9N9wzAp2A5Wfezwab9DvD02k2lt89o179
VhUms851yJY2GtEn6HV4t9BfIjV17Eg0C1qNutIcqx8lVpNF9tMuIM2swVZIYFe50whAoEjtiiqd
ziw9sMUBNoZ/vYOEeru5hZ9/XBW1mPKSS1TQ0zHLAZUdaOusiE5t92Kt66+OEw23mH3qKmI1OMJB
sa5KSMcOqruau+1khKWDrnFTdX4VPBlk4oBKUd0J2IHak2EAf85EYtJL5YfyipTMiPifhbCCAjfr
t9mv9qUOx4TeGPbwyqvt6mBpLNyOgYgPNhV6og8DVzuMM6W0VF/pNvKGbT/E4Sfu/ggFw64GYmJD
LKRmNw+Afhb9CbKkgSQICwkXpuUTkDBmQ/eo9maAKGqb+UXmFqryMG38vhowq5knUxfr7Fudm3jZ
Kjl3a5WIAstxs6DkBCBVi+3OSSKV+I07a26/Y4aCNFuLsukCY0orJQRXosrA2iqv9xawXYYrJYfv
7okukaQ/VNXaCqVLVH3RI3IQJiBbTYcD7YNBgXJoUWK0UMeyp+I0+VPQ1ZhAI4sR9EaLr2WyEK2D
D55OAUhSWtSmCxxm48/O+KkHqrGOjZrFfqul4EusHPmpfOrUIwXN8HOVbG2zR91cwEh57M8gdCK/
ayvf6e1HtrqgYKPZ6ONDsPq+o+CiKAT89d+btbBY2nebmzcV0/kwt3srDzlr8PujseuW1x8C6Sc6
o3k+Ab/stHj6Zck9lXZtgZjOZKbnBYHvlj5LWhjQn1+m0E0ykIJKeThaXlZ+8gWys0b5i0CIY0gr
yl/WBHVIiINmHC22frUBzoR8/ZSDSezscucrdOI0zIsTp4hrSKfYxlMC16U7N/3mU18DXVshIGHM
ugl9g25JIGbiieqGHIQLLSgmf039qPg2xScXSRcNN9HG1b84b9EuWxpCJvyBPojH+hInRJVyZjPH
7yXY1t0c71F65HCOjhSnKr7vEz6/bmYkjRglauNN6lveLRz7cAeWVa89NN9ENv3bCbOxMhUiriY8
krI/T86TDpV6+n4Qb+biKYpqEubJX7d1ogy0J9x1LrJirHcA3Wb9FNg7hioM9DdxxDFRxikSViX/
+0gHI66xGIn9bgK6ql3QSlaelY8MIYyHJSq+gVsCkF5l6IiyCvCHZ5Yhrv/xjBVJccNbp/JrWnc+
F1FJI4wsnupGxoeQdOZzz76cgAoHyMk1SqlYAA6a1zaLeLdYL2ZxIrDgudpXssnKEg9O6kwp1SIR
Gzwxtsp04KgOdSTAABEiPwZmsM+en6uVy6bW6/MEmRkFuRbpl4Yu18pX/zd1vZhWmzMjh1iUdXIr
x1oSTvqKxs9ICf903mklTlWSvFmRmQEGomxGK2s0+qgXmMU5NZHyypyfwl/d9QyHUHXjEFSitMUG
gSWX3a2u37UChvLMZrKh0DTKOZqXYG95x1YpMroCO3DDJCdac/5j/SR6sxsDGmaHfdz2TlIrgK6i
XiW8oGSMzkewA49TYw/7FyTK8S+fFQaSpwlzlEMiRfXvsftpzimQm5QEuRwkBl8hNvWXugfSUDcG
qDGA8WF2GzqgYZtMDNYV6VMAAAyP68mSFdCYeozj9DRFx3+8w9ZeceNj7IV2n7+NjOk90whWNNSQ
b4EYCCtpxzvAtvCKxpQzs/S5WijdgyZeWvAN4JNvmKhQAnzDjJQOkeeXHtI0GZvOS3OeXhC96SIM
Wz0qFNCVRMjZO5WOjeKW8c9fQjl5z4S4ADPdzUELBMtjgVH5a2fTFeL7jFhZBKalsxVLHSGsSZ7Z
5/xPWjC05/vizz0kg1q5kDIwiKfbyUYVRUyYyB/puzIDJv6/jH8FRdyx5S2nTgJw6A+A+xeFqZnL
J0X/G3yT4oUv6TMLyHRZfW5F7C7aruB0YJFQZOvErTCnu8gdkbNsOi/2G5txfAp3WueJMXY5pCzL
/qh+tvZMX+pBE7j/3K2Qb3djbFaVPfoKufMq98o2qqIMnvC1AyV8y44oiRET+P0nEKXoqjakjNcn
D+Wi4ZQOm970S4nj2sQBmZG/KntOiidAsgT1fBWYLTnLIP2rg/ilX5EqF+HhOR0fPTS8SAG5Yef4
rhJnM0Ac5PBD8M3mLJV9haS+J4/nuTZ3srMAgwYmRZS+AJcf0CgXmJ2LZOj4jDIPbj6FIpgA3B+T
y9qjs7j1Fr+eEGDLQSr/LMKV5Y3auPnE1HZTxp0UsfXeSLuHd8dAZHSRW1liZ8v4/2gLnqfdbIBe
qJdbEzs47YlnSz2s2UMLVQrijLARACrxSTHQeHlWeKNOuWU4lLoiWQSJh5IgwWKADfv1k8U/176e
y2z8nDtSp7/k+nk5vTcBsi65a1CkQeCzDMZb0lKzCJOKR0ZmAGcVOJjdFdk2XAxQ/a+LCwIvGnya
is+dv4TRTfHVqPWoN+KbqK6PeXCPfEkaV0+jqBU+rpx4KkhunQzExA1H4xXGI5SBTx7Z6Ilpz+z0
qFEDqg27ohxMQCN7jCg/SzoM7jf7oeebeAMwkiHdP0XkLX7CBTIVv+ToCo7LaPJoHHSe7O4/ltei
nZMcpE3tn785IcPgP9j/uJ95s1A89l6LCV1doYjtiSMhVFmKWdqX49vVCEygova8mx0QuJx0c5m9
qIP/VOEgegqvg0+u2fLDebpdqStscNkvOOgMLeSN4gwgO3Q+Fs7dXBz5ELmL3KkdKejt2FcHTF05
TgC5j8Baa0TNkhSBs4/MDf0Wt5YjqNxP53xHfh3j2WphoWMqagfvie08StkgwYjiYv6nKJdALsFD
Lrq4SctnJ5Q6fow5nNCuurk4VzSZplBjKf/AWfdqbQdV9vQz5j2Qt4WjGw0UHxLzQx8hm55LSFED
XAjxzVuBis4OB2Su1CQaF5WMCwLbpXv9pM/fVUrDoIB3uoBRyKCYluzvkvS2dBC8z80im9FIZBCw
rOy4jtAT2fD3YHHHtE+2qa1k0peR4gjiyBlkCOdyzr7gdRX8y1/odaWyx5M09jLCvltQvTEz3vNQ
XsnD5l7oKa4ztY5NcXJvrAVEwX4iwyKvb+Y6CcfNJaxfzMsc7BSpvlg8kCDyiEmyAWYfARjtlH0X
n95J6UnikD7RmVTYqpASrEXY8fWf8H3Oa6Af9mXHH39PVc1iHx+YTK+x4rGflmD+IuFiazfmZCBw
jy143Raa9AZ5bX4BPQXZ+bEOz7vKkoYjKqRyaA1bodXVLlq0I34rw9ZlnOLJb2/qS1GfiOQCXjNf
3X/tTgjz2EUhGhIc2qP5DSqPqVoQOH7464952uF7ftrQ3C2iRZ3DPk9XTHPkYZMdJcufhy8cEadf
zvBOE2EzjOYlHcxqWjv6Ce7HMN4B6XXcqSmDp5tTkQBK8Fr8xtBWHTheAGrlob98vKQJmSild39p
LRa7Gi8tP3D+BmbBe6D4wQtqN89rysk0f5t/NgsQ3moYPGpxwYapA2ljJVgYXqGwZUZNv3FGXRF9
EE0Y7w2JiR3mRh35nwqzScxjmX1V9NPatsb9tVWvdAkiEl8qk2A5mVYFcfhp5Xsd12dNDkJMOihv
MgFFM5RQ5xIX1rMxMwXCqIqr+/kZvKR0GT7zgNxcB/OUdjQoZWNfz/VUVp1f7n0nbwuIyCyV7jkB
KJ+9UDUwr/FkD7iQJ0bRRz+EYG4FQnYu3EoZIexcqEwN1mEkGXj7OrnEV/xjmpCSlXsqfDe8ZKzI
Ni3RGtSRbjZ/Ed91qehiR7lDMHrJuFfDwxfTlAKSMhgkR9YxtlilIKBldFKy1XbDOrdn9rogmB7B
5O0/qAId57oiDonoy4kQfRJJGMvxdi/q5rJJHC697oEpH1FqS2K/pG95+sfLIlf7vjVJJupqsDsB
5aSyA8zFGuh2CiVBB9Q881p+n5upBe4faA2DHZW6ozWod2Bb0iNdzyFUTIKdyjhO5mmRtvhZCBeW
pmI2uhg4mvvhO4h5+y0nfCSShqUkTCdji7Aa1/homhB58HE9hWkMx685EaQtm7MlRAuxjajZYYSX
KgW/eEqRqu0E4HKtaSkRNMCbkzY8d5TK96GudhrMa+wzB6vDrCBgJsvVjGPGniKYfCp6Sl4rtbfK
B+K8PBKZ+cRifMAMMJ62QTtFnYhGF78UkugBsu/gF/ngAn7bVD76WsT6baarEmqKTKwtXZOQ7tSg
8zbtTrR3EYkdwMm9r343MAWg4tX8FdklQKxoVqlUJvNmwE2lool/+E+DhJNI66092WbOFeik2YDG
njHZDGXHAKltyhfT8Yr9wiD5NseYDpQKs6FEQFGyDFLq2dRMfmA1KwwkJPxi6KbLVz7q3Xa5cyNX
6q62SLiWR4nfFNyVR1nBDUMtviryrr8y7BS9fVVtaT63TsBQKewYpzG1F1kVBhmT56+DwsyMIMVG
OhVhuNwej/T5iJdx7c5Jw02z/wbb8A79cPnHA3xbE+gsnrcdjaKA34buiHjlCStWnGq8STb5FDtb
UYYQL2ZM+bGZVuZSl63Di/NCQj953eldsuaf+yDiesaFq6XM1VX1ME1eD2DdazETDRManHxAGLh3
X0nAxhORXLeaAqI3ZwhawHzOMQrxMNd+66whJZRq6ijIZtyV/ZR9iBBGuMQCJVt4iqEaSalzUr6K
21Zd4SW1TAGj2UMioF5Xy2Nqh1xQSZUuaQmK6tTYosKJo6xKHis1JELCRmKGiQlOVfuxDrD240Lp
TsVN5dB9hLVgKX7Mk6eq2mDmoIpHqXmdCCUYv9D5yoaYzI0PBzdTqBveStlPlZjpr44D0y8l7Vee
b25u/2i4TWhWY+3Dx7//Jkqz6EJ8pA5jtnK2SIB9kqZU4j2lHVMhPt8S+RjeF4tTQjZ7vl6nEY+f
EPdePSYKGOkmwJ/VMIlSJL462yWtlhx7JuI616iA3/4GiGfkXYb0edka5RLT+dZ8SfsyUBcHKREm
HAaPggJFF7hs6JFZG781WC2kcEuYJEEhx4R+cJk8ensWC7LkXJgIX6XpleZlbMxO1RojEL5QwzL7
it5ZZcixceEPE5cOq0eJ9YrwTr+rg5o/P6pTNLBzJe6q1y2LA1tIdbDnKLLVM4n6GRTW0mVU0PyJ
2G5ULoariOlm6fbDsmxMma6Hwj4/GhR9bjW2NDURVFenxFA7p8jI6RLCQ7ahYA05kliwoz3STqSa
bS0DSsqMVc3Ck6Yho+fQyksHLYYh33FLZn6vkP2HKspPCMVH1lfdKe133vf0s2fum8jqYqAm9VyB
H+baeCQDdrrRDVy6QKD9rvfbMt6mTzt8m1alqf3t5pRRKnXQQrKaICEDpE9+1aqXtyLoZXxBk7rp
1nvwpGn+R7rVJrLESdN31AIvov2j7rT7DiKJ1NsiMTY9l9TtUfpS/iqi1Si9swdywJjHzXh9SZY5
1iI9BJA6mpwub+QLgWfeUPwy+t7V3qO/ccqak9uGX+OYubVjbeVeq36VfKELc2MhndKJt06D8BmX
yTg+JCWyYxfrZfyQ/6JN7uCth/SEuFpXl9JhEXvWU0IVXKmxiTR163Nyj0GXyVS8EVhMJvNT6sSv
OORylrasiULx8A31PjZUSHp2Yr6orsLzocwPSSAMFO3sK5JqBOCCCCBeH1UgIXgch/IhJwzfdizr
gIfL+3rOpJj5p5wHxbd3rXGrpAEytK8imgIK9Rs3jl3eEoMiR/yGKtlIQ26ieB5Njscri49xBioR
DiE2RR8z6MWCYhDU+eBwIhypL357kouf5vbcB2PztoRsskP0mB24qAS0gJe9y8ajiwQfPozOXu/M
ZG+b9allj57qKkEVxa/VdecDlrjKWRvhimO4VUiLbyQXgHNR21fPSmGbRPlV3jbrUAS2Rc5dcaYx
N4h5yyWnBJ+3vZu+gNEljYWhoV8J8NBwKsnHnvy9OqY/sxqdrWPtG+5q1nyLFYctLTrpyrGbVt06
hGCDklWfm5jimgbdTPES3l78dx7d+vyHh3Y3dhFAQhE6QOIohrmT59lSEuX3nWNuM7XHzeonECix
kVConsWydqLnoWfYlCGVjmqylsYT4g+CIyCNjtcua5lODi3BdSCAKKRV/yofhqr6FnQS/lTju2Du
hp5WQzrR1getYBnHtpArvDl36c50jw5Pnd0E3C1rh4BZenNzNVRRoKsT9TNplTek03pniN6KQ27n
Fxf4DT/+ZxzDu/blB8pLMr9Rqo0GGmRSV0VGCMb8P4dgAyuxFCdCLLUNb8yp6/KzBuWITS/xvaJY
6VlxKzbHTiCYe4Mn+2ZVTKSUBX/EtqyDUgBRFsixQW7HDd1p/V41xcEz/JplM81Qri87jUEH4tma
8qOi7504ZEXMb5UpjBNaSEJwTE8tISKAsYBKpYzqqvzLd1LgYkInwgLmjvpqZwaYlaulSlb63kqS
RbbdBfds+Il05Mn3TgnulQpp6/YBOaHnATVdE+7s/WoNexIL4M2N0rzB6HCD8JRAmCjBXamMRBA0
7mhGBfU1oo44cnXlDdthIz2C9WEq+7V/i7i2tId+PS3NPgIhl3G/02HZl8mLrcMwhtBHVqomSjaY
IyjoIk935Py48kw06fPWaCHz8hbm5JAxRBRloT+q7S6PGCuQUYvBoISqEGZkgvvc0Iq+ntOSGaz6
XlXK5nNZQeWgpI9AltpB9di6Q08bsa/h83FBm6sIQKAzd2PhV0Z09V/yF5XVQVmuN6j++Itn5w3b
bkgiQ8fbUz9qT3GMX5c6AluxRhUEIt5RWEQotXnnUYBcjOLdFCBARhQbnMMlvmc7MPTU1n5//aFC
jSeIIJ0AlHEY0cjOhLMJ+01j+FTlHhqgZk9jnL+Ao/gGSHwWexzTo+QxyQsrfJrGhhIBxIeSCABK
apNPnYep+RIO41wufSF4MI7sGLvr5B+4r6nXTa1FI/vp0c4e0EdNrzF/vJI6MrLFJ3/+fvQTFhzb
WgmtjsTcjyGkvb+69GW1Ufta+Jv392FYAN9cEDi8OJ/IfJgWusWPYWwvreicbcP/DuwZ1kZv9XqY
due9Vknb4yOnOZQkGuXEnd4L++OkxQibdbKDwRI9qPIDWg+65QA2ksZJcYchgoqFj7Ga+RXSQbUC
ikxg8/SFXvZXGUn35fBK1p5CdN9bfWf33FHJnAumNGwApzx4KOodDrDpSv4yqbptbNlVBlfkqZ0Z
8M3r4qo3oQ+n93jLMpUThxgzcPEZBriAQgCA1GZQIhF85yjzwDszmAWZnB60I3qTiodDe6E9MqIr
ARmUzepOHmoRKmFvsFLSGqJ0c4jyMC83A63pldblcUSR5JLNhJ4XIcpgMWF2VugDkjbM6+Apblyp
V3465yGVrbMZ0rHulUDD4MSitZxf/W8qi0C2vIllDZd0erjGFNNJ6P0jMycAb5B7jkV18IXsqjKB
jo8el53N2lhC0COkh1ZaC2PWtDW0vwuH36kZifkfinsACAIK0xNospc2Ja9gJiyAUUFa0qMX5TwL
zqniGJJUVbnwv7LmeRC7LStF8x7xl47+JC+jAFHipHnSJ7vEejJ7UXRa6x5ZNcISyPCtmlaSok4j
WilKXXb7P3z/nuGKVlz9iEBiTk6zpfecW+cezC+9eeBVXzOy3eGMKTR8qnWdkPvNJxAujUIIarPT
44rXcKBkSECa2iggPYuY8TMpXwPro0e4iMespYzma3jLKnV/oQnbruvoK7++hl2ZscuHpDExTmaC
VCEhwRFPpulfnLGvDyGAx3Mj0Z3zr6VH83wqcUuAlzfBejgYzOxJ962KUQULYy/cQKmSIhoyExQP
f0IF3h0kVdxMuFqvO6uu7e3TRx+dOrJRL4Bf60kzcVpPHSL6ySXOuUmV8FPMyGb5Z4OpdDmoGoG0
8nrkaAhwyQvegeYUDKLZuRAcemQIbrkSMSFCCpSTa7TtxUObP2o7oNOjjoIHWh6EMRuIuJFLz+O0
cseiNWh8rhw4cdxPjqPe6++O9RySwpsEI6HVshvJUnFnR9A3cyA9oL7w0GK7zwnNrLjer6J0h5sm
s5JvfbGQm43+jg9hyN6bD1cl2rcDpybt9uFmIujTwlMG+mO1EWQi/jqKzKriBWexkEB7yJ/mu8vi
SyauQQmc9s9lpkbxA6YpVQdmlMoXweVkKpVKlDv8sRewZ57/iAtkXduuaqbBW4qinPkjvp0Z8Lim
OQBNRCEN31ddnnGPnS0RSNEHJ2whqPC+60Z5tyeWrnC9paZqcus+18hFC4bAh5/IScto0Skvn+E/
bevidFJ3KVlTtu3M4fWeeE7S3f19Pt1RMuqbWBFSRQR5KLlkLqH34xYQhqMrJjGPIMCbAlWdEaCJ
mxK0O7r+e7vjGSIicH+hNgTPu49XJUBl9Lncoqbp9wxgFqV1TsJQzR/R6omo+AwoECeYxsg+crTt
+/8v6Dq+N/GeQHTSGol5lGE6ZNCRsIQhTv7GMLA5Bp/3LxmZ6JJXNdvi+/AvMujjAWOb4PEhZAV5
y0XssWRzCuxFYU7hXF49+C3uxjpad9XiLSZLI2dJyJ+7meo5BQftptjA3JYULzpxFuv/kATQCvNv
EoPro6NXmJCcIRO+Chjv7ZydH4LRKOroTIySVxEJhDpYYB19M5lFvBfhLFMG9fQqXsCbLfBkrrZt
PdDqgJpt0t0ifGGo4SVlyWg/4ojw1T4kVXoXLyxHFKi2qMmE0XNApdeaQ3Q8Il8n+EQbTYCM40XM
N2LVR3OOpiwlJsQ2S01udS/L/mdCW/yjjzQcGhR7D8H1BbCuBBDRCKfN58wkQ2QBzApb2LHI3YtL
WuxbYCmn7PZddS2GnGGxQgmLwAiJ//hdoRMOXZmurjy5KBn0WAo/VSmHy1wqtJwnvi0GZ4Zk+91M
uD5j6WiZN8mk+/7IVP9sZtFaTkcCPzkZX3Qoh51FEp6j/6NNmdpk5ij9jc/aZGjwLTCSz1wJnfDk
bzdXdTmGBko9tMuA4latXXl3jpUrjEJfAWsXbuLTQXt7diZGea3ib+mw7tcaif3XgQ4aNO07+/av
09Lbei9A+x0PxAH7TvALMUDvULqQLLxTVj7SydvpFDLQcTefDUlxU3Q/o12cmv4CVLaO+jnHa3Cp
LvTK/00QPa5D1kfZ6/+6DkqZhXztARGJy+MiPIz20AWEQ0l7spVES2hapSaitREGvPPgZM6KSM9o
PxR76L/L0Sd5ZN+mcRoKikDLA4MZvr/fqbdZQBFGI98RweTOWKr+ArSZ+MPXAodhAnzLFObvcY8z
OzL6vRD2kVXio6A9B0ycd+TWHyRBCRG2Tz9RfO+hS8NzvepdkSXNQwHLTANCWadko4gzzVQr7Rc7
t0OxUQurZ2e+QkvHTv18S/fqfWwv3x3YdL/vWPoUqZtacPlYkmy1dDRV7CEctCailiWK/02WEfOd
TI6dz3o2YFYhPYHd20lcJHrqX0spIuKFOc/yESPnBawEthJBwAglHQeSB5LKXl96gs66NFEoNgZd
Vays2zOqjTn33tmcGlkzcQfuUhA1ziLU/pHHdqQnD8/+ONAM43Hb/v8c8xAvXHZSvkyq+g7z1j0t
WxwmJbJTswFApGs6uBwoUxch6xpvlYfGtbYPL0IjL9ZaVqZF6M/IKDmZOq1c3DvIHzLqQc51ZcgJ
WPY+3B7f823Rb7HUNSyywcOdhefZYpEbkBgdYbWRKjG4jbh6QbH6Cula/GoAxADdd9y0XVESUZix
VdPuX4zTn7mkAffvcrfnE15xvbmi3bLj0jzbrG2TneNy0NhU339gJfT54+1eoEeGtyRHQSBgQEor
t1XDDVGHiSjHFzKno8vBgpEhSJaZ1JfRY5vxCCl19oGHLT3BrzM5fD81Lq+wNuUDV9ZATiGjpJXV
n5uidQhNvzvaPuzUFZrm0D1fOPnWImlYZUlUNFUzN5Z8eExBXWj2659wKUcGYYA+gcam/9jqPt6q
0ZN9lnwddQNfWvplTgZxTC/5vNUqJoTnzFZTW+NLR3PFt4KQcmP+sUwIX57o1IygcRCAnvPV0uL/
y7efNIy8kI1hRY0Gkn4GwbEuLpqXaCFr1LnRstZ6sv4kws7+HvnZLTqgS71GVzv6nraLQjo1stSE
neu0ySrd8G5BWG4rdQanPR9yl4e1oJCyO+JmXAHZTrcNAbQYYR40WHRCmUXUmIcbUEjNYfTXEtMm
O3NZKDZnFTIXrPzELD7jJ4ZCI48ZdA6QwaPAF43fThc4TgC/x2s5fTTJseWWLCxln7KS2pEcq4jl
2KZcNP8fq01ARv21CobDgmxKrplu7+ZcvR/ahmYs/qefVAWOG9JGejjJ6iYkv2eJCHM1P3zKvwZV
DoixAU813x76ElT5H6SVWaRHwY5pW2OHncIABh80gAbV39todqw5N3u6phiyIr/VAJMAz90lLd/1
rLrlaFTEqvDLAP7Loxh62k/gL3f3zDcR5FvS0B1V64PSPwX7UXBZ2GFtW/ro+3Qqe6/AydXGHOSd
pesB198bOtqe7zC3gVzwt9jyNS9jjoAHGe960mvd8hlA0CNE0hwBcDN5s6PGTX9K4YgXcC8EdOaL
s1wUqJAcT0XI/emgMN2oTKPskhWLHyk95ETl+z9aEkbFAoVgi0jB3wGLgEynDgQnsW4M1wMPpum9
u1R0bG8fr+poJXxTv/TFZ+gJAb0ROaBJQjytz3G2cclcZ2+tuVb6zV7M6PlQ6AGJVjscUhphkBui
BL8Sboe9qfqSmkz9iJg4I3vm/4BlNEuViEezkecxqoQwagfRU9FrW3t/JmMm0gXes9QJE6oi0WJI
ukOKxTZhoThQXZbNytLUmhuzN3IrVXYXpmsJ/HQgXD4Pp/DWC13ihcY7nRX8BpGAKwRaQ9yYReO0
EA1REcVGdTzGkhR9FJrZhwPYlKuBz1CwO5PH0Vqn3o9QqYdPeqXHG/RhHk0Z73N1p7admo4u3Gwz
nRyKE+NxJGGqJwartdz7pYzK5R85gZBES5f5dlskCrOpfSdK0vOtMoS3TL3E5iXn7dLZsbz9rjWr
TCBsb9xWyvWaBlsNZYbWrIfzS9Os6TdmiAE93+jB13NUuqXDDPv9QgMZTWG9xl3/TJMgUFXfChMZ
C6AEuEAKrFaMDLEb5slENCjQkjTL47RJ+Spn4iZG/bczDqFk1amqb51CdQF5OzmKY3iCbx8vUWM9
wGIlfOpjAYJQY1IkbRmMWi7R6y0U0WrV1T+ESpwx5hORRqTIrNMeStS8QsMh8RkSEMT/5jCKOTDB
JdEjqac9ZuRs0B9TCDc75oFN6Z8P7jrVQFDu6alHhORXt2NmeaaYALIUzu2rYwfJc+mhtdFyXEMk
o3QoKZAq0RMFx/MHjrr0fQHneagkAdDtbA7mURPwHvnsi/eaxzRh9Ro0H4RaQi0FsNiSm7S8bQ0k
ttVMAkhlCZV4wMTWUe80I8ICVhM40I9pe5TseWRynNNs8M77Om0t0SiO0ChyNiv9nfY3CrxPAmXc
6lWXgdlzkkAXfWejplPISHYg0nzHK8ERSICbY7vv7LU/Pw/+/XsF4ar9sq12DHVLOEacRzCGh67N
HpqC3dh0MQGvYsGsVcPwjsQtbTLqf9otPGShh29M0S/A6fpQszASH4kYs5FZnIGeVnDJkxvzjlFO
fHu/UdHWQ8qk2vwFcnEOMtbhCCjeR279hwZoEHKvXzEHaryOE2hW+DCy+ai17W44LZHJjaEwLpiJ
0z7pF+Rn31zak2pomdTrrp0BX2bOTwzcRprhMMdFCtznNvSgnEqRCiJQDci0bpyJ3+kbeaO8Gak4
rmQX/HNEAg5EDytKHKYz1pHK9BNaBLbmJ2rR3D0kctirIeARg7FbKy+MCaoOf7junhHTK8kTNVT1
eJ0H57L5n/MrVP9lL6dDOqAxQrH2nY0U2BrfEoH+eV013wVZPJ/TayJWrQhrQ1WdAxEfTkTj6KS7
Y2D10zeCwucYMg4Bz6fC44UFQ6sXdj2axm8wd22shKuqGzXaRlf40/Xej0vhzKlGrmOobFt4WuBQ
hjJIe/Y18dxb/X6kHVvdayR36iDUFGRMDHtuS7w8Alc4kKe1LRhF3KwD3jobw1E+B5YYyguRpi1a
1P7I3MF2HNcLeGJcRtohljQ+bkF6bKKDN9GAl6RdhHOV8DiTz60HIr05TJBfgr5HJy3O90Oomj0p
d26uc9DtzV9qRphv55lCLKKhyKdX8oEJkSytSnV01IjdJRqaKF5ASf1q0X4SpThMfSHegPCe0aTm
ZbTSljbYv/YE/UrkigRyGKSQ4QshyWU/Q1ZERZpIm+HUjpC2Mc5lFAVkcclCmzFZduW2qizoJE39
/GIIA6FCDwcZrvcOtJJdOZvP6iuEaH+fUHHxE/7u0UDHRvUiXShGQNmU43QI9MSGocVeOWs/079u
saZJN8n7LsTVWJK5O61hFEJ79Gua7O1ENadfYFqqxrK8prk95QhBTnr5BFfs8C9SgYqhRAhmydUs
TtH2ggS20eWPtWDkr456zhgsFfZN2GqoHkPE7RzurY9tUipT68hzDGpaYo/RnXktqlEIYsdjX7eq
R7IL9AkOmL+tTTNGLmy5EDn1aGJ+iKUlZMPTQn8PN5KnPaqXJgyB0zD4e43JELdwx5LpomRbnCvo
SSwRIpQvhwQzliY1F7I06zidDVkrLeTMO+e2LkD9odtLGWAJAbmwGwXbSt/xSb2ONPOZMFMyBFjt
VebrNpDWwhOfG4AM2TUeJfkvFkulSEI1sCzgKeSZ2FqoQb4YSBkep35/IE9ZjCPdWwLrNKEjzjex
6zJWA2cQOXgplLQlBrAFVVBjNY7jUDnYhkmZPy+vdsDqVNo/YHwKgaNioz2iq/n9drvP9/kcqCL4
r5GCU1hq4mNU6NxhwDnORttXmp3GpTYjqa13yjtMowqFNHH5aGxubjDu14mk0bMShMKWcYLcMefz
VrRal3X8m6EeHTkgLkQ9YtYokqHKNRvmstZk2rRW36Gt2q5HZ388nOZq5lJ3MtwVfBUmCODZruoK
hhmxZqFUG6X1pjMUithJDIa6ur5wBNGfUzkOt1HRmaN8QCwUKmh9nu0Qa3MEIIHGyp1EB/ZZVslK
XpOEe6rXap4C7HnAPX6tLcrK+E6as6YnavB+mzLcgOe9OfActBVew22YC4MjPazbmmEDzfptK+Lq
5RmulXvlMynjiWKN0UMXT0KLsnhMRwWl1ugXp8MNl16e5pWngAYswysN60rtw65+ANN+nfqDgjbc
mqcb1KXBYg4WIH1B4ab5OOnH7lg0qgwFuSPYj+YSDJs0LBsvIFvZ5r8XZAxNLf0smGkPiPPQXG/J
VjH9c4qGO3pstOeN5TZxzrDkYvoSyF3tOTBkHv5tqSRf1ckYNHkJJsKLXGpyDhkUdzGErduwrN+u
61LFWjmgrM/L98Kbd+DNkMUr3i3yYTvFobSLUm2KcRv3iSzqfpdD0zFlqgVhMmW/3cdVkcHtUoAp
ktcp5RFQvpclzqxFh0iP5aDkSwgMDoZKR0qBg+P1MUjy4Tl5JHZFYI0cnoBLNfjYNa4xdjtjnQ1Z
OnpzVUQGiESWDn75qictrYuAZba0TgIGsTi/YK+lkghGYeG1+7HtMOn9+GUNho7pbDRB+ZX7dhUD
AcCcKL15C7mzoVVjUPI3aOeXeiYpIlYDRPSMdq2DtL1fIE4w2mrKI044uXljemZ+lkYDxm6MekNA
W4AUInORinvmpQWjncdweParv0ykmmPR9wGYccoFMWioJs6jAIxBylnlVnV1ahcMwIlmCCihQVh1
vzAWVx2rV/bDYdcG2/nwqHSHInW/+HrI5QMaWdQFvIizqbDk0tedOXhQg0u3WgCxG2uQVsZ3gHbH
XceAp9WFv2t7rBBWjO7iZZZSIS4EsH2NgxU7WyTZuwxUsr0O46xCkGK8WKMYXT7L6137Rz8lzHtJ
flr12y3W/y0sSGaywFu9XC0jCMmKg4CWRGB0b+VdHLYBOV2XHNQmrf4Zx6tVk0BYnYSJU/K5S0qQ
CpWWH9VRKKZE6f6ERRKHYzHbcTnR/eAc3wzeZ++CkuprVAQsfnfeJYdWmsWQHUAbXc3ehF7Va0rM
BUG2trxMK6DDDpe45Yy9aQAkcx85Zr18xczsuTi2ltOIzAm81Z+4mfA2udQfa8L7zqaQdy9yJ4Wt
0HyU95wxFuwpaxxzxw0I3YzRlbG06n5bCw6ez9B9ljZI1nzeBOddMAeCuiGZ3yZo8ORiVBsOOZ6+
9qa35DrAUYqKVuHhdGVhrFgouotnTUd2PMlKULvwDbBu/c05P4ky0WEJfmGo9dlTFjvXFn/fe/nn
xasTvuu5m4M/EzmJTpS+Gvuyb0HbBK+n1jKVXLw6d/qmssH/qJwuJiu2s74grUF0Xcta/kL3Qm2h
GJ88DUoEQlmWeVd0VVFWGkqOhHOuJpCVp1W2mjGVdZZv+YxTsCcWj4oVGSE6c6CsKJBbfhWjZmbL
CvJDTvYmin2pfpPfdYgSnlHPA4U9jGwrAK9l9RlCLOL6/HjiDOaJo5BCsQXgzipdmt5zdf9+EfFn
Ot/Is2mavEXT3t6V1bvnQLDjqr8l5QiFdqdbuaA8yCYiAIjDOyqPfyxcI/RpIaHJVeeun2YLCsiW
vhrt3lGM/QSDSDQION+1LDY8lifYqISGo1OwHzZV1shRHLs7gJKbCy/p9Ajo+SS6sEsXXbN++sAr
nwi+1/9VgIMlm/3PH6r1XVHS7XTt2G8A+zG7CeE9GmshjvHdH9VZEaBO9X3uy8+tSTy4eBuYQLLW
lXb5AiA3lth8nGfdxDY029TPAzTFIWaMuMmnrgXyEeggIWBDeEgY6xK6tFzcBqWTkQrHgmSZmo+D
1DtWLAGcf7X9FAkTfN4kyOwcezawn/XcGp8GraBh+nWxAUhQ770mvTcvQbR8UUYv2xC82H9GG6pR
OJZYzb2u5yeWHMnXDZuSoPn8gESH7t2BIIlqLQUGANR0RnE1eu09ezCvwsM1Hc6mee+YRUaMoy5c
kf6qxquKnjOHQIqWerpDBxr9hX01/QtNWh/XQ7IuFKzWN2NiY4/dl8PTYYtk+p//RvzvenTyX/Ya
oSRHuGtMtJlg/HsZfn7jKS+5cGa3WPh/tp70hVi8YSEHkZXHpKv6JrYAyXLRa6wX61nla1x0gao2
FDKV7CYQ9Wc2yW6Ap0keOxUBe9hK/yCxrcPI97RqM8y02umhZdeE10gHY0BYxH7boDlbYk15oOse
qACYCY9Sdh77s3TJm9AqiMfqx7uLow4lSEnrEx7wvix2JdUwc/YKemMlYzUT2G4FBo0DFbstyDAN
9nq+QitvVaGnVxaPtnXW5x7uHMhewWO4sG5MSJbHEM3MkQqPK8ixm19FKtDxiKegBQFMGpd99WXn
YLLZPKSpIlr79TSEBSs6ha4fwqTwlsaYx2YJRqpNTLYt8x+WJ1t0/wnq3YSM1pCoTUhiGntAYoml
FktjCg7alTnr+AL8T2e0cHyrAoeuLk/aVlLkNBL1MlygoFwyhSUq0Sfe1Ub4po3LVKE26GOVVMXr
ornwZFyQQ3sxuxmvXzkHqKVFvwVe/LZZLm/GaiBa7f9zBRUs+dsJHNNj6YaemHFCPiMxOeBk9cPH
Qtoav9yp5CfGMBYcY1IYC2eCOm+oqThpLOcBgNxF6AV67FHdvv+jZ7osFHT9kero+gxbGpPXRWVW
kOevT5Au5YDOg1tcW0h2oSeQtrmtUOB1/HnDF7N3VNcrWoJnRojl44AX7JtkyK8w1Of+c4ckpE8A
meBnsr/eJ91aCCjbh/Zo+QuZbtFHm/Bb+OY13Q/3HdBLHeeXd+CG+urCS/Qo2Gt38Ys/JMugIbHR
bAx77vLRhz/sKtuUIN+j1d1dkJOI0SP0ZTUMx4rFMF5iaoSp1FiAPF8N8BPLOmmPXYZ8C+gp4lwS
PteVawT/lZewIS98Ilz2fGs3XHsYqyK354TuAxGqU7RlJpI1f56oGDYgWuQlb466Z0awGKAFbRB5
EYinE96uFfFLwkEFGBVC2QQ/HOCLcSfsyYtnuHbCsJJaReMq8hwtSB11pKqUTw0qJEGXpaOil7Fn
LB6VU0fdQ32FCXRHY4WPpG3tfRPC58Yvw0OVrlZE25+2Y9R5lipGHrf0Fkp0sy6jNXgX8TwwAAbS
xuzs+X2wiVubkPf9eMLffSXRg7uCZyq1ji3VvaVGJJtTQNTqOrQ3rgiADLQElG4+OSQBQX43zpBR
RRUDmBMNhATiugZWL/CLQ6yHOhUs1fdeXBlCQYEwXnxvRIO/m4z8O1s+Cqh1IiIAWB/G4CJoemhr
tVVLL6fzwgrFV4rIjtz/Fo8RMleb79TmQOHleQexb5v1dQEt3IqTz2N/q0xU/xJBHpx5349CrLWS
fZYPbIVLgHtjeEmGkg9LWLhXsEGyvEh+j5v8+xTuCR4xsvdirkakB2CdFmA9wben4N+eniL9Ghos
RRDclVMN6yoGFjjoK0p6keY2GRhzREJIi8aRMO3d6Cc/xZiFlmqni5kaqlq3OCmdHbRwCtNXzQ8O
wSk5Ktdi7f1F/Jh5IJ2j2KuVzJdftUDJ+kN1u8dUPm5dpwSGW7odMclYuyFHcYVJvkzDm/QbAtjA
6ylVGUE+xzvbp1C2uF70YZQeeDCVPMtKhkiUCRJ1VQMr2J+TeBiDmyxrQ3WBD6mMBKTP3LMw24v1
+S1tHR4QxZNqWHXCYn4TfCC/zM66Ho1Y7wlbeaRtG1Ign47vgO6V4aClzPI2P/FdQh6+9CH6FavV
WKPvcS0VLzNxun/Zn1ns0zA5hcMJo90y1V+RRXUaeT4i4qPL0NC7DLCxhAsO0mvRG4hlAnJDoXE0
e+3q4as45bnvLkSjsKxWorbRpEIEQrFvh+hZZ6D8WK9ELwvfcvYm/huM3FFbn+e1XlA5fu/Md51k
Jq6IXQkj1Jf0zbsWcUkKtv2YBM3DGFBNesJ8Fb58CGItXwXLJCh7fP2mNKfCfEMUIf/AQUNApGoY
iK4WnlSwloL7xpAlJXtnsJB0FpuFkcbBH3L53Ln0uFPQuFvfPBnw76hXJAO7PT2SVdx9ZhkiJKA0
wICGC3ASccY9iD208c4FzuwQMctsRBvcprp2PwcjNsWKsNfpGXl6krLrBZVy/9hlUSO2yNyWA1yJ
kkMi/dNCsM8Ugtz58hrhaC5PV70hl4dTfnYBJOyBonsjpve3jqqZs7/OdEOARWZS+H0kmeDWOUs/
1EmSkrpLhuVHVgyf3jHNb5zTy3ti5ueIbbhd1wrnBqHff5NFiqzf46ILWOXvy2jp5mw/vC72TVIq
N/1KXdus7sgx/V0qboHqSpk9DOeHPHAI1rHA6eXRYeb+f771iGuzCTm6Tieqt7Z94qeyzHjrToMw
DfFF7hi/wIj5wvtRjoprvSY2F11iQaFClyZmZtTSuFKJLCuUfjjutaRJfHTsWN6C34poRn1/cQ99
pH3DhSvkc+G0Dopo9B9qY7/CMQxNWSERWf92ERbygVKSkdmjQqV+eNtVduc+qdhMJ7P9xNwmXeXq
fzXr4Urma5BTC8/mXBoYsUpPDwamPNcxNw4zv9kQuUKWnrxkFsO3x+jlltWSWGBystZTSvZVTcBC
1sLkefj86HnHqZqdeh9kYU87iBCWsYlKtzMIc5Tf0xiW/vGSxpI7WLzbRQ0DTuER43UQaSqH6XDL
2pPwi9Dn4zJt/UqBCtdE3r6R3EwoLaR09qLF7aE/Y1Zb1+LBUJMgpoT/39ntuNQQb10EFNnAJx5Z
A+Hk2WrxJ59MPGztGp6Tb9hXM0/J1cRyBftcPEJS+h/5pxNLfHvYIN5OZ/1owGsAC2tbJEisJmFj
iVhvQgL+RMRPYYSe9OJNVy0c0r1z0y57SpV92wrpkWRLcaJ0fCYTFe2tBPv0hTQ9l+kVVZGNr12p
blzOq4qqqEcoaho3rbOIpzywIDSu/4sZlJVTuw0TxgJP0IOWQhGg+QYxd16yLkubfJByn1bnMZIX
lhiFKeJDD23s4vIesL733mZfqhcsvDhc98zZbX6fqmldqD1h15TVVb+tg7a40avEwq+vKxC+Fxun
pAqcXGtdPJEH1ae3Wvzy9Nt2k2EdTuTg9cGVtnYLyALkkxVjQ6iq6FqCnoycHs6tp5ogwOs9mQ86
3sKS/0fVgf2RyLTG28DTcmvT7EVYzHeQfsR2+0Yv/26h0Am8SfaF+bvBgH6zULbOpYwe9jSgy6C8
ZlC1V49Xv18jYFx3z7f0vk5pwLLWqWzCzlk9Svl3VSA/w5/Klqu395MSJfSM9modO8kO7Splya7E
P7pJGVEMvuCeWubrhanvRSpxZYUn+OmPsHRVZTN6UiB1Ch79Mpnbpeo4KcAqaxvTysflDlJ9aH9o
HNF0RahPzS90JwTL1tsXX4zcprSjyty3IuALLJNNnFVk69QItHhvQJWRDML7WRCRYSZZh8kwq9hB
0RSPu2oOaJons2o5oLubHLcayK2SMnK2qtDyqxguiVmDa4FCrbye2FwUT2+/vuEhY+yKeUyLF53D
lp9KaghJDHE57+Lw2Fdu00TpA9t6AoGlWt1OkHJ2JXRx88bSmjy/FRKDHxOXP/6svtnM+SYVATSx
b1zGuZm5zAvbUfYGZ7k8y371be6JrAYM0Ii2UrHSrzwJqkU+qd+bifVFKTUW1JxdUIvHC2/qzAeH
H0tiU6jKp86o4+sie8g6UqoFXDND0MIl+Y0RXJf/TqTvUBUd/Pu/ybothwBgcrilMntV+bOXr5CP
M8jlCIASC3CioPLXl6YoQWw+p85dlfxD//ssy8tFkbO+mhXJ7dBxnd2krvdV//9przYByUT2faxb
43Yk8dSCP5M5oGyvKXoov1XcDKr4FKHt2RnMR6LvreB09p5M9hcwEwAR3Je7LMnfGjNiXy3V6ggx
dDzDQhR44EPUCTz2+GysyeURTjprlIZJCJFwntfUE+k182gsyvhWJ1lsgKlf0InE1VSzxTuYYxsu
/v6RHzowRNcftLZW4W8zQECvkg4/ZTcOr/kB2IKQfq8fRaTUHpjnjmkzw/u5VvP8ocUMtP4xW+eu
TB32Td+YH6jT0TmH6ySlcF+50qQfqOizDyvEQibv1cICPSPgbEyBYGXmOH44wpZPpcVq4YFeA+s4
c2yVWYyL9DW1pdXSfcwPCixWR6SB3YHreiGerkv8jEndEJdH9uaoo2ZZpa2olJdSw4TLsgmfqVce
8cF3KLN4DZRYL0quXEW2dxG+hUkGpylwrRPgu/BLSBzIHR1PB8j5DLcLh+kU0LKcHm3do9rILu08
vucFum6pa6ezw+uujkaes8XgjnJkbF3dlzxN5tcSRUmvpJJzv2YRFj5TiFf7obeU5QnqSqfabjyk
wR5JmQIqcYyKpbaSv4omhmxAOzhZqgKEK4ZuO7NMRF32Wv3C2t+/4ABRdAW68WlzSZIg8a8p+8R7
4Hwh0LifpDVDixdsaHwyhmd6nLw2xCTxqLrkaaAXyy8kXJALlsCw6i9mvEdXTOmDZ06T1Xax6dsM
mrDVu/2mEWwl7e2G6anC1xpPBHzbS1Tq/NQk8QqsfiNLmzRrjaplQSpY0N1BzaGylsoWBKlj9VVp
9mcMjY3OLG0U76OZNtneOuQTs6waPlvNOV5PyCvwK+UNI/trnypE8Wuw+Tk2Cw38jeHwnDszaPy2
gX7FgFSU8hMWnIZisPbbXpn3/lTZEyRHOskNflU9zNZMh4j2a2M39MyuqN4t7Yau+UARsrfvYZnm
BqJilEBDcSAlZdDB5oB5Fd7645IXQollqCljT+sV3OJaz9oFRwRIpSw6mdHNAqPdQukcIA72GTH9
k7FWa3A0z0L442LpYxPlKYOjkYmlQnsRkhikC2MiqPvoBUHU2TM7r2b8CynmpzuZL6rK9AmRlw1T
JGpjDbRoi44drfFXvFZs+TrKArlVewTyhwTc1Nc8felvdgBOlnWwN4wkAF5PmjFis9el8v3x6hN+
N5addtPM2Pbu+pN5q/sa3PIZTs5PbQqZtqg9eYlZPNKV7ut7Mg74PxQT5bigih7L3sBwRhOOIllb
S7LRO7JbZzfpBMUOlG2sF9GLS+6fc2NX5DANH54oIRoAIbZxD6LzCi0aFHcOQCLCQVyVTNxJxbQH
0gjiVMWbduassqxbiey9hSNIwFPaZxY6R1wl7H43kDXOeiAkbtIcCRfYrlKHP+V2y/5rZ1nh0CS8
cfBwAcfROtreayrSKu53JtXM1BeYJGS0JZPHOtb718TkiX/eite78z3JG2Paq3kxo8kCA41Ah5Ty
OEPfCh1wPI9fEyxgWgsMPR0rS3CaVnxYLrkNEzE43nhpPa3JAbzPJkg6c1Fl/4srNTl50UlWjPQp
T6Gorai5+KocVuvra62+lazPfD3Hbm2UlS+G305XK6FGcV+4KkrTknYVo+8OXnPhIXuI4uVbAO3P
KhEtIZJgseWleIun9i29Wk/zWI21/wpT08wXamA7MjQ6hmkPk5G48CCEg6XrX8zTPTjAxsvZwhah
1DfX7BlcE9ZbSNFfaAbunO7QRq04BwJyzokCmFspdOHwhRUBj8YiTGpOZgw7T3vutmeY3OxIh8/w
m1GnCmLgnSq4RMvjKMSr63X5vUtK+7updsXaHFsSm61AcdniVrxqXNylytB9yrmmDSiu1f39Qn9V
V7S8HZUYMWdPrybmORLaQ1KPTp+da6UQgcKylLFWuD3SQPtWt/hWAQSntvE7mdpd8Xn5E+Tw+/SB
wl0Wcc4mRvD7mXvAkfKembOLGQv890qXX6iBE0DAxg84qJqI13cz4xrH4t9R7qPHkH+BTZdac1ZZ
IChn9y3kD121x6tPF4kMtLEprfYr/NL79E4krh2+fIQhIDOZdVN974c/fsxTn3Ak39udT1mbXrd2
skIBGWwiBodODuUVrfAZ90hVNzzLSfmumsd5F+4x0eONxgkLUrL9o0zREFM9EUI4+CDvxx2PHgZr
7BCkOcGtlwCalvPsqDzUxzeHSEOaFvNm7+Q1kRAloZTAiWj8bVskr9zJpPCwZbI2SA5GyXVRxmkh
nvuCGGi0JZHvqatNoHZh0hOxU7HhUDmw7RTKXxqnE47ZTSufsJ7WxHm70MCcxRImKRWMtjmSq50N
AyX+/NNDeY00vmaOUkiddPJYunbzk4xXcXgUCasP2BUTGluomlpJG6KHLNuL2vviwwIlpFzSLby8
CQOM/yQ4+mwgtUfbkS6InQrP1vXTwSPrjuVgDwg+QzSjLUWb+9lfXcTwk0rcC7C6WghzWyv9JwLF
5x1Sv7eayhXPuIqHGUWNncMNCwUMWiFgXEbPCQhqNND8ICHJCCN1K4D1RurcsXFta1MxjgDDURq9
WqXlfRuhuQme7/pR11geAOoJQKWm0vfOwYFm41akJtZCra2IgAqC2U6OdxnDbAjmTYcUY38jdP4d
M0b8WbqtXavEhTiuGlD7lRAgQGXtK/BDGZmSJlPAObQgWBHofCMwlcFeskI8xytbSZ9s9D8z4fTE
Lg7WWQPWxljwejBukTLvp1KX+L+URrpvdZZjQ3Zd5vrkPioHvET2Sz6k2x8CEgYk8u0cVxXzQVKr
SaJnwCq+J5swtbTVuTqcfoO3zpuY5kYPLDMaik9L3hTRD1DIQRk7Bl7XGxJJBjOGO78StnmZG4vD
Azggidlmub5aQXd9J16tuJN3+drh80c4gZcnEYIqnOT14snNqIw70+kcvbDCG5a1LEG2RO/T2pl7
bGfx+gPGnEGUtOhw5V+Svw++nwJv0ygwK4XRvtlgMaVRzc0oQWQo2XA/ncN3eMS2chwAk1L/h/ET
EsVRamuKxckthHx9AYezrHYQCQ1KeySnEb1r/sbx3Jp3S0k2CKkQc6SNmBJumF7f4nZXfQYTZEbb
g7InvJSHwjmGSxDtUygIl4BdTOSBEieaJnO2N6jlfYwmkf9Sy5WoHU7QuZG+nEHFyxda7Px/+yOG
x1kzi29/9otyijX2y14zTzaLP3h78u2oilY8FEE8i5k544TRFBra8ghBjT/tTaaqjJdszkYv2oL8
z26oG7fVTCnKIN8sTZfMm0QKASM9Ccdcsoque0n08dEGNUL0e0JKHgtXcbkI9vFwzsDs6O18puiJ
ZiXCzHBC08MIr3ocd0yiTNNj+sF3eTQBD6AvNAc0H2QSPKuxllteGjciUAjbb4PZhmjI2XYj2Rsg
oxVkchCSL3z9eUY5tAY3DcJVSRKM7zhtKHBPU0BZcgUNvJ9Y0AkXPL2VvCSkDXe4OJJT9YXuXiYS
bPHKSn96PfJlShfIoob014T+infFB9UhSsJrivvRURQJrbm4fyEW4g76OFn9f14gojAuuNqW0kfB
1egeRM35uB5lqJG0QBBBUfze8nMlZnFhKOh+LSLPC1Oe60jc/U0C/TvwBbd1F7RklnP2PcIOiTnZ
IzL/BCChiYGC8g0tITvX6gdowRc6WbhlHgjAmtx+5ghriSekbGy7y4nskkkLOxXFAP5Zsbc529Qn
gjCevMJuxmiPEzAJ6iNGtCTBFHfHSBYFaz9Go5CgTrcn0/EDQadpNadZC3JjnN3/eDZ+XgZL+o+u
b79SVdKgDUNaAOmSUGiRazi8KXFJRVekWx72MR2mjS9qiV9G7mUbAf98f1L2ja0YLZ6P4mrIvcp+
a7lmTyMe/DQLTxqN0/e6hPNuPH1q0l/vNAGnBzBG68VzYi8H8w/4ePiZEq1apsghUFpIb6ntODcd
kgVEBtYATDNC50AFO8QHU273VmpvV2tIxXwvgrQpkUvqRRsgOn69+SlEa02dGfm7hB8pcPWabAri
VwFmiO5ki71rlQu3KSCV75Q9Z/sIDRNF476rexMgcbtt6kB7HgUYdfFhxxTblhalkPtUiCHc91dO
N1yTCx70Wou8c2HWH2jFlghRj7wmsM5p4bYRY9/dH+rjLmyPlnTELWLYEojro8pLFt9EuJc4C2LE
mfWvAd/p3eFPRap4+nfvEiSPIsJ8seq1W6e5ZASiX8Kqc0B/adwmuoQbSYAysD3myALKlRkYROuN
whtxSJIjwSG6MROC5y3hiYj7QauTYUfc6RovKsvUEF8uOanocKSATOwshh0yTwU3c3hdcaASlPwG
KYgSepvGgoJqJzJFYtX+MSSI+SeZzGz+48ZFjUEmfUWOfdElmQIcxxM53Y+eTUVV6IlUunHEyxZl
MVim4WpuXBLE1TKu7ZE+fpGLwNZPJHjvxE64LBecASO0U6ICItoc6YrtZpucMZFI5ZgTMeRUFGvZ
XXLRLosJKcgXoE7ZC5R7jWOQIAU6GfYOz16gw9CsEpjJh6AWmrF8IG/NWA6KGuAmylYPsfhvbiLG
qpH9MFPkSXT5F1z6NixPpcFcU9OaRLAb6s9plgjmy3A/WbnhzcrxLul3E+KRWlzMCfrb5stVrmna
HBO1bvS19hFD9Wm5tYN2i59FbqbWY1jNVYNwgIg1cRitONie1UyYyBwor9CoIVVPY7ow6XbKsOI5
dWZLzQWF2nTVgeeo7t8D4slMEK8RCk5Xn4ZYvVTZ1xxR0s7n4c27tgEgMoTcKgduPpdUN8NsYzF7
EG8MMbT5inReygBT8lQo9EwS8LFc1BrWRI5FZ4sA5Y5kdD1b5srHlARixxxdenHqDUGYBEEGOtsG
qs94iVu/UhoX6XEcOlDYdEZd3SmvoxUcVahU3XWD9akg0XEc5bdYoovHdmtlTk91o+vZ/oPhaXJD
04QO4v2uwyPMKmhELwHzJighwxAo/pxTbAnswEtGHqCrF/YgpEK9n6NUiDBoKFkXZeaUs57QfUsW
7+1vfd29YFNjYpr6CZd2b06samko0GvrcEarT4/H9lAWBVvBYdMxxSIJLGjufJ7N3gaKmPusRV9D
Bv7LyBIVwBmPYXOX9UzDkZ9LYyfbT0MnCMLtL1dMNdRaDarb+hEhDmLapx5xjXQGkFhRFqtDM4+P
YHQYV2w7WBCWQp6nysCyp3+C4ybdb/HM6jMc0Bc5YAwFmqrx87woCfcfYkdnwmvi2c792OW9zH/c
B7dceSLxFbQDyVPLmvoQTFE6GM9ksT9lLslRNUxwAb6WWbeW2OznY3SPNC8J3ciexi3UlCeglQq1
L9ZEFQWGe32FAXVl8zaAyjRrJmEtdxGBIlk44S7JshsSkuUUUCpA7mLQBXw5J+9q91p3uPMc7uGh
rwpSxRJEy66egMYOZDvN9gf3MP9rPHnXq0HS55/3kECbegg/YnUsydmqnJtDA0U/lReKespl8a5H
jUgDAudZ4M15wfN+aTvgLJkbuwVYAEQ1zv2KShRSxbKWHgkgb7JX4HNeET9GF/HkQOMVNv9fnhE9
hmipwWgYq33JrH2GPaBCeiq/UBED58myXSRv+txYJnBibzS5FWU2fXOtU5lJwJ8dR4BLKJcmtehT
rj06rpNFXJ68ozEgfIvNYWd2i+A/5GS51bRZ6A6M5tZryD4L0XiXApKv8NFY+sUl4xShm2c2ODdw
ulWwRLdYRFIbraHeDM1dhmWKyH38O0GMbeXqu6V41JMHdDBvjNa6TaVCO4pCtHyjufsuu1RCfPkM
oJI9++5xvrawg7vTteL4lJjRNL9I3oppgcYzUHkKFf6uuCpcT7b2z/DK1w9POUctPvtUfVsCb+0i
s4iHxAOpeXYfhORxLMBGAsFTBCpLUVNihA9FAgJItpHYoIKArNj1Ugv/6RgY4tuUV/oy3DCuhd6A
Kun9kJqBpYe55uDFziOX9PkSflDJ9epQSdpLW/2V7YBKn8y8X3iML2ADnU0ZNBjlv60vnhieSdUA
0ZBtyn2BNpseH1Av9tyLdF0z8fiV7FNv9kvrzDt/H0pFc4N6ozAWOfasm8fCAeU0kwNoD6Hq0HLF
9s+2PeKsiCHGBByn6NhgMaIeanw0suu8zrgZ4FHfCmrwwL2YwSwbS5o1TsaJd32mmYH3Et6KAPrb
6+O5ScMlD477GoBQ9QPw+UkaroY0Hk934gFSCdVUodt8xa6DJQ9s8COyOXmlTliOF+sSvk8VuWmJ
O9DiHAFHE+Yw8jNKP9n9S2EHeDGJ4fu8Hopdh/5l2yZLbUFyoJotUC2AdbPY4uOGT7wOLYhq+2Rc
7bhDD5E0NzB9XnaOryXZg1qKYI0LqYbGXKEMPN/Sln2FS6UZXV3Wl0r1V6e4mj2rLWjreTYiTsHi
IQu0NyHSlYGxRucy42bU6dqkxhWGhSAciq94k55ficQv55MLV2LuQK6FaOst8c+rG9y8pnFdLXCs
efKzSz4+KZwm9Yj0g6k+bshXjcc6xOZLLfSqkcMFEl0arxuSxGOd3ambwH9qfOkkhP6dKgWGvuTp
b/QXh6OOXi5NthPfQylFDUbgqpKnxb0FzMvUQnznjev5MUhbVMDcY0mJUMJcDb7o3ZY0chsSljv6
ro2G3gsVoSme4Ik9dAalEEwkEB6eUmFXyUEROfYrN/F66mBo++NeGhdPc5/i9I/tP3n5m2i3oM+R
QAcXx6ht8EdqsZAGvzn9Bi0y8jTh4GhgCpZSKkwEj2jPRtVanjkFletYsesqoD4rssghx1UTAZ6v
vxa621g/JLMBZGUEx2Gzf2VlkEj2C1ZZwbaXYLhnGMspqzF6LsPPkEPJJQMrAFYobepFiODjg5f+
6gat3gHyMHahkJBcH/1xn6Sl0Kr38eyZlWyYmOluzhcitK6Kmoskq4tGrP6IweUHptXBD2TbFSM3
HUeYuirKMLgeG9hj2VMXg/9ph4WONVtibQeIOHOHl+Z3fFUYRXHnaxzIGTNzyGaW6uwA6ev60Q77
Cz6Tv6lpvftOvzleHsiuqFkNWe7Vx7Ajt0IT+D/dTHDX6pbZnM0B6DmV4VfWuY1sy+etmblpr9bZ
vAR7lzg+WOsmdAtevrRtcP2ghAb9QxAPg2D0GClLwy2DEC3PH3HHJEAhSdLKZpGlo5B8tf/sqHbo
t+RvUwJTO3dGlhM0IlthMwrz8pGqRdy+FqPqCTSedhF20elz36bJdYlK9giASUb5ig+GCj+OjTIk
oz0X8NtY3447+kTATJinrLXQ9GLehBgl8R8TG+gE3yIBA4OWyxStFiKiWH4QXqPTKa2bQzhbZ3qp
LUhmly8zlm/uF4fBbJlzDGF3lGbdMdzO+ud/WAe0xFSSIw7OD+huAE+fwBAQ5+a1pX+KSyuwyI5Y
Z+eeUp6SrjnSBILEi0amDJE/dpOTa3+IXaTwjeVYCF2iZCVZ9kzO5TLH1hx151BLLddsh0U2ZPob
Q73FhgE87sIcZ/MmLRbX6CweLEgCyWJzG6+mmMRrM5wF5wDxH5D/enhCxcjoaZQi2kefZxMMjfbD
8CqPtLO6JmKZghQMOBa5rD7QDxUUXR3ZhzmKha0AxnGYQ7db8acR7aBNp2XfSaYRqIS536p2gVAB
PiU4SuI0UNpGqJ3cAkIN89ivIxXp5omNrw8kkLYs996yaOG86KFhtDOH3n2JYfcUuM9SOyGU+sPg
JE+qfUjTDrDdQgq4iOpJb6IBnNPqUDVj3vmgRelWOm4+A17xeSrEzszvB+IKsFL6yL3pFvmVjiRT
ygJe90asZmJ92uDw+aJ3ModFqfZLofnvgwkqpqCJfnM3+uyCcabfQnJvBjEq8SoawSgc8p5k/tqY
VNSjZcANMDye1hwcLFYmtKFo72NHskojF2yzeIHn+F5HZ8yXGevgCB+z8Zzhs6EoWIA9LQ5v85YE
vJkX9C5aS9jl93Y8aJlMCMtMDxRdTGXgohOY/R83kx2fU1dZ0uy325NE0swyB5Xg4xOXVYawtEoF
kGNWt/SVa3yVrMyu/t3DLQUlsDS8mzDjRIyVGwpnIe2bdge9KdCgxaZ+MhFzq5VbTWcoESpzscgk
FPZ9CvsjOZf2UVc4Nx/C2hXnidiuAIji5S0jtA9kJKYKlhWOrUDryYUku9T8rqrUU1E2hdLx1LMN
qtmglO3xgAY2EktnUzff4rjQ1Y+HGljA82QjDdrS1LBtCZCqLjxKwRbdcQaskABr0TPu5wdykF0n
1ifvpZwVlPOiPovepHcF+oDZsftIZtPtOPAmE6G9MTJDoLT5IQEj0vPRvAi50XLFilaCJbHxA+Ji
wvx9wwXCS/2AYkRpVwH2qGkWsWKlJtzo2KFsDJ9fahmi8TehVqplrajqKSZobTcKfR+A5WulqzDu
kAy0fKhlwhcNdxbCcsCHYIIX3kGrYjEdBp9H/wttTnkwo+cJ/pKK4rzfHFvuUG4dYnK5m3YXfVqX
FbCEAZY0IVdop3x9/umTIomlyK8xfeAsCHTK0eZIYXEGnytYeiNvm2f0DwlgaMDtTI1UyNaMw/w3
B0M/Tz3kqClMwjtqhZsF4QTT1ft+M4Xp12VuAxDfGpQgjj42iumxaTHJWcWOjCB6GVDrLIKiBfCo
i0oVn3J8KMZsuMYjF6GGwOjltDQEFHucIFtriMZsi11xSYjkUi12iO4qwCG3yNwuRwFFVCUGLsHL
Fu5Tiq+0OSRjgB9mlcOWLLHckAijM+AXBBdwIpA379zO9XYMn8S2pCWX+7kVs51uaAQlz3Dn5Ku2
DlgIjUT9GL6U52Do21w0QmvJYM9AZKd+T/yktLg2gMqqTMMdazoXbKXEuHUKWLNv9/xWm+1SDD5E
MLuYJlwB5YwT33M2Ij7lXsrUpdCkQjkitNo4WDqH30Vg13XTU0jWnZP0p9E8lLcMiR0dUUSKteQA
5J191wLoQkr1nucpbw+mJVFr8RZCoUGoBfh5e4e4je0KFtKAJAWVBrekTgOhHfowOWRbik8gfAbd
B0xlDmODTBflWBvAUPHE5aqgMR68aG2qa3JvWM+RAph4VnLhEds6IgvJc2qMpz2g6lG7x10G+sLI
35JWNBWLIHNyAcpxa3IbqKYm8D26VMNaCbltVjGc02EdeI22WbKb9hYqls87QVKxpdMzAG3SsAC7
/ujf6xDdwUOfUBE0G5eKD9lHYUZHFAfJJJWOPVEEuVEioPYguuWztjCV31beP3nUv1YJd2WiXQFX
HE+ok31OIZByZffwTheJw/OjAClo5OIpOKFS99c5TASZKiSxmCYLwuWSYXLMgh8lP2+FB7ZznboD
pp5jju7tS8o6HsHMcrKxsdDnBoGWUnRmJCNjoZvOaDvPxFShZRL7rHZQk2I+XZ0++FvuCynOHrpw
+R0Nyvs7t/r/uyZdyl/1e9+vWOjCViBv2+7Kdu7gkltjQpZRLbeRm1eGHBQDEobFTFz2EtI9NOVr
Zjc2geHI1VUGPAy8BABiHChBDcWeuYdbbLxs8ylSJ47gR2PAwj1b8ZxfcfjCYtQtoy+/AehahC7B
mtbtijunX42H0cGfRAEdQgPGNTXDT1AOkM52nA4GpJ8qgl57vULltAlvQt1gE9304eDSwp1nqOI7
lMxa8fClV375G6S0M03wlE0FA+I37sP9fcapWe00iIsa/q6f6n6WH5s2AlAOthijmCSGE/UyMZxz
Gort8EtsJ770a/hfwxmxw8GppaSHHobeITCSW6d2ALA9Y2S4F8e+g3o1a5F3vXRw87epivthpZt2
TZf8+fd1r+FsqnXOKrk9klQ2UNYs0mEj8zeCAcdgSVeyNzGnTMc3NueewbA8/d4dvpVik8Vz/7kb
o1pID+I1A0e9of0+i9t2/7hiMeM/IrzvMMSE8SBQTTdgea7u9MLbVplaVTCFsJO6NIds3RS+g2fI
yhIIk6Oin7s8nOSmfX3DCHqJbQFlXrHD32giKq76XAZN8BX+CAW7yNFKyn4qdyXO6BEaaz8LM2dU
zXPzzDyAtlzTuj+D5H2UdbFPkpcGR104PBi2EDzP5pwi9Gj07p3q4fa8p8RnAm/tJiQeQN4BcHqU
3/4qkv2/xJRtY1Wov7XTtuoWSoptD5aREFy7Is73miFBtR/82rxFlqVoxGo1c5vfkoSt6L+NRMJv
taKEro8fmy4o0ciixgRlOGWzCu5FhIoXQqyVDt4+2DFTzsOHKmfZoWGFwqLpfmkor41NOCqJn8rj
suFckBLfA9WoN6XILH8JxykbrY4ma3peNJwwPmn+TyVlFzL9brFAxoexDYtjafgPYm4WgTz/ef6p
RaWrL7p4P79Rjef4vfiMZhHH7SBN3oYKEMxNRVwqUbZ+VacjFabACZP4H+j0Yp5ltDzl1/6ki4pX
yrp6O7QpW05vyruBW83uJ2OLqsh+dqXkn4/dE5SSAyPS/LgInVpujOoYT7n3vJa1z4IV83QzRgMe
+uQDh/47boz5dvK5q3jIHBVqd8TbD5GzVn96Ll/JRDrYpH/1MrXyJC0vQHt+1PXTRqowc6uZpkg2
LQmuh63mZ4wOFt4T6q8TWk9MFBAih05vS5EHbzXYD4Ua6VASdneIWIvxFnT7bop42vf0iJ4WLhKq
psUnKIDcPUFojKJTPocFqZNOV+zcPEt1QXhHIqms33L3ZnX89qFEohj0RLCxD/1+iB0or58r42c8
RoNDLa6FXGc49iUUzEN3M9KOURQLCU+pYAJupldoqeA6kNqHzisre0wez98Rs7NwX8ihOpRc8NMr
C4Eydt4lLnSfnDUo1mFS5OTVYqMqw9Cu5L4/ZzUOt1K2GaJudyjZonz4IEh+LnJnDgTKts+DP/OO
VVo2ZREQMN1+ntR3ijoN3wPZ12r7DfeqyuOvQHYwfKXlsWAkfsKWiIc+S8qQ3+Eu0scjr00vvqta
XWhFMtWff+NkcFDHm14M5PJkz6tP2y7cqbICVz2rM0vQdkTUFV958xrME8xZTgpj5PHg3OkLY+f/
7U0UXODsFU5hcqWqkJwsAGIoGI3SjBz23/FoD9Y10d5wpkDAvzmCJhwnFq8lP2SeE+QWgf8Sy8D2
4wHy7IOvgKN2fVnxhJY84ojQ4lDnmlgA4b9FTGBwzK7cbopWH5myB/LdtDSRMsD3slVQXHN/JnwF
xHUjLHBeSNJsivtQfv6X+abuDvbhS9atkquRfeW52zoDWY9xrGSmgcASFqPSpCB9imuhVhPybvPG
Ejdn8EJXNxsoN5Yj2lZR8X0ytAxW+SG3gQJPBuj0ftZEnVu73ni8mKsb+OJyDH2jPw0N85LkRJ0S
T5zrPi0EkBdaKxqai+W4f/0BRlEyjww84GLKynJK4bxzx162lVuxT80USgFyr13dnNHAz6qBy4Qx
quiVNOkttk2fP6CMXOoRzOBGMl0TfbVejjqFpmB7+FmXldDPhFQ1CCQwybRlu3KMcfEfu3RdZxlU
eo0rU6JuvoPj0FmPO2ENuSzOUyqLPP5HKvb5+C899BwAlDCggwIjHIXE6XwaeBdMIByeGRg5LR5y
r2p6ENZX8uXF4QcVZcXkCHVqITmzrtG1OkGtGADbt8l8/osXkesvxCh8CgPOwGxQmkr0/PgT+0xU
T6qmOXr7z84LdSlNdMH1fZo6wB/4TzUaQi4QEYSNbmgv2KhoL2VGdxJinKx7Xe/yx6j+h1n0b2zN
v51XV3dpq6wpNBsIQnhYH/P9Fw7VW4KZXhksgfMz0iFGbqiAV8Qlwutpz7T7qj3mqSQLstYhI7hS
Le0I2sR5bh4L+WB/LWBPkXVdickRo+tZwM78nwdo8x/prjpM/JiibHfnCgRJAvayISV/s+bvQ/le
PKA9B7RFg6eXNExtDSXAZNPE0JmvoGzq7Kucn8pcbJFTY1Hmbzc9Mr0VOTl6Mqo7U1eruYK+AXFL
IsOtxmyNk0mKrkIe3vHl3P11i/FHPAkqQAjydg/jHdl3Z5vxYIygzdmjGyrq1tCNst4watBhcvCg
qIULkhz0+6JPxWLoduB7T35kPuu3eIHnLfTujoB6dqqxT8zlONgQxi+4Wb9w90HE/M7Z51wenqzy
Qm7WDpl+4OSsu1zEr0QKiOe8ipa40+DobGxz7i9TxVMtgmMUt3UbOUONoiDU9rrXo1M9mArlF9dO
Uoqor+VmABKJdoEfX1d7RBHDY2Fhz3iPwRogQj0FU3l1n2QvsyJnG/UEXXB7xGuIWXQPKvIk2+R4
HYq4seu1Ij1K/VxJSCYy8Lp3PErLsqHPfahHxR3grJkjH5wDC1lp6fRkvJUbhQWAFfsP+idR5GyK
p+BZXKVfG8sGsDphLgXymwlrF3K5Rcj0TqMt3ifmfmtvC2SaA4TyNg9gtbnT/DQrNTSuATVlR7+Y
0uJDnccZX+IbesC8jvXae4WmJvMeoJ0WHBcaDeyO5j9AHmjaDXfKPlNmANwVtBAvqouzOLqDn1zr
LA4ibKYUNsf7fHbPn78ZAQ8Zyx4T090zdkNirlYb7RbWLYzf7a9bwe9JHtpuc638PkFCwUea+cBe
zgtxwg6K2mDuGRPSg66OpNEBfCHzS+U9jLco22W44rFEC5OUzXeE1uhY/62fGcqVv1o2Ls7x7JpH
Zx1o+v08m3xmb7GMm9KbqTXv6D4PGVYWBl3prM8C6b5iqxlh6A1/sIMkgTBudfCzJB6aJSBM9i3X
ogZQUKU/uEIvuLAtfTlDri0GyRbWguCdN4VNqpbjWDyJNt2Zg3b/GjulLLhf1hkZOwLo86auGDFh
8pjw7opO/zeMQY9hn+PkwkcChuU4YgiTWPeQa+pQw1I070JGQ6jPRXCFH1ny60eJjsCdVG7UiFFK
7sP5q3eA6isnpfePxINTIJ0KfKigzPqfFneaCViXlqIRNYSD/TjlZQJabGyDHBHbpt8QnNZHRlt9
7jU67WYkysTMOb8IR9PCigxUMV5uSBHz+r13JbhqlNvH7lIjPCQ7xG+QX/GnKZTwUDiqr9sQRs0P
Yj480pg/z1oJBwKFYZ/isiFT9b1Ijn5B+D4ZICPtEvb/JdzsMU/uNVUN3/GM8HiXFahuYESAgGW0
R02EQH77i8LzBG0O82mqP5NMINvU0adQLBDBE40sbXPgFG5cfMv4bXvGIe8MkFBmKxdKGccw3vZt
VR5ooxtgdnbbFBs9eL7fuSzGIy3cxu4dXX8nskXgP0cHAltpQg8dxs0cMMpYLqdK6ugx9A4+y/tI
TVyX4Ui8pe/4LKbyF+OLREyc3lyeyC9ZqeqIUKKX8X2nPNmhDS8KVo69yyZoJ+DX5hEl5G7TOysr
4ouS9Qy1nojrRn4gN9oduz4HmVFVO+py31a3gCm7WJn5SP2yGeoTtNvt9a/TXbVnnaSbaMSMvO2Y
YpMFtpgsIb7gZvqVdO+06EpKf/xiZbW5IBJBKfe2oGXx9OSabNAn/W9/qRaA1NVVAwFjBDpKTSDc
x1NolUjhKEFiCUxInpbrp5gBpYu+ZEe7eOTOw4HEr7XVox0CXZcnmWhwNACBVOBG0ubJPAzkDUJI
pm/veZE3BWD2h6Jzqlujya4qO8Ta7yKCFUorkQ3Dv4SyphxrQusJgtvHr1fNVL/JdvlH1oYUA/vS
K6I+7HkLM5VhHhE+bV3yCx74mG2LPof0g+RA5C5pvdLtEfsCJEF+5K1JsNu/zz+Jk4LqTVXHGEDb
MZ37gRPJsjhsGUhArbYf+wMF1/XnPSoiNveqbidmQmPFFRvo5JJhWLCzvMutgG2FMc6gDqduME8n
gycggiIDqngOj5qKN2yqufk2HkizR0ktxMts9jJXNGjefw3+sehF4L3/MlY1yTEXjweiBJPMos4M
l0E2hIIYCRr7D7Gsmn9v/hFg6+ySHB1hEG//P2kJoj5MkeOTfofHmS+5uwMFZikM91VIzkkMnjWL
Derot9nzWVA3tcEKy8F4mEDPXP2Ymh8t9k+0x4fqg7CqtaPrdOAKAQebsyY3d3lwazPEYprtevTd
KOD85sNv6J1kxRDOzZwEDJ7XMr8SOiPUGlJmD3opwt34OKfyOyFZzdBXVbARLiK85nYUoOyVXcHD
QSifD7gAW7+/kGkKmI7//KJr92UjhkSd9Il2dwccL+ovkdc6o2fhHxdQ96tGvVLdY7lEtRFBvypC
0VHlSnPhkx4PE+bWv1NedMeuKwqS0ljf2e7hV4wBZOwApuuv3mO2dwBDpfH01rZ79ouy8tQ/w/Ah
20wIILCWK/XlJ8t3CEcVrxiIk82DlaF+sodDDN48p/U/w6e+hyjFWcmerDV+9Kg2b/FbGqVoPmyB
K07Br7+TwV29d/KAWSA8fihUQwu+3iJpmG5smIRL56Y/O2Jq2nyRRaWD8rtFOMDne7voIpdP/utO
IWjOND8rz9IIM9AKDF2B2nrcrm0eoCW/E9c8XZrZKT2EpNShGfYfUuZwvz808SuvAIngHyO+WKL2
TUN1iy7AiUsAZvazzK6hyxuD/M6PgRYxEy5uNjWkzfZArMfwysZSOVe9Dc7JAaaqBkZrlgykTBAP
IfeIZc9s1znYB2o2Vy2do+KCtRju3EbvnKuA/tGOgiT92EywCvfR+hJeiC+nIX+zhwMSV/nRpmMn
yybjKOmy60WuxCoVkd/Va7rRGLEt8R2ndHqPXC/gFL0pFC9XaZgR3QtlbhwPisNfF7m3tnxs2Kuq
5d1k0NZoBGyCqVKOLY7EWwC27ScBjhbQt395/R3JhyOy3DiN6r3wvucDfV+0P/Adibw4ejNQVq2F
2OpbSB0QJuxkN0y6EibWunR+k0bBuO5Uxx+Giokhqj4etQEFGhBMK+7PG3YSWikndcxQahz+0KAx
4ZoSYj5Lha217Mp4K71L9tQhyegLDgrBC5gASWRpvqzrscwKCd2onT9Akak4YM/RvoLXi/DyLiWZ
RvoTxWnvAAHWptwwFNmsU546VtnVoHA4sBb01wJ8l+aSkO4JrNpdAsrIAr3M/dH58a62eb3iSOl7
ElqreirCv9LtPo9uC1/uSwLFnpZQn2u4GD1I2oLByPrfdDnrrSWseDxLp71DkkD1T9Z+ZAnrFosG
etLXPvgEWLIFMJYrBX/V2NHz4gGb+vURGBDqP3p6B350tjopStOLAejxstUoYz2B6aGlriYI2TOP
2JOgR3qs3XSELR2NowCLhuA/9mEUUblcLoZIpg2CDIbVkzk8JNyI6bLgl57B2lC4XqLIZ0gNMHZG
fr6oQKMkifsl/BC6VqMNqXhDaYnUzJFmQw7Ycd7KDh4yZH/bCtWDLWu4VKNYgU/oe0NEqGUn6qp2
NSOQOrwZQoYX8Ns/zuRb8djQPRGi/1I1pbBLBC10zEEV2mlr7wZYNGCGsjaW9QfQUY3ziC0caZ5K
eESykKTn7oJO0ENyNKMI1iJrzfbgMih2Z6TD4joju07vLRsFdyj+ixxkY/GlA/+VTC/8Opw2umr1
RXchgCTXXofaMp8JMPK5abNT1KcgqDpiAic0hj8dd4N6dKfObV6cXh0Wu1Q9vO6lONPOKt8maAlL
Cui47owJpmeUH1qxjaeeORRPNjalwLOkEfYhNOmRPxeukeh/rr8SHtd28nQ3iZQ04Pyqtl5u9DEk
Hk0LmcCkI8qC6Wd30q1WGh6QmIrmgrJaehTUSCy1GcIae1DFYWAcZqUTVFeT2VoHsYj7dBgS9ljl
zF91Z0mOQ1+YkNuvWVkWd2dyxPcm+I6N/mPwS68iD6tAv9wVsS0Oh4MkkfebdZMo+weRLUWsf2pp
f7EAIzopyJhUnM9N4a80Dy4vfAJge9ZgRgBtRcd6Dr5vne5dLnhwxUoIeAfnZEgTlE1zxjbYlMMH
FCye98xbCwKYvO8MD7xAglstwsxxYSMSoWl6FLBZCv5QJwflgv+EdPy3PZ7sz9xT89Sy01e1vQ4X
wmPxlxDtiEJh/C07s23PyXin2Bu7LIFu9NxuJ6x8PguJAgCQv4aWGh0Ax1LzDq+7T1R7GG8PwUlL
SilPpQ13jnD8X7SZGchBYYoNwVYv84QaoWWXuPOp6EuQIp0oLMJTx8qLJPuZp2xesJfbZTkferNd
smcBXLr47MAG1gpXuDi0Vv7rNVBZIGgkF7rlrk7sO8RN93DFY/g+leD54HUaiifYw1NqHtx7MU5p
D2Qu1yiQscA+WL3mjVy+Jv5pBp3e42RxuNpKfBGzcZAAoOgrQFW1UDPtao0Cd1k0NiWeY3kq3R2h
APnxj9AqeJjtgZIDo3Wzce5eGf5hrGPdAXtjjao2gc3mKbThfYKpNFQg1hLoH5xbnRIzeEAkPgg+
b6P4k+YKLZjnmxxCZoJ/UHNzaP4VShZM1lbGDKS2MvVsZr+il/uRlJO2knsI1RIk6HidCPaflE5I
5hAuvfWq5s9fJQczRn/RpetRbBWmOd8KC1//RW0PRFPT5UHH5IpGAAZeFNZQOTrztvMvHAG/C+4o
ks78Dh1G5APSPrSh2x2bpd/M6HlwGSFpx9Yfs2F0/AvhVKFd6NknATtrUwqrUrZVzR51K4spCHga
vMrrd+Ytyw0yBxV5CWIRVFudZQKzXHrGmJOzlFTlfPQHyNqLlxwZANM1uXOBQ6imxohF+3kRWkrN
/pCDDF4u7ozhW6rqmNDnOASu70qEZKF+Rp+4BANV6B1ktZPKZHbNHPwGqN4Vod69uqs4xs9upC7Z
9NHD6H5Of+ZoYDsMPCC3DxmXtoF9W6bUTETrq1AMwgaKu/PcdirRNGo5h1XTSyQEEA04be2xnWk5
axEkqXTicp0HRJh16PIRchObt2H7en2b6VHAt+Oykw0T4g6OOy3fk8703VXMxLLJhe/oJexEzfOg
b9X55T7HY9E9nanYgc+OCYcb2fvNtdtS+co6x0Dszcj1DTE5je6X258rqUDE8zOwxO94rmHA8S/Z
ulwBiGDjGAgizhV4jpdZWj14PqfIEZqs1Lsq0sIMQ+pmYfuxw3fVByaB4EGcz/hRINUAx1zJFb0F
W5/IKE7EaVUbLkBNiw7O/xR06CqUBKaW7HBiKF2rtoYttmFINgDdCkpxYXn+BsIMeBh48QRrCN05
0x06YoveUVawzMh5W3ymvs8ABNzIMgPUvELUN/UzLgsSb/BYdiRIGaAjDT3OT/OEqXFFSjjhGvFD
3uc4KwtO7KnnThLDiGXyqTlswSk5A2nOYx6wX7T1mp5ttP9kqAluwjT8uYRCWc/PlfxdjbtkmZyC
NnfF+9mGnD4pGoSiLjvlwOtS4zdgIeHV5LHXRueqviQ/j0RyedWiR6fmyXlpSd3ec39KloGnHVzu
imu8vT+ARKTYhu5TL0dALQHYc/Qv9Prll76B2y7vSL5wCvDgOmnm4nDvoqXhRQY3xM3ImGEBqjQP
+h6MwPCYqJr5b4UbTanm54QYbO3s42I0Mt3J/BVdbaB7quh0Kjrigm/IlHwKXgdn7EnSYcZmKkF0
oVGgbb+9ArArS+LCmLH1+OyD8bhUiCL9zOrekeB0nfOaqRkI/noLcLGUKGimdcsM3dBTLterNXUS
81yvzmi9w+bN+UQAz2eAAgn15WvCKdhyIxe96KmnR73+adQRcvgamdY9yys+r/X9AOAT387bXPSt
MNUpqM2FdGUhGCidpV7S/O5PZFro0d9GplHM1a2YCrp7lBFTIEG8CMFIbqjpCaiBeIDzhYsW+Pi2
+kJy4NlRfDD9JCH9kmNxes9w+93NcKSfyzJOSOn13I8TzpoyAiT26MvHxzOhoJA3SgoHywerqXpF
r/VvJgVT2QPu47NQ9NwuPXsyaydKl8ROoEdMjCQWipufpuAD9jxlpa89xuc3lM1h1pKXUjDUH3lz
BbA8ieOyllQYfXDHdt/QQDmn2B3+ITBSoBy4K2pprXpgXa8NdhCF2xYyIvVK1UcJbZ1f4lT0nIsj
BQqZME68+ESpQFu5tXXEy9BzY0NxlDamt8ph3rDm9STtY1jcMFK25eprrrCPPD8iRGGGyKWfU43H
kiF0R6mJ04RgeOApSbb5k+dExTqQWMdYW+4/3GxeEs4z/R8ALG7qPRfmMfqE0FPjK4wF1T5jYhBy
GOqK2BLaVddzbUKONgg23I4lfwaR1ftjWiIXC2CGNq+FuKqs+yitoNBqO98Zuukk8Xf9//2MG82r
FNa07L4VQ+kE/iWHR0CJkvFHoRIEknw7dWBg/cFPcyj9NFVCnp4GPIfJauKCXIBcdvi8RC+M18bi
e65SGc9+yt/QSqaEy/LpsMsF38R5EI23+z6hLGgX6cPXr0vIsDbNdDr7E3WYCc/g8UakZXsdvRTs
GSJY++g0XCABsqaNCQsVMqV2uYG/MoZcEPh8ZKmlGOtcrUeJnS23xUVuzHE8tE7i+35AOwZCuQLa
H8ZBgRvsi5NEbt/vmA7ukU5kLzw+3zdBqCOvdn8Ide3QtVtgiELTU35p58BnubpBCJAjOVEDTD4u
neuIiS5Fk9swvKTte6G8gH60FiESDqIDlvL3GrD2Eby9uTy2iG8zE3J0Lbfn/YRk88gBir34Q1w6
kG5FVn768RLbhDjH9wJmLVILN+gierfCWFgZyqxbUhz6pwL5C2a0+k49OoGBZQ2UwYuoPwOfqTUw
nLD32Ei2NGlzEt4bTzIBnegdXwvaad2rCqkwCuR/IH0gM8CpSx9yV0PT/OD7jfxc6HunFJoHqJTZ
w6bB9JIilEkUe3rz6X5q9iPXrzX/p4lDPeUiNA0PtiWuvCK3jqk7nC5jncD7NRknSViorLTZbiEj
8eCSbpqoIdEJfhsZ8om7gomlGbC6DP3ob5hMf/VNMviraAlvrUOrFBdd6aGEBvdjasWz4jaQXw6/
lJo7chGgKC/e5D6YfJ2DRwMWQkwihcJdGTndPuNF/3KzgsrxTb9vp/LPAr+We0aw1Qh2YY9YTREv
EHOGkEU+gOQ0mvxHcozstauOZVlpdxaBE73sJ5XRPTvAnqikFVoXNgoStmwMlqAFQNDKj7G72dNu
YMFhLj1P18co/rGcZuPc1jnsp6SvubLo/wkFWraGKdthZL+BvpiXwos2tBbLe2sQS1fL8p9qwQkN
V0wkIlVrzfCAOZqobqlVXHCwMSoVPL0WLdNGIjh2jf8av9fMkpv/QEIcw0SXS/iMO4MlmZ666utl
mIuk2PrhXpeUcb9sGK+gyv9EBsx3k1AQiHaAINB4UAaVoifRadyn0NImlkLVxV3Ai31YfSXz5u/E
sqID2g/ybc6JkUtmiYtTEqAmPdw9fJsPigH6h9Rgd09lSe5eBito8CKFtWnnQYjaIYUmtf4P+Eos
Z+zxLkGSUZdaF1Jv9sIJMwt1TMlu5yj5keYK5GEgdYoqOGXmHDpJDDSaUok3YmL4NPxEQoWpbuq4
QQ4W7LTIuJjkcVetDiLUhJ+BKlklFWKhqU2nbQ286FNmVr4+XE/JSDk3BVIJw8cYaN0UaKsrO8XZ
cN9Rdo+0hegZ3uDEx65g8BFi/sQAGima6+/LhDvtC3JvsLGykmxhJyUZEZ3LhrCquKTNDZRZ0heh
iZ1T5on8sJARs2CYeFJ9YUbbmVbE/ghUqUfxIPqit+0AZdqAsHPTEKz3C3wjBd1NKO+ErYwrqUma
ngesfeS+/t2FCxFpKhMMk9X1QXKaACjDhYbpKh8yam6WeLYoBh9PxuNQ8jakBC8nNY5EaOdYxM8J
my/NViAg0C+GpY1Q14qhLui4eF0JDbih03tSKGYkFKB1R/5H0ZYN8nxPbFf8yYx1Hxs5KFcTYSH4
a9mMn4wUG/LjmHvLVXOTwc4shCf1Ap/5EKH1a99krKrpxxwJNlVxBrPasNwz9a2mnFa+Bf2Ltx5q
DehJ+qpoEuxmqIgb7Q0Spp+cWkHYTBgtCCnSLYyWyRtuCE+MGI4/4C1Gxgn7yuGA5yOM9Q6yb6qD
Q45UY5WlmN3oVTzZOnZX8Bgy6OS0SmHRXrvkbvTobsLTWYNzmX9yRABTYeK7krphlQOGv5qEbnYQ
cwHys0k5Cf0/KGsPA5wJySkS3nlAC2BVOPO5Z+r9x9TmVRrJn3WIomlbKYwLzrsP9oH3YL+BDdMD
+1dWoJxeY0dBYeOlbpYQI3OvqhU0vRVkQPgkWG8W82jq3Q4Tlh02ggjSYXv88OEep+hgwJv512x+
thp8TiV3LEhLKgQLo/Vs1/MXwMgJbDqGPB9bCN5Cjdn8eYoiGA8N1CgLiCVUw97VKxZ43ml328y8
QyFKZUtaHD+b2IM9VthGFgY+5exZ//DlJrbVsZwME8OfjsLo2g2fidPOQ60vpnINYX0D3qFfU31D
fDvdlVgcbVqQOzD9o6xSnynxZWQQPW6WVGAonSut/9lqMACg0tzfMakqVCmMV2wKE+X5AHFzJHkK
Qr/lsceAJAeiAklh5zFdsmr7LsZYxqtwBY/goY62nn23M3oS1TtdLJyWtD41Uvsf7Z2HFuQYKd1f
zAkhmad8kLAYF/AvBUwfwNGQcrCdMHX7aSE9URgW+EOFYsrsXs/UiTLjmmOmP6XQMaekhVRJqpT0
OShyxhMTpPazsdjZUSI2C2sxryVS/QnF5elExmg/lI/+C63608fKicc8cPr81XcftxCddfKdp8e7
3daRgGpPty3rECoGxPmfM6kiG6wU3OB/YOKnZzEZ1joNuAiE6MMk9yGqa10iqJIxTooxfAbdhPeP
usEIP3ZW87OF2YHpjYt8Qb4EDQuiKEsIVggheLI2aPXk9opjnIqgoIlN2tzFZYLHjeGsyavdjR5p
rF8P3qM6tUPJCz+rnR2HQ60/HDok+IQ/gFvtOwLY1IjIsh933Vs4D6tqzs+qmL6qZdDfGHaJloRN
hWSVa6Br1nYdV6svPFs9gtWXe2Ky3hcyX/gMtkCc2g9cP6Zc0oHjZOj3VABMgeuqpEwho0gHsP3j
I9B3Co7M/dAmImEt9SiuG4JZHsBz+yDyss5taFkfAbivEGxC7Th1BjcEXQU037lUrAUKSW8X1RBI
tSaomOFXR+xo17BOhST4+MSEkC3q4omfoAt+4oD8NSzuP3ARMidAW9l7Ix7MrJyGorhs5fZmTXTv
XwzMyAkn32YrcsXHrwa7JD2M6qZXiCAqV3uvzJCoj9TZfq3ig8Ofvx6StiBAKjZ8iSdRhEQx1kks
uEKPbc8vJUVsRGoVKaDsQ2xHqVY1Bo4gz1Z0xNNEFzzKPJ2zzgjjjZMhBNEeFoQRWkZWqeIZ2zZY
NIbdBt8TwVGnFi6AmTYoThCJCBOickfiDDZvTGBr+GtvlyHZjOOtwHR9jfKFKTNG8GC+dcUJbouL
KNCouOdG2ViN1lr5dxkC2IGnacgGejiq32dmSa0K3SvTEEVDBDDB5XJk8CEGRHZoHN7x/OBLZbGB
R9stesi2o0O7N/QsKU4hDVCtpdb3FuRMsSWo9nCGD99fBAw+V/ghfRKNNc6s76/rMcsczgqSo38p
QTac//IMhZdO0ZR0yqlPyHmAOFjtqfOM2JlN1bszVJdeTLP0BZ3wg7SqwHSsBwF1Qt782F1ZITqz
qiYHC1P3p3bpHcSoHAN/kxh0IEajxdD06n0IkV/KwIQfRJN8co9G73sN/yhBP3BOhpbVeMi8arVS
dxOweqLPmBuZ5L3Aq3izX1T4hptUZI4kWFzIHS8TJP1xtFGdH3utwh4twtzGXZVoqsBLib1HCBLv
VVxwhs/DbrP6kCQrmBCRYTdyLTUhO0msjb+OltcxG6f97ITXC1Ao82xriqZch/+uDf7ry4Y5mIdY
+bl7/Z8ZSCGhjXYxeVKu9ttH+WK/GBJPWJoHRWkEncmXtVEj3B4YPFlVctVNN8twtai/NbDvRfJv
dDiLPTXHwSB8CDlG7TGNrruYEczyHKQ+S9sNZo6Vb1ouvZauvrH78I1h1PBwzTtw5t1H7iZyEusF
UyaCUTXyVYAPlh3BmTJfVsmsc3vJrn3q4+WY9WlEkzPL15wWBEHItxnf2K9Fu4gUN28/vv9lOZrh
fF7qrCn7CDyZg97nb0R//GjHIrlDcHJVsYI8HrMzR2MStVZ69FIssFQRwi05W9zpIXGD7kNeqhno
pDIWCxDbrx6EuP88WOQFWiwYj8yaPlO1EiCSFwivIYteWZdxpxxpG18NnnUI17G94bA8NJeY5sOh
KBgIaOIj/qQsEMtmT5Iq7MADhNobT6YoF/URXlIVkSTBRkjcmNTmc4r11wPKBZI72mVBDJzkGj83
leeNCK823SjAr3701fHyvEvSZD5NEIh0KjPSDAeF1DvlbBSmks8Htbenmn6Dx7jHSr2XXuWctx0c
2D2NJbNBsIJygd7vjwzFACBPOGQUtgOGLVUoc09UII4xkyJfNhNz5fm0GqCIXv/kXcAqdYmDdYh8
T+Bv74I/204Nz8+42Bbk+JgGNR8WnOhxh4GfEU2fnWd9hC8VR/zAowgZoxdaLlev4gMbGcgXynqd
LRvC0d1jj2lj1hBC+shiwpetewmNgPCGQXXkMfdFYl0IDoB4ox9LKxHckoLgzrEnpPfFUMurxMWL
icMEIh2rltQLV+uiX3/mln+XCNWaygGbrvamxF8XuEndGv3XWH3cNefeUiPxQ2OYXoEU2xnWrl+R
2I7HTUAZF2Cq4av0eVdOftyKCGueBvgB5tNTSL6QjnaSkrdWwl5zOuGDIuSEbfZSEbLOZasE4BfB
nAlgQpbyNyUcv5nG6MMGEj6HIdkAIZFdCbB9jKafDnOwtpsJpah8fLRO98hyC9oTd5ckauC7dT6V
A1EBjJMqM29xwJxef+lMeeV0OcBN0uQACAN6nj8K7tBLYfnXrPzMmUdq63DWWGl7BfXv1O2VSUay
KzwQ6MruE79uLjUCGTxLzLb9EV2r9yoCCpErYk5MKrJ1TwC9XPo7upxwP9VctJZTQXNA2BuNjWFR
/Qd3RBy+V971g3OyLbti54QKSZXXEAn5D2poNqxb9szu5bAOrXKL3QYc1RwAsINnIjgjoKB5nYPG
Ko3LQSLycxPHENGsg7Fd7ZHK9Dv5uDfo4FIasuFVM0bSaDKxy1D1X7IxcUgezQc/BybXgKlcMSJX
2I1oNMnVafLmze3IDrtEeh/51CuXxniJdvuy5ezqXzy1MOg3C0eSJkGuIjORiFXUUOSUuA/j8eo9
zIqDLzt9Mee+HWHujkMhq/BEb1ycTP4hlZpfrcfCpIExJxOb9W+CQYecY9lipELc4zzCL7YLwjSE
BamFwIkWGkrXmBGlBWksSi6FPpXE6jJjxCP4A4S7mJZXaW8zHqnWOu1LnfB+M1tJMVH9xaCSSFVx
xPJeNMiZzuwbrxUovhDGDeaGTQ0w9GR7K6+fQGhbyciu2HXtORQ9xyB6Ru9LfF2K81GBVV5uf+p0
2pFR86MN5Y9cAu44yjWqcCKCVZ5sryzYukutyaor+hHF9uJskrRzaxkcni4+yUktNVdbPMd3RBAY
9JW82KQ4W5AWqgTTai+6NbCNBJJQyraxpGNiBDV4TD+C+fJ3ndpDeiA8ApH3aJkiQtFvJl/zbqsu
W0f5gGi70qB+tfgIbYBVrmxq5CHkxb6xJ3L9fmjEqb0/SsGs30qXOAEN+NypbPOJ81mbRLPJ4eNH
r6XZQHzwAAZs9syf1zOxQm1w62VhwE18bSCouoIau6KisLTDJAOnBU4luB2adDdL4Kncg1koVHur
6rnCK1zwnI13JvABlyEJSUQMp6DOOi25xPMDJHA+WmTMk2Zil9LCn5XcJ2SHQdGeWeiD0GV3Dlwt
oX82OXIiysPJK1nc04w0nOd2RD2X+d3hcEBZRYSWlWPMA7lYhEKKsXyxALIU5Oc8FZSrYVrosD7E
os/+uU6YVSU5Mz8iMfGGgvAXS6984xZ6G7mU18IJ98TyIx+Zmdn9wmI2JAJBZfskfrJPZ3YpUJvL
BH8Lh0lm1vHNaoF7g83IXsXIFyPWF9+hWji2940eIj9W434NOCzyybKbmp3V/tg49NP5nwB0onAo
cIsXT4MRMK4xQnt97/cDGfEB3GwQnjE1aUDTQ26IW0IxH36rA/oBwohLDPalPE96Eh7OB7fewBAY
sLVoJzabbvr0M2oKXiLV3NPYBnFY+ahsGZkGpox6t84BUVqIOUsvam+lrLwLtmWXlShYzcB4XjFm
ZFFOkfzzFxEnYBKSk4OGmRfi8ZWgvG45ucvvP47WiI96TkSfwUmRYbgiV1r9lF6qpyhueKVjiNDq
0u7U510jMThj2HdpFlmiPxVw/bm6TXvpVEjAbKiKxA72dN3YHYiTWSPprSKzUiGR9SyHZJa11Cwj
UNQt9vunRo6J4sZbnRVG2SN39sL8boCx/cCoXxlLaiGoxXiaDdf/ihY6TGI+31z5W6t4jlXw1o7h
m9/WmJHqo/KQNO6D4/q4F81/M72qd12I2oLCcdGitwEQB1tX84zF5DSAmcJG7RJObGcPtbgM+p5a
2nGUfWneI8n01rKeGpdbO9/Hm0QVYgzOEhCKxGhn4tWJl2L+yc8tSYEE0Q1RcKWHLNLdIaW3Za/Z
qZjSKBP/5hUDiWIG3rJyG3OWi+gyIQ8Oez5m3b/MAm9l3GNnZBA6UCTvXt04rewJYZ+Qw8AH1lqv
mTo26lW1S4JV7RvO3KmEof3n8MkCXNZA15LKwHk9i15piKggVkmuV7SKkytNWFKbjG8gCj/lPMXO
t1TQXEh6gd7B+Mq8np2GTYdMky8b/s1GlISg0KU3v94iVJaJso06BZB5PgbHHcnk/wU2g0jlJklI
yTh/O7pj0bX77FAQ6fG8PkfmQa+FUOwWxfE5xVaMj+4jqNFcyA4e+sgC4p87PADy/ybvQYPiFPNL
3SkgplLxFyjgwViVyxD/0915V04jzuspew0iRQ8JFd4jaA6n4ZShAmMeHvbzKz8mnl7lQ1accEog
uC1va0uEv+RA+2Lu13bTFbSxAwLRWmS3lu4SwO6DIrktx0Xn7GFHO79zz/vkO3ynQ+g476doytVs
5UtXLAb3nOamyivwgbAcTsI7Q0+yST/wtz4DtLkuW48oey2eO/LHPNAYfWNAmcRYU6OZtMmko8VV
Lrv9CTGpmKyJBm9ARuqbLjP1+nH1VJMbmzeDCWfNHYIsbGGrjUH1f2lts4+GatxEtJXypGlT2oEz
6c7JA01TWy8DccAnsXZFRtYTWqRF0XZMIAH9r0OLod+7NNjiQFnLTYmr87QgdYDfDpdTa4DYpry0
rdLXS8awT7VaVM0EX+SSXhvwRn6KGd3VJay4jFPOtTeuph5MBn5Rg41qsRo5WvoIYiQ3xau7GFci
yc+7jdZMextQp4TEOqp9YnApvastLaSesfpR/AWW0db1r8Z1EsFDLxqRzqHwVTbDX3ROdmdRMzS1
LXbX7hEmHpd64lijc9S0K5Kt1XMhZivYqN6YdIL75uyBrB7JiZu1xN3YDtYA3tw2r4p/I5wNoSZG
jNAzzqRjOJK0aFtUSkzvqG4Clroh+J+Qz9gSovdEePdwSitfsebF4S0VF6D+wdCtmfkWcspdLmYV
yGGsBgUD8BrbhamppPJfPa88hDmL1V8fTgnr040kRl5e+tcbUuZKttt7UiFQXRkghLaLAszhMgmE
dLncq4nbgvfhDtGUjcZZ9KG86SHVuqHNj5gMbGxd9xvQ3uOy8BcO/e0TAFPnPBDMMXxiKy1ysMP1
mPzn88eSwT3EMIf1rSczh6Jx0vCBFNYgDspGSkZkpU29LzF/XM3B9O01ubTjqgxjb6LZuX+lqMFu
2atULF3+5UnF4ygYJyiyxqfX4o+U6w4nOdTyCYoUz10yvFMy3bBAgP1WAQ1ISPI0boOIEcQJWfNX
CE74rpQgEm0Fq+bTX9eNlrpffn0SKlSciT8oSXLsv2Lmz/+VPafWLLu/n2UwNLY8UUIXQlvutZ0X
k4wOjZ9gu3/PIy1ytaRgw2aJYyTJ//U2dFNrbN+ifxyuqr0+5oG8AMjyLF9J0wCi+CBmWwYdMHdS
OCIlCNLCIsOOw96IAoZpRHlJewgpcWJN1jQgr41mM0bvnswVSP/AJAabXYotOL6ST0PsbZzFUpGn
VLLhMbU7epEC4QU3PFbtYEBu783q31byqPw7V131VOFCYiK8hpb+B/+gZnoyot3DNs1svp6rlEtL
ZTKJYP3cJCxtVmTa6AURSTEaOjy3gjVZOix148tW3Wh2DpjvXUdjRsJ/T2MZLIVb70fwi3C93L5g
Izj1Cy6piLSUWPvcTVeESF78rVmQloh2Q7Y/v7VSGncMDlXW9rGU91fMSFWXi0+QvLJuKDIfo1MN
a7H6HEYe7pZgMfSjdVfNcfHPVe0LpY5mH8WpLJMIQeCr3QtjDFfUYLKLvX/F9JrapZUCM1QhXa42
6SdHXv2jnvsYu8UPIK1PQXuiNpuJXkOYWc1foUdLpG4ibjD71lAhZQ4F9a/BUXGfq0zPOglW0z3c
0Hr/jt4VE8hbaU+RCRCAv1NwaJoQbvQi+VlqGyfiIu2wgixkDWyoUuKXLJUzCOAQNGzKNG7cJgGU
4sxQ5zyxaWc471Dfl4q1mzw7dflanTKV2AHj3inb6ckLTmkJymUI5lVIasOhYmoJqEyNm7Re5g0J
t3aPry2AJCz/NHkJ1h20gjRQO37BJoEca/JYEG1TQTbot+RKD8vt68svoOBIBdmw8isZVroGIfc4
oq6fACuVAUY2tGPmfX7V5xFzwyBib9V5cHSDc68AChfSCJJST1ccsBX4b5039vjEIcLftcVDF+PL
x7Eao5yeCoEgj8FgYA9YaNJBKGCMvi8qGPAqNP9L68cvH2z7yQDIaDpP0lKBPxMF/HOH0KD6YAAy
7u8UYQSxfqKTfvTwq1bDxZGEBfyOFmh0vQwSrLhgjFz0TzFcynxxH8j2G2QxZ1wL64BKN3B9RvXu
Z6mB0cuMbJ3BkDY/TQuRVJ/8q2+H1CF1T/lbHTdfYxDUFWYpjHrTsfhyuePkqEYWrt4JYXnEr0MD
GN61CtgXP6lDR8wTb+jQy/o3PURcr0vmDWYkVliwAI96l8BaAdh00hOlZOZ/OgshksE/GS5DZat7
7oMfnMGGH28t6BozSbS+3qWFNr7QCEVzXLPu5LEmhyGvi4S2BP6fhF8/LPXhGtF+WHmtaiuoR9SE
PXYG0kVztQuLTvYcvDLVfY+iq3tso74mvlhf0P7gskp0GFugqlgDJJLp876JO6wvHPiMQNtfGQqq
vtl4QtB77gfkcjzhrHCv/muSQMo3G9UCLCXmbqmYtWQbxzaBbLdgFJ46G6iUP/WY9DD1654pD4d0
r5wVlEMFsRyaB8/9esupEKBssoQvJ5gHBqzMmjyAJ8INE4odl+b3GoD1aajTpemfk1OI7KWrtPhV
ND0h1gNOZxV3BwRs6fvSaPe8reVdi7T+rYYlMgk/X3ZDHNl5f2S0Wlys8mAMXueFkb2rlYvMh/qk
b3oKYxJD4fclWwMIT5dgaMiYoEElRBWgiZFjGGCHRYNPxNN29wMuTgwXw61CElOe2ofT3gvlcuhP
2MuZbSVmA1nwZIhsAn6irt4pbIo5fpZJeNjlD7Gkc/pFhhTlBg6eK/e/+f3hSXEskX6Vmvdx7qv2
xtQ5oz2JuEQaA4KhZKxl9JekJi8cfv+yWaah7Kce4bWwPJ5VzROaMyOqfdVfMjtik4mgqRKkLguG
iowsrNFAlT6iETMUAZZez+/p2uFTOaEM4k5nZXCaWp10u6LNDwcmMS5ub/yYY0lXQU3VRDrN4dcA
VHFsKQPetfjzaRBRX9TexJQ7AVyGtnm+RREKJDmI+4CVSNyZ53XTcXZnB9/GUr5EIAHOR9mfD+XQ
Qrgfd5ayg1xmXmpf4bvkkQgeOMImlRjQi/lFMOhFePhOgEDcu6R/Uewmw2KrOjJL47d9JbHOZlNn
XcYPUXFkuAKgDp5T1Hho2uhkkUFTCt/YM55cBKW6CY2Hmlerx1Atse7szPl+GMeShHebr1IedQiT
3TFNsAjrp73gsG9DVpHbQo90QtFoX9h5mR5J7GGTXntfp1IcjD8UK1FAVIvT5H5ih+l46UIUwMXq
4bNvGj8/JW9hJbNextVsj+WGen7JOA2MDWk9edAShPJ07gb9AgBR7hubvNFhEnhOW4hw4ERNjgac
ZiyY8rW7sItTzsF2kNqTOagA/GPdKzlCEUupjfev4tJId6cXb4HDLU1mddR5oLOmrJ3yFbuHnjbt
MQH6HNB0KRrnt3eiWrCdlxvxcdeuUoPi0uCWMmjp3hHbNTG7soWBdEepgz5aKsvEiyojP1yRfBq7
3+bEOXh66eW3f5VQLalD3moSPZH/ZRytN/mUMrpT/+b9Q66nj//rtx+1GI70o36jgVIIVpPgLo6O
A8uh2yPmKywD8xZEembRHDUhd3ED0utqlh0H1t+qzHL3GD9iuZKBb4LJcJFXho+xcAlMOHG6isIJ
em16Y/LpKHS1BS504W0hlbzmxXJuuDBrv8nxJRMW4pMQPfjhS6Vb3OjbX+VaZ4IGol+hIPLLO9Ei
KpmzXpZPHEiEF5MVqF5QCsojXfLh1QvfZghjXSLtn3HwoGgp58dX0Kjaz4WeZLouwGq2/o0lGaJ/
/GerkhTkasSIYsU79hrjdjPBfNoC3iBtQCj/FCVyt9IsiH34Rzprop7F6rljq/dnIc9EkwLG9X1e
UO3nR8R/0Nf5oj+ojsaYLmV3nSi2C+KOa5UJqimIokAVJQMg/wP+eyEspmuO8ReawGqg92d5ZrZe
0rrpcyAuvO/wdPR796NX6js2AiMsH201Q3Kr1Ywfit0bJ8mTLHf0LH5M6Dm3HS3TCZCG2EwNgmr/
DFJU0ljeCI6BOf7ODGBbBvACI2zsSF7+wxE3ZN6rng6dQEb4yw1IJoXOPpFfM/iLssuNgiECL95d
lNqUnZgR033ETk67iKLxjfHRQ0BC2c0KHVFJ4Ws8gTSNLo1+sQK3qlegKlntb+m0V0FRstxEwTix
1s5DaYk7qJzUoJ2adPgKR/hO5WNEfiF3OHa3ZKDir0ERjEJ87LmJfuNO+A0O0gpcIEYS7V8x3rmC
jBDnrmuKHrqteYFtEXt4wmaxMKno1KXzYErnnyD22ew8pCjirUJryVKr+ZGmFSP2YuxEpoStO9Ab
a9bbaw77jbEaDSyhDHbl3e2YT2gXJ2whiFKmBk6k6kL4CV29ifo797ijnKgc9S6LKWv7Vk6iMS7k
btDFNefIzP9zDPmv6cXPqtYIaTU9+Qybkyw5LNngVeaaeXRHU1hJ1LByVqIHToIhHJFxCY/NYVIf
Pwg+xFjzvB2ftsf75QXrPXnCWCtKXk7qAJXxHPK94z/uMpVoD/4ZY1f6fZvvf092KVHisLSj3nGS
hHqx7DLv9YLwMfbyDC5x7RLdesD7Ld6oLDHGO0t7sW8GRgfTvaraso/cyPUVL1uaqjnNEnKzwJ77
cJAyxe1i863tjE6L9o9oH43nn2ld+PCB+H1iOrjFYiPeJyPVX/ZmdnaCx7INqnw9mvgYsXkLtEqK
krX0oNdpA/z1JriK/7oJ93lXCMvSoFezHx5FppwaW9uZkMD7e1IV+TW8QX/yPfPKejV+h+aO/p43
r7Y3gURQmyvq+zEZCz9P1jfkKuLCMUXNdRAnR5dEUgaDVjigc8BdRaBO8c9dHAGooSrj8dolbros
M2/ftjrYIVTnZylWvrCEkyXpvzdJqGivaz8wsRAr+kXZNTdkBi9V+XxJBaCMjeeXA8vsuXuptEHa
lEkRC5uGKOJSeTSs82rYV8WhhRA89cl3Xp6Gun5HFRh4egWPJP+l5wJYRZuGrYCXoKZpZQe/KMA5
LHrQOj59G58tMEx2d2OjNvfB2dewHH7rgNC9c8PZfrtURXyArjTdNTBrvRWn8MQwmNMJ8ycGDlWV
aM9Th+QjigWSI+j5KDZ0ffSls5gYHzW/j8J96kljmBj2ySXbOhnG9xgnIBDExAuy44zCxhMQRhWn
CscsHKtMLc+/uq01OhaSQp7gkTRNS1ANhLTQF0mJRtcA0plFX4TiAOun7kmsnqq6z2ojVaYmPktA
g2oXyruENZOwYxkrGPPA4QQp6P1khCR9aseHtK5yRWPJB8/7qwKYrKaOpZfR27BR8LszVvEoHjto
CCSm8b9LW/S615NyYnN8XP6SfNGBzXfOseawRfLjxuup24SuiAr5wC1tRVXSRf7gNMcni6TmwYfA
AmRjqPpkxMpEeK8Gf0oLurAmaU9LFkJWJt0dlGENlMXwM8Kq1aVsJGezZhOD8/mLvnArYkWmNpaI
A4M7hny48Kkwg7MHJrajesk8wXLeEwSkIcq6356YGhu9xhgm7aAKWR80AZCgz9MKQxzub+Rv2V4j
1dap7t1lr95/6Ghytj6MMMcqy5Cc2WdfQ8LzOtOpAV4N5/DtbISHH0rrIxnvO0/gPPjdQ7DIh8Mg
ep0z8JEDJCSjVvtn8sTQE0zB1UxDtdzXJFRy3qVxzn+7Cj2fgvMZdIBoAz9Frklpf5ri2Jzxzh99
kVPebbKPOp/tJVDBD0FYEBsZ4/WaAvXqee6uOQVWoRl53MtwUHZxIzgZ2qs1YjYTaLbpa1L7zAy3
YaAcultyIRZWGt0pLet6gfDechvGN1rgJpDLhKlOxJseBdeXFsGrQQ4jy2OVn5yvMDRZpxltmdw2
QYhlGEE276hhOYh48+iyqgA7MVflwWUUqjBY0HmDeeJ8Xl0B39vPvHkIUSSmefqJ2YjRq3DHp3cG
Mi3RePI6WBv1BzMVVaIGPHiCzQS8ONMZtpRP+e6MyUKF3U/U1OYF1r3zff5v7OUIaPDUc5rb/vLK
RidCrS5wcv3R9SCW+i0RTj6tSk8jiVluU1arcdwMjWmPSh4/yDiL3zLOvehB8NWsuWbjspaAX4Zp
3f15lmiqqh9oBSD9iupBq0nUT/3bwaj2HZIr2DYC6n/djgYnNNL5SP2jdYMbRcCAkL3RqofT+K2J
zx0UveTN8CoMmwxXLVDR2D65uu0UD6b2rX82kZf76x8tJcEbe9TQwvi8yYrTVfgfULRmf4zzo7vD
X7rVlg77xz8jxmWj70/DuTQZcv1JwlsC7tM5dA/Su4FP5ZJcHaRV21WUfZD2l2O1Q60+S+j2M951
n4Tn2ryPObvs/sGSPDKgVRtLZpB/U3vGbtqqUJghaTV2IgX/yv+E03tesS3Rtc7KHnMOKzjR5O5/
yo5N3sLqEedlQmiRdiNuj5phM9SxWrY4HeZsuV9GuJ1bK6hO5DzYnmAMO53csYMhbzZwniv40AjP
8sabdB8iBzCUe1/Y33DLan/qnLN/xWinAGw/gHIR0ZoLhDrfKKly0zZ5wkwXymtNwKlv9MM06X4e
4PlExBYMEGSE0HmimnvSlhzCRiGAlzitW3f6XxDhk+xfTxReaSYHZoDDlCIFTYNOQ7u/N9XytUSI
AsYcC/IbkKxky3mlJzGhbVGTTCPL73RH4fI8VJ8DAOLIC0U6DNCEHsfsaL2DeC6fAJrWiaRCY9eh
8cD6yreWpP1LnPwKr47yXBiX1O8gtvA2jcQqWtlmjZLSGC4o94zwzAD5zfXyY5BgXpVg2Opy4PDB
b+ZPUfaLuPKu+mLZ8nGWS1S8PE5MXGx40Pbr+vbf3AWmvJ0vAIw1zZV+ZBp/EI54HLXkK9Oqfddb
M+QFp3Uz1PT6MsD/tPpMyR+hEaDBP35p6QqoPjA1TBfU+oO3AM60r1Q0EQ1i7j8IfKHVRBMk1Wa3
yaSKXpPqxBgBxE2pAYQZ/fUZWzgiKL/wCb8woL6FX5kaZXYYYPnWYjm2S2/Uhzzog8v9Z7/gk9jf
CiA+J1uWa3XE3vtalMacREymESgNxRkdleveehjqry6UbV0GK48miBicXKCGcR5bhFYhhEePNTaB
X+i9shq5gyFpIpxHhSHE5W+SQaWWFYc5KKPY0BapeBFvWBdf9rABs3WpnSMX3QHy7U2HEOTh5eNI
B5TcXZUql9YHF2EZ6e7dZVSi43MGji6cBPTjYSgmaKenghPlLY/srh4zi3rGvySaXTozwW7tMht0
C7oJaR2MIKwOagpXJofzq9X+OhPaymcw0X5V2jJ5rwisvJqTaRbqWy2MNrqAadJwziUfK1ptKHE8
sRgGKpy9B2dT597Df8aSOyd1a89WIXd5k8cHoTPiwyo9yKra86VOGDA5vZr0d4GPyK44KxpJheb6
UirKbXyUaPMYZa13xG31J/ANVMGV8DZUZIwHnLneAupqVAesOk9zUQUH9fjEEWBE4AYVTgc26X8f
MRBZM0WEStQEaoPS30cqJTj98FMoSpxczgtYijCcIXAsHLS4ZARVPwUpjDtPjtk6B8Am5gpEk955
bWnEf/OjsfvlAK9z8REiGpfF1fuhbKDjm3Es/8LM7/IUt9D8DJDDqilvxk+HNBiAfX8BYVwGsEEL
wiYX9kSOJTsNv+vrvClzH5PNLVi0G1MFEW5K6GGLTqHe8ncIplK43ffZOl6+0RFK8HAa6Zf0/AYO
xBI6dShjMphJLP8rD+hxdHMYbyv9pkmOeXslVPJrLFSJxp6FMOTs9otJMzIc76NeQxVtf+UtQk7y
XqzsHNRKWV6MpyXcPCtGGvDMlmLuSkyCfaiDc1XXOk/EbXj9Bj3jYD5KQnexunpkfS6TTIW4bdRZ
9qTiN8rIu+ZStojGcosizmI6vEdzCV3XOgePeJAshZuyRuKPOlN258kFwnbTS879p4XFfegXMEOU
r+lDVoW3xUZFuaLgsj2hntu90JDgFErmd7ae/iQkXZ8yr0MzAPKwE/jZo+qfZjZfizwfM23cvkCW
HOpjVEE0eQHOWi+cSaPIDy0ugKddZP+hZ/OcCYAx5LS3GlGV/VZ15ZHDJlrHO2CAAbDYp6dVTMRD
LlESos8yCwJgCfCshC+NJ3PXtvvH7TKfeTCmVxf09dz3bEA+ynoDYwvMIucsJ619qEMhqR6ilLrn
cmy9+FxSGdVDbTEvDGgXXZHq+15g51E6vgOiCsb20Bou1aX19k9OBghPbYdOeYWTP0DR7XoeGY8K
SpbRL53wkr1G3NzPh42Q5AAdSNqfZczh5ILvabX6Ma1fSDuPVZGz3NfieOjWyYuJlrEgG0FjppNc
IgEBI4FcUjCt3g3FL3IXVpnnFchPVasVJCo1C4vy4sWSbz7Mle4+zfR9y37jGB343BlmClMN89I+
ducJsUUMZ+dzZyvgqCbeIswRtSf6PdY9L41Ds1l4r3JxIARQGvj8eXTRDpNymG6naEpbmjAHekN8
hvjTSdZb2vxYBGG3IkWn10jk1YsG+sJlbcC8GVhuxA2E1IqimSOLrADar46DtZQ19ULLDQIWAl0H
B20SE29ENvGop7bUNqincg7AV6udUtK68akF2FtNubhkqroA9b06lZ+hjF9stoarr8qKaCHHnd+h
2R73331MNSEtNzoNoHIuq+wGQ3MOLSZM9/AXnH9vR9JqaBVzYkXfPaAKcUOB8ehglA+JcPRlmhma
QSRGvQZ0kmP1t+q0dBZzdsfm3oX19Hxq8Gsob6djFTClJ3rNSCkhurmNp46cRRumZw06zHwTZLKy
jUzBw+ubU6GujcudDMQe9tQ1EUwR9o2VkAxl+me9+YcRfaLtZ+ntW29FQ8f5Zd1Gqa47kbRjh3jZ
Ai2oDZ1oLVIGn1NnSv0zgi65Gy6C5ukDpv5UVppCwKcnvEGFzIZL+CyGfEyJhMFkufQUm+ZP8fHm
Q2b37evX2SjFas1qlk+8OrpAKYQi45GrHwD3ig042xbLESoJkELem9nLt79sqJ4fcJZUN0K2sUOD
Y66IULoCo1ADyJBFPhlkfnkSS28cxB/z12L8sLzLCRcg4vJN5nB8AGgx/iK77X4V0jWdI6PB+mIB
NPSay8pqxQRMGjGfGqk4lg3X9inO1H0QmolICDE5jRUesKuvhq22RRJ47cxp4gGeMXwlkJFoX3l9
nZM129iRSRU3ddw4OdlkZ9xSwPCAz/iVQpg8iolD3sZZtLNODdZeOuKSfSoH/Po+euHykVS/2Pdl
nlsJJ/qXhh1RWSZjzFfCasu4cZDBbHZsTd2U5nXwQ2JtCOGYel0jhjx0ilPI/rGLn9GsTU8f5pAW
tZONhBSGJMbkrHUYvETIXiRcA27oCTNerrP86F4h9Xn5iuhq+Hgqp4/K1A8nbCcP+7DaNQXyiHgb
Ly2Ak7IF/WtUrvIm4TXS5xvgclSPvJB4H71lygRr7iJxPV1TwuIdzBYZgaHJda67Hwd7cZlN2T0f
R4hLMu84oaRaOI78iSuO0zrqEPoO3akwmfQPtQpFrgev25/Xn9A9bI0yPoNzJBTL+g4atwVgQvRq
Q+mE1LGKi34M9LLASexQ68MaJWxOq4YlPUKPJHTEMrwNfY4hWdqwgbyHZmKZY8pdf34RPUS0B+Km
NIXTCb92YeGs+c8nF9dDq9yzYdxh9f5F/tVpWIKoLAgMCpeyNuBg3D+nlAGWFks7FnjQ1lHSCjFA
U7bxii2rqzFoydJfpMqdayUotQnyVWCn2JGiv6R0bv3mANnE6YXjn0oCFpTSi+8zpDAP9ZLfqRLZ
xuhUffn0hg+Nx8EXD40BbptkzioBs4fEQW06bSShn1HqTILMltaNFlnF1jTlkxnD61Kq5zPsRT28
Z4PPET+Ofy2QZStQ2jOiW4zmpQu5E/lPyM+CnPEt4snKl8eeauKKKO0mGp5NoTzgOx6QjjesjLFO
q9PamfUgAvrL21Xn9Hh/N2SY97qYaNmw8ygDwTSn8SdE/P/HJyn/xq2lnsSW458vlpjgMl+vmGz6
ru2d1zacc2X4aIf83rrCn6mNJPUZvlstEhGfmxpsH7oabnyjp8xW+/3cMhkQVbZIbB2IOQC4CMuR
/q61uwYPvtCtCzggd8EvBFfDiacaRXFn18U2hmcEvNxbJlINy/8UcfYHXqgLFNVZUCXElarJNSbQ
HTFtVwdTOAueyS0bH0H/zVvI6Bdo3gV32jH5RYze2bawEzilNSPIiVaSLleJrhDwno7N/DLv9l0C
cml5lfNLHpOnSWgHm2zBWTsOx0PHF8Nu182I89uVJUvs44FnfaYmfUoyBoIwxYXus7YLLrbJnDDG
xxzBK20YCtnksqHxykH3GrHBc1SZ2jojMUf0eDBhSq+/RVmIQZlOA3kf8RBOHyJOUaaKsDVmf1Um
eY3OK6ZV5VarF4RNc679Jmh8hbB6rfiSqNRi5oFHwVOxMsorgRSv54SaEcEvGVgSZMLApagEY6uM
r5wrQAvBpMS8ZU4FEquRE/4Ry9jZUs9tUMEiDKo0LTkfvX/TV3eR9hu+1sigC4/bF/RkBJPOhUlh
jakWdQo0ANst18Lqe7VsiSKcj4HSIVieciyS8wHHTiSNeKs/vIww4eljp613SwesXnxzlBFjt3kI
w8Bz3rlxE9ISIwf22kAqS0UlTs6iuAHtEHnH9/MXSppwIzEioWvMC2aN/bR1UVaeBy2oydCtdpCt
d17kE5BVYmKhQrNnSEhJ5/Fmj76h6oXuXirZxrKjaujJIeXM6rwhbBW+3QSpWQ3QtxzuYcT4jB9F
26sUuV+pxuxM2wWu0/Yvpd4YuU3HqfTh8zhD7aN/TwEm/yaXRsYgWu9Ey8urISR2KBi0Had0Ajs7
hX9XNrwpzqzCWkNSHE8uxhFLQZoWkV8bISq0QERpF0QjDUgQeem3vluC2QKwry3yZ5nURnjV7Yre
rdvA9ZPWNxnAuy23Tb5e8JHeo049SwBof6RXlWBMNryOLnU/DrYmSQiL4wEpCCf6Np8BM3Gc28n0
PfUPAS3JD/OguyPOe8/EPwe1XZlgxOUE8+75cNBXDOUgq6j3Hfl0Tv1oNOpO2LkCqwrgoB/Os0sj
IIidYsP5fxv37kFA2f6bUziQnFTIoYeJ5YjOPa0UrR8IIIitFSNmwJiJK3361A+ditrX0muHlZ/A
IH5opvTLivbfiRyUXRxC0FZwzxMfLG3ydb0nJb13/Q1rTvfQASniOfF2PzkB4SkldJrsRA9jS+Jb
bKkED8fOKco3Radc1ByeYgCnXfK1LUCUNtaMPTMQewsGgxx1ZII7CzUERSuT2ZwFffMprNPw0JIk
Td/l+ov7K/yYn3OVfdJcqGO/QE9nNyn5xbmQblogMNXpymQBhWVRGOQwG+nxnBK85lKIR4VRF88q
ZfwTyURW1eEdbDhrKCdsUP0fZgjm0Ifn8O9TCZ8ku0+6ERu16dprK3fWbHzgIcY6f6Ck18abGekG
zOzC1wVRqG0wl9jad44mEn/fNn/ZI+M4Q6CyxfazaKNp1FeB0OsPuyEF8MnVjhQoaNSzWLS6bmM7
kUHyM6RZo5v510DmTVlqpWYm3Bkm6utEfec69DDF8q2oFnacPPCbaPwxKFk6hdiRccu1nomqbEkv
SuAycg/6owYaDVTIPYUvYVAo01yZeZ+kx82PsCdIlTz4fmvZieQ8n7eWagki5kVfQH86ILn96e77
5qRMbuWgvfbFBopvKeUpmY3sctYxQzTDN5u+xDICcOM4moULg9us/IdUKUTTlyKjddXfVal849T9
ujRj0wAzM1YHOEIm1DWsgyoxfgsaVSt8r5SlsydqzuPlVKdy+8at08AkW2w84U2HMnkeP5wjjApv
pjdN8qlTzIP3Nrdi2KYUqNDFLJRmzwPnoOwx2H259MY3S6U4NOGmakYv4m85ooB5GQy5PLN8Hdl8
5AVkF6RA8VkjykvTefN8AKT7niwWeoL1V5B71LHDlAciI75ZYrGbMCvoarlNzFdOTlqJfIkkyzE3
5EYfFefwGUh7bxbDc4vBMtlSrqPA04RBSo3dpCyvlt2pk75fx0AfqjfpzZ8jNuyP4fbdPsRnmKBc
NcWr7eVOxX4Ziy9am7EN+tYR7aLtQiax1Sh5s0v8hiVflr13T3hrGXD+71ywyYe//dSCByUGI0BD
g1+op/aw75g9GslnBe9M/c5rKeLpT2MvIhVBL1OCA6OeUqqUaeP6eRtjao0Bl2P8f4Gn4ResQxOA
Gnimo1c8IIIumVl7AHwpVi3YJIlhs51CTdnY1OKEttMuRUxbmW6+IxJd7IJf+pajxsjbMCSXX9eo
lCzsZFeynmhUyDFFcWg3+tNRDuNfQP7XBS74XoDI4zZvA8eq0NKCjbwKcpBY4t7F6cU13hJ9ubrm
zKTW3NLbLygzTsuXMy/LcpNFU8PzksfudSzIb8UPxoUfLGBlB88S1DR7LPmiTCfzlnv6Ozt2Ffib
Qv3eYKogy4O277GmNP7zvRP7YVGfuIoWFd2yHh98VwZlSwEgE2JlP50mTtvXUNoZ3UN6yALpd31s
FGUSOgwm+0twFiKVpKmYEcsPaQP+kuRmjXTEI24PrCe/pfq61PkEckTisl+T5sAo1w96/seTeFP5
iYXWUKjgyhAIZWHfNLOFSB28sl8BvhY7o+/pboz7rVH6WILd6HaRnE7/7myJpmTBjJgpKCreRffK
/mb5+DI/nFfkOgw1v9yVM6UQa1V/rYJV0uNiyasx/lD6O89ZtZZaet9f9MzwIe01twHk+eioSAgq
Be+eT5+v9Mw6OuIhsPAfDlllQFfAAqmtKAADQEZUirHtRHE4L2U4gRozy9WkN398WTEKPl3Qyjm/
+r5H30uFTBPcRi/11NB2db4R0SHZ6Vrb1Vr/rS67mDw0VCQpRMEPBpP2mwudjCUl/Vdk75PAcLPf
JQ7iTN1xHfUR1I7nhtPMgsfwRwGHP0LraF+evz7o2h7IeVdg1ht4QdyCzKB9QsdRT5eYWpQMQ4RW
cwpgogTYbiGjCMCh7MZnCYWtvQhLwBX2up4W4vg/gB0Uk2KlyMNLENt7nY6NDA7qfBKXhKotgAaM
kbnP47I2Z/wU0xXIqPwz1L22TnvgZ6EyOUfYJo8NYoJQSZzpzH/VJqE2vW25IW5YwuZipU1TRkbY
EAzAiqjXHUWxVAfwz8RWaPa6hfHII//WU96G6/3HKjME3jMGENRXgculPnX+7HcGzB3ZT4oZslIF
lF/0wFJbvkdsppyih/QzbAvmm5knPSRZxQ0Gus46oSQAoJVpj95BOWch/VX4Y6ieWiS7yWr6Z3la
iAwCjw4RM1o/3mPfo8FMom/fDhtsBDozJi5SaPgUgmqChoseYHHx41bZN6cd6g/gdV+d1VG0Ql8M
yp1nUs7qRyOQJnR3EOxqJlqih8mdi1MAT9QjcGCCaIr2+Lij0qt5Ls0skX1O8XOq/M2QWk7AgU3W
wZWXr2RK1nzbHnYDKv0yvfdQUQuF4Ta4fCVcpz3royhM61E+DgruDAK1M8La+sTCC6fUwC0nFkg/
/Tx24qDeA8tBu9IT361RU2HUBMmbtfdjp5NiQrCRyNke/1jlydmRw3pWu7mzx7pI8Kblr0znfa9x
pGYEIpXeLRbT+zr9mMEFQrS0VfZvaOPGoItMK5YErJX/D0SSlOan4U2dqYx0qzLN9K5mhY75z8oO
lkJPxuN2MMCmrmux18Yw8F2GlNyhf3+oFFzsBBfbpv1UjkArbk+RSaHe/1ECGT2gWoWXGGnpocTt
2BFzpgJFIGkkedg+M03vxoPLniUR4NVLOf0dXVqNguQ9vGDm1+QnbzHZTbhWQJI3K4ggtKhr76lM
Jod0TAAJ7T39gwGQhcCMtvvoJH7RnfJuzEMGSzmx/GKtnP8UMTCXBO9984xFcJzyI3rnZCfrwfNy
M+DZNtZQ9SVidlcwTYaYsX/MmzcpsH7E3g9R90RMXeGqoheGZqe5XTPq1GTjLKl6F5cKBKIhXd6O
BhDs8F4g2gSKZriCRPV54CxCXdHfzQXtJ7i0WGmRNpHVPRWdfaxKmep1iFrtX1OmWbCI7b2bWCh2
bvLsaNlhAnyW6OZB6UnQjWQBhlLQAwM6ET37vaC6nBPg3WodgkpGB/667WiD5JKOSRTCFSAv37kc
YsWSCU0MOui+jp81hvMFPc+2Mus3IKMhNfvQn3lWpqR4KYE0XYXu2CyNtS0AXGs2qgJnogQ2vSpz
EFTVl9sFMC5Ccql4aa0uTzczE/nf9zXFaJXTnzZ+aFdw4T8zSOPsdOy3GrkrtTd2YT3sjSlbxeU8
0xSo9NSTknEZX72TEipcSOsdlZBHabD2eLV1SekkOdCQkMm5IdR/CGjsUL16bPs7kxDMAro18dy8
gr1nmt/mLLKnbCp+BJ+WwKqtyezSReBCWrPVNrfirTaNkmrdFpPiqxo7ycZMM554H7/Mn89PAPgd
EwLaMRA1sNajayGWHPwQuCbZ3KuJBQYQ43QvMcRb9EGDOG9vZV2LMsJvYS7SCCgzm7Q/RXJBK1Lm
VOWzHxFeTG6LXaSULbZexCuXX4RvD2rciy7UGLvzMQCD5wuuPeYUzNIYD+WOpxLr+Pxw/I7qcRmq
sfQtks3IqdnjGnvTd2MQJaKk6Gk13ON8nUCkojHc6bJCddLmQKeehYGnfahLbpo4/lhFx9Fq8FqW
XF7ztUe617ew1ICqq5TwXGChXRjyzNuPxwNxMFDqxefABq7LRyiIxntjrpC6duH2wSoJHhhqoT25
d6p2zryCqHkvUTf1h45N+M/nydnLrNFR+QTQUv4L/iJZ3d6JnZFoEN+y8UUzHadgmGzj41QjiXGo
q8cPO939BMk8MrQclxi38gv9wmzsl9Irz+RrD9hJXLRpdjo3OQ2uOeJ0MAN3XmIJ5F7ARa19u8vG
qXl/hvGZTJm/vrpyd/Gcr+ZRBWH6H5LK2JZW9e/NSSXGvxAAXcwyxYon1oRRlUjwtXeahCsRIz0k
56QnGjQSUrAb9Cz/+qcljHNjd7uX5EcNcMCwryev1Jh0FY8RimhJmgfEcx+B+ZrscEPquE2gVMyT
gvM8Uswy+mU4sRAzDCQRo9Abz9qNhvCN0rRGkGil1g0DgC8a/h8A6sRYi6YOymEVVhKBV8CgV5Jj
g5OzNeG5AsGBlWV3ePzF9zDZCLRsk1UunxZyxfvLVeiOwso+RNbmGykKtzvHr+B6LEARTRAGrU8a
OJpqXziH4b1oAuu4k53mA/UySfQDskNHzkp/UtW1a2gKRvjkoU8f9Mzo8zfaTf39MpEgh5UAf28m
FJ86OBjLxQzuljVFD5Ir+w9eU1V96BjlOColBCRiJpCrY59X+yzpfq7kGD/KahRDQjiEZgYLFHYx
j1j7viVrUWr7/3HGATqgcZt3NO8QhsziQeXPZVqLh4eQ2I+7nY6cxh2SxV7Jm5de0w8JdU1rNkrw
wh3/vtCAQUVqyi7gbbcmnWmb4dxdgzWJvZFBPujLMdU/FB2K8mtL1PVU9D+1fYyegRBIdUNA4IvM
lcRijD7w5xUL2R6sFXIFcplyLuAkGHSH6F7gUymVlGUf73mOmd2YspHe4woCq7ZY0WMleclKM323
O+KrqLfy1zYNR3q+KVLQUjfFo29KECZWbFmCam0irZqDaMuyrZzaEAvFlos8zi77uYfusnfzGFcz
gH9sc61+cB+2vnoVbLaUThX4A34iQH0BpA4wA+dsd2zS/iU4IIE7ldlSPJVK5/JxDud3nR9LdZmJ
tZCvLErHwCr/7BrFppo2MzhGEGeNcogDrvNhJPoR0jQod/VwfLmwyA3ikWR1ad8KC5dxmNYxCzws
GfLVJLyu7eRU7ISRybsNrQiNJ997Iw5HuRaw6Mrk6rSW1ClxnApwi+pPNR8zXXAGDo/fH0RVKBXm
erYHJJxT0AgJLfizlekvYfOO8TFrQ+hWlW7jbB25YhA+vQ4ta6cPhC/zlOKNm0RwmWzmmZRLmfIl
Fvb0HOxVkZB9Pu/YWBAXsYhsYev9UzcNABRuIALK8bj6cw+992jN8QMLtSAvp97IbIU0Haiy95wZ
Lld/QnrNmla83zmV1M+OGKSBLeWzkI0fuUE9Uh2srtUxvsHbcS3bHqB46uwvnwt2H+b2ggm6nJts
K93S1SPMWg2ikOEuPBOcRseYE0is8BU8UEl2aGjV7NXVYjXQjpB6GBNPZwZdE5zV4emBZ/BNFjvP
4Erfz64tswhbNWoVl0ekFjU0tEJYR6BGLAX6nEUdPO8zAxU0q5BS0FZNDJ/N9zKdS2RaOZGuGqyV
bRIMWhVQRCo7zJUAfXz65cD8ge0P4+ml9yVGAVKIURsNcireXFhK89+WQlsSOSqZqxCcV0cP22Er
Ai5gl4CbUDrbeVEPnHG3LsG2bf2Za9WlqkGxdFgsbVjmneGaT8IHx60kJKzRmguXmcF7zw92lA3y
qIwUR2htstnwgopcZuTTCBsPzYZP7QWPPVurTRCAvDJeeZxOTvf8Rnnz4JY1DNyb+lr+rsbe+12u
nzTY4U6k7nSfNfiAQrG9VlU2QjlbNhp5jzrES9B/GGMhGqL9W8Xxbg5sIAXaNzxleUfrOxkusada
2AU4a9mnmj0ROVJYGhseOSBrFoAZKzr5bJqLv3zadQap/XTBxcr0wOl+Oh8xSz7qBzjbpF0SnJ9d
3tqFjQ/tHBhhbPEo99ux7Imw+7YH/gS8hWndkiCUJZls4X3wQ7kk4N/VMBxzoft4GfEW826UeiPE
j9WCt7yThJPqC3Z5p/290BtYcFtsClPeePWiCUXFnFWFLaqLezJYTRP5d6XtOesMc8mBPQBZL30a
3/ChMKyUGQrwrV2mLZ3siD9G7OGdtmtXW87xTztmVURTLTAOvdxluS3f+/i8STmGZCrTVD3da0W2
cjT8/J8FplI4d6LhpTguimvP45s4EClf5L22f/5hHKfItipJa3obPgAXkutwlefc6sIH813iuty0
6tO33tPUM06Vld10VjF0HDYWqiBBGTMJMyVnBTAruAkgevRqEPTGABDQl4pgVmFf2VEwUVsK6LBf
dWwuwagkF5ec87nI5Hh+wOoIKb3FkEEH+oE7TZBfk3clNJ9qgDz2VDSh4lUexv7VDqRcQ+fd0nvS
pPQA3yQDlLsaLwVOnhkaorB6VNpVi+/+Qf6cuujfrce5CCLbcEc6fQ6MIg+WQxpCOkxJ79QoST3a
RSvHBncp6yt4wfgSCvveLBRR+r9bUd89vgk6BsSUxPtNL/TrhbyHF6wPL3RW38NBRGRlJ425JCts
4+BiREq8XXFfZ7ZqlwxPWqWzdbHxhnDbApSqhtH+y/3HF7hDj4zhoTMhQ4Nf3H5LQ0SXEC5XbhN5
Sol85LK+zjF18nw7/ye7DVBCx1iFI+kbg1riX6miI6LCYx2teVlYSQLVIITKg/rBj9SDNPsnPE+p
teSBq5wB6pRNdgGK9dou4My9ccpvK0ur403A+QqiVKFj9SLkxd8H4tEqu48g7m/i+cZ5ypyDAC/X
VGKG3hm+BJwSwNO+0leiINQ8ODA5x5PQTFi17S9jksaWfnebaU8R10OX/BxKdQ9gI+oP+fe/l4l7
qcva6wa3iLaZRSt3eKUSGLg8PVCxLQHf3zUlNwLh4AEsknxzvGRh89exD7692zN/QGXJtnRXjuHi
f50wL5/d7bpt730n1fSnBr9TqxH7rAySNts8rGVAfkXUvt7IB2mgXQ/A0bXlCnSD0f4HjWTfeKk9
bnjf4sCoc6ZMpjhDeVJkUGoqpGB75VHsaFZQuH82bDvCOMGIurBv4y1pdfF3Mj4ahgsrxTGVxalN
6Ah85NLdogvqDAsdHLU8pde/17f5oRalC2q3OpcygY51lbb8Sm0MVt8YEW024RE6bHpANTtufyWt
Pzs5VxKq+HQdIf5o3qTll4+pLbQ7SiBRdR1svzCg8EmbvL6idVeCUboPy+YOdJh6D8pof4y2UTQW
vAg8loW3aeBstNPU/QdvgMn2obMTYurJva0Y5K/7YsjcUED1VVADN/fkO6t19VNzPf4k/Qn52xjM
ZxlDu/d2vrOzgXl6LBu4rIBxL19EeDaIa1CpHP47Ga13yNoW1rYN8VrqV6b4/fD6vRvjhM9aUrGD
iPr9xgkq/aZq7JiXfMNL6r/uFR3556vd4WqnTWu6jxhaP0bvtKiM8pky13baGLwOoOnhZy8uDl5i
4xD3HEboSqXgF1bYjMv884GbQCTQNt1b/4hL1d/RcfCczq79oR5CFq4kM1FFV0N9QFpMGylB9uTv
KOMytb6jdwpcCAB+d3sMyJvwb3OpSyhszPgpwe4+nt39QyYeHcYAAwz2oM+G7We//NBdXjNjsvSE
ZXGs58bBotc/vpQwxBgUFK1cXNqYXF4xqk7ZS8gdhUk+A5alMNPzL/EJtRAZlKLgLzfVnIykBkN7
W4ThlF9ciw1XGjPooqwTni7WO2N6VhZiZcLf6tWW60dezFk43YlhH6Bvovn9hWLkNMEuBzlAXrMG
28lzjnjFlIKdMdfyDvxilYV9V/c9MZLQUdVE29WNXmoHXkRtcZX6ejWsQrKVor13a3N/E4MqSBrV
DpiZdXZWNu3i5vl4Ec972qBLn59L8HjW/KTu8xPlrqJcChkFbRV6krj+n/bYW2CPB3D9OOBXNs+c
zlXQWpP7w+UnReYqCy1W6edLCw7MLHvTw43N2A00FPONDv6aYTbtwd3yyQDikyR9WL5ieFlCqf2Z
9JEB5sIGgnijp4rNUraSFccvuRbj+EdpHkEE1d853nKkZVHT8WcexWoQyLU+TmEBxlwHvq0NU1a4
Y3d6Bt8tZ0ccan8NR+NwZiCdWWhSBc5Z73k+XbrLoLWlneNuGZN8r7KSBpoF2zYM7dqX59J1ztCs
p007WVkvhJfCY/U+PEUDzjuwPq9bK05THCAhn0eQLmPM0JNkcyZ+LMemrcHvVnnWdVc1KbkFWKvN
x8xlVdVXu2ZTwzf2tiaZfIfztgewidNiw9R0HssOJkHGZy77TbirJRHNAWMhOTQq4jkTfym4DrH3
Lx3j55WTha3cuUdXqHTipmgIaHvC7nybA0iKaliHZi6SAOWpHBRNczkqS/Bevj8Api00CSKjQW45
1m2FbF8hTgHdi5QKg3N+G+VasJpA+M+sLuLir+Wg378vm2EYu75Df6S8fRAu/vrbZpA6qs4aFaCH
XQDhtSu5IVrwlkDfnVf1ByYqtgnFSOn6GxnJsnGmLdKfwhDHZ3ksCh3QPS4ECADb8uHBgoCOOZO9
UXdPOPC98DZzHrAU06g+pqNcBF+4/uD2mim/U2TJrufIo84kh4CSSxAB3xZVPuhY5skjZDgTYkFL
1X39P6UX4RpCnL7lBx53NF7MueUVCaMi4H8rxf/sZTUElILvwK+hBWIR9chLsX3Qrwn4qYzwdhmy
kPzi7h+ItJ/EZ3X+mCSOzaKBxw+kgDveZBssZIdQFdiOCEZ/HQdSjXYoxtoNrS5gSsqs+gocXohe
UM70nP375fPZKEbADF//b78fB7D0ffhWbrB5ouspJUwgpoI4s8sVYPmupZFWdGf6joyLfOU4CHJ5
6Te3mWBS+qUDXd+JjTzjEZopyoqCU1ZhMa9CUmsthc1EvljflTaYIOjN9YaEL00aNacj+nS3I6Qs
rDFDzuur3T9XUucTckJZDFnAtibplbzM8OZSSRI45raGIDIGSo+WSoYR/xVYR0Sy8dqq3al1OU3t
5iX7YIsdkXEwKB50yHAeRMeC6TB6ssY1ZTUX9HP1vsS54OVHY+AGmHsS9xJsvvOmDsIUsdtKZWw8
R8QWnGAdrLsMw1tWIgRK9UisFHw7fuOMOTQMK9oNgSfUADPZZ+/QYvvzX7lE0jlxEV0YwTAZXUIv
1pnZ1/xmAPtlCCGqP5pocUJKw+tFt55mQwkQR1EIkoLml7MP5TA7rmiqhUzF04CBa3mEiHesMYA6
Zir2W0VuoXmlgsFJx1sJ7Xara7TF/lGP/hJBsYUQPf2HLXG/IsQ5//AGke/DZ4RusArj1yBeCCsb
F1r9hSftmEYyWW5DTIYwLpiQXxuUaJC9+7OG4eOv6sXkpVGwItAadqRZ7tGAF0ygcDiEb9WqNl+q
9G/WHNePrtX5KpqcC1zHjw7EWnHYYFeKalGVGloNWzWPI3I/wWlRxTQzl5zXnkkiGR8bGmiclHhS
RJ07rgwFClCgMUP8pOpeGkffRjd4HSaOthvDQIyNxXsFcpqNGmnwCQzxYzPZvtQkLarYsBx6gGdw
Dyw+8SDMxDBBcNdZSpTIybZPcS7370YyIAA9W0+C5zgQhTj9RVqOmyiJp5h611sV+e/bVuYJzMjq
rXNr32187Uwb07rCpNbLmUGTeCSgT/s1z1KxKuxRfpdZpbOP44YvuM9jyO1Mk1wPwiIbllNWr8lc
jrTTuNoOnruq6n2V/qgGK2VWMdgCxOlJZd2Yl5C5nO+y/MtsFwCP2etbw0GcRNXlFkjlDou6c34L
83uNMpwT873mpNgN62J5zTqwi8ph/I8ybjfR2ldj2Igfb3T5gB5SwV+fEvaGKDvNjR4C0joE+aXT
qB3IeHOyXRN3CsV2Xvr24knIlWm1mwfbxz6DnGvz9XATaEVvxhnG1ASs9lJ3vmXjw3uNbeFoMKBD
yD2q79psQy2Rz7rfIYIO4KiDJgUDvPByRUQKP9pzXT4gdeTAghd0lCEGxrkuaVkGd52ODOpJvoBX
rpBH7aBGaXupJBMYnWzqOApDQZwddEQcCpaPXem0Jq2BDOudjH/UgxFxrOjggwwbdCXNOHWP6yr6
V1bkdHncvb3Wx6um/0K/9cXNw4R5Z6TmnbVwEUotvHbm7cuwjGH4+M4cXUtPvdZzEuKB+c//89ya
pWGm3Nmtc6jTWIUv5MofRNj+v4Sy9NT/prOqo9DH9BB6+pB0nmLd/5J2sQeIVtBit4e/QtuD/AAU
759qlNnycvKrWkISik14DQ/hL/y+upf/1Hbouvx3frxlurvgv54Mmde/v7mk7N0tlYcBASO+g2P6
9oJL1ujqX+HlY10LewqLz0WkV58QAHfN6H6qX66rOeaRCi1y8JDdHZHloNk58OMRlvUWaZW2Dt4s
V7lKBl8Mo+9tNlodHX3rctVweBl0BfWI8ZlJbEnxwZZ40b1tUhpGgWGA46xrTgvwNiUXZsWIn/Xf
IPxsVBueFY9726KmSFmKitFDBbQ4HfUqddFDA4pFqHd9UovMuOlHeX0cBXb5gz/XwKRyyu0WB8cT
4OqQ0tV2UOB5nXmbMkppCMbRc5BFi+BXyy4b0tN8fu4+KZfiC2iFMQyy/+z+Q2G5Uc3ir2yfKLnM
oQhtbxRaaamOCJ8N190J7aIik0qzFyTRg0sWSj6tbSg8B2hyvQGgW9dGmDUqnJqr6+LWE0nO7lQ5
npAqZCOoXQmHhy/s71bSvfPIzWo+Qa6m0PSJJyYbaeThK6WnlMsgHBXKQUlE02fqhjQ0RiLjVrfb
TAVWgv4/TydQJ3O7p46uNQRFpHxQEQHHGNwgOnIuRhjV0F8F6+H6z47+FWD5Aa/aaaVszeP58oLU
9k4Gu/m6HuwTlr4keXVdVLmwHe3cPgXI2qGoUDcRbc4L08ZsrRjpvzKcwMvVPSb9+osblERTl3Ol
jC7BCqmpfmk+1RGBO+SENV9LmPH6SLEBt1lxLI+cVhqdeV536v5wunKm9//eSrD/4UJTioU2s/hX
fVNTdsJb2xZbbP1oHVMrQdynvOkTFloSyxdytxUvHxqxHINk3A11CPseJU/5W2UMjS57+zFH1ll9
Xlk7oV07KAbT7eN6Dvdl/LwHRXokfUKpCSMJ4kKwh9tccpNQhQ9qAP/QxRF0kJXEe5FVTjFa8i2A
Cv9w1SxPAm/amTqvK6C9MBd4VBQ7JBvMY2KFpHF76lULdmiFmlJ2P9f+kgTYXQ+p1AedBm+89wpt
PtJuV4GddUQASXb6yAPEfiCpvAEHd2MC6R/CfDZi/PNq1VD8WlF9L4XJOVSbJIlRWEHC/IrC2rMt
IBgejBf8haSsrwy1YnPDs9HkCMVHUNzV479urBQVjV2R+99yG7FD5v6xdvMhB1AsVVruu5nnIdNy
61wl2Mnvf9hbmg0MHXtwViG3XmLJ+Af1RfLbK8t0VTdfbr+xEmkz31Vf5OjTtljOg4nPSU2YTtMc
xCEQBtpZZII8CeX3v689vrJU/Gs+AcHnPoorTufOTGrG1GZgIHinPXzh5NrKJObKh3yuSdnUJCCC
N0qhcVsN02iEcSbv3iEP+Un2inB6tORt2MJk4IHwV60QJqT1XgccYL+hdGemCz2fNsXcXSo5jAlm
1kvinzJCbO5zCEJUgu99R1nfw/wL0kH/CYkPtf/7YMIfggkKZUULOBj/tZ/oOAH7oro4O/jDAxjt
aasoxVpdamsUt3dnzwcWrnuof0GCZxUGmw6bxerz9yTvhZCPuHcnhlJJtPKkYA6HWprMsxrPV6+i
XgnK3wunGY9MCBmNVHWnnxx3iC86wCBqCTsgutzTt8mQqeYT4DmFXyucNqbe7/VB2wYg76Eaik1d
IA9uOsdA+gozihbQO3fAeMo40jfVapkyX/f4lJuBDWXSZ5+8DtFCPFomDVfzzMe+HyrM0DFM68W+
iRP4BDIYudbPvIYe7pgWYK5532frgZFyIltOX3nfwW88Ip8sTB90sMM45T22FjE4sbZ5tSCv7qm1
pIBecdESIAWz3UZv2/znFURKH03FNJ+Bxqn7o9z2HKG0mYdd08Y8kCS3vNpRjo3EVIttdpvTgqUe
U/0zDfJYE93XcYLonQxi3Yy4dzOF+/3uDiYoabVXa26+7ZkEdY1bT0kIFYJG9WPhfe+pwkq1GXtJ
xnqW+LItu+C+sex67Vsr1wSQbQCD6vq0QaNIPuD7/svqLqe8l8X9C5oP+MaYARGQU7lMARKXomT1
7RUlY4A7RU6jKEN2zq3yivxtcZ/zWOqp+V9cLhKksGc+Y49SXagRTMy1pgvxnAutBzkezFo8VPkf
vI/YDcEXz/NEMuQTJE24i3Flx0Kd3wAI2L7JRt8ISDwszB1KPrVXeGTWd5GnJv8bWSsDjgQsYReD
24NMoQ+1f+rpfsFaR7q90biwSvv977IziaRPsogubWSyTcegBReRlv68mcuJMFWbxKSBdlRn+rHh
SMv5ikALvuSrkpzvnVx/UsqdKv7p4RCdbV2msl+lYpLRAZIbqwNegoWrvpQxCt0c5IGC8YgKiQuG
QdwUnMLAf4a6sVxn9slvYpPDp8n3O5Bh1ALNMrLbhH7Vk/kwrxf5eONLG77YCIiKWh0tmmwFV/7c
VxelYqu1rwUOrjw5cq2Qk0SNGoLMw4Pv9M0WZ0MPHg+Juv6TXsFJd2XkzuSJejr3HuMPLh3ACuW/
gT1RdoY2V8wiPU96Jro0Lgt0JH3+vUnz5E1VuaG2+ikNNR3ggAbMFImzaChQaE8QA8PiM8YwBSSx
UfgDt7wXHYaTbWL3n8Nn5VAAElGEn2VXxArbWyCk9Vh0Vd31wwrvSqrO7vYX/NPxN5eq6n3UoZKU
nRZMW8Kj3UYtYhmJKLLKzG2wIt6yN2fNU+9tmCJO+LDqV6efe1Jzjyrn6dsVmiejEpF2j9cNZOUT
i4HONXG1sap6GXslMx6kwByUvHyJupqZjKF1zEXIDQX3tMgxv7uwREkFifLbgDBLMQJ9YXueZIWJ
HESyHyWNewDM7s9G/pjWBb0q5Gc33e/9Q2xFCDmD4Qn1NlC4RsO0MWpfSOdLHEdetdB2KIMLuLnV
j6K5rr2ACHb4Nfsp9Qnl9eRThrmxrltzw+mGKs7zL0BeMUekH6My8+Km7acxUTpeKFtNGoatEoOz
2z5jx+Uij0QVGYcGPsU3XmWK7y3Gwyxk1weeDsN51gFqY3COiwVr6XuQE3ASlqTG586p7B0NV7IJ
qOFufzm+cWm5r3L/JvvdAAsLAdvWdU9DfFtjTNzyVfLUS9l0vuCiqWbFV2y8Is6BT21unOOSOZuz
pN9huBI8zHQ7koecvUl03V8zU5mOF6jfd/ohgSv5q+M1GdrkgHRARg25OSL/cYAFyzQtMCz3mpl8
Z2WJAJkk8Mc/8EJaCFZByKcZ3vATIO8xYu7v+1axU+SNPXPhyz1r4VPYWjcPCtJiFfnDXh1JR3Kn
RktkA8skQkQAvHYQb3I9wmUJUtXn5xfGHQO0fZiknvMyNefYemyjaOAbMwb3mm97RdytGsRXN0BF
z0sYTv2GDeSpg00VyMXrOMxKBLuouep6XEaioHiATzLq4W6BeHKXmNxJmHI+zQ43IKdKPh0hJv6v
wmQKbqbVOoA49BGW4l0ClNOeRdA3pJga5M++165dqgCgbBSVYmqjzdcX3Ry8GC5thp+aT8BsZh4/
tX5bSbfv0IlEiQ+LIO8wO/vtGnlkEdhAXvIgohrClcXgMDgyPOpc0h5ZhLPGZvT5K4rPWazbTsiE
x8DXu9mtG9hUALtsfIwHMFDdOH/gCmO9JFSHf0HeXC6l8hynI6hkF5VdVdM+puazvjf4k/DWL8oj
9ADtJ+qybGn8+getaGHn0/65gY255iBnG9HAeb8BSgKcnAYm/Bktib21dLyO8Cd83H87UuNDce+G
7lpHKTnxem25So6Jp0uifwSYy5/Y2H7G7jCElSVAq5Sy9mp4t4S07jfMtmHzPO0sqaqhnU4nMAmb
isR35Wt0PPGxhKmE61KECGY7B0axwdbv9SL+Hsi6rM9bkHglWonX11/aRxC6fEwlKILOkgrVkkYk
E4zowK0gXNDHshxlMnrCZdSWtjkYMyvJq4QRu4Bm6erwN8hRtMN8EwK34uaaAgQwRgVI0AMdhcR+
JAaGgTFufVlplwiG1VZDSUhwSlSjOQikAjqXExF3ROvA1DSkbrKHEqPwAg9NUyLlJ9kUOFG+sAeF
zTNMvS/0G4IN7Hcg35ifc/TocH7UmB6WvBtI8osNTsoRIw39v/UinNw0iVci4GKEzK6vXFSb6jtI
1IChitb4sl7lXQw5jje4BhMSBjyWodGAshCymVs1siuSI8/H/mWU89ZBZKBvLjARnvb/3IfNZLLC
hFMmIqX+wzgvDWnUUkTAEErmg1Nq5X7fjYJzc78RRIIwfQzhRLstNLdG2sGsksXwmO1K2vzauISg
NIe/t9evmthmprf3cds4e6SIQSmorSu836wmU2w+u0wOEjh+yRIeEkIqXhWgGfSjr+b9YB6r0OBP
G/EgyODwKoQz/5o8Moz7I1zN+BROgAKv8W7nKfKJ2q0B5QYIg03tNtRvPiuGgKC3i/Ozzc3UD8hX
vgcQdMiOFKHGcnxGjPbcahG7FEkYuERGTS7SkKlDeH0yMxONbmhsKJma8VA3F9WdeWTOOGFViyG2
GzDQMVsmcc6Yu/6dXbRuByKyIW4Oa0VZ/ynOraNnBQyJN2pU0cPwOzNyqhnJ1oRLNE117DOrA+Pt
JLxZlgGU/J+ea3yeGDeMA72Qf1WRPZ+EGYbrOO44LCDeG+lyIZsV+koaGtwA/HCN93684SnhfT+r
XOX79Z1R1K4HxP3rzfIJgWHEMsWmLJruq7jIzC1cWNX2pRAXb4Y57EHgkoSdARBDojnKKFSunctg
y1n1RsbNWMnme7MOwML7qOVqw0Fma04GmeX9+Tvx98fdFiL9HS6iSl6ZoeDsvnDu9FCRiTLUyPit
gBsRw27P2ewG4kg2aNCkk9SgfI0S32A7Nvh6VGxHHiWU6cCNVmCxNLCdJV3wEP7S8wx856y9JQWy
bZ+zVIiPMjSf8a/PxifOmyk9VJdSG97ZVx3iTRayCk4m1vKoTvFEefxANijCC3Z/WhUNNj1IKIhI
U1+EPBn8chPqNF1HVsSFyGLTxINYLkqrsyLBzqM0t6cWHyj3gqo5TMRJmJ9r40hOheuTaTkbaCS6
XfcXRXs2NlOIfNB50wFN3+xr3fbPag3nMhb2AyQL7Zig2PYLUItqFGw/Xjj1z7yNn1CUd3VYT5ZM
TSARVyzsQCb+TH7bF/3QEoC8RaGn7qrFPqW9LHCJrYRVk1Gzayy1EAwt0SZqteZ9elbFS32SSZTy
XgEaKueDVfoMyE0BX/YTIY6UdCo6/PPblqCk4Xe+qceVaGuFhbQ1kCe16lUOPds1SPDXSqWvB+WB
i5GFM1jgn9EmAVyljkXf/nQ52apzv4hoblV03PGeWhUSQmLaSQwOcNXzVtioXzY0d8FxPvp+qT0K
jLA8Sq+vZTx+JMFaOYwnfEQIaCv0K/qfu/RfWxl/Wv1wHDi0GhAXgISqukRkHk9KgX6UWC9c9heG
oo1z/RDt+S6yi71DGXuProonicyytbjnWMbA/3fRtTZl2ZY11YC3hL0Acg8oUIj4PniFYuStsGav
SjXn6+vPkF9hfBBvA+EFVagiMOw0XXq6MW9B6xGL7iWoXHT9HdE8/iGM6++gpsHBZ5k4vjq4fRm2
Bj1V2nQO8jmJbHo3Ad+zfoHMtn3lNDJmIqIL1otg5SzrMUqI1J9EnxnmH1aMYTLAD4cMAHFmSYVX
OVSHT78rfhwgyr7JyIxSeQQZzQGTfTPk3gmMB6Zn5+wtPVMHPBP9XAU+7SGL/+1j0xHvXrQPCdfR
GqYpgd+QDbcEXzJSSDEDVQxmgTvM1smR8p0GoXkHzKgzEQwCKh8l4O8bDsQrFlY4Gq27ZcfTlEel
mPGQEbUmBhNFs59XpvBq+3Um313Wfa8SBCXXnfL4GP7qmM+QZI0iaIGkmEqryEJol3XZ8zabGUSZ
9uz7ksgI6uLBdV0IvTx1G+Mn6Bx21UeczwqEyF8GKkHC8tZjJIPeOSUEWuitkCFA+3Z1/YE9LhW/
WZmsCYucOPjmQL5YzUVIvLLNtO/xPivjl37Ha9NDd8eP/VRh9ktK2jPNKchJPLzO25LBtvmwH5EL
p8pAgQF47I8V55T6E0oI8gR1s4jWDS7oWWfVs9Vp61by2h2i3kZG3YHOfdxvmch6D6+hkJnX5zkw
/uw1qt3iSApI8zQarVHu2B0kfjapFFtneLXnhGDQIPvq6QG+mj4S9hS5hx+OQeC3OhBi4JPKUTvz
v0aAffH7adMx7slbmTmaID9HIAWrGj28W6YeI1NhQS4zQR9Ctb2fxz4xUdEz8yy27RuzJWJP8Ozz
k9vIpGU8DdKlb8MlUd9HZvJCF9oMYWAEh9YfxhOqgjvnAlPZBSN6S694ZjTpR+lD4CQ9uH0F36ZF
2W2iVnxCwTbkyu2JSjQfa8Ay+kRoaUvHQYcyqFtuEcGQuQCXWpqFxdZ1raT+/iBy+PDCmVtb8Ofb
pWrm5mvT650M0n7Z5h+woateUouVdvPCijRxxhiIHTlAZTqkvE6kUU9B+brt7zApjTnpD/o0+WK9
Ah2zjbV9Q5oWVljLy8uyu5QiFrLaAooO4iSwRKYpJgf+JW6miSpC3ELdNu91AwaDa/TtX9lijrDo
Rvh1LdYKaKOWEl5VEHP573np/E5mKLvnj9LsGSu7jMVtfObJ+h9sVov7V1u2gX37k1xyiJZucv2W
jwuDNSnW9rkUKKc4EIrubQpDlx0HEtKeqis0bfDASG2NMvHDDjj2qAkDOMaIQQu/OguEctOAX2zu
0K7cJr81edLhM4yX4kxPCcczRnrGQcz1nln+azxdbeOSI8wId+LUlIM5PFps1lEvx0+IxLj4XYOI
saCAIxRhnVXbUkubmnasCEOzkUKGxcjblep+nSmuEhpCP3IwdHKPGVcPJxJ12mFu7NLTQa8HxAqr
yEFW6ouV5Dh13v1ZmeCoVdg9igjA3RvHjGPOSMT3zgRDzldegCjCQkROPsIW/JzJVq3DhmeTEu2L
q4WYun00HwkA2mfMJpdIz/MOLa9zXTA8XqWLZPtPMD6ZiXvNk/2eim7zVXeRf+udvI6UcF/xtiTp
ejehJaa8bQKszJXM9EPZoPu7RHz3YpHFLwEnp6/xzItoUyH9DawhOEb1reirpabX5JWsvloYnVA8
GmJfXR6mTXRoZXIoKLIsjJmgYUROJEUA+2zTgSvBcpIwDoEiNuau3cG+HFj54OzYWVs7LiFdwQ+V
nQDAmNP0Ft9B1/uq4R+Rwgk7I6N/3TLr6h6nfczcwJQEUa+NlM3fNg9QEOAdKyj2Cw4pWwrQBYvc
TSCQFePa9VisPxRmxUgbPB/0dpzpDmq7ImII/NP+Qp2lN8ojh/BnkqDpLFx1njS+p9sbgc69Ivbc
N8l3yHcc82iPJUGSZRwOHdz8c9tghfODjNsBzFpfuhaHNrSiRCR0YnD7vghEPndNuXishhialPwQ
CGXpgqGE4TsaIpX9TjGkzHd43Z/r056fm8IjyoKYFR3MD8WFaWWHBX3hh9jbfh9Hxmr3DbKNk5fq
MJVGPJGKDjGki6IQhnS8Czbw1opPAYFjHwje0kqyv8kv2+jemJQAvFLnPCePfVj3gwCJU85gITxY
4+Qyf2xI0X1PpNSJMxyKurq3WhjmxtBfUurf6TDkPZnlqtSnQHHbNJ5sn+gYEHnYK8VUVMyhIf7P
qKj3TX/G5aIByNs+lR0uzvdEO5H6/4BTnzKB5MDnFPWFX0gEIw90iX2c2xvfDi1SzJOCFX7OaFos
vk0jvqQuxJPAW1GFwi3ZpWym7CrRJXcxY30xcP28PfIOnotJgr7VTzQZbQesy6kMjKURNF975AN/
ERg1lVsUdEEtFjE50DLLv8na/FGBrVP1CGomypOP9Th3tfZUN4IJYITEaTD1a9tNJDxMKeFivIfy
LB4n4H510iX2bEmthUd4Fj9vPlQtPg+NbXNZJ1bSngTXTf1+dTs1heVWtvVWziAxDkWmxcjNzbEj
GwMqd9jZZEmFmEmTESzVs6Ss9bJESDTqIVbzEjIvgGk2pm+tLefOR2BdeU4dR/jMrPn5BjBlOihJ
VBJ/G/MzMSXZQNeOnxN5+D59TNQGyNYe3QRKIhoL9hIAmgcToxexS51oS92rzwVIGoCr/pl/mTee
8zwYMeU2b6T8pc3Zb7N0LbKTTbl9YYvaPSV/Ro9eliptPIf3/90AYi+JuxJpUmM01viARJky7DRh
tO33heTTbbDSwwm8keuRYjiTt2VS2qv8Qh1gM5SRy3Dz9dYqXtf/z9kDxOxunJe/2UQckLm79Fy/
O0izSfCt8nsOpYinbyCnmpFqXkdMbJJo2JkD493saaIt5C52uLfehhNBNkAeq+Wr9Guxxp0u9tB0
qbe43wS9WtCJKdKa/+1gTPS17c0F140QtxYqp4SAkTfLkkPeN9VEi9WOT+5Lv70OajGqzhmyifT4
49hWqKb+6UfgBgz8/QE2fmceWvGtokQSL4B7qTNUZ3UhSjXDQYMgL9dn+nZPNLxdmnilpT8OAn1d
MP+hrBzxERSM5r8fOe3eT6Eo9qKHHLrLugtljOxxgep8mEZIxOL2JdZlst2QEJ+8QESAhJpf+3q3
8nPSXI0qXBpGVXH8mR8Oi+aniImzM/7lVHVzOGiyTbPkNMbIXYn8LGbp8w6ExLobBrMmWsV6P2fG
4PKDb+xby0KEYpNOV/Lpzhtib/3O1x5Xffw4ga3XMCYIROZw5nRGoFPscsev2J9xPNkPN9XoHrih
aVvA6RO+oQfX3qegq2RuNE2bZDivGf0lRPIlOOn6M677Bf2Lqnz9siQxWRQxKnY/ui926G25m3/v
uiY13g6bxrfjTNUK5WPbmWmrzdv3/LqDRkX5eDIsZZ2VL4RNtH2bL/OAYacd74P2oAo4XtzSjclf
ujibxwhIRWs0M2sjwmmp1uz3yojzEyxTt1L6mBcRjWENMH4xM59XFkiDSDLERyPHWh+e3AnmqsTg
DrH9iq4uX6gdKY2icUp+TPKhynvd+sKx9LNvB/o4vyWeZwdnoDzBqz02Bvns9OP912z4nlOO1ENH
/RfNa6Tn5G70sRqY7NKhigI/8h1VmtyUz6CMm8Op7L+D62oO1n11XyUAW+95krOTpSieV2P7nyKl
9QGbEWvUBOYtvKRJ3bv5xMnADbk4G67xcuRrvF92IHfmTyRVtADMzGc++XUfsmUaVSYH081aJTQD
yyF54ub3K3HBaJFXOf5Tk7RQ83NEgYb0v/T8p+V0e5BlP+PWFiyKkTsBidluY911e0jZClYZoVv/
hWD7Oc6hbFwQdJkxnChA/izhFP+qCq3Bakbu474ROp3J2WAo7r9zHCs03Z7nXvoF4+c3DuG99HPr
8uSJPDCam9DeA3dxU+9WK55EsjMTArJv3k0H1DxQCmiy3nWllHWs+8jLMNikGBdYxdB3PVD4ylsy
n91HIKdJ2sNPC/iwK5BE49uAHNv5wKCQeOAG1DwOvvHlSWIyhA/By9a/CYeqCOhTMDsBzX6EjEaA
L2hRNv9et6FEwBTOYIOzylLfppyAWGVsPBtGSD1E317/uZLZ4ES6YD233KCIGQnaHCI38ye97okQ
ybDRNHjeCUabO3E9AoVKK+oFBbcJ768Prp42u6y9GQqxruzChnh0i/dm0h+DV+Bo05/lO0jzm6ac
fBjd+O3yuGaOZ/qptvdjBAqscPhuTOupsfGkVLT9ETOk4eD0gI0Tvhi8PiOUm35p1iNTkVHRiNvi
tQOV+aFyWoc6pTRxpMp2ehbS4Hr+GzFlzUnBb0bVl8IB6IyWU6jvpSTnb8ncQs/CpW/CU7XxbRLP
RedQPa6rmkS/M+7kAiw4hkM7zQIXxAMAvu/BvJnS/MKr+ubfwtDKO5n8qW+PbtBQGTh3Ck3JAJvo
8xYrs+OJyyFklffhivvps+m1s7VdCZGmbnh2ySGym9wTwxbKF6I9tM83NxL1FpwWy7T8hiUNQTze
fhmajHpMKUiQvZfNBdYEnV1qnFLbvi367SlIZoRzVJ+X7T1p7nzYe1WWNNDU3FXmymbtlunBf9/e
FHVxfGUFbwC7wketT7DRWrDnjVUO+MdUdbPdc4CSuwM4kTFTPsQ7oh8PeQAei8N8kDukku8A0dpf
pL15XCQJXXa2PUg8IcGGxD5FlxI5fCYGIbBSL+TWXIG0W9ezQngnyAa2YZqC1crI5bNJut1eNCt4
MYCd/UCB2YQ4u6FvtNLRJ/9cyxpliSVmwYiEkc59yGIbeTjy+LRdAuGBrjCpvX3R5NvNuRAZcF6r
+3yMQC1kpeGiGvGZZ6vdrmpFlz8F7cjSJrB6SNp0IYG3s6l+x+Q61qnD6U46XEzO0X3REHpBySKP
dIACWeZialpwj8OqQq7sV1r5UFZ0AszWi8cs0Rd2zhBsk4cexA36HQ9E31J9rQHloGucmnuPm/Bb
gg2D3O0yhLaseWljSR+loOifrBtxPxHBi9rCYyFBgDKoIzuH9hH9E+qBwPFg0+zEdk9CbJVcyaXQ
kX/vs2s2xs68srYZkxet4jD/9XteBz2BzvJBKBDDD/1kb8fmYvlvMNOUGvNlob5UjevSp8qgih03
QYJ/UjdpITeTaE5wJ5SDEx69R8sQsqnIsLqPNKGdTahxQsEQDPLrJP+syMcDU17Q1I66BrLBhhbb
dTk6Oa5qxW3MWIYVl2zYXtWUq8i+FDfhF0X+HZka7L98nEBPZ6NN14rUOyPG8ncTiF4sQXiAY6c+
tdo/RlC1HdhkTTWfyH7lIxVsZMWoC39eUNx7H1LJNSryZ0sdfIlnZBktAHQLtkpjZ4Be/+HflxZ6
SwKS9hKtZ4GcLgAhrJ2D+mSEHJCCpOR8thUEDG2J+YINBgg0npdBAiReJDegcJDu3VPeNv9rTcVq
F9KhKwWPxCl8H03qoOx54+ElEkTeqZQeJMa5w9XRe+JBQAV+PQHrShjReilz9KgY+tlEu26UmO2m
RC+CFCkt2Oz3ve7XhojOZnUQTcxXHIGVyqv2KIkaWslqCZh5QLoZgG2t0oLavnN6ZK8Kdw7NApZe
BggGBR0+fvjMBHR6nGTOQu4no5Jokn2VcXNSTwk4P+5k+eY4BfhvCi7/TsibvG/LvGDPTKgluqRA
MNAJ52OR3gUTkVLSLroBoSI8g7cv8Ks+8PKLuz+VmzNTKUgVdVcggE0iwwo/to387cD7tdOlujig
LHTrVAGEEeUmr5C4RZwG6jzIAVBI0iy+o5BnCrknNFyKQMd3tdNYJnWCQwaPD0Ah6Rneo8BLXuEZ
b3wBlU4A4NmDAUYePwAb9smKa/UnUp4qcUE9v6+6Yg/6UsAsaXK0+cmJZtqAhuwHYnZPrZak7u6D
TmA1gFYQiFeTUZlfM+ZVeu1H/xHmXavpV//VpAKMa4+qizNnXZKJ5l6VmalJ41U+/QsItlF2Zxtp
j+Vbe7mvXh5fbIYRF/ooBtry4ev9e+t7JkPuib/gnmBGZEBCY0ueC7j8tSWph+/M3tFnlqpHLQtx
ZVpoc4/Ot7wneqFKOjh74wrf7znZBMCmc+AU2T8AyqQIVbnxaBCg4CnmTmdBiV4c6iWPloug867v
7Kkq2VPj3tBc7E6A3+O9t54EzF1JmblrCVxlliudk2rvjhRpoB9LByfXCUT/CjVBMxpH21MfFQ8f
lhbp0lxsERudjZQRAzv1wFRIXRPnXS0eraaV/btSvixAfPr5Dr9QruLUNatkIJWPudFVddvEpIl0
iF3PpvpLY6Y+dBceMEw0X+ljn+dE5d2boCFYyCevbJLOcLfWNQKKC2lB06Skwz4vqgUpoKrl2cA6
p2Mz7c4gJInyRtmuPikY9bZGvNHlu7jcyyNz7LBKXz3Nst/9wnIUXvjNs1Oj1eZqoNGK7jTvz82J
ra+iTmXspz5AAodNocXDCvtuUqPmMj4T1Re9spkDI7e//kTZSKQVkgW7zxSrU880yFC5hZ8TWbrC
Mj0O0q/JQtqSoyeCVF6Ut9koP+Ae+QCX6fPdU2uTxJD+PQxHl3p1a+m2PEdqjAC8yDcqtvLxB3BX
DpYWjQFZAhMy7uitmwbGSQwcEloyIwhfI3r1xMDjcfBr35c5E5TKK2QS/V4c4y138N5ve4NmeKKm
L6IPLgC6T1FNgLeR+v+d2v+/dhs41wYeTLxIuHGoJck4qQdVBJQBHBJnank9EBRRC7Gp3g7IVoyS
XxwMODVR660lzzNFo2hBbAq7n2EX4IOokhjhzW2SQAW9apayXguxODO5a4KU+Q3uPZ0dN/Ao+s3n
ZUq2LPiNuTD6/9PVl/Aaoql3uMeArqT5+WY41afi6at8cclqM/UTws+KH+bk7o8bMjPncvfjs2w5
NwpCg6XLgUFlZeeDkHCg3vzkd3LMtH88LOtBARHeAST24++wTYz/uXZWoW/1HUTN6JTrThIZP6Ie
GsIFIbYrW9UmYnJH+und9te3JVYPvA6ZTRp8d2L4/FeMQI9hyO+ArIjC8+rMA60D3GwzdW5yYn4/
fOpSxI7mLM51SRQiRjxUCrN/jV7cwF7MuQvdCwnh/2WVeKc4GT+lAuAjZfh0GaQzKZtgz5wPKRlA
KPYiM/Y0RcbYrg8Sbr4jcM7UWijiPnM0F0UUONQVqd7J2aEcsJpVrxy9IdIjhVy+ja4xk0dIF3zj
4kgRNsQcImiWYI8QLBeF9HGn/q+eSqzNfYRko+5G1oLXt+G7tzaecZMeGK/ePy0J/j30BQmd6iiO
h6JAuwXc+KJRZYT3i0bryxnhhFBbD4M3WQ2SAnTGIl8aBg8e7sgLGTWtyTPs8HX7crfZZlgPfqQ6
miq+JcWv6NwW1WspWKBSIXtydBZ9Klar7X+bVjb3vGTwHr52aFhHQiMB3itEApXqiyFtXl5a3LZu
b6DIR31k2YwqFMWSdDgM0yZCiZaDeHyT2F0wENB5ZQmDHwKoObjstPQw6lkpBuVA4PJbNT/wNZQc
H326vhfTy+h+ynzvy3WF/WX6B2WR3DrQ1pzhPM/u7wwuMScl7ks11O0Wvfpvt2sNj//WhKwHUAvk
rMOSAC1zno771AScaobvkatknqZTPmxZvo0+1JK2hVlPvQvbhkzhV6i5fZfqTH2fljez0NMqrVOm
FmVEjHuSG1QvTmgJsgQSzyNqs7cYI8gXlhhicErveuRh2l486jfr/hzXxmbmzcqLqGR93tOcaDHV
vHyGr6kqIvvOVJLJ4NVwbWjIFZhb59hTfzQiveKi1dN4t6ZlyZIoU8Jn77LgeICV+2bKy+FUx2x4
3h8jrJEFYPVwvLdEaXZreD1HgKFZlXmX08YQCdRyt9LGORQEsIjzyNZOadm4L294/t6/aiTC5sS1
khEFdIOerS/enCdevrbMUgUd5HVw2+hdM32hBXJ9mBX3YaUkkVi+lHQhxFzE9j1ow871yx4bvesG
4LjHqoygUlty0la7t4in6N4YP3d8JjmHf6ip6LFBwY5Jel1YqrlSxXuJ6zLuxTyLtzGOYcH7egLk
Y1bLCUkE2DEAyEXac5lOTcmwK3TYG6Y54gnb9RkNvpM/yMG+ZWEli69kzNRY+GnqG7DW0aam44JN
2V8QwXBB/4FrWm3i6pwTGCTB8x1RBMiA/PChWKGqFr1YulZKPmgYtisVQk7bN70rE++J3rwEnp/b
RBU8Mt2eR8xeGBUqCSPyMXNK0OBBmyHHMMVbRDYflT+o4eLHRL6urVnmqGp2f+UzrD82ctOID//a
ZcGhUWeFDZWG9L0e3e1UY45sNUtrhnOnQrfomuj/yZOVv6MDkKnTtuYZODUjOstopuvkweorp8t+
4/85UTV4y6BSjI+x38IHZ9lMzcXsh5xYMpv89jabw+v1hynk5QCmLtycMsD0CZW9S+IQg8auhqWE
1jQd0dAm+w1CZiYY0Bbde+e0+v0maAqh/Z714hyhhxfyroSJspSz27QgSXyYUUbvdQVcF/BqDba4
PiJewFyqw9J9VyWRPDWXm4twrYu0AYmv0d9bp5IO3O1KGyNTpbHSBM0Z09Fwz/J4NJTML7lOTr7A
2gkT/2/8+HjHyQ73+vq4VeYmS6cWv0ENBNUFPmdtbBjyu4TNrtCyOi29ymLLfzTuhd3Wm2jY8H70
w0anLdJA97WyFXvihfQYllTFhGJ+QFY8E9yBDLXS/6hjfW90Orpewr22E+SY01cMYDM3lXOyiV5I
LEz8qeBnu8k7MCY2tgkH/1y/WjZ30SdR0S6g+M+eCIN845c4HdUdv3c9AGJ67qLDp6gnBZ8jIieG
i06y9S2xxig0IJ42gfDhtxQOSp0cEADCN7gOEMll2Fav4MGJLmp7ax20hHNt2ESYbtuUde1fXdcf
4DUw2BDnsSQa4EnmKSqwPvOMvA+DP8JIMLjCqlSNTXWCIoe5Xjxv6WBlgKVWme7I0I6h38uHGbKU
xgJ4ZZMr29lmz3veW9HqP0HJvbMUg/Vu87MkLUuKjfJiEHqBWpPOfqCq1+pK91dD5Ac2IWvSRCAS
LmwpsoODodwbgZ4fc0z2Q6j6hVaJhj2d+RrHlLU7XabY2N8S1UFeIheU2v64+CmnMsd6v0ZLVojj
8pDQYk+4SVIjP1/TrJupKumA9zTYmbxRF2Hz8hUivwnlw13oBrle3UrjpXHN3LVxy84YvOnfJeGn
Qwaf5ix6UWd6IvNzlRO+FLYV0KSflOVvvGsPSpLemeLV2aWLq2VLxoFN01hQfWvc7AldvVL6MCem
flHsKpKV6UWXXKHjN4TUDsJSVPW/aU2XynwZ+2SZCvgYKdJGDu5Zwuz3oAEBVBKyE9ZQu1nwZV/Y
bsKLmzBijVflnNIw2knpTo8l2wnDbYcAbkLClmc58Z1SNM+6tbCUN6RFXdoFI91iAq8Ro80uGVMk
jZnHRqtj+LxDJeDGgL2brnXARLOPgmMRzzs3m+jnTGtYcYDIEXBt/3O89tpJDohbn614zWYnyURH
5CiNXv4P3gK6JalxCSq0hlCf/YV2JbRG2B6wJcGeSSKw6ervH1YhVTv8uZyaOhVhpCrHua9MynLL
uArICGpagvrOdEU5jM3RvjmbeHt+EGSDRjqhSw/Pv0YfhnE7KSPFpmavALfYAB34QvJkpVcfBZWR
liZ8CUS4hViMqaVwc+J/4jBltcVWPB6Gg9qa0eiifqNpyqThh+suw37+GxVDnQl+wOAvz3dVQvX6
k4h9cw5WcvwOnDP+viuEoYtnr76qxlBpW2qzv3Ct+rHqPtVQGrKGPlAnVK/Gh5QeXU74d3Q/uazn
/Io5Tm64EB4jV6Nd81BhOFSpem5Ee3Rt7UgzwVaVNPGBJqY0/cE7hOACMwAzS/gkZJZIaxNyq7mA
PKRBbeUj7O3Ljj2InVnMnCnStb1+pdOeBiyBBa4gAtsYewPdBDkm9/kx/GrFWZsXuVSXxLbsesXu
c3fwuXaujtom08oI/skvTj9IU4Mw1FtAXT7Wv9zfrmk/tguODdrc1sRoNRxkgfSw3Os/+zCKo9h7
H3jpANVvzISg9nxzaAoIojMy4kQgKj0aXF5O2LqNl65pssPg38DNxhY5gT8AgmEfLCb5lvB9a2vT
wwD6OE/ZgDr5ciJy9htgMpHMfTcn6ggKYwWGvzeZbGfB+Ej20DYu/9E2EAPsFmt7MFaF+gER2ZG4
QvGUKXGc2Z5sJ8sUAMaeaZZV0yRmyvJtbMeJT3C7H4pwCzwwm89jMRab6t4e1ST+zXQTjXuyaNV2
z83Gn5g9kNAIosC5xfnkdQIWraLlrfOtEkoyTikKXXh1/hK0ZBtGkTiKsrXPc5vfxUYvJ0d2ZH/a
FrUBxAewDtkSye3lnMlDMtFLr7Trwb472W2MVYOep/fW+JnK2j0xi2DLFe32Y1sUhvGulscuAX9O
mEqLBc9v3fHMkiQyFzE12J39DPIlsSE4vjd3sRr4Cg73LPjBMPzA4JSlEEQpxArMsGepqVdI+2hS
re8fVVNoS3p82SgjZp+uBo3CdECy72SQYx9bMJ+ghOlGd10t1R+TUFQ1sSL3Juc/oZRnxfmryGH5
mrA8eokWPtD2g7jr3UnBeOr2Xtmks5mdOrxEzi9XJx+RZxeLEFVGe0SISAxiMEQhwhiN6hI9xQGr
+W4ohyfcgP3Pt0yCla9Kz7vPL56l/U/InS+Rhte8WNYSiQq0jJriIX7GZ0AmPKzaCGuwL0nO4H6V
lK6OnDYtmTehqo+OKYILckEXYJy6J/aDhNQE9fj2e8a7Pq85iaB0hxopBdvOy5O5euoBGC/FvLq3
P8G6I3XD2E6HiRO8Mf87Ta+g9t1EGheuicuaf4/QoGQCWHN5CcjFOuhf5ZTovW7LWWtZXpRBYMFF
cU+116VMzCePRfYjS0o1rYqrOmz07nEEAKqxpeN2UAoOpC+BM33p6uoFzptpBTKA4SORbyoohoy5
z7XnlAb/VxpG8BVcNwysrJ9+PcvIT4M6hLiOyqJRBlbq4W6z8iKS0HSh7ybJmtDnNLOEtjZ2fhYC
HlS+Xry5nclOyWYIa8Kn3/kE7nIc7jJAU1ZLUFgQytFKMbitY+sBv21Mvj6PyXPEV/o0m+ts0UOr
MtfTbsnmyLZ2MCcZW8WFaPBhIyGY9NoE6xg8yuHls5Rb9rsEYdimX5YPBOla1aAotR+BFqjyc/Ny
u108DyA4Qh4RzwNH6Z783Fm/IOJWhZoZpJhAl/7kg7z3UTYwVD8vST2yYP2KnovzT6XHjH4wuhX7
BETfcRepW00JqwsUtkV+g8ymxewWKfeP21pSB0ys+3vbSFT8FmSDHcJ8xKYiGsZOsTuUsbe4/pc7
U6GGcCLBkHGmDMu0vqA7VeFjYZIwRabuZ0VnmvGHzdx5vStrNybfS/G+19WghBaOTbDMe9CuLeYn
wndHXaT/o1QHDtDjN26Vjz0MOuZy3nJGgQLnhnjTff4+Dri1h4QP5NyQYxzzLCJWm3PeLpMgjCWs
PQsBLsrOvk+yQUJikU6cUjUN7Iy3gb78mcMUQU9bnQYW7F2cDdjl6VrgG1HBKl3Re8eBnWGWhfcj
ac14Ib1d+puQZUYkS9GCwrAwG198h3KW8S4jRfz81v5rcVcuftCIhlEWNGiX7A1DLLzlmNN2mXir
ozWGr13Wtu5oN7o20RNjo9zoHxEwq8Ez3mqNQWtDykFKnEMjwU4ZgJXTtep4O/dGztNE260BJnlx
rtyxwtesoseydn4+4pZTldkC+USvwwetCgz+/Q2g1PSfdLd/oAFi4FKzk5FbWEXNtBzNdjifSA4i
aKtXoc6XCRHNtn2pDTXWZinK30rADScqDTQHsMELwxF3fMPCsY3MVo8sLDC2g/CpfK2LiV2lp0pF
waGNvS8wFBEFAzvaDuax9CcSK74DEO5UZWMZmWcR4qnazxjbVsVbRHN1eKXW0cRprA+QGVYh51iT
iEO1DMNiw3iMp7sfJJNxKpinUb932ltkK6x06QRzzZAAKMoqzPmTv0jumCsiI4juCk/NJvLuYr1E
GsTVa2MimDtnOxLlBrep+nX1DB9YsPznx2c6vFitIo5LTFM9WanJQd50SkjHnrnwup+feGH/Lu33
oEsJXx+hX5gGJUtiMgFfkNBI4yhL5y5MpEcOYrOXfSnFJtfX3wDSgNkuDtyBgikcuITD1zjRiXRW
1Re0JwYbV47S8oYZCdtG+knzpShYrJetj/VdBI+v4QkypW8CMXtZByNb9Bu1UtzRAIyRb3esvSsH
Q2PHewPhFaGoi4NBi/E9bQ55MKN20QT7ss5YOZ4TCBmlTz9DbrBj9KRn8XmXt/dtC1s7OdluCJ/n
Xh3Us6H6qpTXC7EFF0q3U7wlue4ENYFFxmPW8FcPxqJFiatlnaaoI9iWOUKoN1hmwleUb5WpMfsS
RZkKunjcOhCIx6k/dSRcXV4DXQuhVtc2ieAaOQCyi+ALDCRgpCNX/BKJZnZOgKTGPXr4U7WGBdbT
4xV7agAuJ1DBn+AiKBmoJGeR6twoK2KkFYulTH/bMGV0IeN/bt4dB48jiVc6SAQeL5EBmXeL4czi
VbtqwDs/tEH58AC1KnkSJPws56QaelsS/Qrppn5w5+48oH7dRLUFnHI7Q9FsTwbzQV3yJi0Q2jQy
8O5iAGxHZ28nJECe5j/le45EJ2imbHEAbCKlGx5s7vjYn+7rC+e53Kg8Ovz5ZLKzfoX5QTRKJSup
b0WLbiHrPOtIm05GGifuX45Me2RO0ZXnc40trkgfeTkpk/4BaXkMbtNpOunIpcWE1elipbxYL3f5
4KCC3J/PxwCODxP4EJkfLDROWsYgwPEB76RrEKcyM4hTQJnPTFSCEfxn8fd3UcTr23a8OUWRxezw
6uTeoi0fOvE+MkqK+0Tc/hJcSUqiS1a5M7AJSwadwwf2d9XCES8Mmp4ItEnly90Bh5oCmh48LC5y
dUW/c0ZGiqXIVz0uMP0CVmuCP6iv3KfA5VYs1hXaSBabJVYN0PqF4jTvSVud3IXk5R4egoNo5V7e
3pm5hhLP2usD8NzEp7iRSfjqg6YHZJwr6ds8f1/D5of+BQxPYbY1xiYJhGNGTDBiM0XJ5O51nR1D
bH7nG4eaED0cImFWIS/NZlixHfsHcASeAQ0SWOWZIh6lU7tplJPUjr985+BzgPrGuWQjoRF4Deit
Gm3O8LH+XR6XTXDfnEpmLyNObyOR3WiYJwt5PFwWoOz3DG3t4s98Lnz7atlUwXqE5UIFNrJL/+H1
As34LspGiWwhHViRptPjSpD0JrKIyFFg6svk0Htf2AgKLB6T+WucoSxTHC8UmWwdcQiN5haNInxj
E8rtDltUKMTHjEUenZ0AirU1NnY3z5h4LPHtJEnHYBSWdK4mTPJil6vOiETSc43ztfrGqlbGMbXO
PFYUSAqhQCqzr07W1cCS8h4gbSXdnvjNjGuQZlw65dC/T7+lvSSBJ/fpFne2IyHG4Hi2JtZ3aClQ
3w4/MfJZANyLig65/v8qU72Q127ya2p4q6dPtt6VE6+DLUNGZ2CVZO0JUOpPutRv9ZA4lVr9nptG
yKMaInsZih3Qi3+hjg/lD1OUo9CDDR9zs9PgI1aiby6lpnTHjB4EjQN+jX4fcEM1cAcLBWMNNrhZ
XhCGUl+9iHqx9fVczijjzLWvRy5dZF4vFp5RzOeN13sikEq+NmrVeSKHKKkWXhr4BYCD4P5a1fGx
1sKP46kK+hLzrcY/WP3Pkh9t9CTxsPvJrISpcwPcYyd0e0BlAxTu37jZdrkp6Wzg8jEKqpjqvWSz
9U2QvAyumiCU87CCy3nCS7UY4W7HM9GPZEbS5R7qn3oaTS/A1xxU3Ix6iNJA89NOT9lncfhAhdIS
ki3IY1uny6tv9NWMlwl2vzPUx7JFXVyxUchC7noLFGcF/174oFHDREKXbNGGdua2HAlsFaZzP4fz
F7Qti5nOvAP5RTJ7C7XwjVlHBk9BJEXNRQQhi9iEBPzLqtP8coHOox1suQTAZo7JSkROglMLMBX8
9unCh8eXu7UQM+b8tWgLQlhoW+4+mLzFDzXIO+M4pFY1T9sC03CBgF2UiMkNNR9/2GEgvzK/0e6/
YFJ7mmnIF2ldQcXp2bn206PVQXubffD81MIooXrFgfOsjXZi84zw3dWgWFBnLjsKrzHfIh883I51
4inTY1/mvi2wQ0TnMAPsctIi7CFjcJMXvw9moVNwEXC6qwxrNuhmWfORD/WEwaIH/Kwh6wVOe5jY
b8tNhVkoRACMRC1WeZxIc32SgACcovSTbJzDSDEzvkD+GSnI9+dwHGINvNPtUDmpDbXxiHxcCWZU
IFLQpzBBPzK689003lNXlJexUblGh9XE+ujIdNi4N3ay8T7JWH0TRpOt/IK+uVo06W8v2J05USyM
ComaP6iBQwNkYtazwbMEHOcqnlaAcLf7SQQ/9yEbTI1vgRfopz+lDHOLQAnd/C6podxzd99eaRWu
TN8HeGk/5XM8VCCXPth6iwpHftusSqPBNgcu3MwtkN1gfGNGqgDw5BhMn+otd7nOIfAkSXojjT7k
foAEP0jBgsjm5nHgKSpTXEds0/5xnKZ67WcG31iHgiM1ZTFaI5w9dxvVBifTrQGHYlHWA8X4VaEh
h0IIZ0k5Gb5DTsylxphCh8c6TuGRCTAbSM/z3wQymG9Woi3lBwD9TERhoBTVor1lBHuIblTNoSG5
ahdfKGG6KGH3eelc58E3z3+Jsbdn5Qlwq47D4qXgwu/M3Ekyfx2m5Z5XtZMq/5NH/vhFt3ltH2Id
NPSUmy4oN+BHnitZ9aPWN7+zyVxy1sxSiweMqe2wM/hq3ewFgNdBXMb/TI+Tyk+0xIpZfE3X4TPq
O7HaDvpxvtDj+kuemJ2P3G5yScMkqQL4OmXHITTNzQLKtVLuF+TmPr+8SKszsiBHEY3XdAvG0p1F
0//ImnOkSVXhrxipxonh//pItSjWyDauMQ9Bh8SRlZwhL3Li5XOK3QuouADjOKpc2QuA65RuUJQk
CWxfh1NjiBaIPF6GrHjosz7H1yDSqtCa7okk8eAocF2x2wHEaO6WrmDvbrY8fGfN4CbbpxCBKADt
WU6gHEuANzc484K5KtzJjgz6JK55QOoHqq3Y/J6yyAsfOXAT/LpFCrEVCkUcaBbLF+799VnI3A4t
XEAeGAmb8JwcKSR/EO1Coj3OfcJAF+KuwvhUdBf9h7P+k1/J8Jz/KwAKuQE1qxXV472KTr0agxlr
lTXzgcmtloJVJhPeARUZhsPUjLs56PPL2KAwvhY29f4F+oWSjJ/vLV0Z/vTGomACPXodMTRqrVfJ
f2NdzOm2nt5Qsa/gwZPGdG20Mj2e1fCP9CpWOqhWORHPpL0Pxb+PhO5Wo5GDkJ1FT/KTIz919Srr
gr9nCK/h9bFLwHjBkc1s1Eqkgv6T1+UD0wzH4IJubR1wg7yflXoHzD43HuIYI8ZnnhzgzTrCZtW9
IYka1GqbB0y6PG30tjwitckWxP4GVNy2oGrRhvKkU1SU561iCvV7Vuv6xs406nzCawou6/8Nyeen
ViKfdRIVvlW2Pt1BF3YL+RdmEHEH3qdTiz8A6iMh9np+gy0EaSPvduXY8GGh1TdV+TaZ/Zh0HhP0
JVyEqcJwjIUzlPYKtZ9abq6l52tXM5TSK5iuBWr93VvQXxtKB+6a4Q525UdeWrHW6j0PaNElL2ad
wCxJ7iBMEl9MkKA4nQ5HokgYVVTPBvhRpjZ/DM0MgIwVUDf+c+dpX5s/KAIMxUVJAHQYsnxt2XtU
qk3L3tX3LqCTVhMGeoUreL0l2qJPaBCHuvt4+5rWrEurew3Wt8iY9kg+7YFfVLaxlOy1eY0VTelF
T7pEsccwZzUM2LWkaKx7hPISDLL7ipNlZNjyxe/n+RSD4gUPLBhF8PSTFB2cw4WrjuydUHMO7Pja
MxQ8HVCjg8l/4+SMMely8TwEIo2QCt2o9f+9P30/1PpR4R8823IhU/RLdtTm+qG/lmwWsv2cb4wu
eGKH4Q0bIyF2kYJ2cyOHEYEKpeW5Yuze3D4zNizmB1bsWysyTom3VOl2Oylq8+80FBTNB0dxyLAZ
hGmJKg8mPxEmCB9sUTOqomsq09FoGMua4Gt6vxlTXxwGpgfKJY5BURINdUuMmYyuLAHTedmr2W9J
FeIuNOIIbZ7GKiI7QZUaIYo0bT5M5XV2SyvFnm8SNd/xx6bACU1w2MaJmSLKgReaDFvNBo0wOOwj
618sQPAkhXeXMLNfKgqDb8Ax/SDBqZ7JfB+NalLF54htsVk/PkE5HM4Uczd32Zw0WzkdUgUdZ4fy
UN9VHTf2eK619tfbiiDq3ZOp4JLn7yZS5RIDzzxQ7Xi41wgWHqeVp/sEJYsFOmmPr8q68ExBSBD3
O7XTpyoJhF3Fh0U7dkN2o5nOQ+lTsqSlRRm7qzt8GIU/VybEiQDngrqwBlB2pEY5Oo/uB8bPxxui
e1mxQJE5SlKSVjbtHtrmyi/yr/oisx9OopxE1gB1oC3f8oKO673VkJnP/ORvlOIkexWrt2XgDmWs
6sDu6AeFjdTPLKUHOqy2YPgDd95HfPxflMyi7JBVNiT/JRilg09PAl/gZkrie+pJwmzqG0WI9fRq
nplewVCyzKKZ7tAWZP1cyy/arSUhi7BeK7G1qLyKIXpegGdc5HtU9Wr1cK3XY16MtuWL8rOqXpdv
+tOyYWs8btBNKvJh0cGUb1eDTb2GzL3K1JAP3osgF+vgedgphHTLTpBrbk2SNx+jZQ6WYeCWUSn8
DDltBzUQcf/nQdHPHYdJuJO/YJqzYaZQwOahWrYveb9lfAiGGQDHSHAsJnn8cxK+rKcOQ7gwxW9B
emSVI5za+VUR8A8W+Z/GM+Gr9VrwsXTZT6Iuvwl0LwKo54cj4Oi7LtjIUeg9QerhZgSUi01zSqqZ
JtscFonDhc3TzN+O1NgynusuNd0gUcEWDOI56ye4G87vpLMw/q553TvIBYkU6+vVqxrIaq8cLEfm
MxIsIqF4RTw1dVmN5wxanmG8q+rJSs0nVxQw0Yj9stXFv+U6HYvo0vEcK3M2QKfo84e/L9AW2rne
fkBWv6BEzW0IssMCxcPkAi2mVsqLJ2KQebrk49Bbmwv+ARqbWm2l8uVguGSvt8+GBJ4768GN+plX
c3xaZJh91v8KD6XyimgvUXVgCCnjJNuQLQr+K56HDDvst/sCNfa/49cUO+3SPO9TWzf6uHfqkEbf
0UMzIpQQ3JP/4Q+5Wn6u516QmqGB8GZZlUdt1/bM391H7nbfbGIvbG6KnVyYGFfw8hArmUQvAzXM
A2zElqTf+HJ4yJXeud0xcF6mMQRa2U1zsvRUwtA6KLn2ONoRdz0yrb6UeApWdWFb3jhv8Hdu3JbN
8N4AztLfcKLenZhJcMQXKPaYEzaJVJpUM3ZnR9QnldakADyJpv+N6G8T1l/bBnD4dFxA4vyZMmsp
+n05PcLxjw34iZIJAisTj9JMqITTPlyACHn2TwpFaBMHDM+cl8tl8Hu4oplphVzaIVmlhBCVM/Ur
ticfVGgxPdVS8+YtrvCKdX8K4CCOgYyADwIqwjPGwRU1wzhoLXci5AajHHMQKv1VILBymkfoeoh+
Rmb3axpdW8BmluFRVJtUyWfIM218z99xLJLJF3EmKZKS7mJIkzOAOLz76oOS5K3mPty6eeO4sUZG
xbwpbKyYOkt4GRsWXCu+UyMPMCpZQgJ7fHuNwLZC7Fn9xiVrMB6xsq0Z+EnJ4ChwgAzHnM/w7gFR
7SBSQ9lYDTe1X9fPeaoue3nTv4fHngP3ShWgXgWQx4HlmVvJZ+LVyFlT7Zw2EyM75nHZN/BRtu+S
GPEH88myrg33mZbD8mx/+DGeBbPwkyoI30Bi4bDbOKmk/QnJc3tS4TVkWUT9XzwF+P4d+VN2WwLH
ZuctnwuP4V5lK7UWS3TfVuRp0L5aCFuEwD7t4PJel7a5ZtLc+RpltFtLa/sW0Ilq7uA9Ax3F8gSy
gte568OxbQk+99aWhbfI7dFYxfNTHo3y/cst7iXfImIj7UpuONvL8h+B1qLxl5DxpTjkS5ugYE5w
/pMBklDD7b1t7610q3rUkuKPqJ9DvN2JxgNkFng7tXYoQpyCEhZ6iRSbdeytyUGLnux/sjHzO5xy
ChYFEebJq/Zf/zC3diGQam3hbHnKsA/FO0FZV1wgQ+zisUuy9UOtKf0nA1c/KdfkejEl2lPfqRCd
oAHwZ/ID3a5SMGNp8qhqRXx6ea/gbw2dYmGvo2352pjfsKGyBz7F9815d5rswVubPnZpLpajowvN
KMSgkenHEbRLu2DzPGkGCGWwGRsViA0C1dR+sEeHAqpK+E+cKOwMMSapfVO/CJ64WvbsT4ZIgKlp
KbzY7lNQ5pWsNpPdaKhd7ySUM1g3ld1uGGHNL8fH7ZCG3VbCIJgLqAdtSNXDcg0Oa0vawSo6eN7D
SwqpH06EkhqPqprUy2tyFM+1AlaLe/rCCbqXUiZgB2I0byZhYDEJkcOkgDl8Yz/1PsA5fa73r7lA
pmdWhIV365h5m5p/yOkVkOtBL58Rtin1uQmrLajMvd/MMrS8hRr56IGMyc41RS0IBs59Q9o/0WZL
6VDAhW1cNKX+A4Zfd6PKD04/qaPKVFD7jZ/qHOpz0J3WDt08aZdv+l5cDQve6dwPBU50MTqQL7Vz
uHQ4E+86tlzchvgCx3GIDEYxi2pv7nHDS/vmzEDEjifvv7A8XEyytYadwhAZjVUjbfjD5PFUnuO/
cjgyD2D2Ai/YeivK82KgYVyqOmspAiqXUrijCNjAFt9QW9Ghv4sL9QojskpxVnutag3acAfgzZiX
VciBprtes3FJjKjqedNTFXqXJ6W+3hSb8hVpBpOViCcXdrJc46UL/dnD5PWzI2wVrPvCcgo6CstX
m0PWpny8BLCRBRNTUWZwQme9HBpJAJ+rKVq5BxpRHJXk7L8YD7hZEEbPjngqBUyixrkif8bsJYrh
U59nADx2iOGiSiONMO74/gujFkYgserOkoTi4Th759oidjn1v/HN0ZEHvMILAVV3A2y8MTuLyV3h
l8KNqiZ5hcrPgPV0QisUMXAg1m3rU0z69ouwayfQyvIJG0cAs4p+5UB3YFMMY7WqcUPxfgwcttlO
L9sVZhTS+StDybll+/oPlDUityRIIbvD0zm3G7N/GwOsHaC1VqYPI1/JGiGvEs+/UDI19Vi82T9P
0guWzaj6wGVllFF/D7rOShVO/FYa3euhLCaVklAgpwKXuFN5rvUAuGFH+gi16dApbcCCpkZkal53
x5dANLYdh7oWQWer44m+rZNXeWLkjSmWLBr+XozcPPkE9FPOx9Xc+4WbZkjU72S3IC74Z3NJO6Nl
lOrSrdvmSPvacXQbKQc+oebX9CS4KrN8uY4g+jeoH9zZ715Ctb3qauoI2tP5bZKtzb173eo4Hpzn
OSkO8hWAyn54q7AxEhRTl4NpFxJVSeeHlXKMtCf6INWhWzzC8L++xJWUfG/PBFdSwtbbMiqnT6lO
Ks5995p+4Xq6lSdoVNdFQ0Rq8tmPvlcqnwdEBGH7L4DSGRCSZLhEDseEiEFU3fkD3LJGLsUOkfVf
SqlHG1yHwnkxCogtAt/9cJrLxBHQ6hivol5dhX/aXFhDt7Jdbc4AYWIFQ2as48l3RXUqcQwxb/Ix
MkrvsI4nTv4NJFik65nW2vR1r0tw4y0/I5o/W1HKUJ7JPipgbeZMGyY6AICF0fuJ1m0YCskOymHS
E5TC22/QmIbXjqrPzUgb5QLOI5d7B9sNcP86Exipmu+qyKU5UqxZPGNHXXR1A6iNywdhEl32PFD6
w8Cmo8FcHdwlyegVES/DFIpI7EuW2wgQghsQk+W4tsm9Wq6XZX7JiDdiZv0Wlb+vECGht6+ynHYJ
j6cQ77R2pGdRP8zvCdPLty8+iFYMtvYGOLiIxpoDDLuTLBPtUKFxxSU4GxcijaFHjuVI0mCGTT1D
NIv3m/NtamY0a98IDEgvywdr32cuGVsop5jdOzHIZ9Tjm+EyrxF5DYmZOMXPgPdThvNefuEX1U5q
Ipz6sS1Gmt1x5gWiY1dgp4C/L4p1PfhusCtnvuVJUKELYCHdraJ53f1/pWzLql/r3Pm8IuuDFMw7
WkFj64fDH0niaqPlhFnFTobHW6JTN8pxu9n4ps1jYEsaHCH7yh3xjrJsKFSPQYp5oMpXAjag8aib
EhI0m901XbaGzdDW8HJYt5CnuNblVGLTKGSO7JrmCYSomfcl76SN2VX2mjeEA5nQxzJpHh1PiYnj
cwyc0+cF8Oi+ZQwDuUM+yb0UWlRtV2Ga2Gujb1M9KmUR2f8UhNUOrH5Ifv/oh2H50Er7/smK757S
42o92diOLARO2gi7efh6s4si1OPvHFvoYEp7XRbZJcZc1aovUceIONTzJ9FjbPzwmZnKfzw95t2H
NSqKr3rJAf7mVVnBY//ugEham38PddmTFFn4Mtq15kuARla0Z6hizLZvuE5a7jjVOwEVWVO6fxDe
6pCmBh3Hc+0eRx1HMAif501mRqNqi+McjmPpCnZUs9j7Xwmdy1bPzjoHtu/hPZmdBSc8Jk2pxMuF
R2Bd9jXhT17bYy9OA8MYncEMnFx9GM+GqXmrf4Majz3oqakPdzk7caJ6uPfCE58DvNRl0Ev4QNzk
FIHIQ3JISTOxDkwJiqVP+sd8NKnPsWCZUd6CVw1wRvCHriaZWxI+0eH8VK3qQ/DQEdT46aRE3f79
WkjI95mw1txnoJVfITBW5RYsiiFC0ElEdF3S5bF8gR5xwWj/xVP4aEE0JFULpJCUnHN+c0FM2xRa
aievCBZtr8I/CT8ZRCrzMEY9UyoyEo89PkMg2b8YZU78ex/11dQNwrAVC0Qy3OofUU6/8eyFaBTw
j5wJgAdErapyFTkB9jHTxKF5wufTegSp+HBykgqEkn+w+5zWP4GWJys58aNl5lQV3od8f7ypTp6M
BQ1X54IBHL1u1MRNe7SBtMu7OnOTw787Ddzj18bcTRY9FlWQEd3SLsA7UP80jdUp5gI/AregaWvD
AIwcZ+RQL0847/FrRZ7AdrsL5iBXccKi1Ut0Eshyw+U2N1VWIIMixjBw3C5sB/OoPLBGcjZ3f8wv
qLeIUPtA0L3hXj/UC0mjYtmVLcKxbIJSaABO2hdS9ZUvWffvf+JFKc44vCAYX++2c0NqbDcnNX3A
IIcYT/ZWcUOwCFDSJBYsSA/zur/ASAWqueZ7APAYhuZe6EktnB6rQOItrkQYeYBpZsLXuJ3dFLwI
hsWrg44EBtpqBLxEKjt9IBZk4fefp5ACwF0xnSpy0gG6CAAv69HQtR2el36NhT9s3+lIb+XjMFjR
p6xWJ9UJWb0XPXWq80uKmSEavi3RBf9JTlbyYG/N6Wsqwv+AuPKLOkYs2Pfr19ep3RpBaOywtpmj
tIBTf+fKNtXcIQfHbYnuB2d57+vMB271Mbu97bQ07gOXeDqa3pn90Mf2dAdOuBN/xBHPhRusSukn
TqlUCvzUHbYM0I+YpK7iJbSW1c4lAbgYDW/uEbzRudWY9tK3Zvv593LmQ6+KHF+8JA76keO+SdWp
aU4bWwoOyiSXY/w5jFBKYnCA9AqMGh8X5vHkxuBHlQw9/nncRkf0A5xDQwregqV/Ad/KYMNQ7KDA
DhjDJim4anjj3IyU9foFQuUCKMqvk/zHQ3SM7x39g2HWsmCJp2KsCDXVE2Gz7M14CfVSAPu9dbCv
gxrOJpzxq6WhtLb3oBJdR1gW0MZoP51xTDk6WFxcnsK+SjOyHXGxdVgtfoYZtmcO0TaBAoSohlex
ZGPaQC3RWagLb8+7milRf0uwPeXPdVgsMRF/r4rnadTsJcCud0sR3JAb6JnrOA1uwBQGsSGM9FeJ
KHq3+JHr21nyy9lCHywNB52vF7UWk1ve4nfJhhK1tYtB7oyuy4xGTND0yezksCN8PvtWr1XkCSx9
rfuNaosTO0OW2Uj9qSK4K+jv+srtMNTtVrqhmeVaJGoLDveuinF9gOE93jX58I7qROaHvmqky15i
iaoS/9CWj8Nb7Gsj2ss0fV9xhGUuER5+aEpyqE0xIisRXRGVqeB2hW+hm36+4I0bUXSxwUIpGqhC
8OO+HjzVZotQimLdVv7ZfARTNxFs7l83OFmpeyKVJrrrZ12qpq8D18vaTIRdeIHVOAn8NqiyaM4f
GfcYCV2dfQgzkz0e+0VmliOkVLLorT9OCz04U9v1ZGgjiPV7nASdckTZ+8gIpcvlnDKnNcVM+Xhe
ghyU3ANyVr72rNY/JBcpNKqMFqNRxAjwoDfm/tztILtNmk0JZ1ZsDCI9gckFXFEuBEK+0erB0kwc
EmML5noYFkJJWWSAGD4E6fBMc+L3V2TjMYHoRKSySulqXN/HnybeTGsaBsPAMh7F+q7gadP20kKR
fhPBmK3NRYLLiHARN3Jx5vnx70/hPVZiqMoutjRltCiFHp/siL7nEbmsOKnVr2qW7K9NB9sbdEeS
5SZ3WcqhktiCo3GUkv/D4ImpQlQ2YkYgJt/aUcg04gC9UjljkN6W4tjMvuGlHyrJGIuhUs7M0xls
0/7a4qiq30k7DoLibRTHmorjN4fszFW308LfIG9iD0hFI75YFO+RkQP5SiH8YrTlSt+PbMD9dQDE
CKqDySaHvNkktRMPFLatWGsVNl+EgubcKhrRyEp9DUpvzRakVbHgw3QrvB9uZbf3GZZmjRMSTaVj
4znx3Wmb89MKy3DEAu/er7mLjuASKArjd+XIm4IHl+EPqB+CvCL+uK2hw/oWDsbaRK4T4EIVHXHE
OIN3pVn/HwX9sp/AZcjhkNUyN2F3w3Oj+RMj4qUOYt51Y0RsBQzhFMXFdmkFfDCpP0KJjKKy3pEV
mn+lz+arL40EYB1+aOYrMkj+rqT/61bO0OsdaoXLW0bD/Sl42HnbCT9ilWv4HqzHRBTneQzSss93
u1YYnHfOiz3PjfP1EulmTf6oEicYCglH9OmOdcYFRTfy0Ov04akIWV7dTm7AUi7xGzSAwOkY5w4s
aJZflJiKms77XAz4ktE+H1N7L8BL5+tSNIFj14FoBXGgd0fQH4XGOoxDnwMDPoYep21CX7Zlmdb3
mVUM95+cIgJlLNOn14RnnQVzCzvyCk+9FZihinHO9b0AvabgImfi4RG1U6c+8UEPxVOiHD5ALoP5
Q48WVSiQX+aSRf+IBrMg4aCQEfJJxHkYVY4uoDY9NEhU947mnDkrFvcdqWPHgO/9LXqr6pvcsrpw
tiBR5Lb8SC+lX4Ufm83fkJpXgpgqZM7zAz1Fe8zxrTI2bfwslHCFJvLBMlVNgJ8ydcOg/1eyzem/
JjZKwmr83iRbjNdwKMQW5GwT4cEq9p37bw3jvgBK/AugXNfyU+vkTgkbvCxHdk7ATxgkqVwoA3Cb
RtJtduKm5oKSP+pYRtFZOkKZzkFjVMS3wsIlYGgNsAfmNpC8gwheORiG2gXx4Pun6fgKrUkIVhwg
qjXadGTBD8SYKnnDGzzUSjPreTehKjpAzyTuiR2TEMdrPy27UsJ0aoIR7o1HganHUUtVpVSZflrk
1zRtMbFDqtio/orraZQp+bjUoXzdISB45961RS+WYiRzZHnKhLYud6EK/ToQ8Wjsn5OkIJiWzQE5
G4t1kVaCAUt8sSnpq9eKCjUIqRoHOJCY0k6jLK4pl1C0Cp/3nLALEJsup2e3njXYKZxp4il34F0s
lF08fBA1GT23aUKWA5IRWWcFzCPSgpcyGRZmeUvqqH2AMqg4M9sdijUzPbiMrtDxWlhwsxsRaRKz
5oQzROu9mkmQriH/T3yB5Y49INpFN8LTOgxC8+8cHkwc6Bqqq9Sx1QNdysCNIWmN3nOAulZqPlzb
BOWnmR5tcabFr7u34hGz7kdkzgnQJfC0xpBEHE57knkhlWDwAPlL+1IlCKHNCAgmBbUevOWTWTrd
wQgt7jywFNeKt+/PJaKr+5wuF4AYg8kb0lwvmWxkOeXK6eZm5MamLzpij0visR6wiNF2DTesgYV1
2RojGtHhNawYZGtIkF5QIv9eV1N2Hio/n3qIWwVNOYS5Kdf6X3qezA/zfCFfMij9YDWI7YcmHv3W
g6xA9LFhN6y660eaiBFazEY9nFSNQ7AGrPQH0vtwJFcLKxm3mokV3IIV7x30pL3e8rESi/KoadCm
HK1N05CPGfhssFwUvrss5xKJOXJmdDOzCCxeLOPLQSzMzTJmi9CMUn9vs6tTI/dEJRU50FiTryEm
uJPkDUmNZET48tsgZ9b6D/1IvN7iYL0PEywCw5N5in9lta303MGrf+4eYu8yXqlemqGXVqTIgePJ
hvGZg27Ae2u8m68udVAaEPuc00vgSkyG3k+IF7GAUYFr5KlKsezbtdA5EFn8gqWOYyHX9jwiPt8t
1rPtfBdtoxbzVFDMoDDiwt/2lYeVPjG/n5ny2Ex1e3q/+cBCanPoI9WEbiVA4dVAnIfLJEY70tEJ
Z5yT4i4q6erY5rMKk8rQg7gNTYUrIFo0EJ0SF2LiyLHOWMXox+mWezGknk07Y9OUUAl3vDJ1Hqks
jDq0hTy8dJU6kqdQAIBCCl8xvrhPudHJXwyx/uD8v1TVMk5EHA5KCgbYRR6VTCA3j9gBdp5v+BZA
Z7N2x/pYeTkxJAE77zMGOgI1DVj4NcbVpMdsEIk+qNEe+tBrte7FsOTBqhMC8Y0VExVqpEQwokYo
JWr4+XHp/NDYs69YqeqCjkmILVeFhRNIHDDZziKKkqMJhSmuYJ7k7fkn8rojsD+OqSrna9vol5QE
gLv5scnXNdOUW9KaHrlX9RruF8IT4GuoahCLagTIpQHePNpIENvkaTKW79hziFVCKPC83G8L5e2W
HFvDZP5LpLni1uyS1xDEXh28nqSjFlpgez0miRICS2zkrWsNSL6fK3ZMV8xhEcn69cW/S0Eq/DL0
mFtQoP7ZWmgCQoCeD2MW+t3W1I/g8vMcsCRrdnrWSTiIe/UnwNcGVi2TjFInU2Xy8mqL8qOX4xOD
WnivkI/uVotx+02xjqIgy0ATxdFap/IbskYuVStCTN2VoFOz0x8NmhacFDS0v2E2ADUJOkcePQFI
gsIQWpBwmBYPmfkkjW8KRPgHQlvjDAv3pAtEQMvuFW/Yxo2KdKhnXSUq87R7XQ+wPrycysrDKG2b
4nLipvFJEuyo/V0u3uo2yDF3zzCAVXO1s7RElwzfhaRovxQMR3y6QgOxWhK6QcWt1c26T/FpWuSX
qguC73ZhZfC0zC0keTd+gTFJsxsJplDDVCgCl6hgNcu8AQThmm1NXG7BYVMVEQxB0uO3qP0L1JaJ
U0o8DSLdM8UG7t+IMWgCERMlBLIL/oe+aHb5Ra+6feZjMYSzubpHztJWGrySfI07m01Qh70ya941
dvBD2maV6MZyywkjQN8RK5+gd1LfLPEUmZ9c/0Lq9QetIqaIj15sKpTLnIcJKKP8EMtLG3c+vaUd
Sct/NSn0m35hAomXgu/oJ2w9d9kHrY9zvKlKRkCA7Hxwv2YNweZjcMpNccuKVxcW7jfVH1p4hIGA
+thugLrt411QKXaUw7jyQYO+XCDy5hY21UkHdewc1gda2y37+7LyDZjunZQftEOI6onYjx6zFCdC
20dgQL37bFWDAaH9cRxYXYZ5R8qtmQAi9YPV1nakhfr1l+Fh9TEl09gDItW0Q5ek3mk5cdQg/jDL
yE1+DtqbNfCC8oee2DsxUPxJySYTrxL8BftPCgSDCKHPvf3MpcxWY3YJBIvVuGKytJrYByxJRDuW
JkaoltyCJeoItUAr7t/E0Vrnz7aYqFc4wroTprnC/rIlRzAwopm0BUWnYXL8/rou+tGH2Hnk6XZ/
KYDjnp+Pm8ALlmEbuwjGxCjeN/zjADC5XU/9Kh5Z6ceKCa2nMMUCd9BLoRGjGVnMHRH8yCv6Fl19
CgkpqcZc4pVyammh47gu6nf1c9P1ccqJzLjlwftkyHrrrOjidF4/0OOrJmTkS2WQsJeBbcM7sNI1
yDkfKjgrKiwHT9JPBPAf00fH8pqO6VlCDKpui1WQNI6y2PpkE69L904VdZOzPkT+kdV63qEXumJX
Zjh0JjiUNYyu6xPB/Xwq9ImLtJ0myZ1xd1OfIKywV7AK/4x3/dpGJewAAFOGecuOLTA4USE6DuwT
yHJR03lBCl/K34f1uauNI11xC1o6dkl90TCZm4/VQ9qwPIAcyT2JdLIvhgSfrzGftZrPnLMe4BjJ
5TyHzEK+26hr7DCkBsBe/YQNNcJM3OrGJYncIJUVkrUMIc3sMdCFubRUlXUN/jpcOuoQ2VovOTMK
vWqvIyxq4ZrurBSkL2nbyNffq7E4FuoQQOy17FermoZhneiYl2m8JmbeT0XMi2haV00cz29rhNbh
eTqnjAEWVb4I04Db9vgL6XVViMSnqm6wF1dKnUAaBmX8VpGgCUaKKsnf+0JlzGsfwOdVBBfXIFaS
zZg5zC843z3QLF/GQEcUcQVBA48CktI4QAI/ovPxL82O6GcwWsSMzwfTrRcad4H9F3xi6d7zI0dH
ykqGzzJmiTsDAiqvkEifu+V3Sae/+da4GB6ms4MvSeza2sQ4FUMZ4560tEE/lvwxJoxCSXBCz5Ag
FrndFfbeiUxDpAYu2CG0WvB0qT6l0QSHP3vYTZPl7DNyYT01fwLsA21XQKip9wd4EB4pxGDvB4YY
6Flqi8xOBa1F2tSkMXldCFRpWfZEjm54nmjvtQeLDUvVVakKZtBMVdv6mwwC3+a7XtQuG0lcGyh0
S1g+qNeG/XvRUJAuMYuqrfDWh3l7rjgs9XbhqrHtXNGPHVlG/KZA82vPz+qXrQdXQPN0/Iy7Bexi
CMKo5s1eokTc7ZtiRQLRf11l6Bw7uoRaO8LReisyne7JFEeG7vtYUTReY3kZJVZGkMUalVvJmoOK
EmyMQjdf3ksepBIDH+KS05C7QsNcqiRBN1LJQMTohqQTPmyo4wpML0TrjG5doBDMcpJL4OATC0j/
dINBp+0Rb+R1BMKSFDQeOc2dFG1n/Uyu+AS43RziqhxaC8NB0emMdpL/p2sPd3JSq0CTE1TPRtgE
CiUd5FnO/PrWC0N/XXZYREQ44Oqgim3+pa9jmCZ98M3g8DHl940PdIjU2vPO4UYuB/hrkY6b4+tB
UD97voeBDMP7cCNQptHY5E3hbtbGCbSTv2znW8hqCMhcsOItuhzfBI4ivSGlut9Zmzb23Soy59NA
3fkOmSDV7q+BnX+96fSvd7/8ujB7BYy3/blhvzwxgzJVLmKtqR7npZCoMPPJqq7JROIi+9ref945
5TehsfSnpZOozi5HBIWjwWGz5MuWlnAUldNFFXlIsBU7d9nP7DTKb//p2Q1Z5MBbg3kZgXrXf1T0
0r8OBtaiQpW5Si2Jr7JrqEHy1ssMsO46UTYmdBMvVZhEcumna7jd99oeTvnCB62ioR2NT7FklQOi
/36supUBLZkOJtjEqtw2i9/6Frt6Ah93af6CFi4GRhykco+lDx96NliauRijNuCnEYkL7tinF87P
8iIF+7sELPX45wnycBPBfJ8WkmhG/Rkkx7Y9FQ7qvn4YqpPQNB6q0BkumWvLRychMHnISOXqE42o
uZ+NlcOtKx/T+6/9nrqhO25CEN3a2IH5LskSprK/53JdHaphR6tyvy61iX92xJYgZYnO1PkDy5zY
7rdFVNDGBhpZu5m/bP9hU3Pj/H7KZM/GFLX9Ic0Is8uVt4BneXrcqUw9iZbfHXdSCfXstL7vYkEm
yNKAzAfcynGKz3XGtOq0LbAc/KvzacLyLWvWytmnslSuUeYO10PtN5W9DhVRJgINmStlL6Hpf6pZ
QyMxyEXiEqgpQxB8VLAwT+2qOujwK0KWyItr11o6rnxYQjGZtZ9p60QD3HHz+VC830G1n6Ys3h7Y
UWAhSHfYpwXvhVTvwmM/1EYpp7zs0wsJo8yj4JKz8T/d7/6G++DAO/eHAXJJTDl/qSAur+MJW7uL
nqgoNQHzl9PuD020ipv+DJkPGVth0tjPcDemlNAqIuccMJ6tPGxbHTeKa4AeKjpZH0qXP9zHG7Ef
zhEUPHJb0mQtgkXx0J5WiKNZDs48cBcTLCkVY8e0VP7pFVjey3rILkSxVCYd9oBJIjK7/XxYnJSn
QJifKzoIuA/jshoszcp3BULbPiqh5HO8sEyBcSXMtLTOHCkVJ/gI/DJsXCHqoXBd9yU23e3px+lw
n9LgN+Q/NdB9AxtyTqM3IDefkSxI+MBhfDdt9OKz3Ki6HwDfPLvCMGW5BCDszo1V+bU2AMtSrR+2
BZVEQPMaS/oWOdhCcgjKpkt2RnRAH64/IQ429J0BBLfPhxpXoO0vXs82mdKiu/bFEZvxc0JmUNiz
xyHkDfNQLghjKZn7oVEcSnmph72CRAzi3xMTWCjy1u7DhT+KdLK1GoJKcwtMu9mgWOG5hhTujoa7
6h/n1u6qaFPzG+op/kC5Q/k7zfX7WGpK142wv2jz4K2J6D4BddVlfK3PDN1PBJUnrX0rk5q5KJiR
2NdB/w7XK+tMpMLyZvL8KCHkKDA280GioNretLTK9vPMes85ojzA6XGPKYxvp6a++fnmjqxsMszO
rOoGxWOjlMPumsBgQF8dRYY+pyiLqUR7BWOCUXyl2gSBaK+/JLo8TVLcDquzJ5lXxdkWOVksEbDm
9aOxA3lASRk3yVAFZ7Sb94kD+3hzXpJj8UG6RgJXHHqEuwBcdBb04NoaVo6zJwAg3Vv0LBtHYB2i
jB7LaU6e3kXXaz3EHlsff4THHilh4kNXfaOuuSlimQqzDZ8Off2bjkm2AvfPreyXcPqBlxXeh9J8
4dWvCd0SMvqaAe4rg1DXBtxiVfPgvoOu99NajqcsN83nL5Mc4ODbJ1Gg+8dmH+uzeNADMAHAuNAt
GuDS5TkqvEDwl2yvG16wgm9TjRtisyBOggl/F3/UmSu9mZybtbQmhOOh4aYAAWl+GQ5OTBmmtjnH
Nzj65RAfAJR7iR+VGFasbdKCabd/MzoWsFTiTZUE0RTP5kCJZRWixIRVdNCdu5V3sUSDh/0dk0dy
5zgpDgBkizNysF0L9ItFjwdM+DQrIpHNNisksTgUpkDWYHBBAeRF16AFMKNEU2ddnzIKn5rRL2z8
CCcfwVHxD3/w1TvF3yEBbwbZqMru/1sKWmmTew0X87F1BDdWxzwGAXOLH3TNHVT2F3jnOHLxL6nq
tYInJC5yGN1wDF4lVg0vx2PNCCAq9Cu7bKlMx96CJML+TvlVHktaGHHGdxLmkZG4gskEkx147QdG
JsQGRDtLMMRVQm7oyV9EngJCKmVTc3y8CyOOp4WLos3Ho0Vwsf35RrIsWnoy/YIayiFFVVebhJk3
tY7IiX8/pfv8zGFeI5Bl/AobQ9BUhljuhvusqdhzbNL51D4TP8hvPHM2ugs9AKy9uY+XBV7XOGXG
ohRDnsW/8K5KmuAi9pqxHQebCn4f8vagjSpZHkyvijUigzOyGOuGmStaFc/RdJ1WSTCbwb9m9xcl
oP+qU46DZVt7J6TD/JIv7atjqUqXvnKfmPCAOb3N4NV3IwXNc/H++0Lgx4UyIkk78vc2SJUV5h8e
XCJGB08VNiBT7rnksbuKGeWKUKiJlrCB8fsnFRM6M++7Cww2+JlI7zW4w10jwZwjKD0b1U+ZaOWz
Sx/R1cTi4Bb00ujUcDh4CHkhcdxuh5WuSzErrDlM9F4YG3MSn0/n39ZQIyvAbcM4qWDVSi/nAz4d
KieZZ2KwM3ntzLsbXVyOb2J1E5H4nbvHzxBW2TW7sssjdMHNpmbOWWOLSdSfyzYJATuxMEjwYFxa
HB2WKWhy3scysxmsiEs3yYN1iCYbSiyZdLQWUGf5FqPX5xdMpNLF1Ryg/adw8hGSAA760hMi1f7g
3dBYOe/ETh+IVLCI1bpnyRQ1/uloevjDqeiyEpNCeRzZlzQGMgCyUX4IR4XnPtmlHqibWGmo9gFr
QeXV6CEstuIF1/IHk6uFYNUfVi63FSgfi0XIgGPKbFOWBvMZdJHmy3fKZTOxmmh4b99+E/KelRo5
4lJHilePdQpTIbwfAWoM+O7P4svAoF/Pj2y4vWbGMgqrfZwbZXyy09EAzyTMOKKLRpAs0/ZGCIzh
2MA6ozmvd8B6KFogIYzZV/3l8w59BEg49u+iQp6/iW7tVL+7q9vTY9MtBXdOGVyjyZFw60Cc87Fm
9Pb1qvQv5RMmTohpDw+7/Ph5zaRNhboz8xzNsH3TgxHyboxgqV3Ob9L88sAZZqADituWw9NSHIud
0twski1ipxLFchQ83QTjlWj0e6QUjkt6YNf7pcT9zK3piz8Tq4zMtjJyBfa4vdJza8TyGJ2SDNL5
LMmMN/fy05S0JvOztX2gw1JXI0Y2tcby5KJD3yiRDTDYvsp0yf9BT0jpsuNHVlAfdILMJvvlOrIR
mTq3ZUrbSqtUqn0KjTBduJsh8sldMNz1taTMbSOcBZoHbhSLkPqP0PsYWstAPBKo5TgCZ/ww2DuZ
bv/uKonnStlPT1Z0gyeKHxbCM6nf4faW+thD/AzDfn78BSpoKlHKJOgPkHyOXUuL6OIG93fgX3Pv
i8WgqPbXK2j9BOIJlvTimXVH4lJP3X2Iq+aKUBw+9VT84E5cbCcgoFeEL5pWaFMWNYyKQ6XwJQy7
TE9wSguTm2m+x+BKg3zEZOWEFnC0TkpGGB2rLazstaGk2UmDgfV9Qv/15dBWsTzcjPC5VA0vSJ8N
PAmRt26JLvBtu4vxZY0VRtDnimlGHDZEsPvdmyZcpLJC83+0kXj1P0MwmpSZ31graGlXS+WqD5YQ
X6o65Yut8q5V3JB3CDr0WpdTrMxb59pn3x5Hq2SD9oMrTIdv+j9rFVRrYCrUYdKSzm6wm0AK1TNR
u/d2wcQaoUShCB6+h04UFQ30XsoendHTBKC7Ak9JaMddI5RWMiBLYXo3m9HPxzvkMX/0xvbmuUkA
ngEgxirCdGZ6vTUljSOPOhy3HwkqpuAR026/Yhrvf/m6HbXSEpapxmo748jm4jtDCjVrWM+AwckQ
WSflbwmz8xMiRjAd35AAMioMJu6LIBKf1/gghvuaTTDZtIRQcAI/Hrpnye5LLMhXqid4bso5Jcd6
nfOOnY21ozKyLJViE0HX7xcx2t2KVjFDzENvFdxMNwKQxYcIKuWmg43pcgm+CdjZCVGcDmOWSnSv
OM7Ulezv27EyBi67oC3zE8r6pcA2wP89mOQzsBKjKxGxoevsxdNd24kcqeyuPiMB2OJE3Qy+yxML
RRRc7VD0GCYFo8yZYCJKjWX5m1aYTPcfFsTNvY5sjbyk9T/s+hXS+qZuCtfi7gQ9Up6zisH8UKkB
BoW7YlLequ6HsycqgVSPsyQKxVaCEI0husTiHK/+eLzS7zHYS9O6kJ60jk32UaxAE8wImJpzPzVE
ZDfSyrGJwNmEnRISVhtguEPNb6Cxqk0AszgAFQg8sFA176FhwuzH3eN9mJjJ9wrraAsDXP5h/j3y
LHra0KBAIDtgHmLUxce+JgxuX225W4Vfv6U4gmbJUaMaqge2WWAbB/CUJ8F3iuGr07sKlpjxxw3+
O9SaMp5f19uxOfkYRKQjPIMUZh1NLExEZCLmo9QdvDmGxw5qau6bGePJpbrDdsIpZTcVZl+5LN3U
Ux6Gp91aMClqTG44NqSdX8M1+UuHYMp/mQ9WKPeA9S12C+IO9Fs4UMMoZ0NLGU6VdSZgy35RadfS
gCYK21l+JOQnGbr3QZeeoUVlqftBOkAwM1+AOvm1THR/7/nAieuxl0LcEEua8bEF0QGpsliyYC27
A+zDe4/0NCIahD48okwEdBP0jhgpWnWtshN6FXrjJrMykhSkTPdFqN4r8NMeIZLuvtK4uencCcIu
okCMUgmLgXcm23Oj3e01o35Pu/K7kJOheCysrMMsFNabUYJJxfzLpqq2eNB4tZILKQu0d0HuNGz1
lzqtlHfEUFuQqPRNaROjJ/C5wXF2Y1nqaxK4UP4QT58M9x+UrMA/rHwSKONpneYvVN5Mx6u1G50L
bYBFppd3RkyYf0PubO3MilamfSSpzp/z7T1/SjIXqt9gLNfK3a3260YAig2aPT0ycmHLFG+piMMT
8fkmy0+F/CjaWas7Zuco7zY0OUC2Tvw087MACZ0m/baV/z/3/rXhP+y2UsaviHbFa+1d78KC4G/W
eSZXtygdI2xZAh0MMylISJhdx4PWgsTPNNJ6YvNUdoGlrqEZKMZn3+l6yYVumaWaIcEnhWJf3KnZ
QtV3FJDR6o0bjg7bTtHFlUfvlm9ynCtv8qf51/0SnKB5Qn8gcbfnPfvlFfjldJ4HRuGzFY/nC7Zf
PIgKe1qlp7ZCwjJVMqsIcY4QkYF9oTY/ZbLW7Zi/wZCAkHHWrghqo+OHEThUVwGLENWA75PVj8Tw
XnloQx79Ag7VI+AR7V8POsL921srRbGPy48EuklQ8uS5mUAoXrVJH/anLzRMOMMZ9kV+gTAqJLOp
Ep043IhYRzb6IR5CYZYSx6V3ASSgbI7z7c3m/mqRQTdLH+xfsckp/Modfc4a9FJXrK5Pfs+b3AAs
v5svoUP09nYnwpO7FK96WkctnxSlufOBrYbqNB43+q+xZpN62GMVd4N7QQLynUeCMuMD14XNInYv
OslIS4L6KXaxKtLL1Sr/KJn/98jNcqETdCBtTihliQ7osv3AZz9eQO+8Q0T/szxOR3z077DyM2L9
DD8q26hHxyhVnBYG3X/qUrtuqCg9SX36q4CTWRDBeW4PNTferby8UEX5MPVl1HKPrGHxtR+Q1zvQ
zihKT5GHcF2wVj0sQH8DHE2e9JoD2GN0XniMMQtVLouuVCw2z2z4ZFzJPIrAuaXdtCW6PXAur4Hj
Fz7zEp8xktRnAWOYiNrbvmLSKKV2mf9tmUVkYYKiSyX4LDUMk/lmUKIMQ97a5H1SPXzbVuM4Irq8
DNxIWG2Qa/Cwc15ooWmG3FQzvxpSz33B/+hp6Nev1ulPvcCyzOvkaTSRZmT0XeEpqFirPDwYQQ2S
kYWrNSpuXQiutCYqbCkxU8s45x98VgDHHndggMOk76Mc+/ic0XmfPg+O0ymA+435S3X+C8YYLIO6
QoZnha0bcJqxjbfGCnLNkhJQwU0hOJaH1jgXViMC6347gtNj0YkmYe2eZzCGZob7F3Qig679z1zz
WirF6CHUtzkTdXhC8Fia3pH3sryY4+mBajMU8jNKFQk3+ftPzTXFhV1rijzdlHqR+W0cKdaVYfAQ
WnctuwiwEq1pyZ2vkMCP3Uwb0WFtmHoGBu65pCzA2AisaQWdoNR4SLlsVUnhkTq8gn8Z9NScdxqw
LSvvuVmglAW16xohOyZmh3IxGOufVNNAQMptHFSpP6hJL7ZUoNefp0lcbYTHSy9PiNPAX6OsWY67
OFxsz1itpwcMAqfHQUhpwZjFXJiM0Zn6quMrNGgGVO6fw9UVS9vr95LrpbIaSgSFMZk90r+1Jr8K
siyht7z1ZcUW1J1a+/2MIt2XXu/oTTE2iyaepurIQSC281cBvKkpYd8HrD4QGjUGK6ANaRE70XoM
WU456YktnSe9rh3ZgxZOMumftIdEMXBZ05/bAwFy7qp7kMTwbU0rRFRa907H00qfXT9wXlf8lxXz
iKN9z1rrLR+o21WvFXb3O2bZ/UdvOEcDL3cUfQiN1GUGaXTtKBYYJh7x3qxJlSH+e/NeGI/MbObC
z6T/SsIKCGcn/lPwB+tTC6YGZiyO2sFcQwHv3yGzjBPuQKr1LvqEZQIcek7fopNRjh7SUZXmtX6t
z8wyHMEmxVyrFiFNP31pvHNTug55DcVGPwcS7ldnIg8ywdZ2RGdGkcD4A9fbXqlm8nabKPVozZCy
GDsv9xz8rLXyOPiux1XMTTGU1payDnociqzm00YSIzSNOc2G4dwKO8SbdkOApJZGu3H9zOkDhw9t
nRUNwA6Ieprw5oXN1V5ey3RvEZ3AgIomOMi5xsaetsuVNolQzQak/0PaK0AYNk2GswyBcD1NDDIl
opyLm+nNKZtqCOdpNf96IcgTWVgmS86aJuo9rvLw5qU8DDSneVIBNkhyp58MN66bnqxcddweXPwz
9cQJ77NZlzBR2q/ZM4Mm49IrWIiaF77bQQ/Xg8vYa7Op2ULjS3fYO+6cF+UkZDbBJMp00eHVRuw1
V/Ak8sPPJULG/jKRXYxJxRgX/MXB0MKHRtPDxHJxWiKOS60OHNLa6iglhWkMJaB7hKViJTL/oa/s
Y31mXAg55SJDbariAuRTNwYwOufLh4yQS9lvQjbSTkIj3rgQFFfeBKKkeyO1bAjEUFyxdB/PzBgF
OSwfXL02gbgUeRGtPIVaxQ6vEiEINggT8q8kGUn1deAYwDmTZOG6xny76fO/x7C2Ih4lELX8P4Bf
H6QWQZE6RdS1N2z04KPFJW6r2kL2r+x9UNrotVQW6Q4OGCSjVeZ9Rl7jx2BMtX3Pud/qx4+xdnwz
yFuCxLHeMLGn9EopawYLzktIlkPUnHnfCWGfiGvdPbYya5IrhKa1fjUF8ZrShPFA6APJUgpbofce
Ranq8gCdTC3Xx0znyJPB3ZVNu9vHJ7iA1eDlC9iC1tLpxxT9ywMR+ViZsdBicQC0xaNRGkZlqAvk
060JRlBAg2cmrnXFh7vwNyWxDNoQHEyja9otVJP0+M9tj6lujLXYSQKi7Bz/kwKPrpYT3PJXnb8y
XjPZ9Xk6c7ZMwyw9FIfmmQA0B9cw+BurQQtyLi2rvs3X89wiJe2nxGwm6Xet1WYPXhFD6F0MSuM1
nx4wHXdOx8i/UccqIiQA7ZGmDzpKurWjS++bBMer9hufNuKog0YGg2CFHmxC1DnFXxQLP84YsHOY
Uvp2Mz4I1o/xw4GwcP53yklxhuVGkfiLOSfy3tvEQT19wsy6yWB7aeOodbX4TUDp7HzqC8RHvuEN
wW2fimlCBOMfujm1HazB3Q4ofVwvN5QKDaPaGAfp+Up4ACndw9UiRRzML+gFnwHD//0+7+/JuiBZ
08gk5qfhA15Qe2nlrhVBe7Di5u38MlcDdkDZFOz9+puhPxxskWJcYRX/ABfAv9ow4yxY8J1P2omf
gHCLR2KUZ5SGYq7wpje6Ti0j9XutgKn5xah1MWMdGjWavsckKQtsYtEp4+3GO3Pswfn+EnBNLi9b
56xbPxACivUKnt32AooaJ4ftGdsbmQhpKLJQwFIJjdfTW6IO0CUssxYXUqFsRnpl4W3MllQrETBc
Gxhj+EL4370Oz8EIxbJgPcwidAQT9NzIus7EbmTc+exZ5SPitQHW1e45Y8Arx4Q9p3Km0j23n7Hy
EIunGg+bDEjvOXUgWXT06HjzE45adx66MkK/bpMlrahZchQ6MNjXBSIVxHtP2+vd0ZSgeRxHWxgc
HZJTQL8bw/ZvuwenTywP+2wkjnrx9IecPIH3NJD6D8PTqlLS4nNJVRAvGOo8sPKEDeA2S2rvWCZu
YCpLSNrPaX3BM4WZopnHe+mTaaQzhYJdA8Ynn/mlvk8EToA7FZYwM2OwrnsF3DyfwDxhVRiS+cCd
pAkUxV1bvEbsRO/mewWy/t7TB7eV0WBFHEIMvnutLRLbOEHyeUtWYcWl1VlT7o4L1snz6OEecKY8
g5MumKcrNRP7ZN3GYJjkDr61RCDQ6klfRlQeaMlYgSKN6UAzF/rE6YfeWulw0qBavdHxwNHhOTtF
AsQruZ1jEipI7ZOBP3i3mDgJxwiACxpA4Ko3q7nTRJNx2ugF8BTfLTzKFHUZCKfGSgAGXuWdnI58
p94DO0CeYoD+ufj8wnY7lga0wXbrsZu1x0r7nQC7PCYvx9HWt4PY+oI7CCK4bZtcLN9e+WgzBejx
mFSsFmGd8RwR4QpmyklQV5byoyijcTcn393VO/VbnNdb/6rZ/ItH+eRU0REhwPq2Tmlwj5+5eoDc
xD5If7xJcmFxtRznLN40dcjs0lXF5vAa2gVKGSd5lZcMxkhpY6a1T6LLWknP+jRkmKEibnhX2W8K
7TOqKklx5aku7CX07GJcO6uVw2djXkqudJzjb2mtMNMjmUTewaz6Iw9kKFx7PxFaNh/l7jeaca+m
//E1da09zInDp+fc+lg01RKTRNcLctJVsIF+4DQLvJs1f5c5/TDxV1wWoozejG6n1nbbsioBBFRD
2XnGbEGRKjD9IFg8gQrDF7dXrxRHOEVA2dK4bEabYYOq6N9RQJdkWQLvoGQUxUV7tfxjwQObUlyh
qvC/G+PnkwpDBZtnY0I96AqXpbzXtdIZWTONlBCUcK9GRK/CcaRPuqu51nWlhEiU6evpyOEvJss8
3oSdDEsMpXQKu5BoI7SikdcpAxjM2KlPF3mopatOlsM2Bwefy7ZyqlTWb63/vuLDSWXp86ncukjl
OgIGb6LK5pG3B/6IEkNY1tYGfu+bCnLWVeJUG3Glo1kiRLucg1UJOMHJon8T1Zxyv2gl7apsLYZP
bYlYVx9npXY/i0lckTaZYDgaNvco9PU2ppq4RBPab/0K90iu5rD9U3xAjDIi0um5edrgXijnP3T0
4YvigIj+jQqGv58JwbwKIg631TN2cZ8TnBjTqhB8fthV7a2HFwygTHi9JUaXW9wrP9dVMqgRdtGU
mFlwWGuwG70otuP7seTW1MZcPvdDQQee3AZetBhZPCmJ9MUMRCHvEjLRWkoDj3VHGhH9Y2yw9wDS
9+mVplfLP8PLE1j+EyAxFFnN2dy0VD9/Ou57E+fPkFZVeYkbT9bh8dFQAppDz5Qx9DCm+5w0EO1l
FXWoOeEATg/vqFlf5RBXU16tNGUJPrySXb+W1x+YVGdQzcsbhYjRg8tF6VRA45Uomj7RamB4Ff3u
0CYcpSrBrIB67Md5JV8WLrDXbEp0dNjYlVg8boV96wAcaPQFWtUaPdCTyzsugR2925qjqhaTYlSe
g/IuPoki1zD0xCCcra+33ePaK9Irw6maI1E1deKhSlBe1NwCsOzf7mQPYj133GHewshdAd4yUDLh
j8VvTRi9CFsZJcJ5vptyszrvbi4HEPEHnVv9Dr4gqAPIv3FUP3GPmv3nX6JsApaJyNivj3Ganc1D
sEMF7u/caej1OUFp1NphNR8czkhNoOue7BcEv3efzpPA0tAUiKbChGQi84ru7jCKPSSF55wtnarS
SUT/z4vRxSz0V85/EEXI8ZZSpOGBKWxdlTXoNMkiCTllRVFbLp16kcpT6lB30z8/Lj6Si4KhUm04
PlaZxgisgO949BE8d9V0ZcQylL8Cihu5I+qVcInO3IgReH9pO2ABoTwzAoryJIttk7Xn4tooaSFI
E9YdsUCZuMFo2zrpLsLMSmkjpmeX/FjP3U91QJHwRSujcvPcvEueRZrEMB4mAE7W1SqTMzn/xpje
ED39rZtp9dVU+Iloy/DCVVx6/kVmdjodEcLMxNmYB3Ku6SYownrk/SugL8lpZfyY4i4UDNKxPI/k
Td2+rZBTkDjQFmZNkpzqjh7Yuahi85XR4r0pFEw8kWn5tF/wpIg65DkQ4XAiKI4hUa40XUiIYHdC
uS2g/PqsAoPq6YMlGcrz3Ggz0+NzE3TJlOa4BrgYdIZZamincA9+8bxOTQ3g6y8eFJxQZdoFja11
BQJHyNrxnXcXsgeRz3I0bPfsvUuWoBOcarhXKNGOMVbFg895UbSZslGz1uBEpaOl9Ay+K2g/fP+t
CAP4ltZ0p1xIrN9Jz9QLxBCWLdUQqdtbe1/sEyMomkGFGoHdP1pqyQ6puca0SzRDVugs7FP1rojy
V1T6GSNZbJhafOf4dcwhi2cofA6tIq1JC495TQj+FhhYre+pS1tX0dQCA4Zx8xI4erba2qhYhfXW
2Sr27exbPnHCoj3W2BXJYOp3RFtI12R9LaE3rqq+QukdaTXPo7utZbOVv44RPKNHjKRDttHvdCkO
8/MatL7GgZLxr4/kxBEbxjD3G2ZSmzzZHV067EQ/Z/qAI7zGHyPE1duJsqOLwaFOAcxreGngLk89
QLn7ZY8e9NXl81D/lxJBvBMTBT/q9mTYPRnU/eOqeWl6DpVG4ln26H8uJBp8wdvbI4XA2aEIsUlF
m6189gn0hVRZnR5Urzxy99iYSO1F9Ivg6fV2A98jGbVhFQc7gq1M57sbE9VUu5OE4bcgzptfVztS
+o02BHlNc4Ys+Smbufsrz5x/umcW52zlkx0zIe3vgJ24g+/KFPa9x7SGwNS8LVUS1rXG/i971YRj
SlcgISvT2tzToys1WBl3e2bSZ7EPX79a7pRsHJvMPi4LXdl/blkGpQrFKKv8vLhP1dje+Z8GOk4w
r15RSEcW6jesbpECdnOkcqeL/h0Aw78kfa5VBj78SEZFh26MXU5RyD3Wit/74jS85ZbqS8gGpLNs
1yTLtyMCZyJfRkjrjIl2dJgVsiYm289W0D0QYEc1AlwwCrx1r2WNbRfqhI/mihYQjIKXpOqBxwR2
Rl5iqmZPBM3YE2SF8oCYkUiwDL4xhe8qwEjZM6ifOzPEBrU0Au2hI7SLz/Of7NusmjOYPFOTJVXt
u1W+NJYmNai9aF20tQp5dn1wR4/Nv+LIHpqxiTHBG9r+r1doAMn8UqZ1KIuQiFWnoxzEqgQpN39A
xEowwLYoo17qe7Xqr+wA+umq5RfAnQsCezIxenbFwK/a4EJ2RBuodv0Mr3oJFwqIIPKuhnjR60J2
8qjkbikOZjHSjOjHTWl+9H/1rSMqoBEfl4d65P6jK/j8deTz5Y4W4AsSZsI4yY1mCoKyQ1Z5o19n
BnYr+/B4lBedZ/9GwcrsoNZJWwiVSQ4/jRpNhakrSw2jopzqfQNnKLR/NOPxnXC33RuqXeaETM1g
dzI9C9VB7XBKXtV23+facTR/DCl9d92RWhQ0m7s1fHizoM8UNbWLWhOF/MITb46tB7UAZQ8pSF19
Y10F/MEaJrQZ5HhjS3G/5UcW1pwI2ZtVYrOU7ln5FGJ8oD4vS56Gg0we/tjs+5nzRmT5ayKccSjl
aZ66yDpvfUnTm/I99SvkbX02XD4dPhJaTaTNxDxD6qaQnRMMqxWtE83YZKqQmTJHR6XUbKIGwsdq
Tg7BZUf497zCuBMGMm3UckJwGv+OG8sFSrnYmE1QJZ4Dh4WOx7aVeFXegancpKlqKMrlTnH5pD/+
twmz/fSM41Y1BkvGZe+BNnxY4U5gokZ6Bo3tQsSWYBDBGUUcKiAvo4ml0ketqgHeZ8lgBMDh5Hm4
YItCqruBOobb1dwxSxzCRC3Ypei93FUMAWpmSJuEOScmQ8wpyR/hErQsdIoK9peRkvhPX/oKU9LI
9HyUZdzs7cF7bi54ywsf1OxsRfiAJwBv5aGT9FYdkSGiyLV0L4bBCEnUamwVWmHKlKUbRJCO/nnd
CbTd6qAz5RgGOtD+sFfpxOsBoqIyjtdTz1npms0M0ONzXTAFGU2Tq1nr/Dvk3rQP8vTDH2u7nUE4
HQWKBXgJ41l5jy1Em9Bx9yVUV5MYlRyHfeiMm/zvl5uvBMnqjKdRpoIeGEgTcodkjNcbDNvPzMR9
ZDhryReEkjTsFDEqDzQMBfL8poD1BenN4eZ1uZRd23MfaBFBrWLI0jzeyBXexezafIre1VJHxEZW
3r4jPODj8z7nngHb1RK1lLNRRp3d/IGFuxI91E3qz256PmqXz0Z48y+yThDeFDRdR4yxCcaH7e72
XqQ9xsEALeQZQ1QU7Bh2ikueQZ8ZPTWdIlUuDKl11wTAGqTk4u+XcowXxhfzI+yYpoxcNEHCrkPa
p9WKHosqum5JpNz5VAzF3B0k4Q1dMdK3AD4kbSc/0BBRiKMk3TPrZq89D69y+oqEG4tzUdtGb+5i
ActGpme2NEURPJiXpT4HJy3zJxPWWLmgEnhPjbBIUl2/5ltidLIjhQT7iUElb3jM80p3vhdj2M/N
bWv7fXw2mFxKEHtGE0WdCB/yzzGDeor8aB8rT81bdi50k14SN7hFHpNS9GfNEqEZMTCzPKHVAdvG
DNVcdLvwj50eSHq7BZ0Bk+GhTBMQh9k+AQbOu9kD5Md9RKHya+NvrROCp64gbqmV4CD4gtc6kaey
QhaMn0MLunU9iPKDXZBGN+ICyQC8STXBdt8NlwzkdebzT4zFCi7h5oe9zu18gYkhBY/jOiAnMw93
s0iNpMj36lsMdek8cH2fOTGtgZwBlafgAedKLBnwa8gg7r+t9Uc+UQ2FBZ/YKfsnnh595YYYWlqP
P+UA0pkJqp6pAWawvqnPHyk28yqP9B1sZr6HzxbmIpm4rvR7D+YNBl+68RsE5RclnCt3QkNP6heM
DKrls57Gn93Nl1jsaiTJPqwqUu4wa1zmJJaJ0TLmxKLEFhGiEFqnK8BbENB/wuG92mcqH7jvhCjf
LYpuM0amnreaD5xs3yXKTt7tAhMuvRlsvukyBfz3BKrG6+2iwh9IhnWuqlOK7LJiDJiS9KfSaGqH
7PUS3rG7HYklZ0bGOKgae3AISg2DQ59cA397VOgZGVyjoDkQWrHiTOdIe48v6ZaO03x15d26ci4z
6LpxeHIx8oHI3xu+/Rigy71O+0nLRNgiXvOpMFMOzberlVxWiwdWYaA0r/zzn3MLN2qlr9ywCG01
XuipC3tFBBSQbqVMybzuBtnoS396mdkoSwXTDsQ+B3OuFLgZwEz/LwrFcx1JEGixruau8Er2AJRR
1Y6MkWNJV+VC9O8+dItz9qZhiqNir2LJXLPlOZE2sU5kXth423kiRPoJqGs7oUX82CfrPRACX4jl
q2WgBAOiP4xZihuAvBfSzo+T8JTr8suScD+Aewf4rKeERsDaRmlOatYx2XjvgNHz2krG98QJTDJ0
IND3euEx3a3WiB6vYFfMWzDGs57h/dXr86EqofmCypf8cFxKEyO/Qe80Pz9fXQJJPOiSdwy9uiwe
FdJ9fpFSUrKtx8FzQAKoO5nWp6MmUpnpOny0hogv6OP6YzDJPvYH8AIXJZg0Pg8c2XWudzOSyCTL
fSZ1YuWSQVQdtSm9VogSS3hyEVjaPrfsjJ1wLEcvSdCSeJhW+uiJhPTrINYKAYBvr3Vvkdnav0VQ
f6muKLk0V4AI1sTqF5UdgDEl95R9MxhqDJ0Qgg9Dwd3jsrLNgyXnFrkH1SqU9yJ7cx8344a1BQ9P
sPxpajhLmEjOxuspKy3notb28f3aqo1sMsMysngefmkNXEEmfsIbElkFKXfh6v7xGAHkJT0weokF
mlZu/ZIltPYGkQ3UUlxOlX58MAkFfNQXtyuIGaCABr2W0zTy/uQXZsYeq5ukYyw7s3EF1qksNEIT
hoMLOtb2HJithEfNlU8bhvNHEgY8Yo2nP5x6CdoC15SvWI2eTX3p+LyK94rV0QDIwbpw7/z8bRtD
i+izYz+dSy41lcYPqGDSnObSFkCsWaWlPTfNmjE6nKQnMV84tkkUnuJeQGim8UXUSGsAvfXfe7P/
5nLNyw+uECToFjo7eIjd6ENS6kNLwU5rmgTD56uPTevH/W20c8WtT+fb+0htTDNRaYcYdMaEjFQv
bjT5uPQSL1XRGb2RynF8WaqoHQAlWmZowKhiLbf2oWTN9ERkguBarVEoaX0C7Lw+pHMeExU1Waka
5APPL2vZP2j7f4KBEu/QUheWmwX5tRW9nyzLuPRFRC95RCXpJ6NFoa3eUv2ALVW8JlqeVsGUOnLG
ajl4ltiUEKOevL4Chrb+d2vsBIs4QY/PIpoWxQzAhdWZ22TB8NVltZbTWqlEWZ/gH5kCr19Js3cw
1Io6vITWRMuN9E2bsXhwSarQKY8a7ROlbkcL1b7dX8/WJiHcMC2NvuZ4zhrjHNNoIfo6lK6gYGQ/
7WFpCzj6JBOAXLrYapptX7DyQjxB2JabBxgQ6L2wmAz9W6jgZjCupgts2Pd0Y50F85b9O1ZWYnD2
shE8gHn68ZAi9Ccpo5/BrUWUY2vL3sJoW62xXqtfZTKjnm5GBLdcFvnqIobGjPa3ZDjKReKh524z
3PIFO3WpKaUO4h6Cc2KTbopgmMG8NbMTiNS33EoB5IF94CvGH792MCtis/yJaITTpcaGMNzEgnFy
3JPyMYYqdY8/yrpz0Mz6XEJOibpGm/EIVOylNz1CCyRyiXu/jXsAflBqWju5loTnRQWXKVxmO+pw
zjdtPhuD76i9erC03Bz2Yfcba28z4RfBNQ6EgaD4pXdRQnzd6COqpNZqd1Q6pkCkRK6DdeG3zj8D
T7JNDGSIcyj/rXWbJQbWeyZylVTFb3S5bf5ugpWbnj7s0vNUgrM/I0y01phcQAgkClVwdNMvKTaa
Tw444aMdvHmdXrP2UmUirhQ9DkGoZVZxEiOZn89kXHQfhpfQDOWZ6P2mrciA4+RV73ducgP/5zF3
WT4ZmyVH4YkrCPPSWchId6hqIylGT9/z1SDuFDCflpNyFTshbn4SiyC62csSyAMCOCwV/mslbhLp
Z8p8hkjloE9MsYBPsq34HGNGrFmm6EmeM62RLLPXoOx3vuvLXvzRmdH+bmFy5/HbSR3YA8qCaj5G
8e76BcgIuoDg1fewPKJKLNsSxdVX2c5g1CFVQIzZXriiSXdd83HhSKduWlUtfPVkLkuihlvBD4XH
oxMF8j7u3asDV5jj8/M8H8XCwnHyzL1GGoJpVQhFk1wILN4hOMjXOVbkqCERGLZGqhnAiBtdJ4k3
ERqIME73NbTMgAlkyxpleyM3XCf+zgJPNmaMpPVcGxCQlUu88rgRmc8PMNgoIXEZ7h2T1kcW8bwg
qeY1qrk2pKIPuEev/eEcS/4T5v232sjaJYooOexItHWs5TOIgdII9PU0rWuEJ3mqC6kzukjxDk/W
52fgnbX9aQWCbw+sbMYgBHeTtwSFrgAhxSHXYI+36NyXZMLooWbMjEOKkdfr1ycwF4/8vykXOhxy
fjEY2uZb/9v/PqjY4hUm4RBsAXE2vv69Q2OumiEM6GmCKAQVudxIskOrsaViu3GecY3ebx8Tlcne
QTmlVNIwpTfpHcaCfS6aCPQwmv9BlO35z9LFzBaIvccReo2qmCx3IUBn5iWgmGHnDZa53vuC9Gkd
8IQ/A1qRB7DWpjSJyLZERRuNPkzx+oCTlsTW94z/7ZiGhe8kRLppFlzx3o7r8YO6bS3j9JD6gAba
Y+sa4YAg1WibniAuIOHA1AiVMmEx3P2QdZztClGN+oewVRo9QKIk4KU8AO/pZbQFY87zwFKjBkW/
LMOVyHYQV57GFKBJ0rPtXP+69KPyLoDl7XDRThQW6pZ5nCO07IOfQuIElx/Yjtc+XzszMMzpBaW7
mLQSVX09fpS0JF7Z2Nle/0rwFt3ioaV+KqFZZqVhv8R6nHE+wIt4Pyyjar5FsqSWonZUu/ZkeC3J
fnTwNVyYHLa7dVLUaZNOSJ+C4huwL1V+cHg1GzkGm4PXQYEOvn13ALz0PxEGSZA8TEYY4ODBsklo
tBFcVrwtq2BJ6H9cNVNxu7OPbB9tEFsYpH8wGS1L9XGkFkdxwrDS3In17VgSrAunuowUbzV2ILtD
cxWyq1IigYPChNoV3DczLIk7ihpLejLca+A6vR9Qh5qZkiQLHLKru08OTTncdFeeops14zn41yvr
GgprttBUX4VTKmrmmzHt61aHgkve0+V/wPYZ8FEuwMnOU0HSvjhJdsqU6tMuXjOHKZ754FHSydPg
jMb+FjRaBNaB8/EWwiyk3Pq3Nw6sBmOU/8mfk7OQHTP2pPrsCXrGiEU5rYOWOu89pFrz4qPbQj5c
qOJxohfiGLg9Y3LH7EWGfYrmBit5kiHsnC0e2OiE256pCfSGsUfUkfVAcZ4fkML7U83xufygIiFF
zvQ5Wgj3zVuyNJ7QFDVYG7aYf7XqWK19gSdaSPSbKVXFOZcvc/fbinBvIVMQM/3G+KcDk5Tm+SjO
IyUycPNFavcxq5VP3SWwm66W60zjeI7wMtB3Vb3CHyx0GDVnLOim+NkDvcVe7JGTswjvJlDWw/Er
AciF6/Cp764eG6R6M5KWGaDBdJPKKxqiBG2TY1rmum80Z22YVBiMdnVt8HYiYh/tTHsCS7Rop09C
hD44uWGczmTEc1kKxC5LjZjoL7lgm4T8NSFjgFuaEL/r3bLnB/wmfTtmscN6RMbiE0rNhDZgGL2q
D+95d5LD0XJOYZqYUMFdt2vuFwfzs1+SIL0jVz/AkM/C+Mj91PIFuvQfZahRBi5y5/6ks23BQ48j
OOn/V2sj8Pa55tI7N/raYrQuqPdmO+zJsRTzH3s19XXdkQYBFOj9yOjDhT/Sf91d7LrFgDL5eY8m
M+JmwmnmZ8nNqEKgmTqIOujtLUYuOEXvN/8beJ7Wyol0bDRsQnCZfQGzszdjctk1HizNllEPmaeC
2mnBaFHBsrPgE67XfbQ+CczZaX//T6HF4SFsEbD8MwewjeQ8+5JywLXtLaRGCNPRfZcbHAdMyXye
FECeaaWc1tidENE+8V/kRm5tqJR76MGvfD+KCFynoKVNdIODa5cgvOJarsi/44vWoZabhaastVTG
OjV1bORW0jJP71jQvprWsRgW1EJUSWXfs0tKJH/DRM36mq2XnS8gXuZaylzwMRGXqgLRnDJ3EmDm
5N1WUAefGyOrvCNiAbsCqSrzHFZqT1OyeoFHyPCa7FLxR3qC9jxNMajwJ2n+KFabxe+RTusG03ZX
1gm2Dw8Vjvz6rObjGejAdc+zlrGuA9aUvAgn2FtBCdcG1YEdpR1bkDBuLCXOF2W+Qqty6z2BN3aR
z23wSAJvo4LkL9fKEkuVgj3FgzWRX71qng1JvV+2UvdU6dUzyX88Y/F0i2VpZr/odF0WYQwDUMD6
QgYDbuuXG/jX3M0qta7e2ufKfB0tmS0hSIgEnX36YHajQZu5Ynr+XIOGlyB5KNbBs2hIFSgiVpps
w0U+CyS+ZD4/Ki77DIhXbrYpSxP4q4M0nlraX3/xhaE8/GKH68G+mL4J8lQbfeisUsShKbMv24/B
RcGt6oxBmQPEbfLkJbuK6L53dkYPUWQv6VaJb9YMyp+hsjxoVENF2E5BU0BOT4Ru3uhuKHwxtN1b
kkK2gPruH9h7+ikqWGWTeoObqDGluT/JjAETjBAj2XOs9NRp+4AlfYY9L3xwl5c73mHJC/WTJKqS
7Bs7u+4g8LLdkV6ELzXDj60DiQLCKEtFIwGyxQhtSjbyoJRm3S/9iJ+f2EVTOCtKCNzVe7yRQp+N
L4jcUbkGMt+2gag5vZWEwTYzqGj1vfGsg8x7r3B0RICvapKRqRyvnn8ZtoQ4329LibWcIjUepeRE
XCADg5C1dqq48Ngqf5qhxQcKq4PjvZqR1zLP/FsRRxx13+4jUF39NYBgq4lgfZmLXGTJB/Q59eTC
mSnyVXsE8v5FEu9STinfDylPjg0ITVE/m0Ki9Xj9ploqUwSs1+nYiwjKhfNHyNOvk5brygRDgK3w
C1imnrP03WkXuQ3TLnOcutdLmyUK/r1xZxNRS/Jy4xXPv2WzC+hujWqiEj3d0avU63nvacP5pfeT
rkNGTGHWfPoxjilOK4r361Y2sPzfPJq6VUPdX9umt2sPSbYa+i0M+is+D1trNR29oCrxpAFw9RTJ
WFmAmL08IADjcfY9x76rob9BwlgWjDzPlobCSutpWQqnriFkEaS98RJBhfZFOg8rowK3Nt0OiKgc
qoDwc+i4ORbSoEISboBoZHh2dwaeuwW0mPClllfDt+F+2DFOvrV0z5FvxAYLFDgcAdRibqgZ/hnw
J3vIUy6U0zgnAjXYnR9kV9Iu7NMuEu8jWXA5fqS2arEe05TpzqawmIsLhtrMMMp52TuJuwkNbojG
oyIoZe2RWuSBv0RT1e/jZcHfdK5o2G5FgTPZfHCgNxeCjboS1x+zQm2Sg5RqF11YFfFzmNudzRO2
kthe9ZQHihTBIPG9ayIMfZrABQcDMytBIxgbzG5Z0fx9FMfKi6HFAyAaJJWzWHZev0VXnyjjK2TA
RtGJpv/BC6wrCpHhcIVgo1gzpGGWS8YSXXvIfiTJAZA1W2wmR5MbrcUDcPQfHsSOEv9nnug9QLrr
HvNgzUqDVIOxLWo3gJb9LOnjuULX8Pu59545NBujQtxHgW+VReRYC12cxGVv1ZlP8/aH/yolVcZD
40rLC5m+YXmLoS8UvrOBtvQ/DrTJlzNREySD+gfS5dRHFl1R8reTwbRFP+I/ftv9VA1IZrhmMfQJ
RHAuCRrU7n8YzUztxU4etMQQvWcgRQz5ijKlso0ziqocpPiIGMj++cd8Ei+9z9L6IbIRRZl5I8M2
wtyggP5hdLNTu3OCAmhT49oCgdEbMMvJ7V+szqUTiN+VZo5a11b86geTyfYNj2kHWhs2emU/EUPf
wi7YPK4e9wsWiAwpNKbcfk1eV1nJ2cAYVadFOzs22z9cgKHvRX3kW0dQSHFlDxthcbxjzbs3JoNe
xzvQb/t+qRiZ4uujH/yCCCfejvSnwewPVPTA2anXpos0AiRIbc8T/JI8VlEaaK58wjyyGD1ehJzo
u5Ne/h7Z/hV2HOBYGXjQiVDaJ5RMrVLaJOVhcXoXYZQJNWUQzp3jocWMJqkCZjhdCiMfcCdYLq98
mNT8GLd0J+fsf6L3Je0yTCDnfTGQawv5d2mOyFIlg7tjv68xdYY1DqiREMYhHNfhP3wpTlrgFRtX
VZI8MPO5DaOmKKe76fJcXXEPhOClWKQMmMxBV4DWX4N4wzEjR+qItM5lNUQ/gp5ZOrvJWNJTx2Vp
UnmgFb7FeD3+TYnylK0EV+dkqx2czgngQuAXJiaPJyPVotI7kBmaRWXvNnWdhzj0JNcyA14c528r
ep3NhIJ2StsoSdVJ9TFKmGR2bEyR3ZK7VFVr+EbDmQc3XnXeGlDf7ui8wQxPjUOuKpqD2dI0bbDh
BE242F0k+3dSPEULam0UTq8cohSSq+cYLrFpx76WHzOFnHNw6wa2/IXT1on0xRyGLsH+gS1o32Px
+cptwy6yXaJtkgtuEBJEINNtpLq4YQYwhVm2U6DP/WM2Kq/UzVO3BrA7Jk2zd75hE3bMjn/P9uK2
/mMLCdD1v3liMQvpnhP5W4PSLqixlsar7g8ZyK9fart+Hc7vBf+gHgJ7PuYlbcrbzX5wczXbzYHV
3l9HGw7DsURvTnVMVoDCPOyB7pLv8UFzezlTV6RHO17p2MFF2K7e1CKjUa5dhS/OLRw2QUEUmDNl
uIXvorefVEC485euG1lU/MVDF11QJUG+BvSlQmggY7ZtZw1toRM+FXwumH+GxIbwsvf3d7NhP1SW
wtNKA3gBmfDlHHsvoz7CZ9Sf8BYlawoNhM07S8kD1loRPvnCnUaKJJnT5i+mDaZ/bcif+dlfQbpv
VZb1T4NgYU3u88ygbrF24/f1JiTZ7Z9saSBJGiA2DWM4Fe4elBNWGYzTZnzE1Z1/okmiBP8Gdxo3
rFX8KAbT9NqlHoWW1UtU3Q83FEt0goc92fa0pP+aWkS3nknsZBQL3hA4pCo1iJAp9Q4IPkTbR60a
p9NA6UxinbTbLuYLS9x896VUSHMpaVrKv6w030IqqYO6LdEo7nkoBcAGgdyBr5Rf5M/eUtzF/6pe
RI5JLIk6g7LQDaHq43DP20xNHEfxrMy4C493UjL88cQpCgZadPSAfHgQtbHYNIAH8+w3pB6XuC25
QWnCoSdN+tSItQ9yL8GQs3wFALNKdnIkgaiT8YyhvqPFGUz8Ivfq4E6keUuNPJfOHWOe/fB/3aVn
Kc2NWYqtG6CJ1dh7tLC5+5OJkxpxlQqA0MX9EtV6R1+loDZoUG3288fvDCi1FZuXQzAj0Zw5qJWi
66lZexSNew/FAFDovTIJPy3/J/xyGEXQ70TPbyqcrqys0bkIVfzM0xWOAHvLc/vN6Ui+am8TD6O0
WRvkdISYjlTztmP9KJKyS2RweoPMMzuuGS0wgnE1dTBXZJ2V644JtOMX/hFqAEogpd/FOioQCzsx
7fAIsKwYmfkO9Nxe8FxO3qfmMRSaT7MvWslldsc6vzxF/Y5542ahhdeB1s5SeKkvSTy+WbofVeXJ
QWQW/5lo32NRwKnpDhoagIMkgKDR+BiRXM2kASVhEArzTmrHFgeYJADoL5cHh0fi3UCACoAIMsJO
7UVS2gyI/90x4D68uZz6Zej/kLXph5PI0GmobfUKt5bB9nkkgINBIxpqtjvaS8TwgdF2uXrLLAPN
7FDujat1LY9lSYK4u4FTtyo0Ly1Y6kJPnzoVn6BA59nA1d2tSbZuZ0vsUHwGQGfSz32omtEnh1xP
hJ4Ip0zA9gNr+a1J26HRCeqhvuLFIixXq/2fqqYKISTJXOKWMl5m+vU65keOp/GyfbmLv9i7IqJR
a2O3wxgIrHstQwuWPI2H6/mfnpZA7MvYso/WOk8KnsEZACB11tu12Ife9Tnf+Uhq50fswQ9k7XKH
kL31y9H7/nZlcAPtgyQat/T8Gw7817xoDvFJLgb6wY1c5FSpGZkCqdWw6iNB39Pr7WPWhyS7iKU3
ovTcom4V3nfglKBN9ZIHyVadtTDDUUhEl6s5CpMpGqQ0ibKv/lRdkmThmB5i/F200xjL2DBVgwPY
JIIcOq951eVbLGijUYytCa5PDElSZybQnSD/ZaXHxzFYQJzNfOXyd/UXlBDUNOkKIjnK0oh8p+Cn
Qaj1DKpE/gO7QGRCXYdsk7EUxCBACEXK7eoVx8x6TlJ3tc1oOJvtIN1Cbn6Iblhgp14H4S39mmYI
B8Uqh4pLyQEOduKXOtr2rNpAF9hbgkhL5bQz0iz2FkNtZg9tXmJchOZdXUAsF+IBz5dTQybiHeh1
pmGjHboG39TIltEAzCKXIn4EAsJQyl065ljfDqtEeQW2P6UeEAMb4QgP78xLQnJDe86ldtiKI8YL
Vkvqy+pI/H+9RFuxZTTdUUjJiEngxePaYPNLr4ybyEBMeA48QxtUxlvwckb9Yw4vvxj8rO0TQTMV
7QAH430AZn5k1ll+fFT+6ZM/VQANBoEgyRhGybOR91bAxDi7iANxJmgyeVm2Qa22K3jW/XMEsAgO
ian9DQ3NVWgvDhLOC8L1ZbeglAgsx3b+N9PCIEmvuH731KjfG4Rla/2pcJYG6U/96opO/UdcYOU1
4XxCySmZvlkCNcp2qTETD7aVw526TeCTj6Jd9z99ykA56tW0ynHMnon3GxgTr4jjrVTzljLioJRf
8j0nGe66e0g7GwY+4gFdhuMuM0QH6xvtrhV2yzoYcUV+fBMesARTeUcjDnHgHz61W76gwwjHMnb/
TvuIGiPvcWVFucZke19uJzdMX1V+1mPoEx8GWuUbAh4MXwGcDSnw+SakIB29YIWgbfBYX4zw3VwV
Tr9rF3v4YbaFTnEM+Aq6NdLRkEHC+LBsdlhkt+ZnxmsYtLoeK4R5aIhhlh3Cr2/TZ5f/XOmUfHho
iS+755nuVGswbB3JOsxID7yU3QTQT489OpqR2QVhXFDWypjSYKcbHKLDphP0VN2zMef9o6/R+353
IEsMxvAME8Q07nAeKe6h3ObUQDjY0u6UUkXGKCLXWD9joV1kAt3/sVTUUseryGkz9Wqw4OiKgGj0
s7aghSMo6Xc6smW1G8fQHhE/ceWJTV5iv8sOcK+pFDXS93OMhP2nEZecxmw1zBxRwvPBp9fl4JqM
jpx5yPuiJcUFHzNV3dWjEYF2v3g2KP2u9gp0S+W36hOkrtcM7IVMiHK9dCNMat2WUZLHuKVHNTK0
Xe+kD+vtnHU6Jb2pnil+uxZaiQK8g17BTcExwPOgWogUmjco/rZH3tqFv1vBwKI/0qBAhnqpWLRx
BSweN72PAZQh9A9PBENRcfsMyPwgQk6aO2CC7+eGAoFlyd3Rk9ia1o+IVQ335fHB7BQe8Hq4+jDq
BBnCtLe4itkbqdt8BiEo0ebNEbNANE8GPINCNrtJEI4IORyMo5eYgumYTqD0y0rZAlH2VLl/MdQc
jmd37BIYRHqjIw1zcm6W1tr5hoDt50mv8zqInCtGY9xLnE7/EfoPi2YMdLOHYu/M2md1V1QDOeRi
+GCPd7Ir6X62Ug8lrh6BppmR1h9ryR//faoS7RCBJchSWma9ARMv/raJnJqmTcqryQyOvzUFB50P
aP9J+PKZj2TeeIAXglekxuEN2GnGLMniT+KOFfWXCmwGVo5nRWYvyHsBtSeM+k8JzARQuNmGY13H
Ej143omYN9o3CzghWv6qPDE3HosUZ4aUxSDrQhgA5yuaueR4SJgXiqByQx6IGAJAPF3lkmJYGpCX
+EddExLPJPSe1MWg7qdRmNaMNthKGuKXW0cXmw7yhgeF2Y7v7katDmaPfZMP9676CAJ1yM3G3rl4
6RxjozGYa73P3KnX366gz+5ayqFQPOeXbe5sbvnldW+2dg9XgwE2m0llBhFWqY03YIodlqsYGjn9
7g1YSe1b5T/HofPArjtceN8YZ2dEcfB/BAx02KezhS7zI448vLRTWNMmWT2cXOp0OlrCZG6HRCz6
ysmbWkgd8ULvSatQhYNRfYs/uA5zid8UPJb1BTu1avz/WId39xTZ+7xr651Mrweq6vf2d68A1YrB
IweAbvqCAXB98crz7PgHxIdy+Y9+u7NRg0m2pGmIGyg2svgCX+tHSnLrnvkUyEfpsQHrPECOkTSm
an50vUW7BfwouZFKKNUsLkypvrpfpxPDNx9+TbLeCec3vSt8A2uX3/OIeRsUfu4PKVMNUt17Xr6E
EdywyZEhhW5sm7Us4/GaQOdrvvTIB/eQbnJmNS3pPlxlYsfNVFYxuq7rHafW+UW96xPyAPG11cyd
odTVSRoxBZskDSUAprC/oS6do6SK8fRBN+7cci7HdWuX52m7hV4oWyKUwzabOXZ3z3/wKSrR7J9A
5mmQNN0c1LRBqBb8QZmts1iwNbP/Tbt5eP+qACbtm0K248qMSHRuCsmQB83zDuqQMuD1zV8l3bSP
uIETRN2qeB3luht+OKoBIOFEDB7RfhMIb2nEvaO83SYKnz6lo/YtQIlpdlYxNk0ImrK5Aj6NgYyp
ksf1ASxTbX7GV1a7Emn6UcnPTeUvM72r2DOoyJyybAfpT4qcTtg0ASmTXhxWzIIAGwym8RTmLyYR
Xh3X77I1LmSRlIYAlgDiN2EOiJ4dklKKO8/YFpuibk2lSVSLwOfinb/RddWSoyDKNkQ3lYAklKGF
Lebs+gcYFugvhz31rpUIR7zV2Cn3awjRFI7dshPKIYMxHcT9b04x6dnTVjSi2T5RxR8EN0hhn4Pr
Fp1T9CsD38QZ367ae9tDE3m7Bdt29N4nJV7Oi5nC/6tt2gHPKoPeydkNG4dJ9l3vqzdT2StpHiTj
hb0AcsZ69aFONtk5aT/f8vQgTdn757KlZ1MeJSOPwj/lHqqfZOqMM5fdeRe0fUpT0GkwYapvHaZW
fcu0A4UDW3ZN6HBW4vZUdvlAsSjt9uvRoDJxpa+p/Dh/3Jk3Ddq+7nGhALYKWWL02jD2PEk8V+Im
WC17oRvK0uKjnuiqRkj4IpGtqytZoJUpuvIpoGcCR/aJJnnuKrIcD36v3XnbnqkvCPqQ9AcGjgBu
hp9A6hzaJNxGo8pLtnXRZLvs4IK7Xen4yxIq97SH4KqmMbLLgWql6D/LGwuFZBLbZKsXo8rTRaqt
OF+nsKaFoZsslue1kyvv45bt3XJt3z+sAvFuwJ1HK4dY+GaUP/zsl0sqdaP+tJDmqpTOoX9+oLYd
LPlWVfG5nvHYJifFBGMLIdo1fV9b3RkL6+l5Sx45uconppaL7hNP2ma9IrGdpWs9bdlwpnW5Eoxk
jwFCR85IzWuiU+RZOt8M5PlO6KM3Bx3iW+yLh/pnCO4VT7A9gQnNUhgimJ6o1QJkV53yrY6DwF0n
tcwi2YeCLsWc+VJEl1S+xf67dm166Duk8zLKV4x45oDsm9be7XLz5qM5C8aGE3D4xPBeS1tZ8Vpv
7OIELvOl5Ey4hZezIuUSydK4UmdAAAn3CDig7FBkgnabkohaaZ2NSRVyyjCkUAEVpROap7p8kb5w
Kwtl/hvRmat//VmRkfx6asc/O2Z+S98IwH1H8Hm5XrrqF4I7MmziLbkTTLtVFtAmtu9nT5ehebwk
UqItAF6wyYiYcrrCB6tZrfZnmozB73tboDuG/JPESz9vgboHpsuDlielgJClHHcxgkI8xEBc5i5B
+YTUp2bp5tOjUhtC/y3oCW0yYIBBJH5rGeCghH75NctInxXowUzLlhM57+ULPYzwvwKzftSkBen4
8Imb3WHvGWvEyl3YHoD+RJyCwsB8f/6RRj9HtrfVCGU+OBvHK8wE9/0rz7Z0MP9Ue0BRlEJSxTKB
cwzkSQlrKjzGVkV9csof3kml2rAPPWAKTTPOEXNWxoe6Dm5Nm+W0kWGiR7sdnVC2upylSq99Qpin
noJ5B4dxxp+nenS6zsxpm1HJNzPP3qpzCYzus4z6jN4cbMd7/OjFUiwn4o3mbmOMKJhsd4+isPJT
rN+oSNSlheOvuGXwd55nawtKURFSK50MNUSmthnu49VoFGSnbfUPfdd2tLV0D9tK3ckVGE19/kYr
xChz2NZ/RpWOfPcA9Fd0Q339R6183IAQ8fR7dTuuKf7lFwXkgNQDjr2uAdCkofUwtsbRTTyzqyKG
51Q64ZbZGDpqIbDvyxPPZLFFri82+8MK5S4N/H33imRphVOpC+GCLVx29jCu9ISNNoKQK/1XKK0/
j3fmgAXR30XgBpU8lkaCfraIeAMH0BrvpjpmAlhytnw1j2D6P2MhaQEGDnCmIqI1F8osDa+6hsWU
5aEFY6NQ6rFQjh1N/bdEf6YRUTgC7UXa+fPuhNgLc5I9TbTaMDIk0ysQug3QCVZrmC8JHeitHp0H
rYcjDgR4q6iE5NFvb0v7o0jv3qLv+YB1CsKfaiPWCrootwNVcE9Q2d68/3K/SpiDHYXKL28f1QDA
pu/AdivzriP9lROJRtVHi+G1PLdLk66uCZ/L/Z+MQFKkZiCwyzNHLQLvNECOox2slyj2N2DH+Be2
gyFZKz/4uYr1DHMH9S58vaj5cXNvla0/+9vHjh7nmvIMIjEApZ6CPJqA2lVuSWNKktp+Y2DYbH5i
MLCjdLV5TaXJD5csAsEB1hYTD/Jv8tEAoSlj6c2D1/Vw1BSFI9oPglvnuxv+hpRntXyy5YJTyfEe
MXKTz2w4nd2isdQtxsIsQ3pl6tk3XbjwIg4knHx1LPZuNQMSDLF3uWfoUZBObVEhls/lYjuVofSp
9h/P9PgKrTEBH+ZywwhKgOgz4Jko69EpZfu2jN4wJHziO9BRKof+scaFrwTPhbW9OmSBYnsYqdEm
Sr+CR+wZzObiqEGmJkIXE9DubYQQw80z9COHBXsdiH3xxjbv7GCtbw5SrWOkBghW+pw39LlNO6Q/
Gd8jAYP5IOQxS+tvsPfRxORKOQOrAJPNGt1keJZPiv9R94VDlq9xXQfxruxfWUe5n4yppEEDKDdZ
10KnItI0bDyOz5BcsWHrI2JMa5+5tpSAupmuN/KnanVTdMeS7xkYbDFPJlzIfEYyMjX091HRptpp
Gi+hDliPF0VhFBTdQSeyH/u4mYpBmHWXd9DkUsIaVidJPaqwY9IZTgJxIBOUj3jPESClVIupxH8L
xGzSYVCGLOXTXnsizgmbzDnGgzo/iBby/R2l8Iap5Hi4zP0frGxeKPlIFa5mdjcEWPXFUYMlxFR7
jupisjSCNypsmUhkUgBmOykXpUeCjLOZSN54NeEQciSDf/s0YRyKJ+M+BBoqRNgtPQL53gWu68WJ
NtM3RnoFiw5dppH4EadD5vO4XfjkxCom4Zg0pKgz7/WGLZcpP7y6nE5NHmR8akiPf5w3XSSDJ8Ck
8JtdCxzhK4LOyCeDmwtqeUSuNbDd48yzKqHdH4ERwpfJKK5KXW6uPmhy+OhiFYIQEQsY/8WSFpjv
oaI39TzFXhIRZUHr/fj4PhwH/AAI55CBj2tIf+UcWG09fAzG9qKYXXVY6Jp/Q6vwX0tikDZIVcf5
Bnini1rr1ilbDYkjZCG6dChjHrq/auhqlzLEht5yDCJtHJskCIDPxeCssFaSb5pfzznEgc8KJDZV
PwKl9WcZEZj2OmnITHph++/lqxODSTo765z5MnmvGDVg2yRT7idnUl0lgb6baVktLyU3MlCig4fI
p39eIXdpw2bkHPdD4+MwZFFs9spePj3KwichBXJLiBQq7s4lRiOLGHPJAuwNeeY7d+MxPMzJ4pHn
kUGiHKfZsP/TJ7/MgQgKlmzceGBMVoTx4aM4uiIOy90wA/ozUkWo6qEXzJGyRrVanj7oNcmBLZwh
rTTrJ8NfQ/oheafYBGhPZ1pj08gANgD+JENDGvQcE1gxoJLzZXiUEUbNdRZYxhuU2HuwwuNY6cWN
OgFoq6Pf4AoGE77zJ9gZNVj6M6t7fyjKRjLUA7/nFlFaGrfDA/xwnLzViCE8404KqdbxR1MgwNyD
yjw6bO8YrSHekouO1eCcBIsS0hh1EbkZaV7RjlRgDLIiRpWAKfeA4eeN1XNqQD5QWatvdyJ7/i7R
+KJJucLiL6ztFGkRDvINgl8cyzMxfHMkbsJoG+1Po/8ys9kadysJGAqBW8KmLgcOkWZdvWqgGNDq
pyd3siEg+xJIAhgL2bU9Bmo0D++It/PaH29Hk9ni59rJwwpBN19pnkb0lO2TnKjVI0rNHOr/ue/i
BEwubqBHBI82IZQ5jYJQgA0CiNAMvm3zT/TjHapEEWKJjM8G0Z23e7dezpxVAvT7abvrXKlysCLc
7nyQlPjfLWVCOOOQAVDRZ1yrevym0ig8+ouHAci7NNBikaelOx9tvMGKEtK7dwqEyzKu8Lsnnqe9
qkk9MGKBJ5ov8VBARdWeVKk++nEjv8QYrQYtQjyGjfixADNVifKsPl8SFNX5P4JvFooNs9E0eY3p
jsLZqh2QU2wMnTuYhv9pkMBy4C0ku/mEGbWrKf/rpv8F6sSqjgdSTez2OL0Ct1Gwi7qb+vBCJJnZ
nwCH0YlOuUHMONAHuvPpeYv1eM/t5/8RdCqb224wKDuAsj6B2wCY/8dKd5ckxAVVUfLLObvfAfd/
1o1TzKdH1uE9i+CQ+ohTIAp/DZeAEC8M32SvuVdBlYn8BaXGzxLci+oiddmLoPtaRIlwcvvcVaZ6
/GWtw0ZOPDrx2Y2ARcsz74KYoR2yQVoAlkByP1bAEYIqkaE8nlgAhFgzi+ARyjwCRQDYSk/PP4SZ
nPMFuluExekB3rkdwpmw90ReSVPPaEHSVOh7U5oWg1Tx75/y58FF+BiJ0wYXGh7V2fHr0LFi3d6M
pQPqNP7G7ecrSRLkmyJpWO6nZbHiLOkBCHK4sqgJqeiKlPJjBCZR22Dg9um3V6qo/Fpx5hd/FT9j
hSIEIvWSkmdof1TNfEi+VEJSGh23pJ6ER41xx9sFQ1pkP9I7kaWrRsuvSA6iRW+cZvw2xUU+iJnq
Hs/5O7kSDpSzLtWa4RIcX2vLP7zuFt+ju1zoUU8sZ5XOQHZs3Ie7e2gtn0f2KxqzjpgG2R1AvrY+
k86GN0Qk8Mcd7cyqZrmgiPgHPro9LQcqlSmzollmG/hnApJGt2kFRBL9biPGxJjGBVWOCYtK4vqM
ZKVBQWsVZVaGhtaYhmqaPYBEBVpfasElDkovyFWHyyaujoR3g34YMmBOIAQH6mXXLzu3c7lV2i1p
TtpQLRWqfG09ooPM4JcwzwS95eZmVEfzd0rUGezrJLW8eRi/JX3tu2a8O25a7azWX6PWOXqtyzQ6
4qu8qNwD2IQxytd2K9rbPcn3GzoJ9VUx6KD/L3nx8LKJUCPvOQRaVRJv0RFP0+KG0KF4+KE7ST7D
Qzrc377+3SaZTkitj7VXlvHSqGWaiqbEKDGplESEMOuTtj1sUTbKoeol+7/vXsdV9LCV5T+Z0TYW
q68uINH6Ve83mYTabyVYfwJVAGRA+9EoXTWHxlpfF51NBpMJDW3I2cjegCwXz2CAp/4ysoo7j3a3
AtIOtU8NriUeBBSDdybNhnGEwJECCPHbgdrP8JhaLwUCH1iXQ6r5RtUpBte+Biyt7w7D7XZgQAw8
95pX0/lq9ueFnbs/CxdB+TGTaTWsvJhqZo0HrWr+7BrDuIdGdOpLn8UhInS4199iw7MZnZ7d7Du5
NqBJM0iDuTpYKgfQDl76DyhQ1p39L00LRLrrzD8jRIsHtopzD5zq21+gvHR9ACWu1wNgzsFvtKrS
CU5S8m3DAQZZ7lf9772M2cq2zU09P+oi6UKkjS4TgXH2YovtiErNlZCETdp7M/O2JC9xdF1O/ak7
RpURGUttt5ZQzedlipBRF+u+N7ta8p9vtHU+TJaOHGJX8zN9Isqu5LGM+r72nXZDuQwm2rdqzEti
h8+mPLCcAH3RHJwZOg6M/ab/yX4tCuC+OAmz9XiCjSCJ3+i34AWqaIcs3qV3qc9+w6aTnml51T2G
Vm4b0VTIZ2l1T9axsdfN4emtmI70vNTL/O6Mdbwi2H73CZZPVycYc90mYvIWOGt8LcrEQnpo1Skr
DHv4U7r6hrlxzzt33+9gMqUlTU7cqgsZloqPStMzgzZEiQP3fB44BemdUtBQg5JUGeAgzzSTN6sT
j6aleXQt7+2IOV4+kWnsnIZ2UwfZSpSa3ZHaR3MZmg5AApONRTM0vIzgX9SrbVtlqM4o5bYq6qnv
ifpMb23SSRgpAGCFkQMk2dnJ5OTK+MKGHxqisaxtMKEt2uoldaHkIWut9C+mThGsG23hBy9bY78K
eFHqIg1duUVjRkQuyK5a4BWSBLl+s1MRpPjxDdry6F4ihGGJtj9VFpuyFgI175fWjm4z5CXfjvG4
vewPxKJQ7z36Dxhikj+ZMxsjuzFYwNG8K4sipW1b6YuTMy3JAWLDDwaw/8Ts3+klxMA47FUN3jll
WUDaA/WsA1RY0uLYr/Bo2quB2JspIEv4umPAiCGq4haZsSjT0tgLq0fiDTFdaB4692W70G8gjLRP
ieydbxz78xJeTtV9HUICnp/8UlQjRfqJgnR43XS+3YR3ENevC2nUeLiedNydqS2Ta4a8b6PiKnxu
ZHPc7VJmQ9lxDZXFuDu0cFH/MwuDhCU8krH/ES1WdL37VfMV8VvpdwO966jVTZYx1QrLNjMgg3Zz
LSzc82rI2TG8O5WOI4hVpCvCKn7FANZSYPZ4VpBrP+hCamis1WQYROR+Dkr7Dlk2rPaqxyZm/arw
byzMsuRdqzq9rdflAx6aWv3JFqtaj6yEDpIrnuR4kwhA5zQ2cp7Hal6v0zhr52+sOWNvAldufPaU
dFa6livgMLcfhjGPD/+dS0za6Q7eqpOE2YDAj9R1/6cLlxsDU65+l4yRt1c7X5skz018K3GQFzkB
abGiWGin8cVWWXFqET82NLkTiPrgIZ0BFyNDY1C1K31zgdRKJovTsK9u2JQHGgS+wSoPQlWCET7b
cNe2yYE01sIT+CfNmui8eY/vbB0yjSXgTvYUG/kdxMgNoUgRYlDtbhixj1o5+xArw++7xQpE0Lk2
SWNWGBJgntmEZONSN5qyEkI6rPhYPDmKheJW0BzzSklO2hFZXjFxYhyE5h/+55ot5CKryk353IGa
lKidQLicGBtom1EykTqyGMAiD+Iv3qBkA8NKlGUQ/zJVdwUL/YqEQTTioQgtXg/quGWY16qwguNo
DOLO/8TBsqoOIuzSYzF5Vks/BBkzluzIvfN+vdt760LymnaAlJrZ8SA89j2CitlzPMpjcM7utDXB
RTRkZPsZoYgkpbcquANX5zfIcrAepuBSix2Nt9pjT+qKg8optyaZKOEj+A5TbVvlBpXvt9WE6RVD
B9XLNJlLxaAD4D7CuZcyCCYyWuw4e9mvjx0UoBb0fGTg13hyLaxniRD2NFY4T+WHWKXNxnPIOcdc
OZ0DWxYcCM5k9/n+1jDP/qdKJu8ZhoXLqXJxD4YutewEYQO3xSUVz3C2rvi9l64v4pETdX1ymANS
LH0CHu/aHufdaIXOi1tEaQjeIxn+XjR7/MPgECPluvJiYIZd+kV51JwQgznBcLxTdbA8K2FD1wxm
vPxaAI6P8HXWjSX5nnjAYXut5jUlE0vd8uktUmfXM69+iW8ccgB5qAgYZQYeNrctFWUTOmDqyY5S
mDYw0W3GJB94MbBpMPgJHbsUFQlQj0y8iajrOqKK27KAnbMA0wJl/fuJj1JkeE5D/zi4WV7U/rb6
5VEonWoJjEItiWSYw3ZwzkeZp78UbkCWxwUCEIcJ/vdJ42yxIF3YlKvIQrzGOKMsm5rZ4D/QgdV/
AKkEQhQobkSdeb0iw+gPkdr5iNvVKP86fUaUrLLv/4fFmO0OCZlCw1ts/RWz4zsjXjLjlaAUhMHk
NmIT1/yloI/tM9vQsqOXtDv1iZF9JRot7kKssbzk/+O0Dt7LUUarQACAxymSfx4F6zrx3davluFs
ehEo5fxRVIVrT0xZgOcrzaJ36otyYUROSdrvkIavY6FoLtozj4rYN8LFGYKNAa+btSvxS0weHq+4
gQfZGKRVXRqCpWv/drthIvUYPYDwLt7e7kCOsPJZU2h3crXujYszFYusF1zABbkrsB1nHNDKt28Q
l14Clbk0IMBOXLHlqaI4gDpUnEIOuIILhh1NaMkyGhiHLnrbIY0X5auhhlTTqF6fkIFx601PYSGS
iXkSREMgLyiGu5XwMBe8bjFWBp2xLMN8Kp0KARr94mEm9BHxYLQvNT1dq85kMJtRZ+a1GQhGld11
q/w9K4RBgyU4OrxHLSXJ87WD/kLGnTm0tApRiAlYvrQ5mtFxtJXaXvJsl4nfDUbQtnYVwe2GKDFY
NTUUrPaTZw898e2JFWS1RWHo6/Hm1i3M7PVNxmowSuZ0AC/XM7Qz8JHPPDxGWPtSfCrVjmUmJI1o
arUBCOipYrJFGUelmuIkdSB4ZKOVYlv909ATxJcWs05unZ2pHdeZOo94p51s1Lct/kgqwF3AXN9H
2nUUkzPUan2fRqNytWm9LE3W5VTgIsKP+PJjFcuqhjm327SRNCn46Ni2Ry6OIG4bPi/VEE9X+xZM
ddFdBf9xclpilz4V6CmISmg1SUQEoNRu+As5u8AOOuTS/LCH7rkwrAOE5oSIFUTk3WBBmqpGfyCx
oB+P+A8rLMnGazk3A7MDdZ6mXAkzlOZd+u7FnlAOWx7pVfqqmTd2JrlTW6rJ2Ds1ZQQgEGt1RKuw
itZ3IHwJuLaUfjsLCAaWNslsIKbcpfRXKPenkX5qhODch8WPNxOdCoxhQ6AaJWVgn3GhbnXjrSoi
6GsBL3RffJKdPm4m03LJIWtQ5WM4gzm42suFx8ONbZamU6cd1czDnGlyTBJbeEiZtnivSR99tlsE
LewHyRQY29XB6ifJeFrXfwwLB77t7GA+yl1eVtswE0xZa4vufU2BF4PfkNai6JlCFhZJ4a2Fd63E
lyXLuEGUdoIJzk/R+3NfCCuO157ckJkPT4++ZSEcK31+43jp0+ATFIeOJPHJiEAuUDlu1SE8W/JT
+65JUV+4K4dMnzaCH6TC/mjxxbT+yHok82EU1wM87K6RhbP0AoNK2lBYp4APNr97HUuG7AH6xMIA
rTpbh4nV+9q9gO4j+wKlWJYWYh/sWDJxHKsSGeKAUF9uQqJQZrxfdcdYUMMm/9RJe6wtQ/TCvaeB
+eboBINa7xq712zERf+6JPx5UzL0mDFL/cvzgvvkQhRcaH8pHsbgyR7jgyyKk31PPhdFi3h+HwfQ
CNOmnKsica4YevKXg3pgwL/+Ywwb3SAmKjApG+Vf6Yz++d3HfHjsDyxC+FMk55G+mqbUE7mg9gbP
EzwO01fKrNLlMfDKl7VwT0oJiKkjt9AjOeQOWoY873LCtiXCrQwZ8Wua9j+7/OPbI1mCj+QgkDfN
z6Mtlpp9g/kIXiB2gBuZRt0ZY00ogkbF7zyqcB0yGbjt+JHnRPVzh6Zz4HC0WyC615imNq55H++l
8rPFQmP0Hh+U/L9Or6SUoeZL7n34SAN6fjFFmu9EoenLZSSNMi41QlboPak3t42Rktoao89aa5i0
LSvCf+50mN8oOqHUHW9ZoRI2L7bg2vzNbH2aeYX661zJxQ5fDTx98lXEAEZo8j6VnZ7w4ArbY28d
z7e+AiZaFyRo6GnNTfAFdX36Is9H2y5yOBTZ5c8nVgotfZ//ZHNe8kt9mQ+1TVxbuxYx9XAO7QsN
IgdooDW0HvtGKGuj32EZ8nsumosfHqWxKj83qDuunGZeVQ7q1oqTMdnlnUXe8GjRNHBr0fxWFOI2
EUhosGDupDAKkHknhuvK3KYH09H8TemNyvo0toUzUYEW/tL7KlT/DhxWwb+9yXNVjFbiva+7zBcp
Cjx2knccGrxZoyVh2V/OmvOL5ZOhvtNLvlAjbunsqw6eL3darzHiBR9BNxxGDTEsAKq94l7TvmAR
i5DDDU2CfNpNpMD1EYbTx6lzRAd/svuon3aYCRRx0x1lQsjWBOxD9XlQu+t8vFJqgIo6EqzUevhg
cQlVwkLNhr6sOcrXeaC/ecCYI+CekO+WOjU8b98HGbBiRMEr5p/74EAKITgijAPoTOGecplXKxBj
mSe5yWfjssnRcyp8bG6oqgFS9eQctOXsMFU0BZvW9sVZSfVpSE8zqjrtqtGAygOA0f8lXYN3Vf1D
p9q19oV9Fvo1gAmxQ8/SQgUFdWImfZOGxsNZxfF3X8UTSWnmXlBnXBaHVVtL5SJZSUL6jAMG3zJE
ag0g1B02PtFF/RB+Ed8zC0fFnRYzpRbNgVhFfACpmWGmODy3D3dLuybfWWiTuQuxkM6cT+SAGuSQ
9dWIKDMYOpkB2n/iWsyVjmNzdYINHeOigFOLt0j2gUw/MjjxvoBYbnBf9SJvX86dfH2imChKChGI
fIyxBl2HDGdbViEKTyuX6GHSl89ydDKBy7aXr9owbTT8xxZqWjBYQPSBfFhmK92fzdKFpUCmg670
4E83f+nTXiZO0c34QSPvScUN9jtYxRjmWoUHx2rR8RuidURlFh6tRSdU5Vk9SDVDPasvJaBAP4VX
d959WhJT9QLy8Of7FF0RzkAb2OaBysn6sdUvoG5aMma0w9spKrReErrimJQf/9edMxheVLJKLaNs
973Tf1FnhEv+z5E+mk9EAQarvfBcuF35Xh7JKxgiRv4yx4HHCi2s8Qi7AzPI4+Rvds5YHC9AfhRS
8xXa6a50JUIDp5ThX7de2fnpnxCtSIVkgGgrOCcdBYLITq/6H1bS2mD0AsKvyDA9sSYab0G7jKSs
T9nE9JZTkyynQ3LVbGnEGCbPQNwbkMpGN/oFca8rLBf030VxWPfr8EXU77WxWoCPQ75KAMXUKnbp
SrrcN1B2okdfRCygo9WYPld9jKifKBCzq1piXNMNvwHMG1CHp7nchr1LXXcnzWfV1vdIM1Ye2lTe
c8UaOgqdsoHJHyzp1gAJ6MUeL2bUEYW47q+WgyaKEi30oDMcxP5/um0MBe/AnXKHQkSvQYQAmPyu
qv290A6UFnN+YNeB8GHHMSEBmDF1j+GsACw7Sn9ZNuDMfPo4iGhPWMvw2S2oKmq5eOTTJL2r99fZ
XCgXttERovd3uJgHcS3vJB2WZTZch2XYqhsr2+dslgIM31GLxHUXm+UuKTuUFfe9pxYjhGq4vzu5
z6Pr8hIhLRXM1GZQJRS0z0El5Mq6K3O6QikastDfX2+W51R6SE7jzz7BUwH6c5/Jpc6wvJUjXaqQ
QJdxOnL27bKX1Heg8f5LOKZ9ksDdXvqQAH/+kwcwLeSfDRPqYom9cQVoDoDFSvCSPHubpMavEzk5
9lYRs/df5DbsaHP/qJKIzHfkp0vwObgyp08HYTuU0RIE7Xx4shnwHPWl5s2PTTp7FkVaZEdDQiz9
ZDn9j1NL/onkcn/u3ownuRBU9PjRVgWH3qFENHI/w79jHNOMB2oM+W9K3xfOQmC1ceeO7jV5Rssw
VPLtDw/m7k3WXM5IRFi/0qck4bf9EkZ/TZkDAljNVccbGjVGjPjCdYc2x2J3AOmZs5/QAbmB9Xl7
3cj4rZjv/IyVWdz74TZMx+vNYw03mJI+XjminXXaKi8E/lwDQkb6D4k+7zxsxN8XjAfkDuPTZ90f
rPcYHl6s3em6lBi3guFxW9fB59SM9PrNexxQKaCAOPbbeYB4wjXUtUQ8iCJkgtxtqbQUkXjeAGLr
svohqZ773OvzObNHHkABxEWdiQ/jMZJWDM+Ci5x6o5Eo1LVnud6iOaeSyACM66XlfLn4v2l3ONLg
XeF/6q5jqzB+9P6EVg+5fjQ6Oh04cFh3LqyfbpqUqdKX+rXovvpzNzCUCmkN/9bRljsVQDu3i1wT
n9WbjpUtBcB8J+0krsfD0ElVWAqHGvrjpT8MUimv7ipW/V3SKaCG1Y0U2j2Nw2SD9JF24O73QJuZ
2YrZ4vGbMKtKr0VUhd5sSHs7TWR1qY7bgFBTPV/uKGHue1oAf+gCXE1mhC+gIw9BiwVu5M7ovCRB
hBsstbJm2ze0ckvVzOoLV8nj5fRnds3K7RyVvVW9JlHN5PzWH0nVbkHf9fuCZL/o3ZX5MaGaWfl9
vA5B4gxsTRoXHxftCagQPnWqt4LSbsiRe2+BnpEv+PLhwKjgaiOeyUNHun0RiW/lIc1McqkCn4ik
f+x/IiWpT3BxVZhdR3xIyHniVntOvSyC7d8thy0y+xYOhqpJhFIqs4+eOd9zZfbNfC9umiaXFJxa
bHv6VL15jOuQbB3D73rnyrHSrx7i1wpU15BGLEHhXCda12A7OggacOLJWneljiq6gOVh3WQeCU9r
9GYNSEpvltj59ZJV4OXu6IE87cREKNHu7z2KiyCroWDcjW3Wluw7baKaygVEj7xJz5nldaS/epHx
daeXyhreQlti89WFKkgdm6QmqPUb1ueqOM958yXN/GfKEUKA8WLYEXvHrusIcBTgll+kDxdS+8UR
zEj8EAwRPJpjIQYiEp8dMWjOyVO+SpoHkpW7sDf9R0GRnaqVsIxHPjkA3KwN6fO1e92IKQItIyUW
j0l9DHJXG6v3PLH5WyJsWGUaX8iqVQpIkqQfLQvqJbieqP96Fb10/DGpgwyOg112zybAouoCiN1J
ulYLAGoogv0ikp5l+Nqaxg6bn7p0y8G1aJbyxOKL6vEti1x6jvdmoShqIT2Vi4LS21yekpbmsV71
uTtHc3mA1BXfYpfbFD+11P5A9QexidN0DmjH+XXUAdrWKA9MEjPdaKsSohIJ8n1GoWcHEDLpxlZh
8jc4U7E4MXHCtP8DvpY2jZcjl/6WgElgZcydJJ9c6mjaQfngwT3rFeNGTBcEKCt/o/vb5SImXqwN
J6TLD3h/iCHZ9maDcaYQD9VW6ZnrqJ/if14L11DpaZEMwa8y9Idsa6J/X3R1Kr2XxjvhxMKty6yd
iJYyN2WNnM+IwUq1LRnKSGt1oIWOsLzYC2eMOjjamzH/73LmCfqJ8G0Cx8SnCV9J7O1bYF+hajFs
0MJbWlat9xP4efwoU813dnOLP9ULqyWIaF9WfUl+6eKp6KdF2d0ZN0e1P6ha7XBl8m9w9rKW59uT
h1Eg98pWk8HmDud76INkCQ3cVmVdlDvC1jouRX0xyu1vgoUgJkMaaapCqi5StLdFRcXl7Zu9yLbL
3ABNPcfimV2shuGYC2zeiXC06d+xUuC+JUqnTbM8XWm0ib7RqENXYiztgAWPLAdzNcDPKHXO/T1P
iQskMpDOM5czmNXlH/M+mW0ncbyWZAB3JasHcxYFWsOKk3YTGjQ/ZBGRoh/0rRy5Fbng2UtO7ct1
PogpeR/vIRyLvp5oT/eTeeD/WilkMi3BnQ1GyHP+ezp4/QHULBRu4p/MzFJEuGQTKgEGHnUCv557
lWzcTWxfIzBCN6QnP8BOOwpOh3WiFGr+SO94qXA5x2i6PudigcOl6arlbXPotjlWt9MxIk93L1GR
uXJlE2/QiLv0huk5PUcTv4wqmIIcTdyR3fkr/+0pFubHcWttZdGb5VvQDyK6vfNBG9VNsPlwo0Oo
W6xZQRmOkE0KdpQpd4cxA4wpqnYdgoHfppo/FsOSIafLoYrtfKwo/VMu+6MKBHQUJVCjFLgKajLc
M0nfwq4bRaUYq3hDrMTZR7mCeuuzlhLHqzzUWd7XHaZ0ycvIMANZoSLwVt56r262A6/h/qS6bfD4
7gODDvJzNh05ba0yb5Y/0CNPgWzWU/TO5aRWAf0i1QR+2Gy14cBVk7rOMlJF9pcu9YUf+7mq+LgO
zC/n0rcHhLskQDLYcbPu+l0UPl3KE/zLvQT0uOJ7NHukCDBlZUAn9ZVgAAXFxOJxt37XBI74OiYw
lCZ2F+gzt2ANfHPSpbXbFBHZKoVo73oh5Nw210ddRZBeuKQNzUxJ7ENEABt0cqBow4lBcDYFgXKp
gLst/6uCGd5HiK5cbXb09uqbJ1b7MO3fNkV/REItCNHf+L0tm1MtZCNroL9o/xU5Aaf7/X551Z76
RiDPBgfJjpvneqGPtcruEWNV4q24j2NaTghQC8FA935H7FpVsgYyBxu2qEOVeAXw1xMJP/vLBZ8P
WAtoY+JbEcMjlKnolSxXd4gCY1OOTPYTQYv9AwxEX1PBleNgBQ3gyrkIsZnIyWnqlDstBa3/YRAu
1CnBhX9hVDRjO8UrQ1CWm9AVQzNu8EcEj+dZarZ2gGQdBDQ24dHibGCvFpigtr7Qblfp4aeRQwAt
A9nLGrdXiOlDWugR23H0FLZ2B1g40cPkWcv56bQw5oZL6toKWtylWw17Et8iCwCShG39QMIUdss9
twEss1hLFWvWk+nOvvH9CaevnHwBL07Jg/Kit/VHKLnVkbS/J1BLNNVPnkeK/PArV9xlZyXzrrTg
3Sp3esYuoWeY16MIGylKOgwUoxQUXm1RAKhJ3nDUVlN6qG8rVL7ENlAS9ke1HdOQO1K1/DTS/wvz
cPMtZUHDRr/sPvX2CrzxKmGubeaVv01WiSOUbLrsSyy+lcbWBOLEqufHqarHfBnAWlgMvBAMFgBc
qz0CPsEm72iLSkVDj8r4xzGTROD1tSOuDmBS4m6av2ubLUXInL3NCPQ0EH1dTLlwUfqjxsGyrIT6
M5/9p/AE6PbcFLDwmMYy3Wc7JRLsTNK+gYbgE7Xo2G1I5+zvyZ0y82E2G0kELPp0FiTn4gnDOJKr
NNfT78k46e7MFOTVWK+zMdKb11b/lhb+Un3ce0bLv1eDt4pXKhB863j1zqhlNETqH8gU+87fMeli
8rK0ihyFKDtKgepcgMw3K8SIUpy7PDufNcvHy7gdSgDwx1vpRNCF97l2AuVYOracc6AAjEFhzhVT
tbb+XYASUTWYKncHBzEHFy0TqbkxiEVvuqXA0kiTip2OGTBFElfhHARucKB2qx76V6eWtNO3oFwM
AI+zf3ibVCFYF8Re5cW0HZuqdbho9TNPE4pJYNz7DVlSp+BQpv6pY8IMMllUxpIs+4F0pN67R13U
v5R4/KQxrDHEA+SmrSg7ieJYshaMYmI9FwmUJRW2M7XY5gY2g76TEr7LtXMwiyhWjhIORtIZY+QW
viVEX50QsQEgMT7lb9xSfjp14L0BVvySfUmsyZA9LyfEqfC/3ZWi0Iq6NQXG4u5BSKC/yckvC6eK
8+bdsuYP2Ec8YCe6WY5Q+N5FF82VySSGPHCRZW6aMUbkfo+VwD63xSHDBLKFc1XMpyVipahB4DUk
UdlGZcHcABBqqfb1yx22ObHq6Ab5+c0jicfXLivyXZOW7hY0GolAQm7fvyxkayrWYdo3EmndvM0W
a5CTSz0JPLh/dWkpUHNK/AQ7OrnhZOuOrpZ5qv0yG0XO6z8CrBDdX0UkvRYyI8ExkN++4wuCn4CM
46GmTVQMeUsKgVS9EWaBVTffb7X9Bdmu1GkpJgvZhS4NGnen58EIF2/txteihLfGfg1eKPO15aRi
9DWppFQLIXCTVo0Xb1CMVm8aHhyl5MIQivU9lVr+8FH/RG07Y72DXNtW+2Qmgh9swD2y8gTcOXfc
eIL40DvQHHAEUXRB1zoualxxY/cLd8Gdwq5p1twQJS2rK8EfN7RsKPgmZcuVsflSsCpwiRdehCfF
ySLfBxB2Tev15Z1+BvHpYB1rx3mphFrJdLBo8I3y8eHHmL07vWeXkLxYSHMcVHFyQz/eWQtP1C7O
0qPmJ9f6ugFGFVYoZreoET3nd1VV5pMdRNW9w8YrXSeCkl4PA1JGN0Wdz5GWVDkdm8rUAaMnUkPY
5VXkBNHxi1+7/bZ0FYqOQbCrjq5ZWfM1AcM9immZZ4hEi47xvrF6Bkyknaj/D2puUVMa0AaYXbcQ
ZOKYmLvUE76QMq54sL0kPxjUoL8rIYgnGSJcQxDLCRDQn87NiQSW+ceKEHS5CtvVNzp3sltZwPLI
mq9T8aNNo9u6wbZ7D9o8pFrHI0Dwrx8c+MRk5y2SRdGad/AR93AUbqv74Q85xIb0cNb0voC1zgGI
Yi1DjNfl7zuQqXtfRMimQFoyxzDowmefHaO39bjtR/ubBxJcy1WvryURR37dE4fLaAQFYT1Oirud
qOBVJmIjNc2mMUlC612z3YzKLa/PyhuarH6GKn1l0YIuL/MSa6Tabmc8gWakE/FDAhoR4kjTtR9t
DQbgPedFQO36wS+2oIvXt3HXLdGsQaiDw6rX5G0mbICiZm4SehOyrbY2w9t+GsorsJohpT5Y6f7Z
ccutU2qSN32CWDh37tqj8zQIEwQtUWMpT04m9R9rMwvD6RVAgfI5H14o7zrW/inlZ16diKUBYJ6f
YFo2rb4myM3tZQ3ZJIJR6YWaELJnpN2VitQJvWo6zZPMTZdFOWm5kfSopoNt2Ijsl8WNRz5iX81x
6Fkg9idHKrnUV0Fal1ffTDzaYzkKR4avZNbt5YRxXAhCFbeskhfbKHJRrTmBk3BaZ5i26CGJNsd3
8xI1mjF2qiwY8+J4ASZfR2trFEmH/pKoOl8u1QqRAxFEHYh19RhtagekOUQWv5elSeGdjNshGmzT
e0mARKK1YbdR9LwYKuSZGDNpwK/zNKlN0VsUrn9a3tYWoVgEwXouUb1SJYEn3CKrxhZeT81EFoYP
7BLBEfxPV6dg8gu3qckeJYsbbMfOzqa4leiucZ3y5KiuOkmoT5sKGXqp6hnNUe1Dkt7W6hsoEoIt
g6quPeKil+MoDqwhaB8jt0doxkYsIwYyEICduWAbnKZBFF8628BnlkJR9Uu1Ng9syZNc2RidkeTX
Qw3wWkI4QQJgWtxeqbyHTTaXGNUnZNDOzZu4uvk0Yh4/8oSODweYCUZXudZru0bbGpN/0g4W/bdJ
VTzre+qtU1Sy3nPg8wwsapRA5knR67QNWhw3RdZ3COEq8XZ5J63vkm1Jewu3GSchyn2KkkKkm7z6
1jP0BrmQa0D12V8E8rjIik9cPR515zi/AjNW8OILVWJJ6r514G4fh83/+0inTwxfCfCVkVwFVM6R
vqjq8h25uxu7q+m4PX5+P6gQr7GMSeYXoWu6s8VlyUuAO5tGeRN4lGFFCGGYJYRCK2+h0zEVg8CN
KCMVaiX7esm1vH6hwN8MNxDz/PwM9YuV2NhQTwNJiqLX29ZAlK7Zx9GuNwr6D3UiXygy3PcevArQ
KjHsG6c+MZCe5PKuSi6jKInzSsYP0ASPwGLzpyUz68j2h8XpX6+oTWLlNIUcEnrIr9c9rHsrQ12u
QAI/YBygpgm+BH4osrdbb1wuWOg7X/wvffEtyFk/61BLcvJe9dep2xrUo0O2/5xjN7GOaI8kMMHe
FmMWdPZS0BjDj8d4Ia4zkNLOaZACfFMxNII/2bZmWWxoyjCB+zLpOy3FSaLLWqMryy7G1+Ed3zru
22OfhnU+b6M7qJGJOZhsMHS/z14+eXX8oSpuohJ+/dNIrBhJQCe4i2TvxnJ3Ca70YMkYzUjTdE35
EuP20jUndEFuPhlWSrIicbe+C5qc6ef98OKyjWnfQN+ZzYTPndCUFw9jYWS3MI+RL2fz6BEJceFu
kzcYut+ArSzaqVAmxBfJP5A74wlgi4OGAkMm51bsImZC9s3GWw4JE2sqLwZv6pg7GF8KrSSl/43o
eLb9ZE5xyr87jDQquOZ1WQW1T3U1GXuGPLp4zUP8LY78gz7R59ylnNJPv6TGxjgmBA7z9Vh0IQr8
MZEVlGomqLVqW2ORYUnD/cI5PBqEiPDZB9eNkZmmu53Fzgt7Vk4INrGcaQ4rpgZv3ujn48/jIu/n
OLeBKoV8thUE6za2XZSxUUsH/YgmMLnKoEY3Ksp93tV9yO0aRgjA+46EwHjb5eKRdDgr8dtoQ7fH
kcfLvMTIrtWgEclw3x4FvfwlGnEqIxivtqBkDO5Tjt9JaTxIE2+FnW//heg3Txj8vTRdRIwme6T8
IPfmVEn2zdIV4sxLWmr3IgG2wJHoYRM2qgqx31d4OUae3JGAiWSnGhRPqg8RgPft0S31bv6k7CbP
qYxFCdZJQ0ge75s/KCh3yEXbXM6Rcaolp13MJN8yQtwA03k6rdOGV3QpeOM4p1YWz1eZznWZB9Sy
vCVDsadEgP/Vrsywb9JT05Y+nK2kEHrGPIOoOwGpbOf35Pmf+T23LSjvAm9V2bo7hdQQZO2lZeKB
VehdHKjs+Eqacmk+jRnVBSdxyv7Jm+PUjEBA+WNYkjwczDsotsspxu+WEE/+fz7bv9r40h1ngsvD
Y67rnlfyTScPvjz9cgASgXp8lNBwSh5N6+m9d3+W1k1m6QSCHW2Ujql+40UoYf0dOliRZGBJeFLO
mX4GXBu4Dx9S/CY6lZgETz3J2LbpSlhl2ecAPiiJkWfo6tUJFEHr4SnKWMlQyKFqnfJtcES7y6V6
w/7qGdVSvSMiGt8MF2XWNlf2crrrO/JBwbdcxNf7QRO1Rm0/hEcz4gmPVjG6h1UDM5EAxtjGzwPu
pXupqNg+llgUmCgFrZlj6KOyCSZ5OIbCqx55k/RlLsAzHsq+XL3mEW+ttY3ApSYisy8ZPJEpGKJ4
OeKu6whqNDKugSUVCuVYyoUDN63Za8shyFX7Kfev+UFBr5rk+fyYlKSmq9GXvxZ6/tiviacSiM+b
aJmRNOUQcDZvwendDO6Oo6Aj8Ag9GOkLHEuck5EA/Ra3UmLEN2fQuUuXoyPzcZYgmlAKiVKXaXvX
RjShQwFGgeA+AUaRdFU4+bRV7peK7Ak4DSKvTqvlK9oo9Au4NgLtLbQPnd1Y0eU/NS6Jg37kaLVV
I5KVbIResrukFtjCbYJLWgzUCzF5SV5+Mvdsmh7iIHqHbJY9UaN3jSVNZjf+wa43Jf5sYJMm/xsE
exdcFaimQMInJKb7NnqrLqKiq1kka2h/XatdKmKr1XdyZ4OvUVN9m+Zyo2kG9PETsJwDB3vToYrT
aPMDENVJ2G/T4xV53zmBP7Gy4Evz1dQ45o5mrWv2OnISZyIaqLXSehxXYstNYdARuGsPvw074D+s
9TXe59ELnLqbFCdJTgq1w/iWWRKoKTKjBY5Cbo981Pb7/4ug2z9GPiFyyWU2iiCxbaus8TIC1QtA
MZ2VtcNT/r51gKQk3+eYC7W1sfcn/HcRBdw4XF9ALJObiIEe4/D1Ly4tQuoOo5i11nWahh/lz71D
Z5fQSwEL3i29mJoa6pzzcNCC25hmOYxHCZXJo9Xpj0WIc2DL1ti8yqab1/O3nSZP3cot0miv3Bzq
gMvuNKAqAnT8wCpm7lT9Rr/q2i9nmH7iuPMPte7wxieIglKF0b3a3jOfvBJT/B3Go0MMO6wBVs9J
9FEItIey4xZuN9TvkcVOpyUXQCqWmGqDFD4zXq9Si8rn9RMOBy/Bjy2gEJ+ripgLoknbZCsOAAX0
sVKcJXjxVrLwy47pmbxqm5h00LNB5Z8sXOXlcpK4UI0/6SM0DCO1WN2yOmkbL6g68Q4IscpL4HSS
olR1rifHFv5ocViTl7EDa9G2aTA8hnjd0jhj3hbxUBAGum1l3N6P3nhk1xJuAF/eG7BtX5syipCS
Ir5vY12VV9IGfVhVk6CxxPs8GjRuREHT+PaomDkxxgFI/60dCatk/9nBCBps7AraIqiYe9RI8aP9
SxVhzrXQewRYn8EOh8EXeezcOS77fyQSzfBuSxiWywF5AWidslu0aMurpI7kpq9eRqnMf5dTw4xa
fw0pKKtB8/9FQk0ZsFwZ56REYFcTiXm2xIZUCk6YsyGi2WxY7GQ2k3MVbZI4g7z1uu3lx23WjKe1
grx3j5ecTcD74LGfV1MF46NDly/wXKvHiroSQGdy5KVvKCpKKBfqq0KWzvdna/fSB43kJNfSsMjw
599HTLR5LNNXNQkT4PrUS+aJ/g+ohVkJTBRvHlFJWL7DHJ2j3G11/TURF5zz/ikdSxDtKrERcvUy
QfJSoL3WZ1Yg8Ljgnd7xSlGQllDUdWXx0wNQisnRMI18Oun0pPqOOfOW2YONKQA5G/868jK+0Br8
vyeCXDiP3wAEcusg6uQG/zzliWkifRr3x7pAkx0xj53swbTpTAQ998AdIZcpdVWY1EqU40thZcNe
fe0D+vsiPTxVLKhJjezcD66QoUSqA1ti3lA6FJXCuB3SA4NbKPbPyu+D2ESi5iXXGs+0v3lFI3Gl
k21sUybSYqkCG1GqlfP/QLVqOSzeKpWIEY7hAOdyt7yGZm3PgQsVkyp+qaLA0fp3RITTSAK0BYDV
pRmusJl88D/HNzRgs/pS8fe7XexDgj5hPDV0VM+CVRD5xjAkq2BWbTvcbhXT+lrBwZLQhqefsk38
ZL6d7/NM9H1p7LuOfKOqbw1+yBgBGRkdKGpECXqIbB2LI4Z7tT4v2cc01uj5zopa8AY2oheXEGSS
LRT9wogLyuSABpZv0xnPOeqi835XVlr+zuQKJbCZhRtNp+d2Jw5hamdIrZo0mVGdcFsIC2mWCkJN
GSZ/Hj4J8G0pDZhAEhEJRNPgSl7N3XDF4pe81gCwBrnec8W0SEBNIO+XhfG5vyiEfKoN9s9REmBF
vpP7XsqKaitMrC0aXvH8rwjKkDavkc8qk2ziRImpvSpUccHjRUhEcgPvBUr5rsU8e69BQAEbCssE
zhIjObx+pRoPiQlbRiohnkXqOcR6ByaR8PAsr3Do1/mbcEFO7u+gMiTDF9n2dzrsiHYIIurTA1FR
jUkfZLRa6dd//HemC52JLt3cXMClUYT41QH+TsVte1O+UD4HjQWMKZVzGyfAS1GyoSBQ/OwfyZTQ
QfzPlUxsOh/IX46iOYPGg7HoWXXjpcWqXwAuGivnIsTjNb8cT1ju++3N9rLE3B6hYGRhxwKvQI2B
ALmSqe8IN9bXIwboCtr7Cjydl4zdrvcVABg7k5+OCcXSJCW54ku4P53T7xkEZgA8d1+Ym2fXJZH2
+CeOdgoQFvN8OTlJdHScsSN2nQ0FVPIKItTGdVBUqo6myPBk/Wm3sx/TmXmY5GiekhLmmIZkp7ZB
mbQO2lqxXFnqSIAB0MZcT+w4OosBmRTuytY3B5Dzr9m/pzjrQcmMfiN4UBCTOWvWKG4QlMkjfgXd
Lsicwq1aDXSB5TftfWXQh3LsfUSfWMPvR4Vrus11sWSRSjlZcN0YOig+pUFFPiSMSMUjcnknxyW2
tELxH9Ne6NjY2UcuW76PoN5+7qup+nQU17JJED+78EYiJre2EIBUTNSIOr8HgY03et0zF16aT1H/
3+leYvK7MUhw0CnyagCbMciHLcg/Xa3XMouNCrZCoa99TLTmQpslQdcCNAbg+Wbb+J6jyqLWHvYH
uKYMo+HJP692dUOcsYYoa1DjAlB1zh9PYSaVRx8qIySShSCpNGsjHBd+SipqLDVoR4bUrGEI/sEE
HXEaL363dw5MCXrHFFZWv9gzzQ6seUEDmtV2Bgkv05tkWUm3RL4LhG7VEE4M8eALbTa1dmvOR4vs
1Kz2LxXjrvGYAOWUoJRLmttfe3NnCmPD4GYjvHzpIH+l8qI72ChcuI5okVqxrog+qN6G2xtuDj0N
yLhJEPhzcrNPbis3jxKwWH7jRmYMSkVmocdfXLJeDuq60uSVFt/Kmeqo9J3UwYyuERZWol4JhamI
eXfciSTe4cR1dSYVbgEAIxaJZs/0dmerqyNJ6D2nbrFR3g4HTpyIup4Qm3qwrTpOf+EZezgyCNLU
tBvHTQyn2iZGpt5Mb/K/kwoBZp9Mk8q3RHrtq1jfqKXfNG9rBPp/e79vo/4sGu2q5VzCREGckSvw
cX3bMfwhPQd2NFJUqr3VsZ9ObgbezoxkTxmLw+zAPWLQRQBapHPH7oBQFi9eThB+JfjtvQb4b5iE
PShOCDzrUsNgeeWjO+Oq+gHFnIntJmMEh/2v5v/fs+g0EtVTIscxFp5+oB94tSZIV0qTUvEWuIGJ
MOlzqo1oBdjdgqF0xZcwG0RWt2O7HLvThqNW5Z1HO5owC0nHKD4hbkohfT4CRGYXA3aX+hcIGM/O
OUu89VTEnK1OIMO1dLEgyfXVqlGG6WIaZE5tK7+ojHo8RQD6wzPeUqlB/oEzvN1rOakVBLloDM4d
Ws+22pge+LUHetFlani9p3jQwPdKaDX08aBLBRqwnp06KVEEEy/+tbsiQAuf0fL396hfY1Nkfrt5
lLwg59fAe9geSwk0zN+utLM2pcQ1z9SkjcYxLhmpsMGm3oZ83DjDsVzsB/n0gfJM0dsGgHgBj9hv
AH0hvFbYwpLG6xjZrxOe4I2C57ypfGBSCS8KY8DZaIvWZ1ZJG7Sbp4B9oTcCVOUEGIM4LhKuVKfY
ciz+Ts/HG/6VOg2LRrsLh8n3Frae3t/vZnH+j3Bus4EmIUweMO7PCtKFfmafCO6jUYCy7Q4r3kmH
bmWKhz9fNspENPRZX4cpOOcEbvfl6ysMOlv92CZo9TKndDixEnnw3vY0FkhReSu4oK2dpUUwJhYx
jDFwXS8D5Gt85BgbgAO7b3Z3C79HMN6ZMoL1eY26Ot3z8GzKd7+sI98NrKxNVYzI8z3oqeOtli5M
u3e5VjmxbbCTSQ/+cCbOfugxflD4WAQ1KZ12D3gLfLxQ/jFhAWNqoKAXXf/YOlG33Kdzhip2w8YL
GmzI5p+ErLpFbwxhkgwIFFWwoflDO4BR3oEin1GBNvbozjHkbd0E814TDpmgVy6U8O9PUQmumxB1
9DzNK0Ev+0DdKpvHC+K/yAutNIWsk0Ki2ZmQThd5Yj3D4h4LsdJ5ig7T2ihEqTiW6Bm35jbFVEAa
p836BDqp7ox7Dh0ewzy6qVGwZ24PoLYQQo8x1eytC9D5r0a6hw5SsbCcJOn08hc5wLBYudcPPEiQ
nHG6YjDzvuu8eoispfy+4+pA9H99Ktc9o/qVRbnprMqBEtUu5czHYxEUtYfN2N8WS3LV++JMuOl/
MeMtQsWznn1MAUsw0dK4KnkRW+kF9bll6+r6ub+/rRkbZAUdPqheDkvhr2Z+104dIz85nXC9STz6
Aqq31nMxX+rSE0qfNBa8bCCgJKt+V0mF9ze0Rv70mz11dAUliO7YGpBUoqTPOjqaRf/E+reqBxuW
HHKx41RIL6zJj44rdPdkQLpxwowLhJK8vcGRYldibG+Swg7fPV07Uoqki0s2XC0ow26HtQM7BdqL
7eHSmIGKdXQuWtcCBctLqylVygTykq1UxcADXt9leaD1JthJ54N5e2AWn+ACIxvgekO7MopIBAiM
3LPfho0Zgt2sjppxFOibpq+MI5q7LhAdHHDmwyfO+WkGT7YLhM+O+MLD1inABFST4qocEe1Uzv/+
sKQGdwn2ee7H0KHmSAg5xzbR9ihjt/b4bpK5q8wMamJEK0R6CBRwk8DOkHWPU5UXXiIdjO2+XEOa
mCcyqL4CvOuZTnBF7DhOFMDSRMRidVIf5MlF0ofsdf1azs5A+S1ysMRgFSKyApsS2TdEgbXppfcJ
KZbnxBpVhDbbLNQiE8O9f2kAldpobr42xazVfUND8+FDLzWTBx+IlbjiET9pEfFeYP/TZwM7rPZ2
7MUI7O8s6Dlynq99esct77U6xtb6sC4vZSjuREVp7FkYKsH91ngr1LQtP493y2IDqTaFoBRDZVma
rwsfha4Y/ws/NdSqmuBI9Vl3mgobkT0IkF8LeM5LtaY6kYGRg8xpimKrBwPt5xoa80H/BHpkn6X8
6HZwhCS9Tz8PB++8XEBRiCrj1j3adAysBcWGfugZ0F4Uyb+C2/MIEaAG9WU6XI6w189ZABszMAu5
qWkPQh2qHjuSnX/3DIXRdMN+yhzamzJwquZYnwC24M+4lIAXQF+LeqqWUJrTjeWoUet/thR7+1GW
hG6t6r7XyGCmogGb5nZbJMz4wF0BMG7FyB4fhVk9iidM3rG1bhZzZwna+rQL88BnMIvhQL2/UYgs
vFDuVnuUJRZYE2XYynohfWYxLwwa1nUke5Ng+Ev1cRe+B4Rajb+mb+UCXnon/RVP/yZHb+3JVByW
H7LfCN+V3VBFXkQPxWx2cILwm/nWn/UVRGFnFxlNuJsDYdY6C1La++zUQmZlCUwZffbSPQUvD4pz
Go9/aNMDDROzyQdgkVOCZFjmlnTHXXATky29P3Tp7ynGUGGN0GX7liUZzKZWKb+DXkVhvfVFIHXH
a3AIAHRtq0p/LoySyj7oisyNOWXLMw70e/wu/wftqeTkY1BOv9EB4eNTU6/3puI1oEMoSlGN7IIg
ijtciLCqyqVHxi1ERoV1A5gxATurLvxfthXYrC4X+IEMAmjcybq3lYlrj8Yzj26AURrJxMLiFRLT
PMXqEcxUzwwzYYPrF1dZR6Sneeje+Mh11nrC9V9kWlaVSuZaNQbJYSEqn3Y5GhGWKgtMtoDK0RWP
H509Gq7HqfZqXnpa8LOFMExiZdeogJN8sFEGSXA/6wNepa8w1VaODTPCpUxgPyToh2jRqUKlM3v8
7d5rPiJ2hyUje4KzkkcSJLO/zZfuRlZeEDe7MFGBfyunLF/eyKj6t4XvTb0CjWNniPEDDctQmKYe
ylHezvjF75gTnsd3e403B7nd5ts42TjmG5ggm6Y9QcpmuDbbmjT+xRbGVFJuKn5biLSD68jUWDoz
KaNFp7qHpYWdrVPryNm8lmwe8A+3bcybA6VRYs3edCbJY8VVRhnfIY2YUa2xv+WzkpTL/hDcN5zP
8+K3sjGv1qs+aypxLBeegdMtXOr6mEDL578dYR09Cc1KXOvz7+U8CIJHSLXULtxESdO5QhmPgA89
OON542fxlMXbsNzdOu8ZzDXg19ABegbJuS2bsrLs/VXA3zzsrnL1rh2vcUAg54n5HgnJOnmRSan0
mMplDvfC84qyyxe62J675W5HM2OaoFT71GmhyP2+mOhyaTeSTO9j3iOxuOhy/SNNupkd0AZ0Z/dc
esayan/Whec7FW0ppmH2deC3TEG4f+AAXzOWXnyfr0owe3CBpD2uyqkLSlfLToxM4ZgoKAVu/zW1
b8pbwvsZ8qWEB+nCk3FTfWRKATYGKBrhK6hw5A6e5/evgcI0VRAsBP/6/ECAzglyG8Fx1FioQ2do
ZuWdX4Xo9sq/DLVqXv+hUrVYoQJ0Svo0rq72wRfCMQfWgoGuyHweOpGlrPfXhvZwCWx9BSIxnQse
pLHJNtf7b19XRV1wiSqIucURHECVmqwc8TRZxBgQhYCT9l/1IYDe884WBHugLsuZSP0ChJNk/BIn
aHIbLRl2oJ2o/GB9FVCyp7rS8Ogy6Qc6LKThfW84QIyFRv68zd/NMn7YOTniX9gRMlrPuwnrzngm
DZuP99JjxvH8ddCQi6m5fzUXoBb1P2+/YE6zJXHW5Eb69DEdNaMHNvZJxo9EPQg5IzbcHApukQV2
Ft7S/0TTauaRva2u9h7KzgaEUUtEwhyKWj7CoE5OmX6Sc8ykSsRnakhAUMYFaDVm0utnNKy4gnR7
oD4Oi15IuVuIYd6csqW6g7AMgFJ9Nuf6McKLIveiZ3H07E8oNboj1SNFsNVeZXZQn8v8xFyVysno
kNElywAzBUgjGk7gdtgkF2BYVD1ScKUt1tPeWO1UYxFMmdgsclYrNSf31Rr9bqNAbAeGgyat6l2G
hwzE+YuTmrb6Dg2NV3SWlcBdkw8LPGrcVgMdOZq61k1n+mYXK52JGDrsHMnjmwF20mc8kMtrTkox
/KkNG/vC4y5JDWZBaGkDLpegP8CNmvh13xF9yBmo4nLM0djoejrzlIvbsxt6+Tjan3bx/An0NL2S
mjTyZJheUVBDWh0YnBBYElUU3T1IBnmh1dnzkOM6EhYLhrKI4gYWSXDsXdUBND1/jyFmV9+sCC9x
ruzbmDccreHUuS2GmbLllS+Q8hET4Xj6d+BXlaYEE0kJLfllBye4nVV5DFV3dovBFB4pQNTDBGsz
jc38hht5M1rVKL3/zT1yNEwNSiiKVAonsclAuTWbw8zJH8zMHx4mzC//mLAnb8DzHhUH6H2Q8VmH
gBiioM65FeXkM7yby3ul3sOdMvQZFIFfNMlh0SaE0G87ktAqhKxTjLsR8G+Kn8NSCWTk9rSaqqPr
jVqh6NxCH8GfY8Eb+VBbRj1LBKk6eqeueJIlukkItnTelxF5u0FXafgFfnfbkiox67rMYrq4kwx9
cz/g6bk/s5ZztB3XoXKyimPNOKRbve7mfGMdieKDY1pfwxywxWeiq+P7Yc5tfVbOI9PzRbBNOZVY
wqwlesf7szN8lW3qPNyr/SN5FdrehrB1hbKV1qvsWv6bzjG/tH4SDZWje99vKPXxsp6yHgXFF6AQ
qhizE8vJEEGBNsAPVzE9rcjYeT+ujpzkl/0FLYQ7iL1yA3TwBY85hIAyQrPoV2Za75A8a8HbOqON
UO9tZbOiGzvBFDKfSyFHZRj9PCJTRRd06rFzZnON8CxQTFOGencK2GnwArBVxvuTeA+SuPkTriYd
bwqPdXKu14GN4DBZNSsUfRREs2n0czGpFc0ddMfUBmBA2OoM24r+qVIzo/Zw7J53owwN70yWkVRN
7cl7N2dK1JFPvs2f2b8qDWktS6SpbfoKDmKtiwehyawnjmSZJtHbqwFqfcVxEA0v7ybrgKs5jsU8
JJmIo7K7lYFweiZzrGZO/jPZEUVGEP1nDD1QYR8bGZAVZSNU9Ec8iJ4/SWFPIrP8CrU9boQOoWaR
JT6UBIrPpfgvmr8rj/d8JcTpym1NIXMYcNHYgZtBiTZ8q3aQR17NXtDGHZjoN8Dzx2T8+H97aS6u
3y8+VQxRHI+xzWbcPwYTjkT31G5A1IpeqVJINttEXm8ffUMdO2qxp/pucG0dZYChBCOTD5SomPSy
JaA+glYemnGx+WRvmvCkypHZ9RAyfJNSdOf8/pTkRdIn9x05Zxu53XsTtj3asIWQlUIVREEqiaV3
IkYs3+OrSuYDN8K5pSl1VVI7rCrETRC/LVl25N7yB/EjEw2p1k0z2ytILzfJMn89YmBoKOMvdTi7
KJp0ac/+NXECBOLlpjQxZP0KOS0uPuUtcLqI1uaMsow7jeXfHnACKL+up8tRfzA20JdBsvOk9ipl
L2kRe+iQ/DTvgBc15Ov4q85QeMU8cJ24oa3RhVmpBhYfQCtjPYkueZZu1cxvtAMPpKKIXhikK2e2
e9EeKng1hC6KDBHUaARYkmGRmqWlixD0Sk8NYRUNCHqix9gcG4cNnbjgDapkyyj/gzt1aE3Unkty
7U9n4gAbQ8bFaJ3ZaC2GcIzfy8OR8fiiBKCMOlR30wsaiqQtaqFA+NLU8MD49y82qhYfydGwp4j+
7KZrl0ZPqdKCE9Pq89/JLbvVCD4SXLAPqJmsA31vVdoU3EhFbu3SzYMGj17TZKA9aXWfkWnwZRLz
cApRdNFIoxSL+rYFENNo04lRiY+1TRdUmjho/7Z3WyBO9ub/RKHRYQaVd4yKgDJgd8Te9lDUXAFJ
PxQA64OW7DY55qrRlFw8HL0/bZb5Xnt2aakEXExU40R6lZ77VzZm1Kdr3XV2g7Zm4cO3F6GCQO0R
FkC+iKi1WluboZB6CuKm1bK9VO9gkjXDDGyg8X2AmANzMlng74zLsnEo8D6qFN8hszTUlLlKZ0ig
7FObe5Fogs2CNwo4Z72u8eKYcBtH2UhJcf9VZ67b1xWglW2kLJn7Sov1iQc1uC8yyQKletQhNc+t
9hpyo64Zxpx6/vrWzlvT64+LAQbqFGTMOIgZb1s/mX/MQATwd5HA7oOKEE4NQK+WFebQp+8C4w+9
+gRmqhIZcaTnVe8Mc8R8pfY2kbGjADqaztnQxSo0K1C602CWAakoX6sfTu3760UN1z3Xmm57Z48R
Wxgazsvfq4sUlHYw3RKo3jSpdSX0A1762Qi/iuWAj0pTM3oNXe25rV5yGVRoi1SAdYiWOyAJRue2
jKYMrObMU7Z8llpxBYFLa/9yic2uE296iEoaM5uKVWyTzoBr0q6LM9OUCysOrlizaNAgC3lWOMMo
jBfKhpZtrowPBMgsG3o79CDc8J6/D5M2l9eBg8xpB2B7U/lPIfSYwyN2cZK7t0pImMNzjr/AnLNz
22KdyCX8fjMfeqV0AdhRQ51l7byTcWN8RHX4pzbLw92mBUN/O08THsbeapuD6ra2oAQ+FtTwQz7e
bx6BKrwyGNfzs5eqkAdgBhnH+RiO8smEac1Qh1x4ir538OZdWQahO5t1+xGN1wLjFn+TeGwSKE9W
KU8FHOHYgqBvnVmsB+TWpGhwkE+C17zsETZJTRpOY/hmvk7+L8K6hGgzwW+8pvYA1+gnf9B3UtP5
RZnTR1k0fhCs2dWYdxFFWFmAWqMIEDDQ1QIzkvhaG8oj1UiiLTyJkbKLRjRWtLXV+ajGbmAzD1pr
vx6LhA2O1WniBZ/UXYW9UMVOWKwDewNnQpBVE0q5mM9pJWVpDvZUV/rhkN4Y4C1mDe6mau8xGcyw
MBw/Ncqlg/ga81+T5ydrhSomxX+DUnD7VuC+Lh9zL4Jg1O7geA6GZykcVUbF8uncbazOTheBQ/2o
KiPIoRDLBHgc9moJcwxH8BenouBQhVmSFxHbjW0KqD4GlGuomlZuT9HXndIg/0GqD5nmH90Anjqf
W9Nk/gXCUstljdQZHl59czc7hMoCuA6yrzbclUfb43iRqa2naWYHnIHvXy4JaVxampmHnfQ65Nis
d0PC+Fcw4AgjtGT1gsBQbptZN2tj1tBr4q6TGMcR8Ms8jYyaVdCGzj2ASJQd6sazqRCemqZK6AtR
sUPPiqN0Mx72WU14EOnlMOp3TysKJEDcBNhfDi4HcHydSZKei94b4Pca9BmeH6qemGz2f7LuB2A2
+CKL8a9wE2PyM4KLjusGqSZMwB+1djEwTUxecpbqcw+QEqUJuMPlpL/GemcZtjqOUK9jfOski34R
pXAiDdA0VqOs5DXAT3d8tKSTSGFpJ7s+WHG+oCvnTWxOqSWgdW5uVtevNznzGMv8b5X4GO/JcmRh
C2TkwvuvFMy1Ps4MMiElfCB5Qa3Tz6+OLMZWlLlwRVLHMQHfNs8NoQ6/011mWt+IkslOgXfw9lXg
FP0hcRnOucrsXq0KW/FKs8NX+Gz4Fp7cKFWfA8X5vhHslv6950UEeL4Eg8/7qanfz0QkFHAGYjE5
9Ph4QyB1GxLvac43oIA/2/qIu6UudUlOGFzDeF3iJXrvL68WGFvbqTvl1oPPtFbvoD7dYXSTozq9
ItZA2M/SYg2rrEl5edeuw7wcc8gfLZbxdROPTCpk5sAEqhWF0GSJLEWu7FUord7iwf4q2hKSOkds
Ww3Y1Un6TZKZbc3/2YryNZ9amUeWKWbGxCrvvSVlU4vHFjXKZrr0wzBBd6EHdG9JzAgjxcVUWWV+
7XGPyvFNd1Gsc3iEkYmnzbjnIcfczc+/rGB9xJaXa2keHtlLkYmeyQ52s4aCvKklRseWBjdmyBep
cIeO3cqgcIn4US2bhrJLEpuMdcmDmYlByOv1BOpYb0TBqtuVg37AFRaauB4T3ISmKeAlkPtIq5UU
vLhdxNvFMUs7Eq78VlnW9LvhwZqC3wo/RA7Z8DjoAje/HjRJxJVsm+AvyWva/1ZHj4D42fsTlZB4
3qHR5xpEqwgisqHoTGvj2yZv3eNumaTFS7hadFW+4xoaQvMxQm4QlUZTGW6OqKH5FCjTAZkWBq5D
ICL7WSZVQ44YldALL5tqVs5Vmf4AEZElvNE5BBpWLBj/15bsvgJJmehlKq0OctLKF8hb/v40t9Kl
GOFxU913eA8E+CR0QdrDvNWi2KKqFL/Rqi+pfWe80+S3ICPafjLpVCYtTSqOzmga0P6v6XbSGl77
lSdF1LhH9FhNRM1UYc9I88es1+s4VCR6nXzcDTApXaxSXnOe1WqC+jKKXGcwqO0AAQEYdVEwrdqP
oAHP6OS/hZGX/NZdRuh100CznvgXThDBimP7Qc68kZL5QLF4fl37IqLMkvItiHNSVrnC3P9OIkcQ
vctjTQicwqnvxE1KyMoqJQq6GM+2Neo+AZ/Zoczx5oalrUYe+hmWKWJYLkt+Fkqmb2hKgFeuValh
QXP3dkJetQZ2eGzrIGja8Cr+yd0SQGclGAVdnnElHNw4CcUla2SeyRQT/rHwxQoyfNQArtKzszNo
teOMdsDjbuvzjZM31h88AlpEFgEAb4oOf3Q6YwqSDv4A82AfQbHE6u7NGUU2aHPqTMBgXHzt4N1O
nSnlA50GP+YtfDPWHAQbEGRsybBAI0GV0AhyTWaKo7ihp6cPSQ+CSQUnBHhoIA+0806ZCB+EHzY2
rO+4Efqx/Q1L72q8kNdTKVJmQcUZS2BdlCT2jGWAb/3bNom7aJ84LofK4JqTP0sxDWk1uYMcS/IL
U7ZH8n6YN+7JE3T+YSOm97edHUCGsHkKCbEQyqWwXT2EmMX3BN5iAYvynNvKGmVBVwsrIZXSDIaa
OjjnINSzn8BSXIHhn06Hqw9TCtjxKSevtJt05SrmoA3/mEkTkLFDAoMmuFTG5UY33c/SxIOOybbG
k3QgJXelYjavmQy0EAx7Mq3KdkWvuKt9KQSFCdOM2P0QepDfJ/stiZZVPGH6+Lal6vuazM20TvQH
5xbxueOIqRRDRwBPCfZfZSXMriVdnPqixMj3qx+671VPyN4OqvIC5j6h63WAJJclEmj455gFxzrK
+dho+4M69npcNT2iF9aBKx+fQw7AnfSoaqb+nmJJmb7vL1DIps02P1PHmbuuwWYgQlyfMVyOCaxQ
wQ2emuvgnsdLN8zycrKFov4RPa/Duwwpg55tZHvKESzWEBX+j67BMNwYJcdxsSKtNoRNlwv2uveE
HHNDdCdZXrLWvFiVDzRzHA23Q2dJYU2Al8v/eQUBSSTtYIJUtQl9zCVXn7XJTdnCkeUFjQ4B6ruI
7THQa/STIT86xGL0q1Y3Jyvl2YKB4nFuo/m0CdS7XJEFlbpnYz2iW3P78dXWa4et662fjCn8MyxL
hIW/Yk6A6+yENKMSpjlJ0c6QSwXC25lrlShn+dn1rZpJooYWpFi5AWGGSg3bYQh9FT+2Ivex/k6t
1t5lH0GHVyP2yMsE9XOTsC6+DoXKO8Zur1V2nrPNoOzaQOktJJbecKEmtFCDn1fMTt/orpFr73OQ
RK1Mwu7/w6JTYLK1ZIt2WVWL7+ObAYskX+AJs6eKpdidvmIYBdGOggGomJfifYlT/V08e44tRgx7
+kUl5xdtnUuItf7d3AjfUJgptBfdfOeUH7hRFaQ35nFUDvXnxfTIsguwxU1MWfjY5p76jrrPtHAP
70qsuCjGlMQlAoJ0wLFHCUqCANiOhtNADWv+mC2vcOXt56u7Ow2CsAkIqjTvwfVpuAv+dNJqYI5H
9rrrtKRfr3TtqM2EC+sBSr1I/am5udkdudNqdjbLY0ezCHmSQRbvmZDfrCBcfXgRxMh2XXgyHa81
ejoch1fXDDQ0k3rwwNGwRJ8H0xIXMbZrvxZ9Un4gd44j4YlHBxoktszhcMha5XMw+qM88SMEqdKE
TnLuJsV93UHcQ7lQfb+nhEMlt+l1GeTm/I+WUIL6ylHrSobUp12ycDJxR/sssoipDsGv150pihio
KqkITeN0sPyU1rkdgSaALNaj7cHbkzG5Bb1POIp0pvXhOOFeKHMTNjjhPPUac0UpaT2TdiSmhFoY
7QTrO66qnSbF9G29O6M3orMVbq/Kh/rOSG+aiQG9Xa3a0s/Gu/E9u6kxvqm/O79hFmXsV5agiPr+
nR5A+RM7nX0B3pt4aeg6MfTYDNIOAcbMETDrL54YN+dtvOm0dLmiU3lp/irAYqEJbttMu2cgHtY4
D329dflbXzflJ6Iytq9Xf8zuBwoYj7TlBdBaQds+BrDFdVrrJuw/90jQBW2+XlS7fefk09LK0Rcg
WJopgcxf9g5ZhJ5wgWFau3ze2IcXE6nDnjJenwIeK0v6+RZZIiipWrEUK1yM03/6eVPVZZS/7Myn
dFBaR37Axl0UfpRYL1vh3YwLbUfcVbROgWSVw4aM3a6JwMYgdeAC9JBjAS8sumGd1moaUGnLzeQH
Y4cmi+3GySKyF6Cgr5rwptc054GrhrgqeKqbiR0nZzKJKRDOGBLJFhaveCyK3pA+oLvckyYUwWXO
fHEMthOTh5ikc2fKgvpHDPMvsQB3aTbvd/GX9eX6z6ZMfU8vk4JbVmkHoeN8uqcgPIMMBW3xwykz
EuAqo3clILloiX90RvE3SP0VLkxBWW0cQKq3UXlRkdH4bRQIkU2FBgzPESAvZBWpJTBu9mG/yFAY
bzjkN7Q/o7TBe0pS+rsngGW49fcjRAgs2gn7cfkezUQXIC0wszWatSEZ3Sw2hIo6nSi5e95FApof
6ZVG+ijGhAnOEcaxkUfGG/+i70eTwZdgeyWyQ6BWjtM22ECFmDYNedlQ9ZpizVsIQO/qd/F1As/w
xBBfwXAqKOmRcMInWDhK8d82eyAMvybORs6IMTjxFb1RDhCzmYPONjzRQd3H5AX2BwgMLMcH+Ob5
tQPmDGVKrIdtoNN9ADWoANlTUQDgT7FfRFhHQV0FeNpGPe2yCaXYeJ5HJX87pEgpfVHC4xVBgdlM
xxnDtfuJ/trAL7bYh2RbxMmmOJCZh/86ugteuIt950j9rcPvgZhSUSVcUQfWntHx5IGrj/fC1Lxf
Qb8GEIOvfLjtnmgIibqTuZznJEsLIbbFnkhBdC45rduGanAnRadLZFw8ot0gxJhk/B8G42mBTtW+
893oRgCIgqo9wlrNoVrgZoD4z0Jax7mPdDBM976DkJyUkgk5yf94KcjG+/DMciigl69fZzN0wCy5
qn0XpoNcP+yvYjhufoKGZ0b+piib4KeB9zyTcRw/RA3SqCf4s6hIymGnguwCgT8Ofq7iyYU991iI
uO8mEmjTQbw9ZmouS4RT6yHyFbmfbdj8KDvIIJT/qGZaAymED+Gd4GcRL7MI84yJEotns7W2pAzB
C6YhyeOrsSfQIaH1GFlgdxlpz7CuqR00AQiwPEm2SYr1ti2dbReZQFxapEfmbi3MqEwFJjmipJJA
M/H2HApP+nLUUKAkoPZds3NqdwRe6wOUM8B1VHELvGHWhL10f2CCMUTCqImFHmdEgG3yntVWPgSF
U0DlI/JC6HY/+ZVhSrHJ/1jC9GM8jutmsJfBWolyPJl/3BV0xCq9ajk2/BNrPy4/nxz+qrQIzGm1
jn75H3pYQ67Q5DmLp7Gth/1Y1FKlSnxH/MBGTdvhlMYwJ7qOfAR6BKcTBLcrVdcddHn7cLkGZXQD
6wrZbKGDrEAjXFSNDIH3doPmBj7iS0nHlI7Jta/N0mvCGxE2YjGkKlV1/C+wrKxRlTJ5UwEk8CRT
RlUIAV58ehj5sYUQ3tg5Pkf/kU/umBndT0avh4X9BwV1m/iyPZx+bSJrCatEjT80uWRrLLHVGvj8
qcTwzF3at39iFLTfNTf9aWGf694qAEJM8Sz/l4txL0aU2iqBIe0y8tGEsVFJsKOSmi9f3qHV+U9s
2X2ppxLjKPMSaH6oKYiatOlYFjDhwwvN6qXaXrGB25YYp8UGjUv4GAuAmOmKoiF2B+Svk+vKRylu
hCyWSWoGHW/BXN/rmJCys0m4Pt/4ufC1JxEjUqisc5AimlLRAMHVRSPBgwwaP7kKArWF0rCVpg54
TbO1w60TD5IVrew/wk7lfKmMURJotWxTVOJuT5d9jvVxTvooFKbr15EMXo7vCE+pcdtyS9uDrxEZ
Zl1VhA4flwK1MS/VE4m3VtlcCfVva/EHJYFD1FAQfjS5+MNeGYh+16vxDTfD+5IFffX9//IG8yIF
rYjG7vOxmydxFBvfNOVzuRzxwq5Z3w6X9PbliCgbLFhcHDCAHzMTctK9IUJYIwoziZUZHmAlL2Kb
B4DUuGD8yhn1H0EAJ2nfFSehMgkAzwG/8lLG+9MLhxJnxU4L4J/QoUo+NfUeG1vOhYjju8DzdXzY
b6ZwLpkrybfj+s1NpebDFkWqf9mMhwhIjnKoaHDLnvsPQ00rQvM5PRmZPgQVi1GzvKAO1wxkgUhW
7v3pj5HR87oXZxBovIlvPWvql680J4m/5b++qX/v42n9FNYCyEPMc/lB//wOZPuNyYTK9q2NrMW1
tKyvGH+tOMTPXYF6WbmP2o7Ge64HOE1pwuAlCyFs2aPbUHOxzot8dZHbIE6xvFI/UsmDr0MjQMUQ
mu5VC+RviSCyexCXKUg88k/3nf1ioJGqn4b/iDUlpOQkIkomxFMUc7SleMVOR0P3YwjUFNdhabeM
zhUIvwedU/FbF/WoQHHF3M/KzXyZtjaiY37AyC6U8jnNRgDaLRFgHxVYlEzktS+6JCx4u+PfscRZ
SGmZbaLF9akxoYem2LeRoDzgBVirCfbsVeTIIV7rdgzLWhjGCvKYlKkhbq4wQg3LGvj0+uhq8sH6
L1CrV3NbnQ7Pe/tWYj3J2q705ghGkLqn5kSxPELmoqSC/0H/bS/a1Nr3Mn+EzrQOkrzQjwadUXO/
sqHpl7yShE8Ys/G/16FFwny5J+9WV5t6yyBTdJ1hujFX1pRrCYICzSBLzLrz3YE6+EtEr0DzlEWm
Mvz48A2YS6FEOSq9baWfaxeGLGeYV+xTMrJyPyc9LtkQLxEP46wJnvQTllQRgGEclj0QCi19ydcf
xnvH5naNZ1dx+WmKWXgw56UxiXN0uwxnf7y0UapoHRX6Wqciu4YY1oFkaY2qfC/N9mt/1vGHmU8i
T6I6Tn6Yj4/YIpCW/1h82Mwuon0Q2aQ21ngvBSQlEQFKoYWjLiKxpR9vUiW7QX9+dPQeLhOLhX5Z
cj7XRKBuNETYXDxYSkBpWecMMoC8kVnQRoJfj5UCGmjZJwl9lmIuB3B4YC8KFzzskLJhFkf7IIAO
zRnkCWFRqVPps5CMRrS52R4uZlSlXGDabOtjnVwQnqaHQxJ/0atsRgB3Crk8meSaBUytqDu0MbxZ
ttnsKh0enUdeF3G6zSkeIJwOsfja7L6K9VycaUUUDYLemzCWaQoAAEb6VFp2Rg138KGtj8ArkNqK
3RDgRvNtSizxKzWKTyP/vqLs0S65cqy0r7oomNZu+Fuk1LkJpsV3++oROsFcfYglDClb4O3WL/Rj
6641KPXCWUaSqUj9qWYoGZtNwGcQCMvtsPPj0BAtryxrGS87q0Na3Vb+nz6HWZ4rCb9f+jH8IM1N
rw99E78z5CfF6LORI8MQc2X6bST2iRghrkwwWqy7pFhE9BI79zzDjopiAGQO7Vz9c3BGqRuZLzfy
sLj0h2m4GzEzFo2Nu09dXSpJzhWLbuM1tnqYhFV6VmAATa/38M/hILSOA6hiwdLpImscFPSQ1dhl
GkUA3PAHA62G/RLaH6M+J8jIVFjL6hayfZuZ8BG1mXqIqCHtGJDU6CppZingKSvuPymMS2Rkj/Yr
FnmtBn4Act+iB4FYioBpzJr6zU8TlQQzF9x/+PfEWP4F+pFalEpBPjpM7Lk9H5BzyW3hunSI4hrs
+zyWsbiLM6M58CvX7jmT6G7xA8NLR4hvWMPywTyRcjWVjJ39mKRVTZeMkX4WEc8bYmKVRpFwzjbH
P2oHfPzM5aO4ogXWck4Vgd7chbI7rgAnH+DojswxI2QXK0Zss7M5x4xCQgWZRuNPF8CtlEe7zAAi
ay29DbULetb62sZmKkztXknuS6+37INV2Ex4UNJD82XbXGsrP0HfCkQWdBsYaVX2HHmV6pBaOlyP
fwMkITwE/q+4lEsys4lYeLgQ3mgWD59Rx5M4XZoBH1elqGhaTbnVdGWvRK8ikRbwBtYKMc04XLwT
4U+b8cZ0z/tPDdIx3t9YZVfO4+zPvsuc5Y1xqHXdqx4HwuRQK6SI6mLY5+kq9ejxNsWxyR8lMLTs
9Dt7gL/uPEc5rR44eQrMkH6Y+8ELcmW9gZCwA+CP3xdAxNe4OLDbbIAToI4P92bz+xRSV0Gb04aF
FROkpaONKmSLgUtVUI5abAu6C2jQzUzSBvHFDiZhJNBTbwnrD9tYelb0Ui5OhT0sa3WrqoL25Lte
z0Y4mmKPY8q4G+W62GBDYVSTPlNNfQ33be7EizBBIJY5FL+Asxd1+QesEGtJ3ODcazAB6+u+noyo
98eZ+WFAWM8I/2VWLafeh0ShuR7Ww5MS4icYSJ/6REO4wuv/1BlnBcSCxpMsv2/D1XILfXqqCPjT
AJVaqvHEiCkCI3iAZL/IYEWhybhjDwu8GxBH8wOAxRUNh4FOemnqEvtnOJwumZxixWEtrMaq5yfd
+JuAV/zZX3VJhdWx92ZgWQW6bpRutG2Uae/IVF6wDdTp9MauDWWkJqE4bgVIe4jTM8ZVeMDnYm7a
JVex68vEnGQ/5U7E3SAXmRPxcNqVK1VFL8GspK+/gLyOWEud+0EG+XcP8MftfdWVvygW+0uYvXv7
b/56WUpLQBOP8ndZmLNCVd5ZJEQqZcGSKklak796wT5RbS1nuwrkYbL/rgaRnpV/IEUm20ITrN1l
Eh/4HLsY68CInW/bvtZMBJOThUzOGMCpP+Vo4VEtWnKXV++J30sGfiLr/uIswigvWCBxhrmql6op
WHX34KynkmU142ay6ZV5jLFS8VP/MdeQdUurjYwH8HeR8PRmEUocAZzoQ4f3a7ppMzEmsW8a++Re
kYCb1sBglgWwLIGhImUFQnGIIcrCN84cRNyw2qHq7UVrBaq/zLWzAidbj389wAHAfADkrlKx2jwh
cecW99kppkj1KCGeYePrZFkZZmpjxVuwuZVg3qfarZBLr/a7TuW0H9kBIQ+Bx056i9VvKlton0Jc
/OcwtddNw6aa3whZsQ/ZLRvrmraDLNcCeTNoyNHYk/WWaLkQebGYaXHFCBBZr3Jue83v6C+adZ7n
/tEyaNsVry5fYnrgWM4/rsQN9n9YGHcRbFl8vTQzMvB0QgZi9skQIvaKy6eJdeBYkuzq2sRGlr6n
+A2285CrxU2DFF96SoxLo7X5WC/SQEhbqRJ3/Y2nLgNwxZBGotvAD//K6f3fkzv1FiCpaIEBrMxR
9jmExfD/dZ7pQewcV65shLRE1pPgBh+D0QfszVPapDD6vH12AGMK9MkJ0a0cHiTqPTIpwfKvqy3c
ncKUd7ph/KFbcTPHmER+q/rB8ATY2THM45c+5IUaAlVN6z5o/3rjRL7RE9TuFzyTJF/bxP7SAFh4
bq8Yb139TLLB4msa6f+zm1UxJzaZOO2paJqP+qMIxl7Yvzx0tH81K6Iu04kwDtD7Cq/g4h1zUC14
JhPeVJiE7I+unQWq1rS6/Xnh3GRu9jopRt4B4XLK88K1EN2b6rQjRENyJNHQIsABj4KLnIxO2iNW
+nG91ArJVFVp1E9Hqf725MCz2qyUTDdV80eynl4NSz88FjPE+PF2FXk2HwUtJXiVC40ZlLVDfkJQ
MClB/3LAyloLgIiGg+c4cX8O/Twmwov498hxYQS1GYLbPlUqeoLX3jbSNrNWeCrf9TPFGbqbR4ME
Y0d0lLn0KeyEFdKWRz7N4laRaJ+FRqID/7E+ncGJpzDMHld6PWen4FNjhjMBM+pnG8sNeeTOTvlZ
l16nOl6d/hPjYmYhsLXFXHXEHvE1x4odrLSMGaY/FTPJF0s1iesAt1XN2xAauR5StHWrmInKSYww
Gb2I9Hrt3TxZb6sePwytC9kQ/buD6bbichDl+xw6qdD8s6K7xGld88HWiB5tzH8BVvOS8nLXT42V
RgONy/+PkTDrtEx0uzk5YRkHNLqqj9vgZ+EfKqwzBZbbuIbCHHqL19hoE1cJdfkHFAN1VvyS2K5w
UU48R3UKTPEj6N+fxr0ipYlvKj/Vh6AY+CpifBqDr6wLli/bWm+mt/9MuSrM1sFhCXauB4iyDf4a
SKoXXSRqepiAUPQLPXyAWawksiWGZcv7tMxZokGPaenAF+L9K2iq2xHM0iEPjTcLFimwfK3rFBEP
gefjEi1nVNyWN4ORzVIYcxq7CfntzR/BZgfH1Um9cs1CB3TSokNbY9ZfI1rdjqpx2LhFufjoVoN1
seMxXaxRTvQKzGpcNM4DvtwEDm2n7if6sEyIRXTRVRYw5jHdj6vHCxQw3f/wpku1Jh9A2Fdj7Or1
aIRSbDotSzlA/Cjc6Fas2jF9RzppiozQONyuifshWaDy37d+fklW1RT2S+WxLVl25hKPIyNVWXFl
NmDLAsLdWCqaEdZByRF4+VoFIFGO4IhHSLn622JphT3pvSnB/ztST6o8tnrJq/XpYJaXd7E9fta1
jm9WypZWiJeuaI8QiFKeOBNeYlIOM0ivQhjWf0nX0Y7fl+/5n87wtzj4t+TgthtJ/eObBBT3iN4F
VGRQm6esoyS7KBswIgP8yD3NGqrMZEBevjykNf7vKOz4976/78ehOxNe78Y43lNxHKqYcMl9qJn1
1bnurwPFkqf6m6MiQxGpYFE+gUHd03xZYBYV1hixSCdFxITLNVyniPQTZqgkpZzTo+0nAheoXzUz
n3HsRJnMDJAcb82eHRbHJ3bYfRbbiorIZEk8+aNE1Fuf7Paq7gqxrODPMpCtPFfzVwzxE4rveQKj
ybNqayEBlJ/tgNYz59ZFLYA6Mqapk/lBpMjbmohBlA6ybYJMPaBRg4c586azislgnwo2wTmUlQTP
OaeRD7Rc3l7HSWnprgKW7RNRwqpKaq9lHaYYgEGP1k8u5el6lgrH5bECU8f4UGiSpxGZ10fAH8p5
NKa4neuNZrpBC62ADpSrAd8PLifP+qpsJ4qiceTyBOe2S3v+fdHkYGZ1Gfms6AFwtQA/ZihyR85O
PNI1TnsIrnEf3CMV3qizstPAHsB7GBQhmEQz5pHjRo62CVRGNWOoJT5RMTeI1jYKjvp0IcN9RuQ4
EQKC1covWm+HLi0wngaJViltKYccRE9NbrW9F7SAjC2MpKJMtn97S6zPJejjFCFijaz4iifU2Yot
wQToYMo+g3lcIyK6ZfDT+MMvkd+bMNazaRtgoGCkokevExLu1E5piFB2yQ4egjb55Vp9iiiCpb/8
NUwkLsGH/bsaTyfAJ/1J3KqIxeAGJg8rinrLoeZ2YfvdSWqOG7PCd7oEzWMGkBDWdq+XEXFeiYkS
gmojkuGB8/EUfT9RMdvsQ8MK1tM2gBUrbJiHccghWS3V2FZql1iByHNxM48hjRZZ2P88xsBmlxnk
E49AvKRaI/bT/Ky5gytAMmTrbLXR2X/hqW3a9dvNbW77NR/TeuQU/1+SmK9DW/DkKFIL0Ymo/kv0
jyiWqegS3lVDxODAEp/goh2siikx93lKyuFX3OTXjPFjZipEaYKZfLNJ1jaNCcYzsiRg0fka625F
SR5GGpvAVVJJadT0KiV+2STC1qrBuM9beybHo8D02jWJxouNEvsV668/Acsso0EHoNv/slq9HIsg
a/s6x8el1+jPF2pZGauWXxb1YMQdiAps/U6WR6OpV5qQQ4HDSlscWAQRSFStvr/vXjlEAxxUqUJv
DZyRvKi9PvKy1X9fuP2ceiiiQdIDg7JDbhV+vlMw3ZLHqMu468zn2XsoAVZtWBh2SNInsGAI9FZN
//etPUP1VdP9jgQjNrp+CVLnTo9s6m2g0NrLseOzfPhHzd1F6aOTb0mSGj4d2ytPJHG3mXa2bYQj
GrRHpbHxYgn2VBqoM/4nGqQHHKovGP7lOo9z1QTNTHEbDDfObexB0gucUN1zsxqA2MljwFi6U5W5
3FttvLuW15nReInSOXZJlEPTBqsuhOpTJl/Iv31zfbq/kcvur5LhqPbEX9QdoptTX2pNJKboq7eA
vz2Zgmr/ProL8JBMtK0b+0Cif7tSNSSOmOdIXDrC4oPqdGxml7R0TIR4TjeprCCqto35slrmNQpr
WJUU6OonKlV7oAWR2CE554J+2WNZfUUbYnU4DHkahrby8IlBmz6KdIIy1yMVWx09qezp1KuJ4r6V
WAZgJN2gaHEaA/O9Bgv/whygo7U2PFP8TxOFrGa0SOPoIZltVV3nKuEO6sKONMCCO66AUnQwBvco
Z8svxxab8vqJmYihqQfAnVB+oGOTBBjpXH4vu2kJeofGKiojDGOwqRLhmwVpj0oSm/m1fEEx4WrI
7kod06udJi1y1nw2bECRJVg9rV+knPmbDLLBixc0Hbq7udjZb7kZUWbow9CxGzHGJnVkW/eMOq1n
2SrLjPNlWkX9O/6WSYLnq2VcSNSIv/cJbeemZ99hSYPUPJj2ETVyM1XFMA0cHSnJpp8ftOkrHH77
W7KG/pVZ9n1cU5lMN4mtZ19Q0/Xc7azcnN/82gD65lgKpOZKIBkt8TV9TXl4WGS3zWRWCqW5evEt
i6K+stCpeYNQqYeckdsma+P7E3XdOsyo1a5RtWssNXMfQmZdNZL2lkAjInCH6Pv1MiXNh35zDjBy
sNrpFpHd55p2VU7lxgPRGAi+oipTGd45d1wHt43MC6MGOqF35YMKAlGOCSgCGZukWgdG0mc8wdjf
BreUq1hPpgNfXq8TPomDqbBBICiNYZr43vsyoaCsDe8W5QCh3GVR+gWuaI8vdd4rFzXpf4XMBfnx
pZUnJwFekk1/YYmUiwAwwrEkwii10v20CmAN0dURPKxD9QnfpybwZAOwpAB/5HpHgee7qnss3p8e
Oskl3mLo49hK+pAArjpzCWccAwiYwLBFwb/9QFE4l7KyXrE+ML/UFU/ePCEHIbyHwsHMdsgAGWeU
9RXtFY71s2rjJYPMeXBT99I8WNesrftHNDi7UVNQMwVc7vEKst5Uqm3fwHD+fOybBIC1lfB0D99v
mSQKMbxz3sRb3RtE2xi1fIbu/QnznNwJsiiJB3kscoFP24PSoZrgih5SkNADfhxqyN1RxYDqSwPS
MEir6R8igR7uLgB2PXnpcNUEg9CkFmhOBDHuXxFx03qx70utInKtIeums00+aZNXjk8DpZaQjZ0O
D7u8yk9kqUhr1pId9cW7E4kcXb+VVUeb+PA/ZsL0zfMue06WriJl+jzSnV2APZPfs0fIjhwL6+Z3
waUjzLhrK7sQMGiXJFLaTueGdwlRw4APajyy+UFHCLQCcbq3vhi3czOhCvQZxcb9zHjKMKC19nNR
fnjNlKDbkmfTtQw03MtAc8eUv8i6COdypeFV6dNaUGnQ//CqopLhrtQhNsClicg9yIsaphzIGt06
8wJBtga7oadOWbLouFwRElKvscxraozEIchQfCQHAw3aKcmJPuPexdXD9Rihf7b04Yzw6QLsH4ds
7gzHT0zzlvcOVNROGgL3kSYWbvMvC2CaEGivVmRlSq6kXp4KjcH8uQPHWGeHLeKnjsfgs963Ny7D
XxPzqoAWyCLoiMH/lwuT7++geqxcP8020e6oiEY1EH8nVsNSXEQRNXvz7Q53JwctehjRMWOz+spX
nZWimoljOC9v1XfcHfQWBxssCezJGzIwm/rNh9/TC9VriRXmmrtPZDbsMrmqLySVDD8+G2z1ybSN
4ftiSgn/CENlDbvs81gHcJ7b09YbZAiyomhp/9XTYwvCTBYAAZbHzX1NYyjGOTyrYgTVjPUQUwEw
m5BQs9QkBaWeBzAn1f3M9AN0CB3zEspvGebFUjxVdHFJQGann4R23Hp/n4Zw69gjlYx2xjmQ1Oz0
S13njSUWT0BOjai4urarII4YtQR4eln3i/P2jjUBHVA36l/TJDUVHmypTt7NsjrGIOc5TnCXk9qc
2RoeJcnXyAEZzrbmZhMufAa9kxDNJnbAUsN8IKUXt++hL6sqi53WqL3MvT8kaDEH03dGQx0Xracl
Ryi9Wmy+6CLNgofa/rP+VRZ/TcuXnYfPukxeImuc2qXTD88xwgXbF1E8xdiRfzUCNWuUinkF26UW
i1tbLQACDSjLlqeDkaznMJrsMBxE3NX//AHNcrFYj5niT7oJIVtSrrCEa25ELdEcrJv3p6CJ/cKO
9y4pUb2GnpzCViXMi3HVEc3cIz6nOi4sX9PppE/X63cJHB13WmJaghe+Laa+rLBCMTTJg1MbOTz6
PjQCJXs8ApOhhqrBcknoJFrJGDamh/S2xpQnjIurgAZovCSjkGANbU16W6f86aDp+LP8iaFdVzlb
Wh/iNWNFbbxI+HDSxN/odmxL1jUDvt4ODCPAjouryAB5e7YXi26JfpNZPVZZl0inr+SgfQD4yFmR
JG/oY+jhAAiqEOHhv1pB+uU8boX832O87gVk7sh466QgMBlV6/SFVV8htnFc8C5x8VGDdmeHSKdR
h+iOCk9ubvzhCwLzWrSOMX3+d/eer2sAbGO3wFHuVO08TAtCPWnZLLbT6GM44n0xlSLdyMnAsgHM
/YV6K9a0dz0co/PQN8GkKFrd6bKiwSA1FppO08AdwUSoHu3WlfjDo/oFHzbN00u13oMMyB9NmDkt
iS3aXD0gTADB7oQnXScX89PRMvSvNC4U/M9ioyQRgOMypmwSUV4Sxk3PAH8TMG1xFY0cKTJKgwYO
zM0bCsOS6IzIO+55tf/R3gYb+rnWifrs0MxIQVCulAYuLNxdOxsCCDFZmUz6VaC0SB4AgC4y1h9N
zXNPpCZ/9kMl/g0w0KPz3YpsB5zeKOnnk4jWtiZH3MXKCxb9TX1Ekp6g/3yYbd07p4M7bRPQu/SY
6sKmhh8r0etgznuoDYqbn/uSl7NMCkW5f6M99Mct4xvZiif8BHj6IMcSHhA60eOesfbFqyTVKbTN
nHH0AS8NZgLnH8R1yG8yTV7OLELMLSVycKO7UVza0rfLC0j0Of5546CZ5cwA4CrcyJrF5q++E5Gu
KODkyM96s5Czwgn+in15Va/jrap+3jIr9C8+U5va9pdJLGUex7xMNEA9bP3DbP9rtWqlPRxw1L7y
Q1BaCYEwD/DbaE4sAwfK5Vr3yso3Ze9ecfgk5zIwsHb5HVcSGl8sIDytNlUIZ1RlrrmgdrF6ZBJd
Z5B20FLTA+YYFpjErhmPBs5Sde6At4gqUbko0yq6/UlJjGn31Rb20obqngnDX32/JRZyTeh7gcW5
IcqrRMfijjmqZK3Ptf9rQ3dQi7m8jOxA+C57lo0SjAbBGVimpMMLGL+FY7+gYP5L0qhWhz36ZG+X
RKdf6Y3mHWnfvtOl3sZvOIIKLEyQM1sjGJyH2VlQw17ay9LIv9er96Hs2d9i0uJaQvV2sVu+jw2d
lYxct/EuEHq79g9z6qajOmzTXsniDuBBC/TGB07AOTnRE0zF2W9nJ63x0sNRJ7Oevy16QN04Gqxz
D5+VsaaIJOv0JDUmNUSI6arzFATlqnY3wuSqBLiNmOjxgJzk/WcyBFQ6jShMXytp7qZYedHOl8wl
FA+ZwrHSyU7qtVpwuQd1lg0YInu92FSdyuv62NuVZfKA5wwALNTlkRjHtkZQZymOeITn1UEF2GEL
TnuQem8ShRuZQ0LjZx4nAYHdyXCqNC+DbobYu0AWDRQWm0sxgRLzlcaYTdb2/2d6BkAyapEx6vOX
9v5Zm+4YjmgmLY4l40W/wrLXh0ftbSaM+A/C/U8JaeSjYK0MBLu5SQu+IiIw923BfMP7ssKmWKPf
7HOB78pMgUmqdx2aULZy8PXJ9Lf1j/E4CqnOqrEg7gnFVGMYF91bG4qV4pH2KtcXEQYuegQ10W82
HEKMMW9+6Kef/THlTwWogDJyEFbi/kINa0ikgpga1DZjNxY+Ni4vpnxet5sQznzYuxPd0mHoJA/1
rRHrV2e4L8KLASp3wg0DXRe1Bi6hW9y7tT+tvfGssciej7W7fSam3nqeLDjw/J8woYkGitwURzSq
iyaadzJfGLyzsdX6JHWOw2nL/c4qQjNq0jKdXW61DK8hTo7vDU4M461ogWdzld+XMu5dIY0/XWsV
TJ0ZDFnGxD3Q5bUX61SAiQt+KdZ1/WXPiTQ+2xsji62O998LSrCXjOcUCd8Q7/MiTAi6HGKYz+At
gXQJLaYuhXLjqjV2UYXsp1+ft/ei0SGlD7SxIOVy17fkk3HNwuEZfv4SjLjlLwS/nSaQ8IasoWJp
Vk0Q3gdlYECdXzjEr0ibshl5qpfspl0O++gRyvYtjd2cMCKzOIauC4g+uim3wuVN9XzxAm8DthJ9
tvUu3J1uUUUrwCyrdqe8348+pU+S7mOKfndoBgCPDmGdgDCa1oVYZoKJPLUu/FEWfC6duY7HXxJR
RftJ60UpSNMa4MJaWX2BL/AACWAfuYynakgV6cwfc/xM3E2q5QrdVOVlr5FI28/EK2bQFUHYhjl6
7htjmeGEI5ZRrqobDz33qwMPa371TkErdrOnCQUyewHFQUZk5kRK33Itm7RNqxM3n5Cl5Kf9brCZ
GTGdaD3IRIoF3YD9uPzzUjDLIg7kcNYdeSodysQlqfMhEdutcLLTKmu/Q2vQwXNDlnaUzScOPnwE
V3V4kkwtkFB0lj+fMZhIPIgxb06ZmmywLCYvA3DfcI+elkQ/Rq28K24yPrIYbK07L3g8sZV4qjfR
nY3/vPW6HLnQ//orx4po5BA0xmtzzvzG8RBYgoqkW6Gc/YEDD3OVbZ4oM8MQF0+flyGA8y7YwPIP
T9SKNJfSC9VWd74UPSOe8c641FTPnUJwrN+mOiZBdLpDwU3yofMtBxV6VDmOnm+4FZqakwoyqpPW
bLF1UQpju1L5oigQWVhcYzDYEWBSrnZijpJTd0vTd/v75Y4ouvVF6D+NJCs9DNnEnNBTu6kFhPKl
C68UHySDhHmzDTMiWRBXSJyEEPDQ042C9VSXcIKECMLkCovA1DjEejqrs+U7QwQGjRVVUv4w+1H8
/5pyKy6kllMpOjRwqXf/OpjX5XWxx92eNckYR8qiwm1HAn+ESIolmR6kN4BR58F3L2/uCSiY4i5d
4NJ10kV3ngtTL6qIV7xFNKd/DH35q9jHYxa8UEyH+mravLNddwcxRwd97p6USXikLNv6qb7ElEhL
uh4tRYqYbXQjFJQyvwwIRgFg1hCbrnBQjc3DH/aUOY/MFXHMgF/cWo5lEBm+IBtn9EIJm0X+lzV+
2Sr3Crfr81wu/C6jp13fr+M6j+WY/OFfpxib13L7zPvv1pkGtJ3sfFO8wrIzhAHK7biRROH5s53E
MqY0kzLrAoUqxaJ1cZRG35BRrxlqa1siYX2mhn2FjCmQ9lL1dHwacGacFoenNSWl+sF5LWdwIsJo
yNxXgKpaN2TXgGKyQVTAm1rAjGnWdj7y9YlwhYwLZbT7cKQZxX15G0n91gVQ96WzxAXHW+iBX6WD
4kT/8qqHpf4Cq1Hhh8SQz8qMpTdegwcQ5QAx642N0B5S6Ad3bha0vGXRBSuRgngLg8VNjHWpIBc4
JHRmS1kN/GtuU0sKKFTRs2GidTuvP2Rhsva+1T/2qzF2+jtcS9Hy77B8w7oBKfGmVtXuSobcgeuQ
cb7djVqfCKF7J7VRC/0e1jWOZw2Thzrb/F67kDXhO08W5UEWKPkZVm3vXduHQIEEVuPECTk5YCg+
vn4LtIZQ/Xfm+xJxV386+Zzi7jhD6iV8plEmNwj3P1k9Gj7UiZlayapwHcnwr/b5BGz3owkrMonf
3pta2gvYzPeOJHtcwpLkW6kSgG5V1B4OEsoD0NYy0kqMeEgyM8+5oURsKhaHVVA3zcFWGvhWVPMa
sDkLEWICL3Zn3pwEtxIrY9sTJOU3ONZxr/lVhQ3wBILPBjblLXRbsfJbgmd0qlkCl4yD7zyNkST7
Ra2pXBt04iDQ5GIJf84OQYjeXWIraEPjTyKboR0RA6+Mlo16frNtVFBxzAMsa0Re/NebfpT+TMwk
jNq5bqlJGcujSRO4wIJfM3xo/kpmxyZpJx2WNCARwI/gHXD1D5rVqEIJ2qdXlHF1rjrFUt1UMnn9
Vg1W+AQ9GYZQuvXmIUW6H875PXKI6Td0yGtuaLBxTFbENvDVMmvVxlmRrcw0QGMTkJBLaLHlBwhb
yWwrmXbGPQGxhnnKKyHMkG3NJGME2BU2CbJMjKycnGwrF8DPkadaCLkHJgKhQ6/F4t48CxxuOSeV
1LdOfrhSNdQ3NMHszOo9y1fnAKiv1KJp5NW8qI8pKROn4rYOIYfqrEV+9w8J48Ws234n2cbvBuOL
v3LVYx3BxHK9BdArNgNupn42PZLqclOciWjObmtozkkfzeVj7zyKD28aLNeyav00AExDbgtkj9zc
RzMU9inEINCVcwGasbfdrKJ8yak7guso3tDAPtNQWl+45qGndixBbkoqzHQKB5Le345AZoy8ub+h
2Y+HPNzq+RfuwDCSLWP3Rly2u4fwMtF58OeNy0bfMWctbI3Q0q/uKavWmYvZtK1Wc9jpNZMpgmSf
ZE93NNsFkcaG45+NDNI7WFPkZzfG2cC7ytwSKerV0c8UvPEjp9cLk5XYa7Z3YoX73nLxVL81lLKx
/UX0nA3JwdqOiAV6zWMmb25ZGzeSpkC/HrZNNfPev3fQMWG+WmcrCRpbfIsxVsxnoPD3Hsc3auK/
oDmfNEqelpGKWm/9nRM6fI6WJbQrgk/7B7CakTeAYnyIT9K4k3tfddQLuOsjZzOVEsQx6fOhVzPu
Y1Ys3qr+IeyGdwcL9XQY1ZSPpEp1C+EKUFK3qOTmDBRlSxswElUzJBlIu2wKFFkoNDphpc+wZd67
nOT+zE1l2EmLJS/tE9N746NxPWcDkFJWyOo3yS1+yUrLZ0EKqltg7e3y8ZbFo+7aEA82fU5Zi15n
2zJZ7Sjfj3pvwD5khr5GCosiAzy/zX/MMFPag1RJq0TJNuCPvCQNUmVmgHHv6lFZckKdJQouPow0
Pk0keiHMRpJ6I1lcTDoZWvFz591AYeWVRmcAegz2o1irs0zDNB8tAjDB7HS0NscVOneQjeDGoZff
Qi8d7586coxV1Ggyrst+Ghm6dCzKa7kPCPZinhYzisRRS+JeInzoipmk9iDaxorttaK0dDMMQy8T
fjDEACPUn8eJSbhVs5y2lt3qrOANTdTDIrplPsmauh2L1LacZM88NUqZ3NMaRctfzQtJQpCHVkL5
ebMYJHAjgOxMkmgjW4L1s7j8wE9VA6HaQaK+CMJifoOuLvrimHGdbPJEwurmpE2SqyVzcXAR8vS9
Ez3NyIGDujXqyYGe1NCa545VB3mvBrGzvLyvQ4K8scDxG6thawtY2eQ6JUlgvTcyFX393QPuzqby
a+Sue4sT3vKhSqY6d8AiIn8XDAp/NH5hRAaz+bpPXsHMRN2j8TDwZuFYPgL4nJf8j+HpZg3n3acI
QHV5UStlB2at9XtVr7OuFjNp/MPXDUmxaGXcuTJOQ8yQ/4/0yBJJ+BwDPWoLGsyVlwaPCH5NlbFQ
5lRPkHV/OZXyv2yPdl6Tefb0cytFC+b6W2BtUUpfACziCxiWRwTS4JPvROMcFU5wxElWmKVGXzuv
ka2teKr1d9o9IRiJJ74uviKHaHCG/pVimfgHooLLbqomnXAm7TMFCdwb/UX5vioojXNNbEn1lIjm
ReuNsb87hVB2AnvomBubrK2mW4smoS4tTZo/v1rU4zud9hH7Z2+HCf+wo8JNSUAqeZG+k+cdJUCl
yT+zmKSzL6xy0PJdp3XHnwb40vKLxDHMwzg8X+iawa/9UQNUBXPMrD8loPepmxP5KFEDTv1d69ju
yGopD/aR+OHnKvT6zL2Fjj7HFkH1/mZIOU8PqAuXDRW+MfuLYKXuK3xpjUBiKzzQjsstfz2nBPkJ
QapB8SHAFjWUIUJzA8h8g0/pshAErutPucjMJUQ9Q5uRKF6ePlbL1GF48+5mvawPaNqjqKrSvlg1
s+43vtLZ1Q+90eXWFuiGLaF2rVImey0vA/ZTpIMrjbm7EdBkFcSc4m/1vALmPu0rwwNTfviG6IfG
mkxHXWlTomglA45NqIj1jerK8aTT6vQvlAPB/9ulejZ34X43/q2VSVIgeUO5uGb0fZMdYSDMecVV
3ybHCh51721ABm/4js5nXGL2qAz+CTmgXMdhGaslF3Zyj3Llz86uQmbyKGv2hnC/+zIvxessSnum
oYvl3OgVUTTuamSXUQl4qDIe7AnsULR3hSpjHjrmsPtgN3U7hMwn0vYENOck8Us5gnKAmwPAgPCk
3Bbse8f9Sd0sfxbQPgPFS9aKBurA4v/CbacjepNhUYzGCJ2Mxx4p1EPBRA2XMvMHajgy/4bFrYmT
QWwwEWs6hrC/xKj8R6PSjyEm7ub2jMCqlSG64eG0DP2SikyLEd1DeyNg8hTYRSTv3bhotkCeFcsy
k/OhPPi7Y9jYgQXjTV1CQh4HEvQGY4YledlXMjMrzQ4dFErpocEbNa7rQSiXhEi+dG3IF79SXNnN
7Bp3JGemYSDc8J1ZEidx7zN3aSHibFRr/k6td2XoMvIuKSa23Ndr38B6EqWAWaGvhp3DgNtcOsfJ
AGY98i7mWKwSbaYhWlNiw0SmnD9oV6j8IrpNzZaw/PfZNc4W8rQ7yYQBcgJYmxrsYhNUu/RqxctH
u/fjTj2JXwejGxC7/p/Td9AXauVn6zzK5p74THipzRaRK604mWTv/GZq9P3l40DRFilBxzC4ml7P
b/7InPgPkuqyVGGZANHTQLIeP9i6IX1Ra0dE7IFyFlmHtPvMR4je6zyy8sqQAKnhI2tFpBWt0gn7
e7b7UD2PZ711vsB1mCiUStpc+2jOLiULzhiJIQtYS10JUhZCdBA79l+49/NxzoXa8kmROYRFdHNF
SiClgQODZtX1Qv5L7lX7ygATDOaGNTUD73oBTzdewixmb3PXMsn1qzhe+rrMupMEfETeIyzus/5j
Ch/O/a8SgGFENNvRblKskbljz/1QM0lerXe2EEFheGiwxnR61oxOMdDtpoWXX98Zlvp/hMLt/MBb
AU1ZvkRiJPnDpUDQfehRufgsZUP7Y7KjtOfzAtQ0hq9u2H9XOnswkY94IIMB7feY2vprph/KY8MK
sXY6fZIwrp9/+FMhk9FwKjZo4zNVfYcAMpVbRuohBxtXtqYhbSlnGErV8pWPvmYs0ZI9qPfXgnCy
wsKVvYstFqwfAh0LHdrywCAnkH2Hqrvfw/A+2OKMSwvAWBp1lQWmC2UT7R8NcSM97lXNS4zTCx+M
IZfKcoyQ75nngCLZMOcZlYOdmHl692kAgEeA5hFDD4Mq08GcspW1cvse7pFcrGdAkrzb42L5zDog
wvwD1hhksMrRNyAEEbrG/I07jFknRvfxLBQ0+FNhWoaioatJFzvJjMEsfvhL2cNIh+vP8uWcQ2em
uT9IOsVgpP/QToRYyeaIMz6D5seWVrxjF4O9c47z5jCevVvHPZWya/JuRB/f+L5owMGXk/kk1oTj
k9Ih0o/Ltm6rGCOCnP3bp4e82E75j/bnFg0WOgQyp8/2PV+9EBkDWr+rWKseo0iINQn77I6ddfah
zudZAEG8OdSYGV0unpBSp47ptAwnHfcwOcAbgAjjbG51jx30hj6YOkMCixEYn3lTtFMMKgnd0tDw
awnPZc09NQqmPJtcIZ1r15JC4mLKwZmjaxTYF2Qv1lUt9xSRV8grw9KsKX2VZHWgcqo0tn7TTNz9
GhXPnbHKC4Ca2AR96kLl98gCn2HPnoGn1BaZzV/9JEEuQZi4nIU+lhzoXIwmWN6m/+ESCeUByRCF
WOE1x2wFtLsVXBX4T7fbSA7pO9jVmfLaLowHER7nALfMfxlA9i/FsQgwfwL2fpNWdyCVVBpJh1lo
a8FEhL7CezSm1HwCJPL7IrvgrQQ1YfdWirj1YdaSacBHzWTaF2wRfUkUD88CqjtGvJ8TSX0kH0Ys
fq0nF0XzU8i1s7UGIoe5yJZj08OtsLLyxAZMfHxHyalxqH5wJmMQqX6VCrwlFVlNkw4VDCJ6D3Xk
d7EklEi0PRW+w3kplYTxViNsCmxnUmkH+EHO03T9DShujo6PGJOGMhpbMiOAsVOUT8c3OtLU8/kG
1x/RHgKN2LxWto1vp6gAOp2fwPJou477MWsKULqqPGT9FVwllQz2VMsQdIOsaumqku32yiSq5bl0
VYxEubFq75qbY1xpM+5pdHnkb5iOykiyISyzj76ba/BiOg+MYyvRSfR8C3Lfgol8qdByVSeTC9Ba
KOk533dhb+wS7dbCZMzb2xzNDmTT2tW4sm5tiZS3XNMRychIJa2ZcVRtT+lwt2F3utsq4yktBSHz
jNuD0xGCu7m92dIzyPjnmSLpIkBr+OGQN3DVLPFcqNtSuZ/t7wPsgKk3YM06URbwRUcDggiaD44O
02zYlOH3rwIJpk/CkEEWrvdGjNrqKXoxTTEKuqDZ6naybiYqFZhFxUpSA+6p/F5hNmQ6cL1wh6xT
FVek+rd6QomEBYOh+XRBTpzTVf5btG/opAqQu2KdOWCe+OxgW5jgekvhJHwjmpTiyVABMPey+AAv
m+vKQl3xd+kS7+oiCIMm4VN1PjkqfQXNQPcvoUXLxDLsF1qV4EbrpYkkPvZQPkchIGK9R0ucrlC2
4+ceOVtnuJowGPXmnwxKxpglWg5XEZffGcBfuHP5VU86P4JzkKzfHDH/TpUyTABqUtERPhONRT/q
hgaqo9K0Vj9viLsOazbqYLy8J/AF1Pn+QnQNj0+CyObMBokzaLFxDIuClq7TDATW/l3i7fZTcOTO
detLjP2x28HkxccgWw9qyhLsAB3tSSF93HiM5ZM3hoTXQPf7JEmJuKTwPsLIakxuKRVu9DWN/3rM
3pMY7eGKz7EiYzMqbN7EneG+fZEEuze7WN3KZRvxufFQjFdvRvNOnNA6dhtHCIUiemTPCIB9hUqe
P9BqC+8tkIilgmjeWxMXTaTQdO1F/U5EZT9FlYUzN39nmO8TN3y/Ogi9H0Nezjj0b/gQXlsH7kXQ
SfbMe1gZMzVZ8eZbTcQYc+HsjWeXUu4oqEv0Ra8l3BH/UC6AiRrPkc3s9xWz+QUQXBfK/+zrkLsB
kXR3jzG9xszqenXC52/XE9QYosvuwknokF/XVkrA+SBn4yW9DSZ4rWDwfxT33sN2pbSO7YX+pH/n
o9Xwiz2NNl6HOLKk6/BxWwLnH2DsGJ9QxLa0/5F8k7IRI4bJ5JZnnjZk3iRUcplAOTskbE5pH0DI
ko6/O4ml6awXLEyQYWPRKynZCM1PKPE9zxk1RIgWu296WnsXGE8QEHSG4GGln0DROnvZwvS9LJqk
4QcmAGqG94VKRLXTOS1R2RcAYaDlcJEaUT9ZwCxvp+tkB9dTPPs7D6AyAWNKDzjkpW/CTNQNmoak
e5tRWWUVCoFtqh1ybG85IzBFusB9YaqPkzr1ZpBHPlsThz7wUg3TC6VDdhm9+ECPL0EEmZmnCMPT
hFrWlcHL54CQlfaHQM7kqKrt9YxuIt9+CjbnqZJrfiThxyuT6BcxO8hoMvFf2D5EHykEM7RiR2N1
40ZzL7JO/REaCjMiRqpLcKKG7GJ/NFqIGSktfW+BG5c+KOzLCYlv9kY0oexRcU6CVWsJbIMmYpwI
oWvra0SaueNT8/tzoF+y9hlDs/I4XFmUnJgEUvwx/t7CxR37SV6OTga7NUSuVUh5Kz9k5gS/XdAs
wn2KFBPxMaONcVqL0OB3MyY5UJ3Gm0EjS6xwK/PevV5QgwSFQv4lpGcRSJ141V6KVAHQmqnVgCHb
fQoayk5Fgds1UeioSbwX7dDS64IIlkytEnwEoCBTQ9v6oX0K4zvtVVxhealXeitpMtAvuAf4cNMm
jiVL0lfGmtNj+CUqzn0PNTRRP+840LWHoX1aJDB9KtoEKm/RGq/cyaA++q3EtgF313ksnZiB7kMy
AqETxGpySIFQjXGdptz9MCRfWa5M5ikE8/87G97rT2pI+JAiAGFWcJgt1yjfqfIlCOyAp0/acPVh
wLvk0igY2M3JYc+RcGfG32WxfJG+7YI5wZOs57WhvbWlAIx6ssQaA/eauB1Mz+hJUo9SBQ1QFqiW
e5KnYR1kiINhvL5P+n/8WwmVg344UmkWCoomTKehhaL7VbrZb6wFJE6eQyKlveMmaw2/CK6MCZQI
WgOEb6VJLR4q5FulXuKvSHZnQ308ZHfXyy7uRHUZeHsxGvluyqjBR2ApI6/V+uIrIYrFUR/DqJoy
73J+9SpxWywuEhrRsP3oM7bsTs5bfue7WZM4fljVq59Hn2+atzmVQtky19qSsPR20REt1+GGKNPo
psmOTd5xDO0OmboMxMQL+oPV8s7sjv0a4ru3jms6pnPCVOY+RpdcG5zHOTvVIdWTgnfYSXniaaWn
AQQcK5h5/ejOBNxJ1oUR8E/hTHQqkbT99nxFRSA8pi2brbHCadEI3HkNF6upLRAQLx4YOESqQu1C
TCczmYHH2wGO98SxPSRRTNfOQ+aMjQYjyme2kLVWn/TC0zmznmvvfhwMq4mux1WxIaaz2agRnsDe
4D/Py0gF3SFWxPjNxOf0SyGIGlzDhE6blm0flbHhNA2+QtkCPvojMZrNmgq37JPtRDggCc0wrt42
MbRcYFusvFEvk+3zlVQWHvIPmlu4cN+7kNYrjGdBU7YedXZf0eQKJH7ZWDSNq/yci6Ytl1PHktqS
i3pvyKkNkUpYmHNhVKbv7QcdEUmxVdmlKLm4iBJDCxQLphfp0iIbTyuk3jY5KjaPBITehWFa5Ajr
+yWbgWArUSEXsPE8JP/hcu0sZyen5ijGjpLTU0719bzrRx89PW4jdti1ozYTHnOHI9XbbYhaU7h7
NuMTIIY6Ac8rP0qjYRe3lKekt4aG4wUcNoa1Hg3+vSrD1D3djdqjw/d1k5HtyCdedd2gjcsufkg9
bBBLQ8OB65OTgp5s/qEQjf9Qab2ZqtiNjWunVf3rvVaa6F61IzWXQUDz4FSdEBZy71LMWmTnS2I8
5I7q7rywIZX3EOp6TSFuk94qMyxHbLuU8e2DYLXoymwIHPjknkKEORJfNyprL75xSiERm17RWWl4
fC+p/p+Hzy9I+B/xv0GE83DU4ALtFN21iXPzbrhHU46qZj91IONTe+DXaqkJ6BcBxxwsPBpRhim+
de72G7qxUFpSrCoCg3+UIpO1yma4Z2KbeCmDWu56iktUbmed5J+THoO2JQl8hSLaPsvXpAfvxMta
DVPk3XRgInpMXSfjZHe4Tg1zWNO+eWPzmm6K1JSv22wgdBZHiIluKAvs8/jVbRqUubbQeLEmJyGJ
6fQaxTOPOO7yQIAXTns8F1lVn8dfV8hNfs4bryjAoznYrKVb1uCw5Gds2rbSTlcEdB+bhuCb6LNh
ehXyGU05ITxPfDOfK7xsewdI9par1DE0RCH4BH/uqGDAobYyNlv9XbIw+QC90Ug8oan0JILbKow2
BQpyPtCnUUmrsw5guAYPoHK+rIMC9LhcWUQXbLQZhW0xap6q/AnkowBZTORbxjRmmEo8oOqypPcP
qJmrdmJ69GzX123OD0SlDFxYR/Dtxx8cT5IFtaYkaI1snjZhb4Th0hq4MQuQE3bNPhBWMgRvRB2f
Lsj1N4TEv47hfYuVgOVI/ir8Uvuvao/4QM5b/ggVJ5R3ZvZcCrDGs8jg7ak7x8RBumzkPQU6wnKz
zs/M2ho0qtIHyqD2AdWs9kZ6hUjIqImzJ/cd2i61nI8tAy+ws0jL3rQwA99Hdj2ottNnQfKV4Y9a
VFcWFURil580ioWlaTLO4S0Nr8991k5R255VAz+WPVfT4zttwB/Z7+wik3Tb8vf0diuEt3+a+jHS
ZDuVF4SO5CqvR56dUVFg3Wt08qyWO5ND5eI/+85BEAPSZztZlZwW/DkwhKlUil9Flebm1IR1W8Pc
2384ZLDQ5c5ZNwGdMXPRueaMNn+R0mgo2+Q9fDMBHDXgtayM6uMOawtABJFS4LlpL2g9WkMrYpxr
eRIoQtu7723WfwyTD53qaRG1ERKfNDssd+44IfGNK1UZxgAyoCf4TOlZu2RAfvRu6kcg5KBCTKBf
l70wadkOnwKBRE3QvMx14CxBc3uVUbJDxAHDsJK9+KFDseI9AjcQdFqTiZO8IPsXop7iYMm1aiEf
l07TFI09o3jLWpiQ9s7N3kqrgp7FFN8FTcYy0AZbYgpOQbg0yOw5xCtmOtxH3wkTmvWadx3paC6B
oqKmKZ9gz6ew52B/0JE2zR7w4dQqvtXAJtmykK+1tYo1fCKzoGzR2ABxlS5LOqxWLe2u67QVyUBb
574weI5QR5OR9LSqFUmdoR9HBH0snau1hKWfyEXyYz3/o1Hmit6Vn+62eqlm2a3fkRkNn9AExBfi
4FCWm/vYDpiS85N7zaXRhU1Ae9Mwook5o64vJrLNcjZjrxBOTVLpS9Ri0AaL+agHYD+fJZoi/gUQ
bykZ6G+nJG4Ww+0UMegmyLyaoRyk4JwhBcthD7vBBhC+OB6G0w0PNWs0FmSXQ1J7x4JF0g4r5g9m
qQP3cjCgmx4k3No0f8w8plocfX416NCgd2ecLZMvTxYRU/Af2BWctShqZaCyd4gQL2DnxKzQ7Gb0
kEBUrqkYhEoQZkxduoAmTMuOvw/SNqYNop5ocWoBhi7CtZYSMYDaplNSlxaskqGP8I4ZfL5zO1/3
U//o77oJB34/QeKLOy6U9Ub2HoCZlDosL12GY1ef4SjOO4Sl9VpcIjnKTmkdWtvF28QLRO7KiCZc
nSr+FdZG6r6UaWEO/eZ79DrLobg4u0+gXWxI0VCuqHvAOOXfIuQgaFEvVByaC4Bd84Fm+mH6X9lh
iEsFmHZVUrxcJxFfXSCiKsxfpmIXlnL3v3odlXEo5XVNlnj74gWMpAtQ+9IpiJdaV4nF2GMlX4Qz
Tbb0NRZeZA2yMJj2dkiBxFB0RZrja5J/hFG5qOLMiwXweZwT+vD7mFdrnPIJez02jUygy+oU38AV
JbUbu20VAI1xTCM6Uc3iiYa9yyB7YKU14lN2ZFOSgtFkT4jJ+OthjgVjYCMFP2kGz7n/ssM1kOPh
snDtCcBtClic/4Qb0qra1i2Sga86WuVTFlvULXaF+mtUweO6EtF4OPDHTddOUhZuawNgSE5Cv6j2
mp9v2rDb3T1NMyrOnXah1ICPZ7iblFz3HdD+Mv0dc99jisNgGJrUBG2qVF1yuZEjsOLrCJcNVEtQ
6fdmwDzgZLkbBYHIi398JuTG69ekhP74EGg6XvC/PdcY7jmrPC9G5uQ82NG/Y9r185APSjnUmki6
nTt3J9X6OYbNdq0mcTdKKZ0JTsVxisw1OJ10By+mHFgWwAEHzJ9KaSQ39i1VFv9YrOIJ2BH3wzE+
o20ysG3/UnFLk99UNmMk/FZi+XLpB+AzMmFiTQ9JhNgpi89HSXDModGbRbyL4+GCOWYoubAiry5Y
pzqFMWp34txwqYZ0qZQDHI7XUkoHwyb2h8hx+rEgB6HTEmcHtTKsZ+PUUlHfwjHj8vjSRFgg51er
BzyDGOz3Ap8apvhyyXdX3jpcZq/UZgFSLe5TZc9fCQMsNWOHA0hmXyEQGwnhmN2o2qW3gMxZR5Sw
Ah47BoJ9ZgywTS7IC6EKAatnA591Sm0ciXab1gDZOCqlkXEoj4NP6bgAKUnGa3iZx3XMgWwDKfHt
BZLUehBIzESFaSZwUKPJvmKpv5lvYjN/f8QoHmJCXabNbjyXo11Og2gW66kp1tiwwoxppXHnsjBe
offHfAX6r95ODECQQxEaG3+c5JrM2ul8wGXfCU3UZGavPeNh09VLjQMPRIYhM21nnGg135eVd5T7
yZgWkDlYeDv3zG3Pvdg61r6Whi2sGcuvvwS3mq7RDzuixkTyDu+LmC5dkNdIBV4blb89yYakCpQs
mhvuJMPpftK9x55G5nuFPUmQteOq4HXQJrIxzm+EI88VnXFocZrYPnH/omvWaikJx5ZUzJi/RmDN
1df1XesH37T6OAiIjvkW8cPQ/xsSRvFxgMRUvXRT9DmnZq8MGpKAQxDZd1o9t3rgBzCuyBa9vA6c
VczPUKV5CDZ32IJZETEkE5X1O3g3bfpsCLberhAdrVkkAboNovBArCvusPWLjiwBwgcl1v/k0Uqs
fi35naimFcBnfFGS+7LgXY6p2k/Rk2ee38MYTxHGC/PliJ+z+LxlcZynWPh0ryWv4Pl2buBV/+qN
i7xeLBQCZYrmIE+9vZfBaYWmHFzNH+di623J0dPvokc+WyLo3Q3VtmC70j6sWSB7HUcEqv0Xa2F7
GguibeUPtnDxbQKmbdlBqOcqu+poEdVx++xFGVvMCuzO6yuCKWh68rP+f+hUl80/aAxqp2k2GraH
G9C88rPXn006lOfswHagV1FVsW9sx2XnDP3IGntIOk6LoeXGeCtJ0IAFt/tgTckqXDXG8nsUQqoZ
YohgHRW3SShhXQ4EUqFvVJmlnkg1zPZk2Lrat8bMUZ+PaLcSMrylTEDeANMSgf32SuiHjhj0epjS
q6NeU8KsAyWHncj3v+hHnVF/hXeT6TZCIiT4IFGySv5+nEJtbpDvxxvFMIsqHtp5dAzFmqJb1Tgm
txoZfPnW+FLbS27+DMyRhXinBVpmmvyRD4NAgR4Af1CvdO+hGZXCFElQOnDiOmZX1xqe3QJL67ra
l3hReNSvmY5aDGYakhxPhJ2bVl5uIgJZtYP+NSURZCM02oZ0xhjRhc1Eziymf7oMtqC9HAlpezHx
LgWPteob5ShTri4gnA6pjqQJWqRZv/sN68cpMgVmstTgMQ3h47uwC4rx95cZHWTqckfT64RNRPXb
beOne0xkaEgmZnh4P2VJNPC2Vw6NCPRufd10zbIJNaZjYD4RQ9hsIx7HT9Nd2f3Yv9cK2DImBna6
nv9LWI+IPblhfJf7wO4znnZw5SQVFAJhhJxS3fLnC4mIMHXDhRPD9c5oAcTzkTdKRDliMG9xRwGX
Ef5iAM5VRmFcd5Zpk8Yty4hpi087/HFJ68X9SUAIUBtjBlh5/2sn77KC1+2tNvt8E0Cgg7XSZOGf
8InmIK1QUdpM6BP8tuJwlOn/WSdL8G48VrH7KhWu/3sW71B1gDJ0kDkBB8i7oTNWd2nMfm2coVIa
1d8PxWw2EtQ/FgJhXmg8KeFL+dxvJrzCv41rs7KEblCiIejdImiGVFToTJsujTG+jFIhbyKB+xA4
g1LrsgngsXq50j6No/062tLnkrReNC32tUxy0u2ZtWeRGZS1KGXSBjt3HG+H98b4DcDJcuZUDBEo
tli5q5roTS7tMufX5XhBptcfhLDv51MvXJTeVSAPz5mciI+rNk+1O3kfdDkTqXcbLyigJFsBWB6S
eDNXP72L/ZvkQvKfe5fH90VmkRUMCZQxodWCWCKIgWQOkE7C+2ZeB6i2wY3i5VjvwUKKnwQ2ay1O
P+XW+00ACvsLo2e4FTQuVfGB2ZKrP2fxz8ZbCXDEbM2RU2FhkZC/4L1RY1cgS2QM9wmBDWrYaVkG
Wav8lbqnNS1JcWFg1BWNguNYIxI0NxLji7fqNMER3qcE0IZoDxmm7jlo44agobSAagoHqZskDmHV
gwqVl95bI62unCFa55djcLSPPhtz+pvQudaV3lzDNUhkFll6LB+r27fZlnlb9yBECwiDHdB5Evif
WeYcdIAIF+pNp9hsRuc4chHzzjt2E95gZmxOt8PsEcDkhFFJKSYcmSIcgF/ZtwLHDS4FP6ltIC0R
4NMG+jFaAuErc5b/VxyiF9iAgHCmUo4/XUQF+fiLUAYVDgs1a/sjA5RmnMlkJHhmeq7gesYmQ//u
4+vAertTGKlpFn+RUpGsnRizsP/dTSar7qa8+DyCChU8e0TNbWNpKEUIs+2Ft3nxLKd1CGnM43Cf
EG6hyZhNg2A+MseJ7ivYKs8czu/d5xbmsI2EkceCgaLHyFQ9PBLHrLPmAZgAsLQPxiP+Ln9fmPof
MioOC0quNExvTaVGHCxbyrCw9yUQM9zOIlQFFYaaqO1rifVRb0X7HNS9aFxqTTd4ElYbx1wguq7G
B8MIgnabKThiRA/Y1Nr4+3PPGodEY7C0ju2SyFdVGW43hLUGocxnOERLsWoCWE/JCKuggFGXJaRl
5jcfPFCnwjs7jx7ja4BELc7NwBsgfRccbg/M2QEhIeJ4RwjOoAEU6GWu3q1UMbq9ybVqJIpPGYCw
juVaBVGib1gFSLyycF4k9z2H6ZDTSIO5/fQL2HYOGG4P/R60oAlGU1KfXD0ExXlQmEEaoKwjZQ7o
lZjKLKuUTzBQX0u34o5A3DxQpj1C73YfMFBRBttRgYf5Of+Fp1/AMK5aJ9+JQ387VXIYRnslge2x
zqIVbkT4WxaZ28Sc+sFeQl7/NVxjEzlMw8wKiAobFM/YWlvgivqm0DhCkyX2VbHpMHCEnhxlyuhW
FchFMC5rk3k8wt3KIs7Iu0WjWazXCztzbhVqJWNVI3tHOzLmovcr2JJhuV55cm/JWnjWfgNx6O16
4jWrHTv45gSny11AjJ2VGbRYO2q/iXXq/IOBseBB4GJdGSuwzqycb+Vn9arxucxo83EULVYbYfGa
B7mPY5ysJvNtsaUa8gWFEw0qOpVVm4dzaKdvIPHp/zO6HNdW9MSgacNjwX7QNAdWl/FkR4TVLSL4
YEYK/8jd+i1nViHSurA54LZBEWqejsEc025yz0uySfaHDsKdE1tKH7gT3w+XXwEPkBMsDYYs1EMc
4DnLfrkkS2bCHM2MsZ5cE+pcA+Zl3d7OSZ5Sk7w5buwA+DNHigFAB3Bv+escR0mo9EhXRDh1xnMS
64lgj5+x2lkfqdDEBj5VePfzZlOANcUamG2BFoeWAmyNf4TgMmER2jx1ErDDcKW/G9XKfWWkvTee
J+Hbc/WY8RSiwzoBn+AwuBBiJWRokcwFLhsObgrPp/oBvjEwZFvt9cvFzyVAeh34lwvAunUnAxi1
9tHUP0L47VytP7N3KWUgzdwzMAhDjMEVKEg43G6RM5uZ2MWo9nBZ7CbODuYokpvTP3+fCuk03JAw
jenHdV38V/BPKqy+YWj9RKHYCjNPTBS/X3XfkVLz59eo7sBO42pOn0XSdaKMnoLWZsxwolNWQM25
Dex7zYBWLUsU0ItotGq8GawpQVk1z6IUJNE8EnCZw0DRFvRdihM2pNgzQXFR3+yN2gc9YuoB3OvX
x2kj9EhydsgHD4v6enYe/+NdZsLzr5pUPvNODEH/5gUUupDln8Dy5ymMwB7KpOKBEMCRn1b2L1bD
bXDDAhZeI+xeZ9GZVLfiPYhAnLwnlNSHBwQMD0oX4IoAF3GJvdxwNTfJlM52Kf9fC2o3l4gy+/63
4clErUHh7x6nGWQJEG9K0AA+VDcLBnAWy8obx14yZ4NPh0njZeWoWRex+UHfMj0CuxTPeeYfivVn
B537hqbZvuHjLfKokf06CD/r+a09kIZHJaLWiAPfHBwGY8KGD4CRnYZuApCQ+NadUNHXIllUKhK+
mschK3dnP5OT6AdjIXJisk/AdRCzd6TzBEpOeCJDm+UuNYKaDClEYFfe+1WUyW1vMzd//W8YmCsB
+ZnYR82CZyud8yThBYWKw7L89KOWkZNfYaZbXUOTEtAZiLR+3Z4sXw+ZSV9Bk3K3k1m0RCzb/A/b
3hC6dmJkYko4RJWAofQjkSS/PtC0E+4WXtu1FV1N4AyYYO9zMyVBe1+ZSRL/3qxL2CaqhoUS+atK
L/8C998sqyAfgT6rb/v6Z7nNt3UHHWur6UFmoyN05tR9X62oh8bkUI4OlsTdtUNf41OuRFXVkca/
j54mw3dpmWwvZ5RGgqZHTYNNbN0nyvoM9Hi4IuZuv9KRsPFSvffJ+xKdG+JfqMqIKuYj13OC5pK4
nkp1WxeIcXiMJGPV3FECCkQ6XLktDtFtJyXXD/pF5zxiyp46sqM1gjEuGYXpJ9T+qv+nKdMHF7iS
xMAUp3NKObPvPuzCDxAbThc6SX6R7YRX+iQ7exD2C/R/VJ21rnC1C7vZRd174ykFYKVWr9bkcjsm
kRUIavbqPtzpvYPyGI1x8yTf5Ol5c6yzy2Eohk4YOaXtrJ6QTQz60EZCNWY/ppY4kya9fpKkKzTx
gUwemF46ZNLD6rU9wUZtAByPPOQ89tnlLtMBBDm2cI2agR0spmG2p0NPBJI7pn3McxMJVayrQ8VS
OsFkuLUCJ+Tn1gAGcFIgwc4rI6T0Kh9LOLBGcpV8NR1iXSH2mJFHl9VhJ0+38D79dGl30edKtXXt
BDGQWGXq1k3TFDX0oAcWtreCrjAfQ935zdTvs83SaTXHtbI/bV0mhJy2wiT4p0ExkBTJYDjuMZPq
P0AYYYOYdkP+syobGqeu3ijFc3hFd9L7WDwuMsK5OSuAeXBKJTXHsJHhe4qBKwD0gDFdiYTj+T+f
SDwlb9upRd5saqDY95O3sOzm4du2ETcWd+w/2i7o/HXW/kZog+0OY1mRJzjnAeeFUB3Fbxt8zkYF
PgT1O3OWGtOdf7UaceTNAz/sLuo7epPF3sJiCTmlbOPEfYoLW1BDsuEqINyWQaaoWMejpyO2pD/s
Gwe5IBn2MrcUmbGkj2bntzy3w8XqZndcbu3olqqFQZCSedFNKxDsMQ4lnW7/rSIMyaPxbxD5KOxp
+3nYipUs9UvbjGFQrbVxFPavR0QBo7YaeXhYGL7C2xl4iFjMtrDz1Ke3LuBvR8jPg3G6x78VvPWz
IHEjTSYJ//2juNIwU8fvTKi+JrzgMmXGn0KhqdVDYhFwKJU0PEp0FoWgrAPPb/Q8w1U0QiZeOLer
TVP1HzP9qovQRwHsVzTiirW1GH3Q7GeRjnC3Yk+EM86fKrcQMRrS7MTNAJhTB47fLj25/foHCNC4
OEhrOhbkilKkdV1qmKMQEKeaefA1fSfCSlBF7XoOHZWfTHxwbGlAqODBQepyAeQkzkWRghC37AoL
9hG1jnMKU2eN87Xkg6NnzHp2d0dheUdnOKlIhbBTP4iidS2goe+nKMhO8jkXpHoGwqp7QyveCitx
dtkQcLyMP2qGqpkLLicHohFKb75etWAGK0c5xlBw45e/xBY/dRPSvamfzL6uR+mjuZVFwtdDGu2V
Uoopu5a+KhLJ8Z5lGY9MFEsdhWL+L2omk4yVGUNEa+rHAsDyT9f57c7sqWOuyjm9Dy7Q+ZIxJByh
DgrCaxZcJbvfOuF+6vT6tEDZnP+/MNlMLDizdxwUWGouFsGl45vnat3MR/4MbLiNi34U18zPtJVM
9jLMSd7zGaFHBB5YtfbDrU6FnOxhKsZ7IFi8+FMmWaQNnVIqJG7jHFnsGklHol1Xicg7qDOovIDs
8t+fPCEx7x8iuhRY2jHWqnVqbZYrRhd76CPh388Ev2r+3sorDGVnoLOGzP71IfmeoTHyhLFQgOG0
8mUnYj6B+RWITs/UoxQ3a3/GTPYMvHLN8kSb2vMSRESp+uJCnYpzl+hTadoFeOKbjCatFHSbAQC2
ge3O2IXCDfmofCcugsGuoe9mdJzQDUplVTjW9OigoXpOA+rx2vu9sxyGM7SSZLL4FMN4/EcRzmub
nxaT3SBgzSbJIXnfL+afDozI8s0m34E9qaForNNFYzvW9RHx1pabcIIxksKqn338Yn6z7KsaLxbK
gHtoDnn+nIumvWOtSHjzENKMk3JDxFQHkl1gfB/p3ejMscgvyMTKHDjh7LUP3Crg/c2/WPSHLvPu
dkweM3LPztIOsQfvkIS3XCnWM7/AKfLZNkkaHzMrnsCD5UHG6QqeYWw+kKH9h/+qx0AIZiRfBa18
j7K0adcUCcnG5b9bjzwzhpIpL2NGIo6j4tbo8ch3myIs7VT18lqYAYzUJgu9N89C4qDoeursaNTD
QkR6RkDP+NQm1Kea+qV6KBMc2OoHDYb44noV5HuEblmuaKc22LetmTFQLZioW1XncWO4yNuvMCuH
RT04J5YtEesEzvVH0nAbjzFmEk5Xn8a+HT0KktNjIRQH3Wz2G6kQ8jDOg3Hy4OqqisTLsnSivFKR
C2yB4zWIH9rs/gEQpa1TTs/Feqz7d22WPWeKW2oCgNeIPevs9Wqi40zrFrVeG20LKvmdatvTzdzp
gtFSP+R91bGhwRDmSB4tYGfXQVZAoi2INfWhfb1AwP03w8Fi2efZapEe/daqgS14y51+/VJkcsXe
Jw1jooxK2/HDZeZ53KGz3+xCJutnIhlhYe4Ulh6e0n98C5T230oPHcaNamHvIfX7YbU+7M0AHnqM
Qk5vjgYCuuAYxv9Kmb3ZlsPn0KGIJMZweaho9QSeLqWqP6qeSNHgHbZFG3OJ8/oVbbrpbH9OJB3X
5U+zKGZXvy84iNrhCXwxCRntoRFVjCecpxIBJCWZoUqnLt8nJKwhF2PmmNrG1IsWtt8jKAPblYqC
S9NlN4b57GDoHG3AGG2+bvkazP2owNg1NCXslcpG5OXX3xtM9J3nj5MKVGZykYCa9FluHdmFRTaa
WN9SvGXkVX9i8NIjWL2L/0usUqqWfS8gzX8xu/YawaY6cMkGG5ZF3G2KMPlWwiNwEGbUjO40dESG
5qjzL8pNtWqXlTYZVHDJ3d4hNARMQscGksGulngh8NzY6Vy3ZEtX+trSELtJrc+M8r444S1GNzjf
A73253um6KM3qyS6KDUdhWDfT1L9uY112oxxnqLq0y9rIS+fdLmopjrFOg22q5SLxE8Y+Zy3mgls
gFQ4UI6g6hU1AWYJQdG6sRCz94nw0QPoBADhsxTTnofx43cQimAcdXLGwMjcJ4ix29MD8Id092IU
mjwUAt3piycpfRUJMwgaQp0yzHZeOIHAqURWOO8sBT2dTQpoyO2khygJ0Mq1Ckz9g8kvOm6eKyRW
90Xmoc1VEAn4W4F76PKnBGtSGOQ6EJrxoVMY9Zb8XO1Jxdl25rmppsxi4M51qKtIZzTHoXIuxpHW
jthoCZF7uL2zOTpxaV8vXwZ/GmYzZkpJrd1KGCe2wT78EMp+eWO3Pp1cdBKUr1Z68T8ceu8pPKm5
HJCmJ2iw7nwBlD/9x4DztQVM71mCLmotd+uBEn2Mwb6SewlEwKkYOxlXv7HIp6VgwLh23Hv1fh3J
k51LudP9U9XHvwceI2863zBBTnU5yRWcdA4RxCbTDBjqU8dg2SDTu/F4iv7pXEYKGFjfujIlM4pf
ZfS8l8XE+253+Fq1A1UFehes3RyV4+jLCCUpG4XrBnCz0N63a4tp/LRZIU0JshyJ3mL8q4hMW87x
QaI0XqaTjABie7tz2OUAeGOyL+xX5wkUtCU3nXFa4CY3y5pW50WkziKJBuUNdWEQohz/pNLDXnbK
OuMW+e0lS3QACq2j/aFJ/08TpADNzYVdda5D5nCHWVjmXRARVK/O1pn6YL3GAi/g7j2GsGb2euLr
RyLerQDMb1YnrGmDjw7yT0D2m6e8JQtdSp3TTob3Xc0OTE4fxItHP02IRt/eyAdpLxg1Dh/LnyXW
7aBv0uBb+FUE2qCZ+tNJkdzPItc978ANKWH8O0DX/t3aSRz1ph/NUaP3oXOJfF1DFISuzB/Q1cpi
MQ9N69T6s1KdZiBu6Be2SI+Y5PoF9Wwr2mDP+fztJ8QehuuASw6L3qXdr22MMmNMiLcb28F00a99
87sCxF3+UjPgVjKbrGtdD3dbEBcXCp5Spx2qChbcSStlAQ9HOUnIs7ukD3paUdgD62AqUQ/lPu11
OqDuOHTHL/PeTdRVzqcLQVTGq3xCzfkta6sntM8uUrMDKA2Tldu6klg3wgCSgtpBS9a6TqGz/LiE
9yLMQFHd5Nlf4rBWX5iqfebSz5T4vI0JUQeThVDmtLPlBAUg1AMqWhmuex7mvba4VohXkvThrpZL
A3GSo30WHSlciyf+paHPme77mjYSPs6YmYwmpr4Kf5lOrZerPE0xJXWJnNFNJreLzqu0oVAEkrkm
7pR6pP9KCGYb4EupqUeepzK0+Mqza+ONA+aWk69ooLwr+Wo3uJ8mGyQzbvSN8S4sl/3b9PXgadH4
f04gQ/MbkIxgZo4rsi2Vovugmd1dpDiOTnw5ZvZhrHoLiQbRN7f5uLORK96KXRVKcIefm1gXFZsO
xitBoGpTmGKgLNXunU1TT3zdK7qDTtednkAn+kdmsN6bDw21QCLaQGbovwPrVT5H90WvA6JSuzJe
UxyEkVxk8blVbU9jx8Q8SjgaFlvoP2z/g2pDlq8lDGu+Ai8lXZD46i0+Pkh3TCIwz1KRhNiFrKtu
5tKOlymVM7qPDZBvDgZxx9OhLuAPjPUHI258jJICPvY72kv6fEpKYhlkp1QOc9ytsIY0EoNy2P28
JoDc8855ygPSsJt4vaBGOBkR6XUlLaEEwPm9EscP4nNOALqORJNFTRQK+RehxwbMRJgbwollWIxu
pNbg3hOUGewwdG5Dq96J7HG16TYMmHr8Ho1oWYEQwAK+42Fzj51Vg98ZCw5aPv6DHjlciCW2DhTq
Ec/S0TfARnCFxYW6Lm+swgWjU02VoYHA5VcrSs2Kh3P+tNzJLECXrpz0lK7nXlluLNXoAOxLdsZ2
3zTuw1Kw3PuwtVHj/CtJK8hDjMpx5dIfSZaI364/pfHJxhW6p8b31+EqHiIL8EXL7MfTnE7JdIL0
sj0P9HGUgCt05lduwzmTd8Lw03v2DiuRSBlBpSfcZswASp84uSH8wOe2/5MwhHZAqpa2UEd+QxGo
bGTBFXmBi7fnKYV3FYuT92IyXyeB+/9b+z48+So/tIw3752tuX8xEasQ26X3LefdX7GxkyTwSqnk
FuTMZ3e0Ibxut0AB7LpR6CNrQl2rAU1eJlPug+l+eo+1zTJBpPZ/Hwu4BCR8WsQpFu2EUzYSJM14
/ujNvcZpkQynlGxFPKHulHZPFbRW8nXeOCjZAQy1MJ+gGvCCoXLgQuzSnpvHH4sCKkMiPei3k2C+
CEC+IugT8Rcm9FouGNah3K8dTUxNIq68KA1WJH0Nybior2uTecQ05CH8F/JQpVgGEZPNfjnhQVxK
8ugfDITJ6q5V2bVe0ki7dyGubkE57o+no8/2y1hVvqyKKyzshNny4CF8LueiICLSZemNPJqKP0nl
wuEH0YFc8u6n/M2qgu4Yk+725beQ15XtrT33bh2TWy0KskWfsuwHPYDQ7fcYV1kIO9Zrp0dFBoTP
4l7HgXOcz+uzNjYPDKlUmJ5GzYwOf/wjsgchYdbShV6skAtJYPP8pfDj0/3Mvo79oGjK+alGru0p
z8RQg83CE1zyLV+o37lzqZ9b6bouZ7T5qQZUmHFisY0VUOFP70Hks+zAJfiL/nTng0WbmatyzTkr
oxU6NknYvJkjeI71cKkCT8M8f+kgikDEQpvV6RXl9RQFraMuC8I0RFkgxculjtE77W418Ve50Lc3
kCvZTJKFp98ek77ijR7mYDvpi2RGKjxzpC2ECNO20uw6nUwKyLRZP9NqsH51y01l85UdRQWuQ2P7
u9uU9M+QUzvTSYiCcrUPZO6isOg3OmT9xEga3DHYxcuMcDWqUHL1GeavmMY0wbhjlOP05hsNVQ8g
s13wP+qCOTMPhdbmHE6hPBBHZ5VaV0rw+/3ae9521wDgCr5altZJ171b6ocEQRcFIcJ5JZY7lLY6
9FwC29cjjH9vysQOaFHs3FV5FPYw/XX4/Y7VXBaB8F1SOkFKpAozezgs7HUQK0FyS9MjK7tQjpBR
zO+kcSEu3omFFjPYXex0BDxikuPGoBOJG19I+ntn43/JnU8Qx8S2II+EDGCD2pX5csL+4LC8XUw5
ZahhvZFabmE/cnS7jIlTtmIWfQalcMiqoJvH8/bm6/dfM+4+b+lMRBl9veFSMmtEcQ6NAEq/Zskl
URqp60ZjZvLSiPt3n3Q+9RBHQMsgCGARSSDBz8LTUENiRNd3Tu2cJ9LG+JKWloHlHJM6hahP5DQG
syb02i6amZ9gT5H4945qMDjkxmwkeIpIr02tpbiUagFyoWUhsrI8mOn86l+1R5Lte2rZIX9gn7PN
Z/nwpw2H+hzPFp5aGQRtkAgigACZmefTTVJxocJUCmmcVgi7ritk5mtbM/KejBfJr2F0IIE6F8q/
hyCCodyxa4Hc9fNXvKM0qCfVyBhyBy47kL63wQbygNoO8ntG9n0hNNTjgpLgRMOW8QvafrC+W2sm
9JEx7MXJQ6dJ84XlBjKodKjtq0GYGtqHil4341uKE0LKvHIFho5sbQYthHG/W04sYyP2bpGeRyJG
DA7FBDQ45MoPMoIeDpuZoJ4speVjPEwS/xeCIDTwfkkitF8ZY52bXwQ7mGWPs1BFmmO2F5IgAolt
qRv0KAwaFu82/3aM8n6cLljkXM688soVVnqXiXP5QGIdQ4d4Z3nbcpMEMQpulZ4t/uqngWyW0D/Y
IIlyS6GMTkPJNGEr9Wm4gOR7+DYw4NU56Nlg7ihozT25lWfCDAVvrMOGgNH2bLuswFwuC2zT3SUq
dC+L4jn4G/1AiDdZWUFc3AXx0Gu7/kJ5E+n5LyXRFi88TsgB7i64Clrr9qv7OxLapuhd24PQFvXh
ft4b22AnkzMuUkgLf5mdEbfLkxZU7uUGmmFdrTXAh3e9+4pMPfdQhhi2LS8X32ZQBaorirD+2CNZ
QWp1Ej3cB6vl13qHV2cfGsY9ctY/1O5NQkZST7emFbGD+8eupIL4fXTVhjsf458CdDpAmcX9LhG/
K/PM5BE1dloByKQ+805iFMOkUjNxt9zIQOxzEwJlO3Hsi7xLcx0ZbQQb2dk6rQvR761PjBDpuJOK
aAtFJIuXV086ZI2xMVSn/wXQKydeTLPBpMcVBeabzU/hNv+fcFvCqwQYEnbhoJqGRJYx7iXwC4uz
dXdiUQRwBl+7TsmZcWoFn6VsRtKIKxLElKdZ4ZivRNC/SAj2NIC43LpBsPWEvF3omgdw7UZ2tbN0
JM04Zk2CRKwOtR5ggT3LgbqKZYGY6IeydmZtMm2Tb2YphQCdyuef9oXju20EWGOGHBQ1QY/vK2QU
bUYz7uZeOwKP1fsy+afiICmiHEk4elnltRGDNgTwfLXbJlAS5AeYVIGrDQUiljTj522atHgE0S9v
Li7d6Sdi+7BdWuo0g+ArLt7ZMSo3Ocb+actaTXNvPpsiJMTz5zdqUo+pTBlzFXXmSLM/odIDMMdx
J80m0CgHqugUtc2jqQnTyioUwtiFT3LODVvA1jtJNOlq9MP3BwtnyGnVIlneJphljDRmd/YWcAjU
5cpU0W+M7MYNDMuKy0KgwHevovruEwwpDndOij63kra1SwdikmPuv8q+n3+UgJLk4K3Fsg7vXvyc
ZVdFmW44EUoK8myyRoGyDgZxrjAKJ9Fh7GVaU1FDNGKqeG48kP7FZpGxjwTyR8TT2+lrKwzmwink
o7iXaOvJILIESmCGO02Rm5qMp+G1JOXWI//wPY1FdtxIXd36Ueir4EhRhqM2A6PpSn/llM57eoeD
K9eJ7hkN4Abt58qQo8d3xfLgcNQ+ivz2S4wLb22pYkNVmRFzs4JPRiaoVOSuM6idfDg3076bx7py
3ftPk4P2hVQp9E9Wk1dwnIM/imKwhmWCoLY4dZtu3oqWvzoKJdYhOit6PANNMc56hQ4Aw62eb8On
JIyZjShCg5p1ZVWlg6ZaKpf5AkXBO3oMZc1SsE8j5lckHIsSnWxBieAkHpiq/aQqyf+gl7PI0qsQ
hywlpm9F3ER+iPqUvRF2/qN5wMzACz0Ti4AIiYcsv+GECnHk7Neo0wDWfiMCLXRYY2jqfbJf3cqX
r67OU1/INEczpE8C1dWmnN31JtEQbGDGNAMqncykyl0Y88PQ/Qi4OZlOZSZrkvr40bekKl4mXTte
PHLGIToOg71SP4DfflvL/ZugXIgMjywe5NH4YeQd6boqBe2u0UPkvsAR6mY+XvTgEm4650mXtue4
ozDH3uKIB+9Agd/JxNbVjcGRteRIT7CNo5l55fuHmKuzzSccfT6taJ8BDNij+OfN5/XxfaX06VBa
gfpakaBjfVqgyOuZbwLahv+VQic1WhtjGuYIgi6ohcrd+TBCVm4t/1UGI7G7n6R6RGfcOCXAwlOO
3uWu16kTOV47gvz13dy4RM8HAMv3XYaPqY4u6U6RnZg1agiMbLOJxfe9u3KNR/M1NzRGNOvRIhYH
JuZz7WJfHmpYUJJCSE9kxt+jZlvKju+3W0qQrrkCuT4CYc0b8SfadwBZ2f4gCLcjZ6exkwtKWa/k
y7/UMe5IfeuNa/S8MBTALD2J6Kt2RMxmySWDCkvmQ6rum+yM8W6nrKbff7nOf/lh0wE5AOinJCYi
bRGDqQABP/BWU4AucEQiBluI5U0x3HwTQ7zkf6dZ1kjkLE1oAilQqro/R+RlcEt/5kczqOhzYHhD
Y9q2UVQZrDr69zASSWepl6PVLtlTUgYV+HDU7KRfD5gMwJCDqkhh7nmD/jBTFuTWSH8bMmSNbdvp
W97Uu2dSqN9E/N12/XEnX7TlU45IcmBx1lm1qyqbRHoFokj7TToFrJeRQEtwS515WcW520/JqcFq
g13yh07/NR/fU04enRmvvwesg02awoFqUNIPg6n7j/ZhLB54t1mTv8LouU9jWK4W7fJDlwvP9c98
6ir7JOB19AcFhF0HRKaGz9GgUdG1jqcAkqHLvi2Pj/lQVwp/WyYtcVE2Vmm2fC0RGXBgmcgx51CT
HAb4VzWvMXnAeWnJuT3LRj4i5vxi1ljsJ/VQXQ/mx8RVIeC9Gkt5Skbb88O8i9gHYQhcfEHvxuK2
6p39M4o/nMF3leT4dtANb7GvybcDjZw4jvLrwiKbraL1vctPzok7oUgmnodh5XWsmqAH8iy+q8pB
ksZJ3IhfY19x2mx9NNTt7sN8e0Eb223Nofpqzqk+ppH8ysg1XjNo1VyLr5+bi51u3wdPYyVpF1Cs
D2z8uB4Ti6mnnNSo+tS0giyX+lJMpPesIxTroiYM6nmAZ60fqPtI2CqiGgBBjij7PY2qeNYIX2Ok
3YLkSeJr4PHf+/Ss6BiuSt8jMxmh+JAfVGgHBaPfW6mQLqOCRvQoJxb8esoJ0hDBp2Hga4JVrnAS
7OpkpitGpktWiuq0hiNaJmGmli7DaSEzk1QVkj+iLEY2CiWEqsoCVuA7MTpuSsd+c3CjqyLMJfHn
OJY2D1lIIoJync4lR3VUDriTzrmdj6gWHVS/MvbrDmChsn5FjkrmgNDjvPckSQaGLuFmCgibuxod
vzlTytOQ14poVk0H6RzGr6e35/oV+CARqLhUE3hwX5EwmHpS08ADjCZPYYYB+ULcDY6zuhng0fUU
4jCzs5fpX/k0ab1Ny85/0PTVnD06/2q3RLX61vTusdbtGJyPOR63NB/nDQHH6w89AV+CVkNmpPML
GbVOoHHVWIF9jAYlTYQ91Z7ySEXu39CstO8Y4j20+JMI7LSnw3A1lWR6mKoxH9HdlzYhebtShy6c
lqCqJskWxWVc+TOp6N1xPCJcMSWKZJBtcdVDXZIwB18tXBNm4cZgj8O9YIm2iPerbyS3oLL+cRum
X77ufb1U2ayUdhvWtUVgYO2zvaq3lLs9QkSXdmubmdrNHX8wW0HZiDQ6kfNx1TmloOllevibg0Md
C20c/XFNaR7a7G6J0A8JiAp5TWfK47AarScGpr91fvBAVg15r+NQSVF+Mj3Upb0syjasBje3Uv9s
P6Sz2aUlcC0CtcprNAF+izafZ6DYWJgJkp92haO11CIvaJ8X56NOJftzn8xjzWVdGNxi06wN6LSU
cS5cXIgGrgkPxaU+B08kj8zg4msMvZcGvCV40JgUVI8ozAJjcZ5+Sf0IUiP0yykxJ9e8xVckk+kq
EA7lLk5nDjmSnW70ToRgIXzRH7iXHxZSaPE7Sf/khS1T0szS0ZI0kT3Es9K8bvJMOxEnd0e2G/P6
FRbehRsrYkZTO8RX0Sy/XdYRHiGJyXncXhLGNSLowxMziH3WkfF/azDMzDIPCvZ3IIGDKRkgT+A/
2wMsAQyJCIUcukrC1af4g6TDbRijtcg2PvRMAD4/XdpPYu/m52ppH0Swykci1lCL0R7CL8+dZlwR
JbVkdEnEmIqdxu/RfWJ95qCW3K199ct2h/8FzLqPcbb7krIhsoobTNDeFW97a+K7/nIvddL70Egi
/UiLF7eaC+lAfFdcKMdy/SnpAy5Vm1OD8ZYoGZsHY+ufA8OvTmu9pa8PTGOuspyQucYAFaUx/jCT
8wiZSEOq2FlbBD3P0mTxylw1yg2zAVe4tDo2TWN/ZQPN75qT9AnGuqatvmmpdKfzzNUI/2yTzTIV
1n+Q0fJZylSzFRTnHC5qaJCDyfuy9ernHCS1RPCC6Q/A6qJ7ftk8/BB5EZKQGaJ/U2S/050YxIGJ
B2bbzfBlKW2GtWqUEI+T6oYTlVOHw2Onr6NJCeiKrLQQXXkn8jMh8hogZ38WC88Ds8EdcbOU0ru0
bh44F8Y9yaUoARJ0rn38psJ1r3yNh0Zy1ctGa51joMCbZ0OpN4xbU/9XlyVTsJ5sazsG/2PEsNJm
oD+93+dOW+CjqWrBn6nwFuyLwBdTb01obgS2f7srDk/UinvmqAKzWXwOeI4xHpRI9ibZSp81SyC8
naScMORYhRuA2Y84HP6JN6RHHTIIUdsHZ2wz0zoLlUEqc1n4ZT/bL7kqlH2aLm6r5TUPcZSd0FD7
g1egEe88AaZZiZPMTrzsqJe3jQkoQyN2Oi+y11JGm6JKcChYaFSqwtuy8MyzK7UpscwExXiJwQTi
LTM/ABPDEAP2srNyrcnf2WU32oP44Eg1D+W+vj8Mig+CguIDRhoZAOhmBikigPVrXGoBzPcdDS/l
TKxEwFu2jTKD1/NWGhpa5mxjy6NfJCPxbqgwNBkd+I8W15cwwa6MEbQG7p5v0zi634HdcKgBouXZ
ku31sYouystvuXJdzwiiGIgdX94q7KzeYzH/HHlenWAVirI7qxDV1UyimYQ4D772rvsUPTPDBmF4
7R5OKA6JELH/6PoKw2KATAoP+sh/lW6Zj4H4+e9RUXu6H66OXr0Kk/FO9RIGkY12hBvCmqpTzwBr
CACwwIjGokvPBsbc5xlmxPmXTWDrB6WJNZv1DnpH+aCLAnQRcMQu0nIad4CrEqvKckau2AKpJibK
yZRw/GXBxQ3TWRtOb49UXVZ08liIjpbB0ysEgADcrYYFQJ4Ho0I8jWLOMolg+J1jQsOJ3WmUpuIq
7Hl+UgCPNGDkC3gkql+hobPla4894CJx+dJErM/Gz/A615CkCBF0ubC4ExFeeRW9druaksv7apnU
WKlhldCdzvChLnO51UUG8QzRSRLHj4Y+Kz23uYf/m84Bl4OdlvF1yiRBluQZWV2tvEZJr/wyv2oB
IeRPMQglrcsAE0qyBd3GkBOtdQpTc8Z8/jAkbi3sXlRQlH2WfIeNeD4wxK+0f8EtVA6H5a1x0lfX
V44XdFklcfQDEKck2BAkp5XtNnGZUION6GydOBXwqRuOxlKzCNtkyvPXIwCLTA+H/PBh9bfIQ27B
AxYkWRCyxnH7VSh2qw65MOQYSKdz6dfsBCmJEd8BtMNZYPYxjmKiycjOpG8xPsCMlfVz7tm2w16R
rVikxdUx1B2KadtEC1vxJuERXsnoT7bgBOcpvew51dpEeHY+0Nd9+xx4h2m9h0D1e4GTPd9tCLV2
6AkhEpVaLcuF4rZao0zdewKVYKmd6XSx8l5d+/89gixPO7AK0NQmifXdzUHHzasHhYaJEcMGsoqJ
SNdKT1VA+lxDiNsYAkAmifsOIaAS6F6FGKr9Y5mbZBWJ1eBhkhB9tHeL+oqQWWMD/+hmR6WZ9f6Z
gaiyaiOeSAPTjtb8Wy+OENVO1dq8QzScmaUuM23gK1bvTw3IWf5V3l0ia1T7dKubcS7dGBv0nMI4
upKt8VZwH8+IcNHHirWwYvPm6P9bn1+f+Y3S0tTNqHRld4qd7G8fBXnCO58UMrL7VIqP3mPIP+9+
SmBuTOAmR8dtdBW4lkY+w8Ia0Ll3WoII5Cs5dp9QuZYg7vmlj0DS/oBXKjbAxHaBv41VQDQ9tjsc
q+iQGqffoACOiQ8VsnnqV3Y6BTYCOogblfnHuADGuCQUh/TPlbOTSqrIMShgevNleak1aWpGnScj
UfTXFdAmL/hLomtzgmT4rV/J7yvVdfSRwVleH2Lz9NGzt2jsB8gNtxJpFLrbWDv3HJvMC3h6vQJG
GOFyNa838GdrPF1pbk0FnqtyIp9c/KXxrQkRh4cstuF6kBVmQqxBRRBnymy2vx8VKIO0JH1dgdU5
eaBOF+ZxWXYq721jwJfABH3xTfK7vILidKQ2dNU9JwtfLtDHG1aadq7EWMWT8Bap6q9+gSFfHcvQ
acs1R7GOz2woU6vLkpdyuRRYy8bPB5cFnFjSkP9OWaXsBi3YvCRMYX2jQeHOfkjYi+Ex1DPPFaPB
Qyh3baXXeLmbJ0UmsD1u3UXJXt7K8JOcavv92iGGcIwn00YOm5e5fWJOO79YJGBJZy2ICA0uF6ia
IZ6k3rslhyouHOKN5SbZDuTSHkCqQPWNAamoMXlFQsb60BUok4r2rxOOX4yl9mWg1M5eX9Mk1enq
ZYEXQHk6+pYZfEuilFefWgblHUOopCWerWCmtbZs5zhMn5sV1ML7StpKYYjvRbW7iCpA43F+ITPo
9XCAiXWIgW7E9+n9BPIlTKJw4t+htOdjX5rZXi1eksZqD7UBHMQUypHhj1+BwdwDTrQhE5gdTMCN
TzI9PI15Uie3erQz1W8PAxx8Vs7ZSTWsq7AkSbmf5qrgr2Svp2wDEgUr9iXIkXLMYIgo5Re7SnQ3
r1jEquzgfrcAglU4r6XnOlMNQGokcJeEg3KEtIlqwTUGxAIJOoTiOfDq4aOOF4HXfa7ClnrXDSCh
VgFIWJZq+2DoAv+UKOcN3OQA/h/rJW5HK2g6ly3aaY81fih8U4wP8v7ma4Xlfgc+kmFuOB6Agxae
dmz+JjpdpokY9d6TYsuXkfK+zrPxBRnmmC1jBomglXAr6nMFgYd6RIlJF6ub4CJqkIQvrdhbf/0j
0tn5eLI8eY8PZ9TBvHnMNLohwg8+MdVKqGAmB7Fs+xErkyM9HcRxrJT0KKQN2GCPwdpczvWPzQHS
W+vOwRMFYZM40xm57RJQYoVwnM41bMCZq//0isBTJSe/sCZ1JhsZC6BVNDceSGZHSt0Z3lbFA3uS
S4jNkwkgMPLxpIv0T9OZu3xoEnVeGmIBb3hVtN7CdjoYM6VLqmaeqNTlS76qqUCond+lcccXUviH
9cxAP4JsZlt5Agiq5of7GPgcm7f8a+jVMow4cLwX0z5nUQZBD9JR2aI8SRMX8MVTZRogAjInw/4e
JgLgtw/vDPdHaH394jbQYvRopVdQz9XxUGPqYj2cIiv1Jg8HPy7/iqPCL0fIO+mgPeI2jbQrB/sa
7UNmMnwm0Gm75wycLzl84w/f925f2BZQMSap6pZTPvxSgU+4szD04iQZ3HI7e1ntxEbNq1iF+DRz
EZzEG7tKAUjdadKE3uhl2INQj182RavP76GHXuGcknkYofBF7cwbs+COb3O2OvC4GJUbaPkOz7O4
sKCxLTMIMr0ms9djhtdm2OCi11NFGuPYrSLoQZONqISywzz1ZXPaVUF8s/X8LkO2OUCXRa17sB2l
RCb0Lj3uoBgSFl6KJdkI+/6dby8dZpglFX5g+XrNanrtB2nQ5AOa1GQ2BqYbizvdy/qMf9JbQ2Xg
glTEiL5RD/YF9T9bnX8B2yxoGwPaFNMl+Xzz3aXeqf9OzUGWIkaq6zgBC1fjZSJLAS3rWpEH/aS0
eZM46OMnCVKIFlQ30+r3/YeIEnrh3QmxLhOszvW4isCgBDOUr1WALPSEDc7XMm45jMGDce/b59E1
pDyHssE0/IyYHlbjsYSvLPIzYCiui5yN3XS2m0YArzmUJSCRBNOoUl4Mb3ErWqKJYNa14t007MZW
CHsxgWLqsg1giTjx8lK8JkhZB+pykqu3tsd5M30+atvnmaaUFHSfjsOqjmJ4p3QZ9aZPM3bttx5t
re783wj+iEf6Uu8JeXxoi90Sfl1iFNAypkze82ge110n/Whvd72aCNOLhZXgggBsDM23RP6GOpr5
vRSs1RbnLBCmlpuj+ocnmGZHigHGZwgV6FCK3BEELmwRu38drMUXZcBV7BEqwbiwQXF2RZSuwOSL
qoJvvUFWGIK9C4FRCAa876q/GS133XETEA5rfxQDl9IP7ipplHbjglM7SKFFtlspWTY0GzzIt/d3
9Xw2U/VHvpuggmt97l/vHLFQDvdlCMc35PDjVeVH7HgjVPnYr/6VZPHz0U5Di9J4a3f17OMp4rBj
ILTCZhumTswc830OlfDOVlKa6fUhgPO+RZijp213ySHyD87RKsLKlOq7/rbPDIY5Jk5Tjqh7+NYI
nZVWSHJ8b0SwSQbVsOOeyhZToh0GvM2cGC+gosSRwgJPUxAotfHNCe+LSfKpmKwvsWrgePOYBuoM
+daNN4c+BAG7u10xA62XOAWOfoi4MeoW7FytbnBwzglYCGeURpDhGXsWV4ESWNk9Ez9kIhKL6bKo
2JolC6iffrnEanaRoRAPfO6dQaaXz383IpSjNyohIElkkN3HOe0tRRD1Nj/Z1rkBMEJk0hw4oAn5
4rXSojU6QdbLPwIVQXvSlXd5fZlp0Rgf/2P2SqYxPeEpx0K8q2DIHtZdTQr6BZx5voGZ+gKhA+tG
yQ/gkgfFB+AfeWbhBSPXkXMhNUYvgeNoitdXVdLLJPNnMOTlnQZbXo4Aeuiw53Zo6P0yyDEXp6kp
4YmMtG/B/NA0mKeVzBIVpiX/2ZEE2/wzXSjC921oJnZgojvtPHbF0hiM2o38/p1A3yc8nATHFD0j
AyDBz+ikE34uHsF2izDbuHW5Br9UqHwMvnU0fjpgSaltM5JiS52PlOVZp4FwxtaHpcTfCTubRXKt
pM3NB/rFsjAwYwGxxuJYyvVkQ/tYVMda8FeToUUruCHpjCFQRiT2pa0Uz39yK7IHywQQQ5MJ1JhR
7WHI4q4FKKlnvPX6+hjqxJfPm2FBwZzod9TeTY+ZbkBW0EKRJp5lU5wu8TZC0Qv/LQ4rPWJXYQFX
9M4lnk/V9idV5EJzX48E7ItthqC/bTWb/AzpxwBvtLmOW6AWp/CTM/FQGh+qeBBq7hNAskLpRAIU
Xwha19ZXM01ZtEfvv5CsQf3LPUHfGzGqfC4KPx6AXpZX6fjrfUQ5+NGUE3mEXYJ8w9Lj2dw3QJhR
OFuD3eUnSg+LFJhfHFZV7eYSmpdelFNOxjkF0FEif7/OGJ82U0N+x1QOx6NzsQLyNXuJRsBN4g9Z
5iY1HLeR1S3XnnI6xp7p1RkHqOS+XQtpFy4N0XeVFHDZpfkNUl/4JPR8iZGFb97ZsP8h0kxdL48e
Vktqe8SYwGwu3JW2dZceLpYwAkQORApKq4KVjuNIOW3HmmuMhAHOMUgGgoYzNKphlGPp5X72pgOF
gAmJRQ0wI6aaZXOLMR9xgzDimG1IY2Ej7HSdGcu1W8YFnYMPq+HlQLcWknJtYlNwWlkDX0LA5310
CwmTspqaIXGzbLAPS8F/wJVTSVdLeICt74IT41qUtb14eiwWtAj6enaFHEEHgjjJ2yXuKJXCwCIL
9b9k0WNhoSOtV+Pr6VM1T/hdd1HZtdIkjU95LYDUoG3ZPzGpgCOKoj+ZBAnkURU+CmcYelXGdb00
lP6D4REKd9Vbw9f3LXRDXOpOd7vD8p9TyowTloXf4M8HwVCRr5pJO2tskfGsKhAWXJUY/fSl2cIN
2QLcwKOEgq2UXnEVkP/6K6VXcwbbRqGorPzptZzPPrAHZ48OPyBDIs1f5eIF62pzI6bOGZUw7NfF
msf8DmsLJN+uXM3efrKag+5wsv11vlYPBe2idsRCoHNztpAozShS4UaBCTtkcVWoAimdyQq8GIbH
NCw0RnkKrrWX4DI5dWBUTYw9WGLCOo3fxdrnLuLGW8YjFnQOZaHAJVYoddD4+OjspkkBrNI2mv2V
yyTiqaKdTp17tdfoDHmxY0w0bpEEBpN07GEUHohiT9AETokdnBNRyjRATZO3JdLfTounKFJhDI7N
hVXHfoK2680xQbKSfhisseVlDdUvWY5AJND/3Nm42bPGb5nliqIOop+iTtm1IrAMYCzS2N/eZeLc
+qk6h+tU4GU3XTHqVC6DevyNsAf9DV3xu4/M0+/WUgvtDCgEuDOQ01kVAR/vpHhYAhSeWFOmwqAT
QTxyTSLSNKajWQviufKcjV5Bcee/HHSlT+m+gSnJACQTRmC+yrN/OT0jDBf63eHxw+7cXP/ZEGWr
ESjlwX84kgRu5owCcPwfGp1ohUq76Md2Ll6AvT7xKnGVF+BycidaDOEsstVKi7griARmFJ52dbOg
ne5KSjDRylCwHK9JE8+q17pMS1sfgGocmkPB4SxTJRr68GD1tAXzrRG8oxdx1TcBFZpzQpwgYdqC
I8xkgfB9KWChyLmLFPVlPD1y+IydIeKRK8Ldsh9Jh7t4ymYF15yGT2IQj4EyGgDM025uKD9jZ8SD
FiVcwG3KFai/A0CC4MxqIStDZrTKbvqdJV3PNwsjOftc5i3kpvp2TFDl5P4ob6dEtpDRMLR+wTGo
yF1HFyQHTKo8VHmngxVdgIy5Y8S0fSfydjK2y77k1S09ZMgNJWvIg4oPoqP/YuOSnxR2tee5bjuE
9l7AjJAipu1kjkRARUQsvdFmFyhNLHT4Uj20ZxQPeO85Go7faYnx22ce/vkkPhaBnz7Q2fCY8vPi
HdeXRqkHRR+A8z7XDGbHxej6JaBYutmittUAmhYX9yPeA4FawMCeqy/hBLI/EK5u6lz5BwiL1zbv
wXJec+DsxB80kWYfpi4mDHQjstTl3xQvIrCkyn3MZVv64X3GPeICTiGkJpJWpvAYykBm8t2QNkSm
U4/dJF1jUv70MKBlx6hNgXx8fZv6yyuxzGepKat/xejLIc5qyt94e++xQlhSwecBzpNl+zlWpG7r
D7NekVS2pXEzbJQ1WsglNVBwDH0LQTWzxf1KfIrPTmc2l4VHeJ44JtsU2ZTVVlyx3j2PoKllTTAO
0pJv7+upMwZxL6Cf3A9WW6zJrVcfvV0ALSV+UUGHE7U07gA6DKQcosI3/xDG09i7hGaUY8Q152ji
uNNOVx0xcbTzQ9CrjbRk1am/BBKICp3N5Dpw8I5jyFE5qPV82PgQ5nQVikMg+tgm6q4KpIQ5x7YK
a8+PTknWN3etyLvPwWs0NimAwHu6B13m4vJG1vwPtcZ7D1B7ejtnb60PxdC/SakfopWfNOiy2yOM
kQmXNbKH7fAjo+gmh+zcGr/Wv1qg7sMMxZ+vGdKXgjnVlvnCI5UBwhjCPJZsyFJwzB0emlrgIPAY
nGA6wSsOvctBW43N5Gu0jGM80zC8iSlrdyQJFldREtkXreu6Jyay3+U1neCd1Hy/TGCtDW6BKsjL
8al0uY+c5rEdCDjiqlCMsYGdUWFhG5GD1JZL5+c6/rF7W9FHU6UxHNKD64kFJ3WxAeMqJCPh692u
hsoQBIBMP8vUdc09IpspXZe8Ok/SK0vIwudv80JFG7jn4Q1FSMdwyyW1EqcjlCsajLnUp1sMZ0u6
Lhtht9Vi5tA38aay05fsaBa7yE4wgN5UbBmdukyqDYPXDZZWSbVgZzOCZ803AzyCjbWTZyQD4ErJ
aSPwx9nGPLU/fNmGITnnOnsqv+gYRSsLAgizY+tru6d+/pgx6EbeF5AqmQ9xrjuHID3GwCYyPxsA
sJS/o7axVDVAyRbeK5cMIYUJklHD5oDC6vjxY9UVv+bBf020x0CiyhLw4j9f8je3M6TDkSOGQQEG
7QYmN/AuejXMq4PTl3LzJQYVemDuua3APflkUBEEvqd2uxMeZjBoe9y3J5NScUAX7KlvCNmCw2fd
+TRnv8OhkldWs5SZN0UBcd4oKDv3csIzS+BCwIVcQRTX4EOkGuUcJARhtqN81sMPXRCi9nV8wdM4
4eLF9taL8bR61QaL76jgECnxt1hfsTB6YBgil7BAaMXOT/zdpwq/qQGN/U5pr0hbxg/ER1PPc46c
2rLP0MnOb4xiO8jARzKLnmih7eIuTTGN9475a/wUDWiXMWwP3M5YkvtX7E+e2KS3UlgqKGx7CdAv
QQDzGVZEERIsLb/MMnXVlNup5A8/3wRV7ErNLsP4vrxxhxc+ZpZOFd5MDMKpNcTd2RpXmt8DCZKD
rkOgsgqcklQuG5FWYiq4UqpEfWavXZAwyHOOwybqvzheLjJ9ISW2VgCGN6gnyUspTOKIIuhuflnd
rgO1IitaKOAHEgOCR343HnrxedMT9dFXP8oQCCY4oQzhEiaaZ9Bc7BJDcdKnbkTarsO8IkAWPi8A
sFV4mWfb/S67fZ1nHTUFTgUeq9MGEuWJEMp4xA4aOPNuiOv/PVCxAR2WaZddTp1XMw1T532+qM3W
XcBq0993ciJ41lj/CyO8ej5V9jjbafh10y8WcrATY0ohkvX+52sVZ9NyP5Dsagce6/SxERMp09yD
e9hogBdmCu4B8uty2yBl8w8ay5OG1cLeDWtp0sXltqABmi854GVGWwXauam6VXK8gi3tT5qv0/vH
vglk9VLCsuvJLwI+tHfBSjhh8n+8J+OtLajUUSbk1djZ6qDYPBSqon2y7lIjrJTc9qH6Pdw0x5rx
YEbqQ6xEs+xQ4EFkwhZPdp+AsP9Mo1sezGiNtO0FKamFgGKvh/m4wZtKf+59EvRqUd5WPET0+Hfm
I6LHdRVq06ndGlcJYsjRRiJwCWneZfN8PmdTAYrBoom3gwXO1+xS0892YIE+Ia3CakhzUoNjbN0l
7+VyNLcYf6SKTjwMzphSQysEWRCT807RPqbrvHGzIjprgAms0gfiFzuybT71Haa6LO89zzBSMLD+
640BkPtGtRjh4NP++76xOay46IvTbGnZOMDk4ZQLiYHY84q9Vm5uGosC12copiju40UR2P4ZlhxX
JIpcfJB0PhQ33x9Vw2CYhgzZXmUocIHPqz6Sm6aaae1qX/5Z/r7g9P6/XCtxxB02p90iBYFGk3HR
UzVcfLx60OEP7j6R3lDZwKn4ZsdsrL6XETDTK5+W/2SssZp+rSlt798ZwBIaeRVw2/XhaciQCwcv
aj/CdlaGXhWTNzjiyWLDidVTEIMmmsJQmjVLVBFilnvtNbxNcTGRO534FZdJF5Mr6+cuXgRYlOoa
A9r62qCMQ+MvplbN1wqNqOStENifGnWiPtkJDhBnRTIqWMmMQg8R7UrHe23HNijhUrSUeF9ip6AZ
DEA2q3YnOWEBPfG6QsH862kNxq5yRgRuifJtjBdm1CAZGIk/NNf8NdR1ilUJCZMQ33OnQ7npMaI5
Z8js3ijtjTjqkNEIJSv58nChfPYZCBr8ZwrT81htoNUHCyt/KCsTsalCVWcP2GgWknlIja0mdiAa
1l8vu5xGIe5hV2yr4LZuAISAy4Z7Z/XfFQjsB/iYSvyy4fPUUaKwak61S/uNlPOtcOPO2gCTv9iZ
GTwlOVb1xrhrdLA1uDOu5JZwQJCSwycdq9h4Pk0B+X0OtEAhpUVsdvkIhzM1+9X4m0bVGVz9Cym3
fdEW6I11odOJKSG9ajREeGwvAAJFIJePjId1gkkASmf8xrnnnaf9tmEU9QHDTytI4RDj+TT6abch
GDPp3g3UalkWvDPHGpFKy8IARjDT6phiUTxqv2AuVj3l6NNjmAR7VP827biBSND6vRtiROdtsbse
MlHX1eOZCmCeDo92IEcnyvQArKQvjQ0WSnIfyJqADmXal55nxOSUjWcHRe4AXmDtotWpj6ajHKZS
qTUNA4W+E8eO2BYVVsBNb8TRbzOw2NvkO+HGe5AT3KUqNlGKoQzYvuLChIKvyPT5G8cgb3Leag0+
5wkb68X/Z1PHPxUevgbApBuiiCQjoapaAT23pbby3woWG+nZ8zAUrgYew+c/r3IHUTIn0tOl4Ejy
bK7F0fa63r9wGRwJ80jtnZRhuWaSE+2d70UW6Fl4H5W4oMku54pQNJbAlUVAsyzAxSaUkXnO9lp7
/gS+PyvWMtdRj2/fQlfmTjedOeZ+RvpMFVBvUB2VE9M+8DI9lL4ud5MY0YqaL9glSb7nVEce7zCh
UdTAU6gE8usC/Uf/nhZNWWUyo0lZsmrbUC03kxK2kAe4ue0PTgSEPdc4cga9EiT7p3nADa6B0LGZ
bihH2JgtdUFd5VjJkJtZpzVXCcM+xfDeMF6GHRA9PFzPq2bAeUtTxqeSMb5whZgs2d8DYFQvZkmX
Eh1bMwOgsLJMuasbQk9fATuBplywMTsDJYG3Sglw3+q7iD9FAXQIpj3T14ccFToOeMvuaKYH2aoC
ErYHrvQTHM6sT5s3o7CmhtATjcgAakQju+g++4lkuEd7d/Yi8q5KSitoXb8xyq676rCDWuDJgTGr
lpJm7R2xeo7NkDUi+Sce6rRd87tVDcpaAVNRQ94XMwltBsPKcyVA86vD//d7Uj+2v8lhSiJTV6Pc
VFBPl9UrfT3PU/pf3mY+BOxB3DP2aNQuU+rXgfyV91tcTxSNwr2wusPN35wnNK/J1OPZVDbt+KEK
ffx+BEwUNvvEP5RMC/JA6/3NxSCx7Ga+stYiH+yS8i9HUBEaWXqYu50ZbcDCNkayfXiRxxJG0Cbl
DF4KTigefziDiNsuToSnzRHugpv0+NhSfh32JaZxj0zmBzb9okSdsflxDY09/H1mEIHQJI0Hk+GB
YTNwtysFYj0HiQdTT5+sahGwcltbseZNzaxGGVMci1j/c7+ELhCfqeFg8sQ3a3IAHrwQpdhnY8xe
MZUBJEL6Hi9PTnXtiShn/b9V0ayC3Zu0f32D3lFrLUaQQq7cEfY/fgvzBY5z7qQbTLQAueHl5xOC
eSR80b6Hmv6M1+Ugh/cevBsGMLAomzL/cfz2wbMSVgIa4ZKKiuEakwc9sYqV479LXVpDcKmZwC5d
l3a+lQem+EEbYLswxpFTqqJY6ESFYVRueJr7u3CvUO2ZFCnNUMz0F3ZMVJ1FU3O21+9BRaP5IxKS
tWeBeXZoRZkIIzMcI1OdJf5MlLnrNd2esMKMhVsmyyNGQxK+VZPfBeQelPRClXQ91fNYU1+dZKIs
sUtcHxKur4wWwvglVncWqFRZ/BetmYXZKlzkmKNUF351V3WTL/TOb3ngfovwHVRe99YZYSw1UhlH
Iv9Ptd581m7GB7WknUQjFbWozxIH8yEohi25tArgYSCWEJjSS1RXEIdmFkeUaKEaEm/H3HplK3ow
yRDS9Xbd8EKyh2wRo3pAwvjSzBH+/sFMdKMPTAdMArC8rUQofi6K0+xXqQwZZ8yPASCCZ0EynLt7
hLb4MtFbqaV+jlNxFLkwVyhXw9k7vldqQfMJOgyQ8Gtdh2TnX0OKIjv3GM2okN3pfRl47FYlCGpu
LMNq5z3XMyW0LuX2mnw/z0ztQV82bp66N1ER/GcrgP1jkWEgQOYFTldMpBoNXk+LUJnNmCiFMBnU
eSTaIMgMVZ4mX3MXi8eF0m3LebCZLOesgVk4+XMiLH6RXHTnCLrEA4C6eBxXy7kRXL2WwS/C7iS0
3JuZIhpRmdf4xVNZERT0PAqcEI9h4za+Q94k96SvXpOz7jRWALCREcR61AkReYNhcxF7NXg1JVf+
QflF/zXMKgHbXtlGDlaEWfSt0/JM8XXD2m/nP6Cmc5VfbZmZQf9uf1CkTmnVdHZ1LVnlkMCo/9tq
xwIsYIpsh/nJBxm+fhj9IARBsjNZhQcW28yCw8jdPFBQigQB1UGd2GC/TCM3dAqirnlrfkzA7ERo
HEdHuQcxbMGu8RO5ABoJtnuVpv/JMiVsWKUWTzh1SgkPGcmKpyjrRNALJifXWK/VZhPllMTkJ72b
vrJ7FGbJYe7gfA8Nriz8+em+NLHCwg4EHIY/gk7k2NaT3oMBfkWfW2NAQkDVjppsgcI88zbUhfrJ
VqB/5RJsqQ0Gb+8TgnV17fiNzkrQK7W6tM7T2wPbfARTakqzD7FppCJUVFAFT15qqK2Fi2IMlU7K
aC+OcF/0hdZCcCnNMqnrNAsxO/RoKKzg6OKZhruE+kA9HPAHu5fFSkKJvjH+KBVPSz8VZEE/4/GR
5PimsIVA3FvQ45/CSo1vUzp4U+aE38ryAsZs+ChR4Az0+25/JkssDGRIcBWDgnU6CEKT949FrDWv
6kOcRYxc02bpNV0oN+s3s3dnI9cb+uz0EU4WaNQvexEXB+HCTC+gYk5/jIIP2htZNR0jgnDBuwT+
ZTzJft1DaOCMTtb0jKAFpt6ipdxJlOGQ3U7C0QsoVrhPyysWcPjXbA0wKEnpUrAm3byb188A7ef6
Y/ZlG0rEsWq357nfNpUo/VdLCnaNDVYYDx7+sHPk05JfWWqBrldN+bJnmf9JhxZancToATEqDuD9
uvTHq69rGOhWS22uj5nEpnxzhPeCm/KO/4KMoSwBvBaVcpyE+A46OgNZDaI9oFuVFAsZatnPSVDV
l73Cm/OM1AacZ7Ubs8V+FPfjvM5UrIo7+tKtQldBcMWmHqB7oosTc2gAg0j2T2RLfcJD6lkxdMz2
LMbL/OgWhw3RS1vWw5flohQr2ODgSO4gGYe7dM1AIhsW99cG08IQnr6w189yFCoOA12HopzKwdKu
zD638DmZZg5j/qVUtCVw92UMZq+AElAVKzqnecB4oZEfLRxiAtx30y8VI7wiep+rckV9JT8hzvUV
WClOUZmaiw5Wyp31FiRIB38SvqnCG6qfIUlvmmYltHxN+6BNMHazgImTEWb50ONUzlj0cv86cVWE
rrpLUzCx0p0vAwyZw0/IKOVOZj+PdZQjb5a58RSnSxg6q1/01u8ucluNQ5Hwt3Et9kWt4llIE6wu
5HmwnzLh00DnvWodAoG1cKpRsRVCa7qwXd8Oy0ayqgJpE5tgeOpZm/oxvuvxUgVYEy8Wyp0zQaX6
XhsLJ5KfRXTFc1uk3iinTYesqxokJ5P1kxDVr4bJWcCH2uJFzXJyl764JRA9urTFQ5myz2jqGniR
4r2e9p7pVsw5Pazx3fWm8sQhN3K807GGFd3vXz4URLya6HRsfTC/vHKmQk9sSUM5O4eO0s+HTqxa
z39z4SvjI761GjHPW29rVXAqKuhF+TdteMGbdQrS+K7dJRJv6wJXuijZRFN0N9keoCjXM5zK/bGf
+jN3PWxZi2zQaaGClhf/WW3wkvJ7z0Sc3HHj/go2/yrl5dxaahz9I8nrartlxQifVh1AnfbpFg1I
LnoNFFNM3vmUr8Vir133dzIN2MYniSn10RfyxJD7pBEw+3wj32UtX7YeZfKKnZdqCWgvJw/5/Nlf
mnUv90H2NLHejMHQs6PCZo+oXJj2WC/wGfuPZx8RN3hTvyK0+s6adc5utRJdgNg9WaaUr3qTcCaG
fCDsx0HKMPml45BENj9Gr9I56MTZK840S6irdql+lfGhR34Ee4WnCeHi+0RLRA6Uoip9d2V4iRDv
kSuYySo8ZNWNBAM1p7N/yeZJAqFvfQfukm5V4YEV9W58YXWESoeZ1TcoYYfaHdE9YILdItE4YhYo
wZF5Aw4nK547ha/W7vffUbCke/smZGx7WQUNmxI/PXntP4HhF+P7vqfCqhSrNRP/yD7jwqPyosix
z4A2WUOLyJhFHOmvF/9VBJgV0af/fLWH9U/AeHeCuUrSnkeK3h/E2wgr7EGjRfxAv0M89o+xl/94
9Ynixg0/yMbD46JrjSTqvqB7vJtmmvcQ8VeEvUfLekM0po1SdxW2ek6sn1e3XvIwwG00RdrcQiij
JzR9eHtlHtAhYTXGWtBHRxPmizJlUw5Dyw9EGbkxAPGjMyustFTM0yUM7z124Ld4MWLPf271hqrs
Y5OF8k5AFhYZOsoOAQe2Me7VhrAdTTE7UjwDjeuV6K1/dOSdKAzEBib9V0pG9nSHo0+vJfUGkgVR
FwnBUg4NQzvAEabN3j98GQz+DfRS4TgWc1ZCalufj1Fr9mUkvkKZUtLffZz50CXfefHBjwqztjcQ
Zk9UWMXHuj2KOM7g6TAaDwkHA3fN7LfanPR85kv7vvNTWX6VyrGaV+qon5Zerz8RcmmGw1coy/0q
2foaS8YHnx8hA/ZSLkqIRLYhsrBqD3Z9OZ11rwgqGnFEaTrQjSdbWn8Sb+SnTBRwbX0OFScrX0O5
QthLTgP/zkH82IBW4KWqhtj6BEOyVTQ66IXRgO0s2rD/VKCi7GvHnYFOyfTJAjorUIZSGx5qbUUv
DC+fZWAcM6At7uepHzVM6XtTY+K3Vi6cS3eaOwhTIa0QvUk3AW66fkEkl02r0vnMe8nFDaBQvJeE
h6Klm39U+fC7rRpDtLlcSFpCDUVbCM368Fv0Z1ix7wNGkMyM8Zn1yuJSsRZvQ4r04TEAco/59Z0j
PKV4UgEnpeO7qKFGSK+kVA1lvyN0KqgavivmRHQoIORZNb4oexwVZncdQwTuwPtWvUAwIKKHpYGJ
5ft0fr10ku7cEaUyDoA6YQUS6cG+5EPDtPxiRmMiXZkcg5mIwUBRX6zUnEEtCAqCeNV3FtRWXo+9
dDVV4++LLKisz828niXLYZ6PLMjXHe72yvl2HGE1aW950racJP74rkMKcm3CZ7Tz3RUgD8s0s0PD
obzs5CVDR/5zzEiWA5JVM7QZ0VbAyizDiwNevrCXubpnWQGwYHRP+cg/r3oDH9I7vKLgqrdIsNfB
xhz7c/qQN9SsF1hZV9BwiHrMzlMSSVQSAmpclZsV2n3Au0DzhFvG4KfROBpvKExe+aJJ4C0dDQXe
aWEOl7QBe6MJBz67RlFTabEXcmTEX2Rs5ob9M7/C/Dz4uoUyraRe6kiXwxbw0MjvJthN50i12Rho
ADjIMVEaZSZLUaKDolrBnFbq2yl3LVKPhbopOQ/POFgUC9j+uHKg6X2Yw0j2hghaFILBCwCyfLOf
pUP+h1ql8KGrBT2MOfduFNlZXwP/I+fxMbyPg2IQICuB5zq6lQV2vcEoS+SvavcrfLLW82UmgzcC
jTdDFHqYK2Cny03tKo8vFcSOJP7jYVNfF7w8MTeNHpofsXYXLu9+IxUiqTuz4nxuRIEyeUQIbyz8
r8wEbHYR5nJVHJQbENO2whmzUFKkRWnJDU7/ANJ5YNVGwpXeBLZ1/wt+shVPFTICWpjeThO3A85i
tBzR6Y1jzgKQp6AFuAPJxHGnBqgsVczC+8VZsh+ONL2GNRjzL/dv5RpQ/V5pizpeTgbqqm7MvFDy
U/W9AIkY//eX1ECj2K+jWJ488v2FqoFvXdcXL/8QFHI+p6ytijO9Zph9GQskERUpJk+lQIonOV7k
MWmSxBGVuYS0yoB5Izbyy2WwtbchD9hHCON47YnptXQ5Ml+NsKfmPMV2Txy2Jdzty8Jcb1xyUOi5
YOo6A+y5XuQpiFWuhkOhsAKQapexBNgUOJu6LRmc8JYeMCeQs/fZGh0Lq4ahZmC5GzhBQ8nvOFVM
0Uo6CFZJejqDTbGr6zWAZOjN/KLQecb64aeOp46M53bbUeoBqU7Jc3rjBU0G4C3nUhkvtsoLrp6z
ZQeFkP0Wq4FU0AZOieXiDIcpS8c9OKjPguQxCAn2IwiMxc4bHP8VN0JbNxaNhxl1Y2N/2ZV4lqDQ
ZcByOybUlm3rI4duW+IPy+nXgPOn7W/GijuFd5AC0RGb4JJ64ljlIOnq6EdtJD6su5j9af0U7aUl
xDStwwgyqY0StGTISiYgqOAoBPQ/VNcZYv02P5pNtRmp0I/FFs26goHfa0oe5VRFSMjxxVhVT0g6
AVHdYGuYorsWywDKyi16CtiTW9yAam+8NVUcMGmSyN8TLEcOsm4LyU3lP/PYh7Y5ZbgZfNTc1d7I
zUFXvZF99Q59onzjglfxZ9nOQMElBjlCyuOGbb42OBgYjW0ku+cMVtwUlKNgRsP3KuMBPgDly/CM
gyf6JVAIyFcQHIWVjPw3QWQAYRZ9ja2JjJ797cG5/k71lJbuGQe2WIvUC2XlBkSTIThu+XvNhReT
LjayuiFNECNJst4r8Djk7xv0nAMmSjq0l8yLL7l5E5RPMKJqF9AqEyDdDI9KZGp+vVHWjA6Kq5/b
raabHArywaWa0cKmpvlLyETtWAFsiCAk3dBOZGa8o1LGAsvvpvcxJb1Gat7QOVfg/VbyIGRz9CDO
z2nOSA31TBFGwhHAbUsSDojQA0IYS5VNHXkesESeBn3h9zqLLGFToJIsgeqET6PISloqHvZ8lYE5
SfaUKg99WYe+A8EmkgbhUjY3x0PY1p6dN+M/V+Ruug+JEwMUr6U55319hTbIrKsRzfvEm5WfHpkj
/3YQibeT38n+C39ZJD/naD7sqACHm+p6RkTZSdxeVywlbwy64pS9PvxB2/MX/RKDt5CCpYJduZ1N
Q0kzCIBmsLFVRLNlNxXtbZ2Zf7LAhsC+6UAkutUDFPxFtymp6aNDjFJd7nsAli9J1x9vZWvJUbbv
gYT6+TU4vsZoJlpIkQUEDcKeq561aG3N28eLPy3s3rwR34KXma0CndaIhIED42DM3JurI9rVkN0d
I+x58FHID5JoRZTF/WHyDYS3/L9ziN8xN5Dj2rXCpOu/XC48SfPC0819MAQG+JdC5fFLoAcrpD6Z
L5OneDUmcmfs4WuodThiHjIQRGLEO2K6makhaa5wX7K+aicRbRaS8BQ3yFL+Uyy09A+hB/5YHuir
mveMeHvLivEvMRsKt0XMexhKXPsd0gGkj6UJCjhiA9V+/copA4fQWK4LVIAuRoZp6cKGrtWL3CH5
0TRCiVfh3vIv5wXuXylfwZJH9o/onNTsIHBlWCZJxlXs09RW0Avz0VbcYZP55Qb0igMTPGIkxjVG
S4AuApuMvfVqqTlY1JaFMsnFdx8O/oTwGmPhtnEfNZEjDfqoWjT8AzMHkwT3Cun5At3uEJeHl7Lj
yQ6OTqbAwl31oZKC+CJYL49CyTD59ORWX4nweNFjzXISDORqHKsfJOAjD7hXrrKZE8/WDlJlF845
N2VGJD+STVBkAWF4seQFSDIx/mNDgYAIswJum5VMByrQyWkmTQAVbsMhyqNzz7fquppkJXTkLkxT
G1yWGKQe3BdHhGSbz6XyWDJPz5N7Qfb/3JrYOgGYH+hDH6rftHEqgsJaRa/bbrefYlIkv4CkjvSg
IUbbB9Hfz9cPSan52V5EpCgXXYYissBbn6X5bnUqAcccQnFpd4Z32amdYFg1BsUTHCTAgPYkKTwS
pxvk8rdhOSB5vHSBkC2GNscb1RsBkHGpuAcsKPfOYHXDn9NueFF3O7vPuKHXmFexebMpW3MKMSPd
tsoK3mIqYV0n/tt+KGfsD6x/QgGKf0fTSpCXj1Al3bTVonNlp4Kj7RNRp4GMkMABHJjcW75/0Noc
zJGUtpjBtJmvFqjLqYxllSjcnr0UN5UuXIPYvswn+lzcokgE2NSLa2hLBuobhPd/njOM+D3/tHW8
oglPzIQLP+JDA60HD3zRxbS1Zr8ueGYTviVDip3WMcBLgcSQ1mGcR+FkBY0POHdBP+Wy4V5zB7DK
jtcukM2HR11RFJl9L2aJNEXzp33J1npYxEPmqrkQeHSKUzJQa6PeGYd/xgMjc5ECacORCKUqmPLK
ma4WnGBEgQgt92V7sbWCogjbRToXXNCQFuG9tlK9gY7BuJdvNez8UXJfGhVeU9ZG7Pqikiuan9r5
rs+XADbt1AcHtgVt8WjKtt5KpeEDavd3ZMjGm0oZAHjZp9fwwxWmqag17vL/sKJ/ZPJ5SyYw/O+m
F9Jkj+qGi1uFvWWurn0N+k2cpdUo4u6J0kXH88B2XmM3xUhOt6Rtj1Klk+dDxGNtKQHT+gj6wzPI
zn5n5DqnZ24OwX0TY9c5pW//s7oztClzOx0LfcBLKsT2KfDbeAj4g8U/vq91TIzkrMhvhepzxw5S
FTfoFNo0WNRbvfrz6zhZx9jbXwgcOV8PUZzg8UwwY7QptI6IMKLjkR3EIkxypmisSq5rNIHwEqSw
gYpd90e2fvtSbre+OBU6VpPfc1L45srSMnYq5Oj6TN5GlR+tFGuNx/zPPMJeKrMQ9+xI0EmcGXu+
rRN3grefOO0S9Q7p6uOuyEm7Czn2+lyfIvPsNdALQru/W78TmPOTgcqPlem2rj0PM7oXmoqkVrm3
KwTb7qYaj6tTgAhgnt5Ep/0T8CAXmDHJkrIV0tcYU5HXa1x+Quc+uSlnN6yg744S1DfSRGYjUMSW
AxWzic7srMqZu/RfoSbAoOaX4jtjLUXfm4aF/nGc2huue5Bk7WHknQ68Bg2N5qIvNsgvSoALdA/j
4qwV5Pr/TSAvQdL8GqhtCz3NEVcN+z1yi9SpoiWtMqVsquXHMbwj1Tg/h1kv90CoKPIRnf6+ElCm
MfzH3Nu6RiIJ5a52uZJ/GSdGBoaah4T8dOv9aozltr1pcnR9nv64lw2jF+qYQvR1cEwlbMTK792g
q06D7n15YwN4+JAQjL/MKf7Gg+uCQozsRtapV1cUE/SdXhoNaj6MGdF7KJKG5hNjyrWOMDLYMJpp
K29cvrrub42XHBNnaiMSGGZeucI9YXVjvtHRyJG/dE41+YfVRkKtBpgLlQa9Kav1E8jHn1pZkiIu
nmra03BjrtI10LfbA180sNlctqf3ippP81eNgPukse/Cx2pNhpiTfmL/jMOrrQlNFncpIKmTPBjA
njKeR1ZGPJgRmHssee3TCf4cvE4P5BNcDKM+amP8bUn3r40WyynbtKTGO+KU6hVuxK6lEq9OhccP
3/n8Q50uomldLM7UgdYshF3DRYRWBCDQxz9iyJzjmBzJJvC1g8od3hjD3tanMoS55NTrmaPgiAbW
OCU/n03uY0Nv0HYfNGLcCyPIiqlxSX69Ghojub/QSmChkxUzgbBeTHh7M/WgHoiHQ6oaizIp7qAL
7DJz2YmtnS5rN+WhRfOMaho8xBYHXUNC3+Dk367mXmZj1yUtAxxjR+n6JBnxv7WBvtabtUf7rgke
UoXvP1p3sj/LxWf+IEAu0f64oQbkESa9pmgLeT19IISrtgTUkc4yYBCIRooBR/gVlKWGUZdhe5aL
3RWX/suvWQ/zK4ROenUoB4cNME989EmtsvfhwG+HGty2KF8VJjTt54D5A+SLM4QZTkKWYg/PX3XO
bOxUjC8SbVuCYR1a4eFolzNZJXgVF7E8DKVe+5iNdQ7U28ZtK1MJu+szuuWy7eOEBwdOtczdAFT7
8z2Icj/HCrG5OYZfleuyFO8Sw2K7FXBkb9eBjnhiPEx4FNI05SDLcA+5xvDdWgGL0HNsl7z73Klt
iY7Crz1L+D6KIGqNz8P5+v2R258mLgFcefZoedA8zW3GeSh8vGRXmtZMsJK6sydDlvjSjxj6Qvcr
DJRNGPGEI+J9hO0XqPa4P47uCZsjyLd7ddSJksxPiXhRttDGwNaCkR51iMOpEkvA6b31Q8U3nipm
OWg9A5rL+bfTKe6bvjbpS4DFuHjgcpxcThr3wC+Ec5ay+6BpsnDmKxkw8peP6Tm1Qssqu0G+f89X
F+AZBNOikQFWbSXB9g1Bl8I+mXckvi7xTLEnYWJCV2oPQSULGRqL3EgdZ78UN3DIhYSREKtlAE5x
9k1bAd2tKMetzWzCwKoZT+dHdL+dvTD2zVOfIvgoUH2AP0WRjsHl9iO5f9UxOvFn1Z10uwLGI+HC
xfnjxDne7j7PbaDltKNwBpBWUjs+yy52KtIsKqmS8Yr1wv/bNybCMuWhQ1qroOnXIhVKoQ+y0e6j
4cDnW2Wtqhb8B1pVCWh1mizbmFZVtZYVostfYnY2hobXwQ+60gbfL9GIpKwGpb/KPLQhakT1L5uj
RhZ2RKHLnqOfnu7gKh6BdkFjN3ZJWXQz4pB1sCe9sK3z/E1j4OFyiYGi/llGjtpwGrrqnjl2I721
aiIF+nqhdcUUBNWKCj1GpH9bE8NVyzRsJkmJJ6X8cf5S9DU9a6/9lbgSS86pmCVfsZIwmfpaG4gv
b1oCkRPtOv8jP4Ktg8BNSspM/DbogisWqOEnPk3xGRu+7jWlvX2VaaHAz3bF0Afow/f0s5sGpBJM
u4AmO9HiXlxmJ+NEy4vdIV9YySdWcN7ixU1O5G5su7P6DYupJ0J0W7hjoefawrcqy/FBrMHokT3V
TVobo+CB+Ok5sSby3VT7AdRYM9rsZSJBUq2dLbKxtKcPSSmSfE6KpvR2ck9MmBV95Qpr4ZrTUWhO
sjO4FoQ0+Kb6YGPL2Dlv9k2ff9fpV8bi81lVPM6Qmz6CQTyLL9FZQhZt8xrjLuCQ4slUPhmRjufG
n4hmTjE+6YsKit36xrymfprmYs3xw92pFqoURTvgEyONbNYsShZDAad4YeF5RsWEIzu9aBhbqJVO
nWPLKHqJ66IN4VIWmGNhfmTP89MQfOC14ZlwzieDIxGTNMFh/5Y6Nw9AXPvITMvgIzOoBOtPqsfl
UX/2/gA/8hwlbyfuksRH0IxxiDkvLaUH3ziqFOw2xp7VwCxIHQdeD8HdNvJoHFBCytDDHmdYjYh0
cdJlxovHpznP1ltiwhTs1Ahtr6mz/rpGtPAje4FEkF7JLDgy+4K0WMJy7seL5QvXV78QjKG1mnPj
qP9/HHDseTq5N4TmT92PYpp+d7bxsp9cN7cvighjh0IkwB+qmluKiEzT0Y0EMsBXdEM/f+rd9hDM
L2/B+xOyvi8J076i4K3S4C7i67jbn10EcVjUMjbVI/R2rxT3GeEAc7yWy1sNUo5zGyC6OLndK71N
Me7dTb9nVGj6wi3WGsIN0+kAzBk51nzRcz1DFgcFRH71nxMBOGCdQoI5RA9cwGcvNZMhe55FsiF8
7iyz8Qt7GnQtr3MQq9ZyNLXP2YYNoY0tCjkiOgy3VgCiv/xB/LSj8Hn69AWhxyS+OloTExTgkxJh
w+yu70mtmjGetTTClef0odWZzKbehREJHXhFT8amCik9MaZgGojGioqxXcPqnIO/OZ/gU2tw/Dbc
BY5JU18qw/uvym2ymR5A60deHCZxZ6e9IGzTlAWrVre8QpF2AMiptq+4Icxb9f1BI9IWOtBeNipp
2/oAAburwcBes9fAyGqOpmNc9OiO6FjkKXqkCyY9KWBACLfrjBkF07PjNhczfmtJ+RnHZBEqiEyz
2JCrYI7+WehOqO5KnOEUiHsCD9xLxvrJ1DKUEEN1M/W+XXy1modzj95034+C8vWAqM2isNRqcdWV
o2KlOnIfrdvhZt8KjaaqnIKGC6U2pOTmEavy9GwMjotYIAhEh43LOyrkYeeccbcXi+ZZDloAHvrF
15golEQIm9aNd4muR24XDu4D1e+UsBc/5OCcmkL3gWQmM5yvOY8zfrMCwTOIiOzDRL5pxHo/W5cJ
1xOu7YFboDz0ejcWJRhnVZdqqaSB2QYpiMPwU6gCCp4uLvGCIjNzTQ/yr0V3BHjuIFqM0/AhA+xS
wVqirY1ZQHLDgu+v71q/kKHQDrlgX2Qj8YjPk38JKHTVdkSkTChOS194EvdiTmqnzhHCF2QgmUNQ
+vNp7sz/YwE0kH+O+56USebislfJACR2c7uggR+voWV4qKznjrdw4lSU7UYOnnmUOfezUpmdUFOe
SHxarFizaDZxUczTp57xJUckjzTFt8xpGH8IAwrtBLaFt2eAtfhacXsFvB63qVDrEufoJNggVmSd
lZHBn86pzXuiw+kAdvSQZJ5oOsrQmVfmV5Pcv2nodiutv21Nd5VqeLVDkj35ajKF3TpUzZX2teVp
8t2XmuVAv/SzUSUK2BgL1IdrTo5UfM0aVHtGmBaXRf+DEjYVJxL3yDOlk80A58gvWNh7NGXg64vL
oR2JxxJrwdhGpDQmEiePSPJiDVuebkWmSI20XvWuxT8m9IiqgWVp+g71gbKbt/y95/AuowVcUc9w
fRfTKoMD4pWNZ6W85yoyI7BcYxPFKgcIfuANFZ0D7eg2ZYvGSZkhZ5ItTGuD9JNqxIq/TwTOISWf
1nNH2wtxq/oKGfDmkAePzeNoWL+0x81KRI3RJIuA55EuOXIpB5zAFz3f4ZtY6rDfyBwWMVpskoD4
vL+ahdFtfSvxRfL1BnEvYo0puAwV1w+jwo/W3LYyl+F7V/GJVYIsMPLaVXEXY/d7Vnzq1qW3yHvk
nFUMMcA9PQK8JWuDnBc9ZM3lUUC+9M5F88vdZsAfOfCp7QuHqdItPbTjE43LN4o5bcQcp7gxJI5m
Fm5ATQ75tYWEQvAr/D5mnF1+Ewkef8OutN6Y53Wx/3NPNqS2mCqJed9erTU6vnohE0UwBP/29qmy
7ksCR8Jnk0PyDNu8+ppuUPxy/BHvfyy1Lsz3DMP0/SikLre4iNDXEN0RnjRwAGdct8Kw/rVAnOR6
lAd2pqezQklg0VZjC7bk9So/28Stz5wPFf+3qpy9ATjrR83L0CHWYW7UumPJ9wchjDfoc+j9X7IR
Hw51rUvWPyem9g/2SQtPg4EKft7uc0PslwLkGeMz/oypWhVCTilRB/iiWz08csGxo/IYqaCSpn3g
Y5rxz0v/yYIRz45rW00EShn+mlrEi0Q+yFGXZcfHTx1xNUVjPykkI6GGubSuUqtGE08YJXdkxhiz
ZL2Ei/4NfeKsW440MmAiQ4jrPAIUMrlSymi6B/bTW67RW/S/K9I+J7o7lFsQSmaZ0tz8wfSmtPyO
Tg6bp5Q/UrIm9O7kQLmhqtYRAmCKwY/oDoAWO0viYCA9vydktMwzZ6vtZQa+VqmGphHUvZTho774
d2qL713wn/YyrSCtruL4m2XwK0vUOBQBxDN7d50HmO5RLGIpdlgnSSp2smLl/0cAwf7rOUTTNdrc
2Is6y/Q0yDcGB2xlnlkHq7wDq9lfPPESvJ0RGqgn5915npEPCqP5kguBKVGBDirFaIlmdvJ0F9xJ
tWZzd60KLDy7VE9pZU9crXymuwBdu2ma+keVOxZOAKoQzAR9JEv8MIfSNBENtNK1F+hUiLTdbJ4g
PBYdZq2PCSJyeMhbEgceJV01cvl2jJG/JEbXTN5+LckKI8J1YuxwFXCZ6uJ2/uqigRAtXIACMqp+
PfLvCSCB+JEFYtoTfhwb4Glmxs8oGo6WIcFlVfdBJwOtiIBiiI/g1BFPplNzy+/YizIpwius4/DX
bOLdHkIgu10Gf+G2M47Cj/dK4dhmHbl9h9uwzrcNtjDscZaWLoMoqfBslcI3uPr0PfwjH1uNokcN
DacJI4Gg1WpbXQq4jxE+bIM7Gsh5UNIykHbzDUEInwBB1KzIvOekN/D47/D1LhS+e4We0YBk/4n+
ytwaxrMyJj4zoO4VHXVsZbnrUGlYwRCsVr/iluPA2pW5gL/KhUkWaNfwWKzDDI0xXLtQe7Sd9Qur
UbTEepZAoxvGVVECguEhMGCQzm3PDvZlZQqzQkyiZIwNipVJ5xd495MgJFVyDVXMfHQajrGDmrhQ
TE6wnLJGmyTlvXEON3/FZnaqYQm9XjR0xAfguy1RUnm2W7sZzRHP/ZJynJqmi2Uw8C8qGto6NWHo
1BB9UHi1Gd+dbjPogZlGfp/asCcanXzOvyzFvMVP/xKovCgprMzLU59hrryT7H0W7tsikkpemcEX
XHZNeFgtDGUik4sMQ1EGMcAgxHeoIL069cyLICJbFDco6QrnqZ6aODEjc3NnLKSIrAji1WnXjult
zkrS/Y5aHUIVcNVQA3do/TPd5g3uXXS59nhenZmzy6jUVD2vKZvrip++tfywexmv9CW8Z8+PH4j/
xGZAvM/DQItcYxoUXJY7qV0kh7q7GqqDX0HyvPUiomPBT576gMvtMxqmwdziBWDdWA6sAQx37dWZ
lRLMfzdKRZ/XomI69hU2liueppdHDzpA29RgAF9lo8BoUZOmSoZJJLdLTESAlgl/RQLsFZnFS/Qi
OwIl0y+/DkgdLRfkhg+orcKFxekG7iL2HHI5E8MKe/Zg+bWFrOCz8P1B/nbsnANjUNffUp0sWvTd
yXJU5PKRq1FvysM2QYG0kR+VuX/0rXrWvnvVsXHaZpx64R5OTO4NzVzsKYTbLedDVZwMp/bPvSlH
dg8bnohwQckmEyEg30+X8BcJ1bXIAR5X3mlwttHLfNTbeYHhrRPXsympdIugiz8Nl/RvNP212gNE
NBl0kQuSTTkurOMQFNfseSTYLjPlayMrNffD8xw/Lt2XmIMIABIvEqUMvpYJPbFvSEetAwE2Vtbs
CQWP/FZn/dgOW6oHou7yuTLRRMFn+daGqsKC6rOrs4lEyqS96U/k2Db+GOToD3Qa9mwDtnIL1Epz
89jZCSkX3utYJ57wwmo0PuozB1HdZ2/mqvZ2SG+MpggbhcBEBKNnaHUKHKb2vGzI+/1YHQ+hRPLS
VoVn9lqfMJwnV4/rmcsHOkODYGoXVFpXlmKNMWAlilJ83zvmDZXa2BO2RnK89IefRrb0ggMM7H9E
S420irHKWYgZPaZdw5Y/VsveFLxrBtgGbLo+ammTC3/ZEfsn+ijKEswEt8SgjeO0q2FTzDSxVn/g
KvWKCoSU1P98E2tuGQiteNPhbE+MDIdnZ1zE8pCsZDvWkwkpyz68cMwTBZwayMPQjN0QCXh70p6V
yOudlW//8W4zF7IIquSpHiK4SGwK5BwpJ+tc1ka5O3eB3VdlYLj+eepFepEYJlBCI2+tKxDfJ6mv
IFNSFYeZQfdUmzofsMLGygCijI6Q7h6mUTJGsQynG0GyJahd7sp1PeGBidpEQziS0kWD/EDGAARS
0vXly1nMvATjNQYW50zUaeDPBaGqNsBRNoTWrxO4UNO2p2HKgak0EmqrbYPPXhsv2DBXSMY3I2AC
YNKSHyQyVVbqB7PJGdJmeP/HUXfdKuXgcFrHFH5uzCD0X5myXl5KzgUEAMkV+DXYoTkUNlK3OuvQ
OIbSnT6f8pXIUcuydFeUyASstH2CExJwhdVdGzNGXiMS5a80nesg/3rQXPgopY+r8kOB2s1yxMci
oFRFcNMYvaCoodprAsrYOq6U+SIzULu4zbHj3PlBQ6ynI0lz06DTexZOzuLslZT9S6/wA24x/HmO
8r5rYcZVCpiozmYxGUlYbMVbkxMvSrw9QqWqDXTxPIxsLvVQnqS0E23mphkE8oDKdIA1GUVesDma
uqz5ovOXNcsfJUHYBp0hjtSo6I+wrHGkIY0DfG/k1ofxKdXOELyEwQlLjRGdoit5bCIH08Cl5ze7
aPuBnpQcNYCBzFYBHGPiXgyZ0HVqMHOKVCRm79OhrYbvxRLSm5MMLQUnTwIt0QX/lbnfS0aFB29x
x4ZAss/xIWbirML91JDZCf7TYhgWguCGV/fpNd6LB+zZyssEIvCQLh5YMZ/E5GUba9IiCxJ8GZSG
WzHoERSFT/aMc1/SYQCIiBCjTakC7i2RvlzFn4Y/AMuXP0ItGW8zw8wk08m/6KOriuEvVsn91KF8
qznF5/HVYzwVoXERPYfsx+HogNEBXc6l+JKZnzeWh/LKWvQgSos87qmPoqafqZb6LuGo1s3flcQN
6TVrq7oZn8CjMshwYQuHnaDlxlBg9GV/V9PWL8cEyoZfvxT+RtJ+101RJ1ccYH8Nu3aKTV7rz2q/
78E4SIPntxw419Z+TP/lucwsW3pT8L6mdIHnDRFIKMmJ+NNM/cSB39+iyed10dzAwumFWx89v/Ji
aIlgTcUmu688Rx7YOIyJWapRI4aOeIpMRSbkzFu53D2KyLtsUHyOjeQDoMLLRPHv/sHmIi+V07Nj
cvlU8bQLFfiumH5vL4wRP9nqVhCrCuj5bWZ17Dxxh8XMAwFGk+qImwwjxCBxzOK5fWR+wBPMY7zO
GlS+a+M7viMHKWSFImUbg493UFTikwdVNbb15DSC45kqkZI8xhjmkUexZxLmdQ3B+P4Wk5tgvHYD
EQoCcCf+G7wn6pUdFuelElVDrvsGpeuq2IOVW/6kPwmIJJc1mS1EHDPBqq4vk+7JpbZNAXZNXm6b
yZWke1R6Olgvx+wpSPFafi1o/kDsbgY0zlTYIj0j8cdq8R1hGcHhkCmf063bAOZJ8Dyvqxmm8rVs
jFBgQK3QonYB4REbe1XB0pqpEKzRMHTcjrGPhgsLn5EmK4NDXwVN2G3uoaBnnFt7bRqDZKhq4egn
0fZsydM+K+DsGrLFajZKQEbbQ6xOAvV9RZAMVhy7l5ZQdGNphqe9hxsm3GGUta4vvXjKVk1K7DM9
ePEPZBnRwhnIMuFzATCMhDW9BHfNh22mo76TiwJo/b4zY4YHKlFgERaS6Ey6FK+bJTbkzWKg6oMf
rTQgtz4YCPFBNyCv35XG+ZV9juB8U3aNMTPl37WbH20qPfqQ80qbOm0FeH4Niy0ry4qRzwc/AcKI
HUGnqPG+5xs0wo8VRvy3B05dibQVEIR7J8YDGhc84Rm+BWDFz+cT9HyXdRxGSN2LsMvS0XIpBno/
CvxlR1EuAZ/TwyUL0/yejLWsKiHDVTEB5rHSyKWq86SrWOX3/csC4yfmGb0CLd28qAQ+JgoA3BXC
4XogxxdhxBCxbpAfIJOcB9Spr465gw0D5tzhKVBuqlCIyt1lYdW8/YDxZHdKb9i2rXsPFmzIdQfb
D+g06lqKdaRisQd1TnXKfwxNB5DAh0tMV5i5LfFl3pNcpVg33wQchii1Kac1OhcM8TNJY34PJAM1
oj0U/YA27bRVoFAE2bWWI2HwdjViEBGztB8MwrswKIqjfNtNZMhnGyerBUnpWiEznwcYZPRKpDAo
1gzUrLifYvJSpGUlv/3Qi0pMS0XCwenGgWv7dfXNr91BDzDyRrs7RvUb9GxMUlOvttw1uJKJHUO8
B76IfK3/JqY9nLU4NjAytESU1HhY/b5wn4m9b19zD9FQT4Qsd2R7hwQbMXU65ZANl9Mz2W/85Lfc
Zd1Kutg6kgRN+SlFLwRdAmDAEwnL/19eXgCyYFum0wDS6qaQB6oHDVyW8SQDPT8wSD2JoZradxHm
4uzzNnL+mqZ1oWzt8vETQHJA3mqwT9XxHF39VGwMYCh89Fvodaz1BnRL+Qms3ZNN9xWbBRPm1Zg/
UJQNcGs/Ajxy9tmPUC17ToMOMCCCrKAMc76O3TBWOyeAhs9J7h63LKOnM3uzTJJTty50++IE8p0y
W/o6ifIcHeIm0KGJCHEzTrfLASsg6g+coOka/Sm0GgiTJNgLFBbt2Vlt+Rs9gdn0MlfLLfWUCWog
HzBTQTQrG+fMfovCKPdlaH+3GitmadlaxUWEoIJ6rl7TpyueTny1fhYqqZjtqmTm1VG3tJjPmGhV
E3DqvPV9KCsSkXYIzanLQiCDFnI9mwXJeQdoMqS1t3LtS8IFjpX3A4Ey6yH8EcvKk4xQXrHH0ExD
tKj2DgQQHdVTH1IamAz/7MRxHbY7fHQShdC77C+xDDCaQlNAVMPxUdQ7bvrZfMgpjLkwuxoHnaEV
GzEY62wLYNYo2Wzc4KK5XQYLUoIgfd7gfvOxYHSGc9Z+Jwv5FX1ElZPVbjAKYCb4YHcL8sDhmXX1
ojDEEJ85wxX2COHk2NAj4Vk7oVqCtWjnRimNLUDeP4RXsW4LWFv0SrWzliRuPTshTkvEdE+2EMRS
NRAiXuzVniXuKukJ658twNX426CXXC2X69mGYerAFSAIruRGlssgEWv6uzjY9pugXhCsNNJ9A9Kz
gb38VTOxqWKC6ulQJuzgAZdWYk+DG8VlFznh9k8mtT6qcpzbMU5jDxpSgr98gO70YrXGV1eZ5v2v
7q2fODIt6DY8oyQxi6Df5bk6BnPoVzis7NoW53QvhYNiKXsC1j+sW1AGTfPxhGwtmj3qVTff2GHi
9kP7w0WGh5zIeU96x/nDW5RpkP8qnySHUxE/6ZpGqwsCAzcGGQPz90wViPrBVrcBALhyQao278RP
1LlGFNf6623dDHn7CcvJEJN8jVLAV4/lwkuoeu/19/d2WaFR6Zy0SiFcYmX+lATnpVR9/27yj2+K
QGhSo1WuMWOsH5ReclYSkI5JFgdVsep4AJwDXxpuBaD13mBAseDrSfqEvmbqH3+msQSDJA6vnQJr
05Mr/jRiLmR8lSaZDE0XFxFwkYZ13rmKzMcWCerJXbkrhFcLgjrow5avdRu0CZo6jUlf6lLMPZTC
n96UktkxFm2DsGk9ex4W1W4MeXFB1NQnbKgVjC6/JWugwggnp8gmlxSmXP+xw7qS5y4F1KA1n/1j
2EmN1pBpdmSplmZBRxCqCB3r6ENBQQRn21vMNSfHd/GKrfbgS7NdgmpJFZ23JGODheQyuPKg7osL
akY6DpvQPaoz7+Iw1nngWRtGYEgnmwiuYL2hboce0ajwo/sDCmJUdNir0DO8QMNxyIQ7C726tbhW
q/JQhgbgWRuH4H0Bjyt+V0gnr7XJvMN9/gyTGI7hr9HE5o0ea2fBvHjv9QPrTep7tGY7ziwqLpxR
fM0hN2JweXbaQ/bv2NnhHgmhdvHa7DoTRTzi3QL5vE3QRkHZV1bbCS8/1KaKIedwW4kWpxI+xjAN
VQjj80+pPepToWJ2HX/HWNF0SZJeiQUCbITxVkJcwjIQkSRvzWXsCqauQXqQc+bVBvyrDvWkQYy4
caeB86oEsFQgCNIDh4+Nbg5OVwztqCuN4L1OEWf16NdSShu4s+1IgXUcZoDoc4QB6uCKTEUQbS/a
TbQngvmbBaB1feKRTabVxKYzcqeSAc+dSnPLAPwsjmkPao2pQcbHIy/3zVQaU65K+jXX1ISSvkSn
C2iqt0u3Kj0Y6iVi+r7BbgXX0+nhAs1+CKyd+C3BdEo1JYXNvz5tfXLT9xB4SkRW3BIC8peY/dvB
e3osIvZeNbgO2Ypof96wkiWwV6PYzDM38jCmRIp1OUPM7RagDWNMFKX1BkQ/f7abNffNjravn103
TcURjaNRZDu7YVOgb0ZkKsPIb1CR23iy0BXu2CRWjInrgV9cFXpMc2LtS2ybSh0XKgij3bx9msGk
7fiYg9ZyTFjMKZrc8zSqo2hC5eazdxqmkhLccEfH0b+1zN4ULCvCaST5vqM3WQ9be9Wral2OEKTJ
lJ+PasvxpS5ymHYY/vtWLobM7vnIa0+0IjegSQwcUB42z6M9Mnp7PR8RAnzbx2np5eNwrQnJKaiU
OIhrd+Z4uhr/fxkAhZuLCfgfmfBHtPj3vo7+UOCY6wOQNt6IlHaqKymJMGEjndwy27g4wEuIQrGu
Qkubj+ExKpHHdBQQQ2hn8zKyntWSDpH50mKnD+A6oLwDh/m53/IEzIguhXmhpxoOXeDfhOfEOEKv
D4rwAYzGi6PvaFXYyjNSFhVQC+I9J43Rd/SVXTbQftoKwCkQAYurgyvdnJpCgGU2bp9INUjkKF51
27DGv5Yy0vUMlH7oImd/yEqAszIuqjaRSf05o9SS0u39qa2sKdJ0NpSmeaFvjxAYWIHXt2Ns1N07
53QIGWusubBjommzHsNps4AVxOCLivDIfb8L3CyY9w6Ee4gPrEhgfaovT26IrErcyEKgd2J6gaCa
akAwX75krLLZsfLaHnOwviixn+XUF5ygc2CvukJA8mtnBlMkZ8IK6eTY4l0pOrZVEEwf15RS4CIt
jzqpm1Nd4c9cKH2c8KYnO6D91g/ICoL3dTKT0vKorfzehmR/kGp4UZiu5MTapQzKcd3amVbMeLxy
TxBf2VhG3ciVKsck+ovjjB1gGoWNCjjoSknpU+RJmTbkHw8Jy192wIc8oPQXc1696Iq4hKFRDUrq
wTiu5FsBM+KJrqXtq46A67Id4/9rghXqSR6GyF07QOUMwe44s7I/uJRfnEwxLo2HVlR/CX35nuXt
UOVWg1TYArdm0XExGqXCUxsxYFf/XeyXZnrlBZRcwffDo9Pc7RFatfNri85H+0aHBZ5G5QyDyCia
HjpevURvQzaXyj4fm0LRG3vBLgwrfN3D9Yn3KM+jIzVABEeFIHRXnVgGHtn42CDugYWFU64NWhCM
ij8nZnreq1xPukn3M+B9DN2X9X3/8B4H0bem3iZUMym4LevxjC3uu00Fdw0QcGFHj4o6lVAj4dMb
uN3vN2FvbW4+Kle/S5wsotJygU0EQZTmNC4oKTrSUcp/cCt8pT+B6/hwBkuwhY+JWb//UVgQyQU3
9BByAasC/Ks4TVaGW7kAW+BxIjO3OA5olRs9rHzHhQ1WnxQGomdeDQsSdQ0RhdeO4qlfAx5LFzUv
eWQF+LvU1wJj+eNkUAIy5+Khqth6mNhd075k3cBO5yJrdZHCmhGmL6NxUrCDjeBt1t7VDRl3oVuU
zc+148jOjITpGH3XuLihfZsQd6DnRVn/HeGuUR3S8O/Zbz0gL+L5zAQhjN/tyfJkIAGfKU7AvInu
PsrgLyG3SuxVMQKgqY0dRpURySxozQfhe83berrnhVkBaaa/ujhC66q4s/kjwGmjsFaJ2oApaslb
YTmxyxE4paOI1UDCXFYOhD2jRBfZAYwDJXZQy1Z4OHKPL4updOZPUAsttq/oPEkojifwzqfUTCbM
mkFoZU5buBdduMLHjic8pdTr+KzC8ppSNIxdiB49qrsztGnH5BIbvS0jjZ73B/4fg3gkMJ6n66+7
WtVoDpNf7RzLq/HfrBAs2UuV/UVw6NQq6zP0EkYFSLm7BIMt/T1APpkaU9jSkRfvNvajqHlHL7f2
cbke3l1F5uS4FnCYtARLFFf6LLpPGaD8NxYLKOgVYFCCJzi40XCxTj2Gt9oCvvcHrwCSZyJZPhT7
UNOzaPhHymsvNCChiWBVLkoxaon66w6Fmo0dFrT8azMGl7iJMrM1Ve4XXRPApf29ji5jDsJzC7CO
QH2JrMIVH7I6efI4dIjGyKx75DXS4HZsZBx/DhtrRrjWgirGsxTyqppKnVic1qnLC+55Ala1kjMY
IbRv0oDt28mT2l63HKddcQTQJ/XAZd73D44kWI3vMeO/nuLjf8lw1c9taFBoarN+inQQJXNzenP9
xzpueDAq8lm53oghx6OAXsQB09RSrro0F69mu14L4a/Gi37GDw97mK+6rzvZ8bjoj/cV4dDbi9BW
ckYp2oxWtibFrhrZug655vJQRQf6I0DQtSTykFZUa8/EB16USSy+174efLvzeP5g4beDNwLis5Ga
Cq9xvviZR+rC8/4pM7uKPxbNQqP5q91LSXdBT6/nXY7u5qx8XB6jxBYuWYRD11ryekZPNKrCf3aB
eZFl7yy/SuBpMTpi0lGvL0swGW1MPfQnQ531wzKF/xTAeyHj+fctg2Ai0qYpcfFAGKzE4isMTPvK
8+27GxIpK0/np9GExWIQ7dXcjaOJEePLcV8gZzqFkR1TGTwtCZ5/K37MhpFQrXgTa4kxq6DEAao+
8JnEuXcSLQ/7ioEZHOJyQ2rHqOrlInSnlg9UoKub7i/kS8/k8zGWXXfNQCdKH96LZakhzR9GeF5o
x8zURyLZiAYPzOjqYEEJnsPVsSmqbMDhvyablYlzgzSuNB9jfEyaV21TKQPEDvdbBjja0x/UoHSE
mQvzi1eQk6pMDG6rHmcjL+1mdQiu+NOpUmM4fxQB3Q9IR0ltSBPIErvI8pMerEbRnQeg+lCXA9Is
ADtKEKGNILp0vaOX6QY0xZTPwVjt4StbAGzBXylBe2zc03arJD9mKHwS6g8iW507lqQ+tNDUBfYp
46naiDvPK6zq71WGqlGNlS9hzdoi0agOOxcWQBxUd/ZAt8bpBZIYTdrcCPNw/sInNFY6FCxdLFm9
agirtnQ7HgzFRSxdki7M5tnbM1eA7ny8f+pGyfDdd0QhTOHihLk10oTzlHfGvYlarkLJ9FojesvU
iS5F+9Deh7hq7TSr923gLBuMLR81F+Hriap0/a+tlYvHEdCjhqBd6IcC8EW1/9qeewCK/mwLbGA3
pEj+6lk0QsZhXzGQNoAa8Qb3OwYfQRgbvk7+RbGLxHGRqwbKwhuIxZM19phIUCcxjRy4nI8h0uoG
oKdu95PVUkY78WNoTyErvtgpDw0bRqqpj69NX4k/ipN3meOLj1dP2y4HtEAoOZDLlFXk8i9LF413
HBR249PZa4Q4oz4VsBw6FZQFw4zhO/LQpWvYf7csZ918EUfSION0jCA36fEYJT3bagGLtGD3In7R
BYT+H860ne0YESj7CazC6IgOpR3Wq4ACjA0sYhG+JVPjvklmos/QS9S47i63Em80W8TUbukdamNj
RmM5u/zC1ZpzqnR0nhaNHK8pnpLEPr8Z5EWyRYJRgQZLE5Uuw41rsZIRxCaqCwh1nrg0Jd/vYQPS
+sDZ4AzXrtEQWKeNFcV8VhhQlh6BRaOkKyD8ihJyyDwzC/GnXRxNnrrrfAMptRJklyL82jw2+GOg
yS+K+t2jIpgfCMnFfVVq9JCyPpDOdXEUB9A6l5x7QE+l+F8eJLVs/KAGX5+dkR+p+dbX0liXqL7o
28n0ORcoT9QMSYBIEkC6A8/34yaFOFjWJ/Z+yctcAUzI5+xVsMr1s8xHnBsOTUWGGyM8NL5C9/uC
JaYY2woPZvbUgzA8eRGKP8eFzHt3+R0ULN3khhSYas1J3GPCgAqm15bNonc2qiQAnkH2tRq7ADDm
8AmL3V8TkQGtLHlwfFUOuN1H8Bcnz+MtIx2/HRT2PD59AfieKVTglxT7JiFcpLX0b3AC9PR9gQ73
z8pHFnrtaNydk5dd0GIA3RdV7Y7Hsp9E4VhYAS6ju5wj/STFAFlIEh/poTpTyxwIWCMuoXSB8ONK
J/6P1zb6Um6L7rfWa5ZQtORvUs5kfgt9tEvFAwQPj/fiCBUz3oYM61J9W53F3lpSqlBpxuAT3tk+
2pJctLLJUXAJHV6MGjsvaHkWmPOABFH/clp6Ik1wBNFVWYLs1S4BGYkieYmt4YZzMJhwyVfDVMAC
Z+byoI8NhugLWxZ1kwWuREM3h5kZE7CvNZwbxNGUlmdC/Y5Q0OnmhcPDtQnVTGLqQfrJ50o8pIU0
xq2/rXMICyV4c98j/PguAz26Ib/2AIdPgb7VQ6KRKUqanhpPGq5tGNYCFGuE58N0VX83Kp8vGqfw
Cv4INslV3MHf7/TT4ujWf13798R9HXKqp90qwSsIiJdjN9sTmqchDy7GA32CppwCeQ4uaC8J2Vx5
nARhtWgkx0s9XZ4og6K35FF3PF3A1zEJ7SKMyJEQtnlhpyocL0dKDNJ9L2FbeS5+1Gahwa7wiKRI
+cwrF9GxKFFH3z3PTxbNYaGaY1e9YO4FBDlQzsTxer6C5p+q+dLHwswFgN5w4Im572ZW3tCYNIEC
9CJsW4ltHLCoIoVv0j51aisGxl8BvCyCubXymZdTbJ70pwcpIyM6t4z90hTank042r739gey5NDn
lGrAC/3dNUCBCZnwBdP9szKVsahxjUSX7U5ujwCH39nEqrExpyV6AU5bFaxUuCtnmFSH/9d4DuW0
SRgV8RJFC27J7rhoAlFEM7H4jTCnwlwEaHysgjLrnlYV0gDAUgJLmTBqnuK4f5sYxLxuSr+wA0xA
zf2ir0E5Z5iZ2vh+87Vr/f/i3KwlSkHh30Pj1i46MPwrEpckK3cF9JvluNAXCXDfIf05+f29QAKM
C5jUXGigWR8mqqyR2L/G9X4cMn6W2NzWG5cJ5+rOYA62NT/XlGVIgwrzPopTKFt4CtSXpAwVvO6k
HgUzsRWLVBzydzODwoUCj3jZWlIL9hMOGlSUIvTqBTzACBRtFe/+U/LBdE3qcEL4wDM9CuzfGyik
xIo7ht+zs6oL/05WDp52wFiy8vm4xwk8YiV9TqQxXyLKjP9wRr8fEAi9e0a/mzsKeDqMFLMMe05y
6JLcV5Rzh5tzohfLmF3Fw2n1/0dNXn2hKLbYH+6DOdmDA4y5jTBVxhlDhqpzklgKF6wU4rYCb12x
0Lx5m2Cn8v1GipofFT0iet9l+FKrWoUS0qaVKA6jwQjmtE0tTQDbdNWd4P7nTcOMdtWuW3z1b5gN
XVs5+jYg8DLmpP+vNUkovSEjKKIW3Aprv+e3VbnUoNsV/eXBC6D4Rp99JMsFZUbvVxIVmNoSpfSk
UTLab+nUHYaZNDScIxGFXx2P704ZF60V2u1aJOy0GWF+wHBnN9CGZIxpzofwNyEtGsvzdUvtGTEN
zt7jrVrH6PmO1OA07qlTjpoy96qN7DjfgVpQkJk8WhKtkEQsGu5/3km/X76wYOcXG8LmzYvT41uF
XpG0uabDhj27glneeHmue5bvaYdE3r6X4QeM76fJdWGmYZ9J4Eq5I7zNFgZUe6HklYuTb0Hqf3n5
nmVFotD5GuJck8ma5184DUwrYNl1ThAHN1dE7Me5dwS19aDlx4rrnNiXQ8ob4ma+9PjotOOnckRM
PrBpcckZBLrfxCa1aEr78IpxJhBw5hJQU3hfhWN3fxD8RLOtgKJWReG3EZp2YvQFQm1IHYuU4rEv
PafHx0vzQLsKoZVXC+9hp9Z4dC66V3IfBvpCd3J+Sbs4/kSfwQadN1Fzkx6gEvWfRLk48bAdnfdD
LtgK1QzcBAloOZeJ/2sdwoHz3sGzsYe+dipMN7DUWIQNDxdiY06xs+cHq5uH8snzCMoS+EjBIRZc
BEfATQaTzg8rHxUpOkjSVyUZ8Fy58WwZCSuTaB9XTFcLlysLO/9zIS+m7H7YAOECjfa1aoXeIHX5
v1Q75im1dPeGvtS4hAUTn7dbUE8p4uLJQpteNZYN9xi0ILjC37yzAqH60mYqJG5qhrboZK1fp5YI
173tPgTDtR1DhhwUXrzjysZpZspsfPzYe8/tXQO73yOSUgAkB4M+xWfQNK11SRiq76mkIN7vOF6g
HSSBGgkWCksBF6AcZLz5eQJ53OkDiQg6uc9qAmvss+FODt+KFQG+PfPFukpexiMNwceAeFaJEhQ9
vPUXK7aP/SOaCjXXvwH1sjjyJ9Uuh48MTeZTrooRqnUTNXQQbStVA0W6CLG3VVTwtk74L5eoG4tG
m6MrpL1p90XzN7QR7nwSOGiBfExcANLo3wcihSjHYjLPYqX+D3RHksyAp5+B5bejDNyidcF+YJfa
nMAlLGX+y4Rl6uPEbbQpDD6CkwAau6/Q6OdQmlgOGRrcTPvYVuPMrmbHCf3mY1+fgwYnzvBR10bD
IaA50+psWTtzqekdolRZfWhj4lmWoIF/AZy5CasGhqEdnIpG1VI36AgPeHL3KGbuhwTOeX+coGZV
zGx90rnRqxm6toofGr5qKhdoGHUK3Hoplsl/IDE+xKEHgM7jBy2McS+Fu2AfCg4Jw/QIif+GrGE+
AMPxIqVSK8+ueP/U4lcUHEXgIMNBYTkcPrpVZavPC4GqxyMBjr7cdKRGtJHF4FZ8wcUSLMc6n0Jm
eqzZ89ANI6LBpqbTk0yP7CSTnW7WiAaUsTosoW7RSIyBD+E4OI08Q39Tw1FVShecvCuBv6K9HTVz
EP/1sBR970LotIDadlq4mJSH7579lit3XPCgdEDIylMgwtpFdVdeMaLBKvtTeCg7rq07/q+dmUWo
Q9pgR/+9N+4d/QLuXOjYAe7ej9xdX7fSJ3Cduz0N3ORhMuN56pP0tfRLN8PsTdQcJxSC/2t4VpzX
za04LcaaVx0rqbpjO1ulN9c2j+yeLK4T3lD7IA841cQa5sVM32jxUHjQkbzWJmI+/AZVcENabw6X
3xHw3eHGaodjpuKYbaSJYBqB2buheFDLuBtcJffErOCjL/tSL+5LuAkz5GPk6QLa8/rhcj/cO8uy
hOt0+QWzrz6gRIHXb4VEMi8sbq3YrWkJrXkevBZHewheQxVG5uQGOChIkwcjLH3JQ9/tIbrT0Lj/
P9dE8WA1jMo6VXP8q5Bd5HlOexW5WqrZGgHusTyXuaPkvrxs8UlRHsyrAHhJsYrUq6zvSHlNEHZV
sjnqJHgf9zGQtsrAJSomDxAxRbN1+D+rIIewlrt0eXqWr1jtv/giLPu/cGXcMZFvUb3nlxxNGLQ1
PyHHi5PsVIZmDbuqfmtrS7SPwX4mfi1VvQ0Ey2kaMItPmA2Invcvj+ab5wlzqoTTcCu7AdyHx4SQ
9kAnipWcJ5rN+WEIOMHLRzVQuIB9T1uLk0Vn3Yla6ZkXSHewm6CDzhpjVJmh34wb1DSJyIY9zVKK
dDtBdHbwTb68gdcJEmv8mpuWZVx0KAXwsq17PpQ1Oe6ZVHvS6Ys1uRZnarQz3VVmq0XZXral6zIg
6IlIWFXjUDxJY5puhQtJq6B+d63RWw+/fZYCv8nIpMk3iQGW7BYQLkEk3egu4B+nnZefZY7FLfRo
SQ+RUA2E58DydIvChq4WLcJrvyKXlMktBNuv2Iku1It0A4TWXW3ZrpPlHYZlKv3vg1HRyvyKuOz/
lJe0rbfQfRNuD0BXWIIn0BFvZXqnY0XRTwokaTunTLyP7Ov/dFSgQVclCjynNe5p3vGAySmYg4z2
Z9pyDw+ADWguznncET5ONcnAaT8LuTru3jOSfUuEkyT1CfZF2t3KzpfZc3CoBHZsZXZvGzeKBcSF
HTt1G0IetYOh91/hbNzY/C3hU8RQKAJ+abwBPtFH2XzbiI+rjHkJicpWL7X3icfcfESsZ8jurw9p
ks9va9u9OU8Kyde0YelQF/vwO3qjAHFKUlr/JSZD4PGfwqpkbdvmTqINgnaOAlpMsoXFM/D45V36
RTNCQ8JUKaej0ezkFVUin3N4MQrqpkdx90XZMkl8jS6pq8BGeFIFOwTwcvebbIpIGX7PHCJ3ms8X
w5E9SSz+JyRZFBJWKCtwc7A3Vs4GBB1Q37oaFOBUqi7lTapRyYL2ED8er+eLnfbDFNDvCxLRd9GV
rxJp2QQhksn6LJ19IKTqr7zziMyFo+P+SOtwB1sRVOIBKV/dSDWGgIFkoUq7u1c/ItNv5y2NiHYa
LziciHcAEEwHfNOBvW8bGPuAXDUk00YGtluHg5WgXCxuLX9Neu7k/EWsMnL8VwNN9BR0J9K85TW4
AxVKz7+U4uMg43yL2WVEPzij6Ky7Q7oRC+vXd1QMsMF6xt+BQqIQqOEGkc7y6W3bMGGxh4SVNONP
Ps+iIVy3xyvJYbcavXxuVBCOytljG7w4KwS1RvUHVtckLSP88T4JozoIc+jRwMFFJkn3R4sihVSb
q4nLKF+mfq6faJghMJQvnCkCgQnPRp/YaJcJHZK9FxCsGbmn72rAYF6rkQR6Kq+UqqAO65gA9sqs
2Jxh8kd0PaGkkYw0tNOm3YvvVKHkT0HNgy0KWw/NL6d26y/m6RarRctN1TFe4w7MTg05QdHZMMcc
Dkpj0r0ZZxUiRKNwemQcjX5C9f8ztm6ngnvhFjHK9nYfHOb9MCQ3UKyVpAE+rMCtIql8E8NrSlTr
cpNMjc01UOAh2GvplgFdxoZbDt1VnEk/poT67n9HQuXf6yn/mpaWf+FLzrVJtr2kpe7J6KVcV+lp
jbX6vHEYFcw25ST8Vnju5FP6h0iQcfCN/JaoR4QGZ5EKSA2ntBpl6pT7+NStF/UCNKTVrPILMi8x
TStS1p2wxodk23/1+XC+MndykHFDcRmCqIO1Bp6FpwuyuZxWP7u9fVscH6UnUU+zDjjDDr8zN9Xe
Qjl0Nx99g5l+RIyVXgQ8XlqPboIf7qKOQM8aAxIjNfcLtbY1KejqPVH2myEdRekqfmNLpgtCTWOL
H/xgoDI/Rtxr/SIyv6V6IPQVIpln5DPqpCYQo1gU5l1craVTOiHCPQM5I9V67RpvxMC4KZDONj+N
MdJ2JeUPnQusSMvMY/+8osL7yfcN8WUMoTRYOKxh/orkpPxvlk3T2pmACWDghfGqu++was8dlKX4
VBGGAr5fHemRPoYw3eSHZ+d3+y5rwq592NLC3yLRRrd62Pz00R0ScCU2w7Ux7UpJeMJNB2XsUmuV
Ym0TU8mi9OwYrwkZ95ghEN3b4hLfJn8OK0AYZtyT8YuDSUjKBFAhVRpNdIBENFO1KHv3rKFQ/58I
hY6Zga4uqnoSFa2E6fsM69fmtjHUCE1tpVUIeiixkg4AuBaGWwzgo14GeZdD5YHH4lT13237Rees
jcIZ0O/LTo3pWorVW2pHnrBJ2Rixpdi0kpwCdTd1dU5Ghw03EMUcKk8QuGEjGf62ICriG4aEpfzI
4j9o43S3gV9d8sVvSpH30/z1WVjVTozj/2YXwpAMp6XQu5mAgazDW6tYHkSQxS1huYli/2cQJe0T
0UoCr1WGR4cnfGIcNegJaXOb2ETXjw2mJ6lp+GJhqS9bFLXOvJUIMbHZ3KqjKWty2TOhTSPXeigj
YucHL7eL8d1KH53a6jLFhfn77TT0Ic/Qw205pwwvsGH1euI4cu2Gxdm+I9CCVl+qVBokJ4PKSUDv
ORc/Q5xPzf4/vhy3tVMX5O0ycAJmjZx8oYPbij4fQflRXpWtF1Uu4JbViHTKEmPtnkWXHuN4M78m
nOjkigr/gdbioOrJTKp+AD9xqUOQ+N+TSJDRbglFmML7nyFtWfZNqnl7nDide6wz1TNyGea359b0
7XkzgPG02g/7aem2/QUhg3k/6EJqDYCqy8jJ2q2q8vvxaI5xYHI2nzU4yTwfyZnMNz1J1/0m/iEB
U/zk8+BZwRkliX8gkwRsg6A6RhNnrwQ15cFA9ilk/BHeOPvrG+cc5Tax1gX39c3nXtpKrxCng0fj
dqmtnZnPAnRWqH4tzDnFItJycAAA4Xx4QKcBKWr8spC8lqGwJuloKsIQVqD5JifXGLyZiXkpScDo
dO6QjEFEG96HENNErJZPhgo5Da1BtyHJyvMXVtKXlT4pGcftrsUZL8DWyd+xJLtJfdSLWd/IYYTO
WKEOKki7tUKm0QJrm0K/KQlib3oxBszB887n5lAqWuP8PSK5dmy2uZQ7FKPyBCWaa1qZRIhX9STx
+Rc/9BG0zI591KPBdlnYh53PSfo4Hyl7Kx/h+6nUSKy/PEUNGtTE9fy7YnLHicnXmyUuVuE8HQ20
SwRy50EvE7KfH4Oui4o7AKY0I1PrCsccEtI1kwFANJzXBWu2MJKyMPPC8gtXt7DYlTI/195a5F33
qm4qOcTyYMhcl/UoegiM4jha51NQxJKNsNBnh+FZtqwVs9v3UW/6zSkWDeLtZLd9sb06Ffw77Ds/
D5Eu8dBe6oJoqJwv0MGmlSctyel/RoeTNHaTPFnVGT8KCmuaxIrrCKwKDajnD3jteitfI2UWq9iw
3LZUi7NZjvFjkUrFIDFGGTXkIaUGV++0KIRUpA0lY4t5is0vJ9rQbh7CIQOKDcPXVFzv4rjKKORu
CUUo68h0h67eFplk2i5u/Jhe+9uweACxbK223gieeIkQ7ph+XSFLAmz0CbLiLUe7ICtPSeNJnas2
UF2dbPK/R2Tv/dBnuhXmsAztE8h9iHujLgEl0BRJ6X0zW9lFDxTKkXjgcjsZGVd+Xtt7g4IP0kch
uNBdo8ixobFEhDKbLCt13Y4nEcIYUdZhBDtyRB/G8n9F2EfZu2TmjEtYRVLRfOd6fr8irpzNzUFF
OjCKSVTucbLyq1ILawaMiHwBNljn/85pDphkS7IfZECf9uzqoxBbMm8I0aKwyR5PEIGDMuUvpKmf
vlBRXGo5YGaSBSzzyVIT47cVOSEma9V443oRiw9RzzhkBX2LdPNNsqkIZt5sP6/4y4BxHj5PqFdI
3lEcCljJaC80ibhxve0EvOMdgFzneXT0KlGELZVt55HniFBHCCB0+FNVDFqdHThagyB7dHeNFfMC
SqpuNYtCM3TsWi+YuhMbmYOVcpgUAOYNCHTB2We37EN48BaupxoGePzojT2SnIEKlhsm/jBNhiXQ
Ew4fU1B84RAcoFt2Q26gUuVst9pYdcRZSbDaAyiExxQq6qxQykRuvO1ptdrFjG/B15Of0K1sRNac
xIOCDktZ59nNNFSv5LnebTcJ0drWrEUEGLkFWiJq4RzMFRggcj1zjivlAbTc0tUht5dmttD3QSPB
RI3fZWbRNtkjUlzaU5rS3V2CFqRXmhIeALO2SV6SQmZlxAP7QKIIbq9JJ9M2ums2flGWlqmmlhqH
1Xx3SJEHtgBSPgiRFxh+MF/gvKL7Ux21IjSwGUgCBYzTDBfXQNkEFTt3tGyA96WNIkfTrmTpw4nW
y2Pm4GHU3BbSsAzz/L5tHKhkKeZBoetFr91g1CN/W29nGfw9j6p1AM91BzICQQwc3dLlI/LyR24E
VAKpWtME/kirHQ2AAZgANKnUZovTqPARDc+fiTi2UtsFfaFTonvttGGyrx0MgMc76hId7uM9kPzv
1M+L7dldeh2CxD75aVdKi8z5+stTxXOzQtfUQYt4fEh+aHF8RDbIkBcFZzPnjNY+++lRhg9i60st
BkFoiwlOKRGu/0hPIK3luy7BmPGtbWHzUOkFaZn7WzwSjYSJfTvm75jrUPxGC+FtKrATU5aMKKeH
okYuFSszacWPhNT1+xn895KRpu9aJxk78zjOZGj3vGnAYODr4OheU8Nc2Zb/nZyKw5DD7k1WCTbI
PzI6EZt78KJUf2uSPixvXJ/+qOEEEFQU8wF15oWR5CMfrAuL8KHwBIHlmipGCGGyXwUctgkUe42v
tBD1XgEWQvdUmeWOiLsNgUwVJjpGDxahqpjjvR/kkp7eRGVjOUd4d7gI28LbgWunv1iKKHUlaZ99
DbUSFSvgq7DaZOJTqcH4J6P57FQlHW2AtxLB4HQigax/x5ct+qs8ehfds8qp1BQoxHhhYgKlrqej
S4Lpghq4n/REBNO0YIKhHFbU8xa5p9YbJjAWExfDp2JJwx7lUZmGMtkjJPITCQudHhwyUhbzuz61
K9zrMa3Ud551P09E1V4A0EyGXARIlzCx4f5xNyzwtG9pGRGtAcEtJ0gS/IjSm5U1FayOsgvURDVw
NFbmBirsfqdD8rdvH8oMQa1bQ1K3GdmviVZD+DrX+hldzaeLY04NrTogsWum7uueBkjohrrF98Ur
nT5rSegBJbTclpsh0JQWgb0MwBtRqwFPvv7wcrLXKYgGJ6qB9UMkDqT0RRs2GsI2gWmqlAtcmk3x
NJOwRVlhtwyp1x13luOhq/lgnoQf500WRwpOhtslu2sxnGbBKUo6dgoFx/D/sbWGNr2eBVY6nX2D
4CybXhhAWgQ4boVuH07xClOSGbDyoCfSx+JINGOmDOHLJQ8uLkP53DPA6y1gRXYMeogaM8Zi7bZk
avUHIie1iM/T/zcXLkKHkjz0TiVJsv7A89gId2Oa5FiPb6WBpKX8SeHYlvPki4sMdZ8aG3ZQZF1L
JzbPAOxiUt6X8VzE10LwhRVCldKw4dBMvhW0qDGGR/pClZGbCWJdQNPGQgn3t3DgssRwlsybadbt
U4AnWWw5QBbWLBoaVMtZUukcEP3BWi8yaBHCMGF2vBE9VHFQ2FhaAooitBtp/atpoJdKs2KwCtoX
T86202cdR4HC62kzit1MYQEF0Hm9JhhcQBsmF8SVPksGPCW/8ihZ1p8/hc8pYyFK2caTzDGTg0ZG
dwtZ15mOYEW6GT4Amfkb7IimmOnsk8c52vFhZhC5IIPfMUFvAwofo+dsp+eyBNGrtLJFCSynl6Ow
7x8hoCbi928FOCBlfGLEeHY1f3qmSxbEHhSE9mdoqrnvQEaW7jcbHg5RDwQp0IJWOxOkkgdJ++DG
VTe9DhAuhA0Nhkx2n2Q5RNHCrvbMsU7CVpSKRhlkE1Q6KgwKeruVvv75YlQWRTtjbx7/JWMoZbXk
j7sml3CPZPpcSuZxOKiXYhw3px0cfwzqt4VJ7q5M2KQwLYI4bD66Zz+fkoKRWWp9XEYx/ET0b74N
itYkJcOMVSBfveBcADQAI/M/peaTObhFxquNSKinQ6VHRTeBG9/8sJRfVnEmgKeNK44spnw9KwAh
LA0H60SM4Xol/Najv/6hdqNxDlmsjYE7Vp9jy768U14BiGhvTBfKCt/ioP9BRat7+GIjNqdWDXDu
KE0q4V0oCLiYS6rnxRUSYrVGvrmbVjHxEenBZrWAGfnNsRl2MT2wy3+iT5ntgqb7bC+87jIXAZdC
RkjQSvIi8Ff0QG+6DxKkASkSK7NPRRbseYuYNRzCiJXkcXQ6yvoEPCMWtVyp3Iz1iXtv6FwDiNps
JEmLNEXrz/HR93+2fFHDtJQIeFmV+6AEV5kkaQHhD177V5IYslQXSkEP1Wg59J6oDkbCiNgIlJkF
6ZoEeQ6UL3J05u633eBzhcAjuNLTNuT4xzGeAXdwGhDh9Bv2gMZqKoORcw+MYoVFd8JHBIKn3Pcw
DZv/jzEypTA6mREm9nFkHQNC6n+qsJzp/c58JludtT+Mshw1pAGwd2pwoAWRk3jLjqEmYcFvsFkX
uR46sKwoYc0Q51CQSCN6RrI/dT0+9k7Mx7xAF3b1W4nxTuBoOB6sC7TGjlewCcs2AojgbrHE3uql
GD1xI6VpB86KBZSqxgVeS81AKv2CLW5+uD/dSg1CDHkIn+h5al47aopXdyfCTR4YJfZgaAjac6si
nmjst1shsxDD3nGpTqHcrGChEd/W2hou47+aYxpm7ds0KCb4uKCgnHCCobJbzGIq/L2SCiEe5D94
9fbiSdWzI2rNhUwT4Y5C77NR9xmb+Dk8GKPbJEOCyyNYXjGwmXyCTdzso+cTQd/GekTXNoOX9jUD
jHx2XKcYfCRX9M+QXnhYaqx0fESfZzJU/AQsmaDkBN9gXHlJkxO4EEMfOAedlCQpi5wYjqwn8959
22mVs8YI0W/vJLDbdTdBAWg7zPMzzoQ5jbQseP8eOlHigeVUmX3LINxUwV8oJ//IHLqXZUCx/Uwy
HQGWS6d9ek3P/xG9Q4JXVRlY359dn8sdh/dU3BZOhySiCFWzlGBan+5p9qnIKS+AcmN5rjJ8fjGK
DLioxnZcIRJBylyJJuZ0mb73pM+pa908Nao2DyFhZhBtUTjEk+tGFxGj+mQTcuVwDq91SHolTgzL
y27ttGHHcTvhXLF3Nz6s/WVImgjThZwdjt16UXtl7UuNQXxb7XprO6tSfXLnOAPUVYzwzV0WQB4h
PajjX+p7CrT7olKjZjaXr4xMjvzw9tI9EA7+9PrusE9GV2tvdV8x/PsmVGa2LsTlvHBcy/OmY8f/
hE4U7KWVcJkLrGCvEfXjLyPPn+XxRMIbCIDX0tlV/tmP7r9LT9PFGk4N9IM78DIwfET9v7TeJGxe
CqMoQeWBy9ec3EfBKUefFXit26fbk3dVEmOx4zhVuOp5YLmANgiN29OuSEtrby7whndG66Rt6Fgm
WXhCs3NDvY0G83V6yd+q9Wff+5juUpApOBZ6ertKfpvYgB73KwzTalAv1k2sMrA5BbJQ8UXjuV5I
kMStTf0a53tNCxOWrVl5zER2noqdywwGANwWSFS3JvFSuq/7sZfd2/zqrh3bwbyXCrKSZ/bMCFZk
qhw1A6FjyxRUVquDQs2lhr3RLCkohRroePIBWmilhsHQmiSw9TFErgP9sCpVcbrh3I0Wu22csYJt
G7aG4lLcESdqv8wBb4sZUubgI/Um/XDojr9qzdbmkof6T8uXD/Uk5LUGjSg0o2kwuR/dBk/TuQhb
WMfeWJmhD8PjyNypHx+qhtb0LVROVb/GIBYU7IbuKPIXi0ip1xpmVeAl61yL4NrQAUzaTGa6Qhdz
4b6Sn9GDcY8MAGNNrYnRjgk9oWVCkm8KOkO12F+VrJUjYzrGdRNnzzfx9urSpNGW3DQP1UNfUNBs
Qe7XYYL30DRGqVF3353JGXhATCYSy4dxa9VLG5WUtvcEcT6SQyt/Z9rYtLRuK1tqwBbKeZoxhgaC
bVrcwGtDVKQHPcV1U8KUyr03IofFRTDHInZZPvZFQo07wBg/d3wKEWEQZJbVHYf3agJqy97c+c30
6iuWoN0GGCYkJ+XoBQkoytU5jrs34WXWp/1a9vemcV4/ChbiBaNwPUvyBUpd8Rkewes7+YWrhqBK
8l7IkAl5K5/P7PIImw4+MNkIiUruZD4xgL2Q6UU+QBwTnWmu3UlQY64+Obc5f1FG9o0qP0FeQhag
ZrMhaqILUs9Pk6avIzJ1gaEDR+uZiIPRG6kop50/cQ7z/2R3K6sVOwsuGMB1qUtpjpvYW3GTHYQi
rJOTNHbGZtclGFslQLQM6R3F5z8HcXysKropxEfelP/u64VIcZ2sniLjaik6JwbWh7+ohBQiu1Re
J45d647W1jc9ltueacTLjc4lxmx9LzwKY3Oq5yt3loWckymUU1pHyhzj/F32w5fMag+VrkDEySN4
WvUEyvBpL/RDC7yLK989hSN22ZwiL/bcWPurhOJDI5lF3i9dNDsu71q8Nk1vDRWoNJ4N2FaFuKZv
3Uhd1nHsl+PMsUMD8fO7Vg98Qx9xUdoYYxnv30CEcTxshG8PAkpV8sGTkckXLfixVYNxluKD/NXu
vdcApZqA9Qt4PKmd/UEX3/Ju01OUplrIuI+ORltYyEhIf5P4+fHl5SsexlFOU+GInz+TvsNTQ+Eq
otEBWqlO3oWMvEIQ7CJOfwmhhZ7YIiiq5inRCjL1tmA7TpWBzx/pHnnOtpp9+M/wGVnJeG/85j/9
h2qIDC8hYMEgDKbHzULJ91jWM2HR733pe0IHdJP+3M7c7Z1IxaCGQ3J0/3fqINRkx1oxhK2rBzKs
+7GTlpdU/KjxjarC4EZgUsnjqrJdMY60tDrgW6CWlxwVX9jY0ZtIyO0X5BGNoGK08fjMbjFGdqK2
lsLFrQhDOpEZsIqG/xVGvAdeRtJ1y9JYMYxTe4HGIZUoShVdweTWaJw1UUxYzs8tnfzRUPzs9xEC
XncRXlYa625TKU8ViiU1yIfRLBwt8JkF0SdHUZusi2+uDptUgkTDhlOgJmlJalZZG5k7zM/r3erC
HazKLVJqL4HApzQRx5gx6qS5fgzH8JwMHOTtk/1xDC3C/y90Z5QP1rR+FIMDCEYVNPK0h60vG0kn
K2r3VMiFrov1I+5PcgXL1TcqVamZYfpfuzk4aPeib8TQIrWK+a1tkoVRrEUC3MlrxsstTHXtFBzT
Pl1zTTB0nh0FQZo7ot6TLb4vq6LKc7GEiiMcRFS5mmdgShR2XaLSkm8Mczur0xwmdDKpLXocJNIE
qJjNvAox2FtSrSBlEUsLSA0UXntLCb+8VSsxDb8Wy/dza5fXxbct6qlJ9737Tr1zRoYDtq7kUTZz
kcILaBoArygtwuHYs7FntwEgZGsmVxpOA0FUo7xIn9kCC9agw6PS05Y3uKVE/4ce+AO9JF3FvMN6
ziEa1PKct6PgbdU0cfaZsu4TxQs9LNZvHE6tIRmw7f/iQP9Vg0tiVIziek0bbml1FvSBpOhg+NKx
FWOO9Sik5J3kjToUg9gpuQ0IPoelVWecq9curlfwsC96/P3EVST1AmSLg05mLDOOmMr3uVm69sd9
x72kiK8G/c+9oaMsq/fXDVrgam+HTyuq1eJcC0TEeFA1AndEMsdX+F6Nb1NjxwfspxgKS941YHjG
5vAZKGl/pw1SgC40T1Dul3LXU8yV9fIf2O7DpLb6KEpflMcUI3R3siijwoFYPfR7vMAk1qu0H1xw
BEAsIFrw3Kto+80YCNdnuuBl6XPAkzHNJQ3A0DszzTXZ733Zlo8KVHAHUlFO1VfJGWXapP+lAVSs
E7DcIXq77iyFgyvzLbgE/xqPg9EOE9lSk6fr4LpL+jH6WNFsOH+qLSC8gZlr72IsaidTz31KToRw
5QWi32y3/yIQK2CaNKn9bzri/N/ZC16p0dcJ9wOm0lK2TNLdsUalqi/BPbKTn0fiLSHfB01YCWyW
6nwKDkIOMpJ2zowSePLss21vAge2LCWl0+DZMNVPywGRJPAC+XUIQNNHtgAGV/ugekwoUoFRBR5B
qe1WZNeY3ZnbsY1dYaCWS1dPn7IJYhDglsodveIe5VnFVoNj9fqVhh6X+GYxriqHgj7oE+pC843H
MpcaB0KeVLDeQicoV4GsONWeIedHwLJQDe5jvCdhFb8lIzo+mSOzbVJuGGM6jO3Ovy1aCCfSBMJf
xbzQqe92SUqCZNcT9k/upKQQ1ZLZ5+4d/KOmrGZLcVf7T8opscJKP6dqO8XX8uD3qPIxjOelKXpf
OW92zVNjF0jwuMMyxB/6Xz8fJ/JVqQrWYVH4DCCW3r7i8aKNRD8g00hp/Pm51l4SFFZ5MCyp+THv
SQtQtDbLn9/Ge3RvtBjQlQaJpMOKCqedRN+yS0r9SfPo7Jd6+0AS4Q9OA2VVLu4DX+DUzJ1gIgGT
6PbnR0ETHOabf6YfR+VJRKbSn/wI6TjDmoRpattgY1anDifIwqDYZP6jrKkXdta2hRmUthzQY5Gh
nueLJE9uT2YUAzKovXWbMRDrFcwjknr7j+dxC4k5c/SSsvhLWEN3rP9CbKpsYdGTZVL77FdEmxGG
JrdGOeJl2FgRMxtHUurxaT/FF4gkjbnqYQu26xyYU8hFZsG0GzQXYpu7nI+J7rTPMh+YFG9CQBMv
XuU3zD8D4p2cLrDj3R55ny/Rw5+zmVmzld+IPM1O1KvEWoKkq5jc5z065/SgMbaMFEtCCYiHjwA5
gFF6qXmlyFKQGqgUhm0fuTtOR9ZraUFmevY//fste02CAZquaK03g2NOF/76NJsil1fBqLjcz7RI
ULfgUo/g9GycoawNJvPF271FmiM++RDLe/8Gc7vplEZFnBYnINdbrH40/nNsnFodZn1T1+qysnEx
M9RrlK/GT2bxGl1pzRaNgyNCMEaBIFY/urCW1VxIRuhjDJZrok1qUzWbPIFUrFD8RigINrteK4NG
VagjVtM/m5F4lZNKciOXef7GC+j9V89mKrvhvG4HdgYCAn1qmcS+NIUGDWfxijg/bE/9GwyLDi7o
llCEDT8vawpU4GpSwyEJk5x+pTi2Wh0LqbFWukV397TKrjMGiaXk1FrnkUc8CBs1mVoFvrRPfftA
RCMHIucxS3w3TOvcdCjkJWbj9G9dAkMiiSki85STLyErD8pX9dogDEyWlHaTLuNISG2SOzWHSWsm
w//8MEhVJK3YaohNXgSvCUzs9bJ1R9Cx6AgA1887AD9hh1u3kjeoiTs/F3VhG72Wgap0wsmlOkBS
CnCQ0fnE+O3tvx/yF0AQybllfPy3HeHoM23AJmGr6rNxDf+esaSGk85jjbVZVbfnpoIsrEcusNNr
h9tnzkQxJyqjFzctVaVwy4Schim9JtRIj2iGDLwca6MwlNJoDr0R36NqEhh7xVj2GrpLQ0wgBDsm
Ay6nj9mYy/vjTmrWZxayvtU4gj8AzZ1QaiHT3dcFEKE1zpSbQ8S7yhs1a2IStLG/lTFJ2jUY+6EN
dqfcSUXHVhRfO8+FF+xWK+NouOrikLZGs4/Fc1QaV46uEqqViewDOHsZdWcb/2u5ixPEqjXD+I+q
LL5eUkWDp4/H81IDMTDZmCZmsVHRIr1PIOkznoZFUHidyGnhmFmclWXK6x3WU+Cy1EezD7AcqJ9P
MBNencLkhbSKDgqkY0sHPYVO+eikrzVU97E2qoDKLVixmIXKTcpltSDcYMxICyNO/146PJonI8x7
Kbol59Y26Q9vmrN7T4TbOdl/Bwh2mz4eAWgJnqtHthIMbWrcc5uFFV/vzNjNA0pMUmP/e8+u13Gg
XQv84owIskTWweyHOJZjvNJ4KAYK+Forf0YhOa81l2PeMa9AP1EbKRaXGDoo5IZZGSTjhx88dmUW
hMlXuDKTq+Yk0nQygiknLgvpL1gjBf6tBM85JvqQTtTHeICHO08nhBccTB2SffCgysSvPU0qnS/l
hYmFThNFb3Bic96r1w8wydDDHaOvUZaR14adB8yaVE6g+FOWFkjGsL8qIIN6+gKOof0d0lrwwq8u
inveOeF4CNbzmqViza7A0MBnoGQGIZgWRxvw6GZts++guzI/IBue7HGykDDYxIhDY0JHDnc4057v
wTTm6my3qQlG4vsDyahsgW42PFzqI6e93iQsMI7wShKpwRRlUp9BFvr7qmbzUnMMy5NtODiY2IMJ
QXgrLpNLaiugEBmiuxhnKZA2T2yZDbuOpPcBThq/uCJyq9UYITf1I3c5unndb7Y8mzBjy4iaCDRt
vU35mG0GHRTiCkN5huyYvOLuX6J+Lt1jVT+ZOxPLf8fACBfBHy4nxKy0kzf2ZtBrZ342H241NVzc
18PHQosTG+ic5K1OO52AR+7sELqwSEcSV7xzB79wtASkVWeaMULhNS0vGG1kcieaRG5OntzMywe4
cK5+C/XcS/PgCrF4yj7wYE6T00ymi15cU29jhEYXvMIP3DjYN1VGTm0mumz/ILT6k2zB5GXekVa/
6JU7vG/+nulyy1JZqNp5/aomgF40yHDqMg3x0Lo1mgHuuH36dWkPSGo+RpK/uJgAicqLOFL6efsp
3/By6t0rDQWKPVyUf19IBUqYBZ5vufKjx+vUDJ8bf95kjSAhEMtZ8KylNvW+EXf+EB1A9w+mLCrc
PV+0/UleLgf+od4SMRWqyZo558FP6iVZm82i9KX7QFTHEac1iUdQfdZYyzruIuk/87ow6rf2rfDN
xseko4ykyfuUCyxxEYWd3JRI7kQaRyY4aevYxsBGYteQwBW7XM5oHbvM8mr+vz0nVkgbpKpVHWAo
7XQIzfr102+jXUzy4EfdST0ll31AMSr9m+yJ4YYW4CC5XgBvnTAEMJwlgTvxpxcH4Rt15XOcndQE
THo4VWME1thQ1ucUqh2Ls2s4GjYMqIJwawmMH8UQjH7jiHyjjsUzfYMd/lfOm7l8LO239rB8gXv+
KQjCiMX/EsbmzDjgund8ZLWFDLk39/LW6pXViTkV3rBEISjzItoKuYnOjm79IS73YMKjVjuB7N0L
7ctcqYtzNyeAcorxFMXUqx7BS6gzlEoBMDf5S1pi35gyTDkLkVW6EdYM6XAHbBUi86SSEVMcdQzR
OhX+9bVNBb097oGKL6mDn0qWYAoBQk/d79ZFjVqA5xN20jUCHhQopbPAMJOXs7R7ni9JfBcZb/hO
I9X8ifZ8b9rChMlqgNuLhpiDBZr7nLbnHPPxOG8A0Q4I/lzQ1fgSyN4kWdPpmi5tDc3Nb+kEXczE
AbWRd5n+rYPIH2321c9CPqw+YCZl99guMoQpkerygiMJPm3oj4tWrQ9WC4tfyzFEvyElKrxUozgw
udQG6o8knKxkrm66AXF3Dce0rJ4ZH0u1qrRIfKalzbIrDNn45rQVnHS1twTuzUw5OAgeQlYQmsG9
espolmiQVaD9q8EZMekzLYSkWUOyYnoZt3/TzFZH2eKjGKK3rJEQhG/wbpAtfvTAFpAK+dF2l9tb
RCIJSUJcjvnXs2ewBEZdQkdLT00IvPvwFqB/5pgKQDh7AmMBhfbHlJAlyhJuUciGah7Xo7nulmlC
TtTgZbCQ0gFF3FTDxl+osWUsFtoKjU0jDp26ZQ8epH1MkOTZhreahyJXYrvsj9q4jDN8eJo3DRRR
h+1w14pn4SPFuOVn4sp9JHWg6LNy3PCfrEkLVUtiND3+PY0rzNClb+djKlQMgM6xWOfnqf8v9iox
lxXAjmpozGOvxBQJQqhDDL8q0iXMCetlRodRrEEGvlrNsAQ9pjFYKNLZiHmrK+VyX2u7USTWvJaF
D7p9TJI6cscCo3P9UgnURLyWzFdQhCfMUvsWLwQdStJGvVPbZfwBuJtGUpPByL5EeOuTgk2MDRu4
P8ZYBuos4HrYIqCfMZjkKnkIUtV8NfbmbQpU+IZm4JiAwpXWz81XmaQ26RoId7Cwh2ag0xc8kQbA
sktIqQQVVZRy+u53mqj1uFoz2QEqkkFvdLdqnTZPr/4q8pWKKgISaN0H3Lpgs+o6r1owNh5xM612
950pIkwVcoGS8YMpmsxeGXu9ETWmLrvQIvg1+AJ5jaKjmNuQbrcQm5FwhUjdzG5IhoXoAVaN9Epj
8OqMdTkl5e/x3Ypodixe87fRaXkokIuXE5EFuKJFbpYdqxQIrNmk9mIeQkl4FlMJIA+pIVOM8I+z
N1jIY9JLaw9uQFCdnGYaAA818T5U489JDI0TQDmqoQObYw4ArZOzC+RhTAuJhvE/qK0VSOmjYmYc
a62aCv74bVXPMbNMoSIXodnBx37gEkUmQoKJMXayiaMVuSv146qe8373S0BWej3VeB3KLEwwBbqz
lvRw8KkN0ZPVhUM9pMUaUjzXmKGuVXP7mEs5vRYs6Sh6xcbr6UZoWPasaHPwPVLEsJX5QoYbSMZr
0mRAUp3TYpIWNglExk8B4HCcrU0NWmiCtOEKm1x0XmA8DYPjDGAITtbt/ohzFnFQcaUlQdXq0XQy
6k8BGo10zlfUikZr9G7NSdHn7d/Raaj170yIrIwBsxAEJ7AHfNMeM21BwW9qijoK2PRnmiQX+kuO
642WtNqzsK4t1ezdzMUOLRE2IIRdCLAtXw4QkXGGXqsb6s/rrWxKWxUmh1zl7EuM/26o+WLETzlE
jBk4onVVYkdUwrKQI0RENlSzjWHyij9E/SOTfGBlGULahKefAN//qLBw+i3JKXq+w29E1OhLj6Sx
QfEPGWz3Z7jKFq+h2pwLKxS6lm8Nh21BbOCnq6gljjmEiHkubvpKEfRld7vGG9j7Ar3KSLufjdUm
/4q9WkQTERG3xaOH6odjO8x1EC49GY6T2RcfBZd1XDowNVing3FbwtLzLGDzUlvCG7o9SSSAKxFx
7KeWv8BqmWsSpfkfkYhKY3RIEpDJ1B8YjCuxUmEW1PSlqfuAZ6n3IkVElvfOQjBTq34ay9kR7XD+
bpWBzmRI6OUJYU/q8YGXyLQ8b/QclC4kXyQazmnzjVCJjhw/U3C8i5oG0XA0enxynUJltfAJCKwk
6hQ0vCCpyxn40eOoEKq8/3KW5UppKhmy88ueVQ/GZ8Roc8hbO3uMAy6XWkRfug2IQQciKZOW1Sim
CMXQvYPXXmVaCctlDGJaBZs8qS+Dd5JEvKvBXyW6yYJIocvznVRJ1xC7KX6ELJXKi6qEmKel7yx2
QzOWux7UpbIURFZyDQJa4n3L8LH2A+MiFt/M/pZ2BgjFLG7jFKNu2GUe9lZeypUuDM5OcWsZ8Nqf
trVXeFLyWCAVgc0cHwC6ngtfuh9bvdpEj7O8WKr5F5DIdBMM1x8bh9cK8rrgrpl41yhuJ5uLTvOh
/4IDnzg138Teq/TrVGYkZI9pbZZJ1lMSbVYhhj4uSAkZA5OXNgdNRPevysFKp6U5sEcZ/TxtKwQf
wBI7WAweFbnBgrcCXghzuuGFYQd4etTa8Q7rei9MsQRHO8+iPspCNAIAyI/uQt0EJukNWnwuLa7Z
rvVs7YrvIT1OMIH3rOSGEMG9vnedjmvmb9D1xvDMGUv7p7/NLhZGslFYTgtShbjZ/cdlCoc61m1w
6oUrK+7bi3ABZQOtpQcYWH7icbGdhQ8W5gDKLM23Io39aOzCq3oRL74KvyFaGNwxQqvIvnmV4fJY
UgLgB3dG0+KAJZG6fgfTzjaR4afzt/AwjdPHdDWLfTfxOaQnJzHq8/6A8FXpaMBjd9/mVmemXGYu
L8iQ95ESdshj5zLvadYHb1iht6casejpwpazO6iUhcLCHqZPkBeMmjChI9BlUN5zdWCQXqnAgGIQ
KcuSvzdk/hqk0yBMRkMz8rB5tpJe8UQURjpHSvo29aieQx4Voy23R/LNWU2j88b9FHpXz1GCxmdE
n4yHEXrrzEQg1wUIhQKfeGFyo2LOCgljVa4tiTz5YnD27Itn9oxR5fQqDz9cG07PtBlB+I2JbHlO
Shm2MyST7xm0JVnoEHBEtFwj7RMaiTvrx5iry3nBtxkLaM2E6Hb11cqPaOPs7tfvugsUGni3TnWY
XjlkzbYqNe2YY+K/wS8StDfhbuAN6bwLZLs64sMO/HAyOouwGykRTzWPBu3G1B9gUxDM/4qycslp
RwnMRppMqWXxwLU+LFHecM21K2m29zU1pKj5uCaMJj5VyQfISS210oCjeqFo46/o2AhbJzJl8fHB
KAozPrGd2CkNtiDhVjT3qVyMlmiBQ1wLqmhJor8NwBsE2ifvEF9SioXS0UpLVdaW/srFQHo5n6dD
jR9mK2cJP9EftNcbBqkMEQaqruLvSNJM9/s2h3WZddh/0WfoGzagafD+ENPVWYqY+/GtfVZZI9IL
TbyHl70q6tjCJSBc8JQKlC6SvX41mY7wI6g7f1Bna4BEn/Q34gfiASnqmFV4VR8FlfjTvBJHNwPt
+C8Z5EsYhk7agjPi1vlFJImbr4bbazuYPpMIx2FdLtvFMV7BVSAnJOZjwaGMUWe9Hbw7FQuFpHvf
OOqt0ebLJ+yaiWKZKDJkoUyxqQWcU0maluVOK2C8i5XwMcIAILPcMqDtYOQEpGr/+pNdzK2qRv5j
ncAbiIN2BZ69R/+l9DU7Q0vGN+E+MJ+Od20Q64lt5e+R5Z8GhO6MWB4m/ME9v3QNY7Hsk9wY85VD
9hlZuKGcPNazdmg6RPUr/CP1r9bHb+bYxIUFFny3qwQRVcfSUkUeY5HK72IYbRSFV7NP+7X3U84b
pjJkhSEnEY2vvSXIG0YAB9rODF4Hjuz7gQJMqZyFiYuajE2gMOU0WX9a9g0fb2yC9DKO19cT2juM
DZrb5RFTQNugt2a2uoTl9yJNbS070lEbVj3sAv52L9EnMwVbHRlbTi1CRSsUX22yDa6J9pD06Z9p
+joYbWpx3H7mNW5YGZCx1OINo0v9Tu5Vktz//tbflXc7GxMfY4IA4tcUiQlXoArp8hXIhIl4BYyf
SoU++MQXT7zPgtfPb079qdku21L82XtwZQVo2AhiMoN+7+Rhi4/3amEgvYAdSjg87Whd4FPNMM3Z
Xa4huyVvjZ/U5yxfBDVuGUBCq4mpdc0xpMcQBjp6DvRUjCDdvn6VY0yajV9tr64Fn333EDO+XeJ8
VjVcupGyixipUcwW8OYYnMMBNZmLaVe0S0+63PTLt493a23Rl6Oa7qwWo8QBAzIouH7SWtWLGdwz
GGhfnQ6ukynpHWK0/a2O4dFkVCzb966ddD6WGZ1MvcXObIbphmUdQcr9tz6XaNP6mGWxS5Gyjsdk
eSa8I4SXKs8ZdZgjNsnoTyT5BDf7R3kqqJkVyTwblYGkS63SEG0BvyKN8O5jgctXE8UTbPshHEz5
j+SiwdVk3+3XTIQv/sXYCE+3xc5ZzGvF/Dtpo29UjoLFsOJEwQh99iOXim/vBdQ++RVMimOkbewq
Bxoixr9L7fJ/HW49XN5WOhNUmF9qS4cKOM3IZXbj5dg6Cv4oQNX7wtuQIpqntGacr6XTbdDMKyNm
I7YkSlCZNFARDDYk9uLB1r34K3MoFwGgfqni+rDGxldYzIOvpNWvQdXD5tN134q1zigc1j4XpWuY
vV2+x4RjC2EZDbQr6cpPUB+HsWZ5p1LGDOdbQWJB6zgUHpiNYTCz9eXQDFpIP58BA8tj4lYD2Zdn
J4Ey71P7CH5F1XV881xDXqXnbqpinqkB5EKWEtJURzMuxys+ISvxfSjQR+Rc4aNtRaMdudzdeimC
sSJQVHAkvBGszQQhE58YMtxrmNMQ18F5wvzmcKpNR2tI4AzNdDqBBq2RAX2Ea0CylBKkKuC1OTSJ
DHCPniIYVGrA39XGrIm/tOJGe0FyNgjrNWr1M9uVRQK+6dgTogcpr2kGZnZn1ozbEfqu6MSTqtjr
wNubA3liJdrwkrXayyjsmGSDlh+FePb1CxBu8yRqUaNcFLmVs3u9frLnhxDSmryY9PrZaNOGFHbW
eSOymQ1xPQ62U5VTsMOE/qJN6vLMTHtRJL6QvgwMMy6TmozAnq+eBDrT8ZmtCJcjILYi3Zq64I7J
jrbh/OIlNJxmVpWGmytoLwrBQtnICbGaUZE08vFRTv2nugkSslSlG+0EwII6EM8oDvjEOLJVfQPJ
4jAcZi9dPG9KEDnbxw5Dr9tOPgdhncNXnkiBR4XE3aE5BSYkWU6JJb3TjNGsA+15+7lptUfoMrSl
Ml6PW3JdNMfeusBMWHDtrYykni0WPA6cCSdyUi5cj0r3TruIhagW3Ok7jt65zp6+QGtKEOSO1R9a
2oR7VzJ85ctIOStAV6oWddtjn2MkDAqdsIMPg7gRJAIuItk4GTnK8tRQE6D0+UxmvQ+K2Q3TEPU6
a7W5QUvBe+FHzi9fiysoPM+vj9lLBZGPkqsLj6RE9iQ+AWPvD0AEEHFSgBME12ud6QEO4mwtKwtS
p9mdLX3TmFtPBtxobuwgCB5BbysjGaU2QgIw///2hmEjTCJxRFQl+L0tWQ6yDDjv4jZACm0L4SHu
AsKOkaeYPcbKd9Gw/+nDrKN9SAz+f4U9RId5uj/QgWFO+Hxfbp9y0hwKWcoyBhANC0MvHmzuhNxO
VSqy6BlKB5/yc2X5oBSEViyNYup0nDyKaV4HTTN9SM/L4zeLvhirMicCzLr1LowwNAxIED4lgxqy
uuaDWBp6MXGn4DL88bkzD2RMoqN/7KwOLEdvuGeZL7TI3/kduAQeAU7BiORWYeUi8Vr3KaOjXjVN
qH3nhS2oxpBEq/ZxMrZO9oOfrr6Lf2woxXP3r71eoCnqsdA7kUGI21KPP7dlS1VjEO7v8kcvt3Ms
yl19bmKWa7qMiU34x5aY5bylFwLjlbU+3jCEw9P+LTVv7AT7B/AigVDv16JhfisiMTMnshrxH6oc
TfEPCjFiSrxcpCHxR5mlZr+8/ZSnLArKU4rgFU1oOSZzGxAU9cpTr8N1RdKub7bzkYto3mtmUlfJ
JHMGwpQPBIW02IU5UzoD2Ma9yOFotRvhgP/gbJRENzLzj9U5jXUII2hcQOQWUM0CdWEij1DerTmf
vXEL/7KEPTY1XNhfhabv4CpY7fQOTajXrx5obI5wDb/1SZimn4CrEOKP/vHruVnYGPYpQGpx5vi1
qpzrEdwZICE6xMMsfomjjgtVUYjnXoJeHrudhVIWourccZtO5xf/nLzpnOzuyr+jPHI9VId0oH+1
s/WZ7s+832frq+thbEcGD/APNZyXZZ547BrCsGrQXdcNSjWogLy95oW17stcZgEBV19BajFeRpDt
OKYngCaR8gKuFlxBO3SbjbjO8dcyPhOHAZmSeigMqadlGCSnHIsIVfbHwcSmopp1HBGtDtz+xInX
SQdSzZ2OuCYMuyRMdHgupMWv/7+H5E+nHMT3e0CtlfAiLacjBvdkHeW1592zcZBQWQ7k6eE6hWiA
8ltRUIO9ot0iZ1nACt+Ezo2Y62rNp0uDLfrdU7LfGp81T3/bdkavgochx8gOnibxrIYWsMlMSfCG
oYFXDSuTBey/nBV7uly9PTItr0v2inxhc+a3vbZiWOwlbPO77ATDYI/8vIobjYFXRQE2U5lemnhk
SFm9ey9oI2Da1Y94KqiS75TCCPrhiz1TizAQQGFkHKXNJHJvYeypwNh2yqNXCu1/W6fG6fCNs9TJ
9IGuxTIPWgvY9on0KV5Sa1z6jPdmu2xDu2MMtLa+sHajuFY3PWMW1H/FmxZMkRQsA95MNwGnX16o
21WiqHWRRrq0M1NMyyBKXVyuZFp2V/Hh+1DMYiItII/PUEg8wFy01QUC3rvOx3Y1Bs5CHSgDZBLX
XO/fhqm0iAikhGqaISbPvjLc3MPtdf5LBlHc8YcJSN0oecF9565cTzjUMkoCxajwj4KdLbmr5SoO
qYnX4clhaScSPBQAghPTLRgs60kwT44vu0adB5JkVM2mXlQ3M9CVszOrZ0ykxv5KnNklPjiLLkGt
Ui15TG7uhihgBuXQ0aneZ7YXkwSNKA2u1NxvABELCQAZjAlatNA6b/Ke1Aj2jXcw8swJXtp8txJo
rNR6yjcew46iURRqh2hDFuL8x68Cx+/Fi7V+/u5WSqf19rAOtMsFT0d+NpIIwmA+LrIRHT6hUl2x
ZA9HIu7leDISEa4Pmsc+sZHN9Oso6Lc2ka2rKcOfmcgLcNi0qYqwxBA/dz4PFNltZQF2E1bp2A0z
zkE/QEZH5/v7rm3ldhicoXEmzizyD2gTO1snvtrOs9eEVTxb9JUXSNfsjkQD7iQjI7NesZ3GiIRt
ehCrYQa8SfmmB1tRn4MLUjgsdZcSeOz4Uv+dh/x43/ihPI7UGMQh/vz2K3l+ZgFmTRIjbhJvHdEy
EBKrE+NagqsTpxKKJDHK3W/f+QTcSIX/bXsBeERm6SSm9C3gyYSDIvLBvOIsf1Zuq8dHADBTaZHk
ZotjYaJmW0uzZ/02I/AEmEA8Bh95yh9tJ/ZyWgfDy228uvaBBNNR7Q0dJluHtAKIwxqXRc5mo7iC
iUooEHT/UwcUDiz5x4fC5Pe3qFPSqkFcF+cksNOEx7qBgS2mPEwE8BW5BI9zaHTC9nPXw2zY+K5s
++6vfAWQgsYJwj9jaeQglzibi0b0xilEA57PJhzVS7C/6N/KIbRKsg1x8vb8ILs7WAr6tSsfGg7v
oOCafxUJbeZFb9YCqLpUBPP26mOVnsgsqoswj52q47xKK6LAMpu6M16HssqFn261P9RWSE8QUUPP
2H93r9LKniGdzNDbtSibTI1Wrj1WMDUkEW0da+Ml3LH3MMLUGi7/ZgHfcGsP3U9ITdB7fm/diF/b
/5M/SPEjKmvbDbnrF7OIBXx+kKJbZX/f4Teu7keG6bvUdX9I9ocvJG0WbbEtfvtp/4chn14g4dVz
+KtLj+tv4uTP9t9p7ghu4pkQcd8YJLTG1u1mo4Js/K6YMp1mWsmqGJjHo/pDamNbaQJT/E1nclc9
dwip2D70nKSMEwIuX0AKr/igHgmTL4JzA4QqfhU4ej5a6jB81c69Ul1rgBNTS32c1tqdhL3Y8oID
gZr3pukyfPcEKaYQF2qFgSIm7zyRIIdaGF/C8rOf5fMXo2rvWrZeX90DIZI5GZQk3g07vlNyYRmL
s9idcg3tEZ2QbGGhviU712DLIHh9YP3FRuL4LhWe9u4alir7GqUA+vAgubmBPcWiRJo1SXysB4PA
D7qrM5HNEyw0EtD4Hs3j1cwQunVLSuUFJxNr3Qv2AJn0r8CrEX8zg29f5G3DYvgnDr4xuxEwDwfz
S9wjF/Gr2K30xLAHV7Ij8GPF2SAebw2hffOLRtBjjESlS1+N8wsFlDjNKWHrRqjqTXRRrnB/3Lky
uc/vdRLjuiTORXOOPRCM3gynASeeWkPFalVQqLmfATAuu9XaX78Tdhyf9SB5NLHRyITFF7eyWowx
lWZPXP1wwcmWZiV86H8CDPNVyXvkhtHXb5ZvNvj7IiQUqrFUjRa2+yxM5YKx1MUn4vUE7Yv1cgnY
kWrk6mKdNevXZcnbRAMjbRIcDSM23dF6Wco5yg04f4BFxCIjqkHCxCAKmRUf6lVjG1o5aqPd70L+
RXLZsoeRkIJX9/SGRJwCqm6fUH862AXRJjNEBXOR9Inty028tC5+q/2ts1H4mN5+sOITw5v4Rq/Z
2Ylj7ajPQ7RnxBx4fIRpLBC4gaXqzMkCfrVYPCuj8o706WWO75A+4hlDy/6ybmdRJ91bRKgx7TVw
lXgc7Ixzq2YSGpVmf6KFC/eCOj/asIPJwrM23skiT1yGwprU+kP1vvAE2I1ABKqo2BmetYrD+WJD
QZPvpsnmUCjH5PB05RzQS7Ezc8EH8hfx1Duqg8H1yikyZn+a2A2KtE6fGCnZUOzavMAjBaI9VUp0
mHicz6TJl5DiBW/1JX+zYW7YGFB333UVSjPrbpSzTiPjd6x6yy0+HPzUlj+r+XLYW7e2Gnx6q6BE
tcQz7FPu5OOGFtTiPg+gtnvemb94/LzLOnlZttxmGKYmr87PnjlAcaRIcnWYBw1337p8/TqGAGBg
5tps3WVPZQpSvh3MEj/Es6lWH8Nx7wAihPfXWOvKcZMaNNURBERZAQGXLE3cLOphc3hIP4HOONPe
0sIsljeg59u33RFpqFw+WxwyvLH4hg1QLQGj3QwANPKICsiZtnZa0qVmwYPafBppw5OK2K2c/9ja
KCj8Y1mF/3L5dzLUC2bll7bKENg2fCu5K9o8HAM0nwlqBzl4+/vaBu+0zljBIL0KLsrH6knjrkX1
MWXJ1v+FzWUDUcL0PmRz124bZGr3wnkDmMqFyL7NV/aYkWRpwO6ZF4m4Qp+Xc4U3MreuqtOzVuXB
tG6kExOlYWmZFE8Tpj9u1k5goWMbNOrnoxSGe5yX+WdwhqzCAZd9TUHzm6UWTI5Xoxj/slC2Bbme
0Sea7B4X4NSGHXLstrt3wTMiYexPbSeAS43enl2cG3uPxf0R9FM9cMmw7DaQnHsmZhDeDcKQte8H
/M9+Y0Ig3gpid3wkTqzmzc20lEahNAzViuPm5e8cd4cfdlY0BPFDmtCmDEYHpkorT+8xYHJNJSZk
aFTH8E0LRzDRRW8uCp8gADM5eDmXw0Vpw8i3IVjQEpY9wgeUYYBFiJocXMQINU/NKl2GmbaJy/Rp
kVwivHbJZfW3jInjeTXfGyvlBnM5RJ4SVECb926I98LXIDlh39up5PgTurHqnXcxPCkMp/j2lrcG
uSzRJqzJ9CdZnQAI52/5xNGPNnSwtEtCpCfuSHryRwUOGBWvrxzyKR5cy2PQscK4PTScJj+y1lqL
zSQDncVxbJIqRd0RK2t85bembjikVK8k4y0je9DRfHmK8fpmDR8ZBGdhVZ6LCMHgk3HIRxEb6TPQ
Zd2xTKxwHpIz4hzLp1ke6qV56yoBuqodibJU0uN3c57bgqi0qpAhU1Lsbo1pMgUMXtvIdyM48Crn
U+VwTxCpU81hv9j0Y8FsEzx42sKWW94PS1zPtwsxxzYhI7poZd0vH8o6YbhE0/f8OtoNcAlPSELd
Q98Vbi4Hu6yzm48MxIyD+2Gsea/0RYQvwx9jgNKGCTzWyz/B6KDnBRmwHNYkieDgLIK2XswyuhhC
PdMgxybkmzSNf5i+EinauEWBD+HBoECgjE4gnFfLTA3NbDhJoErKBBJ7OMK+iS9NRoG6aZVzrscz
rbzGjpZSi8Zld9BfhgZt6sA1zlFLCi5H/O+1U/zkOkX93zAFId96Ej2JmcfwemErUHlOBhkAGRT7
AtU2PGjqiYFh3XFe5/J1p+bmKgHe2egPSWn3KI0jKaTulhiIl2wD9dgEj+pLajzy09VG4IVEcYEn
yej8IGBapsgA9VpZ1uJO2umFB2hQr3w3DPqLAeVs9I6Y7Ad105GM8bhxAydowWxLpl0nhldHhSe/
+grPzAg/LziJhZCI6ZhyKz6//A1HoWH8Ex68Hnj2x5Eo5n7tFVXXuKWpTFBRAz4Frcojtd1C1Fcr
BJMa3/EgCEjN5NuogL1gf9+8J/PLB08llsGcZIoNCrBI1ZFrRJwtkSmIgGH5+9EAUN/H42QBKgEk
H+fdGZwjDv7BFQQJvc70fUnsJt6kjLZGETAvlzwAQ7ucj3FS7920AfcoSvAlS3tGwLK/kmMq0ffC
BXXl07/lkNenXoAsxRwMiCXm9ZjsJtozDkwqyePVs59creUwoaO1EHGWNTza5nlYNEUtsTXk/ALn
CmYt3JvxqLYuVZtTaUcuU/20A/tP6jz2a8e3EZW/1wY80lu5mzdio3JGUmkTvcjH05K4BWERs0e1
giNCMdf0I5yHPC/s8rUqQhZbj2Flls6li7CzTnGcT64Caw2K13KsI+L8Vwq1E6gFYQS/7bmJz7Jn
VXT0/WF2ZseY7AzodDOEWaWC+gjzpgm7IbPXPrTk5+e02k2D7enpF4xk5BQfcZ56QrlwXb4jhnqq
6hTlDbMe7hjOfrH5sqN9IdFWPJDOis5FRJs6p8hMYUYhD2yp4WZkaCzXc0t2kcE5EkZTmN5/Msuw
69dy9HhNu50y+2thTduBV0SI4Eh1LCVyLlewfpN4La613iLA1Zb/Colq6myqYKnqyVITXg5If6un
ueMSp5HC0yb0s90b8ktIHXAsYgiCxpdyVPY4n4aMRGWwx62rjqFgLxaAzEoCM0PEP4eDvTanZlYq
NDtrH2AtuVW8KkrcAcSVBub7qEMltzdg0UA05rjNTHqy86owFBvrlue1enTJjp5fo+eyOYvm3tmV
hbRvBwFRH68e0aifQ+MlTePIuTO31yP07c7OwIWo704dAgVNbgYlOQXy40MxZD0K0bxJVlV5mrEl
BC3MqlruSrKLNh+BI3ynNACPZxFZycfjxBusJVkldWDMxfev7Pl9JekAF51CTKfZtxG+ytsinjbk
hbEDj2Whdov5HbNIMjMJE428EtqcFBC8pndJ2EBAQIdIQAsiSTbsRShKdEhNDc6lQA78Me2oboJc
10MgY/vNRcPuBd+v43hr3q7aAsNcf6M5s2rPdU4cRac0F1Ajci0CYB8T9GQZmzkgZzEByLh9NZdm
sD3AEdtN3lporBjbifA9xO+INvGvJNIivAXg2TA/tIK2+rcjEEUVG0gfvovu2K5CcAw/muQpr9tB
6bwhZ053lNuO8TxxFqXySAWT5mh0BcwOKhC3ikyJmuDEBI6nPim3D99DB/4GkgnpU0VBUnBvuNyF
D1i9U+wXpLUvCmNlDv9yTi9MOhnCXomjv4zKe6Inz+5yamLRlAZSAn4313I8TIYkeEkYco0t/IGn
t4yAz+1XBJdVJkRGiV58K+FsEadyuIMlWYG3VL4nigx6ptqlaUjk/GfTdd2UIC2qycnra66ZH6jT
zoYXE9YYAZ0fFWd9DK4u/tUg5Tf+Z8zUhLQfqoY6XrxIb0FeGKIVPPqWVdJQjFnL+yl79b911Lq/
CV0orBIWahQfV2xcKxmgE4QG0Q6IbixHt+xyDQdSA7cbk1nxMD6WOsdy4mn73tl47fvo5SB7HReA
nVssn9GDt3mFN/kT0PJYIKF3eAWdWYJ5LnLNTXX8TnX+W5w57xZFebSaIg6QXKcAlhl8X2NO4nZ1
sIW/s7krxQZSyTS8fNACUSl7CUCcpPJopuK7z7T9dT+lBjyKTDpQB/lV7In1Ah4Y61+1B3py1jNi
YfLW7CW4sIV04zIVAb72doBqmuQRyT4T5ui5z2CV95PSFIl9m4UIocw4qPRDd3zDzCCanSwr0SD3
lOS1HItbgoPuOUotQs5iCbEAq9hHn6llFfML7OLP9b0YEMstiXWpDDQJLAsSiriwUwFFZqewzcr9
Pr5omIg0YZop1ZG2x2+NiSGpSpONyO3OzWTsZym6ctWaYdQqaVxct8OLu7j70vTj4Vb7BtV6KG+s
hS5/G6Bjya2KCitHGn+iVrgtOtRoHEca4Sjl1u6S+m29ZHS8RQG6dNI4zqY9qpzn51TRRlZdHrbQ
aBa4DNM2JO8VIzNjLt8XPQkuJ3Cilf38T9YAGTF5q/PfVaICgxH4cSTwg+4C9uL+6eLBP/DpSGNr
65sssiLoED/x1wwHVDLkJfwU4RosnGznrDRG/CxKqNVcyb1KmVosTZpEvLV/2sQwoNIbTYKaStrh
4kJggr7E0IOl1iGi+HbykYYztSaqqhnPC57hj0CBAWFtKGQ93F9GDH/8oiE8LDsbVSzs6UTJS4DS
qcC6SRfUjBZAXykG1UUMtdsuypu2wLSvCSYdcg0a0z6PkCpomqOiJTZJPGfFeIKkI0tuhFY45Nz2
sL3bPrBCGfvzQzbsoqcT4ZCi5vUfzvZKNSDdoknPa8PpAVhDrYjHycRQRidsYLHHxTNy7edT4Zi8
ZvbFdizJSBBfWuGsKaYcQZPxCAejfcjbvMdVCGWhwOLrXckc5+suADCZ0zZD9cqq5h8No7HXB12w
ZpphSTTFDAeY1v14IAxVrz5VP4+cgn8n+x5c2DF/3K9XZmXaa2i3Aqv1q8yRCeQpydQlQcJoNOCz
APH+S8mKKIQHcPZ/qaC3L0Qsv2ovuaCgxKIACSDI9iUEpu6aOoY2+NA2BmABfirtp2MJXJYC+Jfx
+Ox/4BYEfiASImEPcjbyBTt9PZc78GrT3k5WsAK6RdXSNRJIAuhBehPO/PsHWUj+OvyoiOAPvICz
7VW8a2vj6/Ycw6gnAbxYVsNziM/j+2SnKB5BxxSigXoe4GbA/06oauSEd1TlPfK5D8p7Tv7Oae+h
vFRAoayBVzXNve6zcX+2q7hK5r0IwCeiimezsxT3xpTL3xJblJpd6DE+oUDOWX8bal6VXnxcd3jQ
85VJA3wUUHXWlwLI3YyIdANqpgzz9r6ousHa4F0EIEqos4+VrsI7t79JBlcXDl+W4VYStRAP4YiN
pN5vxGnnrUF1zqkHRAR+G7zXb//la5pKQ81GMzqgpySn6/4DFgvccljnnC6IlxH9NedzAH54onaT
rfTckf78h+7Liy6Aonz9U1ULS7S95hsoUAIc6H9IpGwyOh6KN/1/t1YnAXZ32rZw1B8ssdVXeUXC
k8TeAJ5h1Ovd4Ok/O9pn69L3PG3x89G+mgfpwuJKICscne9alBaXSZ+touz8Tz90OQgxl2hr1cj9
11p6cJ6VPyYs+AJe0yj6PWpLGGzcLaum3nkziFRzKCo1PEyVyKFp/MqbHIysYPdcLg9LEZyfBZlQ
YlMgwhGifWOeXXChGrSTGuzTzo5rOmTl1fUcgzBdrp8dhgLUbvIyHg/q/nvsK/BZz5RiH3u+7Jp8
g8qFb2kqleCymMx726V18UlV8kUpKaeuGjTYMNllR8ASgb3MJTKFQ/nsHmdROgbvQwbIgVqXIR0o
aFdPWgHitpr/ioCLz5Jj30OdaztBrxAulicN8rNd4ij1KrkvxsPH2VsuTmJ+rVk7aWevM/JAs6sd
upRs+G+mp/zFx62clzZaQGumOuLPdK22MJ64U92mrM+9P5juavzTFqUWukCs9vpszjm6jVQtPZlr
BtnVMqS3VDIZTGVVQLzMdA3V5FRU1dDzawGS20V4xWA/HWe+6DfssIX1X+YOESW+YjcIfr1DHVbq
/3sBxzh29WCQalX32Tgf783cyyM62Cy3XgWNqShJG4IcUnv9dalnKSRBByRJK8y825YJpNsuv/5/
vqRnagi/Om8xJ0YR95jJs+QydJFcC9s+fbvP1AZiboEOz+7oh/ypBYUp8M1hJ9LzYkj+epyZyFhj
cYbqZsYs7SyILTNps7clkkhjoId1aLF/Nx3FytUZ79JqBW1uV5FQWHyUhnzsiaKn54hnOrPTDJLc
wS9WFviP4SYo9DspeIHsHP+wsP6ZT5EMTovBAmK/q3faAzObDZg2ZEKz+F3KGiJERBbkMCBTLW4o
svO5Ky89Gw+BqgPcGqBA1gv9IESjuk37Vegc7HlKUmGuLsTMA0ZyCDOgaNx+ACJySEer/hVuOkJ+
OaiBCZPKLEaUWWF94BZucM+znaEnRU42VtAMgy9n/dE2YOoKOi98yTQeM1n3PmvPvMfCjhMDw8xD
zOqH0zdrw7UHXQf6X1qtyIZwdL6yVaGLDUlUQJECUDLU0t1stMfZCUTPKvcmXl3C5ATN8ZZmLTJw
XBNbnWuKYEv7flFzrPqRpz917rHqO3mtS7Hp7DbRXHF9eYob8e7LdXZ5XnfnKEUS5pdeVtFSWUWI
X+i/0lrqe6Uw9RY1Hboxvmx896at/JZapOqC0IVDeTsrjXGO9r9P5YKZ8FZLqMc4sEZBKUfnSxEh
rpFtN6IF9rtMfa9sIgfNASZBgWqX4ZE6s6OuWKDpnMgE0vRwrfG08NEdw7SNYj+E3JfCnwrOebTk
P+Yk+JnGRCQwniLbgVIhjlMPTQ4l7sdCZLyxqn0bGaC34+devqlzPvWI3AYt00f5OdGjf12ax2n9
jULVjuY6F4GoIxSqAwQwadXwc5Yct1fKTcmCerwwhlQUKUqkOiudbGKcRsvmxnlQv+gsNcwhhDU0
hrqQXp0hhVFRJJbK4fuo/biojDTS0MJpq99Vk2u5XENz42Ibz54F8YE6dqB9VMxoGhU+jXQKYD6F
jzfd3pH76zdqA52i2TeFurHnIqwNGrBiJrUwV8owB9D9r3gHDsVZQ7qnZ75pMZyKdbpPzPouKDRK
eGJ7nl32IkvNOCCRma2Fi6/1w6enx6Seooqo/EXBQNo9z2xBP2JYmd3hWmu2AwEYHFcU5BP5Qap2
4yB1Fhb9r6wGYv4qvtQfmAMsKMN0Mxjf465nykMe9BV36HNoy/IIZCfJKp/PY6rXTgL91axsVPxj
brUaG12XJbVn1Gk4IxsaP3OtngSdJsWVYyesoJ5Em5Jt2VEzx0Ytub/Kychd+u5tT1CSl9V8OEwG
9ZySh+gMwkFD/tc+c9F9h58HWoBN8BmghSJbBuC2uBcEr6TV9txl51DzdBlzPFaMNcyL8jM4qPNi
OhtqH9wFRH1EjWxquu02K3HO3e/+VWQusRQGXlpyneUNfWYKFQ/cTo+VVjniq82aI/QyQZPRF0g3
QADAobCsLsn1vA9gwZCh6Bud5y9DMb30+Si4sMSsAX22h/d9BHzJTnydmWo3e11K1o3IP3yerPq5
2JEX49GKJwoljrf365LNSB0pNm6IEL4pa3q/cU59xsgTTq6CJsVV7ro+UmOma6r63rWaExR6/5vF
Qb9/FZxoYO8/E3w105+5mzaJ+2/DT1GMgE07MEpHYQH+V57KXazkHA2RZi50RIIo7MWLWrh8XJvi
iKXcUZZNuZkVk9Pwyx15/jsnuj8znM+ivWITfL0Bs5Wd2cW0O6RJRyYYOVpvawu+X90GMkia7Gub
rzpmaT98uZZhy7WzMm7YamP6Oa8o8oTDG2fVJ+Cj+jjx1jU/Eu8p0PYuskepY0nS+91o0f+oGRJs
oYOwz5+X0aK+mxBMAwna4UskOYRCt9Pklnqwa9MC0Syejq4sz2xwJwrn2ybjKWUW+PO3zKvMVvXt
NYJexWOatLv23eaT9kpdcj40supt9clm2/qDMg5efDKIyCJXknTiOf/y14+QdQTaG5B1OEkJ8j2q
GsT1kLI9UIuMgRWe54iOP1i0DJ1ZEE7apkzACy+6H5lIzdRtZhAufnp2P/dQ2wzj4+wFAIGoZxKt
ox00uYV60kpH3O1O7W22t5DzREO/8Ci+QTCDDtTvSewpBGhZVXXUG0nzJcem7bGy4QDvrCXAYeRw
VAkQXpUAM/Qe0PISQKYP4nQTsy2d6qMyervumO/4H0FNwOD49hKRKTJNSxAAfLmQs41HeVBFmArW
VmCWhhPpwuUvwT/1jvovd+HucI3yamXm/SobC5p785AwNf7656gZM7NTpDJCu0Vdrf6fx47zSKxa
bM7VyF5DJKkpe75dZ3nFql1XzCj1uT5iNEXE5heaa+5Y9hKRWqA0fUtX/MdKnusEflC02Wac1XvA
hcfO1ryJhm591pyaP4wt9wBUPoXD54HR0/Njge9XrLdkbb+X3XaNy1h9n+o6/QISqH5tbklTumnH
YJrcrMs/3BtWtqAIaS1Dx0XD7Xu4HVT6PzLIMojXmL5/ekGk8nlDKoQIMqzNeZZybIxgsVrm6q6V
XpGhsgeZQT37Wp6lCMEkY86cPRFVgeTNKYSEf2WXPM0PmiJWSkn2FLTAq0oSOID6VHYtGrXjanMh
BnL3OWol4cTEsCO70EnTGagY5yytI78vKyP7F6rm3JzTUcDw9EMpokeAoauo9cB9Z0C3wfPLxhn8
wsIiOKw1CEhIQtW10hPrrPKO0e2uHdENQiU6mA6pYWtmqADIeBVsQEuLg+r7AuEfXS18P6XoAe8R
Tvp6xCzr2Qt8qgZTVWhMe4EDU4S7qe8rioP/3Hg3lQw+oEyf0V9QdRZrmsY9iOGK8jn7TdUgE9t4
j9DLuLnPVvRoX/8zcQ0BJBF730UBjsf0IBzw20yMKbxUe/4AHlQPTncTtPAPFJ2yf7FnwA3Ri7UA
zZOnOnV0i4nAwPxb7r+UFqvmjbV6s9cdm124pNXlmX2MGIlEmmgILxQzigrPd1y1NcZyKkczaoAF
g+qQ1xQyTiYyFMAUebLto7BMpCTZ99gbvMzpYxDByCSjteIHSooWo58NdS4+LmBocbcMfI+llrYE
Dw1rYLMQVG/qUGzlrvYSjBGFVEZnaLxPSv7Z8AprMCb3L04KidjWa1+axyIcoN+njUFpzfa5fDoj
0Qf3oiNvelEUl7Tzgj1Pd3s0gFJ2fKfY2z2iMsWt1pWhy87CBT1cC57/LezMhmRi3SkIipPOVhvp
qMLzkuJFMtB+HuZYsBvPL89VyFG86/tR+5rwsRecn2OOkKZ6E4NYxDaRI4RKBRph/k5Bs0rHhXgT
OYvX1lDtuuRqi+W35y1YrrUxB4+shAp67o2VagF/fFIuFDknbAxT4etAJBdVxA17AgMpmC2aRrfr
C3HNpYujQTlJEwqluVPUYEK/kKtJIc5PSjD7J0gfvkFPz5xMAuviMHeZF8ZxaV2yC4GtqHs9dEpe
beax/eUEeXHXVVJAKkLVL2KXgAx9WZ2s8NBSiLWY04inDfbuMubVJ6bL+YZOprouzECPxILe9Asz
9QJ2/7aHxChWqqbTsOiwmcytLyDDM5hPgI00o/Imfs7n7RowvhoPSw3MCglmaeFgWEsFb3cuQR/1
EhofMRG/aEGRAmiRKCsMQ6ziRAR6GQwck5+2bOSyjqEoMdnRO0yKf4rt6YZy9mGQLXKaUT53jsdn
9o3uNJJmvZ1KMuagMvV+yXHsdiY/5XNyZbPkVo53bzCNt5/RWDtel/lLgb5XmNxDLBLX/DjGvjlo
tG6RJHza+Va55ddN5B+os3N46Cr5fGjyBE53f04NSOmLet5mUENuwVVgIUIgqa0+JggS7Rp8t4Ud
lhWaH4QJUoGbHZk1PcjPVLwpKa0iLLOyDSAa+jiSkzRoszS8wJvh1OmybvELIEXv5yPA5Y/+hX0G
YSbLzdAYSfY1f8Vm02Dx0kLEVpkar3FdQ+4eGy4ZeypLcViUYUcHx4p6HUSeCiZC9f/+8VFE2c6b
XQgKc22pMC/8pqjLOL1P1jLJ6i9dP7HKncaeqmR8WOBGZZ10Q+pbrw3HR9Pxh5sVnQ3RFqraQbuZ
tQnIQMVbs5uBlNQFIfiiHBisH+8socH56jjS6s6IHayXx9Pny26Z8S6dmuuC76IcBBZiaSfS7i//
uqGSX+0VoLuL29N1/t6hAxlolzS+DUwQfmULXfbb4h0ZjRfLEEZuf1pwwzuSrA+Ij8hRxLmJgjOo
EyCWRWj+Bfeod7r1UJb6jAv8/HwaZmFhPU80oncAr43+X/aud24+GiyiI0SzjZTvJDq0vQxifkin
OtSCcNRqSiJl8FYx7gg4h30CCc2c0V9PMycs2JBzFmrS1QL9P17Ps08Kzy8tdvcajHXh9xAjioYe
TnzOTFMCF19/k5xaUCyISeLhckMWN9yIE/bB8vNifk0SnhjiQCUGLokkNGy6WARfniAjGTgkUMsa
/SYDpmXWiRyhnXXzgC958gX/q6nRVrI0VrSdNABVUKDyuCHb067AfJIp6/5ahciB5BapttfSPxN8
2qPjgfqSJymE1zlc4GpJ1t51IQr499wXb6xTvSRRscKe/2jE698LU+uLu+sR4mliJ3B1VkUoxrbw
WnNzEit5z6gO1gGISF4GCrMURUBWRn7GGihI5MXOpswkXWmysd0wx9lvS0PDH1E9wF/S5D/xWo/e
C5kXgku83VoJZusYHJAcBbqU1/sqBQUX7aaTQPdCsRiU6S8Hg78sZAeStP2r3KiDPtDjLs0Yy88P
KS0bA6f9v7ywAoP0cr9FhunAH4dMjZgJyva/Xg7o93Flpl+qslyHr9YiF1KKvetLcgOY8VaL4ncy
ahyPqHeuhk3PupvrOq9ToJJeyybbuLy1HUrLNyCfvSejNlQRyQqh4YprJNPUjREfTeJDRKQz4oiB
azg+uZIYTq1iOB5vtGbXV2gz6r6WzLCze9Xp7JuaKvgttyKFqUYQNfoyKNBAXgUMyXFBqdsKPM2m
v993uBjyhMH5HaLmYQbyKHfzjOLjrY1m90apYk/v6Sq0Po59wiUvE+r4pi0DsMdCHZJGKvlB/Ev5
4dWQFUcYfa5VUAKtKm/Ms5Nj22rv3spUlSEhCTHOawE0RyhlVa1M5qD2MWmURwxb4G2uIvQ0pj7y
r/rBruF1B2JkpOw7vjZ9lkL4xQfUZ3EJpgLazTJ7uVFOzgsUSRREZn8wcg3yiCVr1dKUaS+fjwDX
8Ba5hjoO8ahURuoWiYwWtMLPR4w1zIb2IJmjKngayZc7dC/S0dViv9e0rp7q/RN3FHhTznlUcGBJ
hnfXI8SaFO3KF8HkexsQg96UgmsUabveJbNC4vCogl45Pj0jZTnUSMrvFNZ/PYa+CA83fVpFoich
3SO68xThfGxgeQ1hmo+H0ME47LDYTPjQDYMSpEMMO4qQda2VTG9ysdnmmqZqaNL/P1f2IehJ14/W
90ePWu9LoqyrcYdebEqOLD+UklrbadlZBqRvnKRKnTvR+WcmHk2dQbvPYZdRDf/5KIY6ns3y2lHb
XvauNI6+YaMxJrWweuUEyGWClqQWZsDQSWXgR9IMFXPQgaOaZe7pOn6pywK4Jbwye2Is9WvQ4wkP
krrNKH5a5cuVhtK3TkqPyn44OJkzUCbMT9RBklD/MOpHTBxUDns8MMrRqlupe2cJDvyUCsyvNHEn
Lhntr0cRPILy2KhnW0n7jbNeruNxRHov6VzUP+Z09qw5SubFeSexc5BE7w8XtYues2sSwu1IJfk7
OEqCQA/RMi70Wd9/mV8JopmkP9Ufl89VfEVdfDmoLNu00+FM1eOKKUVzOs4UJE6wDR8ABbSkgP93
5AyAytQULfusSIrrvlFeE7an27tKf7U3ImM+mn2o9MjdODRr11prw6c3zXpn9+6aroMRu2KySrmj
q0G80m710XvxCauEfCZq8mdu3rAoGC7bbtHilcU3UM9mh1nG3a4v6n2csq8TkWin2Diw58HW10Ka
NPA3YC440X90hqqlbVuediJg9ZdI6Eal6SkzmmxqMzqVbADMKh1og2ZZHDqSA7SXHg7eqV4CJi5B
0b5tG6V27QY+4isLOYyEw+Mii8KPb6HECls7KZfES0rQly7JUG/JECKd2A5E5YDHpOgvP+wrtAYN
ewJtRGv/tKnWtz+HPxIUJrwuFPf9WPMEnYw0xgASpKe5M6VYcx1HcxE9mh3TRXNyQR4m9lZ+YRWj
FwVe5aW1mj/+uvmXAazlNvbW9tWBOpMC3bj9kaHP47ZcO4qcMQG2dwo1gyax9ruTp5QbAtWmsZQw
gArtzhUdeMcVga9lRFFwM12tE9Vz9I3hqWZgprhhLQsXV9SIlt1D8Pzegee6Sdqd50jFznb2ytHY
vRvCtT+kdJJWVSFX+oFdZt/WCW262CRSl4amTlH/wpNZrZ0/41TFpjKpI9k4T3vn5/zNd4XKuF7N
WG5UXUdWSTfyhdXxfoPMQUkSrNm6AazCHAMVc8Q/U/b9cO97kukNmPDhSdqjpPz3TiiE9Ttwgv4+
Q8ZB9PVrr9YOpP+ftjEs0GFzJDGgIFdc649OUw8mbLvVlzJu55ea+7hBQC1hpyI1OHYNHK0G29Tp
vdhHtzGZr7R5sBRpdVPdfZHEvQGECGZPHnOnAgJwKFtx27923SVnCtSmhC3lESuJyaU0W/ixmzpp
bE2EDozsy6ixbhTfBIQmZw71BVuqlA7j9Om6yqQ+oP5jT9YmC1oqvOfnEUck6cPse3im/h6V/uth
mXVHwWlg8yHpD191THkVCPiJXu0CySQXQtn0G2cieFy38oESepygnq3ZEBPLAjQdO7HTUjgUbHR6
G7khyBxbIhilFpvOPwNUqKWtCKHPeZZqBO6vUJxl/Wk7G1BolzrIRtecDrtl0QP8O6l+W0/QO3E/
6XmwpJYpvuALwxd5oDEWyhTsHZPQSJyORai+2nuXLr1qPNamvaDFgDpPdUmGsXc0srk7tERwmAmP
xsoK/yo6dynq+4NY20Q3aKQ66LCQB6u9rspkTH1RtvGldMjdJ6iFoWOr5vMDAK7RrgaCrn8/q+mf
UXL/3llnyd5/2a30ip11LSV9pQEAWR854Jcz0zTGgVvizv+dqE4Wfkt6+m12BbnTLYavgKBgSSlB
eT1kmZLCR5vn26ynMDglDdQ6PLlwUQV01Zqv0ofhelnJILzoZAQiZqhQaKS4rSft/OjD/G/8RKr8
O0eBnYKt4+nKAtzVikeZlch8SzTgA1v+I52XgsvDnNIsfdqwNVXPnjP9x/3+BFdzCXcbrYwdIrIL
G/VZErkG2PS4HKlwcefyUcEFiQo5gnBfYdBmedJ9FwN3cXMDKE5E9S0Oq2+ROiWx7QKrXfgwQpZg
ijmfzMokDthKH8CoLucmvvG+CXeHlv1UX+pkW6NGfjpKpHNAy6FMK1bFPeWNyQGYCVxiLVO+mu4g
IOJT3f1wdk9XJGU6fgcb1T8z3DdygqixjGJJn2NBj42HVAFw8JnZkkm6sunwo9Vp1UPMAG1pHiMA
KBxSssMJxZ20VKYg3BKRmOH8rlTDxDboQxrz4sNA9sWzYK1UrqP8otK0m4e0+T8o98EmrBKOp4gS
XbS+esN5lj12sMbFb5KUlnYWvA1PLrG4g3hxGwyvlVdRIBXD97PBfM0GP48zq9XZx8ImYOTnK8ih
aLbrCcS0lt0ZTAX01wVdxMuw0HccDyOB5q978AYPZBCaJJ04VH/H5rWJxoHmNe7JwJU910IaexwV
YsgMk58S/6hubRmeyBlpXHuOzjkY9Agf+AXqNEmh7ktSxaP9n/aa29ntC66fD5z1T9F2lDqfteNw
OBTaLzhQntg2bYDIuyKs3rynZZjvOSBVoBOL3VUAbDwfinPxZpCQW+xowOrkEIahHBJGP19UitXb
auE3YwC6LphE2oEULbZOE1r1GArP/tcsZLkbpLo28CodX1YZNLEs2q0N1k5DgX2awzNw+wq5U3DT
RLsOkNrzo63RJcuWLaG6MtEuKQrJhlSogcymKqRrV82Sm+jCucP93o1iW5HzBIPliRw1vsMnkAqK
IY/oLnvJbBzoXSIRLxLLCYrvxiMOAIy/Ydq5/o19Kbqi0xn81yGsRnA6AC5/RO2NIat/W+qRxTGu
YUR5Y6djo9Dqc8RTHrJdxt+/7glh3DEmMg4dfBx872uvtYK+hkkaLNT5SWXlskzmDK5qH3QJMLZo
sltGspkwvXfAouD7bdfRYf7xQfuUY+sSeLhaoiEdlSVzrq7pl2lndRxc8+BlF0/Xyg0Ox0161OCn
Z37hCVaoLNINj3ZvhxM2n20EfwNIufx6FIAG/Ld1/jr9q1Kj8HSxKzxaO95ylD11OKSxsh1XSOkH
jLSvDAJoxyeSzM5Dj7yXiPYSpRxojh5xOISKHK/y6ljgcHFBeDcpk7hw+wgI2sXoSIxjE6EzFxye
XPH1gj7L4mdjHE84/G62lQrrVLqwG+055fl47ZRuY6t0AUT8NHVqKV8EdxSqcmhvOXWV0JY4x0P9
HkZAUu3vdzBJGJziBMIspmHyEdEilazE7kUAAjgWa6t14KHdOP/woC8CBldIhgf1sY1vojEFKVM8
A4ZyrolBYPXiemAYdGrTV4Iy6SUsD4lboZyqRf8MO2sd7BzUUnkNjNTdgtugn/WLvz7P+XXrbkzt
4vENkZekkaIZUTwiPxZ7n3q718+n6Cz8lXN3jlwPTFiBKIFH0t9ZG12BbvwPY/FLuKPrERJpdy//
L3IhwB7nqFwlhNzwDoFixwG08qAgTPtud526A9vnUc6pPZNOOsAyrTMF8j5gijEiGbrtJ28xXf4w
NUytx/HKtAQ02BBgI0cYgNAXKZ7OsWxvuyUfTj9Rcf2J+BAV9zkAL3n+H9M9NtCpu/bhl/epOL61
/L0/pSTmpfr9K60s8KPIOBLwguBrQZrI8BnetbNOV8dIckQ+rz+sXh90UUpoIJUHFEOHpmLhVR5c
kyK4JcpEDCW2SZuf1U/wczrMLOdkFqZz/NPI9+Cvf6ePtRMaEmo8nai4DX62dBJ608C0V5sW2ANl
0hD1vMskxu4vWRHOK/bf5fJPFHAp4vVeQe7sobCd78wnf7p8smWuAVBNTcosiy5k9a5EiL7u4LhB
GdPoDZ5mww7P8tKw3oFyCQ92BVyofFOS8hJ1ZbUKUtLFvQs+DWr40uiijaXjCbG6SwBQKAzXnjpe
Jd9jYFGp5D8OGlPSKN3gYacyFZsxGI//DZBVpGJ6ua4atonbLPUOLMOy3Modaj69JYOZzCfn2r93
cDTZ3XLGz1egeQWtrvTk3bnYTSc2rb5qHSOHSVxE8AzJEODDhP1zQymab/bD0/dS3qjosMBQ9jTt
6KxL9BnwqJt+LDsZkdMl8/WR1TsiUeoZk9Xq8jAPSJWvCpgz4lKrl0AMlNfvSWAOzOZr0D9KkFq/
vKd+S+cp+YFtvtScUiz9HvcYPs9KWPhlJSLHUw31CJNba73xdLybog+ymJF2lcnLOVPqD872fWFy
Du+q/GOFIU7XyZRFC43/nifxc0xtWdCb5l/s5z5oAsyIr09FOmWGst4kDuYLO9VHngtm8K8PpjoB
RftmEifzv8yp+xQho3zf0KHNZXP3DMe19g+YVfunnb4iij8GmTo89zFLV1fG/P4Iw7MXqP5NcHl2
buzfAu0JOjGQm8bVLjEb/KxiGUL4LoRrYwjBjFyHSQupz/pxamncqDDQoV4ioEWKvVPCfr039Vu/
PavbzoBs18FvSzRCki5BXVXtVwMFjD+nJHSavp4BlhFnUtzivX75UIKMpBZptxOyE4GQKAGm+6id
gpsu9B5TDSqhFIK/3sAvvlpKu6U5PYVDWMrImURnpTLCC+EtZwo/CUGwLLsqnASVABFRxoHLt/j+
pPTYXpvBSxCzyQBrKXa/SIwDy8mPKhOOeYYAh7ukKd71FpAmTjAA8wWXyMtBBnOIbjfo+6dGgRzD
6/MZUebGF/KBXEsqtJlh73jIdlc7pGiKnCdOziOQD9WmE2GisW/7Uba3FDeY3Gke07a51MAus0nn
g/NaMbs+jgowzwK41xTi9T8T7WVOeeXU9tsr82Eda2s68qRSZ6SvLn8mUnKyhzhnMWfrlJqslcHn
uxAOqNchnMMoEcjrmrGojb7RGTbuKlEf1B+Rt/KZ/K40f6yZW6AZW7QkkQpsyj/Ox78Ta+30RxwQ
VB2z5ZZm7Jkh1Z0Q//Iyd+VrhV2lV1HCJ1z1xGBSiv7tEjLo6GYmSiVkjURrWGGbAD+Ivz5I7mFK
c8z5CSnd1dsQCWQcK8ZNlVFt7ocuLJO+ZsiTEsyh3bO19hjtngyhG+N2fL8r1zkOon5tHiUQVJqa
TTGiSkblesj9tMYfGbu3BAP3em2jjMsRzNbtnzmtUJHN/IRO813/86QzWhgUixrRThUvu6ishi04
fpjzGfeKbl7VA6vGOcLgFF9MspsG6u4tAznUbmIUInugFjZt+b2Hf4jU+L8nvscf0bwlCt6EvlJl
rrAEw3PTrQRANd1IzzHQY8LjdMx7zsRiObO2IkG59SrSRbtLdeR2S+1nTAKjkMD+jNGjdLefkdKR
M2eijqjD2nBmG6nS4XdjPouOC2Vza3lM9oJ57t5LzvtT8aKsRXnIX7maP9G/5g+hcwi5ycOUfT9B
X4TJDoS2E522Bdi17m+LPNL9aBVFB+Js9htwyoJjFUSDUr4lyGDGtp2ayaQ2i/SdZZAqD8OqeR1x
Svmyk2ZhJMKSqbpc2DDXYYsHEVqrFGT3Z9b84CkDoMgJPPfSAaa0oIlnlHSi5UV7PJFXaAe1uFf0
26Deba6v9mRqfZkHRCV3Zo4E7CWx9BtPH92t/rezTRi60zwQKfhCgTF5MVM62XVIvNMQXqYIhs31
jij6UrHTClXwx4+pJR3NvID3ncPIcLPpSlCzxGT4i2LT5K5cHYYiDS/EpKLFEsKF+tCrrxaUrp1S
F8ufuYSmx3pmfAYhFNIsIVkrSFpZhKGsP5hyk7hnM+9I8tzgLIVb9bE0r92n69PWkkXQo7A7NOm+
/pbc70fMsLhdIBPzsohaARGjwkJOFpL9IIfPaZqUwuMZ1jdnn7L6vIWFRIKqdNVIM4QdApzCZv0T
nbOPPqcsCfcnR88W+BVA5en2V7bxourC887QhQ4PS/h2eHdtWTCNh7H52PMQciAAU6r/uMbqQPIz
4LeDCAFRg1fSCjv1nJun4tR+HgD54tQmVZLBPnHi2HcqQVesPFzxbTT3Sa6b/eWh9DzZS7LFP2tS
aIQUxZzgLMyvBBpFOByR5TzKKmwrSDTHpUrXZHXz3OajSZaAUlVIWiOinfy/7HKjIEyfp1WwbwsC
GEN/bk8zp0uVk9zN9j9biVEWE6joz9ByMfqT5smX+QrIqXoxhLpSdGWgcGhUx38YsIaxnOgbe9yP
WK55L2j92nDiVNzE8SUm4GLboNEXWVQXmkb9MS4tNHcwbQVK+GkMIRY3ejgcFXylzSyavZJDs9lY
qRB6sqmBzWK75dkWSQXhTPnFY1SL6hdvodnv6MJ8XF/Wauvt+ILNmLZ98/tQSChbKXJCeXSe4ijV
fcdqPhU5HMveVrvpbS95HUrtUcMBfT56gZClkwZ6TI6N6GYn6Gg3zu3cYl5rzVSEXNWppScXay4x
xo0smF9JoVO+YE2bralOw5KI0HOVjLh8ql9fISF0+ln09lbhzzMoA6exl0kWIAOyl95qDoo1K774
zqbXoP/9zMrPOa1DDMzXXR4KjYjOx66c+it/tHBLt0o9H580cMa+qia04b1nnMuKZ2umUj/31AtP
IbowV3Kkg4tpGbIkv8McAKA8pn5LdoOu/WobixZRamJ+fedRyOSfv551E+HiQsxN+rztaD8qPPaV
5TU5tH1+ofvGDyfahWP2BW9b7+7DVh7mKyLVM17nHsHAJbI+JOaoHjPYoHFCZW8DRC8KTio8eH4p
WVEYOsva+EybT2V2iyEzH8yguBbLsE0QNQcmKEHOH7lDFK4bLBxX7feO0TEAFvCucxsksIndnrgJ
a1/FksaZWZnTBMZ0bI5lYXSARZbHbmLKeHmM4ZDEJOZWQTJWXyvcGWAtn6cWvR6rMEB6oyaAmL/A
r+RLOV6TLMo6jY3gLGlos4xdq5Xo8BN26m734AorxCgO1tygf5KlWjtRo1p+z+209riT5v0FnU5l
AqXHkAvn6ysB7nrELP2/QKXUfJD1g+9F63EGg7rHkF1f0gqEanHI+FbY1EqWM0JHv4CfTKvtNkIo
kAh1/tu/Sl1iNNsUki0Law2TnntJ2mGLyvn0tTDiLzZ4+EIpoBbYBNXZIPnvomIs2tFeWCd89bTf
UPm8yOq1b6JTdyPeoQpSOmcCCBoaedET2kVcsMVjwwn0VCmhTwcpEQFAPh00o4xxyOy5MBcFFNMU
3D713LSBdoXJjoqwV88u1C+pX/DJ+j2AzgLwPHPGLZDQY5HuDw+/hKLPatirBemtZWJ+KZlH4NPL
fT698RGY4uTQnnbRslS9CdOeYWOsPqxLzbNq3pP6p3sPsICit6JHcFSHHkh97NeT+ZPxsY4uS5Il
n6cHqEOXa/S3PWYh+ZR7i/gAnCQ8dpQ/Qjv0Z4V+MEq6BDt+cVTpi1BUqSxGGc8bfZqGfZvGL554
i18i43Ebv+q7frXxvtUq8Sw7dC+kBKwfHbqEq0gDm8/EncorwlipO2E07yYcmvbYeclWgHOl+fg1
S3J14Uyiyhm2pbIfQ2lv/40/ugW3Ge59UEsVAjM9ailIVSAAa8hXu3zQiw/hKuWkT4oyz5e4XtTI
HGR1fX4UqwwdVxSqXkyJ7oO5BWn84SjwVDyHL52DquMgmU+L1q5Sj+BHOHSYjmwfelb2FnBnmxrZ
1KirLjGQ9pgD2Cuv8l1g3gMhcgUD7ZZ0gV0TqLw0fv5TZwTys7yfuy5U93HrOMQF1kZVNvg3zvao
Pf3lFcS1JfKQIXjLTefG+v86NNjb/unyrZuydMzmN5kRU6kdBPSuGtoqSKDkf/pZtQQnOFI4aruu
rtVQlubyyBleoHerBmfdIduID7Y0sEsgYbFx2AOkEtIQqBnBnRmApOfhMe0+6qZhHDtcpCFtEdXK
PbrHtkQP35KGXJ2iyLi4ovfBYwGih3KxANPGrT3LJMli+UYuelF4505RzcsLDTuV/3OlYcsgGkX4
8BNzpwq98pCYarY16Zy8aPzicqa9phiwN2osAZYbDTBv1CIbxhaTGkyUTDnVbMi99tPa2FRT3kye
vrbOdBXfkdTOMNAKyqj8dBr6xQOTr8/2lLRi2PF8obn9ouv02BdcNO15kuez2p216ErZw2tugeq9
idzTrdWgLRHx3Kh+D2Eouh5Z0/jSXnS4Vv9LsoGxRb0DyEMafVFBVgDqt1Clll7hkxITOqw2qGMn
9IH1zlVZHES7zLgwvWNdubfjSYR+19IzHIXSP9LuzkprI6TFMjc+PPtO9HOHEB5Djcf6Xdf+YFh7
LOk0y5y51+UDw8CT5IfD5R1pGXzRt0z5DV12fW3O+x1DGiMpUg4phCuRDEkTlt2744h1Af17syYD
5v+lluNlwpfaGMz/3VArWLYSyixQipmRReUPnpErXGXoyNDwWLdkGy0/+u5nF4IRRlTkGVKt0IhL
LJ+26FQjH9O5qFH2pzov301+zIO3/RXAuPpaO8kTTyBgXockSefTTyi3e4xRRMKDHmpxAvLU3wLr
jUT7uPMAUOSKmf5vLF2gLh6Zs4m+LnzEntmfPGPH3CcHi776FwZgn9jBEGdOXkHbGRkmc6986Cty
RDWBY6jhbtKyM8sgBELMxPlT1V2zJqJd8PPFpuvBWi/8cr5Bx6uv3xdr/9vPUSOFGxUCBlzl7/Nq
GqCc2Mj0vqc/dU5MrfLYZ+LUmwk8zecw9nztkkJ+cjYb344etWhkCJBgM1gW525Hh8+Enyae3m5P
RQHqu92DODvMA+SfBF8CieXsrzZVio1Sli9KtPgVpDKpzzxwPFLH1dZxgIQZkH2gc8W4piHPGVct
UlOBM3eeBtAerwvlHh47+4ZG7J/sm2FZb1g3ET8mnsYkzYiSQYmBmccg0cpXTW8+UYd7udmolM/M
1ng/zkjZfKd8n9Ko7gc7iQvQZ59D/niusR7lDLz4Q3H06dRBhGlvbysYP22dzo6/Jv6uNLPgkS9S
5RgczeQpcsoFPZBMSWvtjipcWlQO/uNJACSiZ2stu0p5u3RyQ6cQVI3sY+7HbnK3D81HbkttVf7h
XsC5zyrV3Gkc/AhUczO7eujHPdA31tmHzBG2Az0EGZ0vFyKKtHNACqtiSLPnVft7bc9+jAwefnyq
F128c5Z6tdr/YEUbQX8gvI8+JiftGwAY9NWBw6TIxTzm04WSMNOqHmy4zVVyZtnYgwucL+4odDzW
8xCB8cGlznS4A+VWwZGYZAjwDwa+Uga4y44iFDCoWVD/4TudSRikNvecvlHcDn2fpxiQ0ClktCiS
TkTsZW6Yp3+CTU5HY1/W54W5xfh5eCqJOqNx7TjHRYKSple2r7uqtBw79ZxQGZkcd2XVR/2wnWY1
5/oxbAFknrqausPEK6vN/xJJujFnYrWF5shHwhe5C4OTm00ho0S11lF/qHTcMbuCRHsifG2PD1jZ
GU18+cX+mDU7jJ2Ur/XQ4RpceDTc3e4gFQq1vNofBmay3E2iTq91aErDHZgc34h9fAY/2B0HP9aa
4/hPWho4I9Xw4TkLH0vw1yxyG8cV/pmJXvcGvnqMxVwIiuQcYl+CjnXOKUtPDpgwHAmYZbUxuwSC
H/s+Xv88XSQ90pt2eR7N1UAGu4vdYJRHj3ZdErzoZWVqn6hT97Ee+i+MWwJL9ftHuRuGDBVdRsam
p2/8BetbrosXDz0bgdOQl0PRgwvH1Yiem+/LAhjbtNqjOrIS8VIITTRsF549TI6PcAxO/era6nS2
zwmowdvNDkc4s1hLgAAQ2yJdADvIDDoKXnCRaNhybPr4n9MsrRnRNwZBssHwWPTtYhESrwsC7bMv
h01uPxGq+vXLsh9DfP4jQDCKG+IB/oI+oaf+jsqcxKwTK7XoxvPWo91b+MGxbqTXf5vhRzTcnn0I
pJYbEQ6TiZUwrpIwgtNuaueGBdgEOKQAGbO7imUsVr0cDM0M65sZPe6lwrL8HmXhqIgAONeNsajK
hi4bchnhxibwJIr7X/mASaHvWw415J41F9Yg4IX6sv7GXHJ6IZkVngztImweer6+b/BnXnnWujZM
d3C0u3Ui3MJI7NdlruM+YJs1M9W9sooZfKWfvvMGP6cl7BHa9FJ5fN3caYJ4mfb1VJ0mYwm1fIT/
Dpt/5Yw7oz7XD+pJ4u/KEAD/c3FBkM9LRvuEryGtI2W0cuTy6Lk1z4QE3DkVGTo9PW6hhn8wOVlE
ClXCrZBWvrDrR7qkI97gmsp+R63StVASSrEzDYZVKdXrg4ye17aIEncLwh5fQMNaPrgpSLPQtKzN
KV+t+fqmbVqOzBanFOcdi5yULIiw+9E/4yioK0g04ZL8cktrf+WUFvJpqCBzkJ2eFtrXq1IQFsKk
zCjKmx9t2EqmuCCGE/+/LWCzKoG/yxGUK8/3xFfIZrROnfNko68HQ7Glg6/YLUgaheEq/Ik8Kwfw
L7lyxMFtjZtkG49zM235eZKxX9nkj7lKlsDEMHDUq5RQ3LScUOZRpW4iocH9OeUwvG3PGuIxnkNh
gr7V7T/RH7+wRd/80eQwnZaBW3eykqk0E298PA6zye4V3ljy+zG0/4Ia1fwvwYAJW3Lpewhf6fRC
hl6FhO8Vv5BK+fzDX7w7MvBuPuBChX2Yw7mSzx92sduF+fj4vH9XpPVEag+z7BWHdE4MVV7h7M1Z
zzLRwMo+m/FiS1j2T81Ddj7Sca+L/OkKYhdnerhhdmGNtZUld6aw3gnlmhsuRNwYUJ1ENJ+XgJTc
uBR+/NODDtdzQakrsxw3K64kjAvU7pMNYOpAt6jAOaAOSRyacQmj9TfyohcmccxBe/tufR9ZuB7a
Z4IR7/E19qlwgBCWUmp6T7zl1Y0uEhwO8VDL3vFcXKj2Lje9tgcdD5cq0lKBWVQHNxNGzcuITOrh
OpmV/XAd7bpXAOXXqEK2DV62pQj197GdNYL9pNBIDqonBgd9dQjcF6hjCllyZ2OtKZdLJMwUDBfE
M2+LNNWFeFbxwaw5pJShd2a+uOoNBbj4Vuvl4AzH7d8shNB7iD1qb1XGq9osQVVILONDpNKlJvli
nUAQjmRHA4feXd6mGGdum/ufOaxFEr8EJwwVYjE1Tm+CUL/B2PnWPgpEnNLomV/TgbmoMdUx+SKP
MV/MfgeBcEZmtNMZkSGUm7Fu8+Py0w9TZOPmj6car7FCS+qghwHEii13GFD2Kd9n8EAvX+FmgCwP
3BafKYLAKeklrCN7ImSh4d38K6cVXs9m1wRJau3lAV78B7NRRt8laN5V8F/nv3Fda0mXYQZNUUMT
nvJqUqj9ui+7s/WvjEIetln48GkR8jMWBLfotbpBoHnavCVd94l6aOnrk6l13SlTiIEMMrmsoMQI
V16rzmOiTHy7/JptZ8GzvcnXsSCezb+BwaLyr1wxmL9/o/XljAEVkw5bWKDJUZqy4BpU005bY5rM
7+Ssz3RnXSA++e4CjKEPuGQ/uH0+bSJDnRKEwG5VADIUi1q49w82ERwvLCX2b/JwCgIKDdvZo6S3
KGOXtHzIgKKEDtNRPgL/+FE0F6d1rPZutoAa5e/sdObi/bv08Mxug6X3bfv10kN56zTMusUXQA1H
i8/UKhW2USwbq6eBeJ04Q3b9LKdppUAEqhZ7eddjWzRjYxUWJMiF8GigtU94O+gqfz98yUp56go2
DKlzcyhl/SbQUg6sK10jL0RLAksSAfMLjmdk6WmE9XWlde72VlOhZ+Kc4OXai8SpyqRoMI6Pi94D
g7u1D88V2YzFZit+VftFgqc2k9mvG/coVmVHU79iyxhNlGMseinH/M9q+BzZzkUugd22xQkPZ27m
bs6le6lrIfzUVQq6k9Sisb9ZQV8mzCXVPmwevuOjLNlmoPsSFUqNdBxYBul1JiUDo86Va7LJ4DUR
mEYjmmSJDjteBCPobTps2PsHk0TCS7Pm0nO8ppxwYGDqZ6Xjs9TvE3EWYbnpaQjyebTvKnJ7c2HY
nxJ93ILmH3MkXXbDZHQsNC7IeTzpxGWO+uFJnIZoreOVSca+/6EPGg+Z/5uRhxQA9Jt7iJhKRVLv
XG9dxXtRz527A6oloXgxOFwZ03jgoIb3nuzUbgVf6kjUv8DdLxnSET8iq+mGIBK8waTrH/wqyF44
eyFkFwv6EwvTvayZjwO3wxIqmFPVkIeTkDMI3Z4Kj4bxMOvoLKYJK3B+v+EbpmCiEosVf4FgB7vh
TERCYgjMV6f0ijoYQO7d+pU7S/8/s3MergU3qR00PT2SJFP6x61aJJA4sveLXoJ5jn39gD/BdOzZ
M5A7TlbJns6F9usiozubRB9V4IaOS0EwToI9K4UuVzKxCUQNv0VurStptWNBUmcM38dT8WNsFNJJ
azev/hz13Bxf+QyWmm7rDcJHVt2TBQxSDzYqnNfkaQivNp5XbOqqsLv0YBwlX14uj/miKju67W17
8VRuUSDXvEJfvz/By7/RRiCvsnqUfiqJDgcnQXyn9802sLrFt2lXinyns5Bkij/g/Ib/3S6T7wbQ
hsKGV14cuHX9EI7XcbMcD+UtFm39SC8eYUwfktgW9zNX5Yo98uPiwI1WbiDdqC0uzhLHJOYZW524
Y6ROYIp0WBmRcXqr/M8a6JxHWJDJMMU6K1eoad3x4jPAU4CL6IL/BvjP4r8MT694IQbXcn09h+wS
C81p66c7/s9sm8kW7Q2YcB7DNlMDzjS+GovtdkB0ndyTFrujDXZs30ztfSg3V2PaKJMZDSwrKALT
BpJEfoZIarOYxhg+XFANBYaA0RxDrlDM0aiw8l1ZlOHygpElScMeci2GL6bmowWqMvwAZpg1+18p
9vAoqzYby92N+xy7//FWN0Qh41pUGDUK10sIaimB7omsFaY8DPIfW6aluuF4AXvTFgu+pTsBlD0+
5rzvMTpDxFjKPZFSRiBG9VZXQ75shiKDxkUpdEYUFTHLHCP2Krj7/ROEaRvgi6GHOL2ELnb0ZPVv
44i8wXMVMVbjFXbNHljIZEBeqybESFJwkPOlMrBF5wcpbTrruw5St4rmv6Ll2lpX02kjVkTWhB0g
WjE1XlxVopfrVidXRoN+PnQ+GZETDTS/wKYyj3ts6kOx6T+vRfK6j9Zt7EirStoVjidA6WD54ex/
HO4dzHgeJM0OChDyF99XvutfFx6umVO5upNVhStgjHqbNSNiBrmL8R2Q1R75PKIZanE7axWVpMfM
g8twUaqvPcwd0ehNSwkrigk4sdEt9heQHTObAWgUQix9l0h3ewUSV9hKfl/xA0kkrg7088BGz2tM
kZiYIiXBn0WfeyF5dgMprheBs7Bny28f4t44FY5wjTS4FPEQIYMv4opTKE8rkkOXgH7hWXEnnnl+
hL3bN7iSQTEHvoTK5aV1k3avH3PW3Qdl9EhaIOy20M1/4Ep5IfcAwakAhc8MfO+6G/j3nlBmcZ/2
5RllgwyA1cp79NrsiaprXARfU0vZqoDw8EGwy74S6YWFCbHa5+YmbZAnzAPMOxgD/i961mqx5pYP
Z7C6Nk9LLUnMR8fZbKZHUux+kHRcvxyQSIQfXYKVyLc2suKH8K7ix44DmeCvS+IADQL0owegPY2R
c+XUlNcbe5rsR0iQM3KJs09yVFsnyqwn0110Ck1i9tV+TnQZOR0/YeNM5zPUuMkKKVH1Yq8+/yIV
PZ34jCqCVi9RkSBYBLxROJpGSmBjFsdhwe0XTF+D379z5FMYyaegLvsJrFVksx6xtIrv63GooLWB
kABFVcihrVMHHKcXTCIq6z06HI559+XRPGsCRrAdubnHsTDcDc1r2qePycAnWqrGIzM/Udm2bG2A
b/1MbbnZafJEGBtepKE1yhuOL7/uLYxjvRghG51lrKZc7sAj7UCNLWzcaMI4du3Xyv16SCcLzMzR
w7GdIVrkLTTKJTl49nDewfl/mnv1NHUEn99KpiDf4c+kvzABNuE7BS9M/a3CJHuMQGAOIN5Q0FPZ
/SGY/hQsie3TlJG5KCURbLQhRsMhKE6xs6yZ5RLEUOHoRHq/TLrlbt1FFQvmUjXJhi53vPtPF6nh
76JYctR80RUlhVpxv2p+UjTiYKsUAapapnYvJgIGP30Da75VrHdntz311+dSXXb6mIEsHKqQLMW4
Dpt8sBEQUDD1jFetB29jUo8Rpkgg+zbWSlHNANjoavDkif2jzEKtzTO1hIgp2eR386s+EKpONZyq
GBMvEWcL46z/0tfj8+SXs6jH5lgQibojx7/aUWLkwr7edYOLRWeqsmM7ZFESbAiYoiyKZHEglikN
63piCeOjDw26szuj0oZOQtakNAy91J6yCNMkjBNtubYqqmkITlAFmyToBtv8Lt2JIwFuFly6A5Rg
4kiGYZszIK6CDXbsB2VSXYqt/bu4NuM4ut3ulz3ZViwF5kgb0bpT3dU/NTfODfEnylVhEjBtyRIU
7b86XGSeWzXI1RuwNbuBmqBq35XDVmjiHO1MGcv2LkpolpWN4TZq8l1/n+RpS868Lvpv61Atmf+9
psux0Xq5U0kquzTxitEt6FjbWVU+SHHOicNVhaJH0R5OEikv6vKCUc1KMQ+ZBhU0QZnVS+UiUKGY
CTS77OfJcvKQQsMepp/9LbXil3ZtoLvjE+F3WMPKAMeMoFleJ+BaSHDn1JPW2zdu20rX7Aw5qyxz
DeFU2l1j7r5VIC0Or5owIZXgqwt1Re1tzjES9OSSlHWzBnUC4HAf9II/YQwYsNlC4GmELTPc/OFe
jWqn/AQE+PeLC8sMKkNqXO4dIa0RhsCJGYP6JUnzDYkcPqaIlJbuhaejZCaMn4f78h3I/BmVAlbq
KU5DuORzX7jAGuN/FK9O4ybNxG0y4zkxKvbUN3Lly/kpgavUyvXMTL+WnyRYNeIqe9GztNbRrcjX
UaCwoWzq+LbuMaBDbOts/53hNyC0eNViqeVZdEpNMKAqa3Mi6LghPdOOS4i0Fw5AS3B0Rmv8394f
WdC1DMOLSF6zBb3fBwE9Vvtwp6j05AiL9430qg8VOY/SqJgNgRLW7uX+9vFfNYP9ZAMt1GprRtcr
RpGWpmLd8MiNvDxYR/rmtfK6Lt1s9KyyY8dQAOSeTiUFn72UW/QCI2PDuF4p/M9zb47qQkOCbXcf
CCnxcu3kvDByYTeydipwLoJuRJZhmKJq4kiWxIxHDQDg9fMhDiIoHpE7dpDPUXfHXDRwjP73B5Tb
XvQ0i6adff2xiGpOG59e/0TCiXeNO71n3gVz9kPbiFG0iTam1WQlYEHOxWvtL3v4v6oZO9aCr7nO
U5mAQauo5FnaL3dkFWIJALweIF/y1wlrBq2MwuSYrH9nfnUycm8HS9o7YEQAHocTN8oe94QhVEtF
BPPh7lX8GSk1j0ITZpQdWrPGb+dPgNWH9SRcDASS3s3Kz84o/U/sLI2imiMfq4TUqCrF3aMVW7fO
iWeq5EYZBehoyX6DyHdbARb3VWippcs6EpegXvMir5gbtlQoEtUr0HZc8q06kHYUqYTUrzY80AGN
G0piAQch9zRDyBX+mInzBW3dAw/XPGiQRSyAVM1MvDE3v+vHmkhk+2gkV7wozsrFhSqh6B0lV6Ap
hG5nUFCOA+z2fuIaehYnlWBjXeOyDeeyxaWQaW6bK4Ajj1oofIHTHcltdXDfso+tolh5J1/89TeV
gYWpVfJz08sPxzN8msAEqZ5E4fPxOWo6GQInVYkeCodwChk/pujFzd+nhLtN7vqwWz3t2R8kbPCu
ufHctpIU66NlDkV1JSd9AoT/Bf4LQZ3O85Pq0NqKIV7ycnktwhInwrxO8v04B3cOzGGPie1pO4zB
BZf0o+1ZfWFD02TE2oS02sCFMQL4lMQXfngMNNPtS7cGWExRNrvUvvWMTyswt3kehfJZx/qYtapD
5YH/G0tWwWhaMYB+3s/Cw+8z3SF/efjItsWqxJXT7e2Lpxe9GcFtxxA74bJaFuUkMukCH6QeeHCM
Q3/bhdtviF9A0NZ8wdxOGPvA3MsQN9c+9WVbjdXuGk/zJ0jAzCA+JrpbdDRIXinNkd26HPeur1Gv
4ki9EtkyeiVZc5Nf79hDTtLj3U/uzALHL+fWPCcJ8s7s1SUxhf/k+b/t7GAxolaq31Uhz18ET+oy
cL9feEBuDiRRH24NShnqtlVI8D7IWe7YNmreilHvpg7ILAhLIdGE+YvvrMlCvlZbV6ln7kG2lyGF
eTQ/LqY2GL8gNb/K2zswk4cpaWnFwG0RsTDm7DEVWieWR6ymys1uc16F1MHEsIdNRJjZHh/XsIWq
ymr/NyhBk7jEfEqWkO92CBolL7jeT9e9pO15FapOXviT9bNVvGOMUQpYm0Sul/C7G5O35YKyBJnC
BAWUkxhVQGjw/pCDBZug1kc7iyhQNUq7kGW9nD3r8QBP+j6L3ZgjkOeEZqMCo/pqfHSFBcceV1AE
+VqxUowq07OzdYfRohNqgKNVOdrj2L2iwW5IktUOpUe/sBB0hQsEQqGo3GibDDQ/w51W110bTXow
ZbLHHSPtCR7Ac55sGrrzIfwuvLa1LJHLqMY+gdoKhgxnA7uI+xqWntWca77W/kdTyca/nm5DWEOH
ofJ1TbGnXRMg7mqA5c4rgLAOVf2tdA7bsyr3nojA6Llkg382M8Jjtx1qWQ6xIeAIB6aLIAphRrHJ
D2xWGdaEeKg1mdzF0IVw5T0Ayb0NICxDNrnP3HC28yySsY9qNPUt0GEKB/8cWvyE26BCGfpH53U6
78ss1e5nerBgrIXRxKIenlUoZHha/IJmepnHjD3JtHvywnLVD6QjNwKjs5AIG1Bl6TLw1lNibma1
IHa5Fk6H3kepuJ2UZdAUkeuAbjlMV0tlbtzkqqY3ZmoxNjj31FvAQ9gvUBCXvaanNAVsEN3FpnfU
UWOvnYQIW9ydfvsVYN8PkXVxQCgbCVvab9CcNxzmbK2duPd/BOpoFglHibeQLXJK0Y0Kj58Haptz
kan1njHZcgj+yuDzUc8Z4L4O7gG9+78KzoKuvWvNQh59CqWzdVbei8xtmHApWYLuTxyLyT8mZOM+
ALftN7yJzNMhx9NNCmEIxGc1ibWeH8g4PCw0a2ywCOyCeKH4KTwwKDObe/8u5eGl5tTQVoWVGXdr
+h4edOcqCHO0hJ3pi66I57wHf0A+5teyZXS7qATYwoHJriFDipX+0f+p452RF4sM3sE1RNMtM/D4
b/R3GKskYJVIzSmnnIXYfAr18fiexFt4mfqAJj8KXcowWoGcNj7eBJnzHnbELzzGHhVZtbTQ4auM
S8zN9d0DOkm7pyk09r2VIsHAMb7YIpX6P4NYeyZzexaT8ZSnk0UJfAOaubcej6LIkC+NuRM0nAhY
JwM82h1IfITawO1r9F/SlL52HQlRiIfos9SRwzyP4aCZr5GXbJNqkQN0FZtuprKManfZ518Ge8E3
QM4wMX+C6vBtqVfMHtsQj157wWyimJsQj/sAhNLVIVXz3i9mdMXwTro2m3a2Rx1YapxbiRrixZWb
DK1K0ikaVds0Wx2mp7rWd7u75B0LJonc4rLev/KsOA9Iqq6F4AZlqoj8PgLWBzhv+AGMsC3SCNxb
chihuPTzBnIo2Hk/m/+h8BjqtclMUoW0uUajvn0dqjqH4Eo6LvLdmkpbE2zyoHQ9HOxYRRv1Ts0M
/Vpn7oxV38sNXEWSDZgfQS4FrsKncKyMSYwZ16BYfX8opKYn07ObhTiJ8IoU5xrmLuTbuXSRH5ZE
PdwU2dNBzNzlH9OyMGGJy4oos/siqP8D3Fdfx3qa+t1zeizIYIPjkcHT8yIiM0Zu7KukTI4aYIpU
Hj5S8M2wGxR3+hpUVmdNCwqcwporCWjC9JZglCggK1EtqWqocQhWlAJtbLLxWp/bW0DZTJhBDHUj
eTaqSMMJzqRAgWpEsQRUz/ulnZv/c67bnSh6LQb1Tl+o5PG6Cr+BYYf8rTZui6rUxdsdCwTaXU8u
2Koc7Q3d36GKoe6nFsd5VQXHKo3n9Nbh7OuUAdtTecPPAIHIbsUPbyMHWddkuKZNoozM6xDZRExk
FkZZKeH3vZi4cNc0pg/FfxZ4fpRy9HNguxdFQLhOxLtJxBBctahtfmuaKj2V4y295LvSTShP/0++
K4XE2OWyPDT6Jn/rEzskuqZfGKz8mjpXOi7qjvb1Wn0JMwlRVzNWR9i4bYW1bb3X9jibcJYCVVOI
zub9FRy1PaM9/0nCa2r93yEP4bwjN0VmF+pjBCpD/hLB+TWnRx9eT/7i7eCzM4usR8aop9fPgyUl
IRcqCLEUpZD8Qj84q+MPDEM607TKPK0j2O8nn6E+3nQhw/KWYxs8pFAh46RXCWeU1Vq1h+pm9bLt
mKio0enAvboxIASkFOGBcLhESE5UVSnSEFGRq8kZvIDiB/yQ7K7D3/oAuDkD+wb9FO5db7dG0F8u
6+K4nHFa8pY5QrpqJUfr1euZ9lRjUGxl2ZIK5A2UI59pJMAx6PwTW0UGi+1nxCeSr3GnChM+iOSL
sWz3lR4R3iNvfklDztP7HCAkpBrPyCHtE8YOts1FBt8TzaxSWX5eje17/qQgR4B34kXR1vjm1lXb
amlMRwN5SuGtVa1/Cv9+y4qTMAbKMNqxvmDaF/3gIyoTJFiF4PlzkcUNgFXl73rrrqXmapm+u5JU
0J8I7E7LsEzg/cfvBpUW+v1jj7r2FboZ0w5hcGROFJCdh5QjMKDwn1EGszz6TkHeigdzoiuxoo0E
pmda3YbsY6uYKtRz3+lYXgmlrNvV8IPQIad4+yxYqU1ecP/MJu+xrHe2ZlMtGA6CXtWwST4Zn6TN
otTa45HeBjXwEWhY6ip1cG9+lI6M+D9FC8dL4Yfg1eAwxJzJK+xHeJXx0E0IHjqib42FviNpmP/c
XKlCueIPchVyRFKFcbMJepR/kmb44hkvUly0vW2yNJ4iVYH3j/XqzJNHPJLPZipMJ2qui0g3tfNa
ypGjGL+gcNUyc6hBUIGd5CNM5VliAJBoMf0i2hjGbG07cD0kpMrUdPL4422czuOE3IjCNBm6Es3S
OoGywoUr/+z+pf6blL9xx4FBWlMStfemQt2IyIuJIITam1SwMvhv93Ik7fjzm6npao4YiAyqMs5K
CDT2lmwNUTPAx5SnesWvMqttv/qBOmlfUh9xHmkV5PUQizCkzcBTs+gD8kg1ReOxXdyIG5AoZYrc
cuTF6n7vFxIx7C3Cepkxxi8nQK4ar8OMfuXGkFB1/zM2KgEcebWbwVU9ZIIjEFi/YrkKwHbO7lMs
ahCEhXUa/s4IoPN/qTRe6p2If8j76E2C0q0qsjM3qvDTc46Kx+2aKruqqrZ+OcCSTB2cXIdlTpdZ
UfyvQFqMS/2eTOSc9nXV2PHjeQa6Keu6fMTz9D06GKoHf9AObzZ4JSxmGrwnXylL5EluWz/vxZ1I
7H4b9ae/jNeXWVbSoPd+saN2LoSiF5PuyRPE2PBsKRGCPHOS6A45v1DWyeIZOiF0+QJQSa+7PVw/
WtJIBb27GZ0ZsyapoOKJnIEtJfDUpxID1vDfwq24ESBcjZd8NkHfdTSLb8aB1qaoanu6GyCss7UD
7/EmmUqHBlKzrATHI+GmxYHzuhpIFGV25syaisEzPskH1AG99FL9gPeXtI7J193prZ4aJMQ5nnG0
vabl4QItyasmMWXXo4qlknZFqzQtuw98J4eWLn8gD2HgcOJty3eOmCio8sXkXfeyETobS0Kvtuhs
if/Avb2S0EZeKf9rt7eNBPyojD8NkYNCugAmQr4wy7d5andiOcGJTZZQwoE4QYVkbB/SUJKvsr9p
jLOWdB6/eMS+tEvhyfVa9vwwdyWU3GnjOi16b1RvWEgGZewljdtjFUkXGV6ok4VfKfGkN0jNtEQW
8du53qkQlbDWGSMBcoww7Qi3ppBYdlG62oOhoMQsAMS8ju+7FTp6hTGmiqL3g9R/2N7nEhA+9ekX
7tnyRdw+bI5IIiE0Yvg691bXxgnvZdTRbYoREx5C2TXHN/OQVwvTEt0ryK9l62v0mhY0Cr4mn94s
YErGxdnrHy+see2/hh14Xv/PNAlaHjkMdJHxCd2DulyquRIvf5J2ku5fj1eXjwy5bm6uQvCycv6e
3WHwonjmubHc4o3NiNfEYW9VcqIS2DJ9hAMUAa++KcJ9ZPu5SaFgsuhxtkxd9RRNNd/DduJQZa3G
7Jh1EKJo3VMxCAhMS0Tf492ij6fNlT9AHy5zjfSyH97tTKwjY6rxqjc2tfDS7q2aYPQug8bXhGSV
joGzJwJx2UewK43Tz2PP+fteGNqkwHNr0WQ331FGcyVskXXZntO6X6slwNTPaBdOrGRfQgLIbxTy
U2ePLhazGv91FuRXcV8TG/9ZdPYoLIi/pmcQW7zvIa+oMeVdotz6yh39X0spldajnSVMmY73V7Dw
Q3BDBBqMLgEcEuI3Ldzcm9NELIySz7CBA5qBv3tkMBfGJ5xJlNDHnbCk/E82/17NErhd5GinGvFg
MwEqO0fR2p7EcXeHBNhDa4hBz9UNNSJSbU3FEz/+J80MI9Ny1VWqorh0MqIGb2C1CgPHQtZjpY25
D3nLOzm2q68df45v8En7nD6LhhGVeL4jaQtl2w9taYnxaglvlNH0+PFgX7TSQhpVwI53Ajs3Apc1
ZZV6Cs24gHZUBk4ZIumqRazO76zCi5NI3DxMyufoHrSNTSpIJbDUXBujSDBXhZ334pfuluqu41VP
3TeLuz2cw4rDY6dggYoR/OTfdMtjkI7Uo2wN1SyQPkvX5ZDz7TflyqzMxabR7+BVmmIco09sTRUI
SywzJVSBF5Gv7CGxgW1TGPOhQ5/X9mhUNeagDNdIW4apdX+FnBxumyU9JkzoXeWCk3fiCerd7fmT
I+2apmUr8U3+ct32jn1ZhuZrrVpBEBGMfI5T1F6CgNvBN25Vh1VjRtiz51g/C8L50CIUih/7rDqk
zXnEXYPn9ghZNkSIu+Eqi6U6yrTKpJHPoMNkynSUjHF2aZ+37+JPkdEm3LbliAN1oTdX9raYaBIq
fJLVArpm3hh0Wrnj0QQhhCOskTOwY2qQmwEM0c/GD9hM/FUYOm9SP3l+5cSf6QRLyhXXthGtBwk7
ycUkcTzNhZl+mfivdpJuRHihfQllTLRuUM78VjL26kgsGDFz0V/pBiY7xpz0Zg4y1/z7zZPu+wls
ohh5Jkh6my6SA3w4wqVujw2ATXHcMnTqxoSX/zzanq/LdbnwNlYXDOA9zqP7PPHEJinMxTTlpnar
hWP9UGaaJrgqIKLwwIrCOvIQ81PdC0NxZIxztlRHnPjSmzhzEPxK20Nlle/e6Wv9G7wuDPfUSpPL
2VTjqTbujlThEkk9l/yJfdWChiW0FRuPPRyheFBr2oezvObI1+qcUucJ/vaKqKi5beQFCGSRQoc/
TukZJFE66F38oU3sTT4v7/uaJxpawWRarkFNNzkkfBkyzqaA9uLyP6g868LFumwhCkml1RI4tsUz
OpGGyRbUmGUBNL0TAl308krhFUnOBP9JHqSCTSsddfdczokIW4p+AtokvCiPDcdd0dyG1/brfa/0
fHCN/5quvAcv9A6U4LpeZHDSF9Ysbz0OgMjhfCH2o4rIKZCAIHcq8QVkGapqkP1Q9jwtgVjpWlAD
maAsHWh1LsemIG3ZNmCtLPlMSYH0zR/m9InBlLoSPsY77iZGMNrlahM5PV8Xmm1VBWFXuhc+JyeJ
R+Rwl4Rj544TUuoW8KyvCL7nVoXFTfhhhb35oRqTrZsUAmOgM46IR6+R+6PGwb8v+EUNWBLLRLQ+
FFJgSAHo3xGKvf0hs3PuNuWK3hommkjjyUV8okXkAmLDHcr5xibEXHityLkfOes2s6X6jqGmMA3h
LP2lAjt+SeBTIGYCymoNv+8fjHzDpfi667tj09UraoIrjIavCpkkjBVjm8JQ7jGKcgwcqTU/JjDJ
BYagVqYG7cnB16lrFzj02mhkyieX0O0XYjDfuxMypb2SmwtCPXb6qDOU+IlLnrGbZLbHPaM31Kam
bLZkwm0NuNGV2XNQZW79nxWbNTHaXLeKW1SCu7Z6Hnke/pjNW7EN0LJHMU6sCHtAz1WrAg2BWMMF
fGCzLXzfje+aIRtQxuyeDyqkAeLhJq9DKFwv3cJrm2hGbUiKJW79wRb0skyhvZU72SMP++pHJk0S
JVEsFp2xbrZFSEevQ/iagENXGUS0v/XFnJydKY802PoSwwqUMtSpcxUFaoYsfTMK3Jy3MXHNFyiT
6G6Px1iSKedXed1HDTc2d4b2BUrOzlw/lPt0tLE8DyLXR/rcLWQKg2dFrrr5pXYBU/KMOseCPmfX
lbrUVP1L5EsBF/UhBLOsS9bKxLUjkpjWIwA1jSTs1+Y3qARhx2a7QzAZewbSf1QFnr22EvmJd40Z
CQYQGj2mfBge5/1dY4G2BSpCqcNqjjXThVfNyshWcbJfuUBX2KS3nXz9vWikFrei07C5RBGL+vMz
d+1Mu01hKiFsJ9pplLRxJCr4l4mbPaCYGJgwe0juJvVPimEsEEUW5sTHFGg7l7qMGXYtg8ywFXw4
jOuXzRtc8z94z+DbMArthn4SpJfwksIVNsYMPUfD8ZoCUACqXBUulBDSo0/gPs/SW9dMi1KpfyT5
ByrM5pxlCCp4oAJfZP/Fe+iiW63uNf+oQ/5eChhbbY8Wrm33oRpdN5wzbtp6RnhSs0C/xJA1K9Pl
Vd1H+n1atLVOzLr5fqQuqAyvSo2wwale7Alduc+onkzAm9wYa6MeD9yHksIhLVqqOi6bEOqBt+kU
wC5Iz7W0kDoMyzUGZpzpe97KeinXKZwfQqIEHHMwsaY9cRhJlDVwis6/TRizuP9WhKeFcgiMHszy
ZRksLf8UvYClwEppeLG6nikmQxf9wNKkDg/9XUf+amPylXrvCDcLfg398lXVGE3L+5enHu9+wlk0
JkqDDnmPxmzj1zESgreeBw0t0zwEbRtvUXguYACS7GO68/Sim+S7pBG/SXH0/dGqBTaTFEEXXaGh
JdFf6xo0TI7LNs3ygWrbh7FSGnQe2kxP4/h0f7gJWlTs2Ctz/xaND8WIuA6MdH1AZWEQUEzfOllR
IhOpPaM/d3Vv52O7G1zmfMFUQtwhI+o7+dkBMJaAnFaRuLosVaW10kB+H8GTmZ3Y6hjm0qqtm9/b
QTGqdLHoVD5bJW7CjspqGL55xzE4BNPyC2TAqRwXOqR5pxbiTGW+PCy2ZfmjtswRq5g15BykjbGR
dlu4MisrWUyO8Qtm/RtwiJvbPRLKUB50M1Ymt2NwtJOZqzdU1vGyuo4P0iuE3l/UyivfGpAKN0Vo
2NHlthsNq+jTZpGhDrT5VmIdgRfI9RIjFbL0jEJWFErqCZd+a37EhopyBR2w6GRYX7OiMv2LVIeT
U1g5rQmReInB9PhulSVWbXzL3fyPQ1pJDw3vBdSKM+AgLyCNUhhSi/Mqr3VZGzEKYxlnJ3mUJm0n
tAe8g9KTERT07OBJQWxm0Lh0wISIGHjw8RCjmZz5quyT+qykQZRrOPjxCgduV9gysMGF5atpeR/H
+Ow1IsM89DqVUYV+yXGBpkoNHNmdcpJNXZ+MlMtEzCW3WOgPAQ4Jmz/gpRXXJnN4pZPuCUmtducU
cbwaKwUeimh6ueVPfzazmbsuF9cP3YyhJFf17a/dtCLIEvdWV69LfG8jweRGJDjkU1pZxVU7Rc0A
WQO00in/b/bDArFyXDNrLrdjcgtPARngwFlctFu8Prkn5qaXrqPzgq4ZnoaxsHTKtItBunBeioJz
b1P5h4ANP9z4lIEqo+ujCPQOxxPCCsH15CTPkR+NhHTMBOMHJCSTOP6VWBdIDAmCLpxhpu9s4MlJ
6I4NcCqJjbbYP1RDpXqcOFU+A5APTkNub6O9LVpj89gq1EdWI3JXyn16ePrOpVKbKioe4z1M1IlA
CYx7h1MeS2elR3ZE7wRnNYCJ+cMkH0YyK9AdQpmljoitmNlXlHr+M6+19W3pw8DZxLL5/cn36dLF
CF8HzAk1iwzhsU+0bYckXr+XETCUT9NCFglAu3URwZSenS5id0/A7zXaUYKntqbbax10GasERzPE
r6ljxuTO3/VgC/Fh8LNaWjAeF5zm48ZHthxC9yI4Zsh3nhf5CtXAKv6c3bD9k6XTxdEv6BwDv27c
wAUsc0kvX4yHoSYX+ewM6yOb/fVkRrfvrceNCu//3+OkI99Pq6bVjdnud9Lntw9aEKglnP16vBIB
Bz5bL5N1SB+Na8MPLjsm0Z0kCPT9VlypEW0V9MgXeox28p3aE/lZkdH/urVoZ29WlLLdkF5/A+8x
n3EB9YzP/5pLqFA6q6dIziXw62TaSTLCiTCZCR9eL3QPfK5Cw0vf4LmQnHv6qY8f6e/8zBv+snRq
LMYTiaXp9ZCl4m66cqU3KQGzTQA/IMqTnKBdG54k3RICIF8/0anvOPt0mbdLxsmZtcjh0Yysn+CZ
KQleYgdVuTSRoumPNQoUiH++Jn0JdJ5TRYqcaYqaXyitpxrhaQunHPMbMoY7AOGcmKb2OcS+9i2n
igL53S2qiyEQ3TcRuQ+YYq1q66zlPijZUzJ0YbGYhL4pljebLmUmo29xEXBefH8s8gngwM45pp0y
Cd62fzpOWfQH5WEc70eLTUOLbx4zJeF+1+ZHEqVL0+aALBrC6jg0s84rG5uyM2N14papi9GtnSsm
eCBWE8y03i+RnhAiGAzS/MJK4THx45Cky0/kX1eHJ1UpA2xKZNm1L7ijawdGn4jUcYaB6FUcE3un
KMtACakrAZUjBHOqMgai1720mjZVAbXkjjHGYX6dIty+PKKa927tgWfDGpML+OdZqMpPC7gr0q4X
9L9TOZnuTOgK3kJklZ8fRF/hsfn8Yh8cKoRh9yfkUB7MzfE+3DtJBzUGfSTqs3+yQCaqyq0eyqAb
LXrNKrAU8HkCmqvAqZ4L3eltbhy53Rczdfe4z7m61IUBUMzIL3OyU8pbXimTcEuUBIgKwuO8QqWP
pOGJSREZqyXurQd8OFDTU+PnEkYt0NPI0WrjFqVfwwBy+xNjMysngAawQFLjxdAwYO7qR8+pLD3y
iqHtDHWSZcDpNnKatqUFi46sBZi9wJwbJ9d3qzLgNn5jwQd+XtChL3rT8yDX2PwTOoy7io/1dGT9
F+2soLoTcWPeBoo9Y7FlN1MyVZHRfk1ECsf5+z3vyc6cBxrYYbedk1qaSErfKg4ZqR18AWxQqJ6u
SbdF9XkW1e2TkWfFkoWlxxS1pVfRwFiDjvxmwASAxDmYHXY2k1xy2s8dwwzvQHLFNpIP/MXNpT63
HvDVjgCnyV9mLeVlt+ahUNC5+w8bWL4h+Ue/aWr3EHlw2OdOTmGED+KN6Rjuy1URuDlQO3EQ4E17
t2JwxXD2wylFGFcU4lpyKfRL4F0PgnJlWMOkqxujiWJ1bRd27t798AeawTnOT/u2KuOeE25gmMem
6WkF1qnY5HpngCUZfQOJBuVq4W+2nNJ1DojCW36YdCMfpmWCx3TTqQNHk5K1aWbYWqkKQ6XZ5b78
CEZDgB3+/fqFmxkuL0E0OaGEE8XYBvfX67JYQQdQqLAy/+cI5JikYTR06m4bid1Osle69KrD82Ed
GRDU1TpDoP9wFiyVfkk9eql0sQVkmig8qx7ZJEe9C4V27Z36Kn8utz00/1Yxt6DCko8xb53n62h9
lzjMkrl0gDBctUF4F5PchwdS1vyDKp5nyOfslOWiZZxB63uJADWcTEjQ2pjNpmaNEcx1eMYc0mFe
wGxtw4T52dIOMp/9whvT/LfnHnRyBB+kppCbI8gryFsvE/v1St/+Xih3Pbn/tEb9YRC7Prf7hAxj
QEN4wfGAu5M/KpXiGIgznYvk9LvkVzy9YNhkeQwK+/1g2FQO4qqSAF7zSPpAzuF55xJiK4Z97RqK
d/n1pojGR8hqZ7B7lsjkf71s3yf3crhV0sWr4s0TsJg09Zuz92Dy49C0dwVhORM1IgprX7MTDnsk
f4qejbY3lDU01/2AJJVOgw/tBfraOq2kmTakD/WQIAPMSKNKvxCkJEtoV+DBOMEQPp1vFnyu2Di9
NKpSoSJlpGUQRIEefAiIny5+pYBk1y/lbtTrsijIa98vJOgVe8UAMq7iXJRC0OKlVVj862OAQfrq
g73O5cQ0c5ZPYlzU+HcRtXWlS0N8esl4dT0aUgt9+8WyMa0NJNlRoOnI4yGHE4RIgawrHZ957kc8
zSUfltW0Nvy5AxdsulIEGJf0BJsaCivBa/cw2JBmd5dDMCu+UwU5mPHZmW+9RYRz/wkpaN2xIVsn
6/Fn8jvv5Vc4IM03L1eVvJ1QX6/R/eyGDo1fnDBmDTx8FSMDJbgmMoOS4r6a8PgsbfrOpgQOd9HB
9kAIPKawK+HaqTh1rLRZz4/HHA1u9mTnf/xybwh1N1L+Zgo1IEglqS6wilT81dVFCxsQ6C2ZC/O4
Vrd1CyS/AGQ+4I7sLvu8NUaOwDiO7Vpi/sQAI1/arHnK33Sj7LDn3PBXO+1+gY63OqKM1aYrE/14
J75g6smL5JRJtsKEf6G9kQhYSJKooH+CXN4aTehTAm0PD/O+pU34EHHAObJc9qfRoPODPc2gUH5K
cncqG9lqi04kMhHxXNnFnu/azzIXafnOtOTdm6mwvx1AKPkXzpCeXv1eeUEvsMJP/63ljg1frQbu
31v/vvv6X4DcGnkmBvhl/KwG9jPQUz3tvfHhtIAQtvp5ykstIX0MHB97+1+XKPQEdCUJeiijyj9Q
kL71h8JVev9MIBe4knGB/3wYK6qa5ZiX5s0j8qgpBK/X2QsgxQNrYfk0LOcBOAX+QKBFF6M7skno
lB5vPHybBB9Ny0GDUXT+aNfDUZ0CNBBjs1hdxBTEf1ZjRhQZMjX74QgO3pz15Hi+4swxc8o5TTFh
jjh6NuKuYtCcK3N4VRGmLfTyvXNZwNXng+L/+4iuWsdtdznCI9iLF3CO0kGKg4EjwnfInpsfK9J1
MEW2bypvZOapDmVAMEG6JbhIzDq/ag18ahvSiAxH7hyO+BgDIF2rRNQvveqFh7UQmn5mxRggrmr+
XL4jDJoxBWL/wqBdHfnWod4CjkFBuJNpTOJtgcWRtzlCX5tMdXM6fvYIGi891a8NdJ6fXjDDaiW6
fyA44Nidjw1cZxATmQyRrTJPrUpkUVQ6CIT8XTmiUyJdIQBez4J8xddSXqo9YZbQcmFvnh18iQRq
hcJzng3i3KWs3PDUwkD4ruqNCxvtC5WmIi0RoxRh2NdZuRVOrg7Mi/ZPdEJcNe8m1E98Y4OmrCcP
qs5fyDXp3OB3EROEq75ew8FSK632wt/P66BibwOY5zKeJTFHMtXZ4XWo3LnNciyyrAu0iRga2EP4
mvfr4Bqg08MrkFCMzYQbcNUAfPUFMN1/GW+zq7MO35f6YSENrzUUtxZBi39CkkIVQIje0FSc8aLg
VLlza84kDkEcJJZ+o4T3uI//HTdRDEXRxkq8CAexv7DWWJkfViAUjCUgMvaoF/KJY6fBP2rR4JLh
t36tWl3K3b77d8a3yPDFdbffSNt67sctKpJ2rBYbJfsyrdT47bQm/TPbLK3Zmi+Eewn6XqYNs+yf
JtASTqf3UVm88AuNM0n2gLgkEaUH9DrXLKDAk5V+HHx1elTZOLHY/d1kYx6bxtEg3Z5pyfKObRzO
gxVituGkIGMmFlyzKlpxJ4VHoqkoIYcwfFhxQ5HnnF8k6v7uRG5eNzRc0eebMnfdb9+QFCA4VUBe
0h8h32QS3cM/folAd5urkg2FC8C3qcDsjf2gH3+I1bUESx5Y0cTsk0tc3YhIACSZaKPKuGWjZuuN
U594Aev1NjBR/w0Wcg2+R91BG6/j5KAJ4OVIz/VASigrrfk5BvkfDPGuIZY8eRkFKuka6EvlVae7
GTSSynyawlrdCfsA06ZSXPIfmFFbNlff8N/oJxa26Do2JwZTYqNMmuMqhveZ+ZWTeSLjJ+EEUW2k
gGHw/W3C08wW++oVGbeD5S3YV5xEzXtUsAOksZoSIWFO736zQOMqD9cH1PUEzCNkF4yiXzcKtxaG
I9tO0EjPVOmKEAYFiduQXeJJWY/Dnfj3010KorBOu5mg/ZIX9z0lJ/X+vvKpCKuXtwG8P+FU643p
7MQuXNe6rsEwIbsmLqkvEa5jgIav34C0DadfFJPXTDX+TdnDcypBFdqKzxeJ7mHjo4dyc1nkeju2
Nzp41XBPzvC+AqJNUe2uphhzFV0C9qAjTEFZG7K1cVatvtsrDxmjzOLQqWvH9uxediwz3wIDVkw9
htPvNtr9Tgm844GSuoRkXLxn+33yF0p4IkwEqBcsKMBzBHlQPgX3wPIADjUUOyVEmCxbGJa2piiw
hELPVFT3NON9WHcGACzBF6YjnSBY6jjn50KGy6WoAuKlTbjOK5n0ku6u7td9fL1MSR1lGa07wpZb
ijyTSIr/HGCE4Rcd08aDKJ++RqM3zQiDujHwWczZOuhX3IO0FoH/zopqxjHv8UgwP6hVgfChyGEM
dSLUJfJVGTti0gbyhVdmTvZM7vu/SRKRQbtaAKtCm7SwKo9xomEiKFCK9dBCFV7/A1CPpkK0xY+1
MvHoG7xoh5tbgbmIWIlek4sTpsWLIDZOv42QInSygOzVnPJvsAQDy6dsbYQCiBCIZmKAJKLd7sDR
JgoXP/Sbc1Scfl9eT2E+fPt1gATdNxqUiBGfN4u5JPHQV/iyNXtDAN9vTQKkalMI8jiJDxU+zdyz
FuJazwOV9IWo/EgcdIB79zk5vcKRU+lugdV5bmIe05xbdWg0OL4D/fjkIUC+fG+4Xb5NZCnXKqLr
hWuUYHrUojeSX2Lfk1llPHmYI4k9MYU8t/dEeaGbikX9ilh38mGaBK7OQXjV/m1PT9L442LL4xdV
0YSxQxnGXf9CVWnkZMmSjfI+AfaMKRS5ZQSLREM/bZu4YdNfc6dSnGSiUXXenuGhSS4U5BFve0TG
5cowdoRO8AprSYi/id8xEAJ8+5zSeXlDx8FW5wDsc3OA+wT+ZnRkj1w9LMEjveOfbBGhUHIZfAkg
O6qX7/cEEcJEcRFt91P7f8MpxrS5ABST9j8HHaE0Wiml8JOp27EpTYxdPtCLHtfY+Kbr4lUbIY4N
YsnId30nml4IQbZQqlNYkLI9woNGSYklgGwBqA0U4cmhbNaApoaXlUg3dcN4J1n63u3dgyXgP41h
AxK8mzhCMj5gusyPW3G8KxekLWyIziXQ/HE+HwF6QhJ58ZhEyezGC45kiDHNwpJNIXqdMw89+jA0
/jA1JLj8U6BR1HK35krLUMgb+fNmtSlLtPOVZUIBP9ihgNXN7/EsnUCNGx/PvbjAwmp+fZR2A4wG
nb6Lj1CAGxjBSDbTtlbHZjZ4LoLXpfTunlA64+YSiMVB4JV4JW9xqRFtyeGhN/4Q2wKZIqoY2Dz2
V/bWQu+5qZ/UU5YllqM8Or/YCiiIHG8Jn2VWifwAPiMOZXWa3yFohwFzkXuhAicATEOBCB2GD4cm
Ppi0U+XkBAFfpnqBl5SbOFdnF5C+8+pucyxjT10HeZKRxQZqkHlSPLIsFyQxFuq7JZp5bKwD/TxN
xr2lC2115NAR6XX2+KNY7ao7N4hHy8c9mEc/XJPb0uiUz9LdrRWyU+Yot8rE/Z1PdD2xfC/VyYxH
6kLiM1Aro27ojf+xpDK89edbUBnXNU6dFmld50j9mssvcgSADS0cQTmjwe9G/lfh6HaTdqOTONQY
h1x4oGUsPLPaN8tirfXUQYo1l3ypFxCWgluG0MOswqpa599LmLMKdq4IWIveOWJ+iDFYFD8mjQ1l
fphPJZ+hvOgdGiYHUaCBMrSZEm9dONxi1XiMEIQOjHVAAudHSPOIqCkewIJteWMwTRnvI7s2kQfn
zPDmu6ez9BSw7Pq6+NNbYNrSkn45Q1x3/9cTwsZBMxUUpl8BIxk4tKkOgO95Vn5ZSr+aXiRDFPwf
maOqzfhYB8irnV+cM3j+YqbrHPWdHM2T7lhRV5AIUDhzlqHRzMrpImKtt2Esv1Y9kirHXIHPjYWq
/cm99aVyALzGRndDerjspGNST4OCop9mDDXKFZJQNS1wSZyV0iegshXiuAnTj1Qg0b5BDi6679UM
N3x7bEMVI65bfFMpvrEZcE9kryogTiNu2SATIxDk1RpkX15pvvXmMRINkVqHc5zS12CJNwVfWwj9
0QGt384wYM25miiDmYzBQgR/Q+m1KHQ++Bn5/IuKbTfm2onf2JJ12kkO5ougL0oOH+VPGzl/r2P1
tp645f7BnnIubW4k0j95NERJ0wQxESF/WBt80invaso9gVbZGMUW1KV/OZAT98aX5JubtArhJcDL
ZLxsOiAK9w0StPLG/UhLw+AQloM0vEyaq6YM45gZLqWjxhfHixuVZwdTINnTPFScuu2XvY3gHNO/
hoaXZzhf0YkIcIKi+pYjFH/HewnnEND01zKC22+/ukVkb5XB/ymNXrU42LLgCQpyOty3aSIVjnVx
6pSQAe71NzyHu1tlhIE1/lISZHyYTwaXMHfKcbJo+iBaFe1sTkb+Jy5y76R3x5cWNMTRKLQ2XkuO
hrHBxkF++Z2E2Dp3m12zA2t++Y6QwLyRLXq76P+2AAtAm/0rJzYEpDm+nPdgSBFaKoWK+acHlQIA
tkO5l0vV0gJYejUzYea3+aAuMKrpyLQSCF250GVr+2KEfxgv2ikGE+wt9IxV7ygevoEUulsPJ4HU
4eHyNsBOc0GuEo3hH+TJXf7Tzdbv5wJjgHfqArlnu5Lu0RjnTdefmFMfQCVE4ZH6oKXb+ioTTJ6S
nLROhNUa8HB0MH5JWvG4I2Tog6fL8qyr5KyYXLt8plE599TwkN9nLROAGTL0ciyLCP3BLB6/naDh
YaVFCg/IVEGgTm2LXiVbHXMEqssHMhD2iZTSZcGcAy/5t8hQOj+eNJOrlvH5FTBTvgRueT0kapt9
YKufjttUcbs7ne9A7M6n8pG1K1t2fxmlfLGDpU9dMxtD/2nUiBKFxi4cuwkWgK3r0k/fnbVF4Bb1
CufPi++M9uKHcq7FpqHmewnpTvfLR0206X0IC0BA3QUnMYp/3Tu/smVvee6kQKXeo9uCUZ93bsCg
9Ae+irXUU15pnh5Lzs3eDApx0kCsNE3Q+L1vPd5Py4IAC45wQxei9NW0iYy7vq+Z1kY0SGQCqnDL
VNcOtnXQJ6M6M1oTLPPansDTK87oU/OVX1ttr/i6H1EYDaMrp30p2jsfgqjgJQKtkTCekf06xKC3
YfkhxN8zupcI1Io8P8uYMG02n95zSUR5EFMcPhsXlIpV7x81Yx18/OZLFd1DrWs1lH3g3XqeuQde
pg60CCvUi1DnF7FaFHTRATc2zcLfCEf33pMzp7vSZ6Z4BtwwYWiw7t7UQ4yoxFeT3qRrOg2cG2VJ
2J3Gp8WEmYlR1zX/JlAJKtCqlHuEpXSWsdZTFtqEznAAV9A8ZCF/vPJtJrCQaykoWmQF6EFkavSm
c71WtSr6S7mpvRgTQgvLFoBrMR7nfBjv2NCJdSfR/iSLhBplPuqzCUG2MDFbdX3ltiS1coN8fzCr
talGdQOMghMnwfch7cixE3JhtZiFTM1Fx06kpuEHfr9en1d7ao0inDMbk0XYp/2miATISWoct2F6
R+XZb/Y4AMXIuf+Xvp4NuxV6RmKX12MY8sif1O6cSmqjM/1reY37GV2awmpuor2bQ7EII2ec9sdE
BCM4Bk1JSD55cpMIUTCSUn5BULZNne4GvKMvaXNmRtJ8gMVqNb8qY2vDH02XJhjwL7pFS7ea16VR
o6l6ta5W3WCKySIFXoc8/vSZk+3j1k7BQTrW7Rsn6XgM1ZUILLWWvRuAQmAWSZXdLpM01Y7E8SAz
VV6vNF8uA0xxWEfeiuUswdUhFF5LW6CvQjPLJVzUJOZdKKHPA8saINbod6GDOTyVhO4xk58pLJ/+
ylMpHyLnwJJBu+Rb8kZfj5cIhy0HUveFJMyc1iYUZeHovyIB6etvIhhHYH0HGijrAkSw1/A8xOBh
493lEucWNLXA83RuDTyW4H6v/Bypx3QOSywqI5wydN/GJg/aOIzfaXmISCUqaWZ/mr2ckKi9ZLIx
IxMVPrL6baIznmFVEcQVXYwsS+vsPbkZoOQr0D/WX0Bp+WnAXcDfvvCUztRHhtrKzyUSjY4PZ3Rm
cRfr6D52HVbMxGshM4Th19Pci+lICVEPqf7l7ofa1JLULmJEGvGUIddz/AaX2qD4gcjRvuWPtZyM
grPYMxwYistmm1z6ZUBgqnD0FKbkFiCVqMVOvB2DCcfiMwjXYR6yN4kcqTvTSYclJanizXpRD7+B
4HsjqcSAS8X3G1o1L4AgNB/hM07kMYWhy7Y1lV7+zDvmB4JoziGg5Zkd92rj2gJbW8p53cwu86YR
lYSSyo1b5TIaM0mrRulkZVdr+FndiZbTXwjmvmuaGHUOqsJyuIrQ+ejj9LQh0fBugcx+51YYVLkz
q7kyilxe5faySHgra90J+qYNNhgoPNQ/B2PQF6TXGOM0cbySWdcGe/qaakxLHI4ZzoVnNCeqMHAK
F4LfTn1aytdJClQo/IJ5TaHUBUk+6brZybuD90NFk/OyF9FQgFrGlkci9TElE9bSDRH5aBO09ZF7
bGtpdFtpJhFTjgv/AXb5I51/6LIqNRq1X/HARD5/kQTpcdDwdji2mCEQG5ho9FVieBscIqQOOFKD
tFAMI27lqiuxfs9fbTSy0cgeMWm6r6+Dmuj8HqCUk9/JKZifSzqkB5fNb7J15dhsV0/tzFl1tS3Q
rjClBmr32grdl9A0b1oLGBLGvUFc3jXDHD5ZjWwaLKxkcB7GsdMEFAoqkmYDGaQd7SpkVXnC0/TF
3daFiMhBVpIscs3+Gh9sHbCgmhOSqzeT3MWcw+Q8lbLP+pigoRcCH7kOVF4M6qevehzX7bV05vTS
EI9OrkR92y4naRv6DnTTtp++WjfV0mKRajnhQSjud/KkrBKSVjgvifd99vcOmloO8NDyAGwGGhS4
QGePwJRAqozcOv8Iam6nFk2oVQVwY6SVyDa5oY+Lj+KsZ6++JWoiMoin82NbFnpI4rtYVAMIOaC1
oqmLtPkYTzz4qz0W13/VfatjlLLEX61mXChJc4S9d8mK4PMoA+SeypiXZyzp+DUCMbd/BDqJdxZs
0iCtAHnSQ3e7PwhVQYYboKiVuDnXwHWbSFp7gH1f6bPYs18VUDxQqpBzYnqp9odsLCAFvKww9qJm
VTp5V2lOI0q5M/yJYX9QvDElcjTcKgwCrfjDqfxW/BLK5W1P22pQKZBRZY+i6GZAnNO23/aer2vZ
1xz78xl15PA082DvZYiF4eCzOrq+kR43+h2qP+7QSf9Uw1mzn6/h/lVkw3n189idTcWylg47ZDKo
33gIemd3pOpEDK322znbSNScOukDKsWO/l1SlmoLZ4zY2HrzrelmmsI5SSnW/9yMnTxRCtw77/K9
TI5ezNZ5/G+mV6C+8IgFHrBnZWFlX8OsrvL1DgCcFKRMvflxcAO8NR2QnQ12+nsSdslh7s13z/IV
Wq+ORV6sqL69kbfnzUzB771Z82x0aVx/7eHZNdo+HM+QL0J0p41V9Lji7sNXdbJA66vZcnwnBiqf
WAXQSSchJ2mvU2p+4oA/zEufRDBC/+bFSPrZWjWMeGyMLAsN8hs+mMyqB9yNiQdufJtddSB/DTKx
KolVRwYGgT/Sm/Q+OixANRJXHPIq3m+55PyusngxWmgBvC9I0Mq+fy8YqBc6W53L/mJnGfwPW03b
P3po5KtW5R1cpQn35XJbwjFEH+jCTA9Q3vukI9MeQ00aqlP3FMKJtxB3sSSeOutfG7vLEWFlcnTu
dp+W+Cj0gAtneRHLBGDk3i3gh0d6TqpaNWvymlkQrErRONFo5YJPvTp1InjT13pjSbisdvIiG1DL
/kTdmAwl6Fsy9OCOuDKMs4RPjqPSVhAzFW5rpSkzPIs2h9HSjtIfqqqRqQmeoVxKbXlB3fqeXYuk
oCLfSwVrFqUzzHL8y+BFlMxo69JvfCujXuun4lX313b07s5LsqojHpCO1ek/+zDMuoqI/VCyjd/H
naOrGC5Ati2EhfKr97xgVO5HkVKlGPf59AmwhWGzsaI8TVKFrITjOCuXNVFkY4gMLVVcV1eBktTk
4pUzhfus4aCYYKv1/zkp3FsYmwNTRPbxv67aodcOK7ie1qBp9VtakrBrSqLS8dLeuH+RcsNEwnAp
0aduT8lF+Xi2tdF1yZNc72LdpKSOf08g4gaJRwuul0oezihnQowNdDP+KBVq9g16eDFLx3ZFvubo
ADMUZURVnyW/+MV4mM6Wl92GdoNr/peVD/I3DNqAO5aWM2Fd4hL4FXCj8sr0JeNKjOwFipr1/IAH
S/5E5F7+ANnbxtmPaMaHiCIGDZMLBS1ICDDfhqmyOiTRyKfVDvlAEAF7psJOpUuoa03r/sePFJ6b
/QBoOgUBSSSG/SP+U/y2EHpalDZN2G8ZasjyhalQqhvMCmufUjjqyZvWKv0I0R0APH2IOD2lVx//
52aGPKpsy8rk6Q5KEFVpxVLdi6xCcWav9YRhW6fbu+Bbu6BZkmCE/4s96j/EPWOwbpTywxxJHuG+
cigu0F9RTZQssQIB7uZR+td5BD+hEHs6fUUDd051OOxloDMUDRyH7cfYt3M5aRbhxYdJrWid6aFG
DURJG07JF1nrSNOsDXrc8MQVUhuQiFCdmWZsI4JwlZDT6K1V0//ljcRdKZlalM+P6Pxv7HtzoVzG
Ww7jqENGhvWee4nbZe7a/GN3DJ6tSVrLZeh1xqOqkyUsLKc1KOSw/7h8y9PYRW6SYgrBOpYrdfw6
/PH3KTLgMxDuGr2IEZ0fWvgwBUcVwh58xfhOMa/PluJVQh/CbZdcIXEXIKskvwnGmNZJiUjVqfIr
NoZR4t2x8ti0TdJ1ZcO+QRziSglBpLUHrsVENvuNz+lR6EonlNjvD71q+6tdvcnOytGNvov5Cl/N
GdAFLO0kWwyDUIZA1yK/8LTkhZPmrbEF7nBnNh2SFQvpsK3IhCRE3mi3duI5PqkuFyQ3IpuAl0Ur
dwntcEE0gWpBQlrrywJrZ4UFLFCdhxATbjnI2n7pEUIZ8ZgAaVpT/vBIg+D5n585et/FD1j9WmMI
/7B11B6YGAnQGcWnBHrb2hs+14wwBTMSM0iFXk3o91nBVa5ftsMubJXpddqgze3y/J6ZswrXjIXb
7knYemIi+q3da5icBnWOa1enwxvmyIkrNtyPQz/LLjkD10L+Uo3qahxU9/1QbC9phfYFUALf7Gjh
Q92Aj9j7HKFlM0eLjb/5GAYRPPaXkW0eRd81Jkh5ic3DGWuao6OOnwextneow0qqyT3IYT2MBKPS
5hbpRcWHiYjU4+nhldFx9MxvWFZIzlGWHBGJiS+BqNJ9zvf3sWjNtVNxlo4DU5MFc7TirMYjmo3k
Oj9hU+L3XRbSzJM8RpOmD2LLnO9JaN+WmUgRv6WEktOHRsGMZWS0aPodStQZ0OM8y5eGs37HyVNl
pPQKsFe02u6mWK+rg/1RHmGtm4hMUfAARubZZ1/p5V9RCISuwdnxmowbr8s815ftQ2nJt7n7H9FN
ada6NSuFLojaewHjtNrSQuUH63uHd3AaJHF7UAxE9rvnB5LG1TUV+zF/7bA3sfZlLvNKBGW8Aoq+
dASKR09t5ymVzRRzxwFyyj8FgEjQXBhXPXGnxsidZEx4kkdYjwaULwadwqYs/kJ3Z45S3+v/mTyG
eOzp/fNk4JgAe4XlLYJ1zNCqYQETF13xcQZMgFjedBM1kS9zCjgjCW9wra/jLWhCbzmi7cLnVVLN
03jHv1piRnGWW06vql4k8RTLXeiYyXKoGFQrT3SlRlb7qziK6D8MzZ+Z7GTTTPNKUT6W6PBkkQuf
i6diD4SYS8BDrb7gwRIUDPpshciVxIHYXAjhKfz0/DrvG2DH08XcYURGlsbYyXnwkpUJGzZw1dMC
US/61rUnRdzaxunARrDkP+1Ne0ZU5mJW1/BVglLq4oNtr6a70E2c2kzaKDvhp0hO/Ana1sYlRhAw
F7+gKQ+siuWAlDr3EkmeOZ44PG04AoeK3re0WlYC8hVD8JQLbUICTQAiX8sYBYEzmrFeN6MAHXFF
oyqtr0fx8Zllffx+MdTHBwlqLLoVZ9mi9ghv1OG9QFJ6uzNWB/myVPQK0bRBLXhq0Esjh9deMK58
ZuVxbJmfjo659ySQ+KisGkw8Wa9TPFhvqfDu5WHbpp0o2HAtTT2J7JEOcQRLOVmsjEOVWhLw8N01
foc3IJu+QFl3/nvHGt1+U+Gd1rY+HO+KAmDzIlrH1hHAVXh2qTiaYTDc8ea6/8VbJHo5TAtIgrel
iiI1c9luZHl8JgJk2OH4+mrVCQZ4UAyOUvUCqQRl2KCrrbSoDo4KoB3G2EV1h3FJHD+yotNa38+c
QR9SpdlfMTUFy+MR9dCv27tEBqmamfEEECTMxpv4EWwU3Dq5AkinkX/XBrooR8XT+eRO31FrRpxf
isYKv8T2KdoNA3w6gGFQNR1yfFhdO5wLATCMG+g1l3DzxmR01SFE8Y02ltujqpxOrdOCAzoVxiFR
CMB83SuAJWSsJX11ieiSrBPvXt+VRRJjRfnoO4+l3nW+W/rIM43PQS4sRf/BQnDCJbfdn2Ap5UUk
VZ6dB9gEv6m80nTdsOLUBPKd3JOA9qsn3mmTVfbZSYTOg59yFaZzoVTQ1+XLgfkmxecwFlhlDjwk
oDHTnvoulji/Tk9P/ZR7e15ODfXht8Mg01Xh4FjdGs7l+wI54WQePBtC597PLrMzFerlXrfl0FSb
QzYL+TJj9PkVSilFaEWGkqJ4AqV0y0PI4/BLh4DTn2Axv7msbmHeUE0dwOT3ck16G60kt9xYbZvB
DKhiXYY/LbuBXNyuEBNsDjWu38Fog5HooWNmtOchuWAOXzkppZ3Cf29kedQoA7h3dcg217yHJPGG
+XcH4asWmzjOK+gzrQTaVG1DZ7pg6X6RjXvL8S079Qp3MDUprEJLwexwgiNwvNoQXEfEBeDp7DtI
93w9vo4kEFl3/BDj813TZ0hXC+pmaKAHBJOwDWTkXKolnlI9LimqtPgdTDJv5oyUBX9DL8nVtWHD
thKXPZLrOtnKw7qjgRN5Ki8jIUzpMxlfteS/sPf3RuE15kmhzt/DYtzdIKnYzzEGNp9R4eNLgQvJ
bLt1qbLARtSa7o53DAzyvVwfC0iCVeTOxNuXu58qEc1MDsjRwzhXYo1ZV/6Kl6k8erF9f05Nm6pf
soq+GNmof8i6MNS2gYPJU+4Oi6zFLmhZ2NS3lLr74R5mPUGefr7ayIT3OJMX4pr0uSJYm5iO0Ted
tSGJlDDePLO2LTk+XHRuWY6KuDcXJL/HGHSmsmiUehnXCnzMqNbw7mhyKVLTqLclnVSO7UeAw99u
x8FpnXb1Qzp067hanj2WzjdlLp/ExGC19mnu2aHfMd9p4PNuWPzko511aMH7rL96uk4RvKhfqK8+
xjSVqvsOty0PdqRaoepAbQ4lultC/LSctNwvdMsHhM5J+eDKr9ZRLWUmrxUnCQc9BHM/t4jEObZ6
Kl1WYYgxDWsHK+4DO6VWIZtJNh6bGLtFtghgdAk5luE5eiEErlJiUPRtMvQ7h+pv/VzLpTy/PtkF
OjWtmpsZqloAUm9By2zjnTrmJ8QTZ85laeLW5rluNlSmGEgUZ4JldE8U/hBcUQA4iST5NSeDqs8l
opZm5NjATnSLNIUY5oT6bso2Qk2e8u0P5+4UN2ugfFbOVRbpoLv7bA7eMFv2wtYohsnpBEWGBL8T
96dFVoy6yQQzhgr3msBy4e2aLLkgqEtNXrbuGESsqz1VAwu9/UjB9UoPD48lC6H8Z/6LzTFoGP1c
HUiThrfQ4qvMgFb5xqOuKsIHIi/DfG8QR2Yqgas93qlBO5LjEjYtytx10rCDoLUsghzjbX8Pf4NO
E7j6tmNO1q9GPVJEDx5Qned+drsgsq8KoKAW9OWA1g6cmr+rjUNWrRoMbSB8WUpUkOGOkZL6tZ2z
f+H+LRTTnwY7FEDYf04fM75w8nuJLTboZOPnD7NZY6I9p6iH1SNRedXiAaEk0tQDDRTlzYkkizt6
9TbG0JQRzSi0e/C9dmMnGpXvwAqzFaEaADqg20Dv9KhCAdz54oA4aY50vsaoGT+nMHHQCwkW1/V/
iHlf3Ah6lUDqrD6h/36e50zQuOJGsWnnnX0FWVF5djxAwcACOYg6+POJzOuSfge/rXLDMkPj51UL
sznq7uzatYyJtUSOWa2HiI1oexoof1AoQJyKXEkNmV0qVZCbqlxhqTbHnJt4UqOft1RyZXKAkPXs
l1SEtpRHMMR6LZpEevB9gM0iEcqeWAFVFATTwAYiiBAjHyyULyzShmKUQzPgzFjs+G4kYNxoPto3
2QvVMRDV5JVCKajGcSNgexLvYcDL4oAX8rhneaGSitd5eX2k4JNXSPvoQJ2Dh/HpVDaErH6sKLMe
rCOLKmxfIxfP1H5uiIcr7uSmggTcx8JkAKdM6e0wEx44M+ZwFd3vKnlTDPx86YO50v4D9bK3ZNKU
vBfX4mwxBnnRMdNuQJ+rJ9yNS7hvX4t+XhLIap0WQlZWQn3C3vt9mnvdzv8VdJN4fuL/NNRPiXDY
bby1mTaagzVGqkJa9uDt8sbT7kP0rouYvciwwuwrJ48GlfrbkLtvKokEsGYj58DAcMqLaEnYnsSF
bXAAomVIVHNzpnWsnskK9S7WN47+oj05ZdnFG1cnwesE1+wrKYNmNUl619HoefIdDPjsHzc7XpGc
v5SHcnSTybetK1+T35LNOAV8S6POPMAAQISSvSHGwwTvBMeEhYvOmk0USdvX3e7jmqPVYY59I4gJ
62O5eZVICpU+dKs+xqgPJL1eBvhZpfR9sB3VB1HFjUOXlrRwlFAAWO5TKsPl542Ih/pCXN4QqceD
AxuZGbEn0oI6+jGIqXfnvkowFjlcY66CHxhanNh5KuNOmj15jSMu4qsvDvRn/V5/725B9+W2R++G
phBHSuiuQ4xOcNP+LCNUwuEMyu2a6NonQnE8UYnuBRW6Eg05yItsrEuIGFjYTq5sJdr8QofXIVP7
nKPEMxBW/2q7zl9PVDfxU2JpqdFK37CEn/ArKmsJryEzot8PzdYkWmXZmTgKHjJtzvZ3um4GH3eU
aeNJgM/NkDPHHqwIJXyW9Z/MxObLOy52IQc4qcNMO8F6el9HmMR/c+C8TXbOQgFFyT5z4vIV59w5
Va5SMp4HoASVlQW+UhsPPN+QOhG0Qae9r7IS+u8QJBWEEJ49xBjVVESig1dDwNu9uqzlnTYC+ApV
ycbQkSdNX7gHYC+4rxJZ60XLrOx0hRJNL5JqIieTPGcqkuy2M5XHFcsc04AolwnqP6kVmsNJWgML
ytZkAZDD9mDdh1NqFKzfYA4aTnInV8tkQLA9IOylzZcWjao55qdCHV1jyL/LJSNGY/q0mZcUPp2K
hmbwkwX3ViIxN75kylDBr3CVN0Z8VBxxNCAsoB7wbLeQc6WIEA8f8gx5qxNjsqRzW9m0xiK5nRa3
AlR9iDqhzckLgtIzTIVVESb5GuP2CfEKvpeTgAndjG9GVmdhYe8v/qbsDhnKXHdq2uWxCaRNkFzs
jAO83b5A8XCWyqfYPsSQPvMd3Pyyon69cWEJJPVzjq+xvR/xiGXtZ7XkeCV37SHOMKZbarfAH6Cl
+SAsxyqdUWMMLfRRfgXk5xeJZDkN9UhkKxWc4sCMPTRgk5hmp+sTOdb/BA3E63YT34GwErd21CIt
4VqQXgmmDl/95N0FRheJ24uqiyU7dT9fgejFjxbfSD/u26ue1S04XDx9+FWTHRZ0ghO32HqTDvVZ
RcLOVYVcC3WKzVTDsqJyuy67cRFANlrDoikZ3UlfmsvfgEj94oiyxHOCPP6tLP8SJGXaRbqZimIe
CbBAoAw0jxbeLnI1DiWG1bFl0J9Hq5zmJIcqlKmhSegZkZ8tO+wwDBkL7nVn1ia5Ivz04V225nse
hzwu3FhQtzpzT7I4pFADwxUKOLXOgU0+p997QMsgo0E7KfJMzqncC2141B+fdGMpP39btAhA8AAJ
/WEtJfecuUj7Z4tpOomVrPyh+48kkRb/+672FAoXU48/9hw0NU85pYoY7yLM+S7UmwrWNfV3iTp9
JQsta5YyIBCvxWynF8EhKvRg3KNV5t3sNDt+DRi6Q5dt4OMMTU56ogFMumh8rF++ERcRnewg/of5
dRRPSblwMtvzzp9MfcK7A7RAaeYjwWQ0hWqgPllatyNPAnax/hjz9k5onn/uBNx73ByK2zlm11/F
H0CbSWDN19jv4WcJhldDzSkfThLwV5J+wj4hFjKT+7Bq/bNtIYj5DyJA4wQCyIlHmZZpUEHsphL0
ZMLcXV9jLtcI/oWA74ahkfQedB524/hLPSbYntDUap7ouEAmABjAvpgiEm5o7qbvqpVQcIYUSGyj
I+nPaPrJoXuOlHRmExfJ5/naWSV5473cRCs1ZSww+0rL8G9ot1VIIUy2PRytEhTfwxwqxV98FErb
lob7lrBoz/1KNWixI9gKpOOhl8rqA0lGUB9BHmc/V6EdVdMVGjD1DH+8T99JZaajiiK0oD9sMUJ0
NxPodWqnm/S4OC55DtnColm1K9jtOhdNqqRW0zI2eqYDfbafCh24m4fEyiYWvjeKYAQT38aXgJbP
GHARVf3S9VQnztnjy+Pa3TMWbenzzGfg64d9n8tsq2NlGNOIWiHRoWqF5Cu2PyWCkZ0WkOZnNZii
nrzJE7BcODFpFjXCiOFZsWvErK/G4gL0MkFzqc+cJqyZPta1NzAHGQxaOuO1kBA3g3Xuxdit9LCE
MW/ow1hTD0z1mRrjkHXq9m+kDuIxubAQWi3V7Xlt/D+QE/b4gq01NQePuPL87hMmEo4wOg6IPi7p
uZA7AfqL38KQgFjYquHBhekaMTC1uu1gvLT+07pXMNxw6kcenF5WxPlBQZ9rks53fwpGp43ZIpll
Gret0rT6X6oGYLfKaXOCqwi+8xmpNNwTa24P1v5M2Lpa/u2eptv+Jho4DKOzd20uspcpxLQQSORG
pEQGR/U+xggIU4KhD7a574U87BWCoak865eeSqy2Xxe9LGAtPO4pRTr9El8BXQV+QLCugLDIqkNv
Kt/LEeSRXQr1zC6+R89iaq+FIsoVyThKFyOeMpKanOagCMA6KHNBHH2RFee0WCJ8GTVQDkZbIxpd
n3A4nPC7mTY3EfGFLAGP+7X8IvOvpN4x3Ty5msOQc9ZIE9RNB6jtmNW+aBFJvsUI58mXkcr4FHdC
HeJzHJ7AbtHA4CDbAUYAg8JDedOS0p6qqB1//dognDJ4bU1aD1Cx9lD+tAVPCudFOaTanZHqWkEy
osJcrWlfKJrnoKDko2nzEexC9DzcN7kS4XgJ0XYzSyqIDMNgRG01DGZs7Z99Og6Reoi6GBAF0ZQf
loPOLBOBWyII7Ky3O5YtoMWkS4Ec+kqFaRtgVLDln7mBtNrQDnfD7Aag65BkNePsoVY7zD8nqamW
eyHdS0hHyxLF0ZU/eAmqF6jFU52oN3awTaNEhkypWunLKHZcwgPGadKWo7uIKAYGo6SfFXTAUROr
agMmJqOq8Mzin7hzV2G/+vdSbWt/j5hq/hny3o2RLVVoxiixv0fM2Eeejz7Yl0cIrFrOaxxbEZrx
Ed8UuhdOpgTySd/syZ8rahnMSvX0YnLBfU1hQ8okutf3fbuU/4UJyAilf+VCgF2kt45CxmKDc/KQ
VtQvUK4OPQmLi+RCM+IugNc9Zdkcy4ehC1vYuUuDF++qIWlo8Y7hf4e9MnQSh0vvsg1vNKMGTFMQ
7sLJRQBUaA101kC0G7cn91XaLQcehilzva1zd3x/0X0hJtYMvNbKWmQOhEuPaDY8Xn7mmYW6a80d
rCbZRWK0pf/gVL1ZUCG6D9zxXH6WeHf6jJNY9IorEadz/7FQ2HcqtiKaWy/ag8Ur6G6WH5rUn0Ry
r5V796eTNZRSwF8V6CkuALmomN5M78+J0ublTmPlEzCenxsAgVYTCxYn/4osEVwj/Z8oiH2owumi
WCbeNDAfEDabRsx5z+ONaTkJGnjIPjvH3cO/4PRpPojCkvKtauWBdnt29g9gu1QbdmriWGFnLg5Q
h9/4jf3EQAqQIASqE09vA7oMkw7Nq+jVBXucygGyXRqt+jLKEgsqcijoqlJbmrN4jcExXt4q9n4t
H/jco9fs0xzbTMB4u/0c43J0EAAUKplJjR9pGuEMF5Ehw/fq4tDVG+PBMXgDlovLc8hBkxrihBbI
J5LxxBSDCv4ILCKTcfl8K7UFEPyiyIrg4FrVGPtpSegNBapefI/3cx9D84biiN0aLah2sX1gsW0r
uOHBi16WSrX5hq+E0qMX5L1IUX04gRe2AwURvOUSKA+mLaYkeERLGB33ujaC8KIPhvKdyaq/tJd9
PCy24xEuSFkvG1SJsoI3Ncaw44HyKtU7VPjYOia/zcEGvbitw7m8P2MpIykWHVo3Iqt/0/yQeXAg
3owiaK9G6upLJ+QItVxcx3Fx+JgYEimBXplZiGUdsx9OPOREGuqcf3D/5LrJjpTEGhYkRbzzuAyY
/mxxzHTM+qpkbZ8i6+mc/dWmQx3ZNl9/TemuteHTqWSJAJoqiFo3pjvlrPNqxkmN7wQNTU5msPuz
170TPYL5HYNK1c4nWGzDCs36n1xO8L1fE1Lud86v6pTgy9jwoYjKESn28IpUgWJI1Qirn3LM5tLE
GjcC/vTbuTXm4GJ3laGF2Gq+u0Rdkk+J6tEUoFKklsno9i8+xQGTMqDQTZYgCExf5crAVIgQIHnf
G+wZd1dG5QPVnM8mXwfEHPm74LZrtds1LOGWCZR1f/iQy+e8GGe3VJ1qMzpBE06kPLaWKnM+5lPv
lXErkdhyx9biXXAm8d/DWKWDg2nKH06NxbNHCFKXbflBO2A4Z2wTSJsj8UbhjJZyfQJbitZUxINh
fzgvvNH8C5QPsToo0ZPeflvYgT20w+YUO0LybYhEhyys1KabNeso94iF082EeKrs68rVqioC3ZIf
rCn1/+rXr6wm4Pn/wUrybbXye+IdsPPZcfyUiPZaaFcNNT7GwYw2NB5nDc5Ayu9QuAeRWpSwZRxt
1biuJuszvfjw8Pdg++RX944pICvoUitQcAruuVcEqYnjul+PvAb0ag7gDB5hIVF9FXIyO1PxntSh
dmLDzikB26V9bwz65CDX44fjTOg72GqTDA4Sx08rTke4Wrz64btVoXtoQw5LjJIVy+zLmR53CFPE
ORLezQQHIV8IIVSWetnN74oc4s1+zdWB4Wus/HIPuSV0Dk/+L73xlETg/k9Ily8U34tpv/0mZ1V+
VEu9rmFUTH8JTas5+71a0KtzpvUq24WJPIapasaQJkH6qIM0NshtEpLjmgpBwU2/pxo3hfZoY3b5
HfK8kRvL492P9cehh/V9Atf6uqdluTTP50x/NakExB/9oHIH6eZHxgynCYkE6NwEOpUZ4G6YZHk4
SAtQqQ91vhwKEDQJM1AMYmTEBCOQWuf11iqy5L1h+q5m7u/4IpcqRnmZtk+8FwK6bXSQrd+1zxRJ
GOR72gd0SpTzSy02tkYVoxvdg1CGrGPZe5qOJ4nV7WF8u7P5YL9UHqVcyBkyyHqUsLMN64DwInQN
hOhm0d7gPPVtdGPX2iP1mY6RVj1edmpXg6iZETt3fM+FAfFQq0S1BoaxIljBiko7wW+s3exbOQ6H
oWoGjdjhof3UYJWO4HI5Uq0X2mMN5+Msd+e0GLt/6VS5Qszr2XbF+6yci+EgauN9njrxQ9aHl2Ps
74G02Hq9aKPsO0vdwbl1u0F7ydGjvCUXJbYLmvzGw6JaR+xeeM1MD/lKEflUxwXuB391iTnuUS6q
dyDlaCbOvtoxYcwKsq8jvmHLqKMgbqS7caikBipUz01/HWk3Q4KrnMOXd0PLm635Z0Eddd6hkJKL
k4gerETdfhz+32oBqjzutxo3xBvVfuiu9e8MLUHW4tHwDxR5CtZtain4N+PNI7bhU5dwSfyDJWCQ
76piIF9u/JOt03Wj1HAvZW20Rf+ODuzARJ1yFkrKBKz1HG1VQ+LEa9t/dTXZbOymT0CcWFDTwAQ/
7Aqt9MVbNfdSV0WfEH/kB5vP7Rg5sIv9GUBkD1GkpiKT6Rsr4i2omuk1rkhJLBcepoNaTbKnZS/m
1R5SNjGozMRUStq7X9UC2fxbNm5phrvTSVVn7k41ZhTJVunVjttO8vAQ/qO6Ax/FFqgjvLg9JTcz
2gvmp1aX2UEyj7EqrSpnphitSgzPXjo7ej9xT7ieMmYeS90QovIF9OLW5dK8wlC4vRjbtqrr5l1p
vZ8DEsIIoAc79haP2QcoC2Y2mXrsn3vPM+c0du4lOBTpayBUyrAH7rqQzqbSJ96DpuF3wOdzTWdI
AKrcEsrGnpxBajrWWs3frB8mD9pCEd87IIp49xS3fiGbLtE3Aa+nqceTyoj29i3QA34C44RF1Dl1
dNmGXgnj4NYMfvaQ9ADiVWCnyyFpTBfyQFiVJHHrkW8SYzf3SdCGqRm3DqQeltNdFExltSA0/cju
jzMm/QvXa6Lvl1kYOuWVIx3gUKCyhatCk4AwyP+wOXCCGaNbqJq0zBii5iIxjnzBXGJR6yvdX2tE
J0aXeP4WC2sS3nHBVctn6P4Hjrbcy7trAUQ/7z5+gDJHfy/VKUvqM5rCy5Y2ix02LleSqmWP+6f0
s/FveKp03eLMopjd7nJlKiEFxST9yJNgg3EbR/8wrMENu9aOd+nzKgwOgGICUSkyYZ2lIpOy6pHu
UtK5TyWQuaHdZS6tHLBRhV5LzpIBd0/sG45eGN2kCkflhKjvBPHXZ81DSZMxiZ5mr2ym0hEIHM6v
uJ+lVcrPNXDRrMIc4Osnk2WPffFF6J20x8bu3JAfqiW/1O5npvLWoCnwt+Tug8LO7hqKeXMyzDEl
hsbgbcRdiYTOPa9JPSkpMgd+0pwKrHO3w2LdXey9xiuYZr4QfqyxT7TRTLKcDXkG2EmoE+HsbzOE
+L+emQRlLIOcHC0GorNr6bqAojA/uZAnNjO1yS3JaAYpf4fa4Z3p39CyCFjlrWGldj0llf1U20j6
sOIwXTPeQn3UR4xa6Y07QWseN3SFDUh8WU9kis5U4/AKwDtL0VPWzsfNYyp+Nq8zPZisWv3T+roK
4XWN6VSbgEd5OIdrlGSYwiFJtv4w9/C8kTmzDyfDQZ/awei5ci7jz5O6ge2XYEGfhyTDGsbtwv8Q
yA6SfkJQU79q6xakJNJCA/Afhb7XRFlZlZAEmPIOZF4n0jZQ0VGvk2jqxiULYtA3K3HUNlOph7mF
X/9/dJXx5B6+vb618eo9bUcKS/7H5N2qPNr91DCo7TLwz3KIVMXjlY2ejbPcRz0i8rOLMnaIlQca
ut9tCAgOgKcViUQvrMQq8Xp8G2ZGVdiyiMBmNOxc9Y/SITqC7lMZMuq2ww8KPZdD5fzXXlk0ZtSE
efpYrFkiykyIb3DaqQ6f4tEGKyceAQpBzVtjPMMdc9OWvBcMdR718yNqW5YxTN9BmppDJPA7atIy
PiEdnrLnYnl4B5v56ikguqFnF5mAqhOjxDBFKUEesu4iDbFA4bSZqGx7SCMXznXniQLQNb4P53Aa
Ql5izPpuH0kQJP4O7NRbsWaFv8KoRArqWI505uHh20CMNG1r08a0B8EIYeBGzrHKLDsb6GUkIdoo
726YgrUBUm7tapK7519KRrZGUVEVcoTyJReiqL3wys8MiwdoPciNY9uoUyaTQInWuR2S5CuXAATS
7JTYfs8j23O+rsE02e+AXNY2DS7Nlyp7vlSpoIwYR2oKbh32inimFwYfPAeUfX5TR5nVE1FPqNgN
cZHbTSH7bfhw9+ZehGjULT6B/SFpP7+HEDGQtMJjxGbDL8QIDVU0VmM7xjJlYLWi801BIMo61TTG
9XU5vosTl/8CaVE+Q3cRysNmjjCkLBRlcyQftLpA02vWEe21bZtzhp1zAzV/2P6B8oZYOG4/i/L0
c71EsPxXQ7o5VnO5n9IjJPPJkjegbepNzuczNScTEcO2TK1GZ621DrbVUWcCFC1E8kRxdxIMuoB7
vTvnKTN5si4ak0R/ZDBkP7WOUzqqy23mnBIEqbD0yWbyV2SgDsW9Ur4LjPg+zPm5xeynCasbeTq7
klrzKQDo07Pa+SZ0mnAEKqe9Ud0kUd6LgS3Aj0HBH4dWBk8rc6aD0opB/lCzTIQ5mJllquuEWfUr
HSOLnYBQiiI5npIHu2Xf8Fwk15HI4NhLM6Gn5gMXZ3bGgIUQyGgTkQWW/YPn0roVBxSRQEgpbKXU
+da/o7U7Onvvl7m3Az6LYqAGlwFA0BnJ6cBub/DM1Dik0AK91lhbOnmewSeUQ5wym4JgYTIOlIiq
lWWaHl55QUd255dA/8ERzN36x2FQxhTW2OkSAui1XQya9zihKXbEBl75vYpLNkG4C8EQcZwtKIPj
yVE+s6fFPAQKrvfoHVyHHSg2sIae3aPiKZI0js/Iw8HZuoZvNTC+43BoqxNCRUKm+QbwRUbYmOjT
43Oc6ObnnpFcP67r7LYEzeKxGMoAS2wTJTiOHsJLYdy2W0hIg0bfWhhuhj9+qAt/1qTyrug82Qg5
9HmUou2xmlpNnHrDOX5bJav1s4o0wz+RzAppZrY13vbt3faNhAfsMaRZgDf50a4iLIB/FKTUb3dW
VY6SEG8jmXgIH4g53TFcezdFqwZud9ORqk3UrQjgHe9U9OX+1jYvBXC2yN8GuXJ4Dgg8cRP5HXVP
H1nXgVVu0Ep+OQ3h1tS+BLCOr6CdIqTXrH81HiscqnPY9VoEH0fwSOFqYDNg6Mn5rT+wqNPZGt0n
F1RLJN3yti+ci0PjiQe3woP7YiszJ5l29IkuZKcZcfMQ/Q7Lw1E0tfmMvfceu5LQ7COUJkAhZwFv
SG5qVLgv240hjoevesQAyyIIbPQcVS926nVyg73wOoj1ZdIuWKNq1tg0nh3saVIf21CQJ4G5h6FW
WpZbCpB/ysMhN4MN4Q2fiwZlZRZlnggy0MU6FyorLiMuuoCADocdY1LyTI3M9L77rOodbRkbbOX3
7YTDIVxK2r8VcDMW/CPMs+JyQvNqISyEpCB+C/dCGNmJDwlBwfXxjDvFpHADQz3CgC+w12+Sdikw
pk38MV31nO2xnQKXcwFI3TRPpHzy1rpsQod5YaNEQXWY03E8GAsSFs45hiIiRGsH2rK8yIx//Uo3
0V51/ZVX6aF+8sf78hF3HhFdZow8oLgjRYz4VOxIguj4C2gYN+5Fo7iEOxZBC7F47CwgrPBua4PT
u5IaiI632DIdwjAFLZs8CbMaX/66OGvQELNGnvPJhaqjwMbs8jwzShY1pkUs1vF6Ns67xKCmG+o2
ix9E1tgPPsnD9fk6v1CJiZGSTiBtVoDvnIKGmbFn3a9DSIEOw7J6kbnsJoHCFd/YqigAqfqvFQ6U
dcwn3Pv0vBYxwqS6pPLTnX1CcbeGBYk2+Tkg+fqbkQ4oxNZh504DE12wnPBqERPtVKv2UNYGI4wU
nHCaeA4QqZHF5tlsCkF+D2mpYmB3w01oSChqerrDQLBY+9RYYZPTW0dSJpn/7yq4XwN5Uglm/urq
MiVW1kGaSN7SD/RarnsxoKoW3ZrK0dzx+FfYxTTsIZPDnQvyrGtk/1VtB9sRDONubc90IqLtkFHS
b3O8KX4rpl6kLLW49QNqeoJoCCk1iQabF3YI2LiFJlGKbAT9eJfqO+gn8uw1Cvq7FhqYhMSw/8yN
w3Ow9qt8bwKnIXUCqAmN4GdXkbcCTYOA493Ch6CsxwHiFvQxuVaPixBsTNn5EEEygeRVJ6BDanxJ
F4tnsyvE9JmNB7wozWnabRwXNrwSyLYW3IZGcS6qniMS7WTIIEB8M4lCFS0ddlUxspzt1F1t9Uos
+Zt/FYQuOBvRptuvqJy6fWCBT/pwN3HXYjwAgpkr/pPHUqwqg6PXL9DYOTXc9CZIEADTDXWVt8hE
AHOh6POhtwBp07lnTF/YgLLydUbJFHlgpYDk+tEUiapnRcBDZllFy5GWwzM2xgneSotyN5uxAeQy
TCkkU8NgKCd/1okhpcEu1UXxYbNMZds1N2oeHg+n3u+oHNGX3bIdxNsWoCu4nsXY7Azxao0f0TlP
xxNArfZP1BpqbPY1K9KQhp5sNJ8tOpTU6uA+C3eNSY3sCBFQ4VrSEKdK4R9Y0jFSc+yeg44XTWGj
h3155kPSyMxnbYYt0HLqP7JLykEsxQL/HokQqWlDFQ4byzZBG2AqzdctJVd5GACG3tEi2VSySJ1G
zt4ph1JC/WI0DWoj30NDkM1nt9qjxKKEwGChWsIhCFJvr7hmunPmOHSv0qaMJKbA1MrGl4cHIFYq
mOyJv51t3Pj8PEl/hLkkoMoylseRZ4oNfa3wp1Z+DrQyri2Ssi46voREIb5fAJ4vGeZ+4UMTdBJE
YIKR8YyOovm4WY3IL3rVs46vutbw32nwyGWxIsIjRli2DdGQ8WfxtJf/a/Xw/LjRuKBaU3oWAYDn
5fele3UWvI8BIfqH2UDBBXPIw7FDed9/KgAaZVFojOBEbhNJsJzhfO5mkTVD0/FTnKT4cW5Z5adF
AXC86ZdvHbCetraNoRYCyc0HdrTdStkB0vYwZIBIDcEA3fhYet3VOYWz/jq/tuPtXgKF/ljsMIbB
D28vLnq5dzepXeIBpWAR18yanbkxhlUJ1YGAiqxuQexK0143Voy1v1iBnNxTpCVk+paZfk8etYe/
KTujNj0qAFbINCdB5ZuVR13FULudDph5xuStjA1wm/3F0KPtaGa/HQuhxj3yBoq6wiwXeUrLKCr8
BsQMeFfB1WuXXmtXtpgyliq16nxjchXPv5+3VTKUokIBh9UsMnM3irnrcRe5cSe60gpZ/3InJqGB
l8HjmltC1OHnkwr3DYFup32AOntUrglpJTZ+01/Hc4+1kNIFPXXZqS7nLYnR7gnHIKAuTnG7CVeN
dWFNFFUnfWSoNJrQVZ3iZ3Fqz0pxuZ0r07O6ne88m0rmfyVTDLaAStfFpD22fIoYg7xKlLCkgDH7
pZ8czDrY0uqr9do20jCMXPpCRZyGwseuGTvqG1HLaOEf3fq0Z6DrbaMTGPWfI/r4L3GHZh1G2gXY
tBhZsqFLxorLL4WUYc+il5n6+whDlyiO8bKEV+G9LIvyNzKrTmeWUOWSx8VfNAe1btuBwSBLa4Fj
0d9AvQbCZpqrZPzIF1336OKhOi/scXjiayeZZykP/OpFLNdBCNvWt1+TyCsC2R71ZlGs25MSaGcy
TjTDNmp0qHWloP51jve89ndiXq/X0S9MYc7bRff+B+lh9yfrKXjQj/NA/+GmqzxV/NMC2oWAur9+
L8u6X572BIwZ8YuknMmJij/1HQ3ac/eyvEgZR6sl0mIyxkGOqgoiYYx1DKJTZcfdAzuMzFwiRr3V
QtiZJeHoebb0SF+JgVpufOqxy6wVufMSsM/qfQyFFJpk41fzPjrDTlIh6ZoNuHmSDJVnH6RIoxY4
FlssJR+B5wi/YMwOtbpjcHXmzVywjQkgKLrn0CKb+HDQCDh9suiMUCPMjiXssU5SnVx4Y1kncXUR
0VRPvE7IhvDPGse5tPPYysUZlIiCMAyXaz7a1Nk6K2vMTIXBS2cAiOq8GJ9iEwoFJ+2apQfJEQhJ
P7PVzYCzJbu0XB1uUPu5/Mej2yEAB3SKl0hG2Ih4s4HBPdjPEPFBsTlybDHd81PUFARJoCMahm4E
2zMo0+juIqLjX4S8evOMrDz2hgeawEnkE1ntScwTztYvlpzTFDooQkPA0tXWB9eLr8SEJyPkFBar
a6dU+YSYmCoWjRRi3jtE0c4xZoETl/I70rq08MFoThFQesNFL8J7/cu1hCubJNgW0Do/1PYe2zcP
/idWFEgbTyyexrFHJXGAXnBdwpsYW1UIgRvGWrmlNpyWbzQUW6twI1FMbwOhyv2xuzoAFQM80lVm
zlMrr/ipNEqwdYhTY5C6McZAg7yU8r5k6scOhKF8rWVpXDR0PXq/aU5EFTj/XWcpURns/QPnnmmc
QjgGJlpqQeYfF6ABhcU4Ft1/G0iAJJs8GI27EU5vNClEpscn2SAFf2qI506pfrUIBcfReb/Y6U1n
iaPhIEr/TlCCnPbXKct6NHwaWsOM7Ifx9iVqnUA6lup5EhDnqfsylLKoK1DzeV+/qbpHyMnjIpeG
bbgAgKP5ZFMDFE60FUgIoedVQ2sCzQqIi07Md7IHAHE3qeOh8BgnEvPNDk97+yI2Stkar5ChPQaV
lEd8vSHPnuiGeN1RvRKO39jn3eFIodDxdS1IfZEAYgi3R/7Nz/u4b8NzoQtnTPcRvPYwRXiGl5hN
JiQC319C7DBmBtBmLnzZGmUpLxtdy3+V96R+hz4Ss2sNGILWeVCcxNMU27OEdC+deDWUjJ6yhHgb
m/eTFFypU1/WKfyD3UqpvXi473K7Pkj4AvMWwvAS7lfiqLFP08FVcM4L+MP/znSjE4pENTpElVZo
IiT3bmPf+BNk/QZc8MwPQBKHJs4w4FckP62bjVGJKLAo3F72dgk63RO8AF7lr77GUj3wEkCB94iN
oQhb/YwvkHZd830/ul5t2Hp0r6kyT203F31dU48AjQVXa/AKXMwMxBFtEID47PKCNLcsAfJVjYYk
6Z/mcD/R3kVTxv5zf+YQaL0Sf2aSenfIHP+CcdsSSk0efHDFjRL+h18nQlVXjiyTlSulyONa7Tv0
1Xx11GMSmKfwoNDU8NrokbwRz04euxuNWvS0OTSdnU7YT4Z1LKau9fE7G3xB3G+hoxqitdamceVT
zUViKXMfBKocwOARDY0nryPb9TLPhz/Lp7MLAtJ9ZH3xS1nFUKYJP+HlDm1oZWk7ZvJBCDojlICP
kwtLoKrQqnsjQ81KP0JF0Qhhu0a7Wgm96Hb1MgU+8T/OzYAV3qcnoXuME94/fMUBCzJrQ5Ag501b
00jVmKGFYjdohpD2mTXSQTf4UiVILldtasSonHkTTTxeLguq6a0XDdtJCg3Xbxg3DBrRPjF7KQZF
UORdmf6WbEQlRPpHotvu0dDb3prt8TeGXCg76VPk66QJCIpwpkbIZNnHiklXYoSt8Qoxfn6tWN1E
nI4TCyUcHx05fR6EoV76TN6c3yET06rvgTEw3gutLne6zzeVaNXUDGQnEs99kxwUifnvtBXPiiWA
yvU80iKkETEHRiPROT6duow6VEGe2L7OriiOCN8tRomObN72T26DglJP+un+zsgAVlooYyMmF4sR
vJFV32CZv8FWOfpHOZPSY9Ptox8Gj1iM9rJFlyd4c02rL0Ydi9PyoB91aYDTN2ZzhvcrLdedC8zW
4FgYPaKmqJBj46rUaI9QyNcWxdMEnEc3vxP+Bz09BTIovtqib9lUJrLpdWdLZZsN8XLLB4513s0m
WtSK+HJzxSY8eREcNVJaAOKPq1egFF/nXXuD+zFZwnR9zBVVblfYb12RYU0cq2pdPR4cvqDlub+t
0LAJWV5QlqQftiYAWh6m6YuvYTlwwNvnH70HA1eQe674eR7/rC7a2FnCTJOlAb71mpNLLl/RGjFt
fiQe2kBO1Ya2Lz70o0eo9Nzsqvn6I2pSsW4bL4bVuRJ3fTI1vjumjF/Mu6mfJtWp3baAalU38Kd/
oLiHa8vadIUrZ4DmSvIOTUeFHk4cHeJDSmYet/6ZZgyvgEvUI0Sm4xXDw8tQSo+VLlClpBSBC/3k
7nt6P4ncWnAfGEYIdcdQ30AK2lfKiivB5VCEc9EWYTeh1dyAarHtNmoi3ll/6fYBxdsXErnBaLnM
UZTgEf9k3fDsYoaFqJ9ZiAUeuWFZ7ZvwjiaS5FXL1h3hMuuhwujEuorWy3D9kUs3Kt+jMNJs/h89
VaHwaq76evzLR2hdUZdWKUkomNk4B66Ev2qt2MgCFQ+CzBke2EFqxreXMW5IcCQSu+t6MaTnPvu8
GfU1/xHMEVMoZi4IRUfkj9J7ytwz0pcdTJy7fL2i7u66Jp5KjqkJljyQ0Ko1zc9TKGR72Fszt2vi
GENwLwzm7Hj/w6Pw7wop4q5Sn3MxNXNUDmCBdHqKBCrPPQIquARLPqTFvaYhex9qCoflJ1goMaGn
fUj+t+WQ5/MtKiV2YXHJoXPbu5tc6T/TCn48bnrsjz3G68SviQwjUqFZ9kdZ/CN0YtMbB3m+9c0+
30poQZOAffBIPD2iderFEglUv6OAfzh9i2qUXUankfH7H0KvqJofWL3TaZXzgOwqkATcB5w9H5HQ
ZFYkqXo1kgLMWMV2QXzLTwTJPVZe4yj2gUKPirgBhbQIyXztAOBQVXC/gcA27AfT4XwOWYPrSlti
0gyULsqlVyctFafZrjAbJ3HfQC5D1GQECJtDPx3nlovsljwISuUP1Yt7H1nzTyxTT86jQr5XIwJx
rEUtVTGFRYKSw8FOmFmpWW8g2FV2KwFtCUrGM/Riq4mkAWQH96D+nYx/J41pjvaydHYYblkODBZz
p4jtlqAdAEcfoZqnmNorPTiAOkbseH81YMi91iZ7lFe0o7+KGhGbUXe4wxrHUyi9fwMiaVp1hQwd
e3lzroPUJGYdY2GONVDqBjOm5g1ISvU7d7SIc7INMQ++Wb0yh5SO5fS+6oQ9PiwpHkyA8PHfpsZg
KEk5rYqb4LT3wVlbbDKRd1lWExzkyNHpfnKZqmBFKVnQelLO65nbT3n98s9PkcKDdAJmGqFNnopD
D3MvguCspegv4M/QFCnmoInBwfiUjxCipSODzLDdkytKLp87fWg4x1bVpHxELtBXs2lEm85aaQ/9
a/nY6VPBQRwDjg1b7+9zWUpJVonQni/LB/o68epzWL4CnGe+Tw+mKlsGBQjbykUVlx6OlZ5hP3qN
KCA2aGrtIOYjV5c6Gly2LsLvIDoGDNOBHov7QbX3DICbOlVSww1CXyT2rV0sENC8FDbPav9x8f+U
emLM8OxQs3CmsjxU/7c336R/gDkAnuiIdLFfQpDVJPxniLzVu1fruPMaxwq7D0pFM7iG/AdSbIN9
vy1byl7QVPavuTGlQmUIU6se00eSR4t58KtUvkGvGZVrN/4Jj2uvO3nszWhWDt8WXnPjRM9IuYCU
4DIgAsU4g09wv/YKfKuP6fNJ94pWIXnvyhIdvwncPkp7FRcu2/Ulr3Krb2aP0cMfh0JJDAD5695c
OccoSKqu7Kmrec7Z+qc8tJaG/YufpAfN0WzxHvLmEaKNJz8xeDhkmims+FiYiQwTmx+jAsfDxqXE
eBZ332KW5mpgba7591qtEu3CCti2e4vGA7XPE54+PvLroflpELEMcoNfWN3uFr8xxpajb8irhw0w
9EFjsjrWSWwRIcqCkaGiAjpr1CWORjAkJuRpQ565AVcFkpzUlP54JKOom4M3PhpctDBTeVTbzPQ5
Xl9GbkGTHMB7x3Rvflc9NdbmWLyM5L50DYWvikGsFmxVdBD4BXm1peltkq43a6vf5jjVyNea7S7G
BR/rhDtCz6ju9nWWuoP0NKWFjebmzgOxQ9/JsPrsv6FuqK81YIcQtFFzczsOHE5D1v2lCUPhjmm8
DZbcf7DAcYGC4CB4esOOLpBGuhCxxj3tANTzxJ8oLbLzoPamvLg+cht701t27CLdeERLffOZMrcq
+vWqHxDfCkOvRDem1AtIcuHn5LKUy/ufMbxkeOq04yfioIEzrGjXVkKR8HrNClStBTeTVmUgX4YO
vpVAqHgKClf3SftD874IozQeGtJUdqIwbg9N8F7bSGJ99N/o3eJdqyB6rJYUUJN15EDTynnLjPcR
YnJrgpPJ/s8+/pXj64RZATGJ3mdcwHMeIU8s+MWCB/skWlWAqmxR5iIsVxXKYxvNrn1kZSkJLkXu
kIDuzh97GRubZ1irvB6hRuT0lPzR5JesUooXmzP+zSmK07kVaytL3dZWKhSetIiDF+oqoVwoNfjd
WE6OE5RX5mlGspLezUCAy5m7gpaykh4aDoJFFoYq4dKaunjphFQe7ZxAN3GMwlBEpsiEDWgN7X6S
diN4+jD1HCURfcySo83dvzzb1MOrohneZyMt5SPENDvpYrbyuU8hCRxY5hnUlw2mqHc4p5MSn+Ms
ErH18jZBDc6AoirlMqO1E3dV61ZlV6MttWqAhFOBlLMiN/VUECALVb5EC6ciaYyuORZhoPg+8AB3
bFUSbojm7pUNsc081dg3oVCL3tGHI3DNcch2ob5WG/bnKJbEOHeYxobT4jM7e/l6tzLd87LXT+YT
BX4mCBcQ1f4rFDT3tL4pWpAQQaR7TvDqXwDJxf/MNhQvdveFnqwbZ1kvZ5ap+4OXk4+BFI1Mbv8j
FobWct0pNpXd6J+X9p566RdRkHF6WTdvjYIqvVIxvPKm2iixpG0NysizMxS2bhrq8T7HWdiYwlWF
RHITSJxXkNn7hmWUVEOyjO6xGH24i9YjBS+H5GeVUrL/oPlgP9Aja8xkCtwAqPTxMEFga+Zc4hj4
RaeR5pIqzYQZsFA21xdlgMrv7zSwAyRFr5VRRJs0WpsLRrBwF5fCXH5VKAVFg3wMUoeqd6NmTUN3
7B7lVAahjCE4nQDgqZgM097pupnoAccXpE7W1VkSklmbIL5fqYVbf3trUlrTkk6UKIEN/GrVDrBC
riBRAByMzq8kSerFTBoj7ADhdo5skDceoP5pQGmlvlepsILp93VmLdnuHDZzKV0K3T9aSaoskw5/
983nkac7rTaArin2qzs/cLEnSKg4YGhd/6Mj9ykbBgoPZDhG5x+Vt6zwxkcKauXLrE++BU6hGLaY
mquHeD/HZ/faB+1DXXeWV5sv97ik4IPzCfdunZ2FbYn3vxlAw+AJUIW4lruE5aErM5iBTtBdBkb5
+Ef/1WyzlZIb/W+oYsWVQ9PQ6fIjd6rb/ftJiHak5d8mj0AWPQQjJd46OB0WGpyMNKYDrQLtei/Y
yOWMprdGlp0zQRBejYoNheY2HimTckasimHh8ki2OeH02YMBJR2GuQVYXtynlRHP13w0jDiTjmSK
4PL0NQw6/1Sg+xiJ/xuq4wTeFf4A5+Evn0MPEuM8Ipc+OiiWUZABoJAvzBIbFsscvtxbLBqHcmrP
ro5qySXkxDZSR38Qez1GoBzvi5PVBqJFL0G4dmBbgcCIuqTkbKLZT05V5ruC5wv0heDm/jHjxL5d
u+/8lm3PCgrrfnQFCpohytoW8DB1bLB2L9BzUCl0xRTEQI3AWGkUQPgVF/G3C8G/bgcxeFeZ78uP
V9wwwYYWB6HHtSqtj2pqISgE4mvIOkwGtYW9kigz9ujEp4OxLUbJe20MS0/ra2acyxFtEFnNOX+c
olOgFdR7YG3NnMxENohKXz6/Gr9KWt64yrhxTtyYkAKPwy/AlZ1rSVl3opGkYUEGGnuXM/r6JebG
e1pXbF87vOh/LCqX8EJ7KCE69kLZa4bVGUm8t3vSebPKIycVYeVFx5Vhe4EWnYxMWUYPtBhIVd16
/J0LrcqEIvFi21JeLJZ6ZTNf8u/ZZebCJ2AQn22rDtrD3LkVeI3/nq2++hU0cO2VJTKmbbJic0/I
EVx3Hg59b7AGV04D0DmhnmATn1hKGuFMqVXsIokJoDh2ws2gFK0kyarc1fUSLCklSLOdMdVafANA
eXCm0bAxlgg/lESuXphj6GDSaRMGqSgzax2nrTcieWtx7sLnrqyyBXFp0ta0mcRi8LIFzCh/IPUx
ogG/6UrRQSYMBZIm9NetvNnvjcZvy+7OVwwQ7d1fE8CFdc9AOzo4bRLmU+F+93hTTIoZNgjHu3Go
+ZZBgXBGsbL/66toUItLJaZTY5e1BPQeENjGVA2AuZTHtxHSCmjWUSppha8EYLdyzONXUQ8htgG6
3yCqeDNg059TFzMV51tg1o8DWvQjRmpo2rheTn+/7VJai06RaUA/bE2+fhn2b4TX+OK3PG2I51jF
FxNz6489pupPeHNF44YNz3J9QOM0HSoIIiFeI5AWzVb9ILsHdcHxsTpvFfvkpm6O1tdJO+4y9wLk
uw75m9OuYhANRA2Ar/bL7T7V581+JJv+6vY6cZxnxkbRJpFpLnjQSY/ku+PIeUzhjiCzLF9HQFX2
db4p+T4raoCIYg+CvHoD3JtfsCbzy4qCMsdylJsIdR2v3V3G/Z/nxs52YIHS+Dg2IF4cBHOP+Zd+
rCFSIAZRs7zC80B1xgVS/VDTZ6OmspZ8ciLwWDadXcISRsRBz32rfsxPuWDAA6C29laZ383Ko8be
6oRyv3/M74LVlzEzUWy8jZbCWZcjPhsh3YaQonXFme6IkYi5svK1Ct7ajHdYJlh+Vv38BbOOqCiS
fdxRfNSErrgsltoUgYJMVMALXt1S+l/21E/oAiZPCWQ3kPhunVQepvkuCe/HTf0nes7au3MTHt2j
9OtHoZlQEupCkMl7WxrL33WI2PH4oLe1SgQyL1gNuasy7OTILveH0sGZE0o1R5z3i1SUKKvQileO
OBRynQvcc68GRN7WhdReUfajYE58Kprb9KS3t0mTTRsZK6lxgt23prRvVqRvxJIBrVt7Uugu25Ub
BaecL60pX6omwTVepzItXwd6l2v2YyE9g2E5hROjTKn9awkeAiyreatLROlmi6YClmo1YPPY7JHI
5YQGEJJ65Nb6tGcKZrsKSuTaYLgoCB3A3YwN8R2p2fL5g3kv7y744bYCCGCkO9fXgbHPjmIMxSwf
ZAjhPN5VVe9vwCy19oAkrkWAYEV66G79/sFzCvEEtW8nGBSh45wzdn9i0yW5QA1nhbTh2ALVfxkf
xp85Arx5fuFYYh43VyVo0W85cw0UwDluhDVoWdaFIeVdmHzHw8C38g8LApC58BRNBI+xZ08vcFOe
5aUalmuwJWc18ol2gb5lIlqOVTlaVYJvrXbrznfa2aN3lD0kA70kNGz0Vb6u59J4ijEsjprJMGjK
7PnA5deyShxN3oNAT0Rm4F+y5OJbBRGmaxsE3jUhwlDljact0h2vxMgzM4nxv1TJ4OJEz5xLb8fC
StmHE1Mxf3GuLZNArK5ZNfaVpynJevSLm+3C4mxkD//52saM6Dw1UDjR9ylVRouGRikuTjXl5q4a
whA4a8siqibmdd1W/zn+2ozPs/TJTVSQChIi1EdBbgo0zNbplrpwkI5FH6M6pM723JW3apMnz28t
mE0cunm75/WzWV2A+ZEhXXR5mFebPSDcUJ0aPBXuTMGxx8n8mVCKIDpyfpXXrq0RMBPWavpQARz3
6Wis9JsXlaG7MvzCMa6kdHKev9C5dRqgB3+LDvXpsZJbXl5QtFhOwLaqqDMyJhX2IWBKshAoTl5Z
FbIKdpVymFWe0MrbJlhJZ6uH8w7KO8r6qWbUPxrgDAp01AZZgIvN2ZJxCLjWVPy57Q3Igqgc4Dqm
pA73oywOzgrh93nFdqSl5hCHLD6Nf++ypHmCK+K+Xo7y8TFffVBnVRdHmpTy/2pqBOj7nTii+6Ay
vyeS4OXQs72VdMRFqlOocjPMFmr048vqFFaJXTyq0MhsaPQfnxV0FykgC6Ml60r10Gw48GI43HSv
KOo+xo7kMsu1qa+ymqNx8EK6xJ+QnaKmRJSq7m1ijOwEuVRKKPA523Dhgfb/WvQD+XC7mJ38YfXn
/EhG+zAWYpw3k+JFpAlJXcDwYqQBph2ytqaqa4O4u871bEEsH6mO69kNibbr1oG4FhlYVPJukNzj
xEi/zd3WbPzfMrBebCFNqWwXNZiadJ5SqUPqoErp5asadOdLFnPL1Xb6dXCTCZ0HMsCApiPwx68W
MjB/ln1hDLNlHf46XQw1rHiEZ5oOWWNtc1Um5Ix+st0Cdaxuvm4dzq6C9tFe7YaDnLgW8e/CGkff
zBRcwQ2adgteJMJyepHakjpSIbph346A078HKeBHdH+S9cuV+xJbfqiLtlEBcRsxANjiyNlAoSUX
Awog2eBmRiDlgwZfU0cwhxcsUPyGZONo46HnF5cOw2MhtBEAF1xLahlqPLxxcDV0Y/BZQE5q1YdC
441/9nRBOdc290c7NL3Qvsu4708B34SFZL1/vVL3atFQW18CRugfOciXcnw4ldWTIy964YTMB/H4
dwXb9kyqeYVPqMtCB+L0uVU0OmoUuUrVdQ8PydMMjDhSTz3J4F5JKNBiGFx0aWnxbHcrIW8KdwT6
aWodxGTOeGFlszodBDH9/4ruTgJHehth1DG9fmaZm/uXbyg8o5skVbnkLBUDhBfpawcKL2reuLRt
KWZteZlLWkOccuLHt1rTjnYw1xUoVqz+x1DOP5dYgkdYgHx0m+v03DgLfYr9PtLoWQZh0fOJB9dx
jGsJJUqTpPDeLgUcomMoIrYi/et+MYyhJBhOM+mHH67tHNSJpKxonfrkRfAW08xsTnQNlt57Wl46
g4XiU3MJReEIJuYbeLbvjGw5TzVQPpqWCU2p6uVj3vfWWg3OTzdxqnZYVZJ/DoAfpewqQ+0UeMGb
4ZtzP5FvZya+sGVXVAH7t4d1BHH/QOZXaNw6dvH0erGo7EPStKTkU4bY31BlYG4zngx7IOqZUXP0
4YfYEXLPPOENDUaXIfP1LyCPghh2ZTzhFr54WJyMOfsk1MoiwIxIebU1hJaVSe8z6rgjLVxz/tAO
i0Z/CFODSDhRT5NYKHqt+B4o7vgjpsRaCeDqFCBHVuot8o25JXuQjvwON4nnC3wduj4um3+a3oAI
J9sBYVHBWsWGtlQYF0TMpDkDc2ucT2apoM2A87P0QOIl03jK8i6Jj33cSLmp0XxxlJlQmjom8EI7
269tClDB/fwkM2KveYQF68hYFdATtJspgx5RGHb8WPSUA83JRc7r34uNGJUinAZT7Tr09AeTWmsS
be9kaU8zEpJ9xpv9+8iJxpxB60sGU2SXFk302V/yOphdpEkTUHNSqzaP9Go8jmcVTX9VNSknKPOh
5/nHOIi51BMurpQ3D5HkXNNTUJKyRQn3DCZ01Hj5HQ+KwWweG3gR9OOgYcYGOfolbnHu4vl+/eLN
4tsDyzdNGoixCNNOLmiEz2ibv9phM/op0WycUoEb33+jGeJTYVtRnmWi04sN6mL3r3MHpwRbQ+zz
qgTgU1tuEDMP6KsJb2ZmIOp9SMwBnD8cUqn/Z95USCfuOtxxxr+Dm07vOM+YuiMI5Y6WIYfrt16X
7sqmzkoLcP6WJbHRcfTWV1KI0qDI7hyidrNfuuoDNUCTlatKXCqQPUdQ0OLBHhfViEsGmFDG7bHq
fbs0BoD9DkYNJoe05MTzfRU7rYAAO/LxtkYhxTdjhGmCcGNPIm/dsNshaVD364J9VpGVJHN3Rvy7
hdNMUcclWXF1KF7SekSsLgVZwKFw45dA/NMhvT0WFurCPP7Coo0AIlO7wKDAU2lXp0dFj8BGucXe
mvF1tVjnDtntdmf9CD3EdE+GpkyDriksXgW9A858aVP3qB4ilyrPymaVWaJCX9GoYIeUug7UPNnt
jpbXxsiBlN5L1VrrAvvGt0AiMhvEN9xjHXMXf6joke5VSRrHa7EFz5fMWpzU+CyaPmPkAtl3sMG0
FNIvFYpbl5rwwYc7GqxUZQhyMEaJEkzROyd1ovF6JlFLFfTegJrYKzcsQErM4zVope2+7R0CdN8r
Pt5O3Hrs2RjZqkkCHb40EKvOq+zTJhC1J9txSN9I5gnz/EqMLQtwjNTmEMi8IHgFziOE2i5ggXBp
/blpdMxL/dHmWuRGtzU8swsOUeB8sX6WLKN21SkqeEISqSLDgl8S20i/AARAXAB9tlV57o9sEJ1x
/dwYGsWJYSv6//uEKbBub8Dj7gNwf/5cNX6uHgiAntXsFbOkjar7YwAKx1wXqXzrygLaO3YdC8/l
3sMeLxz0pda3OQjzVTEyJjQnX6LIidmWd0GIyBXz4X5GHNioO182PfAgeKd4FRVCJUqNNt0z65vk
4LNE5KUsIEgq/0XbYC84wqibEtwAvjoVMIQor7HKIQNvhwzB/85iOlogAW3IYAXr7vmBS9y23RXT
R20cjRdHf7duI2OUTKmdsWx/QXvzOIAjB860mBDxc0PRsGM5ZleT+jZSXry8WVSAzRmdshKCvWBA
5ljBH++svrC/b27QUSL/HPMUeoo8WDMJjJFvS0d0Qm1It4bnsAbXSqOMPYmjWBhT7EIuEu1ylmU7
vFacXz+NmRwDgY1eKcEafzDs22HkkqUlS7jaPmt8BQIEjIf1SPEq1LSNmSltk0yGvJb5dotFClp/
u6hZH+E0Y7nD3Sq2x3kG5smYAfMJ7zzcWXDCVb909SBSJ2YcdGoxJnU4LSyTrKuu3rvH/7/DBNCk
nw9b5UXZ9Jmywb8CZhGT9aE82xyZbsAsxEPlyh6FuckdwOiEpIhn/lJTeXy/4mAa4PuQbDRJD+3F
FRVEeE+nM6TMonu9r3pSraGw6uWBmqWe1CtHkZdqnPTmAb3btNL7GmMZPHQN2qmXjobD64nYzcr1
9UxakWa4qg8l2aIArFLv39IivdQ6TeQ9cUcmSuE4PJkgGSbFLK+vZPFrxLFh7h0lYJPabFQIPzlx
1a0TdOloI8hSi/PCnSaXRspQi0yMW1oBHVLEkLz9sdyNaJ9KpqHRG7O/QmQStY+ri5jhxylyMXFZ
csiyHMn3FtHUokh8K4iE9aqMGNRFhQbOhVr3wqs6pJSznfTx3VVoA5sYB4GK/sSAF4Gddk4cBcSf
huvi7M8I4gmFydvxD+5gdhqdJQ/g/t/c2iAr3QAUYnqGOYr8lTAl438b6wzwjFpezbCkTC2O08UZ
TfGxss6l99OtLCtuUs4EY+wGf0StFP9dQj1WsxKLOPSM+N7kFE3KoyxKkq05TVJ+rDMiuATsmyX7
1HapYSjqVRp7ISQxeLZcxdBrv+pYNPu2KuXmIftYimvFBkxnx/KUjcyx8jNj5TcBSqemLBGkwlJg
L/TuM0YvdniTigyO++rKOPQdlzJGUrd9Kei4Dzr5to4ibS4TnSTvLCw9bvjEyhSrXHtZfBy5yQQO
9h3LMc++A5ur0IVJsa4noko2xSYT7zPVkFa6XoIu/63b3XnC0mxfl++3Ho301LG14cGlIsVQ2wn7
6wNd1pOGxSIR6DW1WactR5a67CfN4Ta8sSzsuMqUdHew0Z1FuQLd3aCS2Xrr9DJ7qqgxAKXWwhQy
4xG3XnPOa9QKh9+CUQORxMVlK8u3tceaApPdvC2UTs9Y2Jfsbndas1oot6LXqJD5E0om6LmeAxV7
Jx73nzGhGiRljzByGhwr/Jf+yJTW0HiaWNdF6C3JPHyRmVWW0QIYH0K+acO71vLoayhtyF8oW9io
Jldl321ArY2EhCj2A7KcR5V8ztx5UTfo0mn9TDPX5UHK/VWw3I20dP4Wc5dEdZ3gAekobbh3g/Mn
KtLx4nWFN+FIqtLpncs6a4gxE6N/U65mTG68ATQZHPuIfqd2j3+QB95NikSlPFTKK7f+PfbycLMA
pKQJlkDtTjdArH1jBxRG2hdlZdw0eeECbtrKp9+Dq46e+7ky5qbnwrAl+FcPjBzBtFGfj6i8e4M0
RwNwc9IsrvEIvJEVtg6zilyQETNLxxjgebGkZ4FPSbAcKbTj0EmF8FHJaVytBTJDe53Hue8rDUPo
1ugeY0bPgzIn2+nF/HCL+FzfGW927C4vV/YJ1djJaBWhiXkUqULivS4lEwhFGqXklR8VHC8uMT3w
+wgcgo2+mp53F06WkEg88z9wsfBL6d32KF8lYgyeb14r/33uKujeWmzWB0ZiCI7pwSCWL0U8ofdm
9ZVc4T/ptdRYfnbDU3r9f0FO56fwY6AKyEbv2/LcUPT2fyhEdMp0KODM1fvtwB87tkEXKNR4MgUj
szL9b53Ey4Cya8GZ9jIsys+ooR0CQ5ksI6ZdN+n0jYtH9gcvxE+XdW5LaXfTQ8FAGIrEZ2FCYyhx
skRYSSjZGoHG6yIpjo7s70DawyZk8ITQIaj0GcKPpTfWIfmWmd8IeydbS0R8hg4CchiiVZHLIiXP
rcdqSMvvy4g4q8WdggiYKU6tH20RDiF5Vhg9N9UVaSFP0lhlb/Nz/KwU3bbrRBbabbjfccGkfFLj
dZJIa2b18ckqSm+rsaG4zmQfmEtZUYrHPgD0HST+rHF96uvhNGilVLW+b2FRXL73ndhY3UbXJhE+
FTJf/y8ZP5SvIWyrDXR3Ky8SkmvWOqZElyd1yHGi9A1zGUAc9HlnQgSynqACppp6zcM55pMRzy1Y
W6Jrs13U8V0F8ywjZSGZjkUKHpsoD7SbSpjBXBiwgesxaia0W6HjoMZo/s+dzm7dbmehozd7hBqx
ukBki3Fn5k4pZjHKljNbGicPJr+rg3zBTKuBrY1uu0LfvGYPrMb9MUAuVG0tw7Tri7VPTM15AFW5
udWLMl2rG44ZUyuCoUTxLs5HoMkx7PnCf0N8feNxUKuzxGW42vKKAmOQANpSs/7byGNlqrVBXeyV
5yImXeDCcyU4qpiAWLHzglynJmhENQ/lewK4TVh8DwhA36cKjO465xd1b+iaIVb7SFrR6HYI31Ul
40pemYfEe9NO5TXNi6/sBvj4gDa1Spz691dF78yTaoTULPV4NLLQ61TyvatroJEM/BcSCFK1uX1S
2+xmCbrytFHp4HZ8IvEAPGB+cwdf5gyNIpCQss2KW3hCsHMKZ9y9uacyyYCeNoZ+j+i7MJkP3DwO
mPCSAvKhxYSWoAspk/SK13JZcVQQwzqMTZYT2GrnATj8/1dqRxICo8wkuQNHl1gvIOkWlETit22B
yX3kaJhl6Sfx2Hda213ngW+8447qOHmh+qUdFoQFJ7vXb/5P7swdgaLW2CS1qUzhFI2fJTZRlmpJ
UVvp0Mofr+v2CA2rEa4F2M05BAf8eIKazG2wJvFv3okGcYr9IspS9AFPYNBgi/vbPmlY89vO2asm
+SUg+V7oQUInSoTLQtEL3DUHi609rUHUMCAoA571R5EhRo+XGIsNqD/F3UAtZZnje2HmPZwUzvS1
F+ksHCnrwt8F+hLvjqLJg3OjXErDrB7RxGMF6SNwMONkCl+k0D9pmDpo8DS2hjWD2Jw0rCqGom6Z
GXI+AgO95Xyjq2M/t3Oh2B/Yys3bVOJSCOkwXb3qKgTS9C9VjWUyCIpC38W87T0ruxo2fsTyaeXY
CcgNfY2rOx3lU/CzQd7omUmILTaohvXdozufcpQkoRaMuPyDuZGy8ywiC/zORKDzUvwoMR6Ls+Oo
FZT1b12z0Pv+E5xDHbyDUNPL7cPaTpwYsvYpyhnpUUgXtxoFRrOTSGGuy9aV3n2hM1fQqaeNMc+U
svOjuQ1Qdd41Cv0Z0DYjzDG6HG/LBV/+CJXQomPBq5VB6bIS2cDQbWWUVN/HWcrZYwg+XCLpZL+L
SFlH4MZ/hGWkUwjRqbvQByQ2scIQdWUZ60VSxidsY4NLnMmgBK1Cu1v5hxJCpuGnCpvcX6QSRCIR
w1QMbmbwddUhgK2y8ub8773WfNVwKu2fbsw6tVm0V+9iZomM1eMJw0Dlvp2/JZi/vvNxgrEIYRU8
QAIGBG4Ast3BS52Hw5U79IcorYDX4ZH9oKA/GFT2AUbtuwSedfJ2KsAZHXBhxhiMk4Ayzy0fJkKP
l+SfLYkWAquzf3cdcg15QfilMtafy4Ym6+bRohXTkFoQ1ef8MZhjVc6y4Igw29RRs/vmwMpftIkq
jFuwBZAj9UJL3X/g74XIcKLe4j7Q7ImdRHPDSiHekE2UioKkPWmvjEWLW9GsBstwRUocdKj49Zoj
mGvnF/5WMYrlDYglkGExTVaLxzg9ib9rNjz9p82qetZcBJ0MYQdxD1K4FE3t+iPXdW3q25x4aGXS
JM3iJU4OzIdJ1nKhrMudw1W+o0eSXRCdFRFYoXvtyJ1AIdsYv+ZX9RQwXiofqVIJGXM9aI9BArVu
GHcFrO2Q3+NCAE15h2jjZiVOGslqwvWcucxUewJw2lCu++aKG829UsWAl6gFPevTda3akqIhco0N
tGT2hwGbc9VOVgssetfw8mz93HWl1rgHNrE1OSIm9Lhlo7/0xIP9hGDGlkP+n0sp8cIEqFQwB6un
d7sZKl9L4buqwMJSWNEPjxc41uzQ8O0HGxX2i2pnLC4sXNV8IzwUHCyp8p0VEVEv7IFyREsKoeyl
04uTaEeQUehXW8rutUXdi6+gZ/qPP0bICKkEeA6DhO8uLmXuhMEeb3SOgf65lK7gzQIGkk6WJYe8
eUChmKrFm3hkcqCcL7VZ/OkW4ABKM0rpHAwR1QmR2Kw2hSpZPyrfa3Lcg8oDTx3LntPX8lLWPV3B
3JcHHtlsWkDMEx8asPe4Qz5ZKGg7G7OHLVVAdVKtDrtOcv1JHqPUx7A7fN2fWbkfn8ZJdMNz6y+H
9pgTXPa/+PgDwyd2nJnVqgpStxKfEgjw1Pbau+h84lHiLhVY6+iM3xeLqwN01CPF2PQRjWmeuejx
kMbYXEGXKrRCubdl0agoA166sjvClYTM6TRC+o3ki9ALr62AGHxqy2aaaBLGUKNlZ9WliUWSJszR
tnqm/+KE+H626DMOvfvWYT+dyTCZ7a34nzgPxZaLE5mHvS8+KGghd8cnWgIB5uSopwOObrsLpPCn
wv8CPlyOxOaroAPUbelj54gcscDDdIL5VpYWjTaIGG4VSIva5P1S8JmbgjtZKifwWmpoXWOgtWxx
lz2WJ43UZv3GZleNFa4BbEoFInCUcvuDE4WpNPkvkXJZoq4/i8gLfaXZbkC/MXi4xbO3aci4n2CJ
HPaYCX0UjUoKsqxFJa5PHjZkv2SbJn0HjaiiRfK0x8Q6CTQxGljR9ZgFQUZcCZOIQ6cr773lFYgm
N8OlvLmF/vcRMvU6O2t6Y2flJDZV/V3RX0p1UrRkBNoxjsNErep+bTcpsZ2nSKgqGOOlMxIQ7K2c
02inO3LKHg9ANFe1QOit62g+1RHqlggPz0xFcfnAbVHV2914pKRXy6hauprXKF1xB38mA0lSCwpn
m7uxFlAQX58ddHAOuK6p/DyNmnySzXJIqnCUnOUE08QrkaNa8gg8X5X/0xAN8pJasVeTa9KcsKc8
N/F/ZxgUAJn/QZ6mTB9pM65zSmwFsKOyI4RLueeXETbraMUYZmXuPHXnfSMO8u4bstt4ZXEplVSN
+Q5pC4/zLKBxGpe/OhHwHRU+RnXy06onaQ4/9CRZ6tbxKbGZx0IMEOAioVXEWzZNc/6fiKftsmIA
nYXK8mA7VIqjkR+jqfYeGmdxcx5cKlTjeosCyH94lTx/MaT5pRoPj4RhF/9WEjAwjbdSX6TbXQpf
oHskOyL0kbQ8hSBTt9ZJW+GSMmUVr3EQP2xmQxSfz5wT0KdL12mf0yvTF5aE6VcRjoZ2QMbKUDJZ
lztyPtBTrmxjhE5KnMjN+l0vx/tUDTMGAREtoJbRIY1fzttr1kHmoO8J/7JTyNyew1RWAqnYhc67
l0aESgYHh/t7VYQVf14Sx2nSh2Wpm7Vj3h+SN/66pe5NMX/WH5DTWNpY75U2UIxLhA5XEeC0mhWr
yJcVH9YYQJBFMIw7wQT4ioBZ6DnQq1QVMAVVSuhsfwMq4/J2NJevtgKpP+t+1lFCt6YDl4LmxIBH
m0syF/5tY6E6Vtz/GDJXQsLE87tRJvE6AfUBAbRgWpVaLCkgsEkBAGsBO4tuBCYWZ1QV2zYrBQz6
mhzalKpOeHGBKF2Z2aL809yFX+PLTOhbVHJZiGYknQ985R1gs8Xk3zenYCCOxTdmp4Q6JLDoWUMw
/ECl/4eZNUUFC427+ol4hshPoUOha4DE5H9/ETjRALX9QqVaYkIjmH4AuwftJtvQ6kT7KafTtzKz
Ewy4aGd1XsmoM+5MGiexQkMG9IBIHqm3v5jXMR4WTl5qgJKsk4YBhMIAwcqUBrA/x02uxP+GH7AA
R0MHSwL+Pt6s/28SEJ2BhEhPdJy7D1Uw4T1bINJMqylmZxCWPey9H3pNAHfumpLyUrlddwluMvUM
NIZn/i8N5x4r3QIBnN88yP+v+1RtVIVVnWfi28tgYWyzUmdOPT4/5x2BcgkwV1ENfwBqiOQldjEG
5ccmXy5JNRnYDv8Voz11q6zCj0X6FQEaRuNMcTsHZBTu9E3JZ0MaPoujQbUCzSa01LDVUKL1UrJP
aQa6vyoBF7V60JW/XF7CkU04JKtG6qZlt/c7XXGfMHsV2gPSsB59QjS2nu2ezfxC1e4iOCZeGOEw
qbJbVo35AwnaaHn3zh9F6YBrYrwNApBREdmPxn5ib5q4i/jQQSmhMpbhVaKLflTGJFmAlG8YAaxz
Z+1gUvRcktO6nBV3HclOWiY2yO8RNWjzFwhP9WNWCxK35EwCg26XcHIn6vjRy61yn1YCGMeveHHK
zOxYUjXK2dRAfxYgLFtYPydEtu9hijTQIxXnNHZNl8ozjiLw33F5v/mCt9wOpyryePslrr5J0JRe
h+q66YXDjmBPUsDA25HXhXTiRLwcHGGUGRb1Ex/AXhAYVG5CMljZWiwutlCuyRuZtap/oRBEBMeQ
HnndDvP0sa8oVOF/m2IL8BFGZakCWwF5ciMvxbb+8FOS9uyS7cs758NqvtR8FKhqQlx8x7UbgXLl
weV3215GeyE+FfsGwk2QmbR+bENNFwrs72zg4MweuRCYhWlSKIy6gjvZN3yLIoYMMq6WeXdHvbMT
UbbacXbknO2u8QyUFOm5v7+c64o3/D1pAHrToUTbEtB2YVBLQcN9oVl85labN3/msWQEeg1kDBod
rx3NaeM9pBTv3XGo9OW858yZcFGWRFo/BPoJF6aiITHzNzcdANX+gvmmfZJIutOC+Oo95SmacOgS
Z1D3spkJbRFGrBbSqYHDF9x/cL1qmtl/AHI6XbDYq+n3Dv7N4mm8AvJ9Db5QFD1Q9exG4nD8Q/J5
c5Z+OMFB4IYWvGW7jX8S1cIgu2/7BT6Z+deR0XFv1AwgSZO1tkfdeT+GHxv8AbmlNOFwNBnce+Kc
Z0MTmy85bPMz/QRlaa/HtWM8b+61TmiM1+88gGA5i/HnVaLKHdUXyyYABvlcexQ8tQnsg7JJ1bA1
GG5reNPSoWNmcdb2+X9fAtYyyje37pNXotl1eFw86uBUd9+sTT+OZYrq0EOAobE8RduMeA9KkMZc
k66PEtHx/biyOBB0BBOOIK3Y7mS5gGlOD0Qnbn+Lk9O8Ptadm3/JaZMN5ka3ZVgQMZHf8RnqOOFX
y5TP4l0M48vf97qotXy+RqdS5bvJMm6ri2x1MINHZZXrVziZ/pPBYHOJd29pORFEy6rohR6A8A4o
dHvi8WhMPD07jB/R6D1PQcwtH5fkwtAOReeB5zuyKriucXATbr62mTO0xI3tg3n33rp7Oof9v7Q3
IL6975P3rpiKkY+KDbfj9bj7VbqE9KNfKj0tnvissEbfi+L1ZFSeXrMpVZxfrE54ZtkoxOwZRcF2
9Tpo9pxrIYnQzNrumqGuVJhNErtJtBtlyXJ2rd5Km0fQkUzFPqDN7J+bjlsz7oxMJ9O5LQholiDq
ohSGSraVX6VdHIk8/WtcWC1JyUyQEw85JLd5zvQOdkFtdjO5vlbvrNmw3d8SP6kWVFlgbOOhPaDN
SUA/rJhlj11z2dM0XarpcadOk+AmTObjDrjIpnIdziSmb7YzVGaDFe3xl28B3iVHj+SLPl+nqBru
ARadpS4Bh3TGhv8bv1QwWADDRNdccvITdtWfjXyL1WS3ascvgBbzCIIYiYC1e36gQsk6fFDQybAe
s3sOB2SsiHGCmn457Z0QL3ZtAa+gNa2Hl5cldg/rtcKOe3s6wfC1ANCt+kC/RcbrvQ5AIEZEUyOg
9XusHTq2afUSul/jJJKNbiOEqyZwbisC2Oph6uXRBPLLb7CaYsX4nTzOiwYab+bV15x9zghIaSI8
DCi1bhQk+tLwTq4Myu1EweRLuU8aHaHnx3t3iD9lwGMrSSjG5pgyMdEfCrsFDOUaNZWIU/NC22AP
aHkO+Zk/H462U3JvOPDK6dRv2sJ3No9YTz8DhGhVHfeFJbPlC5wb/WNqoCXFs/HS68Icfx1y84bE
tNWGD9R5qUwbQmFq461L3y+VFGt6alIwRyN3NlDeiNhxmSnA4UOcA+zXygyRrr7oK0iV8PWxSeT2
lGv1xK+FnkcES0GdcO6EQMWqpVIav86FwDErJp2FhaqyBObVzJJILj0hUE0+WdUzkR4ZqZDkyyA/
rLJIlyOsEfjUA93AIPOyLMUnUQOFKL9DtqaBENEBigOgmb6GmrLwSXe5byk6cundrSGpoXfLX3f1
/uygh2jrGAuLZw40GXjujPv0NY3o3MIKaCd4Uocf6WNYYzDRxjNmBM1X6ejoOTz1YqiNzOAT0gMW
YfhxuSarM/yKh+0IMFpDbdEt9nkRuD2wcZEiXAbSsVzWpSKpISDD01MS/ArLMOyT0xvIJJZQvqxw
snAtgZq4wnBooqQ46ibX0Ld0YMKgw3puZBABYlQwHNHAoirVm+kOR6puc9BitoxeyPTKC/dpv8E/
kh6JSUxIeBA5X90T4QYnqadLgm71q0lY9oGVjgBEf704Mx7A2AkAosX7Ljskt7+40qnBfrJST9f4
aoVGyqKMfBvORdTULLyJMM5m63mA9yYH7km41gPADp6Adj04Yy8UKNbkX1e5NXWAUBCjUnBQujpd
LVTSth0Lj0AmVWujpJcfIbvgD6WVIATU6sN8ZDbLRAMRvkeBFqqZkptMOl6fsATasy8FH0EPdKCZ
6fa4TN2ZhDqUGp99zqmuwXb9nKWJeWUT1dFY1Yd4SdanfAlBaN0hW+o1fpRm3I70KMvHhFd0Oqa3
oxAzg8+YGDuU3Dj98a+p/W7C6qP68DWXEpWQhLXX3qW7e+kv3vDePCSytPgXhEFkDWaGetNkvqT7
xrNMCqj3EdHkEQjY7WXMEBlz6XIYqe3LDYOgw/sEeAX6t5UmxFyZ9MhTtDv1UzvxQuRrmJGS+euf
H+57jZ/lw8UK0FnTQ8BCtqBHRjlux4uBIsF+0rw2Vin2VYsc+Cp4+5bYwuUsZK+fbjw3gB9Yl2EW
eG2Lv+n81lXTlJV1hp0/D9LdkB+GlvQaUAOfTWVToApobUbByRECpuCkUspgL/by1rzbOchhDn13
LZ7+eDljjx2aK0LpG5D5us5SqlbrXtCNIJpI4LdZ4Xl9gnVkYPRVzn2ZQLNqqRAdihIn7Ft3+6BX
WzF3P0rijtwkOkznq9FMnScJMu+S+0ABY9+937oSgnPt4nbz5OQEvXHB6TxzhBDAnmr+Fm9uQLPE
UaCobaWoJVMaGmOqkxrph5Im0deJOPR0ZL2L1c1v9eTHgiY9u4aiPjipw2m4nasBXy2kJsHm54ft
qtEutvgWpWtmww+iGSwYLbrjJONbUuMT3Oe7+gwrev6iEXi9bhrgImXn3M0KMYXDAkPdqUs5VkIy
LMnW5GQRFeULeKSIEUKysXd3JyLzdQtbRn9Oaz9mGY09NSRWa9nmgu2AYOfWyw0y4ZpctzxWQCsK
6cMtL+84rcXthsDR6Qhx+W4YEj1kNIXFIzoI0MJhhukqw7+oyIYRJ+LsyX8a32S6rSPnR4whFhEv
FF9BWOW2ZgVAjKf8BiQRQnpnvqTzWQTH+Gd9fqvKFC/QYKFf0mUNPOPGafT71DIlDNeMViIkw+kc
/l4SSVBrUggkraS4Ses+2FcGGZG1+1vPGVjdng0m2aO9NA+LLKd5ngNxqDAHmVufuAVPmt4VeaH9
8oM368GD/rzRmnSMC3M++PFDcXHzPStJ2UDLpzvwNkGBITuVqZzpLG5Ku2vbQMqRRAU0RtJUMDqb
KE2mepbF0m0Z4vx+dFoks3zSAG8dYU/YnK+yfBE6kH7/aWPGhjcDV8/gOdZ7E+DGkALvzk0MdasG
qvHuBsTo5jvK/B0KxWV1bHabGOuc6Tr12TUPPzwSGXyEe2wjR6XMHsLUSSpgvRmWOfd3p9FGzCFV
DjSvdpwXijewmdSHgSdSMbxNlrs5iGcop5j9vFMZkMNDgvrcJhyfgbTTgL11TPuoEL319eukKYGl
T9jpF6QgyAq/CWUBnJtkawf2IF1cgQEno7s3/wRTA7PyA3T4UvLOqFgWt+wVOInac9+qjugCLqAE
sz3RusuB1dm2w6yh0blhFIgTLdJjahkbTvEZ2hCRFbBJGEEbgDze0dSP21mxu6g4NnTgAf4nLg2k
or8+BamZFLVmyL0XfWMw0ym//2Q4kNCk64AH/oHyI5dZN6gRaAQf8LtJoGDFctkThhfNB9ZukUpk
u6WLeEftHmiDMv3Bzov0KICx8G4d4lqiMkLJCtjPCxx0D1gEvR6qbCwe25VA2otJKhz8aFc/Tw8j
blQEf1CKBzQj++jJEgDG+RH1K0BjkpBGKILuYsW9l9SZsnD9iGd/9WZUSSCDRqBxv2qaizvaCJgN
b2C0fEtmzLP7BFnd5HR6MyXEMcOTnvZUgLBlLhd3IgS//pw+LaRauhE84GzjtT+5B8Ssf13/7m/W
JyJSS0pk+iqFSVOOlnI+8iYcyjX+E22kyUaQ1WE4HnLFY6TUdED/bXcqs8ybGFitR+wux02UaQUF
rJ2KAi+OepJ+XDpa/EBpF4hOqF6CszIw0C1RdYhM7UoDbO6mkvPmmLQyDKrkhY1sXIIRd/yOWqAT
ujGoExDxyu0WnJqsgbJsLDy7H00fZj4uVjSrnVSxJvjBcVLz+FfVcnchGhc4B/jQmZ7jMcfb9tU3
Znwao9Dleryst+7AIKQjIV2WtmxHmxFfHhPHRIfIuekF3fixd3X/nQHlipaQ00hirxK/chz9WGKR
KVVQAUCkK64iU+qUZ97ilY9Zo6lUHV7zKOIcLrD18zCeUKos4GPlhkkm2JprTcwb5pfYPZ43erCw
+WOf6oee/Y4uAdK0tFGYEQSTlC2qDGgzi9DCRLf6ktSSQUn1olcanHqIUtZ+aMhO0ysyEb7qVJIS
qczLTdgmZV40ooygvob1YWpMhoZpWWOyX9jmuf7dyKXgEtv4tLzmTuxJ+KZHWDpHx26LZgYpaWYB
AiAxNRSFo3Y48wQuAMl1Q3/kGVX95XZGetRfAmYZYAeF5n0cjUAYb1s3hk9hNeTCCWNAYfZYNu/L
bXFMA9zqJkMS58CE9aQRCjH8v8hSVAuYn7otUU8NSSmTMtk9sWs5g78Xazsz3S74n5sOg76I8XeG
DUG4j5UYeXBYNeLHxii3pqW0FKFdQfyRfO69StjaXRVEnn5/Qnyi1PJnf74XzSeXU1fNNrSiVo/H
lH/tZkS6dUF3nAVemrjZjT9fcWN80++COU81POB0e6/T4drBGD3W5lUP6Q7JW5yzNIkLq7qrs9y6
0LFIs+vTJbqjxghK57Rw9q2aTNPa3aPNXiULmuL46EQgD1/pAwSb93BhnDFi0d62tIjeYVW4+RiV
jjc/NRQRfYLlfeY5Ro52jH+S0VaTZH7DRokwxF+tF6UHMBPFxKwgwYoWLM4r+b5ilvmi281x3Z6U
s3mMyJJgu/1EwgistRZKdL8HI+He72NxpF6Nsa9uosXXWx5bsmN7aZJEVkBJ0OqckB/s72+1rrQf
LSU49+j9izrkgXOJQq1fK+9z6SzUzHnXT8M36DhFnxY2huqlViiTs+zE3kJ4pSjoSM8W4+g+Gjg9
7URg0lrcx3WyDnc9lwj6qdHqCzN+anq+UTeBBvc1o4K/F3dzzhg4Sse8CZsxzRMWab0/cNC9yjKg
8xPVJsXifZ5kvxdvTmTMbzOGzo7FrtFX76eX5T10Fia7MB7caAvZhWN0QJ1b2X2vpuWEp/3bd9Md
zbrVUwKSsc2BUQa6MTaKv0RGbhVA0Dj9bJtiKz8BJcjIYh99CeogBWs3178q/cbUb6OU/3SqUKPX
KdPq3U8WkOZU3aERkhikcbgWH+3fLEnBSjFhJe7Xrr74ChPLArtpbKKWtE/i2SoURoUDlbl316bO
05lx/5QCQlx23alPoYvRygGbCa4npSh3dGUji6EGBgEsqDabhFjPfBVL1WfNS8j5dXpQV4e1CMTi
NHr3L0BbNk2iHzZkk8Omdj97XYYS9nX0yQ5Ufb1P3JtBGEIyQqUrZ4uIMlvPZP1hcZ2zESEDMwDy
sf1rwbBF/knDJK4kSyoOMOrcUHMl27zRx5Ey0pIwKCP8Dkh83rmDUxUtjIYTttqoreOPsLPvIDiM
qH/qis6b0v4IoSGjTe1ZwptAQuB4cqm+/Z5OON7N7qHJo0m8rWgGhRWyq2h+gBxzaNfx8Q7jc1xW
1JG/GrNRMSSnSsiVsjpET3rWk2WFUG3Cy8J9mBNHFB/1q2ACi/aWU2+mG1clDTxW6npczhEfCaBp
DkrPve9/NnxziQlLugGpBtc5MPftXZBi1cezIx4xpGSqbuDGbTysH6aCEGu8H+mtIs9ab/M8UCPh
gV66rh8kpVIDozEj+vGgcBwoNF2d7RiO3JhknFlKJALLFyOpbUK43A9OxMhmtEWmyz/ap56w/SxL
CxRXXkPzED1ULbVWcdB/83cXqmPgPwUnKQUBp8Ucyp9EamjrSh4iNkeAbO3ednrXVtDgGVo7s7qq
DZOcZbdAwLZwHoU3YtzW/MuYQgw7PZuWclofIRgHmpQS6YBJ56UAeA57EgOn47MxIZdoEcYI+aKS
R+GdM3DyjopIK2T9UtnZmDsTVCS+Jm0DVNVFeh8rICSY+okDHchtuvpJhPyKWF5OiiPtTTiQPO8t
mwPBCIMN84MPMzsQB9F8+yguRmLdy5G84jSpmERsRi7THJLG1tVkCvcS3KgIS3LWlHI5MNsqKEkW
P8cNjPLOpnG7Ebtdlu4Y6d2VuE6W5STvQgYuCMRbtXNAm2zNCvc1vtCAOACdJ2oyYSt+rTrYGDGv
bSqPJq6sJoi0kj9JUSbHPL4/26UjVNTpxFDZpYzpQoaj0f5HZJkK7z9/7OIHgp2LK78+En8Xu1t9
QRdFUBlrxmVGNeIkfLlqKfHFXeF4Ipsb5jhSWZx+idMc5cEMxG+Jz0FKnvhcehefc58JsewaqC7o
4Fy8LSPZOYnrw1ztz8l5SHmCZRTB1VFsIiP5sFOJLAgtFYa80muNkRi7bznqWWfBYsTgpWCuZeIe
1LHeKy0rOYQAWrAJiSKbwocH4gB7ON4h5Ie/an5hmoOQgVDQ1k/uNys7ncSJcPuwZK7bvvt/imbD
5R/1v1LZ9Xd3kAvyHtl4rM83B1jkc9qi5H2lF0eXGYxelFC/WGSy/zQWKJx/WxmFOAYTWOiVChXS
FoHuux94kh52E2G65S91Xjcq43hlxkCFBzvVR9jDKp4SLH5eb6iFtHrqltGyA7i4J6KvnLvYDcXY
RTGoO4Dao9qrO0tVKIxFyEzvvo6LONranpQ9UIVLqo2Xo7NZIld9AvJKlNnZqoN2fkB334Lsykgx
x6T/7TN1w9P58XZ22RcUM3+Ow3mKfLYLQLPrM/eSr6HjweExLtJ36myiJr8WlzmETLavFR34s0lu
e/Q2X78wgphvr+QgjZIc7hxmiMZGSG5T+skTHWTvPQ942ExIy7Y54PKhv6KOOAquPwVZjKS1IXD4
vrQstDH91z0iH4md2vOxzlno7ZTjLv6Bj74E+dxQAa2tBUze+xRnNpQGCBCFXbqbMgExSsnysjmx
AbH+V5+H3aY89b5b8Nb3EvyfvJDPaFSiZHf3cI7XTRpNN8AWFlquMipGlOlwKLyOzfzsfymkhi21
EaJwan7U44+zXgk7hk/fRMMG+hmjR/cxjBY6pTLzKZKBRAf4ojSXM/CPKYGcHpXXsq2nWpoqz9+y
qMr4AubG0b7JelctvDzCAAD9Hyy0V4DeWsR5Cwjz3pfJ3C4Txlh5gUg92ce2BUDAxHhNUMMaxCxf
m6f7DLcHoEVn41+KlI5F1kZgghbclJouqP1qDpRH7dGkJTN534GmvZSnm9i4qRm95t9cpQ0kHSCY
lTB5J/HwvlQtwsbyOunR7M2EwdO7ga0RBZmbkEZ4qstbru9I76pzkCnHh4+C3911B5swTGUB+LH9
pUMuPd1f02ZCJWAghLtUqPIhXaVlR+AK6wYmtxgnBuyE+8vm06JPSIKG5wzm3nW/lfM4KSpIRflM
oNdvb6fk6+IZrPEq1dqMDctGmfyzQvDEJByCP4QpvF2DhFgr+GQZszahuwhclqQxY9cxcdxSv3io
pffPlPjsfL7bYiDXs9eJocpIl7riEsf3eA7PAU55H5I6tnNXmkohjvJuvrpfjbrbQcTGc73CaY4z
bwPH89wiB40B4AntLu3Ft7EShzePd3sIlQWs4lRaVDQWmPVSOF/RVALque6WfTQPRPGgYGLiOslx
gMLQF8NgD3L6uHPCfApZL5YzgA3p+8mgDnE8fnfmcXymqByViaVSxI6Uf97VrJhNSH+dC63wf6yf
Ns28UJhiDb/aqH68T4yXifyTJqw5xLk3PgbVzZLyurRhet5VoRS2/BYA57hYxowZPF1H56w597nq
Wwz2knIsMgHrrlSmp4Pj0CbLcXv1FVzzqrFytQFLi/IB8V91GoFRgPnU1iy1aUlIkdemic9qTflU
TgbynHkK5g6jCB9b+mBZXUpiQP7jTwfh1nWhEYiEp4c8YUweIvlfKSGqb0eRXSvNxx+GwqIR4iID
RrOhPHv09Jv0v4HtLxwf6g/B50uk5FodQsbWmzJ4JWdtelEJpDJcPIogOgCs4e1xlRRfH0OR76PA
b9gTOXzkEr1ujGjDNlt4E9KDZrcVL+wuJ1ODHh/e90FRk125sgQb4zEeNd3Y2lFzmtqVITZ8vhyT
YYfTb/ekAGNkJMBu5U+RChHxKfxMv3zYYrPBURzFkvTNBod66bYeYDTCRu6bVNSP6zB6odAqoUJ9
/1sq2KlUwkVMx/S+RzNsZQSMMTXr8/T0b6TtLixapgX6U52AAsMfGYiULx+UsmYxTIanW59sNvTR
+ZKprqrguoaf/yduCH3MzpG1dlVyuu0z+yRGjz1UZSou4ZuI3p+WBH75KXtzCB9nJlp5/qlRqZ7R
VC2hgsMgTkQZuDQWv67fOi1xZ6si+1QIP56wSVhpeEwZ7ENQ943Izh0F6k9ocJC/ZIvAsscaXiv8
8cN0PpNLbLSYXcRc8OJ3waLj70mjCg2QLB/XX4DCj7jT0dtH+X530Us1NKS3g7oFOtKDoVtECIkI
HOlVnsVWPcHJOUd7yska0Q0eI2zW1gHQwN9jQ8u2ZsWdCyMcH6MRpERFALRV+bknPZYsEBjSOoye
MF3VkkxuNE7TYau/KDlNEEeLLDoEelZMq76WcSSBRg4bRH1ILxg9VXKpfII3OZf3OFCvMAIYq1d9
R7f+bKFUjMKiv0noypGhhndrGT9rbZ3Yrgfxm0DLhGttentBWJkJ6ModU2o+2FHlFBzdvkggRKwI
R+4NOn+OHz7TfmQ/2SEz4oWeaDlK/XmnY6vgizvOyfq9uhmisY8u143OqCBe2pbpzf4uag0q0cbg
Da2t1s/y65odiyybLo5YYLVYgMKMIohUNp5qxHUgaeGDtCKXSheJLAargeuOACRh/RFtnP3QX5ZD
XKBWXLaes1+q/FT4fkT/5Utb8/5SQr6xJB2kADs3pi1HM84kHd0DO56eFao8iXJqAltDFJdjstle
jTqmRjgx+9yUpErVYD7OcJCcz5dK/xHZEQIWuEwEcfgxqnV3n2dOCTn3r4OZkDTj5qu6otXuEy7K
dFAnbZvDvsG1mGY4EDW4AhF90ktU7BEP3RRoeMl4aGRf7ov5GbfhD+8zI/krVFIyKgrXym458iuc
wm7r+EUKuBNyE540lsN6pgSnafW8H6d4ie6TTc/lDQLBrCQUt2vu7PUbJQHPUqKYOle8RJ/oNY4Y
LZYCL4SfEfmwqz+0r8vcG9Ch2inA4ak7niyqvR63yvP8ZRA2VtMZRXFRIjKuPbruziDxWsr3kYoY
NiuHqwkTkREZ+DXMz0080afbfAg7VuzEqrG3SKtnQsBTthq2wmhUUMa3Lxi+Ml9AnyTudU0p9thF
TbV78dDcKDcZqpyXC/TlCPjTtZXplkwdzhO6y6e2UeZ4k5NotLRe1g8dTNTvhWbvSIam0zPJxK8V
XgSaTz6PtlVYgcdpDlqCdISieK1E/lWm5hPjIssQPX043slBLtD6l99Jzjbn5AwgUPo2q5VFLdHv
KzydLbygDB79y1T4/uu0KaZV9ChOtKZsJSWoAkLcGWTVJsxGJaiTSInNRmZbVvgVOFR14PEopUzL
zrAIuXNsXNhKZDASx/0FBv0h+Z7bXy/hfUepxXfsC9xdo0zEzm6kVzWG5+52Lcr2jrOmWsucYWib
miXp5PnCje0EnBY7fD2zt8s8MiWf+mv9UsbeExYYeTW1LOCLt5hsIsOP+PIeSYpe2wx9RO6XmII6
0i1kTXM0fRnjgF8wfxWD9vZgaZAKDfwx0qFoi9yaYjgs8Ykv6p8mTN1GqUtbNIwqNo1rwC5kE6ux
5qimbKGKPxywHSGgDOWil3nhPZyPs+r03S3WeTHC+QkEIAVHeKmC6KRxz56wvIUjg3mQdIbB8D23
ev+s/eUF6D7s/fNOBbA4XPUPOlQGBjy1/9yBGlqaocwSh83mgUZQJxwE8cS4+6wFCvmmaAys/Vwa
jc38r7lwokzwImDOeDOruKp5rgoJ7xYCEBq88Veyw5Igidnk3oQuuJJQ1ynRRuNh6pPZ93OEZ0Gb
fFarL3T5IJXi86QLocY8t+EpEtRYc4s+wFFUPEvdfiBn9QWLtZCxMrKkMwfBAtNo2knOF32lqTaF
aQM3WuLMDVOL2bUI4cRHWh5DUk3laa6lXtmYUrREvnuHLpDKLZsZWCQEswDbM1muULCwT03rqfKz
KeYkY9LmL+hra1HMXRWgNX0sVBfp3Nwu9uQIZjz0S45zyECvzBjhcTgkg9B5PRecsSWgZTxnB8L2
deYNgRixtRwft7t8bUIgjhaAEzP1hu9o0szWD9+3wvJNQtCMdaotEHYNiHWFRiev2g31xG10A56c
lRCON77G7yrajsv8tqJi807EYSjGjn3hWMLCA+xa/RNAJOHFuwX0lq4JdWRBa5MINqhUYOtZ8jzb
M9lhvjcF1fO3mLf5ovj9bR25PfdpTmQpbbQfg5MBR/guDsYwK4auyrp7mEt8GXOuboeUswNFPuL9
CsWwDRj3fYYcLF+jXbvgdkH5bPRqf4TCd1TXmMBLuSu5cpt4xU4PioavRgkOutqtyBTi6XFX33eZ
/KUta5ltk+kpLj7U7cu2DudvUwxM+SJoiD7YyEZxLLYRvPf3Lfh4MMhRHYXbHtNXX5LP9TKZNQBi
hf7qoDAcu68SahzUnae3EArpMZn6TTAyFhveNNsDR3dpPOdn/phcXt6Yr8rZG+khdpwda5gfDRsa
TRk42Y1Re3YmWhwEIF6ySF8oRljSDjcJF+ED68xNQ4opLmD9jNw6z9A712N7oZYxZz8xGxfa0o2v
WjkG3d3ac7PojKu+xUbTR0z9260XNOAriJzgHt7FEWdygzIhg84UGgm7tJSMdt15oS6QpXXK71pH
A3DbPkAK1ahX8o+DscIiVdPvmrvcWhFRl7fY1vK2LSXbEOACoOd+EI81YR5tKUqBh0ukDkSV8HU4
PUScadZnUgBd2pJyzt2x9RaONV2byyGAc47td7kSxPAWMCB1axuPbK3b9dlroRqC2BNhpD0PBMRd
TFiFaANt0447B+HFt7Bi4bBUSsVd7IxMjARbpDN+OzQspQ6r096zBmZ776qB/RJTPafPG8Zu164E
aFvTV6JqdwUTFbZOQXmM6aYF61hmNQzgwQe4BLY0ibfKNJ0gUIdFsad9zxLf2PPafTh+qWfHvgCE
VUfDOyuU3/phGknWd7wN4I+rB5efFnfouq4fBNkuYASKHaRyJy5uwu425G1ceaZq1nqpyIaGMKqU
gbciS7n6JTr4xz0HiwSYSkQrIOxO9jLD0BRLwjnufPqj0jgWXuDFC95MVYufXeBlDtUk63YqSHxV
Z5FLahQCWkWh+oXOrPCvwwGuPYzFpfpfRFLD2SBnS8ZUiY1H8VhuZ3e8YXadWzgxg9Ac59WnCQ2X
y/CauJ2sQRPsBsciB0Dg4jo3IdBaNRC7J4no5QUuokYax2DvwwVGgsljGn0GK35TXBDBlUBTBrJV
06jGpCYG1N4AE0g+Jg0Bm133RmSwMTJiRpFmRl1Hb953/iYdOIxRdAoCbvCtz8H6l9LQoTH7VMWd
EquuuOWPUyc4VOvuhJLRRf11zwT0OyRXxqtKMpWK5NoGSWaGC2vA8zGhCeb0R/ESWpPtHqJbwbXF
6moc/pyNFLVcqavlIQpG+4vp5Mve8ZwZxDXmkkQypciBA+EOREAC3iDF4uCKKKDmv9cXKHqyX5zg
Wpvp8N3MAPrdx74miMeOHxXZIiTWO4F2KMrYvQPP4y+u0xh+IbHAHUraCX3llCBGVOf2QP3wMg2a
wUEfyD0I19XSwqcjHl5yldOvR78b5jg4zrl/2c8Y3dAYJC2XK05zrcf61u3spM0BK+DAo7YIxVGb
4mODKiWBgDrcIaKRs5Vkcjd6GHNFvHxODBG1XGVrgKFvBkrem/ToPey84PERXhC/Jcmq4wJmGSC0
exMsXafBAIQRzzod4oxK33SH99jg+gZAMEdYy9tYzmsm4SHw24ilU+pDQgFClsoj0yqUJ2ODe5Sf
1lJ3MYjKi4QDezukKr8/rW3N48PVHCZmEkDDsBS4qnaAK58RTLyhMoKBcTI2jYZLxNx6lYJgBmft
CFyv6xPaJccQl4vmM+2XHfGbb1MnvZ6YcZEdW2Sbsk7px24oqONszhOdo+cXn1DUDQAW+sIVsDZZ
9TvlSVcVxSU+GXAJDGYXK0OTMvnEl8IPkEkiBnYf/ySqOZWbkoJEH2ptkNbjlyHmn5CiUB5pLT12
DRz8kQnwYfwPabTEhEasDOhnmB1WdfrzJo8bAiIoENdWyJuGddda3g1y6VQVcvHRhp3DNUCGABtY
UePokJ+tzzAW1FRtx2//dwdO1JXLEweN/ArwML++/6xxWkTDHrPH7qsoj9p8ZHxuppzGGUG/6LMi
6rOBX1TVYShTmY5djCc1y4S4VcVtgbMjjJKarkD1xq/UPSiDCZtjiKc6sOnCyM0qrS7EuN4qV4wx
XftgY+q/8C2JOk0iApLPe7M5uPU61oJ5ObjnENjlEJ/HNACtkB71wsp5eBg9niNWDEurygq86ZaH
sTmtCuddiet212AAbpvLAYEpWk0NHjumvmhIXIpRuCb86Mo61gH1+s1InmX2lwVeJGxfOb5P/xdU
5G+h6m8vgyMxKjRUbuKWx+OgkldB/A72pv1usik0zRYqvq7b0jWIcanRg0wFKL3/k9Lxi/mObxK0
T/L1F2QoQwai97FxTaGSnOXnwx8eeawNMtnSOMUybGBq2Yru5j+7UeYI0kk6ZthEVlQ9J/y3r7z2
PuKAmjadV+XXjvlPHeCoUfkFeUK1HhJOp18ucI1fn/0g/TR19kuuETgw4xU9e/Y5AOjpnmkLG9JC
61g6XoZBSA8lHK3ilfOEWSNUKgnL0qVWigxFVudxm5ktN/jTxBsOPV5lMyk4uMZuqW70s4Ylch6W
OwPZUDu7mcO2gBGdebdz1GEgn8kfu08EkMTZTfT7540iUCiA4Z1DANF1cWzmRAQmNqcWtyQsB6Ll
D9L5zI+kUxw+mZZr+jCMZPCwCb8eNVt812fDNWVkqlRmysQIRIm3xEc5xrRpaxx8rI/n2nbQFZC1
ejkklPkfrMd0P5htVJxmHnKI0RRyDRGOiKdhvr7Izugg4qrDQy0iDO7PySQWkUt2yTP5wTUhVWN2
oVn+awnFvAJaoQMR7WsDfIAiLRvpfDUBDJtslOgxSy321nQkdgGWkGul5GFhDlMt+aZa2yADqa3t
I1LIJ5Fyvh03lHTXzQZ/FfbRl0gTY1PX+O0ySO44gJiZRbUc2eluxOeA0uK6SARTxEMGG4bEv+pe
giALA/3gVCZTma6uDdsUuHqhzVT9xKT8cHlDQGIxBUqJ9LYl1u6NLst13UoC1qJrqKsT+1OFRW8f
W3bejNz+ZbVqHFTSA6+Evr+K8KPYvPrv/pS5VQYkh7kMxB1EGYEi/1r70iEiHg227YzRk4rl62cj
U5DYaiK5cAMC5AfJ0ipqgbsfps1tDe2YuMPrGKOe3z/q8VtFkU6PajsFb+9azdaTaCnfeCFW9tQo
M0jv7UBL+nCc6rgtvLn3nBxi6t7QeWfvSoMa6Lc9oJxTMqVPiabKLBJOO+GfK4rvC4t5AjRMIJPW
ak6BSCsoYjL+87+9+AWPP/hVVw9GMc3Y/M1Jlvm5wN8asuD3HwgIHPAtAXqmcevf/bL+Rd3jHYgh
DFsJxb1of6WtYG1WQdC1CLxjm5XEYfGBb3IFAMa7jDGUDThawrmTeq4xN5LutDPPUS2RIqNjBwhz
tppg2fw7DW+ir9e3B8dAAb3BU2/Q743zyQDp/Bz+xIG0Pk7yIqnQ8z7pp8cGslm3l1+YvaWNv2bK
2In4vX6BYkVjWK5pbs4NC1vCBVWk86F53zpYmq5WoyEoqoKoEfW/Y0II/5U9aMHDEIchGl8U6qGL
LFOFFRVShY9ns3h62FO5I2wclaBDT3QD2odEAYn52rs4Z3vrTAgrj5RU7LgNSNnWJC1nbEADS2oK
s18N7sJ+eTdosPdEfJ9tH+4Gcj1+PLedk3xHwDMmlWCwgAs2ZIpWTh21hPrepuTiA9oolFzXB0qL
gkR3IV4RJFeYzzldPp5pOLvcpN6ljv2R0BSi2EAvy10k4YbKaOUoRrgMif+S8r+3L4hB/5uYl/c5
3doWVWOcmsDWCFx+B3SdcOOIq7wJn9m+TXcgAroZxSudB8tlcdDF6r1v56+2OffIH4P1xT1vCN0y
7U7Cgo8U4Hzhctfb6ySnKvoI5VqI6WFSL/NCCj6+fHMFVr315qaocrWMVhStzBi2CU2vdnWY09HN
qE8MXabJASM8Mrk13ukge38471IPFLO9YrSqen4i4GtEyLEWeW0EkFlLiSdFUnLvIiOhW4FcjKEZ
NhFoGCbIV3m9i6SAw7Mjbg2rT21VI4eC+G0NR9hjzsVlyHzKzXh6XaekpZWGRg6DBThkSKp53e64
ao9ZS2gAPxf33aI3AEPFQupLljD9+jFmQB9XmaEdgZbdmi2GD3hkwiI9tbiXvPlV2afwJ3PhrZOg
dsTEC3cTnp1bAekKWgcSq7zh9eRZPoi+Nt9kjpky3IrUYwB0iKHh9wCB6X9U8pqbnAzlG872yaXK
al11zopbiu0jBP+rAA1jXmicrR1bBMPc3RHtJVdMJbMD8q63acgKf89UxdKs+05m/Xk0U2c0i3cj
J7DqSGEGWK8JJ+CnW29cTw93IGms7BvM9vnbi/o6pcQgUS+C26FpyjWWAGCr0sE6L6IaCFHtgEB7
ezv0nBdUrBof6Crr8kYNZW1UnPd5s78AWjQm6Q/zx4Y/kYgVeuUrzO5KfKDWiYqud/QXGHMD6Wy8
P4iJG7qwrnyx9CFf9DcFUmFbrrSw51S3hK9t+twRe2qQYsoovjLx1iPm0kBJ2HSgFWOAlP9EOK3C
4lMcEIP9Z3SBmDo1UrjSPBD2KEfETiM8lBe8ILHiBCncSZSBZVo2sWLE5/TeyGlu57gO+Nv1Os8w
1i9zRsRwXbTXJSQZ0eIlcxcIQr2I8M4/B88zorBWPE12jfazymhbGT9CEt+w5i1dZTST3gFlIdb/
3ylfx+/ETrr2hrHCzkXnxKS/DWU4tnnfBk9KPgkGpeZpCAlTwa6+tnuDXoL1dWd5TAWCaduJxrVO
B+rQrLdP4tcMrNziPgXwyOAs7DAdb3eNtsqGha/yJsRM7i551JAgr2v+PV2VXSFEJlChZBhQJshs
5dgtzqJSV/cQ3K0pDjMufgMqO9CEAHfE4qVwWhpC4dD3FNVKCaQ58H8TpULaOcp/X7MEkjPymPiE
V+bemjjegqoM3/YIrbpuICn3GojqTM2CaV1qSXaYuj/EISVSlhlv0wTIpRW9RSxg3kEVASA1+YmC
2B9lB71QOgVstHEKf0PKOaPfl4b8bDjAdCUeX97sgzkB9ulHAROgtrZCqE60eEJJKFKuOJYxNn/Q
Rk89i+bRlv5UdL+QaiexbQKl+i2FFFddh65ZVnoD/6qSwknR5nY6Jaz53Y2CbNi1iEu9YgBDMAVH
dhowWr9EhE62qCzSLRR5dXJdmAGG1HgzT6ao7c+xPfDl83tRBgr6m9jQNU5It7FXi8BOpoUeldJ4
2H6zTz4nDIXO/avjNvGxrAfPOwaWL3lkNAlO1o9W/BQFv/12nL/vl5Csvg893b0FCq0R26DHEEmD
DtD5i5Gy+XJTn/08z7xok8B6pNDYOWRIcqVvCztkpfb20/l8tsa1ugRzF9Rr9xDscWXZh8YvL4B0
sBW89Cha3YyQIn4o7FXpeDr6og9hwfiqER6oxIfmk8O1rVTPztzQtiqKi14hYWaLU5QSd7bpXTPh
CNcVo3Z8v29TSE9dAejVclO+7til815mZ3Oe/g0NP0OeY5TN8zvSxH2Kzr5OYW+gbJb1a5ZIMh6E
60v1Z/mTM2/7eB/OPqu7A+k05mu6H2bTp6ZSFn3P5GTA22DFT7mqPlelOx1gLTeDaLVnEILNV6FA
nvCyTdCIAaV1SjAroSf0ihfqH8TvarHgRaNcNOkz8v46z1qkwJ7RVzkFjaWkX3Yzse56MI5V9aON
3aiw0AwE7bomLuUvQ0aehXWyNJm3/NAw1nHkf0YM97p1BCoBsULOYPCHySt90tqD0btKrdZG46lc
ggYjIq/ircuB3c76Vj5ePwkmjVB6r1/yoAXhra3DlN998SSVHDsjM1xmnKbEsMcuvzjHx+M/zjAi
98sKPFNQzSfKdZOUjrSksFrKN6ZfeOQ33vbzn0UzfxhZREn8FbLn6NEmnXlJdrKhsMf5XehFHGnJ
Xhli1tOkGy2Z5PMA/6+aO9voCV53LzTUcGz9bt9/yLVRp2MZpoQ8Rz40Ti213qkVNuHsm6MX96iB
zhi00e4qNolt0zCiv5sp12zb8wid/amSfD2aysBbCf0X3AIy6cGSD8GzPTtYjtSSB2lqeA3YlFI6
ZB7O7Frcubmh25jTFZmW/0zH69RdesRCyLPdxDJ3g8I2h66mXCkFPW7DIACXMoRnQKuwB9ACfz8o
hSJAhs7OH5vCc2HY69rSPc3p4T5DoONwKZvRND/N4IVlE4UJX+EVO4bBxe4HH/gQ8FRxCWBqWnFw
7NaQDMNzXdM1TeBFd7n1KgJWi0IaGzA+cHQFTIbOAUReWlFzw2Prt12Zg7OGF6uWT6+tvfgzjtNq
MEzAR5rBQyMeoAc3nN3ZPGEKdaoC8GH0g1EyxKKjfQF2UyvolIeopmWq801KXrs3yHLeqOn1GTTI
f9bmxq2JDfGY7v4I2bD7OWhV1MRmjokxy7k36StxqcLxm5lMYg/vHQHSYh0sqUBygUqNuelhMWPQ
ZGysfvLIqRT8mipKFmDS9h1/JLdpOKrwZxd0OTu4Mk+v0xWQIQNQWRM0dgcbqh9y1UoljJBoBl6A
J3/hEy/Y7hnSBn0LXV+kcr4Y1PIpF8BIAiJMasRDeHwb3HYkSZdVnjaA/U6X3wLI/nr++IUj5CNf
816h/Ad9cI5lFwBkPIQaqznGgx34dBaGZOFV+qe7cl0JeqZpNn5l6848h4Ej5i7BoPDDA/6B1/D5
a3XBsdKnh/UMaTSgarL8E/UWDsPi+zqA9vBRcrA6RZjOpPV9bKpASjxD6ivWzGO+kywkAeAHwob+
uO1vKTcQgFGeh4Fmauo+1IlgiPOL1yZLURPFyziwViOJvVyMrZF3+ypy3iS5SXxHoDNJlC7ajMNw
LaBa2kkGiJ6/I1Te0t7fAJT8N4v0ZGZ5mf/8WQDnPsuCk01DYpriosLV/eWxT6EbevVQR0a8cXo6
F9rhBM/kz86kQU0w6W5Gqk/Mp3AgOJf8HgxOpZkLjJNVM6kro8QJqxN6q3thTtrYcSvOQpWAs054
Y/uR+tJc6auRAytQEIfbO4gURqZWtW65msr8C+ebh9pmsT8oc84pRTqBAJ64DWUqgXYBbTuHb9vL
/IiSCVz43AX9BG6uMtNYFq+sCmp2TU2FcnFhjJQKeA+baXuGzveq+jTASivGlnmHvPlYlKXFeEjQ
36y9sn78ebFyhU6MQgEbKOKm/ZgqZskHRxQn4F8aDkDdtCgJYy7bOVDBBcmZdy3SnHL8LmbmMpnC
0fept6iZyewVw40Bkb5SabnQOBeukANvsr2mNSCZGVejaWz29DhVgN50zR5KjmAjw2I2Fz4WfkNC
K525VaE7Tfoas9sri8B3QBKdVOFbeKCnyJ1EMBuvJEZCdmzrP53GO+27H+ig0Lb5alzyJmQ8ehmD
nccLdKpVHocHoMlkPucx7Ogob4QMPB+KXeXOWHAuEuoywsZr2G5mx+Q2Bmwe35+r6bfCNh3vkvMS
KyIVoOupmdtVN8s6ZIB9NQRIbAlgtQ6y6jRM1Dd3jz4W13rX4cT0aRGstbkpWun1BVaPNDqLd9gI
zbNbTiMxGFkCPMTOJg4P/0/iAwJtqa4U0tfu0/wJQKqHVIg0KL2i0OktXEO5DbmOPcORZ3/VVONB
Eqi5syhhIUp9fYKyj9GGSIB5r3hVEEKvNRzFfLTADu3AAv7K+0z9EEMfadrB+hYf4rvOVXpeMKJO
EfElKhss7/CGmpt5kPdcTXf92SyziM+8DMLTd3jWfpy4UC0l80ueV4xcdahcLVAh4Eb+RhgIBvhl
2mubHRE/mONtQUi/cvNGpE2dwUGugqe4xTXW3ZVDubqPWc8XSntJpSdQj/B9E6f/aasIgfEW0FxD
bmcg54AZqiqtkQRPjdf3XR4mFOims+ajhJpoim1KsxFbxUMzbob9dUlURVzXnUxKvvDPNhQqVO5c
k8rXvSCE8uOL4j+SDSWjNnE2jr08ePGbCzob2kvERi1/RVK8v2RmCReDbT3seKPbfbvB7bPtBY0n
UyxQvsdDwuQrTo0R7wHzGSfzPOqgTLlOu+Drbake4T3nq+1ubPqKZ8C1Yxb4QS0+qrNFMYR7rL75
SuiwivhirwxWMccki8D4zCWCWkTq9L+aWCuIpALOZNR3B2oyTeTOGxlUVT2DeqOQCZIAf7hkuu6r
GIJSslkRzxmp6mqjzBX9fSL1oSbmTTJSkPjGplVkezi1hEEu/WifsUlcmCq9cbG26nYTe6IMhbHT
eepGALp3L4+iWgH1jQv1uXw4k7ONtXWXappCtmTs7vRJLj2K6/Lfe+imggwQXRhyKeukDiIdZ7pa
NQdolf2HCGd3qxEq4g0riBtrsfxsBL4S5fi3WxKUe6a2qJqSYdhzQG7pmEIzVhzAF9CWlUEJsFTd
4SvNmzfune+R6CpB5u3U/lh9iQ1V8PB5trwaPQu+0WOVw7sD2GO5Va2frGF6ZNkwWsLdr55cZBr0
4QHgxN8IsIUm8BfRPoE1gN40p2jqzp184oU7Xq0QL4yX6qRJRf0DCxAloKQrTsVx6LZ8SqbygIEa
9m9zNN0OVmhKviHo72dcX+9jIZiwe+FcMNk0tGnE1TNLHxY9dTj5X7cPlJn/4o4G8QJgUsGTZJSQ
44d79SSjgxscC9ZWdNlpSY9qRXU2aG1e0nI/nQxHnIjGO9ofjE1NZ9v7ML35rYeZFQpmQZKf7hzZ
0tOYeeLczKkYu+tLNbg9m77DJbORJZ/4gNFAtQNp09tFw4O79P2e2r8SyInKv0nRJU5AmvK/7uVh
QgtsU9tsH0SmL9olBdTt8D3KAFH61aWIRx2tvlQyF459Zd06O7oryI8ZEE5TjX0UspHDam+hpc0I
VkrRqRv7KbU12whefAXPBkbV8ZRybltZTjeaA2tjYYlzng8kRhzojVUL61RhnHgjjBUKwgJiqpVW
GeGUu41plXwJXl0xSYF2UrnU3SrT1v1mmr7DETinud3Pb9h9YXWAHU+2n8y4GU1zwD87u4UQIJo1
AtZWdYUs1lLdZ5Q/UwOBA6OXz2rLYw72NxknZpMrDeSYEmJfCMJO+b+KL1RA1lFrwlOEtjGaYawH
dYcrW1o/RPgjYWXcF5fF0T8h5SuZOiDHG9cWM4hrDCS9m2D+VmuUXEkU8CX7YVE1j7N6SMu4JvEt
NRQrB1INt8GjEyTMCSuZjhqZrDusSuUWgv95rrFGP9gU+jR+JgbHj6XczV8MdnjCEQM0rPapABFy
qkR9JaSGTKzrwAb/dJ7S0AIIEnWBEmNONLej++4BtpqekjrCSjhjLhqFnBPmhrAPCS7IEhyjuIk6
1l5DHuTNfkf7w6bqRPhhHvJPw1ktucmMGOLlHQ8lKR5af+JoJJzUkfOKIyoO25D64j/TnTV11mn9
weaZr+G16T921uxYzL04uMpHY8eB5qDkkKTnG7JxnkzvbEgK+EoCumiplSZE70JzpmtqCbMAk9gP
0oGIKNvgSD+/urg35Ry5zZgWeeouQn1ys3VODZ09DMj1Jyg47MHqj+Fyu2MEfzkX9BDj2GHvtcH/
ChnY6rtY1pGjiGN2/VK0c7/VIxFaGk1aF7UVBkEV37eMNa2ntq717S6Lfe9n0PJMxGo2X0a3Y9TB
iD/eUSqS8DNuSN1Z8L21P7HRcXQuzg39RXhHWVQjhjg3AsBPUrFxp4EXP7Zp+hpeNdKBoMELbl+G
xnlfF6afJd/8yltFkMIoKjvXzJVL+dQvdZFszlBSQobYiHtXjMZPy2whfH1F9fT2zI4Nm91CqhGy
YDUnp7EbU331taEFanE+qhwI7c0fjcPd6QuxgfGGi+oSPIbS/UrK4oE34y9D+C2A6yQonbulImOb
xzKjyJYPl6HpDd5c6mQgijH/8L/sWUrdiTD6NnbyZLqPGx65NMkfE3hbRhyKGmfGk7EcQXzW0JwL
MledEC8t9rk7vDyf2Bniku59bPSTbJ4n6URdRBWZNRZKPUZ4PBoJdKKbcexujI6QKMhmnMd+hYLk
mC2T1UOmzOyzbbUPz4NBPD7ojn2cU+Y10IWay+Z1kh7/3OK1P/xTTjkBZRDd47p3I2lrsXhLYlmS
vcHZKsx1XqA8ck/BYMUQ8pLXqnDWJ35hF2uOEHrl99hVRQLkIvoWrZ73Sgsr1UuiBu7HtTVLY5kt
/ivsCVmBkdvP6suUOTSQZjYaTS3w2joqVRsekue81nOLjVRR5SHEdQyVKmysEeCzC9iifqN2JI5D
neHi4wL1+DZzLt9E5J8akYKiveAeGivfEaU2wAamRYPjLYwWYlqCApkT72HdL0T8p8CY6yfBprM4
AhnmTpOvH7Yd/cXzsZUg+AlZJungTUFMygy/rnxIDGHcUHP/oYj/mwrcfl6E9kuiOpjl6Kc5S20N
+SDYGeMH8uka8UoufKept1Pu9F+hVSDTBBiaaJht9/53c9udDTTG2wqz7AER2pOOooMvEy9a2bfg
K000DrPkr+fHrvYeXTAUnG7R3NQthKLShLpo6qVK4wDN32SsDIUI8Zb7QKMTkVK/emGnkQXGIX3v
j1ObrNWasKiXRaGBYM9hyqNQFkMk9MHe0wMY9v2yp/GCVaODritYnVoeY0ndQUzuCr2LBZfCAmZk
tck636DcSTpljwBS6mOpf0e3Tvru+jYNnR+CwGLXE4od1yzOs6fQ77aN/A4/6PJ0PeZUfOpnnWjC
y3Selx759ETg9pAyh4EuJbQTLtY6QLtyh2AXIPSSSVNstyQoVl8zBW0Wg3jmHOv6uMzGMi3IRPIT
fAOb74++QPw9H9r99E5o7IYYiubarUL/VDf7y1QPvfbf8XN2S86Y+y7fgrRyaT/Sigae8JcYo2XM
0kWJLmfxBidOk6Oauxiw3cv6tYeHKR7mgSEU1PV41dvxBXAuYzKFobZo63B2y0GeHVKcbscPCJaR
xZRX0r3tcvaUSCP8n7BVXz6VP5TSZWz3rLuin2x6HMJMNPWZzXVfiw8kduYcq7p4PkHHHkI/gknS
eRe/z+lzVZHzjgehQANyYK877rsbst63JYqqUHgzU1wOw+g/rfYbgJBE663yTPH5bUpnrFb38kMr
+W0Kn7nQhfUE4rMUh4Vf0G6/iS0ous637W5VVp9yb9sv2K60W9Ye3i/1ZemVSpATXFIx1IxmqxvX
raW8au3UHJ6EeX+dpZQA4ayskY48GpoDAEwzfBrBlYwUAqPBXZnNj/JBXqXDSs/n0L1S4l/YFXnJ
7Yy/dAQJF1jN4iiZwoAAc/kgRzTYy1iwe+2054VY1ar6EXu8kfBP/jXhSHoMs3x2iLlswGX4M/VX
MU9XDKWIpvFEhIFR3M2EZxXpFZckJ3yuItIookBRtBgKbTfxs5lSOU3RJEAIuHr0Y/9XctpK+WwW
z37EeCWoNZKAHUl7xfPDOnLooFsIrLFGp9cLCwFoiN5K4t0MikHVK0Frl/1hJbwMuxlvsVLykivI
Eo8vxAr4EHZgVHIAycJr5bG1eXob7ZwTQb6Esayp2nWYwbR1zXWtu2j4KCabn6Dbh5B6Ou6Oz196
KVriSOrlmgHFhafNR8RZuL6ka+5TU7pg0WAlx12BZT8auVCAad5ArYl6OSR/SexSy8xhV3Sd08Um
TTJtkypeyBMZUnVFRKVfcOLCHqTCNTBFoJ5MoMtYRD8befKhwyZo3EBxMsz8d7tPmyp55i20u1wn
i7GhwHZr6sO+OOSQgXSQB3tGdlaGnE3VWhLW0ix9nR9SI7PuswlKHMihxEwk+8gaif4OdX3c79jl
2cjdBn/nv9KDWEY2qXaNI+tgNPTaVc+H6gc+xYTlE5PvmjRS6gCzBmlxYayIz6552ZR6a1OhKd7m
1+0Ro2sVrXQPxXhwucfDE8PEG1dgQClYX8oT6mcdL098yW9MrytYVoXiF1lvmPEkdEnkU6QQCNTw
W9eiGGnJW9IgcruDtOVzi9kAZr3lbYenLpG6TdWuzkhjytinwOpUxB4w1JVgdF2QScO3LFuZrxBh
eFxSQkYarraX6wqRSCmb8k1C8hKpLDCyEPbNTsr8gMhktbfpDDvs4vfYaP7UADLIiYjolopeYwil
GZFlPVy6Zfv0fLaHw70GMsXPFdZni/LNRua11gyRRQymeA5Q25R46R27rgDp9S8Jiupc9WqKU1Cy
zDSON97sIYFw+82ANndV+l45xqk0X9QtbDb7PFWvyL67zi1mEUbUVNz6BfmJ3+No0/it1KKLBizE
XKTKyIQTs4m2qT04Q770xFVoq3yvPiMCBhZvy+sv6ZWeAqyTa0BQHJCcwKUWVAtn5iB6mU15ZwVn
zOrErpkwQniA/OX4vYPCt0DLzSD1yKJKqPOKqAn02JKIxOSczRXYlclhvX3N5p/2oduG13RqZLJP
aPbz9qpMR1kDBa5qZ4uK4pfsIWFnEU8x+4ssdKTcjpfU/GoKNHEYfMBN1aot8eWOa9HEdyrfr2NN
f+urljhLgrX85fCwQn/ViIW1tenEZVxtKYPXFZ+F+Dk7uXGjnH4PmFmymvcDnr0s20hpinK2eAfI
dkLZX24thLISbehYz26PX1xf8ilZLO5ytilYJnyA8+LGPbslE7txn9OpTpkSsci8tavIe/YDKZ1a
l1C0EzJD+kCDDP1Rfb07mzb1XJBneU7Mbq1KCR6JBa/QioM3bv0w/clZPNYi2SZrNCNHtKVzrh6C
5kR+q993IcKGVQxOReeKR9CEk3MJ29rQevyO+F6zYO59R28v0y22tji1I9Tt3dUnGpfq6b3+vxLp
/RQloc1qt2nvVPCl4X4WNFhBRmu0GfoqPqZBuWGPc6NJg9GUCTgeIOK4KC57kDP6CoT3pRv0R8qf
pb361FzztKOhSm+RXL4r5f+T9gkXgJDEyA4T3N7bxPOiPSfpPr/+NsF22MB6HJKUhmEcGf0cWa/6
rFpHQ4DEakfWUTdIY9OzXpda40X74ivoZa5MhkCHNXgfg10/CWFa5vIit+bRmBZ805dQrsqGlZwu
CJurpdXoOT6AZugZFM1YaH8sLTPeJ5dXDmUyItiCTpT3tCBXM6HRAdEh21QcwO7BW9Rk267mlquX
Xk2ady6Q1qa78JT1h5jeLJpJL3aYkBOBlyOMPW/puNl8y3zm50IttdidD689wEHvCEzAoAphxK5n
7hEK8TTuPTjZoBmk+bBZ1SBAzpLeZgLhKqvwkoP1msHZ5ppK6YX8zrOSeXorz9CqDaVRCUUJtMrC
7nUm6gS+S1KBpsxf5dTsh+P52MDhO75+fgfETjFkNh3iU72BtmcrWvuGuP4dtziLoQ/ZDW+wMjNl
QyNQVRKM5DED4Ima0upsa5xxw/AnnkXEab6GH6rbF+Wkc+5tURSpkopjhKx0lPXak5tzzY/t09yq
Hn1zIjsIniePpoJPLcyI5C89sJqusph6EbAotMNnEWQvKV3ThP0VYIEekbs+qZiJ5AOlxA9MZEHI
xgF8Bx+NmMhqqmTc3TyufCSQFCbm3I5vdUizi+AVsFhWxobDNG8Aszxts27XSwvqFU5ul9N02ky1
KnxjgIreWqip0xjojDQDl7mFg+HAK4o5SnYFNoIN11DoaSt95qSr7fi+sexsO+/uQfvfo48IAdnQ
MUf+6SknLfzjTRtDud3s4fdRS+53Wrs70P2RUw5LRFpEdg8p4fBW0eoqeMgzDEoXbSton8tUGSoH
HvuJGhDeHhSvhkQfFCl5Yj4MgOfJK7J+jpPrdQvpKgXqp5W6hNtqrMIzovBmki/fjdK1cpMUnthp
50W1HehBxsmkk7nOcvz+2WE3/crsC8Mns5Yfz7+3FUZjThCGX35UUpNvld8nIh4OsIXAs4T82P97
6bUk6hQxiDeVYNc6qdIMSS/wkkIQ7RE4LY8LHSbkZz5DsEd8pnmCXQVbY9MlVFR3JOy22dpEasPs
QlDPoGVI6dYCCFNhiXtwCY/YRxA1MYVMRip4W5ZmNwoa/mrl9IOJuGxqNsYJPX1+XhzXEzATzMBx
dbjnYxd8vTqKFtcsy8eqWk46Y9PYr4FtdrsLy32Oywq86SzrAlKq2Qe1iCRKKFt1baNhA6hLDvBZ
GlQvx/9yQ8s+wWjQ5RnpHDL/nOtx3UYT4xdjH7/v0OIMCrhSPeQgLjvKyqdvIbQAxSJdpsDqfcb/
ivWZKQU+M7fz2qw28c4Cg3RC7PCDFHtDEjFl7e4sJqkvVMt6DJfcHijthgQwIFwWuCjzL4fqAkRo
Zfwvxnf797+8raFhOCBiVMUO9Giah4HJEJguzxXMsPynz0ciBEcMJTooKsia3wReCG55cdmReerx
Yqiww7M3mPYexYFON43NrnwYpFQKPcZcHdKhX66ThcC1jaBaQGpaVFlJCHrQyLusnKcYj8tA+D4A
G0b6qDq8wUKPLTKhlrXkcZUKKygQp8hV16umhRLnB+T41cP4Ng2bW2PiqM++6DRKW/ajbrcQZ4re
P+ag/EsHXxtJuPuSONa/MRk8OxhsL6izUpiEo4oVlp38FHgLhP129Fu7N/ciLC8ZZDjfYwp+hDVL
s22O8ppsvLVCHV6DR7r89xPTScF/veW3LXUmn8E/5TwhVwCZEA01sj3nHE5aeqU9GS8t7kdSe7EF
wlsKo30MisW0XyoBInGQojY0Z/CgwHn1D7DTiFHw+P2kcgcgyBr9R8ed+0C85wTg1UNR/YHx3Xpb
ic9U5hdGpj/e6KAV0ir61DHfY/LbJ3/oS61HkfSd4ybj7gihX7E1YKM63YBhVg/W5mL57H8Hz/t2
ji4eghVS18fjjUvWLgDmkGH1ZRQA2c2AHHsFz9jOMQP11tZImD3RNpGVkS7FcNuCogM9/GXZMxYT
4S90vBsYTIHRjaCUB0j/LHULsxTYBzWJy4wm3VTZ5eVBRNyO9ctrJC1CE+T/Y4ISDYuqclPa1U5m
0A2+Rs0kBvUNrF8Ae1txoRngLBiA4Zz/en/ehlgEFYRpekBqJ87yNFpwUtYtSkY8CORCWkVv5ZeQ
fQB4Gknmo83N2h/1X3iYgk7PID51KKEll96IkEMTkCoXgUaHS6lXOO90nHDGTbhL/L4I9a6qy7jl
soZ36qJ7gJHyOa3GcMofSkGWiI2CbEct+ctXlRmSyKp3xrs4fx0iMzfdHKQj7AuaG83Blfi3I+/W
6UImSpbJo3OdlRGz0fZrHHn9N7GufOBcTY+PmwAWd6k1CE0m4mbD852yuUPkOuGiUmnqcK19uAeJ
jl9RCdXrhX+hOlClw43K6KBCmMIoTtfNPXVbZT/5vu1PeOnXrwD7qAmWNjejfvzX2zbSl+lSrKC5
TNPGOVOejsBwsW0hiyCK08Qu/Zjt8weBXnzqmJmyaXkPOkxScCdAWDAN3u0/azu28GLupY9R1lw3
c5Ru6bpUpX7R5w174BoSP4QeeZEDjQMG+IOApqxzLPIENwsGvxo9ZKGUFIOD9EF+KplkAYJ7NyED
Z5Qgqvhu7dunbmGWhR1gPEZilc6TNTvnFYpIWrNIJWkoCSYBqgrWjm2HtMGr7HLOcTJgeMyIOQqh
gqq05swVzJZmhhuVoc+tzN/hsA1/i4+ITO2EsurkshD4D3x0qiIqMzKW46rBXmNiBojpGv4NPbw6
jztD8uI0biD43MS0Sg5oFxpuPEi6xTTjbT3LCQ99dfl374pkduYsZh6hFJqcT+tiepLAuQL9JO+6
4wDMgmSR07gYqHXGf+0Q3TlmEwgbqDeaQ3oVE7F32BG8P8PI+cHEnIPvexUyQiWPGOkt3X/QiqwX
JCijawn4OqTJawOIHTahIk3rikXGb6kX0yYr2KsiIcN/NJ5G3FNeq13vvjR1HJUUzoNTamoiyO8e
Q3djhbMI+EXiV/5o+Gxhemr+HZsaWvLBDun1lVctrm4ShVbaV3F0Mkpp4CFbgmJRBEMXNGKDzJH8
IrGGSF8sFTMaZ2zRShigYdZfYl3zO18BykMiyHVAG2wZkv/gfqI3ta5bFQBHKq4GLIHTmswiVxsX
JsBk3gRWSFHFrlB6DOQUJ9c/cq90tD+7ZL3OXfdRj1zfa5FXI0/XBOeLB0lIP3gD1BN1WyizEFRl
D6jFr5peDGiOHo6/+Vz4eAa6ne+oBNV0L/VzH7oYm6VmW35X0fbCSl8PuKLGPrxDnw0t4FzfQM60
HlHoBGi1r7hNois0ctft8bOVIJ2hYB0vgUzW7r1Bp61hDvJQOqXq+gwtgSNS5BzGHBNibsWgoiFq
umtGIJYowBdJE6Ukn1sBf7tfhhPoMciOaZf7zBzCulnHe8eEA+SqHIBSTKTbmsQkFgpQkOwWFZDm
SW5Aymr8eJ4RhHD4lfJpEYecoREvi7Vmid28IuVN1I+UXAsyIlIcBsdz5efuq8cCsM0rwBq7n+HJ
jAxc67zA/2HkBDMrOVQjvehAU6a63Ofyx0Ahqfy8yP1g6g9KZmgyvwydMbzdCiFjdrw9H41fI/M8
feK+bpdZzFpAfMfKJxkpW8V7/octn9s+P6Qd8R3SZhEsu2IA72fWWZR8koYqnSNuHR0PCVnRCayy
qHYfz8+b2xHuvLWLTeNGqr9pJvf8GXDwjN2iIvDuMeZ7f8w7y7uOMC031QZVHIfaaFdqlPHzYWA9
coyoGcFVT0PQu9iRoINJveJj0vbHWhYeRYYQi5f9aKAV7v8rH5f5YH1BCPnG9rKuq+PchjIhVv6A
OkavyruUHSy9w3D9pa81Qms69CgBMXAjZBGBP+swfVAzsNO+YG5N2nC/DkdMoN5Ysb2dG/en3S72
8721yrE2lCTLLT89/jgM5FNH9IKJjjmdAOvqQDDuV/OS1HdfkkYeq06Dn9GOogL+zZ1UYSaW60QD
CL7d5WZTxdZaW9zDmXpo8Bm6pXG+kf5NAdo8e7at4FLzYAE4mlLv9hwhjsNZFE15g4ABG0i3bUNR
WdXdxuElLy3/gztg0P3hHZRxgSDyNpy+u3c1j7p77x4tUe9ALg4oezKC7268O9zVGyJ/xgx9b1Oe
MDTBoiiXa/hNy5tqvy6lSpdvuqO27JS9ivqt95sz+Uxvq7kp+lGqMjbzxO3MH37U5vDlbVPWs/+r
FZ0zBRZCiW0DFDe8xQHZzComdzWtZ0QfSu/6SOEkHfuCXPZ9Qsdh57Yy4mAZccQo/Gw2PMXiOi4k
tK/vipghdJhN4cTCyEPzW8O6t4V117088wuRX17KOzNtUDHJ4PK8+cN5KHprp2xZiuF/DFjm36G3
0yyZZ0QLbPPvdli56CC94r+5eYipwuwqxKyZ5/oxt0pZz5d2ACkh/lL6O/s6blwBeSz6FDHFf5vR
ExU38fmcOgjzY9/TPsvqfvMbpc2qTsUHssTDxpGVMRXG6KZvtKH3v8QEu6RU6Dey3F3Dut5Yr51H
iECSdTthnMSqn8yDi+4kyXfzNotYVKeCYqSoeSxHp5xciDI4Kf1wnEDtO7tNJPr1mzY8DdknNMu/
u4H7dVPVR+M4PKlYA/tZi/Ovq1vs+emR3G4fhbF6EQ2i3keLu3HYkA8An709wKGkVYbFyuTVncRw
edIrOwktjvJX1BAGXeRpKFjyBBdGuyNppDsG4hZCJCbNxc7CromDITkCfWuV/k+vlXJZw9+isrPD
XptSqJjT5mUpnrhf2/YwY7pZQt6s/cxg4o4pGzzqEsEfMe6TIaht4pMRd9T3uhWzhmfQZt3/JKmr
3D5CwPCKOGjm5xsExSwHyXreAdSxErN3fuTeTEmZ+7trfovnJS06x+XGWOuCP2DgQcPhyhreBGxZ
dNVW626F/M/80bpYZsUSE8+4RyIkDboKZTht3dDHm9F3PJEGx6WC/q1AJ/yNsVl0nO8nbsOVWPRt
FklBpTmXfpv6lZA/+FUeRRuaraBv0oG6siMq/82gGi1LRcXuOmW5AcHvz5Zxe1emQw9rT3c4axFM
BZtfgjbrMd38N3rXlNDgJebmxWlf6XazkRa7TV+Bj7TEp60cZENNJ7+NOHzFZ2IItm2Bwd1HbRlb
TPYxYcqfdXlNyXzOxhDyDWwPwtzSRerN37e3WkP0+ULzImUpWz3JDDRGXRuduzKyl9nsuapy8mUn
fQPO7QCMk6NoobjFHL6uTrNAq66vF7sMmKE3zDvH4ZfR5M6m2uoTggWBnHO5xtYgSWCgfR2XMNLQ
XCfEaijxjsj/oDoVBz0CTm+H3ieYeZ067hAgl3bJvUTDZId1x9kFLQZixNWBQ2wHx9EPo/pLj2Lo
JtDUnX0F14DEIKvZTEGOyt27sGn22IDCkL6s0o4GDIQ52ZVavvb44I+CclnifLigaMucDYkvWBbT
d8uDt64e2dP0+Yd7TNwRtrGE9NvzUjG6GIDxs81OLUZ3LyEEKXz3a74gT+ubtp39KygEsb5gzMe4
p6PHILTKfPyxZLKwsnmyCotdfqCfvmtEQdyy5FRxKfVnP4PIQ/Zm5L+K36nwAYVMCRESn0R89Lt7
NHATI/Nn8QLgN8anbrwDh69FU9aO1VjpWkpf5gttFWyWmSDrZu6IK/kbrlYAGmAs7eHZFGLICdIP
+A6HSFp2kxktOX07Ul+zAEBNY6CcL8hadYyI2WOwhnfEN7gPRHrpBrA7SdEMk3OStpUqn3UHC093
GmI4XB+LBeEFfzi5NG1N5qysdEkUK0VFpcprg4A0DwmDgovcZswhfVO6gLkft04hvT2+zy+99XNP
POZUy76StoT3DolD7B8v7dp8cxGpprCmP1pbtgn2CrWLmLaoFANJnBRKxG2eawUelJepsHQpgcGV
h7Bc6AC102QWHgYR/O6VQJqIY6PdnbYp8Rspu9+mOJV1dF9ESOOQBSrQbzd90RPoISdBuuj69PzI
Dd7OLquwtrTrPqbxFkYo//PocE0NdmuuxsaenWdRnWRecAbU0gHv465tBOqoB0MULBWMtjzLDzd6
eczFeCBGslUd+pIZbzdMcLsf96U3NynFy/frBuzDzjakZTHbww2s6HTyO3ZV6WakeiyDfjhUjIIp
isUMRZKJURmOxHsvBHq0mrwX/qLCC/TXw8JgzRsOlxPTE85pFLUEoP/Psqb0Cj4c33bjQKD0T5UY
CEaq0nuTEyzcnOw5J9BE0zrOhswdbEWsXskaf2GeMFR0EyMNuoILNFuJjm9t1mtqje0lGH1nNJn0
9f1uWSA/2AjLRmDS7c5lV9aeMoEZrBsrmFtcRu9V4Bq6zCa6WZehDcp5KBYVqrHfsJZzZ6eJ2fGE
Is7sTAKAhsT6mIKV4Fyw5zYCjlqVKSkf3Vq2n6agsFZ4SbhTi0KDVrDEh7dkSEbPOc+nFhWug7eQ
kVoPa0cTgWinbXN9lwZZ2xnrmSVByTjGjQJdrmrCtmce8l1CltfXSpaQggUoQWwf+Cwle1QNB/cr
+1GAj1YIsQfrtLcDXquu+orUUs5QOlDBZueXn/5v7HK74ht2CkiBJ0v7q8vNQd+gLzC1I2S8osrP
QXSjNa/cZnZ0peybZHa4HJ4OkgVxCu4+uIGG0NbkMOujurkS4JVenzMV/7e/T6Z6SRcZR5tx4AjT
37khkyJfYs+Fu/IkV5hOsk9dSXy9MFwEEqhQokvKG3tebgcoGJ/2KqVsaK7np0a6ixTWsdjDAlib
tNn/XTZqdaIPSfeb63dZjMh1TS8UpzimpT5asBDs8pkN0ZuysJLU8od/m2EfY3fzChsDKwgb/IFs
DdZBLG6dTcr2AkukqCnpdldTSMS9ABKE4k3vVRl9mHA0hkVXO4ZzbCLeQ5Ie5wrpnT8p9xeKgKzU
72bInD91frt797SKFlzV/+Aa1JZw/XwTGzOh0cuVSklwsVQPNpEyP1ESrqMF1fZksAghUvESneiU
2WTs6q1ykdOOVWFRRRbOr9lrS5IeobqF89eXrl8MROI/bawxVLRhbpsL1X0mR6GKY7R/O3vrdsJ/
BSFggeqViG1DiyWDLo3Lqj25sXPNlJF985DNyIlXvgXM2DgC41gATd/Cn6GeIcG56TOnIX8kZW4+
XqTEOoWZAkHRe2hHDcy8P2WC/QMhr60Umoo9PwTKmagCyxGCX5BQ7H0UHGzIulm7catE1FQUBXH+
705FGu2GJWz/joXT2R/hmTGVgoopdRuxNn4ADqymK80o1W8B+xJTep+LbJ+pBNsS320D/wzMuBBl
Vx5D2XDDHBBQN3akwhAWktIl3LF55f8tgHLdhQZzsbr/ktue75LmV+Qa4u2/efbrziraiG8GNMl9
JvmDYOdaGTAOTWttk4sOmaD1FQDNJnC++zNjheAlxpgQneKZMmb0r0bbV9UaoJSyubNkyOfIzYwE
UYRk8QGSdxzUYAyHawMnw3LgWA0XomRa4scGIjjF+WrtISXOhdhEr0OK5VViIr1m7IZ7K3t/ED0Z
ZBH4Ida/UTsWza+x3kKn+EepL5w2esfH1cLguO2r8BMxmwPwlX+eXL2giMqordSaR9TQqEskALxi
3Tl09D8dN2WEecKrhlsx51EWJzd/T5/0AiAaxxWh6LC/nhLhRuOqmkAP65qkKeEkl70telzFGAHZ
02Z63/lfeXLR9cMfZ0CR3KaSaAow/zXReZouztPiq9gv2qkRK8P08cZjxnkgyxXECbHbOjP6L0st
xcCe8l2r7DwoyxZQ8qaoN+i3EqZF+NVNDVfvOHO/633OvU/PAl4SFyjTREhwBqQsF6V28e4mHeRC
3tW9QX9T/FX+V9zz8VOsLNMlro7YxC8jgcgpk33qFm9XWnSV5pH1HMGA0ykRFvzuZ6c/MHXz8qht
zBx62j8ugTbDF3hIPAoZBWGydNNB11SIp1s0GVtp8bqg9nQaNjXLaXA3uJBuG2FO778EwrqqvPOO
KwUDv9gJzbVtLGGUHAEBJWk6WwhOvZA2ZiCBKwG5vx9gsySDt8uWXw57VO+wuq6bPEE4YMT30Lie
An18ccn5Dp/HadMXCnpP7n0vQGGwyQW3YjfqU5Lolj0I6xMpCWZwDQ76X28WQOcP1hbHRuhdAmeP
VW5duNKDrzhb4aCbazKISHBc8N0KgAR17Ek8enW0KlSvZba4+Plcrz+Z30T9F/fD6/zkOZIE4jvn
NLGjLT/KY3z7o35s0RS2bMzgtGGNK2tNx6pE8os606r1F2StWRXet+O3zOmj/5JUgQODTzF2/ZJ1
MiVtOaDazmfCEMV9umQpuOFLlhqDP39hzbYawxbkCks6Ky7u6ntUeW3pqvzQ1wwYaRC49P66o7Sj
DaOYHRYshHsrfxaBHJ1fGn1bSAsds74QTat62U1/d/UrHCYRpgXptg3eGOXwfKEWfCNVp0E8CrUN
TQv/l3yv+4lwPEMUwaeN2td9NPKAMM1v+qxaw638QFQGFxeYq3PFcwX4VxT8S19aNEFU0Uktd8No
2ZNpIDfwMafc6s5kjolMYOxb2wvJV8r2MF+Irlfqu7Fb8d7zZLwHz5IpuGwaaHjfhwP9d68H+moR
wJRDEyR8Fpw6dv9TCNdiCI7rnEGfVux+ALtGKlJVUeLyRzgbCQhUAvy02TnR4W2axa4Od2og2LMB
SUon8FBIh6hAf320Ua2nKhFBhHoJ4tjOGJ6Wd6M8V3V6GKtJIIqFZNFOaFzb1McYaZ5aAcxeUp5C
MXhAhOaZbtCsCS5YFVQ8IHYS5fykAnAnLVMLWoWoch6y1h2KH+ng+oWYJ0dsAZuelC5nPE6PPpn8
rZzXa/iR0kSwbxdDz4uFl3xBoJxEO4j4c4V+MePl1NKZMnsstqdI8Mia0N6NTgZEQQJfwaF/QSLY
0gT81TltR6iB0QlQ36N3ex2A7yt0Em1In/aD0SEbM9TWFSoKVI/eP1TZwV80ld6Z5g5XXIqicN6j
sQMZaAJWuzsJeSkj5i2Qfu+Vmj1uEKWuqa7zN7zYK9/7zzrU6jywMDhxc/URiTKz3dLVSOSxilNf
7cDZv2Gm0yq6Wo09Px0l8fn+nFojFHWP6CzxWwHIHaM+uluWY7j1rf2lUco/1t7QYzA+Nd5uqvis
WvDZYi7Wya5Pa7mLpBE0TF8IBieSU7EfEhHjAGTKFvwEU+HiwDvmcvZlB4SAW1KDj5qlnn1LmzqE
5KnuKy+gfl+f0vzCjfW8vBMshFANxHTW7tzVvSEPCgIMC09T6Qo8XIhtKtpTiDdJV897x8K4jt8u
+smSN6Ag9oMzz8ceUwmz51AXyxchv89kAdUE3s+XLACLk9XZxkXndeQhaUgsqNq0Jgbgw3tbDGcc
fEblcAPpfcEnYa2AIwJaZcQYO8s6cL9jH48ZG5rTkI85QGT8IdquTQpDoQXonqvPhT9a1F5fTxr/
f3ZTS5JDHfrTbZo1J/Y2As8NplfAMTLY0GrDHxDdL7gItFJKTOQm+0JOuh1N7M1ECs24dlbwVwMk
JLkKTemdUX3XTot/ezlywTAlmYLoLto7OjXC95YVJcPxv4mJmbfNoewCsPRQQzY1EN3p4S60a2X5
idi0304x3Do0pH/vxOr/22+CfhmP0h8KqfMvlKmXisr+CVKXCB65iawCrw3P0KHa+gSmifL8/E1Z
gsTlYQBDCZEZf77Pu+aUfImF71YtPTce0HcguN2o5r9ahYTCpGNJ3ZFBbL7UURUHfN5OpLXD4hqy
HRDWgUgdbeyeNrE616sxf3+hlWenyKamic+b2It4cTTVAjlz/jHlxXkEYSg8r5O1djM1jOM9+XK5
FsBuq+SdWmpGqaal4HtdB4m+l+siwuuLzjdwSWOW1r33a1xf4F4gfJnEwf47VTpKzIz+4X+SnTBU
82afYBjgBAEZBM9n+5WuV9k9qxv5nZllP/Cj4CZOs1gATc+BolPSR9Bae5F+GouvPjK5OxJRjzw2
j4Ce1LAvH0c2VDkH7KRZqdrz0W4jGguwRI8yGKz3xsOBgbN1sH6NdEwH/uKqiiyV6y15+jrhoK+x
mYX7YM6mhRrvrktKJ+UNBIPCq1+ZKmb2hhUInYs3GQUcxnSiADg6iDpLWJ8O2vUVE5gE+ICniXMG
biyyIcCPSfOebb7Z4UujsjLbNbqabA8VZ3/g6jeDiPySOSHkaooj4V1QPVvRFy5Mg9RQ3b4FlIqK
ZBRdpatMrBPucjpv/OCHJXNY0iMe7ieCViO8kF/EYk07OTLxRKoummtcwPTX2IB1MBUcRS6PFxN+
VoMlc+3sXm0rslQuJA2YpW0ON+NOBFgFOGdARHDlkT8VTIGekPNpeQFr2uScqleiLo4ZTM10jvGy
o8j7N0hFxH73LlRJVzwlKXM6b5LC/guK0anqpyvjVUnWrs3k8EG8FQnYkYJfIbv9h5boXkGEXegS
6VaJ/pAT9ObnuksC3IOuMTN02QjF0omXS/KQrrNzZQNbT4aZzQtqlyXAiw3K2U4d7HtTB1WvZ39d
yrED+yuBi4qnwGKMvCzVZ5iJlsBlxfIn5cIeOs1iys0R21vaEiUkHsqAodNspL6Pos8LLLnqBmL7
X69PaXuCpp9kE61FTaoHw7zixVoW3uxS5LpnHPRy/B6KN2DH5krc+m68RmDKHZ8+wDWOCtxb5ur0
mxq7Ir9VjQQTRMfXramhS0Efure91fx1qUV7TKFCynnv1484cn+hgeKial6p9bRfipCNohgWbPcW
/CygAgRtfGfzEvBgpuh9ZAUm56YXyHC4j+8Ly18tJWi+nXHqWXpV9ADBNuL+58KMrG5zlSGwPtIg
1KiJ/b/Am6SYNkFDeJ8M3rrAMu+2s0GgpDNx4CR3JlZsJnTjq3FoyRnQn648B/pg6EBoInEyIx54
ytRT06Q6kQDqbjNrPGKl8s6M8R2WvjbzeHgn8DmebfRd8+obQ+Kjgmtnhx2A9Dnr8CryWWwgpwxQ
IMLegqsWQSa/+eDklhMbJLJJPA4/TLzZRdjdLdytPic9wVld2ViJ4sdT1QZzICZz0BGoYBXZkm/E
bL6tUDJXX5ZNwy2VKpivoYVwJ4sGUjndEu5BSbLDOJfhWDaHSjZANxrKYcc8RhVIR/+wmUXeDEmh
bM4olYyTjf6ssHD8zIbdGEGMIoYdHyLfDLs4vHZoWlDePz8FepIwGC1Kl5X2fLGGRXIXsZYHxhHy
HN2h+0/pn+qG3xFqIwH4tmjT72i9Im/5a5d4xKcRVRWaUfD31z6EE1tzfa1ArreFFayLDlpCzJD8
G89CDpAF9bzzeLbW8/4w0O5hMxYRjLQDi5QZEq+gRDrzCGS6kkSoZs/WsEEykAbkrdNYIhSZqHYD
cHvqzH9d+P77rekrUKBESR2/0VG02fkWTJp1ca0cSyiAoVWwzvKZRrWFz6rZgjwPbRh2PUE/7EeH
PQUtPu70PiAG9fKde19PYefRT8zM4IgT4XAegEe7o4aA3FUsTBvLanaddq3uHRbS4j19LqymzAXj
77tqNd73qWbcJOU++mz+YIeplSpbyEjyDDG5JDtZPbAQoArCmOvLrTuYezQBJCX6sNC1stzSRuc9
ehnZT9vT2lJUIpaj2mZ/hMW7tBluIHjS6xF+ioCmWsaM39of7tLUsFi2Vyx2CPxstIovAOCTyoSo
j+qHqjSfBD105BhZQKx010miptwdH4O5AtujGVKPNtsgP6Lal+iha7vJLLEJbBBnDHd2VQtGke6G
We87FRVBbvDM6pvusiKHb3buJvummvvYRu3PLnXma/8ipJZngnDGvf+KF7ZkHAn4GFnIBHoh5cxM
sUuogfqxkyOdEN8TAk782Jgz3XTdWRNiHQ5C4kWbCVO6R0/4VtB+0Sl/bZExaO2FplEGOo7jl9X2
LpkwgCKqVXC+fADFd05+VJW+RBpI1XjDl9R6zWux5Ef6X3kzKdxyBqxZxtlp50VaqkyEvmIMDGWe
EFpst07vpBK653Y2eAqyrFgOcKTcbb3+W8jtxBV7rueJP1MDqpc1lPEPKa2rRSrxfQvR6V+6CRGy
HW0XHVowXWcNVaqVPGaPwgWr9X11zh3GweXsA1BjSO7+PYV+8xbc2N7N4dPI5I16Hsn3TF/zZJto
mgeM+o+N558Y+FsKKyyuBoM7z29xeaNHKSVf66ze35SxItRRCZFlDIarZ/sE/FtQFiA7SVPGimES
xA+ZMP0pfcwOnI52zE3Vo15sjdUDeuuaeVfzVkA0DLBKq6dESeNfqLEZuyvG9lq8eC/JHeRi2e18
Vp08cj862jjxrWMGW+/QbuPt9vEBtDgl1Vohi6T2mAyPSwB0fd1YIiejyKpe41FvknPQtPAkWXxk
zY+AbqZm7N4M2C2olOvKvU1KVULBRumZAMXoIuoFMnw8jvFEvNMLqTJpciMjd+CX7PbssG4HLxMe
L7+ezkjD85wRjtXv1qo21vbX8l74W+7Ew9sIw0qZJ1hp9hI+FMKbBGCNi/kyE9jhkWGV6bFDkgEK
WtbUi6a5E6sNYHXqNX/cuE53Sa7DMix41X2rZPipWDudJvMW0Zx/170SI31JlfwexD1adXK8PnFq
4InwCuN9GyZR3aot6pLw8bGfv7+EqG3plYuX44hp0Rnvq5LT+ix1ZqE+B+MT7x+FCFLJvdpfgbCB
H88eGvmiIHuP1XojuEYZhXpjfSBYidYNhTsrFyVXBLYlkEvT621oEv6/wnCwrVqsLn5ADPPYpBZr
MgulDpMUO/wfubKqo0XTqh+l5PyQk3cFzniBcKw7oeA4THYeOOfcgqut0eyAfLcC7XEjZ7UDiLAD
ciAKgNjVahDrvVUr22PTRpM24Jp9FQfk2t9lBhJK8EgiKq2crer/ywbMvdsAKJ0pQAd3d+lbe7ft
HotIVy0mvshaxODOep2bm95Q3U/kInEJgSAc1g9SdPfoEoWX2gAQRD33T3PBS1n07V8dANysQNRA
m7QugU2xkZe0uzWf2EuMC7Rsrcwgg1t6fii9/MNZ3U+h0t+Mn9lLuf7pZiq0g5hAHiKliPVyapO7
1XyGYdv1pg8RNm9nSYCOqZn13unnxSeWWqHYKyX37QUktuItDabbk0peK08Z95bxxSP6PEyKNnnx
XoYm21PaF8ZGND42gAJBgpIgoGnjMQqOilH59aV1DDzVW7vLeNzSTrGtI+S4hIiCI5TCCagqNHvP
7m1GRkH/mMebONoMJIXBSD0U1iLcBSKo42fuOaN3cLNVjC0ojDBDfdqHmbS3i68V+T5bF4s1oGP9
xKbS+EAFNdnnNluftlxciX0qwdoTdmwFb9rkGNAC88/bXyvU4OGw2PUJUCTuFFuDkL0ZA93BIVWw
IJmWP1BtRrjqgGZw+FlEij7Pch3sWjWE4nyYYUWKeYK+dqBsZyUiGhbPsyS7cT5F+S48ZJm9Arxn
yHJKrtMuxBOEkXdIZ6iUZU7UZaDi95BAWX/+lAK44EYH56Wi3TDb5f0d5EtoB6S0TRGHAUZdXc6n
UZtVrAcovyrPmrA8r12Cj0Ek3Z8iVyKijm5lFuE/SdlBilvSkKuBiQSaCb7DQBHOruE1rVlRC7fp
5YBJHMlJS8DADT1NK+iHag1ctobWkdfyRlDKnXewSN8mpzM9cdTiqwgin995L4xofrO5eS3IwWk1
v757M5jrs1NcICeguPTe+Ejo7dg3dr2bKhQ4QlWbTw8QOrc97qnghtlLIKSREfAArSU3sKW+MR2Y
Ek7R1rSOFFmhJcjlbeydNFxjWwlTO96ydsteKIjlV7yq2fIINWkL3Hc2/hcOUWJijyv3Kuj9Kqic
8OaLbg8NWWRENL3LK+l1CKL7+x/mzrB1RV0+dGrn2/F1icumlYHh4IbjbbUmeygD2Maxwe8YxFUq
82qggQ7Zw/c++xWLCX837Msg0jHNE0RZAZYUI922cNpH9V0GXt7WKLmrpGE9cUvjcnsHmVbd46Tq
cL6HMPNWrQir9vW+mnDV4ScAXV0/R/jW35e0pi9mn6VKp2fTmDQaI3WfGLjJyNrh4ps6tf99ww4f
QJ94YIAsSChOLKweUQdpFJH5ZtU/2hseIgdPhYjU7X0Ktu3HnSjLMk6crT18KZfLlA6yi0e1U3gN
Ap87Z8kVf9pmSoUCZXYEGi5KWtwWxiYga/8jO83mgHPhm4+9RLqWsuhnKbN8Z00Cx+4gZ2ZQjV9K
u/LzyMy8YIwBbF093h3bf2fEbYveuGqPk51qQizZSkMfSf89Ts1bBt0jyqlnw7IBszPVenfovqtQ
ClmNX6YIP3ZfyCazNCtVtD1/Ta3Br5RPSIfh/TtiSn5Lml+QWbn6dnHwPkkXWoXrUftA1XnXa6FE
9z8/QABIwpwwKA+z8M66tJbS878WjsYHhn8XhDUvhprAoK3Nz4xi36JEWacSIcQbahV22G25Vik7
gC5PrOldf+4pb9KGYEnxw3Z4qeaSb6feFQWsOjAIw5ngnnfgU3KpQRL0VJIqGS/WKEZcKal/qKyn
gtRrsmlW2iFg4YMZ1xkaNhU6ov9Qqn28OtaSJjkuUIJPPpfyBGMXc0N/u5z6XcNPmpgJFEDWaBYR
l17FoTGEYNyxjIXkco3bV/eOf0ZRme5eJLq4lkrqRWiISZkCskO0NnoTOGA2OUbwtKX0GmQnJMzT
KHj//TulkjyapFGTM72dc+1b0yBTSVJG4HjT4sFXx6t1uZjdDd+/AlKOEWWyXRpeaRl5L0Ivx9Aa
+iWqUC6x6kn6LoLEBWM/VBgHUoGGD7rxU3QTBJXpvvEH08qCWHAd2Xihbs6XOJx1VXEAq1fZhia6
d4vodwifjVnpBwT46PJjk7xl3m8Pi11h/fM1bUKqkP82wvveE8OU+bU+OEvPvisj8A+ISbPA8Y1t
fqNUonKKAsfQ3fNMYjOqw3B2Uz+h+kO4FOI11etjdglUonOZnPROi4F4LTOUCfA/J6lRLS58Wfzw
G9z9f/p5dM6sOO1tMFvmCWgIjj8/Srp46iYR4WbPBwf6z5lJ5iwd+ChC95oaiIwgyCMr0JosSLFG
xA1Ovmni97MaAba3Hiyb/Oqw5BHyXRjt/zIQc+2V3JI0gh9qCTXQl3sJcTodUVJjMvg9ODdurb0U
4Nw8KSFwvtmMbmyfWACdRBzv/gE5DU5rWIIWqS5YyJRdVnOhSIuxR1hR55rP7Sq8buSRecO0RuIT
OAlG2Yr932y41TWXmGVaqRq0QpnPhKnsWWidmnmi57vm6MLYWcYILmxYDKpwvBnf9O5elQiSoGiv
ZMJv7bL5rYDamGhL5sm/YFiF29K8oxSYNUxfhi4z3vBwCcuKTL2jQ3OqC/JTamOqNrvwjhiYm6BJ
vfdFdRbZE4EMW3jQVlMWnOUgHBP3oudCRHYcNC0FBrD7JOQdlrd3uk8Tgz/8i7FylgCtr5gYMF1n
nsBy6uchg9wHRri38nwivxPQtmZBY6e/3Nir8zNvu9dDREy/YNlY71sT+RR80u//DnPAGKJGgl/i
bd3xaY219prp7lcg3dnzfWPAOFxDEOr3D0oJTDrEdQ52e2Z4wableb5PGpiatwkXGqoWqx4bV+uG
Zog7tlDmO3+5kRD/7Lz5bh1Tgf5GEQjvumKBKYdXMHPjWFKhIhoEMzqD8insmYM0FIuEnQlf2g5l
SkQiHmzVYJJR7caTT16jTbf90HMLJlFZNYmP3zKxamTLT4SsakYhc5aEeOpQc4qmYLXIjppTOr53
RD98rUI0ZK5W11R4oxZUQBzN3wzS1aWPrPhK2HxMdGW7/DCfiDBTBAwqNxd7QHuyumFygB9KCr+c
NQuzJGxYswzRtHPoVk5/HkR11UzP4PmVjwOuBx8PFgSlhhDVrSepFRxeR8yOnoeF3PpOrYoxdLhe
eNzf5ToD1+7eh2MQM7BFm3DjiOHLMaUWBjG7sasGP/GcR/f8Skp2IMRTeSVMcObfjRiCZYZ+pgld
MyPlbqQgfaJPLJR39tTNJNpfOJLOS0sxSeJU2TXIan/QW+Y4WfcjCp8IIhQdaDogQSQEDHEAeV2l
FT9XqXV+yqVB8QOaRo4XAGa265+M7mnCc1cVCRINijVgRFp91WxAw3IoR5NV6j6PBQX0DLjhUtsL
21ynbFfHNoHEKsAYa/ieTpsopNheQMsM27wYAx3zJVoS6Ho8SmdSB12RqvF3T067CjJu1nR66BYd
bYsU5r3d4N3cKcSmPKZd1Kc+h9GOtRMvfgM7riekeny17xJUjrA+SMWJ+PovX57RoD/QJ46WsaGn
a8mBSM//oLW9ut16DWMyWx0Q8++ZH4vNf7XInM1dpmctm1VXf+OevaaQT32bqTSDGka3JYWbvM4Q
FedYHlwbzqA8nzoNQqNjbjsL+VpeCv49SpVIputEl4P3pwGk3tEe4w49yR3h7TmoSUTBJYJ7e2g5
p3AcWXLRzn9F+RbbevOKi+9tAxcQvvPOY09971o0tRKrmLirdJEe7A2F5soKMwGblS4gOBZ5yk3s
hBAxZv8Amf6CDwwad9HfaV0ucOmOwMGw0OD/XVyYOOIt98M61vqMqT0fRrXOZZ+FCPn4iN3y7CHS
DOmfHbAD4H7pKXbpW62UGaZvr1r2UeiA8Va91+Iju7WKZycW2MOmNo28ySeUQa9R9cHnHEpfugp0
t+hIlgsiBOc8fzeSMmZSAUO/X3Ii0UtDEgQmgF8ubfECUqgmVnqBzQAPel5AoqxWaCtEf66Nj2vX
8xo0VClw6xW4FWS5MfQOnVAqLyhKQq4d0Z7wxo+T4AL98IwVpQfSYV+oFaMYFWaSoWl/naABy6yp
gID4TSd+6DHp8tY3rQOH1NkOECxeIewUDg/r66hbgEfQ5oP6MS1oZyKqCWrQAsS/YuWWfwZJrXrx
AUNpbRDXcTZnJXiUOuE5Bk4UawNu+rTO0kSFcYR9CkUkJtKC/Me8RfHgSZ9iu1hWekGd2w7q97Eq
ehmXLMplVj/RZB4kHqFyHyfbMXAKAP8Ypjtllu8v1ImDK69YKszaN5MTZOZVtydbTIamzzGxgmGZ
xV4ksVnf4iXOguYEdEcGvESqvpefiC1IQZf8R4cuxvUfn1xEtqx7o+zRENFWMVyzOoTye7gqJtfm
I985hQcbKDTC2l9wNStHk2EtT39Pom/QC6LnZNaguZgyyxuxAD6MbUW9+zUk/MStwMY21nS4MPvz
RdU606p8ZbPXD/ql+09ufGsbk5zrkvLcHpmMiIrB8uHT62z/0p9ZhRbtnoPUzYUS0YLffPHDRwpN
xw7IquGWOVHPegFh5XcKXfKMhvwQ3q+R8RpH7iJP8Y7pO1PsN91zWCqzpC8Uer/esJKUCqzc4LF8
+kkWMqvW5G1N67fGn1W6XmLCX/o5rp0aqYp3XRlaIeNTYphwskQXHhNxVH+2W8qhIqVqp5DHKSAs
36RburxQWanvCf6QbwKynOeAXuiVdvn6S6i2hNYhJWXxeftrEbCbxao30aEGXjYZ8h0PXIi3BeVn
jsQeV5XHF7TE5n+zQhNyy13oIofPL8EoW7YFueTi/zoVucG4g49hkkL01f6aodddtQOavdeXFy7v
aEAfTksNEwjj/tZxcOgNr7U7fR7YRZIQKV+JT04qXTv8zLCeyh52PSHds7JHEy0jWGDRPuKbXz7t
tljmQPjQG9HWJeqZkRBhsshX+tzm+rMi7yWiHT+nFlYS4wC7q3WEBnyLNE0dI5HZEfg6x3HeFeQg
aVp9TVb2exORjJP8kep2U2R7LHgz4PzZEaXpTsGAHjBPSQXXwij9Ag5O/yGGhh2zU/bJ3edBJio0
ex41s8tSxIR66JCiLKG9/dzxEsBSRJK7lNDfpaIaKZ9k/1P0AsWXBeMXpgSHEXe2M8n+SHZLPlrO
R1/syVq0yGYwwnT42h4+AlhMfpB8v/7f3URZGWBwfLpBB4Hw8jJgvPbDb8GaqZ97lbb5m2hjLXHq
9vkw0fQLeFE1ud4utJmEpFiBX7I/ATpOet0SZecP/Zjk4FM/eeGBKiPERHozFuZL7mexBkOpVS5a
3iXen+TtjUe/AOnuqHSscKZa+HA9fh4i+t9l47MaDIjIJ9JPpNBy7emZgQsXCxlvvDQAp8EKohV0
QW/8uTCv99D2NyU2ZG2mvgIWi1v1iU30ZJP4WmA6TcAT4vRAd2fyryoL2eFu5IZUo60MGBT0/jUw
7Jz2RXizfYDQauH+aBqwqQmHoS3LhIjHUk4EBJ5PIkk1vd4sw16Ez0+tMAaivqPxucIMrf++L2tR
1NfxMXJB3nebO4emYm1ptoYb81zn1yL15QxYFJoonBPYWKbRycaZjLqAHXfBaypj8WjC/BuaGIz5
lQuWFLPtVZK5DnCwvO6v4CTq0epF9O3jU/OFWZf2FEBaYt5nI7mUwltilcsjj+BvAQm0KAK91at7
rNDaOdZNLdFsgii0qh16chBFudieX0qUfUV2uEi8axxNRZ224sLqEic9WOUpC/iuZDHuYw6che5R
Gc1Zapg0kISH0IWd99qo0xEgyyBlcqINtyUBjw7bOxiAEGDnlcKI/AR4B829c9elLElBMbDWGn7Y
2Ypn/t5fdgvoG8rJENj6eXpysWFb5zqy+jCjkFE/z1eXt0TcsF+IQSnAVuo1VF5FNU6msxbm2t8T
I8SBF3RgWudnIQtjizvshBZZjWLY3mT/KP+CdqxlFUeIo4QrCyvEjfOFlPtg+aBCNR4T2YJ/3Pun
DK2FYN3gdvgj+hys+jzeCwu7O2tmi1fXvtdEiuiCEEaIIn+z8G6cCf/myWCU/k707zcHNnThDNRw
Z25UZboJdSdFJQ0DNd+Eip1HFs9FMbIkD6EBDjEpcevIvMYfz85vgyU9RHN763HPMezLnL3emjdy
rGNbIWYdhqSlEpCf7yWXV+kRUTFeTj1uNW8gFcWi/BVPtz/biVIerTfNjSc8Fy7G2eyEyWzyhqN0
v4BNdYsvLby3ehcIErpU0UE1BPjDW8JaV7QJCYY7waucqvqvAUCynQRFI7ImVwZ7zzSwk2k0A6Wb
MqmzE6Zz/FP5E5Hwo7ypBoFqtV26V2ZLfUWjdiQ98FpoLV9Hvpt37HfMrZxuRib81xMZk0/Crfdk
mdV2YJJjwl192bn/pk+82K818cmBJAIWuK09nzQpKDxvuJ/426Z8MkiFeRiyMmRiMcr8KgvkVi0L
so0CE/gs5UDVrA/4U6RHnoxuMrlDD2M7YIwWHpGq4qHdI2jIkwzzT7dsa8iRoKeVHQ5GLxZ9xz7i
x472BLeDpSxDTuAkHGKrRZexXnaxm7Zzl+jyTCPpXvnEt9/chR0TWeW2F97dq3XUVymXiYzB4XXo
nKXS6pFOJi7wXlBPjVKhoImjiaz0IOd57Xa4v5PMrhi69lKCd5kuo6d0IXm+n7jsyY8uAYLT8GWb
MgjVvZdjZrvZT1QQ76xe+sowWXlixg2BHCFvpOMZg9SB2m3O37nh+dNwfRXRAKBCCU6QSCCCPYRh
5sf3nX667RQZ62EC5dtImYgYV8jqxjzuBSwHxR88XG1WMaV9KDaPEAZK42De9f9p5a+8AsQ7n7Zr
y3i1UEFARSiRuyqz/OBSF4PX+sn9M0XWlX0K7CCpR3jmW81xIOoCbvPF56xvHUP73PYNT2unV8TJ
MWlP+sCvrYdB9On6J1NISFt8AC2BdlnuOKAQmnzPh1tKvEQ1Y4KQtMAwzg2k/Ql2UzyMx1p8xQzQ
FTIW+p1wcrIK4ox1p2Dg2d4BnazY3LEmN8XMNIJabsQMjjb5GBbfFA97DqeiSJOOHn9+8nJPn/OC
vCCjcD8f+Ql1DOIg875neQ3I+O+fpiY6Kwnm63qCYNR9BIqvSUpswzxG/5DmTTIN/2Bx6C5bKII8
cSaTTTMu1dGnhR3TmYOnTOfS9bG9x7C91M1sDI7tKa/P1wGwxwAKxWzDARsdmHeWKfIJxcnchop7
ptbOidhdRHNadbpv7EWlSZtboUpCF3GjyH85etg8ybyFdGA+hv0T1sWjZlGPfELLMcKXWbvLtzSr
2AlA9tpQWD/GJi0BGNiScV2uuhWhzCg9PkopfBEIYpvDtPCh9Ftnol5mp4EQ7g44xzQaE2L+TlGb
9gPovoYoET9DCWOa1C5ZAh8J/B2ZWx5kS8viTC7K/+QDrBsoQnRQOF9JLv4buu7VZqY91embsryR
fvxUBcR5kzUrzq804Ar0bCzq/Q1JcX6ZnHECrkjevR/bTTggXTfZ4WS2SwmkeyGmnwH/8Z575Hi1
8qwOVwaLNOOpQGH/KwkRZeT9xXEfVPFSs6RGlkh0sqRbuGAv7/CwDRd8jqBLUh8++YJp+s0F1VOE
bE99pvh5kxTzQVUZE3lnrnhiLJkXU38VNNWSkQh22h7Ssz0wNxOdb3Oh81hVRo4bajEhIrw7bb7Q
Oma0wH/yhESUuu+zBFZsWPzsIpWQJgexeWt+MNQImKQO9s8yqeA/VreTHmb5OWluFiqrBac8EtBi
JNXvfOsmcNYSP0nlbYPfIQvT/mooJsPpkQjQrLW2gUe8jDcUEHJZCSgs2Z4s7rQTpR43POBLlPzl
h4Gl9p41yevmQsO7yNvRMAyFQludC4Le4ylUsM5owLXyctr+N3VGRDSI2xVr9BQcHdk4BiP8kiT3
HoZfoYDz5MX9/FYR5ZgKSfMZZto+VEe46jo9Wy7/DabhSya2HeInfmpqz7mePzeHNaDFARlA0ovN
JLQIPVo2taqaAT3tuKHKs7sDwmBsE4gghV+2k1dQA30cFuBgkm0Rr4CfSctnj9dJdKIpAzSOE/KV
p37pGN/cBSMli/mqnqMdWkgfyDptYGx+B/lWV7xc5NTDvAJJcFEwrVzbZn4fvId6Bb09ftpm5b68
APwh6RnamxAbVlincdcuB7T7CORDzDH7A2f+n3xG1as0jmm/YpoZlCYgVVmbQUpAHNmQXdSkLxhs
TQKDZv74wo0rRxhd+23b+K/EI6eDteSOAuQXKoahsQAwYN7LPHx1UpUd42KJdJ8ZoItaoQ0aHuG0
piPj9NQ5ZLBXrtFYETEHwYUf7TQ3Udfjr9yOG4nG5OWYbhip6a5hbG7kXYHKPV9vPhan3zxWQBCS
IMSrbVdbud8AAVa0nxrlQTZRAybQuBej9u29Utv+GqiEKSgAgy2U+j3/jmPg0DCCwQiXyQxBnPwc
yQZckO3KBAzUULrl4NacK3y9w1JclH7zNZ9Y3PiCNrZpMGwOgN2UjLs/JUmMZEmtuK7TORjOU9s2
CS6ZRXmvZSdFaNHCQkP7H83htLECNa7qrGmh4vSkOgrgJ9Oi8wj6huMhd1B1R+/X8BbWpvbMwGc9
grZ8RZb4KmSTwhMsOzqJLS6xTVQ8cQDGI/t2+vtzD2rsojRbgtw/cEMCnz3PKhuiOoB6xgN4JzC5
PrAoxRbTiEIVvW9pJ7fjErdhYdgHB5HILW2jfIHQzeBAQ4wZg7wZcyr3QOPqcp1ZXpZ9DCa8E6KR
uLxYyd71bSm0/+wHuwsp8XbWfXSHykDreBeLPehF71GgRhgHtHtKEfI9Y2KJLBIiBPhvgMjZyDCm
bCFR3dP2pntIpmsw6IP0LRShIBUicoSYTXP1b4ZGTxgRH5UEmJV0BkL7hZaXDRPFLgG1FQDylyeL
dTIR9QxeQEDEXiNOte31HFBZSEIL3llHh4nW1B+PJxWSWsMzXcy//mfweeoKDTQglDCKReHJ6P/a
nCv4jrSd6sAqCaKW87ZhQo7i6Cmrr+pmthZAJOpiTFcZvrMIHmkY1nDDMYeC0R0gU7SJ5qRsYhBy
nezf5oSWNdxvd9VN1CDKYaRxvCyimr3vkv1o+M7lZqWvmzgT618mCORAQhzVGt81W3Hs1wYalxRL
/bqPzZn0xirYH2rRsxunqR6C/9hjyFqgdS0/7zzbJIWr+paKK/+Gak54ferZhj8VisliDhak84Uz
+27G1JquXTUPF7JUKtZloFFzEv5wPsM7GB+I5ic/74SRulsjLGj37gGblnpJ/KOCe5qI9l87JR9N
rvpJqYHGyA7Sslde6hPixLa130Jl4Z3pvEDjJB+1pDPVXFfWBZULAPT4M7BJsZ6ZbLSK98R5tHq1
HHoHV1mFc+TLklejuWY8uwySAJzo0zfmL8mHJVxDjs0NIIFytjJs2VwIGolSbPvLn5tlIQl+bS1E
aXfCl2IxKw7Nh45LDPtfOc876bnvuDrho6N+L+g9L6p4M4Uze1wSZQlV9m6De8dt02XGclpRu7K0
iw2rdwx74LaTKICmfoHnYKF8B40xsEGleCRGIDVnUweoRLEgEiuzPZL13W0VtbgkDYtcf5r3utiw
ZL/TsxumfotScHQGJHO4i/94H25OS3KJFD8rJT4jMZ2Zo1U9tLwise6Zh1dDhgy5hjj2GpzWq7BC
tWXAywLGSP5iBnIEgApjcomms8J1cx84lTwwA7cA/n5BZXuoYMKqqMD8CzBmlHl9lXf7p8ARoghh
UmpJk4ma1voEbS3fKjmOXoAm80VB7fuwC54U4/kOcDNu2vaPNwAfq90czcVC35dXnjSJMsjo5xgu
h99baLaioBBcfB+CPvv7tMJmHDfLfSRB88Lysv6VD1E3MA52R9kM88j60cIr5fXAn0hCtFtxpsjM
bB9/ewcAysrUlgofBQO0QkYPHe+Nq8yBd1XddnWiPl8Pglj+vxIqBjW0kLaq2OxhsgWqvp0XFB07
zIkRkE4PYINo98e9OWDdhts6uADEhssz/O2IFN/E1kymreaSdeMznR/RrXZmNdZgtuXt2W7/HRfy
zuGqxdsOTxk2HXnTUXIYhPzYqLHqzZi/vR3NQkc7wyhWBKyKC79MmVF/vpMYn6OcDpcPK/eFxsTe
WDgWKCiAXsR2vDi6xQ0hwgyjpQVhbtsRCcSIfM7Ys17whvTZk45MzVfuHnKdpPddejvvO+5btGi5
FcpJQp9jUs4rMHsGxhxo7uh0DfsXjfuuL7kucGNdNQYnswkidFLbv9jZ8jP14zCJqRbWkhsEuQ+g
ToHzYg7F8CxTu3WuN0y/dfcGKNr5vKXzybYrPKO71RtMOjv+pY5z/mwK/NGUX5A81hr+sEfhCARH
Dw+BZZydu/LRDSBA6M4GTyjQQqCgDcdi+Z9d7/8hFvZ9Z9+00Mp6tl5/puayZNBybi0ky5OujBLw
juLDJfyCEfNLAphuHT+Bbj6Ixv3JQdnYPa95zHLpCQNSRDwkyXL76H/k3rtXHPEBPl3ub7JRIV18
XyXxlRWelY7/bcK4UGh5tITv0kQMnKYFGd/AhiJ2dsi+mRq06PREwhPegYuXKaCnij6SoZU5IOSQ
C+2pbatKko0R2SW3J6cDYf0EbswHtQL0mqBoURS5Cf9zgsWedWVxDYm4Tu30sRV+Gf1eqPKkSSAm
/FH7WF+XiRJVfoT6x1o8ZWqx1f7P/06DDlWUoIRXrfP85vTqzVSDAzm9PCza891Wrui5INtDc7ZK
j3GSy2/vwG8306EaRnW3+qJtvYLuzJXVUGM+JKy9EEotmk+1L5k1CrKEmaiMYb1nnujRKsGny0YX
klYJ9xv2X9jy9X/x9xThYBYTJlV5J0DpDn+AKIg5+HVjWUtCtEAYApqg8kQHsuD9NcBXfPjtv50H
UiZ5ifdI/VNci4QYwrC1+nRukbHDpmdasTt39ICHcZLAR6bouWJzCKXHYaGJE2wvMopjPjAwZeVY
n0Yo7+PFv9jGxMcdZ+boGexE/81nkZqYTUukiOLgqIIf3daoeE4eueKm/65A1Fm427stcV2IKgTa
vm4KNkwlEdKrF6ELTml2ucXDYoW+A6EvcksfuLyCQUCNgpDU7IlA8LXXbY5h6h8Kw8SwJiqtWgbD
xq3PTZXIZBeucq+XBWIgK1nzSdyAflJcFyi8goZkAkaQKkfI5NM5w8DwhPXV6mQdbMw9zUR0dEkm
Y+oT6NxyVro2fuHJ20ajSp99wcWbPJ6G6lwnsjJ0AKTe+MOWQSOdBDoCEHc0IUWRYabYNgcIqtGn
TLqRat9KiHKA+4yYjB4B4RQ2D6LR+miJIew3DuKXPqABOSlUvRzI3v21syIeF9PkLkWCxkwvC7pE
/Uszi632gU1U+f5rr+g/gkpaqlG4LMjifQuW/0DIMKqfc84Dtj/OIs6oUBj/TBmARa57n5DCdWsm
nsjCmfE/vPrd5TghLJCq0knHHHOm40uogVqco4r1O5Lw8oi8L5b8gpfVwGIrYUo06C+a9uZfQK4s
Y4nrkoPeVO1jdF8mTzN4SJZxyVJ4wFMY0a+FB11Fb0L0TcOffaLxVVDtEhQe0VsYv7+iETYamIi8
Sr5VejigDDnImj58m+peIq7l6mZL5CVjwgGgwG6tmX/SXPiN96E48QQqQw5l6li3L02bGDU7x1EQ
94Y/2RSxkkO9WGVYlV+5HkEJBuuAD31pQfEsOgzt3sKkpZ4iBIzvlPH+NAL/+YBM43zL3tsdoQW/
l+L0y67l1Hm0DN5D99RUjSj+uUP8LbVdIzh32tvV2o1tc0RDJ/AG/61Gu1O68w8Ddyyp3ZfYdwRo
3FWHBCeP+9GSnV0dI9D/Sx0GYCY5FvILNayspxdaMqCMqaPwPmqatgfi0RE4yHr8mE0Vni79ngSu
+P6kAT7CnpOE4ESqgNa58iOtTRY+ED69XJdcfA9PCMuk8m4jRUBq0g6oyW03+jyJtV3az0VqEbbd
AOmLnHAXR+c/W2b8VRw+9W4KQ+qq+fzPKCDikpLi/gwwneCuTEv1Cv7aO3OURHak1bjVpdsyTrYV
0IXjM5DQIxPO/HUdrfc7qc2wEBq2d+ZeWhjalQPZXUU0K43hRD14ELQL3VtArmHLd5DNqNK+Z8gd
l7PZgM3Fuc2TEGaruNMuAwwqQ7vkQXrSon/aJqXPnZetCrApm8QsQZYA85Ge7jVjehxPzemUmlKE
VqZA0AzmSjw+8Gmzh8im9RNNw2F6k1OaK9KHotncKYfIuwhI5nmlOdSops2ABjVG4/EIuD9jTjWV
NkkpaaAta4X4kR7lMqEoBxfp+e4V8o1QBNNJJz2Sk1DrfoZQVd+V9RS8h+lIIAHdWKIPY0HazXYN
Mfox3qtuM2tFNwLz+wfG3SBeQhabTt4QbK4uVL6NjYaZLQ1DDyw924YgIXHlQQ3um8rxqG+6htGi
m2FJmVo0WDgnuqfcBqfbSYXp8K807aWQus+EOQJZNrH24D2Wsok2eU7INxcn8JVKBmEJaftSuHoo
1bd6WF0bwEaqGnFcTYc7iHPSrumdCiQ1FRJLw55eMIeLgh/Jpcy2PC5G58qxRZR6zWGwKpcMRN4Q
FLB9vMWOnLMX/P4dG9itrHopLOafqVSutBXz8LLc1fG0fjG0ThreNfh5qzg0UU0kgL6xCn5bC8wX
W3UtnLCfwgNb31/1q6e3xnGdM251NQNZjNNNKz066UswtEVUm7gSt2qWbfvnfP/8yA3OCcMt26PZ
XLy8SXGk0/kpAphVhdgHQwskofyHIWgc+eRy9eBuwP+sd0okDVrVBTQ+I1bqglE8VQA4JWh99qi5
DJS4ByUeRuMYC301EEZ4PrtuQJpvI367fy3Yefa4iyrT/hStjemTjxq8jS9YVlq6Omqea/u5W2xB
yAPMf0CpGBlXjqp8sB7RhytkIYc7HWt2lQ8um/w/76TdokZ2ONC/cn4n+eS2A3mi3pGZNz8DZEiX
LZkrQ9EhCkvsX1KNpx/J8mYYCj12jlVCzUGRbp1dW5Bi92EyrmXFf1v1b6o4d5TrY4WVfJDOSzQB
z4aVmWI2Z4Dth8uxaAq9tWJ33Uz33FDUT055+f5Se9slamdc+vwSPlJZI99jv2+Su7mlFczlO/5n
+3sjCNrRbgjjB7N5hqRE9bdQa31gm6dujZtcwtpJV5dLRfrJJftDry57HePjPJMuVUJH/7TOvsEB
+9PMFFzt4ZnyKbYouu04foCAG1dxKGLuzlnUFIP2UpU50R/TwhzKKz7WtGBtr2LneNICCSzdhGFS
kMqEzKkw6NE0aeHMl+O4G7XzArkbRRPb7FMFfTEXc5rp9vKHjGlwRtFrTfVZr1nuXbwd0F3WlSdl
/MbWz/JvRc1Z+xC7G+FGY3RIqrjJxwOR6MlzFkd/Fa+Pb0Y5FmJf65JwsBoX6aQe+B+uO6UqMphr
hHtaL1SJaDnGQBOoIKcF6JaU3V+UJvueeWHrNiXcwIpzOXcEXwf14WMoypz1O7UUdIgPvHFz7r1A
xK6KbARgjznLe0N5kWxZJ+TELUbo4lqOGWSt1ujN/yHaiTvcXCXntGdA627IpW2dW4uV0/TNHtKH
cwB+eSdIx3rj5GKBlMh4FXetIDY19pblGtOMdwGXJeGX8AZrq5J5Pl8SEJ2IzP+gVHTN+Tr2zI7p
QWR5TGmxAKJG/8gBHRMABnm446ncXDyD0HzKGoeUlxegWBiB/FOYmTDODhuIst+eEuKR+a5Bw4Mn
Wv4BpUZuuIeUH3/0gJIv9X0zGCIdDQWjn/ModTKSkYYzxwBp0OitSidAObelOSUBpmg2twcYaLvQ
IH+GlYTrXASMSO06OIM+X3ONd53DLnJWO+0USt9Sf3SKpeJrXNXCvmqDc06JYic94YNDKKlM8CE4
ZITcwrrlN8z+QFaqfC60X8gkhBSmZoitTTzYR2nO2ly5m9e3GGmmgAsmeRoKCxqPhb0cLt941mC7
9xXn0pVMiqLZgt9GUxUTVSYfamG0wATc2vXRq4Q62AbVww0wWb2bDMOriGDtSIF1jMe/kmjgcGTi
Az/CvfHJV4np4YDI5VzhWyGw6MZiyY/9gJUoSo5YAS/FJk/VCZch+L7PChxZ36NUMS7mJMmc0Yfq
UEPl1TkpcizeU16QlKP7kxcbqwrlXzcF9wlMojxNzH4yxsf6WRwGubbIGdAHTwmbKRIEUXviVrFd
wwgiTgLoIxMeOuD2N0zzgklhchqJsrH5I1S9tTf3DSWujNtmatPOgitfsvaR6JcTmYWxmlD9tIuy
DVWQ7ftnyTqVPwHLeVJAus5HkflcV2ACQ/U/hY9sUrKKUCzHtBlmgqAzKK5oGUDcuUchm7u4QDVI
jZ49s0TcxOuwVQKgtJ8ZZVh2bO+y0fxuuxLLe+6oGO1DKY/h+E+CqEQGAVy8F5m5D5/WMFj33MGq
mDWs7LsHQeU2Xf/kwfyDBEd7x80pQAPUDLf1jaxPV3UpVTKHJNZyu7HMzgbt64pMGNK6an9arAfJ
k5JXTGJyAN1ehZWVa5w/OwjNxq4lsbsp7H/ZpbQasv39zJ3NjO0QCYtj0RbQYou51nF5YG1k3GQa
H4US0wXXKmQuXUdbynldikDJKFkjx2Dk+MT8izjgYCWLiROWCFdvroeUcngiiK4p0Z9wdDctD5zh
icP6svgfaRFHK4sbNDPri0J6U2TWVtXLtnW4WLwMppdTpHhlj+Sl/WOA7Lu4PpsXr0q9QOGWG8iq
Acn3fOiVUUiCA7WUjpmk1yWoGZTTqg2+5mpEroQ6wG+/TWfvaM0pDWYytS6jFeqE5z4wt6DbBYfU
UoGXxRQiimoUKscpTTcZkbImidLNyvedsu9g6NBSVZKtSSrKaAzhCkdEuMKWzDavCCvoIwRp3YoW
zwjkGWQP0YQTZBMopO/MTbv4NbL5pyPgmzwsa4xU9rUnQD53cDn7rIY9jN4aOUQXLsWzgcrjkfuB
hHa0RRqdNxFrdh1pN/uP3FuKRH/dpqHRNNu5MNZIkawAnbCQP2W5dtn8+3wGvVjKotHAiNKi7KbR
NJNeIADPIPOO8u+Xt00M6uTZNYHJxKGL8XeNm1XkWlSOyRsiY3nHyJXIF/jZw4nUvWfpDx6sPqJc
2yaaxGSquCxy3ojAGMdQHHu0o66Q3lCXJPdkXodRTgdVa2GhLIxr1B49fIlRKbKCZn+MDLiHtOCC
2R7Nd5QoLYl9b8uCUSQK4kbgUbQ+L0PSS3OiSijT5JrSD0dlSVEvQwRt4F4Ut/LRHGFH0k+xGMd4
OIO2BSBv2GlFaW/2oaidsVIZYHNQmJFaylDb8XvKFhMoBSRTsDHa1yHJbL8QV64rV86/YtnAX+qn
yZCrlK5VHkusSMyyiaNMJqve75EYOGqqhf1aUaD0myfL72aCmYLQoPEQEwfUK69N9OtMvV2J3s5z
Cl7NtrNRwvWd1UQAf7fBND6oWjMYY2xN6yEFgyaPdP+icHpxM/q9nrAV6UJUAwr/2LBEFg8eVDmA
rr8rDXxU3ZPShvkxUX44TAVyQSttNnsmb+aqV2xqly2/HBb4nxIxgX8Iws39ap5lbl7Hg1GDTiXI
4rtVwWkLkCdGiMM8JxWg2H2Stz8acXqsRFyGtqUTkr4VSqgZgaUwSbBQ2yxr65/BRLyHRIGFIk8b
wuTxNInYAUNz5z6bh3sq3Y30VUwGBoAcvjN+fuJM2STJca2Vzaojv5T3VTcGzUIhDRsviAgi2NrB
gmTIkjFZw/zXe3obngJkFRhBt9sf+lGp5C4KOam7f/SpC+/Y/bLc3wn0Rb1EdLrAvzHaNKrFCI7U
iquxudAl7q6AKfrPB2Fcg10RoMDonUga8Vgc3cdFJbBa0uDzosOZKVCKmIjhiv+ogzcNNg1P8yon
UtEMTrYFIUOS/k4ZcLPjb+8Lj/cNIegW6s5mpOg3yynzAFNyv5dKLhNkU1oxCJ/jhU66KfDAtMq9
QODhhpcJhwlXiwY3BR1f2JEWRO5q6dgbaM9GZPTZyWlrUwYpkohqfHZKVbecjF7aFUaZU5tvt63V
H4jJBF4RwqcxMVjwl/NQXIDSNKrn+x3ASjDUKQpptkrrZekDDuwGVgvgc8FcefMKL5A1DKFNHht3
ubYVBAGA1yJilaMfKc0Z6xXx3JLaKkXdmJIsjj4mHzWuQqKGdQ6HEQROFOUcvRhdjVlvLiPq4PY/
jYEZKWkpC8XXe1pQWtKnCA3FOSyfXjAmVyDclRw3IBmagwKJ6MIv5aKDKiGcWVUC1OugnGSMnOVS
/njls3YC9HuQjpGfmfMg41RTFGCfVkUasYxOh8rVxKWbfJEFAo7xTOy8SwZLjaJB/ZyrRcHAtdPc
Dqxj0vI/WYPvDW4YwaADYZ/RNohKtrs8HxQRbeucLeYbF4Q8VuIw8kV9eypdUnbDUYUu6NlGO2Rs
mNSMlla7WcGIv+ruxxxAvnXqqHrM49nnWfIKP6v6CtGs1SpABdZmdbdzgAQ5+3NVqJGy5f/xafjj
36ieez0pya6Y7+wqw57x4+mnuLaI2C2qZjyQ2iQ8kYj/GI0ZKnv4rjTk4T+1lV2wV5kjmKHHBNAM
nF0R+xBWxRJ6IKySXUbwXjbdQXi+gkOBUFkmXnuhKlsaqC/xCBirU0c4OH/JrsJWCFVlM5df/BTk
FtaeJFJ2kEu/MXdZsQxGCVrhBRTNHnTniqVkwBilQ+dyd+66mfrxPmRIsru9Q7L0BC7oYMpMx8QK
GO8W/3GywNyUhJNYszguB4zRuRUQ4t6T8G8O2yWeraMy5Dc4tWycYseQsCZanSVvdoXzk/UPtiTT
gXU1Hg0k4EKKjZ3aMAZUsbmfj/BSTIwaTQj/vmQkdPUYIoGo+QPUwyamAYdiFS8mm00o+Q46vtZj
xz7yD6kYJcBlqzH9bbBfpTVIU8RD/RifoyKU9MWrPhxsTPxMxLg+gVqq78qmUWJGVKD3FdXakXXq
OzXjILlHyMLcHdif2IweuiwxtpPd2zB8scpn8eaKXloRtkm0sO+XszTjbF38f86h5bjYUIyX+DG2
3S8gbh7TrRIAd8xFTeEESOmyehoDKmTzsnff7g+MFQXXaAGlYykiHZz2n4r3TVlu8IOH0qBZ21nc
Quy6jAxl1VerX2me+P9aYOv5AdvW8rbFLkBOeFxmta/AnV6G2M3knCAAfdtYGD+qmZoRUxF/Vb9O
hw7JasIO96HYnwD2ar6DLJ3Eikd5kLzmRFcGvVqZqj0nJSMR25nqWyczyXa4i2PPVTNxk74DZIoX
I1CCFMkPXAQfH3uTlFxzEVwEONIkO8hAmh/6kADn9A69AF5WWiB2dzolLErZf0mjBDWp6pLgn7Ap
Y37A2c4fY/XTUhDgzpSdsMOONhrnJLg4NTS96Ch8OCJwmG8gbVQj+csaSKZjdddFZ3UTxkl7MTWj
CcG9awgDF1mIuchTS8iEGGlz9U93rL+9o9Yv+FojSCrUHGIlAcDTA3omOKeb4kqNv2VtXW1MRcu0
vVplfNIijaDpy42Zs/0ldESThhDjNtahNnNkAFsAyD6KbmlVyTUU3dOaqiR8Y5095pSDxJyBMnMK
u1uMH+GVk9wq1YeP/PxarRQebb2ykzP6G9ZQCUBIgPD45ElYY3muMMiRK+cAnMHo83H98/55XHks
UWJS9rg5T+kLxXeURcZjC3Jy1nCorvffxNAAVezokW1IYxUb/LD/YhUzkxYebLIT/gRAVok5PXmY
WqKo873QkldG8bHS0bN4XxbWBD+681bICOiqW3H3lhX5qH5CtaCcCCi6A6hHhMAkJ65YbbmPYIsg
1lhBfhfBub7KiduwrO3VkeUBFOUkD4aHRwtAhKoEuyhnZTTEkyGXAepo4Qbn8Ve4+dwO8r0xlQS3
vdB/CM+l+MtFoZRTYPZ3sWM9WT7ie1paIzx4qSIO7xKNNfqFbXkYguuftjnGUCO3k8lQAAzd0ajr
Q1HjM+HL25aWDaBDZHE5MnMVHOs+hq+el7tNt+KHaOYZkxPKOXaBMhbKt4fpF8xwJy6hSGM2VTMk
kN+5RSbmfRRxrIy96RgjqO7BQwUn4zBdznoPtiNL5ZMvvU+m67EJyshpzVz7UlPM+rpUBZ2dusfG
NQXUfjSNvd4isyM1ToEUHIIU4NeJDA4iVln5ENEHPOEX6kLCgn+sGyuLKavgmfR7u5/R3LmDbj7i
kDueKse91p1b3Nx2VDR63OER16srTQNdp5HG0//phPqruVcaJxAvSyyrdX7IVn38tGOoqBBe199M
dYEbL+z6mHemZlK4xtfRIihJWQQJbAH7HHNIQq5ekjofd5nXeI5QCe+f0j6h8Pj0Yi6llF4G3ZIg
6waW7lw7/eN6abdhWcsaFB4OxyLw5mg+V+yYr6hlJAUk0k+Ppm4fgH2rHv5vMuSRUJZMlW4g/EQg
3JZMx4HjdhfNI56TCk2QUAxCjIqi/pesYV2Qi4O1nRW4GuEF+wzlGFQRThToQTnjZnH8moz4963L
li/+O9YwOfWeZArJwPfoPAzIkw4NQimoMMkYiKkxCIdduUUUSe6lfaknJjy+gCDkUU1te7fThpGk
9uea//94r9ip2NdqjGtj9bWjF2sUntWfJMyYyfsYcvOtCVYdyv3P9zGgdVt0NzqIdyfDn5MxSgUS
XJIilYjzYULjqvJFjcF6B574MY9+2RsUgFruUQ6VNCphSBUbqPc9zdfy5tBRWdyM4TuwgXVBDctT
AJ5Jl9Udoqwj25OpFjm8UVFKLNsT34PkEC6be6uvUCfoT9JTYJESoB/M2rotDzs8hMF4g6O4Zmr0
A823CclNgPQCj817cGqx0rLTVn5Cb8Qrw/zFZ5cKAXkbXobbkOXAsNTa0iIi36Edowh8Fo3HF9iY
0pam963KrL90VD4XX0uKWU/r7XkHW0KN3Cl8K0l3FCLaqJqvFQlArziJvRQS7d2RjBCbXfSdGRTS
icwzW5WlfWeRY84+XE1UGf4glygF5Qwa6ssif5q+mdlzWLYYM48pO5r2tsQUOs+aF5za56ndnaak
a+RuaWwRuyHBME2Qg6HqW5gxNC4CypmNGeA083f0BPlQYXWPQNNvSU7Q9vQKhFNyqvX8Kp+MQSoj
Jh37v2MZRp6tSjeCd/NiNq2t6h0LUj2gQEyT8w+3ogmKO49BrsCBElQvExklQ6oUTshSssVNwKsg
CIj5Hl+3Gh9fhwKQ1S4nIpXvEd0d2wYUfiPsGgKxlH/GOlUq5tM3GwnFIAz2b3Bt65lg/hUYYnF2
DmgvOmxz+3U3JeoFiRY7xBrsAzh/JnYVyVaUlNagYbcAbAHEWgxTeUTxly229t5nk0m5zUXqtRFb
Du0K5bHa3gcezzfiHJdw4kvJn+fKDdPMRimlg74FuYxwBi3Y9z4STYRbL1WZN8Pv3wma8i5PaXYB
Nnqi6SYcaGYMh+tCMz41+MMjqBT9MqfD+OlWM/II03KWInHKfxLzrVO4/IWc1gSg8s5i9O8GDpar
OUXmLIQcPTt6AK0Ae/vMbAJHnIU8aCQLa7k9s0o9EnX5u4ohC4fgGVqwma6gq2v7fRvsZGc3QMba
Mra9SUQPfZmzTA6aSlMsaoVgcmVFhqKajPyW6aoqSCdgw512/UqSYv/1CmhwL9EeDUAHtOscMRL9
Fi7ZejTXQU2b4hFleA4OFSANN9aO1XQJkkLcZTIZHeGXiJ5kSMBSKZ2ONmiI6gU4mlwyqPCJx7/b
fNdL+Uu98FK8c78s+D1B5u68hWssKvzczagUD1pxkoBKR7dpjPHLue4W9VhQMBDK5LcxjxAytOrE
VSaiIZbylLtCzda+EG9gkzDVezKoeTnpUzCSxqbKLSzRR6NG7ZcmR/BBeTbw3kU3PhuboOJokEnC
fLxvUiWJeNTUF9ddjLMwtlQTXoPDVeVtOFN1aKK/JACCHZk54zkymLXk7JgAjsi8gR2AH+WQvCDv
voOPrhk8Qz+YxIcnr2AswfzHuHn+45wLPoHQZJHSEIhXjKRmoDuQgnEFycPazT+6ZdEmhBYlkhtk
skrYVL1UmwqnPh1rJ5cHeprE5l+NWOiuXfM/gao4GggWhw9O5j0mTwHPkRB+O77ZFcV2/w9AnVR1
SV8PjPUaGapUfUv+6+hXafq5Dwl+bzTmoG5776hZrOLPjS35Gb+K3QDwkk88x9LCLMwJ5XfGwWiv
HD7ATuomqkMp5oPMBziinjHo7nOut6YFtypWhgbKD3qPGPTsfZMWJVGhhnsyGbt9BlRi/tUBqcGe
Q20cTsvNF3l0T+DnwTBzcXiLO6+bpUoKZALCTfE2oUz6U7HB2GunUGje9LgbXMnFWsEifsSFmsCE
BXwGRWlwZGB4M9ofWqJjPN2gJiGM/4hZ317tedjhR4qz+0NOKG6DfPskIwWf9jLDHynyfUei46RP
TNo+V6irQxV7uHZWh38p+iplbfZsAyg2Fsyf/bLdHpScvSIeLuJvumwPRKf8iBtgORHF5+G/B9dQ
LN4wblj1fkFPms/GBCRXgCq6AAAZRbJJK18XL8klUZKTrS4QFAZiqMqIN5lkifmxWueYNw9A85/R
dE3J1R7YdrHBwv4upJ0HAuTHMfnhCSeR6gnPQaVWOl1lOll1f5p6atKNJ69RLXaf87gR5RZB9l/Q
CLLZ756cuEQMEFPg95QB9bOpftVphNogcuekhLIQiXL6Y2obfDby4Hxsx8iccCETuYbaAvNXnvLc
Q/YQSCIV0uUE1CVR56+nOa/lQMRRS6tDVpcpWgglvpazZ17Nf3ddJEnBbuKZC5scA4g7vkNiRIo3
eKzHs9vYM0mlXvS8Vd9F+R1Z99MjGqtVdW1+Org3/bUEaIr5sMkArWIYn7Sm3zFBzyzhQ87Lvwd6
zN1Xr5ABX5at4zZXvdyjj/pCSaEqDeBCXgntF8ctoI6aCdmeFPX1wly+xiOgf+vmneAet7wUbzN0
c2+skzp1Bx3QCYK88SlmoVwjaIZy46QPMvKHlMGtjJdqQrmrphiP+JMdRV/MJQ1/AqUp1qPgi27A
pq5YdYwC2bSwCxxxfLKYT271B9VtoieDP2CNC8ltSgkm7+e4noBivyEYy83y3xhnFKDCfubVz6qT
DMr0a1sljGrPLiRRGJxJvykqwMeRhQYTJJqNhbXPdxeMpe3rFAKNSuP9tjmHDh236/ib4Er4uwhE
CCq3bRc8qGDKr34uECWr6ijRpXzNygHNwQf2UAYD0HWzshHa8TPhzPD6QSdpFzqovKz91guOwvwq
Xepxv/vaUGkomXvrevS08cKq28Bn+VaaeinGm68vNrpzVz3mIQzeheepVefqy4I3URCl4zd9QsKr
Itnb+mZfo4ewANeyiYhUevuXcwhu5zIjZJGUYnjvrnUbRn4LV1VGD6JHPaA0m8U7Hz2X/q1lZzel
4rLLpMfI7LGvCVWDVV+TjEuSariWa92dKZ1NL/uKvcwyY3x+BA2uzJGS2+nacxNfowq6mjRs/Am9
lzXKtmpgIOewUNmAaJ6Wd1ZSmaTMVdutHuZ0wzZtDWb1QaFZGQg6Bk6JV52nKn67RkSkvlULac6l
N0BqVPBrr7tZZQFpHWwb3OwV7UFvXTLDZAKqPlN5fO+TKc6dFTRdH1ow6ZPLuyPcHCHAFxw1mefd
79YCvcBP+nfAar7DAF8N++Cq4MkYi4w6ykyIBnSYkCyQh877Um5KC99TrdXh5FC0xsZ2na0Ei73S
QjNHIHt4MzAlN9z+buqXqKKpiBS9ibw2nstHre26nh509yzWIqwp6Z8xNlaWRvCXuP1S2XGbkcnP
qAn2EMx5hH+KyuKuNv1ztvr/M/e4wZ6ctTwwmbCpeeT3cRCyqgr5ESJmdDN5togYy6HFla8tyUrC
hq9nv0mE96KnLGwFKlc4BJAkZCSXGlTNWRtK5qvNxrA4oloYSJOAzF7H98eml17B6WMerXWKj+OG
ndR1ghcoOSgyRiuyoOO0hF6omymOzoJ8f+7D9E38pRUlvG2xIhBu0M0/+HDsEdsWUke75O4/ORaq
ih4RTZyzLQrCw8UMkd900v3r36SggC8BDyb2xPSvRAuOGc5IlRX03ufX1KLEIajgxf3+x3NRGnSP
P4b61D0lP8v3E5vph33yy1IHoias6QE39X1MpMtC5R+2Ai1kh/M6VITslCq02b1T2u/mCi9ouho8
BMHEf/Dk5L3dG2Gq4Vfc2SmUoUFrlUb9zse61ta26T4zvKrxSt0qUm3PvRfFYiY+9oPTuh3ZT3HL
LJh0XVXU5UHE4bKkKkWGL6hby9Nar91WfaDNMt0WiCs4IVc9jkf85W2YRhDHUCtnK84CzvYzXam3
laxxXh13kwM5JwTM9RpmTB8K/TwMWO2EQnm50u20BFUv/8kdfpk/Fi9xOSpRBJFfRvSkZF3tX1jI
BJq1SurPExpnat14P8MLkYHwuaMSuEWq4jFQqKGT4qcWn89IhQh/Pkji6cm1uzoVoNYClejule2o
AchOLyyQc/aOne/3KwHcoemekx6H1MmIeegLIAdHKw8d1DhZbMF0yNZsHbMOV9dZ3lewLlZVjq6n
uwEsp6d7Cb02Z4fqJMMymyjqyTYD7O5kzOxTGy/0q4/tyi91/pDct1oVvQz6WCTgkVSbEdiRnKks
A2e4g3Uk63bG55VAgUXtIQlBDSk1hJChtKEXFQUeyRkbxqV30CaVzze80DXr576k80/tw+Pp3Xse
NZG3cu1Qp4K2+Qx936SayOiHfGw9N7JS9iNQV/PqMILILGnq0HVLu9yg+aEpaT2DyHeOlTy9mrCD
g0dsUiKTCw96Ux+IAojGDut92nZSMhEBS7GRBwGnEo1A8d5qy4BWYYBKjBqdvScwVNvbPdnzKSGx
b0wqXoTsw8SDR/J8l2/zuKVz4r0zCCRmFZUjdneMaVRSdurgzmeB8KXE4fGp1eHwXSqJ/CQM34VB
E31xe68dCFEW+J61+Amm6gHHrlJF+XQks3+PumnJkMqDM0b7sqM7TDTDbUw5q0d5CdOn+kh+pTku
YPSwpm19bbo0Z+MrZhIHTOYo3kV/qCqomR9PZQu14EXzW35A/rlVudzavfIr8iD9fbemi8Hk2/Zc
uhhaj80qpUUhp4yEWqfXJ/uQyylofLCX088BbygkcuUj8WVnwhOISOiuvjrsdmsPyE+HybfSwnOg
eFIVIfpMi0wU1pFj3/C5yjqV/q201S9Z1VMStDZaRS1QPXnbuPdCkYWoBm3G6pp9aCIepFN3i8gQ
tPDVmEsk86YY2TlmnuO0ruZqrDpXf6g6AKmLyUGrlQ8Dmi9rYnYQFXZSlAgg6nUus+R32VAENdsM
U+oT67EZFf0a+9kexrIrS/SZ3TAvLPcY9S5YaUai45NlO5qZuhrhv8FZIY49O6Xw8cBUa9TsA1p/
3f29jpSsNbz0Wva9rOSeVkok0IZbQVASPC68/4TE7V7djXrT3En8q5DY+TQzrYN+xAoVC1Muy1kR
ilSdV7WLL2/XjynU1KkZUu9kg1sHvEA5wnsWsBHRmtbiFDYdbIwHDBsIw8S85I2g0WX+kZDxPqm8
ljGmwkXIoGGTJcvLQAg2C7/PoAtNzDJOmxfmHmZIzO0/QQdUi6W8Cbk8QRYWBX8ZIJNeIY1Q6//L
eTggK/Y+w0ryYTWNYEmOYCyyvkmC2EyGmKWxJU95IMs7bexuOJgNi9svx9tP4wGPL0Fl46/QchXs
GXO5vJKPeCjbaYIUefQGJyeB7PL1Lpl+uI/tUgbEzKs9NNGjTYRjwSyCc2HjpTXC85qR0gSYxbKB
jTtTrgq/+VNJrx1bhpjFO71CwYz2srz9HBXuOQaxUjm783JKL7yeWpV74Zcw8zUyjGxvoFC7SjRk
sV8N/gfCyq+l+KM2SZmtruSZzun7V5N13AAd24flkpkjY6r6Za1gmG0pT8/izh3jRMPKst2T/F45
F1RnEEFwRm2MSehBTws5NqBtUgZdwN0/okCgDGFy1bEbiw6AjvtB6wv//SIKr0iWEgikmD4SrDhL
agOtPF5KCCVmW17USsMXnn9CSmVQChWhG4Jk0CAVGRxZrSr4SgwR608yFahSqmTXAABNnZiXDajo
SIwTyfZwTzJSF+f6EahF8fYov7Ehznpbo+iXIbZtPwCUfl4/mSqfgSEUFv5heA9nfUpKJuALn3x6
ArKB+TWVL7dSHIpIN/MvE7pOrBtSMkPDZoHcHzAOhGFYpSPilcQ6a5BStc0g4vRn1zyViAxmN72G
kK58erDFauSRSCDZlYWk8yJa3QI9el0ZfTNtnb1PsLH64FYKV7aRH9bJfZIyXKvv8shJkkjdVWtx
iyq1saWIcpyjYuZxs3OPQ1RExWUV8pLUYEKxUTAnUQOK1+q+dJYFt5aAlxHpFUYT7u9smZJZ+SM5
TBDmc1VX5bgp4n2kF8a43d3ZlQk1rNyYMWl5JyleNowwAO1MDXd/H+O2fjXMS+swgy2lgm6SQheq
ei+J2kKCZEhQqnfdcqtQiPqpR4/YurIxcWfAQ0GcfaPyaE5t8lRu1MqRdTgozZmqtS0uS+lWDf8u
t6oD87SC1X10I/JJPjMnq5DLawetwNMVC+qouNZlqKPCIuyMBdp2X7/QqdqEqedrYQNuJT8IisG8
guQmUfC+L3YIbjQYXvH9aaJzMRKqejQ2BiA3XFXv3KpVdWUgvL+MZxw6E7okg9hHQNvp5Ms3fyjt
aKfqbeVkpcYRTE4lO4lKcc/zgM8DRzpFOx1ibnhCV6gSqW1DHWTmKMpgkR1CTa7T8y6S1f+jBVKF
xMA7PLxJD63S6ilGVNjRU7wlRG4zyhypFIGzlkOLRGJEM/tDcAzCYXpw2ytfCH/QBwLM8Vdy9/Z9
HdDN7+ZJLaY6JmXRoLJd0uMxwi52UZXQ5rQCeOnk2+7CfoWRXU988ibv+RWXhAyePCUpZcSc3Pd9
wsIriUiuOQxWKySie8Y8cZvwb6Vv973Rjccwmvx+7Kgv6E0GSq3PWBwX/B2PQG3UEXPB3d0emjJ9
5LJFHA6ELRGaxg5fjx2/0iY8jKVoTAE7jda6im+IQFV5jF/l4y8CAm6jSd0sbkVTaFvGVAaY9KNl
xon64EsGG0/IlihR4F/N9c3tvL1gjmA9O0ujaiZ9j/0HLepuP+wduKlCWFRjhBiV3ofbVKKnU3bg
d935/2am0YKhRvRBDB63ih/EDKAK5oWY0PAe467YDwYETpG3PQ8wwaPdnlD7sgDtDeuowwVHjxA0
pSXurHFs9WciK2Ah5rJKmEL4Pflxq0kjXSUqb9Uui9QMO2ybhWnWWEGiR8Ioj9PSHLt/FtMe5/lS
Cu48r096tivAKnzYkn+4pS6qKQFY58agwLPEUFyDRKj/C3BeL2bbJncWfJpnYoAPoaXaqMEz8Jzy
NQ9ftPhcyS+O80whWIOEE1eC3MAF65iOb3/Ci/T/gUbuWuVTAaHiPec442QS405pIe+f381EhAdo
7jvbera4vEQ2bBM9c0Pa6oOsf4iDkdKmg6oVreol7klij99Xb6NnwfIBV8gSAVxnKCnSA7ZM+GGM
UiRVkNApKQ4pkOOnNNPCO7CuLjjOcUi5QSxsbbJETY45uBdeWAyuvnU65+nk35wd8gLv8q6kOJYX
/KvkBalyE3UALslid+UJPXXWkk9PKULZQvns41r3n3B0tYJ0GEFRSJuYNYdGphi1iiv/MxlSahJi
UF255JBzEV4sckdJnS9R6QNabjPI3JNfPeglE0deTKd3+TWuOoJp8ER0HqyWyFA9+43GmEHA3Ps9
R6ukfodH+AO1QR01rT17oJKzoq8JKF1TD9AUKKveQ3/7WbTtS42l3H7tM6UKAbSlXu9Xq0Z0ZurG
qXehoHHrOPb4oOrTVOx858hzeaL75DYwkRgRquT7GAKoCVpchv3XPRWFC9eOgX/Uoc9blOd1Tucj
B0pqH1Ux98aAUSt35H7hD2kc6U1cVtKY9kfpiiLya0nXRzb2fMx56YuQljwuD2Qp0IT9OZDd91ie
622oJwtuIx8qdCporM/mtzCAvLlXlhIxM9VveHVRm7VvfwBWwJu/CdriScY4PZmzJHDj5Kv2FZ/f
Ud7IYk3bDfSR97hXl/Gek3NDBix5iXWERFRSLy2B2j0TRcdJ9BJ7HE34DPlrBs0Xo8Pn9/Wkg7zh
0uzQvVIlgd00mVsQhkAJX+p3CK28uNilY5ihN8so+AqtP/S15c04dosXolynBx4qhDBIMBPK9CaY
RELEa31SKxUlikm6pn5udfgLFYDc+Ljl/eLdsDREC6tf1ZIkQGp3sFpKigKViWJCjquQDAUVCfMf
EQnFjt5k57O0/1KWz66+jxq7mwToMkOOm8eHdwYLFs/9OB1cwV+KOh0FFT1p7W14GFRF8YDhpepR
CzG2Q8QVp2V3i1o6j8UBoIAnddtscWtcCm/RyPgDIFKbTtHejAPD8rLxouOPYzZ1KsR1ZfOWQ2sV
t185R/K1xMRY/UbAdi74F2bE6JUnBo/20A9ziaqQqN0gPTPO4pyAdaU4dIxbstbl3t7PmqtwBciB
mVw7V2qn7Ge4De6evZQAxHSjfm8uLzefzVmMULpxGRDKYjiU4xdBEFncgxmhkNdVfNPc00BrxNFu
sNRO2B1UhxdJmUdzrVhbq/B/fRNYNBiCUvETq7GcHqYcTf8GM4Jxi5dBtl+ENsT75X36o6tSFTCI
Iv0nj5fEJrRBxOWxFK6LkYq/KQRTjMo9JdfIYDrNgYBM+l0n5aBHnGL1Ll6YZlEGP6ZEtrAgYVsF
Hsa4GVbBfxOn6ObDeymSEDpBNPeJq5JLZy/I3R+O2eJAyhIb+Fr8GtDddWUHGIrzBGnBvT+knhpM
vQKanOfc15+XezLkykDMwE7yuSpwVErYR0JNP2mEjTijJfSCpVfKiehpHeeybd4gidSfsSy8ocsN
h11eEJQ32KAMUpZAoRamMcbLlcxEjpsQpQUAwvXU3Tr8hK/o56ZqbFoYEEl8/2JMF1xDUs3OC4O/
r9/PUdpeD+gtBl5ZGjbDCn78CKXtHndJFX96+Xrttxk9DSehhR8wpoC0Io68lKgr3G8NkzBsQQjJ
RAQOnJX5Da614aTmVI9Mb5L1HuMg8kD2ZOekeaE68i/1vNMOkDD3FDnOv0SxwuoYcnt5N4ag1Dzs
172nT7hi1ieajl2Da+LcTMbpGVSVGv9BKIX9RIowtU3/YFIokl/FiCovD+kMgKVcrKBP8Lam9E/j
6dOOfbomHQyPbgaD95JhpfYuFqrSg3YCM+9xg6Khwi7gBbP/TdfRxX4/4N2yJ3TIbeEnzwHwFXFw
QM+B22a48UInhm2JP1H3ly4ny7PLYG5cjGYpjeE+Msw4k8JRTlUxBLUVoQT8vMpssB41gXgt0Rrd
6VFYOiQAxZ39UY2b9aphk5Ha63cNe1po5nwBK7MLSiNCGhPFoLbUQFsX4PorpCvsKvbwpQxLyl2B
/L6fvuLtOVlB92ZaKXbpDb2ROiqt1KCwuohNppOaGp9RjCDA5YAWJnWdE0VzTMfCTCXXBXLiwIjn
H75xEL53W+LEvhbuiEvOWfwZ6NwiaWiMSdIVZox4omYzlk/rtRBFadcQgJEcA10Jnckw5P5YYpsR
PYmkLwFaFu3GW26Tm8Pi8dZyGpvGmBB2yOd6BdRZPZYKv7dky1apb0EWO1b+alPigiyuTmYi2M8M
2+73XLawfTQAEvarT+7TD3M9bH1Zf+x3S/O2r36NcWsDFinvcOIZvXktVJTm5+wqNabM8d3uP8m7
0uvQYdr9wlgCtOhe6Q2gAxjfskbtQMWfFSl9rr0RrdNO5Pt2/Qqr78nRboM/Wy6/s+l8rgYnvIpQ
au4pB2UmrpGPkhKPywlck9U6wTANRyrL4ENgZ9Ca4GT6jF1S6PvJNf/Ax087ACwfHG5xDKY7pOIz
e9PqdUWsEnfxc7/GrTbRqDBR53r1AlF7qau8+ixSYt1GZxyLsA6av54ZuQgSXXveZ1IDQwVyq6eY
ahiq20bOcPHvOnLFVR45GKHEDpYtU2qud+DxUlYI+1mvay1aK3hBNkkDFBWRligog+1RDVfMtMlS
5xZ4/rxz6HRAoYPNL7SENEvDt1aEAWTLvCxO7cgHdivWFpwRKBI5Zo5MnTjMfUNpI7z2W/1kGkF+
01/eDaSIowG2KlI/OTy1i5uJDgQsvBie+OSyeJnsQuW3hWEJN+sYQFypE3LNZQ5iAycbe89d8C5C
9lVQTiRIb6xGy26Q5ILZQywjp2ETCmbO1w2mMZrxkmaICGMyaymza2zeIf/PBw5V3UzaGXhS/OkS
eSkq4lzr3qnBCGtLWnt7vttL3V3XMeEKtsryULARN210ODVyj9WMB9dhVFN2WTkoc5fTxsTrxJ8n
melsgaFbtzl1WoZedqA00h3zSRyO1Pv/M/Lp8aWvqIHx91+OXDQ6O6mEks8HwBxutYX4gx2XDCKn
0ISIEA577+a9HALC/V8TKWEzJYo/+L/ju9y4oDU2DKtQfby/YB48xkinXfCSu5njVr+R/m9vWPyX
rAhE2UYla3pTuJ6WM+OtTUITMEB1TtjsoXuorMJ9WJXusPeNDkJMwrgVwHM7IjRyVYtgo6aHtdun
Aah79QQ/O9YE8rdovfV7QQrXspy03sNBiTT6BthCQtBhARwE4zTzMZ/GHg2xOkg71oopNemgcH2p
b1NADzcpjorjRXC/y6OeUpIt7OlECnokB47uDSc/Axcf4vi19O2j9bD7lsS4RuSRaIOcioVy7vAI
8zj90eYNzucOX9D147uy58W/ONoM3dDriOBUL0MApK3/LdaE1uX6oWyI+ZYeAdVJYfKGno7Lub9l
CchaOx73ddx2ZBJQXCvsyTSrbTAevHseMLnlkeba2vpi4GbhbIAfVPMlnDMLJT/71oA+L3aG8U4s
8YL782ac4j3f8kg85mumwNDPaFb63XyaVH+M/hfMCIZWHVVTqjWjsAMJwj5YH6yCJB4TvMkgWSPJ
dpPZ+/YgxpLiWc+6LDbpXkc3t1gKrXwXahgEaA4Z2gY4tE4pyT5Uh/MzGRzhFEG50NfwqeCHsGK0
H/JvgTQGIfFla0GIbdBSFNCN4AG0rP3IQ6nOVEBqSpnvnsOIO7rqf0DpOhp0esfawgP4iDsyHUj1
0yy/lfAB2KYF+WhSt37DMpiKlXduk+ZxaTysqDAiHclkTFe+PfLOi6XCvm4j4QPuT+Qv85dJEJNp
nNwXjnWZxi6BUirVYZb4LWsbm4xlZ2DzOpMQznCSnDAi5OHvSAAvODzZzZ96+xRxcedz3zkz2vgd
jLW+3TfUu6KnW+9UupvZRHNJGQYH3ajtgLWed3oeFQyAX3dYoQeoOcZDpEmpJrqxYmsH5ofcMbX+
pXL2+Oq6MMmKZewmyWISZLluV8a5KOQSSlVdEbcpf0i0FniIeLoJrqUCuWfHyfd/C/XZIxlWFpI7
1A2pyCMxplISmN2nM5AX2m3OSdHtFBecGfwE/MN3F8rtGnwBozpw7OvmtrbhCu3J//62bPJbQ740
SjtTZc+qEbre320aAWWbnHJ5jDPhyYb1+qLUoNMjgeCHrXC33MX/L6SLmbMfLNcZDUJjborzg61g
eOEhpxQPov1OQGeQA3pgpINKQnUHIDkuWR5xBPDviE4LTHKbxRi9vgnST7aEElF/S1AZLiGxu+rS
F5mPf9OcwIFDZw/RRFZkH10bV+d4JutjK2o2qGcPnaXR/5y9grWda3YzuCDHUFZDSUI2mR5Uo7Du
FzEVMdvzGpFjP2ButMTIxjqQmS/9vQGQTWhQFu61BmBw0jPmRrG8ahnUD4SLgvA0NwlqAQbtifob
oRj0PvlV4HRjhFNQokZUG7jo9hCIVTVMdrAWRinWvu10XtAZ6Z2F+3VOLRmvlZADuJtBHJILSbwE
sFO66ArSKtGOzDtHi/rign1VEO+HTsH3d69aBlOWQbjAZzfyQG1j2TOEiCWfSJfyThqCDqrd2LQ1
+7RfkzM9i/UbNfSUvDnHEkFtCXT4MQiSItz6YjOTANpfVjLlzKj0OH+FUBVtWf67SLgzZ6alp3o8
TV05HVTGqR9R+kfv+DPcOyhh7Qy3V+HsDqvJU9GWLrZttVAJkLzzZlmp+ia2+7nfg6pzGDe2S+j5
3kZKiZr7OG4JBCHlS+Sg4/QZiu040WI8XO68B2s5emyiUd3JereQwpNtgVRKupPRr6yhBMxIk50Y
5Gd36ee3rCbc6IDj4cejQUUjemNYmwY+dVl8QM2xUaK96x2Zl2v1dDmiragrWDE2W4zhXQ8gaybR
wtQZo3aOpdQLdQ/pUQnzccvCqjHm7LjYiPyi/Rv2ozx+ns+09RQE/dDgEfSyhlHXb5UqKEKKhFAd
Hra6jSCEEmGqjJbMtQbQCgavWJgjOQ9C+B0+F2DXmhbw9it8g7jIiclUH79XQSEZSNzwEFlijEW0
uYLdzstJy44hKLhRo/9cz96UXc0N5TnExbXeC5T/u8J0i9wMuN52Px1EXwbufb9GYuKosQAQoDvf
6gyPOXlfxWI486R83UWNG0/QeBgf1FBIiDxNVamKZhCvYJCXkjXl8Kw07fH3qqtwNG0OUbgVK2+2
TY8ZBvvKc0Q/Eu5JRyoxBFlbUZxQfldjlvyffwd3m+xSkMc6JjdhwesMivAIpgxPYkjLWRZI6rMX
eODs64YwKCxpnEAmBdgSxSAyf5kwLqZTcFja4tm3IimeP1m05rjQIHa1u/nMQP5iZjCbPNBy4w+v
sIVeHj0X35aMzZHenAij8KnIsh3T1Pox760LNNDQ5Zpx9Jnj030Sca3uNgHtEWz1m8fpv0Nck0Ip
9KvR7o8O8SsQPkQpWWPK0qv8THPrZXBq4+sFmbA38RKLGqARcnVEQKujBIPENnJpESzplKp1v68x
+2h5ROF/OU0xSAqNkmvY7Fq7SBJ/Fe8k8lIdfpWUlNCSkS7Vx/LlLg503ONlmFsVqfbY9/onRRlT
IuCbvlU5L93iBC9nJBVcTNFXxBgOoB4jWOQZSP/rycb1rk8740EptEbZdvmrvCouw/HEtPnW1ce4
P2cpKWH7RteJTfobOiDz7vwrzaLItmiWJAFC3mdnQAwUMraRXyia2jvTBfpP6+YCIq1E8GB1Zik4
+AEImAPZyt/0RAozfYnGjWKQraT3K0dIgR7q1JmacqNzmrDOOquu1f7qjEwmifYv/gHjOqjb5nfh
XPeOzwPcW5xJy5P0pKja6drR4rppQ3jE8AA8grmSOOxt0XLakfZjdDCYOnBbTtf3baW0B0rFpGTt
h0vnaBGqWhbZUJoP59SHyCazrSXFztcbrKBFtuVWzT/DzZR5FnV/L4BasFQ6zFYWKgB4zdvj3FLt
2xvovUHkDztlIx7uTKVw6XfHcjCvTqwRSYD29Cc4U0M5Y3IgEs8lQq6jbZxnhBr7nU9sb262MejE
CIRwgjQpKNnHwCt/jgxm9uwOL14iIfbTBOUdAX7UfiJHt2NQUeHu81G0rOmDS8zrZcwArD8Knk63
NT2Toxcvmb/pBY5yogD58ldf720DLrRXGlE4IPz5bJ72i24lLqCrx3cVWW5oJDtyjSh/HtbLt42N
ic5wFpKYBFBXnaxg0aPmnsHTUytqFNpajWEVTnv5jmJNhwNGlFId59RXx9tcUWiNXX6/U2TjE8Wt
6G/UWZW8URqePuqkI3X6gn3g8x2m2p2MhUm5u1nkBroGqCB+zImZSj8ROEi6RS5eCYSbG5tkHeC5
q+sOY461pAAoaEGQMlPKweJuIEkHHqwmS1nMSGmeJEyjLl09GlBTfWJiaNtDqTMCftlBnDzFQLq9
j8GDF7oKWMW2+KbeFNtXaX5ic9gSmBujWYdOIMniQrs/iLJWLOUzUyFjhq2UDjFON0zZGVNYJivM
qDb8EG0mGYccjG67mImzHxG9smfvuLLh0sXNgCe73UBBg9jPy9boLs3oPFLtvGVm9dNEOwQ69P71
QVS+zxffEAe9wy5Qty3S5iJlcbKO3hUwWZUpNb8xT52BeGXmcik1HYZuLBjYXgIU2y0zq+oC95Jw
a3yEHr82HYs+IW1NeC213ZRrLp++wWGfXLsYiMcTU5yVfZb+sA4B/APe1PwN8QCV1dJqugz0MdH2
hNF/3yLHRLTOsUCxQhQtPJSqNPzm3GfHWEOiDK/iRofu7azw+lG9ExCvPjUXxYt8U9D3pUV2+g+0
wUPngb6qsADtDyEMg/fq19PUS4YubRZeCLBSGsTs9/hwLT42GJprLtDVDl77AgqEvUf10Sm7AT+M
0tDvLqOjuiM9aqFTtLeQiFSr3eX5EaePnw+hJ6CH2+sgYIJ3aq0LgaKEjd3C/+p+Mwn8g7EFwzEr
u8LwCrcduN4dDmoZpB/oQI00H5a+WnEEvcTe5oIG9NP4dBdZDlpwpxPCPPbLjUSziiGHB7wwxPnr
H0MaeGd2/ltKWxtDA7mPof68MQxN9ZhMox9traJ38gRr2xurAZtMat25K6dWEsVgc22PURksedIJ
v8LCZZZuNXDhr4gv99B4XxZIEswWcpKK4/jD8si/kzVM7zzBsx/rmmvXHetrzdy02+4PDLsVBJpE
QEd78BSWy8g3wRpmyqgff8a6hThHuN6bjfz+qFes80iww4vtDEFI1Jgy4+3wjS7z8hfgY0OBbjaO
znysOlst+nFz2asiHFJYJYsAt67WXx1FVDZXRkGSxtx+5m8nnsBh+3q814D6QfXEXOaasKTYZ+Du
ZJNQKNpr/Ss+WTduFoWhn23IRolENXLHWVHmkdzGJSGYzFnbBwG9gqfXMzSOOrSKwYB3fXcd3zrt
7sHXHyOu4ShJWZyowk1vdY783UjlGw9Mvr0QdwaXC1H17UrDT4Jw4DoXLhrInPT32jxkgpi/pkoB
pu/Ba7wV+sVzws7GhEAAYaIrjUVhY9AX9gMXXiK+utgTRoMBI62j8gHSxSsjRsW1VFl3J0oKAeJ4
hHlenzT+pOEQZWPs34sBFiPD0xMVmWVbkAzkG4Sxf29ay58vM+NiMk6EjSVf1a0aOf6uJviOtmlR
5wf55+GAa5ko5ZwmgEfv2xWSIzxsP5ajY15KNFNx0uOpZaFa/QXPggHauH395FRFAt7nkLyrWDZ9
OOAASKN50dACA2AmWx1nPnjWubcoopkiBA4u+obge+yHUqlLoWe1foXwKDjSX5S3AmXfTRLLIWw2
WuTlx2HhKd6SBFdenTcB9MGFQdWeGBHPUafHDDJh4edLVtQR3k5aF0MOITvMHF/bUZxyvtmWcZWi
R8iiNOvCP9K3T/CTdk8ICr7csh3SHpF5rRh6t/0zFUjgL6rFHInEjdN7WFgGq8EsjT/floGSGR0W
qZBOGZgbS78vs8l7F/XUSGXMc61/8xTPAmu8PGXF78PVfYLNgvg9YuuUI5KyEvzJqoXefC4RFylU
iJXmo/ljY926dLrarrfP+DlczUTG80V7ouUYyLYfw0QWEEYAkL86xYb+3/uCQu6WmztZLSfdLuYB
SmQ2F7xtDhRipD25ezy70AsV/M06YTT7T1OS3AmZb2scLUAHmllujyJE8fmOukbI1jaR6Lfnu1OK
BHfg2F4zvqr2a+9vbpCeGh2L+iqI7Nwi1u6Uc7J4gAScWKl67fl8orzmFINodbOBMuVzvZ5x8fIW
OIojBJZX7PebEU1z3O1+NmH+L0qs6JRJwKtKlWtoyh0newpXqxYwc0lRfU9NrjRKnsDuk5x8nfW+
h8eOQI0J80Y2OZMSf3EGVsA2Mc5cxpde9lSEBIsrAeKqeQWZP+oCfh4OcYFi/WHwxqiS8RpSZLPH
PpYr+60uBs3B4MMH3kJhQa5xIcLjFMSESljEzhPv2UOVf+5Db1PB3Lq1LTPOoy1e+dRoqujGmPJ0
FTAWiqng1iyULe6xTN3p3qwsZLwttiUcFOFyyYHxFnRZKQpe/1HzI7v7i/XrhsUYk8qn7O7K8RBl
Kcmy5nFUySuWu8KXf5Ck5fkJWpIjCbqS/toMBtczWkHQ636xBDp7e/wcGdDpcoCpMC8WAnsGWOzF
1E1PgD7V56wuFRGYfi27Zx/IvnZmjEWo8+x7ij+l+VU9Kpip/Rbn2zwHOKRYjnoiBLHwYZjAia8B
wI0F2RbStXLyZ2LENMyL6hf6e/QiZH67ZbQeOOL4G1aO7BC6QYsWqCssps2ygp1E9W0gVqqO37Kh
hKpvQwCeXDNa5T64bpLBb/eooLjlc3gNjpwCVzBCFi/X5oVUwPP6TESLJclseEN92Z0Egb43LJdm
geODZ2Jf6b8s/3bEhTLtkcYLYqamfsF6rCyjvum5xy8kQ4Za3GKdI/ym01wNl3Sgp6UvAlMBIAs6
37bLoS4GHtjtkh2qstY3yM32jpxor+UFTMVjIotUDknPn6XTRiTbHv0lTTtGAFay4Qcm6DHcPton
ZAvmPCe+cFr35Q0RqsswozOsbt3MtECt6Wu3R5+TW4jGJYJOyUjOQM7fyMSgVM77QyowJA4nVzlR
OO2GqKPD/uJ34xt/ZapNsjzJ+Z4cGVc02sCv0iI6rrP/1E4fKK7VVhk9vQ9oq7cT6O/s62googlW
cFrWYz24Smh0EvQhyxolGN9KKnGRMhXA8antrlrVqfAtnhjDKkiaL6mHIPC2d5ki7heP3IV6WKjQ
jl+a4qVb/4j9NTWiUNEvfWxbxaogPrEdbEUSb1W7hovQpvXNCJxfB3tR6L0RgdrBerNSffKtv9Mh
ffks5+ABlKKTxwzBn+0N72MWZoabvPheg0TwnDbLOy76bOMGBQ+/MMVKqZR7zfkohR8lNEAKnSbJ
wacPdmm+Tna0Mo/NWmkdKfnVZg7PNeH+a4NtDv/7q+bx+HT6Jpi+ZelwNATlkC3EW2d2uMrJNXua
OGWQ9pBieS9V2pPZqn/Idey8ovreiS5PbRfnYGCJL65sGdJaFce/hgLSiWv37VMjdheQokUdq2DO
SGXJ1n7TP8Zi/K/ulX9HqECfbpxmG1P1C3Deqgsaqym9iIaHFpkYR8P1Z4YQjFEE+7RrtaiTm0HV
MdPpkHHEctmPOUhNlQNJRq/v5WCj9TOLB/a6jwCYnuzB0tFXsr4EL3Xb3ZalVFcGaTG7wLBo/yTX
XQZZwbXqnDN4roDynu4d0UwLsEx03asqv9sWuTuj8tRChDISJz/08nXVc7w7GucIlVTWiDCenAfm
wVVMpTg1DSPLNFIOFMGqRxTdBy2snVqvdAviFkIkGsODjIavK3i+0DgTUe5MEsiWt5/kbpc4AyfM
dTVg+iBUc3MR8b6tiwibFmRWWi5lQF/nroMjplG10Jko4Wy7oVjgwc4642ml9yj/Jk0rbRDGu4zx
zVdYEorTVhpv7yFJjpW2y+e4mIn6N/vFIG8aYN5AF8i5Y3lMMmi/GbL9VMLVIz8voGCWOA1m+9OM
Y6iN/5WkR59oZuS4P21D/nP2GL35ucQGHSFBC6D7FsI6VeXyQTGnieacU70gF8d5mVCCnrXTq5Fb
ROuzKpOUcOq5it+K7p17v2huecvtfLZk371EFQcsG1r1ljhKThTG8e29+vlsF7GxTAZG52l2zc4F
8mNGvCXwLRNBu/8bp67zZgj82KUtw0lO+cuioTKO+Y320uKJeiUyum1UELjtrt2sI+wYZuPTly8a
Mlr/OMSBqekqQKbl/sYLDb00YWDRXZxHIda8U9D/h5W+vF/jtsNG+RM2WCcJ0oSZ0YAeFJWT6OAB
LyCSvd55BBIBxkhmebAzGze8IsGrexf+2A6waRRv7Me3QPe/IB8R6jAqZnwvgzXkVoEGl4UAgpij
14GH4ePdZiveXthnY6MEbYueqJqOy39VjEQXFcrEVnwHUtoXg3AHoLuAkdbd3KGCF+4pf7k/pX3p
EJLkm2Buyqkp9k14rc0Y9UR0FzL0IbO4AMEenFvIBSuXWjgbVUg4MVGjDna3MMJS4HE5cuESLIJC
Amst4i+uvj4hJSEejj2n2g37zpyYo11HshRysOOK+dogb2y8hmymeF+4ybGx/3Y35dxL/bshOZ4F
fyPsKNJWd5UnV0vN32881BErKLoK+ro3qpL/hQbwvnHr3zD3m+HujFTzsxnPrG3xFX31uuP5ZajR
zeNmTRelyyyW8CZW6gpAXuzw9iif7EIVlVkSfwvYRouxT8E596uKftqlzj4LvDLY8p3QuLLg83wz
cSIwbgin6BXYVUYfbAaUxAE0dp287vCAepkDTAndNh/RH8OOSLaRMhu7yeouEd55zFogDWlOG2nW
F7/pGldwt7DFZ5oHg3IVJ4+HjNouerTS5unn+RU6GcTNLBXUnpmrd049tURjdG0aeu9IliKJBIxy
hnfzIxa0Qp51XvbPS6RLzADpTVQCF+0OZuW3uH0+tgW6dtzviUAFu75ePlwQPe3Xxx4dqp+72fr1
ABidyP1raKRWE3d8nt8Us5thy0m7Nk7Zt8bNxxN0EmSCRwevxP8z9dwhX1hQzTvB0Wo2UbaWWNBl
A/qVUBzzSvsm/BWX6dL0WyvsWcDH1Pu3kRzrEC2NeyJ9hKShF+OZ+ad71QXH1itNMHH3Z7693kx9
NnD2CZEBCoLBf68kMPDqssleT6AGNuTCGHurQWrTfQKUonksC30naH7be5u+tfKwldyCk5qIJnWj
LZv5eYbkCywLbLiLR/ufa+cCOO3cZVrB1yhAENMjTwtis7cXgWIg7nr2G8oCTj+TWQuE/sNtUgR1
pMIfr1WPiNIqQxFzZd+ootZd0wSfMWpGLibZmjj1Zpgwmhdo3O+StPpfuj2VYOkSZ2K9dpED/ppt
eI/clkfsWhbNGNHdCitdt5uSlLCfotkhpy8c9PD1I7dSzVVmkW/Q2D3AZGYTYbCNsGcZlrCFv8cI
7kLIEx6EziyP9hkX7bV0v3X/9SNaN09Aa+qQAi6/6XkYZ+uk8JNiC7CQ4vVAi5LlGobr2naySaM/
GxYRa3tqvlB1RHlqwVht3N9Vv6UIXJ/WcSzVeopGdxsYnC9UAejzQxMsOTA0VEa1e2b/aTsW2AJI
6O0D6yzLDMg/ADOQwht8dNUBchGNOh0fpXmRzxXxfaJLDRd3q4/8Tlg/qaF4+ShYxYhGbPIwBH5N
/gVhZYG3/cMOnb+pPoo5yWKT+624sduyP6LYhRdgqHrlXrWglWuuJKr+Sd61NP2LcOvPOkBnWsa6
8u43wmr9hRaa96S+wczeG2ZeHwBmzeLuB/RJwj+EMa1d5D9SmCagbk9IOZUL95cf1zyQElnvKu4z
oe5+MVl0dfF5QMv9FMMjS/K1uE46IhVTbDp1UOsoWTfpqkMGIVx2Nob49ff/K6jx5TxUv4O7zvxz
2JBXRtBrIqzYhmC9RmVUkUe1u1IQl6/6ZH3V6iMCFs+gi847p13TmxlbmT1cVAK7IdiJAxi6rkYz
ZLO9I/DdqSv2s8T9Wa2xMnkie/8jVLcy9Hv7hz5ZI0Cjk5sqyH1heg04BWJy1ZRMsNt2JSVyt85R
mh4iPkBPWum8pQkBq9KhO0Tjl4O1dB9M7wWiPjGS3X396tnl7JwSSORmUWL6NhNssQXMVkWVxPmT
6FiwIpI7q+QkxbQ7JGiB7RaRYNM6nuMBvpkkAKyOrixL4LcKNBKyJjwnOxqb6cI7yEBd62Nut8KI
UzjmhcTBI3NoQYsCCv/tZt3hnU89Kf3lWUphVYd1UlK1BjliCde/UeKhnSM2m9GHXF1vq4mf1inB
MR3dzRCqM5Kelg/VHwIEEvXMCyPktG2n2uHhBnHYD1Cz3VabOs4ooSGbHRpPUu9HmKXWT8P/VLqN
DrEgYF3wpRHdYFOlboS2uiIychmHY/W2Gwxsk0LeN614WvX4tHcF0DiPM8XpGTuFXt9JP7fe95ld
C0d1PeJY9P9AAvBO8ykb5ilijEWUYp6AY3GQSRaj4jmfV58xdt2rL+HLHMgiuaB12FEcAGZomld/
e8tPAFOyALpp0jLdlLGm1xfxfPeWRjZ+eJSvnljs5oBIlPLgq0XJU7CNh3wEZNKbX26Z7Ky1NKRX
6nUscT9i5nFCcuMqwR9fcpNVX3O+CTLCWOE+xczmdaaaLnSWHuzXUK2kHoUnNe4cMp24YiY3jg2C
T99fTsF90TnIG5k49ZhQolYxXh73qhIRvQ4446p0pYeqYu7coRIkUIl7310EjXo6Z/gzwCZCbM8H
PQdIgUa0kuBPZx3wCl+d9BzoX6/r68uURYj8oQclWzjr8qh0No9JsU21FOJqiqBNfYKZ6A4drRYE
lEsJ1WI1qoF6o/hAqR3rxqsJPjSfIcONpeNnV5zdFPQHKq9rbj3C+7OUPX4kfVF9ywB+vrGqHCRp
WoQ5DkSYgKvFIH2wVV2ZFTJxf9I3TW0YU01B0aTiXOezaNLYFS980Eh4r6K1dstVO5z1m9SFnO/h
GZnhUX/qkOMU1Ps2bv5a1CsLMcCTeBycy51fdlVljRhFO/Cm4xLfEo9s4IeLTPh+BrSU7HAY94YC
ZUoQN5vuH7GdjrzqeUAXJCqWI1miU2bhuMcaDWZ+XKV4Xe4lyO9NF3sT7mOmRheXAzQpt6laG6jj
9wVW/FUZJKHcg9z/Bm9t9Bk98yUwk/azHCtUgU2insahdERpnL5awuMF0pMd6eb3uXWtPaxTt0Nq
M+U/chDVtpro9hsfKVk61GDJC3cXALYc02c4GMBwb1PAQy1xuxR3C5oF6lDBiIuCdwzXpOP2DbBx
PKwC0mzGrPPMNo8/wb3r2lbvyso4BLUeSXJjQ4nfzm+4NLKkjgAu76bZO2qm8ApFekF1yQswEDEO
zN4hrCGkNAw9SfYHzNewpHmNAcqy5UvbVIPw+IcLIzXPg/fjMoQyU9XlaHg6XNEoWUHcsIEJ3AQu
IKGK+JHr7NQqLl7hy6iBs1XrccG+eFBwwya39/5pDTtFmpa0/Mz6PlKveungrJvNzxCurnJKcJRT
DlEmA8uvagSKUYsLK2AShImLpkr2iIF04Vfq0KAVF01RlmzlJBcMVslgoCppwm0Gr2BkL6JT82mM
mhfcJOSnULA6FBs22g53xPaB2LQsBqSdabEpJiGwqjRsovxQ6rVBmt9R01EsWmnPguXh8n8lMfXS
mbjNofQzkVeWglx2f4I87fG7PAQEZyNm5HFmiY01v05sCTYzXUyhPBKMrGXgkzPulaAJaFuf879M
6VXFIKUA7KT09nMEdHZ4b5gh3eaC1XTBCjoRYzcPVDhhxf0vMWsJtZ/xqfR35M37XED9K00YxfRh
6Rmq8xmsRN4EUeDlAk7ZTSqXBhViM2nzXPNS0owWHWuC5v7dkisCFYlkFtukFhjEt0V3ylafq1ld
Ni+rdUOQT/fXf2+zH8vZGtS2wDKbjrysfNy0jOf32YVP8MynO1E/QjAIi9KZPGKgXFHSWOtjh2Rb
HmbhE7TtKPZxFZf6LX+f7eOllsXiwdjLpVd3OzYMeR+4ccp5t24Y57Tky0Yb9VfZsBwPsEqmG6oJ
HCUIgQOtd8wHjWNMisDHerAA2fbJuRJaGzBvikG6y6XWwRMiSr4Xr63+/Y/0SBGFWjwMyd0uSad4
UU7HCzkvU8KeSE6S1mYoqT+LDsmULyhFuO0GAuGh4OpsP5MmLk0CMa9nqD+4ittgSqZJykxSSzgM
0jo4mO0gF2ePKZnDC9OnMXQXkQ3VZBkzm9BVK4ssUlEIu7AEtE7Y9RqvHk8ay4GcC4Ag85tB5Meu
EztLW3la7gCgped7CsLWrID7rUwsVATl3fp3OZscIi2OPV/w2xFXHHinG4L8jav9eX2yTXaeNJz/
5MZ5xAXOzExaY+e72BugvHr6q4eo69NXOwyNRmuwsMzQRe1Ym/Nu+Di7Nhk5jaRZ14DeAf4TBHLM
Ltnqoqy9NlnrZbiCydwH5Ap7JpVjbLlMyCpXlGfMEw9/ts0V/lSMi69EY/igwdGVvRaoL9bEK8g0
+vu7L4Vlgc3+Is7W7x8Mp7Q975Z94C2sg5cN1zD/nmeP6Z9g9kpLO3JE10Jfl37XK26HUUy3ldd8
DLfxyM+2PHHklwpWXJhvIjeOL7yJQD82inchbXDnNbylg68iJ/WRygKiY8rc819NYpGVBh0Do1kF
pUOdGaxaAk1ZeLyrN7pxlymVY0gv3gETV+D13s6CqQONL6HoV1cXPfOjadOaQ1iO0vxEQrGjW1x+
b0go/H7DBRlS07A7grzSuvqtx0hd9LXGVSLmbk2+4kEGpyA/IGGAf1kYWXug5/8RAcgwJJm5e7hL
mFiR0JgkvhvZkMS0GUWtpLoihybzDktYLc1lEmWRIS0MVTD74YBuvTqdkSG+sQqn1SEaQn/DBQtb
2ilwQyNIvrsSjl4UFow/S0iwx00LdzZG9edUOOh1/qMHEHZNk4QLlQAik2lvdpJjHNHWgdHA7oFV
dBlfUPIXzZRik11HklHzOthGXwRZWfmHLJH1cANOJOyvwzqW3nCsCPJyuhxwa6R+zh155LPht+sK
peMLb/FVACcpSkugG0JGa+x/fe3hPx+0+uYK+Mwhbhmo954Z0sLoqMzUGGhCtZfTttrG6Wq0NkIX
JQhwuxaTgKkAB3XJZ0bYYE07xtWY7aYABuHpZPZWRpgBn9xFIB6yb6gSyBaaTdgk18litWlIKK/x
jDqbfD4uHdSACX4MZoCq6ZKv61GrL9lPyr+9iuwh+WFZ306Xh5uzDDiD/jVPKnR9JWLD2PVptWCy
h246toxjlRfuhhDqqRb8o46haKKuqjLVYKDPogNTFZIiQ8zu21vBmrNef7A8ZQmOFa2JWOU0WLUu
dgvQnHakU1duHBgIY7RTKPuS3oLxBWFJzX239KYS5uhhoshtbG7CMmEh1BBMoCQE2mpYzO6Llvgl
QltpCu+f0/ci0IuckCzbU0XFp/GCS+TxKOhQMFnf9MfvHBMzAloQnqaF6gW2B8kqkfxEDTkiGe/7
Bq5Vet2IrRuv7GUnhkf1JXspJLJhG6GOE/mx40ByllzWO3kqcgeWS63jiGQyItWrTM3qfqsH0q6M
vubnlLscqccz9/rKybuSxSZNsbFkX2EA3Hr3A3TvFmi9n2BQWMIsLh6eRvweLCxdIH4c+dClqQwb
OKKs1tgd6lXEK3XsbBDKrG4hGQShW/IAW7lrhzNHQm+47NBhp/TnnafNqkPy1Nk8D7fEvP45UJbw
RMojWwd9qvQN3fFyGVVDKCcBZx9HxKftcCWCXWCb8jYtCgVpN37jJGH26r4FmudbhgYMA3WR8ahD
ppfoKa/rT+gi5jyDf2eBCQ+xL5DchDqatN0nY5Q506RL9tIx1ry91Acm8N1cxar7tDdxcUQUv8Mu
vLq+1K8KwjI2hYbMSkFZfDkRxEbDDFZQa3WE+TC15ZAx72qp4PdhOqBUdRuJqKbmO9StOc5OvFaK
e2TCxpebEzUVBsjsybNgz9Ir+9COEA1CeeXVVeiLC0ky+I11wut3/ZoAwHehilXi/WMWgGVyEtVB
lpWce4qHguqJ/elIEaEpm358pPG6Q2yzD9EZevbOcIClnsn0XeceZN+n0Htngf0JWk39EMSm+UWh
v0MGm+cDe0zBcJSB2lMHRtr0VM9rMg7/VJdjwj37WVtG0fE5dW0oOQp1EJI4LthSob5evu9XdClh
WZaOtNT2JdQYB9nw3W6n9GQmgWWqMLQgFcobPgrIIUwttIbmOz7jWhwN3ZOJ8yOZ6Bj/xauJr/F0
UEFQhMipJNZZP2IjG4OB85+9C49cEde+AwKPfWI6lI1ZJKpM2K7Mn+At4aJrx6UOR1sFik4ccfTt
CTp4x5moKwUDWY2pWFlGgL8JxlskV2EvDLlZD708pTDqs8ofLD0o58nEkRmnoqmHl9Wb0WaY6QBI
ybYT9dLTH8K6cwt0icCgDj2zw/8Hmx8vw4ZmzenS/a5R9NW8VNe4dYybcI03BiaZPtR3Own4LqXh
8mYx8WSMZAJqII4dgOp88+SigsNIuCFNf8AAT5EgwF0dgw8zI4m5PAB3D5G83Txz3fGlEk7CN+Vn
3QPoAq4GSp+RJS1gqfhJOmtiwkuct+WQg9Dm/0VAj6rNbgpr8pD1b3IkxeHmB/yU1ooIJB9i9C5K
GT1qhDiYQVkhIIfC0/GP/RzbwPCmLSbeeWHtgaYHVIxtNfFh1TpEP1Tqj6o5PrTlM8+erziuDwnO
Mw+7Sd9ixBFhP66ClEokEhjOxTa5uwR75SAU4SeUIKfguHdoTWlbNnhVjoovSTRbkLIECAHMHXrL
0jVQgSqyrSGQtb7EaZWutwqj+vnUhv3FcYdg1GOyXkEQXaK4GAqH6wifMI4+ol2NRNeXb4rXoefo
1Kic/2Zh+uIZffITRkxsePfKH77kVbHdrkwSiM172btPx9FEJD+qcKjcKPlYbcJHNyJltx6jgZQe
2WBJCWiC6tDxNbNcYxzv/NCD7/rKc9hyjm1RTfixFyk02nx9wXboo7Gr1EGo6r4eebQDA0+uOtBR
WPza3qsd1bLssRz8jtl8FU/Ob1cnW5YMXzZdIeL4Sz+VFXUoFZ60Eb9Z+puwga6Yf7HEpD3rvXOH
Vo/esIH7mKp0H052k5GlQwiB4Gjm88exrMZyli4sAMjSB5Vi1yk40/ANoyMIt7cqAulEx1FopyNu
Ezv0sq7qa1lTdebfmlncUoRulI9s+CxHQySrIhObmvcb9le70+eRY/3wf3m2y6WHrkkEU2aWUorA
s5oSuH3TlQ5eZNSH0Cph5iQoIImT1w5tWQWSY9EWxuRPmmq0Au0Td27XdvlTUQ3d77bWMRLgH8l5
HM/UCa9ITPKSZ1zAUjnwsJjnsDhA5iOzHQMo2stBA0i/Iw1Zf/Lt9ZkLe/PK1VhR+Wi+sqAUpr3F
QMrS5g1GlKFUVTAo5cf6++O/07pEMBFHohHa+yC4FCSxFeOdEWQm7NWYlxDNAUJwGVr0agAdP1WL
jxQxzcpuAEnAjlVUqinMDarargc903BDFIIymIhNObHTqc22PwYl0w4xeUq93MRfztwM4Zz8ZEv2
VWTSe5tuB4OOCwcanyTl6M3FLCpmnupxqsikzjPfgie8m9KXg8AMpXOdvRTs6fgqN/FybOr3735b
cu64PSk81a9A3OnSH/ny8oTrmUJaV0pcENtw2zIaucGMVxTkHJnwbu9DIFGDPJv+MiLd3QrVM6dA
z6VoUWD8RVl1hu5DHxafTRkKhyQcXor/84wKYTA1Two32D9OjoKRzYguPOhfLGozTeEk+SpCItQ4
Yu2SpjmIBYcYdPVPoKjO1gOwMZGNBzk+mzjyrCufyRvxFIqJre6YjAuoEcTv14CeU1oY8dvSjBeF
jsujDRxq5s5Wc6iEF6/i5AMBR2nmNXrb3omliIrlOP/9YbmQ3fnN4HM7UoVxClueAouvLuwNRCVa
tJlyLGr6JAez88xc3uPNGjcscrdGsYOgWzhRg7rrtrDP4Ugu9Q44R59R2K0EU6g6ANdprnheOH3W
DerPX6FQ73ZcBnsEFyRugRDPXv/RThqvtjBrXY6/4Pmk+v/ClsdWRI3tLJCFhyWFFmmJd3wURr1W
c6ajp78JOqEb2cyTNORSpfFWJfdqpo4BM8XjAAB9yWGg8AjqxofcVrtJw/V4DRZJ5JLuSNc5lhzI
Pro1vZjkMmtpYDZxsdLHv+ei6zT56FiWjYzFCcL86Qwy52HVxw6kZz9qOrnvHVED6AArZvZNFGNv
nQPq1dzNJLUY0AtUal1cc+P4kKME61CYf2Pyi9xFLQMmfZeICFAHXGvQZNtw1MgAUZdDWLWwZiu5
xKSdzWrvyCV9zP/XG+X3lDTJ5CtxHweea13lhCCAXJxkyvfBrL4qf93CpKmGr5FmnjIWyaM+ew97
/zRtpCI8y3yueh2aJ20viuvV8XnnCHjEw1HNTqDzYc1iFq5HcOf1uIc9LQp1nVkMo9amA7NfUPc6
KcCSUZ/D8C9Ezo8zuNGTjc9KeSuHWrrJtc1FVXccgL6iG9Tn09uaI9KJdFi34LXoFOwU7y7qEbnV
grRfypW2xaTYTiZnSPS1fzIdwZpwwvYpRIJXx+nHLloayW5C2IPaH8sVEbafjvPdk5X3ci4I7TT2
SHlVWhfL9Xnm0zb/rBcqmmG42wauUGR6miZiar4nu0WvWSLZDGC5xDXwNcfxBEI8QDhfSmnXR14q
I/pRg3eUvjwV6wAXrTRHAT/fQw2VyiVSAaUsag5Tc0sEs6q0AVFUMS6d39Ok46Mw7HV2w9Tb+PGh
AbJpx1FbWHYc0lsgveYNgCxBAUQPF+90sBRV3DiaB+N+OgmodByBmdkcNtmbumwG6XHplXnSlrOI
nrKC5vB/3s63+uOqORQSdTqyHjqs1vMGmI6edQIAjzhSCQA0AKClzvZDVKdyleJb8G3RfvIifqoU
vObcWHc2HcZomV1j9c1+xbrTs5rt1MuN/8R4U1OMHbErIG15FfwunPeW+TkbjOYD2zS+ESxuvGpo
rGJ+LQSyANDN2ODfNYKcPJ1M8Pnr4x1WDLlqbUmg5f1HtNbuZtkSf8fy867mBW9FahBf+vpxpHWF
/66dT8bZq4A9hdZAl4aB0TYz6oLJdwF1lZQ6GB2BcEDjbD3wYXKnB9M4t/jj1Xc6SmWtwiG3upf0
r28JvD3U/l5fdBpBciWhJh0t/WxxNOyRW9HVxBfHsYNHiqAZvE0iUNGMzabUH6RrHc+HbcOQppWq
EN31tsBGNgDTfaOxZZgpmIq/VGoJv+elbrhrXxJqOXQfOnRUKGA2iI70/cuwflgesQbj2jQEHTtP
1PEy+LQmiOoIhVDXRcWberJ3waZYmYScPOipE9hr2dg+zB+JPRAiYfIyGKtUpCJwjHBcKugKE+98
tw5Na7PLTUga0IBqhCc1vZyIMLtlH5voKo5ST74Ee1Q25txWzPN2O6sG4tCLJTqhzbOvUFcD87iq
SHeXQEnijsN+H1UMXdEXirwGvfo87EZ1/ju6fFs3pDt217beinjBWmKAhJsi7gBmal/qd4WN50iE
82H8Yg8SJnpGyFI+9aiirh1Eyv8KQ6ABPyJ1B6QIjkQJC9iY8cWy5W0EJl+blTn5gCPYAIBp/Uui
UaMsgZbdgIvlMt8MAZ3Qqek7qu8LbKn6kqpqWx6sGyFS5tGmw8GZbtZBoiJcHo6JyY832qChLBDo
mMxSa5e2FJZx898PO/ymVdbqFyBPewF/KFgD9k0BZLWhS5dCjp/sx8SQ8LPw5LU/ryQqw6+ZEoUj
aen/k3V1NQTnWhQmq+RWOnzNOzOXgNuRL2POE2Y0T1CRgvcI6O4NN+Hrzz8AYnSDFozUhC6Y7S/X
xNbtWfjlO2Kukf2AXeZOJtOSHdHCIF1fm8Pf7YCpVH31XZ0kjoeJ9dkzKoJbgTToiIe9Nz8KYI92
19Go5PpICRIMjCdV5J5pHX01G6Ekmzklft9aHjkKimi+JTUco9NHNmQaSRXzje3kSSGIjg192S82
rmdvaJdHJWFVTQJ9hEJHVSxKhomYW18edg0KRRL47l9tANFJsJOmQdI4d0nOMkWBXDTkTm5GpQEy
NIXnVFD4vOzKi+0092dwvf6iL1goELvoB4NkpU+2c2tvd8DVAos+zQgOgv9i2a7Va0dxIO5kZivd
BxJ2JH2lSJcfPuVYQovI2vI2J8N7Pi1xTdv5SXPe2NqHEhHRDWtgA5xTdljyjHDAZC0+PD9jwN4b
dNYvWlNy112QeOqrHEvoCBYZeqFPkz0ZhM4rei4Pvld3Pqup7B4y44ziBuPpMP2wmyZYdg+UvbKW
Et0DdUtQ6Ndhi6OtNs9NufcXPgmlsLOgG6wHgZIgHYAK8JgcKONZsj50t0W9DzvgQt6Tq22BzCM4
36/ZS04lB8lyrxe9vj3h1TGotFukzEe92zIXgOWwjBH1TfFw4sl/B0YKG1dSdfcSdnTcBnjxNnVx
FGAYdjdbvgnTdUFZeJex31aun0ieZfQh2YkHhJhbzPGFpCr4yzP/aXYTVoo0C7UhFwOW+qnFwnHB
aLJbJZXdOEG3M3GwH4WL85PmXjRbH8697j7zzCJy9zNDlM5xtFS88Syr9b/iJzRb7QyX4MWYruzF
b58yzt1yvDTUg901Sq1pdTJvcHEWfmEZv6j+ua16fzW+h3whU2JHxIR3tFII3jrA8fxwnLBJYA+5
3MHPuy5sxuUqfviLg3Hi9Me7wkT2JdecfTTQcdklUvY69yQK7EyKtGU07Alru6UzDviD/NmoiDMc
9HSy8nEwM6GcmVdLksCWyNddFnOA3jxpnncQZXRZYrKkC+3fbihjSzD0PSCIO0mxEUZDG6i3Q7Cw
lelXY+pwIypTBEBin3+uVB90ciGnyHjFVSKnnUe7N0R5YrjDiTRXX7kZWLI2fcdT7UeJwMuw493D
oIiSAQtHZ8sNasSdiNOw0rMLRBF06ZoLy+H85Bq7WNS3NiSkAFjQnOm3cW3fwV82ZsvRGO+8hUWe
RT8CoCVuIl0ydXhy5Zi6gn2oZg1SLBI265t+8exXyAJeJpLI2kjxGwh1E4HGzAg3/hXO3mU0PUYk
n1f77NFQLPm7JKGi+67ez9mXCC+jeBDsjFMwIPpbiNOnd4mjbm5gDnY47TBSlFQZcMNv8x7p4EUl
uw2aC5Jrz0ASklxUtMG1Hd1e6WQAo60PGKtyqi1tMuFhM9QMc8TzwkM1iCN4aahGzql2Ul1GinWC
VNO5KyNfAVnqFH0osY85V6ryuRoitCtTezXDcwJTsEGBS1SkUDQdJ4p+Xn6mybcmmW6RnJ4HoqNp
J9dFQlrZwvt+KdBk+2UO2+w/xd3tF6J1kTpTDK4WsqbVwiqA3iXF6ovyl3ylsA051O+rL3MFYkgm
vNh5D5gCTdMjoy1v/2xTbGgu69znP/zfGI2F2T0fjAP9CMsqeFl+Wh01f40tDhesrNwc7V5YbX0V
4lP9CMf61A7loKBdMMCGyagEPCRmj9Pi0nNEZ9fh1fUQWoUjZJKF3AoIwgU0BX6ou9xAeCg1okQ+
t/MNCCXl2j8OEOJRndWlZvgommteaDtCBn0FP08XL7F716J233M5LZ3lBqu3DcNzmsqQygTEOtmP
BTj1ALlv+mmUxZ8kOCNzkNAFOzUBf2GUySjAUMd6D2bQjuHc6dPIx6QnhrHigElEnoCTSwBnC+mt
AuKmo8X5YWuncRQ8bzzLOVsKb1f9wQwT5kjeMRNbPAH9OdPzZi66rKcsrA+Ops+FJ1av0tT1gnCW
fdqh2plfBEP/mGWG4O9HQxcKfIX5EipxZv57gP6wIpUInQRasE9pXF7V9QHWXWP76XcA/Ncoo5iY
unci/NyqipJWyxxAWLHfmulEI9fBpIZUVk94amfJS93fo/ZcZU1apuqmPKLHF+M/qyUfLVmOzZvD
yFXzrpZ9VOOs1jvfbLzRC6GLb9B8+2t6+DvnAngoz+ihy50r9HQlCixgfRkcfdf/qPRb3ZCmbVcu
LE3IVqg5QhTaVZkkqVUH2WJQyGgDyVfDeRiWBLE3aEkKZjDcO4nXieA0ewH0/aKy/oH+RF2WbIsr
TAzJ9OpedHVC6fN6M25UwMzLh5Qs5uxERHvQX+WwC5UBpyS0gB4FcuJtNCX3QsoGF5yHAQ6fv856
LLaNkhhBGsQCoe9Ik1Q0Jrjiq1Mr3Zl952CjZ5GbkS+JDF62OCeOvEb3FMzr+aOanlVJ1lmAQ0uR
tzXEVTp1Nea1nIzmBEH80NMhqmzPKdRG7GZfS8i4Do1S+EeY7kc9M18OFeU2tV8y6L4pg+XDR6HU
94qhmcMLP+HlZ5z+dK0Yi+Hl3q7PtOCi5UMJskEjd3BZlCBnYAtTSYwPdRw3pnmo39/bErTkSaVY
r+nslKAR82UqL/cEm3HwYnx8N3dPnW7spi7s4wJD7gl9O9w3NgMz6Q1C9chNcRweWTqIYZE4fzqU
gpWMBiBY8woWhwjR5uys96v1fIpCdOSckfgBIamz267ZSH4tZtm8wnBKWVGOxyXbfWgIk4P7NRtR
loStoTc2R051ioGUuQk96VPzyV8eAoIUjDZJuXzp4mfQOABrZNxwGM7NkYqnob9dNwnnEkiQpnFQ
Hlbu5zlkbPmGf0whdARxgNeBhfxrU5+Oi+CSBmlA0wxTGEkZymq7iwOIDNy2LdKdMGK7vXA6IKcj
0iDsWIRoi0iBjQU6GZ/2KstXaO/A6vAdaP+LZigkX2NH/b5FkUwdxRoNk7gFnzYHhegx7u6XSVAo
uDca/GLlHowj+srH5g7v9Ooje8kfmZbZoGAJegbvKAkemG9KX5iEzMI93d7ZZrrJPl0ueBSGE+TX
yNDyFgydtCcmuizrFeC9qBc5B8I+EIsc21NHuBiNgyNLLHxgqHV0fcahFUKxq9uV6vyhzNiAqACs
zZk5WD1dYqqSpRIIuRbDZn+wV4IVHSTfaRgGP8W6oRCEL+8gTDojJAEuRwSsRorMpUiCsYmuYCSk
1x0cims0jdWjLUTY1qWy2NZ3Pw1nTO3hnNUibNAhKBVV2/eJm7wApkQIgyJZI/4DV9Zt7LVKp/hR
wmrPZcv/dDmW5Lc1tdJNUkenfz7YbJLDLHMvlSUg+LlhcfkXRStwaDoFdt+5ZXeU53eeHidx3CmB
uE84A9HdPMX0Kq4ObsREBJGIUKIYxEFhvUQanY7C5jruY9MT2Dtb7yXifIszC1f9IE6fFVeo6bzr
n5JMZhBkM/rdWpTIvzCeLbHWHvSXDpmWegvthYc/jvPicWXo5InaWdDnt37lgI/nG76Mpf8XLEdf
2BCXWQkmIGiAR4zmgt1KKhEu430eAtMcT7R0uHl7ahUQPag3VfHoVUh6lfXmqS8nFI8nn5a87XU+
aiJJxx00oRHr7RBPguxvIElpCAV5rKo2rXzZiD550TC2WNb5EWxBWaWynvmA5I8jEsFbVI81nO8B
VIT7tWy1tBIyLIx7OZuvR6RbLYH7arObpyMRfe5lBMLGnNL5sGCG8dgTYPkqLFucOXuxoANuOVlZ
6taF0AHQ7t5deAa3WzYuSd0jj7e/C1dh2tSIK7GwV6yYDYo2R+bj1jtiwOoiyISAQuWHNEwZn2eG
JCAsY0q47FeNRy2YlT62q7D/U0Id34wcEPUSuuGkSDirqD1MkOkcZ2vRH8LkucaqRl8v+Iwn3ggj
84ABc0e787CiIZ3EMZUWrPvyTJAalFZYZY7zeuP42ks+FGBhZHGNIgnPl5lz92OUJ6iwcqNg3ftU
ubHHiXWIoqJc0oMrxzvilMZqEiJpLPkcysmVchHn9N+VxMAEkJNpPIxbLs68+QWjuDRBI6oSc6zT
B9NRQe/q2+loq/3HuIlR3DP2IPbbInVCTi42LiMxSSfWTFv0+vI3YoXo2RlWweb5FNSKInWxawfY
sn2MaVMjqQRvoWMtX0N62zb1sP6+5NIbbosscWVSUkNfErfNa8kgpyjb14+U2fEeWdhT+mdsxjxx
+zgMsALhkzGjiFpxPLyZFBkwWT3zmja6PodEDD97ORZtzknB8neyN9c3iCk0GROOPXMMIZWCFvP9
j2in/1t0TXIEZEg3dDskGSbUU6bO8V6u+iYLlDtgPwufQM2qdOM3LL6jNJiIMKLG9YR1x9GcwBCj
ZYrZuFDVsJJYrLaDBtmDUiK08hCVrYJYBilug8cKWmBt2j1pGYyhNn53Jrfg6emrVPhF0sPd+H3M
+ALW1pEHbgcaYEqMB8sjjR5CMbTmm/o0Am7vnpm1dazoYecOJWIgi6kQ2M8Z5md5/yWmijEsNPBr
oEeziEIUvQRvgehbL5FFT98f9Y7Doh/s1Z10eVCXhXYcf6BfivBhW/nFByqQaodiCZCM07t/xLjK
FwfCcyBkoZ2vvdUkjMDy3RnOggUbMPvYgGfpiFPxgkfziOHWjEQFWGe+GPwGgG/6dgAKrHS7h5Nz
C6KGJT5XfXnQUrXy6M7CIeMUVK2TXv1mLorkGjXL2pXCoU41Oi8HOuggiojpHUE9DW3L9ZDYLhZa
TmCJzZdvqvBQKwSnBlGPZsUNHARu4ZNpC7Xqkqh2Q6cOZjO1pn2CHZZbvsxaX7gMPTQuy+bvIHhx
EiOHkr65Sr1WqN9Hb4JBrD6N88psAtPptw+A+uYnxAYNe6d5Liee4sKgnZPDnKNb64t3RQ4q7LlZ
5ZHdQjYeiWiSau3aYc6oXr9BS+p9YWuWRH9ATrc99ADGmrDgSw+C1tO+Yf+pNTLk5Acww/y0+0Nf
GrDLuOSmL8XSVhr4nWjrLjf7wZNMsC9bN2/sIdu6p6X+KvDdhENqA/wIJ/LcaGscbmvAHdhIB/Q6
4Q3AZO+ZZDLXTkD741Bvo09+yLPiK0Z5NOoXqv803I5q8XvBAqKdXAr2S4qo1gj46VWq9t25JaAV
F94la0JYeZjUMp8u/LNtElrvOg4etwMP9Bkx2QIZlqVSO4mYfv1Sk2OM1muSamexS87aRCaaH4Bd
f/JUK65IneBtMmhUXPoGsBG0dtU9mO5gCZJJy52OXV81aeXFJGpoPh3GAzvk+gsa5uijMvoXXvXb
W3k4WdKJ7jKIE9g+yjJzUbfl/H55hVEpdN0rae2ne7h1EJ0MZd4Lnn7UrRV7UQx3ByKrX7HKcZoA
nJwVAyOqRQXOzbU4NuWRbLnpfr/LEfiU7g2c/w3o6UkKyxRkbsNGHMYzSEGsXdRaAaeIIwYndwKH
wUt7vLwXTSdNiIRWKHdntsYkxoA3mjh9OGjb6/eYmhD24wgwPgVKcWUQq82+bxXrPHH3V5kOA4AY
VzOWqfSjbfKeQn/aDmh5vdSPqaNaGhAbWB5VOghpGu7616ifjKbsL9291Ly8dBpvx8MsV5TbSpK0
HUnx/rNk62a4pEGHilHVuFP2XsXM2/1YShqj/j7vEZd6+I0RYU3qs4Giap/Nzog81o8M36S4GxYM
DAFf42KJbwoj17wroZGPyylrbE0QcIsvcKUqFCZ0SZygqOUfH1bfOX0ZcCMFW7++YS2UbiV1rSj0
X5WCZlTgZELZhCiwzHiEPEkOHnJiTlQVliYxWW6RXFbzz0cv7FCwiW6p02N+1JcRDX8Ni41i/Bfi
8VeTsscwfYby6B4EnDRU7//T4fH/NGGlvmdRmw2ImoJ1CdTRVcmA5MYGLyfCKmB/HMtYzMUf4hW6
f4W7+vHHT9gkx/Kzq8+vesjBd6B7oM1jpQscmAAnxB2fnepiQRMb39SiJtJ1SKvDANxNy1coMp3X
beIGyFCa73wgSP6SP74wcGI4cs7f1Is1cXaV9LYNPXIHW16a/q0FoJUANUxcbDwq2SqJ2yvVrHpq
H8QsaXdaf9ph1S2bYfJkrNgizISAtu1k8aO9pKJ3Im0r7QIJlhFfTqbG6y82UqM1/dH3qr3JL+Cz
eCQJQ3gL2d1mu3zth1c/rJNQ8JtVuIoN0kwCRqcax123aWPw6412Npyrcdkpu33V6B25JQso2R4Z
Iuw7xm/qTsXF9QOR6LT8FILxZl5U/5K+ILbxhEwHAeL1UqcgD5lsSu10CKEeJj6J05Z0T7QZn33W
Al/vCwy6St08WdtlHKjnynvgvKsTeB+dlWoovsIBU7hzbVCcAEonLcw+IrFA28rmauvTij/KbVLz
PHbyJS5cmTj6z6KIGUtGWFMl0wVgmpptMgVNjYoN4fIrAkmM0qy623mLgxoYJ0+tpclCzre5nw4q
5BGiiN/fjS+PhEY+HuOl3s7FO4XoUPRm7I9RONoezz/gc71Grd77dPZLl41Y9io8eWiIdnwGhlGn
5lQQ9uF8g4wT+L/abl3aaMbfKtMQNLUbM4zSdvFj2BvWBO8rOu4Em8ybagRWZwI0VY7pa1H0klTs
tm7XhaXdBeSYEws7QhWWK0WXdV/deCsrE4ZMxxPwC1H+KPdzc6+23ViRQSqrsRX/JOt19dLTGV9D
MGWfbGKHOBNSlmJD8IRhEqVA35pXoClpC4zcBBnfMf3jlVrmbvOVcneNr4e9uZiASUm2QJQuRtfN
QgElkcF4oT4Y461+O/uYfAJIZmy8jVibVOBEmJqUqj1HI+48izH1b+ztQ9Qo0DkKATwUUl68sOlH
5LjKwZOvXeXR8ppjGSnMvlS4zU2aDDOwLtoq54WJNMdSJyf3gxanCEvbW6CLZWT4M++VbirYsOY8
ZrpZq+wbB1eSw0sNkls2JCXJWCS/0ZvChM4+2RK6Uz6gBZ+yU3kq360XOh3MrQZwCsWpkN/S6QfH
VI+oc/FB2ZXyNM92vFuzNR80os8LBampDoVonKExMLN8XTmSBR2Xw+QPekJxWtVeAFQL6ckq30uu
YS93EDWAYJcHZndU7GRtYi2sj+OBE1BPAOB4HkSRqWY9QBSuJmmkMRGxhfucExqTXbtg0OsQ8F3n
Z3DGL9URHeSVFI3LJKRvrGpFe85qRPixWFCXPkaveEZ/3Cg8gKFoXr9S1UckhUHcDngSEKDUq/dR
uPTtwKhjXR/ttPBS4dhWY1nliFma8qVFL3vA2HZ8P9wMaDTpUJI7sL5Kgl14+YZPwJqrikSUCg05
GpEVDx3Q41GonQrwRl1g/EuONP8xCX/uPvMNZz+i1R7wIOZAHZVQLcpkcrSXh3r7ZXoiO4dsqRIe
KfhgjyDfhxNQ459XZtEYEHrgD7/NdUrUV0bN1jFqFqBdlMoR2pkQ4SOotF/8bkmuv8EiqCOps5bf
Enf8+dKvKepJ/4NUt6yGirt7WGC68h6ZJyfmhWIXMpuVowNKDKBjNpFdCZeUViVjZbwzLVm1AYmv
0E0sUnv9dHQ/ORszQJ7Cv3K3kExbbET/0jPgfdXugV9qVkyjewkpqUFkxDKAHDVJQC9rWVlQvcY6
eNJj03zHDIKebT12O6hXOd2o1argJ8hCaPbVUOkeL6SNSE5FnPbBdsuDpHaVouBR32+vD5ZjIktb
bM8DMk7Q1jjNx82OqdiSrWPjhMvIhptlkOeL0G8LeKcuAGhWZJr1lfwpDLNuS1cUMqHFMQ/Dyaws
rCkB4G7KZvAs7BlDEXcfyOpr4bwRunWpHBowAd/TjHvCEi4dit7RhcHAlKG1ddNr3iVzCaNb9Sk1
iM6Q8M7A3HpC0j7pN7H96oqhAhyzPoS7byM05L3gOKFZ+k4AK4kI7RwCQlG1Iye4yr7HMRoMhhQ0
eLyw7l9/TY8U3HXNnVYojrUzuMUMrmjqMmyhOCsI3hsIetsCDmNApCQDdk7t63J6sVSB52k50r4C
VIc+TsPzc0EFnpUYpYdCtvIPf0GeBqN3nWc4Wc1FAIKDkuGOweGGoNbfUE9rnp+cPt7hC2PKifRW
1hFbPcojx1xTIwLo1sGplOpb7AFMCDn/Z7yTjy1PZKAMVFOMyiTfEwJpksD/iZbEq/khOCjz4lAF
L1K6Adbm36KY4GAI2jZbLUqxgKe5njWZL2gnTa2px+1qrnRmBvQOShiFtPrZ1UB9Fy0gpW0muAAs
ZMn1FS1CFxhc3YS17vH6jNscpAMwNtLzCAs4xf3rIELTntz6J0TQAipTBTGrqZouZO8XQ8iHkPyb
9sB3SAgIB5kaLgbIfC+9cVNUk6amkLQ9wg43p41MzgQnt41CKTle5OrsQLXcjDXkWcXOVALFM5Bk
2xZNKuazy4rctRHEDCNGSFmDhNhEvVIwYgkrQIVjY/jR05huw4Ngd1a6eismilKzpNXE+Mi5TGUk
gJFG7KOIz0sPfRxUC+W/g2i96LgfZGcAcXnUUOL1dZ6unPnCfNWMKhtbqQYAo8LGI4qoWxbfyMWi
8bVYbgZ3r3vGEfB6Dpii9sxpAncgp8sdhZZlINhVCzjVtA/C8iPzn2xe6bBgryiHTZ4PMzfX81b5
DBDp67aMATnvMokVRLtYC3CMtMYlP35/fEqgBw0mTXnx5VwukMOu7svdlL4JRt9o6iEMXJMA35ca
eKM5DTKw+zuJ/+Cco3b8F0ZMwIGQF/yD9iH7E3FUWTH8/ziHVrN7bTWek2c/bh23Dt2tCB3XyGzV
e0cqwIWrochqe8Kkl1qXrs+QwhJYwYdLYkSU8d5C0aHippZPqJtEcgjVeOQ7gXv0eHFTj7tbXzBj
hDpdmOMqYYTyC0oA5HHsWAY4WSkS6FNTsKOWT2Axz/rCHcPjbPs5t1wiGVgLPFt1r8JVgbpc/IkG
VyANhebr+9i2rqHKbAXfoCjGmASivw8K1DzH4e5ZpwmRLjWxjPVgKHWlqp5ZSgTmw6Wg2gvSqf97
PcKp7qAJv2uFjJ03ZtG/vBJNv/NmGtn3wHJHuIkoEvUJqh0MMLx/c5McWPl3Z1/EXGTVSbsoa9xD
ju1ULASD0UYdIoq/0mYbQFfqEv0IKhdIfVS5xg5ZMxVk/TMM4ktGHlBmtEYiWU19Y6xrDXYzKRX/
eGLLJKok+MDgeZJrGnEDkp2JjAE3POsPTanl+DCML7PX/49ijqKz3e8h7wiYEgAx/ghOxjfyEBes
ZTbRCZ2SkVRXA0fjlAUy6P5Az61kIUK7VN1Y4Itu9Cq9BtXFKj4BEEKJMCgG5KRtbylU+JKRJWyz
BkD7fJzACxGBrfFgnZzesdICaKqDw/3hvX+67Au3T08ICQ1Bh6Dm481F0y3Vyws0ImR2/PfE/6mF
R6pEg2mPE7kYy9A2Lt1EbTmGcrF12V8doUNJhWrLx59buOCGZb2wQsrQHm3Ix7+DU4i2KhIYgWTF
uaOJ8NZDN+iOmA/aeHaYDVmxAEhnglTDEGsLvMFA8XHRd8fsxPdv1eTUzLE6ByryEQFR6mPiDszz
gd1oZNnnl1kYLOXPB3vbRoo6KYxL1GuFjSAxqpIBfiJaNFYr+neGtZlKaeKSDdLSPY3RukSt8yIP
1b7XAKziFdBOxuz6NE1HpxShrEjO92YDp0uiBHawffkLgh0o/+8JanffHsPsoCyiKWuiajntOuIr
TqEpUy1ovgjPWxM4HVopqeApjCjgMWfCusOmqVWm119lWO2Y2SAmhTIbAh919ZmD4y3p7uCAM4SY
/2yuMGbMpzaHfCktZ2t3BU2uR2nTHZ2QvgahQoVOrHtidowTQwN/6KemF4nRW4+HeG5xJpYW9Uby
oa/yH6n4IDLIs+Yg2PP64LIOG/7TNn0BazKRmuEg/J2fArhIfGdkbFyeu9I7dSkVJEylon/ty8gC
LKGZ8DALF0HQmYk/7Rh0hq7zQXLRmXolmVBjv0xpe42WmCZfDZxfIUBnEgM/cnPQzLm6jCtRte7w
ek1Q5+ITwWwN7ssGDPBPCAAAWlJZpDPEFAQYzEeiigNe/3b97pG+YCHnQ0DMscelOJKUJX0a4ja/
38VIWRZJwVBLpgz0nwHluChSdSV1c9fTrMssz7GP4NordhXHPzVHYfETtWPLAdS9qMr6MJKhY1dF
rZ8CTQX5sdil7/vZWX3fk48AxYILUJwj38Dfan/WXh0AQcA4xujJZPUe15gRt+/nTCwmAzeMEc45
fV3x/rrloIv+LqENNFwabvAT2RZlKl/K3wM8yRO8bE7/Wh3Liu5rHJXkXIGtgRQ9C4CPkrao8/4s
2wPFEIiO3SBTbYRat7zJiLnxyUWdxU0uSB0A3iGddZHedKPBvIWoPoI3k2CC18uDefnbbLrsZxYn
6dXXEiN/kHyOmakQuu/fsQVQhj6QKBFuzZaB6mHq/SJCFIPh4l9G+gnNaHZnl5Q6RNv87lyaKfvC
IhSRtO0K+j61a65Adeyz1vmfwdj7uNgd1K1nXSrrjpUALVXta9lycZM74aTu5RfRCrOI6MOvmhd1
sN7hDSPzg3wdsz9YLCQULSkFbvudCC7JTdBIzknTTs61r5v3iAabYWFmQxARdc/yMU+7gMHh+G2E
x4h4d+vuj1xEtWkfeQiACjJAoTTDPh9egJqcbz3SCr1SktbggtPMru7fRji/acp2a/jUecNshx0N
O8UsurCkn6IsN0CL5TbrSoMRNYNBAapRyF6vNDjST8+7DuTfJ2ZVT/l+XK2Ra8r0cnxkfaFIIi2W
i/nroqzZGtXDSjCig7BKgsqhlpqs3+34ibEkZU+Br9w1MwUKi+lv1m9riMzeaKvAyCJXRNvKwpY3
28l6t165cDhlCsf9PxJhc5q1ePrmg4YOL0oYhCAxOFx2dvzhCNN57OVo+APkf/til79UanG8QaqA
XH3Q3A7+Lhg5udgvH1ga0xTd7qTIiBzp+yyz/NSwlXcMN6eZCShkdXD1XfTfw8LAn984QsEGfZHV
NfzuM2NHCA3K5yQZ55hk9e90IHK45xxEKsCPfh/98GD/pZuX13Mz21Uf+S+dJn6isH9bfY78EpsG
+6BovxPYz7hjATOnqP/EHtrLJ79haziqys8S9O0CRH89tdgpu8ZkvmxM9pzKkvw5fppUTZVLmubT
MayDdr4e28QULnoZNOY0zeQB0chiGEKIMb2Yc+vHfP7fKZG62uo6Iszl8zEP9CdvTqiQsao6iqCI
5EwKVWlEA/dXhKD3r9ONn3nW+boKyxmrmhHuG0K82aLbOQ9vEgxwwLOKXsfTMOHElBBrdU5z68Ch
530MI0h3rKmNra69HzRpNXQ9Xp/kPDloI3PIm6xD6pXnYf535HlskaDYnlqpivmaZhz22eZYV++k
yn1CqZFyUfMvT2X6xR9eW6FLyZhUv5CoMr785t4aipqPxlmkkKOegclTLRWgXoZy3sWRslPYOKFn
T04fFv2Ak/qKungQoP1TmI9nQIB4xKJSHBYpdub5C+OZiMNPBLSnBQxHGfX+F7ak1JIXgUbTghiI
viuA6U6XaEcv/cWycHSiegRDbDzOf57hkH28/uwQ4Sl3tC5fbolxDg9Ujxj6UnxHyrJOB/SZFiCd
VuzMNOLCcQEgek62/hhx+LSSEIl+hhgvoGsIT/UNSaSpO8ohxrpa+6Jj1zQHPgSGngoTL563NKiO
rKqA81ngWBWZesIo5YJRHSTl5joaYrBAxf5GB+kJwo8oYvHoHNt9JqhaxzeuwHEPcdyVTZKUQNlC
TWsRmT3FMJHGcZWt2vzi5uMmGtz11D0q+ZgJBR3bWzix7OSyakEetb6a+oJfI5VBYJRhuc/041Bg
/M3BQS58fKzMWD/FqoT+yXg1na63xiqHhOkZJs0mHrqlr5t8LCGfwlp50aFB+NZtwjCa1AZLijo4
HYZ5uqog7j/0h88xRrPHcoViuLn/Mwgv9c5S4oH1m6m2NeJOhJHUGQiZgkhK0rULn1m/5x7QVMNL
GOJkvMtiNVVY4RQSv9sCe6kfm7WP726oMNAQgjuLaAWnp6WbMB5ihvewEJo5GaJ1bQmb2nZwsaM8
lUB31tS6ItQ8PddWeEK6Kb8TNnfATo471TPZ93V1fqWN0fkzIGptHEao89Hm2ojXgf6j61JMWps5
RFjIKyp02hzX9ETa8kPMkR1rTuQiicxMQbM/qeHupRPfGwuwowu9HQ8T8ux8svC++1KmuYRew1QJ
72EqmsOvkT9KnaqQJKSZ5KB6cfGuRh/6uxrVwQ10Lqo2Hor77oRRuYGRzBlB2aCIyjJbBZBC1/5S
d07bGXeXmp3n2/O90Jz+PWYam8eXkYfMjHY1AC7QHiUurm0N9hRoPTi6o+rE0/PZQVZPEvI1y0uP
HuuU3VynllrY6QirtJCTPDztMpaq9C6nYabDBDD06oHRadLFWfTa9ZJUh9WPqxKrdNCCmJoM83Js
n4HcyR/B3FYvVRRpPMTa0dLoLBpt2RwWfxSAdjgugo4e5gSHD4CRs9XLcuxsJmwxbSQxPgExD0kb
/10LRb54s4H174+ahPgogPuwQ+kQd9ArgHTRI3Zx9bnwZ04WnW+tpjjDVFogNuYC4+vT3Wku7fh0
fSU5SsCp2rAqLcNwA2meq51WWuEMS0iHAY2LCDKnve+HTiGFjHD1LrmGlYQKzeT1+3/YNPKXUpbO
xmzKyKHvfReoPk/OUngvRvSzQckTiif/NSjf7ambEzb0ALZu+i4T8MbQ7V/zh3pk+sVEBjBN9roV
VtY42RZfTM4Fhcw9rXt9oi2rriBhH/ccw2kXcdiV7K1IHv+7G0XDjwH5iuhAORqb8qJqI4xkFu9U
QmjhnVvdL5QSq7SOVnGAU2d3THcsTNx6hsHxxvKrtynvO9acuH/3eXFMmKRwCk66MZm9/owjI9th
mtJZUgmRnWgFa5LE9vLiHpSnHiEh2N2mnTQQHfFtFBqSLrNP8MFkb31SkP/u4FiuaHVx/uHg6bRv
IULUaTzjJMSjHqVxc9vKYu2RFIhKq3lEoa6GoGpnmTWo46TEr4RakRi7j6rBa4YTn/JDE+4by0vp
C6XkLWvEMzn0fn9JK4AHg3bVHcjmZT9G4Q/FSBdJOleu2Ayl2rDGWTS1HkF91h8n+J4unl6+lBq7
P3E9W1BuLNsytebWqxrQnNQtjQZVCnGWRoMMU7sIv+KsWUpzrcfvWAWyUmqsLpAvts+OFn8Tg/I3
jahz5kSFd2HiUrz4W92tXd15cAx4861u/ybh9MuzHTRmfvayxiLNuH+BVyRfOekkAy661P/nsxlp
AcEYi5kU6L7PgBvemFvpMyfs947G9aXaEerN+UBgnXU99O2jzMQiPauubzodeD27bnB+UxyxApDR
RsMRoC1JVCD4NN9F85wlCebpuKNkEMl2oicISSNj2xJSGcbRICid/fYMIqUsKAkktK/dgXg4JS4a
zL7z4zriVM7u6gKTmoonYVJB0N+yeZavqoPQ6RiSNXzFG4wwDaC6jdyhmiwbLalnYbPAf9CwFsvT
YdH+BMOr9sk8mRZeFBR0KUKI5Oyzufnxne1lQpJ8hrfWBAO14cXNr3L7hEYZN+NYYTRrFcUfkci0
24jfKuysLrDhexlF8sR0oaZ173oToTaL4AE29o/t/hP2Myva4ywvey5QIMqTxCXVxqoZ83cJbMac
20WJ3DzPj1SKVb2Jys1Y2bKSQHQz9XVyLBSr+9WVOS5JzR6I/E/2C5m+eIX31fpOsDMdgbUB4//V
om/G4xpqNOLB46EPj9El9LyjgLrUgFCN4AFGhFwDJBrDXI1qSo54sWZGft3LuDNkO8gpKGdTFnam
kw6yofyTvNf/pnyJ23crAwhOcRX3c4IkawJB5p1aOFu3BRxPokG/WRy38NdxiZANZAC0p7BS115U
iZ7/HF82/bIEyCVAEDf3aOpY3D1gnYX+h2qw4l8mZvlL/VrItwNXewW7NBvU8JVVXq5u8S2M3Wad
5fYpFRmrwnaHbD13zEHeSYpwx2YqyCaXS+/spVC8SpRdhtHb1rPWa7rIzV6+CzB6Wyp7CGgI6Gg7
qA7/krOhE+SZnjOFkuxkQb/IOO7IuZ1N9M5+NrfC20wRW2ygCpZmfc0P/+xXWWbSXNy29KPQV1in
neuJ8Atl91d/g2Wl6uNKHeS3nSbZ+NaU4nk2p2ngmtBE5v4NxsauRA+C3o7ZFz8LAW0o5xeJE945
bIGt6borO4dxwJmdValx34bkzVN+1BYnP9vqRP1783ZcIxHMIaSYkqZcyrW9H3cTBRfnocYbY+K9
R2iBxA5R4afZ2dLb+lFkgA20VSa4yVEoJwvhCrSNivaX5KYP2lPcA/JGRBg9CtAoQH8q67QtCl7v
rC/WlVO20uWgxS9v5SRZwo8Bri72QSSH18Y947Ep5CmTjBNHneUcKDVxC+67a7pj99FpDXuYFu98
neqdOjb3NCQHYjBm1hnwLikmVCrbIZeUqnrEuZ3XFHoXbVBHxz5HUmVRCZF+FKFrIhAKyxhESEP3
bvabdSKM+mdTKaOXey4MtiyrGrUM8AlWIv+f82Sh6rtedzGqxqt5VwJifx0c+J3qj69wvRzwomfX
TkQcn3kid5/7gZGnTtMkjl2eCHjvX8T6d5KV7Ric7aKnGPpP/tOBbIiu2PjcbV9W+IfivtATijWu
QiD7ZSCMuIbV94KcDENr+2Q9xTmFwsgSykpE2a0+FLr4rGFCSHBr/z9rLbRxU/U0pDRV4TR1DXpT
mXS32U8rs/fWTHkb/t6YSaywbBDD7/V4lsK1btQ6t08IH9kqm4DB8K9SS87bi8q2qw/9QoHxz8wJ
E6D/FjGIlNvTsdoiPm78yPbzwHkXHmsZ24n/DURmt/Ow4hdRxhQ1XWeElxIKGPqWFFMe0GcVZcJc
9rNnVCH23E0eLWvDbelJTnV3eRtRu7y8if48mtXXl4kRBf+J3269kBAVnwaR8VnUXuHa0QdwTZsz
IhGPHgUA1aXMJADNvOptM7NzG9lWENW9erVD7C+LZ4gTV7+ZgclDADAyt82OyeJaFs2xHdri0wPc
g9SOaV5VFCIJUp+jRiLMt7icyPVFiQeNDV8wHSPfHbHp4OmqaFqQq761Ge5bDgJfnIr+VJDheaqY
MqWE0PhKmWdx0RW4dNKM3yv2HxJwk5nIHge/1a2opyvs0OLq2GVb8lcmGXJHeHBpAqtKyXy+q0zy
DLJRq+aFEVOxvOoRwDmp6swrQbrE5Qs2ZQSkJZBzjVa0hdDFEM+cL84dXvLXfJO2rGVd9XtUf3TZ
HnIF15DNPM/x15NmfJVSftwjdjwaqZddxwvthIeKeCLha7oCxfNgdkPgd/JUSK2Dj5hhssR8Q7b4
mL1ZIUn6GPAAk9Nkpr4/cY7u+9U1NRZH9JsxpvR7iKI8XW49OEqYx8K4357Opdss4HXFMymStdzx
d2NYLObazeVCnkPtIuigdxezzoIgca7UX88Crw/QYZqfME0dtGgqDx2ML9pWdRbx8cjUJUwocby9
I659jKQryQx6NqeO224pERFHxuv0lG6XL5u4CoCOONlOtFhZFM+iJrHAkGLvIu4MnFhQuEbpX7SC
hRbtpFtaav+f0TSA/AA2RGBFl4PVK6tQqW4/UBwWwtOq/HKeMeL/NMxOnkGESJDbuwRX+boScZAP
eraWAuLsTjGv8eJ8GpVXS82TDfP3SostSoYZk1S0/jpaWCKo/yPJH4uiAlVIKOYl4hDaenwP4tsm
gg3m6NsQc3rteq91wk9Ywj0JzZQ7qCNExY6LLZCZxKH+AIMlpgcyH+bjOiXblEwVS6XdfGNioMRX
Aa8HDdESRMuKHF6o/VbKxD0leYTJt9hE7AyINFeq4bMzKc9ei79uLkQV5H9U7rWctLAr9iuax0Oe
v35HeeuzB6oAbtnW9KoBc0iVuaCuqflD01oPWjL433+lWRHtraj0tzB34eQ3VF2tiQHzT+J/qU/c
Vtb2MDPtWbXE73h+zvnAuOenEndDgCFtQ2x7s+TyULkgBusZlCiiEr3F1iTUUznnNpv8AGuoerP0
loz7IZsVNoHEa7dFFsChOyU0tZX8AAEU04ZqBRoiSDw4sdLygYzU1Wsd8eBLUuoJjU4pbFu+oQRU
puZxHskFDpU9xZsS8xr3antjkO3HxwLDAE7Rj8JbDCbgMdgVNA6uJgjUE6GRfU5UIpKXBibyS0wY
V488G/iGifxC6xTtHZ5t2vpxZlO3KBciKzKMPeKHtSw3kCYJqYCW+ACGIwL5/Lhm7fcjdGjB2Ib0
F5eqWPmesEKdVDgOiqSVYfTxHVkJrI6lsBKDqSExoHY6dw3Q8MV33JhUx0SIvActJ2rN7VghrV0k
mCEr8pr8WFt0xxNRJF5mTMmnQzJF0TymIM0pqLdMXScI4KWoxYXyTfWI/4Ksz2Lu/81MgmO92NRl
003UqOKtv/y0m1mZkxRv+ZVDz67KEZbZ6I0ZO+9NJV+1SI34VqWpig5R5iUMgd25BRiHHX2h4yug
jkUn+FofTLpuUKtgbKJpUVL5FFzs9xKDt8a7xsWJVlZYx6uD8TR97oQNNnv/2zvwacPswp6ijBVs
J+EOsUobVov4SG1rV1X4S/1HbwDjRJZ8WMJeH/A9ZI9uZVpLymMhggl0BKeL6gS33hcQcvwv+ZmO
qysFLVn1vNVloKM9DO49HUG3wMTYp9qoXaIcGGD624qtPYL6VrN8OUtX2zgsr9gPbC8p2nA/5wsJ
BnYKD3qU55fkaWJ6VDRvYrmSKXcqWe0Lh8HhpFPZFwRivsDw20570xnWMr1iJp1bDUd0/YD+j/Sj
4zjYhH/rI439/L9nmbhNRq4IjXh7wgKdAN9BYYCGqDrVuMZPwrURZHpviGSqBavLF15lzj1p+nQM
zWiWI/ivIL6cpC37d9UcbfqJ9xxViO+w7D1x38miTLkq1o+WimqRV9gXjIvcpKm5sdVz9FU2Zz1y
5BQHVQf+zNSPZXU7rBOuj8r8ILXC4UeT4n9tduyVJA1oXM7BXGmlM3YU6RM4JGd3DNqNPfe1LvZ/
OYt2nRCEDBJaRROycyMEs9y/bcGQrsiOpEXESsedHJVpzJENYdYJ1sFJ1WOpN9jdUgVumbzzRQ8Q
t3KULdhDzxc57yV3E0UhLHoZBCURVvBvrUH+Y24HoKX7jWVr9gVe9twzcliiT6L3ttGYglG+1Rpl
vMkmk4YB+42wb6d6JaL55qPe70GX0Of+C3mLMxh6iXsIA9HApTRKifBxDcLFHt00+qAAfxO+K0zc
0PGyLC5Nkfi7q3rg1qv8djfttsO31I5KkBWIiPQQ2Xsjzuf44FIAoRvno+mv3FV58+XJABYZty5W
duS/E8r85S/3hEDLWLqLJNy99qBvV7PqJcQkEyZcbjZJJXB1m7QTkgzSloNhLaDVggzvLId6OPk2
K4Y1jOgn1M+SMh/u3t2PzHRszoISDKHeg83W7xwAqnr1uXsMTA/FiM6KDkR5rdny0lyqye2a4toD
Dw+ihME+ET5gfuljrbetUQzNcfu3+nnfOqbRhG33GoGT/l1/mC3+dqWipf0BOxdAi+hv317mFZBx
+kpqt4OipU8xOeBdBVqXGIdQo11f6S3U9N531BVOkAEEyaXDl6lV/MiM9Fl3x6NKsZVwjsx9AvM1
0QG+urJQNPYkvPrEfbZi2cC3lRqnWU26ye0Z58XjUhmz/UTWenwa/iN9GChBZclBsZEiI/ARxya+
EJXlMi46mApYASOJ0Kuk42m+Jq9B6lGvd5RnyS1WjrnV+/auGAfJRzfGD/M01MDbGRAVhHvUiqfw
s8xUJMsQr4b8YkM6TSKDdQUl6kTdqQcwc7JEmEQfrwXphfk2/4oaQx3g7wV2g35fZqawVLHr4Szh
3FO0XW3Do3BZFasGP9hqmIDumSC0XyuCVOvRQYY9HXnlic5/2uuENZK64BxkwWliMxdiUXbJvz2t
XL0fFqVzjcMhZCPUE5bDs4JXIKcI3vRYQJuBBJPVKkiMlA004cCkC3j4zYjGFPn2G1tn1LOv4vQF
ItSV00wHirzsfmkmwzraKvjCp3ZswtBWH+hR/csa2MMswAGRStleDIudQwrts8gbZmw/X5lNqXm+
c4bEZUibw3PHZL/zppfCvMXwE1j5+7oritLS9IQ7E2CqdxLmthOwcjueY6yiLK3PvqJtP0UESXu3
pGTfw7l43pdtmPZtDvIa6+zz+zbYKk3HmNawP7LGqp+7onQqbD9kJV1f3nHnYr/luR9WCWURWWZY
AL7hFtCzM0IzQNSvnAkNoidj0vEAwiL2xGBLp+CUVTE5E6hp0cEn+URYTZUkrk6dPWblFuXZ2lQ8
9e//kbUcLuo6jPQevFx0sGyQ3JHEk+qhZze87wq4XcqnAJ6kKbfBKtmKkMa05/nOutVBieXnS/q+
/Ll694KlNI53LGQkXSJYWYVzxP5FFS7WTFeNLVjawh1lTFYfMvwSICbqyQ0Vbdt0bEm3820aR3Qy
svpET14ypOx3+7h3T7p2nvX4T1ThKGm5AcQGQqZlGQv+1ee+UPDnkGsVQJAmmx111+iWxZO307wx
l11q55jWd2dfik1zTMm0dzQHhZxAiTEZL78Ce4Gf6I/7OF8XK//vIHJgaq6WsuJ5z2Y3IzhM3Dio
bzJhGSbYPkkyi7iwnKLd2EXFEYe+GldaakBy4pPxum0Msl2nK16+4d9jiijB6qy41Nn27cEjbrou
scnxI8icphPSVxeWQjp4MFSdc4HMoc0nx0GuzJ2hmYrYXoY3TiBUHTetZfGgur6C/0cSTZ4utehU
kDudkac93Ze84R99NR3e54AVLuI8iW71IsiWI5SfrcjGfVpRVaH1svRxuwiPkjOm+Ufj+KxDqRwY
MmpUie4TxQY0ko8SjbPdPZk9kAdJDaEvmxFy35CwMMf6TlWm1Epec59POwiRL++MMbub2pUqYhL+
GMjov7Xy6SprZ+ghmJlPOGzrZcEJzjY24O8MRE9PJkZi3EPOIwKPmjy9wT1TcbTEoe1rXbDooG86
WjfoemSzo9tFK7UbEtYJV7b0dpPHyz+BIlNsKJzdBPlK3/3ONBi6sMNrun1gaRmYzhhokQJgf62m
r7ELlDRQdYD/CNTCPl90uuoo7mynFI8HNgMdotWaMDmleisTT7PqbI/geMVlI8djcrzPlhMhwGx4
7UCqwNgvbxgLZw+3Ipv8Feg3vhPtDkGql7NxUr7sFLF4ch0sU+B70ZVPZ582sFnrCKm0jkd5T+9t
fWtWPWwXYEwN5qnStvyb2xY01niV7hi4bKtoXdw+S7K2dRcn4SSmVHJNpTetaNNBC67KuJCQS3Ay
/kpLVWI4rl2MylvwYlzIf4KLNjes//+300lu61MmhVbCRfwl+PEo55zGD5iREt6mLAF3jeT0RSiN
f6TRwl5CHu/IEAOO9QFcCKLFloigsEz8fxvhXAN901+ge+K2MQ5QEDL5EdeTnIdncKBEj7HZkoU1
bbfzhGLK2hum0qr4vDFu78Ur8puDLO81B+j437wUrIXw4Lskhs2Eqm/9v+vHb0nNK0voL3ObiN3v
tKo1+Gs3UDcZy0ltDtD0khesnzi47rIKVOCMJC4irwIxwVAvattlrGbX+KZvR6iPKqXFQKf0C/o3
dsUmFnzpuULnhkYSiQV9/bMoSdj3IoEYpK+1lq+h6FdWhg5nctdHWR/PzOd0RK5gwjnxd0Nki8Jr
/0sN/Uhv9AAieAXEkFNQc77E0DsHNsrP8LGoZzlSDHWvO/NboWGIUJBM0KJrl7drkpzYwbER96/h
89O64GoIOeMLVto5EdeT2xcbyHk8WPkaTCDJs+Jt9r73RkLF7h9dmGnjFr2JpaMeq5Bb2YRZryjv
vz4iAjizCGXJJU5WXtJRHuQMGpSHGGqGwcBcz/7uumR3ccAwO/2DUMK2H7ahv7t45N73H2vDS5WD
/K7RAubhYkeUPjc2H5lByCbU4LmRGtOoO2nRw6FpqdZNfAsdhwbxaAWElXB5zAdDNdtTZ2fNMoVp
Q1giUkSm/pjnRceOKjc5u/JfXpNMmEt9v6SjyK0Cov2ae6AZvtgn54diUfcNuX595OpaAkL9OrVr
aAe6fyFiJWXTfsBuOLH8YaVySWikpB9eiobscI/sPExla3AOAZ+fOhr7w4fE6qF836lN+8FR1BbX
6Y9RH865s/eHzWIm9KksV+Y4s3WzEF8zbC+qwcFKXGra11dZJafQ4zAxARXdZ2jIO0lgdIww2trh
Mf/Szb7dyz1DFyOb3VHfmaP+9r4bO7fesTsMDQYxrJFtRVPmUsXm/zbFYklLf7IuaneNLC29QMsw
eNRVgu96kEnSlZVw/neLE8rFA+f81i5jk6vqC4ML2iMc3/w1zSO52uF9tViqjsSz9fpBU0GdceTA
O55tn6Vo2FJqhGFxVNhGIGlEJYTEEx00VTe3VfV+39ZU2Ydu8dJYZRbilpU7zYdZWzu4lrEGpT1i
o33m/rcVOFqSXGjKeNldmJoqYRK/ykLBhibl6C0Sd2Vyox8YsH2xdfFn6DSXCxsExPYR1r+hih42
bMwlCaVQqqQVs3rETxk97L+O0On+aT8jrL1Qp4J8vPSEUzMPgx0mAYVecer3icihkcIdSeQijmYM
Tlomz9H5clVONu1mp8+pu3ob3zkPDw/JKVma6VD6a2pd8gCd8jmp1B+ahw6qcsmTxQsykZqa6Nuq
1QbIAff+pts4qrU6UO0gx6/CRf9731tpSFFNiE8ZiHIF3O3AMRIw5DaXKdhgyqa6WwS/yWGs7+DX
KsPD24WBp20NFjuXyYDunxAw1cJX6AimCzRtW36ujdUo0LVXDbdYQOLvmJavtxAXHcpADn3f5xGT
z3HSvIhjjIa7/suK5wxbJwYuj75LDjKzg23FLyBQEA1WKx0kyp9bNGNU8DV27aIXfL/QNvbh0A65
UT0RAfC1XBYfCavCDNiCV4zLZKvIX7hOh7r9Xalt99DJ330+nTL9+nzm7nSsy9w8VSVk58k6tLE0
LHec9sU57Ofmz33FNttAZY5EW7SEH1uo7XYLEsyRyRjthE7rOfC7UkajIiU7RNCs8xMCmAREEPoa
q/4Uu/1AcyAiGXGUdgdChVPhgkPSjTuVAZRcn65hq4zAyECwatS0qC6WL5YdvkdOueT91yTZTA7Q
mm8Lly+v8PTiUZdhRq6dtPrkD5KPLqHADtu3gnaJ3LGu7QSGyrnnnmh52WcpOc6CBYMgNpTL4c8s
JIkm/+umJRP72IKPsJIH1TGhqgN4hExcGiozz7C9Lb5DBHn6ZMGZdeYHcMHY3EmKd/FxCy/OWyvt
c6Xesx2XILwPxaKDSucVrJ32chPPjJ0GTqphs6i5LTijutUKDmwCzWFlQvaBSnJw3GOABB46XQLH
f2/KDzSTt+VdG4l2QGDaFJC56PXvJbgYX0nDcfbu0LW+YxzHLfxlmipBiZg4TXYLNgzDlIFHgzP1
ig/wyXRTdUiGGLg0spWhSdQp1GWkDyOCPPF00DsbvYVO1oZig7dHqKXW/PECymnfpPFVzfL707LE
Qs+6G3VpW1TRv8dfiaJ7LCDF0sJOb5v2rLEtguahVXJy4YYTjrQ9CLyzrdXn5NVTb9Xs4zkyaxMW
RZQaBYPwAe03d7U8zXF0+7dYy5VZP3HHdiQ5MgHk6g+f/Yrj4ZG9fxbkIRFsiyCBRwF9IGUhASGb
vSsdpUiWc8DUpm3jhvBJePPI0blTAS7BAQNPP0x0jUuc5EByPRC4o7FwuaECd2zcQMRuQ5tqgaY1
rYj+QfjKD9/TISXO4K9yRdewac2gJZSxtUoIfYe91boiy4r2ieHe2igwDyf4pMDuL4ZcUfBvVNr7
7jWHbeMoglLVzcPFg2PRLNrVq6lbceHSGNAIN5UWJSrwa4guUpfYXPmK1DIuvdnqWdSHI4tUj5Vy
MwN3EKqKRaMWzXbOl56Cqv9lpvXYMl0mxYghBF7fS4a3a3AB2iLvs2B/7S0y5Cx3YzGsAQ16sEPo
eTL7WkX9owV/jSj6r8vy+dfrIAMkmGlr7DL8PDdCEwfeeRYHPO3XUqCxKBDdmkWXyQ1NAO7aQpWf
LguN7OW50qY+ndCoptn1yvtFUsV0ZWXuYCVfGf5AQdbXynZ0LT24z0Wi6f5YUmwBAXslT+4FpRoL
gUmiePd+iUWB+NcW0F4A8F/2jqhwLZFbCxOnZpf7nHNUnPpW2U8QyzCAD+TVaYJ1ZDeju4ynCr5U
BYFgyOY5MzFKuDRHy46VlPnpFJDBcbhroK6red8PiZLwvuLcyHfF4zBUpUjNDRMY0IVKzmVdoW26
xTpjLcH+Xw7CRUKnl6OJ0PxwZnjpurblkHNl8+ykEN43inYHVksxHOAIce8UjNNmJMU5m271Ki1E
bXDnm6rgTJUepwdph5OPol14dZ8J7Y5uTn6qdVwWGabLpqcNy1+jJK4SoueJB3hFC+GKz0K3aPPF
t+2aSQmsKGqKVra0q8vbtpC33B6+njCB/bdcKQhsdh7VVi+f/1FbVKxv1v+Hsn5T2b+ZISU1TzyJ
kWrHwOJR9GAGLkeiwDDHBcTUN5yOd6h/ER7wwKmI1HoaujXgNKEsctWDJXHiNjH+zhuiuxplLLWJ
G/Gsh/WiafJcljJaU01z/IP6GYrkaUHFnPTAyUnEy0C1j6fWCh4Ht/3jDAGVPV2GRMyMawF6JGH0
O15cBT55XzdutbS/XKPSsc4+YxoeKP676xssEp4CyDkKnbbUgiEcerpSLqmZR5FK4WmJjS4/XEst
yFY8R/I4eqcpSL3QRZV1E7Gy60xtemmhFzY1+k6JZeEVkNAu7h9+L4a+OXcmK8xJDtmtqSvASdV7
ppQOOOB1z8XKU2t1cYnGNkXp455PkQdRhcEGyxYGJGn3XgYFTGcfKtGebP/9UrBTFSMIK7eqekDL
CAOUR3PHhvXgelpR3Bj5TIst9EMeYrkThdlag6fYsoq61OlnIWnZzXjhDjCnukysP4zBLL7oH7/d
WtgMyTziSB2oxINCmzXMWCZEqTz6pDmLqvH/llZVmog77N2JfW1ewtJzADBz+RS4cbFMvYGPjkdY
Jm2V/kutZi8a2/w4jjema9tiIMDgJPMrE2d5pDGH/7GavBtgjz9nzOfG3nqTbo47hrpPrdBu+Bsg
ZSfp2yJaJbQNe6lzaNyiSSfDt0VV+lrwxVskJ7/x0Z7vg1BRn1TA2ssLkwANVhsiORJmc6oE+w9O
F8qwUCUXJ58k5TSi/ejbzaA92Ok/ppkHJid1CY5TV3sZ5IrCPiu8iR40iwoXvF2FvomReHhXExGl
X17QZ052WrOM4bPo3Bg8w7mTmWX0LvIyBrjR/DyP+9OGNLHIYlrdcqqgt9p+y8LjJhhOR+c/E9//
DdMWc/ELrxQUH/mgNrbXdHwLu1ryaQtpsAvusVPHwcwl9o7SB+mvkgvnWyf6VMydWD3nPhdfTief
n8o+bBWEXJYVbgSKbZB8ZKBJU76qrchu11bnpWWjm/PGxIS0ey7TyckrYig4TbKDCKHMC/L9qh4r
0bBc1h1h1KK0hL2C3+WdmrPEGBRApUxC2MnurZjvftoS27dN8D0I3NuuuGFSX7uCq3GutyqUH4Hp
EvzO9+wG0recVgJHvXhvVtxeDKDNxJeluCpbGrX/Geihj8Lr8+mQrUrNW5yGW8GVL4j3+mMeY+FJ
DBsRlFxFwQAtWGGVSEf0fFPrQfgqRI3WsyLFnqD/x1uIOwmO1gtR4nv8ZN38p/HNQHlw2WB0E0mJ
cKmoeWBrcIwKqNPs8WRORKwd3N/+xxybTOoUjnjK4Apvd/ei9spDJl1jeW9UTRnduzhTJnQ/k0yu
c17bLq6AjgLYAjkOpI9ytfpK3Sb21IXfu37XaCZir5R3AqdZ6iiJcrnezTj9jgOftGI9RebWE7zA
HiHSaB0SoQ5/Pwd3wTtqH7O3lwX9MiztQzdbqqQi7Y+NENAZ89yFbAtVoNKy8NO3f85WxQAM5sHF
2dJeMfOl+lLEdfD7qn6mGOGZhhNN5bLHX2CZsv35AdJMwoOzta8wvkk7kPf3b+mJYy+mmp3AFqfc
qOEv7EbMVvoCuGKvC907olUHtl9ZtASYEwTTSbZHhgBlx2xo9821HPEuyxaGxPbpTEUG5m9BM8bi
BC/EA6Wi5urIZJLilHwB5WRfE30jCUxEid1/Yr3QIbUSVY1E0nS7Iu3sE6SgBd3vTsjLtmQYFHD6
2Wgo/nwwZzFjnbREnjW6MaUbUmWLUK3dnqsWYQnjGijkIAscgbTCMe+wYvejyS8rdKKDJ0BBfN7R
ByeZcOX7zA6IdjPdJRbPlDd71QIWpzUdi0Mi9IVuAdzn+M0LRZDKCxq8Jqe4MwqLQeaXhYxFvOid
f6iRQNy9OIWmWDuodDhNpkd1bjlpC6ZAtdktCvgBbSBEpHDIvUwzXALcP+QHyDnKHH1T21BLjuqG
818fwEmMh8doRkpF9cyRVD0PmDepf2VI25imVD/S3YysK3d2SVFM6kV9czghRVsVO0wiAW6wnm/I
+BNd9AJqFY2+xn3vnHY2VFewxm4j7KX0Uhxbtz1IQr7ZcASPGuAOzUdLGjQXnFyo6kzlQkj024mN
NHtUZxuKaBrtnKFh8KMEMj2RywF9QG6b7IqdNc+lreDrcDwoca4adUNnt60LkT7WtKBKip4q/R42
i7IuKCtnVJcY9BJykjCdt3iw7vT69hb0Z2DMxz9lNBDQhEm/ZoaZPd33QEwtQt8piSNn+7wxsJHW
LIPWyNInZJ5RKU6MjNxFULhS177pUfcUGWL+4Vyu/PNH8ZYgH14rv8aq8iKrCSJz327n/h4sd1VO
W5dYJaTtszlmNoH08yh4vYe1Al7Mg/6hMME/oQF93X5wPAxUaFk/VEi5Cgb7fGl2nJKrM7zVlLeA
IiBuAZRx3oFU7VMSXtIBJ5aWR+SsCbPKYRqO7xAq6FTSOVsjVZ+OTmSaMgQp/v+fSPhQWQm2O3TH
7HFxmXd5cPDSt+UJE3Ol1M1ONmvfUPM0z8eKX1ahOufUO4iGEljjbOMYalqNbfC8m8P9CeWT4omr
/9NZsURzVT2Zfnason2mQ9nqgSFFsbs7hv9Mrqz+pi9M5yQV1jqjpKLC+bqaCE7jr4h0k8D4k+EL
KZ2F7Bi3I4am797ufsLoRoMX8Sj6Parni1c7uv/6pRzJVNDuJA+j5mo8kxzKjD1WsKwLzdqwrnAr
kzwUP6YFvFJPutrzyXHZqXYm9id5Lyhf+KW6/DSCojlSkoo753zzeSS2CdKA1KBSHXeUcqtPJrjy
Bz03QaYmzbniR0UfxgvqXFhYbWqlQHW7GrACrR1hyyPvKf/CwzdrtP7vix7H2s7ychXC4GRQz9XU
h6YQ0XeHc5SKmvfPOgF6NcCY/DEqKwf04S0UpxMnZhE6Ylh2+a4Zimwl9D5aGPGH+RunFhxaDcVk
Ux7h/cu6AWe9se6Q9BQgHSCIJSFb7VnnJeOJY6ASGpML0/SewPAH5xTotyL/ykszKqhcX0jPtO7/
Oa3a1RzWFy7dqSM86l+5hRQa1Yct1sCoG+SlVe71EXuhZvRChL7htx0oMKjybn9ioNy3jTFUNu4M
Ras7am0yOLxDeLp+zIZwWaXHZG3zMbimjr6Y9nuxdXoUBWghPt65dN/fWbeUOPVfW8WkXn33RPoG
iYPCCfGbpljiPRmfnyzrofLRAshmhz9viOOOIvCCwVSmMqSq0fW59ZeTShu/pLpr+GbPn9KG50In
85t8WIweZTjQlRPcvsDHCHOl53noFGtxVNjkTg5rTx5mXL4FA127Jg6JaAz1Bf/hMCra8p8hbUq8
EHRQR0fymMOMwPZc9EishnkqSBomKPYjXgedFrDV0SzSA+wm96a4fF49QrTIUDfNv465AW+Umdzc
12cbSdkN/NDyMTtcakI7+VFhLSErJXus/W2m8OHkqrcjomeyHBHKCi0SXGI0cbPE7SADygtP2I0u
eQO2+jc+8diY4tcOkpJV4KF6ybtu7F31NEt5kqoGdCPM1BEXwoww4QIGcv/OC5edbi+j9oO2Pez0
xvXMbiugZ2rnjwgepfvRSrxDlggn/gMPdJo3t6mjgeOsOzV95Jch05Xhafj0fxrV60sHeLpy5QpT
RWXXiQ0/tHFQYGVQ8hUTOXpJFfvbD+bKf2pNqBnkbAY8knILZ7yqsUQNfHpDbtsOo7Kcz99S/ihN
eAoShNBk6Sh/LIDxfpKiwax0FNzeEC77FLmf42XzjwzXWnSJ2Gye0n+xS6tlzIObl4sDFwL67Pv1
FeGLgU+rBrbtycVQgLT4on63X1Ce0uj5R892QoAfJZzC0DIsewRXxVNtK4u7AkY+Pixf61lvzF+y
4z7OwCu5cVpMIVTGj+8nx8KIatQdd4HwYnYD+X8ykv3G4HumwsEsbejcTweKXIt/OYa1wbVoMuzA
i/h5ZvwgNyI9Jb4NiSM3jTDX2gYYK5r7AlaqWYhR849H8Wvm8xewC7AagUg1MuV8z+TQMzU4RkpN
ONB64kOMyg0qe0Xy9s3lUi/jO/olkJ8mYz8qkyhvzoyrHUQSP6Qhdi2gj2doNYai0Lf2lp7HY19K
OgXP6ZZ18ASLGH1lbyEPIVExf95yAxQGX0N/mUfYKHviXuPJtgK3a6jQNsCQ2C8Ul08wDLVyX9ur
FSlWwS/Y0EBBR5Z6FUvN58chDo9HUDidpvpP7WO3sx8TeFNCgZJc3TZReiG19NB9XGD4G6LO6jI7
KQAlooSDTcLdsncCyqluZ8URWLX0LjnNDZsXAcFt8SAst3xZrYUM1QsA8cTBj5pwMmwQLkNNT0TE
zUyIZ8INzM66tLspJxv7qLgxjaSMQkd0Hz+DF9pZZLNb55anzYCjkL1GpF5Z9yEC/7qPOhBzDf1+
AwtvRTaVA1EeuMwPy6eSv2F/8UIqZ/D1iF93YSymqwteQUyZEN7BVfWBqAF1wgiux4yN0SxwLcTK
1tLLQNBF09cV8sTH0DqIXqGur2+Robm3P0Eyy0v8moC4V4Oo+I34BdWR4QOjqVS8Cq+tJf6ThWdZ
XEOfafbDg1OhA1qUAAhx/V502PDwYrvxVMu5D6xpFoft8C+eXrt5efWndBtaTntGnRH9Txct+79J
zUEYjXUc9vG6HVKVE62o4Hc2gkRdLjQrTFv31mYoo5RvGpSqlDGQjWhcLzkz1WfCZKvqrkLZp573
yZRnhSmTwjVVoPM9aDj7dXbF0yeR3J1g+Mtu6i4a7vaSrXax9vXl64eh1zsw4+mZNUnF8HSCNKOh
JE7XD5GtGFItC52ehi1eSJ6DVhsMxGNNXjlpZLm3UNlfbYMdlHlk8chCI4rPZ4AIBmrHRZMlatHJ
arR2LEJk2FwLE+Z3Id5y2uv6XoubxecrxGuvGtQhTw8vfyaXPjLJ3aj41Za/IRDNo76f2xfp537a
lJQWOWISlm8QJX3ceBNgutKZa0vTvXRqEdlWrMAPANZVgNI0PqvqJzVGo9EPPOKRynHtHhhcfmww
9Ew6T+W3RF4604UJ7nDURjpz623BZTifmwf4evpSTWUvwzyLnN1GBI8JgHrsFtWWT91uQy/URt5B
f/RG+TpowQLSN1W0VVJhrGemYAT3130k7Ku5Q/B6zubWVDa6NLXWDZjWUsdN7mdB1nAmFZ2fuRIV
7E0IJPEola4Sb+RQLdFC7COSb+k1ynVOmNHU7omUuPQNaeg5vHwAqwiRLWP2PZ1uyHewi44RPhpO
wD7SSgin2PbsMPwkNW95UiCuLB3sVMuJJLGS4zJSecEqdJfVfM6A0FLFS0xbiGsaJFYIQ0HUjudX
61cHYrty61RVSq98uz1DjHMNw4n5XWoZ+pxkHUXtwMuWgEdl0gLlUYMiSHNoPAbkhKE8ok1unvao
gKtFzgBOWBLCDkj6NNcS2syb7u+QB3KCSzNr2yB/bv7ViY2+1kIg6nhp8xKRTYNHvdsUN3W5Nu2v
CEDD53/JoHywliYt1YzZ5zpdn9mZiBzcklNPaOkaOJa4LycduYG1RVG+kqPln1UvzXcEvnfiEH+h
Ga/+VGeZjYBNs8FvDf4VcjVfAnO43ji6Mlu3M84t7ofYy3T9Fbh3Y5gLuI4WeZuPAjzMi7aIDrX7
cfUkMr+mVBcdhFAGic7dunzUCVPZx2Cv+Tc6U3K/0lrbQEcadmBb2ZLcT7GexdtA5q6gFWdFOXWv
AfdfshvMD8klg6GZa5HD5idlpMoHEi+TDfvvkpUS9dQHtUavNhIAXtrf9sk6FVvo36rVmzdGHgJl
z5I3Ab5g3Q/1EDLImClf+G13XOTqLCNgJYyX64zu0c0glrIHrxv2Q/CvTcC3lXdakmJ066EhD2ls
gjcqjqBxpqB0k8kDqg1/TkdS8jZ4F4TQh3Ss+68G+VMmMYpUGBf+QtWi4UwkNSz8tJ/DAOefRsoM
qqtGmoom8vk2F9Qe/jEpClmePeUuU0SNDi4Xq6juC6t0YcRUpzM40oBYvfXlLgzxfeFwvUncIA8b
zbPKJV7rwCb05s8gPQxRXqq8fUNPWhSpsXb8GJT+DQkxLU/wDEjqwxhaQ2QsnS8Q7w/+P0n7c4Vh
D2Vi4fvpQWm6HXMglLpWdHgJBMM5ge9H7eftFzx767fUkA1iTha7ixKOpAx3gJcYI9uuirYb5RUL
i19UqSFKYDwSZtDQTPiB82d6hVQQCA7Qne8z0yxpcNgyjKmzXafVdIwBlsJwJeoM54Hw3rGxAPjo
KeS6YHQg1JMHorWoGmcRTmdZEIQC4Gzsn8aYYzXK7a8n1KhhYJVidN63S1Fxqon4WWtRpwZDYjsH
Q18+cqi4bvgjiIpfC7HhVLl/y/jw7Aocuyek4DJm40wl57O7f98ESmwla0wa/TIxx5IHWyLV2Hy/
fUNClz64Nu24BHZ1souck2y8q0pL+3mlKdvSs9viNIxKd1ZjYo3oQkrigKNMYFsBSX68/gl0fzwC
EL6b61uN/JSV/IpzHY0CMSHajWTvnT1CUMfLEL2vDmIFEnfIrWbEbXqY0WPd+m9QH31kwL6qJqPx
xVW0VVXXBbMLfKJvQCILfezkcjw5uj7D5Y6VTiGPGtgmAluTFJucSXHvapffb9LPnvsdJ8AFjdbi
tHVBEhyGSYrSMESvFCT8fWANeIhwz3Qa/Yk8Y2gMEDjVv6h04ftDUsdSX7htoGtMmDEKfDwPdB7y
4G1HbzAcIz+MG6GctgBuB8L/Lo0P2MPPS5zTkKawz2PRxFwgbW4ibvnFHQqtv8nB3sHabOdjaqEl
EW51qBx8fraYzI13eZ/HPDeujx/yg4WShPNlLO44WhZFzkZREi9HpKBrlW5O6C6wgEfF2YtV6ky+
Jqs78qoDjZZHN9fcZNEOgpiBYbrVffIkjRGPI/GU7MSdaVVv7TVsmKeFph92eD404BpEwYa6Gh2x
+CrC6DvX8FOUu9+NSBszbh0vEhRSjlxsrkb+Qn1OvA+y+k0WIxAABJm8kQbhBoWF8Jx3ROXljjEJ
WCePuW1Ssgitki7GpWbKhvkBjOmd1pdy9LhJfur1I/7xskFccp379mZ25tyHJE7aeA1mNHJEEN9D
g+AZoC2V5wZy54Cyp7XqCOZ/Tt1hHYe8RvQ994fHAfSLVS8j19TS9ibiqrk7JHhx95Z/ny2CwOLQ
Cf7llA+MJDcevRP3BlBBl2dtez2UYxyVqq+h/nf0H2LCWEygrhyFeeSFKfpDSUN6AHrunKfKoKID
Ffrd6hkql42xx7ofjx/a3Vn/4K/whx17isVoZVRhnx3MRfqO1kmpUWbx0FdJcX8z+Zk/LsMdF+Tj
tmTTSacqJKJZhWa5/H0j0Imgezwwg1mAc+CWOXBS91TeUx0nuY2ZtDDjS+OkCiJcrs+PNjXoT9rj
3DnASKxTyWwpmD2bkZ/kv0YEsT3l93EvIXACYIEGksLfEkJaIxdo+dtMtGZyXpRJr7clCaA0wBPj
1zBUahXmK0RwZsFjF1y7CnX0zDwDLsGEOaBIR9jBQhmszFR7Gqgluh/ZlV4MpyYZn9Jyl59XeuwO
wk0XzGqHoOEItHeYxR6082a1nxrqywcD3/Q6Y7/1r3vNWV/ZnhTMDQSRlcqk+Vk6qfOujPkFUkbR
OjcEbnhea/oDwmqXthzrITg0BOsvHb9ApBkfz2aW+qqpixuDwlBLXoelqU/Ly3vI3aWKmJDOh3/0
YvrfxCRSrnbeZt+/ghRFSYV20KqlLA2S2ZwP309yQLxa7kMvRjXBNLTcdrhcMAXaE2aBOAv4npNc
bajcC9l5VWoUBQyXo92B8S0/a00XZdrOmIgmCORmuUJ4yBIT/jEePibsLWz+/Ww7AC+kBYP0+RO/
cQ3tAlWOaaiLInIcoFB7aNaJlTi3Ool9DlI+5qC15pTT8MQ5TyoEBzuxkeDUZcdwAjmRAPRS6umj
N/BNxQFjZmLjkmxEerOfRZwP2A7Y1FKc6mXTckXkVxZ5Gw5TqvbVIN7jWbxDSwuJDti1f8q/AdK+
ZvJ20zT4/qJ8z9KGaH0FrTUtmM9B0yPokUXKrqXcu+2TQ7Pyfqx9yYn+Vw4gorMKQrc0baD+W6cd
BpE7nXEZelGh/ZnJZyNSW+qjvzodXdbyYMVIYOcm60v4ibkxGUsuQC9gxBidUyFhDNmuLXP86R/U
2G12XXwzTp38zDNeufHVmHPxTirExDxwggxWY4gEgR28EAypBP9de0vr3Hb5NrxB/TwEa6gVKUuu
kHw4GRmjxfGpPTVR8Xfpww3tUOAT8qKQfsrsJWy4fx2XE4mzV9HYWHLLNH2AtozDbSXYwRS9a4WR
BQqH2YeZQ8GyRL7cQcTLte69gzZqc4a1njTEN7Xp0SCA1OJiXAVturgda4WJARGEOXgdUeSkg7Se
FM4HKCfTOwxlJYshxDlHHn6+QnLTl6c9TA5yO/Hqo+mciOV9bL/61rVXAldEMcZCQeao3+IZw4DQ
rCbINNQD19ExTxMbBa821xHR+LXFXefLFdhpCuyBWLxIiEv09kBQwND15Zb7DtbE/yYeJCeC6WvI
Wg9u3G2bu0GhyovOveOlJ2rg5sRVaLdoIWn6qCvQfblMhmZrS7pwqTjAftBeJeHeu17b3d/Z80C9
syzp1U5P6fY+bFb6lHusJSQmgQLsGXyHriQ3jUQfJAw74JXcwmnN2Zc7/7HQE7Bo9NwOHyXkEVPS
AJ5Fwp3N5zSBirnUNjNYu33br0QEw9wZwUpNRRi4ff9E04iqQ8QScPwMOkgVlb/1+zmyImbTKrn0
iVNuet8l27vqH2sqAvXer1XS3KHydWzDTFd1NU80hoero/rkYnViBIDQcaOB5pILaFeBFYjbys+s
MTqJF8jjW+C+IBDZbcSUM5HFW7MsZv4dTZVaz2G+qqlbYt9hY3GzVQeISdkKi5G9nxM2oQ4OLtO1
q0Mgu1AlXgqzpqD6tc3htZvCrbBg/hln4pOoi5kooGZaMb4DeYRNUpEkaH4i+0vJ5f3Ql/c1NVof
RcbYaKmUSwauNPFhWWY/CLISSu7MLwRDvGe+WBdb5LToX/+HXAmwzl5LN4KHQQsbh0Yz6CSuc6oi
6GNDWMRN0A0HiZKq/nEqE5FPW22sU8cjZqg85RC0DuJNAJmgdIqct+QUAJ9wCsjaP66yTOZTxF6y
eU/FdcaCcFrhDHHWfzqenmngg2qJmHjSZT1KQdze46iJ91E/pmt9juhYuZge+8hPGIBO25iqd86m
YzZsCK1qZ57/VVPhciinHE1yzuPq+L1ZLP+w+vf2jihYpipoYOAwwpiLRQfSm3okJjXoeOZf/5mR
tnxhy/Vm3zhu4Dp/PZhDUaWRhasxvF3Kob1FX7mb1RXyp/zR78QU2r6ZKUll2myUDhGxjvQJ208B
M/SJ7QVqTqQZOvAjTenI83dgP7eUpRERJFJIyW21J6iswXJAi3F09obv4zVpFIcxhBIcOi0RnUDW
Cs5Ks5HiJT/Afa/HFDYDA1/OYW4zpMkJF3igiJUL+1+tELEuIxUZuFbZyKmzGDr/gKjX6eDFMxUE
tH3/AGPbuTkJk85mpygpHEKQB1RzW+IYWFKC8+/s52gZiPgZ1N9qXXZNubMG9ZUe6VZN4pCm7g98
MM3s9sUFzLaB2B3aUIin426WhAbnj1U/raB7+Gs1k6VTUhQCaw3FE/j7FL3LnaI9Km+ydIfyzGgF
cjWHucsFLSM+BHmWdObHqQd6l/vlu4mtw+Y+wIvUe8oo9ffS6Fej+r9FLtZPJeF8G3X8plDTMrOn
Qx9Sf2x9zqa6ANI/0ZMKrQYRv6hADm/8GLB2wN7/NZ7Ek9gP22nOWGRxQw6f/a5gBZ2KJJooyaXr
FbCtPrMPQjZcqS26JEYZtiCWvH+UTeuaHzbtm4/FxGBjA9kv8RMs56sjLuKgKSRSwJr74W9B8DdE
6wB3f4mCViQdbaW3bb9h6Ee1+n4yfGxAsjD8yY4ohB8DuFW2J1e18IwnNHTFAmPa/mk6O3FeoJ6c
i/6L+DRQoaEKDgiOlcDn/ZXzWuDtZO7fioy9bnZNN1SnDJ5r9f95MCq8BI4HtqgZgFmfj3QXeiVJ
77OT/buakydvDQRPJbMpQ3NwdHIVe1IBDZLrUaMDcOFsik+bk57wpEk0JWSXxPuWDLcBGUHOxzkI
drIbMFDNgkvCEN6A5wdZyvblfrZqcEHRu1FIKlx1mdWc2g5K0KSRjCK32B2rlYe8b9fNvSUYS5oX
Zh9mUTZ5nGqgiaLIQSLlPy6N9yrGoYdhMm1zTsSoK5wQaO/GJ0+uz/BvW1asYh4nbCqVhr6P4stc
kLIUL0kDZkjyutuZeeE1va/ngpoShZLbp/Wok7FaQxqQO+UVmQSqCG3HD2huvo2uXIkTfgLNfAJR
o5V53QfRCJzLLXft17lIlBblWbR6a+d1JDGJParjNIELw7v48uSpDfg/cypTRK9tVIqXfM0bKDfk
+lluJhsbd0yOruRFzYeS0hcbroAcXwExlJr4r6a2rPh8B+bhT6GWtK4DnmaqXZ1E8I9U/koqe2mb
6Sa/AKIIvYYRUJkqk3btusMn5mh3TaiHxHWX2uAKGMvYDshYQJNys+Zr/i0QPpTQxPK8bd6jGDD6
QG31hQ8VH1tQYXN+W8L/AZZNF1qhEcvZJQ61Y1CduZitMwngAjVWvjsoir+pkKbkPMnkU7/t6MWg
n59fh5u9+iLI+VRDF0YdFxVi0m907bNoIV3Z7CA93fBhvNK+hDpTn0VlOh2KOZ85CLFVR3KLbgcc
dXoVEPfUmI5sqfw1O6C9rraae7aXvQy2A00Ydm6z39pdFYTuJ8UV0tNlJ3yvdN9NP7sCEGJ0VnWN
Ekgvie6Kg57nHSk3Ww1aZgc8sLU/4xTsfxOm6BRP3N0oLEhq2rm2w0QLIAB3/wwPUzfhSMZdFEdg
aOD35hBK1JF4D3kl45no0XfosWfIHjVnlzZhW2Ty1rPc9LPvi83rqrq435yVW0TvnYih7abql7kU
dpemk6D+zuZWNhT0kKbWEFXoQjrKHv3dPDAgAkWKDOrlvdfuxblHJ6c6ORlBaXQALnfmf0isdiKl
5GMdgzWNTpNiqRMO67KHrpW62ESzVgVogulszKDs503zXgDVKIm1B/kvG9MP3LIimg7ePc2GN46k
ek1IT35ocQqT6bxU5nzAXgnKZqAidIiqWJ616iTcOZ1tPHTRJsZHcwH/RietI8TNjMRLa3LNgW4r
0ceZHwXeKjOPb/J9rcvwrKwIuOq9bpRswA/emELpi9OCVgQ/aYYhmXG7dqENtIpQdy8JDhQ4Q9jP
5FuW8Ee9k+/Cg7AH5Cvw+qIKYzPrO0GqhJyx0+f1lKLss9egF4cy3E4J6U4KF5Vy/CxC8z+23ef7
ccCICfSGOe7G/3wAxrAqeT/1H8Emmf7VqA37v62dnh1bOKPM3hoQZ7aZ+IQfj3FMsp5UKQjTYiRX
vtyJ2R3VuUpbao+Qhnx5Q+CN2gDJ/LywtzkoxvlEcHiD3cRdKIOY0IxzPdLB2WVqxLUm1/7qfCYs
mjO8RJD+VskXL249ahKjUCQ2N9e6bNvJpLWy0X9kriugEjxhLo4zUgkr9rHjfC8HYtvJH8uP5FT9
FpTUBQjZtL2yE4ooYvDmuydPPPPMDIVRzOszKl9WSmfBhLEzh45pAMqx+XJC7RAi6t0fTuP7EC0z
vge9xqkoThOhZNn5aCIujfM42MWr1NX5nf44ntIMyifqriimT73Smva1BiTt67mRGxjZu6p8d8/L
8oG6oMT/yTz6P56gccHzSSC1Jkea7aMKOnQ2Xq9hQZCpjty1akLGwckhtNRkNaj3U1+7K6akU2y5
J7SMQqL3INy424ZKoyE9gJCS4Zn0bc/ABo1MYy5c6rnEl23Zjmx4t2YuBIwmHi0loJ+xA76zNGUv
hVR8yEhhxKXM9yUsaQbTNxKBm9zvOddnkd9mMEiYyuhLiY6+OAiorwDPswlwuBK8F2i40n+WbVju
qXp/eEZXhsJjLxLog/64Dm55mykDk9gqo1vxfcapdMkmkfD0IHe9R7M0Sp4RY215MPTqCssvNMvG
DU2Kp+/sBVOV+h7hT/EW4ZoyBfpdIOWSk7Qazj5abJ+pEmTliRfedQMHenS7vkLP3CgOZvS/5Zi4
HOKfLq5uUoI5V9MgbYI01eGaSmWURj+XkDjyaZ20XGd897u5La7xIyt2QKJGeBF3GYx2tANqAhIi
Fhxg87hg3miHO1FELH6i3xTE1LR08hTcyHzP5JnicJenSKYnreVtdJ2zg1JRz4eRuAv6TnAvaPNB
VD1Zl1qg/LKzdlfTlFNgiHuvhm8UBY3LT8ndehWnYbH9juXCYhHTh6aljukayUZVAI94c8do/8GH
Cu2qsvW4NxFiwQea4anVIF4+XGotUc8VWkWPRh6d//HBNuGBI+WCFtkrtwDDE/QF6whdRuD7i7Az
TAHUcZG9P6CPespS7t7batrls93ZW8y9r1PFBNpriGZXTMQEtCOvOdeSdkZU5yYs6AGkb1KrSeLl
1+QY0LZpag+509fj4e1sNVL5Dt0oJ3lL44qhFn1/alBS19X8FJKQgZBVN/nxhSMfzVWk648zYdJl
EExkQvCN8n9XFA+bB7CR6CVRMUHPeDKsS+ydfmix9AbtbQ9LLgyu/sLKvhH1c5fGTMseImwMKcrR
akgVf4mtvkYm9onG6MzTOOkR08OdctrQESYo/KWhpA3c4kEDLzv9nSKgquibJ0Jc9Stq6dM2i9En
FbjmzWjXR8sjAb4hM+kk7ICOwcLN3tWeY8cv61v5jII5YQOOyJbKnpNRnBc0H8o8DGM+NAQ4le/U
2qQ0UwSsot8RDsWgqHh16MuohcrG7ALmt+5fSyxRRZiry93AuKrI0Ds2SGQ78Aku99S2Q60X3vD3
Vo0aaAjx0+gvDFKfzKz+DANyvyQJ96SgC8+qDIGRz5LeSWyysQpriYKWGYtmYjbCPJ5fkbcrus4j
c1wFhF92vEfpkGir9+S4b/ADm+xnlIALBejBbOfMbGcBkkhwVVKz/WRA6xiFGIDYG2YBY2GhWbZc
7hO09J0CjA3wCCH5DsYTva0XK+yytr9fkWbwHBB3IBhPGwYBZHOB0OGVn2V5cXybvhTlokdDewWF
YotUcfVN2IuCqk/vZqgIFT524taRU1EjjPf5RUcRyCTGiDlkoShKlu43YpI938y//bEL4TKcXL/D
wwNVlL/f43M6iQgej2izPk2C2VEQCulxpnO179rrr1C0BjAStXy3ahaBC0ywR/mqaaZfs6ZblbsM
eVBJDewdViXstWMmq3mxjXos4rvyavNS8jhs5pVf5nT55Nm3/ZUV0j3+UKXeO4g4+Q410MtwoF/Y
oSe82V9VPObZltyFGSOrhksJdtLggGdkRR8f2V7hSbvo6phSaDMZn0WD9p4R0jEg/AzWnEbe48kr
whxj8HV2svMT/5bh05NcOsQmZx4HMuQzSUAh6OHNnTAPiv4uUOpgW7L6k1HGCWVo9Y2TDwC3n5FG
t7RsiZJGcl5yPECKAanJ8ZFJudeNoTGM0EZUbdIhoL4zaUBsTbmbiAiK6FSdcnZ7qHypygi1/ekv
GsjseKT8FAeKPrEkGeZ7Yo99a/Ou7zqXGJ0shzP8l0zMd/ekR1ibPINkV2BAV5RkHoj/6gERboqF
BVxqpnlx+DsldaF3l3Zw0Yo40Ax96r3+a/9lmj5l/DVVV/4NfC89fpqEBfCiEW8hDkST5OMJp9RX
uhiprQEA/LhnkuSfKPNZuvlacu6+JnHr1TrmWxZLTXDGHV/QnH8sX+QDo7RAUOboty+vBD+dQg3Q
Fd5NyY06xmhNfsjKy536S+h5wViV/3XSLmpMkbAPG6RM1Ht2BbZO59TFGj4uSHSdOk6vl8lnxkRq
jeDzGe4KJqBbB/ZFWaBUoH/53FDfNl9WXE1NPBq6bGgPVmR+CiPLM8dfpoXBFyuFo7b9KS1VXOwF
mOSzLM1nEzFo/7476m0VBFa5KGZS6u2Wn1jILZJjafW4c/16wb8GFLyijY+okBVIZFh03TxZB4hy
SHna1lPBRLMELhRUMna54TBTNR59XaAgx2aZOFwuck20F/Xtm6GP0vHphnbcGB/Ft+VpXtxNnOhe
SV7umtGBCMUGX4zDZzG9iheG/n1NwxQiVnan9i+8rjHezg7IlIL/awodeS9VyxU5y9HIZeMbxp1v
n2wde/FgPv0sSqsuo2tCaZZhIrTC64eGv/r5f9CdVtgiif15jd7IaySfQ2XZ+t5hPvmRpFUtcdkO
OuAPYYbabTasdh4he60j3kcU8FavbQSSM00Cb49ibEHpTqidNLDWw/sHdniyvUu2cgJ16LPqIfZ/
hxGfovxXYV6DMUt8AL977YrwDo05ih0s8aYjFbCh7WPNu2f1MTlk6wot5mlk9QIymTQ2ynmutto/
wqCBVB6GJ9UB6RgB5e/64GOEqEDOQvUeUhcdUzzkG40l/gbJ1cGnUfOoErXjJeCXfQxvG7K49zkP
NTn95690dgBZqOKCti2quYi4iAt5S/MStWQbN/L7mOVpUi767rVCGoTCT77Tr5RJTP/hFIU7xbpy
qnZ7VzSg0N5canJobxQxjXa4Gy34KLBoWPPAtkkzjOEqAvm4Ukz5Lb0uNDUPuPxyLKGVTXFrb5W1
LIIEQKKn07W682s1L/zBiC/bCazJRGx28e6gVufjv/oTYAowF/NorvIXfxsbLUGuAg5kB6T8qp0k
RGCKHCePo4ulJVeHCnOoHEiqjEp6t198fDEBqKsbW8kKgbz9SNI1NtwTQ6efQnWTMkhd5p1INqog
hNLB/Bv3Wr7vrXMd8d7IJV10tbP1p4JyzUJZ8LvKeZ+iTKEUwXhcisZ8XzmXLQuFZ/R1ZDnBoqc6
zX0FlRN9dqEmcs5HdTXRWkHpx+I2OBMmKWNdf+oby7ZSTaFtJ3Ds/QHLOf6cS43fF+H6DUuoEN+w
deM4QqMugLu8Scful0Sce97OonLHOVX94d1Jbn97HFDwLlQvsXbKtjR3dzevKQHb3utwR2VLlR9Q
xXMLGsLZTN7b9i3M3Im+mDVteHC7qnhZrw/O4xdUq/ArjaR6a9V3daG0Lej+895e39gC9Fd+cOgS
4FduEivNA6lZKd0KHF2mGd20XwaB9kI/A3ipjis+FI1wadO1Y2a7lsN5G7ZO84mCHuSUKoZy68lp
3aJ1ZmUbAuXMcz2uHf4z3kZqXFE5TTCvVHfF7DA+iM6nNeTDNlc0UojV4IkhAKNdfzcYSGIX2hkE
WVSaVAplHxtVIumJQlbCg9GzOzuZ17G5h4LweSbMQ0eJSsvbOXU3NxGzPHPsPRSAuw4XEThKPlYG
SIMg6RE6HGNIL9pm+l+NN0L8c8n0slGDApSwnWq/Nc7/kq2FaZa9SiU/1UVot76ycfAgc+fEfxP+
3s8/Ux+Fws5ZqzefhSoFqAruPc2Bvh7mQR6QGXdG1MSLw0Lg3KWdcGs8l9T0ewQVzC+Uv0LrzhG6
qxh4Apjr/m/kswShSq7Rs7HZlPYTUePwFuWFV4HPk9CL7ai52Jl/Zaifwroq+kmpLaO9kIl8TO2u
oE85seQ0MC8Fpv8nEby7/UGQpuoJCcuRODoUwNHGPFucK0z6f/iGPvVF9YHF9+lsfmRQ3cMk3/f/
a5j1TOpwoFa1cJIznLl5r6hiBrWg/gQDfrnFFrlp1C+Q852HNEqKY7vnlA1vRdHhwzZhTBNX1HCw
IXrTejY8Qj4c88bGwY9uuO9ktwB+9jl9nB1tKM+oU6a3vR2KSr/SGWaJz0o9xSCsEz5gZm5/PZ3x
9Br6j6KfsAdYChyqGxELYbdnxfnqbqBFgp8YV4XO2SPIsNVWuSgANVdoztH0g8+RwI4xV7vcCv0t
2WaW9FEWZ9BjihWkSPROQ2DjdmBOyxYafTe39yd+9rlevGoMYAkqFspDaxu5GUxmppWNS5Ut+vU2
NZMZSBmyh/wIKXG46doE7uesGYJahA6NEu8pwvdKiDlx6iF6nD0PbfCMfjRBRhEkny0O+5NotU0Z
l+QqMCZMpzOoPWnyineM0vjtowc5b93swXkUikmWUSgHYNz37QKDSTMcpYyA+x2hiQ8xqDH+VXsW
VSpgqaOFCDiwj4BPHLr6rrYig8H5GwyOANs8IUVLbLL1wWcKC5gpawDRqckiVFBOlPo0b1EWN4Lq
HfLnFBfd1R3++ezFqrlg7y15UBkx7vE5w6gdoMwFasoIHB2vTQx/bjQG4A2eE63a1sDb7mZFDecc
GPcSQRZi7zgyIOcXygkqgVWbdI/y9Swf8w5o8aMq4s2w5jLa82NKZ3cqEN/dF2SeWkvzTpHnIye9
v0aH2fsXuJDes9ycVK+Xcv8DUIdwKj1MIYE9pCNoEfZMFhFEFBHGDUqvWevs9AfQBJpF7wZ0vavd
pXBWxjeqpK1X0iacoz9Wjj4T1YuHtA7jXy07Bt04+1pJwCNf1gGL5/+/dxKQ/9+8QUuMNnhzc+S7
wEjnSCYGShQE7TkSsf7s+jI1OlE8MkPqBT5BMzrslYTZnsBU943P1EIJ1f2W4kjwi1Vw23i9Smbw
wNBsktev+vU4c6ejYy5XLcCkN+FLmsfSYSF3hByJoUQ0gvk/DQWLSDb+hSHZ+4PKrpjpwEuuVQLN
whrKt5W4ZAa6bs7Rw/4UcaRN+yHJ0U/v2XZy89cQ3UKeKD6rEC5294btXgIGZ7/Q4mjLvYITD2vG
mmMQWLXz2rASVGXvnD4ec8CZTNiZSRFipuN153EhiyoOR3Pdj5H/XfyW5ASiYjOaRBs4sbwbd1Zn
cXzwp5Rb3B2rlNsUFTJarexZLBgNt4jj9IJFnSMHST7SMi2uVaC+u5TpEYaL8Mzr+nSbLXpsy96j
JHIFNgUFP0LN7lvSeCtVLIJEKs6dU169rvc7j4QGqEpXVqv85XYns3+5W8VZNUsHYiJ09ULndPhe
PSIzvvJIqJB5HKe3JLx7sfDLMB6UiH0PAmRi+HlfdKh7U58VrNAVXkIv6adjsW0vJcpl8ivaE4YP
EtI1LTNCbU2coXA7wu5C9pfwbj0iVG7Rfu5m/Msm3QrlAJ9+j50rwfC8hTJQZcQC/SG1idUm5Wmk
RtwhSgmu66l8dZO2RZtGNeBfBGHketIeAmqmWBXmuOd6nk3mJv8paDPK9WE3fggBjP8Yyc4KATgP
ClRQLRQICo2PS0tyZ1EqIigxsNWpOqk04MbCvzpMKEDLB/oGspHEiaq3N9tjLJ3MwXQoZ+Omyt2h
tbitqVsu3Y/q/NLh4GFuDylW3eKRsh82mKhLbZXtkTsn/uV8AIBWkS6eo0ZJ3/DiYkjXXSLTP9yi
EYN5DhLYGgTnksCLMKIPiUquv435/6l2O5t6h4p6mku2QFKYJ7CJ+PskgwC07n+R4NjjINpHU6q3
ztSD7NKcQUWpZeNm/nfRc8JdGmCX/nTWzExAEOyxwk1yo02fGyCR3sNngB7yBxwbfoPf2zfddEnT
s5SuQNqsnX+ffwxb3KN+gB0sWAYxHo4BmkY27xyJrmy+9EbDmt+G2ujAW7phBLCU2HxClvNNqPUA
YzC/oymosfYlfLreukeZQUfwoy6v2ScknvJyjRD9igOnukQ6Pb++//hp66FUdF56Oxfs/2I/93UQ
ktORsmTRRDoEqu0XPbzY0K+fhtrTJxsKteC7iYeQ0akgyGYex2e5lxTEQ86QgVkN33gzo7/y5yh7
kBMqr/W2Au6xQwxCBqfJXOqaZ0PrmLlSshfa69wrWxrWkuGAwi76Xq3PPbSpKsX/ujCORvfEEeHk
JHjDy4V85feWjSEOHAuwJObIETaubQAyi9AhG2AInueiftSHWIBUwZbK6NiyCBIfUgJT+qkv6i43
3NXqbuVFOzWYFYWJCa5mSYDLbXwRW5KXXzksrp5BldcT2nDPyn6HIY3aRVD++MKSyrO8FBjIw9KB
w464BJ2JQFI7ztYxTz/oVS4BGEH/zj4p9sthdwpzlMDH8k0ZXHxq4d6f1F007I0UMX29swb0A4td
+fhG63/WIZLnH774K+Y51TCFS+U7smMVUmhuB5w+nFQHXISeMwZDsEbwrju1rFNrDza0ZD24kVNG
s1UM0jWBgwu/SjjoiIgMC9u+dI3WTOAthLB/pQq47mvIAX5+0qYNG6j51qaRGB3H8qFYCOtzB1Pc
GkSi2dO8Gk6+4z5ZdvWT/erb30T54+Fz85OvtzkKSaiTPXDojbKQXVVF+N4Ic5L4klfzSatcOmBx
f+buhFHVzp35raTVf/cJI1NwIwp7YBexe0nJ6wcYWmdAK3pVKLT02OvWey3r1lLgThn1ioggWxAc
PHQ9xttV6jvtF1Q6voOJBC/0uidq+xRLAvTHUnDqfxuAMfBj+7QWLbPcZI2quLGNAhMueEkTP0EI
cBOvQmd1Asr79/brKYaVZCJTJojRtOp3CSFiRXbmAEb9etT23ZTWCxTsfxG+1eYly7OlFwV3+/JC
p2ccspbdfX6/vf/EY82Aa4CPLuaBRHx4/yoNTJD1tWs3q7NGkVzGx6frZnK336ms65aUHcEcSgEe
+yNXuT92yZ+6EaTTTuGygOmkitIg9s5SAGbnJfVqyhqM9aC7EHjNXNGHYtHPPmB0bJKibm6kN/wz
GIzCC62XpDDGGcjU10yFz28EWnCHA9UCrOkeRfJujz1FR7Tvj/HJanlFxZ6sO9QnhdZ9N4HUtx+t
5DM/kWHIzmsgr0D0FNlvN+e5FQlkCeB9VldSiRGBB8gDYjyonhnBsLHpgB/ZA5th83ukaWlSMKoW
tof59xmvIwv/nIiUgm/gpSg1tD5CQnXUtSvER3XVFqhFaxpS6SeGWlpdMxCZvyuGge2mh3EwzQDC
D3btOWQFEV2KTulKRSA7R9CdmuBstFOn1ENNcKqBxrWffKcuOmPVyRP32QgJz/9BYZ2tiFpkvUU5
YcbO/zM4Cb3U3R85uHb9TsqVprtu6rimkAj6uR5gDDGC/YWjDRhyTBOmHx6DI5xV6UlJv7mJEfL4
YSN8hVaPXeZYv66PmyreefZ0iPgQnTPm+Eypy2OG8nSgqyP14/eKW4CAF3vUTZJYXW+UbyveuZ/6
zqK8aIkW85I0diDabqSC9lwKttRBiFW7wZKZbrrgWrUkP9lHN819MPjvQ0alvFOyYjLMMRB9fGHB
dXLNbEaNRl5hFhAXESaLob5UXLNcyK7PO6usnZvvN7e755WnWnuxoTCJh3A5GThRbj7C8s8KSu/0
u+LmxSk89xr/QE3TWlebnTYj9KsNrNlHcvwr22CXspz0NzPiKOlzlb/uRv8fcwnh7UqCioUwLmuE
Um1dkOel9a8a+Gt3RHDB0AMV/W0lekf1ZIiqgXZb0p7/3Xob/WX7RQ0vZz6W5OeKvcBgqn1DYuUH
8eMdvl9m5nTgXbCEu3Q4W9MTxkQg8Pwf5pRZSBMTd7wMuoRKND55eiOC4P1GWDK92kw88sxBYUPb
rEK2yXwf/hYpSynnXnQLrcaC27hA9bZ0NJU9l3phqf926Oah4w/KzdgUiT7Wyg7uf28133glqtlC
IIN72MzW6RvVJbugi3moYTDZht/P49tfPu0Z5owdZAvY68IZ4mkPpCe3JogL7VfbeE0hGgdsHURJ
184hoThMcH+VeHh14eFmhtwgY9pTcnfq0F0bOTsdHYhURSWobsq6xXhSawTZGAuEMJBYHVdnG1+f
eAx442M4j8KhmDxI001UOoMOBKOngw/pdLwXe0UHRLl+fPYPtyvCxWv2nVDg46gter1GMOZMFNUI
JYbfF7B4xlLgt8+eIiHUeur2UEy47Bet7aMxDaUMe4rkyL0SsENO2m72xXgAPQYgTkbJ6NFbqke2
Iudzsrspr9yxflH/KmFpZpF0Rw35ltDA/DzlXVlDXz3dwddvUQOUM9ZUcFAVUmkdYueBZYbQd0qv
Dnog2B8cpOAz67MBYbvfJMTmbQHmOhgCccw4AT/fZLYAwp01cjk3NvZtJMQoYNEfRvHMEnycD4IG
FIUko2POmf43RMyK4phV3CjD/eHDwO+tfO7Fno3qKwqtz9QHT89p7mH9q5QIWmAoaalTFz0u2D68
Dq2ijWV+mOBsi8wpUvSDvbA/NEMUSaw8jRR7gM40gFB4EQHYtD4UEKVQH9g4mx76d+D57yDtpmTb
zD/YhS9rC0yrh/FoQ9LqqQxf3m9VMsYVOY4yfnQh/x0Q0675a3vQ9Z+F8HfnGteR5Yxn4W0fWb5x
NFW9Ufc/o7Wpvj1StyWIbSgKuUAYywl3rv8y+mygiLlOxrR0nmhWlr5OIdLU+yj9GjIzLpx8Zq9H
LuDW4QjTkjfC4Y66HOFDhjiDUlX0kvXEe2CQNcQWt5co+HbfeNaAoRQfTeMmMUc/pJlH9GpdsDOC
quonfL7u6e6KcK3wbi43BkMPRPy7Bu+BF9cKWS8ykcYDoJ/GnfiShcn/R09qrCdrD1hC1FcnEwaR
NNRRTECCw3txjWFCR1GVyXKjjZGfi3N+459EsM9tZoheiZCACpNd1hoJZ/6Wvl55L4tfoHngG1zl
73XfvZHCvwUBSleVo5Lt7InFBGLw9orZAOSYEwSI5Jw6v3n33KysQ5u7/kx6RtYzQUVTWOz6BvVy
CypjHq4F4eSlbgZSH0YgofgocMNA+XXg0oAGkGO7BYDnlIqMG2+YfIu72CX+Km0YdW6tY9Nhxc2o
U5C6fOh/3qtzZkXDdfbWTp8vN97nw6HUNMInFXyX87t+EpuS5VGPV1iqU21Pj0sPP3LINgnhacVO
IiAguO67hySOHawe/bkyUwLYtZEpPnGZPGWJkbBtGdLknFzLRKhm8OmG2RUGb/NL5FJFOf8wXECl
IE6l33gZx01XGcQGem6WvnO4OYGNRE9VQmezxNTEakEIsNLJCynb5KICRQ2M6H2GA6XWjlhCGZqf
PRXvIdnnGfSTzhYd/By5Idy7ghK2GGKjDaqnFQtw/NSuvTQxXLE0uMQIiY7RbPwaJBtCySy0ZiAj
2OO6WBUvlLl7c7ucDOT6yDnQkdDAS9GYmx/7HBNvxApCUeVgup9W3iwEOkKxuO9IturMlUMF7Zr9
EPf/yITVaGpOpuwex7+oicxwHdDuJCNFjoWX0heTS3fi3SIhmEEvUSQdAI+i2dJPAY7q5/noRojq
ukYsnczff/3QdOeo6FqiKbNOfU+213MXd6OZoxmO/4uUb6KrJBSNJV+aiIY5It6l9zuFh0v5Wjc2
Sh3u6IR9qoYy8lk2SCWMuPkDspFxFq2Bnpie9ZoisogmIR9n1VClYl1o8u2WKzv5F335bvoYGqhp
PtIKalpP3ANA2Ul1rIYfuQG2+BbZo7MWydoEqsEHJAe+ghmpC1v7huaoUS4rKKG1vG7vv8KcGr9b
TPX/gzVRZr4e0KEsegFhJmJvdfbWRzLgyfvprr1A3fnqja6ejrwI0/7UPAtyI76qEWt3M35qFyQm
t12ze9i9MYU0173eyH7lfh3nTJP9PDco5p8jdBPEmbhTuJ28EHKfRRTq0rrNIduxMdCL5ZDUiUj/
w6rqCnMjoP/QihkTHuQy9jsLaEbR7tXjxbvqMXwK/2pAdESwxJQm6XyPGA6hGlaLEgcvKNNvGE82
ifBWHgZZ8lnM54pIfQm6h5pJPhNqoAgPh0EFLKxME5H6d4mvdl4E2EnuJSPi4lrW47nwr/17GfOr
ZLv6bH+bJ3lUpbAIVaLPe+CNUMYIQDhwIhqpKOTjXOlM3+lQJiouS/qOsAYi5tBhShobqBQ7d7/Q
rK+4I99Frl/HWI5I61c4Nxzrp0lpbYWbRsFySMJ+y2JWfDZBYthSI9/wQKdR66d/oTPyZOPX46hj
BbylDOW+omQB461of7dGAHbVvR3CFJLEdyo3Zv2oweE7CgovK9SnJagjUADDOQWsq+K7v2juPxmo
XMnIh/NbgvJgDdGX/e+xqnLOV+x5UBEt80Uc1Lunsj8HBGMeyn7lWWFT4t+ANRAo+lKnSNyHgfbS
IGCNRjeXUxLQCI8M217QMsuPkvQH2fN5oCwgp4gpWmVPFB+Q4CmYlG6XoIhhUNQZaB1ah3Gmb4o4
dRK9Drka3axyPN7nh0qw1IlJcFSbyVzpS+HfTTxDy7XtMUwWcTPgrpgrW+eX67TE0j5xibNhyV3M
xYTsrjDoO2/hyG+gUNr4nGEd+j9J5j3v+/Rol8iSX7M5RETdvl+9Mln6vwHxmiXssdprZxavtKp8
trWa8YUI3HJre09nhY0OAxGU+mU15ZyzE2GXwVDtQDOkPpLblk90LjZHgvPu2a+rZXtkSgwCYbkN
NzHW2o5cHMRgugtNSfi1176nv7QyKJpZGFKwvJJseSEBzfbfueF2OkUAwS5zkCL9QYpEjaor2c5A
JV/93cZGEt2UjraKaturbGte061QKSu+8i5JS66UH3mlLIzW+TA0WSwq0SpNEztVc7eqZijGgQ/q
zrDog8Dvj6i2okHY42x7oSJ+XgPVX9Ef8AE3089Uv0+Ky2bXC2gLo8R3eUXJf6oZCvKZSzfgF0rR
1P0nEGq0cnMAx4wncVt48VUuCic7n2wDphWunmAT3bA6bAX66pWz5pEn2IJVzZSC3X+RyHxoLtnr
z7JE4XdOvErtFTkJZ7G+z1/4SHqHPYWRUJqUyjAeTdnfY/ExYXAG7u3nXkgOQbw1WIZyqNb9r40+
4EkGOBPvQsg+mRqJ1hnYPW8+LKcFnIT+2vqxgirU/m2AX7yGuBhdj0znuhp4SHLwuBTIaGvTj0Yh
IsFO60nNtp/ImHLEdXOS/YjK0kwOMrs1pEb1QvwdzcbwBvcOp67uJB5FoQnm7kd4ULTffKDFdg26
hphNB5H5M/F0c6GKD3npqdaI+xgtqjQHBBf1iBde1fcWUovyELHMv7+Hz/viZqoHJFN4OX5fmC+k
U9zTA2duxI5XzPUCRMXquCzTjhtQ/KRMbgMgMeQ5l6Mix/HhYU+tWjcJfwZR++OZpCRV04J7llxd
vea6U343jlh7R5v81ZNzHZvqPamN+/uZvwW4aSSlnxBWncebjYVSI9NWeSbX5SLgKoSoB4IQZ45p
NXKvxiMJzZ/BKvRILcKM+QDe6IUc9jctBAkhs6BaHgnLwsO2bMH2D5LE91zGfmKQAfwI/iUA1vhc
BPCYRmyVcx+E4NJlkb5uQQJF/qMC40JB0PfpfRSkdCksnYZV6HTV2c2Ia1pkz21+/MVRQuqB5Jmy
Um1kP6tVhtfzttiih7SqP2Si1cWkLQTZtrtmFITQ9lfcYlBagsQNIZsngEB/nj8NEvqT8/5D1H5f
SVOgsR6i+gjru7RtGDYufccimhnmYuw6FApZdn/vNHLAf/ox0mKhqf335zqJmz6AmiAxGsj5j+SB
Ie2Km8iyNlScwL7HekeBvstufcOp6OvmYSPRLUXretv9qiN51KNKnNa1XIOP5ac7q3QchyuzMojt
awaGHcoskZangHyHJXa4dYXtVCG6fx0FxH6z1yNVWGEcZzuc3MIsjsPbOyZGxdB8So8bU7lW94C2
uf39hvCzg18S63lfErqvG/1AV7oqT0TmU3IMWB9XntslfdZpEje8mNMx1fD5wXdnH8khC0iGel/y
SZGYx9kR9+dWJc7caDMw21JmT1r80tllHbMQa5/+Kmyp0Cpir+3EISVmOU0h2VrviKaI5Me0kdwo
NV3hZceph5FogcJTELYpfTJtZ0EX3RIcvt+9MqgrFdaglgUc6fZcrgA/5lTB6uiX7/WS+xPsqMJR
n4IddAcMsbcJVBFrbwDhKAFH+o7fGtb8Jpyc8xzHrAxE3i3LBqJ2xnG+TOFDvmNGFLaHOshWy6Hb
Ml/mIVV0tQ8gzMfs9hLiy8+Y9AzXwWLj3TRA/Io1IXenMWU7mLQhnEGcVL+Dy+PU2K2MTeDvzI74
G/K+r0k9Wvaz55vwvQXE76nefUDMCNlkgefTL1iC2at88iT+R1mIqyUuq101mvPKyCYdj4s4G/cY
1rhb7B0/kDELu3qk7871K6GBhflj30rIb375B4wpaS7dqORkA2hwl1xx7xcU8DwiFgNZYnaXE1Ln
nZvMnKHHjBNf6W71GPBbobZq4eJTJT+duT74S5pwTu6xQphxHx+1EegDQxi/ULFVChgvfqdgAvhX
oDNcD/uxWh0Ok99YAuLmR9owALwa8PYIY18nyYR/l2I7zI1hh1STzRplNrXVQ9KUK8NC5nPyAwwT
wuDbxAKxjxdwHqk4yPrpTOBpziZJYtgJP4VOqryv539XzCialw6Q9wgMcRnqeF2E98P/wUj8FpCG
W9mrpdSwuN3H/8KfaazC1YpXNLmiR8JaH/2Cy90xA/kkJqQISKsoWMLMoY7Gcj/oDqFoiyQcWRi0
Bk6nSLPtEreTOE4rU8locdFbc7lNLeip9NvX2cAuZSs7bc6MA265fM8sNFDVDNvMkROV1kwq3nNb
1BEwNCBlQDlGq9axC63Kl+zXNAo4zhU3YsoFmNSpL93hjx3f4N3avqUgGZqHQQAQdqGEzqjIr7PC
U/bsfkTj5v4Ln1Eu8vqcYT9+wJYwQtgEZ3XJggq8qukcHKQVp1tHvta40Hs22EZA8I4MSdPjBthX
/YMFSopTHviwtPpVead0jjYyCvpdNlHgQUFRrDBePvogdbCUBxrrBFrlZkkmnYOR2Ij+QMaMDKW3
8xJ9yOOysceG6xh0vzBIqiHvvU/5WNbqXujBeylNpe1zb2WCLWNkIuFhdw4X+qla0m8uVKz7Tepf
c+zxdeAnXZ+BW/m4yUH45n4tFDLyL82DeNVUZEBGlNuwFEYxCh5pvfx2+EosnYWGfVIHoVmvVlQO
Cl+FPNXfNgNADLOMrCZ0ifg656LIXJo8R0HIN3pjbbFMOG334c03x5H5cG7OfYamdCutD0BoQbEN
eKEeG1dpEDdtBpG4Kx5sogXsP4HWB+iITI3Go+MTs5yr3mpHN5G4Aa97zDK94Lvc+ZWSyhj3EZlR
kzLnVFK17LTNvMVA8CPBOcKXlsa4fcv+MaNJBw+xEih0yLWGcVW9kwY0+CJSH7ArQeUa6MeBbZxq
2nee1RTP1TpFqmyVD55USD8GnBvmevroOxIZnZD1i5EfuJinTsYECg19D5EO0iorNV7F5NSOpKU+
k9Fh74JSLxCu+lXthZvDzMXZ7dwQDaNZrjjAuniRrZD1Q4rAPBYNjVco6ZLY/GY258wyedmfz50k
91JqfPGtfC8FEimBWo/lMBvavGN23eNOU0ErlGqYAcS5kjHyp2Qdsab0Woz0mJ6civg7PS6OBb44
GjVPWDHeFVB+yEzMyEtvjmf5o/R5X5r0Aao+S8GJREfXTD0q1DRmgevO1ohwKvIm+bvkBSoc5n/N
d7pPDxzkSupR1fYZ6DLuuFWxTpGbhvIcF09OUP6/jIC/EykYCypf9ZERTs0J2gmvCj4ijd4JJnpH
gHsH+d+ISzjT52RSt3mkX4NdOYPbiIG5acSHF5s3nVkgvVP1e5BFVCdz2YL3zTZ9CL0pbcshlJxD
cjnReL8L31B8JXQEWVBFU9N0IqBZ4Lc97Z3VdwjRxGcg85w8QFmseNQ22P0znTsomV+5XVzbxS59
FDaQuP1jS8moewnyZp0F3L/+CDMguOilJt+0/gLo7ZjJ5T1QboEh+s1J7h02iUiLn6Ozb60maWfR
vuSt6HUGXu3BphAfeIEeYslBi8Sjols4vjuOrq90VXBdur3uzjsDenDunLEy462efcNQH9rqgCWI
qu4jmlYhkvmCW2TepBhatWsiyhtj1lhOuEAE/NtnlMEYb3/wKeOx5PVg3Ik+5QFTZEIwGwqIyr9F
DNjvaXlrMbEkDxlbsYin0rgmUhxEE/42B0Ky5bA980sSMOnD7acnV8JndLhqcz6ET2ivLZl1dYbE
++MRAoB+2gHFXvTSlGQt+hRqxuxehnah2fqtnI+qYLnvfYDVcAha7OmMZk224leV1i6DmdZoX4jM
yYLn6Anlz7+NuR3t5wuucNZncpteMI3zR68t3xknQEU/Q/jsXQzJErJnry27/n5HwQFp4Rm3aRSE
5zko7Tbt5ikkV8dVl90UZ9gAe2H+94ZWGX7GOMQaWydVvcFiRZEPKg/dIrgrVDv7JfTdJMXVjsd0
6REXN5wQWdK0AATP90rFe7zRTZWWoX2W/DTiZP1c5oMrNknjazgx94M8ED9gS6B+vv9LfUvCZyCJ
GvJy2MFse1j4Pa/zhPRQvPzBdG4UJNE7Y3yCwh8jYaELfggEv3/l8+aTp4b2ywcpAgqA6sR3USiB
gtPcr9M7+Ce1WdbOzKjKMcZg25AJWoHc/vNOjD1KbCdFEoYnmoqSP9TGfivjcMu/yUXyNfA2Vk3e
7ySktwlwmklHJxjqpRXMvOHlFqMFHp2FQHR9tCG1hPEHCUPgiC+tsdYjF6gLVdYOIkU9OBnuVZeg
08yy2h8M8A0QylcAiiQJbh8LcrB3ZmgBjnJ3MwnsiyRo776dzNzRdyBDnJt96d8WbTQDtJGS8YKB
JSv9xpJKuKfgpy635fNt+N75umVsDKfs/W9OAnWVYeZ3sfEGGiTgr0v6pSbw8s/6UwKHApxBIg6X
7jL17Iz8xh6ytIiXJhREo0MbQDl5A4zk23SvSL7rLbMe4uVp3APYISYftFywKEiSeCTqyPOkRAdq
uHMgJzO7l6vvNJ6bUUs15hdpN7MgQ+hPKonhuNSP8lK9kScIb20UxCdWGtfFf4sGkkv9bz6FQqRp
BvRLpkZfd7uqnqmCLFQl/G+Xrs7uWNhghykOl2DzPRmM3nm9S/10c7CaLvq9fNchnqk/u2b5suG8
3C5D5e3c4pQUTUlTmqxbGlQ16y8sd7iuUhb0p/rWxjKTC6k6rlS4qg6cn1BaB5uKlmwrPI029Mdq
oVVpyUEyf5RgKJOlH29wI3zCAIDjm3ZH0b4Kl141sMi7Y4TqeEjtGqsMSZpeg6BFFY8WJsXbbB6F
snSXOK+Ba+HRHk5T3/rNgA3uvxsPOCP7zBgMzr6dMsz2xDZSApgt0dEG55SI3gamOOeqUOQolLok
23Lk2s47B31+X4erK7P95KhdWPTiW693EP8ZsvYGbVdQvpLJjeh7ML+6L11NwyoOTM3Hpbb3JOqC
g7pmilEQ9pwDF0rZAyhzptWL5+EKsf8xf3NdPcG00Cp1Lx35kDHGPIfy2CSpB9FasSRwYdYPNXrF
JHWod5/+0CeyfHwo00jh9ez2xKNmIVAwETZgKMVyjDUK8cAXMqPSFXppJ6Qy537+meaGTKfLLprv
h7ItldQFNUe4RVweM6aw8gLuiVdMZUbET/ILbwRBn+ty/MLsIu0zFh58Fw/Y7o88z8qhg4hNQsHO
3WtMlWdOSgI78CD3AgYgjWIVwDdc/7tiBl+AncwSyWGvs8T090A4FY1a3Pci8vFjBH5ou80KlhRx
WR7NToJayIiFAMkv8lKqsRD4/779PhCYYJdq3eFXX8ltHcOL6cAgjmHy/6AwPzDOuF3EH+R+JHkk
3s9EBW6flhEdJ14RpMCOrJFpJb8STNu94rTsydtj4vogUiatBKbKkf9Rv0yYxginQyTufuaZQsTK
ywUfePM+/RjKV2zByyLJGEh8o/OMl+zi9O+Iu7OUJQxvNfCH/PJEAqnjx3kpuAaJDIPQ2gS2u+wB
UQuRTbQFN2j44yS1VPkP868PdvsRRjjGubiCsB5DgP8t+yd0UDwsYp6Yf14m15D06r5nQk2lgQ4Y
d9va2CoOTSfoz2rJtkLU5hxhaBN2FN5AZziNp6zOm+kqxe6FruZ9B+sEm9OvJoUUWfJbASRDJGpw
Oj4xVJj0JIFBrqDIzZ6/O9l1GGNgLNQOrj8oboaYwz7llPxK6Pzf7S+VXnzxbneMhXHsmI7jeHC+
HVvVGG9dOPsGJZ+YBbo8rEDvUV+0uHu8FcUbgbWejm7RrAkmz0QyZilMZH9aBMaeeEasQZg66EyI
LkstqLKECBlxvEZG0LuwwiJHnBiwY3jrM11L9Olvlpru0jkrJvBZFDax6cT9fU0B33qBRK9Xp9Bb
/X7wTcgT6hx3jd16Hz94r6iigumfWw1mw38pjtafDh8WU0lzlcqF0SbWiyjXO0es+y15qlJvTNJb
Xg4BQ0BUNLpOPNHn44y7gbYHuLqL18SWYwT0x8Cwo155DURrq7xMQCkLXQn6vf3TMaylP062qvJY
niFXw3Zvjq089S7tjP24nrZR4IgB6Z7JS2m2ZGvXD0s6nvlczT5vzHrVoGPWq07P66XThesiHePp
n5IxhTHNPMcvugE6eeWpG2yeR61NFlW15kKJEdCivlsGUiKKMKQuxyrUP9cVY4fooCKunwIUXWr9
ZVGZm/XBp8iijSL41R9RzCzP4So6K4528v/NzGpeSz5xr8VncOh/pQuPsuo74YaokhrN73hQ71NA
6Mahe+ox2p6WziGHYgPEvXuyJh9iQ7eMnpYI/w2yy4D3dRSotTBYinnDO+9PwRR4+qIo94Myz5KM
AjxfuutEHTa1Wu/6M+vntPBghGlWE19/HXjGoF6hXZdhaRrJTz60pIpDGEg0GAbr+A7xedvrdmTi
UiYBZaYiHrQg0Csn7fwcu7SJ71sQn+iDvMDuqBN3sK96DJomgx9eV8hAkZW85hAz9D0vTNc2H64t
mx/IYGCBjJ1htvvb30N/L7RJxI/MjFXpgEbRs8xN1gETXY4Qt4o5w0yQFtSwMeAKBjGMR6HcE5oL
6ZgtRUbE153+CpAPKq08tDkX1izKAP2brF3IHom0mIv/hbULmBJcs3ICyHJAfmk7mmSxHtjIsz5Q
rcEZS/d05VdLPro+QeK2ovY4mxcnPBoJd5Q8iXdsjX/CZcWx9rHRiH56o8vYwIsekwe7iREW51/Y
O5rG1ps1oPqPlY3EYKB/Rn4FnI2cZzLyOeDYCHXyBa5nnCB6V9kDhf9ap44BONsTIvv7x4OzzxhA
D/J4LD0kiCE3RwpPOOa/Zfh9Z8KG4Gf1IS/ZRVCwDw9CF8DHYI9a8rLlFbBj4Y67+htVkZgEAU4e
dFFlc2Eg4YUhaRNJRg1S6QVS4HzszPMNki/pzjF89aBLmGmUfYzjPsI7b16lLPr0/nNyeKNJru+9
YXjTElDENu5avJr+PaRVi+GVd6Kqdl+SmBzEDsa2GXUkwU2F0PgCR2/5O9XxL/2oXOalq4F+JSsj
lw7Evpx9Jd5OlyIyX1ZXC/r+rE6huoOjr3H7RHU18fW2b5ZAX+oS8p3teFYKGeJuHNaM/4iQ7nTq
Zc++htpcTOs7kz0JYUCdU1kf2bZKqm2b1/CROx2eGpfuTvnkM86BHE/ldIDW2o/yz6tVntsocxUM
yqCHPDAO6IB5pgmLELeUjHMPhS06xtpMHxFYBEII7RBIeU0bf03iqkD5agqqyzRwSETx9tdxQmCS
E15Ov7ah/tjNeBRyHRetWRzyWgPNvdTUOFqDOMI0Vkw1HxiGoNf/O4buT9ZTR2JxXWUUyFYK1t0M
5/vEZc9DC9Auwex2ZbSNnsEgY+e22ykj1aEV1qzJiqkPEvKeiS9gdWgcSuA09GOkePqD4/X6ZxJM
TdjefCS5OK4kr4jNXF8lJHlZjcoCAXVjNJIBSZ4X+8gpbqxcdOETUxpmN7scGgRhKoVumq6l1JIV
8jjVYDijbsWfT0POGWxdoa7gQGSEkPONrVOKs9vXCOKZMqrix18a5Za56vhBB2sc82cAe4r3FBdH
p+j7cIt+3yYONeDIgnpqkZA+bUJ8m3cgUXsNYaw/trnjrNRsVtGtxiQz8zjA37X3ZGa8nX8oXIKd
tsMuTl/Y+mk5H5B14r1muYfwzDqc4q0dAaapo8rnk97atfYotsKwI8PtgzS0ecH3EByIGoKsHxrF
RhbhOajFIeosgEeCIEhhraSnPQitMr99IX1+Oe66ySSo9EhEXyBpUaGHRrA1OxBODRRwDWD+2hM5
4L+cu+VKwp8sYp8V9QNtc/prHm35vxLvy8dZnTU1dnzLGve0o7BDwO3e6On75ZD4KucPIbUsakSG
TYxEb6e2VAJGyuKoeQoRF4T8YlxnZMtQAx523xy6pbzsKxgMFEnJFWtKIMP7eW3SyYgIfQus2fPk
RwTFUrC2KDPUVXagari8Kg47LQ7COtaI5KDov6Qz3TDQskJPxE3VHpVoZAslHB+cKu3JFevF83RU
x6TnHkJv+Gr2H/UIItl9v0pTrwSirozffzyUw0FX7HdeyrIqwP0TuacDNN+fsNX+NPh69iHWRvbI
3ol+NuSRpZX2aLXXr8sgW25okWAMZ61pDZwiW+VXNWforD1prC6w3SE1mO4BR+6YmXq9eZch+Sny
cKnjbm9Y8c8UG/MmSdVVqWRZj333uCZAYKpi4LDPvdtlKoubvZRStQNkISRI+MYgx+EWuZTFjn4D
PwPSe2HgrqM1IKwBfLjXljFvZVBBa+M6ZPyXc+5lAA/xjwGQ0wVRDmlSItzR/WMM4vIr73Xv+/Xj
p8tOHRAYsnqnpiMIUgI/ZFv5iSP43/iLJ4Ipzt4DuZrF9HqOZ3/YiADl+GG3q1kF0GrhJSjiqk1N
wg8bjYJlZMDVzk3R17Dp3Dxc13n2edP0GVTTTFYnq7E/GYOwSUQUQk89OBie15c1EYIS3jBK3zt1
f1jxCU2y/P4dXdeGXv3oddWU3LNfEy5cZORiu/GFDD5Dnt4/OTYjJt2UpgRfTTS+3Kua1CDhaIew
Q4HRnP1Y1rLHSKiGx3WNVIyNE2OxWSKfIQ1qNzNFci0TE9dzAxyzkHQc1q/1YeJbnpi4eFRT6JxA
IASsbxpgbnw6SATdBX8GgGTayDqHLvF9TpYHwy/CrLbgg+86S95F7Hnjw/Y8nJW+IKbFFCK/0k9j
LvNzkyEbgkVnFUI15EwHHfGcMQiwLKnUA+oI1bIVQRVd++qbKNFHo/FCtvFWXpcjZPYgBR9iM6wD
yiZOeXfuhuFKPjf+fyCzd/uvUV4qe9M+0FoB/2kDvorFWgn6w4diAZXJdUl+/Xf4yXNdr8kVa/mR
pBrrFZ7476tjyUrFF9QwSDoTx2xjuckJPO8nwATu1V6F3L1Y2yX/KYOENwQccDrs03XrwShhle8e
HuW7dBzUBrDzpoCtwgXFSFgibP/VhQt566kRyPhhIMRf1pMIttQkmVVrnUB/Fr7mc2hgoQKv/bvs
xdu90zzSGIfyVUlck5RldWLMfGie6Gekg7ITubxYi0hknRgIf+QsNQB6R1Hy4h+P3CKQ5meYM1Yl
qq7I3tqhiu8gRC9CfpfaxU891IpqYDc40xxBtTuazV1ID7FsNtVQTHf+uMHk0SxKp/w6BAay6Fw0
UiuI7GT5PSJHRln5IsqOBDNhWiuztwg0UxoQeN1MMXlx5xzLOylC+oAFUTDPJXWZfo8BFO6DrJ3t
u+wryphHB+z71j4N2Alex20tc0cOBlyVeBl6UgdiTZhwZNeCMHeukRqvGHW09sbCMjDR8Z46PJrA
IZxK2AFikwxg9l1XZzGavdRnCqFKtFBgvEbdSJYMJEBPZfOHyDJCagcWdTsCce3TeDhhMPE5ZpLD
Mqs8/dkCF9m7zlwqMn9GjgTr5+LI8QCkcEfxUgj2/RI+bA86xujw2YxrzrPtI+uMg0esmmah+9r7
9x8okvhVj49A0rP7ViN+e7BV0Ngl5LJf6dL4z+hfvxUcbA2EPZ+pAa7W9CtORNSM2lMUBV+ZtoZS
6x9KFIDol4jy+cflQOf09+8o85UfXbDrRV0DJ9lvP/slSjbUlJLLZ8xVvWMDdcP/aIBWrj41kE+l
XsFH0fL870UoqRUoHttfVJNuLhxtP6cgz9zjHqp+Dv6i+XWEC0PUMuUFfgZkdK4UgC9uAXgsNls/
oA1UYq6tpm3sQhOMT7dC1DXoqHdSE1mv4qdCD3sc6D/5M5IfJuYSKCfk1Iiwdk4ud7l3o68WkjXL
D9FsF9njfLMIoDhP9k0YJj2Xlt+C2yiMDWrPEL917ZoHPvfjSZ5cMqzQvaOL+vj5ifWkAvQxpoIh
NlCLsoXSzNF2fOKfWNFBUvvrPkDYH6vDbaPc/ZjRREs4DaIYzEqke56VDKrAE8jflDzxhY16zJ3o
gBAfNpS6sdA7Qq9+RDDjd2CO2RX2uGX3PCNvEfWDLB1CFN9JttX/uUyGmC8UcKsEcqYQU57QfmkR
CWtf+WsL5hTNDpvZr7/kRHm3cGEjmfqP2uXnjxwiC2yVhFoMHno6UjeE6huvrI8y2gHSYSb2mAzu
2JxZ+puqP4VYla7a4oNymhnRnk7LOCXOhuW+M11HPL4Hivl/Nu5R0tO5Ha4sJYuF9fryW7rekB4R
I7hGLPb3EFVYH5z+Rl4YS1189Yy2ABJ7x9+KnKOMnEBOsNhEm4oSAhTPNbuUp9gHBgXCylmE4Scu
rzAXxvezli4k9h3VQkz0wenffOwXFg5DFc3mQ1mX9ICn2+3vPg1G+HxMTVUWTuedl21lKlw3rMmS
y3HJo4XJ4QEOooqJZjNOOax0EGaKjyUYCcSKxVe5hS3oRheo1MZcnhaBE6HOhRv1Mgvw8lpJQ9Rx
ZxVcmj0Itk9px4ecgpkPCGfmQR+IaMZB7xNfPAjskDU1t9dpDl+MXDAHWXTn3utqrYuKpYYoDMjS
sGf3WvnpqwvgNRh5XUjIWS0a9F+nVS/mweZm3isUGSxsXuMdYGg3hGBEcEdDJ5TYKxZl3O4szKe5
2S0aPXZBoMJKUtlsDwKRKXWOjshVsRaVY22i7Kt5xeE3cqdCN/qgBLy4dyEdBQohLhE9lENiQ0nS
qo3XQggUD9wgMOLNZJokpK8Fb/EmeF+H7ahFtnH17CQWMB1yK/l7X7C7kD57F6MvWn7dxGJNjxzV
u6oBBj95BXAJVwUpP544rcIH4QsrQuZS+rbeW+V25YYSPFYQSvSlvs3Txe4KHzihJ7aP2tqX3y9I
/+s0rkVZNwGXoEXxcIvxFbJUJ/NtgrCm2V4iGOJEz4C4g3V80p/OYPWVm+n67UQrQaqKs9gLV1LE
2S00Ka2Sv8qoj8lEl+4aAgG1+TA8/Ozy4crBok1tluYxu0ibcJ73UXUOKboK5kKLfmUgcP1NL+pB
bJsXLNVe6rTlNq1nw+j1iGm7SDWpYUGVStJ+Nn9ZfQanAB5tU70eyr/uIz8wvP6E1tX04R+Rnrfc
zut8fpPIuh91bhn2PVl08IhL2G6odIZOZXklhdl6YwKgcMh8sUTXbOlv2UYZJKKdbx9bMB9znDDI
DYTkeT2JxYqv8lLHF2PNhk0UcD5n13zO8ki1RqK+Wjijo+DVqpkn2D7YOQAvOmN4dNlEdOsEQpxV
ouB8HE2Bu0RPX72M49fwLlkqIDw2dnrQuczakYbTnsip6FWtNSNN1n5gmQs3itHFuwyOAUmg0Am8
rsphNfRtoD9lYZT00zIdkjOS5BbrGgZxa02uVYlfi8sfhISLCmHBEA/HrjVCjV0/5D75z1O3fhT1
1mMPAScdg1yLbzTiAY+MCvPGjqFYxC+oUe3UvILEGkbdMfNO696hRgxGgLxQbgpNdVqcBScSt2qb
xXRhIjudwOJUpwJH/1w58fQHR01UQR3qPc3auz7iyIOW69mo+Z88yW8ODk7otitqLOV32VL2WQoV
M9+CK9KRNv/z/e87APNDNrDYR/AzYHBNpocgqqYUkkHf7F88LIzTubnNYDXL0fziMhas4ZY7y3dR
1b06zVHsQinKAVq2NeKVvjSM64aL1kVtDRcnxbvGSbHpupq/sSVPYJg6YGV0F+NkLp4E5C8Oem2v
ySBRjUELHqsTRNiHKrGer7QyZXQVeLn7Y6mWJG1Yk7u3bDFwdMdroy5QA36qxh2UDbyeMYHnPhEO
Ceqi8+5d76f89QhZ/PNjjkxinX3FyjlEMDjE6zZeJfSMrlh7p+L+nbzXYMlMFd3Pw+RExE65Lwyc
Dyv6Kh0Ta5eEonvvP3vBcKQVGUGlGdsxwtivdiqdAgRGR/vQNwqrp6o3gY5vbODUugW8a89wfNsn
3oMOvWn/4Jrja/w+mFHUuEew/jGVPA53ct/lbj9eH5rkCUpMonpmykLE3Gns1VwlioBU7dw+3M7m
HznN1PLu8SHh7ENYHuCrzg1K16if/sZUXDlvCeZTNbrC6n5dEkSz1IbzNC1cUcqcylMkNezOyjcv
eUw8zYf56BhGdAqKaI/CZgidOY14yht5oxrqo351R1eY4c93gnPclTcI6Bvu/M4gybQ/+XnBXfrP
XE4Wc/pQxfCCaP8INQ2EB+wPw4UTdi56FduBzBuL5EXh/h+ONdbHGYC34F9HU9VeiKAqA9Tacb7n
JzjeD6ZnbIXinEd5hTkJad4qxw5LI+P8czGpvaYxlL5r5EB3Tj9G6feLw3Hn+/f5iTolO27+/13h
6JdFgyyphegCp+HiGs7IuisxESy/WuklenuKllrOkv/Fn5xJty+KCDYOLzr0r9igNCyEJMQBozGT
dcCQaGSf4uDUIeYeDcv4SWyXo1L0IMbby716KYvPm1WIFC8zn/LZVpONPZMQ/eZA185TmRpNFBsG
PblUE2i5VmwDwVhy8FH8P44JoCBM0gZ5I5uQ9SRuqErMhHLfqMdl1QFoAEeqdnGH5HcNGrPjxeKb
sw+9+MbNbwNFH5p7MClURBpZYxDqtG6ZXvh8BrV3sqmlJUQbPXitKh1Z9hfl+hmYvGNu2JW/i40v
Kunolfc3fgNQKrJXwbVvena2Q6Tb1Q38n1ZwssyXbkj0/xu0xKb/q2TSqLNt0es3K+dYdN8adn7P
gHSuIJcQ4Xyh6u1FhFmRs56X3hs6fEQB3UGzh05k5zpAPz8Ese6niRAOP1lVngRQ5S1xsTpkk8yY
Hj/dAbWm3oHzcohlnG9FUlWBo9btW+57oAnWNYcm48Xcp/yovfnJX2BO1RLb65gT6bSTNIydyFUS
nABtbGdYSSuE32bRjEyZahTnkrotwFD64upUbNhVq2K2IWL9gQ9tt/RivSdDNbl78SKQoQmHcRVX
/epfIp309aNJ+/2JKZy23NYz0QuoRr4Ix8K+G2EErBxWztVQPqOFUkkD/KqVV5H9w6pYHL7JraR/
YhHP8XVy5uisp9ThStObJVOzIltSDBUjMjxTMPazuRq9iahTwJ4GtrhR8icAJI/tPnATXzi/aPBY
ZBn5YALb/qezsFdgaUx5xJsum8FxX1s8HW0lJ+p8XxXWkuAkrolU7boX9LQJoXRlnBZccayLef6h
ggL09SQyO8LyIjgCNNWja1uKBzAkWQS19gtdedsQSu97MuwEaMogWKUfxLLbLMgESB1GzA7+tWq3
dAQGmxSraSJ1xetNgGucYPq1CZwzjx6xURFP1iqtBRYEKFjfA+qxR52lTZ5EiMosMC4MxfeGcB6T
TVJdSqcKYz3Anl+DcWtHim6aJTZgpYKKVbJkn9pAOsZGfza6b+L3uhpshyJ85TG+jvEMGewZQqW5
kjBS53fbsrrgho1ZqLTSahrWZcpf4q2wLko4BdthrmVvUd/7xOmmDWWOPuYPTQiG455+KwcJptG2
CrbvIOheXsYVYrS4eA2jQDcre4FrKgGTC6Sus0Gyjut5aIw2cRlGxLCGOjvpLPewKKamyQ2PsQPv
ff+zXert+JkMrEpNxh79HkMKLzsW/Ux1YYAeuLsTx1JQq5xfAs5jVvRwjEV6V/9yG5YrR0wR92Ie
83PYyXWyToExKIi0rq9ATOzW7Nh8QfEP9JG9TsYgm/v1ogw9mckXLMAakXdKtpRVEAN0I7CQS/F2
e0CdduTR94FqpmQYaX7EXteMNEN5P1sHl4pUZcPVv+auZZST7ewSWvGWu4FnR0HoEzykByRS3kIL
ragPMoULU+/PjXLIMT72wHA1ajHSufqyOu3Ip+mOY9Y4frHCcY8qcNYNL7yLgro7K60owxZdD+Ff
qLIF4NYNs4ESBCIsMlRdYs6PYSSdIiOEpwFvkY1cx5c7UakWvyUchCOuYGIWmqF3+Je4WG+CcaFy
4FmEQrx+FKJwxsnxFyxP9fUs44z/YFxbXGqY4NUfgiv9gxLdJvu3gfyD3BiEOfkSId+qZTNQsxLp
IHLpWz6Wzv1t4tz6nII2BpxNLwlsK+OmMMXjFNVZVppyzhEiq2fBF774eanfoanK40EoWuHlcHay
CtHg+M9rmvMVPSQGFn6nCEJ0mUD8oHmjeGkQkgpeWVp6WSAdUQJtH12DBxgBrm6UMpPzl+J6fwyK
r5py7B45VUXJ97N/t1R929vNtw3r3pRuRvobT+1q/4uzoo0hxxrkUu/3mCSPRHM1Ra762zKy+Wve
TIpBY6uekOIkHEY9W/OeoGPGwMpGY4bQOBDBHqRJrzrTO3ziEiwHQzBKXfW7xtnhpCWVvXZg/Wu9
fw0XOpmXnLGCoC3So+svLejbmIgaNV0TW5BBsa5TINvWqHQtJ/JMSmJPJbpDmpZmRbSb76PRlN6L
ShYuyx5IHbxeXW+OBxkrYcRIE7zNv3r45e/LbjOqPJWm9uAPISDXzfZ2kGG87cXmuOTcPUFCwGY9
jbaGwXZRycjsYUmrpK4TM/4bt1RJlEoNKRKPV0n32249X/6r8YpUbtCYbc3/jOodW5QJrX7MXLgR
KHE8wY4nCqs/2wwk0E0piHDnTtzR7XBvsf3JYvtyypMeXgh9pXeNOqkXNtbIS4sDeGeIAdPDauuV
9/A5BN58J/aWklAtz4ij7iDXZwXQ72Kb+aa0X5frUarpmTiR/d3ClaDSjtPpZ0qtBj7QN/mFDXup
sF7hy0xcKnnup23a7oewkBlCl38j6/zAC36ipYN3raZN6HZ6IV4nYsSMRRG3h9DCf45BZZuYQYe1
ESN9kCSk+9Vo4rGIfbSF6WLIjJM0jSvFZ5ld4jRdeT3+TWk9OwntqcM3bYW2sKNaRtni5tzIp/qv
1ixVREKWIzSZJBxK5nN5UYEXXX0yPIEjZ5uFOFhYFaw2GJySMxvbXywcFF+KUvMP4X2s47FpRPcO
H+oAGrQQAvIahDeOagvt7DF0NIvljFB8xWs7EtLkLtpDvyDDpu456otX4lTUVGE6elc2VHkgFinR
K7oY+0knIEqDilRswkSdhMx2iVyvH0elGOntFu/r64pMaKodyzANq50Nd+QIGpXzZOZbXoI4l0lu
0DE7/JjVGJB+Kyc/G4RE3ngbWFCWMaJrnj3MI1tDwFf7QO74CPL8cMwfAtlG+ugv95x9tPeDPUgF
crfZwiisKFcnEQF5gdNFObXXK2NMRQgDoBEgvtWseqQ2YiFbry9oNqlxNvIuB9yeS5459KHsqMu+
bxPX2Oy6Io1mMY/LsoCv6TeJaf8rW/y8rzSiZM3wrMxWgu0xC5zb7C6Mu2uJG5Odz3+I8ugsV9ES
FQXVlcRXVtbT/NU7jUANUViz9pMjBtaAg5JITx0xj2takTwhtj1CH4QpoQoeM5iSmvvzQVwVTuNd
khw7eJVIDNZGk/aLhZukPMWFbaHl1nc0euDV16dWkAHEnGgwqsVvnE93B3iFhTmVu64mR1KsE95y
TXIcf/t95m4ajTArWrRKzDolyYr6VYyODuTi1StxhPekJRKvw3iUr5a1g9LwYyVS17G8biBHOwGz
em4HpH5VLE9LDh1qaHCLA0Y1m4S/tWSdLRB47oBj/Q1HVSZGtU6xer7hVc/lcnNYZVuJStuyoUkg
wcdkLAvPPRZAUPIIOQj/qUID3jzZncAj5/GH0yrsxn1g+95dnDhvi1VF86EZ0yPhiVqiGgQu1Vmb
fTkk2advNYtltmlhZpTgjezmsj1FJwLD7NW+IJmAg/YpBSsECi4xyropjbBoVXM/qMlKkL5FwFeP
sdcKS3qcPym9+qUxeJWlK7dB4hryicjgJUJJUEHwVCQlk1GXO6dODShxzWSei1fvUbRIO/GpLeHK
CnOQwjar0jiK69sIHYEW8zackZr9a6JppL3y8PW28zl0sCHRraLp89QjyjeAod1kjmy/q3zMaVEz
/H7cn6FOPHTfLTU2toRn4Stud6LcRjD2o99B0Qt3BY29vfj2hmpqFJ22rNfEsV9yYDTiRPV4bDtn
UejX8VzscxMsmvYz6E2BcsIIVC0daDHErir4ETR9G8QP7O2s9SDW7LB2aqGwe8zYylUmgaK9E36+
rsFWQvDQivtkL+s57lmOQmXere/pHAUK6nCFOiftvC1YpxEDnFgox3zf+lpQ5/wB6BRhbPhN7txZ
Iebx8E4nqn7m89vsbLej+rYvDsaFanga2OTHVzSf2JvEviKnerbteeAvNXefCA46N+1SikcJjLw2
fUqH2DETD9G01ZhWaU/dBONeqph7AUYJfO8nl3c+p3LDmBdUwJsVVzP+xZ34QQo+Yi6k9On+1kTn
nGmb6sSJJLaBMuMiJ4brUSWKZ5/C5Ne1su2rAns8CQQjI7f4shJSi6xrRhQnJJmxT/yagUhFIFPH
Dk46dsNA0LZs9GS50QNIc6lpgqpMZ19SsiWXEID4lZrOcpKYupMicDsK86bRQ8B+ZRDkRS/QIQR5
pga4QaRYGPiPsWx27mUzZNUnbpIlSqm2QaJBoZmIrAUvW+MLeLdRU/evDFAg2MshvqaYgk5H3DI/
gT3IHpP30iVo0BRhOvMXMHzQ97HOtIfr/ryvIXef1r6XB3rABe3bR3p5Os4blTlsRUeOLEcuH35Z
SCo6P7fsvJz2TLVRI6EqZYPhhW7lRyevbMIMO7Fm6e5PSXx/vkcpO71j8iR3Pdr9k6Fk7gtxT/C4
M/v0mQz5SIU+7NnqP078544iH9iegkpPAY2IhzbnZ+JRsdtZzieS8RbQG9qzflXY50O1hAnzeR94
lhJ1mGMS7dF/mabrTwvE0LwWKFXOCokw/e6IhPNV72wmgvcYnSUsYW65+BVV+2EInIicTRHJpuXi
p5o908mWodBScjRNDkwVQk9pJ3ZxoawF0tdgnBatImVZ3cMPci+K8pJHoddgExhH2d5vePr+gBe4
P0jpFfj9YUDA4CxQ3qpfZHP2gjBWzYb2KxBXfUKHuDIf9vmHk6+Q2i4VPMZHkLAHNAPF7WGn8dDt
1pkge6EI2q9U/vMc8ZLWHaPMpcLwPbXmq4350HggqAF60CfOijC9fhIrohquOsZ9MSivonbYdfo7
TSqMNL4c3pgYA/PTR6F0drdwp1BHKbw6Ui6+7auhPfwTF5cNL8UKSUHU2650xp3fGYLxO97psBak
JvRckLJuX6PXHPTLW3g4r5MdkWcCIz+zuhzXuWiyzI4fXDBkVTlocqM1cEThB2cg3890FWmZQyjv
PfAqHXuAQ083v/H1z8o6ab6l6zre1Ro8t132gkFd/7ZjCsFAvR6HEZRZ5Rn9sWjXrBJAj+CHkBuu
YtEd/YMVeVW5BHsTyvWeXPlIhqrqvuUyJQ4x21rnG4tDfvI/j6ket1VKZi/GCPCiVKZYwIvUJJOp
tGDjOHVfyQfv7A0NXKs0nujwRGKgBNeLQWTp57ARHP2qUXVirymWbB84rLwJqNDi6L5qGCYjiJV3
3FW8rVlrAsFYnq0vVXJWN0rS0HCqaZsAosL78/qXtSsCsYfMFB2gzcrWMJew7gmBb+FAe34e95l1
4yuQU9LgDh4kSxsIilM00TgTBLw8Vof9TL4KELrEfjw3uR/ntUc224ETwSR625CeYGqvXKttuGJL
tWYBk7Nebg5QXPGQrOLr1+NDkPylWiIPK5qHH7kkqvXdxDTAAKq23yiWmmtY73TFvHct+cnlHpFW
4Bf1D67SQLFU0NWfv2k8iKZWed/ndvjnhcSkODqyFfjepQcGBK/LNrPMDZ1QGatdCfSTBiw2DVSL
fXrDAWbb+LNywsYqh7kpNvjuDG9+tBlyqngIxtFwrP3UYFkMw9+xxatmp1O5vUV6FPlhrUkOvHQQ
RkMjl4JoXPPJrigKwx8jivwVbj8dx+msFXGmBk1mACZGvlcdmklFbdetnOokoBYlMjtw7QCF2qiA
CqpwIvI9BMIZpZ0tFfVdbj23ZtxTVDBibvmCkVRG4tXPNBKI6dZcgEHKGG/dfC5ML56kBro9f4LJ
4q0sHhqStKUN840KVsORBe84EvmaDi5mA1HOrRUEJQod8azqCI52fd/KWSBuQ1XzfsbnrWhsw4i+
vCQ8ZEf5krizffWTFs0Giiq+Iudhi4aiRoO+oTIsIl+ULI3YrU6qLBywPFiA03dIOfnYI36cUAHJ
ng2d3oKt7yvQoLsKptayIpQcXUcTLaS2c8AN4ihIPP1UDQIxt1v61tQLuARH7YKGYQssBDKRfvlE
suD4p0Leqk+IIPUjYspReMEi49TimV6RnU7hfzeuQyzQhhLa5hR5dZR4+b8xSbeXwtNef9ZEFGrF
ORMbcDXy+ZkVg18Tytnz03L56VTXFHQf1DKOCEU0r0FyB/fM4gSl5e2CPGvm37kCss30qu5YDDZu
mg/c3QQd9IZEl4BM2etfyJM7aHF6E70IQPwcjKznyc0fxP4/AD/k5Lekn6OVrXTgGwpzvlP8NMN4
ldD4ImuaR4JItXWpBAl7ruDrZb2gJmfRWx0qqDIQDALJKG0mY0m96bms1IFyjlckjIWTtzR7/E/Z
XLIupXdvV9DdCyXT0pPRExGSk+zoPANNYk23QZyiH7jFwOmJXXVw4GCyTTGDmmaXRUDQePWrCQhB
agaztzVc6Y+k9YI1y54Z7gtgRaIMPlTCdLTTDrNLIApuWltki+YocoQfQ7cQwt2huaaUhZ7T/W86
RVaU0QZR7l+lPRsHGUNL6Xp5gby9TbhaNJJJGtZAJTaM1C8QIPcfDd1Y0cpANE27LMZtqGEZ7BVF
mu9IoJUClHtqP+CWCgmE1JGa/Qb4rQ7LWpAQz2sHeUu8tbaZf5XY9O7zPS0+hxuveaQlLQwU+AWn
Ik/RckbQASPqiM5WQMlwWP3ptnxSLcmOxEStBXRJNLYwx5V842w3KX70b2cSXLOo/A5yzaTis+Sd
BmuYKHuC69/iGbJ2I8WxCOOk+YhHQddhcOQHaJ9f67ihrCFB5X/N67s2WnO8kmEnE4NHPF4WOUzO
pXm28rf4KLYBKuiw+9SiNlxWtq2C78eem0cHcX6QZdItYdyb3odFnlWdWSR6jKsiFIKGUFw7vcfs
cfbkXaaU+ZXZLjDDBrm2wrBqkatERUFQXZO+yDPHV2lKAXo2vUkGLKzpzWYZa0NkIFZxjn5piTCT
5pZj4KJqnbop00nTXoM4i20hdVVd83niLYqVr3d9P/JnH7yA9/y7VKh1RCavHHSIrqGjwLuVyQ/l
OlZn5nxzTpe7seCAMK7gxKLNC2OBX1jhueUbWg0p5zi2zisQ7S5eQfeHVjUUVd4WJ0L7ck+jpjFG
AS/Iw2wN8sJWkZj5MjED8TAi2XkBg9Bk5NdI+2vhO/y38TUoVxOpT/ssuW46J5HlIWXFEJNR9xqq
42kUlPnEcSSv/DJU1+0/VEBOaTzuQcTS0exRR4EZB6Z7qzh2WFOkYCywUTKEclQgt6ZxZui0dxtN
Vua8VtwKOqWlFUrmK7z4iR++AVXRsqspGWAh8q1JnCfLwux17iSlsLxmlbLZIMdSUD6ljffJ/SVt
nOqZEdqLxaw/T1tkj4oCe8QMbVEkIdTF6jfhnIwZUiCEP72be8uWrlknWA7fB/AKZnJ4OjqCgRyl
Yx3QwJ9AMWtzOcclKk4/Vsu0gwYm5QihFX6sPB2GQUCWhgXFVQQj86sUtc8/4VAq3GKMhqtmYWD1
MjYq3lyOERYA3mFyLc/J5BA6SO8zx3oA3HSR8pMaaMKVMaIJp0ayjw0mYbdPtp8wArtOuH4MC4l1
j6g75fMawJ0THl/pAVZEvZs6OTdDttyAFltnCKnWzNFqghwrkYOIcFpnFqulI6HNgrCm6LA2/bnz
lQ62A/WILgy07y8EacL2N7NHIn+3ZXEVUqA/mLeU6ahRHkAFnSSHBGPETn5kLMpIQGlYG3zMh4yO
x3nUE3Wh+9RPXGVfHLnB3qOi9uoNxYLNU5l5usFugkdiCvjv6avq8zZ6Xp3ddf/ltaOr4BeqsGpo
+aVHVzpEGP4aZpG+qE9OndWtJ5tJEJc9dtZyd+pdnMdaHu7lBpsNscCddyCnbM5IvNz7FEJJNeaW
5fag9sSdqAED4+fbuwILCMbe5B6GlzYXUIR4B807CWbMwHUhQAAFTb5Epw5uICD04h3Na5WcdRpk
9ZvQ3Hd3c6Mf/Y1vL05LUFgN8oho9LK6YWxeZbE0jtzoTanPe1RsrMD8oVuNQrGczm22aCuL7+RO
kZKfRvzoQtapy/dcD0Q56TUcl34TFLz3zfoZZYIxoN+xU1kdZN53cPkx+YGhGD6pHnKdhDKzWfrS
jlcpctcxVj5IhgAQTm2FI2nyHFLwNi2j7of0v66ZU2dR7bR8QJaL2CJrmtWn6qcvodWt/jI2fgRA
eKbkKO872+7jJqiOmeXM3YIpFTyGXfA5FD2rAJENCOAMp8ocSvhe4ae4qdWLA2VT6pfFlwcWp24f
fBpJP5N4mEF1k5+UkE+oxY1wBLQhTZ96vpx4sYrGe3jZNNleRWKn5qDQ93bTlmH9wRFgioT89RSA
q1QnZoBWT73SAEAXY1sC5pcmZDFkIxwovnl0+t5uuDdymmgEhjB//hkyUCuP5su1bVsuD3tJbboe
25Mp+QFd8v7hj4IcH0JrRAdkL2dy2uInXgaAZJ3o/LbbLY86FW+hkP5e8w1YegRga/X5Hk6KT4Iv
04YkR2LSGvtvqyFfhSCCTqeAAQW0O5CwcT6n8zG/g5TrPoIGctZc2R7Rm55FnZZnlSSGnMo00Zl0
SrtAT6UD5cyEmJSWEutDZfWiDGpFJNFFg9PouJNazJNDUyRWUtEwPoQxOhjZaNoGdoxE4bCNkNR4
I3zmUJMpYtkI31WdZZYtxPkgJEPw88/F4rliPDecNzjYac65C5cEPt7csvFzhLT/oqr7eT9ffdBx
eCjlBWMaF+G2jm8+eV5+a7xgKbIMyGlHPB6cYdUkPpJ+E7MwdWinWwcSUhDaiIF6JPigJmHnpJJI
5pXP+/d5r7O6nV185c9BXVVkjFALbesZ7CDwrLQQ6YZkuICKH/blWGLOwRJu59Njtt0wAz4d1mjC
okZ0vyYhQ7fQGvtv0ophEV6pCiWsgp5ZqxuZzkh71393XU/GEcSYRNZVv2uYuAKmNPG5TApp+0p0
9HLldwtVg7jjDAeRJQICpqfp2xSu8Hz0ic0ju5RSkUaAz+78AziWsTszGGUvppLYn0ri9m1ECM1M
R5wdX4cF5sfycccldzf7mNwbOo6l4VO0BXteTeg8FHC799uR7X0YJPTg42JLzeH0coY0vuuuXCQo
QQE6OgX/st7F7BalmhjSxTQ2JwX6D9Fl1GHGRfjk+oMmKHrjV6zaMrbo9AU+TXAm+Fneb7IjYyYJ
uawLQ20UqY3uzUsZfTSh9+He/a6vCpifQMnh/TpSTrdn8caRQiFbUOv7AJ2nEnCZnOjlUfYKpkac
QKXve7BvGlDuCk6iyClsoDMI72etw2TdFVcp0kFCW8CcPgpSZDxYb6c2nim+1yWd/vDrLq6xoTLt
agIAZICelYNGIuIBNCYOyN/7bkOXO8m6gva6su8Gv7qInBuMLnB1OUOWZugh8B+NT71Ff2W7WA1M
TXSNf1SAPHyfURh+wZeMKB6/4bBq0OIPOOF7NnvIWOeCXLSkoK3eokoqNTYCjwZ04iZ3LjoKMB6d
LvY2e1+iJjmmMsCbYtF9/kXSyKB/Ef1xHikjF0xWblZzQiqHjuktSHTqewhBfDjsACtjgKQ/ed8z
WpQl61Wr3+sLdbZ4OyF6/q3zRm9+eiyRA48ai8Jh26H/bUiD7hu0xdO1Dr+k9GGGeA6hHoMQupUC
BrMG6LMHdSK3f590kfclu6qARAiBS6KIwytEXoTttogV9dFHcWm/E0Ilt4+5N4ASPVgADZ4jlz4H
lGxf/Bzuav5J3NnEBDZ+Wh+/mCHWLoPimcABR85QBbQD5p4j/dhXWmcFFaAm8ynurQ62MvlB5HW2
IzByDmYLg8l4mcNZrZY9WR0DHCxVxgWpC9iQXF5qa2Yusx0QuVkvhEGBcFJh7qnFRORthI+w0Xft
4/LSaC1I5q3ZfNpKlVxTST8Bs1Sleg9gcY+EB/N/q/7i+cVvXwezIJufyYisVb8c3Gan5QGGQzvn
Dz/5QE++Vb24iafGsRSiph42MASVWPiGbvK4S2EdQk2YXS8yEeqdhgcr0Sid/8CwM2tsDIwy3V8B
dVsbYwnXz7Qh8uf4TbxH2gwrirkfbHTl0aTqQEzHYEObXhYbdBalvpFXxk4tKsGqqN/y9FmMe355
kSlObhLZ0PvW+domZO7xO1fZCsHG9Pr8IE5jheOBvJwDwyTJRjli+T0AZbZRW7dv4frshqM9v900
B3qAWxNKYn5f/YQp4VuDL+POXsI/ZGUwO2U9EpZcjY8TwTQZQwQ91L22gzZ3ZXraw50Sn1fpZkQ4
/9k9+Tj5RBqdIYrdUdq6qU4ZSywEdhwe/kCiye++mVaLmAvLrwERTJ1RsuzGDkbsWzO+biPRYawb
k83k0dIQUSYGmk97rBdlLrEIHu2Pt8DwyIC/cvHqpoyyeHemWAOlmiWzPFUJXL1pB2K1w2eyVyS8
Q+oo+shhmUWWJRt4QWnhd0PMY+3n9L19NN1yxYym81qASr22cAkw3kn947Jy4bESPPwWXY9V3irz
ub75Bqfz34jeKjaBC+3yAK8FequnrK8fkzghJDXtauoGK8xaHFsV2OLHSL7iR3y81C0bTs5oofZT
k3NlrucA3BVP4XJLwYNXk/nTjT89OJAxYuHws6gnXXPYKD5npfkmTCsgFDr597sy6cfKXBAyAQ3C
+7PZB57MD6kIbbVTzl/3ZtI9ey8H9IEb8dpyeU+xDfMQ5uIAJu3xQUO9j88NVPfa7tWiJk973T05
TZq0jAByvEZ+g3QAz81JOpQPZLX5/dBc9Y2JMnpD9tJ+PCikDfPkf70xkeWNSdxWY9+hlkks7cPI
aXYc4/zalpndU4Sq64MNNjk+R2Qusja/pkXDaLhDC8dUzDGhRCPTtz70xLSVfjugNA6VTeCSR2DU
4Q5iC82gWt0DesQ0bjH7uulwMrZcP7/aCZc4bCpuMVzaqUm11tzAVTDRhCIGvyXzLvX0w+pEip9u
M9cAo5B40auM6+shVsieovqCSFXx83ONW0EepcVmFcTGm3KTTJSpp9ZqqwUDCTEiMFx/JDE2aS2t
Oy7F8CrbaR4g9kFnuAlMSfzSCyexBBakXbwDsRilT2ufoPtodI0M7oENMJDGs1yarw7Wpqr1pWjl
tLXGo14+ISENozPXnxCBJR4KUhreYSTpLr/ESFUSLd18rMwOHaPHzNrLUpBZV+6I5yGyOXsmGm5A
sNQgMcgdtlyH9ORr4blW7sY8zZx3H2ZR7dylblP49IEKVjGd3erdlanxVe82WK5LTzEOCxbF6Rk2
FeyvPY+6JMdDZJw9RGV3Y2vIFyndvP2n0M4ndxbMww9eUszJt55lL4RIcc6mx0QTRpiF4ffAfzXq
cJ4Ou0NU7eLhmH48Vv+QyfZNnAPMmJao8oNrATBAQjap8Q9sRmETB5uoBZQ1ARsLGErLwYcqoU1A
xE4xY1GpqPDL9Cow21d1C+V0LgMbJehEogAkFU8EDdhFIC26nva15zFNNVHmmzYqa6PTyw0ie1B+
EZk26y0XT7i60CplCq0vzMM9c+XcT1CUrBOVglg9o1ghEHDOue/PAA/+NkfDlNpAW/esGuiaN6rb
GqWsNIpNqhnN4d+zMfeTNicMcqoSuToex0f53woQNDuBp4NHaSi4y0sJQk8lTHWVO93oDd+ttSkG
W7dor0HMU6d5NwD2/Cr8EyB8vpI7S3dqJrv571hmhYZK87w4eLhcsvTOGD1Y+3zfewlM7nvpqbBv
X1scBlD46ZoPhVy9gITnPXQSHEncji/ZpHHmdr4fziyEZy2oyrtlKrHknwE6gaasFWXnIxSHXv2a
bIFRKWl2aAOiWjVANEzsXAnFHHuO8/u4umcXhmatb1hYWh5NxOMGKyIgqRnTCwFqfNcASCWB6ns9
4uvhENuJA3XE5NVHbvjvXLJ2E6CHVWMV9saDIuS0FLX5XNJhsDJPpFvYz5751ZFqn/TB6/CzMcQU
JhaicFz3ODgSPNt/7CPKywWnt+WJ4bqfSYd02am8LH60ikPoRJy0qgS5E8EkldeZ2cKeB/rDBlFH
EADke3bYMErMfMMGoyONzNtYzNZSa3fVnEgmA/tMpX8n5ZvxDOc5HAC7rybAlY9h7F3MGOoEoEEi
x4Lva4CkYcdmNooqLd4ulO12PLoq8CxxLln2HD2V1JU49nU/iieb2K4+/l9VOjZEkUEa6LkVxy4M
wLzAbRrksLq/FsckmyzfJ5uuAgsmzryEw/zRRuCfkU37N7kYOVaPk/NivN624Twkuc6KbNZ6QMsp
eknjsEwW25to7Xvu6IU9QD6PyeW0HXt+VkqU7HazsgYM+reHKMI8VUKNckJJpk+ASQuba+uajrGz
FyMX2HGzD4Agx5VSauFunhPR/LhKuv1YDyBGBrmNRs0H1fwWIcb8Rnc+VAsJSOXfV9HbgFtMwQzD
YPAj13hXzRTviCs6tS7T7cRNHhD1homMOr5YOGV0kYEN7m6WCBtaGKfvPGzY32rcHiWHcH4D0Ik5
ySXnJ6sIN/yLytXovytkdhStgdT6UkyFDO1Y2xBRF9+ME0dDt1A3SIAAuVePji6jw8Mb2qLKUIKo
N19poM2oaV8q2+bfQHuKlgNh1TYOS7yymQmTe629SxoNJt+/0agyy8g9smJruY6kVf7FN3ViLR//
NfPy86ZjFfmrnpoZZzTAuf11slYmZBHgSG4JUHb+kaKIsF8ZXWRdIyzDE3Y0fgrFBj1aUz3R+C/l
bmGB1a6QTtUQCG+3VWitfgi0dksiCmCiHRjoaj9VPwnFk39KKQnOiWg6fzz7YWuDFSab6jcZoMj+
KxtWOuaIZg18hQ4oABLGu6aHx5+f8pyQH6LIeg0zzgBghw3aqmADOE/lR6jkAzXOKiNfaDB4PRt8
6JhzLAPsEjYi35wqsp1LTatWq4sT9xCoFoPt8z/F/EdHE4zJyH4EDddMQXO3i8Cz7cNjwRU1O/4s
aTMHlQMB5zy4fjb5ZHe4/aVVIPHR1EjJ7XobyxfgMvOZaQuuII0c9U0hwONfrxhSlBb3k0vfIH2D
GFAnTWdMmFAbCD7qDGyCwF5PvrlJcXEn1tjUibKO2d1yIWtzaYrbpPPASJc4+lvs/4bJCuJgEek7
11TjgwUo1SIqQqHtyULolX/ANweqnJyS0xL5b3R9vFhIwUUG/oQx2IgX+zO2qOOMhsCyGvxrCm1r
4itYrCspu2Vph5leb+nuLjuQmJH8SUvB8kKgma3N20tUkVw2Hq6vdxjwj4z+a80Q1UoHOnF6WmqR
HpysHwJ/7dw3EPrhxlQdy40+eZHXNPSJkE+WrVVoKOtsqut7Fnp0qrdrWrmFRhgLiMHtNAPeZ+Dc
MAIuXABMTtu/dMuQsYGfZflyn+PWBOnXQESQdI47oU0xz/xaviNO5Brv/AR+RHsB5heiqIZDJ6BI
3MWD8jUVazNSPFzQrnqIyfqqxqjqPmzxGp96Tj4Ya9gNSSC3OnVToagN5gRVNhFH3HpsuBOc1Cy5
AHL0SBekd2TTHVZxmheJDgkSs2eCREYjkOmJSjsmamLo4BrxKYinZ/J3bRBoetbgh34eWV3cbUsP
hd018ZqFr3xtcXuHkOfDkMglsj9WwmV7bBRIAElKitn1JBdzoXiqpUcDSM8ODPwu5jilE6KrE1qN
mNzCcXLLpqvTtaVk36d33piH3bnDMC/dZ2Nh6us2MGLDDzyT6OlnY0KPYt/PYZnI+w8Q8haDbV2F
rPj6xGvwVwAcoIh5NBri+J0tyVICqrKwMiwjAPH2F5lPtoknOQao/e6XShTfeFfk4NDWRpc8l94r
vHhwKP24w0SUwRQSjjKwKfghr3yNKpxSvoS1lWlB/BZ9IV7A/6VL/esNUHTIG1BKXJnGTABq8/JV
9kOB3KDvMCYQcMFuphHr9dY8bVA8IlK+/l9p5t3wx2WN/39B2fcLm3pwRsRPHs0wd8Qd0wx/Goy+
iYRuMJ8WHpGB321D17Da+IWScCj3K2JrxZOyoPAUYwTSKkwe+Jd3clQU43ARmXzGFa4Ht1Q6IFry
d1ElP3lVooKX9t7O63t8St/G6uVvsh46E7CVeyL1Aa4oifGJKpgW6TFQUGIUQepWWchsu+fNbI/4
HqtiKUMXUbf20VF2cnBsHcv88mrS8UDNtBW84oGF2EUsvZqoS4mS4htF/s/G8pZ30Qt31PleBFNi
Oqxi3cQtIMbdMiWx9sYEopugz2ivwGyNpKh+dypkHFulJSAbM6e5NyDVz1fT/ic7dai/2TLKqGAM
7c7WX0ZJxUxamsNjaDIuLI0MMZFwzAmGc7VNYe0bcszZwfv132NY3dUZMIvS6Uf049Km/GHhQLhL
EmjW1zHrBvxWUh/LBZNLN4/lzAwXOgRjXD36rDoDvfRhZVe48kQ3UoFGl7uE5CE+bNNQh2PlNpVp
+a9WL/DTyHIUqATa1GzgofOxNiMj+ONQyW1hCHA+Qvwf1ajqS9GoBjo8lwQTRaUnce2nYclQ2rZX
0eXZ24vm87x0z2aH+iHDQ8Od9hDLxPtrUQ0B/cpStn6F0IGvnZrIrCOQpvn/4xSJAYOmvhtix31j
MJ/MQL1i0IOWYEbUTosmy/OO6CMPC4Mlzo6nMUTBoQ/l4MGpOssTl2fb2J2iDYsaVhviZs83h1PF
isNN/6AWoTmH/I00xGrhQjXjgKg2lo8pOI565hBjGL5iJh2bOg4ZObTthe14PxTYAPwywQfw7K07
iR8QGHNoJdhdHgSlzAQ6vxZe4l3r2c8it5XLz5FBtR7su37S77Htrdf0FrTXr41iIf1kXRm2wyL7
qnKs4nOGaWKYzNrhHuR00vuS9IMHWifbOGHSVJH5zY+L9K8r6eK+SB+oT+zRq6XOfIy5K0RU1WwM
1D9dNle85KNaDW7VbX7YINnsIvhI5QfPEG1o7FC/O7s+aee9BiWMEqysQjTyYcZkJErrRB9REl5e
ANqyymf6c2h6PaEI52nbZj4GAOyyaD2lNUZXaV9i8dlznd8/J8+22rikCoD2GwjiIJEF9Gu5batY
slspl67mqzbgtTAsZKA6UHCVSBGjyGDTB/57ACyOOOqEc8AbXn/JBcfwcoNRp81pyh5up2sie8PO
IbItbRB5S2iZQpnnHq3cmRSXlZZcPoQscoTsVi3/8budbMAzoxgEFSO/DfqTVnHToO3r88Ahs9z6
PoCktKJoP/cDH1ym/8xhNywnnl+4yr7lbYnfEUQrfynu9SOrp/dtd4YcQNbR4We2v3qJNrgGVYpw
0r03QCe99OCGCGq8YsfU5vGWlh//iHNSca70I80jVbDp4ry3bc5dSU0co1eJJuVv0BBk+7JYEImn
trAQwhBrT1cDey6CGXMrE+HEJ8ZEzMAhT1qY9rAMJ2B7lJEwKxIRL8bosLi50aDITZxsYKOFYtLM
H+or2EHv35gvp1sRfmq0dG0lXNY08snL3UiDAu3Jd3s9JKKx7fJkY87jVAsPJX2X6VNLj9UIW3xo
GbkBncUvYQi1i0Y7DAAprEJtWS7LCpxoVeXsGwjJnifkrhCH5EfHRt7lbDdv8s6ywrfoxgPjkVEo
wO5l+bw9pPA9XbsX78Zt0Me/xRQV8iZjF4ABArnQ+uGmrri8YmUl3wgMsTHRs0nFKeBgDPE6UAyT
Kuv586ZCSuxDC12AoZ766/Jxv5W9JbDQIHROEuxhLFIRufrIiWvuSFZ9by6YyG3ijKaNDxgBmqvq
JOmbRWg4hS9lybYGdHuuUNhGbjRM94qFXliq3wvITnwmTJYYeqDHOnp61nbTsVIAb/dvlnJPP8tg
DutREJDNnSBzRNQ86rr1SrXXG2nABqTTrf+Mi6DUwXcsHxwh3HV/AHyJTaifdhY/4JFr1LOwLcZp
mfIDidtYHjcnuxpneg9cOJWZp/PJbBWrll+4ATH3H4nRl9bA477N1GzpHW6R6LB2kMek5v1zyxJi
SuB4fVJv0xxMSuBaimu6meSyI3RLzJ5MC15ojHg+TNRGgZ59bjoaP9NLexun5H3I/eFZsCe1ghp0
F23iOARKg+8vHdv0vXUTgP98w7Ds2Cdz8SDt6JoRMdiqkD00YmpcQ1+UuD0jMMJkhw9KHTxMQlAt
5QgCvv6WA0zEc2YS8jcv+tyXvgxpGSpaoV3jMwm4o2kD9LHtPRdoU0lpzzDOBzY7oNSYPqtWSVYX
Yjbr4hCWWOdnDIh5mzciEWkX5rF74wqD/h/+pzmOOsAEPjnprsR8joM0s1pfE0IF57MZx5jaPIIO
mudLcKFnRnTeWI0o2wTl4I8uq3GEvzCUoRuXcvoyu2AkMwTiC370DB5XV6/LM36dRD6phCnwuuU/
cTKVlzdi97La8u6JzMRbMA5XsDdXs6TSoyshMSnIduYFu4pScfCB5cshp3v+/0+ung1J2AAu2VUS
LVYv0ygLw+J8fs/4+jwTp7Cvi9M3AyjUe/pgbPG8hVwWEZkw8fVR7L9a4I8Qyz/GpElLO9CN5abU
9+Yfb/Hj6ffh8UUdLO3HXp6aiozt93ypxFDnlU9sXpHoScxzoRkbvD9mQhzS/Bio5+UgDisQqieZ
nqtJ5Su4ngGjuhvqkl3VLzaf8Of/rz/xO8/kZYIVhyBwY2j+iZfNuhNtQODylzcZnr1+Xy2oUdd3
roIgxyrODAZ0J/c3SUBy4SJWlo/jDzvtuGBoqvJuxZUhUSU6Kj6pJntqDbRV6RlbwBeQ726mABgX
dD0gdo4Wb8kOprqrbJBP1n8nvSZikdSMCpMx0tO0cIs6o6sGAaGY0wNozZ54dxcqU75SHuoZPCr8
dNVj8XQwrUaNxS8vIYTyogYegTtENyXbaa5yBGTbZ1Za0bCoKBO+ZNNLMW6uhA5YyW7+GfUJ4oJL
6BKRl512ZYXVD3aH6B/BcoYp6EfpUgTMHAhJnIuWxOnlZDAhCiUGkbxUumagtEi+cMn+iYRfR3Td
gbHrltaxECD5SnLAussPUxcrh8UlT+3EYS7eLTR1h30UTRffjKDLP5bnroqWNSO+eKE3Y3Okgagb
4pekkUArX9SYPJSzrwHjKMNqIuWTFlz0EEg1Unzi7Jg3hvBedb9CY8EZek4cbQNkAyx5vqk01YjZ
dxXyk2n3mNdIynLHAFHIU1eaiNjTfbOdeQ9Nafe80CvCJ/vC2g9WOarvXbZU/bRvDhM2QfkFAO/s
vr/o81xFItJya/qGUUd0VuRr+ZPhQhaqzlEq+rqIrLTtr+KPaTO48TnYHzW4UlZPTx9kbRYIWJb3
d7Uf7hrf1B4PourQd6WpSGl5NNS6RfYne/h6cQpCjjgrj96OVeqtnfhuKRJI0QUU8uGo38a1ZxER
gHfgMbKRa8gyjwJs9RcNoUJ8/ka9cWpQbk0tPCk4dhldUnz8nTtQJ3txsZdpRQWQZEe2CzN4Jav1
UG9FYC57oSxG5aG6308M3JYA1oZtBlSYaiehSSHmHp0Qp4bclQ44Zy11lMThmQVIWkMIjatzQh/z
2ojmq7q58ertOsJ1QgJPBtfijY12GDbJ1i57XMhCvZjzLzaYmLjTmCNjhfM032fSzQ2zkkI5+xu3
rpfIlImO3BBADB3PHEwTNx3BWcmBtiyXguCtGGpLg7IU0yTZYnymRRpWjQ+E21IvjJynfnekHnU/
Cdq6A6DzWuuvfwy9hvEoIHsSCVr5IpwYOVAB5hCUh0DANDslhF3LMfjd8wCoxV/FnFeQDHEnm2mG
t6/ZaADs0iT8priOYxcw9X1xTtdrmDapJk/e/JSxJ4Juo4mh9hsQgnjtgKCGPXFhVeW+9ykovGdX
u7fIVxsD+k0/RiKKrmjUtiiXP5ouFpEx0Lxkczx9FWbfLPdimhNiRF2PxW8/4mwM6U2yy5cYt5x6
1jcDTJUMBOx+4vSh+L3upr1NwVleyFWMG5x7mYkQPoOxJIx/pJaTonGVw8fLv9qFouVtQsJ52KB0
bqtrfuUrJ7OJ7Ri/yOLD1J36h10IG9m3G+QPQDlf6EU7GHzYZUmppdlRLNhtMnvY1j4bdyC5SDz0
rwGqjuU9aoJBfsM8L7in/O15xUnn9Vx5HZF4ef+RYqpcDCcz5kHaBTSCC7NNtJ3cM8EHsa3ntPen
lDZ1x5JxRoXEjBE5PDOfoaQybnWy+aFth5q8Hg48A5s1TDFjumTFJeCnfub6Fw3HD6F3xKOpZZjU
RjNBOO6kRoa7RG6V9CqPFpAUqBVy2EgcbPzRh56NWOeQtQ0pUlPKl56gdC+FzvfviHj1+vZSwa0/
tePBIh/Rm7rC808o+5jwuL4PDPgjja2J3W4VP3SsGmOLqFNlCO5kmp5zrIA4x8koY11Sp7kAEfmF
ZjTJgUVjskzezajYXwtNSSPeljSak5tL8Ow8PNbyT3fPV8Hu7hAcG9PQls+0RUv3AxWdKPgEVElu
au8CUOiWjg5JaQYTt85mA0/DrLyVkcTMte8USUlixq0rnpPIVDCr9K888GxqFamkLTxzUeqYSSdS
PmjyHVAOADDO8QrnsXywxentqj+FgFpNYzryn+p/tafjg/HMMWexyAvs9R6CshMFEGHSk8doeQtb
Od7tWdmlyAH2ywTWnxTlJBO17Ro5e++xNCdJJoPEkTJOp09FBEpXgDrUgTnKzyrmgwExbhi6iGjz
pvL8pAsuszJVhTYlw0u0L+GQFvQNM0kYrmUtLTMZcElrBlI4nxz21606Dz/6ajoisVVRzX2iHUmz
cKWDenDYdhPaNSR17nk4spoOmWw0x7GhI0KpPmhL8lBhdh4DcB27Xx7jhIG29p+CoK4lLbRQK5OG
Z824FxXX3e+ki81BzEhBrSmsGxHRAX320FWkBzyXj06frQfklT5P30BvoeO6oAw6ZphFP13QMRGc
ELvXvXGss8SfvHj++2mOJNgHiPnCpmkamVksEhRGu1o/nhLnRZ+DuWwHw++xMEjaBFd/q9KwqcRI
CMlda6wYW6Hy7kLVakG0KJbeSEh3hb8fv2jkvR62mDHeTSDPZKXot9X9y3ENpO/Q3idsekFdNepo
DSjzk7Hy1AKMrJ4Nje+11yxVVJXNqiBQlOoY6E+wZJWetiU/kCCQ36I3HoWQsVWZ/8vcCxqNR19r
gnR+GbmlYOHwl6X8Cjr58I6z6OaUNhl6AkNSICt6g6NPX4hK+cKhgd3ngLuEsv+zYHIT9RcRIlyw
0JX3YCNjPTC60QcwZOPSZBrChf02Ym3/S1RueAu47mJ+cXD1LewGxSX9N9rC+OqAFmPn0zgYra1r
7lMMAvu1Yi7B1PT7vvG2gakRNwYmwjVxrtYmjH9Mr19Ds6E2XtBaL0oH1O6HCax/6++VUgy3TNQL
hZUhi0lnHRcDxzR8TyKRraAbLaVJibcdIrFWYDqu1CaLGyOv3EYlnG44aGu6aA0FqI/5AB0wBX+2
Lr6RIty9W59GM+YV7H/42Rc2ovsEN3xmlQt5fUnYbYbTgCOb2ru6f7pjKC+kqIpu4IysPJBiU5iW
Lpqh/rMI0K5SiqDzv9wNptIE1NccJKdm4Ub4tjG9xKvkCl0T3bF1xRUeVjObL/XyQL5FcUnHr0x4
MV3Qolgge49gtnzyaQ16KmEk2pEV3RlEpLz0QiVcX/iZmmoHU7YUo6vbwS9Ag7GLp882Xx8tpy4C
wy9IzwWjwVqM7K5DV+2JljcyHPuP6XVdokAgbgFNo3fH53jO03MUlnMuSG43wz1c6OUpgVW23BoP
wN456zRuyGUsESj4oDl42u1/2UVZGHf+/dYiIF3NXOmNxu+l9jDtOzR8dOhQhOyIrLeaness4Hh9
iQz0OMTu/Cw6Sh7avKHKJP1aN6NMZ9l+23IvfkMzOueZGJlxcLwRqOAbVEvVttKLNJqoRgQOFPBt
k+BPqXI9IJGsy78+aseFMnAAhOJuDfgzXGOD89HduPl4FVZwjZIQzFn3B9Ziw4X0szSZD5MiJ/0Y
PTALeXplveKt+X0SjmFKB5mWCSZA4iXHClMLZRCp0A+HGr465v2ERoHnggsu+GNPt7WFofAGMf+b
xylBtl19C9uCR0pZ7hHDFriYJne+Gc+14MO1oJMQgrbOkjh4sXJzqY6rUv5/3MwSUIZMcDGTpAkS
HksbUC184tio0p228yq+Lv6YIrDIvZwnkBt9UPZ0U0LEEgGATrtgLqgo982j8A9Ax/HSjeWQzK20
ySXmMLjFIBxlU/gwVL6U4pT6nk8MxqfbRKgNtXOw13gbr2RKUzeew6voag4rKikzqdVBnKtklGbZ
58YRKs1BUkHhbRTkCRzw2M1L5pU6JUPWaHJfJhcj/6HqK7iZESBJlSRf7iNn+Z3M/3MBYa1ngopP
EOyKSpFZ/2PVqp7md1Vs+vRxDHwl2P8u+PuJ5VK1l8Bo0SIESdmlins02SFaPNfF22x15N643JL4
4GvrErsNisa5IwvGR6rH1trx/nDIvPr+QA8fCyg2m9Hh+bByZqS2B8mlqT+YZb/+Objt2FqEWzEt
81g0Y83/vcziv5CUqKe9wm0nCMTb5nT6f3htfQdQjj42ri1W2KUou/pmApeOxPxoDmAcx91xIKih
4Z0ml8oX7C3pl57PbqCwS9KUUADv+Qlxi86gc4rs3pZhtpvKCkJGnhB875yP7ceTIoOJARCRkMu2
OP1YGoQz3t+OTZbY4LB1NJ2RF6SdlH01TJTf7ZM5cdBPwf5j+YjGPV7c+rAs5b0bZQ79KNAQzcHc
pWxe7ZfkjKO38U2D+CFyTwZ/ywREUiNS7qgvMSoe//qmsKzNHPDIO2K5LCn7XpXCNfj9YvfeAYFY
TDXwhgxOPmVbKDsG0sgLne70wXHiE/t8raP6xfwdCzrC6/I3jlbPA4+k7rkEqWHz0sdPdDrzYxWh
Mhdg0Fc1+V3eDyFOcaP9urHt8MQvDGZO/C4xfFC/VJnIm/n6v5nlXK9O9zlDozgYNtDLXWfoLYXQ
wldqMnxFfnxkLARdZnGj3XIHDLZoeo6mb2Qfz2al5IBm8p9we+pZBTaGg64hjtcAXhCBvnZeVZ2f
62w5M5YReA5VnWnCFybtmO65sRatMzjN+Z0gsiXUhYrZedarrJcIeIwH1uTv3yRnNdOY9pMUN1EA
c9wDI4Lx6ZOTrL3OVZT6q4XeN/YmBSp5NKb1TyTVP+yjTlG9JzSP5lJ7B9B0SflfkOq4xLoDaQa8
Bq6eZRicQiYtVYcufXGe5xn5tQTEDBLqlfxaBr6rEfQcqGnUHwSfkIW2GnKSDx21SOBT6BBXhHNh
1blo81exeKjfLODsmePxjn2GLI3lN3hxendMorqejrC4vofggjb1TEEqErBQT/uqElSJOooxxHlk
fTp5f9s1nQC34cjwCHH/RzBsV0q2L+GWT9SSqYwYy/lk/tALGzL5eEXaVvXKzezKOtR2vbSxtAeg
sqkWo8+6IiZOXd3ASGQN5wSFdZQrKRNZhdTj4ViEomP8fWmpyWvD5BxABzzF5tYEWcWiRwl6urSB
izuNW744Ipw8iaBRwPQrrD1aalWItC9hB3xRphv4GtkftN/68r1SU2nDYCcUbuV1fJrmbB5JmFXY
UVByOFdC+qCp6x4mHMstyFH8P28p3fTDTX5ZEAkyoK6oVDDfNanwlXlDs2fqy4EFE3CyJDcnsVTr
8r44JE6CpXyzLaQO8aFD5+dufyzYVgloGD5hkPfSI6pZegSoIVNdobIRAiho3AuHB0Ha9GMlpwCS
bYNt0v4tdVCZP6R3nrZgnNuSOdfTBY4flsHfS9AM5MNpxTgVql1TK7+dZq7cV1m58nzX9Fs59lzr
wD3wu4TaHuMdwOLJfU6ycokYeyPBNuBKPxwZJQT3F0i+0KNMnSY9KNCzPOEFXcZ+PbNj25Mb4gdC
y5Xal+bw810Y2G3/HIL/7GPhcyc/HyW9Pomxb5fmXwyanenye95bxG5x2+1AJqXHD+s2iCkw0laH
pzOhVgU5kdZdn0KqemL2HvQauM6HxvhRFUfO+SZeFjlAR96+N5een8tjLEC+Tm+pOGEOSHy4akKQ
knSLxmazMI+f/gvvgkev87cKWp9CXcVs7VZEnV7UJ07CCX1xrORT1NxzH77udml5CpY5+vmmb84u
QfIGDnaexWK01fJgT3tmGtDIcrywtg1OuMgNJGxN1wG7MY5RiBnFGNJlasDu1Uhetxk1cESjGiW/
5PynRA8ccKGJnVe6vMKslRUVb0jsEBrT8DMrtY0OVd3wvVsTvk/sRQ0l0deVXruVGI+whmbAgO0g
C1RhHtFBFwxI5sXy/vpC5NW54QqLgza8rrtyCYFsPD7GIwlx9e0yVXnNoGHWT0gDgefnBptDvFZ6
96nuSmzY7n9+yvPnHpA2nKX28ypR5dFfs8riGOg9hI1ldinEL+oVLxBB1Jnom1IgrHxfl5Qc6cUr
0nAKIuilC+2zHBaR0NbH9GyxeYY2dLFcHDlqlE2tWlYSV958alG4QG/tqfcZG8ulBsyuwU12zWos
i8uD/w8HitXWWQjlkiULF24PRF5M80gvxwWLrfh55DMoe33cmyKGEDqnO6fhxL3aI2kL9RlkpHvR
/RpoBA7UxPQ+BaKFqwsFcEFiVIaE5iq5NSJJkih/lRwj4zbcshHh1D1yZJyTVgnnWgBTEEEBoE+B
NOiBTIRWYyarPuI+K71YVFbpnB4Kdx8II14pu9VF2R5PpQFroAdxn8GwsaQ7zXUJn6q8rQhPIRGS
eBnckjdVMd7RmYoRYaPEAwOZG7v+u5HRQyt1NG+yt/3ulo6oEBDJV4Ry96nZS+3JxzkQ22YQ2u80
4zapNImRq/0EVLBl7gcQrCvOw0bvFARdUCK1bQ6CxYlLxrYgKrmHF5SfFes8xxDe+/7LUss+GeFV
A6rVr9EkuMgYspfs0ySXoh80TOFiKWKoYmUnptMzsRTekSXIYF4uE+LJkP6U4uww+cEgdNBBRFF5
/THIZwInjfnuWcyLGyTx/LFNLEwxopgshZcbKVpRISCKVthOzNE+LdlBZd+TbV6fZJi6SlvUQcld
md4b1xKQWbpmacV2fZ6GhCWz48F7eA7Zj4MQDDI9uO8kuChA/Q6fDLkM/kOHPVM4evriMPxeWGHP
wLu3P+lE6OcqlyTIVgRtloGZzsxlZQI9w4hCKsGQEyDPJiWRXyvHJKXYbrj68enY6E5psbn/dOIB
sIfkIdi5hD6+lfMakOQNXdNoMcYsLC1H43y3G/ychW5HdggQDB9uagjdYgeWMtTWewGxGoNEpqkF
iA2ZMESlU4HGiru8PUI+kDmadODXrJoo+hFEY6qLWy/I5x+FfxrmwxcZ5AuuGd/WQrfRC1kzd5d6
/BB8YIyIbW+7Z8Trqy4zVn4FhOLG4caQ80Z5S0kLofy5WIF1+GvFJfB9z8jwpjEfJ3L1RDXeC5e6
bVWxwl9sKSLXdjJEBpIIQjBPTdU+hCpaLgzrc/r7lKGS9z1gI8CeHKhbM8flG4SSyyvXubgcsVmc
GZMiIW/l73InemWGOZCCmWff+JOAzhR5YuErzzYS70N4CvJytnRo3tFW7CUCrrTYLyJ04fGwwWkG
f7DbeVaiG3fhwopzwo1raFQvctwL1x0yP3Xx1pvGeCVBRyaSF3qz2xT0jjSeT/JXGXhOsbV70ykI
5qwkEjnO9bTv21WFVxZR3YH+en14bXP7pLrw34D8V4AvhAj2fYiMmzVT0LFSYR1C2LqjQW1ockFj
oSRMH+JulV0bVv0lYRppZjJ7jilSh6zTUYV3ykYtHfSNvIEIFNtyHrA6yGAtXzAZdeFeVCJeQKv8
qKPyLk4jhzJotDbTdZNM6+Y5RgvNIGObpV81InHu8kN4YhXah+Qx/hdPX8y7A0EWt1W1ZdF4L0Ob
nGDpcl5X8d5GGcbGkmwL4K0XfleoalOB4szLrMlMcE+YPrG9s2UjGZWI4u5zFLQoJFeNAANxDheh
BdlUqm5dadtm3p4uOWfGmmXQDfb/OtzxxU9ASU7Y8E1hyKGSWxKkf72RLokF5lzS74fRlKLV0yvy
5qm2nrq1LjGpS/y8Ea/pDGEZaMIzemQoe5KKYF+DRxHGIPeGDnprtgI27MXf+ITmjYTy0tGDRNTj
wJI/nFZ5wxI50XRZ5gH3BglHXrYl1Evzs0uRTgFK80SdLYceyOruKtuirPH9lijjd2pPO2gj2phf
Hpi1lWoGZzHhbbbt7e3hc7epCPotHd1VZh8xEe/ftYYfOKsLhJFSC5yRgzyPCnLbKfXUtGWIfpmI
X3717zC41iI8ASxGWoc3sOn8N0aBJh6KuL0GrbxZGkZZmUxeI+KMt/Jy0HfDN4OcoqNIbQpQQWFJ
j6CXei9Idfc5kI3pQTyeT7mknUjDj5Ce4ILUzQMpXcgLw34/wWp44Mc0yZHDkMIy40JF4TaQRTK8
vVzOeRkrBfM5KmT2196FyYYJyE/nQL4CCtWIF8K0F5TEAWt45ONny2ExUY0L4sHVzRErXAQvCdak
B6xfQ55pBDyKM1rjOmLmWOKuKIFq5NLJLGCL0rvkaPRLGdQum/6JOe3YysW82E7F8MVI1rQ6rhYg
Fs9gekiPdPueyoMkq9OVaCtBLytRhpghhvmscCP8/1UToMtreF4HLqzTkkPDqpK66a8iBO/zNiys
L7yVKfP2dQOYUZhEF/clrjhDB/7QzeLH5nM1wIdVe5qOlrWZs4SXgvIgJenIqVNrvH1vx6KHXbLs
k6ShXgfklrNtb3kqbS2a9K+Um24It8BrkaghWW5XZ/uVjKZnXoCDpAAQIiDtzfSKCdy0kzOQNSDP
2G4o6pNwweunojbLpIP29XhxQBYCDku2QjuxMZy7GD4+WdJqDjjPSssexnWwTYkeEhOygwaBEVz+
zIZtnCpoOC17cCnGllpe1SEl6T2rTAluD5uD0u5mfT4lbHzGhAjWydlVaO6YVhxS6Ys7GeibOYWp
SUEslgrsAOkWeXQ1Np+VlEPxSDzYWllscWtzf2DeFsfMHhvUtU952Wd9XNv3Gh8rMB8o/j1vhrbm
ZToLRQIMvnTb/aR6hV4DcjNubFy+Fa+I4X55zZ/FZ9TUncEEnZLWx9pCc4S58sEXDZZenLCHk60Q
iKOWh2vyEYjhx3miFXJ9s8ORbaHsfjKuT76Gv+Yz33wiLMs5UsuqYx6xc3H0O2Dkg1xMSp3/Bldf
joqYt6d/7yO+fvQvFCCYSSRQ5Vo6r5IknkGHfQTU0cOY71rUgTsR/+I2UerWXHBb4wqlmDDEOu1U
cdJ0p5g5BsIbUpB9aV8bvyfXU2pNw4RccTC7ppTo+isnSTdBhxn6pKj8vfc7kiWKKO2R87xHl6YN
GVqSCqCuiAW3IIL5xC4ex2KsSGNj+r2+6LtNaF98jGW+moX2CMexQdSIKxrKgj7g/IR/nt8fcO34
CtxuCnqxCcwkjBVRIBVECS72JyLhSYm12encVIBg5wFLgLHZYmyEkli4zzYVlrl9+ak8KHNWgcjd
J77Snitms3lT3l/N/oDkt02RzxkEHUxt8NHm9CL4KlSNf1fwWEDM6UTFqSZaghggZvF9Zi9OBQCb
ftE1LZmFkFhcRqpcl5HJQBc7+aSOVsuFLWda5M46Hi9+nk9DDnZkMlgP2WTRdVNspgrNx4NNiu1a
i8DwOy3cnxvXfPvWUzUkhFrwZzsgZ8gduUPXr/OwTBwz49P7Tv63YMXZM3iRRcYGt094EqU6PkSo
ev1Rzt2BXGJ5qc3woEgRTPav1eJWn53AVB17bKuMU815RYVvm/lVEI1Z0yEpXa+phGTAdj7VfWt6
90pWiHTjG0/H7clhoF+MqCVf8C7TTqpLJ6vdAf8k04/dBUghzaiOmAQZ7wdHUo6J8CqdyYSVE594
Yu4J7QeDJb6h6swulB0Kg5pXwhXUXnK7sl4sWgTPPfo8j/PH7ec8kKHy9vDV1bEwgwIx3f9SKgdK
KcO583ZK1OV8A9fonefEPksqhU2615n7Nck7ABwDzVXskm+4swnY7FsLRswp+CZcN/aUNBVkjguN
qgUgNkqq0J5IvMgbLzI3ESO0s3be1ZTPTYB5LvR2iZsGNnnyLS2KhsnPNjx1WeNJjNioRVKop92S
pg7exNxmDq6TDJwrrqWJbmI51AUZ1xXmLJFP8MfjSeHvFA9dpWveRhm1mQBDuSHWv+9yHwFP+Ga3
B/QoVlrtKbr0cnv0p6wa7hR41YgRoHErLgP3db6e/gqxG4ZQqDzMuciaex02HGQSv+kzltzWki51
KXohzVT+F1g5QvVreBDx2ylDIvpDuda8HnzQq5uMUiaU1SRKs1FH+FKIGlwEhjaBQZSL6zdQdfBY
eH/0DMKrRg1deUX50WuvDgia3GyTuEXsbDzTlahlvByD/yCYgGAzhsS91HgdiJ8nhzEQHE7jKXM2
vNBfQ15hole5Vo8kIsSbTI0Kl44sF1uHSPqXBIpflUukO5157vZSa3Abvaji7dw5l4peLvJC71OV
cxuO7s4WZ1tm47Pyvs30Y6pi+l8kMpk00Cco42K8oUa4mea9rd5GFspx8zJ332MgMsGdEtC13ERp
m7pNsIbDws+H6kN4mtqLWq1tClW/q3Y5nK7T0I8RrUZqsF15OoaZQVnsSNiUVzYptHKFRqW0VkFD
gvHhdcgcZ6cQQhW50XBOB62QDKHjxCsLvEroQB2s24/Z38DPiAy3TDwazd0kvGuUPASF+vuiXd+7
AuYRI/sd9Q4WVz1ZDkQouMXIkCXBpqVoa+fjI/lgxmuOxmP1CQiLLpWsVUUi8SKbq0OgwPY0iHnA
9jF6nLh4mzeSY+Yj3SNxUHLUITjZS6YtSW5YCWChiHmQAGu3tIwuXfRcMUKMXK9SkkDaSB9CvQ17
AV8HP+laGmqEnvHOL15VLraOyf8fp5nl1Zz6pUvx1gM4/ozEEEjuN8IRB2aWF1s3H9uXAAr33+xQ
XDlkGPKDSekBPE+KLHqHEDcwqvDnoFXXRBu1lH1FauSDy4yXSS9HWzlOsH1E1aYxKJBUokDgIZyR
8YlLTYkCKbRArtPftvjnGdtbSGTvwwcPhaJLTyHPQhKap96mmcHWhzaZ3zTiMKfZbGkbBzIVzTQV
J+MOOYvr2DfntWv0waSdOzxsqFJhS8P/m6kM2Hb5Ldmjw1DLYt8Y/6jcLZ6ULdoyaYczbb64YjCH
wO7fg3NaJtBfCayDltLqFeDu2ooDhEWqngg5XHVZjhw6c5NdgYFrZMEEEsfQy6Eg1c1UPO4Ta6fR
b7G8zMD5qKMzyFm0cFiyo96szL0Ou1cyZ5VCtK4YEzQmI1ZmthOZCS7KtEhP8oOH9xgxwgb5ITbF
qjEBUtErT878iQ4wvqPWJKEqjrrF2YZ+WoqakvbI6kKnNT1Fb414L1afEG/YBzmSe6yZSN0cTBiM
nXBQzQUcKNlaK7Pq+NZIfiZIX+sdonbOAVLoMTy74il2RXs0Fvoz0fSCqrA5HLcGRQZC6CaHBkzi
tJ1KWpEWC675zRIgaFdgIXm8luZVcFiDFqaWh6PUMHKdWVFwiPskxcOKee7BTKNBCZa+JxifUNK+
YwtUXrzcwv7HeA3Q7hTvkYvx2KEKJhZkcaxrmRTm7J44lTGYbvurcVYjqlZCw729H/uaaEGuWofj
q/o1IM2oujdYc43qIxDoOjLw8yg0lfCKoFlP4qs9Zh3/Oj4YGJZ8F+ORqARl5h8y2o48C+Q1q9Rq
KNdsUyQnAjmV4enkCgtFS2OdIfMdYpJ2pUGK3qcPn94E5XIOvDJuulKiGSUlnW4s6OJoU7bCyKfd
FnbsQlCDekyFvBO8BkEPyGoSWpQTO3vUVKt49qbzWD7OmJH0Xnt8mxTWvY1q5yDPMthmc+GnJiFc
go6v+wtgg5KdCNW13RCJoW1Qpnw1DzuQkM5UBz/PWVSMoARP7OD8hOztH1yB2zswhBrl+GO03GJQ
wedIEneWiuKrvgT+4H9MjQsTf20IhtFALCSPZyb+sOvIRkKB6fPwwCvD6weIXSuTa2hp0s60FdUl
AxCefN+3b7+9XgKxdjYKD2FmQU/haE49uOtijou4NZ71FiqqqqTxmN+/BzwqqIYXT7XRWwHfMv8Z
bB5hJ8xVgWZ4l/tVd23ffze8DYlqfKXLzEWxNn6wrHTuOw72f9zkVgomUHDT1tcvtJtxAeWPrX0S
NZ/ixwTSEL7mp43V0xtKycQle5J4Y7LnkXUbJMouaXItHHZBVC6rTS2qQx52lIJia4AQX1/x3IkR
t87hlq86Sw8y0lriY+bevF+BDO2t4rjQfEi6ockzY2o+YOUDj3UVzYIo0rEzjR9JahJzki+y6FRv
sAG3UI5RNX5d0YXuMncpQmj6Gjixfj2/AKdCsois0en5CJEqJ40Ki+DG6JNegw8BzwRsqS1s4i0X
aWt/H872BYYBBgk0DS5JpYC7o0yRPYS50KSxLbIn6hI+AEs52YLEae77m6rzdFv29CTPZzj0jSKz
fooXeSMPDwJK/ZHPIPFdJbChskFxzyzUF8L4eEHXhVDPnAabcnHavYXD0I4mjnpvefQSpyZJcNoI
FnHVeFGnUUuhvAc5nLdSGlYw0lxqpHSx+0LPurgw4d+9NKmdGocu0p6ZMCNmJREuRpc2vCHWFHjZ
YV2oNdlE4ZP+egJqMvjUPorrUN/WQSKDGIUBYqBqHraFE53y5i+SXoKfchWu201tIyot6xHRgFmU
Bp0lQmEzHNyxR7UtyxCJ3fhe2r+fABsO3iaYTfrWAHdDBLGAoxGtAAsJOjz4/76A5Bhj/1+FPmRi
L73oJGlvZnfUW9MEBy7Wi1+vKZUtfGJXeacWSPutDDwbh5827JjWWb2ZHwqYAxTfRxu+dZpTu4yR
2r7HzFClKAanEj5z34PvKOE4tRyW4AsxvCxcZ6GvxeVJR6tbgcAlS6oh2Ho09+F5UXHThgzIgedU
73T6atZ/5yC8mlZ5rFWxSf7eIH7z8oZhnpyBNMENDIUwLvbxx3X6N2LFEP/5VG4vcgTxJ1dHq5bA
UaqpljoNhFxCIUkm4M9+yFhFgINjKOfSXiFxzEcK9whwQ7wHsmUq1M3VKdfeRk3hXZ8z4ui2ZJBa
cJpDHB2vApW39JkR/x3Ss1DIenP6Pp0VLKbomNtHBmOQ/4uK1LqT2W016ho77PwqCJ4GuaCL5Voh
mu5YE87BEU9Ml2cjGraM0dGdqDh57FZfqdkc4CvdRGpaoFlUrGB4djLD0tU16ViOrFKMd47fpArG
WI7iO9ylOmLwUeK0pH1O0AJj9ciBsWYzTLWA7HpVgArJLF8MadM6RLe82/SU/q0kW8SqT2f/elru
iu5USUtgY196ZfSeN6GGUWKStO7Kh0tJJdTqfZGGitZjZiY0/XHdkBA0FQ1Iun0b6+G4DSnbjpbh
+8oe2K1hYK6HY62vNXkV5IxV4C1kgzv/dN5tXz1Jcz++q647467UZGWpKh5D7yD/RpYviykr8BIY
FDrjD9YQVQfVgGPbMW09hVDQ38q9W/gs3erH1WOMDE7VDgeXSlCRXoIosyGbDPp3YDDCulirCAeB
ZF1KdN7HZDHeo4/2Lj+bbB/IY4sDQJiWTI1NE8xpJg2FAcxSEpt6iQrrAb2g8NuuqLv9vcfxLR1y
hPUN05a0F4rTa7NtCSsU2NscZzj1lOiFiG8K6EkKkSc13nOlPZN1DfZo8RJ0A3hVhoz9vYn/ndY5
AxzFlg2t01UnMoZ53NnGykLiDYi0i45lPEEh8FviwVLVXSU7Vzo0S8zW2WaOx0nCwlZzUuRZtYvC
xvXnCiztbosvxWE/PFL7eCigYSNHO/UamgsALMTKfL7rZ2XPJq2FYt/7BvPZF3XS6rilMCGzRlWQ
YsJrjlbigMrY5X8aF0PzvFW+O0xfEYmoKwxtyBzGWjKloNi+ed8teUYS41clQhf/EtPssFT5tp1d
Ieclepq+jErMnYekaXNjhk8EJVRkMWwpAtC68i6rkHZEB5lBLlG67RSJhqnZab0mrBWtfLNktogq
inpRVgyCuk/5wUG0AtBvddPqwr2jUtX6Mto2+FSdVlM0E7KEKt29Ymh5krgAFVEE5Kh8PSzgGpnv
9GpsQb2XIbw8IFWVgFPVskYSAyW/1HO6l87gzofYaVgxLv4Mn9DpwG7AiffMaOyny+o1R5VAO6Fm
fY10Po3/lL5/7IlKiraz05DtKUii160iuVQE/ujNHRX9YfdS/wMYl/5D8cEwguidoBt0rV5OHUN5
4c9iFpcDwh12t4TxZw0OsYyaPLA7uTWwSeltu4W9BcHiM6RbIIvqNaJoP9VNaYqdqpxnTVVO8UFk
WVxrqV8GWc/I0QU/VTYM0hBD2zv2+TWLwgFcTxgY78xpjQLP0gEUO4txg89jq/dp6k2kVHyWqzRl
OCYYmkIHqCQcezhzsrntO6J6sFY7aSGp/YUGq/C9NiYiyGzRI7sIaI1FuDTe+UHo+x3GU+jspde3
IscSL8C4g7qFbbIi43usJ1aDk3/TypkrA2teyFPTxnOvL7tk8/nTVcAxwWrBf4IC0dL5eVg6dGLH
wzDCgwlMNaKQwi1yPwk4fc8RoGuADnQY8RXr+SS7ZohHSQpcYwHZCO1T37QZ1PV3pOJiyc9URAYa
x4rXOE1nazfL0mDXIgwDwaztyKYJe9SV3n2UFo8oqv1YaVGJe4PljdPrzbHFBmpsQaXXUfsOWyhQ
mQcN4cBRcn4GmxfgqZ/eRIl98UUOc0c6vyxjiTKfE5Q9HFi+UTXSx84fgERTFTMb/7kJE8ugOrfK
fMyLrwXrAITwUmhBW6by/cizpETh/G7LE6YoEIced9DbumNLllpWrF23o66P1roAVLP3YwnQR2D8
oOrPtf0jYBsiGctR5lBkPfWLzx2IjmLa9KnlvAs46hhQpEeyzApoPt0caVnGFBYKdxQhilNbG5Po
yfb/9jzfNvCvXnAvTVOb41PyyyjVSX5/RPg5An/KHihboEgiLTjVU7OShvAUGHwXsXGYr8PU4Dpf
BITwheWDPAhAGCyRUWPFrrSJ9vZA/kJSQzcbD4Lm/8x1jd2k6E/vMLOI5/z54l1GWG9uwXUAFvAf
JKqpasKzIViDhz5pgCyedG+2LO57bjyxS+pd3fNaYtxskGKi+AL4ntLH+giIhLXLaXweXA/kgTCP
gEi3QsuE+bGclvDVCw80mZrygrEphISzoYxIWarmjL4OU4s/2uaUSaOHeW/HI2+yJFFSgp55PN/M
GIkgCvudeKRlDXLOuwQKAUAgefxXzSVm0u/0m8nfRrEu7BJqXORgIStDWi951ApEgYUku1fD1IAJ
ZQhMpM1X92RA27CFjlIw27aDHWj3mkADztm5/YzN/cPcnvmHO+R/c2SpWjjNMHAndaO5+2kr+LCb
TfUpRFbh20ccTVjhDTvPfHqKWH/Oy/dNeCg3KNmFLx770cdCU9Ek3Il8Nywt1z0zYZyIZHxihNlM
ElbFjVuCBTgH3fGmf6SHUL0VsE71vKFPaXyg1qwve4ei3jPwIpv778+oz/GcwnR+GOJubWzAvtFH
W7G7YuFxDX1LgdlbXkI58JbajrdVF1MQqVRBzG0ED16ThYrZB6y7+d4RtC9S0pN0r4ECdhyya+4e
BKpCxtToATbP6NaoWnzLpXAmS2rhQymrWAaYnKzc9k8ib6VW2IAgoBZmFAkwDc+AouTT/Pa3gWU/
1wS60CfMFwCAcH/XcTx0Y81YcCm9/XDGgs+aIfdj8/5mpqQou/O3kyXoHfLrZi82FFaAcW/7Yu0s
Sx7u35lniFZVgQZ1DyA0Wq9hv/sbKDq3puVFosB2njAqv6qDJ8CFD+Gt/lENUEdUfM3uuq/4ZuTm
86EZ90Di1trEUK9WCHHRyQAWCajn0q4KgHzCs6bFtrMZZUDdLO2gKv9RcNoaNezQwzIG0thLaqeT
wgajf4bdHsSXFTSTaNaJ3MpHp787L7WqEOkFnySoyvufCACYJ5304we2OjVrq8zFTrPcohdxuPnd
EYWCXhp0Rzc5WNDKFs1bEOLWn+iku66NEbIw86Pam97dLodxdXx4uwuGUJH5PxjvSC08XdiaIvHb
OcXR6hfD0L88ufxu8DU70mrmk/r6Eh79ZutSO9N9X+6YUJHwqXRJmTItu80pPzvXtbxpZZQIOUo1
PvvfmQXMg/QS08fryDbc6wdgcXQ/Sj/4q01dmL8I41IxJ/LywHLL97iJIDDyV3fuKF9Ca9ONbDBx
QD9TPXsH0lhJuQnR5DeoFbGTixbdrf1ehHx1pgQBQf5SRZpDGdL9tCmITGtwkZe1V/w/fR8vwvR8
IIgrJL96C/FJKZPctBRc2u9WDIGco2y2WxZvDu6ULnHpM9sfiBWzvB3Ou/zz7qVbYG6HSLrhz4hc
IdlCSqkqp3sSoUXrXJhV6WzJ1s07b0Ejg5MLao1SoUYbJ/LupzlXZ422T587ULhXpqu8xNrwPS3u
SpcSmUbqOzvBqidVSiO0vqfY2nhAM9njYzLFEyjQNZaOSyO6GRa5u85gkTVZ/k9cuQ7sXiSt3ZhD
iha0UANBarubM3CrcXd+dVW/A/IVKJYdUCaf8sJVH6l8Thfycng+/+z3OdWxX5hsVWS84y4zwKIm
a8PN8OI7mYms/3pn74qdgaBEa20m/zoYOqv/Icc7AHOjABcmUiaxZT+y74EFT1bsAgIfDU4ajPff
kUWeYVOFRHguOFsPMoQ/WtzE0fnwcfUt3qWKmQXBE2o0UyuL7KEcmS6pLb1kzbskhgq8uHDORFk9
r5kZDr7vu5C3COfvLIpQ7UotkeFG/Nq+iwfJdiC+gB43HjFLqN8hCppb77+HlO0fZEYbrtCyBg5u
MZ0UvFVppvf4dAb1WVC3fBgs2ReQPFz5QYjzmSURFPO9QdRqstaLRc6pX7HeCsUOWxpm9YyeLahb
4xc5BTjDfYl5meff3Mg03FXkKoCVEEX29eLMz86s2LH0910va7zcneWz3MrwV0gKiai60M4nkK9E
X9ulY15qD72daJabMModnIrP1PqA75zQuDXlVlZR2YxWa8WbeB8JIGxsKbh0WRXvaTXtiPC7obPL
GUGck2zAwPU9pvBtjmDHf/kD5LA3cBlcMHub289XTVxBL6stxDmE7X2IaGJAWyfXemgSwnYdJYhW
iCG75WUiz78wQgwaRUPKKXqXibb/TSAc2tuIzeWYd9GrB0mU2j7oCrJTTQazlHl+siNFfr6pngBy
SvOS4pKbdMoU3mmffQxXsIA2wRhlV2k8mXfFX68KdvEp57iQux3sCEN30nLdjBRRg6HB4GVMMqmN
0ZFpc1FOY5LwzQG2F8BMihQm6g3PF+LsZK7Hw7hcPIijZZ5tirYGDkzli4prkiMDhGuBvEzaYsvd
g7cXacLTw/QPVuNCnnKYY3Ps9jc3O9QZDAzgn7PCs5CF7bac7Lkz1lZsdECCqUHs0ZmELCP+iOLN
pVSw9cvh0Na3LghXPglFoIOlcJK6zu8iNPioR3kb52ZEZzh6yXHya+Tb6e6g6AI9kl6Z1W38J0k7
4D2Sg+m1k2uce7/thsBtM5cctk+JaE9z96Ro2+6o5m0hpvK5RJKD8lOL3zJv/PpwdIqzM3J3XMim
Zpb2ZCvxZDnHUfYs7S5fkkj1PmXWPC48n3QPDa4KUJQZSKnkfRkfkSeeMOUvgM/M3ajWVwpl8oIL
7ZqttJe90ccrRDm8TjZJyqPyLF48Ixr46S+SzICf9yYR3SvDbDiTozKvziI2jylmWhBAwwEgNpZV
lfnPywP6+f3EMZGND001uoc6Dg3FYbeWtAvNWGrxoEiAqdCLSfb/jsp9bYhQPE1Yfn5HdM4Zx/AO
FGmg//fKW6xc9LR1ZR16tXs6gVPICMLMQBOVcXbFTdsUZpBLnkjzN8KhYp6TPbyXmRWA41RcjhUt
GNeiIss+WaDwI9EOtMhn7uGw7dR79s6JrBQvzYmoRS4dNUhSH9lykGwsQilIS0cv1a+D6HUZ1NKb
BbrZVjJSbdtBC+lI1PC4z8eP1vPC0pIkP0l9te5tv880EuRoGSHhimW9Yh7cG/5IQ9NFTpOT8QLR
y2PngwSsqFBVB0jeBk8e1y0daDY0E874nN+JTJsokzKrzBALgX2/B2i481fiSGSc+sZNLWFj+Jn+
JgWp+5Rg+zaT34cCN2cBr33e/jJ2NjsJQCwjEo5idkda8lAaMLpnyQEfxaEfvgyIwaVxp59Ya1SH
jy2WjTFY+KaA4LJU8XklRY1ixzGPaDxZQmw4VTXoMt2s7sFl7E64K5mct09BB0NRrd30wQrvIeIH
7lWt/XHxhiXurLtd4slSo8DobyAzVvZi6fhJFsRXn4CFOScHt3cG/PShkrZBDbw2RzpsGD11UZh/
B+CyP90yChbsIJX+dxgWL2R4FlTOSSg/Jo1pYGVdHyJyilSUxdHUecw3HnMt0S9/RdvPqc5vZAbN
5GtI+g8oa4zJ6Erl6n/7sEpHtpCjlRGpEIgvTXffnXWGvRvx7FHUi0rSFLm4Ku8f+kt0vWuntWNC
WHyviViI1RMnFLmqNBKl7uaFfFJ8votyDCkW29qNqrQTOzWUP3DNGxIyn0J2ZeoLNVrXb/F6NlNK
rmUQc31TXo5LB+UBnYRTL3uMV96mgiLAHarscC0nW/OYQq/RbEsYUG3QAfW8wnq0exEp/6hZv/7d
f+f0/bem7mQn6026yuyeb07eEwKVyJ3WHyLpRDTxy4zA/xYkLBkhBs0eKD2JgGeeTV/pvC0dFDFZ
/ba2WNZEBc2KMAHqOyeeECyEtklzs1N5J0c+3d8OY2zXtX/km85dpfW3nEYrPehaEAZe/IMFuIaa
Z04+xYOA+xqJphWqQM4BajsAQU4FsaLP04678B5aIjBuDzFBj2ASExAjcQ2ldEJDP9i+XmGsnNRJ
l0HeUVZ6XA5j6m8ODi6LRd5liivsNBLNq542VsNM6fzCncz04G64Kk90tGKu39lJYFngkWz+lkzp
JRi5NN0sctMw6POMNFxjcmjui7ZCajZyFsrilpbGly44des2t3pQk1g5n8ZEoHMyOsm0HJz5/W/i
8p7tUDXIVcSc0PkIk2ljfrtnA5PN/927Acn7BOnAw0EsbBU3FeKXGGZQEI4R3lL3FBw5D7QOhRDI
Kc9SxcbMaLI1tX6aeK7nBiTl2jUuzJN7lU72n+SZVluaPrMZFe3eIfn3fb+rhZ6FU9UH0SdLE2Hp
4abt1aemRA8KmNoIjeKRkOXUt655Ip1amVzEw3Usy5hQ26a0dP24V+iCNVDZIDmuh1Vi3TGlSysW
el7Bw768dXXUcSiBn3WiupfGRbnkEEU9teb/IF9KSo1kIPnff8fEauhOI7JmoqBCVggNtD0qlNRU
t1FY8ByNUoeynSYSYxDPSy8DsXdiC7nM9nVwVa2ym+XR/ZZkhIqnVvCqLySRqjXs6EHYd6MPXCUd
boWNg9cXOCrk+EgauY1jYj8Kkt/iUADME22/8ayY0WuCMVIP2mDltYE9WmWCuFgNMJnmEJzYrNIs
ygC4RokmlccpdUf09C66PZ2C+yQVXUHt+ADZix7tZiwK5c1hUydkgA775uAC/WFeialSkWd4Vg5T
SZlN7uTYuswcg4AV0J0GlMR8pzMuEzoDG+Ege4B9ZnmXneIjgQQZlyCoqLt71tNZW6if3MSoMdX/
MqjQD2JOBtMZZgLzPjmg6WLRdJkd/ziksI15+bsGejztBgMrpT0CE609unDE7o1XuDe2W4LjOJ7x
jsm5uEdwM0IZOqjL754DF+/rkWCOENBD0/nwYHF3v+7VVHsHr2N99QXoRBQn6pjfJoiklW+bMWAJ
Dz1vhVHx4m1QHUsrRMaik9yP9KFm4wJOlhbFafphU0g2EIc9gLhDsKkQ8mo4FSt3RGAKC8nZ6Lcs
fBi1bxo2JGc4p+UyPjk5C0AUL0K7XhXJOwlgBdD3TVg4kHSxS8i47CsRUXF/5OeHl8OXb/FlRZQO
gEPistOYdYao+zPu1fh7PfEQYJA9JSzzu1YFTBZy8wQ8kVeuLj8P26EckbKSaGUNFsWwGu1AXsNb
mSvsc1Zs5ucxilGcavYCb1ZE3gOE77qc9S7Mjths6PuTlZaaR78FpIJIpndYz0izdzc93xP0220M
Q1b8Tx5rmmekV+8CPSvHgAdAmEVsb9vxKBIG/icP2ZttcVzbdGqkKvuPpaPZpv9ya60EutSniTuT
BBiVNdUTsQiB35zaxm4TZpesD5nvrcLKW2la7igEWEtQkP++atmkXHdqe61tTjRfa4EbFI+a5I38
HR9QV1a/WUGtNgdrQ3mt1SZcZFDP5mjTGVlUd8HZGQhqGe8zoNIRiuxwN35KBxdj9fUQn4YpTgNc
02lF6kWXnKQlNQ1i5yBvYNmvyQoFIQ0+olMR0HQOM7j7ihY6koxY2IDdjJ4vsCLBG5QjLiIJ6iWo
SNPqLQ5yVyNCK4VQqxegeVsoZmL8FmypCRuRgHVmjRRuVuMSjEv5pNlaKS6JfXsUwMtf/gQRsah0
ProqqZGrWixCjemWVJsdvqqOhUv45u5LhVryKc4pZzJalzimyKrsYG89qKoiSGLQrCUQFcCyKkwB
MWYI2MibyiMSk/WN4cC5qJu4djmskb3ancllhyI/DrEVY4+v4XZFxFennTHAC4Atkw62GT/nqnZB
i77mqPpZcWlqLFZzvcUmXTb0YtY5VHgT9RpEVVZ96OFlLwhA7Qy0aOZ+BQ65qbWm14UVHs8v30qH
vuIidISFGKnic5r+CQ/sbUApLJST3OsS7X/cv9RNgvQVyHTpnQO1/aUIW8CT16G4yZYb91oAE7r+
84hHdbOkAJn1Sj8EM22trDw79XOG20eiRQ13W6JHjG2kN8l0XoGGu5G9eV64cyd6SWAfSd1XitSm
w67OEhsnhYiUiY0YC0udgTuqVrlp6Zvp+q5CAsVniKLNl9fhb2zH/m8zFpIeIEDodmrgLyXWA3vi
4roI7JKX4DGg1aTNRA9a/iw65oDqYf2ko2bnDcamIKtHnsGkOesb7ltTAj1ZSfaKRk3J3ptLfCqk
aTdJCIJE253Z/0Oot0jvi3mM6yaiffsOQF383kwjCHJJEtnLASsL/NdamDr2DUwhjfmHOkCemV7f
+xv+qCoeXgFzd2ejmW1EqmzKuvD6koSXAuX0auaBlEQZW+a7uufeBYXnhiMng56pz7dJLQFXfOCj
qEvSJJzPKBn11+hZO6xj+rwIYSVbM6cii1T0pM3WsdVYCb7SlUvfSCKUoM9ylXlTLYbAcRLzky9m
TlvDG9yTrtJRTN5HzND/gyGl0QPxWoWWA7b+gj5fjPs0+8e4Q45z3D+rFRKzxneu+rHgp9WTwCB0
D9xrq7ny9G9YW6xgxLHUSFH/ljvvtlCXzZZan6r3mRA9Rf1Zeo8DBeXHcO94cTV8YAvluyLSO2XZ
EqRZmtzOLGtxdYoKc2WmngHAdvewCO9W7/Lt3LK0xSMPEGfaL7cVN8otpAXCQ0w0eZP1cQPZTrXo
vtpHVgDh4vpdtnq6R24Nw0d54T3JpVWkzsvcoJJvJ/FjIdiHzEuJn+mIFNd9fVIm/RxwUEGG8fyz
XIjJtCV+62a9GIv85Zrx+s7uS47pFLn6vrO4CjILwyqp0GtRMUH1mP3t7Iyc0G+SJYjlzqKzPPbx
IX/lVBzW9dwU2zWcBAVBT9DTwU0TbvhgUFhWkGM4M8BhtpUCOGmPrDZub8dKCnYp1LdNMXQflSNP
iDzlgwx2BJ2Xskb/Cw5SnU0lTWRTZTsgUG9afBV/fFnTwwc8vZ85vTsUYNhoXRxPWzNHRjMJ+dO/
xKxQqpAaK3o9s8wV7cgRfuoujnDqUUC3Vw0Hah6OF01cAkHU9Z01dAAonRITcKe72sUso/Tu6JV1
qcYOgVLRkQJnr5k3r7e2numgCwMt7muK5WhWwpdWgkU9NHHT5l7iLhKRINx4IP5zbxcaBbCSdEyW
VLHqRHr/xTmORf3NW+uqD6IHQ2+PGdOrjH0J9x0+vI6ijKFM6+uLXe7EDfGczz9dLgwfJJ8FNDIR
rfTi/wMRqC4DDMjHt3ZIELFg2J2IVkghFxH8yGSMk9BZerYaRtwf7I4r7u5nqWSkqEmmFLEWtwlX
ckTbkG5X8pPV/SeopL22h30WCeQ14YL+YfOIzmGVHH22HztsBTP+rPFL+yyPPR8EevEwahPYBkor
LO2Zj89kiaAspf3RsvOK+kzbMuLosvBLnjZFCkOOefOCPQfc93SzV3+bWhsmTk1AeGLsXJmkfRwq
4ddENaXsutVC9FntuP1llsevgpGlfjapxCeYtuIriZQxkLyM9QFtktCDy6PV+eOV99/ajxXPniYg
AifrKG/yJxeOmDKx02WJWIvkLIJP8bBBgJo3ZwubGW8NrOpJngx3jbAfi+wJEjT5gQlFSHkWfY9n
5tA9rDRx2zqLU2sF5M8cD4So4RfkDyX80kkvq+wMQUFeazE+pZ3EvAV7dYTLgVA+zMkuV5VKdwyg
mCG4U4SPCpGLmIwjBa1XocX4DKTUdl+WWLraPJtI8BfaiFzkagKmBQzPHAL6NXORzmLrQpI1ChKk
EpBMPkZDvizdr8nOdrLLeql/9D3hO6wVRcOgUAtsHy5M+h0zBaW9d9aaRt5pWjNbrLyrVtAZBnTl
EW9oRokH5AIzPpM7L7JvE9IPheADy3xe/l3YvAxNODfsIgz13nx4Es5bbeDKtCLMaf7oJev14CoG
G9B/CQMJVOK7G1tFlxkLRXYLhTblKZoB71ZDzG37TrNLI6aQFEsrOQRoHp+dkIVdo9ir8Y6Rhd/4
4ewP1j+eG5tm2LiJuHp/+2Aa9gqUeZir7Sea5ML3xuay0JUe2DwMfcLIfRiHt/bOYtfiUSjQr2lD
Kc9acCgs4v9ziu7CEyILAI8km72goF6XhdfBt8NIG0AsBsnCY0lRjvjb0EuXkVspcNaw2QUrl+85
BURtLO0OKJjlORTAgsrcy6AunemGPjx/qgijhu3pQZG3rACSDLriCPQVUQ3cyFdoa+wZBsP4YPMB
pEmiKZQBin3UhH7EDH2tJ+e7Nf0JkMpzxOICs3y5ApQRc843EcaPZ4EvNHDOt5a/CygN/uiGNFjx
+UipxytazidkhS1rxuw0W9hXr5lYhqdKH+8wVWcWNK7YtIDwNfC4QusuxksYB61n4SGlAxEN+L3u
MaQWleYgkgT9ay0wXK0IufFoARirvCdQAbv1f/FA6tTkWJsCxQyiuKBA6U7QkX7hFQA/1H+C7wJx
j1ybdX6wBXxeISaouoB7d8lAt/hRPXju3b+k7znoR3O91hJlXs/cwyV4DzZNFK6vHUzweqy5EXEb
zv7uKQLzTpb+Qar9Sf8j2QAFYZp11yU3A0dZcVLhOuHiCYRIpZUNdn3QmYGAHnw70qEWuzHVlNh/
C6MyFNl2swqQhvzn5vvI50PMwmaqbIb2EizoDYi3J8KTst8RJMOiRf4SY5J2XzldXMlXnSCBufIo
cryN6MucUSXZMUUTEo8BvfNFTgY4hWD0TzOE8i5ynC4pPBk2Ti/5tHnV4yVk124CoyaicWyNhB8R
qoVjiyuaA4/zlNfv2TKmkedBPY0rFDrEk063YCoYVfSywRdfIDgdzFIgvfZaML0Q3XteZLOAK5MB
8EKwCfXuidQNVUEHJzEyksp7+ofgdlg1xLPiGrQOahvXDJDlO+vAwiy98ie50AhdQcI7jCnU7Rdn
gVqUowgJUiPI4+mV+8qpknK1QEvAlF3ly9IQBENU4OpfWp2rPxMPwX79wCPvszD5MHIwO3xbHrVj
lPiT50vVXHc3KOojMJcdWlD8ZF8lF7mWo/inpWh2NV1cybVdxNyg1FA0dZtS6yLcU9qCySlGl+T+
sBwqW199tKQkVQCxaGCp98vi9E2GUUWbtzd8ip+5USTY3FxvLzcfDPaOdGCv7kFgOs0wX30bqSG2
BNm8AdYwo9ZQ1DMU8N0nDcXXAQ48Xvfayln7QMS1QlIf9oEOywy5UPhauE5oIG5sVmLrAYvJw5V0
N3GacMUmSeY7c7xMflea2LPZVdVHA/+k8vcxwrnUt3PYIvywg+zmjqKeH4RP4rFJ+oUAhxPhDB05
wEGaYcV2BAqyCe8r8TD/u0tCl1D3GLd3iefVxx2UGSWyRhJrphHA92DYnT6ZlwOmKvJph7Kf7exF
PH7pXgk4s1ImOt0faxonKbiUnHKW2vvijaQeZHAkN3hsaoOmod2wyKefIROLvP8hnRinyYDH+Qi/
9b1kKHUG9B1ifCszz59BFYdyHhc6zR/a8y6e2ckcmR9xyNiZ1/+53gEe9NksePBkOCCt7us2v4R4
De2QIOnljI2IA8riU1Em3wyfuJ51+IFttkBhgw7F0Y61RWdBWgpmj7h/pAzuepekjhqa8+SR6YNg
ecv6v560XOiPw1STVRaTv6Z7wg4tyK3hKggPM7jwRf2hzj5bX7fF4JVTKwXowDtACkeybg/RHaQj
dJ3cXLduHpNEAlIwvuxenC9O5XOwqRejFdGLNfbLKuZAAIYokP/ppLUzQDz67ewJTQGRnjxdyqrB
4+KaJAN0xYn3M75rhIicFoJriBaVetVXZ/+I//fsDK2CJut27RS0g53QOR71OxgQLoTtIH52uled
8G2HD+1Pv2xCzxxLMIymdYpsucusowaptsZEq2/NwyFirvPizUqZJwOh00HIlAaAV6OHui5kwL2E
MwjxHeh7+qXNkvU3GWM3ze3/QDr1/B7qJQom9qimnze8IhzDRlQFWQztCO1BmQhkH7huSI6qj9ek
Cr82Wc+MtUIWGOn9aaBpI8Ekeij01eJuz+GVt/0Mcrvth+5bRtwdIWp1jHht9xQ2HBLAGKgANNwt
LxZrKC7Kq84oQY2utLPCFC8P5KsDBulh4ep7pFSpYe4lYG91jRsU9MYb4o30JOFYoDErs+XBd8CP
fNy2X4hng1VsLXCeMjbq1sgl5szO2b/VjvcBVKGRzejIVeFMIJVE7TO3Ct/j01M+p13tVE2VEhnM
HSpEDiTpy0l11Gg/lZgYum471CdhsKOZc4SJtz8WyYLwSbpd+nsb/IKrVhtx17i0xDfEfwCUZNF8
Ohf/IT74lp5wRI+HDhcAV7/A/9y59rK35u9WtxNive91E1yMiJ3MSQQmnWhYMMXot3shOrSrOlk7
sAnpRQW+QIwPJog9S6DL91/t/djFZerH1Wy8E+D1c1qguujZc1PlCAHpsCzC0vrZDIU51RYmrCGp
Ku1l2eOUdWbJ0TSH8WGVh4mZ0L5FjK3JxFM/YqCaLlP40TTtV9Fb1vPshZ3w6zzlUVdYJw38yfCz
TVvSeTBM939+rp+7CI4BsaKTZ7uFwxpaP/lT4i3RfMvhSrC9Z+Id0wtLdULm2yZ80LF8+esyHhsq
83dT297Das3zd7JvSKurUIuglCqxISxMQgHFHDI72RVUYl2X52E/4bZhgVfTCr0u8YO/lTY2DQ+4
6jCl1kBP9uu2R2Tw9GFKwKwbk9n0TgZDnf23zJ/xnHCZ4zPlkzLh0o6s2uZaBZ+YGrYa/bdnM7Wj
Nc5sQRbPE9HjlQUA4ajy5aYhrb0RGBM+YJDg+M7Joly890BGNhSVgujGFCqOWqJAAJ4Bm8szwWRc
qVJH2f0+HOJBo7Vm0H3LkHtz0DwFffzNEzjJMkKIC9qIZV/fvt6QzAk0FIoqrhV/NlvxtNcFT8vs
mumXJHbZAnXR8oHOum7BFYvUyfQ1A6LQuq0DacWt+gQTn8FGh2vFMO8FvCvZ6BJ0r6PEKxrLQEZv
HzTubyKIDThP2lhYk58G40pat5TidLVY0IIj3N5md0zkRnDxmS0kEr9+hf5SdLgPCe5SPh4WyWmz
C15jqfAv4t/p/B2q1xy+TlRJHkGjSrglFlW/dXTlT0YfyGUlt8cwrIyi/JQv4mubM9BdMLrWJdhG
TN8G10YrEzT79WO+32LLFAur6OxiOMEU2YYy6LqreIAwCAhsehRsgCoqIboXU9BL4CRXa9zVuzof
s7hrRYx7sOG3x7/2MgzRYaohLmQbcvS0yN5dFhrHknlLzTDroUMNt4eTpi3KRv1wuRvxJs8hNGTK
jAvrWSCGylTPg+POqN3moB3eU8qooVYdB7YCgtW6epzUaV/UNBfjrlHkDbMI6dtW7B12xdgFRjNX
Uz1yZBjRBl/YAiUwAcHDpnUlEJpQ3kBAqcGjcon43Ak61+3zXkQXDVxD4HU7qrKXtFSAF2ztD/aH
k6ikkP+p2SFiNWXhVG5csHfCNHnj7QNi8f90ZvnOE4VILW0Q9KJedCBsYwQzUPOheBrO6sj4Wl4u
YSWpB/BkgeNrsfypmVXXYtBFnl9w59gTqRWtlZ2yKqH8/QcPfSXFogIZE1Mqr0YF3uTHH2sdwNG3
N0wbV3JhZq95ANd7KdQcWkPHk4xQw4r9HI/S08rhBCMNH5zz6t8uUMdVurD6FJemuPOMVSa9v/ZL
5BGJZ6ul2bSQw+uuxw5YJZbeWfAv2SpBiLRhZ8NgS5b9BY+0d7DK8mIGyWyw+qhM+Veig9vCeu6a
f/NpbSgwCw62VknjNJ2T+WQfIOHYyfPRtYd9adsAwgoy8nCTICgDITaLohTxP6Rd7W9G951ZOENK
2+OhJOl26MYWbKbTwQYrhYfriEKAaxmU1dV0a2wdMc0UsmruI2mHy/yXUwBbZXUjxh8GcQDq1XZu
6Praep0HteWO1TF0Q07eF/U56fwf0lA1C4bdODj5QVFDl7CQC9lRCPhM9GoJI5v4FlNY/fnIiU/6
lsp2lVM5JetutVL63Hb+L5IKWumDQAWojxXgCnWB5miAoZ6e2Vid5zqHCwZ59W5NcXNX09bqkxRM
9Haah1hfUPGPTRTRYXM99ccd/hs+O131EN65w6xFX/mnX4iDEpsouoIdN+al7W0qNUBuHD9NjkFC
IXjWy0z5IUnkuAvIM0450CVeSbX5oDAIiyoR3Oz9OPDCdmDV0IccL7H1Z30Bat/5nokJzTd/aYeo
XtvNBvdjoAy04hyRstVcy1a8lxz0CIq9zrcQCXfFe9vPuDBQCwa9HeLzrysF8aHA1avmOCRMrViD
mRwcd+dB1TCE8sSrnVMEn6NuQr25nt16Dye0YRKhge+/HdpjTo/xiFpb/ySc8PK93FO37zOKPRku
2LTCiRUS+LJfuTo5JwVB8ZybvqNtC2J8Or0xyFPyH7e11HwKth+Bm923kTASQfc+c3r3tzS9ILo9
mxaXNngaXX/D4kDJk/y/jxFlQ96q6E1vLHcBMeOkcH514h+u3w8qtVeUuOo36meoy/hMZRVaobkY
9TxTr30O3FQoZZxH5VN+P3ZL487XSrumhwI+3r1cHxK430QMX6HVVqGq6++J8Kv9R96iKNkpYzO7
dRApUM/ykaKbOl5fIQRJdsIES40FefsrQBmknM7oy/oMT2Und0hlmr2veteXwEUP0TBC9VI6YFRq
I+nOSamHJfCWY9AB9yku+JLLeIqZszDbQionNL54fRw7B0l5oQdLL27RH+x0hs0pc04zMkGM+M2a
sQ0n4sTK29XsO0HaxIb2x0JZ5CN0Q3AtSzW81SKUY9b1zmP3mIu3JnrQh0YDw2OCG+PB7J2HOIvq
MdbOLWzYibtyQFKP1kuFeyefz9jKVW61Rq31ue2B6y7v2rLb+59S+nXQRBUyJhkVREXor98rmI/g
uiOlRugdbyZm7UMimLhasGK2tEQx0+bqr/fv15N2XDbx0L5MTGYJqSLssWYAHm+2MDHS8/yR+JF0
b88WL851caZZ6mYTqhHFgVlg7A7/7GQAURubcukK3YLZAJT9LBKqa8vOdgtj3N0gDWnz4mpcts2v
WTnpB34X+wfR4y2Bo7bke35i3gPqHZem8UD2G5lmeY9uTTb7B9AoQ3nf53NsSAMJjMGFmtTVMl0H
K5rA+BWAcj03qTD5Fk34A/G7GDdkS8wPSmMj4Jp5wLzdV7K+SMXl9o3LopIKOlO5RQFCtqYTuKbt
+nSEyFiiD6mki0lMvtFxhwdqkuc9Jfy2FZb79wOJcWtv6QPPLpFbYsUvLk9IykK2shvfh2ZJqaCr
HlpsLi4zn7UQwWV/r+N6ohYQbzbq5IbLQ9XxHjmSlMVpd5OHcnVWDsC2P4HdVqP/lDnU5DmcunH6
0Tz3sbX+3hJRYGQ8VCNwUvsqiwO2SAdBkI1aTgC1LBD6lpcwEaR8wXjiZwddyO/u6LGNx+Gj39hj
D6x9oa8TP8DBiA3Sns1mqbrKftEmjrfl6D1ORE/WfQkCFQO8R8DSRTnoSrdk0zV/Q/48H4hO/fQ1
LRLp61fDGD/BW/xN7wEyqzmBtI5iOisA+0aKVit3nmhXW+Zqo8Cmw+Qj+z3bLTg7r6RzIgOQlxmq
f3tdvMsIDayevTyvcg8AHgvY5SD7jms/kEyeKqtSTEyObaUvd9cGlJeNMSCOpgDuatmX40sacvo/
ZTYMSqZUiT9aHxMW9WEiZMMZRMzJuk2Czvz3AiUHkAW9UN8Jh/i/D3Cf1ChY3LYzXLyOiHZ+4Ch7
Iu6RfzlqWWAdpIQ/vOdr8uQtM3ZZ99WCNV1dMFlTk745OE3+lZ+indO3fvtfy9PZni27BJvuZwW1
VISCZAy7WM61aAFtL/WoCUQeDR1Rg7wRcRRNnqnPFU6RLaCcRhvvNOKi+eqmSmNItNTsfcz976b9
GsA0smTK3JaTfvJIXX+rzFfX6wkiG+4fnrwgXPLh9j0y0Ey8M3aP0ckjBOX/jX4vQJsI+qozsdIz
ggKQNOvVhmQAapNk0XHIFPU9AXstgkij++M8+yOLxELT9MtgHT3TJve4s79lT6K7cP4NY0LfpIhq
hdkMsrRTpqRArAiIoWiXR4Ky3ZYU+YVluqTySAGCD7y050ziDH688TNRgYx33SDbl+pOxEsLyN5H
epxCPa7OKbVRWgJXL3OvJe5L4J2nEkMNZPH22MhP4hd5PsIX+ru0h4YCQ7bN+yhb7r2XG7CUZOts
W9qqzRoRdjsU3+VeoX6N8FZLqsUgwmIcicWx198DRgyimlOiQJ9MTxLKy3K8fPitMZY0t+6CvjWA
8FmvHDyPLCbZeBDFUiHwZxry1NZj8pBl0tWcQFSTlQoj2SKk7VxIpI3zW7tlyaij6FsSYOGmpxHa
vUEQhckHlJRiMiCvvAZhGwD1wKwdRZxR2vCZGMQVXsUNbfBiY3M4I2yNrZzLKu1c1WbH4v42ZfHR
6Op56qlK1gSFJabc8ik73Fw3Zuk9Oe2xaUImugDpUtGmnu8+IIH26HNHDgJn5nw7XP/OVvg+ztO/
QT6stFL9WlA+iV5Fu9u3pcRdDh08WMhbY3DdSB6v3H9wgpZo7clx+kqKpTVqobMjelqYVT1xq9dp
e8s8jfaFi5u0G7D/pBnszpJJjYAab4cTf9bD+eYQhygdE8FMjRTi/R22ueI1FDj+kr3p+L2N4+AW
24Mr6xt0zV3PsyptbM+a4bFLL9gEZcwGPyxdn1kfBKaY3+bk1/PLRqn0DFcr0Ys18S6S+LhXXiD/
RhE6wPcjfsaukV4VowEurGBhmm6Ptuof6fBpPFhxZRvk8yqFx6hNmjFmvRr/+yLNekJX4X4YOI03
yEEFScvuXDAaPIwJwtGL0Oz0AORTb2myfjrHgaUzjxISl6CO+uS0Ym1naj/ai2+SSfiG6oxRneS7
MPzuJJFDyHBEUv6bc3jgQSqtuzJRwud7IetbdAGiEHoyK0ejmZfuR/NBVv+zh6zi2AyDzgqfgeRK
4iYhJpUfABUu0gjHvjy79Qh5W2x1sN571z68uylUzKPm58+PPLqLmVOPwboQA7WLvdVO/tq0vzaj
wtWY6hWesl5W5HVFlAkI+mD/qCEKNLN4F+b6JhQgTo41XJ+cOoefX9biLYdKaJVUL/9W0ysFxBKo
JmskzVKqQ8nswNJSOBaFR4e0JPHrfCWUA1PS+OMX+Lczl0rDR3k9p7BmHlLLWoC9FNCgvNFu0tg/
HA3Z0lw6hpFi6cQRcUmO/fHFbzkM8gurPy8w51ZHaTAXWv+I6RCuB39L27lCXyVg9Mbjhe5NatYl
0aFW54vrKUHPql2EdD1qnfv4ThcG/+npbzxrGeDdwTNxT6YvxnRD2I1FeZCiKWij5hBibZG0SMCP
JzXNw+3xWtw64gyGVbPGlqJMvN9os/TUzO1hdpbpSHtk/rEEKeO0x51WQ/HesCqMw3VjL/JtYM46
32Kkdkq9dmvI+VmfK3TcSsxeTB8ZIfHZKpeUBXJddxWrI5466BccVHuq/ayupTA9SN7eTMcfOzvf
qojIfgyH8OeHhHLGkzOTxffQGKibrFI24tMvTLz1t8OG67vK8MUNM3pFDFkFS0pkD5Y57YzhHu1D
8zGImmeLrl6BZVX3Xi2YBWfPSuftn2ywWGTjuT+k3oNb/FZVz2A006aEpqfOikTcreMYJRVEHrbL
Z9O8iuaz04X42MGrxGOqzS6g9GNoHFabNaRizZLungAs1A7cnYNgd5uc3h9zWo2NkFjVUogmTzyh
HrKOahFyI5Q4wJS7nf02EAcy02hIozxB98mai9N9q7MlrDEmca+XRVh2AltO+TIoCUVIr1UdMAax
k5DSgkp8iShvQbsrLnSSLcHWtyZSg0q+U0in93LlIrlYMa6NA8oCAYNuQcM0+OuD4R8j2QMYByoA
+s8e5XXn99SnAQlYAauuPYuM8ZL4OvhdoFMRGhK/povkjjoa4M7HxZnThUUNCaJ7Sm8Ktf2yjLw3
8VkXFFoVwlQpLrBws+kQokHxYcImXfD/PQM8KSqurLJvGHmhDFn6INQxXCHwYnt+6TcTnc6YCAHW
LdSOlHITuvj7J+fucM/+UHkn8c9a0RM5UdvuuW1GLpZBA8KgptI1xWKfx5hImsYIIkQOvs9DxuNN
7xdJ2ezOcgShv6oys7ddMUBMBde7j4sE2MeLw/iluJ3ZOxXy/1mWGPtRH96/rHuNOoI/NB+kAYiW
drtDyAUsS7z1qv6GEqefWzdAbJ2sD8+kOpES04mKEdbJMUuzs9W/fDduM0mF9LZadd0Xz6jbewgi
Xe9G1e6bAsopSOrbNvNXpkA54GgUVDPz6d9BhhQa6mgHFZ76vY/yKanRxxRHTD0u6p/OfiOZV5oE
SjglmcKe2Sc/xUZjww30kkxUmbPzr3pc3PHstN5fc2xb3152Ev6k4a9rpLwNecTPFBq9W7ue/A/E
CUv3UkgS4sHU+YV1Jy0VlrMlO3Sr4oOS+01sSzoo5s0nD3nOogpmBRltiBLHBfbVb3XxqdVQqhm3
dVZBoJajS15yubF5usOUg226Yb34y5Rij7Qqw5XSQzINXslvG4n33gfpZwhb55SlhbhEMI48J7QE
AMAIcER2kDIcixKBmcO9fI4NIaK8d6IG0AVNB+S/vUBZtnHzdKVYzPfAXsGsskv3bB1oYwcL3xl6
2lP4sW1D6K4Ty7BlyiKxAM4F4V2eT7TjHAxoaY0ycyg2BwCTYmPnhk5KYr5NscZ54DqKBwkr/iBp
rxLSggzFOpc+g3bq1eUoYtke4pSGTeMgUjM2gL2HVrkpNiI9gkJR0aazazfufA4S8zSm9TLJKOAY
gOEI+LH6NI6mHRAS+z8hMrZNx6q7rLQmZe9sb+0mwcR+pqBCkLyU8TUbHQezf5ByuT+zggoUXXxN
0EcNjCZtPF6jUPVnN09nuxU08rYkJce/mGErkou6t+xnce4Mi/SkwfuPJnY0oY6f8vLnARIJFobP
vvgRJML8jAcmi8pK5cxI5Ajz7nen1k6cIwsp+LrueG4CGqta5vQoZbWIACW/H55dkYvhukbtAxDK
Ficq//3LxFW6Uc4qGgwSX4LgTYaxD4ujdOgZ5LrBJxVrDKbB8s2QJoLHg/1MNLm5FFgVs4uUw8ih
OoRePwA5Jkaql/wemIEOgQFNjsXxXFcVrMxPtTqcneCuGEpRqUV+BfeGAsuaRo/EpNvQzDV4uBUi
MH4DE/auC7KZhAsxbA0i5AWROrHvmkI18pfdjWTYm8nV4dvhN/M43d0YCEgOlF+V58r+FUs7zWh+
iqiJ8w0TGOD2wGFEfdUwDm1Efou6BL+4bIIJFMOpQUah0e6D0pHBbji6NmUl49nbTfb0GeTARzg1
4dx5Yv4R+FJQN3MQPwzOSx7B8eM6ur4c8L1QnpjOmJ/4jMqmrY49KAdVQ1InMq1/bZkL+KleMZw8
e9N0NCjzcsbdvo1tMwylPYlcHs0Sju/Dq/4bimta8/pQr1wEAZK0GdKNAfNpmivc+r4u1jmV1VAr
PjtxEyAXmoOUqqGoqXVLKIuDLTON33pFpngneYKh0o36URR5Gmy8k61EBIaf8qnQxAhsUMh9ftVW
RDnrbmb0JdLy8KZ1j+gGTiPbbIkZdjiFXM0A1DYZUnOwn4kPbGId3ltUgz85gqC4PL+wr6QLGDwg
AKIrYE1aaiESg30RP7YwoML4RQSwdp94H4+8Upklzllab03oOg4tv+Ir5aWq/r3lRiEI8on6N9ZM
OZNIVRBM82Cn7YIRV1tyYun5zbHgYycZthacJsQ1Y9Nlf8wBrTeyY6+WRlfmIRY9hhNnLrVlXNbx
5qdKnFoLS5/z2mptfq2jOgCvrZHYyKnTixX7nKSOjyVZtEUuldC0c+tJJC9BFvgw76CfJqGgQyHZ
r+bJrzIodndzSqcNLGm3LC8Ud7+I+sulbgYEQxFff24eTeN0V+2Qa4ZUa5uia9p8gzvYPxtXmhP+
N3BKssGhku8ewP5znxMpxGX+lA45uVbKHmyy2LK4K6iYG/Ri7d6EJzg59hPMrxjfFkxgYBYDl3bo
Ao+EvotP2YYuVDDTJSKNBJqvTs0ZXL+ccD7ufmbNfRsf9wYy+ASFpUee9LztEtz2iIceTGacpi/L
x1YhI87VTgv3yP9dCbWMckdW2EghFQUlBHLtOe/ops2MVS31RrGfLuMkxnnWnh/c8Q84qqxEYT53
1AHP1lgzaTIwijUIL6/uQb8enG6EXIsP77YlTTi81MT238Yy3UzJe3EmuPKgk1P3WBRvVPMl2/Mg
V1OZrYCuck6HQoS2+IRFbNcPPzLgHz5lFCWtQicP2t8uZtiYLjkkBI2175mXfQ9sD6/dPd+Thad/
fL7e0IlOr56tZqyJ4Fd7jrs4iywnYpNJy7j0nbmg4wtZcWoW7YIG3qsxsus6qvK/8ttw6FLfF2xx
bTiy/M8oY7nGXns/bDR4VtlQWvBPBEJ+1GIEHUvdkfIo3FkvsyjQVbxZwz/PkUAYNk4rz3hhnlW+
kfqnfGVrqledl2amVALlRb8teehkFsIgNzj990mSmWpzkEtKT0Af/kXta8LWa/tUO5q6oDlTFbON
1gdx2o9xdVrFrHAjqnjYkKpx1zXbvNbKVryjNI9iWW+txEBiFaZjtQLl2nfyB3nROJbHj4P7yhCJ
orNpUzae28zvA8oDvOyVAgu1CKGbyvL0l2i6uV7Mndu5ms85zhLLPbRjGZh02Jt4bFiAPC/8i/QB
xyqdDevPCUn9n3vPBb32aFcNo5jNFIx1wUrwuK8KD6na/moj1Lt0A/xUreTt1JRa7DzEI5TPpXSU
Fvm21Bl5SgdRzAaPhMGrSjwvS6Jcq0FNb51gdqj3yeD7C0EgR9Si6IKsv96GWdAlHZ/gJd3oDRu7
B9IExNRT1Qm+DCMWVlZzkkysLhZEV7flAptkXnRsu+YOXUsnqaGYFG/xMjIFfNYEoa2YBaLUGcZe
FFSquLSnEfYDCvDPVaW+3qukH1t3qO6xbLXImC+y1DuO3wZyIK1XuyxxCbidcD0D9WCWPIaShFU0
Dz3Ll+xVCurkxPy/LnMiHKw7krrUfPXuQyxsFj/yWIvFqUD2TTWvKqmLnQ1LHBvvKVJwZ78C50LR
TqEFuaWfrq/x/ON8C2Z5k3z9TTXPQKVvf37EJORSH3k5i8pyy2FRQ7TrmIvyx53Ktw5mRke4W8Lu
N0fflaotmXKsxhPwvKf2Fg4SG0KIqo0CbbNofN4Otsa1WJwFxDSl7b5mVqStwd8TCsJhOzkcLkWw
KzfoLO7vOFpkVegqsCFxf+9BZWG8ByZ/drtZRrK9OaK4pDp64TdGoqiEnCgDzXEYdimy49XF4/gW
+8vmJg3MjhbzI0oxNJ+m4/u+bZOwmnuJ9HIbsCYenO56bl8hcPkrkJgEtr/H7Nm/0no0AjdpCnE/
BP/+FsTe4qZxgJP/L+LPX5iY0II64OcFZbGN0MdvwGUAxpjnynwE+nqbu3wZUlihbYMTmrdO83vh
VtU+Vb9KS0FurloPMrfRO2UYQy2/+dr35e/ZIDDALzNIdhP1iWCnIJCmSFACaRd6FR68NUE83lbL
rFTziZf8KoXi8CQNoUAW2hxL8wvk4+61tUJE0HklxsYQQ7HysiJoTkn6yKKWevruv1IpVqHPtMLK
5aGZ7uM9cA1/FD/kou5pV6uh2Rpm6WHl+a919A3OZ1iyFqz6Mn5hF1E+BtS1cfkwTBJ/mcY0Xl4K
goj2dhUnFd1jo1HLZ3veLrto7KiU+OnESpK/hXtmizSv/ASwss9uPYHKwpvm3lRbymaefZ6O9ye2
JHYu8VLkPBPRmFW/5qxnf+7cIi9Lby+2kSEX9rwXXbHuZznKkoNRcx6drpy/QNif710nPE8c6JrG
xXbuHFmNj9bYZ+HSe/02bmn2EJl+u41+xKW/ACt1VHTcLlM76MRg3v/ZzoONDbHe96Gy7hNQreaY
qdkH1FwS9DPT5is8inXr/9wYJSEce0Dq69tls15yjEfp5SBDhA9mxHjCSdWRud1wdL80Gd0wwNRU
w3MBBRXe6AiIJw7+8X9qMJl/fs8MmzCWzWeadTAV+zNwssl4WQDGM1vQ2x5sBZy/c/SdrlIGOzCu
w2kcrgbuQnigjqMAQQsjM0moACm70fePDBXxsKR/hMKrEuq8dRb50Q70jb6hHR+JkIDkVYcTUcGi
PYinMDedQGZaaL1wl7PAR9yo9l8mGPJ1OkIGkIAninAnjWIxFWpNBcSbEB58chhbx8D38DjWIkCT
tvmq/1euyn6cTW8vb8YrBQtRyhHNEYsJLO73+hUMDoK9GyHI4x/RbCmUWk5Hk+J4V3H4b6T2ft1u
XwAKJVhmGGGii9zUr8HTKFaoDmB597WVoMCJ4AO//E4AHGgLoKE1utmlTXrq0vzCrsAvjfKOV/Od
oy+G9QK02KwatNSpZTuttrKxjU13AIWSqcygg/qKLQbI23JcsaEpwfwjHtDWWOgD1Y9waVp8DrId
OwNS8PEDxRJmNw5FQNyOho/0UoasPgDKmYea8YaVJ0twoQHdwriH9+/WlRJb4w4XZAQWjCckKtkp
ACK1kg2h63B6VyvTaj/PLubPkfijlqgoZ+sxzwbiU3a0wi0s/ki81ySnopaN1gqQGB78oxxGFRCV
Uy6oq+9teVhikXoLNDcQHk5BeRNgeJx5qcBFdkSo0nxgljGVgjD6/n3XHSaD98hU+/u5ta36iE34
mWS2riHbr6jPFyTs2dAZHYV1Qq+rmjVP/NNAvr8N0S+tWllmbzLrxPk8Uf1JDQAXphb32roz8l8i
mEVVed++GFpxtq0/t2ppgaVpTQcfin8vFQzV8YqDSqIQSoxP27XM6sRLcqJ2XH8JE/M9wXyg8rJ0
AXqbEskm284RWV0W6gUX1e5QEQlqxYdMGg4DJD2HUqMbCD0rjxGAzRExp2D7Wf0lG0JpKlaPbB8n
XbSJUvOeWpMq010VUqfFXYOGIi9bU1x4I/rI3dUryly0fSNT0ZC6EobJgCXCW+ad8WyyAVqL8+ar
PbIhldmTdaQFplwPk6yDnlESTQDgWkRuf66GNBJggQD/M2UsRgb4B2HX/dHLlHg1U9ozSnpXHVwI
CDlpQLkstGvBT0vtFPNF86TKwdn+F8bmKeihX4gZ453OhE7s8pvftcLR+HNfX7NKJ5MsOqWvpnjb
mvl31cLicuLJXHxbyFxCOdnmrdtYb/MS3pkQ3Ub6ucWX1XgQfaT2UDrkXx0n9WKfL4SzueHnOIKu
YDKEGQysKlTlTuCeHvJxfU4/GUu/ulLO5A7rmFPyVZEgw0Z4TPQpylg/If0uCsH2zR/0uTQLfnnr
7Ur/d/R73ezdRLLm5FkB01efEv8g2trVLRwK2N92CmeQfT4V2PWO4W4a4qR1If3oPbhq8S1FgZ83
621OSg3ZzKEIBH2GPoVUA9Aoe2d1i5t/Nfja5vCdLzcczY5NIo7n1bQc+oEqYRUCuQTSyOUv1TnF
S3HKdcCX4iRNLr9Q4r+i0VTjFYu8SpcLSdh//rtiAo7ZJ6D1RJBL5tYNM/tJMVNpvFVtAgyxKNov
YUTi6rgTsuPqNBnbDXiELaBlJ6HDigoWgy333+0piBrE9p1PGPcC+nRcTbdi3NGazbkeUJqCY2RK
J8OmhJIcmW8GdMgoa2WGa+CajpVsRjldsHV46gaIZFyIvVMd0gDwNfFmc+Qy84MQQJeVkqzZ6GKq
GTPn+5kr7W1+ES6oLGGOx29ltitdUEKLaUV7fyc6wBJq5daBii/VcuppSNRzK9ZIiYwXrV6NXnse
wZ5CM6fLgb5zXto9AjYWPrCQu6mjip7ICWJtYAcdnMjZbifi5MVzKMzr7j6qUufF8nGJSZPguvf6
XVOkhXyIfTbtoAKqoNJR/jIUURQkPm/ga93ZL+AZc3fBil7+8gQppOTukfK92RtKvdUMfig00+7c
QVeJ2OO5S+m/3XNc2A8sMDtnPWE6RoXR3ke/76NTaa8ynI6VifuB7BAow5VSeqaRf7w9ufvf7OIu
8MTDcDqSKHMZAzEoUKBV1GmwbC5pkvgC+dZ2X00tcdC9s6g3v8vignYmkfKx7iz6Pn4Dn30LvRCt
aJezKa/ztevAEj+lzMDwPuhNLNtaR2ZkoQCT880AFqel8UleDeMNXHdMdkxosofHe6tZZfVTLBth
hasKGC6lr+O0ByvnaS6nqkEE5k6woHQ4pJ+2wR66u3VQntVH58iaiZd3siSxpCTfzbBvnH81iUUX
GQ0xFovIywLx8PRi+C+3vI4ohe7Qeu2VG8SPDG/gRTQpGq1FQ07ruJHVYpMIBnwb3E2rrfb9Asb5
rf1JSXs9G3W3nVufyeUjRO6YDlGTltNlyBBsj5h5Qmgpme/aJ71N5rr/4YffQGrLp8lWdM0T3SUO
61qkG/B4nayKaul5KIM5npLdLvHsvNLVeSj+ksyRt96Pr7FzyWBiccx1h3cwvUTMUChFNLTqg923
/y9kmhVp2s4MPdraouMwZrKUjX3Fi72lzB5pMDVIyahu45WmePMew3z8tjaLuMpxdK2V5W6yjh/s
HU7YUs+W37SXVyhp7PFDi+qTVKAn06AAIxSkxXM1GNRXO17S7wbyq8710trJm9+F3mjW+a2A9Pw9
zXM/mWage28AYkLBoTy1dbal9vR9B5McL0FHCVXy3yQTyCInWT2d8EwKZoJU7oj8XriAn/cjIib2
q9O7oCqVAvriHIqguspUN8A2V4GE5hhqEalAYUwsZZE/NCe9C/IebMVr1p7qTtHEiQThxkvmJS9Y
LVMgrV2j4cgV2UHyuJBzosqTjWs5pOSbnI83eowKTIVHKFhMT/9fRvzRCNXmhbLXLkn3qXkVF7IY
hnWWNgAfwvZcQI7RSV3dsBBKISlL45E6cF5pzQYL3l66px8XVJ0jl4Lp10t8IUOWm+dUfkFiCEOP
FUYT5SuT9dDnXg3Tu8I87uQu/WkDWp+MFLV+9XDDcQsIKNJOXksj+ETu8CXXsEIALLLbFKdanCW7
35cFtNxxwAFeMx78aGg1LrkP5fhH6Jz/LkzWOB5e+QB05HqcjcXyaQ7uOhgVgsuP3GvDZm4ea94z
tXQhB7hguJwPMFw7H/u9muhc1gtroS+e3eag6MWj6Pq9ZeTZE7MmqdofgWnvVBzuaAfUiwXzwSrF
8yedOKAIWRwFhLiGt6hkhPizga0UmpSHHaMcMPudFO2bDEECimk9bIxHyT09bBthwdiDe5VZzL+n
MXc9adot3sxR2hjJpK20gFC2zjk/adSY6hlq7MiLu0CqImJCewZf9vQURwOKL46TfHFvPxJDDJGb
iF88S5XzcJO0W4OSUtskunsHV6TMUr+A80fUAR00f0SFHplj6l30/IZ3PhpwKFPRoOxvBOMojQUS
xW3D1vklCie53vHRAYMF/UunkynZBcsnlfkHRiSIKRPMgMBlqBlXyDzrQOGY803EHhoRiCzrr0Q9
mA1sSh0IsoQELWimIQD+NrQdSdpVSmxfeUz5s6HsYx4JuXrS65XfnMb56VkkeFXK/HuoxzDzpNPQ
Xt1b9SOLt4P9RCJ23u61CeXPPYRUGKY3rYzNRdyFoKmatTZkJ7vOIr8O2FTeuTZ5FcKEWWbTQoyO
ZpKXuoEJWaK7N766CbzsVIzCyIj+GDUQL/LDpf864ENGP8RecSKrzZSt6nFNWhAO8DoViVh99zMg
xqCdXJjW4xc7ngTMlwmtHaLf78Cqg3tXZFck6QuVm8eHC1RAseKKke8I3s7lNtguIUTxGyGy9rGu
YHlJLybjchYNNGqiUTYYLn/gF+9RtNUorTNBkTq8n0esmuJ+BxRLHHpYeZLpumpvV/eVRiGyu1OJ
xIZlENvmzzVG3eL1OyYiL0jNxnMLxby1lfJlECfuWHZAzVaV8zMSVsNYzcB88EusOwal+Lu2fLy+
gMs4wTBbwPEUcflPky8q2CkTqGJfKTpEqEAnDOIy9N4+j8jjhDUejwEvDPVzZBKQrUA8G4BuU26U
mAli/4nYcBM9NGvkHYHi6rIUzt8VXW1XGIgP3S21AtPGWZqvuYe8aH4UItTKU1ncPriF4gxqdML4
5m8Y0L27g/nRbGOL/T49Q2GA/70qpeUADYNGWwlc2AEXPyFvIfY+DpE6pbLWIXAvMjkxfsvjc0LD
vNlVgnZv4Ru4UWfxlPtryFQhSouYWm8kC9krzXFmfLHwmjhrLQCm0hAPZ8Eg9xw7eImwyCy5GRRW
VEJSB3oGTNm5tmM96Zt7CVk6GFXZlu+QIULNO93P5XHJDJbnfe//kvsrS/i1iU1yGLC3ytp1U8jQ
elpMcBG/Ekhh7Yfp7wbOD0iBh22fyu5ZX0fPHLW1F6Njs1I6iBKCl8lIp4fTeAhPIiSIiq5eECIC
tQSWNpoYjhpxMrfAiu43B/LylkI6/yy15FNWymq6cFkIRGh+fKYb2Xy1bEnaf0DcpOlGbGL28L75
x0NVMpdKsyV0PTVjm3aoaztMOdw4RcEOTexFt49yAEFJ1a4NNvmAojvLmsvE9a+YIEYerIqqWnnF
aim6aScGJrMBAN7m9OsmtdEty41XzbgUNbpF0vD0DKYkB+uCmrR4kpU8zInWBxAQMt0JLuFxXF8w
6Y2RbYKb0vHbX+eaWrj5FDnweAa/kdb52C6kwILJ1u9i6mVipNyuW0/IaLVB43QQZLiLsMhtQDRI
3GrP+/PZrEtgyJMX/WrFFed1amkPc98ERYJRi1LDQxVjy8LT5icMhpV6IdonO6Km1a9ychloypgm
Yb1vV5q4PAOlLc9ioQX+VDU98mxNP9xu6ZyVrzK0dCMNCNfo1WZuRF9BJ6DHtqsnBoz8M902trqm
/Or+2Yr+fh58de/l+y9tCMTBTzkJfTUG/9tlOIaFfn1OqCY+qEkk7Z61Cu/Z2184uLdWqghZjm3h
BLp2LYm6ZM7MJeIDyZ0FPY8JC8IM1Apr7n5A7v5lyGvjoIvyAs/bOMt/XiH03csxHb9Bdb/d6VjV
k2f71jbxWtYalGMi7IvLY7pZzLY7ecHmg7u0Kg5egDXvNb99Urk8XGlXhq9dHaEgSdwcIOmnzYDn
i5zdpZkQ90Os0Duyi2Q8Tb0VLPVFkoEzH5ArydASQGYE0MaBu/xdHQcYGgsPmVzPu+MF1fOv8XIk
gZF3WMck5Ffa+TzEnelG2hGLtb1pXaS/GNNQ0iac7qAUcGNSTUflDIFlrLr8fMKykYO0PWvXvBXI
kX4b9VlBzp/bvtrunmltufyp6MPj9Taou2Md7EFXj/BmGoV4+K6aFhugBXZIT4VWT5kngHpW+S7+
Ba4GxAFh1IgTamAofMGR6lzatYsTL49em1iEZ+Ha9zbbLDggEXldLi6/MWzCmS76coKYuHXl+4PH
OVl3r1TFcssEildeDNcpwABR62N2IfaR+XjwKP+EOM6q/MEu0gGc3NpKVPDxjjVCOoERtP8YShBj
jGUKstrHAoBOxNy0gooRQUWBa5eMLq5c+l5rVXBtJ9C3cmxWbjpbl594mDIZeQAXoxQgAdvKsCtm
D/I+8pntA+sYYy3cQti6P1Ro4xSIB4VCpZSxwiMdsCaLKYGwV050rt8647K9ktM93SAN7q8MdqAP
Xqs1dQgf+Dxv1yoItl0qPT7JcK05sv7p5VRZd2Nd9SStSrH7qVjbH0p4CNWF/dYy3F2MCHHjslT2
x3UUchn5+HoI1cfvNUZFhVPsjxPTSXmfIA7g6kG2hQjNokqhHWRuOEzRunBzp9fXLiL9OldiuJCQ
saPQDFKlB8vvm30jgHXuo9SKt1vBRgEWwIc5dB+0WZibMzInYZCxKmxEZe3EO9lJJHL0NOtKwtb4
sIx7mJFY+RstZ13sg6jOlkBuiZYrzhTF5+07PNihKsNJT3R02f7CmOE+TD/vWSnHEYnqnOvxtCr6
M4ezdS2oWCerbbutWetq2YK2dH0pQ0UDF6PfF4BTqwUVedIBn1SxYlD8yWlkPdTqJmhBMAFRynVO
WlcqtKes+XsVLwYwPb0zS6bHAcSP2IYxRdjQnDvF5mew8ku8+K37fEtltagSr85e39qg7hQsDySe
guzu1TtS2RzB8InizUveT45gw1UdgmaGP4HvkaXZ0+gQVjg/pWcR8Yp6xHyAETOnbTjuSB2l6DbQ
yWL2gB18HOGy7cL9OjL7wFRChojcnWYDecIkdrnAXDeQEx8OYmpBvpEFckmsc57ykZcMsyi4aFVw
bRAoebmc7m0j8wAOjPbxnQ2CrOTPkv4itk952b2t6xfWUi1I5vZRMGg2B5En/k2IRZF/LLuTA4am
Ms4s5tVEWLhAbXOMLNE5gsNBJfqJ137qLTjpQBz5fPhVa8v1HwzwEkqQwYgHJnzXLiHtVFzvn1mV
6M5l5X/ClfgKiuqNY5C1mPfJb+1e69acPuhPGuqlUTMm2kCxhAt5i3xj3ej9gNx4xwq4UOY1o1CV
VtnnK0BDETG8w1SFIO+NNx/d8AsxGjHIY/0MsT2GGFm7XI+fQxQeOe9xlkaJaCyd2KQLLP8H0YY4
qBu4+3u7ixlxcxlrCgTkxKvcd+N9UZTjjNzWvVpKPawPZrHcU0Zdv5EkXf2jNBRU+0XdOAC1X0Vy
tw8swivnjW2cQYfoGgONnWY1YSbQXREBCkdQjR8kNZ2uQYjZsrFZHSH6f+b2lD+U4itWE+GjDOmx
ueYfuVIGyZveyXzV4g5SYFRaDEpq0MnmCss0RjvLB7jVAuIwWVGmO+lP0DclMl8zHbz27oYhpLFH
rR4klO6SF3uQ5/gHI5TxQI7EezHK8ZHweq2YvRFCzxlnTcL91kwmSRJDNhITYyvs1hPsLUyqEEJh
yMG+si40zb+tuoaScy8zivzb+zjbR9dFmKAWtcWxHqGp+VKCz7Tqu9NN5ldqytvrrBMxvEBFkcgV
vca+H8w14D7ohB7XcuuesW0MRz+xYaFuL3GFEsL6BA40WDIgUfyIMbVc6S1R41+B/0dGHrScIozf
6MUd1PIjrjybVHmyByz71daALgfbDycLG7OuR29nAyASx743N/aVPy/XltkoN9AN6Wjob2njAGIU
dZWk5VDaKFQ61M75K7UFnaW6upkVctV+oQ89ePW6dUW5nHr19lD4mZo7fnqDaLvxYoyMCJVycjEm
LiGwCOkEOehx+GpkXxZ1/YLsJLmD0CqvLHMyroSRBepE6cQ91XL8mlmnJsZEQQM2HrjNZ7TSGuyZ
fEZCG8SGmdDBjLmd4KsH5mBubJs6bY3t67lB8BFGfogmDUUnZMI9ffwQhl+S9J4HDyiFnoxo/D8h
uk+i84OmU2ak1TBXG5R0oqn7xAyyIWcMZR7vM0IQzSZc9owo6og0tDiYIUCKNBZGz+rvpNWnLNaO
TH1v98C91YT+X1KpDBKg864Jf0C5WQT2s/fKf4HXevOnfcbQzkXKQtwaxXcR1rcNeUvoIGimAPEM
i84qL/SZ5V5QBVdwTwehk3pundp+9W+Seg4dTRAI7pw/v7rqGZ8B8bilE1+PY1mnlS9YpM/vc+vb
55bsCY/5V0J1SUTAIfqVv/piqtk5OwJemBF+/Ynk8reCRtNMHXgUuSJKaNTA9Ka/HgdORsHLzt1e
MOBbeK1P6bHpy27P1k3b4Agx7A+Tb5m8/OACICa1IJCujYitj1uNwwFG8aLGxCJlhOiQ/D8g7vkB
1Rdt604QR+O3EjSFc8dZZFiaKlYLob0W5IbQu+krGWMqR+y728X7kgbVlmINaqZvKeo/LaBUblBK
0oWBGLDenxt4q8oP8kPQYunVcHYPq8kWxv2EqDOT5xmmfr+H6xsNEgn9BMQGYnmjSxtSvXnOhvzf
Cu7KWdXhqoyckjY4ZMf8W+949ZoVHwLJJmR4X35YEj63oavuLKQ4T2uHfGD0Y/FgELZ6r9t2VbCf
Hnht7lY32w3KhuCXYYBHWLUbwye1rH1ELljuogWkicF77961IxMs5k/i78cZbltgaPw9UejMbQSD
VuHEaHQKRFNqj6jOBb9UGs2TDX5CEf8Niym3A7mN74V5+sn1EM84dLqZmhuKe1SW+ymzaAOhNx7Y
3JBCqD948Ig9ZqtIAWq2ODxobb4t986CSj/DdAGu1uHriE66idNufNCiW4VC6mHAf7WnDrdWaSrQ
4QeisMiijsKdASaJ6dVQfyAN+YcjM/EcLJUed8qN49mvdZllIXMQfhe63IqARPpSOZIr0vJJekNy
XQZC0mb8WHLc/D+dfoxgPXF8hOfbRnSEvdNBjbvzTKDGC2XCfLOY+o2/K3T505nxdyVOyIhw4yHC
iL+rNqnOlfzzMQxpstuoxUos+JRYDkkAfPq4oszUsJwrD80qApPPwK/2UzE40eAS7taSltLegGK6
m3Dnzi+oA0MVQK6ts3YsyaGYIKafg6FqeUkKKgwnkExBNTX7z+lPsCCaEea70fFsNwx07OZpgheh
ZFfSjB2Fp4QRT6jQ+nHPzljDfIwMpLvFnV43HV8urymPJ6Eh4/2lRSBi/5xVCuFrlchY7AYxYUUX
X1OcgJPRI6F2jjl3bTOz0NVVIHQPfiFf66pDG8Q60ffRfgdspt/MiTD7SFkgAni07Zkvq49P4ghq
vopj/3DGdANyEq8p0Hjsv2oAIRUvkt5JukuvGDbn9aq4j6zsVjOlgclvV9EYx7h6KQnQIs2lmIDl
zb7aQEkv4uXYieOrCjn4iB+2USau9l4WjQMdPTNz14xkHIQKAWRnTDQkNPqEzlyQQ0PFWAn16seC
BHT3VFqbD0z7vaiihoNjqjEekYlOnLZePVcWEskc0QTgrkEbG8+or58qYTmwlBZVjSs/sMj9DHYs
AYxHNrRC7bjqvHUOaygmVWS/zN/IuvhYMiEUF4qbJfHBXaZmNkU+Y4+4Cly92zj01IGFwnUGXMTT
cfdjarvAF/CjjhOXS28UiagYbVKk2Gw0hPYJd0/kpufWC8dT86S2c+XCzRX7yildze1+ZRMgasw4
PmCpPgSfd9M+pmtrLPWkCH8wrdsd6VDWRh8El4oky8eISPKmpzr33mzkyT/G5F88lRRfOQdwj5kb
xIuk+1Jl1tFPghjDgSk2CAsgMIHRJFbAP1Yjo3dkcyNFSf9HGRwyUXoi4MUjfBde8ROhvXpSDJrt
feR+RTNQLItyBWCLkKhLuWpNLv+lEIxG2fLlUbsuEjWB0/Ss+3491RlLne0ae5uPiCAcEzNyWcNj
2u9nYLokH0a2rQigqFNoKAcVjfwa00hDu4KtFdK7E763DB+KPOMO4H9XLzpsO8+KULZ+x84jL8BH
3zqrEfUeAfGlcKhEpojww2DAD93H4fn4R2EhjTQBJADSb8vCTKcqBPmkotXVBS98Z5LTSUZfA6K5
FrDcmIoZDkqOMAjt5c5rinetgXm9L7j/ubphhm2x/9I7yZ3XMxZ3of04mWCgO64gZMgaY+cLCann
q2vJaEBvp4NVFSah+4J7+VDZTm4tZhSDhBA4o98V+xcdYtVXoUf9IBIr7Ogfa7CvQPFtd2exURGR
Ujui0QYuhFAoN/zwSehmCVHXGUBYqeEPRudsND9hMPJekBrYSbNjMslu9hnTnVG4oqq7cElrjGJd
8Mx9z3d9HYpw4zkx6H9DCwV2I181R/bPbEomHyVOilYrfzHaTZhU7YxZc9d5vIjRfktGkuq/yc22
0p5Kotz7+IcB1wxIqvt4YR8c3ew8cpBH/8mb2ghXVsuNnLm/7Vh/Lk0Fc/ayYAT58eob+EAVvO0M
S9efL/V+fo4e3DdRgOv2LBhnOimoVbzFghL9hLLaXCTzL+ncgsufuK210NepvkoN2eYoAouUrb0O
3Mu1LmbUJviLuENDxV7X7Pa1C1V34W11Jv5yIGtBvMcu13OX6W36XdP3dv+gl9GgXLeGtYVrXq6o
d6Nd57DFqaIL8ERL8jDAmtuIQQtbZ3Qpu4x/ZNxGSgllMbTe+WWMvXRSRqkaMCPheQu0AAOBuRIQ
H6YCaEXnTAur1LZYEgxCbKV4Afi1714wNNr5yi/bmEPI9nUm4dSmCEQo/ul+SXYoepYNPF30XNDX
cKuuQTeb683qjWjoRXeQLzvMXfMu0dHNxiUFSBFVsHmtSl72L82AJ2fLjCZh6dh4ApTkm7d0TGF2
8asR1DgLQX13uEIEV0yNIZjIMOB5VdzmTO7Yoh16pph98Vf3tkPiDAIANtiPlax57GckaMvZJHwv
2Odpiaik/XBHhom5aYt6+DkaDc0YLE9lYoTUu1rHKBVfiATr8Xw2/8t40lethfWSu8C5X1r0RFDm
0HKC+p/Tm5ekBbU3FPxrB67vtb+WGZfhlnVg45bs5rGuhURanRBl8T5yYwvxaSPaeuIPgjL91vr/
pjw8q0tQHd7Hpe+Jf6F8NVveKkJotTRzmf5iFALg3vnL3QdFIVvOyOcvlxHKNYHUQckG1hI0IxdF
bS2jbrJBcdPmq+t3yjIB/PBWcqMPIoWmVTWDzPWSfESPeL7/FycTKr2c4Bv5ZwldxBV19suW0Neb
HrQYf/CwVWJk0cLCh5r07z5RSIy/9skFJLsT3n5tgtR+6ZYdXBvkZH3iAuKykVuzXoOaWpzZrysb
49jiLAdE7z1jGZ981eaWSxQ62KzQBxtb2KdLxSG5FQzLsGelxSD3RhHAWgdp5GM8SAifvtoMASho
dGAJrtyG1hKSq59PYgUxhkaJiwuY3DZTI0d/wWOyPuryLBg8FsKmGtqa3cEg0WLF301Nv+7yzbaR
t8cXvmsv6QS7YPoF9UT+6QiYK4H3GZu9ZSpoP1zhc4ncsTWth83gJWp0/rf+492tu4OwSqPoUglP
bqvR/Q3SRtwReLLnAtdJnW1okYUbNlD1v/D/DeFcS97jYtZy6dRCW6+bS9c9sJQoCpCBIgm4eDEW
xuMQUUTEnjB+k/yIXOyYQkC4eTNgaGu+V7FDnCe3XLsjnzV+/x/sqyUff+iDjjmN5FPpW8fkei6K
jsPMAykE4oaqJCoQgtUtu6SS96cwcXdt5MNLjJnFgrjD6y5eG9g9PmlI1ktNKsn8Z45MgYDouqsl
inUuV22CET02BVeLNeJ0DZuql+6W3ffEt8CF4U7jejU7r7Hx+pTd1uRlZyzF1GbeuyVRciuRoMSK
scML3DBIIMOGonL0imB0A7/b/TXrba5Bc12sdFKw6hHvbT6tZoIzYVr7qGJqno9TE3eEt0C6ZGHm
NeJkquzAVCr3iKIx3aCyGsUAXVASptok6hyXxT/xx5rT7OVkWnnVNF6Q9x1rvEGf+euuBX50f1B3
dLPR+952NRyj06YOjcGlw7bJy8XYbuWAc+w05bmMGSedBzACR+s5FTAqiRedr3ZUqjf7J66rSK+X
JT+GwWnvEs3G8J7IVfDLJxe7QYwA8BYQnbJgxitz6GUPQEf1VxyaJFSZLuWIpu++b9ABocjKj6T7
CZd+ptCzvv+VFcW+tDYG6py5GRY+Y0CIpI96yyf+jgJMYrsYmZ9cmjZ5x7TuosCAkIRFYNdH2R0q
k0YYpWqTopuslxhIfhod1uL52NlHp9gZlC/fSoOcwP18T1VWsgsnuCeXEuF/BZSkzKpS9r4V2wTn
Y6itz1zPv0Mb3uaheZ7Feai9eEKymBF93cjE6HBxOXjcNWX1Z0uXOL72p1QQ91anKKM98blbcl4L
0Uj7Omm00ui4jkrUPzU3jrVzuBA0+UuD9KxcfFR5lD/hJg4ma1/0R1jzR41bPSdSn1zbRNlIq0C8
MO8Chdcv6lEmA0uTd8X6hOVEK3qJ0jGaimDERpLd85la95pCdidqNQAOXz9ds8jn31AWIljF8zX3
LIGN/KuB6yd2zvgPNqYFU8e5KBtKdOk26O1IZMGjcG2alXa5B8HPErEOobXu6xfS2br+RmQi6mCJ
mICqIqM4KWesLAIgokIns3OEfoc1k3IkVFC++P8SI4bKkVZo5Ts72lWM7gLeKs6NnKtNtseu8jXU
9I2N+uqLs1KmQPjnaqui+sxIEtQLE3N5kRu3WchOSm8znaumIsP/U3Qu5qHy2P/zvtDrkn/gn65r
jieTsfxDWdrclBCzxN/zrATFFJxWzB1g3IL6APlk2RXwcGbGkGCC7uby6wkyz3Saoc6Jz3oLjOK1
EBabO1owQzxdI0KMDz3w5KS24t3q+HkS09Iv8hQ4YxaVIsH0gd30r2hY9D3G/et9crC1VtPfDWOg
t/7xWe79lFOKEdW9H7gIqBr1yyQt8EryPNmliRswrrQWJEy6JIL0cz6dyS4mc8odgF/WuGRyG8MP
7o+93oEqi/xfEKnQ5LQVLPLK/SHwRu+sFYffHoMxXKSeCDgAyYUGaH80LSeSgtGZ83zfPxQS0r9A
XZGSqHmvVoYVl350cM7YSNfMQlEWfueDAUOTvWV+8Cw9yJyHIyEaj7HnHh549bczZjWys35r903f
J2TowyiV0s34zYzHCWMEoPPZ2P+KwE512VB6j/25WpNa0SFyfFWj5tKFe5alLvPKEE2pEXz7AgoO
uE59FZ6F47FB7jZw4UszsIfi6UFaqscoIanJFKzCiSyXT8QQ9LyfCmr596O568lRs1Kzwz2V4mx0
Mhq67X52MTmcLHXmLItZLrqH68p/95jxGIO/PHwsIhHiPXe2HSO1QgfeVA98RnYI1jAFyaOs9XJ0
myvoqeTx/tJrujsnCw9mFP/ZVN4IJPjGdHCpCnfTu9v2u1SWVXzkjNyjhPZBNOwUrb4/tN9SaTnR
rCUIepAdCnLa05cNN+gLiSo0ZId35VGtKpm7EL2K/4LCOO1mpUX4fy8JB2jw299K2+vedNtmoewl
yfsq+rlfYyKgGxUw3ASdZknON6au0ZLge0mm0gror+CUevXFeuiuxiUNpNgD/Zj4wD192i+In5mG
FDNXV+4nYXLyPQb7EoHjBrL+v4AYsbwhGX6B0t6V1LHtI44mFMdpohu6Z7g1vliDb19lewBSmp2o
S2QXXGtmWj2QMjeRZXSA8kJlloi+mg/CeQkanCYk4ejwYJ2izbvmrkqXFKu+FvK4xn5njTS0u2kt
jzF+CUMQ21RBqwceFtTV08bJFdvxhKRtVpbqueM2LAmhGzBOJ1MFWPkyOjvfNPOQXwNeR0fpddpP
Sy2HF9hfZwTNWh9/ndXGP7C0hHzWZeNlRDB377VnIoo3R5ZMO/+fnzPy/N8l2d41BVVAfEmE0pcx
/VCe6mzHyk6+ROgOSY3ppVtG/9XN2S5OLMzdiUASoziWhtVN+06utNXvkzSXw13ctxg3iF6SvRGT
ZtuggDsQQMUFQr6TMrwWrivG7KhwnJtCBT+ohKWg4e/vuSEBIrHSuYPwDa0ckCxbSC1IWfE8cpnm
uaSm8bvRSU7wNRkQxcnxRR6pRb/d0L1nplomlexCrpqWfoyjH8gFU3Bx8Bq/9jFkfD1LHg6idPxg
Ry83kmocLtGbrY139/6LCCnSr8vPd3aDyMHxgrI3EYJxFN7Rj5BtMPkZiee01gQYmBnJxJ+wKriY
7kA7ikfAYOi49Ngjyt9k6iK7gybWsuLxyxrBgd26F7PoSjnb7qkGa0wHDTFA9fOI9AkMbDa6E3B2
PEKwYqHnVTzGgW5icjWFeH/Eqi2HQbo0WJtliK9pe1wJjUBHGBlqsKNAeLQeaNy8B8DAIYj/Ozjm
3qU95JToh7lOOWVsEu+JsdD3icyrXC4uhlEdFiaknrzm1rSAxxOvfJjUDXrn/TcUjPMc7uQfW/kS
eoTIQJLSR2HO1dQpqEPDts6IT1wZ5dwG4wFf0uuFZwkLgvvaR4oAX7R6jCKeaBezO8mNp8JDgq8y
PB4Mh7tARXYg4LsYNCpq513MN8pPLfxuS8En/biHv2yFFPArWgI6l3HTKS7MdpcwtX9PBXMImWZx
cCGoB46B5RPI+Qyw4YKZnTGDarP3Mdf8vvAsa/gU98+IS8MrkF8b+cjNFvQqBnajb4IHmiDpNSSd
7JeSTwRgx9322jfO7WgjEFIds1ZWaYM18hgfVAoj2zVOy+TgyRieoKm/v9zhRtamoMIQKxsXvpMB
4CQO82UnxsG6pylP7gSVqadjt4iOyruRC9tWvvmEIGHLtfz3ZoLKLTCLC2puJjb7Mj+juSvfuifR
QKdS37vp28IP+LE/D4oGbGbbLuDPL3elZwes9jjh6aniT9wACFRrd775TbxbVNMSBwKZ0plGelAT
n+xPnFVkOEbHd+R5S/nxvHC/stYjoxgvmgzcdVBIwJ2eSN8ssQUdB41JmiPjibogpQkpgGT08d1t
e+CMwiXJVd5Q6YXqp9cAYIMdnQI6vu0V0KX3NN/+JJ0JoEz3fbFpBvmQWA4BrfeIbd3oZxXp+myZ
STUzLJMG+/clNSQIdDGkwyNKfZ+j6O8vOBYhnQh81kUskvzmGxEFIb95P+jxTQAM06ME8IkifDzY
kValg0JqzgzmrIC+3imW2rOkWfBV8EURtcmJdc1EqkpgP5rxmX6ssxPFPIaLbziD4qMW7u5H2MZZ
oVZEAw6R0k6Y9lJoMbYzzeFtlFAU1YwVYThUYu8fabuAY84Uk0qgPbk2iGLphPmYXNfGBRsPzoFw
uFYXkLbf/pALfwd1N7e5TGPqePAxAlln8KMdK68DfIiEJhg/pR7u2BBfSzRgMHEgWNN9eeLtA5hs
Z91Z1z2iFx/iY4b8PalJ3ER4H7KgwRPaQUDAnf1PboneoCNnzHvxPYGoP+0lWrD4hL4OjIz9Igd2
0aBx8ixhO7sACJOrKZhfGgWQwQmfh8t1epYgGxZadQtAE00MMHMCcKDhe/qaEjJ6KtKM99l7Sa2+
IZN8B2Z4+UVs9WQKRwHVo/z+ywP2HPr7Vyz8CtoMyqXrMQaIu4WpftwVzt7W87qv8xL56C1W/reo
5/vEv8Q4zT/vKcEtgpla3G3ZVEV2qOAF5hlFlBjm3amzeP+2jbqEb6Ud6W/hGOrQkwJ4uBBIkYPf
DaPRgRUbOKJ8o+YtoePJcIkqAS45PTGyn7Fn5UztEFnlECioDTtdBRYAyVOMgs9iihxz++T8AUNu
ZA/tVi1lsv/980hnuL1SRHx1a5u4DpMLbjWLQUUw43YNbkXqBShhU6bvPGbJegwh/Ifdt9DC0lTi
x/GrK2oc+IIsRmrVtBPkCz51CxpWftY/c49C+RaV9zbWvAC2aONrLazNHxpEMx2SLptVbFwxE9xs
cNNxAcukN/2+YrkB3lInzxGS3ErSSdG4H0FMiNoraSUFbxaf3LPpddd0MtU9XjnP7Z+WKoE3RVWo
StOq7dLSqccGgk5lmbjU7lGnmPBAxQD+Kk4SsGSAEhwkrADAv4FRE/pkf4ahN1sVHJtYhaI2rjJp
HRavPvK45WSaDI27oz7Se3sdEMyQqHkX0hKkFcQZKfLU6VuC8CeV6QZJc1ZTtLKoVn5qg72v+Z6l
gIxDsXgnoVXcX5s0R9d9SE/OQT6jtsUVk+uJvpkhKcin9PzVNz9MXWBAdGE7BzMHAu2POAyQc2Bu
W2j4I2eGNv5L34Um1h2brbv4CCmgY9pt1JjOIy/1KtlqZC/IutXhazx2bYysIP0TQdiAqGle1C2y
L1ZzXfmV3Vu7FJk/Fx8/cPWAhU6ozHjhAztbr0lLID6euoQAY25GH5GOXEf6SMfueZgL4hKm7bnQ
2Y9QeCj2a78nBvKS/UW+AFX9Fi8MekF1DXQEv/umZMpHCbIy2XWp4XxvCxzZEAVT/ZRWizG+mSlf
KnYbKq4+X2pmMd2ZJzmQdDYbc8LXatKFnGckJtIpjhNeTzJt9YoWnmi5wDe+tVg6+A/IYDozr2cN
CXt8IJk8nhVDteN5MTlLVsZd8wp0WIq5dpvbg3EXc+WyEodLoUBDhiO75LiDQ/0FUSviclhcRGyG
vJ/YCKMZ3l1vuxLx3GikHEPAglB+6UcOBpz6DaFXoisYzDTVrau6u7lvY7I+oLkMAILlkIK512Ku
dNXDGcm5kz0adud5d/KY2oxLdh8J8JGYqVgho+5WApiqmLU/B+ynWhg0hrKt5LJU0mM25BLgvOps
SK7s0km6fGnG+k6fEtyq5ytxIeC74WM2nn3Kcu3Tt59tRvUW/xVqk/ZlwuxBCoyfUsnt/5PseAiV
akCDAgVf0GywYeJzaUQCHRa8lvX1TbD6sjX+P2wlWieb+cmJwDfyHMi4cnfXHZ8d6W9oxiCUC1AV
6m8bYsOWwoaBCTfkOor81P0oiJF2U9QCs0P/B0oFNoVQumZW0ojXnRFn7AaA+FnPy+yN+3t15I79
Bb7Go3F/VkwDwHUCV7mo1RtkfJ+fht0nXKrEGY9CLzBsJRTHAFlo4N213d961NDyOjrkT5YjKgoM
CPvq3ANMeLNf5NIHgepPnTtLOuxVVAdO8vsC0uBjSJtFwyRTHY4NVWbi2KUJEkTs4x4n24c7W//V
PzW4KChX6Cb2S7Fl4bNgB80iNerbHYFZGOzYYaHsoP4DWKYTyHZxX7nxFNnjOCU017UO4mVfx/7v
EmcXRp2/bLkd9Ty7PMFvGCEv8xlKXfbYW0Hs4gRun9IPavutUMC5qWFdwpBF1L17ur3lpmfmYkNT
195e3/JFPScyCmjj0qbs7ZyL8bnurw4C/6ooLezHKX86qsVqHxZj/yQHVPYClHvP9E6Gpisvbqyy
0tFCLDH0O94seSJPG8MaSlDm0FNe/s1cVwOnsKg8fkORJ9P8Lu9/yqHftVVH5PymnTm9tGLoCxoH
UlvG1+jxRKzd5KtNdKfkRgyO8C4fKg5malZ0g0f20vyu44Ijui8wh/5+6Fy38OyORkJW6V6NdiA/
HS3XEYic7AHqasbYQaXbq/hoiZWjFpU7gRMfzEwH3LKEnfkbyxTYIZq8ErD/cbBfPH3MhmgB5Y+K
RwrqEFL4bl++RHMFlT9GY1PDR9iMCkGp8HFmv70tuqOCvdDfXECZcr1D20+rTfoMv7J0t2zPVZCa
uukE8iJBe+Kz5wSMTQqGTQxDqeHHLSWC1dT1HjWew6aHbPusO+415SGaFulbEK3zVGc12QPe9xhj
KL6Oio061T6uZPhZCx6idgHF7cOtDBhrzjb0ts5j5hQvJxKYZq4vCctJMixtMz+DNjEcMCHOEm+B
qROpMpta1KMCc5qxZRVkql4A7KFUIj9RnS0p+YMsKClkQ/a3QxEpwFqw16ztunTaHy6GnS4vn45Z
WSusfqnx8LAjvhKaVuFk78oQprr/XRSP6gEyJAsbbX5rO3TuqkWdDWG1l5mm7XoULC7uRxq/hu2h
edabgo42RgeDKlb39xMM8dWnQ6if4/NzYGeXvmOtiYzYs8NKl7UpMJp+X7CpC/plChO/a2/CIakf
G4DifWm0OTowIob7FJwsxzu45aZAjqSWWJUdHcxtBDiPzxBzzopmUdx4zFyUBKsIzt6zKTjaNp/2
wEYfNrg6aAMvZMF1q2NjRXb0iAGN13eY7Xe1LfXFgQ6S1RBlJLSxniVkMsxX0bnbaVBQWBi2AQl6
xwk/Ci1QSk4TapmQd2ajquyqM5jnJrz5RiwBnrDMSY5Fgx1uz5POYizwilujgPKAb5oy3Kh1rLs0
5rSlA3phQgspmw0VyEaHyo+dfRyOlkZEP07Pb5EkgGwp72FXWhpWBbGlSUvfYExGRoFpVmR5flBI
CC/o7J2+equa6iZC3i0eKSHYqsJ0gMV7xBNamtjvQ5Wq5PrfUfnaK3dR045mxiDYMd06ARbS9+lx
UlhuB7DD8lqfm4rX/uzQCf3XFozKZsq0o7NvFBN90Igkd92HdXYn9JRmtIRwYjdGkxc7TLEZd4bW
xo4Rha66oQBPLhF64jsQcjkzZ6codhVDO1y/2+ZNpAhgKCdJXcZ0AJXhWDwn8hS1+037zHrpaTY9
6uyXN/w+leXj6hrYX1VOYz+pLNm38QAb1wss2Wv1/0RCQtE0vKLy0ChIExZZheRLWbciFhtOpzEB
7LsnWvzaxlmPd/KYgqxtUMBIGuC3MxTSrvV2xjbIpE9kwSGIcAHezCr487CuUJS7UZbWUBbaHhJW
ond2WLNnY+0R67UWC8ZKOrc33yMGESbYpzV03eYenDpgx84HCS2uBT0qPS8DRG30dfiDxaBW0Xfc
wUaRf9zoEeLTc2kJXAHwNaeJMJf3xgSk0uAmWRd+0G9LjGN5A4eIOZimysLH8jVdC5b/kouW4Wqz
Ps1j6RpNk7itcujzB2xSLsU8wYose6ekU6l+bgrN7n4Eh2V+VcjCFLldh7gp77WSf/UAShaLRq6c
bhvqz5s8Y5fRalTVWHpxnRkarbP4Dnq52ylew+7SCM7BCbpCkLg5hRVih/Q0gtRO4vtbDE2dYPCW
qUqOwK5v9yiycsObLM2NoWDlRWY/GBKEIDU5IWF+tDqYNmi9k8GwvuXObq0zuTCK7r9IPWpE2vRb
dd6BlGJGaSmUb0MQKkRgIyXaotswhh9fjKl6A++rdbKmL0PLPpQEeBxdpfLq0Gg/pVdFJza5RSec
kh5uXrRhsaje1QoOdR/aBiLfb7rfCMyZZgOaRqrIZ+8+9hyVpRxUGxsgJJcRIpFb4DYW3kCEJb1+
56KeTda/zdyIkCchzp3XzJ+kID1UYVbdOBpluHRl9e1U2ccQgA7w5W+NUMLZ3AJc1BXwbYQlgrb4
3rZ5+P1z2h7tWTbbPvRpsKxE+DVBG/U9mZiV9tFOVKlgEXf0idzrX7tSvfmzRqqyvYXibel2OzdM
aRdmj9w+jsIWxQU2q1nO0BgRTxUIHTavl5KwYfqXSw1zU3PRajSZyvgsoirhGEplH+N02W92+cyZ
XlLZ+JlcB9m9ec+tEHXlSKGSx82IKvrdw2+fNpf3rFCW8+Oa+Xlx2yqw/O1iVmVX25fG2NGioCk4
d5V8CAx5z3AszTMAS+MXuo4qkhVUpuahk7n7kM3w8hSzLmgYzRP/HNXkq6Yv+Vp/g59VzxoyTqMN
WrECuGQT6LtyuL9mk77wAkqWaGz2tLABBqGwk//PoWCi+0zHAsDVk4J5y2rxieZfVlvfJOZTwYRT
1k1Osz+C4cwOt4pAtEGQxwfiRNiWBVyedzLPrRRH1fpDzCxEyeyJTnhCZOuqPznt5+MJC01JiI0g
uQ8wv2tN4yKpcVhwEwZYPQFcWNgwkV1usxWIxl9cIROz4iXYxaWFo4kp1nc5FffPQkpjOyt77ItG
NQ326ImhfeG+0xg5Oj3TqM1L32bsEjIO1NVgylKmmp9LolpvugMXsKgnMvVva+UW27UPP2h+mvYt
tX26i9K9occlbP+wQ+J9gJQZVzN+19NY4gGHoDR3/6v3CaWsHP1++M/VgWz5Roau6HnJuIRu2xoo
TFEeLrxtANfQafb4oYsF+SF8TXeI/BfRatilb2ztTmNHvSU1gfaEmbJlZGqcED5W6ObE7FjajXeD
/444uvJcpMWtWfxcgpG/dwp1ymlb7SQBmlKe9ousHXe/kM8aHJIo6y7EeBswbpSa5bdJwsI/xRrJ
Smj1DLwDQwHqXyLIz41RcmOa0SJMUFdQBHMCHswiJJIy2WVsJz/PWHES/dYA+1gic/khBv20V+CN
hJQ9c3Dj2EQTHz/3PlCSzHP+VnRqKj8cMhPW5KQLCtRf5dwl3S/WHRES5QCssnfN0+6t+y7S4nhm
RJeYZSJAUOjFusPRLjYsmZFRSUGa3ocNhY3VqrMAZQQL9Q9PWY9H1fID1U/gimRz9PvvZph84cwQ
qOeElAZxRVhNuRb0rwPgiPjXqwpOUToI6sNop5ANydVkcfzjqOj1LUaZrZ2JYy91U838JB1HmABv
djrtiN/94OgqUChi563XI9tpxIY3b98xgJk1Jzp6vkiYeD6sMalOqAKNwsKP7UPbUIotyVK39DPh
nhxWHeOUEqeDxtyQkOPzbI9hNrG/EQRWmZtU7Toziwt5YuEAXAd/w9fVhzswC3TBlb2KdLlrNaQk
3BMCEHHUccjwL4apy2Dg0fNroFEPnx0V/w1YPLK5Tp7acLOv4JsESa66rEmBc6mCvuzV6E70LDhH
cUFxd3tnRy9WcTdIUal/+b3GuCTt+v8KCKgMdzHcyzJMO3wWaCiZuZNPeE2Bes3fH8xHQteVpUio
3UkNqlkqsHQP5MvrBu1zPhmjyOj8jLslak0uInKfsPBaAEiVI4MgTQtLgifwUimx0Q7j8Wdg+rgT
E9DSCZdsN/9FM18JGXj6OUaLmhZCbUbOctoMvbPGnbyisvPrgdC0FIkgsWsmdhJQSeod4u4aj9sw
hd4oZNXlsA5NrQ4o7YcM+TTAlqpK6nt+hF+xODw7GrlH0FaTtRJh1JVgwTPJHrnMPKtoZF7GSYPy
5EjQE6IdAhXONBBq46uIkwuX0+AN5wsRUMPZ1Yr68jquSZqcMb29ZxSzdBKnJ3mqqs9JOKxDIcjV
dqFemXtQs/S0sCPAmdZ7AviqjUFa4gayrdJWL3E1clKUL5ph/SG4BXxXWJq0wRzJfRApigvbSXuF
HA1cYFFlGQuaMn50/4Vyf0AVxXr09ejOjWUm45+pYRs1R+14VOINhNfT7k3fyh/tuolMJVuoteY5
8lzbYCjB/3qTAR69ClQ1jbg16FlInlSF0Xbodd56Kg+vgbioySM8sQPL/3/J6OuMctY+Mu2/rNmy
nSzM5QB/McyfrHS3zS6MqBCqlWKgZHQdFkw/vLiVVYMvl2SIkTXGsIc0c66fgTqOGxjFleuUTHLk
IRdv4u7edsiAa4i+MS3xIQPXFescotsXqwv6R+XsbcsIisAV9wMD36xBjn44D7M46DVjVvv+QKJz
HLjKJpL49VLnb4aK3kWduQWEWGsr1Vl7mNQjHrRWIou3XkbEVUDHlfvZNJcYZtIEE8g+tF8J0qoc
TFdYDQyz3hCG55Yl5LHZZdtiE3AEDGaZWZus0UpNLzuBrwBWDLNR9R47kDtCPAjlFf6Uk+QuFzMQ
ZI+rLBWflDov+VGp1oyB6OXg8VV+xkA3VoNxqg1bG5lxnH3qiNTaL+o0fajGM1ownnloK4HESc/V
VfYkwTy/Ux37suRSOxIcY77OunKtPaSW6TIIFP3XDYBq72mr1UzifVcQTlw2+VaTw+iqigMsULim
3r9Swug5f3sgkwQKhekPRZDet2iNivJvc0awmQXdYKrARhlQYc8HnnqpcBUkvWjeUd0TUdqcutsi
WzdsczhfHl9q+3HJJCv83gd0AqOUe1uF0IG4zjY9nepTtql58f0MW2GpR9p85pCZ6jCLiYgQN8ac
sMfvi+ZCYv9TBaZWlrw50M6eq5c2rzYMvONyotyuFG07+hj3FLQBzS6PLmOSVYe8G/3eIxhaZUZn
R7PPxKst5+LB329ZHd4JtcFzi0/S0LjzMDAEoHqdJQ+ht6VntMaep+TNbGbbRZaAl39uuBUUa1sY
6d2Xf1SDTmzrUHXvsUoq2x2ItIwuMAvIE5/yBfnXBdijAkgRdBphsx7Ry/ydv5eATtaVsFeU40g8
33hZlcoonJhNHuSbXy4kedQyQ/3p5mwCx3U6Cz/oZdBuXjodvtBb36M7PDLRAB+iQgUH8QGAsQJe
DLp1iJMf5th3IQCkww07CpkM0qPnvUWpExQYN9ggh7T5W/wfIovIlRoeERjGPOvNXSF+4G4Xl6q6
7h8KOGmD/WUCfHRvLbHVF3K9zMiSmUSK14G+/zCmfixOWfs1GVuF1OTp9MV/fnZXPEqpaKYGM5BZ
ld75pqr9bxhETA8VTIdA+K1zEioTyRJLhDOiI6AOTORqSPX/SUptWxWbsIkNhsZMpLnScTQzzFZV
tdQVodJiqfQMmTtl+sZLidJkckrf4jRzXxs6ZNacp2ykhBMM3Cht/RM7FKn31c5qZaphYxv7CDBt
yHWONl2DPJXTYkz4jNsgNnt1LvpPw8t1s3U0KFBE3IwYtjR13bZveLd6us8djDeOodFN9DP9HifD
kIRGZWWgRaaiCesF/b7fdnOjQV+SZOW5LZSvB8Gl2yVN8kdkW9mkLl9XIrydclMyg7mYYp8CFeQy
XA30OqcD7jbvUJahre97L0DwXGFvX76JJ64BsJOrswGJZ137bVF72NiUVdfua7lu0ECTdzs/Pz1d
qZNlNjEAPLF7SFpNw8dEF6Je/F8k1S7YGmg/FDtODOJ8ycbH4MWozKPZjRkSw+IP0pvbYNcHKAjf
eKxOW3J2PUYSL2rRroDT71mQHAV2xx/uZnlerqATTcI70lcBGgr3uqBstYGqyTgAJhWU/sbH7Hy7
OU2rXEK0z/ZmPI/6wqRz2zbq7tr7AUEbijFzwWHuvuGvrtT9PRyxYslVtSeZWXXFWOKTUZDEFMeK
HRssYEjOLXOskMAKdF1BmpUOpPBtJDrSqtO5HVzpAm0wPBSRdSbL6gY2FqNrfuS7JNkrEifSVs9A
FppKiRc1Pt2nkRXiJNWf6r0NqpzOYM/WpRxX2z72UyNbGl6obZALpUQVnmq12l+tQghRpR2USdv0
oDkKKcYH4B7AMGajm1QocYqstzQAX7/iEk/9mPXJAIWPFUQ53jiCoW4cfmZ2I8mOAu/MSya2R6oX
55/5iBWoxPRVyWScQUUeXS6Pr3q7Xll8FXSWik3cXnLdnQrCU6g+35XnAPcKTZ4XPK1N+gjPCOK5
r3/ualll4oSsWylDRedVpAGtcCzndjIacSTAic2YYUC0lqd1t64YTB9fIDMyGZ04hW/+GUsTWf07
nwCht38PAXZy/Ycn1NcjFgY8+TUvB6L0DGlLoYP+RxYR+J/wz6ROxKyUgY5CjAVhoT9hy2K9ORf8
WuNnLUXR09dvJz3B+l+9cGxV+8Y63/3eShkPMOK25D2ZVpoiUyAJm5mlu4TiYPiIjRDb2s2JQbXA
CxYT20VA7Kq2mFs1S/A0wP2IAMLzmIdKhRo3FzNL9YRzXkbIVvddQk71RRgRjsDeu2h+UFkRgoGJ
amLg9dIT2DCiRDIG/Uai1ezvRDNb8o8kUFbMDWWUSzxjFI96jKAItP3LAFrQJn4IOs8FJWFnn1cE
bWSpwKbP0/NONSwplR1/2OVldQjAkSe3Z5hT485E6viEeqQNmLpoG4/y1gp+aIAwF5GGJvSe+VST
t3PHdnjwh+Ql15sdo99UPTsLgJUQWX6sVTHzZWXCM033RWynjDpSLIgGmmIxqROmk+SIc5jle0y1
MgozxXpApic+H/R0hGQmA/NhmFnQYobjg/y2GzT24Q3tqIfSJ4CMAtZok3rmxYn942NWIlsKZ7YL
wy64wXZpYPhu+aYx4vKQMZBUK1MegQBziiEtilC+C+Pw7761Z/C/yS+gcTNhmfkYunW2HjfInlM4
WZPTbRAghlHqxqYZ3H1cb02n6e/k4FZwI9hRFEiw8aPqWutCf0isYD6meyEYmJIZoth7LcdFdG/o
OD0tFek8MYf+PnMR36gpgmiFHdhiAHVpyppM1MZN9nIZp/xTJ9ZdXKVoHhDi/H/SBmVaa078RIl2
REfG03pqOoNfRCT9AQ20HnPMLlp3mHUNsw015SAosFppDYhT/BnDF9nUXN8I4vq96z23tcsP6gUf
6QTcRmHaaRAPq2iMEpYtRjmPkrnugydRBTZDW3USqM0x3KNLvwSGfIp9nq7K8yqYPk70DOErTWDS
X0bdbipyZvKVTTmCSlgqRmnKRlWiJPmlJADHj8Fjlsd5oNEttWWq/r67LYCsfMyOb+BK1pV3xiu/
Gceod2M4vOyh87BmJgX5RsFtAyrzD2oMaq4lxDUdA1a406ScA0tH+bqpwN0SO/CjCOb2ONRNlmHf
pJGFNJiKFeu56HkoD76mwLDUYrybKxHhh7qgkchHc+mwrxO7G/ylS2bkqqPmzKS/OIzp2OTHhTaC
AKyibdZAuocCYtX+AIM+u6K7gJGQ87RpHEYUEce6sHFAG2xgQ7m4NuHghgUm5DcusjIbx1gk+fNE
cUyf6z+GoHDei/QxFI9IrBJMcmJxAxUAi//fsDMOIZBn2X00nMmE03SIm5JsIZAX6xdMzSMRwPHz
Ydj2+KD6yXTp7w+OwH+gcc1bLEwt+WJBhHqfS7q+dR1dEGHcL4Td9wxxobi+07I/GGvZT5LDRKAS
O/jc5ilS+hlP2Z0K00x5h02UzE8wlUgLZ8iMCgPzHTEoLNRQWuu/h32B5LRNxeDkF1s/hdHhmabI
V03/L0G2CLU5jrqHnKdRxHlL6v6hQe1muE5s01winCLWm5QoFUMbd/54Pli5QHCce23rLsVyIXOM
NWTxJQH8ahu0db3u23asSG94BAlUXGvcatV3MR6BFlP7NrJS/NRdsAh8lPLFUuYJYMFflTdRcQGX
RrGvRrG16lGsHRGGDSU2T9pO1N7no93xqjXejmbelS8uXCAerURhnynHmerw0cv+Cf2HaA9XzgJS
1vqPDzt0PHNCygtHoyKdO1ydQOYVQmihPJFzlm2Bc+B+wZ0plLX2CWAEVnmb2r+CYUdhD6fuYmVx
1GCX+kzfMqGdg+INY82nqaNn76wmA7qzhkpfncM+4c6QVJJ4/gQUHF2jue23quFBGuB1FMkFFNf4
cjRON53uHU48n3ra+FQ9etUf+iwhHAtohCwgXKX6xT0Zn6mA+jrCWEFZbQ+1FDCCAc1Qfv1z/VCX
24RWvPeoAD8d9o8diuTo5QKzpDnePUmkl6VTKIurtsEOemZ74ZpOn2QbTyMfjUO1RDj99EgJ2O7f
isUEPwEyRX3+EWG7tMXMu4y5FXtyNktnSNWhD2HR19LeXezIcBg2l3fHZUeZapfTcT1QUotL3Jbr
QjPcOWlxw0Ru4bu4ektj1AlX5zmSGRGbCt5Mb2J+W6XJbTRKb+AGSY4ZR8NMOXYbggCmvs+t4CvT
OH9OXxx7yQTPOIF2dTv1g5vAiJldXmno0MDJppiKgM1YtZPPzWqbL5nCtmKEwKtLeB7ePX3y6dnp
F7xMEu6IXxZGM4ZR8gPDUbF+8zytQP2SFSFDxp/08ZFBeLjtgX0cA0JBjn9Vw9wJ4EnXj0NfdVCc
sAlKNaDv8bxvrZhUUbPc0zqvd9/tQxCEoMQElpqWtefSbsMN9Ax0HCzdcLwOUAJpVtyrLTmKSQmz
92Wfnf5s/lCgbakPMqyjoyRDScd1qi9SoDIOZczDQlw9NBhRf8ibijqD2SeeqS2N2H5UFK2fPyLz
CEgq8iC6MLq/vXLgJr0yMGOhcDnXU1D1oeEl+J10n1pokfrWVrGetFEJ3u/s9Y4b9dAzsYJ81rz/
maHTM7wtxMGNvEuKo/XxhRQljHIzPhLSxA3zBliS4FxwJmrC4aQADdXGDpHb5o1nyJ7LzRnBUAmB
tpiFkh8eNOac0xrxQHrtdBfpthRgryv1bWiNXCt2cLi3O8bMaWX+Vyx1XaGgsyRi9v/qQyJ4H4vC
ByoCT4WVvS7/Vff38TlcPigyV41yI3cR0iVvBR1ILOvaHncFuqNnPd7VQqe5VVyCLhB2fDRV8aka
K1Uj4ybiv1v4BaHfEd8fdoMiW5aF1tCp1quXlUmCtdEYr9BB3aT5Bz9/kR5q1mRH+tWC4/Hi5w2A
IY+ghQQEqc8pp4Ip6E68MahjL+t0E58yQNDudTOnzZYF/OGGYGRRP73Cqagq45ohAFtCDvWeZ9HG
o+vqUd1wDxAr4NOGKlZL2w3UrokLRH1jMv96hzuXZ38Zn5klTaZvE6yrbwVZ+DgTF8bJf41ieuca
kZRi+sBCencmlliPTnqvcCPvp+yLVMx/PS2cYYhlb5nK26QqHr8rz0DCTrNbZ+DthelGC8WSWQTO
+osWCB6VlZPNu7zWjbOYjw1SAuXrg7/NyPD9mUwWZINUCCAqicg3DbzukRmhw130aLflI4wqCLhH
O/Og2t+XCrOF145fryQfoqDhHLfOBEWDf7mZAWfky9FRGF0g5e4ngu5PF98+t9z3BArqzfaO/hVm
KVNv0RHMxiHfuY35XF3/C61XhzlotTdRaPKyeplxldd3EtSht0+6xy0/kRi9BpIexQQqlusSpNAM
8kIAbOgvXOIFtHSutt3CvHlqcpnBtD2+i5quONVR7QFnxwj1uhLjxWKWS3qTQq07RgMt4khNvmMm
Bjt6RKHZbJ41iUb1/9/+jzVPETJ0W4ys7trV/gc/xmOdV7qzh4zu+3NJBi40Aymk97fqTU2nX9E7
oF8nxjIXDFtHrj4cu2OE+7+E+dcG03zkEjc+5y3MnVbOei5uWByKlLHeE6PklLTdu34ZvXWd7C3B
DgD9dnpODGxHmBTBkBF8GjVPWA3Or6X7HpDbsrNWEJWnijcl3Ks4fkpraWk3A7b/QTu3sL+yirUl
UiRR7QZSeiU4XhfcYx8Ib1wmoiG8LuTBTKYaw7El255e1rNtZO8KSXL7lzn7DIe1pjBfBarjcxTb
aN6B23LDc4BoU82KJIiAONFz8oxrvB+OH/7zB+KSGmW9UmxGOFEhVTKEqPMM4nYAbbaKmFmgyDF/
uQB6yoX6n8J1JlUxDdXVRXC17ZbYOZojcg8PrTYvWoFphuiPDAN9rJuiz5H3AkSaN6gtzNV1Cdeu
MyAUBaEWk3ondYzVeTQ9qVG4MnG3ThicErjtfPOL711wWNOmEjiP9li2NCRdQCMp1PF+K1iZazAB
0QA9zuaKQoA8GLOQ7nKFw8cjJQTy284FogtZH/ndqTdrqcEIxqdhZ7O5FaCo45xLq+smDoPx9ukJ
Sahn0Y9noIRCxjk16np+bqoj8qMQLBJjgaCulRY5w7jWpEtahRumtmcIyhzf2noVZinqbPzw5zfS
BBLjGzdwNBT+0mMyrLZ8iRYNt2kFA4vX6afq+Spsq1mHqbhSq9sQZpTPxz2z6BcKE65+K5im8OJ+
T1GERrXgVsIqfrwDxpCgBY2iKdO+rM7i5pjACpUAYy+KPfh8JnwRmrWtZuQrI9aR/gTU0LC5VjSi
tpTFKXSm17FWKDFgmM1eKJBZEqv7KZYeT4B5c1ZSnAtPv9wqIAQ0Ho1Am13OhbauPi5AWHhOsDhN
CfqJJbIcExjGg+YnwOja18Lw3fHJVxoaRqdpjCZCD2acAwbIAz2PyUOuFKjDo/2JPE3q0seiGUwQ
pkJybHVbZwBIfcfnIE3HssenJn7e74icFunFbu5PqZrftuu9AqNSpZOMDAs5k6YKhkJe07sXtjnH
xy8fZhkl2J9XHPYcGPkdgeNaBNAXBRnKMa7vHDvi/Og7JiBFZN30W5qvdTFXsm0nucSzxHdRdGMJ
FN/9kYeOFCF/uzqA49QuuaT1j3w8kIrJRTRHJ7td26kYCr0M8HXcCFZq6kuqfuPliewf5Ato41aj
qaUrVet6lAbsccLyKm27/acGcxCkBqvKIo5nqqjM9IvN0o23UePVgYOY1riTff9ft39i22FXOdOp
/FChPrbqWC21iWPnZk6fA/PVD1rl2ctv1yuP02fnGNT2Efvju0eANss1ez8DslhbXfsft0cbpiRF
9nlT/oZC9745PHouDsqHcuSckUPVR/ontwubyWaNC34X00cl5guXXigQk8gIUFPh6Js4J2nL2kEd
X1u57jsrNnTQDf9JGagU5WCnvthjEiwWsNw8z8Gc+LJRHBffED0R8ButHTRuqmm/I6t6Zp8rdeVa
ZDS1hQ+Mw5OD6U/101sr4Ph/5T6WZLEFEtMt1u5jlkweZdBg4su8DK7TfS+w8quNfzBYyWb7q5au
8YN29/DAlsKLYah/pbvKV/ipAqHYqrYt7cpufsm7VB+tHXJetp6lTfKuEqaLy8q0TcfL7f/8seJ4
jteBBW+mRsUx2/Jplkin5xqSP2oIbqDafwCJCmlUqRlAV74b9CTRyfTIDrRoK1H50qPhXcGFbXox
7P+DZsgmrjR5KeihVDEXQ7Jv7Dregkq0KrcA0EPCErhT/CQbLC+AVIEJDv4jMkkoLzWh4nnjreTU
6v4UqfneD2k12N9DNbOQ12EHGdNaNbcK+Gi9giY9sOv5OZlz+S8y23JmORCR0G9ZWhbtSPxfm2wP
0Ncl9Zob7xdKdJWmkDPlX+Xz/17JObxHx8x7DsgKB8GVZcjEhDzjUPTKVs9KRf7U9SLcc1FaEQiK
gl0TkDoWDlwlpCE6dzhPlZGLwzuCpp7MeuiWWz8fRy4LCoaASh+83TzYWqzShSolc/Cnvo5KXuw6
Apz/2sz6M2ym41d9dwPbg/LMQqqp+gTGh3MEBtAf3t+Mgl4E7TFqOBu4g3YIPj6lKkXdejOGL01O
6zOF+waOetsIsNyYRrsQ5z1SK7OdJtMDmgQA++/fYi9uCwxGCN2cb7FTu8f8lOkzzx02Y7XDRvlm
Iz65S8vME+EMqzwff4CrhlIZeOgSAqATvE9EPGn8hSn5ovNmiRBEel4EpMHL6BWzoLlJXZnZTjA7
ph2wXDAi2IPMpP4sWjVbwCgKJd7W0kwFdcI+0loVn/Pf75aYe2qAS52Suv1k45R1h5b6okd0gg1A
aEQSW07qZtwgZBPTxI05adbMBKr6WVu5asU+dEfK5bz+JE74uZTAB+8zuminOIQ0vB3A7Phzm9ZS
9Prwet8n1fKpkxg2a/oC4QqePMV6bEjoH661vJdNTTk+iga4gUIindrOEkoayomOdAm4JTeQx8cE
8NWnGryzabnt4oGDtugVWNzfhpXg9Jad3uV2osMdxAFAVNQbwy+7zXt4Yv/VQPkfVza5YzH3xAFM
uwmQ3fKiGahbEXc3NJzSc/vUy6mnQrRjwKhGqG2UtGRCoCu/Bs3YEn40440Bmhl5wXEtljDy2ccG
wNS8RbeFFB9APDydXIR+uGXQ7A41JO3Wc9Kn6y9aMw8SU9J5BRV5R4EWtZPavyeg1ZVcKO4BWRFM
MzkhlP1suWnWR6e1w0bMAm3C05MZvWlBGLwJ+kiN04jD7DW7yOuph3riqBbXWsxBqbNcGV67kOW7
YOanKgl6miUElMVOcZAC8zkrX6a2Iid9F3Wa/swwcezgQHJnmtrfE2DHwZn5fDqVg8dK/DhOaKyz
fYziX0f5re6CWKg2D0UgtomCKfdP/sUn5Al7pxaWE9demaVGmmfL+PgszBgN0VjI9ovZ1pyxb+mY
289+b++N/ncqzWOTwRBykDlYSnrZJzapM7uoUWYqMLTS9VHUGidS7gwLR5zKGEcT1XP+CFnP4liy
pgUab9pWO6Rb7kRLOrhbcJtr9YxWODd9QUHVw3PAwybiiGkNExESo45dyf9w8BpZ78zlfiU0Q0oO
9AIrMJJz9FCPdKTrP0fdEMt4sP35qPOHC2Dg3cb/i2a+hmkkcYwvHPw3neaKsD0pbMPJ2bA2/JVd
uzAOQz87h6C4zOx/xD5VOiUgyqMvhVCAiGfYZt4ZyWMBOsV4YsxbKtBlo1d4WCTDHlHUMDusGRFH
lQYm1RHg/lcb93pSqjXSXEIlYC+GvjlTK2K3p+q2Dx4p9p4wUfXDQQm9k0ibofC02028IikYgSuM
MJWA82a08uD1DajCR063Yzn4BtuZ1SJQPq0SuAT2lTDtMHh1vDeLH5D6bHFAWLQFwq7XIgD4JK6u
qj8fQ8G9b63ub8fDGG+h/NbY+4JiaEcUWGn0klELM1TU8KcfPjQsEfgbc6ONHr1Qzk+dyeylsXJn
dPqcY8ui37EUlLmITWASFtOtEokLxeNxKgIZhzjQ8BuMK01zc05Y0aK14I3hpD7TUG1MrUcKcFVy
UGW/UA7xHMqF6g/QlO5hP4ErIZuLXGce6CAw4nk4FotCnFn+vPZc+OftAKDaTKCDfue0BTxrUBFu
gsCFqKES9RsNOE2bv09f71CoE3C5FP2dZptma1OXcGWIJKCI3JNFjGqGGYL2mau2rXoLDxeciBLe
+0QbZQnsgFtmiAuTq9i59OQ6IrZgWre2ZpU20jypkgk+LyQBG5fTgGX8vnNLgiNuAUjOsrHWFPSB
l39czeZgWbIbnFPTf7UjpwfnfZhWCdlOOHRc/h2lSOFrT2Xga+1O+vnzvJw2qs1NNtBY9HeAMIkM
twTqtlOFog97DzODc1cSvgo3PN0rTCsNkOm2X9xP3Eof4UnCslMaC+mX2iEWv5zCwxOcTRPkQ1Ow
FRTboyk0mTfA6ej8ClMuLb6BUnJ1tc/sn5e1cieEu+6YypUrC+1iJSq8NDYqVHwEU3j4wkwo5AZS
r59kpRdTXoK/Zkn1LPM5MHFb43E+yDler4ypTltzcVZfv4RqCJDMz4hIn0r7kf0YtxWIxbcW5UMT
JYjtLxITbEK9obQkSJmk8OaP+vwxThF7g+aWbgLtvReiAVaOQQAeqcJMm6h7+8nPXDVCaDtbEoRq
XJ46BfH7iVn8uFH6oDmuC0MletjIxHCjqkyQKnKDOpNyjWlRtlSCy+Gh9iyD5DRHtjReeHrmgBe/
r6FnB3d/Cx310NAerTlLUVSXvMdfh3PJyG0NYY4Dq+seUzA2z/p60J5lBWp5QdF1Z0P+t7v8CNcy
ADbORhZJshWBC3rW4mqSx67brToyToNi3LegfW/HRYXWa4oJafW2Jeo18vnS13WIkh8UxLZPIcKU
SUi3Ta9jiFTvZTyHdROBwlZAUNqeV73sPPVmrc215y9X30OXUa6AkvrdZK0pPQ53IcXizlvlcEAC
Al+/ynGCshrIrp95Ii4yypL0/Hlxys5EJLbOQOyefGlkLGe2OsXvn7aCjM0UNvWZ/vVLY4XeTsQC
+GKKjZYRKTrHVeg3HMPrOf+ym6PmDbmyr7cKm/WP2i3Dj+uTq2/KkoRDoUh7NsTK1YNu6h2VgKrQ
uRTHasx5s/xnUrpdErjXTQJpAGMD2hsqOQj+msSFgvYF1Ry1/KjYyTidmFOq4OJbceaULufvOo9b
81plKDxhCM7X9GbQHLUplI7+UZ6JFWKVNUKTzVELm350Kx9weAL2Yi2UhtAU2pHLzF9OYXoOAhSn
eynVKHtqCN71/ubW2Ao71sNJlGXtPf50iTaeJwLqB1lf6+mDZWU8bmK81Mup98M0jPg8YjfcWGPk
cepftI+0JVy0zh5fCyxuXe1BFctgsuc6gfIHFjuKXnZ/vWz/owFCUSxS096qAMSGZ3qe38fgeUW4
lGKPVaC5ePcCMjUwVujn0Hf//goXmxq4ItANe8EDz3T5fJ43z7DRzMetdkihmhWLw+xMYZuJnOd6
wDAFR7SDd072kgRT36TQT1Q09y6sM5z0IDyMor35pASXYNGKlpc9pR/9rYylUpE824Jph7pazYxZ
Y+w0IR3Ix0KPsIdQ2gWhszha4xSZGohy9vXvUC6TvWDvNselsTppT9e4bDwOAA9T0wACKtx80gZq
fjZYWxEhT4Z3uxTK7xaxzaKntzzdED8EH9oUH0ZV9nMtYx8Et+gzR5vcF+zwANfVIlZjsTqr0Q0m
M5snI/Avh99YH2VzwykBofuB1zJd/wjfi3G/3QQ1kI5bt5V2u5m3eYpEbJUBMgyNLQpT4nM6jOT7
a1+RLs5pFB6n6i+ZvnNnE2c1Yok0TPAKn4VTbJwhTkAyLdOS+WupB1jfJNyKH36mn5L4jiWc/UUj
OZDVzCkENkKrDpuEw1Emz3L46O2Nz8pRNvdz++vpnUKWBTv0+++6g2sM/m1uGTprI5cdBFqFGBqf
bkl45YRYe1i4DwyA8TY6PHM+9tCUJKyP/l52j5eu7sweZp98n1Bkzrr8rlHhgCQhz+lnnMwOsUdP
l7n0hAL7SxlpYhjG6lqA7OT8CzHMLVz/8BFA5qtjI1HHNUk7POr+x2Ru3ZVgVONRQsNeMv8P6rYc
wysjZ9mAMRrsyXCZb0x/ldazHcHIpojGV25zdTPUIXTp4in5xFbppxFYArx0zB0MzBfaDMU5x6ue
UGUt2jb2e2VVVkvTnIU2GSGPP/6RLV9/Dg9VqO/RujbX6g+cSFNO0uI0SM72uMPOfcE99pHhcwI4
X6lsSpTzvER3S50tj9C+N3Xd5DRCxCTyGLTw8dFkWvW2YCW08cUyOHKTlMyRqRaEV4co/8dbX8z3
ZUycUwdV+YuoyMyfrI/m/JZv3Ux0VxHFRZqUsgAQrSNyY4CwKamt6rMKfJ2N39Xq3quOaJeDRQuM
GlXL8NeRGZg9hkMOAamwXEvFDNCmK6oX35/HRBOXBqXYwDadF5RsROpsl+MPzYQdDEB36dbfYXoK
eqCoYT74KA7oPr7nWUiSsu2U0mtFhlBRupJb9Hm3MjEeGv/fl7tdtLuY31VKdd1dH6EhoLsmzGxa
Rb7pd/u2f+ccc2/fzdhLPqQqEO+RottA3ApDzOhm6oi1jWCBYjvFtNpMjhtWeJ+9dIBys8SFaqFX
EoXdj1Uw5JhpQZv6zsY0YQPGNpnhU2ArwXGV3vrGIQz+wF1vdw0tgBTZud58qecvAnDtcp7J7ObQ
ZC/rtNS411YY3OGHTn3jYRX3QJvm0+J6qBhef6E0TCHJ04HanS9/nn5va61Pb4ISZPdS7IaZftyt
a+8325Pv4r9gmhTHycb6eGi0oXz6DsDl7DicVHuCZRZ45kKWFHTKdv57cuR4CycZOeawkFHeBw1N
ZnOpHsmL+kqCNIeZ9PEWCUI9YNrOSK3PwwE5H8Rb2yyPJfFa/NYVe1MlZ2hA6I3I0Tu+/ZBS5ZgN
v2uq4bc4lXY14FwpjzVFdNP3SpzFEABsUULg4oio0E3LUSXFcvv4Ezf/Tp8zM4gsfw5psTkENcjc
tu0Furx0ydcjhsG+STGeBzvlkzWKxKX+d2MOR7+JKato/lJggNuzlPuqKASx6KHrNR1J4EeeQOJ+
O7xcNwmU0+H597bFozu15+VzvVEmfLENhxZfuA4Dv4Exad9ewamUg1nE7ayGKkEqS21IJDNof8uf
spvDtYXg1wbgfRgWe9eji6FyfL1Bfi9NRPAt2+8T+/XqLBT/Ok2xSOttWrdF7yhfjb+jrdH89eQ1
AEpcVSKIiUSIPgEdsOI6vkBAmalIBul5bDSD77Jk3EjIay+8grK/Q1ppeLMJAs1lx1CR8Iz4BqIS
zGYsq+4BzGpvp79soeuyou7J3x5moeTB1V7EMtJzHSqE6IxKG8IC8ydNz5FekDPYS6c7E3Cs+YN0
Vm/ZAYE//8Om+40FJypCfCVfvMdavtEg7sZpBkfzyXt9sU75IpnWyAakSMoTU6sx8/NmS+A5NNhN
ejJKDj8DtdhNJyNs7FEHw17m+mxS62+KWpaR1/rd14IDrmcAuXYLyAyPXeO9LLgugXXN9+u37bU2
n7qPR+hVwtYnVg/CE23dlyidPgc0kAhAhz63c0gDBUg8UN4+J5C8gpQ6mAg0iOyjYqytJqvBFd7j
9ZUW3XmVlB5hpe/87YpuZhp9dNUPldSo/VYVY881FLZU4QQ+x0rwSFzA+3Yi0ou0FvAJrsnW7DsQ
p0Wa6eJEojnmKsVhu+dE+VlZLelHHI8iPWC5mHyUOpwzT3vKdZPPX1Uews5m+rVfT2XLqu7qw9xk
4VwQkDVZlD2crXh9VLT5xFShLyqb2c23m2Nfere2KTN8b383RcmABry99kkcoRf6yQr0k1CIkyEF
dULgC9g6H2hAsQZq6J5xOEf0wymdfscr30hvRufBSeQLCab8g2S4UJg2Js4pCxmwoxo4PInH/J5l
GPccYaaqhNG8wDBeID35UT1RZCc5WVJTsdeObDPqBYf5NDiftCO4oc+tTxDYeWXe0Uj/sM18u6xy
o1bQM3b8pTEif+33hjVrZIBGAO2cIiqUiv9IYtVu0SVos/6zPvhW7Y938NHfwQ+kalW0ACKtnyGi
6s8q8AJ5TalW/ik0L0XcaUybK1vvLbuSMXV/yi6iv63a7iaTxf5aFOnKbK3Jl6YXLpj/NvXl6RHi
+cSGvLo4/a5ibu7yY7QkmK9k8b/inP2Cge9q51iehOYSOCWlC4uLwNiFU0M7cF3AGgR06QRO7Rgm
Wd98e9yKZ0smusNQM3FCnXCCgzzCiaV+7Y93DrFYtO87WIxksBv7owld3F3EvAVwAKjBDoTpAYg2
JnkV0+nNcz/oBe3GdexxngR1uNs8CX+boliUGPQ4o2Z+Bg8OvE0c9LkhzC4us8JAXZPxVunhBo5n
beTPmzKYXGWh/ACmT83KiMWYK9lWSFzd8UKlp8ClF46fliDQ65K7OQc+vZ8JtcS4pVi/H9RUAf1D
yL/k9yvxmPSKL4ROAwC7A+72KFp/+ZWlx4jdkkuU5bULsv71oJQ6yls8GDUZW6e3lh1YLqCiZBQ2
ObAD7aWca1vsZNaA3ozTONLkXe684m9tpuhLJ8BZOx8pTqMGbTor2CqR7ybB5UNevFLeVHGimIY5
lqsQLIdRZWDATZq5d2OHAs12B/MiCfY4OVOIpgdS865EviX1XpLrVyEuQw2gBqXKubOEVwa21Ah+
QXSEI+pAfJ14zNHDomS0uwtiuuCxVPngYKOdteMTR+UIuvfvEawWhfbP28BZr1PpILsGRdRl1ASx
h7b8AhJNNGiW9aHdPJ3q9MXCz9oP7yOpwtmChqmicS5dycng0hPrYrq0cnLyIfyo7S6PTqylvcI5
g5JpArRNtYcXpTBV0z2ugl8mkT/3oq4sKDvMyDoUUOibtJbEhtnql9Y6zLa4QK5OvmUZz+2s1a40
EFce8wOiL1DD+wSPe5/EveG+RtCvvMnREeJIxf8bM+poSHvo3+R53bFTcldY4OpNwy8bd5x2Iy9+
Sy7DuT3HqCzSYssCDPm3P1+A9g5vy7DGp9+iBsYDXvETnMMdnkDNB2xDqEFE1GnSjqKiFxhOuz5G
KO+1Ku5uInhU0UMPAHdrv9BmiUcQl5ln/icpVHHVtSua6mJBXuIqVKFYUeOQeGLtrpsfR4ZIYGDp
Eij1QdaIhx9HXdwDmmIEsZmrGE2smphEUYlzekx2+wxjZya2+BHAJA+8mVhRHjIoJ67JxYky/0ns
PNvsIvbB7HhEW+nETZU9h1Vw7UgJHvczA4KInQSqAPT8GvSSpJ4sXKHeK3BEUASzYQ1CnGbIEd8Q
OM0FgX+/qr6mDLbcRZhtifWBQMLiXBJ3RRPDkzUfwHyGZxc4ZlraSQ5iMKlpj5wwnfSnIMRmRTUj
VEyY2zwkinVQutyzWBi/ACXuT5ccyEgnPEs0NqGpLT8iNLlY+7QulDG48iKie/Yd6Ap1zZ+ZzMHa
WKfev2mnE2G/d2U8ELydw9FxlEnd8pvUJBymUdnB1q3xCk3cMTIgN0q7Oihw4GmkcJ0eSOBQIFdX
vHcdroJL+SUvJnL2+QO9odAKLWzM0lubC2XG54jQj1Glfwu0UrBWIDMIz6ZZ3Pf4/+Bpsvxn3WlW
RYl96Ah12lnAeXpMkc2iIw/X8EGmtAEjC7X2Nvp54gWsesh/rLyhuZLX+v/UYv/OiJf87tcibCkK
SmD+U/0lGBJ3BvDgLUpgPBVFeNyS2OzjCL9tHjaR08PEXU1HKRH0oL/h9/jnse415Vojv7bo+xtq
1zz/3KK4T5YUwn3wzDupLMf7V2MZPItPng/TithPeEslj8SO/f6x6ARyEdhb+ETrMtOz31z4Jx8L
4Bfn8Cai3qWqwdrqy2b874OIFjP62NcEXC7OoZ0WzwsBvYqHKh3jAVCO8sHnDOlS/bthKtYy3ujV
9v9dJBHp4uDacBb3jErGA5ciwiFuuNT1ZWWKKUaeCGsd+jOdn3fBBUlHOlxQFTzXoa/Cw1T8vEJ6
M8tMmpqE/EP54pmEVBTne6rgmRYGcVecrOeHGKteslSpUUuCPJ8m+cZLPJG4xNhL/ARluz7fDdPh
ax5OHV4kqSIkYrr1+2BWdScMkODOKfh1+9c+7UYKeOCi67r0Y9fHJftv3N/XZHhxuuOL87L96cgo
NG+AQDo2235nk4270S5rGC4+1ZJ8J9w6ENJVwg5NlogwnZkmPHsBBiO0Wf+q/5uqm10i1qO1x/CE
EEzl+fKIir+P5OIIxEzDeSW3CbySl/rBb/oK2PaGodHLXEDeq08xRAgCG3jnYRj6yuqOxg2cnBAV
I785JqY8MduscgWGjbbb9gfNZuwhXWd0AD1xgwpn1MKr6hnUekzPI7mot4KXslc5n5gBwe4vZYr+
HcObkD5rz5VY5XWTfQ8kJWB48LWQY3QU2ZiXgB9gskYhHgGmqRKKf6Uck9m31EdVgyFMkp8W3gR+
icibg1QzrMKgBg77msaXAdA2fvNYdObPY4wMTrMi/i1MePvkRoaQuk3yaUM6xehgKheeC/J/GHHx
LlfKP7vjmTlk1oAfuoKlu4D0YqKwb84kMBJvCABHKTNDEhMBjuj7k5dw6a0sfiyL0lrh/bIp9weC
2VE8DmhfCqIe3T+B8NsU5htQt2+HE1S3yxmO7rdtMfCUNNNJ+u86NshUNxTUMbbcDdTlQUC7VvhX
+lHsnLgJ2XWoio6J6AqjY4kauy1OyjsuFC3ovQjzluldr3AwrkrQrftNiJ3AV/MTI+zJrTFf1w2r
h0s5bIzecQPwTw9RgQqek8bFWDLsEkv+zwp56V/2L3I+4El0DdV5tMo7/4u6uXl0+6Byy2rVPWt8
+SUSgSzRpfZzgzVEhrjs79l1MLHKc3DTAPpxo27k1senmTQe7ovMUPFuecJiRH59Q2gbgR+Juzji
1abuer946M8MbkgXnWR3J/PZuHzPMELWcgXFqHZJLWOm7Ae/qXiA75H3F5ilCC3pSqaFFpP2XL1y
mWMJW0MaRbBFFtXJnuUNBLE7CY1amE/q6Il/JczNw+M2VpfUZJ/A9/ryg7vtSs5TcOY0gW9gkYzf
rQo36caycm+28Ik6KG2++OcpLia2Q6WxsZgcokSbEsi9sSWX3JlaFXfWvHOyM8SNbkhrbpIvN/DW
GaLGtIyRr4Ohf8g2TJ793OJh8nVOBnK315UZ3fM9WT9b2YzuSc12HmfNrIu5zIpQpVOo2zC6OFbo
Ll/l9Ad4ZvFJEw1jvfr1KytUcbLY1hRpuQ6E+zT2aIFm0pGhPlYf2EpqP8rLIb5eUIB6R3L1LWrc
Eg34hJVtqqylmEEwHsje8CMR11QdPe5/5Hw0KiybFlFbA69vzfkvQ+DoLLaocLDz4GgsQj5JdyOZ
FV2sBsVE21Z8ObSZxPjqaWcjxqTiNKeWY/KvmPD3TYR0Is15Tbiyhyfb3AmWjsbMkhBcPf7/ZA1h
b9Wp21hwt33XyDNg9TtBkWR9ZjxXRHkWxCDBgGmeSGw9ZoJPYTvF35zFHAP1Uw0FWtrIFCCKeENn
i6ShbiAxqb1CKm58kE3HLxbhe/srU2ymQyuhKh+3RBRamxcObAgUz0ZuWDz/xYpDc9ooY529KuMZ
zyBEqe90a7e8rmsQqBDMGdie/3FamrP3CsvlgRh7CTxGsgbjqF+OiNVrxK/F4BDwxKDabNNV/e1E
sbTN6MxQkxjf84y3+veUILbFRAHDBpiRTCJnwdh6tbp8EfEmY2Cu/uptDMYV+Kci5xd6hH6vvIOa
xhKyz3wd7eVG+HxGOzqHThzW+ArhLsZBOLLAXKfCMZiJ9KXLdIICjYhGHcki6cXxQsFkLJJnWKYm
nVvhxECpnBL5TxwXUGkXlMLcl6Iy4deqF5PrjsXkCECxzy4QE81CfL8vWuK4gVZj5LpDkVa8OL2h
3d8VcaMBe2JeDj5scwCAK/rzbK7/OHcySMaDNRmgmhJfbGK7WijXq0MoOSaZ8AfU3MSfgSAgvB/N
KwvSZ6QpQWM1R/4BQK5gxr2Qt9JfEtaYs3pQz351AcY+bqhKd6+Fv9Lly15+eeloDyFNXWM0UKMh
oKXduhQJ+x3KCZNZ3riIW77YUqywJ8AWjwMyImOEX9CitDsUWez2i9ocF2FIlXtICpEtO0AXWkrw
S/0x+4wHKJceWdRC41rMEZHfGUp0+PB8GFFPFuUX2/sYXxoceBHPCGnuinv78wUCClJ86Zbg/rM9
b+EKp79X9FSaN31JNzBsobpIYTzE+qThQO+jTrh93zPwbZL062yvRxz9hVnlPpA2epNz++DZwFE6
+o8vXgu/5oTgnTjCm0DVagjdqTdB/o/iVn+A/ITObOUPv4CXqtuZxJ+yBHzxRpJYwW4aRPiEGrH/
Eg2tW0NhDZQnrcTuMIygdNZCE2wodxLaWoam9QIJMMOwe1Jo1tS1DeYEIQolcLb1nipkg30x8Bar
JT8oa/hXz+SWMU95ANh7L1rkSgP78CMATSDfe2jOR2vCqcDOXaocFuCw2jqu0//ZQUg9BNxHnhkl
hKVuS+hoz8Rfqg/I16zkPEdwU+ttByWQ4cUnES4CtIh0PAE6egOJOo34yaumaUWZmnoF1i7nU57w
0IeaVdrWOoUG/G8Cyyix9rLbQg0dDTe+ZC/0AYfBSRKpA9z1on7UAByMMf70H2TNBu4vDExmpNo7
5ELTMi25R7xDEGhFhaE0dLKzluRCshOP5X3V3fQXeOqmpm34f/w+Yf1o7MWlPXJSw586xiNnmKjr
hYD3oVlW1pcIryb4v9F33D4rOtlLYLghQ3vhLTCDGDwE7iBu/rA8uMzzeQwehRwAodmnuNu+oT7A
BtaBBCAcQALrf1vkoijjXq/KpheexlaDgdbAsf9g2wY9K5WIaNcdJtO8WO8WPK8X1WTcGYfnyKjH
JMiGKAwpYHxjDVk+wEYZxSlWbEF60oSiZwReRFeYfs2nOyPIc5avJDZiPKNPAYIVrjaPGzXv51bO
37TSqESJxXONsf5aA1gYgj3LK53gdKA0OJ8oec11fPpn0i5NWQk7pw7V+CbpQDMYUIbIUFQ3yIyo
PnYbFZekDmUCck5xgu/8TC01o8KKoDH861DT+CNr8LAGteaL9KOy9x0fGTwu2xTaenF/vgESlBC1
l6rD3Q8Uh0FPsbcGIs4JVfOMF6VRo1lEDJ2kDDJ/Mfvus0ip2IiHsvTN/51ivaq1CpnZCWfKVAOt
/Yv3bpWLQ65anq9CW+I9/F3ADyzqHlBg8M7e75yPkMuJ/D4acV48lcFEOlcUIfKPQhcfVkaIEF2P
Du4qzTVUGXKiLPjXgv/NVQ5nSnfHJk97v+CrpcOdkOdjvXRK6hUVO2RsES+UVbmm2dFdsmUDf+O2
EMYOouZlFKTIKoVbM0BW6vAVmI3HBOTFGnkGdSTb/Epm9T3H038lbGWK679lBxKcu//pMLZlGojx
keUugbLC1mmhE4jstRoYOm8Z5BrUv2ggiMTkPojge+gjpVij8ju7pfUSCRKLOSGiWiZcBiQRZiMe
Cv0nk0X/MM1dzsTqSkd4XL8+Nn4RGWS7j24Jb9SP31ZyOk306q0Tkr4jK1Q9BmdYMWIJDEvaC4di
lGlhq9Us3PvrMZFiUiLAf7LPT0ZuNvxnx4Qq/y6FiVP8UXdKOt3LZfdG+bfBLC7HWNST/RtSGWwQ
WHrVoh1XS+7ttMhn53/T3LvxMdshY0+lFyHcFcPL0QH/sRcNeML0KB2+MYldKZ/3/Ro2N32Q5/XY
TB0w4pCrjA8mwfbYOsxziZ9HAlnvN6/k5/ODkSrzP+g+FQgqWh7uNYo9nQxPzYWbNfoT6AN2b+m+
GrVhz6h9ujq6ATANlgUNsckzutM0Bcgajcds3x5OXOv1eEGIOWaXzfytGOF7YFTnPvjibpAFtPeF
xPRy1ro2cv2YBgjyMPtlFgL92SCZZsJ5S93hrcGqlSUclIo0R6dU1raUdEWNzhl0u0TLg+Ko9JWo
m/nlkqzHoKfHj8cmUuF5IE+5XEMeqpYFgWqRKvJOSHNTozwZN3XeA5qeGZqcY9UKbXysWNTIrbsN
UzEUgPxaL2qzLSnI2yWAe9K9oCfswV02BOFR9C1OoniUbIFRNFscJ2vNMIFWbDmBWZYCXnzldwRe
CMOrr8swg86OYLDegZ8G8W/E1wNQLTIibcg7MYRm4T8Y3AiuZmJ/7bqZXDVjqAfWJfdHdwmJEWDf
YbdyDsTChV8G9cLbW05bn2t7gNRzPjcaM55KjI3mCq11JECErFTRtDR66R687QcS9D4gqfV5n2bp
wqkk7h0E/GyGugvFK/5hh2Y4AMCOdGCCAVoJL+jWzHRpjWFyf92oVuUkuiNizlpxHrXu/X0/REGR
G8v3AFKzmT7MwIOle9ujOM9y4owfPjS8fYuFOg3Q3yhcD/LjhqNdxELdX2JGiZjtcQHgTz3ZxcWW
d4BFfEn9OKRDkAAsZsv0qhRvyTyyK+JzpgWLSMvJcbuVCM5qYgxVr6fkSZzstdQWRj6kfMCPry8D
3Rh2Pzw5jR3KIRZnvf7wnBqzepdFD/msfZyV5E5mV9o/dxNJxEDeJbLsQ9o3nqfmDX7FbvYWAeHS
EoO7xY1zmj6qK83Si376p2DspMoNRlN0fNCwsWg+VJ1F0tH7lAuJcb4FbfGpyirh43W/leMU+JrH
esWFOoxm+H3pKQSPoHHzZdsyaXzsJnx7K5CEOl+uaRYwSCClpRZ52+8c9x28z0QPGeOTMGLZhciD
8J+Khwt/yLX9OtHD4kz/ylsBChvImYzYq1CFNJc1YDfWnK4sg3INPJ9LKFzEx9s6a//W8vNC5tag
ksM+z14YcqVvIpVR/sp5m8srQYDr4fTSNkwY3/p5xUSZuWfXUXqgkI8WY+N8VaTi9jlLNb8JzHxt
8BzE3S3Tj1x5b94qpHBFKHEG/PSM4+InRVrUnBRjbf/l4aUpVannrBSt6WhgPsIg5UxFlkIkibaK
tzdb1kFPoW2cYJyX48c7x1jVmWc5lG45V2pHbH0j52zITaTzwMrkMmH6zVpzrk6rjom8V9xetOne
O2kjvOhYs7JhVU0f7XuhHdx6iK0faQcceAYjDeRq+l+7JS4loxe9euIBgUW+2JXk4Zv3xf30zdet
94fUyYjVpscuQRdf9pLL6v10yqgTqV269sthOSjse1hnL2rtkjqCdfXTNxkttUmOghTc/xNGjn3Y
zKsqJSwQEPS7UpUoLIPfZR4TrbYLcj0+e7N6RevW+A88I8fSO7zvuKqOjtgidA6SqR6ZfptVREfp
VKq+hT5++aI3ztlaZhiimIfPoAKE0tLsYqX2HDKYKkLwMaUHwTI6Ksfom1B+pVZnE0/1/E63aUzZ
E23Beu0qhcZ06xcJNwnsgUFrG/cN2a0qxvxcU+UdPcOL1uCuBNEkrOyljD5W43NHNMoYBp3HSS1z
84pvznYrNsOxGddSgnR/zSm1MFy52TtKO+9st4M7/g8SR/piGFZle76qGCSjbqK2ayha2ZcjRFDV
EgnIo/FzXlo0XsPORD9WUnRPeX4FBC3L2/9qtVrqBZO04ZHCAo6yUre1ZEf82LtMHL0oz9qrHuXj
X+BhuLoGt592QVssCLzjvWU06BY1Sh498180PSTVRD3vnpOg4+fTLKUTOiDrdmIKRjzhEWVmUCEI
Rprn+clQ/mRAbiF3JMDWkGqTgVxOTNqi4siVRZoAGCDDseDj/ci9DanJn3pT0FvIALnZ6I/q6Vlt
1hRuDMYFL1qeKlEh+y3Qwixcms9qt3txziKPwv/Els+ZhQTLC1ODYPj4mdmXA6fuGrevhgrJFGXo
StCKZNREN/87QYywTmOJ5/rH0dfQKIWprIItWuSWVpc62OD3JYzTLWcZm+HWxAIFtWYZt68cfTcM
kW5YGZ51HbdLnalki3JSH6RFhbD3pAIZyC1Oog8CZezjlIEmaYzm7a92W9+HjGI5seReTF6Dpmo3
TM6fx9+GaGmxp/eF8U6qYEnA2e0TZcmZWwVp29WpMuB1X86LMYkGtwt/mgHQPwrFBpNvNP+kCQ+h
zfVoSbzNPhPiKqbPJFjB2YrVGtCV6vgvvGJHMIaMC4dFArMcbzbjMh74jvIs1CDZsPQZeRKjFg9K
ce6ppQNW51zysjdNL6R/EOzCFLlhloctn8RBVhbtzE34yTnCmEgYFJM9A1EC2hre7mTCx9NZze8G
UfNpxSPzAmRG3htvnpeYu4tuEZeEGr9IQTLU5icEcRpV/fklqkHwKmcku2sRqH+0R/iw+OIDO99k
D2cOawnE3P7vYNmSEZ7B+yOhi96TbeVujh6DFAZ3xg8sNBSQ0bvF44q4HtdwU/EW3zckE8RTPJ8G
pKu0wiWozNEQzmH0Zl6UQND7/8tEiUIVRWMMJZxhx4/3PeYqQwsvTIZKh8Nfcal5/cAT7rsLexwc
IpuABdgzZGumdDrmd9LzeVbQ5KAOnDey0ynR/Sqkpwsj86D6idfYGjjSQ0fuuJj1nRIIKqlv6swI
87Beanga7j8J8vufF4cupRnRsTFVni1sd/yY9Nqqc5eEmVF8JevaoCKZwfRO3cP8Zu6QyQKKlBfg
PNMkjx9EQVLb+GyRaV077s31FVPdOwuwrH4ahVKbknq9T5Dx3hUxTolxRZzWtC8uB1taWamwjTQh
wA/WHZ5F5YN1mzz0E0mYqVMRiEUr1ho13LKZd39DtZneOSPDlYW/I2qoic4CUqpo43er2/5BZxZi
oI/LSB4hEsFIWtRkbkKD6e62Hfmxviokm6sBWxeQUgSQw8uE3cGbRHji9NqsceykO569HnBHytf0
NvZp35N0NJ9bY5sw9JvwDQgV5rTBkPZIOvY1K+tr8jBNfbYH1f+bWCWLgKV1WLllA9itN4nRBHYZ
FIi/rnBu04RJdJwKL4dOQhOY7uP08o7PGbDQLK+CEbj+dCdrpQ7u/gc6NDWmCpBWWLOXEQ1ilVUh
/nr8W4V12onWG5BYUx1kipMjbKRJ9JwvbNyr+jWUm0DBgaE1iWlYJ05C2dlGq7cKG88a/RI43eUA
vd7v1qddHUld6BF+ss6LYkENzkkYZncm+kbwEzQbnKv458sw+15MATZ42svhcVIsMjyPRr8o+HI5
Z/r3SB7VYAi6jEGjiuf68bkPpZ5SGp4xUvdvhfKAacC9GVM3pWzWEm5qt8aND8y44m9wT/2+Ga6X
isUMgkPx+/h/bXrClaSjJkqM8geVBd2Khop/ZygFsmtvDZfCCbNKQgytF+ufW9MqUikUzGwmrHxj
mRj2SSVuLSCkhQ1EDQpGOzEvsrktbB7wwgWZ6+jCGuSC0jsNLNGkAWY8WNTM7KpAZwF6QCxC7VJ6
ALFmR3ILM0PkivrnG1L3lOlHsxd4Hr37HKP2yRWYjawcFwT+bsVT8uFv7uyZsUS4EG1nLg5HqTvR
wbpVJxF/5MqY0JnS9vW6c0DPumG7ELmGYj8H2aoy5In/3OafTMTrkPzXnSw+8E2Eda8/KHy6RofB
VeNeVPMJ/WXUZrCnGoHbCa2YBoPZ2URVaaePIO6LxJRNZAEfM3xNPDlns2hQQYqih6xVunndqJCI
wvYjsNZt3K3FVLZHZNcqths41dltG0swJQ1EZOr6wqPuk+HCKCWshwiRa+xSrKtjL9i4ohcjWW8j
j8G8Ul47TZ6+Sctx+x0AUa6RQJXTPYIePA60M3ar3junn66pa3Pk18Ifg4zn0Bn39NeUQ1zBpX/Q
Pl2ergkSO29mRN+VdBr3UugqNAS/I9RMSSP/EI2OARjt9cKuv9qi+lFLHvuHgE1MqWve2h6QCRKi
PjMb9a+YpVZAIbmEQ9d1l1u3yvR3jywObeRZ3Wl1nvkxhUniJqQ8TNW/jGfWugMnSFwA8t2mlTp7
mCj4mqwLL6vRacutTPRqpN7OxAkL6X4P7LuQxCGefxBvm4/AW2JFeZScfyqDbaK101WkMXojwP9G
IQuB0O4Ns1WtXfd1WOo7G72U8ZapgVXqMVmozjypl/aeVL5ajAk9hDuV39dFfXtjTSL7X6nPwTYk
f7Ihv79kAOGXEpbMUqMrT+mwhmJcTXu3lia2jruHvo685Pu1dj09zm9O2lbttl/9pWKFLLEy0JxD
1l6+uaqayWB3PO0hZhZ3b6FME0NlHxRH5+8aBYaRdwL4gDZmlceAQ1AIMZJz2zoVxJrpAgGyKPED
vk6s1SqRgEOcqjea8uE5KBdEburpoUSOLZaw5Qrr6Q2PRulABfa9CPXUH+O2H7vbThiQDFWmIgsi
Q1yTDuqOrxtIG6xX6kHKD7aGw66wfVagbUUrWhGaUH9VDgBbaUamWMjPXtYOhmYCKH8NgR5Jfipf
GlqbMk1rk4YKR4Nw1UxUe7L0WhZ1rdcePwpi9YOP0q+YdO/BBrj5ps6Y/vNKG1AOQJLZ+Rmx9rx1
oK8L4RpYa+Us6+R8TsQS4ebuG3n8Hsp3zK3ljjGKE8Ww7rnd53l5qw/7f7Vs5MYf673Cx6lgWFA+
TBjpIbwNeGMpKYV6ZyC2HmGkUWeN8N5Wv8lzyc2N1qc+s3fBvDndTFoZ7HlxGxSX9Q9GhqHvVyT7
nSFjy+Yo71chAMxAXYWZ8U47C5rCRhQIwVuhevzFl/yBMcx7fmpLzuievdmWujBTczeIk3yq3qix
PendYxonfXDhBA5ThtbsYK3lnDQKVcSWC7S8q+LwakRmIEF3IE/Vx8wb6tqZdUb+V0ZzFReDcsF1
5eec70zTALwBUlZR2ibY9O9ZN/B9Nc/BC9iWvKeDnCoZ/G8ZDOh+xH/agWMsMMGhirqKVdkAxeMA
Iqp6AlvGsMJp754XNOEzE+nXom8AxK/kYXMTANxRpnDosQI0Op5MzREaJV6g5UMQxpNm8r+vlIQk
6r1EfS910o/QHQ9+bVvN35m3NkJYIGUDRLDdmSDOJN84oMHYtb7XG9jPdpyRbeL1qLKqIwA4zKCJ
1RvZCkHV7NJJ0kEh2IBKxJOf7MH88e2yDoExlxSUsbpgZtIXkI3Gk4GKFipckVH6gbte8rF65NxA
1sfrIVNMPcix/sIqqf08gsZ+MObosdiykxiJq7ElfYJHjUo+8jbtE3jUJWDqyskCIK+Jni2Vw25e
YAxNeCRXtutdGmdu2VXNWA8BTv6AwPdpOzY9G26b1KmVumZkRpbmGDkjp8j7A8rKdhuEzsVLH1Md
sEwSUFYl0BKpBdoB1piPYbRqKinQ9xL03H6nNwJST790/0xuM5trf2FD7PGIRSFz2FUn8VW5IkUQ
srlpjmXiP2mctQY724Bb0KDqvw68lHMmtk806sKV0Dbu7cUI1DvX2Fvfp8I1EpeeqXlHAgEntfBQ
lurAAYFMBZUxwaP94epijXjM+/gmThDF5IlEoHowI4YRFs0rNUjyV3q5SdwAQ+KbXLE7/HRHOIw9
tJiP3LreRP51txfPbK4eMjXqaRcbh+rOLx5ME2D+/yTeM9HhDrYrgZq9v7wUfGL1FxTwFRw8jgja
0QrfzqvpnyPHJg65dA4QCMcLu8G480jzYuQ5+7jzRZHfbzugHBBEAu4O9GvrflftXuby2b+d04f6
GqAcNTPqsezdM5P6nhgo9qB5gT9nxCdED5/vrZvJTnmhyS1tiigQniI6if8e31VxbWZ+rhu9trnn
tzMNKf/VklK22mAE+ASdTMYRv0uGqSlHr2fiJFu5+goNbsGMnZaryQmxXgBpSMcTUmfJEqGzbxcI
8sqW+h+MamIDVbyQSgKMeluzDM64iweBIl91Bzge1Fh4LpjChx5C3TuRHgepJKLmzTX5lHEH8aVO
RP/qid+eu0lKxNg2OHNq0+tNMUEZbAvklblUNZfE0bFEeBAVugW7WZXwkELcJjjIttUE3MNjhUR3
CQpQURInODbAXQQ3ste1SoqbBD48ywiNOtqQ91/XtQSSFSSdCWOvo58QJ7HDaET5euID9z6IHowY
b/bqDqMaaaaLfFmGcQMCyFca12baI8lLp3J2et3ZfonEz5rurset/9pHxazCjs6XOYM26lpGVCUx
sdR/VGFjKyOULIa3QNGaPgF2wJOZrxLQis7NqS+nM4gQdkyyrw8bpEUph7wi8unUjeudX/X/Q2Kt
sa39RAB6xpuHXUnJ7q29E2GVJFrxNRGdv4f8e51U/uLMpaFXnhU5XCWFDCN2AAJKTZxleSjQv/ug
JHNzynNWYiRWo/PA6I8hbSa7bYkmKUyAcamZP2w5RGL4y4+jnt8fHS1hxnIXp4fbIaHex9sxSVhj
oUGqQ2jHH2M0uffSuvPEn5ByUsq1hVaFoR+o4Ckn5fnOR6jA4OFs3dcDGW3G1+l+Q+yXmjHm2DS9
X+fErhxNtsEnYHbcRFMXtYc4rV1J1j/thCQB9GBJ7P1TXLHg1W8ClfP1spYYYtttTXP0u2qZLFzt
gynsm19Hb1zGkwT6IJmx+8mgpcBuFI5IWhxRJOZBCJLus5802w1vV4sKfT/gIcuzbcw/1XxnI2ts
oqpt9vJKxhKxjAmfSmDWbXfp4WI3S9/tsZZQBiMWgNbD5NzSA5gLrwpD0HoqT+1gjnJ2yu66ka5j
auEcLuEJdbY6DhVXSG63k+T+YzIFIlAnLMhblO2qEOUhp4MZAqDzqHRRilUIh6sosmQvCDHvdClr
AVes8koayV2/Y/kJ4FLPSpEchh+iZKPIRBhtiQmYwnKxpDky4pnMmuJPvALlonxQ1MtL3aLkwsng
6Gzre4CBJ26/nerso7HBreq298FNsZVUHRRDC9MCpxIFP7vSptQv7fSnHBHE9JWarkqYdwK+FIXQ
gVWB9+Ye3LkbYJVOerOePfrS4Y3mtAA4QwCDcJHX4czJB+kaftp3oiFywoGpf1tuPUm3ptOkGttz
zeKx55Xva4oTxA0mORPklbsdepwjghNq0SEge0WxFX8/A7XFQCVomjAgolDTbiW3GttHAkFwrAbh
rrjiYruCEn1ARmgO9Xo0HX7WtX61zBqpqRX1rKK9q+z3Inx14F94a+VDh8gLuSCNx03lVasQwHuh
iHjsExEkXAtKzFW1xw3t8ocfmy4HLwHHZGRvmxJuOJv2PlbVfEUqcQA7D1w8jsaqnVC/vMNonq8q
WkVF9cPjQzBjeTZ+oqCj/aPlZF4HavsecQV55UWh+EIXCifrrQiGZ0PGsJCbyQIHs392Q98YmLeu
24dfHVB/E+rA2BAs0E7ksjq9katHQMujNCnEvTZ5Ugkt8U9SyY/FGWFUpcMYzj+bgqpXvchGEkmF
cPNTBuJsnbNvqOsGW6n+rpSLDpoj2DcG8EClvJHFRYAqHjiWfBYfEnGc4r+yXI+8oNzkQh+czek6
Xu4mYRHIoxxtzUdRZTQTNypMvmPVN5gsBtpFeRLXh68epTOckFwrAR6hH5mMI3tLZNN7CnQZ/UhD
NJcEwCMWu8k/HxteqJE632jMSaJlUB58Tt7OA4BTAFLu29lVvIXQN+AgUmJ4aVDUzxKW33KPlBxw
Q35vi1e+FiAR6dRci5gg6pdC7S7gYjNpoDjfIbTYBDsJiaLjEuCEYUu6aDlWvzGLkbZ2Lj8fjCuk
octk5SlAEuNXHSkJY+/J+FJAoMTA5XvyHMc5vB2nhaiYRRFpT5wX+QtSxLWV6vjK3H54Bkzh7lei
6Uj6IArLhd+B0cORv6ikfYn4RYsLaWN0Y4ZdEtD3+yZEXaMjh0l+30xLZTdn4lPaSyAF4kJExkzz
C+mIcNz/p+SsnwMN/mahs1PcKSS0EKCHSI0gKuCz2YoNExfke3VSqFIzTgqyVv4mq6zzN0hd4G0x
uFqE1RLH9T4t7GJ59+Jzu68xo2y/KvQ5w6n0F5F958cpuLqAuaA9wPDrc5mTUJjA+U44xAtR8UoA
L00kBNNmyuK4ULqmy7fgjd97Qxd/M6khNFFtFhlRusHTT1+EtKVmcu8Sl1eRisrnxINlcuaMEy1X
jV8vHDSTX3bkHMn0wX9X68BfiJohcmr6RxiQfCCe5AdXzKKulUNI8kDS/OmIgAZ1Cep+5HcrZ1mN
+D2sGfkXkUJtajEVPeHwzSn4eIvfNmXoo+SCz7svc0zqpexj2Ejy6NscRtYcaOZJZqiaGkWpFVyE
yyia6bsd01Mcw6x/zl9flaAoIG8UbbR20xS6G5n/gwIAoOERgPyZmNYPJ14e82O4f9tBwcAqoZj7
MgFeLyEaaH+u6Y0y276heCz19aTnnD6c4zGxaYuPfCQdrcj+5k9jivTMuX6C4VAQ/6eqOfKLCfSP
JDafgEXrcwJ/lovH2RVQDdPuybE5/xsQiW5jLQ8ljta5w7Fae3bdQ3PGXGlb8zRY0qoxAnFgb7vt
d+36qJsySY3FhwYJIE9Tvs3xHAdLsVd9Sj0WamAgdeyExQu4h5ZKEvqUVeUWwZGkPZx2ZV06jrrc
1VoNzXy/Vk2BnZp85mAMJqptwWKEEr/qxl3Dwb39QEi9Z1RqFdizjHBw3opYorMcFkMrzmu3RfKq
XiOuEjeQyodXbwzpo9+3ZHV7h/qG2kNU36AuB0izW5DUs83bvO+MidgWPxy9+e5b3vU6Lny6nQY0
Q7KKDyviidDkDK7NTRIzP38bV630y9ukaL3hwFOdQJcEJkSXgQsqEZHbw3lNfErslQYIQ3QbVWvQ
M4dhqtxPdhCAaSMFfQOHVWwZrLX77snGpwCbOdoMGSKGZq4vcU6BuHxt1bOstY+b1q8HLT5BD1uN
UKZd6n7CXHHOi3r+ezxus6wFvD5UxAlT8vfpbgZiSi3lJhKHJCrgXdGRUBgyDPRWEw1M9wmQqGmM
6uCFL59prApjTRsl97aZY9ZNIzPk0vXn+OJXERGAOKnc02HeDlkCQKpK2gC2cN4JXjzG4WXZee52
d8mq2dt9U0W9sK5r2AlG43UrukhOOz68PB/U4QHgjOqF46dzXySJDa3wfqgAFyVTsgNWWEaPpNCR
WMn2GRGjzqocf5AEF6iCC822bqb44WV9nGuAgHJT6oeqU+65t80WfhqCHYbh2pEzi9LAIrVQ5WnZ
Rh70rEjeH/gJxx5cyt+UU7dqSTquDtAnwpgjhKzP/ja5p75klgTjmdTzcQl8WCVbx53YJUgmvfrJ
N2xfZgkZiQrEG7OheUYTQn7mPC302sX92ftlXDoJvZwwG+Hal9HIztpoavHGkHGVDEq62Iu18PGG
qPleUJPTiw6BC0gFw4RDsWVfmMVbjQDbXzYKT6OpMYyS7iF9uCdvj9ZPIYx5qkqffX98KWpNV2N0
tBLvhi6vWMU8cbN0a9pVQJbKAvB+eHiqdKbZnh8jeNZKxNDc0pvSyQrqyGpo0l4uPysBXB7fn6y3
dD7wT0qJtQ7eveL5GODFaIzof3g1R2h06TmrkTofcdAZzGFVSf57qCvOXE5l9B2q+gAZhrK6dZfo
NNW2SbbD7m8xXEmGRBHoGao3SqLoHBLV4wRQ/SEo20LMFBsacxiEwm36iOntnSwlEQ0MMk8BrITp
9WwStU9OsoT+vdpwLWM7VT1eE+r63ACX/DqyFOgfKWtOr/oxPfRFWg4PhXWIwP+pBAohgu6/uxes
W0hHD0R/K4PcUAJLjSF4DTa+SDC4LItKEdm9MgqGn5z1YSpBiplHfFjd296L2tSderkL0Zs3PzM2
m54ofTR0PdZu1bi9dc1lmm38K++Gx4TyXxiBXNijR1hUgd7pA7g+2hQHishq3CML7A6zev0mT44j
OYRWQWLx0jy4x8cRxihddGKxWqtme30Icajk533AZEGJdmabZze8gIT4gUUEiRaReedXWVlIGNUA
GPPq7jF47frR15PC0Sc97kk94ImebLHI/cAXjSRSs6pPE0KVqfmoLQfjNlMd+N8TDiZ76plZ2B+1
qI1FEOft7JlWJaC8QKQQFD9xhdSqNQxX+WZYzCv7SIIYvDhI46GRikE1LGOD9EMoPOHSRnW3p55T
PGtZqDd059/DlNdZScvpi0/0Myuzbpxmm89Y3KKNF09WI8XDK/+fvAchCj4SYa/7rLYwoPs3NGAH
gUyo0D2EFkEaiMitX1bEhUYM1/zhNl9PfYag1o7V8nugwOYB55OWiZ4DaNLAaVbj05CsB5Uko6ZD
IbTXDtUaHZ6iYOLxQ5SltUTjKru44oJFfuq4U8kL9Go+2+fAh7V1dcHkGoDAZq/ffZC6dFTbweKe
eGCL/WxoBdV/Ct6KDnxRfNQoyT4WOsKtlO/F1Bm7IMyP+ETM+LqMtH66lw8FPzfKEh++ElquxfuK
N+Ov+ayg6l/gpr3jyTDJI3FSpHeKzS3KfS+7+YdhRfM9XXybHaO0WeVtoU/qrRnsQ2Ky2Wrw373K
+ZuaCuQB2k7Us7M56Z8iXQHZSv+ROm04bc/gjBpeJuO9rI3CgBz6stSQJhev7MeLuhpArQmocemd
s6DsdxrcmG3rUDs72Tc6GIupXCSpxDppy91mUXgc1N3M2Y1ZkfKl5jjSnnvy3r6f63/B1cL7ayl1
bvq5fzahmRshOHQJnAMqj3X9rt+bQk+5QT7uURiL+VVa6axK3GDp8OLxpkbo7WGe2I3LWaL7ELQi
iCCOELVaoRTkcQ5sKUKac9AZ7AtCGAuA5sMfrg46Io0/A6ZGITojO3GXm/Gfh+nCwLdIdjChuTq3
F/d2unKDN/wXVKv1zp8AE9Yxmc5HfWApOLYSsnBDuoOT6ZbLCJ9Jqbh78edjUVzYJZHfA5fthI2z
78g1NYeq4WXvLXndLpIRprmWSE94D0pE0ghlZIY73Q10axi4oRArNLaBJNXT3LL/feRzbEsRz+5a
HPCdETETbbMjRVD/phbJ1Yv7P9L/PBb4PIhPhWO8d001wpnrzQdh7oiO2p0D5LextJsQAO0TDKHu
MKbEZYqwYo16g+jOJRaH3peVuJJ7lDhTi/wDtjyVjYHjnJcPgopO+Qgn4LSUssyAaUmAUjk6RAEw
YXBKbKDqc2Mq4LBw/aUIhzU5x9GNa4iwdri9jVmbF3kWrzODC1HYYruimsE550lYS7piuKMBfj2L
16oRJXtv3EpLd0FrzBHH/HA2PTMgbI3XmLKr1dZoDUvKHBeg/FZA24BomAZfDotqZfu7lrmHlJYT
XhXrlRyXe7lLA+dy65HRYPLMd76rWdpy7doGxq6X08W3VA5yiJPSWTu0dI3h3TFYZiJk3etOJXsC
nzWzf4SVy1cucA4EWo93UAOEHUzjxvDwMbdJOyqk29od39KOsyt3S9VF6Vwi6lnCDFnb8loria0x
8+VXeTtjEkhzQd9O7GSgG//unuIEvDlLTTRAeNCuqn7uF0XOcfGGzV1wjDomszCmKJ+I+9Rr1Xwz
qzPQrOZ+cDLKnQtIW5Zf238TpHHCQ/g7jL38kJ5bzXs5x0jhAQd0yLiYcG9ItWmKyWtuKGndHN7X
RAJIh9Hrtg9f+HWT3o8voxctX3xIVS3/2i1Kamn5mt7HyuOHyZo87PfYzeGCruRb1RRgeQDI/hGv
dqd8HchG7MhlEO05LDQJ1n2ucNumpiEsWQkAHYhaYbNqYDr20cZBvrpCAhsderhOZH5I64N7GSRq
MgkotyHzZXMjeGCjSVYsroYQ7AjR7acJdsmQmtgZ0RV5uxQ4AL98EYP0zy77Hwh/xKYqlVftN4Dc
oHUMnU7ANJ1EQDceb/DH8b3jdjIzwI5nSZdrxzghh0QclVWck1rs1OqKS2Q7bgpJ6NPqOFC8Vtg5
zbjjiJ8mklOsxz5RV+nnx/exT0yo0dgcTKDuiVlJeXsz1pvidYtbrbxqj88riwWrmSXmw5gRvQcU
LKFE1bimEKRqWiaWuQsyUUdkWDQsqPzkVYQluC5iOouURf1QZY+lALnNLqAm5z5pLETOR2fJy/a/
MNwvV2LYL3y6aGyZHha1Rr37kI9KwSvaG2UWxZilCBgEojbFgRmWB5nVrBoV4AAIC+uqytXoc+NC
vIujPtDtZN+fnvzRbD0L7Z7s6iJd7OYhAATT+psdEzX8Bx2E+opG06UAvAEsUMXYx3ToPm4fKNgj
EX0BmIZap42JBn2Bqgi2IAxst8jqBnHEZp2SY1fgDSo5xJZ2xQYI/5fKePGx+4QKkbrEA25SuLUe
FJ12w5KR8EGP+5Z/a/zAjw2Rot/7dWYUMQbSVtnBHiRZALi8P0zU/s1C5VZBS44So0RkYkdRICrd
FTFmiFsRKvEOvTGewwyLI+wco9OLzg7N1wd5GVzasMA34e85DC0JSq+DQ9wo313zzj0l1Vw+Uogz
Lpn69AbQeemT7toGbYgIfRa81IViwP7soyoJZjgoC+i9Ge3v+GvsV5P4iOkUOTqYBcltSxCSoBae
Lffotc06d8Z084SJ6bCSt+iSN4w+axTKpaTZPlt33JXDL9zMtAXaMZD2traNRKk6xB+KhafJ50XS
2KF9wBgcbiCiFinMXV50RnqzmK8dI+IpMyueJmiS8l0sm3q+NcS7rMedV/IIp0/9Tn1flJSc/vqN
nAE4FBFG9NmqZGkfb1XUll7L0oz+WvCBu4FOaue4lHQlY3aBdQv8kfAimKYofxpGO8bayMatTyLl
czF+RGzlOe95eTu+5rZq+MpyRoehIxWoPilJ/zsAVdshqRWWbbpJKnxxY702G7AOISJ7J+3JHigN
lif0+FBSVyLlU98SWS3yCp2OGMmtyVN6dnJMfFixe21FTKIIobvqXlfl4jay54wy6+OenTUrDPGD
4LyATwcA/nraDJaCzTq9zpnqojD1mcZ68biIY+hXnFgiZQWyNS4JCV4Tcgwy13o2XuysZXAvHxuc
+Rr01lD1Z71/s2yjSJaUbO7M6kOM2MOPDj3dgjJjIfTJuAZkZrLOQAV7KCKWL4/ruaPstvlUeVN5
kd8ufcVjjPXvy1aMxrpkSqBhXZPiN8iDB65oELJb3W1SIK4dA/24v3AIMNbVYdOR/uIiFH1lqaBs
qbexDU3w6uN9LUxiUwPo6TT5LcU/NuNxwS4AG+nDcj3dATwUtdgzYTXATN9iqwNdC6MXz8Lfhp0W
6VCdjqRiKrPMZR0uZWR4IO4RBh/h9lXI9lQTuRtemLBDhACVqYMFT+zMm+GJzs6VHB7Za83xheHR
zKST5WVptuY00MLncdKpC8TJnt0K8hJohrTiEG7YI+WpEPir9maiJTBG6cHirKwfDac8WsuZp/qH
DlXCErfQenrhV8BViIy7WY2Ll36aCSRxsOi3PB8xA/DeX2P8XS9tvNfJD3838UsUKFO79ZM6c32k
QqtdV6WN/nY+X/l+gOLpV3oHn7G+00WSMIeDAQFF0q5g5kc3VVwXkErkfReR0LnMzA8M0vDoJdwm
gbxGz6KoXahrjCFqbYxW/I4SU9d7dXM1RI1U6LJ/IwR3aIHMEFsJhIspWRwJmBXpg5S+ovTOJO6/
MZWDL9MpcNMSkk7moacMCEbmaPUjTisOzvz7F94x1/8mxJ8MKkErH2fH8/fghbBK2dKSpahfBtHh
OS3jZRpqXZsWi9CAvw/LOyc+XYqtDiwVb7CYfAUsTBd8FUe3v3VYyZM4h43oibxycTozI2uteEm6
YfAR82bk1OLEKr7MMwFF82Fu8KhN1uXh2YXf/GBsJ0LqR7h9ywN4jJOvNscIxHeqKav8qeDKd9za
GYQ4ND1uvBw5FbCSM4DzutJuSPEcMGN12RYfj2EF+E28PjcKPENdjeffXv0xeIwllHhjbkCPKkjU
jQgI1crmHpItz4jZavIXhSEHS4EbMHuKxwYK2OCZW5qtbii/8xuyn+/y41qPfu7YjBC9hxgjmoD0
yPZU/WDGo5fRUxW5gV52jup5HH7HtZP1CZqV4atiRE2kXb2w1B1BfzipHdzFi05TMLH5HN5tC3RS
OHi+pf9OvdsqyygPFB4lYFA+LZZVzwWuR/uQIMx2X4oFLbg30ynXlOyka5vcrSpCnwCyNNX5Llrq
I1HnMlitprSyiRntPOPlydkvxysN4/UNwX8QP+FIUPbCwc517dkLGCcwkoosRi+91YKEmjLmbXcb
SaGgrHr98P96Rp6ULjt6lLnkaylJ5olQcO0LdkrP9nsrU5sEsGE5eBo0pPoylawF15/EQCMZyTHn
MbJrQBYFTzUcVMNiLibI8vuJRlUBnicg+1bqfNqEGqAWUfooOFKd7z15374yJwx/gCyYURYc0QnM
lD+aFVxGOS/cntohIIu+b5qPziRbjypPeC6TDFILHxT9L5vQ2v58uI/ZAmpDn2ApY5m62jRXUXr4
RW2PlEjayTE4igxKLk1ZvLMe6M/ghHFNFrHN5Jzyw2KmTcDS7U8yZCC5z8wfCDr29sUUPywtOgSb
rg8h+y3L8XWOlVjPQd1whYJWApfUtHL7YU3iACmJ8qkWa8SEQI6p4kBL2rAUVK2/P+jY7oTkVpwO
3ZYDI8dn9sKj4fR1yAd8arHEPnDO+GgRzXmQA7s+ADOOYxJkOwmhMum4knuGNiNqRGSQVlb/uJJn
SvKYcDs+NTQnrry+SbdaSKj/CklVfMtcQ8zXXiIqxaN7tVRDh9vu8iyy9LMS/WB/APcrPDgOlW8h
kH0L6gzE6XJoqpKOH6TnRK2pIhvg00XGo/QeiLTqUB92uopiGU8Vucos5U0Co2W/2L50nizOfyp3
+G+OHB0dTf34vkx1UtCEvwRQKcNMEP0DjhYvuUU+yhIjCcYO9YHwt5FE7VokTJ1kX2rg6V2YWETu
ilIUPIaNJK1ROn8zb72HOdUGIlmzT2QJGMPYdS+n9v6y3Qe6rP2pg8ue1TGXxSlO3LtMQKCM18cS
fQmr+DXZ6DKVGXRGFtt69w/fLaMsqZYIynL+tDMfAWg8OK/doHirb0LXTzEbDgnjiev2g6T43eWk
hk8dwoygTn41ilSd/W1onVTh960C/uUzboG37azaKMkkVvfphZiqS0gIW8Ae/tEu4cuQSowTbhzn
bLv4lFBGr94J0J3l7T6C4nLWhKSnnRmPNltMoOEy4LtXM19y25xDpvr+83wzDf7MaToAV4SfjQfu
9ju317wLDgeslt2wzMecG7KKb6sci30+fuSyS/0dIpfSsZCK9fOd/UfrvWDE/msFPtO6yJj0YSYO
V2h+wqIjgAiOILTGlVFw6Ae6W8YvMSpDbLlWtw2iSTF8EQi+R5boHHL6+VgxLPLnyAypmBUcIjRB
BprMnmtSgLHmmugjuF6LFRvKIWcKY0ovgpNszBJGEcYVI5svqDVPMrid21nbr7N8QbD2XBs0hkd/
mIpSijbes55FZK2a+VHmR+/OxkvmJldk7ith3Y+fH9Xlzq/bI4r7D6ZN/SV1Z/aMgLBjQ9X0iHuA
jyOtvwB52cj5EgDS0FSuak24M7FPTeVSo5lPvtyRv6nVfGv4WiYeqP+3w5ckIlsswb/uW7rvG5Ea
GD4WamMs7FUd9N4Vb14sFQ0JmgtuVXMw5QRcUc8oMxuaOsYkplf5nqiEwh75H/gEpL3vxWF310+m
x2rrlkDz3sXjPio07m05wPVGVGDETyZV0rCpn/fbkSNRt0vrozwJ0Nfc/MvgKhn5XwDJx0BLfbAp
lFWc4JR8K0mvy9BiLZKi/+pSA1XhLESDfEzx6aQ9G7iVJjsEcxVCjQ4R3y+osvT+siyqLnS7MWMy
s8ek0LGE9YrZriOxgpoKOMMSDqy4lVZS4yLyxWbeDbejDYhB3XeSYsviwJJDgGAu8n5q9R27Bu/3
KikANpTgR0MPEKYZ2eZ4z5wh7iK9hKDuduAKRHDevZMhGY5YZajdDw+/dyiQSYpFP/dbkC8DuISi
0qw7OZF3wnPtxhpxOB772wot8txsEG5Iz/oECq8iY3hjO+fK0PvPJiu9enELGPlsg+CBQjrwfsxx
bvuY5mNF+9iam93pdQDsDmtwNL370bTfVO3jLhKO0Ytr9JQXII6W2CBgPmAzlqDIi5bOQTDmQTj7
EXRtG0QiYPUDrQ+TKc0EnLaxcsepHZR7p1tglt9PIpXZGMRzMYPppu9t8UNw+8f694Nr+ItmJrx+
+1n3ZWci6CCWl6Qw9WccT/ih9IPfxP2Yda5HnbWdFl/DR5fNb1I9XEoZZMlvtMgORc/M3kcJnIVN
8XujRZb5Y2QkCerp/iDCSs9lSLNVPbUWkL9/wE+cLKuZLGiT3nZA/iln2GEeYm6IR+12TTfH7mIS
6JrKyOrSQkY5MGyS3tODA7ElnJIm8kCIIiMwSD3ZhGdJ7IeOynrr+B7VaPHr+yHrXrRg/5k3BP45
dvzXSt9jDaQaDi1b4P3+y5HoAbmworTXnoA+CUPPxyX2RA7Y2FpFvbxhdHYA5GMbyJ1DAwMm0H+V
bAzsSCTVM0DE1xqpMabjAPZ7aOfKaZstQda0oqdUs/FQIJ/J6/v9JZdlDNn7aVuP2gdyxIh6E4t7
NtxssXesNd1zaaeH4OfTDSD4pZ45+yE52a3sQNiTjU+uoS0lTugwPKYjrwW2Kb9nhTBoyc7TZX/W
/Y1jCiixO5/qusBXjNPhYtief/vGXKKLYRy64FOmD6fyMw3YUutCUujX8mB/423sanorhmea9Lmu
S0b/VtE/3ozcL/1501LzCk5D6elTD4oXqFqhIMYrW4GY0CRBif9F2ZRKJVonIzlhD5oY7/119oBr
P0QHYmFxTiDYFvfNFhLICEfYN0O4C5sZHUHki2rtIpCq+QH6z7Uuh2BYLUQvm8RXMu4eg+cYQvP2
06DUrwp+XicUIOoxqm20JoENYdHNDIOdR7IbFFljJhmha9wrxVXcP2jyV/J2/EZ3KxMD+KKTmrAf
N5KnO28PUrsSN/9JG2qV3pn9S7fqNrlq5yGuuf4U/2AfVbaPhmsoUJD8vdzfU/Kxg90H9G3fiSOB
g4c2IhoIgYG3xzHibet1JqwLcZ5+L8ZHomtfbnLHivtx6mIElFWPFpk4WHtSoRrYBH0ZvyAWtvx+
Uv6V/xlVERDO+St/ANC080CO88NdTVHja8r5PUJMAW9uXuH09Ss66Ou+Y3+S2P3I3amKSnoij3nx
gA00MhLrTc7nY4GbULOLkbbkOfrdyY2zkp2+9p5WCsuucH2aDiCGZQsiQRMGEq7QckjWfxh5QoNt
wJAgRqPK4d++cRko6KCrKyOJIykDlW0Ph1Mnr0kJ4yYqVQkP9krKhBKgtLulC/q0qJa6y2/NXy1U
C3fJ8BrnW/MeTH0e4xMaSnlvhzwYXW5nZU6IDvc+Lk/bdT0waFIjxpSi8tfqsXocG8n6oxkBa9Gc
xntvYJyHwfC54neI43Yx6zAZ2z2VlQmKHtLw4Q8cU01GLYCd0RsWLqxecvwfWGyxUrj0g2uudZd4
0zeE12UVxWuV32uHUURA39lTTD74PwsLa0WnAKhFZEqYkETrAfnr1iLtBlM5imiIyVBjf65Ckauo
PH5e1rJKJJKNmROKBOufWrzpWVYNo48Li1SILBuhzieFhbHPCHtsSscLY7CyChd7KlcyJ7p+fkWD
izkXLIvGTNOJBYXTAPJgbHNhcDExqnQDqeZOC8k2MdABSUoWWOF6VW7VjJOOYnCIMH+qR+PH8RPQ
Yz98jM5M02X1bC0/q0opvX/xwD4UbxRM/+qndQwMEL4KRd0G1BDnZqzAM4siZx3aCduZaMefmEA3
VtI/YP0DpBcsiUd3gXdAA2BPpF4ZgPDv08ljzF0D49UOd69NfUI8KQwOKDbPg8aDNmtUOsadUBJ2
dubSi6a/SKe1UbVXBajOZAX4JHsDsiVnhzlvCD/DN9+XKSA96FtkPKYckYAWyX91SgV3PHjysPl7
oeU0QWNJQzaWVHOs4RSayp8A6p4fhSozrklIGxOfKLDFJtoURIVix2mixhV4WXzVB4JcMMHY/Lys
/ucGbuR2BqsinyFjnmRI8dndxsN58qPYy/0cbVPLyWFqWhC7e2Ew9UNkFWHHsAjjsjmrD6IK/O1U
/A2XYlLrqOzKvWdcOYO0TfyLhYQcI++lTN4rIP7stZ5UGb4Z/sLk9nPc7nb7vTIoSXZiGPCJ3REO
SsT7Z09OTSQvBXNDWLNqw3E/rcheFpyB9qPrpai4Lqkm80bxciI4DVkanFo5R5947McFn7bx/efM
ptAgIaZi26Qozz4cBK49cSWO9xLzZwQZ6CUsxKMVtbLn3aSLyAOD75ScN0bzsdQNvj8NiJkcXNZ2
vkKApSQ0yQRqXty75qucCsTJSTLA1AJbHGCJatL8/gVG/3WeXCAkJ1oHUafU0DdQB5vQaHyDcWJg
FX3Bfb0sI4SLCMtsJ6m3VfHyvpO57LOORzkF8oXOjWe33O55Bfnj5gwJyGjlds6viY6evMfwsmEq
IjxFqQPchckNHYsGywgGG60ww9dCcUSm827KwvP6Ur8I0MYRyf45HHSDSqkhHaHxD4n7bwfik0Cx
cunkRhRv5J9Rhj/eLlVNNiPHB+tdUMNaCDvsfl9kdTjVXK82RcfBEOfepBroUauBQIhM1jYrLvbT
0nrVfMc9Wa5QFQn6TXctxzTDqFxuRwIcdiHih0UPNtpt+NkKUef8yLa1loMO2h+Jebmhd1a64dMT
jo7s67qCnFfsns0rhIkqIaP0ml5GfJsDddH8AweI3LEerGNX5RnVAtiPiepmEGf1Z22E8Dg1ARiT
GTSWVpBTrhZUCk+ANDjivVGV38ZCJwMIL6eW5RqDOTplj5Lsrk3TohDN7wIKrtwtRO7YNUw8oxEo
pVRLAgo8Mz3cF1EVV2MH3kr242IVwX6VAVZVH1tRI8Q8P9L8GQZJPWVuzJ2J3S7Ws/ewhagT5pI9
VDSxfMPIoW1Y6ydtLKd62i7eZP7NtEBG4+wbzQ4QW3GawfEb35xtJlipWZh19SO9bf1BSbVrm6xx
etVUJlovdpojLE/l2h2oIkINYyQI010hAL2MKBSjqC9n/nXQ1A5g/WghQccJm8qaHWlfemYeTR/A
Yq1zpB2OIpLYCTLdIBNMhzBhiBr0wp3Qrxhgfb+EdACXH+J+rqqrlNMBQ1CnlgyX5f2PQkKH1RA/
rkqfk7pSR4KaQmSXkP1e4UYPUy4HrdZTW98CRaB/0Xgu2NL4MDmfDzErAfoCD95TmN12ZsXz8y35
vg3X1dnWFs3y+1zpg0AuyBREsugAr5yvj4T9X2qB0iemMF70lix60ajDlkx8ffwZbmq9B734EQ34
MWbPht9iKt+nBkIHkP3P7mgfJkaIzNe6ucfMmu8ZRdOMf3UYlp/PRnDxH69AwDDDKSL+obOW7+UV
J5TglqVL+/CLnjYuP4L196dT0EgkcLPEdAwPc8NyPnFsLiSJiqLisElB2enKZUGuUDfGZWC+IXqt
U/LG7jRu3hTHU2heLLZnvkr8yfVL9isPF0FUw6CmfO93JZkVMlnREdvQRC/3LzLSiYwyBEH9KYId
Wk+4RwOwEHnpW4+8XE/xwzPSHHnoinAKcv0uFFb5opB9i6iD9QdYfrrrEMtSkSIHjj/UEcP3byTA
GZ0m12WCVBEK7YS7Mxn6Dn2H8B5dgqo2L3E0TMbTp3Kd27cghQCBHDxW2lHPCB8l2B7msbUHJ0Cs
JIEX7rtd1h60hSl/puv+GkIf9AxSBqO1peQdpca0umr8hZ2Up+H4N/lpJp3ZB0Owb5LNgxw2EcxL
hqktk+rz1y6e+HZPKqbt4ZHibrAMioVwP/V73mxf7BAqkRI359o8fnYTV5H91Pc+Zfne1BUzoqMa
kFzLsc/LfOrAv/CAvlwEjZynH/SXA4HIs+FsDSlOEaDVdYIBfaplkUzlA01BoNyKrEnDbP/2kBE/
M/lSuhXdwru3s8Myv+g5Ig/wLDDD78ctZyhfQLU5jKZd/OCbPNEd3W/BsuZLTYqMheFfr9MkMvnN
sEzF6IZR38eEEd89Xauf4oTZzni6S5ipf9vXjE27285jjQF4/bOhau3/wXlQxQl4vIK0hH66RXvk
ySloQkPCMYkr76G5hkyb34dCnWoAV2htEgo/hiCleJLkCksvRurh1j9Ovu/HDpM+hS90REx3EIhF
biBFoA1t8s4hHLBuFgCpSCwTguyyxzlzTaed/9zzgnrLNzU+ixSOHAWfOjWdU11eYTxB5SDAx9EF
qoF7QE9FefhgzYvnfqtNBvFb9/0WZoC1tgcrHh1tm/5QKjtyWwmC7WKDGMOeNNfMEBnEZ0UW2S0b
dBvndUGeW8xfxfxYs+XTXhwlzmP+gfILOzu7NG5eoesCu4dHMm+mnsDAaOPS9KGRr3lgFoLyV3IV
/Pog7jeDyMFmNuqvzZXaF7PHaTIBcI+KnMyo+zduBd02QrIClzuq+ntJ8QKmQJXsKnnxevomlXi7
twGvUO3VEm0yZ473B591nVgC3v8EDb89DR6/vGrKFT/U6gagddyeqK9LC7PpVP7xuqK1T/PqFDNr
avYCB/BNx4G5HvXcUV0ZZfew8f1wwWSf7k/NULOYznhPcsEeJG9RMQu9CEEiJ8MOl7VNGWcd1Y2V
4Vo1hMS0f/09LcsS1p9d0kSVthmDg6hMP771/+eEilWcYtIUq1bqnrayParhfOj1Hh2O9NeNec2J
OFGEp6MvGc9cdxebN2U+u4aDFVdvL6N/7cpwgkBfA6L9DWvIZXe892uEnex+vwcEKlx8Uy4gO/xb
VX2XjIpl7RAs/ZTJxQmFytYrwB5GPww5lDxEK27xVviM76pmwNjP+VrEBt2H/aL4p3WE67/bhyjw
Txa4xSvUIxk7iiNcv0dr6cbsw3giPJkFt7TTDZ006VmabEg6UHZ63AIwbFxFusUv8kzscrK0VyG+
roDG6+jqaqWJU6MH+zWEHCyx1Q5yyNNvMfxjc0kPfQeAD2/fRBHB+oyTw2UxlgZGxMSESG30ZN8o
Bqw0NLU2zzlPyo0HguzeDPv3SZTSkLjKhsove/DKehFCNT/h55eMSTQtZ0UI05QnbXeky/jQ41NB
Eeizqq42Ta5WmUH9nekiGK0Y5nKuzJrOHYDi+tPA9rXDfVSdg6fWiSAXHJS3L0ISDg1TBIjA9+at
GHLSWu5YxeSWftCf3WVr6cC5tXeavlHQOwF4e/LEzEBULlYfK8K8aZ/RzitSc8bZWJpcPkDqlcqA
wuL66cMDAZNPWZxKdcrlT+96xoNmLCq/738pzB9lB+pOXRElIF6kocAPY28si18j/98Z7kXy3r52
lv66uoYceb/MpzIDpRfd6ZC1nh7wZc15jKbJXdIcswQvi08ON1DgzblNZ0IEJlkIWQTB6X8mUqcZ
ADtNJxA2r6vvhsJ9qexm4gbAcUxjIJEiX2AED2c6JOveA43mPSews26eKGlmjZ8lADc+pNxpfDSh
TKtOma5nHxm55hMWdsIujLmtZ74mWTMZfEgz/Up0IT0gICsFMDWFvfvLHwEh+8TrjH6vlLCg0N/7
N5BkIVFbllFohsGNI0I2m6DyJWGbkcrd3c3BZ3ukaAUTOqOk8YwlTFyUy9CBvAT6crmkOWN4XAhN
UpdSdxOP43Etmeju6TqoGDFvTdc8jqhFy5mdzUlMKiQ5uSePCWzXs4LKOpoyENH6gGBR/Tr12NLT
p2o6tb/qC9EdIxBPa42m2x5RiRs4xpFcZWCGP0UgAGWelr+RcEaG8YSmEQvu5lNAxgyVvqOtnm6t
3VKzlTOae83h+3wC+v4iEEY566Zmy6hcQmSeawF2HGxEUppKeH1owckTM9dU4VGUfzsH23bO+New
l5qIJ6HOg8lhFatl6mvI9w9tJ7J02aX1FjgckHco4DH6a3y/0QZvnDPlEm0aPO4vhYNh5MsPX95E
QvQHFd8BEBr2z69NC7RQX6fSj4TMklsUlX1IqAB3sWKi+McrUHokiah25azzPgl0tyg2Q/eAB9K9
6l0zRSJWXcjpCor1m+igUi4VEQK/URDpKpKUAzdychD2+B4ZEWDwxWd2C7BEZim85ZwXog3ZTKzR
P0fnkpqIoQ4c3RTUM/RoTBc7okjVt6oRiZtjKeUhiNvTkNUyYZpoBUMLsx1WCxOFm+iyr3MwWI1F
nibBm43T2um5MQ1FMQ2FW75S+zARHw0y8U79ZQMKBsbn5ndql0oREC6Q1q2kMVPpsa9hxpjl4qSw
32EtMb6bIjlbUzvyQqoUloeeZOjmJT1V6g2VcsqsAR23dcd78/Eudlwec30fUYvMbboGu4Ldkh9Y
DxnVK7ulAfKO3AY+jykxVI5F8xN9yQ/RxJt0Vf5pFvpoN+6357JPK/I6/YXHcyjTFXyEhmQnPz6U
+8dEDBkajACENlmPrxxQd9oF14Rl4e6JBJlgozCPyonkHKktlumIa6raJRjvm+sft2FOvQGsbIDj
QUjNEzhSnY0mEfWD3iLal7sIA7vtt4jTUhguWAvBhomcbfaupzssoQw2is8VZoBSIRoiLp70gw27
mDNnkzIfWMf9asLtfuhPMF2KNhLGrZrw5ocv3/pzGUyx7IH7rywrGh/DCN5ZFaFrAr6qxWO+9TLT
A/orDiX2kAam52ZRkE9sZhpHj77Y3rQl0jxYNX1sLQund3e916+dK1MwaVoOlZ9PhFIvsmh4O0FJ
XFND6ufAskvw7f6EfPLuqqKCLPUV8AeL4IFygvhYsXkn7omtH8WoCHTjrbNZG/OffDh3dW0ogdZH
BGmWEcREypUNftlrivbzs4RiPyZWkwUHC6g1FXQXorJInR7VAZ7UqcD7Vs0m+b4WuTUayOEDbwiW
CPqywX/GDdrQA/nWludiLJMulrk8ptNXl3d7uCWEpktutVSy4dG5kCz8yDzXqfd48gbVqtJzWGab
wK4O40ehq1t/3GGzMcfMjlaH9ReIJLeiLzmDJtcoUsvT6YvthbpYzV1cbls0w+PzSRFe9u3Aq3Lk
1k9BqDVUHUYilgb3cvLT/TjT5dyhaGIabiazYAfcC2cjGnEhHZCqyVLI6d/uMoJTt8co1y6dvPLR
/ruMUKbKy7/aBK3220gA284DrAdynGKPA7Zq/AT5tj3Q9eSnjHPwUHV7JrnAlgQvN357za7rg+YK
e+jYdeWVztJYRL1xsmh3aiUU1NFyOtIMHXITnEUW6F5l1zhkpq1jSLpB7rITaWimg0gx06/Z1gGU
OCLjFTOmHK9zPM6r/C9pRTltNkKyAWGO4Uz5I/T69PmX9itisMH/yLoz0BxJKfQk7TFNv/b4mMXS
ybimazVp2ZgfMsDZRRRZAPp+6+Rjvj01thQMLa0Nlmyt3aS2yb+Zhgx1v2zVCc5JCoj2H+7N4HP9
+tP8Rfwqy7h4cDIgloDhnGw3NuY+Bukd1ZwHlkhzgFmRUrgv7thEtcmsiFH2dcuQun1mtcr91joC
mrQYvxdcUcAXqxrq5/he2wtiFKBn2iXmFr0hE09PUZk1BlTj8c2uqpHuzdpQuKI+VJYyCkTaHrMf
2+TXT2rtntR1KMDBo0a98ocZzntlvI47ICLZE6o62bPV5HurtcbsaoOcM0xXa5hXnwvcYSOEaAek
KJU0i65vHjkPLdNi04nKy6rXi/0epanpceb1Lz9z6LT7mDpaYx0Zq7w5x0H2uTGguzSB9pjuVU//
vnDg1cVqC76+PFSTBkqJsL35ig47Ir25AC6pscIdjbfRIRvK6gkn3wwWs7bDIBCyVIp+g4gQKTIn
Lchvri6F1uYtklducfl3HdeZzPt72LX6kMMLtXuXQSbXOqboBolnA2EiCdfZAL0eAZu/GZfjI8uB
MoSWJt2JCcwlaLS1xUroDTuGypalnxmjRrm/XppeKXun7VnMrBdadb8xCMZ/d3eZS5pVF+S60/pB
86rccsVmALojx9+MaFVH1o14mvRuEioZvlJ9VYd/KL1XJnWucXk0Vnlz3EAgQxn7fH/wuboZk2z6
yUG2r1M0ojTV5jzDdU5FmEJO7RCT32pWP9QNnZpyEI/9/htoGO9W6jPpRzD7xBT2/N/9aW+5bQQ6
SP1m7g1CaDzBKvRCXkWO+5lAk1vv0XQ1s3YVR2ZxZhedgpurBdeSfKwFRF0TBAd/RSnVu/c6oMM2
nTMZwVp2L+FFOtasvCC+1SH6HBON+ELXYhvDslRXFMBm4LE2n6P8C1SHkiVawVg6OzXKezahq2Xj
+JImOWQAUsNjOCWA30T536EY/OwZwv+JCcTI4ddx1yeMAISIxHsE5fPvARLxTcXjFK59cnkHkmuX
tTdwsib/WYnab+z8m3cjta0YaQhBNsMUU6DcYQMtNaMNDnp8uEm+avZ40jZkB7OA6N/xbWOlnXVE
RZrdUg61ht+c/aSn8HrRKNSkoDXSiQpKVWd0p4oap6WMYFT7MUdPsIVVRGqtXFod3AxtNWR270NK
B+Vd1olpxA1XoY4Pj3wUUuFMoOKS60c1E1plcWvCyxs/kixLlRIcagPDhNDif8mFqiyXsDz4qh6c
xRKkaYG3B1D19fAju1xf2wh0vowzEtqENXfylnHoU2SS/2bEw0iI9kLmHkS0Ot12JaNHbneyp58b
hqMA+EDQQa8YGI5y+ep6M/7q/SngnGC0odprdmW2a9+QUadtAz0yU4dIs2VPIM4uwZzssjioJ8s0
n2DKZ1xJs7MDcxOeeuFg+M+DdSS0EHxYJVOwKJtz4OGAyfLDhjpEwE6rOsMyPYhhiP0rRPDjeYKR
rI/BsMMjXh2HWyA1n94CoZ1neTQHA6JTaTlTeOvJyCWBCfUhS9dRFR7XjNYDhkFJsdKh6SJPeTSv
ak+5qMh1Dw0VGPM1hi5vfY/PH26Rm0xR8sJjHbzYwqa30mhqhyYAt2x4D8PLolrPXgk4qko3DVGF
JIxEBuZK8PMfm+Hxg36JTtyULPUG3smeNthZXjrthO0rjvA+2nG1idvc7Rlq0UL63vqs0k142xii
NUsDH8R24EXKglq2JBlD52l2+zOYwNYef8KMYMFUi8f9D5xnet/KOnasIet9UIgEEEtAAK9zWiGc
KwLOYcdR9fQUQ4Mg3eeSsHeoSaKmxkFU4CX3j1vhfDGRR5DG8mAwFq8UApTreENoqrA39YoeMU4R
GdlT685Qy7BTNnZk+NDO4mJjibvjy2UaXaDQgEcyrVjN/eSqpfsJOU2+CZdtLecqsEOm3Y4FZ1mj
SvN215mwzQ/Jkien0qobSJniSIZozFCPVw2BAVwjeuG5rtIeodMVm9WOcUPQO0knOobufVuCUwFo
PEgFiRCpBIlB50L7HyExwaVoVbdBIo/2F05kkVqrYzz8Q96VSvR5tLLpcBNYlKeXe2DYCQ2ji/Fa
AH1axNR1pB481DfC3V7yLttLcLeUg7ZgeR85j4EVS7iuYVG+L+HISlYN8livUG2fosxHCBmulP69
J9ipj04fzu2UC+hjXvFta4X/7RVphpc+ROeDEq2x8XvGBUgD53OCQiLiTKc/dy8hTJa+ydvhvUzc
3FyJ5+nfgGOGNSvCdW7aiA8D+pSwBBe0eaIue8WSuWZ226Myud0//Pi6fhUbG3V+INRH9IvNspZi
E6jVlVf4ILyO+UAFWEh7Sw1ZDOS+XdDvJizHmEs5qdmNj4rzVi8/ufE7odUA3m8N3aLwN/hX0KBM
Y15UjAhre34d5YmPnC1ie8v/CuvGi5ofbkV9i7W9+Zw7dewGCGpSc7o4NwWy9CZGiKrPIhweBXUx
zuvVPy0tQcm10gFn2V6q6C95ndfu8XP68DY7EwUu2QH32M3tKRud4h1C5A/+9aQHswAFfMEIC5wc
ci5xevQLOxN0vrQ8Rfv7bz+0edCRt2AQjtEp6NhRBKUpCM/zG82LnAFWWpXoQXZhghpWO9TLTeyP
X4AcuQdAEY8lPUV7aOfyH0QZuhRs7BRUKeeiWXUqL9IRc6PoP1r+gEjcM1z2BYndci/HzTplC2SR
zPfRMxAot5/tN03rLTScrzsejnDWCfGs8zhAXTTCnpEqBYloLgQT6sHHEz3s7ZiIlGgXpk+EDp1c
yoKKcSI6BMnbdi8Wqc/TUzXum4n+1XPqoc1ZwB7e8GbwMOhLvD08T7IAgQTJdttfFVrsPu+ipg1s
OIKzvW1tQfCm+YrEKvvVC0yYEgN3T/b5PpylAnz3kJ55X/E0a91qhnXYEp6FPq6nAe2lQH8KPkOv
xvYKlwTkbYwr/D8bA+YFKigTz9W4sx8iGhz8Zdrfd2otiq9KxLZgJRrZc5Nt8PPagrMbn0S+UoXs
jCVu6XCoXDEZ46AkNjTUktMtPdZ1vHDkKFK/uvc6fjpoSGFo+q9P6W0tyyKUjkyseUs8H3uHmjSA
PVMeWAYn7fH38L8VaSS0QExQcbmvoCSbG/r1GikAzraA5P+J/PjOxqu/ZM1Y97u4afr4EVjQEXuH
UEYD13dd+A0WScsFAbs5xiIG3A0J1oSe3S1+MVJxN58DvNo2CDf+14nToK/ft4hV6hzVT8XrAbR+
TzuhdHQZKR6fkAnQfluQZI38KSdjpR2TS9zfQ4o+L85HffW10tjocIWQdr13uTpK3uHiJxGvP0C5
YISio4/EWbVXtaCiiLvuiqLsmu6pkoVDtDLMNrANjSuBaGa4oAVeQDaL+A/org3NAUFa1tGjXIqN
IoA+Vm+Oc6OUQOHpGdOtFfqci1HcmpJYv+318aQUcSqnqRSMFGdrE8LJZgKBIVBUrikQ1c5X5Bi5
3DB+/ciV/1SOVvB1lsd/8tVb1Z3SMCJqOfbp0XBZNJOtsoFCJdMiFODVXaFnhJiSg8g/zn6Jmw9u
kCKKOKLIaBxFCVsrsgtYLpJWq7EGaWZEBcQpvyrtxLPqMIIrdWMqU6CMgXcp5Wh4RvhvdX/X2YaY
OiC3o8djgt2lWug5KYeC3TTqTVPflKxwtjhk70/11aoB3fPRp3iDho3/QJuL8L6WtsHmmqUCeRCC
zSeksJkhjBxoBrhdgChrKtK9GCWvHO/y6kh346iqY9hDcLF3oran9R3ZMPuRgM1MWWsr1/jpebHJ
6P0krEjSpV+DoSByW6WNvMfdwi8LjU+WBEZ9nNqm5V6eDEG8C9Q86zBfQrbKdHWs9GgJokr1jE9w
1XROuhuCVaqB6yqh7N8SBt9nMyOERE8ZLl50WiF4dylOS5AZvsmzoVc3BZnKaxBXwHX3OfZaxVyL
b0STSkVyoBXWoRDBdtg8IfYjNDgYw9lUulLL/DhzvfXAznu3wTDXXM4pnBSBUTs/+ih76r8FEaXq
iZR3dzMaJEDOcvIdYXXemfi+MnPBBPeoxYpnM45/A/fz6yfpqVGONB0W91wQrhW4gzngHLFgUexg
XG/cfCQtbAytX3rRhPQXeK3Mx6C54X35EZkIACBcsYJkulprZbYrQSB4iUz0N4PonoufJYMmpeZg
3UlmZc+789BjvtftTlPCfiwqPGF6qWcDf5O/b87no6aI9ZP0euIUSDeLsot3KICEqY87trg0eVfQ
8W14pbyllBY77mZ+0EJ2xgrj6pyEj4o/WqjTZBA8pMOxeEjCEqPdQk+hDP1HPEpatoUSDRLsilis
XHOEj6yNAWq6NFT79WmgZHj6Nt+LkHIyAIftovWvaoLvwkZjObenczBm7yL+5Htp1q6S8cThqdNS
hvzB0L+75pJrGVCS8BejZwbIuqe4K8QU/MWQtW7vVr5tYNxkIme0pP1EbQ+mT74i59UijuJBHAW4
9rCyntbqRMllnib6YQ8YvU/CA30vIC+DUwPynKNrD7yMYd6wjDg5t5pjhc1Gb2ivs/D6E/OxDqHh
Nl1h+QWebKEx5O85OmndKX3ibo/r6u+aVcDe7VauxY5RG90gTDHGMQCepld0ZORedUj1o2jEthUV
GJKTCkG/gI/nAlHeUUpIDaqkQW/Mt/1kJVH+u//nwlIXSnWdW+aYb7cbn7Sb8DEToRkzobGA9mYB
FjQ2j+ISq4kuA4ZYpgXzvoMOXnXG/eDM2nVLSbLn1R02dqSuMRgHoO78xnn2RjhYASY5ZaErZ/Ik
guuFciLiC4fatkqFRPjD4AOfIRW3g9o9n1uD4LN7zLDfHS/ERaVIUPr2PKjr65jN7q17TB3yUbzS
Zc+qOn2aiDEaWvoZxlryH7oPgWRnddMddaIssFnZyvmEdib7ypCWjFkVEdWLf7SRkjkKlLbguuL5
OU8bhnRTO/yR4VBF1JWuBzc6oONJ1cyag/3EPkPnvQsdugjIhDthvOeyQZg6GDPyxursSqMTI7qL
trUpzpPEQXA7BR0MWi4iw1XSmxoNu/ZlzXQV44W4a8KAlOzRum95qp1AM4gpOC/GfsuCJWwbdR2m
4WNdayD3NiXyGWexPFQK3jilM810DEmZOoWq2XgxukHRJsSB9Z4zzsv2Sk5O/tNDN9KFrJh3R8cA
t6/0nZgTbJz2yX//JZCNYHV4IbcyrGM1TrUg4RTlx33e77R/Kr9v2dGEsorgjo1fRJ2/WKm5a+xi
n/fmyXNyOkflG2ydYOb+hzf34vAyxJGUbOk0s3KQSZEGFgwwfdzFy/xs9YF51AoJZHxePIj8ZxcW
selrj3kXFMy+xVR36ouzVuMD9ILscCNzXiz5NqK6BY1nMq2fTgXaFbOdk7LYAUoDPP+SGYRvDrEb
1ImFX44Ue7zCuRxpzgpT5GAR7UYkAvqPMSywai2csTDUlp84kw6tZN37hQRZsVFddoEGnjLetBIL
FEy8B6AmjeBpFn9/5V8lXofiCyN8oLBdHZeDfRFbmyFRrVidAJ6JXwRd4fyuG/doDb1j4bGnsdbV
cRjfz/rYu9JXiRk+CHuatiS2GsUxMojcVb+NqOU/aSIdpc9ypeLvdfM8xsgYZmiO5hT4xEPhP5DI
UtjsHbQE2wMIyj6ZYCV9kI2jDxcPiJZgNiXhkFa1iHmvFmrw/xvhRrmisybyIGzj1GS7o6c8tiaM
YvGNlq8wQe+Ahk5qwJmUBOTFMoZMRP5Pz2H0T+A9v6igjW6OKBbuFUm48aFpbXkTAH0ZDI4uR+RH
Ad2fGlyETu6TeaxIBdnbbROfJMgCQJUGzMy7hrEivrrZCEXAOszfBIOUMaDN2eP4ecW3D3fpgyZd
nIg37pXwBaLvSiiwvkSD3tdB/rqBvX6mEDfOkuFraINcB6xiVYKoHSDhMZiYXnK/ky8hixgByZkw
Ey+ZS2Lp1R88b7N8k0k3DQk2kTJtx8VwtTqAtgU9wFKev5oVxq8wZjqi/awx8dPD/df1xSz9Y5Vd
44A21wzEMbfqVQxNzBfLu7TsW+nf2oo3w6pgNDkq/mGukJr7/q/1voMNa/wS+bTeiNVJDSlI6yDe
ptsA3meJX1/DnozhKrhLQaDyTiAh5Ei22vJY17DIwf0CROskl4yt62pKz+UF4J3GjctJGWQtIxLo
8LQnuhuXylsub/zts0hxwlk8bF9yWiq74tOhHx1AHawxGntHiGW7t4mt3oQJpKD4duiMUiIoxHBv
UPetNJL4kDAITzADwSJqgm8MQ8YCj+Zq6rI8XJ1V4HkBafxGbtSYuX1WXqN6AVRoMUh2YgiwdvSK
gHWRKw8Gxxz1SnaNg7I5NXfeZAo8Wb7MHdWpMIGnJJy1nAFDiIw6WrqfsJSvqEQZn3cBmfXnKzqK
ID9HpH3BYkdNiWrIIysM8xsH+r+TYcKBVWt9oO7sW2ZUdK2J0ZZXK8pSdtLrKTka8pvapElB25Yc
WODLY3ACHv8wWaZuSzYYmleU6EUTAzPYR2b1uZPezJTept8cZlHeZksTvDsfRC8QWGqTmowKIOBu
WyIGZClEqzzCcPb0KKRolHd3yHSkdSSuj2ZrXR8dX+lXRyrj4Rt/raCpihXQF41wIg4tygznaOE+
UGfTdi3+iSHLc9td1ID/LkA6UyqPo2TSqj8NgAcHGNGqbgllQajXegBebCnnFxqPZ8RFH8BYtZUP
1IEZ0ttn5WsCZmkaZmPz0K8Be+xMvbmGGUa0OLWVMey4zoGwclmvlK1RbIhLTgXF+jYb3ya497v9
9kmDYrBrdDH75gv6lsdrRYourfZUPZkW4V0PjdbSab4r8fQKei2KK6lf2VPCn8vFSLCfcN8T4mqV
Rp31N1Wvmu/B7geYrx5vKo+FX3JQA9xC0ghW3wAi7eSWvJFO1CO+Cwwx7rDtEl05GUueluycAcsW
LJzng/hojmAMICKLgvhJq+Q7tty5XwzMbpK+RkKIjLxGiwLKqeMyiKTbE9mwTcjgNGGO8Z6dOOiT
+Awz6IMkeLUWVNQnunw2TCIfna4HvvvhabdRmCnu9etzdnrukXUdMDU9XIpq4KQRQYBI+dR/cRph
8C8AUu8Ft26yhQS6dIzQJXJmMFadgs3pUBzreHOjLUtfTcAvU3R+Por+8R5+Mb9qSYFSzxQlRtrX
j2XtiOedxklCcU7712qtA1+I4RpEJns1emvnfebDZ/br/nMXRPbacaTFx/h0CM5sNM2NtAf4N7O8
KmBIJlsfbn1Ez2m5aTG71zNeZG9iKq79SmkVlt8P2etwGEdQ4i4C+6m99aLcIQQZ5GmQW1k0nPgj
N0bjpt/VH4OXFO2pSBTZMchsYM8KC44pUYVDEZK9pY7L1dqDYdLJ0QDZ9ao4oM8Aicv6JTcF0xvi
E59jLRmtDMrAdoKIot0m+98O9pVRepMeSjUfxEwlxW3SdB10qfLPlc+HhfzO8gzR2c+479GuZ82A
Afx2H9E/J8W6Xye5UYT0nQCj9+DvvmOs+1iiLkTMVSMOKYCsFTkZnOL9MspuxPO3TldLAdaiclCK
yHMjAioG7J5wCEoeFzmigMly0k7YR3n1ZUfbvcxuzUADttr57RAF7o5ZfvBH2Ap6OkAKHuT6W94t
9eR6HIcasjMbcD/vhOMOsHWYDBxk3lhxGiBtIgKh7XPCh9lidcmjLxO5GVQkXunDCMkz/2yiqkqB
TWNeP4hctTsnaZW+G7PKoUh3rb3My//tur5oUYf5VTxSjC2UAy/XCTInmddyFO+NKdIM/lDZDxPx
T31fIpsKf7fpiqUG81WN0yqzL7DQH3gLN/BO7nmq4qMw63zgKpAiGdC07ybPwJmXfkaImkIcVmk8
yqG/9v08Y7Ku1sZcdXxc/0GvgM8IfM+QtHIOh1BS/uiOBrlOoxIB8umFeFxlQENENLwQ4cVLRuHg
OJhKRV/69hhpB1zhxbaSF7mASL8jhCco9r3/NWakG3bvdhwSzs0o8mLEI6DE4Zcctmd3P+8uSy0g
QdkJsbn3X27ke5ZV6biLFUnmUY7F74KzlhoMhV0CzYNKsD5NTYEZPq4ffUhhnHY8538cToCnSKaQ
VOBT6AIFlkXZLZ6ygIDMyITgazCEvphH8ULm/3XZBpPDuM0HXqjO/AzQ+cZ0Zy2uekIYy+1KlrRq
2Tckh92yUd1Lf5/WrPwNerUoEty5HHtY+oqiO54CMTm2nrHn+jIunZnt6SmVYxZhaZyhl8kA5K32
mw2X35AzydDYjpQ367cD/d9BeZsEb2/ftLPFLD0MtpAvlUlyDZPED5najij2EUmiOfAUXc6GRdF9
k7OdQRV3ahRnJaoDt+s9LHzJmF5SFLiUtkEXCdSMDU9HHyvsv3L97jelP6CzRQnZr7TJ+AtL1rCj
olWJ7bLmLNi0KsdZOqVOeZNxuemnesY1NROGoOKbYuWNiAP3wEEcec2mN3IdwF/iYlgi3KTE6Ar7
lAETvkr22pu9TKlpx82f8QfD+pdMWOP+0eHPt31ZuVplyGkzKmBWYHSVXDsmDB5TENLx4M7YINUA
Kc9eA5S2oWYxHjAc3AGrhxzVP7ZWdsemD5XFfOQhCPlwDDnZtV+dI15VHl7MbD8DrYhFjBJm6B92
qocruayio9bKLh6/LbVZTfNoWaf71ueBAKlp9ZfWINKSfWK4jKkFewSJZLZmhLmpz0fAwS9WtJDw
OvyW/2SI+2jCoVboiTS4+lgNn4aCndbNJowDNIdOp8axZGvSMUwk5H2iVBbA/0DGcEeMCjL8BDFO
axgt8R4FO08/izv0Vo8K4eLw5LnCTFRbnreG+Mjb+/1calZ5hzfKHoTgYFEIDEHjZcCgzrNwHhcD
I/7mwDQYU6oI76+G6ZIp6KbqV9fQPQvL7NnVI6bZuGZ62hlw6EyYNV1ZYNYg/FcA+lhP7Wrtb/K8
2JMjXzE53gRp8S7D4FTXTC39wBvJObufYI2cIimKf/H2LA+RDmgKENTrvm//+uQ3s4fRu59Ithrm
VriKoU8r0QU6xO/zj6FQWrKVGOox1lfx1bC6Aak13q/DkJatbWafah9F7PSFIVaG5ouKEzQNg1Mi
eEaylJmO0eyMogyhJC3Gl9TkCkH3GEoh/OoL4X4qR85kccsaSDhVsW0fSKNwKPVDgF8b1SO6otG+
0abac7wJRbDpDoYObatbl/r4e514PVLyKYpQ0iP2QNqaf9gcKuydyj6aNffW1REeKnezh77KMHTN
NnAoR3HjDyrdFyFnWM4uXc27woLgjxWt5j/l/9fNUbuJhScnQF0jwgO3t8NYZujjLqGY/JDrXzs/
BN1SlAL3X2W3B/ZHTl410/BHDH/fU+wqUuuKxd39Lih0g971TE5VKrUEu8fEACmeLPK84Dfb1knf
w5rrmdR5M4aLKC+iMh80Mkb25JNgS4NF3vxVq0/EKsOZ7Ak/BGiAJwZ8YaChGf+fN4TLS+OD8HxW
A59AN83oTTbJJdGFDzeiXQDwdZUg4d11m4aobBENJ9soFJV50Va8dHDPM2mQIpy+yXJitenrpUlP
IYYP4JiVPs7eY7vfeR8r79c9kwA6wBHoZqSjvnWGYVTqizSJ25kkDYjxItbELB3ZiRhQ4ihpkZxa
+e3J6ozW1c2eG8QnVtVEaFH2HBZv86s/gT4riqlKDIUoLkgSCbFiGnanTw2SPLmzT838pwXcVgYX
m3Suf6l6udtYugFKJRxtYO4CuIB6QwcBzMSLFfL+WGvQvm1EpalK4JR5WVyY6jmXO/PfI0pEWvQC
UNUQJkonIKIrRnmd9ADBzt3xB7lv9p2AAwZJQ7g0mHcDquXEmsgxQqLPIG4QXVFtCB1tP34LwP3W
R/UTrVdcvug/pBMBjUt61DgHeJ5FnunrzHY0Pqm2B+gEBMTAjoovYQkiJlyAWXYjYugzTZzC5yV4
NWYl/ji0cH9DySX1s6lmSV7n06L0dXTPqCtA1btEnvZBA5ujQ4sdSZycvqzlsixXPLtq8RfMCsfV
5LRFBwVO6GeIS7dN5cPYkz313ZHCRjrFxdLhBugjl6KGwxC36rxdhRUqBODdwXxAHfgjysGB3C+f
CSM3VYClJhVf3gck0y36M63Dw+wWBYyuq2kY6cq0WwWYSgmsvjdlJ+DPm776r5Otumfy7B2ePY1B
BRJ8js7nkyObdv2apJeRKbPqpKjxdhB9X8V6huTMEuXa4pBlVe8CzAZHFppagbOIm0LY/g7gdoe/
RqvGgP3bJhgA0CtTIQwUbtjuCcUo9T4Poom6lDVvE8Zk0n53ifF/90PHS2JT+mVpbff3/5UlVXZ6
gMb3QSm+i270drwXSq/FiOXC+u6vytreHt6wNobCvQVTF8ryviAE7FxS55BMgL07Ibm7JJ8u41Pm
2K/SJ6Ttd/W97kMpGBv/ZM3vpR3wisigXjBpbve7CTqmnKOT90N65E265El2xrvnMz7WUjozPNdi
QpI6gXepfHiFgN5FbW7jvtb1qKPbPhwxHDquDh2vho/MBAY3N4JuichUQjK+pLEnWJG2PVx3UDcm
BOciHWJxl2sYQr7jlTf3eu/GIHTY+smnxEhsxnaD7qrHOOx+FTIUorvhYWvcoNvzlAE8OPbRwcgH
y+T8QtbgUZs+px1w5XRwCJ2ZsfsTxcomXVddWQBaiA3L2J0l/7LLj4/RFadAborSOlMwa4VbLWnN
z6rHy3SXU+uR1XOGohtWgq8wfQaFE3xJaFwPt1mv6Um0eH6fcMTKftASrce9LZa3XqkxrWt9dO23
Lid3ZLzHlJOz5B//Ns4aBgjPIIJ6Wob8E87b8x1YpNZW4iwzBwnpCs3RU49vJZu5EO37dX4IHH1I
AmA7i1o8cJtxZvAFeBibVWgt/Lc/gxiC40Hr/BnofdeCUUNA99iEgSICkZ7X6bnz0jBIBLXFTe/8
C4jOtHAl662eLXHdOWpYkZcKYycrtwsE+a2TLSNAiXQFihQl4FLlr2u4zJy1HFf3dRIxAnNes7qy
2GmEZuJ0BToNtlaVtD59VOY40RBemgt/+xj2dTwQWb7s6H85ceVTADxJ5uZoYkWjeffhdYD3jxR4
j3W0C47xKpgevRhgWCFXCLCigreyXv0uVmXJ49KELPma5M3nl7JY9lkTHxl/J+KJUdmCNqgSq/UO
eFJLrotuOSS2FcZV59FsztugZ7ASEJB4861Eu8qggvxcfcwA7o6dsXpL5+9vqqjeGl2d1SyztXRZ
NMY+nNsLf96NhakRd4/HUgA1moHvdgsoFKVy9uPT8jlsTjR4MUrIEb2mDiHImXdK9Pk1CPZob9hh
Y5ZZv0d4XrUDQql+u/mgLqoWmfnKCHXg+GR/wHGBxINp+RDvYI1NtDPSq/FDqJY1vsGqWjeIPdrj
tbbR9dDLFeSSfytt4iE+3t1zfuhE/WlHl1d6pYi2XvbkiCFxuFrpbELCkVx/eocHf1e8Ed+Mk01H
yfI03nMhBqeoKb4YoXqDpvFmLwfXVo16yuuVShnBszNN60DhWwkO0CyG4pM32NYtY90RBiIESqog
jH2ms8CrH0I0DanogLzU0c13Esvjg8uOM1lVX37M+JTNUs/WmegoZ5TrNeIErOXaxaJydtfzWCoR
joe9K6awlR4nqM1tBmOhGbCiiVw5DuZkN5zqxCKjnqqlPwkRGQ0u3MnNIPLPrG9M5Lt8zXyV8Wsa
cJv/Jmwkvl8Djt7j4RxmtaTWWZG09HwT784/Kczp0+yJcs3H+a02TJ7vv3JP7JQAC3c2rL4fWPxz
9+AQ5zGjFOiBr4TLSHqzpsuMAxP8LsKuM4LDbt+eRLgCg7cYW+SIgyY/lNr8v7MMrDNYsffP0EmQ
e6RBW9mjJOzg/cgpM/9u6PgRKErSEXC7soyX1QIXo9Pw0KQBN9RPZalEPJSvm0nAh4wIrj/5hhYh
12m0XUJLw+ORGU0OTTgSpp89JhDxVsAy7TrY3ulJ50kSZOkj5RlYWJSY+M8IHN8O4vctVg9D16QI
4JFWumBOJvxSyzJhPGVkSKzT6dPhA6TwnPuK+J7FVZs7JRfuohzs6g3Xqd8Gy+M4C/qsUFpC9Uuz
bNx7efCcqm4HDV0OoVKhyW+bON68wFRtN1S95FeAW/AteRsCzigFABpYAhF1sxs8iSlGC++9UgmB
mca5NSQC2P0j8B207ZVjFOUw4kCJuTFtlyevOICZUDzuO5gjVd7CIf95hxWuvtOEhJFXw2IB93cT
1YFrk9XcZ5AAOkTcSHSKNkXNw6tpL+tQP9KKRN4yuj4oZc4JfSlIaoQWtf3HxbEXnF5Qclm0oAew
BMR1w/+w5T+O08jQAQ06wZdVbV2W9TM0ffmQpV9kBWE0pfWcziDt1IXkUiF6ysJOU6PQGZ3LHiKG
tU0mLW8JPkR5OfbXGLjDlfRUyqfMlt6w6VGfaZMaSFv5jasAxBfm/EX7nSHRFxRyltQWXiQY0lOo
hhtrSmW+DdmY3itbLQHvDW6NQ9lPQFYYsIbyyVOETColBhqj7H5yJll/O/vohgGR/dxAr2A7V/QZ
Dk/pVlc3rMnX+wtvoC/uYygb4sN6ENTnBHabT1E1/Pzi8B2uQlf/EIYDgtCUEmeu3VN91zt3bQhq
nxZkRqZHhE0Ytk8gK4n4qwQlJ6isC4WSFVrj2nV4V0eohLwgnFWLUHI2il27xghLM+BCUvA+Bt2K
atyJoethUXSsEC2aN2wubwGyWplYBuHGidtGaP0tImDbhO3XAxEXT3BIhfuUJ9mIFFWsL9EH0hz7
F7/FSFiFiqHHbMG/oZX7l8YkaROgaBZ2Mz+pZNZwsZg8BFEpC0dS1/Crmpr6u6KvC16xPbRFgH9u
vvAu0cqD6KjoqDx++vG9Vp8YyHu3kViOyL+5aMAiTZEpXrL5QdnZFdVvv7rxSQ3LXP8QM2TTWsuz
dJIDnlWBHXwBhAly85pDO2hHfUWqhbsgApgd7yesDzN6+eSdsHkFKDPisgCva+VsZBO25HrWFQL/
MNxhyLPVnoOExBPT5v/EJAlDIC28gvtl1x5BLx15q05BqkmzYBsd27ilS9FOXSWW/SwBUJw9VX9j
Bxzafw5KJJr9mZlQ9ShCVrD2LChsfBWB455n3pRqfLf6CHe8pgmKr85M9xlCGrhJrLKzWU142FQx
lF0/CywI1a3K8AtKpTAkWReJIjqXDpfo3PaKKUqh8/ow1WFARDFR3PIHa/deW0M4l2+1vW+Bxmz8
U3GZM/DYzOI0U747oCujyD4WJtNosFNGlP2AzLWu21jtR+XfwQtDTEIobfWcqqPGx1uop4HaOZ4h
1gOsAb4Xky/dFzr+tTHoEq65Y6XeO/6YFp+yvW+SiVqFQwemqIYcwWF1PfRIPRhBvQDD4qhHgkyP
xPSxMTVVQ83fE+sl9NABH1aPICddwjYkwbIFQCabYFeXNgFf+HGO14N6hsuTQHMwchObM1oG1Equ
bF1cvBiH/lPCg5TQH4oofvcVfIb78AB6E1qZuOsvrHEchUMhxvtpJDRfNqjuSfAv0g+q/nXv5JmO
jODQ8gLhYLoHChPMMGo4+6i63SABkWd4XJ+EPRLOzNQPF/jQNnS8pHsJdt45Q8T65tv6i1Md84Im
dP7JMXzcWEkVUMLoqCSDJh6eO36QTN1Fuxz6FDRgLSm5Bse+xwx9n5ZBWAY9OQ5/GCoPHs1VmN7G
Ramzb1kL5P+qpUXNvEUocWuw+OGY6HuuOxBT8lsuA46RWSeIOyjTcDfNJ7lSM9rKqpwP9vMPrcnn
oGdKD23XuUqBxT9e67f+bu1ObYBYRgx1AqbVR//iC1xmJlPVYeGjJCI/DSAxWx+xY0ApVuks1o6K
GuScfpm5W3qyKjG2DxVmKrcNstbjsQKaULJHIapgionB3y3Gaw7nBLTb4EZDXLnf0q1n+FrrZV6U
MT+aN43MzzoI+EDcwQR6IPd/1ZMVGYwRAFnbBz7YZvJZxfzR8rSMbGVTakXUvAYVSMTQRe/931Wi
OvD+vRHxZb8xwXxCskS6hIn9sFAlgIsXwl37NMhQE3dF4+rc/2Yv2nhsqnkA6O/8COC0sPJw2YTC
8TPuDU9prqwL4+50Kw5iZzsCScWmNnO36v7oXyoOcyFyJ72fv0JLf+0hoxcWuvqMj+neNc/vEPA4
gMU0XHN1rUxwO2EDT9nmO6/0mSmgxbZYDzeFGRibGrSzy5u7aWvqleB7fUIFfnk1c8yR9Q50k6pD
1UkrY0uGVtd/J9nhypZusJSxuv3mFrQGSB3/e5kLDvmoN0K4eAlXS/4lNwv0Yx9lZDBrg46szTJq
3mzsRy64L9gB8jkQ4ZuI4MYQUVzPL5Dh3Vqb5jg20QlijoOx8yI9XO2Djy69fw2YmNk7bhBFc+JB
LDfKaCzMU5z00It9jsN6IUlEc8HVAygDABIYt+xmTQCGwqVtnX6n2zl6GDyxKC3N4hRCtKMlkgNE
QobA23ec5EVWs65hmPhWRZ4YJYm2qRc0wscnRr9MN2CcTTRpcHoh4cXo8dpl6og6ML0D/AsXEkdV
T5G6RkAz17rEiMvm65db30lVb6lKenHwFGlm/3ns9ETZIraQlAH0XGflROWu2n7zww5iaI2NbCzd
3i3L0EPyXsUhrlJy49UU0forPq6d09KlsBmS8Dkpab5MRVXn/z9B3HF4D65GJ2JJ1S/4JoJeodun
Ni//wza1zfRv1+1af45bYvOOFbC8SOjodAdyDG94N3WL7oyZzylwgTKbCoo0wQDr9BX46FRsiWpJ
AU3m/q0O3DOJNzPtTvDUVP9loJlQTPGPyL0ODdkufcDLH7/y5vgZWE32P1tX2JSnFjdbrWalIsX5
O0tSbPH0QLxedE60QPWCAcFlrYzvsTKwfPZjNXs2b8FGLpzUO5UE/sraZzRU3JNKluo3HA0VfXmA
qD4O9afvwMhuY3WkJKEuL/EMXPjCENju7rhXam11YE6ecU2BeoUUNsO4MY0Z1nSQlCzvb+IK3EKz
eNV2S2tOwgri1gNL1dlZ0g6+KZwr4qTF9pz37JZjctoAhPPayIKHFp6edAf53c+jHDD3TCAKEG6/
Rx5ZFXVWCEamxnapHHQEr5t2Gl4S0JmEGQLI1tC+vy2xDDIekkAhVTlaoqEFOx0XY4R8ycIPvfdk
y7F8r0yXStWd+7Wv99p1Q8dwJpVFuOqo0Fddp8CDMAxevu/eUTmZ2SJO6fooYRUTuxiYWKmVG+K+
/ku0lPERkSBVHQLYBIAtkbbJUAZR/4N52ZKcKI/Hcf2xyeychBKsmiIdnfnx77QrQPfXVgUbm+JR
20SpbtWaXZF2bXAB7V+8LVNzaSagTgak4DxFRQmNoRaREzeFJt5UCTyW6l7/MPtzUUBIArlA9QjI
yCaKJCGFpR46FMxfmEFadiMh+BRmpiRjtPKv4Eb3KTYUVCDwbh3FrlWfaR9tm/2MnAtRkVg2YFB8
v52OGtvYDMY8yunqvhI6w9HSHjIME4FYzg0FlYqJmmfP9wiohyNOs1syBXCHigUFw40/Pdg/KyrT
hMZrOgYs+VIASGBTXpRcf7zLHRvpBxsylXhwMYv7Ja7uJojMM//AxSiI7SvGPjp5PKEInnEeRDe2
4aCdbTsDnliv3fBJWGEpro3qm6Q3eJTn0e8WRmNOtFAFndPbkx/9Rh0HWc6Zec7+bh6Vj0JeFK6u
/bIcAen2TIJquqx4fnq2RVc73bZA1ZHrkYWVoo5oXC3snsfNUj/YLH5QI59/Ywraw4TBe2xIuhDM
wFnT43h9/whRxb6p+hSES5X7/IWezRvkO2Fb4wgprQRrxmU27Pf+GXXC2qHCU5s5JOP47P68c80L
UN155XYuiUWRkjt4EaOTqRRhiXfdMrhGSuPbDny0acpUB89HXEpEBW+THNDjtn4dBu8rPYgaIFK1
cNMbD57maojtvBoBrf/OdVEu+GscIUY4JI66jycJvO5elsxBpkBS9+k2wvt5DRGR79y4XAd/VEp0
WQHkLTboK6qypyf2imGL+3HmZ3KWAS4YGTXOcS7IwS6hfeSuqZ/yn4sPuTX6S90C4C9RjsYXehA+
oItox+BA0tT8IwrNECJTgDpSUIpR0Bg3Ta8P4AbJMUgWX51rZRwIGFGjKJeIwVnhOxY8uOLui2AU
NmJTQ31PMkaWVRLDKach4FKZyIEx1NHj1rvlvAlcZv3wYdsMs2bbOI90SYpcemnbjpja4JtUjCBW
DvjCc1p1q/qJ6GFK6a6M0aQF97OKZYuOkPnl0oaLXWcr33Omih9k2nyiBKuTfQFtx7bxwih/Mj1d
PaujtDcAwJEuq20WAU88pkAPGe9h43smqFr3uGN24v+EUOJxnwzEtcSRV4jYCNsAUAu+OOlaDJ8M
xUtz8db+OqtYPb4Xw0cCFfHZN5ZlA9+NGUWmIfL4AVuBMRRNhpeRmhrLrKZib2sKPJB6fDem1In6
o8vsQ4tTC4UBdauw+JNULgSwehAblGkcipfWeYiwIVx0lhVnGaZG6LvN9g4mrCUCCPPJ4v8jyfHq
XXyBifowcZhdC3yKMcgnUv3u7mPajmfdeJRAj9ao3kNqAzjJlXE/QbdlmejtwLcDgconpab4FQwZ
686kW/7PdzBhIMvpDSmsd4imOq/31jYs4umZywCEpQ9ReRgdRIaMp92oPLCzpzpY5CruNf6vbNnZ
zBdO1DPvNFc+/AHXL3bq5fNN7xnGwIheJLarjPp4Fam186fOBr83+u0LpVesH7w6VN/nkAVsSEwH
cfyp6aSof8b/2DVyMAX34rBqOlWvaMKTqFyniTTtUVbud6HdVU7mJoGHEvBpeJEJsUNFqyDS8kK1
j8e/pBT1fr/184f//A/9kL0RcGPvMKS4+Hx+8bL79qIVfihW6vOsnn/lvKHWTpAeKLOyQgtLYH1c
flwc82uzxK9ocVT23y0RN+jlw/IkudxSgTWIXNjjs1+Z2TMhSD8JyCwudqGxTQNgiswm23KiX+VC
9tHAGpKn9bpujA9e/wkNxZpljXDwpTwk18tbX5ROLEtJtOB22et/GQy2nhYTPzcTwBKjp5nD4STN
yv1z7SD8nuwewjFw/G1LXckzkW6Cd/t9/19HoD06EsPUH6T6jqV1geNZawvKfDOZ9XNHJiH5iQjY
6kau6+3E23ww5c8z5ss/ZriGpUCWHIIR30aNDi6YrpGuJequ9/sPdYUhbDD9osdTtDHyWtf6R/ky
McM7WRnxfdhTyZUHBzhDy1TKvrXHNgF3BV3v6E2Tezc8H20wLYfEZemwdN0IcW5FgnTsnnoeDLlI
pBORUkqvSuKY+AqQnHojforG71C9KeKL9ABFrwUTv0ZhnVyRs1hIXl/SJfbdyP8c+ZyemJqS+fe9
N+mPVnos1ZquCSbnb4ailo6IzZRC3XCEc3NVR9dA28ue/HPAgFj3iNA2nJqUlrDp3aRzuyAKhb4/
sSYmBhDXoYFK7wQ+273XssXn8AQrS3yixtIQSaOCDqrpI5DtU/ms1vHfpv7ixjy9v4KxH3oOUHvW
puYqL1CZktNue5TPaUXBq6T6Ad5JHmADP4WKEuXc3M3I8roejgtj9gXnwb6tLxpIZnv/ug5Km4GQ
DElBPYdpxgWigIBnXO7lX/KQKQIu6XvWso83C7kaE10Y+Zctf0HQMY93bSVZuZAsIanz3M4dUkyh
iuvUU0VSyAAhabUwZeaV6yLKASGQgcgqQLhikGB2EqP8ZCSfHCSxSZ4+NOJ20kEjckmrz6nDXlqV
VmCKjlBDcjkuq2R3u0w8KrVo/CR+OX91DZnN3CRXfqHXhJutimjsk4+8GQdjaKRv84Tx2vBEXUrW
0fN+YV3nSY5mOqVMNqDhRS6dClfeswWHOFAzZtMbnelfMONifTZfBJwwyMpJeMnlYrsilKWcGgEd
2MrZKcmBnB3A7manGvVhzYXnDYEvPHOmA2h1+vVlmHbbWerLF9W1/KZMzYwbvbMyjVdNTthsMpct
01PWhqE/eXqRdZYIftdx7R23eup6jEu6PetEqsMa2Koeeh/U8gIzjvgOdKxuzYgAO9dkjmNNfqi7
RY83opzrCw4nFpQqaqkMsxiaPZzRnY7rWB+eNsmKpyadPHy/5e9NIb1oLFmPDTHJFRKnf6HQ1g4C
07JoshBWlH5lwescJd7aOO8y+3QXoT0KwJbOi1MR27y7ZkWfELlu7ERQY7xMcnD5a499GefCbijm
JoVt14LoiR6ANQZtTZiWk6lZfOATn+DILmtH+XY7Wqg+b3/q2UqtuA0RnYHloxbEqnyRka2x6Hes
pWxRhJ3Fl8TIB4bHEPQo6R7cHxNu+LGMCI9ZOfVS6ZwxZS95ZO7cjd6S6ia+S1YYdlCkn1bwlwku
7vDaYj2OzojF6OkMwnrMYAlGHaB4qXkbsu16X7CDC2qHR34C5LEZlKAhha3zMqvDykhLJOFu/rp6
QtX/6UuG4hPxC2dGLu8dH9k5R6u+Of7kkyYe91LascC0DN0DxvLA44FhTTXJKcYPbdudri7xX1e8
Je5J+Q2EOPXA255AEpGQjFCj6iRXrSRYGKPm4SxAOHOFzLqlAUz7VNfxY+PwoKpqQRS0C6S7QUAO
I0XfHx+qRHj4c6130Q9qvXlYejT5+7Ky7G7wFJUxl7izcv04wpuKhS1kRLSRG1fdYFlpFal71SvB
o9n8ZEZJNCoz966yTZb5kiuB8OyN22R3RezcOiGPk5Lno9mS07sD2ZMNcMjQQgjsbAWMMr8u5wSB
0jwsv3o2tPqGAMAQX7c1M3pcAA02mfNwkoil8sQ+n5PAEYqQLPV3bSqDKHwhWAiIxaJoWZLyL1+6
XO4xbzCuH9f+tDGIgR37L3Lu420kLLvALlQZfpDvpaeSXTAkG34giHlkujgju0OP7hZUvdzKVKzX
r8Q2C1PUtqGIWQoWBZ6bkrhAwtJEwsTQ8fTVuq+L99FMf0H+nANWQpdSDXH+vQVvTKqXIdv0QyoS
u5p6HQbDlB9Kg95MP1TFnYNgLKyXK8T3ilNv+jNKWBo9k9brmGzV608drPLnHc1qQPI2Dptx1pML
XQUAm2a5O4yp+tSTrh7FOsr1aLK89LiWS7sNxFWl4m51v8n/Y60yFJnXiSFCi3SVUoToapp3TzZa
0T38dD8yPUXrOf5io/Tj3KM7iKDUoop08MlNUGFWE5UfpIZMkzIuf44DTNaxn4IDHNIyV+RyQHjO
C22BtAD3Fbp8CnwxLK/uo+WKr/hgnI/fyge5wrKUlCUgOGs944OMBVfkmezz1A/FBO+dy+/N25nm
GXm8CQs0NWgyUOCgSJ5QfA8FRWp0kLPZ/vAnADBsSYE3pb3YIfFTRf4nKCk7YweduxmDD8QP905m
ZLkk4R48olXVk92lq03tRGO387mXU7di+THeO7IMLuv2kmWeP+8eoDVj7Mqeru2jHu092CVs0+xs
ofsNTyR74IAA8q7AOZws75XCwCt0ip2QxqpfVzTPoa+vKucdh7MfC8HwCOc9qYGSuuoT9EhhHAzJ
kR2uUF7WnrPEV7ZfmvzTa+7NBk4CZDQU7yf8mbFRe3MZEjkGnvEnTecqcgz47a5OR7AG7adKc4lf
r9DRhirEWxhYbF7rSU+r+L847DttmX4sig6owRRgSNPnw+ZkdP2k+z+vILa+oVotkq8feV14+Ssd
p1RwZUatDoZ6cVC/IwBZofme25lCzJG/6+b4byTOWDFn30Lvmke7q2j6avRIs0n2tBZDhNGXGvR6
V2ZWipdJS7JS/PdRvYAKcqRRzUWWnbye2NKgMrwkwImtrNHfAKJl1qeRwKKIQDiIuFOZHix4HEOf
/R95rHncPXa/FUqEWAsoCmFrvpMwRRNbWhwKRBGouswqWeOE4QIk8EWzSTGnDCnRmMFiaMaiSpsT
MmqnKoMFo1E16Q6UL58DCJSUqcSBSjbw9J+rFW8V8wsIvB395xLuB9njStn8xvFweNm5DA8bto8d
Q6QP5Ts5BzX966+xmMWhiKGCJoBfoRt1g8fD5pewODcQAexjZVEx5etBA2z9t4YZhRfJi83qfS/9
6bhYt8GNnHqVcpuCPZo0yiPTFfiurycDRUgZkVEbVd+hHLdpjvxZz/LmQogTvb7vNSzsM5HKCJ4/
oPlSMxRjBJXTofsYwM7GyrjB+n+YcqsHySuBBCGnrA2o2nJ50rnBr+ZZjm2Xt4veTR31iKp1Po/W
KyaBW/XwSaUxeCjiaEOGOLaqYJQ1U/aqdKAzEQOaH0ErMexm9Wnsd6Okl91C3zBvhfpy9VVmDou2
D1kFnCx3Jx7iBRteOGvzfgM2QVaPDnBPbtugdPo+pP9o5XoditsFlCH45seZlT6zMVhiEBs1BdFB
ODqoWlJJB/J70IxazxMlE6WdGuwOiPcr99knY5lez+i71JlUR5J6qz/vylfkjEJEABTiMQ3OP7wX
CpN2Q7JNLUSvrvGuYMky6heWGbIhq3K5Ub2ZJKfTWxeB3y9PU5+6P4Nm0zsEqd+YvdlO2TzucANk
iZttw3JqK910hsHsloC2IPc/lZY1Qqh4eyh7Wq+BDgj/REcZwY5RtR9aigdRLZq0Z+/9x+JbE1io
dwnkgdbROtMHLKdVxH/TSM+QMjpSCoAhLMAynUZGe7GmvBbKeU4ug9ya6Cx1LScMyQ392RX5nLAR
ClyFkv1P+htUG1Ox1hSzIGfhTpfSLYEnFXEC45rMWFdCk7gUvQQ7gp5zdNrBdsL6caQVfA6ldgZ0
KoYjoVI8oGlQW1wWQI9vhNs8VCanMAc+PYdfhY231z8xsMLE2vmSg3aAKqVsyknHOZqAxzPlMi+o
TygPVOJfOoLSeK0EHsXqb1ltev5yvd0Kq85IXVapjZHYZ38InlVkRZR4UoKg1zcmB1z63iDtiFed
+pgN7+4MTkH1u7ktTfPzQHp7xtWh+dLcb5gyMvCZPZQlwt886ISglSv1fYeQYWdoMNeGHrhwij7h
bun1c4q6s66CSMHOOA66nc0Vd//0hr2bW09gFm31wzBUgCOlrfM4it64SNiXXdU7t+727pid03WH
LVYxcCwV0IJ9U3mYlQ7sPkaBdQKvRZPJ5Rgo4I15NX/Zqoa4eQ3Nk8Tf+PhNNhV3+iZgWnWCC2tg
wy0Og+WWmSbYjC0+RvM8ZOye2GhaqBQeuq/8uvf9eRLbWoSIn0jMCdomzGTAuakaIXRjnBhGCZnl
1WcEceNNiSG15Q4q1eqMSg21I6r4S+KK1oTeC8O/iDA4uPJls3ylHBB1hybXy6AqgcaTxyXJq0kG
bBPI1KQ4sL+kN/1PuhSWbOGkUThOfpFdEPITWFDcokYNisx+vSERMBEnBukkc/yjSg0Wi/F4ooLV
qQWyvl6YS1OC7A6vyrc2gyh5hRak24ZtUme3elx8ZIixMb6eD+OUjBAC4zdz57IPGc6t3gPgyCHI
i0zYIMRpKBJapSFicVQv01V9MU7GNgKLPS4nAiqfEQeBdoRPm/W+i6gQ63Qqt2HRWML0sO6QkUrR
WPJDtxLs5QAYsdkCjKffYIsh7+etl7wCfiU8eopuH4egPpTbBfW6m5hnbC+6R191/eTTaNobTA7a
oyt5MmzxuzqC36ermV4xc+5rCASPtUv4Nx2vMa2YThuwzfn7OYClmiGhlmVm7/gN1vovYNBvxAKi
Tz1cz+/I+Z32bP9Dun3CQ1A5wvqwMyDHvaeIB3sGeAm8DbkNkZveXFlBGARUYKf8ozmuOvNSK820
+cBX6/xf79ZPihosFPWyfC8bM+ZtiIPsGcFfa38EaKmE4tsCxHJttl2MoIkssA1oPiMBJc0yd/Mg
Oiwd5yHipOFJan/q7Tv5DSy3nUtO5Mw9AMeoK9D+Sq2tgfhEiX8DW2EmS7OMCpCKWWCdxt8ekZKz
p3MPommwE+9wI2isqOb9UhjsUdl0boedbz7PBV7TT1j07FOFfTlgkVxH/blFlnjaZ+MAgCxGsFVd
yeKEj20oko06y0agcWpvgZXTyDwg5oMukg2rRYeP2WBoUdwTcePHEke3Wl1Fsqx2Ea+dEk0MeKQt
BiXsdcHJYZcZZREocsqTpsOL4PFm2v/OstWdz16S6ChIonp/dOZt1uwvHjzqvo8cFPQ+HxdzTKi0
a4YTfvU5RohZCiSG/GukVwXRa9kW8lBd0ovJ4iFuMnUAOBGQRCvfZDl5Uxmvd/n8fyOX/TSy9aGn
Zfklh6hex27ShjsZq8cJfa6YK61BL4evPAA0KNIiK9wMj772i8Xqzk2+gQ/bSvDDl9OOFCI5Eeet
Bs/waNw209XeO2QCmJysBlpkKZGfYCEgQwnvSiC7/5muUKWehwap8cQOwaNYp+TnaxyGC8+VmJ8c
5uyRRmJL37xx70jxESF5WPFAQonNR8Dgj6EdUu3tq8mboUJJiqjny8TwIZ9O5Z3j5ZQ0poMI5YXn
IpSYCmrbQCF63SVqLHcXB04K5Kt2zuH0RJ0KtQVeg5ccyIx0Xf898RvvhXrjBJ+kg+6ztHcVwpaM
BOXP85f/Nl5VnPnm/zCfm2F4Tikz9iClQtZatzxw5xO2TMa0KMk6b0By2cWbELkkws7laHIedOWy
D+vL2U9cYDryqFe0tBGXy0wZL6eyf6YbDMQcj7MLx2RBRQpPIklOu+IxvvGGIdji8siCUNnbZ8Da
3ucR4CpYWLOjLMZa4PFTqldzmCZontABwBXOyGkahdFh+ffOgZYVOnknAOP0GjRRX3aI7siYYBUh
eu7RLaXdTjpr2KkiVm77CNQ72f5THxv+FVp27ysf4IMZ5t6GidLZxcNk9TO79BXMfllet2msetut
guglFk8I7ooVK8aLTbB9ggpXQQsUHwt1ev5GgwRdzJ97/OCkOL44Ubo+anYcjM7QXiQ+96Zc3Lvd
FdO37aQUDXBL7aziiwh3qJ2mNWqdVztiWUKzIgQOwSSpic+ZkIps8Cm7qn1W3d+zMnTQ2GU/AK5T
TNyMfxF19r6dw9WgAHyBmU7Dqlyt2ew57wGiH2/ZLW+6fAHGKwGx9TZL1p1Z+COrS15V/5C7hX97
1T+dsMUHUBz9ASha2L8nvQ3AKiZsp3IA+3rn/BwFUggoh4ANJqq18yGSNG4Mmm62T5I0AQrJSxae
Ai14A12miz9FxXgZYQ1Y/2fPl6vxMHiP9B1XrWriWSKR2wedr7EVe/PkDVt+hmd7p/Pbh+t7vbtO
dJlhPz1KoQRjVPbm6RXzkU+CppMpeSidABhC9axR4Ufdmwzaqz3jOVgUGu5zsGH/yKmen86BdOSj
UHzNnjfCFpDcK3YYktpUfCO/6EYKx2CDSzA2AN47F/vjbW56lXIvbeD0c+wuWLW2ZgklW2r2wXUG
0Bjr8CaD8NnTxTS/6hXmuCgdXflnd9XCUYR5W9nbxTNz4tGKlTb0Rv7536+7DgEutqfgYfle6wFY
dZwbUdJY2eCcFrC1vNwNeavJvwQano+yvMeaoPBC6iTjA86XI9VxPjyCgZk/sqc54CfYESUay6A1
E7j/TdK4tZWRFG2+ltUgLYoik0oiEX04QLJnh/PjatGOAo8chzu++mEKLrTgonX7QZBARK+IOrQW
K4YgQ5AVgOQ6uIN0Gt4fksj5l+3dCQ1TaQkZEi7IS2gH04tnX9Wet7ofHyhUlzrlVujzpayta8Bp
0DALGvcW7QmVgxJ3qSBwhmSgBjh56zBftwLr/MhzDrwqvbCgogHv8/jTpZOsnWyb4es+pba8bMm6
cPWHOtmF5/2LZawMbQCNCMViRNAD73eMF6/yR7HX5oDbRYmzjnnGNEQIR2mLRHa9QSmAaK63TeMZ
+JekZJ+B8ajTzzZi2TVw0V8Ry0h9f4B9g5uawTCMRPkxjG12DE+H2l0OY3AKgEejwJfM1cUKecKk
VL9I/SSnpuu5iNxsKJVdiaJ2bAgyc0xM7aI9Urwbf9SxOKDjerb3/U5Vlot1zbSxna4HUT2Nbu26
h/fE+T3JWl2mwZhohnXS1I4r0qAaGHBOWhOjdYOkDvakszStGCIMuSrbZEgIHS8rLCLs4ZbZPbs7
bKP74MyNknwCJoZuPwLpIYJKSynjVenB16v3FHzsa2S9FKXGj5wDuWuBLRXvXqLs07KFTiK+zBtW
LjoHWg3I3vaGTWplPGcQzKv+V0vbP6oHIqSbWop1vw9Ed7Vmw1KP6gp9eZ41tokwRn5fVIq18CZa
RFchn782wIUrAZyNDAXDC7OImMaHdwtqobivmURMhbEfwQnosrxo8NyFgiWDakJTlkdEAKVpT4ze
W5OZURV8fe/tBRy6kLc7BkctJHWKx3cOSaJ/Br9p8do7hoQrpylI/DvDBxg4q0TOAbVVvUyyTKGE
xkXMuPwZpQWF2ioHGzW7Sbr3TMO68676MlqPXaHr/WUS2GqUcDhKCreWMGuOm1+ynZDCqeRFaEb2
olq3sXTI1Hrb3LyNIOI7AHm9ZF3j6h62DpN7AGIxst7phrlr5Zcs6D2gKAR+lws3KtKtE8NmtZQF
cslA13NXVO8okwYpYT0wEqs7CcmuH4Kks5PMKwG0/DCM9qF+q1iP9QOcJ9mbmAAEZ6c7mgJLclTp
KwTEy+2m8iKfs4qQECbseYLuWvqXcE1G2Emts/NkxvGjlSgwe2Qz2qvSJF7D7ioD6WizmzfOlt3K
v9gHD3yRjcVopHK5tR7s4WD/VL2hWtB/ZVX66UZmghrqEmgEVAOqV146KPzpzj1fabdtzxFvBwhi
aumtN7+PAiiL6R2Q2RggemHY16KzA/IgSAM6IscbRO2h4yov6RkHfcWRV459n463TxepMihBS9Sl
To4G8jBJxsC2iKpDmeX57zccswm3GHBjd1rMdGBwydpN/flNK/3jef7z3GCANrLOhawRDI+aGcP1
DgsT+GzGUxTgwteudDf9X+qGQ09l7Fl6723oTnBO+9N3rcG1Wrf9BfxZObBvLxJaooO4wl3KH5y1
jGeWATPiHLNz2mUPYs4MuSjPdhUA0vGJ8t8N5BhWU/a5KYfx2ifzzgE7bztRHtLYISnyHzQ011/B
PZXa7l54pDrevSaQPHD8fXg01ZYM5CLkeMfKvFFrbS0yDX08wTtlfmI7Au6oN3k0OhMnal72EaIK
DHoRRQGXBn4AAicmnU2GvAtBXlj/bFNB9RCQ5ax49CzffFCDLUkEYctfVzE0nOaEE+6fGdVq/5sk
phaTb7cAjxj2Zd8osjhcLkz2RNQaeVSVDqaKneJNXZvhJ5tr52WxOxIVCS/+5F0h9D4AYl6D+BJH
QSM0cODb84TUiNFdaHoiFVSFmvIpVdZPT1qO5jaWeVN147Q27zrOQI6Ne++15VXbvkfMxVsg92YI
Jog4aAJ1/01zJDhpDE2Yvwc6buO4fnY1eGmmeXdZzrIl+1Zfu+W9yX8KxnH75cZ1LwxWUL2Hea/f
Emz0frrE6BRcnNJa+cOXdzw3Ted+U4Fzup4eLr+U7zUKkwjWvymvHNOWXYB7f1+MK1mf6tNlIpyH
UQnUuxDm04bL7aUFphSvGQzaddmd3uVMWhoDayTmXS2KBgujg1WaOV9kpf6dtzg9y97kTRVVXOYk
nVhY0tIduWVF2nbaSUIjUwtdi727d6sEAfdcg4IgzD92mWBo7XkQU1iMjRcJknq3aDRE19XSVQNq
LrKWhb3BhU4IHhCaG8U5sZj/HkpLs6wO2aJQFJiZVcnafI0FrrTx4trlAO5+paE8zYJE5wSWhGZn
n6YROBItzkcBs0TvXyMeTn4y+h7hAt+nbT/ySicWSvUpPQa86dlwWNYJe8QvS4LV+3XeJJYq75aw
N5rmTeXeRlQ51F0jj3e92iBwkCPCiBEgTipyforR6Tsd2qTfLmA4GYPDKGJcF0Raf1lVOwsl2ovc
kOGx08cYnKiQYkFY3d/9F0ZvJOd8d8zqP3PXNWpQSBFvjLVFPzXTxxTvcuqK7g0GFyFBKg9a5dPy
RWmi9VVNgzrhfj1NzCSunasbRE4hE7H4E1QhrDi89nmBdbCRUisK4agXnJgflqNj81iFdVgUlu9h
U5q/6tP8B6utDzucewxtnxphlSjQOmBcNri2MwFB51dzCztyn2sTBNTfvdSDhxXVMczUwxYkWZZG
3LUXguUntLkmasQ68vXiR4a6XOjjkFs0Yje7eOYyLYZoZpqpQ/uAvZUdky/ZEb25V5X4ikUS/jxK
zlIpb4QnHCBHbFTezfiY70QwFW3nTs7xRMBOrKLLi/giF/gO+ItrklhmK0Hz5GH0A8Vlgs5EkFkI
8TLZVHAbI1ovz7zzXS3fUfxD7lMK3rOi6HWu91y+bvaeB0ULL1PUiVShr87MjaUUlmfxTThJ+/ky
Pmk+QVRIStkPppJKBiD63lVpvtKf5GO2EbzASJjaoEi1yQM8wx51zpJQ9ePPA0c1/mK0oNmpzuo9
BXZGRvvRKuv9AHBtlxa8f8LB0KRNsac3dUXAvLtt9wAHe4pO2y/q/Cf+yTlYekAW9ap6PJsA6DkY
+w3VKtRzvmS9s3cesOoraHdw9Yxd685JuXCZ7HytmDGXMsJoY6nQODMdCOzYAeknQJMJvbQtCcTD
MqxjUtrU60bx2V9uOF0Ch9wjHLPdrNeVWOkgNzki420y8jK0nm0F1kU7HspQxc9tsisA3DwcHb4g
TtjcWG2DfOeanC1zhkx74N55cQtJm4wBmWux1ckbjeEAc1CxYOv3pPvrx4YHKNllg6b2lF7wBC/V
PFF2H6lmwY1HE0hLDSyHyj4BWgiWb3hUCdQbnq5yIdmcb4kzBtDUuPEFQLVMtY6JMuv4WtT2mzBs
I6JoOMn2DGimYwrG1lDbg01TP7eFqM24xyggNwqUokfLgFLhN0CzZGfBwg/eLSH07bUW5Pp4uI5B
i9GKNp/RgRSX0VJI1hPV/Ie/HNZBQ9cxEWaEZG7e+YU20hLZTf+W/PcWYn79SOQXbFo4LtZistk6
ZXrhYnJ2JgztaolJiJlmqcKfd9dUPgOqrTbl90wOrUc+iHSRT25eF9WcBWFB4L8rgMQMEeECly2u
2XwHCTYKs+7J+wn6mt7H90v/UjMEDOll0jf7YAc5+mc3ZtFtBIH6RbyjwIN3OafliSoKUxXdwHXY
8gPmBM642L4PPspHLxzIHSr6pMc7GYLgaBonh0dPCfzTJjaGTunXWmD1ffTiJ2OQQc4DYa13Ukie
ugM23IoBUEO9F/lIMW17IQsSz77DUo/MTSkemXNbtpOg0T0Kq2b9stPThLiFnPluJszmArN65Dxk
Pj/MHERmTzAFmeVl5y8WXap2CEWJJPBbz4iTAsf3GDip5Veo2JXdhUE6U0eR1jiY84mtCB3Qf6Eg
55urP/zf2PrlNldDZq4vwfvtCRqqX4KRy3mbvsy80+ukfCO1otKGHg8vNfxLLEgs1hYNQ3oI9r7D
p7R5y6BkDUDz64rI80BhjucvKZXVFp1xdsLrThI8Cmm4fyn/glQMCp/7LjLb0Vj3wO6U+ErUpKhU
xBUpkm3oJH042JaRvfrU7B78KMTw4h+1tKl7d1QK+M9oBkfO3oShEiqRbretIrwxqSqEZ731hALo
LxwSerEmWzyj3E3wjFEDv44AFQlFwew9Kc9vX4XM4w01HIojLq9uK2wvsntSGkXtBfyD87in8rSf
RPfFym1kvCvMupq1I03i94554h91ire+QFf35aDoDNkDq7/BzK3JMglMnmgFzatCw7l5WEXJXUK9
BGmZu1vUX9QKWU8gEjA/xlT7QqVONzA2uog4OfVK1DucFzfow5ewBreS+P7HCoN4tRroFK0sMsH8
h1jeVXm8o4ythgNpFVlAeAPMaN8QNUtk75J3dYqdokiAHk32LIzFhqCYBk4/AqKmCOy2Qgf6HcPt
bY4fiFBCAIrRqNP8i/hiCSwff2EsDlrlGM/t/xiqNLC5aAnWGbDDcMVIo8KFWMY3RgWSwWNsLmlx
cyl8vhy/kTb9WoOHNs7NlaQlLb2itUc5l+bo9vfl1t6+OMW3CiHjASNo1OfaF26GX6OmXuIT1IVc
iGJgreGpOOArMdWzTheopM2pW8EdfBAIZ8XR4D52leO346jp09F86D3JYIoRAt6ksaYWh9I7G90C
rIfuQ1CWfZHNpf2L6Oc+mFHGLt8XYOGQi79agTe9N1Mm+SaKQ3J8YyjG3n5F23Pvnj4pb1dmnFfB
L+ejs/xjUwWSBh/1V+n6uucwHPnAmxdAIfRGaGjUNFyIaVOo3iznmyuz6IvMnuZ+fy7G4HLImWDZ
Wgj9wW4+YSNSLatGGStV7juRUmyqmnCkkdw0xFpCiy09TakeaMqLEr3Uss6ISqzbjDQZUUZ51UmP
DvYE9Da0YaDNIBic0DoYlqSDRG6alXBeZIlJ8vkX+jcwL2bB6ihhbcxg2DDAnHHyKQSyWPGQgHxV
kRpUmih+MzGA+ic9X8QTxMmHYXXPHPun8snHJjx+r8oj3aXaYB2oqaf4Hy02FMbRxF4xzRyCUfJA
GmGlmycTuiS3Xt+sxMWyiT158qK5SQJiE0u7Fcjjtc2U/gtsB71gYFNXxfpGYVDfkcXLZCdLDqe3
x+8LYF22/z+oU97MLG+WRhdbSYwBIPMJkdP1SjwEMOeeStzLc9ov0MuCa5vJnw0EXiEUBT2aAwtf
nez1BWo6YrWfH3EhwgUQSc9WNgnuihPkZfBMiLun/5sGiSgr+A1aIvIlyOrhYSAjyXh/rZ8Appkk
dpyn4gk3G1ZczDxGh9bFrrd7O91SoGnz9RIgq9H7qr4MTeDweyndE5u8gxsWW5tT5G4xOh6Lu3wj
a8MAmpoCA2Rgj2PmcusWxeNC31pj7dyyznlzkfGhbsnXE7s8dbRnMnXCER1GrZPHIrNF/wR5T3kH
s5/jR8L6Pbrdof4gGVCH3DZFWYOnMwJzOhJq2WQrRU+zjb/m1dEqipbvGaVoUmDIdWh5EMnWV636
VXpCLCqA0/1eluGuSSf3qt7rWWQfRnKFzp/WHGFfG+8k4VOFRS6tUSrxLx4pFpv/U1Pn87CkM5IX
jdMFo8jRNg6ZU7Ll52FmJnSk1Ai7pm8QVTUY6mtXv6esrTtHzJ4BCQ1aAV+LRIAZhvjOEgqgpEFa
aROsQnxW6WexeH4aL/s8UlmaeE9gbAQ0IF1Ym2sBfUTFa2khtXwbjQCt5ph/9LBzw3L4sfncx8ZX
cfGWWXq+WtENA6xZWRCLzP3H+LNdHuyJQaRmO40bWPfUb/cFilMcxO0i8nLeU0REl2LZHfk4dheB
vp5JVCa7CskLUI4rfKimfcGf4o3Q0+ANQwcSn08Jog6QNvyceA+7x0SfpCP6aDDcmPn6tOhSskYg
6SD1EArIv024T1vo7nJ5EU9Qzw1JQLnJ+d5K34LpcGCgvxasG5N2CMKj3oCaLGs8sUhoDFGmZT6u
aNFnNCWGPdFi1puzr3pz/wvJGADNG4sl72qahjPUDyXzMjfaZWyS0SQYyocrKYeWhnlhLCNcBbfK
nWtk+3c/xK9+94reaJwKeaawzN4oaMx1qRj7k6rTlTA1G/z3fgVAdxeoPp+MSNIVSRj+MD/fSuXA
0XPsKc/Y/A7pcpZYlqYlXACiM7hGoBk0pPpjwet8e8N2DhCV2mJQ7yUTwAcvaMNPrTqX/6UoUnI1
0nGRdz81EjlgjRA5HXSCOt4JyCcWm0Ie1+sx2FWCj0M/RU2dQT7kxFOvUUz36wByB2kNx0yAzSa9
hB6RbTgJD9HmzYB/AQw24BkgaFqvIxhZD7LOMwxCMxi0oE60wcqMl7M+cDg2FBFxdrP5IOwS5vex
J+OEx1k3M+zn7C9bc4ReWxOsWWWol1ynGgW0Gzn0pgf9Ie6fMzV5IYKbqQsc1FpdkdYkhyFtze9X
wclatfvgV3DXoiy3V4wYGPZ6jG+D9hYa7A5UcES3uMFbNVrEN8z6MFKRUPZp3EMi+aqxFdjBjQ3t
uD/N5sq1EQG0EEAYFw7aymTqybDqvsePRuFrZ5CHN7RK2xo5GsVytBoxiP+BvUij547uMabYxcS9
HMFghvII7QP189+uS3xSbBX9cmNzp3ElhGbH/uCaJ/li6BgDqOuy2Jxi48IgeN8UM6pdtGGoKj4O
KpNOn7ocZQbB/JlOz4HKG67Z1//cQssMRxqLKRNneNw32z4HTqYxkJ92/eHJTSJ1sqF4Vdh+tZbT
5TxbLYrsqTdA8tLJDX3e2BEjUctdVlN5cD43bM40J5Ck10YP2uXiWJBF289Hd4S6Ucqs47GBxhbl
0ytptau3PfYjMNmOjnaatx93X6lv8AmmQtuBlcIw1Zsi2UBr6fXTnZlfXuI4n4N03XmPVRmcXQ8O
Uhia1Fx5z9yx4SlCzCbejKq/1kYUrOCl6h3lOaw+gndhRuw8i2V7xovCKxR4Zc8j5boqeBPASZAm
ZeEJ+qyiaC5sMjwKf9JVya/d5g5icY9jbkREpFOcuUjnxoIpkpyvwJ+xnjAXMVtzcPXPLPU4Z56U
xn2HJcRjMcsqBJUuaydjE2MCg3ZMAhz8tk2JM1nZC15dGM92tf9fod2T9V/5TNdLoWHzjhkYq0b6
RLQW4s0PINxmafnrLKzsI6vPEzmcfdqtgXK7oUNayAo9THpz0nIyR46quRyE/rByxodIwNAjWN9u
FLHsisl3moPBCNownwyJuvAAy+WXeG9apgo01yotoHsEMAyGCvjkUjLEkFh7PBq5X3n7CxrhV0SB
+bjCocESef8h29JwiCPhln/d10yid0pMpQfUJ6uuc5zsjpCjBzOZNMbN3TPQqZFnZKwOlWbi2TDt
sBLUU/yPrlWrDqCrQVEfBtT//jn9ZBrQzByixIeYDgDPHROK89+62DBHLWjrhJcuzVlNCqAf0/Vz
7faDrP7bckElE4oSmvF8IDuC61CbkfyXo+D2D2glO6/pCS5mxVseSWMgSEIc/91Ek++Bf/itZfVO
i7pJEwwkIZY3hd+rbjTg1V58no9AOxmyOxsAVlMxQQ3yOt605glItDVaY7qrBWPbHCoQ5K6TkrnD
ybWIad865A+zrfN3yjlQ27BQKYI9oCZTWbWUTYe6UDdVqVZiQTN/KJUOacVVP9QBjs75tJ5Gr8EQ
LYI3NcJUsZrOATtuf5OMhcSSNbSIEDW0ASxctOCCRmSGWxumAmD5dYpI8jkyE9zvCYhVd4cyidKY
CbcD8nWIHiLp9J4Sf6usiPHhjGlp8wcGfnFYFZBdJ0CVnGcKrPD9aXdsKn6o3XOcVv5bYRyRcxRj
fK7MP7YUtcRNczfI+25w+i9XUMej2XwxxnJIag6DMaC+pVqJ6VVaQbpCUoFrlk+bfQmsWScxkcOX
jFp1EwM5Kub288+8LrRNYmsVHgMfpVSvzxV5bRNakorUbPjNzUeyfBu1th0FrzwpCL9yBHSoGmYJ
//x9e76xe39blEnuWggipGhjyBnmpLr7wFUKu7P29mdZ3CRXKeUWYZd9J0XczmZrCV5RIWje1pdo
k/6RpQ38c84mRFhNIW5A9EgDmwS4t24wpv9GlNTMwZVtRFA3UmBf3Icaiw+A42En1Yg48lkVYsWB
6m2OwW7kceaBJWLX8zGTjN+ZBJDzlWUj76c6R7WZ+EmRaCNt3LvT47ykFq1t3YpSUDihuWx1zqkq
ge3egjyqXenkeyjElC7imye8Iqi1vJ40Iv6YMpMdVa5h8jPuUksTzIupNzB94/UXJd6pQYXkWiG4
BGQmOyCge/tH0M+HMgzcW7n7dSOeYuaPNX3dZte7/3QXvgcCeWgA3NvSTnYhr8kNFZ0g/QrSgbEh
KJuBDS984cOQnbjJOZ42ySo199XPaN+C+Gem4qLLcvPjYxf8vk/cancbcK3DyMPuq+2YEqs7rR0V
1FqcvVV3M4SUuwlPEJZFdSZZF1ZEfNyN/fldLs95XdGJjSXKXJVIgYbM2t/kndov2ub5rWh2qTd3
OMGmKatE4/UfYD/Xclca6pvRFwrFN9c4qhF75MAJvz2jEUcDRQwVcrdPKp0hTHVd68x+vhwPQtMj
FcbvX0yXY1T/w+c6QUsPi1Z16BUnL+soXXjieRjsDRB8L7TJW6awExJpVWx5O/5huuvTFimiIKAG
4HGmTLxfXAG4kUtqUe8HkPTE4boxT8LwHauLsRzogvPkdDNb01PLsASNKUtI0zRQoAFBVlKy5hKM
Xz1/WJZ9N+oXW0Socz/L0AnhUeZeG5bhaSVvvu7JNkNUqYpMtUkjDODJB0DE/EzEIKZHGfpvys2s
e/LD6WVI/99LBConLw3J4c6cBdHKPDNpBU2koaHukxXXZVtz7zRdpA7ct7mFHAoP/MKMLY5e3wUJ
PSENnSwmmE7IuKrEk2iwIE9mFbg5obfR2AGdClh65ZbsuEfk/41DGAldotR7m752ej/8Mwp2Ym1a
IEukee26dsVtkD+A5o9FpWMJOoJqN8Wu/KqZnjsgtiAKL/spSCjzjUa3wRo3qOVuQ9X79+nFqoKp
x8G4sLTdrwv3tr6lw9q8EQm7oNQ7G62KbnrniV19y3T5zHQcY+dVykuGSFJWVbLaFc9ZrDKA25oi
x+LQh63AXQXrWNuvxim17F3NCyxpfcy+b9a6DMOIUOP3bq3hbB5SW/Iu0ZS9rYW6SoTOxp5BibZV
FjcXhmEDQLnMkBJn20YdV0Qx7fcjcWVFO2unLHncLotwPuJl/uIxDNWYXtiSNnUhzWyvl9MxhMY5
Y2fbHvkfPI3bfhEOsLcYzHOxjjovz4m3Kl6zAE2l3VZjdOc1ijYrYuCtoixLU/DRlSA100JIPwy7
cil9AEuRqWQe090ONnFQSkA6XWDoHZjELfeiwJYBjIKUUdHQowgTnKCvA5GZnt67/woY2e1F0Cya
/tL3TYs17RnpkGoNiW0LjcET+iPK1qOK3f0JqO1+mAe3sqTVOkav4zCCla5aawgGXtysicMoqfEO
Zhv1/8Zle7WsuRi78SbxNCms6qyrwKjdKo6sNPfNnQNOktng8CFJsp0lCnsMzQGaj4qR/YTTMwsK
uK4dK4AQjfNpkghj2f2Z11XnNrz4pZ+yaP/tXAxood+wQBLHmiqwm9CAgy8w6DMKLjQBfqkSpMMe
iklCre+h3lfbPA/UdwXiUrFYIsDhSpYrkoQrwYwIxEqokefKz6klBwyeoKwElBPgLswOdymInPeQ
5bup04KiPCwDWkyEIUFkoaUDL3KRvFMlF1ICwk+Aq3Ce+Z/lW73jDUZcZfQuXKxtdp+ynLqg0Rll
IaqmJlzwFCMeJuaIsYCkURc+8MGD1Z+KOzGAGBLW72G/xSV+V88GOg1Eaoav/IB45VaSkiPTGtIB
O9mdx8lpdCLeWG7k99DBKDTZin7IPwtJ3B7glUnV8Y5FCM/M0omagk3Yf/0DBHfa3bRdVRaK7UJ5
g4dG6KGaXYggScjRy47T9KA9As6TyjXvj332PGxk98QrIGdR2C6FiSD/7SuIa90/RcLxSkUY2nJJ
w2/KYYBEnRNwo4YlppiXh5GVCJ3Oud0lWeuCxAz5MhjewJ0fjpnT1zQKq4B2ewmJQy9yMPVwDafk
g4twn0Rv590p0vvkJLxeV4jF+9iQVWBCML64vTltEByOkkNXwmE+7CyiGaCFjhpLiddkcY+NhAu8
0nQ4+s4JVg8MQeSzUB6HHKHHa8SDbB0vpNciZbVEPWnl+CsmvmYjxHcJ+2LHDKGnSe9Q1skmH4Cz
WQFCHXefCl2UOM7ATrn1b8ak9/KFwj7n2WeGCXBMu/ZEhPR7mPitx20sjvtJk3Gh19S+Qg/cx4Tt
t3H7lJ5/FXULnUpEfewa2CB9RMGinssMFji6ddRytEjqpbb2ONHjyuQQ2hXuQLOYlTnW7E79E7NR
+Eb0MVEWw2B4csD3xXrBY2moOB4SqEb4VRZBVHGBHEvSaaUF/TauKs/ZChlgk5jUV9M82QqP3Bbm
iarRh8Iry+kaUUoFjj6GgC7TvSr+1CgLHD/wS5LYsRDKkBgi6NpWhex3sGCE4s2Gw+yr5OZumZ2s
iXnw4CQfb8Y2uXFtJ+yEUVBnxqij5iIcL33q2vscXQlkGE1ylQJ+zvhxczsGEczjDP2W+AhFsY3d
gQTd8yEkBf9WmC8+KkIQ2Mgi3EajL7ldOJRDEiedx9fmgKDFF3M4tpeHVkt3hEKwYSLTRIe0gagT
QUgQ7mdbOn1bjm/a+g6nFnDhcO6Te5t40GW/OvmCUHKFjsKermgAe2G42BIDceq2anwz5mqvi18h
t3gt14ZxdEx9bRJ2r8rX8YplV+K0OS5wlbpRANx+YexlO5Kzl7XCNtK76hSXoAdedlIB3FH6C9f2
KW+9z1ZkG/wgEi0UsoT21CF7OSj/V9JND4kMAKiPCHsKdgO+XkGzdBuHmzsE6WoPTNBcNuQvmJ6E
4mRkdH65vd1helsVc0sHJbedShnZxzJ9DbFRHiPWIZW7KMC44KPGqieiXXQUtKt4rRID1Gn9dHkr
ht2+H4W48mUP5BwVcjHcVcKt7cgjnbX+GMnJkbXfm3PN24MCq96GSt8Qi2K3pipaUdJsHBIpnASb
apIVX/ow0aVhtkyOzbaczproPzKb3ZAMe1t03HJV54GJFzQ3jjHGGxZ3S7RXT8d0wD54rn6O13yo
eTQ7w4B/mdORbDNBLSLGspuKGU25zP8pBN156kc+t9XE+Lul1e1RkaXyaviNFzW0LAz0G3nN/rKf
9q7BmzKfBoMp8nCJeiPvMJVSRfTsFOOQG6FYnQf7XQ/p55MrxvC5BbShO4gUG3Ab13B62r6Zuj8E
Q0wZWLnqKgqBm0W+G+bsMhjYqWJGh5TFbF0wds1q6HdGD0HqjU50HO4Z29K6jEe7gS7/oCWwJYyZ
gqRTPbP81SFYK0REW0IckzT8aU+wa+Ssi+vX3DV9B8dJlemtd2hyE14N5V/L9zsII4nZytQ/6jMx
kcBGpNQTNgt1HzhlTk/BkYMbMdG469CrBCsH0jX/b2ysyik1nVZk4NHIIAmV+N8af25rAn6tRptZ
IY54la4X/bIQwXCShia5x2hrcXBs0F1kaBCMEZR8pSTj2TU2A77GXwtROKMv0biwQNmeDExKdp67
kuqWKvXKtixlohPKNjwot3OG/SUGXhf7Blg/cW9DKbO4mbPvFRq6BIIqFoSn/FTORyyLhEBDmyBk
4SnQe5vUuKHo+wbJehCOZcsKCBxDV6jIGbsFbAxqPJ/Sl4MgmP5GEpiW6wYBKVjMcJikhQxytzYb
oi44OWksvSAZ9WTgPD0IL6RB6Hem6PkW7e5nb/qLbPuhAStVdiv6m+pkQTGCFaU6AgU+P5EcS7Mc
JDxKMUptpTQDsfGlDAaPvXInpSIyFI80vOcADdxcXudy4qIu4qBQYitkBg+RG/f1Bx8if6wZd9Sy
JAEfmkkHuDo2baUmiP8y8aoZ6H1TfOCiozyyphfYHCnUvBKkA5oF7H2ApFmAJW9ic0jsBJNszxMS
jzIJpcnL21GmQdY8kugxiXKzIS77VWIZs38VLfbzpknq7aD5sPQS1kjyAlhhRSxSbUPIlEfVuPr9
P2d7bSzspbbDVGiOtEkLX5X6Y7qDFTKw4Y3A25AUISgWWs7GRg+1xvKdG3qJ1bZWel+3XgMUDPbs
k5PT+RJiHaJjiT/QEWXYhz6Xegaynsau14q2e1eJY6r58DrcACXNdEL5IP4qfJXkqol1dsY3594B
e/bdXSaOMTpGfecRE6oyUiYoN4PY15z2sDWJmt7N8PKvsKrRH8Pz206qj55iZXx2mu2gMJ6Wo7/s
YrcporbfawXgr+N9GBdZzTodoUUqLgnIP0i+cy+leCypb6i499POWoTl6UTCbbwr/gq/YNbT00xj
WDiVHjaKSv3jFxfaahQy7x+SbzywkPU7w7QkfesQIZ2ojMiUIZrs2iQ1m2ZldhNGdYTYjyiPEF8a
q/4cFHhOjfZFDXXJMRMFIArzaLlItkSkGLiHaznPB1l97/gB03p26YNNylaoaifFpscoDwgxg8ur
ABEcuU91AVpZ0ZbY35K5hb9s1R8dHgB8w0SwcNtq/7aBIDTjUejSpqDoOPkhKUeEUyQYO9CGI8e6
LjMVqFYpa800roZeUveWs50iz3qPObkK5vCwWeFvcyPCG/XE5p1miuAnEsPMmUVGvj36tGbir+10
PFzxQmAJ645DAgXoyKjoyivc0Y0L/TdA+iqGPWM5lEMyFKuc9dgr+Fr9AUsJngNTErOC48boPTPK
2K7ARqs0bGjcb/GuwR9LU0dnz4ME/X9lY5crmtT6O5m2ZwTUfX+9JsL7lxXix4O9172utGpfr8K9
kLivERKuxo09N4dO37UEMdX4GzcS/YVgnYGLYuRN+pEN5atokWvUkPg4LnBhbsWf1zQptZuPj3BO
DmJrDO25wMdxwlimbwwCvR3cyEzaWCtpsEEm6ME/Jf0qmWMqhlj3tGjiLAqyqHJ0Ml/eYNBQ4IYN
awXqr13a9+i4j6zRDrHVKZ5l33er+Svl5CSAfo6BUg3yJfK0Jz++3NkQ3/1AYO3IAv2e5qUNoo+b
R8mKZMG48xoCl/jaTmjnM/VjtgNcw49zhO89wXs8xnugufzVFxkAXI0fPlcJbFkWh/uv6ci7AHDi
ARV6nR1quMcqPEnhAT10raK/0Je3IUsCZm14TtGoW3/RE/uFwAmUjgow48arK7npZskzLfrgY5cK
Az3e3JhW/2cH9qcFcDOhkmWy0SjTNeino01nXeCkqXlK0d7QGcyr3z8ms4fobNGwjuFMRHaqxsLC
iL9LKIlhC/LynUnNs5uWpeXLGRuapIqs5/oBPCSQaORdSH2whc0sg1vDn7wnLgS0QAeFkCBsOLcH
ccwBky08vtpDRs+CzE6eSp7I1iy5V7YtXhyoMAFfKQUroollC3hFGd2A1BG7BF2v3opMui+uxiH9
IkGYYkBlIol7JHpT/1A+QpL3GQfPeZl1cVesSjuwySh/5VnWwrDiKl8TBsbanF/bi7DkTO7IRehn
HtV1eJ12CRbZ9RDAcNZoXZGrqETyE5kCvTUCJzhLBxZEnNQQBmQOT3YSxmZridW5Jl3orwxhNSAu
gyQK/gaSWTSzrgTpJthP7d0vlY3aVqV2d2YD+zRapBkbEN7w8OS5HJNaJfwRvgaRCHU4CdE5rY75
Rl/RMUqHah84WQshdQ3Qn4sBIcQrS4PsEyxp3ZP4bAT02F2+wvBlAZIMbIw76BH3eyLjJglFWIPq
HpW7KW9KQ8OJH2rBzVqmTPeee+6AyGAmWh1GgLALsBg54XwDP0AfA8KtcAQJIL1h3HrQ9Q2vCUKd
cxDxkpZMiX4Hf+KyZjrlqe8bM3Rm5QYWdJ/uLef/KcL3X4r2aUfe3oXJoZgi4bzOm3qc5Btb7hxr
SNilemlj4qJPybOTC+4QM3GEyKsCgUzDMGYAXuHKQRSFLzMif84Q2+y956NA4l7ewh7oLqJfRXat
GAz65/a6AOWm+1+0dkV1HeJrMS3NOEZNTn3LT8oPOtyfT9dgJ02XPZYs0AhZaZeYWhhmaGVLseDq
znCAyzxcQWk8blTdGFvTacTmd/urhbope1pKZFfge2FtBThAOzxBJuc6jFOBInVxJA0GBAn9XJdM
xqJ3s4K6zINvp2X+ZtAGh3sWvokup8E3LLUH7FMGVtXFe4c5SQbKJxW08xoOXJnXuouqt56S3h8B
P65pw8TCvBSse/OiV8L4MGRXiDl5mXGiKXscrRv0ILTm7AQgpL2cO1k5o2L8+UN+SuB1T6q92dae
0qOIovBvBBl4673bOD1fLiREjhPoia6VgKlEhZb3uJlNDOmF6Csdrv9duW4IdKbdocaVb9xpAvLD
f2ZpG2I6BnR0U++lDkq9YpUTDUuMflYryI6gR31+ehvlQ1x5F2gXXseWsIIPMuTCKyM17TvDZruD
5aKU9GcJ+LbR8bSaCStykvU3iTTK4DPiNVLXoLGMa32fLX44Na5d4Cz1WAzOZL53diznoYer33yY
Dk63d2xrs3BVyTj31O3pNSCGS5PiXi2RrPgXvtCqY+8i0/7P3dolhtKlJ4cSM1prHtVEc2kbl0LI
lGrvSws+1tBiQNIdsobItdLt9YvvQKWS0PeQnd0zWrtJm/Ty2bLUqqmZzkx2feZ8WdoX/xyDslmf
mShYD8ISCBl5BGb2anmrPyaiojcJHR2pVi0vgFXGctbrTB4koZ4J0s0vJKMrFTKwrMIlqHHbUWRd
I28+UISv6H5R3QrdrNTKXEo4LPmjZKU2CJXixuIw9VyLmkZoWYf00A8R8eSsjhsTg6xEEYH9Uzb5
S+SdiqvOyf4Qg0ufuKSNOsLqzL4FceIAIeL5BJpWSFTYdTX0p90wdHva9gL3uDzKf++qUNV9WCqP
zekZIbsgBmo6iPE5GfyN2bb4UT9A2J+mbBfdOu4N8zqWXf4GleHOvFbT4MqmDC/h6mNNlJLG42Oq
CV49Q2xu2dQBDfihXSIyjosg+MCfI+sfdWv+rQIpftgYOZoUg9nshv+1lOEQgM3Ymvt8gbkxWVeE
oDmOiiRZ1VOVlyqeKvCWtZ30se1RGxpnoIwaciYraF9P6sMoGBdrwB1N6rmLqw8JkEBLbR34Yazt
p66nbYQba9Z3Wd3dnaQqGh3La1Qgrvtkhh7Zq5dzNDr1GMDJrteBu5EcRNrF4Ry6RTVs87ya+nK2
DaIuf67xWlf+3UOyCN7OnO9+vPlGzt/jLVf59KT41PMs0eH9ftOrEeaAjc7ofWhoVnKm7E+cCtYT
kjMZ+/EM93YthOcUO833tFMWXI+muVe/fivPR4MceqqiEar7pkhGYiXUoqgKUVG+RsQSu0BpUQBF
gj+vo/N9vXdmBccaa6RuwWiSjEsqAxTxYIFyvjlMY2Rm07GdhFZOV0H2glZ4EUebix2ihTf9JdL4
Y76eM0tkF5noEDLM9Jurs7MfsUyQSLYkui+pbTbAfX34UQTLfGx5s2NlXBNhX924JB83+ou/BBYs
WT3TZTmVqYUUs8aOq1xxiS03yuyk+usCnWDEep34hDQc0d0ZEmA8Nhny5DUVVMcDV4rWILnJr1uu
XTSqZ26vDrVhCflpSET3ZF1br3qEKcy25CE/eaD6AyYgP46EZ8b5BCQhKufFj2VzcEQHYz7HK3M9
PETWYLijMcw1xqtFFf/OZ1qmheU3akw3XWo6+5Tt/xGGKTvHzK/EAvLUffH84SqzfS5U05zKJ8D+
NO2tD6rGf55s6SqjTF4VMwDa/6wv/e1jSSFJ61ev039yK6XsU3Nnmt7a8LYQDqoMVeEW+Eu6horg
uMPZwRulrNHkzLpV59mSPpvpCXW1QWKM4N+29QGLzBBFtaOBnXerDrzBzPRK7gQjnqt2ytkxbbNb
1FVQMgwAB0zNMVvpHrL6ZFmmXP7b9d/zmxqhvlGyyh5yjiR56OFY0PSyk72t5uUgVGvRCNLFX9aZ
mRlJtb82XGQa0TazHp+EragW/TxTBVZS2fOUDwVDxH17OmE917yUlZXZDdTJ99e6aPdPOC0gjIVx
JoMXQc9d2AkgOSZ2KJxrKopxOMiczYeU82PgDHFXYu1GQqrmNDluAmqeMBsc8YKmdWHqoBkFbisM
Y76KmnYclji2yQG59dODFfvPETXdsB+2mVWB2SPuSDNLQNRjFWzv026mxRHOo55ezfZtur7t/ilO
/QTUd7wfe9MG/EhhsNs8lvCgfg4iFBl41uSrQAENBGKDm8k/zoyTY9wouVTT0SC+zpYLnXUdmoiB
xlZAzKn4shlUEjdlyfjuYHdtaZUPMVHFzG20SxSz9PISVVUXCWeDuiKb0KlnVM+DQXuqF+NCNU8p
8neKIi5neOJzWmRZVMGlNcAEINa2eMQoZ8W898Fwp3eU245crUOxsYv2F8O+mPjgwpkRDRFMnjP7
rJMTBtlWnQ0fZji7T17hLzM7q5O13AsFrkfT/CIOnzUPuWtxdBnsdlSwy74sXRfq61y/CQmm/jlA
lmy44bpY56mdPKGl++afklcHJESV3PBOZLtjEbr3Qjk51nOCa768Yghh356LkNCbOjGjCTfax5/H
FLckdCQX//3FXxWUVdsnabEbymv8Ps0i1Lx03copau5bDgfjhntc1aMa9u/Gl5S4gJ80m87rQM5x
JuekCPWU1ycyE2sjpxyoYkfm8rlld9NBdkBmP17VDqzxnGYCfTkeuIyC+quCIO2bq1u4YG63ZPTQ
+dpHFZl/zj5Lpb0EguAcg+zaa6+PmPYxa+yUZGzz3S4ncQP6KXdrRkzAJKMjxeKmot2Fj+7CD2KS
KJ8CIC5vCy1sdNed4azoCFgzAbdLXPjbj41zvwTZhdYvZEbzzpdENNG4dnH1a1yEZkDI65sfz+3h
VPS0IZikRYnkIL5tgY1mQ35SXX/396XN/YuRhhPZx0ko209onMoMsZ0PJ1UenBQVka3rxVvq98AE
HXVcix5eRUq3TDP5lY2mWl1IyL3YIQ9xzYT12wEITBgT0Kc/dbWGWsnMOguqzB3KLA6WFw7HFljy
ztoJfS2HlTIFvDanoXuSs4EUAxIq08kNdU+pImKIol/PDdIT/SI+usvh3gUPPMxeUhbEgq2fX8zU
d2aUr1kwBxUlJKHLmdtobFBmS3Todclqj5HbA5l4yLIpTxoM3+JlgvJLvMaBCZShMXxZARdprNiD
Ww0xJwqFJt0BHDGqxQNH3lBor+VnRcoTY5kMKrm6TNfLnohpE6stEsfyTKkvsk6spcbQs9c1bmgu
mb1IpNxlOU/zAQB/Ckqkj3PdQXTKMOp3B4VwBReTuk54pjF4UDWXRxrl4WEWQi2xJUQk6Oy3PrE8
2dh1uPLxtqOZh6vyWohHW6uiT4bFZnpb5NeKZMjEpEAbue2nHd/6zY0gGbHlz5if+Vr27pmuFIr4
Idi/zYF+dRa9ynpDBPQnflf7+3nx3iT9cwa94a8teOfQqX8XloiOJ2jhe1aynYroUTVSdE+6J4NM
XDJYLvFDrQ6vG7YEL3RNNdqC2sXsj1Wyfi1U7UKsAshbdCMvwANTa2Fda8wns5PbKJacaDl0vsXJ
NFaC5QskWJG2t5kk9wrTBJRpwwZ4UIS/yVv+9ab5CTtroT+KhD2ZKIW4bsirXtRT2mubHAoROEDd
dDztGPOOOrQDoXq+OweRdIaSRU8k9oGNx0uyoUVQR855qX456WUW38G61i9EQORvc21lqcHYve3x
yrUL1/ok/C6M4oZ1msEVT46bBtpf+MZYBC+a6f6s1hkd6jJfRIPZcmgxPViPhn3S8PLFO253Zm2L
CTPzwQQGl3qMtsU4082vwALP4PxXVoCSy+CftrWrL1twfVGQuh4V8HVVynRFJ9hJpg0VddqCy8R4
1zeszeBiiEsI0hFnN6Fxn293l4tNFg5Yq+kaADyTaiNJ9SJdatG/dPwJQvyuOE4EGVFWdnikqORd
k/rp2fdFYJfLvbmNkeIQoLhFTOVePZ64LNDY/YeGyl0RMm8jQ8r2MwmzcQBCBqJxaCNGtp7HYzP7
0GIUBEprhFrooXpdRfQ0uz3MJ8lkCFQ+yoYLrCPd0bCW6l/JLbl0fuvp68kVNIaoK+yLGvVfX9UK
lxJpe7RdXKIfx8YsqNw5/nq4JZq50ctUPlbQ8az9SMhwq189SR9WJ62zLyRBIxIGPHGfHgT8CxcQ
KjiWDXWu6yeJnns3Xcxn/HrC0/NP3Sd+wEdzQoD0q4GL07IV1GMk2tV/8yJvHPEWs4JelNBINjvH
gnuGu6G8q3+8IRXH/lGgwey9acVgQnAzEq7bLP4lhzanOcb2ax63N9K7fPGf4wTcVIP1+RoOLOdx
hLWFeeI//ASdHsZZLaQnZZEY+b23cmhUWX6hgExJe89e95dZqUc9YNHEASXh/OdM02cELtaQxp4O
kwMgozE+dl79UmlHbZYpmiZwWRn3MgyzYKq8YLtTuZ99dzLR7FFFVwnog4bUwyqvoNAtwrRgCzNo
LXaJCW12R4MHh/D/WNTuCKKd/FnO3+Yq1u5IdjxaMzDEjkgvUj6GN4PzNHwZfEWn7Tx3mA+cqN9A
eNJEQ4EmO9wG1JoNEAAK0d3V8aPhmgYmquKXdRl537HMWRnPy6CC2hzAP/oJ5Cg5rbJdlLo8nn0O
U1EddV7pECHfSO9IOE7lUUs1JIWzq81+h6kyaD2mb464NatB5PrPbgpzdQac3MZ5vE88aDRYpPEr
QvGGzaFjO3G+xaTcrn+b94oyOkEfWV6//We37JWNwwvWlhqzJW+NOrqchF5jNkcGpShiRcFC8AIV
smDeeMvizAM6V6AKywgSUyj+frSF1bVgNs6t8K5wIXg9QKaPIsueBDXqMjmtdMhHVlQVYMNqkPOL
jt/x7ZPM5ZArhkFLVr2apUkE36H/lQxjVE2Yu5qgX10RpHYb5Rn/zLwD2BO3t45knPuKrrlrypUb
qhHRVr1pJLgms5CTf5zvfSpMZ+AaJUafPS5cif0WaP3UW94SdSSmEAnueLSQvYBgwJ96Zjyr3+IW
x2iZ95h4Lui042MDVqb8kgsQEixB9DB1FfiSmPQs7YcY6C+u/mgdEVrN3J2XPzesJQoWexs2bi4j
I1QacP5juukv1GELYON6YLKXN3H8bs/PQdoCDbud8uvjixBIxO4HPJK/OR55HBDK2EOl/JSpU1xJ
HVhgHdlHggegpaFW0EUZeTS6XvnuVnalSlL5jNsTz+jl18KHLKyXv9L+R6lGdKCza2+VrRhgLOCb
JokFX+BbBqvtCO8ccMST+1OqaZgrsxOdag47J+ytZ8k88tABH5qxCiqNQvx+17ychDSm9iB1oYKF
9R5hl3XmIkiCvglzEXg7ItSKiYL9zIRon1bdhord2ja9JblroqSbT59owVeahO4vbCpyMX/ABvDR
D9WhMkEkPFbgfehUkoYCBMQhSMans0ObZWuLQdijvdEeKSOYUiQhiH6LHp3JHvOvmSsxjbRvjvje
cDfIJcpiqA5GLaYxuVD4vQmbyRQe27kG4Ad3q4jDgshfY+BoMR0KpIXLN9LlicMHFDHBnvBWL953
DKrnn5iABuzYuiDv425f7dESwIUbViQrxNONmv+h6Fcqavhl6q2efvwv+CNIBidg7gt+Q5gOELO/
28u4Bwb5xsJlhphQn7kBOUSsiLM4XYi7Y4l6tiMI2L2Lr6Iw4ntTHFtQzK+L+G0j95TLWINqZFkD
ExB0GvvYXF+iMGrduCKoAPA4ILjLhJ6ACsR49/AxXl6ayHc58dYDXw+clFatTBj3YQwtWE7N9Gq+
wbok4OqWmTY94yTiPd9H43fEvM1T0tRCm4jNFb5sgQQobgClXxvdqvlohm4NidTRUIR9CeivRInD
4ugmW4+rXbzott4O/X+rTgg7+MbjmGeyIxu9wIiKJ/gRp53JMKEHMvlpLo6hhv+vOuU6tcN92Dbv
1bQuBjZe09wHw9CCRIpuC8pQdqBCOswEgaqj5ppdbEt2NP/1t1Tt4TGSehaezZTKzRRc0oo+dbxM
+FNWPtBF9QFYHnTfMXsKy9X7hWDblT3SGvtxCprlbFoaG8MN1Fj8GF3yKVtSJvR4f1v5c2QZNndi
7/cUhTtFkkLEXSbQX1JTkL+ecDR5NvMcnaXuzUb4hAYh1E1RnMYpG/AampFORpbwiRCtg/X4iBqX
2nJagx3yDkyB3PnBPRJgOe83ktTDa5K7SPIo1Lu22CEOmOd/9TR7AT5K0Q1lRng3NAVMdr4ekIrJ
d/qWTSyfH+CcTErvI/MM2eLdkpWF4IL+Ezn5WaBwcSd19WL7DXD7ejvSCaFgC5O34EIwmfcE6gHv
uWfPNM6CTCQDf1f8Jmh+cXNlKzWWSWLrsiUmvnhwWV7AUB1YIo6hMWme6lEjrrA8wQtqeq8SiZIX
Hjbw4EPrV82D1zQ38Yv2CIUvx0f+N6pBzC1azrhLkJtP7AbDiz15tGhvIE8ieccEWBd98ZDIl9IP
KmD0TdDYjO9PykplC4WavGaNccKsFJeY6AtynQY+7YK0/W2dTTAHqy6cupZO661by7ezncYYYbRG
lgtFcWWqTC6wPjZJxAcW/lhuY/7Gzmu9cKjwZKnVjCyi9TaTi4rQccvMKvmIl4xrb8UNtpZLOSTZ
SKMV2541GeXVwsj9XBfP0ohFivZQQsWJ0cmIHfwuceWjjz3utbCUSKJP9zYIhTNMUYQrf2Ca9t7i
VKHssKE8yuBIy+ApS6Zt1lBx27fMtjX16rQZ4D31ya97DvR6pMrvFp20U2W8Wh3LO8oppkBGtvtd
1p5YE/gJoRniOP6AsmiB/c/8hFSNMUa/xrR9YM9qXNRXpWOIv2DPgtLr8L0GSQEcIF1cUmfeq80O
3lSNy1K30YCXK1QmEZaX5doiUrn4iJMmPYgzlAH+HOfGfMs6HUuFaLgPH4BcriT/axFUG/YbhB4Y
2oTl9+5n7GcmOQTHqSZCOXpRxZJnV8huy9uRsbBGIDSwZZJvg18SqWtLezGG/M7EFB0Ok5GClF6b
30JkhaOJ2z0rNYEXQ0d9fJlMdntvCfpAr/pvuO+hQkHLZWNUkbFKkCYvvqKCWxywGieyUQqNrkMS
ljP0dI6h6LbDxocy9M3/G+Sq9+7x7yUxH3yxAC46W48eOF5SOsrT9pS3WoYnAYlm/wj8vRxSKA1R
J2/BX6g/PQURcHghdID3UCdDXMqLn/XkN6DiRAGVUoVluDggJP9LyVlaHWpQ5haX7DF/u57SdQZ1
4WvxU/QashxqkU81dWO2rB2bq+UbCmQ6iTnu0GpLhMZew9vV1ty2jkIGBgsoOcAVE4UsoIIZkHEj
uA/IBBtrs26tXNa99UMoulJgFa87EQaxhfz6ufZI7lc4bwwrwUt1wCeNjQ1bUqKHyMceNeppHhpU
IhGmnx8p0TZoh/RNFFVownNZ1tlM/cNTCFVAqhgtl/LnIEfoN1WAkAI4OxdUx+DzNtuLqlgep2x0
/ssn/w1mA8IpKcEz2Pzy8jgLXz8nc1LSKEE9Tg0H9rOWRPbmwAP6/gDo0vyn0uLO0sYQ8C+U7hAK
VWX/UdGro3CUQPV1pRt37KxYUN/0Ov8EmDbXbxm9G2xZ8flcIWVGm9gz0OFb6uB1EC3Ik+hNhUFG
vXxOtKl4C2P2lgxlWb5ftamc+xa2l+ZiwZAaMBE2gGCp0IQnJYs1b91IXF4nb/L9StBHJ6wPHhjV
pc8z31F7GNmIRcnRUY/c5iMOVsKd78ukI38vtfv2HT1GHSij+RvKM3wlQW2Y4p/xdubNQ5qooav7
nbp0qy7e9TL50TJXU7Y7XQEBCyvvVa6QXAavqPwPtPu0Y+HfIFfMsgDPrLCeI1KoLpPpBu91Bl5b
CX8LQ7i/FOKZBu2xjGU9rkbB/tXcdNSAGxGmZuPv2e7iHXe4J0+8/0d6njSbzVIwz7bzHBQqjMzm
gkqcNqsCTt67TpzmAg4wK2MJUQEboffeAK+gXtUzZQ7qkrwkjXtgJUTf2IkA+oVah5yaOXQB0WYr
5wJ8toqYQj+mpJY1Nhiw2R7jd0GjxafetXTh6bsTmMWnXExPLUHTMkaKdSQ832UcBD78RS2P6z+T
Rtx1g3+7iMcRcVfxbuDdoMN7ly23g0MhIIF2MPO61lT+OEObWjkmRxcGOy5sW6UGOA/u84+K2sbL
TSQOn9s1MU9hyscRvyzVDFHndy5EjU03WWaRzYlLRPm505zCZewm9J2jB9rcTC+CNNylBd+vu29K
HieoI99LbD/Pz14E0hM9ppksDix0Z+zHBLBdTN5x9ZLaYNyelJIZXfwlTAi7JC2X8aEdlnjKYlcP
JJGhStnyWljhoyWBcGC/2KpUPqpWSv/R/LKkSPPeyYeXwi2M6QG+PYa5ZAIhyP2b9TXGGwTTG59c
XRyg7i1/hyXr4ZrM0A2wKI8rdGeAI1lkdsneIOJXWArJsUXrrdAjsxCAJdGgUQdmicUpYiP54Xyr
dehXMv9Pmftzu2J20MX+96fRfbdNm4wJ1iwbhCz28iskmpR1mz3JS0dolGXvKdw1PVSkat38lifC
OTomANtZTR9xKS6J1JRKpPGovxhqqYCqZlP3FrhwfF0I21oltDGnxiNPIzrIPiADhWcrJaBN+7Um
TKDcEQrTQWfnU+VdrAIgDg5+Zm4aGOa6qZiALwmfMJZE2vfI5nMzN/OBKOVVtC6qx0gqzbXGghXX
XypBWJ/G5PClGQY3q2uNtmIh9cbKXWfAwb436+y8gjIzmDfR48R6HbsbIYG9K0zCOgVZnqnziiUn
Jit9IRt+bVawRddAJVbN+OFpFiz53oFCPI5UUbtmOerVwVt8VLkif9dYJD8dHdWgV0AN7VQLdT+b
K87dz8WeakVB7wog+uaqsjMk3PCLtajxHU098Kf1bJ8cErb5Dd4J6nWkBfLTYgowJDc5qMk28BAY
afx3hhbu3PL816YHpn0CWjliFsHf9vNIOYKZn3ABR0QYn9F2piw7INs2bRTjOGR8LJxija9/NhPb
Wgq9gJ5y9vtk6S/AamF9IDd9n9nets9Bb+Irdk2obIK0IORBemnIlNeR6k60y9+zEWLFI52gIF6x
5inAm1mr08OldIH9hmfcKzAQhVzX0SbGFw4+r4oO/pLKwguKiiexId3j3BZ47gTx9WhTrbr5KQP0
sbDKgX5dtq4W+jI9B9jxivg648RF+xdKB8Newvh9CGF3FWfQ7rVuCBRY1DTx+51ICkIx7DKmssj9
7qWTGLAJWTWmqO/Nh435XycyFKDqlIilvZdIVUNPkolE8vXBZqXUQbGnvjapqf6asRzpH/lhApf5
7bOtMgu/07+E3dRlGQhmvJ/yQu9OemxdMb7VAvQWIFXJmXuu4kADBQLPFqnj3JBaXV5fTVGNYvYc
jY7141Msgbz1DCDk96yoT+OjiQ86M8WdhMrdPK0hBorHFevNv9EhCxcqLuIevOSQEMvUupXnMb8+
s6QokeCNIMjosv7ubzv3JKKRW07RXtJDL5VDvCDOXvVRW3qaeLipbo1bbGIVzfsulKJyz4EFuD8V
JMG9cjX6PDOcZapFy+ugGYbqmwTeuTPlm1RQiKdFP0ORyUTDmCFNpKP3qIwFQKATHN+ltTzk16wB
Zr187ZNGN+vOl1cTFu5oW05VfUZ44bU/iAf6cwj4JiD2fq+GD/Y4a6joRdFBiE8BrQ6Kj5DEvmW9
pNcZIXSF3q0z1rBLa2WEeO3fRIETfpxdjw3sPFapBayHThAtWDPSKpUXiYdNPrMh7hGVtYjSx+tV
bSc22H22cZECEKtRwVlj+X8g/PgpWRTw/9Pp+5J94FI/tLZDFGKNmgfBB+3/J8bFfu0t0h74nv41
RtBlF+myVyx81E+AAVj08HSbkkHqtdYNlPQ+lTCmWMYFucXmk04XkNoiPAtpIRwtJ0fgFWTwAvlI
p0C+9BIR4pkzzhelMhirq80xWr0JPQfIjeQLE5fG9en82V8qgvBCh9LUtDLEgkgvnTdEa0DfPCz5
64H+lLRPrCaftX5LgNtegDxfeVbokWJ8saHgtBugwVRBhysqh7IPYatCuS9D+bHlrH+NDvOIa8z4
qKqkW3COjuiZGK7Q9r++FKqlGguK5ukrpRbGhspQLKwsHZIc2Ps4GCK52B9hY9ckQ322yN6d28Sz
imk37XljubmZjaK2LiWWssnSQDNSQm1iYvzLACN62GSdrsaog2tAKt17JuDeizfJXc3vHnyVdOXv
ldZ9f+7UZicZKtzfyQLZ1uUBkQuiyOlLK7UlSeESVKj0G+RIuGN9zD9SKtrV0W2ZwZpVWWPf7MGF
6Pa3JBk3XIXU4IM6gRxr6luUuOfk7TBWIQVKqYXQKxMK+4ClJP6piJe+T5P8XVFhVC8HushUWM0K
x5pHTNkP+a3Cf+jOgfGbvrZGloptAWcw0Phi62F7JZKs1CkuEd50qMh3wxIfNK6NX3H3fC3CGjD6
sUxF9916dAwD7kWkRaVLkGSZAi9sbIU22Gf8FMJQBPdgf9/xYGXpz9xqk1tZL414FANtFhlar+po
iKm0ZgXfKPFx3m2Fl2pjrno6IbJKLRG2ALG/eYVbl/1IghINhCAWgVaB3SAEnbcXqEJue3jYL/Ib
fwex4v4KUJf22MHa1uyAdYTahMhJl7JyAGpR79HnxazAktMqkKnL2cNyCmL6M03PVyRrOhITGf89
rnCSrKm4DtGJtiqPCEoH8HIRFY2VxzERo1PKK2eWZtG9aafpInuZ0ZscpIgbg79zN/redwNrUQie
zVGEXVw9/jI8B7IID6cozT4UdD4O4m3O6/ORyvxYUeWaaBJAnzqa3YZnxuVN3GZHiieY89ZIWfeH
9Zts910sVyFMn+r1kCsYUboGEjKx9On0di2H00Rogxww6gS9keMkU1EQOPCHGDpcGt++8BoIFPrn
76UpNXaCaJ3VXd9wluaCaNAYkIMSsCsPoSoAEcOdG3/p5+LiHLQEJCkguhrPGKlAd4O6DRHFJZXf
3zb77I3RFJJzQOr9hrTrfYorT1MWui9KTlbJtonBC2YWH7TFlgXylidw6FJgn6c8oRW0CNxv2dc5
tDvaMAlNv6lexarLNYBnpoF/3hJYn2vZ7vkJ/MyqOIdgaPSP+lOqvUELl1YvrNQujoNGO5HQ7tWE
5bSZDpkDgK4TnQ3CyUU8EegVXiueM+nM+T10WgcZu1NzUzOySJn+sP/vn7zmTEkjAGCfw6bv0+QS
2Auzg95EPP0Up3KW7OsyzckZh6xdKv1bwSQrd6bMf5w8u5O7h2chhwPR2pHqJ2aOAfrfTfGd2t63
7QZOkWq2ZsIQufsj+Jx8PCRoLBM446zgeatQZVpR7RfkRll5Jd42k9yjjfrkX099iHh5Fk0JujXh
Drh+59KudpdScungHQ2Vf7FH1hZ9ITyIavzDqePvhXCFx1MFObrT1iHA7R0Z6UNL+0lC3HWsahTz
/JGPhZz0yu8+8gF6/f0/50emHR4CozSkFcLJWhhl09pjlSsNHk98jslgX8kk9Q8Sa2sqQIDdWj60
qOxPjJyukRWUEXBFyvIsKpGq4Ms5yZ4NbxYa2H+blhE2NNlwQbRFdvSyCuvwGkzQOWs+Q0zS1msm
YzK6ORyypjGyv7aFToQbizBUcF0WIrKuch8fUo1G4UA9NzadoW8pL6xewLQzJQE8DWCBdIKDzxRS
yDZczjQ/ALCKsZJ7likV6tyYmf/Er45hUkwib9HCBqlLZhV4cJHmxxbxGodpO5IpwB2bDEqOew3W
HflGgwaL3icp4lOJyuuDTZ97cU5IeWi6ZdVxHIyjtKdhW4ZyLbW5tKA3Q1zvN9rTeaEFEXwqonPu
RZeePwe5hl9y/flKpUAs2ufV7LilyIXS+K1k6o0F71IiS5XyYLPOFSvZdbYzp3mDEfbfI+bKeFt5
uCBLgiDY0AWmJzc3e9SxkB7FO2ZV8dV37UfUBdWJrydJ81Hh/+p1+TsofXnQ+36lNc30QEN3P2Mr
xoIkJuH5/U976zK+GEJwbJ6/OzEE3Br4KaogJypLTvAcWXJDio1d7SSn/vUm6CsE94CCW0AMQigW
BTT/lzcF/702aJbJSLbSATo6xoKC9UNBbJpAyFTxmWWQxYO6Qe/csOkedo93g9vc5KAAYiLvZJEw
roaM31Q+XHcQB91Nli+oO3DddgQIoPSRRXPfMYkgHwPezGwNl4m1wYZErhhGxprdRF2lXtpVrEDN
ghrLp3kACkN5yuJIQ7Wn5JvHOLsAg3/fa/qBkGmGeN1cX2YDnxS61Q0cBcnys1i3dh3R4ezAAwFm
9Eir929Neum1i/5rNJ6JJym05YywnLrFD1y5LwjjsF8jJZApSvAZdsla6sgMMVkQ05gtnmr9aJTH
VUarXfog9iqapXd/l4U374C0D+k+cJlRPLyOgxslLX8LrkAahxmJluRu5O9qqssK2w8HIPhG1jVg
OnLOlfBqyOe1FD3ElQ2r+OdPp+McZdOiMajuNC777f1OAN4iP6ECNTTChwnVaLnRuPViFKua+tH/
Gzw0naOig6gq6lpQ4j0ucPmH2rmxSogOWLVcvqkMRt0zu/bSKNjFtN6mEeFV90SfJ34Hm6DKQSww
IyzoL4sFERRwWxby8wfV755WVQ8xl9cLXMAGDKUIdM4v+wVQtCRq494/o94+Eu4MvOOsr/MuX5G+
Da3SFYkCHpKAJh5gQvIgwQNGIp2t0o6y8prQbmdt6lnepETh1OsQvFPDvFzXvVEUBobbluONF+vZ
6OLlbH++O4cN12qb/csSHlzNuug1r3NdroZFUhkfCxKjT9qpLLaVxm3je2QIcJqsI8uIWAmlW4Uo
BPbSHgRbMhcdlgTipVLBAXZuzWnROSNDaNKpdAmDS2G8xVRXvnvyYFh+oBOXOCdJ1PMklAwAcogt
5YDCoCdsn/lJKwy3u/MtdRH4y4O9at6DQVY2TOrsCk40qQXboxsKjNVf6K/EN9nvUNzzkF4C+vUP
yEPbxx0Lhtr7p7m/0Jt862M6QYxEbKX5z6ZOJXgqycj7CvW6KiZUfpLW9Rsvp5lNLQL0eIR1tBxO
X7qVJGs7+ifWe+Jc3+S+ac1k78QBZQV4OzBZ2VP5SHpXW1wyYdKuZb3QBH17/WYdlkZaDJw2zACC
+2NWt9RmX4fXtnrbk8wJ5lrZT9dA2qeWJ2NVy7fPCjE0DPcqTyE8AhtH5oeTWbKbbzKfSJGOQUFc
wSVn8qpTzQaRlYPyfk306b7nmiGCbize2uFgUpEplA8mwaq7IAaGKaHqPCppygAZSmLaFIKTJUSz
BDoT+kpoZFesVhllCUwQWMij6FB/sr7HuOzx0d1jv5AgfMKAW8bOBLUik111FX8ietE36mX19c2l
slA0cScGn7/uHw9FOjGemtpvOKnQIcGLwhWuLIXJPdZRrZWUMYc7dcxM5F/cd/gxMbYNU5r7cwT7
MWw6zwsVbQBfJL890pfCRd3XA3CCWML/qPWNjzRJpC+M1z+rRZ/8vrJx+n0AsTHMSNnZhKG7kf5l
2IXcZGu2hgdx16AKkRzFY+MF9PDyrJBhUqXv0Df9fA3ovOnVdACZChzAV4t5An/Ho8Kllm9d2PfA
p/DbtjhXIZUP3rgQqfbejxplDfBihGgVQTsrncdRPe+3DdlffsnkN210j8DzK1ad0kMgx0dSxr0n
EcSVFyPVUcB1eWqMj26QQ6IjdO7LVnJ4nlyQlP02M5d8xwubHl9ndl4tEDl8RHr8uXedgNO7HRvq
/QhC47aftzceDB5B78aLMY6QcBFF74CIcJ19sJ2BSwYswK02vPRYt9VAHJIvr3NozPS2Av1gCmim
dYrOrp0681J4TOpNs/6rTSUzHanPfyVjUfTt7P01MPSxW+YEImgpp03y2cv0svvBLpAGdbt4thD3
FnwLu/GJsflIf46K7vrjyvtXH6Uyc/DmuvQPQbdW7lEB+NQbClCs+UKOmxhMgd5yDoHWHNF/18TX
xHbZ7HXKuNx3rg5hma0dFDC0ur11N5841iHvP5GByB7lqSAEJcKnkQkVJd1Sx29wQDNrXRNSqbQf
G4P2IqISlA970uhpKqoZpA1D+dC1SoyGR5+L4qTFl8x4jsUJr8SGRKT4tS3D7UO7m04364s6STnD
u3vgvkw7xBkfGK5N+4+p+B+/ROJRlTE3o8zw5yt3HdX28i9pt6F3IfdVV1HhULrQY4u5sci6FyCP
kfL+Y0YSpaJ5zav7UfLLOVgCTo7tE4EKO6mtW0O1y1B5uJs9J107eMEWexaKzostSUimoZyCyB6K
reg7Wl9XR4riu2ue9EvVg5wgsOCbLf+0uPruaug1C2ZV/2+jhc9QtYjquRdPWtfeLu+YCVRZ4tO7
4bbDovvUupSCnr59Lle8aGAGD+rzZ4OVfWEo9PwBVTawv+RlMhIhTm3U1mW0jq0xAml8S5ftVYgJ
LWOlHU2h/AnuJRB20cQOz7WYb5wIAGh+6eN/LT841jukoC5XHE5HkdZzGDsTS261PROSL8iLfEnq
2h+xwPtgLX09SrGMVuqQyfz4JoTX5Lm+6ReIqJ3fg6eTs6nTwhUkrUGIhTD8pX69K1iqM8Gd10TC
0yX1Vf4oVmgdu4WjQy1lJAqow/gRLPWt/NOBwxrcioAVTfAB/GILjmLuIg5QN5MZiicCFMkxu2it
Xi0ir16ntgO6DwnLV9v+BM9eCNCewikZiCpY+cvboVJMR5kKQZuB0lCDoEapf425SKLGatzxL6Un
ptqAmfB4sUcZsJ++KvpdIGbn1zg1KCsrKJ77DssG+6xQGKQBwu8mT4bdVgtAsFJTB5g1S5nL7vj9
hInLbylwAKgHjPUj8Uulqm7h1HTqQI+oVN3DaV3FNvejHKMQpRj+gBUPWkn7hlfW3SzOehst5Cdi
jurA5EDCDCkGAROc4eOcJKLT4sYL7hwgBkdsbFq8M0fr/wYVDe5m3oHTv0yxGe99WvgO/C1Dw1r/
WLBTFcFPW+QY8qq2ExOVVuq8xOEZaIJtBJ5PxSpPKTib/8Ux3Nl+uCMJCJ5Mkg1bDVL63mxlUnvZ
g8xxAdTsbqiGk4JMtXpDbsort9z+CeSTMl+Gri0NBDRpO+9UVY4NahjeDoo5OxSIiABOyEeW5O2k
S6ePpY0kRu3eQNMhfoqg8hC5uZ1JprPPyH2EZcIVMmgjjCwnwOMWdBq22voP+vgNxWcNfbWiCnuJ
gbPQdCQ4B1usk9qMisnE2rtoLo2htIgyXU3g7tOsOcHkLvEcDKtI02146uqeHjdLgegqLYpWsWxr
2NLE57oDKicPWLKr02y50Pi/i6hVDC72HWBfKzVoxfWjWNwqmZ18aXxlkXwGlULSyS7t7FlQTGhN
SIky1rF2eYxloXyJ6QhG1kEtjOgSstZlDqhripemTTsKrXolqebE0PATOFZqdAgnBOz2fTWs8OE3
WzpyeRpvJYToGl1LMoj5tUrIRubCcPJTewo0HnFLikc50esQB9IdBbM7Ir6n8IHYHUjSyUzUI9uB
HJkga5TggIFbYKcb0vMpy/kzIi3/Ezjm7Ve6IuYtaqmp8aMCYOcd/aSB5JrQzz4EopE2H12MObuE
9RdHtYgw22UMwLxCKRbwOnuvQJkfpmet2qjePmTFz/01SXWbD6iEckBTIVRLrvaJM6sXxW1JQC3U
UlZFhKJfyprgtEUjEG/5ciEP+3HXR1FyXHEIonrDlYcn3XubQM0Mc3y6TgZO/fzUakaMRHayVoBd
O8TJEWwwlWxiW61RyHc9TpUeKCXxD/7T5h6sKQijIApYVTTbqlcjHIvTec3SA1Sj9fGexs4fh4bE
C0LYnEhtygqR90XenNcQCU+PW056XfcvWXIlSo6blnOgklHapwIrM4MT2KEBphZfMAYWp7VyFhLt
VYXw+2cW6VFzaqY6e2eRaGtsB5v4HWG7p+0AG470azLJsr5hCTU/4Tx2tK1rP+inAheGpJQWvqZ4
mpX6ug0dvPAr5OQpmJYTdQ1rh4jJT1crVCsWzyPZzt/fiAFz1d/ttoE6xu5liO4XCSuDkDty35Pd
qomqeN0KL13UUlOgy+UsuCCXh7jwsGuqoq2gfsdclbXtNsRkuf/mxchvCZ6opDQYgyvu35teC9Ec
46EilHQfTVMmH/IXlAp+rcY2Vm+AUwTF11cs+Tna2vQT3pacihj2YO2gAIWG2qODbC00IndRpN7g
8+LT2gl/FyWq/PllmNow09oqmVKMd1DO3FHtfSN4aNCvkplfghBmTWIrE166VU3SVg/hqpgvsO9P
juqk/U/FA3d0fI6Rr2+HfzP7hq2fCcc2DgecDaxWkcc/lNU3pm/dHH+T1WAR+bXEkAdcKccjFfCR
M8kkLE1YVizz7PX/OCotopCDH9VTaU+qfRucvd63raDgWmCxcri3LJnFmpSpIskrzlME1Xo4FiRX
1IdE2aoU4CsnH+G7GgpwcZHxLmQQN4kkxnBLchctba6NSHiyD+wMzMIHGbZfMYjcFx/PnEtsaald
ibUlh9EvElryOOaQ7oTZeVF9wRkONRytx2SVzGIrPn21Jw7dJe9hBbKm1CscV/F+zQ406OQpvTJ2
fFN8qbeaobXwbaOEEEBV8hGwcv8YvqnEtzlhBqkHsqT7gImARRxsLdA2rHno6ddzXHmEgtJDdQVZ
UDURnUekfDWBJ8K9sMWJXr5n3L0qPI6Y2y/c4HRWvBKG2mazcu2HjPz27lDnHdIWqyviEnpIPUDb
fIGPtFm+1x7bCMCjt0gl4FMZ0mFXCJJByKhL06eDZ4IP3V07bkxH4Ct2aEKCdBwT843k1ZYrNUtr
mUYUAotZVg7WVYg1GjqnpnJ3jN2hwyYLY4scu8TrH5jbV3bd8mEdXDCiQoYSs7siqFTmG2O+ul84
xIr2LVdD3+KN2jLrOx5ckEH08DdlvVS3WTLdF3v9gJUhHv6yrpQo6n1hxi9rn921Bc8g3iGx3Va/
pOMSQZqV2EMNElcvwYnCbsFCNmxZ5rrqJk1eF0FZpM4GOlESJn1MAXJMaW0YJRlq7isH35VlGS6t
2XP65dWx9+0HgCX82piOswsKvTz/i8QNDP70r3n9w5NgQH2KP97d5lvsqmIuvelkjFoyDc1TknEU
K0WvLzKVL9Oaj1BVb5z8WiJ8s46nh5Q580essnhTdlzePqRYe0RkML88meZ+D5DDYR87O4+O4Ztd
TGgFW6EJNY6jHrO3SPAo4ja93W5/1RyGlmfJg6QFwRLrs3U/v/2rKDy78ftCO0hx5vXcCqY7AYpc
rI1Emcliqzyjm9coIBOe/Xx+VFugY5P5lrosfuukqZb4vu/JhpfPOoLK+7/t1OOx5m2vlDhs4Ic8
lsLlZ2rKKf0+vEDy7BqiTIecHcSJlvg4klm/1++18Hz5gH6HOdgkxuVW1IuovDJyi1xKd/Pbaw8I
wRRNTxMjcCmCm0YvGr2kusPGTfN+0F6m8IUVqg99cvXqVGGqdv9bWeE1ztVRD8vdMhLUFnS3l79+
ceJHXrElXB8vfA+HqWoIIaPYVvdFOKfkKaymmVddnYRx7hKWsbwFwkspL7RLPiO/SgaQLFZ+xLy/
DXRsWzpGe3yO6k828MljMvwMdOj6+twloHI48Po4KjAjMRoRUvA6kSrk1aHEYkyNP1YIxm1dPF8P
yTnPZbV1KEJO0z+jl09hHWpo5zXeu+5eW2ks3odwUMwJvtVM/s8gN4w8ZGvpdto3cmOaY3E9T75v
QEIFM08YSjyliabKhOprb22dOFAKM2IEnt9TRP3PXa7gPlAGpgwSQFQMvNr7iKg/MNX8WYArXFZf
NMCk3KEqLacnspKeT8pVRm0Sow0JWfK64rIPapzV/JmKr5MV9LFrJxLze9Zw9UaaDlf0dma6n7oZ
hEPnW4stsIEdYOoZl4GFie98G1S1RyoRtZHz31cqyhg7HOUkZj2onuQcxr2Y0vkkZiiP3utiobvp
tnf+CmgoW9Iku2pOpY6BGBmRxln6Oa7BPf6RQaW67a1kJPfplk0qFIeJukiQIYtkLBA13IRtvciL
iqDuqTFg8OybEOBU6ZP35XXJd3/wo1nMnFzsETZOQaZt5WDpOWUr0w3zTV0BQXvjjTi7qLhEpvqD
W3ppUDbieWclU6JtVikSzBwMndrULV6Xvvoh0VpucH2IVkd2vpTuKkYOIGL0eazpb5dL7nVKKQl5
BEVvE5CcFwq7S0bOx6xRD/lWl4gSvtxtl8vSgTtiNSz0BRuivOQ9iVA47OGZqAYFgBFcGJ8PqR12
MBtpk6dXEskivNlLzm1rhb2rZgBBOmKPBR+VIyXgfQYdbn4+ebipD7opY8+jpfmu8iI8QCDvVG0k
viwQBL7R1ijeY7NRTf803wZ5l2zFIHR9Ns1o8c4xlC99NdTIM6MiV3PdWHaDRXxJAMRpH7Ogfovc
Vzz3OB59RQPkg2whPdsfNgs9g4n0Naez9b1pAUxU4Ymo7H6zo0kN6G+cT4zwrRuzIGcxD6ZOxOIb
Z9AmGRCU3BDMdSmFDwA4ISnU1IrzawFqNA9bp/70FQz968sY+5hW2Nlxo/5L9uXF8wFsnpNmpaii
qJx1Gd9Wz4jkwQkJo6ie87zK31KdYmKmXWjSuydL4QBBtJCuRozO26xEUfUkeomAleQ2/nWnGbin
jxBmNU3hTbM1M8iksNbFqjh6sIlbyN5K+DlPVas9qUMjxv6D3JuE7YymdpibICp10aMQ06NBUYzl
n1AsOGr33TEZAwzqnkEJsVxYaEH3AVWmvMe+So6zPEqMj3T1rfeV/Ocl/qEcwQkJv7Ym9aUVmrmx
TBsp5KjuYx+ED7sosKKA7LWTDB23MrK3Q4UX0OvIdYtWf2GbPTE+w1iYMpaNJnD56wsZFo+MeZM0
+mGGUiSs/6wvp/6/MYiBI+r7KCvYBlccyJ14AiMfN7LtbQwYEur9fApwQEhPlGWg+vulr4oH3nbr
cEwJg6Dy5sQIDXKspuXXNDSrBeH3GR/seOctBcDTFD18pN8KcmsQp5QgpOFX0zbiJ/4p06Ey9mal
xfzJwBQOrCW6MVN+cKsubSOR3VZ3pOKJBkl0HW5uqrbGBXvtfL3uXZSlmkyS57VtHVZGxN98F9oX
RbDsSz86t+2wtn8x9YSxrnyInGznvhNbsxIEf7YqXJQZ/18NmbUyDfDTnX9+j615M5bY1lkv6uHK
hEKb7xfsvhsfd6yqlxm2uNfLJZH5K18bkZitK50TKa2DahkOuJQLy2WqG3rNYPKwlZvTgQx9FkSf
3cxA+IYY/1ppiRm5xf0QAF3lreucZekZmNd63FCGRAVQB5v2CO2PlZqYQYK5jgsoHZLZUY2rbeMM
1/+RHj5RWboGBg+TMjRvyTmmBc37mbhw1uQk+09Z2BUDnXbxZ4fhtp3VaBUkRkzPtgN/UMB+L++y
gDWm1nNksyvXdW5wZUXg57HCVfkDL5//y753KCowNI7miakO06ugwytfSf9w3vto+TQq19QmHXj4
pSxn/vNHBZ1Ao4HydDOPNBI8m7CKw8wpFl5BtrNDIrueT0pWo6ZEQFJkb9JEzdmt9ymwUuhMQgaj
j/WQbsTRDj6t2qq+uqZxVSw3a7P4iCom33GAZDpawd/wh8rbdkDMfs+V6WA2MWIuLA1pkTvmL9nc
DoJ1a+TqDd2CfjcB/4Mwlq+ZDV54C/CIJbZ+khxdcHKunSkVSYV3ezblLHCcprbSl+Ffu2glPqYH
2ObVu+Zse0m7k5uipDEq3dhvnUItMld/59/J99tYR2Emxyl3HVOI+JGd3WVUFqUtH7Naroqyh9+v
AiyimLEKLIdK1GHFk72dgbKXThh/rQnFTxyWTne12e7zgyqa5FTiDLbiQRVzGnjWd0LkPvGhKQDa
6vb6lSRldp0L74iJOsxINCjG1t54nea6FjMAqojN8kfCdJv1LwRbt7R8WUoUDx9BeZo8L5PFgdIO
LsGSIy4yGrkPq5BNZlZAOQ2V8HB1qPiBo5701FioGGHd6F+IG8Dg60FE50UHiGqy/t3PNYGrLX7d
4Orc0J84zRiy/1nUl+MSUc/DkxXdsmjLCisoR1vsQUfb7VHnkBCx7YJDhJBetHp3mqyld35SVExq
Q5lewbVYSuRjGb/MtuGdjh0aHsYXkeLMYDHMgDZcM3zAciuvFTypErxU/qRSL7ifUlU330PmdaI2
s1sR8XbfeF6pFsxDB7E9Bjdy28ezj8VAJDFAkEWVSJrmN2FsPO/8R7WyL0/UNWYLaNtAxz8F2ICD
52ab3wKS75VO5FUHUK7tbVIY4eQLhYg4yugKuw8YnFKheJrYjVrFDZcpEVbewoOFUbtzT/pL6XwD
SqYGdLNcog9rUssB3w5fgNgcuDwCkl9dNHhp2vEJ13E09WjmLDUDL+8+MxYf6gm7bNIrwtWkn7oi
XAbx6e0+GNa+FNeCOArpzU6Z7hIODbEQ3d27UYHEBMxoxRYIKrKId+VAW+Ms9qmgzL2hjG7Znhfz
hmpXgDXbENb3MfjkHmGi7ndDbBK7SfJzAOhEezcbO8ZNEZpSTstccu6NPIOr51QUPb8P0g/wxABs
23Bo5KHvazTdUYXOrW9JqDDxa8Hewno7haoHcBH59Y2aHW/OxHvh6xJnJzF9N4qs5xdNTevWofTZ
mnJsyBIFE4+jTNNqqpHRtD41VCOFjflT/LpLEpHKRV0yjdNlLTVZ6BWdhHiZcE2lFIHmEF+QfsEV
O0Sm8xZtP6zg69tMqAWUQ+pKxX8x27gKE1nRDnDgmZIoyqmNBcP3gK/9TyrhUL3g207092T9ojKP
SHSFt9am0z1ObGgHHXea3r4btQmzAx1kaE13WbhzpBLr7CE5D8K5P4Ta1n7xL1zkS76ZSa2WoYIC
+MQC/TS1IJ8qd4ajxM3H9u8peAU4us+xy6t1THMQsDnZRz17I4Abg0PZ7hrCDzm9ZbVUMFTzj5Lv
0WhD0BzyDQp79IgfaKYaKZEm366ZPDEx6oU6WoJAOoXwiVJx53WA/52cuTUBLnnkNvtXodE35N/s
3SoIb3fHvF7/RO4yXS1+BdLrOQ5uCqQ7Rdl0KGvOembbpE9Z79yXgpkLM3EYCRkNGuuRDjGyBLAZ
84M8o2R93mSxgn+56XIjC0ypmZBHRb9+03osl/PioQZuGpYNOZmmZ61LJQkbCoLGval+KecBZ7a5
0kmUo33Zyb/W6BupVAE+cDx8eYJDxwI1PSIhW3gQDHYqBpg2GJODvRqwHauzozGJc0AbzyO8bupp
sKhJ91Mh5Jhk8QnyNAvyJD/BHroGwfb+45NGd3FD/mp3KennFoVXY1z6BJs8Kh7uM/CdBZq2Tg5x
GvF3H8V0Q83CkWQZb9bBfhqvvN+FXRJsvC014ZzkNlyZPzI2Cn33iIuCdlF/xDurY1UWjIGTY14F
dC1nODUHeEXXxHNAtK+47ZVR6f7Mrxq785GbScSvMwRRCNfZHV8iX4no3bR48kcmxBMWZBXKiMtl
QusJ9JCHfFKs/DogMp2JhKW2EOO7tYNdbSdozeRP62Lfc2rIKzoUFo3fPGyCwfUrJCalBRIQAgMl
rPtp4U6nb1gLV9cEpxczdUurnb7fhZmRp/MyinTJ0mO3MOsxek7Jdu7xgqRbXRNc5gWpRTBfagHK
3qzDdmykVq44UoAuK5M/WnOZFCfsdJBuk+9Ew3K8QebEWdQo+aA58Ep+3CpyH2SaWBcg88el/uuY
vPBs2Z+nX3HytspO1ejWzqzQ8+zPU5BgsA4gDFoDEzwwn9mue+yDAF+jGo5mS8kRhQW1lBrjyPRJ
A9PJ+nL24+09a5XuVj3rz4KD1LHDqt3BRAfPewybDKzUjidC9xffho7ET+KgHX7ryslVsyA6fBbi
TYUmkTfchDk26SGsBqJmsnyj3F6cgo4xSEuRg8bTKkFewAjksKGvIi331ZJdq9qDOUgrrdGGEaso
xRltWxLV/sQJR95hKCtyqm2AXtoCtIK+xAsTEm3RCJxqACOFlLgXLcIgVHZ3gwwW4uvpKNYnnTvW
01N7BLXyoFhmctlrqOqwT724TOCltejL4aaJOphkqGYuTNA6j0ygaF0DrCFRBCmKpEgnxgbuHuDg
bRBvj1zZWt6XKvzS/9Q1pBGzfMbaOBv7bjyIAWTg5fTUU39w7WxkooQbfOsDpA6XWc6DAXtYtO+S
BQkwRfKj6Z0qPBbFVrP2Qwd1psbInx/IYMJHtFj/SsjC+UbGoHTE5v0GxzyKyiaRf/seaTsWsvwa
w1cxV0+1sH8QcGZtiBrE84RT1Ut/89HPvjAfPZxVzV8WVWM8DWZ0ubghSLcnkFNW+693s8dXM1LH
uHMFe8MilkP5jz9qypDF6a+f55OmNCWVCvXsF23/g3mwXRgZUSP9fggBI9nEXm8kXLFLXomzOnGU
JPvh6ga+UdadmbWONjlEf6Vt1vpRYytyhJQkJjKs/wRR8sP8+tgf7NL6du6lZOzfOQ2wTMzy9z8H
Gq9k6JeGsPHZPyog1/jaewRJm7Xf7aQUH7ullPtAo0bMb78TADt8K+TZlpgY4xSe57MEMxu7mMBL
DVG/hHGbTIlVIR0a5nvTV/tOsNoN/KNBTjAQTzsLmBK1jEurLJJeJ9Mr5btEHdRiShnhrcWZBYHe
IZlwaApDxdLDOPe5n7iC6C3A+ISD9b/1oJWIMwqPbs8F7/My1zEUtPw4ec3k7bQO/Nl4pZzvyZIA
sq9yZk4+FQQlSJ9CrvzHfmWEfdQYhlL6PPH+9x+nkBvxOsNbn528Lp+NGu2+3hzNenzwQR10spXd
DvTecotAiPcEkkd/sR3fF7CmDJYtO3QMuUJ5BfUyUnJZ/97cHRdcIFv/F9RjTH7PQEiXvrdWegrd
UwKmXpoanVW+nWW/yx7blG9ztjAK2N2p7FCBR+HJaIFHkslu0NCm8oYhfShYohSNBPCsliUpChNX
I3BLMFeQVhHZsQocrrKLNfmOcAs00obP2mymbhqFrWf4uDFtpn90glYwhc1AglQBAfwKQLs5IOek
mfCzmO0RRxVnDpl0bYWvQNsJVazrjczFRDcb6dJcDH5LYiGDMm2QfSZciaZRnGlpI6LmV15Nz9fE
2bbcOskgdAn6Q7+yC5YoDfOK2VmtYfOlLSc4y5IC7koWpKCgiw79mRBG9eFSKbMm/Ui8eA4HA4lj
Xw2vGaKC6yAGUyT2Cx5XZ9IOIIxoBEozp3wylBTh/SsQIldVs/1yxR5WTLozog+qdIGZVdUw0UwU
IBW8KP5g0FqQZAZ7y1qnLsYy/kbP/HXDJPBWeO3IdhVwTZIAZnFKvkP5//Fbn2bQ/AeVW4VYofrO
ejJ4bdKz44zCVm5KsZhxi6JJzsFtrWHdqs5rcu8zNq4aJ8509yWAsilAD6yUWNUQfIkstN8BrTGk
WDuExcMBAfE+w/9TdVW7uzARSpOOcGvVVxxFfT9X3F94wmx8qWgHDpoMHM5FpAjV8j2sWWiZcNKh
pTzRz48q8PCivc8al1t9xL+/icjgbc08P/FXkARwmTn8ss4MeaDO5rdFkAQkc5V5yNcEI8i841P1
LLUihpgdCSguYktm0DuMWyabTtfGLVhu8qNgCTyHJNB7EWQkKwYYk8YdF1Gw/7QyyN9XEJbhLlPC
8MUYFkN1zo4OAzflIrR88fprF49KHr6GmtKimQ6DDzAtmobwFekZAYQqnaTFnz8z52RTNpjptCXP
9juKs0Umj3aSP8Eawo2NmqnuFU2ps+Sm15pMU3gUc/mqOIZXDIKNKSlvAj9hoSuMzZkont6LjijP
6LqLqeQcDSIgFSIuk7VcmGC68guwwFdkvheFbhQyheyAKiwnUvJJopCPwNQIVcUKPNf2gEkKkDQp
ziUt6tU8KFRHGwq/NE8Vj2XSk2lf+yeFlclL0+GKuMxJnXnyWbbg2auFd/bIXNWWlsjDNEDfjPvn
J3cAND8xCnqXU+TfV9GWpPuc6KAV1dTMWAP276rsnUF1PC743x1P+k602Oyj4HyWuxctu/Lnwb4M
xJr19tZ/HFKGtj2WIeeRJgm9B2ffT4yS9+htT2mCAIUq6oyes+tdPxFR7vkBa9PFeuXFqDEsYU5q
Btaizh5kbRpwJeb6k4n6zjGbovagPMBoirfz+8JljPXeG16C9W9DC6NJahfaYBh9N3WcYePYFQhD
3gjP2CsbFFfufTavZIjLsgT2ntcuQr+qjeGH8obeucNxx4w8vk6QWLTezjUrHejM94+/D+W09lqV
dxNMR/jB4iK51PmJQQUErNoTAl2rjZPmIBixUtg4iEm3+zctpiHdGPyfhSo+E7brhN3tKqyhoNzZ
bSLJcVcobgWkq5cCx0M89PjXtKYJqjQ9YzvsaPXUTYQGBzisTRAO7mqT5acVTNOHIMQDiJz/PFdF
gk3A/WhZBGjm9dHrnuiHOR8ZRIwId8A4r9UxD6/tGxu5zAUg18yXFJhXR+BOosCkVIhhb7VDRqO0
Gu4PXht0KPODezXY15PKLBBfxcVVSqVDAAc0dBH2ycCbT6U/rwdFfIApXCKx/x2Wzs4QQ0PEK8nU
BI69817lAwlOOjqXjIECQjnkRuA2y2CC8AxV6e3tR/ySIX4XjSLWp8GeybEvvHKHG2Prmk+4sdI3
R5X/b6PKflw7ovVVJWvUA02v5V+2cegPWo+aafcJXGTYFFjXTDX2JyhGZXqhJnFVg/b77KnZLT5l
vfVgcTFyomR0892XhF3r+EiKSr0ypH2Gi8QfVuKK3akJ3FLEKO44zueE6kI1aR6+oXw6kFbauQ5S
Y1/BT8SSoNnI21x63UKVaPwTlCc+atZzMJB5P8bnRr9W/Eq9Q42WkAeO1llvqTxBkGSQJrGV9+eE
0quGTF+cz/Pl8Rciv3+uSE2l6zuDIaoEOMW2M51R1SEslspP8n1tmfOWETzWuCZWOB3kst4VhdmR
LHKNcB6EEoFx+3OxGjwMOS8Ikt6NSGhCyupdyeofFZVnG1efgPwhxgei0oyMqlfRfNPkN/30yBho
wYFEL+UN16tMsQ3+RxsERlDF7wKHapcsYOLDZiTvNBob/jbBV0j+Dvk67gyGPf27OhzyYk3E9dMv
M+80yPMoHnVXPMJfIfhnqN3U9KzIRsKhsr3SmrQPoEtAsRwvfePCGDp4TlbizhkX2dKhSKQgTNrL
jyZoDvBL/WWmBMDYoHxQMtQ5IOI+EWEpmdH/JA8lbiF1GMTU6CXzi2bw9zsi/gClD20SpLaSC/9w
/59WSYK2oLfUVa1ZvQLhgYEFZn9igGtiVNgqwMJOX2Y7ZtQkrbWy6eV7o8frTmR5z21qRoFwcvxF
6Yz9Mbw434g8gcZG8Iyiuv+VsJ0+UgL8bF2djcQx8h0Fz9nFtjVmU+1THSxUA5CSjXHq7YqPjZt5
bMD0sdiEVtW+KElJhvkYwFuHlMbDPXyaouxbHOpwVTDxdCR8E6BDUln9GWkkWlt4BuaigFAKcQ03
IStOgV8jEEZ3CjP87ULptE8JrYSrafWWUSr1pY8ANLDaUc/XogpfAtkj/MoIcJOEOvcI5whxKRCv
/15YvKtqxr6OMOC9gY8fyprpVBKKIxrilX3htMnnE47FKAf4sK0A0yV/AdeB1OXNBGgQm4+5pnMW
zNXMkaWwzctmvILvNerZs4pZDVqOpmFso5bhz3CtBphNCpUfCUyc5fhQ64OX+5h9KuM4j+5hQ4C4
1U7G8D9FGLFzFVGq/XmBx8cNYmepv9m2c+dyMHfSRZ/9UsB8zcb+NY/UPNsoFSLTNQEZCgAp8ToR
4/lLxXgcIEeamPl38IuoCaevnE+RFkHL0F9AFw1gIzKGVpolTUCr39PQEILEqJn13ovH+poqgTOj
HNrRtOJJ8ojuv6bzYrrbr2UhuhqRFy0diOiFAg1UGGEhB+z0Xrb4OVYdeG++RSilJG03D6RkqNOA
n9K3h5uESTuGtvrVV7euMyjIeWmjqawxV0cehODmc3mwal+ymfPNEcF0T/EHpNsXL3ur1CC0mM+P
8C77VMTNVJDEORTPAI5WN4nbETrz+lmEKzcpYpq7tyXBpNqXEEzwZAEk8ecPpIiuxKjhfI8mOIM8
FOkWwREN5bp6UkuXmNa/4MuObaNs7WkMT6pFlh8rwBWg5kouDUTBZkZ9ne1nZtIwQe3wmRuP52FN
Yd0PpioPqf3DHdr0bZOXCszbpDKsZARIi2bz0sZ482y+STINIP+sJeBMm0UXA0ps9akHge7ozARP
Mq853qjkv3iIgF3V2Bwrsz4FOpWhLm1Naaue9ePFSzd+pvipp6J4ScPHAmNsFG5xkJwbFZHsF6P5
Dp2ZSRIhAFdTeAtjGh5uJ/OaTV4RF9e7Jfsu2sjauZqA2lFUFckc7taQSRa0zfm8T6T3R3IbE3od
qFjh7C4iaoQui9RHbSYUIXD8syuXsmoiL+CTEstRkB+ulShFFUxBvarQ8GWunoiQkw0XtINtEdo+
ISRpProM+9MabDF+CgXKfigFhhAoQroByxfL3uZ+qZgY+GXO5xFT6bMXOW3wpXnzvHvMMu6NIlHp
UgSgvWY7mVIcXwvtOHdDWkIEqnojMYRVAv2XMszFdkLzmKUkzfoWl/qpK2BMhxnZxDLXptl6SkdM
kzzpI3Gl6gV3kQliozCwo+RsaEhNLiv49rD+2KjOLCQoYhvKqI68wW/MpArBTE59lXFzXwpX5d8e
t7ZDJkF8ZVfUq8fAg0RnnWq5c5xUr5nyJfed5aLo4C10jJOoYEr8HtNJMxJp1htcQCrQCyG3ibQq
nrjbzPYozHUig5njvbSplYPiIuIKNbb1JBWJKGvCZg6ftBPK7HsBaB35K3nQjZwHXS4dLlFmfEkl
fbt/NXWlN+eFNxMVzM4Ej9/pqi1ny1Kw6frhhT3sMHNKKbEj/s++RZHDQy4h0FqAGPKMCEEMhQYO
sjzQdG4XC+/hSnFP/uEYc8Gbt4k07LIMPSM+rmwpHhctF7+DwHn2UWe/0/tgpQ6s2SW7iOEtugHm
43YY59h+j3+N0sM6Arop3SfVZmKcp1D9FvvCnaxCeaALiLnS/PkvD6IWwsOU3+ShyW0tImntZgUf
f7UxaQ6kTKO1GAN3jPAHDAs2VPL8d0AYNrhX99AlBVFNQ28+QpQDk3FxDQ8jXNVHlIFQ5E2kBg/N
3HAaLW54nU6eakD7gd5tiUw2qY2D455v0GMQb3/P1sduGJnMTsy2EP7N+Y6+vw8LpZ+CW8rd5gnM
v1GsMvKNePRMFkhefsDdAf6xbz5zXqmJcECl2CKWXYghMGbYBcJLlcPqdFSbXCNPg9qr9Gd7p+CI
aTpO1JMhGCUiWcosmx3R9hbatl0Z0qcmFxW0h3dJ+Liaqw1o64YfiGDAuAcgZy9krg/luq97I4oP
2DjY+mQ7EUgPMet7RcR5lqsAkOwuynoKDkA2eQaM2GOJYlVWpAMhSkKfA9HKI/mAkwZyIVSABTLq
Vc5ZzU/9RaQI3OadtTzvUarwYIAfcrLuzFnnr6HS+vkB7WEvr41GMbqGj4QLvfxS9+MLMp1GIa+D
5XnEHA/tiRkdQflmLdlVTaEXKOc/EpyQfCD6FGHobPqPDaHCIt+WMwVdhut589U4ZB8hlbthLsYe
TxIpJHt+yEQwlSqQ/vYx+aTfHnwleqB0MN8FQbLdwcwLrBNti8AKmJSjlwmnW7jN7wKXLQbpn0Zb
co8AqQnkaQEUjfKABz7BOKVZm4hEOKIiXAEyJPHC62BmwU4ZxUSVUuJFcPnd8zF4zSdGDgI937Qx
o4Mg/WfF8p2HHBtUnUYRbm9Sx7IS4Kp8/ShhIxWZMnV6FIs85jNlrrJjIMmIEEx7YYIdwKlTNcUf
vBTJlVH0sBcckUdJfEJhPmQUvBANQQyMNH3FcVKGTqhiCe2Wp6S066DPQO412UT9FaMTh8imbNCL
Jc2cdDmdYBZhDPbs5vZCR9BpyDpJNMkD4c+hh2B16F+WI/92kSpGRM+n8nSLG0mQGwzePhA7UGwW
XSthXLfcdYirVxsex2RfzqfCKeXfj/mcpMlt2kYO4AYAjWlWw81E9ReOQDCmE9PLZfS9SDoEstqp
u3HTg1SwBjvEXJEQ3lczDU7XDBHF9WvwtaAMZ3zQ0W0piZXh2gOrgYX1CAWvdcGPa6Kv14wqAxp/
gTEySQyBUmVXkdQS5tWQ418cZj681szQyhojcfaquOhUMVUYCvQbhTi0HPgaEGL7EQ+Ls1bAXZtr
wMS+USQRBImx/nWB0qydBCntw5QLVQOyqT+tJXmvdn9uwZEqnr8nB3FZYONXJzvClPJpAGunjLm5
7MzdGeyt5F1j0Wa3fljGfqwR1t24oZjNOP5Z7V/w0dUnwo9aNdDXfDqj1MsikKccFXhXv66jWTIg
xT0Y+GJkUOIF5jNzD0zFHDn8bLZpHrCAi512IJ/ld1VChSlF7yWHIF+EivS0fdA4doRh8wmHS6yH
QyreoknI5iCsJ4a//PY4Nd4pu5nUhIts/pdAPfz/gFqv+j9WLH09ToOmvabLbpuUkBGyHx5imAdP
qpccwsG5nnJEIb+15FdInNo8PQJm0qHS2k+Ks385hhhHJXTU1of28a5eDTDE32sGkR5PffvxTIFn
SZ/Sc8AcsKlgsJ+W7AfQooiGofK1tAzxFiY/YqNHUqcXY73XTajKIKavUI45g2KqqgX5xRH8+9FC
A+U6IAWdeYTpml8o6ZNTTW5AqEuMik/YmaUMTHr0MykpHCHEmkSNKw980KTJ+ZUQssjx+vxj9l4Q
zkGtaT3eGyMM6V8jnu+ZnQVFx64amYCOroOvgGZXn7gpuJhsOZMCNucUXvCxL46k+PqiM8PHr7zR
Ic63Mow+CshXP2sOhI3QaF7sOIArwcx3QfnCP6mZ6bmZG7dCDe4LUIXPgIvmvU6nQeeUdTAtwOfz
Q3wpjp0exAOvDLNJp7HVG7tO/+1Y9d2xTIdmOU9QiZXKMHiC5uvzcsdsIscBMSyPcvPNRCfqQkfv
n3L0KLb17+N51VrFFiXGRMaQKwtwUlYyfPmUA0sLTESHhu4F9yLEa4naIwRgc9ey1noEMg7i48nD
ythRjVUqxJMfq7HbXi82eGOuPb6UFzOeVAH/GWvq2X/JJyikhLuu1f2EwNZG9iKJaph7uyLrC6LC
3UROo0GYU8b7JmdJvJBXYlih7y5XY12DPt1LoGUWwVMiEg024w83UuKkDiY/7pDZJiJLIp+lomXg
uH7efCdqAKsr8RRcV+i6lyAvSC9c6eTOxtajQ8NavtnTj0sWXnrx/2s/RvCMlZMm1y/IYabsFBL7
iOCXT4gdb3IAxT0eFGarhgY/NvtmL6pUAiqGqFU5JQlT4MKku1ipaYfUVXBsLNiWORhUifjjbFA/
tPWp4sBQxdVMwIBPwOEQIquSwKFHUW1k2UKErjQVTPq8GO/zCbeC3eIpFmzYatKl+XMU71cwgI8r
db3Fvk+oovI6iVu2cCF8T8q4Oj0Ro0JjJxRNecL52z9CSi6LUsSedmTAHKNgNhqsf8KSufBqKg0a
uDSD3HlCT/r7hFkofv6sL1gDqrY+bFk4sR0CwnMEUxJZizX83xKWJjFZIb5LGKlmhhehltL5NYNd
NST5QkQraKu7404RVaTrUwQEmFsPXis2WRqniUUbyXRGcXs05Rlx/V2iPSzMs8rf8rSVEiDto2DI
vbDF/14G50S3YfEV9U99ZJR4RIgHKtwhVUSsU9JqSID3eTZ35wHb4ChUneOWBhF3dXlCEYTz6cHU
eA9hetGgmhnOjuzcfYcnL5viJ+Zzv4Ip1KmdQ8epQ/r+Euu+9uVELN6cI0mCR0iFJfHxah0eUHW3
thYFTIFHdSaHVEjdcT2H+oKzDIHXK1ZY/xT0B8VGMwjgt8sjiiXJMxbjlitfvLIsFm4uBcXJ5kLO
fz9P7RZo0S5GT6I7ORpV95ZNin0QkDYWrtu5gnSpdnj9qQz9fOFM35HFIBP6iWRT/C7WcJbT1Wtd
QTydBuveSw29OYag2ik2ACA4MZMzAKgC8vljrEkzhBFrcMfMukMGPbfDbo3LDeT8/Rr9Pqh1JFGW
nTP74AJ9qhBOJGEONb7WTASCvsIW+B3b8VBFo+yuUwTa681m790y4r+oDoLIlbas8W04T+Uy8S2Y
0Hsqb6F3r1hYue74++SZK4czW+NTMJpE0U15vtM501Tsv/+eNebhtI53+iS0PX68XznTDpTLXxir
H2gJeBfZ0ox5tTpYdj80od2ojCPx1YxQeCBWu0IzcbyPwp+4P+OcQuRNf9iMgmJK4aplwIrGIbMp
wpjnkfbRv6BcYrZFM3yUbKkc1O8n3JdMIM9jIMtEtS2zuF7mpXDQL8b022fN/0ZS5MJ4vAH8IPe7
1GJ567UWMwixZo/gkvhIWgpavDT8YsbkLs07PcEMbMrzamtYQO8V/oIwNXch0EXYXSLixIxPqXLa
DAhxNBXfZUjJPfQpYCeG1/5F07gbztm7OcpUoYpE/8Mcu0mhbCQsiHLx2RAVYGcCXHOZwKfI/t/t
QZJAqrLIVcIYpKQ9RfbCNC1m02WnwD5Ya4cLz9iN3+GQvq5dkKyobPSyWENMrp6WiUlaepYuUaCo
vXZ9F+S7xehez/atO2cwTt6XeufgcGDIEjTjnKQOrPFYeTgGy8IdbosJtgjfA88oW/3wXWEFuHnf
5klHKrPDiAP5pCAdxlIvMHZ2oRWqLeV10jlvdmWqt2tZON1CV5VmT4sdKVF6ymr8EY1fdCR0kku8
4zygdW7jmeMQAQvtc9moNMlV9CwN/hY8zOehIgUuOvrm2ZS+M86hvovBriNhga+/nqXVg5jGwHr4
vDcBpZgI423invGEZGSBLo4kS6sqPIiKLr3nMziZZONWfi9Ijmr6POIq1acImD7OAMhkKnMUcdQV
ffl3jUyYJVK0SpIeJaw7l5TInbHRHN44Uq/F4UoBTJ13+R9q//84E/rIYoR+sDbybwHoFzb4TOC/
9SOu8JyO4cEZ0MtleOEc7t5tjepDN5jJtSgRizsdTSvJdLbGcazzKTEh4WoRhcmRwnygUe2ymbwB
iZ55s9niwJ4bjgLZEue0QxV1AK0YJeqmW8wg3ems6YAA1+hR6EDNd0Pb12jj9M8uWGsaioTSWk0Y
VEEeDvXx2In7JLR0A8nTxY/3BeGhSVVua9Wz5SCQ7wxb1jZeXl8z4wrkD2eN5N9223DDg4PxxHE6
KiXG6c19MoZVQc+t7Mk1lDJGjsv+49nDdGQVY6TE+pc9+sdgGY5HSyiJ9Gkv2ObD6mlHeb2XmFH/
2ywRhYWoovxRNXKgf4dpC5EDWkmTa56cBMFVtv9Xe4ZnW9oh8a4WN5jXFXAcwrRlCZ/n/aoNvHIk
HYoAeM54/LIe/SynyYl0ZQLONwK9nWokmaXKJfvCTOogRVzzzjp/Aqc/2qhxVHFcDHNPXAunpZ4M
20CWpB04lBRnJ2uJ5pSLEAPyybM/9hFZDLQPmATIRFIgDXOTqG0GrNF+QUNhpqLBoE7vtcI25+Cr
HGXYlVPg9GOdzTX5zjPBF05MbhqOaxyYh8i2phkzBSjbItNLDQeDyvT7lejiotC87icYKnzpZMFO
MaefaR3kOVMHy9glnV8rIrX+9vUqNQnf1Ifh+1oNcmouY8Ylrfau1UuaDhTjfQ+AbNFzoFYFSBKr
dJatwDz7eCpBxfCeSlV4dwpWnikLKi7oC05GM0r7MR01lTA0et9ImAkhcnoyCjsRIxNMQXamCXhN
YkkrZchm/yBwiITkTf09r8G62pWhkI3mSHG69M+nOYqYfYMkj2ovSWF3tv53loilUQD9juGrpcH+
wtz1UEvALY26cA1AaCQfcFKeH7bGQ+a0GexmWuHGaZAMA1nHNMbuLnFDu4u3I+M6ngnkZNdBr/9g
WX95ugAbBpJcrd5cT3vz+6mozMbzNHAg687IOJbNqYoNjtMUrUnRJPGvUJMyEPHCLXw4FbHkOxOL
OoBTqYafh7PA8Syx/dFBmnLr+kFwhB/JbGJtVYqDLXxpSOthI9QLw1qhbt+PL6lT3YzD0XTqwwWB
C1anC4+KlcZI+VPS6tsAIvJgjNe7sKpTXxp40h3CGsZPW+lqxZ3XEvqFKST58ievx/KT+fnzcLdw
0QSyWdL/AqpuMSjdgj4U8Uwtw/KAbT9J8ImuxmVjTwYx587GDY/RwWTLIKXk0gUXhhMMNSe3OZIX
W2VrrqtTam8uAAwVuHJY4RzJbmqwRM0qm/ueehQ/rNZ3F6XV0d9MrYajs+rEXASWIRSDkootOg25
Ut1i59dp/n+PAQEkrAxZxNvxkQf3O+BVcZp+TNd/JmZVF7GDbKWmIUAh5qAtp4vzrD02X0/IRS4v
r7Us/8CFzy3LwaXrdXOLBmjS2IRQ+kkWeV9Z94yDBnbWY3k6eHgPp0bCFtPZA0wO++LFCuaSKb6U
hI9DNtOije69giMSsI6hufI109C2pi536eeBt6eCWa264Z1hXeENN51wVGoI6OizH2NPOhDKV49k
6B8NVOwPQHP5fcE74M5BMK1q4GsYyoPS0lgOnkkQtPrLuR1Qe+oy3Im9I84ORxvHtBkKGjKN7p+h
KVsS0V6/pl/mLhMOY0IpYIiXAObSxqF8VzQkux7+OD1mHua/NB40BQ8GPkgWFM0zDXb3piGSQY6+
31ap8PkUUHBdYjdRnOdSVw3dnaNwOzPk4Jze2U9ERKgURYqdX9arBT4mFuTs/6jpBZIhmXZ70C3H
NFpV6a3OE9x155X6qndyrhxX26XuZWw/XOZxBdRdVEavmLSYqpT+jmR/QrJ+UyjWqZMTXbQIv5QA
DwDW/JkCI1ZDaGQreYJB1pUKjrezIsVjR9KEIlKCHOj/q3r8jyUmwC4AGs6XgVNK8jrsxelIuTwI
LJ4N6RoZk6EOkqeovPGZNyzKdtaywAzkHgYAb3TRXbaBGu2BbxrAFJc7WO1I6UclzA6v1M9860D1
7BNLuthEMWcoRAI8jFawEOn8chP8t6NCeLksYllcWqdlwwZxhnZPndx4LiaaJoVT96N0++7CzVpY
NPayo/xZl/fcA0bSbOu3I+H2gOF9F2ADQP6l7x0Hi8pf3vyJVDNKn46oeoOPQdZNcmkLpPGrIWMx
CeE7FF0YECyD2MCNEIQ8/w8SAGKxFqndf3mxxfkjtaRRh9UouoQcaCiVW+vZrQ1/FQOJFO5ILmdw
5yQyoSywvqkiKKd/9bXBTeik3ZBZBgDGgYTMCt0LKVPvEmMW9ZWPhmirwVMk1HO9FvlUfpaZc2mD
XMs8J0rf9w9AI3Jjrnn5MxeGk9Mfs0QjNvSoIjmXcQqmA5tWqYLGUKOrJH9nVaz/CviQyfKjK9gU
2zhk5lcbKwM9g4FNkZmIjJ2v2TJq+05xEK7MXvPQ6lPCEne96524iRjcfg5JTTX5C/dwq52FUege
pQ1ZqjXvZrH9pJP6Tyoady1FzeRGt86wgCRcbJh2BS1lXkECqR15sJbOlN6KnhFFzqU0qjjvv5OL
H01SIh1T2wdfXncNCODVnp7TFTUJDDkMCerR68xYPMDPhvsXlvZMgxB7KZ1HlRc8Ky5iub/hSQzg
MwQGd7mHoCrv/WLkqq/cyQcfeaOtCRe3DEgzWJzO/L5Ff//DlrLeJE1X0WrcxCGoROI6FhVjhhLi
Ce+ZE5SXyGlRb8SDamA2XdiW/9lw0BnR65QtsqVp9BBjQA4YpplChKd7Ms1/9stijcuHK6oVVLA7
yXUUyucXV2yA+QoB6cS48lxG3fuMrdlif17Q1LbYXDCwF69F3adyxQezqo1Ykuf5tpvAVoB8TObm
NXaD7TsBHxzXTezZtEqrUmLi1Dv4LtzkRBcU+AnHaNZj76ktNKiFVeBrK5Rx0OTdnkNVH1VTurua
kxkqO9M7BHqH8LsXmNeMC1/+dnWlWoGHhYP2vUyciDLHYd0SxBDN0iIpjLMp8cppoVr1J/kj0EJ1
rcGPI5yF9kjqAl3Z3QfhM2bII5dilTzsJ2ATZAYd8iKf0M07DVN5yum5a3fi+QiXXOKO50/z5vbU
v4G1ATI3N1u0j0a3rZurpB5hg5w4FHCFtvBZxLpGFFyz6JGu86hYWSexIVbQqqXxknrgyp5ZPy68
10HljJIFG3nSc5sThNundz0PBedDHNIc1XFXw+1W1qEOOTYRvuat6x7oyoE7itiYOSM4vboGYd6R
eOP+Fq/kRL4Y47ovZB/UHx3lzsbPSD0S9DmVdEgdT15ozIk944Z5AXl5O+4VwXjPxlwipiO1B9Fg
y6AQzhYkzc4JizrZgONL7GLd6o7OQF70JSx/KXAqu7QYgud1f565V9qvxc2hlEgAqseFSZkuo0PW
aHMzy5NU5PjZafm16OykSJaJPwlez1QfWEU21Am7pPdL65JZiPZlYNwC1G1lqi5Bwni/3FsJ8r8Z
C1HnVqM0b9nFEN79gGCnRAHg/vgRYNfTYKJWeCwNnGKvALYaiZYK7qWWzC0hImkoVGW91gvDFlCC
Qeqwl2pyNy2FZKURvwGuWUUbbrCEdNNjs4btVg9u5b5uuFwzRZCqyNOmyebmwq2psoqSPQGgroo7
xJPyrKGw7GXC3AhMCnjpoI/6xQ9dMWe9B0QbtJIVIf6bwpEelar3miWSop7tCelCJJBPhe4uLdyh
7o2QP7whi79GzZTKs//rNdnlaeOmINUEFffB3l0xtMWjRdyM5lOnwXIbQHuepJM683ivzmpbiVh9
+XZILY7B35k34NZCxKumomRlBV7pIjHcfm8IsY51IyoFFIEOslYwmYzrtuLMWW1Gzs3PxMI2OQKc
EPUAcIU6j3hZK/SqEzb01SYGqQQJhLoIiKNul/wXApvCJQlSDMeqoRtSEkHbKfmRSQBTWjE2m/nS
Sy3+uP/kgBM8hUl9EyoKhmtmMZoOdAfxKlL1NmOgz1TGKADuJyM6SINmA8boKe4XnBqaAqacqOdI
cMXqo8QtoP09YhOwUC3GDtqR8n3fqN0vsscj9ZFZQ1QjCaKUN5GY0oP2bElY76aCh0BDkMKMpH93
Xzclwq99GPJdrEDd4k+I0DU7F8+RVnHm0BnDk8OQXMzwu7KpiqV9x/aDcyAgZQIDEcpCSTFwiKo1
26L7gUw3MO1sT2P5ZwbqJbMletdHS2rTI0QjiEd4rz05Z6Jcov2bWrtot8MvkiN0Xd+KUloEEcjT
zkYL0ahL0jrJRdXtxebcFK7qB36FyEohR0TOY24ecHMUDe752J3sgPh8YcvTuAdcinBJRsb+i+C5
NuZx6DMbgjIJ784ZuoiMl9wftO61bVB8qGwL1I+yNPPfXEwIm02X0u004Wyz6zg9elYFeG4N6hsz
nyIDHY3xYtnpJuB8lQR5/roKpYgWF5rnEtsDVVIINh9w8pldrrIIL5CA7sV4YVVeQxSG5kvVef38
jwEqbfTPQWrm2yx3iCCaUQnV+2fY/oXppg8lfrtSuosUqF8rzFGWTYKIDdCm/2dM8WG+8Ud8Iwde
YebmZ/nV8Il4Cf/yBh9CF3/HbWJ8IHkUMI0p7dwm4QPT1KgQK+K2i2bEss3u1SuJjSqtufjC6M83
788Mb8hDd6KTJaxuh5Ydn63FVcvl7WUTlgOo8Zb0yRudYy3irIt27axbjY1Rrb1xilP/4sDUEDLI
N7rKPps3E7jLCLKNmPFqPknIA7ysdvswB2n+FjIANKi3RU65+swP3ukGCoqqrwK/kRwKWDNz9v6X
to/XLP83FORwOl9Pc1XDbgjgvXWOBdo54493VcESMCFV0kGVOF/B2y+Ht3I8wXgSVP5bOwuWKzjn
7K8g9wBlZ06fIR6d/NHLHtbXZtZc2a2y/3xK67y3Zi2Jd99geJLnvJHFIiY+xqI12LzwpGmYAtHm
lGPj7oSe7VMCRTXd6XqH0Oa8XI8hXrkMfOcCokpBaNah+JHhWqBUkZkDBDH5F9lCDmHfYntEZiC3
VZb00EOo7RJKKtBsFq7JgdUhi9ocsb33oKZAeZoX+VFSPF7lOi+bzXFuYuroMnapp+DVLaqbgXP5
1QRpN2h8hVhabsc+mYLfbVkIeBzzdESvtVMwJ1WPKLBImA8LnYuOl8aL42Wy3So3nwk4sGyX9oDa
U5+8reGs6x+CvB/X5uDhd1YDjG3LfT5yJKTG+/6GZybRzNFvfMZQohjxFvnmhbzKcZ7pjH9IjdB1
XrmHYNyOKS+Eb6g2I6wO2Nl/1JslbJ0bzJD7VsCLf2QrsDfH+lMR/R4HaLziNfji+xFmBwjsmTVZ
wBnE+C9tmq6iQ+a2jpVeScjX7eAkpzICk/1BAjxuJJeRau+2Ktg7LrzzT29IzgMcJ6K2hic6bzPA
rdFzebxKRTyQc5+e8qNOq0MZIoHCTSZ75chhMng8Ow5QVzhbwIAswkNlHoThTEnxsEMAq23T2iMT
+0VbUajlvmTIkhzmb1rgKniK9gINSA9uOZvMGIe3ur2FH51KvfAD39xiyzWN9ayw44k4N5kSaQV1
IVZUhqcn9z4x8I6uX4rVbw+DJ0Ft1OWH02hqGlfpzuiAFsm9qYM4g4QqzrFDMFaANFhZxE5Mteqs
hg4pj4DAF1hTza0aLt6LwCKTsnWHvhQ/rD8iaWgJTGGFJJ3LBBh9DgLjAkt6aLXtknRdTGIKvcCl
tqLgEzGemEcjxJL6qOjzbNTQgQmvZnYk7O6z6h/GdOvI7qobgbw9oiFp3Ecwupt+NbymmGs5Q4XG
5mQZxTk+xejM08M9BmDVX9ekEkOFQvx3PDm7ptaO8bqiPPPGKMRA0k4zaUR9uKfsHW6A/W5igx9g
YyiIn8o7/y6cc9HQIuacSYXrcpGd+M7dWGlNWjRROtd1nmoM0YGbuhbfBbOdfHJ1IJdL8Hbact3z
/ucHPfoXhRE3ITzMq7OgahyPvaL8x7tTCv4DGhYRXnVd5IwblUVFd8Vaxex6PRgrHYtfR34EShFm
2EZs8Si4PjHzkR5FWQtN40k61/it3Dyhink1Z+P4ykyg/tBysmJcyY8sXCMUamEa9W/ZSxil7CDY
WmTWDPJ6UHzovIt3gPyDomcJrIAQat17H3/60IoVmi3k9IIKfkop1J9ohPUyt7fOz9vsgnqOjKPF
RClGNLGhf4R669s0q5Q1FXqJMw7CLYuso7hIwFYd1zZjVPeyz31VJIeXCtof8u+slSTAZJBle2xf
UjtcF2TeEwBj8RUrKsxy++Uy4kzPd04mt6PK+OpHTAxPyvoGdG5NnzPmSv03TIy8uCY6TlhI13fX
D4y6ZPyr3LetCgU/ijeqzLSUXrqIdk2pYpW1eDPePTbmIJRSPUgqUSFMofdbkhDl9e/Af0BO/E4p
swIVrHII/Gb3WinMoXq+UY6kAIaB1kVSaz/6XYDjZl5kIrEcvlNc7+QLW4BeLWNyiGOAu0rLVZN/
uiC+xIRgHY7/8CnUcuNy1u6S2Yoe3wJD6xqIaksslSH4UNHWwoKQfEWRRpTrftA8byw1etzDrsLf
u5erCu9Xxz/I0ISNSDxsWxmRGGt7KAujXdXm9TfHl0y4v6ZGO8z6C3SXVTtmFFOtA3WUOt6HzPtV
05by6n/InktrGtRHmo8zdh+JHAOTrVN838c66z6k+rLapQAKeJfg+PM1XIHOvEzNSKlu/pkitXrv
zRlhO8KKL5HJAFdB5mH0kj1PJALJnDuPq0wOQ/KSSpRpOLO/IguQeDQBfptUik4ikZlm7AeHErhP
5YLujwJNCR/a9sRx/NoiH+gsTJdrxWdSYuLSDh4qH2tSwP5jlPp8fmHsI3kd/rjuw0I6TMm6esC0
lmrAYHyPpsm/xCZm409DrvaLKe1X5cr1w+V5lNBXhsArQWkheEQugfEvOjjBroVai6vmQVFQwix0
9Sa1cKbOMZX5o4ZWQgtdmPIbdvBHdpyZt6aMG8h7lAGorJCiz+NwCzvsEy7w6GUhppLwo/kMq63e
CM5RYFvhDRsC2/c+FwWYZlb73yiVqoNOkhGWOLTRc+BXcryIdqs3r5EZI4BU//AlQSFoK/ATEbuF
IJPlFUlO4RfsTLWyon8mVMbfe8POgseXqa/cVBT+AobUZYPqljHSKG28FmPqmZdIgY0CB6NYIKjf
IN1tcv/U8/UadwOnTPw1+bBewC1nSGWPYl/umzNBSIpJKqL56UlAr7dJrEdWv7niBWcbhgY6dMdl
aVqqAuh7vxl2pJE3xnfzOKgJBCJi3bb9iiidW7T/Equ+QngilOGSNdZRGyDvJMmCeWqw+BMdh1dM
v9LYprzhowA7vuZzGDNLJR/KYyzkrco0L2bJSpNjhud62qV4Dq7K9KFbFiXUBJKI8BEASOIUCgVo
H9YqEwLQlCEIwSRiqy6YF6cPXQpnYdsRFSpDt3iMgR0PtHv1AKim/JxcHLfHkRsaQiftw7WkfRWI
6che3rMGJ/CSInxYH7fGqLan+L4wLaVAB/uuZwPZDfM2F+CPv+NWY0DkqUc7wvOggX5wEBGTtMxX
IkSLS98wEpApe6Gsx4CFZmqbyQ0eXRyYMM1Nu1+PdAPzO2wwx3fcoBVqlzBMyEChWRl8wPUSQl/2
qXXadeKHU5xpG+KuLXCQSzqcnZHpj1Dv9106eewAsVRTuBEJcZS0W20MWfrQUabTmmfO33I/IKpH
buAE43G4UXMg9FNk6De80G3/CVk+SmHprCBi7sXvaSzseY73BwVOKRq2vXIAQpai/GIPMagiQ7gn
Q48xHlq/78roYxSSejw2EEtHN/ebAq4oxQWcL74ynMYfBLFrUrkhIsWx2XQuEAhydxfu9S4QZvlI
9iJvqsq5A358EnVuMGKn2lxAWFIAqtjaf2h6fBHbe0hK/BDfvxS+DdeuwPhBYEU1PB+g/7VnNZ4M
Mk0PcOI2o8W1RvOPIagFvReyvMfE8C8mSvFImsZBrKsfsZD6mcC2kh942BoH1Gzpl9fqoKuLSmfT
iPNE8sacrCZws7xDjp+usKnQD5vK6qtk4ncr6SWTuMPB0DJh7MYYaFihVTyd4y1PRzKj86+CKwLT
VGeLSI755rzUjuML308hp0ww9Io0uIAl0luMMN7toYlV3wM4H4V4e4DNpEi1/4Ux1qgbPdrN0NXT
uODaJ3UuDhFZ23/OG/9bbomTYfet4C3uhujMrvLOahp6qX1oGC4ujMJEEHf17x8hgc8g/9bp2d3x
RBn63t/U6X8qqnJHuyDcdX0y7pjrj4CpJk3AJRbU73RGjGE1kRsbpZ7UQaGZozNJZCcbFFNvBpHw
UKY5AY2L6LInCoIR84fHXOQrKphCMFfkP9lZJJn2OBr9a/c4Wz5QvfoOc6EJuloOPiDVwJQhYCQ4
/V66hfc5wnVuR3mCLq0PYH3P8CNJCZutQFL7hN1WM8fkjY7hVKipl7v5TG+qifZwKz706xZtj8Jt
EcElpzkD67gphK+qNizQN1/uDhIFrH7YVq2ciLCQU6OP+uTBP7VFzWTk0uum7ued2RvswSg5ygD1
D6URW1oNBk/AYWVSLowZR6yHTTrKkaq3zsvkL8paia2lUYOltMy5BB8cd6JGkd4btBCc/3vOi0BM
C8DglbOKRpbZwi2tGVfPs3SPjCC4u1+i+z/0/mlbM3gKT9DiQv+88ZugaooLfopMpLz5n0PeX7I8
qeSzNKnZ84Uabf139dRGAVmU5xqTSsPRFgOg0yj8qL3586UiEb6w6ls8Xf1VKfjAEOT1Rx9zjZuV
cE3iFkl542EZX4lOtKCd3mC+G8sJQEDQ3XFCv9eam0ptHjbXApnykxGPTmAbDwv9bL2wzRQ2kwF+
5CXaLT587HGb4dgn6DlzSyQ1fXOT+UXK8YxlprPEl8wXECuM51pote2einCpwUVHdHF9HKNeN0y0
imcQxT4AzUzeqPUjxCIBoq4u7T3uLjWjiEgXZHX9VhjV9Lc2r+roQqWKV2OBwq1pq/Gzvo2GlMf4
tiYAT6q8UYfUy+zNlB6Q0bNjUXmA7xSJJZCoyRR7BjMLedK/dPfMbPxsNFzFnMj7VkIZjW7RzQ0S
jLBXrU5l6bfo4NwgZlLSVaFf5p5dQ5Gnd12QWFufKDHezhfHJZxp8fpEoqfewhkxaNeRuHHV7jix
AzlgvrGQW0uRo76CC5Ka2x8vjn99RZau5lN964dRjBtuApy3VkhuNL023iPyNSsh3kb8wqqZCaOT
HyPFJ7FuRQE2z6r3aQKSp85mE+xcCxbCvV5q7XyVV+hhiub2snR9ozMwUIoo5FXOsBZ97O7acDGw
9beRNfbnR+LJBBQ6Je57vk10JfoVGs7hyOyiHb3tCBzir2DEtIwpV6U55MUiQK5DB7RSGdsMIFpL
UnfaCyE3+8Ic31FhuQajg1Dk9nKqE0GhTHeF5xC0s4iIxKAXOZHqUKTv0Mk7PyE1C9ayHeYWRZ+d
YOn/FMObxUmVfowyd3zdBM/sQb/M6lCUtobu8SQBmuaEGF/6/SMiZR65QZOV0446bnv+TwSrOb3d
s20+HuJd+So5mjMyv8HQw6W4715iLnNTe5azIyC9dqTjHpsr/qOu4OjTW7lyyu9ODgMPINSK0QZ9
gFGsGsB116RZPMbpRMi65uUh4htXsIfijYLc1M/ELbdKd4CldYQ/zkMk/rdUbecKABNgaZH8A/Qg
LnKpey7zjgVzO7O6gu1OuOkvQujwWW074iEFWbpTes9uFQG/bjrXVvOEtA0shrFgXBTHrxjzC+Hq
8O+/FZNbq6OmqkWxvcovnUfbtGHVn8GyQMsY2g6hOYo4TtNlbxfNumKu3CZAfjP17ENcD5oh+i3u
mSYbKubYKmBqlZqzv71L7NZCM8XfHefEHraJYdSXrBd1FbX4HcmU2duBe22hfNERfENBJhu1dyvZ
x4TA9Usat+w6g8Q2CyI9CPfX5n9l8HBH4HF9kJx6xUtMFrQOib6lHYXyU9Ixt2xdW3tm9aTpzqPf
buDWprkYbyuOL/eNplJc9kZMwvSBa3c0VWNsK1ABRdzoHGObU2fdXcA7qV4c1h90cBw+ixNyPxe3
LFtUCVbINBk2yHXw9+XCAD7Q1clY0M30ai076vqbp7DAlY3TOtTS9sTLWAbQCOsy1pgJoCcJ5jpo
FjdYRHyLz9YEQLHk67kIyVUVtfaItvpcn5DRwCC9mUhNb2ENKhYkavhPwSwyS2gRABZsktt7SF+S
p4v5XTC6TuTQc0CT9Al+SNbuI2+KjKJN3CraOe15hmLA/Kx3wIIH6m0TqWkbbdnoBXZpG+IqadPd
kuY3hUCVbjl2NjWU21ymUwpI/APu/IexZLREQZGxRt7GuizA+n2+BnGVoXS+sj7TJO6pbH0q9zA5
MaSz+QUW2Z/sf9trKF7nbed41I/GluP4DnmPYhmkYlyWSLIASzVR+t2h5UljAqKgX70hnKlLg7sb
QrIKBCGPC6yiEFA7M9WXPVJ98DhWYW5KjIx4nKeMHujhZD31Liomepl6lKeQNXgUmnl7qbYGkUmM
e6L/kIuP3hrYXj+npqipaJxk474ETTz8bB38c3Z+SS52A09wMLxTyXiUkj9Lm4dYBXl4eZIme2Wd
esWlYzACIiqkbMFnK2vda08o6LCeaRWqTkA6i0+XC/I3LCu9MV1T4kWwY43xkEvaOuDILQUtsfRG
ckZxf9c9yio4u+sLn/99GjDgtFwZOkuIhxPl47C1Mj8kBV0D9VOwVsJi/8YuwymxL8JbM7oeuWzH
XvXy4q+IVw3scn3tTxryIbHfvkHLsUsyllgJjZjqAfgdwSN4ZVa2LE5KdrwPQdhGUS0CPjeT+IPr
2lCNJzRmnDmKP4fri/cxvqR/+PYkjIyWaUd30cBjIuTywBW/uLEujTcTlo3J76rSlWy3ljH2a2xh
p4CG1avJVstvkp/Wvj5gKvUtaDKd4i18gEXh+4U/8pttWtat5e8ABs4uOtADIoCQvnPq+zO2DDBT
P0jdJRtx7HWeU57RyG6iQrfvagBZAFCr3go6dMxJFIPOIaBCaptJVa/+3v1rFlWgzx50ghd8ceiS
vSmEAn6klKf5QjLE5E5wknlsebjqNL0pFpbE4kezvG3uog7/soG9GDtBaVLU26R8kkWbeyeTbC66
CyTNOh9X2auIBRhrNUAdUZE/HoQhXJV0qngKp8ReTdekoqjulBW5SGof2w2OXRCjOKn0J3ZNx723
xWmBiJb3b/7yo8uhOxYB0hvHZ9jCTPDZsx+xpO3pqnLb944d4XpI9KYPiDlIuiEOnnEMjl1WLXoJ
l2J1UNU5FJ/uKD4BBG1USy1d2/6fRYZvAZhZB/tJstRXQ2X7Uac2M+Fj8n7Jn0fGc/U5nNzNQuho
aLTOAFd/J/K/gtv1WA2F+bCX3LYbphJDmgYiyudV82BlMFhbrMOqVtbpuguYUZYsTjXg8jvqLxL6
KIRdQM9pjMNbeQfuBh6xkpuVGdoTMaYQtI1vv7Yx9REbHoFD3i2ZAVgd2Pq+7A2DwUetjuSxeBFb
BhtZ69ELvnlHWWvakFCSLW5f5O0hmibEyp3O54gZnzQXjHX8RhDP8Hm9ViWK+vt0Io9y8Fahzhvt
T9BKdUhxTZZygl2eFagtDgTdPgSYPMIaTsI3sqteyFTCPM826UgBn7boJ2FUtdidiVCq2h7f2xUV
hm71CJKnQkDQPjXPNrFavgkOmBKeny/0nmZFtiwb46pQFz8lqgPFdp/w/0nDU9bJzKj0FlAQx5aU
poQj45HwCUJbysKEaBtUkoPoo/01yodZ+kh71Jfw2j9ubT+YKVXxTTz5PUd6hVWRNifh66f7Kfc4
7yi/kdKKFf+rCq0wNFU4G99vbBZpTYuN3zXn9/hOoxGMozSEYGNnPISF01/Zi8GzWhoum7xCcnXK
W5MtRA+jacrkAPGSjgIaWL0iUsxyRiM41Fh7jIZd9E+L7ak1PpmzSRakzzcMz7ailuPYstNGiILy
BsOYO3SBpAeOZ+I/z9w9pLvWW2RJuVWVpC3HDplfNWyehdyAH3E9KabUaMu7/u/5K8c8fajFZyfC
IaZkh5igH3ZD9qC7lZRCwH1EXYQBEKw4ib9NYske6frAaKsbNSz5rNI/jEAnymw1NX/hOk0fRvCc
1UvzQewMRP0i3qgVGRxtuj/HlMzHzL0kFkGaW8Fs0YuLUD/li9qkW2PQH7X2uTprbcgBkt/jJjrG
jfaPgq52HUsz8zYtBwpBosjBa4eSrpsKORhzBWJ5ybbWEjFh7wrKkfquW76tUhDDuwzNdyvK9oXO
lKgnrBWsSS7EAgGh2IUS99+nEOIdDV3GBUy2SuY3LHgE/0QKyCxP2yfHNLioiA6SVV8WhS+539rV
zj4RldTf2eH1CCy+LuTAhQ4Ncu7bEW8ELq9BAQQdCHbOv5lLfQg/D/N5OW0rJoqCkp5++xIr+HJu
p5Z8KJh9NxMC+dylAmg5Bc6+nWtKs3DIsyYnrwQb/LUoeD57l9pmTwKPeH0woQEvs3OkgE/iwnNV
QTVjgYgbXtbNq+ylM5md0yMjl5Jx15pQ+orrAF0mytZV2WBU/q3wBRj2oWSJEDVLNRmk33Bl/jrC
9Y51yrSW6SMf7VHIsWV+m2u2MR6sq2C99IMCJwCnEIWT2hPdltbkzE0EbioLGfLiAXI+32MRwGf2
bGL2Qq0idgT/lqGATbzObl814nqi8pqb/LQQyqVUBFXezwavhW9B0i4yIPaQ1KJRSgRngFJ2Anom
li3zFTayjMO/Q2HEdM2xtwzfVRxXgwY9flQV4iEIuz9g4v2fJS2SMEJdEYUrBiXQyiQlmNzSEMrn
716lMxXpFnvQmKSYY70JKbAUjF7JuBSRWtvIVAr1YR1zyJKIngMRoYJ1U5UzaWjpN+ZZogQt6FUd
xw/OU1mc3ch90X0qIvB4xKKP9LTe88x/EwbZDFYphhP/Qzft4IEtr8o/qjjS5hEX8ktnDGVNykW+
c+fn3AW6p7BVM9uDgi9iJNfkN64I35BZIFRL5QhprfAPJ6rlthKRgmyv8xNySC9+6DDBXVIjG9wM
APgNGAqOys6wn1IwXrdXNPM8t98QQv+45Zku8J5J1D3YFKAgl5NPg5WibSKnDACq5gSkIMTGebEs
U9XXszMw/LB+DVNuqSDDE+7jtMJiJFOiHCVHYvAgdJn5J3LUnOQmtnJMgeY3QHNmwGDzmlvojLvb
BEr0v3MmnMR2GqMpapF2pXkS3ggqpGPzwnFVcsNdwKmlpi+1DyUb8tEIljnxOtaPOIjnpD3t44F1
9LCeyhIFpnI6wRTGod5cG955Hnx1a3KUxd1gZC3ZY5YdRQxvXwInc2ZRpsV1O53ycwWWLRjrq4Uu
95aKWZUGH8NdF26eQ+uSWiLN4GVG41Rk17PVsWblP7Y8OMmKTYSew2mJxzvHKOKIh3QoOvaB7T/K
/AsohcoivpHmO+cvCNrqDvbQyqNaq58RxxqGrSYsHCKCv1FAUWeqMW0zFzNuON5De++RzVh2YsGv
nH3FuamcGWcPxhwXbj9plRe8gNTRDEHyZypa9+qSR2hBK2Gs0ITfkbLwRNX6oRNfEQj9sCQ0Szv3
vMXRQbkpyNZwyCx+laAgtBhRUyll6O4KN7/yEk1f3oakoMwxqvj7p7f6SA5bB6UdyRqpOmeuR7eG
66pWdfoEcvmBiSM3PxlEwZFtQaWEERS0AwwiFaA9lNRpxIMulwjLxk1TmNKaQmLTS3GiLaZj/bPD
FBDaDQkVyemwwW2QTE+P1ztGHWHsgjj85w2evqlFQSk6ocSpUS85/AHlt4S21AgOh2XEIHfyN+tx
qP1yqnfz/pZGp9XKQLzoBguY4Qt200Ja04BKMqZrV5k8lvGhBunpK0u7nx2MNgbhOgwuS2avsOTD
gNhfjx3RDzvP/ePuR99BzIYn2hr1B4AeRsImZZAOdSIRiT9aL6jwniE86LvTAbyeI60GNe8YgM+6
TJ8NLql0o3cHOHIvpUTuBoeC0WayZIoGzJdOuw8j+jPj9WCL0t2/sdcTYQBaHR+JC9yH0nGy7cR7
JgRB9HKxjO6ry9yb+MwD4gAdJeJu1ICfCreiMqaXWoDFkRVvgf9/v7e2yfJdhw25EMpXQR75eQCO
pzRSt2D46gPuIeCRBbOLmvX5TlzwLffJOjAeF3IDRxGHTPEVHIRw1swIc7n6WD33+Lf50/N4mAjf
06bR712wWvKdslq2rK7XxyMsvNs/2oQbDF2Sq82IqVvHxX7kvWnRtih52njRtM7cBtdpZYCuMOXL
0RxsfgdZTaIKdTqSrRtuA+mQQIM336X1ug35uUsO1btzJW6bXOU+l6nfok79NRc8gj+dAMEDQIX8
BhW7egXcJeetjAEFPDHbXIsCm7pCXdlAIfTKzTm9kgeB5eCXtswAd4B1dO1qI+/jshpgP94tsjPB
TS2WRpeQwKpI+zvPw4KJShdOpdxTEFp8RRtRXNAsCXz9kGJqUkHOc6Rb2p+GZQtUd0o3QFuZE0gh
BTV+mQLJAO7IVQscTkOCOK0vL3Z+0ExJNIAyJ714wosKPZVE1BF5w11w6uZeL/V+Bh/NUFRa6TBe
df42E28/KelwZSawryROp7DNMUdZ7R+uFJXVI6lN2kNeZ7NFXTvAv955dfViWwYEwKpFITKhu5Y2
7GMcpb3O+jdurFTKxPWQ5YJMcsj6xltko3+Xr8Gh1x0JUFvq/iaR29erCslMj5nkc3mBIbBiSI5w
dNGZee/bwJzxSY3gQNbXR29s3j55Xh/CklkHDLetFO1IFTc/6wf6gofDNh4VAWHAnhrMRmbb2IWQ
ntSuun8ibO5T4FFlkhvEluaWPhZHXaadfNzKGxoHcEN6Ol9IkbRVa5yxPS9I3Ejv0paEJJ8iLUlg
ryTiqgyEOq7O3QKEm3DbGgsCTJGCru50xYw0DcGm2Sfsd6yg2RAMxMc4465KfzxUCMVB60YrobaS
D9706UUjVOu6ZMiGrXxIWUEB2dufhhbmQ7/VcVLrFyvuR8+PV+F9AWJCmGZs8TypaGKHpYuhzoqJ
b0iul9LP/gIrEtc9SbQHxlD7E02uAMY0hSthWT6nhWLRzYvK6j8e4HfkmRu7p+OFbfRbJDTKq59B
eB6AqxWsLLR+O3TkTkfWUa0Fpaxxw6BHsDgqRsiNv8DSHFP6qxF/P/bJN15SnLr8DySctJs/QLPI
pTAqrQTN3iPoHk0MdOllEvsGic5bRVp1llaekg0pJaCFWoLU8hhxF3qjd79+mPN/bpaZBjhdoDp8
syfaIvjUu558OxGNQ6kgZagHpO6TvxSvVFAJohxHjU+O9YVCwesa6vNj0sGfqHETYWeU3V/griAz
jHuQC6b6n0lMvI8P+b0Gooxu061+Zfsyx35B4wvZ8B58LbSLmMGDLUCOTCL5LziDo5BYhlx7kyG/
dZbOKYkWaGj8yRMULfowIWQBPGjjCHsRlkYdBS3egxKnOP/HOcAGw0T0fiJ6m6NSCtaHJRHkplW1
86SWVX/pHeqMnET5v6WXziFwSjbnq/dxOmte2NEMC0sFUjVF05cP6hh12AZkBjV3kXlgcOFL6wQa
oDLkme12wJ+wY43Gpmz26dw1c1TPlgEkVmCHyd8TVMdW1n9QO8XF+/bDHXEYrINPai6QszIUq+0+
sqEdIf3GwHBZj3L1bKe6sGTJe0mCxknSpqYteHVAFb2LoeJgILblxBzLjQSaWaU/ciNbQeabxtEB
w+qbSwCR7i0sF+sRw2RQ4i7Y7U/mpv6/xQ0PXSjigbxCVEUtJJUE3T+fivZEI8eMaJ845MmLg4Ey
Ygljuen0OaNbSHYe0Z9vcnLxTYKL0ywQYxb7rJeAehQwEbs+WlJu7alljGx6MUcg68zESjaR8eGR
jk7CgOR7lEPPv7PdFhFaYnkNjQgfG7Yl6UgRCIImg1m8wm28POeo4wi/OxRkJyDj3+fAEETs6dAi
zj+/JxvBUdrrkuQbItndN/PSOTtng4eD3ZJ1NFa2+nNfX4aoRDo0WPFPsn8oAJKCokPXDoT02Loq
G76qzixwTB0US6UswgksD6EIuHjnOIE4NAAysSKxLKB6BMxrcMPMdpw6xv7EOVPHDgf7iSboIMX/
zHwQgS2HJ0180qMN4EcjljFuX62oK4sCgKB4StOVY3x5Cpkd34muTnKc9xFQ+epxqMua9csNyVJC
e7lVMp8f63D2dUjrS/dTRFVCchVFjgEL8lulw82G74YHFSrrydzh5TD/zHU6u8zFB5F0F1u60VC9
gbRQTlYsz6wZS2zHp7rvNGWXdkITSzLG3jEyQ00c/76tGbe+ri2KOtcIy7NNWbCJiWiJdiJHIozc
6XgXln0EACnCLqjaTYHOTngqEvD0puU2Z/DyaNhgIMMWLbiwy92uPNescWy8pIoAz4y2sSqQGLUk
p6oh1r4eetI6eHTi/21TMKeqd64jZQ2nbUNARZZnBt82KAwwvsDRV3JdJYGkJb3JpIpL6t+/c7Fd
Mh7BLqd++6z/5jZdj3SSd9XH+cnfZBwpEwOiSQA4VDSfXmQlYsDPNNTTQvbtz3sH2G1S7NboCjGY
GnYi1bFS2LWv3lQ07fBQIiliFv5Vt85y35zd4Fvptr4lkeW3SFZKqGvkGGQAkTIefS1crXSbaoo/
NtiI4qrW1wxH/2CMHWeNBEYtGFuIAuIg/a25dk9hGcVHbaXfAFh0ISLpW/XBfp9lTBJoyD5tIH6c
2T0TvQo3uadakxeF/B+Dr7lJNEH/HbJGJNsqa4s8dAdfvatq8txbBZGGbPux1leUN5u7ZswxdDoq
tw5r0yxcFnlL1ggg2/ip2UhRxpUwJR55U7OWepji/HeHyJorQBUJnULW+WH74j3RTJIIgwVo9lNK
QqLtj3VdmQyImh+vtlSVc0JtgaRLaSpuCrLIhPb9uVbHTGzJxxekjOLr2clmARYH09r8FE6D+9CE
avw2LI/v0Ps6SNj/3t1q+yqxCpxI/72Sms39/M2VmA3qkiADTUvmRrTtYCcoUarWfWwzm9LYzC6i
qqSstjTYqHy/Guw2OJoHStD9bikjhJ9cnIt55D8CCuIbbUmT1Zf3AGuwWa9R4lLmOu8BmX9+H7Qi
OhE06ETdidfDYPMdjTD64kcWVGPglQcKPhAew4bClt5hY0r8qdt3PqQN/sdIlp+yzsZhd7gtOZOF
4jxiCQ/GrhI8iudYrD2yAEeIvdxeMi/xANChWDuN2Yn0jQMJjdLcC+tYOUnC2Vp43i5oBGdkZrvF
zrnLI5ANMgfEvc5AQji5JS0aESbyAkOPx5yDcFOb9H57HjQ6gGHi9tgh/s+1x+pRzRxvxUNVAeT4
GANmzC7buFNn3htcRw1SuyuUBQC9+1x3e1qlb1ftxaxEyRruHIgtK4Nn7DnARVJDoGleWWsbYZsn
AToTS2dPCAbSOxYRQcmLpwbJxwW4ppg6AMWNzumnDDn7KvbKPOVDvnzzO3y1wbqVRV+fowSG6qrs
K8Gk7iFzLD6RJZ3nZGLH1JgkJvZdcmYaDGOEynb7l0dkgTOSdPSnkt0FMtNUN5+2zp9SqWVK3zJn
BnDfyz+jqgXDFWY5Q73EdKifR1byppHewX51XVkax4YkHTTL/6lmS4buNLKGvDOGirgoq+K1WGnx
3aVvvpXm6ogRiWm9rfcMtr2S9nNE5yPlzG49V3pFDS/c1pesDs+Q6vdfNQbcLz/4/HMBTJC+jne9
fs7kvyJOzuc2nzvMHijKsyhQOEIuOFuY3csju1n9u8t6oVlPUvqTw6f7Jt+ofva+ABF+6LETqPBp
r/nW0fPHPnx7OPIdAtqwNWKgrFBCOlMQ3mxfe884Cqlaa8QU7Nu20r869HQET/xcmynd5yTCUh4q
zi/7gHFALOj471qXPtFLCsvvFWQv+IH2Z96rVcfHH2I82jQmgwmU4jzxTwNdUmkBqLrx/X3qVcs/
nAgrW38eISLKOeCA2Pz7U9NtpQCLcjBznnuX/KanvTRZzhEmfhf864XljFIIeWmaTT12STS1ov0m
92uDqsLqMpGcLyUHDYUXI/2+o0Bcc+yo8dzrirPzsCVYNSECYCWyP4MBJvPY16KDZwqINMfSKFbo
dTCS2rUw5S73MwqAQzhk7MJj6hmCaCx+l52VHiMC5ZfGuo/MkPW1YuWsImBFnoGJN452Pkxj1rTj
+L6tntUH6UhEWzhWSYbdhkbA0ExlxNJgrZ74A4V600LzuoEVnNdEBZf/8+/2xWO6uNDFW/ZN2KgR
D2lym1ZHtx1/pylRmR/3I0z4MI9R6l6o83Qcf+BMN4om4V5aHoU/X97N0myfKxm7cs0MQSRND3XA
ulyXQ78VdkT13a0bmA8aH0pP5I0ojqxHaX6GiFnTcAJKUyu2QgjVKUS6eVa2x37LN2iXTsFDHVFa
N5sX8ukHfKh5TXmEsR/4i9TrG/cJiL+bene2VW+wxdDqUukNSAd+6y9WG8hivVlSzSrYam0nRnk0
gRHszgTwyMnDsI771TLrzgsWEiegL0+DEZoOPem6O6vPsgx71E4ueXDCfgdkSsBREs1NgB4WjXml
jWX7AL8vIEPABqyd3h7Qi0aJxzer/Ii6V2HVlgKTyVjy8Pdur5JxzE4/OZHa8Mif+wz2E8KPCmVJ
ooWQmdcnDOlvJ+xLF/9lbXeqyfv21BpYpVL4Vv7tQTy4gXbNUk/a7x42nfvavWJAm/1vwuCA58H7
xi6w4Fyz/5d48DAk+1XvAR1bbSdt1Wiw/2YVUdlQZsTWvFkwULvzidTHOd1qyZpiP8CIbnSXjDfS
mAhaI8xXw/C6vKrknsh+NWTngpi91ygcqJyebRaIDPShMBV6EimCxeUzgvbHc75Ts0LRdjWGrIDr
snqdnmorVFyuli7mcKghbFW5+LQnLgU3eDRrl9eAjkutJTWlo7owdgX/ImB7SSME8xtLdHwuk2Wc
19x0gX85IC47i7gB7ZEmzN6VUirqwrHAPFLh1Sevou7l8EYL8OLEA4lL889mzCA2Sw9vuUt4TOlR
S1WbIo2uJGxi0e2x/nKJTew28cjXZ7wR4tTL2pvSDrTkf1gw3/R7UvjuGfzW4oQ7cqUYiHRtiWZU
ubNFgeA5lFVY/gP/GLmV01Pn9xJ2m2FsigigSemwXymw4VBQyCPBS8OCsDNkJapeESGKzmqgjg4x
8Ol7mE8OtEEY0hWZEnfp2jdOu34pGOLM8ehVCY0Uclx2C+TeY7jr6eddYbwF8DAZyrVH4HBI1RmZ
+EXUfusUtTF+EmzALbRs1gh8Vyl7EU1GZ/ygVQuNotEzCCc18ZmuRRnktVyESm/duy+GoPDSIs7O
c2FD8B5UGAVHyll1pGDKH5rN31YuIOTWlbk95VPp92DDDz+gjMt4qbAlJ7HaiAPNkL4sKHb28edV
5THy5KnrpXVV6MR5TiVpgKN8k6U0NUX6p/7kV6GdnFDj6JDLFcR020QlyVj/PhkPQ+EX9c1mgi5K
XEKzcn0HUMFci3jMg2wlb9escKZMFUvpquMdyk9usaq3YhCmvLS6TOkmGazf8VyLBdHlpPCKclSc
W59f3q++SyGgOOM4O3lzvPktse9vWQfR8hmhVv2ZgNcukC2kFCa4PdZ89HIUMcWKWFY6k8C8Wbcj
zKM6kcixMAxlt+511jLLuWQ5rgjx0h7T8VcfPn7xJuHrvWk1191fYa0Go+YwshuGbB7vKbD98p+k
5dLODXGBqs+Jbuog/B2pM/Mfgeo74hZYHS1YGh4WvabEa0ogec0luPreS4lVtj6qGkGTrePmk9zN
vSRYvxD4NzkHaCzOXYRCOLkYlBVQ9QRDzWQISjtDfsrbGGUkrJdHwNCphcgyYOX3G/iJfIhj6Aep
KIXYfZUwyIInKSH2t+N+/ljmjPHgBcQk3ZVfzriybM7Z8O62hsQmG/CRGekImCF5bBTm2SDgnZUN
8WKmna0YUGR4F/IDcWy2SIHPEmpo25r2soaN39efB8qY648FpWl8T3Njo3DxXqnjE5Gr4hNe8QKJ
yqbMa4EwNMHDW7MyYsmyfF6rp9DNwVT/xUaE7VIZtTNo3Aic7ixeIWN1TBYf8Xtp8UyfLhjqNSQ8
3SUGuy8f350cqWv5xUPgsdVgvQBt27v2W5yiRXz+D8QBtkg75P+D6l0e134gCo6c5mhLYxBkThrG
sBxYwL3/E1a82vkfN9sa5Q8yrAmXtr5sJXV4z1Nt5n4wltQV/5AUVmPwoRB5WW1KH5TvV4x+zVfM
OtETjiJthansr0VTZM6sYNg3I8SpdqugujBgpyZqRGeNM81YBnEKeb+Dh27ZSWItMo8ehLXgfJc2
dn9gmaou3Vmor81UzEhySihKqi4WsZi9nOivl7lxRtTujChSnGU9GiFd3oZ/Nj9AEc2EQPT/VE0q
G2ZHc+zpmZ+pc9FGzWLsCFFDleZ8taoNSVNy/BY/ZgQUEIwDI1xyWUFH8wZRoLdeQcbA6kqtm2DG
MA/B8oXpQs3y/deUvHKOkxeCCxgpOVI97NPOywTjDBDRPe0b47+KXPt2Ls9++QX6XSeYOMPMLrPD
NAnIc4nj+ls1neMmeinUr6X9eFqQSY9HNZct5/lmFnMdXm7gblP7CitqDjpW288wjdxZj9e8L1Yq
pyZGvP1nuzsuXssrmcqU1XgXaxdM21sl+n/YcuJRgKAETfzGcIJtJTbME4lRCEEBXfJ1yJEWPRl6
C5CwBbGccv7A9i7P7Lt/nGvGzsZV/z2fAtC5M/BmZGgRVqOMPkdRLDemcrZIIJRhvrlGu3dHsQVt
wNOPgNIyoXp40YUonFR3dRLXMEX12iUwDzNF3PsQ/D03EhnUP39e3QPRFLzRRUqmQqdkzp40braV
72Mpal01A/itLPRdcFpNkscyVhb9Bf5UDWJ+4zNOounQeKUS1LmuJMcDF3Lt74bMK9V0Y289a1zj
CQug9Bcm4xNn5fuzQ8kIwUpEJnbIau6VAwsc8iDvj8t1l58rNMjx7NkitgZnNI4WD8UO9N+w6PVV
3x6rvzzGgJl+a7T3votBBgwJ7t3R+ynP2mVzWfkQB0DuHPb4PbHmjdFhIZC1SV73xSMTVgyRQzJk
Y+/qFoE844oPHXA3A+uX3EW0o03J6H4osQ1mBKKBgIMlAxcsDUcd0AomjyGmmnRcTiCyQHtjITDn
MbjbPO3XAwPAbmzKQQbqECAEXjYCTqvr8hRrZLjY8fIvqb6JNA8o5igR+cpzLklYHvpMKZP3yNMK
j+HIR4OtJWKpDtlt/IPS8Ka1qvdDM5qC+kUw7SlDF0DsVQFlxyJSPqVg4/73XojtN82ixP0K4ox/
u+2fZL5QjxeuFmfQ3XTRoNUkafgUonccElYiSSAN7zK//1xHiBaV/c7K70PQM9o2bilIsl7EVv7W
yiWQAVFJt5Ie9Gjyz0wODDo8mYEmFUCoX8h80JrtahKZxPxwfaqMnoAD9ddUrjGkitx9W9VlUmWY
NyR2P82HXbzIrfQ41pnHw9GZiTSzYuuu8Nruodqu87aiaUaGxi+skr/q6VMrXzicWCIJjsx4H0wU
pKFUisxbvNSytRwGYAonNhBitCRDGHnHUycGztz5HaXP1I6xRRdTaBF5kJY3jLy+aHR24DLzUs6g
C4ManyyyxszmBZUazDfBGBQGDfBcIf+S6ASvMaJC4Kz7ozVguLVFe5afH8x1NGjDHLW5J5PLKyPJ
aOE3OwEXhDfTVL2i+Em55+TE6HZiUjJAxeUOH66QVymGmVvxhKvnYfVl4PRjmL+jOn/6VWqcoZni
crDkeuV+AT3FAQp1MxFBU58W6X0Lzu8wqhpJZOixckimBErUpD0aAL1+XVAinXHqGOSTfsfL0C7+
W8/F42J2Oc2/6FX7HwHxKjdcbbHpuB6261Cp2xfHUFFuIqfIPlgxKkAQRK0MXPwdqV0ImT/JLqOe
0+3vx33H8lMs2nwyn4BxK7mMvyxxUj9bSBluePu/w8pwTCWmnb1lhc6UjwpP2spbT7CjCno3Cq42
Ns+owg9Z9xSvrZXVHh53b5RWdCW3shL1Jy5zlB/sjiObO07L0MuqPoTpEne2bhaZUVPEX+PvhtZs
SNke/QsCKsAj7/4hOxPnETPj3LLZrRcC5XbRT1HPD5AbNvjEsptVCjsepyn6fsu1EMlzpDTJaA43
NPpG479Ag0WpxNwqmqYMX/ESXQXYyqE0Nn6Ov9YS5NgJTbNx44KoCLW6PMPc3SlypNkQi8tL5u+K
T0bprrHbOOy+HosAbjz8QH6VoHJJvxpQ552dUSCtDM34OC0cum5AgSFIzURbNwbRM32dVEKp9tbs
GhkbkMnPpSWl2uAGkAqaHQQB9YN4Ve/F3k7hdK+FthbonIrFGenL50+BUk7qaybCdnkRNzr2Wzqr
LhRJ55UVUp/JUGfOP9AnkbuBGMFZq1iGTLn/HsbUEhaVNW2lG7mIJDMrGBEJUVBtyrXgjyGvAVlh
iUnQJQo+GOPLsdVanzJ+xSMLgc2yJ+a20lDuycVZb2el5wWX0i7ckGCiN5tB0qwjGeeiA6Lv9tII
kNXTKiuSm0T40AHkgsgCQbGFq46r79B/fidt2QZgGdee2pSlTDoPziIVn8AjpNGxmouL7xE4fyP8
HiRHkmkViHW1nUHuZ40OLWS8SyEy18NKCRTuYSIB8kKKFzBMu2nEIcoRq+xMmsCa4O9J+yXu1H4C
SkiXMLBve03LkYq1Kl0KN3WVa0gsiTSUqYmcAJUOOY5oBDfNtdst/dWGtxZyqKHDfOXb1AZ/VDuh
jmuRdiPL+FsXa5w24J+Ckj9W6P+RruGv4KiR1i3+fNjO8MSDXVliIO18UJl8Jyv0OP5gDXZeSXWl
AFN6x2Vv1Q/r0Khmht3A4R3xtIZEUNRieRntcYlAUVhhmfCxVts0zxSpIwsk3QSPdmSM29pLsa7Z
sC4r8Om7GPEkOICROg0xWFskGhGBtCfQ7fY6JsJ+tM5VhYtQjeHztSEdWWB3vEvaou/ELYjuFN7r
reyJHCso2jvVbtkr/KIc1I2iwDgFh4QsMTfk193/qMHF/eIZ96UDfVOQmSAewiFE6yj+eNCPKnDK
CmHQKn8IXjaElcDXVlFAOTMmMU4KwxqEy7VMv+3HJKy2PYwC2i26IS4IQDUMYmyGwIY1x/e9ZCRQ
yuFMJJ6bD8V0zgckUI85vZ5h8yUq25GeMWF33OebDu/By1Lib/+KuEQq7JSBp8o2Jr36MLNoYfK1
Fq8koD7ffwaN13r1d7zDx8vH3LOz/U4+tr1aXp/e/iX8MqGEXR2c4nC5VLa2SDsV0/UquRcqlu/B
QnJE9XCA1xd2eSCmelQHZIME5nSJgYdEY9tvdJvVmK6MlPmUvnpYxo6NpCoaLNtMsaa7XZ0TpJI4
0ZrnOS+pV++/kYz72kZDiQbDGJmt3WNFka1fIOBpDXjRToLQCtpatV9bAAX3ZhXxIA5vBQVf0aMx
dZKzXPDQzE3S25Y3VajD60MG71s1fU8H25bQ3x0v5vFUoym4ahfoxD+Ydl0AqdO9A4t2IUSQQc+P
2DMy+19glZuui9CO6a1S+6FRSjdfp7LQEZCpup09DvUAYHNzpiy10MPMIFN8A2G7K+wgN8BhKm0+
I5D//JjVdQbePdwgKIMNtocjXFTAGInUIS3epSZwV23G9BIdBg9sWuMPy23qM1e0DfCtY0nkP6A5
lnZ/pYOBSY1hr0JG1xsrF+2kaic27tlXqK1RY2FsaDGVUsHUQvpkVIafVmPaSIU8JLdm+ET5XTMB
evDa+Gtp3t30cdGYYo92VTQ9DqPRTBOX8oc2J5i9xEn5pxRcFJgCQm5R6E7Vu/aTUVGM1Y535595
1iHn06KMVudIYEgZsz2MSR/Bx3wghGoFncCbUrrZl+iZaAlJXUUAcN0lAQLI1syfJa3NQ3eyxnpt
cVGbg7JuaUNB8ul1l+Z1DnAJMQW0sfgmpcaatFfUuS79sTOxxo1Qay43ovadj+5RQv3NmIu/GJUI
giMG/3pOfT8wKdlod0sRUbWr0PcueH8LSUBYdZiTr++NvYciPdY7VoyJbdIaKBo4uVCJXQuELcvh
ifvz4O6HIxYNfzjTLFlsdi8Isc1ok+Nps8xtN/blSd1zcXCdnQmt+XDR/a317cDezgtgd7ZT2bK/
IqrhVOTT1aBTcG7vbGzRDdiXbsdgI2SwN5TdDH8Pzf5nvWxiULtjQXUtG80oaW2UwKDnCTXWthwt
49s84ON0A+esVhcjR68saFkU67LonUjVK9iODv5pWKRLh4A49bKs3yS2rO7lKWaTgolY+Mbsp5ZA
r3ax+4abKikyqvJxl/9iVL0Orvqp03W8kfd8jkQK/ZNKhR5Qz1PLQ2FPcSIayGo+Xa46mAcWZwQg
7qWrVsMp0jq/OUoBhk9dL84Bw7TN/XAFoVkBkaitiJNMvTEVrCZ4VJoEOwpW49DucO+9yXnbzcSl
k8mwdLZWl3RJc4Nr/jtS7xCZ2sC3sRSt4So1nUhKnOLv9jjtJ8jdxXrrFTrFA2ybltHKcMdCFv8/
2CeYk3mvEWEKTUXBNkEtB/aWfNFCziXHcYnCP9yMQLAm2mD0U0Ngv+qgIJVMMj3Ykosi8LOhIiRb
zQzhuwtcrBOTBDXFWqlPNPCvtQZz4YsvsIVa8lYScSwv0NL9qNqhDBkNeiXy6cFIf43AN6OGSN38
7+vh2CEgdotbSV8FMC9kuNRjn/4Ye0rfYXuBrNsT2GAh7bnu2XTHR3AUND5BRc328slp5XT4Zbnt
T99ZTzUcXwB4M6EbAj3Xj8672DWbJl+kZ5B2ih4GDcDrLX08NN2y4GLtDDtWKo6gpHxbg0aT6XPT
xNm1a9zHOrcMb5xkvPQvCb2olyNh4qnE7umq6msyLjFGjbpakwyWg3sa52Kv5GKtHbAoEEO23TsL
oo25cRAkQIV7KtsXviZByQgL7Gg99VzlQ4gGFanQSlba+6orbxRmDI6nvRXa0uSIB1fDFLuTXWi4
sRYCT5kfKZLjxP2Z46bNrsEgxZxdz7MyvPwjlQ4Pg+c0biatw2W2ZyUCvpuUCzRUqao2C03YZMpt
OndgzbzTPX638Bctk81+dChmGIqqrsqWyw0QmIFwFSJiIGcn/RgV1f/vYLSKTJ3S2khXhfX7MdGq
ryKUtpQBEoJK5ch7EV5buZs8azVCFmJQHGyNgOpVPcCWdtV1bmtQWlawnYIwxhmjXv/Oim8cU8c2
zNqFhQUIG8kjd9IlVsyPBpyEP8Rgf2w8+8+Tg9bwW22neRECrRomarGwc+npL2/QIkUZiZnXaim2
DBHBLOlrhR+c2ZIq+MF43nwwBITEY4wWEDC9lFh7po+afUwcHSEe5NFPb5cvvNjUMIoFlN9OE3Tg
urr16ocmXgMycE7+nQYBLrizOcqcPYjszKAEWT+cve7T4mmap8l0kJxVMLUI3bZp433zhPELH8jX
NFT+rNJeEgQWmkJnoEYLmO02VI88Y1yP2P16Fhdi4Ev2uRpGUhzWIUTEtL/y6n7wHSJnFUtnIkzx
U9HQDa5dUyTdlhKNQAxgGsj6+KKdHk9JTgVM2vxEuH3gASKOwEWaPAM9EBA1hVF4QDnN1aLEBWYX
ZaCUHS06lYi9B71ZzZibr19X8FxCvNf3//ZISo9Jj5lM4FH9JWxM32A/p3IJDWLpCOTFU/W7n1hq
i96wT4gNtMZJHcDKF/ofipNM39gjKMVmlmZcrZ+b0tG+Tjm4yvz0D4BZHTxvxOh7Zhk/HrIRVV+2
lbJalqCjna0hXIUWb+agBQcKNdkw09HV3RzTc53AFNbau+nWad81Xjj50dpARyN8nY+o/eN7Eijp
P1yokciPM9NGaKghc4VOOaJ3lvj/nix7HLYitTbh9y4rFdwO8mQKASelmXxFEdyTXA/YhGsXLDdm
iiYrfysAXNqU3/5JdycPih90H8Lil/6usM95eZb+OURdY5KM5ka9h1DyyRp2aZrQatnGDCaXRn9R
AXlM1QxTkYjzv4vb0vOK072WL1fogACahw2miQ06OsNDosCRj/9ioEFELcZEM10lDkvvCD/6iL60
3/6Ku4tG97PtXs4wHdw/m3Q+hIkhUWXW6QTl1v49SBcWRlF+U7SZmMaDQBsTyrsCQLeEUJQrLra+
Cn4xQVZiAgAbFNDC84HAP3qlgkgiycARcIhDs7WCYpB7CvLliW3Jk7ihhlOzfzy2gAeOek+CQOPV
d7Ql2XcSMOLl/eBe6P1We/kfjMG6gQjcG6wTG/nB7X4abwd571gbIe00C9jq4jVnWvlpcPEDHaB2
ihkjrpoSMkbznw2jSzi1x9ibvaGpUvqWoCaRye74tQYKYYazrHBERN2KRq92jteLwuLCud/qZ3BF
5ksfEEr4sslpzuVj7uP1me0adIWFHAGyXgKVWD5+X/WqcEKTDd5Tx746069egvR2ZaqK14h/mcli
xdy5N4EX8CwpfxXagxWbtZimX3T4GxyGgv9CEzcqbZGr/+1lKDyniS79rYJ7daEDmzfG7EhkKP8/
uFYjJ7VtnMplkqsG/Mb1x7dBcEgLzwu6h3JNDCTt0FfB8PWhJy/R0/7tlSVhgBKbBDfhnhiO200H
Yh8GmEWHDnTIP94FvcJKYmKXkyUV0EPwKZ2NNd8/HpS+01PmZv9wHMMrIFl4lDnaRhedyW2YboE5
OJOe+D6Dtmy+VzKSwn5vExfadmF4SxyrCpbLSlE3HCq43/fDi4dCYaZ5qGi2bp4bPyFwWKySzRlE
6pb+1Zm2xqkjPOcX/9mKLU83FfieXQOwKccN8uPX3ipxCEjte9ZUt211fPdNAKwhBvrpwtKUBCzx
HAaXmX53/szXTE7AIbWSL4KdAIzhjmMwyuPqz1tbR9/iUtf3an87oDfKH9FYayZ7VlWbw4xk9u5l
iir2FRwXJkFQuSZN08EeGLwCWbLQPrJN71OkYgzrfo0yH6K40fiLRGc73xOjqd20rds62UTkWg/6
QEvTdQLaJL6ua6yuJ9umlWteiV2Eg31T8nj5Qm0eIseHxqx6dnGp+bWqAXSd50WEYMVK4EEIejH0
iYh3unhmPJ1Q0aIoZhgQVeEZ92fuoSj6Bh1punb/07vDa3NbW13sjtk3yWft7zCqYNKSNAYLng67
3xHFpLAVBiu+ZyBKrvNRnMa63MMLk55XRl5jKHvfijZBGqVMGsCdiIhiotAXHaVAfEJmTmp5rTpe
rKhMPNGMft3BzePym7it2ueul5S9slVuH2VF8IspqaTQL7htwDPe2YyTN4lPcx67363M980XC5KM
sYW2wkk35X9AbjVok69bvwG0Q9PA+JQmT6Yy+W4qMtZlbtxkDK0TWM4hgsorBUBVnvjPG48xxhAh
rfaBgne8yTE/Z+NcWYv1X8aa5Rs+W0UlnnYAFp8M2YMeAS8ZYbOWqKG41eLI7Rk52W7jowjpwRWY
hCXJXJi/J4asQ55XXxWfzTHFMlv3Z2C5V6uRpNak2D3dT8gl6GQpIuQ088veU1s7/nmplqSUDN9w
29VWV9L30S80viBnmuK3tm/diCaXMuTAAodDPju7RnQlHaZwp4atxyQUt/esDNwBUnq1nu1U0kXB
3EC9UMnlX/FP2C0Az31VFCR2yYsZdLFVF8NzX3bIWL1hbNEbADX2PczS1u/n5+JdSLQJcC7fWoVj
x0MsE1NLz511/oiHGg+QxAJ5DXawe5Zzh8Hjjo8fWlReO6OU4cZcNzxTghvJGPP1tOa1K9Nfynt9
+UgFKvBGc9kIEH7c8HKlesqzSEc5arEseH7ymQsnzriBVQXcUMxJf7bqMmZZB0tddFIyjfW+hb07
RfqXDA8MgmhuNRyxq7cTC9ghBaUAcJLeapMKPqjPYrX92+tU1PyHDcvQ3YVQUYSDQ1BvToulw4+g
KQcc6NPf14+mMewJ4ZRKt3YTbkLCpBJ+OVTJBX6xtTx1WnWmKmTHTqMBD7qunuQ0S+cQOVrMD/E5
g6+8/IVVdTpZOUkHWc6bEL2o48R3e6DWt+jwJZ1WWHcRQZ/OTQ9uISGT9v9eptESLhqvWGZHbzXJ
COyh2iqThXsQwtTnjCTsiXbCbuNz+ksSz9FaPqDku71rAa2MZIArm0yTJoqsQsA/O4D7y0u8eILO
fDsa8zrWBbIhSddouxrMQ1QAcz95CVwS6w0Tufr1of3lhqFZfMgvMTKHhP8Df0ah5vLoUG7RZk4s
Qli5+UjyhXLwc2a3mVULCbk5Mxq/z/zcnTiy9y67XPR3DaUVQuqiuWKlrIZ9oUulS0yVus12ZMq+
iyeDiR0sUccy0ysnk3U6Uasxe/DrcUDqgSqVKu1ftVkTdpmI7NntT/lT/jFNOdeNcmPxH7/gPmOA
x8ckXX3RTqXy07CB7spb6VtMLmQP0naLuDWPULggiSZ/k8DBAIAnDrjx0R72N0YTRLvfHHxreZAs
twxUkawIbaXHkAtKfvqUoNn1IuTwlneB1B8xrE+QsJykK/AGnBa70GmxVUxJl7TyyFnbkdRMEG4P
eyh91LzNvUCkCMZv0i4Xos5+YIM8ckNPD3eDB215XXX7NGJwQXvAwZWpGdwnf+gnHSB2P3l5ObME
Q/FYqPLfeVZs6mIQRkZ/dEiLUUyofOM8l/Qt67rNh3K6IuCYlp7GaJGotE3mRE3OdcTOCGJO4fHn
G/kn2AiqHivrWcf0aUTTewqyavD+8za3eKQWCuIr5upZDiDfpv2DlTr6q7rnsY0yzRcWszB+MDhS
Ub+HTfeTOtaqI4ujJXHU49A1DCFoxR8zzAsY4bpHvzmYstltLM/79hw5c1uSNY+nLv/VZO+ESbhC
EGm6dHrKXEuUuskx1Jdi1DKHJjAJrneQTThnCn+aL2nzXd30dF3efKjUh+UbZ3gfNGb5Bp/XXfPJ
pf3HMBTvVs1HNnLzsZbTxWnuoF1nr8MQo/AP10Of0Re2R5MnvL3mPIQosx3cJMCzC3wovJPn4zC4
B9EKSR9jYM8dZ6KZ2RetzrMbF5rQVsHhZmJgBMswcH5IXXw8DnAfymSdUOZeLKXdE3YmZNt8WaBN
yVJwt9tKycfi60WIqDSY5vv46nRVpNqmxUX8Ov2KYn+U1jXeCmjRDL4s49N1v4lDOhOTM/k9b8OY
z1o487Zqb32Q8HTlHRD8Ng4YYaLOvQyWFNq3/rvqvgJSlWSBFie3m5OyvbLf9RNy/R4H1JCCwVEX
Wb3E/+WYA8vbpUx/46MOTqfjGXJ78b2P4/zJnLo6KCny1EVRwEbr/8pEjGKL8IGRUnYEZgLYRege
27bhMY+M5QFxO/y72hG9zhfpGdI7x8Dl8RNINMauhC+uEO3d+hIItD5+nfJ1LiRkMcmOyNQB3G39
n9RE1hA4WPyProP0Ydv4XLRAN5RXFaNli7nlwPe0ngs83UyJZWEvQW6QmFyibKymAVMq0Pk6E8oF
zOoN0wko6OxokDhg2nydfreHOe1PA+CoaD8PkXyp4XQOgc6sLLU9BGxsWHf90g9d2hE09jwvjlLH
pXLSlsESX7StvX+Lno3ZoAneoNY+ke96GvR1CigkADTGu+2Wtd+QJaYudw3d0IQHk+j1iBz5T9st
O+Wdxz3CWaMtoezjjjsly465DFfWTIl2UuntSAOLtHM/bf54R7A8ygwe6K3Ecx/eitmyoCWaAWmQ
+ZOJE8kO/gR34tWZDbSxEzrhIRunfW9BMr5LqDtq6HKr1Rj8w/YUxRsHAhdjI6zvfj4ijvebKuEL
2Y8GKHHTNi33eqzjmPXmjufxYXmD194LeRBg0aMejrtEftxZB2PuLxH/DgHXRwKBuUqTEoWUyV/j
X473jF0OhnvnBDIcFtPe9mQrQhsYcM1b6gm3vbHMw6CdML12+lS4o43GRljTBuj4fWkDAywfPkY8
V4YPTmoqwvSapt574vylPe30S+IwYXquhpeRFrZAK2Hgx+MT3+luFz6YNmCeC9NZgtjuKovQvCuN
4L9FrkJJwNbyeH9D6uvyUz2asqQzAsBMZenhET0pmLGls6hRluBH7ryC0e47XZJ0h+1pJg1DqLMy
VO3oCS3H1SZRT6XI5Ugur/9ghw1pzsUYaWJFg2UZtqyHThMu2BjxdpQLicJzizFo+12Fpykc9a3F
YDGs4PnU8vlLi4yff3l6dK+mHmXdPsTeK6A+LBVPIEHJJshURfzi1idn8Cc37TnIKG8OpJ431P3v
QCLMgJvIvF8DgSuNgnUi21LFEmKxk9RAx/jJw2Xub1xqRIh7nF2NAFlTNS7nBYDYyC4YnF825ZQj
1P1EHofxDLY4YZTAQ7q4zaIf9htKO1PhRhorU8otXaQlqJzTzaDmMh0xM5/AP9xZllORZkJKyLyD
IszM0CHhntIzZ3U0C8jDkqDAyAtQ4DbmxROZNsayULqJS1NsJaRBn1JleW3O387BwpR+tg7T6ni6
slgS8ysVeZZdXX8tIa2ZFvf63sRuQnd9z9aQeODDqObVU1wo3gvJoYYVWmGpCkzXIVUCFLqSe46t
dOC77YuIVBcjQ7697GtgGDcwqeq2pDcZtCpdpLI9t7D98BHgNwN91M5VxDKF+QrXHq13b7xl1Xfe
Zt+8HXjNUdmY7mvvzThjvO5zAC3L871HFQgs6CBY97jpAFtTfFknzmSxNcPhGFqXzVzarw7YsoQw
vA0tPGnHdYiFfkZPJU2PQdHXk10Fk9hUD3ifyJhjJ/XYLVW+KEj5lzLD3WqBSn2KcuFqDVA336/B
7NxqTr5yOsMizkMyDRTy6DRBCCS9d15I+Mv0LeRMkwWNvrRtu6p7Jub7Qr2x+cuTtKivxyF+I4AT
7qJfl+XznlDkUzXXWlP/WwLwkU6VkihrkjkghX5ywynw7NMm/ohZ56gn4ZnfW7Q4Fz4djV//Kad0
5dKgzRWbO6O4hA4KMNzqMQKfNaK10XEfujCq5RbeC0qy1a4aMM1Z49HGGbi3z9VLepeEDavC3QL2
g1X5ZkOzFG+iE40HzZYCCIw4lbul8ciH8Icidr1T8+oFJRBPGrYIW8YwRtVfE9Ph3bAIzH9Am98b
NQoeHGLysHRgQLX6x1XuuNshC1gkFG3XU/XeWzxRgKfn28TiNygoh7j3GHauJaBmpgSUmvGjZ2Dp
3gIJhiah/0AP99JzjUQr6IePna+GjVzvqdloUdhnTkCiZne1E6Dmglx8JcI+gQcAJErVkbEOKO1a
s0uzkg1+284btc0nLIaqABPEh1IMC0NtDeBVBUtK4n7eoh2aW5xd+D9WAoFAKIv54MqjBNGs4Djk
EU1e0Ue/twYucg40cc++n2Fsyh5qd3YNRU4x3wNwYlzc5mTOvvAt9aB+sgK9XBxMP5vkbMHFHgUn
u7ZmUZu/ObXvsuZR/7umAHVaNl63g2alOChy3kqyeJoJrjIkTxlgcgmA93DsI9zH3JFc60M7hYYp
cmMOB59oLgSMKKPQNog+SCZHSj4/HD/Qoa37SWdDfBdHB9wcnxBLoIlrooIUvkbZKj4/9LLccwZa
MRn0PVm1F3hnpAhIhsOEujt1Hm8yTtlc2R0u7Irj1gWWmba8TJOV+07OlFfz06JqzLoLR09NeNK8
21mABLgNUVH225Gxa5Pfcaeq5nGCMKJFZxQhGQpmvXTEUn26MOMBSqdIsfWjt2PZXbiPGSmN7AoL
rr1pPo1S7f0Ej6oyMJ1HlZ2JzXd2pNQSPe5d7Oa7BrPybuLVNII1O6I1vWTDBwnLiPtcspooicuh
VYTwZpUzcMAmEzRKNY1N/3ttnjPONoye/DrvvaxrlVsrZeIRVc6NCK3YksH+bVDZxm1ubDhxN9rL
OVvyFceQ4cdHblxu4CMzWuor8KBrTaTXilaj0byb8Z4zVzR/JAy+hJnJfoJHmlHdEaRmBQzIJIVP
2Y8IT2R2MNMoN6iVgXgWRnJ6F9IDCwJdzeAwCBiA1m2uWjZB9FRk2X8scqh8Ob6E/VHKecj96l/z
rFxzXD5rFvSCQh7KR3Jrg9gxN7FI7yTblHGZz+Sb/LVrosciQyGmgzfoOF3UqJ1ugp4/r6FGRKKP
y1lbIhyQjbckuGi9s1VsqD4Ei8aHsRT5EMJhpttiWELwy5DJa8zb85MSnsjQjQ/fZSnltcnYByvA
+bp79s/xWSe3bG/VYnreNozw0laLJDZdw/Iqf8CO3U0Hx8e9FNoe2PizEe0E4Uavs5/oXV/p81h7
vIfSqu0NcRw5B+imilHN4qJFpF/wfjkDvr/1gw5HrNMu9PD7Z6UhXbVNCVKwnf60CoT0SG9+Ffq1
9l+cZjLU3MJMQpElH4hVu921yOfjB45bX1syI/uMtHb8f/X3cygfQdYns7clfFxNfD0wVdIsBASa
HUlMCbQAKI1qwGgEsGk0Bh2TW547cK8DrhBK1FjGZ0Vzk2ZrGXTvA6gSFCfUhajw38YF4eFovE0D
Q9vbfU9nhOeibxsFBxmRpFcbipquJIkIYbaG1GBl7DxkuU7cvaeidLasM4sX1js2gWof448UC6NA
0rBGjYBSZ++Hz8PIIUjSfJ21hwZqrsgM8eUDotyMveqxHwmazVCHT+xDy79fcGFdA5mfdQR4bHNO
2xzDB7TkdQFiv+05Oz+SJhHA/l6JYU62IeqnmCe5iRahjoMIXFiRZLxKsqRSsZHwkM3fNJ6QrHlq
1tolCO3HU5RW69rWLVffA9qqe41+3sHaUowznhYVhvuEM3+yZWnQA4Adt1s8/VQv22QcL9oopB0w
k++nAdKRoH8L6+RJ08PiZIv3Bg9AroocGvMhfnNrHGI3ickSRcxKyChQxGS5oI7Y9cV3XaTUwfzJ
eis5VaY1VmPtJGavjqLPWZgrsg5l10p51WaIsvXqQACJe5DoCAwOYYT77e2Iny1e4wnIwcyWy5M1
q3njJ4yxdwKdQusnd70+pgfBBJmARnOXOd2/al/TzNw7txwgtRr+lBx+8dvu9QhsYXFrHaGViFyd
dCxYUVCJw7fqIHOCPpn4CUVdEfM7EDCAmiy5soCkynJgD6GtLwjW7eiZsI/gdNZkMF/XuWlOv4JA
BN+WIxyj2yarb5LFe3EmrWCySedAQlFwfiSa1m0fFYlHsPtekHN/7cYX/Zcd3Wt1q1Mgjn6k1PCY
gOi7VzVWEMWssMrz3EXwhS6Knb/SV/Z6F7Ut97yw76H7M1CitpCBA7KOVX4h8fN6bBoh5eVW3qSM
dt9HHm6w9K10+lQCRDAQL68n5SrPZ1jgWXtIIuCHPlGWvypksCDF9VNzMbYP+WzF0N3UCKgBKpJc
Zt0Brx3AchaprQ17lwVbUcpHVpZNBw8gM6g/RH8K4x62VmlR3PslUmdLoF4y9GvhAo/JCKhYJo1f
Jj9VWu56Gf7IdhEXqI78gp0yizKYt78ugQtMDXFcgY6UPin/Ye6n+CIIAL6yDRYcMbBAz3Jopusq
/zk+lxpR9ybXaQ2grL667iDMy670Z2q8T8XBGJYeA+BIAmySH5DSkPV9bTv4Ijdb/YCh2RkqwqUQ
vjQ3t9hITF2ho5xjLxEnavMEjGXMeLxqd2td7CIf28CZ/zPdQ7AANqkjdNCKA3DMOWK6dJuLRVvS
dhEkJV6jy/luwf8dPtTcWsHqTkRUnAMEwMwVe6mlod5s6vE414UbEs3q2pwnndRqnjvRTKYFILu2
7s97YjI1aDwURzmgSKcHvMzYLNP+BzdGmX7GgmJqTTPpqbXdYr5fbkyei3hiW5cErZl59jsJ64Mf
34vb8K3X00BC815tqxt+BzimY8n1bT580GvU1UkqhjF8GHQVKOnVay2z1QbNGTLGSdO9sn5eUMBQ
nuprGxX+ewnfg8QDtr1OGqGReW1tlE0N2fS9z4g6SKQL19LK+2l4RjeJ7GpOk+UQuXHIfUIWIFhy
nOnQty0Gp8MVPwuBMJeY//GhkSvjZ8w+KmUpSYbd+avkfp3/1hh4xuLfg7q5DiKVoZ0V2hYgcH9E
f4ko559bKNRTrV99Z4dr86p1oGpeCh7ZdSgTJgN6B1ThCTSm19VsZDls9A63EFgA+RnqrleYVGLp
IArzv6AEV1LUZebDgsmxx7SOcTymeKRM8Ve1J8qgblPl5BqIDEzl4I8rCYt8zmphamW9CALdREtu
mbsojR51rhFLcFwyo9TJLcp/wQbwhz3iySbckE4t3eNX2S0Cf5L2tY9vAvaPGqz8kT/u+ArL6EWO
nYsQP1NaoJsFy2p5+buyiRAw1EgbqeLMqRsKlXNjVb/cWINvYtKhZBLtZjH0SMfCiyXGvJhtmdI4
6VP1HkS7s0gFxlgdcjdwLdY8+UMt0yPWKStCITQGqCmxieVszjbLSEvy+Is8JfTPFfF1L7bv2O96
mKuemdo/nBQ21QYD3NNEXceYYKHSTci7W6FK2kGeMhlfE6yMJji+U4sY8bSHBRQEHypQZLxZPl/O
I+5Uyctjum6VCMaBs8aYVpK+4/Tk1ChgxxY0Y/CZvxUspPewCYJrqGWNm5DCgTwqoBeKJ/tJOwGh
c1NIfdARs5bk6dStZ3H2MP/k5MIuEsPJfufQMUimCd16RZbLouG6SNm3opwi2ELDQbUaPoq4bfqG
yKZrMXKIMiQVJmOU1iGjkFk4oBkAxAB1lwA6GTg5+3Fh4ncLewpiXauoMlBZ7am5r2Coi1bdfwaQ
gjsQR5CVUBdHSCPLK3nA02FyWvxeB3Fu3HotkkIdPDs0X4TOg6ictHAYs2FIsz6WBjXZSLw7vCy5
+4hLDttAaBveG7DD9mOaCsdx6nTbUOvi1Nqk7NMAgsS9Okh33GdfSbSTCKF0llwjJ3Wl46tmh3J6
cUsTZD3xW1rL2afOBjqpLIXfbOfBXMU8UqgXbBBBpEo1x8XxM4isNXZzSC0oSDeOFaf71BonkyKB
C+syZSxIemIDUAazgQqt3djId8Yf8RAGwU55hRTseM2h6BOWp9nkXMA6cSu2FnGMli9aRtSNtl5I
lfm9Z8S9tmPO5t34hn3aKC0SimBOZX2AkOWKbvNlP6y3u61C/V2SKacTi8Qs8J/2Isf9AdZVHlbw
cqb0XbU9OpLNw4qX0+Tu6O/9MY3cxL/Gwx2JGcUslOfd4Yf/kSZzLYEeNHQ1XK+gWFYBqrlzL7im
qvFQKpg8l7wFdwstzkNnDB06u2mYi0At3e4XdjZ7ccwHbjgfQW+cA+gDEMLSPz/LErcAxgZxU3Er
3lbhptraBztTNhEt+82JUWp9Nt3qhtdqb6QzmRoSoOEPnfCK7rEEya6gJ4l65xuSIkH3yxbCQSAn
m7kOBSxrtDKPulT/c/2uNkSo9wPU4pzmrqqowfaZzkZmzibPzGJrxo41/9W4CYfKKH71nAPQ0xLs
fULz4RqsMQPeH/KNAltx4BM1GQj+m259pvyLkt7rn2Rjvt8tjOAkJgKTNtzaQdFDDd6X3YOxuYT5
PtbDtB2CuHMTpoVozrjIvmk/p5rtgITANUKlNscn44LPuColpmm8uyKnLl3u4cQpyVpexnAhDT53
LbHfM4bDg8ccJxa6+F9pYByC1Mha2Yzn2tO3t2Mu+qwgu+Gjjdde82Ub75q/IfrmhXCK1KlCj2X8
iXZ0zBq3ZQ8Qu9gf2ApxK6vDfVSkB92XCam7fKv5okr9W8VxSiYm+Dlmhti/tN3BMUpac+ibNJ8Z
9pbKtI3krixVgEsVUrTrcMczjWW/J/ntOcalbfoYIZkIwhDJmIlYSMkeW5oOfwBz/clmJebHBoR+
BdEdylQ+2J1HqMZyIA0ytKleBzGxO13MsR5ikEPC+jXY/L7OlMmoSPOzY2gdEKI3QChTb00QcoBY
0LqqMZtY/nWtkeiI0JJSRNaJvx8rVaRLuWDUScIGC3QYEdxfaeS+aDDRn3tguctvKJ0zy/hiYI2I
aaOI6WS2qDJBUO5dunJc2kMZ6914vMO95K4l1/4f2lQxN0xPewFnDqWJ8IhGAfXHBqlBFU6VNjbm
7M/1bTQNF5tuk0AyBikGEYzu35uqbqBoeasD0daMu1cBCW8kHAPdjmuBDiHddpQs927L5g3QR9Zg
MDQFHKODo8hMIJNb66Mi4VYZ6sM91yRo2DDIImjKVgYRBD4L5FZAWwbHaFtpgZBgitqt5UiKpqqP
Y8+maveFBLcdOKs5WPfWpGIAjqo2WGG9b4AEN+1aE/EtU1bP+z4qZHQrjt2YTNVv/3B2G8BAdyuZ
2CYuKRKypy8SjpgK+B4H/w9hC8YQEjeMsG93lugGYnOQNrZLSYOsd2CW9okbc+CWTWZ0gWanHKFg
UQ1tZK0svFtULKQpTZJ+IfzohOvpKPoe5rauV+NujQVYM2xUP9yU+mfbBfG+61Eb9h998ehGpaH1
0nz0Y2q6Z6AlGXKbc21iQuLBUuYQ3rQ9jJM5OeDNn176f7OvDeD0EW+Utd3j2NPtG9nJ+CwA+jtl
RVJRKpKDeWxp9R+3OPbk5oL6wGretKIaITcFClcdDWo0qdajN2fiYHd8/cCNoVTprnT0q6FI/XWZ
PBaY0HVf2ZUjUNUHfweF3bCNkWoQ7r5HaTPckJEOjEkSWpJu8qkA3ZeIMaCuMbdkkcfk7d+Ehl+5
gGXfb7ceU3ngxVjQmZmL6zGNIUxszeiwVYfQf2IzcdQ7rl1q5JEeIx7LXcZmYTtduGK5RzXl8rcn
WjsPNBcHl8mhrF59SIaRBuzLD4eEKxBN9maWvqwlfGLZbEQUl352mEzslXHBjb4EG3UqpMwIwnNC
o1c5gaZohPqCqRciCLT1/fZXJ4LKmXwMTCaE20jrlz0/24ifeIlWBbKsFKY9wNoW4rlcstCsygCM
3PAUWwp/byYJWJ4g1/uzE01uN2HgE1xgUs/QZhgIInESNZk+zpz2GkTD2nhUtTAZco/rQrJZgHIm
5UEE23EPOushUgx3csdA1+1nx76ksZGH1BPommsmNKyZIDqswQPqS9f+sB3z21ylWck579Huu4C4
LEzk3skLyzdo2T5dVff/vmOW7CUlPLmudcF49GYa3v52jIrUbS24xWQndMqCxTv8yxa8iPdXmEWI
rdmXT399rLpDY/1l2FgKmrSywAHTYTeJtlVON/9dfGAJ3/lChN37q0Vl5E/qHzq+wpfLkfIjrXcn
Bk20sZv6rDinD22BeaQ9cB2XhJrgiu2n74bN0EBJ1xu7MxbTSZrRH99hJRRkl/TwfNcSZyqrdVet
1xa0+VZrbORArejIrQUcyxj3LgSLWt38KA0rgZdJudLONflhd68CgaczOx84qfGn0m++NIg+sjvC
6BxJdLjI7IBHRx3f1sibN4nBFHeFfVCUidEXv8d6tS0zbdFs53IkOUYCLwcrHeWa3ebyU2k+mQDQ
3Kg2V5BLNgCi/2/uKJJ+v6SOmUm7OEF7JsU3qowLEFEYBJwmrxTluEJXLpaLc9H/nGq/pQwuX4jB
6z0KZyjtA5j38dJ8mdMNcOu8UY06zOYMbWRWUsA1dT5dSiva6i/girYcFPY4UukDGFiXHVVJS6fs
um39ep0P/2s4nNKoonutMl+47EKOmCMCdRVj3Qo/RcF8ViAMq2Lw8zJw+OYepH64cShJBTE/GI+T
9+O0Qs0x9Qd+HHYxe/4ZhSjxMN7hUhAMSej2m86HA+CFtLVT/4SwHb8C2HwkppVfmIgtYKjd5jK6
uSaeDPTKJJPx4XCxn44ihLBdrW/5UfncLmMmaFZVFYJDvoADgWVy9CDXp+Bj3MgNNxRMl/FFSrDh
LBEZaakbDHbDLeRff5ju34acncRx6XvX5kJRUULS2dZDSjf6a2tWoDhDtfiR8Y19pt8zcn0fOisi
RsKRunp/49yEpZQerrsBkodCTCyHV2M7bw9ucqC2/mnmLo7OrZ1JFYi3rUevPmCm3qmr+dySbXmX
uEGehDIUveSFi8CtAgJAuW9bYaw8Cp64ky1uPbY2UI/3hW22+/nFadv0uE5nRfJ5RPw1otFm2u0W
joNxdlkBrdevQaP1k9zg1RMN5wOH5n9XQy9/UuP0ZP6b+BVeJa43PQAl7uW64SqVXWhU6ErdmHnT
pEIzqfsFbqpi86ZGwbX06+o9OuMxvHYGMUP6JYFXgAxpLe04bFQdF2i7kmBx7J0+O1n7R3ad3C/j
NPytexjqk4ymyCWU7JgeIo+kxU2/Speqqp1S79Jtk2hU67G12F2hp3yBVTa+VvnYKGHQJwZ9qZBa
TOPHuSahFXP+et+P6rNgEtUvbWo+y2DCAoLyxgvESqUSJsc/TpeZ0FGn5Lw1ttN2o3MVjc8VVoHf
Jrj+ucCl7NbeBr7Mn41GbdWub46fDvkFv5ci7CcqrgpicTws3YX4xI6lrX13VVrNdoMRN7U8PJNQ
PtElsrLV4WiEflGjboTuhAlVkFEvaTIGH5miwJtD158GKxQXmaLzBixbxH41A1p7oo9PkYHjAxj2
FqwC6Aw3I6x6oAt148t5Vd8suIGHbhE3ReiQs/zMnN8zKr6Uu7LGGm6flfkxFZXxhqe9k7Y985z/
DFD2d/rOdlPVf1QuZ40I/IdIxmqDc/vIWQY7Jw2cgyYSPDFPaxOhXS2NhqeUFyqzo7Gyn7HIEmCv
Ld0/OpaPkAiX4Uu1wgxw+izoKXaUfb+9xingLUGbo4YQXEmS3wpDNRGmH4aCcSt7fyHS7gzlybqq
YVlfZInb84L1QEQCCMizvqOatUlFa5WwLnNQclkU3xF5N7Ktd/NYT9/1Kla8bygqaIvMr1wyc8oD
FtEdrdeTODVV1ViOF76uAkceBhzubkAvYYa5P/zVg7n3Jhc4D+wMXGfwFwQxsCLEGK1DmoJZlAZP
1c6KByfZcPlGExfcrEatKKLXYHsMuS5IlmdL8n3GIqnGrFdccAv+Yew+KpGb/NNfGM/73NfR7YAi
Gb0j59nhKQm49BP48Ce1Nb2KJjzU2RfHDoiNpfA8bO3NtiiXJy79RNtqtDIESJZ6HbzsD/g+4FXK
ZMfmIrdS2YHYn0vFGH0vVwhqfuiAAiQtf59P+EM6DyWt9M8Sk24A5/2zIL/ZCYEQ6tuRlNL0hYi3
Rj/3Ad3ENI/kwFeQBvzE7GbOmftNP9u8uTl98h2DDFMxfFPDbbx4LoV+d6yE9YZ7iLTjMXjBCmMD
CZihwa+Ofsq4uWtnFC+4BG3Bi3Atx13y4q0ihCYcgUjZmNMGth/KWXw6+tlBI+s+SsjBsjs266te
2cB2dmPfCOihfvYcwWqJppdvwPe/GDy9gKd2TzZRYKiqVsrcnwHvWuMXQ6/zjX4eO/M/fxF6rRvn
Tm2yKJ7UvLekvvT86wh9Ajdw9UeQs1Hhw2WQJzH3iCShmwqL2FuyhPvCERVACfjSaRJR9EcwFICI
Xrb59BoG7A2WIiM5qgbhFkGOTAEd717KqIB7jzKmD5bIMUi/ekEVng4mojlglTgYWaGD2a2/rICt
x1K3cdI1xmM9HOqWoFww1j7ospcChBqGIYoLAEmINbeLphHV3EttxMgxE8LS6susI+XHZL/xaL4i
f9MhSxH+Qtcet8D7nPB2yJpZ28V86uCy9qjBQAcRyhU+uxMexgWqDXywr2d5qYusSht5CnU4qaz/
Pr9j2J7hi/W/7qszdj1Lbr9l6GYU0hbTbi1v0EufkWPQRox726sTyM4e81LovT8N0iFdD4xrNRsj
dsaPy8jFmAFHKL9pm8aO0NCSPEfa78rTw9MVO3GluFdyA7kK9F30fsR8loQTgGrt0CGjhuDiDyVm
LzZ9aN9CH8wE0f3Nq9tcN/qoJBIWjERlJj2R3hMMTHOHVjNq9WAEhKKSNxMK6Ol4ANrxZrz5bW+G
sMPduSvkdSfDrvLTvHO46scKn/gsF2aE6hxU8fL4lXQ2rUFFVkNeGXqwvMxV49pfLDRfgrFlfTKC
m5WsyzRTsAUR6lXWJUzFPfuhSIde9IC/tlqkIRGSnFNY2ZWScNdkOwXI50GBwJ3gAG/+k+Saebc+
l3Y+Ksj6JdQAouOpkxZcSlJpMyMaepiROHs8QaP6ciSVZtWerNwjykq9KZc00CQvz8IiyuzejnkX
Z+VYBRyXdFwBnyBFE2VXNmSc5BBlaT/BLjtHjhDaYu2fe2/ZYNEvpLzfvNatcaMvflRtebODuAxW
JqttP1uEsY3WMTudBaZxj7VRbYroiXM7pqnre5ckezR9pu2G1J1zj1aOzIbml4qO7x6kt9Cv99Yo
Vxlpnqtzlsb+xoi178wSdUQmPPXLagtd0WyxNah8zr32SYeOrIZKdnXbVh9/SPYpCHnPVv9GgTth
07wxNJAsJhqs/oNSN6eKL92ldJDajPialLckuS1cH9pdqsauptvWBQ8EssO3BYOMs+dbURoOymhK
K6c+BnSmLEzIB2Ol3FGrF1zBxN4ubzAeqvYFaaDc7C0EIRXjTrmr1rQMrmvgrBJ9ytZ2mL10AGys
84RFch+0I8koIpAPrILJ4VLYi/W635qDz8It8jzyyUPBp0wfaP7f+nK92r8C3N7Tqa3PcuRBUVdy
4Bc3ovZJjBuX5nSNfHiqr7EnVcJILNAgay5Gw0E7ezLfuM5XjHlBticBgtrmBwXQRtsZnnNhaZNG
8ShCfNKUQMvKoKTmVoGkFBK0I2jaMTZpR//g6ebJr128eZHzV+JC0njqxabXHdklYNUz63aeNaCZ
8voNeITphpbIL4hLv39LZboOZYWQQPUewUN28PNptOsf9vV+8vpQHCPEGMYEoEafOjY3vSOAgC6D
qXCfgWM7N1Cz/3/lN8mluErmx+ajg8cooeo3RFUPuaupOffcKxzfRV/yiziPSNlzqmYb0eajj5mL
avogX7iBl5eJUgM0QykmrJvtRBxXqj9II/8oGxHEv0thXFilL4d6eJKDbzeLXhUCPQEY6WGniJfF
ZEGU1BsVEnvJmaTLs8cUO6cMJSn/gM9+v+5G51iUBRpBPNItgxy2TD8Qr6SmqrYblsANIOPwQM0d
tEQkv/ktHEvxmtnWn9wEwOjiOXDTW+pg8QNMN13oxcLQSvOgz7zIAPvWkFK5ZPaiC1VL0QlWCEhf
ELxw7Mo6Vy5w7auydZG4trpZHHtEJFgNlcZDAXdxII1fnzn5RI0qzNMd6txanOU+xaiPM1Vbhb8R
WTfZEQgV0QxJZOeFwLICw9ZDPylOgqUR1qF+5/dwC5p52Z1uBD7WPwKCAjC3P/fHc9z4QNkvhuHH
+Hw12xQbWi2MFA3yqAJL+D0cSLdE5NWqjGUOJOT+qMWI51dEmqqeuXbmnkdY8s2BI0MKH/60qbKO
RaZeNe4qJLO5DV7suj2UbyRHiOFVOsZIm8Wtt6Mp/VWhqzFCTUwyfYoCV4NWkpbJSnhdFDmE9qas
a1EtIiIuDQhrcV6cdQspMid0LYS8NpqtYpsKPgq3/SABQAuvrn4HFl81dQHWzdPAF5NtlDutYeek
GQ9aP/Xrnb169JB0I/CBtWhae+mXk9SUuRYdtd1pom7Oq7dM9CXXSYdNkcnYqPHtIwzrxHrBuqTw
rNr4ugMuYzN/lP9rMIv0JSd/IGNdrXHszsTPvtNpE4aF7d4ukJ/92+3EXLAAe407/svCaGGmsGB1
sQCnnlJ2QEAl9LJoynr3rh/h7FEPgpn6neJRheV3roxlNLLSDcYDljYmz2HSabLRtwiY6fh8zvPa
SlnWTc5HfO3yfM3hNfpgiCeTbjbtmIb37uNENf0fzTJz1nF8HU9YamAMRtv43pU/+7DdxNQG0/Ug
F+jzDCwQUj34/63c/m1b8EmNMKZUnZYy0gjDNT+5WuGtFV4hga3438QP2xYzoB5kiGfo4vjIlhC6
d4UYjxmjIjXwxgd9Tty68pec2TquSMgwZKfl9IbPFyw5E89PAScvFh1abufYSbvngpFB+lE2yi2o
YRvHj2KqkQ+pjLT0P3ONr6CX0P8kyFTRjrqsrrhS86h97F8OkqIW7WkJjXVcki7V2+PfbLTdY+wf
faovI3p1F7C6KsqX7mDVr4OfTL0yCYAPYcln4WmWHcVHBxxeAixuWAN/2c9dHpimbGsyBhomg9YP
5RmwUE/n6D0CHmuq6s/P9EDIR9JtNSVgRxStvSgcb54UsEioYkwKijGY7FpiRzCdja6GXv1mnpLW
69ezw8Ze4d43vjtr0N4VjkI5pFpkQP4OcsY/Dyt4Z374iT6Kmnbt+6HFqYQcA4DtOC5FxlHx3/SV
RsRnBoJUjxJu5GxNrt+UnQrxY2zazbLe1I6YXi5Yp9QRvTjX3yC5dUgRHhRBGua0VYtAzwULbk5k
ADb2FQxaqkv6pogrKwbq9zkFsL6OtmdpvhuRqQUZR/8zaBQnfeUbCzzWktuIRFvLIU0E/CzaqRp3
M7ygvpQ4oJUzr3p+6M/jgqt34tUSckeS9mdQ4CdHcgI74aCRIuiZdb16YDSNaS2T0VAukqc7fIMJ
/KGUx5fjYHYBNGRGG9veJD6ypRJ/6AL7l6ux1J+Vg8RO7FGmQE+Z+9kE6xGZXyDsjZMtktEz75aW
/IbGxb3e0Mu7K14WzrGoD3shO38l3U4XevdPfIxsj6+9Rze2MpGThTM17cKtBkjJWAWBjK4Manhv
e2qMn4QiW30eWeC40hsa2DFqUS0ESCE1esCk6AGUSX9e6/ffy5jnfVvNzr0dtt49CjCYmu+vmIZr
KVQSSYOF9zexPWKt1JIMbbE5J4xFODNDt55zOqNjIrjDeIskozEXOMlMTsH5PWmMm8bSlI8DXkr2
fV4VoPCFFsMabA5jjBCFAuAeVp/YkSs0/gtfap0xOylx7JrUr0KJl1eGcyVdpzTseMvIL6erGA2l
pQY2sCL6tCphswWkbvX7zWmqRSxQcRTqxGf3q576C2LozQOziRdbywevN84MmAyqTJdzpD0Rjwiz
OpsdxWTRAxpMeTqUbQMXMsuuET5BQoPhu+oUZDSUY+HnNu83xpyhQFjM/xG3DYJXK9MHVyzcI8FE
nEDYlRydYgCGSYjyEBxOEe6p7LmUiIU+5KRkO2P1NxSnrYbpLBja1NIeuvp7DcMudvGdiLbG7bb/
cSGrg0LPauY1B0qHcFRvuEmxsMhAnZLgsyM+/zyN1Tm8jNil1m6PSNG1/dU0Qai4wc0VKDVe+6DM
numfx3NLbazA/mw7Nzj0Kp3GLp9z/ahl0mY7ADELf3Esfc725BTwtu+K26tQVWTzN/M/4k30fj6z
juBfKceAJtxiY2sYuJEErlt4RBl4InOHdJosKvrkiR5wmjXNVcJMaG+Io9sXvEXHJKiR63zC1d+q
RyMxruVCoaD46T5rEmpqb/2kdOW9JIQ3iCRvWm9BU+Ed6WNZbl3lOYG0l435SGB1jsSL6bhT1uE5
kQQeO9w6SxruDa0kOzpNxEuBYfb4XzxLGefHx1WhT37x8gYiRryZkoLE19MhBN9R3GZUkfSzojKG
hgqFZ68igPLNFB0QksuaY4B7Ed9uDD812TkOgmAfVK71TyitjjelxYSVwbTaoikbqeRlBWi7cELD
r5jrlmKNqajZ9TlN1Zs/6NRL8Jfq09/KJ6FzwkliURs5RHfc0hdYB3Le3fY/lQi+kGY3GPCFigNU
L/j2o0PI0adeoafUyLVgrXLtX4Ecq6vKIg48YZVxXgoHsQDclKHswlZE1NkTD+cj/wQAtK7Qye5g
lGnxcPdvF2y6rqOIpEUPznhOHMnBH5TEhAsDv+o8LQjydMxkDZYsCOg2AgjTmQm5Vh/+Te9xoBaR
uJIniH0HHbdvMmGzkJ+JLy/vBFhKNPMmU/ZLj6Li04iH8e/ObCbZF8qjxhulccVDnuiK92KOx8A2
JPKCXk6j+9HcNc1IumTZQYMKSPcUZAvnyf2MMBxgyK5/G+iO4COJFYRgeVU61AWAmgYem8pzwrw4
YYVgVgdXVJtBW1RDNOhnDbbPwDkJdfIRPEjVy8g0RvcHn1Od4J0EzHmcVvItvHFkEyUMsmUO4ANo
Jlypr3wdbPtSDqPtDcjSOE+1CQGBG13KBcqianLWcqKJr5G9R1K4LcZPhdal99dgJB05RQOZg2qu
11HCnK34KwaoadCEb30qP4cu3e4Rpb9k6LT6jVRntVmd5cSDFpDvz0gPjiGEBWOMmE7LIjzmB/5x
1GajnbQSWAQVUCjAkaMeI4AwZ3IibqXizDFE3NDPN6gxKED0ELVxoPc/Na57u/dyVXeWnz/jj1JM
QbVBHLRmNZ5lhTx395hmFkvqoE1lcrMWIKXycf98KN+ybRYs+3Auo+Pc3BnuU6YFR6C42S1JK0oJ
3EaIXCVADqdpuJ7pKbhjSLdE0sH5TjfEw0jWY9qRvZwVRlGYFh1eLh04dk4XSVtFYDh2vTv2t4QF
u3XnIuQwmTcOMKd0jjfr42xuvgbvhzK66grRUV6HFWQl1QlfCgvDFV9psd88huzoIiu0KPVeHSZt
QAq8T1do2srfev58laUAPrKzjx0FpJxfUO9lXIFZDcALhjk3weNdJAwCGVTWB3NljxASSi/by4f/
OSuLF8X4AtYbcAHKLbkm4jVl+GjBqspHJ7tZESQq46J3yk3OsWTQt7XKfrDsIeDTAKwHLqo9jym9
ZyKkG/nRGvKSI/j+KTWuaSZ2Pj876Mr8liq/G6yv4mcq5XUOqyO/9czQoZnGobtURaDd+jGrl3Px
LjwDqRUZ2OARd83NdmhL/oRaBeGryL+4XSuUO2KBEhL4t9Y+pb1KJvFg+epOpXw1Tyq/FDdobNuk
Sphyfubke360AU/Ch7ug5pId9+Hy/KQAsCl8Ap127xrVbKyw3lmOXwmvPoVAYVvqeHJCurMAEsc2
LI7hbhzKad4eZPQtMna0a030Roahq+MYq1kELrbQNGc2zDllPYG798gvRYkF4AB6bjtBwxjvTTE3
GxYBZBx7E8nmzs8aVfglY64Zr/RGC7YZZEucxNnlVhG0TMPNbN9N1MUL52chQcMHMz2XVi5rm34d
3dLI6UJLV4h9EbjmRNc47FYpoI7O8OS/EVSh2eKoGcRO6q459y8Z61YBGjRWynYBPhlQ/Jqe8dcA
WEB4eUxkyKIi7L4Gq7N1b5XcqhmIjRlHBFrmHhH6HBg9gLbDPVZkVUllezXD83ZV+g9L4rpoulkz
qgsZMNyL6pjTatqoeh5cvQgJ0EcK0dogCqG/3YallqjXu4dt/RUqaHiRY0/3EX03a+PYjLOZtlmD
fTt1xBBMPJnoKRkJaRMkNl9Emh3NNt5wYrMZjG7fKO4bLJ0wt7//eQXM4ztvE9CGColOebQuMv3P
01DnlDpK6/os3s2W4RUJe8FzgHyPRRIiadrfFrSd039Qj64PvlEuOnceWM2HazdcAbXdpyaN/ffC
wbV/QpSsLdoriXv16UMlLLhXUYGpEjcBS/VILlquODA9cW7oKXDzdZ5zXSkFXW8+TYr2WfT1arjv
XFlMtCtcGdxbOB+BrPhTkgEp4DWU3qqUSGMD6EmWPA+8qy5/Zkx3bHXTLU0ClPUgmJ38JzkjBuan
lBweofwxZjyUAkwEy6sHr9peN4gXkNqiZInqcJQ+bWzBc8MYiaCXPU8Kk2A2eB3kX+lGhMZ2TMf3
AwjnawOUbXTvbahQ8PFsQDr13REqkB80NZ3EQHXECCf082JPYpIsmznPbHXyyr5rdPb+iNNT57MQ
iC2EgzBMScaxA19t2p+8CtPmmgmUCEEfWtvmcoISg5AJuvT9dd0FHg8BsBdSjE0H0kmkeIABqUtj
gZQefvOfbI9gg50rHY8NkC7jyYe8x52iCUV3h/eIpsr1uoPEP/iwyRCcfTVu7woWiKgVz1MthrYs
1nyrycVju5Nui/WI99kkDIVKehf97BjQhrKmViW3R5FGda+ZIkN2X80wjnpl2iKXE6YPtXSx9I59
DKsVg9jIN5F1gjOW8R/8rCAc2A51EhRstTWu7rE7+cQnYUFiqgg182Qs3PJThA/nXJG7qqckayDg
DlrZw4uZKFU5o3b/coWsrzn5x+a/ptTnU2OTXgddMD6He+WegGIrZuz3AsHlj7vX/NK2MbSawcYo
KqmRMPN6T6SW0H1rPuEvpQtYD/3OUJOWG56pYeozBhfzljEaQ2i0zpzcrmHhLKckukZbkkZowxuu
6hBQafY1qehkR2B9/lUKAReGhBNF6ne2T0EiSnvT45+AzUU6IJPHlc9AO/Qdp0wlGadJJxmcioaP
Bkom0F64SMacS9ZfMoMe+3cavsRwyCdHoTotORdvoDWm8hLdMwZt7QETmWqLowCzr3ycqN5sFF48
Z2JpvjmVSm2Kuwveddpj0gKM6YQ4xdsmt5Hv2WqIkASuYPZkri+gZBa4PrueCp991TO2kE3vGKyk
/Szz5mS75TwDwBXAb4JgW2L9ZOqzM/LXRqS/5nbsy6Ga2v3kLBA0igmwibGfsEYXW13cgw3Gyf/w
36LwIAy/1RzCw+1x5LbqU8+qDTASMNTzLeqyh/9+J41WwBS+xHOoqi8jon+bbtI+gi1F+m0S8hHo
3uYFUXB+Uy3P7/twFC34fT2zNm9ZahuNBJTKsi09yJ+lzkOr9WHioTyxCFgpMU5H2R5CN+6352jO
6CLGJGzC+4R2qN/KKXu2tUrUep7klEcXpHY8oG0Blvu1jFMn5V9n55BOchaKbg56RLkh0yZYsmqu
2kY7+x9VyHmVxWIDuQOb+2XbhvpfhqJhVNasVxFcObbs5T0uSeBVUb73z42k1EUDypezLryUrqdR
HzDxRrmNSw6eiAd0DTM3NfSAnEwrYWWP3XXi0r79w8/NwjfWuLCGqPJWxjnQ9tXYqhxHPo2JEh9h
MC+kWzjVcz37nM0OWDcPwD9f8CentSWjUkIVSxoRSGUVq9Y+MEkb3CVVxModeDscJAAGyC8srFZy
oz9uCMnENopFG43okfeAlfIot+jzRUB8uwTZA9apPNLkMvzB0OJjx/9hs7JB2pNoa6N6OvF5PZQW
EEHha4DDzls4cBJ8+h2vCYB3FPorU7vX88hywZ/eqeEdEaUXsp99WrNfgWxKZTWRXbZAhHeiNAFJ
zeCEx0FwbewR5tdzlEjeTJZY/MFCmRl8cYei9xUFNEIJVOpvjkQhOp7cZjqeSEwEMtEtJkv3n22o
9lFNuzFl48jiJhIDeRydabeFEEIQ9nybbWBV4JoDcc/lDZc93hbHpB5i2SViMZiwNxx7UIAaVdQe
/KngiGp/MP6EiRWgRJizGhe8wk6dQ3vyVSZbe/e8UrVjHu8JRS/9VaNywM4onTYYGC8WMleK82dM
kG0MlPSt10/JLF+4ygo161hlmODCk0OBwrOxBIh5AZrmFXIx2S4kK5DGJAoqVDtIeaYvadye+VjH
2MeeWZViasbr4xaB3uW6Siu72ocHLD0ZniynRKIft3OfZhLyvLQq9rIbx3/b+fakLj6cIJ6W7lgD
z9gbgLfmps/gYEORkgLTY0QQALHvr/wwvRlI6rSn8nMQzxpcJr6HoKG/8fnZXf+PA0yuGMzBzzdk
FKksH875gJdGLe5VRatIpAwa6rhOcFgxQPHCnZ0MjqlUu8Cs57+IyZx7FR6drs6qtm9+fdHbUQI5
v7ss0IeDwk+3CXuIfnxm3KYncCXRRrzPkpbSiMK6DR3LDzjfcrXMBdI783XfBBzaIbdsLUB4nnAO
WLcz3NwlHEAyAlP+Q1qGZud5LaOSCaAk7T6hfUwGFIMuOHDeMJuZSilbzKIzKEzrZ2fmC9usZzYt
VEA+DdRkKswnJ3rayK5M1k9WH5sXhXIX7GGlkJ1j25525iV7a06C//hWDeANFPjPM9TNy/BuGKZU
NCJYgwmShZzwt7XxO6HTU9GffAg2zk4t8+TYQyjcpY/wA3M+Ulx9HSijxoensAlukG52yVdg0fNU
uApwkFiI2uoFvUUgHTtQkRwLqrjcO0KvDqeOOe8TeOQx1IPDQIQgbuKMdWaR2exNX87W/Z9qaHVQ
Y4ggrkl4TVBiQ7H+eSEuTaO2onXboLi3K3iAY44j01Ta+Oh1OKEN3H6XdoOVxBOzZaxnE88fzsqG
8iO7FeLgOSASXWcWDAfntXpJTZt7jZ44R0MY+ICloLE74RcSdXVgVsH5mT7OLnfZXrvQAm8OOVHk
I0GnTDKA50c3m4OpW5wIjp/SE8+z3pxY3O5QbJE0lCzVknG0DwaZH5v7JzAxr+Bgzai8/zFPZxXb
xHVq40eHWhlfhEapuoc6NC21SRmlIkgZsj5l7+Rr4BFjGPpuIeOjGzJPaiCSEGBwpEyJJzdL7Hxm
NryYQ4RKUyg0CR5Dp78i08sR4jex5YKNnZi0BAKwAyDklrr2GTCwfB4nUUwa6Ba8wBC4Hzpdx/5e
Cuq15Q8GGqEtb5GgDToiYfhZ4mczorv3/J3z1kxYbXJnMw3SJbG1QZzVSe1BKOjSsMpUrdj61n23
z15yhWrYeGNZ+xf9veialfB8MaVd8RXjNpgrXMlIAtQ1UL5yxldS1pNwFsTLeFZbTrMR8YTuFilE
xAgnpVQnPOxxgaeVvrUu0cJCPmHI56NC0RpL5hfmn07fJj2Eb7+y5l5Y2e/8ZBdKZyUwlAIvpcxu
lfHyWd/pU730lBgx4+/4pqtbcRDZKkFKchmpt9nm1ESijJUw2iUljgHVmPNHDQM0IKAZw1hCCgb+
GSZ60RjgV7w8RroKIl9mAyxFe8WRvn+2IJutdxbjXC3Q2MayoRQrarbVlPW/PdFFk7laHLkzh1v8
FZjDY199TRrjtmuq6a4q5WipkC35FgdJFVtM+vlub8IOw3/xjs7dH0UrSwil+8XhVPNqw5T/YGXG
juaZQYFpOEUx0MmgxbVhuQEGV4y4LIqhKcpnAkzNn8LezBg0mGZ327Dl3gj/9RAvnuFdLUNzHy+g
Xy5asLlmiBYAsl+/9BrAQiWovwd+aCEbXZ3q81yDJWg1T07SxVyaOr0dqm1rfQ/j3dNxwiwZ5hbV
U16+/esJrgvWbbViijtxIA+Q/YT3bwwDLvtRq3M5WdJHrmiaB5oVbhHCjRPG1UYpldpoIXFob9km
b31U5YYZhGmU45c1iAqot0+17CKZvgu3J4R8vTC3xuxkIwcBXfiENX73vLGlubP6IZfKWuXz+a7y
lEGzConm11SKTOAM3hn/Qxy3JChRBGH0/LJPwL49zQOk+O3nkdHik1zhoOGB5nzfnPHHR7opglT4
kQ8EGaskdsiVY9kgissadwrSwHv72Yfp9NaHZ/JNSwraH87aa/FqdHVl+5DkTxpQ5M3zfg9/8mu0
Oir4n6rEXsEYDsbWxyDF6cvZoFwSIhFIj1Ex5AO5+8d6CYbPPMtik5Zj9XpZASSrLMfeTdDwBRNI
r6zpN2FwiIal4W/ZH1/VRoWD+iXtaRLWt9NvNAUIbGPSgSYDpNm/Z+hA4ey0IWHWnmXNqPFcQoA6
MqnxrMWoYDT8cARK/NudPWxZeQpKbJcilhdngX60ACcoeSNgHFgtd56SwOrAtz4vczNSDCF8wGAh
kehvVPZ5GHaVpozHroYUFb0Erzbx6j9f+exV+zUYEZf7XW1Nnge2i1wnX3zYMBv/is0Sfn/bNvnt
2mYobyS+sJRx3XKUG5BxJGMef0tZEStsRVwp0PaNb/B4Yq8ZJUpU6ciyPVNpQZthF9h52ACl+OxU
y5+5r2x54pP/iH8t+slZ7Tnm1lg/nZ/blpn6/FU/PomDZC61WG88cMjsKUX+GEXbvavcT3Fo75gz
yK3I8k+RKiest15xrEsR5ri4uQ/PvNZrm0mMEBgedh4Z6epfbwwnFl6fnUtgXTCGkEZ6Av7HubBo
MuCt9xDy0Huh6FEl0NpRFAtT1webGpiINg3XWxuuM1O1mYdGSRreawKxnZeXsXq7n0gBSaS31Cd4
BRexoQn8eTp1FENR8ySMMO5Im8KPUgSnFUM1+vhT72qSEnBDGB54OYrLbPfutYpw3X8xs6XOZotE
BWCFaEBR53YphtBQzXWv5GRxnFM4cRbG9iDsZ8chhODBNS5BOlhvFFcGneS1Fvl2Zt2NB/asUzYq
sXbVKOhOL55v/gzHxAgMopiydsOaM/xVAcdxiN6K6fQzJwH1sWDyzz5jOdcta9C+RUUl6g4Drv7J
rCSG1e/+4rLVE5Kskb/ETYpndw8lSGsNMXsAAF2nrNa4zVLnp/mfktjEt2OAHhdOQ+0SLICkYdqF
CcLNMZfJEceZF05NPpugE38m/L7jRxBmwC6kJ5XIEJfgSMFXwYo0GzlIlUkO1ZdiZeUecmFxKZJt
UfBMHeabOOQgXTTPH9KdSov5Wn3xJeGmevP9r25hGWRRZ52F/9pHy23i73SiX/VV58t74NUikg3a
sjYuUoTNHwSYAVCXOdoQxeQL9ryUxi0xh9sQ7HlKzVqAljiKmJwtLHyxn7wZKM9PkAVyr0Q85Bpa
q/fGLAz1dc6l1Om5XVohNIdG8MzqBkdhYfCndzm8rKPRjFIOLUQJtgxXHW5AoZDs/OVUsmozYED6
aPeZ52gEZv7CPyEA5jIdWN9CBSokDantocQ3d/o7KcRTfVSvWgK13Ose4jCFVOdcPaZEEy/Afn+4
FH/IR+4Fjm/m6t69A/j91y+e1bOrvz0N9aBL6Ks2pPq9d+KW8x2uDhYquqSs2sAEs/ahGIhlPGT3
BkiGylQAJ7yA17ZlK+aNVm/bv1n6yE35PETXnHGDU5Y21uEZobzzHg/l86uWr9EaX5yqspq98RbK
jPpr5hhAN0e/Suv7E6ZkQCoq6pVd0ygLOMgNLtiWtC9CvI3E46kAh8UsxjZtezMYGRqGlys9UCwB
czNCj+/DUt4aBv159BWPGwcHsJ91ymfdDDCgsN2kHh3ZInAS15cpn/bzPu2bO9z6/61hoWNgvT+x
RO0GrI71HPOILm/3+LtdP1TO9B9x6QFZCjtXcRQpCLmee+2KbgSDFVW/ZjFPqQjFt0witN+wdpL2
f0VxTocoQ5YZaI7G+d424ARC8x6ZCVJgWVQkD7f+f/ayNKfL4ObTwdXaY8qcn2eFwXGvuJ72yVnn
EWohbpzLDNQz57gtwlRaW4tUpkAjkLJjg8f/DhxWUelFz94et6nqB388oR/CvEDSACxUdjO4LPfu
zaI1uKgxO7FKMyy7Gth6VxRNSaMXfLcc/36kVuHW+ORS2ETuXB67m7FAnYFuEqvJDWnikulciSs4
ZYyf2lTueyv3gvMkFZiZoVH8alAp6JeF+L5tu4xOJk9KnTMXU+u1lvGF6C3sxz3dgUa+rP5kYXaH
/IyCSHIZa3RPLsOV7igCPyP9PWEOTSurFHMUSNmwQzzb1cHdiLmlDhzrcXkSrg9/xPHawYG7mFhl
+C1w73IkGr/wPBwZSCMfADW5ueWR0WXxU4CBBKxgBr22i1zRZ2DAOnlbvpkEb3iYxO+SCCye3SD1
OfwYYyXSCRB8oAL0k100tZrTZflJONT7VaLXe4Kz7MJzTy0KihN3La6hrmwB4SdJXxNDgYE9TYYe
oShaGwDflzjmjkb9wjJXOn9jNqFg8OvUWpfQD8+WTM1OQpJtblllqVgGQ1uJJj3DTVpyhKMJm/bw
+A4IaDHd3r8MnzCjlWK92VDAgwUqHDB/okDadsnk6BEiCNktXN10w96mu+cEV/J7TQzUrQy4f2OX
12EIluc6bhikL50E5FMqxLpRpf1aIgb47zhLbctHLmu0O5zhVb296KKnrbkHeotM487q3b2bl9kV
0SDhVcbmIXBUJgsGpRJSq5Hv+9BGTQdAJRFFol/0UdiGMsuI4dgbnV/3uJw3lwr0YSz5sr5dSsVP
xHZDzpKQUPUaXnGKJHNrim/x40MLYUD1deqqeuX9eBrJvgGZ8jU44GW1V3feYrtHAb/8dinBdpua
I6ZHLiUxJEfo2CDpAp7GZdQoQdJjDv/fWmykjbVF/K28SCbHEUDKJxtc1MVkOITKar6OlXrEkOl8
StYQtj1xevbGL/IkC3HBhlufq2aVgLdaPCt8yl8wwgwo0hmblGjDXRksokCwZBc6yP/xM23RaBQK
dF1USfy4YcFiPhNncmBxsAuxTTtnPN/h/ixJF6StfV5LAritHkNI3vuF/Pk0hjRUqbmrI7sYIV12
EzfCX0PgUGWz+1pGCKEDLvmPyWMTGwjpTaNjFEvTJYXykNOakwToRTNdg45M5Of6/hL/6w2tEdxG
fspTnrC9WXAN61wJfLIoCuUlNg0tgLoXqpS4F/GSCNDAjK5K/NvkjYdU89j5FhmgWN8Me9E1deY9
9GI1HTnEoPNG3FIWQCVi3ArVRENajr1ydDGCdkqtZt5QyxVmdMt4mPDOAVx7XPCtJ92qyPoMSVSl
HzkpYAfMGY2C1TJLI92ORgZvXpDiVOo7Qb3MnGXeGThVsLeOZGzf5ofHoY5RkuWBzJuke1YDQlAK
7/qF9BGodP9wkg13xA6u7Rud6hD5xTSpju7/rzN315dYO4vHkSIopExnhBsnBV00deqh6QsYQEBa
m9d1TmhzbmK9Yca9rLtE9VuPY0/bKaze2oMTOhadgvG2C3AYcpJn6RZhV2/rV+jHc3JHpyRNFi7N
Y8IKRlOYi79RQ9ziuSI8Bqzrod1T2e+t8suokey6A7txdjW+/e0U9DCfXMcye5TFB9JSSq6XQ4Su
HGHd8asgeufzuLSjBMh3nACWy4QcE4Q4yfIsLl8p89QT8HZav5NoKBqgStbNwxUSnbghibZpplEa
IsTGMDxrY5Mq7wOSyTzocuQI2QpkVr1FDpmjhzD/XfiQbL/tG2z/FMBlgRVHCJBdF2R71Pz+woDo
EAf+kSq/DIRARMZRt9ud4qUbr9z7mRT2+fq9/H+qtuf0hPm7K8qkEEdMJc02GgNd53TTqsr2zTID
46I1PSvWz3r4nUXakdIimMwk8IRB8TQP7jQ9Iac4hblxu97FmwWpvLgaB0C7SsEvoJo4eMfPlFqw
BtiwFRjUGFL7PSIYyvdwcqymtuIfQXiOWsTF59ldOc/qO4CGpdNtG5uHjsQln8hIrlXnvBLeAawt
dRSVL4M1L69WKuWZRiKih9WQWaejW3W12O18DeFTkysitdFaTBGiBjwbJw90dF7poEBXZCHi6GoA
8jeXN8pgggFy6e/CUnE6woRdxnjgc9K/LFvHnZH6zyqm66MqPNCDMiZRkrDOW3NtxCE/xZEjQoOK
y/IG/xQ/kL/ZeIx7JKL8uS9dQzNYfl3HRORXb2+vpw0YEHWF/+sR2LKKS5KVUco6eJwDK8KqYgLO
hvqCXonRm2VBOmM1BV59UfSoha2rkDMSq9Ym0cia6c+ZnzxmKPBsYLFCiYPYbVr+AFH/Y1mcsdF9
RY0l73YWMtr8zUZUc+cVU/B1Vtmg27mjKkN3Z3hmGDYCuDWKjad3nxFGliyrFHfHUV0d293uN2/j
hqCy1VBiss4YX7eD6lmA3ezPFEZXHqX9w64rm4J5z7DzsG6rUAgGW8S2xC9ghOHAnKqqzZ0ZLfQW
PoEqQjpBFoQt1xFUu0Q+SS5RmxulIJPV4ZlHS9hMD4MgLsQS4lHroWRmUsvFtVewGLav21GPJClF
ylpcEOXRVcYf8eNPBbZdJXu+KF+SD0zN/RO9xa8H6l3otA+EU/qzrzqHfPgcBat+eO0U8S3/2a9p
t3o7d8tgmNlNIjl2eGnIl8rOwW+c4IFGUmUihsLTROb3bjmo2byZf5/nf7hDjRNXv7FCoKcc1IZ9
u4mrCYJXDhP5748WovsOzEOvEnBD76f54oan0MvzjXQ0fOaMrhXagw3R/bVzmQrVPyWPfC4PQJ4r
jg25x2OuHAPKzsvGRbhCiRZ5eG9JnkptIwPaQgmyaEywNrBnZDweljYDenahCojnnxZZk095x7KS
ffpvDrp+a9X7baIhPogty8BxBQ073RrGO11xorHO55cD+dECCS6tO3NE3ZCumE8hZyqNM8N+2QLB
3R4ycRDdSHCRo6da8OznFn1QgXogwLYUO8igJpIedQGbRfWB0rCt2QKL0rgLVinukTkiAF5p6i5v
9mrPVDXylZ5ob3g8zH6Y+flN7ZRh51G7aWr/+ynNT25Aj1aNB6zz+OoJI3hsbi0aYST0zGJuNmnW
X70prVBe3riEypGk73kmoYSrmXM7Kpt2V3ee3q9lA3cTKnpL8zmATsiEy/iu6eQhCGDS0nwaoSuB
w+RGxoOmoKE6TT6UCIU37iyyXQmyFjQ5FwV6zOujqvt3WAth15ALORLjsU8z71CFjfsDfR8CuR6h
hx1VWfwAM7XI3RVpRPIJnzHfpFo9hvYNP7aYbO2clHVHOfxOjRmDa3wsAqBvCi3Byt3DvWIz8EYS
RbrKKeij3OoNfOZyokkVfScPGaMX4PyL9JdSKaoDuuuLf8NPPVPH+9ikTQZEXYNp3/hJxDA4I9mx
6chQONkYyRsMZjbLMqtCKTLzpHsMCWU/cRWVRMybxf2WXtUMSJAqH0NljCiKqo/mF5peTro1CJ16
EGpMJTRAY3mBTsT0m1P4RG8s3u+P7SIDy8K/B2ZNt/GojZwdBnV0pXrfg2Rmt7vM6TfjmJ73gkT+
32MfOjgdVxF682LIQ+wcLX3Wlmc+BvB0KyP97XE8JIp3EQsCEo44HEM7a0fcWML7VamTa0Oy51bZ
XfaPATJBitUhhe4VNJWsgiDlnRjj3rB/LAVEkfGUvIxJ9iFv/ZUWQq/2qviArRLWLt/2/2b5CgxR
AOGAJ0lb7J/6KgmKmqZLil8jjYE7j/7vZNneu+CzIYJiZsU4bLZWDNTuKDGN6MS1bYlIwlDEIMdF
sKsGKv2Ti4qk50r0ZwfXDOj/Cg+o96hVzTKm2ut7+9Ynt/drBLcfbYTNlvqT85HOv2wp+/jSrlgb
LcxzK06n4AxqhC+6fnjDFPYcXtDcminM3cssM9G4BImQvWPgJFhnjoXddWBKMRjUFcpSOKzYgHEL
YKe3xYeIY9wqi7AxVH1dBjc8axOHQpWd+MKRdHwHVnmmtfDxcGH3L5vXo5H2fGQt/Czgow23Fb97
SVzaGBRPAKtb7zaPe471Qk8zgIzN6JXAXOlxwu+5SKmrCkpBE0Dx61crF5UrEAvIF621noFqvrDw
xIUtTmq0pMT6klR3Xe5KwqAbM3KRQ3RMkL02MhQeSrDkyUsZHCSuAFpN2OBjfUtcQPW+9q5z95rV
aLjPVpkTT2yuqyValeTYYY8Ro7DWCARZ1urjVTdqW+tsIF9j3CuzcUvGlwG7S8wzXP8hEFTBohAs
zYmV4oduhFAgqWBIW0JEROjYBFmbYyPYdJf1mi9LCXIs7o7QbGCC96sBV515NmsVVOOgqXrrfX5q
A4jq3LWTr7yXHnaE3nQ+NzksH/qXZfkHnBN8tcwZDZUBDXZJX8QfUgi4I/+jnqSWBLnBItR3qK+7
oJQWAIAkxskRB267f+fMt2Z2hn8O6c1IzyASrDMPBa0jIiDlOE3I6FbkTJV5vwRhxrZZm6ebBdoF
CkbOIRYePc4CA9rv7WNUWjrngcahNuyqy+wN/cNblj+jYfaHnCDelGeqID4KcM5XTQxrc9XGDPQp
RdxI81ISO6OFOErWSwvkrWjpOEKFIKeDsiQpBv+BIVKZxxf1EVv1nvN8/Ct10+ISEbx7yy5BsWRy
E0p4YzqpaeTkxYDWZhqqnPby7ohS/YBdniyrkomqD7J9JyQW+ci6YhiWnUfbZ0Mr4FSz96PpTQN9
erKQsJ0qngxX2ZXyQSoSS4aZbFLTViYgjl9kqAJypt6EMiw8iLtUwnuTLhfopp0a5gtGlUCskoXg
+Loe+k11l0MJ81xXLW14JJjU09rfaNwVYUKhxK+wYMLxI4Yw7HH4Hcttna3vCSETspqCG10VmIsB
iZEF2JLBGI6jf357vvQYdCNdZPnzWz2Pfg2Ygg21j8Fsttzb0l6Yl/TuI5NsSN2+IaL8Rx4MgZSm
vOWU6R8emgvTtvOsTwCuaEamTgHo6UanjVAK3DZDW8hg9eKTswVm9U9Zxi6LAAfelz0ZSMQR2crL
o2hALzOq2KHD63xCh1u0zKCUFA6I98zIvdM0sjl/Lyj9wjD9jM441YAVD3xqZl/vsS6eQL0x/h45
zxPvDbUI8VwOegtTaCz8TpMfLgZ9UdXb8bIDKEItDkcf+yAohb+/Iopkwlzevmgn+MYbtx2tilRl
wsuUTNiFfxhX1xbvNLNxf4o2/sgHo3Q0NtesywRSlU19D+NlxsizVCXM9N0U52ixkoQZPBUP0J1B
s7idrgUhV4dzg87cbRz9Ls0GDPa+ThtEsYthxSzRJeLFY6umtwcyvz5NevrjrVoBHXv+n/GcR/fr
DRCmczLBmvX8tXq3dfZDJlMEcBq+f/77SkoXOKgz5vMNQU90kIbwEuxjDN93Xh7j4xW1CTJJp2cY
evFWGbJQC2HgUsUiMDyf2SWYi9WyLecH/HgODhO80oJt5FP6AG15S2833gBwLzEwSoLdDpcRbMuC
c9wXSe0ZQ8WbNniTC6+mIC5LMglcrD95Mvpdyc4eVsHpbjQ5HlfyeLG/049xuJD3eEutJvg9fXiz
1GePxmjaa0NKZ/fgqiZfwjVbrHzVMa+v8YC4bqazktM5pLYpcK025FiDwDUw/omXBPc72YXyIhCl
68KcmNqXbg47S6vK+lqh17Z7CeEjtHXrDmDWm8fXWfhAT3IvIUaYplwe9vOfTWOz+1TxrAJ26uCm
AEngN3PlPIbQJWfzg/i+9eACTjLqyJw8PGI8SGI8TajbQp8Wgg7+eXlIeKORQYFoKm73ohjvzOF6
YJ0ds6XFczcIUTKAKISseYRQvLwOB5r5SnvemC+YHs8HW3J47VQiGGe3the5L0AtSL2wfH2MrHz5
2sgZVwnN4sxUUF3AobMqFKrY89BW8D1+/FWLwT489s1GjOMCGnPs7Ni/h0a97vNzCOBlPH+swRle
mvP/WX2SAr4ecoo8G9vMcPjWZNOin7G3tDkZT90DlYHV4SdokHc5xabG4K3Rk4iJWiLbmiam2PSb
6F47n+y5i3UvQpHwVKb9FM6wugCKTFP7MVP1ZxG2hlFfMofuyKLE8qINIjHZe8szQ0tIqBqQB/ob
jEbRepI7XLRRz86qGNETlTOCdnzEkwGDut/H8tFT3sSeShvQRbPSzXu0k42gt1/ZZVWDoTp3GRRS
yM0/+JACtyYT50jR7ZN/2CTnP9xbQL1mCfHR+Wk60xKtBPrWfc04Z4NS/Y9KvqkLGuiF+swpKma/
k8ePpXC5qcy2k5HB12qixiHn0xOeD5ipi/eHCSkdZtbVLLtFGoFgeYK+ig3XAT+6w+EN/WDNR1GK
dXP1AHTPt+ctT5p/UBggpaBVlh/NvmO2erTg9PCbeKhgDgpalAw1vOoK0F+6gbenru76IUtlPz1H
16NLUePVhSLhpVJJ4cnHkCFPt3tOYVmWvcizB2QjypVhoxejWooxwpYGK3JJ5QxrTAq6xG2w5+6S
2tj2cAJV53q31XOG4Bmmt/gj+bpjS4mwptfhDfcaP1R3toDRnaN54OHXMdUY2NJS3Agbnz43X6mp
UrrsvzjiIAW+QqfebGNkz8Rrhw7PO37yOkcTChlVuFCr1OH9Rr4obbSt9oYy90GHYoV+H9Rz+svL
qT5R972ihILY8E58TLq7N9WS6+AxiyVU+KvcXg5JJ6eidXe4n5fQqI2pfyQn9c5OH5i6vKDUpEIO
JAlR08RgeBsP677LimX6xUxrXZEhBCT6EvA2LejbsuFaOBfP4M+xi/ywXD3RhfDhsiQjtG4ixM1z
y8im5zv9EVBdGVf+05Go6PBl61w0+yg74nlJyqtgmY45lrAQT6gLQQacgoSyM7KzxILs6ZngN4oq
qrYKYvzolP4vmJ0mfXoyTcFZ6ZuA0ow5I7Nq1TZvwGXaAwsCTyl+aHeMwhXJkdK42syIH/Z2hq5T
n241bP5kDNUyZ2JCKsifkGckIf/F1kb94M1MmTsdEGHpenv5czt7NoUBQ7AMQ8uSUyi5icM7LZod
Ru3Du3CF8RwlUvHGJscVA1/wWCiGRSGoA82W78tbKom2/zf+RoQw6hOkY2VcQKpBXLHdHkyJq41E
ovKlA1HfD8pZPZuwibzOXFG9mgRr1Ou4nIS74pgDFKAZZa7gTKiTdJ/PkINei1TPH47Ik9OxENHR
tG7He1VZThFmy1Nz3wj8ePP8Ykdhs+7KoQ/5wzzb9k/ItsboC71HMndxv6YpZ10MEw4j43rtwHEd
9w+8BxiJ/91Vjanw3vkheEVfobu1jRw46evcBK/qQLKVhNYgyZvm+SOPVMWezxtCarvA5ZR0zHXO
xRKSCGuTh+gE/ZmJtJOcdog0WGr8Q8noiBiLJvBs3ihOSDZ1ykAgDz41S4IxqcVUjRAjOIKfKZAi
K6/aIRLwAm0H4RZz3nVP+1x5q3iBhcLgl/bWgnttKcuuRymlFiszm4z6s7f2wNU5nTeR6CfbqX2c
aLGsGvpuTe0ZZ5HUfFE6J7xNWVZcRQZxC5yZmQDmIF1SiY+U6V1y74ejRr25DcCQ5LPiHKzR/dyu
fhWmNOs3z+RCdU1MpIUDXGQkVIJWrpm3YVDgGvtgYMrLG2DPkV7U2rxILUdHGoV8diiMEzTw9juI
66h6TxpVMTBlP9LuM6iKFnde8Nn5lVDxTXbZMok3c9cJ8ycvwTOP3n1sZcJoGIePnc7MBFOoSzaH
CXdcJM+S9/xWZZh3ZrI6DSUwcCmaJkxwWHQaxPz4SjhOYMWahJ4QjIKuKF80D7i9b7PqpE++0Hh8
9F2QK3yZMzN0pHK53dP2/v3kN6aTEzORzugs7QDvX3WIZ0kA/O/cuo8FgpT9/5uzv6Am8kKmUlqL
63PFNLcx0jk3rc6YrzTTRtrKMziEW7fRrswrwn2w0YsJajyNc7MAckSFwX09R1P/KtJLzAvCQqr7
W0NLI80dnKbHBeD+efeOBj/cP9mZ03LkhHFnwSEyzb0mWeJ3DIEIXZdruvWOaf9HNQEIL/PinUeT
IpomcpaGYWJecR+TaZKW+2QDnqh3cQYIFVs2QxmUvSDLbuQc5c/LQ+LxWTTFhSurHfr7ZWjj93kW
yO2UNGFoqWc6E/rBg37fvEj/55KoaD5vIYH54UjfR9d80FLtphW8jQZI+BMGfmqe9CAw60riUs2o
OFQ+7ZJrxYUbrCLESyJ8wy4pWcNCDnGVjkPe5PRZukB+qkVQIbMsl8xy5EGASPJKCYe873FKPQkk
HVgQwd9VULWF7EfcBalyzcIDVqS3Lz42GWwR0WcdLjktodI7oBEDSa56HP+qpEH04alRfbJbGt7F
qKVIi3N8H4aKGkioync0jJ/SWxlXAS05o0mokXbUWiZxZAHW0EvGVGUcXXI+6oxaTvrM9mfRjg1w
kvPEnt92xzda9U/JPuwbN2cvQNOsbRyO9ketJhNsUvtW7Rp12s06r5tRkDSxHuJ5HWOwaTO2h+Qz
xDmY3LRw6xnd6rtvrnURJBPAVtEEY9FAAZZyLm9nGXCNagEU9aZznEna1EXA2uAn3KCHYrIqnPyw
YJH3x+cgTku2agotRXuoGcG6aFpLpemq4yAr03ON9dCPqStzUwOtaQ37dsSP+UzExtXCHmwqBc64
3nQwwu1mrYkyVrWhoGpdsmdm5CqARMydKAe47n3I94meA5k7agszIvDj6Jw5asjVVnetVEh188po
ROEM+Pd89fw3ARP8Qc5v5Vkzcwk80MIYGu3hciTpmXrKAAtOltCYLfgGqj8XOWzx/sJbf4qeXJK1
EsjlP5YZ6ZnjWfCL5RoQrc2Fmf3H7ABtzm4YXWFpP1RBZiS8/XzvhPP9N6LRbDljT4F2oe2X8kqG
3pDd9dbep2fLkDutuoSJiCjJ0SI76+2c29Pl4z46Th9Z32owRypVoCuYqzrs0IgAEug65ujT5Au9
QivBYXvxpBH8LOGQZ3JpUw2Q5L+DiRhQ4NnNX1r97648MZTTo//wmj2XA1Wrj1tvJp7S1qB8o4G3
lFILCNTqbQrsUG5DPySEDEn9XbZFc1Xw5NnfYE9c6xoFvDfO82IybmtTRZgLJITcqm89VTDPdhbY
2eITDbnGUSomqQXSItS8nTcV61ECwZbBlnRr76hJ1xTlVmnFJxm5OH4LXKA9q5I1yv3/587oomm4
cZC74uAmpzB3izyoSFdp/cPMXQfJp6CoXENtlFJqprFNkr1HgTmrEpkcAsp2zHxGmHLUJcX1l205
r41j/Wkux1fklZw0jaKOYz/+8EOOoo1Ndi3g81DGL/wNVDbJ4fC+jcxeDwt1Fw12mAnD9Mf9YvDQ
AAAOWQ9+bHJMCLGXrkZ/Ejav1HsO0Yjo3/e30GmzuMHecsW0EDTZXxKSnpFvGB8erFuiUCdQ0tnY
yMafSHiLyjA4BLuiTxGUprLWQwzeS4p46oXorx52IknCGTj7yEfV2mjurcb/6zZwlS2VK7KNMp11
XdRJEbkOD1sjfOlZkL5sWABzFrvyHOieLB+HNmDVzWxCBigxQPpO4ojowEJG6TTti/Crm+zHv4hy
3VzROSuEg4g75lbPnKQi/I3d2JYL4Fx+6owIbgG7LZSqCQMgFSnHrTHHual7b0uCl//9Nnt8OsxD
sG8ZJBIGqlRk+5dIBqrtY3+5og+AD62sh0WN3siWP/GDgc/nTftoPjCMOuREQiqJDcOOtJVVT4y7
JA+VLAyK9iO52VdspBUejkal9hp7dRovePzUDDsy/2HsH0WPh7p7dqhLTlhxGJ8rCkuuy3Bq2Bav
ykY+VxE1qGsNLBlFEXigJEvYjZgPP17XBYGjBJkXf8GNi/8m1xH0VWQa/m6XfXxUG4dIaKL5ML6E
dMeVJFvM1Dm17DgWvb2peAec24lVUgq+iFPq4WyAdV14Q7//RtWGZVH0CZuA7VA5XsXkOtxPpOVT
M6obgGSUbhg9h9OPCwPO3hvEOc0OsvanvD5LpMldqpJxJf0sjsoa1DEElkZuCQYxjiYwUsFBAXF7
f5lnSRwQoO2llA0cJT2+IbhwKIwfbXhqUufPdTlhCe81LJxl4WJlg5jJJMBl3WDhdmWJZcomHFDQ
OxThA8tXRTg3ssVnqcuRjEHckI9Xt9ZnOFoK18rvZ517gx2yaCg4W0PoujvN3ennRIWtoLgC1+xP
M/haqCHk/OIIsYhudi6cX4msdKPwbmzvf1J5FB/AItJf7r6UM1wfIcOKhEfXX0cYMbcFI8hBqY6/
6hIbBUG4Rrzva5sKGpGk1/OPVC9yN4B77nbbfblQ0tf2yPbGukP5c6MerQw27i+wMb9+WzXk+YC9
GIoSYzPaHitlQaCOP7ljGjc2ze7P8kwPM4OvvP4PVNAUr6BldNl6o0wIBhODqVQJaYuMJiBK7QDe
YpFTjde4XFm4aU6CqDuLKWFFr3wFFA5AKUleFEzqTQbjXvNj+NMWF7QJgiRmOhgjT+NwYpUKOH+t
yiYY8TsNXcw4tRkRvXONn8fkhwYV5u1Ih5P8fnPHbrfuNFiUOPtFKpSOA2E6Bn54xdJRIguwNwTp
uxAPoDEYVWjB0vVH276rLBNnD6erD6YriQrVKdfnVqDZfguf7DSjo/sHaGzLnfEays/DtJP2p38s
6Plmy05y50I3md9tV34dEWu03T6HGkoXUcpKeihlVbdCT3462XIZxXk8Kr2KOSTCGuYKkcCmeHbM
AHFBfR60etDqK88CsF5LqNmpAttNfn+0XhqH87H/fk9gJ3zPNx2SZJcVClPlXjxeOHagefmzlgy1
UBGhnwDdqIsYnacY27lej2iJ+uikVPe1rtqKlXVLAJALJZgKhNO3D/rUCfocc3ieT/6rCphCIeBq
upilQnRbiDA0a0DgrwAtY6iJ+S5RzKF+4GTRsEVCExx6K37EkfZxFkg+bFvWAs+W7gjFD1GwPYb6
FJNNsFaQ3UKmEPKDc6NX+MB3Nv0+ooCo9hLECNFwfAOmOsbFzXGmucDZeDTsyOuEj8etBWOTvOz2
HO0L6oP0aE9oJ8wO2MWNNQAWUWVIQD/MkzrR7rkD420PhY2171Ifp4ZDjgeYjiHmM7K9Ry3GwXEn
jHJF9xOuesN07AtCE6KxSw1mo+HZ2bHmy/sXpcAxWbZ1cyxsuQ5GwZUIP7gBYM+RS9kI7CYn1eGs
bE78m2vUT7NkemeQbu076NfuD7LENwWwOj8oLqdAi8/k5OjZAe+O+klU+A1LbXSHlfR2K9qwExW7
1SyKm6RHQtCkOZe2AIGQ2S63JF7wc+lNR4YIc+gPhiaZN1dKJ5LhU3DxGd8uvr7WYNlacR7w72jn
+jlr1S26m2Z9mrqllJ5xL8zpuO2ZCzZRU87MCu1vsTVD0x8wQvRQfCN3uFiHoIWsEuEmaW2G9Zuc
46rVFGfra5vWrvEQPOeDwVcu40IFfEFruEoYeY6utZlLIIR2d2MHFSHh8yHFiQ5mw195AIHJ8DUM
qIG4Rq03TBCgzHgIekHdqIgJdmQ2jomTpbb4Fv2x6JfmnrTXVY3XYxEhb2I472K9xvtWnw17WxNq
ydWGwa7xpZS/Q6n6XquwxDX7ulCJtdhyro4F2LseIIZwa2g7ah5gwohsVO0a3pxrpy9WSzt9I4Qd
WUpGvMduTW8QwJIQKZeoOkTmDIGlBJzpbRsmMKMqXsvj/jBGb0cWyHj5I23eQMF8NRLwoCdUN43y
1yPnghZFUVoFenPN+NxQVXUFIFToyETRbgm2dRozPYh4HXYNub24m/HX7D6m997YMLzmFHlKw9UN
1294+LUsZVtm8p5UpBm4YSBLt5v/eFWZTnsztmFgBHzgDl67kBkia25ATVtB9Jxh+I3jvDuht1UF
ZQXzVT/73WrrzCkPmrmWO08Jao9x0QU7DJiF2bXGHyBio45cjudMHrYXGX/Prs2kbAcr4GIFKF6v
duWYEsqHEBB5TWtbDIsqbz5FJ6mv7DxJi73PQUk6fPkeK+zbQ8OLw2CmhLVY+yIEfvNpjVpq+Itn
rn30f0LYjdQ+jCTu5u9Wzeomol5W0TXTJoTB5bhU+l2ZTpnuK/XvRQE+sZ0lY1dkXFC2i4fzKHTz
uzz15FvMgUgzAZxHDLj6YXisTSS2SEXS8c3IANhVB4tVwMVwmUV8qmX+dQGFJFM4ARRSTB0Che6R
WPlWFQake+0qL5kMja2gz6Nv5e/TMx15IacoKTYeh8kcjxc4pjq8Cd4vezo09jJuCxvPxxxdguhA
3+49rY3qA6DYbvaT7zvmc0/Xraw+1y9bKe5/AI+eJYhGP7hGqPNDbW/sbKLcz5B5MxnG+JVUpad+
YvB5BjDI2S/OmCJz+bQvltp2eU6/wud/akDsNL2wa9Dxppg/Jt8946nleGPuGvSI8JBW3kSUvPp9
pqIVznXTJJUe4yiipzmVWP/TaHuJphJZFhIeJV7AxudJ1sn5Q4oob9IsUjJTlLoownePTYWwaEMa
mvK4NLR5ZN4JK/uMRzwZJboMe5I8cb6q7fCQrsdVAyMmGS3cX46h1ZTGw3Tq5L2nP9eibylkAuKY
lkXF+nTR7lkXf62nQtl6cgZnSCGEc0vJxMPg9LiBamxVFsFwm/VqM/OWymOn6wrKwsfbHheVU0us
j8P2+Jp//8x6QPieMP5bqEGzq85de/xkMsUbzce3y5xHh6GV0VFb4m9g7kwEb1QIyVbR+l+F4uDO
73LVTkvSW1h0wujjAyilaT0UxXtTY+prnxoz60ZzM49a9ORGw/wkJuOXnVvHG3XDB4Xl5BMxE1Xv
KSK9YQCHkIRT0F8rOps1WX/WCO5kTTbsPZo5igdj4QpXDCeJfNQ6wED8erXtxJcwYzuZobhgruYq
pf+F1tO6B9wY6oUStWE8ekCNt3YdFnwjoXZeBqjHYp0tkOgc9DDkrq9NkhSoCj8tHfRTt7Xi1OFf
5i293o08mSS6VWpZsOoUhiIXVT+OsDAhPNN46mzMP0L34R7HE9scYjd6eGQzviiJfBPPriJu33Yd
2zx7ANyJKzTCkkCbhu3fAHMxGLg2DBXPKELFQgPq+Nbyvgz19cfuUU1U0J1Q/4U06dIewqOwp+Qe
ConU3eRf/VhRkzSSFlBrFnHidiRU4AX0vZdPJgt5gB9rd28xifoHa9T6DFkA0bqgBswEQPuHmfYi
dtDVmDvrSjmQTdEeKjzE/rAVwEAW6/W2Ca8oJj3p6erdRcGUQ8l61eQJ5DsuQWEBZLv5A38AwTdp
jUM+LpKsMTjCWXAZpUU/c5SDCNDKElX/rDLbNspjQzJHmLjlp3xDFAmFjF/c0KpjC1C5SDIAb+lL
ZrPXX991xsgO8Z0mQQaSzjbB247qO85TmMcPYJV9g1gSDvr2pFJpcUVw6y986NCOwmBWLMnKAVQ3
Sv/+j+O/yr6FXjO4yBCBHdk9GAPYwuYO9fx+dV/y2OIvK1ZFhxO8zcj5hSBbrhIKRmbVuc33LUk9
EWkFdDivPUUDRY7rMe2yzlkMPlxpGBXFYzryRie5hsXflduyhxMwsWkGrFuARUH7d0iv+rsQPGi1
GaAp0rir2KoB4LbxEBks2BRWSx0kyfTV72kRJ6Vy8lGjNT9HrAmD20rKdLJb7l2ohDqyqS94poNR
HMk5r+t93xZvzFEtv2+iRnbs+Jd48ZjIhgP/T2s7K9j2g+ZzfCJ3wKlyQ/lRc3iMotoUIpC1kZn5
iwj9rscGSSMaasXRnO3jbYB2Vths2u2CF7uso07G4YXlszBmwvfQiJnS4RYk/a3GuDjLqeqAbsQU
O8u8Wr11s7DxsbYyH2nIvS3xVquNbCbjo2EpGqk05uP9fgGSE1xy3BcPKVc3MHfk24NztxGjZ6Jw
H6Biz0zYevSpzyISJgDPGP0BGKkyYf+nLAuFHl4r4Nr0WaxO42i1P/AYrHE54YQ/M6LtdiNs3z7f
KvayY+xRhw5bm1ZwSn45SXROHotDl3jE8bTuH3GIx68HaYV+BomRaUMacrsHjACjs+fLUYGz7ob1
Z7iWzTnCHTGqs4nH3C0TZBail1IUInvR9ZgND2y9qyzzj1sUdCcUte1g+/KjEU0qrco5c8oW/nvM
24U6OhGBMmlGK2p1OzF0x9NRne2D54VU/G0HlHOHWlK2Vb/slg+rQ3FB9Ani5Ez0t8Q4l2pgwWwT
6FqrTudI0M5XqLr31UfAz8FUJ1MV9laCEKd2tiJrrWNg76pwcQgF7kb6SjHam8clWeI36RWtS2wQ
wJ+7NZ5K6Qi36O2Ucz7bp3rLBgChC1wM2YAOoTgS20GzRLJbl9ZIX638sOmuRqrRUJgeA4QhX09k
UfAHYa22Z8LBFzz4aQZJfjV02ny0tOpdNFs5lZpBgH5ZY24CMZb+JGjQKtI1jM6W1vGNEBumA9Fe
A1xhRsTD3X0wCcG+Elbi3vN39ssD8sjRdelA3/it1F7A+v7W+hT4ShNCkDOI6L6KJu+GzAVaiioh
j7AGe38n4vkgxb4HVn/nw4LnCoHDxhQElff0bfODvCjVVp2vxEag17jOUX3fPy6DQ8+A6j3YVqRg
4IEfIaN/Q8QBAoIdEUuqBQtpR7QOqqm/eXJMDVWUvFWbDmXPJOwpplWVyLV+2PbGBG7ujZ1UetOV
eTFBKRhGNiN1dvMxGMpJ+eoKzNtiAJOeueOqKuScMOQqW4uia2HKgsmRwUW6O4qjaaD06JlkVJgZ
HamHTCyD5RDF574h8fqlQy5pCX6Be2Z3i0NEkGRjm7EMr1Oc1b7IQzx6mOjc90joLw9CeG1fJvWf
RRU1t35++jjpq1dujbd3Ykr+DLT2eF22+E87HZR2e2uz1KjsEFP0TKHuoU2tgjYkZo6LW4UrCeQp
yPEBCiKKxAvaoR0lqlQKqJ5A+CdnKS+1RfB25//de+JZy9JPWVDUnGXhCCEo7JW/WjSihlQtUcIB
ZpNzp7475ZW947xWMwvqwlBr+Su6S680eH73bFeWCADit/4dMF2B4gdrxPOvKdM18g6JPwiLQTmj
pe1dkagFzc41d9khoyxziZ1OsXnUH2p8+Ge+rMTBV7/gde77DGo/VVOYWe4+GZfJWxpc7PpLjSNT
RsOxepNb8GombWEye9zZBrUOpwS2YNDzq9h4rKNugB9pNw80YdD9KkzeT8ylwVSfL1Gvh7v//nLn
/ChZR96aceci/8a1X8GRQgWzYDwKpQ2HkD4XB3kD7sArp9gwK9YeacBOJeDHyRLZL/bx6b35vxMo
Rg2y0tB/YoYDhRHNnipzXuzs1AfNm+vxlmKU4YrEOxbCqx/5NgHki66ZyPTtZtOdHSM5f0solBMV
G2TCZmwmUaI/qStqPl/qzNBIcjdQOz0xqSsgaGHPG1Uc2iahZvKKt2ORtjp6FEUY8z1T06RN7yzl
1LT7ziXp+bdDjNkcXTgcOEkbh3dJZkuAVJiMx9R9fY1SV6KGD9frsyC1zQopl3nnPdBk7PLWKnKG
jOnFcdWD7vM8fKkIXsVelFZPaA4ZVLunCmoWVoOvDUPoX259XMDwkXApamVsQmuO+dReOlH9AVJt
wx0STOGkNVm9mJQvq/WDRyFfWChyAVV1/H1/IEraQF4cl9YS9WN2X0jCZ3sXj0VzwBtgppb++GW6
9bUo7zHjGj7X24DdCNpokl+jSB9AN8jH7kIjQzcXs9uCMrCUkhgPnDAqd5ipswuyagXZGBIS/E81
b/kxKW3aLBD8bzDtTheeG8DzIcI9zW9b/2Awf/mGH8b2RN+6IYIBnKgm59Ou5gpLXWXKq4/CtjO7
FFpKwiDndOfAN7O4Jw5N1ps4UiNJunHa/DYfj1JszxbZ8vgS8vpAuK+PmyWi5KmdnYFpKpcgnobp
XOpxOYVerUFo/E8A0llzOxsd9OUmAeZRSeSP0vb9nA0MBfN4FLgWG0DrhEH/Rw3fVKdXxzdm9bQ1
HNquuP/M661paGyzgEzvX4stHvrK9ehB2zEnBNbywA/swV8+TsL2nOAEuKFHifqsTXHu6zNoKgEW
yD6aJQH2+jlwDLmsUEQbjL864wsyNI7wVyp9LJupGN+rSmyQjJm9qv5JdcPgO/zDFLwgSu+/Wdqn
+vVU3RbdsDceEu35TKfnupk9kv1iexxfWXimmu+aAP6csk+QMtDxvhOWpkR5UmJldddezc3gVI5b
nIjX0TnKAqyHevfr+c9XPEjsDa95RgA9XDkFxZO0NR6m1kGBAzZ2qCAg+YJ84p6YB4rArzhWWYwD
eHNzIKyqcRBbsCLEQL/FBA4iQqrcfRsTjdiCsyHiHmiQa5IyOScmG+BN6cB04YGRksbm2SgdCgcT
Ll494uhJi+qwXdvnZ1ZIpRw1omeh5TZIn6JkjQJnz/UgU9BSfTzjG3SOIArpvniwrzDDsRHZKfOa
WrHsn5d2lM8Tv/YouwAH6NTLpD2hHlGtyyHbUBMbNOV4RlZjWukecFdsSuBpsvvnShcfvZtkUqLW
U2T997K5VTaQSG8zGfMdMKGQ13BAUATtI/HD8z6IEWqb91d4+gdFcN5oHiH7qqts9OaGlqDoVupD
xQLNYgxftYTZ7/gHvr2rXb7Gg9kND64Gxt4z16WjTEQitS28EDR+sd5wvy3PcacR+iNqXdfPOeKr
i2CMbJqXytkCyQR5HC3LXNZfFJ/Ope/Oa9waIu9rAXsuvJ5dLlbnlzePHDxqPzc6ca0mIAcrKFi8
pwlzG++yGteaqb36N+k8mfoegzevCS5F0XJ6u7p5PPMAp6r790UhYY5hSOkBQK09qOUpZH7hnkWy
5oszUL0obuLahu7IiLDGr/OKTaEDYJ1Lz6wP2/RZVPfXi69+l9O4rmOFS1CuU0PxuAv9LQuHfs3R
RD8L6Ch5Z5RjL19bdjQMcE6BkTmpEtDUHD/XRYBi9/vdCNQWPODEcJEvK8NzEWqPdfHhiMNJvTGN
B+agVozpyReO+iDpqZbaULfFC+Jg8eeplDg9VPUzHDwGLUu8CaWBLFPI4rJqkpyW88+FkHVVLxDn
+4TZOmVUzU2po4wSTtnn/CCdk2G6zeWZQmNdMIruXsyUfLo4jHgoyCCOyff9ot4aKbwYjUGAqXl5
aPXRbCqyhTuIq0u1Z3ZWD+fM/1rTcgN1JkEPlpYk9LiiUO43UmtEn0ckTKlAdKl+0sdu205/e8bp
FKC1SuOB+6X+X+GCR+oHTAQREv70fmWA02Ks3d7DyHylLqlf+CiMwNzLJ3ePMT56Wpk5w6qjLD60
1647i7uUsp5gs66ueo5/FmBSKyMJwty8kvL0jrdypA2JvEbYmi+3mPw9uaT2+VyG7uTT1zjurSUt
f3k768XLjS+4qI77P8d4S2SK7NraA6uTlfjoip+ZltlI7Jp/DXYyR5dSRtz/uSjVJOg16ZDtif4z
6ugo3QV48SJJ6zX8ixqRepVEbNqno3arM0YPvYxsMaljmzq1Eq/kZ9i2Jo6jGcgXloQKyo4M1A3s
kfCYni8yTTqXkGy0rjcZ2bn4ecNzML/VrM87SwgB5f6KECeiq60EU7hblycrJMtJaJ2TNwFE5bi5
/cGu3Etiea4vx+RC/srGg8TDSqdtPDHOfJ+564U52D82iLpbD2f/2jK2eOIR9kbR106oP5Jxc3K/
nekuUa5SzMmhOCEzx+mWQ5EbIxC2wryS5BG22swfAJNQw8R2mWFBsUBk8MtPZdKdcuDyFvz0EaBA
P7oqz6yWwUabiHxBvtJBmNvf8lO8b+M8mDh3NyZepHhqrHRhdi0SKXeKVIaJjQIaWjacBhgjRAin
Q4KJoMhMvdmhCtbUYbjmX+nVt7KacpA5t3Go0wnGEOT2eoCSeHBHjQdB0k0CuCJkQzjG56RtZjeC
DE6wYoT+Ti7OtsrK9tg1DLfJPLTyvHFAUQUADMb3PsmznxAPVL9QYineId4Hn/7PTARSJbu+paQE
UFCkH7SmXogygPwZJffLYwmhWAMkwjCc+pXyf7qI+H6JtavjwKBAzLWC+f5I4pId3GeVYLdcJbNu
Bs9ebQbBlvzfQuhfpX4APkqNx1n2jAi+fEuL+30jqIF64dxaDO4huFnDa5weBR1h13sjMXYPJkN0
MOjIuAmPD9opufp8cx/wNb77th7uw5L6UXCVC7ch4QZilkuIkm8AeLgw9k9fd6TzEAWfm6j4o+R7
ojUPE+FoqjRC+riLL+inEpMdQgul6mlRUnmsvp/829dixKPL69U9X2ZzIzL3QglRtVEWZS0RXsCE
7bYw3jtk6RmF2A5qOcSk0Hk5wDYApjV6PMu7Wdp05/YLwbnXnmRhCn07wmVOOX3Ye6odh5U62vGI
MDdyMIaIEE6yRmJiD3EZYDxTbSGG6lqRFa9vFwWFZz7y2CGJ9fB0P6YTj8UCBmLa5BnavQh2lEsi
Adw3UKDkgubVxUfMerLGt4zsbeCWpUWwRtSSFSoAdtCrnqrDqZqgn2cS0QzpQdQWtwD1UJbs7Q9j
GD2ocxGzMz6PDigkQFaC0SNzLm886+nY4lDPOAvsWvvX4/zkI3B2VwMKEuy5NMzNOixew0ne4nPM
6ORsgnMKiD8tFO7ztKGHcW+BAlgrwO5qhDkdr8iHyB2LMOZz3ugBy+rQNyocZnLGxqdBjtzdB2uw
o7J6ZC7ZrsILYp5yYQvPlLGpbVdzFhJz+5eeZxv/f3+ryfUZ0fHLTzHsW8TmKhOdEPn+qzPgS6tI
RnqAvCXwGie2O+erI2F6/NrtfBLmii61nKv6D4ce7oatZCDWdL+koIMvn1tFUfl6h11rPiueVN6m
JpJhmwYdCbV/FVM/W2YwF0qA9I6BeC9YS1AfpN5t8qBh/6wI9GW2jwSI+kn2SFMJ+LKII3dckYTI
xjoI9wbOU51E2Xg8dkj1BGNC1q1UEgZkg7LsxEW+a4HIutJajD8ocXwBrlAprOVazZEPwFpauQ1S
rKXAHQToWKff3ijoOGIqO/NxpOW/4jyqEJiD0Au2AR1FSss3PnYhm3fTFEZV1toO0ZYbR1qku/kn
BAiij8krs8Op+JhHReTsRoftzyEH/CWo6v3b4CRSyr5LV0msUgpCFk7/S6jbqpXsrhgyirS5D33w
A5yjgYHttMryfZwTNxyvol9quOYa+CmJgKCkhaImZzHUI8VQ7dLt0I9DNGslPR5ZnM9YYPRWq0mf
AjEhhx7ckSp1/KTqcGeVazjU2+e+7OUzgXOJza9oXklg5liZAXwAknffxJzW9k6CGa8YWZRV1cgs
xlAXD231tuxLOq47OC4e+nJ53PI4CX6Kj/d2XgK8vY++LYDNHLtrOHsGelY+A78VAYtRFQ1/KE4c
Ou1j20DClvaME2hNtVQ5iuM0J40++3TMotW1h6by5RT/vlSLpADvaQNxpJJTC8YlnqVF+vSLIS86
SiRJ6i6/fPv4f+D4o8fZQATqz7ov67MY/Ti2LlApoKiM92R6Ow5PnbGvq7qmybRJMvUR3c06sVHV
xgEf4clCymqh1UFydVtK7Kb1Ul4EfOiV/e33QydBlfn1qtTL1l0glciMr90bOI4l4YpbCbhkgJiN
8V/miXDOCR9cybRoLnhBFy53iIn1nVjXoTA0HVa0M+1l0nC6W6GzDJ33PhD/gTvZiJJWuGhqEhXB
2OF2CHHZYpk2lot79ZCPlhV1M4xEVpGefFJdlcF1IThUdAObtkhgcYUipVulMS2H4KzCkdERrNcw
cfkNpZpw1gFFUEOzU8JSCRg2AT9x7pI0gKHYwcG0ePj6h+fOJY5ySm5joAmPXN7vidcyWqMtsVnu
LvHTRokJPP/j00PsiwODtz5NXY8MowPzGEMuWLAtkOkli10t+Pjm20Dbth3aY3GUwMr5z1+HC7YK
IvwGQOYI1j4JR1yfQOOcu6WJ7y8/+Wi9XWZG8U2N3LuUyccLfWtgYKEew/P/zCzaCtmcrOK7ipOR
tpbyUH1sKuaiWc3oCMNZ29UkZKfnYYijYsANff9F5WFPwq70VfBRV13B+Qp9Kbb49m7VJjQXWJBN
xmry3A/Mddksj2561jQplu1lhnMOnyN0E7XqLKz5c8xWH27NUw/nKqPiqGlFuf7eGOm5phUkOc7g
QX6u/9iHhwgtH5/Q9qKqHfa42r4m4WuztpEiBfKcdvWdyfFO5JbvVC4xe7+yZ+SAyLsBZBbz4QcG
mM39uc1EpuCTv/uGdKRNrUxFgVXteFELmx4QYOBvMh06uLsmorSnMjOv6VDprEv6V9KujIxTjIEa
Fg7KI3bOV6SIQoPk0NKyvp0FbnvfWMNpIRkYCXeu2FdhJ/oHrk2ODlxi13OWXedWj+MQSI8qvPBB
zoOVtGOxc4Ueibk/ltM9A6brHdZlY7wqcYx3cTolUNYoMsEjSNF4lpYagzo5hEgw07P/P1c8tRe+
QNycmi/ZwfeNDZ2D+UFV/sE+y6DW4mOAmAyBv1MErPZxdhVrbTbKqqnHNnlTsVd8RIyDbLb+iCVh
5iL6DuKLzgC1tAbwLc/Er/M4ZXYry6/FtrkLfdDhP31fy9EgUM5ywFPu+OD928xp4BG6lzAeC6Mb
nC9Fnx0XIvd/N0cpb9SIpk+FPmdpYYoTEvDy6lggQleNXiOVQHojCDOw3iqcWsStPEaVLjrnDgwc
tGJEjjREOh9fv5Pjtx8q4iwIHzhSbAP7/Zo46OrU4OsR7lc8ITys9SL9Sj8VEHd0UeXNFXRVqBcH
bC6e2vvdJR455KAY5MwXYELVdCUq4qS73xHI8Top6sJKYghpbqtaGQ+NblHynotya1zZ8CMMxRbB
H2QkG4q95N53pLyG4ApvYxw8XDgkMtLVUNq3Ho/bnSo0OofK4VUASDR3xkmgOj2DfmR6Zwcm4k12
loAqs517127MJ/6Tdfim2yQJQduSqBaydEKgyrkPRxXJ5q9A5cUmF4ln24MIwyCE5gsMdjWVzaeQ
MSdVLMWkyFmcxUrn7M1qMLd4pRTv2qcco1loMCnwHpqDjnPf+l42vAEJY1E9PiZFnfkGdqimUHmC
PRnnD/MJ/+/jKEayXNit50MGp0nIYcf/APn1BJuWa0uRpIe7lTHAqgnb95o7PVA4yJglb/TMVOLW
i/QrG79vHxfqIc/OZePEx4mDeMHqe61PsMLeFlampPDFHe//JvgBXMkiOkqzss//5vVfgGNGAv9m
YURfyqzsRS1Yfjo4YWxgrsdc9cxpv2mPu9Rbqz5Ia9PODU8Nnl90+jflyvdM3ZZAYZwFytEY/EGK
5wfxAp6p4I+SCtL+PkQ/2caakvOjuf+dZVBo32D8bOb1fl8KqtZrNve7dggaTXIiW7msxq0mbHY+
Snj/XxGtTbs8AXHCt5nfDJQNyZONk6YGuOMdM8HMlwLbmPJvimyFou+XsiFtOLJj0F44fwJ8J3+W
PDCa34uRmMrb2rGayFX+l33eQtUghsEGWj+zRU9yQC0ot8MroBrwgTiBDvA+2k5qkKaRpYz+WUCG
d2p4rPIo1PJIgLgceXG6kgFyI3q5iwqiTYKZEgrlnLo+eVbmcZ30ZJ1EgVBzup7x4AWBWtBaP79v
nUPYuv4UhAZYi5ZmoaWu6MkoEGmnJIAZUeVV9IW4MVZYLL7Qh6BpHiuD3DuVTzOZYc/5Tkj5eTYK
/q8nRpQ9UgkMd/Iza6rfm+317CNyybKayeg8ECKmkJ23bsWv++UrnCKahVVzRRKXSZnRiD3/unzI
sn0JkKct5GlMtl4c5EOgevUm/qOzUHrv0OlBwtakUpdP3GuWyFxOxu09r7tyL6D0whc88em6e0f5
kz1fESd/zE11I/1Q203c+D5g0n0RsFJX+fIG1rDETD9bgfybmJj+SN64kspx/Z2dujMCLszkb9Nj
/DhMPnblG8Gj6pNtWyGqhQcVGKFoapWNvJSB7rzDMglAqfDdpP8fHDwqf7Vv2Y9V2nR+cHf4TZIF
4PVMaHM6g0UPxRyc8M7slFvu2JtcqXYeWxYYOXAK7pRt87vTjnizkqaYL19XI06OPafht+BpZvU4
GWhyI30e+BIvNwQhCp/X6imIJWYV+9Ep+cLap31Yqa5KFVRBM/PwjF1YuyzN1jxlG8pOc7RB5JH3
8Ciqq1FVixc1OXxwaif05prYfyBcUMvqNqsiRLxjHswN51vbbXVHzZ6/DJOvVOoe77rQMRnK+7Wx
UkBvKVAypAMHsuWoxXwPILYknyi5wO8+GtqkSIUXXlZAdkujpe5rgAHSX4YHwjI93xrS0+XSclMU
8edZnlGDhbl8LNWRfgPc+XhFqer6Zc092jn/hgNkwMg8n2M9r4WNDFwp3WuRB8MqZT+EEUo4KCfH
asY3sdDlCFWXIufxyWvkWPji3XVLH2ptAVYM8VETsJCtm3WzZDEl3YBCeK0fTwjbVHP6mCUSvHKY
3Q1+ZLLMohGJL7hWYFoGhg4dP0Fkz24Iqj2SPvzpahk3XYOMl6Ubc9V8CtElB3V/Wz02b/AXlPVc
f3zSxk0m0EdGXMcsvcFVyp3o15juGaBsXwRLiWUMdpJZfvmAWHEDH1CJpBAjMZZnqnF29iFB5zp8
XNLgs5YgEjJ5WC66MOhjlKhuSifi8VaTLKTIVFL1/LOr1UUAfq5E/y9SSqbMa7d2vTmLSSFYlH06
dF8lAl8wfU0NczX0UeHkmf31gqkV8Qpe0gmgNT4Vj4HtQQ+WS3RudX01EwMALn8fdcPr2TXoqlxy
IfQFJcguixxFPkSQmEj5Lobe1rkIacWyBhDtGtYaTAB8d67mcODGiUkb3nx/ERSvOM92O6RjsybC
n2GQV9CJFzoY6KJ6YcJLQkX+vl4dC6c+21Hc8YjsFcU/uy+e1DFWk+k7cTl2u3mzZEcMFjREY+Lk
5XINtFx2QGJ9XFIaf3snU/Z7EsnauZbEN1JYzXJ6VeSZwofodV0ylLC6yA/grL5fDZas0a7bdloW
IB8vCt1kHAJIFpfVtHQ9qDFADKNntIvuQX1fKFM02nGj13k9gIo0Dq3WwpH33zpS2Hsha9VFjohM
41tht6EJ3vyOVnHjbtk8/fDVTJbboswZukA2IR7uJStlzOVQ/6kRSsONK5hnafTZ7yxzy+I/UqoB
vodSxVMAs2gCoI1WdqJrWDdHbCTLTku4nOQXZ6jufGnri4plHx8yVT0VlzrZtPLff1cUKIhbwYUP
IXDNsCoJzpXoCuNMO8J+L8FzcQV/Ld/+E06v1iKHsX83tStIh8mvqwVJnXxrOVysF1HJFDfBjNIt
JSMjK4q2eSFO0t7M383flnY5WaZMHRwrFmpdyY9jn7RbxNB1NaRzWle369Ley3XVQ30pGEpFUqOb
hjeph2fayQmY86GdCQ3fitO1ovZdbSFeWHC8hf7JqgaD0O40/UgxpDStK+P06Ek47Hq7uCJoPKvm
Hs+q59yZsQrYmQt8bgMKvSVoiUtMsLqtfyPyykUf7z4Y/LuP6E6k0dwYvp7FQ8PxUEGdPNjhLSaM
qqkBEh5N0iAhjY91rIjsPtclYEjZ+V+Jb/TM5BuihrtMN6eMFOD2gZF0kQPNCClGJIp8iWk2asDf
w5MEKqRxYUfwfTyjdrF+/vzX6H3u2p02ifRY4GJ1bJecNJ+wcSl7xNfKwvHmAr/Q0vKd6yOouJuf
fxpKcBpNF/fBozs2e3Ht+y2ItUZznO3RGBgQcdSBeZKHnlFDuVF9YTFz8p+ulCDIPUm+8aBlbpMw
qDh5gi+zgU6BNV+EOSXJ1VZPk97B/D7Wl4crsf32EQEPBWi/P6+4845W6eguN8YRJkP6puGDIAzZ
N8FJl0pNJ37tjC0tzK53YiWXvnsRAaoVj/tOAM1/+PR2AsxtjXwpNwjBO3unL/SPkfUdXaYLDQVK
Q3DBiP36fiTqZ7ziuhXEXOc5Ri75pMQ94DvNwDyoMZvDjMq5yeBpsChK9vsZIkHvAXAcX1i9aRhu
BioD06IVNYhhbPMf/fZlMA0Fblj+f5ZNut++ee5NEUtYqWNPjj0+nNPuV68AGQAXdRgJr0uMg3gm
d8jcWe56jea/Z8LPgjVvnH/1ZvoI//0u1hs3SEaLNd0/bTUbH91nmS4TdJr90IgeDO0RJrD3AfsD
P00AkDQCh0yUtcZ25wYrU8oVK2xqWlk/gn26RxjfmE3/HWpeAlLIXim5YUKkHlTfkSPU3OHWb7/r
O1LoUYsk4++0aLYD67tyQVsxj65j1iVV6+JlcKn7IT6HmqcUkLvi0+dHNX5yze+SZHNF/HuUCX+h
NdW8duRAvLpqleCBZ0WqnSLY0VnTtVJnLnNjyqF9THerJ8Yq4ut8QPTNiIFwfdIUKb+skC4FX1a1
aiH6jPYEigYb5N5ju6VuM8xiTVH0jkvoD+yATcJZvKt7vkDfiYKGgB7N/eQd7L3SkWI59WzQwRqA
GjxSqxrLVU4H7k8R752cVWBLpCGVtxvBxiDW/OEtx9mEIOHE0a2qk+WcMTkPsHK1eBPy8ND66cTS
DdKRw94lCSWSRnPm76wB/bUGIqLWyELmFtz/ygG7qWmbIWsoiLcaSNrY4BGVHa/Lg2wwghL8WV8M
a8vH/ibxafPu0Yjf8BM2DxBSmmBardPve6/xhra9jFyozE0Rnf4114xnh5QpPcLXsoVl/C0+QY07
J7vGwXZipXVbIYtTh4lGqrr1so7Wj9JhcnSVAhZlhI2wO8Z1Ft38nFR4rb6TNfiMwz199hwLr+At
Cr8JtOIu2QwMR0oR9nW9zp12me2adt5zKy63RcdgIiSRplnR6XkmbdyVBr0c1samEAqtb7/qU4cN
8vUZWfYKqA1QnE0Dnn5ZLtcdIMbXnfypeL9C4CAh77LK3Z5YMUrHIfEAzqnLbKH2ybvNI+bl5C8A
s0tuZw1IM+Xp3eVYEzz3z2ysMNRJHfYWqgNAn9RWVOrs9HvZ3QRg5IO46UAQKzQP902uFLfsCwl8
jj2u5d94m3OzQAsoD013GJKeLN3prUOWTrno7N7xQxaMNnMWFUrab73z7W1V97WU0ATwQaA8H2hn
2JQEvg/PfXdgT5hdRlYcDeiE5xd2b71EOkdnDOUuDSoUHCz1jTMBJDMRWdXkEJ2QSD2TWWmPz1cQ
PHwihPJy/89dSrSJEGkGTWntmgRPkOhNFsKFUkjsGSHxICKvIypTvktvdyW2FcanHFXlp6A5CqsA
9JnfOq9hGSibXURMw5xNzZ0uLRV3QmrDCyxoCylVeOxI5DEqbu5BtkX65lmGCjT5k0YbtDVZgM0W
xRGe07CR9lSEbdesJngtbtl38Yo++nqCBXOc3mVKgWrJkOALZeOApRvAFXKZVqKjdISpYEo+ql3g
WIJFNNJiFcICTTASa5t8T/YxkmYHlc96SgQmDTZyThRyPsMKn8JrNbmnh0UZC5I+zOSmHnTs4n/9
ErPvPnZDdIspI+CBtyOjxcO15rfA4v3w9HFCcBXaEzrGu0aBeRJiZLS928oGAh5TeUPuPmn9gpCV
hsbLlSOZTSPi0iHAqxdAAOr9BIjEp15d3/kXMEvlhuY5Ju1j3eRl6Hl7+8bQCYiu4fd6OyoSjGE3
hyx8ic29dUlHd4xmk3laNN+Co/oEDRakmZ8TeSvUlqDOhVep+sdq2TvvXURb44/Vwo1e/UHAwEws
meUj3prhKmplCvtRClPjFRU3tTsrYKLkOHD2xC5ciZ/5XrIv4osswxEahwaJ9ExfW7LegTaGyz50
MhDdj1KhoDhjdUDADNkdbHGJ2ave/QIoNHrR6AUjE3s0w2Ve+e1i1QIUtYgm9C4FufbmPxzIZnyN
pAVvukdroSA1VzGRkl7r9MssbId81VbZ2IkcIWA+wamDvs2CnBKxzoVgfEufCi8dofYGlhL5FNwe
vxGcIGgzXX2HwqiG/PCDJIDsIpnih33FpAIjiI7goF8GZ4nMZMDi9tlkYzN3lOD2us8PR5oP6mOA
y/PXqzfyz12dcq8RPQe+Do5cHKqY59CzvJ3p6hUh37f0Lg8XjgTc6txW4EtMwQX1HFaPntWu/69b
wltRBhu6+tZPfYTblbAjy1lxqiOks9KoGWEOIVeCM5GPs/rtVjM7Im74VlBpGbwrvscmYz9IiOqg
B1RTtXr3K3BYr9OkKnmmZ9liS5+XSGFFb7mrl23t42lkAd9UbeMURcjQcxNqwjBRJJvn6OnLMNlu
1oqPbgRJo9oATjLlxG4UZhkGi30fQwbaSmtrheRVytDbzYq0eb1oOJxgV7fQ/reDt8CRx15eMmQF
h0h8FpexJZL2XiE0ASDj3DHz8vC3weRHgH1Y5p8JJLqsiCaE48tvU4JwYNr29wlhEg8eP5QF4beu
Yrpj4l6nSzLt7B7Bb7/d6LmuHg/bnE//IZUZ/iu58PO9RrAnwfOQ0gFjRjUAuTdPnChu1kgiKayT
sTvYXf2hL0Zh9y6ohL9iKq/R0qrh1+iioUA4qmNaGGMFtK3hJ7SyLSwcufx0eAMLNPmNy9v6dTNZ
1v6Vz6ZgX8ULlgCVGFGmTeMW9F8LrH43H1EYNVBu4lc+/Xsw862z7CQV4cQWw9xB+XupTE8eP9WB
fCIcU4zAnjxfl4FncEuAFEF65zGPiMTnO59XeRGlWMOaCE4yhOJ06NyLz8H32FArBi0uZAXQV9iX
s3CaVGxtsqafUv7Wkw1eSYz5aIBQO0WbCM9tK/jixr4b4WOZxTiFhZE5Sc8eilKyZU/BdWsY2kmj
wsA5j/uzQ3cgVNI7tEjAFCr066qU9tFgsGoOWs+Psh9Nq7nr5c8XtNkdhaGPRNYe1RTJr+vX8q/N
b2kWsDgNV4PiOQBj1+1QUocC9VX6Q0ZjFMlcjTC5C63QwuKmWgZV3xIdbcLXFoqcb6H23+J/tulx
PCJE6zCaScFdBWxQZ/F/dFilR8pOgsLA3exjWFDSvzLNZTmwj9rgq7MI2ov7+KkaL0jsSlF7TaEg
Aft4GBgp30XL4L+clwAuuz/O2KssoxzOk8j+z91D+SF6t2HL8ep7SZTq9ldwf6AGestbB9hXY0YG
yqVy8V4ofzipHVVxxRjOgMespUdqmRtieYreVCxYsRQ5v6AdIf5LtCQATLbvhGg6YYnxfF5p0foQ
xIb/rjGoJtW1R67D03ZxeKKarR2akIuq5Hbh8RNHkoLUsYi6hW66OGfDj47LBj2MlvC9BbU3bo7y
byJT+NjoF5hamRoTQ7NU1vo0GNcdVgEVX27FK9GnuKaWhGo78xxYhPL1kMTTFEsxxROVCMfWYcq7
dgRfKcVZx6Hi3hf+W2aFlSxT1XMAiG1IjAJ0nR0IEHBgAJbbMRw45VD5vWvysKgqeQw53zWBbDz8
yKLkoNWno7LaTcdPfA5BksyIVAN9cb3OLv9TwPkn8Au6IyYpI1z54NsCJN6Pxi3T7mzu2XP4KO4K
APrtAZoM6zfkC++b1LughnJR9GkhvptPPNkqFsnh6pJ2Dtd6xY2DIVaWirm+mSKbppQSXtWiTZpo
tun8CtYXpy9JU2lIWMn4UDLC58SFNIQ24y8BarjP+AmjPLv//suM4hZa8Em20IC1ft4MfMnv9P7Y
2kjv4qv3RpOSJm+Hlc+R0F13/pE84IIslRyru74M7ikdFK32uDyUWxPzUxeNiASxh8McHwbOLpex
jL5IiqbLXEDCK4gpZWPTMvOOV+Ejt+hmQGVMqhDKpPFv313+UfOvM+4caWxS/PYKHM80DlOKnX6Z
d+rT+vjwKr02whetgU8ARiBfsZPVXXAEoNwaIsJzoKQ1JyMC0PtZKaIFIVFIuovbwrua1Zj28WSD
+gdTUu2B5jSQqBAPkNowd/d0nx+xPciL/ABGMLzIZllk086Kj0qpwxdzIHoSYg0RmzrEb+FBICCA
OQsCHYAqivC0gJli/rt3ncqN06PXS9nZZ8qINukn5eM/Sezd9/OSK5xq4h9d9fXAbLb9Qw02hzW6
VCPJASUYyRNsSbP3HsCTd9Amzy/BQAir+ybsc2Y5eGxcoLWr+FM3YiqlxOE4ICwifQZfWBJKRK7P
qHWZUi1ggqZVVCnArZaJnaXaUQblO0jlLc05ocUaMpqoAJZBH/bJt6HT6RSVxwo2IsQYVlvre8ue
jgHthRet4o1vy4zQIvnA7Fogz0w6nHLUhJPQCqR3AVEjQcN/sYsE2BYOf3tCs7J0aO1WctjWrQ2u
IJdN9peu4DgyhANKa3DyqLBfUeGhL1WeTm5zS+VUMfrK+BWi1BUZVCJBpy/I2rPcG8roXFnUvImR
jZRFveNatZIl+t+do0kgMFTLuH6/vdbEcZRAVZJOcTq7YAKi0ecbc/f8CCu7aYElAx+e36ejRbSC
eICZceOYSE1zjNpsiuQsubpSoFoB3X4yfG20H9ZzVL2zaf6FR3uEe0lMM9blpS2tsNNfGfb8I5fA
+THkJ4VSNI8RQ9EFF+2R35VS4iASTYuJqRPMkpTFvsQblS0yDGxtJ0z1gOOWQN5yXdSut4Xx+Vm0
qyrCFYkYZS+8x99z9EVzKFus7TF0dZ5oQn8SGU1VXqFTFEXtcBnsU9tI7KOngFIJ38TddLAa6diW
6JEV48CpPD9yu4Lkj+ZBwg6fwnpM5VFlVEz71ia6UnE3aSmzDHV771MvNHzo1aW+GXTUunuS/iTY
X0r9k/G/vPjQxOfKZRp62uZq8sNKqamnqrAvUwmR+Nzo5oGgJkx8QLTrFkeHXPPcTwyM9504CtXT
KjaMiL6tnIl7Wp0tnN7EUsVY9HLJe5mnQvz9PcMNEd7wGJ8xveidJT8EltOH81nWAxss3BankNR6
kJ24X83HRpKliMof+S9JD//If/wt4XtHPL8lo1ucWsEKK0LtPc2OXv+wnEPapepj5EYCh3tDYDPY
4Rv8aM1443sByd5EJSAwRZ3Ibe2f99t1qwD67Rbf5cM1xes0QY0khEH3s3OWCHayiXXYXIK2az6T
mcGSG2L7p7+E2haDdOR5XccDffVE3VcVTFaGvJ8ktIq5EjUdSfgZOu0S2Qv0M7EEzcWI0ijoyIhV
15fV9Yjg+bKinQ8+k8LfZoq0UNV3jqT3Jfg2Qg2NR0CVyFmiz3WQEvhHelPjg9fw88ril+AOxokB
kUTk0ToXkeqVy2Gs+l8Hz5VX+371JPHgg9270Mr+AfjWaLUuVk6VZ8NP+Ie5qXYRIUhBLaba7x28
TXY192UaFrmupUUTkJgmLWzDy9c8o5VzbL4Hr0a1E8JxCqeeToQuk94vyoIpFNE7Ah44IxxLRniW
5dENi5mZOk0BekbiMSizLW3EFQVwPa8MnKMRd94o4a8rgNEfhO0YMNOERiKHwdD1YtnnZfQdlqyQ
7/q9+0tXievgY4Xsohqqlub/C4xVCPSeL/aMgNxdi8GiKDTHFCaU5i95cZrLzeb7UHl/1rGzLoUY
xgf2QefyFDAZg2ek5o5ouW+CYTyJkNz/4p02pBdZJnhXZU/8aGSsr3KQ6xeG0XZ1RN0ynN56D0LP
L/NafV7i1bGsoRrVAwjSmb7HVJr/NlMJ6KvdTSPq/UBSHXT7Ot+wvTzjbrW7+j/B9mUNUWItsVbJ
ZY17TkUJ725cF95wTNYPSDRw3gCniiWINV3sCk4yFR4+c49hGh5Nsc3jxhimS9cQBpvQ7MJh8Y6u
R9ArKpFlPsmoObSWKAlHhTEWlsDjN1CgMb9GThoCZ0iUcOOS87677e14vIwr/138wm8zG+cHjOXt
5/ifklNBOM8kpueIfKNZmWOf63/AGjdNpcLIUJR1dRgj1XtxAovT9ea+IxQAvp1MCNwSi2jG97Ap
U2KzKJuCRNp5cT7nSW8stEFuq2H6mtNCMBlRDPgHYarP9UEx+WAqK+E+460rghU4PrXdZk45apNX
fRfE6dNJfKtp+ygOhd4BUxn94egc3l2NNmsAEcYklU0ZFILqTdzcskRKmas4S0OV8rBq4JXDLW1E
J11h64PMZIPrsLudMoWeMRLFMIKozr7fO3fnNZkIkfEy1egrcM100z9D42ROfL+z4AQg/1NYY2VH
SmXah8pzHJ6bsYuLtxXX7heLfmXkUN3/6lRHMzxqcp42etMtqMSi9C8t31ZOy6KGNS2YTg41REia
hXBHSGB/cop9Ynj/KIIFLflLBvTemG6i+NqQ8A/quP8OOzEPucvwXVn/q8z9dKtCd9wJJvQQxcHD
zw5D4HSU7vcpRwMxGp2M+qWyVpDlbWrpEYk+NbqD4xfYAYResmDYf1K5VHej/8C+eD0kweCkvDpt
TueucFiAijkOKaZh+3ey06vV7zjqAeNY8xngqUWLnFqscL2IgTkmCwRoEboAS+b09wywQIyZJmpv
UsyxE9ZR3+ZjsBVAniBo8NAa9pMkyT8WyhzBfXVIZnbxcxVwYuaTolVm4NiTDnIVxt5YvRrMR1AW
zWmxW/cd9T/OHTAUCba+MqjjY0dQMxGFB7k3KFK2yYBLcQRpS0yOvy4UtzmzvLza6+GH8AljUOAM
FBREJ6mwlXHtfAYiSkUJ9by9oO7hJs1Ll5Z8RAyUzwdJFVtI+uAKo7UUY5lr0yYPsf9COZRMyb/q
SOvuyh1ur8pZHRgYBZw+LnizGj7RauBOaQaoEPVgZIajcWSanaIyhwU841zEt7almmpUzUJsLr6a
6XKwc9N0UoiqYc0+XBKC5/Vv2jZJ8KKMkm6MPYD/ibGZHpDUBVVJ/8BTDSSbD+NuFkgVYn2jsfxB
rI77FA5+MzJofEI+vATbg9P0m/gKMAdVvHzN6NlbBpgLzWm+BRk11JPI7v5jn6v+hJ7tRGEoKDwf
Im8KB4I9hlUZ5iRz5eps3xyjznnbh+fd8jA251mwl57yKa1ZHPUwdLqMm2spglWGbfT2njj7PHoE
typvs/fQu2YWwmBo96B0EBLbeo+m77XSgerq96kVLmEsl11wQjIJDdsCPOpMCHAPbIXhmiaxEHAo
LHJZlkwoxFTfTwdOl45gw9oNrsY2o03YMx2TBZmMKfEVYpBkvG4SLhgEC7Wz11rLfeGtSWyl8rPb
bWVNtaN9sDF1GdpSiswAQLUnT6YppQo/eqqZAnztDLP3pFzr9IFQmpFWg9FLHwYql4jWbV/Fzy+T
cZW8U2PQuZpT/UNT303SeFmCHbaUKt6cNslrBkOb9Q7oMtbK509GnMNbP3tg3UGXw5Yfae6ClAqj
lvSEHuN7wVC6dxmp5ec54qsJBr6slQ9fenRHF4YST6dPV0dpN0I0E7wKCQO1F04Ljjs0baIMg1AT
6M3dP3kRPJlX8CsNn0Ym52ZaBZ1akGpYZ9S4NQU1Ql8MFNMoJE0lFePMKjMXUoeiUMCoIiyZWkUt
ZuXLULKn2EDsZuhquZHVKXcfGnRIG2VWiiXPDEz3gfKod5jdQBrxNTfcgGE1Ydh+rNJxjAPB4Als
jh2vl799ZKan91ddkVoB0q9ZFl7frmK0vlkj3eKXGeju6I6D4eJ+bpP4Mz4y77Cze3w7Z3/Xd30j
Yn2CjliAa1c6kB+vFFZNubjcSkbkzrizQAP0Knp6uUJaojX5sjZpruIEXQwZy/3hKWq3sQQM9Kgk
LUwxzYJ2qc9EWJ6ib39Zcesa50F8Ri/8C4l6ZuHXx8wMxf9rMGc6ffq9N7JobDjdUybNgwDfczRO
GVRDfDx/Rk3H9O0yYfg6Y+ihGFvDdA2b9WWVBMWTHA1iRCX0n6Hgt9pnorZh12wPmGFptiulRdlZ
JzOl1Ud7W5gfnlRrgopGC5QTRiHNbD2QGYCGgKaULT7oXrerDRgCyZ3tEkKTHbaHk8GoL8JhvVSg
DqYq4ILINBPKyOwZdDqRkkEmWuKeFt+A012wQZoXB/zVOVUb20Axcog9+WgnaY38Ceodl/IFQMoh
OS2h1V7TFOKuQgAVLPpMuFw/xyxHFcFWEYYv43mNcM1AZ5kVMRczf9Sl9GVHaxujOMDCOCvQi9ig
TBDIa+9zeiURtbDkqT7+SAafxQdPvKJyhtcC4/yZ3g8DPqjZhkfeI/Vh5tnCe9ZKhmNhZRmdXQ00
2ZOnT/+RfIkxjpkja5Df9PwKFjDZAZHUSYULZxTjR4Q1WYX5+iX/mSxjA458oOuOARIQ6Roco1Nx
7A2fByXU6kINOJoLtXCdHqNK06oVLV+rTpp/XzhnjTKbvRh8MHwN0BLplBonANsAp1TqT3ct2bUF
O/9of0XgJZ3Sw6vsaskyj/3Jl2gru/ZsvCIcVuvvUfzPrMBq3VYoNKuKY+yeEGBcvczjaaLVepPB
bCTC0f0ARZ4rrCmOYyuCjisWvoKptK/vHALEAj3BCyN9fiUAdr8azc4fo4G12NE1iiyo9mtCWMIP
iawfLZcjXTIMSzoyAgdwCxt6xCQ/3rGBmNil+Zt6oRvXbC54zz1Xyq8DAw0qJ7olk7WEcbmxSepf
UZvuVVKc/ew/W1xR4h/Yi+Ea1Vr24jNOaaxKez8PSj8C/z9/i2q7SwDeB9zAhJU1NTPiMg4dvWTK
pB2kkTCN+R2FduLu6d3yr4RPxZ8rTA0BPoDZtUHKjkitKGyxN8CyjzHDrPIve4whWnPpa13Z+ZmV
4dHeCL4qChIkxrq3UPxm/2jc/ohHef9Pye1fCLsBmkXIJuB93lq76I+VP/hu+GCl006fo/eAWHhe
9UFneQvRird8kpp9gQ+oVckg5F1x6xN9VrMxCK6TPMQUbD5Srq4+VIC+T1gtYyYU5dyKdN/IC9uR
iiB4JIZqxUxavKcdzPprcT7lkFhY8yNCgRK2qiDOQLiJGt4+MONHAbDXpph0xYdfb6vzEY9bqbtm
o1vkkvzQJaRAdmy320neppD1GzCCxJ7etfavxW7L1PoPzgKiOij+NGfyEMIhGK/Np8NPOh8h5n2S
9VOyQGzMAweegKULBvujyMekjq0lj9XIQZcV+25dyF2invupOkglxUSKhhecoVWih/fL+RjRualz
PON7dKKBCtInvINZ2d8BGyWjBvsam/wh0VFxezkYdq1dvGAxgYRXJOLWdEaTeA5ouCrcnBEk1jhB
ODmoWr/pEpFLuvMLCAS8q7U2j0Q2JZobf1TjrHU93tGa4+fAXM2UgxmIltM6GhueZKppR6ObTXPJ
FIpY2jnmH5L8FY/OEio9rmfguD5djt3jTCX8kJGJeJulbuhWw0yBZnOakE5C9iIFx6kZq4O4xGDw
2vymPevhAai2RlciGze8Bg4VKboCPDQFleslulxyUagxHaDThUmlnuHer5I0JdmX/V880hUyvUmv
GH8ZhlTURagv6wwWTkelkXRw/Xt8f43ibd8fXrwX3elgc7yjr4TES2ucq6PhCgBpJnyOxqhLsLp5
lLUgWgjS6oec4GeNrpj7JzxHxUHwT5Wb1AzhGWU3XuuDMcFr0QsMDud5KNJpeRYAm3a4x5xmJ8Pc
CD3AdPyqTX7a/wsvYv2/+4gTdvNwCCcJRyXHz+DrzPgf8HCdKbYd8PUEWFCa6sIwTuelo9LCcSXX
L/3XGpZCi1mhU+E6QNcIDSueR6w89H6swFA12BNKUAPT5/LsXQchY29QaFtiryzprrW+05Ai2zZz
gsiuRsRZIf7XbnkzCdJ5to7929wAJ28W2Ln/Xe1hNzOEKeSEG4fDpiEqqAiw/Pk68a7cT9SbLKov
qQ4QZZQJrv1rMn/nz3hrLieVvaFFJeCJhW5BaoB4C/8P4pb2y6UaLZNIMp3n1Qfgdc9hwT4hkQNs
n0Le23JKffy+NVj/x/y8o6Og+ks4Hp28Jzt+X3wlBNGmC9b4O0Ryc15T67zamS2NB1KwNrW7aF7v
H+oMuw12WgKCU70LJgHjm/BFXc1vS3Sagh2x+ipKKI+unkjHmqBchic5vYqmx9Wm3vLUtbj1tF6w
L7zeqi7zyPHL4Q/cCsSlgNxQynRP8PQW1EBVCu03ZeVJFbkDICM0A5bXb/oU06jkz9nCl8p91lov
9L90RpJLfzFN6VJzyJuGMoLeuTRj9FespDcutjsgMuVHGZoTU6iX/cA/8nsbLRDVS2fAtNuMHkbj
K3YrJNy2sCk+mdNQrcC19pCX1tLrIh1QPjhpCwRtIgJEosKe5Ft1NXs42NzNHIsRpncPcph4zKtb
FwBcWzZg8ehZ34ILX7EtyxoW1rM+JwwHyQ4bsdxuutQJZzo3+eXAgrz/CDR54saYdjT4rlPcHVxq
qA1sP+hPm5fW+XxlyMAZ3UxawHMP9+OHqBEY3nuVgmyT/kWJtncS57+EwfcTDMHOQ08wN3l/Au6t
JNQFuIVyJKmF1UaylyJYLs5/LKLz49W3BkPKBl+CHEFKK9aPECpLcePlGKGK3Tvsk3Kd3WpD8AbZ
Z5gu9CTMZjXsPXoM+4TrS2GAM25Gel/yjDO4Ba09lrLoLQHN1oFHtML2NuZH7bD7+78cunuSsYMj
StzHQM4y7Oo5GCIuRYufOyJWw+f1FTgg86uk4Pbkqilq2SoqrOes3pIQk9wh4o9SWXqDDSnIdjSV
I8d2OfDVl6rxFWisoWqErbrGuJ8ciEs6yS8ogJYmkQbDg6tu1/oiSwxxs+CMOgEmTBUWsRhCtWPA
oGCgIgb3HyDwb91SVIQmSa5TnFIVGLRzazJIEmAcYLzrYkL5DMTkB2lOlfjPSLkDNwNfEN0FkDDb
Tkwsr4UID9+qGD0Znvsn1CDCIvZn1wfxw538fxaehJhgOko7+QY+2yk4YkdGLghumY8DYfc+VJjh
e13tAvhqS79/gtrcli42yhLkcqvKFkbNdPTdXibI4Z6h3C1InFyWRFosN4PLrsJ4KqM5cZ7q3XEM
3MRfTXwIdLiGMLRVJOl5cUjpMlATV7qjm7ctp3mOXoYy7r1DzU1ec5AnAQiv0ORx8e6ruIFxbNJ6
15N7GLyrnscEOkBQ57GKfNSAQngonSsQezl9idEmqG7VvHA6mW/ODVMh5QE5b6zVUz2c6JtKrm9Q
Rvzty3o7i86DRuVlQVdMRUk6GB47+yZh2BL1cRs2415u/LtvE1yrg8X1tXyTFMkxsw95Tl/XLd1m
eRkKnC4gFLsVG1nz9yGjRv2ODxmWDi2onjjpHa/5zrzq+/8mMRNUKvyxO0hl3aYqA6RtxcfRBdmg
Qoa32RBl6y9X//z13YdpHNUVVd+MKZB/gfx4ltE76n5l7CeDhI7ijB00MyaIOeRlpIwvH/4sJCaW
seAuC4XCHLd1VF+toi4CWNw53VaZOFmrR8zDehnOdedI89BAsjHLtxH21ZPsXX3vZ/cZrY8PDSQK
gEk7dCMw/CFc0+3ePAJm1aA4O0K0LujTZw7ecD5EsCydq0ZhWjao8yTqtFjjk88EAi4U1IFcCDDJ
7o4o/CuHaSPKcLA+lF39CWYnEErQS7bo9P86HMPVhVGuBDNJ19xWmz572yY9lZyP1FpEv6ScTuHe
3JWhyHC9oqNJ8mDIsiPr7S3MjWqUaaT4BitPLQct4DSsKvqFKajYnwdA2/d+j5JXg8i+66bf1uRA
YqVyzrMFxcRbyZXL8+jFDLInfwnBRlJZineZpXTZCo8yGANltKrCR9ZlUK+YIWNK6PixqsY/4RE+
PN9qod+5AUv3n/2hQE1ihaROqW7nkuIo/BcXCbyYYeVmaIeJ37svQyrTWMY8iLxVl+cqV/gAfU83
psWguuZoeZbjv4NObJVTPw/uFApd7pGfDINLXPxreErjWgvP/HwxzYNIEfwecG1Bwgcw5y1gvTwz
frQyM1gIHXUuEdWAx16gfRElnrwHnLfYxrext3eQKlhsafZXhdJ7LE75V3KORlQ1OtaJWbwBPLeX
w2ToYoqzk/+/siAzjj1rkX7T8qBfT4naEQYwQa38BxBYmBveUV2TssH48Y2Dhhu/bgFf9wT3vRYr
KTqWsulRXFlLC2ZSV+zv0fTYM7uYBfPeAWMfhEIeAQfinHj3nDs9qrSFK2UxacOBo0H+gVue+42M
TV6OgyvPqhgnNkQZSOlUtzErljkIngmb+Fgl18/KQiXbjHNPcG0lZzxVV5ZpXjatVAZH8gll2B2O
RBDDdDy/shy8rMP8M29sjbpCHq0w4hqvXAMypFLn1ndDzTUQDBfS2ji2FT5j7afprbtXRG33lDku
8u37BqsfaPv2V3x/XPZAZ0NgkiT4BnKUtCnTWJeoug0+E22EQvnobNN4z/YDs5SDch02nd+nciPC
2GmTkwLoYXtvlQ1clCFdiylyz6tFnPBgJxPNakIxRO89g6oDsjtNvrSiceVwVg5M3vXbRX2Qzq6c
beD+fARJkBHNcrTMBkWrbIqyqWwVADrZX8OGSVDQ9nw6S6S8WVMKru+j0PE+xoFWA8adu4fp1ehR
FG4gven1z6qnIH2urXEG3USfIiBRn1PU4SRnsHGLDFg66AK1qtb95VnJhZnTQvRSy2Wf1g/3zcG6
5ashXmj13aJXgxzs+nFNVxy9jFW18j/W4s5zG6p1FOAkQBSmHHm3tURRyWF23BSlPSNyxpN5JH8Q
lejKuT0ATQ9gEM7EBXeG87v3vIX5WT1UpzyGuOfN1wNqF3QvrWjpNiTircu0fGiUIDs3XLIW/UMI
4lMzfYd9oTMPxtp4XrYBo1RXSv7pbw/yoGqLDe5XQxGR5gcEB9eeRPKOgGmrYEcv/Wnv4/N1OrZB
/rDZUzjzGn4dEEuL2rbMAjhFOxdEk7pCOZH9kG0E0Rc7+EHWUDyHcUph7yZ7aOae+kd1fsv8gcY7
lahDpHuFrmtzUuL3o9v4gBpbJpDnR0TyVS48COIjJmq8I639+2ywW/4Yyu3s7LqmQvabvfuJpy4V
rlywOZcoV49cOt7tvTlmvg+vWfhbwkEpFVKrNi85zobCSUZZkQHVLNU42eiTLD2Qp4hPjEZNOp6z
Jy3mSJCbWI7bx+rvQzI80lr/iup+NzEjtmPHW9hWUR/8RHtoFKP6vGKUpE/ijDze5hU1no9rrzdP
cXQTlHztyIB4Q6N2BbPBP0S32Gv+79DlD8L9rWp++UYS0wPmPkSwMg7tc7BA4LlmYnLuci8tRRwh
thfw4aezAQQV6S4goJpKrctxjijPMveqFDwCl2kmrlcoi1IFpcoli5shLZoFqSHeUeb39Nbzvjar
3HDLCuuzzBzExJP1GQuyRsnQdPFb4QMGzM+nuYy1fJzuvFNtRl4ie8y6QUKJ8/g+sm7KoTg3x5Fg
hS6LyoewePl5dyhk+cWs1+N/jTk5IBFtpbWwerrlElXvzSXMs27pWnA18bB5JrnyzIjOLMpCTP4a
me0zUAPy254cZK9+IjEeDVaQIeIndQI1VWHWv822ju2LdNXf7RTHzi5hJtdBHthH4d2uoMp/lSJp
mXxgbLaTJkItMinz528OEQv3eb6RU149RluTcgQdACokBwpe3fDpq14QsBuNtMDh3Id4lnGnH3Z9
PWDahe3oAcwfnIwJww3XgCLA84v2rWMN4Hx6rHQgKebTfVaSyrvtNJNUmtxefdupTaEi9JO08M6S
o64nIKBmdjj0fn+qg+s/STrI9Yq89Kooz5tVI+htVakHgLUCAOQB5979DyfV4/pTDBc2ZCG3yf0a
lpiWJZnswDj3WXFu5gdebjyFhDDiFMkMTgA71tUvNLbbkkOE+aZ2jJG4i+T7gJqlPt4gDUj0oyVt
sjunMWS0Nt77+ZqD9nvoTD1lTi76drIeTvP2l9Z2cyzyW4pLP7Elf45bd5j/+2uzDdoDMxlDLkDq
WJn5tqwIoBOjiTe1JscH9H6SwsN0+7on2gZ0I+5TxPxo+gZarmcbiXPurMyYjX8LyEv2quHIsIUf
BIfoRKJonbkolQHJC2vypF5JDX1RxTV5TThLKni3FKuQXcz7dMPF+aeD2oud46OBT1wp0Ej5CUCo
6D9w92MXViX4F9rECtJf0UGhM9AO11Jh+gK1ha8aN2w7vebP1jHkM6Zp2HdeT5zdbVkbxdjN13ke
WvKj8PZdW/FKXCdKRoCC6DFWVMX3orwgdTXfFz1Hxi+cmVMuMtOJU3fUAL2G+lFj+G4cLOsM9akc
V2Wpvx6trktzx33IOeGzKlt+aHQtlxLWVjbYk2mfy79u6WHFu+DVjgkWgJBl2VaNhPZoZwAxfu68
fW01dV39FKCJmiTInWTj5OHoEfC0NzW0I3uqQlHy2xlfUYHCyOnsbvLVZPofXPn/S09ToggdZDht
a1QMJryB59JTriPGWnReAZJPfQ5htS24KOrV0LHaC4UneU8th6gPGESUjgP5/VWomxqXgqEdh9TR
dLe3czBlXNVq+sOm9ovOzABE5/nNcgw7UG2F0yexfeemw+9LAj9Z47pz+XDvxJCDoZjM1Sfh8aBB
3qtBjN2Lgoe5hj+aou1BO1sI89Owlg6niBULbqQcUL1JVRVJZxSyF3DJakBNuYfYp03uXh+RgTBH
i7RBDfo9ESmvFgwmfZTaQgjjKds+xTmBuJ+gfHGRqKHSpLHO1EO1mUYLEXMQ+U4iVIUmu1kc/XQy
U9H+CEZBTatIT3Vl0W0PxLG5wQTkAop4jSGNVmNhS8HlA4wSZGT451lvQzvHSGQBrxsjwVPvpGRt
1RYTuwz3jT5ezUFobw2DSj5LcXMwboIqqdllLeFNscTvCs0IzOX69ApzDut8MMmA4RctUX3YtTZN
WgCnPlvOy72JvC0uTyVS9hVPrC8rIr1bGXKJUw5fqYZ4n03VtXAP1MnZOJdvWMaJCCg1lznwnR4D
TBGKGm9435slEB74Rj4OVI4ZKAP5ur0EBbt+7MB7ujGDJgdCEDaklX3jqyznHqrqYgAsAVgtbUst
Jyk8XNFWWvjYc1jPyw4Gb6szZKafER8MBChL29i+/4b+cY4xTjsGNdCQU3KG26G6Iis1pqHMoDWT
J5hK0fAaRkzY76s37Qg+sy/EOIQXo/g00hAP7QVE0vizwyueb2AltcY8JIOV3jkh1rkaQN5bKYjk
4XtTHfv6/qDzTHovYOf2IIooLViaIesuc5L5w1dcMXL7fbRCjckz0WoaOoFkasHCqwPw/S5BwV8H
LkUJizr+kvafSN7rrT32FkfFp0icbB/q/ZD1+xWoZUbXca3Es5C4/k/qWljhpcZs1ytRldb1YbpV
tcY4AKJ5pFJP3Qp3J/6U1Ul7lLBkFQkiyJ286uTM5BhADPtdrgTHaUzj6E5oyqktox3FeezjcsLS
PUMl6UVBF5B2ghlfh0OKpORUP5op/TNIwFFEclwsdMlBW4ux6p2e4AVMlNOLhC339azAdhgZDFU8
xg+481S/rhLWEhg/QuCgtuqGsvFnCtdKt29w3Qi+UVblaRpyVZW5r4j1SHe3NuQ71/kVnQ1bFOPL
9HBhlGSt5Wh2hJOc1RHyhs6uioWdMho8ER0gMewu2+uIaGkj4Ff/OzH97WciK0k0nRYucd9ev7Yr
u/iSZb7oasM99z88aEOTcMP5jBeDnkKo2hOdgCpeLqA2BKdIdhqQiNVqyd80/Vw5WufX7FxOySuW
mmfV7O12gcOiVMUM37aEIOUetE3oI0uUBhokOUC5v/F7UEYtOetwXjFK6srtMenl1k4hbKygubuN
aCDJvaf91QFufaYuB9XEt8vHtbTQURwjgQJ6LwZ0/3ADmHI9hsqdHwRlt/2boJEut2RP7/YH1wym
DF1diuLwPRFqtccAGO7wMnY7gh0q7fyN/qNfdT6gvJl6X/kq/HfhRNmKJ2yuj3rfkEEKpnLbSr6v
1TPtC/cQmbY1qSOksDLwhzREosuqBUXna6DJsAMsFdKVs1+FD8fht8IojuaoDb7pFEdfA0U95qcK
mPXou05ax/I9S2TAT/AJTi+RMybz/h4IXD2FFtGbOVwDoMoPmotgHzX4TjDhrFqyO1/aXhBAf5ge
/1BoYdHyJMtE+XpfQb3Zwnq5Pft+uVyUAxWGkCGMjpRx7XoNXJglOOZCr5jE0HcTD2S44FDucg5E
Hgsva7daE8bDCq7fF8r8/alYmx6OQ03xkv1C27sIkLaxf8/6jruGyhmwwFLo3lVZnoZLjc0FmFcc
nEZww3F2kRT1H8pqjfLg9KApVGisXDlTK6p2qZT3SjeuxmyHx+nDNkNmbKfHGMPPLcHHhDjtq+91
IY8VvO5or10/JwpOj2LAri1vuLwHLBEzmqNnKJGlAiIB3xz6uj/Xprefcnl9gcvjpf8yU8OkDx1F
h7bliLgY/x2eAL5gXXbfMmITWTf5IVWX34fkHd1AncudCxQYAqjeO4GrNHmvz/jdgmOKI7zONZHP
bg60CCooQ9Kzfp2F4I4kzLeEYHZdTsqpXYSMiOJ3C+WxlOuH9yrJKjVOxQ0shnPsEP8x/qH6corg
Js1GIrkPJ67JOU9m0OocIcWzPBGr+IZQt0Xty4BG3WQAAl2Hd/yKr9kSqq4jVd2wKu8btnOe82wl
xgIu4Twlouw3CmliUybfVh9bkT1wvQhOpYER/fFNUOI7T21lXnD3RB880Q4k1cHdJqvYaJEa94Yw
Ya9B/+oOXiKSwN1e+Rqw/PX5h7xtcFB3MEf6wD1TfAYF9gqDL+YxP51O+YWCClEODhy5wwzb7+Y0
7bvcVYqcK6H9XMWBvhNZLJ/iJx/bgd+ARrpHcoCdpbc3TtzjvAEdiL0FiPt1Bz5T/zLmQMcEpoLB
D4y/GzcoCOrgVR+ndsp9xTTjXBDbquW7Yu4KX6KbM2SzSi2b1YQ1NrZn+YZMFUfDxWPQaFCKRqLN
zPGVKZIBA4IcgkmaP6rzOwLbbl0tRvBJ5UTptawJ9k3nDW8bdSLt9Xxtw4kSfmXJM1UU34Y2Gu4y
h5lLhgL3I9HICIQQd1Cvg9ltHWSi0Ux22E4OS389eRl+pPb7nLbjmnCNs8zM4GwkJhEG5TznqK3o
ezXW6dWo4b6YGdH2Q2lW6Ue1qamHgk7dlCeJpmh8yblhruB7j5d/65ihuUkPGJ05FSLPbGNcn7D+
eBWWLduH+cnlN3GrQl5CUJZj5pdfAo4t7OvyKo2+dfUmaf6dEYiTKYluVOm2mMXTvV0zLg3dJyPB
YYXbrgi/LzPgz+3n2kf7mnZW85k/rihNrOV9bezQk5ZAb0ZHJDsc6EkcuS69fw0/HwYmJCH/5sVD
h/sqjACT7ySsg1MA8nwo1EhnC2EXupSYL7hCjTMdN9H2xh29Z2RfGH5eZO9lqata3ucnbJ/gsSQ/
YwE74RYE3hps0UPO60w2bEt4fQ2Q3MsK92mX1fiR9xc+e/N3aD+wAjrjwRiIpwfav2V/ivQPTz5r
pNQiwlDEZKrv3nv5fb+ePjFdEfV/tidDdBtu41SoViZq0aOrODXImjfRqVGeHBLnS+rgXH54PVpr
1iLb99e2qr31PpaZKieO385aFG13DaE4iUm3rVLHZiGTifZxSNFOfSwwDQUbfzmmUJTLxeclo9rA
dED/hshyc1LPNfxL7HQyQysfjsrYu5U+Z4JBTCPhcg7XDcqvTcfp5hpv5kxK6dxj1kxLPYPxNIT4
ZDDi+5gFFSDCaAcIXV5IdcsXlw8GwEF6TSF0GSjxZEa7kZfkAco2WiMXwoAOGFbeJSMtNrMDdXn0
9/t80b2T19mKDacw/2bFPdfL56rLqldmii9N5XFlUqf6NRW9RZca2FrMqLTc6c++ZUPKC/C0lbsb
hi0TiZlDOx5lmJzu3JVDyMNKRiZ9ufrNDmRFVU7Kjors3IjPyg/YyYeXIMCoQRZsFjPu97+ale/u
zVyslFJ5dC375RSrq6Wr3kVp3rJ6fz64vW0Jp/oiyhbD7E+qvt/pxUdtuFmdVbh/fUrCWlg+fKqa
omgjBC3dvIjT9oJWB57ro/NCYuW7T7OT+f8+aAp1DbHX4zJU8/s6XKMxyx+XdTFjCAljlrOX8HPG
/3wRHePNMWtQr3PLKVBO+1cKU2RQvvVg8+Nrdm8NtSs5+Y6mBecpxJvcmTRatvz2CkqtmTHMltZY
Xx2/2mVmqGY+96p6Z7rOxjgm0Acs/GS7ZtNzBw6VNeDSoi9xQvY3hoOIymvgZpBf2aHT1i5FIvg6
yeVz+6U538PrA1E4fNrRIAHd6XMoGuu4pNiEZRmvhJ1qNWjBGQN3SFGs00srr15/myDrBYUTdAp0
q1/W12wyrlprvUFJtAYs50cHJ/RBhpy4r9UHS7ACQI5EtLFxeTDojoh/+NtBkMeIThYsPREwihHi
WOon6RXqUAFALm3JsYc1AfD+BjvgqUoh68gyKA4IsVc6rVJY3QNDUnQvecd85CMKKnyA0fHBr2hq
tRa4jpzw3mhWmmV94xPqJYo5mh6KQkVeWKWjW9CKCLwNsG8cBgn89UzF7xRPAq2jqgpqPh0+LBSn
41eeJj0aABHA41uKF12Hl3rruAvgkqdmOI08DKwI41ZpYvmSHf/MhdRYqiM1A8fqRxOna76XQmBw
/4fD4Ftrjd5ONxVSs2FjxG5Qtjcc1ffeuRBbX+XFsl9rK/l2W/0mNF4rlQqlYS9FKtsu+VOYKXnq
75LnjeAVxoQ/buI12T/LSMxyboV00Hon4xhkj6uUxuITkSbYXuLVvFUPbM0J1XLZQhiTgOezjzT9
R+zxtbJPeFT5IsQ7IYU6+du/uf+0c+3Zw5lTGIGgDa531O8PnseEY2zVk/urIS8wBOhBCsuibnoC
18sVuX1Z9NsYi1z3EkwVDjT1xt2xPQDt51ZfwMjnMCia1r9d7srn4kKMkiKdzqKsgG/ukrpJwNeM
UCHY7Z+x/dlUnQD1IASJn7B3DlCVaR7fYJPiz9e+YxBnj4rhOybKpsFDCulByicOVGgpU2X9nv92
C8KkTdFo+oMwExIXFvtuVForgyMyl6NDQd+C7r8yk1vbIMEQM66isr0FlUVDg4drDcgWPEUPW2pF
/TT18e/e+cB2vwkfxtwtshJ9Oc9lLMQnUVQbp+cKzb7woeKm00vgwfVx1IWH/Zk4Rsy2jzRPXruw
uPN44fM1ZPhNdK1lSl+Q/3TQACxJ4UlbqLK0H3Ak8XtSpXNkezlfXFbjV9YL0GGUP/EUpotpsuP8
jIXhQzAmBjXAKda14u7BYKO8og5Ioif67O5uf6Vid3kFuOCRROZCGC1tQNbDbCNsoOG7pzTK63fz
L53Y896EW2bS2EuaXenkcEqgIhcAKr5lwao1xNUQcdUwE15KjkWuSb8WBH/RrG+MlgXCos/AOhm1
vWULc6xTUJnJ0Q0ZFDzaXeEHbHD195RvLnxkrLyrFsRIs2rkA7lWgojZXzfkmQZ8WHandt21YDU8
Fxszq3dCJkf98E6W+VtFhkF9dLmL/oJF8p7Nj5ddu3gZ9VXvIvtA6W0NtVNR0XlgEPRdr+r3TN7F
dmOuzn8NDuPQiqHVfGOxAwvJJucVIJ9kjUoqDzhgPB/J5DFmC9gvjU9pEvPKpn2IMwSDolxphYSG
3MOP1GiCTK8jbFSKTfxsrksa0pyEhKhmZYMoB6QAb5V2J6h+qZ7Y/QmA/QF6EjWmcvk4YJ7Nf1Zz
ntFfvK9/VKMB/wj6RCUYrNyvwk0TAQXypYYvN02/+zI3k00fy6CLfzdUQawVg4V7+YtuaXmAwArj
qME9JfYq5zj9nfRRa5zWFTlrhgE+of85SAAjc1EUADVbCoLeazLg+BMiggrbowAE8FqktPG+2geE
3A81o63SyUmuGnNp1d6E3QolPzigwHzKcMZtOFJcjFP482JY6DlOPIccPneYNp1krGWDFR4ykp1K
wJR4eZTlfrPtMsw6aRra4ZNJyU55xHbp7O8SAf+i05JQo41Ymel2yaMFvzO4x3uQgzUeFmhHITRw
wNV8UCn44FZsLHlJKJgynw1Su4lsugiGC4mNe9LtItnzxRpupnhSIYwya8mM+l+dqYrSRyhlSGG9
YJNeR9LMD0gcG229yAYw6M4b2lXKrDqnQdGX5A7ztPA8BPdjI4DCkt18hbJV5sKbBNqFdbJFD+vj
QeiMjFtAtaelZpBCD09H6keGipa49Q32lrygXh7kUVedKZvZW33qjoBtRMwfC/ALx5PQuT8ROm3E
kGjcf9TTwQMWXbkJfnF5FWT6w7HG8b9ijKXy2j595QfegOLfJ9vRLqx+W4S71ZB7UuSJd74Uo4hi
mUWwHBe5wNEA5gOLWdB9waZB2cOOaOzI1iqbu1BKOWyNfcYkVYKjtQ+AZBA0oEqaZ9IbrCRhz2+3
ri8s9Nhhd2RFl4YOVz7aNrb2Y53rlb9I39SvJnNszwjyok25IIO953FMySQg86uC9UOWkq13MWI/
HC88LgY4bUWTFgGQg0FWGiNIerH85Tn7mnPu45HXdcaIuKw1BvEQxhpVrSjj8RC2Y/Ach7zh/CKs
bKt0w8RzemvGQmQYJPjf9QaEnFodsLsdU6wkUYdMEnylD7t13ot9KsvPWaWEkRVB7fiyq+ljEQhk
SV438CvjYKVC0z6Vu5gK0E7jOKolSaoNqM9JHpuTw4nK465PONAKhpc9ZCHEWmm4gwQvnD3AHUpa
glplq2L61ZEonXk7dik0ZWK1E7yMZcMJWXzWfHjg84sjP9zuTiJuGMx0cXYt+RJhp1LWGMWLZYeD
AZp7euXEoG1Nf6y9s3x3bCtxQYiBE6WmL9/oPwe290xcm4paQAFqP9UC99lyTNx81mdm18sjT9TW
LdRY/ZuVxuguGDYr/h++m5828FLiew4p2n4APciliqE64PoP2lL/gbW+Oy6dX9gDCVoHNJxt80m9
hsI0ANZ7hCAUj96h9VqdCTeW0V+YkeixJas0vBd8jmUwHeK+CQuXQP9fvoejB57fw+Mf6g1pkwCX
5knnWyD+EUrJe+Bwvdaucqk7H44m5ydm6/ApgLz6STMBFPVFu1zNOSNNjENUDiVJM6we7eQaDE9/
z0ZPFKM786UE5H2Fxa8hgi/+THkqSiWxNRP90tOv72S/sO0VWv2+yxngKxNy0rrpPNOJ71Hsc0H2
F+XyY/dopQpyUYbaEnyKoK2Rxv7PJlwqV0dFifolm+EEN6sZeY9kl5Zndn7rFcxX724zfHFpPkBE
1/K7Em6nOl2ywKx94q4E/8Ymi4yCz3rVRMcun1Rn6jQVhLlk5Y6Rkju1Rg8balMlCeuUkaM0zxfM
LlY+uh6hw9nUfFCNNfmhz2PuwkHB0IkTTtfr8dWW0XOAfDhpPOby5630iP1unOxbzw1sWRTelE+d
RsACira/g1vSjd6V8uJGxYMJZ9PXmS776mAYkIckJWIWijJkmxAVMsxQDzrjWuP5kUwPmEswNJLZ
AOgM05mhhgnJ1Cbzwiw5uy4k9/0V/P1IZ1Qv+IRGkUhkgCU08HfJGvvTQwOqIkSDRaZTqKUjI5mM
/e1ymputt8c6GyfXhmsnCyrIX2Cy42yOJN6khgVEJ+v3ZT4b6fAK6LopnE9v/i6RU6FOFmd7reH5
rCrbD02ugKv/hUtOO8MKyD+Ew4E/vVX2b9VF0n6nHQepkfpedyjcBuOOQBPnI4Gwmiue1SiPgPAp
3qWQ8jIpE/yzItDAQJaQ2uhGJu3uy8OPVLAP7dG49U59n52fyh5hQ67Nh+p2ISMtnLW//HDpsYkn
yi5ee28JN5NFExNRoS62uUOiNR2zF2PQZJPxUvdqAt8IcvUIi0tXr0rsHg0YbUxjKHi4juS8zH4N
22+7Q29E2lBH73dUEpqKrfhRZQ3DhfvnQsEOZ8Rt/n2bQ/i4G3RyBJp4MfpmgF7SZwN9D65EbfnW
VpbjROwaHRuDzhm5Dn0r5k7s3WdjOcjtDMhdXgdH7+6+eBu607M/S/2901Krms1ofmycTDKcoq5a
MoK5AX8XwaC6EWhXLznELv3JWowNB1tg5DGZyQg2ImpGSfsx6lC9PZ4DGK87X3E3AmJt7Px9b5km
5dYHOBM49QU1keJ9lcTwFrwLVGsQmzPhRqfe0iFUqswtCwxWbOIgQOSkft+n6xnXbzbGNBqvI9Hw
4vHQsX6cwEWWLP6Zxg1RCmE4x0IkY0swRdDhtGGbWghs+MD2Vfy7iY8J1c6unqDNXvI46aDEGckb
K0/q5Wv8mQJ1kcwht2RtF1R8D7ZFdltu57fWN/fnNqTqZT9UcsHeXNs1RoZfLxgmAkMvVj/pqD/h
xTyw+yS/GPO35lz7ps+wlwkOXUIfa0artJjf2WuScTBNchDlyWCOjdfqjG8IpwUtAr4NgVjKfn5/
OIYXYRJBvhhmGAVArGhcEbU6BiEaSFlqHWQRsxPiYVuq2v6J4nG+9yPrzWD1vCUivetFMzH8jVDR
O0Wr9mgkZ26PiSYmdV4XM/v10oWWROwUS+ny+R3OzCRCDOKvQVnddMUe9zRaKyjtxSBcqHN6Z5a9
ibqJwrfNLZfI52teZ7Ewl+Sub+UfcXpbG1io0hLlUXQOAlv3W9iZ0yIq0uZTuUnUVPnMMyozEatp
OlAPdof7xDxI+CMi7UgEVoncmqGIJNTT7tXmAkahtPROhSsX4YOJgiIYgfvUiGzwOGS0hp1cYfj7
lD+mNraT4pjxyAYriGbb21qAw/5KshdOPiC/OTLg90pjCpDEs8D91C6A9CySMTcI3sz554vo24o5
5SbeRNleTRo293A+zrX6F9KPP0iLLlivCITjwqJtgTD9Kew5Ze/xrAVJURhJuarZNAOsIi/YhP6F
h2Rsj6+DVZ7wV2mMdbVBQtzgCVSVEYxLF8u64dm5C1yOwYWBsHDbIDiHQ4JvLgtvDusBPzHExlzl
TXTksa9/2nhv0hVLQhnanLIRvc3UCGJR+yWB9i2H4bVOhNQDdS3/j+8RvZXZCgHP8ob4JwFsYe83
/m/mMiqrqCJy1zw/TEBWlkiHlgtfbtC6DpLs1y4Azq8LfLxchWtsp5YV2oc9pKL3kVd9C1awBmr7
ItZGHiA6GavRZV1xSyld41KMP3QT+K8xrCRNvGgk0b7zIQR8lkb7ASmhtvN1vAjRiuZtyqzLpOxk
AU5J6usuZIP/sliNmlqs3inwBKi3HYniOPoDKpEl5drEovNNisvjIhJ3Nb7TAKiGBLEIl3lzOgPr
CapWztA3PRSz9FmIrwe+683hSGHfGRRFRgrzUAiXGP2eevTsQIH9eLsi+uDgralUthxG7Shg2jbr
8LzmZxw9COOtLR/1sc9l2CfxO0fYqs6kUurqj9KkHxYkHlNp7q4AahHRcbT3lajWIwiVKDNxuYmu
QTAFQl2fScwKREUk/+IulLy0NYrQaqmVHR/WfEgCffdN/cyNJBDp5d+wWGlylQp7W7B8BKe7drva
5MNIFyKnbKbQCcSQwZ358EhAHHdpsFAAHaeOFtCfBR9oMHwqOMuQhnGDk8MfTVQ6b83vnSmUFLqF
+dP8oP8JF3mAfgJoBID11MAVYAfjxg40JQY/xnHJeQV4QLei/OPRZG66YNHz16efhGktReYJbRJr
dYe5wcNE/1bLyIt/pW3oJyIRSxqsHCqnLWU/wTQpwIqqbzCX5xPYYTlQ1QxHC6NrE0AgTq3SCZDQ
oL5c733RKcDXVm4QyzdgBdyKWdav4tMwVGqg0bxjFFYBpJyYuE4OB4BtjkSUNLHlG9Rqi1UqbxkD
zh1mQ8fEBXcLSboG8kc/7K/rkrcToHgINjrMa+cg/2LoUIvBg2SglLTVq2L7j7/qMzrbjj17ICU8
KwrIY8YIY0VyPERpPTDtkAvdeE9t3yGuOIxCQHMMy9azWxV+5xKqTno9p7zNpmdeJUREnOnAaMnp
a0qCi8CI8SFSHOoqvQej23eKF0EO0HEwFraWakmFoNCxOODGDX9ku+m03StD6SZ1O6EbEiOMzO4O
B7XoHOKhIPpTo+Z5JOXjtS0kqhnH9TWZ3WSxRLvOnT2tKW2QRhrcWTATJcFAYcuNBfUGKdadCNXq
VHnMnejuQL/8iKgbmWsCgCxhqCfkCedn7ydVQjRDj0DU71XFfKr0+EG4Bh8Tp1gzuLHNJ7QRNG7q
Q6ghcsmxMWdILezrUFWp1ls4npL3UiU5qqt23j8FaZGsn7RA8J/13l0ysz1/0v3KrNJAIddZhubo
Q5MrDuFuivVTL7hf31yXv/Q5A3ELs/+ios4ChCqTwJT7Gq2sXVjoKXz4ykmuDghIVS9qlzCCQ7ca
A/JKFuHFK6EH5SjQTnX8jUepc0siHOfzrS6b7WQFq8mlWpMLO3UNQJs0n88g9Gso9fcb3nai0Q9y
yjz/JdZPdynzpbuO4VJkpxc+CgSMMw4d2mI8lh7E18L30edjbx+lr2N8CrDigHUOHlWbQ355Da1d
wHUp9vvT3nVroNMri7HtbCxbeeauktBbJwO4nVlmz9PWMzZjXy0LKIS1VvQxsbvDyhyAtwKzDtMB
QZbvA8qWDjSLD9XHFIbClcIVD3Ojr1iM9PPzgnjQ5D2A36dtPwgUILsVR5HaNckYpmihF0QlMCnc
a8NHrNSieh6cJBCoDwXRWibPkxAvr05TyjEhcJMgG71Wl0QobOemgu8qBEFtYcO5xyyx0IUeqWMp
Brhsyl5J1MQ+2yl46+7GAK9KFz4r3QuEXJgZCzal8O+JebWlqDmVKvT86BM2tCBjHi06sd3qS4Xy
ZQwUqpgPJe+qUUiV3pmzFSOfDchWQhL8ds2nLqC7qfZcbmULgiZqrEnPwuC+Lb/+a8FsTEbNWu4h
8Jsopozc3fWjFV1qpu4xiajkc3ArgqqeQjC/YtTozWKHj2FOYutfjnCEXME3cXhjheF9a6fv4Z80
92BK68s8rHb/dLm78AasfUJiwYFyj7jRgTxwWpQLHP2sLKXtJAxaQHR956obzgFKpW56lrasiL/i
ED1nTXhmKEPX2HVw+ku8qzd4gF9B0J2W//6D3r9eCIKzqr4HG5Pd8UHzYCK5u8z4VvtMiCk+uwm9
lxhRdIZLJfKB81j1Q4FWWoEd7VHO2UPv3NdGAhOQc7PgYM+KfH67M0D7kJdWzpSlwC2hOpoyIeSv
quJEKLC8VVpOoudcmWZHHKxWDsxdiGi+xfueN8TQ/vHpBOWJKiv2Qfayjkww2pEojv5A+ks3UiML
CxnFHmbE28wXdaaSwa8x3B3oikwqk9e4JMOjmyKqjtJ78Ixe4+9x+zuqg5TbzeFma9gNJApeB1wM
JGfG7HrUF4MbcBZijK5YhxvEgkTXr9eiX8TgJkvKRJ3hPTJsOxizf3RvwjRH4GGB7409UFEKZ2s4
iA9swh7dm87pU8tDZURBW0uUJMBYqUjlK2mWr74ZywF67HIEozrLgs76y59Xu479HlB+/7mkYPF2
vTwy5LBc+Ykj7JOHoZXg9hZFBG09Qd4S26FN/f6MmBaQxk2xTF/8v7VaqNhXL/hMWa2ChXWY2Bg4
gln1KgtAEs8s2vYvViYEIUG0qkgKAeMxdTzzzl1NPKQeWFZ6XP+ZalPXupt0kmERbmjiuzjBkmy2
K3fc3rGBFJdPQjVfdpm/LJPzyLyrcI6f3Ignl5ZVeRhaCWa6BpSaHZQAGmJZUr4ulJN1JBm/Sata
TW8IGaEBxkwu6msQ1aIzS3vGYjqklzM2DRCwa38M8fo0Ap3J02W9Dgv3OEzdSU9DeAaxrYhRSR4D
zsLSRtq8rv2ySWOTsTNwR6CEh63UgaKfhr3wuj0g1k/4SaHdx3gvSGerGd0PCnXPOfPJ819CZ5+B
EhM9ucIkrIyHxezSz55uy1Wr/oFEU11B+HCeDAhRly4C/j/qWwCrXdW3f8v263mBDJrh9PioO6CW
EZjMP9v5ySUToJbjjWH8gj3wYmvu09iqTzpEQN0BrFqTsR/iWHdgKh/Hk6xIcgCGEIUNXxKgWCHO
sq9769VxVSK7HQLI0IjaZoHmjfzreiHwFA89J0+1TyyLYdMAK3mzcuwFzxRwtW3pX3nhfntyv4ur
V9DmJYRJqxhpLetSEBJDteHPHkoMpwZxRgqtk42oYyYtLLtG2fADq8675kOIdLklvTVBB3EQQggk
tNbuB1w8vajl2X/PCFfT+VNsnuhkWrSXOFV6AiK5ieEZz2zzNl0p0S9mtT52/3fCDqOxTyViryLi
Qmo3cMmOyXfhV/N/OFIxQaGFcrj1vrhrR05oeQMJ+LOWcDqdPwvgt86S0WaEBQnKp3kCizNPYbsz
K8aEk3gqGDfKSZ8d6acjbur7zfL772kzulj7WFCxJBwTEKjvZtTtDDs73jx2wiIYhgWRIdLJmp5c
cK69fGbNnNjh0MkJh/JMgTXllKK16eK3mT5TS7IiWWrUgxGjG2/H7V3YNOqA3nMQnRJHSakS9BBj
7JVBaUUKLvp3xae2joAOz0qELXtxDyzD6lx5wRbYqbxQzxjilcmP8OUH83i6npE2L4HZgk2ja4hr
UmusUn363OhNGEVK5pyJmy0YxJqtW94MxmtU6O3aJe8a8pxJs2uvwYRVa6yUspzjbiC8Xc17fwXg
zFH1TMnTyov+YbSG0MKOfqoTA7i6+UgYQJuL8DlHuB43mF0QWjh5641LTCHB+L9Z9qJkf9xzcQ0E
HQ2nttcpyevd/CPuZsOrxtm/E1T4KnhJUpBLTuW99IU05r1toQFocDmmudw2lNTWdfMXrVWYDINB
8I4CJKXWUs2wZ1kS8HLzVcvyDu7dFFOQVbTKM8DzNDxau2+hmKjgriC7qrIFKt8CF60sDJ9P3ZB7
xeNWoWWcTAdrrO9lHfQnFw7QskCSZrucY3hZaaDYGYCzmfsv2hVh2UJxQqx5CjvXgar+2OfctJMI
4HqROABab/B5N3YhdfLhAo0jwAfKbTnKrhSUT2tGsuqzXIxC7x1kUW+MT64PODfONedY+M7BFFJV
6FV7y9EGJQPmklcFDgpHaT4v70CS39E4W6r22L3O7XTfEJm41VaqJy9mT0YqTCGtW+410v2RS/3k
gSCRtDxblC+GQefl6TUqPkPI6Ho507MIlYggq/ILjQATfnuqZYZhrYDYZPouBhRAAurENHeNwbMa
ntkjb9L6z7oICVv10BGKNMoYMHL7TEpzjqDcdUMAzaVIyurI+aFP6EYMucoExYaMpUxYNyn/JPLt
EPeU+lWpsTGLv0EJSDgUl0iw2/tpVFNe+Zv43jqb0zU03i2fdbLa+5pkVqX7/LQuqMEX5b14U1ae
JBCRZ5YY2JTxs4j6zrunuV+aa8PyJgMq6c7IA8Hqqh+0SlFA8MJJxjeiv22jEytnPSG9N4RLyXyg
vwNsPwKTMm1endpQNxKE3rcvrU8s2Z3FSp/wNG206fh6NfIfRhrHBh9iMBvKFQ7hSQ22Sq3RMVQj
Bz71pd35P1vtRwN0PQayQwVlrUnNazYsvs2nqIORDfvshFtzkjC+MiO1PSxoRByp6HDO8JswrFFc
Qp6c1pFoc1i42J4QWqasT3PEQyfU2yEVlodI6CleKh1U2MkviVIQGsCavF53PVCn2KRClGQPThd7
7LwDv3Qqo/C7pWV1QCxYomeO2H8gUqTYF9Bqd7koBV7tFFw77HjSLppusZBxMa6hxvIgjqa0eUc9
9Moqup/MIcJyQjgtOlJ6pPFZi3J6AqavfqlmaM38vrFn0vPlDeRd4V6OX8WQJzSc5H7g/8EoxRgp
eFgi95lJzFR3heE1XEMjb1dkfK0bxDWJUGQMcxnPW7uws+u1ctXSDvEaojxIbAnUGPXH/yRXx7ev
Bp+m0ApqdCwx5+cW05Hlxy9RqpuNfSna8IB8Z5S0pwLixTrRtjxd7obzphPVSUghhBzdf4f2+1kU
i+mtZxhmLsmEMpV1Bpf89ybcuV2fwhYqY/UT26isVTonzfOCsnLSX+30vVxS7MfqHNZsb8ZztoZZ
SnadWmtGTqZF6MZYXAofC1HILVVAdrLblijhgRWnJ6CeJSQWcuKYTxJ71Iosk0dwYh9ZDPCKmbJs
LdhoienDxo/oO5otAsPY/XK5xUM3GnEIY78wQrjQyD1yf/fZFQkVURN+r6xK5RbIvoIZXJmP14y3
T/IqzQYF4vlNxNDO4ta4W0o4uWb1mxLX/xuThTY7rxAUfAyVZZM0iax2gnx41SFqvjv3FCCgKnqC
PJewthFnnOVyWt9y4Mj5kxBgoK8SlteXOVLgFLHFTpv1tStPt457QG6/XoL1EfnMawKFfw1cT2z/
ZcM4HieuFcoI5LG+w/C9W2NbZySFr6JRx2PA9VOwEHAc+gvRyGRXwYhFrXreqkjQHF+hxKtyx82+
aIOMJxkrfvmt2cZT7P7fBYaisg3n3zyZhcLCB04fkja/LNugGy5nu34h0pdAGcIb4Cer7bSHwaxs
kCw8K+IqZ2czAWkwI6WGgDqb9xuT+0aspdadbjxf0MiNnieK+PvktJ9SoHcMOCq3MNeKi9PNz03Y
fUpXb+6yEVI2dP50Szt/NqCN0WLYvqeIbxpc+NSOTKEOW2GCXRBjehlxMCNP8jpaQZbpBTakUj47
7hcDmJzC1L9Ri5Ia3vpZotal0QZ7PPufMNmQRdAjjnvD3WLlind9Tnd6b4wmgdrP9YOvNaiBylsF
thuzKYH1LQdrPZm0WorZdjhP60oY2/rDAWoUgQcrTdqfe4qgOSbJGfKFg0kumMRQoWQyDjprOOOG
xxOxXkdZ52CtgfrETOLpC0KcfzpArvcXVpOUo713Inv3wO9q9AY9o/JXU276ylF8zfrk5oSggoqP
XKkdMCu3zCkCldpawz4Nw/Vsh2MXwlvTFzZwQEhShjTAvDA1fiwKmcWSWhodaYrtRCNmrKG2G2QB
5CepAY4jtRfiZwdSSBo4M9XCOun1D5wAkKaOxE2I2NJuRB+0BjyVCsB6xjLA1Ou7iR1tX3ZDbSC8
8AkV9lr1ycMH+mL0/m9HJbQS2xBO1PUfgiDACW6nNDj65M1nOg+sNaMzG6Xnp04GKxBPu2zbi2Eo
15k0ujQnXxl+vBGHb/Pij/9mO/TSgFmkFzPa5kat0xBnZemY93hnECnCsw0AIUQxOUrGR0GMN0zo
GWgdDH5EMegeuNVC7uqmknjaSws+kNkaG1OLn3mjR382B9ACTdvaI4zhmCQ77DV7CRVMykkDzvZg
JChw3IPWL9zAbE9xsQ6IpEomByOYUEReJdiZcEsiHDV+Kkmz9sM2NXwUGWv3u5A1VkRCRZ0BWv7D
UK0lrBbzMIXAGL21WpfrS55aFgxSiiRAMqetnSXeUMRRHHbnDLuQ2+Kg314+88sCtuxAUM5+1FP3
6EKIA17GXt0Bzs18/+QuNQvtCA+rcIu0Hw36L6JxpOqTvmMRowuUXtTPUNgS8b3z5/+MF75p/rAh
yVcB5UKhyRIZb0SPu9tnJsrFqdxALqibXK7E1+c5OC/I3wO3WL1zZVPMDQkf6Pai80/WiDCiPQPI
1lOcrXIuAw5ysD60Cd9bkzalumCYaoT43FKNJ7Aje/g1FFB5vFFzFnOedr0qUhqdR/c5xeiVY2cn
FFh+SHTE9R109TsGTTRQcDdkiVdPFUFOe72o1e7xTl5HlslQ8qy4PgvxqfdsxNfWbTsj7P7XKslx
kY7NpUAMvUlf359UllnVUJBABpJ4lfdN0u5uwhCfdQO8bd0U0//slRwXrbfvnLW8KHmNTFwda282
kZ7N2li9v45bFQtAhuDq1bxyGuEgcw4Z+YOfS4sFL2PSdwu48bStMDocKxArwz6h+BfIn49ZNYXf
eCkrWbIrMM7EgFE9W2CEWZdZPiCZrZKys3a85ZHwDKe0EnlpB15TQP3SZmedtr1suT3N8cbf6pKr
ZMy8xDFyQaDjiwVxl56M+De20bd0BikGLZJJOgNKCZRz9XNiQ3mrpIoMQGWzNhAzOMHYDmCfQmbk
XIa3fHzLCGGUrVVNNKHMvCt5Q2MJV6hnm4Ev8ncH7gg+qQFUAv/aFO7vTyGMlrTFW6+D0qZxdpc6
7SDugNfKXHPY6pl6Tjf0FrFIuUuKy+sYQxIwFFLnXQIv1yrAL6AKo5Lkz0x8Q2BwXowXjyNKvrRo
zE7xsgDhYylz/L21B64XUMP8Y/FaP7hRvsRVFaGzBpydYX1HC/v6nPeCTFMzLwRmjmmgl28iqMQT
9JSrPiqvEJt5Lg8EnRIaEtpd4+Y7RBXcDVJQkvwKmR911NKNERxYHQrlbhMtVrDf5l5nISBvH+JM
yQlJxJjB7Q32ZDVa6udM5r8gaeFwZ3s2SBx6gGw1V+JbOsIrk0nUB1FrxEyrlMYjXO4T+50vssxf
f/JU/iIH/zFYWtnCaiz7vpSVBJd9qJRcEv/AKsBz4TBnLJWp98VStz4i0iGdmkQAcqjmjsejwL1F
nHmi1YHwi2sHjeGr/ysfBuFmRHLxxPYVMy9z8RAgv4EMFn5JASWv+fXxGeMRJzV9bACjJJnjeeZP
HIVckGLOJCfB3NtmEeJc6z7lzMwBnYHjl0G5KdebkO7ZfDxpveTTp2dCj62w60cKTMdQ01GhATls
H8TeqB4ZhztPriiI6cLacZ8RgbhYThJfZ7XbJ81KwXvhWS+Sa6G/u0ALg/rKctUfpX5OWEtRoaYy
Qpzip7sknh96ww0jh2SjSWXOEfyDksDF+jssQ/j+NGte2NhCqGoKb4k5VLscHpxnXf7n3bWOL0M4
o7zuCquFjEvE2FGWRWpQXcqex7Xsze+stTqhjkrnTwY76B7nFGmpdexSvD5dghPFr2/SCrnuef/w
9a8gsnSRNbwg7tS/fwLNsSbqqufVoMS+X8jVyBodGCRh6bCO6j8Ph8j0D8u4bMmR3/yeqFbceGGc
MbCXeXPCk2pkqioa/pTnpVvx6yVWvTIKLFI5/sWCgATnP29E2Elj8qoncmzcSbcRPo6kpY66kXkL
GL2iZZ/rmCMr7GWaZyWG/Zwazi2FaFKKCce/DGYTuGAREE5j1xrZaFE19IRZCWFaQuCpikqxDRQ9
pu+HRG+pz9UcHBcWlswdoZCuPIbCM+PGnHzeXybK5JmyZVYCAcFwFnjn4XEfZWaZYfgXOhUfyDtc
c7HZ3wpfoagRoeGaFOTkk8tzlf8KjMOFZ9+p/HyKxJfIIfXkws4GCRH90eh9L0jvpOTZ0JFFpWBF
cML92wP/zElvmVGALq+gb0GOE2tzKqofiM4dJThkMp94OkEldkhZoE3glRWmf4hkunCmEtRNrars
h9vUi53ZO71xu5+zjXTuX2QPV2VpYgt3uTXR2/z7qC80MeBNsEsUSMTWKWyeZxXzVQW0U3vvz8U1
ARxOdZj6tJjjrYZLP2N+UwPMIGyjgmSifrBCPL8ylz+uzQQqIporwXK3FuuDGfvbqt8GgYWsEMtB
ukzgR2riOEO6lFGyS5IdO0PhhRrs6Q/JqQaubrFYgPxhbuy5CBX99uj9KZosYeyD6IVkk2/oGByp
93ijWopuUIHJ084pWBbhQLgg39GTvcwnAFPFYfctw28kjWnROsP8+PmugELYsO5zqIv+a6ypjGV8
RES2eyclNp6SCvRGghLAntKGHu2B1HulG5bt+LzQR2udRGFUq0WUralDbUpmIF345bv7uegVQaBV
w4/vZr5WGDdKiVMFVTrhuW7b6x0DpZaN76XRcW0Y6d2uQL4pVxda7IEuihsG6AeQIwHcCRJ+mcC3
eu6OkU7+JiPBc1ivUCgNMp26FJw2sPtav0dzmMtFys532Y0Ur3Gz39A/+VnmpggtkjqQTwF0p0rk
LAonTe+orvoTzjre44rPKwdJ7RwJTzQCmSZr6R2rjO9JdFKWXPyHCrjL3cwrDhstSJSenVdF2Xcp
oyJ4RK64ELfCMdMkaKzn/jw44dYxb4MAgeKPxZdH/5XnEvqzFGjReXkzRjWuBj3DB7LXSSyIudHU
NtkKUuJlLsZdL4PZJQu0lZ91RD5+q5FMGGRDpkZ7RONW6MK7qP0xO7uPGBKu1teKQV4voXCMLLaW
5VZZf9i2uTtw0FH90oL75oGOALRHXHh9J+2bx+pdfnbd8Z8LskCcXgQ8lfjJlf/ZYtFmS7Io6eMN
ILUxDQXHRhSxSp/B5lEQK0EsHHIcD526BjysXCAoKBdcESiUbG8C/1bgcgOlL4NUaGnIdHK6r6UQ
cFGtJ3wRDLq3e0I6/5Klc6QqcBhECnzn9m54R765dgG3AQ+L5eB8fr9/2gtwhosjRTp6rszoKN4w
E/C+pg+08r6AEfDy1K48gV+o98Y5jDDTfJcAordELanQq+2OU1XH4JXxt6U48KDi6pEuHJNHZEPO
uUph4zcLuzRjLcMBX4WibWYVMWpe8SlLAmEFvE9mS001wnWX9oIPvJjO4nEyZqP56hthAnXhbZXt
1VQp241nqcOSYwQmaKLdql+vtqnMChmJ9qfw9LPasADQ4swvSZ9lNvSseCzMTTer6IlKDO+rcYQJ
Hj92CuOliZGe3+zKqyGPZQxPB7XB3/gTqE9xqovqU5OPW0jI5JJhPFI+xjXrKtDh17Kmo5wVrXzh
Gw22yYgEK5bSZU2VBIgHyo8ANk4RyMJwMjq0QCwORrFCWnmoxzA1qz3TcmbcAGST5gswbMHYIYAk
fzsCu9xvlkjxTV4KiBo2W5drZZLzgxwiLOQU3mFWIVmKOUihMYRgQO3i+lRX/Dh+zbUuUbXwVi+g
waKB8unuTu2ULZTt+vJITizUD0xMAsCPcRCmVT2XGXU0M8nrVdteCLIMnInlFj29XWf/+k/VxpTm
RXo4t5tbwGO/oZUDqO/6lIxG3WLJDpb0cNsZQfkv187agmAhMmiCQ/Ksbm24Dr6wdQZRPPpl+wcJ
PXzRiOCRTVYZ+cr64YduE3SvtVev1DbquEwbycpV+vrIcBNOunw3Qb4NxFC4iISI1WUnNCeN4ASA
PpMVgMviTe3Nq1qzKeXLVIePD5qgJN6HhbtkW0xIWmuz9IHQxBWpewv14WikK0UG9pVl7fZhQ5Ub
TxFgfjiC1nFdZaP6RQny5wG4yomkYsICtQAnm3q6xkULYcpOhzwJ0bqXSDP7uNzMtr22jC6E5ft4
9DkvWmEs+N8I1a51zBOnMuXUsgctQJbKq5/A4JO3Xy8Cmcfa1+p6QN+jryOazyOs0DUPfIUTqvjq
Ze8EzB0iizJhPJBxnOx2qsSmrMgczeMB2D9ALXiO/b0HkciyanWvgHgRPhXQxymQo3Y2qNqOWmvW
GBlJBLRRcowx95nty63WhmGp0a7KeTj6uLtQB7RXcOXwRHnUVDtJV1VwXyUUJ1hLrYG1N4dudsSE
Jp5GQafoww+W9d6Kqi1jVUUl9n8l+LTiLpkaD917DLr+/VdGOnNPIoC3dEMped2z4uWmhdyTfm+o
7KtvOwrDo/rVudYjWmzg1G+NVNy0KlMG4eYw9A7Vblo6+dXNJcTuWrtdB+7Fohc9bgTWLBKMB5Kg
Vf267TIfKcSS+zlBTaCgoHtHigbsBZjcIHzrOt1LvFOtSuCBYWoqoy78Jbn8bm0fUqdh3bx1hX4y
jQKsj8VsMy6xjaDJxHmVZ2t0htWNWLAbL3Zo/YmCSkj/9pBMon8U24XbulU+V8cR1sfWQn0yEmy2
QwaYjAp3mXPqo7gNmtKqo95Dol+PpZGGYEVMYT3bapPuyMFQsD0Y2EgxwG1Jm2vy6GmB90GOogU9
SR2jkQyGyl3mjMTeVXtmeTsjXu11wSllLNvZ10Fuqwsd6MUgDLpeHdWSyCX5DfaULIGGKO7Elfym
bPr7Bqnu+DprkUWvALZFGDwAz5Gs/9srZy4ex0Ue/Np7mEl4DkqePlTjQCsN9HYzkqeV+GIFqqTN
x95AtYWq1DCxBTzHiYk/xAhJn8EA1ZTTtdHAdr64Oqnlz1Ie5d8oiSWXfuD0dADmIfcDE7UGcOMU
hqXxsKN8VK7ZKdZnKkCOBDePXCGI+SF4fFZ7qbj/uv3KDdGpFnOEidB4eliR8ObJLWD0tiV5XCtd
VC94xo2yReEs8Pi/6NLbu8yF/4TAihwwwYXxtHgmoC4+cz7DxUBaICBNnx/35MVJXtnFzDscjJ8O
CUOBC5WGO9vkPGy7VPLNRED8lMEqmcfbC/fx1slFO6hJdlsAiKD9fYjnvEz5zjqP7RJoeUhWn1jR
wrGG6CvOzX+rIBsokjZqdtMJpWk7B2Zh6GulwThGYQrrfZYuQMG3LzeWxJvE49hWpDhctskv+Dbf
gV/JrAgoFR7Z3hp6L/ufgfdmZ4iXbBNbz2bfzpGfh6YrLiu6ebT91GvHMYm7UZjrTNc0+H1Y2Pwm
/BlJkvC3J4cNfyrpFpUcdnWuFrdUG/AhwIXdjhUEXoRD8Wc+QndgAlcBzuTgZf/KCat+uUuLkR/k
K0aU3zDU6NXR3P49Q12nCtuShchdc5yDf4Lf6XokwlCIIwU9MjvIEof8WeFByo2ISTOq5KVr6wP7
5BwFxG8QNyLHJZBDzySto5MSvA92FxQQLUupPmDX9vDkeuSY0uNOIPO95U4G6I5iURTe07Z0foRk
Zs+04YuGGSVXu7nRRM3Jx/DM3BugJNfqrAfnnMfgpkddXGufV5rdfaNYA4O+jAfuX11gGv5v0lri
V7yr+P2luERCxdDGftAh6WfoSux0gsTYNlSPQFTg6IH3lWSgKrRbQTAU15wu2yCuWm/ymFRf+BTJ
5mQv0teSA+TDfjXwSCfMHsRSge/ycpo4kQUSj9TyRBaCnbQ9LEwxGRCMILTNEYzHunn/C4sfsgwm
U1aXnqo/KZog7uAPDTPsDjN8ETyKVy3/0FKIOZf0UIk+ahRyXuFFx83MGVlC572mTxxjhHSy3q0M
KPejCJyzMZGO5lM1IkWEc0lwWBTxjQqgZdreur+2xzclrHwwC5IEUJ2OZ5e4ZZMoNFtKmei6TQ8E
MXV7yLAqSA+ct+KLhI3utXEGnB/n8NhSBEIWHS1kemlKQ1qmlEy24r4+/J8ZvbErrlO31HWp6qFR
/AcxmGK0tOiKpOB0ePAcQsb3YvbXERb5v+yrLN105mWR4d9P8L7YTIhueBh1DYnYrwokyCHkeEbo
jQsp3HGv1UG0q8tYsZOMKW5tQL+YdJ/QUgN+gBsNki5Ze5BrJOA9dqS2scmu3uRtwWpz2FBg0pAb
90KGJInEWwcgD+z983HTsh20pGejKHU3RLOg+TNMVhfOn+lNd3yN2xEVJcpjfKRLo3byrbSn1GX6
1svAyxRO7HUekSwbca1kYYNWc5j5MlYJnouY13R0a0S+vcGTT5XRAizLryBPtZDzT3tuBKF9pGzH
M3+p4znxCx1xDp350jpMYpUaNGhZm6VuVvGPE+UC7yJGvNp/tyvPIKWMd5CONPHGprwpNLybVe8x
9spclfc129TMYK17NEEJ4TxMzhQLQAMvLBwibQrTx6Cz14QME3lbzzw6NtNKss52bdqoeipH4QYN
g5DsXLXaMmQl7NbHixsheWPfo0TAvcDAHVwLmoeKaqiDZv/gaa/TEXlpziknivAkVt8LsxdRAV4E
53EeOpLxz+VgQkkTcMbcUZp0J88tigSWq3kOkPQ8Llgf8CslWOadYjnXv0B/q66LXENHJKVQXDnv
yJk1fLmqMg+mUTOPvnyqsOBlewRSp3A1Gqet+vM/jupT8H6g9N6fDG2pbc39aQFfZQSHKo6bLnjK
5LDKZdYe7CXVRPxYu+wzJY9m3Sh5rXZlQdd0KqSOjdPsVU38P6ORx2VtpVmErmkdzoVF669VtOEu
sgVrIy+m8Jk2XXIyEQBvyJAgkkIygD5c1KyRssMGzvlKfAsbyOQKZfgE+fk6cegLyjRkHFjIbB5Q
lUs9I1Flwu8J8RTWHTrRuaaIcA0yOfpPuXTcNKogqvtyG9c6p2lrSc6kVyGwOaz1dH8OjGUhfW5G
7ufbHWaUqq8BcmrZzQkBH/KxLPhxYI0+J0bwnmXIBU9/vYr4Zoarb39fbtWpzJG1uurZjHLJJOIb
DIIerjlblSydk9deW0S0R6sOxgZk6ZI7s7qh8PJScDkgGXjTl5EcQYXduTzEzL/uY0MlgyW+fDCf
9COWcl2+vTq6jAceGuoeKp+Axd7nzCqF8NoonWAuaiYYSdmIEGaJn9fW80bmm/qKtjbPsVgbrYgW
gnwuBSxH91HupZF1+PJgUL1eFM8ZtJR0GQTzamdWP52sg6jJkoun6knbJBURcm2Zh2Dn7kOLSETK
0yVi/laBH08LSTY+klK/GKDnLKjGsnypuwojsx/2lydvM4F/G4ESDZA0zB/Clld3WChwlv46GEKH
uMP95O0CfrM8GVuIyhvNIqFM4AReBP52rZ0R87Tobfj+LPxnCFnUCGhvbwepE2UnFb/khCxDiQ7Z
E32Q5p3Kw18D6UgteJvdV0XjltM8PJFYEcVQG3bJEL+JyMC01lcdFagXPaBLV+qpSFzTfBR1FJ7Q
gRIm3kxKFlhVrTPSPFmVy9BB6FQub2yrwKI9c2b9Xa4q4KzIEhBMdHAKwF65ssEHoVbyyYHASO4K
f9WtHAe0I2LsYZ+eK90t1RhfuI9UfGhIP1NtVI89hGEe1tJLlp3c44MC3KxIIV1/8IPuzxXafsar
MVc4YCJVX1p7nAmlCqzrGtZqFqiYL+CaWJ1ZU9LAzDv2a00zl1vg4OsfD/czWJ3ON8T2c9iCkfzZ
EmKv2uSryOFFygtH5xh+1pb7bHXDeAj01c3w6holWXf3cZ9yjOI2Ta9SewmFf8IbruTeMGYIkAgj
c/mGyXUWLdA/Olskjb1LpTaoU1GGfvCwBmfVVmkoexdl1MecbhJTkxQZmaXhsPAMM7fpHKWsSBAR
MqJ/Vz4MSbmS4OLp9pGHpHMH/QoXaCfGCKNkKY4Ee467NuvHFTyw1KjhOHTkdJ+JLnfVHm/RMMKz
NnnCeqc8Ik60ECCuNceRxMKcow5me5AEyWAksy2yRYfrre75We8dsobB77yqbNqlArqxGBWuA9xo
P/gOf381KiPaPBjGWeH+Or0f6nRZ96GArAgI4SMBtG14b/kfK+RUBBd7Yg9gYba1oV6kHmjN8JCR
QN9Z/aTfACzlIGTv2efbRuARcurwc2utsz/1+VoHarPi9qKw1fOslztkHFtkFr+JRedrEZMfKQlz
ghGsJlCBee4V5nzkjgETIX84tU+YFctY1mt56uSmacgfzl2zchA/NzVms7fUI5f3NUSoZdiFs5iR
ULXlJogH1G7EIqO2+mt4DZlafXqOPxIOfGI1lyfx3rYhuRlw0iWUFjSJiU2yVvRr1IDw3jP+QtJq
VRGJwFgfYttGZjem+G8KOpScXCUsseU35EHbOb/hr9fMuMXA3EvZPZuAKZRbkyQ1iaTV1H/+qpE8
bP19MUd8aX/iKJ7gb2mcyLyexH+cT2URxAo5gUA0oNop+WF4cN19Uyc3z3rpRCWHWHHmi7JGYlHT
hQTlHKhk/d0YDbkAqFUlmg6k3w4+NiEA1wXWn/ezADu8ig0G/skX2p7kyHocnCKL/ABNBL4wZbkG
CtOecHr3u51heLkmfcEx6owrx189QherEsj1tznjtKRXH28ndEEj827AIvIheFLRPUjxAl8ge9U8
pDoMKlsIUf1A2mNOmK/qzXCjWBFw/MCURgqQt5kXf0KCfQhtjmtxjzqrjM4KeokYRRkKbyvFWkoq
zqui5acLVzfKqJylHX8dB5rX3z0UPwAo5Ak5xVvKUqIuXi5TQiEBsT8gJnH5D0Vnknf3iH0VTqxY
zCD75heiKIv2ixrALPS2UHNYB3nx6MGUX7NXeexr399OVTDH/a3a+pbUCrN4nWQsjNepuHPoWX1U
oKTOQdsTgSlnQniK4Kz4yPxCxxLga6oRr5G0N43qx2nj4PyrL5wjwzNgh1JYV6HIrEapNSvd6Doa
qndwv93NtXEYLTktcPokaiuO3Ttu1NMWGvPj8jlW2qlXQjoxzVOJCqqCiUYcgFUPpmvNDkFCW/DJ
fczYW4Cs0Myx+BTi6rEqfT280uhoFX8pDzrQexdRM/tzmCxSmwK2pdIf7spVWHs8garCd4TNJI8B
jeOA+qClzZhTFT10yHS0c+MTpwez1bhR2IH6Tv281zgGxaPCcRwuZGdnNGM4OntwIkalTUAOMJZd
/d85fo2EvwaSWAjnfIsuBfvmQ2Q0pQfMtt/Gxlxrq7ebq7+LrAG+M1tlVlI59DRJH4VH2d3CLi79
PVL9y+RNw+vNRbOIKro6B/zZbQEx+SHtgnlBFCvx2meiRo4+Vqw8yqDrB4yN4x+UrBy50htqaIAZ
G0ocbJtA6pHBslFOxWcc2MN0HVdk6tQQxfuJ1x47Gnqba6vILc1bx5V0y7Y1y5nqAs4HM+SkNVHh
kzhXSkmP2CRJ2FFG8Cxv8Y3+3kEsXAPJgltv+BA/30LqNh8ctLDCbSGGjOLjLSus011zLkHVHgi0
5qks/Kc5PylEQB/0/NCGKwnIrtVYoLKgu4OXqE9QqCUtpBrqr2M1i+Y9iwU3LXon1js9vBFcUS/B
YrVOx5cR2mVf9GnfOTm09HrNEAdihu/wuAdLgNTUSuU2h9Wdg8XsHgv12fZWB6z0RyiV2NZ0i/7p
Bwy5Af0wzuodCYM3V2bbceLqR4dxPuryulfETWZMWXPe/yhPbYBekjtUfUSiWJrMgu3CB71IbzQs
SEYJCr/OnHp8LVSfv+GMx/vuAaCdxL5m5GIITzEdIa+kX6wJxY4aYP3+kzmFrQfxoUjH/f7v4baH
YTdHOU3xG3N/1bEqMd5T3LhZb14fU3PSQZUZK+GHqMzXpN/+IiQGMQHVR6A/jeU85xjI6LK2XzFq
yHOMV/DbEercBA9xP+ffyF5w8ExXjhoP+oMvORrI6zRU2+0/496hUqgH+P2mCAdmpovI5XbmhICi
QOEFge32jfIGEbAvBGrL22QVjSzz+VcFlvvlJ7yGpMw3NXF6AJDG/uq2l/yuk35UhxxNe14MbVP3
1wocO05KiBiIBUrl90vHyxzdsa5+yhmIdAgu0o3jbt1cIWN+6isng8HFViXgWAmZtovPuq2d57Gt
Agja9wziahVXBSzAYP5BwykYlu60++w4nSVBvZsDG0eRSpFBKObZUHsIRiSQcB+Vf+MKbSS4yFmL
Nui4pBq17vNTqMSq7knewQJHL1iQHFdMMyT6+xhvxnfzfTU/DB8yoCuf5ARICch0yUgcSt0p9ZuS
s5MH2pnp5MmBm+dpSYa6ri67lEWvTC+1q421Uo6znN5pBMGUcurjjbBrLIFgIzVEIsgJTzdub4PP
ZC2hUJaE73I3p9cCmfMxNH0WvhlQAO90WIJW5uyT64v/Y2p7/dB+iCybuXo+Ng415d3w7rrC7zpG
Cj4U6+l3qrTWg1dk08YJEX7C3EUmmU8Z6ZbNyL42Iu5suLSRy85pAdcZFbpo0S44SzNdwCa3GnPh
oGnQBl2yv1ycpS5Lqu7f1h12NSTOYBDU2qrr2W0pRWo12jSi3RIwR0Z95oy81sINTCPUH74awFcA
aHzrt8JtnOSsms16PjTXU98YDMrHgrnNPcqfbBzM+lyVQoCZpR9ANZQr+wCvRK2X4zJ7VD6TjtLS
RTHhmiwycezXdwT6azayJYhmOBjPmY3FVps4nV/8knVDUcwKLTIeFyNUKKszJnOKMFgo7y0wO2OW
k25e6Lc6HwWNdVD96yAZ/5PP7QXM5H5OS2F5CSB0IhCL5B5h9RnEAsj6VeE5+3iQCZRURn2NQjkm
YlfkC7xaD9I56Lb/pDAwyRaruHyXRTu/1aihAFiUyqwnzSTs58gGNCfVmEihzfsi/tS3qwgZ9CqG
BNdWo5ryHLyoy04dI3ZTdFmjOYTLKh5fq6Yki1U73ZNaNtuC+rOOAvwvpLEeQp8cG7gJqgatO/AP
vOqdmnYAohCWIEVo3+TFepCdmBZWM02zSgV1UrpRVbGVt20xIo5nxyV0BCeZAucuWR2+Z9a70wlk
nyT1g4aRGWgPLwTmE0OcE5wYqB3dc/WUWLklMb+hqCMDLYty2eBtnIfsW1PU0DITZsAG3DaiX2dV
XZdlvBCIV5UDY2fdOZCvP/CleuJ2cLKXv0pNJzTp4Q6MqsfYwVKAAG+lhVKehAefQGrwLPkQ0K2X
diZDllxyfZLADEAmkJkmaVJ/7WbEw+Lu392w/Qb5P6HBi51rh0yjD6PmijO5NjLXrNp/zoAda9mh
PbmqHub+8PF/mNsTJYYuc58zPvJ/HC3cn1bzZ1HSdmetZWzsr9W8fY5YgY+SXkfY42sCejFOdMYM
HlAU77Loj+w+9GlXpisihEGt5E5vSrRpeLPHgCZ1bbYgD3mCjw0e703cpc9WFfqvNcsdwwMk/Y8x
By95gf+ej2xrrMcr7cOyqyB3NGHID11JWKiGRTpTied880QLlB5iAwNB+waPq813dbrboa3Z7JfT
NmCznEwzKN3yR02MJpYghyyDl4EM9GPZKSwuyUUd/pS13Ja4cVFHjAw47wwPoIw+RCvsw1pxSUxw
nKjJ9rKSTqa774qbY6zzwyxXNibma4Edp524VY/1SzFL2PrW5dLN0pKr2gMArVhca/sFe2Ml2Vgn
4PL6qEXbCsQBsRapF1nlrcbkeory4bpTTtm5+yV1HVN7eisVun/rPoAXyFlZ3qnt8YlVZt1MU4Sb
EM8Q+/7P6RqLOdorGLUXhQ2jOay14koLVXHafmKRyzGTTRECXRw6S+Bz5kvqCMM+uvgQa0QIfEMi
zBMyuEnFm74uuvgl0BLNr930gogGAPkztZoTeG9RXyHLnQ0lB6ZCdRMRQx+Gzyq78zlXLOIPnZn/
sOBxp/lqa8LWTMYeB6w9o7y726EJi2dfRgTwCPnZcXA0V44yMXt0YdLA3/GwZ2P62xI5TnN8G4Zu
14YD2231EEFGEVTxi487HKnEytojNjh1Bhhe8jUQqhGUFgdukR4l84TdHyT31O5SZ4hy23MIZWfO
lkaZ6gqHksNkS3FPN7srcaG5nvOOoRrfCAQH2D6zR40ytBZH8rEpgS0fQegmuuIPyR2jSdpNWmRv
8GXEIGdUhqxE6AEvQW52hwaC5tY5ldWl3rrI+iA0H88TL3mHXO5ftWcCelC8M2ppyL2UHm9YJtpz
xB3jHGMGplhSKOw1tIgGlIROqxxq2/X+lq/COl9UqEh7uOGZrjZaNwDbiWZ8K4yJLXsHcwMu3OPA
UMMjapOqSi7ik3WkxAiHEGunpmiiOvo2J1+biO4PBCymOudU1b6jTKRkYtVComq/aiERXn/HfPq9
1pAqny8EQMgAqVYlfqxsy7l0+T+yZq7Bmjn/Whz/OLk27GBjTF+kpesA82ahDEjIdoFVF8qMoU4r
/YBCUo422kYNbny6+qQD3/TMqWTd0XiP0UZdnPLbh8zx3NffXhWyeICSPwH7Fh1Gp3WtgRRjdl1m
dVrEghIHwDushS4pMLMCIo45+P8JSt7CCOLuTXuTlRh0UoH4Utp1qDH10J5G1IyWLTnrLekfjOjo
HI+QMzBIeimbQwoVzh4g16BXOs4T4BHrCwxco7qtMkRg/O5T/PvUX2CVgef+CI3MeFWwRZ5v/MmE
VtgeshODpW18ZRwEJjyNdGZKiIJ1XyRfMz2xBIeoa8OoruBtlyaBJhZA5Ce1vgmVfoxUMkjGSo5f
vXY1k2hO+6dJ/qJam2t/6ihUelKguEAR2HDXDBv4NTAZsVrs1TRPCBDwEIsWbrsxAeoYXEqvynlG
mGsoRpu78ZDTLGF6NR2tIV+nVy+/fxFxv76wdG+BO31Z413nZswWfSg9mqmIuPB9NJRAulBx0/W5
uzKv/IiSTAqbdeELdEA/XZTCl7Bjb6TD80+SFKOMtXePyhZ6lngXc5YHgpw4IOCPgK1V/Wv2MZCX
SsmsCZzbZhHAV3ESHIVUJcrAOcEYwugmb6FN/1OPeySNcWL0XemVLzvyEzVcs0xeKPSlOqdlvP78
Rwk1xrPet+x1kkIffuzRW5bCD42HuIwjBQxF2RczfNX/i6rusvtFr9+GMEix7ww8/ALZCUROfI79
Akhr6AtFgS4haX8Ax3rgdOgeqhFij7C38jlXHkkZ9wc+20TwEq87HTx0vKUw0YLe20JOYjCK7aC/
LwMu6n1VttxxoB94np/SsmzFcQaWrhFDh9YDb7tevhEmdIKsV0F2j30nwK1Kl26NljY7KBX8v9H0
t0mrT5AUT6UYx2Mql6mUygWtynSltFgj87QefhorD3kPy72qUab/K79F4/k4GVjYe55a75PykKrq
jRw6P3K19LiCJsbIslcXzB8cqF6gohxZsxjZd+JNErSjTqaC4tp2m8v7ZudzK+HhPryvTL8btgJL
3TwNqqe2D3c8YaJC9ImQOJ5U+v2SaFVTpu9xAKR6YGlJ3Gr0HEG0vLVSF9bQVVLBO3YulKJur0og
ZwmdHvQckeIPBXy1iAby57qc9BKL/MUkvsYYATHCxa+HmXQQfINCoO0xOC2RWZ2CPADCG74KluLo
w4sbZ2H6WPQO4fW8QojeGX9bXy0Cv7BctdUm4AkRarNIzpw4bL1BxH7SBIad20WSVQDh6D4mu4vd
hGAar2WaD1z1U8PTwVLWgeZvJN4/psqu5f3SuusLszxkUkHXhh85p++H5lqbMiD92xWenZLlnAOv
XAt/8MgRg9j9AzlXTPeWRBaorqrSubKBtB1hTBT6lsgceNQHKE5dzOz5m/x7YhuOtzErYN2QyUzn
n+VvjDtmhGRHZILbjOAB1X/Pu5MjQqlsjtz/hbv8XoawnAc9y9hkU60Y2fTSjD9gokApm43RFF0W
+bDodDBpCtq/6OWakJEAlz6aJRTOTRCNjfeKJ2udJFpYY+uBZEbU/1uGygHe9lv+cizVakU/vTY6
jeRa7rbb6huUFirWngzYedyUtlXz+rBQScByzXnh4gDFuCj+tW+ndVXMD33Q4rMD3cW2wNEzNEB6
ktlKgbdrj7I6hjKF8vf5IyUVkM95F998/hF4zi8LDZb36IzB2EjKg/d+rE7cYOIsrqaOtVlZCb6q
6PH7Fn9TsRixZkxq3pk8oKRipyOr+RdQVgbl9/rQ7CJOFM2TQdTCbZD+KuQ2cyXPZijwfCO/RSTG
b4sY2aO4DyyBVScCwlEf/YFbT1XrPAMIHqs9X94P70hXdQyYPJlPk7PfphY2q9vrGzaQFwKzaLuX
v/c15JmaFN6IQ3GmK4JiTXtLSwI0mqc+jgUK3oniq9UJez4Y4XRmdAYfUtRRYw7uZwT4+5yotb/J
h8u4iSUCob1Q+76mvS4a0YScacNFwmPhjTFjoRfdnl/FDm5hUADmYLf9m6EMc8vn7YlHXLX54+ES
OBfB5eNOAKnscZ2kdRYjHTHCVCwo3yb3h1oLhkRFvU9cvC377N0lpwhJj5bKk4hpEmh54KFTx1zu
rFOaH8WZjCH8qEhDvCKLdYptolPQJSmFcvz3OvuUqJY3e0SF8Yz53X73GaXbO+SJWMMmJIbfCwwa
EfkLXk/yI39DRppSusEcLmBEWrRwabllOg9/TgovuUfbO96Gozjhl8LVDc0rywo16WdW54Ai/EhY
81en0Q92JHG8sCNw6IPgeFy+u6w0m8Sc/haEZ5tnuafMIqF76WrHN+1ViPZ0USwc2FR6vkF2ftIR
mxE99J7J1EYlg++2q8WcEJzRspoKsLNvxc+6jWfOy75Pld6EzqjeCSj/f1Hw9mYmu9T2GnllTrKi
okDyBZcyopc2nFBGsAHDg0x0A/JY0DjzAU7W6WSxdRt8YRmtGmBaBjB/0sbvXcVvf+/ndEzVBaqZ
FQo5FCPuISO/ulkCDwgOAz5DMJkJvM2mwWPaSXfqgDtAhKZuu5Y6amVnxKWUxlKjRzfDsq9uUxmF
EflKNAqAJeV/7QbZQNBW05RBGjy/vJnXZOBmsWVnhORDNQgoUES30DriBkOm0qx6CAelzDGCKTUa
TPK7C/cBzDM38pfHf5mmWTyzQpxoY5rbzfTH4GDbJCxSvVhk6QpjYBlVsXafnWfWaEKcE48BGjWf
LdhNtEa0f8329ebH4g/UUlQ6c01zLfdgHD1spDv72r12Fq2zM1K+kZLEB5g/05Oh/SgukcMamZI4
UO3Cg4jiUFWLXKBs5OQv/biWNeC2AbBBPo1ldTPgzesAWUKrLQaVzsAag+g6Uvl2MyUniUryyI5m
fd4t6Gft5tlvcNmVB+D3FzL6tIZz3aZluKmdxAafYHCUUtZup88bIc0sYxyjVrd8C4n5jcoDYiaV
aPePRYF0+ycF3TZiJ/0lynqjR6KoCwWHbEYgRRLr40zgz/ExEaqUvRlnEeuiwmDKuYeqU5PgcyZK
kBlvjix/7+3r1MoXNF5fzpd6V+vxUnUlE3XKeVrRhyQxTEsgCsJPnhqBYHNoO3zZwMXletOD9tlP
pxAxQ4JZj0lDZVQiZWpXYqPfj1iGo29/WPKVRylftWWnBp8eAFmuBCrs6CE9v0ZC59Bs8Ytirk+Q
1weyzjCy3u7begoPpCzWQOUifryBERwLBrjscWDIzaLcLYa+KpuAV21oCSk2vTYwr1dYWcVNsCZc
ZjBXK5qX1dFA8jqLSWzNmIyhtBssa7vBUx5sItRbsC5okk4sINlsDohM4fNkUxogR+VfzyhyreyK
OFNvVl+NlhohzvSRzp2c3nDfuOj9fcfHZMH4BQi8wna94pR3XNkx8wKzbtA711f6DYD22tg28vzn
aFSnqPhWUgTALRu1LYrP3vBUBV5E+mwDHLutwJnMiOnrnUxvMFNSkCJ82CRyb7j4+ywXuSTMTGZz
P0vfoTbVnsfZdI2VjXoojm486yQvTbNSiKz7YRvy6gIKG8eYZqAJoA9lz+n4vDgjzwTzWpcHyMB2
iVi4DmppjWsFKYIuyJnMT6xGWuNHEGIandVOXprkUGFwxdMXQXLyB+WCNy9EuM85DgCJoj70wxgM
17x0RcrOyC53P9qkh8jeShV9vTHZXshnp4rTI+UX6M3/HA8lqlnl4rFTOgz02RarIrJswtw3CqQR
FgiqjvPMwCIBH8DpIlUwe7DIibrgcg/8vsJzT4s9gtoFX6jFmALWaHKjGmdWHA2TdFMjsV0nzMFZ
D3LlzwjJzThSCuxzY6FcBr6hJX9VI+sbQpZwEh0SaKwsjzeFzMp2srGQH/pk8y08Elxnrw1f6rpm
+C7/oP1kLY/OBsBNybq0p9AfmxEXOBGq0HOBlaDxpXL+EijX5Y8jPbBHUkbBQFQdhOgIMaX+1Fdk
4tFcz5HWmtJi2CrkjG+TE+DA6dqs08WZeq+XNUaj010OH7WNaysZUrbjNukgS8VboGwadv74pxRb
+Xjiv1HsyWmtCroI6xBDyo4e0QPCGKOKK+nx+hl/YnMP0JQPIbAKRXzdNCJqk7rzG/wvMiYfTuV4
Gw5Ni6YF4oVH+nTuia0kI5uGS9u168RFYB2TCGqPSpUiL3OJpRB5BRJ2wIigdTgSSkNO0EzoW0jI
JYjcvLF/a4j+HA5VerPJtVSufxcKDHfb7KCZy+pCV84n6MkY3hMaD68RenoO/FMEns4BYyz1rPKe
1TGCatpsIhMf/VcOvecpVEAF8rL3x4u+FHw9BXcv9M2saq3X0qWAla3xUVYFj7Otr/N39swKRr7v
nT3LyvUmWXrqa1CxUYz2/SjwAwKeBoFI0xUZAwXy3nmgOZD0o4pDQZ32vkt3jYEwubPtVp5w9/Vx
jm2/+q8bKN2zq1vN818m3m5h0gzvhacmm9c7SUMERXHTGCQDInGxD14uS5MWxygubJs0YDTXCHv6
gbYGVlDUHwR/fw8vP/JNDOXJ3US/gOTogI8NU68ELTgTmnW4oRVtHFbhEY/82azp7PR8t1o/VWon
uANxEuk1TBNhHbgqz7WlLTY+Cd9IJzXfiqFIsAU1GMMCfWtiL0NVf9+wo1Po/5iXw0vfLOkF+M9/
Q0wFVHtSBjrBedsg8p20udChKaXtIimzR/954WMS6NsCgumtSBHJ0j34jgCiKmyKVJMoS0KGefXq
BnbpyePxz74hge1GeC6bcKMrAjFIsex5C2aSwTDcRW4JKv5gNZgnqAD9jQQmL/h/QQG0VZfIXOcx
zhS43i2hRn2DNxxSOvJXzpleSci50Ssq6yIbqasBstCa+DZP3xbs6XmdBXXq437f2Bzsyni6y3Oz
0u8WI+p/eVhHY+MOhI30jPqrcRFc2+iFl91bX1sJAkdSJ9KiI+tuQzfRT/YLcWa5vBCsCpRUdGks
RSpEqqPI4MbLLp98lo/3Qg7nKzmFtP8Gpzf1Zj9HT8PXRMvYh1UNcR9avdtFM5EPtNABBEfkZ0uh
rJDXvjGc0HcUvGknj9G08hqi1AFBAt8hNM11yzjwRfzwlgkUGNk9fQ7FTHo4lRwEf0Sp6bMySQ9t
IkxXyIGxvbrnBWbP6c4OSEUwUGgL2HuOTEDIiyta/S10oPvbs6X3UKb7m20ECEF+8+QnYisXM0XC
NpKNn5ae+iAWbr1W8cKhfC7ImdqUsyM8FpmXHZjnae0b6K/7dnvSwvrVC3/8NL68/oG5fLMuxH3o
q0y73ZMxOy+WBKbvA+3otvwqlHc3l9/7s13kFIfOmHshp33jqMM2QNunc72m5QkvAnTAeMoBTTAR
2r9t9ME2HU32E56bMnIQ/XALcMhKsSu2/V320GfWp5v+x/lJfsrxasBgNC3+SDquSN7SNsVsvXtL
a3e/rmNm4cwqPuP1+ORLRNDLoVDJksU4w8phVTUH0+PVJKaDJQU56cNu3r9HZ6Tvulk/gyRx6q0G
o9cG3s1vwz3XAwQQui8IaGS5Zt/PNr3fAt5DkmQcEgAvPq7eUZpPdTFtLHhHJAyd830x/kprC4Lt
i10RORP0jUS0s+y8y0+NEPds0UgraJHwHDDHWdZbFS2sidqwfZutl7i0ZoOySevRANQDeVTrxx75
jilWrCgexHXGSYhiEDuq8EUnFVK8I0RSPPm5q1UlH1K9mskFxbKh4m6/phf5fb95DvuBedZp2HrR
soHNhzPulYkWpRKefLqUKTRPMpPHlFC4VbBb2NczRqTnnS6YBhPqDqg+4lFtW9u2d3O0yKhOZ4WP
ZF9B2m+tqshrnNCIzjB7vgUfRxs3my52/FBworsra18A3bruZoit0NbAJ9C82mWXKwPfuSblb5nb
Jc710XYpcrp3mkC+JGfrVPz6aOwt+mi+2hJys+91jtgzVPveLB1raPWZbTO2aijRY8BrOdTvFGJM
dznTLL6e9mD3dfDmXbKW4csyAlt9aRxnllsRUjgNBvln7NEUiQzh8c3+0oSlUoo78zezJrJMmWpP
UqaQxcc4y9cXPlqJvGeeUHEMzeF4fnLg/t4hxIHEoSc8TtizoGSITmDU+jXXWdb4nzTlzhUf3SEp
yOX5X4CW0DdiXn15PTzour5LQubtzMh/QDt75BmMoZG8yTyQOe/hnag4+oWs/xPC7hCoxl2qXszt
QGnz8m23Kpg7lDPojUrhqagWaU4O0WvhLQ8lDEw++a4CTUTkvhtUMS4GdZ1J7DNCRc0ANdGtW/iH
mRJgxyZg0RZdVBkjd4HPf69zLu1u3rjkpigDw8VCmsLitV223BsZvsKpFjve4uZimdXonerlWZGD
eA5uG3OlLy5opPDWQGmr2OFF6632Pp/i+gN5IGMhWPnWwOiqlO1q0tR+wocmQnH8JvRKE6Xe1WXf
/7Iw5TCUwakkysZenbTs1MYUyE/Fn0XqurlTA66xUoJtsfTHVs3VE96DzIuRmR2l1F3LcRXy/ppX
CPUM1eLbSQoHjs02qB3NoRmpNP1rF10lmyTDfDe4EU7G9BtrdByYrTTM47lJsn/GDDIlmS7Xym4n
3lUCNG+1CCN69WpVNTfFGla6uBGd0rI62p2dbpt9JYwLmJuJcQKqipYpjaxVdAaIWmlwH5c7daqI
XauDFJ6zM52ic9WZAg0dpxfs6iUY+8/kE0a+ICSeVLXb7U616n2PUYSPa7hQpo5tbVHr2BohQZZW
Xkpi+wA9v+RC7y3G8C08BPCR3DvYXb/JWsI/EPGclPqaY8K6lr/AqDfMkLYfX8FuUiBKytWfiHIp
cIaiPvY+9ClTq4zbKuU5RsUTHNAcwhdVrxAf0J0AIhZ7cMp9ol3rPR6qQFH2cC5aMRLiZZ4xv8CJ
nlYvlybPjOBgci4vlqecmgqZ16sMuc+aLOxVcTUKhuQkDpLlWOOXHJ4Bz4rdGLdqQWB2nGm9YBFB
37ErG2xmisl09+7jx2ng8YzyoMxw3q/N98y5pPE8StXCtZFKcXhmzNRCz13To0HtM1XBvYuqRgI2
ApMBywWTi7NXIHhgWo2Z8JbMbOs9aa1CnfakvcOAA6qtsvgK4WHHlRfINLXDS8VDmOGxWFUsLVub
2aBUsN6efS5BdQhY0OtNmVtCZLMyWH6PylPX/6WibmrGkLKYuRbI2sWokIqtcaA2Xx1z7ERA0ePj
umIjWxguhb+yJbLP/JxXFc8XyUjXbLV0yr1dHKdtquIO8u1jFR2+bNBBECVymk6g4mhWQAhJfpun
uLAQRX2js1GXfRjbSQ4/aebb+U5+Cro/5FH9b8ouhZSoqVD7n4tf2rnRIpgl0zWXTlZxz4wlXxqX
SRfvA46Ng7PQt5V8/f9SezuW2KzHmnOnF8OwsRb4rYpsihCxISlLrkIuGyy6GegTnu9NocnJlONN
8v8mrBWwqPYYaqw+7O5pu7YbUiE9egXOrTvaN/646vsVE61jTVO7FLR2djHZO9zDgkA+/CnUE8sK
mqNytldMU6KqFsq9T+C1Q0NS7RatcrmIHzoF+1veFzvVL0DdbAxxtUr3P6v0khK1oSLWEQq2zuel
hGPdvrpJ7R1mrbuL2BSNlU0Is72pbZe7L8gORTO1vnkmcYpdGrSPEt2rDJsZDlImM8116+DKI0sr
suLfx3wBbqYak3GyES0DJOmLjBOcp4Qk7dBPYZmiS0W0xERzcBg3IpjjEAa9y8dXuclrvGPdRYi/
JOOyz5PDnRCMNVBKSmddyK4X+YfAvFiiSpdmaHGbO8NTS06OOkPoGx75ZZISQxKC0FAsVpvJXAiO
qd2/COaxpGaIwx6wumwG4D4KffAK5+XRKC5S3EBiRFqq3V2UVm5/fEg01ua2UL14M4w6xrOjblPK
frBriANQV2v/o1gGYjbr9qUjzhjkNPuyKFBozBXs6dUEL0txGbez/1STD/5K5dIQ/QYqiNbJam/8
226IdT+fPuME2x/iks1mYOqj9FVRZFbyIuJyXDqvkSFx2y6Gx2FcgA9JsawHqQdm859gQaaMqT3j
hVpiIyFuEGksI1uGIEioTLB9j3Zi7EM+fVr5kz2ONOoW4c4zRaV/55hDIkbyuH9mdVEGROgDTnNI
UWBPzJ5bOpyqfj3EniyeJWz5NndObSe/9sqkn0IzAdLW3ewrSAIHqc0Me4vdXAMaTsuvHWuKkZ1g
RO0NSEVh8d9RdFEAmjCzKJspNOH84FCYu5EH9D01XEFr7EJOCdtWNqJtED07YLL2hvbzLP1k+4ae
7MnodXE2WgrOKm4F6NTR7d1v8CICtpV9DEWVDi8KeN/owKtggAVV134qQqI0o36WzW+aLdWUFVYi
Pb1+lcB76PI/oBseDlKyUNBMDGpP0oM2dIXUIk7or/U6fLI9voim1j+jKbph2EwE6MkcCGe+9vrS
FmMnAuHuKcnywRQwPUMt3w9hUve8yir8XSod/EWDjkDzk/WRpmmfGfU+GLO7O6FiZtm0g3Q3Mn2J
c1MGYZPPjDQ/xX5XisszQmm0rHuZzReCZb6QDxvDMwyysavRjBXdSDwIVN2JLy1Ii0qJgy6rnX0h
rxVQFvEgVJa2PwSxn/IRVLIOMxAKcDvRE5h6LH7F9Nm+DgTGLm5VSEIIvQZCnxpdt3YPZWC9XMbS
H/MKkgk4XjYGql5Ha1BMTz060btn4/cCvTEbm8aPzfhsn1Aup1sDAnldyxnEIMCQRcVGQnNTjQM3
S1n1lCVNl33zyyfuNd5zADlhuZ6ohiJgeuQA/VR/pMX6KrAjlA6Z1jhzzXX2msa5YVW8/9LnBOd5
SROdQ5bFUm0WrDM354g4VkI3rn5ZP+ZADEKUIX5An5maHlEvzHQ8LduXYVRWwmX9pR9RasOmcyCT
rQw1SikXi14S86Rp0Y+UCKmoiYwGY+tNZjyMt83DC4DubWdqgAswkChxLRO3Q1Y3kKDKbMukMKWZ
wOQl3Qx+dGRXsZBk14zglC7gBOe7ufeholc+W+MGaxElM0X1MT0uJh98QOkP/w94U6sraf333ULh
OG0E5ttU5JsUG30KckUe4F/sSFGalm8NxeWZCQRSEYhJ3MKFM01J5peGup5tKuutIx6+LqgFobby
GRWzmqpTcH5J05OykcYWS0iJVUOfLsaGiEaLoq9DhGI6tq5xHRlUUGOtO6AnQugQRccQUk/hnD3j
QSKeuYP0dk+qsBCnR7yruFWvaLuWYtgxlgDv/7v9vDZuGt4TKYSJygBCoyLDl6ERjmkjJGa7IIza
7sfHVJHGujhGcuKLaAQ60wvd+jNjQ/9/TqJeqjSG5t1jsmyIlvfEM12umTmU1FyCkh1JX5Xtl/3M
OnBzrHHxzD1tY1nGXF3u01nJuVxglfdXWHiBbtNF/skNDmBhx+oRNgDKnS1/E6NssjZYj5xYeOP5
3TwplaE0OyziqnXLyBoNt+Hbjy0xRLHda2E0FYJ8X4InItambKQweqr3M/DgrVCfcJ+tsd1UlQI+
4oQ3aLXbzQZLhSa7GGO2rxXZRhZefxM6UHuebWR926R4Wi/PK0KSv6bx/URTjb0VSQulGVOP5VkW
nyV6Q2oEUdqxsN29Bf8SfLSGehgbTFzdwh7fGm7IbRd95JypqsjqVddehoqZZGC2gYlXOvXHnx3k
PrKo1xwZ/XQfrJqi9RrTdfEcNJAhC1yLLyLfIhg8ssmmmatScSujTAD/EIaLQ5fBCLPZRoDK8rDm
19EmEaiw/oiT5qJeMHRhBbmh6xJgpeNv58s9TIvfQzimhSCWk0L1fskHStcBG7P2lmSFOp13Reob
ZolgKSgmF9yUPCJyt4Sf1e2URGvPEfa3W8shyXRHZ25f6Zmua+E7p8/M0bkDoQHCPl3mAb815+sW
oqdZd/CvdsdUiWIeSS8ROfacmfL47bNfKbN9HdeR+r8TgnudgJqIl41oE4u7jAZOYy5wOMzx4Q0K
+aqfdHEP7+bS/6YfeQc0qf89REAsJttYzyQVZxLvVXfZnbEMExELlHrLU7AtwBeqRMnRfn9re/jG
ei89BS5cpRINp0Fxrgxa/DuieoBXRSvTAfIRKCLFUglopH/VL0ONmJLPymE74OMqucRfCIqw1t1L
msaTCw/E8UMGVQvigRkthgjL0GB9io5hHj2vWpE6s/sISTrloku0uijjq7fTXWMJyGz6B6ag9Zyk
iI2x9tSB5KAltRpiVhuL2AfkRTg+jsUlvd7mxBKDCjf/8+mNAvyVEzAqVbgLU/WiHrkOuPgTxu+p
xTeUzlF6xTxh3ROszPmc0WAyJubDMrNh8/rAhx4y3C7zKbfh8OAlDopLmNXkKJ7CprJwfqQ+3aXt
C5qsb3DygYwfa72ObMYvjyf20XMt/GOV7rFenSEABxsgO9CwmxKepETdG7MInadRj+MBB/PKzcll
YP49/TRIU9f0hoZagbj6gzYlbOBlXQVBzBlI3JygptrEoCYVwa+VXx+v/do3BOnlI/eB7I0kF6Ny
LAQvEG0th75r+v26oqdFXZmZR1zefrxqUpnGG0tsy4w73vDYwKlHDW74jprFGbcdkczWj6B1aXZc
DZRSxc3mZ1WzSo75AAGuQiezpxz2V84E/SIic/RPJKyfxJdKJbsaW3dqaG/tMkvxTAqNjJYvI6ad
RWDl5eSqwjwjPMYgLEDmfhyc1GI90H0v4BgVwam00cjitTanxfKeTXg1DLhdhuHP3TBDS5pBbaCn
lRqKPnXKuyOOniXLBEUp2mxpMKxNHO8OHp8/DF6zBmrYarzV+7D9cfL4XQTfx9HB8P+6NgOCcUs+
1RCpW7FlKEmAYHdC4rS7JHSqOfzj93jPHTFXA9xQe4z5J/+GPe34i9AJ05To/BDNJn5GXLJkHZs3
EWH3rnL+2Zon4rZu1PmdTzPVtRxO1QJQHGdpPGepBtS/Oso+vv4ROQVql+HXhhAuCtENVQxuGkun
6qaAJPW5c+mZgDjQqBW83Ym+IVj6uwt1m1fR2BHwfUTFR/FngD2938VL4yERpHupfifrkMz3VDdc
PIQR/amZjE03Wp1SzmVU0iu8ZHOSEpi2tLyMSBjsQd31QzRFWT253wsZEJggYfnDmGPGyV6dUPMj
iOICijnZcZIKul8aq7EzK+fZaadkf7cANU2eGFGPppImWfAld57pRVg7LTRvGy4bX+N8QvjoOJt0
LDQSO16NRAR8xU6CWnTNDTDN26uPqk8Xwnibh00Xl7BTNCpNhDB+8nCMhhZTdXpWKdPg0HkMcKaM
uBK4L+/WGcaCBi0nq628Tzk6Sz6Gwl9ikFkx4nI+hZwjz0+RRFnoSzQ7yxIKiyzEGqqFzQdA8SgX
iB2AkWXXiRH9bXgIBDlso1xvUeXxYJme0xPymI0/5zOXGL9GxPs69g4Q5uPRC9UAOOOY996ambwr
AFGCJo/0PKW9TtpudlUQe6Ja8LWnfL/HcifZhnZG0igq8COmi0yD7miy4Uny1ga90iFIKkCL0Chs
dsYvfsnF9xTjAgaoytjXPnqlaCYTR76IdqpB4SZKHlyDazZHB4W75LBf8Rw98hIvMGcFG0ToIxJc
SxVcyYVSmADno/Sy76ah4861zMGfnEGVZvWEpF0kw8inCHOWbU2wZQnXvAE+kxdoENgBv+hGNyfA
obNlFuHbRw8GNWDNiLXXjYnzfdDL1aq0dF8uqTHS5X/3x3CMQQtIQORjgzCGp0v51xsa6GCeKUtO
puM19bwhOxTOZCUbCIrNHfFYpDcOYtrMC1k2J+zky/B6lHo2ldQBtgw5SXQE1v3c3fOkYPRjj+rA
ziqXo8yheRlW9gzxT1ZWldYzX86UX3i3GhpkG6OHd6xU3z2IdZG9Wamg1DVkwbRPusADi9sm6hgu
GvdQEzLEZwJWrhyc6M2DTzkI5BcBLtlJpElrFAbcBoh2uVZifa0j7Y2V7X0cMGkCEXNTIKacQ5BA
1z2kWcg/4EiifCQwPdsu/ly9sWJlATXimDwZXhNbPzWnY6I2zgDhPHTwiiJW3cKd1lbmOOZYJgfO
iYpOIv1bGnq3j9B5oyik6epC8n4cMoSgRmxZi3zJwCwu2IwTIe7su/ZKe6AMklKu0VTizGY/EO44
1Wk7GVsHrL5+W8uLMNrZ2R3FJmHgE7HDZTU1CGs9Nb/1g71qujEUKej/vqOpr7nIR3vFXio8Mycp
9w+n9ktQrJcEd9JW2+iHWN8nv4r3U+cOQyx+4L6otHBkEL9MIM+VZu4oC44wQ3YPrjZiScy5YmRD
gRyp0qxsznfObBmcU7+uEZ+rWRA7RZhdyG7GNtlBzfV03BPrPGIKppUfq7KqJI6lOC7Hs+/Fw0eq
WzoJM7/OBvNxjObpvPQg2Cliyq8ytngXcW+nUv34lpzuuUPNEiYXve9IuhX7LeRxZz03dHnmalk3
yo4lnQOV1CCpFpGZdXLjuQQ9322n1FWzMgLOjMIwfKOjvENITYnfiEbJmpUjaAY1IRyXR+24Vr/N
XQau2cUbEaC+saxrXIdTpC7QL4gcQBG+7F88BqHl27XxzZ3uNWAWOgXNABnkP3gLnhVShtaYjD+y
87Fp7K/LYINQsWlnGVPamjg51QiA+CQdFYsgu2R2nSUFmJt6tAnTvPH76O/rTF+RhKDDtCjztcW7
Jy4+y7UtLQa3e/tJ1pu3bB/8/1SPhgysY4IMO+m9EZhzeMdcCDUS4ZrVOGb2lSF4p4DNgAJGyMSF
4/fSfubLfeSRfOn5GiR+X3gmc5dIqJ2ME332aPPP7sX0eb3i6KwQ9i+4JyM4a1YFawlislbR5kp1
2jRVrNqhwDvEycaeudHNEWlDdUDeCeanCr9QrumgEci+UX7CagbNVpaXNM4JndwcgiCBoVgLGRbi
8mztAScz3LlLxeYxGdx/Ak65y/uD+it4lHtrGzIyEn1IPnBjEbw46InmpaEoQUi+XnGsRw+zcGk/
IIyhq5zRDc8FC045zYw3X7HkckulX9vACAjTayHkQJ5xQHmiexM/N8a7WO9os1l+qJV8Z474FtGl
yW/wyVdgMPObIs8/KFUpPFOZDeyLDyASJLclkyLYGPj9HsdOwfS5/2J7TFJaJ+fU+lrXwIS3AWap
FxeKSzYlE4g+IFAw+SOGzazKcYW9TeqbW0V6KIFCfIXb/0fPRktp7+MkL8k5Q4Rn9qxIZHBvbMFC
gHH+LWw3j5mIJAXQ4es+KtklaGR/waPcMFaPGsQOlb4lecP4D0cJWt+otXEnfwnJb4NiJ1p8ZZPz
0b59UgO+NilcL227knMbrDr330QYYa6aNH5Iiz7bbYbGE0+Q7l1xbKbU0nwEfz3JtCWIPGdDVNdb
2B8AQhdXBYYCbB7EIjIo/1lK466uvADTVCS9A05fuZ2glEmSvBxrckxTDc690Rd0S62kzCxe3Qt9
DEIqsw5rauitigvDK3EH1d3yC0Hd/d8ug9bSTNjxkRUsG/O0Qgc4GY5TMi2tm3aiFA739Y5j5TLo
00Cv+dKZgD9xq0bwTSJzFvy5fCFwpY2Kys9xcvUcpkW+ZjvbMZyhsNtmF9edUuvIAZ4zq99W4bk/
/TypykZhE/EPZGzdVHh0B+DFN68RdH53d5wzdxfUwFWCNOSopx/mhJw3o2VRuwfLyajIO93R9fPN
a6UY59aBvaHmcMUKpjYdXH6GGoaNxGmyo51dJ4RpMSWcKCWAyMozvp0bRwGY+jUk+6bb0KY4pHum
PqQF0Q80g325780OZCL1WXZmZYWGkfisO9XqwPHlbYpEJCcj4KsGkFLoF59WujzqWDMIbMG0mtAe
d7q9pYWpDcuzd4fixhOw/u2jne1+RaLdBScfeS+zM0WjLo66zgGMWeN7b2BNQdtiCvhD9qJVD9i0
It5vvLDz40udFMPFA+j6Uh4pzM2W4jRrIG+DPJFCvE0S/KKXTBK/RDZRU/6inEt6Y7mQdRpUa3dP
ZHssubA/yhQVGd+XZHLMTo8I5Oij4197Y1bzdYW9qG5OKLKcaoiwspqH/DEQUd0oWqe/erj0fd2Z
P7hSnOzU9QCgvHCiDbpbf/gemlaN7SQlwovKEpypj9hCZJG/BytVOfpHoLeekaA4V08wsfG4/vte
ijdF3WPtYIjkR6jez+iWcr1xaicrPEhdbLQgfmyV/96oejWWvGohTxWw64uWitVdD0Dx2W9Aro2/
sRK+xnDDWBGpNjU1SNsFPX4P50xOAL002wzVQ7c4nqsVItChmgbgEdXj+eWriockG8v36gsqd3LI
l3W8ldQgrOsGWwe0kI+8BrR9oGwERCj1ak6Y2OZd3615DqM9eaLREm3uDoDCJ4PDJgdDZK6usOqe
PecvWC47/DyAFEgQfjhTx7n22j0XZ3MxoiewSszMfg0Q+6KrpRyhN25gv5YZwDv/x80bX7b2ksKG
QC+x/7Osz/Th8XPcDpj16LfTO2//BRIUj37UiR+V33KkCTvSyCGQef7R1qCqaaDgzWh/P/WjzlZA
WWvbmM/hQOq5tKgo7M96BsBdIjXv5ex+EReK1F1yiyTrNUG3sCxAXce1Gfl5B5nPnqxPBWDGw7Js
PHLMTkToGD51A1el6TB3oYhS2oBuXK/1r3gCYQjS1RUe6eX96kvLCs/14AZ6scVgWe/yzHPPaHJa
F3yK/2ghtirDeFyNa0TARCCul5b/rpmASat3nD74EQyAWDWlt2A5K26tojb9sm/LCbbnynRIaQsE
c5UFHEPxDAPrGUyumi7zoAckah9YP8WYUKOSC6zKdlv/2FueQ1y70fcXb4X1LLwHn+d9z0HyrFoe
3nA4qgdFDhRmXEmKwhFh2Z8ZWVJYfFh6ipag52bReDkUAd2EJ61KKNJs9pgWuWzuEkUCEBtYQEI6
zxNGH3vYPfikecVIZb6pvg+VxJJYQ9AejyoXKmf8SRvWbOmvsXRRtFQdI5sy6iHlU65WVGuucmXa
oi5NP6O6ZBjpKP1k06yhyezT6HdmkieId9l5e2eYfsKoEtVdIX8GmaNLLrku4LrzX/JYUw1IwdRM
9T6jCF4jb6hzmXYStIY4TkavE5HGHXsXt8UHLVBl16z2/eWRneC9sw/AuHGrDLTqhJbdjLdWCNYC
KbGRziWhjudtDkVFoC+mSD7eOYBc/bL6DTt+00mSUj5latJjuo5DF9x08Y5Fu27RCLyfoQVVWipF
OH6ERTYQAoy69IL0ooyuFeHmIb3TR5g0mIBVjJ0oh8w9SZCWyL8lLTsgu64CxEycAJnPfXE9i/CG
t9UQbsrfGs0Hw+S6x9ApLByyMfQR6mDah3r1yFoCobRBrJOK/TevSoZLpFKgcn+imN+BW+q234YU
UmW0T7fKeCP/au0puZgHI3UJ1kA0W2L2dqrx+g2tinQUrvgFUMTVuOjijsevlgl+8dZEQ3OFMula
xvjAHJ5p3CH68e0VFa5outmPCz7Wu0ptsLWteyXUu9u2ehKOPZegQ/UM5Dt8YuRAL4ytgyIt7p/4
tfTKp9TNq0IJ8wutXwoJiEmGSC7CW9HVeypHe0w9HvPb09vE7Jn5V12PCLIbLCyIh1bp5GUJgJFJ
DhemHkieP3ha+d9Pg7Pv2frpI0zwi9++ZRkSGYJggjnZ5zdvB2MS9Czh5qy/oNXnri15xVcnvCzA
dx58iSiEfdN1O+T6rGbWcA1A0+oD672lNvHXKB5x1F7LcyQUfDk3a924J/RsZnk5WWPoc9dYGLU1
Ud1qaIbROvKIhD4WcMYsf+HAh0bmYs4FnC6QzwUOpUAFVpCTCp6FftEEhbe2HHoMVPsli3BqZ6Iy
44H4SASqceBbzqihMWg/ZCo7p8ckrICKXgTWHDDQrUhUnyC98G8b5Bet1DGQts303iZwq+xrNehV
Remo/9GOWqOnNoZtUeVHuYg9Ddy+7s6mCf1jEaFAyIryp1K1fdga+tmmgBAcMkQWIDMDc2vad+9L
oGQW8yRjjkoY9GJ0ocgFh1QmQsvIuliVEMT/EiljQPGgCfKL4S8Ey7u746rouOzxvvQ9Uk4Y+c8Z
mr6dI7mW5veCaJ6PXGeSR4BSynid3bAW3SRzDQXplYxRDGvDkM3z14T9Obo5q/jCjfNjQsxMcwnM
YPV5JdCbR50SRNRoQ4Nl9UZ7xP8aqlgFxYO7sqyuRJHbMx2EZJe75WipvxIm8jHYXmS8o++sr35d
Duxpe8XNp94NJLf90c5dHmc5W/xV3q5lF3n7lwehJdXv+a/PaVs+KOxsE5s8NRduD2q+Ue8rP5Yn
nn1JRFayRbsyEV2RK0Z00MTKBTFm/g8DfosgkfqeWWaB2vgtrZ9TrhC163bM58zUqSaQo7w7e2u5
UMWuZmdZk5e5xkAJBhJlgB+9Bc7WlVUjK+5SRBgaTwK6KDZWUPHZj6ErTM3RSZz03ZJHPkB5GW5e
eiArCPdpeg2lAStrPhuSx10bmmTd3r9Uh7zn1GYcsN2K/jDb3nzAtY6EIeZLcMMmSZQG8vgL/k1W
0solg0QFa9BCMPvl6Tiv8KqmUv7jm8QzkNucBPspVXd05Wy0HZxZ66wU4GSA1DZ7XHwLorcLCYTx
MCRvc7SoTA/0Y462no0pa1406hOGLtP/YFtNcZ0Pb1nbNt2HB8a6dB1G5nCH0RuQPtycBXP2mOOl
qvx1tAHem+Q8JeR5a7tx0MFcaxz92mGplZFoO7WsiNcLZl4evGbr0EyfS/Tk7sxeM2PH3ON5DJUV
eseQduguvmK8ND44ND8SqbzXbCV5esKQxYLH27FeaEMH1JcsULo7qDQrmxfXEsgfy7h8o9ETrLdI
9IIqUSHEAPZH6w2qLo2+nvXBQoTf7G+e38bZmofM9tcWi+AiwIWIb5WGqeh/eT74SkcFoJhs9idf
RrCR1CewsZOSxyuw5H5tMVlRJ/G6IsUk0odbJgteRphYicKYcd5McHf18x9ohW1m5ct3DaIKiqrs
+DHttGTfInf67ATtlsojMAz6xARY1pryUjnRqS6tNktM83/5FqB2kSQ/zGpYqywb+Vd/B1YpIFfa
AS3NQI9qAfGMxfT8VDuYZNERkSN1PVPLV9hzH4lKpLDGbWyyhKRQlvBpdL7ZNLRtWm8wgUPsoygV
ACB3oQkZtCnNRNFFOtMG48YDBDJJVvPTn09OUi9DjhFL7hFFGTOFVL+XtvXcb5j1q70swusJusbt
DzsAltjo9KL0F5OT7ER5AHabmLDxa9a9eOnvyh1hXfe/V0mQ0jyNugBcm3FscQoiCp40rym1xbel
QlMwpgXo5PUkfnYtPLf0JnZjHuqJZKFnFnUHyxS6es/3vbhc1PFGRCuIIFI5rx9yOhqGVbLmcWeB
eew+4c1GdEz1PfbgW8z/CfeBvG3LF4eJsn+/FDmRPBGzAapurR7/HMSBGZ79Y/2DL+aqn8Gx8fxO
muqlSWBUTCig/KW8cl0UcdcOfZWugGlbTS9F72r0515Im7CliZSp/hhaIfYgkL3BCfCSbvmmlk76
qVezHuaosgCesAGumqKbg2a4S3vuGEE6qkoIRIdwjoV0W1/3kKP5C309jzP0eZiRVV3w9lOBlmdv
WpjVwHENj8TgylWCR/HRjbwO3dHJCu+D6PM+dR5hg1rbNuWKZ7lsDtet2QV2vVzzv5Cak9kdHtP2
/PvCPKBal8dn4t3FhkGW3h/VmdoP5GFqRiSABCC1SB1kJ73xXI1To3rNKhm4ZmYnEQfR0gxB0hg6
r128cBeFXcBhqd37eR7uPdaTkK0tb8eqBJqqlU7/f4rihdZXpBQnAZ3yAYRWV67kZzg2ymcPgKOB
+jlpRLnGKSkizAJs5e/rwXvPF1lHe7kTrmAnDryBJHjQUIuvN0w++B+WUqB/DCJCmnakJxx4DjPh
NknWVoYTFCIxjUfozWaiUrI9yNSamJ0m1KXX95wo8yqy+4r6tr3CJXtbUTyNuPogmWF54cBU2lBL
ZxrThi2wTBcucoaulvx7RUP16DOBkWvi6frfQn7y8Jt35Gka4H9NtCB95Z1HwOmyuBbehW0Ltqcp
Jq7hbGLla5qIJA8+ni/anv688j8itIfhzJ1JLtOErU+Py0jX5SYGnuSScV+aHi0HzhyTB7YqLXHS
y5BPb6RYRyDSCfK1+csuKFn8FiRRByqshg55wB7CwgzYZa4GebBrldtDOdLVB09AoJ7Mn96agh0L
V/9SR3MNBFNEe6muVfJRks4uOfrev0942Nnq0m/FqsMNlhbGsKjcdmhw8oN33uYI/jOFuvLuA7t6
tZLsk+1tFbuPzSy4tgLnw6eqNJ0On8tVs+iPi27lCtaop2pY2kLWJ4DUwsJ1lk0kMZUtvgSmJRv2
imSsaGZ/1Hse4jjx5CzTDzuGkyN8BhN3ipeNgQhxD6uo38VPPaHog9w15D+xVpinRppSOwJyL8Zk
/UEwh4kr/wnpKs0lRh2e91u8q3QF4XthAvZbn2JbM5pur3BZ5qHLwQGuTIW5XKLuIpvpl26T4R80
ifvaq5kLrv/Y5YZKLm/sftBewkB95+Ymik6mPndi8Qa4OleXknBfux8YrWFYeLN0RbiQGdih/sDB
O5xKVGrPmWWBs4LSWTZEnUnYFW93a1UdWFv1jcoKAQyZWMpbZK73pBhaP45xMAaDX/YoonAXNECN
UHx2rIoNePh1uUgQsvHUxX84MU9FSzBwUxoVMzTOiM6rDd9MVSIYp6I8XuLaCuQTjXQDBdpj4Qof
RY8QFnN5lRGadAVcSh43Cs1ejnD27n1PL60DuOMw0uC9JTdnv/AHPuYeN/hYdArKEnoTH1MNZSZH
Y17KMy2bLCTTFWcdbIJ0cfVNejlPeA1w+QZuM9U6VnGyW44ezL1UVn2jVrY4sAf2MW+TPJzN/V8q
T5Q5sLuXPRIX8KABFIQji3ozEWxO27LMJ4l9nGSlWS4DYaD+jJSk49D8r3mxos6H6PXDbgE7nSAd
vEHjK7VHdi/hlPxcP7rai5xRqJ1wwskIuQ68/wdn+sBA9eTia2ALK1yMfyYP0291AhoA0GlzWvZU
K8a1E72R/f+ghGRmdUDz2aDvP+cMckGhW34Cte7nQ+0k2krY1SMnGAY4H29WUi8KDrq9i1pqWSYa
oSRCzo4VSr7Vj9hUC4/7PVCeQIL6MvF33fpeI2S9oOhcngXyE7YX+pZpShtAf7yxAVnV0VxHCNuc
vitlu60QLDyfrgyvAm3+ylquWDf1DX+0RD/bhAbDrm3+PEpMCLO4+8AhMS6ayOrz6+L+HHNB0t+C
O5kjm03rSKUtSFqFd5J1dsloo48TUcpWVHV3X+JiW6m10adhwYEexrGniv1mohH50ihjiVeKY6cB
Ce4Wf3OAIuQn17/PBtJTeKLioGDGVStWj8InxVLHGiv5ngWDU/d4RTomDaLcg9nKTQdjJKruLrpY
SXYq1tEs/tS9aVad3pNiNGvA6Glx6P6mSRtSV8rQqf8L4kQcqxikOs6y6iWbd+/H1Od8l8+VC+ow
Qm64F9j86oelwP0SsWNi6LS5jTwLoxkEUtrk9s0N0HL7SD8tqKATxsfg76Kjmx/m3sKKx9Hzh510
8WJhF4uWBTrHU2FSZyQhwgDGJBM79yplJydW1XhdM97BcrVb1TdtVTpdk07urVlBIf/J5GaEWOeC
I+Ylwjv4CZRjHKuKjusipqtbSx0+yR9wtPIg0cxohZZZj5X7wt2lyH/envAzv80T+C0pRfmZZTSP
1wcZZUOpOXJ+BC2tCx2VCViUSF4sxpwCuB03XCnyFjFWoFuCxQoMhQLwMCXhJd9TLCJ9zt6pp9Il
jftg39Owo5x52hYKP4iMYkvoDd15ssJg4jm7XNJiv4xEGnY1WHwdWy5RAbCkM81bVe8Iu64Jy6ME
khZ+qgC4GXOxyLIsHM59h79kz/QIPObCsn4viXcErFWUnKWqaBJ+fMmjxseoHasGjUmAQDGZ6VEm
h5QE4S5GuDH+a5ynNZAA/cgUK4nGaIoTd97rx15CYjvdwgAfVwSsY/Z/XHKAnqsaG40e7Boys13Y
8rILRQwWoyTbViEFp5Xz8MYB3yWB0rYIUKBAfXhBUUIgEZZaQdQ83aZs0iq6pKYOdbhddMQk+Amr
N7HRWMS/2D87/t7kLTB9DSZWt4BX1oJt+aO79YELnbR0BW0cmN/5vZS0rQTHIWxyOG0CDZ/8ZiL8
bpN0na/waO+dkPD+xkCbpYqtHEYlO2v65UpUm0h/mL1T+La00C/N1VavY00uwM8vbsvZcXn0+GZO
+hhkNELpigrIq40WkIrrJqdMtBPWFEAqAq7HeM90CO3Xd2e81ej8QyhkJVDJL68eqKs17fGPK6t3
+9EocUmOnosW6INtBzXrcs6PLQVtrveifWDiCBuVPd4h5rEvuP6egGTqRjaOBI1zy0UVnPQSvMKv
yzkPVvpFgDPFOp0u6X++Hi8b9I58AjItPDlXsWyq+2ktXk/fsKBwpvB4gxFIKzpKryMV7TBfa7Jz
ZdXNm8CiQ55Ft0dLXdB7DCyQ3MW4mVktVZex2RByoDkDD7W850Ov+BJqXecTD8bMG0mQuMg+1Ncu
0irbQ2YrjtRrNro0H9+xlqMy9HnHwcLD+9MqZMXC1QUkswb7UhsJ9d0QNev/G6Ihmac+r1XPZmmu
PqFGzYPdXlKV2aIfW9tTHebfD+wq92nPs+VdA3On8Sau1wtot6HVTXo4ws7nXUczy0NTscC0QU5i
GcFsX8kqEYYH8DMkaIEmt/t5nhlfVNBCDiX4I9xGWjguLJdm70QHd5gd4FurGoCdR/46BBiqM4AB
wLaoqAETE0ncVAPbyG2IX+o1CZIu9xJZtkiNPjLjKBWeSViytBYhq1sf7F8IcuJuRs09G1wCPY8S
X1kY/fXATw/Q4pXaJwC+kjn9z3yHr7YpT9QnAnBSPP5iqNF9fTAO/Ie3yKMV8+jVraGO6yeNo+Ne
32b786AvVLkUCrpA6FAJXVWEcMIg+Bf3wSXytJLvQTvb9VnI7Cj6+OOfjK5BhAdEM+eEMPjzX3v8
jWlowieDtQ8xDiotLk51a990gf+dLVfOjd0qT60K4Sq2mrBNLyNogepo3byfPmvds00xAdKcuJwd
oZutS3wa2u+ZzlDStdDkC2p0pwseAalIjzCKexoiJJxjwbHo+MCkgrXgpMX+3MZrDULq7h/ERhr+
3RP9wJoN8uZgd2S/Lp5rN9cwu6YdttEcFmGCGyMI2kO/d4Fgq+53aRt2b4Ks9BgmRXzgkozz0Ecn
f1FES+ToptVy/ZGJK8mwucPC7gAuu731pXj4jj4Cw3UZGlrFcZZP8QLEvfCuOMVRon0tJsKR1G7u
ujqUSw6bwZWH7GiqLoDcGvE0mSMeXg95Ph/3eRkE6FyIJBJCjWJrgn7gK70PQ8Avw50Ax8W4eVVO
r95nTVrj50/PXPF2f+xa4dVOMpH62mwkc4dgAjvUnKXzkcQjWwdntkonWD82/7GF9zvIxlinq+D6
Ab9cR1hiM3gFGYDL4ZfgTYyLCZkytDG1cq+HRXEmH++Dx4xVOs5/ufL9tkRem51u8Mij7onz6Lcb
KikJiBdmGFLCNfQ3QeCA7qlyXlbBJzYNmaL7+7VJpV6owt0+oRHpJV+3NVlVfL9H/yl7cUCifR6P
L5zbSbUUigajcRi5ionc37tvUlUgObIr0UmVhb2ESu4BDhMYYkCHyXMbR7qkia+8Ba6jgfMpdSq+
Z7LbA/OnNRTxY8jsKsxvRT/7HLBPe9lD5zFnApvgj3jpjrAFHgSHpsabKkYAmtwuL2flDgp8nBhP
xBHitxb81321ej5QTYVaLCHoQ1hdGFsr/0yDZefpWuA/P+OdlhYqN3Vij+A4+dnIG4Ehh0hBzKUb
a4C9yYVprvb1mJGejU1lW+xRE4n9Du7u7b0P6tcyCoOkMJAEmiyTP8D0DQNP2tRorcGnV+zx27lu
VgYUOr4K8k/cv4laZHVOV0BDNLEjVhhD5h3k8Gz6EGqGDrOGEL6wqBjlMQNM1BcJFZhAuhypVn84
WxJweO/UhdHeC2ymqgHz0yVWzgT7kMZGXeR1UPcR1gmY4rlXgvpTfwsnaVtdn7QIv4ygivnFKNPm
gJ2ynNzXsa5ydxY9PI744WDoTo+s0crMLnqomtp+W/lCHwgmydxcM1i0joGmt+Jsz6I+scJeUctJ
oCYjLHKvQWRMyA0PL3PdYErkjF9O+sRB9ZPKPkBRICAw6yYdVm0dy751So5fidpFYeq4xcP5cNqr
vzJYMbY1OnxrLFrSO4c0Uxq5r2tS8R1z7dCGye1fS6uHwNlVydOTAnvIZjkyuvETBG8PFb7juVUc
2DB7U/PNZQl+AWCX5LzI8wb1ldg9ErNU3GtXUE2542QHvHiWwnEy97tOylYTMxhB2EMHRfhSp1os
bM728vjTlWmEfHd0rXs1WfbQP6LRvlx/J2JMfbxCJ7d2vrn6Vwe1QN/yEqk6JF28qwOWywvhsYVg
UdbZWNCuaq5JL7PBMDfw06UOc7Qm6jhV3ZQQX/uIzsnfLEBIZMfjza6sVb0l6yUwKDPlZfXgre1O
SPPVV6dZL13ypUJon/mKv1ewM2Ba/jsWF84RR4GiV2Piqpjg+Rt0k3QQRA+cLXhnA1GDxqdWXHR6
DzrooTJJSKdDmpgXeudM2/Sm02VvfZAd4XH9sQJzh3Qypo9Xkdzr2h0Arue+2qmrX+O8hyX+Lv3J
TIGOGTRMnYi5IrRqDmzXAR0ne1PHeMEvZQY3vCeqj6mZT7BtekqZ5X/B1FTS9PHgSL1UAwXNxfU/
ZZ1lcovsqJP+sCIutz/voCuayen/QpI3QrjLJZ94gJZyNblEV0vgnzxqGQ371NyOHi6uGChhTNtp
lxCh/moH9fEr/l5jUO/Vb+Q8xU3BJuoMBPODJ1Cs3rlUMv9a/Z1QsoVClMlEUZxtForBN7bZA6fr
XWvjXr/jMp6s/U7Xhf6UKUnJEeAUDJGIg/3n2yAawMpFvZhhFGdSLgCD5Dz7sct6ASAjs4AxaTcA
9xirWUUss4nQXTal6CBMEW0+2PvpAb6uZgw8MEtQ6x+yS+LNGjns2EdbDK9ZeJwiWzj/viAb6Xgh
nWFDVkDc2sE7dz8b8VNuFvhbbiLIWdeIlChl8vtwgu9mnrS+u+nQ1iblbflEwtXL/ThergZ3enVC
Iw03/lYry9cfg/TpP38UxxLemxWjuluRHI9kbQxD7BM1V8/VKgb8/DqSfMbjbEwWrEaYVa1lRoaw
6I/KpA/iptxK/KIokX074dHv2QMaJ095a4eaNrfnvi4ZucYUHxeg79YhD3qD8VS1nx5EJoSqGQ4R
S0ssBubRifGMslt9dLBZS3GAG5cQvj0VT98RITFAlTjYOb1/7YXeafu+VwnXD4ufTy3fuEClRsT0
D7SunnEn/JvaMkZPllV7oP5BuC7mnT8tbziJw6E/e/l1Eck7TIb3TAvf8NNsUiWVdpPy0xV6zrOM
egTGP8KIADXnkWS7z22KcuvGvo9JVaPRqW9ZxzyulzQx64JS3zarddylb6FJHNXX61YrpQoO75FN
ivCx5e+/Iqnfmqulecqp5B38AKwFozCKRTENkRPTf/SwildNol3IMHHSkHdYI21LLmh+PkCUDk/j
ZX0McgsZ7EcNVVWalnvNrFBzYvqHQbQ3czmR/0DnzLHso25E739ZVJVOx8kTp18nI7Dwv5GbemiA
5G6X9ziX/7Ex1zrqVjKrD34lG+wmc92avcyu2IOXc1q/3jrq2Qt6HhC8zlI/y9xg3YPhjoMeOy/s
okCPEPxF1ULCD/GBY7Xg2EGr8aRZzG4U8VjspgzaueRk0hMjtLuIwt9v53Tm0hXyoELh/L+JAdRP
57iDvOsSxfEemeMfU5m5daNrSow1eZWG33HAbHFjbaHMN04zHFnnKJQVDInE8FvBdEQvDqv+u/E5
MWtIccUcT6fVBeB/J0DERAZoq5GN58EWGpmOV3DeRnFpDKP0qKrqmVllEaJbHMJr2wxTQQRwVPZq
Y9yRgyw+bUsxVY65SillcRC2vjPFe5kD46kZ1D/28mC/9x2w3cupgZTvytlNd/eklnLLSraseZkd
fk7ICeY6oj9RS11r15X7sK3QeFhHUTWtA3pkmXuoaJkGvG2wi66L7lyyr2Ce94QB+peaP0maLBuH
bwZo1s1imxJxeIpbP40G1x4ffYN74JvIFQuhk/aktOioaJw1yv4pM2htc3j9GUVISSG053bDtwpO
qxjM13lkDF/3QsjXsaBVX8owWLM16Y7cIqr5JH2cBv0IwpjpmlZ11X3/Snen9wr2MIQbIwiJ6HeZ
kW6rUPQl7NkBQASwYaM3oqn5EYO3hx0l/bgsYxn0586YaLiaz1th4Z1qYG2/jZ4GO5t3eNuyLOEx
Ju+k70gPkx3DHNuYOwJ0ANai2iiynQHVDTOGu1WYxv13AA7VI8Dds+C1XZZsO1o9vyM2QcGxr1F+
vwZvB2UASomPRT28Zpf7Y0zVge/MJ4QVXVxVAnp1hKeXffvIVZJhbgqunKCb8r0WGTIqgi7lr45d
Or27pm1b6dOlIg5BrKMPKMG3FwMuT/wvRWCMMDAgiJMYEvTz/GRXnpVWBdzyRRHc+OnlrQ1VVafu
73pOE0JnjHSFdQl+sukYMNr6muk4l0sPJpusYxzs7+r7iSE5yX+V2D0u7kl1o99R6O1WvnarzAoS
ZFJWKvf8OuZCCANtUJR3S8AsWGDNIAUFwqd7+hmwTxmsYKZMUs1aUUDMkjBM1AhBzJ+BBUmN0EFq
BFWIJAnfwbfllekTP/f1MQdolSvmCki7H2UrKAUa2nHnoa9du0eoVdJyeOUPaaHK5hQPyorvQrb6
qBnm19+tXlKMkG9rv10LjGeWyGRoSQjmnpX3ETa8DxFAj1UpgCmhgh0eDZxLIbqOY1UkoJEoEWWI
4J/tkGbLz3hApsLompW8Qz9rm67b+E5YKwbBYdyc/uBfp5UahyC626pOpKAhlL90MRpHxKmMrf0O
qLm5VjhOLGuxBHg3aKzVBTXo2V9qPt8m0PJWtc5rXtW8qwApCPhVO+iOXqJP2UJAeUFFWJq3Jd+/
R9nWT7obHAJCNodnwA5tzr6rhTdlmW65kZt3YVjS3ZY0b5bOmQ9erEpD3bMfD5wTJtkXZ24tLf94
DF8QJvyZfEQGfRSqs5cC5sepOjHH/+rXK7Qmo/K6m0tm1nEPQ+xwZoBMLnCxocGjqQfI0PYA50je
QyJk/D5Wkfco54WeUlAXyNyBlRFJofJaz/pdAzcPoKSZgsXdkY5F5IhPlfkj0qNYXcZKCPeXQHeG
TbGMmFAC2E4SPP1v51az/Si/5JD3zcyP9MXz73RlWwU90ASCuBzVoikoC6N87wLa7vCLYdaq3a/7
QTzg2LGUo9BXCdiPXFWPrgvG72HCip46umTiQeojkRoSEM4qYDcDnJwgr13sjXefh3Ch/SmGAZJ3
/iO9IUhni3QwWCywJUncV6em5BYHmfCn4DeUHXXMXUPWu7OiJChGEM/0xxUlBGfFgYrOmp6oVQoL
tsYAsEDerLL7Nb480oeoX222tlWYaarc09AZQnYMUV0wV0sbqiq1y2RI6BYENDV9rZWmfCy2lNDO
cAQF+yBe2souQJ31R5PIPG2x0dSJt3DPp7ZwiLExNLxVTUXEE11Fblg4XT+ixWy6oIPoAboBJoLf
bPhs5dtMHr4lzj/rJI4r5Yp1QA6tNpqENFiawhxO+Vhn1wMXIilazBQH1M4hdN+1jRlPT1MQ7jlX
KLG3BkihRAOfqN90D5ybuJfc+Qe3KKnfKpU35vXrEvH0ACbRo9pnp9ANbajo9UnQ1YvcTIU838Z3
IQgRzM49i35ZmAL1hgE5JRBvLtkR73J8SGs/yoBmM3q5qd9dq/hafYsIBsAie9gDW+CrdXw/EXdV
OKRne8u9+OIm4YSsLbZqjHdm1xZGKNP2e73aeQRF/W/LO5jQx2tba9uarByg+3uhRsF8KPHSbsiV
y0jdyKWXU68YIyUiaK+3GkXl5PRIf2Tq7tLSBfXVClRM7Ctdr3i5+y8bbht2LHFAuOd2+BRrfAMn
hdl9YxIbdCqtk4RolS0xFJgUtvv3+1B1INZ8EzHrfjbGZ9+0e437H29WwTpTduoBM5j6ZYFXR+Kd
MpVZhgJQiCRxV10BylCFHWNpTcFxaMgEvqNq/xSmFT+mgxD5TiIJu4s1OVswc8/bFQhsatPAFaop
8n3aooy8ug+tuJWq+GD0Xd6aPB1CfRQ2301SwwyrVWYVY8e3wN0Y4ncTrACnsxe8dm1vY9vh4USH
m93wULMH3lCO4qe4aZjQtH0th1izRboc6KRTmzjxYnrZ4Qs2s9zrSH7QzCHpv4LxUJbwSXqBzRmN
F85jDH0ppGINcEKFPKJg8dnd1lejGsSPWBPFBMxBjLqflHy0S0andCUXN8rPj7+14lHDi5Aimign
0uQNQ5ZCo786gJfoXg7jw2PWs8ZMJxMGDEVyyc4WuzwdfC9BsEB58DrMNurW4SP97MG95GXjwrX9
0agD1SDIRNKyOSsatGeoXuTLjOFO156Tqurgw+0PZRtPR5a2E5pscLoY45clFDHqD+AbvCONTU1R
b0Le1gWsYhfxoyFN5kHG6JotBjegUSbz/80W2REl0D1YscjynsXsbD9MjucAOFi4Am00/Hefm+Tv
ls71oVylFiW5/Bx1mO/ZeX6RUcmYuxHocAS9OANBuyCJRaE7MF2k/wPgsBcjsHH34+5Rvtw0Q/xL
vFKQzbiwZOCaASrgifRfVetM+1quw6x/CjcsqX9egleMB4lWhj+PoM/fNRbjdv1Uy3uw+rugbnzD
WHH0ClJoUcHLt1gEOSwiZbz4jWPcj/+u6ZnN9KAIyKY33kit+YODmrWxCXHSGMzWxUUCGMCLdO9j
tiBbjRE/c/0soBVw85qAx2dC5+92AXsy1yPJqB2qB+kB5Ws8b5fb1gaVRB/qN2brpnWBLkic7y7m
asjijSM0DXt5SZMJCJEhJASjcV//uQSaXqs8ofM3fscVb+kENeRKiaK7yYZFRhHXAMI7sX3lWC9d
JstkchAwRMLIta52oUQZMWitbX/+0J9UwaNT92nFQ1KSS5JJqIpday6fMgIN8+ZMQHorayBN6I7Q
bsydKcwyaAMAeScaUzs65Op9F/dVojH7PrJWkt+wap2UQgz1g4YAxZ3mWIWvqVrVO2oyzbWbZ/nK
5CIxakDVGsHiop1TMWvW1+f1MtmhMzyTXxG7nqDdojs/tLs+CNHdTWt0+Z5TB3BQ0254AQP8XSN2
0ewd72pKxijTDNIEgHSEvZp0VZLckCCW795jege69iVHYJFrWMHhvoJw2zm7sTCQWl7sFtdi0ICK
nXG2ug+x8hBmuKALBSOWagECWRiUO5v7CWb/oqIirBFDAZ/GUn9ZEPy12maSqiiOdAHCUDUD7qHh
KjFNmZ93wk1mYOYTBCLRHOdbYZfgwS3kk6tiSaymoBVUvYrub3GzGmbGFL7anJTJbZiVWoKoies9
LvX5bd1Ky0NqUTBBRR/DNglBG5xgj49KyWbg5hFTTWk6YcdqP6o9jHVvRhyICrOLpqifhPF8J3ll
9D/8PnyFqzpM3/PZuQAPIuRGhF+LpFgq3pMbSk0w3EWQXX2XB9hJUDGhjf3y1JWfT09fg+Ghdue5
3CZopxkaIbCt0oCJ9bvBT9cixAIaMQ3qztuCmOXFtUJbI+2ztXmjt2KiEiBeEVsaNZ3sbHMSyNGP
Kyian8mJkl0SlXBt58M8WWtd8HHZT6jnDIaHXH9J5usyp/BsKuAWqMqQ5UfPS2CO7aKFoSnuHcyk
LLBEpu7AEAqD9RfzkswgDxR46c2CKMGozKNDau6ckdpFnpXWYScTuncDJJX0PWsh5y7ag8wXEib+
VE/HTDUsy1SbSZe7Nh4qVHk5umpEUn5NjJKX+CDJiTee5mgO4bfqLJwn3gL5SB6mEWYwN4HV9Ztz
oq1mvaySOOAsmtBE08iBBxNncZWa1pvaHe1cHnwfZSwCcT1ygU6QeBdB9ZIGoMS4/FXDSPk5PRGk
NKN/bGFoAHj3TJQoCG5LUhZre3OdRkSUj5JpuIWIGo9CGOBnDHQGu7HW/HtzhLMlf9HtG3r72ggq
daWEwHEB0VBtg1KJ6SvpolkFBW6CTj4Z3HrOiIOQ6CW1VxE0pgf5WZvLYxE4/kuw8SG5VdB/wrIf
DLiy3qMnAGbXEnf4448CwUcheKoWLDScFKalBFKplYXH5NxRWVRsPxEW2jAAHrwMOXzGwkRe45Bc
8M16xog9bsmlA2vpM/CC/xr3umM6Rjf92Z7Fk7+9Ia5YsP06shkKsabuAwxBXlmOnz25pash+JyD
CyiSERr2QetC2T2mvhlBrfRyfcOVxiPF4Yj5y0VGj78eRCi4+IlzdrVph/O8FgW3ZlHxvgxOeS1Z
1c+Ac0ZEtXaTZd5ZAx3QmA452OR3ju+KsmSWieQgvNmrUv6mVdfdEsHmnie4FaOjYcUwC2UcgSoi
5Z3b9ieCzwQagEy1iVzHBE6/TZpjWfbMrPAweDhE2g+lSKA6dCBvO32Pf5SLGhSybTbaHRp/ek0f
GNlySoBsC5rSUUacFLnUMocFQdUtRZNTjT6InSb6+N5m4IOxwA8czerTn2wKBth0Is3GU4O7OaCJ
meU+aexoGJiMNxE0FvzRFBn6GK96r4h6qZd2JTWYDlIB+hXZ9eTytVZKcKFa0Vzxim8Rj1rD35dU
pd2Va5Vd1OPFvNTdewBKrTbCdf46og+tBuGCDCX8pn95kxaniNc6Kemqz4MzwV2L29Vf97TnNsT7
155VsX15/Tr18T2uZZ/azwZOdUqdNrMMiog2gC8VWj5xmMi6PHLFQI6nEZHyKIjIVkjx42qMX2Pk
vGDptTbKr+C5Rv+55bkC+s4a3CjQBUMiq5oF1dhbpxcXsNTg6LfI5qBuMUJz0oK96Zhw/cBUVHz+
oiS8Qrm5WZNL+cUUBa4iZRH33Q0HMY7oauFJKTkROId2zza4FXJkiWJJUOCvV2ha1T479GbNJdIG
YLIbB37TNKv2DlANRbXWCWFqCq0epqDEnJxtjIAN5feXO03zaWlCwVI58cCzv2XFfY5KBTLBGzVD
IKxScar+7X30sJ1Ae0uiWS1RJ/XYOFgi0vMtflJk1aK1DvoBD6eV4zhBkq/SXEDew78VfHU2OQJb
SffTegp/l3s8DdRlvFLLGAdvFG8WoNtdzAdclXyrpS7rOFOojPc6xHYlw+3ZYLdaOlHc/sWh1LRB
02e8hpdgBgxd4A5TY/5aVUaWs/zlB96unENExBEFocyBmPQKbEyEJa2fORezB3se6VolYzfn2h1q
3bxNJFlVsPk0zxqoy/YZLqAjQcMMlSskiWnPCLngmxC5J9WjIL4KdgJgYxbPHf7zVbqOEUFpIZZ/
0suAGIVoKGh1G5rJ15KzWwBGUbitG0lZIibtzL5LOW3TFaaZltGLOXXWjPaqlXEJ/mwK8P4rPSXx
hZu8E76lnni+gbW8ZRTsZ23BBdbtckwq82KJODBBxzhlO45YQWCTCoYBV7U7PQUJEZb/XmV/KLoQ
AEs35xNja/jD4RWQ58z4vD9e2Zrb+Zossvc82ZvTscYVa1ZR7cjLHiXgO/e6xbMIkEtAift7Xzu4
K4ti6Txy0or/wJcCyCpFOmnn62dz4fnp6/pCvIWJWisceuFKgk2SkEWDoUhALzCTVGorI5fAqeZL
elFPK8JxumTvMEKAxo6ZBy5Rzn6lEKjdYGm5xQsB+jKp6WINXN89Nj+ax16kqKOAZHHJTXJRLrxp
2EYH3/4VVyKFx/ACn6yZcHZ+upDqn9JgRV0dYcuCiaOMvjG9lvkbBcqlrvVXUSxguzS6xdM10R0N
OVA9oMZ7ccWbgxDiv1gG82MkYTnDjAY7vzd58Tg2IFbv75Vi4lhuw/5WTLODLMuPCspJlrF70k5x
uZbPWWEbRpsi6c5lmOyF+LPHctRTE+lFC9WYwejw2aZSD8YNo3kEfdOgYqnWbefMmS6Le9/DBuGu
yEq3MngnnMAFd6dTKAS5Yhr90OZDQiMaTaNBtozjTTOl0IsrmtwIfJLkRSi7WTSa251r7xC9td+T
SO726E9xEaP2LxlXDsnDneJh6Ov14ZWl3Vh0ledguxh1az7DKBYABd5sr+FtDVCxLYcb7aZ0WzFq
bgko/RezhG7ofSz8EEa5AH8puXa2+6nJmLUR48LJ47rA6GZns7YoS+TGmuKNR04O1B6PxPXE2U3S
unSsLIe+DTYwdFoGwQuZyX0ROqxL09I8O4J+UfXE8Wo1Y1QbrzYaQU9ac5cjrwgnSnvv6vRSXyXS
j09uL4x9CSq7LVKfjOK2S5L+R9XI8raAr8BMAYgebQVFOHYZItq/L0rvGqEMGQ/KYO7wDhejKRee
gCtC+jIepn+qA2KiIWVhu4HCYI5eCHxM2Y2gbqp2PMonmRxbjdjNgtBFi0N0F0BHQYFMukP9Syin
OCsarnxthtpdQWsm3RuDk6Bx83URrqOO8ZXlcijtIHbgMTinS82GsRz+MJgYzzRuivIFukhxVBPk
5zWEC6DngeaAQ9T7sX7c7sbEjSzlsSczeOqepS2YUzV6H8iROxAnxQgUEf1zC7by1N4ZQLHPyQpn
ZBifgXl8w4851IJrEfzYwIEhlmZghfeZ8cjeNrZTLGSu7yoHaRtv/mFOix5i6hHgqIzDj6o9Bheu
1CvgJiF4L00u4MuVveE/zpVCGrW3mFp3W/eMtLKJ6DviDJ9jqGMDgvGud8zYy7senzSOBdnqInJm
1+5csJSB4N9h72E+PHwZk2kh3TqR3rQ954xTPylp1esXXGRBbpOFx+9OzTIo4SoJ+qR8+Cq2v4ch
4XOrC1vmAG1kxCmcZykPTelcy7WXEw2IJb1j/Kko8r2oD5JhjLA8wECA0Fgd0tBWKJrXtIoqoc3W
/Q6b4O+7Hd/99Q2nVKX4/nE/pI63axDGMMcUESewUQumhlt13TINfBZIXdFOJuxBdIVbib2hNuX4
5XF2Yb3UXVu6BsoFjdmdJgehxgsdVUlHaq3P1WbhzgxmBnnKB0AxEo0ZtEpfsU2jtCzGPRl3Sf5F
yZfaYT8yckNEVKmhRQ9Dl5PgN+ijOzvG5oaJEkyH0wBBZakHDBaJKWrrPieLYwD6BPsysNFxlqjW
HaQ6Rxilf3pkqk4q8bSHlKiXFHpmYXHputUi5wskz2wXfd5QXYFSvNGV0STm5KxYSrjJkVW6lhim
bToJdvghnCs46bLwyNNSSkEHKb9+RzbRAJU+j+Mt5kwJeKWMdT1NvcwsVSbVSI1t91ioXjuSiZdr
qF3ohcon9qI3ZHPUVTB07wFqsRdFVUSaaKvzf1+a+tr2x1g20md/873qcEg5PX2OFRxoiULcOnn4
sdy5zubjx5knzH7nj1+AzLDxj64gbuZOPjTC/zL5R7P0gq9qUbJ+RgjzJE3bSthPMQY2+NEsAAZd
GpKLZ147lH6yiaVvCseHwgkQC4LiYDU0VGclAy+4BfHCEX6CxF9MbpN4Xj3lWP8yc+szuI8Vnuca
8CsUp0w2t1Kj66Iiky3TdMpxBzUQ9KS5R8kp9kT1TALn8Gc40M4ewpZ0zQ6+74C8J4mmPJ6Bb4qJ
Uz3MB+2bz6V6mkU2w+ouWKAZCBevGFSsbS6cMcy6LdbL1SQkawzIT4ME3XcaDu9DB+UVoRxVx1Hr
gx7iHQe9vvJyii9S269YbtRXDrlmIkuVdMruCGEAU2UeCPay+1lwkD5Gh8vvIlIDd/vbx/gQ/Var
8yjvAuE5reFam397xeZoqQAGhrEeTaOOMA2UhA4PqBGvTCUwnECHivZkHJQdWT8/wlrryCVmWwpU
hYwwzzbSuUD32080o8iKIPFJpTLTNeZ7lClPQkPjEs/rUinxvxDAsIV0MDMkE62xdUgWWAxoskjB
L399/d02J5QofIqlOslgBeNymk/XKeTixA8c0G13bcLUqTHVdI6Vo3k5nxa4bdjIRpRp1v6ryLe0
JDrPLvvPXaSXWwg+t+SmcYf2wcQt3cuiLbGArcoAEshbWsnK5ak2q9K1WLPbh0NhUAQWRx4c7VWi
ZLLk0yULVrcRo+gT+pexCQ+Y3tqnoeGRsKwolWrM9Ca1XmRzvOSeASm6mFiJ9valSAGlncmtt1Pf
So1CdqjIuNe/3QUH1Gvk1K5sVpg7RG/OpuM+pYrKJKyGv6n2lcm3yYlweW5zHLHRUDJDRvBw/9bF
KKiuGoG6Q53FUSIXFf/+3RgDV8UJ1tAFITvC0Fxx42/6TRcZKVwy0j6H+71l2nCoUtEKZrh66s+/
5Q36gfUzXpFIbaSpmX/UZbJLnIJ32thtftKncabCHz/ldyf43lIsoiZS/dYlOMBGDPJiG36rWC3T
s9JoBnpqdk86pk4+mKUSTMV4eJNlURnGulXSGXMhWRhdo566N+pPP4uA6MmYcnqDz0e6ipl86vP/
kJPRQdt+foGUVwkr1jpw/pwwF/O27kUF6n1WDULjP3Jz9NbOQ/MPJCDiDfo0enMkMcUdaQou1Bv9
8OPWZGPfT4QFgLz34cfnsnNMnKVTjXUgidiGP+7Mj1BPe+MZ/bHWg7iqucgz6AV8MwkIi7pn4GvU
WJIeaSZ/Kld1thCGH62NKWUCmVb0P1WUCBAIkaVideqfmvif92Ur35cVUKMOWY7ZvSOdYatqk2QN
FxsbNxJVV946k/wowwUPFGD/THQqMDA1Dtn/FqsGqDMXrFzcThhXFz3E7DaCUVso2jQeZD1EtnaP
Kzg9D2vAyxLXs62n/xpSxO7Qmen6tdQF/0yTGwUa1JNg/L/uyrnCDXwdpIBfjoI523oMk6JekjL0
xW6sL4Qy5D40E95dM7oLGlTR1XOetVfrKstbIxao03gYQGxc0fvRxnFq9V6HvKPgclqKhCtDA+yE
fsKOyP1BbL4ZrGAHGJr0UVGSQFA0mdlSTEK7R6f/bWiIQOMJPrE/Fy7hozFM8ncFMBDYUACcPR3l
UxrogstfSawSOlncZUEGRZU1vgzKyv6HmvbrQ1dyoqT5a1nf14Jpu3h0wzLWWlAnVjUspWa//JjD
7HTl+yWxJchXseRk3eR9+3yzWyMqTzB/5eR5nv/DkskeyI6uaFs2ch/IA93S5QY7AgMOrgqUlmFy
cYqHwBvVJTzYmbxnmiUhk6mDjXIWqGdKzZGuH2Qu7K2/V0FiMM7D4nNrb0uZ886SVwhVqeFZs6v7
I6Q7xeXcrLxdDwQYUM++IbPfiGfFlTEZpjqDKQsz2CWDGUAw5EU7Ofw358HxvmNvu2nZW/f9x/SS
xrqC9TuxdOcf+SHf2L6fe+dO3NDhfwTarxYmX/2XQ1yz2UV5duY5FGIrp4H3wOyYO7G8D4+lQaQb
hc4/0ZR/B40Wob6lYN6rqgAkpZoqViLhuhbRy6h543Q3NTtOhHgek9WALm47Fzjro0lVhz/uLXiX
o5oNDgnP9dIVp9YAf5MAPdMJyh0CjjK9r83loOUo2DCChi+YfOKljDw1ohbid4EOLBmNKdlrOwnj
yGd16UgKt787vPVMeSP7EQobVBBP52Vk2ZHBcQepkq+UWfwr3uJJFR3Qm/2aSXsGP13apeOZ5Dgt
nFtnjlH9YEVxs8/L2VF2KgtEJj8cXTcSQn3F6URXTB7olpD9ytr+Xh5QjN5nh1/lkgKt9NOD/BYL
sr20DmJbX6opeY4BC3RPruLYgopP8hLWJNnoZ2AwVR//OFTkFCmTB70JwIYncHLiWt1FHKII2NCE
qihHv+9bhI6DWXibCR89qx87BsKDDt3fZ9iPjbYUqfczkLc/aL2hw9q4QoHXfrVknLbxjxu0Wd5l
kq0ZSsEIHRgbsBNrF5JyHXFgagffUEcsCRuUeaNSaWBpWUIkTNmroU9+XbmqCnFjKIu6jJqNfFRw
lfg1loWS0n2nRhPP0YvDz3ntUSVfoby5JxND9WbwjKLiEtykJN2u8wQ/ASAk0VZxFVzEufpL6VuE
sb2GVW1FqLsSjZpgxxRX0XTfjCP8EEuegh+rVIOX7qlv/PjdIglAzkzgGfv1dn6FsRf5Kpt154ON
4QR8yO4isJpHDQ0DxkCEBS3kOtv0lkUV+Bh/R7dm1tsTbTp4qS5wfFevscG6jibnp+ZGAqIpDoXi
/zW+6egyqyrTwHAH5fppRt7jOpx6i1gaKrNcFNQYjAohUy/s9Z02mv8ZdWuPTJovV3OeXJfFv0lC
KbasYu9Cuhz8RdcR8WnV8LUq5pR1IDhJ0TizIi4/AizpsAF4pKcTLv0D2zEfjpgJUUO9sH7/boPA
HnHmH9NNVZkfVphy+eIkR8zsi69AdGx1NwqnJqHMIf1zNiKuRxnZrdt3UPrYkt3HO74BGrkhW3FZ
W8sGHhLjr9FZ5XjkvwVAVzsE1Zp8lRma7A8Fd91Jp+aSisE/fFOVlgOltNuvl4m9k2RSKzjt3+Ll
zpCi3O++yeQmot35j6F4QahoEofoU5++BwwF9MRykYaFGvkrw+Rve4oFzToX4JBnS8foLiZxesFE
KplaV2E4ia7A93ZAuO3YaUQiuKmruH8QXNq52WYxw/wGcQ/ZNMe8CxDkE2+K3XXcn/yEc8qI6135
swPYUqkUjwmUjWmmwBu2CeNJuen7CLvf0QrdJRoWFBRHxGvvj5kXcGPGv+hDB4NNy0mHhKQsOzSl
yWCvq/U1UHGP7QbgrZwIL6W56Eo8DvyY2bIvdNM8zoeYI8jhY0sdCaMW+HF8/zdec+owD64JgW79
ntIKxsVHVUfsbuBfoujigkUcj75XpNsODmRCRfrAxW7PmXLIz8kvqY5bYwWg4W9EfT2o9c479x+l
Lg780316tklRAIwTuxNezaCo63SPdfcnsZQ6abpnjb8LRoVu5laR7IRpYNJygegBseVPnF0ONkDE
tzN1aXaqj0Fr1ZkeuUuCqNb7BKCvqhd6VLp4K9jO7NgSWdKR5VNZC++tnv73ZZ+7YI94P2z0cflD
PL015dURUMJTwrvo9xVt2dzhAZSoPkbKeYjLmVyCqT8KIQdA6GuFpPj/hP2bCJ52ELsGSqRWRH/a
f5bZRNq3hFczfpVur3j3ijlrQ5Fgf0eefMEV1g/K4e2abXczkiKBVdd5gnv4Kf0HUUsNU8VeE5Y1
qnVzIS0IavP1PcZQXcYAb4t1VEtcmG3R2GTEuqGMmVj8edWJbsxcgh7SXWqacovsInbXgSMiXm8z
gvU0cZA+3MfXewrRKWxc/m80frDg24rqcBBNmOQDanFjDTvtrYRMMaz2lQCUFsawAFZt+3+aw4MZ
W+yYdnqPt6Y/PpYZyV5Et6+Ir2lzuU+ERX+oZKEyAvS2PwYkl9DDgWcmGk2aaGZGixzUUGK3otiA
lJUeTHvQXN63+dTVC/jLVF6V7lAWkVdm6hn2WNs9yc8yPNp0mcPhPaiHs05P/YG2IvncSqA1Ercl
z96/chi89jnU4ToZYplxemrPLjHJaX4Sah1WOnUwJxwUCrW5+C3nY/U3omDa9sIQ5kboznd+INkF
l5ERyrg9PpJUX0trfMWyb8DPQquNBbGJAFP/4Y8j1WIaMLbUzSNxshLGRsRPpAqv/hNSydXAvK/H
+oNy1KwWhWCP0Ubpw4W/K567CGFECglofT21VUAogQTvaSs9ZXFSZ3n8Wy83gb5mptHPd7GpvBAq
aLb17fsJrfpq6mmnTWT0ebyAy+8eNY1vrVHPaM07L3V36HW1BqN9Q95ESv4czm6UD0EtJ49TVMnk
FRSZdAD4MB1ta1qsHQVgfq0EvrmGUE6MtqOxUtYaGLinKDO8LEhnSS/tH+XDrT81gNK+PD83ZsPi
fGpVLW8kTJxzQlZCDB0WSp3lGnv548GZ0kTx77RasAfyCNwS8f9yZhfDS291zLp4YN/YUn/BlB8t
Aa/ITbkC2OrveAwXbtYOv2YWWuV2cDnUurlAGsI/zi0fGXTDeA3hhYVywmNKkG1JFCr3Lly7MWqf
xhSZ2r1xiQonkhfhl8e+EZV+FoVsVEp7OU1cMpj34iAdgsXDBFPbVSDwJXe7kisacl5fCtV2Z9UH
idQa5g/Gf07rB5SkIKDvZ/go352XypS4jAMYvuKZwP+ENf9ge+0utPRY5uGuVVYZQS3tGdth+88t
8rl3UgHTPt+jE1fq4ui7k2ypRFMf92MVlD72huIYoFD06ijdJ1PqR1Sqiu86KSuB278BB++BbatV
RJT4uATfwsDmLdY7LwoU+2zIQAnh41Lsgmt38CwTcZ3+s5tyw3QQ16JjDkBx9rwhO2jcBWJSFhFj
GVOpwSkQ3zMF7zDxj6pyZgWww/jfWtxYrCwQC/8wTlEZCDJsnLT5z3wngq6L+Z1oCrn3sU2UfOr3
bs+R/GClRC/Ig+ImmDxQDr2Z2eEdj6INg+6heKX3kXutqaYKhIdR7MFOQSF+7GU7Lg6mzLMOwIx/
il9lc0gFtdfXYldtHQ+NR/w4g/EeGAJ/t2ur7XbKMOKoEWl8jMElHbE6B85u0/mlCCw92ryj01AC
YyUSRAwBAx/uf+pc2ScZJu1z+UYoCbZgn+lY5gsLkbg6QR0/X5I0w7g67DoN+YM+ZoSq1Mh8Cz7C
T7SNApGOnOPpCeqcSk1wUWBZ+vnZBVOplA/tTkjcgKPM/kOzlGSaSx5FoJ4JmaeeE6nHZt3lSK4Z
qWDIpXCs2SJJRtmSB94t2sxICRuj710Vp3yBpHxDpFr5NEtC2tCtlKpYE4Y0yoo3rpEuo+fukfjW
lOQAoJxVKDcI04T9hCRiLc4/Zc4MMPY4lKyIZKGss3qFDGxqun7SHpb4J6msh+p6JGZck82M8qAz
nzchHkU8X2IFJQpsbpg8akrtb660VcQiZfruSzTO90CPT450V4y+sgKAWW5cuL9gUCY+DnTN+vf/
ZLPi+buF4YlzawTkEX18I4p9hFvy61XFbBF8SQLgYLHfoz4GYruygeRo0QdbcRLfsUJRsbr3/Z0+
aScVeatq8fUtNDQa8lPVmcOnvbvPxI3KMTAm8+zzOAfPbAD54UwumI/A7qWwF/23DOkKmw0nFxyE
39T6WpAYfsgRlimFYlavR3NpJae1U3H98J7l+d+USFeceXEiardsQd5k+uQH/n3nt+PZfF6NxHif
Y3UwuJxJYYYwcA2L+Z9VkQ25QnpmrY2Hfjh00ZKYaY9wmUZ78eWQL9FQYFX/rlytyt6vcvJlqT4G
dEBv4epWPZDGX4QyQGcnofjxHWYI0HOBJABk6NLqJ2DSMd1yY5ED1o5WMQslzIAU4/Cez0+88Nkn
0q2qEwlZpoI+CcAG5bNJuCZ6V5S4tnqusctC+SrOPPoCZcvAVuwu34L4nfQTHM9z8HZrRZi2W6nc
mvtquSnTqKDvI4LjYwsUQkioSESKWq4gYQXMQsiZqBUFztNiNfoRMFOc6ZruOOQlO1mA2QrhIWmt
mukxtLjLprHmK4OcIsGVoQ9kmMZ/5k+nEMwUcgCOFMLkGft6qjVsr1tt0Mi2RFhyqvOCmMcht1sS
L9NRkw9fC/tU8B8/ZmEL9m1Kd2ir9SCd11VT1kQxe/UWHdNw6LJcA5d9cmj2jlU75QKG59F5XAvF
X76v4PHhg2I/gK+JMBz4wqlykeIVSX1FC+5KYYsWIG21QeG0xUt1CA6dAWJP3V4iwbW7xMcEvsRh
S95W58P/zqEXaVSeAKojO9BXQhXO4eWzsA8vDgSlUuzgUDB6TFJdwSrOyxXdqoJRwBiFFAS25K9J
Lm33cKyAaCCHiiiG3/pY7Cc2xyM1EiI4E54Nzsfoq57kjtr68dbkmbXTieQr3Zt5nAYRPYTMhPuM
R+Stbc03VFJkY2YstR4CytE+jyAs+n2Umwh+/oqFI3IBnKJUFA8sv52rRPGswGbmt6xS/8e9WpW8
BOytGqckphpv0qGHJo+SJxEJWWNuz2Wfvd+vTJYOHik1Bw+EPRkCIo21ZiTeYWSn7tkaSgVBWJWN
vvG0bwwYdRnDUOrbGhTm5p7ZmkKCGtKuPd1JGsrCJLlFE69YLbpbOULQn/XvkMUHv4tNEVmQZ1fW
JmG9sikgBmoKuSVw4NqRTkjmwWu+1d7yJakjEThu7GqeHrMt/QgH42QH+Ay9vrsC2b4THbaP1S3O
j3+k4sVG6GwbCoTpqHt4PTD+LFLx/bkJVjio4bH7KVoiwDfosmDgjCvHBxlNwN3Y96sqYaiA40bc
z4MWpUWpCudRamwzse2LdLLonngvn7oXCvko11gcSv783DqvR0Z6lOEwFwrXEqzOru4kyuI9ZGS/
1nNnIc/l37h5ryR9WutzIgdWRjOPp9FZGYnT5GH1UakWElsVul6hK4LYSxDDxNA1p1kiGnYzTash
z+gXMbG3Smf/567OdFYZ+pYEuUnzL7ZVVtXCXPC2wqai62YaLU6L3k9WeaJKVHf+8hnRy1nAEmf3
DrHKnx2PYaJKZp99U6KC0nhTsJo1ngM7uTWe215wbGS6fNA7bnKIvOhRMD/l+VxnutI3a9OF4BKB
XqABMOuOgHRfNXw5LHHGf1BUdGGrT80/j+s6yVNXD9YqovwUS+vGAGfvsn+la4iHnHPWVmAl7DkD
8oUCghqGV8OaEnTuHXHOayC87nZz26PvsSb/i9NU5j3dEpGyy4+Qu34sQ30FhXUTsFWD4GJI5MoO
x4UAAbcQBdXhevwXuDz+KijMjMKaGEmYNIh4h3Hw/iuw2Mr29BIuQy+/ZekQz5y3c1yKsAftAyL8
CgzGhYSdoBdAbezfATcBh6OH2cG3jggefvYVteQcTWwyFW7/Na5GXF42czkK0/OIbN2LPiF9k3vv
0chudhekIEV33qdDJ9+3WH3BOAgunLDUAvSaTKLvG8et3s2Lij0HWVV0eG8S+XVtKmr1yCCPl/oy
Ovu/7BHctie/63XbVPvxq5OFaPL7QHQj/5g3jRIc4066jYjqxK16jxmt3X2lspiGs1GH2KrBms+2
Wjz8l7aXsm49OLppHjE4+9gaDCTFxtUmbaoS+asr2g+Mr3glMhH//Ni8V9YQkpbAaRJrQy52iAWb
/VVJXyh90jyMtAeemXwmNxqJzN5o6sOKtIoL5c0zPT/lHiOEZ96+FeKEPMFKkeRgPb3CAONiwWiP
ZftfMLqYkur2fXpN8z2mXHOuuCFhOHZu6PzTwtzfrkRiCj9CVBgbzQCGHLsNHdmc7xin8uFByA2P
zCe+1eh9asvB0S2nHq2zB/E8fNrBhnkNE6RBzbhtCjsYAqY6hAfR2AwDpuo6uVkclRllDkK/Tr4Q
s2khrVkvM2rN52/oR7qsnEGLgI1HluAnyLeBa0SyYXbuYwSF1RBZEt2DYo/fkJaz36Ji7CPFaoqW
VtZMLBhMTsMqC3ZBrOx/3r/5QjaHazWzVg590Oxwfzv0ApP+0xIq+J5Nzm56CnXdLPRMglkJZ6Rv
4TwRuTL6lcYtEuECnECpYwxqP+weERm2GTTXUa2+xBI4lIIv2sAiICXcqvcx8yF6LtxBORWihmuC
7183m9+gWHZHqzZobYT9A2qSDy4nLpv7SCw8wzOYn9oYhkkT1C/syGvzwq9tIF0MhRzXuNQC2rW4
gMbBrPTBEVw+Q61LurAuaukAoWAqx/qmr4hj/2y0AsWS8ZwBB2nU9IFPgQzg5dz1TErNmvDjznBG
VWdFYqd4Defo6RlFwE6/p/pvMHuuhfcQU1++pomw6GIDt2YxKegXs1fonr1jgpQrTB5CAM/dCRnr
keWukBv0Q5v6YgZysbcmvX/ziPBFQ7V79zohS5ag5GlVxd2K6GiJ4rOAZVX8nrod1yz5dcH/s9mm
axTdvKzabklPw9+l47+kOIqSMsU7n/NhpV8pp8wFdGwsOmXGVuWHQPTvkf3tndh8nE60RCo3i+5X
1fLS5vZQ2IH+cWg+rZkOFNVn1eqJcAjN6D1PNcMKjeS2mdH4sZ+/zzvYyxXNcA+/KAzNtwcmYzk2
nveG9Fh6LdjPMYrHNlw9JWqUAdQiKgEWOnx2NWxSI3Zqh2i+Sc+pRnyfSSuPU6ZsdEbBellHL+5x
WaRzuAxQeobBpfyJNHhROEZSMYxQVqKS5/TozDaFz4ZOyvOlp2q7g1BlpXEf1sZWE1m21nOtlqUx
l4f61g2OM0HDiW064qDKXmYha6Ra06uOFrUjqPC9jnSnXcTJb4ZUjkDUTjfyjS+6HTkniyE8nJFX
awObQ9I0l7eTQuHkfLjIWyQcGP3RuCVHt6TRNLZe48dWEZxeEgbsjoQkZDpxBmmkmfgWvRxdin+T
gUcvSoGNKF2bPrPFP8lLhzl+Id76m+tJhc+3fOsBEP4B6Oo+hNscPi/h8EjDycGPyuMTtnlw0LBn
416RDSK+bNMbJjR4f3RcKTzVBlY/O8rgArSdrEAHPVmVh1yAIdHTzJH7JRp1m2nsBpziqpKYGXor
tUPIJ0o1zg3V3dIhpAupIo8BIp2Xzq61mc+USaDFFnspJsZo6paYIEmgY1MibqH5ib9q4T9gRkOs
74lrJKFWlIJa4jcbGOkwhFlRelTydGrUZujnxD7pA/W8MBrenuU3ZOWLB9N1GBchzG3jXGnsmdAb
1gIRV/R4Y05Znku/DkX0wBwn5ENImS9fbcGg3wRBUqyq8vgogDJPImNX9aNYQ1uLI80cJCxfSjJl
rxx9fqXqwINxzD0T66vy3UVxdULc8PF2clH+exiZIyA6oiS3Fbg6jleAcecOjIgurnxblcwUfO7P
9ke8AL4bPRrZjbWSMfkOKc86hV6SC4hvdN93ozwwXKkesMBJjT7o0UDordkHtZI4cIXTaqS9sq8a
cPHY82oz4RonJE4rpIyDfbZXTK/3DK7r7CovT6vu/QBCKokzf2fsYCH/GAzvJHxVRKokSmeAr3ei
8wzetkOq540KJFylJ2Q1TPsJblJ1i+UiJqSWyWXtZSTAtSraojF3uJYp2eh6sZo3hbCH2105X1Up
c6HjzzOZ1KBKM52tiKdadzUjb5JJJCeE8mCmz2Wi1k91sqxyRvf5YP1m4jjFJbz92l6K+S56uMZu
ABSBaRedLrtSLwyTzauFcmw+k69nlPz/8Nfe/QWbWEyt8rfdbaG/7mOTxaPQhIddmv6mc/sLX5G2
yrjNwk8A5o50Al1udLc3RDBPwKhnTTM/gKg97Q0rzWp+PNpy0Qt7c5cETn6aEnmjflARz5kSOFAe
yvDtZ3P1Ev1vDLQ7v9WCUbOA62v/5Nci8OSh/mzxwP6G2SUw1zGVt5TG+dahQc/CY478YSARO8/3
k8c8ucT5U6NsLm5ONhIRwrEycOGODVs9U1xWxCdr/XzcRGWMXgtA9nxWZSQl/iYXww1yncZNVdPF
WE9y231MXtK2EEu7CvTDP4Lbv8CNFhnutqJkN0cPptW1opxgkARR2FamTaSseahxsbTx4W+wJxVR
QiNVFIk/ZcQPVrZlwc1sLvMQwa1SZpNhbHZG9tjfLvh/55Mh2F74m5MgTNfCERarK5nrc+u3SLZe
+9LhdIQTBfVkC7ZoOO4HWQHUloEYvfbOAzbFwQn61qDNLISDqO5VjotDhM+eqM2uvPfa8JDRgc0C
N77z/geYV9ASc3jf0ZmxxKGwyPj78capZEQp2/Y80phc9meWjRclITcfxBGHVWHTaVrG1R4fNG83
vq1WERGFXFw2LuNiNYkmR0Os4P7UhqiDHDTJiy67EyLVDGMq6Cj0nZiU4pkC0WKiI3RPVc6nrweR
Ony2B1+RknWSL7pCJtCrSev4qW5xaSJTqvzSy14Z+aZsdAW/WrnQukjRJEQ74E6eORKJxlNaNZy2
FrY2lQJlCosZ/NCAvM4gALzDFjpWMdACo03tf/rZmm98IxkNJSEmB7MkCbnL2ozMUWX8kiblaHeD
old421k2sStYlmG/4KCrasvcGy869O8NUUmFh5bdD16nwInPtXv8/neh7uPYPkBIUAFR1JZ+ggDv
8MdISYR11UOj7hubpe9vcVWxFr3dVgPD05kW9biqba50qe1hvdShnjNMkfGrhK2BrYahzlwFwOMR
eReW/oGhNMyLQNT+KP8rltIhWmLw3gzJnKp8cVQRM5by/YP/GqbU1EPV6PAGwQtg81C+pWj4Mnxv
TCmfHTR9/V2bBfBgN6tIf6LLQmZ8gJ+tCWzLYx5Y111HoOJqtnhM+5/RRXAJ+/CwejEmadBTPYxx
sXCfqcZvJRynX/DoQfai1KOuabDjyFVhKweYFISoO8hzQDhOQ9Mwlc2wh76r0tbidbCkSFDagZEN
ILTzVl14q8yc0v7wFgXsJ+oEn7ILK3bwQi/WKBwfZDbjSpAEOHaJ0/5RmKRa53NOIqjOEwBmk/0D
0i8Y/SsH9fv7nYkoh2e7fckoqzIeeDrldla0uBIEHMSMNWgFGh87Zua3orjWfAP5+h881qZCHDUB
3OthklJEDcg9QHwwEwNZchhhFeBhbGMJeRoXYEUyS9WAap6nlPomP0FDX2U7WJ1vYhk+CyE+HrU3
C8pVPgti0l8Y8Wwqw572Y0JqivNInwazAhDnGBmv4EUx4hssBHLiXbasUtfnkEsyprqWi8+VL0Tn
BPE5NCwA1cisG9CY22HjMc0BK+6TnfgYdxUHKbglHxIjdsWVmweW3Ql7GZeFpXQ4qrJOfUCY2D1E
5PclplQNAzM2NxbFDFFDUGKfn3T8M7ZD5p7HC3bcrSo1+c2Tt2Zmf+5ONjRQJGmVq+19VnuxoBV/
z2W4KXMmvGmmtrlAHjWvdtcCkJRlq66TENqud+bc5LsStA6xWUDRC7NDJc2E9l/NL4vZ7jbaEW+U
K3T5Q0IOrzHVb17DbmCWm+l1gC+26ZwCEHMy9/zmDjzKlUIPSWT3RrwreepsnNWwwWY5/XEdOCWx
yqMbSiFOmbFXtkMyzGlDqrIUa6vOvsD5U/qwh69z2bw7sM7rp+oEFX3EbLuadjNgN+aBl+9ywbOM
6t35F+kkkTV+rShvhmEXxvLbiXMFzEjGNEcmKvzzbyjRiEU2sVZ3Mj/mHcF6bmSCICF+IF++tR82
X1IKZzj2UMQh6AkW4jBhxmrZ+Z7qc+5wRPj3NPDMDYVH1YfG7E+9+OrZyCIVDXBZQNu3iHJxjeQG
+Z/zHL0x+tid9OiNcHisYsCuTzT5lcPEAnTdNMFqiuxBrpcWyf1lIbCkw3PkBowdNXaE64XiHyow
qmBxSoh9aIWPxFsQZmew5x+G25CGef2LPnQeoQ7rFS00Fa7Zi1sugA7RcbE3JxwEXvKxIt9uMEB7
3fYIPGBN1A+Vdw+1M/N8IX6vdRPPQLDXE7gwHfSXvotr9ddNSr/wu80MjcCLm6Qk0dXPg8uDzwqF
jJPLUUbESk8IfgkTt+A1kDx6rr2OgAKA1+IyAL4kQMdYLPV7W4Q6NF/7iX2WxuH+oqnQM9xI3JU1
iCwNw54Oi76NSifgSrAzBqUrGsr6WNYebL9YRfUz+ee9G+RVtu7zGUY3TIyKN72g6+idLSvT52Mb
gIeozMp/XCpEeKm5m8KutZzJR4QbRB9pZen0JBmav0mugBB7L/2zSb5YBIvRyWrUASrzDXJ9ahEh
3aJh1nrdE6Kape/MPIWwLfCGdUBfWJyA1gTEOdjNebl8OkeESV9eLn73CEy4ob6ClUvdBQN2N0tM
T3g9hMetSyanG1irD/hznSIRne1I62k072xtTOyicdq2d2DVODf88eX9BBMOE4m5vOPWvyQPVSDG
gyskk2hbpyDqRD5KNfxiVvPs744uf3HXzexhZjZyzclm7TtUnK7i4xGRiBzpBAulrB/p7gY+z0mQ
rmvjUKdvINnrGWIW1dllo07Xfb1BQXo9W0jLJDTMrrTbGDG16eVVPkFbLI4mZ6w6/j/HsTXJv3LT
A7WKPux0EOSgLsy5ORxDwldJFSAHhkwItvdj4YQoxjw146b6Kd1T+Sy0Dz7a7B7rrKsUCv7z95ri
/IuZmcQTb+Vxguz3QOYKuaDC2Zi5QQLTcesuGB1/E9KOuTC+YV5mBaOT083vWF9n61lWElilcS/A
dldqD9B0mRl5lLr++cwPIQccUmwPfYo5z3UXT7NBzVdWkhwnx2N54YsCDioPokbQotWND/ni4uCP
N+F5JZ2eXfD6vvkYGMO9zYoG8igrBrArl1hBCyh0ZEN++jXlYBj/jd7oUueIoN2zYYs092aBvuTg
OLzaL/kXZHh4WkLF9eW0nhm/dh83zqw1QW0vcI7CwtOz7vwE5oAj7U3pxYOslIp1xcMYdBRelZb/
XbziCabINZ39dc8w9bO3UsLlUtpDJdaTVRu27YMYRfpbpX2qTBl+Fkr5DQrHddbVgePnPPBZ/55z
Rb2qboYroNUrwqA4vZDpHjCSDKG1wf9ehN9XzRC3Lxvk46yMhxW1JAPVQfpc+JwnNV9DjfkTsOSW
OrhoCOhP5y0vdwCI51QhM/8labOVkRHc6mu/+jvIiWP2U2SHi15wiII50QuUhT1A14tSddtodnLB
th2iafqBOqsHKTzsL94IO2QHIqS9qEEsj8xQWT4tcap5nzmqcWoQnbrLVE3W0cMLvhF5o1SbXND5
W6wu023EiiXKrof4Iy+FB1+Y11EogaVEvfeCgaq97DNRDsxDHM7CrijpwB03SvB/zDOo6TXZ+Bkm
ofGJck+ZuJ4SD+31Fd8F/VaLB1VQN3I0wVENG//m4Uw9q5u1cwTFKxevS9m7v0/rj5wxHuUKxl2j
M1Ma8LVMjrEYrpIlbO6A/XWVVqpmktJdbWRmpBJggFoHUPJwv5kVtXDfpfNj5bELIvodtC9m0tiZ
loY8j4aGdX09DwsJP0x3EA4bimKHPpc3NKUsrtTpBi4jq9QHohcVMjgb01lppJJabdJ/FDloxqyA
EyqlpNiwPn1aO66h4D/5rdUfhiL7cnAlBNy3SXdCckIFBYMTVIRGLSYD444wa9foEKCs+5Z4Ubcn
3yAgCPYttPS/YKTiNxtKhJd15t2OtJvRT2bEP7yoxTcNpon/ARe/lc9NtDxMZtB4jab2TuzJxpkW
BvxYeTDFmIRJGGSK18v8Qcvc898ALtIKmrahm3RUBUjIsnB+IHX5tTBHV//cM6+bl+0I69Ub4jjr
xkpX456u2qBl0i2W3CvJ+BUOwUc7HsnxlCCqN9fOpgA7kjb1atTESKcCPXfGD+YndcznRSQNby1f
Qn/L17inF9hsU2FEQ4oVQNFZ738cuYT+1G9aHJW53bGODdxGJ1HKMNR01CHsWGcKQcylCf2P08CK
P105QSN0UbfLWgdQd4IXHiSAVBzmnrxXuMJSJQTJfdEPH9dzQ4Bj3sNjjhVX4sjqlxnCRUFUO4sl
ARdNpmFhvrtuvlcyV70Xl30KfKqPDlVPwmbnlFmsX097pXlbpqk7mPybCzrLUvwrw7PX/DKCoBlo
/64VP3lSw7hflXXDh1SByaYW7M+1SxemJgTtNyOpm4M/UaNWDimwldjZ8oDuShdlf+lR7fhKYP4G
ccbdwkOi9T8rI6tn9z5yYPC5kKOJVwupA5CEICLOXTvJ5/xRqQ3F1ajklpgB3Fc8f5e71+vXAxgL
YLid0CCY8A8U/aPVfFR6U6rr+hQMGiepTSFxMnwnq3lgdHcmVf6a5POOOcUdrH7RAuiZRox4E0RB
GVERGMzofwNptqqiq/PYNfCFwRW8+eLGAkHVdOdl2B4Kzz7tehdy6g+3jR1Kvx1/B1PVVDeE1/zv
ys2wynkS6aUw4H68jGDS2gCffRmV9BX/eDLEPzTngcYU3RGzlQvtuXlU2UBl347V+ifRo9zU8yRa
NOj5lI1WIvq4DdQ4ZFObnOGfT3IG6OKpSTvKINEtLGzGXcn7e4RWi4G6Pr2ca2yK5/nKEIdci3af
iTk1GFtNiH/KZYD6OymJq/7JWVFO/owft9Bte3SnUv43AfCMtZzDlGKghy1KvFs1q+ea0kDqB178
VqXxIq/sNp2/OclxAadnSpazjW7MJfA0S/rH8QDokdyywG7mNBtXrzVI9fUomypwj1uie5QzSnQZ
ekBBxji9ay0VDWJjaNQb+zbB4yynqWHF3UJ3qrY07CgS6+NpsZiNTzr4jt9QS7eNG7uUPdEWivsA
frL57dwWWMcu457IP/gSEOlcNAhdMsDCViIF00+fBvkCluiMMRVbdISoSmzqlVj4IfQzBIOp0HTB
98RiO2ZQqTuPLIR9T9V/u1IlZkZhRsPRA/T5rd67z7FqMAcuBJcPrzhKhXvqJZR7mnEmZ53sx7DF
BVl+ZQLfP1vDQgA5PlczQYsWGFjjph+SlNJxIrbF6rR+LyarcD9UrfVKKEYCVYXf36yobu3HcRAp
rcjAcghMzlGkxad/IIsbqeRIkC3bCdGvVUjLfXl0PuqSpfvgOkJFawC81vyogjWGZjZnkfPqM8Yy
qkl6Wh3sM9KAcQ3n71eLgsO/SAEIlSrvGDZrj4QNWoxN7Djh3fUwiGcsDGVRBrj6yr+sd2Pk/KoN
04Iwtejn4vTzQ/qggL1+sk61dKrcYbWCjp+4MRvCrSu0Wl/vtyS0NIrfqAQqbTYhRYG8VGANpq29
HxiRPq2zyGDOR/JGGof93PZxps8lc+lL5QYp8XLs7WNL7CD7u1JRAiMuJlq167nKnj7wYO6DtBTI
xf2wYrwiFARakvv6Q9f4/fCJMoPnf99QsXHA0jSlfHWCrEKeH5Xb1g4vijrDgfsWHll+K3Qu1AHH
Jh8EHbhi74QWqoLdynYRiEh1HpUqoAhV6R8E5p76dEFv+CNOuRVtqID2iKHlSRCQihihVweBBAkJ
B+hDBqNbjYd8bB9ojEIZjcKYWKaPk/PMRPrfY5Iq76O78dp1x7zrtrR4NiCWybTHq68JY4gkpLBT
3MvTn2y2WAfFmr5/Z0ZLntcJB0heZuMRriR64+MFnkrJ04Pc75/pKoudcpgSoVq9ufRRORbNoKfX
g67vbXYIWQO0vYkVgOdMCLVHDxTVvLnBI51+D/mti4u1AP47w19ynaRedvjsGuwzz3udVlPQUnrH
4yCpmDkbDPk5PnqLVqJP9jDx10911DVbTvnS5ozFzNv4fZama1g2mhKLhY45xzqnmmAOuVOnsc+X
YCfU5Yks27TTrkGrmkUQ5D5IGvethu2oW5lM4A4lFTG5LwyWQv42WxvM16MyyEOF7w5+jOWivrOH
MBk4FKgsfVimw1KC0GSxfl37fKoGtfzqQjnkqopDZZLFR3WG1ioWdrN65qp+V+P/KNBBpKfdtdu5
Dq525qVUL3R/UWpDsdSMvyHHsDGYG/Y9NqnwhcOsypwTcccc5CyF/CrdyXW53c+3L3RktF5gtxlt
5Kw8DUvwkEBO1hxd+oLc3FpSGpCiuRiATN0ZJ/WeeT8XXVkGBIdAZ7mel4eWrLAYs4+PxQGBZBGe
myziGTFrfC3rp6Fz46Ej9ls6+G8AXMiVNTTG0GQgdp3MiKurjqlK54giJhuxrDGu5oO6pSifW7wq
L5unzSofLtqYcAqUcgKM2XcPXKk1U9PKddSqu/hrYrcnL6wUkEuYaJlm/C4vzl75E90bNJ1OLnqB
FUWnBNvOLpKqJfikZghY9NfLflVbg3dorm4lTOHge6xfsOWrDx5Cb99z/V/V28VdifAhPqvHlj+o
OkqslKtaw5sXsXO6SLs12nih9/uGd9vFzInRax0DtTIcxYw0tFbsLhdqs5zLfKDlrO2Vgr/yME/W
zvYmrViKPO+7mFQcFC76hidMenVMNNv6fsVLMSGFu7RXfVu5qKHJr7pOh/LPyWsZqy1EqcN7gON3
4RxiQcOn2xwU0O2VyzVhV/afYq4eZe4AoXAhG7XJ4Bqdk46yZeQnspQ6pLizINHKImKW8zr4pj4+
YHhoMXoJ9siaxANi9C0hw5iGMfptstwbTvdkUc3RwqM7wNn9SDnhdKuMPC2HdSlsl07xdygDOk81
+l9GE7z2B3Vd1YF4pGnDvPze0PNow9g3q8L+z7mEfvSuqUfAa33wnEQGcfl3/PTUpMKIcdXtQwSr
sQLE2jNEj3h2lNPov+tCbVZ9XZnht3FP/AThlf+iYBfbUC8nkSukBDI5ByZQ+MH1Scott7V+YTFk
ISaaHA1N9Bvkxde80MmWO/R107zA/337gZ1ieWiZFrq/DQQnBR1KSg31UYSeAGIz3HO/QZIweztp
Y/8yeXFgXjfUMtypH5H+87gF1nExhExjHRgWeEdtnfXLGpkoARBgTyqZ0fdST/2L3RXjGl4LMFKi
//h7T+Dd8ZG/pHR5sE6hUhI88OGYKt0uoojwsqku9uEDgCKv4S9FCHaU5f/kdwLVPaEGElCAjfX2
ZlAqskyH56zonwEedLYg/KVHP2svduOJgUr0mW5AEkYTMB6ALwyaeM+Xd8v1AAG9a+NuEUmCGdxH
XUWZ3X0EGJSEYmIlSQFfmY+oyJSu0H5Yux37Hfq9fe7iVnScIK80Np7blaVwXecwmHuIooJBrZRe
uzzPjJQWslphLjXAtdcnqnIOv8E44TNUoxNQUuTVHmZCeEdgp/xft3BZHgIFKf95O1nGaCt+91wN
YQxv+NPp+vjc19DgZ52E37TUX+h3C/ZtCEpJ2Z+qxiETmqfzN6HpFGshTVrxhKGtiDDycyhYlE0e
ht8BJBYxGGnZUmtrhC2fL2TkVj1qKTsEbVNKhDNsMh/498tS0+wHpSvCDOvPrCTlsaE3+yRo/q+y
R9q9o2cY8XW2AlRmylcptyDm1d/UBTJMFjoCb5Dmq5D5v5kJ+jTRj6PuDWt3+nMi4Jc1A0IS+8y+
I7wQPhhd6hDhAh/sWtLDarfAUwE26DfwDCsDSKaPyJS4+vOktfzL6Xyxp60lh1EZTkY86kYxPrFP
PSQ/Sr3iPskyhCPxmQDdMwJL9XgtY49wTR/A5mzZYMdKX2zh2ZXP2n907eqeQhmFlH1vdnZ8I8u6
EqSTI2mfokF2Q6zOMBdtwzrUdQqUooHdYhCsre76Uc9YevxaaveiQoULQyG6cCZ9mN3xugN0JkPu
7DNdSQPCFeKVGhQ7L3uL/StHlG6FSYD84v0NsT6shWoflAPE3yUtKE9SKO2QW8wx2yseFvOQf6jA
rTU0XR5DMp16l/cZpG6f2JO36Y2XElkLyW36SIVr13J6aksVTn31e0/jzXENqLIw4ToBGC8+eNaL
CX25ZGN8e/wfa62k1cikONJW8EXVe0PvgvFPYKqHpjlLB/+nYjVL8AdZJI8959tQUyrBlJLnGIWA
/fLvg7TKDpC/wRkhfffx/BPd07rld/zwzWPll2AuI0Jit9MTR05Qi///7NnDGxX6GzQdd8IGS4DP
vI6vm73knXcCJTM/EDAgi2yuy21f8gEEetBOanh6zZkGCjRH608DpKu6dJYUENKDGvexcyOmchk4
zXWpdvQQoVXvxVC5zicgsviqGwb8oNbxMgGcdbVy9vfsvtX5tKFM9tdZHLuKnR0QGaQYbJRYxPf7
lo+Qu3xZR9C3/4qG4O8R23tb9SGphJvh3/CT05dCyFgSK6N8MRoIK+RB9DJE8iplZGQNL9bTEtdB
0moW2e8EOHeUxV5f5PlGvecUvKLTGX4FmtR7/I3v4/yXKHGQ7HUt6rldSXRMoUgQI0xNfwWkq38m
wNZjXRC6AZX+KVQEIbOMd+w6/EMTAkhFExcjyC2MF9PCcwCIbu8FicFrVfdb6B12GEIEiZn/yg5c
f+0PDvtDM0mQJ9nGOcL3ETsjmFDBeuZLcWAqQMuHlsCflrtk3wJyRmNMejt0dpGkR0ayH9pAYcDn
L954KENVAVfOrev7GmUNlmIjrJS+NFSkKEmbN5hZNHP69gIvuZjRfJvyEa2KbYnC8XbeTgiamesv
ao2V3cToy0sUsCQHxrkXRpPzuhIau0ib7KbFI2Cuf2ZP1DDrureDvSpJ3dzYZRsJimvwsaSE51zw
79jSSysuRVJZ3aCDCVTEgkI9F5hQsUxYR29Rc5+/l+9KIiqRFOilX4DUA3IkWdKfr/4SW2/JJpMU
JcvC/wOAvEqRneMXbY65PwOgRB0aRS12wKSyIj3hzBvj75HG3UwxZiJqTuy3nsHny4AKo8d3bTsZ
SKjmid2Nz3OmENcIG1p/dYAO9j/oItEMsJkn5NRfcGRrN0sKbjRMwA24Zxiu2mYGigbXVYBKjleU
58WvBN+w8rGhIsdpYC0PgneCviDkSZfx9tqKQoDWvzr2AXjKO+qhZtgTXdfRwBXYW8ZaceTm52WM
JTWUwHMr1AhIjLPmOiH3lmrdwDngCIDBPibccFh1lebywWEt09fsG2sQvEU8GsniTiAKnaTDxMcS
Sqye3mKlv6l3G4dVzyCM8ir2w3Qo0p5LM49khan3vmhtOHESs3PJU8ZKBA1iQzxY6iytnXNgR4e2
U3nFjJpCM1VWmG9xzIUjkvpLIHT0OTgc1C/8lSSjpf74Ma2bjqYkBj7K9NPayUNUacAozSOvsw9x
capC2seRod7LIxA+SPQUtWKS57zq7F1eGqq9cSh7La5Chb2hi8B36a4bDDM0cDifv7EkCrlytrXP
9j2ROA30ahlTBDe7kwskJLYNTmfBKg1Qk0W/92iRsAGrP65aGp+FaMUuuhnhcrRAH+tImJXCBbAF
StsUDaBXIRXGEdQIPxnEoh04Eu5VEyICyHbGJpRxXjHsSIKzd4K+O6p3v3zkROmVNf+ek8LtU5c9
ZdVxEyNWdP41M8nw167sW5FT/cyPich4HG5Hjd4bFtrgl1Jz7VVcvZ/A55uw9xTQAZbS2s5h1owA
n7SIaQhzYzZbnqkxpE2kHD54IbnIZikZWwug27V2r+bZEK8a3wDqVt/zgU+ik7t4AFRXlRczlXRI
QPZEezcNRQzQ8HyeDScd+XL4EmrMgjeEhIFKaAzPXva95/Ix6yD9abSe6d6K6SbYHaxHjr9m4T54
Cu6U2FAI+AZR+rsfVoHMkou0/6aj0MaSG6iKeUGZObRX1p+32mnjt7lqigdGGeWo+R9jmA5XmMKl
Qs75RO5o+mfqepcg5mRO5Kti6eFQQNBDipiVQHlf7pvK9IobMiy6WURZN8FyljPVTAkxrhHApqcR
gpB1qUW/3dStVyOOOE3RvWVCNh1k28SM67jbRRqMVYTiWqQI0WyIaFS0NcGFs8JPA4Keh4MeVj0k
P9eW3e5e/wV+IDB5uSYnRHlid3iMK/yOuFj1AzAZUZ9Qqo3frQZEM1AL9QSl47wxgS67+VKDGC3c
4UN66tKtWSEbcAMrh9/8qqOz3G+qISAqYq6a5NTYSd3Q7jVyrncFctpEoR3YRKYKN7i1CENVZwhE
WSEwcGBOTn4CH1DGBv9prtzh2riSylPDK83DK9FNbbE9nALJ8wz8ZF7Cxf1pWnzQlqL2X0DuEqPC
U7OFCrG/cxji1Cca+vIqfIkv6jO5wC2B0abKtFlIMsgYAmB0VCs83gt0d/m8ug4D+vKjmUIKZh9a
By4LZjxiC7ge1QtAIG1m/dEuw42zv7s4Vb91UULkkFZJ9zYMW5YT4P2q8g1MNCrC92u+XbOkry1a
1YaCsn1Vyt5yHwvHi4O0f5ZBbu9VTY4P9+1LhLAdRFX2GAkGsx3qXDm8a6oSs8PA4+T931JRwgav
KCwCfv+rwr75hYfmoCXGCIiEC4I0qExaEGvTlCSxUElAenOfBmf6W5WYkMmGumkO0xxxAWpuDpml
cTSKLzJ6vyAYofXX1RzVnMKnDeJZH3jNyWRAv1RJiq0BTn7jM2UMWBQYAqX4yNzvRVRb92SUNsSO
605Vrgp559YGkZLNbM8oMno9aC4HQ06VnFOpjFUldseKYl13Orv/Vv2A/dctCS75LwgGawre64mT
eG8UuY267/RkYkLr/fz3dp1NlGGsRYB/kSw1UgnkakFeMsAlQ4YkgDFltFqW+gAhkqIfKxzYwBGd
7kBCXwG7RiaVrwpovgJtLfmJ+7daecJbaT26VfEOqD8Rkst7csRjbI5OjuWjCeztEErFjWOfdaWx
Y8wKQCz5Gm74vDvrozFTOX78shfXhznBR3yTBqBS/Sg/1aDXIVVfS6V8HFa906KBRYWhkavwBq3a
VpbIxGCZBwOZH3e2pQ7WwaHudFRt3pDB/SzrdUaLAVc+kCjI6GBJrlem680SKnQ2aQTMHhKCbGnQ
XAP1o7hvf2Y9LFV72SXwuPj/xwWrjOLJLKN6x5MAAJxgP2VXJlFK6eM7PRfFgp2u56OlUBNHuPld
hKQDwhCAHKbBLMFB6pNzqgq34KZje58CzgUA9yGHwcO5S8bQQbJK9jSBYVngoDQeRAMUID7CGEnt
KpXIn/Eg7zTcreXMDqUQu16RzgJx7vbTKWuuN/1ZBe2I+9d78/xrDDsRH/XDVBFjCQmiS3m68VGk
Zavy6Ds2R1blxbmo+1peCdUH8RobnPYSdYiaKfi5zHkBT3lS6NIcM42X6HamCgtCkM21IxkjxQRx
wfl7MdMiIp0I2cnkz96c1UMoeUnMynHaAL4mdhpGfAhrfYnQj3ci2vHM1yHK1tNxYTZGzTRT6tPF
yw4XbgyBtMZ40vWrOceN7wRLJIeq4nmcj0aWXfrsZ2BQ3IsSOpLiz6hQ+bjgd8YMvbNw9WT0y/uJ
l+uJ+wP1QNZNkQvhkdtfyZh9BxWlV/8Uj5EuzAhkl3balW6EhgMedydFano9E8Sy+aRq3Sus5C0s
F3LWdjNpVEJ63md5hkOxC/WUjD5SB6LNyfi8SqTljKmr9HJ/AqHJgBl5bJczvzPMxQvA2/SrROs+
ONQ/YwV8oI6xcnujAwY4AkNcwtJWV3CutwpR84DGG3KOgBU8BSX2zjsFB1Bh5zsMnX6NdLUPEmhw
1Xc81h0/+/5pZsVzDfwsU47KyDOFAhkIzo4sT/YrEI8R3tqMQwMWN6LHTLUMqIMu4C9xb1++QiI5
NsZnifVwkjNlQpMgSCpLqdjYmXaWGjjo/ZTHtsjrLEKb+GW4m4shopBmcows77I8rU1tnh8QIDG1
I+rj7bCMRyfLEusFyEcC4YGhwdpBpKShTb/KYQWFtBcesYhvkmPPNap7s5A9f8DV+UaN5KwtmZ+U
3aah2zfEpj0/pksBjJS4bUAwSgynSNaedQbqD9qUi5tmfTrGaCUvXYk3Ozt5Dz3WVCMrpe+vhl3J
CTP8OVrtAJZkM3YcmEDulKiN7Atp12fIyO3LWX7GmmLP9/FLxwNBBUhHdMoeKrCIasZEVq2s5x2+
SVmrMu0Q9eyG4hatpD0mArTxEwyGVKGulZn1QzP9MDG0a5Xv7yCWvXB0fMw/H3vsXfLDpiS47qd4
lqA4WaItW1tC8iPKrMdWVIY4oewEbE/WikxkaPVuUOEB8pDAPb/bmHPqIx/xLK5wJOWeyXYTWKSw
SeVu1I0ZaD6QOueH24V29HizUf2FXIzqtebQZZULb1imL/eJUdKQdSq8o+Oypfb4xNxjgi46IQ6o
J2JWLfpDxZJ444B4EZaRXRPMR0eNDwn125O5Q4e+B4Rt1NhBhH7xf4zUeMV88OiNKWgTpU7IEQMW
89bulLw//IC8wD2atUjfuokYx187Y/I+AJk8FHnsZah2VajAPx0Y+cbnxkoOJ474JmJt52LyjoOt
o5VzdoPB7HAOijcjcD8hNxsmKR1nKvswkFg9whQvvyBQ1NtPvbNCa8qFij/8+nwkQ4InuIKsjmh3
TJRNpobLCBTI6mOFVhB1bFPw5OICCNvu9/50wbdLu1QGEepe6MYggCWUdMr9SBvvRsXk1Kr57sq2
zNTosYlTUCl7qHGjirFnCjQYkCRADS2deTAheFdL9K62QrSMbF5JynSEmlT9z/kDbTnjA85o72Mh
KDVkZ6F0VGzlclNcj1J00U0kj7kvtgnYXcwgZy7SvIv4G6KlPEeHMJ1aS3PlkjIyeQkQvuVVJCj/
HPXl8kaOaXNtkzt/Sjpkuh80LMrKdYIUcPNCbM1LP52Q8EuWXv6K1HhOEHF7WvcqV13pR+cufr1C
LqYsZrL7mcz6TtVEelydEBXyOkK9qx+DkhP9fx2gEhYOgKfm1FHlu1sfZyZbY120Ncg8fijbTRxT
1AtrJKVoaacdH1mpCyaLK2DmkSM2rRHA3GNWDK1bPwef+PrAm4E80hHdZScBHy+aQH3ljDzJ1z3h
tGaAreHdWRkhGx2Vf4PfFtYqRVpeEEOsgR4GojoxtNZ9zCbg2sMsPlWFLdCLgIEpKL7DvzGVMRT1
PnBl6bnD7OwmT7sjcE61gjI2O/4zx9O7Tiy/ZBwOcufY2OtW5QW/Obv7My6stXWXVeHmAfzofYpl
iNwUd5g4jSx01Iavd7pB6QKsu3x9TRZXTmou7TyODAm1RUgDs3ykT8RPaRy1Hcp7tyEA8Gr5vfzH
xeeQCZ+rQQZrVZlIf9W5WyMJKV890lz6mTOJJZ1oehYJNBMZqvILBvtdnrQnYPoMqPFbDLBPSAAy
SeM9kPoXfdu4XVZAY9IQIz2LMy1GK5FmYjiqtB4UWZ+F8j/mcRM393uNird3thIlP/6Ufv49faK0
qij+UL2YqP8a5f8fG4u+WhrScAlWAMCsbtLAqnOWg1r2uhadfa0anFsRXUr6nKxswGZAv0URhmPG
G33lxB0H/PJmc7Ri4/wdn6jI969+0rk9NtOlBC2vjHUtfuLbpMyv5moau78pNmHRiJAf2E3jVfnc
RRzeWGHWbovUvPbZYK867e3MRZGoMjTqWWEYLLHVwJEm1sExwsVmGNBjYyhpzDIMOhg4FzADfCdh
HxUDPN8cCiEjLWNe5zwNh209GLVLGjMRpFsoLW+qpXEwQz7ouuoEXTdSxqkJ8iZAWdOBlkMKy9GN
m9OBSTvUl+epGGTsWDdNCJbqAKtCHh9Pzp/os/y441X61QyiTmjrF0n2s1cIX071yg5LCU7RZxDs
QujjbuiTNIindW58afX8n6jutyZ53P95uOGZf/fuEjK0Ox/j8t6eWv8s1UtQC/GMxyVgh3qsHDPR
TWV1n2CKEoGGAtO4b0XnRf7DsjI6DahdVJ10L3wRGdEBxNkGKlfl3iGeoNUbPDIaX9v3Ej7fVcMb
EE9wbhdJRxFqdSwpJmp29ElVwWn/3NtrTpAX3n+WY02NkV5Jw1Nf9m/llXcTKYm/E13mag3XgoiY
2QmQVs4kh5HnDErnwsuddBerNqnlyGRbA4fU2oP+mxsY8RYv7gx/ysUe+svEPFCOzy0sa5UZse4i
KXnOOiWpiuy+yzBMMwwmfrx5is0wOcfpxfatMe29Ldkxm5pSfDV0pOsddQ1DXqSSVyUKGDhlnYBn
JExEt04VVZRtKOzyCy1gtSws/zpFquzFw+t5MjnfsgGdVY160m1WMAiYBjAz9x9meRFmqzAyy4QL
nZoex5bdH4G4GPsjwBTV+UVqVi127eQMK0E2+zz+EMmfzDTFzIypzT3WWP8qqLhgmfSy/1dJAXSV
9hxsyg57Jffv/hQ67YBYlxusOJ9P808LGBWGZLCWCs9IQPK/V8JHjsF6O+HrDo0RuPuo4JDZryrE
n4bs0Y8FP2ZRtMrf0E8dWO5R6TSNLlKRMV4Y8/faOG5p93lSEoAJlFwu1VZ8Dbg91NgnVBjZWA/x
o2WqlNVRsMFMq5eTN+HykHphD+3yMZYCS3F6d3Phmj0aCkKZ9+60vjtLLZfDiJVEBi70BEMkqeZS
zGhoUxs1fAWdTj/sNQdI8ZF3F0i4wbNwlEVJUXHCsDvMziWO0/QRXRlboYIM7AyCRFZdv6SZKGjS
NwEiIRkla+m/XCLTGiKtTkIxaRSDWUAYQBRXoh4b1a5DNfxaAqNmsZxRS+YUlfwQ+VEPMD/jmatI
ckNaMMAdNVJiP9+uyNGHg6wFZABRUw6v4kJSRwrg88fB3xYbQEuw1K9Z/Y2uVn+4qD6PtTlQYnJi
qTtsnIWtF9oMeN+B11RdlyKQPSlKOZYqCni2FqpYmUXVytLvK3fxOGEjudYYw4mG8Ic2n+tHLSOa
DciCeWvv4/wVU16/JOhcEQSv3VbH4bVqnq75tHoLU93VF6Il3gO3V7OolwCs64JXcxfbY4PLw5ho
zvGVxl7rAhMjjhWeLaC4uQKtrvXGfpVV9uP2cv7JDtiYtBY3AS76015wm8CvbFV5oXdKKWlVMvfV
dlMx1u/6G4Prxz+CmW1TPkkgNl8C5azadFpTjViYVcHXfGBOVLzBq7gLthXxTfj1yyJrvHpVkj8t
YBlddnSRHcJLk3YaR6dfZmuuSbxbx/77U80kTCIr3WKBBcqK3UsSn9sSRMuJR5B0LedFOe+cSQrg
dZRAPbrOzecipfXPzonRNDNBZs/Dw7wyIJE/MSM56CxMot/7n58GdY9GvCxR7e7nXFqcCm6CJV3K
uYWpvEHwDP3w7m2t6gWXGO1bAbQ2PE9ft7DAXCztMNb/him8pHB1luQvNEvMtGF8Pk2iJmRQkaFP
fIzBcyqRThUITRKMibnZqDiscfyinAU7uEACMXVSbbT3x5bUUo3LyDfbYq4Pk/BmuDyNBT+7JkSt
ZySnaHTIiL4gw4zgMTTvtonT3ZSJrK+T1XspQp57F4/umsjP8/+HMGSN+oICtl6srAjHYoOmLLG7
/9QszYhMnHXt1HjEgBd3xXXvKgDbXk6BUbyvcVbFxFhKvrYv0BrvWGrEPYeK67FmPxNNNf0ZpvaG
T3jg7hHFkV85isAV8MnWpHZ6Ao5DalH3/ZBdUZsYKJVP0XEefqYtRREy2wEfaEnXgVj6g3py1Ri7
7yuNQ+xyzOkOfD0pQLG0ccItGJtOIFtEscaxCR7iY8T8Bbj7Ubk74J7e9dYjAA/vlRuX3Qe84wP/
V1xCRaTHU8XqkmOxDw5b3kMaIvnqfWoRP9CZaSGI6SrsZd6ssDd7xFIdtPJahJehFIwgDHLpWE5x
F0OqP1fJYYa7ivY6llEh7XeMcLSdgjDxohZ3WHEJc5mPpx9kFHITfwFlKjozWGvXpcfjy4sgxlRj
G10UqcipWQT6TUmWzzOCBnb/wQSbNtllW2livuJsCp4LM1x3vij85Dce6g03mLLgidIp6jvvIn4F
pRv7VZ57Vi2LnW0fou0/o/HXK9hVWH0O501tj3K2SQNHAx6h6pudEmHHBr8X7wHhd9WNZjnkS5Ym
lGFnBezT5T2NFCRoOBIZSHkEBo2Z6/X0ZBQrJPEy8QXjKb0EnNWUqE7Yg4g19f6xZaCq9b6pW2/2
+IKt3g/46efvvlbGS6MCl3UV3YjEcVMvXD5TnK4bTLLdlzzhH8EG5jIlRUmrXqq1U03h5q+ll8Up
XZQnuBSAuaWagwRu4orp11JTTH3qKa2LTEipZu8+nTP9jFdjN/TqonGDAqFl9nHQB79sFrIpue+i
dzwvX1OZbH/V0c9YnPkCO/OokKDDh31KbHVypGCQAptlYzPLjQ8T4vLeOvNO+SjQF6WYcNK6kIx9
ei5O7780CCtsrTK/3tNpdfedV2dqMWAw/3LAMP0Ljd40KjXJquOIElDNXA6f8i8MVaOQQvj3hTnf
Fg8gZysaMi60ibIpOThi0oSYEiPWaa1zGPiFJ91M/pjii0RAyXyQHyDJRq1i6ooY+NMw5LBUZ7cY
eI4J+3elweZhlAsUY2+5Qee9Au0k1B7VbHRcD3heEOnjVBu+Fn8AJuU2zHGgTL/GPshtbHlBsGPE
2d4OqS0jsxI5IdSbBPhKTKdZiwwflIVG8C6jlqheJbBhcVGF+DwCQLU4DUt0DJMbFj6xueYka59q
cnrpYOMaUgGj/DCMN7uMLySc2BrQK6Aai2ehaktF2kgivicLQRYlEBdko//Q2AsvNRw8K2EF8v51
j8D9oTbXMb6h5sObn0zdD2A3+uD8ZJ4fHW1qkN9T6cviY6yeF0Gqv8wWbJYhYasqmdL3POF8qFil
Wk0eJszs8joOMjdrMXU8ovzHtr9iQRpA3S1DU7j7FE7p5vrR6uoVtyHIzzrtYxYEpXtdUjDgkinr
xnTp0MaM7M3I2f5iN6GJGsjIZnX1evK7CT2BrlGQLcyoFooHNTAWTQfoXjRySrYxInUO/53Pwm8n
i6pNI0/CxL4idrF79GfOyZmSKNTpUMxCewzP2cRTLT7eKxuzVUZly9P3uiq50TdcUOa8npuotnIZ
GjnN34Eva4gRJMvNt11T9UzbL1OqcOVGuNdHcQgpXwkIea6GSFdYMleYrO77LOPETShAw1PmXNvU
W7PrTV8+v0HyiM+0SSB4VpKixbI3DbY9SCsJ1sWCiV3HUwAR2hTz7WWlFF6nEY3LPbtwXUzxaQh0
9vHW5H+N/oGYLTrbEpttU3l+XdJyBgbXLl9YNmpI9TttNjwbdBfKk7h38WOlGZNG08LUwKkfv/dG
b9ySHHpsoJgLcothfyZTCRPDQDCd2+VMnPgxcoagvqI3IMS5j7vQttjpZ3OWWtQZJv+n+bHiLT52
xr9v3InS5fJmDhTppftik2wQ7cm3/g5WbbnBrVyrZFxtffpwbl3GN44Dm4mdDK+7zX9JoNFzbhWk
UFb43oaiwJ2UWgZ/A6PYyNA1sWMTgl7ZVDI8XNSsK3mLwEofPTCIEfcHCUIveaqjW6oYZIcWUmR3
YHeBGVRrULk1peKn6yHoi2jevj/Hj+zZ4OVLg+GrlX0S+Q2QVxIAGZ8Bz3TZrCwjfkr/ksYecKyx
AEqO1xonTzh83kc15RWzOWJtkM+N95c1cwGmKzT0KEbZQNGTLodUSu7JOJTPzWiIPEasbm0Zdvbw
g0sfJLB+aO0g0URLltULPpkB5jT6jFz5MCtbGkSFiBJ4wG8lW5A869JO8n4bBziNnoJV4I2pLEFt
V9AeEa75a+cMYQX2hNmsXENkVeMZIwtwmpoG7PFgEhKtVS09ucgMOfn176hB7jZ8n0KX2SYac9bs
ny+Y+EOeqQsvLx/cfOq7pFXtCU8VXThbe7OiaAuGdWOAXzEsv4bKh9JdF+5BXlN01kxvvrQNpmXS
lkWDCTrFMfA/tOMHnnPzDUX5Y284sJPMJP+GdKOpi+T9J7wXzZazCLE/fIO7/RzaJPhzzSf/VCoi
pdwc0ZgkO4J7MxLrwoeXNCIJiD8OfqQc7V6Vb1xfUSFTz1g0AlwO75ZZsncGj9CsHi6VUE/UVQ/g
Xp8fMQLdH7Zkz9Ta0bBMvmkeNYmGwj0n91AtQ4pXRXCC7T9zqsXDhvQI+0x87XRsDOQ5+C14YnVq
JvnTnJeq+xNDe6yMCfulNmgEZZN2amGSN/aIAKMSqezSuk7B7iYvJeGsIXwlPPwvcLqK8rcYnuca
XABR4uMD3grNs7UO1UzHvxacycZi18G4hhvE/wsfiOAwRPW4a/wUdFfYtU+H0zq75L3IRqdD8KOG
SSSZe6DmNUufxh/hQly32UAf53kjXL/RTQrgKGUXHJSIUrnQOmiqRvZaERWLx2RqzgJGUgDllPOW
0Hp+/ywofGncAfEjyA0JaYfhHs+kHzIdENR/sJQZMsiChphODXuEmmL2RAswau4B/JCqeAa7KbOD
XVp7MG5itsnJfH90ZeULpBVRBNvbe5AiDCYhcv4HSL++6VA5YFr9BCndlq98Y9JMxMe6Kdu4J0Dr
7LEhn2n31n8f+wX8BVqAj27gqCTbpOJjbx7bMehPUYLpi6GPbVkIn69ZSoDUHtudw3UVmgUTao//
+4DeJmyxaisv/6j02LLyTQqY+7RKEgvHgLPBmHnAVgfzZT8hixPGhQFTvJE8UlIHkGSzJLOeMyqC
lon9tR6ApksonrB8p2+63R8K+MG6mF5dleF6Hv40Bqh+pCFJ4Nwt+6y3YUjnJ/7TcIvzwDCDuAPm
IFZR2NokH4TQOnsu4S70dSI1N+Tr0qNOJZM2tQELXnKjAXw0zo77HSGOgoaMljZnLlA0SMsVr4UU
MZEOXuLILbNDapfuXhJs+4Lc7Ux/gPwPjt+iJWR15JxCANXa7geIlrBa6M8X8G7uU2wodXbT+Z3J
PHZY8T0DCX7W1cGVa90wxPeF/C/s6lUSwbjvUMI4Hy2Itsi+GLjU5xjCHBVChFdvDrE2lEqLaJmK
4Hn7NjrTBPIZguvaUeAVToCfHG7Wf8lSmOU2kc9PCFlLRWYnzQHUo4enTcTYF9jrdwi6YZE/RLJB
JYXuxHzJvxGMx6G9tU4mMThbFPRy1ncKxNYpiJ9pau9LoAix+b8+rG4KpwgHeSQbnmzwgoPPsnXi
C/qjp9ZW/FLwYbjXerJrLAL+CYzte+OhLlYDUJOxikU+K5GCpR+gQHLvlt/h3TFgdKDwytAbgVwr
6d2SuFLCxf4pl5QXrNTwVGS1UZwIBYHDBaa8YMWe1wUqoVe4L7aIhnA9BCxVYJAPv8XakmYta/Sb
vtuHqLbWGO5ZkRGh36DwLpnrQigYgBG6jluuNuWZ9noh/uj1hIjv2dp4d+YQePdKlSnVLIpWF1OF
gqwL4FUIYOvSRp2IGQRWXznMyC9L1XzwS3hUNL+B2dw8Y7dWB37AJxX9AtWk8eqrnHoj9rlzUb79
z9kiOnFwvJX3cCLdy2cIDyTjC4GHo5yP09M9DepHkj2EjGjODgRI1L6xNAaEXsgMkVcdJQk7plGQ
7XUKgzMMPr7Dk9HUm5x3SXUPo2b2BCna5cSO/HLWkb8m1Q9goeUPCuwpdgWxJVzuHj6333VZznat
Uzs98N9idV8PD956pBlxTPp4rExqUufwKCLE9I59QLqchnuWASNU1tXbhMmsvhvQGc60MZPP4Pxf
evFoHCGogpbkhk8ceRM/Z/BQLJF+A9cTWJKQsPdptwtQrp6zeyc5f28s60uAdXIcTCoCc3JRcJOQ
C3usaPv2OSkCVlN8Rn0w4CamhinVrXEtvWbrL45zB6GLLPyEgguYnVrrvDNg0gON96EHfvVF2OyL
gHaL5qy97OA3NgddCjsnUiFLZT9kPJSSNmnp8mI3qpZ79huOxGjlabCtJNCcd048dbAnM9TV6Kt0
q7HpqRgSaDkco8svC5mOkSuBYfa3ocepNwas8rOt5avgN6740jmG5p/FrrHw0tuTJFoIJm75uSOk
RUPWV8M3QCskpt6U7/aujbWwzKHWGIRFvCwLvn3Jm8pub96VuzrAlKN7dBa5ZsdPfwPGYKpp5LmP
DvR1gtY+tvncc5MuPeT8FLnaPZfmBbuIeUgMBGv0YJOVf/Qdv4Qh/HjhX7g8LZMm65llBjRTLfYd
U+Pz0BkNhg5E+EwqSFDWT0OO1F7RHrcK3m+q6/ZHp5lUr/YqD1TGv00URhDrLtuB8kAvh3FoJHP6
dNACCN3v0HD5kGXsO961JW1K65Ny9i2DHMjYSkf9H59yRy6O8dpRVq1ggT+ptDbwZm7zQR1j1wy2
gEd4U6q9/7E/0LeHFyyf0Q0RCIXwn2rZWUMUrsxoVga4vM3MWItEczKbf1oPShOjgfRplStiipn6
L80YqXF4PwVU11JOJ5ahUM8VgpqEi0fqHmaM2upCWfeYlz2nM9MrioubFizS9477cS1iDwMccSAk
KQMPMHZHQlEgIEaj3cjntchIWjr/n/6IOFpAYdKiYU9EVtiBWjoNYvEvrg4KXeFm9oSJ1s9UHop0
iZcHaRVUc/LB6WeYfV1GBF3D49DIRAfnR1dCnyXL9L4/YBZM3N52kl8OvxkphVwZ8L/r4WKm1MMj
mXZ4JZkIdxukWf0fGV1dtFWpFdYNGnsb8bKW8Q3usQwNFCyPnW497NRo/t5FVvyVUM3949xOmSy4
vTYT7T+sfcOzBTh6cnu7278uEEqqQbxRturZnJEA4xJpDrUHSdxof99aFi+foUTVsHVHl86IWtBb
LbAsuFkml/ulCFN1+0TtnajcsX2i0hT56K/La3RSoJQUdv9ZpH1gentBMbN1NdPBZdInRhxMOf3n
65hc+EoQioqR5ML31eJV31BpN99T6QQpR9wK6yzwLAbvj4pvk5MQJSgqv3FpgpWsozRIcBFD4Sfc
liH+81LPB+DyQTtM9Jg/Xg3gaWScvtpnnIfj6heu7Q87qhx2mmY1zlwzI9/hdWbvWsheU7pwEqWP
xDriUR/hjAhx1a+0XjJK473sxbAkz+c76e7Zg9mJY7LIu6O4Dy/ufqjm8UGr91dEyZJxnAFH1hK6
x5NtsyLtw33sTfInlXdxBVTBxtJwWJzyEynFeEk2qJIs/eQrw9+u3p5Fial23u6vYuA3GD5Wcfjz
DLlKwnEAyTFMYyosTo4RvWifE0tQCfdrgurKVmJoPM3E1bT6jxAYBZGtUmrdaG0eIvEPAwGL0wCQ
7QRQnWSuncxa0BTjGo5ii/zOEtmI3O9+vmkjY8cc7AhPrhfJcnHofjy1VZdo8L1pxJVv8eoII9Nr
wtoLS70Ncg2fCZQx8kk7hAxcU6p2zIB5RWlS9bF38nGKBu6bU4JqTZbhaB2gNYj7jCKLg/tSURNE
pl3vM/FjeZR7Kq5XOR3GORcqlWra9l7C8ahX5OCaJ94f/sJeW/jB8i/tj6GVAbx1/2YfclYvvQkX
togT5NCNI/gNMSp9i5j7aQkQXwHEwL7A/lQUi3RUpOMqgHpYfZvoiuPbC3PPIXe3H1jK8PKQAVMK
JKURaw8JJZ0CbapastEwlFG4uRCoarOuCUXrvc9NgNhgR7CZcchjHYzuFPHIcLT/mQT62KqpkKyg
NWQOcI2U2FlOCszgr4vKxpFO56sUyo/pcf8DNloEgN0Sl8vsCOfmqYg8rceeo3xxUlDwe9kBxsW0
t+UxWUapvLZBC3RT8muieucXMXqVCFdmFedC4cluzjoAa19jInR6JypvjhHakBp4Yces8vw6peor
xqolpy2ZwoXpGlurcnXRparLSXR4Cu4JXDHCPxoV1tT6VSJE3/+l7KqpTXwkSp7lT0bCiqI5pEUM
hciGnVC6S4biaFW35SVFgFZcmSd3BfhIn0XIdQeGM71V7wuVatd4+qH6DH6ZxGj+xGGFF237AeV+
bZoSAHWVZk1riYydgtjSy2UjStTkM6ZG9Cw+toOIa43MNn1bvVkleQ+58AzX15wSU5eAl3oXZswg
HW9p6h0x6/mkV/kkq/0VCvGdErEDMlpDwqkedimaO0edg6UGCPFyI4Mgqgxe8ADFOul0HIVua5CL
auilzhv2S2AgAyS/1PL4rey0ankLltsqdO335HKIuwjYFwCoLcwkE7+ogG2+Ns7+AZ3AxXBG6LAZ
ftLTZP7NlxG1Q3V5eb/o/Hzk2e6Vrm0Lxv4dmDd4V7zc7Q2jjBU5uwcdGy7b3t2AblXQt90EcpAv
BsTxioJsGa75dAQKWwP0p3nkz8UazNsBFQOG+y5bCRgzAWbWAhL2Xybp59utXJB9ZRJhqKO0tRtu
HfwPNzb80+knC5Je8h1LRwatrn/26ZnABggS5E3HvofzdjTqCicSK1EwVmQP90o10KHfsxG7HrqV
ccdG0MLEWtoWctSTZdACVqLiSIvmxQBR/MKcZ5x+6CZLlFve9+MXp7A+WrNxqYLFRhZ7Z3qiBdu/
NeIKBNTyi/V6JbMDseGF8pXLuatchuIYaJsD8Th4x5Po8NvFSQ4vSWcbBheXbhHaHkfl0Lggdkgz
T/lCEeBP1K8790pPeRh9kH/S6gzt7SXk1eB2BmNcqVDfBg6+uNgWVADRW3lOXLYplSeiRte21dyL
OI8dEjF0ebZ2+QjAoEd1/eT2f1npN9xCzPA5k6eeIfbP9zBxWN/na6i96jT9fQOgvicyAjSwQjdx
DBJZZ2FEuJ6BlU8VwgQltdrXfLdKhix25UL85E9yG7kGKTH8dqiUD9aR40baGCGwz6X7zDxOHept
xINf5bEiREqm+lPz/JtGiJRoFQsHuMmU1B6+PbKtX9s9iOf9jNL/cDg8niSVM9mxvtB/bqBdV79F
63XwglOX4qcx2lnyd9l2oN27igL7NzPZ8h6jP1dYgS11qUqVVLuDafOXqdWTikX7sK8jwgMnLQ5u
b7U2+GSZqweOr8Duo+E4nJoCi3S9sgV4Rfr5/ZUHayXwaXR+NAAol6DmZxRaR+sWUKnxJuHE/hxp
afjTucZ6SIX2N1yt1hkdEnBNZI/y3cq76PbTmONIV5I1H1mIc4RKyBLN9fH9FSuEnZqjMAegWDRN
2wERTdoYNxd/0u7NDo8eMOAberVK5MX6Yz/zp4/ONkF5vKUe2hzK4h4bkhkRkbla+3QxcZXdYgnx
0mqKfI0L+uy08FJNLGOjaD9kp80WnCJU8yssZcvtiEtDAcqVokGsEGVKOY+AxT36WsLw+tBhMiGV
RmVX7Bj+MPbjE0e9beySYGHb96NqFO0pMb0lVudtJzTCIqFO0tAd1tF7niBoWVNoxUU98Zr0P0//
QceiaagadqtEaIO0L8UEixE36Vi5KV/xEk81h9CS5pSrTN1qN/sJ2ifBgmOyZ7oPBmpYxRV0MetO
OhxYg1u40gYOvlYNUdF9t7p0jx50TFbKHAkGGTDP6OqABT2wZi0lfGQvlBT7TAaXOjAUhtMOZiKJ
9ptFm0fqH4vg7/tIq+GLZ+YmAXGeRUhq/YDuU/BlnCXAOWcZ0BY990wcW6xQ58NhsTrOhG19v92z
jng41Kbsd6DbYWPUfck/h1VkrPyXMeso7SH/51GZXrpHTaVMTQT4TJ3DtdIEXoYy6AzI2F6uEGkw
5MC5oNlEwtG2LGXKlAmrF+nt7etbVswMhPwsCtJuqoqwJdaSHm8sNwwfIv5cAlm7JYwjINjlF/SO
TKrmwMwhQXiv/crQ9RvQl76uRzX1PVvxdX6VcfygfA+WYRcgerRigBbnOPdBDQGDfVoQgVrtp3Et
N3ItfHQuhS+W02m4bmPSlxKksgf8K31KkVL0aWzpmi0jYcgeKI6FWUrFjJg+bbikZ6O5gTBrfNrE
xdsNaOGx4PjKlvu6wZYCvrtZvT+QXSOzRTddSx3JagDq7YkhkGs3Fc6FIjRQCiz7pj2S68DnBn6J
nJt4WuM1N+QHiU1csnyPVg5HdpmXftASlL+a/sUZzZai6aNwQ1hsfTYVbnl0FClP1Vn4jY5RBUoa
i0VwRdWvTUhzqI+uK4aFB9oe6N7ttIzLOTFMAS5UJPFp4X11E06z9grEoYaw7YGdFiGguLLmGwqN
Yk13yNq9k+LO2Fm+kHXOFPg6JIxEVdiqRD3MpGhNGCt+NynK5vGrFzUFrE6WL6ciiTWvbJpLc2v5
xTflKu0UhSA9cxKdS42VuzKuBFQFiIE4BDONGb3Kf8uxEGAP9n0S/L1z4x8RSspz+W3aHUY3mHC4
7oMbGpRfZJVzUSJIqxolQUuDrZs3Z69gblXutfst5FFZsF94lrhjGZRz5du5pvG+XrCh/4yMg7aS
Le72Ovy7tmzI/d48gVcIn/QEfFdhVZo9F8LAAP/IulhvCvlaBO0Tsbqq7+HIqjuNzSiiJv4wQxuW
5oeNKKI32GrYwyQdOIHtWEaatuHEiF2BcY8AOREunsklOaoXGXCw7FtdATtEr2Kc6NViyFSLHJM4
aflqgrC0zgt4t5mN33RCjimSJZfHIfQ3JOqOr+s0dr8eY399EsabDyh0GKhos3F7aBr2nH4Hhtar
rVgW0bnBPZlqybPXHJfSJwShImrQTOalLBhbM3Y56STgfx96lclt/k7zSwGm0L692uAZqnsy2LLd
yzW9stpa9YcDSLiS6Yjh4xQI2nEnBNLYhRh5O1VY66hpIHK4P8ujRLis8Djvgqj2yQF/iMkIsqT4
8H641ae6FMLES8Ib8g9zHReyK6e/C+Ze+ktp+0uY2jSb4EWA9RYv3dPeq+g4ZjJUqsnVJxt8Poud
dQjSt0bsNhyo3OOWY+XSrzge1bDLnfylv1BYb9NzT4ecyyjLq/gpK5yfEPsrH3GpwX8g4DzTudp2
4CXK72YMF3y0B1+euochVi7qwH819wn8UIA5MtxNR4WQZLyBb0neb6UHIE32bP36US1jbV9PDAtH
N2p1qpvmmfDlfPyEdFSbuOn77A1Kr0pu9z2ipBLapJPtTqSWegbpXFTNMa78S29M/Fkw/Tskj+FV
d8NNguPB1ZlXLmJEL62tWRheEVIGle6BQqUirSoYfL7lxtLswTfFdG5c8G8Y6UkZPFQIuMr3xa61
SewSRX/GcSmMxpTvwP1OwAFJXGrWPBbfXahFn6+DPieZhtftdtvpWMjRh7P9h18e/4DOvF30thlh
6j/qGf9eGHFUzyWNY9IE3KWlyDZG3F4PtvvOEsOM80bDNVpFV4JSS8XwRWd+qLEOz7ySBVLPA1Y6
UBwvnLARrFIZr6fwPdR2qs9kUfmv63fk8CIH1bbSOZs1snPo3xHhDbKa4zInzusbx7A1SirkZpRD
jxDy3wEdDtRSmICWmXktCVAVyTXYr5a/0I4E4nwX4rVdpAY1tJVmOp8fpkDSZIooVUvCZIUK0OpL
OzoCuhgb/K7NSyKWz387i8RPBDKrtRH0cXpAECB4gDI/ZqLGh+7tqnNKl0AreanPS/g0Q+b1zw7U
Rhi/X1Mi2g7zsYOQkxl5yZZX2TlyK/IWe1jQOor1U7afNAo0MJEU9JXJHYGy9EgMaHCuvmNiFkwR
SQzR+rHIwrV7uB/wzltqPo5XIlU7WzWbQZ4odFDxBGFrmkoXYoSNMVM8r76SWsI9I/AZdTk+vywL
Vf1WJDhAoclqhe9Z0wv3pbe+5W9jxd5ITpDM7wIZbdGdiNKwtb9A5ugd98Z2jbX4laklnY7vr7sy
BZXODsbHHxae91S9Hn7hsHt8gMwVkFtSTWG5qLl0cfGD2hbfTTuze/d0OG7bKxQIF5xVPlq1BPQp
2qELxebct/fC19W6E+EjGJuBga5XWlnmRYT3Ya2p+eAiDbPEKUqoLiechw0c4C9r/DbVvnF6Syob
01l05F05WFnXO4nRx4TDSPdxjSItsOyniMUpMoCKjpDRKdnTSyaZFpXigYDIj8YZMkybAjvG1V+3
Tv00miPagfMZZsCqdlIV5PhVfsSETT1Q6aefaSDXMFX1C0UyTbeKMDOtEF3LowU09Scy0zs5ztiU
l5ETHHW38PrM/fxEiOeUEkrtHIIf2IZcxaybX1ZszcrXneyZ24eCmudiTOmd40re0Li8ag5a2zx3
ujJSoRFrGliabNBgu7Eo/F8UlIn9CBcf6w00y+b7+GuN6qK4tRvY8JoxmiYtT9FglJZQ0A3oXGbM
vQxtMly1hEvNsUxUfWFVKDd7Z3YwkSaFuQ7jr2HDqIDKGUNBx7zYJ7gjwwWgW2L1d4UTNM2WMtYr
o5k1nzbp56qiVFH57xgxYkpKIuWIym3XpKd7cZjM8Qgzqzw8MPVA9s0EIRq+u8vf37w44+KkPCMz
Z9jsVlQ/Yi7GmsWaUpsU2jvtdRVhOyZQz1lxDNR/pC6JRuYufHo8iXLCIeEhzR/7X2GHf17d82w7
Czn4QwB80lM6E7gyldv/Q4YEmNVkHbzrfKc/Qa3vpkZwhCm0xGrjjt/r4Y+S+8UiJaeP87pMFpcx
rUogHqxv2lMXmgY8Y/7F4/MwEFoPxjqG2V+SCxGL5QFxyfrDl6ZFtj/VXldJVnN6l/zmzHM7poSu
S78yNNs8FwrC/d8EaYbsnzzONYwO+qV69M8FuzOvEmyUMdzw1dmmKtFuBLEfmXzlwSlYQ/TZdnMP
6ljhrgID2RoRD2KivBOL5hyC4QVu+V5Zs+zMFYL3hSp17EgjmsZpsOYfV2Sqea3eTRfQRMQj2pb3
Qv/PAKdtu5oxO9DWu6fzUduu+P5xxsD06zMk0MJyVhGRimhzTRdMy7lJC4mrrA5kdUPKS1t3YCG9
HMRfaj+6khsv6oDWJ5ACPYgpud6UEoXXYGeaJ5npKdcndE83AZO7r+Rd2nqCxbir3NEC3QRH5k5I
NbAxe6KeubmiUvoimVTF3RWCS9P2CjQqMd6CnYEfJmbm+r6LM6ShBg/dMvs3OnBsOCM+GasAa4co
lD0cwVBo+LXT4qKmXo4O/KwiTZEmD8Cf8ROrhRSrmLnGcLG7P20YPlvxAcKV7kBux01uc51nLPub
D9oJJXKmeo45F5F6W9xV5OPwhijRyhQhEIGSQNkXNWNdJ/SI148RF43SOE64Dnm65o4QxShBYGgQ
xT8xKvhmn1//fDvbrRQkA/LuGB5HSaOlJ5D2u2AZ8nEajFEIQQjHDjte4BO+sEXefXxjB+EAwSOQ
e1JZYo1h5+YrIFUacLDB/+lUH3oXZhKMqfeVQg/SrqgBZW/fSoChuI/W18wHo4fclcBN9DxIlVVG
bdLcypiGyqGOBGImNdSgikStAdJg2y3PbdmX38dPkWtybyNZezwTGMqGy7WSzorZs7xwd8U3Rj1u
oWGM768AFT59FN+z8Xxf1rUVizfreH0KyNkafbZGfXTr9alzBIUDlaKkKaHVG9w//TdFMfobJBZf
yyImp7Ubp9pQHSjohneTg5CDjxMrXz+wSgwucN4/uK+aF6RgFw+PMn2xH3IVW8Pd8C8rJ9skphg6
D7Q3AsYkXPZD98cqwfL10Cd1h+EMr+t0qCTLrU+giKi+4Z1Hio6ikwry5G6vJvC6aSRLfECTgUBS
qmotgun6sX/etgp3IEIED3GnLXen44B8IdE28rtdlAheEdqIreRkv438r0Q2iXxMp7MHeDlkjk4/
uk0UaKc/0k7X6C1Ic+cNBZyjloMzdj94yDqoR2z+Ofb+nFNKVdjbJABZE/wWR+J//+MHKUiLeYaT
N/jBI4OMkuLaMcV0GEBk8L4gkltqltvaIjRfoAIefTa+Abyu1pRFH2L312986rhiV7xKL6SeG4b9
m2kdm6+WrhDrKrVF0snsZK8nFf+eKYVOMQaKwo5bJonMux1E8JK21wrPCxAuA+tlV35Wzn3Xkk2w
TnDG8XuseGRSH3Xf7vLhRgm/BnCx0iOyMHxBWBom3Z38XbRalSzwiSmv7Va3jMmbtFVnt4aIk16t
LWbJO7iq19qSC2Dd3ibyEliTgR7GPXjc0dev5pdoChnrvC+6CNVVinHpUQegj4OvBPTq2AizO+pc
ZdMEZ6CaVr1rMw+Nm9wQ2x5Wc/zQVWFKhhqGszVOCQu9yzo+H1da6RVirs17y8YRw6qg3xBBo4bg
HD6z38VfyKOtv0nXJ5rv4xj8sdOJetv9NJOLKxDMpWi6wG3F2NsbSLl6CfqteVmuW+7EJrxNWaO7
JvtKNZQlwD7q63+bSO5QD5VnRYd/vFvk1j96WAKkhwvUVQHhRxd/c64Mgmnj/pa4lE0RGxWuX2NN
bEWOta1bD5fxPbd1y/Z3v3c8nfSYFlv8GUzoRrjsQclGiJukQO+XsZ7MJTvwcvFVITmnw3QH+qeh
UT9YLPixlD/bU/jnHuPxhUOnuEEmjknNw3/y3NbT2hwF/XV6pCZ0ZyQFNeTHP3HHcFcBneSIThjz
JVsKNPwSVwmnzIHCialDoaGSTod02eUa/E7UVLVekiCZvfk+iIWIEqFwG/9vnnVLnSdtC6MehDzn
3k3CMf1YztktI3So3JfKeJjJnZe/cLxumGMZD70YcQZJA6Wjbj4eddV0P3AIxH5qFAdEgSXbcKM2
x25orRbau6nnppYk7x7t1hPz8jZhzIcezCjVfZcaUJEsvSuWr64nl1vVAXV2fzx94fbhtyr7LQlL
bqfJ1nnYYZKiXH85qaIS4EonlnWPh9qFuERWCJ8QjKNkR6K4AoPxOGdoBe+tFO3DC+aBTaqGBhJe
mQMYXuinJQbzFnn1NL7zM6H+OBATlwOHAGxqmaygWVKR8+Zn/ExYL/nC17+kNYwVy/099diz1DVM
nQohmGIktd+fhTkh7p1umODVQqk47HhF2BEseOlcFnFeUXeoDTwHrDRSeRdPRIffh+kxx50MySMa
Y+2o0m78kIyPFYLn+ZNrt7VuV8cwT2pvED9qgp30uElOzfHwb3OSQGZ3Dic7CI033BituHDI1oVa
6F8l49nSEQ1ioSSaNR5Dq26n5Yk0t10IdZgmhUp0GZzwS/iurxCpKQfhU33XHHZk+Kl4v/DNXH9l
DV7P0I7C8SydHBcoX+EQjeFaXm6sc3LmQs8/DGv00CfgwX/K6GZ9weuf3mKQD0snW3MiaCZMKfGV
DV+2nsiN+EEeAvkUhoDDGFRdTrILWSPA1l1Q994xydOPHViaQ1Edezm09qTjr6RBFW8+xrQ3/RVr
xsULIQtyV6lIhGV1o7NBiLEJQHKgphdzB47DwHSAD4pwNkqjIb9F55oj023AF4TYnAYzUwmeLkK2
Mi1rZvMjh/UgPG1ywbRM6iyogNQg0sUhl6zD5jdTIEs2t/UFj+wGQvn2MHx3FtATzDi72cYP24Wd
7xWlmZH9xTvDIprc4cs0Kcw33CITKr46zdB5yTQBZ0ewlnNvszZtv3l/k/rqsV9pMB1AAD9MjoHi
NEgdnoDtFktzDWwwFi6K6oFWccGmgLlVwGn6XNwGZKNi5NytmgrAPZcMEjrQnb7PO9EYwsGHFq1m
KNN+W7DQQUD2AOyMbw/x8zgmcj1FCpUqakR9QY42Og4vNrN1GPqLvTzd55eaE358GoPqRdte0wDM
Fctx0uYKY7/jXQPkqFNQNxpFY7N/URl4h+R4Fw3ZD1sfvenB/XHTn805DrIX7aa4tA8E4ybKvz8c
5fayN1CGBd7Yxw9qvE1LQ1UMqnH47KsPrwmmfc3tYO2QU6ZymriMByWr/newB5Tzy88nKr/f7266
6Ausy9ZhDhbq7ShyWBw178XvDeE//7lL7laseAv0ri+4v/y3nwFyQOgwxEJxrez6r8oVuDMd3MeA
auxl14JncgpINevZiyjGWE2xczkrXU0ccaIjLy8V2BNA983/Yiks5Dn7tj41mEEKUS7iuvZeQPiL
+hzzQ1sdgf07Y4SSe/AAZs0+pbJs7vnNHyxMpms1uwDOwKRqkz6m8RMtngBmuorhQZJupMuVPjv7
qXAbDi8azT2j0enRqhvQRaTA/bC2inuuafJRhmTRHfhaF51MRjjheSwye5QKTtWkvFsKmk8aR90p
v3ubqgH90oceqnvYiM0WZPlczmNwR4uuBtI2rzVP+3A3Vfop5o/MPLhN814IY5jegudX/tQrvrKd
Cj2vhQicSK5t1Mx3kJRr4Qz7ey5X3Rdt+HOEPNt/uZnVRx7NXGNYY9f2jt1i4+pEFAXr55h2pkGf
bmQyhnYX5XpPUh9YyNSjuVkoonI6XWpxLlQXdk4K2PAiJtpX9x9IczKZ3YPRIp7UaMgrTzsC4sD6
zsC5r/hF+F5HOiya9H+F1A182enDxli/axzZ3re+SWgf9MrzAmgtMd3cAnodIcPSm0+2o2ToDO7q
wtjJcPTjeCjfp+DaOF7FKLd1OyKu9BqqWroL/IAGjzmrrb5BAXzwVbc+658ceWBrsy0XmOANkh6r
lrRCquCyW9yGUdD9eV7iNtRbPThUtHZzc2VyZfqzIOibGFVeKnDL/2kxAh+ZGz7EAckP2ECVBsaY
KBizsviutl2sSJsZFgW3TEjiJ6g8zRN0sh92PjlBOUGhiwLZhDI2dJmysbkXgr9iOZdMR1QHphjV
AOwk4Ls3R750ibUHgRiJ2XAZLusbxAkPR6WqbAW3YU6e9Yuo/SFw7kmfAZ+lA66XFtP2Uu/+fHOT
ES/elfVH+o7HlNZbw2npjqKP4J735eHubW+6oCKOxWaP/vr0aO6Vd1R6Gp+WY2oucUNx7K/CJLzu
8Qzw0GMaZ/iib55eNrBQo7kLCWcmykrM8LAFjiu7B7qLYclyjJf8oR+pJUKQas/jalF56GxpAR1q
gP/Y4cwmT9ntR5O9b02Fy+Jfn7uwqZRGr9zRLnQfob7HwFwb5le2i7p4W9+zcCNqGlURnrDBV4m6
icHqqYouOBLH1RzR9XaJubXDPlZCbk60ofy6PFcyg3bYmyUHjsweuq2bF3GTk7GEiQXfBxS59iEK
n71jFTSuU0O3SeOHfT59RSOnDQU2AWw5ThLBpaVNCvGdBxt8E1OeZxGWrZzKZuH2lDIM0mPhYJlv
HD4all+Vvq0Ed2HiON5Q0hc36QgaYhQlC6GtbmMYzl+x/DD+saA6l4SpmN1PorEUhy+rh672t1Md
se6YFd5fS6lmZfyUcyIxfPzJHSdiwKL97g65HPr43ViOAiw8gNCsAWfJNOyuNDKnTxfUoIdI/73c
E76lLu0crQCmnBZQPXjbK8Z0ycbUtpc6877mTOSTfnx1n38o4imUgPgbrwJoWBkTiRsi70N70bsY
+HXir7uTFNSROKDsOHElcSvmhI6dj23fUzUC05v8ttDt0RXxp51/eei6MpL9L16GjMyYh1vOg9Is
8rGD497L8KmPB8gtT9E4H52WU9JiKZRI5VAdwEVjpmPOIB+Ymhuie00znge/7Qm5Wdp8EyKg6DQ4
D1aoPpLNlQwRJPToomwCUlovFpQWEpEhPNZTYXiyxzftmCB0atUwkHzeViW1/iH7PV+qGtVE1Bvf
iq8SDyozOEweTNJvjhRotbltNIigO37zG+NaG1rgdMwuSQQCXidqRnVZPCEinSOo8WQaSiPGU5EL
j99QWZ0i5zWOQgIlvH4I62FpfIz3iSoxg/0mhXvqvWGAVrYcZQn4UzGouIY86REFzjWNC5FpDPNS
FbySMbir3anm1cqHJTXL2Dx2N2OwtUfaq8UOzOqZFX7Q4cp+EK75txrRrj2IkksR2rCDVHqXUPq+
WycC1cAL7fJEpEmiU4zIjLOEUHshapcAE0kggn+nAQbTTl4V+eB26rKyqYSLy6rKtx681sq/mM1k
GAcTMwlXDigTDTylSK1NiLTOT/JlEma27XUYQY9JrVhzhg7ohiSyBVCpJHFX+lG7rD69Y6560ZmV
clZ8oH3CIWIAidPoTLxwBAOA+LPMOYcB1BIc2rUorqLUWv8tRNP21sYMvgdXX4PmqOlcBPhXb2JA
xmyHgspdqj/hT+6vKmRACfkU3JBMJIM2v5+2Cfx1ZNkX4es3TIKM/w+h+EHWENKakPXW6yRa/UqS
krQMX/buzCIkknJxAB5fMrpPvoYaIKvcsnUEu+tLCIcJgqzqVT3Aq/SejO1I615zSCNYRfCQVWoA
uoMpGckLUbKKKVZQU6PxvPWFw/BU/haw5KyUSS83QG1Rf4B8EdlCq8YNBbEbNKLUg9Hz5+QhMcye
8OOWAduJS1MKjRAeAvrqcQO7DsP41hhTtQyjfeOYxMxsrtBY65GnDo7I3cfI0bRMCskFq3dcxtmN
fDm8RXnDwJCv5ZiwNEoIjs9Wlx1ppF9utjBZQCSatMkZtqc6+H88BxrD3Y3ONMr4jd3IKqPgNF+B
PRW6LPQzeWK+EDdtM1GG9J+CsqiZQbVuXatSAZibPnZmf8fRMSFLKdvlqxj31x8V44qNk9X0Chqf
Mhh/XUwu8171GSzLI5ozyLr0yY7ysPJdEYR1NGc90AXfJHt8gPbJCiaD1/5+CvAZLie6upoDz6KE
HgYEpRqDeeN1BPPjYypgId4Yv6lhhH/3Kzrkelpue+dPFgBcrzUtLqWSI1QTuxPGgBaK/OCBZDAT
48Q6gwYhjRJBn/H886nd0QYEL9vHuevKQoJiMdpWOjBDjSO3Ku9yl3gwm5pjhKCqgrSgQMmnucsl
K62x1NRvaWKf3pq2HYLkO1sFTUuBeviRisM4l5eOVLFJjqteGM4akGqqP7Z7JAlY0PE7ON3gNoQs
gwxOX5BLEGARIRIBRq88V2Q9mlRglvWifAVmCM2qP9dEjQaBJRmhlTG1SaKBhOtE5cT+kR0Rl0gZ
iotz9VE0+tqhnVlfjwDXprEHkP9xPITA1jGowKATmWs9rlzOfE5RDbyy9tDdm/Sx4mwKy2GYYA70
LH7gLo04tCGTkgeFAlw/7mWcRywYz0SkgAtGuszlemoJlAhwmD5acABMekYx+HCrWBl/O5fdxZqp
g3JX9g7dcBl/bST5j9/3DxEmAK1Wq4C2QeRziVRZFxTqrTE6foTjS9DLnK9McPsZHxuTNd/XA79v
E6Gi20WqibaDgOvvtTb/Ek5hxSiz1ibhxU3BppY8aRkjbJx7VvHMXfcXwWaTt+ouUUzaq7NPCZtU
HmFQprbRgtSX4tPoLot0gv86oBUnbXPD3/W4Q4W/I6F5tecdCEdD8cHrJkxL2mHuo0nZLHLt2LwZ
3VWtwWbdRj3WN/3nCh+ADIwJrqsml/JH6tMxUJv13PNQuyIYdGSJEQzOLtzv/FD2W/TifRxmFWnk
XewUwiZqCvyWJUU5KNjBIk1qgdfbpK5pM2mBdDqqosdNlSyOqZEDF0Farq0LJigX9x9EEivLz8b4
ycDLtNFCHl93BiCF2PjPEuXlYF4SjXUg/OAf3mtKjjwfmAy8YSKbTnWN/fjKLSKIIFf1FdPoElK5
jWgmC502jAOmfTxzUP2I8J4ebxVOY7m6XiKt5rOslGUAEisn2ExTKbyARHhoima6aIkuiILj93QO
UCQVtmGoH04Dqc7h4peP6oJ+qWvRVsyhANjlqDqksBINX3EbwjSk5dv94tcgc8/557ybh+OneBU1
UAmFyoHhMtcvYZqDEPfQr2ehl2dACAqDAJKe2xAHYgGY9dtPxjOmIn0bsj3Ur47rfllVUaIZWGX6
P6za519vG2f5xvlOfeawDthPtI0yjt+XiVvWOnpFf48e8wzhX5agCrLxZQoh0G0w/GjxktecLWsa
eFbYwuOw6JbYH4W+L00I8ac3EWpaun/7BQNrv65OoeWCuCColgIN9zXub8pwzYD14bsrr03BIUtV
/JrUrB7ckGZkNWLNAJF4VR/165jQ7iW01NQ2hiiVA54mDrhIK4Kj1T5e6pk0dc/O9aBmWZXxLkvk
IO2x7wk+nlf9EXWd4/f34Wa23EucCVEfxngVsnkTGFSKYBJi62AEHSYZ4gY9ZEN0qH9muQxwJ2DB
HYB++9xrjCMm0dUlArJZjA/Hu7t8cBNbXinLeq9YSZzAgAp87RqzmY0vxuN38PIa7B4g1/CN+ww2
ZKOKEF3YfP5a3gHaFDcfjU6iTPfXn5904M0bwHBZIhGS+sMHg3I4taJotsjC4dxQkzxu9ApFq3Gt
2TpIzJw3i7gxJWQLMPf46A/JunO5FjjOFBLfeHdylY2fLeqRlBhblW3ZySSvuRWG/yjkKMyAsWC9
WUR7DJEeyPMtA/KXc3Ww9rkcXXHhT0yEmsMIletygTTnLx28T/LMiJYlJC32hW4wASZ1OhkDt1M5
dpb90E7DVzxZ6rGbFHVm7OT0SNZ2fxHgRIg1KpOvsyVhqLBKuJbj4ZN5h3pDwtjFoLCrdxaxJrfQ
3do1iuAJewhXaOyDSIWoUxNSv1B+YdGxVODtEPOItIVo/KBOPsW57k7SCj5rynI8UWCsw+NjE9ow
NeIwCJT2VI9gLYBegOTrlv4F5DO4rtuk8uEZIj4YGwVaAdjGkqneoqJ/+0xknpEKfeDyv5f1jtUx
4sDkUet1Wtkiph8QuiDIRDRvKNsZO0oGCSg87DLHSVNs/rvsUznOakYomh7qv5OrM0x3YAJ8YN20
IONLoU++45FyX+6Zd9p+BDcRBWG88ksFY/MRcbP4j7fU04Hcfo9LobxK08jpKTbNyTo8KGyE/OhC
D9h4AA9o/hdErA+XotJiArfHC+dQeR++VOudc3/we0s5gZtz6GrSIDA8JGziISpOyY/Gmx+KBHBg
thDSifY/+XvGWuGukm4WVyTNQMqScfyH8/YPTdUx1ypFHMjDz9nBjSo6VQCSIm0pTT64/Nht6V6B
flrkCuDjvGDwdKBiDMClKzpJxjEgmy0IPk2gzdizXIjiPRJQ02FmyWSJV3e+WUMlwOwl4lof7peh
IQoky+EeizXud6UPVXrIRDQlRZRP8szuvLKQCyI1/JXDTLRdIH1G25cIyXJIqL5CamlWe3GjapHE
5pKJ210eEQ/AIR2F6yvhkZx1HwYLMjj9Qz/uqJh2h9Rbv+oS+ftX9xTnkH8ccFbKnGHYQh3VhhgC
l/mLdDwlEQrDNqSpZtCv/GNCU0XpnAZoWrUV8UiQjCjGBQV3BrS9MENnWiQOOCHe0pYEWM7xf1I6
+xVpI942mWHh2OuUGqPxcXhrBBKkYPlxREopFzUMHFihswG/+6eLj8xycIC1zuZtk0BeHcI0dYzl
eJrWh6cYuCcgwjkDaXlGvgcGSVIY71gZJhmiSy1D82fnEfhlz7G0I+sKvmGr1O9MM9EZRc801Ffo
OtZLhH4/YUXQ3v/BWUQde3Vz2mxJAgkqBQbEDzGB3qV8XgoFzI7V7kfArGmnTJ1xgbbxxM2DAgzB
Lf2mEWqe9PSN2Q5Jzm6pagdPlMXkivPy+1jqs9ooBjUMTa+OuUJx/jc4tP5ahmCbSMi+u1xkcQFr
watkwJc7H12G/FU3PCsOuvtqKhEvSmc3nE8evDzYkua2iLFeueUCwFKHs49pSAJjzwxokRrRplzy
axQkouwM9ZBEFsapez7F8CdNYT7+YqlMJnV4bH0zWQfFsv6gL1kEyeATJ9O5ywlJswJPmop6lP1A
r0iseqqHm2lu0oUWELQ2DbcnMh24TBKp/RFyrpTglWpNhzSK4Ok4F9GhhvRl8ttb579vnhivNfxz
w2+irYnXhSwsIx1+dnfrnKQspdAg6ah8a3Ffjo0/qq5Adf5i2RTIVOo24vazvBn8MvdkiHgEH4Ar
uICdLCWdiOGExeh6OcuMin46unwdMVjv9XJnSn96fikDz6lc2xJCFOUhCP0zmIyJSFH6JQCmnj9A
RjZxG4H9415W8MBJbjGwQrLi6SDtbfNDkNrTkvTWDU4aG2aMoVd5vybL+OahMjMo26s5ulUnUsOI
zAQXziwyUQ+5nPDBxvFcvehRbUTHNRoZ46qdhD0apHK2OCVpLboelScSZQ65OVZARqSAS9I1Bh/B
U3kc99X9otyL0D8ihLRepSyS9b1ZfJCzhpBT572dvrTHsFwKySXQYXhm4jbsMCe2pR6DR97jVklD
e6LCUS0RvSDyz2fdO1sW1hyBZksl+RIKhiuHjLJyMwH/nWoWlob5IpDYE7F0fkYBNnBJCXjMH3h6
m6yF5vhxkpickOtzxG/198bu70PTQIe8wpI7zrORgUG90cM85hYWPC32nghGmYVUntAftldN37Xk
Chr2bzzY9Y1vJw1kgwCEW5KM57MBTr9O16lnDbb+KZNZkPyBsbhbphOXnF0jbB49gmmS29ipaWRV
uhxiqy3l5opyBLgateMlZQ1NetvA9Z+cOlpVHDuro9LJQ5aYoE37JXln7eeJ2RVLJX/MrHml+CGH
pfngOQUQvTRQtLXjJOCZXYZNZV0pPqTQ00TGAWz6gJnXp121Z7pSaUxEOCj6IGsMHfvGFD2fHwLh
2XvbPhkE/unXi4OJkIJ9KX6xbokBNax9P4BZdJokv1jApA5dNPJOYtycaP9JGs921fo17iKd6DNb
oBI6qU8QlRk+/mlR4c18mDrSPB73Gha9TdlmuH5v1V6gvctG2SZwegIz/O7hitJ/8ozXhu7Rghti
lTZGa48uEL9k9pLvF0GNkZCAJGUML/RfI3YxYmxHUjBRNa15uy8ejLz7fRajXH4xilOkpuU3Vvnd
EM7J28daMAGHa57MyfN8EpIo2R8QYQXyEJcJ7XJDDRK3d93aFbeQTWhbnNVTAmWeAfbkxw9mNXCh
TbAaZXpJ9Aw+vxxpsq0DHheJszqXOeZcZUZLrsY1vjiLV/7oKjWbYsPj1zmCbWhuytIPx0deZMb9
ZoZRclse1VDCiIVD66WciNa835tRKdvRbiI2Pu/HbRrf4KpgJVS8H96T1lbZmho/1+cJXX+X/NO5
yu8e9+urJV2FOV4nYQSqAalR2n48lbFMrgli2jJCjGFRd7medUhqLZsxN/zdgPo4G4J5tuVHs/Vv
YDfI+wdt5KSk+p3GBPIV2Xml+H0TGL4B3GbQ+5d8Yqeb2m3L7MzB8GpyZ8FhtGkxxXskoE57Sdif
tCeNv9dGIXo7YxO5ak/q/uV/9a1srlGHCVMlo1JfH8j7qCSOpWj/FihQQiittYkPs2sEyWMtfbE0
m1Z1EG06UfhhGJ+4cirJc3bNoNd9lk18TiJHJiNM1Cw3p+kH9NqEiZum8uPFzPA//BsTh5EZd/8D
hho7OMD7H45PuX51+Zz6SrZR4mwMgB+S7RuL7t1z6AcmRhQ9vfR959cm4cej3gENmTiJfV9FcTh2
OsKb/Cqqy2DTew95OmLFW7O4/tSnYtE8WxwMp+eFhV4CTmt/Sw9/CyUaZ2PszuEybwLVjmHjvYf6
LnDAmBcyqJvWDJ6dSHRuKxWvp66OpV+8qiAtXXyzWcK3losf2bvToWzLyk2xxJQdZojSt5DK5JxJ
DGHGFgTUHtbN4pl7wcZ4g88/AcwCJnbvjDmEKyXa56OKxWfEKmpvnyYjXevFx6JeCdlF/KC+2D3s
RYAxg4TnJq8M78h3wPcqalbnE3rN/LwVbWub4bnNOWpHXsvKEH2XhXOvaV3fAqoomYQL/bIY5keq
T7ydFmELXXdAfWlmfdWBx/bDnOYllW07ZzO1T5zV+JxqOWcb13+eY44xI6T1L9wjUD0v+oxRtf4d
q3Z4A0ygDgSEeg97APIGf5nvXgz7ekeq6FzNmXOa8iW+nPAhZqrizczBC4I550CxgQ3tW+mhN3kL
+/QgDpJnYswCd9MJjSrO86v7C+kPqNgJwl1yCaGy5pvLJfR42hPhELg4DukZ0F91JIpPTwJgcR7q
KXAwKY8MFR+/NEDV9tpGe8t1RWmZ6fUIVWhvApCLgZCvyg+e1RKRQrAhr6z+2SSgHsgvl7M3Pk5O
kEVl5/+1FlqhUd6qybxQGzUhiNiiXI3tdURWF7WZB1WADg/ag0t1AdTAsOYFGww/lIJ1bKkBIW8k
dw4AEAxXM4bypiwHLonT7CvptsBLUmU80jDLOpfd7qKgaKhJZUDHCUtU4z2NRk48mLG9F5rM2eFv
o5ozYkxNKenJTtBEGZgHDWqp2YUFQ1qrAQ0mPmpMmfDY7yAQUyLkwHe1q2VvDDpCd00eODB+oBag
weMvoOXAmFsc3dry+WE6+xiLxkNl9MUBy+DNZ3RNoKHemCec4pEOVYPWIUhObzgWYsolp0rV6flG
wolYDrdA8JcnkgAJiVU2I8IBBSfi+FXkSs86eAT1cDgla1IydHkU6LiYtpeoHQ6cLc0gVwGFfWmN
FXFUqzFiCW0IQqv37lDBa/mcaD+e+E4qfgausIJCzgYSP++3LDj22XKCCv5pC97+rlBT9l2CXdWc
hu+fhAYARe37H7BzyovYQFNG8T94fpTsrhS2YZ4L0z8lSyCP/nWj6ZVYzOdVy4oZ5Sx/s2W00XDr
nimU8iNz9ltZSAJ/1E6Wb89jCG2B6QutYdVWXVNEKb6UJX56BZoGrugiDYDxT1/1+oqu5toSYN9s
5JFv48ucsVj6UgfVu9dzfV93npZz+pe43urmr8qwG4NeOo8ggm9KZVh1+4L6wKuTxXHBAsOp9uvR
sL5g50PL790oPiksyLe4qooSu8hnJRp8FMN42x1X268bWzkl3KnM+XfiZQ+LFklDgKB/YtLkVE6u
FKXGKDUBVC9TyDZ25nP0Tvm/XuENIRAdYEQ7x80QJXMiFsJXtmOO6NyUV0gWAkJETRBcxVNLr8ui
RmCkql0c+c+WFkIMJm6QkdPdq1NsIVYLlKwKUdHdGOoh3nh/VSrFkzQKFqGflcy/Pun0iSomUDwT
0xzNk2ueICIriLc2SGFU4Zab+h0Ld6s3Y0rDWJ/xBq/XU9IDI0vF/sS2d5jWMY92lDST+8mDopS2
rXERq2iD3dBK+6Kn9DBbsEc/+iBJAnvMMFiToAwlZFm4wmWGp3CekDmKc6g0Jde6xw2KjLkOtsJD
uUpSsVm1oWt9J68ek44VmO3SVU7zdd8yCajp0h+jvIiVs08j209HI7TmKysZe4/goLhm9DfNFJI+
7Yt5L5nFjteBuDe4A6eqJppev9UB4xhBHw2LjdSQJG1WsqCDuqn4KF2FM59DTegGDJb+I7BdpUBr
YyqNWCeeeR8vJi2SYLvZGx3gQcyMttKpC2ty2YN35pb4iDWFggsOKOmOg4AJdngaHlOxB8OaDgv4
+Kfvd9wMS8P3dyRM8ahSO5Qk+TFJsDNsjJKI9Qk9VsgWWkTyxNQ6+H3Vr5ADOqSz0oU8YqxGRhc1
TvGWZXsEeIoTFzOJRU4dwxJA1yPSUfz0AcIdBaQyXl1UIj9cVRCPki7ufr+oo2tNZ/oEcbblu7E3
hoIXvCL50YCxFl3F5wqlzPnOWqMUJE0KBZS0btGVuk+Zg8JaTdrPuymmv7yZ0WAiqyupTBPMveKA
eaYAyoOyI9lG0RGQRA/knxTMwN22g1CtgNzhWJsRmjpTqMyckpT8KUsZxWMDh3VkZG9hUne4j+ex
kKrmaWAFdNuulTb3+UYY5QSU5ZCijhIi7AY+YaEnO2eX++fAXWnWARVl9z4PtlmacGPaAUkiywPO
iNYCKR0G2pB2EdLXSV2CCeRyVCl3n/8cfj/zTmOTka0NI8ybbwDZB2ZgSXddd3ZtK0LjOpNEFJHI
Sq8D+y/PUg46623kzaadhnLxveZLygSSEu5XCaXU+r9/uPT2q7c9TTN9dUg0GHmVwO+fuEYC8AN7
IU1lwthCpQl9EGOlzgoz2nlzycEetvinxD5nBUKEBExA//9h0dNCxk20gK4BKONZJGjKqOKOj7dE
iC1bM0xMhqmLI1AHUYG7+oAttXMa/L+prj3vGWjujN801EElw3rZrc69bY8mDD5WVf0bZwgAJSxR
pQIkclqBUBEgaRmvMMKNOlwnKsYkKVwF6C/6OQOqKTR2DwSwheJC1yalRt6nILlYgH5Q8JOZkann
WkYjIpkGxC++sczaBkYgCjhmIIA+3kbr6QoEL8/cut42phmS71uOkO7BlxFsFjqOq2An6ROr7Ag2
EOqbVzm8c4ZhtLHxhEnJDf1ququwNrNU2WFOfU4Xx2T66GgE/oFe8zQbTF3I9VfWbWNBIxYpvuOs
Xld9aNfai/znPCKJJG4hn2WKLCKD61u3KlX6/nVyuX91gr6weFa6UBQl4EMUm7m5uLVlJxdzLWc1
1MkEZvOFUt8TPqc1CCq6zBZimLhvjxV5xh15UrLHcYO7COg3FXXgOoqkhXREYzDHe3RI7Tn8D5xS
/2eozzXRhGEa/Nlunogi65dskoJN4xws6uj9wZZhqDnXz3kv3foMU9jrOOJ/B1/H2p3Qzg8UmgA/
bDXPs3PgVunEpMZ/bbS2kDzcqwGuXjCZR6Tyena/Faq9WSHHQEeF9cN4vSMh1wQLidpl9qlaSWQZ
+InSPHNibinJZ4Er7STIBexb6t+MqGOkoQDcj95DxdNdtfYnyXIIxZdXfqcrxx1v8LlmFKw4q/O8
ZcEj2QyAqw0jDcfmtLdzmRLnlJzbpw4vL5rLsQCDNW7bfGxVHjDwQqSTjTmz9cX8F3gJ3vpR3Ura
DgvLG5erGjos4eZ2OUQUTu6D6NDICPYGyDASOuyLY2IGTlW4Z/E4X2xD4IKoSqvWZkDh6ADZqyR1
/DsrTjoCCfGcz3dO+f0WrzVQ8CfPzbb9x40o9tkDwpBPbe2ZH69Nhbh+LsI8/HQ3gWnAIfaC6qfj
AnFny4Qzgzp+bDmB4+zRx0Vuwreu7Rqird3af24XbbjfnR9D83AQN8qeCptiZKFEdY0C2VCmbASq
cnyXK5/3VS2/y2qhz8i8eziIHfECetWY3Ur3PSGqDkOy5HRQ2wSnx/NFtCFvLXtUBhBGdyojk2DS
OpgSyCXTjeKhkoleMhRct4Y35TBz2gU5SbMsd1eRKw8HUmkFw8M8YuP3/nqvp2cxoMaVoOkdtuI8
FY/xNeRwUvP0rGO3Bgz9BzX4qAQc7f0mXsyR8iJpjyG3dAsyeuGTLdjRkDQ/bhlxKdnqht1LYDxp
lbyxyATH9Ww4X6Tk1yAS3Dgkjlscom7gBHkDBeRP/KOrJK87nVBexAmtwV3SkB5UvtVOP8MGaqzg
2MwoygC3aTwZMCzrcgVg2gDa3OC5jsLn48d+jbq9hB/8hG6EpCRdh1xRz+blymfIw3kciXA0JbNo
dUHxN6Lxe/PigFG0YstTxtWpJfZl6gp2Y5KzKOhbwmn+xEi/BwcxgP07TZcqfn2llRWSRaU2bpAm
GWji6xTJIj8Y0otg3lNpelwLYX2Ar97m1jk1jA3VAp+j4pkQu8sV2KscmTtbtiEOB7UEAEWQcKYM
OqoDahybr6L59g1ZRnUYV9VILntQdNQfV9xjXv/RqoVPu3l17AcDEColaJglfhXrTbD6/KnKHzIF
Qy7kRbPWllkqv1+/CEqGAp+vw6yPnQgdfRk2XespeswGj0KIDBQP4Qb92+NUTrYO/9lhGpY5h/og
uqjpMlVfpdHU32yAPivy4z5mKGMUA6bUIRmu4w5XhZeKSJ7nzmNAA/T20qTpKHKXLU4R2NfX30ej
IA4GXwqx1n1Syj/Fa+tVA5ITy6hcVM9qX/w279DhyCxR8DP7kuHwREXFj6gGQULB1Nu1wvAa2ZNg
4dIew49hcPall/9TK287pgIZs+hp0aEi0USLbMWGdNY2l3uKlyx+eg/mv32WmImBg24GR6szHKVM
5fkh5JCp8bG8pcVlU7Mdc/nC64hnAABmoUH28BaSm6NGJGMNFUI9nr89yiWSZGwnn73RAcEDXpUa
PFb0VXI46kE1Jr/X/2fTkz2DaSQRKkktRacMAuPfAJN847+tpVBpx5dBNcECFI7WSnOyD4g6TPQ2
Nh6zzJelJZjbAWrHFEqof4kQzK6M8erRztkMIwEigC4NSf/S1HXCBJ6Kwoos0zRI2uQNr/836Zfj
faIj5kG3GWrhWk3y6XLM3Lkbu77XlsrxVKHyyVAmsMfMgdr6FG66ZggujGu0qWS9QT+atagr76/K
M4X8Sw06cPYKv5OVP2vAz3sOaqweI94cRcDBRsPcR+F4TolYAnHHW/zdI23oDZdW5nwMRJ7KmR8S
3qWn7a3yV6PDdYVyF5sC0O0UYGP7ERuS8+PqylBV4P+nEEpNYV6VhGeK8qmXwxZoAvewzvZUbaac
ayj+wrTNBAwgghvRK1evRAew3a+9sa6atIKZa/5QID5M+zDlsPYr273N4PYBOft9m60X7C2iBrrT
g8pG2xq4fbjILh44Oa3rbB+DICKMjwQ8sgtJQNJyvA7J8Enh7CdDlSNzCh+D/aoCXSiNrpgg2J24
oYO0N/tbxexhaTtX13g8It/ZihguLNCSTS3xWwmg0bFhQ8W207lHCUwBXIo22VFAxEi2zJwS+kHd
ihIOwJibYm4R0C6iw3jOkj5VFBX74Z3XuhMuadIgPAkU8HAjmJWYA9vbYQZzedOc5MuEhE3aw/wq
gVqUEiRn4ec1LaEw7bYNb5Wr3uAvOdzHK7mh5NTNAY5KfWn5ze/E433sWEVPBqIJqaOb6o4F3EEI
c6iT5heamtPU/PF4j52w86S4XvtodAdvTKq6IAlRk3P1BSm31UyignH/8mwFhGT3y5fRQ9TrmOBe
Vb+tUb1nckenhwekRxy2/hHHl22WD0cRHZUNrwj0Vj9St5VjcLjph5SMxTm/Ui+NLPyKUip86flC
rvY0DYuxtIgxPhTWzs1Pkabp98g+DeyNIVnVDjfdB+rXNJT7XpKJDw5hNjtXkM5WvpTQ3etTLGka
tQqQGYaA/ced9GcjlLPU3GZgMdgtoEy+riIZIu3nD4K8hASXcdwo2NDKLF/CccR347uOG56IQIW9
FIQyLVrewZnzwnU7uMAGy4ldsYD4cPWxzTZ5xDmiiFm3j8JVLEG8EUx5XDDZzmYsA4qFhg4fbFZp
RNHPwaeuEEznhzDqv7fufbTqyU6r1VQ2xaIuCZxeUdJjRWgA0JjgzGPSLL56AfSv5jvEtq+spul+
iKorm5nJVllPmRFdfKrs6sphmZhnuDyEICAYaaeS/fMG709hXXG4WpMd/GnC3bRMFF4nen0ZlQig
dprFZkwmslDFeZLvYMK9USOH6S1yRAT+xMr/WhGxwr+INytnb1a0XKvFEhbjtyV5drNvi7px2K1r
R3xwXnXBd8BcKIBDda+IjyyMjT/SyTqjREo8R9ThiKTCzOXfsnAQLjij6mpsaGOF0/Z7AJArP1si
GCNB6XaGOF43BMwepS9PiqQnPgspnQ/+74VYyup6k2UP+PZz7+bXhVMrm5AXAKAe9hA3+whd8/AF
377sAT1gOPWBNPby+x63JuL3PDWHRwyOhIAUxdBKuQXA8gCRjnsux8XpumWMEPyKB3jAZMhsu/aX
6Vx25UE/kOinLNsynqs13WkGyKn0nIa3+h8yPP4aF75HUC1iLrDDdSwRxJ/020U7219rugwhXs/N
1lKH9ZAWKXWVucBAC6S15S0UirzimRPfl15E/99ROSMBkmVhYWapoYgrdOOsM0tOFhiN9APd+DOc
T6o5bEIPnimXXgTgwsDTGSh5tQsoxBwPHS2lJRUUCu+a82WI+Cqdc+eOHvDZ5Aey15+jtGsZ4noA
EanBDf+g8sunzWXakmeO9CJF1Q3xyXYsI6FJyXfyWz1oQ2sBiCOvqVM6hp2p0QixkfQ/EENqHzhI
lzrbPxvrO8YpJGKFuKpURoMx2Dfxsd9V/JfJhsqVMSCoOgfJMaACbCoqRT74oG875ZojuMCAbiZo
ebe6LoP2lb+6W/t7iv9hQFksJpwi+zFgt6LRzBy0+TcGWRed4cNQ7YOxEX9GDDiEWr/zBXLZaCny
MavXTQkNj4/yhbYcqemCq49j1DwM0hCPi8/hd//s9RxwsYShYpXpvZ4mz7t2QR8O+9BAmbqPvgWk
Aobt6MtWsTdbvFLVxMEJzdnFEcMOQdxB167s148JKYVY6dBJqrIHyt/RE5xapU57iVliyY4r6a5o
oW05HndAYM9EFC2jXeHdrixm7KSTPuDqyXFLWnJ6d1GJJ0G+AUoZNIaE7ECUYtf6ONOM9Q+KQNLW
x+Na06/o092AwulBD/Mp9zBREaJpcc/arTfDGZDUr49+TJijfA12AxQSnvPH64QGs5nUAuc3b0nV
O2MXpt0kNjKn2CjnsQ/G6ZfQiQNKj1pIiZKnIagLUwxJxgIgFUYUGPQ0Ozboq+ndOoqhmKm0q8qK
UGAClkBI77wExdn+xmWe4BfYjdhdr6fMDRviBztMqKYhNOA9ePNntSZcs3LWDZT4eSwKnnLGuQ5L
uh81oJUtrSPV1BlhEcttT/jkgHMoxyoBDtUVGlaFxaij/6xqdFE4+bROkaUQyIyW7MMGCIi3hLq5
ejr2oUdamypq2paF8cFPBjrbWoJ6mvVPtvWiMiOQG7lTpApw1fcJqd+q/I6oD1DUhm2Gl9Y2lnyq
pttJb+0vjY3aTfoOK71eT/eDplgVEwSI9X5Exm+8y5TN4OwsDch881jtegHw1e4h4peDcm0vpvFm
ALkZ0KuM70kzkuJd+z9jQ/QGeW/k7aM0uNO/nriaC1dyjO6b/i4Faz2tMAvUT9IHBr5rob7yEAUu
KUUn7Gc+YTI9auufZ//7gjQdZuJOpAXpk22HCfJURMgJ27qJ7r4S4xhjNCbjeU1oIgjNizBpdf+6
cow8kB9iTIYzuraApwun2d/wKLturagCkoVD/XpvSWVVV8hqo0GGopB6iaplMZ8USM4OqGS0DwKU
J6bnpsej2gHCQB0vypH/Y4ZnbbYFdnX1jGTYzWftEQ4N3/o433Zi2xjnjMwO77NB5Uk6S3dyQWR5
oCprBUFW8o6v510EO6Ku9LBE2OAwUzF+8B3xjHz4ubFeUwVudgztRfPlNAmbAtSGrU/SDlbk/BtA
hm+0Q36VMw3g8hCQRRLg7ncH8uDYzHJX2VOrFa1ftTx95Fb/9j6hAJk5Hg9DoiF+6WgJ9wNcGm7C
ktst4E7Xe4+jLk9mJ0wnkB2s3hn6No75ZrWpyL5LDguC1EFx7JH1EgmYYLIu2qqj/UZ3Ob7SHhAf
+OLaM9ipHDuU8BFsC+GdVlRJXvl0UREngRxafaDic7/ShTtFJsbAJhC+T0vYTxfHL4XKZqTI60ZO
hGJhA70hR9q+iofLgVaQPvhMLXchmfgfbljDPGLkzazmXv7QCM1GhagcoHaYOzHTGOnd2JK36YHv
YXbKMQg7WX3NujL7RSXMlhFNAUENuUF/NR8OqvxJ95ua30niNAcMn0xNsOJYBXPvs+NbK2lhXO96
uCngevVNejmIvzGVK1HYJEvGAO6cjPynqzG9cWTLfwii7NjB39WnMllgGwME/71xkPE2hgCkGDN8
00CMY2FklyRl8izL9aKDOoO1zhhEsocnw9Dohse8pjD/sg0qpjK9UQAdjoeckFyTOZaqLQ+4WXFE
l7WYLn6zwSLjwd+D7cDnATGyuU0oLJcMfvtQtqoPWp6SiyQthwXO6qfjH/negHm4NbVAL+xNVz78
HZGrp/QwjRBOoFu1+npLtySoXQgTULfrlRUikJrUFhBER0QdsCK3Qiu7mvROvnLw7BFVRjxQO1aB
l69RnBmST3ean1LGu8BIWqojLz7kiHtmXw9hfI5JWh//ch1PrGU3PzeTyv6eEkgT2RnZZ/9KXoqe
ApWuzJrJVfJhoZJwLuzw78NdAHgPptuSa4mOYSH9BzfFuZvEuZ/u1CUUlZ+ffJr/2HkPr9j6rntI
8apjL6PxENc8hA6k3JmMEOslcL0fvE+HtzOvR4IUpGRBpk4hTw0Sr7rhntIxard8FxVl61nOPgLP
7y0jW+99kvf6Aom3njBGa3bgFWgbSBN0mzXTnNf/4DyLPVuChakU8LZ31DKiOZz5/xxMMiJX2uut
FXSefbhY3VjfFLSzEF2ZiuZWktaVhC25aDrblqBo6NroilY8/UKJPxKHVh7srYAjxwEb+EkSzxpI
oiq2BinzHJKdoeGudIxBNMZ08e8cLad2U9yNKtaB8OEgr5wtkfSKawLviiBEamBYk1dKpn7d4Pmp
aqsrIQUDges/eOTVmEYglbT74mi3RcLrLUDnMM9wgmaCL87mcGJrtrxM3hx/MFc14Tuzr0mNLRS1
m4oY/Id3Va2IfLlj4didjiWEtmZm+QG3QQVWJy0J8byVc4dxRog68kRlCGGmnlIoHD5/fw+p6DkD
vlgSKuBmRYzb7+NCdZnLEYR/Uc7ZgZt/fZ5WnlW80HgdRTT6qSyA7W+e7zqDsFFNKkzlU3C6/8TR
xgE+GeQO+jj2cbxnbj0VOXzyJM3csPeDGB9iYFdbSLCwsNWGezupAR6hRyxuaeZ51mO+Ux/9N6zx
JPRXlgBIvYzsVWs7vGDyC6DkI8zcxVAQCj0AFcwAkV+rZldpV3WmODEZcvr+8zixbdiihNL5zE4W
76RirjRXMaWX7lerNE1FoHxJT2kgPxWR05kcI82fpK4MSjM1sHGiNMGzYRHdvo1/mke32USKYH9I
I2m09Y1Y3ihiCySHZOE+8QzH3OK6lSL05X1RnOdvzT9vKMYxysCUIyro51G2Hf+dZ1xej6mfWoPs
XWhyIgETb2hcQRmvI9ZgoicM+mwEmdHFrzaBS5CLkUNntIBctbGDzZhPpw8nZsEedH6OJDLYPrpu
bBwbZLy881+21ARJjvYn7+2wuAduEpH3L0FVKcvK6bgGmfiwIIHW/Xu+bQS+M7a1mHnwUsv4oLnM
dRYCi9wDuXWO7O/ZVxKWwTffz0DpKfsZo6bNGEpSrPHyO+o0P3SbPbmFaxi+iuVzXrebqXPdcxLX
GcSRH4iZIkcfJ2U3YCnrimIYOtkhJnfLuJ94ClhkkTocywx5YMWC6txP/YlndclpiMl5yZQlFz7K
z4wlu3mzsiRH5psmGfLlLFgADm7gFSoW5IibHXHAcr/lCOe6QzvUaAGYOvOkHI7qRr4IU+avnZSD
2t4dFwZDlS4lwT5rXGdRVJdEL1bKpWe7cCtrSMucJP2LI9XmqP/QVHQTom84fcSaPhpJSKYFBYB2
MOvsW2bYYSmrcEv2U00NCsU+qefRzajbZlEIDl03HpasOUxlvNHQrR3xstxIYUqCdPvAYuQatiXk
zoys1t7G4lXozr44CkGqDct3QmBoIf+2Ac2fZSUOZQ4IXz4oYlZ9zW03YrLiVs469Xsa/jNC1t5v
DHuWutSxX35lwopwz1yS5wsdMecRrLRBvWieyjQd6ISU6QbzB2gj9mcr1ZlLFYx55cZoWsTDYRoh
RFEmW1lB1t6xPcs+UpOXVsbQFvOYnPLp2QKDnF+M5nwy116PRAEzczTV2u5DoOhlQGAGy4/yUQ+j
kg++02S+hRXXJO0mRX8IeFoFBSjGqwXdTLLf5Q6avM7u1m5uZzmvbtKPz/DFdqMXg2is7ANBZ93n
S+DvBUXkfCSwqEe9bgVx8ZOUSum49bI9+eeie0fVj5WrrAt52krJ6cC0J2Vxm3oYW1nMbKhBM9Ra
E2QXrZV1RQTOUVhCjCFHWlD49+6LSR1tYvoG6r8ThTtuanjekqhlL+GbY5WqUQtV5cQdSLMlrlEw
pl9TAMfULnQTTmvgQaFMJZbYn9wrbO3fwatAzEasfGwx7vRaYnc+69HjvQa8bs7gzo+mzhXLgCwA
PRHw/gdmOxkpZLhmD04Fu7KH7HlmDBtKotO6Zns0YiYJAdkpWD5UjIjwJZZhQnpV12kzk7KvjXIV
QCRDoIQCVAjnk6z3OHgNpoPifcHmUNsyVrgG7bdbjF38McH+Ej28Gfs3wL3lPjfwt2dHW5zfyEiR
JDsa6+cZSOVsX2q7/9sGshF2iozWNqRnMykFANAjy8uEvrCvN/5R5G+Tf9V2lrA6i/w6iFu4RyPR
/8SOH6siHqlnC/ZAKawUaXikN6zo565GZMdSmZV1PpcWPDPMANAPW/LdArPgJOQexJSoJpCUmLTL
FZfFNmz8qCtjhZzIMAaakWgTKDdz6DSGtO4EzUHMImylaehijgpxqM0F5lXPwy/MmeE9itL7qARx
WLhP/nIPozAn5KQGh8g9HDh3Klz6UdK8NRn2dZcCoibb8o1kDMTpPhktHm9FgBs6MRt9ufD15B4h
nbRu8AsxhfRJkx0hVrzfJZ55m4J7LIPeoF68ud7eEU99VhrPjucGdjr3MXwYhpSQNtstHAI9h0sE
MwDzH3nBTcQNzDIx5D9Gye5QLuliEpz9LzWVt1LiRN6xYhYbX+vxGf7QYEavUOUqmgp89HxrnHhw
Q9qwO+uUE8FrtAYw3uBeUyO0Ah0hfSACa7ceh29M1OkHaxgV8kfBxKbe6Tv3DoztursQjkPaU8pb
UxUnS3ORXZrRUWh3eHR+QnCktECmF3+oR9HLChmn94YksgtYyATX8VrmrCpCZpJk/Xx6s9iG3OSt
rhiB5ZCCInQvMcca8lLXdAkW6uxLpSqens0uoEzKoRtSjM00NbpzCJOnE9qIexl+aBqWWMjnsf2c
Nx+P/9a3ED027Geg4qAcCCIZUVLzlq+IJoENwx3svbMXDy1OiXr7pXQ7oh01UaRKE2ck1l9A9yqA
K2x38aI0sNWtwxpDDGYa2PRttZu0WcMAfPVyusKlfaElrnj/CxF7RHpTYPcoIi0XJyrhSg1GsZdj
cY0ZGCSrtuqrw3eDBVOrBVlYtGPf8Jj1q8JuTGhAkv+dPa0cibIgIewGhip8LMxOydJNreIqCUN6
NTENl0KIInkoFv8H6XxuD6PGtHEnsynJIrlOyH+IRRx9qX8EQKGjN2XzN8HlwkzKZmwbpxa8egeL
/dQMLz0c72szPNNiHzo+TI2wsXqvp8J/kAiL4exghkP7yuvbmW9OfMjCpA+r8u2aQaAFzGUQa8ye
Yw7kGyEoFCBNc9QdWQIlon7/9gb/BMLRDWtSGId61ZnDmUSFynXTGXoja7hI7U3BX50F9gFbXbHk
MA3o4eNYOvTj1KHTQmGNi5DDQUDYdpNGn/D796j9YGfKHCzENiOScRyNI6/os6/OEZ3yeZDt+XRR
FLwVnoWeVRZxkPij83I9aJzoJsaAfKuopmO2i5Qu8I+L37EfB8Fm8EAJs6/3xYCCR3UD0/8xz0dQ
mi/Shm1m9mg40Ve+9qVw618whbYnMsv4osUHKUoxOB3lS4UFAapbIqpehjb7LFczH/w+nH03HomK
Z3KW9m9YJ/XR4qMhMg6vmpOY0Tw1zWRf008Gad28yWrVihC1sOh+3K4hqtVEftwUUb49a28xBttT
BghVand3j2maBCeLMNGZeKEn7VjSkaixqEbZuxn7jhsS2kmWhrwz+TCmEsYbeEJ9JQzXh6+fP1xN
47Ktt0314O28HErdtHPXPpcTOZYA0TsTqNkvgb9FMhx18O3bJ19QUiHKxyXa9ErD2aIbUrIrMS1P
VE94gM9rlHINJH7qjA68xZV+Qi5+Aeze28HpAVC2BAowWXIwGkoh4RkvgQPD6KFfhwCP3ed/ClMz
rR0E3tzz2OVSahF2plo9DdSC1DwG8i9FFwJjNzVKkb69J9xbQRHzI2njBcZsdiZb5PiT401E3ifK
18E501sTAdDs8IBNEPLKHSvlVUosOooO5FvJWpFPBefgdilBDVzc201lLDAkFq8B8yh+x8Y/RvaS
fX1isfGQjzlkcWnUMcZzWg30auP51q+Mpa1W3xsLvYrYySXpTbU0I9Bso4/0xKKW2r11bdrC5Y1S
LJGKppook2MoGp8HDfj3dWs/xwwnb/BwA6mISutwLAewV82IqvCAHlAwsJh+q7Zq2XQ0vXS40iSu
e9NOXlkXQ8c5j4rEIakFAPgwdAe6Qt8G8GLIoTCI6yKr/XE+PyA8Z/rBDF7JHdpGw47koOD7p5N0
oEdKjlVNl8TndKRMWJnUI9j6RuC2YjVH3nzvaLGDjlmQhheIEg7W1yd4HmtPBFD7WggVIgdsVXBX
Nzy8ZZg7pKGIbN7ghWLpTUu2B7rRqXioKh2hAhRxP/nNdNehazasyhoHKX2IL1vbGRfsAi2SZPV/
DqtDsuGEMOGzfkfsAUef6ifsNe/rrsvGfNizJxP4epDDNs2Zw4Ldkxb+1KQHlThJkRSwPgtjNDFn
P6ELlXrtaE+Sdto7E4eH1iMsTZ47asgJUV3hkW+XByL80/En9bLpLL0athsY7LLE2HYeCpzCgjR8
Vgjq7fSj51YlZWqiFi0ZPl2hWwNLJ1msOnwD8lshnekZ/8MyeJ4zVq8jRD+Bx+X8jXstC3+u8GuN
HJ9xBwy7rmg5ew269BE+v9U0uw5s7jalWKZiIcOK8lcmt2ntshMdjTvtts2tK93/QwuhS27toN19
L1A86x4rNPLkAsXk9H1yGsDr5euJeg5A620AZE1KJAkMl4ccaL+JT2qYWwJtWI7KAzcGfQV04koL
Hf8B/2xGvbtb2iFW0CNMEWgBLrBjOiQ+LxHhJZSRb7n5OwVcmEJVkPkY2gGMpR+qdBDC8gG/bNKk
t6D+FQcr52WGzI3fuxXa1UpY9GjBRDEejUv6xKbSYmS0MSiG40vZlCp8i0kJLpQtOgkGAtcGFApN
KpF9o5cfah4q8XkkzHSegLr04iwpsHpUJu45d3oU7wlXVK+RFcxs5Pif6xLO4SD0v95dHe3ZBYck
Sv7PBBKalRf2p9KGSwdgX0f6ZTMxfbaYhOvHJ+icJlhbvLa8ImKzyO9k+fVW7RfTqjy7hI7BnVkY
XjhtAKwxselcxjhLThnRz4CXx8ndRYU/YvEg86z4+yh+8V0TcIZ5WYDzWOpWBqU294ZFrxYXN5RR
NwjDP/sw6KowHkXNKVi9iPFhlhZcYtIBMDGl6I1o8yKoK2fToOuslo8In0PRjevajyq3QybDPyBe
RAE7S1g0+eIHNCbf0VgKNKT4+TVl3WiLhtH96He3SxMKFFi03qdYEh7VuORI0ffiKG0/ly4bMjk4
FTQ4U/C04jgEg25pw+f+hWrP4427EwjodfwKJ7DufJL9/+M8oRzMZQKRQPAkBoVlbpFCiMaGA2rj
eXV3vtJR2V5/uujz7B0Nba/FS7S5o/vKzM7RtaxY2bkiIJVnsE+SFpETNXMUpvh3FU4MJe0F1O5W
yy2YPYLu5qZTYAcLJ8atx2BcJPIcqBCTUDWhPKNDovp8+9zDw6yQ1uD78nqnb6VvfzPWggAwOmlj
om2J1ktw8txIUL/OD4izg+g84HgbIoyzi9pjEEmr4oIQCkhnkHu7pRofKFMn+hweVq26TpzqK+cs
izFV21GEslILpqGl3RDkLtFg0QZuR8+ph5cTbwh+3b80P8+PQfiXerDDydbJLYbyZmrNncVepotz
5a9X01c5d+1ry9/deshbHFlwq7oC3iLQPduYk22NI5Jx6ufU1sqehTVfvoQAZNMqaZVCCXM2PFjF
SisbHhL3NDdu0xgvvIcMBQXJyT0H3FZtfCUJ6BbawOHLT+owRRSYheqtJ2OU63ggqvMS+5eWL40f
1YfVDXyDb7jYkNvfU3dGthlW7c5zMYYQwWN3MMiPVCGZ0g9hh5jZZu4ERCpKi+gYsRmB9DWfhK0T
BqqeFjKR2aRUSyn9eOJuxPoHuRpc2pa705rlIHTnx8+wKiMRpUrDBnbOfC0XP4g+Dddvm0KaEUrZ
9p7BQ2ejeKKXA1QWmQNDlVxL2fQlr1fU33mTn3hxEoI3R07dYu6y3PObYOkjFIRLoZUMPoCszfKu
ShCQFqrAIkJI0zwwydFUrUlHME2wDXTfa5MXyf95kzp6Xf4yOP/arZ6lcW5CdzeRsK9Q6uY14OBP
EdD6OPxC0JnLx3XW5qmoNq2L/6Z1TwZMGtE4HJCwkglKyR6Mvc3hmLygy6wccD4cSS/C97RXrpt2
47HqxR2v5AIDiuLTky26KQpxY6Tv7kXFkaPVO8oNvKxrjau60oNyEUU+xaMIZnU6uiH5WGQjQY54
vF6xkjXnDskqVlUv/tRxhsaY6lfMLm/GuK5ZYRaeO5OUAV+4PmQab1XmCE/LImi+bcPEpse3yCZW
0sX73P1VqJBUxvRo8F2FV+Mon+T0k8/cyNDsFlIo2KeVN/1VYub+o7Rqj1Pg0ARDKPqKF+xKA7Tg
Qt0wtVUXrvEL3lSFHJDgjpJIc8+dOgx5kwatrd2eIR23WRyZYp2FeRYCyaJrEVidgBUsUdhc1zLn
+giuMQq7LUoRVO707yMUYCG6Nqk/HRqvDpoIy3iUb1rlf5qwv9+JgOq5mwDWWULVdVKq/esKmm6S
tj7EyOWSHutQ5b3mOijWnywM74WqgxjhVAiK2x6rrVmJi5cr61ehSXrJM9hSkKvWau/R3tUKa3sq
ujAM0maPZNY/v098eoPUJnLrQ1yeqX/9irOsEtC33+3HpylZKwmFwyalBo4lH7dGw5YiZA6aE7vO
gGyQoHxwbe9CXQMUjt0nhuJUpq5QddevnXx1bjyeY3nXlyDHYecLTe/rpQcLafitdiX93wpyHjaY
R6hEZ2BZSsU3baJSeJhonZz4aN++6zqxrk4rjN9SIbYXJhaZ6GU4Bf7ggVSnSXxVO5gis/+MSfyL
HYJCxq0lY9oQKHRgmpCsXUOrEQg/osB4prDmisdzAOC2s5ACHgDbPOZX0B5/Q+T+uD3rQ22TIuNq
wRz8pzgGQcpSgnrPytCPisQrIUms6y+Puc9SkOfiqWaN1Jd3M7yElTIUDu1qx1U2irbhHLfw4Rh9
7bMku/viY60c5HhVhGQC3wawoekoR79tu9ph/cpoiWlC+M6nZ0NWKzKhdweTqoo4G3z2H8TJJH6q
kE1YwYSPiloHrHYUeEZnhWqWDRg3Ueh8gsr13J36dv7fBoslMEEdgPhW19eSiOmH9M8uGdOzG+90
20PAahgYcj7YhWIXcWzoOEfKzhh2Q31Nwon3AWPDN703JFakQJTStIm/4lU5iYhwMT3CHPcdOdU5
AU6+pp/ZMCyBeMp5i0Xq7Zkdh1Xau2hpw6lQh0fYZ2SgJospAFTRe4q7ZKKUqYpM79YpEMsnuigr
hsqst76GsN733fyeCiLVv+vWBEZTMopCOtGIYTl79qPXv3Sg+IIrxlqjSKH3taKNCBkaU/YK1jFA
XoM+Gr3qDvwapOW5cWU6WlJ2oS4K3dk/+oGrrPkmYjQFXkrE9W7IKvovPYXoyec+z77PYc+juXC7
XOcgYbO7jw9wZ33MA3YDjRU/bSu/I+mOEZiFNsAoaOnowlpCRtqYopmHZRC9YG58nxpBA4mlMdMA
FomnvFDD94H3WAwiuDP58fdZ5JxE/DLPSMXFddGjfYvkjm46TGho/llcelBj1v0TH+8TfeLo/Aie
d+Qm/Uf2rD/fqwDRnUlkk6/sIgX+w6wijtrS+0/uFL98gpG2xP7g7410+E77T1Auu7DY8knGft3B
HyzSonsfNShFOWBwuvRWhgZ3HUW8gmkouZ2N5VzzwuvS5TEYQwEg8JHaVMfhVcgxOsUQa4aFE9QI
3jasCJnmRG2DdU+SQzwZCblogTKdTKubGhrpXSHAI2p5zn/ipvgX2fyGcFTA7b1fpUuR3rrjSPbZ
NlscwbzpvtFc2giegmqhQqcvWH3KjXEerFiYWy10OUP5/aiHMUttEkoGeVC5OOrFQ2K2V6pbukQ2
+FWORxu4om87ElSM/yd4B6WBQxTP2HEmWhCoPtZSHwZFuDyqex5qs1O4jO8c0ej6Mk7fkPm8kH49
Z4YYTIEzLz+ZvLx3odGCkpzD6+unoN692nMRYSI91vNirtI8QclqwEGqio4P9+PEaHQdaVmeYHqw
c0kLOxanfLr0AWSAF0COGoOWh9B+3cZOcif1N0k7B+FKxLqUqLjZrfVBea8rfQ26xIN7+NB4q/wi
7W7hRqf/x05z88S744uo+8nL6BcZxjSj/c6X/83E9A6psPGcNKFllaPREivLfk1hx5dMij71/j13
vSXF56ula1b3aHhAjY0vLS+r4pbxd8LvCu61WgvRCtvxqYiOYcd6ZM8ao8kBSeBFnw6TlH1k0J9j
if8NpJkAR9zWwHf5fvyuFkR2m9ODKUcGvTmUy00suX4OfsDynEBR3+EOCDKVRESEi13jPkdixNeU
tdY2QWWNZks+L89TnidN6YMoVhTt2Qm3NZ/XrdyqlXdTUagpILyaEZDGbIHH09SMALJajc3WACgl
T9NNET2Uwrr8E1FjVSfPMVHV2Q1OGx3kIh3lSKlSPu7rfrtiCTOLS63MqeBp/GyBt2PORGFI6cIg
zUC4E497eRpzICfxlE4ruKWP1cdHQR0w7TIflWEtVYHmFSad2wouFEJ1URt40clSiBY8cMfN+z+r
CvyL4d+6dmH9hZBunYn4tmZJpiwYzzUR5ArDLRQ5lOq0CRPlXHDZevwMMr1IzxPe9LLBoivt4L6g
rQZ/+UMTvY8J+0jBjP8R5TGos6l/rUK6kzHYr3tbwputhzUdgLvVfKFzPbQ9vubyHHjwv2TgutNz
EAbKSpNPgn/xpZk4Ue6Gm+hX/U3xKAjJWR0rotR3lQPEJQEM3lSFP06W8vM4s8b+sI59Ao9Wh+IG
79WP12iY6oVcJnqfaJ05HJ7ycUFs/syTeTADjnpqy6dsf3vK86fyShCFWIc2oaNOUhCYAqzR06SS
+7bZjBvwP+skgWNG9eQQkR/+mFbtxxlZAoeABNAoYnm8RY4uJJQiPftBUG7XQ4WgpGDeVaAjaG9f
zpkg6O6cNBD7z8rcMxvg/JI9PmlhxoeEF77soH7ClQJNnZze6LLITBX7PGQazjJY4Dm2G83U8Z0u
RwMWKhzTapzZhUoAd2kXU5x7irmOLw/OYUY0UIJcDFwjWQ5bsmUcsGd3Is6nabEdzJCO0iUyNaTV
8zy6ObzwlD8zKYTRVyeJDt3BCAYD2k205sfl0Yt+a8UVb4KBaXel9ipLILPTpauuG06fG98GAIeI
Mf6OYLXNTXa9mX2KhgvCcx8giUw+snH+BnZCzQXb9oPXDCm7W9zqgi1whUX1h8IpDeIg67Rqahde
u0um3kBwOHEPQMKKOTq7gHVQ6OK+2PN2oW/D2gmIo8KLkqLixJxNp6JzU1Kb/2bnxTDQ4N9cAcOV
9Bs9g2mN5naNMRbSEE2M/zkQahmGbenwyv2hajq6h79uvWFU5Rc/4ZaTkJgcTgiIKgeET70Wbl4k
osJhFeJA8f88leLS0jr+fW17MWaYf7x0OKiuVpJOui0yx4xuPwK2khcJGjJYkQ9bdFbqoCxZNkvk
7yFW+O2Ie+vjGC1EZiXa5qODv7MazG5iaaOon0Np36mCMwUYXQVmCEjsRdjEsce6IVr2uuaBcc39
LW8BpiF79mr2JyPKe1KaDuANp9BjcPw/o0d9vzeZa1AOYg56IKhwPgaZ4ULJyscAjJrSXho8QgT8
2Z631ExKjmYI4KkV+HxXgHpsd4mYJvlmh3+BXpvhmN3ysLP7LnIp5SYAxreq+xz+4BBO6/Jerfx/
GKCrBQD2k2sGFKsUXKW2tvVAqQGkQDZjwIP2xmv80yC955usZSf1YRyJfVKrQbp0I+BoWePcP+H3
vxhAoXMywZkOPUL3p8Tmdl7bi7tT/akDMnbQ5QzLceTCwP/Q9Q/ZYAsajJGgoxqD8I+QQNDUT2Cn
I0HVYFOVtssHC2hrCr17Wz1iuwgf1307VdAGZ6uALDIF+4yXaCPmsVKmcgcjiZvSlUwrJ1HoQxJz
2vvs7zgyhBeDJvTDAYjLy/q2amqSEDWQh4JTf0+dGweDqF8YcFRiJioT+PNo2oNlINUlHNaguZcR
tHvpo/JMANYsy15BZAyPWuO/b8jR9uOSQzmhYJeH7HzvAh7nwiqDoc+4bYOaORVaGw9MSD+7TLdO
b3fxum9qGoE+zLirLN2kBTZhmiDidJnKo/4gW3HTGA69E2HSsg4dV2t0lzvU+peTHlQcpqb1tKW/
+7nm4e3QBkyVorHzeRpA+BIdy6N6UQeWJGap738vjoIUG6Vrn76gUpKk5p41QNMWeU678kbL5wiM
zyN+7mHGUSjuM2koo49X9Bdwzr/jkehvB/uturvoxIJpim6inqpteyiisJsULkdgKQAaBxqw7EBB
aox75D4/naGMjNjXiLAK21lfI8z+rK2OcZeZEWCap9YKOnwBkvOnyVsr8+sbxuJpRJAu/DvD+/mJ
3s8DVFMWArgWlemF8hO/Q8pd5/kfh+ukJZbs+TNGvZQlHBgVcHkVK5niMMW74efkLAy/vfgK97DU
8gKs0H3DL8RUBWGyIbhFszuS3OQByMVUxHv4QDwJGVnuHdqmdotUymubHLuvnDwYMRDrTDihrFiw
EdpXc3VUxpr1+h+C5M4k2s9lHUzxowI4MJOqN0yubG6FuYhkcWaQtsJBXfPoilb+EEmSYhs3g6pO
c9Huo0nR7FysyAsIXZKjjiVE0NPy7chChdmD+B+4JRfGkc1FqsYmWMSj9RH/Zvge13PA0sE/PPdZ
HKSK1anzymHxXtmfaaq7PxNMbw+LPBmW/iq+zaqivT34B5zp4BwqtGN8PCYd7lcj+WL0+R96qX9n
E962BLZnkz/7K5sb/0bUxil7YG6ZDwSPFbLdqNl2frwJRhxH3CWu7WyZ1z2vtUl2/6t//4lvV6Q2
ZeHbJEPtCmu6FwkZjlm8zwh0ELoQuNMSLqngNPLeF3sINCsZsvSBcyaZdYRGEaGP6cxGytMAn2w9
nsL3PQzINWhfOzCVtEtTTgUNrNiK58Pl6VOjyVy+xCrCLApO4JlfwZsTDCf2CrskYirZP0xe1GMS
wyhe2IKryWiFRKP+LOp7cq/kd8n8A6t2p89ZLxeilXyEczk5CutgJHVyHBx/5NowCUvN7+AfSQll
KnVIm17X4ifmPNdj8HJFB14izKKgvY3hb5VK52aBE5K+PQa9bpwAOIbooqVIp2COdJnbEo2XTXTv
twpdMi4O1+G7WyRh8VzyayJsn0H8JpFZjgp6aDgOgiBqsBZe+j5ZHC1ZJ96DfrEjZZmim1bGU/Sk
c8fri+UeNX+hKI7b323LrBOsoPOlQcLrAQsyYJQTryrENgqc4bREBm4fcswEDxi4z0f17j3dUxjb
uUz8PM4mmUSGOTrc7TkkShbVsFlad0rhH/n67ZrElZzW/GyFHjUuefZDGjWKqiBiUOSRLJqJlAs8
SF92x7luPHqrGG7uMpE4U3HkUc6XmDX1YJvp1zQXx+Rg5afVgHUKXTYzoRJ43Y0ciUQev8fv8IJf
IVUSLdmmGGt0sKK1dcnES5UcasqmqW/pnsHPbo6RuIWpb+CcMahGugatkvS/UoPnBXjZhUHySstf
WH+o7KfmYchaN2vxHipCYRFzQOmHyvf8qWN2JL7k6fqdydNEZqjucr0BIW90OlFSlWmvPo8m9i6e
PqURYqz+TtXseUidJ/cd20AvlVTQhxlVUDKydZ5Qpm7PHdecCnU0glEEYGEs3PgrmnP8m9N8l4sc
EOq1CFPPu0ADeq01yxqTSp9F96AsExUn31g2zfE7LjJ6ouN12BRuoz0HF3RLyEoP+DB0hV0R2gdQ
JWmW6RRVH1waqjoyjJXRSEtU58BpHyr9ut4NAAEyfK2v7UVxUzMMu1j2Zjwa7s/oab2R8hNUEFrG
OvzBSCAnvjVdNcSxSotZiYTcZ/HB1AEzHQOndQKIYzNF7tWA5yR5OMvb4etBoyF3ukcJOzrXS/XS
pT8JBEBHljyW3VYWXi4AXJ8JDOUJH+g7srjDHbqGiDhos55KGMvfWkoEnrNfxeyu7UGTotWmGOQY
aznIigAY/5bam1RyZsj1DdsZEcr7dVjpxth75gb3cv5v9RwnRykL9c/BSzrlH3RnMYhE4BhEMXUS
DpQIEqPyzPBfFQHE7IDGNKuoTacswFIA5hkhFlZ1+Sujl6peL7I29U2ICQK1j1PFcP1DnNWgloVT
Z1nGBY2Zu55zva1TulRYiosID5ad0jWxmWXEx4hB5R6VREaZLHHNMxopd2ZvOWlVlNGDmX45b13q
WuTBJDMlbS77tuFyyTbqZQ5f+Uk9bxzgu8gU6oV50EPNbj1w8GCOlv5fNw2br/71CKQcu7JOlmcL
4nxMp3iZ7nA1Pm5i6UZRMQnybJG0wMTDAjmHC1SUQnMN6sl/5BLnD5eXyhZwynoN1iriou9zopJV
Rv9N6m4jMGG6EgkGBdx/i5iMr6NNiT5aqRfNr1kJkEP+kg2L2k3k0Zwu9H4SvN+0c0+SSr+BklNf
fookA5KVtGTTRwDoUjK2vJyhk/mi8Rs10ykLpiaAuB/7rwKFCiVXEC2e5yCpQnkAMM+3JbepWHiQ
QHId/3lJKPPk0IFOr/7zSlhCybWORC0tnysJha5FqOYqUMqxIuOoynlohAFRIV8hM71lNubNV+WD
ru6EHKJ68Tit5Lnkzn0/U/XQTylzauv4omM7D4xKjB2ad1cr0XKL0MlNnDDJRl0tPY8BDNMxVhgX
qq3ej0xNedUoZBhpWGO7fK0T602YW0/JBez3nodrBdLJP6MGOkDX/KzLm4p8TMaiPlWN5P1a7Zss
5AGJu20Xf1uMbilGDB2muDmiHTAH71ad+NWT34WPTP3KbxxsWtSQmwsz5fB/NyveHD0gQ8E71Ltw
W/MPz8RpYPdwySWUKaCErJALot9ahaUgA1Q7Ay2Iuo8HweKp4wjFT6hgmcvbQP0OX51WU3dBkce2
yl43tC6dZaLy+I+65KHuTMeggF5mBc0LkqPp2Zg8y6a9+UGD0cKR/p/vMU7WE8B4v1idep9QwOq3
v2y2DKaFe9IAc165syl/OyMqubWVrN4eZ4WAoFSLi+rMQRLqK0mfOf9l9zSYOC4Qd7OJfm8K4oaI
9ooSpgGtJUQvn4gJLKYgl/VCw3Gmq9Xlp3DL2rObdQcRUGHqYZ42tn9UM+NNMqxiIWgcJnWDRfQB
CEfD52HOPsTcVF3LoqjxwEHGbj4HR8XobNJR9i7cMsnMa66SaXTCz1mNheso5QafifmjDhaEOhj7
u4pFoXMBERw7/a1fvSQ3stZ4driOIQp/ASTJBQEs1mFg2pKOHXZWnOdDYXMgaSbqZBckAHXdAKyG
cQ88MeTyAT5nSRZpwVHrG0evVkLLCcK4CT6R54tbYuUqzpMSv4TDp/Fmu0ev5lF9MF5iWUo4UErB
rDNFEct7BdxnPKN1dQmjnYjftERicvAZJYuuio6MLaM2o06sWHPfH9eH+glv0aonK6Y46tjqmLgO
KBMnON9hXGNqrA7Em/dMT4yFXu2DVL7oTDnOiNGCQymEHJKdBsGSL0Fs7BEiKh68QweTJo9ZZ+bZ
+0+tu0xuJ02JzlrNCBwuLzuKKrPwDxZTcbcvI6r6eZrn+t+afaavALwLF9snr2EBEajxBhTUokr0
pYR3xllMtE1QGQ1bciEgYYiIktt/hdgs3ylNpEur1Sau5SnBoTZUedDl8ODPCzrmrqoludXW66FV
aJwRoSnbgd0EgI5srlbxz93w8J7U0xyMJXCFr40h+8y+ie+ANTK+G0zHdUwBRXUyioKjIwhaWeSv
wIMNYiZtDFOQD1G59kHUb6jgRjb/y4IiIGGR4Q+g5S5vXBPqS6oGXKGTeLvXe/udhAXGVGsHDfea
lP+OGnP8KO23gdw/rGHvv8YX/TPHyUNPF8z3OT+/lePUZbsNJEiQtkyoNb3p/KLxNShxCvn73qI/
3bE7+TfJFngASbJfFPsHW50DalqpskqFsYdnhrAhCDC4Q/0rjNr8buf+5ocB1npfX2VFO3whQNy6
vlpLg6UfdLB4M/yl68vGoVjH4K3TIYDaySFsQQms8chqYYP13z6eVt0UqCwPmfuImuzIfsgkRqSd
s4NY47PHuI3V+ZrQWw1fZyuD0ijd/RfbaoADSX0R+QYxIwlvRSiearFIHVvUPrzluvRp4YxcT6VB
BQfkrW4A8sCQrVb/Xd7beQFvXE5gwXh+pkmFMIGHJZOmNg9EFeFkaTPaoLj6l/cdEoKlPneUMhYc
oyf6mg+7fXXGX0YO3Z9Ztzi6GIozBMjRb/2KQ774WNwos6wU2ra0O4gq79C8B3oPmqquhrbUscb6
w22DFe/Gd2sqFUeYpUzsJqh7KTj23+McKz4VeareKMZMGnYu9fGge5YdF5BdczyyHsQTy+XO8S4q
eRG0daNM+dNVvrk5xExj9Zj2q4OHVc12JMV6PthB+Tb2Bjw8dpwauwNhbmDSwLraeAxt6YD7B4na
tYOdZY1W1ndgCIKa2bloEvkGvMbBiuJn1/XvzNfxUDM+ABecPrTNZAwHiqTEvFHEpwo4YY6+z461
UC+p6pS3SuSIavCdU280Wla9JdMmBMECK7sM5jVndQ+CX7VFlVSf4ZhFTujI1pN8S5m2Qo867a0Y
o6QK/r5lmsedYrHSHbnkNcl7npepw8Tfo0hHEOd7HpnxctIdrz3aoibBAbsl/2X5ysZ9CDMG9KdE
t6bHaXMjr1r7m1p5eL8bQECs8BxYASt75r4PY8zCsNtc+C5aCwwxcSGqgf8+DKZFDht1U3c7MMV1
JpXjUYYBygI0pmMrhD+qCxpAY+rhHqrFlwV4TidffqMkZLBT2GGFkmB4DE2JQsSEgLdN+hWMHrOV
J/Wsr7b1DHgdkjLxpKhJ/OBIsy6b34dwYSbuhoj/DAn33R2Q8RwQlsFSLgEVw0JIhlPe/3rKuZvA
Wmcfig+yFbEydb5i9V3cTg/m975fRWZrlVVGMTwCbuLDDJMlkrssf+44NP1r1DpTPJCrGg+6NGNl
FphPIeGMciijDPcp5RR0A4W/3/Flc3dQHxFiLfw7AUD6btSoxz/93dg+kUfUaaMAneNeeVfn2n14
o8SkUgjgofJCkskZZcFF6P25i90O3LXSQJvbMu+LHH7L+6kBxVIOSUw5c6dNg8Q8p5RDGRdF6jwL
mGwS3XApiaOmkQa+qhaQOeLDWpBEZQiE75dW/dn1wOhcsVWrrVM9McwhgxxBJ3PYuN5nqG/IshAE
5Z3w3UNEM7xWHbG0D1YtCHs5eRAErAPjocCCjBHibuiu9JuByUErPOt6RJblvlDyHuDzf42W414+
09ZYjA3ASq24+3aZvdlNGM+0BvFLno5kgVy/Jh/6LDgYiwnE2Dh2iWLhmvJwxfJscIkLjoEXJ1L6
cm1x/d3shaS7XX0J1nqUOfyhwm62w0TWi6zld+FSJL6n11sNLRmJO19AGBtPJ1AwBcj844+cPHCZ
1fW3mddreffIF2OMDSSlrwI4NMHmuLH3gxuJ/Ae4qOzuK4X0NxwAbqrlQealu/pR40R0rF+FIN0i
CuH7SD4cT9BJkr7Ado7p88mmIhwa3VwTBeb4mkECKVCySLabESsI7sTJzNZb+R+8TDMVMqbpIeij
bweK5N6Vd0nJYkZFvr4oOBKNJNQxDOCg7uPoCD9w8JThhAt00D6SkcC+0qMpztNkyZFSEjkC9A/B
Ip+INMXiKF21putpI27adUWXkGEJ4VzaMZas7ynfK5XvMZ4gmWQNepvAE8+LC8WmKBfCw25eTJdx
RKnwLVn60BrK82D2VDcAplPb6Pwu5NutkG57JMYkMQcKedYVMJjQVfPlTLtZEwZQrBl5pnXvRPqv
R8/5HNhh6/Fs+pocRm4RKlrhw4VHaU45xb6NuVzVEv8pUXTIebnOD3tWobLGskUT2HBPPJ4d+txz
utS/WdlfmbugCdCgtI3LYqA0Zse8IhRm8NFCQJCcb7yeLjyjIXvJmGs35wAhWX+QQpef6Oy7+Z7X
jN0E8o2RalhrY36LIlv8dzm+F48owRI4CMN5uFW4+FYDuPrL53gkIfT8dD9528/juqDnwd2koyvT
8TiUt6ND1RsLs8ifVKgnFB0RJxF87q0l2PArE98ehZiVfi77yBJweAl0kCmJS2hO5wsds486He+q
FmrtD043fRtyNaHspf4/FHnYzeP6mAD8JsBeUNINZkZMW0y7A2xWByN53X0CZaTlj5fSiOFbqLYo
cITljKMMME0b0B27ZiITh5pPGw61LkFymRwydisS/J28bijdUkU9q1BYlCIE9B4zzGbQloK1lWST
NAt3sfwtddk/RK+MDIeHn0iYnI8le9z46buxQl0Fwrh8p4U50my0bU+3qaRG1jpgnv9IIghf/jYb
HNePGaHN7LbrKbsa4fAp494d3wnh7ldHtajFCaM0qzFyNKv8QRWLxBp5E0Vfenn4YNXumkW8jM1p
VR0foBM3bB0n/HFq3Fh99d3mnhftKxbOvNclZ3OHt8/sVOTL64bX9yDhRDkSZrIUgfNBou36Q/44
nsKYLEzd5PdE/jRCqfaEPc68VPWfvEGIywLf7gXP2HlYOneVHIT4Wn9PN1gKNnW8LHBkjpc7Tsmk
EyR/MYiHeYf+9bpMVoF57Que5u6TQ09KVVGxQ1kYARDa5KQvDmg3OwbCyN0icSs5LrbbP2aLHBPz
sCiILVGfbYMmrkco94UUNZjNB0J+lr8cV3fdrzdv4Q/i+Q8qri4hDulxlkgDklgeAPBX+o69tzrn
s5QeU0B4aLAIrT1jod65w/97sbAU1UoIUhE6qzaXqFQK4+M4oNy/hLvdNt6YznRwLvxPar2gwikf
Ntfgb0ONHDOq0OxrRdh+wZrzGfo9YebxWSf2qkNoMToNibvPmtNCSOFrcUOJGb6g1HiHZSrcxVVK
LavRchhQisWCRtaGvb9E0SX5JI6/gdHu85bgElTM6pcTdLqmMfQefihpgmGFmmKa+TEvUH/SHUv2
5Vzaqq2IcdUDkpAn27YAiTCTywm0o8XMSlTmJdukKlP6zwBsMmpZVwETqbjQ+qifFyAkUMIyNJ1A
8RbKbfIcH5GthqF03uRMjnjQlWP7mGyLkhWeuBLPh8RNaj8sFxM6NGz7onz2wpta9WzXlXJSa4Ar
pr/X1vT/5zvZztJLcnOMlGPycUlzjKQA8Wc0zYSg4hOPrMzTVDed+tzbNTlV/CQqLWE5sC9G8mdr
0llQBjcy7q0z/3F//HVKktMuMor808QgQHyITizlLFoLD5mnXR0u41HSh2hbQk1fnhtYPtl0Vv0K
vc7M468EA9tCZ8o5WDKZyP/9v6tOpF7CFHcCcjCBFOrf9bWH2uIw7dTgbxWeJTi7Yw0gojc+fhGF
HdjSwOHluO9KIbN0iwsUcfwFUwmrR4UVhPhY0Qyt23oHUKgl+wFfNFFwHsOzr5o4M0gFVAz75KSo
9wg973xsavQc2PXUCM3aDbeBpD2SZN3GhIdGkqvOQwlFpb5E4B45hYHK7oAQh7v1R98saGvbYKhC
C50p7iUzgzMD3d5vWu0kOVlAFJgMho/uFQpjvxy7+sGyzHMe++obolkEAsmE/3Nnp9Bv68PHJzUu
LE46f8Ke0hRL5gshQf7ruMumsz+mwlOGkYmIVcDxeaYodj82YSucsEAkmIVBYEk2eoNThD2YLh9t
YPrGfLnKdJGUdUScnRWGI0gqqK1cT7etW50HTokwwYiml83qwRVZIB7FQSFYPqyfrh/V1UmF0NJf
IbL9X4E9xrI5nNhG76L6wFLSFzSg5XNBzzYR+qiPeVMI9dYaiX4ea5QRH9ltH+juYwgI1otRpWaf
uW2cQA/N/MxOmeutvCvuJDV9CR+98tuxV0mdZ1tJ8Q8XdLx/lCA8qRHLXkQWxXtnEqGghcB43ePm
Z6ZFGnRkSt8BZCQGmvJvUZrZ1uemTtyoJlRDLQUznYWcyUdXXApGMfCQMI1R8fSW+8ZgkLxZO/Ad
Hdx2KaqHNbwC/j3cLfW8jSRBuiTTpjNI5nZQhMyWks2usBXQq6C6Ajyj+mRmGlzUPuAK5FUTJ8Wv
PY+v5DdnUX7HW5xtnKnY3bhZt+AAL+N0fMWnmxVbQDQAUZPrykyf86IgWMH/JnFfJ0Cp+M0/B1Fq
kVJS5Tm+Wc7Q9zhxDHt3e7vZ0cyU7HuA4OGvlmAGqpHCNgeYtt5egsDIkqxWkRJqar2F9h/wAdHi
Y1RjAxshnC7wvP+JSPVEIg+a0uGyo1AxGdrBeMRH3rW1Ih+aGnzaY//RNPktgHxtHRCcXui7HAqh
r7sQ4hDggFhjamR9UMhUq33+xRW/7Y38YeRBoZ5M8KpxvggQESImTJRapLAz5BAAJQWwsEQoR6/Q
S2ZK+XiNRB2h2W6x1LRGgIZee4HlRGw/vmNz0Ry6HEOAKisFE7LvtDgRAxXrfHECpnpMUv6Eui21
SdWhWbOEDX4UIXN3180emGZ9PUvGaobafcYweB5S3Y+AzKp40/tLVlC5w3zP1l79vtGiYMhGhoSd
giaAOUMdT/0+EeH8QiklvlxuaHDefifRPxbcXnyxvElcwa5+O/Dss4CZFaM/Eu3ZLTqzd5S01icw
BL97M2dQALbjrDp80vpB+oOgF2JwWBHDcx0nezSHS30wTHl/cnpgVR9XvNQ1GYnTw4AH/DF0CoPN
9qf5Ua7BwZlIfT7gbDDSDz+lIY59RiBmb/g5j1ghcXJst3RYi+JP1Ji8uG95mf9JC4TF5idksUzO
lo0IzNdw1Oy2uXrXPFJNwT2Fpqhu2DCj4YBAcSYJD1Ov4cPqkTxj6xjcqvx0kKIYra6/Es8r0Kma
9e6fR7vbtL5FCgbr4f1qrtHS5wqUD8nlzRsqzu7rIu37s/l9LiAcqHPh9KBZk9tS2RN0UQRbQhEb
ddb/9I+9S1SHwr64pcXnqQKmgnj5JqdkJZ6VwS90uBI/m/mK93n9zIRG1RLVRMf9pFSfrlbdxTxZ
0HytuohY4BFGIQHzPW29ZERhaeak18ZLwP0gKp/4LxKVCV65I1Fihof8BFJl8k7TGk9QDfh77Wkg
giVKGFXQpHsPBDNgqsqYLaHm1fS5j7ltiawh54JMLA3j08FXIgYI9eHAxNOEtFHSHmvfMvqfOnlh
Tyqb9YHEKJbIJKw3KixcuHaCqbSn83X+Rr/N94wbHCE5XT1S8TwXnxXTOKUr6BBBGTQsvwhs50If
KdpRXFmFcJBfrVxrwXBFsIVNM6XS7QzDKDVggrFDweKOe2gqHPenwWcbLrehbqq2Td/qV7zY7+Hz
Tuil26lSHSGTHL1yQPOlVFblsGnrFK5fv2blAeHgUUjcNnDfdlsMOI4aJ4wfxPVF3qy9k4d+93KR
Uzk3Wi46Tv/FWQg+C6eGOqX3ja5ULU4tjC0HKriDVniE9LoK0innxvGEyw2VgEK6Qtu4NKc1WV+E
F5XbDt0YAlr71eREFia1w5F/CsIzvIg5fS5lrnWUsKCjc81zxa6TMi4zMEKBUuizxQ3HciDttA/r
PMQREBW0Gdi6BopU7/PksGWg+XB9eVcxl27BzoJFuqc2H9+AsjOwlOhUzGHeVHYf9gZ73gXShD6x
68Fx0WEE+LbQSwnPcOCsGh+R4ELOddGzA1CSvhDNqW/C7OHpTohsQWYpTqd4mNsERLzEW5IffQ8z
yNQ5HqfuPieyQGhxFIymBJZKN6u/HoEY01GsQ6jEjyFOKiU+ZrlYUj7mG70QhT1Rsx2W92vuzDrZ
wil2djwCyefwEg2harS5NWLxluKTQm3N3mbqwoVAFbhYxvTy2euNs4tSmyhqUTfOPBjzFU1skdDi
iO4dxqEQ8OxaqLIBEP6CHQ9n8LcRuRYsFUZi9ZD4MZwi5OmzCn86baWx/a27t7KR6Ws1C77bjXF/
dTPGy4gnI652amykIDDzuLVmV0rAjRskk4F2ZCF4G0BX2tO+d5Kea3NWV0bOvHt9B+xmpLhOW/NG
snhb2fqgA6thlSwO+zYds1QAgKW9r+CehoLdPihDef1ZTtf3S0M12p0aM2U9xKca+aaCMo9lBlLN
3mNbpWiswhgLfKAzJV5EEFZn4LejEVlIKRk7s1LJplUpPYHh9NsJpdlvRS3HrdbfHL3o2TCdK+CF
i72CqWIGS6JR2fqIEgXLJ5OMQypoLnytTZyjR/B0RZApVydtvy/AsUlzm+ye4+keZfFKuhfNJ95d
VNZfu8iNYuZ6L/OdKi0kZ68+Vak8RkY1oCxuQTD9ouvpxxATGLOMFYaTG2CNUDhpKSeh+/SIg4ul
OZiVA/JUk/Kh68gkaBofplGxIeWdiazdemS0eLFN7F/0a/V4opMi2fswwli816k9yGFyBldgfaxN
cGfmUAA34/Lz/puVd//SUwYaW1l+rmnMQ1Q2Xw0Z4UPztoYKn08vl4DHAOUR7l9NepPjhDfJyJty
jvj1kNgzcqEp1oU/+kOZQnafehgIpov+NxfqGuQds0x941OMkBj1p8gSsLjs7elDD+1lhiDjYryV
0uslZbjvn7Z8G30YWA0g6QK5MfoSFbClI9VuLZ3hi+pc8hxoPR5ObciKGN8/13QU8K2NKyqOccT4
YIU9zC/+0D6IWnr22o9X5ctIHieP/pS//y04EG38Al9SCyFKOYBAO7HqWSBVsRA0Y0NXy8YvWr7e
xoOpdXbl+og/g1GvkgVYIGlmYVRngprK0yZRmRWKfOBoMT/tSAXVXOzaVIUScnSb2LRSapl/dxoO
vBLNvHWEjcyLmRTOuaad0zRrK9zBdEi5k0r11ulLJPszFKgQwBT77YioVQ4YxAiLuDVRSQWVD/m+
yjlUc63TCHb03WG2NWUfi3QHMuRqvhMu2E58Hn635re9E0nPtFPFnhl/aZlkBNpWYPKUT9T4unkZ
ooodYkYFT8iydRGcrjCri0nTe0EPTgcRH2ZoKX9GjOuwtEjVKSIzaNtQj+xZoAi7kq2gc1hpwBWQ
bWi9kWe4dpAVBxz0TJR2OvJK49Grnk4FVaRrBTJkK8hqiYroWYEW0ZLlwz1xpUr3+JluAmvGCpcq
3DMFGUk+EehidG8RAt/cXOjkW5dYA9Lqj7nRWjqNdvRGZ1/sqqCU3Db+UGSR8+dfjwDC9P0dtI6x
WYrJ0SRH1cGZXlozlMKWaTheEGlbMaeEPNih3AdokjWUpKO/TfOnMtaZQCZ6y7l149oNB8Aq2Ubv
Q2fuDMU6CCn/r2O4x7WE3TaJsUhznZVl1kS0blQ/WN6wNdBa46GlpUsafZwzU60anZEBEi54YmCu
SCVFSVwEsOrqg8cUFCDVAyy5urFhA/csy0dUsi1S0IIGWaJUu5zV6c8j4oUklXZ05hZj5ImXVs3Y
CzQEyBSfLd6e/FolHwM2tLXRiUZLKKkYQrWN6SZNB91QbDq7uCzIQJ+ka9vfb7PdsjekmvtYrVxv
V6rHQJNyLMJy2gaYq/dGg6vG68URzcpQaSElu/HuDgq5IyGV8cFFhWCexv9hnjt4WFL6WA6erXbt
U8l39HsRVtyTP/LYMFreeN4tqD53pTZ95IAOGVQKw8uiPQAjd+iXJdt7USozZmrkNzZNZpmGYNQ7
+me6zQVTWMD1134+BS7NoB5ozbaiHM0NbgyZIQmdpy65zn087VgpdJ5yyTHvpJPnJejyRoN1byCq
lFhyjQJXyEVjF/WPyHkA0Cv5qiiNT27uBLj0n/E7f9+mUNt87FgwLKt7ghclr/FvkNYmDClraQ5T
qK/Xe6IcbgU+rSyBBiJ/t0QabCkATBPf7+hj7J+N+nU6hGoUJZMHcGsiIyR2806Ipe4eeWrVKeun
UmlkDsH2y1NHM41YZqi5Lwul9kJzzIFNyHlL+E6mL8VD8Z3pxICY/2gTIiNf5KmtBFQkp4PfQNti
solLmLNHt2xubsNZ3tCoW/VcTJCiUO35YlLqwltJsV7g7PNXNR8F8TGDJRgKSbRFKJlpasFEn3qE
+Jt6+sey78tF62RVTKzZKFP3Ktx1E/47iGJ4NMFK7dZqQBc1OTmPwcHvmXnuvQD8eHH8ZS6GRmgO
tAInnjMY5tvD9Ydif/2y2USzkRptW1kkEzrMg/i7p5DWatog4/y5YV7/Zlu7uN0uFCaXWXHOWFrc
CyadRHtGpvw9WqpLc/PQPonri2ibbp1WA+5FALFEsmxJPS5EYHFlV/gwRD4poBW77NgRzNiWyTRh
y9xucznDgPlpSpRnKVIJKmrrkutpTy277vMxQ+pdBDAZTvIKyJuaNJk7UIvznKp8StFoRmO67yFT
WlBIGJJbFe5ZquVecFUeWEGV1/VmaUEKM+jJRmHOQFHCQ2XjCSKP6p0/fG7a1+uYlBePWUEwX1B/
h/yioSpBFEVy0OYyazlCZGqXskd6nA4qd3HYK/G0DL9gybnXBkWkgM4gozkNLPETFIiVSwdypVaB
rkAq8cgVdgj+K3K1T6P5qrZjx7ZR/hNWwJZy1ZsW7gTqImcMqzshMKdK3DPF7tp534v4AjBGXjNm
M6v5OVTIksXmlkpmwWXWNweGPjx2mv5WrsZ2sdQWYuUA9MmwltsfKfUcbqay/TQcr8vviLoxB8G+
f8YmfI6syBcD1HLkPDIkdDF9gRdsvsonW2lozti+a2Mari0mya1a1mwGJHS/NipJO+CJcvHPZDt8
+9ahnycFqWH8kpmZWhtQJk0toD0VMOZchyWO4RamtgDmA/THfHD+vuKWImfkjmRyT6+jCmeI+Lk2
9dhar6QtV5Ddrt8fIi2M0N+Fl75QfRWyO/vQaSd2IZJAB4qNi8ccyfSqiSyMXDaOVPYsqSHkSUZZ
/kguw9Q02/FsLbPZqbmwIJ5tecAQmqTz4h3OzFDvLhGR/GEjpZ2dMbA+uxg1uqMVGnD76PX7J29J
BGhYMalsouUkoXkNT6hu8Q/ASbTfxIp7EcxSz111pIjhtnJGeY3nxeH2rUADE3uG08UXISA/joq7
LhXx7j1C5+w7VbA/rEpdlKy7nDJ6mwoQcU4gs+71rECpZ9o7WjKB5ciyq7oYoG2tooBA0QvZ0DEW
2DhCZxjfGqizyRgF9pJLuq0flUzBwx7vcY7sMnucOMirA8Ucyzv6XJ3XdR7JUbVTz7N2WTybvYEc
3acppnL4TCzg2v+Bwo0fXGQzNVh0joUxG8yRyfS2zOuhfrGbjmbGF20omPl35DF9wZWaaQN1f0BK
518XdROo4opDG2ufjFQ/ysrNjy8vuxtL/StaXNfemArh92HZQ5q9ZTD06ImET5kZXP0H4oyt9KK9
QqIHrvHoonHELFe9rPYLonmv0jgKiQk/SKLqIXlWiGu1tXuNTovcOgF5cCvvT8gY3HyRvEUvLwMG
hPfdRSfLtR17Lv8JUtQZO75ogKwYRY2IfKFjz4mGR1c6N/lrmn9uaO6vT57peY/Y8XzgjWbS16DS
QCWexfu+h97raU1jyDDI+RWXxlh/fy/E6qvRqmb1eGLEzmN0EhV3J+dfOWUvS+pvtm6C0r7CnJGc
LdnC5bjBLakYG8LwSsRfh7Q1ZTwRlmKfHa3yV8cWUqR+GcrIgS9dP+jv+LxRuQB4MOzYgf/YThF6
VjPeyXrO2f8V4YtrO7Dc1uFk6D0CjHIyQlZ41urkBCTTg/g5Aop8Z62OJQ32LwnxVgGpRVNXbYcJ
JHTaIMmXC//bsM0/OwnGV8nCetCfc6dsIBbkaFeCBxmual61coF1JWQXAli6qIbf69vXNxiK2bGQ
6Ct+2j7T1jzxOhRGhYjc5zOLURkZyx9Yv+qgO3/1Xs9tzJbtw3iHWVKMCihDPFFS/DmZBtLr2+LL
LqRXi//RlPkgpPKPImkK1dVFH3VHUtKnUP/BI//HJ9qiC698r3Mhoao9c2g3TLf3TkPznOU7L5TG
7AMHk+XTNn/o6P/RTw6ZhpVZyQw7xHUrbQOD9yHPJqk+WrnGd1GMGxCKJRsFv5PiD1sARmdWU4Hi
3yz17mOsnsSoJgd3mPkgrWss2LZokas30yUYGbJDx1rrJL89rF1h/yI4Kmy4wO0b4DzQEJx4/eWw
UuYisRI=

`protect end_protected

