��/  ��Q(���]G%�B�C��G�1�*�$�^�Z��%�������[�Wq�~`�	v�.@s�Yꥱ��+[q�~�����h\x�W�f��O�盁G{b�]���i {����~.q}<�	���`�� �)���(�c�,��e�طɍq�޳n���6�����������HZڠ�I��Ƃ�b�_��c�hd��N��q�f�M����t9���཮�l�rF�$E���`sQ��<#��:��嶺&$��pwe���bcz4��fZ�2��F�Y�
�����ϵ��r願:W ���9�<:�N�;|Nzy����{�_�юw�]�a��Wv�}�0}�,�G���pm�Y
B%F>�YV��X��-�����<0���y��m�-O�1s+����4��� bD�7߇�V�I�_��r}�L�!��t ��	B�������)�������L�B�@(�l߁����%����3]��t,������@Mi�ީ z܏�&����u�ڙ���:�E�éy�{߄�(����MN��c��.����R�m�Z�%���T�?g�Ή��C�N2̼��U�8z>�>>I�o�C�x&��;�jh���ͳ>y�-�#�tT'F�y~�Z�
KX��o�̚��X�pߘ^{1=��U��Vs���30{'�:��s�e׿�]�����C���Mc��j/	KǊ�Oe'4����<K����i( Y�y�S�w��EaGW�Mˍ<>�\�R�S*X��,�W�_�--�E�M'�6Gn��Ӆn�:��)�k����G�B����)%Mp��}��9}�"֏hih����Dk	@�C��������;��"���N(B����69�Ĳ����{D����k�Z�Y�������/�CԪ6���a~>�Y����� �r=�e�i��? 4�u�W'ᶤ�d����nS�������װ�X�
�ؖګ�H�"���Խ1��Uq��?~z�	4(8h�מ�j��-8��c�Jw��4z����J�Paz�G�%�*I4�j���/� ���K#�N���a D�J޲oX7* Ɉ�;R�����p^a�b�x%U�7c���pc7wR�;a]��tk�B}�!1Iw,����I���d�'�Î��rmHݵ⅜��r*~; w�ӡ5�G���t�Y����&��~��:����1(i:K�9�/	�&�z��C�_���	�c^b;�+�%;��/���C�z���s�;�]Xy�3��%݃X��@@���l����5� �h#i�hE���QJ���/P�B�}yڴ�ly�������~}���FP���س�@��Ϡ"�c^���j|X�j\f߀���p����lW@+=�.���ٷHtS��)՝��g˪���x�?6��]8�Gm�J�X����Օ��}�/9!,ΧX�9=ی��K�%q�C�dy^&=��%s;^Ȟ-��~ /�H�T�T�AB�
#�6��Z��8	/�M�Po��b0&��0�gG�]�~��q?�b�O')=���6�F�e#Ϣ����m�R�>� N��	Hd��~�L-ڗ����y�RN�V��%wH�-.`;��F���K���:��1�����T�&���"����6�ܣ���8�T%g����v��iC����m�	��^gÄ�6�I1�V�v]@�"U���Z��ע�uH�W7hT�?�:�4�.��b�Ä	�߿~y6$WP�$S+�
_9;���]&i�S����6����&��;-��&�'��X>l��^/�"&V�޽�q���M�e��,9sWRWt�Ti^> ��:��#�\.�ff���e��M[�Z�nqP\����:t{Mr�;#F��qQ���bL1�B��<��D:�m��w�?]�u�Y�N)�jT���"�gd�W7J��j�[�6x[h�]|�#���-/AeV��gC��a]��ř]kP�����O�KP�\z1�n�5j)=8e�c���9,����k9���H���
�N��+���^9'��{rm4��].�wVY�;���$Lt=�=�T��[�G�ǅڱ��R�uG��/�A�,����(���F?�U���\1�F
dd���0��L��Q+E>�͍��J�yb�n߲�k�xmp��DRw�1�[1�-�����%l��iL�T�)p�)�J,ˊ��$u],[�9@���=o���J�����|ťu7�m�+"tf�8�	�����z휙i-r�LG671�����Z��x5���?���FL�`o��>C�%�}mp��~�Cr�J�;���HBi�֙����/U!�Ǌ�{iB�+H�Gˉ(��=�Uh�G�+�+�P_�|_�%j��|~��BsX�B��R��{
_oT���d�����#��2��Xe������T��Δ7k�<~��b�b��1^���nQӀ�0VHĸ���Ñ��g ��f��QIY�?T`9q価�V��󽧡��٣�5YY7�g�`�k����A��=��2Կ��X�c�yɑJk��柣��{��I�3��Y�����Q�|�-�)q���|�b){b07�U����l�7�*��2�JQ��r0[5�r5CE^�g�6����8�������z�����{Y%����t��2WeS�$Q���F�*k�IX�����P���`]C�d����fG��_0���[�c�\~P4��{��w�Ä^~��,���3tǨˠ�i�@`.I��q\}�o��F{���w�M�:��hX찍g�Ejv5;g��=��U��#� I�PJgB�!Q���>Y��=K�3E�����F�<�S$£��\�!&����^��l�R,sR� �ط��e��e�ɶ����d��ƝnF�Շ�K�����1��$��!���փ��^V���YV�9�b ;��$N��A�C�]\z&��A�:�Pu�^N��dsp��(<җTS�{^�� �>U��+z�CGC�����z��߷+�o9HBY�u��:�����^��zg������ �4�['�28�E�2��y�K��gǻ�d�#��N��@�_X�����Eֻ�/P\(3�~~�A9A{g-7sBȭ�j���t����>2���D�AG�ˌ[�qB-H�������2�,O��IZi��ޏY�P���M;e��\����04pyTs!l	K "~�C�|ũ�멒\:�_�R�6��k�ڇ��qt�j���~�ɱ�~��TM�t�?��g�e|�j�$���:	S�Z���-�ۤ� �B�Q74.hǜH$��2H(PE�����f������'o;�F#N��t�0��̒�`��~�����;��X[�H���]�Y:��Qĭ}.zoͅ��� �WuH��E��>%{5�X^ܓK�kL���=SNY�U��<��*����1y�.����l:�y���N�����^���dB�n�_�<�ry��;/>5�4�dj�̖�7&�y ��|lu����(�$�zd�X�p�� �=:�Yiͤq8�t9m��,%4~,^��	��Yn����Oq���/_'��H�"�t>"<~[���/�̃fHsu����9y�\ŏA:�  ���}���@uUy2<�V��D��7h/zv��Ta�x�(�W양��U��21/���a�{7�D���.N������
r�f��x��1wetꗛ�2���8&|vI�:�a�Fبf��a���N�5rp�>I� 7wd;+�hC����kJ�
����g��g�y�𥴍��}2�X�kHV�rhXA�9�	?^c��I�НZb��X��2�R��滁_��3m�����X���ƃ]��x�먽�W����ھ��#0� ��b���D�'�o�;n���iRa��=�ܖ-V�C��� �T��9+�ޝ�˓SP���n�W'�cG�D��H?�+<���LQge��a)����$/)W�fd��\2Ոt�B*��G����d�Ga�D$�Rc�t�L�?F�Nvr��m����P��I;d�MPl!:��2:���z��������a\��I`�,��V\#���$R�#�H�w�H}f��5~��1��^�2�P�)�+Y���;�& nhu�h��3Nu�c�>X%�c1���@��3Y"��I���É\�d��E�g�����\�Ls���ɲ����d
�ժ�s�J��싅A,����'8^qP,��Q�~��"MB�K��Z����tϹ��dj��i�Ss�S1H���%������zώ��?�xn��Q��,VN�R3�l����m�.��D�z�.w�����~õ��B�  ˸�$���d�@s*L,G����9��"�K�����ic���Ī.+�)|']�=�!Pń*5v(���zg s�Ӳ(d[���@&��ӳ[�ԒƢ��\1�_��+� �Fc*<���"l8	��Xz���"�l�� ,�ss�byʚ&OC��b�OO㟄�1w8x�F�T*��e.�j��%WoLt�a���:���c�~5#v�X����!�/A��Tl�!��:������VG0�g��x	��Vi�v�����7~*�8����zj����t�6�TTܲ�c�������Rz����i�G|��S��T�&�2�8}��]�27�z�}s"�V��P���r~XJ��%�
'H@��\ �+��0��:����3O$��l�{Q�>,�|::�=ը(p���%#����]�&��yM��ג��X�|c-������������@�<>Z"C�"��C!ـk�l�H}�ʓ R*2nx<��6��S=f7��(���?�yN�q*��,�'��o�}J5"���Ä�ʛ�ؼ�g� �GM�B}�X�z�F'4�&zh�<��u���f��dw$gʾ�\�����Npv.S?=�0I�L��-շ����۷���v��-��]����^9԰ŏǷ�?�yi��s*4�d{CZ�����y�&>���~GC���|*U�_����ݖ����Y�v��7��G��C9��)�[�F@oPu:�az�tU����GΤvl3����.��mH�@/��I��r�����
f7�DE��4_��`�)�NFs\���	���э��&o����lj�w�6*���g*��c�q8ٶ��#W��%Ӛ�H_�f.��V�爵Ik�AG������^Z�q�;�I�Z�A@��}�@�^3)��
�	�7�N��2K������Ӄ�Qa�-E�b�	�Oޱ��g�{寔�V?���G��u^��ŝ*���oh������	���:����o�z�0��*����t���l�}<q�-������ſ+�/���m���-��bo^m�\��G	`���)�"���<�ň�pl�|_�ĭ��O�W���ǦTT�w�8 � 5LƵ�ab��dicr����:Y�������b������V`��XUTC��rG��A��)��������{�����6��^d޹*8�ѐ�ǁ<�����xd��U�r&7*�u[��/ө�O6�<j�t�� p̰e��5
��@��1p�?��Sb��~�;������Fn����Q��p��G���G��D]&E�����x�R���+ö�CG��1ui[#��GI�y.?�)҆!�M�����"��,�7��fV/��u��b$�B�� � oT�[G�0u���01������*b�RO����PܧNġ�%==Tg��W�����խ9���[��Ȣ78
D2d��c����Op�-
ed�V�={oz�&3�٠ /�(L����+21u>�Y7�R�|X�Lro�L���3�������?MÛ��ኦ�I>��B���MAڔ��-�P��U�DI��%�ԛ$�m���ߐk5���3^e�u��F�2qq!zCsIQ�ޱ�p0Aw�Pc�z}&e _俫*u��"��y��J��\���iW>[��\O%��}z�����|��	J�\����ZC"�E��d�U�l�b��C�`�����^��jc�&n��F4�G�S���d��D^vů)�TpZ��-�p_p��t���;��(��QhI���X$���x����رu%���C�Z�� ��c��I�(����L�2|T�V�Ǝ�[<�@N����<<�ժ�e4���x���0��,��dEl�HtYJT����,�8F�׼���������g>v�{O�h�o(�q�+֌�%Y��|���2<�xbw3E{ׯ���T�}��_�Tnx�0���i{ջ�{L:~պ�t��<}��w�X�tfL��#�����P��8G}C�y6.����e{��i�e`�P8E�f�Zw�$�b쬰\� �/�|���~-u��r�^J��I!V���|b$Z${�1� ܤ�����d_��6�<�c�%ԾΞ?�1ч���1��6�3+nk����T�7^�ā��}�4aMh��J��${/��2�㕖-�̪,���`ƿ��&���D,�|lz�59�Ā2�qÖp�i$@�ITV���&<>?��EAn�]ߙ�Ƿ����3��#¨�`�SS���d��T��Umi�1�&1P7�f�C�ά'��Q�W
ԍtx��� ��c)�G�뛗dzRᔊfD��;��Ҝ@Ll�Ԧ�\�C�~�G�RO������s��ge��|]������faJ��f;��,���,~ �8��X�G��ƳK���ܪ��K���v�r��)y�G͖^���m�����0���p��UO���Q�s<����<�\.nUk)�G&8DfgƎ� Q�r);v�sX�y5���iMk��qh�P��Q̯s�b��{FN�!:���B������ &5��ʺ��Ar��O�������0�a����w��;jFDr����V��2L��)���3c?�A�=�A �@m���B��{-ZǕ�]�!�<�Ò%-Z�ЯKz7"���D�WSp�p᭹�ӊ�;�FP��+�o��y3��l	e�fe���#�fӟ �8���U�g�P����@�ɻ��V������t�S��������@Y�C��5�ٲ����_2H���"���o��������[�m�Dq�&�`!����Y�}i�������.�����a;8��S��|�q��>�K!��o_#߶�+�"�Fx��خ�,�f���16�bޒ��Emc�{&�hz�#�(Zb��a#�j_�����	���(�r�q��M5%�qY�#�ěR��$�����c ��]ߺ?�W��I5��W<�%�ȳѷ]��f���C��@�6���X@>�B-^��ȴ��T){ɬ�h�^�@yK��ˡ����������9S ���n�t���KH`,���=�c8GW��buaD�W�$6)�� Š87*w�<��X�$�dZ[��V��iE�G(�oNK�}P;�C,�KA�p�{_�����Q�����݄Ut��/QP�}��*�N�ڀ甊T�JS�����x�Ca����~��d�I-E��V�)P�����!҅ɺ��vY�I�G\�!
�����p����T���B�E3J+U�7YS}�4���|3Z$�_�B�c�Gb�"<�
�Z�aA�zmħ�i>�}+��A)�W��Օ�:e�����ʇ�����yoK>�u��?�WUS��%�H��u��?��M��C[u<�lq9@z��Qܛ�`X�������K�{V%7�����]�˖ۤ��K�j����)Lj����om�*��{�$���Ԩ[V�{"��xm�K^� �؆D:�G�usk�-.���gVVyEV��~F�x�S)�/�gt�9ll�P��#۵�Q���.4l}�L,#1����Ω�F�wbҺ���JM6��v�I���}��q�[G���q.��b�{t4:��7,�p���ة�#�Ƙp@�D[z���+��n�j @�8�������O�N����}���E��}���T�ͽ�1Ĺ�`�}��ZQ" 1W�\~I�D�%���Op���堮g��T��{���>
:"M��_p��L���m��Ov?8��`<�(�H���~�0�zw.�N/�
6����f�R�U��6�{ZA��w�4�_AX�>?|w0�>�5�-��y*����7S��9k&�@��|�>{
!�o���:i�^U���@� @���'����6{c~���Ü��(�_��{��z��/�m;�3��L�^�X���������;f8�S��=];,�W�
̔0▥�V������>Y~���b (&�����2��Cu]F��֧�>-O�䔥v�6͏����a]�'tᱣ~7�AB�gRs�����;r��M{eP����*+�j��;i�� ���)yAZ��9�縯5�x_��l�1/���)�4qp0f\X�1m?mÕ)Na'�}�3r�r�}�l�I*.�P�ϐ�S�é����TvV��q� ��l��H�M��-\ѱ����L�<rc�mUh]N4U��Ô �����N�&F4�0�Bc��8h��>Z�k�����=2���^_y��w�kJ�⚥�9���o���*~�j��G����שx�q��Cƫ0�1Ù��*{h�8�3=cKU`5��rX?ݐ+�t��bg�l���[�t�� ��=�d}�.!�dg�~�-k�ԉ?���}|�s�����O365�6]��J�*Ч���WY��)���.�h��/J�)�)r�V/Üt��0�w.zCj�ߺ�D��Nx�a='-�S`�ӛHi�oт%9�eE!@��[#*�s�d�J8�bW�p6_rd���O�i�Q��?bW���;�D�s������3�>���z Yx�7�E�>K'�г��4���b��-�ʼj��%`�����}�l5r�f����?t-}�Eé��/Y�ĪV4��6@}���d$fU���i
�����Z%wy��4�W�l�z/O�W��gx��d�]x7>C{�"���z?����f�5����%o�(!� �!��C*��V?���y����vS�B3���p�eC�u*������B�0��ܒm��,�f@���G;s��Ns�s8���x��ܨT�§�s�w�W�n>�a��:�lAk �,�й��*���z�i�\�e �A�O�	ᴅ�1)�VGc��@I5M�`uf�I[�h���q�6��X�vVf��i����{^>(m��%.�K�:����W�}�"��a�7W�;OzWȶߝZ�<H�˩9�J�wU4m'SvG�^Zoʁ��ŭ����1�eK��WS�i���C[���^�L�L!�Ih
�B�Ȓ�e�!Av]Y�~�t�F{:@45�?3U/�Z���h?�J/����+/j�CiO`z	�K�b�(Ǐ3���f�(E����Ļ�� �xC]�-�-uK}�#�VV�ӫ�o*�n-R$W��f����%�@����Z�:\��SF��1�����R��Sc��W�]�1��,���:�;�p%��W���0����G��xARg��)<����mj���+�2��)�`g��I�ôy�WU�z�~z�Ϋ�~���M�Ԝ�@'���
S�	�F���� �M��O�( ��\7)� �^��d�\�g�+Ku���R��`
�B ��7Ǳ���C���E$�s)�/ݼ��Ѡ�S	g$�9��:wR�w��:��5�.��$9\.�h6a�`�>E��@T5�/���fB�=j�"�A^#��ȱG+>��"W��H����_�<OG�?N���ò�*k�Ά���H�g0����L��k�"�V�h�؅�0��Ws��½�zx�S*o�4H���廔��@�P�te��%�ro�׎棘��D�~�'���n�x��_�Of��<w1��H�G����Q�w�ZaH��.���X���p��!��u�=��d2�� 7=����\\���G]�Z��US�Pj���~j���ec�̆<tpn������(*�^Qf]]V�_�*����"�RDw�f��F�r��Қ�����kq�|��@�&���	]{��FLY���ZU�[(�f����!��R�H���8���n2���ZMmԨ��۩�ꃮ�p�
,Id�l=����B$���$CsV����Zē�j�+Pʹ&�Jmȝ1�V��L�LO53x_͟W~��b������!���H�XU�����)K�1�J��>
.�,���A���� '�].�A�����o/�!qB���uX�M��7�\������	DB�V9���V[���aL�/�Úm����ϒ,s~�$n����jlg
Ņ��7���?��]�h�V��p�Dh@�P��r�5OROY�Է��7Z�鎚,�J!�誳�#>3��
iƓfr7;-#�,��w���$6&ȣ��~ЁK {EG�"�c9X]��k�;#��y�	��I߱%v/۲��\�����i�J��s�;$���������E����!�GO��
Y5�t{��'t�U\��)�*��J������&;"j���˃[L,�U�R���)�x��X)��R�+�<�LL�f7���u��ϡJ�K8�TmL�-=��C�p�v�#^��ܙ�Ζ.΃��Ж�ej��(�x�O]O��+k'�[7�#d���d'�gdLuI))���T#ʜ-a�xMJ�v��6K�g�NJLv�������kҭ���D%9�ũT,`f��k,�F�����DFQx�
ύp��6з�z��9��>��#WΣH8��֬P�O�=njQ<Bmt�F�� �+�[��sg#+S�j��%t��\��G���-݋�$z��j��E$J��������)�E��F��%�������8{�t��p;-����@�t�Q�I��Pᮃ	�N�x
�$͵�h���_�&����wW{g�'-]�2�Ҋ�h�������l�W+kFk�uώ�J�TP�|��}��еF��E�\�{�M��[F;��9ꮌ���U�T!��jOy��^>sU�R=�I��9!�p�X�������B�x��]܂���5�P�.�l��V!�k�89�i��W�"�q�P1L����5I��2��˳���ؾ<�v�9?a��P�K��|��>�a>[�=��1	����v��2Z�{��/�#�	<g���{~�v�ʫJ1�(�-��>Zs��Iܧ(��t}D�p2:L���G>����^��5��ü��H�J�<�3���g6	�K��~��`q4�G��fր�nU�˱am�&��wEr�Q�Nvˁ�_�j�5=�2U6��М��h.n�B�T�M~�kVKt�()��P�S�(I���뉉�]Qju�ϛ�$������e��(�al}6S:��D�9�7�O�%��f��]�.��S�V�z������Bʁ���%��ؘqH9Kv���B^����Q}<'�L�=HM�VN��x��[� qoXó�%k��vm�����l�Y����b����m�o�iwr_d����RF�xo_��s�5fr	ڂ����T$����P9�77V�ª#V\��~<�c����Tyִlh����h����{�G�s�ҫ?^UJ����S1�]{Y{;F�x���'
�%Xb��\�\s�o*�9]���Tfҫ��g?��!9?&������ο㔎M?��y4��g��<h��Էa�	QfT��z�Q����[��	ܱ���JY>�;�V������iq�Z*i��ձׂ����S2㜔��/y��4��gpz>>�O<ؒ�\���C��[d+)b�{��0���f<�V�o����%M֚�N�
_Ö��+Q���Bb��h�,�X�~���3g��[ĵ�)��s�p#�#XC�:�I+c:���l1����l�9��&`�i��	h�Qh��� O�eI2b���������-�^ޢ�&�B��<�����KƮkk��^��j�$�{K0�!�T`�e�'4�;(�D��=�t��y;�K1t��������H�Wl�c>S�]�U�ū�"x2���h��I�E�8���ɕ��33�F��ź����x�a�����w�F
���9�>�?�-��,���u�v)���e~����ϲ2E=U��A�C�['t"��7~&��ǘ`�t�m��?I��F9�!���<5K������\��鸽6�ܣ�j�T|��_�7���6H?׆%�e�>�V��{�ԩ��S�D����i���瞧�R1�R��O�\�� ��u���V��
�K��4i $�K����m�꯯�1 ��o;�����1�.�B�{�-ŞORDWw?����t�	�c��b�d蝝0_d����#��+�U�l� �"Ϸ���Dɶ;�¡�KD��~YX*�Pٝ?8�D�}�q�{c��?J�p��'d�M$�S�~���͝��k~W���)��E��n��ˣ�#�䑺!:�%R7k�h�Ex����#�U6��Q��-K]3{l�W��kK�����󄏣��X4|Nu��e���|!��t(�H�\P����ӬO V���쐏mz+&���<�I�@Qd������h�Ƅ/�]��ڃ��t뼂���&����l��@����W͍���������8�G��JTI�Ժv�҂����{~��4�D�_.�:n�[&Y�!'�&�*�ҍ�#t���,: �OZW���\�c����)����g�?�8��:���f���s�f�[%�n��3=�L������uә-�n�ة���O��`k�(�J����P�At�,VQ�'ەI-^@����[	�ЗKv�FZ�!Gp�e��Z����n6C�	�݇��ù�l�~�:��/�a?#��]�0�O�^�����Fb�шU�h��v�$�����s�f��/�hj#]����������S�A%/��?ٙ#�V��^�0��̕�o�������D�ss�A��!s�@�� �Z��;�P�j�_�*R�w�bT܏DD�����۱���'��1����"�h$���ЎM*BB����Nc��d�=����~eZ(BD5�F��Z�y����d�5�p���Z�N@�����&ڴ.V��E�YpTѼ���l�	�f�Y6J���i�u���s�E1����F?�����	�wP�����K�+�:E$�/�;E@Vs�u�,P�i�����^��f�7��7#-��DϤ��V@h���Qd����g/�?���h�|�r� �f�tى��J�L�@��y
����?Y�Dq��W�#���&�"��e糲C��ժ��Z5:I2��I���(;8�ӈ�l���:3�Sdb�S�R�vo���޻$L̛��ۤ�۔A�R_�1	"�s�0P�"���Z�)).�`�5�M��(��c��oHn!C8:$�-��S	l�f2�!�t <�d��v&�Cy!T���'O�
��<Ǩ��v8�3���$է������x��ᦤO����V�����&�Y����º/��$�P��!{�2x_����nŬZm���m1 �kM���1��k���!�!���-����V�U�;`��o�t�k�=6�
x�)���b�{p�~�o�Jo���A��h��8a�@��h./��Ϙv���c\^]6=ħ�{,�6�/�"��ұ��~���\�N�)�]�}9F'�]-��+8���*"���
y=*?ڀ(�)h^�����A'oҲ���h a�!�]6�^��D�� �=ː��3��Cm;a��1��E�@�4_�Qꆟ�����Q���TI�0�v76���^MFm� �__,���C��"q�mJ�N2'��S��#��K$]�B���P�u&4F<����F��_��,hCn�
y�Ga�n���4k�c�\%I|v'�9�)$����[�[Le���qC�\�`�b��s_ڮ�jE����h$�*�T���KO�O��L��y�)%n�y�<���PL?�`�o�]	�\�Ԕ��ോ�xض8T�A������
�����56�z����&(Ww9 zbf�$Cn���bY|����p���}��̘��>l)��6>��r�4P-�K�z|'%�Y�`��5uR|-H��حI:��>T�)�%�Q8,�=L�����Wd�VC�WRVkM+PQ˴�P����,"���x"�MN�9� ��q�9c&Ǟg��]N�\O�tW�;T�W��þ´�����)�cz죺�-�tM�C��6 hu��\/�BΘ�F'��0A:Dv��6��D|�X�yr�G#��J��O� �l����(�J��cD��q��� �k`пP�g�d���"E��K�ǣ�O�K�+�X�5��K`E�w�%N4ORtE
b��U�A��]㠌8�Հ�b�1����s3�az� 7�ƭ�Y+k��"谏�������%�T�����2�	]�g�j�u�-�2g�D��wsi�W�fH�F%?8܎"&7��'�R�ݎ����	df.^ȽP .n�:u�>��
2maC����tZW��Y6�<]�Jw�R�/q-6"1��W��7D�q&��|Q�s[���K ���}�'d]$�t�/���z�Z���p�7�#h!��������[s��e�������m#b�1ƃN��5�h�����Ԃ��ޞ��VB�S�������*�.�
���M�[p*��ˀE#�⤯��#㜨D��:�]�`q��3�'�[ٙ�M`�P�J8�83j�g�&�B�y���7�?��bv%�Ur�=d����;�0EX0� ��_ǱѠ���ٕ^� %Fo�v��?���4�w��-5�{Mw�!���I��L���fa���
&v�(ZdSa6�j�]�B"lB ��é���[�Ӊ���gz���!k�*��8��(�d*�Б�����fƍ�������Gwu�pHd��&$� �aЖ-������
�U�n7A��Z@������s[W�Fe;M��8sI�~�a�J�"u���{\�l�\T�)Շ���[H�}��:��@w��Bzvx`�ca�4��75a +-a�o!�t�A	�V�����C��Lfs��%/��*�j���NFS���}���X�pl�n�J�57d�2�nz[��ɂ� >�q��9`��r��]I���/�ڙt��(h0�^��68x�i+}�y��^6�h��� �,�m_��y�:�Y�t3Nr�R�%!�Nx�t�D��9�g]7��� P�+[H��x9v��0R/%�l��M��L���-k��JNCB�S��M逅��?��Ofz�r.�Ȓ��^��� p�I:�u-\�Wmc��RQ%�\�;%����y::>��mo�����6b�,"�uD�7�X�F$;|V�vm�*a4#`G�2�7|_�x���U��ڔ,��A�N)���-�]�6e�8�ϲi��YgP���NI]����q�M��Ǧ!�k�B�v��5��R�?ѐg��8׫Y�y3���O�)B����-�R���|��!�W�T���I�X�@�*��Wnڟ&�^��f�-s
��E�^.9���=�b 
2��r�y�9,��j%^��Ψ�=*P��B��s�cr¥[�HdQ��5�ZlZuQ���&�{s��Z���,A�X��q��l�_]���Qr�K�P)Hk��ʽ�_�(���,�@O]�T@���xڎ���E��KB3%�;��w��g5����jՍ�}~J�~`T��.\�G�3� ���,旌r��^6ߗ��tCMI�VD�}#��<6�*bx}��?��.5��{V1$L~=�)�.���Z�r�o;�����ϗF]p�)�� ��c��m�|Ĩ��͜	]�x����z֩2�����:�@Oc���=%�.w�������O<Q�g�:N~��<�Єo��?���:�������y�0��(r�����������_,���T�;�������
%s�*BV�����f�]��?�u����Yΰڳ�Q+*��Q�¢�4q	��EE����İ-� _�y")=���1;9�7��o���o��w+A�i�E�7��;nD?��k�aO�d�Q�j�Ҿ�>F���l/y�X���%�cL�k!X��m�̟�7G�|�����S
/W�����j�����.�n���T�O�D�R�֍����)*��t� տ�/$�ú�����0K�D&��>YC��*�������\U�F*���:�f޲A��:"�ތ�Lt� _�E��Ώ�`7��?K_�z��p��b-=J,N*��!L���5��U�y�#������k�;�L��8���O��-D�I`�gFc��X'�8�a��}�s��:�S%����JB��V��d��GaeՐgsPs�y�h����a�
��S9?��b�,���⼦�i�0��V���B�pEDޏ��M�p�?��'~����1<�Y�||G�+�Ȏ��V���џ%��&"�3�e�b���4�"���U!�Y��`���*o��d�lSI��a���C�pj����' n�Ϟ!�Ec���y���k��4��~1+�*�c�(�n/�<6��pʐG���z��ax/�JȚGD�֗Tcl��T���s0<��
��%�5�2p�:����b�S����`��ԇ;t���3�;�q.��3D����@�"��Mu���@e~���.X�D���Y���C|}�2�SC�z�X ����ʺ�03��R��S�5����eW̪�N��4� �鉀��<��D�Q�h��O�ݕ��BD���z�}3ݪ�:+��H�i�W�N�������w���K�rK�}I��P�G��Ϙ9XD�-��?�9�p�iv��g�́kz�a$�F�􌌻�JP���!��^g�_*�I��H7�=�C����P�ң����j�9$t�Er�:9a�(�k�������4F��X�7���l�Q�7|��Yo�xbP8�ۆ�v��^w��Q�����#�^�k{�4��Ibs�
�9I������.̬��J�>i�V�9+)��Ӥ�^��p�]��AG�+��i�e�w�/��-PNM���Nm�R��� &;�i�B�U��5-��!���g��b�{|�Y�?܏�u���@���`r,���RT!��'A�F�[���W��O���~64�*��4�D�iX�T��  �h���y���+��.�\ۦ�@�I(�귏�f��-J��1�.6&�����G�3��*�o��8�F��&��I�W��.*`��LB�G�G樉Dzy�J!����)$#ρ\PO`ˑn> _�{��O-"�%�Gt%n4�vͲ����<�Z��lR	K�[��=X]D@�6=`��&Q�\�c6�z�ː{��b]t��41�%�Ũ�1�A�~�	�5�Ԭ.�L25��7�K�~]B�aY��U@u����ε�&խp��-,�O��[h��XG A�sd���2�lO���xG�J+(�(?EP�5�S��C���7G��Q��ˇ�z+�|�A�`n�,&=��(�J�"cB[�}�. �
�	���>4d��c��A���x��N'��9�6g��{<�E�*�g@��ÿ�������uT4�J�]�wj�`� a8C��G����ުF2˘��o�p��݈w�u���P�#I~ 1�^���1�-��3��r�nk�_����:g�z���An#a���<�8PIzmH(�J�-�L� 9�ɢ{�ÒM�*�$ to�l��h����j�����]��a<��)Ë�7��.Cj�X�]�-gm*�I@�0����ϴD��
�/�Y�����|��l;Y҄�E�h�����MN���&3�'���y�!݊�itT�� ؘ�Ō��%���a3�0b��w����L��B��v_Pɴ�Q��G��@k�0�~�G���
��v�+M�8h
��޻�Ӆ�vU�U���`�Ru�3F�Td�4EsV����i��/Xy=:�q������,�D�����i�*#��N��{����$�:�,}e=c�p��r��w� �֧E���-Fy�ip���?�C�����X�Z�0���� ����.�=bR�XTϽ�,M픷�E�׭4=��+_*�x�%�c:@����w�"�}��|�tY+bpx�-�g�\����h�՞��
���0<�_Մ�V��of$z��V:��`��t���:�H�f;�V���t R�1mI.��u�	��x��h%�����]GR�q���RJ���H�?�j(�n����[#�
w1�Å����s��\e�J;������6���t���"�>�����ul}�xv�c�0��A��7�W�RD�m�#],)S��Z�
[��3��W��u�uc�3@Bt�X�Z�z��	!x��Sʗ�zYc�֦h/��ҕ�}��j8�H|��+r�O�G�X�Ѕ@.�o��f_�?�d��,l�pSb(���$((JsK�_�S���CM�ފS��oʯ��a���,�jq܏����4@��y��,jt�}[��j��(`���*/�3:��T��J������4�;$����z�$������u|����2^
S#}X���`�/ �����5���G­_1R'����I�N�(��.:◎��9);0\��ѱG����M�aK]91yq����4���4����J��8��u�7L?���SR6��Co{�Nv
��5�y%��Z������,�Za� eZ�,�8b�}"�λvC5W��Ὺ*�ڶ��j�Ҋ`�u�s|1���i�`xtm���#\����p�稧��ϯX�.��`�׵��2�c���o&d����E��Rl~s�F�F�O؇p�4.JUo�� Jn��%.�sPkDQ�����-�׬��C�v�%G�d����s����~�SBzV������(x]:p-@���S5�\OyU�ey;�|D%ڼFnDZϔ9m���B��o�Po��'�"sSv��'�Wi[��� 0pB���e�5>�[lq�d8��g�ǖa]���b� �Ίg���W	����K�SAB��b|�]����I�Ho=c��xH�)����\�}����,_1�8�%c��Q�I��+��2�����BF�ӖW,�uG<��7�ݮ���9PF$��Q�Y�-aI�D:�K��BͰ0��Ԝd�>j�[s)�N�̯q�@}�5	X[�Z g�"!��A��L~� ��Y���I=Jc8-pǎ�0|V@N�����e����Ґ	�|]1�^ل�\z�U)�:řuD�9 �4I���8D��g⟙vv���R S�J��*��Б�@$�գ����XMKn�w4'�TK�c��tav�U���-2U��ow�e�1�&�uj�:_o	]b!��\)  m}2�1�	�/�$ty���u�M�N�go���%�������J���ۮ������/�W��l���]8u�|�x����@�F! ��P?uA}-j�ԏ�bHe3K)����%V`�}Ϛ���N?�į(�*��6���|��)����a����x6s2B�,P�;pz�w��Q�g�"�[��R��q�+٬����3B�	ۑޠ���;"<��v*��u�KA�It=�7�	%z���%?i��8�x$#c:W*z�/fm�Q�ʵ얭�&�?yut_%�uHR]XG�Cj	���	
SД8�&ɋ�XJ�7o�ya�3����1�y���l�`*�a�i	[ ���#�z/�x�qVK������K�
�����f�Mca�,]ıj���폸�0z�sAo�S��G�f���Zޮ�o�
�m�M��,� ��N��0JeW�%r�v�/�'%s���ذe��i�ot�o���N	ݡ�+$� *�H�L�@�ܿ��ЧG��X� ��2�-�S��*�1H=��(C5�4L<S�φ�O| ��ɗ�{�yg���<�5���������,㎌��D�q`�ߓKU�9ó�!���b�#R3���E��"�h��B{	�gK8p�4h3��߻���p��������I�g�$���=����t;��f�mGK�Q�7��TH[�̾�l(�"��j���3Y�8��
���|bq@x��_v_�Bd�n_�G�{8q%2ȵ)͚��+�]޿�?�\4��?h�:� f,�W�>�gwo��<A����Bn����/�D��\d��̣6�ڌ�����R�R{��v���s[���@�X%�B��b���a�$�8"��edĥJD�x#�����1���|u�� ��5�,]�QS w��S:�������f����j|�IT�e&i`��?S���nQ��?`�jV-8Nb8NX���ER2�+���)�=;��ߓ�t���.�.����Ur_�/S�"g���@����(l��:6�k�)IZ2�<�ڳ�PYx��5X����m#G&�Ko<w6�a��W�)��s��?G�i�8�V��V��/����!#��}Ds���#Y��� �j��I�����[MIt���W�u�+��)��bz��F�\�R��|�<������Ly��L��e�+�Io�{4x0�p;��_�8�FGՂ>"���z�ojf3�ck�o�����8�C'x���#��W���H��.���0��+K<��"�Y���%ڍ�(��z^S�ZzB���TK�|�x�#���&?��R�q����Xn�W	�{���C�?y�5Jv�԰��^
�X��=Ӟ�)y�4J�uW�P�;#��~쀰r�K��2Z~>^eڠ����ޑ�?���i+0�m�m�WT�r�|�%���,����1��+��f�Io6!�C-ʗz�(v��&mo���Db����a��{9�6���!�����60�8N�]��R���
GvfU z+��"�]�"����ϯZѿ`G(9t?�`0}㢺�7��~WQ�ט�0��9�a4ޑ�|��w]J���U�9�s�T=J�?�ʲ�9z�����9�g�)���/�͂7�j,Q\�j7��!��R,M�\�z\�+���׭i��@�<���B�'�eF?>�
���ȴ�[q{R$��2��	������6�%-�`�A	$�w �`(��!T�m�=�����f��lP������s��P�&�l�_�\�z�5n�`�&���e	S�A^8�YJsJ_�8z�`֔Px�;�/7�֑t����,�QC*~X[Y�g�k�' [�?)]*>P�^F���C��ӕ�/9�� �F�#��a�޵�!79��Y �x��&���,e޴M���E���x��(�d�ǀ�6\��\m��I�k��3���A��'7�Ǝ��e�d���ө��BZ��73f��t��\8-�������Y'om��r�,ZF�/iRg�)�e�E��q	)n������@q��{�f\_��#5��x���`��Z��B������
�,/���uGN�6�)97�>��]�m����^",����*|t0��u��e���$�&�f��g�J��,k!�@O�5@�#��S�߷W��T�>�Qd�R�$�#󓽼 �H&�c־v H�����а�.��0�❾<C�:������~$9%�#�_��mZ��tf|��r��ZI+X�&��ġ�N����9��/K"��gW����u���d-�q���Mϊ;�W������ٲL`�uo�d��^Es���y�����g�� ������ �]zA:A@��ʄ�·��) -i�v  M`�T��L��9:�r�(�Qjo�.h|I�}3��(�]��WZ�}(t�������ڵ[�v�!gh�t���t�����̝���}}L#��Z�|8���L��I�%��:ہ��䝔�'Ӣ��ki7��73�*Iu&�@˘k�p�䗂D���K=:֭M��Ye��1���Wt��B"s}K�]��_=�/}_��J�d��Ͻ��j�������<��4z�D�%3o��ډ��5�$�;�JF"xW��Q�k��
A��(�S�ɛAå�˗�ӹq�c������r����V�he��2ŷvr�.KH?W� ,����%9�P�_�)�H�n�ϸ�2�-EV�B�!��?� ���>E`8&�F��O���(����QK���=œ�2?�ec��9L$�W�Jn���J$D��3?z��ĉƍ�3
H��z�|ҒB>Q_o?`X�p�ԯc��WC���3Y=r�F#.c0|tj\����O�tڻ���H�'P<3�Jm�u��+r��j��>��zr�E���xY�hs�H$�k���lO���ѡ�0��nF��i	ui�>?NH�wz�	���8�li�o�:��F�ʚ���N�h�#��+���Z��Q	a_�؉�/�[����ߵB��P�->��(�-~,~#V��WĦQ��rç�e�ӄj�
-�t����C�_/�<�.V��)���H$�|,��!����Q2�3s�B8�{��@p���m�c��{��9M)��vy���܀�r{+�L^_��8Y\�$��v��*(Y�ʑ]1i�:+v:�.�^_�G��l)y͝.)����*��br���p�R���7�t��&�L��w�#�$�@�w�/xPX�/쟟!Yf`���J�lznY��UJ��{�|��$���=L38D�����b����Y�g<��&��+�Aw�pY�~�-��g��z��*��6�A���nxeR1J Λ�\�F~��8^^}qn��N#�)�����v{WG���K�[�7��|e]���$B��|�7�� ��,&n��mP������?��i	�yq��E�/�q��@SR����g�V�ݙ��Ge�f��-�U�bsҦRhˠ��{�����֡I�8" %s��]/j#{N�T��-�`]@:gf�,{��ф�خ�;ئ��ME��`�![������������G��HvU���?�b2��66W�I¬��6�A�K٣��=̝����G���� Q�T�ԋ�q��4I����X�m�����7����R{�i8�g'����O�x�/؀���J@Χr��$��{n	'��~胲@h��ZH�E�S�UV2��o��p�����Lr�}�Z��`#2JS�P��%���L=���W��9��sjC�u{���T��)��Ӱp��&:_�b�n�_#,�_'�B*��φ���	��K�Wm�����6���ݝkt�F��7���u��J��t?O���텎��Յ��'�|�+����?�ݭ<���B�uÇ$,>�ձ��:<��,��TG.>�ڈH�ٸ��� B��W�X2��7��1Gx1�,֒+�x�ݶ�*y��׹.�F�u%:4̂i���轙��*+�!5�!t��T�#����i��۾��T��t�,ܵ%��>B^W�s�mΟß�f["j&���"H*"��g���Y�v�VS4�Oz�E�A�d\��?���1�2��&c&.S���n�%OV�ЉeSgE(�#�����bsUV j��8���N�����g���F��)����w��/>�j�>�A�>��b��oٝ}�-�0�M7����y�4Hj��/�gh�a������Пp_2�Ӟ��J׼tI��d���H���Հ�J����\
z*9
�1�:��>i�$��$ɦ�Bh��g���P�'}�+f(u���k�͹��નc��aS|hUȑn�Ekl=ʔ��y���XH,C!���7�W�ΐ�f}�����/�a-O$V=�](����:�S�WXeHS,q˄�L�0�:b�q�Knڅܝ�l���so��Ux�h�e������i�Bƾe�o�u�5Iq��#��f�I|�p�W�<p�k�I-%���ՎW�W���OБ��i��S n��8L��r='P}8΁$\l�s�vQy�	A�}k��ǀ�ĥ��|P��G�T� �Ҕy��p��W*#
������^FW��QX|����a�:��S�aI��"/��rV�۾�++�w#��T�@NuW��� S��w˙�t���翝��/:�-[_��"mi�y�Q�߿��!%��'��e�[�Y�>��Nל�8S'o���d����5g(`ҭ�3��)�}�3+뎴鍘��@/H�Xr��EC�e\���k|�/.�<V�aë3ԙ��`���A�k_�Sb���-��� ����K��!P��vw+�;�O�h)�3s�{���4Ox��d�/���'y�9Ul��:=��/$�G�I��\K�т�2⤯�T��i���9
^�G����q�!+۲e�M��n�I�ٯ)Y��{yלȰk�.'��H��v�g&��U�4��E�����ئ&��1���; ��^D<���ùOlC]|��:+A�~qfP��*g��@|A����sBXݵ{"vr���W��+�jqc��~b��C�ⷛ�|�6�]� ��'P���s�q`��hK�K8��]-�I+'�	i���qN��B:�}�屽�:i���"�if܇�t��£�kF�Wl��|��ަ���j�9&�K�fO��A%�,�2�ާA)5�=��8S~���2���ٻ/#���4ǐ��w���-]֫�����t)��������|ݟ�Hǅj4�}���J��}�D�]�����o)��;�Sx�E��b��f'�6�q�����#�$h�U���{��s��u��+� g93�r@��+O$zPis�иhA�D�y!H(B]V:���������6�J��YF�,�x��aG1Mu�I�<�����V����׸3#D�"��������:סST�3����w�&pI8LP�w���	l-�1�	n�T=$ ��&�KrV��C�C9���$��q��4��x����2X�����۶$r���(9>|�t��d��|��$���|�@�?��F�13�.J�$��I����!��$}�����^z!!���}Ԩ��_;٤�@<�3~,�]�0u>zvJ��>�n�T �~��p�2� ��Gz�{z �g50��8F&�Աra�!Vȏ�}�Մ?���c�X�����a�D�h>��|��+��?��D��R��S
�8��\z
_�}]��R�۵o���*���/B�ƶ�N,mE��`3� �D�8��t�!4��{ѥX��$o!�)N���D�S���>5+���QL�ZE�O�#��E�a#KtbX�&!2S��e$��Z�ehK�>[M��g2ټ �2ZM��
S$W�B�f^L��v�͚�#eqN��W�v�B��/0��i�w��u���Pq�y40eL斒�!C��yhƵ��@�ف����j谣}��Sr���|��2���@rJb����oF���/��%b�����R��<3FO'��*��4����$���E��M�
�c���;���d��k�V�����MP\��<�CA/�ɍ��8�hĄnh�c:� ���7��!����=���1�z�~�e�yc���ٙs����'tmӦ�PQ��I�+��N��!��+��K��A/Z�z���^�¨���`��B3z<uYm"D"&u�l��B�Z�1���,����<�K�Ÿ�������+BU�~�U5��b��])���L)Bw��U/']�\���Nzh���.���k-����t�г�A͢J�݇#����D 輁�q !ͯ�ƈ�>�5e����J5� ��y�x��k���3�hx&��(j� ����ފ/�q�K@Wi�&T�UOj �|lY6���PXE���^bz)�������q�g�)/9W�Ԗd�YX��eG�:
.#�k;z˄�86����(��͚�dK#�Xp,���lM5�}Zɻ���n��>
�%f-�<�)s\ޜ*������A�#غ��`���Ê|a�&0��&�C��nt��mj;"���-�0���+ܧ<�~-\8��RS��{�5�zbL'��p����N�O*�+�zB�&�<	q_����1\e%���{����2X��&ぺ��4B�,�/|�Y�sP����R󤚅V2/*G�&P!g��N��X܃&��E�!�6�����,8��b�	Tڱg�lC�$�ۈdd �6~����z�~5ȍݮ!`k0���֓��DIf�F3!���:6��M��Fc�/V�hoKp2F|��2�	Jn�C������Րq��`���ƫS`��O1s��|~�fQk��7����Q
� #�<���ĥ���	�B|>&
M�)?5��̕)r�c�A�aT��	��5�ćޟ�]5#�*��u,�E�ς�k�vRT��x�`��F��f�}�[�4�ݟ��S{��DK����jC����к�H`2p��)�x�/��ڡ�X�A�_#�� )V-޹�ޢ7x�l@ی6v9�o�R�"�)MTzǟ��^�K�������vC�����e�O!�����$�UB��-5�M4�H�����}5?UE�Oean����Ӓ5�8-��l�dm�fzU�IW�.���*�W,��4JM&�m��R�߿�Z��������Dns�a���?4[��U^���r�U Z�����h�B!�����2u�Ru�k~c��ѳ�,��'�����X���&�|������c�c��nV@J졭�#0%%�Tm��˜�)�:/�m��~-��4��z �C�dvs�"|���gt�{�p\�f�B�������<fU�Plj)k�*�V�{�	��_)ˑ���1����������B��X�;BsOh��6��uQ���ĸ��������v�{
#B~R������T��!ѣ���;���X"���슫Q���%���?��Tq�g 0��rbO�
-�㰺{�9�����gJ��Ioi.���Ӏy�`˜���2�Uq�n����y��Ь���B�'�'��+�e��Af�����ק�&��
��Z����M6XFQ��w�H��8m�YO�/�݌^d;�OM���1�,���M�0�{��&[M.�Lk�]?�F(�w��9�5ݨ%^����7��,.pz�(ȯ�\T�iN��ڥ�׎�k�zj���UB�V�s��~Aa���Zm�1�/����I��7$��H��(3S��B��z�=��%�A=z5���se>�����h�u#�L���!�.=<<~]�]^�	�y�>��Xr��L������X �~lw��{�H�&E/4db��UU	�{2�&��YUE���J[N��?6�2��"$�:)f���pyX�ɰ�;-��>�f�s���ٿ������l)�@�E�� �;�D�ʭ��JʒJP�q�0LT�M&�<��؅���cs�֍��A��K�γ� .=���@�lfrÕ���|c���i��ܠ]�fQ�wǷ�5б!�J!��w�Z^��ц� Fͧ�����a�|�
C�ʇ;�]�U�Mwu,�~�PnH��;=����8�C������>�+[G��K�bI���	�E�o{å��n[����4�q��jx��ĮCl�sT�/m�i+kRE��6��JԜπ(4,�O�Q��'7\ ���~AN�Ӯ�7�,�-��o�cX�v��/��C��JN ꏋ������pe̟��]��sC�9�I4:'�kI�M��Ѻm�v����
��PA�+)#~<R��e�"Cxtz�ӏp�ܩ���7ɸ�EbS�U2=O{ ����I����C+y&0#	|We �*�/ב�YC����S;����+�`���-$	�px뭫�����VVD�ڙ񋑛���y��L����$�Q����Jֶr�Ԕ�n��G`�����ư����¤���O�ar{�!Ϫ���nL�Lw�ߌ��?ߏơܰ��]��}J��`Gߜ1�����J�B��Ͽ�v���gFl���0���(���"�,��H0@���`s�<�J�u�(���!�R��v3�*ۖ�uH�Q�:�|�O$k,�S�eB�^Xx4���,�9�Á�{UyO
c� ��1�T���$9�tܘ��G4"Mm��e|���B|�h|����o�.�(���	���v�[�U�}-��3t��!%�/��J��~�3�֡���T{��͆�p���߹�c�&ڊ��*���!���r ��D cJ��#L���w�"G�۽��&��۱��bL��8�r!�\@HP^����jg1���0d�0�~N�� ��B*b+�J���P-*�
�ͺ�ޫ�:�6+H��xs�$�����%E�����3[?��� �s�	s��5kw��XM̻C'{�۰�J�����C�j��b�{]���Cgx��d�����ot*c�q��\���V�ZO�l�o��6+�e�	{�|���#d�_k��˼t����q�1:�/��:��e�7Ϯ
(���YJ��C�Id!��p�C@cū|'o2a�s-��g�6!��ʒ�
ϓ	� 
�tB����V�Tws�g�iQ�&��+鑨�7�D�9v�](9;&����6�:˺������7�i�l �ѝ;��<���;YeC��$O�ao'�Z8���pR�b"���/4��`��c��l���������JSӊ)��H�]E��[���/d�f��*�aE;ן�JS�)�w�\v��7�C/�!�T��i��-�+�M�o�詝ˆ��b^�kNNiX%�y��6�"����\����R4|�9��fI���8�����O����Ӭ�����J����2�ZѲ?q{���8Ɯ�~|_�$_��Q:���ğ��4��;Ѝm(��1��#o�A� 1�����	���J�I�N*��?�_]:����M������7������ֲ��Q�<aBP���c�Tܾ��J�����5"	����C�;$t���yW���e
1�p�E�G	_�D������{�L�_��Y�����70������#Z_�şl#}_���]������^x+�g��y�)��Q:c��N�{,�%��(������>�PF�8���)��|���GP�[׃�B��Y(�K�=20_�Oc w%S
1�
��ˀ�H�i>��@Q�B��T��*HPVapr;�HqN����V6>j�����q)�)g��]LC�w�?��0\��	"��J$	���n�-w��Z��<��_�!١cf6�vN��LP;��?[�ܳ�i�_K���~� �@�2�Pv]U��^tX��J�N��g����%���t*����B�3\q�Z���f����M�p�%��[E5(Gݶ���W�%A	��Q����u81s��S���}_�G�Q�<� �����p��2Ae��>�D�lZk�СG&0�[˵U����"��Y7G��f��aUQu�\�6�v�|1$m�og�V���%8u]�	׋H�2
�É�ΰXx���G��s�Zz��<Dl�?�y'vc��1�c��<��.6��^ٹ.�&w�ǘ]�s�<$�J�!��cltЀ���S麳��E7%�!l�M�i;ovo�ؘ��ˎ��A���]䎃�y����7���BY�^$�=y��	�>�9 $⸲���8�!<�.B�?�C:�朋�����m2�2��>��</�K�`$ot����mX�1��w�>���(;�m���B K^���H�I0|�e�@�H�Ep��i#�ł ��E0�{�S\����4�?�,(bJ�*u!!����l�s���'U'v�Q�����:iך���F�B
-zU�K�����������hM�]-cۋ�8���bp�A��&D��|�J>(��	9ٜ>��U_(�4N2u��f����;�ȍ�wa���Udf��JӬ,Q���ί #��g4�'n>=�~G�b�.���g=/5?�a��e���[�
�Bv���0�=���Mr�m��� +�k��7�2+�K�2/M[�*�Lo /�oJ����e6�c};�9|0�nZ:�d$*[���������L�r�V�aW�9��&���I�pQb���Q�\���L���~A��<:�"�Q~��t�u�� ���!�������ƭΉR���АZ�_0������V���r�����6/��+<1V������wlZ�����L�KTU[?.a�臵����D��2WA����`y�%�І���_^uq�c�uP�]�wX�M��4|���*��z�����`&����;��O��Шn2\���!�H�����I������{9�n�eS���x]���>����E[�H2��b�KB��Ce�z��c��J��g�3pîT�`�����8ݮ[o���3w���̄=��|��W�l2�I몽�sX(5ߔ.���q\���y2)I]%�y� m=�2���4�S�CW�^U�g�Mч���d���31}kő�`K�Gۙ4�����c�^�o7����5��&{�2�2����Yar���!��SV7���5���O�������&�QQ�EE>%���Fx�aFc�㮜����Q��îi���!���Z�(D
/���<���������=.��l6���i�8�wd$�%��(��,Dd%󤴙)%�$J
�`�MU�ˠ2p�x�L8��	�"�!M��R��w��9��L���i�ad`"Yϟ+H�06��jӮ�@�m?�q���u��h�f3�l3�e��f $Y`�w�K�:
4\b?}J�yg�6�_�SҐ,T�\{E�b���Φ�H���q�sѬ���u��Ğ�!{{�s�gɗ�*���^H�&�>s���y��٥T�H��q�6l�˶o��Q m���qT����]�/�2z�3�&�)�K)��.��D<���Mܪ��3�1o���,zݽ�!:0�0^bG'���uy���֘r1����A`ՠ`�:Ix^�}L��@%��X���Zr!�~�Zt�l̫�����'zhH��F0
(0��~�q�zgԢE�o+'Q�iIT�M�-=_�� ۬����7�
�� �Aۛr��dl��dx[.D.G���1嬋$�]�DufQ��rq�Z*�*8��ܝ�0�R�gY�)B���dε����s�����~~�������;�?���a�@�h'�nZ���Xz�����sWQ]j����NpG�=�H&hzl%� �� ����g/j�����Z���9+��^�l촸M�t0Zү����6���&qI^l`��Q̒v��r��s3����P�G#�� �H�b�	ˎ�QIS�jH�T��I�窛Gb{>u���+�]����/e1e��E��7����d�f����%~�� �V.D��e7;GD��ؽɎOd\��f1���8!ꐞ�[�D�'��L@,�����B�H8͎�˛�3�0s=�����Y����K����\fN�Cw,�,]�e�2�ɸ�e-��.t�0�܁):ig��Ӳ�h�p<ܕCOH��ɅL3�83]�\����%
]2��Q��"�t�z���*�^�QZ�=Z�灆�*r���in�k>e����@	��ǭ	�EiG��I���j����]���
�������<�CA�J͖J,�4$&e�=�T����%�Td��V�[�������g�|���V�V	����p��
��)B�
��B�g��t�#@�(���n͹�-���r4�d����%��0�,o�v�t�1e#Uo��L-�5������J5��) .��C�jAߦ��3XB��v	��C�D��=���3�J3�彖�ɗM
I���v�̞{5�����>��?tJ߂V�u�λmqi-gX}�/pW��rS�[&[�փ�1D�_��:/$&�����w@���:@b�pe�/�zyUV�wɩd.#^&<J��e�'����2��j���B�ӧ�8�g�v�*�ph�����!د�Cp=�����'+}@d�;.�B��	�X���6��g��\sr�s-\����l �{�`ԠM����ي�"�AawE��֚(L�KVTؠ\k�ʅ�-[�qg-n�si�$֜��7z�n*��f3|�Q�9��'�!#� ��*/�(�������芕=���]�w�R՞�����Ovա���
pU��Gaء�	�1�E�F^`����zr�XW�=eJ�C�8}L����}+�W��s�\�6�<����E�$��<����aD�Y-����Q�p�$&�<¬�y$�RT�
��i*/��k����9K5;W�8U7�j�K��f��1P��s~c��:�9{�h\i�"\�j�����	嬧��-������hoy��D���
�eXE��i���`V�*�8&i�o-k���T�Bl��9%�O���=.�dқB�ͷ���!�qw`ߵ�=5�<?����8�ȕ��x��=�S���yws�,s��)T��q�|��M��m����
u�	o�{��Y#�RHa;�Uc�������ֆ�4m���h�g�qO�����=���e%x��H�WO���T�W����~�B��%>���͂�\����	�C�K�0�P�3��iHn9w¥§��\���z��c���B��C�y�K9��eA6!&8	�����6�߲Һ-zm����*�!��|��x�����S�]��Nί??ƣ�\�:��^f;M@��ʇ�{x~��5
�Y�0N �����=�}�*G�%�e��RaϞb�iZ����xɉ�+I�%����v|�x?��V���Z��yƳ��w��C�N�ZHe�q���q&`�T&�.ڡ�o1"�L_�.hz��� �+��E�>�m|�I*+@��Ek���2f��FW.�T�� ��¿nhT����хlF:�W8���ANӢU����V���+��oڋr�ܟL�^�U��HD��\	nAa@��%�`��_�d����.M�y�����B�����ӨLԜ��#�w���
h�3�C���pR�2M$��I��:�Ep�� Oي[^w�wBE��0@�10������xycW�_�i�u�w����팰]D�>��7��� RA���,Ҵ�t�T� ���S�kRI�S��fFlQ��F�������~�n�\L��JP�?�q�6���kK	��BY\����FRb�	\9[ޱ����T.E��.�u.���*�Z�fp�����I�(�de_����~���#C��+Z�XǴPQ�� ]����Y Y)��)M>����n��e�/�[	5����b�E���`+���~:�|���o�?u*�ܸ)�'�O��	~0kmMRM��$]T�5Dp����T DEoJ7
%�c\>)���}_ 1�*`Y��.`��bq�G��w��OA��������ދ��F7�aDf �ug��v��m���r�\�J'EH��Ɨt�N�9�K�=���X��8����Z*�_Տ�1>9��,���xB��M��f�Q�O+�m�C�hp �(t%0����rǃ
�[h[�x#�D�M�����ytR-,���|$��@G5�e̐�Q�<!��y0F�B��^J�vGmx����B]�4���a��|� �L�,S:*{n�)��@,���3��Q?�x���KOg+y�M[��}U��z�<�@�b�
cM�8Q��Q*�Ӟ,ob�>���%B��B9��l|ԙ��5����6>�s	��IԞ�wHR�S _����-[������P�K��JH�L�?����O+�rO��d��d�p!J?NԌԯ@[u|���Ŵ�I��K䓆qL�K���u��a6��S��}�?��]w�~X�=��-H��I(��Y���)�sM`�&t��p�t�G�3l1vC����i[5}Nf��&X�@&ߺG��߻������L�G �j9%�����N��&Q�p�":��u��8�T�"�plg�3�� ��5�  �{z�z,xWf;.�J��P�@Lg�`kH�c�t���`ǚ6�ܿ�+a����f��&@+�2��J�$�D��!�}�*>>��v��_�7{�;��8�6���ſ������* ��ꢇE��Ǽ�e���X�Q�0Q��y���HV�#�P�k����΂���]�H�6R�-�$��34�M�9n��盢`GҌ3��/m�c>fю�ҽ ��F�&����Lg��h���O�p�^�r�b�w�9��}��{��;c���<G�s�}6e��ʉ�%{n�O*����=��-��̄��D�ց��VЛ�p>4�|��U}�΋��Z�����p�Ly���V1='��]5j �Fګ|U[����40٭pi۱�����2��l&�馲�e��F�	���� u�;?�p�@��{��nS�Y��ձ]�,�'�u�����|O�Ӕ���P�ݺ��!�,mv#��[�V��_��6�Zb�����G�F=bUU�Q2y�}�d�8:?�|�x�댢��<<0>Z�݉X=���P�;{'qˈV���Ҵ��F�*�$wp�5���Q����qmW�Ǿ�o�̊�դd���������2	�Z��Vy�TR��gj��^z=w��㈪'��ϴ2f�:�����`�Hm��-˃<gztT\hFX������eoyc��3S��g<_mU��*Λ���i��as&��>����#���r��/;��/h�;|A.�2��]6�,��b�}r�m׶��X~G��\[7G��\�B�׸i�~�Z_V~1�HdK��5�l�L�<���9�s~�I�G�~�Eo�bAf�L/����X�~�A}`:qR�fU�(�5rp��萫g1n����x��Em\���N�8�^W���K3�>���a�\9�9m�XPz[���cT{��<k�T16�����Z���t3����;@���A�-UU�8�yUP�P��;��\�oO5��ڕ�h;e�o\6tp���c�t�FZ�/.g��S���iH�����\L�Ob8C���м�Kȓ?+��?���
����AA���F[D��'�)��V�t]����`
姘��:�Hz������3Gh�Z��B�rO�Ǿ�;B���Z��L.�<\Q3�A_3qw���ÿ%�ãe��ť�
ݦ��y\�p2��W�]���]���}���$�l���ZA��`MZڭ�� R\��u��*���4�q���"=�6��H��}"Xl]��_��VS��B�`�rE�y���V��2��] �q[Խm� ��Á#O(��c1�5w��ѽϜ�F���v'�n��Z<�)���cp0��h�/*��
�qU��c��T��A�02�*���o��Ni��'�	�~|[,\��ʏ��Xqn��__��s���\?��妥�.U?�����e��K�3��d�%$9U��� n���t��,��.a�_R1艁���̍Y�-ZH��H�5�+	ӕ!²��ٗ��%�<�n�����3�OsN�x��z��J���dh4�Ԝ�n��}�Y��>b�?J����ꢈ��Q¼�����9�RZ�f
���s�7���H�>yHL�`0Nv=u�;�Ok]0w����>p�,����y���{���4�#~)D_���SF�p��Xv�Ֆ�5�Q�_�A��p��)�R�ҟM1��Hj�k���#��s(D�a@)N���p�V�̑���� _̖:� 3��O�c ]�$��U��b)Z���n����K^T-
�Gs(TH��1�8q��Q�u��E���GT7�)������Ğ~�X�KH9ʵ��'��k�$,o��E7�?p�;|6"O��r7��%yWp"U��l�mmG)�TϠ��d�p%Œ�c��E�>��EL"sk�7�]�����RB��'6��хÿį����e��T�,1�kFL_E�їq����xꥢ��+"!�����ݙϋh�HCP�4ű
e+�|�i��	D��zL± �/>�{�AX�o+�Be�C��OХ��H��)�,���-	��*��ؠ�D�fa�'ۡ'���ߢ�-� j1��w-u|�11	�ZD�M�%�z�y�����,�Ɩ9�j�H1|�����h���H�$䢂ه�"Ͼѧ�ⴟ������V�,��Қ�K���q�3���������W��7g�(�j�$��&u���d�x�
��î��1��;�u�ܤς>f:�� 9F�鯜�}��w,�[_����8&?`�	~�3�xi�(T=���r�%gF���^�Ƭ��^��T���sk����n�k)s `��Gv\�]�=`&��e��c���C�n�;��V����/�9Ӟ��F�����	~]���qx�M�	2��ɫ.�-Ȕ��xUpW)��(�Y�,{����C�� 4󨊿�թ��#�,��%�Ãx�ź�u���R;/�!�Xwt�7�&��
i |�$@��/��ݾ��(�e�{��Ib�)xnF����� З��*o����r����ú��bi @W��(f���쟄��>F�.c�2�}���1��Ԧd�|���i��	U����#ǁ�v¹�0U��M}�1����ID<�ϰ��7fU?�I/����w�&��|�6��>P~t�bt�b�f��� @ع��-uv��K9�Or��&֛O����s���n�6�� �6��3��h�zz�F�E%�jy����<���4R��:�g-��us���ﰶ� l	�@d��sa��7�VT�_~�<����C3�F|C�%[ ���Y�x�dFR��܊'\�h��
R������$ly���*v�JIğs#����ڞ�j���$<�*��v*��A��D�qC��*��7�)�¢�)��"{H�3�=R{�����Ѧ�s7)zѼ�i�p��~��~�2u��%�#C��Ub�Y/ٕX����GE�g($'HHn6�k���G��컬<
Lb��*C��e�5���y��M�����A�P�k�Z���Vz5��#��Nd=���3B~�-����R;�}��\��x�}?hg��-��vKM��%�F|!L��2��a�lև�p5Bar��6MK	����ׁsKb"����{`H�3��M�N�T�A}E<6��%�n��r�_��?��. ��
�(�eIY�UÆ*�pgN��i�P���;��ăa��I4��M(�ږ&������r_ʝ]�
p���,�`nR�{�DЊ�2d4�H麦/��;-Rz(�=����������u� �Y a�' >F3�A�����W������y3/iZ�Y��8�f�.���C��>p����r{�F�F�{%/W����Zp���M��i2B#��$m��(q��]�w��/g͑ɚE����`߃mG���$�Q��r��U�����g�[�,�B�p} ��Y#�Ex���قh�1Sz>�y_,#|�y�Er�j���YZ��h5��\�^�H"{r'��rUBg�i߇v�X�]��/�m��ه�-��oU�F�6op���]ng�(�e�����%N��X�®d\·�hxxfY�b�T���$�(�����6إjR� ����?�ӊt�� ��,j�E#n��C`��]���|g�݃֒ɷ{aL+i3ٽ��ȿ�R��a���4�`��-��s��?��L��P�ҭ�O4A�ZWT�Vb+��eT�:�������~�v���})�<�����]q�i��a�p�b֌�Z�1�s=�;��V��B7�B$��ҩc��79�%USʈ*����G��7�VPm?B�轻$O���W.�}��kd�� �1��\�]�ڣ^������]Q�(�9b8W�K?z�	O#�ܔ�	�wpq�튳��C�����V��#�
!?���Z+����*L̳��eN�1X��7 ..���sa]ம�w�"�i��b&�mrw�Au����ec�Ѩo�3a*�XS�KI-��];{�{*@�^�"�c�^�S���K�N|M,���t�L�����U�{~�����vpf��b��^H�L17I[P��-'{��'�~ fi�]���:-�~��ay��	�b�m��ō�T��(noV�s�W�"wFb\,ā�lN3�@N�-�Dmͽ�6��Q,)�a;��}�����4)~��[�4@�:��P����Ze�D�*�&ֺjk����X+��p���Qu'oT�X-y7Y^k§:y���I�蓪��U̥v*\"�?(��(����\"���>�1�1�un>D�\���0��!�K(�og@0�m[��ʍ��̚׀�%~�*H��2�u�<.�O��O$i`Fݘ/�T��N�S��~���|A�)��nv�~�|��\J�
NǼ���O,h�Ѣ�V����kVоf���@�ю]�D~�zd����o���F<���a^k�:�(ˍzd��>�چ���wP���*Ч~fN��N�l�<�-H����(�b�QiC���j�iv�0ĿJ��r�x�E���e0S*3�
�w�����	��ה���h T����'2#�HU�@�X��!"�?4�o��1N`��&�[����JǷPEO�?X�~��\������'��9�����?VX�Y�l��c�6�ēXX�kS�lBYЄh��N��w*d��G�]�����l�j]�Q�:gM^z=-��]�n���<7�.����Q�b!B\�Y��m�s@-�f�p�z�����q>v�J��%�����u�$���Ak��6�u�h�s�x�Ň�#��svv-��ԩ�gA�S�Q�%1�b�:hA����hy�V�H�~��p�G+��y�}��X]����(X�Nym,�7#��G+�'��x��"QAW�IG���$5`O��B%q��N�ތ�5�=�~��
ߨڨ����m�R���0���+�w���?�f���Y&��w%�AbJ��w��������A)8듰�"49�ky���Ho��'�m���i����y�k��N�er��Nz�%v�| q: �S��qEQSZ��q��D��+z'�r0����o����R���1,C��z�2�2��l��ٶ�r<%|�يHm������P��:�T��� �o����I |�VT���9k(��,��5�����З���>b��N�6K����t�|��p�d'^`b?3�^��h";��x�����B� �Av՛�$��d�N������-YMO�ah�'݌��m+������@P�{�Y���� C2]X.<�`��EXW��K�CG;s���q�������)?(tD��ҌK)��W����
խ4-i]r):� }s߸��[����#F��е��K&+���?�X��,(��5l��E�#˧	��j,!t� ��s�!����jzʛ�D� ?�#>_M��pg�0{�"1�nb�|C��G���Y^)�kGe櫁�����^t@������$�޼\������8�k�A�r0��%�J��%1�������)�GWؖ�٬�x�w��H����Oi_.o�1$^�R�D��?��Z�ꀧ�XB�'����i�Mc����2�׏��SI��-��Ú�MZ�%�e�	�a�bJ��1�o�wuJP�C���\���7,S���!D�S�`׷�@�){��f �V{�Y�!��x�Jj>2��` %�/��o�{r�i��:�;�T�T
 �m\�}#O�1�\�X�t:���i�C`�Wgq���j��u�	[�{jݴf���y�}����]i��NB��y�u%��"���B�9�p�����ą
�jX��5OݒO̬��N��m�z���)d9�����db�⒴��ع�,�����@L]�>Pf1����e���鎟@��BE�#�QV�A��<'����t�=QMԫ]oTurK�e�9�.�����:e0l �+y��[%G+ ��YE.�AXw��]�[���O8J���GDM+�}�	�2��n�l/�453�E;y)F=�YXu�R�%��F�:��tQk�v��r��U��޴�k��Ӆ�í �t��Ɠ����c�*���(��%i(	���bE�����&���̡��:�,����;�(٢}�<�C&N5�wx6[���g�~�M�ְA��y��x �����T-Y�c;w�F$0S'Q���R~N�����d���1�<�C0�J��?�5X�y���9����򋉤:x:��b[ݓ3>��f:���ɢ�_��\Ə߻H#K�M�N܄m���I3]+�ii*4t��z�G�8�m�QQU�G!ʐ0^P$�R���>1��0�	l���0����}p@6�[%�S��_�-�{3�	?a����
�w��Boz�kf�iNpY/�_���>0��b/U�;Y\XS
��*W�;����>U�"	�5wј_/�Ħ5�u���1ْ�	f�G��}�g��� Ƣb�褔;��i0Pt���;�[��*���6u$��e	�)�B��sc6?]fn����p�E:�H��� }��Ϝ[��qh猊�N�����M���p�p_òY���?ٯ�bG-yH��9D�qB��g*��Qto��jT����(K�fAz2cȪ���M��Bc�\^NGɅ�ph�����5S��P��BM5p]{Y G�v*��S^6s�7��E#���ǰ�z�B8��~���?K6�3\|�i��8H��51�:?�u4��eK�p�K���HU?V�靳�>T���PU�����n,�Ѯ�3zM�p��tY��/!���E�vo�q�}T=���10$��~Y��B���&��Dp}.���{��b���=� �u�A��{�1y%&���3`��L'��-����|�5�-�)��8�a\��2�^9�P��<TLHґڶ[����,����I�3L�%���'i�����c�j ��O�T.O�h�]��L�޼r�6[������l����,f�K"Lwޏ��SJ�.��\.��;���&ִ�I���t?�a��ޫ�`�"m���I���*�l��F����.QUB��`|w���=-�LZWd�H�8,a1����B�~9]>���v+��]�|�f�N8�A�؍�,k����>�x�`K�Gu�q��0���5��I:S�/x��(�{�$�nw]��i��v���c�R�>n���o�k��V̀�����a�ơ�(z�F?�έ��Gw����v�
�|і z���n�Z�Aw[��躥V{G�F*�o��䤉+���4�9����.���q�a"�~��ש"X�������<�$���V�7;ʈ�Nn�%8�D�=�Q���V�֗-b�R���i�%�8�h�Ý'5o��)�#��M�ca]Ǜb�>��1�K����4"��OS�Sĭ?��$|)�Nb\T�X��a�0�l�:�NX����?��DMc4��`�]� *�����5�Qͦ��WL-��K�ʻ�=�T���ߊEzβ�l�׀�����4yC:���7��(gi�JIE�`���4sC�^�t�al��z�{�#���BB�	[��\cd�%*�Y�j�\R���A��-I풾ˮ����8�yxy� �g��0�j�i�tg$O�մ5c������i� �:ʗ79�̮��צ��b�C����ǈYF="���f�K!�!��3�Ť({��`�δO�S�e��L���mb���<�[÷�Q����b�i	CH+�����ם�m`�_@�����2 C�o���EMZ2��'g�כ��8�H��Cs�N�bAs�7/3']؎���í�hj�z��?�9`! �^��p_�-��aƮ���EV�1�� ��z�[V��K����%@����U���; I��� U���eփ�ZV�� ��oV���Lko�½׶�0=Jz#]:xO�aK�iK`hߥ�=K>�7�w&�7�-��,�U�B!j���̭�}zk�;���4�����?�u��V�?�9���iK��|Cʚ�{5dE&��(�KL���~�K��vaņJ��+���/���za7Ͽ=#����wB�R�ĻTx$�;�L�?�OHS��5R���Ԙ�yՏ@WZ'^E��.l�op���~˷�qeѯ�ё5�1���+��^��*)MiBj#bd�}R���?bΨ;��3t.-�!	��ъ�� X�&^�h�;\0��W~�e�0��f��k��V��%�sǟ'�1[g��=ܛ9����������s�މ��l-�%E�!�J�����?<;�jB ��)�`�0���햕�V�����=�`�Iٷt�~R��v��غ����PuXER�B�Jrl�F�<���J7�U�ւ6����}��'eR�v�f<����kU`8��5��XK@`���c�1Le�&�q�Z��t�i-�%���c�?�^Ř�J���	��M0)�7�+}v�0l-�zno8�)�7����=�����<�տV�Ȏ)��aCh�e���{��ZdguAL#�&2��	�i���Pm�'�"��j���@���?�z�#&��3�b�s��$p����Җo+M��D|KjOXڿ��-X�G�i��#��}���D� bM�#9����U/�-=VXGY����9GM|�^f�}l���2j����_��e*<�em)�2�r�_k9�MtBqTH:�^16�J�"�{|������}�{W��Fj���U��������YZ7��4ߖ~��d���t�D�2���0��c����8���{h��7���I�Z�c=X�譤�Dj��w���"g��X�	�$��Xoo���.%�f4k���X��o�c`�]?��B9���q�|��$9�ֺt��s�!_rtr装�؜�� :�C���߰h;]��[�}�M.�A��o�d4�h��
����-����u���,p�34]ϣx�(Q"��p��(nc!�jS�ݶ���6� �:�2M���;S+�*@�7�m�
˱�§,�*'m��qvs+D�ީ�!��&#�+Х�^{Ԧ�_�k���Į����.l[�+t4�ݘ r:�Sl���S���o4J��W��Z�������;*7?M#�G*fwav����A룩{1PE3/��!hL�τ�bV�����'-..d�����S��;.{�@ʈ���-��xU�3��N�?$S/i5�g�]g���#�|d-u~n�--���������f�E(�4�a-Yk���3�@.�5`���ߩ��~&�Ja��~�$�U�	����j�x�.�eʇPk��a�W0XI�")o�JW���N`,����ao�WRB�T1�?#�n$����k�z�ᵟ?�;Dw�7.���0#�bO�jЇ*['9>�-����|~8CDd�R�4�� {�3���`���l���Z>'�W��|w�1>�õ�K�k�(�a�̶����$�z&�Sn�`��|��/ �C�z��W)y�������|~���/-���sqZc�J�q�v @4��_��Vy��ڑ�P���X�SRXsP-8��"y7B^�/�N"��9��W���SST]�s���(l�� �s�BK��	�W��
t$�
��ڮ�`���4��W+٦��.���pe4���4�G��Q�(�}�D�
P�F���KI�L����P.�%��ZO[�>q�F?�b��lu"���T�J% >1O�����P ��A���0ى7�ωO�ѯa�*Z���"2�Mwuc���n��h��	yE���5�^��8_|<
�Й}��i��x;��_-��y����;�{�Cg&�漢������8��j=A���99n���*{�/��(���rq�����|ԑ�tlˬ��ׯU����o�G��;��yK��Lg�v:tQE����:Ӷ�э��0��bb�zY;~.���e��3%V9��jP���%�F:,��=_�>h�T��"��E|=��6g\��� �r� ��>��m��7�0�A�M�+GZ�O�a��bc�������E�^:�=�4då���c�J{�M�с���
�%g��`<\ҥ���m��a�C��-� T�,gN��.3�w����K-��aM������ب��'����h_� ��8+\�ނ7��ұř}~�XXf�K ������É��t�>��D� =�=C�%G���*�b�#�D�k�9���X���3 "�fR��J&0x���B���"�(�ġ��bT	0$l@�Ur>�	�y�MN�8�$�24�?����6[P�U-�'��`l�i��.9�H�i/}����	t1�������i�����p�.d�nV{�	�c<�n��&�mt��g��p����'?�-L��A�G�SLȆMO�j�	��M��`���]%��Q>�3XO�� �\i=|%{oE	���QV�\1Q�"���t"�BQ1CB�����1��[�RFo'�6���/�H�q�˾jVD5"�d@��_��Y~@��V\�JDY?������%p3B����?f.џ�/U(D�y��aJ��)پ���hH(Z�T�y�y����<��b͠Y�T(�1���q�2+�v[����p��̒9t�Շ��6�(k��Ȃ�������F](��Ȅ'���l����8�˱{m.@�i��L��d�{CG���l�k��F�����p����wb�Nk�>��EB���}���O��n�'��?zz_i�s�`������5u �ѳ��28Jl��?�\t����*��~{"��.��X�Ʒ����8����3U�9|�$ʒ�v��'5q������.�O��_���j����+e�A�5��#��S����{"	q/�o�k�Bw��	V���{�XL�xl�Ԃ;�דɔEOEi{b_������{+Q|�Z��r5�:Z����ö�#�ɮ��I�,W1ScD=8X鮢���ξY��{C�2�'/�lvS0󒷆�We˭7��T���+'�CzorR˦5��Às��8�B�N�5�(��ڐ��E���`��Y�!m�W����Cp�O��\�{vQ"B{��ХjZ$�]t:�#���d&�8�%>�z���b��H�hyvy��p�����]��u��O$pX����=���3>z'��o�b�hQ����V�P���3�7 ��K�r_��"�|�1�%d\��P�+��x6tG�u�m~��=U�;�@��|���{g,�3O�6[�4���W���v1����I)?|�g�o�W��N�_%26J|v�U��Ƨ4(^Q,�
Z�@O��l�h��)ik����[��l"��8�j�8�S������u��X�������[����n�y��N��r^����F`Œ`��07�������Yh����n(.��9˹�f&h��'i^FW0�H8	�eZ+�
�D��2��ph��A�d��ԫ��Y��LE���ݗTAr%꘴q ���"�DC�e�'���u�_V���^�_��^ 3�'~Si���z��k��l4��a�	�b"�_���vp�4{��kJ�S�=��D��,y��b�)���:푱��l�^$���F��\�p���x9ma\�\�1�[x!ܝ3,��hx��)Ң��k��d��;$n����ŢXj����0*�5JZ�v���������ٌ� 1}(%�@ju��ǖj�������_��g1+|]ڌ��v:\� |��Wύw�X]��C��
M�7���(�Q�D�l+� #�XJ#]�k��c��}��`an���I+Lԋ�m�2��3Q)��`��B�u��㤢��p�h�J�{�����V�����~i�%�ԛDU|�k��Ui��X� ���kh̎���&'^�usFJ:p��r9�S@mTG i^�(��=���#�T��� g[��_�;g� EC0�9zJ�0��ݠ������1�dj�g�C��4����D|����ɨm=�7�3 �18�$I��\��y�P؜ДjȪ�ȭ{��ޟ�j���K�A�>�b��׈=�Q�_��_��7��b`摋�c��*2)��L_-e��Bz=<��"U���1������I�q���|g�}�󭀗aP�I�԰a0�2D�����2	G
�g�r 7j�棸�����=���ak�d�(݀͏�M��$&%�yl�n�4�����<-�(;>wʫY�O����T	� W(�m�߶}�P��ȕ+,��P��6UL���A\���V]oy��t��f�Z	<E�E�З��%,3���܄j�,�v8e�L��������e� �ߋݹk~RZ�E"������l��A)��v���PwL�x��t�0n���m�R����ALineMi?����/
�!����aI�C0�s���Ii���Ʒk���!}Uk���� X�fgp4��\�h�룾�k�r����|@Ջ2@�@�&��U_�Sdd�o_^�*�'�j�J�d�ܧ�6I���U@�Ğ5G�;_�������t5ė1�=9���u�Em9�M��jF��6�`�zH�$\�(���ꖛ����dU���A���7�f�b����{S��(�*6A~�QR��z݃�(ay�A�s�@=��s�?�����R	o���r�{8 �Pe&{M�g���ԂF|�L�wniqI�~R���ʈ���8؎>�Xl���sC����Y*��LY���T�&������k�H(L�/�BCL����J�r��_tKk3��&�;Ȅ'7�1�NAir̂�/e���m�5�h��ux���W%��S<�fD�ĈB�����2�	���GDP4k��K� ��	��xZ��U���մRr"Ll�8E�u���."j��i%x�������mr1�s�2K�'#u�f"� ����뜊��1sZr������A�-����`_Gl�aj^T[Jrp�,^���p�"n\㷁��d��Կ�m$�(
~`��w߬�c�T�B�6�0�ߑ#��P��
D	�u0w3�2��7�T����x5�lŢXF���������`2�X���@�,i
X�g�VktN�`�f�,o�O�q�(ˡ�Z��qz<�����E����L4������CX��8�LdR���7i�I�}�jzE�����}q��xZ)�d��@8���X��I�����#�K��T#cږ��le1B;q�b$������ϟ@�+������:�l;sÝ� ���ŗ[��K�
e=�G�1͵k��rOH�*�~i����!�T�⨓�{�� 4L�N��)�mt�E5 z��>Sf����/���G�x[�!����m�l�����!��#G����R���叴��_�ճ��f��@�>m-@�ڻ�x�b%O]�� �eK��/�T����s��p��L�\�e���!#��[��N���Ҿ��5�����b�ͫ�WٞA���&�Ύ�,ƹ��VZ�N���<�~�
0�������qq^%�����N�
�����nT��c�a0���{f}�˚������G�Ǡ�JW�e�����q��:͇6�U�����c㜌�|s���@�X
q��ܼ���#}I��0To%}�c���r�IV\������\���;��6���5V:��'�k-�U�w�gz��%����T�	&�&<_?-���P�RA8YH��}bO)�x�=*Aұ_f�������<�R��b�	T��T�Z!t)��=h���0|�����>L{��\�|�/)Q=̹`{آ�ֽ�s>���/��o���_�ѻ�{e����o9΢�e�U7�)���R��GM��sΰH�mw���	ݿ���:�/����׻h�?���J����Ul�e� t=:9�}�x@�㜬	l�d!���Ekʩ��{P�dc�w�Jey_�?g�"�	ڀW��I�=�~�t�A�64s�3��ԅ������5�*Q��V��H�=ޏK-(�'�ّ?�I^�4R��`Y2������9:Aue'r�>-����q���h�x_��;$O��u(�6O�( �Qf�oT�!JWמ����m��ԁ{���6���{���Ҁ)��ܩ^��B���C3�Ƒ���p|~�P0oS��'�>���.��i�@����X�Tzܪ5U�]^��x@�/�	Y��k�@a��B������ی�L\��62f���o���*�J��w���I��j�w�����"ή5�����(�?���<����ߎ�?��a��/�t�}\�l����4�
3	'�б�ڀ�����|���8���f�{֢��C�q�C�c�p���НQ���|WuY��u�l��K(y�!A�Vc� ц	U��s��6G��o�]J�b-x 0�cTuW�h>���j�z�i���/�� +��]��b���2|%\q�{�mo�l�yl�fTX�B���n�����y!���*Js�s�y֬��Aa<U���p�Ȧ]-H�:@��Y�K!�_2����f�1����*�)Y�?2	fU(2b��^=���'K��t��!H��%`����5��4�[�X��
/٨�3�`�pg���ĕ>�Sґ{����M��{���5�^�y�GV�D$p/���Y��gz�R^xG�f�ڍY:��S��㿓3������S�+��J}/��0=P$m�n�,pe�Bl�ξV��;щ@�sFJ�� �:��PZ��|��Z2g��0��l�N��}m�Z�m�F�I`(��{�A8�]*������/�Lh��X��5����K�˩~�E��P�PU��|�Jo���Wi��+�lS��L�K�TȮS1(��(Ͻ`�-f�ܲ!�74�XI�cْ�j'�Y�6�v!���pʰ��t�Ҟv2��YB&\��|��>UZ�A�m�G ����4��UD��K�DJq�"=��g�7�9�);�I:2�O��P�B�r86���Ӈ7ۣM�r��>��w����q�|�e��l0��J��q
@�oU�g ��뢲D�Dp|^�<qq/;j/����ۼ�G&=�q��W��^ue��# η�y��^���!qi�3���s�Qs�L����g�+�������C�jPM���.޷c7�bղVN�z���@�,FL0�#+tS3��$�,)�V���&4>�|Ņ)^n�	��O�#���T�t�hg�]��R`�����=z��hp��M�ba��p�Ǔ����*V�Ø�X�3��UV�b|w�w�j{�����;���
EwbRHȴJ �3���-�i��u�UJy �=ADN&�o�OC��AY2� ����s��e�$���M�c�R��f��/�ߛ=��S?V�q_��|'�e��~�3�p��F���Ekg኎qF�AZ�`���滶Ң`��i�wz��S�Ew]��%��W;Ť�\±��fSXz1!�1�,��]�+�G�"�n�c�=�l៱9��<ogR��'��,����i���ˤ�]L�B)sP[�;����;��+�K×��8fР���#4@O��ڕ�U9Fj|@�b_x!�}m���f*5C�=�D?���T�&U&�1�*�}���V�]�;��lM�Z��Bֶ�Ӊ����H�l����2x����v�u�_:�r�+�z5�Q��⨧w�)�.^���\<y B'���OH��,�-b(�&�m��
	��X�nK ���:�^A;s6Q5��sO	j��7���+L��c������A��o��tT��x��Ĭ��U�.�2�s�E���SR�͕HD���Z(�Ir�vw�e�3ޅz/j2F��/P�#> �A�S�mε�)�6�����8V��͋�� �Ҩ�LK���g4S��SObB��uq�b=���4��
��Z�s]4�y�ű�F�MBK3�W���X)�4�ۍ7�f\��`v�À(�ܲ�O� jg���U�����H?L���I�<���@H�:Br��k�0L���^�-l��U{�U�zr��!'�Mzhu����F{@��V�)ٞ�.s����+�d;���%�� Q!ͮߤ���}��Z��%�}�Ë_���ڐC��k������K�\����r�!�)�[��zk���V?��� 4�+�B�>f/н�6�,���TN9��̚�~�j��gt�|t@�d;��H����f:��@J-T�7Dd~6i?�8��� Qg�{]n��d��%��nk��m�����o���D�C�锯t0��M@Zl��V�,��s(�Z�޹���E�+j�i����k
R�trϔ��MO���AԬ�Nup���Y����i������t?a����-�6��<�C�g�2qn�Qm�`���!��ۄ0fB-t�2;�*�i����	z�`�G9 x��nS�qثp��^�I��Ɇ��m��<3��U]���?s|��^�yN���[pU��Si�^����e�;�f%!� P�ɭTN�PJM�4�Dt��CYPѪ���e�j��u��ʲZ�ߠ-t�̠_���Oΐ=�p���P������2��!�h3O	"'�oJ0�T�ڊ��W���`
����3ھNH�!�1g�=�ۗ��1��ŭO!�T��1NH��[R�������Q�!�=�۸(Ȑ�de�'��I��*����bI��I,0���O�l�QLj�&m��%�5���5��6��,(�X�2G�e��iHXziօ���ԇH�8P�­3eF{�e��-���¤�IV�m~j(���jla3
 {`�yM�>Y����($��(VI.JC<n�]�L���xP�ٕғ���U�W��Cx�P��ʗ�U΋�9X�J�-Vb��j�BZ�g�@���^�ټD(��ƹw�rV�з�ɑ��������4�i˺�jT���rJVl�g&�����c�A�jhD�+8d��4T����r3�MB�,k�ÍL�ڄ(z�M���6`�Q���(r�_�!H��;��b&f��z�硫 ×�	Ֆ]��J�)_�������B���fNv�~�I�p �D����ٽ���qye��� ��lV��ƚ�u��,��ޕ2����E��
��'��D+�h�ĦgX�6	���N�7T������-@��z���Xb?*}�t3��6̠�w�B���Vrm�̼\Tx����ז��������Ϧ��?��oTw����ڑC`�fZ���N�u��R���|��:T��[ݚ�}*L�4���*�7I0ǎՓ;ߋ�X�S�V�����9w�8�&���&�!�N����4"��Z٪���M�8��~��V�cơ:J�m .��d�ֶ�'�wj�;��w=	�0�-�\����&�;4�Y�s]��ՠ�S�2���NWk���Ϳy���<43����e��V�1|uVz�����I?ӅS+�gE��ohAI]+��<��h���(�� 3NHt�o
*����-Y6B�v��,.ܴ�V��<�6��E�&�p��@��ñR~��υ�8���WP���;P�@�і:���'����Ɛ7D>�Q�6bcM)�6��A�l#�=�ι"���bP���P0��y3�F��Ui��Ì�H�zN�[F J��fޙWC%;K�%^��}�y��n�X�e�O�S�əc&;��`�n��Z��8{LRQ�
a�{
j�tg�!�������.�u�+cqu���.���R�ғG��M�4:U|����?�D`T+�<����.����+���K��
}/��������}lA���Ht���3o"͹���ȴ�9E5�+b`jJ��o���].S�UBH�,C�w�����q�������� w��d��c���Wm����"W|+ -���'k�8�9I��4�{�1�ķ�m����7�~��$k��m�h!� ��N��_�$;��]P\�f�7�B%ԉ���������.�ŋ�xX�Qc@�z;0��O�.�W�8#�H���w��E��;�A���RUiRݯ��Z���ۅs�g �;"n��C�ߥ�/}�@Jd��^�?�:2��g�����;�\��J����d�^��M���ۍY�<ޚ퐻���I6���z���[W�hI���S�/ϿSWeVa��l��J�X�SE�DS�����x��lv��C��h�W�ֈ���P���鑳l��J��˛f�NKW^GeGE�<+�'%*h#�����5@$����azAI�L��']!	˿)���Fu�:���Y�ؿ4,�,�!,,ϔ���J�4h�G=����E�P��ÑE��t*����79�x,٧��S��{��I�Ah&��lߏ~UJz�S�5��[f��8�o!�0���������c`G�콂� �gp=Ƀݚ8+x�q=�H�(О�irמ臦���j���h0�ǂ�^ZI��IW"P�%LE�g,����+�;�2W'#��QR���-����ʴ�r	(G;o���6���EG=\9��.��k��p�9K�b�����%B���+w�G���y��O����������_
����D^=y�|`�X�%=?w��9�C���Xwm#�'�do��äbO�*���'i�������1��Q+2�ũ���3�+y�����hǴq���0��ƚ�S�v����w;�s�̄p�^��XZ=�[\ʿ煫0���T=�|�-7P�oPW5�_����x��+���@z�5���W�(w���8h!�L�#�:ܹ�-���9����D{���B�WA���h�h�%��x����5�x�\Q��s��֪I��Ǳ����AR(&�������r��.�w8u�I�Ien�"� v�4��L�+ $Ot�0�������u�-uuP�S��[����8�8j�r d�� �	�c�R���Ec���i�;D�=����h�ݏ�V{3���Y��]//����6U�'h%�;;�	|�6RV�I1����o�>�M��Vu�����l��by���~�\I4����p���#ذ�@$x�8q�?Ҟa��}a�9��l����B<�ԩ%�m��\:�l��X��M�ȑ���IuUcJ�9Ҩ~Re��{��fY� X	g�����o�g���G="�6�5�r"�֥�{�"G4C���`n��x��DƔ�{�QA�����as�����eU�o�1��c�AI�u��~R����\֬y@��<�A�ш�
M���M;�D�xg�z�ɝq�R�y�b��w�-rgλ��l��T�Wɉ���-�-�ϲ,�q��Vf���X�Am�ڷjɕ����4�7�5��G��@�ߖ:a���kSR<C-�V2�y�5F�A���0�g�{�r�������'�� W���gG	--K(�}�����#���+9��=��4<� 1F����دُ�P�WȃHe�%����c�t�Ro���Ǯ0�]K��j�0/@��{��=�4�(]�蜻��N*��aUˑ�7̱�� ���oT���2��T�?aw����?3���G:� |V0~DS�ދ]�x�9���4���}$b��`�p�D��������rw����͗�R&�B�͸�m��U�kcN�0�j�A���=��hX�D���`o�]�02X�:f8d���9���!���P�${Y�k��MY��KL�Q50`P�xEo]�!�t��2���5�dUɚ�Zƴ��:��[%�$#{�� ���v�ԓ
����N*�꽂���Q:fu{Ӟτ[��mv�
ϰd|�3�m7'���×IA��e�&�"1_���7T��h��}�0D�F-�P1�kf7(���՛��;����3��%˲*-a �Kp }��pRӼH�G?A��b�gcX���P�W�ɓy:@rX��L������[�B���Sr&=�����P��^�?%�l�1���B��ۂ]��X�|���_N���'<u�Yף7_��, �9��Sn�`�TIy>S+g�'r�"�pOG)�C�i�o���3\Z�~��n�T�K���`68�A U3� �H#��/8�\%
{��c)B	P�����qr\�ޱ��_U������'��'՜$���R�t4�_ �p���Վ��8J�f�p�8��NZ���s>u8eH^XРg3
���cz7����7��u8�۶�[��.W��awWl�M� �}�CGYֆX�R�q\�$��3���[�= ����v��a帛^���G��\������rv�]�j1o>=(��gpg�C�нr��E�~�i��7��`�g�|a����]��z2� ��X��I+�
=��DF��.7@z�n���ZL�[�R�_\ݷĥ�~?ɺf���#�YU���U��4�6�~'lg:��ؓs�Ɋ�W�S��}/4�7(',�\�+��3��(n����^�VNq����X��e���M�!��Bc�"�1)�J @�w�����2}7�ѥ4<�f�݅�4�bYm=C�#ϗ�97o>]���OƮMcϟ��ăWwt=�Z�� `��,H4:�jC�&��V0� �M%ĝ�� �R��Ӣ�^Z8P���S�clY�-f2�r�w �W���1�����y����qɈ�+�Q��m�ۧ7���7��gƶ��td��*kJ�`�Xl�	r���$h��p쮠�C���gE*������𴼑�F��l��ؚ�I���5��b�j(�8���-2b���0�i#�0w �r��-y��X�#�i�!��]��ߚ�[���@�g��_]��֪�C#����a1�^[��,H���	#���F�ѽ��a�n۲$�B��<k[�pv2�Z����g$�EH!�����D��=AxM��jaWDxf��}���hkؖg��x��څ�)$h0΀��l���~L�Ep{�4jM��5F��4�%v�}�L�O΃�]/�K~"t�;+�ݓ�[GV�}�=�� ��q_h�.ڌ��{c��W7���N����J`aތ�h� ����of��BZ}���@w�	��d}�Px��6�� gLg�r�Ç4*�l���X^��CCt`'FH�M���<R�=�|�:A600���Ǜ��q�%�a��0SI�g)H�uu�M-�Ԋa#�<���zi#��A���@j��v�`Z1A|�B3��MƄ_��ư�_5�*b G���=�@s�����s�hj�|J�U�aO�L�*E�x45�H{��	��*��ؕC��2��P��CgAOEj�����bY%��hX.��9bJ�DY�T��iJ8�X&D�
�����]���tۑ��&���{ۡ��0D�?��[CW�fG)�к8{ ��+'O�����Bf5ܫ��>��4�e��3{�z9�{	t�7CA,� �m8-ȹ�'�t�df��?�=��^Бd�N���Ec���Lrz�aq-��;��y�$��+����A�h~���7ipn9��l1�.�<q*d4묲I��N=D!	����s!KF7��ǬoU��V�u��o��8�I�����A@A1i/K�G@1F����^������9�]�2�W��(�j�I,&3<��O~��z�Ȱ�k��$f�G��x�K=���"�IQ�.i!*�wG;v}(l�ס�3z�[��LQ���_�u��q��;)Կ�!o�Qv]s2������F^:�|��"6��[j�f)�w�f����	�T3dfc'+)���
W��2�ƥ�p�5N�	�k��n��j�l���=P1�z�!t{yttiu���7.���25����z
=b�QF�Ὗ�D����[H��`ӄ�hP<2&[�PN�zuh�������W�@�^J�̩������]yQV�8�s�긋�b7:�BI�P�C�ꊫ @�@l�?,��urn���&yhc�|���i�p�lf� ~�ob�B��Z��g$�ChMuޅU�!�b�=��G�s6�I8'q�Ɗ^��t���?C�N�Q�˄�;���Ah���C�b��'�s�z�d��ը�/z�܉�?w� ���pl����`8ؿQ�]7Wz��L���-�8�8���LoUT��J�1g�M�'_27B��9�p������"�G�1r�Z~�ఔ60r���H �a�6�t��5����NNIo�K4�Z�h�S?E�������L�`#�I�Ώ��r���t��J6n�F@L_R4�ۊ�Vm%��R^(���U� ��-|�B��X�u�@�ح+P%�i/�~�H��f������B�*q.��-hPx�)�����9�����B�����5׬X�k"�1�JȰ���U�%���D��
�ww�e�f9�{��Q��UW��|zw�[i�"Z�5���,�Wz�ВK�����^�1����(rS}`?j�o����p��Ð��2���Q�5�!�����nǬ��y�n��B��"ڶY�E�Uָ��g�@fȚ���p�b���`,��JdLv��y����~���dl(�P��@^�iLC+�H��D��,4����U�c�j�0@yi_����~\��s̼Q�|��BL��/��VJm��wkd>���>��	)�} �9 �j��qr0���(�D�u��XPA:�{���W�3�0�ӣ0����琲"Įh�l�̧�I���} ��"w
��F�e篣.*Qg4T�+����X1����j�;�!�����f�q���%s��ʐQª���]��/����^�8{��fvI9�/�)��qJz�%q	T[
�D`�v�1vu��,�N|/����k�7�㏰����wʺʠOA��N197T��T��j��k	�v/����V��&�|+b�N�����MO����r��t��&N�������X��yލ�[�L$��P�e���F��ioU����p)��+u�{Q��`~X�#O���]m_x�[}��= >�Wv&@f�O�Fg�H�L����7����t�l���,ą��O�5ݝ�M9%Н�?�[�=�Ąb$Gh �U(8��)�5NLʿu�s���A�O0�����v�.f�U9V>�%�U36���D�!b0%k>QPH]�˃����?�d.�剎[��# {x�@R�������6x������氭�a����aR��~dיheq�opE������>�@���κ�����w�
���O� Z��k�����?����:�f�`å�.��	�)���h��$C'�C�Za[�]̑T�R���!ǻ+#��g�ا��S�=�0W�l����Crj���t������.��%�+��#��f܍A�6;�K{5F/U�%2(C�3�����Z�!���\���c3 U� ��?��40v����&&�)��5X��nX�%��Z��|�^��[kc���JB!��+�^ƚ�t*l���K�C\�ƺ�0���s��z�q�������BVY�ȶ��4���*�t�B�8r����zD��.��dLDPQ oN�lh���N ]��A�I7�Sc�5Ȗ�@��nxP���ۦS?ښ>P�A+����^p�ʆ��߀��A����J��.N�H
=��@�(	�HǔJ`��:�6�)�����b��l ��i�?6��-f\�e,2��c<oF�k�����]j��U>���o� ���Q`�E0�XP�[�ot<��#�usqQi�-6b�Wv�Nt����p�x��`�T%cu2����-p�ɔ\^^B�-�8���v��V��)ڰ6�(̦/�b�;Ƥ���"���ɻ\O�EG�m#���A�����&�ڞm����Z�5�>���敹�!\$��E}��DП�>��.�٠��-�`a���M��no����q�@��[����D�� Qa�G��p_9~l&S���kM��>��gO���G�^�JM�/�����x�B�hی�j�ICi���z�s�I��0���K�YըG���d��i�r���2�w8~�x��oY5�@
�{��a�k��4{I������0�|�T/CRrh;�(ޓ�JU�d�(4�j�����!>����j$	�dX�O�����+<dӹ���V�V�0�a�gp7@�h�O�6�>��TK8iM����2A3�t]��6^��<h��[�T@&��:ߠ�q�A�@F���,`��4�ǄPTB�/9b"=f�Xv,�'��eu#;�b�=�t����a��	�ł	ǣb�U}^�ۘ�w�0����,��ڂ��	9<,�&Ճ�Ylh��6[}z-�����z�$7l���a1m���Q��yVvڞ&��Ut�[Z�����7=��y!�jr����$��h!�r]AP����;����!���� ��/s�8��RtL�����sj�Xշf3�Ł� _�3[��M�%qJI��@���I�C���!F���B�k�݁�V��(�Z�6�:���]��ձ5�ʛ��QX��V0	��q�7�O"�KĪ������((�	3'-���3T7m{�-D�@�g(����H4�H���6��ܦD�U4 �Ô�E��=V~t5��R_+��ʏ��ER2�G���,F�akh��Z����Y�v3�`�w����?�&3+mV����ь���2����v��O� tR2��G����/�����j�i��7)ȯ%ձ>�;	A]`K8�5�]W]�S�7�R�XdZR� �S��n��)�;ʚ*�H����KO�	m���\�o���5�|���c�J�nt	o����O�%�7�JV�X)E�׊�砝����&��i�Uݜ����)ͲHƲ��F(l���-zRE�B��T>͉��Me\�\U�T|������'�3����C�(%��q�Ļz��y�1t�bI�<Ԅ7ѵߐ� <����E�{#��fo:�'�H�㦋U���jo�,��|)��_���U#�W4^׏�rS�$|@�|I�/��R�]'��+B^\�-6 ����-n�1��YK&��GǼ�j�Yyhi���[���k���#�j��&��� t�"�Y�S���R�	ݓ@V��싚 <Ǧ?{f{6�IR)����Up��}'��:�� @��hmQ���8�~�߀����xo����X:���ݭ(���a�,;�l��%���Gn���+����`�������vTV�AOn9K��q�C��Ȓ�jWzά��+�s`�z	�L΄d�㦪�����80^L���m��]*ԋ�C��F�������v^,W��7�ߡ8�����j�םù}�� ��"AW����@�n��󪏻��\�@Gs����"����E�a/�*�:��Ф�v�u�9�I9�{��(��j/ҁ�o�1׈ܺE~۾S���}�m<�m/�iF����B�z���}'�v�`�ZA�Cyi�E�����v�5���73O�Y�Q����/=D{Q�Z��N��R��m}��-���
7��K'+I��6�,@����ic�en��g#�Uc��~�����@cy�x����W��2�C���il���o�A�������֧oj�b,��ms���F{�Df��b2��E�W�t��\�~+��j֝�t�zpo�)PY5Y�=��/�
Y>�,�S��x��q��YD����|:�g��O��c��Л�}�慉~��#}���9_�*��[��2֗Q<E�|7�u���$�@z�%"/>�>` c��B�àV�`X�VQ�����:M�p۶#�GpQ�n����Ei{�N��\q��KZ.M7b~��@�W6͋�p�b���(4�H���;_\ƀ�&�㢦}([+u]𠀡�dbN�T�6?��.�m���@86�^�/{��T'��6�O3�t>��������@����t��漶��{���2�W?��M`�B������aX�������"���y˻2���6���G�+3�ϖ�?�ch�e�M��%����_�F��S��*�	��h�`V��kƙC����Q'�ܳ���Y�.l�vYb3�b0�f_�'�^��j_�%��j19�B&�'��ѱ�vO��u/��7������L� 	�����u%Ȥf�Y��d��TK�Ϊ��X���4Æ��󨙸Zx���I�}�o���+8�u��5��J�@�#�Y�T�������+�sD��!~�C��wd�JȰD?��(���'��4�����_����!>Pf�D$��vE_�ʨ<�6x�5�"^���K
�'�pY}��F; B&�w�:��)�;=�u�U>ɑؑO�XQ![�#�
�B�)L�f;�=rh3�:�k�hY�����]D�`��9���T��I�5P�s�FQa.s��=���6[�;-B����P�������d+��:�iTE�����"&��#usܣ��=�zx��U	Y�nj��̍w��4Y��OZ�z-dR��/�r ���o�� z�,�̤L�{PL���E�����$�N�N���3_*3_��	�`�0z��z{�����锳������;��޽�ݝw	Ni�R�(]��`jdHϱ{k��Y��E�	#��Fl/m�7�`5�P��b��������qr����0�����D����+���� }�:����y�37&�+0i%~LY�@�q���� �޼�e�!��vb�V��������U�Y���nĘ�8���k�0?��P�[��
rY���k�H�E�H�-�3.��EY�����(�M%,�y"�ԣ�p�E%�9�}(�6�&-�mb�1��8lG"K�d�gg�>��:.w�GN2u=�@5�X\���l�Ck�,�AE<uPC�n[�<���!ʪ( �k3��*Sv�F�־6vۇ[Eą�Nk�'���=o�f��f�b���sG�
���݊�|����n�?E*�Y�� �FV(c�;�Ӳv	!%��z]�����I[��Bϓ����1Wbs����mxzmo��!��P`�U$����݂��M5{V��
��> �'�C�c�K�7˵�L[���=ߧ>ypTˬ���;-��A�����l{����M�C7Of��)I�F� ����8�K�6�z�d<&�U��u���2�T�Lft;���W��G8?�<����'/���X6�%�󅷖��g<����k�[���U��h �`01��m���V��C���߾�+t�����˪sT��y�~�Ӝ�,�����i���v��ЫO�:�|�a�iPT~>��b����	��������%��}l@+�~�e�l��㈱��D��dz��@[K�*�`����EN�(b+��3T@�?~)v�7�f)R�/4�'`H?=N!ʦ+���x���]P|�f�������ᘙ[�_yu�__6m�Eei�}ķ�><=q$�w�*uǶb��8��Cfa+�+��GK�zlxm,O> ')�J��L���.�.�/�ɗpyZ�b(?]�R,N�%�K	<v�c�no���(��p�Jg�-?iv,wJ�IFZ0��]!c��m���q�h��@)S���҂ESˍ[l�ڼ"y��\4�ȢOL��Fe�e���̚'c����� �Ʀ\:C��OK���J�q��{LO����2���A��jVt�n�,")-,����U0b��`��n��k-5�g�@�&+�V�������:B.���1�����&��3�	L��IR�Iky �]%r�9�HNyr��:�[�j�x0���N�U�Ɉt��7|l�o�y:��
	xMq^��=�<��1C/2�|�ذ�w]5�\�<�r��J�&zPK�z�01��+x�!D�A,��7�]���Y��[���,j�[�[��J:t[/H��/T��/|Q�Qć9hW���P�XTtnY�X@��o��v���-�
B���{u��z��8��%����@�
r��q�q�5fX�����Ki�C��)[�])NY��*E蒛�qZ�O�X���.�@�&=:v��S`N�jb,6s�KҪŔ
ho؅d���`��H�����C��D�}���僥0;�����o�F�@j�RB����7��nҭ2��`c�!\/��[�;������ێ6;���$6dOuɕ����N�y�4q;��<Ona��,EN�9s�x,L����=yPI��z�41�.�+ u�5y�����"S$�au�y�P�x�Fa�;0i![�S�-h\9�Ap s���dR����P�6�	E��E�b��;��\�qa]�a�J3��}�ٝ@�Q�7�l�,"��|"�(uF�Ϲ��ιK(��}N>����M�E��K7]���b������:X���$3��y�@Ұ �3�V����c�����γJC,h�;�ݥ?|���aG�Cp>��L3�'��O���x����*��#��+�Y�����Ve�]Q
���A�5���-���WT��ƙ�H0p�, �v]ڌ��r�}��I�p.�����e6ি2S
�<�ha&)�
���dQ`�ٿ�vԩʸ�|Uy�E��.���E<h�ƩA��m;���ۋ��r�׌��۹��Ҿ�}$�&��oIȞ�7C�X+-��A������r�G�E��k��ǋx��-Z7�a����|#���@������`����P��w���r�Ѩ,,�U�~������ׁ�so��)��N��7r�Y-�졽5�p�q�2�o�\h�[+hsAN��ߐ���Yt���H�հ�AB<����p��+��={������;�pno���^59G3� Rc�A��hk�i�1vE�&�޿�wo�,D��{r�Y���}^�J���Yt���v�H��Qކ�s�F���rI����P�j��J_i�*���2.2<�\Y���iXn-�j�s�fg��M��e�t�G�J�M4�p�Xd�@�nt���?�����1-����X���F )��b�Ƈ�$} ���h`��*�ɸ)�l�]���@����[�77��;T�L9ZG��^��
�|�&j���tV"��Ժ�����n��n�ީ®]�v*{/3"�	V���<b�(=;�+�퉩R���Bސk�$���9�`��A.|�p֛���K׏�t��R�'�k�˦t�l�Mn`5^/�������,�x�ͮ�A"jM �!���p�βƕ�V�Z�JJh@gB�9�#Emu�[�(�S����g[���(�n�6�¤�ɲA;Y�0�R���G����ro�h�!��ֹ� �el�5��)��@CLʡ�g�|�w�S���!����|�HA��p�X���*���I�0���g�z�_oC���U�^<MXO��Ф���ښǔ�ƴ5��т�Bk��8X8ꎢ5��i2�����(@���K��ap�'~���J)�����ĻX}��K{���S�F�q-m�8+�T�1�
����잎p��`#		Z��S�KY�ܗn����P�C�[T���Z�@h�T-��u�[���<�]2z���1���2H��(�!0d�m<���fr�*=��0��\���ˇ�cX7���]��q��Ll@���,�V����JV�w<(/�v���L�ժ���D�����5��w7�&=ӢNg���	nA�|��8%0�� a4!�wĔ�;l���Q� ;�?2���(bfnz��w��䡪[-�@G���ӝ�V����Zm���f���zQ�wd� �<�e��,�\|񆦮� ��2��Ji{3��%�sxA��yR�������q=�Om��3͵��'����0�ʾ�5 ���;w��0��Q���?��(����\�yI����%��B��N����	���7h�.��Y4`��~ "�1�tOJ�#6�H�.P(m5ֹJ"�`�ī�_�󇔲 ��j�~�����R�A>�M����_���k֬OU��[���x�W��.��Up��L�~x�� �łG�R4΂�F	�^�;0*�.x��G귴4�VL�A9�ܰ��*~L�w������6Y-p��ߪ�������9rv
�t�U��( A���K�M%�D;�Ҍ��i��v���w�TgI��Z��5�gz��e�`�0��oC8:�*�F��OP���wwl,<V�>ȭT~V%xe7sF���B�ĕ,Ky��a�$�w�\�|���cv��-�{�P	S��"P�E���)�z`�/�O�#P��L/+!<@p���"|ѓ��i���5S;�j/��đ"�=�QUr�)ϳ6��qA]��6S�?�]�
���mJl^P���������NCl4O�%\3�o%<?�9���Ŏ
��2'��5����մ����ރ��P�c�)u������@g�m�S�M!�è"���@θ�^�_�6ԛ6����?�<��l'����><y>�`
`k�>ğ��W���U�M,����²�PH	I��-mNx�7s��V�et��b?K�(��7n�pU��eoK0>)E�q��q���`W�����LrV�R�*p�T&��E��	�c�ة�[����o�W	Ba:I�z�r��͑�g�ғ�� �Y(�|������6�0�U&��~'[���$��\�xE��zj-7�����>�(z/~%� P�+�ͤ�_��P����B��'�ǚ�O�4���T��e�c5�(�w��.���Ԫ�a^��P'�ƫ^�i��w����`iv��'-�?�G���wm#y'Wm��ɦ<<L��M���yX���!�߯#��� N`IY�J����K	5�7��1���țWg�@�x�|
%��j"�?�M����v\25c��jm4����\QX9�G�`��� m��
����k'��;f�A�͋��|�~�SD�<)X䠘=��x�����?���Q�8�ğ[߱j��C*}�xBT�Sҕ\6

.�tp�p?��G�<����Ex����f8�Yk�N�B�����#���.�}qZfs2[{���V�����d��l�Ι��d�˘�w���i��?=�!O���ꂋ�Հ�O�v������x:TN-���)��b��� n��O�,@�B*�H��$?�� �~�|XV���I�p����6�2�r�Y#;��KD[fTv_j���O�OR�Mr�%�m&��
$H��l�2<�-�|�ň4Q��FǏ�����*R�$p7���B:���>S�eM��*�@&Bo�VM;5]A��V����M_N�7G�9H�r:x]�R�3�d\�'hB<�|jtW���N��]a�U����kĢ�L�u@��~��k#l�zN)kɼIa�y� $~(׻�S8�y�<<C�jjI�c��k+}�7ױw�
we%}E�����p��֦�J���On`c�Q�J>V�b	��#�&e����|غM�2K��G�	��m�qi�&O,���O���2]Qh#�ݍI�����îq�9͖�¨��t�N�qH��-C㩔/F���R[
rg�(YN�y>�f�}H,��΍-!���v���2�'?�1D^���z,�h�b�rdHA�t� AQ�K���8�51НM�,�����L�P*ok�(����U�a��ue#�O��ip�SP1�%Y<e.�L>�'��>k�))�����ӯ۰�w�`2#}�@P�)�oV��S���0xw	��4-�7<U���w<[�Y1�I�j���n�Eo��s������<+,��슋��uTp�X�#$[f� e��m�Z:���Ԇ��0|ᙬ>gvJ���6�s�<	�'�b&��o������Ug���8i�gĶ�݋�xWH�!VkA/��	���9�X��DƵ½a 	A[�H֖�0�ϑ�����I�ʷ��Ǳ~�(�I����R��_��X��o2R���/���������h�3�.�ٻ9�枢[�~Nx@'���W��!m��E^ݴS�/�:��U��U���J�#������C1�8y���l�����H���0�@�#���A'�(T��G��+�A�'���T�E	�c��=pvFZ����9^�dw=��%rF=�${s"�֥���67"9���cޡ��ɹ9���6E�ǻ��k8O�f�vQVeJ���+���{4D���4Kb��>�}���5_z3%~&�#5q���;�-]g�n�'�����OG�2o�Ϥ�񒷪0�VXo���fi/���)�HI�42 1�1�*:��ϥ!��`�3N��M���9h\cO�����ϝ����?��Z��׵�3*�b�F��tzCm��Iú�p�6P���I�O9e��\?��1(�N 7$�X��Q���4�Ť���v1��)~y�J�T��UkwS+ӟ��_xS�޸�˟�+���h"O�:�)*�����u��	J���֑;�_�p���������J~�V��r�YL���-��sbG��崸�.?D�acK���-�p'{��	ҳ?Y���͖����Eu��C%%��&?GP��M�sߕ=4�}C�Ϯ(; ��Y�r~��YlQ�R=/����ȑ=t�p�P�>��aP�ae�֒��Z��|�1�o}M����1�g$D�Cƥ�8�f�f���*Zo���Z����}������d�e��rz��#{�>%*����Z�ʕ�Cf�e:�v"骬nw�`Bjls]�R�ro�Z/��@.%�ƥM����z�ȋ���~�f�8��܅R���iy�Y���e�1�h7��%s�r�*�$0�~� �:N����i�눺G��([�������HQ�G�j�9n�P,�L
� T<�3����0��������I�w,H�i��o���?�v��\U��ž�(�]vr��z]���C�y��h�(1�K���iew7JK.hK�)g�d(�Nb�+����x;:&�Nl.V�=[�H�.OǨk�5�z]��-Zڳ��_��
"�FW{���w��o���/$�zT�>�ꈍ�=p�U�\ r2��B]K��A0L2�K�lj�@7[-�s���8۔�{�D1�ج٠\��H������0�-�C^��T�!�g8�e��9�*Q�_��g1x��$5���"��Rˆs�_1��=?�j�T�ϚT�"�^�gIn��uݷ�xZ4?{�A�O��r�~��z@��������{�*�h����X�'���y_#����T�	�T��p��Gx%I�A&�#�K`'��.�Lwqc�i�����{j����*�L��O���d�6\7ќ�2�L�)uO�Ga����H^��������A<Sv{���v����`�ף�I)��E����`Ū���J�޳s5_3~��B��x7~�a(�OG��)qf4����o	�v�4ZL@R�Kn���ѳ��A����-y�d6�Zy�׉h���C��(�H|�!N���Tza��������ʷ����Z�e�'S�N}?9X<^(;b@�����+7ctɫ:gF���Okp���2�˥U�=V�0���I��6���������?o����y�u�ǩF�Y�h���c��y�у��C���O�Jp~����ēJ��i�&ΫĈ�SL��qF����MR򻳸j6α����������5�)��6��n���M�9�s���V��L�v���o���͠�:�}�kَ���&�0��GW�.܄*��^u���5T�D¨��=S�@�������6d��!%v�s���]K�$�ׄ������|�<;�\�^�2S�2o��.��C~J�Cz��į�J/�����2@.R�5���h�H*�aZ�3D��I��"�Ӟ�'�ѫ欣�Y�����R�
��{M.K:��Qy�W֗<��g���'L��p�j�eL}��b�V���gq�́hA�����:R#�vY�B��%�Q�wD\TA�����c��*P�P˦��3�m4p�Cs�� �Hh&�]�T��m��M.��Ա���->�6�@Ȱ@oX��mx��׺zT��w���GmS���G"x� kV؄7i�(:z��P��q���ŏ���(׎
c2�W�n3��'�xK���M^A�ۇ�Pa����aQ����c*'������w�Ȅ�iH����a���m��6x�;�#��O�0��u�?�XV�z�q@j��&�sD�j���3+\�cm.�O��X>�^�����l���T�3e:���0F�U��1�{w4x�)��x"Y!��ݛ�V����9DL:�p����IqB�P9L��u�ܡO�
�@��x?P�6����,(~���"�Ra�:����H}�q��A�:��DS��FD$����+�~�������>؛�uU�s�)� ��A��p
�'9���A ��&�C\��!�Hc�V�l�Ҷ�c{E�g�Q����8�*��z=�����D)���vp����h� ��j�C?Í��b������ׁ-{�2.�þ[��kP����Y�&}T�u ��/_�V<�`��.;V��K���z��"I/ K�~|���ZW�Vd7�'�G���G�C�f�ɖ����G��hk�	�<�m+��(o�����<�b)����r<��:I��ר[zL���Xyk���W�x������'��!�,$�1��-k�sXg*^�a8�2�o���+PޓA��t�ڝ�m��0��59�K��5������x�]z�gv<�})�O}㤀��9�ƚTp6�XM��w��Ywl��`�.`
�W�M���|�'I9�8��~�Ve,Wn		3���x[���4�.C�V�=�<��њ˖�Ax��/��)O�	VM��%<�N���}%�nW�@��D1��缩��e��
{ٟ�i��R?(�1�b*\]�������~����t����Z�R^����f�u�R��y,*�`�1#�Tm����\N�����	����6XNmݢuS|��zE����^����a�l�f@m�d���%�8+5�s�
I1K�������C�ȽG��Sd�l`��U�u���b��F(���y�֒A8:)-�A��s����NU�}�W�/)p��_�3����#7���H@����/[�f22D�d�a��Vz �I9w�L����+��s�:
ƍ@�E�_Ûq S�Qi��8�׺��B��,��n�&�����ۈz�����[W�?�VE�~9���s
��VL���r9�����V�p��.�f+)a�;!9D�Uԑ��J�m�Q_G�ŏ
�fk�c��I����������y:^�ڔд@l|LD�ߖ�S�o0P�M*̹/���P�j$����А�_����$$��p&l��9_J�Fv�i|���B��T����s�C�.+~ںH[�V��S�ZB�5e�!�����Ž+����H/�ؤ����P3�ۋ���+���b,��%�mz�a%���������6$
��uY^_�5I�M'�X�<"�?��t�d>�D	뵻��R��3�lN�{���Nɗ���:<]�}D�sR�ۙ�d�J�B�f՗7�̊���;Z⻰�V��W��ZZĞ��i�Ў��1�Ɇ�"�H���"�j$�[�G�E4���L� +koN�?��y�8�&�~�����7J�E�����`�f�"���!@��a{w"�6�Q��+X���7�
�Ϸ�M`4j�U���h�4��Ly��Fm���p����%�I�����qb�R�� bX�fmy���3�
;�8豞��V�d�X�Z02���k���B�Ϣ])�6���W�r�����6�RGG=����D<�Òa}!�d`�:J,�\�P̹)=;\"���(�A˒�@���3�a��
��E&6�,z�
���G�=N��A���:��=�D�������`�dH�@��%�tK��l�ۙ t+?d��ħ��+��S��~h���#��V�
�9���X�dWCn"�⎍������z���8h"ؠ=MJk���'ʀ��f���	��i��K�F���g����t]e�w�h^	�b�-���,���g�d3q�wY�I7X3 ?Yx�����H�fH6���TJ*��<?�H��żTmڤњ��>����!3��i[���Ƨ�'Eo..M2��5k�ѡ�Y;P%
�w~���O���� ~ge�Q?��3����h�$tk�@�9%�O6۸�i�	4��JP���CYW�z��Ʌ/V���q�ɔ��9�Ä ��D�}�0���"b���ȣ�-O�B0�?{�#Q��t�4�'AO]���ؓ:�;�����tܺ�?��� �G�U�&Ȧ^ڻ�����+��� a��J�ÑU�d|��0!d�=e���|u���ǂLr�����^��\����<�+|
<��)�R���0��M�yYV���-������%3�J�(�C
�p�_��c�K���&2N}}k�fC}>���G�BcT���ޒu�9}Z�%���|AJz!�)�k�r� ��*���M ��y�딑��ݞ!a��,x��'����$ry��(=q�|#e����-�]�H/N���?T9b��̕m�������p
h��<"�7jY�&�*)Y���闉o��qݦ����Zr����Av���$�ʂ-걖_�5U8��p�"����|u�).�?���F�l�U��!5L�O���Y�7����z�p��@P����������#XT2��~��u�EQ�1�CB��^�2��o���v={��ߔR����$�^�jiJ���Ό�Ȳ+�8c����Q-.�쒈^>n_n<��93�ʫ=I���I&l0+M�f��.��.�ȗ���]���t0�5����Y3T	_��Q@'̒R�_�ĝ��.fH�K�{�UC�Ҡ��
m��ڽrn;��[a;�E��F�jM��^7�JMN���!��H�zo�[��L4z�6Z����ƅ$4~1��Rċ��:]}w%P����ޱ�v���A�� l�ʒRâ]b��0�
=tp�l���o�n/!mBU�`s�&�l	�p�	W�9�!|�3fۀ�0�&������J��7tڪ+,�7�B/B��њ.O%Y�@���y�J����ME"!ɬ���S�
��ⷪ���Z�ؖ ���'����a���O���0���z(�i��jce����"(Yݤ(�����Ga��u<X
��0��1��"!F�$��8[@�G����q�)���JG]�Xӥ��]���5X���S��R�Ue>�/<����2=���~,ޞb�p�K= ��&����v0�M5�*E��j����dV�`S��ل��h�̉U�d�u�X�$�pi`�&gk�_��}v�I��D�vAϹ6���%������_��W�ɀ���Ws錋���A�4��� ��s�M���hk��*�jm	ʾR����y���g��������_���{/KĬ�Gz�s8��k{�q�ٍ�2���=��TX��^*/?mt���Ö����L׼_�������|�fa]���dr��3��Th;v��ࡴ���
M6��"*h�%�/�
} �p \�-�	�h���\��͓h5"vИ<IC�[����/]��1;�%�Pm���ɵt�l��O��ѿ�k�34�^�.���pбj+� �(U�����]����
ڈ��ΥT,p{H�������	L�15i�dGG/�T�t	(ըfW��"���3<��D2a5q�	��a�ݻ���MIi�`�P���B���|���G$#��V���u9#��t���i�/������8���O���v* ���<�
�B�%_��Ya'e����;�m���߈��`��V��=��ٌ������d�G�����U�-뷲H�����h�3�.�w3G��:a5�ʙ`�Yj��^��a��?2dg@8�ތ�ߣ?��F�w��� O,�z'���0��0��oQ�[�a=S.h��|�� �A�Wbbq����R8��u8	�'�Ǟ���0f/c��P����K�η��Q���4Ri������Õ�O��PT4S����g:m9��YL��F���'�&Ӑ����0k��vqw8/ML3�mHr&��<���R�N�'p;��k?e�܂�f'���%��8��d�	��ҹ>�O�gr7b���4��R�r����q�%�36�T	������~ �C�ayb0�u����*��}}�f��.��/���y+��w�~l��j�(�'�I&����)�c��PJ}(�h ��_�{Cf8Q�tcZ"���T�)�(�c\�[����P��Q��{�v�H�'Ru �k�� ���.3%��K��2+����r���q��*�9ʙ5�E�F|��z�W7�����bzݡ�)�%G=�!���W��(�n���s>8�M���?8��UzA��uȨQ�ʑ�J �� �&c�^ۉ����.���1=��|��}��z�~
�����;�_��$s��]��xbSU9Rr�mt�V�Rm��`G���46�5�S�
t�߷���t}��f��Z�T�巢��`� ����'�'�"&x/_��9P ?��iq_�e�O؛k�3͎f��N�*O�@Ϩ�yt��ͯ�
� 7x���%DO�QJ�~*k3�o��w�n���ؔ/��-̀^Q)�B���4a��<�Ҥ=o|2���v���o��^Iɚ-p����'of"ymo��~��@�?c�S�B��ûk�w�R����#a#"%=��(��ׯG��
��B`Л0%[�d�z��`���A�79���Uo��$����0'+�Wn���y1!X�����d*$�Ҍ7(�[sr�M�¸���b�KRY�s��;_�G�>Xo"Y�"u�6�MkޥR��(;u?�X���I�a�����(��r�ƍp���d�����s:1��ap>W������ᳶ�:��v����~6ϳGkO쿛Uh����~�\�'�k��Eo{�۰[Z��o�-��D����;Ұ&ik9T	��W��_O�}��4���_�F���0��QF��GI<�d{/�둬�RQ�_���m��j�8�4e Y'3�L�	wTx�������/)�<��q�+ð��lx���$�&�P�Cǣ�Π0s��P$���!E�ړ��\)��$����W<e<�֜�G����R�1 E����r�/�I���օ"�!��2��t���"i�Q��2kk��9[�!�^`(�E��ӊ��
y�����L��|t��)'�O��C�9>Pܘvr6�`�/�+����NT����d�Dš�d#�掞]�� ��-�����W�ޅ(��/0ac�1p�L5y�F�$��|^ڐ�u�,}1�����:_<m���lOғ�YHr��Fc?dk�I3ߠ1����O7Q��m�M�퐎��|@h�t�.~L���;���d�!p_-��C�Fu�/D�L�.� U���h&�^ow=���I~o�7�A����5�hc���;�������9P��n�:3Uv�VbUf��Ά��&�	t��s���H�����#K܂8�e���mOg/x%#�3Ӱ1dэob��qq��&�@���k�ҧӨ��a�ۭ�?t�U�i�<[ @�G|�F��`ܥD���˒��&A����o���#� ��`���9��C�­�F���}�NSV�����׺������i��y�	<ĸ5b���NJ>G�<�!��D��c8R�~en�P��;�!NY�l�N���9�(����	��)�ޓ�=�a󽱢��:8�Θ�¬�
`��Q#m]�5���	��ا\�c���Ea,j��c^�m&��@J����<�>~��}�!�+Qש��s�`ۢ��+�J=CH�����R��B��,��Y��E�D�!y����@�Q�K܄=tu�?#2�HK�ʊ ��Bom!6�/ox�h�΅��} �q�@v��8�Q��/��AIK淳l �Д�xI�#p����ӼG�unŬeaxت�l�׾[pal�'��m�['��=�}5�D��.P5z�-K8�L�Q����f�J��[����^Å}����d�;@2}��0�qz ���JB��G�J�O'��T	��0(|>��-�Y9��f���#��e�*Fcg�8�q�Ge���T\�.� �FC�$�����{��8�x��st��(�8�?3�����1C��268���C��u�F�A�3����RP�(J%{��]D�i��Y[3�������(ki��r�*�a�=���k�@�4�'4W�&�E����5D��]�7S���q��v����r���"����{e�r0��jC��ѩ���kX��S�\��ON+��]>s.���g�3��}<�Ib��h�J|,\X-��j�h��e���k��?,uYR��wL���%=�c�4�� �Y����i|K{?��k�I�_ǚ�gVH<j������jkS��QKj2�i�g���Y�s� �*�M_�"�j�Q�;����AtmIH!����w�Tʖr��^�T)��(Sb�vK�]P=�2:%{?S��5piQj��~�r�v��ˎ����.��R]��ԅE	k��wr�_��G�DI���^��:)�8�����(C�Y+M����Vp��ź\Fr"xu���z�sq�!3�%� ����yrj~�+*�s0��M8/�m~�+5'B�,o!?O�/�>�	V�+B�V?�/���L��1�Y���?z
c��	�����Q0�>1�f^K�����tG�w�8��詿�>��.˚_��+�A���R$�h����>!��ׇ;i���s�<q�-�2Z��K(+��Rd��KyGl�����tTO����zm��v:RD0᭏�����E ���M�ʭ�+jmEH>�묠���i0��\��̤����IK���:�m�N�YCq�����,[�����I{�I8{�E��C5��-Fc�ݬ|�|��[�E	�:H�V�x<������+��,Ĝ�3��#ې�.��e�@�<����9�8ԗd�gP(C�Kb:$��Osar5����z��o&u��A4ƶ�vuS�a{��w�[�����q�F�9�:j���#&+�{�_1���,1�~q���V�g(<֛I���wR۟�2�?~Ѭ����U^���{�nv���1�k���_�I<ϪA�G�&R>���g�>M&�����pd /� zp�]�x���U6U#>��j��#��kEP<wN��J)bڄ!��22�[�@aC�k��A��*����r��BԢ��ȵ�u��:��*A+�l3u�جV`��_��>�l�rs� Y)�Ge��ptD��}��u'��&��c�sY~;�#H�Ӹ��|���C��[M.��ȡ'��^
vT�4�2�-� ��2�;����Ř�P��7�Qzn���l@��$o1锪L	4T礅�1R8'lDwr����!�APl�3�B��� �ڧ��(�p&���`1�K�G�\{��%/Q��2l���[��|�So���QLU�� �l9 ����;�*2�-��W�`�n�C�b��ܸ,��%Sf��=�r�_��Xr6�(ܥ��w�Z��R���_�	F�rj ��c{��Y�SA���cۉE��Ǽ	=8E�[]�.�X�zKɡ�(K�	���$����bς�D��Ħ����b�i2Mp7|��a*|��,����/rD<�'��w���$�m&	�{h�ED�?Ƨ�����0D��n�K���3�m4�-�*����ภ��Ki����z �>�٦g����Q��S6���7��e��7��*2����x�p��N	ܸ��Y�:��՗Xzp ��[���݅�}���t����X��Q9�����)$�K�	r���+3�8�;����ybqT�f�y� ��G�ju���F=�Jd�P�ڹY�w[d�/�u�'��;�)Þ��A%n;�А_�$�3���Z��ե^�q��ne���@�*�C�;?ep�>��I*ç�J+���Lz��OO�|/�Q4��ˣ��6FjQ�� �P3;�
8v�]�s�z����M��#y�r\�c���#}��{��RqV�F�̌�V+Ch\mZ�S(3Z��0��D5�(vX��j�1��OH6� 6(OHZ���!�g�nVm6]�F��cn��Y��p��o�;�'v=�sZ�鴠���䣁Y��O�Z�/�M�6nQ,�`y�n�<��.+/�%�4T�7�8�isf��X���O�,�O4�/�����>��i�>$&~$�r\/}�4n�=Iz�s�f��:�qv/�pa��K�n\Xo������=�2K.V��d��.���H4 Y0~��E-���I� �VHݾ�` u�p?���`G��Е*���\U����D	�̀c�t��
��0�央mj���{{Ի��2l|����l|�M�t`��3�y�?X���tey�.�T��
��\ߓQ-�c�Z����=��.�"5�HHs��^�B}�u/�5є.�U�ꂷ5���'#�&��;�D��E=o//"�,�3:��_j�z
����$煴��re�Rl����x��3�c�cW%�1���|G^��}�Z���0m��[�B6��2}V�ؒJ�*�����NO��i����5>���r!���{m����[%H̛�	n��פ�{]�s��O�`��X�_7��7S;S�d��������R#uVr�~���x[A��꾩�u�Q�Z��"R{-H�T��_%0�ʞ���c!���E�X�ŗ��]5���F�θ[�?�����6��_�u�,8DqN;���bכq�W�@�B�Q<8��B��h[�qQ3
T���{�_E��9��j�@���H��hzC7U	|��ao50�U�i�a3�w8�$������)f]!�8og("��)a����r�c�yj�tEB�S���U��4-�� �ܨa�M�k��I�Zծ;<N��q�-�J���9k���Ī�u������[��f�C՜�I
��K�EX��T�D����t~��ING����v�3<(a��&KA[��ϭz!�*��f��F�1F�\a���u&[[Z?��v�h���,��j�%K,	�b.��|Q�	��<�O�-�7�
�I��G�b�!/}�r���*ݽm�������4�t f5C`�p�ῒ.z�2l+ȠӞFu���';����&?
���Dl����}˙�A��x��x�;"����&�1��v��|{���ǔBN�wպ�&�rVWu�KѤ�iˁM@�u�]���m��Md�~`ѿR��)� ��Gj� �:�@���j6���Ή Ҧ�	ɍ��) ���E̮|h��@�`�=�I\[������~f�Z��'�[�8l�f�FG�v%\��#��_�~3�V&�*op��պ�Ğ�O	[ ��h��tE�s����&�`�b�W&|�x��z���
�)D����������h�4êrV����ُɀ0;
�lH��[��`�d�Z[$�Q�#��H�9(-j]]��Á=�� �^|�k��u�Ik�n��o�L�\}ܔ<D���W���=�:]�UE��bB��W�������rK�t�����u�Dۄ,<h��Vt�N�����>,]tþv.>�ɑώ�|'�L�m�@��t���­VR�U-���61���;-��W�Bg	;&[���(���}�[����MU1�9��5x$�0�Ju6�L7��#DNh���>W��%�-v�\��o��P�K�S WCs����%b�V���S�2��н�'�Z��&R5�na/�C��`G�[��}�!M)�����Y�cM<܃��5�����tw�v�����\�柟�$���#��5u����'c�`�q�XYY�I"�
��<w8����EE��,�N�.f1�ꕁ���P�N�{g�!MLeJ�:�R�y>dW�7̡�e�m��1�+��F�o��cO�T��S�V[�'*d��V�1��R�n�����gU��[�a�r��LŨ�Q�I�@W�=xa��HE@%z�E��U��[z��ϖw(&n�
;�.%V��D�D.�lg�%����a~Z;�7B���H�4�bö̋ꠦ��eE�9ǃآl��cO���|V����_��^���	É�����A˶��� >��:��b�*�n�Pkf�8��)�F�X�{�'�Z�"�t�r`A��3�;�}W�EH���f�v�;+���@k���0݉H��0m~:�|���7<Vv��K�E��u����L4[8�lJ�-��6���KZ���d�x�L�᰹��v\,��]
�PLxá�HM�����&ܠ?>�2J�nw��٦�F�h%,�k�ҵv�X�lM��A��Eo`:�dsr��"R�b��V\N
&ӑ�#&t�_H8�^�d�0�<�"]٪ULc��a��X��l_X{&�W@�J�6��2�2�> ���NOK�o���2=��*��+�}�{GU�Ώ�[���iQ�h���@��Z�-m��I x��"�g	��(���m*ǡg�j?QJr�-kIq�?���m�,�?��Y�.�p��Cm� ����- �'�c�g�F:Ӏ�w0��0W(��d�����|
���#�D�x���,����:��dڱK���~K������j�P#{�w�������#T<H�4�������g@�L_.�����Q}�N�����p^�:�+��r�[�2��V�N�F�Z��S[g�q�M��$���'��ӻt��(�y�;�};��H�Xfn���r~�s��@ ;�n(f�0W�����ټRR?�M��yj9�JtE��(&�s�G���a4�'-��"ō`��I���x5�@��j�j��[W�*���1{�.CV�f�l`�<�J|:E�0�W�g���5m�Dڧ�Aخ����v�1�����T�3�^���*�����Q�t�����>�чL��l��pm@	Bb6�Y/���j����e��_(CU�2\��F�Wiύ[QM:��7�!�:VB���m�V�-�R����Y�:�kv�&ޭk)�6��Az���[��c!�:	k��'i��W�x�=v\E�m��O��	cy��s��m�xߥ��1w,U=FC�3��b����m��˞��`�x�X(�:]H��Ꮶ2�C�:Z�?����Xb�)��xaڂ���[�A*�eQ*:3��roK�Xh`�R�1��V\w�q��l��jD��w����q��!4*�`y�D�&&Pz_2�ｯ'��%D!��-ׁ�F����.>�#�D�=t+�q�}&��0*�����W�n��⇈XLi)[:J�� {<MA.-��d��<�Z�s��4y��.�M��P-���� �L|��$b��`I�5��'����!��;���g��F�� �F�c�a�I4�e�Lԁ]��2r�?E|tM�DJU���2����O{:OM��<��H.v��0��6`�����H��zͦ*%/HOL�PkϢ�OǽԗPIP�փ�v��࠹���o�B	��I�g#�Z'}w>'e���&(I�S�ے�ȿ?���WK ���S�Z�-���3���*jo�u`��
K��r��jq�
b��.�p�e�a`����wu����j����>��!"rds഼�|�@�N��;4�T��N��`����	R�ʬ�t.����^
ۋ��Kw�q�yv��<oփ�a�HR���ĞI$�6��$�|�6��u�a��B%�!�Gn!�#�)ԍϸd��cki`�*��_N�������Tu��$wM�~���=�e��b��c2����-Ie)�_�W��%~� ;�%_��k�HV��:����H�����/�m�xg��-M�T�`N�����9L�q�n����0�_��V�K��4�-&�^��ldd^�Agmt�#���B��N[&��`���FdmD�D�"��	���S��2"ν�\Оޜ'����Ts'U��q���ю 4媝j�hg�j�,�h�6?�"=�2D+�����E-��$� �g��&�j����J�ʸQ����sSD�:XCF_9�<+�=��X���o]� �ʉ~�FD"(�":?!����r�Ō�����h*,SPk��r��4p�=�|+s;cͬ9�0��g}+Y|��`��;ִ=��-�n/���R�$��Gs����-ĝ'	a�Y�h�-���`��&�,-RE(�AG��v�,1qJ���Ő ���/-hV�33Mh���*/R��V��E^���cBq��
��DϠ��dķ�@É��lT9	�o�!o84ժ,0�^�9�b����H�{)^����߃%�E�W就�z#��Z���L�<��Hv+��R�ޒ^�T����S[}�,���(��ǯ�cr6:�n�'n���C@���R4�I�j�p�8��7�`���^Y$�����0T�u��~��?[�B�($�nE ����A2^���'��T"�|r�c����|9�N��#J�?xH����9{�S�RXU��^
�(�	�^*����}�$�9��{�ϡ�8��LN�k퇏�4�]*;�X�6�f���ԛk`�z�����m%���3�O�	�cR�6բ���r���Qa���0�A�ҍ����U�tNaC�=��Y"@(9<�)!���������9����LtU/\kh����'O-���m�,hn��	]��۫�IM�ʭ/�#�	8�ݝ�ȃ^��"�K)��f�Q}M�l���s��V�E��T��.h��5�^xo�^-�2��\��eI�y�:(�i���l��J��튜��N{�-�'ZʝC�{F�TWG=:9�p\@�8�Q6[׾�@Ū"M���s6��P��ɢ>�N� ��j��ʖ AQ"�V�t�tt��dcC�,�$;�4�RA��E�8���$EL�ڥ��1��/�`'n���w']P����F�� �Ȣ�ZmJ����̓��@KWȗ��$�3qt�.5"�ɝ8�����\2��˭u��q�E�@�����ۥ	�Rȿ�*��8Q�i��4`�TU�oE��If2пZ�%��!b��k|W6#�G�Qh:�X�o�B?�<�yT�̝KA_�s�&𲄸�%ɐa����T��[�1��fl	�|9�����N5R�g}ɻk�p7��Hy�0��JmP�)v|�	E^c���UJU�J$d�=� ��c��h������S���K��W�1����᡺d\�n��NŐ�?<�+�=��$	�s�4l��'/�NX尨�=�	�T��@��n>O ���DԮ#;��;��4H$�Ws�.���)5gc_�I�����]$U�dK?$%PB��l�w-�t"�P������V^΅�����0�vBY4��3�[|�!�L�P���@O��I0&Y�V���LS�����ϓ���gk� �Ύ��vg�����MY���3���Äy��Š����pV�٭���������s@U�h.���+�/�����r��R�����h<�%���1�A�s��u� ����g]�\F��kd�Lq�Aہ�B�Z�o+����0�X�%�5U|L�ױ
8I��:�d�Q)�q�;挭���7�e�,��p���DZ��#sk=;��x���9�b���#!Pkܓ\h3�>�Xn��@�MK�q�'�C(�';t��4�g�K1���i��+�x����S���D�Δ�ڜ�j&D�֭ � �.Ci7}�g��A�y�͖<��>t���$2j�UQ�(~�Ig���eKM����}[!T�� H)y`l�u"�4���t���h,V�Lv෇?A��"Aa'Ō�|�Tk�Sh�6�����LY��@)���sl
����Jcr��q�
��TOm1׉�U)-k����vE���b2��0D�6���4�-�}(�Rq���V��"^��05=Z_��O���ǡ(���}3f�[�����ނ�]�sP��Q5e�oJ�p���}N��f!M�GBYר��ʷ�v����:��WN��ar]4�׹yʺN��ZB&��t%��܊Sn.4%6K����>�S�$y��s��w�$�͔�	�[�F�����H����Õqw��'��x�#����0׋V��R�.t�F��)���+� �˱�t��Q���W!8���6���͊y��7������- ��Ë'�Z?m"֑,����Q���ř�o7�l����4?>�2 �J�o�2(N��Ź�L��M�nVYK�|%(_yFP���eh�v�i��"��P��(�������l}��LM����b�$�D+B�͋��l������W�$�H�=��6|����p0I�p���Z�ߒ�Z��@�1�p�3bu�u5="g/�:K���С>�`U��KR�2��^��ֵގ�-%J'��Q��'��	&�g �f�L�%��G��E��Z,W1HG]�����R�dZ��`�E�����6���]�)k��8yλ�����b,�06���A�_:�����t<��6�Ce�/�4w{X��'��uY[_V��� �R[�(��M�$�Z�>���\���h�ճ�נ��-GM'`��i;��;�}�rᙢl�Ys���r̭e��{u�DtW� ߀�:�P� 0��oL]\�ǯ|�w��G�z�z8�s�܃�e������__./����G�d+��?�i:���_�%˜:��G1U��t�b9�͂Gg���r��c*��AYss�aV��R�'�w���)LB�G����I�;<'�Y��X7�� "�po��:���Ic��!�`�C��8�\����>A#��'�����K������'��4	\�F.M���P�+����#����p�U�(-�at�-(��O�G��P�r[8i�T�� ��e�r�B��s�p�V.Y�M��+HF	b^8\ک��=���S'YG���*��&^qn��\�O�[jp,�eK��|����=�0����J&�J�%�sQW��i�^�A�x3&8]��OE���m�W�6eK�"�ES�aں4D.)u�ss�e��n<���\�D���p�p���G7A�It"� !gFܢa��~7#�L���`�@�s�Bv�I���}���"������:�b���@_躝P�\��1S�n��in��¨8mZzbN�]�5�Y({�7��{�����[IGp���׏�E�7	Ȫ�vc�� |'$a,�����yf���W�tN+�� �~�l��2�^>c"��G�1�죫�����>�I���^0�@�5<n�Zt�/F�X֩�����9ʀ�Ky��	Q_$JZ�s�'Էk�D)(pz6]��M�"�1'�S����O���"Ӷ�h�i���5�R;�Xb�r�ǻJ�x����b���_����x1KP�M՝�+���J,y�q���8����:�9�����nd�J|ŉ׼0y�Q��sGSV���2��ԥ�D�Ë�ϣ��_K`��dFc
�ڭ�����WZ?�g[��Gp�B�[����3$���?O�ԍ*:W�`�N˟7��U ~����<Z5�P���
�+�����}Ԋ�F¾�&�w��M�:�mOK`@�5Gg��&�U�0�P�u_m����vC�:L����T����_KE�4�^F��� u���7�l�۫�*�c���l�m#�.y��ϗ$YQ�q��7� e���җ���`5^X��:S+�"�L��oW��-1�K߱�y
��~�g��M���2S+���E�iHv��X��,[����\l�D7|@��MZ�E���>�����@>����d/|��'C��	x�$x{�$|Cj�\LI�����ɞC@|����W���� ���`���J�Q��U�Y�Y������Up����6�Z�w�w�Vh��h��b�v�h�h����7��G���ߐF+������(6�r�j���7��T�p�	,�=�͢�Б��U��ڮ���ڡF��lzD�k���EO_ɔi���ٷb�� �%�T|�����ȜѶ�`^�]���o�g&�Q��| ��c�Fߌ���|>B�����=������o�p��ȝ���9J��&$�P�/h�Os�f��;d^��gvZ��H=�}��j)����J�Z�R��s�݀�.�N�,���r�ܨ?#�`�4�̱�N�%�d!a��q�7�*Ƶ��W�Д@\7Px��F�����@t+���h'݆؞`�f�k�����#���Y�E1+?�;$���[aB�h�v̷m���ϴ�G[ǙiI*^����p��U^bi[�{�.�h2. ��+?����찉;79��Y�5���-϶��0�z��އ�m7~~�i���4j8Qf�@x}�q� �Ά����d��/N�t2�����abݝ	��45	�e%�w޿b;�@D���x�"o����3U�
���7����5č�a�4[��.������N�`���n��u@a�q*����P����Z̏���/���j_2Z�b�mN�~�ѥ�� ��<->^�0R9H�$(TZ\&��b*�CÈ�0C���l�a�pQq�����N����=��j�V:ÝMTX��Z1���J��<~3CeF�$k#z�?fO�C�T���-N��T8�Y�LS&�z�jD6�kW��l�H�]�P$j�9=�����]�e���e�jDT����Q�*���-���?��-�q"�։d�h.��s�A��V�b@�����KA<ȻJ����^O�Tb���^���õ��Aos��5B|("e��s$\޷�R�n�������O4�!C�%R��Cڀ�ܳi6e�A�n<�: Y�ɌJRjB?s���7���^�jN��?j.ew�U���ґ��������˴�ޒE�~�G�T��x~<��(��uG�N9M})Bc��.�q�T�݈�ϫ�՚�xKr����5y�Pu�����+���CYs�S �f/[� �X��)���$�GN�S[bs�ʱ"v~/K!�&Çt��A`�K���b�!"���ڶ	!j���o*�h��~��'&C䠫�I .��	;>��7AF�� r��'OW_3��~���(S�^� %��W���?��E���߆B3R}|���/�
wQO�[���(P�#�*2 �?��y����\���_.��&Vp�"�q��[ )�ݚk��L�������k*�j�{��� ����Z��/�۞U/}��w�X���h� �}*�����0P�A��LB�L4�H�A�0���[g�����Y���\�k+��N��2V��Ȳa�v�����N�Q0W���z�B��՚to/���!|D8����%%�e�1���D1,H!�I��D�u�Uz]Q�n�����m��ѹ�^X��)e�m��[(�cR��5	��'����d`�\:RĪ/���g����B������b���+8�d�f(}�Le�h[������<���o�*���9\�WB�uB�i^N��}v���Z�Oį;S������,�I(���T��Qh�^�i�S����>���)4q0�(ׯ��Ɂ��9%�� �ƶ
�;'eU�$�p�2�9Ϣ�0?y%>����h�{��������$���m~v,�D�#�7��;��L�<���~��Ay\���S��@��8\�*���(�W��x�����u����,���S�R6���%�Pg�)Lɡҥ�/x/JE��-�W��s�K���j�"Ⱦߒ�L|�ja9����E�����xQ��`��)
��	�Լ�;�I�	�fh�귶�&U�L��V�|O��{�N�hXD�b��l������6T뙷ލ�^�}h1�8*���H�1M�}��3?��������f`�u29N'V�=�_ۇ�
l+�h�8�Ͱ$�C�+�`/V���:&�̢�#y?�,�:�=d�0����i6G��!�4ץeê�[����;e�Z���z�G�߆#(�'�%�?�� >z/�,�7w;_>Q�o���q�����C���0f�K'b0�>\V��oH��g60Y�w��۸��T&�&��݄�%�lMY7?��|.C0 qLU�}�@�0�(?�66��!��K2�]�n̬�\��6 t�w���)�H�0�Gj��b�e`�Za��Ks�.�磮���ň-����")��P���d�p��gJ+�/SJ%p&Fh������%SGT�>D�8S��G
,.��f�wGC'I�ч ��&+�`���z�ł@�S�����$�J��+k��jH�@�)���"�B�H��ݖ{�}*�H�Vc�O۽�BX��_�����Ʉ�R��ֆ�6�q�L��p9�~w{ll�t�L{�F����.��R@xw<T<�ֲV�g�Zr���+�A���U[����%��*X�Fa�v让u/���x'�Q 1����e�o,����F\`���ʞ�/�v�b����Xb�nS,�q�z+.`�-�Wm��/���B���7ʵ%��!��fG�� �a����oi;��|��p�3o�cc߷ړf���[�T�B�dd,}��Vr��0z+H��Rܼ�6"�����@�I�M�U���/7��&q ��c�֭W�$шR7Gk~�jFd;||7T ^{c�F~�FF>�͝��x��gT�.0_>_y�fT�)W1؍��Ǥs����2���p��x^��X�N 9F�q0/D�O��Wh�/B��NҊxA�l���%~���@+Q(/�EUs.)�8q�A��~ ��3�tJ	���ͫH�T�xC���[�jKϞ�b}�rGE���F*fN��{9�Ӵ�x��V�`��,^���&��X~��������	��4=Ph��Nn�.�Μ���`�',�*t&�-Hi�!��{��u���\���C�"YγKaW=��M��vq93�ìD�*�!�E��|�c�[J���4�kWS,
�K^^�XJ��ӏ���
E�]M�u�W���#7��j�B*��u�]'��B�4*e��''8�>RK�K ��̉��G���X��c�4.8��ig[�/yW�8���L-?�|N�1�P#eX9]l��"#%)C��\������˫��1^V����Y�4~��7�-�� �2��>;C��BOB� TVI����X���1Ds�i��0� 2sQ�ʚ2��p�Q��A�"�����C4�nT�ß�\[�����K=S�uA'#�Ӹ1�I��=oUo���廎:�(/�.���W���r�h�{dI��]Q	[ײ�kV�p��ƃ"]>����o,���M0e�	_�ȡ�!����M\V����]�N�#�b�M��$46�/|�2���{�Ѧ�����lL��?ƙ���׫ªt�O,�����)�gY#8eK�o4�}��<�?t�~�մWfo6���)R���m�)|K�m�k�e�!�:{6^6�)���O#lJΦ�.���a���|0��h~R�E8��}o���7ڞq����Ң0����pk��;F�+Y�_DL�4)IF��
a��Ov����{�5�[q�lG`!|�8S��(�ʏ���B�}n�3��m��@�b�6�`$N�ʇ��P�g�I�(����d�)��=����+d���H"��l�]��(4ç��n��	'Qy���W���@>�uo`����,j��.�P�)�J)>�B�!��߀�����{�h���g���>^��0]�&��qf���5��xѫ �CZ����{�i�!s��8��i�s���TlV�a�g�7e�o�j�0������Kо�=�)'<N�`��e�����iNv�<0�X��T��"��!2�mjԬ��E}@&r�	=J��RD���,x��Y�代���H�`��X 0���N.@?~��jЃ>r�w��¥#J$�@�� �� ,��-�_c]�?;G���v�$<�u��~ �l�T�@x-�j�:Q�X��ϵ��h��[�.L��a	N�B��jMN}��:��|���e?g/�^:l��s$B��{�m B| �̓�>��͉����|9��t��A��>M�fYxЦ-j�~��>xv�<T�A��bwW��#�4|�R.��1�L���AX{(���� �Ew����ܝM{&_�w��t�o���[/��G��lO!:���=���zM�x~��P�����$B��)�� (X�����_&Z��?���>�-����Лa��U���$��e'.���Ȑ�:bt(�sX��_~ȝB%���z�[�Ʋ��yM��#9D'P��h�]��L<���a#(�tǽ�k��������}�{$�F���E�K@bvT�؄����i!��Q�t�c��X�����3>g&ܩM��y��C��9�z^��þƝ��w�H���+�U����ó�R����/q�D4��o�4gH�m�JBVBʌ([r��h���
z���`�V�����T{-*r� �/�|����1�K�i��ۮ0���*Jl�8L�$�e��L^�I�,�6��=7\�|�]����H �ϕo5n�m���!��N�\���=�S2�3��iUIX:�Z~�g�E�]�D�Պ*�)�/O����zj�����H˯o$��<�錗�	�Q�!��a��S�n!M�����l��<��_h���f�8�Xф|�	�n{Q�n����@�=����gxb�e����f]
ξ;)I������� ʘ�q�'�6�>��k-�'�<�l��풮�.�v��}��� 3 6�Q���!<m9�iSEdFu/&]>U�6Z�B�3>��X�_�ƭ(�O�/�q<s��z�y=�u%Q�o����w?��/5�sN�P�[�o�G�${m
F4�=��<+!k�ﴪ���ۦ�}�^ze?v=фG뫀1��,{�h�fg��̇��D�g��BV��~���az����ش��z�X>>��՚�
��a�F�0_�؃M��Sl`�w�!��H1�O		�ꙁ�JWM�o�lH��_̉2���� ���W��lmم)����j�e���2��Iv�dR�@�:�S�&yl�<��HZ~�����M}L	t��.~f[�]�4��BQG8Y�!�ˌ�K��<��'���<h::��0�QAk�5
��CMج�
���!.)`�ླྀ�.�G��'~��\��>�4S��vC��1G��S�r�)�18�Ǿ����i�7x'o|�Ki`�{�4�c��%QQ����%3��W3nY�gɍuR��U/�H=��^���:IN�Q�a���Y͹��j�O���qLq�A��a��:"�d���H�bp�V˜�$�}ѹ�ɫ�s�z��D�d����ќ�#k�����C�/����7h�_�%��*U�?��^�.@�}Z���*��#C�"s���o��IA$�����\�?������P��HA�b�ΨIWtM1���Qz��(�4a�;���y߾�W��6�Y�N�� �TN��y����S�Z K��� k�	I�C��z�ۦ};t�lQ5O?�T��)�fi���)]�`d�x�5l��r�+�wk�,�c�
h��ш�w���(�}P�+Se�RU~_���~���r��F����r=���]�)aJ�a �[�5|�m�������2�c�6�3��
�r!to�VY�5.�&q�Kc'֠p=}g���=���o��Y��&��W��6Q����_C��Ӕ�X�g����'q,]�����.���p��x�vE�� ì���e�������%��W�� 	T���b|\a�ْ��)���Q'��TO���%Av�X��滊��7G�8����G��s�dI�ݞӑB���M����Ck� ���8ʡ���y_�G���®f�)X�/���&qѭ�����h�:��'5	V4����
��գŢMwU)��ꎀ�����M �+��6��.C��(ೱ~
ʗ�"gȏ�p67dz��I<~����r�V�&O솲��.`jj^|�[ՏR25�"�"��^D�Qt1�3Ҏ��M���i��]%��ӻm�}V��@��N��k� f�\����Ɩx�dh&����4U�J$��4�?�bk��\�8p������=/��܈?�Wx=sp�I�D��2S��AX��	/�MED8S����>�"��̹��-#��j�y�����3���H&,��oɂ b�L��aЃ	t{'P~i��3l�
�K��u��f���9sSI��ȭ�\]��%렃<�7+&�+�P�{6f��Llפ6y݅�B�I)����%�vL���V�Dg�B�e\�N�҅� 7�{a���������A���*�s�8�q���+o?�����H0<Q�SŸ^{j��,�h@��H<�gK_���Ə���'A��A�ëY:!��þz�WI
��FT;_���D���d���+S�
��}@ {��QV������n���:.}���ߔ�=���ޥ믶�W�r-kM8�``M\�M����vL���F�_� ��S�Tsڑ��Zн�_E��
%�}����R,x�[r��)�(���{�ՍMd�{�y�`�?�����Kl�w>��ـ:��0�Ӷ�p����z���\S�(�^u٬�]S�O��	fǂʶ�ـ �&@H>��T��挖~�e��3)�tn+��Q�Է�B��%9�����s��~�%oY��L�mi�A�R����H��`��F��S	�Mذn����B����32}ܭ���k��U��3O9�"x�:z�:��u�˱�l�E�9C]��3���p�Q��>}!�i6���@�%����%�G_�,?�o��W{=:��]7�dB�IF�����4 r5�����rge|�P1�m�p�\aUBwa�6�,�n�8�܏z�	�?@o��vP^��	��؈.��ut�Е��P,*�^��uCh{!Z��@V"��Uz�0�T�;�͏���0����9�Ӥ�A�A1e���²'��5�z"�����`n��z���q~"]��|�T��нaW���`
���`������%5 ]����4Wf�3�4e֍&��W�U?�Y׭���w8�4��@8.a��0K�Vz�B�o�ʛ�1Sf�g4j��G�n���Ё��ъު����¸01i��⺄ u4z�p��@)�O�9j^�g��dP%g ��[+��6�D�X��
�`hr����7�uT�^��Ƨ֥l�B��zN!�
�+4f�֮�z'����6G�
ä�BGa�Y �����D�. ��]�BnSɨt�9U�$M_a�	�V��0*Q��>�iH) �Л�5�_���M�f��J��O�.l�h.��0�CxY;�)�Լ���Zg�g��EC�]�pn�������=�
�d�����x����1�|�T��B�r��H���NG:ߘ�!��2����&XbZ* &UWB�ڱ��p��k�B=>����R��Y�"�wbH-��B�S�-9�(K�r�Xr-�X0��/Z�u�|�AƇ0;���ugdP���]�TOga�*���}�6n�K�@�d@>�1\1m6�~$C�g���$BiD��cA`_-h���:�ɽ�.a�
F�G�)��z�>J{�=�T�xw��+g� �pQ�,�\�_�	~_�:s�F$�H��^�K���K��$���"'~���Eݭ����{������]����?�wo�1�a1iYvI�s�K��k?��T|�4��(�ј�3�����N���Ҁz�.�p������:6�]�>�T��ӉQ���Z���)8@'�ݥM�xٵ���lH Ʊ9ڍ�jds��
 <"	z��e�fndW�H���'Q�W94p����[n\�[��k02�ȑ	73])��6�W��?n��[3�5���w�ι6��)�yG�d��6l�V�
�@�cƙnD7�z8S�,�R��xH��EN�,@��΃z�m���xDcD:�V]����#"��|pd=�Sk�t�[�a���@�8� 3_���΄�SB��T�a��Ӏ���Űj�I�.�!y���j�vJ�T}�{�w
�jy�������asF98�}(�^5�-��జ��d'c���Y'g�0q�"3�F�|*�̱z"�</���ͳ� u/5q����k�����W�H1��*���{���ŝ dѦ���2߭Ŷ�%�XӖ�}#����(�e�u��G]�3��h�)��A7~�������k�-��e'R?G��2���t��WT�պԧf���n����|��x}ުZ�bGw�R�~g�Fջ#����́m�s+���k�6�{k&��C��q�w���E�-#>.<�r,l��J#��<�$(��FX���:���c�I�!�@ݬ�?��$�K�ft����i����+�w���ѐ?ouQVq-�EHp�T{�C�&WM�?�ݹ|�|�R"��5�#A=��zHs����<�L��Ic�<uB^��HP��0՞���Y�c�A��"��M+�n�I�=���|�iЅ�N�R����O�ɺ�y��V*�	XnW�W��ѣ�aܬA5�n�����%���}�z�G	a�I�ըP���~\���Qm/���`��;��ʙ������J%�c~y�*�o�j=��r~Z���$��#�m��4�辬����ŭ�v���A��:��6�]��Z'g#9ޑ���F���C]^�l(0�4'���r����ҹ�ܕ�7f�'΢�0�(>���{�˥����S�7�řn��2c�Es�숝:����'*ss�<�6�"�@p#����`Y$���V��� U�^ĻV�T��\fmޏK;A�ƙ�gLc���x�EU�q�
G��q�4�����tʗ�/�{c��ц�����,�J���nD� �>��ϫ` �JE�Tu"_���#%���MKʷ�C���3�����9p���+��[h��.~Z�'i�L�Y�~>M	�↷>�yi�\��R��&o��C&����v'����	ZU�c{9'�7|�a���*Kb�;�r�̽w�QG�تRj����8����)7<рj�OQHd0�+��Y���63wař��9�h��*��u��,�N����MY�{g|������YJ�;b�#��X�E�������H�e�Y�t�/M[~�O(R�P��s@�M]�t0m\�θ�c�I+0�{�Z��8X�L�J�Srs�hÚ�~ޱ�����z�܄��[LfNY��xZS�y"���2&��pj&�"ڡu�^ʬ�(��;L?��������Θ�K��7��y	�ېM�Nك����Ӆ}������R�/ʁ�x��
��W��Q�8�1+���C���٩�E>������c���\��Kf�R(؄� ���]��鞶�ً?�� t+|����$[2��c܄�|JE��\�⇷��"�K1<筹r����EP�)ڟ��� 8{���+�T"�Z��w�WDS�6?e�5n$��&�?����^n]_%+r��F��m�&K�Z��T���&)�q��py-��SG�b���W���K��P{���1��8I�Xu��l���n�h��#��VfO���hX�_�GHJ%�"0����ȎAx�-�c��u�c�ڈ�w�w��>�5���+���|�U�Wf~;��Zr��_�@�N��yDY��Ь����a����kr�Ѧ"�S|�<�N-3��y��d�M.	,����iTz�o�������[ʒ�M�7����"���G�=M�գ��d�t�Y{�)1��F-�}����J�\^�c�Z��v�;@�1ƄeԪG>$,>�-�>=nV���2/zI�d�ʂK$;Վ�]�كtʯV���<̵ʃ�4�7I�4��u�Q��>;�9���o��h`w���&JMդgl�=��
m�y�����ؿ;�XP�0��aL��!����F
���E�i��	�q~����ǖ�����ra��u�^w>瞟�JR���t����6�M\`�W�T�X��!]�;Ÿ@\�bR�����\�,i�L�#е�6S㼝���<��py�ī���{�WQ�,��Ko�H��o�4�3 DmB��&�E�!1���ۜ�ڠL�}y������� �S�ۀ.	��3Cg��</z��-XPˇS[���!�?�KF�JA�=��~��ܦ$T����zi4�0`�Q��3�������K���sq��Z�@SX�=[��$�6�<7��.��LN~�r
>n&�ݰ��߬�bK����h�0I'u�u6��"e>sb�5��zC�Dpr�Bz������5����>�k�}�:��gL!ƪ�%;��U�`����0�4zW�U�4VI��}�LZ�L����F��V:RR���P��Mh�}:Y���b����c�K�'����3'0��J6:���
��㯖G ���v��fpTq62"ctg��c��b�١N���h� ��폢B�j�To��U�թl�t?Ƞ�-�(�[�-4��{��O�,�@Nb�^!�ɥ���Zi٭��˟w�m�͐%��?�(<��>Wxʤ�{�)`P���xiH�:ٽ,�gl�P
��_�E�Ez���d���!�*R��#����A.K�\�^0e_��]�~n���y�pu��s��x%t:�V�ƎW}��ϋ�C�h*��o{�4_��
�_���*^:�˦L��!�����A�Vg�~4g�
o��Z�:%7�0����\[�o��#��7c]��W�ud�]��q�P>�gk�~��u�~Hn&�u�����A0er nbG��U�o�F��b��[7�#�4�!	��v�NE�L��l���]n��;�8/��瑄}�-�&�^�"����Y�츅����r���(�Չ�BSoͲ�������P�M�k�(o�\�j]����VhJG�aҐцk�²�XzՌ�X��¡��[��M��e#�"��7	�L�/�ǐ p3&_>������d�j�����?�����&���ֽ��se)f�{4�"M+S���O$I��`�.���N�"�Vf/XǛ���u��-�i�'d�Ii輔�=��y�� o2��6���JQ��؉�d]�y��Р�J%R[����Z�3�%��VKnY��������:��@�Ros;/G�"���[^7��X6`푃�N\�
�-^��y@��'�R)kئݍ������ӌ��R��[�VҴ�ڍi~��j.�s�����E?}f񘯿����\���]y�ݶ��"q5�IXQ��q�[�܇�H�n�s��9S�yh����!�̯�V�*g��ԸjE������U�S,��,�Ԝ��.�ò��zLR	�J�"j� ����8�������9�]u[�KC�1'�Ή41�'u��[��Ѻ�)�4�~-����A%�W�n��H]��?G��x��l���U����k3Z�AM6<ƺ��W�W�ѷq�z����ʒ�(#�&�s��6�b���`=3ODP��i;=L����	D��ׯ$�R����9�J+,���I!�6O��O*���U=XE\�
ߐ�"�)����e�m>���~٣�J����e���N�燃-�@)0Q�ҕ'#�⒆�yHۧ�-df���\E��3�W~�<CT�|��m��/����-p�EN���4lL@7輏��7��6��R7��xz�Fl��j\�r�_H�s�p,�� ;a6[N?��4�WO��훴F�@�m M���+D���d�">l�&�ˮp�T�q�~�{�[��য������0��#27�b�W��𿭫,�to�U��Q���*}�
��1��~p��P(ќ��l~H��r*�fñjq���+�:����L<M �Un��Wq����TPtQ{��&pF����ͦ4
7�����\I��"������D�#xϕf@xo���vm�Td's�E5Ќ�ipoؑo�f�it��bT��G��\��u�[A8ט�����,!�ޠ��Tw�X�j�7ʒ�t�~r�E�p��z���)|%.Sn�۸�����%��+���b3�$d"sź�6���{BH4
�]t���RI�K�+��U�F�����<��{צ� �QH���|݀�r���H��`0|��l?M��Ka�Z�dľ���8Ͼ�#?�	?��1�k�
Ȯ��CI��ޤMt�4{�S���~�C�Dg���-f ��)u�yQ�w��gj.|0 �{�|��� 6��U�}�|�h�N���r>G,����������j�mX%Dk�)����:g}�IH�W9�d,��>j�k��X�$�&>����,���B��QE5w����=��j������ɾ�՝ķ����;�}I	S��:U�Y|[��^�*���+�wo��7���5$���"�/� �<�Y�BWARq�dįa��
S2v�zj�dvi��+��;��+��\�lI�+�4���E����X�̘�H�����>#�]#S�����Tƴ���Q� �;7�R���q�!������a���ݏ%�lW�/���O�EG1��Y����<�������m'��"�DO<�\�H����ؾ��A��R��/>���h"�PSVH�1���U�QB�2�����_˦`�~P̸9���h�Sӵ[�� %V�OT'�}º��8`����e����D��kb�����l��
���2Ǻ�$��c�U��xq������Ū^=$���=���5�<��I���,J�Q#�����'�sg�Ae�<��b�XX�v�o����9��p�G�?�?�3��2 ��2��1��AҨf�2�@z��(z�M��LEx��,K��=�N}����������D@�y�Y��Ɍ�>+y*���@/�� ��\��`(n.�����ؓ
I�rȥ�[<���I�"�僾�&�>�|�6��8l:j�s��ko+��sj�-�F���-`Oq5�z 'b��P�cx�=V���lIM��=��C�5������T�Gi��E(��BT���#�Z����4^�����?�������GV��c������ødX�AxO���x�KŲ�۳��mw�X)�@:�Pp��r�)4,87�:���/:a�}	]��b���b��+���::�뿗��^�D�8�K��6��p����%����P4Zȸ�q%��\� аc�|�*��Y�0:jڐ���:�	���A�UO�Bg앣w?Y��wl���U6JlV"�������l�7�u$�,H]��	�kᩲ��l}9~[�kQ�%�oâ%���l�����e?�>���������A�����H�TfǠױo]u��p`L|����>KƢ�XE��$ L�@��E�͗��=�Y�U6O��5~a�9|����)�&�U;��_d�d�t����r}�y���'�%��xܣ�Y�!��{�����#��az �����v�D��b�R Gnm$W�?Tx��@ڷ9�e�-S����5^��!��k��ϖ ������4��c>�B��t��*s�M� 7*��@��Z�.�je�����K���甴`=:�*�2s�?�K�"��&ۜK�{}<bA�5��L+�4�})~�+`�H�D
�N��#J�ϙ�f�Dd߲��K�'��J�A�1�)�0�K+RY*B���qx9-���*���}fM"����!/Jqb�%N�[��_���e�74��y9�g��H�{$��֐��yN�7B��H/lCt�;֤Ȝ��J�	;ڼ���%//��
���#'��$p�5dl�����n_j��AL��}-å�̴nᎪw�ɦR ���]�ܘ{ ��^K�������_�n����d�y<�X� �/k�!o��uq}��&4��PA�fx `7B�4���?.~t4}lY���� �*W����&��fW��^�|���n'�*(�g^c7~'��ɱ���K1� �y�j�k�6Ak� �TJ23�������sx'���������uȰ��3���2jvl���΁"M��.�V�"�	����rU�>�b�^�g��Bx�PH[�r�b�a���!b���b9��B1�M�Pm�S��b�')�dV��Ku�AF)����ė�#��m��wL=���LcQ��^�?����xF���~ܼ� ��Rz �rȐBIf J��.��r��9uE�;opH�җ�1:Q��Y��ұʩ�u���?!걟���/(sJ�9j�3Mx�w��n{�>P<VܽM̂��S!�ŋ�.@����`37����W`Ȑ@�������|�K`齀��<V-,���_^���Ny����]�H�}��u=i^5�L^Ǒ�e��*�L�-�7��������\?qK�S�eg��%����b�M�(!x��֩��?��J���݊
��lu��q��$8ͼ�k���G���s�o�Y���#�\�%�w:1��a>D=9��*<jSJV�-{���\ �G���|�������@\�[IѢ�!&N��T�N����
�	'U,G���*)��QG�pp�B O����n��a�5E��
�â�����J_�y+V��O��eoPIWm7|��x���h�����[{�hg��[܊���M~L��g�	���歅GL�:p�%����f���0yf.�zcV�� ��+���%�P�0�Jvju�vipw$��:|��'��at��Xܮ�#��Z���dc���4KA^k��,_�P�볪R,��n_gq�8#U��'18x�:�1@���T��{ܳ��173~>E�HB�	eϣ�?��Ky?RI8)x/5�sV�e�T�뙥�T;>|���m����*�N�B+��V�]21�Df
ۿ ���oՒ�C��0')V����e��y����PA�W�#pa.d�cK��.4H�Y��qy=#��w!C &M}⫬M��d�]o�nRM��$ �"��<�-��y
�"������D&�W>�V���{�&�@�{���o��@'�Q����0�&4
�
u?�j��s�̊�4��^�X��ؗ'~����`[���&��Тx���[_�x����-L�S���]��c�,�8�&��,{�>6e6ө�i�,�A��aY��l|ZU���4	�O;'d�,[4�ُb��l�b}�	���ïuf$��������:��fI��ؔ �x�b��T�y$E֚�Z�_�v��������:�}f�i?����B��-�~�8�ewNktf�>���@�bW�T%|-?J�O-����
��&m�,f�F;���y-S�� �{Ip5�����.�\m]��J��M2f1��>�R�<�bJo�`�L��*��Z��f����{V&&���f.��;�pYH��X�lf��F'zZR:���m�@0��13C_CQ{ULR��L���Ae��ό�)��c��u͆��B֖�_ZǾ�ܳđƙ҆Lv7Eݚ;�l��t*�]��|+�)�bM���gJz���f:�9��(1�r����1��|9P���A����E.�Ǚ�"����om`�ǯ~{Cq�1�/-v�v���3��a���h��4�4Ga|a�ZY�}�@��N���B�Gǥu���tjx�1�\�*�$��ӆ�g�a�����	k�Dh�7�z�|q���l�&�y�X���Mo�$4��K��8��zR^|�9�KU�G�����@S����_���5	���O�s{�\!������^�?[\���%:�)�$?O����z���P�ź��T=A���M%�="@'aE���.��i����(��Y7�mw#Z�\BC��>ތIy��e�:�M`7�J#|T�#?>��4�h�oyb��$/�PY(�M>U�� T��ĳ`���o�/P��rPE%�C�[��[���b�22�pG*��x4|ܮ��Le�]`�O@d1�$���b��sB+Ʉ뾫�BgW�3�=Ǣ�R�'�Ÿ(�zR���S7_����
�e#�������ޛ��v F�L	YŜ��#�IVaľ3�F�1����"�o�N�����t
X0�2��:^�6�BW� {� ��˴eWPb�8;̝��v���ng��o袊Z*~�}��?����_��}d����f��s��s�1�o�R;�P\2���f�&2���K�U��&���,$���~�-�`��q�r����h��$%,M��.�=�n�Vvu�˙,!Α�:�믝�]셬_U��`��r	�FJ��iB͆P�<-Zn��:G�mvȐHn���5p�o_�����sy�ʦD�:�%��*���n��a��"c�9����|JH�(6�3��u�T���Hf�l�r4@8z� �g���|z;BCi'܆��V�p�u�����a�_����[J��{�9�<���1XY�����U��)��W7���<HS�Θ�٤�ܢ��.��,�)7o/��R��h-q♶�Jn9<�uVq��.BۢX��M��ÏoH�x�#����jG%�c?�%X;	��Z@����j[�Dj]����FR�?�݋vb��_���J
X�	
�d�(v j~Y��-���c	㤐oXu�%�0�t�N[����C��ƻt�WA��ߵw_�W� �%`8a0������=��6���2�\2꤅�mU؁�\n�5�x��~�B@���[�-l%��|���
�IY��'֋d������]R�U�O��;|[bɳಓ�e"9��]ƍO-�� B�Kj�U��oTad��� 0����%��
��dOg�BHg��}�K��^�;�_�;]Z�\s��~ƭ,�A�$�_n뽸KCU��""~MRD	����R;�f�7��/{�i�'~]��g��[m�vɝ`�� ��F�x[�,�.��W��b�Ύ�7Puԋϸ���xM�r�__�'�=��+�,B�6�
�2�E9�+0Gl](x� �r>�G����ތ�O�Ѩ�H�JK�R�?:!+� d�2w߇K9�0��]��%��r�i�.�ѵ�̛9��⥼��Պ�$��{�lF��ط^�܃�S�YKT�*B�����i���۠�t�]�s)f�:? �]�=�屙�^�Za>@�ЧsjF�J���E`g�P�rʄ��[�˔�|�y��\F\4�c����7t��e�tx����̳8�F�D{�Cf7[2P����(�G�6pM�$t��K�$�O�W�)����0P��[�3���PN��NlMS�异��6^4]������I��>6Ԩއb��jh=vj�r��F��yB�R��Xҁ�㿷��>ﹱ�����]]��+� B?�%�)�p��O��f�;��G
QFZy���N,����V���̓�PAM.'4��0S�%iF�0��v��u/k�� B��Tcgw�(8��Thѿ�A�M����*�us�s~�o ��2�(A��ƞwj(��Rb)h$8�&ڝ�0���kp��.����^��e�w��|v���$l�ҥ*b܅)�!�
��7���\��)?��0Dk�v�U^��4�7T8���ԒH���+�S_������ �@���+�����.�~EC���lY�����%�5Z_��4�F	�����+B�ET��\���\f�F9k���w@��W�he�k۾����Q�pc�^�мD��N3n�G�:�!�˾K���L+N�!b��`���q!�V�b��_x*��6�H^N�b��9����'�+GI���d���V���L�u�	av���V�%��_��������}��&%`�8�J�I��H�I�MN,����J^}$H�DO[?_��ٴ�q�ߒv�~GJķ-�PSTd�eWǲL�5���^W9M�ʮ2��D�A1<����m�7���=7!��k�3�nư��e`r���YO��/6�c�"B��UQ�-?���T9A.hh-O�S��M4v7Q�	u�6:Gҝd��-���
6&����I8��f=L�����J3ӻ�O����(�uR(L7W��W�5x�;UgW*��������� -��@�#G�KU�?a8� �0ȗE�Y��H2�T�.}�\U�bD�CYW�� ��c~�|V�N'���oЛ{�e��ǹ�YԺWRE����A #fN��+���R�?��9�w2H��vP��/�u�rtC�.F+���j⭖ݪʿx1=Z
��lqQ�b�췪&� :l��A@��mΙ��X\��~��l.�)�iٺ'M?Xр$�ki�L��|�E�O����3p�ۢ�Ã��-��'�80cs�YS�W���rm��+7>�����M;>���ݠ�pw�����W{��̴�k���]�]GHyԱ��9�>���ݛ-����q����r\z��	j���|����������	:.����@��q	���*��I�:�Sc��M[�3E��@R+��"�5���h�g��kZ�pb���]V��'Fz\�[]6�&��Щ����
��ْ���B�$��	&��\'�Z i	���,���ttE�e��m��Ӝ��[1����H�P�YKk�5߄7�(���(f4������#vN	IB�M�'0���^Pb��� 2Xwd#�:~a��6�OJ9-�յ�����۴�G�P>=V�Iq,�B�|���/��[�� �Q*�_��c�"�]��Ō�� �}�� ��Nv��o�f�7>���Ko,��h\q�B��*��2jM#���"�1ގOT��LɃ�vo��U_f8#n/!����	�ж�Vn������?{�y�Z=y��o�hC��$�R���J�Cq�Xv���!W�F�m5C�~"��#�"�#Y.ԫy��F�I	'�3WyzEp"^zU�rϣ]+�8c.J>cen>s�V �$yCIK�?�4����-`ѻ!uh�Dn�����Ԕq}%��mP����giФ�����?���@�_�$��>K&�L��A�xV7�;����+��c�ιm�DNc�t�Ɇ�d�bXՋ�����^���P-�[�9l���@�E�ƌy�k���4ɍ3���+[,��e���Aꏒ��i��	��T�|q������/
<}�9�|;�+W��P��j7���TŒ�
���h�@�Zp�S3<C�Eō��Jٸ�Tj��k����ol�Ė����pm�W''�+"���z����Ww潨Y6���Rȸ7g;����pf̅,���ab�g:h�M~��>M0�^� ���lu�Ks�/�gy!�т�@?�c�2V#�u�6-��!�|���[��Ϲ#�;�Z���\jS#o�Y���-$!Y����u�%=�&��V�~)��S��K�{I��,�J�<!���<`�ݻ%]��|p驂��H(
��?���dm��Kx툶���ǒ�w���\�Q#��y"��"x;��%�nL1^��-����o��ᄀ��n30�;�?-�V�g$�bf�4_%�VP���ع��I��/�f�XX!�q<C���s���$�M��F�7f�3o[{R�a�i�W*�_�/��g������^z�����2���C�6�)����w�G�}	��s�e1�l7��TI�Hi���ͼ[N�څA���X.�?�Zvl���'e�:���kE��ω\!�S~�)Y)c�i���{+�M00cП�E�W�Q,F�y�JH#Z�B�"���q����P�������[��r�N���N����11��Э����������>`�x��̔ފ�W�u���$B�r�Pr8����=��Q����\;�H��iq�`=�zE�n!Tv?�4��Ip�4	(&�N0�d�
mJ<H�H��RW���69'����e'�V9���&HZyd;��/�'���ӦN��1�B� Fԣ�B��� M��y��oh�xyFV>�B�3��M,m
?����j�	vzD�Ҋ��Z-aLJ�:R���Z�y�5s�̜!�|k�&z��6ꚓ���&��a3���nrL��<چ����fԷ�|c�A�ҷ�e-s�V�G�[����ynڎR��$+�Pn[����_m��ְd/���'-��7�W�Q�8_�$n�9c����ᔘ������r'�����<q�d�Sf�-N�0�Eg�H6�@Uw�(l�gK����Cm��.i��s�Hn���q�W/�����7�]X���?jʇs�m9���g�/4��� ��G�"�x�ƏE[��8T�6;���c�9��r9s�����P����o=_,i'?�����))
�R�;�!�1����!4�ᭁ|Y0�m�F�yh�mʽ�Ɨ�a|�ܻ��#��-jP?���{=���t-%⟠,��}8�������xw�^�e~ywS7F�G��gN�?���cS�$��t�Ua���7�������b֦���T�_��`�������I�\����x��D�qo�� v�������z��t��yeʰ�H�|�M�=�Sc�k�]>ِ���G�<
�z���A�Ȧbi����/�|���%z"�=��.�*c����䣾�q�^х��[���������;�pA�:�@�s�᩟9Q�#*XQV�5��}
q�\@�n)QYl�U��W!s�#|�m@��7��\d�ЖɬK�	��aN߳�=fm��ԝ=;	&�bt������a�%k�`�/0��V# �����e+�V���gNr;�v1�%����$�������9'�*+|�yr͆��A4�)�+u+5;��� �@��u�T��~X�[��!e�v����7(䈠d���vw��*�/F�Uʹ�AD}i���c�eEw�c0��R
G�s)���sI��L�8g�`/%��Y�Vc]��H�;D�Q�ǣm�+�X��=��/��W�hL�8mtn�Ö�9(����C�������|�p�Y#�/3��Qo;�ɼzAp\�GPү�X)��p�e(jNi�ޠ�$	Vf�ާ��܁(ѵ��O̊Lw��������A����:����P�p�p��ki�����4 ����k�[S����ܡ �HoL���QZjP�H��~�M$֚��e�qhr����o%���6�9.��BB�?�c�ׇ���9Z�g |���tZ�����dK3�:��I\��t�f_��;Ŵ�cM�0�i����47��^_pj�vt���w��C�8Ĺ5E���>�|�58��<'���ڛÊ�Ɗ���_ߞ��4���u� я�_�~S���=8RV�{��0!d�:��rj>/�JH���=�hx��H,��G�d� ���
�@a��1�_u S��o(�;�'1'�;Q�Q���j��3]���O@A��<���wD�7��j���{���_����Ϗ��W��z[ű��3UK��,��_���;r�@�-�<��}�%��`vO�����G��,������{��@�F�~�xÃ�j�=��~��n�2��~Yc�T]J*_F�3fڣ�N�$*C����.57�#!���S�o ��B��Ol���n��4�~4^��uA�c��*R�=��&��q}s�H�����f��2%�Z��\'�. �a�TW@^~��+�!�����}��7�� :0��5���l�P�c�
��X��L�?�r�lc�-�A��s"����0�����n횹ۇ���r�d�5L��g���8QJ���^�	Q�Q������f��<�P/�E�_&u`�"(��P-����h)� X>��E��TY �f1�	���)0n}�f���Zdf#���"�w��N?*�E��fEA{߆VڻC�;�,�e�1P4Kw#�\�w9��ݍ,�b�D��AǪj�\p���qVϦ1!Kz�ب��EK�`r�}���y\~L�o鰄����^ᅙ#�u�|u�/u�H�=����,���O~������0.W�7��)j���?�+ߐ�y�� )A���\��/2-)@d�x�X��'%�2$�kCZi��/��ko�[v�-�Qp%i?��.:>#2r>�|C��t|ڥz{Z��
�?K�JH�Bӗ���@�v����	^L;�3S�d���~���I��)AӰ��'6�`UR�V����G8��p�_C(�]��dW1s�m�q�|/e�3��1}%�s��E��e��/��驫S�F�mQ���Y�������/�g�t�t�7�"\��M�;0*�G���ը>��nD�F~�rwb���_8i�Cf��cоW!A�kb�q����(��Etrf<�I�7������Gu`?�9�� n���{�ό��k5�0��u$$����VlS�b�k�A
�X
� n�G�5�߄����c4ME�x�-�O�|۱�;�>�X�A-oW6�u� �S�a�|.S�u�.AL(!0$�z�������[��@͒�R��݇r(�
g�P�<��9�d|�*Z���sZ��>E�b�����^���D����;U���\sl�p�i�J4k�" h�8s�mӆ� ��jF�J,慩���d���0��"�F�j[O�ulU4���ő�ӝ���5� �l9F�����	��2؃U�2��
D1Vع�S3����%��6�*�^�u��J��9	��ot�r�Ȟz,��p�6S���H����{���>˖3��A�8؅E�"�2z����� �*�dؾBe��ke^�\?�2� � �ϔ�Ĺ�_��t�cc�=r8$�'8���E���/���W��G��8�a�)�
���p�$�9�&�H�k]e����[�[Y���K~4���[٢fR)�����I7�E��g��Gb��=C�:�~�O�ؤo� ~�+�Wid��c|�Q�v>W#ZD[�q�R����EU��%������;ݩΨa7���������k�$1Kڥ��&p��Ey\+@��H�C����#�:uE�P'TK���h(�TO)� |��*ư	Q�~�.��V��#�w!�2Љ���3����y�~��j&�l�@f4�>���8���"��G*oqR�6m�Z�����R�V��1�<z���#�Qi�7㿅�DS�Ӛ14�T9��4W}r�8��n��mn��oZ��P��tſ-���2 �/��`��A��&I�IE�׿�E�'s-�x��Etύ�MG���K��D���N<!��]d��XИ}�m9+VYY,�<^+��-��A���v����5
�45�.A�1�NGEq����,����%��Ȉ>�E�l��w�>���_���k��d����e�:o�'SM����e�D[��I�i-o���&�	ڶUH�<�n>"��c���/��EP�~Y�ه�H��cN�V�lk����}|yH���V#ib�A�ɜ!��e��W�=p�X��s�-3��E3�D����8��E$w�$Y�~
c_V�@�T��Z�3N�.�Kn$���z��'�r�(x5'Y�w�,���u�4x������j�,�kĥ=��t��J�w�r��_�i�{�5ɋ_ `�M�wC'�HVp%!ܼB��7mG���OR��#����.V��O�Y�o�e��l&}�<�!H煆��B� ��3�v�d40�%��{�M_D.����?~�@"���Q+g��!}�4Nb�}�Ho&����	R�I_���3$�V�A-5��4땈aјv��M���:0�4�k��Z�}�����ё���/�C�KҐ�Ii%vRt��� �������M�pp� Mښ�lFA�1� ԑ�}��ؗ�~7P!a�u�����X��Z2�����|�'#h�2��,u�r�"S��[��I ���M����s�o���b@��3UN�$Q�c�Y@_Bn�s�u� l���#�3��"�H��r[h���M]��3 �]M��w�g������U��STl&O.WE[K}0�Ӕ��f���Ơ�Χ�o�'���s-�
R+Z��Иmi�a��=n���)�'��S����~�P��)�nҧTc���2�����Nq�$����p��7	H����e����Er %�/L�p�A��A7X˺��:v.���G%��)���u1B�{+"�;���4���Ď��̋�0����u�>Omo@Xs�3?-��}0�jK�2�ω�!ZǙ�X%�-%1������7@;��~㟙G�+�'��g��DSQ�<�f�ǫ�8PsZ��4�P�
�ͺ+\�k94NCV@�|��o��D02�f����t�8h;�?��Z�.^���OC�]�MV���畔�l?�^kl��6)������f����}7�H��8� ���1�v�%-��Q?�}}-60F��[Y]L+9v;��&�I��1[���p��@zy:c''�F\J�Z�i��'d��#T6��0թrһ �d�] �e�$�d4�μ ���v���)�V�� ���-���[AJ��ƅKdF4e��9�qu�B6�yGx}K履Ѱ�!�
�$�M|h=�_1��y� 6��%e��+��f�)-8�WV $�.q��b�? ;�#V����t���wW�%q	h_f'~�����>,�l��dn��N�?RӢ�e ���<9Ѻ.{�k�t��[B�zg~&
6Q�t�Mأ���zQ��km
&��Q$1��A�����^ ڏ��ӻ���#Ч�-b��C�����?��lu�<��k�<����v_�f�^9j*QQ犩��I��(0!�|�Q��x2����퐌��~!!z&ڛ����)��F.EGP����ᐶ
����0P����]�L�B���ߝ���Ë����.p����V+	/V�m_E^�����C�J<���3���ۈ�U�Յ�ܬ�N�ƍ�N�zJ�Ȱ�v���Ƶ�V:1��?���:h)�@�8�!ϯ���t�|�qw�9R.�!�b�� �{.�Q�Ū��4��x
�����휡�\�ϖ�M����x��z]��2K��ݯ��Яu.>�~��Q<���W��T:�{��}vAk�a���������n��E�!h��?[�/!�Կ��^LY:cX�S�{ryK
c��9nM��IυPO��ճP�}�,X�I�uٛh����U��|�=�θ�
.I�Ǜ��	�1�i��
?� ��%�,
��rn���(��H���p��驓�1�3�Jp�}��'�� �� �ԡ>���B4�I,&���A6R����#|�d?��Ð�#�)�h��MGz��=�l�ʹ6y��7�fnfO?�U;zW?	�qǭ�D�v�)ߍ�"��L�*���|��㍨� �Y>�	�����D���3��n��)��/���F4�J.r�~�p��6�.��FCb}	��pX�hr2c�APk�&Z$&���,����~��}�m��/���rC��f���V�&�т0��XA��}�t�,ː�-ۭ�H�R"=<<���F�9���k7!���[ޖ��`�kj��v�	⦎}�����o����c6����M��rj)"B��ؒ'
��0�0h����wǤ�=]Ôz�bNu���w�h%��)z����2���L��9�	��(gwȗ�X��s�<��$�gYB�P���!��tNp�AQ�ӂpw����΂�����N�̓M�����z��P��M���V���w9g�b=���K�lX���/B�t�T�ܣ����N�eůp��e:��"��A������`�a2������q
[�i�:��3j��?}OX#��5��Lڄ~%�b��3�ѫv :��B���+�0�eq��!~��'l�1�^}��N��,s�"�#q��8�Y�y�\R�����B��yȆ)p}{�jمY��EY��Xt�H�fӆO���w��B�[�������a{K���C����$���P-�M��Cp��uL���i��^�-��N��B�[-���x������o�Scq?|��I�vJY�n���~�v��p	[�F:�5/2ނ�/�p/�)mBzɤ��y}JMuK�ǡ|W�u!ӥNAP�[)�*��*Wɣ�h4���������0<S[�Z�1�&���hظB�<B����X���)��>��m6���L�r��k)CF��md��u�4�^��j���F%��-BN����N�EV:���i�;��zg�+�����bUM�4�!�E�
�Lb�X���o�v��<!���ǐ�YC��yMH1���� ������2�����H�1i�9"�eM�f)>�Y�m�q�� ]�D�I��m.�]�	�ٴ��Eo�^�đw54')�)���M��l
rh�����m�|: "��B.`�	`�M9�N}^Xi�I�r�Ù��bB�&��A��"Z)�����g>�y���\5��(Q��o\�6�]����J�ɪ�����ߢ�-��L���/F��q?��v24Г�٥e�P��*u���7�=Df��CH��ҩ��^��.���f�R^���"#�ͷf���s����#���0�f��`ur[v�Q'�W>�Bt�*5�@�Ѯ*�4l�7�C��ּ�����HE�t���C������9y�fI�%B��uWId��a7���	:����]T����t�ܦ5(i1_>�Q|3�����H3�;%��
@PJcy+�@��i1��S�Oj@UB��ː�H��}k������C�h�&�an����h�%(�T�N�'��b�s9��X���Q���i�y�ݷ�9���=�o���)+|��O���wő���	@&+2������
�ա>O����Zϧ�8�(ζ��2�Va��!,|��D����V��!}������}W��Fg-�߽;�����yE�V"-��ʐ��,0*��v�S����IFt@.���'�>,uV4�)4D]GKg/"�T�S�J��R&����D�eK^v���D�r��I~H��Y��͎\�Z`���#�#���B�%��&�E���<
A�jK�=-��-�p�Rm�%^ptI��߁��A^�Yݙ��@¥��+3�^o����Ǣ��jH������<�)L�P_��j�=�7�bp�&'J'"H�v*��6�2k�X�k̾*?~v�yeZ[�[wOt��|�蔏?�?}�:�j�&�橃�5���j�1G��㶫A\˿�_tk�YX16Ws������b��u���E<�Vd4�[��T߀f��"�	mvfyL���R?Yo:�^.r��ma���}�y�O�� ~E���3��c�=O�W�{��by�t��<Ou7��Y�NtQ�Ā^��귚�H����@��}�S[����$�[S�FG�x�2�.� u��~��~�<��9�oVa}��v���b�:����Q��v�>e�*�ˁ�!9yq��'Nu�V�U\�����E����'`E��Z|+y IЌ����\A��24�
G��v����M��O�`2Ʃg|r�O��(1<?�x�UH'QܼY��{�%�C��l& ?u'P	V�RR���ȋʛ_�:p^���I��ыy��3W����A ]/B827Ѝ�[v��|j]�����TJ�~�$5�j�8�A��.?ۣr ��҆��R��k���i�x����� *zԑ��5V�E"r���6"�sR;���T��4h#��	��< gi׽wKШ�te��Ӧ�
�X���r}�[�)�>�p���Oഉ�p K8a��"�����{cV�P�b�l1z�5��L�Y�U��#�0�O��Y���og7 4��r���s"�(߉=5q����E�:��h�d�ĨX�]&���:B��[��A�( %�� ��c�^/MUz�v0�k��,�ԣ��0�ú}�,0/�߄O H�|@h2�!��b�F�Jq�}��v�+�.�0]�>�q�����:᝿&�>��֦�Z��MG��C}�R9hL�Ex����_��碂���("=��
%8�02��T6L�M\2m	"�
y�kS���>�e[[��^��uDLʶv�]+���'ie��!QU��	K��:V�j z��!n�� /"�o+�*�Q�NY��ݕK�����֢<-N� �f�'K��?1+��K-��D9LBx�^��)�i� ���F��1ɋ*�Q�8a�y�gf���
W�Ӡ����8��ϫP�� Q�@�R�jD� �hFm�
�d���<ptݗ�8��6k)�E�ZOy'v$�� gv�޲@@!=ѝj���~�pb�����g=v�Da��qs��T���4��@��A�\"ɂ:/p��-\/�݀�*�>�v����d�K���_�t7�gmdv���M���2�k.`($v�C>��'9H9{+�#8���������C��teBO�}�%Ԭ���X�#z���R�$�t���V���>!Q3d���0a�OPᡡx$\���,�C��fM�j�V�ߥ7��-%�3��`��1�G39?O�2jk���S����E'�hG-lu����ᅂV	�C��\qN��������\օ2b�>+28�j ���b���: R��"6�䡴W�yH@�NP^|mÒ}�tc���0�܌A8T���CW�ew�͌��{�J����l�D�nǦe�r�#�+غ�XD�4�vŬ��m0��1��i�e,�d�_������EE[^�c�Q-H�~`��x�L�4�v���3�@�aǪ';�ҡZ�1�^}RTɋ��*�&����>x�l�<T�T�+0؁	�tY�$m�i�XhE����G[���P�޾�|���Վ�Vt�"�w�Qi_��K��X  �sDX��B��{>X�q9��yR��L	[R�+q'����>M r����*Qu�%�H����bq)�W���ܡ��{��rfY2\�<:�YQ)��,Cl�����:i怆S��7(P��o��
5`�xrzN �N�]�&�GS�̈��
��^���.�*}�Ο�`�oc�G��+�	�zD��6�ƭ��h����\��ڋ���_W���
3OL�w'1P�ta_U�_�oU��(6�Wk�z�7���9�����)�R�8��C��/��|Y\g�V����=��	��1%�����w2���P[nd���4Pz���U`��^����#�L�V9�¾��G�O䚟!���)�;H���晦�d-a�a�*�FS�3R�R=��e`�jv5�J6�����g<�a�v�	�k�F�)�d�)ϫĖnX��F����{^07I#
�oΝ��%"<9��n���c�w���E�T��5"�X�uc(�ܗ�����(2G�fE����̱Z0��*��r�[!��r\2N�$
��q��!���g,^�k����Ik�xB�]R���'巩I��@e��F}>�>���Ո>r�\�����$�PNx	gf��f���R�h��q�Mi��{�p�ډ�V��a2,yt�zD/��M2�w�q�,G��V<�ɾ�����B�MiX�CeX���C��JE�}j�h��?ھ���_^,L��s��v��>&_����>�74��S���u��
�-�ye<���W�E�����{���GO�m�OA�	���B�5<�	��qNP�x��c5�t�[Rbp=�p��k}��ݽ�8"h�2ҝ�����9��S�*C�(���r���E��w!q?��0�d����#ūf�����^�Oe`H�K^�]�ʹ�L�Ne�����N�I�'��鬒�)8���p����ro���eKR����ss��N|��eȕ�73O�]���6��}�򂿍e��^���f�y����aH�11�"�1q;OU3%m��ϓ«����j�`�����X5Ӫd#����"Eлf���nI4����}��F��m����9����t���p�`�?C8����JO�s,*@�\�.Y]'�"��. �Eʻǭ`����!�.2����ny���U��đ��eE".�|��ԖϘ�|f�Y	c�9z���0��!�H�߁Ēgf����H��T�*���W�_��Wx���O�
I$>��{�b���Օs��{ii_<�y0��M* ?�	�V�	m9[�͸ƚj�~ϯ��X^��.����e�]C�������kR��]UJ"' ���w�IjG�E ;��������e�D�6M��<�\y�S��t�3��rA���h]��c6@(P���n)G겯?��A�J�A�g��K�N/��&s�я�˱L�p�.�G�J$a�*D�r�o+\��k����{�VY�[8�˹�G�A�.;.i�\J?D��Ĭ�(��~C�$��Fo7(Ap|�8Z� C�{����o�/�ݙ��$�ѡ�dc�ȨĻ��{}D��
�+g��x9D5�ܧf��>5��{�/��6k�ŻB��N����`�+��0oJ�;@4[�	���ؒ �)�p��c��_��'�:��x��Aw�Kl7{m#�W�vc�k��9������q��p%T��{�UVd�b6����._��7s!ȤN!^�`k��DZ{�11��W�s��E�(;�FX�j����- �#���}�@�%����eqӗ�vD�M�Lf��{Y���\�ԏ�Wzi�ڔ�L��H��5-��*'�Vwɭ@?�T�a�	���� c�9�Vl (�x�z�tp�xX�g��K���$��l.���E��>�-
�ۇ��P.�)=Z�h��b��˪�"2��z8�����	��@�eW�ast0K�7�Yg�T��|+6h��'�\�&QD�`��駋?�̪�,s�I�{m��r�8��q��y^a�0�/Ս��]�ĳ��4_桨��h�V8<nkc��x����	/e��' ���Tb�MK�r������d�"owE���|y��[p�3JC�����T=#�-z$��fw��FI0 �9J�B��Mh�h�����s@�}BRL��fW3�U5�&�c�_�
�j��ۺ����+䕒`�q�a�t�7ޝ��f+�P�z�G���1��;��|���¬9��2��cr�y���byA,���C˭6tDi.1jIS��°at��P����T�ry��e��|��d�1�U�P����+���:��w(i��
GK�筨������a�,y D8g��#�]¦��������(�jPpCv@4+�mIv2S���V�f^^B�ɧ���
��z9�c�gRfG[1󪐀9�_���-8sPQF���D �x��q�n	"��b�������i��6y^�@����\ا��o�ʭ�t�O��?� П�֚���E����<�]�M�������]�XxX�{M��M�={�4���݆�UP㉶̚�Y-����^��L6"�9�K�5z��N2�`�V���A0�iA�~X�Q9��������hT^K;�gg�Ng��U	��b(jxF�O��.p=�uTb�c��]��o=d2E^�C��=�O����F����3�m���?K��16���1�xZ��$�j*��`���/q" �Y�op��8��
����X�	�o7������ �=f����i�9%~�]�����N��"�
Z\�slz�DW�u��"�2��k�l��\~��=�@�Q��>~Z���[3�>ݥ���Q�ӱ�sN[�¨���@�v&U�b�I��>��9����� $/�G�[x���֠��^�K��M,�5��@��Y������+�<����|����4	&�%ײu۴��$��$�?D5��,&���~$���%t�8�Y�%:�Y�P>�D0Y&�0`�h�{�G=�OE�U$�5}#�"���/e��*WT�S>W�Y��VO.�-̲8m�a�i/�Nc %�o�J�!��<�������,����t��0<F�A�{�e�����kȮ&��3yf��"�\�w?����_����Lߧ���P���N0���q��~[�d�����Z����3���U���� �<�W�Y��$z��B��4ڴ�跹RJ����w�j����6v�VI��z�9�N��wh���3k	w��bۘ����1	O���qADư�᏿m!ro�YN^%�*1xn�a�ɔ��U���aЇ���i�{%o�&Ń��"}?����ioߩ�x���0��oj��#��p�d�a��z�S��՟x����9�7'�C{A/�;�eZ1�?�"Y�zz$`U�o����ah$�l��*.oϤ%�P4��W�|h�є�:dJ2�q�dt<�	qö�C��g���Jz<��جe6�5@���{�%Or�N^��������#��q6#r�H��bȂ����-�s�,@1�bF008�l�9��C��xn;(���$�����H��Q�ր�l3��c�����S����k�P9&���iJ�^m辀;W��t�[��^�a ���������ά`ݵk��+9p�5�t�[�i�}���+{(J��)�佼f��  x��|(T�Ѻ��!�;V�<8oN�/67ˢ��˵�Y�	���j��n��~���.�k��I�Ē��'�NW*6h��wc!'dTkTi��!0K�sw�S��0�����RX�3`҈�4M����k(�αr��B7��0��Z1/�m%_s����4Kg�!�0n	��i����l��1�P	�凞��]h$T�2f�3��9�f����k�$e�}F�ڡ���l�2+|?߿���c��:��I�9L�,���w%���ny�7�=KD3�A��m��O=5W̳	��Y�+��$bmn 7ծ�Q���'� o����~�%�� �.5��&H�W���R9�||Z4����T��h�w/f�T��$#��=@c@!�u�;(ٷ���1ń���o�|{T�~��)��������SUg\X����K)���ӶA����څMPvj��
�-:-����Q�$����ִx���R}��te���>�̩�1~��lEͺV���4�)��/;�f��8���K���K�X��'�[dĹ��I�7��8��e?��U	�Mr��K:�7."�3��M!�?�-�6��:���j�,�#�Z�\����=�J�~=�n""|� �:�L���*�`�d�˝g�O�Z0�(l��|��r}���V-���ɯ��+l�����(�J5��΢��
������YuG�16��KǸ�ⳗeg�9�?]�Gc��VŢ�u�D��%v��"��z� �tK�W�
����rw�97Q�4V؛zn����AN;25Z�����4���H�KE^�Y/u]Q"��]d[�ay-;�K�lv�pT�F��W>4Wv�qC��=�d�U��y8V�-�,� ��� ����۩//(���7Z�(Wg��e�Ç�>�i��"��V'D�����yw\�:Z陻V��0[rQ����gWO�I%h�ԵU�3�z�cm#5)�VɎm��?z<&0���/�� ^D�鮚�U"@��^"�����b�x�X��Е�Z���:l��:�7-��p!�#y�Ƶo�rX��	;.g�Q�u�d�-��$���k�3I^Jio�="<���l�'���G���4Y�r�U�+2��b<����n7G���6/�k�Q<W�t��a���ω/�>S�=��z�z���a�������x%��2T$�L{xW�0��� ��Kh1Ե��?u=��s�Կj�,����KE�<��~�lB{�c�A�q����X3�l�}T=D�<a�i�O�~��rA�H:ײW};t�*�p��'�ҡ�5�-��Nq�� ��wMxt��c��L���7�����[U�������S0��X|t=��,a�@�=_���v8�Ͳ�KA��~CYS�2w'�I��ٯ7J��t4�	5D ����%ԟZ@>>}�8&Btխ��'?� IM��׳!��(�l���ZI7��@h!�B������j���SXc0<����G<�_eJ�kf�N�����T���CWIH��3a2�#�[�C��	���_ګF�� @K�/tg4;����*�6�K�M�Wq�6D�w��/����6w�
NFP55.��S!��R�6_�@4���Ъ�/�{M�^$ˏ�	;w^��P#h8X����7�0��w�v�B��S����;l�a��(�T��K��.�A_�Zv��D��M���������s�r"O�.�EP���1�A(T´l�<$��G\7iʐ�8@�Y�:ӈ*=�����/�!�;�����͝m)�����ǂ,��SQҊ|�Z�����	�P�#�/���8WKT�ʵqz`�_tbS�x��&ko%���TA�r��wZM/��ҿ��q1���Q�ʕHP˓Dn��S������ �/j�j=H�$�4d���x��	�0}V�~���ŅbC|����`��͔�j�ܔ����h�l>i��?TCTC��R��2��k����m���-��/p^Q�a�7JмR}>���C��j�٣���|Δ^S�vOa�{� ѓ-��g���x�������gjnSy1C]:���R�kZ�){O�q`�N�1��Fґ�E�Q���4�g��{�,L	� �����Xl{�#���c�2"�=M���#;[�
������G\�-����#'-�k�����׬�_���p��}��7�G?��K<ʩ��0v��U�}g�8��'Ũ$Ư��0=�7Q�˵Z��i���e�>���(��FKy��`��OK������1��j�ŗ��X�!rH{�.���G��HŹa�%ŇKŜ7��0�G�R�GB�[�0Mh	U�pP��wa�e���â#����|emў�Ϛ+܊>$QLa��I+�����/>�ut<iQ���Q�T�0��z��҄J1�b�������0õw0l��u�����WM(6�!'�ix�	�f�h�"Fg���i��E��U���ԉ˶���J��]��eE�����s4�^Ou��ey1\S�1Cv�䁅̞��k"���LR���^@wV2� �kq��glnQ�����D\���*�S�,���p.�
`�^�����L��Ơ�w�fuyQ���A���_PPZ�3�'J��Z.��yp?Qt��V�p�0��@�OM�K������h��
�E�
dv �H/�H�	��i�h/��0�N���c���EL�L[f�ƒ8?N�L_k9�1�
H�Q����)� �_f�kM���+f�H���OV5����������;���"H��s��s��,�悥��U|~�V�]}�4��!����JB�2���1fU�Nu��P����U4��v5�AY8��E8s�RX$_�	�"B��\�9�@\���^|҂��7BK��奇$�M�V��[�g#��B)�=h�Mũ �C�y��Q��nND�b�Z�K��/[����=7	zފ��*g��s\z�6p����xX�)M���c��A�Sb}3xնYl�C�@�� �M����b�Lo]6�˷A[FϽ��Z���E'���Q�<s��CF�g*�p)���p�ϓK��}�D��[t����9�&Ṕn^iv�?�m9��dBW�ǟ1�C�ᅜ]��$_�f�R6���]�������^�A2l�'�Z��@B�n�Ek��	��B�X��(��m�O���{�=D|��ش8�yng��K3��nV�<���&�CU���ڕ�a	�o`����Q�/*E� �;`��������t�jf�A�aC���8�i?>6�h'�$<ȏ`�4@P��y��&
:���H�,��E�Y�o����oM�#�����ZY���j�3m`K�@ �0�>o��`�=Z���n��Ҩ"���k�↲5|���Bo�����o=`ll�J��:Ԧ�uR�T�8��mi��	�oxi�"�VOgf.S�{���4�P�@�p�{�C�����-�Z��Q����^��Y�t�?�|D�B�n��YmS�,��o�K�D8�� J+���.��s���)�K*�Y��-���5�x6��h~���E�`�B)7�
� i���4���q;�"X�FaĻ'�PX�H�e>�P��S���:
3�*�o��}�:xNC��B�Q�ظ�3D�����������'Y�ڋ|Ҏӌ�h	0d��1��ƜC>:;|�it�^�m*0;o&�u:6Յ���TǊЀ)�w$�Lø��L{j&����ŵg���կ�4�gF��~_��'`�F���;�p"���[�`lng�� NLo�e�9���S�K� ��v58k|�ĀR�g�5��1rމ�z��T���m�DÔ�����"�J���9-�=�/[�eQ<c�^s�`�%��ax1���#���U���9�D\d���C�m�,�[J�J;�8C��cIt��.$5�?�ڏ0��q��Y���ݹ�V[:'�[��P�fj����C�gQ�Ud3�'"g�!�qg���wE�2�>���� �|��b��,쎔��L�NK�Sx����析(�er[�?���s>��J9�!f�"���e�����B���Js�BvDcU��3����B�����c&Z����uB��\��̘��"^�/�@J|/3}�d�;~t1k������>S��8�̣�.�\��]�@�y�d�������!
@3�o�KĊ�Ϩ�в(	�����m�V�]	�5�vY��l?����N0�G8�z憮�
�}�{�����o�	 ��4)��,�f[)i��`E��2H��q��Q�����.P��N���ޡ����C�QXlb��>���A�h� �Fm�B�� �|h�7,,Y���+j���T�������!b٦z�?��ĀC�xtp�u��=�f|{x/��}��5�������X�^�e�,�l�v�ݣ�<�4nL�"o�H���0�;���>ߣH��!c���` z��*'�yM�Z�=�1�r��QƤ�5L�f�q�r�!
�Pt~"v��w�����u��YQ�8a5�ʹ�
������G�Q#��!,c:�0���ѠE��&L0����{ˋ,k�RФ����8��9�J���fc�~�嘯 d��~(}��6���y������&k�u����n:��V�*�_`�����/U�4�(Z�q�̜��f�)�I�}�"�OP&�h�,Osg��햺�P۔�BѨ�,�Ϡ�GdK\�Uz���P�L#Ā��6�D�;.�LH� ��f�,҃��5�x[������H]�2�W��t���SҶ|�"^�7Ț��Pԝ+��[���.[y�{�"� 7(L$ �r�Hj��Cv<K"�FL�?
.���P�_�_��9��J��_ft-(�t��6w��l��j�v2 
�7U��3��0�����V�XB>V��<����a��{�e��Т>1��{5��~}�˗�p�x�_��=�����c6U���mV�%9#���W>�E�٩���B���u�`��*����<�G����y�� T{�c��jG�@�)��Zv��τ�?��ěR�j��f~��-K|���z����0�����V�E��s?_ɻ\��+rpl�S̎�jTT�����
���x7�Ԕ���0��Wtv�u�*�%�b�E`|c\���]�W��r�^�Ebb[Ր@ՠo���Ë"�Mw4����S ������y������p�81�g���r�M�y6�ޓy�0ħv�`��]��-��y�0������Kw����2�Z疀-�u~�Wl8�*�w��P�2�@�tN�ug�~�'9o$�#?������?�B�����'��y���B�2�����7������&���J���ѻ��Y��x �ʧ�Z�U�H+,f��kf�o_�B�����(]�	��Y(��tR���gF���_>�
����Ǹ'pf��[�KH�^ +�X��=���n����P��YMDŷ��]�D�-<�!,�{x�3]0��8�
D�xR!lb7�$�1�y�n��yl�>$������xQv !�{�y�lƈ��>��WҴ����@�԰��?9���f����<�z�W+ܟ�K���vٶ)��,mt+_H?Ђtn��z����$N��4ϴܷ��"fc�<Y�t�s ìT�ۊHN����)�M�e�t�4G3x������k�*0Q��}�y���2�����:nȨQ6DlQ�c"�4*.	�m؃!i��Y�.:k�<��8�����<ٶٕa���;����`��dX_2��@�69Y���/�w8�p�������$�Z�:�B:��m�t��<����)�����%j��vR��n�^��6���=����"d�Dꓠ_��P�(_��zfD� ��W�X���F��L��ѭ<֒�D����nŕ���?�J�8#����\4oMZ 0ӗ�"�[$�c�%�U1#L�5�F�J�x^ԣ�f�t[��)�0��L���vD�e��p��	�s���%�h�O���Ϸg�L�C�*��qU2�����g�����WL��L�L���,�N�5f�뛔4����{K���H�Wk�<|�/�u�!�����@�}2oN�"X.32��3G6<`�ĦL�ʲN�6���5�xec��V� �&��uk��;��P�˄&���o��8*JJFx5V�j8��l��?�U*�$��ċ �Z6���G����דa�:�Έ�Z#.�����to��Kd���8ɊԂ�QݘC�9��AկJ�|,@C<M,�E-ZOlWz�ȑuO��@=���ݳ��Ph�'+����f؋$���?f��э�٨��2���*B�2]aVg[-���������(�0��a||d���Y��?ux�*�n,y�����b�m���~:�~���y�Gݥ{���'��e>�TA��G�G��`�d���Yb����Br��՗��l����Aө��{����1l�ح�!
��Syl���,}����p�&S3'P���|�\�~.��J���X@3�鈔����!�u*_��ա*s�EB����A���i�7b���C	^.��a3�Mp���߿�4Ǻ��@g����㖛�E# %�ߕ��چ�{y��u8���Δ�P�<+p8��I�}}���BR:�<�m?@,�3 П'�al�#_���utd?��u|l��b���tbw&���Z��b����(\�M��T���!~Fxg9S�����<�3��[�RN����4���pի+υ��o�y��n{�[rڕ[�G�7@g-��u4^q�^�'Y��/-t�&�'x�u!2��=��Ϙ�J�]$t�,�/L�b��y��8d�,�P��p	MQO��ney�����ՠ��	w�&����� SeR�q��$}q}��A$�kjϟ!i�'�c/�ʖ��j+;\Y�Os�� v=��Dl�3���66��s�����V�n�SG��U<�o($��B R������C=�������#l���r�}>*�\�d�{��6� ��h�cϤ�S�-WA����ӯX�bJ��{H�}H��D%E�o�G�-�"��ئe��%�}�����I����3g�?������^0�,�D�sy[�mٟ
�)��Q�.�Ӓ�"ɊY�Fh�pj���F;˛4.��DoA��³��_(7����������[���@����5=!�_��6�+,RS�.`-S��߇r��z����\���,�%�6�j�\8����җ��S�=��|�_�Īy�[Z|��U�������S�Ds�#r¯4�9��L�ke��M�|Ө���)8��� ־�B(�m��M7 �(
u���^J�̓��f*��|��P��RD���2���=�`Qͦ���Rk�s�f��c��F��S�S��s��/Q���S��[V�3�g-��s���&���LE�c�o�|@=?M',ꕖ�Ͽ����;����q��f�9@��\V����*A�ē�,�đ��e�3��~��.����iaG����P��9�Ԛ&g�)x|c��S���X���d�J#B�<��NK��^I�� Ɓ[�������+s�K@����d���^m�-h]{c�5+3���*?t�����3�J�m�a��M� ���)>��4���?t�a� �y��������r�0���e�>���OhZ���x{�N��n�0=;�B�^U���Zg9P��o ߡb��U�5ǔ *$�:TK�,Ç�d����6�<9�@_]<ω���xHǎ]�]��@�����GB4�W����_>?��Է?��O;4�S|�13��c��f]�Q�����T��*[{ѐq���x�
��/*=��=����Z�����em�Հ��%/�G^ڞ�ʧ�W,�;q3U�k�C���4�5� �F�`�DX�D�N�B{r��D��c�����ZN\��v�ԅq`-�z�{��/�륶ү=='>0s�� b�M������O���|s6� �3��7	���ШFEG1�u��Fl�����8 �q����sZ�TSBX)����V�rc[���Hɢ\��񑑶����8-�)��7�=%S�	�ܦNp�g��2������T6X`�iQR轹k(�Oq:�����M���"d���Û�
�������<K��R(ٱZc5<�.rJ�Mn#i�v6�M=jB���J?��;}{��bs��S-�^זZ���0��D�v��ec��\H{p{�t�j�0�U=v��lH5�e�����0N	����8��M6'f��b�]�%�:\,��D����^�6E�ȋ�7��8�.�03<���j}�}3/�jV�}8��݅�̡�r��ɧ�g��[�75KeN/=�\�B�ʢ�C}��g��4�F�	D�ڞb�0�	����[�\:}U�$)w�`���t<_P�-Mؔ�K�����O�3<"N�*b�~K��9,<�����4��!��NN�^*]��*�%vʙB"��q-*x��vA+@�Od��Y������u����NseC��"��Ue�����x
7�î_&�&
P5;^�_Q�id$�*%��#����70���q�nU��+�́x�(�R�K`��aTn,嵷�1T���]�p��e�p	P��WeJݶ�_EY"�u-��OI���
?\���S�[`��w�o9h��AK��f{����4M�#�����a��KO:ى�z{�su�r�,��%"Ր#�Iם�k�v��
;���z8Ql��w�fY��{f�� J��qV���G��,�>nj"����$\�D�
C>iKR�ܥ邂x�9�X���7�9E���1��sR�g1��P�h�$Q�	(�kY!�P`�|ݷg8m}kA��"��¹V,!����x�O
�^����`#H��<^��������5�=j>y�3ҢXw���q���`�A���W�D��$�禕{EC��aC �V�P������)8*$H� TWv��fP����)5�WQ�{w�YҷBA�!��x�0��-<���1~^j���bof��jg�!��|l��5�*[�$�;����o�{�W޵�ڑ���a�bݺqg��J�]��9�`����p��R[{�D��w����L^����6׃�X�3F��~�� ��E����l�W�;��5���L��~�75A��������t��q�ѯF9�%u{-�U7հ��ذ?`B�lZW��#��%Aɛ�;�spa��iP���6��}��FW6D�����״�
������K���.���*��*�h%���

�_X^��g,�������\4�]r��gv��ے�׀P䍟ي� �̘
�qah��&��~_jB�Xo���R�s���Y���f���9�9���6���c)In�?y7g����i�MQ 5դn�C{�Eȿ��;Խ����F�h��}ubp`7�;�����'�p𪬳��nv����+���	^�����������2u�GIEE���Q����Y"�ӕ��:��|Z[������2k]`a�f��w��駈�q�!��|e�t�E�T-��m���������S ��"y��tĂ9�S��r�\V�e��:@"I���� X!�
��n�����ʰ1?-y�KU�uH�8/�<�0����)�#ʹ�lîA®R�t���MB��[h����o�đ�[�%��q�ܙ��F��'C��2���_[uPf@�2��{�\��s��w��H����f]z�_'A9����g:v�`I^c�*�#��6�#$�3��-o�P���TPr��m�#��`�S�:�����_��׈KY�/͇��Zj��_Ӟ�6���e��q1\jq	qE�iU��iku0�'a��|�����aM�z)M�H��toȻ>���>;rV䬭T�t������M��Yop�<�(AK��5��P��?J ����������|k�f6��Q��3�ᓜ����.� �{?7��Ѻ̔ח^h�|y�Q�v�D������&2����Bv�,� �����Y#8\cVxO9.��'(6�d�bm��n��	��{>Z���w��ԜbZ/��ʠrc��w)'��Єp+J�1+�>�11�S�a}���b3�D|c��`Tc�`����¼QAOY�~9�R6(/sb���f8%D3K��v�S�� X�Ǭ��қ
�k�P�����jf	4���fR{D�uoq(���}^�v��cd�צ�_�������!�y�\Z��|/�:�9�Ӷ�dۭ��)ao�9hFw��dP� �<7g����g���'���C�#L�t�1�C�������Qs�s�w���]2?��I	 ��j2�����AN�^܄i�T���h�\��.e����@��U� L� �KXhG8on���>�����6�����;!���᪥���X���`p|§�iUx0:�v���k���~u�e��M��iR�mK�Ef`��Zxn'81&O��u�M�&����M��"�e
�؆uIR-ls(
!��H���j�쐜T��G��Wb�|lΔ�z`P�W���1���u�B��i�p��{Q������5����e�{�6��m�b����
&x�����'o���X;Q��1����0%�F!�~}�����_r��S-�T�����a�<�pYp�,�sd(�-(��	`q�>B�Sv���K��$V�0	s��3
±(A�.�D(����6XJG'��{k����>��[<b���h I�Ж���/���iA����Hg쨸��� R�w#pKHڔ+���vd�[����߽�c���>o��f�zk����]a�A-��d-ӈ�t�P�Д�"������B^s���eT��v�=$I[נٝNkOt�X�q�
��%v���]���z�N��L�-��FQum�ֵ9������N���	ڛ�3F�]̟S���9_v�3��#\/�|.��b�+ ʔ~�����J��v{�m�1�e�,V
 &�$�ńla����Q!l2d�U5�J���Ԋʕ�����I��P��h�|��ש)�K�u���#u�8L�$��]S����|�Ƽ�T���dK9f����sQsK�mTdwp�G��~�
�d506��a�[���n�hR;�gyN�BD�>O�6;��ׯJ�28�Or�������} 0�B�٠�����G�5�9�.o �>�z�}�ǣj�Mi���O5JN(��oB�"���@�ҫ��b�<�r�T��E(_bm x9�d��{ݒ+��&�b�Y{QK�ٝ/z����̀}[�oV��7�����Ox)@�O曇J]�X�?�Z��9�`e��5i�������5����$�G��	�8��˰�At���p���9��;���a��K�����!�Wr0�B�ځ,
̝Jj�_��юI���<=���p)��)-^o|�^i[���dE/���Ъ�XoY�3��a��K���l	L���+��4��D�}~̀!�o�O�>�T�$�
?͝�&�И/q&�I.9J�?���yD�y�R�6�T� <��8�@o�V�oģ���z�X^��c����A��jq�{�:�0��d)�ǌەջ�D)(Wa���u�!�ps^m-���\`Ӭ�q��!�L׾���d韁����OX[�sr��<)f����-�%���TB��U��Q��f�	��X�ݖ�����dIcE5!���;����W��S��"���.��;���#�/��fͱA��	���P�Gע���)X57XGNt-�t8@�j��h��:?����i�����jw�g�^�����_O��	��a#@�
�nlISV�N<.
NR"q�i�T��$�W��[�yx�TYa.(�jҜ��kll�83��sNid�0B1A�~ ?"|^�]F�ӚߖLDs ��e �Q�ghL��n��8�8�K���n<MY,�B��,�D�/���[i��EQvK'���p�ۗ-ů�+hl��i�|z������2d�1��G'9$�^>xN��Cj���(�##���]<(����=�w�� *�{-��mi�j��\u��o�Ut��A�7�9<�@wym�;�K�z�:�{�pӗX}q�֫����z��n�<t�q@-62�=�f�k)J��X�`S�f�y>x�̤��&e	��%r�s�=�鵇�8a}	[P�����+?��l��,CX7��t#o�`ш!�3E�n��M�pp"qgV�8pN�Lf�����I>G��,l2k�l�����oZ�I���/1$_F�ȗ�����i�^�������2����;J�v)�r�P蒯,S�Iv�Wr�׶����X@xm��L��Ϊ�m��՞Lv�SH�������}�J�6rPqG3������L��_y���D����A��d��f�����h������Q�3��ېZxR����%1*أw��1��Z�GT6ڨf��EU�ƞv�4�Z2��;[���sD��y������#����Tt�U�G�|Q����gL�K��$,�V�o�/G5x9jk�>'+�^rN�$�e�.�ɻ�a�{�,̱ulrR9Ũ+��}0�')!ݾ$PwF�ܾxYF^;F�\ʇ��ou>�OR-��9�i=Ȩ����q���,��^4�I��G��|�\��6#RE�+=���~�B������ʹ�II��QG�(�n��mh�!Z��(�ϋT!����r/�AF9C�����i�8���� ���^��.Op#=I�
[���g�,9�>��,\����{�XD���9d*} ��0o��&M�nr�����q�*!�UAN?9�n>@��k��� �X�և3�m���J �k�B@r:�!�x�/��[�-���4�C�	 ( ����RY������e��M����R�~�8W��}��ʺ���9a��~f儞x����3w�~[k�3�s�"ƃ�6�k�U�(�'zzB�i�ju??����S��pe��4̠#�T�A���b
������]��]Hl�{���ɿ4y�ۻ���e2-�յ�$&	j4������J��B����� �',{�RP���8Zb\"pc���d���\D��� �H�:��ǡ���Ϟ���m�A7���������l$O2U���A`���@�C��紬eQ��_(#?������^��\>ǟY5fw�͛,������⋴�31��y����ɳ�Kq\G��ȏG|/������u�7�φO��s�U��m_Hc����ȹ��D(�����rv0Wn��I�>�y]����57�q.����N:%w�V��Nch�f!���KT`��a�i���}���K	(_^�f���zh��=l�L�U�3:��&@(��O<�L:lq�k��fj��N�^�D�q|�N�	H�ov�E|k�{� T�@�?��X�m�߂�W�NP�`�y��Ȝmj}|��r��3�$��U�W	^k�	A�p6Ι��G�UП�$�<{�F��UC3۠g-��lU���β�'J�4�=s:������:��V<�Խ|k�M��f���5�+�|m&r�	q�P�x[2�㣚W�M�4�v�My.�h��A�U��?�^�jfc��?�8@ 	��nLWnCL��؅��7cb@�2�Ҩ��=��s����Y���a�TCu���2M-���TM�
۷ Iރ��i
�}Z;���Dj�(^ak�
��+p�,��)R����)�S�@����r����32�W惙Q�w"F�zOR?���ψ0[Q�FW�����4��	���q��m�'�q���T|R�H���V=�u 1��~
��ƸJbTg
t(td������Le�=�o��߇��������-�O�B׉dXnۮ�WrŘO��K��/�]�?yD���ON�x����V�+�m��BdMaV�Ʃ+:N���v��F�Ȋ/�4����cϤ�S�eN�NR�Ⱥ�;��_��]@�6���hԣ�&���ʻ{�Z�}�����.�E���PM��c{c׮�$@�Z1��h������E�$cKu�\]�2(P�?;2�F)}�� ����X��G�7�M,lXV> $��S��b�}tX�K�B]Ǥ��/�b�Ex�Wگ��>  ���J�	A����Su�=����n/�W��_�s�i�#�P��#j��h�?�XM�0��C�c,Xk�.�ƅ���G�E��xk\�֩�$MD��MQϘP��bt״�����iRQd��SdG�n�x���[�J�q��Q�t�` Z.��}UHr�ϏM�A�/01�@v���;F�
�00�w"���k���� +�M����2���V�8��,* )=�߄V~���v4I7�����o��	���3	�I�/��ĸ�NϷX�
_:�A�'��y{d1�A|�����ҀAr�lMO�Lm)�e�@Tܽ������{g�t�I�W�E�m�6u[i�� s���)R�,}q�T�ն#L��u���w�tt�";�z�g�@��9�U�=ؠ5��l��U��i�ܞ���>3�����)J	�Z�>̞�C]�u������=ʕ�&{�N��]p�Ľ�V��%t{�!7�Rm��Y{�_oS��:wiN>DZ��#Á�*����z�+�D�b��!t���+\K)���2��:�?��F^"���bUY�����9Ԯq)�K(ꉤ����'�Ҏ�$´�cxV���.�+�p�G��pcV>�)X�z�\[��z�?�ZY���Á�[��m"�}|�����L����M�ݼ7��ͼq֚� i��h���$������a/.�{�^��ot>M����k3��N������Q�P{~��	��: �$�cd��)�b�p4�rh�w������QpG\n��ƃ��ؐ�ݖ���pD����fh�h^�'�:�*���9_;���ڈ�M0P��[�Jx~�ҍ��w��;�����{�ko�3Q�z#�\y�{0�α���.�Z������^yw�7�n&�;,��+��`3O��R�2�d,�l�^d��K]烘��$B���0_�X��]�!�E�깸��0 �6�7X�!���"`i�#��?á:@��"��a�-.z����ל��Z=���˾��D�&�Y�oѸW���04}�I\��ꔌ�
X�imj3ϖ�m��k��j`�v�)g������W�]G`u�roBiP՘>7����gA�zGS����W݂҃0�1`��e����0�@���Y��8ΪTLL?t��?��Հ�Oh7����MG��Wn��@퇓�5ɕ.K�y��)��@o�6�M7y��V���y�4sr,-�U<Q	������6ݕ Ӛ��Ϯ�3?-F��R�q��'�?p
�g���Ŝ\�+�.��1~�����D��I�{�8F|�V���u�'j{�}�hv%����g��i���u��-&}ujm���7XJ�`|��l�n3:���,4�s����Q�/�!�|��C�,&9!@�[y����>���,ŵ�����PF�H�8תa�F� ��*D\K�3\�CR'W{D����\7��B��)����߅�~��V��wPy�؁��6W,\/�eJX�zʎ'�O��xz���ЍG�?��E�N;}��,�a��#	��U�.6n���/�u�}Ȫ��bOe���`�F W��9���;�S7�i������<��ul���V��+?��v��q���I�w���,S
�%�M��3�툁�T�y�S/FƦ	���!-�ͱ��W��BM`5�J���gߊT��n�2��8�N�����jV$)�y��$������z���s�a�k�!�+l�X���\�ͳ8"���O�~���G�c��2`�#}\`����%�&7�4�V�9T�B�s�ƄO��]QO|�#NCgI[x����O��EM0�� eE�*��B�.u�OL�gP�q�n����Q��f%:z�{�eG2j�����N>�g�����~<��4%3�6��e�7�vj�ӫ�:������aFŹ71[��I�h¦���(�;-�%��9eҿA�<K��	^�������������Y\���_Ψ��Wo�	���.�(�O��u.C���JWI���m
�h}�ﱺ��-������}H#���+�*����*��c�3�a�L���QC۽����QV3[mQ�ޱ4��	
��F��� �nVV-�0rj�t�㋷UI=�ճ�py�6& �F�hmȱ�K�s�N~�E�,
.�s�a֫��D�FJV��Wx�b�7Bf�]]S���7 �"քduN�zW��cͭ�>�-�e�|a���'��R;v4�	���@�1���/�)�����P��㠺O��Q�A�܃`�U��(������n��_�5�7���I�Csߠ};ۉ 0*$�_���<�<6s�p��[h�cfɠ��&�' ����%����<d+�ΐ~��1��^�ԹD��c�JRg�b�]��g��Ev�5�l�R�PHCG0=���R�޲(���o|����A]���Q�C{
�(&$�9
X�nzx�/D�`S��t�p�i�7���I��Gt)��kUKi���kғ4�	l?WQ_�9���VQ�r�DIޯk;eA����!��Oy ��W+O�� ��pEh8~!�Q�j�>������^��V�?�&�X ��\�UZ9�4���[L����a
A���S!�	<�dF4���_�׼��M@�9�A�D��u�e���[L�;d�c�<ps=P���t��<�r7Qn�d5���J�F�r�?چ5�D���Z����$*��m �<+0��7��oxtu��S*�TSg;V��KeB��i����߱u�2n�F�e�;���:j�D�m�Qy��-8j�B)��|k�L^��ۖ^�)X�� �i�$��@�!�Z=���� EK�<��%�U`fLbj=����M;���,*��W*�����: �ه��{��t�1l��
�JB�ET�t�΢��Av7R�Gl*� ����kO�|����ڊ��q0������|�8*��s돨��?nM�c�d]'����ǆ_,�vM)� ��X>_�#�p��+HD�,��E��������J�D�Vi8����@r�ۀ?z�A�o��L���v���F�����|���p����,,%�OZ������'썦����C�|Ժ(:Q� <dq�S���Ǔ�w6�����r�-��:]��]��M��bQ�-� �,��Z�SDHޱ)��\�nK���ҹ���&��-�'�LQh�l%pIôCU;t?.Z�fpi�_8A���T��6�O���-�]�"��&��}E��C�ɱ���3��`���߬�t�]9>M��O�����l)�9�"v���$S�q{�=*j;e�#߃���I�܋�/E�?i����I������r\cB�÷�\
�F��= m�F��[p0�C�F�M����;��R�\j;�����`��P�0��f ����}�jI9��w
�g9V$����P=�O}�'5��_�8:E���0����u�;�Xز��*���O^����F�-��3�^�]#�6�f���'7�P9���Pc��_V��ڪ.ՆAK�GmQS�"�5�g���f��L��G��h�7�8�.�?d�-���0��bT&,���eB��Y�O�1�?q��������ٞ7<�FNЛ`Z��X�I����z%v|��EZiV���S7�O�}m��"���Tk� Y\�	v/V�G��+n?��':�]�;����d���#�L�4"7�ZBpQ�mya�GJ��SC��n���\�E�@=��hG.�=���d'W��q������+.�������죅j'��#�3��m������Q)�1g�1@����bj*����BRE���G�I0�9uH��8��WQ��ۂ���� ����膇�.g��gj�C���tM�F�3��-���Ʒ�j^�%���Ko�k"�<h
����umC�I6�o��	��Y/~d_v����OK���磔X�����٭-��ȕ��e��~4��LHss���9}w\/ǕF$�A��f��?T�/l�>+����o���&������,��CG�v����Q�U ܮ,�z�%��#Z���;ؼ�W�� ���L��2�7O��	�.�,DS%+�OÐ<�~��ʅ��Q�4�y-������Y@h��ߚ-�k��H����|�媉<����ü����ߖ�cpA�@x���>1i�\�����pݩ(:���WҐ'{�$�h�kRF7�;Oʵ�������s �ʫe�������� �d��4)��4��@Q���%O�#�5����4vMq�J�5�'˅P�y������=S4Z���.Q����;��.4��"9Y]�mAPJl�{a��p�2H��N:.���~����j�����N�~Z,U��F�A4uu���q{�i/q)Z�UOu�O,�S��Al����ڹ�&��Tav�,���0��=�����~H��ޛ5N˷�X�=�)�_b8 �f���#D��P�E��x��dG��o��߸���\�&��=�َ��#'=����})WI/��=ܙ�1s�����iT����K��eц�}�o0����_1��P�Q��0�����e�(�tV�i_Ne��~����Q�z���VPlrM�d�EH���#�����/7�X�i�qx&���նY�k��,��;�vV�bZ��X�0��3����-*3Y�wZ�N���1�&ng����9�/+3vB�%���,"l�~_q���qQo�t�7[��PǺ��(dA��uӕ8=X~�M����;u�Y���r���H����u������f�0yi�u�_��C%d%�'3ɘv�ݘfM�`5�T<�Eܟ��n���֐m0?�7�`�t���T��5��_�H�d|H�������Ǧƿ7���(��˯A��$s�3l�d��!�[�nŲ�G��,�ēt�e�CO�C��ͥ�5�"���J?�����>lU�h:۶�J=�ܙ�p�7�/XW���!t�'Ϩ�n��u}���,a�B*.�l�o���35:+�}����7bP�%.����x��3���0.��}�'�';���a��q���T6��5]�Xc;W[��+T@�r�M��˹� �{�򿶄.Ã�Bv��A�E�����EY�&��d�r��Q�f��&y�!.�j7a��Q:����R��ʻT0�"�LϿ��d�3؛<���m�W�I�{p�E� GR��G�����j
ɉ�d�2�c}�c��"+����H�g:gٰ
O�K�U�_�vM�S��]����+����ys���[ʼ����=C6c�kEz�5͏��s�����FT;���墍a޹}h�U$k�᪌
���{��EUZ�'y�DB�$6zlR��	(aά;�w�P5���^/DU8���t�������}e��uח��p�q��i\��V�t|�QDl�>�����ٜ�B&9���p7�8��O+o�T��,���hkx��g���s�����?h�n���D��Ӻ�-]e�BNf��(�=�����^zۆ3ZOJ�����:f�D�rC�Xf���-�I��H�& �z�FJ(���lq��p~�G��VIR�&�!CE]E>>�Y-��}���F�W�A=1�kR����xd����u�c�M��i������i?0eH���dna�����ch�=�C?|"�zbB7<A��<*'g���o	`U#���6��JD�G��h��N��r�,y�\Ȼ��/l�dJz��䭗���ؤbEQ��=$�Ec�uc�� <f��[����f��ʞҺD�k]@��Rb�^���ͪ���G�����W���%7rἇ�<ׯ��F��Jy�{̺��|t���MN�o�Y��	a\���'�@JYe�����L��cI�V�^�9�Q�F�tf�+�To�����vT���So�ė6��,�	HTQ�[o�Fr|�h��y\� o�W_��j��*�C�&��Y�������=�&!�-���4�n+t�6�m0�4�A�-�p<�����Jۛ�k�!nd�B�_���|������׭b�Y��z<B`a�^�@�� ����H�/��qϷΓ�b?��]
���y�2Kg'y�B�E�\�:S;(lY��Y��e-.�Q!Zȡ9�l�u+i�Y�To�g�������z[�����c9���R㍩��l�6U��!��[�;D��.�o��m@��!R�!e;
ݓ ����O��bڬP� ୅d�B9�l�1�2�l��/4 ��������!�����Uy�#��U�σv/�.G6�6d��	�Y:>���6 ��qtc�����u�S<,�n͹�Bh�m�O{�a?��Uq�����]8za�sug�/���P���ru��ɔ��&�
�'
���Q�{�{��ZI�~��J�*��5�=
x9_B��z���8+�+�����h����x�I������C0K-���u[��I>����~�����̞P��Z���Qġ�p5$����芾/$]��-��UH -��aɷ.K�s��64 �}�������t0����˜%Wfŗ5Ҹ��r�S>I1��}����L�{�@�^��*�f֜B�v�'������:2`,���z�zz�>��F�Ij�/�=�{c4��\.�\���ˏ�p���b T�=�>�IΒ�z��x�#��/��"w�L�E&O�O�r��9��Ǚ�9�4�L� ��ؔ��&V�~�	�T��0��r�sHio�����|`���6xK�جv�;Oh;!n\�qS��E�T��� *¼��=���4���������향ra�L�X܈����=���43�%V��:D%Je6Iێ@��ho�/�ӛ��C��-M�%�$�o���},VJ���W�(W*E�薀�����y�v��u�U��d�F/�^��
��U���"���� a1��l�x�;`h�%�PS�F8����$����M��]�3_���Y��%����ӊ'��>��Y%�� h�y���gӊ0/�H�"��pz]L7D3�����P��}�	7{{��-
���ߤ����,cJȨ��0��fv��Z<�M��A=��h�/KM�����8�o,�P�x�@���y|�u�6bѠo꓈	f�0"��0��iP��l���Y	���
�.��<a�B��{^)\k6O�����#A%1!�Eu��_ӛ�K�<����7&k[�M�H��z�:r������e5k� 6��>��0��Z`7����[0������i�/%|yk�R5��$��Q��3t�S�[F�Q@*ay�}
�ھ�6ѩ�QAf{:�K�n[��XN,\����X�52�N����4st�R$�ݍk�3��$�wz��BF�!P�f�!`m:����K�,wb��V�7�#.�� 8�(��W6��5����?�����y�f�מ���T<Tv�+�`��"���ŉ��rW͵'5����2�SM��@͵��1�& ߇̥��t<�Zو7����c�fkh
*�p�7�N�O�'�G2��,����/�}�b(���6��y�W���s��G�Z������s_Y2�����ip��1d3_�kY�N���=:)  ��C;�O�~X�)p��y��gˤ���e~��0r�;�k3$H���� ����i����c�	��F8�J��3�h6j�T������>L����ײO���|���D�ě+��2�z�e�cAWM���Z�_�q��
��	p�k8�ؚl�	�>���J<���K���q޸��f��_Fh`�s�<7-b:d>�0P����T�!aJ��{�x�m����T6F�o��ۨ�6�H��=�מ��boRW��Qۚ��'?��6�F���/g֏�6�X�˩�>u�&C�<a�T�t�t���uP��볋�}WdN��կ�м\�x�1��S҆����2��H�OP
F��Ʋ���11dQe=�F@�#��6�Q�~a�A>*wS���	��_Or�%�~"r���r4�l�2g~�!��W?o��"��-q懚o�ы|��Wv��
���Z��/�p*��X�j,�Yk�ҥ��!w��ZK�;\dyhzÕ��rw�Ε�����8/�3<?|$��=��
u�=-Wc�)� +����q�w���+�LY���ML���~�V���0�r��6����8_8}��Z�s@���D�]��,|4A%�gTTuuo��.褹wJ��ΰ Wk���O�픣3��c~%�`���<�rj^�x����l$��@Ȧ_o�9�p�Y��Ɨ�o:ge/G�X�0t(����ޣm��=Սѓ�I�^I7z�T�O�p�󼺘3P,:.�CmN ��^�՟}����������C���K�ŭN�H�S�㛆/o�g�.�(&2Qf�5�P�B��E��6i�`�i�q�7�8����o�ܭ��C+lΠ�)�g:�B�N�%�s	�]яǒ��`�9� 	��gXd�C��I��ݓ0�m��������'8��dz��fϨ�}{�xa�
3BHX��+�R�6��6�H�_�����g���?0�y�m�+t �ѦHz�F��Z���d�i��{U*���J�?V��h$U��
��y5�0��,"�C�~5�����1~q���Z(�rU'2�B �
@�zfQmS1.:��o����19����4��*�T�j&C���=Fx�<���.�RV�(@�Z.�����
�ށ�j��6�H_(���-B�Q	'xp��P<�"��IC��%���[�҉�D������Ov���g������
�v�h�rM�15S�ha��2��s{��6Q�Ix,O�A9o�V�(�yw%a|��sA�Vɬ+����Xv�7�˗��g5�����1v
_�dV�q%�3����CeN�9H�����d��� ��v6B߸��A \���4W]�^l�#wG�H�"@�c@���i)Oc��`����0�'����H\is6�����A�'�A��H�C3o� Eۂ���x��������u"���_6��?i�������L���]�� Ť �h-o�pr�S��i_���j( ՎP����c>`f�0���=>\-���o�i�� Z( C���(�Bw��Ԓ~�J�%�y�ć^�M�7�"v�@GV��WW���h/�P�
S�	�T�D���H���%<;�X�m����5=�Њ����)�����c*p3�>���T!�*M��>9囒׼��#��(�\��?c�;���fohc^W�0p���>�_iמ��o��$t�S=]őId�;j���Z3L�-�*A�3���OE�	Z<���-#*�<����X��N1�6�+�|jLVU�@L/՞����ʧ����5s�*�ϡ�ݐ��+�r��\����CK���T�.�#����t�t�܋�n/o���U�}`U~	J2�5��0�:K�|Ļ!HDN�탬ԉP�d�Sйf<7!��H;4?��n��Q��d�q�$�	�~�rG?~�&�ǠO';ɬ~��c�����rɈ����+aA�K�h��y�>vmCe�e��vK�#��i��{������Tz/��1�t`�i�Ֆ$�g��ꐊ�㛮|6s7P�r��%G�_��@PGl���G��ͮ#��N������_�t����E�12;QP��A<��~$U����|iԵQd�wW�|ᰟ���h��#��y��g"xb��5=��B��U�<H���p_Yi�"�q�ʔu�	7��8ϕL�S����W۶˟xS�8�c��?'��� R�x�X���̗R-�ي�F�Y�	![���A��5[SϺ")]�EБ�IQ���YQ!�ơ��Ic7�k�����J������An~DE��ꅧ(��W��@4~k1ڂ��U���,�d��ױ����rZ}#<ާ�a�Q�x�.'$���t�$w��0S�P��i����1"	y!-��|�6cՇ�����
s�K|<T$���[�ޅ!%�ħ�4?g���C�~ū����:'y�1�+�x��~�����f0�	I��ly~t |cSb����ȶTN �y�����C˚�m8��'�-5EFX������cL���EԼn��aJ�������z���f|�^�/�тˢ$�$J��������.{ ��pT�:�t9ãMP ��Y��G�Ir��@/�A�V����N\{�V�9q��7(�=�]��X஠�;���wg yp�������M ��hB1����K����'�E��МUqX�C��ݾ��;l��br8�yW�Ki��U{���Ӂy�ZW�|�d�1;�vA	 /vN��۾��_�+qr*�� ��C���ibO~��K��1a������Ѐ�
�H����+D�f�3��2B�2�N��n�C�:I$j"��e���
Xr�����mj���6P��R��C.�?k�B{���P���������Ң\<L��bJH7ۄ*^F��91 ዼ�H���������T0��`6"9)��r���pH�Lz`��D�+�.�Pd�Ҹ��5��->����D\��!�q�Y�*�/�H����۳E�1�(�ok�������q�[�6"P֩��>�B.�������:=&#(�m&����nb�WAiܼm���ʿK�Դ_�W�Wߩ�N/�,t2T�B98^Uue���ӟ0���/���6��ǎ0˰��H�;}���/XxE>���Y�����,�o!�70�Á *17�)��M���(K+��Y��M����F<NM��������]heCM>s�y�[�PVL�,0�R�Z���YG�,nF-���ZVeN��dO�N���G���f�$W�2��1����C���Qp�jE��Ku\��t�����'Aא�]�mm���=���H��ʊ�e)��Uwq�ɤ�na8v�vk�t9*X铷%���U���>+��q_���[���������Y9�����e!�él���GF�{19sڽ��rW-�J�ҁ4�=ĀٛW��,�U�`��)c�VbMp2�?�GB��f��M<�'!$�����_~�Z�}C(1�hu-�%jGg�p�i<�X43G��Q��B�o���"���]�:�/Ug�.KLh��q}Y�¹(Ṳg ���R7��()�߱ZDg$����� �&���@-+[��\�-�;$֧�	�b�N}��~�>����7,�{��{��k��C�aKZ�1���?"wJ/@鸓PVB���{��\��HV(@?ݔ��n�8r���'�|e
�Y�3�=��gP���3suԍ�)�b~]�K�7�%RLU���~1����|�-*��Q�|S����3�QA,���+Η�9El�:�B���p�8dx�������_���n||�|�u�SV��_{/C&�u���B����3D�
:I�@�(������^�48�Z.�Z������t���;5*J��;3��UXSF�XP���' ���E<q����W�]Ge�}�`'��%��1�5Qmz��� p&���,�]gߑIS�Xqq~�8~���wYPg��6�8P� �d�VA�?�C��4�W"q��|�He�W�GN�Rt�j�Gp ;c"p���J, #׸��z�V�V����W�h�꒎ [_#}�a5뛗S�n*�]m�z����?�^�%��g�oX7 ���Y�b�۔�˕]
tY�{5�$-�~8:�2���aU������E�bOC�R�}�^�u�2#��@�~��M�Vc)�^��)4�����fɝV�W�<�4����rh��Iu�vc����i���=�	iõ���bH��%ӷ��y_���o�Ϫ�D_�GvX^M�R�+�8�gX�5J�SJ��p6g�m�XW��������x�� {�ݮ^,�^�5%CQ�����Ѯ��W)�,V�
���m���3�yP�sG����T��|o1�V�U90��{)��w����V�v�Y�'Y�55m�i}&������@�k�\�;��88R�V�e�
թ��g錢jb�%��Y�W��m�ksd�u�rK?i[Q&,ML���]� 8�0<=J]�"C��,a;�q]�;Js����aS����v��*q*u�Ŗ�K��L�^����U��
��J���Nª��h��Ma�~��^6DA8ĩx�A�4��봯`�@���#�8Mk|��aU$�I�#��e����?��[~��-"���9`d�%v!(X�@�<�7�N1���C���R��e��{]w>z�͂[����$v[j��Oʹ;�Rmc/Nr�b��b���u���o�=׭l��z.���z:˷@���>���+��3��9c�X�[A�-�6��=
�o�ei����?)��h9%,����`�3M1&?&���W&F��E	rI���"0��ʸ����	��fd	�@z˂5��EJٖJ�#�d������X�\���/�3�N��x�����"@�'o�c��Iq��������ݗ�B��Е�(��?��!��Qx�R�	j��?�5n
b�Kk�"�6��Se��M������k�·Ty� w�|�V��E�;�ƚ��7�Js��$�hSU�j!�PJ����V�в�e�F�P����$����� ��5|��l�ȶ� fw��W~Y`�Hňֲ��.5^��c�|��Е>Ea��ލ��Br�2t$��80�R]iX���헣MaD&\�F�|�1]]a�֧ĥ�W�ڱ���&v~�o�5N�L��5��BiҪiV˂p���V����f�O��L��3�Ty�Mw�Y�o��ħ��8��T&�HGM�I{e���@�ׅ�,�P�<�b�!#��{���@��u��
�
(F�y��l|���l���ق�˾�	i�8���)�jxU_��m�\�>/�:��2GK����(��+bG���9���[�0������3��%���pZ,Y���ʕ�|!os����$�?�;�lt&����Ue�^ڃ�]�����>���7��C{�o�f ��?��n[+��\Φ�՞#Ξ��y�����hf�E%&Ȗ<^���layX֓z�>�M���s���{�����zHl�z �x^�ګ���/Ă�z�%`���0{��M��S[�%6��֎kޗL�D N%���v�a"#�N�}���4��h4V-�2gJj�����4� ��ܧrv���XT]��m������t�vb?U�G<�V�kb|�X������߄+ Z�ys�W�ݺ��߹�i)�yYNu��1T��#�
�vS$����h�s��D�D[og9�"�.�Vx���5@(���t�]��P��ꕔ��~��]���(��i�$�q�ˀ��!���	q�Ѽn��-hS9�k� S8w���m�CQ;'��U�������t!e��?�]ti��N	�.U����绀�?�,�>�?p݁�ACHa�&��1���VI�M����
&F;����um��ۍx����}K�������jS��S�f{E��'Yv3רu����i�\2N�K#8�8�`VyX�IuY���&�T����/�n�8���z�� 3
;{DS��!'�6�g0L]])uy���L���5m��Q&[��MD�ඩ=Ά�w�#���<>��q7���\;])6�dg���O��w���4��$`"�:K�����+�'ܤH�ǹ�E(*���c�O��.0�:@+�D�][-�pE�u������/�m��N�ug�i�O/}ry�|��	�
�r[X�
�D.�{����L��)h�%���r��~!νC)��;s4I~)��h�@�A��)?�XN��E�4�+���?Z�q4>�-*p9�j���Rta�m*�#�Dn�L�w���o*��ޮa�f�e�2SV�V_]�EI��Sz�Z�i$w-#75y�YP��	������Sn��U�o(�P��;r2��S3�O&�_��U�ⲗ�\�9�H���@鴃����ll�3��+�O�n��`��y?96{������wj��%V��:�0��h�s��/6�e3~�i�`V1'���Ɉ���1^�CH�}�g4�l������,������ǗV���J���)m]~��U3c�%�p��4�݉?,(r����(�7��&F]����o]��CB���z&�	�z��^�c�ݘE�L�y?a�e�\����>j��dܬO:{aI�D�S���6��	~ȧ�����l������G�i���vʇ�_�A���G��R�~k�	��qU�՜ܘ���Hվ�yy�����R��T�!w�<>m�> %��=Hw7|n��"��~��Ř��i�e}�9�O�i�|5��z|JgK{�� ��D%#�������A1�|d�|��Tt�V��+�R��7��1�-<�.|�)�@�;l�!o��>��;�x��h��L��D7q`�ĥVz��tM�R�XCD��9Ky��.	&��;���w<3�A�˔�XTɭ�P��a�d�SΆ�@���o�Ӟ�H\i]/9�}�x����rm��1�OqC�����,Ꙋ8��y�Ƣ�u%3�V��s��LfѧM�@��Wx��M<�<�	;�%5�8��N^�~{:GQk������Ϋh��}*�j���d�@�3,�Zh�� ��'���`k��A����[�u�u����W[�U��@�:�|�|�E�)G��F���fCKA&���U܁�A%0p<��N��*Q�6������R2��\�9�A�!w���Nv�޹df-�$)�'���,��o�U�}2�S+.��P�Y�7e�`O�(vfI��5�蠇.�:f	��a_dR\���z�q�*�9N��<E;���ÖR��?�R)�[�h@�Z����,�lШQ�A���z����/+����<�t��������I�<t�z���n���~*|������� ��M%�i^�� �hL�����=aOB�ez{�]�x�!C�.P�]��u���8�F�϶���X��gt0h '��n��"�A������ oP�tDÑ]h�6��pn"�F�s5�*UzeD�^?�p�ХA�U��C��Zu�P�I���p�L�=y�	'��YÐc���,�O�;'��_@�X������o?�<���E`�����j�?y �&S�˿�����d��[���٘=K��Λ�g���8�U���3ۡ��W��M 0L�]����f�+�[�OgWo�e3}k�$N���Y���[�ZM�
+wn����}'w�-%�@�>�*HG��i��O��:�mW�o��O�	'�$q���k8ʚ�./�5�b�'�RHg"K�Q�L!ğj�4����d����٥3DN�:�b�nԙ4;�)Z��q�ڋ&���3�d�#��WO4�d��.pw�C ��_;ԡ��Z�iIf�[,��Sf�ذ�l�h�B��04e،�x؜1�
����E��Ir�AMP޸��9���}�����l/�܅cوlV�x�,J���O~R�w{��]1��}�Y��7+�(F��i	Х!P�����dTHh�}�#q�!�G�^6�)ec�O�L��q�<��׾<&Y��T:Ѭ�.9݆]�+9]w�cq
6����|X�|]A70l��c�+��\�	�,EWy&��ڎ\Y��7���}�5媉u�f�m���v٣�����I�G�vS���bnB�*��C�.���9���݊\U�wZݚ3���y�f`�|�/���
װ	"�HL��1��U�=��������	Kَ�e��jx�.�z8���M]E>��v�
 `w���|P�no���h����<�#�`���h�|�.�s�W����ы�g%�A~U,Ƭk!�3�j��F�d+��©�;��.�� ӱy��~�DLӦ����-@k��S
V��Gk����Jf�b�q^����|VSV��%lw��K�:��"��D5�q�'��#���^��p�1�Љ"�0��gJ(��W�tʔ�V��Xo�-pԺ���# {���c�F�*�2�ӧ������Dm-)T_UM����D��|*�3�%'���1��]b�(�Л�^T&�2�[d�#� e�UBW}�m����b_qk瘡�(l�����]k�4Aϼ-����Iß�m�GM�}P�u)q����,�� KѺ���1��)ŏꉱ�X�F�~��-`:��^i������-��g����oݵ��\7���y�EO�����c�&�G�W	�/���O�@�! ~�9�i�C�A���$�9�$î89|��2�. W[�'7� �	?��o�y��<u�9�}L�wk���>��	
�3`0r)q>���Z��@��a@G�cMJ�7�R��C� ��W����q3�����:K�L7��W�e]e�pM�z�������[��}������1M�}�R�g^Û$X�vP�q�Б�v>��j J_9r� ��0��Uۤd�^�oÕI8����ቬm��r�U
t�đBHpgF0Yw���X��֘mw��p�����t�b����~�`�V�Z6�d_�7BK�ɇ��j�)�� :�A(=W���GS; �DB�:��O���Q�w/bY���GĶ��������航{٫��6'ॳl3�_>
V������Ҏ��S5f��5ݬǲM��d#�
���n�*�P�M:["�2�w_�G�p���/ܝ�A+���D{�7r�2�����#ג<�J����(�l���nht9���7_�@b�'�/P���rpè@2>0��`u�낶����Kҗp2��9�w|_��d.��^"z	�/�	o6���D���0����,�2�Y�U!o�d��@�����W�qe����D�+��(����򴧃�F����)��@�H@���*9��6�<._��'���iLN���Sm4�$���XL��EP��ص�?�L��>�.X�p:�IȂ�/�\?u�2���!�G��![O��`:����xt膖��|�twQy� џl� S(����,˯�~�]u{~=C�ӭs�0�I,g�B�P�iGR��}�)H<��BG���eD�Wî$�b���D�%E���a_��A�HMQ�I�\9U��-�Ψn�JYaO�� �Ί������ǍN$-�y��
|��<ь�3���7z�b�km�h�z�.��bw�	�{$������3g�0��>��4���V
*�A�.���*��\"�Uy"昒��q�Ϧ��v�d���g0��I�V���+�py�΃3�H�@��#n�OG�0��H�0��#��xNGa�:ۣ�9��y����nI�2=X0#,QaW8�-�8�^U:i���D�s"���t�Ԃ,]o�6���;/ŝ�U@��D�)�{���1<j��@?tO�z�
��t�ĩ?��~B���?92�����z98���K�KD��b�*�������R�E�:�f��؛i��z�
u�Bkb������G������:���WDW9�A�����6M�y��qU<�弙q����U,;2C1x9���d=�e�p����(Q��x�NI3���t�۴�c>�;V�u�ȿ�o�UQ�m�c�|��a��������_��#��~ߪ��Z�TK�#�����I�1H��Ê۲���l���u���>V�)������u��*�f׋���)�����/�Fh�]Cͭ��4,ܘtZ�<��eL�=h���(�Z�aߊ�>x��Yu<ϯ�-Y���g�D K�3	�'G�۴��3@B��4~����ⵛ�	�6lM��CC�؀���Y��M�%z�;�o��g\��z�r�߅�>_����e��kM:��ռ�
M�(X�A��(
 ��Te����F�N�By�Pp�p@=?%��8�8���������/��Nި�Ȟ����৯�2j~�Үa�)kA��_�'����_�"Ķ�Ñ6�%�>LeG���@gd�Yy�T�l��k� P�����녾ԡ�)BF�ؚ���cn��}{ai�r�����L�?f�T���?��Me���#�&�[+;��c��l:L�.4�j\��R}��p��_yA!h0��[=q ]�.��J�2}��R&�|99 ۻ�����[g�s-/d���A�w ␾��/��-Ȁ��%�
��b��I�lL$����2��c��7��R����S� h�D��NTDLBT!˒θ���f8�$���]��%H"���L��	�⩔�.��e�ޔ�M�uhBЯ��&��`�M!_��!7�K�^၏�8!��S��*�ڔ�\YX9&�ę$b ��mW�S�ӛ��-糡�sLm��0J	}´(�}�	ZEG���F�/��8|t	T�Г2�ۇK=���VG�����}��@�?yE^CR�APQ /"߿r�d�-T�2"�V�9�ao���V�zL�I�i���t�b��M�H�6
D���Uc��#��A�g��mOܴ�^�o���g_����Je]&hI���((�$��~�۪P��F% }a�0k'S����� 7Ff����:�M���A-뗓��:� l�mU��D���96����.��=��2���t�k�ҏ�-ۥ�C?�%�������`�*Ns�V(9����I�4�`�`c�V�Φ�<�o�t�	�EL���m&�h���/��-;ѝ�������	
V��%�I��&�%zJ+����J��k��`Yl��b��a�Oי��I
G@��Џ���o�vs[~/=�p*�i$eR� h��~����8�q�~����K��1�H��;������ �{"͢����dƼ�~���n���w%�6��"�us���F�j���Xr��L���W ���3�Gf�Q�̸������Z8~���c��4'�9�*f��J�	�e�u�L<MEĸt :����sü�����S����a�qi��W�ih��ԣG��:�~��J:s�Q�ZW�[��p�T�,��6����1C��K�)���t��e�ysK%�;և`q!��FI��l%�9�t���S�W�&J�nִ�N���z���P$�ٳ�j�<���|63���x1��x�x�?��(�0=�I�O�	�ǅ�:��=�L&n��ʽ �`�rdJ)�K>0]l�RQ�i��ϸH&�(�t�y5�Ke^B�'*��R৤T+9:����:\*s���	����Q���j4XT��i]Fڻ}Ԇ����ru�U�{$$� �G��9��Yz��-������O�k�)m�̵!8W��D�����Ͻ!�vQmX(uϣ�Q��@�ipR������=J:�
!н�bk<3JA`H���P!�b�@���:ݦ���������/�`�Yz�e�V�1U%^�S�Se�5�$/(z����W���Y��[�����u�1��Y���
&!��+��m�n;p��}Pe��ׯ"sX�uxJ�e���[/�j�q�~�~A�7Y��Q
:�H�#N�[g*l�a��#0���7���ٮ���r,T���g��,7<��
��C�]��R(H�[�:��'mJmCZd�)q�K�!�WM_	r�j�U@Y�>��ږ���V�uILCR�~�&���A�g¼@9�a'��y��S&=QM_���$�-�����h�P=�0LF0w?�&��ִ�[DD���kN���Ҹ�6�0��.��	s8pOL7T�$,��3��#D�8��� �n魂L��`Gyf��h�FWA�v �ĵ�c��el�oC0?ee�Ĩku]iA��Y��U�HN��>����ю��S���i�0"�V'?)+���m�˖W��"�h�����`G�$}�K"_#6cѱl���{�����+t�U��ޘi�q���7.�7�Ey*I	�LJ���i�c�A�9��9#�%|Z��^(bfi��P��_5N�S����T���zV�_�]�X�M���5'ĤU���F'�Np�chk&�˦3����3��c`c�a���R�H� ��{�S������?;�L��"U�#��ϗ�o��+��8�P�և�Ӟ���"��n	�bˀ�8#j�����sy`���%����&ƺ�����ާ
ߡHd�p>��]y�*��Ob�{d#F��e�2�B)e1���y�證-���
{�q�QW��ePQԄA
إ�X%��{�N��Ӌ&�?˿�J]fq!U{[��E��������*~nk�1��L�o�_�&6ӞU?�i������<�d�ȹ�T�nQ���[���1 u�߼<_�N�:���p���c汀^��%%�}e` ��SHf;S��h%�$�����v@�v=�ml
	��ڂ��W�qI��݈/v�Ig׿��ui
�q���E�D:�\A⏛P$EB Ch!9d��c�Q��x�ȴy���oۧ_����ù;7?ڸ��<qʾ��I��f �/����4v��������Xe����X���T�u��#�y��G��H�kZv1�|�V�OlS��#�[����\��ݕ� ��Q��g�I���/&���̲~ģ.�9�����cc���YB�w�l�<L���<X�4���k0�zu4�͝G�c�[�_tg7Yd��p��w�)�.v|t�E�ǿ��Z`# ���
e�+#u���/���2��'OmGLKd�$�S���?&�=-�~����ւ��y�]�P�ҳ����� ����'�V*�'�Y�*�Ś��f�'Pْ�U� v��#	K���2��s��_ю��x=�H5hw|-��;��)�T�NLo�#xM$]v�${�t9L@�T �E�޵����������K�{X����p�� ��;�A �W����d`���F=�󧒤b�`���-O�鏖�e��3�3bb�=��E�m�gߛ
l,M�Y�4s��o��K����z�ΛZ[����:0�����I�t>�S!�V�@��}�RDIDd��쑰d�C����A��2Ƽ�v1�*���?i��a"g�4�S�%HP)=��$�i�1�p��'z���+�2� �Zy^Br�u��c��lt��m�+�q��E�]�����J�����Q�\�[#L̻a3k�D!�<SEl�z��T2�����w*ދw�����1p����Yd�yc�N�d[X��;�0�zľ,��`<���N�# Fo�4��=i�©�GM����9X-�1޵�⩄�.,(ƾƧ������A^L#QWO�r��/�O�C��E]�����_~1���^��L�H�T�6�sd$6N>pt/���]�'��׵5���5H*�S��Ɗ��E�4K�;��xk]���l��%V�jΧȳii���ԩiAǈ��2�V�z��I�����4#�v�]*����'?a�����gC��d�A/��y)p`W�ѡ	'L3+=P-�?]�DZ�Uf}ߑ7%j��Wl�m��<�+G�P�ƿ������e��a��h$.`szX�$\P��W^�c�Y�bQ���y���[a��8����-���G20�᤯�L����u6m}5�fV��,��M.�^N��WTo�^z,i�����mX6-�c�/�Sft�\/�ňaۉ�`z��$����b������Y�D,��>#a�X��S�k��Ah&���O�U���j�ˆJUIBu��Kz�����un1�^��X�<�pf_���J@�Q�\)��&��T�C�HY����m�<Ħ�X:l���r��i�+%:�?;�2��O�5�g̲��QQ������c�h��߿���p<A�E��t��P����g\��;\��~r�+g�xJ�ˋ�5e�J\wj΍��*EW��n
�^r��R��)ڠtI�u`'�:b'r��G1�r��0^�!Þ֌�:O��Ef���D�ԛ���!	jwcC%j����Cn£wlݽ5�(b�mȱ� =����b2�
QP�S�S<�)5�|��n8��s�d1�X��u��۲�^�o?�:=
��J��:j>|���K���%�(�A0P����`.��Nv�7W�XS�V�9�/���bї-�sM1$r��M����q��#,1�݄X�e\��bv/k������ٲN���&�S��9�5q��h��P�d�`���ڤ�BW�.����S�hv����lBy�U}¬�o����S^n����Pp١�<�b{k�.�]�{����-hh�+��Y�G��+�F����P��ꬔ#w�u��T��"�Δ��eV��rZwM-Y�`D>�������к=�'�����A����w��೚�%g�Lq۴p�b֭	���7��a{��7��_)���)D��EY��9��8�]5:�A%6���)�����i���� "p0w����1Y����=�(a¢���h���x��-���й�"��N���M�T�{8��R�ذ	CS2��bަ�1u}?o��fY�����'��r��16���7�9��ht�#yց�c�`��GLo�4�i+��%lp�]|ԃ���j���W?=΀#�)���;{5E䝩ʃe�7:��v������H2b�0R���q�B`��od�ҫ��
+��3i 4����������L8��	+����T��y���ՠG�D�����}n3}kM{��Q_��r�cr�s�+uy�S8��YI��Z>��P�_��A&E0�
��|����A8YZ�����v!0k�����f�9g��	/�Y�P�4��������_�h��ᒕ�Y٬��!ﺏ��� ���H	�D�x������,t�O�-S��`��_�b)2`&�o��6�{�)�/!�����Λ���0�6
؏��Q9��w�	�1��<��Vw�1��o �Yxk+^<�ڶm7��#_�#�} ~t��j����[cL���g�t�q�m1��xj����p��M��D�<̬����⌧�V�+��:�>��C���}@�`���I�3�HO��	 ��²�'�=8��O�$��pƎ�c�٣=���l�j^�19�tx|���!�K2}5��c�U��wH�f2��K:&>w����~I��������v�R �oOٌ�
�����hR�nͳ<��2?	�)�Z���/���*�XC
;���[#~y޽'m�`���?��/~��*�����F���a���Tr�\L���B�	8>��X������3��\��8f�o,��@ui��3�+ٜ�4ʽ! ˜���^`�LD�i-���EN|��H8��!TZ��}�MsȌ��&OQ�W��{��\%q����"z��YlK����0�&WP��FЩ�ͳ��mF�Eő9e�|<C��罷9��B��(i��-�e��Z�v���o3�b��5�Pb��G�Z3����op����VPQ?�c�bVo�2��?l�����U�%����5��@���&]�����͕W@�$M=;Є���=��'{ٓ����=��x6ә��A����A��F胠�%��+�gR��s}F�VǾ+���ƕ����2y$8��՛��n��ϳt�"�#2�����t��Z�Y'u�����z���k�_Zᨫa�SΉ�f�~�����=d�q.n~p�6!e�0"�b!P<�V.���<��HnއĊ=���nz3x�9���od�解'#�����Z}k��^��"x��'Ĳ6@��4��/�V��w�6[P�#�/�~�C$�w�v
"��f5�������������޾J�����+���|��j��y�-.�����H8m�6�F�]�|&�'B\��A��7�+R���^k������h	j�q�0�D���pw����,�����#�n�a?I���O���w�k"�����_����<��i�Wv��t}ؒ�\�z ��l߭�^0�c���� �+e
ô�Ň.�:��b������Z]p��0/�T�aS�(�}�抰D���'��?�5�3�Mhs�Z},���� )�~i�LW���9�ǈ�m�Ɵ�M���.� ���AY������qjI�̶��S�IG��`Pׄ�a^�(eO�
�#@Ϫ�^c�Kr��f�Wa+y��#�vũ�c�.�,�+N��R�Qb(�����`�ob�l����Z��<����%�=^{��g����v�����Nl��0�� �?������ܖ`eӱںEM�5�<5Җ6��s�`ÎRto��&,�3���l�Z�Z����z��?�/5�����3ٰU7VA^�v�;@O�V�6?�y?A�����N�y�ۓ o�e%>���&��Gx�!�\����>k�vY����KF~�g&�&�/��Fϝ��yo�M���V(�)<��H(�����z�U���$������N-��/م�G���n�ov ���By�85�,����jt����~�#�irF'�P��C��E��Bz��<grc$����=��$/�l�z�o���WG��̱��F�����sF�oLE}��(��c�[Iw!Qr��?i�0\�<� ���ȵ3����9fN�b�)��Rv�o�`�[�[5���s��?ɀ�W�Ao¼��ȿ��)�����^���^�����T'��@l����(�z���z@���-)NU��lMn{]�����59I'�������e�7���M�n�����wQ��3���(*�	v�L���|��h����E��)T;�[i7�dN'�Nj�A�3/PF!ݿdds%N�R�s��ȈC��Ṹ�������p?3g2(�׉��.�roR�ؑe<�w�j�M��@Z��X���g�Y��T�QZ���Oe�����f~4^�6`�XY�S)d�N�NxC����|��hH!�j4$׍�e#�����4��B��P�h+{��e��t<���9`�U��G�� WI9�;�	�#c��DD0�I�SJ�$1��;齵�"5�.E�������d=`���r�5�50��_�t�@��+�pU�5˭�*fz{��y$��w�0���G1��ϟ�`b �=(�����dEmC	:��-����M��J����N��v�^���n}�`A��St*w	��Ɍ)G;��❋�%��<�oe�ۙ���/�����F�^�ou:�l6g^�A=k��+b��Z��7�ڪ>T'N7 �?�T�l��k�\��e�n���qac�k|}}�.W�\�lam��<���I�9[>�A[�n�ۋ��Po�Rs���T���k���g�~u�>hP�&¦�ʴ�*3���Ȗb{�
�P�b׋ņ*��Y�"��>��?Ҕ�J�q�tjNk`Z |��kX��uΥP���_�S	���
ڗ�lfE���"PD)���1�=�T�\alsrm՟�M���\^&?�j�8�	���X2���J!T*��U����3Kck :��3C��+�'��	
��Ļo�������u�8�V�w�"Z�H¤��M�T�
�}����x���֮�r�I���8���d[1���r8�H
�N�1�7���f�q%�5Eu2t���0k�m��#�i���j�뎒�@�kK$ۼ?f����x��.�6Ɇ��i|�ˋ�g*�@6��oҠ�U�/
���*pj}�YS�����!���\��A��9_մ8�V{9���8��N�&�!�q�E������@�Q-&�Ьj��I=kX������IǶ�^��;d-zh8�&���23��G��>7oB7�} Z�`���}ϣpx�"�fc0yK��ӟ��=՗u$���I���N�:g���\��Ǟ3��%~�ʈ����ߑ������ȀH\�4Ѫ3,r�Cڇ���|�<�[I-U�o鍅���?�&/'���J~KdE6���r��z���{s�'�ne��,q':��c����� |%N��;t�`4{�u�M		���ðk}S�&��_FEp�dѦkZ�c��{�R�� %d\��l������{�'��f�z�"�+(���b��n"��XP(E�* ��p���RKK\�M��+��+շ�0�����cR�Հ�W~�x̢�T���#��##ak$쀤��IZ��FHG�B�� "U�L~��{���5��bM�p��bg�أ	��ȸ�d�Kܣ""I\�u�.��?�p�Jj{�룝�R}�59�j��b/sFf[p����<�?EzgI]�)�$k(l��̾�j��@�j�h�L�G���Z���~�w�#g_���w����[>�D2jgz���T�Դ�Eգ�?���΄����=j�I�E}~�o�����6�SO�N�^m|Q���t1�$�#k_��u�b�� ����+��"7�����ְ�Ы��+l�B��Q���'�c�caۙ��D��d�(��ֱ������{-�bO��2�\�ia�+@��Se%�й��B++��; ��@?�w����j��mw��`	� d��s��,�1'�H�c~;R���bc嬫�u�O�5�9�o/������ ��JK%���9!���6�\SK�����+���
�X��J�<�T��~���x|1y�]��փ����js���Y�P����)M)���TI��G����Ȳ�Ԡ���%����&�e@<{�2��:��cd0��y]�y ���m���|����0�p�MU���[ۧzV�@�Q��K��ɴ��e��ܬ��y$��!�ͭ���`�<�uy@ѓ�.s�y���C4��Vԏ���u�X�Ïy�Au�bS#(+�0DA��q��A{��Y�Z�0y#=k-��n�T��o��V��ݵi����b��?���9lh�0��2<~X��6.���u7E��.j��7N�s�W�\�ϡ�`�ρ�yI��d�7�?�k�O��Sz+�o��go��`z��Q�A~�s�a�݇��)N����Bq 4w�jB;�q�;Ũ��?���ʩc��h\'�w&<u�wƨ&?��ƙ��Ѥ�Yc�L!+qĆ[�'����dQ~�T��oY����w+��,K�z_}߭��Rf^<�?;���`Y����A�����j!B�I$%�X��l1yO��e\�ը���$��v��v��q�P�d{�Mb�ǎ�fK�|�4?�*dpu�2�������v���gV�ǥ
�K�K�4
�W�F�dv�y,hy~Kq5��Wt��(2O���E��Q�v6-��L}St�L_@`� PE�Y����e*�l��bF��V�Fo
V�~|1��{B�S��I� ,���B#2�U9��<i�R�Rq�7��n��l�p�}���/�a����.�7"dX��_�u�,Ƽ	�j���ot'ݼC	@���^7�
L,������6Ó͖q�)@P�*/��:�c�)�V�*�+�#�:��N�.�B3DZ�Y�l�
�v�H*h�!�ACy�F���s���cEh�V�J�[8Sw�p�x��읒)!X}r�#��r+�}�sq�4(�]����'qˋ���J��]Ȼyk�y��c���Xː6����Q6��:�w�/(#����v�f�'�͔%OG���YW�,�G�7�����<�1=UZm� %��E������C�<w������H\(����IQn�Y�'���s���r���	Z@,F0�<��h��{�6iNW�pl��u^skМZE�61ry�9.-V��-�� �<���vG��<p�����;��(���7x;�1�WaJ>��=�8�oO�j6 ���a��!�fZ�2)�����঍!�ܟ"��w4M��[����`t��=�Ȫ�.%�?*�;(����U:����n �)���W3`��� ������cΠ��|�b��^4r4f�qꏔ�&�Y[��F�����z�Hj�?��uD+���ݲ��
w��^���Ɯ�l"�����%,�1�S�cWly/�ռ�!��O����t�����گQ.�u�г������K�l�:k3+7�?�I:�(�eH4fj_f���-�c�\�R������������C��n!|�@c��r����G����L�)ND.��({/�]A{:�Q�;m\U2c�H�Lhd{�P����%d�i�қ?E���P1�1�I��oq�Gb�^�2L��7@V�@�_�bU|���֣A+h/>��U�Lj�y�p0V��.{�;��[ھ���'m��W�"�E5E��^��5�y ���z�.�ge���i�Q���y��Of}�	AK~6#'�T�Ͳ�jK�O��:B�~zbD-��2���tz3��[���D��,���fJ�Ѐ���9"�*ڎ�2߱��'ws���m�t�"\쯟7*T���&W��ӣ��hy����^p3��|��9���[(��x���m�U��|K�F��?R�\%��L���B^���{ӊ��"�Ra���zΗ
?�&B�4A�_u"%��=cΥ�Q��z�o�`��M;���E�!���nf�;ǐ� ��������ȟ�&l�1CO�GjP{���k�4��f۬ό�6i�3J��y�%�+o�Dv��г6��tP�	̍��N�`j��2N9%)#-��]+07*�+$`���m"��􋬣�[6U�P�6�x�'s������v E��D4k_8��f2p�J7Ô�"V�,�0�)ق޲��a=����1�k���@��y�z%�Պ�Ӯd�v�_��|�j�@!�`�o9�ӳ%S{�����;mu��~�ߙy��,�۔-'��רu�qz���u��mO�A��!|Ei$�sf;&M��$�+���Ht����������Dp#A;X6pq��t�}��Vt�-���8����k}�����u���C�q���<���tX8��B���I���� #�&������մ.�+�܅>%��.�D��/�������'2�Hw[����(��O�����"F�O�\�e��-�� 6�;XJ������:a��˦�檲)��f�0�K˚_�Ⱦvg�yY��ˑ��H��@���&-�4ֲp�����v��V��غ��fyFW�hc@��ā���Α� �E<��D�U=#_`�*c��$��y���ɰ���u��n��֏��M�\��� zA����կ��~,
Ƶ��U�}�.�!@��:Y�y&p�&e/xJ�
�u�λ�7sccrW*�֩8m�� 3p�SFI0���a��ǞEYm&��H�ʾpF)#<�?N{�ڭ��0r(~�j�L��q��[����9���MZ��K�%��@��B����@���y�,i{{@�5��`�眎�_�!zw�f3��Q�zD���=Y'q y�N�- 7Z�Y��z���/[~Kg���DT>�T�w ��a�(��C�\��5�����y�z�x6遯NRQ8�g	m�۔P7��䒌.?�V�@Ŵ��7츣�B뺕��P��x�A�T�&��re��+��@��̩��n��dK���ydVs��Uj�\<�$D:��~f&��0zc!I���l���	�OB�p�>���i��k���$��
��HW���鞲Z�x��1,����nץ3����XP�U�<��[ߗ�}��S2�>�r_���t(�l�āE^�Ay@#��N�j����1!�>��������FaV�#�ͩN~�����p���i��<1</�\��Kz�;�1谜)�ܫ��wт����Y�\0��!w�l��bDb�&N��Oh%��i�W��j6�{���M���1�jCG&d�g]H]+�=[+���p�м���8:}�V�|7M�~�$����=�}�L6���K�9���'�4����]�L�'b�T=D]��@ʈ^����5�	ʈ��&/���h/{��G�Dn�A���d�&L��^ y�]�S_-�V��G���;�����Sa��E[pAO ����5�S�k�+#�S��F���^��ŋ ��42r�'Z���P�3%G}�^j�,c,f0n�U`a��w�R���S�ZW�T����\�&�<|����B����d=���_�V�cEn�.��D�)-CGaӞ����W��S�����bx)u�#�b�����B��t�A;oJ���Ҩ��=��
?�H�퓹��%e�Q(±�Y���5�F=����;dt?�~�ߞ�P�	� ~��lp� <+���)|���O:fj�B{�!K� l�b:Z�a7(��!�]�4�9�v�,4è:���V͙a��_zH�w8_�1�o�(�V���g�fN��	��sL���gW`�����f�z����n�=�`p��M<� fe�X����O�I�3�Ɠ��v���R��;5�]�m|��	��wE�TFrmS��On�kh�?�)\�X�c�u&���}Zz��q�����ͯ����`h'���0���6���Dx0���ݕ���xߠ�j�,�$��y�e�I2n�dq��K���ʧ�݇�T�h*��H.�r��rp��PY0˻'���A����}0 .�~x61�^�;��40��9Y{��lzq���ĦfVb
�$?Dv��51?��O��~gߩ�C����\<�lXP���;���}�<��f�{����^�WTo���׸e��&p���e�춭\�d����c6��	Lck�ʳ �*��@k�S�݁��N���
�/��:�ܝh�^�--�S�pd9����SlCS��$\�e�V��oƑQ�\�"�coL��:�r���@&�L~}���gf]SU�����M1�+H?���G�"���#�bG��+����4$6�0��5E��q�_���$��S��+��CRKb ��N��/"�5�����j����۴5Eɥ�J�v�K�f�"���\��d�L��=�+;���5 �S�1�
�E�4����H��.�V5�9�;�@+�f�#d8��_����4ZL)C���@��XѤд�.��(����eN�Έ������GH7���������h����t�� :w�����&�R���en<��Y m�I���\X�.x����w�'&Q��g�g��l�C)y�6:C��g5yQ3��_������o�7g�1�ݒ�E�G]K@���7񦢡�P��B?�����V�V�Q�����I�:�`�����Ow��cSفE���(,�R�q���Dm&��-C�D�2���?+���z�z0��zD�^�@�ˉ���ɖ%����Ⱥⱷ`�5b�d����K?Wm��������u�+4��&~�+��ָϴ�m:"�Tź�a=te�5Cr]����J�|u	�*�R]�y|�R4SX��S1��p���w�ga�:�
��P�&e�nI#1�+�(ﷴ��$���'��u-��^t��Oh�kKW�F�?[wk�"(�Z�ω7���������W�l1�L�?n��z�Vŝ2�f嶥�%�5$��N8��SH�M�>$�RAa	0�V96e�ʓ\l����轆���cE:@ k�Z;P�<4��U�ROG�s �	`
�qV�?'�`��PMUiJ���xe�~��Γ��r�g�a��-�i� ����ZS�мT���vA�'�T�+&�H�4�ƪ�B�Gf����nC���S�ʓECJ�E�ƝGj��sk�kua��i:"9�zj/8�����~[SW��Yf�: ?m9}�M�=L{{��V�3ئd
�>Dz�]�L�U�팲�0b�̌E�[\39��)?T?{/]�+I`�D�&:F�($���\������m���O�ø���%��i��יpbyn�w����N�dm��O�/b��^x�dL�d'|�^��d�v�%]b�.eP� ��9U�9Œ��_l��	�r��H��Me��A�i���Cp��;�9��g!o$�|�` p5�$��X󨅰���Z̞�՜�/w�q����ጐ
*�\�^�0z�z��TӇ����Ё��u�\����}�=��*FgRԐ��MԒ&������rdjM���'����RLOͬ��);��1iGh����oxܙ���E��P�Q�8�}<�Bt��2��6f��jbG�,��J��Q�7o��:�lo=��YܙϘq���$����C���/M��>4�F�L�e�d8K�l�#\�D�����`O�k�*��A�q,3����t'�[�?`|9���&go᩼3Ī��z?�79ٜ���`���k�B�/�m������y����'�
A��-f�%N�q�1l"��T� �ib�>������w�_��MC�{	\xk��(��Q�7�O�ṧ�� ������6V*�HV[l��3���j0s8�͘�=�$��b�H$�p��lNS�O6qR���|��r�P�5o��	(�N�����|�G��'s��ٰ��X(�+[Hh::`t�����HٽD3q3���	F�&)q�HX��d�HV��5����`��p�\�B�˅2���h<��Ւ�e ��W�u��J��ȏ�{fو��=gJ�����'�@+���/YH�;#�+) �D�Cg��n�0��W]��PTO����K��;���b�y��R��R���PM ��e�͐�,�����Y��[J)��u����W`�:������F�)�n;L>^U�0k�`����9�&���&s�L`0jE���:��6�Q�ȶ�4��ݩcw/42��ڙlqew�1�8۞�9��������wq��e��2`�F	㋊I�=�>�?�{5���4��?홂�B���*u��iD���[so�2̾�cd�!���&�/�`�q��֣�U�]�ӒR�s@�I��C/j���i�I.4˄o�WOQ3K�����-�$��R�Oe��D�/2$T�:���3\�\9CH�k�8�|m��59�>gv�a��4z>�JQ#-���!�� ���}2��Do�SJ��ÛQ��DAʪ���#�:ȹ�bwiqM,��
�;��}���6�M㬨�%�w9�����N�����L���Ɩ4��!�����f��3����,=�S�����e,#�H�r��)E��_�Y;��Y��3g�	����h���,��V�	�i���V�آ�N,ŕ*�Wnఎ��b��_D&��E��+N$:U�j�b[ۑezG���j/R�ѥ����0��C��-d�- S�`�?�f���c�Ƨ���_ �p��QWuY��)���1���V���9'9	1��W�t����C`ÿQ5�E	��1�A�I�&��J�=,8�#���?� ӗZU�e�%��[bQ��@
U^���U���/��0a�ր\:�k�	/�5�ȡ2�����5SPX�ƺ<��u8j&2#��,`��`j��*˖F��zn�<�ds��X|�^TC� �i��/��oB��3w�X�^�� T�2�n�/�Dݣ����=�_�"{�H^Ue�:��A��	L��wĩ"��#�c��e�F�H2ܥ�Il#H�fcU<�E�K�fL�Z�'�LcF�Q٩ v�i<$۶������Z��#��o�9j��������K	�]��˱1�)�:�s������Z����]��F?m�=l5	��+O��@� �ykO:WD�	;�����qRNrx���v�g�)օ�Vq�.�(�20fD�ػEP5�![��rW�DZ^��+��Lۧ�<������W����J8
�
3{������ � ��=��a�'�qղL]��yԙB?���i�ܯ'�V��=`-�E>����M��A�=|i ,�钳8�6b���#G���p�����<�)c�����17Ud+iaT5¬��R̶	_1WNQ�8����z�n�Q�`�Ļ�C�H����o5��_l%��PW2�����!�=�͂����n��nO��_�B��_��n���<��%���%����{�tN�a���\VjTw��#-X'���aT4���`��<&�-���#_B�O�3$�j�v"�݉HHE� v�3�����e�k��)Jf3�K��f�+�zC��̗��y��M+d��D��?���W6S7)��:@����MR-/v�/Wjz�3�;(?|Ԛg}�-Tb$�'4ڹ#W�"��t�)�Dj��S��} w�i��_���눋����DH��E��Z,c@�fڲ� ���) p�*�G���U3�t-**޻(K�̞����JB6���i>�!#��;\q�fs�^����g����)'�m]�����ذҺ��$�Z	!2j� <u@r͗WصtL �O(%��-נl��=
F�m�L�(�$�~��i�q�9�3�r>��_멷\�9G�Ao����ȡ��@�U�4T�����C5�����!zJ�۽˫[�F
�A*{)@�a���Ԙh���PH�u����L��`�+��`Q��ř�֬��F<`�{�́�F���]�]��V�$�W�Gg�;���j�	':�}F���I�=��{�
��?��nh��Jo�p�7+�jۂV0���[p.�\��c�N�J��'�Ty�;,��zR��Y9�5�̙�_�"�>v��B�#�]�e9?�s���-w3�+��z�--p�7�~T���%$�Hm��Fin�[��_%u�q�k�������o%�Ñ�f-f���Sw�'Mдj�8��4����1�W��C����'��w �i��w�� {G�$�Xk����w������*�� \�I��0�]U�,^�!k�����/{���0 ��o�|�ΆA����ޒ%�#����/=�"�x�E��"�����T����;)�!m�H8�j�Yʬ�F-���'NJ�������e��s�n��_E��RW�%X����	�쯏����~5�ύVg�Jn�E�B�69�7Y�?�NK)ݻn�)��t���.��";ң�~�4gO}��1X��@�.��1un�uDO�z5N����y#��$�Ϙ�l�~kdA�p3ړ���uc����+��K<?@�N�hjFK�Eu�E�,lVlo�՛�n]mcn�f�0tP۳������ͧ�z��:�-�1l�tef;^P�1O3��oh��$>���׬e���*m�(����gP�,V��kq�|6ރߊ���mM|�t�p`mَ�=̂�ld�ߌY��ID��>�#��w �T�<@m"3��ΐ�B�f	'Y>��*��,Բ��D�V~�Y˧�TK�f�|6�8����m���RX��6EՀ#�w�Sج +���d:�,)ڕ����t����w�����TK�7^��uڊ�0��7d�/�5�(�8ȶ��O��Ȫq�Z�"��5..$N�t�u��*<��@]h��G6�]ȅ� ��¸\}�H��{��GT�_��4\�s^U�*���c:�$�T"�oi��e?�'ԼƮ��5C��%��T6�����!�� �{���3�h�meKS�vz�|S� "l[�⬈���z.F< 1Ӟ�ߐ�� �7�>�`����,m孳�ϳ-����v[-}~�"�?��p��}wÙ�UN4I����`���$={wK��$su�'���<(>��r�R�n�"VB�S=6uEX�5�݁�5ֽ����v>�T^{�����B�Mu�~�S&����&%c���;�H(�0�'(H��)�S�1��SgBV��|�;��1)�VB�,�MCѴ���=�۰���`��J�O��Az��!qy� �F��y�&8�u�{�~ h�fG���1����OWB3���A�F��`Dڧsq�	�&��L����F�zf8"-0;�w3��Z<��O
%����п�������"�x��(�/!��߂Plo h�\_8e%H���&�6�wv��Cu���.��?�JUy�c�h#c)�G-;�l������h�#ei�[����,��]�2jJ'Eh`s����>RᔲP��O��/*��,�T�hGy�6G�k����߿1���H%�|ǄϸY	��\tx�kO"�q*Ȑf1!�/����k9��N�֔6/2�џ�C~a_�v��Q����}Qf��@DS]F�}��:�Ɔ�
����|��iKƲ}vy�9R|��) ��ƿ����ni�߻G���R�ڒ�̡�>}Le�|�y��15�:+�o�Π��s�]_\70MvL{�,o���Ûa��|Y�ud��[^�c�+(H5�S�>��<׵_!7�rB*W�<.��j���?+}_J�_]:!��V0=ՃˇK�zC(�\ .����Kc!z#���l��t?C��'�B3������+
���i��-=H f~{0�8�ﮠ�*�]����lX��(�հi5��!�f_qk��
�k�K>��U2�qǫ&]#y�����ĹWij.�|ͦ%�*W�r������Q�{X��=��H��s����
0 �H���K�����S�i���g;W������-Ea+��´��h�0�3�i�ka4r�*�ѥ�"�4�C9dpF�Xwy�cF��;~ @�jSo-)��-~"��tf^�vGFUHhl�b%��?j�4�y7E$��
�l)�tA�vD)1k_��ͨV�*I�Iȁ~�rs������9���J�*㇜��p~BϠ�R!^�{c�&1�}���Be�0���;G8��XO�q� a���A�6sԩ�
u!�3��������G����������[$���^���;V�@3���KV�j�m��#x63�Ԟ�I�F���D��[Q=��a����YD���*�Z%���v�_��S�2�*��;h�=��%�E�P�FN�k=�s�	)w#c Y�t���������;��R<t�����Hi5��E���e�Ti�;��B�2X	RF��o�Pu*h�zO?+�w�K,әh��nj�"y��T�[�����K�������Q�Lz�#���C|��i���B.�4��V.\�}i_�2q$��>=̇�́p���fX�0���G7w�}��*��\�&Hs���8���f�_�����޳����H+��P����u�3~3��������"A��5/�᡺�nWՍ`�Z%�J�|���bC��f����P�g%"oo���1�����NZ�������C|Q[5��'M�x���t W�u1��X�>n�a�nN#q�k
߁ls���Ò�9Tn��_KD:e���Wz���,h��K\���~y㚲��.K���f�M��Q��9@�b˂gc֣'A\1tV��P=&�B�1�0eb��7�U\����.D�|���H�8Yl��7c��*K<�V�;-������E��-��#qv��Ò5�P� 1`W�(>��*oyg
�	%�3~85�&�����Y�Pe�6[NDTs�%D��`��֠Щ�B}�wQlgh������|��ŶUAl�w7����>S�/$��D>��j������^9! PU�*�
%��1�d�|͒Z~e"��D���-)cS�NP!��hvi`�"�Hz�<z���4KS?>3|��*��y*�7�/�c��Ty-
����T&�p��%F�W�?�I?�O��H�뾵��٩��� �E�]��������\��Oڡ��T��t+Ke��ۦ����� ��;�{"�Raq���5�?λQ� ��`5ˊ�P:��U���ߗ�1/I�S���@�8B��uO�Iv�� �}�3�a���d%��GU��Zi�ac�+4u�S�aޞ`ǖ�c�E�=:�{y�.DU22�0J��:v�{n*5So׼�Y7��GXijǞ�SQ��(�)�8�7����!c�^���Q�s̊�UsL�G��d�q�=T��XSB�CF+��#�G�?�O�t�Nc�����zT��ө%5sX��yj��g��%�����4����%됭�$�U��f��e�N��S)d	->��W��Jg�vϤj���9������гbw��L�+T�uW18������6'��J�I�\Rժ&�W<O�Ђr��V>�Wu��(V�Y	�X���O��s��響xյ����`�����R�8$E����l��-\�@P����)�FMe�d���ȈH<��AX���RI�b|fG�M4a�њ���oq�JXu��?5��WgP��>꼪�xb��VGw��Y�8z�u܈ut��}۵�|���x'�p���Ŏ���ZRp�ڌTN��
�i'�"�Խ^8g X㊱��M���+�E��>㑝݇H�9%�?^հ��D[j�	�ч����鮗1F�9��!�VɩU�2����k��X�K���h�);wTv2k�,��0�_�2�����\�%����)T��d��^3�"G[ž(��B'kC��+�ش����݉�h�4��6�O���%�By`��V���︔�	�*.r�'��y�@����m���ʁ>]g(et����c��{�&�� ��h�N����L�#!
��+[x�ef<���7�z��_��#�Y�X�M%%<dB��ב���QP ��ny��~T��3�d�
$	po�{R��Ѕ�l�'9r�`�����p 7#.h�"���
������8�@����E\���󟇐�����_ס��!�vQ7
����E�#����yF��Bц!�*��@��?#s��-�su��Lo��@��ځ�ӝ��c���7v�	��U4��u����L+޲��/�kS����)
����S�'B�XI�~R'"���-
)J�dW�69���l��
���߶�b��lmW?��E^f�
���eymB����	�<OG��KC��m��5J�_�7�N���k�l��Ml���q��u�v%�Q�1���8l�}�S�U{��q/��vU1��a��J�&�P�g�����B�6�WP���n�B�N�S"����s�*�Y�}h�P��cq��P��NJ]�p�?�����
=QD�����dc�?�A��.����V�����1�/�j��`���Cb��=JS��<��n����m�(��I�+����q�0��d����U	^��2��P����.����Iu�S���/lo/G�2���U-O��a{�c��EyU�vP.v8'|i	����Rl��%�i�=/��HAh+����M7�~`ta^#Y�zB��W ��_@�@��P���P>�T���B6��G�*f"��EƍB��Ƕ4��М�L�T�rQPpÍ��T�?̤B~���*>���S�H3�8�C�8;���!&��RI� ��ȍ�.�^����Ǫ��XӧC��Tq����Pbd?z9ŠDѪ�H�Epy��Z(�V����<��j}�F��y�S{��2�3ݤV��(H��N ���*Ǜ<��Pg�N��?UX��]�LA�ݫ��<��&3C���.Ţun<��MCw��JY�N���X�)�( ^����{�\mBN��P�L�8o�i)�ia)�r����|��*%��?-���w��D��>�0��Տ�����N� 3�)(}I���$$E���Y!�D�����1wp�y}/�H4�?a���)�4_U�b�w$u�nbB�%���m^.Rc��HT��+��}�Q(*���g_pApv�V�a�ߐk���EA��[�
�*�r����'��P��%[�U��܉�b��m?��S��$h'(C�}R���e[��@�՚>�8�y@�Y���
���8Π[9ȁ��}��lp��!��n��H��H?����l��\p�&;�^nP�he�9��R����B�
M=�Ec�^��Q�^�wBE+�|�Uf�?�Ip���W��HxVp^eSu5\�E�5Fe4#im�'FeT|�(���ǡP�f�3��߽xT���7�yEO������	yЊ�Sሶh����jxN�S�=��� ±�f�}M�t������`#)���I�Z�d�J>Ьd�JKjv/K�.yqW��ַ��u��(��/�j��'tN����^�%ڊׯ�3�,E.�������#��--�Km~$��o���^j*�P�9k+o�9��1��L�d�o�2�U�A�]:ۚ܋�[��;	�f�p6®$�R�GMެ�M6D�2p��~��g����r��.v擳]_���.�X��~��6�QM=%1dc\�*M�ʍ^P%��kV\��ձ�e�(��B�v|�L�Ŧ��H�> ��-��i5�ˤ�%|�,�L�t,TRoZ�T��F�_�BŹ}�"��kaG��9-��s9�ܯ�,�o��++�q��8�hn�[��jYf��<��j�ht<����ǾF�P�+�kZ���p/XHO7c=�+�޴'`v�qd��l�=�2)��$V��[K@�S"եغ	�.LyR�0o5'D���d��>Nv�����r#މZ�,Q��Vi���	�BbAܛA�1�>�<�EXѦA�>�q(~������n�-=����9��p�z`�F��N�A[�P �}���4@���~�\��*���5��7�3�@5V�o?��=��F��'�+���NA5�*@�_�K�J)���bH28��x�p����oT�i���ؘ�
���硚D� ;F�`}��k���4����� �����^b)�����w�G��{d�R���q��^��`x]>ʣW�~�Y��y�\ۿ���$q�ja�S|����^�:��>����R��<�"d6.��q�@��C�-�v�解4�. G�icR@�m+�FZ@V��/v(U�$����s��c�:��la|�{�~�JNX��<�	SP�L��m*�b	(�^�<�n�󚬊��i������ٛ6�!qNn�T0���%&I�o:���o�q�ZPl��P
���S
9��pL� ��x��4��?s��Z�a�������v���˃>�]&�8^Жp�S7�;Wp!bZx�O���q��-}C��2^n�G'	�X���[�ݟ�#�/�b������N�Q���%��̴,�@L�iz��K�^#��8V�f���d�w1N����(X�.�ⰿ�j~�tab�7Q|}�p�ﺤ8\�#蛒 ��V������/j�8@(ĸ����ʍP��r�2��E����["�K������a�D���(������znLm
�*bS�'���/���?��q���ʾarSM��Zq�k�i����D�r�"�ܩ��Ҕ���z��P:V%qv�h�N���.X��pip8d��	�@�	"o�HG=����RE�W�H<����mlW�à�p�r/���|�t�qjZˌ�"���CUU�ts��Su�*��!ѐ�o�p��i%��wCb�w�7ү���X>�' �R�k�����0�!H�H>�t�Zr��(���}O3
'�h���}�㰄�
�z@I�����7��������u-�-~Pع��ٖ�_H���*�D�)v�Rg��AI�F����/�����:/�)E��A�)?E¨�5]JG�z���rdj�1���w�Q�Z�
��{g�Cr�L�`$����(�2X�-�Z��6c��E����������=ﾢ�C<�:,2��;=&PKã��'��,�-wM$Ded�;t�|�-�3ٲS3���ƾ�ރX�l.��=�r�T���!�Q�S���]���*���h=���m�~��
�RG�ݙ��k��p�qPW0�����k�0�A8(���r)/�n>�S���4G ���R��D��t���^��/�/�e�����/JA����_^w+:��R�5��˕-���j��q�.Đ�h�V�Rx�=��з��e��V,�����K�睂d��d�� d�f���<��C�xV�͆��PmD�^(��\v�-�>ю� ����Mܗ��j
 ���U`����p�ߛ���ypN�����yQTs7f��a�G�� �l!�n#9,� �'��}$�R����Ty̰af�	�j|�0�Q8�4(} ��k�;�1�L� �2B�T���،yqHQ;:��^��p�t:�tڂ��{]�ʝ����V�v�׭�~�5;����P��-���7��d�MpA�l"�Np U'��Sh���a�'��;9�绞�s ��Tf���ݟ�0���v:�i�]��#E`{�R_�x�Y�M�Bծ ���*��1�/���y(��7��V�hcS�9?r�ԑ���D[DUà��V�`��<�U6��
63E�e�A�	cH�(���ߠLM��O(<z9�X�5Murտ����ʒ��^b?���I��j.8�:�P�|�nhi.U���G>��a�*��@*�� e��i��f��n����rsC�X�&��,�������R6zL���wL��X��BY!�i^��,8�(��߭��'��%|�OR�L*�b��ŧ�$L�lH{�x�V��rV/H�Xu���P���m�ɑ���H�F��_+�ʀ���u���G� ��c��r��s��.V_�U�Rb�KA?�"6S�@VH�q0u��W
��p�/�=6%Y� p����Tf�8![�v��Ņ:=�3�jyq�o�v�G��&�c�4c��.�˄&��u�N��ɒ�&�P?�U���4�>�F�T��W+�T�~j�CnW�]Ⱦ�j"N�7�,�������l�Q���yȬF;���Y��3�@�gD�%��i��
��`����EA���lt�`�$����%:�8��^ʷ���!�*�%R�4�[g�S�Z0���\Z� v1�U���R`E�����W��2��ZS�/\Z�ˁ�1�;�m�y����K�*�p
��ê��=��ݬ]H ض��k���@�T�'%)��yaF�)Pa-4(=��l��\�@�ԑ'��\p����'���ǿ����?4c�� k���2���%~m��e�w9�+��Lk������ �XK��A�$$"s���!��={�n��:�oAdG�VMQ�7gBA��L����k���'=K�ݹ"��>�X<�+�S�m9�o�p�E��@�Ra��!�qq(��)Y l-M�I�S�%�Q3{��㢔�~ם�cO;pU !�x��}�Ǘ7���Q���͸��9Y8���I$|�<!^��#���B�\��b�l��^��r�����d`KL�/D�{����ȿ06�����<�\7���nGT!�h�
�����][�b�������ｙ���w�~�"���Ýo���
��b�Lщ��gq��Q�ig�Ad��/�T�O yի�3�w�b�0��;�	�!(��v�N���h��,�`W�� �vK�t\J	�B6�s�41�� �_�k�ظ� 5�]4:�x�pF�Y�D�9��o��Gmy�C���)�7��2�Ĳ�a��>{�����&�����ˤ�����)�p��Y�b+��eo���W��yD	��g�"iA�`H�K�[�J���t�s���)������S���i���FMwe���OOݬ�Q(+3c��L���H����9
e�](��N�@=#6-�J�L��P�(^sy�ҏ܏د�|}�.	@]�L@�?��l��_�Ð۪�'�)S�8\-�*ȹ+�ɷ*�T�V3V��ӏ��U�'�-�?�x�p�"�a���/I:�#�$LE�@QE�	I�PsFY�b��:���o�X<�d5i�1�p���LJ�z�����i�֫�K2g�:��+6�%&?%Rq�O�#�5��U�����Uo�wc	T��ࡪ��3�k���
�$����ۊ��s(�gf��= �L��qG��*���]-�M�G��G����5~l�ɩ�)��g�<�w���f,F�;���� {�h�T�W3�[�Az�L>)=I>�t>�ٝ[<�~�lD	�\�����d�>o���C�cD�?B=�Ҟ
�mX��o�����J��*Yl�2�����53�Wg&@XlZ!¶4��tmx`Y������Ps�e����°��r�ŉ���ډ��$�%���,��k�����̓k���5ѕ%���\��u��k!���J�q�h\�f0�X�h-W���]O^� x9 �D��`z��4�<Y�o!��9b*���I%�r��ޤZ���#�*���.��uF��Z)���M(�i�"��Zk�ؼ�_7�I��&p'o3ˮ]z�Y��kMoy�I�l��[;�k0j�Ǖ�����pƬ��k�hD\�H4|FI_a��nPK��2�a'��5�:3��Ћl��6�C��N��Ad9�"��ϫC0D�"@���N���a�5=���'���a�	|�s���Z9�fBν��w��퍼Z_iF���n\׈���x�DQn�%?���[by�?�5{qG|
ɲ{1R "td��	;��[�aa
b����ə����E��*��9�f`����k8~����@{jL�D�*_���>���f���x���o%?ֺ��5�/Ё0���\��z�1�9B$i7_��o�ߓ���|@O���K^�\��6�CZ¨ȉ�p8A/Z��}4>'���E3LD��&��'�N��9� ��u	�
rf�;J8,åGK�
<#��+��Ǧo.�B(@�@�(|�<�c���1h`seV?(�I2�;M��4o:����0p�~���9\T{[[n�!��1bأ���|�3����)�V\㱻�ˣ�P2}��#�
��>���p$�꼣�I���!*H���?1nY�og`L������lڵq�6�$��o�Eaw#��C������/:�,^���9���9b��Ld�b84y�~y��TTH�8�SO(|˄qC��+ N?+Ix;��el�lKd�T_F�����wJ�Xp.]8�u�בbbb�av��zQ��u��BʏS��l�P.�}��8�\G�|��c�N���O�e	����M5$�Q"�2�~J�w�Z���mY݈Y%�����13D��#n!I3�[פ7����͵�� �YX��\\R�����A�S�A���������_�P̐�w�E���:����En������+]!�g 6��0��7�S���6�b#;��%��Lb�/��h��]N{��E��3��38�y �K���	A��y�R 7N�9���Y;�,!���"��e�ڢ;���N5����A�L(V3������vl�$ �!�N	�B�|݈Lo�"�{�y��F&Y�q�eۥEo1��k���ݻ����]��f��ĚٞѸm�r����� ���i��UB��`^Qm�7�Pw񖘢�.��'�5��:S!���K��|_�[YWߋ�1��$�U&rݷ2zk�}}��*��DW��L���h�j.��&�A�.��&�w@j�e>�1��j�Uj�'	�O��M}�~�䑑v*�+�I�M�B0M�E����K.U];s��;��{P!��a���T9��&�ߡ��R�1�����ފ$~2�wd�ǈ��Y����ӝ3__!��6���־Q�Zkzy�|?�f	iT��I�>Bt�\��rI-k�_�ŐqԂw97b[9Y��v��|��)0��Lts:��p�0&\�%u=f�Z�'2�Ð���7�L�%�븋��]:^�GD��w�M>.���"�M�&�w
��k%S@*��J9|����0�Ayc�1M?8���N��e|�y߅�; �z	�8=�� Y7��g�:�&EN$K�[�H6��5.v >4UA>�-wf\֎�^�Ҷk3߻�5)��v,4e
l��81N�4z�ɪ��ͱ1K�����[ ��\�B����O�%<3�i4��M�
���'+BW�E�OB���o�=
���d36�&iq_S,^)C�l'c�� JObSX�x~��T�V��0}�tl@v������&{���C��u���J ��ؽy��B�C#Ӡ�2���b�=}}2��

)5��TW.��Τ�6�	� ���4b"��|��2i���3�I��v�a����ؑ�1�9J`��'�Ǧ+Z�J���r:]+��-\��~�'���{�b�[�dD<��W��D��0��mQF�> �m<Yأ_ $o"�~�����jG�"$yeT�v{��U�~��� !�>��lS�U�Wef��Ri`�Tq�<O���	Yt�'�r����W�H�b�0{��7�XL�WgngG<� ï��B9�������{�y�z_No����0��*�#��1�4u1�=�1�l��7e��5�J_�������5���Ϡ�F,YN�gP��
��xѡ��/P�mΠh]n���2�*�X_�"/�|����� n2�:	>��Cc� ^x��蜁����v�P
 � �O���r����<�p���Z�z����MUυ�F��d��9�a7�ւ��[����9������m*��k�)b�ޗS$"~��X)g8��t	���.씬x�JcE��y��~�\O�r�!VkҚ��Z��T�:�B� �]nՔ�80t�}`#�^�~��G�h�#�F��!�}K~�}D�d��E�+��ߗ�ck���^��F��%��q��Ex�A�(��)�x�zK8h2B�_�p�6fd�3��^�	���O�Ա�f�� �٣t�ה��|� �A&1N�����"���`�&�
�L�A��j4�T�e<��i&��ߖ���7l;Ъb��M�ݿ�I0yTέ�2�.M�����.W�y!!�A���(5�U��o�s�dJ�#$�����6<G@i�����qJ�Üo�1�/{ɫvFE�g�#�\�lի	_��ǯ��K~܉����^$x"�uKb+��ӄ0�y�?�{R�N��+��x�je" �Hp�Ps|�[�h1bx�m��ƒÉ��,�`�@ؤ����y@	/
g3����������]�����o�q5���J;ۍ�YO�0�!�q�bq�J��_r(լ��}�C�Z��J��M��I�/ӷB��ߞ ��E���`�m=y��u(�i�wႹSKL�Mk8ߠ`���2�O �7��V="�ƓY�@��/���{Ex?>VOE���F9�UD�у������r�ʷ3]���C�+eN��X|�7�56�P?�;6�p��|�H03+����^Dt�C��r����\���7�Y=��	Hf\w��M�{c8
�B�	C�M	���-T'��,�CW/��i_��5�R�v�pG�!��07�!�F��v����3aQW��8��W*���kev�[_��>�q`.>���%z�d���Y���s���p~�m�\Te��/O^w".���)n*b�c�C��D|��C�ZmRS�|��nD���\An�B �!Y�R��y�b�/ϐ���L��b"�BE�ڇ=s���Y��wOL�B���s�.�ty,l��m�]�Y�plxɧ��,�i�OB��tp�$�����*�i��N�i$7:m�����@�r�Җ>!��jsQS�mϱY��p���+U˒'���b)4�������iY��ݳf�(��Xܳ,�JR�,�"�ˑ%,��SkPM�%����JIH����\3B ����:4@�g�$����5N�\�����U���h�\&h�����P�'�9�A� �����4�jslc�L|�0!l���"sv0�6�Ϫ����i6���!�#��2ī�5��v$ӛ�T`�F����5���n����,d�8<���g\�>c�K�];f`�\����b`D���aFk~�o.���x��q�p>�|�W�����Ĩޚ�ŭ��5�pW1g��`��m�z+���Fت�(������]?�PVU��.��jD�rocK�����&a�3Uu�Q3By ;�S7�O�ZR�]}����S6��-G	L%m#,e_��S��\Ǹ�\S�
ې}u"6|2�|,�!@��y�n���-ҡ���a��'"F�)`�qQ�7l؆�ة_ݻe�'a�ߛ
��oV5?���yu�����ػ�u�����ө�����C��+���eY�r���|�Y�bݳ��Y+��ُl�a��c�+�Za�#�=ۗx���,}�K Q���*�HRЯ�R�,33.&WPJLn.^^u }�;Z� �U��!2�7����,/�ͱ�']&�oui��(H��WjY���gHp��r��f����"���3EuxE��ix�Fe�Y�)E"Srm���G@r>�����]�_X����j�<<-�;1�1l��qi�w1�� �i��Ӽ����d�Gsz>A�nx�D��i��Y�Nj�����l�;KiFtl8+�����B�l17$O`<��3&=(�`�&�{O��%ٻ�	�Z�$�l�@Q�F9�ᬠ;`/$���x�[��G-[��[t�0pu��/{�T?&����fp�\�ך�֡�Z���
5Q�@c�}� ܐ7��N�����l���#wo՗�	;>N��^0��9�*�ǽ�Ĺ��ڝN���f�hu{!��<��:�|f;���O�1�\���O�h���K��.8<�-�����5Q�IFd�	�T�l�&�H ~�k���gc������AC�e�Ʉ�dr[J�O��ڌ)��j�OÉuxN�YN���L6��8��j#Oˋ�҄��}��CD8�׍#ȏt�^"� �R:�w�ȑ	o-�3�	���*A����b�X�Tr&�9�R�o����p��C������SP�_<��c���[c3���]ݝ�I�fq��_����ޝ?���ۼ�{�eK��_�Ly7��ӊ2��̴�^9,�����?��o�&�k�8ޙ&�Y�*d �ќ
�L@� ���;J{,���hW
B; ov�UC`۔�[�Je������'����q�eW��O�Ɯ�R�4��Зk�{���v�'j���<��`O���j?qОzZiD�|ڍ��%�������=�"˝��։,��#6/a�ԫ�PBM�	J����;�q$\�铊S?M�$�STYA߿�X�Ig����&�� B?��>����W�cɟF�t��N�j�jLμ��Oѳ�[���c���,2(��ar��^�kHi�q*ӊ�[�"�{�DO722�_��m��Ӌ��q-�'Pr0�䯴���L������R�Ǽ^��Ա�i�  �v�Z���,q=�����,���ů��vԍ�5�*m���pd��v흘���W�WU� a�ϳo�hdA�#��zp�����1��U0eb5D>a�*��k�t�"U+���Sf/e�2j�T3�|}�8�V�3-ܖO�~{���f|�;T�ֱ�=��Lz Nɇm�B�Tw�'ܗ'2�[�]H���NS&N�h1J&ȡ����)`S3eS�H�� �.��x#��VI�/�؄��^�c�����,r�L�PLj_y�����g�+�QI�v\W�"�^xtW�1���to��_�D)y�BO��$qa������pM�t�n+!���r�<�r� ��-��i�%>6bB�D���Zm�V����f�L�q=�f�p�2?��]���[pE�����o��F+rq�e
)��f��-o�rC�L�0��P�ʅZ�`=�q(4��$�޳nԞ�1G?p'�d��Y�'���uե:o�y7�^F�|7�fl�+���@�B[�)�YZ��ꆏ���	�����(�ֆ���m�CF�
�к��d-��z#�q�_.'D�Y�jeF߽QJ�Y�A؟�����=�8�����9C�X�� �~yۙ m%vp����;�m�#ݜk��4'r��L��S�y�D/7��p�8'vi�p�>��I�(]��(���_F6}�>����mT�}A��w�����W���`8�@Y���5�L��i/�PV�6�P��ͪ0�U�J�O'ŲӜѶ�?�7�I�hVX%����$rj�Iw��؛A��"�%k`K�&�����LPN8��qE}���50"�b���x߀�����İ����o�]N.�
h�%1�0� ��XNs"�i����&�W2�[�Z�B��Ǵ��-�2{1�+��W�1߷�bNR�F"c_P9?S#㛛"�·�lП�g��t-,�k2����޾���6J`����dv��*��0��ytȓ�/JİJ�E�VE���1Ŋ��8�E����*�"h��)�]�:����z��\h�Ԙ>R���M��Aƹ�#�1Y몱%���>�D�TKjRj0���f�8�jn�"�f���*l��p��e�/��N�hB5͔[�����|7?��H�>э�y߇U��G��o\/	bTؠ����A:T�d�����c�F
 ��q�K ?9��&k�h�ǡa��;ƞ�I�fq��刈оJ�c���0�Al�M����+M$ؖg'ZN�RpގI�����T�{�`��]	�,����y~䛁%����9v�c�E濛k�:��c̘��Cčg�q��QőQ<�<<�~��C�[�6�O���}�m�P������(^L�s!k�d��i@��"�M�g����y*�HrXa�O}�oU�Mj��+xD�inp����A����_�z
��-�\Ȥ�P]��Ǻ=ǣIF��>^n��_xFNn�/��J� 2��\XO��ty&��{��H�%ļtw���͔)B.���M
o��4��B4���G��"·��y]~��*<���������0�1F
�*܊�g�o�U�$J��s�w5\��N�P��&�ق�E�0��wMir桞��-��F#O���l�F���u'1�x�)��~ܩ�O9s�$Z�����"B�R�a���;/��_F�I�i�+�:8�`�Ii`��x�pJs$�^��@�1���aM��m7�H&{��(P9@OG��ܓ�9�K@����C�4��p&FP�0�޺'Ѿ���^���w�G�� eQK#\�Һ�w��Ag��î	hY�|�\�1N#i���>-9�ZjM�ݬT����� 7f�Wrg�|s״���[�J��
[r��9�n��;R[_�W;��d<�J��!�J�y�;7�^�����e* OIP�NDHB �#�Y���9R&Ui��e�7�u\'_�Z�G	xuY�)%��Gn�F-~ͧ�����e�s��P�^�_�r�=d2P�_���!��@o��>�]}%I��A;﯐�t��#'��΍T"�ua]�MR>q�]swz�uj�Y�A	@�����9O9��G�����.Z��>��s���f��ZۢJ}	д&����[8��k �Ա��.���k��z �	[X̛^L�2��]�iH�b��pڷ6ee#M̴N�n�m���]��zO�� �΅�J�2FA5�?#�>@UR��ܙ0��'��&��&5�G$�_}H�l9�9�8"I_�I��_*hul�^��=������+�"��|;l���J�K���,	���gxg�}_D�s�<A5^Y���|&�x��N�j>&�R���C���ekB�+�*ޭ�kJ�Q�h�C�&��x'�M�Z�)N��uX���X���Ic(A��A2.\w��?U���5wx����K�3��Rh��}��>ĝWh�I/�����S���<nR������� ��v�%kH���I5X�LmЇ�Hv��
&�'�� Q�kX��)���9��G��γ��9?�����ssu*�N��ԩF��]�|?n}
�ve���:�|$q�k��!�笿I�� b�����)���ӫ�^��y�x`�3⌦�%<]}�SMcW~�nHy�x�7=Y����X����|������=_�q�k�����2�C��٣$wˌY*�є۫��eE���B]'~�q�"��2}��Fk)�g�L_A���5�l|z	��� `�`��Ҭ��qnՊc�ѐ ��x`���g|��Ӿ�"WD���p2sr;S���"���Z] La�ʖr����ts�MP{Ȏ���w� ��S��_HZf�^ �/��q�&!��2b=CQl���PN��)�n�s|�a�\=x����c�j�̓�α+$qwb�&�Z�E6�Ԛow(zj?��6/~F�:�����\��ʇ=o��k���'L�/���w���R�m&jPfL�R��n�@=
�e t�u2��6"�X�P��l�"n�E𒧑�PF��&0}��%���`aJ����tqK=����;P7`J
�Q�2\�;�~�ϩ
�����n�N�E�ۢ��be�l�߷�x��)�H��4�ޜV�x^d�<Y�N���;b*a��5��B�8�a�P�v�����iJ�a�9��Z�/�4_�L��N^��Q�z��ѴY���a<|p�$�V���� ����~�	��)�YC_L���Y�0�˝S  ��R��V�E�~zvi��q�,V�ŴNLi�4������ӿ�����ԕZ蓂�@yV�P���0�
~^�j$�8��m�����5e	��ޮ�U��J�0!��|�t�8@�}V���C���"�H�YU�x�
��%	�S?J�����rٲ ��G��IM�(�����"9Z=R�K�g���**�X�s��S�Eyۼ���������Jz��.(�)u�x���ă�����t�����I��PO R�6�N%��Q�I[c�Ȣ�Bq�M�~�Bz7��&��#$��Gd�X>:��R�l��	�����I��.���P�l��q�O͜6o�Q�ʄ�p� �Z�4a�6�PG�<��Ou�!%�)��JV���;>u��r�髰Y@������h�� B�p@�������C�_��r;D��)����5cu�rU*��ܿ��zCuͷO�B%������1���<�j�<�f3%&�ɟ�d�@k�_�2}�ݯ����yP&P6��F
'#�}�`%<���3ws9�8�{�*Lᘒ�:*������h��Iո��΢c�
�=Ean��M��vu�h%��L p�v���<BT�� �Ӛ^͹G?PI�_A��M<ew�t�o�/�(6�e]�����]��q`KQ���r�BCB�|��
z��;sh5�4��C��M<�ZCy��<Y88�%R �!d�[��H�jB.g� ��M��ͳ.G�B��>ϾzJ�����}���
�,Rp��`K/O�Z>��ʅ{F�
�,f��f]7"Q��Y|�_�%��I<�8��ǐ�F�^�0��V�����]���1Dj��(P1ҙ�LM�����:�O�ܒ�������&ʬ"|e&Ϗ�߄ �<��: ��%|�X�m���+b�r�H��xRO�&�R��������R�g�t�B)@�OH��Ədu��J�M)��� �gua�M'����3r��Ew�pނ�ט�J���V�l�r\ay.�T�� ��%�i��C�a]I-���5,�SO�+<	��AiɈ�5ޗR��V�̵pH"���U�h��H�l���_���c�B���]EA�!���ҵ�t����dj�5:_�,�9ۥ����U1T4d�_Cf�zZ�H�VA�r�̿v����W���8���-0#�+��P*z���n���<�F�L�?L%9�]AI��H}�f<q깄�n%�-m1����������#�����������1]wq�iʔ'<�ZY�	�11�jm�;D>�8�@�dnqٕz����M�o�Ŷ��/<DG�^����3�h<��G�#p{�T�s���x=_�7Pþ�&m��r3�{�*���3�L'���2x|��7�*E�NӇ}�d�Y-���{$��������e|>�|Ņ�W'a����뗙��%�D�4�]
W��OM���$3H�XH�+)�ǚqJ�|�%R�Z�{a���k �b����+m�HZ����bC�lq{׊��� ���%���Ϋ���IȾ4YR�2
9Z�<oס������&�ђS���UN���l�|0��������^?#si}P/��y˿A���.�Q�A[7�[�׈�k*�Ω����sbz�3"A����Rb��R}�@}<�@�gqB�+}k��K�g$��ޘF��*`F��J��a��W��+��.�)>tVs�Yhzo�.����������K�{���m)�^FH6DY%�A3"C��տ�++:���[�-͐Z���bw�/�e�T�f����X��:�A/=Z�	��C%�7���7v�9���$��Ssf_J��lC���'~�W�c�'�*�:2Q]eQ����۹��kB��ko���8u�ǚ`�)t�O!�|��!��2���l1p�7�ä�H�
�Ǖ��Md���Ԥ鹤22G��=��US�������?���Ѓ�V�}i��õ��!�nd�~#�\�����a��(:�+�������}�J�E6�5H��� �("�l�Y�� ��nN���Jc8��J$+]�����_�O���D�.��'
`���I��\d�:5.�H�6���(+TR�?��+3lʒ������3�Lџe<���QXq��{�ʴ��:.��&�׏-�m�m���U��%ǘ�U�E�xm�@�/��\~�AV��&�$)7�s�M��k"�|�t$����쑗� ɝ�m��������h�O�j�����tR��1�JU�D��®�!q�+�����L��EOM�pR��垑ß���叺�?��u=�}��E<x5'\UdҀ��O1,�>(�Mq�+{67�7��/���_:�S��?%�ћ�m�4�w�U�o�O��!�\>g�v��ʬ�%���YW�4��ZƟ[-�s����Āyp:�0}���ߟm0�	uE!�c�7!X�&��$�{0.`!�W	E����nw���
{����tFy3Jq�l~�7��"�g�	��~Ƣ�������{��0�� �wE'�q0��Ϲ����w��V�+-
�=+뤢����^�*�C��v��vN�N�����ڄ���H�:�
���s���Q4�p�֮��/(��/^Smg�Ů��J,�w{�l�������h7\�	O��A�5����)��jhwO��� Jzq Cڎ �x
�eG����T���."�Y(δi"�No���:��^,������F��UÍG�Et�ƭ�KN�1h������bnmu���qP��٧-9��싣���qu�t��u	��2˩�DdQ%c�9W@�f#|U2F�x���ge�������]��W0����P��� hO���c�;��7�O���	W�f�T^�yF^,bE�V:YT~[������#�e�rW��� �V������>A8���tֽ+�l1�b7<J���Gӣ-���|zx�u���F͛�@�L<�]��>ry����~]��s_�K� �h�`�nE���{m��dB�����W� N������u��}��Dժn�V����֘e����+��z��·��v�7��f�XE�S�V���%iT��t��IfWl���mT��v�hI1��XMɔ�@~Y�¯knQٱkd�ہk�08Z	����Ic.)�f�p�-�bQH�ܚ�f3,��Ną��.j�|�ǯ�^�쭹�+������G��\��ک}Gr�=��@���:-T|���	�L���/{4P��o֡�U���A��"�*���L�-t�[lJބJ�Ņ�zS��_���G\�>x�<�&鳒���BK`��"�49WGBu�;�C�����U����s�-��sG!#��_���0ӭ��iݑu�e�*z�ڥ.1���8���ז=��'��m�X���}W��iu�N�+��`�Hw�g�����LO���
Y�!�`r�)���G5q��7�z���R���0�>�R��	9��L�`�t��q4A��Db�Mĺ��C�.z��E9�2@�Ja�S���DK�q�3d�p=�&	t�Gz�~w�-�}쓒p�aO�B�;��7��ΛnR���i~-�� �l�L��myU����:�:�&��{v��;�����ԡaN�G[84y�����s���8w�۝���اB�	��Nm��"E#����i:���u$,Wu��9$�;mC�ݣ�v^&�&UB��
�ECP��d=tɲ2���*���q�-k%MM�5v �V�$F��{�9(�^c45,��b��i��z���>dU�c���d�z��+�Z	�Ø���oT�T��} ,�׆����>�Y|� =�D�c��b���#�("t8�.��[U��g��A8�Y�Y9��*���}�a��E����7$Mw��f�g���0�:mx���k���`��7�-Ixh�{tyz��=��ZOy�����,.�P�F�),	�An|+@2oӺ<���4�i�fr�ig��z����^���$��qh�m�����8�����K����@�>��Vh'��0�i��p2I�5�+)����+vx^�$8�$A��R~i�N��3�3-�o9.|���� ���G�!�;�����n�6�mό��_Jh�oph��CX�sN}˶�\�t@p~��8��ܺ����n�342�yX�@hm���#�a��7Ȼc뙗�%c�e�|���?��Ffl��'T�����T湈��}�愅t���&�����g�d��X�B�֐!3a�x~�&%����	d��F�j�n�"fZ�I>��Gh�q�@��X�=��q:"?C��7E��q恪�OWe��)��RCj�)��,(�]S�#�$�bQ�j ;�Z�d��4q��D鳸�jT������=��5�{gcٱ�TF��l��ʞ��8zFB!��*}��qBR���>�M�v���|��F�@@����7���kW?u]-ߩ�G
�#�1X��ym/��=O]zM��ݭRÂ�f�3���S-�֏� VN���L���Q��$�AhG>Q��	i�ެHw���W�1�=X���&�(](]���!/Ӡ+�H�]p֛OҤ���|��p
:�䗌��O��깍A��^�5�E���LVG�On&,�� �0s�^����z�:>�'�!�Ⱦ�.�y$�1���:�2�iXwE�;�zR
�=ҙ]�&�����Z]�	)���Y�4S��Z�|ˢT�}���$ކtM��^l�Ǆ?�҆t��Kˌ+���<��	׷;I<S�\��%�kj\<�gn/����~J�p�=p҂Xd��+kq�n6T��cȦ�|q�@�:S�W�H��jH�߯�̌��3���p!�5�]�.��1Y��4�	<��@ӊ��.��#[��yp򐽜�:Pة��[rl���� ҧY�bx��#��D�;J��Ӛ��$�qY��ak
q���΁z� vB�
`��$��ۂn�b�K��J/��*��ǭ�1�*��*e�5:L������ġ;jX)�k5+�"�(��װj%�$���Ph2��v��m���Z��p�&��p��4�lĐ��W~�bI�T�R�jޜMb!�%^7�y-+`�������.X�4гE����r������Sǽ �����Q�m�A�E���/"͸M7�"q���f|Nv]3-]㈜v���t����Ⱥ1�l&���.��a'��6#.�ķ���>|��g�h-��&/�ң�\�uH����1ylW����I�GpלJ�ГC�~��I�[�]�`��U��a	G̋�R;��j�C�-���]�iJW�3�1���
�\�3iA\�(x�� /��ܔ��.�8�:��́��z\{���X˦�k�
���9���|`�7'�����D�ƹ�#ȿ<���QY��s�(wm�/��:�U���wAyq�����W�A;l��$���U�M�f������aM�k}�8�$���i����ۦH ɏ�(��[ð��̾2�SV����c/@լ�s���!m2��'�{��i��Q�t�a�r��i��(%��2jчq�e���4x���t�]�f4�<D��Z����L���F�a�Jѫ�?%���~�k ꛗ�r&'�� ��Ls8��k�,����6�S�E6P�<���O�(�Qi�VMS.c��]��OD�*�*��L�[����'߹���rA�	B���m`= x��vZ���Leq�)C��Z��:΄���6���t�~��8�M�sQy�E �ǭ�~�tpD�����K�5�����i��cv��9�����A�Y��~�oT�� �}8j@D�e�B� q���1;ɟ����5D�GT����r�TZׁ �X5�U�}X�c�/# 	�6
��'WEuMJ(t�����)�~C��1uW�k���O{{����^�f��.b#J�&�cb,�`�|��&�g��A
�n�z.�8��=@�7������aNx���e+r���2�\���>)#=��8��� E`��y.����P���N�*f8p'[m;P��`���}�VUQ�])83��v/V.�d����ۯIr�.Ϩy���a����+�0���?�y���h�r�/� �R���J���S籱~㞇k����6��F�!�V:�B=���g�_Y�R 3��e���x�)�S���<���W�W������Ҋa\��C���Ҟ
��A1X��H*�D��YPGe�i ��D6�H��%lěu!����lR<Dx��1�;�4�t�^V\��>�T�u�W��6g lD��8���֌O�V���.��Wm�i��i����8/�~�6�����5��'S��������NN����'�İ{�^k�c�A����l=�$�X&� k��_]-	���d�㙩�n�X���.�̳�/��n;��!�3�Kͮ�h,ݜ�<�J�P-U��QrW݆u�5׬OH�!���aw�#)��L�-n}�g���S� o3��d�R���Â�Z�������6	%�ݏcB����B�������VT$�aJS�y3��2RQBg�JL��ҹ�%�d@���
oWBH6s���7O����>K����+R�
s�߷z�d����4��>�/Sp3wZ��+'�EF�f��YƏ�/�[�lq��~��t-d/�2��.x�b��U��Bt@5���
�+Y�(.�mR;A�$[-;� m�d��J��n�.�
��Q���h/�S5蕫�b��HC&��t;|��Ň݀N=k�"�H�ճ����b�֔��?mE����'*����_蝩�eo��v=mR6O���AG��g,����[��2�E�<L�1ۤ8xx�߮���r�����]��`���λ?���o/� ���ͦqMڴ�BA��w)h��="�G�s=�4){�O��Ulb�_�D�8�'�L �v�k����6>�G�n�Hc*%U��(�ITV�������p!��ϲ"!ŋm�\t-�c۪���LZj~$n��ah)b�6�:�I�G�NJLˮ 8i��.�6���u�u��7j�����w���RB82��O������Si1�x�4 ��٧���e-k��wg���`�x%��*�����i��~QA���W�+��6f� 2�ΠɁE�R�9�� *B1"�<�\�&���,j���T�1��3�^p̅��dB�rزE�r�mB�������
�o�S�_���G=��ehJ=�vl���{�ˤ�w�Á�z�I D�^
78�f�轉n0�����s�^�: xRy�!kT:F�_�`#e�`�!I>�'�,��fB����d!��-�-� ��pm���k@`�mЗ8\H�o�`��kX�~(�`��9���kؽ~��oQ�E�%�֟x)�ؾ��a�C(Uy��y���y^�}�n��6�8� &:�%�N�1�ٰȦ/�9 &�u�[M�A�x������v�0?���$\y|�q(Xld�e�̵rn���4��8��|Ǜ��f���h}�/�\�o�����-�3�(Hˊ>��G���[$����H�uL�	W����ݽ��ͮZ)�uޢ���p��Z��~e�wI�����8�{�$i�Máu���V�jQ�Ӄ�;�Z<8@�w�`����&	P|��CYdT�p���ڗ+%*�Z�*JP2��G�v0��z���i�aݔ�D�Ku
+��w7��4 �o�vK
�2T��RQ�;
�N%m�PUt&�!���t#��9���Y�9��8��i�&|�[�L	8���,k9�aN�7��2k��lP?���`��t�$ף!ѯ���P�s�2W] =������M�bGm�9�E��?�T�3�8�`�9|\"^��)�[�Aӟ6�i�qiB*^4��}�e|�w��6�G��@~D�6<ڇj�������8g4P~+[x�*��@V����m-[6Ĥ��XT�����\�s���ά�Fz��%� �|p�����L���kH�I2Ѩ�|ԁ�[�a*'	�Zﴁ]ۗ�F5�&�nϋk�E������uLi��f�u$���i\)��f��Jz�#:82�܌T�Q��3'?�uA��o%o�	�z�e	�Q�}�S�@tl�bI��S4q&R��-{�N�3%���6��i|c�FG��(O��X��n4):��n��};�� �.;�h�.��>��N����͈.3���D7�7�x�fN �\���A�3=ZK�'�X���p}l�����p��Jӣ�e��K���\��k��&�\$U%�$z�f���!����i�ohCeo�rW����0z�
g��� R�#�Y�OJ�����]F�^Ȓ��ي�!��Q�oQ/�j�F����R���`WY�&�l�����[�=�!��+"����� ��D{�<L,A:j��;|�yur+���֡���I�6̽�@�����Z��kx��BWm�z�p_�5A�3�\����^��?C�J�8W@É�A8y��Η��Mh*B�0�gMo'�m_�yߐ(#��zg���=;؋hAI���ޕ����h����$�����2�-ū��5�@~���}�SA��:\ǧZ��T!�zw�|.,����ѳ�@ڌ���9�1��u«�r�y����^I�_��ʌv-��Oz�p�� �pT�<B"����b�A��
*^.�^���ׄlxU�X�i�
��[�n������k���Q{���B[�{��C��.-�sp��?'{��t:�`�P��I���uol{Ԭi��!ϝ(3\����9�O�	zv�W��X*`��lF�	�vP
�5 ~v����G���ݥ�\e�ܮʒ�念L����m�5�<B�}��A��$�����<R;���7 :�:��GN8T�����U"���M�u�q���J����)�Y�lA~Z�u��B�9)�ܾ�YZ��@B��R`3����۸�N� F@)X��_��7eӊ`I1�[FE?{�������dz_�ܩ�,�Ƨi`��~�����ɴ�O�%��3���k�HƠ�T�Wɲ|[��&B�:�%+%7U\;�;�!nN�
$B���<�D��2K���h�l��1U�c�[���H���8�����:�D\�Gf�إ��=�2BOͬ��!�v%?h{ԏ��dT�v:�����m[{���t�:/�"H�rK�D,�Gn(�P׸�|ʬ�?��/��=A]�l��J�����ǐS��+o!�Τ�}H������X樸"�==7�$��39��«5���|]F��ѩ�	e����,�v�o�G��P��SW�ͤ�A��ć��rh�z�>��+��΄/ �h�&!Ps^Q�:�ϟsɩ�:8�YcQ	O�u�J���\��s(�������NW�������ᾳY0�M���MDt�k��L`"��XI�.��{���b	?�Zg ���6[X�/�)�w�d�����L���<ֈXw�����P;�K�)��40�O@��H��}kf�~�P����SYg�X���M���F��pEo�Ґ�Ao���-,���s3d��a�E��LDC��>{�`���sS�tu���]���ూ,��~ċX�!0�����s��L�ʭ����x^�����q�AMX"˟�̾q�)/��Qݍ}30�DOԸ�z�8�2"�do{_�CT�Ԓ��,To��%/�*8:����1S҆�wܳ�:Z�����<^{�Z���6�(8�� c~ɝhB�<3-�Y���G�,���F`���ij�ӆ�ط5x \0�uU��um!)�w^��7��<���Z�Q�>F�`�\p6%'j:e3D��~��紺���w7�\�""Y��u]����k���97���ܗ!�LXM��G�0�r�e�Bhௌ�MNp�
�z�m�ި/���Pcw~-�B���λ���5��Z�jn#��PFK�z��d�]��V��,"�8�?h,��:̢T�T[��0{��-�4}� ś:��nX�&�����+P��3P��o���ˤ�y*��*������;H�dˇ
oVMA`w�z���n9�~�Z�@8��ק��g��t����̎�%_B-�@n���G���[.a�.��1w��
CU�C����c��@o��_�`zD�捂�j0���a��!~�U2�:���A���:������ӛ&���KȩmPp���&?^:�|�B �aǊ��^�Mz����]E+�:H���MW�`�X���m�f��w��PP�gC�E��'����|{�7XV�v�/�'�sǊ��֓��~��	?b#��@|30�ۤ"���҄��P��8'�#y��Tf<\)Dz�1d�$�ͤ˱�W�ͱ�_U��᯶�* N,�h�X��º[y�&[�0���Euن"�ʟCH�����J��?ɥ��{3��{�����H(�ߦiꌬ$ \1EbS�ƛ�������64��h�/�n4�Yea�ěz�3�4'7�)9}�8_�S/�SEG����G�*+��͕���4޺����m7�}r7|0t��b泩	����g8��R�0���n�M����}Y���&���S��4�݁�f3��\0A���@�3ЅHy���,�?�߈����FH��>��_*)8��O,Õ]蹝Qo��V�
��usw���Q��V��N�J�� �7�5�)��������lb�_i�6��uUV�+���!|�}�mEψj��u.���Y�w��,�{B,�O-���^��E��\���p[t1pC�ސ{O��N��zA2�9�HPn>�m�ߊ�v�)U�~C��)H�=����	3�-%M^0�H)ݑ�y\�;�:�)�h
����K�)M��ǐ��Փ�9�Aۻ���CQ�W��� �{��6��W�n��{О5��Q�ޒ[;i�E w�kC08)�u�.xA(*��&4k=I]?+Y��I\2�|WBH�Z$���Z���0i�.9��FK6���)9��j�ۯ�T��=o\����F�"��,X� Ņb�����~s���ʈS��b	��B=6�U��z���`�Z1,�#-���d�S��M<F# ɱ������"�R`�	��Kቬ85jm1�/F:�QBt�H���8�x�Z�Q<�A�Z$�²2�Ta�*���S9ٕ�7G���`,��L����t.�H(��^���:k��N!m0}X�S��l�����Ӈ�Z��t����,�����0M	-מ��X^�`�- �!F�Yn�t����~�Ma�ĺt%r�2������#���q�u6���-���cy��V�+�AO ����ËP���'-'�y���|mJ��������I;�DQ�h�㱇�t�G��{�؜�����t�,��K-1m�Ծ��N�׫
��կ̟����5?Ʉ3�>�u��Ttt>P);��=�K>9:o9o��E�Qr?x�:��Q�eܶ�dr�3�D�k�^g�~(	�E�Wb}�
K��͓��f9֙�,�$R=���.���;i����q����k���-c	_vu`�i ��SÊU	_$DOJ���b�l�j�Rs6�@$(��Bw�������:_\Ԏ\Q��_��U�G�Ԧ#g]�P��W��"�e�`�sw�l,d����0��d�h�8���#�7���|��9��A9?Ȏc�=G��P�!,#}��b����f<譺���p�_tx���$ ��O8g�D�ws�X��I�vE���퉠�eؖ�娆�Q�.����i�H�6Y�N�Z�ş�gjy�M~{(ʪ�c!j_;��[jEV�`kGW��"����,�Ѧ `2'�p4 ������}��HW�$��	��D�΢�?ze�
�Z������ �0-^�)0���C���Ȇ��B��w�ߙ�(��>�^D2|U_6�T>�B���t�ôM��ԒV�(%Y9�/F�҉h����̜J*m��G�sK�����p8k����IN���!����r]?M�j#@g��=�G�r�"ܶ�ɴB����0De`y�ߨ�W�C)���@�ʗN>���y�D{�{@����^�J%.�q��K��������~E�Ix�w%� ���BsIvt>Ӿ���Uֽ������:��w�&�;)�{���
�Rӵ��`+>�m��t���wέ�Ӹ�~�o���	�8NX��Za�8D�,}��Gs�儬v99�|�o�es�}�� �`�c}S�\@�	]�G�ٮ�Ȩ�a�c�o�� �f�~��t֩%#�[t��4B[���A��Ul��C�ż��͵V�Ae�|���i-�>����)'��ߑ���Y.i@���3�K�����x�߱��?=�F9bI:J8�.�lg<�_1����t+^Dr���~��z�7�����7a� 9ϕ"C��Er�iS�c��*|oOAŸ;�B�?��ȿ�U��~�͕o�9��bNM}*"�Z-��T|q�9-�/�j܀�q=s�eBа�:��{��p��:=c�jL����݌����%�_��v��Ƚ����2D�B_�e�;�Wt���>�l`�q`�2���1��ÌWjib��NΣ�rkJ�2l��wc�$'�.Y�P��A:��p�n�)�R�_����/���iP�[-�G&'��~�՛b3*����E͒e�<z��?I {dD�@�(���Kb�����@5�������Q���yF�ML7wg �Vvd�����@�(�j�}�4�@PS�S
͞
$���0L8�c���D��9F�X�*�(~�/�h���N�S1��]Y:[M�Q���-w�3�w!��\^]fC�g
��k�JQX���d:/����/Хgx��z����?Jd����t8l/�v[	�8�5G�4����
��������l�sZ\�NЂ8X������>��O�G�/c���|�_E�
���]hX�r�g���j]��B��#_Ti3��q�* Ć�:�5��?Wn\���˝P�D���dx�}�/�'��2�vV�]Z��P��C�JD�ŘE�zpm�x!\f���pnĒiC��:ƺ n^�N�{!��y [���E(ݬ=�i�����Z+�~��*V�S:8���zẑ�y�{�|��w�'��a��HU$$���3޷��� ����s��ʏY(0`��>�%�	NV�!�w��
� 2"[��@��k>Ku���Ò�7���G�Ӻ�9�����r#��V��͠t�dx����Z�?���$��k�1�o3��~W�(�<����<u�&���\:�zPZ��s�lj���פ��Z�/���9�ơ<��q���TU��D,(bҮ�dI�SY�*���u7�D��E}���@�|���6�4���v��L,�"�>��@F���Ř!�B���Q�37��e9����hc��-�uxD��%��J4X��4����-�>�u�������g�%%�ד��W�Kǿ��y��ȡ�YU��P��B�%K�Ku�|�"�:�<��a)x5z�㚄yk���Ί9����/��Z�O���o�~~O��9�x�� ��p=o��|�����+����+X	��/��$mAƆW͝Nנ�<��9&�]�K
[��W�V��4��:v\�8L���vm��.nNz�[��u���ݫG`>�����s٪ݗ�i$h`�8i���G��i��`~^�<���F�ծ�9{]K 6�8`"��)ѼYz�8��C	<�s����Kvf��K�� o�_�u�qv7�2oFn�6�"ٻ���񵵂�e������FJ1�42�ĕ^�n G\-3���H�"	�����XM��/[�~0Y�W��4rM�"&#l0-�&t<�q�d���O�!2X0t٩=r�epw��F���=�FAv���OR���l'j�v�Ѓ��,ḽ�Dq� �礣� �l0��9Y|�(Hƈ��������_x+>aIԵ�/ꠠ�)����Z�Ùe;����N�)ױb�N�X#L�Uad�s�0$��� ���t�n�w7���ݬ=�a�3�B9���FQw�o��aG��G��Q�	+��+8�ϙU컾�uJ��_`�/IOo����n=����R�G����&����R�����	�|���:�|S�m�?(��]�(�H��zÖ�,$䤤��(����.�'��Z�7�I�1t�리�O�b��rଷ9H�l<OLi
� ��ⷌ��7��7X��V����-��i5�H���.�4�/�Kஇ�?��e���cUA���[o������7hޛ��í��CW|Ħ;��椣,)M�t�c��jS��zFCCa��a�J.X��g1^�ٝ��l�Ov�W(����H�r����U�DX��7�5]~b��K�49x�x<@�0����:_���x�����U⺱�d�k�}��UkT��k�xw��@�i�׉�4���=>GW>*g�Z�?��]��#'��j.fE�g������%?����5��S�cƿ�$t��ru��?���Q�� F�Ț)nL󒤣K}['h���	H|�>Ж��`��>a)��B�f>��<��羓�QZ�q�DzZ�U��;��:Lu�k0�mv�R��Gz3��# :�Bf"�y2�ՕhLU�*��Ū�Q�QKQu#���x{jo�����~�4��EĤu8ʣ5���|L�ũ!��3�ߟ�b��l~q�z���C���6Eb&V�z��%��r\-��� vO�Uͼ�ULJO0�8���
�E#\��`�)��`'׆�Yv�<2�	�\Ӏ���ؔ�v�&�fw�S;��8>М�PN�i��}���Š��鲀�Y`ފ�6�I�5�mO���7I������� 59Z#ʅC���/��_Ɍ�˿����)v}�Ǌ�껞�3UΣ^߀�X�xa�ņ���wl�;�U��-���T�[��?;U��>c�R�Bfq2o ���8M��_&(Z���h%�%#��˧���0¿	��DLw�@0:5s⮦T���zt��B��<�W�YSɐ����V�2V����a�Sp��)��P��Џ���+!�s���j���U�u���_�UڶE�����$ �k1m3��*���g΃��(\K:�Q�dKKt���t�#!�9��zչ�[�]�!�s�t�Ӌ�΍�go��Z��x'���l��<`�ߠh�_���^痏�p�X6Vf�
�;��8�?��IG�];�E���>c����ɽ@�HQ��{6'��#4۝������;���Cw�HV��� �����;�Y��Yl1����3�Lr8[p{lك���N*��1��
�C��bP8����n�d^�\�e<�X�4�7X����Z�v����½��{�+L���
� %�8<je���S��NqHǖ�?�#�Y0�*k�ݍR�z�8ғ)�o��1s�*�ϭ|Q�XTP�s�����ea4���[�3��p/\ 6��V+jʕ�M�\��-�����n6ٍ ��JQ���C��v�|湝�ay+��n��d�W?Zr����G�bgGd�;2r׆_h������D�����	���к�j�D�	���vڼ������wȀ��nv���d"]�	�O�(7Ħsd��x��l<�N���-��;{�Ywi��=պ
<��r�C������1`}*�6Ec��/���jJ8�sʷ�]���<N�8�8���g������5�e�(�z���w��W׏�˽	��O���X��`9(�;�H��1��a0�-�Y��[��?P�k�&m�F#��H�3C���bS����Q]�$zM�e���qt�'����	�P+<So�$l��)܆�@(T
ɜ���H=Fb� �t��P�2�;W�q���иQ��	���}?6I��Ј���?V�~���	 ���يXt�H-~kV�s��.�r�X��/9�Hc�c�?ۈ��.,��U���� ]�2!X҃�6B��PG�ר�D�Q��Z������S�a�
+�� Vu�w/=��Nض�>Z�H�o��f�mlz��$BlaaR	�& ���X�JK;w�~�7GvO=��60�S!������/�sLW5�l�7o�1�~)��������:�Ц=����H#�d~p=V'տ�mV*w$�h �c�	���׶�����|��������� W�ET�l���A+5���Do����F���U�mי���`o۠�4W��5��<)9HC w�l�}���j"�t���6��d�S6M�Fם�l���T��Ƿ���2t񴜅��X�ٍ�7S�N�f�@ň�Z�y�Ra8Z@p*���������m�3:_➜}��s[�+C|�h�����=�X��Q�M"�56�% ��t+m�BU�gp9-�xa"i���^=?�5Q.k�#���2��8�p�R~�fc�@J��*�j8$hC�C5M���xmo������"R�[n�qF^�mM,-��R�"���U���i�AgL��B^o)���r�r��	5�|8�Y�;�Q��]㮝�1'u���x��"��D���g���Q��Lci��Eeӏ/�j��U,Z<���̏���C���KVr{U�:߂�hm]!�|~�HƊ�?��|��sU3Q/ֳ}]~=Q �����~�ӌ������hsՠaU��Y�0�H�?�Ǽm�}����Th����:g���^˹ �k ���Z��v*,d�娖{�خ��=�_���|�*�s+�th��ҝ7��&_����<t4�NB��5��m9�;���ݍ�7	m�^����ʟ��[b����%
��7�� �@�j���_�E2�L��h�
���w�o��M��GaG��@���Z�}�# 5��a�%.7�[��0���l.���L�K�q+iX�b�i��|���0��D��]��T�j㴦��t�gO�
'�d�w�i�n����gh64�o��c6ڦP��H6��r�D�������˥�&�SU��1E��>��֕�߿��L?D�h�� �@�Y1t7S��@����|��Adǡ���I�L嬫|M�tR8H/����r�n6���81w��hT��:İV[�8Wj&ۍ�Ќ�o���Q�e3�b��+GI}�:���������Y��/`���-C���d�����a{B� �N�V%f���c�߃Wk�D?F\(�>C�*V��䫄Q����y{�K5��3�M����Q�by�K��jY�Yll�^��{i�׌0g��H*��즌��b��M���O����å����BÂ��x�J`� AZ0�_gn"B;�֣�M,�$��	�&��5D����]�ͮ�L׽�)$B"n���J�_���e"�F�@]��@��w.3�R�:�*���A䛫ߟn�V�?�P��w?���q泧i��q�D��T�J��k?,����֭ Vog@�c��
�*d��)�$3�#&L�y�r���2��a�����l��VN+�M��jd�a���F>��8y�JF�n��6�60P�/_��<��SH����,)6A+�/�l�i̘�e�'�#xxlJB��]�m����<�{�Mo_�!�������1`'-(h�^ʜ.�Cx7�8W��:=��c���'���u�B�Q(���ƺ�}'��#b�_xg@����Ï��^������}�f�[���yr����	��J���@�)^�eل+�)���A�Qs^=����_�u�=�V=�O7����KIٌ�G:��J>��ҫ�1��f�?'],��>8[����=�aϠ���d�ʿ��Ecƙ���6��������ʜ��7ӵ"�ΛR\����
e�H�&ŉ�f��v.[u�Jt��n��T�+x��x��P�D]U�Lo�H����	$\�'`쥚���{#�ʒ0�W�r  o��tAl5$m����ȕogr�+� &.F^3��<s3�V��#B:�Wk8�M���Y�/\˿�܉�"�5̴n:�MEG��2rA[;K�n��:�UR-^��'j��Z��"��
���׳���}ד�����B@���"�k�?�Q!;^�ʽ�,?�ȽE`~��t:!3�z��S���_�Xd�J�r}�ˣ.��B� �+W�5hd)�S�A�sa��b�"� ��m�u[�\���������)f�z]-d����	G�W֡uE�;��<�H��XJ�6��,�HG:�VJi���ך$)n����q����e((��{�Ï�QJy�O�3?�&0(�h��w.�R�W����PTQ���߭`�3?��v�F����.,���l˴큔
X�ߜ��M>d#�������]�A�r�ݐ(�T�6�Ԍ�6)BS+���H��*��y��ui�������&��7oV��l�n�W!8������53e�	���<L����gP�S\���,�5,����(���*��9�I�"�k����������MVw���<���kj���t��q��pn�':�ێh!��׺��Q?yG���2F��"9rN-��k(��bA����<Jڳ�p�,,J�ytd�����>8D?k�q��i�������3���B���c�|x��ݶҖs���x3�]R�J:L�Z4r'� 3h�9!_�9s�?M��Hl��<~���,�,��珯�mx�\����!I��_���Za������q�i�]Kɵ ���Џ�_6�#�LX��Aݧ
N;Xoy�s�8-晍��l;ژ�h!�=ԑE�k��_n�=ǯ�ȹϼQ�t��/(� g�b�D��y�+�|����"A
�~^���Ġ�,�
��6��U�z�C�<�V�����%���� ��6dd�gV���	_�u���,�tE?�s�|v�n�����5ڑ�9��H^�)���A�a��<�Vׂo�6*&V�'������R�n���/��觫Šs@�9���:�0�#�!Ɓr�(ƃ_<��zi�^���x��1H`չw3y�)(|BZ��!�s����t-���M�/\�!��:e8�l^\IkT��u�Ο
Fk��UJ�����{I�Q�O��<�f'�vyO�$�O��O#�U�a���Yf31��=�B���=���I�	*>�=��h�0���n2�n�'X������wZC=��G>8Bv�N͂��cpO���`4�¸X�6Y�U��+,͑��mMo�)�C0��WSے��"I������X>1����	��V�>*�`;W��!V�ta�^\Ha���t)w����vyG���ѧC�Z!s�ܦ�h(l�qܸ�<.����Y���"�1 �Ա~�=۷�LN9���@	����yԦ�@p� D�)ބϯ	Ջ����a�l�~O�|�FŰ���#��e�n��z͂�b���,��&�2�?�xP��V�-��T�C��i���5j��T����8N�|>��%�*3z����T�!��S�Eo�	.$)Ciܯ#�0~+�ϻ�:wxx�^cH���RJ=���,�d�`��g���0) W���">"��'_;����"h���1�-�M�z��1�c�Wzu���?�l5r��>�,!�_�i\9��G��ߩB,L�6�`W�dI�u��YmL� iq�g���C�E=���z�j���gB�U:l//oF]*$�ٛ����`�gn Th��kN��ןT7U��^KV�)�G�o[��pci��:>^q�������}�K��O�����P�6����C��W>�w~��C1)�������f%E�ٲ|�g���l��(��6B3�@�?��o��1���[dAkglh��
gv=��f0�0
�/�%Sx}d2�kVE��y������{i�Ѽ��+�}R��4��{�9B��(5g;�5J�RO�v�~t~{ޔ�N�����/�p�5}�s�7CU��j��)˦I�N���������ar��X�#hÏ�.M��C9vtcf?)��'�k$�;L`�1����жjZ$gh�
��K��,�H��Jy�Ԭ/�=�;A��f��yO��#7���}B3a�j$x�ئ�H3��}�[���J�^D.���LwobB��^\J���	�;O�;ź*����'� y�Yr(���(���C��K9q�^(�[�"���*��^��x�[d�em~��;�L-�A1B�,��(_�2�TL�h��ϝ��;p�D�R���� �H�^����љv��)m�86
s���p�n��*"#�Zz��!�FW�3��hT�QJY�,��/I�T��|��� ���깔��ml��6����)4�^�͚��x:V�zW��:$G�O�.i��ia�_ƈ՞&���% 1B9\L��r�>�d�R�)R�Q�D����1���g�&T>Ha�)�X���m���V��)ߓ3�.�u������g�Zs��:�����e䜱9|��Z��A��?ad4$)꾡a���|F����S7p�R̈́�t���'i��\��Q��p�~�0Vˬ����w�9M�dͧ�P�n�#Mx��*f�袢��n����Ί���4�9W�Pk�$Uf�;�3�0$�*�������R����B���`�A�)�	�GOǯ�5]&��_�в3�IS��A���|�K�b��z5�Ȼ{�h��;���4�.�?���t��U��NxHT@����j���^���kϩqPR��=8��3��?SR���C,�Rk����S����8uR��W9�JR�T��"�~_�N�V=���@Ķ!5P��׏��b�2���c�d�H)$AQ���Xrp����BBM	�I{хj�j妦3M��N�<����3�	���h5�^���:�H!�]J�k�X3-2ĔM�7���ע��<�܋ֹB�b?��	6��/� ��TEEuZ�fQ|�sEc�A1f���G>�HZ�3hucd��t���xC恆s���B4m�)��v�qvo�03��2Y��VEN���Ϻzt�ؘs���>������o�\wD$2�]�2B1}��Kw*�VH�Ͼ��H����m�F���Ƕ9�Nڢ��T�1F�z(�x�Jd�?r�������;���ʡ�5�1��ٜ�Ԗ��}>k�A�@�3�]V��<ce��ry�����C�f3���}���<?5C�Kq��nC�1�l���U��0�zQ̫s�1E��IB/�3P���Q�f�G����8p�z��Y4J��=��N��n������RJ���gҨ�%-"�\�Y?��@�o@��?������{�xd2X3C�7҇]�*��9F;�lVڏ��1[��ۤ@���X�;��_����!�_I�I�d?��1�g���Y������Ҭ*)���ٝt&�Ѷ^�au��Sw��5��j��7J*�٫,�,��DQ������U��'v�j5a�=+����=���:�I���r<�Coʘ6�[Q�@k �Y��{� r��fK�-�Ż���ϋs�����kc�G'G}�������RY�{�!l#ܔi<�>?�������~��L�r�^h�����������~O+.K�7��?��נ3�i4I�����4���ތe���%қ��'�h�d���.2hob�������m7���7��>��,�7�,��wO�>������8lE������OB�q��%:Y�m���J�R�*\O��_�y�1Y���g���*_\�E�f-א?�������:�!�ԍ{�����ekH�H_c>�����j�*+�m=DX�O�_��>���} E���z��r�p����H�%'ȏ����aT��@�/5����wY�%p0���"�F\��.'���[�1���lR �B�A\�}�����9�9��@�U�q�8ߧ�E�v�����Й������(�>��B+Q<g�U��,��&����w��O��E����zա�P%�?k�]���׏���1,6u=�kɪ����&bc�G�g���Q"���}�(�)��\6��cX̊�=�>X��G�l�②F��7i�;��~e����6Q���z⼄'^"��+%��L_���Nivv��ԅ%��\��F�������-m/��v�%t9�'ޫ��#�3�g���Qf�B�??�Z1����0Lo��5��������q�o�,#N���#�RRGҗ��7�w��9�<[yE�6)�g5�,ď� (�Ӧd5��ϊ|�S�Z5�<f�<��E�p�FȧSIa7Fī���3�`�
私�w���"�"ȕ�����u�i��
d{�
���4�wJ�KX�����;�Qe(���2�Dk�<ekf��+�oɃ��S�����q�j}�A��T��pFO������	�w�Hя:����xC3O.Aa�P�bj��E�ϯ=���f�Ml����/#9>_U: T�s�ZF���y�b,�ɱg(m��������f�]��R2p��ۏ�֓�`��ԧ��{�G���~4o�'s�'������K���o��.@�nK���O3녷x˧t%q?�:Ϝ����e�?�T���dw�04��c3�i��W�蠧����`,&	P�,-V�`w�9��,t�2�aӉP�Oެ���$��ECʖ"�k٧Tn=�4Xdq��\A8Y�q�wt�,8M��p=k�{�ş���ӭ�5�m�Ek�)̱.1����$h��D.#�?��>:r�>>w��Y�}v}n7�&>@��_�;�]8A�5���g
Z��9��K��R#v���ܩo���a,��f�V&�L�o�=Y`�|`r�\;ٱc��Ͼ��c��s��Z�H	�YS2~A[����M`�0�5.�o���"P�5��]��@�kY%%��M�V'�l��������sz�d�_M�<>�n�p�B�:�r���[�g�0K=��[�mT���kk�Vb��P_h�";��H~��*&�9Խ�Xݓڶo�Cǫ��Qw�4'���,J;�|#`��FA���A0�~�JM��g���(�#DF�75�X��Q#�i��~��R�>
���Hl;?}R0�	�3=D���p�� �f?=yc�'�_ �v�\\�QW�?�-4�m���r�K���!�@� a������ S�$ NDh��DX���uWܱ4�V*m��E�C����DN��u,็�f1��U"�7θ�]�!hx����t�dBT�.���rIh�z����Y^��PTRV%���IkH���z4m�-_l�]����$n9� Z��@?�N֊$�}��˶MAN���
sL��,�1���Fۦ����8N.gGw����X+'d��wc,���mS[�}��T3ٍ�V��Ǆ��=�<*PI����$�4��}+X�Z�^���d�o���	�샩�3R���#���[H�LU̵���#��%F�hM`���OK�x#ٙ�/���J���E�X�}yHXf�^�u�� ��i3�,�Hׇ�.x�l[yR/Q��ouq�{��Fl�w�<�<ܽL_�?R㡚���SS���[�d>֜���?b�)i����W/�Gw����EA��B��(*��ΡE�\�%V�$�p
��3�od�t2��j�jzr�+�����m(̀A�`Ef��p��A�9x�J��t2 Fi*�i�����}6X�C|Ɲ�|�C�c��"�ny�J��_��S_\/�5��60`�Eb%��}abW���Rb��fHv������3ƯD��Z���se.�Nl�R� dA���,���"��۩/>#�q0d�+��;�C���}��ڣ��͒IV�c4�v�I����c���m���G��
�#�$��'��ө����\�"N#��%c�%JkE�b�� |y����? ������u�&$�?����<N���i�a]�L�������������I�5Ӻ�#���nx!27 ���O����kT�Q����V�
�8��Z���ot��_�o�� �>�6�����XR�XM��2;w��`J���d%��۞��p!�̢��Ti� ����ײ��u%���1D�ܒ���3
K�Ft.�-Y���x?sB�}=���0Շ"rTĩi�D������v�2!������Pe�0O^������\ZH����;M�z�9r�7�blgL�ݙ�2gh;�ÏP��z�� ��9'o����1f�	�^���%�jن�Y3D�&c1���^Q��G���XiS���3���-���;�.	`�ө�󅱲cAg{P�H.
� ���8	+�[@3�ވ�l�I�5l�]�%'�i`��V���E�f,)��B�#m�*�"cuuo��z�%���o�Z��dF"ś~�tnKW��;��Yj�{�����4� �{��A��SN���#|���<�*�o��/̩0ʮ��s����K�3�k���a�c���Y\��4דX��'	����J[�M��R�W�H�&ol�k�hQ���Q9C��.ִʪ迺:Y�ߴ�۵�i�Y��މ^V��kA8� 9S����$�ab� �ڙ]�7���y�AW�%�C���~̩|���`a"4E��*�]N1�ϕ�@b����O�\o��F������q� 㼳m��a�����bGo=��/�?��v-W��[���1�����k�����ǫ���O�vI����fT!6��~mM��,S��D��
0��.GI��CzgF� �m�(.�~���N7�}��[���*��n��%��yv}tc�Kv�x8-��Z~�pC<B
���>���X��[�¿ �<����K�v�3��r(�b��M����-�QsC��Dg^?O��ӏޠDj'!;���|'�B��a#9>�J�l0�~�k���(�C}��F��
��zg��Qsj�-�h�S��q2�f��1Ȣ�.����؍u��*�/H���ӕ���ɫ�i�����Ss��$�?�P�	F�E��Q��r�Y�����$N�J��0.K̉�!�k>����6����-33���d#z%�Yg�F��'U��.03�g:9?���}��K܇��@�t�����jK01s�t�Emfz'�㲍}/@�*�w�!�ZR������	t�C�J(��K^��l�~U�)#t%Պ��f��#���>�'�����ӱ�v�.:
����D�g
�y10P��
��^L�q��,�y�����j��p�����4wqQo�c���)D��{3(�%��$<�Dd�;���R%�}`�p&IoÛ�h���T�0�<�"WM����mB�g��A0�5���Ȇ댱��֔�܍�2�պ�9�>"'�h'|{��Gm��N/8=�	ړ0`�,�^��-b�j�	�w9�T "5���P�/�G�T��C]k��������Ĭs�F�EQP����ۼݝfb����� ���K�'��割^���0oNC����ڑЄ.�ɝ�c�ha+δ:yS�|�}P�VS�ց���`b�W��dS�%���%��� F|}�~�Y�q����	7yU�R���ü��.F��a/����yV�ZC�y�*�~�*2E���9�v������%���3�TŔ�_WD|0x�I/�߃���(��0��o���V�j�ݔ4M1p�!�L�(*�جq~�!�
6��5\g~˫F����#8I����\��q��B��8��_�і�f���~X1��_w�(Ou�fb���D��aK�P9ɝ��a/��ݻ���HU1�o��w�Q��7ON�
NZ�RJm*ŀ gP0��_7�Ћ?�	�%=�wz�#�}�7�z�mz�˸�)bv4J�Z�9m����ן��奜�����5�@�"h���<��&c������:����c�s��=3�Vx�o߃ ms
�_��ϯ=���3��?��U% ���1^�Z�U��08u�U"ej�O�	�����˧���n�ŰK�t�fD�{��D�X�ST>_gFyD�8���K?�_�͖�f������gp5C�ۃ'�k'��lUQ����e��ɜT���H�gT��1�[p�>j"�P����BҚo��	P?\U�Pm�z�a��2Yr��gZ��CL���%��(�:-�p����,h��2�&�i���l�`���1���tTH���s��!>��O�	-�DK1uj5����I�r�e�b�{��kKд�qa�!��=���Y� }|5��iA�u���֓��j��8����,�j�H^�bnT�uZI1���Z�G�㔻�ugT�Ywq)�^L]�Hv^���pěo��;�~x_u'��5� B�k���Ϋ�V�7����KOk� B&?�99D��Q�����3L ��{X�hyrV@�B.���w��wn�� ��W?M �0=�~�*S	X��|�mYm]w_�ڑ��u3xv��&�k���s����|2�R��~���K��+8D"�����&֞�ޘ��� �O��8<b���Mr���^([K�bZ��+ڻ|д
h/�v���)d�RCW��J�*t$�C�7S`�]Ɇ�q§�	�^m2 �9�\�g@�Lrj��̵�;[$��M�]��*.�5��+R�`���łsi%�A�V�
?��Вي��X +��RJ�^)��i����4/�3�@�~Ԋ�.���:���p���A1;6�M''�\�(Z�(�6�ǉ8�eLF�]~�����O�%��-��H�����a�=u�i�B��%��sp��܇6��Y+�����͇Ð�ǵտz��ﯭ�f�q��)=	__�RFp�(��|�v��~������8�J��JQ�]
<���x%Ѻ���63��`"��:]It�@�
w?��g�"3�)G�O�.�u֑��1<3��������:���[Cŕ�C�$�vM�., �bY�6'����\+C����;�E��1���X�Ndq!�xV���#l�d=C��a�S��E����¬����>V�[g�Β��=bڿ�yyt�.�!�f�х)���3�54z�`�%����ȭ�簰E(nr���%�bR���&s�[5�u\=(!���R��ϟ�'�y���F�v��_Z��N�0�
L��<�����z[�Kt��o����sY�"�XeV�K�2�"nu��mXȔ�M��e ��>�c-I�m�I��P���\�:'�����lN�v.�F�Eӆ�"�j��t��G(�Y� ���\��%\�er;��[���߮v43h�n,~G����l'��'C�w�l�}�#{�*Fl������|���}���G��ۺ���T�ED��ޫ�s�]4�ZZ�.�ŮJ���BK y�E�S���nb ����t����N��(��
_,rv��kIUsUz�j�-Z��hX��OC�> -��9s�<��D�֭�i)hT��H)Q�i�(oW6���`V+o�|����19�q�w�[�&��R��E�N`ix�	ހI�eWf��}3�{���PVKS�&{%���`���KA��zT,i�G@��*�4L����X�]�zV�C񦾃I�ؑ�[�Z���/Hʹ��5N�������.չ�i����,D�e�f6�M�Pg��\��2�{��s0���?�5̇�ۀ���rH���7
=qx����Js�Q~](�!�y:{�O�K�������
��_�@����+�6��z�!��"�E�6�bpƷ?V�L�]�rS�_^������C�GZX��AU)�m�	v0P��Z�ژ����ů��Ҡ�בG���P�3n�����S��sSs��.s?�` �Ņ�dv_(R*,I���t�z����G}���l�s;(<}C%GJ�a��9����f���d�aϮu��ެ��+��?g����V	��8�
�`&�7RXo�Mw+?��c��4B�ޢ̾߄ED��P�"�M}�}��q�J�/��sJ�;�kud��+���W���z=�WѼ�a��H>����4Gk|5Õ¥�"Qp]!�S��"��l>����dh���V�i����S��sU��/*(�椽c��弥s�B�h=h��O��>=m(*αM��!�Z��E�'�+Ҳ�s�_���QY�r=���8![!]�Dra����d+>��u-w�9-L�η�nr�`�"V��҄���d�Q�x�+�����`�$�4��n��g���Z/��A[cfcs��~���#~��[��0��N�s�2!�}Ӂ�zf��+�*���g��������m+��u�0Z��vy��|dqG?'����B0���:Z�>��+������#��x5E�5��j����U����� 9�'���Yj>�8��F���r?Rފ&��p�� ��_c�����slJh�[��9k#�t����2�%~�qw�q�x]x u(6lC�NO;����l�$�o�j�{�o�4�H �ǰ5V�K4P���?����Е�8:[��:ͳ� �\����j��wQ{�E	q��\#�ac9�0�"i	��O�[(p��l�[��1�K@����8�C���;(F1FS#t}�^{�X9T�)��M<� ���P%��y���XѦ�}�.��y��ח�.;W��-�JH=eb���EG|Qs�����C��,��s��t��C�h�FD����KL�=��Gs��B[T��Q��(�ֱnYK���������l�mA�K�)"�<���((ٶA�u]�0��CB{�	|~3�R�7�K|�j)�e�kz{��dP�;0%��c��]�3��;����I2�MAR��	�[��0�{������]�YG2W+\�!�Ũ6*F>�3P�3�e�����6oe���IegU��u�O�bK�rM����C�d�5
����~�~�mr먛�����QԌ�*G����x����Ui�k�V������-�j���;E��Im��eʘ}m�_�8��>( �瑃�
�����HwG{x�%����M�f������$��^c �_���B~'24��M�|2�H�n�mC�0"�azs�	5���f�5Q��/�<%�뵅��&o���3!�h���9�-���]��MqT�"�dF����L����)ꪛ�_��Ϣ�?������!�Ӳ+p��'SIOF���D2^!�E�m�ت	ċ;v�)�q�1��v�����YB�]TP�1�v���*�pXԞ����t� �_���Z�(/�GG/��%1`G�I�3��XFfѥ�K	����qz;z�bAa��7?pҠ؟no�:��f��'�@��MF�i[W{��S{���^�X�IXN-���^g9���g���p���a>�������t)Y ��e��K�qR���e�	y�������������ɇM�.8�8��0=n�O�\7��4Xq��#Llk~��`�C��|4�Qs[ӟ�uM�E�ω��䜞��Yb�s�@`��k�����<�a�3-G~`y �h��j�e�N��[�\��ye��x1i�9�Q��g��|-�p��n\5��隹yb�m�#S�������ﱳx�� �c�9�E�i,Ǣs�O��RpeR&h8)��S�4�L��o�cI�����\�M¯DF3*�k__t�w�u�f��kY�.�Z1G�,��Az)������:�T ���1�aۋ�za�]Ȧ��g��ԫ�bh_`�=�%�����gҫnLԻC"�4y��%�I z?���w�)q��u(�+_�Ԓ��hr��3�i�%��=N�g>�R�Z>	(�ɾ������PX� �B�e��CH�Ů��~m��7ET�$a(,��K�ԋ�P���-E�Ye����Ҙ�o�m��qғS��Ĕ��<A��j&4�ޕ�B�2<f���#"U�dM�Fd��i���*J�F~u�JC�%��0�37�;��3�V���W	�zO��#�L�����Af:�t*�M����6��U�[�s�IŸ�WE���9g]�^<�E@ٸ~<���Y
ۧ���8�XO�}��U�}Z��oD	_�����Z�^��E����i�5Ztޒ�Y����l@�0!#(�	�cV�� �Wo��f�](	w�$��uğ,\'���0��r<��=��\��&�3&�v��0�8�+R��eVD<�	�7g*������������ÝA�׵r�UX$�ck�
/�MS��4�Q͍͂!���P��}Cvv�t�veX����K*Ƈ�����o+������F��:9L �^��O�t��l����q䖵K��X�6��:j���lF@�ަ�R^��1lR�!�Ѓu�<�yѠ��3��B�R;:b�X|N&���Ƭ�� 7ūM��T��\@�0J�;t$y�,�Gv�e�'Ȅ��ǝ-�U���O�]0�.�{��h�C!�,,.��pJ�"����KAxt��C�5�����1 �5"?�\�fD�YjM��_�]!>_�Vl���L�h���` �Ck#��_��8��7�H��7p�p90���sC	ϊ����;�~S!��ԇ53��c�-:�����%���S"ks�}sp�vm��(��1��W�u��֗.���v�1�L��\�o�����#���t	ML��Q��Q�m�^F������͑i�#Пw��>�ޭ������<�q.h)��|-�P������f)��0��;�a9
�P�t�ϓ؍�X���F���w�\��I�ΟU]ޣ�K���l�E�����)�m���S�I�~�s�t��G������v.�(�tG�+���>���zW���g.N��	,���\2Y���':8���Mb�V:�ԃ �P���a�{�Xl��=~�P
z0�;[r��]���B�@豚T��q�Bw8�ڛt0�w5����z��=	9�N��ky�G�[17����w�a�i'�@�o>x�B��I����L��?/�~'N��Q�<w�v9�YZ������(�8D �Bc���\7��l�:jTR-��M��J�r_��!v�qimzp �z�#��PM�$��tg���7���_.!�P�8�i����^�5���|���7M���U��	R��Y֒��5�ɑ�m�}� o�\�tQ��0�n��(�Q�B
��0����ң�
�C�%.iI�Z��mO���ɵ��ŀ�UU0����9-E�Fv�i~�;�u�6]��Z�cC+��M-]���)���kC=
j5Z�r����Ѩ��_,�Q�� CnQ��|#xG0�A�!�XP��,��������iz�L��.���CU�ftE������6�()�
)t,F�>�xq-��'�ju�>[��_�g@� }�	�9��kf���;��a��~����u�!�0�ՁWZ�Q�e���u��?W���4�;�.~p�Y+���ZR;dqK0��f���J��N|��v�Q�V�(�3��B��t��R}"?l�C�F��"2�?��d�:̫CJ�k���Ce�R�
΄�k�(B��X�8�F��ЏL1�f؊��X��7�z���zW�?I#�7K,.�T���E:Z�#J/Hq���˱����|��.q ��lxtcd�\���L�J=�T/�uV$�ml���2�]�[���)�?�H=���NF�EE5m�D[8��}b�*8E��D�,s#.�e �e���^X�k���>�Τ�<D���^�w���3߱���JY,
hpظ~P��ô�����E�B���"���+3"�]@��t�M��y���2���.e.U�[�8�2i+�E�LP9�Tg��7w/�e�GE"��/�x�?FW��=\��Y�1ZO��2u��H�}N�@�b�"��93G[b��U,�J,*{�/��$�>�X�L볿��Z^o�і+fc�9e��G0�xۧ���9Z������S�D�S4)�䶉�Y�bpajA��S�/=������C&�
z�5:�ck5��L�������{�<�/��ؽK�E�Z,�}O���[֊-�ȗ��dK�ѯ5:n����n�[/vCbWt��"����k�S`/��F4VP8�]���6��xĮv�\5Q��z���4�����G޽�`u��t�϶1K�TfVɬ7�.�A�Lv�Հ��dR��iצ�;�#�O�|)�g�T?��Mfߋo(�tj�T�}��V�iH�)o[�Xw=��UI�J����
;���*��#s�>�ٹ_>���V���'w,�}R!���4�Xg�r�#�I^Jq� �M��Zg�k��h:q�=ʾ5G��=WҘHu�4XP�̫S�W�2X+\�c�6����H�x.�e{��3�*h[C��,jQb~�1�7{����yb��2��j����pn���8~��ដ�6u.�3��T��F�����J.�N��� >�wS�~��8�S;�O�JC����=Ѐ,�'=!wn�aÑr7�j�K�,�<�}\\���[�8]Z������Vs���وf#~�S��t����T*�lڔ~P�E�]�yb�����qU�P+&�����1.�3Z��e���i[9sF�fm?Ǚ_Q���&j�n��^�R}
�4��nsP��M!\���Q���s�<�("l�2�R��$��a9���z���Y�1��$�����7>��7�뀿h����{����3KΤ&(O�SD�b����A�Хl��<@�řV��d��Ղ����E�F?��j;�h�� ���֦fR��PbtM�c>9ץ
��� L��������Nh_���N���ݍ�l�E�a^֔�-�N�uNk��Ҷ�o��m��rF��(�g?�͗�L��ߊ)j)7t�j��;Q��!�z*d����m�Y�9L�?qȲ���r�Y�Rꈊ��������&��]F��]u���X��F��>A1j/��=I2h�__Obzb���j�[F{R�2w�Ze�2����q�Wp�������8�
/�)����2�Z8�����J�߬k�wBڅ�h���4�K��`wJP ^��g��nٽBN�㩏����&(u��s��U	r1�@�
���%��}�pa�;�.�7��Y���.�m��7��ΈRӭ��_��\0��u8u����o=|�wq��{]4�KZ�ed���[��$_+F�n���\O;]4ܭo��G�7�}7�`6e#��G���Uqdb\��9&�f��G꟢��@�t�o���� =�zG�k8�}�t��-��6l��wsQc��h^�R�ͷ�I����lϮ/�|���X�l�Τ?��a����6���\ZF �(�_���I)���k/i�Q���#� ������"�����:�f�R���0�L�����Pyu�F������x¡�զF
��(V��{�(�oU/=�L��V3φe8��#r�����@�J$2�<�q@�}V��u�?��#���siЮ�l����eX{���R�m�����[/�ȩ!��⸅sU��5�k�S�.|�
G%r��_IsDM7���	$�p��]�~7�~�������ϊ��И�Z�#q|+��6=�PX�7�-e�	*�`����x��@�Q^E����L�^�F��~j��M��� �_r"�7�	�-I�̣0�E�˪��}0�"�r����刿��=q��`�u�R)>�҄D�Ѱ�[Lx��89���BU�AC�z��@} �g�sm<d���S��hf�q���v'�Cb@-�~�iG ~m`��w!�C��d,>�]ʏD@�.�	����o�V`kC� ޥ�:s��Z��%��k�r�IZ�Q����</�x3#�|������Ry7���4������+�SM��^<���ba�Ij� �&��)Y ������_a?]���lsGuw���?-��t��;��׃�`A����o�u,�'��H��
g���~wT���ȯí�sQ�)�έ_`&�I?K{�-W��:F�<'���a�h� +,`���:�D�ͭ��)�B��̹N�Yb<�g�m�s�K1e���U2�,�2q�����;&�3N���Q�l�B�A�=�1h2�G0�~-qr��fZ�2��u-�_�v��Bg2ZTc�U�N��{�� *��^��r6�����N�� o��,��2�]��軨q� �XF�D��ޜ�E��CA��Dp��>�� ~�@[B%�s���8 ��Pu!����^�<g�u-���W�	&z�܁r�p�x�]w`����PαMcp�W��y�ȤO���P�z>x��<t���,ISG�æ\	��>GX�؈�%�͉d_/�rKu�Uc�$j��W	buq �YG��1��!ev�V�����&4��mx�UI�u�[jA�j�A�g�-:��d�SD��3Q�4���穩.5�]_`‘+���������W<c��XH�\裡V�W�֖��v^?�O���s�lk}��=L�/*��Y90@"NB���AR(�>�R�,��j�G\,-�t���Oȏ^"����.���X鹴C�S(��~	Y��WD4�*�i&$��W-e�!}䲯�Y҇�i��v����i�R'!/�M��c����T��d&�RK���2t���
4#!�ሳ0���N��Myܷ���--4��:||ZsT�Ue��ӥe������]04e�,AyX=���:S�*���ǚ�.��n'�l�<�E�>�!ѡ���rR��;P "��=�׏N�it� �bQL���
}��Ze<��^��@^_mȍJ$�?z�¹��d���]:8���~!i<�v�`���Ȣ�0FvI��tֻ=J0��Ź���[u��P�1�ǳ��9k���(9
�����'
>��.�O*΍>e���4��Q�۔���3��I
;D�Z��Bq�ǃ�je��t�K#�s0`��7P�uf�K�P��#�epgD�ytR��6��J�iM���]�\]�l�x�Mm$��EY��aJ�F�k�D��_�7��x�w��"4�gQG�Bs�R�s��UY}
�uj'1f+�R��ùC��&���+�)U]3��am�������b(�c j��)D�:H�@��[L�P�J8�V3N:Gw9ExVf�<~009��˒	!Q)�G����c�[ ��?+�����7,p�,g���,����>�7}�1���-8^��6w{YL�|u2��Ƴ�$�&`v~J�}9�ץiA��V��~p��@�j*ԝݞ�4���u�o4?8���=��cW�OU��тv�͌�`g����S·&�c�"������	�ϱc{���S��и�:|	㿬u�|W��%,N.�y����2N~�WW*@�S-c``�Y1���v*5 &�)���K�����<�����V�*�|wkE&�챆�>~����NS�ۥ�6|yA"�� !����B��kC�r	A/XB���f���?�ٔ> 
�Z4 R��~h}��v�O$!���*�`�B�?�ĘWD��$ ��q��=��m�O>FHP�
b	rU�Us��\��dj],Z��k�G#epD�0A����)b�c�����ں��
b���~�
�ѹ��˜��a�߽�E���.�]���p�-�R)�C�޳f�ߎ�����Z�~aȲYEP�.#pMBAR\���aw��9��'&՗�sȻ�s)0�W�g�F���Tk�*�
�
�r,MrHcI�h�<�H/er���.HdiO�b���"�#a��������OV���2���7�X4q{O�[�F̙�y���S��Ec���w֐�1��,��j����2��r���E�)�D�V��Mޱ:�ɼvk,�,**�M+��>'nF���&<�?�2x�����[Np�����9�Q�F]�dKh�J�k�㍋�o�kE.����6)�4:#_ˬ�6�]�_Z񴊁
���cO�.nA#�:I�\��b	dy�x ����u��z��C2�~�S���l�/UYAӠ�7f0���	i�I!ō9�|Wh؃���j�a�k85Yl8e{����_.UΟ�����I���&�D볃�Pf0��;*`?���8����X��ڋ�a!\��if:��"o�CQ��~�s���9�#|���e�n��-B�_��R{�![Ԩ���L�x���E{'>̛��{�)���h1
'SoI�L���:E��̬k+��\��sG�M���G��%�-mqڌ�'kj#~K	y�  �c�$`�d@�.���s"O�?�8�a�ɢ��C���oS_���C��)ܬ٪%��`H�qa�C`b�L��V�%k
�T\s��ՋN���u/��_�j����Y��]΀m�T���r��^�t�x�'��c�
��f��jD�=�Dstb���'�/_99�lAdH�W��F����F��h������-�ĭ�2�w�D}XTP�#2Ҡ�����oT�֧���X�U+���GBNI0ҕ�4*�X� �_zp�:�[�Y6{ �~;�p�P��>)P��2�� ��0!OҾ�D�u����2]!*!��Z�h��`�v���}�0p��B��@!�HU_)�7��Mx1�Q��t �JJd8lv�I"���a)!3���K)�9�&�7@ٔ$����SӰ����!٪�D~���hxõ:�`m���ԯ?<ND8P���%�eq$#"3&
�f���b�^�S&����@�V�r,ެw�"
���,����U�u��(���֔�R��F.E5�D���JO��9�[Lz42�u#ԝ�T1��YOFZO�2s�*SR!����R�KV��[ŗ+=v�8��=4:�F=�O�w�T��;��������qLR�:�3l�s��f�zZ�)L�p���ћv	W��j
�Al�Z�=���Op�a�����m����)A����A�.�Cn��c0��=������j#(~mlX5e�K�{Ų�M�Fq������Tk�"�^���LԢ���m2{F��u�i�Mj=�R��e2���hJZu�PO�5IX�<�~<�oC�����B#���,���)뮽�[�[�{�4�z�?�쟐B�t��`����ؘ<J+T��:��O��n��� �!WJ�&hP;�f
�n���"[D�8����G"�7��n��ǝ{�U,~iE���XJr��3�^���P�;�C�)�~U��s�4�$B�ex�Q�"`/�[��M� ��p�LTQ)=�g��P�,,��0��@�sz��eIy��^�#��gxy�G9��#�%� �!?] ɒ8ᾤ�Z�;*�Ixǹt��ҽb�9�B?��iW����$+a��X��^^Ve��v��o�W�:0z�Y�v�ۚW
�����³�d	���V@�ٗ^-�UV_?�#�g�f����$6��,af=OaRZ��ӭX����׼�.�M����i���B� ��[*�+�8zmC+v9�@ 5�� ���BN�o*�BQ�DC�-�N˯��0�{�����Ҷ2#�D�)�J �3���o.�4+��vd�<-��z0��J���j�ٍt͸���ldkX���M��K��4�3Z�L�?�t��~}�A2L���!��=B��>Z !�A_���Ԡ��c��y}î����݉x#�>��!k��!��<���y� �A�|^ȍ��'D=!B_���@C��~��5��n��6����2x�b��L�JAT�Yn�B�M��%����M���a���B8,? 6|D	`�b`�Y�ud��a(y��Ge�JRtN �����쵓9cSKc����U��b����ae��v6w��ħ�ޯŁ]�Ǹ[4/�w,��דc��p����}����?5��f�ط����Mo�dV�ۧ����s{�F�F�-0i6ȷ���kU2�%G^�������Gn�����{��3��U����ì�h�� J'r+�L�A��,��'���R�d�k���2U`�)��SU�ť�ISf�Zq��$e$Q2����$o<�DP޵���������3�ZΤ$ ��]1��l���7� T0�,���F���$S��a�Z֑58�(��YW`�Bm���=��l�׼b��`���2��؃u�[��B҅
\�]�­�6Q�t���@�gc).�.]�؄4L�#��ʋ�@bH�;�D>`p�t�\�b�P])4���S��D�W�����ܲ�i�t9ʸG_F�_��a eIw%�ކU��%-e������
%�gO�o �L��^�sF�����;���������|35�̭��i�cp[�ԼD���7�F| ��b�����Ea��[ �GB����t����؂[j��/p>�C���H,�˦Es�f����1��d�J��[�<�~�!ng�͎o�;{���I�C-�%��x2M���P����>i�Aʈ�M��*���7��c�:���)��Rr��#�J��Yg�;�����J������?��,|���b�#�y_�fdr)��T;�U�^��:x\BZ"#����Lv=�-s�_�h��}�}�ʓW�*.��E�|G�E�GJ��
�L��v%��	=h�g� i�*�_J�`�55�_�nN��.�<
w�G��4Ѱ���5�Ο+��fc�uf=i��H%*	�l�0Z�c�p�UK����W TV�O��3�	��Z�.E:�R�����$xi�g������X�kvp�д�1Ac�	i���9���"p���!�vT�U��{2kҰ�7@#�w!��=���8d���.��G��Z߮B. &��,��r�^��?2�%��U֢�X*�{�͠(�,���1�h�1��|G{ �S�EpL����/=����{A�=u Lo�,������@o���J��x�@.�%����h=}�"��wWl���wNl�LĖa��H��{<D�1��لvдKr�JA�|�<"cj@1p��r	w��X� ��Oe����p�8Mt�&a�SD#�M#2#�\��jÃn�{:�2�v,�!U6����g�w>*��=А��u��h!�阙@�}���@��T�a��P؏ ��q�m!�u�ݺ�+��0��wǟ�i�Ҧ�j��U��|e���{T$������KM�R~�J����T]$z�8�݂��(x�OE�!���K5��0�X��9��J�W߅ ��b)�{����,��Kl$�QF_�Px7�����_�ɬ�#�f}H��u��g��Ay|�����O�s�u)�s��&�h�e�����_?u�o�C-n2�� ut�[���A��=ǌ5v��J�14PHpVج!���w�>'^u��RW67F��U�o�wof�[�����(�O��("�_�`%g_AW�ؚ����L^�h;��t��v�Q���{��P�}��)���2Pd�rs�-�>��*,����"��|�`�c�4Z��ҡ>�G�7v�-'�N��a����"N���xD���޳�� F����^`����I��s�Z(z�H�q��� �o�E��J`y��CB@��?-�z�7ٺ�^T�d;��8�����p_���D�D8���4Ρ:>��̝g��Z&^9~��~r�L�68�����&7A[E~���甃4ٜ�.�sh���X�"Z��K�X�����ϧ����(nI�]�P�1+���;He�DA�!�d����ީ���)eK\�G��Aw>�!�m)#�E�6)�W�]��Ft)�����k�μ[��e��5��_�}�� �P��;�Q�;*_���!uH��OxTOU� �M:]_n���l�;S¡z�*_�'�ƞJ���&��-M�`\0�^'�i�<DL����Î����˲U��^�T���@ԍ�0]�U���a�6��K␫Be���k�X�1>ס�ֲ-g���c
j!!C��+o�\��A*D�x憠�=���1����#�s,�3CTT�2 d�'s0/ې��B��%0v�h��h����(�jT�������Z߽:��9-�j7.���z��[Bt�m�ь��̱RU����%��('�M��ի.^�g��x#�\��>6�yN�)*@]�,5��f��K���e�bݿ�Ϻjl�A����s�K�ٙ0�ٺ�q��K�(Xr����|��L%ٶy��ouSąi4,=��x"B�Me�6��An\}B���A��"�Ơ�/�N��U�G���*o@6��%�:���E�����=���!�6��1(*ja��4`Ѥ\���T��`��Jy�B��t0SɦPl��tz?55��}�=I����������vb�ϼ奤9��V�EЪ���z9��}����
<���n�\�;/��o��
�<�'�#@�(��f�j���|2�pu��uԱ	E)}K�����L,�L�H���_g{�*����&����rqֈ�H�<��ը��\w�%1�S��������7@��N�\Ҙ�Q��Ҷf{��=�lkI��&#�8t3^��X�r���H���$��( ��f���_~50���ʡ�`V�V媮�@����I���n��!n$(���?@g�w[*ld��;��cB�O����r�#�m�^ DG(K�\Ah%�ѝ�`C2CZ�]�L4��;���u2��Ft1��a�.%cnu4��Ȝ1	1�K�v|�ɴ{͠�M}��$GI���(Ec �*� O3�I��x���H$�l�E!�����������_#i�.U���2_�T0�iL�0����$��y�����H=R�aC,�OB`口-ڬU��m}H��qW���]!������a'J�r��=�(�Ն<X#e�0��_��G��>�[�
�L���h̗�q�B?��+�Oo�S����U��О7/�LZ<a�v��{LF3���}��ZR�oOi 5X�7e�q��dT��ڰ��E�3�w t�iq��6��@c�5R����/K�z��F� �Fp�Ѧ�ؽT�1�YvWK��m������Q�f?�-��;T�G��Ȝu�e��b����t��ʂ��8�hk,����qA/�j���Eq�Ij��I�^`�#�l�?
J��SV��O����M�ą2���y�p�?SF؇��:NJ�d�b\�r����Ҵ�b�b�@�N/f����FT"����q��Ze��t����0�#c��n�hN���R����>dHC�ڦ'\�]$aa'�G�
�[ġ�0"8�E�Q�<F)Q_�I�.}����F�
���1H���e*������ӬHf4��V���<���w�9��3�<�U�w <�@�:[6�z�*N1G�)+�a:����,��cˬ�k8�D1�N��fح�j�(_��� ��D��Bk�>�%�*�����yH�����'Rv��_�KP~#���Lr^EI�X��P�X���\�о���Pg��WBBT|s�r���]���[��u���~�J�E^��9|�l��^'���VB-��U���+�ɞ�?��0"��wD�b��#���V�r��57ڳg���v9}
&̨5�?�4V2��7���p��x�"=+��>�>�!L����JG3h�M:�bi8�/;lͺ�t�$�- Jv���`�H9;���K�,.�n�p
�Ţ~,A�ԁ�"��D��i	�)�k�3(���ʐ<���E�*1��Vݦ�"2�#4�����c�f!��~�lAXe���c�T��b`��uB"��r4��F�D�{���ӎ�~��������<����} ����]��7�򳯘�+m�t�f��Sh�j�$֜XQ�I�|����3�=�Ł��� �4�DF���H�=~�1�Pxܾ`d����ځ�q�>B!�{
QޭKLD=����Xh���p �RuUR�B
+_i�W��Ak|\_3�Kz���G�H&��"�t,��ֱqA���4�ކЪ�~n�����yV��^l6����y�
+2�'Zcᯗ��3jv=��[�$�Za��+���5�������w��{#2��^��u�pg~����y��x��S߂����vd2f2����l��w�$��nE����6���,�)�Ԁ�!k�ϋ��Vl�G$�����I�|{p�u�g_��<Hy��~��O;��6�)�),^�[!��'tjk�-��9xo%���(�Yn����Td *��n�L�^R����Z/A3� ƽ�Bu�IeŦx��j_�)�ƍN�OD6�,�?=W�U�©d(2N�zֶO
[(�`�;`ø� ���"�󻾶]8,+o������-��'����9?���^�����y�,\��%T��apn��rC'	�_L5�U�)�@��E&,1���S��K�~�*�c���h�?k��q7-(���]�Yb��j�dV�?�v2F�m�\�q'D�xC�N��kT�Ѽ���q'��S8P?ҼᎬpj�82��c�9DHt�Y���i[qD?�U"<�X)0=�ޔ)"�����q�a�B$�P�R�׳��-X!�� Gk��źs�=��)�!��n�B�L�!I�� �ao�_ϕ�"k��O?h��Mɘ�2��!c	� ta������Tp�w�3|���$x+�)bM�͐����DZ�O���ԁ��[,+� ��E�]0v���ZHHB�V�"h�a���a��E�ɐTV���P-�r[Fx�qD��u0�ё���($�=4�dk��<��LŲ�L17<ф\�Һ6��%�Cb]tq��Z/����'�=qg�`��N����)��U7�f^p�Q{3#(��F_���q���#�?�)����7a�|Ϟ��j��׶)$����a�^3��ƙq��E-d(]�w�(���~�c�b򂅩�������$� ������"��z>��.#��SRĀ�c�N���yJˉ8-��1��̘Z���#�29K�ܩ�����t������q𹥏@0;wt�W7����Bd��Ț��u����xWB�Vw,����{���Z���.�?�nVr�����6A�@�r|o��5Aݩ4J}�0�U�e��G<FDՔ�e5������'���p���5�ydC/#^�p4DN�A��#�?OP]�2�1���m�*�wzp��xF�.����;�����+����2����QO���N��g��5������	�49�ó[ψ�I!��%	��p����I~�M�Ȁ��������p/�C�< �jB�LsS��!]�ږ���T2�&�h�/3�֔����N,�����kJg0��i"*��C4*�m��^�#�'�ͽ���(-��b�A�V6�"�/�:1�LY<'�e��ǃ���V3�\�&'�x��0�`�� �?�4g�����AB�򩁌mU�!�!���\�e;!�>��ͨ��T�sӥi��p�}��җ�ܻ����>@���%�A��Z揲P�fS��a�upr���3"��`d�|-t�cp^�"?`��NҒ��cк�R���H�� ��!�Ȝ�՚�C���D��ϵ����e�z��2�����صO� ㆔����g����v~���2
9Bv�y�^K�t�+�M���2M.��& |T�Ꟶ0��a�r%7�
o�� a*>��ƃ�������� �
�Ğ�>9�)i�9���qW�s ��	J3s%D�J��g�H� �ֶ��ϝ�}ۨ4H��=�Yް�e�wG��q=�|�?�Q�qI�tj�¶�U������a� ��
4Y����Z��1ӕK�ie�Ĥ���	�=/�&H��°�RP3!0a3�j������\$0�
iu��M�=s������T��y����l;۩ylgk��{��ӮG�k�&װ��6J�oV���Y�ly��ڭ��o��zj4`)<Sk#�g��|��mc��~��[��](���6��o�@Ʌ�1$.<���^�E���"��J�O�~�[�n:���̤�ig�3���+ɭ�X�
�a��(KH[=���g���VQ����s�|PE����Wd��=6�������v�����o�{c��E�yT�ЂɁ������"�q�FwF��z�3�^��L��K��Jz��چ��l��S+������%����Hc����+��=�X� 鮇�1 -�	�(qI�N4��9&9rC��n��7R��i)�����![�H�?H�,�[jh�}��͘ue�2��������FϞ,����X�y�3�jpB�Kd���F�z��yT��a��t�A$N$-5f���a��[�.+_O�d��+�5h-��/�h�l>k` ����խSE�X��?@[6a���C���(��+�<���p��w9<4�#eXjc��L�Τ	�9c�U�=,4�ߩQ�-Y_��u4l#�6�?�U��Q�Xh�kN5�i��C�H6���oF����~=�L�����IB�DL�Hh�UX��M���B�Ѳf┳�Q��G�釀7�;\2{k��Y��m;�����`��Iidi�[] �jsK ��3��%��K��#&d6<sͮ��Кߟ��F�`���U�{��6�:l�0�>����� �JX�1ڙ>�T��o-�	��@a>����C�}�Db�S��зm�@���������M�x�������"�w�	��g��}�ڞ���xJ��][h�H��lXâ�`����_�9�o̝+���Ы�����$á�� .�7���Đ�f.|�h9R?�x�Ga�^s�Ll��/����Ksw~R��>�>��������5)Y�{4�`�/��j �[���rZ��? ��G�3Z�ɗ�EJ���?��1���ˁ�HYŨ�#{��<eD�FX�_F6���2���6�(ߥFc-����3[,v�j-�ֺ��+�l"�n��.s���c�܏��"-U�Q�����^b�P��"�E`8��4��h$��{�/A�D��`?�}���S�3�G�ڎe3�$��{�������Xv$Bg����Tv�'�e�Ap�u+b�e��,�c8�<\C�t��:��P�#R�,Ŝ�r��}�o��3���'��|���_�?�CPB;Ai�$_��${� x��'KtY�d�������f[�>��sσ�ڀuY��%�A�SI\���r��UH������.Q=�I&���[��=4���4�a�����G,'=��
Z�Rv?�V��}S8�[�#���x�����{@�"AL?��0՟3%`ɇ�'�;$p~��,ğH�ù�4�9���_&�ZDJ��?���*hG�Q(v��p�}pT_2+Fk(0������Iʮg�QFէE�T�.���#(�-�g�AW�ﾂ�	x`�ӈ:�4FQ�0�@��nDX�	���/�e�]3G���!�s�s�'��?t;����*�(Z9�Q٤7�4ܭ�	�0���3�W�yW��bs`�y��"���� ��eYs�gBOn��x7bUO�_��Y�����ghm����Nk�뿡�@�Џ�L���_t�)�Hr�	�]8�lT[�'�cIƠ[|[�˅�4"fG9�ke�M��aݨȊ��93�����P�RRZ���>E�]&�N
[��E~�;�M`l�JOΰ�i�r�}�(��X���UD�L�NZι�\�@(@Q+��(��ݚJ��Ũ��tѬ��o��{N�'�Y##��<�W������O;�7p��~�F��g�Y��Y7TG>���U�	B�?�Y5�C�6�`�NZ����?�f�� �A����]�ݲ���.E�D �����k���="O-#П+]�1K��.>Q�AoUmn�tH�2ri��ш�n}cT��9ڸ%��j3h���w�^��b(����y��C�~�����:�+*�����l���N�D�+>��|f�-Z7�a����Ty�)4|�̆r���RjȐA@�}�W���o
؋�M|�~޸�]�e�Z�O�2R,�����J�~M8!�l.�Ls���uq�ց(���%����F�0�;%�r2f���1{�2�%x�N�O�I����c�2���q����s���^Q�9�{�q��r�:L��oV��4�:�T�	-�)һ�z�Ot�o�T�-�:3�щ�c�g�V������ӕ����.�_u��t���ϯ=�+.9�Q���/S�8��3��
?���O�	ӗL�NN�ՊM��j���b��K�ҜK��dd��	���|ƽ����զ��R��w"{w�7�����2���Ta�P�v�F_oJ3A:�y�\��ue
g�Q6M�u��v�f�93ZUIGi�/��Si�>!��߻��&Ec���֗.�uC�A�P�^Cl��>~���Tz؃ �aBnJRq&�Z�4��a&#�S�{fw	��	AtHY���4��ԏ��N4|~����z7U�a~P���k��2��`?i��Ԕ1��0����u�C�Y|x�${3�r#���602=�ez\F�>5�5M4z�bN�{�=f�뇖�~���
u��4�ˇA*6V��b�q��_	��@��X�?
9N�Lf�?b)�=��L�vӵ���p�h_�lp��Qș\�����-'M��w��	O��3���{�M@��y}m5�����ߩ ���57�?�jPI�H�q�ȫf0?����wq�!�zM3�x;Wf���R���[���
����ozE� E�z�r[on����R�S��2�M%u/Qڕ�(�����Ҝ�[7%'��wMP�+�մ����xC�`Y�¶��^��Hf� �!N9�/�I-�[	(|�~ ���9]�y�5��~��#�jYҔ�/�A;���3�����|�M�_v .�AZd���@h��h�Po��$��4F&Y_��H"����a~8�-C�+C�D6�M�W�R�>`e]禼�U��i�"`�A"qݑ,�$>� �j|Cu4�CF���[�Yl��i�s�V���j�
d>gC�a[����Lg2��|��\�_/G�����#�<\z|{���%��,��q� ����D���1�u�s��l�޾i�{+�V�Y��%�bN.>
���A�	��0���}�2Ҹ�%.�:��NiU{��buEr���5	���I�(�^�.���4�oz�Si�Ɍ��TP'"���ؓ�O��L� ��u֟N�:1���sWVZ����}�u��F{S��3Y`.筽��H��J�c?8��W<�\
T��}dФ�TF	.rb�Ju^)]�1��:���"I|��K��hJ� �A}f�&�ŭ�
rDmjaVB���fP�vX4xB@l�P�A�h� �
�ё"���@�;��+�+_�Қ<��6����:�G�Zh)�hj��E]���2E�	W�c�_7��:�,��k �(����p�Tڔ�l�D9�()�P}gC!SB�� ri=��ׁB�O��ٰ��F5��@��ħ�ʂ{�V���#j�A��V��:=������Bz�3�áv{؞tIU�k6�߻粧,#X���.�RF�^#��2(�y��j.�%r$�!)��5�/bo��Kp�-�i�Ŏmȍ�d�dS�"�<BQLo��av[�z���l4��	\l���O��E��H0� Lݝ��%�v��Pc�o�:ۧ˪����R��7�wTK�0�XKI�����f4�&�{C�ˆ�u��o���Oz��w��EZۮ0WyL_]�{1{�7��r�Ml2t1_h��M�!��5uRwX(h��O�p�� ��HƤA-=h7Wզ>��\���EU�*��i
.�XƘ?�
{���	:��c�J�/^��O��>)�Ç?4��-�ܢ�(m�i�}?���n�Q#�N�T���0����r�h���9=�M���)����9e ��Ԁ<'�j������k��q���.ϡ��䎇�;L�/����Zt��opl����a5��#�$O���C�s��c����o���o�y��T�8/�;ţ���c�尝�p�5)�m;����v#v��ex��w��/�EE@����~�.F;��	2h"?�Pt����*8s������$�;�B�%ޯ&�ki��ށ�+:�Ώ�8}N�f)����0|�wG��>�+F��B�[��Kj�8,�]^L��J�މ�(k��;Y���)�.Pf���픊��Ӯkg�	����c_Zg䜊U2�]_4���9r���)2�\f�s�%����+9��[��;ɴ���sE(�̴u�O6�D�SW�'8�����aܜ[4��������@[���sc������c�u����k���4 ����@�rT����qQ�[�)P�x�Eɪ��[&&�ŏo�t���ċ�\��ö�+�8)^�''f�QL�O�lS�B��ǃtF��5T�){\�g~��6����4�%��v�s%v��z_���2�r�q���D�q�B��͟�C}��a˵��I CP�|Q�p��ِ0�mQ^ij���-�H���n��i)�b}
��D��px���.c�
��TO�xT��{q���<�d$��}����Ewp��g�ϝ���/��z]��+�:�~V#�jS\ �z�M��$���n���wPx�����3���4����[D��8}<K�
&�<Iq�l�R�������O{O�,/�I�&�S�S��;4�7��tdz(l�W��ٕ��d�B�b��Uj�X{a��lg��}%�^F���"q� �@6y��P+I'ϩ��Q=��c,��'�Q*�9��|�zTc�0X��~��T�q�'�0��g�}ʇ;�&;�p�k�'C܎B�,��/����5<�X ��㐺�=�}���R \�NQD٘b7M��}k���͂��Y� ��A�(��*����V}�o!#M˔����D ����p��<��t�cɓJ�W
�o���u{�|%M�U�5�y7�{�M}��bRS��̕��'.�Ų�V��@)�2|���j�c{^�/σ�έGAw����F1���m�s�!p�e5��Z�Vo.F�eF��(���8%%#�^�T�m����V�,h<���z�7؀3}C�ޭ�?�i��r�Ul-�htLwraXYyĖߨ<dms��\����IC�B��A���j����ix:��7ݾ�t��wDY�e�2I��TV4- ��\#�M0!���:{R��6���f�,��񑙬MծE	�����'X������<�Bvo?�k��ej�"K��vC7���*��@O�᥼��rcl�����Yc�ޔȽ������̕�bjZPZ{���3��b�{�{�G�=�0NQ��y3�BD�j�:v�XEA�QZ�ɿtܬ�b-����>��E��V_喐-ܻW�ES6<�T܅l4�W�� �J⛅�`�\�R�U�'�cZ"p�1+���<zitY��D�v�f(N���ꏡ�Ç�������īð�u(�$���ꨭS��:�ϗ������Tr	����p3W@5Y-H�p��@\��1j,z��8�����J_�|��5hCZ������9�l��Mwj	/���O;��i��6D@G0&��;�RPt:m�T%��)�>	 ��']��ӕ������lm����)�7���p;nkJR�Rq���M��Y�N�z�f����Ɛ�)x�`�?-��e?�k<��	­NO<;�Ҙ3y��S���G#b]ţxiHy�Ց����D�F�ХJY��P�G��u����ᒅ�ȶ-C�	V�"�V��U3Hw����$2/�ƢT�T�Ⱦ�%b�4@NΥ�.B�`óߪD�ݣ�$�!�|�ȝW�%�� ����T��}+�C��MXYZ��e|� ��!]у��68P�_p������pQA6
p�0�*����f��6�6S�?������b;
|���k��6|1W�d�ß/��Z=Υ��70��U G!;���H�A�*5l���y}V�U����ɠA,r �2�91�3m����`i%��eT	ðhyr��A�����o���%<�Z�Ҙ�:�a�90���5�QW�Q|07��Cn
�ψjҨ�!_*��ӄ���6A��Ep-d��}(��iNl���SG)���V岈[ ��ys^w�)�-v^��\`�Щٗ����V�B���x��B@�b[�TKZ� ����KHcfO>�{$+Td�0z'u>�R8����q�� N�*{,̊���&��;Ⲹ����ݣ��>�����BϮ�/�^��ř�����?_�NR��p5�˻��3Nb\<�$≤Xb�����-����Z�c�����1����誴҆����?�w�^���ૡ8*I��,��Kw.����7�4��2)�����:L�wɾm����xzko!���ܞ(m��8h*��җ�{��'q���O�=q:*��-��]z{H���H�~�c�F��l��P��;uP��/���}Z�Vq "�YI�#�R�|�,��5n�W��?>۲����2�������+��(�V?G@$Oo��`������*�|i"��s��?�����T)�T�S����A�!����2	��L����p���;���p0��
2U����,���T���~��`Y�V�!,�	8�>g�׷�Q���ܗ��q֍���U��I5�^u�}����Ɖ�����q�>by�'�J���
�js0λ�}���3�p��k��Y�zZqU쏌�MY�@�n6��-���{97���ޕ0%*�1�-U�5a�
`�7Me_�q�=�t���E��bl����q��:�3�i+]��)@�n��+���n��gT}�~o�$|o�>�b�U�,�(�3��i�4bO��H�~3qji��] ���aᦪҨ}�:V�]/&b��K�\�=2��+�R֤�U����"��}�0U)�QDw .�t=Ru�/�F��U��Uq_��"�P,��Y�8,���G�f��:��:��κ-�Ɯ7D���s3��fj#��)l`p�&��ZyL k�x���"�78%h��2��f�U)�����JLE\R�K9M������=-=㠒��px�j����C�g�;�ށ�i�w���չ��*���$
�c�rk�7�pḡ����}��m����:���L��x'��ڱtG}T�e�o�h(R��g���H&�]x�]7}�8���d1_�PJbQ{c-͖% y�i��FŪ.�d�,�;�y�b �S{���Բ�"�K	�.T<G5����Į����-���l�t�
�Z��EL�V!CQ��,?�R�( 2�)
E����V
Vu�~��i��H�����m�æ�j��:4��H�0yI2N��@�ƥ`�Q�
ķx��˟a�[�E�G��������0!����%������ڹ0Txl_:Z�׼˂�ԏ��}Oy���=3���5F���ҕ�N~�0M����f���o+W����a0k�����p��%���#E�" ��V���TLun��tT���K���Q���t�菙�c[� Ho��WF�H�:`5/��d��g���O��a��V^�YD�=�L��@{�ĄXKҥ���<^m�J��@�7*��l9T6P���UY d�l�#ư��W��g�f�� ��J�l�,T����s�VNO��v�~�.׼^�tKcJRQ�gO�{�*���vZ*���ٷ=���f)�����b^:����sّy�%�� ��^�>D�<�����}��aY�Tp�����j� ��H����%�l�m<`.�%�(�p����Y�	����CYL6W�=s� Ϳ�S7Яɤ�BT�vuܖ���Y���B�ْsˬФ���e�P�)Ɇ��3�=K�8���q�Y�]-��/;�4����k�탭�v0�I���cl�T�L�g�rD�4�G�&�[��΅��5��	��6"�d��?�dd��]z=ޭkK"�-��v�-U��9Q�Q�Tg�.���:�n"��7"�H+��i9Fݒ ��Y ��6�]F[F��d�2+�� ؛�q'}�;��޸X�Ɛ��}b�O!5���p��bm���wӠ�gQ�v�k�+F��V&Ƣ��"�t�󶍒dUCU�l7V�:C�� iVs�-����u���t���q/a�jzZ�mq�orYp�*�S�k�{I�+�55����)�É�#avcH���W�	E�K�3�)A��d��J%�a��I�ך8h�4�u�n&;F�@V�
xCjs���
y�d��Y�N�9��N6�c��f�vl~����I,P��&��+�B[
}M�l��%�h�2�n,����n(���94μ����A���	fnSNB�ӯ�L��&���jsf�z���9s��0��+���Wc �jI�m�D������6L�E9pdZ" q�m�}?;����k�ҧ�\"O7Es�@׋yu�	��sH��kI�E�6f�«��pF�5%��Q�ܷ�1�����0��3��a�Ft����K-0+!���]SU<�Ҩ�Un��b9#q��I(�θ���������c�5	����rz����4�ԟ��#�pU[���_���d�UY�?���,c�k���?���5�N�b�'��\��'7e&]�5Ý�kh(��`�-t���q�������D��ͻ�Y��'�uK2��mn��`����,�^��sg����ww<�Kh�+�鶳l[G.z/0U�ΉBD�n`z��/hr����YV��8�\]��hoO0;(vy�0;Y���> >�S��`��L���l��s���Ў@(��B�o�}���"'�kյ�5�m��Ӑ��S�X�?/4G"�8/�3e{�U��c��d��K��C�wx�(Nq�$�r��:e���w)��k�J��]H�&Z�+���G����`'.0a΃O�'��/�iD���"/�X���<{j���Z����%��,�%Vɞe����y���%4,q:T⁕B�� <`,�� ��r!�S�|�����K���$�f���
�0G�VJ23R_Q�3+�����kj�u�`WB��E��R�ݴd��ưEn-NA2���,qIF��Wd�LeW�t�5�P�����v��9,��w�<ӧ�а��'V(s����C�F �*Vx*6�,��bk��o�����9 ƥ�)y,(�~�_#��A�{�KE��%�y4���GWɽ="�<��껖\ӛ��������D�-��zD33uKȃqqB���gq�%�M���5u�K���iy���^�Ｈ�Y�Ͱ�"څ�/>3")�k/9�̣F��$Cx��H@�z�B0j�Q����S��D�0;��,Dy��Խ4���,a#�ʉ���ú��{ĺ�������H��8:�hfU��-�������[���)井_�		f
av���ם'�Z�?M.dz���:jt������Y�����'X���`K�[�A�gkt�V�}�M�gc��R�^���h��o�ݢS?�q��0�n  &c�8=����g�rC懿����"�P��2�f��]j6����)x5����D�V#��s^#d��J���e#�!��Bk�,�������wt��E_��l+�l	/�x/0����Uq�@/ޝ�55(u(����p	2�+�Bi?�C����y|,O�����?�g�8^�#"*2�&�ߵ�O�o�
�7�<��p�.��U�r�]M\���.�����Ď�J�W�/��3��
	�����jw�eB4�C�d>��Of���zb�W�U�x ����~}��19H��Ѷ�1 ��p�_�X	��:�Q7����.�ʆ��2!8ˉQ�nfyga0�����ٔӜF�TH[~�& ��h�-��¤���^9�]�`�k-b��y���?��MȜ(hdZ婏���_),t��HP�G���{>5|)���:Ӓ
�5���E,~s�K��t �U�W����q�T�5S��H�ۼ]�,�C��zώ+]�FpN�Cũ��w��Yמ�r����$�޴��c(Ѹ��|)Ѝr^�@�����e_Lc�,�#��F�rb�����$Ԝ)x�������)w��C�r;]i��r"��G�t҂�����&nDg}�p7L̟�6Z��x�!SI$�ؕ�p0O+^�{X�=Y�֝�ykz��5���0��2Z����4Ű#S��`��s�8d�Z�"��^$�4}m�����_a�y?�N���%a7/��\$��sdEEج��Bh3Գo�����������b@�-΅��ԗג$P�mǞf��l���2+ .�����$ (Iv��@�In���+)F�$�[Ԃ�QJ��?s�b�=�����̓��ڶ����%��k�����M��F��<On����~��r�6*+��s�4�Y8��T�Q�ȼ���U�l�%q`Z��Ё��B^MM4�U����X|��sw��B�T�$����m�����@W�nLԴ�.Ѐ�xfM����.�%C}�h��}�m�{����1?�,�x���i�,�P\c���*����	s���iP�#�R|� A����[�Z>��1�zO���6�n)��I��[NF�z�ơ|�v�C��0��n�j�rt��"��2NV��2���V�z�v�x�U8���[�|����ʊdqL��9�5��7ViS�#V#��h�k����͹.Eo�����7I�g�9��|yy~<<�J6^��U�sn,Yw�!U~�'�]C�w6�
���z��p�3ws����f�y��A^왴��)��BB��`�j+��M�H�򫅅'w�g��k���57�������u\�-݄�/c�1>��\�a�g"���g#"�2b<�_t.~���	���XP�@=z�O�����q��1u�x�oV�&R ���i�a���J?Y���L�\Y�@ Pi�\����m�C4��&&��8V�-Q��Q
8�>�`{tW�ʄ��0�RHo�����"������<�jኄ���*�cK�_��?
�8�Tў&���(��n�kL�4���V�g�q�7�Nɝ#��}�|	L\I�9���wa�	��x�Pl*�M�u�i�9�����ڸ�?$'�W�@ys��ed�u��]���.���:�ށ�	*��b�
n�E�-�:c�q�[c#�c�������y5�{Ɩi@�cKg��ڳfn��j�R{)�%VB4 qLSk��4,_	�b�K�FĚ6��o���>����ڷ��S�q���j����Z��ʋ\��,�;����#���I����`�D���E��Ɂ��F��=��B5����P���2���U���^���u�]Pgˠ� �}M����J�[���n�$�(�!^B�u���۲
>l��q�Rh��iK�9������(yǸ���򱇍M�0�{�^�)`�	.��փ̲1���S �y�!���q8�FwH�b#�iu��ua���!f9�|����o���ؒ��q;~'W��	@A�q&$5x��4Ǐ����'K�Z�#�Xp�Z��M��oڧ��pw�Q� ������fs���o���vs�dͻr`0Ħ�I���i�b��7����	K�n�~dmN~*n(G���U�4����8-W�&
���d"�=$!X{�w�F�2k��֒/���N�FE���B�t5�*(���-��;$��mY��#�������t�b)wί�e"����|�T�%�'�J�Jz����1�R��u"�E�A�}P�_U���4��/�3�*/�;�h�%��3���'�X��OR_�����7Җ�.�v�[>����zQ�IL��
�P��dPapT	�q{bՙt**	�	ݰ#?���$�<���I�#9��]t�����]Fvk޸�7��s>3�>�5�ް^������62RA���c�ߤ�".^�P0�U�g���V)�-�_�˔�|
��<��	[�\�*q���3Ս��@8_��,����{k�xy��M�N�f�*���W�����ҹ�S��+����5O!!G����3�c��-\���m���^Uc,�K�c5������){�`Fk yL��=����e�ao���m��wK�y���%��V���(�[e��zxD@m��B@�#P�g�4~����!��g5�/r������Q�*H�и�DW�d܆�3�-�*��K�1s���2h�.�-@Φ��G���+OS������Ii�ߝj@'���b�UX3!!���z2����&���nA��eD�HR��0�YH���F�M�]��bt� ��5o]q��6�qd�s@��*Țź�����nji�����gd�O=���8�K�8�����C����,��	,B��{4$>l��g�������� X�#jY�T�3��Hۛ*�����C�Z`C�/����>��<J{[� �}�w&'�Q�䯂�5Ghc<+�W�y���R��Н
t�7獦�:Bh�P�e����c� TpH
�����?y�J�LJ�I���(��4V��g��J\4��j�I-�F���M�-;z����l��j�h�sϝκJ���#�9`:,^���Nq�rcH���q�RT�z�ڌ�:�j�'�#i^�h�=f�E�i�
��6���|�cj�;��=���WY������3zs�]C�k����v������Q�Y��� �����0;\n�jkcA9Ъ��8{�
A^��Lv:�����j��mk�b_�^?�n�x�K�=S�H�"L�d5l#��t��� =ݔ6��
�^��;���yxB8A?�Z:<�j����ט>=қ)��2L4�+����˅��])/D�"`�f��o��*1��z�q���f�1g���9Ԥ����|d�2�c��^�	��ܘEN�۲������4�ج�%�-�^]�Tv��K�rm�i#1�q�sл������':�S�k�?k3�J����ECZ��d֧��&�=K|`pd�~�|�l����$=4p�d��h]��Ήz�� b_�O�ZE����	�w�0�	B�Z���L���#�;�.�r��w�m�M�$�JZwD�p\���AZ��5�~��E�_��\�_I�[��j�	���,q�V�)�욲���xd����nY'<�J�w{o�%�oU6oޣ�K��A��m�ǔo�����Hz�豲ǼQ������_���F�&'+N�@�d,C,,~gS�G��q�x_�Op�\�V�V��A�q�����RU9��6c��\-8*_�ڟ�OE��xH�eE��s�kْ�UY�M+�&
��$�m���Ǣ$U�(����j�v`���k|tJ���9<�,����ϐ��-
�bE@̢�3Y�Y�E�e�BUFp�d�� U>��������z�Z���M3���k����\�=�\k�Ɇ*��[��1k|��DEd�zΊ�1�V���*���^�"'kz���p�)�-9S�T�Z��/s&@ۘ����>+(��~^W�X��$����C��Mt��ҁ[���0んV�E�.�/����K$M������C�܄ˋ�V�!yV�J3dR"q�E���r���W�3/ ˽耗p�#٪��h�_��q"���v �����7�i�d�T�j�sʻw���8ӭ��Kp�a�w)'�:۔ ��wʞ�_�������8�)��G���d���a�����Ȫn�c.�pP��jko�VW�;����#~�����:���~p����A
��K�Y�t.��0Eb֚�*��{��f��O ��ӷq��O�+n�M�A&9�\�����4���b�v/\l'�뒂:Rͮ����3�s�ԅ�6	J"��Q��q=4/H��}%��f�7� ov�WҞ�߂�y�4o�������K�Y`F�
 @��z^�=��ϲ"��@	Hy�8p�y8�<��m�ɢ�H.���Rj��Ow��`w����Չz�PHK��������l�	/��g�����׉�K,��m|0z̲�$(sX_���q�e_M��E�R,��l{@U��V��[�+r��J|I
W�tO�'F8 �qM����8��:4H�,@V�/��%t9<�"�u�E�v�k��ԝ�p�yp�㚈���
P ��	S�s�aAaas"_�r1��ݏt"7.��i��:e�@4�Xo��(��#� �u�܋�,����T��b�2� ����m�S��)D�0�[F<@�޵��>J�y�ǝ��h3��)���Sy����p�Yv����,>�'�'�Օ)� ����/gz�'Vx/�؉1�۳�e�>ϴ}��	��2摙�h(K�!�5�Ƕ�
m���寍�N
����G�̷�u#}��Ї|]�7ķ�2��pjfM	eVT��� U�ITXOϳ/�s�$�3!�d���!��/:'%$G���.���x@=g�;PJc��jR��/��E������!W��˸l�	h�*�2�.�ǕHN/����[X3 �!=~>�N�*��QVj�[�B6��4���\��9��CL|©p�U��S$<�0&T{[�֠�c��Q���C|�`TC��ǭ��!�F<�u�B6=�S�,���5�d�*/?n+�UV��-�Q�"�; *��ZO����[$uvx��mTr��
˘���Og�	v݆��	�Ű%i(j���$�s����)}=W���w�z+*�>���szT6ّ�8i��I'�q,��D��� \���HJ����6��Bs�������w��t�juN�Q����6��﷛������6�)�]K��Z�$%�*��޸
"�87���^��r--�Ce;�p�	�~�k�6�s�ik|2�#���N�u�KX��`��l�>N]�;�}ƱZ����U���@R�=ko�2(�͚�(of�8��?�uh^.���p�G��~�KJ�Y��)�A�fB��_�:H��ox�F������h"� ���ƕ���瓼xǤ�.5V��h%":gt��� ���V�󛷽,�+�B�oT��s�x����:>4�����]�	�V:]�XE��A�K!J��c�wfz�L�L��AMM� �[��Sa�k/�l7M�{�0,-�N�t�]K(�eVO�b�)����VG�QI�e�ZM�aSe��6��g�G)�YVog����ќ�ccM��3�{n$�r��;�A�R#�h�c<�[��Vϵ��Tu$����$�'���`���jP�O�D��!�|J:V��V�h����w
�u��>F�~���?�����N��s�}���Y�@��3�H�BxS��t�3f����*S>YS�"�H{)��ecI�i�s "�v`�]�(G�4��hv����,I(&�.Wm葐��le ������ɍF��z�$���f-�l\�KM*.�?��^�k>�x���v���A��hA0�;U�v�ӪUf��s�U�:���;�l�W��=�WG�?��.���������kG��傋��7�����-�ڀ�ȡI���U�Eg���?^�0��$L0�r�[����W����ϴ߿i����83BO`��,�H��c�-�G����_��Ế�}-?p%5��/����v|
72�� �!=Y�1�����o*r}[��?ܸ�ˀn�d���n9��ރ&,���'��ZR;�g"�Ek9p8�%��� >)J�%v��4Z�U�SsW��1��5�,�,R ���ha,�CJ�ц��r>qYn.�G6A!D^~j�)�����d�v�W���@�P�t�6DNyur�X[4H]��$�{��� N�`c�6s��3���zGg���%�S\��v�WS�>O�:�P���'X���2ïű�.ܗU����{MC���:2\���~V���cb0��v�������L�	��shCB��]T�>�|=܀l��Fc��tfĔ6F�P�U7;�w,28�3�1�Q{��~�f=��s��۠�����;n��;9�G���\9��f���B������h�C�����-+>=@�J?M�-���J?��ُ��
1��������D]EBj����ܛ�$_�v�Z��͇�;���?�z�L2��d,��eH��k�V�k��TG�î�:��}n�x�^qy-p��3�|܏��qQ��5�RT�"�M;�П"��+|!n�Q:�t�'�OK_)�=�ۺ3��a�D�r���n:U�p��o��6���'�����@�x&b%��� �ix����Qf�^�e.��g��G��a(�t�^Q�տzf�FB^5��ל��0�s5hę�;ϡ��Lz���ݡ�Bbrn8aQ��1M�ɑv]s�����M�/z>���Qq��IhCt��;���d�Xܘ(���`}�qql�NY$��'�#��������T%��Vʍ�+/��T��#?�ψ\����֊ߔ�"��0�"�!)+>x�g魨B����	�w�ǫN��ti�\ԳL���xԣ��@'@�Y��n{s��fE�O>��]�g�(/��qy*?�^�Ps�)<IU�j��\�}B�m{����OfZ��}3��2���l2�;�C��f?�?g�W�!0� �����A�#U�?^S�N�@F�1�{�ܯ;����{Ɛ���p��xm�M���J����s�pj=� �o?���ys-������g|�Nd�)�4��!V!���g��`�>@*E�θ�%B���7:EkuPO�ԏ��?iC�<=�ː�;Q=���+� ��kk����
�w���Y��eq|q,b.�2o�tcE��b�ݟ	/Bd&���䷄���z��cx<f�@9��kя�����Y��c6�ǁp���P��9)��fna�9����u����1�^珺.�&�W.�i j�"�O�T��R�*�����K���#6aJ��A״��57�hl#>y�Tm�+̱� �ɵI��"�/�8Ju��A�,�J]Ü��-���UKwA����C-���'�JÖ!�;�>g|�n޶O�(��e�.$���|�}gw�Ը�r�v�t�S�KP���*h�,��9g�l�-<�k��p�ۖ�('�X��󟞂*�v���m��#I�s��$[��;�id��\a"-@�KͿ��p7k΍g��,[O�τ{B�l�ǻRO��j1�ϲE9����>�q�@��bFo��

��gW�+O���	V3K�1�9��v�j�1��8�[e��<X!�+P��פ~��`�|�C����\q[P��:��q�1%��>*���ڊ_�
�г:�c�X[̥:�c:D�f�kw� '>�Z�WW����r��`a�Y\�p-e�/�`,g՗j�rWmz���7L���T�r1�.��5��7��>��g�z�	DL�~v����j�2[���9��.-5
(�Lc�U�{�Fp��.�<t���df�c�%Kf��n,���h�v1��_E5j\ 繢7G�ي$85��߾uO1��?q�_b�dY��hN�)���O��]����Gy�L8.ax��0��Èx��N@������Sfe�HZ �KƗl��Σ�{�$�q$��n�+,�K�lx٧8������I�i���${{�����ڇ�o�@bç0ߞ�=�h���ؗ0H��j3��u���1#콟ƙ�lK>��D� �y�������5��s���~���\<��5T�48�e��S�P��$�k}A� ����f�A`g����峀�QJC�E�p�{;�|.�������9-C!�d��L��T�O�K��Vn�����3�M�:��MI�%#�Z_��5�띹����vO��u�#!���S5��A�W�:��4�m�s�Hƒ�DW�O
;
��l��Uz�ZS�-ܚ �RW)긱�e֫�'�&��+�u����6�G��ӟ��^�gK'���F@��{����?�?���z
���6���B.��:��)H���O}���ϡ)G)�C�+`O�<Ȓ"J*ƃo��d][���C
���r�6��}�{���|���a,@N+����O��k��ŐZ�t{��)_R�x�sc��x��53��l,G�Xe]Y
��:����?�&��9��L���θ��a�����3z4�1�/wj˧� ��:*����خ�K�q�̨.��b!��%�B��8ݿ��_�Ĕ��~9x8�x�e +�=�ìD�$e��m����\���[^��;����q����V��k#��ܢZY"�$�-o_�I��Ӣ��W�G? �nG�Hdg��W{��찈i6;{ŹW�&�c�2 {����[��TU!��+ �rDg�������%B�XՓ_��$�-�J��TpXn�%�y�vm��9�>E��g`D����5�}����,�J-��$V�ҫ�u�V/�ه6��D'�������Ӳe(�qc�GƇh��E�+��V�а������3U��jm�+Ǜ��u���n_��pU`أ����qh6!�ƣà�����[}i��O�M=�3)���'��0�k�o�����j�Z�hC�m1�Y3��K���Kw<���Z��M��#؀���G^�i��۩���xTd�Yrg���SRh���m�a�\)��'�1�#`�z<��,t?�x�m��k��6���K�z�=�%b�'@����k31?�>u�Sa&��QVUu�R��f��;�C�I#�-��~k)��{��
� ʉ��Tɠ��� 'RUd� ��:]����"�I��v��۽O���SU/�?V���Fi�SPD�Z�v���ڀ��o��o����'��`�7���{��煲y	�g�,8^ı����P�����bc��}��_���� L����
���1�x�T�Z9����eKjnQ���ur~�]�L���a�b��͠�Ć,��.|$��"n��\Hl���(xx,7�λ��Q����\�P�}�G���l���x�M�3�k�ʺf�B.�� �������N�;k'&�&|��wT޶�s����.n��E	������)*�dM#!�V�3P�t�@�PnH���`{`������q�8��[FAioZk�0�2�Ү�q&��0i:{��T[��%��lţ�/@Y5_,�m�L〗r�Z�r�i<����xav�1�b�R�w&���� Ux�Uj��3.cd��t٧�q��'!��h��Pf<�8�dIr:'\��z�F�I�cQ	R걃S�0vYz<��/c�eX~۩�0\1��)X��g�x�^�n��$�T=�jJ�Ϣ9#'�3���y]��o�i��Z_�YLg�`~�i��Ls`�J���}�m0NjRc���W��ÛV8�K�"��;�R��\2i�f�� -L%��˥s���]�X�姧ٔ
|���!��0o��d��wY���8LQ��a&����'��)>'���EZq����b�/hؐk� [�u�Z.ݗ-F-�� ��~�OJu�#@����aM�&i��(_�l2��K�Ó�V������ l�yk��6���:�Q�a_M��*.iUÎ"ٞ�2�ߋ���r�Jn�~ʙ�o��S�#�ז���V�o{Pl��F	� ���ݮ|�j�/H��ңM�NagԪO}���.��T����-��Bc�v~ɐ��4��� �a� �Rh<w��/�4N��o%�*3cl8����nP:u��_��|le� ~/���7��fY�w󺝂����L�#?�֙Bv��yF�<�7�8d}��H|f��[��q��pe�m4XN�&���=1��L����U�H�8��\շ�5r�b:��Rn�g�]l��# :��>7E�ޜ0����ȇV
�Lإ���眈1o��"@�Q���A��\je���S���3��������G<r�Z��M��Ŵ|�v����׬Ǥ2�2��mWy��|�Z����z�DߴB�dLT�k�����]x�B�`"Z��C�F�yOx��>��*��y���K�Y*���$>J�22��nʀ!����ni�cse�;�"8�l�)���as��-Q���_�j5��l�����nCk���R�5?!<����U1ʿ���!!��Ǥ�^EcU���C��%��>�`�U\�߄�}O�Ć5n��[����*jK#�T&�"_TL-wB&�L������by93��_�������H��9�vL/@����~^\�kA���כ��o-g$�Y��'�+"�z����ޙbi��72�n��0�
�t@C�`;�a+h��T�򚘈�B\�΋�ҍa��3�O�����d���x�+UЫy~[#\!2�R
���Z O�Kߠ�&Xj��h�,��>�蝙�˫�4 0o���ۼ�r�;V����Yܒ�A��R�"��KY�ׂ��)u���o[|+�~en�.�O��AC��e~0�"J����s�Z�mꄉI����DָH�'���󙞹\�U-LSu�*2v�47b�^h�4��`+��۟�>���o$3�/|�:e�I:����Rh
��P�{��>}�~q ��N�Jߊ�O��H��%�؋S&��FՕ��b�pMUҌZ6�\����S���JRۥ�6N��޼R
!��:E�AF�����PD.P&wK�sL96��5ƽ��l���=��q:\B�����dP�`��O���衲U#���[Aj��"[1b���Dv��V�+�|D�C��\C/�r��h�*�.uƨd�{��� �e\H�d�$D�j�P�1&MP��J������w�dV�~I��r*aU�C��4�$e�@��+������ɼL2"j<[T�h<|��#E �>��k�IؚqaT2��}Y)�����{��Z�W�a�?=��/��Q�: ��f�]��ț�ѥmLw��q����Xn����;?��F*{wɫ���K�KM���PH����k`w���a�#�����@.���n�tVv���p�蛐�6U��N�����JD���LRCRm��i���0�g�'�NͿ@-La����9�*��s�:�;�Au�����:4�A��5��+9�)#ɾ:>9|�1�\NRs��EН/b��19�E�0�+đo�g�z�o/{�{��_ϔ�w\���oD�V�����?G�7RZ���5bR��d:�(��"j�?e�� Q�8QL�S����;�軑����JZr��R���̯�G����sAf�`hz��%��.Vq�piŐ�T0ڳ�z�b,�|z\T�Ɵ*�Y�a=�}�ط���H�Mv�����tM��%X��
�d����ω���A�PL�{����| ��:D� �c�Kk6^���I�:e���/8�I�l��W���'�^����2Z{��K��H�K��(���V��tPPg-Ņ�D˼�g��qE�L�FAS������4Q%Åfp��OL̴Ꝡs�I ȶ��q���	��ĜU�k�$�++��G*�=	�&esﴺjR9����V o�g�S ���ѪmU؝�LƏ��Y�%37T�2�'��Ǆ<=[|�]���I�!�v��ho-l��l�t	%	:g�2�9*hz*>jT.�C��ڙpb�����r�v���u�e{c�Z�t�PV%@�� 3����*��ˋ=�L"�.�����M.�/����
LQ��o�г�p4k�����i���	�kq\j�	n�l}.��P���e�9I�uC#�(eڻ�-�&�Ě�*6!�y�F�7Ĕ��	~C@_|��r��M�T�H���3al��D��+�7r�bT�%��tv�Cc65��C����R�#R����J�������k��J�h����{6	W3_u7vk[��O��٤�.U���S�n'!y�"�ԟC$T���y������qn���ew5�3�j�1�Kx�ئ�[,[�x$a�Z�x�O�E�����-��"{c����a�k��@�S=	��j�.�-\}��_�J/�V������B@��T��v�:��x�ix��o��NMUv�'��2/�B�0���-_B�U��z��h��5m��i�e�6/At*�y��@��m�~��/�".�Cn �T.����M�`���R�R0��m��ˉ%�.�tm�'XH��>e��̚T��GV��Q�=������+Y�W�J@��T�����X3�Ocz��4A���m)�{��=5":���b:�w&����`鏡�ԑ~������r��������8��~�!��*�N�̹�����d��z�D�)u����țH��>@�
1bf�`I�Qٽ����W����c�^���JR��jZ�=[�&X�2��pOL���6=��}�e��!VT\��Qp*j�>#��5 'N�����At��YL���pv�H��o�FZ���	1�Q���耇���V�6�_�#��8���s�oiɦ�)k������&�n�NK��1��#����J;Aj�F Ң�;<,/;$\0�]�0)ݩ��H���ohZag�N`I5���NVgM�a	�!�[� ��)dE!���m�&�tlz�7T�S֑ ���_0Ie�h�I�
\��Π�9�/K|r���,�k 1��Z�
��>�G���K�t����I}��#��'4�հ��\�(�ω�tTHaΜ)���	��
Ľ�,e�{�<Ȼ��&��1����g�ןb�B<��+�V).��(*�qՋ��K�莧����b��c���%@�F\UG�׽���E���tQ��
ۭ��Peq9p�ݎj�B�E���g�[aU����A�Ҿڞ��ȉ��(gKR��Eʞ4��:�f��-�7���{�!fq�A��� [��O(�lɱ�M� �F����T�3V#0�1�?7�z��FG���G��T�x�#��-Z��ؓ��yt#B�������������-���m�_Y��?��1}��h�)R1�e�����ߚK9�]H�p�b&������y�[F,�x��Q�^��ynƸ�b�@��*������/�dg�/u^Î�8 ��.�(�-�eAT���y��8�ht�WC-�p���%�e2�	P���uHj-����a&��}fy���?���-�����Lz��JG���2`f�'s�b�ˋu*��ֵ��R&:D��哗�Z�Ѣ���w�Aڊ~��F�'�����6�|�h0�ڔ��|A?=��D[6"W��ߵ��m�S@�����ܟ@�v+��$��	��`�����=Eʘl��Z��G���!�9>u�k�蘾��}���o�偓�?!��^	��QЪ��*<�d&�M=�A���+�a��z�~��2OvzwJK�Y�36���bZ5N�n�|�^qy�4
�� ����٢���z5�fɋ�k�%A�<Q  :���Td������r��}=�v�͸�j�#wu�d����@��`�x���*�	��$������"��Ú�q��ak,/6�V�>f5�G<�-z�=έq]�`U����嶞7��(4��S��3�w�t�7"w&�"�f���2ф��Nݥ5�Y�v����[{U<��<�\������!��:��= 0p�4C�*eW�
^�����?�_�ױ��6��	�;���d�����ڦ,r9���(���BOӼO�uym9���,J5�.;'4V+���"�iO�����Ik����2#r˘�s���'�eO��Dl $$������y�-z��WXje��qj��E ���c�Y�����1S����x^Bj:(�Y��_�����h��I�r0�	�ڴ�D�Tt���ʌ�c=#J~~@:���u�k�Nc
�&~�q(���DB���θ��$�/����Ib�\�`?3�4�M��L �
(�i2 Q:*���G	��g�[�V��{0v��8,/"i��KmM���v�Z��Ü��H���a	`�Qg����Ҕ�T�1M_@�Gy�XD!�݀Q��1A�_�g>�êő�F��ڋ�v|S�>���w�|X�p�/2�(��8Pt�%G�q*�So��5��hx�H��R%%�����]�6F�j��`��XƔ�
'�ƨ��$���H-�����ae,�B�^יqϜRu��lUA%aWcD4a�t�=ֲ�ّS�f:�(x�=?!rn��	�'�	`�ŋG��~�d��TjuI�v��-o/����Hc��,���LzA8�N��T���&�<��Lwo��ս��K�=��ل}�W��Ñ���R(�tk�M1~�ݳ��͂J�Y��'̍����z�+$0�S��{�b� Դ��R�ul���0�����V���7�ND!œ���<��+n �J�k-����	`�\��S`�%�]2�\I�����|�O�sRV��!��r�u��1t�ÇxY��~�m�s�ӽ���?Y�նF{���C��f���.G�<���P� �÷{K�%�ވ�����=�N��Ƿ�PO�Ht��S@�����_&�	�����К�ȟ�k�m5�d:�j�9��7
T5�4��T&�6SB�ψ�&�x�~]R���T�ƃ2%�[����r1�L%�qJ�8��LY�ܻ�֥ ���v�%䀀�ao�F�����ìɚ��tѢ}�	�r�曝��h�.�$�q�i++jj�rTsH$'�!;�)܄d��"�!��@��>f�(z8z1+V<�2O�����a0�%4�(�@�U�nJ*+�)�EAp
B!�EYC�g�'<_qsu��D�]]GW^���A�L��"&D�h% e�_�ʐ\�*�_�Ot��L�f����<��Ѻ$�.l�Lr��,^}����賍,�9�B��:��N��A)Iś��L�Oh'�l����5���@r�#Si���E;p+�C~$olV�=�%����N86�Я'�\�Qv����rbԺ�=��:0��q�ĺ����za��Sw �6V��D-���%�6Ml�+%Y��/����כT�Լ�����o�T���V[��2=c�܌�	��*ӱT9�g�-���� C�lȿ����U4L��������:�!*'�V�Ri�|�G��mk���kI��2V���M���g�F���F�d��/��s�n�{�ؚ�{�-Eud}�t�yE���M�&#�RYZǤU��wAMf~��LH�d/FV�5l�G�}��"OYMe G�M�U��a����3�6���n���!�ͅ��,��K3��#׊[':ڏn��wd�ك�D��[�ga(����:�JO2�=�u�2��(�e��Vzצc�}X�-e�-u1�o�&����1�ƺ�nTNˋy@�s�w��y�i�\<qX�_����9�<}9W\��p�%������R�������>h1��~��z�7[Y���p��=���3/���XӉ�*�mku7fz�����=�eS��N�̦�F�ˌK�Q>g٤m�\����N$��2�niu�LwG�\�҅Ӌ���%��̀B܂��	nY�N�ޓ3P휹��D�13F�a��ZM�]JsSJ]FE4z���l��`=���Y��X%z�C�Өl�S��swjm�M�7 W�Hr?I	7��N+I���j=��������Z��y�o�z?"��a_?����[:���i4onCm��e�o��t
�`4����Ϸ9ϠӀ@Ips�L���:F���g{��qk�~Sצ�N�Ut��+º�����d$��@P����sB1��>�Me���Ήz.�)����.S|R®?��! U�L9L���k{;ِ()�7]�: ˛��U�����\e��=oH)V�Q���g돑�
���nԓ��zM�۩�����w��W�͔V���mۧ˶	p��H7��~��l*�~���N�}M�i��}�˒<�x�_��b�t��-aZ���]D
��A.`�~QTT��Q�$ξ`�7�υ������enQ�.yZ���7o�W3:y4�;�M6U�`-�c�	Y��K���G�4�t��I����c��?)��p)�i����I'kOj�˙�Ų7�3��"�<��1��36V.��Vb�iy�Kv$�������y�Zڶ�z�J]s���T�P�{�	 ���GyH$���_R]����U�Bu�h��� ]�Ud��x̪q:���Et7k-��̐H�{f��J=rsh��)�b
�kD}K�=}��@�o,�_S�ʷ�`z�[Wu���Em����Ak���8����OX���V��Ȑ���O�>x���$PF�h��'�dD��^�r݋8�䫁���E�r�4ꦿ�n;ot
�7�?wu��*9Π9����6f�I���CO#f���&����4cT"�������-Z�l0���ɮcQN^��BB��|Gj@��<����)¯����
,H���X������Y<�����O��3�@ T�����w7���v�R�/��L���*'8ީ�Z�^�yg@� c����`�^8�Y1�����N7��Ba�*��[���7�q|hဈ~��F�j2��.�jC�-����wj�q��ܭ�he�Nm���L�F��n����aT���ͺ2_�Ü�vM�5�Q��g��c�ѠZ[kW��d*�5]��J���R1����bЁ������2��S�N��w�� ���L��;����~�0��r�@f2�f� �\����SNws����'E�a\q	�OԟC�L������;�<�NH钟��e��� sl��IJea>\ҀR�c'VM���a����|�hv���>ܗq�&q��|X���F	?��~x��Fy������u�v<�L#n��Ͱ&`��ѧ�E63V����O̴85-��.��i�h�2	�ԭ�J�ؖLN��|���_�	��h �C����t���D� *�z�Ç�Z����\���F�%��0����ڎ@B`�Lgo�����g��9�пc%D���
��&D��U��=�C�:�rh��5�w�15��O�M�������y{�>�� ����t1XGj�4�w[;ڠp�I�j(�ʕd�E���l�M�b�W�b�8	|��Ё./�X#�ure�P�Q%B�BS��x��zy~33SwShR
��^	�&a^཮�_^�>/��,~;���u��ڢwAK�f�}�
�n�T���@���OR����g(��wT� 9Sk9[�/0 ���
v�
�%D'��߯�M�3A���h ��tq�q�S����ɾf����x�n��wi�����[o,ob��H�0�"��#�������	����~1�)��8�{���$h�&�Z�b?���,�����&����Pq�.<����'_[��V�mk����ɩg�L�>i��T���H�����7���uP��obn�/_	���=�l�����N������&��w6
9;3͘5��/J���<q��w��ʫ��$��k�f�F�Ka��Fsw�Om�9���̇���OH�I�3-�e���z7�6�%���F�*�8�)e`��H�X���] �#B�����J5�f\�e�� ��۴(=���2�nCki��/=\4se.�z�� �g��� ��a4�&i�D�w�q���N��⯂�\�*�u4 [��?d�uD��*QL-<f�����@�#0��U�},� �B>��4�g�JΦC��X��V�"~���q��i�3��-�z��h֘C�J���]=�����%��ڱ<ǘ��6l��>��67a��iP��ؑg1.�룖F?�J�
�$��p�^���͆<��[*η �5:g�µ��;f^�:�����(
�f�Տ��J��X���o��Ig�-��.�jm+�3�,Ȝ��܀P��3���
�T����[į�KY���e���wNY�ch�W�1�u���:d�Dr�P���~��p�,�6��o3��)V��x�  �54ًF�m�$��<nA��gH:	�uR�W�KY�v�h������x%u	e�����SXBW�u�X-�u�E
�K�����S�W��H̶�	�ꧤi�#nӆgGǅ�q#�q*����W��aa��#.�qVx�JO��t�\p�C6>�J�l�^v�-�z�u"�Ǵ��G�x��0�-�8�D��
S芜��.�(���ӟG����ȖPɢ���m�}VPT�����9=I�T�������{�~/�s�v�(�AR�Le��v����_�!��N�☐{�$ֆ�I�<�mh�k��󥵀H���v��IG/M���*%��]Z����n�y�Z++��{�+���8������RZ|J����}Ձ�ā�%ӽ���;�i�8�W�n=�TV���S�"Ȕ��wnʞ��"��	�c¡xP�X�o{��,�+��n���y�z�����(�����g#D��t_�����]w4����j�*��ud<p ����!�6B��aq�y4$��8�&��1�A<����Ӱ_�HJZ��ϭHq�8�X>>#`~F��~F�i,�}r�9-^��˱�~l6����{gSC{���{���·�ۍUt���qz���}0�u{�G׍QM��_ł��k(!M�Y�\����#s���q;E�G˽����\9�A^�̻XF3���G~��B�K`>+�Mh^� ��,�?T�$>6\S�l����5��s ��+oKl�p�, �%����A��M�^k��/��F����As�"s7��P#M�<
w�� ��q�G����aʋ���V�p���I��w��hx
�o�PO�I��/���꯹�ү�iJÏ4��A��m�<Kń���8�z��A�$���L���i�+?� ���Bư4�m0�87$�a��y�f���J�X{9z�1uIW$������4`ă�"����r�"�N�7ǡ�Ѐ�� Y����ݭ�̇:�,Wa�5��`m٠�	eb� #�(�CS�����4)��)�so��:7�hVVQu��Yz�Z~��6YaB�QH��	��~.�j3=�$R$̛�,��c��*�DAz����>fy�)KԊL�����5�B�K@~��$��p���Ξ>���$�9AU4�9�++lU�r�*����s|����p���543�X�;��u��!�z���=�T%e$�zR=e�����*�
���}�I(簍y_��:s�U]��,$z����N��Ī=pܷh��M�C�?�De�t�\0;V��	\D�o+D����tr+h�0"X*�Y� �U҆��u�Pr*���
Pw�`U�{��%��	�����C��^8�ӄ`ػ�ݞs-���}�^y_�ɔ(ߨ����z�������M3��р��+�L.<7���?=ȩ�����&ؑ�V�H���ek�t�@��r�%R�qYϜ�#2D3�_�"k�,\If�c�g�#f_2�vWf�x��M3[w�N/����n����H����ɜ�i��,&�ą4��rV�GP���6��8��PZi�@�
�#�f4����D��Z~T�Z��쥋e��&6?N����5�H��ۜ�ق����8P������6�#^�qʲ������`G�Z��|h�ΡZ�z�I=7��P�93�c2mA��{t��(���36� ���nj��L�r�0 �^<���B��	H�U�7F�� ��T_f$���~jO�С�����!�j��4Eǘ����[�D�{���2�d�R��� Մ�����vX��\�3"�\���bٙ���y����'�%J������T�ˮ< h�&n�Z�O'�;���fA�[�ޠ����o�^�=�i'��:�?�j�h��ސh$Ig�0��	ۺ6P�i8�B���V�k�yp>Bb�6CLM�W���CO�[��;�nz��t2�t�����~S X	��ͣ�S��XA ��}�N��N��N���XRb�7J���C�-�U	���f%B� ��\0��{�-�0�2iI���
�V��Y�,�� ��_i��T��N.����.�4�T�v��Yl�	���{�-:P��+K���Ұ�i��-aX-�Hx;;�	q+f��z5A�Tm�z�f��x�K�t#�-�qo������L8gs�qH��`l<k��	���� �L;&tUh����3�c��P��۹������
���Y�s|P}�pV�D����>#�O�20��>�͸b��j�ɶC5��M:�p@ᯔ�iix�b���	h��[�a�N�R؅�^Ɩ���S���Q��bOTK�S+�HZ,�r�ӽ���ݨig��ԧen��Ql<m�$��V$�,�n,S�ƍ�{����Q�q�\�O��c@��$�O��`V/k��I��2
�E�J&gh:H晍ֱz�L
�j���FՊR,?�?����DZ�cD���t��1�!��	�mx+�:$Dz�E�M�a����Gް-/̶��GO���xֶ�w�mg�ރ!����CK���<nΞ��f���H=�=�S��qXj����� �xK��A*�??$��n���-��/!P	pL��1���V]C#�����>hIw���p*����c�g��f�$�-p�퀖K٠B����U�2-ս��b�Ȟ7�*��w�6���I��R�C�YIfG���\�.XmxE1j�_��߿��������L>Z9��򎱏�D�UB e�V�)g��K�Fx��o�fd�k���]X�ڤ�"�-~�y�����&�V�Ͻ'��G�b�t�(;0(��P�α��mAϝ=<�ȩ	F׹=����E��;�*�A7��-,&f�|�� S���U ��g��깽[h@phQ���V�Wsv	h9&��Q�lj�yMg��ӫV������"�{�N��:	��� o��s��t��xvy�w�#�>LəTB��2����h�sT�0;��C����� �_Kx?NI���#p�n2�M�C'�'3?&1�k���K�)�����XR�><���x�&V��Q�C�y
�[PX��u.�
MX0Q�Bi_�ϱc%�����$+��X=���P�³��^%����]v2�2�b���W��n�n�&�%鴀�>����+uYc|�6U��:�����;h����0�li�o�~V	Q v������fa�����~Z�]����Zh(�-?�zfS�ۢ8��[0�f��;����0��L��:�b�^2��i����'�JϜשK�ܢ��-^����d�[�X�J�J���H��h�jɡ�GwQE�C�ɢ�v��!,1�w����t���I�`쮘�m� oԖ��vx�`�Ɉ\_�OGl�#l��U pd�hEpb%�9wcV�Ž�?s��_�l/	�w?��	4�����H�<0*I,���,��nZ��-5��&U�D1�2ȶM�W�X�|5��M��,�o�9ª\�t�ʵT+�NI��֨ t[G�Ժ��ʶѠ�z����-������Z{�����h�1`"����Wy�G��;0��h|y~
�Y��u}����3gsbk'��M>����.��dtޢ�e��>�����A{I�	�һG���Ӹ]��8�cE�G����.���p��or�s�=�h�¦>�$�5�=�vFa)�l�Y�@}�h^���Sk���e�;=�����|�S�65�s��
�$,W�嫄�Aq����d�����H�O��� �S�>�]#��@(�pל2'�F��C�y�5��~B�&t'�B�	���Y�� ���	��?Sa9Y�N��� �����w�t�X3�EY�����>&0���v�}ɨ�g��8(�yy�1y-#�� tmiF_ݳW&���߅��68y�?)J�%�*����^^�ƛd���ɚ����Н��L�c3�+����l<p�6���U���g�ŝ�4��ߖ~O�`���8+� �^�@F��7z{���z��ks�]�b˗"I pp������w��u�Q����y<Lz ]&�)\�}�����!;�:���N�?��j��Ƥ�k8n��̐��)/�E�T�9��^%�gPuy��tM����ם"�c�I��d��lP3�x�\��� ��`蝸��5��ꅄ�n9�1+��=�
��y�:I(�iM�:jͼ.=�J���O���γ����X��C�o/��+���|΋M���	���a�ҽ= �~C)��PF3�[TqyV�����N�� ������K�#B�<p�4=�y ���.�����!������y3��#D��
Yl�L�̌uI�G ����^��uY5NC��G���]w������_�3����B�o����^4���	:�yGp!J�~�}�︣kK�9+a�/H�[�{7�p�T_��n{3�z��`�hKhClul*�U\yzTj�A�Nl��g��Or�$`<�+��j����9�[#�f�� �{������'t�W�N��3��R�v;��52AaH��o��{��qI�Ә���=��B4���"�SA�j�z6LV!<M����O3���%]��.���O.6�[��K���#_�6����
��Ѐ(:��1_��M���t{�f����ѿ	�/M���w��1�7�s[�N�v����!�N�6��FHŊ]�� ?�{
؄�0�m?.I\��+��u���j��n���ν�w���s\]����Ǧ�WV�����Y�	��Ȍ�A9�mJ�`��Z��7_Z��}�@��c�t��s�4���| c1���3H}/��LX�#�s��
G��9���QG��|�wpRZ���.�K�V��Hs�k�O�g6����bb��Z	�s'fMO��� C��(��Fɸb\�����r瀔,ϑ��������� ����Y��|�bB��et^rU���V^��:P��nW�_C[MF3	_4 I������Z1��f�{�-��������O3�-���ϒ��88����7��@.���0���m��v]Y�㸱n�������p��Y��?�Q/O9��TP�0�sI+��}$��l�s;Q���Q#ɳ�M�*
[|Uq�J��R�s��Z
]�B�?ae�G�?�Q�s��e4|
5'kv	�5+�P�ݽ�+��V��
�>T���T�>����O�9����ͣRr�B��m�Q�$�^MB�BƧvD��{�Nm��r-�Ei�9,}�ƥPV��r��LagM��Y����S�,#��E��Vj�_���+�����\+C���,׃���D�_3�P]�71��-�vk�!��YO�����?��"C's蹪���8����ɂ�&W��M��5��a��ç&�3�Z��>CQɑ�K�O�o#k��R��9�iI7�߈hEG�7����ؕ:�=�}�."k�	��]�U�):,`�P;������b���H�dh�v�~4��SL1b��?�\�>����>����,P2(��Vkȡ,Nx���Dq&W�4"�N�h=?��$�r\��8�Vt?��uF�<���3{�L�8xP:l���԰ѫpm�a9^I����K��E+_�����S�%ψyjp��"'�w�R;>����_��P�GǕ7�qq`��S�i���2�;־xT�Fo^o?GR
9;�����$�=�(�q��p��NKV��=MpU�1>�k��]���D�I{0��"���t��e3���6��2t^�O$}�"�Ee�܅�D	v,�BvY�����/�	�Z�dX�Ϣ��ঊ�=�M9!�O6�:�u�9�3hi��ZN��~��D�o�j�Z�t�%��E��G�2`H¢��@X�i���Y֛�~M4����Բ��@�v�9� ���a+��:�
�����NW[nzᝉ�&��d
Y��� ��Էy}�|��8�m�!|��!t�
߆���$b^+Z�-`4)��0�^�	{[��)|�}�1��?�d��;�׽ֶ�V�����K�J����(Jn�k��j����}�V��>AN������2I탄&~�O��gfX���4ݧ0��HUߏ|�f�*RVT�F�횉�#[o<L�dm�<�Y���J�x��4-�v,{r��[�K��w����S��E��pܘ�C�T��[9�E�"4=����-��qx�,b���l�E���i�84|;8/���Q�*�}�e�-��%$iO/���ݝJ��}Ky���$�%kk���:��v;3?}��]/��Ǟ�$� ZCN}�"4��ř�j�X.�5�J�J�6BSIhT���L8�Jug�c��Ž�h�N[�ᮭ�o��[��a�3x����@�ܞ�pNe�
S���^���Uџp��;J(̚�-�C����*���#XɄP����JTT��;��k5��6��<������*Kj�U��P%�B���k"$]2����}�U{��WH`X�p�Ib ��d7�R��4��(>ӆ����ƹZ "�^柭=��b�IfsG���%��p:C��u���/��T�wh�DB�����J��g�-��{���,ql
	�?������Ȱ��ul�]kt�ݦT�yQ~�p� T�Q{���&�>~_`���s���J婅dW�3i�*vΝ�l��9�Բ���i���n�[sfsh�Z�m�ȯ���g��uC�˹d�9����J�wKmʫq�'[P�\����x��.�KT7U�2��hjP[�hh�g2m�Y)�`��c�j����h�~3��TX=�ӫZ'�ET�Gz����K-������s�	:
t��;~����:��=ֱI�3��_���_��\'�$��	Eu)����O��I��|\C[ G�}P˰q���A7(�דY�E0���+��끫����.�qgF#Yuxi}渦�{ޅ,۹s��zB(�6��[�8�P3c���ݞAW؊��_��z���ڗ�{<&)Y�7"j�m�	1I�z{X��Q�4�`v���`�U��f��]
@DX�K5٫���f�O[6���tQ����N��!5�村&@�znw%��+(�$���!uv���[yn��d,(�qՙ���I;R��D,�`���V����
=��^isq�����6� ���U>�/�J�*�}��:V�T�k��:��\!�a�k�i�J&��T)^x��zr?���9} �F�L�W�<y8��:���+����\�d*~����)->�`���S�:�E-����!���A�uw��M���#R���%_�p��b�����V�	`�Tkkzp=BvÇ;Q�}=	4�&ѓkg��t34te�1�q���W�)��{E3�9�m��n��Th� �V
U7�C�n���%��"�����������ݳ0�L"yY5f�7����W�����  �9U������D=����d�x��-*�rN|�ZdB���Ivӕb5�́�O��Pͭ����ɨ�Ls]Í�Ͷ�Z�Ѡ���5�Ͽ�5K��O9%L܁�:idtY���ޓ��Ә�d����b�IB*�P�.0�ޗ
?&�;�xH���Lp��V�@��vq��?�I>��8A>�6�c��=) m
�]��2��V����/L*
�t��2����j�R�s������FC�3�Ȇv���C4���3E�C���"Z�����%�R��Q�!.j�垌�b��!���uJ�z��]��`�{���z�+���P����q�iV�Q���1�E;��M�MW$Ԃ�</od�G��%�M��X~ϒ�3�*�	�d�y?��?�����Y	��G�wz3U?���$��<��>��D8�*����賀��շ��`����Ժ,Scb�h�Ͻ�WDa�G��F����-��f;a� �#Y
���G��'Ng�1�i��r9�l�Y��p`
�4G!��U��6�y�q���?��6�Л�x���DT��z���Ot,���={ 89@�l���<ٲW� 5�#��,v,���t���8f��EH�~6�^�b�����ToU�0Ǥ���B���'"D7���*���J�?��7�������Bsvqm��D��f~�` �MҊ#��'� ���b7�dY=?L�g�������?9�����1,4d.Q�֌!#���s`#gg�:�^�f�0�m�,�˴P=6P6�;g؄�f�ߖ7O�!В<%h����=q�6��O��1�9��_��3�"�yũ���F��IQO�T��Z�]�%g���\=�
)��l
�RI�qvtՋk�!n�K��l��[ӄs��i��M�����}�.�����5�A4���o�	S���16;m�#*���؄�2�����@�u2����#�����j��L�hk�dY0�B>C����^J.0f�Aeا�L?/IG�~��,eN�%[eL��Y�Y;ש�i?������Њy��o!�s�
����gG�� 4S -��c�b���^�A� P�x�G^❉y!�Z�$���Sw�~�v�N'T���|b�q��I"L�m8�߷��T|��*���0'�l����6�J*�A��rg��v0�t��k8��V�Nn�Ex�X��SPa�	ךP'��q�H�"��;�I��]�v�m����_"v�$#�4kj������<(���.V쬗��0�H�N:���Q�7Hl���F�H��PE���X�q�3�s�"�q2b�=��jP�!��_� �~�X�B~Dm��hG�t���G�+q�pÒ�����/n;{	��9Q��)�w��
�������7&�o�˄�|����t+�aG�N���<t�o���r�:�XY�+Z�S�<!��K\r�H���U)�X��N���O��H���zR��?�ߧ[��9;���\����m'/�w��f%���<���C&�a-U�RD�.�U�*�7�Z���;@z�G�&���m78O��2�^�EE��~j7���t�HR��MTLY��J����(�_Z؇r�Cy�� km�u�����ޘ�E�j1��f�\�,�3�>�#��oW��ك�6��8{!�G��o]������p	���^ߣ�A[c���r��u@s�����輳�|�O"X^	��"���8�D=8���N�8|�1kc�p��V���Ɗ�Rd��ֶ�:�0��v����ۨ7����R*�VZTku�㦗Z[�n��(��f���JF$��XWFc��B�b#3BG!~��[A?���:?C��޽�Xɺ���RN���e�&d?����h��u�aU2M�8e��-S-3%�zrg�L��.O�#���k�ID�jo��Z2MM���Ї�:�O�%��^�9��Mr(3�v3H��{�ڔ�K��'ֿ�#d�>���}j%�b�O#�B_�Y�ͥ5C�j	shA�)������U\�<���s\�O��Ӊ+S�A���
�v>rW��.�*��)*�U���71%��������w��p ΐ�dAs9�g���{fH�g}�GJ���m��g��"�d�������F���uY�k���G�+��r�����%�!�>;y\��Q�T���ԟ0����Km�$en!Ze�E�&`؁� 2l���J��d�������}	�=�X��>$�
����N�C3u|O�o����'ٶܷ1�ed��Q88	�Y�ըqN��	�J���A1�BXR����I���uau��T�W�ź�CkЇ��\��q�+AKƴ��	(�Wb�amCm���Т=L'��m'y�)3�V! 0�m���x@(b��Y�e�Ru-}���O}+j�-��D,U�\~��,�h�����iU��}��z���,	�`�������5t����F���x�Ɂ���!h�K>�aD��$Xh:ϡ��/w_�{�����	�ǵ9���j�$=kFL9uxa�3�w����c�x��T-��so&n[�7&��?�ڤ4G[���?�5���j�q7ɫ��S�l�{ ��D��c
�2�#�y������mgbEk�X�H%簵�ֱV�*�r��`M�+�	��lW)��I��,�1���F�8��Բk�-�~FD�iÕ������>�P_5A�@r��RKŭ�	ؖH��!�>(ӹ�U�0E�tx��f®�x|���,�f>RwZ��|�q!���aGF�,�O�D�})�|KX�����i�s�௿�7��̽�H�x�-$�^ު�A�y>�~����(}��j�ᔠX�|
��\6u���Ƈ�{u�4b��d��`�x��L��UO�\^I���� �Ж�{�Ì���8ڟ�xAMݔ2�K�<t����2#nS��������<'B�F)����p���}n7�nAxU��r�F�C,��;��kj���$c�p�4e�9 ��-@�����.0���u�h���59X<V�r��c5�Or��I`��Z�T5@0�z�[����gB`�T��N���T{D%���By�`�MCN��ɳ���B��0�Nh2ܶ�oh���D�����~=�{�XÃ�Ѹ%M�gt�1����c��I�`�NP5������|G���
 m��'�?�g�^/��Vx+����C�*�@��%�W����~�Xr��wc՞�-2��A��n��VP�}��L��M�`�����If.`;⳺	�U8���&�i����*����H�m!'��;�G�PP�F7zS���-�; u��b�[O�;=󆜄Ήd�^��Û��������.}ǻr���9|.�
!k̥��]����j���L�Ғ^�}/ee����Q�A�Wo1	�	��z��婮���`e��#�����9�YǤ�����������VT�{�h�/��/L��9I������
�MX�궤��!���N.5�H��V6xxR/�	5D/����1J"p�R�0ӳ�թO��(��9[E�9$��u���Nu� K�#5�n����{��w,�0Iܵ�M��$�x���r��K}?�����=�#F����K����[c� �`24��\���3�|>��gFתV���X�3��z���	z :͙�Rd��$D���4��/��X��[#ry�aV��ҁ`Ǹ^1-iٻ&1��7���r�T�D%�PQ����v��|�.#�ɼ��J�ҿj���x���*�}x���A��ۗ�B`X�&!d�L�AG��GX,��F�*���<0�w�3�ڼbPX��)��w�Z��D�|��nN��d�td��R�F=A���͐δ��C�JK��
^���k��o�#}�{vp�����j��y��z��ခ��W�,��r>dLC_2��i�CL��U�w��y��K��xc�#���~���N�>Ɂ�<�k�J7U�Y~AGR��=b�M�R�p���ʯ��.��k�b$d��S�L����a͠�#��l~���|]�����ƥ�G{�AӼQ�>'MWͿ�`[��/�9u�%�����L�p��M���J`q9	>
��佄m���9z���92:<�����c������o߻�;�LK"�7r�tNdS�o��{wh�n����i�hh��a��h��E7�R�z{���~C <�-�|c���K�h���m��Rhq%i���+d�ʦ4��f�61�PB."�@�}S[�h�+�{G�E=�=�1#�R�2!6��(>�A��e����F�y�e��㔩���O��so-����B_���ƏE�A����D�F���!�t���{�B�%0�<
�+]������3i:ޘ�
m�ןƽ�?�"x�5�' ��u���*=vQV���t��6f��~�S+�M�3n�V㻉i,NՌ�C�)}�&!K��x�nQ�h&o�rk`���+�9��������V��l���_�b�ނ�ޖ��,�����8@w1�2��s
�r�؇H�xN�Z�vz�_�i��7X�/xeêB�����9?�)�k�'����L�L�9�L,7q?�E�|��(�W��$@�1�h+�[l6�!�
�v*���'{�pBA�01���<���/��5��s�]��8��8�(�T�[ފ3Y���f��-����$�b�!.Q���z�mغ)4���]���z�o���9;aF�]��i���E$��UT�j�"�@}�W�+ݯ�-��vk�P��@�`�7���h��#�jC��P�t�d��a�#7Ș�):k�Ffޱy��y�^��̱�6P&����6]R� ��0��塥�]p��^n�Y~l\vaz�"��=�����^]����x�F���?i1?^c,����{�!��Fc���T�}as�0��QL��n".�V����N�)H�|��F>���C���\z�t���}5��� �pR�r:X�%?5�&�+4��j�ӚD�a�������	�2�h0�;�;:8��g�������6t/@�fK�x�yM��>��8�K��oW�67��D�	ג��a��Ï���{�5��W��uoA_��y�����n,̾��\��gSQH8k,%�"�(�L�ׂ��SMo��~���'tŲ�{z�7B2�U2Y��u�������><������ʝ�;|*�WS]���)P4���g�޽؆�b��P|�SK��K��F�c�V$p�</�n�G6�����g	��twa��~ț:9P�M%� �18*�"���̇\t�r@].��#X�Fx�p��^%���w�^�[9䧿Yy���G6����1mZ�,�z>X�����l��>i8�P��L�w�9v�JO�e��%/���U�$����B⦬���ULׅ����Z�*��6#?��SaAϛ Z5���t�I#�3!��¦�<�~=�,x�%�����թ�q��:
�fjl�"jl�O�j�lՄ��l	$��)���[����UӾFnedd�����)5{r<�eh�¹H���|�j��ᩫ^P���`~�OU�<�E�,���6�-�82�G�G�Gꘇ���3X��=���bI3��ڱ�=z�G1��?�s�"'S j�}�n���V�*r����x����-��`y�x5)��M���Sޠ���eq+xp�p�y�DsGqRg��O�_^T��樒5�W�$'�9��ޥ;>�������� �X�O2�q\�����}'n�1���������㞿E$y��_Q>�;,�ky�36a�:Q�O~�2ef��ۧ�p\�h@7BjB��Y�%��w 
�@k�����7�|������ʯ��DyV��\g��~�j���4N�%�-{W��rp�#w���e��mh2�[�4r��F�nQ�Wb(�����n;]�����Ϲ,$�͹�NFͨ��47���b-�ޟl���t;:)�>m�%�B��׉�ԃ��ӂ e���>�F��+'<w�O
��ǡ��`�R9�<�H�7��r�0R0�}N���D�j�W/���4��S{Nv�}�>nV[�b���h��|�݅1�x6��yZ k�akßK)"Ts�s6u@�R/H�?/���^,:J�/rs;�u a�?���"nr.��.!2���� �:7���#*��B�2�-t����n*��ń\>�+r=��E^�o�'���jcRA����i,�����n�+5\��^�02���bo�aQ�C�{hvs�
,q�hs�<����a]��������mo�GVW*���q��dy8�����U�5�kң����S��oע�_'��l��� �-�7l�C��`0Խ�:�/D�����Y�]��i�H��b�n)���Z������ٌ�^��R ��܌@�uQK黿�G��Ɉ�����V���˷G� u+�X��b>^���d����Ou+Y�#o� N��%�^��j�!�d���zv@�h}�1�nfFF�6}��;��HU��?SD@9f:쪃�.��fx��6�1��J"��"�?�r��}�+�~j��*#e���پ�ɖ�!H�H��_�w��k4�����,3E�"�V�Qk�����"�F�;�K�P�y#��{�:�1̨AB5�ȡ7���ei6��_Kg/�S�4�K�����;�+M0�2c'�"��-c��ɍ��\�m�h�j���d�h��n�^a�x����G��8#����z�H�s�%vOH\�~^��;����l���o٘�j��ju�`��v���F>bt��C�k嶦��F(��a=�;D���@%0g2�-��z��捸v�k����^��Ƕ���A��K��T�e��c�r�����~Ȫ������&T5���z]��-O%ֲ�����zL��ʹ����{����GrYF��HB9C�ԃ��K�������V�ȓN��>F�ru�N��xȪ��@C0ٮ{���k�l�zU1\�}�J�O��*�7���J�&&��[�V�l���p�%�I�w��gm���0��ih��h:UY��b�sc�V�ɚ�ݒ��yƍ�� ��p�{J��q��V*l��]������&T}V��5 �TvˠI�F�4ӛQ���Yd��5"Vy�H� &@>'*a)??O�!����CyD���s�L-JSG#�Y#����k�����L���%�:(e=Q;��R8��^� R� v� �Qdj�mN���%�E$M��Z#� �[�%��'�^	�6��]���G-^�"0�C���h�VӓYb��U�F}�{�
���~F,!>M��P�� v';���|�2.$4�jea�Bs���;�'g����?��	�Q2�ste�]cHw&}�QM$$�p�؁0i�j�k~J�<���]�\� �Gt��G7p*���5t�����sI>lU�t2�#��+r�d� Nd-h����/F �NQ*?�p4���s#�	�{�)�sbA�ϙ,e�.M6��S�C��ox;�w��j��ړ�7��5��E��`���#B5�A6f�\2��g�)�ƥI]7Y󓛃���	�� 2�� �33���ki��Ɇ��9<B�b4{,yW�%���Q����Z
o<���T�R 5cHBbb� f�{�^h�SL��j圗����d᫁(�z=r�<02n.�X#��"LS)���Û�P�
�ۃ������[m�'�0Ov�9��;o��s;��TWZQCp!5�[+���
D�1��I]�G0��go�4�A�^ԣw��>�?lv���2k�2fJĤ�`�=�n��&��5�SD$��;��M�wfwȑi�L�>ae�"�.�>sd�xT�
�;�]�?��彥DTa6���|���T[<L�=�=]I��ff��/P�~�����^$		v�����C���S�R[�J\cW�]�#�����$�)���F���ŭ�*�>�D[����9ќ���v� ���_�����EZ5	��П�=z�Tt����XG+�2��[�B�[�P��Í�A�Կ� ����qӣJ�sg���q嵗o\|n��A��r��H�w\w���ѻxZ�0�3�e�?��� �j �tt?�(�@��+%�BhnOl�WycT��څ �a�SH$b?�c&��`����;WJ{��|�&�y���\����fM���Y���`�����Y�m2���cg���X�B�ϊ�q_=�a��$�Z� I�+C���V|R� ���EQZ�Q�@P
�="N�FO3�%92��r;�2����/�^d����Ҏ��2��Q��L+���\��^���X�q�5��S������?�-�TJym?�	?+,�` ��L���>)�ʇ����qZA���Z��	D�8���2�q�%�U9J�^�q! E�#�:L����ڕ9R_6ˀ��1n;�Nь�F�|����~�[a�
8����ŪVS�Y��.����y}"^�d�+qp��ol�@�YfYT�g;d��χ��3�(�`�&cx4��	_n����=	�~�I��z����_���D���v�,0��3^/n�i?�Iϐ���ebyl�EP�pݍ�F�-�j�{�Z��a �{�ީ���&�z���.��ۮ�O��A��KJj���-ױ��FO LV�Nj�A���Wu$/|�	%�����H���b�*�l38B�m�M�؇W��v�ʲE��r��)�-��uAX��
Ü@��Iz\c�����iX��I0��-j S��s��U�[��E��шn*8|��+�c���1+��u�E��5�Bw�p`����,��z��� ]��;���=v�n[ԕ�?k��Z��B&����@��fK�5��]��w�
��-;���О��9/`���/)/��ɍ�%��4��t�:WL�W^��P8�9�ڡ���:yw��A'�qrt� F2q�3��Y�M��#���"�҈=��}��=ՠ�mV���-fB2`��`m�Ӷ�l14ߪ\ϿDZeߩ�ӯe�/CT�Ic�ʅ���FQZE�J�-��M��~��M#�;�2-n�^&�9����5>@3z)��skM=��eo�p� �8��"���{]Y��̴��{
Pꉒ�#�Sy��#��l�]Ta��}.D���A�S:I�f1�t_0�9-�ӁW�`Ӎ�n{��YO����{���f��*C��9���@�C����o9-�z���*��A�e�)j&�<��}A�Ȇ�s'O��X4��տ徖?�?C������뇼��	E�x.�VAF|i���3�$G�L�1��I
 ���#.�Lgf}�F���#>�9P�xb�,-T��,�M��9�A�m�SЀYQ]7<K��bk˹����D�c�ŨI���-��z��hc������`l�7U��8ߩ�N��[z7�>P´��i&ھ���hu�h娩D��A��?#;+	"տW�R�s��y�������v[k1�~��~���	�n��+%8��Ո$�1�}����s�`�]�y�"L&�`r�H�ϱH^�v@��Ӛ=@Kw��TF����gZ����5RH�N�+q���Zl������SU���Zb��34���?��#Q7o-b���3D�ܲ��%9��S�+�S�B���6�|��ҁ�ω�]r�s���c�ߓ�̹2�*�Oq!�Iy��&�{�, Lh��Ď �lawY!��E�k}�#.���No�����Zz37v��jE��Һ��}=E�ωQ��hl�ړ;����K`l��LZX=e��r>�"�E먉�ݲ2O�7D����!�n\�����Ɓ�i}ݒ4OI��+���^4���#���.T�,�\�mʡ�i~d�i��/�D9���d.�IL8�L	\e{OݧY�5��� �QM�&g�� ̣���F��rpA%�_�Zdx��6��|��2��8��EX�CTTJVC��!��z[R�3��[;����ٺ�O
�J&0$�c`�Լ���j�U�s)L{�C/�7��H�a%��s��`c�N,=	��P�,�c� ��\ؾ
"	�@TI��yTc�Ǖ��8~�x�KJ�s�"@�O�H���沐3�����Jd��⪍�����І�t@��塕b�КR��74�h���
֭ѳ?���ƞ�%���Q��P�~�кG$EF$
 ɟ8�*3/���
{���ۏ�[׵:�Z�P\���o��$K8��J<6����ϭ���Զ�����m����vwex9�^����X�~�^�	uSr)-��5�������n��ra��v+��*�������`F�nW����|}9��ǧkT"*9)�!
��{X`p��8,V��Z���]�T�%<�E߰d�׺Ps��>�
�3E�E��sp���?�]��<�_rÈDjr�{IN�J�G��*gXg�"A�A><tp*�\<���v~q{�������t��S��?*L���O����T�Tnx:&�+�O��1�~q҂��e��iJ�&�C\ߏJÆ>{�~�L#l��zc~�ΤL��߲�$/t+㋤��<9��6k��m���=hb��P[�\��'ђ�47�l܋��WǷJk2�;\�����"��={s>D�!Յ`�]8!�n��0�%�U�46���Ͳc���C�@�hN0�Ic+O��7��R,�Ң'��C�d.3Ȧ,a���˔�� �S�3��7D-YZ����&�<O�>b�<�(R͜�D�f�n�e��PXs�AȐ((��y�Ž�^��b�inK`��\`�F[}�\Ԭ}'�q�|�y����w1�-5� *;60�o����F�)� )�!�~�$Y~�8_O|M"�b˘~c��ցq^�ѧa���$;8}�pڗ����ny� ��	}�`��� �`^ِ���6�]��,��=���i��`G!`�m}!c�U"~��-n抇a����4^r�o�U~؈\�������D��*O����{ܒ�+l5	.z$$�2�}�
���#�֕�;)�JE�c�%���+��c��;��aA/}�JT�����͸����UW���5�D�/�l4ǪvAG��&F.���.͕gWjS�W���q��[q�qD[��P$X�E"��}7h+zy$���.i�pJ�~���X�%	�O�z�1�8Y s�������'�D�ڹ�!���)�H�J�t"�=��L�8��,��DT�B?	�/A��L
pK��7����+��n�܆�3W(㯷�<�SF+d�a�S�S2�����_��)������@�f�4���P�����g�%	�S��I<~������N��kHЉu� h�q�*�D3�/7}J'h��K��%Vʰ�DH�GP��C�'�z.��;��y���?�S�0����<o�_[D8B����u�TJ~��+�v�ʘ $ӱ�CL����Lĭ��~]o����z�/�l���wGe�|y�YhB6�W��}�� �*Jx4{�}�{��#<OA0u�e2���[k�z2�=�r�ݡ1y�Ȟ�g�d���ǩ�ؑ���]��d��a��'�(�"{#� ����3CQ��0�[�K?<e,�k�G4q�������v���?����wS�y*�����)�p���8����ߨn͟�`��wS�w���щ����l��_	83��� !����,TV��wӟ �yj�:c���S(*Ԉ�D�,���%�M�B3� ��Z��j��A]A��
��8�<Q�� ���L2,U-��20�S��=�s.�N�R�#*�b�J�X����©"���vcw{��חÑK�+�rȼi�������<,q���ό����Ss�Y�L��I��*�g�w�vEgM�H���|(y����*�=�U���� �S����`�r�"a3Y�V��h<l!jj�k,�)�P�ט-�be�5f*������_������@<5j�l��CuV��-q,��x9�".1�)���\��t�D�=��yrP芁iJT8)�H��{HT�N>i# ��0Il�ā�n����lIԡ�C��%v�����R�2d�iQ�9�h1��,s�A18ή�d�ֺH�g�z�s�q��>�o��3(�<�z��귍�̵d֛D��k��l�&h���]}��#���F���ϋ�j>\���N�2����tpL�#�$O�ǯ����(��|#N�C����{C���z*1���W"��Me��@?G�����z
�����I<mk��1L��V�;;{D�h|�[2���vP���3.����h�,��6�z���U���Xqb��&��|m����F'�PN�_��4���i�Hkh:�l �Z *�����k��M�5��	��h�W�-�@:�xЎmO�;%����A�`�)��.�q`=h��FI��
��HU�d���  ��my��d�ڇ�f+������P��7B��(W5+9�^�Ji�"[QF:���_C�dȫ0o
�������VͶO�j$���m%-�u��݃#��ٴ(���:թ�a�`����s_�?��l�q�ɋQ�x�NV��U/�e0���T�`T��˩t���������屢*��뒦GA~jTz�������u��Q�m��^ �6�9vM�A\4��Ju�=ڛ�#�B\"5q��s�z��og�ٔ�B�KJ|>!L�MĪ��;j���'^��7������F���Θ��rfz��n�Xt���8�s�ű�W"ܿ���4��<N%:��aȷq�6�|8����|�=K��\��D�Q�4W���z�<8#�*T�d<�/�Ȗ�@$)��-��@.h�vl�<�t�?cOGf��Z���r�K���g��pd>�(|Ҧ��x�}V(����[1����I�O�I�H�w� CE ��\2�L2���2|�Zװ,^<�*�3~�LȆ��b4�;[0��{�!�8A=��֓V/�'u��a��,�i�ϜQʽg:��vTJ\2j��l��������}���jN�V�#7�EI�9���@�[��)��Oik�l�۳G������xO���(�n��or>z�tcw����ڸ�NP�pd���y��~
���T�żL��Py-1�ujz�:o7�%��+_s�-��Hm0�_��O�XZ�����n�4v��C6n�p�̴#��=}�������k����ݭME��&��u�ntQ���g���mV�a_}��hU}J	K2�����k��2v���{�ލ�А<,b�/�H[{S��J��?��m���'"P}|g�c)�3�X���n��E��7���P�^��0V喇08��¤9,���09߁��f��C� �$
�F�����n*��2�
K��W*�Q'��O`�y�U0��)�M�0h��]P�;���=d�߄t����L�^�Op�J��aL�� ^�-��|?�>�:�K3�Ă�|�IX�����^��g)��m���{U�a�2��Hڣ�0
}�);z���?jt���!�zf�����>F&Oʎ2��жR1����!1*pɥ�#>���p%>�l�����L��B@�ft�OZx�������m'C*(��F)�}���7ԩ�rR�p܎��F�!VF�10J���_D�<�T�Q�K��.pH�2����1�!��%j�����#v�����kNs?奚���4������w�4�5�\P����bp�\��Y��2�7_�]چ�e��@���������X[�����4��*�(x"�G3y-�dSZ�f=+.�}�4gHK?A���cE]r,ɚ#Q���\^�y
)w�W�.T�8d�3�:q")����N���S��!1mC��z���8�m�͸A�*H�w;�3.�{��Z�Ů�P�mJ�[Ҝx����T�T�#[����4<�P�;:X���X�'e/�A͑�O��]�d�=M[:�9N3��z�8L!��P1�q(P�pm�S�����D��ﶧ v"k�F���8�����2 �?��<Ob�j�z%?!��i�v7���dw��K�<_]�����n0ܳ�m����r�K*{^˨w��������q��#p�3��~��p�6~����A����v�R��>F����j�2��(k5I9?���
?�㥼���!u������ QƈA��#������Y7�����ߡ���&b�fӃ9rP����ҍ-��Ƞ-i���;�U�Vp�����<��7�� ��s5�eabB��L�����'>6]h�y��<���m�U\sT��:߽��{-=X� b�ü��ae�[�����-k:�(Z�;P�ݹ�/��_/fG�+j4rDKt��L�r��� K��N���i��^LQ���7z�:�롷R$^J�+F{A�]*���!���_�������9��K���x^�By��&��>a�rL��R�yV�����S�e'����ϢS�>欼����[%������_�zPn�˓�URAa�!��W�\Vh95�?bt���Ï��o������	J��y��}�	ʍ�?�|tBz{�?��f�
�6���dHcDt��J��m���Dv�Ƃ��hj�}u����b�rb�Ժ��H�M�?t�jR��&�cٶ��4q�9��Ύf��iH�E@��i����K��BVe6+�	p�\�u������4Y�]d>�%7�.��^� Ge�W�*U�����(�3���'���1/	����ebV֞��p�^t�o�ߧ8���	g�R]l]�\ɗ�U�2H_��<lHA�gO|d>�-�s~�II�J�{/�VA�vX!+�Z�hE�,��rP	��W��>����6�>-<��/�گ�C����?@KIv�/��˭>�8��x�;���Z����x�g������H��Uk�$�.GU�"K�"�i��=�F��k#`
�h�7%�f����@�x`��� "f	l�~��<芬Dg�g�L�+��X-�U[���^�����Q `�*bڴ�P=L� Ro��@�����V.�ɞG�k��"�����qO�SRX�_s-��ŧ���T��Ɋ�1&N܄�g�^�`dLh�b���.��03�*�l��@�L3�V'3�N1��wD6�Y��41&�wv�EA�8���Qǟ:!�#|�%|���n�E9?�q/��R>�N3�� K�`�JgN�q65�<���T�^uマ�{� ����ZQ���z|e�� ����I�ip,'���:\f��sZeǼЈRjpO�oTw�5S��ěhp@k�V��|�ݴ��G�HuV��8�����O}Щ5�Y���/��'F�^`��+	d�>Ha��YY��M?i�i��!�f"�x�_(>�:� ��T�o�7F��gm么�.����晤AiH�[����~�� Q?H�X�B��
Ȕ��X���N6�Hf�W����Z���B�4��n�ħ!�Pݸ�4��ֿ{���I� �
�%���U�jP4��M�zZ�$�z5���E �E�������>ؽN�A	�ssG?��J�iw^�F)h?�^���K%�^qzKZ:-)%�/��!��W?���]Gܺz���zJ��)	��j�x։�5�2��D����w}FR�T�*�}�WǨ,y|�p��VL�'1�R6_�Q����K�0���2����Vax�8O�#��\z�S?X��,�S|�$�Y�XXH`$��Q��zh�K��ì�}ѕ�2�I�\ӛ��<w���aY�f]���C�D7cO+�-��ɺ�d���v�e�� ���P->�k�p�G�؞�����H��UX���Xy�� T� ��\��a�������b��|=�Uױ��^���Q��_z7�3M��$�/�Blipl���Rq�o����t�㝺�$Y���s���!�����6f����3"�H�@pMmᆛ6���(MJq�E+�D�p�hh;s2��YZi|Z�!�O}P�/O�LTm�J�'(;G�������n2����;)H1rj{����G�=`�J���S�bV�W�f1���U����K>s�etKڪjdT��Jֆα�c�!j�5�QHz^����6-``e�y�O�X���edv֩QE� ��D\n�?9j-�(@�%x$k#��O�eG\�S�͑�E-"��؍nׁ~Z�������� <�F�m�s:�;��+������c\����P�#~i�U�@)Ih[��(�g�IEF��o�is\�{�WUrą��G#��b�xdS�KfXp2#[����g'rR�7���s���Z�A&�z*0`kl�G��X.�7��i��rw_�ڻ?NAz��b���A��� Y^؄U�'Ud���riIY��$G׋���i�Hdu8��(�� �% }���qQ�{�����7���4�쑓�U�VG��k�5�IW�>�-d����6Mz�2М��g�0�e�H�;c�
���d港B�4�ê���G5�$�@׵�`�&0U
�c����`t���%�����~��mӘ�_d5�؍�X���iqӅ�Y�^���c����Tþ��u�l��<ѩ��۝�Q�9��^˒8�8}��=�����@�s`��7gz3��W{�!��� 5l��Z`@��_JF���J��(�nj�qѝ�ά��<O�H�	��|�:��^�����;�����IzVw��>��:{�ȇ���'P�y!M� �_�d'4RwS
xp��(Y�͢G��z7f\�8}�*ҙ�{"�[>���3tMȃ�Mt� C�"6����(���'	#�/M�����rB�[��0��?��{��n�o���SS�
�.[K�Ă4溲���Y暳�Զʬ	&�6�;�!Rŀp���R< ��3��m���,�ό��UIV�@>�,��8��\��ơO�!�
()�Y�&�̴Pw@�A��z����a�	>�	��n��Ip%��n�Ak_P#\#�ȵ��=�pL��`x�h�y%m�f���h�v�=��מ���ʉ,<хR�A��U�=[�omv��c��y0om�fc75J�X�P��p�']`�#��D��P����Y]>�*�����5����p���X�*����p� @��˘��. O,ek�A�I^r -�7�8����n�H�}�2d��4�D����ȭ�Er��|�ڜy��~'��R -b�Β4{�;+K���EחIG�ā}�L*�KID��/t�a`�\0m�s`��՜u������'`ƕS�4K0�k�э�7l_KhB��	��U���s	���a g�r�L�k�hD@�N���E���7�c)m��Kŭgm�;���E<c��MO�X����%z�ǭ���9gb������0���8nX��o�����k�����,��`�䈆��n&>3��5V\�N]��,��C��nL]/�kV?q��"ѽw�)������{��>�@���F�c�x���`�I͙�\���-�Ò�o�
XQD�?��(^��&�zaԸ�������|;�u>�!nNB���'��V�7{|	�6L`��!OJ�՚c�I֥i��R*�N|�d7~�n���\xxkO��`iL�Ӷ�Szg�>���y�/�څLȖ ш1��{��^y���}������6���2Sh��#
&��to�5P��P��Y3$������v��%��@�=�m��/O��dO
=������_C�6"��N���!����D4���@{x*f��˦�G�N�6�ƕ�/tG �]�q�%SQW���������R�[�T��!�P2��~�`7��f��d�V�_zͮEg�#�Q�e�]>�Գf�-@s4Ԭ�����^�
[�c%\�bj����/�F��&�� &쎧������y�t[dXK�@ ���d(��:F�T�?�Mf��'�����L��2Z��]^qāT@�0�����i^-64jHǍ[߉���������H�0������B����?��V8ԗ��X>�ݓ-��s�0��C�qP�P �un$OC�ǣt\��,-U�m�(�.�DD��vb�pz�,�E�ӟ�P��D?VH�	��m�����xXTOXC٦Վ^IFg̨�hʧ��-;5�/����R���@��94�����y*�$���[�/^��o���M��{%�K��0]�����@'�؋̞�9]�W��������!�#+�债�IT�##�3>:˗�®�����������-R(T5�2�e��(�
���]�{�� $e���,�������W*�w�1�v��.vj�lG8p8z���׎;i��S�1�y)��-�8ɵga�y>a�I��h���R-IKW[A�q'���D�	������
�M4�(��_Ql�����g�Nt���{�%sN+I�`el������p����i,{N��bK����z��ELe�O��=��]�����ֺ`�B��C�N[�,�S�����gN��8^>5���Є�}��}a�?��O����p��9�_�ٝ9D B1�,C���� �&ىZ�\���.E6�
�OmO�T�����W���Y1���iEh)7��8��fWh��H_�q��C��t|&��goy�$���c&���Hw\��I¡2#2'�R���COG�	���:j$w7u���`s#�wW�O�<󑐯:j�X)v��0=��!���d� 9}�\��F��Ca�\��6[��J�vw_�1�:%"�M����$Z������%�ɋ����ɯ}0X�sY��ѪO��~ �'��ɩĉ�e@�9^z�M=Q���.�pI={�r&��(�N}!,��?I,��2�����"�x�	LT��,#F#z��K`ב�xf�4fJC_:y�Р��Jqлi�A���es��[\E���3�>�͜w��X]�>��f����a�SA(�ߑV����F�qm�!�������dx#�u�s�K_?�Fw���d�N��'��N����=�6.ӑ��>w�sx&0�)oA�[�miBmT�P�J4R�&i�N������s�x귑���U�_��\�[(oT�#9^���� 
Q���E�q�v+�a_̷=�ޜ 폇�g��,���z��9�⸰���(/U��&�7=W2ZW:X��k�.�W2=�Z	{?�⽹E�9�%����a*|-�~SU��XB/��]�a$뗓�9A���@�}�5��b�>	wE���<KR5X��W�����m�W+�O	�K0��5\z���^��++)E�	��Նt-�B?�Wr�g$
�q��k���1t�Ҹ�#R?�l5B.E�T������E�nЛ`A�gHN� y����dO���k�#�@"��Ns%�s~tY�r�È�<%O��6j(v��Uj�:�`��R��T�WI�K�I�0�}T%�,�~U� �S�?gqQ��e1(�p�����nC]��S�-A�iܘ1�J�ӵ��?g�2P0�ό}���d�Jd
��5���L����u&P2kbn���*p�w���4F����0��2!>Zp���YI�H>��G�����a�j���^�f0�CN����Y��2��k���gp�7?h@�MSr���Qh�,t�LD��z��#�e?��N�>ډ0-�Oo&���A����O�8���D�!.f�e�b �V0'���)��݊T�=_Ub��P�WE���K!��-(x�;i�?�����2Y��WS�
��s��;�� ���Ǝ�댗��z����6Z���������:oPq/m,VG�����3N7�����4FYr��|�ˤ,�����;�.l�n�y��Q#0� �}^���0�QX��O:�#�`V��.0�k���VAhT<ve�sJ������'�%v30),y�+[z���+��z'�� 6Ņ%�8ZKʌ�rf�ؗ�V+��;��O /�$'�t=�9�ߨ��x���٣�i��E��/�>h|��Nв
��4��ZR�&d	��D�VzD���V6F%�0 �hoe ��oRHX��E^�о"�n�������'�2Æ�Ȅ�1�<^�h�s���Jk0�䭆���WS�%�i�H��q`5�,��z��aE����R���X��ӌ��4r�Y@H�.�c!��'z���"W>�9G��!�α�$D(�g�`Jxe��1k�6�c�G��W�Џ�-�1�HR���O�vs���2��~�M �Hi�M��y�Z-"��.�=.�^�<r�C�Q����Eכ�� 8e�u��:Z)S�r�}�X��B�Ѯ
��d�(4@�����W��C��z��e�>���7�d����̴����zM��*�#V�"BE��FK̢?%g�4���{���_NH&��;�ӹ �?�D��ϣ
����$r�-�珴��n�\m�h�A@ӏ������L���kW�V�Kr��fx��b]�@xJ�R>&B��C0Ð��΢�~�\�����{+���2�9�BORl���s`	�	�櫉])�Iֺf�TR�VM � �	*�Ntj���VzeVT��ɖ�5��Dd������G�r����T�/_ĴJ��l f&���|���U�c�e��'�"JYۺ �,k�v�� �ANo_@nwc�O�@�#qGw�-�5l�q�$�����tE�L�������J��%�;�um�����H����!|nXQ��������y��4kd�|�W�e�Ѹ�w�f��.�66l���:��^/?�_I��� n)!�t�~�T�<��{:�wO�_�a�H"�]��송Q���{�AB�U��}Kcם�����B3���(�2��B�D�"��s��hN�d��#�!�V����23q�$�Wxo�Y,%ǭ2����<ٸ�Q���3JXᡑr	o�2�XO0
�z�&��q'��:���#^0D�]U;{Z�T�l=��,�9�p�"�@�:�0�1����( 
���*M�o:YNJn?��O������S�)��K=*Ft~��~�*^姏��̃�ۍ�Z��
�Z�@��q�ϔ}�5��,�ۘj�_l����px��&K�I��df�=��^��ѳ��1t�[����M�˃�	N���jҙI�ZǪ�6�7{Y4yf�ِv+�h�r��841��D�;��$��̘�8NM�B&��`Z$ki�.)P@��jW��j�h��������^3���/T����@g���0����ß#�veݺT��K�k�N|�E}�0(��.��ǌ[�`�5��4{�Cu�f\J�>=�4�&?ilq0���>���e[RϜ.��c�e4��vk->��\��D�q���$	��X.��Oe#��ǋ�|	/3��{W�)p�e[��5lF��d�<��_��Oc)�(���A4w���os�������0е�潖�IX��']�ʉ:�$j(�n��~[��K��_�īΡ1���Ք�znj�-�S�zy�{yO3�G/�C�w"��!Cz��SU���gW'�x|�ƿ=X���|톧?~`=���I#��'y5�.a���[��%�!�d#C����8,�t����]n��#29���M�+$cR��p# ��#R�c�N�}�E�2�a�-絭�|P�h���'���xL|ߗ���]0�b� ��I��a<��ߚ��N��Afa�BΑ!�(2��������]�I�{,�ln�G�L	�4x�48��f�߇��;+u�S^SW����J˭(n9��|7�Zܤ��n�����/��+${�&��ϗ�և��A��Q֞��r��>���ZD<Ѓ��D�}���������$�X�r���S��To�f�ll��5h. �,Ϲ���{�ZV��aO>X���o�{0ۅ%����"���)��:]�����p�Z���L-�:F����~�z���j�Y$B��N���܎q���ɉm�Ni�)�B��v �,r\�wK"&��~�h�k�n����G_6��=_�(�x��ĈFw��? �M��	�����	�L!�6�{9SD�6�T�C���oB�@��U��K��k��[�������4���0I�u�V�u]���:,˒�"�d�\�E���W�{��c	7��V�a�mDM�S8��/^�<���ѓ�:�GHO֨5m4]���+��tO�f�|�J#"yV�F�w�-ˌ�+��^��W�eG��V:'Z��y�����e��N�\�ɆT'&.���c�*�~�ڐ���o۶�Ķ
w�xa:6��,���,��eR���D��5S���O��R�l*x��'�
=����E ���V{��"�������nH��"�v��0�b�Ұb�Iݼ�����D<63��|9�C�ct�=o��ҋД��ΆWFv����F��Sj�Z�RVڶQ��4@ɅU��oUc�z��\�t�0F��DX�Â����a��UW��#t���Yq=��E���q�7QS2(���Ȓwrr��lv�- ߲�Rp��9��<Ԋ�~	��ъ�����(
RR�>��]�;u��w�V�`\�}��: Fw��L��T&�<o�����L��h�١�XA��9A�'5U���y�5f@��]�����m��H��3T%Pɢ�n,ެ*AuJ\��͗q�,(>A���x�� O�%�D��t�\I[*[f��t�$cT�uM��z3���?f\��9I����m�7���O��Y,����@��
Fn���ɶz��y{�G���ބ;*�&��z�����Y�� S2�6��W#�h�(���-��ǝ�Ŧ2-��������=�W�U��$>Y�,������~ڜ�p�!~�^��O."�4#l����tT}��b��oJ����UR�(@X�i�I�H��w{
QS�[�xӸ�*��*�O2I�n�m�S�n�����Ua�*��NW���1x1!�Y�Q�0�YSW�0]=b�`W�s�Z%k�T�����a�#�]��	��(m�c9�p(�	�_0��Y��M"�l�"�t��څ��%.g�"t�0P7�A���dl?�.�Ո���CU�2�݄��F��x^ğM�&rc;"u1�>l_��>4ϫ�k��M�L���+�6M�e��X��f���>y�{;gO��4�$�m�����7��K�����=%~ Q�&�
1�hi�)T�.���}�� ���G��)��y��͎~#�7��o���U�)�,)Õ��O�s�T,�����om�wս�q/^W.>S��OԈS�+��j�-tf��e,j�ʳ,��a�*���A7��q����"M�j�S>)�_�,��< ����-nQ#�Ï�I�w�������8��ub��7v��Ù����BO�i��$7�3�.X5%P-i�:��vX*��ݎy��54Kq�,��=#v�086˫f_9o���>�
�P�$�}�dD��ul�9�8	~s1���[S�B<L3��� 	PB&�	an�"6O9�P���J�y"V���Dzj����Ђ���v	��MM����o3�Y���V(����s�j{�}�=�_k�\n�:�PT�馔�n�͆�\`�^I�R�Ɉ��[�gT3��߆Sk�/��b��x0٘K|��!�����V1J���ۿ4���5 Q������^	*�5��`]�n�φ�p~|X��"�Q�[�T�+a�I�6���<%�tsן�UKYUs�A|Ϊo4A3;OP�*�I�{B�}���Bfs�۷�/������_R6T�Xu���=��7�V����B�-^F�zt
��#V�
���~ip�!}M-�I��+_��b���2�@�U�"�Jz�+�o�
fXKi����	�Hgı�����<Yi�K9 ��8�O	W2Y�o��S�rK�Z�ϧ�mX�����)�H�"�iKǊ����jVU�W�G���m8b]S���R�YT���p�_K[ِ���c�fXٗ�۟}/�̻�W"ڊm��L~��D�P���d���D#oǸ$�K�4�����*7����Uz���_0�%���Mz��	��i��|�S�h �@�|��MA�?pƧ��%`����>Ci��}�}�$]z �:�-�3}����V{��	����l8��� F3�C�-d8g�p���j���ܘ&��(Ԁ�rK����z!�KV"&F����<�t�	Vcȵ�^���� Jju���Ȃ�_�?��x��Y@�l���vd�N5��+�̮u�Iꤖ��Lhȅ��'�q�#zo@���e\	5^�@Ҫ�C�r��4���aȧ�ّa�/^���v*j�IUF[��d��}{�6�/�Fi���M���Z��o��hq���n��Z�{c|%�8�����7�Q����%��eE�x���TQ��`��#�xF��+�_$��~6�6�ӫ����ڃD)y�w�N��h�T.�'/ =u��ZhM⟯ez�d���1j_
쟫�8:ȴh����נsTL��7�&Wv��0r�\���-)<v$)�z��YzNf�S���
.g��VPJΦV��;�;2�Ӡ"�o�!!������':xE���=�9���ɩ�h& Cf]d�:��t`y�	:���4_G8���9��,$����,0d{�}�P�D��(�MBn���+�R��w}�����Mvtq�88zu�7	F5%4���_\䩟�US���i��s��iY�m+��5��I���������)#�hI��M@6���u�Sh3p_J��Ad�$6,�}�����ɵ|g���(�c5��[r����b��c���u��FBm��/	�3w����`Me�d��o�ú�̪��)�Y�&�(���ء�ʛ˩�3`�/�}��=MJ7x�z����˔c�)ɏ������n��I�JS&7C+�?�7��Bq�tl���4��!��[q�nD_Y]L�|b_]x4�͠!��D�d�� ��Xj�[��!u"U�*S���ްF(�#ͭ�W���� ���BA�� ��� � ���I�p)�����<��`&KF�}6^��
�k���S��VhkW��YD�'�G��D�6:�wN$TOu�@:6;.ʊ�!Â�@a��0&�����3�E����T�7=/�ʜ��6�xvy+1�C���b �~a�nѕ� ~����Cb���r3�2�]����*3�b��ɦ_VMZuF�`�>�g6��OqN7N��J6\��x�Ϝ���� �k��j��9:�]!4@m�Hl�q(Y��o��`��n�\�D!КBmQ��K��C�MA�z)2���M��ȍ���J4-���d?�5��2����B,����7�%:%jaK�����6��*��D�zՙ�������!b�2�</�G*�O���i��>I[�Tτ�Dp�0g2|k�����L�τOz�1��=�5wTE����p>�zّ���JrB���!���J�����?��t�3܎Nή��r�ϴp��]�*�G���|�Jv+jZ��e�)I6̜�������W�.@�c������|~����
����\�貋���&�3�����S�xy�3h�	��(l�Ẇ2�*5��p�՘k_�b����_�_�J[������QTj��={����:�:�����o��e�u�45��}i!�7��#� ����?C�](T��`�1����2&���ν],�	��?�K��ka�YVV-�]����f�("��=��;� I������ec n���}l�v>���_8z9�i�[������A8;��k�,��M5ʲ[����A�H(�P�L��eS)�;y&�롰�����c%��5v��wx;jf�f���Y7��B����8��/
�<�]LI�9.ٞ��V��	FA�jjP������1�-�%e�DNa|'�����m��ƫM�'�aM�E�xc��`�K|n��%Nh�8 �k:�BP�<3���U���������c}d��8^�(��ҵ���l���/��+-��Ή^��<�kK�r&}��3�M�]lF _��pW�ҷYR:��QȾ]⛟
UVqi�N�0���,��3 � �N�?E��rØN�p�Y_��^��0����٫*�-�z[���gX(������Y��N��w�đ�s����cH�e�()4��Ӵ^���W�uhȡ��"�!A�u�'�l�i��0�8:����F��n�e��J}W=E���ű�fu�Ԕ@��=���������n�9���B�Pp�^ݡ�6˖�5+��s���� �����MX9�,R���I yg�@;�	o[�	�b����=ʪ9��2�ػ@���O� 8V����\pZ�݂U�l�����b�qD=xN�����g��X��6-�����D-md�@(&����?�z��by�p�mw���z�i̳ �x��u: v�GD:�j%��Y��Gv�¾�?�Ԗx)��wǲ[�Bˠ�)�����f���2`ܘZAD7l|T��ԛ�)B.`B�b=L1�s�oS��%�>ʆh;u.5���������׍�N����G?�֟]�:���dǈ1����� ���Hƿ�t
�vΧ�:��!w���Fh	�m�&c(��.���*����[�M$e����D��h���,5!�
*Bq4�1�B(َ�h�����}M$�sI�l��(s��Wzi�%aM�>2���<zR�P7|X'�"/9���T2=K3y�9������b�ݎ����D�dނkZ>)1�+�^a.�/��C�K�����bx�tU=�t����s�%,<��5G�����=���J��PgT���5|x�F��)a�X�n-�\Gџ�^�H vxH�cc5�]�����9` ��=�i:;�� �����<������O7�/�����z�Aη&�Gn�X�lLÌ�,t��'1���7ޠc�TLϷ��3ڄ�֬-jw�M肁�ꃸ��o��4A/XH�_;��**U#��M?�������&)�u������YiY�����I�Q�x'Ccol����A�$у��?�Io8en|�t��O���7�'��Q�	�J:�� �}((*{�Ls�����q�k�)��{�O�g�v������:A���l#,>h�I������&c!�?n(mp@r�9h`e��6yA]��	�30;�{u�'�܉a���9�^�� ;���=��G��9#���(�!b8/`���nC%"�G�.J�h�~���J_,�7a�="�c+nPź���������"��n]u�����К�ﴘ��MHX�݈���D�'*Kn���Kk��
' d5�>��7�Tb��N@%J����T��R'�}d�e{�0��ŭ�� �Sq�̯��;�Y=��'����j�,��:B��hpf�[�Wb%���	���6|��/��Qa����IT�(���M3<�
�8�뀡��a�P�&����U*.����֤\��J��$y�y��r]���Z?�BX���ơ�V�����:T?��
h�$)5�j@�$2�8�{*�_��d��j���r��w4͇ŏl���u���ߺn=�T�W ���5��U���5�c�?�^���u9�qʠK�7�'��8�F9V�i��}�'�} ���ߥ-�-��b�k�Y���'�I�uB%� `���5�jr�	��^�mO[\��`�2�O�".mK�S��"hk�9`o:)n+E�/k��]3�9�:X�����飉�����Ր�p�KEF�k�a��#J<������,���n����yrМSX������e���y��7�b��:
2�����S�u�z H"�bH��|b��?N�+NqS�i�&�����y7<Ge�dϡ��|���o��CP�^w,��c��ot6�M��nr+�OS�?*�X ��G/�C��	���27�h����]�NR�����h��l���냗��0���wE�L�#�P�k w ����v1��kP��0U#��~b�ւ쉊ڠ�a�^��y4I�E�x�Y�k����ʓ�.�R�	 ��}��<{+4�ͨ+�I�4�7�����gB�?�~P���Y��tn�g�vu_v=L�t����������B���fp�i���^E*��%�;/��@& ���vv���  ��,�m!����a&=YY���&���@�wp`o���6��E�)��c������-�'{I�T�$���#Β�s_������~`�WZ��8QY�!|4�]4Yϲ"Ll���U��!��Qvs2ʿ>e�f5	�����Q&Kx�K)4�M�َ���EW�������r2��9��������*��M��T�{c9, w�j�T7��u�N������(Nv7}RWV5��wai���j[Sh�g�
�0|�܋#�ߧ�������@�羘�w�b�.,_�%����������,̴�۹_�Z�~,��ۗ���H0�Cg��S�jJ��=� h[8n�Ġ����Gb�s��F��i�ڛy��aY*���k�I#5�`}��Bcj��7�9�u:S�P�aۇfn3�� �}��Z�H�Ⴠ!מ�8����4�v���o�~��:�c;��O�O� Ihe��)&+il+����X70R���	��FZfԇ� ����Q	�ń����I2��:��� �֓}��F����Y�?d�w�h�_�e��� ;�wPBǼ:0峐�U��o֗��/~�ݕ�����n- &�Q����m�]IoƦ�o��U9n��_YX/x�Wo���~*guk׍#�b�+�ú�\h���n��1yA慈�U�L���;	��
t�DS�O��N���(y?�*�B8��Beo-�ź})o��ϧI�M������m"�U�����*,;�c�
G�܏���!�10cXT��6��|M��Q.T���'ꘄ��8���s���jV,"B�B�r��Ri�Ìz����zN�m��_7�Xk��˩�
����We�#ᖢ���#�,{��\�)7�1��$����{ڴ�4��/Uё=9l0?h.ι&�����^~
�P�y��@�+��<�tNLau�������MrI�|���6v����5ܿ}�q�W��ޥ�J�3���
�9Sh〗�S�A���^ɔ���)�.��,MDJcb�q�����<G�wID�Eg{��,���_�_%��*s���ׁ�{M�����L����Y�H��h�SټC��ı������F�Fi�N��]�>8�2g&<Ug�� ^8� tܣ<�=�S�ђ�S�B�J|��:3�vctA^� o��"%	���۠+�\;�B��Ō��C`�S��q*�R'%���qG0�pY?ҩ�͆�tI�� �b2̹�h�Dl�l���e�rip��\�Ҁs
)�K[��İ�1]C;���O��o�V&�h�����i�i%aQՒ��WQ`K��!k�?��W����H(v�׵��]ڹ,;!��S+q,�Z��yk�f��Li�*���Q�+�bq�Z�^��-?���B�#�p:@b��*�0����π'�\W�\
8� �d� 1����0�h�?�4	�����뉪�8�'(E�"��p��z0�o�:�4_`>���_�?�Ѵ�[��'	��HoEC����'EdݼY�p�t��n(F���@�yq��3C.�l֗��Ɩסo���!8��D?E�R0Q}�Z���A�
��ƠBǋzD���ucT�f��t*��8i\Ko�"�1��߁��� ��P) �v��/>g���m��ґ{g�ч:�(j?6`ȴ{���;�����_��b�U�����[�I&[��;z�ΤS�Yt֙���l�ͤ�5irfXq�J4^?)��Y;پ ٝ�)�S�|[���3���Y�;<_���(t˰/bǨ�Gk[���6��'5�^��?�07ӯ�u���������e�to�X?�#@����V�\X�	4E���*�F����b��
<�����Zj��d
 �d����e�Ǧo�`�gfi
�}���h�	}rdz��bU�Pb6!!7�,A�St`z�<Wk�a���aj_�0�|/�g�MA�_;D�1P�c���^��Bd����J�0��������@ͫ�R�E�Jlkd����+����~|��'7��YX� C+\x)!�<# �{�濯�������C�@��ܴ�á�Op��5&N��i!�ݔ>���V��`�Ƃ��"�˽��^�GvV�����7Q�,���@;�}�**"�a�
&rr[�(�1E�s0iGH�����[��6��WO|I5�$�#�jww>�D�)�6�1Sn��10+/�^V�3��`Ͷ���h~/���&ٲg�
��d}w�=��cqG�� ��hy!V��_��C�i��+��*�I�P67��21�:� ������9����Ç���u�f����3�Tش�C�^IX�f���&ՠo�nk�&����H��S�M�LQ���;�TP��>8߸~�=�#)�n2xΖy�N� pe6Sw��Ot�����YK68t4E7w7��~�&~��Q�W��o$�@HcL���O�C����A��2diH�o�PL�@��W2�k������a���G@	�i7I>hÇ�l���R@-�/l�^���f-u�O��/Ҫk�b�3B���G�4��xf� ����	>���G,�>A���D�X�;����B+��R��?�o�|�?r��R�aG���cǖ1c\@��9ۤ2G�8��Ƴ. ��64�����{�l��|U�2x����q}��,,f���'/ ;[���Ғn1p/sB��-�jy2TE�<?&�'�s��yb�&����L���i՟��U����W�4����K� ��/}���0���Ӫ�M ���G��h���c�y%�_��Vβ��3Ƕ�X؃�U���i�[��P�@�[5lK#'��6c/m�2�!����2}D!���X�1������O�?��R�pC��t�T���y�睊��ۜdi5<?�����E�!i�[1���l��Q�įXAwBRiH���(dK�'Wk��4ޘ��1YC_œ	��ǣC( ͮ7���]��+�d��kyu�� �ջ�z�QH���E땎P2���Zo��7'��-�~��uśv�\+k�m���(w7�ot8 ?���y��r*b�!8X���͟M�I���k��Y�9(!3a��R���딋�u�'>���sGa ?����������Azc�>ÉZ&���Rr��Ϛ�Q[����@��
p��xl�W��Ö�;�5/��`�qPR�^B1?5\��@W����.m�J���nB��f���50�U�ҥ��8}��HB�r���?�*MoO�f,�I����U}׌ĥi����d�3�̈{���J�M�BE�-�@6�I_��C<��k��PBAϻ�ی�����Y�2�
W�J�XqX����֨��h0��>F-��-K�����4��.ܓ�g}x�`
.��zz��a��:�wwbBZ?�b��͋�Sl����)�C�GF'����U�/�t��39�	T�4D��3���ޤ�uŏ�� �2�O ����L����',z��92�U��Ѥ$�fE":d�s��\?USxv�x(&*����@��	�[ص�+����">]��ƃ3�F����eU1-��|��6����{�����\萉3mFy���t�-#���UU������(��J���95q��"�#F��U���ڸ��KSo��XvZ�L��2%��(�R�<A�s]�)G�VSh���K��7����������L�Qk�j1-�c�w��U�c��ag�D"�F�M�k�'�!��	/��!҇��9h��Ͳ���qF�$��|7��M`�V�Q�w�m��9� 62����7l���ˬ���C?=��]K��wFEt�,����m�ay��vbUK9jq��q���˾��68pd�N�
 +ˠ��D�@��)�����M7����M4f���[����E��ҀF�lJ�#���Tt�;�!�x��kk���1�V��Ql�(dl'r�+x��
��߼�~s��Z�.C�]�E��%�1F�W��c�HP��#tp�c�^������ox��l������m��P��j����5A��!�vP�����gR܎��q��@$�k%mX$Sfe�s�P�^43F�>Vl)	�߲��NӶf*Ɛ��X�Q;��V���kbu;�[<C
����2��	Ձ&����1w��������������-�,�����J��J��ܨ	���ù�32a~�i|Qlܷ��
-#�W�\��3�j�_�m�8�F.h�ĳW�~;Q�z���%,��/D�������QT0�b ��)�(8f���%����%�)��e�l^���	�o�皘��-+���U�I>���H淂$gSĒN��k���ȿ��&r��m�U�a�g�*J�i�}ɩ �wQ���F��ҖYD�����տ�7��pZ;<j����T�s�Ǚ�ÿ�y�3R����OY�kb!l�h7����k�D�w��&))�8�> ��C<��U�	�F`ʺ5�S��������DH��u��|=�W�:.a ���gX%��\	�kBi4-/�ۙQ� ��@[�X-q<.a�Rgޤ�]�/�����Cx|Q);��Q��i�JG���N>�O,��rJ�]a������}o>.��=\�F���f���ω���8�%D *��J��-�E�"[d�OT��&P��� ���0
$��َ6P��_��؜6�`��	�d���Bw��)��Ϭ}�w����{���`u����ӿ�\[Cp���d�ZV<��$��� ��%˓L.`�W�Jb_voMG��G0ri�˩�v{�`�g���F
�*
\S��\�g���B�ª#����xq5c��=�-�wK�I�4�T��3� ���N�����x�k�����u��7�����pL{}�TPj�p���bb\U^�a.$O�/4g2t��8)c�c�$Uz��\�߽���$P�Q�{���#�?���k��n��q8�!1�)�̠��w�|���C.�i�7$��O>6�o�I���?4�k���nj�{{�Q��ĒS�L�W�NNz{���6����@�3�Z��$B�u�o�|w2�5.a��sp�_��W�{�cI��΢L�b2�T� (X>���L�v�#���%vưY�HG�i5#������~cl����~J��d�r���Z�Y*���]_dn@G+u�Q����h��By��B��.�E9���� ��5��@C/M��C��x���`ңv��5��<�4.�a��a/}�6�����	��G&xMi�]��͛?ܾ6(�q݄� +ƫq��;�l�/]�qBH�o8����Wd�_p��f[� b��y�z�6&:!�_׶3�0Ǣ����V��:��Ǫ��Fpd �-�ʥ���a�w�~��?%Qu�k���s�_��RI
��=L��4���	��֐��I(6��k:`Ve=D*es���R���_j-u}���$��a5�0;��S��9,�(�� di�S~ !���/V��Z;��Յ�7�ǓN��~
�)l3nc��Tz҅��g�Q�^L����P=���lH��S�ם��v�U�A�D�O� �f��#V�sAt�U@���lg��J&@����G.����@=�R<�x��-V,���q��K��A��훢Y�`4�v��:�.��ln��(�r1Q���J=�6�`/�Cf���g�5W#/J��"$�1��M0Nb�&0������Lr���i�/�尐Ty�U����o:��wZqPc�ιs�t��� >}�K������b���J������E�Ux����׾��Tq�����f�#��))c��C����4#�a���v@w����k�]`���	m��F�{�K�5n-
+2��7>��gj�fs5�'�$���&SĂ��|��P<n��G{���6���;$�U˨����	v�����/ ��vN��y��K:ˠK�D�{	1b5��0E���f���@S� ,������H����x#����F�~�r(�=Z����38[�g9Y���h�����Û����q7���"��݌_�JP2֠��:��r�t�-�i+��Qx�,��Y�ZN�# {9C*B6�*�z����#� cF�#����e��'0��Y��������z7l��һ��֜����*���ˈp�&f���&F���Gn(R���r�As��#O+��J��`���B�B0<"����¦v�%��J��c@A�e�vm���g�ji4������F�Q���*�����MȤ���,��H�3U��h������ƅ��R@lP4���@��ec$���@��e����[�~��'*��y
8��
� ����Jq����!��7���WF�1tiJTѝ�e�]��Wr`�G!ݸ0
y���m׀[���b���^������s�626�?�y| � ��2��4W����#����5����f��$���~�.�`�o�C��΀��i���H������C�ZC�!��C�:��掞h�iʮ��vϒ�b5��DDͺѫ�,m�v�&�4����eU��F�̍��4���J��0��,�3�E�
�aT�& G<7]�D�⊺~�淉ZA+�+b����K+`� �; RN?�1���M�Po+{	��Q��x�Vz%��-�"a�*�-t�I��%�^�Pס\z��J��<�_�jq��	��l�ܝǐ�x&��@��iS@j��P�C4W8��ʚ�#
LY�߇�{SeW���"w�㕻��>:�̫]x&��fX�j8`m���,'[]���cp��H4L4);cb�������]��iGYf�ބ��4�V�	/���R�`]�
du��a��u��U���f(�C4	
\����^ q�vL7r� Yre�Ǳ����`�'FЏ܏�ċ��,��E��D�ZX+��s�>,}��bY���N�У����߮v.~ϰ,+ bь8'ӄ����F7��~P���V�B�#Z[ى�r���3^��[FX���bϩ�Ȟ
�&��?1�F]�N���?"ggyt�pK��HG0Og⯉���MTǀ�{��R��k�T�6��r�p7/���I����V�ϡDQj(����tf(�n�s\��k�xl�y6�u�z�7HZ�Ԇ��2$��.C�K�a�0���9����� ���E�`�NU����C~�۟o�-W�h�~e؛IJ����-#����'��'̂ŕ����F���P�c�������h�bĖf�������9����|6u|�c��L�ZU�TP'�r�V������Mϣ�3�������.�ퟁ'ݷK�`�?ލ���xqN���־P�,�*�h_�
Wv	���aF�k�27��0���8�a�,U����O{|��9f�QGf>��p��0[�*��+���D}Z'C��Z��ؿ�(�cy�e�#��'���F,��[�蹾��r��k������@�L���QO�0'.� �AE����]�Y@�|O�CDO�(��-��Yӭ97�׊\0Q� ��H�t����@o)TԈ�am�CLN'�L_g��͵C�MLc��l�;��$d����t��/gh|c=�Dq���.��z��5�P�Q��M���$��j;��u�͌���/o�#ɚ���W��RrF
���(�������-ڢBwc� ��Tt��M;�G��6�݁�4lJ��萪+�V���1����M���,�G��5�~���iZ�M�r��;��s��2��Cc�!���u�خJ�-b36��ݤ���v�(#j���2��~��w-��Qz���͡]�A��hC8���{n�ˡ�D\CA�f�䳈�1  �r!�}@Ol=?���gS���5����R�.��q:%{���?M;-�$,����4&N+�*���f�%$.� �.�'�4�d03
w�����h���* �X���W�N�A��������B�8%�S�����r���r��A���r���'��bČŅ�5��@{G�=8-
��f�����)�kC����:H,�iJ� �.g�/�Z&�l�)�[Fiz 4�"���c8��7Y�~N�ߜwA��>E+�v���"�h]~+lk;8�O�Y�Ɠf(�!>�Й��l=�BgE ��Z��5��k��l6i�
PrI#���5a{4�}TL��k��f��u^n��°��Na��d�V2\�Jh�r��'H�j9,������"����~�x�Ϝ/S1��q#,?J�֪.SY�H"7ב�O�g	8ɛ���d�M�)���w"(�+�)��AB� �چ�z_��$�z�myll��G}�PM�������q{�wc,�E����oL.��������?Q�!� u�.2�yC�����^���Q� ��#��ͫ�:�G�峲[jH&j��p�t�i�/�-_�B�+�a4/ƹ�@%w�+��3���.�wk�F4�ȣ���s�QYp&q�(W����A���τ����<���Pþ/�T�z����A�6xø1C{�%8m=ɤ�Hv��C��������V�s�Zs�I��7�4��jF�ع�W�S�<�D�ݍ.쁆� ӂƶ����p�\CÒ_p��e�������F�g��ѧ��2���$��Ӡ!��k��svv.ԏ.�Q���x-��3��e�))L��G��FS�����u�'���2T�6��v��m)u9|���L��9�C�.^�d���F�#:��S��n��@bpw���GԾt�ۭyQ� M��w�����4 /u���"Ǫ�Zq�r+���)��[�Y@wg�1��f������3
���^s�N-��F	^/zLp,�xt�ER��iv[qq��$��
��#��&c3�*��,BY�Ze-N`u�44��==�`	(6;�����B�WW�V�$#�M�6^g�֣f��)W�r;?b���D�ޒ��k6@�o&�q�d��˲�BN��5��VX�	���ˌZ��7�\W?����!	I�н�{�������_���4AI���|v:��^V$�)�G�!_���@���X?=�@Y�5ee>��V��2D��7��>1�Z��pX��n����h4���������-h��z�B��o���������B@ �=ՇZ:����z9RY�c����%2h0!;�6zGY���sZ�Ṅ�=��>�Li���^����yCi���̳3|��i�{�A���E���f�غA�idQꙈ˯�*�M�@G?�"$��F���-s�ߡ��E��Q8�pߓr �Lˢ��W�'�u9�XL�����R��QjZ�,b���N	�<��3����Tb>|��k��Ew�6�L-i�o����xC�_���䈾��C�v��m/\a_�HRK�E]�� RK�w!�����4��-�%1��H�B[w����S�#ā�{\3���y:�fB16sO�*���{�)��+^I�ב�>i�;u܇��+���o���	.��C���X=�O(�^DL��J-�6cE�6�.��b��rI�d���`��<}�Y~D��g�qn���Z���B|oy��@ �ϟ�_C �+�0� 'UE�_4�̪~�%���d�0ד�d0k��zt���%g?��W!�I��$����/`Q��3�>ox�{S=��
�s�f����H�a��z/�>���ʳ���l���/^^�M{5cCmU���q��]+\�����Ҥ���8��l�_����JJ<�`B5� ����9��sQ*S���j�z�]O�n�<���J@��F${��o̐�PP_=�!	������L�ʋ���^�/�`��/3h��}��n��.��DspN�/%9JTc�iH���+[���1�s�H�#/0���M�ͪ�|�]߉Ҁ�y4����p����X�%<98���ES#)�sظ
ǔ�9�ִZ�C��OL��\�L>@�A��^���if����!k��F��#�����h��o�u8��R4q�1���(&r-��� uHł}�"k�7R�����
�oYO���{(a��.�V�P3cu�ț������3����V�@���_�Q+1^_�Mϥ1"I���X�'���-f��t�V��)�^����x���/;h��,+yMx�h�N	,�|y`��{O{��;����?͟�=E���%�� �]�"�rڏ�ޣ��Pҙlg����闗��C���Έ>+Zs٦�{g�3�Id̻�O���+��w�e�W�j�ҠQ���;�Uc:�$���Aٶ�Ѳ�]��z�Q�t��;�w�������j��B�m5���j���+��s���}����� �,���u�01�P�����%\�@�j�i��*�}|LM�����Ѕ3�:�|�k��~�-Ԁ#�1<1�{C�-��\����E�jSڽ8��u�N�s]?���u��Zp7Ge��j��m0XU�Zho�H��:q�9��b��S��jp?�5��[V`f����{����R�U�$��~�f&��u�Lms\q��Ë[���eg9m'6&�,�A�2F�H�%Nb��~�B��B��������xS�Qs��Yl�b?bm4HK�JS)o��� �+$���_�E��X&�TeS��Nq��kXB㨓���OeE$����n[�$C���>�;�L��f��������M7�b{�����"�d�5�Z_I�n-aDp���7��uZ76j��<��[��m���ȓ'�x�P�mޠK�dN6P�&��]!�[
f�.��؝1�?:6W+��w/��C�v����hM�z��k��p�G$��{��~�
D���i�w����}�Nn���F�����r�p�������7��x�@��5���v�_�1]�J�ˤ?�������i0�P����~àP���w����!���^ @����0Ҽ�{�l�-����&��+ O,��KB�y]D*��!͗�/ ]AG7�LOC�C�����!6J���3�(�/��0ǎx�v��v��M�z�ڴ0�����&	��B���W}���M���?��Pѻ��#N��k>x�5{��k������I(y٪?�?g�z+YPߓ� �l�ixF�O��2����d2����K�u�R<Q\o��Ey�w8r��N�ҖlĄ6C�y�z�+�}�6����)���c[� �ɢ��@��v46G`"ju�rB�	s�]"V�����4���3Fŕ.��~p[�1rG�+���\0UƩ�y��y�!��%H�P����"^�k�,(�� &'���"vG���}\mۉ�Hc8�^9��\�d�(:��)W��{��(�g{���t�|�X�#�v*T,fR.T����`XLE֐��z1���u���HB��O=Mi���_ƯU֩�H�F
��g��b) �x�@��gݘ�sՈ~�� ���.�J�N�'c�����(K��f\��>N�7E����b^%;�v�ZF�����)o�νـ,9�L�<a��~>@�������uǌ�	����96��ő�o�6i��L����L��}���u}c�3�������0��� ������9TR\���B�*���d�ߗphB�.`��!ÂmZiu��ƨd����vCf����x����Y}v�W���l�7��~���#u�>喠Ǜx�����2�-0����ZM�P8T����:��C�ת; 﫟"B\��N��p��C�9 t�o�-P?b��K]������˚�����mH���J��'.��Ө���3�(�>���T!�A���:ا�U���n"#E旯�PaЄsU?=V�	e���a$R	(R�G3�D�k�A��M��M�L���1���<��%�1��J�q��K��
F�c/S�]�dB�_[�ռ�� o� �SM ���X|�2?n�P��.���w�|����!^�y��V�߆n�<'Y�8j�U��MNꣿ��Hx�"�F�HP�:�^��l�@BX1J�ư�|]~�]�4D�d���uK��x�m2_�m��Eɏ�� m2��N_���wC�	���.���-1��B_��79�G�m�Y,G�,/:'�[��qT��_b1y4b�����<z�p��/�����Ë
&n���H��Ü�?����'�>���HF[��=�D��AtS�L`�Am��/����Oaf$����.p���scי{�Yc�?Su�pl��h�9/VSkfa�Ad�#0�-�Q��g���)�[i-�jd���Ʊ�ƣ��4�d��-�D�k,�G[Vj-�Ώ�AP����'��{��$t�C^7M�Q����!�{T ���+q?��_\K�A�Ŗ��Y!#�J��֔_ � Qmȍ���Z*]ۤ^[@�_���0r�Lh�.�O�k��n�#ÿ&f}�1:
�T?�||���hD�~��7�Z}�g[P�ͯߛ�� kL�O�^ ������e�Pͩ����_dK�' �X?HD�.;��B2G���o���{k
�6�� c�@��$��L��X�����_�3����	��#ys��!����ycUw�����zO�k�7�/ctH�S�p�yl#��ى�.�Fx]�C]"멾ピCE�/�jB�[�M� ;ʢ��~����g�9o*��@8�ң	���؄VF��W�������})V�`,���h2)D�gW?�|����I��)�.y� ��=gE'`]�)%���L4�E@�		<M��m��O��ޜ2�9�����U,2.# +7XVJ�dF[k��56'\�5;>��!���fp�ݪ�g��5��C�@7�q�>�:]���l��P��f�+��}t�YA!a��
�:
�H��j�4p���_���fJC\dFU!��6=0���_1�r���"&�:��h�`5��2cIW>{ ���9X�����ZT:�Z�~&-<_O�]��rʴ�b����gH��H�H��z6���:�a�lW��z�%>ȴŞ�����Țo-{}��1�PCK�}�>WS���hA%"�<�Z�e^8x5\�o�{�j�`�7���#Zԃ.�ĂE �ܾ�h�e&	�׋�T�P�^�ع���.��\!3\J2��.�()�e�zgY�8���xa��n4�{?�<_++\E,:r8Lܢ
&��6�D�/O�e|1�HS�I���x/�RSa�t �����4yU��o�X�C�w�Kj����l��OK8��B8��#�^;<�v��H�=,����^uo	������8"��	���;EM����v-���Q�g ��=:���<��{Cj���_��r�%w���H&�;<�N+s�k���>[۴�� �
sŹ0�A$�:7�I���S��ݗQ��si��4Q�N�껙)��77A�2�D�1����~b�-�_�����v��#>�M���i����� H�A7��A'�(���!�X�ei�C�e2��bH0e(p�����/�C�Ü����x���^*�b��,��,�p=�y���Q��2��V�}kOh�9tY�e�
[Լ��?�������6���7�Yg����?}��5ᮢ�t�n^Z��wX碏���f��$����
T���3)i̅���� X�ףa?���M�q��*.'Z������^]{^m�A�7��I�J��,3�M�$��.��k���ꉜr)F+�,�zh�5b��8#?��2��ɍ�3��aޑ��t�=1��%>rlA[}��\ld��!Kr��β'����AAҥ���Aq����w� ⪦A�^�
W�"ǋ*�Ŭ��X:x��M$�Z��=[����Y"QP�
:7�l�|d��^�Bpta?��[ϻ42$L�fBD���2w1�&�?4� ���[M.?�Pp�r� ���|�S ��C�-4�h�L\= EW�7��n6@ZD��Jef��<}2�H��EW�4N3H�9Z&JQ	6*ak�V����ԥ���:���=�Y]��Ą�{)�ǁ�5��+k�_eRe|�e^>C�r}Y�.Q���FU��7�Q<62]�Q�^$�~RE)���2	q�L��{gg���v�>������v�~�URnG����A{-�����B�݇��?#D��"2�������27+�qf��<FL�EU�s>�9��
Z���d#-NT��2�"��{���6Zj}�&��Px*�Cф��W\�l?+���fԀ����RËRz9m\��HHl��m_�YEx�D�x������^�o�)�\�a@�*�TD���^�;luk�&���j]ԣ�S�D�b D��7��Y�+�Z�~�1м�B��߈Iw�]
�د=�7�'�XZ�E�b��r���7�bq�3f֑��W;����&�T(���2\����϶p2�;�%���%�"�����y�T���+�����=b���DS_}&�r;C����fn����5�rO�J�l�%S�Ϲ	�%�\d�ͥ��j��?��0{�0�����b�j��K�ɝ*Q/�\�DK}�ⅭD�R/U1�	nTz76����mr�F_����+��� �2AВ>����Pj.����4g���9y�.�x�o��� ����~ �Ʊ���H:R6FO�x�����FN�����ú�y?�(�N��Xk��:Ou�Jp��[�����)��a�5
���G[�iܚf�_��/6���դ�-ES?;y��SL[�Ǳ��ȵ �|�}]B�a�-G�]��'�.ޝ�*09'X�+��՛��2o>�Chp�[� �cp��>ev"��'uB{)Ts��γ�u���i�m�/�7�5��9;�V���u�� =Q`j�1�5�`��q&��--��<���B�_�-'fG0l�}�x�'������ֶ��)$��q�� #w�CH�|�1�ټ??.���&��݁�5}�P��J���Q�s¿�龎Y$wP\B�:��ui�=�_�%`k~B52��sn/R�]�>����Q���I��{Y\39�a���.�=Y8dG�=t�4����%��=��(��bɮ���Gl͊ �e�+;����>�����4������>�Sr�o���ǀ520�nw,ˏ+-o���P�Qn������(���߲j1ȓ���sE����a;I������N���K�����<�lv�
�h�m��G����$��w�צ�B��tFe�Rb	�.�<P�5����˩��r<7%0�9j��YYL�0Uج�؞�J�H���1]{�T[�VY_k���-\�I��L��"d4g-,�K*��R=���,`�|˼�e6� ��wɃ|��y]�:����,���DMnn���ÿ,;���h�l�f��6��cpa�"��w�ٓ�f�&;����c�=˃���~�X"ca!��/2��� �C%Q�32�3�-6�Cʡ�����M��\2�5�3[sd��ܽ�ڹ�M{%���,����U����#�c����fƶ�B7֟^�6��C�#�'�%꯾	��r��>�� �3 �^�f�O���w�^�+Wa���k}>���+�/�Ajg��i��&��t.,n��s�ǊP��$|�~���1U��J�
���b|r�8��3��"3_��c.�f*
[�z��F���k�"�������V�<T�g�{�@�\��:�J���2��;^) ��{4�#8���������z�?� !Q����JHIg��<��c-Np�둶�8#%��d��̪{�L�j��Q᭻�Tj	�����C��������Ç�{��s�2�{�z�.$c	l�L�q�&����"�.��_���d����K��w!�PG-��Qn�-�T���ӱf�ɊSBB�a,T��k�j���`~B/Ht/�$�[�L�/F�!�A`|�\�> I�J�
��KejeJ�.�lᙌT��}�%�H�JH��<�ڵm���ڢ�����U�/Ґn4G��nQ���\e�a->E�.�[��ag�ڠ�z�h$��J�����~n���.fc���ya��9���V%�o� �z���+fd`6��s�7@42�b�����-!�?��i;cIn҇NU�	�0�c-FC
M�ٙ�m�8q~����
Go/��j�p��'�+�$�ܘ�Q�d��1��u�X٠��}�h��i�EN�?][ʸ����fd!x���0b��2��:����Q�	��+8Y%���O�'��sz`?9��~�b�l�8`A�S�л�=�=���]���&�h�Wk���B�ݗJ��P�GI��唱�W���#���"b8҂x!��cRG�r�M��6�j�y��;qr�u��npv�J��Oh�9WZb�5�-�\@�q�U���mP#�=m�
�ވ�ƭe�z���T�:c
*����D�n-����vmdZށ��h��<��<$�AM�2���vL���I��/����=��m�|��8�m1\Uy`A��ԃ�0vW�lbPdg�Z2t�S \s���gs��E����u��[�du�ɤ�ŶI�a�׻(�o�9��L��BrF��8`Z���)�A�<��(���mXy��~y����`��y2�O��=E��ݰ�*�dm�O	W����\�Z�0k��7��>�M"o�P}�Ydc�۾��SOq���N�Go�}��e�^�scw��?�̪؁��F�p/v��o��}�Si
~H8���Kgm�&�cg������I»|�5�S��Sf�ͼ��D����C�ӿ4y��L��g��p��������E��zֽ�0g,e*F���U��i$�#JZ����G�Xn���_���)]��\Yxv_�<L�:��R���*��?&�<ܯ*�J��hAG�J<L�y�W�]s��Yބ(��{��ȱm�X�D�~�=ΰ6B�9do[���6Y*�hE߉UF)�؊���gT������4���/��u �W��~Ɉ�zYn����߹�/8��Ϝwg��^ʙ+y��41(����z|�@ȉ^���6���3]����OM��C�q��߼�kv�#��NO�JU;��S݅��� ��^2����	�u�Z���(�=���W~]����|>�+)Q7m��� ~}]�ג����[]����U�jU�0X0ac�bm-.eK��
��43�j���q��4��@f씰��y����ٵ��5fI��=�W^���9�I����tf�ĸ�3��ez^A@r����q��M���Mf2���i��˝��b3
�Z1N�\�Y��d��p�v���d��<��A>ݢw��S&�\�Q���Ey)�|9-�=�"lI�B����9&�C;�-�M��`C�~�.��ڒ�0A��PZ/"�ҡH�Vl<䞢��DK2�����}-�N�c���;+�������A>��0u�-���Z�+^bV���(}���(�Ɠ�j���~�/���dUE�D�+�3��GG���p����	���>md�B�no�2���O�FA(��>y�:ØAe���
ו�$�)�W����^ssn��Pȟ�Y�1�a��v�r�b.��D/�f�������b�Js1g���-s�v��[�A%�N�֘9K[2�	��o^������BT�١�nE4`X�]�-`%f�+:�v8c���8:�Ґ���s��"�ddx!�/[��{;�Ur	��@.�m����D���������s�n�B�w2lig~=�׻V�N��C
 �zÖ�w�[m��7y[W�P;\L"��w���x���$���.v��D��P��(Yѧ5�>�H& �|�d&Z,�g3���W_C[�~�u�� ��J�je���{�0���wI}$)aJ�|�w�O\�V:m�7n���o�"![�����u��7(�,!��A,�Ċ����ܣ/B�ܻ��&�H�i�r�a%��I�t�" o{��A������3 E��e�/�w����B0���͊�F� ������&DQ"�0�֯8p��ig%nC�`���\8,�CB��D��2][���)R���k����"�sn�+�6*��>���TJb������A=�'�H�n�M�񼁇��g�Y&_ٶ���?AD�Y���X�AxzR�@�^�Ň� ֆ�!�\�i�JN���ʧ��()�9!���,O\	�:F���	��(Du����+��H
�~�b}]�ٱj���1l鍰�l�@�����"�0N����M�w:S��:I'0@{��R���T���xڪrV��TB6��m�=���W ^KcO�YJsTڐ4���.��x�ׇPڨ�qQ�!����Z�H��a?����^�x!AZʢ�n�K�F����q*�D���\f�Y��¢���bA���;mN�:f��Iv)�� �`��f���#�6��S�E����Ԧ��݋W8�`DF2fj��OĚ��L�4;���X�k[?�����'�B74�-�� ��&���F��g�L�ʰ�%�q���S���n;�o�Qn�A,�:��G���Ĩ;������:�=N�@�b����@D�B�
�
ǔ�r:Q��t(��3�
ɘ��>A���	oS�p^�{��9+�[�fv�ہz��K$ۿX�)n�Z�7��Ք����s�MVb��
��{:�`��'�9Wnڙ�T�m-����gR/���ۭل~)+�u��k�h��(��T6�W&�IE�:���]�W� ]4��5�=�J�R���q_�E�K=�!��hI�C�ќ賓0��~�7�H旫�jDc�<[E���R�齷�:�:Lưi$iS�e=X��_�(����Iz���eN�}�N?��i"�~�r��Ċ8����$
���` ;#�I[ ���_��UU��S9�2��S�qRڻ9�6>՗�*�KCɜ��x���:0B_}'`u- �#�b�9��.��v ]��-5��dsz5ep�U�7P�@��ԅlߪ�����X�$i��3y�����bVdܻ՚(�1�Je	�m�O*NV�7Vj����NW4=���c�˰ݹ��GW*f~V�\[U�����~�}�ԾO^��Ρ+ �����u(�?��?N��
|�Ϩs�͔��k-��1�{kE���O��(�Y_?��@@�iW���dT=T�5�g'�I�
m梩�ۼ
dЗz����qs>�ه�b�N�y�'�����[�:��{x�c۾GN:Z��
MBX��/w�|L�G��i�1/O�����2�v'�G����ɻ�l��C���⤁�h��71��7g��;5u�N-1�B$�?p�=�$.���*B�������L ������΍��1���t�!q�JV9�� w��|���6������_��bLxp���vo�`Ec��K)��$S���/΀�V@E�?�P�����gn��@�U�>5�,�i��O\(�M��e��vO�:���Pz��,��G�����4T�9�W*8�ֈ��iD�����2�ISU��D�֙��dM�b �g闷�r[Da6o��7M��"Q#I�EK�,Py�.�zcz�2��C�3�Q��wDEA=��^7��-������:�%H�p/ԣ0_�񚶂��nP��kd��b]���~��_f
T.�̕�x^�we�󠇪�E�Cu�7�yac(�}(�w�`֘7) _��Uj��Ѽ��d�۞�ࣛ�^:l|��(�j����9R�J�T��E��HbM�(��uj�0Iy2��u� m!n3�΄R՟������L9lY�O�5n�PY��,A7[Y��e��}zWx�Z��_P:�����z�;h��)��
�]�!� �S��4�o�HA^@#��(~Rv^����hmZ�:�yGq#�?w�s	ɥ&����N\�q�F�?���j�������@�"�G�Z��9����A�c���M��W�͝�=�Ԟ��n��89�=x�I¥G�{ߠ�fХĉV�.,}~��{1�������uAd%��y�0��u	�-�"2Ct�*"�� ���� [�nX���#A�Sz27�f��
�o���F��%�?��
�}&q��YC������غ�����O�܁$�&�aiƤ�J�E�N'���\F��pd����L���h�7;���x�,��?o8g�AV�m1*C���W�+���ɚ�d���_�W�!��Jj�[���?�RB����Ի�^/zuSE�";H�e��ѽ����w5�d�f��d_d��Twρ?p���8�z��y-�i�{��8��_��Y#�mg$�T��6C
S�$KAՆ
�z��E�a:�3a�����¯/,c�^M��s�u�����&������4�d~�3� .��.����R��)=͌+�w���H֠�2��.x��12��y�tْg��4�|�\8�E��j>��X16:-/y��	$��p*��P��j6!0KJhq�.�A�|��(S��*?��'�������Q
���h�e����#�b&d�u�*�бs���Qo@VYP��f�:���|�m-��_�cD��K9R�K��.�Ay4)���1�x$H�پ�t�Ud�����g������T�'h2ـ�7���""�w������;%EH?o�s�C�4}3��A�+@#��>�R�P��ǝ[���4΋�4/��_�A�#UY}Z�b���Зc-����X����`�[s��c&2�8�Wil/����-�n�����6��R��U���Wy��o���R%`L�����jz�|A�m�=���)�+_
$���x��?�A!kz7z%�@w�(���#Dp-���bB���)�k��SI_a�.sУ&DK�S l���t�	p�L̙X�Ӵ
s%��+��7U���l�.:C|z��?��tL�,��+b́��	Ed�����"������4̅�|�S_i��q��jK;=�:�Z�*a�g�_�.���<ڌ��7C��m���w��g5��:֚��V%�\��jl��K�~����͘�������W�������i�{�%��0���2��IiS-nf����>&��e������b& ,)D�^k� b�@���|��G�1B�t�]��W�oB�B)�]` S��TS��K���O�8���Ϲ��k�5Ew�y�3m�	}����\;YӁKE�aq�ʗ/�] ۋ�4Ch���vRe�P��_�;�-�ޛ���b�{�0E��_����y
mq˖�D�3	���A�1�M�yi���H����Zv0̒S�gV�4�n���ו����d;�5��_(�y���t7/T�� ���s��ߍ�u*q��h��YĲ�f�
@�Х���S�i��E�Jt w�@���N΋H�Ç�r&_�,#.�U(�{��=�}p�1�0�|���%�/��"j0z���P�b����,�K�eH�3a�LC=�˸}�4����Pw�v.v�@�=�b�.U�+@	TF���w�I�!�pd���9��ى<Ǯ�:/��P ��/�rnz�-*�$��G:�1�7��Wޱܹf�z��b%+��z���5�I��z�!@M��3|���� �Ն8��K���e8*/��嗥Vn�j.!pt�-�^/� �%�Uy�g?�`Z�
F�,*���^������T/�5���v�w�KϕΨA_��t��>x�ٿ��Ϝ���k����`��)�����M��%�R�����y���I�ӑ���Α05��p�_d)E�S�.Α�#B�3I�?l[�W3`
8	4��O�5}F>�͇�����`5aQ�턟�C����m�,�B: r���|����&����8��T]�n���%���V��\l��{1���]�\c|ܝHH��#��"��h�s�y���]���t���LR/�3���Yl�ă�B�kV���p�8��/
���6G���M�-�G���Ёoz&1 0�a��%�Lcn��R9�^kz�7�R$�6ͭ�#���j�\r�M�Sڈ2;�3��٥���5������E�<�K��0(�c�6�<ե�#�4S__��"�^lU��K�L���7���Y��o����'���0j.C���f���⌿���_2�,�[y>kC�O�]�wxp+Q�؄� b;3�"P!��;<{y���A���ܔ�B�[4͚G����T��gz���!-�K�<ע����/�� ��:��x��V"vK�j��F' �0i�����^�����~�@�ok���v3�B�c��s��r+���Qnⶭ;\"x�q[�[̭N�PvK*����bʥ�q½�Q�� B���yaٲRj����m���aQ������y�i�M�7�V�w�	�:B��u������6S�+
�� �lu�
�L��mQ0P^ G���!!��6��!���my�����(p��dp��=�x�H)~a�7�v��?8�w���"G g�z�+�U5{#�_Г�dh$t�����p���A��W�["����_���L���8���΄ͯ~�`tK����NWR��RM '�[���8��zF$�8�ْ���%U��q�}?���'my/�k�`�>c�/T9,Ʈ�c������.2 ;�b����6gv2��$j݇F�=�0�jE��F͐(��rCZ�=:������Й���`�h�G�}�w��w5n��>
����r��`n)�Lu�/� �n��,���U�V����Am�0��V_vhܗ�%�9�#�.}l��W�H' H����3Q����8�<�Q�_o�֙�1�[(��K�[���+��Lb$�$f_�jtIZ��Y�S�$�g¢�p�����Git�/����t�_�h��C��A�c�2֝�n����Z��P/le�ri�A��&9zt��<X�S�����"��%d����|IӾ&���b4	<[��fC�V͛Z����9c=�ΛG��k������-��W�5�5���T&O:�[��<;+����(�íM��i뿀3^�W���v��	����P	���xWh�� ��_N }p�n�h6 6�X+����~��Z���ȼ�N���O�wߐZ��*
?�@;1G=Co¨Ǌ�.�Y}b��K��}&���a&����YtecG�]�b����Ƈ�0�2��3A��)��֊�v�8����V��������.o�cJ7�|��lɅ�Z)ڄ��eٔ�R��s��]L q/n 2-�W�A��X��P�z�a	J���q}^�a��O�I�v�[��^6�AR��{�6b�.%��I�qz=H=�I��[���ݗ'Q��U ��mO���W��cb*f|��af�&X��{_�\`{�j��zr۾��>w�����X�KLs���W�Z�f7;�����{�����S�r<�{�����Tx%��+����H�PX�8�X�c�t�q�o���H�l��w�)7s�|�[��*��<5�6'��b8=ߘmv'b2m�����Ҿ2o�;�h9� m�=_!;�Xz�uu �M^鵖$TC�o9�h��w���2L��C������2$�p rfB�%�GX���i�۵F�	�@�pK�8�3�.��O��,�/�D$3�C����vz���@x�Z�5��ļ�kj����wo��V��'�F��Jt�~����¥�:Đ=)�"�V m�PT䋁"h��b5&����I~�|5=(�ѵqSo��M��"d�ud?���lݖb����0�$O���^�a����3�iS����W�Y�cFBD^�Kݺ��&a9$�`2�$���K���Vi����0ȤU7�p���ud�3#Q@`yU8<7T�U��/e�4��� �͵��a�N����;���o��F��vfU|�C�T�}�3 iڂc�1,�準ƞ�i�xp*Q����+b	ԫ4w��J��,ʓ�~?�������q<&v�_�2�<��h(my��S�¥@x��P�}[�4$�	�r�rFr-�r%�g���b剱�?�P]�(�BM@̬`.+gT #.Ȩ*!o���j��h��5���.�)9�^[���r5��샣W���W�碣,�b!}4�+?V��C�(�����}"���b�_/�ɦ�0/"��iz6S-I \+ԡc��PUܤT�Ku�;���/#�ә��n�O��������gm4}'�̩�j���9qeڨ'
(Az&��}�(<�,�1�5y��XLr�r��5�9��[��y@�dW����(R�`	{ɜ0�=8�%��Ofxz�4�n_s�`䶴�3[J[:_�U)�:�$����t�)�=R��G���A1(Rpً�X����J[�Hd��#��JC�ú�Q`�������R{���YB�h�v&ڌ�o��3�D�8� �S�-�Z�f`}�;����qN��e7l^;F���B�B&�
�M'�Xh	�ƨ�� �誦6�ۃ��`'��F���x�v�=�-�q����"@y𛛄 =�&����f�6}�{��zjeX�1`�CJ��u���]`�(j���&J��`�E��8U��Y�����Ζ��������-�!������Ȏ��R��w�v�9v�C�������%��&y��̃��RT� Jc�P��&*ӫ��m�^l/��&֝1/�ZZhP�o3~�{١�`@'Ӆ�
��O|��2�0�V���R�>����@�wY�{!~���_��p���~��&co�6'8���B�,: Q-�*���T��ηW@�/z�8,�6X��[�|����S[گ��8:Q��Hr�Ϗ�9�H�{.�mZ8� L�/_�Q<�>Uf��XA=̼��z9�T��7�b����'����ѧ�+��j�m [_�#�nЇКD�`$�g�3�9��g�Ӆ[e��NӖ�硂�q�õfF,��p~`��	�53��
B&���<k�� ���8����ܡp� 1�̶䨞��f+� �~�G7W�%��/�[x���x�s�;l;��-!��US1:r��Q{:�>�c��g{9��3e`����~m�cD;�l����,��[��k�N��J���QϚOLݕ=�'�\_��4Z��c��_�v�6X�H���B��|�u(��x.I݄_%Z�*����N��O`qmy�z0�F��I�	��0=��Ԑ���ʻfE`!,L�a����=e�B>w�70Hn�T�������Q��+�-΍xa��d����(��R�,"�5��=&�w�8Vt���I�D>]�� ^�`d��=�����#qT!��'
bK��>Wl���f���hҀ���0N����SQ܁Y�� s��P��lӾM²�ah{_.��I�R�n�b�8���E��W�A��o��.�P������{D%)�[�k�]�"�@��T�n��5 /�u�|d�9�cj�����e�.I��C3��v<��Ω�Rd��!Oݰ����b����<�|YM��w�q����,Q�\��'�i�v��Oқ	���6�&��x����,��+ԇͱ�p1�&:�Q�[;I�y��u�������us[�Mp�4"f0��s��%�c;!-�@��}"7PCwT����Å�u�6��"�:տ�J���8��C��٘��~)3a��G�q�
��N)���n$k�z�i(����[j{�i��eWۘ��XI5z�ܼ5Wi-8�:&s��hg볟�/���t�]^�����=̗�*<s�Ol/�*?����b�e���)��K;��oo�n��Q�+�]������-贈�Es����l�i�|ów��_z�:�����L�@�%`f}�(���K�-������I;�O��mXb����|��L�R�V�͇WܴWJ�m�F��z�O�쌌�onR��?��82�fD��gP�HC*�-E���$�j:dn��^nc�@�ٲ���G?��H7�ףŮiR��1U���G���;e�M�fT7<�_GADol��n�5�<'ݓ�;ƈ�Z�=YRS���	���U��F����1�V���P�;�>�h��YoN5�����ۏY(��
%����#�KC���/�;�K��yIU��P5_�
��Ivq�Ɏ1.�i���N�H��"�U�6a?>-�Mj^$'r,t��/pA�׫N)�L�]w��y��dg����{n:!аh��I(�_髩@�A�y$ն6��]D>���A�V�(Ұ�����h�����JG�J��&7Tտ�<�
r�NV�^��T�GhV,p���&�6�kOg[��C��E�Yȴ��/���淪ę����STM�6�OO\>�c��L3�Em�R%5X,t@'^�ʝ	�&�.�U�mur�t*tjؙV2�a��(
6[�ҐXK���.+x�"R�]�
NF�i����Ѐj_�ٙ-�Rc���q�5�:wG9lRl��&��F�U_Xڡ����	�&����ԙ�hWY� )�-7Jj&�,��6h�bVV[�R�0ujF{`�b��d#�E�1 x�RWmU�zq
�2�wM:�+�\��y�o���Iv&*���	(-�G�l$���Ҁ����r��#�K�60��#O_g����f*�C�Ep��>�t (��1�ە9��� ��BI`�U	���^�����F;���%�5V�T#C�.$I�7���ڃ	�2�Z���`
�&�8�$F�u?�;@���_ɏ�/n�"��nΨ)E�@�E�G��)�G��Z���1g{2�`Zmf��$�Ч��B�A�c�y1���Y˔1X$�Sƅ�}Ѫ<�1�WHQGq�\�0�7B&u��!�S�*��� A X��ِ?x�N�i~�p-����(�˥-�[�� �L��Uh�D큢��]!�.���ɉ�ڏe4`�,!L��40?ę�﫳d�*��G'r��~G~�7�.�B�VT�q�'ē�k�������p{в�oŜ�(�T�Y��\�5Z>��j k����[��vQvٴO�B��T���<c*o�*��h���Ly���,	:X.KW
��/�L�fpe۸�5���)wK��e�@�ٞl�Xk ��I\t��N���[&�Srmdo��&:�8&J�ȝ��@��*�c��`̒Y2Ȟa���G�b�hS6���}�g-���;�J9/M����Q�8�P�n��,��SG]p�~͸`p�:�+��s J໫-+Pyt{O�@#�c�j��K�0q<�J��� �WO���ɌԾt��Ʀd�#�oUm�*�AT�MD9=��/!��x���_&�]�3�q���A����I����VŇb��I�����(8���{)�y1\���Z�IlЂ�+���7���`����4T$]6����=����yWΙ�n_�[@�������~�#�9�K5�6��4�����'\e�Q-e:��ݙ}�N*i�Uq|[����ݜ,���D�?��ْ+-3���#�����_��.`)ng~�h^r�h�6W���[��'�?�Q��(��B�I�rr����΂2�g@ݣ-�Zl�(b31a"�� ��bPf��Jy���pP��(�C�}Qb��͠;'p�ȗ���`�.�C�j����ł.��ev�N�j�`{�dy_��2#��p�s���s��"��6�%+�L��:<���b-�6Ms m'��1�1^�ش����8m���f�u�L���(=�r�uww�D���B��m��M�Mt��K�����3�Ķ�L{N��
E(�S��k{��up���E8��#f�:������i�Ku(�S�˪�Ъ���7Ft�� c
وw�z�=��5���@�Aĺ�LW�]�s�͗������h)��֭M���d����{�����vY;�
�K���`^�q����<����gWRu����x�5������k*<qeA#RM ��
�������|��/܁�lФϾV{µ�KH�/�������L���?��(p)LK��()r:QMH{Iô��E�����j�W]�ߙ���:���N�x�+n��&�q�[��́1O:qyy��� �pϼ`�n��쫭
�ױ	YnD�(͇f�Ԙ�_䕐�J�քcE�<��.U�t��vCOm�p�]1�{-�j�H^n�t�^�nע�җyAI��Y��a�3u�Ň ��dP

����a�;����U+[����aa'i�����S�Q�Pł�."�A�K��Y��Q���!���R�1�d���E#�p�����H��xZD�k��K@{��_�5��LR�����2њ�W��X�Y���~���8��؞ܛlLI��f���X��Y�s�jS�>�jNw.Pi�"b��'����U��m��%�:C3�ژ`Gۼ�x����Y�i""I^����/��W:������)Π�- xnr��I�Q<k����p��ES�B�1�J�#��T���J�	?�p&^KF������瞩�J�T�0��Z ������X}Z;;Y��!��c������c?D��>�q����55[n׶m��]	�h��eG/����*�b��_��y���č5�d@���fO�)�^ŜZ�DJ��-@hC���:��G�VQ��ú�-;>�V�	��+��u�����O|��T��zi��C�3�uNs2f�u���5QC\J�,J?ﳗ[K
n��}�j8j�`�����m�<���y~�{���w�����'�n)T����P"Kc��Á����Ff$7.�1���I�%do!�lCvJ� ���|�
K��ѕ���-�x�t&r�ߴY��Y����H�Q���%��Q��׉�xPCwm�&�ߟ�Q4h�j���QǶ���E!b�Q�1(��\��$��M�Ӿ�kq���}�L�y� ;q�'z��/OBp8�"�n�t�F�@��*�����^sG3ZHUk_ĭ��p=d�hR ��DH��2g�Q�	�bڈQ����^5Q�4��|�:��,+/�]�"U�"���(9͊�m�7t�� Oh�C�Hh��.��-�1Q@��i�A���#/�P��[��xL�Xk`6>?��Z	��.�K(�[+شLV̍F�wS������b�Я0��t�5����;WɅE���%��~��	�>��:���Nv?�]�-�J��j���e�(��%V�;�
�(�:���HZN|�5�+$�W��bDE�)<���mT���������(�6$6ìר�D�W[1EXl�C��Q����G���<ٻՕ��>Y�᛬�C��/���8(貢'5m^��BWz_I�*��@vEc�5Z"�	�c�,�UO��WETY4�ƶ��,����\���#xm�~����L�l��8�oF䰷�𨨭���j��,��3���\=D�ea���"���_÷Q�b��5[�#�He?�OO����������ú!T��WJp�P~�s&:'����%��	}w����^��h�J�/{�_�D��\���m�Pu��o��s��uSR�QP��X6E�
Z�4�MT>s]%n��*��B8�9ٗ�ơX�hٻ�98x��l�딋���;�7�D0o�N]ɸ'�R���Ճ�n�j�����ܾa(����i�{ֱD��ĕ(������p�N�)������8d�4a�+z��{Y�l�e���(GAF��=���D%
���~�Nb��?�Q�Cg����{�]��	9��4 �;�U�ά��d�����wg�d��}�2a\�����+ab*g�Q��%������1'j�':����)�̬���_x�x�M���ێ�˰F`������������ih�B_KD (&N��|������۷ss�p}����ʛ�]Xx�B��Wu[ql~�D�_φ(E�ڲF�1��w�cP�:�q��2#c4b���a�͛��7I�#��U����CP��:�01�Na��䊌H�x�u�E�?���X�����dt�.�lk�W(3�r9����7��h]n�,�G�i3-S�Gvjie�������Ҙk8�cYe+V�N�Sn�V�|�Ԙ ����`$�[��K���u��U,P�*��K*r��uMkEQe�h��v}�)a�qEʝ،"&�H5�ez�ޏ�ɋ9�M�/������ag�zcJ��\�e�	��{�J��0��̎�J�H~'�!�,8�:��H��w
�ee��߬���_�h�Fʋ�B�ղɯ	N��D�K3�1�8Y�3�R ?5��
�:6����h���i�ᰋm3ݙ�b�gSFuI���w4g�p�%r���f y���l� �dӣ���䥒��<<���eG�5K.�AY8*:�����p�������H͋�F<�����\V�Gc���S��L/#\v��#�� ���:a<שc 7��<Z|��n0�Z�Y"�9E6��5�����\`f������T8:;>s�j"oS�~�%�s���n�Fq*��P��+��u�+sm\�4�kw��5�|�fHߦ˅��}��3]��]��k�Y����e�;�'b��"�&
Z��M2^�\��8��E��!a4 M�ׇj������ Q�|Dá:�қ*����[�8PL�F��^2�
�r���MTήa�����n���A���UN��z����&*q�0����QG�{Ё�Y�OV�$K"�+��S�{�RN{�U����2A#X�f57&�Q���]��VW���}��ƻ?���ᇏ����Eـ������E9E��{��M�Q��O9�/~��B��01�,1f�?�>����Z�F���K���?ŚѬ�]�X�|٘����&�V�\s愑[���K?�*����ݱ�݋Z�R����Z���M�Iǯ����an#;���{�������	i�7����|��P���g[Q�a��}V_� �
�Ѐ�1�f��K�Ydѵ��Ț�L�Ŗ�v��t��K,N�'�7���`23�:�U�������k ��f}M��Vm�9��Nn�/�niJ��Ѱ�7���|ZP��C�L�C�XE�X�X7�������'dC�[Ku��7\%ԣ `���6Y���z��;d71Zĝ6��o�s�@����M�K�R��5y�����̶�����}��H�2�J�V��@`N��:ve��j�}Dc�e�8�o�B��N7�xQ
�Q��k�yL����h?��&�;�F��q��2��	�g�/)np�&ʧXvz�5Z ),_k��1j�#�&dr��\%�i���LɈǂL˚��]�Ti�u��g��e��P&q����ݣk�D�9鮊��h�*@��s� t	cܬ}g�CsO��|��)��G�$`NowǬ�g9"B��/3��:=6;c�k�B!��n���(L��#q9������"�p����˼b5U	��1 �V
��Y�Vl�l<@:�=�4�Ԡ�c=[����=��(.
�̫�`b^7:;���?='�/�
x�qȆ�nDG�#<�b����(ٴ]��3�y|�Y�Z��Q}0�F�%�8��1�N�g���١��X\����`>Pֽ�TL� �w�x+:��wZn���>��Q#hFTz^[��<��Ϭ�F�vBt2�<�� 9ۺ|�U���s01�N�%s�Δ�Gk�Rl��ͣt�]�&������
��s����J6�Inƣ�fI�a~"`r�!���z�)�9��s�N ���ペ���W�.�Ŵ��m�9ë�c�<���_$~�y�,0yY��!��.��> �zS��n:.�?NϺ�@Ue���;�%�d�\��e@/
E��cs[�PrS��!xF�f�UڼH�3|?�I	q���y�acw�ͺ��?n�w�^g�2�Y� �P�����i�� �S�VC��mi�i�02�k,79I�7=�`#��1�	�8������^E�w��tA'
�ls���Uß+�_���9n�&�1B% �Õ�z��PNo�����@�-�an'Sy�����2��PZR3;�s^�����W����9C��;���gL��v����L'[.�q�t0֞��O�EJ굳��d�^�g=���jw�ܥZ�n��[���������z7j���`���-u=�I�_'S�� �):�|y�&lkzc�z�|n�Q(GM���v$��	�Uv "��|ّ��VNd�F���FY�Զ�q�y�dw�	ӱ�?�+P�Zn��Э�7�����*�U����.�r��{�֫۸���>v��	S~>I8n�۬�~\Z�1�h]7�;�׿��d�x{;}]&kuWH�eb�����fe�f?^�0 �y�,��������P=/��s3�˱B���"�݁?�֯��<�u�eC�Ȓn�5������Kn�KO�@�h{I��_zU������#��8���{��S��VK����HXgv���rK\&��JU�@�|v�Y^^�zT{�';��p�&�͟���F�i}�DY-�Ty�{ij�8�?��(����y�uc���:z U�d��)�.�&�����D��Ht�ҙ�����|V�W䇯�K�W�-߭��N�v���-��S�@���VjM^�����v�+�醹��7/@ �����G��$Lpkk,��e]�!O%�'���'�mſ])4-LE��	�gy��}��
��3�}��[�Q�Ū��Y�_����#*���w��a�w@�gśy.`��{���T��*�e4��ψk���������V�g�mu���[�~:�ڠ���X��R(հ��\��Si��q�X�i���cri����4��^w�.�Y��P��)�����B1��UhwtN��Љ"rR�f�����mIxy�䡭No���R�����zj���6HO�lqH��. ��@�H�h;�E�E�}�3oZGB���Lo���{b�T�E� ��GʧЊ.2k>rb�U�b��Ë��Mb��դ:�� e+�8�tp�(���	���Z8| ]򫗦S����T���Kyf���Ճ&G�Ċ�l�?nT�FJVy������/�Ā��if�B�t�d�@K�<_���H,�~E� +�dףM4Ea�� Lk��̠���Ԣ4��2�/�O��J�W�
�B,���@lV��q�+�Ё̈́'�׫��08��iT|\�
��z:�3����to�������$�wbV�5�s���a�0nv�^[<�
�dC��v��>��Z��C��>�"C���C&6M��c��좫�*�"x¥|��ᅑU�K�m��]pV_��oJL3}���fv4�Q��N���N�|�`� ���Rn\�����D��R:i(b���\� �eq#?,s�^H�˕]�'R���R�²ؚVD���Y_|�Xc��7�~@M������ˊќ�Ҿ�73�*�.n����d7&�@�S�BAj"�F�q���6	W�ذ�����Y����aLH]�?S��͜�CQ�0��XV�7�r�X4l��L��`ϧ�L��/��v�jW�7���͛���8�!�^��R�~�R�/cSJ�K.*������@խbA�ŻP�ɂN��;�1"�R��p�9'uM�U�u�H�� W��T��2�r`l��t��=��wl?�}���'��3���:%	�-'m���ցI,��� Qs�0cֆі.��:2Z���+���/����Fr6\g�if75���䆦<N-�\}�.�b�n ��
�S�\�cZ5��Rz�2I�)K���k	Q
�{v�X,U�W���� �󝖆����a:�f���
�˝��ş����=�(B=��/��Ӆ� �z�~{Nt�lj<�Y ����ھX�/��
,�ƫ|���R/�;�<=WIGd�T[u	w�N���=��bC����.tC%f�x�8[�z��ΜUz+3I��(�~� S3�Hv�|}�/�W�t��H	-Kd��/�;,��aTS[�r���BF��L��çy��4��p*� f���3kT`�.a+҉0e�`����F�yr�J4��Ĺ��x�Go�Iq���i�b����	�r��-�h�A��Y�wDΠS���q�]�I4Ὲ@��r'9Ni�U�Y���:I�7�&�/��_V�I7����Z�\
&�	���i�۬���Z!�D+�����X��:�
	��#.H�F�ga1z)�*������W����s_����ش�����0[W��1��)�=n�Zt� �`�r��6��@��+�P�kr��W'�;�@��K��5�;g��m�Wͅ�t�p��ڹomτ�����uu*�U���&ps$2�_!bc���H\TAk�-��z�֑=�])��B�mY/���n�Z%�3�Q��@�E?�,�~���O~�֞����/�AW�a�:��H�A�IlHn$�bs����ba�š�W��ØN��W�WI1��ԨЇvA�$SA��m]oܿl�������W�)�C���0 M��	�c�?s��|T���O��^���J,��A?��<�C���O�a?�:`"p$�����L�J�����S�~��*f�$���%���6@$�mX��q�?�w��l������)v��?�3;~��\�'��A��U@ٳ��Y;�K�!��Pg+� �+�{��T�4}O�v��ڼ��%	(���D2O���e3f��	�1f��Z1�M�.fu���o>;����A��e�x{�4��#�o5F$�b�&��[Z� zr2]5 �]p����uyǛ12#&�V�xm3�o\Ǘ��փu S��K���Q��Vh�ynD�N�*�H�z�j���D�YXC��ǖ��5��'����Un����y��"�j��"��74/̊�ڨI{��,��|Z��;������_����j�p�O�6 ��H*��N��P?H�~ʙD�'��@C=u���<L��� _���U�s�'ؕ*�cxn�m�:��u��8�|2�?ĎO�@}���2-��N��>?]6w�B%�<S�������,vJ#N��!���]6jߍ@n_���r@#)�U'a���ѥrqi[>s��a�R񶴏��R-�6��3�c��s�Kj��~<�ђmPT�#w�� �Bm��e�?�)�����`W�@Kəe�f�@a������Ez퍧��jI� w���n����bl����N�����̊��
���z�� �b6�Y�s���g ru[���\��`y���H#/������ߺ����\��i�$=yȫ87��7�B��>���=���)zkH/��
�$x�����H��} @�yL�7�ߵSM��p�Nѧ��m�ah�ol�}��g��T����`�v�zq0�c��w3G��!�:}v�q��U ӗ��AU2�'�C��~{��w��q*6R72�ymK6�a�i��l�_X���TZ�f���o���"Y��WLk͟~v�-<�����nS�&���&@t���O�����]/�Q3��֩�;��})_:B ���X����~�9=�����;�xn��
�s�f�*�B�@�$h$�p��lak��n�Q4
����c����ň�<a�;��֠���mR�9��_����9'�st��To4��Iq�3	��uY�}L���f�_Qfg�_Q=�e@=�\��B*^��U��Y2s�,��r�:��n������q@�蠱���?�M�7�ɾ/��vܽ|D�Kj�ѱl�?�~�
�-i,H�o	�9Bq���9B7ȫ�Α=�'��az�n�ĘK�s'�\�
p��n���2�˓.�h�`M�cNP�Z��X�zeE]$J�$�|�d�sԫru�rV��E��W����:
���2��}heR�B�G9I�zH��Az�e�Q�ya����x���(��w�	�i�f˿�����V'�:\#P��yȾu)j�.c�T����Zsr,��d��6�X.@�l�c<���7�"�3*��ak.�;kej�܎����/�,H[���ݝ�\�ix`�<�6WzN+�����K�ah+ewP���:�Yϳ�8��`�sP��w�&Z�6ᘱ��77$��lڼ��bq��4�[b���~(�:'�+H�Zh�O�8���
��{�yS�^
� ����f8�\��$�Aa����X��m�)��A|��(e��04�?��%g�dƍ4��6ƛ�3�MW~ �˪=F#B	m}�I��X�񱚍�&�_O|�@�_������B,(�����s>�I�t�םZ�P�����Ƕ@���h��W���Nf#\2�����m0z�;��]4���BA�?�ʥJ�����G��FF��������!��/V��$j�q�����E�s��}�K�5��]��B���溝0�$��Ċ�������Qȏn�&�w�\H��X��q��^Q/"D���nժ��Z|cY"��Y0�#��wn�;��!\E�g���Zd6�,�E���.��L��|L�K&��Ԟ�ԟ��ߺ�����V�O,�V�_�,�%80f0�iէ\�+D�+i��h3�1zc^N�F@��o}��B_�����mBm���W��5	����|�^eB��ٱ�Zdѥ+����~���X�@�U�	(sH���n�2%�dĶEf�`��s'#jQ����?	E۾8gZ�]���uN����J̘�>�*�/���Fm��x�YpiKRy����j��k�F� y�q��!�_T9�.F��QId*r�p���T����R&��>�����T�&VdϢ��1�{H��!0ƴ��Oe[�6���[�^�fYV`�lb�M���a,��l#Y2��R��� ܪ�U�ժr�,)��DZ��E>�w�@��g����.�tO�L���ܲF�s�򵜖��q"�#���@&!��4Ket]!k�B|����m\(֯k�/&&�D4�t���4/� 
�B9�\��'��ՏH�Ԣڹ&�&23(2	���[Ob���W��Wq�>����T���-6T����2�uZ����"�'�y:^��jQ��<�$�*���	S��LMe��S��!嘯�9��X�妩���ՐK�z��"?6.xo5��\%��+]��'Y"c7\�	1qW��
,���,�tf9�%q�xIp��@�F9JK��6�L8���fx�_*�;��G�`H�Q(&�֙�Ո�ي��0+a�5/*tNH]��a��:/M�ݐ�bQ}�w���p�UY��j��5ݳ{P�G������ҳ/Y:��яGNmP-��	2��[�0]?�AKTa'�}2n�·���bw=)�c=���Ė{��q�2tNB�+��&U�ͪ����E��損��/���^�V0)�����1y`�Q�&��%V���J�ɚ���������D& �.�$��q���7��Hlq5�]w����Z���"��Oe���D�8~宗�4�P���C|c8�����Q���i��;s����y�t��p 0��H��V�N�����B�J� U��g�l�/��d���00��R}h�-;�G�j+(q n_1�Ъ"Et0���+�eJP�BR�;���Evo���:J3z#�-�9̚U�r��_IԺ$�7�֫_cڟ�Q&��l�*�{<�M��l�]� �����Q�'��H&N�s�*g��ϒ�il���B-����~X1ё���dS׻#�2�٣>[��r'=�#?�u�A�E�+^Q'2�0XmegS�kql������o�+"�|�\mp��N�1;Kp�^�b*H[�jDA�.*�^�{�x!����>Z��Ha>r�q�YF��<ݢv�����?A��LW� ;*���op� }��s�9jv�׽b	�Ǥ�;yj� pSg�~>(��h��}�R�_�5k�PG �������o���V��S;iK��c#'!��?Vxa��N�B<0I�<+t�v�u ��52�,V��#��Zl���ﻹۣ��6�ɴ3ҏ�z�دR[lDh���{	�a'�$"{C�>���y����oJ�,��
���_������/�)�����e\��TmD�Ԅ(�>u<ebIq>��2{'��ō�ȓ����Gp����Rni-z�|�3\��iL�⾽e�|�in��w��@M�A�D^>
L���Z]_o�">ن\54+���A
�Tָݦ�@�Jಋ*��Ҍ����vO��.�Y�}���7�)�#�V|/֝���O�F��I��$F7}W�f������5²�2�m�L��.o�hH4�ё�ȳ͆~Q��ؑ���#٪x�y�g�,ض����<�Df��i�����<�A�l�6�|2��U `��>����* ٹ�|�4- ���~"�@�a�\�'؟Ͼ��_;
�Mn¯�P5"O�+�3~uQX�*�:߄�v���	y���]o�x��BX�x�Z9K����?C%��93�!f�XNp��5�O��4 WB��NfZ�>P��F$t���>y!��$&/H ��Wc��j���@T����r6-])�8y��z=�Q]J��hQ,�iƐ֖��}	��uU�ޡ%=`�PZd>8�a��kL3<ѯ3�?�1!�WTUg,�'`� B�"/~�$�n��:�q*=�u��
X�X�#Z�s��N�$p &��}����W
��	3\8o�]�%�� ���˽���f�[yǎ�a���1���P�P�&��*9:60��v�����x���D��������`'�5��-�ƣ�P��&A�-��|�/���[�}���i�G�
j˾�F��]���da��D-$�
��K�.@|0ϩ�f<�3�c�D�b�+Q���[`x@�Α*�f�X���6/wP�����i�=0��x��oj�S9�t7��%o�;�m�+� "�/�r�����pp��?�]pZ���C=�"�{z٨�_�R��Y�;�(7G����k�A�'x̠l̸����HX���K~ruR��M�w��j�_�o'�yG��&�\<z]�9gJr�3�7#�i�l��<���L�� �q$U^g�y�ɥ��mB!�� �=쩶w����o�7�l�N]ᤁ�4�;� �����C�,�6,�HeQ��|u2�^<�9Y�e�I��/�o/�.�cb|C��	n.0kq%��1�s+��b�R��4U6c����34"�P�S�#����dc=�/	�,Ls��yl��Z�)(���_�,+K��y�#h�p"M��{�ʳ��^�t��Ǉ��1���|{��#��������!��U3�0FQZ��y�=Xiw�ib�Y"f7��h�30F�ou�4��y=��'��׳$�kX�:\&|3!�|��c�Z�m�m�e��ZgOIi�L�)w�7���1Y6��ٕh�$?QǰZ�Mn�My53�[�c½j�N��c ���|l{��{v���J��Yn�|����W����F$o�$̕���~w:2��}|*z�tY��&�pD�T�k�| Pf�JMku���u�����4C�������óm���.��'\��衬�?1�ͣ�P���Wx�Xt��;p5O���!��l�� h�e=��g\�&�a+C��"�t	P�%k�w�×��p�
�o��H-���P@�(�^RY"��9U��N�L��ayl���k�B������I�		\���Է7���m��}��&,݁���0d�Uܻ��ޏ�H��PQO����*η�bb&���=l-��a�kΡO�E��+E�!:����7~���咡�k8��3�V�U�2����W���tEL�o$#-��v.^��:�ս�f\���oL�H.���W����/�-Ă�T�IAȵ+N�˼J)ƺ��Uk��"��IQ��O������Ə���+{��*Z@�[�Elns!6����_�YB�+tQ����w{��(s��ۼ��>+��;.Hp@T.G�l�p�tg�5����eܼz��i���wƮ�y�� Û'��'+��س�ߚ����L�|��ٷ�0�f~�!V���RSV��������,,ty5���o�<nԮR{mf��%R�mY���[�hD�u��A����W���	� �X]�� 9ӷ�	�D�����Y�s1naOh�2��r6��� �"O|l"GY�y��,*�P�R�`ig���N����W���aMw���4��;1���^�"�5����R(s[y�'�?��5�U��t�z�x^a]n� oO��	x���`,��&������0#|F^�Rb!�װ��w�@C��~���/'�u�G��p?![ʿ�e��1IX��~֫LP�m��	�!�c�0S���~x��� q�^����Ƃ^{��KS���w�v���9��k��O����F-n�t�j�"i/`�t��@�}�%U�X����vQ'�Y�2�C"�"��o�!�;>���K
�2b�݅��G�H�ɩ��ПŞW�a���������R�jcYGb��f:w���n�m)aŤ�b�2����nm�h�ĥ�P"�U���А��	ue��t�m~�����?��-�`�,ϔ��F��Ƙ�|���ٴ�¶�1}���Ls3+��	S�%C�	�>�ْ�D�5�~�Ѫ=,��sOS���)�MX�\�U�J%`@c4�H��GoYcO����=�������N���*0sҷ�(��E>����;��'�c1�?�ͦ$5'z� �_xy����R���-�9j ��y�Y��|:���9��?�b���R��O��<ğ%��3�fZ� �8,<M��k������r��i��g�w�:+����X6���9��x,yD� [nU�S��*lG����%?�,A䆰\����z�k����"<�̋�����՛�-��_4~z�Φ))*I�#�}!)_���`������ȳeJ7����&ܶI�:�,�����3MV�l�fm��6�'�w�h��߭�D����*����oK�6C(D?Y���-���f	���/�����G$�oi4��=Z@�okV_�f �(�]DY�4uk�&b&��`Ex��9`[L���3-�>{c�o�h�6t�Q���$����}���O�p�����o�ed��G��j��5�\�'� S��{�D8P�莥rC�N�F"�U����mqe�v�T�_���2@<�����Pd���Q�<|*u#Mt06T�f8���Ø,㢖�j3���0�ϊ���976���R� �kP�]���qp����:�9B�P�ת��؁x��+lo'�����ָS�TaGеUr8�u1ĝ�k��S�g�G/�
��;����pUiЖ%����A�m4����
l������'e0h�L/�o�p(�Y�uꍪd�>K�����D���W�JU���Q�B/��$+�/B�^R�S^?8ّ{g��=p'm����i�A#<K�4�� �%�Ͽ�]�����\>6EQ� Ar��|ʰPD8��Gf�l` �{f;�����D�C���t$���94sx&R����K��4���K8�n1��cz�v�e*�Q��%e�ׇ��cr�3D/ylN|���3�>�=�����S��8���a� �H�ؽ����t�ߞ]��`?�xJ�42h�Uҫ�Ky3�+�2%(c���^�a�:p�V�~;O������n�y�w�*V*�q:�9 �G��n�
'���t�(�a�L�U*�F /��،"8���m�O�X�4���&�:WO?�~�����0��[���*�AܨD�����Q<��UF����^7�X
� *�Q6H�/*��^���T���c`N�M�u44����0��F��(�Ǫ��E�:H�����D�6N����Q���׾W؅����w�5��SY����n�ָR+(�<�N��_�1,���v(Y���;���!f��a�4�1 ��v�u`�M�E��s
�9���ŋ>�-��sPp�(?�y���ڣ�d̳^d^;"�����#��7!�#.@���C���x�B���l��� HSȗ��q��C��N��[ʵ��d��q��@��k�SҠ2�b������GEN��@���� ���'�'f*��ӌ��M�O޾����g�>������D��n�\��M�w�H7"0⹸X�����"U�i�Ҵ4~8�^0�5�������i��}��|<�;=��TjO��x@���{��ls�4O}��)���-���J�����Y�1O ��31�֧�(�.�q��bW���M��� ��	�mc���_�P�K���Ѵ9�x�9g��pCD�*�wa�o�/xCV\�9B��V��,$�M����y�_XY"Nc� �"k�� k�°�m~��v�{a��U\s%6�>���lb��#By�&�?p�g/=u�%C�:�Rvaº���f4�Lڢ�j�0�|���>a��zR��:�o�a��q*�傽 �������!a��s�j��&Ɓ��i�����P��6C�h����(���I���/l�4�����On+�=	�����-*o
Q����'��x�X+X��֞*'}�s#���#vT�k�/�-]Y��.qˤ��f*�(�2�Ԩb�����K��n�K ��$ -/��A���j�MC{�.���Zq
+��?�U�t ��������Iè�;�Cˀ�(r��߆��u��x�0���0�l��R��򎣅��}ݞ���݌:�[��E1�N`�1����d�ws@� jY�r.�|�y\(nn4��:�{��`Lw�	(��f��^LR#j����q_��˘�azH��G�N��%/'�ƹ�)�FG��Q���ϵ������$N(�0�;�h��˃��N����K@� gb��B='�j�g����UMt��R�����i�$bL�P���F�U~C�I��%��f�qrs� 0�:	�d�]e9����|�>Rŉ���E"��/�o�@��}�UW�*
�=���	��g
׌.��˒��)���DO{&����T���$/�9 �9e'nv�o����~���)�$����|��a��-�	9�� cZ[���f�#�l%2l��d/z�'Y`���#=WeG�C�p�� P�W"@J�w���5���E��_�C�+J�ސf���ڭґ92�Q�2�HDs����bN�]:�}&�����3�z(�9N��ܯ=;��� �I��N'�P8��I����ŋ$��W����OCG�y�LJF�X��Q��,|���3B�S1�e��)���]��C��8���IZ@��X�b�hF�;K���b���;ے0i��O�6�$�I%혦����mJN��%1$bVޚ�9CW3�l♞c/����!$p�YG.�<9�Ox_tٴx����o2W1h1MT��	_��[�]���+2����)ۡ�%8𙕗;�"�ɟ�*!�̣�/�ԓ4k.�
)�B���1�� ��R?���fIZ�8��bC9j��� N$�_V����t#��g^`�KН���Gfk����YԘ6�9��"t�8��{5?4wߊ_��e`�>��O�,�}=:��ab�FNd�^}����:{�B�P���,4�{��;�ؗn[�Ƅw�M]��U:
~G��_"�>�]���6ע���%Iw�g�p����ο�ض�&��-?�+��+����fg҅S��������#�?ː�p	zѱ���޷�C��1�qB_
 �Е��X����[W)8�<�́/�ʔ�ZO�
9�/�%�����)��u��|��Ugxn�`U+�0P@�.Z����e	��! ֜ċ&a�|悑��ŕ �w]�P�7Akl�T�B+@���-�-��F���.٬���o��Ax��%�d�����]5�ts煴s^>niA��D[�ihtYl�����A�*���T|ѧ�N8�{�[�����Ԩ/����xg��O�F�ϯF������	m���OX\ƇY�xl�ف������1T���0k�w1�?��8���փ?�ܸ*	~{�Ĭ/Ʌ�k"��	�X�>�_����n���x�+�jv L�C;�3�
X��\���Զx\|h���2��6�#q=����E�נ�RWzD@R��u�5�e�}�e�����i`�ܖg ZA����8��aOPD0ԛ��� 
�����gɯv6��+�G*���M�]u��4d� ����Ef;5I3KRw�T	柽��(V\��d��5ȡ���G{�k�C�V^"���P�0�6�V�bGۚ�	�0��l�#�f֛e���|�k�4�bq��Hu�3�W `k�/��=�f;�\)��4�/�>K�SvD���m�@�䖴��0��ӳ�2M;�m�q�s���� ��R ��q�E%����m-ʷ�G>�9cw��`5�Z����k�jPk��u�]iR��Q,�$��)���x��m0�:��Q��/�I��P��jI�2�C��j��o猙d��h��vt$�� ��H	���ܱ^(� ^e1NRf���w"|;Y�m�)rj-]��rD�I{2��k�����!Z]/ݼ߲٬y����(�2�z<׀p�x<"{�4!�oI#���Mi��-a�Z\Z�� 2�O�k�c�wז�n���v�\�;�`����$e.u�.�~W:!�����qT��4~h�v���J9�Te��d��l���lT+r��?��q�0ƪ�T�j�N[Hp���;�lfo�m�$��4Q�Tq�����0.q���1z�O� ]�����zd�TJC�G�i��	 ��x�������YD�ˬ��I��XG[��ؠ�����\��3�
k+m&D����8G���l7|9���5�����!�t+lW'_������a#.X��l��Ra�ó�@�Hc..�S�h������&�� �:�L�z���2��@���ni�d�c����jࡌ�x:5#d���ž�2�&�|�%�;ӈ�$��5�K!����,���)o��ɟ�%�;ђuǪ�pe��u�*�gZ�QB=�A8�0YG&C�#�?�>(��Vx-޿�� ?�m%��Y���|��%�eD���ot��9���&�25��+����2N����T����VΖ��̓L�$��	1�A�Õ�J;��*�ƀe�ϕ;�[�q��IG"ǫBq�>��b���+���K^�^Ue�ȷ��x�@�#��ӝiPb���}��_��&m��'�cn�9�N$�É�Ln�
P�(�ۏ�'G-o�)t�:��l9p��y]S������A�ջ�ְӷ��L�C�%8f�H�]�%���*�����6��:&�Q��x��~�O��Dv��Y����EuE~<vm�dUﾨ�JlX�}��d�����6��Q����:�Q���5�A���)w,0gq����^h�X
)���&�*Дe!-��խ�P"����j$��Yc�h�4'*읅����?���#��d�"zi��5��-�/x�$�#O�w�����Rj��$!|FԢMU�t/+_3�U%]��hb�#��Ŋ��>2HG����}@� 	ީűg�dl���#Ys�D-95kj���[#��?l�$����x��d���Za��Rj��<�z���W�J�+;�1�j6�9u�v����-�4Uc[i����Uj�>�=/
��(����i>���m,iH���p,�hO
�U븡�:uMX.
��2d�����+���f�+�22�
p 3[���n���(w:��vΊ����p�M�T��f�B"�,��b!$�_�i����{���a��vf��ɿW
�r4}����A��}�l�|��W��Bb��U����V^��^[�S�H�uߐ��''�>������SNzG;��8.���eR��Z��r��d�B��PO����w�d�3DVӃ�[/��m�k�J��� �p�������莮�u!Q�l��Cu�`I/1���H���整ZЃ`1�-�{O��C���}�$nJj꾑u�����mҁ�~��e�>�	+^�tή����*)����ϼ�񏠗�AӼ�:�!�i�k��4-3�X�D=e����
�����XΤ}�d�X&Uh.�\�\4qe_��L拦�������~��&+�vN�>R�}oP?��g0��C�8Xm�d��V\9��T�pn9I�$��B Q ��S��]��v��vF͓������fL�Q�/m��d6��=J�͝����x���2E/G��,�=��Q �z���"��h@��J(=����0Q!���o���a�M�����~���YC{DVZHSr�Db��S�Ķ3+��b.Q����}��Z�����r��?bG|ʺu~�؝���R/��Vn����,v�����mU5|\k��b�h�t���K�fZR��`൹kH��/�����/t8�	�O��Ey�(���n@�0q �	��Ϫ�~ÆxH��aKB��ff�O�ߔ��,���cc���3}�j����ŶE<����tQ�m�+�n�W��.�q�z�G&���A��\Bܗ%̘��}$tBl�� ;�����k9��p-��K�WŕO�DM�(�m�į45"O���5�����u���>�b�g��.\S�2[�^�a��؞�ب�K���iK=4v�4�p��^M�>obT��/�zx�e8��Z�)������u����Lŷ�"M�%U�PҦ9��-���@�.�k�dTt��$�*��1ka�vK��\����9�X�.�;����'�-�(ʏ�I=i�!
�:Ls�`���
����y�3�T�ڿ�#F�q���L�Al�����$!�D9�G�[N�]���%Z�N��o0)N�,�uLX��V��1乺��h�̭�y�E����.ys����tU�����M?<�!��в�1+��
�Ʌƞ�D6��)��+�黮~�	]P���cYe���!d |IT�A�%�7ܣR̎# ��$��1j�vÍeFLIo�8;{�#4�S�oX���o�,8��x?:P�-�Nґ�"�,=��u\��6�9s�h&S��a�(�: L27D�1]��$�GY���&4��6�`ɋ��Ւ��0p���"���幦���]W<����@n@��$j���l[��̖Sw�ه�ݖ�f�>C�!2��	�'�sM��@�Օ�+O�sz���p}�%�Oϝ�d���y��X���
�J�r~��/Ν4�]���~g��6n�ve𪦜_)�TM��y�g���F�V���E�Xs4B��!}Ik���C��aL�a�G�L
}YY��@���_�#��])��mfȓŖo��sP�n�Cf�7��� �	�����GJۖ���-63'��(���:���L�%�(O��j�*_j����"(�ô�E�3!�������D �+K~n�®>S�Mw��V�FvN��T�s�{�./�4	�u�5�}��RT>;� ��E+�	��x��lɫ�Ȝ��
�6�+_����3����_�W}�%�q���z�^�sƇ�"���L�H�r"-N�M�DL	K�����Z��:��x@��b]��Γ�М-1c�n(W"2j�"0�����qDx�F ��(¸
��BN�r������j�\���Y�6���w��Ef c?�m�$��H9�O�5C�[}0#%���a�����'�!6��=��P�A��Wu&��֒1j�YoN]Z�����H�Ɉ�"'0��=���i��B�x��q�	U��O�=D�	�׀�{M(H�6��㢁��l�ّ��htא�.�%ڦCWA6�&q�;X.J��F!�����k8��*��ag������s?�`Ҹ���_��!ái���W�e?�)�wH�
�E4@�Z�=u@d��)������7p�Aj�ۛ��<��Asn�6���Lf�eb�	�
xg;9�
�0d�u]�k�c�:ԬK8�L��W`PU�y��5��	��x�5z�lP��1O�!�º$'S�ň���W^.>�������oiy�����������w{HV�&�gn淯�_|&� �$Uy=�Ͱ���0�$Q�nXW]����ۧ~��ƅ���� ��z>��ܞ��q��v5��gF�ӭ�����\�<@�*��.ºE�O�[W��4rR��z%֌s߁@`)XL�ҳ}�ܜ��}V���^�!� 5=z�˔w�؈d��X2#�{M�j7:�yFN�k�q�|K��-�!ad�
��4�0Ȏ�};E�&R�W��l/;&��Fә���:��i��_d�M�דX,i_�N��^�0�az~j�����>�;��	
.ӭ�Y��%֓	����33�bn?f�nד�r��
'G7��۴FDY���޳����)���n�T��a��?��z�F�WI�l]`U�����H�Gș�a�c�c��w0sh�!�EUp��PҀD���j��D)L�[��ɛL?B"|�p�eT��;e��b?
h#½�>�������E�l)��.�o�I�\��?핋�yv .�5��A���WBL�{EDۘi���7%�ʿ��;���U�4B���k�q /��g�7g�w�RO���	ś�3�kZ�l�)�IA'd�a��u��)�
��Ł-��N��Ħ"�\��m�Z���p�T�4s�QN���wO
�	.b��J;�\4M`�����o
�@�%r��7��G��}-��^�]�˓�A<W��T~pњg�r�A�H�Y�SB�!	�4-��unpߠ��q���
\%�m�Tйf�"[wWk[��k�c+�ݪ_���t/ܶ~�ڈH<>�1�_�_^�ݺ'k��rC��<�4@���6�a+���uM߱\2�IKxfʶ���B�c����a	�t>yZs��0��	8�;+2�Տ����t��	�|�>4��5�{����*�N��F5��
B3�����Ԝ�m��I���F��	mqt��P?a����� �#c�1�P4�'����o��9x9��ѷq�VAA�￦A��f*�p��/I���g�`��B��L�n�Q�CW��ܨ즳~�P�h���g�.���
T��ܡ�z�h�P 3Q�� k��s�pA�7+��x7�3>KI�FEQ��[=t3y&b�]|�����0�@��w��j�@VA���"�d�%p#�k��n�gF�t~*ħ��	6�?���N��6߁�!4y1h�y>�9��y�~@(P׸��
h2Z"b�E�8϶��+��15� ǦGp��H�y�A:���6�,�7��	���̯��I��D�D�8o����y��'b
�(x�զ�;'�K{rӌ�;T��h7U�M�W�x5�ɥ�Q����d���G�|����ƂŅ��-��w��Y�(��By)�W�[]SAnx��<����������G�'LI����3�Z�g9�;wp� �^�,L�����LO�8���~�1������J4L�2+�e��w�X�6uo�q�Ju���,G5o1��U���Du_A����[�>�?3�G��_&�P{`%.��q�6�,w�o0��f\L����:B9d(�/Tg��m��8�U=�=r�󏅫�ik���@ 1�}
P��5ARwb��3����W w~�(O��㳙�����?�U���e˦�!��V@���a04M%�H�uW�Έ���yB�F���6�!ȴ������ҁ�O����71�D��ˇ魂���]Y;�.8� U��8+���u��p�^gl��a�������f��\T�|�g�i�fR'��JA�ՙ�'�8���';b�  �r�f���Yk�~:���-�Ѿ-䐶.I3�kU�^0�w"�iLҿ�cW�����v�;cbc�1i�ծݹEzZ�?��a����^��g��Y+C����2\R�¯Xs�c��o���vC�4��]���I4��gF�v�J��0y�|:�+p�.�M�TѕES+u��Ww���w��|!H���sT�����~�A!n��5�k��t�����A"z��|@�ݤ�}؅-����:{�A׮�gU�*<7�\�!�#���η�6i���$�Q�iԬ���p���6��c�I�Y|
��A'F���kd5��|�:�ym��=�aɃ��{)V5`�c�fm�hB��/�6$�oܰ�S}/IV�Q3�uT&��n���͉r�'�K�{�4Aj9|�&O�tm�\{���e|�Y���,��p)��W�ˌ�~��Ic[
\�O�#:�kL��[��
�+x�3���f__g���r��ȊF�.�\^�K�#z)�쐨��r���ݕ���Rh�/DYpzA��d�y��� �ŧ���ID�Ȍ[X�DS�:�� Sε#hΣK����zP�?x�,o�Щ�nP�N'�W�9��&���?���F�����g�"F"U`=R���q�3��!�M{_��˗g�Ĥ�4qtw���</���t����t9i=�\�� ��q�y�kr�}���d]fD@֬%7C��ׄ�w�`�D�>D&�~�|?/ccDm�0�wK|�I��iW��[�u8S�2V���y;�My���rF<�8r����EZ�����]}�3��4�S��\X�es%��4�m����ApVQ�lBM�9cN���$;8p��3��K�,�/U�����ʦD�cy ��$�n9��OԺ��OH����sb��X���f,ي���g}��_OE��� �ۇ��q����yP�2��>�YZ��,�y���w�q��b��ĭ�l�r��B'��g`���KE���칇c�-�	��n����ʤ�7 -�Bh���O����� V1�t,O������O���<�|2������r��u�ip�x~E��k{��ȎX��9�Dۨ�Y&��Z�	 ����&�}��ikרϧ�%�\ �&�%j�q�hK�{�����r��w��m��2�� �6��|�D�Գl�����g�~�5>wuڛ���1s��a���F[Pd �����/w���y�>��FC3�h�娺E}�a`�BVS(ʅ�	^�9
�;Wk�o��~�����ʉ�\�Pl?kX��(�8��xW!�\U�`'؝D�H6*th=�J��_Z�Dt�ܝ������^b�W0�Q=R��r�;E�ͥ�%��u?���E�=o]�O}U~�PF%i�"���A�}R�fAK�
Fp�������,�����3J����^�5U�# �ֹ�g�%1��f@^�?[ǴN�L� YT��S�$Z�#��>:���*��"��j�c����k�G�QȻ�R���������x�q<�2������5'mpY��b�=��AL�o&Zi�CRXD[_gg%�%���X�K�.��#v�e��Af��k�j-%�q��N���I|�ī��PCF4�}�4S�z(��4��ܩ!x�I�_a>��60�*�dL(�C��u��$����1��c���H��`A����5���1ϴ0�Q?��:�"?)V
�a+�KrO������7�^3� �)��:��j�ʡ�=s7�qZQ���x��֚;��-�I�`�&h�?J���H0��l6�é� r�BYF�)�c��Js|.h��I�ހ@�xg��[�(�7*7Q#��"i��0~˗0�jM�����|����3c�*eϭ:�Ϫ�m��j<��s}׈�>��J[l9�>�-�&�Pש�kt���R��x����.��hl%U�_>Rŭ�=�l'T�C5��Z����D����As]��!۹�7�]�5���1��$�а�b��%��S,�X/ϓy�g�������靾1��(��P�����F#�*|���
���IOr�Z4c��a��(J�	�fq�i!���v�/,��cZ��ұ�$�/�����.�`�R��d�Ä�
ak��O�i���{<���5���T��Gmެ�Km�i
~��7��R6x'G|#�L�V[I�T?��@p�*�� ������p�I�dVGR'O1y8�CO�U�_x��+^/�p���c0"��$�&.Z"�2쎍�>��~�rҹN�ⱇ�n�>�M��e@�˝��}6Mh�lv��x)�/��)5�$��x��X�������������e8A�fξp��=���K��6C��/�i}�vT�r/�Sј+�6�h���C��i�O�Ga�$�q��B�;�� e$t��` �T��U�/P�1ꡝ-p�%�ƺ��
v�9���c!��������М�?��p�_^��0�]9|��I��%sti�Ң9�$@��w�W(��� f�Y����5�br�VwsL9 �l��-y=���}y���Gt�6��?ђ����u2�e��A����
P�"�J��%}t%U\���?�ka�[�	E��myrήl9L�7v��/Q�hݖg�%����f���S���&@�k��ğ�`�Uu��j&2�Vؑ��F�?��@�|k|'&�OɕM��M����%%���.0�@9>	���s%U�k�3#L���fD<i��K}�%u'eQK�BU��r�����	�E`��o��!شg���Fv2��W�ŕ���c�h���\�P��n����p��4�k,��V�	U b���T(.ޯ��UE'hݎ�p�� �h���cB7�8�M�Ӻ�R#c�,ʪ;�
/@�J�G;�*��G�t��O�yu�ڡ�c�"
ze5�?�����k��	�����whk% o����*�`rI�أL�ޞrm�Աd��|4T#���uп�U|�/n?��ə��=��N7M�����g������key�<�w�n(�������H��˜9��o�;*��1z�����s��"�[��mk��҄М2ݫ��D@U����+Y�Ӣ������p�q�x|�U�ᰚn�۴w��w�Ų*hI��Gb�	r�F�dS���߈(^.��ճ=*������,�w�C�.>�L]c�|ŃE,�0#HB^?�w2"2�AJy�򅥚P��*��&���з�
��7��v7,ӻB �:��So�N��Ϭh�566�o;�$05�ȟ`�5-�ls���/i�g-���EImR�����`l���0���#^�+s�G��|J*��>^K��f���6v���4�Vk2Y�n[|���InUբ����l��9q�;��=�DM���RT�'��ZRB�0{��b8-����1-j}~m�J�e�gm����w`���ѕ�V����:��qh�o/Z����&7�P�']L��[迃5�f��@n,�E	��٥��`�笠�)Cd(R)�e6��
�(11��ߐT)�(0нa>:�X�yǓ&���pIK���y�〽Nqta'�+��o�������aK@�?����@-A�op�ɬ��r$��@�������J�@
N!�M�7������ X�)a�vG����+<B�I~��u/�,��N���y�����D�,j�ȉ�n�C
-�՗��jc��' ��t��ָ���?�ۃP>�G8�4��Ṭ+4t��	��?QLr}M�I�	��cIu&f���ۀ��\l��3��	�K�;sj_�{3��c��W'��e���=vh��]���rW��ӱ����Xb���_�	s�qSi�~d��Dڨ��Ǆa*\���M,�(5P5�ȵ34��1��t�=�8W{��v�M8��̘ia��e<�1/-3I&��8��J�[��l���N�W�i������t��-1�ǲJ;�Wݚ����\sD���D�"a�yH����?֫Mm��+0<%<�Dy�d�>���qJ�������.{�톒�A<}�sCGcټ�ob����!�&��@+D56Z���jԽ+�Ⱦ��è�n?K���s�<G���#F�u�0ԅ�~8�Yp��<��}�e��V*��x�`ϲ� LA��\앦l�O��q�����F:%Dq��g����-���l��É�g+:@��~	U���I��V�^U�$,�G�1 �B �zc�W��MƮ3���F�lz��]3�����2��LB���s�1p���(���=��st[SC|T���*�ۍH�'�kL��}�=��6�����Ч�aѥ�*����o���J��XfnO���ʕ�}j�~���ng������{̈́� �>4Y�ݷ}��.ϓG���)��*����X���� 
�� �g	���t�j���� ��I�V�%�����`�7���b�[ѩ�����P�[��&%"�	@U���<5�8�}O�2�YQ!S�6�����`�r�8t�5���j�ղ�a�|����2�W9�X�¾a^m0Xp��!~�3CI�	h��
b�na��]6sP�&/��`@�[Y=,��vs�e��X:%5�pM	H���А��,=��j�_h�&�TS���:��غjJ'�¡SJ��םA���4����Y	S҂�.|��S����~��Lt��ۉ��2c��lSu����cwn0+�'�H�N�%z�g�ǋ$�3��Oe�?&B�ҲY�{'0\�R��o�1ZD��q� &+}P��aGf@H���(�q�U���Ah#������Ӳ�/rVd��}�=����i��&�[����-�eh��-�cF<��))���p��<y�Y�B��$j�"Dt�k8�x���T3^pkEzR���2h�0�����������8M�*�� B�&rH���>�0v¡��V�c�-��8L�p+a�x/j�E|bn�w�����zPj�?��M�Q�2��~/�Ʉu�)��ή���Xp�m�6�3~��*�)R˵��&/�L+ޛ�ĤޮQ�-Tj�����-�VI�c5�>�>��J�I��+��d�Ơ�//e���IM�x�5�� Ɲ��:u=��ۭ+ug�2�����u�ݤ�b��j�|y�R�Pó�Z�g�F4��N�B�W|���>S��?���e7b������~�R�ķ��Q���L��J���2�#���JtHE�����CR��6x���P1W�dA]��Q�дq���^\dNZ�f!��ހTh@mc�y���4�Q�Sa��ԯ�����R��^�3y�s���b'W�֒1#lL%D���ݑ�Ԏ�F�&q��L�_`�t�O�,y�߹?�C�~/K��=����b+��0L��]=��s�m�x���cIޣ�S�0 @�0�V�	��L��>�eJ���RPi��OoMLhY!�N�X }`H��
�@�~z�;��e2x��J?��<�
T�&�E\����X="t��tG�����)�N� ��ȳ���7���w�૧��d=C�1ŵ�\�&���ZB��g��I�(Xs���Mp�y�W�]:�:�A>Ҫ����)^�T��w
=�6�!�Q��7�IUu�!e��8x���z��.RW�3e��j~?4[ͤ�W%�4�g��]��w�~;,:HM�>?�pig8 <���l^{L�]wsJ0Q�W#�WK�u�!.���|��4�3EV�,�C�����)Չ��#}e T�!ބt7����~br�DQ�C:�#":��(�Gvݭ\�Ll32�.���d|Y��V����w�J���Ȥt9��JR�5�^)��#�P����!��T~=&q�u���6��*�"F�؝�b��~�-]t1V�/��O4@eOX'DR*���m��l*���za�pU+8m%s���V���f'�F�nQ���O���DNAI�N�Λp!,K�M���/�l�[m$������yơ#�톛��!���䯨i??��"�v�f�{m Ԟ�j'��@�i���]S��ͧ;�B��L�0!��X���/`s-nE�U�c�u�����~��-Ԇ�|)�-���Ȝ��_�?���Kpr���I(S>�������,�ɨ�g�c3�M>��y�N���^=:Q�\&�λ�a���(�R�h�o�g�Ȳ��őu�nX�19�xIA0�\VXyi�$�A�_T\�LX�I�~��%�xċX�k�)�w�rZ5~9� �VZ7V^���
0Wfdi���h��Y�V��'��{�Y���������#Bȓh���Qs%a���d�c���_8��}��=w�yo�6��U��\A���r����UKR��\�!�E��d�`GѠ\Ā;�#v��o �����w�r�ܬF^@��@��G�g��,g�?^7�O%܀߸���7���^��LH�쵚n^ڎ"����m��?�G��p�N��Dx�LYD~�ɘ�E�X�)/ɀ��Q\�7OR��K�������
	�?���Khb
�2u�ۑ�P�I�Cv�m ���������8��J\��S�֋��^�����e�)w!��]�S���8b�ڥ1֤|�P�/N�p���.��6�R|���e]%R^z�r���\Ҏ�9���������̏�n�R7u0F������L�W" ���A3�i�չ�Z�+��_�J�9� ����R�� ȃ��4tU��%Q�ےM��?����yUD�;����K{�4_ڱG>�d��Y��Nٚ��o�L�">.��zH�|�����=�̹�Y������!	qh�M�ձ�0&�����rr
'����[����y1�%JC.�/����V�Hd�in%L�����ä�(~�
���WG��6��NR:��m���۠\����S��O1#����'�]]��|
�rK�z��Ɉ!�V���/�_�2\��������1�$C��;�T���a���vp�H�� }w��z�pf�.��R�hC�u�v�l���N>q𗕳��*����_GH	���`AW�/��8}��6H<Q k����{�%�u� j��6&������s�W��J!�ww�A�x�+]���4�7�,���V"9�@��M1@�+� ئb���I����`�#�f@��z0$�6��+s�G�P_+�Wm�F���~��UC;i.���~;���b�@�������h����v��	��ω�6I�fC���2CX�;��gf{uV�����OD�qm�^/G"N� |��^�K��#p�=4���a)t���Q��c6�C\<}U�l��an���"t6 ��H=���&[l����Ғ!:��4���m�Y����/��	�D��dBZ�4{��sA|l�)W��u�뎔N
w��E��O�* �mŪ���q=���9�@rD"5�����x;��u\F��墿\n�I�`��h��@�I�d��ĥ�Bw~�G���dT3�L��[���Zĝ� +�:����i8r�1�p��m�[ΠJ�4F�u�^��1_)��T��t����x���;W}�9zW�{�M�*?Lq'Я^��%�j�P\~5�;�	�o���u�*�`\�����uyI*�ҝ{�BBL_� �[ɣ���<��6�D=��G�M"o����T��8��w�pD��R�V��M�fMS241��_���F턧��� '��;	 �j��7uQ,A�*��Ͷ��n	��W�AnL��E�Z@�Du�=Xܸ�m���&
�.
L_��63��b�H���5�RNcR�{��hKl=q�;���q����p>��3�)V[��Q�3@V�pC�ˎ9�(�B@5N����cD���(��YB/�ĪI�Iuc��[��� 녾R��g���)�,j��C3���0������������p���J�qH�AG/�\r�B40�t�����B/��ՠ��&O҄n�i�e���p�zW>�ܕ7q_�����x����g�]4��T{|e�H�)��n��T�H���� Å��)�(�8� t�і���W���9RN�fT� ���>�ʦW�w�Cz3ڑ�8l�'�S��Y|%���N���G-�'b�Q�6�a�?�M�o��2CO��F%�w�qþ6WU�"모.�q�{T�bŪ�W�"peu��NS,�#{�eS�!OC+��\��2?�3���w��V�̴%
�z,�f%���BB��-F�%>��G�II.�,�
{ S���h�=c�����߽���Q�\;6n��%����E���E��k�HW(�cSV}'m}��|����Ƞ�����=�k�Ŧ[1:D1[�X7u��'C��?�o:f?��Ҩ��>�ջ۬������AaJ"".��E}=�*
�QH?��<i����޾�C�Ke-���\�!��%�v��%��k8j�+Ϊ'
nR��q0Qr���o�K��6F�����A�^�^ �[�����`��a7��;n��z�۩D`�e+M�)&J�vG��4(�I>T��l�?� �j@�}�fu|R>����@N�D��~������W�aG�BM1����+��OO[�B�%u�ne�%�:_�>-��] ���B`fP*�?�x�L|��_��0#�0�H'���g�O�Ә�`/��w�F�\\�D���^�D��1�)��$�]� y�!=�q;{X�}�!'C,K�Wi��zްQN�>�,C��\�,oO`� �iٝ�Sl1����鉴ID �^i&�[{�PNx��C;���d��pmK��g���iV��`�i�`>��ԣT�69xp��c��é�	��PXvȟ5a�1�	���K����⑤�y��=��:X�8�%��FW���3ז^�usF�ºs������)J_г�T�J��k�t2�F*�6�-|�f$:0FLz�����t���S�
��� ����pw��U�䦉]l&�>[C���aA㡾T�S�J�=�l{샮F}{�F��e'��JO0��f�E���X4%�q/d��A�蚣3��og�����e��;h�V� Y������vO|#���x$�NZ��XFbO�_�IŠr�}{�^S�_z��:��R}���$�$o#��k�F��+�r����]jW��؁s��C$.�m<_fI���ض���:��&�p�I�`^L�o���g�����W�9�L�tz�R�qL�<�پ���ڍ�﬒_�y�W63CAb7�x/$�4����0�g#mo��0�/��Ơۃ�*g�fݫ}4��J~��-7W�NsΨoy��Ցy���X���_RF�O�K�M��@�l�J2����\�6�ʌ�]�x⷏� :T���׷��Fvąݱ�S٠�V9����g',�*��_h<W|����4�/<��q�ȀАQ��"�7�a
K��y:%@M���@䖻�@��j�3�i��1��Y�fW��X�;�r�|�S�g��8��}�Rm��4T�V���=�����U��Y�=�΅;LX6`p���҄j�JDY����E�:�sf46�O=�ؿ��<UxЦ�Yu�]]�%.���8�d��:�f$�w�D-�~u��U������`�C^q!�SHi�(3:2���r.�Y��$��r(�+����ܔ)Y���C߃;���t�,b�>D*l�XnrE��K<���tB,�H�9e�������n�'��x,�s�<� �4 �=����̙�Oi4�}6�@��G��!����R�0�iw� ^�~�S@=��R-�����:U�*S��،/��U���B8o�-#�e��3��;��ݪ�������aF�ܔYFO�H><We]0�L�����u[Ti�l�8�V@�F�e��,\r�a�>��'v�2k/�?1�0T^��������gֵopZ�I`T|���R�ɟX��H
"K��ݢ�O!uD��Z�/�,����*�>��4Ʈ���<��g�0p�H,Z��ؖ�=]( /ZTv��wF�'S�W�a�H�W&wU�m>`�y+�}5�+�-0��b�oo��2#�3+�Yύ<rM$H��غ�ƄّC�V��y������hB���dļ��uV�H�?��G��X�S��\�������#�HeE�N�r���)W��<i�����'F}_�(���w�1��(c�_��V�IrO�ἩP��յz�/�/9��==���9@ةl���AҖ�ﮨZ�1g��c����VK���/�Yɹ�b+��(�	��&�[�S��Y�1%ńE�y�`3e�.��Tv�x�`�tK�TZ\*/�5�5�,m$�'�u����k�ڑ�x)Cc|��F��l��țm��}<�GG���-�~����e��gM���䦮�<��Ǆ�}v0B�b�"l]�[��ܣ'��������-�`�?I�U-�x(�F�����z�*)`fqz	���W����L�D�X�e���zׁ�:�6������-e��P�_
).p��7)��!�=`��rI������~���ś��O5�|	K���X�T�8�njn?�b�V��O�0�{&=Rq)��^6`
�������?5&�5A��0�"�����{�!������c�L���k�F�X�Kˋ�����M�E㤹+3��!�B�u��-ЭofJDY0�܆���G�?��S�M��*\5w���r�$l<k��x#aY�gQ�
�u ����ׂ�&m��9N;TF��{�$5��f଴�)�Ln��g�(�fO1�Z#�PS��q�d��J"��~�o�]�D��p���Y�c���/����R�8�?��m~�c/���=/ؔ�i�QP-�b��r1響���RK�9�������o�����y�7O�r�%���8�R�2��#�d:��f�}pl�(ܶs�\H��`N��-��p�����s_�����k<���F;u�?�!�b]aB\�˖<��0l���o��j��-�H�������n�<��#ku\i~���f
����'ֵw�2sd�)m��E��N��Yc��gT��F�N|ݳ��
�1/����>��jM��k�z����hx ��зoeo��~���tqS)xO%՗~[��OR���ѷm �R�����.�ea�:4�/	��@�6��V�X�1m�Z�:w�OU�J+�/U+Ă�Dg}BPgw�l�<�c*w��H��~?���ΙWN��P��5�̾P	�T,�3w輕�{�A�e���a���Ң̷�Q�ߝ9�ER��Bt�KbÙ�N�ߐ�-��p$�j����q�	H��F��0C�M��K:�k~:�*���b���Ñ�
}G���;ٔ8��ub�Qʏ� �V�o�ߢC/��J�Q5P�Y�(X'3�W��3�����J�ޙ�c��H�5���L(Ig[�2���(�RL���n?��b,��k��jK���6�#��(��'���+���E��$��ǆq�I�b"��nnÊ�(=5\Q�	*��~囥eh1=�ǉ�1_�I$�`iO>�v�#1]��$H]BB,~���Նv�e&(���H}�1��;�e&'�<�n�u�@�I�\Wī.,�B�+@�*A��T������F�"�H���e�0�_K��s� DeV1,�����/�t��q��'����"���h$IلRx<��Z���D�w�c�˥ΊXZ(��ά^.���<���͌���P���_A�D��D�yR���GD���`�4`
���P��m��,2�ȅ�.s�)	��9\�<��?�2���x�T`�7�N�������Ci�9��ԉ��]}��W����0������R�g���e]ꨬ��_"��\7Z^��M"RM5M<ˇ���t ͐h�{n`/}�{�t}Dp]xb�*���%����}�Q��T<7�wČ3mv�G���� F��],OQ����w���L�ASZ�����WsjD�~N" $|�/V���S#�}��g�8�켺+�s7!1PPw�,���7:�L-���.�2x	�H��Ya4[�V4j�CwI�g���
q�_Z��p���ez�ĀzM';���7s��Sx��0�f��`�xK2F���Z��G�=S*�<��v�n0�1�N��(�9�,#�ʴ��'���nyJ�.��-לK���ʆJ|v�\r��ѣ���52�v�,3B%�Ɛ��
�)��{b�?p�PHZ��J�7{;x��;d؎�U��>�-�]j	��؅��Q��k��љ�Ci'9	�oӯ�p�y��] ���1�s$�e+�N�U�/9H�w�5�ER$�Dt^��wG3��Tz���u_�����KZ���%�Y��x_@������j>}�bVd�*JyY��]��k���M�f��UF�S��������N79-�1��-�x��V����p0�w��rmJsO��+7�.�Z7f��ʪ�� MrN ]'������x!����8���@)�~i�f����:�����E���:Be�)F�}���܄kJϜ%:љ�m�\^b��f�O<S�ڰS�|??��{&�[��H����igX�1�6��<,�	��/�t�⴯v�6��T�/%(��0PF	�h����\H`�?ߨ�?��&����Qס�d�>�MLѡ,���ק}%���U�B!oG�K�PZlp�!�E���ړ���)F���z��wY@=X NP4-��xB�q�O������U��-�y��A�X#���$舥�9q��8]k<�^�֘���v��)s�]b>��:�7Ű��+�{�gNV�ɰ�c�Ru@�[%W%k;L�Y�=2�[�u�)s!�r�j���E�Sboi
@eg�j=�F@	=�P��y�p!?��͹6��^�E�P�F=Q�͓E�6�Lh���c� �j|�������G<���>�d��K����L�F��A� �c���=#�i\C�x�$��h5h�S�+w�O�����QN��)M�A>ܘ�7.�K�i���@~����p����!����V,��3孩� sc�|{`�wU�R}��u�?�"�K[v�Q79�r����=��wE�� MoȐUo����ol��͔�܊���/�^%}{� k�} Q˜d�/ou_�V����}��
�x݀�T�>��϶���7<�k���-ԧ^�s��>*W6��g��>�(��L��x�">h��������B��Ǚ��`c /��6474���A����w�<�#�N�I�n�l����f�SJ�2Z��yct�Bq�A'9y���;eKT[�~\!���iuH�b��U�W������:�/+C�B���e�F
��E-Q�i2巁���3P#ыeK��^��i �(�b��`�$Q���тaqJ�)��tTv
ʦv\I�YA`��m��n�P�'%�D�7�e�E�w ���vG`����-�����G�A��;�K�9pn�H��G'�6�	��_؆�zi�)�[��,���Ra=����7	�L����v�Z�.��PK�Na�6��y))�(�l�o��`��b#VѾ��W�S��IlŨ�(�hY��fcXC+s�`�P�N<�Z郶YR<�Z��0ُ.�4�� X	%�Q�qu�B��`�
�Q�$���&װ�[Z18f��'>�8$��^��#���8L	߿��#g���d�� �0�͛�������Z�`��5�j�B� �Z,��~����!
݁׈)��kb�s���#A.��T��Q"��[@m�Ux�dy�1��^�d�帇,̓#ͯE�e�6��!�W��Zy4��\����P,{C�ia���}�w{�(���"����&{�A��;�MR�"ΐ4����Ṉ���R��jmH��]��Bf�Q�Z�_�^Z�����fw?B ?��X������J���y2���ׅX�!�i��۾�_��ZO櫶n8���w>oqS'��)��b:y�#<���$. 搤,�H��S/GAK�:spi
vɥP��͑=���S#c�M�S�|���pQ�>n��و�w�!w!����J+a�p��_v7�=������4��~Iu�{��Ф�Mi�y�'�W��pbvN�	��G2�kj�T�h�EE�`հ��d���.���uu�U@Jf�ŎQ���3��Ě�젰tߘ��~m���lQ�2`��ƞ�+-��7NUO�:2�1�qg߰ -\����&�?Y�bO
U�a&�0��*E�`ƃdÄ/���-5wslQm��������Ѓ�j�v�TfE?�)泈>,bt��M�y�� T��B1w�߃���bWK*� �H��-�Z���R�(���F�iqx� dcL��|���׾��@���v����D������}�qo��*���FPaA�4��\��zЅ�N�������Լ��-+)hZ�6��eq���y�$��i� �{���~�Aᦼ;��Vi�"�g��j�}`e�^��֥��x���Nmt��|㔳y�J��c���<p)-K�i-t��GRa�t' �$��)�f6[��iśT�/Erb��'Lr�O5�yaX1�e����8Շ	^���h�~�HN�6�ɬ2�@*$c����]��kHNC�My��DP��e�^+�������A3��h�u�sEB5�S��`��"t�ǚh��A�9b����}�}�t���^(��ů���C#E5�E��g̴�:�;�q+��1�*��ᗏ7 Pߖ�؏��I_M!��
�]0G���D9�o<���	��UHx�&L�^�K���bY�)��:�w�؄����Og��չ��:w[EU�����������j=7���k��Y����ֶ��c�B�DI�x��t����Őq���0yL�퇶�����/�T���3ف[�+�/y�9�) UgA��W?����݃��҂�������+�a�&	T����$�ʱ� �ybKm�F�]�/��w^���2S,ʐ:G�����;/���Siwk�뾏@��-x�\��{���k���&�)��� �H|�:�8'�0N�YNBA�T!�F�]��D<��H�ǭ��vx,L���nCn���F���P	�G6$ѼBm�h��:���m��o��<?4Q��6����p�	��!�P�P1oQ@�7BQ�W`�|-(��&�R�R�!�J����Ub}eFN�T��  9W<�В��$ �u21��'A~��'��QA���%��cq�����L���t���h��2n�r�@����%��ς(�X�{�l@������!1�[�Y�j�5�H�X`^B�R��m�Q	��m��;"����x��"W�I�H$ ����r����sˋU�7�%���4����t���i�#g�{|u��?z��<	������mW�$�b��#e�9������s��	-��6
��"&���od"�4|���Q�&)D�u/��}	(���6Z�Ȕ���>��s�]f"nlD��XZ�cT�2�2H3�ιd�SX�lP��=,cU���ϑ��nk�'E����w�>��a���~U㪽�M��ۤ�:���&6�8�����7h��c&�4M&&���d��#9Ǣv���X,��2�_����� 	G�%�cqC8�4�C1���8��7����ͣ���Ɋ>
��v��iaXɦU�������a��(�D|�z���̞݀�}%�5��jM���i{��VC�n#}Օ��^Tqh��S��R�%�w9^{�T�G�$�J��b�Ԁ{��hi,����GM���؁���?�1�br�Th4MA�%���F��L~��Y��i�?<��6U٩2�b��U;;pi���7D\6�뽃�/qa
t�c?#�
�F8���/�u�M[�D*�Z0o.Djʼцq%,�t�0����h�S��T����5�����'_�ϓ�`�rh��l����;�5Q�cĘ�M��?pK^���p_�q̴b�c�緽���WS�Rz��tt}ŀ�ҮH8~�A��gQD���Y:J�i��n��&fc������1��+�R��KВ8n�������t�o�U;�GoA.�iCF�q�b,O�up�U�!F�;4`jүa��GGLk��ގ�����RT�U��#��[�(��s����B�w��i(4�s&�����pd�F]3�o�bН��l��rG&�Ӆv�r�_��Ⱦ����Oΐ�}��aV����kb�F�F~��[����s6��Z�+�+���xѩ��	��C��ק���`>�h�R�L(K�=�e�7������:����#��Q�����ԥ� �C���HK�P��J� k����T�;����X�Bb��nz���RF���o����i8o`��ǯ�"n�4&�_�@��q=�隳��Z�w�y���k���C�十^|Ze���E����?td�����w:�U�lK��E�9-��}����}��.�����%�ۈ^.-��׽J� ��8z�o!��p͐z�6o�UN��ag�+ѓ�\)Q�DÓOk��C0`�\
�Z�2B���Y��Ť���� �4!�j��?V�ʛ2����q_���{���C�E\w������s]����r!������*�6�o�\��ΕV�*~�K��h�/��u�~lƢ�en��dd�l�v͚؊�{�C��v
�lR�1�b�Ӗ8���C)��}DK��\bzu�8��I	�@��˴&�i�D�߯y���Vi�4Y��j�u�(@8%�Z�����ev�� <+r�݆�4���gS��a���Wg4��y4�8��B�2�A7��׬�D(���!|�������Z�l'G>�)T%g!w������j�E(�v&�M�߶A%;N��t́+����w��E��!��E�]e̬�!!$+Z)O�<�R�ڳ��_`�p�d<`����k���b9���1@e�Vy��F�[�1c��H��{" |U��y�_����@��`:C��=�\�	AMz��+��cT&֨�C�ǲ~X�I8K��"7��Q�C��8�D�?������N9�r�4�%cs�B6�KO&Y�S�mS�!P���Y��ca��������� 7F�2�I�o��%�H9������x�F+4���v�a�R��y�	f���x=�T6�M�i���0�`���5��[a��i��y���f�T��9&����0�\�����;:��^:�X���n���ٛ��fNw������q�2�"wJ����zs�EP�6{h��k��>����t!�{���0�kI���~�2<��7���`ۈ��4�"�JӶ��ȗ�O��
∳�2>F�RY2m���X���C��~��pZ��<���,v �mk�N� &�AbK���j�V�f?F�)V9M'�F�+R���hn����j�η��)�#��xk>b�nj��=���\�� ��Ml��K��}8����㯇8���L�����^�T�<�5��y4�Z��)�m$592e5Tb�]O��j��ځ�tg�D-f������O���ぁ���}a픔5��7h;y�4"p9|[���D���Vs��q?�������8wk��dˎ�7?�I'D�Ԝq�[d.����7�c�c��`�,w�iE��n@���Δ�h��L%zX��[0i�������3���T�}R����i��ͧ\�^���beШ�W�8{�����W>�ٵ�a�}랐��ַ�Q��r��O59kn����5�?&�\�l�uJA❞��ܿ����F��I�e%�#�@<Q�Fů4ښ)�W�؟\K��_��C��Q��e@�%ЙcЈ(	]��O���L`A�B��߰��Ʋ�����A�V���Mʷ������à���Z%U��D�����v��?�vW���JO>�T%�����8��qQ4*��eOw����%ީj�oJ'�>>.	�	p��o,6�[�"D�S$��҅:L�����I���D>�Bn�l�G������G�Ď�)LOa�#����af�c���)�����42v|�d8~镰��z����;U��'W���D��H��y�]ͻɷPe�I)Յ3(x2RSvS�:�'\۱��SÑ��)�5���x|�h4�B�'(��6���'`hdL	6��*�ҥ�M!�;�W�ӷ+`�-`U��Χx�uHD��U����Uj���TG�.0�>H��M�W��m�*A��2�UCc�D��t�!�,��<�tv�&�	����B�d@�e�rx��`��#赝ǱE
L���يP�)�lFDz�"l6v-_[��;�DԖ��Wo�u�C;����뉣3�O�`�+�*u���e*(��Q��fQ]1�aF�XC[�r|��4�<���^a��8L�p�ٻ2Ԉ���o|��]�MISǚ���A��[&����^������!����#%@�妬��Ȋo�M���ӓ�fd�!�8=��!j
]7��>+{�a�Ij�IF��_�� YNeZ�uQ�HI�����+] ���[�`�ƞ���%�����dĸ�܃��;��p�oOa<פ� ���h���,PҞ�"\�a"?x�?�K��~���@D��py�u��Wy��|>y��(V��0Ƥ����^)����✒'q;aT�ltړE�����m�W�Qm2�_y�Զ.l<\|��r�U�g���c8�C�|I��zFUj
Pr./[�c��`���
(=QɬF�	ܜ��sn��{5�&���Q<���>�I��ND�p2r�����1�Y�42Tu]ǽq���A� "O�6m�HsXa��bK��(K��n|�w|ݏy�����YXR��Tq/p�����㵄�I�э�OͤG�@|�"���.��ieL`+����������#�e�����:/�I�����		Ɵ}=�lf-W�=�|9-d��C;}9y/Bڝ�0�K��@��5ڤHF�7p��`pé���Z9��ugb�Vn���S�U@)~|��\R�v�7��7��Q{+�ǜ��c1"/B�!��'�t ��c�yHr�mx<��x���p�X�vfb&����?��_�.��e��6H*;�ճ���R�2��p4������_�{�7#E���M�Z76��xѶ�1�1�f4���������:�o[��ۧ$N�B�3�=��J�M�e�(jډk]Ҏ�/M�A{g��\�
�1�u1�
DM@WG�g���(�G3�d�izB�
%~�sdc�ݖ�w�:��&���:���uB��`�Oe8���{�ȵ8�SY�ל<�VN�2����F+�	�O�F��f����d������TCG�A�X��c�4l���*�JɆ[E��{�M�,��c��MƱ�7�w�r��MG��C���y�0z�g�b���q�.�~��`+ƴ�|ԭ�2���|�5�+P9F@u�e˙Z�s��qH
lC�S��������C���@yTq�/s��l!�x���D���Qj�,]�6EkN�OM^�e�o� ��ؚ�Z���=�l������S6����� �4�y����Ce��N�:��9�<�QlW�����8I
/=���r�C�W}$Kە&� �VL��i5�~ I��ڣ�	e���8�m�zq����`	s׵O���"���d��Y$�)�"���>JO0��q5�IG����ؐ�~�F��R$��2f2_}��z��[�tǼۼh�	����ʈ�M:�/Oj�R�l؃�VNا�F'�s�:p�.�M��.󢧻���˞���鷵����������Ka��[]%w<�Y4)�_�"��׺�x�����V��
�^���,�@�O�Mt?�I�(�'�ƒN��O�,��4.�2]\�=�]����X�qЍ-U�3�!0I(��(v�\�hڋ�Ԋ�y<	H����h�h ���啶*�E|^�KZ=�+/���bJ��l�9=�'����`��Fr�an��Q�]�$E��Q��i���q&B�u��9�T���yյc@����%U����4l(�"�r�&>���Ӻ)���KG�f�O3�>�n���NV�4��@ܓ&�!��V2{�ǳ�->��u�p��!��Ͻmg��Ġ��ћ�V; �~~l%�>�4�_�����J 	X����h<�Kr�&��f����Ȝ����@������Gz���dl2�A=]N�{%�X݁� �mT��	Mge}[�u�4�D�[�:C��gζ�Ԣ��I���U=lk��KG2�@S�q���?��DL7�}�*D�iG0$���I��5"�-�@�G��Y�� #�>"Ev�O�v:O��n��c$/R��Z)��� P�3�uV�/����/$fX��B��Pl�#6xX*`��
� �o���(�}������/�m 0,�[e]���B
&>��nE}���M�g�/C��<���S|D��2��Pb+Ŵ�c;��i������	��Յ�2%�l ؆��l�((�گPj�!��ݟ�3.�*�S
!so�o.e�	j��B�����Q�7�15��]Mڙ��֗��Bb�X�)�Ģ�Z!�i�S��e�I��H�;4]���P޷4Da= �Ҁ�	��s;�%f9�÷�~j��o}��>��2�lT���3f�Lg;$U�^�W/WѶL}/Z�(F���������w/~�^Yd�W�W߬���zY�G𸛌�ʭd�&ʃ�����*�!^�e�˞l+��g֍@i2%��&>�p�T�`��a�b�f_GJQ�{�붪�Uв�A��a�OЫ�((�6��
�߄�|�����?Kn��	=�w�e������
:���,e�Ȥ"�y�����m4}�))��B��]���-5<��ܜrH��+U�@6x�?��tH��Z�k�8=�D4�?9�,�H�����r\��3��٧P7����0���o.���)�z9���.)�h��{�[�x�'�tǀ���b<� �	���H��%1I��h�L`��a�R�V?���~PJ�`J̹E#������w��Ց��n���6���"��^�~��ƫ��*�~,�J�{�v1i@�o��y��!@��㉍U���|�x�XR��I!�RB0\-w��[q��4QXy��4����{�7�D��E�y�G��E�O��x�wS�$p���ʖj��e��vW���{Vo~������>&�&r�����"�Q
}�B��
U(`�60����w��7�h{���R��A�dw+����ՍG�l����I�2��Aut&�/g/@�� jJ3��h�%2�'��o�=���y^������׎rt�gFR��ZK5�F�u���%��C�\J2���B�7?ȵ�My�b$I?T�\ Q��|M���w������V��v�@Jk����uI>d�lLǥp�[KpB��b�a�]UX���'���P�e̴���ÿ��9�����Y�6��];#�A[3��?"��F>V<����ͤ՚.+�[o�^�@z�� ;�/�,*�0%�&m��}��]���j{T\��|~`����D\D�����#z�����q�M�|�F:I��Z��S���ĶY��ğt� �f��7���".@��0�7D{�Tr����7QV����&+����uw��@j)�TgH��k�AӬ�
�}�{�޵	<I�R��+��A�t./kW�� �(�'9�b��k�g��&���~�x{����Ӎ��f��ɮ�
6����u�Ȕ̫�%�5��H��&���;��>GĪ,u���c�F�V) �<8�F0�W~�$�Bz��� l����c�_/���,���S�o#e��q�97~���b�yUP"����e���n���KRTjk]�p�$8�ޅ�.袮Xj�jDpY�ߑ� ���&�G�T$�j��he�)�����f��Tֳ��*V�<��� 1WQ�F�iѮ���&$��
gwDy��e�aV6� ���.c�NE��D�g�����
�.����h+��׻䙗eqK�ZAo�ץI(Z����_î~�c�s�dN����3������T-��.��j9>�<U�Ect�$��J|��J���e�SJ&�g�R�_�C`�*b��]����Ʋ3;�
�Dѕ8�?�)Z��	���x�m�x���sk"�+"��1w�*[#*��I>J��NV���3��E�VC�����tz�B�HZ�Ah�������ꢸ'NW?��VF;�`���AT5�:-}�a ����|;�a�#�*>���G&��9��zr�3�c	Z{\��++�r���9�B�Z'���1^�~I�����(JG�2�1�fI�'`���V�2����#�}�k��4�!�k���++z���,
�\R�"a��+�F9���Y�3��G�*� �(����u�g�)lIAoY%ü:`�94|-�3�`��v�rp���	�U�H�i4�
Q�cM�'��E2X���,�k9��\��B]df#��
r�����|y+ry�r��PN��v��8�d|` x�/)H{�)���˺,)be�.me˘�pr�[5#��X> n�/�h��������,O�g���V�z�xc5	4�Z�8��m>�w����U���7�ԣ�����,�qԹ���z�=�����_YQ�|�`�B'm����h�=���Lф��5�*�@J\_�?g�{�u]�|N%��Q5��m~�d~Yz�Tk������\��',�3��LgKn�hq�X���g�_��$�S�ę}*t�~�A�[Gn{	�-�Q�D�ƦNlk�����}�?��K ?�����.�wW�z�T������Ce0��85��$G�d�R�Ւ�	�Tm?���&�	�ԍ<�����$Y*!�}M�۱�M�����3��9��ӟ~�ʥ�`ú-0��ֿ�Ԧz4;����P��i��8'�̿��f��-VL����~W<t]�նL���B��Љ���|�R�����~]�3ļ�{,b�9���h]C'���f}�&JD����.'���͡;��7������_��L� �kT􆲞���k<�G"F�o5��on���
���oh%(R�`	��2��j�CH�_�2N��>,�E����O@��(��>N���E��h_y�Gʎ�RW����j2g"���_�Q��:I�:M���F@ѱH6������ݗ>����\@��+H��PA�۰t�t�]�QǱ��`~Yn;�2XT &�ھ̕Gβ�I��e���4�+i���Q7�?�*Tf3;Z�[�y�ڣ������:d������<5	�m3�
 �\9����b΄�}��(W��ba�O��`o�C�K�b
��]�G�����d�9h��^V܃o2s��v�A�FK�u*�~��GG@��'�.�L�����XT�.��3�/��0�N.CΛ�\ڽ}�1")��bu��Gz�,���v���Z���ͪ�ܠ���p!)���\N�'��`}��D��^1�WB��u&������<0̣�ϗ�}x���J�`����<�ޞ��>rBdC�P:O"�H7�(�!I�^�ޤ�/���~/�.I�۾�K�[K��H:�q��I���	�=�*��`�rGJ����`!O7>6T3�Z�,��T����y�FT�;�ԯa΋7�D��7�
��"��Ҡ澖X��mu���և�W@@��6Ŕa)�^�Ls�Y�˷�!'vƆ"�HT_R���Sq; ��$�'F#���4��-o�V��j��@�	l����i����
�ܓ'�U��\�1�V���Y�>�"Z )��5�\��z��R����K�U�6"YW 5�����:�nP�[��M+o?=7\zqW�,rr�T/�A��G�H�9Ld�9j3�;��]�Y	��OZ�f�6w��Bٕj����ʠ�t�j�&�{9����B�=��v3sQ�3���`�C�����댆��a���~���w���dμ'|�����Q��92&<I�=�9�醍qY��s��LKiFS��n��k�q�*�3{n�19�V�������3���s��
+��}ħ����|Gk�{I��ZBȹ25-7(�lqؓ��!��2$P�C0@)�6��z�!*B��Is��YG������*,��wQ�-8���5�x:�8YL�%Dc��G�{�c�$�EaݻTf��%V~_���c�` ��|t�D������dh����r�mx��Ж���Y������L�
4�w�ƚjv�Q��0֨���g�Y����	�~d����I�n�nۼ�������Մ�cq�w}T��]p��.k?�Z�������������7��-���NM�} 1n:JA�e��������W��l9me��Fp��+�xD~�W����VWU�ȅ�*0�d{����P�7�{8p�Hoh@ժЯ��H�z~oϨT�iC����`,�:��C�ׯ2�]��;�p8#ae���m�M�k���
��z�y�&^_+E���^�:�Rs�̿rHq��M�TGT�jp���cCV��A�w����ː�����ԕ�b1���cY�D���E�Y�,�yݹ��-����+{��*?��"�6�[P��Î�C���'S��0\��8��O��Py��Ct�M����>��tH�*�z�21�4?��5&a�Q:H���@�o�^=Qk�a��z��)�OX���[U����S��v����>W ��nm��95�������%of���XճsԐ�"'Z���&ڄc��`�q�Uݹ�Ʉ�O������Ks���u�(�i�M�\�|$�	 ��>���C�����X]�3�:���q��p�=��?B��JP(�3�&�@>�ϻ�ZO|�=H�I�_	g��@Ē����=E҆���Tf省:G��DD�I�q��Z
5wBڗo�Y:x�S�q����Gt߇�0�.FW�9%�;Ӳqęh��W���9��η�Sq-�6!��q�Ś�z��U5����[�hB
ƍ��8������Vp�!g�6�q�WMx o(���a��?�s����S�5Ü�(��J�ȅN�J�J�	�I�߈�IQ����
���]>����ؒ(k���4j$�hW�Ӏc	���^��\rN�]]�W�j:8<�Ё��yC�Gem�p��B�7;,�$�?n+kw0�Uu�A��^�0�#�����dk5�� D���� �|m�%���NYQ.�\G���p�?:ls�ܩ{�y ��6V9��� �[5�Q��m��	]$�!�$��V�^��@a~1lh�e�ۮ�����?��&���pm+l����AC�0Gz�e���"9>��ɒ#�4<�.
�R.��d�ٳP݃�!Sl~x���f�|��ƣ;�*���I�&Şn�`��r�RXm"���v�Ox�0'�Q3f�,��O��b���dQM�%7���61���q�fT����@�	�w�O��"�̌�)�ܩ�J`(f�9[���X[��V[5��Bp�'�₠��><��5ani��#W��<˳����GX��Ű<Y|[���4��\�Ю�Vy���%8=!h��ҏi)�d��ƱBj��~���@5�n�/˥\�/��%��'���T�0t\�ڷ���M<�K�c�j�����m�~�!�4o�:�V9��y�g:�Ŗ��		а"� �d%$�c	{u�כ-��&7�f���ك,������f@*%��CԊ^�dї����l��ÇΠ�=9è�5[y� �^�*$8�BӷҬ����l5������nP�Xho��2"�\�t�/�,�9g3�ͬG��hS��=�hT�����>�`�h�f#�Ǝ�b?�S\��?�x�ch6:>�;���@Chl���\c�FQa^�𜈥�@/�$P{�6Sc㕦Vh-�V!�V���H�?�
���k���o��B���NX��?�I�l?�Z���I�<*�p��6�L|���`��]Q�S+t;��N����8l�`^��Z�Mp8�� �o\	1�i���W��`/\��߬����ptP�[�{g���}�[���8⩇Θ�^�������w����]ڃ	)�����m�N	9�!"�I5��\,V(�.�4����>�����O�N���p���,\Wť1ZE�oe%��)H���N��dВt��#ΕuW�Y2�2���
���Ui�����������/�X����8�d�S�AX�w���j�	d?���|"-A9J��yQ��
E��Q�m�������$�#���)]/ؗ�J��%��R6�P���j��SW@o�
�kU��UZ���r��?�������}��63U�w�!��]��[�3�q�}+)��v�%�3'&K��/�o j��D���]��	��Jj�K1��gK��TN ˞�"�c�;҃	��:�S�W���ʍ��gԠ�:�jlQEyb��X��?(M��J�@r�k�q�Z-��Zw���/��]$K�H�$�� �_ �P��J)��gD
�T��$����3퐣�P�Vߵ8��6@��C�� q�y���+�	�׊�,x�p%�e7��,�I�z���`~��Ij��F��T�q���_������ᨙ�n;I��{ �EM�ﾀ�\�Ɍ��uXM���F�\���7{�w����c�H�/����7�2%b�{Aم�䃈5Gn�6z���&FW�4FC�킷w!���k� q���~��oa��v����˦���ۑR�B)�^�x�Lk0|R��댂�Xg#6d`�Ø�cu��(#/�J�����f�3�`L4�P�?CǾ�tRo�	r������_�6���������x�Z����y��Q��K/�)�,cUԄ�L7�|��2�\*@�E�����K ����i�&��T�6���U�#!`�2�9C���
m��[���nqTr��ϾT����]�j���ڵA��cBrtP7��h��<ovz�R(*���������A�i�����BZ���|��o7�`��/P���(Ԥ�$�v27��Á�/?��*	��n	G�H�#2�I�����J��{�D(�L��4a6Ag��v
;d�}@_hH~#z>�o��;߶�"����ɄW��r�i�>ւ��pq6?�n���y#��r6�OjJ�_�P��� D��u��qj����� �`����"����]��3�p�<zE����m<�p�nl�՝f��]�v�Y}P9?IJ�Ѭ��g����Y:-ޗ�v ���g8	iɌ�s�yi� \�uP±	�t$���j�.���[Rv�$<��JhI�nw/��G'M9�T��\}������W�V[�ԹN~����y�כ�1C3�$�s���^b��U~�30�y�?$�L�_Y
�ASfa�D)�;������� ���e]Cw�ݭMf�7�"��4IF����k�y�:�+��۸9p�q쀅�jڐ��RS`�D}��Jm�tt��I&�!`�UX9wyB������Hf��7 z�D(��[��;��Qר������;���������c�
v����@��v��$!�f�����L�S�6uY����v�X��r��@���V�Y��J���'jdIV��	��=�z;�$b��&~�&�)MY�!�uZ�c����'|��4rL�����x��tߡjVN��זK`Dm��ƞ��)p#F�0ߦ�h�@���p<���y�*P�*}V=�Uy]R�enX�F���Ϫ��ݙ�d')T����m�gΊ�� �׽A�ʔ�BEa�.�2�e��%t�.N��;h��hi/[,�h�v1aPz�~�mYtM��t6cϨ�h���Vi]`�#;�%��9�H�B���%��Љ����Yb4ɕ�\�=�u �1U�%�!)Y9k���'�2c(:Ih��v|���"�+LD1E��1�¢G;�޹�}f v�w!�����#�ڑ�K����OYXSv�;9%��U_������%��8�ʷғ��i��{�|Bӈ�~�^V)��#)�Z0p�3�j�h�TG�;@���M7����g?�%�L>���'��͐2��oi?�nCYC�����¤�;q	���1n�{���x�afb���_�" d�˾0�� ��H2�mU��`7Ož�� ��e���-jO��QЎ��>i�]�z�I���z�l��q��Mf�[;I����
�m�2J,�_H��K��� �S��thՏ��U� -���� Õ�e�y���;@U�#/9'7����.�)`�λ^j�_��֣@&�Cl���@m�H�UcăFe�3���d���(�s��9�#<[_�p<���d�R4й��m�������*"ޡ"�
J�z���O�g���J/4�+����gQ�|���$x��}����d� n�^?��+��� (!��Rv��3�S�ҮK{@���}G��G
�5�Ws���!�;�Q3V���#Y�F(O���ݶw��x����,"J8E�vU��3H�ct��ȓ97x>���>��r� ��9M�5�>:�O�J8`�;�]<�g�O(�(�K ���cU����$��2�H~���_V�-�����i�������|RU�q-�jJKarJ��}E1��B`K��
�_��נ���0Cۑ��ZP�sm���W���z�u���=m`+<�ݢ}�)ק��hb"���w��beI��tO��}��������@e��u�fe���31�Mu�e/J�����������'=eU��D�52���t��7y��Y�c�����o�⪃��ŗ��Τ�}�܂�꒽��7�BN������	��i�s�Cj]�+��e���s���,\�;�=�Aiѽ,0�h�@�/bc���Y!�"s���c�K]i}��v���u0�2:wa��Ua~�V�<Ń�d��^���~����o\�����*�����V�Fm�����m#�f��!��+���%to�#�h13��
QD�	���1R���:ƅ��)1}E�$p�Q7-�ĽK�ܱ����D߼�v5d�6�{�kXT����jի@�n���VK�(z���蟗n���� ����|��������ׁS6��8O��{�济qZ�O��`~U'O,'F��=ҍ�?7�����k��ډ�шV�X �� ����l���Ex������'�o=���Л��o'e<j������ȜU2C'�0B����v��=F������U�`Q�\g�R
D'=+KB�n`��G�n�Q$3Mg�,
�Hd��2��͞ P�%Y�a�Sڽ$����=9�Jh 
^a���U/����r ��`]9J~Hф���
�����O�j���x�]�l�М$�����9mu+�W_z��6� W�)C��4���ZT�Z��g�� bx���)��"�}W2��(��6Jx�A�1fr��V4���`��r�Pa�;Sͧ�\KŊ�w�A@)��;��=�n&JO��E�����a��e�i ��Młv���Fo �`��א6��������⺊�_�i�ױ�e`"?�w1%-G�Q�}�� [�&D�w������U[_�x����q-9��V�p���v䡋O��]��i�@�mt�?N
��m-/;����P�F0��z���4,!�pQK�I�1�z]Qh�ca6���� �%P��9�rn���%�@�q���*{�>YT��=��MK�=�����W����V̥k_\[�ok�<� ���)���N��!���`6CZ�b�z�Np(Ǒ�*���//\ek<�R瀕�`���瞫��RNZx
&�j&h��:����\A�NK�4�Fu1�S.��H͡!����	P�uV�.u��l:9�E>�z�>�c���&=�u�Le��ϡ�{ȏWHδ'�3�E��S��G�=�xx���D9Y�r��C�pDw��堍�'`
�n��_����#��a��F�l�E/UM4V]�u��a��������g��+������^b��#�d�����Z�D��b0'���~��@f��%TAc8WD8ȕ���h�U7��@�9�� s
->���?O���[��?��sD����N)�Σ�v�|˲	�stJ��j���:�s{��N��>?MBk�c�	p���q���d�$�0�_ǳ��P�!��C�}�ȱ}
�]z!Gz���&�}yEBBI����BoUS߂�Z�� �l�2�Nb<�]_ǥCV�(�݂o���>]��Qݕ���PwW(IE���cd��?����Ɖ����7�Pϵ�������)�.h�  %t���6O��M%�MV0��l��sC��guC��>[���#�s����-����t�/���H���J��\ߓ�e�R���g��~7ybw&S�'�,=IDr,e�����+��ސ��syz;W�a�}���\7,U�X������R����&]uf�8���LzQ�#�8Ͱ���ݏhT:���� ��^���DLA���0�����fC�{_Wd4�a)B������y��@$�)�,������3�Z���rmO�s"��b�s���R,U�Y�x�`�czMm}�?�2S�,5C/�n2�����^n�[5#�]�B�aS@Z��eP$C=��0c����*+�z����j.�"�LN��-�פV��+yWdWX�����A&jHLO6��%�Mۣ��h��g�pAS��@` U����r֕�_��\"�۽�<-h�l�'v� �ߍb��_!(Oo�0�N+��h������\�U�8�v@ji���AN���f����N���P<���j�?8L�3pɗ�������m��Ɍ>(A�$���X���졲>��0|b�*%�}�k�w�x�"�p�\:�A+�G����h�_�x�tt��*��,:qѴ��3m8a|��7SY�V-�ʲ.'[i�G������zR��4$qG��J���Ӟ��~h�E��Gt<�aR+M;-�ɛ� �5V��	Z��T���<Ϫ�#���DT<e>㷾b)c{��������Q_��k���;3��%�,P6Ш�Qr7�=��MznȢ<X�t�� 3��hU�ą,:G��@���+N�7ĕ�vc��Ҟ��fDۆ11N�$	]�m{�P��jG}]�VZ�p_��D־]�'��im�*x���n�o&od'���|r2����L�e_E{Ƴ�;w��˚�y�a'�2�[ޛ���U�V��g?�C�_�~c�[����5f���t,��
�OB�$DL�Bɝ.+ss�bϟ��9Tc���Rŵ�p�ড়WyG�w������9[ڀ���� ��$=�!�z�h���{h�w�Of}Y/�ު08U$V_�;��K��k��fw��p�z:N0%�l5"�L�:_��
% 	9��{�lt��X��dqd���A3ɏ=(牨���hX*� �������d !������m�^��ӲV0��v�pc�i\�G�ټ�$�l��s����1'"���q�yX�q��!*<�p��2��4�s��)5<�(�8�M�U�|��|��C�6&���3.��%�c�,�e���F���@��i ���Um�OO���懶�ļ=޷QV�D-5�e�n<A����B{��-	3gc��6ɤf�\[���?A^�å���~�A�^�%VBR��[XBP�ǵ���l[D$
�^���@K8Q���m\l5���`���7"�����`�v��wW�"���g�}���Q�gT":�]�SM}�æ��i��@����;?JC�����tufe�͌]�T��z��T�07ޤ�ƈ����MW����������A�$����o�H"r��=�����F����iq��]�q�&LY/+�����~8*�k�j�rE30��I�����6���P�˳�0�%��������]0��|�昁�q�f�|�WX>%Kt�.�m�|l0�tEj_!��`_�%L{r�u�����t1K��6��U�9��v�8G�u��"[NS+� ��O�澄�Ns��so�Yr~�u�rސo�w@0���=�KL'#��nC����-ʛ&9b��������,X9�|��c^��#�#��2ht�*"�j834L�V�Ng�?s�V�Y����6S��tO�L$��=���4ڴ-�1e4�s5$�"��!	�CZ�C=���e!��d�ȿ��	VJ�qV�"ex/'��z^�h�#�3e��]��4�/k�0r��ODO�0����j��i��w7+�OV�z���y�`��X���z�����%�H�PҀ�gЫ��\����wK���\pIe5��`ńğ;��@i�!��ؠL�}��P'DV�}O/�����!�qWs��9��+#x`(i��1��l~�7������F��LLcM�T�kdi��B�L����<�&L���k�+P���+�9��^�Ÿ �ǜ�#M��	t����	aZ�d�q25� V��fw�(ҕ�J���B��Y�)�og^��5FD"�Q��E�F��:�-�u�k�cjGu`f�n�&���~�W�� LE�KF�ZK��VI߂l��fS��ܪ�1�2�gga� �n5AX���ˇT.�ROH�	�N��D�ֻD4̨���L�{u�D���I�T�̺O\@ol/fS������=	i��n�Ͽ�"��TA���]�\W��;��D�i�Į���s��n__��W)��(�:j����p�/d/����ScV�3�����8d;]k�d
�G-��#�Ά����zp�n},tYik"X���
�;��J��ԝv	#%_��0���^E�A�+�Zbs�@D��"�ًW���]M��BӛAa���Js�LY�n?�5�H�C��QV�1py�i���5����Td���D����4p�_D��x�t����;|�9�W��t�LbKƈ������� �^q}�ɇ�Sਥ�]�X|�5�z��k�
M0sEz�P�'�2� O�O�g���4&1��֕�{�/KYh��貎�L�T�@�B��eRȳV�?�db	GE�f]W�\�,���!�F ��>�P������!E�H�m#9[T��88d�g�	j���՘�4�u��+'�@�)��j*���zB��)�ԾH�0�D,M��
����#�:؍K���R�dA�d�L�z�Af�fX�����@�@�~���ܗ�9���Ò[����2��P�gBfO�#24��+uV�b�=h�eߙ���a�(�gp�H���C�����_�b�,��a*c>�)A8&5l�~�T�O�?@��ZZׂ��5��F��@��P�eM�U�!��@�:K��V����(���yǳ�F0G0�.�rȢfpm�U�@��\A@����hf��θLK𔞉t;}i>��fF�JP���9*��W R!۔*W�S�ATB�ʚ�F�1��"]䪚R�j�+�BAs� ����=7�+-X��0�8��
,��ꏾS�o�"���q�����x�	���&�W�ác�w|aq���"������9��[��;�4fX㐦�Ô�s����=�E@�o%�������f�!O�i��ڽ��X���=`�):;bYE'�L��(�	c��.���I<KG´��׎�2i����,6���>*�?�c&�baK����Sͯ:�RM���ώ�2ͽǷL�ˌ,�������/S���n�9�����c��m�x��9�ԗ�����/�L�!�y�c�X����('d�'
��j2������0?���i:�hC:�l�es�n���]��'1��Z�Mb �Æ&��')G���ͱT���F�鮨w�R�������ڡ�(�P�R� σk_�K w�)��
�Ar�)?�L魏X"b��Rx۝g�[����X�,
�>Q,J�D�򼈞s.��$0�dAiT��@�'=��?��r&�����_��f��͌pGO�ca���ĕ%�B1]F$gz��/�����.Y"��ؘ��}�"�������끗��q�޶��U�j�":e�t�W~貕`�ϚE�ktx��\��b{ԣ� y!�̵u�����꿟�/��'/��U*��ϳdlD�x��@L&�;F~%`��:LD�|���~	�d�Q�>W'wп�/P(om,7�X��}��y����~�U.��dѯ���1��խE(��X�77�n���+t�f�@Jx��#��͠
m��!Z�O!+�È{]B���P^���lү-��Q8eȹ����zfӶh!˭�#��ܣ��R��i�	�WC 	�锣g7�ny���LͯQ�#Qu��NJˀ��H���̪:�/���ٹ���O�u��ds-�;(3�⛏�"��ѯ_���)�sx��C$���T��.�z��C+|fsқI�_���mϭ*�|�āl솱��.�J-r��� ^��Ql�
�i�0|�n���5��YC�m� �ĩ�J%)����<�1��Z���?%��
+%�l�����@������®�dޝUݣ�F�d��OJ��!m�0s����:�N��BAL���8Psq>�!ò<�,���[��S��j*���h+I0����8	4*�M8�-y��:�;�[���R�δ�}1�Đc@�/��M?��ᔪo,�m>�>����vz�2;jw�vd?����X�e��hϏxO��J �=���W���3����|5�����R�D�WGuF�Rѫ�Au"4B���0�W�=�Q6�!�C<H��<_BlU�r�ۧ;����&&�DK� z�R�u� P9��Kt�8�H~Z�Ms
�ve6���VB���x�$7-��\{-3�'�{IJ�.���y$��!4w�v�FW���SY��}|�a� V���\~��W/I�H-���:L
O�A�g.���l�$ϲ���X �|�6��/[�F"����K5ܱ�>� #�e��b`�L���\�('�H��~�z<�#�X�j��0(8T74!��V�ZH_�FM1}۬��ک��i}#�W{�Ij��	ss���z﹛��6 &;��Gg`�Q��������H���\PI1�#��'/��@,(��
\݌ͮG*��|皝z2v#��D̴�y���8����r�$s�O����S�1�+��Hm��>�د�|S��Oڦ����"��޴�w8�����\W��$ow�ɐ׀@��4Bl�0i��=��"f 5�F%����� �X�G�����~4i5�z�%�_��]ȡ �Aw'�7��n�0��8��.
�C<���S)x; � �CN �v���~(xG ����7>�}nh$����#͈I�z8�$}�Ƨ�T9e�^��E;c��ְ�z`FVݹ�Ea�64�֔Ey�h�/�n�^�_��ʰ�'Mm,������$�]o�4��q�7!��/���R6�Ht����
�\ ==|�,�O��Q�ȳiN�ZB˝�kgl�{�rE���&�ћ}��a�)u�І�TH#����c�L#(=ŠA32"���L�Z�{�A����f��y�c��1��R`YV��i̩NuQ��,HQ =?�0�preG7	f���H������^2}�.�H8a#�.�!K���%t��I�b5Lo���u�]IY�G�u�`���W�L�S��&�����	�_2r���\g�m�,'E��X�z@}��z�[�Ž"Ir|�v�UT�D� �DX[:�7b�M� �˛�s����&�ER2k���'�*T{�Q� �"\��Z)�4`I�`����舺`"G�<K�j塙�W��vLN=ϰ�̱m�����8��1Ԝ����O)as-K�V�b)Tu �}|4�[�'��|����.sl���O����c�8��
���H��V��ieNƬ|eJT^��*If���*pL>���AP��;��K\�~�ϵ��A���߶�[;sB @ip�,�L?a�!��|D#�R��=��N��"�4ZW8�I�k��G����e	I�D@}����K_�O�m�"C����&�"@�!]��
���I�����Z]f3��6��ȍQw�c6��#�N� ��5#�.��[�vlN��I��F]͢����]X!i�7"�^��x����a/MEX�����C���;Źq7k��X���{0^������W=��(����@���|�`L��K�R�:t(�>F�bk��l���έ���u^�͝*3�ekrT��9R�N��G��±�d.�3gE��x	A[k(���Ob�Ur�t�/���I�_��X�,�ǒ�
؈[iLk��U�>T��'.��߆-Q��
���g^j����	8מ(J�Cz젎�M�X�E$	a���3��˝�fԈwV��~�f8��>d�s��e���.su�tp�K�-(���~�+�����X������u<�`�βB���4Ţj'݊T�#皪 "L�rK�k:��R�-������Uww,��$T�[Vv+az�-�S�<�R���@�������pd�%�q%��D )�q&*�4�;�x��BZǬx���BkW�t�8l��b>՘�]{g��Y��vf2�_sR��b��bZ��׮�ټ��q�{�6��e�L ,�N�#�J��p	N�B���S��u�^(�wn��X���/>:�U~O��-����)��l���􈲞�դ4�e�/�q�������#��a�⑵㫏�U	��/X)�G�U3��������)^ӽ�r�b#3G{ڷF~�ά�b���$"g��IgX�Fx@GT��ௐ0��=R#���[<�V�.f�f���ޭ��8[���m�;�3٘
���6p�Ӯg����y�,/u���e����{�[IM	C��>���5	�\�+�օ�30>������Ơ���#2[z����B�o�bGyx�P�+�Or��J�u��3|Y�5bHG�GYauX3��j�Е�#J�q�J���1��D	�������6��N��0.�5���$��ı|>gi�v~j��?���t�bE�����GM���	�՘M�+��Nu$��A��hR倍�Kቦ&|:84�3;`��R��C�=*S��،��(]{�ز�X��cW�X�Xf�sWλ?��Zl`���>����Tl̻��P�6�@:�D�����g�D/ߠQ��d����������VO^�&5��"�wL�M�	ɛ����1�N��ȥ{�W��(�y��=�;!`�!@bg�������zY���J?/��LJ��4���ԗ����=S��F��ʲ�W?�f�yHIZ0��M��d'g�<�<�J5	.���0VQ�}�����	l^tQ��^�e_`������T�A���r���,�B��S�b��z&�W��u�÷�0U�5)d���8�ּ���3a��sV�,�������vy:cHQ�ȋ��[>2��]�����KV���G���!ίPģ�h�I/" h���5V	��bŕ�Ë;�"�3�o
O���߭�T��]��&B�~�IP~��!弫�T�Ǫg�*>6I�GV�f݄���g��)�告���0}��%O�}0S�{y�7��|0�Q�Ֆ;6֘��vM���WF��7 �q�9��2[P�g=F�b��6<%�0�'FbO\���o�l �MW�מ�y*�jG�vR���5{]��o�b��"a�t��Ƥ�f��T�	�=-�)I�?e�=|�qt�i&�&�_�_XmX�	jA�";U+eE+'i�~�̿���D�����@�!�e�W�8��8绔��-(n���b��q�r1�1l���#� ݄�ߊ�1�d��LR'��I���!ᝒ{����ND�@�ګ���rd�����py��E�����N�o�wO�o�e�}:js���ݾW�!��Lo;g9!z�[$���<1qp�s�e �F2:|�������ۧy�[^�-��؍k|����E�~{�T�˼N�w��_�mc�)1��$���"f@c?K������&�8Ç�����@n����GR��j^��d��>�XEd ��q���Pzm�FI54[���/f��y�# ��rw�0.<�8PQ�%r�:-�G���{�c��GP_n#8�#�d1��~�ซ��H��*�-�� �R��E ��	��ZN��UnEa�uGzހ//��U6���<q�i%��z�#�?B��B�%����(d�\�s���=��J|7,����S�9O��U����4桋�������#/���N��l2��B7�_�ȩ��sX�  ������Gn���Ѕ��N��һ����Qd�>k�^V�W���\�Ps��qMPÑ�np�nS�M�=���B'���ࡷ��peQ�(���K�}��4u��Y�ut�;��&Z�&'ԍ�R�����C�o�MK�sT�G|.��c;h���w�b�/�=��v����i���Iw2q�������d��;��C��*���0����_0���j�~Nq�%��Y��E��\���#Vq����
�ǐajQz�=�B?�=�"�~@�&P�
`j�v�̂_T�D��h9��$���C��l5�65�}�D����8?��xт
���L�{�&��M���L�{C|�@����� ����p���I:�N�������������� ׁ��\�Ƣ�_����[e)���ۗ\�O~i?M�%%EaE�`��'�r�$X>ﻻI$��0���1�2N8���R��������T`�
OA-�/�1�*�$�Q#���8ݬr���}�WK��t�;=�o���2o�3�|�b��̲��dr�Jxf�>@���*�Ŏ
���\��6�T�[��e�3���ū{uAaH2,.�ڭ�owZ8l�vg1������1q�j�u�d����Ϫ"�������)k��"N���4QЇ�e�Hx�˵����vD�{Ս.���ml����*���<�B�c�{��H��I-,T��'���v�M=J�,L�#5�j�ꣴY:ƌp����u��}?zK����B��΀t��ml�]����"��oq� �<&���);򤎔����)�� N	�}y�W��4v�zK��=V�#$���z�U�Nã �>�t�!},�*>ư�]�� ʲ��%�����P��:��A���_Wgܿ���FП����* ���?�R��S��r|��E��j�IPw�K"4�ϧ�z�]��IIc����R#6��ೆ����)�1����>�p*�� �ZF<w�9�9}#��@�.i��L�<u[9qQo�&J�8�P���B�Ҷ����J�����h�����K�DC-)�
�R��z�K`���fZg%Юc�%�kηZ����#�wci0[R��0����k�_6Fv�t�.P�P0�.���T��FY͹�蕳�nV�&�s��ue$?�] f�	*8��i�8��#&�N��O�pK���u�Z�Ѩ?\�n�v��+����^�	��~JP�]�]{`��5�,��{�b�j���K��+�e�Oq���W����C�q���#�6��Q�gu
�Z۶ߐ�~6����?���1��I�x}�&� i�u�?�	�,�s����RX��W���K�U�l�Y]{���Wr߶7O6�v/�rQ{?�KD?�#�Г���J.z�f���/���޶���A]��i�C
|y �y���44M���a`
sM(i�Z���zm�"�r���xEf�V����#��T���	x�d?����\:7!X-c]2@)��l�;���7E\���	�Z��Gbp�vY"�;��o���P�_��p���=�U�[N+[�X߉\�&1��dd@$����R�hګ
�p��4jCF�R��N���a`
�k�g��&׫�饠aR�9�y��� �5 {�c��o$��̤@Q
�@��m��ج��B��Z����H9��x	�-�+�����4kp��FvL+��%WѦ�:p�4���֒ 䴴af[<��!�q�K�ؿ�b#��Z�Dx'�7�]AK�
ط��uKz�ڃڮ���.�0E2ď�A�����	��̱;)9�vɧY�Ƒ��a��Z%k4=��#�P��������Aѩg����Cچt�wy�X�8��i՜5�@��s@��T'�^(���[�/6S�&��E���GS�d�@���?�Bm�k)T�v!�V)��KX5C��&t�1�RhS!����T@S8�ZW��/m\������>�c�g��	��^כ�J��4�m��iE�ez�!'_��P[����gEטzL5N4}��/��ް��I�CK�5M҂����w�bw����d�EE�U�$�q2�8S��d�m.uGBE�tf��Wj��ϻN�xcR���� �1MI��sU����O�.	;'�'$��U�Z�F�����lnY;k55��קp5��>+EE Р�
�.rT�u��`�l�����9,I�8'��ga�2�N9\�{��JE��Š?�'y��y|�t��D�*h=4�[oh�]G��\	jĽ��M !|�Y���i v����WW��,c5�	��m�aa�-t��D�%Y�����a��#"����H��A�2z;��8�Yw�hȄj�yd*�8Q/r���I,檋�	zĲ�����e�w�2��;1��E�%���z�W��\�X���qԍ2T������Ģ}�^��]�9d-���A>�bzd[�~p��%L��x���:ꖘ�8����Gm�M>��^;�iQB������M�ڶ�#
��mخ��h�
��ȥ�Kwa�lܯ�xa�'�&�Nnb��$C���R.�a9;BFD�eӯ�Hz���@'C?�J% ��a� �x+�������H9V�kG�L�����zehvNeq 
��Z�\:+��k-/H���Z�VG��Ka<W(���8��ETG �4��w�fr/���VU&�m�󳮝������y^�c2���HYK�6LB�=~��u�^�Ǳ�+�Lv��P?���ˀ�c������%���1|g�Ι'md�.�a�|�	�c�K�7g�w��OiIm��&ӳ�NyH�
�g?�q��T����`y���X�xx���DL��~1쥌m��ODQz|vV�Ng�R �����-��l�7�@}Ɗ�le�?dq#��������Dj�	��DH���@��/�g�K��6�Ş��2G
��I �����%�eh?R���0�T�Pş� \�oE�1�@�H^�S��b!&�!�K/�I�E �v�(tq4v���i�i�M�8�hL=2��R��/}�,�keU#�O�D��x(��,R��Z�5�}!����c��`�b6�S".���r��~(�{k	<�p iK?Hu��Z���)v�^e�t�[�}�w╀o��ġ /g� r"�%Y�5WÛt��.���#5l�z�Sn���iS��éZ5�Ю��X��(���e,к�X�'fzeﰈ�\W�s���e��|8;��,_d9`��V��3��z7Xy��*�CZ�hF�[��̨3��3�x2����X2s8�|��v]��ڨ�BP[S���ܗ�Q �8aI@��ۓ[��e�3#ԣ��n�hS�AKu!��M���)���P�>w��/sP���%痦,�'~ٻ-V�h2���E#
Gz�y��?ՠ*7i��3��_ك]"ڸ�F�y������:Q�!#���q�����y^�@*���ׁ5�)�����M�۝Ϳ��ҳ������Lv�� ���l�~n�֑A
��\M���-R,�r���)�}\�q�����/�oM{��Η��������6OG����V�8-w�1\>�-T��Q濙{��["+)�#�e�9��p���D7�@$��Qi�AK��y+k���$^��#)�J�ſ����h�x\��(Eu�I	ZN)�b��?���f�5笱(���WC�Ǉ��������=x�2�b�@W�/���.V�S�ެrM~a��5^J��7�=(����]��Q	'|���܊��=�,�YA���heg#I1m|��K�����f�m�HG�hm�AP¥��A4�L�#�~�ƵB����gA���4�0d��a�&o�,s�>s��"�X苇�a^)UW�"���S�|I�B���'�k�P#�����	~�T��(�P�-r��Z)�]���k�����6�-y�E�>��1�ڎ��S[���]
:�1//�z�#�L�e�Ί�D���If'���	`�,�L��ӷ�K�ڦ������W�,�r�-;ڇ8��`IͲ[V|���$��^ ͗��ŧL�Q�4=+�27\P�̷l�(���m�ď?C��P;��oɚ��D�xl�A�~KweW%��WB^��z��&�谴����������n�^�I�;���Z_���+��M�b�07ʣ��Չ쎒�kUe�������5��6��)�E�Dņ!4L�b��٫T�*"xF<�\�a����0r�Bc�lmz�^���:�zg�� �	2dz�H�ǝ���<�4^7%�����@��(o%	se(�ss����X��Gԉh���G���T�z�T�L\sv�xo��=^�E�1`7��CQN���ވf�b���(Pm���LzZer1PA�]�����wj�w��T]�w&8��#�Y!��G+f��j+�h�k��d�k�e�[ŋ`i��%����G�8t���/�h8N�ע2�=��U��l�C��	� TF=�uk��x�P��]*A�L������(�t�c��Z|ﱥ؉Aǳ��=���sq3�e���a�E���ݛ6O�f�u���>�-���k�d�_�Ȣ�b��_S�sH{�F��z�����`�p'�vkI{YJ��=#*�36϶���t �����.����4i6d��ň?N�w_iM��.V���O�6��Z�Y�d;v^*��S�z��E�æ#I��>CH��$���J�:�Aǝ�z��aH�%�ЉmprT���ǠJ���W�%��W���� $d��aX{���9���APUqq�>FTԲ��%�#DL�����%j�ל����ӹ�8�o�����Z>V�l����,^��K~�]�h����9h���z����t�&��NK�}�U�4�:B[@��w���>�m���o|�:�|�!��h��[�T+~�?�^){^��҅�N�\��O��9ty���Zmy�>B�Xg�lX*a��8p�"��]�hx�ַM�XҶ�V��*e�%��GOF�*R�e����s�?`�;?�2]ṎQM��Ŷsarŧ/{R��+�4G~���О(;&���:"4�1�fr�gqhU���^n1O*{�%���z��O���)�P���d�H�U� �҇5f:��r[W�[�rX\F��0�jDI'��pl�ԧU���O�G�{@����*��V��ۇ&uz�)���DE���|�;���O�NN�/`B^�~�)���,�4���P?�-��os��=�r���t��Q� �5i8�M�����b�SR�o� ���a��� C-�����²(9(��2R)v�W�Pk|J���ȏ�/�_5�:�W�ӳa�<�����q�rS�^g)���{�GW[ď-A
\�ʐr�򔵹����h���!7��ل��x8Չ�7@�|������$Wy���bPv��9�m�s�a�Fl�+�o<3�'/���5��0�"���.�\����A"�S�8#�=�i�p.�6��!짦\�����K�g���%a����������6�	��@e[�YB�r��FP
P>(�+��T���)�ո*�����U�
���Й[z��:�r����n�VM6ge�-"y���S�/<B9)3ʇ�b{�Ί������N�e�Zk��8����xN�G�p�+�;|bf��O;���䵮[x�6�n��Ϻ2})J�A�Q�h�Ȍ�L���`��0���i`����<��:�y�~	�<j$E��-8v|x+v���)��I�P]� ��Q^5�*{�:/��p@��axKP����pq1SG��_*��6����X���[��0��4�����Eo��}�L�R�f��59Q��"��L�iE�o1#ݾͶu jN��h�����]���]y���1-�G�#�6�����I�׊�%�����ʃ���BJ���w�K@g��\j�>���X#��1]�Y���.����q�C��eՖ6�~���,��c�M�c��3�Gc�5����6�1雭Ko�D�t+�zK[�����O�+�R[+�A����1�U<&���-��K8 ���b_<��g��c6�K��#�:���z_�	/*�y����j�2퐰��Py���x2�[`%��Ho5�b�?M#ɣG�o�����{N�3k��|�������l2�5�禰Bd��:��h��޿����{&f%:�����+�l���hY�`9��_���w��|�5�k���}� �CBG�u�my��$esx�bĭ��f4J���C�]�B��5U��85�Kt 0�mzw��_��V�m�(qr6��
͕���|�%^ �.W�ïZ�;����_�{���2,�R�j�丂d��2�M���U��_)��8���6��ΓeP�M��I��ʏ�R��=_e�����sL������]��d�ۣHR�2mK���
��}0�YݳkHN�m��6�I`,�U+�X1m%�N��e�Z*����
װ�N&��m*��m���9}BV�����?�ՓuA���'��Sq��Q ��1)ޟ�J��i��5h��ؑB�UMw���(û�?�����g� cE�ڭj3�m�g��H�� �gbW8YR)8�F~��iȬ����r���\��҆إ����b�AZ�
�u����7�|�M{�s`��_ߤ�o����վ�AX�l��gw�)�n�v��$,Ƞ�7��#��\�5��P}\Ѝ���-J� �w���
<u���aU�%>՘�s�)�����&
�3h9� uE��o�N�u�U��p��|����+�x��/�F��H(�w�eã�i�w���Ӿ���n@o��{4�0c!�} P�"ua3c,-˟^�$�I�3?x��JM*��;��IO�ΰ9�o`���׌�����h���d���Y�գ���M���CS�����!z�=.�K�h;ۄX5�A�=;���VS�fϭ���[>zy�`LAn�h��ǈ��V�˒.c�m��v�����"�b��K�b(���2���~�Ė�O<���˸��+�M:����󋩘�a���?)�\���ToA�J���`M�d!xK�6	��n�c��LC��'�S������[/Y)����rZ]�B��W.�6`��܅�TR\��ԝ;���C�/\��+��l:�^�0�_!�P�gF�g������e|�v�:�04�&�IN�^�k���{�Hl�?� �J/����T�UuCbcF����㐐�!�)�t#;��5?�P����
qg|ke�f̤�;K̭O�̝��v�lA�4�G��CŦM~+։F�d�˧H*��"��A�Ĺ8Y��3�w�����*�kg�C�>���Q�X#P:\�\��n���7�h�c���I��UkIpUu!�y�ꨣ<f��Qo,�g[8��·Jk���h��"��˻��}=�E�G��&|:�>���R+9mHr�K@,�w��6av�q��hUC]�۹��������m��N*\�#
S.�|���{��P`�77�T B�a�m*G$͌��+Mⓩ<���\������2���6��pbk�8�qE���{�ö���������+��.���>ae�k�zw�'�w`']���Y%	x� $��pˡC�۞��	��DU=f_�AJ�5N���\@X�k=�qz�9��0	D���
Ĵ�����j�\i0�
�:�F"�(ϭN�*�7�n�A)�� 1ʖ8���@��v	��z��lEƿ2Vw=l�n�{����Z�����$���lFըM$��l*@���Z��Zc"�7xjNi4�����o�,��ȸ�I�3�~fQ�}���+�M��؝:��$��)�t!L��9�)�R ��������yO�!�Q�)
��_ff���w���@�6� ���wq�WIO�u������i�=)�BI�[�q-#�ŗ�ϯq�I!ZX��[��}�p�w�'F��Ǌiм#L���%Eth�&��q��	FM����:">pzx
��N�C
�w����-C�`r�]`�V��	�E @��,�#��a���R5��p�������g(d���`���)�/��h�_�o��=�~F��܂آ+e�a��%�[^I�R�1	�چ2}Q���/�%�ù !�;K�U~�#  ��K;�����"4Nԓ`l��~���s���u�o��>�0 h���h�H�!W�cQ�Y��;�q-.�~����{ާ����idOڍ�Q(#(h���[fI�}˅w����ڧ2OS��2��!�7@=��%����M�4<��C�%t~�L��9-����21���0s�X�*���i&K��ŹL�/���-EsV5f&�z�,7ܧݠ:�)�Hd�׳�>, k�oR�>�(3��1��Q�I��# ��Ü�e�G�Sߖ�Rl�)�|�ު6b�ۙ���?,ɐ�ͼ��� ��r2Ϭ��j�/G�K�֛�0Ƌ�Yv]�9�Ͳ�\�����]�cC=�&���Hb�?ىY�a��r#�ل�����)�]���c�cw�ܝwR5����1	�e$a(�(���"�f��;}E`|���@�#0M�~�d	k��!Y�mo�q��a3�{��C
�����f���Rq���q�K����S&�y��ن�܋�:�W��&�Q�γ�u3k�-�KV0P��1��m��حG%����FE:B�@��)�<���뵆��2��n���$�=5d�g��f�DN�4@���x����~�_mW��ꝝA�FF�Áv���J��nÀ��/~fU�dEw�{6:�^;e�I�:��s%{������g������dƦk�Ad��m� �31�(���dZ�82�[�n��]ƹ� @xC3���f�*;�Dⳉ��P������3�$��C��z���ksp<�d] ������&�}��ȸtT5��㉸av7!�k��"����Zm����W�9�s,�u%>��3ò	�v(�rE4���Ty�Lݘ}@��K���?˙�̵pc}�u�V��b��)��,T}"�F7�\�k�2���숂GK��_x�\�K?��`R(���4�-�� �l�{�g���B��JAׅ����Q����D!s=�:��޷5�y��l[k.W�`Դa���?���a��2�o���y������0%�m�(p@=b	]�,��M/��`=�V����9��=�`�7�*�"�0��ٸZ@9-��}�\�"����Q��<��b�-�DHN$�P�2�H��oe����>^*/K����}{��3d�n�i�g�"峦�~�c�1ܻ�ߐ(w%��-_��傥7����s^���`t��e�խ����{ t�T�*�!�e�7w�4��i_{dJҸ�(E�aL�%�U=�]0�&�y���c�\��·@��_���ozy!�UrQ�D(2²�i���
S׿�6���=:��3]��*q���d��E�`�ff����ix���h-���cx�r�5��'bUC�@��oU+h'M���6�ܙ�͂��<����� ��CkY�~%��:�(Y
;;l��[���Z����*Z�7f8�;1�^�����N�u���<mP��]w^�#r{7�ݸ�A=𙙹�E����M��#�*�x�w*]`@����9��o�x������6eZ�R��zԌc��t�ڜm븏�!�X釣�N��6ók�'ֱS��2;�/�e��Z�F����ׁj~|B�ǁ�_� ��s_c�FK�B�(\��y��Q"c�_YR�����7l#X%E	
$P��̝��xjݮ���>B��	q���P����Li�*=đv<Ӗ�"��=WY`�/i �C7V��D:�����+r:$؝��\��]?�A��[�]z��	 /߲u���J\�@9K�A͌3�XY�yMS�w6Y�u������zk-1\���;(fh��H&�f𞁱n�CC�/�c����\V� ��`��`�1"h�l#��5d�$�|@�&!fP�mt��޽����+�����\Ep#���E��� ��p�w��[<N>Cw,f��D��W�@�+9A�Q�W�����V'��c/!�v�[�O��K���g���'��c_��F������B�Ŝ��P�k��eO>��%I�� ��=5~��&_Ӭ/������.�e��ZȨ����\�W ��^��w���FI��3QtK�<��G��0ft|>��-/->�9c�\��)k�/�z�{+��8��!}���=\ʘ���։H���D*�bݥw�K���M8��l���PRO�buu�W�ݯ������������Q��#�Y]l�F���ֺE��������� ;;����3����9w��;���,��?�����ᐜ�ƅ��МhhL���Lݖ��^V>:���T��v���=̻	���Xez�q�}� �����r�~���$�/�Q�q������� �M�� C�>[�^ �n�!����ts`~y"R���� 1߁��qF뚖�2_t�E��N;\k:��,2}��>İQmPE5����O�Z>��qZOJB(2a�Y�nSF͖|��������!�j�'k&l%�݂YC���rb>� �L����3��r6��!%�ͨŅ���u������dWq����C���A���/���z��ޢS<��������j	\�Dl���U��)s˳3��U�do��
��~�8g�:���[�?)+5�,�hk>EC�ip�0����E�b,[�,�?�X7s�!M��������4.�V���qm�H�>έ������νn?2��u\�ʔ@�1��w%��
(�6W4T���{��?�g�kG�������<�Odg4x��|���y�z*���|�Ӽ��qJJ{�ʲ���K�j\	lyU6dP.O#b�sڪ &⮗��
��{E'"|4�~B!�}ل��8��2�E�����̢V�������w>��V�wh�:!�rP��	`�?w%wW7�ǗU����߃hF����o��.�[Q��X�R���� ��v
vYG#�}�"=�Z��2L�t=l�ކ��4��6�~;�aU"�����Ym�U���D�8L�`�G�y�L�xԍ�N��hnG.�
j���̽�A����iU3�\�U�Sh�T
G��tF��~�%�,&fS����{�0�6^mF���F���?��>w����s�A9O����^���x�o��H�,1Z:�0�$ :hx���cY����P0���=`=_�K��r99�>LA�=�:�l.�Y%��٩0q�	Ӊ��i�݋�mZ�SN����h���r|Q<L�X��>&K��YPJ�^k��~u�W`C) 3�q.���w���9���D�%w��d�UN	2�b�������Ċ��$���B)��%q����Q�6Ma��"K.���<�W ]��)c�=փ0����-oV&�|qM����T'	s=�R������?��\�����|�L����sR)��)��#&$�{m8�W�ٗ0r�!�ʿ���~�<EyB�Fn�� ����C��]�?|XH6�ｶ�9����	�W�|,�xOэ"a�o���d�z��c�'>��ĳ���𖗍�}24��1�-/8̿K���h�{���Zi��|�p��ߴ8��	���s� Pt��W Xd�����v����9�M��Q��Z�C L���q�}�J�$�X�9;���d0�Գ %�C�g�!�m2DCWc�� �e�0'�*`Ƽ6���hΚ�����n� L��=}a�-�v ���XF'��Po�B	��V@(�9H� g�'8��%2�U��Ρ��{�SS�4�B��Cuh�Y�g�����A:���8� �@�.�1�_�Sf�S� G"8��I�BF�"��|	�e�r�en�F�7��{S�.ֆ�H5і���&�S>�N]�/ǎ��ʴ*�����t��e� I[�Y<L�'���6.4�1�j)�S��Jg��婋��>�*%���\��v;�%�mln��Qz�&\�Ft�B�����}m(�����}<��>W�P�����W~E�]���v`�c�P�h�@�J���+ݓ �*��2�PE
5�_oF� �Z�k+��7;Y�tj��ohZ�� �������&��R�k�ʉ��ru�a�9��[W��I�}��7�2��g+ʑ�>	�Ak��y��	O@��*���V��'���oT��A_�A�E�b�f����ќ�w�d3���~HH��^6�\���S&�|C��5J�#gt����Kl�<�����2���z�']*�bƚ2���f"�#,s!�i�B���׽����\-���>��:V�ޞ$/�e�pY����Q[@߶1���yC�p�����X'�*{93$U�̉Р��ω�%�����q����P��.I�:/cx�T\+`�gVoN0-���N���̯I�P�J�8����F��=��S���l@���]�J��ʋ�����D!����i�6����u{L��*s^� u0�j��Ɇ������}��=ķ�N��^��8�T`��Y���� ���b� $��*f�G��՞�*���qqJ��$$��������QY~y��̻�M�HG.aB������P��^�NQjI����U��jڙY������f���EI{�n��xc_�*,�:�Q��]����#ݡ�H����W��O��� cp��&)���^7 ����@��"ɸq뜼����o3�|������]&������u���{BwJj`����g��Z������`�
Y&�<�E�x���j('�7�u/����U+�wR��_ ���r��c�Y�K���c�_(1���|�5:�#�*��έ�����Ǹ�*U�8 H�<v�7hM���+��K���V���H՝�tᔚEh��N �I&����F����k�k�c�X{��R��Dl���ʖ�m����q�@T2�	��bF���-s�9�6j��6�"��}���W ��7�m���y����>m �<���*�	̗�?�$��|�ܢ�+� �B�jnMB���H����}��B��$�!���cؼ��#r	��s
�����Nw�Nm�O~�_V�juNꁯ����VA6� �x=.ì�R��Z��)~H�xaT�f��"\���R���#�����i6��5t
�*_�����u�
�vA���s2 R���!!�ڲ&I���J,J�B��tV��`���r,�Ӂvz�Z�Ոj7�1�и�f� h͆���i/'U_���%eRi�/��DK7��t��8-��1;��V�8�8 ���3l[;���2w�ч�Dd�ִ��1sN��V<�����ɞ��>*��9 �I.��s��G��_��g��wB���UKb'"�jD��kk$�B�H��2��0�>�(j����f~�,lb�>�b�lR�Q����L��-�/�����F���^��&g���L�e�[��5������7���>@�gG��SՕ�e�r/鬟p�d7m9JG��a{�1٦��Ǳ���!=�1����>ep3�� }-��s�5mޑ$����@��2��}�z�s�W������iՖјF�-����S�����I��a51`���_��yf������_���>��A.YWJ:\�L��q��e���$�@HK N�~!R�߉&�<:3b�fEaoU�������<:�a��'?�Y�,�#����61u^��r[�$g�G��W�+2����5*�$�1�q��/���a%�\2̓����+(}��u��b���t��[J�Ȭ��>�n<A5/oI�G �9�f����/g��4��P]W��j��S{ϋ�k�qR�v��z8��\�?�&k��%W�b�����룚JyӐ��&a��d��B�\5'��SM9�8�H��]�n�%�(N��6������9 E���^bb�����͗M-���F� � �������)�в�d��t�D��$�O�f���;�;+�]M��O�������\k!JZ����!�_���U��&	05��@��w�/�Kȷ�]Q�r]��]���Z�Ԓ�ٵO��Bڥ����z^0��:,��w���=�J�L"�ZQv7��i�^�Y�ܚ��p[��)#f�!��zO��ͧ�g�Z��-��3f��'"ē��Ok�&鷘��mJ�t��%����f5�UIQd���=�(	�����W���=5�-%0`�<a���>�D}E?!�����B����HB(x����`ĪB�LWv�F�au�u~P�"\u�����2�sg�2�w�v�IC�Z:�,2�� �D�,ɼ�n�j� <�v'������#�H��M��v ��P�f������+���+Y���o&hMn�l�B�o@�/ל0B�3�0�)�;B۳a�x���O�������G^l"߲�m,RG�9�o��B�q��|�ɚˤ'K�L��*����;)�x�k����"Yq����,�x���K�!z^s��BHlu|� 띩4oGא1����m;������q,-f��ܚ�h)�Pߔ���Y�̍�Kc�!�9�[X����U8��}��1D3��_��a���h�� ۠ф��K3O���f�?l���E��#����QЬ_E>̘g(`�5����+T�7��Ԅ.��_���Ct��S䗚�,"��0�XM<���2uy��(���$8����3˛k�aǐ�����
� �_@���gm9`SY �&+��&q�\��ߛ���3��dI�t�$��0�������z�n�1��2 � �2��D��$�G7~Y��PϿ9��y���䞂�w@(�9Z�����h�����F�E��c��$��� y�ź��9�ID�ox����j��V2y��:�{J�z=p7T4���ϓa��|�C�c�
�I�{�,	����k�����`��3"Yw��w��4���i��O^tbz;�f����x��V�Vu/�~
)�陥�6O�&&#��Ð��N�Âk�>ӈO&��ð�j���u^qR\��!���gL��~+�R�F0�':�e�og0�(�߆U����F)�*;�O�Y1�&"4Lbs�~A+V��H�I?'��p��&gg��=��!����L �u�}|)*�Jw_�Qe�QL�^(rP_�7�`i�{Er���(�}6Ԫ"\_j��E�V��8A�A[hEу��o��y�Rj_	�7du�3�xc�{���&Q���y���c�I��UU��+�\
-��f!�V<%�1�\��[�����rD�Xmr����P���~FjoRd�@����T�:[��*��
|�	*�&�$����H5�(:o�1GN�AN�	4�C�)p�����8�����h����3��߼D��JȈ���e)��B��@b"�1D�N{�K7	�U��L��|)�8ȁӞ6�n��H�� <#�;�(�󚍗�޿���
H2Y��5-��*TJ�	ӏ��4�� $�M#z���Vƈ"Nξ�J�d�Ԙd�-�k��W���{!����hM1�K�����կC�2���2�pB3�@��F���ANR���<͈A`!KNrI�\��2t���� B�di�PK��U��j~E��-���=�4ln��I>Hl�H��[T�
j/�؛���x66���+�@�I�P���?&��N��a[�����&�lHNڷ����A+4?"��Ic��p�����!�Jaf����f����s�f��>�Ec̜}���[#ԘӵpF�L:�!(ɗ�}��fB[rS�->Ap�,O��t %�T����/�Xw!����@���zc�	ov0�*fͶ��HY�,$�!���p���hXX[���m�p0�<<u�Hu�k��̨���̱�ُY������
=x�bPU���]|zqβ/zu� �K�7a��Q��>������5���K.�u�o-�ˮ{{,v��Rzλ]�͒g�^� ��ap<��b��'��F��7�[�fR�'�K�%��$"�Џ~2��������\#!d���C�!rꭩ��p��>\P�5���5<bN���F��Jͼ0��O�����>���j%���c�V	��E��� ���x�VpJ[����z�������w�g�F u�V�}#a,���BC�]0�J
ը/]C��1�ͻ&,��ެE�6ޚ������P����[��)����΄+��YhU�wq�*��d��
������6�}J���Kn�x��"��)@�K+"$�m��@G�1X�n��Y�N���1�G2�:�v!��1n]�_����i��A����˦ż�0�[X%y*m�}�p�^�8�Ra>u�H�2�K���������W{��ˑV����4;����Y�F�*N��/�ǽ�!�K"��li� �,�����I�R�1a?����ty~�*����m�>̿�N��8�B^X,���9�;9<�ßڶ���*
�6����h �����ɤ�ca�d����=?��HR9!k*8 %_f��3�0\M�~�Z�
2=�8-aHi��	��	v����ߝT���ﴐ}J�` G5Y/�����ɧ�^��a-2�}|�����m��o�_���F�&���o�
�#5�&m��f����g���k� �0��ǟ��,g�����������,�J��&g2�觷�`�� 0?���hXr��&;V��/�&ΐU�z����Z��li6Ũ�1&�C�I�/\Ѫ�r$�@�L�j���k���`T��;;�OB$�I��_�C�<�%I���$=,���m�o_�?�~ے�vs�b5s��V)f�Pc�gB�
Ya6d����.JX`-x��F��K��A��>?5/9�M����?1���&��D��iV���Mr_�nC+�����G�K�9�/�4j�*��	Lw}��݈�)���lH�Ȥ4�����d��;�kl�+Ke%��oc��a<���T7�m�5"�;ߣ�̣�p��c�XF�����q�5��n��x�a$�9��>�x�X�ٳ��pT��l��ld�iu9qBQ�Q#R���G1�N�C�O��ֻ�o`Hb��;���?�8�\!r���]>�����C�h��O�-Aҵ��R�2	p���f�X�s�3��g\��o�+����~вq���hY��pmG=�6�U�S9��Os:ϋ[�
W��ڠ�`v ��T{�x�#o�s��<��H�T:������N���������(�YA#����Hgݵ<�=S)�.�>����W�f�NY��g�@>�V�oB]|�Ɛm�jw�/�3 	�0�aƣ-:���r��M��S�,пZ���=�\Vv߈������ɵ�f�`?����g��;��ǥ-2�O�Z0�_�����x����8ǭ�Z���i9��H�3BEqnG�T&��`����}#&���!��J}�҄k?��1��M�v�����5��W�Sf7����&���mT�ӹ��]�&ސ�
��j\T��p}w�t�D�V`����t���04�Ò���P:�\ �����)	k��~Wp�|�H��f��Y�h1R���Z��Y�D�R_���T5��H�l�o�D�bSȂ�Y$��7�/�"���n��dEAf*c�����,?0���E4R�>��|�n��}�~�UtN�s��=�e�gз�O�,(.��Wr	�M8J�K���{�n���?.�؜����e�se��^F�v�p�T+{��%����f�>\v�C*�[�R��*��zaE+y��n�,9Ƃ�Gٰ�Sev�X�<9�b�Zɴ�����U:�E�y��k]2tL�P���[9z{����g�` ���0<l�ؕ������HS��t�1=Ǫ�(���g��֙�u?~Y�O��[�ޙ�0h��s�
 c�L��p"tU��B?9���r��;�Y[�H���*fNu|V�����I��i8��2;G_(k���`"�?�ȍG����ۢ �sh����x/Aw�Y��yu��i����~���h�"摆b:��#S}%��؜��접�T�ͤj��JS�����B��&0��0������[����Tt��$��O��i�j\&�tυ������0�$ǃ�����a���͵ɇ��{���T��(A���VS����#�k�U�z�	���vJv@�������N��I�R���L�>ɟY���:����h3��8YH��fYe���Q���i�����r�;�|:ɷO[�uT�H��)�ꭸʙ?o�9v6��q�%?�� ��+��|����ԙ�>�9bZ�JJ�Z�Jݵ�g=��#�;p�ne /����/���ڪ�Ḋ�������@M(��Ѿ�x
	^K@�;�- pW�M�}��N�R�{ &�+�=b���m��ϵ��:�+��=�0|��9i��W�:���r=5	�e�o����L~�r��
��GY���Z҃��TeAL�Ϳ`x?&�h��I	e���0�CVI�quљ��Č1�mP7�Ӣ_"��j.�O�F����9�!�;ʳα�3�9���B�K�s���ఉ�䑏����	l՟.��F�c:�]�V�Z�_�%������� |;'�6
4`�e�ҩ�8��W1B��f�$�v0�yIf�j��"��Q���#p5B�>m>��e虃�N<�-Y�{U)q�|CD�A6��gͲ=S�@'�,�[�X�2��|�/'w����z���`A�.rU��/Oa��E�����4)LF�Oi>4�s��W=)'�i ��P��W������;�"�c�z�/!�e:f��˸L��V�=c�S��!9qteR�ǯ��H	�#��.�[�	q_�u?���.P
���.R
�%`�������*r�̲O���X������(jg|���wi#;�(�F�Q�*Wz�Ԏ�����h��:s,����rF�8v��nK)Y�;�yV�$��)Q��_��=�3{�7�Р��c�H�.,���E����떦ڧ����N\8�B����j�Ǐ����4���l����a-%;��Ak�3=�g�|O��/!Q�~�n?v�j���c�)�T�e�~-��ڽ�3c-W?�&���N�}���y8 �G�? lk��5^�ǉn�Kp��%6���&�E4�W���*��?�4%0eG��U_���4�c������1�3��_M�M�{<���d>j/�0�r����|�eЕw��5G�c0K��QGVdS��Z�a��#P!��*��˰�9�_�b�|��9$�qj�Cje��!D|d�yi�����ƫ��8�_�v\+�H�S����Fg:*~lZ@A�����L����|��cvy���߀�7�������q0�v?@|�~�?)�L�Z=�O�Equ�)�VQ�'<#A�t�c8a{LY��� � %"�>�(@S�u.��ě�,�Q?��G+/�य़Y�})��z��u����u),p���>{u�D�'���+Wq�8����Ưl��P����egN~N�0�w��V����j������]�.F�*���7(-��@k����a'/�{��y].P��!���=����۶�b�8X�ז�Bn)K)ݲ�zd��@-��k��Ň����L�]��g�ݧ�\�݁濲��nJ�����/1M�&J�րwpT�;M�R�c�y�s/��媬n�f�� ����]��Cs���r�{�HEVP/P��/8I\	RB$?�lVXM��n8KB����Ը�0Qdi�mB�*<k#EV��}�k�9�z'|6����1;���y؂.��C��DFBUZ�fR����PŢشƠ]/�O�.r�>�Ϝ[q�텝^�_� �?�}�y�}��؂О�Uw쏷���ȕ#�p�"-����W�̉�5���GLo)�ӭ*�腘�9�����U
#b�G�F��˔��p���,>�f��"㬿���Sxͤ�c�w��j�v�3|���I�z7wd���#�艓'�/Ќ�SX�]������$iIꢼ�ALUĪ�6��rq��6 ���W���� �D���y��Q�7ǒu���%���5�{���������H�h*]�I~"���&KG%`�v���d"w(b��D
�{�IJ�I�(�G"l��٫ �2���Bi��~�>�鎜��="������H�Hꉐ>^� =�j��}E/�,��:��?yJ��2��1��S�N���O�͓��F�<B0~U�xle8�B����xH�y��i�V�� ��+"d�����n=���*˩P~������;{�t�-�P�K�w��ء@x�JpW���b�"a��]�U��8t�j*�Z^�vn��ĲJ��ۈ�HU3�Am;�����~���O��ך��,��޳PƂ��c��!"�t|�Nk���r�'i��-Д�k4`����>QD�`�y`��Q��;D���g����iժ�W��Z��._�e˻����(�~E���Y\Nְ�����+��e�'�'�F�!kZ�%6
<Q �IH��->���5�e8wA+Ƞ�Zls:M��HR�ż�{����}��Z�2%$�~��Nt7y�wm�+���JC�$���gRY����x���{��_��ﵖv�9��\{1��C�|Z��ky�c����ֈ��x��'��{,FL���}鍑)��rZҜ��Ю���3�ݱ)�\u�n�>]�%o��g��B����S1���V�1��2����`�Lpy�i�� !���$&�0y���G�&ĈÒ'�H��I���ML�[�H�w�����;w�jy��k<�N}Ҡ������D�t�qTL�	�iS0�J'�sϐ/����/&8�[3���4_�n�1�S2/#��i"џ�C})o�8��?~�{�U��5�:����
��3<	0om�寇�ū���4j�����A_H��}�k�?L�u.��sr�^�u|�8�s�˿��]=<�$��Po,���&�.(��tȈ�}ƃ�`��h텫Xx]��E�3U4U�ص��}��'��$���c��G���0� ����F�HX��ә�\���Y)]ɂy�N Jy@���*�V�����e�	��D/���g;�hO=�a��L��D�.=���m�ԙ�����W^���Hg��<�Cr��X��p���g\�"��R����y���k��l���y{��t��˕�S@I����d���wp�-&g�,㊯���!�a��i�,,bErq%W��~�D��t~B��N7-�mKP�x��s�J�U�w�y���oڀ���|Bb����?x�JlM�������s��_��.�Hݟ�
��
��fΦE*���`���ǯV�Oc����aens��=̭��9ͣ�\�炙�ڙ���p��k֏�J�m�|KR�E�,"z�Z=�#p���@X�4S����v��T ǎ�\���ˍl��nf���u/����!�'� ]$��{՚��Չ�Nc;�tw53vwa�.��k㵘�ߴ5�=�\�Y2�����	n���V�N]�A��s��ڛ΋5I�	�d���僟��i�I�(�)	�&�M����.c	Nއ۫\���2��:�1g�ޜ���V�o,;J��s������T�0�h��B���d��^,�t�9��KJQoR�ۑ��]}$K<5�%@ԩ����ҕ�`C9�=� � ��6�Κ>���^i�_-�ks;]�c��t^�gիo$[^/��3��3HJ��`	?n��g�>l��Kݧ�D�����Z���X�e����)��j�'A*���iSi��u b����R�F��E�n��$5س�Zyb�X��Wy��Z��3M�D��s5*e+;�/b(�I���GS:S���D�c�>@=�A*^��=D�T��E�pI� ��y{R�7	�(�j�{�!rP��G���; ]~��c7E59:.>8u�3��f�����V'�R��o��~�C��l3�!���t���E<{�"*1��8�|�[��;l��G����W�Y��琁~�>-ߢ�xv�$|�EY��L�a��<:"8��G1T��UϮ3:�=uT_�>�1%=����椱�ߞc�B�����g>{�q�o�F� ��c1(>��P`�5�"G���l�_���p�3�>���އ�Xb�����;� �9�d��KϦ��RSkZ�B,�/��68gq��4��s���HNޢW@�}U.һ3��Է!(,(�����\�ڂ)	�	l���w����P?�3�1��U�4���@?�,��-�FlC&(qW�� �V����>�$i�'��)l]�|�J�c��N�C9�`���[lE:���U�i0�r&�rq@��3�HVd٠��93���ڑ��]8�Vv��[(4@cMBҥ|$�2C�V��'�@b���tΨԱQf����:�IQ��Ǟ;@�9�xa@F1�`���p�n��)�|iNN�!���* 0/�}������G��vKQ3�B�:��eH�|B0�b���L���zj��q�60���o[�3�|�g�{��KuОp�e5A7?����G#"���`�E6��.Ou��~��Ru@����z���'�/��7W���7Irw�k�w��-��fd�*bd�)�0[�'ġ�?.	�;h�Dp2Q�@(s���2��2�uej��೺^Bc~;X�٢/n�^�����%]�v�{D� b�xPD�L�U-h�E҃��F�Sf�\�G����%��XnUWD���^���}���Zy����R"�+���u���|JJ�_�
��fu�آɂ6"\�|p�]
!�1�A&��XX��=G��|)�2���O:61���/iػ�ާkQN��چ�Wy�֥NE�����^��Vg�y:���\r�ܲ�{��.O< ��g�F��iҷ��ς�%5x&什K�`��jO�O�2�	�:i����!kYKr�R5����CΖE򽓽��Ӷ�򁯏k�BL�w�Na��nI���H�UN���`Sge��-,e[ ��~����V1Ǒ* ��[��9L0̬Y��-,J��A����y$>�?�e�XI^Ŗ sj~���[*�"Ӿ�������bӤ��u��������i�>�J�𻏈��2Jk�~-:ݤ����Y�>��B�!����g*a��&4�A��rʌ�"2�����?d���ˮh{��b�#"�[}3��h�� ����c0iI���x�>��'��"��d���{���2�?��z����%�e3Y�Ɂ<g�!�Ý��k����������m�]���ƅSN�5�w����f�I2�������#$�����V
���W�K��݂��4���]VʯM�E�
�Yӌ<A ���.M��*�8�H�h<����޳�T��P -�:�`o���E�3i�k)o>�E.A�j�$#��Ͱ�{��"� ;Ļ�L�C�Y?q{+��#a����	<z<��z���&��l	�H��8�F^�����?�8�O�s4J[.���v�z�Jd���[��M�Z�ᑱ*���Tb�F)5���J�9h�I���de�o���_�R�z��:���ٴc^4�]<��+D�/u@����k�G$]���l�����G�%Ree�����g�����Q�� ���(��������ˑ����-�X+=��怩��>~��	��.`�%]9�%'d5[J (%v�`fҽ�����9w�&�@Z8O�[Q���p�;0Nlvb����e6�|bo��r���H������\�Y!�qy�:�/lM�F�)o���lz����8[<3��X}��#�3�m�bߋ��^ Bu�z��v�������#�vk�.�j�e���~��<�a �o��[�t����ʀ3���e���%c�*����s�s�NK'Wv�AS��Ӽr����p�:��������Xbz-?n*�.XJq�1��YCǳ�f��j�
���ΖfA�|k�����VM�I��O��![7I��8A��t�k��Ɖ��~���pq2���L��h��D�b��`�y���� �����Zv��0!��ml��5��H�l�q
�ܙ'���w%�F��>>dг_����A}]�����6
Vj�lu�a�
��"���* �h��� c>}a��<TT�L�5��:���k����'B�1��p�q%�r�7E'��RObhѷ*ʶf�h:&7Cl��"��ey��f�^�@nP�*�-��X�D���^[Zf�Ů���Ui+P�7����,�P?�ǣ���O����%S�Q�� ��Z��H�V�q��Apr#,ޗ|���]����%�O(Ks�V�`�Mo�� �|���!&e�ZZs��vh.��J��h��4����
4�5"VX�g�Kf�::�>��^�Ҁ���S*;�H�o9a���}v1ߕ��r�e��s�X��R9��e��	��B����v�vO�X����7ӷЧ���y�Z�e��s���=#cM��n_oJH#%!N���ғ���ė�3:L�%�rNIp&��`��W�2�{-!�(���V]ʖ����H�Av�����p]����DL��Ʉ�jh8E>��Ɍj��,l�^��n�c]��O~����E�g��hD�F���|�M5q�}��ߛ��?lGx���P�&�9��gk0����%�E�,w��������T�^pgr���>�S���6��]�IwgsF'A��w�>P[I�e�F�������Dŷ+O������_Y2��T߲I�o�_�-̐�>%9w�1M�?�5��Af&�we��$):���6O�0���nS'�'����Վ.!d���i���,]DY�e�}~�>�ko
��J.��ǣ��E�͟�c�%yL|�0�Ãƀ��Q?(�5� m�w�&��>o�|��7�ϱ1��}��z��,\��1UJw���J>���XO�"�o�(��RU�6���j���ތӯ�wE�����g�-]�+T��5���T�bK]���7%�H��v�pΔ	�^�I�TOil7G.(�����J4`��������wyF��!ukpF���m�-$|�kk"g3	������_Έ��`�sɖx��J^�����c���s����9V-�G��E�W?�rt.��<������wB*:O��0f@�������o|��w�\2a&sTྖ7C�z�K+�ԅ4I��H���

Ո���L��f����n2�k��ڷ!q�
7x�L�$�`��b�F�#(+�ݺ��zҘG=��/�j�_n�[D$o�3�!�h��]��E��ڳ������j��P6�6����Y����g����]�����`�^؜�J4��>׫{~߻�|ᇈ�=D���@=2.w�E��PQ��vC�j�>�JU2CztN���Lv��b�T&�DW)��3lHR�f���4�׭�%��)no�0y����se��0
��*�[@�,҇!��G8��T�� ����A��`t�U�Bnz�j�;�X����(��)V�Я�nA4^98:��͆��뗰��bi�$�sx�$��8Mol����g5�	��/�A���ݻi��l0k����z����m}~���p���w�k�q�e�l���)WT,�?�*��yw�K�V����i��,�9Y�RW�o���0KK���݂{C���+����IN���P.�^�C�.K���X�[=$�+�X��p� �[vL��ۜC�9������Cُ�`�r���%C�W�-�r:�^$A$�)�SZd�g]?D�z���!Lh��y�QrW&M�����<�}g9I���9ZyF��Bf<GU�Zn4~L�\9���:#ZY��<U�[���9ӕ�J%XYb:ە��.����O����'������W�<Zrxw���p�I���}v��|sO���)M�$&�|I�o,����e���'��	��~�!%��τ�H'ɝ|OI��x���	�M�����ӞTm� �m�K��]j�}���"�֮�md'��p��Z31Oa���]}�p�8w��a���/��;���)s�(�sK���J+���R?B ���-e�o$#Pn8�X��;���.��w����↲����}L��@��ԯۍ�1�W͈dz~�n��	:����S!SFBޟ�в�r7Y�&�n���Oa,;(:��&i�Y�pͼ�я���ps�?��f��'@����h��N��7ߛ���H�Il��*:W �*�1$��$J]w�z�|��H?��Yu8i���j+b�/���꿏G��;�]^V�����U�MC�]���>�O�s����1��҅ᬝ�]�%xe�������'a��7E�0�z���*����������"�0��H���ݔ^fؕ���
��D�-���K�iDM����7sY�T$�s����:e����>�#ǁf�^��UZ����W+��˛��:�!N>�`��"K��κ7�c��ܺ���}�y�~� ��j_��]�2́�\��t�Z5ƨ$U��x,��IIkDͶ֙�xg^���J`�A8�dNu?��*���ޟY-auG�H�y��ủ9�(��oj1�����s�Q�2kw�G�����`���J�Ni��5�坙!sk�?�ާb��,������KӜU_�����^���Sǉ����ʡ���i.���֖��Z~�p�Al|�A�q�� 2m~��X�����:���/_f���X5>��x�>�z�-怫��L�چ��s�����#N���̻�����D�4�?B�1�N��[���.�6������0��Q��A�5�w�76h�=��S�*�_�]j��[��-]��3,,7:��(q;�u6T��5ڟ3��#xŢ���8�o4Z��s�N$�z�Չ9q=�𝚼�Ǔ���dL_\1�\�æ�#����0�<��5��d7�V��nK����8�;kkY���21ؼ��@�n=fց5X��@�
/�-��n�fjo$��U"[p��GL�kό���A�����M(�d3aK�\�.B�g�\��_���|��ڙ�@�����B߷�V,f��]�t�]}�b�nDڦ��!���x��ĺG�89<#mX�;�OͶ�ϯ�\'�����鏃/ζkP�,�.^P��3�<�����8R��<���)�V̊䖟�D�_�\��	��X�G��MN�_�S$	sz�%��`f�
�"Ca��W^?��[����x�iG7`��i�C��Tk�z�E���Y7�(����L������4��F_9�!�=u�	ˋ+$���.�~=��Hӄ�G�P{m�a�i�� ��o�o��c�~k�7K����ع>ە3.��J�������o;��`Al�wQ�M�?�����Ն޶��鶽��m=pj���v�t���A��+�!����ZP
c��(�W�1�jk"<-;�bd��	�I䂑Z������4Q�Zk�s�L��Pg�#I1��8�be��N�e�b�3oK��MSy&��� ��,z#W�/�\0�zm�8�J��8G��,��9��=��~�)8���#�e�8v�oeB���*���#�Q���?��o�`�{���4�q;�+lWdI�P�J��F��4�9'�/�+$�iJ�'��6y�@ˎ�s��>��!�AL=>�柄; �����V3��s:�lR� �'���ꓡ�V���,G�.G�t����B�Rã��8� �tVt��6�Ȯ_�ï\MS��Ɉ�鄾p�2YfF�/g򉅁��Qd{8b�`{��ϻmS~��q�'�� ����+�l��<�i��\�U�ʟ�8+���Y/��.��#*�ǊD���E٬�>��<Kn�P�&�P4?$����H@)��c%(9�Ef�����(�ɨ�1Y&W>� �T�D/�,:s����i���<����B���=x<�����D�n�������b�4ػ�5�V� ���N���H��IR�ѝI�G����۽.?�42�(�o���
aIi˲�����N*����t����1��w�צ"e�.R�)�U
bRƔcn$Q5���n(��~�E?���/ �U��֔�H�"�%��rY�Ȇ���<� �V��+i3�v��V*��?��p��j<�����P�
�x��o���?R��ӑ��z}�{�����ut�����w���l kY�F�����I���g�����_V��s��X-n�7�N�OÜ~Z���9��ޠ�����m�j��"���r�І(rԨ�Dѱu�Q�mA�.#!PRR�+c|*ϸ���w�VM�Y�&���.�˧������M�Э=�`'��7�>,�U��R<�����&p|��4����{�A��-yXSe��\5����-��h̞�e/K?�<q���,F�E;��V��	����n)���*��ߴ;qٿCS�QB@�$1�̗�h���e�U��̽8������!�  �Us�~e��N�; ����6ޢ�d�^�ۥ���(�|^\X4�#G+}���V�Z�`V������5A�]�^3 U��r*,�hvD�����V:�i���g�w����A�n:,_��=��u�Y񀮫B�/�g�M�YI�y�;���(�`
�D�u�7�J��,F f�+@S㽃��n�����a�U�y|���W�u�M�J�'渣7�ؖ�D�M�)�s�'�s����%�f0g��թ׸T�T�B��*���&�7�9�C�璾a�)�^o,��
���Z�=�\h?�Ԣftk�$���G�:�.�g�/��M��gq̧�ܘ?��������yy��Iqf��.�#ݩp�3��W��/]ׂOs]E��㙵]�"�Yg��˼����?헎rF�U��!�2��)��-��n��:O�ɂT�1��1���a���ٻ6#2�j�������UE����!���p2^�5�z4LPu�}L� D�c�X,@������"8P�,��W
˟�K'4�1;����Jƪ�)B]('C��a��X�ǣ/?N���Y��?%�[,)�&�R|C��~��E�N(ǈ>G#�ƚ�[̀zoO/�P`�i�|5��yţr�:�����V{&o�y��t��� #ͶLC��?]`�^mF�RWU���sY}p��Ì�b�I}��k�L2��I�TA��t���������ˠ�pC��X�i�8�IQ���$M݈�Ç��cW��b���i�*M�_n�_,z�#�n�W�:��~���,�m_ƕL���d,�4�\:>��:�YOT�p�
4�����e;�.��[�t��vTE��	A��b}� �����%��+[�������W����Q�h����0��v��ԟ{�3�I���1�s�{����+C�m�dVx��j�`�7��3��&�����}��L�d���c*��"���W"�|���ח|a����y�,�[���@���U=IM������
FX�A�%�XΙ~�YJ�T-�:��3����y@��&�С�s��J��|�P�=sSi���MRXuJ���%����>���3�u�.��|�#M��,��} =�G�+���Ӿ��R����y�`�~�g�z<��y:K�`�$_��UCe� !����`]�	�X�U�"��qTc�K�x��ѫ��B�Y:=?��pgؖ�Yq�l�ai�Z =�n��f��c,+�ݙ��	�F���ƻef.���x�O�:��F�BB�1��P��.&�M"�n0?���P"|g?D��n`l�:X��8�Ӏ,Z5�{Y��c7��djKR��tA�霏�%yv��SV����.��2%�/�<��G�Ʀ�p�@I*�x���;��JF�>�6��p����$�&���HO��iZ�T��uB���nֲ
��Qf�b$Hw/a;���I�|���q&���ˎ\�l�f�,�Fh���! �[6t��4�8�fF7N��)�r(����W��c����Þ�N�V7�]o�z"9���M�pα��cK�'�2���peTp>��Nf_�A/��
ݗ���|��QO��cM{�年_�0ձx���X�m�A��ƒ��ٸ�`M��3BtZ��Y���mm���6ou��Z��~>G���'�0�d;��5�>Ϳw����c���-��b�Pi��]��ϣb�����c���[�@����\�k�3��r�AS^
��a;�J��I��C�M��D��L�V��ĔDB#z%���+eM��Ӑ�����}������Z�b��i���1jk�� 7VƜg�����(�Hd�p�7ü^ؑL�/��2����h�e�Vf����Q��W�
��i$-Io9'�y ��MQ�gx�X{�c�UȺ5[��O�<���
!-n>%%�� |�'��#�{���e��Nm@7�R~�`[j}������v	�i�^�&O�8��:� ���{�
=B4|?��X�{#`Dg�&jT򦹇ں�����]P��Ƀ���+�A�Z��{�n�G�};�l�4a:od�	C�k� �y�C��sD�L#l�������WR�/P������$��V�r�PL@��ۀpXS��� �O��G�W.��68U,Ox���7���o��8)y�Ag���(�c�v՗)�z��x-x���n]�Fz���lC�&�*��6O-y�/�V��vSiܫҫ�y���²�(�+�y�-Ws��V�|؁�I�O[��S��gpk����J?[�c��o�H��{QrjGk��d�ԅ���yS�3Z6�����I9X��#�95r�@3p/�jW��� '�wr���q��8R\��C��R��j������\"���{���{�g\py��#�~52�-�P�`S�� ���t/YAo�j\��p��3r��;�8y�&������hg�ݛ���6È.\�ґ´�A�9�b���8�:�,�w|0c�������hW���1�u���������e|�Y���ukj8y���c���ೈ`�f�L���PQ�?y��7�K����2�}4�ٵ�"&�H^^�׊/�����W�Ʈ�ju���ўK�w�k>����a�J��=�J�ܬ*��� ���T�>;�Bk����~zٹ
�K!(�[n`m�Ǎ��8�?��d���G���.v5�P��ddy]�tA+7�S�C��>*ƴ�#��F'�=|2���,��(���)��[ɫb��N������l"�2?��1y��{�6�m'��hV�Ӊ�)�������WF]�z����w$�	)�E3,N���e�RH:-��S/��:�`��p��'�B����S��W;��y16�x�ե�Q��|�\p0�g�qk�Plao0�6풣��HZ�%�4�y�H5��š�3ɋR��9UW���Pt�����1~�s1"-��҆�8��N9b�����Re����1n9�j��%i_�����b.��T��
�d'1���o�#'%OӣlV���'
�I9A�/��`���r8�Ob�ĥSߧ�G{�����:>p9y�C�Ց�<	%�M*e�V����gn�w��Qf=2U{&������ђ�k����v��p�L����[�7���j�j�D�h��~��H+eX�EK!���A�L�pJ����sW&2�77`���צ@����'�.ӳ3�g�����V�m�g� RQl�Aiq�7��D�7�\ˠ:M�ab����T��8�J*��*���y�����QXF�n5�QF��p�����1��7m/��7��B�=`���b�z�~SK���fFL���wy_�%��|���gk?,�Dp=��.V�X{Bp�ܸB������)���Z�C�o�D����+�)�֗V�6��#x78"���-��jD=�Q1�Ɯāa��%�h)�ލښ��y���?g�"F=r�3^�Ҵ��I�H
63�g��O8�{�h�^�22��}gޚJR12�aH[*H�ht�IS&	��['N"9�C[͕`vX�����q{^���n�=/�������UP<*F�0-�F���C�WpTþ��/�La7��=B�^=�|բ�Hu�+��g4��E%����5"8��S؈���O��C��N^y�2_���*v��L�1]�sJ�85�߆���,Df&��mzo�*�������mP�v�Bg�M!����*"��Ku]�W��׫@�����t��d�1���ID�n�r��<iފ_B��1�JUxj���/a���6�V�&��1έ�7?�d���H# =g{z�C���4!�c%�Թ�z@���)*�~�@-	�b5��� �SЁ��(5��pO����	,Xx<*)��]-�_��|�7�~z���W���8���O��*f	��F�D,�H��p-f�h9�tcy]9��-Ԍ�!鴷=\�:��^�F�k�|�<�� ʜ�=����=v� N�@�۷.���?q��#���~a���K�.�B>��AXX�{��`��cZ�޴6�q�`
{���Ѕ'�?���k7;�O���ښ�y�^��y�W��2���m��Z2�eQj�����9��'�s�CǼ��`�m����14~ h��[�=f%�q	S��DGrS^j�~��_�iH�V��9�(�*(�ڞ�7��"�t4�7�B1�xz�rm9�G���2i�a�Fh��[*Z�?MA�@���3~v�qȔXJȝFuz�6��@=�V߼�wٕ�DQV2^,����L��'��}�x� �W�6[�Rw��&F���!4Ig���.l�?O3�����,C?|���ӎ�y]�?G�(��@��L�Mk��!�n�	6���*���(U�9����lx�`&��;��*�]�Pс��Բ ��>��c{\�R���t	����h�q7�S�e:�i��J�2\��"P�p�<!<P�b9�%o�Q���{��v�A�üת�;���)�RM��1���k�B��գJĂ3+�U��M گH�ɨ+��@#<��!E�J�%�):h���
ߊ^li8��kw
���nm��f�4��uH++*@��̿�¦=t����9.��+������Huep���K2�―.m���>�Z���^��ڈ?�$�*1�]D�O��R�y�m쓶%c�$#�??}apU/D���frS������[�x�u4'5�
��\ถpxw9����~�u�C�\A�20�X��P羅<�3#�F�{�U�gr�L/�8R؃s|���I
�w�~X���KK	��ht�0?�UU)�g,���r#[�0�c֍��t�������徊��ˤ[B��T�]��MW4����Ɖ<�q�̀�J[�o��G�$>JRY6��5����z�!��MˊF4�׳�==�1�K����zK9F���2�	�����|\Z��-�d�$Wmu���b�:D㹪!�K�.���[���I�A��Ⱥi���W��\��Vݩ4�lf�7��S.��
���9^�Ňf�8�o��*�ފBM���J�X���M5��q�O#�3)P&jj�?�:j��A��x��냍�=�##x�8mn��,�J�A�w����V�r�Y���'	Da6i䏯\��������pC��+�S�#z)>�U�!g�.D{P�g�����C��I@�W����w��κ߷��9�*����t��J�j�L��F�<i3��I�r��g,�@�i��v����^G��FIy�#��L�[��0˪7���O{4t{s���%�5����f��3����O���CY�;:(߭GX*�e��4�:���	
@³Z�L��`$��=�8������/wjF
����ǱO-Wk���%�?��%x��DM�J!��R����(R���3���S�w��^2�>;u�n\o�$q���T��kqYxN��pw,Wr���e�{=�;�0�c�����O�_A���S~�I.k�`����|a�J��2	�g��rh��|�0�����m�2<#�o_�WUY9������XeY�M2���c&�����rQ��O�6��������:Q4FǱ`xG��WղeFCR�d��Ҵ���戼�o%�Z%�ʆ���[Z�	����(�B�V�����;bL|�lW���G����G��f��=�_��@��*�io?��V~��)���<y�� ř�G7� �XT�.��/a��8��:B�rvCSs"���S\�p�ٱ�Y�4ƶ�H���j��瞞M�.��!*�ҝ�7I��g���}R6�\���FBI��P{�
J�A'$S�g>Q��� MݵxT��V1��b�$�h��m��WǠ��s�*m��/Osa�3��f��z�4d�'��_h��"7j�y%T�\�O^	 )@şW1�u���y�ѓ�>y�� ���=۟�w+�T��&X��=��'���}��"�'諶�_T�7w�A3Kr�V��F>�.��r2g@0��qwY��f��� �!F��6s�	���ā��3^i%M]2N�|�6!U��.H���QIK>q�-^��Ld�@�0������g4���]'I��T�$�k~(�8I�9�Z�E�a��Ԙ9��J��������X`��e*Kj�:��(�t�u)��bP\e:��y`�(�<�X�S� ���g9�(���y�짊�'s��a"z�L|�Y""�O"�[��AS`$f�5��\ĉ��x�A��Kѭ���j�=��o���ߧ���-�|x�WΝ|e�����eR :���c�L&Hu~+J�)4�逸��L~s�%������ڸ�4��\����b�ᙏv]��O�Df����y���%��j�*)��_2�o��,l��*����b�=>7��N�j��6�0��|Ϥ����.�
I=Mx{�h��7�{���4PB�A�K���05�nc%��[�d�ǀ�S_���k�\J0��V'4p��.��夒ȫC�5ݶ 0n\��_��2�{?(����wG#no�����W}47m5�\UJ�]���=��7k1�A�i����<�\z�T�����X��l�d�j�K��)8.+?'���])?���HW<��'N��8�d8����?͝G�Y�r�R���l�����5�������8#����#��Y���{5ܯng���:�-�vgp$��8E.�P,��j��*ꓲ��)od	�:�/�{�x�o�jv�`8R������-�j�(c��>f���,���4�^���=#pDʞ��h�^��%*��fHXi��B��u��~��	̺C�@EЎ�Jxg*��<�aB�_B���#w����:�����yVx�y�eb�������vR�������U�C�0�'\5�s��F<�埕$,�@om����{q�<͋��7�u������cw��S۞��|+����.��9�p���3+9zcD��e��p�3�~G�+̎��}��炠}���RhC���3�7�}]I����me��S�Q��F���.�Iw5�J!�\�.�:w7=�T�랻J��H.����wbd�?�L:���N�+L��'(?�o*4��%��7b�f~��@z�E*�^j�sd#짥!ǱY�Y3����V �k��~R���%�s���&��"��+ų�Q��T���{{(��Sb���6(ہQ\pF�ځ5s���Ώ0_a���p�n����O��E)��;Ő�o%��m
���$�����O��0O�;��x&QP���F��(#��X����D����@yB��Ǯzt�v� �p����� �נ���(��8��������1s�w��x�lO�"ϑ#�y�uZ;WИ3v�)��Z�0Z�����Yp�'��|[lNR[T,>�:�E���פ�P���/~ޯp�C�_f&�����K���m�2�"_1@+�V�.<]Gr�-^��o;,�3�@3+�fr%jErO51%�d;?8鞺������r[�nbڣCY5��Oc�B�N�(�b�
#	�3��k�9?��&���F߫�~�:����)��&cY�D�9.�G�+�{�|~>����E|�Oi禜��XgZ�;�9}��Vl^�<�?O�_v�a�J&_(�Qx��\�k��/��p�%"�ࡀ� ���@���n�-���߳�
9AK��Z+Ȥh���&��=%��q1�3���OOsd�qֺ
�7u����n��r��knXL��w]�P����K��C�&:dl�;W��{���,[�H�j��c�ԯ=��j0�T?|�?|Cj���N���P(^���b�Dõ����w@@��v_H�4���� �����x��n��B�o/�0�̿��<mhx�We@y�p�\�]y|�<a�զ����Ss�݇8��c*�����4�>�R>M]��"��S��s�}nFx���hu�d�@ ��e�X4x»��
�������$b=�s|�y�V4@q�E8Pg�Y��~z����ϔ:��� 4Pa���Nh
|Oq���x�*y��oθ4�,�m��T���ѣ`�JGt�\5�o�� ��Y���[���7*3�6�>�s�d��x�	bC�Hz �]���Uw�(�+�B�2]X��G�j9����_4�Bї�?�p�±�R.��YT���c�f�5����I���Α̞$ʄ�jY��9|�m����v}�Z:ښ���Bk�nw��x��!T�`3TM'ʛ�	R*w;R׉�*;k���e���5oQ.��1�Fm��,|��s�R�i%7y�s{ �ḣo6\+�ަ�V�ŀo��ˡ��Q�O�o(�Z�ft�xU�X�tu���y�f���)�&�G0��Rn
^7�� Y�f�/�o<s������:�5�{=����֛ap��s��+��?�Zj�N�8	���p.|s����G���u��S�uY��=��CB&aBj��x�Ԫ7����S`rq��+-Uݧ]�p���	�D��p�D��h@�W.����L�L!Õ�Hps�})�͉Me%u���.�����uC {KP7{͒~�)C�d��4�x��qb#2(�u=�[��G	ެ�V`~H��ELqۖ�7/9�'��/�$� 4
�Z��HZ
~[qQ9&���4���1\wI����n�49nqK�;��/�������7KJqS���פ����2w�C��vf�O4�D�D<�a�'e��W��f���0sٗp��D0�^�U���7plZC�p���w�Ȟ5�u��6��\��%#��_�؇�r"����JV���X�GN�ޅ��)�˄����Ħʶ�%ޱڵɷ�t�0�.f��-k#�X_�\�1M�yk����o�=�[�@�d��nAr����rj�.J�B=G
E��w(��C�Z�K���D�3�6�Ic���i_P�̨�a�� �#���	 9�\��8�Ġ"��R�#��|U��E*��ťh+���䱢F�J*�gi0u��]���+���م!)lO�hO�v���M�>�a�<���Q��sS:����E,`K���^x�d��㙡W��gL��SJFcSa�kL��Y���ٺFߗ��|�c#E��ج6��HNl���mi���̏�ʽJђ�d�Ib�p+����?��\�/�9��	|&n�.������s-v���T�w�f0l��.��khDh6^^͈	x��R�u�i�:}�A�����W�sz����8�v܁�������K���H�Gx�J�5�4;�<���Ǳ~]mVP]�X_P�����K&����	J�U�L��`����ijdheH�RN�)ۊ{�#�)�g0ׁb�U���>���Nu��.�����*�exX1��	�J�@$��"�#t����!WD��f\�����@��6���񝶼��-t]���{�Z�m3�j	�,����w����X���i�X��rx�F�a`��~ڎb3�I�u�"�C��D��I��dc�9�������� AqzG�@�h���k���#�v�P�(����!�ݙj�g�&�vKh�"�%�f���01�����?�s�Z�pǐ�Y��Zö��~�π�#y�����{�5�N#Z�#�x櫪�t�3�v����������<eo�{=x~���[��:�QC���cd��)��'�L�؇����s J������e�B"�� \��"��0H�]�o+cq�R"��%HҔ��$�ڍΤ]j�l(�g\�E���(�~2�U$i��DaWx6�k����:
G;5jY�I�P��˻�/���*?Il2�,fYx���=�\H2�3+���B~:��d�
e�-�l!�on�~���M?/�W]�"� U0���(h'II�����q��{3�&w?��b?�U%7��|�5O�q�8�<�<33���3�Ӹ
x�tuSW8�H��N߱�X~_�a8�فW.+O��֙�bB�{3��1��r�:���|MYX�Ň�\�}ި���ͬ�O�3MJ�6�;�8��,�K4�Qd���٠L����v}�����%��F-q�����#�n6��[���h�R�g"���� o�$� _j�=)��y\���܊2|��ۛ�t��[Ҭ��n@�{�|]�&�� K���S��c���F�k<N�	����R˅n��Y���nA�{#s3�8IQ=��n��� �=??`���M�\�n��
�5�cy��y���9���ȓ�Fy���Ꝑ�$��Ͳ��;Ϝ��	:�RJ��pi�������������+��=:�nZƲ���|��h�Z&}��BT��m�E+�_2�n�|ޖ�U╙ݯ �������]����஻����{|�Wg�#���.2q�(�1⓹��u��zU4U[��>s�BW�<�~�Fc���,@kl��k�T�]�����boqi%=@�~�f���$9;箩���-R��傩�eAp|2ρ��x���.��h�̠f�$��\ �@Q��=p�ä6�eډc���||ء ׎QCL
͋@�{m���ժm��������LJ����@�4,�}�y�]�j���A2.Y�����=��#���\ɵ���쉎Ь� ��c�A�`�u�jH3�c΂��"r��n�� �/���3�ҽC�t�M`�-����	j)��f��29i:Y8e�7Lhŧyv(73M�Gm\����r-���� ���_濜��@\wV#*�o��_��?�(��:���E���V .pz=�[��Vȶ�<SeAA|��0f$|�5����t{���=��ϳ��@D�^�ڳ�0y$}�K��J��@fT��s��&C�]P.t!�.$�b�t,�o��l����"ܑT�e�R8)���tW?&_��M�(��Z�v�1s���Q���'Vynd�\��V/(;�{Jc�X��i{|��u��Nз�s�IH�H�;@0���F�l>�irx��U��|�U΅��oa:QQ����2�C�y��ᾒ(�N�Q��ߴ��/�<�$r,#!XD�m�j.4�k��wۋ���AX���#����D�>�*�@4���S����"p˄\�|�-����$b\]�y� �~%�J�hS�If��t�9N��2�b ������V��Wgv�w�M+�#���y�ۂ׺�J�s���c�8�,Q�/�W�	�/ޝ���֞��l98\�pd�.�&�T4�p#GD5�B�t�Es�M�戂ӄ�=��I�\��/��R���V��Ξ�<��R]w"4n�S]!��=�G[Q����g�i�� �$����w#P�K��f�ʩư��FM�eQ��:"�Ҝ}�=�|��GnW/I����u.ÞNw���鞦 �|�
���'$qc ���2%���eh�ذ����X�)���1�I�܏�\�F�Kx�4�M ���_"��z�Q�(�8�E��a�/E:��V�K����ݪ�~,��w5�	��M$Z{�����#�g�iV*���1-���~���^v~�ˁ�'�A�����q����f�θ-P�7�⅙�
	�7ENU�Q, �í@l}JE5�&Tj����豠��y�&�H#��L���
�0���H��������c{��P0��%+Y��z��B �1H�u0�Q����ڮ��%��ϐU��~y���R��jSWW!vֿ��7EcFR$+K�;K���֡�F� ޞMe��r� ޑ�Q��%��4������-luЩ�����E�p�Y�E.W�۝î2�9䋿by9+1���o���-KV�Ss�m���K&��=@�МL�ك	P?
�	������t#k���y��$j���b΂M�������(f�����0xk��J3�P�ߪ �`U?�Z�S��#;���O�[�X�(,�W"KJ��}�*)i$u����&�gj�6�dt JzH��d�#G�,S���Ȃ�&2daSZ1+��Ze�#�T��F�0��q	���x�(��*�@�4��*e���+��a��$���)w���Y7��S7�bA�Oq�	����Sq������0��u+�s�y�M��vZ��> T4�Q�!�~7��b6�R�H���d�h��
��@)� ��@F��J)�d��_�A�}��_+�S��XZ�r%#I�+?��B�x60�뙚�)C��v>�%25�5��M������P^g7�V�R�������;;�QMX����Z	��f��Ja���0�c��Ik:jI�*�K>�ˀ�e����z�WΌ�"���/��ա��r�rVa^��yT'5";﻿����)��������Щ�]u8�������,��C�R� �D�e�>9���0S'���9�͜�yc�uYRL�a�fq	�=� �U5<�Ձ�� M�T�U��"�S�f&�v���0ɟp���[� �I�Z!7���>�{�o~lIZ�!�">�յ	�s�6DX�g�4�g�_>:��e�,�A�(�)]&�a��o�1i�7�W>��ómϚ�����K�v��B�#��H����4C����ܭ���%��$�CAЧ�ƃ�5���tw�tV`|�����q�5��`v��6�B�?d�"�f�T1��ց������Jȋ� ��zȌ۽NP�nlƕ�V���`�kQ^�� ��z*׌/*�_F����������� ���arS���K�����FN�m�)b j�@�@����R��6��gl	|�h��pfUJ�D�7�r쭱�Q�����b �����[�D����&&ÜjX��n;W�BC6����yH�����/x�l�� $d\�j_�x�bM����4tp��Y�'b�o����,�$�M�
"���H�>���1��/N�q���2\�+p�Z�ƶo�+g��(RnD��څU���f�(��%De�Oz5���E�$)$�� ��,W��^y�Ł鹃������h��.�b J�t�!!�ms�\Ĩ�	|
K�з�_P�/���:K��Kx��L��2����f�H�X�n��fE�n�T��:��_�/��r���ȝw&C9�h��؄}g��Q};3-��1:,�!�T�������*(��	:��1�K��ȵ�eY{n�W�ȏ�:�Z�bs0�����!�?�9��t��ys�k�F�!�H2m�]���;�ʪ�J�?� ��2��z�0Qŏ�d.y�HC9���ԛw���,�]\>��"t��d-i�X�^H]��q0�I>��4�����#n�JP�A��-�`s~�w�+��
u4���0���CZ���^�l��Z,Ʋ�H�0K��3!��_�v��W�[��>=d'Q*���b�ޡ��P9o��4��K��+H����k~��Mإ�eH���^Zo\ʛ�#�ũ��t �;`Q,_VJ����O4�c��Ig���F@)v��S��nO���0j�;d`}�`kk�w'�߸�}*D��F5�Ѹ���N3�n���龒�:
b�dwrf\��dH��J�96jy�g��ĸ]����Hjx
i�9�|��X�rؑ�����\��Þ"dg��`}')6fZ��S~��x�d}�v����pd��z�so^6n��,JڬQZ�l�<1Op�jC��ܸp��4?�������A�Ŷ4QE�g�5�;xP�_K�89����c��b���3��hK" �~_v�0��i$���b���ߴ%Q�2��?���ju�T�W&V���̣�΋gҙ8DL��BR�z�l��=#���q,O��1�78��� �z��Q̣&$O��d� ӭ8o��cX�^��:��O�4>Ҿ]����uUj[��=��b��:GX'j����b��V��k�iv6Ay���� ו�������E��6��#CC_��`�э�U8&���ruzIٌ�Ĉ�O����G�4�z�;1
�������q����;��9���b��]~�C^x���ń�Ň�v萘�OD�I��R�Ҡ�G־=���g��-���g�Q۪�epG�D��R��On�m£�'p}���N�K&J�	���䚏�ؒ�ζ	�Ze2���@CA>�C�`zPC��߈��.>K�6�'�>/�$����g[��Z�o�w�A ������9ٶs��N�>q�`���:��CG,�t
ot��r�ݎ�)%�h�B�]����*ݻc��Ҫ��L��|�,��ߛ�`+���.	��T�c�y��Czppv����bӷ6i�B�@���U u��-5�+����*wq��|f���v��V�Knom&�S#�}g_=�
��	�Y��e��SN�u����f��%k� VJ�/�@���M�W��C�<t�"�mD�{]�-8E���c��_�� EțC#��t]�-z�#��	X��Y�]���N|�щ�@|�iMc�f�'�e�UQ�<E�����G����lk��߅�+��m���*IҪ�[�b�X��O┿s��HI�!d�18������>W�<��<�?B.��tC�A�S?H��`e9�
c�3���̺�8v 7k�ۮ��W��L+��6Wlh���c��2����RؓV��*J��*q��k����g�? ���f s�3jﴜ�?�Y/��
���A|�X��+i'�(��߭F)i2��g���0.�/�d��p�ț�O���c׵�������>z-��� �P2F�-���ܗ��$6|�	=�;O1�^O1L�)~&��w�w��ř�uf2�2k>0UR:?j���ͬK��lDZ��<b_�?���']��<���<���8���Xow���<�(�#5��>����t��\ �U�VI��ŲfAvo�s�����2hD(� �^A[@���GiZc��v�~���7&9_T?.�É�
�|���t��qS�������m�����d1.��>��Q�/����a1�>��覮8��� Z���0�_Zz�A@O4Uzyp�\?�_눟���п��	lg�p!oO;��x�iT��SO�(S�1�k����P�D�x/���o�F�p�k7�4�ΨL����;�N�l��ǪM��Ib���;.�Bu\N�h��|�2w9����U�=N���I�<&Cՠ��P��"*0؊�z]�uDe����Y���I�1{��7�N,n���c�G�%��>_(�=X��&^!Wͭ��ñ����"�fXAǤ��r�)��~-��5�����4}�VP�'zw^��ҺlXg�eA�c��r�bD1�Ν+��K�̥>���ԉ��!�T�9�͟��������|eQ����?�
S+��	���x��>xf�w��v ��.;��K*���� �(k�d�&l��p�b'ܳ��x�%��#�O�*��g�U�}��3T+ᾧ%?C`��x�%�9��S��i�Lб)�b�S�}�tį2/��@
�W~�?C�"l{H&��<ƅ`-���J�%���!iL&�������������p{����o�ޚ���N�ղer��~��b�d��b5��oٖ�(rL��;M�d����yl��j�֖��曧|�GI2Q�l���>�n�J�*�b��,�c�f��9�U�l��� 	�8���{��1�V��q�ck����.aZ9�
Q=}A��~��H-~U9����p�F���h�ͺ�&K@B)R̹3�'+1qܫ��I]`iٿ��K/�jD+}�h���7	��X36�laBb�:LZ������r�������g �bF%������n?�KZ���^�c�!�'��+(8b��4J�* '���shԫr\rBЕG�ʺ��=h7���Qd�n��wqJ~�>W���v��(mck )�Y-܇$Ј��r~	W�OA���X;j�0�A�"p;I��}�,�1B3�wuc2��ڕ���Pv����d�;�uzGA
�ʞ=D(�7���0�Ϟ�|�Y
�Nç��`�'�����p�]����A���D
� `��{��c���/q1�9�)�Y��X	i�Vrq��U6��A�4�4l��/��$�/�4�P�T�������캛7��0�~�<�J���z�qЭY47:a�������i���ڌ!�,��I�eV@���r����.q���w!�Fq�G�8���%~����q"v;,%��q��6֜L���M���ef�w����m��]���ä�;���9�{zD���W�m@��:7�$���!�)��ҏM:	��z�����L֘���P�W7V����̸B�a ������ߺ�+Ȃ�Q�t�U��#Qy��?��nR�>��t��4 �)Ë�푝R��Q��ck�#o� �)�/�M�`*�Rsp1��Y0�w�b�Ԣ��pEms%Ϭ|g&S_��!���t?��1rs����,<�V�X��ڦ����im��c��}�~ ��1,#��30�]�;��өdL��R����^e�u޽i�H	� ��k�}��L��@7�3��|J��Yv�i��X���ފ�!\ZP�Ki��d��̣��5�t1y/�fQn����¨~#%�<��_�Bb�ݰ��b�t��&����B���W�ѐ����I��f���K��6W���K�[{-�!]��e�3�n���g��A���ƕ�ݱ�˔��d���Im��ĉl�j��B��!�.i���W�����T5� ��YA%���R�9蔆j�Ѝw���#�+"��@�4B��A$����4�%-��Dx�F��L��N6{$��l o��$�D�$:h�_�!���fۮ!�H��~:�!u�LP�����7s-���O�F�4wa5���{?F�|�4�5� �G��_b�t��+�_|�es�#�S���5� �&ƺ9��c��*Fs*"!����3	kJ���_|u�IV0��'�C"G�g����ؙ?J�o٪���P>)��K����.WǁS[]� �u&��$OO��+ɀ�:���U�� b}pq�d-[H�����ʬ�ĺׁd�J���bJA��9gy�+��܆P�A2�L���鎦�5wF���&MAG��`Մ�g9�މ�1��/uyF��'d�g�]Y�"G��7�ߚ�����C)�k��x@*d}��dAf�4۷�0@s������j��������bh��3ѫ���!rڴ!D6����Y��Ō6�(.����	ȓo2�\B���՚��]�m�p��ZtM ��+����!jLV�6Z���#���>���2t���m�����S}ӣ���4�/6�*f�f�x2���Q���o�{����8��Pwؘ���D��na�T�i�,��tT�oWty�=鷞d�D��H�������%��z��~�.�qwG\�T�B"�sꔰ�1��*m*�M���,������;P����&:|���D��]8E��`itJ�_�SgnS2N�y����V� �p(j�����qY�o��d�|&#�A�U��5j<�8��t���X{�^�<�>(����~��Ƃ5?�����Q�v�'���Qlk�_�ݴ�m.�W�ӂy�!�e&���l�X�p2\���~~;vZȫ0H���^��@��oF>�w"�)����3hH����s�zM$|�}�3�v��G��d|~��n|H%+���}�B�ؠ�m1�����2�P��6OXF�cDр*�y��DpU��1>�]�Á��V��k̒��]>߰��;�<�Ry��?]��q���'�w9�1>,󵙙b,׉Z_%M�]�=��{��4�1��"В��q�Qy���J�5�㿢���iVA�\��y��}phs6q��>�j�>4����y���;�f(��O�4�0jB��Sѹ�m�_�[0wå�\, "\���M�����VR[l������e!�-z�<4����!��~F����F��f0���s�������x�=���c� ��H���L�k�瘥в��j�ī	pq�%��� y��K�8|�映r��P2D���ub�G�n��b�cL�.����~�M�!���⬾��1�G�7E?��5�{�����7���o��Y>@凥��P�R��
sI�
khrk@��2!�5��@�$��,�x"#�s�ж�o�y��}�|��g����tt�z�(C�yYz�Ӥ@�itw1_�Z��X�:so�K-��Ku?L/|ó���U����H¾�<�`�&mi����Jo%��:\���"6��K�{�չ�	e�LƸ<�;�XY@�@9�4ߒ[�^��B!д� �%������3P�p�IB�~�g?�@b;��:¦1��*J��I�=e��F�g׼�z��Ŝ:O�Ұ3�b%���v�|L����������z��eSޱ���S�Cm=�t�'���
�0�1
}N�"�LƝK%�)sƗs�1�8�d��g�x�Nk!�U�|GǄɡ�!�:��Q֔v�t!���X����R�P�N���3�[�>⇥�J�KRON��A����H���O����l"ԋ{�C0������J���rk�ؘ v�'�e+	g�y@��;kO*�������c̱	eIu�ʴ�i�Ȳ��
�s���V�b�
)I����qj�%nEv���P�D�g:�b�?,[�rN�pě�`��p,o��t�ڧ@���l�cƉbK=������*�S�M��>��GP B��QϢ��f�&�@��>��S�R�����ך� �2.a�}Q�?��I&#�cޖ�D:`���5\a�i��U�ۛ�,�<*�ŧs���T� �� {�A��9������>Q�3>b:�=p�� ��y��py�\��|�e	
	�C�_���հ'��I�`�O�.>�DdD�Vp�)BI�x-Җv�������	]���jױއ�<JxG���@�'ʕi�2�=񉺐�N�)���U�/\���M���)nzI��BGӝ�7ߊ������:��zK�QN"��v�h9�������;z@�q�1��:��}�,� 8|O�f��qu�%I����ٗc\��\�p��7�u�7��{�<T�W����.�bX� �#�8���R����Vz��Yn��ɯ1��_�8����s���ysvt�������]ʁ��^��Ǹ`o���s�滊z�ԀyĄ�Y�UɅu�������}E5��-�)�[�^��H2�l53����?���%��G>�;�F�э�*��g���9��v+~:�Z>���S���Le�����Q��#�o�bY���#���{��Su�2�H6���C������l}7�-�:����Cd��KTlj3
���sV�p	 A���=܅���ZF�n�l�!����0��`6�~�p�GRc+R.��/�-�7��U���X�e�_��C�?�L�j|;Fƣģ��;�Y��q���=�h�&B�;*����JC&��4�<��\�ܴ�*ҩ��΂-����9+��e���DW���H�e��k�X��ވ���L���y�6`0ԟqoS���3��d�MתHx�>=�u9mI���d	�bV���� ��ь��Y�
=�$�h�ࡽ�Г!q�����������Z�1LL]��
��7H���-W��,��7�Ѩ�捻�=����������)���c/g�U6x"�-O�e�76��p帟��ho*��x
���)�� ��;�$�Oc}�r�]y��3M�m$`<�1d탘Y��<� .�;�����@)^z�Th�B ,ü)��V���m��8���ĳ�٦�<�U�2�*��e�9~�b̸�Y��:��S@Ա)���5����뿘_hP���"�����-
[���2,62AGtTF���pӔ8U�e�y�����b�x����Hci�G�(	a~���e[,�ݾ.$�	�	g�������l�DC�֚���C#&��ԏ�]&���]"_��}�x �.i�9��J˷��R{��|7�#�Xi�9���w�lfst��|ؙPr���ۄQn�incR�j���_����ְ�Ba����lo*Rb�Hp�O4����+4�a�ϲAջ�@�@m��?o����|���-	�!Aw���� �뻖������ƚF��ȋ��U5�+�;�bk��I��y�z(�E�lN��ݨ�*_I��b�ׂU�Z�_�%qny�L�f�.�O 7L���N������Ȩ��[����_���'�z�Q��8c}�e��.�9���+VDS[��V��\��P+ ٙ�1��>mA}�
]󣤲l�L��#���N ���]0�2G>4ݭz�j��Ao�~,�$��_�w,Rx(���--�0�=v&aSq:fS�꭮༞�]��d8A��#����oKmQcA4�� ��0��`��N�@<�%����u�a��$[�c+�<��e��JrԨ���hC�AY$FH�G{C�1;�c+̽�I6�|gS�ПVҚrh9�)"�Qcp}	��?73�(gVԉ~�aL��±Z�"�o����x�*0�I9���{���N>���̞��	f����9�i�j����S�0��z�n�:X�-k$���D�M�^xt�S��4��h7��zY��N�S�Q�8��G��b=L���H��UL��������� ����3*0��~z2���9]�+ү���'����P�w�)�=��:/C�Wdep��_�l���{[X�Οuk3n�2$�@��|��dc�'���E�ur�Q ���	�'��3V��f� _gC:�dj���V�`g�>����
1���Q�����s;�g�e�W�e����r�T	s��,'��ᢘ�C�o���Qʒ}j�e���(�A}��M��.�D��'�	�U��Y���'���Lx�V߄��#2�Kc6��O�>^�!��0W����J�0��3~A���}d�S/m;w�7A��fq��\��Ыtі�Kq`��![\ Z�;��K�"����·h���U�Rj����bƞR[89���8F�L�@}��Opg΀����=��?�����@�P��>�-���0d�.��M���-���3i�O�/�E�G�7x>k������Pv&�O�nh;�J�L�M7�)�x�#w*��'M��:�Ž�	Ή�?78�H���sɢ����	�w�ki�ߗ}�4�$h���+8
�����D]�Fm�lHr���2O�}@|����DPkf��D�:&F+u�ԧ,�u�G	��Yʎ��z*���W9q���	�2G3�j��������lH��c����M.� dJ)1�oz��'K�ObK�K��:n�Tٝ��l�D~@~��q�V�rk	Kĭ����}�n��z��$�[v�d�c�r���	�, �W�.��Ӓ�(�a�S��_�7�!�֚sÐP�!�2Mwo�39ށ?4��?U-ò!��#����i�_g_�;��0CL�"���u^Wt��@��i?�2� ��ɯ3$���t����v����Yw0��Z�_ߌ�c��c�v�������R><�F^�-\?���36��HF�
Ix�b���b<�S@�C����t�k�aTZv�>@R;9,F�p�M��tm) �~*~u�b�1����C�'��!��!����C#�W�!�8��_e&߉��d;������GpҦ{.���%4տ/���T��3ex����O�w^ܷ#q�GBO�Q&�gŇ9okl�i�01�tZ�d��J<���>C�߻c=8�91�/f0���qG/?�S�e)Urv�O�G0��'��֪�^�\��r�/c�9hC�
Y�2}?��)<k�N��)�;w�P���J�F�XV�_g�o7�CB<�+�'/�F�����,ܜVvJ�M��>(�O�)����3��C�ttΫ�t�)��E�v�!�ay[Ȑ݄k4.�ͪ�/�������Ƒ��@� ��`	S�����_����u�:��<w �K[j�v���NN��-�����0�Iw�DŬ��\���Fm��	x�wB��V��w��#����KV�PQc��`���5�6��
�[�[X���m���с�����7���E6��[������;ԟ�M7�g٠+��J�L d��j9A��S��o"��R`�zp�H�9V�[U9�ނh�.>Sv�aE��{,Y�����1��~�O������>����1�;�q(�5���p:Ip������:>����^R��"���
�^�1ѳ��{��U�,���F�uhb��"�΂,ދ��,]Q4pq����/	`s{!b�(_#�4ԕ�����0���E��|���,���`��Uݛ*���qs��o�� d��ur��Ar>"�n�NH�}�ql�Ї� y�:{x�����ˋ(��J�D4�b_&gS5;��.����N�;)�S��w�?>�\������!CK��b��<��������s+*����f��a7���X_Z	��)6�7֜|nc5wKu�v�o��i{{{f�:�ۚ�7�r�p�ujI^
�.�qkد)Ɐ�J:�:�4槩(�"v�%}��t������ZI�Qg/� Z �b������qSQ۾C@q�(��R��m�����|�R�P����z��e��=��T�$6�"�����x�=B�����(|+l�
#s�CX]�I	��ҥ$��<������q4gx������E�K�{̵�R����z�F��-!��.�� ���r�u��hO/r��Ӄ'�"ŀ���(�W�4K��$݇ŋZD�xN���
ߔ�zK3��#�f�q����=�lP�\n�-�=S �u}i�,�����$F2Vnk��a�0�%�=g*MMC��[��7g)�,
��Q�7��:$��j�4�����ys��B���6x���w�@��ם�������
�0sw]͡2Żmv%�|�7[D�^�/�y\��UW��R��6	vb�e�>�:�D1�^,=�bkқٯ�E�	bI��!�M{A���}���@�uY�cy�?6�1|9)�V!r��V(�aA��K44�~���Dz��X�#I�X�0R�J���S�V-}�=P���r���]�c�3��a#�e�����D̶ƪ�7ލ��9���\;�8,�<�A������F]�\��� j)����J ��5�+�#|�C��\��'��,�}��ޣBHѓ�:��RӡK��3l%�1(��x���o���zuѦ�J���WΆ�a���"��N��CY��C�1�!�г�>^'��)���S���W>��/s�yqהOY�DsL8?�è�-%��q��l^���<�an�@-����E��P*΁ܐ���&�~��UŘ
�DS��U���m���[r֍i݅�oC�(1t	=AL��U���T��Q�$h'��W�r��(��5a i.φ��*%����#wl�����tqm�V�n��x�����i��$���4t�a�^U��.��d'��_@^��q�i�q�go	Z����-�}� BA/������_�_V��!&z�?Yg�?�(�T���8/��m�I0�oڄ7��9vS?��i}m ���@����;J��,eߖ��?KxfY������u���/�:�T���t4�e�b_�Ĵ$�}����̓ :��AY�m�F]<�+��|�N��P"|���B�t�͙1����ۀ:�Q=D��V��X�Vޝ��eWiMF/k����8�QWU��}�*J͵�p:C:\&�=��؄D�����r��X�0��T�M�?}I�ձ�jj�������_�a�^u���9�݃��B�P��>-{RLBݗ�"�QW�7��H��z�~��@�>�ķ��|�?�ʣ���&B�� l�ãZ�UI�E�$��W`��a
�aS�WX!5߃�y�_Y���~�l�̮@ZSc�J���I?��/')[��>�I�G%MK��j��(�꽑h�!������nw�:�����Ȼ�``��I���Q�}�Ib n��s�`�ƕ�)ױ˹��"��L�!���~:���m`��RN6�V���`Ɣ���H~kl/�gj�o��(�	����65�`�Y��i����AV�	YC�"�J�A�����?��Q�C�4^���g�d�rދ�p����hԙ#��a�,����H8��5iߥiG�@_�G���M-��lO��
;؆��-}���k��Z�����D7�RHksq�r�.(��N˄����z�K�o��e;���&���.Ҍl��t�k��$-�n�fit�y�KHh	%Z�2��sy��^סd��VW;��0������W9s��ą����ބ �2�7l��}���{ÑĖ|�m%8��?(v�����V)	�`f��ew����o5@{�B/I�(�����N�>�~�̳N�[w�����6~Z$�$$�%�1J�����̂�2P�F�,50��7Ӳ�i�[o�^�f��z��.U�w��DIˍ:�� NKu�$���ƶ�N���1�;"�l٫�ۋB�SHggN��M�ci��LeJ��nA��n�{�$HGU[�xL��#�D�NZ��lQ^�l�rz6��5/I���]W��h��̕2,u�/9�\����b�B�ֱ��0o��Z��r'W\�x�=/#���A�G��N�c�}�DaX�Q��_�TSb8<>��w�kM'��洞�6��ZS�<��$��7ԴW��_�U��r�~j�e�$�� 9]�u�Y�d�F�:��*8���#��8����%��t��G�*z�����dQ�0��f�R�k>�1$�
	��!ze�.�Z�|\&��Ƣ��KT:)F� pWFN���[sBf]��(� a�����L�*�&�5�K�y'*���P3Z����d�y~��J���ya�e?�|�����*PIO�1��f��@:ˁ�C!u����9�bI�v����&��-c7���/�
��Bhd��&�3��)B����%6��컞Oe���hs�z��o�:���r w��2�,�5q�?��3?Z�c��2XEh����cfZ�/7RkJ:A���"Ϣb;�Gƈ����\���� =�8k��/v��2�������@D���w��iv�도�АP���]x���	��'�<	!!=�����:�VB5�q�tމ�Ua���������iG���z�(�(H�3?�������N)����E*i�
.<���@g�ɚdz�!�|sC���0���(���!�ȟ?�n�O�Ƙ#D2�+�j1~3m�w@pOƽ�����Ȣ��䈨^����PO���tE\��wB��a.�ע��z�x~�-��Ĝ,�g�O$C�m�U��� �H)��Ϗ@���|쾜��A�s{X�b��y���¡ u,B�s~��N��e�o׶.A�x��(GTWZ����si.�i/��n��������X�qr��}� ��b�#VKB�Q7*{	�@Q�Uo�\�\[w��>�s�Ytc�Ug��/ω��-Z���L<5,����0t�3.�6B��un��4�`(�;���iIՐ䁡���5u�wO$�)����x�������V�����>a�D��#��[	����5��+|����@ԫ��7�,U�n����8�s(:���Z���'⮚kWH�f(�J<�x/I�S�o��U��q70�t�A�������0觑�&���SB���6=�q� �9�p�6C91e��?����'~���R���؎��g� 9NM���/SE��{Dn[([{%�M�+��Y% ������p��̟������*��|�[����]R)��2�M^q�qV��m��R�:��*��DP�!F$O8{8� t��5P4�]��߁��ZN�����O�;���ׁ6�uZ��+4�����!Q�F��c�n��g���$a`�<��^ז#����rP%#[�ء�}��ձ/�_k��4^���B�B6СW����rA�g�Ug�C�����
|�/�?I���Ы�ˍ�h�8N~�)<���j,��u���9Y3� yc�ۓ���8������4�*$g���oE1_U�Ty��J�*�F��(?��Ƨ���nU����Kx @;�M�{�?����x�.��r�*c�D{�G�ć�����H�;��C�Wo  9?��v�y��w�Noo��s={7𲯋�z������G
$�{XԔ"�=�ͱ�\�OK�V��f�T��n�[?N��~Q����$E-/��%n��]��nV ��ē��Xo���H����4��t��36!0b���4(�S�?ʣ�;=������{lCZ��֐��wV���"��d�d��都U�a�s�p�8�٧�{F�"�y9�"[�c��3W��N�u2�`�!���7C��q~v9-|Du��di��e�P}�/�r�gQZ��Q>ژ�0���<35����g�@���.o �L(�yM��mS8vve�c[:�������W��,��V��F���4C�;������Q��g&�#f���D8޿o`6��,wWs���ٓg�l�Q�G�<P���钡��$^T4�f�#}��R�K��,��3P�D�^��[�hKwʷ�&�TJScNx�D�le_A�(S(�M�Y U� �8�ƈ�_�=�.���������7�Y��У'))�dV�r��L3�����sc�6�@�fq��+G$�[s�nɟ��'u��t�ۅ��a�"�8��Q�Y侔m��_:�c0j=L�\	d��Ê�B��$"��v�._�J�-���ٌ�,	@-Г���3nH�a�(Te�m����\������G����-G�=���$����d�~þ��R/��y�
���s�'M"���Y�r� *�8�l��|�!�e~�"X� ���u\o5�܁���P�R��[�9wkЅJ#�oAߌ�|U�ͽ+>�MLP��WؚDѢ�z\N�	14ZH����:`����/���'H��� H� �(�-dh�!�
}���q�����'�D��&?��:��?���zN��M�["��ĭh�4�z4|}ϱ�xp�c�M:bN��'�����]5t|�����40y��t��\Pq_�W�JF�$�8��ыʉX�%�B29PbU�(���^�P}qX�#}�>��S��9W��3�E�����]�࠹�\	s�T\V8mWn�R�юv�ɘB�����QCl^g.��s�-�֋>�|³�>��"���)�#�c����/���1�,�p�"��Y�-���	.��8p�0��~�]���JK5���Y�h~��h���"ýg�v	��j�{��u.:P����[Aؾ�O�7"�4"��cz3`ny@�o ���uɘ�%��F��"�F���&tI��"� �pP���_���na륁�i�K���`������Gz���;m�F�:`O��m]��l��G�;	��Ѩ��F˹�$���3&�gZ49��$�=�]�s"@,G��� �q�G>;O*#e~2ƫ4#�d�E0[x"&�P��؂[VFԑ�~��O�B��.W)��������z��%Ja���X3;���U������J��ZTš�m�{�-pDBuYҲdYj�Sq���'���$!��q.�᪋_b���eJ�e�j�����~� ܝlb�)�m/�r�OXb�J 6Oؙ����A�ҵ��e�2�cd�5F�iI�ASl
^��|�I=�y��X�r����Gɀ�5��(����t`���zpNj�a*�5�09�>�.��-Sp�<���gr��*sL?,���Bl�|��k}n��xi�<8��A���F \�g�:�����:zzz)ntq�.��}}��U`Z�G���L�����%��T�O.fᚘ-����Ϣ�`�\	�E=���t$�C�~LM�	���������Q���A�:��/�����µ���4s,�IֹR|1>4]1��[_�Q{ׁܑ�Ϻ�7�d���'��D�|+pj��k�ʮ�2��s4 qF�Tm�;��3��0�wi!��p��M�ci�>�K�~��F�0�RK���V�W�B9����n��yP��	��i7؜�Hk�����8ڱJ�&�I�L����PtJ�t��p�< ?���|t��N(��`��)v�q	����
�͑�Ki�w�&i�&�&B'�z}� N�����X@5T������K]a�:�|�&��Rw16 F'`���U��׾b�39�A�%�`���r%�a� �ϔ�-�����蠪4q��L��P���� ׹z
��5=�����b�\Q�������h�6:�a�~�d����PU��ߛ�s`�O����}���9r:��?ۏ:�1��u�P���$v�>�]ޝ�+�����~k�e�s]�@���>�����,�XV.����2�c_�5y:[�,|*C�M�r,
�U=���SQi&��CB@h4j��-e��^'��:�./�>����cy��S�sBY��cN[e�l�|�ӳ"�\,�m$�N=QC긐���H�[��^,�Ϛ�'�?񾞌G[t:����	�/m/���q�4~))����%�<qu�/����|bМ�e�+���
Q��jS�;l�[<��GK�w��>��K���޵��?.8��{��^U��й�j;v�������3�f��h-֪�<wٹ��2J�)���+Jted@��<�o�ӵ�C��H?)tGLg��۫��w�=�%Ɵ�;��"��[��0�d��U+�X�f���up��+Ҷ^-Y%��3�̦�)��@r������hG�?��d�0Qt�9���>���B��塀��n����UH'4(*`�#:�~z��u��[a��_���1����n��EK�n.f1DfM��Q��z[�Y�m��'dWq	�u���3,��оA�f�����D̿d�,7���h�[I��?��r���le��VNpg�>��sJЖ�s]�H���:�#n/���Ǡ�>�ScZ�R!�=���P��h�o��y�����j�}so�w(�I�A���T��)���{�J����G�(�A�ڥ	�3����"V^[�I�̅��.����X�J^sI9���!S���T]�O�0u��#�&��mp���P�i՛ͮNj��A�!T�{[�]|t��!�ϟ<�Ч���cp�����2�b2�V�V
9�bǻ	�W�U4��\��w�4�Aj
:�Vs(��.%�_�l��$A��鹸�c������o�wʎ��G�g79q�ӭs�$=%�v����T
�ց��2	w�/U�Ԃ�R��ꘙ��[��!y�`Eǟ�zi^��n� .G�%�R'�I+��yem�p2�:���5�k$V`-����k�exg6��.b��C��u:�����!�ea���j�����5���d~��*ɗ�HKB�7ɒ��)��G��x�����d������X^���{R`�@V�onԁ᱖���m��0�=��1..d�Q�����%�7�M�]���SBB'[�*%8���uO�amo�j**�+�DG�rQ�+8��٢��[���l�6н�Y�S���R.�C�kQŹg����ࢁ���> ѳ�q��Fp�g���+z\�
�n(6���j�d�x;�6A�i���3hZ������E	��9�/�L�gvv�ĶݍN��c�j�F��ß�I5I���S	��pt��Kw����U���������,�V�#�~�%`�b<7vv2)xʩ�7|L?�y�k�+;�R�*?h@P��)�8�g܆B��Hk��p施w�)�����}����vy�c:	��w�����ς����J��u)�p��h����OHG��f�s��������~���'�{��p�V� #BQ��X�����X�e��� g4�p�>!���OBY�T�M���T�;���$
:�|e��c���m���T$8Loܸ!Q_������E^���K�C���ݘ��Q�����S)u��c��C��^/H�	7�nM$8�� �_�qA��g1�﨓��&�w��=􎲽K�F k+)'��{	A���-\v{�n�S��c58��"����Nˌ���aՙ-���6r���$9`i��TV��J��)vM��8呂Z,�����{����\�xu��P&�|����/z�e0yіY��:���>%���g9݆p��u"��VwX���1J����Q����1~k"�����]L&c!W��	���i	��0��*q���n��B�E| ;l�2	Rd�� �~w��+e�=�v�/�}�i�g�w����X�R
�Lt��lJ:��U���k7ۗE;���^5������p��c02K�=�C� E�R�h�{��f����T}�+�Z�?�ۺ�/X�w��	l"f[�Ӊ:H\�.��-�����N����J��S����]�)��"�1M�h庒��p��	1h���4�O�����YY��}Q�[�{�X���s�}�V���,Ol�n�٣�����?�U��4)��6�x�K7��<נm����$�/1	�0~uı;����ᆐ8RW='���>j��[�w	�P�q�0���,�����lB���
+�oa��A�����ϥ�Ț���~�2���m�:�m%{`>�L�� #$�/�r��U� m]�����&��t���=�^^缐��}�s�o�P���sg�ݪ����N��P���_��#���Y����S�y �������F��	���*oɉީ@�<��L�|�/%�@�f?����W�����D�Kε�H�\�����&�s�<q/�߈�_+%��5U7K��"���ﭹ2��[{|�kR���PK�� ��/2�Z��P�XL�T{�O��w�>N�]���^��]��dŝ5�x~�������O�п��j�3�k��^�J@E�����w�"�j޴P7Ӫ�"{�ۘ�*��/2��{��� ����&eº��{���F�H>��/��x��R�{��qh����A��XNf ��!�ۚ����~�s6�����@�M��R.��T�ޗI���"n��N��t:k�<ȗ��
>�v Pe�=F�F4���d�t��45��?O���Z��2�վK�hu�%��1��"G�N"�?�`A_ږtR��L��lF����J�H�~}��/�]贁.e�1�G���`I��i�(���sK����G��W�P{�A����b�U�Ňy�hF}�����H�|
0�|�Ls�-3�Q�wyIm��M�ǭ�v�]m#�aT|�X�����4s�Dd���t���bA�o�a%02��Q��hrmS�D�`.��r/�?��6�P5�ƺ%�
eE��'�sP����� F�{�[W>��ut߹�j����k���*칩J�	5�~w���s�:u��t�������#�_�4�^��H�~��>R[�Qgr*���W��	�G��9j�e�>�#�;
�qڶИ{����Qn!V�3-�) ����ů ��=�rC��t�
H1�_}�TS8�^Gޔ|b�ے��� r>���Z�EJ�����th���_�#x���FiC��}@C�ՙM�]�'K4���1��~���K��,'jI��4�Ib�Özvh��)�����ț�li����ފ�l�O��Յ�N�V�aͧ�����*,��Oe���ѱpվs3��7��M��������z�gc���=�B����U�ƺY�3�G*Z�-���)����2��@����G���4��@P:Z��~C��(X5IP"�7aP�{C2��0���z�K�A�?�`j���ٿGy��2����������zgq~�Z�����#F���*�%���W� U��8�SA�Q�{��;��A�rO��Gz��+�2�a�.��{�0�� -CS4�P~��1#-5hQK������F�dEt�kv��2��&�zb���V:� և�H>X�T�6&)��n����q�T�L7O�l��́��K�]|��..�����_����L^���D%�QO�ԑ�;֫���>��)�U�,n2D��`i���^tŒ�FBN2{�f ޕ6[J��mZJ�(��e ��v_�.���x V�"j(6S���Ƣ"�p�; � �>)T-�i�~�$���ꠛi�<-�{��B0eXnQ�*qz7c��㪳#F�k:����ܻ9��"���8�2,����L�%�Q;��{1�ex�@�9'H��F ��[�;4s?'�*|�M��ijP�j&���)���D���<>s�ˮ��b�A⳱��O�+�z�T-G���C�Yd��0a�Ř2-��$��X�8A�b&�A=��l^���4��u��ko�����Dh�{݄d���˸�D����P+�h\��?�'	���U��."^G���2J?B���I��}���-�T��2s��(���yz����/wB(	H����f���B1�4qʸ���2Qa����ھ��>Q�|Z2�Oz�٩	�s���9��d��:��(�9{C�s�����L1|��R9��gv`�a�3+	���|����*u��?�99Y_(_3���h�Y`�G*a�i��.�[8b.�� �#��mK� �giW�{w�*��.�[�8e�8eϪ�>��JZ���J��"|�'+�.�c ^y�h�0OI��ݏ6ᓏ۪���I9�?\Vn���E"�o<ڎ�O���@�������a���b&f�T��76^���mPI̢�qʤ@X������I�u �S�����Ik8�t�؈�J9/#]N�QL��g��{��Q��������Vj�NT��k��}*�v�1��wٍ���W�~��Rog�)t��{��M*��}�k�h����t���c�<�hw�|����&��R�+��2�Ƀ�ern����{VC�3�	�f�\��î��5"eR6#鋓�h-�^��]{��Is�ٿ�V�l�5��$ub���/�E^�7!Khjs#P��s���o�%�2k2:>�mRu�8J��^REldRO�f�b���7�(w>f%i+��,��g��,�b��؄��Y�W~E��֧�(8�kw(��EU��3Q�bSF-Z�/3�`'����K瀝 j����־�V|<�N������x�ƤukJ�k�B6��"�Qa/rشɼ���O�\8����R�B�^�f;X*��I�7'�� poӽ�r��?�n�W]��/�S�ܪ.�-�S�ߵ� ������T�����:��ak��r�j���:�k�]֖�hpcW�g�0�0uyC��󮅯�+5E�x��#�4�k`�D�zt~"�Jҭ�/LrJ�f��s�|��+�`������� F7]"�� Q��%��s��Sb�+6����q_����m�Y�e�O���#$�hf�;�ewr�в`��G;|�����Fn���4��(��	��?L@Zc�r���Q�>+C%�LhB"d.���ò`{��yؠm����+������eF�37���p�;��o��=�b�[`LWX-Pݖ���8d'�Ap�q��/��
˘ᗲr`=zLb"��(х4l�7�Z��CO2�Ҳ\�������4��m�.��>���##S�Ut�&��y��X������H�[Y9��?�T����)�]6C�����5L�����&�p�([O��y���e,�$oz@��ۦ.95�b��;�`w�:����ȥBjL�sw꼈�.:��j�q�<�*��f�{e�a���3��Ӓ �h)r/6S �~t�G�59L�cl��?��uV�ȳ����S�4d\�V����������v�E}1��^�i�%�w�S߮��9p���˹�����YqO��h�j�b�P�8�~�,����*}������ڰf
a��(?*.���,���$����ˆ6l��!�����򫦜�EAu�@}��|Kc�氓����6b�f7FW&ІC촵�jC'�����/fQ�s� WNѭ~l��S��"��h�͝d}�Mr���v�5v%13P����rp$�2�	"�Ƌ��3�G�M��z��X���D_+#8iU�yӔ�S�p۳�#�$�(�]��0�p���,�h���R��V<�̈��Yz��wGi���E��KGf�Л���6�>�ӡ�il��\R�u�ҕ ��0 ���r�?Ё������_�:=��[~�tL��ܴ������e
^&]pu�(X��Y��1�u;\�,��	˹YE�8Q_,?Y���
��۽����0�#ďV�2E�L_��#K%;4uI��6OQ���Cl��íY�]p���1lSc�ri)��+Yh y��낟�*�n������[r|y��>�L��M�~�x�Y1�J@�j@�᱓I�xe�b0�,K[�-|��jr�+��ai3f[�U�Q��{�fPI�MV2r��������;$��|[nOGG�I�X<k\U��	�-Q��0��%H��gs�١i`?5Ȳ�\QyA�i�������S�+�z�(i���F8� A���=m;Lh�����H�������T5��ys����q��i�[���<x�m)��n�< �c��O&*&�^)gݾ��HwNE���tm��i����	 6����'�Ja��]Q��s�6�Mn��P���@̢a�n��.��Ɣ>����O)#�]��n�xi�b͌U�Z��/�w��^�A�U�4�I
mwB��A�0��A�%��1|�,�Y&�>�Z�N���ce����Q�Ƶj��ʽ�07#����'����J�Lt��8ࠋ����T���ZP�H45���\e�d�a�,���u��y3�.��B��kӅ����wW4]��ű�Ae�PV/��$Ҵ&@,{�b���1��+2P	�E�{����� 8y��b�e�6SV�YY��SN�]��� �TP�үĿ�/�.�qҙ~�-��g�)y��n�v@�}�%s7�~��qɜ����e4�L^H�|S�bN0r�r&Z����D5�3��3�r��ּ��1p�D�=��܄��4�k8fN�3�S��'�����@�}����W�`�L���	�^?1"�i��E�?�w�Mw�r>�Nœ<*�$�)X/0z]?3���K�7�Ԣ������/�{�m+}�`t����+���j��Þ�r��i�%��m�ʙ	�N�D��22�7΍'�p�/x��8�eb����;�؀"����{��3��s)� ��9>�G�KD$<���k`�1�����맚ca�A=L�0��`/ފ���ў�Eg�'|�S��V�pn��B`�����f��I�nF�x�����x�5a�P��G���-��ͦ蹈�:j�:�4��k[,�����m ������z>&�Y�[WQ;c�N�I�Ən��Pi^�C;-ݣ�]��#ڎgP��yo>��	4��q�,�E���U��7�Gފ��(�o���?T��ɳrb~%��H�w�S1@���A"�g@��
�����8�x�uo3*;��|�W�0�N�]ʔ���	���N��AK�@G@g,���\��ِ��sz���WP���\��WZ���9ۊ���5,���Hs6�,��C\/8l-�p!�G�!�-�J�)#�MS,%���؋��jB���\��|��֜�����o�]|�Q_�Qy�r�v��hh��V�����B�|ZM*哅�=4Rְމ'l�uapma��ڣ�λ�n�z�C$s��T��P�_� �$��q�P�nu�~�mP�T�Z�3<l� / ��
7W�N�=%�L�Ϛi�n���(�6�x�,&�kH��s��q���􃋗���PA���`�ඣ_N�P���x�M�s�1��v!��6ڂ��B2�;�:�Wc9:�{�1��� �]��O��L�'1i��Ә�#U#��YY�]��<m�۸��}���d�g�5�;��^HJ����:��4���5.�В��_�rd@Qy��WPѓs�S(�2�풷
�I���w~��w�����K.Vo�� �T�M+680�gФ��jMr\��-����!v�bev;����Hz�rt�t�8�X_j�ik��(I�����m�9켯Ħ���w8`@�V��{h)��o j^��.a2p3	�?:8:v)Z���#��eXˣi�6�'q.���#��H06�qPy��F���F8�YF�M���R����mI�iS�S�r�Gb��0��Ƈ��4'S����ș(�J����|2`$-ج�L��ܼvf�F�N�ɗ9��^�ύ�@�]Z?`b���=�n�����Zr5���W����O�LÅ��%E�B'u�Ȕkm*�;��ٹ�ۏ~8ψ@@��ᦿ�|F*^'�-���Y���0HEX�F����tH�*�Ԙ⮪
=���C��0�[�@�3HB�~=ፍL����0�	�l�|:���d��V�����.��!-݈��D�Htn�f�4_����������n���gI�8������̇��TYj.����$4������$���|��hYR�N�~�2t����:b���ߤnav��4:�&��2�-����
�U�_ �C�bG��
��C��.`'���%��Yb<cD��V.�ĿV�,�k�:W���[�$H���R�t�GX.j���@ΉLS���ƕ�����:1�P¾B��9��"^)`�,�f�+p9��z�5��շ$Ǌ� �����!'Ih
����r��M�IhB��;�	���}��&�	�g,�����T�����C|l�>:�d��b�:�?F�.�2�� @jP�ս���2\f���l�::�<��g�R	�������	��� ��	��Ԕ6BWq��ϥ��W��ʖ,M�A�9�|��cI0����?�&������ACY���{�mb�7�a�����H�����`�2-HV&F4���B��2h:+��[�S�Z�Sb�i���Ѣ�S��r�0�dg7��|���!���=.я�ɀ'\QM��s�D�b�)��|C*�`z��7H1ҳ�j�
݃gF�����	��gf+7�5o2L���kf5��0ŕv�P��uA������4�%"���T�",!������(\��g]�p�򝠎��wyMЪ J�N��K蜄9��W�?x�Y2��E����-�+w�I>���N��5Pa��G����V}��h��.��b�d� ���W��#�e�<j�f��}%1g�kQ3۔�nB�gYŶYE��q�ϫ��HE=��e~�u�N��	��/eDD�c��'V��֥ICJ�~�d���'����uΟ�	���=!v��㰷^ތ�\\�ُ'}am�VUI�Aq�vv���:7����R���Io�{wT���[��4�b���%#&�
�8���2�zo�4;�R��J����\>$�����|U+'��H��;�o�*��9��MhGyzLƖ������8�)���?�|�e6�M):��R��R�@�|�Wl�����EC���j�I��7�|�*d �����)*}3~t�{q)?#@N5��Q��9.�=V�;���n0UM)��~?�fPֵ/B�7���ʝ��Q�bY��}��`�,*5���)_`� Ӭ���0�8:J�N��G�D���h����8ѐm���tXo&��..~����3(�Ϙ�)x6�=�.��w�w�q��%���m�����ym����З�_}��8vÝ�q��\��r˞�3@�W�ח��y�(��l8�gZMbo)��A!l�2���L�$*�@��#o���w���%��&i��0����Q4fI��G-
�~�5&CfE��	�w���8-.&r��c�5��/��6/�\pa�\_��P�t
��{����D�=�V��S��8nh������[��ѝw�S�"jEoR��v�,ń��F^��dc��tq����ʝ�(�l'����4��+dN�����'@�(�m��"�����6�t�is����0v���[��~H,���@&/=)K�Z�����:���yF
���.R�l*G~R5�wG��v�M��U+X�;���=��i���|�]��?ˤf��apa�&R�Ra��k.�����$�-��T��>�&hO�jZ�͈ksox����������G��7Mן��_����c9���&�a�(�s�����Դjl|�&�ɒ�y�{�?X���w�@T��0$V���J�w|
�h��
�B��}� R�hV} �"�"���'��;v⧪d蚞/�6��a�h�j�L���E�]R�y�]"\E�P/3=K:�_g��n���	�{aq�[�"�:`�)�>�!}���~�t��qm����T���v�|Z)�J���j��HuKr��S���A����i��[�+6,�u6`Hi��X�� su�ܔԅl�������^���.Q�|2��a�y|�San��$�2e�eG!����T��M�'ӵF��&!�-�C���s�Pw'�o�G�˲�W��4��*NL+>��p>���LϽ�\\m&8��,�]fV�y"���$:�1ou���U_o�A����������	L��8����4i�G�|�e�ў&ͱ9�'J�����v�_&��}U�*8��qyDf(�_��=~����0���>fn��8�u�6��f�"sl�d�ű�~��>}��N�c�.̑�o�գ0�8������y����};yq�Ӫ���v�x�ћ��H�d^P6��O0&����ڈ$r���W¹��#ښ��s���vE�ӑ���%�~�v:�4����}�X�$���S�8���� n1�?��X�RD�4�����>�vA��j/��6����Y'�O�[+(��kn����O8��a���h�`�����=AdE�yA�i׃�VA=�f����6[�~�����C�(~���W74i��:^�6�Jr���o�
�Ca]P+�d��^� x��C�/̧Ǜ俐������+�x�Ai��,�|-/MS��awd5��zqE���3e�P��B�!��bUo5UbІ~��H��a`��&���d� JP(�hqA�1� X�(ڌ̮�FК��WnSh�4�+$�X"�Y�
�&��a�otk7�9�JIĄ�,{�r��k�=�ޠmm�zD�f~P��$	L{3��Dݤ��oU־<VD VQ#b�r��"(3�)\s{�#L0���ca��x�EsD�shn���W���{��a�E��3�u��XCv��D���z<����$v�����k�$����3�O�E��jmhM��<�yk��c��ژJ!�szl0���4�0M��v��M�Kzò�e��g�0UD�c
�gGSA3��g���".��J�?����� �l�%�퉄E�u_{������t1��u&6�/�����7�U~6b՚�L�� �[-6�A���Qn�6 Ժ;䗯^a�$b��Yw<e`�Y]��[�;d�O4��s"�]Q�VјAaK�y|E�j�[��_�<4�5�g�K��櫕
q!��ܕ��1�����
��.r{!5`�qĹa�equX�z�G ��y?GTA�y|���ml��c-�F��+�[B�yB�,�v��7*�f�^H|�s�1�8���X�z�����fA��P�����,C��%�!)�M�����#r��,�F�qP	�I�<�Z�3N�Zl_#��4=貍�b`k���'wQ���[���T�o��9ŏQ;
�����Ҝ��R�?)���˰�xȣ�����x���k���9Zr܆��dR�!�آ!yw{:��2���ut�k��nx�q��b�W(�G�N;��:\�m�����o�C�<]`�h�zV&&���Q$82�)���s�+���^v���,g&��aF��A�X����j�K�ن�!g�5�u���-
�Y���F����ݣ��'��׮%�ǃ�eU4�:��e�U{yܱ��mL� �O�&�	�L�nG5�r�� ����F��S�R`��K�*�YL������u��J�&q�#�{^hH����]]V2�:�Ƌo��1�����2���W��|�-pԘ#�8�ޚ�k�<�Y���^���K騨��Q��=�)��S�����J���9�fM�-K���Sŷ N�̍��**��ֻV�ˉ�O��F6TA��m\{A�E�d�X{�l���Ex���@9��M�#j��:�.b� ��n�|��l��Ml�x1��ﰶLk�ЮS_��٢й�e�g�}�}�`M��fY�o8=��la��n�����ҥ<�3�g��OMj)����CJ�i�?`���5	z�k��oUD�ں:��e4L�s�K�c -) ��J,��GF��GP?���J�E��Fu� ���fhY	����h��l-�T���y�O���մ��Y��GΏa�����T/"R�r�羦;TKv.C���u�m���e2D�f|�֟���q�#9�����/(�v,��{2�ha�Gs��y�J���`!�G ����v��$[��N<�� ���+|5H�g�]���<j���:0��S!�R�(���Q�y��#��px�I��,W����j��4�LZ�D�	o8F�Q����mL���_$�~���@}5�z3G+6�V�5l����<ܮ@K�5Gh�
�����{�TW��m}�=��YE��a����7�����\���(��p3<7)�D����	GiA�ɽ^�iNB��2��W_���-��E�����޲K��l���,9��}A��&�O�9ѫ��h�ʆ5����O1����d��lD�h��M�\��MJ�N�|�od��_������M6�EY#)>�}*�7�伫8��yB-�"��%�P�t�>QP0��?*W�0h���z�I�hˏ29LK%�ѻ�x��ھ�U2�ߙ���B��H�r�O��ỷ��lEF:�z���,�'��
X�r�"��n���;��ص9��#@f��$�U��R ��+���ͳ��X��A)ʖ5�s��>�[��I,��M�~6~ȡը�X_!�L��	iG�>���(�lr��zO�s,�w@N���`}���������S|�>Cf��I��)�-ωaڊ�����Gg��#@f�Ho��c�~-&,h�x��)�&k5���
5��`�D��FG�i�5�G�CvMxx��Q&:���q���#NL�w������	MDnd4����!�?`��>.%�l�7�]ބ_}E��D�S͢A*�[�������4��}�4�`1�j�~1�|*��q׹cI�)�nʬdf��AY���V�d����m�-dUo�=L
��� 2+���I�3�;T�2~�}3Cړ�$�����mT�!��m���a�V��;�P]Q�*�^��$̆1~��.t!�%C�١���X�:k��*�t!��_��Dϫ���v��o?��5=zD��4���ly�sH-��Z�����O�l
,��d�h=���;*�&vG��$߅18��[?<�GQ�7�o� E�:��� ���I����N���ˬ!WAe�l���7X������O����=��o@M��Ћj�<T�j>*A���4a�	
p�A�	j����p���u	
�Ϋ]݇�˪ ��D6��D�vlJ��"6@�����WO�·�X��Ӵ��^ܿ�b��﹏����[�9�"�4?L=S�;�jl�ۑ�]?:�)0)���ϳ�����-{�����y���x��#C;����R'ݩU��dI6&�	Yo���/[,��۰K�y� �J�b���п�,��-A��^���.F�U,�ֿL�<��!����FV�=�"S�q����V2&�G�s�'h�BX����Qw� ��̀�4�b���Xx�tƓ�G ��k���(�c��Ck�2!i�3v��"I6kQ/���;cOGQo[)Z��a��I��J��i�{_*P��V�W�qO!�O�D*��@� ��uRr��z{֯�54�#0�J�đh���ɖm�GFڑ�y�]�~�e��d��2m3x3��������K�EZG���$z�M���wk�S������s�|\֧�.��pR��-k۔��;�uG����֟�ӂ�K�g]@����\����mq�t��Kߒ�q��=I�1D�A#�r��sѫ�^&"��d'�/��<�oG4܎D�T�?�<��4mi([��GL�pU?� �R�eXh���b/a[<՞ {����'{�X�@�?���IZ�S�����C�~N���@#�9h^�_c�W����3I�Tp�.ݫ�@��T���A�l�����/��lu;��<�4)vV�H�[eE�$�l��N��]�N�:�
5ۋ���'~6uH�����Y�X����n�?H�O�8���=Y`�Ժ@H}�/\��~1�*� +�cs�<���`�q�T	1x�-���̷��I�wvEe�^����WLHI5�������0*�p�|�nŦ����\v4�!q�oʱo��$��d��
�t��t��L��h�_�X��p�gr4䫘:(qij�	#��/�ՉDEw-�T�unCL��1��d�Rw�DBr4[���i�,2"�&Unfe��:к"WY�^�j�5����ps�<��o9A��y�vSBs�b�ؒa�3l[�g=�#��2~��^%��~�떣��eе:+[��2���A�G�b�^����t��c8E����ɮ�F,��� E���˨_��=b�[#�[�e2�O'TL���^���rQ��
'p<�[����c/��}p�J'uT�b2�����U�xPm��qP�^y����=E�bC��N�	������]l\���$&;�8'^�ˢ�l�n/(����M���AEVa����8Z��0~܏aEA����4�v�7�����Z_�0�	fM3e��ZD��{8�p,�d�>*��ۦ2�+П>sb '3�ň5뤸�ov6.�es1��ø��̅�ŀ�,%���������f� T��P�ېx[�Sb��$��,�,��0� -�f��^C�KVm��$�ۇ08wY��Q�N���a݅�T����b���9,썫7S��
ES$�+p�]�nA�\C�����Ӆ���J���gu���û��&� ��ץ�Q:,)0�:[zq�uA��p��	]�����إ�=`6:�'w�i��G]���Ej�����b5DN�nύĿ��й~�d�����<����҃T%兮��ţ0�̂up�[�����s�X�c�z,Л�"BK�R�c�q}4a�U�,�0N�縍�q"�Z��:$d�Z�g3����Ă_�����c��I�ρ ���I:f��L���/��0ܮ�h��0��$�5`�n�H��Q�h'.J �/�����.��`���,T_s�RHO�Z��m>_���As+�_���R��_�9��,c�m�{t�i���Ԟ��-Y<BA�3G��X=�A��+�[�P�v�dJ�nrF���H�s4�� �8���-���g�iv��M��T$*�?��|�#'�}�f�(�����Of8�jyu}�Sr���<_��,8��i-=�m$`��l� ����#���q=�Ⱥ���֨ac�#B\�td1E�0F�Y�p���OR���|��Qّ�\oo���-�ť48?�I|���~�K)��3�(�RY�T��Xe���,���6:+'K'���u�i���X ��������.1��F��z��D�(Vd�A��E3N�٬�wA����?ڦe5��rV��&j6!�X��.���V����,�%?��2�%1����<p�l"Z�f@EEYΗI�fzzZ���N	%���3'�`ա�E3��2�Pt��G���t*��:~`J
��´�3џ��+�t��A�y�]m*ª�Ք��-nk�<6H��a����^@T��4�6�Zl	{�(�����tK�_$e�4�L�f\z��GF�����[ry�����h�ڨ#����S� i�Ł��?��������m;�e�>�d�̍�I����`hÎ���:=���}%N)�S�Z�@|��DߞƤ�h���d�^�u7.�5���䤕LbwƊ(k��e�<|x�?���-?L#B�u��d�Y��7���7�2���k���XN)�El���熳�E�{o���V��0��j�������E�x$��?i�9��DtZ��}0�Y�G(�GrjAЊeG�B��������ӨzX�7�����d�+�P+���ʈ���	���J�aB��/�N&:����B���F}"����Rw3k�`!f ���O�Tl�ҟ���\~�&f�����CÕ����z�*�Y�E������ ������#�,���M�b*8�:�|��J����@�V��f�|�h���7�v.��y����H���d`ޯ�� 1�[����9�9=J-]Q>{ج�
���n�z�=P��Ƿ�˕�*Mk5�-	���u�'� j�un 1�APڒFM�Ruҗ�F��}��!�M�
��<�6r&�I�-q�@IeH���s&�j�+��/{�;��UsK��� �G8��z����xbĘY��7�K�:�V�@p��ح�0�X�&9�\�U�J�����Dը��ѽ�kK<u"<I�״�����$Km�NF o��q�{��y��!9�e����w1��T=�>G���(��I�B�>�K�Rk�s۸νk����)�J�\�P� �[7S�y��d�<�I8�+S>D�Finuy��k��,;�����!qI�X�(����(�_}u����bE!����F�X�����7wGs���%̪�.�Z�#;5�+�Ͻ�w���~�?1��Β��n������C��2Cs�q_��Yp�\P�_jy���6c�,���S([A��t/銝��4g6�I�ic�$O�-�~C�����N������-��E��/�+�x�/O�x�5�a�`���h�<�zu=�����T��qŊc�LA�_RX����;ړ��K8��j�����b
��4��U�sDb�'@K3��Nf�3�"�)\�/���ؑ>�E�8C�-it�`�Q��k}|A���t�~ϰ�'���u	�xEjU��pM��BW����/�y��E�ʎ�Z�h�F	߽|zBJf������pT�i�.��Uih��I�虙�G�En�rN�wʊ}XU�>�'�s.6L��`��	b��ZHq=�0����*N`7����s����SQ��b_�A�UW~q�>!����c	?��|R򀵨��.��� �!1����Nl4�m(��u�b�]3�D7
Y�pL�YP+�g�?m�k5��.�^�x��/��VSJ���o������d��&�!�=��R���J���&b�1�BC�ruȭU�X����ܫ!�_�,:�����4W=د�>D#h��2%��m���.�r�L	�!��W)�KG�!���^��e�9�����YxR��jJ��Ϟ��2؎S�"��ibApp.?�L�d��/��SE�S���8���O����7{[��Zw�T_��A���	�2��W��[�C�M���S��7a�R��etz!�exӄ���Lc����Q����vj�W��r�gڐ/��8��7�ɢ߂�u��R\�����g�"+i�.��\�K7��lc��F�R�8PYe	q�ӄ�t&~��f6aL�S*����(�u�KlaV>J�8�k�%�+�Y[{Z8��n�g�%k6�h�e���J�C4�A1��^���|��l��w�qS����a�}� ��y������0#�g�ߠ��g��U�p/XSV(1D������{��Q:+�X`�}(G���	�ͳc,��X��6L,�#�n�mYŋ�)`iXx��LQ�%�^_�ʝ��8ss$�I�,W���E��R���V��Ч�q쭂��u�x�	�N���iޤ��h�W{D�z��I++]��<c��Eq�Nc��f*��n�}=��N������wk�Irn�d�H߮�Ds5S9�Q}��?}�t�x�z����q�>�y��MaIh{-Ku�G29��F
ۓ݂E��^�ie�GBX��� t#�b	�g��bq�:"�� ��5As:��x��ȥO�K�5U	Eo%�lmny��B3����6�=|�_I4�h��.�T#��>�lBd�ȟ�a���s�v��W��y�*<j��۱���>OM=��9Xn1��Dq�-�pl�Ib\��kMZ��������n�D�������hE�#�q�}#�6�>�e<$�Ը<0�΂b��wT�[=E�;a�~��?���yl�D����뜶V�ku�e�h����ܸ'7�[��
�w�Uї�+
�֭�C�u+^�f��&tҞ����4gBU�n���/+`����
D7=����b�S��kƷ�$��q�%��S^����-�\r��f��9я�c�@��@������{�;�#/qc�1�[�6�S��N��J9S�tf=n,X�_���M�U��^��K�{��sz�S��`Gn�[���e{"w��F��Jz@�d����>�Gƥ'*���ch�ݚ���OS������YX�(�v!T�N���HJ�>�L�cE�4HY�^�𧩘�o�!fALˠDK�g���a���j��r�6^�
"b����݉s�� R|=^k��aM��&l�+�G(�P+S4��Sl+ל4N�υ!䙢b_!�O����"Fٴ��W���?\n�O��<��r�������#��2\��
���i='�d�d�@���	��=� ~�`!�ދ��ʈMn��>19 ��*vVD�@�k��8DUߥ���S�%�%hpD]dlRP	{�=�,����J��Cϩ��W��g�!�lI�u\	0�?S� ����K�g�UX�����u]�*_�n8M�v����I�lr������u0'	�W)��ҭɭ�����W-���qK�x Y޲2<g�`�]�Y�IJ�i��,K���J�⼙���ox�q�N�K'C@t�Q	-zo���md��i�.���W�h%I��j�Y�	s�y��8��:
����A>��X9���/���n���̅�>g�#�De���ֵ7
r"p;.=fT�y��lN_��`M��|��|��iQC4����������OP�b��gJ̭���C�ʻ��z,w9���{H�����u��IW&�2B�"6��d�Q���yI��.�C�?x:���,9=����T�=��^{�X8�$C5��|t�LmJ*"��8�Q,��]��̧�[��h��b��2D۩��Ia�j��/��\�v��,y	,yv,¡��� l�&WD���٩_��d��'��^Df�*�:#�m`Jmpk{89B��&�GFUY�_�ǽ�����YE@�)x�qp�/ae��''�{�?V��.W�f�������=��-��/�:8�(��{�:hoK�O2�w�(+*1q7wHۍ�U�k�Y8va�z'�����,#e�=Sx�ݡ���.�x�z_͡�ྖ�����̬�vsW���q���(>8� 
E���|���E��-���0/;b��0S�0o��gtp��% �vF6��R�
] hQg�S5��+|�	�pw�����4���d	\�o���|0�u����A�G�2kY���rڐ(]�.F�+}ͫ)�RW��Pt8̵͑"���[&�����caF�V��@2u��W�]Re���o��#Q{�<��hH� �6�#��
��(�F�;;�e��vj�Ä%�&�!�啲M������Ԥ�x�'�C��!Z���vN�I"��F�%<K�a����Vu't�p*U۳�R)����ĨIE�3u#��[n��_���a�<��٩=�'�	�W�O�A�� d�����S�c.��Q�:��ׁ�X�V[�Ff�v�M�����TjSQ��ŭ�M�I��v=��hl�A�%c|s�������y������O5��YʙkU.S?��:5C4U��p�Vr����X%GUp[����M?�Cu�=���M2������!z�j!�"D7\G��E-&>"L�iu�O#����)�rg��ƷQ0�;�n����8�77�ɷ��Tzg>�Hp��DkKԎ���$����[��2!o���}_d$���&��mj��a�p�Sz�\�P>�vH�,�Tϥ���V�i�ß2�]�=_kI�x�9��Ũf" #�{������.f�c��`�GjCqtu�v�t<.h���'���*���[S�'�=�1)NJ�F��л��Rr�VX:ѿ��C��>:���v�4."��}7W����V���S&cJhu���x��͆͢�	fVj����
�G��>�j7Õ���O�gB
):r��Dw:�q���ܒ�܊����J@n���pd|��`/��6,-���8��g{���a��SV��������2�᭔A����\l�غ�mS�_���P�%�(�Qb[G�!Va��Q��P@7������P�;�����	�"�1��\.�Q�T��.톘��*+����j}Z������ՍZ����W/��c��q!M���0���0��������FuZ}n�����pJy��3����1:wBh� �ȅ�Zn�{D��ҫ��d��d�\�VI��I��.�R���'��Rv�A���Û�G��Z%�;C~c\	�r[����<��{�M}��Y���M5����1p����������`�mS�c���g�:��"r}>�>�@V�c� �l��>$�y���̱����B,2l^��a�n6���!�䢠�f&rC\E&�������Y�<��Tͥ[r>܋8����H@�w�s����p�:,{���E��H�A�[�g���w��S��:�c��'��hN����>�3�ZC.���TC�s�<X&��)F����K��L���;#N����>J���E���?�	*H}_��k ��5`sK�� 4�>X�F������$�J�!%�gK�@LMaYĻ���0�\�ՋL�W��rhkW\A� �G��j�������,�[HH��� �$a��}o}��X�*����<�Lr��$?��?CSpS*#�h��[퀻�m�w�e%�}�ב�c��(�/n}��ł�0��%��ɥ��$��g ��.�i��7���;}�#��-G��U|ĄIXt�u��Xl�>-E3��B\�X�;B�0j�v��ham����4�����X1�j�#X�W��^�p.i��0l�-|U�����v]���R����&�tࡓp�~�����A�bL�R���H;X�B�.nX�G�Nz��J=�}�Pe"��������{wfFf�*���dx,1G��&��6�#�;j/F�/t(������n�]�d�pcH��Dh0�Z8-�z6@ѩ�U@�s�Q�K�7`����u�ź�/���H��<��ރ�R;���Z�)��W>�<|���_��P�Sr�X��)�s���0�<�l��<��4�l�W�(I�\�}f�L�̮l%<WQ�(w��tWcϬ[����itL�����6�i+��"���Ka�.8�/��m+�ejQLY[ݘ�3���M�ѩ�y��({7�(=�>�ߘ~9����	.�7�A-)��L�q��xa9�"�X. ;_S~ˠ��$v,xB�zmTwa�!nN]A̱���m(�Pf��9*��@�o3j�&���O�v�������5����]�"o_UA: պ|�E�j0�o5ڽRnݐFJ>�+��E"X�eh�0��S��(�/�n����"����d�>oC^�M. �u(A���>M�(��S�{��5���=r���f��M�AC5Ǒ�J�Wϥ�۪�ֶ�<�e��B�a�
hOC2̻'��ѕ�Pgحn�%+�g���;�H�"u�����Q]��f��@��LpS&7��+R|�;� K�!e`!r�S�G�����ϊ���Ǿ� �-*��zn�yH��VħR�|�2��2�C9��K�Ǆ�On��SO�vm�1����a)�c��܀�d!�*�}�#�\�љ�+ln����+�e�X����[[H	�c�NM��,�9���N�B���@�G�{�t(Y)Z�I4T���lW�wr�VeHR(^��8���oB�����;~R����/��q'\Ӓ�W�T\�!�c���$����2*��<�2�����oI0ӼT��ūȖ	Zۙ� �aFw�@"ke�+ A[�E7�ʠd�^�Y^��$��܃kv&L��^Ax�����rRi=3f�z�%+<����=(��8���B�+���T �0��ɠ	���Za���+�%�l=.7�NX�t� ��/�I��Y��W�Sy��B&�HI<WW�Di�C#	��H�vl��K�`a��:cG/��Z��!���ָ��p$.�&��ʲ�վ�~W�3ع;�~��8Ϊ��)o�sV`s�J�E�;�� h��I0)b_?ĩ��Zm�,��e�"JzZv��Z�����3��`eF>���zR�j�wW5ٶ�[࿱X�ˬl����0�|"�Ʈ�K�]ԅֱ��iγ�8$��z�o�r�Y_D�E�st�1��H��%G�V29ta�{�R��;+��8s��0�+IL������'	��-*�����;=�P�;��[y͞B��ͧ��`��W�G`�+`[-ݑ�yF�e�N퀳U��1M�� �F�g"� ���b&��r�� �IXj?ȗQh�"l+��N��G����2U?�U��V��ʈ6Z�3�\BWy!���$r��|���bW�t���+���eB��&L���ve:�a�*�x�Ǜ�B���~7��s��{x�_a���b.|������_����ѹ�wd�o��oPו��}� Ů�u�-��N���r��u�Y^�A��}@�㒱��M���7)��/�J�J�nX�)�u2>��/�����렏3�|Z f��=?l��� ��ȯ�SDy��uס�%6�KQq���U]ĭ���kBϥlý�Q��U�A>r^߀�R�r�K^9��P1�������Ϭ�W@�gH��q� KW\�+�ؿr���ԓ��(4p 1�����m���q��0�ds�fS:���CKW��y�Hm���}�)���l�+�����̜a�1Cbj%r=�Zy<IuŁ+"����on�F"�Զܐ���*��D�$��:�L�Wlt�T����)�jF�
g���1�X߇���<��+k�%�~.�o7���Q�S��Š>Zg�S/Ɯo��uyѲg�/��QM��[�\B���j��D��xӡ9���`7�УI.�)����T�r�톘�E�L0��q�������MѬ$'C��w�K�|�tm���$�'6F����g.��1�<��sgF����͊�{�,2������Z�~�\�2&{:	���@��D�ʭI���v�}WaW�j�*�>�ƞS�δC�Q�1l�����k9��$�\��+M0ob�|Q��&	ϧ>�m�1��UGΔ�����-��2?ǅq$|L�H�PK!,�������m+�[Mm�P�w�ٌg�_�����C�?O�٩�"�����2$y�������o�i�������Hka�wQ,ҹ�2g����J`w]H6�)�
d�K�^���.�].D��UH��Ӟ��[�h*�U�1P�*@��o���Ex^�����\�"�Ϝ�v��V?��E:��2�����ƫ���ґGF��)�y1>�wM�A>�T�Q\9���wS��A���<rqlf���-`�PV™��Vs���޻�Hn�.��7���h�Լy�7Z��>��k�x��|a�K�_��q���X��ܖ�T��&�:��EX]Gvd�T���J����n5�ꌛ�u��GHs*ae�Ya�O�w�z,F6���@�'ng i/�v�� ��y��e!\u\.A(�GS ڳ��+i
M���jd#���8���i�0�q���t>��)��Csv�3����GAk��h�[�P��1U��Q&�w��@
���2�[db_��VKN��z�LC��a���
A����ws;�Ƶ�$r�^���BH���%��z*�H 5�\�*�M�
G�����n���;����s�� "Q�8��L䣢t{�C����4��m�)��g���f�ec�J���u����KЇ�gJ'����Mפe,5[L�E��ѫ��@�ʯ�In1�~"O��>T2�`�>���fB�.j��M�)4����X��`�<K@���q�_��3��/L�u�U,K/��"aa=2v�����L�����qZ$�@q�(�wf��D*���_�v�����Mk'ztF��|�(���f5P�q��FI�X+�]�B�Kj���dd��0��7�R����#;�*#
�:a3��'�Y����A�Q���|o>�clz4(ֶZ?���]�g81��/���p�"�@�����b�L�'h�#�����C��KO�Rj�����0ӑ��06h��Ä��j~��b�UKR�����N���>hn0�B3!��|P:wC�Ų� CCG�8`Ϊ[�N��p�\`/@6-??����F��R:F!��my���~�$�f��Ŀز����ύ��M���;H�����ߒ/�B?����2�����夺^�r�7�g�z%�?���Vi�j (L-���{Z��چ��B�]0U��*����j�/(�H��P�3B�����x�ƞRf�{,lYk�5|��9��
=p��X`y��)�R���-b[���Mx��eQŶ��O?��)��$|v��Bs��2��˟�ݼ�2sL�کW�l>.K��Oq�2.��Ν�2�o��D�Ϫ��l���@0����WQ����Ie;3����=��r��C�v&��AC���&���B��lg �U�NE��@�1e[�\�lnE�)#Р�s����f�!�������F�b�J���$n�D4DMh�	4~�S��Z��i
P�mU�:�fc��ж�e?��V�0E���2�Vםt,ZS��o"Y/�C���R��I�9�su6'�ҔS%Tݭ�������DvQ�+ q�K~�� �a�h�E,�R��07]�6+
:A�iz%n�Ho���eK(e��j]�O�2���	�8؄ΉL�pƦZT��c�$��Rn� A��u}i�.d����O|��H͋0-_L�Nk
���L|��M,VҢA&��uV9ދ��)~Ϛ:�T��	X�o�.'5����\�wS��2��b:4<�0]�Ww��&j�;��V�hYT�O��E����@c�M.�P^5�e॰�d�`�-�.�i��7��M��L��1d�&XӰ�Jy�k�"_~��9��<�A��S�3�^L��o=�$mo���n�Ye�j�k�B����}��.*�mF�&Z]����`�����7|�\�I�S��o�\:a�!ag� ��tX�Sas���)��(`��A���S
خ���=�CW�Z�K~��ҷK�4��fk��.�!�}k.ӁL�5��	C����"I�͑�N�=�z��1LE�(�xuS҃��U���#(^��kk���B�ş#bõ8�ҷnҦ��ʂ��nG�7�:���g6�:.[�V�6}\�)�����`����R��K�B�8��2�����n���Υ�r�ς�!?f���Nj��[��2���F)��_��)0H�AY�S�$� T��Htc"Z��n�K��4pPԘ�H�������������u.B���.��$�8>���٥rO�#��܎�H�4X�(�fS���L�P\'��$�������Z��uS������]K������A�e�'�S�߹��e)�Ip�,=���|B/Y�,t7O�3�Hw��n�~�5���l�!�M`�n��"�h����>���g9~�R�u�_Dj{k+�ܮd�*����E�vAARa����\��^���ײ�t<�u�&4�p�+n�l�_�;m�簫�N�#�}T�ˬ�'ȟ�o���&[Bseh��4�.X��s-%2� 4���:�Y�b�a{㥦AZ�wLZ?h�*©j�`kw�t��x�I �;��}�6�{�D��^&I8�9���l5}-#I��7�Ҥ:#x�Ao�~��0���,T������Ȇf�U�H�. ���
LA7���s���^���&K�[Ŗz�� CC<Uc�k4���nd��� T0�r�����5��<Z�ΐsEm�f���K;	��b���(�t�cy�h��1s�чϥ⤢��w��~)�X�#:ܪP�I
�=^��ʂ�NR!���J�����[����/�}�N�\䜑��"X�f���w��Ӹ��������D���Q�"U��dq����~d�+��R��f>��X�u�L0��6�q�j�}R���j��< !��I�`иۇ�dy��ս+�9��m'"�(�^�e �P���ܣ��F
����k��c�M��=Ud�w��ry�GN�fM\)CÓ�ƒ���q�P�ˤ��k�<����-��ˉ�y�����\�Z�Ch"*Oap�	IQ����[Ǹ-$������={��3�E�̵�&�\=)L��5{�\�VQy�</�3_�j��J�A\J���xB�_A�ݏ��a������u�#$FnW6DE
���0�:�*K�e��N{�24�敍�::x�,I��j���ٽ�$J���l��X'������C 	��a�'���bk�#6V��-��[���#�h�`�aȥ�Zs,�X�ir���0��i$@��ݞ.z~s�X7��N�*��S�	jy7�=��
�R-7��/�^��iG>��A�C�����+b\��S�k��4S蘿m���~�ʐ��	Yӳu���(֟�����U������u�Qp��G���T?�`uX/��#���w_[j�=��"��y�UL�mJ�p���P�#ԭ�0�@�ָ�B�Z��w�ugM>zA���HlL�*l!�z��-�ț`��3/e��J�;*����bo2���)3�,s*�k�j�7��k�=�2QfMnВ�������oz8�]��)`j���op��s
q!���lp?��N�H�����>�%L�T��C4(�OL�(�^s8\];np�4v��;�v�y�QP~�U�Z�[�.XHu�"�O)6`^  �*��m?�z��������0���4���e�[�v��s! 9�]�%�p< V����U8��\�Y�y��~W#��=��
Nh��������k�X�i nX�*(�(��N��ᾣ����Y}��:����ܓ�����f'��~)/������H��!�)q��₈������L��m��t�� [��@�t�"جS�C������Η�QOK����n�*t�}�O����#΅����L�������=�鎡whV3u+�-ScT�������|���Z��C�`8C:�6Mؤ���0�8
����/�cI#v��wT�b��o�D)��QN��	 dM�o���Ci@*��`]$��֢��B)e��r)!d����OM-I2Τ��Mƃ�R�U�zHx8��k�\[�j���i�r�u��ȅeٛ7*FSKs݉�C��������Z�ĘМ��od.��>,\�+�Q`�a�+>�@M}2�Ac�w;j�E�2�bP�yMX�E��6��J������ �/�͟��;{��C8x+i�p�P.K�:TR�qw�n�J��i�6BG��ڭ�>��9ል5��\�;IY6�E�s(Yڸ"�@��H�b��hм5�_��JJ��aA�wА�/d�C5i�?^� �~+b�=�$P�ώ�|O�puϾ.S�4_wʄ�p*�R3�-��b%vo1��G4���w��#?C��C-|[(��LhS�1�|D��3TϞ8�v��e�G;�m�dc����ݎ����z5����Y��^2?yq�i��|��-�5"�"�����BcP�E�)݇��>��5�161�\;,M+�����Q�}�1y��:�L����^pԎ�n6��w�'�G		�,E�FVk�]�D�-��n
>�9�ߓqΊ:{!�V��y{�6Ć}���|H�%���qϿ4�A��9���6��4\@�Bm��i��jF6�����R)���q���J����"&ht��{Fn9��]>��%�%-"ĨFgŴv�β�l�7{ādF�X���a��߰��b���"LK��[;	˟�ǧ��C�*+�C�;��hOฑ�ޖ��]]�����q���h�����J��O����/�]�)A,.��נ�L?~Wxwۥr:�'�����ٓ��;�^�c6�#�ۊE��؟iu�X�~�2���l0����{;����+#����{?aoq�A7]��F�8s6(�p8�����q~r��:?VRb��8t�@O��@���Bf�h�s,�ur��m���*������D}��X��k���i4+�5�r�VӺ�YX��*���=�YP�i�X�o�����4�z� �v��"E�w-��}��a��M�U�'Z���f��r�o�?�X�TlrN�]=�r��e���,8A�2B�z��cc�c�ps�H:Dy���Ip��<ҹ����#�g�#�Ҁڤ!Tx&p.Fa
V���"Y��;ݑ���j�{i��8��>��?��vn��L���֚�mR�
$F�-��׏�N�x��WE�8���*���I�u�z��*�������|��R�" Z;Dܸ���Ye.��$556�uU[���&v"QaOmP�����y�k$�/yڈ6�۾^@�Pb�5����p�q薷�6Y���V��C'��<��Hq|�B�Y�!n��mN֔	Rţz�� �r�,D�N��Ov�D>j�*�_��{��;
����������i�$�m��W�Ͳ,^�R��MpG'�.g���w��u�7�	��u�����w*݌7~0�Q���L�Pg�����qµ�
Hh45=��N_�<f�܏~(:=�ц�	=nmd�>���Å�Ą�/�8��^�XJ��E���}��nlj�����8so����<��pK�d���J��o����埓�y��Xs�D\�P풜G8�V2������NאfQ�e�+-0*���t���2��vinU�X�c�pΧ�]:9�~�N�3��āHi>�$�����>��l!���N3���FֹY��I%VV���u�ۥ��?D
�˷"����1��Wu9���>��MS�{Q�7��ژ��Q�%���+)GĒV��9/�r���z�A�#XR�����{�:�>��k)��fC��b���g� @k<w���n�����}�%:��b]�=�0n�̺�T��f�6	�0����$��ڭ4��-��i�S�I����M�ZSe(�tC?�ުw�zc�lŻ�!�Ssi 1�l�f�ט�5�	nz��s�VJ�rV�K�y^�����Z����vHK4�(�V�~A[�C8矱sIܭ���v�t��G�����I��j�͓/��@�	��8UACj��t([O+����]����щ�ѡ�{��a���Y���*ӮAGo@��bb���~�"Õ�I��3#�y�ߣ�B׵�J9����=z�!@���v���1԰���o�r6ax8ٰ7@Z>&X���|���jqr��엚����>�z_���:opis�s<dd�Z`�hH�S�z�/z��E�t�R�e�,4]��Y�V �|/��U֞�'��;�<i$��X��E6U�[�7��s|�#� l���4S_-m�Q�4'� �z���A��=�z���g���<�2y��^/2�i�b4�L-Q�ɡҴ��w��H�q�X������+�������$IR�?s�R��_���d�fw� ������=J-�Bk�i7�c��:�;o���w�t�= c�(��ǣv�Q�?A=�����?#�Z,ɠ|=Q��Wj�d�̥<x��S�&����2xK�C�X���کvhG��z=�uU{n{?Q!�xq^7Crsћ��^M��OXՄ��kX�n_*ķC�a�H���d��:	��5@���nM� �|��s��vQ�$���Z�,�� o�|e|T��9ҤF$ǐ���<շ�_T�G��*��Í�j�� @ɕݡ�kC�������d	�5�7V��q��(���۽Y�����ŝ�_�yjM����]Z�(�3�6S���0+wV QjRrU+��:�3�DZ-��ι�F�|�;�;��_,��K~�"���w���g妇0i:��F�is�JQjҎ������9D(�>&"3Ķ��$�P���vhw�lG��4�Q�'<	�%-�	a���q_��]1/�)5��S���X2t������mIVOF�u��
񒉺��S���܅Γ :XQo�A��f�O�k�Z�f��]bCz�{���,6����x$�oh&��ӺB�Z�����< j7�fLU$�
*��o�k�ǩ�y�F�3w:���h.mI3p/��6�Uu�rSt~�����L�0h��hk=�5�E0�\�-9eԘ�ě����=����xv/�Qc�s�N���>^'9x	bji� .��-H�G�k�5���(LV��D�L�j��f>Nr��&%E]�+o�e���߫Gn�f�����u�$\3�N�ZS7�Λ|#&��g�鳬�7(�� �N�wF��H0���o�#�C�Z�?�:�����|���<��:H�":��KJ̴R=���.m��WQ!_�-�����St�5��w����}����R��<� ��B((��Ԏ��Cث�@xG	�c�?�QD<�hj�f��:���"Ha�3��G�	W*�����8����󰈓cFɐR��^^���n=94,���q���k�YE�_F��?������R��	gkR�ì�)$w"9�_=�B!�|Ϭ�޾�G/!ϑ6����
(��W�d��ܡ��H�E��E����9������P�"W[�NQ��,�ͺ��ӕ��1����%�Z7�	&h�;�k��qC5�Z��Ql�e�dU�왺.mȋ�W�����ͫj���"^�|��d|nZ;Л���+m�d[
�iD�GBz�|,��dŭ�k:�X���hј�V�0�Gɐ�|���)��njҟ�����h��Z�>J������o 1U2���ǞA�l�'�r�g|�����W��\Jsy�qQۂd�:�.m���2�3�+����/�6��|6��eJ.���x$��,��Q��ww�3=�c�̐q&��"���Duz2֝�̓v�7p�g��Q^yG7������]��Sc)z�w�H���T ��R*#-��P�y����1��Hlꫳ�=���+�RZ$��y!yy#���U[�ɽ�����m	���BL}��H		h��%�=�v(l�G��Rs�c�U��f�I��MX$](�h(L&�9���ێ,+���\T��0hq�~T�[��bs�u"C��#��ݟ�1*q�&\�m�;�\�:��_i�Ж͍h<<��������1��l��LM�@Ο��h�z2�Yҳ-GѬ��fL
7
QM5àǏ�d2����]RR�۔_�[�*�P��gT �.�v���D�	6>�xO|[H}�����s�Uri_�LOe�]�p-7<�l+A-Cx��A������M��B d��0���\��� )H|7��{5CM��(�1��Ga-;)^��~"�5�e({�
|}*S9xU���3}��p�{xgsm�����>����ܬzÊf�; �d��**�'0�a\��/oh�w+n��@(���٤�\`�Ɵ�JB�:E�S8��x����Hd�����5ix�]�(�5�Q�P-��,��>Y�0o������Btsw�̦<�]�0�%�����}S�Y9������V�� .�I�K/��g+Q1�撶��H� ?K����x�y�����ܔ<-P�"��Ȯ�&����wY���n�?Z�FxC�m��H���;�@k��(����F!��?-��l/�������2Gu��l9ȫ�.�,\���� ��lG�@�t�5HG����ж�b�'c�w�͢���b2��M���i͞h�-�����,�=�M���)�{p�A�tIW��Ӳ�X��͗H���'4j�7OIJ��< s�2;�t��������+�G���r�vˈK�
�=cH�Cb���gu�f;]
^�����HvV5�n�m͖�E� ��I�FĽs��Y!�����/��f;�$t�VD����"`_��E�Gx��L��QM���J�zl�t 6]鵱�p6��@����Y^g$i<!�����\�@�Mvp��?��)�l�*驨L)��0B��R���u }�'�2��&�FgK����D�u�,E$�M�/h�f�{p���l�:�e%,h#�Iӽ�b�;���L�Ri��6	*�&��Jp��w��á6�� �s{�v��cM-��_G����:_a<��t2c
��qk/�e��&@4@YˮΙX�>�;��'��)�������`��񼽩�=�^�i��g�	�0u�oa_9Ӗ��瓠���`������T���>��6�j��9T��2<R]�Y]l�ק����ij�4���g�*�wuxUB ��'u����\^B�~��( 坥�y�CԼdǋ_�n�X|=������E��Qq�k�x� ����Z���{p[_��-�F�oq����?LB��ţy���9L�5K+ܽd�	��ˆ�I'8[��\�@�H	��W2�G Z�^�/�_��J��w�-`\���r77�����O��X]k�������*�E����|�Rq!������:8�E��ͅ����Կ�E�#�+�4>#����S�"��U�$m>����q=�)#髊:��[e�e����?������B�a�� m�䉴��Mm�m�fv�O�

��ݷ�c1�f�ۮ�_+$�?!D���n��x���Qc��	@������%*_uFK�p���� ���P�T�>Nqf|�����x�1�{R}��N���u҄g���&�����e��1���G��\(+�b/U�o{�IV�ZЉY��W�fe3e�.ix
������J�T��)��q*�E|���̵�(j+���*k��%"0�|��w���3;���@Ͷ�&*��4b$�	-�4�Z�(n�/�Be`r�c����s������Ģ��l81��rc6�r�T����{P�Nw�x�s�����N���p�C,�D��foeӏ�dn��uI2n���В8*£b�?��=*�li �_���Y�6�o`��j����M�Z���
�&i����?��A�,����Ib� 2t�zSv�P"�7��C"�R��=���ls�3���IƹG �]�dm	��T���sc�����2��;k9)�H'wAq΋�f�<�gk-��a�k!�J�k�>9������i���9AZ'j)5*4?�0��$��T/04�k<����*�U�Z�i���a�A��䞑�	�N�� �T���O�u��H����"�����>o͟��f��<���@��skɘ ��NhVf2��i�9��ihO8�$���8�Tq�#&ѣ�5 x@�x���=BɌ��{5����P�Q�d�����ค���9��sX���_��M�ME��r.���!��B�h�A�O;�6���t	fC�F���^�Ũ;�����֏�2cg(�6$~e�Cg���)U����� �⑗�Dl�^��Kr�w�s��̘�A���{�"�ʀkP�kT���.z	u�_�������L<���lufJU_�(�@��?:�(��oo�=P3D?p)��<�G���C��$���F�D~�A�[���v��y�'Y�4��N}�MB�q�\5�a�����(��eR�7��U\�Bl��z��S�WBz�Y�,S5�����I��q�i�0	�)G�-;sS
\m����a�*U�6iو�v<�Fx�=aD�m픳����w��'�|�܂ӤW�c+n�hD��k�}�9e��e7��w����U�{�|襁ˠ��?�b�+�Hn%���M�y�	�;��*�7�/�ht��P:b��7ݳ��P_�FwG��?;u���[1A��~�gf�$�]�w�|/�Bo�F���b�����6��G��������#�T�h��{��I��.��+�A�Ȑ!�.�`��1ݎ�l����Weԓ�����H���cykπcu*��c\���<N$C�I{�C�O���e�l,�b?G.�_S��|���A�U^V��<�>^y�}�����.�e� ��O$���?;��i"��J4*lD�yՁ��Y�+`���uJG��d��XW�� A{T�ʔ�����$=н�n�e�%��D4q�G)|Y��:�⛣G��qMZ�p��4m}�ar�b.߷9Й�Q��?P:	�J0�B3	?F=���Ӧ��'����Eg���N�Q�X��R���*Q6c�7�w&�i���x(�Uł,�K��t�_��5o�����mL�-��mU��Xi���f�]�b���h�����,l� �p�TA��Z��6$��}*��R6��T\��] u��7�&��Ά��'�q(��da5�q�k�4�Eav��b�Ǹ'W6����B)'�Σ�?��3O��y�sP��=ڄ'������h|׻Òզ6׋������E��w�(�Lju34饏Cz}�\��4w�{⡰|�$���5��Τ�bK�6����An��e�[����!o��R��t���O�(KV9}�@��p�n{�^�^uS �y�����gY�,R4�bՆǚ�?L�l�S&��i6P�B	De�^~۴��C��,�٘���p֛��XY���4��Y]��웋2���Q9��N��x�|�<������S�S^|I�����: \�i�}btl ipme>?:��jpW�!�FN��:)�_YVPo��Oѽ��G�^W�e��0`O&r�<�7�(��o�%A��֮n��� s�2M���8?20�~� �a�h�tR�/SԽC�AF��P��/����c�iւ��H�Ջ���#�ٹֲ�� ��х��J���r�HSZ�7�)��q�L�O��j�])'�0"!ΰ�`�#�\�{���l���FP��
Lϐ�uhkˋ�۱������+%�1J#�3�*t���?��t�s�!��o�+N���DtG ONzJ9ae?Wq���|GG$�>�	�AE:��ɤvE�J-�����{e�O���qy���Rz,@'`�6�pY$�:�D�M��E���K/�����G�G�:C����eMp���~���=#�ի�l����.��o��Qz.�����i�0���;��KNa/�P��.�ՐW�ꑸ�$���w��W�����Y�c�e�/̍V�#S�!���Ͼ,�H=�� ���_*}�ﯹ�0N+�zpu���5f�Z���8�|i���o���U$to�cNd��]L�5�?�6�M&嶬���\:CN��Mké\v��݄<�Z��H����+>���lK��4p���h6��Ӕ&��#������[���n*h(/��df�f�?��i�C����vW������ ���d���"��M��[�1�]Bh���2�	�Ս�J�5�R�H��+8�f�����f��xN��s��y__TsX��U�Z��0�jgr�k_�mj�Qw�8͂�1��l��p<TX�Rx��U����p�N���m�IUQ
�W��H�#��ys#{�iP�kUW8�+�^[\OZP(��Y���0o��W�E�b��;K�[!E�g� x�VLe�z@\K˜�,��#ؿ���F�p�v.����(0��<��%�k�7����b"4ޛT�cj�ȣE4��:�͎&z�c�/C�wղ�ȬTb=��!��C_����:ē��* ���ɬ1�?�_�s%����[I7��5 � �3P�bf�W��� ��ڤ;x�E� �Ӫ�]�$eiM)�V(��������VR�(}��#�p���CP��Pd�yˤ����h�T�
�ת��I�d�pyf�~�M�49?�<wMX§1��|@U+�j�.4��$�q�a��3K_��|�9�A�!h֖z���[?/F"��ľ>#��s����ܦ��0܉���@Ԝ򗉄�on#�ܼ�u"�p}�:��ۆY����0�r�X��lW6��u�8���}׳z�1%�`6���!�ZM�y	�����ܬ���B�	-+��Ѻ
���VAjLt��v���R�Oo(gQ2&�p5>DZZ{��;C�]:�+n��r���Gdf�QaY�n:�h��u5#2���{�]s�CN���'���̏�B���;a��Q�x�f��@S, ��EȐũ������67������U��ȒS�G���L��z'�=X���:�0M���^�ؘ�7-5 �{�14!��#sh�ibXImc��P�(g+�K�����41�_�V���=�����]Gc,�U-���9Vf@�sg�HS�%����KJ=1�� �ƀzG�����e��H��&i�FGB:�W������-�,��t���6�jǨ'��K��0��J�c���l�u)ʣH��>*���:G5�{!*��x����t���!^�6,�ⷘ�.P֠wܐ���4�G�yyq�w�4�A�lX���8���0ή>If��+
b��̮4Q�1]�;Qoa���t%�t�x��W���ڨά_],�L9�4�}����\h������=�S�#����v�U���b.��^��u�����sS�:�K�cE��x?JH�x0,����90�����`��dRv�����D9�F�_>o����zb��U�1Ϝm]b�tk�����@�џe��D���0@��9��?�SeJ����
�x�5����ᤛ�Z���m �*�圃����N�E"��.#Y+�Gɓ� ����<ͣ>\C;:!����a�+�b���*C��|`f��{�UrB������я~V<�E�[Y�;�D��l!��6�f��(�VB�����*=$,�������tt�=�8	B�ťq�����Aդ��l�(���?��yܼ��!��FrJ��<�Y�wކ9L!L�e��,6r��8��-nU�U�W�9]1��$2CҔ<��R~���RVe�fKZ+������?���.X�u�J��S��8�K�,�S+�u��ھ_K�n��ݺ7�9�7������Q_��M<^���;����`�-+<�G�ښZI<�o$��W�ɲӜp��%}U%�j�;eT5�#Q�buJyqoZ�{f���)����c.�\0��H-QӴ?\:��g�n��=�����!k��+';Y��<T��S�X�A�%fc��%o��!8z�1hZ޿�H(�8w����p����ൡuF�|���N����s��钶�i�D6k���y�u��o�mre#"YUnjq����ew��a�8"j'�vI���>�nBϠrrP�����=`�_�\���Fi���!�
�����Nc"��?�	{��3�Q�B�'y��]��c2�9-��7�ԓ�i�t�i�����z��f���tQ�PD���a2BQ�H��-9:6�Mg�7���CmD�-F�vs�K���I����>�lf��#�i����ܮ��2��f���EZ� � ' ��z���	;]ʩ^(*��9^�w�푝*Ib&����Ş:X��0�����@d�����a�Zً�P'�����K�M��RwW�s��s��͛E'�"<F�
���[Z~(�;L��)���J:H�#�Z����A��u5�g��+�|�w��W��"�}�s�������+��������[v���L@!x�D0.��NX)�Ni�Y���e��%Oξsϵ|mn�/D�����r�-�E@�KQ��t�3�x&�~���i6f�Z3�`'|M�8��������IԐ�Am�A�����%���P��x�1��.2�A
)mH���IqDEc�`�߀L���+bi�ZG�Md
�qe"�U\Y"��V�E���s��#��B���c��r�8�ӕ�]���NE!`☲Sm�6B 4�æ�WO���o�g97@�.;]vԆJ{���A=����������6`zS���%f���J��B�ƿ*�����C/M"��y��G|�9�h��VM��{h� RW�Ό=&Cy%�ەం0E���+��@�5��)�l�\>�5  �������&�c��|4v0�Z�u9����bZ�����֣X���<���wV�&���#uIL�����Pj/�5�YA��A��?Z"��A�^q�!7���)	 Sq)d�{�1�Xs��n\�5G�L�|�JE��\2���k6<B����I߃��=%�J�V�f�u2�'l�M��WD@���ct;8�ڹV��u�b%�����QC]���y�33�-Z�Ҥ���z8g�K��f�M`�{�e?�������N��%'V��Z`ɢ!�ӻWd� u�/N����E�A�H�i�����x�Ɵ/�_iG��P�Y� �\�+/�HW@s��M�-(e�PGf��$z�,�Cˁ���z��I^�1qp�$W/�ǧ<�
E�[״������%�2��3�{i����'V.�͟��^E���F�A�+E�8uM�5jg?n���?;&`2��E��P<J�n~R#i>�f���#�\޾~����*�;)�M1���/���x�Mo������I���tW+�C4�,�d�"*�m\�=w�S��ͼq8��M0���,&.�z�k����zP¯�`~�HF淴X1��zy�T�K��K����.�q�&n�ǲ������G��X���w��Z�v�gKK�^�hʓ(�shbڼ����9��6@���-+�������f��y�"¾�઴�ЊTl��gHN|�6�vdI?r���C��=Ӊ���a4Ȕ��8ȓy�����)�hHlwVh<���(BK,?雅�$9�\��W��f��`�����10�����J���\B�˱�����q�	��-����hh��\d7�3�b(��Wߛ¿k��ؠ�Xܸ�Nds��W��A3N�~g��������J�F�w�e���6���fbm#Kf�2��4}^ ��R!���p{
2m�#������=�8|���i�<��7��Ea	��u5Xk!��.�v�AH�=V���;qQ����$�NC���o�����Ư�-("|?��uB1I��X���V�߭4��he���z�kKE|%|ǵ˘s��|�)-�k�z ݫ���F�(��UZN��,��x�Hn�<�N��P�@*�v�EYN_v��~�إ�K�i�G0���<�C�*%`�;�G:ex�ޯ�Miy�:B8� �%�:\ęZ�N$|��F���Eْ���zw�Bp�,�p�.Z'�nM�˚n�蝍����.<�N�X�/r�� �(�A6ų��������j���$h���-�5�0 �|�&n���J�q��zA�Дc��8��A&RСuK�.�
?�'�$�O��ȁ�v8=*(���H{���W�I/��&&��l��ZF�.���h�ZQ��#	 o7�T&���������ጣ.J���P�5�g��5	�������_l���&lm�.���>���uA�$��U�g���%(p��S��)H}6�>�,G�U��?�m�X��l���Ag�{?���CI���no4ț]�!�X����'�A�!V�����e/e���#g0�!1���1�\�:�Z��iP�AFy��6��%jq4ѐ+D�͢�P��8Q���>i��H�]-f+%y1r,���7YI;Ķ`���t���M�/����W	kڦ��<=�'�>�rTe�Dz�������^O�w�f��~$c *@�o�h~ѹ�\�w�#��y���PX:
^-���#�@��4+��*8������U-�w]��̙DU3kx�ے
֩{"�y�b��X4*z5�������Z$E=m��&m%���մ����<�b�FG�<���-jЃ���*?�㬦˽ky�&9'Z���܇��X�B����A\:ᖁ^k����teMhbuoC7c�^+�=7j�5�%T�w6�;f�%;��&}^������!v����[�V�l��ٳ�rE%@^ �'�a��ψ�\�'����پ*UҖ�!��P��� ����_����P*��$�eL�MM���������C�I쬗��"s�6�B��e�_�È#�[(3��H��,��q�K.��,�#[��V�OL�Z�0&<�ݷ+>�g�	���֒*0���������"^]���M�0Od�
�o�o���I�$k�T ��v������b�ʣ	�,sm��ְ'����?�U���B͝r5�_n��B����-	T�K;O�]R�bGT��w�������ƫqe���lK�'��uH�m�w�^zQ+hʥ4m/�#��$n�fCIA��x�;Dd�s��"���h\�'��sUQd��#��mL~��ZWUؕi��l�%p4�c��7z�t7��5
#q��<Mt�b��Od��1�d.��}��RH��U�����)Q�<#�7��YM�-��ݘZ�9S��Y,5TBޟ|�g�
ҁtF�Q#m�T���V�y	���B�{Ge��iD�%V\?6��Z\���i��J:�p��)�=����Q�O���K�U���s͞Q�� c�^���Ǣ�	xdVtY�u�6 ᛫g��K3��DhF�f�c�Se�o;Q���-����=����Mo�s�^��ȑp1֓�g�ul¤�<X0�H�Z'0J�]csjz������[�D�=>O�hc)��q��2��f)�<�MBr6:T�r�qل
5�}�D�/�$/[��|@�M�<^�}���!���K!]P
��^%�[�Q�f1�N|ih�Y�GUY��ďD�Q�귃���� ��2�YO���y�@ ̛�����X�Ɓ����
X�ld�4�:��<t*�mTX������I�Z2�G�CΥhY���c�3i_4c�<�0#�gwq���­Y�0\�h��'w���טz(��xzo �a�<��q��ʤ�GT2�!0.���G5$鐉�4q�g���w���K���Bl'Ե��I8$�8l��ԕ�r�o=&&b mWU�M+m{^����|k@�(��:\�L�x]�^�)w���S������m�@�|��|��4 oQMR ��<�(u�^�D�E�9j���Ԋ*# 	�M'�0������k����Ċ-�Y�&��2�	_�{�S�2��Y�"�	f|	�&L�������2B}�m!@���a@J]F���Y�#�f��Τelk�<���߾0��f�+0��%�D�Ur�O6����ǆ�v#��I�$�p}�/��B��>�~�2�$����Zq�6D��Y�n5&����CR��fE��a��2ے]$ސ�	c�%�j�D�}9P^�(�`����Pmv�B�RL4��������D�I�'�N^=���l_���	�Z}�B������=�����QC�(��YF�$�����7�ƈ?�
����V��jK�q�X����C&�:��#J�Z'O.���tw��[��;��u�/��Q _�m�0�F�݁��`�#�N�V�-HQ�U��e�D�`�^1}q+��2$��ɊV
�)#_L��`%��Ѭ]Z�}4i�7�/H�z��F��������$��2���i������`�fփ��<�o��_ݩ��ï��������� u��LX� �f�Ϧ^waL6���Y�r���J��'��%3W�@/�G���JP|p��z�m>������2νe�[�O�'_AZ��;dP3�ap~R�ƌ�!?@!g=U�sÇ��QgR�7ֶWn�~���y��K����dOᢷ�mY/KS�'I1�oC-h���I��-�.'����묳�@]Fr�E�5Yz& 9P@s�`ւl'	j��'ʀ&����\��P�%�k0�`A�n}�$;�=8**�b�͉^�o-�T����k�sI�F��ڼ�������X�Ǚ��H6)ar ��K�Uj�b
(�r��M}���"PD&����{S�A������7�X�����_����+S�+���u�ؙvm�0��jIܱ9I�n�� =RW�V@�rթx�U!�I�\g�����q����6u5��`Ѻ��8
f6��^�r�k���[Ȳ��ÚN�7��]��I_��6�i�Bi����) ��=l���c�e��~<��_Z#3Mթ�(>V�q|�D�jΚ$$�H�t�߅lIGT���l��/)X�����
22%p���/�w6�Jt�5D�� �ds�މ���b��6��c���DM��6��b (�<��6 �~〉�B��X�L�ԅ��ඣZNwx^-������Eȏ(N46;��lJ���T��'U>��Q���7��:�/�t?M��?�Ʉ�͔lE�!��p�o��O-S�Z3 ��)0ȜXhۖX�{��'�������m�8}��mR׌ �
5J��+C�E)�)���K�I�&e�ן\J��6=���.hC�v�v�X~���L
�8�DQKn�f���o7����|"((JS��$���=�C�<$
�3|2%̆MÔ���k�Ԕ,�6+�gX�\l��\З!�]%��2�\*sW�^�;®=��ȧ-�ۤ�5�d�J�"(�ꔺ� a]�
7�!z�TBݭ�潧S�C���A��ul�7�����L�cb�00����*���iZ#����D�х�;6l��ES o��� ���+E�,jp�����hG��sܻ�G�B��ՙ~j������8��P���`m�vbƠ�
Ĺm���0����kz�w;�ٵ���͗�.YMI_]P��Z%��ym�*�6��Yeɋ_l��{+ȟ7e�r.���y���������rT�8�n����TIyW�7K�4��0x�����ΓQHl걌�^o@(e��,�(2w�&���,r��YֆK{T��\s��'H4Vތ��+� 0y�T"��޿�i�q?�����X7�UK�:�ۗ1f��v�НDYV��.���zQF����wDo�:'R~@0�v�`iv�ܩ�βQ�
_j΂C��!���2�æu6!]���y}�́��[з���s�Hι��9y���Tu�m'-��&G�����V��_���l�$���ǰ"�К���9�@�6��^��rH<�����EҦ��c��PH��аG~u�7��פp��܂�@�Em/�2��������Ϙ����"Ⱦ���Vrfc��v.-#�1I���G���	����mʕ@��U&���p�x���g�C��_��q���9������J0N Y믔N���o���m��N:Rq���}?�(�$��2�{B5��K�G�`�량4^Щ{� �k��'šhI]9��<4�i֎ 2��C���������t�2���l�E�����{h�t{�����mR�l�ӽ�����8���-()�t��]	9�}�ogQ�R)�����U�nF�䑾 ��N,ji��K��8;���Wuf�B7���s������:�hΉ8D��<!�}C���o[�\���z�ɜϗ]@��#���@��E�h���/��/��2 �Pz�<7�"�T�ˀ?�w���0�$�sh+��-��n(1˶�F�ik�d���iH�,������X+GZ4W���Fj�pV�(��~lӃ��:8K� �L�<և@˃�D�"�?������}t��dX��m��i�����A�7��|D�+X��=H�]�M��j�/5="@�r	*(���ҡuX��G��K����/�9/ Ɓ.P�rg��8��꜃�$�����l �d�����O���e=�,�[	�tm*t_=�W�@g�U�:�n0	��>ibo�&��P�?�Z5�[8��m~�Еj��&�
�3"��I!��9�l�1_.��ؠ}�	���#� ��� L^6	i��`�o��.]��M�x
�����g�����Zc��4m�&K4z	�V��﫠K�\,8�N�O������H�U���;}�<a�s�����M�5���bg;�,p`S���L'��`�N�V�)ᶪ�3�<��E����N�#�i���/����;��FF+X�i����MUs/���W�5Z~�����J�L���&F������U,��`�`���z� dC�W�:�9d�w�-�Y-n��>�U��+~6��7�µG��4�c�=�[���cИ�m�;��څ���'������Yl"��?;���G�c�@̟�u!��̂���%/y$Є��ma�(F%X(����F'��*h�pF(��~�m��\t-1���<��3��wmj��ah����5~�I����^�FO�j���ls�+�~d)@��?���!�.ܻ�M"�c +q�Eƒ����/ �Z}}0��B�T�8�!�xxq���t�xTP���Kj�����%7IK��b/���p�Y0�#Cυy�5%�C&��.�� lS�92�x10[�9�Nf�f{���׏|ȩl�jH^`�W����S��&��]�#w,%��H���}��ٵ��|ű�4��:X�0$T�t*W �����Q���1cv&�.��Uy�����VY���B��,ma���#�[�]q�&?�����L���*W�`[~��S;V�(㙣>�˲	5�X3���*>3ASK8܀�l�"@+�7�{�o	�f 9o�r�|\��h��$�!C�-ޣ�*�!YIٝ����6SH\O�¥�)�v��g�y�+S�cH�5���URJ��N{d-K�s����c>k�&��B0զ1�Mf"�x�96_A��1����-�
�p�,�7Z�_�x>�2����?Y�z�J��z�����]M ���
ό�<M�Ҥ��G��=~���m&%��38t��A���� �:�%���~}��o��k,>1G��{�u����HTx�U K-~����v��L���xut��ЌUғV�h/g������
eJ&'>:���^��vqfh"��դ�z?p˕8���V�_�+��䥾�}��P8�oŉ硚d+����&Qϐ�>oà���A�����w��7ç��`g8Bb���z�������Kl������V���,ʩ�C
�2�6޿��G�t� �+�R��C&���b����,�+U��:���R��p����C@���i�H�
�'�g0�����x�|� B��t3/�J�����h��:,iY�����h䢔K�D�i4�]�J��l��#�a� �ߺK�6?\�,�R�T@{���- �



�	s%�*ھ3�ɿ <[�|+�yߐ����j���q�j��e�����eR�v�'�Egi�	1�Wŭ�@g��"<�xt2f�q�9gةD1�	�m�>@��������$�Q<g��=]���.��v�|�[��r,�X�^u\���a�� z���g��;�5��������7~�w�c5#n�7�jZKŷ����ܻ�T���|�.�Z��7���U!�{�Vj;f�˓,�>��>�m��k�(��}dt�\Aۋ��)�/�̚��8!��ѧ�xu˹�Nף�uq��t�}��G�v�5uY.P��5�`'������Ɯòg!��X��oPu���}����G�o~mJ��-����Dȟ3�۾��GU�`�6�(]�����v�������B�n�!"0h��6uYr�� ���5�������=��Q�
���9�CMdh���]]!p:szŲ���<{y�"�0D��b�1m/,��zVƝbv�݇I0���������/������&%V܁��=*�>mx�Bcߡ:뚝Б�B�=�\���j*ː#�М-���1�6�]H�{*%��J�<.����3)X��kfF�"�J)F�ݨe���4�� �֟ƍ9�E�_��4���VI��r�H�+dS'�J���NM��������x$}<t��D�4ݦ=����?e�9�MeOcbf���e�΋t�$u&�p�������� r�6^�ޤv�]�1���ЮC���.1������>s$�P`�H�׀���$
��Qp�"9�#���`�L�+A�B�u��#��N����`�pQ\G��	72���X5*�ZO>O ���zҵ�H8E��o�8����CbW x�m����C�EV'|��F�Ц����c�2!4���mh���`S���3�E��EA�ʜ�ѧ�?���Ai�1L��6=�`-DB_�,+����l$��p[ď? 
D;E�s��W�+�G�$�SQy��|-8�0Fl#�(w���'����8�p\@��Xą+]�7��*��.�.g�ae^���4�G��������݇�Zqn�)�u2�/R�e��^�mI�	5(��HlXYy5��:�>�[kS�N3����]\L��-��Y%̐b$}��oe�
�a�������bf m	y���noX�/K�v.(�� 3V!����B��<F8��Aխ�KU���:@�ӯ�<�S|C ��j�fI�r�������zl�I�������4֛��~�2zdB� D2�\��h��ǟ��HAN��&�8���m��lυ��tA���7�<em�A�R[�395ͤ]�Tӯ��/cL��"�d>xYE�ZK�&L�.��|�Q�����>s��34�(<hz|4�,�[��TɣVV��6���ə�.�C5?���w3i�;egN�wE8�d�>�h�x�^F��w�Ⱦ�`��O�=��N�G��)���GULxȍ��mޠW��lЖ�_N��Йo��`o;%ۨ:J����F�����Y�&	d��,�p��s�0�d*7�-�v^��x���]��`�Zl����y��_��fwY�K�%� O*��Mb����$!�~�~�@��Z3����Swu���k��q�O�Ҕ.��<����HӘ���,b�~c��^�8 ���O�mF�8�RB!-ȳQ�5J���Rc�X�ʍNί��.��.�Y%$/��<S9�:���n)�m�X1L������6��������c��3�d��݈+d� X���j54��Z	c�r��p,ɬ�g���x"��m�� Ɓ%_�2]�¢�!�o����5�x��e7D������x/u+H�BjL]�x�E�R�HF�wK$��p2K,�y���;�5��uE�y��h3i��=25ꗝ�(2i�/�hf�uM���w�y{�Y��-ku��c},Wq� �k��l���,4�rf�����*#k�}We�9��kB�<����5Ll`R���:j��HkL�d��%���A���hA�q��`*����4�O8��5'a�7��y��{i}ˋ�F���ՄZ��,%dj��t��\罚�Tv�ֲ�	���}���Z�(,}�oc#����k2D4a��\'0�^��Q�q����(S� m���(4�;�We�)-�]O@:�&�Z�	rj^��]��N��\��b����&5&r��^��G�C�LuU�#�(T��ab|���j5>I���.�
/��#T��2�R�J�k5��;5�g��,�cЍu���ޯ�ꑉZV��y'�6��S���T�#=MY����H*�>^JL�����~��|��~�l)mӖNnq�M��F������5�a���ݽ%��c�uz:k����Z�ˠR ~4f�.�+���3e�J6{���)j�`|YX�5���_* �Ha��\�"�Vۧe�\J���3[��ކ�� �rXw��N�!Ι���)��9߅�D�BeP�چKJT�X���8t�gl>�_ظ��Qoj*�6����:���"���r/���p����T-��ĩ��|�oƓ_W��o͢Ќa�}��r��}I�K���?*��C�%�h>�����n��q�{Sv�,��هC��ry��������%gSwz�����3����p�	�`n�����*��t�����,t�dB|kF��	�F���\v[�� N�x��g����'�0����FͅV'�o�Y�I`�h��x��RN9�a�n�Ygfk�Κo[���u��0kã=Йs�5�����zbWCHx��&�	&}n�ׂW����\�$t{��_��H�w���ZϢ�m�m���OEi�wW|E6�����`ɘhdtEXgI W�h�`ݩ�Nu����g��6��,�S�]�A׫���Bl��}ϣ^�?�F�-��⭳�ȷɩו|WU�~�������weXR����h��Q�	�?y��Av�cGR��8'$N��tT���#�y�5!p����<��g0`�N�靉.�v�����sX�n����f�F|7&y��!^f��M�[08��dlպ������mRS$;"�M��/�俭�*��<"n�]"�6��6��Ot����IR����ތ6�/!Q�.'�������F���@瓥��Y�QF� B�{��'xFP˶�H�����;��f����bR��l�ǀ@0�O*3�Q�G�����L�+�(�c-�"n�v���1��-4�E˙�Bp����M�^uF$��k'��h�S�	m��O`�O��wJ� �VY�Z���,�[�����_���'O��u���2�ߣ ��i�ױ���&�FD�ױ���1Pq�wK-`�l�@L{�38GW�hp�U�����;=�c	�4���z=Ʋ�E�B��1u�|�tZ������3�8���q�|v�T�I�Ֆ������˯,xt����	�]����rS&fN��S�^����	�F�{��>�F�x��������$�2+�4���� ����@}'3'\����[��"Ds!S�����AK:lۡ�s���z�BJX�-���:��y8���0T8nVbd g��?EA��R4�m�d�	6�)�I
��0(�\���ij�Z�F����mTJLH+�JX���	kO?�9��ĕ�BE��뮗��K��/"Ħ��,b.�Z}�ZZz=y��|DX����܊�A��Z���@`�9ye���'�d+4f��o&̒g����}�_��ؒ�Q�q"�5��'���F�

�]Z\��E�y�w(�p�xsV��h��IF��V����R<�N�C�|O����[C5K��k�t��j��q���Q�z��mu�6$|p�`�ۤ�&�:��^ǩ�W���� -R���J�&c���O4�S�6���{�SMQ�{.4�%˪R� V��_X.!���d��i��z�g�)ojR\^�p�З(%+�� �և��V�nP�4Цw���a�2�X�D��<��8�\��R
ڭ/�o5�ή#�\nMo�Ϣ�'0nr���圎0��12)y6���f:6���ٝ�m�t��`����c����Tx�o�p��I�y�mq`�9���H,D�v��j��CWp/��RY�Ĭ蛃���d�ɜ�d \�`я!^G�2hΩ�yɁl��
?/Zp5ؓB��ƃ��<�T�e�8�(�5ȵ*E�%B���Y6T
����_�=Z"�����Rv��W0��%&̜���GB��dD��_C̑\bZc�! �������Z�L�݉���aF�s[-O�.y��u��$��Cp��XP6t����D꾦C_�r��@/�(�=Ѹ<�@�_{e�R��o@fl+c���W��?��e3���nZ���	�P��!i���l�`0�ڧ��8��R@�H�a��
d�����t�eF�'/9FÓZ"}��YN*����|Ω6�f;���$��,6��F��ͽS�I�+xi�����h���"V��i$RNΥ�AE��R�`�"Ʊ,��~�{��\�����ݨL�bk�CO�w�rسDL�`&P�K���E�B6�\���*��� ��ᡟ-ݛi��� ]�/_R"����8lG����nR"��t$����h^#[�-8<��o���d��%�6�:��
A~�/3�O�.!�2!8e��F��V0�`{�ڥ�� |���kS�/�=��e*����:�m��|e�=����I��?��\"�D���~x�[NYD}F	�C��8�������|W"-2��s�Y��Ee�NU���@P�iu�=��A�<"�M�B�D*d}n�C���Ѻ+ys��p���HJ�J�yfA_��֏�����Z�J,�~��um4�W�e��;�@�s����=5KVf�\�`1F�C�����.y���aD�)�oFWN�	���CIU*/>e�{_�����<�<���W_�K1��hY�=�n\��w ��󰺳}p�Ld� ��L~�[���}��\�hF�X[�"�z�r�bAû�|�޲�|+��e�L�+�y��T������a]�#� a��8��-�M �N�x���	�OSwI�z���~�3�jh�Y0i�T��|�ע%�H�ʝФ��EW3���Ǒ�_�64���f�_/t����p�P�S�9b��3�<kl�Y�7v�z*4��|�c�_s;�� ~9�C}j���o�DW|�AB���O��,|Xa�ӱ�����d���\IM�2�ZߙŠ@���E�Jy*:����p���C�>m� '>;���������/�~0"�#z�%,z]��VKO)���wKm䪆��:�����w��������=��{���4*2C~��쁫���=�Ck�G
@R��`��ۙ���
tb�70gb�Q�2�CZ�1C{�_0}�����8��_�O_��?p`��[e5�d�A.\���Ո1�c��B�����nʕP���Ą"�av����8�\ov1�P��~1�	I�~m�Ǹ�_��SՕ���[Z�m��& C��<���� P	]��q����"Іux�AI* ����Ӫgkw��y��c�Оslp���^�X�9�8Z��#���8r�W[FHK��ܨ���J)��RfOq0S�x7v ��8K�� Q��3��XPW��m��9��Hђ�뙘m�H:4)�z1��Z��n���W��U��E�� ��y��tڣ��f*�I�#�-Ц��S��7~B�8#Z�~�e:`���*?<h��t숟*�X��=48��m�I��[�D5���}#x�t,d'� ,�[=�"���M�!Y�k�k޽�xD�.���.��p���Mb-I�~c�;[X�WnaӁ@a��o7Ͱ[�e�K�朲���F�ku'��8��:�j\�I�GmL���4�N-��� x����P��2�Y;�t��o��M�2K�O_�w뗁��o涒��f��A0��hS�9$\ޘ�¹�y>��	������2����B�C!8�.���@/�M�LU)��Д{�R�	����B��@���%$���kX����(A�)BK�����̜���7p'�dj����	�[��sg��`��7��'˾���|�q#�ǣ{1�/I��M�&��~U��T]ՉP׋�!-mzU��e�quŨ(h�H�����q�X,k��%�O^q�S�m0�I��¤�n�ҷ!9P�l���lX@��od�TOӗ">�~"~:4�����>1�����u��5���J���A����
0��{uDK����3B�s��h�:��-�2���.�5|e����g|!��q`��i�A�^��>�ײ=���R��(�whVAec��B�U0��� f���R������e9b~�����_}%O<6� #��!Ց(��F�����U�>�
nV��>K��'% z/� [|�`z�R��@���ft���.LH3�5"�y��%�������{��o7������(�:t77(�R�\���#߂��uY�s��_�:V�%`˅���Z��)��V&�m"��]�u��#q4�O�zE�NF�n�틜}�����+�X������$�����0�t���I䧰�cn�dh��,h���R ",��&����$0�7��V�9̣��w�����-!٨VCϞ�s���Y��)��{(�y�*f�OIֹ&���[˰ӤZ+z@�|���o�R������98���uZ��{�!���8	����igDݦxVe�"嵆f��<ww�>g,�7:c�E��\E/�qH."2����/q��\��t���e�a���c<q��6���* x��I	T��:k[���5#h�,�w�b�(����(C���r��If|�Eu�p)#2~ƈ�^dt1a��jD�׋��
�4V�#�0}F;A�Z�`��*:�A�>�����c�z�OZ0���{�u�73� s�c��\0Z�{E(���[Q���J+�!M-V���)���_ӵ\й�D�U@��xRi��Ij���<�5 �0�K��+G��*��E�<'JD��DT�GO �K��=�%�#ێ�I&X1J/l ��S�߁�Ylj�yKW1���t�e3e�7È����؎
�":�4b������&��a
��>�6� ���4ۜ�����SYĕ_�D�0ܟ>	��J�V�sr�)�U.ɮ44��r�Da���{D��C��c��=��q��`���(������ &b��w�����?i���a� C;�{��2("�T��j�3ҿ#��1q/��ӹ� �u����"�_���_>JgE|�`���Zx��q"&>�����T[�!�i�`��% )�Qԣq��~yK�FI�� U��i�\�lT]L`5Q��������e�d��nG��O��-P�x7C&v�xc7���Y?��6�E���L��`���ʶ�%��6t ���8o�7�nw����7��8�u���d�_RǠ����9�=�^׽��{�C�{A�Em���0��ew���4eȻ��Z鏔Ri��r��~'5���>����^�{X�����'p>�O������y��S��j��כ�.f<?��.i�	Z�v<(�m���%��
�@+D&��P'B�L�L�6�Q�!��}��@�a�kU����g	��WЃ2v�]�Ά�������v��n:�O� (�a$�>�	�;|�-�/�r�L�3������_q/� B,9�`�[��d����)�fY�p,��|"�Z~�Qba�����o�`R���se׵{��oK����BAA߲�n^`PR��j�Vԙ��4�&�&ΖU�C�7P�}<�w��+��ˣRg!���`s8�m��O������k2��F#��1Q�8��V#��0�L�/߈t��)3Q�y(?Y|��A�	!&�3;�(r�X�*��Sza�o1�pi;�_T���׎\CI&�3�S7I6��8y�z7$+%���h�p��D�L���|��vT/�̉w�W�}CXY�f�5��n&�A���8�oBo"� 	X�S����
��f`uj�� ����F�e֍�U,�\�4��Yb�ġd�`"l'� Dņ�6\P0~F��7{bi���c�o##FJ!�j7�ܲ�Y7� !x�2G�_Fëp��c��W�c�jI����;J�}¶����ñ�Ф�L`N����$�	���oӜ���2
ӣY��v�� ��3�{�J��[2��GC�r܎%��y3��_�p�1�|��IaS��1"h��i���MA�˵��K�KYn���r�c5)��Z�֒���!����v,s����6��M���#6��6�u��⺵�;�*G���G�uQ�6k�v�dO�#�j\�V��F�i_c�ď A�����>�o�\핍���`e�T�BU��i:�F���eu����o������.I�c�3>}T��QZ���s��.�򄕕�v�6A `�3��e]��>�A�.�G�oN��Rwg���8*�m��X�6��['"s�7+��(�Q*�R��]A&��������v�s�g���5�`���@$�3mRh$�j~�(�^Æb�?+����4�$�G��oN1()�*�>��	�
!S�^Թm���k�7e�Ubj}��|��2s�m
���U&�����	閔H�;���Xq��ӟ��-Jx�ZJ���J�6�r˔��o�guxa������E����Ȱ���'��G�`R�F��J~�Iuژ�*7>���\~2���ۑ��:����vѸ�HS�q���ՠ���]|�2�4׮�o�3m��I`��!���(���h�[�"��E���h���u�=Ω�s�7�>�c�8���-Z��"A3i����/V�V@垲,�5R��c�:�n@0��m���S��i�ѓ���.72�q�_�m�<�,�5,$����q{պ�#�'��Sw>T�r��x�'�����ܼ��S������ �Z��&QV/'��!*��#�+��[����k{'�,P��-u�P�NE;�rG����pߙ��%\�ިu��;28"-d�U |=cV���;�>��f�t���gɊf�����LE��3����@�j�l�gi�:�&�D�5¯צ@Bi=R�r	�{��X?mԮ��{�b�����ah#�K9��]/����+����V�����w�����1�bi�=}1 �3flF=����.6V,2y������J�@{z>�k�;^���OjX��NjO�PE�vw?�T��Xp�x�l6|z��X�ꦋY��+Cɤhi�6:�Y��- ω�*��lN�K��\�u����G3��jV[���Ф#^������C�$�/�q���R�����9@vͭ�]@±�ʑ*U� p��.���ǭ�_th�o�$W˻Va��e�Zw�/��j����^�H_��%�'[�*��=�����+?������s�&MO ���!8��c�;Y�9�W��g��ɸ9�t	l)�S��H�L��>�K��W	�r
`�M����苜����Rm�6L�`���^>�]�o�o>0|\4�� 1K�#�C7��]�C/���i9��˕�l��p��n`y���x�٦zl��~��u�F4&x���sf�S(J�~��έU��^ W��p��6E�PUR��dTS����v��p�I$d; ���K�{������.1hia��uϙU�O����CtrJ�(�19����Ԡ�on���羋�t�9��t��*Ĵ�4��M��v�=�G���'�1Y�"��M�Z_G䴣��b&W`�c��YfX���(��Ut�?�ScrD눸=�_(�|/.}�w/���> ��e�o�{*��!��3���,���Ep��'�=Ǟ�N:gAN���	�(���	�U'<�E(���̈́��Ę��ϛ�0�eʶf���ӜXUt���-v�x��$n�K8���GCz	#T���8��o8U�T�A�����D%�8'��)���M'&�v���$�8r+w���(t$������ö;������*�6�'���LpÜm}�s�AGQ�7&A9(�Q�>{C䢺�6�Ho�Q��6�� ��Sz�-��2F�G� �9τ+�;��G��L, G@�d��L��\o��LBK>�5�r��I��ʈ;�8ɿ�k�-g�yPT��'7�P:K.Μ�Ϝ{n�&&�ijc��
.���/]T����yz�vNd�Gڈ����o�ǘ�K�x{K�i���C�f֭�x��̎��k'�f�E?�W���ϭ�ټ8�x�}�� �����\�2��10-�5��ڄ�t*��{7"�O�}G���dNo6F���<��#L��ud.sthd��8骧�Ɲ��*����!�K8X��0G)�L�7� @%g�hx�'e��S�,�ێ'�cʻ�<!����]���EMo���"��5�VR)�s�d,�l��|�sz����L��\����n�Ķ�����u46����z�ل7��A��N��A�7>�ʌb9od�`�1$2@i���_զ�)8yn��]r�*DqP�d�8ܰw�����Ym��vT��
G`!�{�0�����%ǧ2�F�Z�%H�4�/��_#66�<�C
x���{ԧ8�|W2A���}"��dfnHSi֏f[&���p��o��q�NEQ-�,`�*)�jvr��(�r��uڵ>��-&+/�O���akS�|�R��WT�#����g���i0A>���+�m{�2�$|Q�]�dc������kďfݔ[�[��9�xm_qm��E�M�A.�F�+�X�l�S"�����#�,���=wu�߄��[�<���?yDb�d!�u�J���Ԁq���)������$��f�I���C�1'_q�Ժ�N��ᲂ�^qu��^�{/܄{a�a;�B{�&|5UYӽzPm�����!@4-���h��� �Y��Yt8�+8����5� �R�ls%"�z�?|��$�a�n��_��yn��
��ֽ����C��t����И�'�Ȧї�'�׀��ġ'�$�)"Ɩ���f���h)�R��A@m%����ܷ��۶���A���=e��B�RBb�ĚLFM�o�{�cdC����W�Wi���I�ҁ˜XH7#	��qv0rc]�	j�����ӣYtx�����"@7oU��u�0OT�(RU:����Y4�����*���Q�K*�0Q�s&}��uyxd�M�_+��@�����W"9��������g�|����W-b�Z+$�1QI�t�#���1�{/q �������=�x�`z��#0�Ym7�O*��1_��륊h�ip,x*����|�t��.n���.��d'���
��p	�:�V�A�
7�9���%�c�3iKr�v��	��P�l)�,��q�QrH���pr$D�@�z���=Ӂ�jp�᩽Ȁ7�{@��	��Ecf/�:�|����-���_J�Xʳ"�s6Z'�>f�66�4x%�\�u�"1���xo��BR�Z��h���a��Ѽ�R�!������dr/���b�d����ɀo����,LY�!�l����U4���$���3������"d�n4�� �n�t�)��.X�&C����q�KגҵX��)�h��ћ�T�j�.6`p� B�e)��v�*�x���I�5�)JEEϬȂ5�m��;�H�������#s�(L�|�x���pMDv���E��mN�/KC���a0�g��v�vS#I��{�1Q�>K����.�����~��n���	U<�w�@P���Ui�7�T����9��,(��63�.If���yCE����.�-���j�ճMV�f���g�DC��_O�b�(�BX\���bk8���C�x�5�[�)X@�A���@��x$v���>��v�%#��y�*�(���ޘp�$�&��M��͚�y���6���Ș~?��␝.M�B3��a��I��\�A&�����[My�
d)�M�Ȏ	��!��\��!bI*hƜ5���7�E��O� ���No��cy�#tha��)�����u�ƹ�6F��Zrv�x��/?�&�q�q�ZF�en�~a�x�3l:��R����%�3l�$���C�0�q��0�B�aL��+)��bڈ���:O�y�J�2��9��R����s�j���g�M�4�%�B*�t�AR�ϼ\ �퓮5�K�9C�|�J�3Q!?;R���&�*�<S,����B�T#C�u��c����,3��02�gG��o��#�8l�7���"#g���\Z
���5�V$ep���޳�ͺݼ�v�%�� �)��ݤ��F!瘕i-{k�v$�?euÕ���ڷ<�e�w	��%'i�?QSʝ��^$T����&}cϥT+ȱ�[w^�ձ����1�=]�E�0�	 <�[n���j���@�t�k*'��/��YOLȎ�F�5�T+�U�����={�ZPO�U��v��$�t�������獄[��1�{)RB���j��}���	~����6�r8ܜ_DxuD�� K��5C���A���g�Z.�N�4~�rԌ:Q$Zrȓ'%3��"�9�7�^�Pˡ~w�7�{���|���&s��A����
<ǜ}��O���0�ԓt@��&zc[id�C�mΙ���U��o��=�?�G~���L��_����D:�,UE�w�_�K�:�j��u`���z^���J��ˏ�=���9���up��>֥�ǖi�(�Z�*g��l�׉y��pu�K%8e�,��?w�������%Z�c� q@�b�y�����=��I˵�i�ڈ�;��{���P�!_�0�!�wk�;�n��LH��M����3����0���ȫ��kX���z�O�I���E�r ���q]!g�-#�{NL�$_���M��l��  �"�.�_�_�õ��b!��i7,���B\�g�������>�N�oq�����KAƭ�;j��&<�2��_D�i]ec%���%��*���O3�6�	F!�D�K�z��,��� (9�<�&�}�|	��"8���ҷ��-�W�Q�P�R$u���;w*2wa@L1g�h�����gBmT����Yo�U� -ZĠl���iD%���e>$g�Q������Vl/w"`�9��k��B�>גZ�z��1�b(������wB�����P˚*��
�v\� ��S�pY��!k4/�f��+Fl5���ai*Z-*"���G7f��}�R��k: �O�?�Ի1 ��,E@H�xS���� '�d^IE0-�qA{�dVE���G=N�=!��碋#7�NA���"����g�KB��;���!��^m������M���&`[Bȝ��7y�3��G�o%sbV.5R������������9���,��
v�Nh��J Rk�_�X�i�i�J]���; ��h��v��`j���bF�E^�'o�>;	��蹴^7aP��JT�C����a�&J�_�v�H��̂5d���bO�	鬫��٠|��Y�*]{G/����L���#��*�ee�f��
�Q6l������,���ө�%���Ғ��rr'����00�ީZD2s`Z�Ѱ�و�˿p�%���E
ZU�ɱ���<�C�F����V��lop�5��	M�c��i�3��C, �^\<�T{�ۦ��&�Y�.S��qm����6C@$~�6�3��zt�Rg�s���uMRP��Zt�I��u G����d��L�"c�N����Y#�2Se�����v$�d��;�����M�~vOt�bm�����\ݟ��C�t ����;���6Ul��خ�[cgn���P�Nj���F����mu��:i@a�_��'��\�훜��NJ��S0"'[i�
PY�6s�W%��Q_-��ʼJd`��_22u�[����ߒ����䯒�P[j��������e�3@��A�拴�_7����n�����R�ʽ�ٶ�"�^72f�{�c�Ruȧ�3'��!��Ɯ��k���_Jh�^3����}E���;�sN��S�p6�2{g���,��Ѡ����6���X������R�sX����)���q�%q�tI��W��P��0��@��D|ZԲ*���~� r2�+7�o�U3r�	�����7z�c��q���u�K�4�]i��Ɉ��<k#�gG�s(���Ȗ/5	5�5�Ws�=s���È��~O��h�ƙ�A���mӬxM_�c^/t��~ʹw���!\�#�-��
iG�O�b������m����q~�-���-kͪޅf��xM]��۴N,hqk���4��-4q#m 儮�y��PE(�(RC�@o�ֈnᇶT�裏|�ОN�Vw�ý7݊�K�D�k~ي3
WXv��[{7-l�Χ%�Jy�4����pT�AO|����bea ��?����IM�Jٻ�q���x�A��~�֖���F9d+��rY"�\��������&�����TX�t�!���r�1w�gu�}fuX&�������S��Q�Q�r߳�OLn�W�����+U�|cfY�R�藳���G�T�u�R�:
ô\��J�ܪ�:�5q�"p|g�ľ��=����K����}�⪪���RZ�6������&�1ښH~?�с�=���:^S��8U��</o�\dMT�ڟ�H�Y.2����tr��W�����>�T���*$�����9/�G��咙q�]1�H����7��|��m#8���O�2ž��"�����ݡU�"� �b�nL�6ڿ*%��Q1o�M\0F~���{������\�f䭖��e��ѫ�RB�L� �Uq�����_���Qo��Zp�y�� Sfr��094��	�?tmN���n��:Wl�!�w�:�L���0}E��!�Ee�NGi�1탷?��7�ѓ�j��b�����TjϴG���e%u�]*�;|��_uts�jTG?����xa0��jb����[(6�.ۦ�y7-l��O�z{8�M��L�����`���C$Z��v��M��P��������"�����ڣ����a�ل�����6`�4 Eۙ���/��X��U1+�TQ���T��⁙H�{�b�oA,������%u(u���5�Sc��-� 	��h�C���
"����$$�ᡲH��K��c�W�k����7Q�����9������(�1�VR��@�j>�t+>�k݃���eK{(��� ��ը6�
�	�'�Wz�il��L]��)��:�[}�/��A�b�����)r�'n�+;r��4�E���,�tc=K�0A߇ ��e�ӕ�����h�$�!	���?Z����b�̞b
����,W���|'��j���ǷA��0�ғ���T���t�m�BL5�f�5�$;��}��1�&���6$â.7X2���H�e��ݠ��j���!s3A�%�] ��y�ȟ6C��θ-%�?�ǿ�lU#��2q`�Ɖ����&��O���6Y:�{�Ө�n$}��	����7rU��淀E�ה9�G��?ŋ/
kĪ�XUq�Er!@�L2LRe���(7`���x���/ajlh�,	g/�`w�4o�_�2x1�; �S�<D3 =&���`8��q���}��G� Ȉ�:�r���N����@��<T�����T9�ԓs��u���,�Mk�6y���*<nnP(��9��tY�A�\b�?&��T$�P�����J4[�v�Wv͎��q�*8�����o_p6�v����v��B[O\�]��M��mD��#f�bD��9
to���?M�pD��x�s���fs�����A�S�� |w�13���JW�]'��A���Q���/���z��JJ�.<tN�.�Ǔ�g'�P[���}�%�kD�6L|����}	G2ʶ���o�����������n� M��R*�f����tU�t� w$֥���D��͑�n�K�:W� $*�2[%¹EWZ �ȹ��W掹yV�]�Y�<z�����2+�A�j:�Z�˾�;��u0��=�{~��m�2|�G�!n+�B�EeR�N�rۺGw��zI�$�4�K�;ͱ��Ew9$�a�����&`�J�c�ߎ�1@�^3m����_�L�#��Wb4���
i�($��'�bU7����)'�F�u�?0��h⣁ű��5����;�4�K�'�#g�8k{N7�Fq����uO�	s�Li��lzޟ`cjs��VV,͠�)���"妻,������_����2���U���X�_�	٢Y�u�yX�"B��<k�FK9%NG	��>ұ�ζi	��v���l�Z�G��A2�a0��?=�ډ�Ǧߋ�NX��x,Q�V�Lm˒���P���� C���_�ߕ���˳��������W7�O�+���Q�U>/쌿��dҴ��csr�ᡩ����+_jٸ��_��j��HRhp�<#x����G����y�椶#����O��^;���߃���r �w�S6v����������*i��5s L�:�O����2$��|W�q�~\���dl3���ɘ8�Y����� 	*J��Y)���\f���Zتh�2D����Y1@!�� J���E��FB����;Xf�B��FB�3���Z�K�ۆ�{�f�K��)?$a�����#��!/EX8��7��~D2��GW�\h�JѼ�E�W
�b�F�g7K嬮Z
�
��׋��5S:���ÃZ^7�t K`ꁇD�l:���wXj^1qN>F�%K�*Oѱ���ɤ�J3���e�#nW  ����-k�����������~-��|����!�zl�8�0�ԡkO�z��9*����P�Kf����D�Rs�4�;96.�{�JU
o�9�vS������zÝ�r����-@�<�e�okS�>���|O���	V(�;ꉤ2�C��x3z�|L	�xM�u=������j'���%����$�g���-�D�YBSOQf*Y��h��љK�o�/��Zݞ��ش�A�V�|��_a΀��,���#�˫4#�+��8-�2z6f�qҮ�.�q�"�NT�V� ����1��hn7~ܵ����|a��k�ok�vVH�(	6�Zm82�=�1�D�q�e]��k_1rͧ<uX������&U�l�����2?�:de�b���`E\a�s������Bk�Z��f����}�j�(j�ysY��Pb�!�$r�w�0�9��V��u:��G沄�9;����zw�R����D��~@�(�f��kY�Q�������V��-^7l�ԫ�ծo�i��V݅�;,{�>�)�A����9?��Wis6��~w��R��w��`�R������_<?C�km�Ѥӈ�om�ն 9e��T�y�d��8����Z�Q����Lג�-��%��orV��>��;0Кj#455�j_��ZQn!F}-�~����D6J�	��&��\��N(��B]�a�p�$��s�?J�C�3�����Q�h� ��RoN`3U���(��$��*�FnHa)F�}��xq�L���8�'�S�t�Q.����U�2(��Vn8�w��P�ƃ��H�7���2
�
���q_�Gg��n�]̈́b�i��R	�ZA�۲ydSx4������V@��/��TQ��<��	Y;N�"��u+�%�������uӍ��|L�|	�ڎ�!di9n�n�;t�<���I{�oyrz��v�P�u����K�V�s����t�Y���S;It$uS�S<��4�x����L���bIp����'����_a!�*?<a�-��n �Y����a��bM��:��!D�[���`��-*����\,�.{V>!|W�0�HG����|��3��Ϙ���@�z�{.���4�&��U����m|{0��4N�����	��i��ҪEϻ�ﹹ9�Ͽ#�������#�! QGr���T���g������p=�~R��Iu�7:r��e�/����4az%p�@z<)A����>k#s��l�P�]_�9�oѧK�x�Վ�GC�I��܏��Ѳ�V&�<�98�4����`���=E�n�.a1�O�}�E��j���s�2W��g`��w�grM�ᔩ@��=�I�w���<�2����=�{g��J�y5�q\]���W*G�W����`1;!�a�2)B\zBҭ�=����\�'�?za��nV���.DBT�X#%4�A1�ŷ��Ԭ�5�����j4N�+��}��_@>��?V��������p@>O���?\�C#�����S1[���?�8��֪,�z(y���'�P�����`9��͏�za��O������xi�Y��Bz����*)i`_)!�
�[�VN���f��L�_
�|u�T)��B���<H:��)��v4(^X�,�!��1q|#�<�|l_���;V�Q�ua����Ψ��C���,�h>k���KeJk&*f ����+9�O�� {`�r����fX9�@!�Q����X���?�f} �|�^�A�Ց�	�p��N��u���6tv;(�7�{"+H�Ϙ�<CP�-*Q&��A��'��93��B:Il6��F&�a���I�,�c��qq��$�F-��懹Bm�H����׌�ත=�T��0x��Tn�TGS�+���e�<�:���t���*�׸����s�?�gb-FO�64����c=|��LB�v��;[���W9{��[VR�4h-�WĮ�Q�KQJ�G��K�m�Ug��yT-��H��rL�~_��ĉ�CK�0^�뀟����1�V�AU��	�T۹�ɾ�����=�2�0G�	�Y�	��q/2�!��s�gd�!Z�	���)c[�b�Eqj2��b��IUr�����#�\z�P�l�����g�fSn1k��&�i��ʪE�N��A�Y ݼj�B�@�rPT���A_�WΊ?-�]z륪(FJ�5� �$t�2�Lfbo~���ɚ���"���/bAث?�H�����yg��r!oc� #��xB��'[r����$J��K;㕲#J��h�X ���IJ�8�i]W�T�,�-H�9�)PW�J4�b�W�jU6��1�aj�|�t �}݄D���(41�[>�<�6S�ɣ���]�Y|�� �Ġ����%���&�'̆&ѡ���!Gc�!�z��l��3U:�rs��Jr����$�gx^�O78���t��ȹ���O��.�\����v���a~��h�vS �V�\�PO���?�����'x".��Z�w�+"]~���}vT�RkY���LS]yq漗���&�V�~�2Ǆ��u׌5A9�>��?=�3%����Ӗ�����rcIF�ѭd'] �1>��X1���&k�]��m� ��k*I\e��� �	��0�}�g��U�̥ànވ��`hŦ¼Sf ؚ\3K��v�av����K�̈���ǂ24�� 9��<��tv9&�4=���Z�i\o���sk��NT�o���'����@v�楽�d��5Q+7ԾϨ۫w���2uC1���C��w�j3�L;���PQ-%��;�>x�V�(�clO��
�<�����x�f5��C����Lb�N�;{[�i}`��8�a,�ԓ��mUe�*oES���z��I�P�������r��Kk*Y���c�{9 �]�%����\����La�J���l��_��Eø��[a���h>��ً�H_�(����1	<�e���RPKbiW�Q,�F�0v��F/ G�ec���������n]E0����{�gdB��Z��F|!41���>w$�|�, ]��������sծO��}C 
�n�:�]�@&�r��~]�`	q}�����L�U���yO�X4�����n��LZv��0��Dy��ќ�������5�R�R��A��Bƥ�|!u�������s��.D�#�a���ܛD�2Fq����A¹"� ��1l��"�H��Ⱦ,�,DbR��,�WM�!�DX����zNw˷B���b�F�yg2�¾�:	������
�q���g�"�s �A�)#��`#�^��O$��3/�w�+��z���0����L�D1bߔ��t��#�?��&ʫ��\�	и��(�����C�����2 [lSB��;E���Di#B<S"�u���t�w��D�/���عH�ұy�P����N��y��L�7T�?���iQ��Yv�y�/�䫀kE��ͭ#�+u�2�����ѷt��k`
��ʳ�x)� �.��IW����a̼ikY%D���JS�D��"%H<p �)����3�1�ÿ$G�1��jq\<!>���dG����w{Z�q��M�����gc�,at�V������=�������P�S?��H�;�X����k�48L�+CBW񱀓7\��*B���7�6��^h
0�
�m�:9�No�%Ā�H�h��"ɟ�#<�ꔞ^~�_XV���@�I���a�c�r�G|�ώ�"O%���s����N�9J􍰊�	R{���\iSr���ɰ�l��(ҽF�N`{.B�1r��Hs�H��V��@�(0^G^ ���(����� �ܙI����Ͻ�b7o;{����
^O�J�>|�#g���s���(o���=u��D������-D�3l�#ޡ��oe��^�狛TC63�;{��5�<�����pA>L����7!k��@_��F� Յ	o��r��M�}}G1Y
Fө6���"�M떜JE�x�N���e��a�v;}���=+C�k��B�3[����+�O»5ހ3Xs��C��υ_;_�\.Hj���� dՎ6&�A&ia����<��?"�t���%?�*"\�<t"L��@��a>I�#Z���|�쩵h��'�P��� U.�_�!pT,i󹶦�C�u-��e|\�܊;��z0A���6�\'��М��]����
���'�Z;s�a�n�8V��/G�?�xM�m{ʐo�<��F"�u�}9LR��'"�V��Ҵ_"	|d�G2]p0q:w]&�M��=
��<K��j�}G6��%����:k]���m_s�ɱ��3��6�-�æX���B�MɆ� Ɛ��U�K<]!�y�����)8��;7�-���G�����'e�z�{�_ID�3��+c"��_�� �X͋.�f�3g���a��s�!e��z�'��Њ�]����$L�����F]գ�`�q3�5Ep�d�b#��udF��<)$+�@/�J��
�p�k��[�<gz%̸/���(§q,�ÐL��/�� ]�	�EWAh��_-��v���&�Zm&�Q\�{j�/ߍ̸q��i�h�^�\�o;��mr~�GT�߰ſ�ͷ;�g�� 5-�J��̷�*�X�<n�82s�*Xo�ᴇ�ᅛ3��À���a�D2T����Y��8"����͵�y&I����K���慕�~�,�y"�Q�ũn��1m�r�>Q�2�MJ�*f�"��uӁp�pݶJ�%Y�K�o;�t�[���;�C���e������pzۧ�wL��I�͜/1c�m��3�~8FTe�4�o���
rv�e �&J�.c���z>�*CBL��Fӎ����+w�5�����z�{u�G�m�W�M�=c�홣��������㐶�N�O$5�i�1>&P\\��;d�!�_�z,�-OL�ǐB�����X����zn%Qǉ*��[�
�;�?\.u���X� J+Ե��~�.��[=�+����]x6�%�=�s<�!0@�b���6���Ȗn��\5�%�<P��^ $F4ީa�6��j��fS tO`�!�ig�����A�"�U@�rhR��]l~u�
RB���z�[s�Xbm��L��/���P.��M�PX�4�H�O�$,j��ȉ�Hޟ&��/^[4T� 
�o�"7��F����+�����P�����Y#�W���0�.�?����Ʌf0�rF����/���I1c �ĵ�X�[zس�u�>}@*��^�Hs��t����C�O������h�\)�S�ðKDY%t%��S��B����#0�����of�y���&oV4��ޜ�J9���7�[A%���%��r��]tt�դG�J	��$�@Wb� �����p�K�Zq:���:|���E+�z]v���̥�DӦ�Y�.%'���ݍ3,������QT1^4(Jf�>��@L�rH?��ni����U6.�>�IL��CjqM�,X��<�K�/V�m�,����p�9��D�1K�}��ݎ�L���� 
�rnP����9f�x�V��I�ChP2��~�ocC��8���_��+l����;S�SUs�4�������9�d�wm�I�����u��>րu<���4����{�J_�;�3L�I�0�!��V$��`�v ��~2!�K�/��*dL��a�P>������i6����|���v+�#Nѵ>�������J"��s9�y�Mc����2Q_�|�e!k�rܓy�K�",��z1yL��_O�4F7F�\;�����b	:�l�YR��4<b��˅:���]�>Cr��S��ڋ��D�|�򨮭I�<�2�JbI����'f�z��3]ăޠ��U��u.s60S��5��YN�f0���a1���u)���v]�	�c��V�^d�&�?�y�/�I��.�,X��L��*c��D�Wk�n���A�Ɍ��dw�<UP�.f�{Y�,yb�~ނ������=��>s���$F� l|~
J���R�x�M�o�,=C���.�xE+}�Q�B�O[T��A�Q�0 �C�
��K��qbQ�s���!���c82ʜ�=����k[=
x��]Y�H��_4�μ,c<�E!(�chƻ{���#����.��6- uy�����5��u��h
E��ײY��y��sx>FEp��BR޾ʑ89sm�	��Xх��c�8nx.Yu���e��Q���#O�X�f2�m�����M;fi�B+���hu���}��Aο���	�̣oЗ�{&�op�G�x>t	����:��N�D,p_� �hx
~�� FĎR&��@�e�Y6&��mvd~�m ڴr�^:ķ��@9������Z���@lp<��``�C�4m�,vʠ��1M\տk��S�j8{�๯$��bUs�$����	�j��-�MT9����VB������d뛤����݉���Zz<>����yl�n�����j���m��t�n��$4c$�y�:T2o/*m��Ɨ���<Z������8ڽ���l8�G�%#���*1WC�= �=[_�M#�o�:L����lr�lQO�V%��&洁1�qK�O�"?��7�'�V����A�g��7x�ԧ����}3�� '�p��ïo9�R`����A�0P�8�������B]K%ݘ�>;�,�f��	I�G��/�C�U�F��=M����E\������ �)���qW�e1�ś0 >�^	�4��z{x�@6z�o����x�o墸Uq,y��=�<��{��hW��J.w���m:O*o�1�y��z
>׺��� ���ϫy����R��`����i	<��m P`.��*ۄ2�i��R��ֽ
��S�(Lp#/���7�����m�vI ��V4"�b��+|� ��($A�V�^l��,��W�p�{�)��fnB�e�$J�<��/�TD;k����uG�/ՊY��#�,y�s��ݗPݲ��IaW�7sɧ��c;?�z*��y�����>j��Ŭ�12k�7����)%u�.q�<ec��x(�e�*\��F�Z� 4ݮ�8)�Hܭf�i9�T��J��7�[��jG%؜�x���H,�dՕUˬ/�I7ʞ*�I��f#�A�P�~�1��9"�wʀ�@�m�t2*�U_kv�Y�Q��L����M��~�v�a;�hK%��O�ܞu-&#�iXg��(���yw{t��0M�`�L ��ZyTp�.q8��9�x��D������I$����"S�]9�T4F͘j���D_^�R��ҵ�՚:(S�J��ZT@�)��ͲE�at�T�r[�2�	4����b�E\o4[ā  ���h����s/�3���VF.�[�EE�7G�M�AwM+`qH7(�1�'�R���[��6]��������h�Y���D���d4b@B��>�W�M���[�=Q/���K����:�OO�"��Si	 ����������f>4�y��Qp~��;o���Q���ט�ZzI�SԿ�(_�t�
/��]����;윊�:� Wv��>�ȃ�_��i-`�F�s+�S��I0�.:W&ܑ�� �j�X����G��M�6��)	 �I�q��]|��&��T#X@+�Z^��m�2xՃ�{^-˭�M7����"$�rӆ����c���"�9M~�,�|kQQ@�g���[-���Acs�ʂ�o��q+J�۶h!���ŗ�#��F����G��]����,bt�^��^1n4Ӿ�)���s��5UQUl��ڲ����?�����Q𞜇�Ҋ����? �'�F��Z��<�|�@*&'�X���h�#��Z`�o�M4A�L@��WM��U m���q�:n�L���ߏ�������$�������f�^���+�}�h ��t�%F�ן�B�D��G+;���C����.�/� )�J�׫ъ�C��H����k��)<`0N��?G�[����z1�q~�r���r�*�4�7�O$w��S{[n;��t0�YL慖 |�.�[�������+��J�����9��K� ib�~��QH�W/���F� X���hS��������$��#T7�� ]�ң~����J�G����(M�L�s�u�qJ�z n�Y8�|R_,�QϚ-e����T��kk������-"Mآ�O'wo�r��TA!9�:ʣ�-�F�?7�]�a��a�����1i/��l��ө���Њ��o�8/A�B�����,�
�'7�g)f,�>p�^��5������w�z�ʰ9��{�GI��$_v�7` �^�;&'����&��N@G쭍�W�!��jِ�tI�Y<���N=(�ωKJ��ɷla��z1:��A��o	i3Խ)<n�n��X��o�=��;��W>�3Ե7��R]���w
�qݓA�y7~��b��k��S�V�AD.�A���$�CF��1dk�`3�QF��>�[(��h����D�F&����BP�?�NUO�zg�J'���5�;Q�
��4- J[{��|���}�/И�@�O�ƿ�>�8�nb����-��Ƣ�������vqՊ���\/�G�&/��A���ʿ.f搭�(;8<c�!�9L�t�Ks'\:@�dУ
���F��']�~Fˈ�F���g��6�!C���G'ka)���l������Dp��*b�� �uA}ͯ��n�8����k�b��gH�[�M!6w������̬k�)�\�y��Eݡ_�|��ƹ?��{��`ᨛ�E.�Z�4���ـ4�D�����޸�Oƭ�*�TH���/א&��8+=��1��9A5m���i-��e��f [�P�J�f=j�e/va!1�ٝ���c��ZX��=O}]�Jl<�tuT�܍�K�:�(߆9����ނ�QM �F�o
�^b��ձwt>;	���a^Fמ�&
�=�J�geP��v�Oz�y����d.�Y=���&����8
�U���fIQG��Xla�Y���B�;ȗ��� G�q�v�H����w��?C����׌G}��!u��s�,��H�S���!�=��Y��g@��/��o����4ٺ�$~�@@X��0$`�0��h�&Y�����D�F�'?�U���N�$d~�jӜ��jr�Ģ�cS�,b\�'�ф�&�m��>�]q7��l�F^9M���������Ib.���M��b��q�?�	(��|Đ��33P�:߫Z|ZS&w�)�DKd$������X���ƿ�9�zͮ��e����d�0u�>�Χ6n%�W��k�T�KQՌ�k�Е2��Wn�AhqsX�+���T;�	xQɸ��K0�<>c��_��*��p@�Q����"�R�:f�i���Pa{�&{�:�A������+0�~
c�1Ӡ�z�D��o�Y�[�Z�;$'?<q�XH�{T�x�3O�eLS��K���m��2u�\H�>�&������^�'F�v�8�m2��|N՟k��+*�d�ء 47��Hf�y{�0p_7����B&j.]��Ee���Xif��~}�4�㺋��vĠL��r��j$�3�D�SLPA�����CJ���k3��H��e;ZE�1�ε�j�|����Vυl�����&b���߶�kh�wےyd���XȢz0q�)�ԬB]��oE֖D���v��]��#�g�,�����DKN1�+����f�P�	��µ%C���.=U�t��va0���ײ�Wk͛Me����z���4�#�A��ĺ�{vê�����e�i�)�B��v�� +���~zrV[K��7��X�@���Z��+7�3��H-�	���/1��M\����cg*�n��}�G��+S��![����w��0�y�A�y�L����Y1>�7�6��H��㬀�(̼�oY������^2����(��N+�o@�*�	&�#̎��� �Mˌ��6��LpC�=�D6a��p����w��iK�j)�����-5j�^�e��
���XjȾw+�D�Щ2��1:24�,˔�.�-�����?�[�eܕ�Aޟ�p��iW�/_�qt��C�4
�=Y���,������_��jP�!m�3�骫;�<k�	S�xS����}7ѓN��&�%�J���G� �]`�c��U��s��1ϻ��v*�p@0���)��a�0�Y�e���AA�H�$k��,(Q�k��AY?�.'�N
K��>��I���1�f��<�ܟ���{��9��tܱ�q��r��۴�a*�?�Σ������(�$p�.3�Y1�
�� �)`C��Q��`�Z��Y�J�/��6�,�&+�;�4�*�2�#�yǈ�'f�r�E�,"ner�;=$�9^TA���O�7�9���Z[g2����V�����o^�gࣨ�Тhͻ)�+]oeS�$��hǉ0�v좦���~ά�z�3�.�a̳�N�P���&���}�_�\�W��Y�D�\Ζ�7?1�O�o�׵��`>�A�����ML�M�F���6���YL����߶I���ClNiW��a�@��27����q�2=����	t��|�����4*�����.xq����g�?5��&E��)An:�O&�kZ{��8��#_c�*tZ�pf"�J���#����	��-�����#�S��X�9����8���� t�YT�5�ŕB� �o��iRT5�W���xyp����O=�LL�Bh�ci�T�� �5XI�~.t�3�!p�#|Hw5��"O�s+�jo��(�:mύVDY�3�Zv���h~ZE�h�BR�����__8A�����9������"�O���Lž�ۣfM�}��|��po8�kp��QztI��bH�����'�rt���RY��P�:Gę�~�8�s�8���N�?������9p5���+zIcơ��X�n��,,�}/�:&oZ�Y���F5�9�Ǯ��w�1iڎ
s���Q�@��ڛͪ/��@^hVp<��wTD�)���O��k�: dZ]�O_l$�=�P3{�2�AYKL�R��1�"j:�8��L�k,���i�gUO�Gn��)�V�ۑ��~z4�����"�n�x���]؏�Ow�w%[ځ�K�
-.[�̢���d�Kf+N�1�b_ȴ��&�
�s�� �'9��k�x۪������$�36�wJ3D�#�ĒMK�Q�:Fښ/���k��az<�+��Vy���l�rRbb���=�m���`w!�����v\�]2d��v���M〲��P�:��g(�E�޸�#���'�{C��Qo���ns���ݭ��/G�c˛$�KUf;%3Iq�-@�4�ɥ�xf�ں�M��jͦ����n����#��n�r��9���N
�\l��bY�����:Xp£����Vm�S�|%�i������9�*�y��VS��HmE�s���Q{�QA>�e+w=����/I5y)�B�nwd�_�MԬP�����$Z������C�Vt9�z��)�>,Wh�x{7��MN�_�j�_+�����,�:ݜ�f�O'P5Gyj��{� �i-��Z��3L���$t�shx�yG݂T ��B[��zDٚ�Y�*<&1w�sB^y���E��#��״���7�F~%�
���GrbGQ5���Gd����C�ف�B�9�9D��Ė�O���}�p���������Q(�\��'���/$��x��/g�e�UK��H�ՁF��Lf�*�ׁ>����E�TҊϬ4Y�ܿJ�e�F�b�\�Z��	D^Y�{I}S�ʳj`]�G�����4:T_)������������^~��WZU��a�dn������UAi[�ĳ\�&g�~��:�)��
_���Oe 5R?�T�� ���ț[�����[�$��� ��������`%B�U|�U꨻��n_�H�d�ƠZ$p�H
��pf]IB+O��K&	�X�G�؆�f}
?���|�ꉡQ�W[� �Tg��g
��<��_�s��t���֠���V3����ˣu�V	����;����h�F��,�s�w�s�/ѭX�a0޿�F��pU�.!N������_b�H�h�E��:
T�:m�fDQ���@�����:�\)�`�==;�6OJ/��&�i������iiӬ��=�}W����)�$m�,�C��*�[�Bb��%��Abka��%����C�XE�u�L?��p�uy~���\��"�e�L7Ex�D�Ɖ&Y[S��A��^i*)��5�#(�RocT /� $\O����v;� �T,�΀�Z�?�ص&C�H�'��o��O-S���H�t�}��Q�y��"'.���Lr��	��m��y���@��3��j��<��=����:������Uq�WH�j�p�;�pW�̀��Tk�"����T���d���l]�W0�cusw�N�h�N�7�O�� Nk>x|9��`�EQ�bU��X���r�Ȏ��x7o9�j��^�Z,��|�=�$�
��T��Edl������@Զ����;bJ�R�N�]X���/y �l�$���F�zTݢ�%����,��3���5kR��ď
;�����1������CN.@��,-�0c,vѢ�`����c�.��Q�+���T6�7r=BF�-f������/U�y�T����4���N�V�o^����h)�`z�<��O��``���
�Bw�+�6�2l',�m(Ch���m[�j����o��t�±3�e���yW"\Oh�$Fa՗�����s�=����
l��񮗗� �htl�ο"/�����'�E�#�'s*R�:��~��h�L#�ٿé%,Ȯ���!aȚE�X�haS�B����	�x$��xjH�}��g�;��H?rdMM?�AN�sL:�P1�i�{��m͉�QRS��փ���a"ec��jH-�7�nCx�����Sky�����Z���[)��/�)�+[N0u�[.�w�U���]N�k�N_��m"��+&�������܌E�P��{ױ\�M��Xm2"�b&&�u���f�Nx ;V���PYO%W"g���ӛAV�~����ֳ�؀��ֵ=�"=?�	�Ru����,�GL��ӽ��l�@G1�YJ��!���Я���fn����Fkxa:�R_i��w,!�J�ә��0߈��M��e)�r�?T�s,�6ҩ�jNs����ѱU	( ʐ�^��myk����/Ψ�Qs���O�$�KI6��z R�����`�0��t���a[�$xeH#�2�E�B�#�� K�a����p��-�Xa�K�����s3:E�hv�,�	 ���Vl��QoSco[�4:�O�L�\c�t3f���2`��n��q�I�'�^�A;�ҷP�L�rsk�V��ŕ#����e ⠱~PG�j��^`t�U0�<�1��!��+�G��36S�T�o��Y����yvd�b_pZ�\_�z��#W_@xe��!j(c]�F�m�W��"sÌ�/�W�<��Jj�X흗��򷯣�M=Rzp�s�������|�l��M��'��)��{�ΒK��Ӫ��̜��Ku�P�M��� \?�;V`�#�=z�c�M�7n�ϋ��������+��MQK�'4��~��������n����O1@���6�hl[Ct�/~7���-T^ #E�����{HU���D���o��J�W�o�T��!d�ŕb�3�˚����#�c�A܂��: �5����~u�FZ`��ƀ��v���{�!���`�菠l�>�����Jp~2?e��(G������ގ��M;�b�������&ƪ)�;c!�;/V<"]� �m�g�|��r@2w`�ȶ%��T�AjLzc q��h��;���|���f()]ގ�Enљ��L\�Dd�1�m�:U4�y��ĝ��(� ���F�]��tƢ �%`(��C�B ~q�Î&��ہ%?J�xZ3�(|��=��4���9D�_44P���`��.;(�\O7aycɎn[��,ԝ�)��q��6?6U�d,dd����kS�@!*4����1���(]#X�`.h�75�ӻ���	�EM{������CGG������f:��mV2VJ�pxK q����.+�SA��2n�m�R���qq��:����L�e���)��q�1X���%w�nn8���7�G}��L 'H���<0�ɧ&�s��}�z`	�8/=@�v���CA[{!�+�e�\C�ǃǗ`M��?�JOE뺔���W�WQ>�̎�P�!������υݍ�d��OēP~0�k��F��$�&@�(d	�2�o�w4�Y[��$F�ed&�WQ���!�gD�GI뱐��Q�̐�z1N�+��
���K`�4x,a��>��]'d��P��D�덯K[!6MBvAaʅ�]k+>���󧘕�{p���#a��q��ȗz���Kp�&�kj��.�2����{��}U[s]��1z��H/��G=?,�����u�!o1rd%���{N̵��=��3@�%���o�&<�O��}e?$��ߚ�;!I�د�}#������{�c�*I+|~G���P����
&g�2`�u�X9|Q��{D�uh��
��|'�(9D)����xt�ߜw�:��Wض6���g=�?�]k�4��-�k�'}�� �f{��Z]"Yl����}�@�����T����:�s�eHL��� �x����
���`P_�*yhIƑ�����	������'�o46u�����/���X+K��`X�b����2�.�������'a>K2���RP_���Za�!=e�Ig�@$z)�h�ʱ[�&���x�f$R�����24�K����:�~騆^��&ļP��m�Z��M��o���'�4{�ӊ}70H�z�!�j� 4�����d.�ɳꏛ��'�22W�r"�@oeJ4�J"X`�'���(��h��6�QNxa��ٖM��iC��2��x� o}��E�����Iɭ��)|_�gǷ���(ܹ���År��6mIK�o�
o8%���~v�i�@���~������W"��U� ~�!sC}}�{/?W���FR���k��9��5�ζ��}��ض�(��S��!ض�?_��J8h_K_�54?�xoqc��+��9�x�̈�����W�0:��j�j)NW=>�\;��H⫶w�pf'�ss8��R���y�B)���(B���H	R(X����jT�Å�	c�=�za���N%a�lVĻs�E�6����pz�ړB�d_�{n��JVc�<f2��"o�p�[b���Wkx|e@~fϾ�\iI�OwP:&���`��}L��i��/$��4+�)�G��1�v�̗6?!�D���l�%�����&,�ꂦ�������Jy�#�]�H���;�60��}|i"N1'BH�~Q�Evc/�#)ywr��{2�<�����W�c1�p�~�6��	�FJl@ l���V�G'�j@��^�E��zI��GQe<��uj� u��4�Wo�Q�/�6�!z��q����|�BiB����#�d������<�WpS��1.������)[b7C��Hޅ"NX�A9,�C����ڕ���Y�_aE�W�������ĎL�'`GsQ!�����U��0�1�%kd2�#B{!�;�>9� j�v�.~Y�?��x�%(6D��z�ה!A31#�p�	���$���� �*@�~��8�V��3��U�4}��?�"�^˥!��r�!��`6۲�Z�	#�������)�])k�k�x;_���^��D���6A7�N�Z�E����}��B�)�����E�y�Jh��c����b=����9�J :�
>�8�E��4Xy�P2K4C�uwJi1C�M':x���W]�gt�vC��p�p�j,0VV�w��[^��f�b��NS{��u%�2���:/��}��_��:�e�,�$)�8L���4�h��uO�'5���Z�1�&a��E���GNd�j ��Y�sX���yPT�����e@�IW�S��o�s,�B!�|=�E�ǜr[�`C�1բ#�"�TDF{��l�7�fe�2�4wa�Onn���Қ]�T9�_����;��"F-���Ҙ��P�E�K�b*���#P�oeȬ��ϐ�ٹ=ؖ��k!����w]�n^���ҽ�6ݜ#��i�y��$�0�+=8�4���w9S�id��>���5~pRϪ�7�U$�Iڙ��'[�r� xp�*,��sB�����U|l %�v+~�H�"hŬ<�l�4tZ��!�b��$T���G�PĒ�0Q���O��b>��d�6�3IW"��,���qڵQ�o�.ǳ-��˃�<C�"g�+��_�{���\=7��_�Dr0�ܭ�ju�E0�;�<W~�"�M��?t?)����
�K��X�o�l���0
 ��tb#C2�`����##y�Δ���G�:�}�Vu��EZ[^ý�h����p<Ǯ<jz*�b��~��pwh��+��3ۅ&��+�����"o���a�&g�N���ka��tK���O2i�y&$�S} ��O�G���Tv���M�-�^�_���1���lN��ݐ� �}�H�M�-� ���"`Ӄ��)=)ӓ����9��&��E��bp=܀�_�%��2�'�z���2xvi#�p�
Zł���n�k����[�8A���m������B�
oBxPBj���,�~�s��bjҬ���l��u���n���1ȋr4�.�$��Ϲ7�!8�T�	�k���3 �+xiج�$�覱 v:��u�H�Zo��� {�"�^}ս�\�٘D[�=�6L��Q(�|�z�U�l+LX�C�{�D���6�mz^8�y��������`���y����׀�f([�x�g�:'mɝ�7��m��6��J0m�24V�>��+�+r���!�����B�`60����+5JN5����'>6�������i
��)�����u��u����+j�I�4I�@g�u֝k_�JQ'��������0�'@���unC�5y$?��/�0�_O;(��Ѩ-[.8���^��
�ҢeWd���+�8�\�1�E�/�#l_�>`r6�So`�~�F��^�U��J<�t��}������viq�$J�_�c������:�MW�[�ʿ\`����&�v�i@n���|,z6Cp��<P25�5Ù/�k%�1f,�פ��+��-�942�Uq� ��޶\�a����Y�~ơ�J7 :!
aI,�`��M�����U���'��4ʰ�Zߍ�F^��0��&v)�W�K�-d�?yM�5f����L��V��'͊������AFDGy.����M����N󸜼,0_n�ha��F�z�O���,@��{�76���2;p�m7���D4S����m\���vG�����͕8!�zU1��Z%�n��
cl��@���İ�æ4�\]�.~C���X]!_�k{�	Z��Haq:��S��@�0(�V�T�����aCMYʶ�s#�}��Q�� �eZva+N�n#����4'�����j�N�pF���J���RZ"�J��8�?�9�����Tl��T�[��
I�O�L$>����z�y�]/��(pm �gȘ��k�Ƀ�>WT���?�F�yhݓ0H�`���ϊ��?�>�,k}wt��z��M?����>��[mEio��T��d�V%���J�()�.3eQG���%(yP�!n�a'S��SN�4���\syQ�ɉ|z��8Od̝u��Z2㰽m��@���kz�ܖSZ�bQ��L(�K��vc+q�=W��lQ�s`���.�o��A�����ϢEZŌ���t-7`�.�Z�|��fd�3�Mhl;Ëeq����W�f���'}�#�(�W��G{�X�V��Tk�Dq����u�d'M�v���r�nƩ�'�"�p�Ww,}���<x����,}��[>?��r�\��l�r7������t};��
H[��8��o����>2lR0�mLJL��Z9�Z��C.��Si��;d�)���Yx�!mX�� �&{�M���
��F����Ym�����Ծ>{:>f���(kZ^�k?.?F�'�*��t��
]|{��2�3�K� _�`㻰�y/��`̌��wHvx�2�z�$�mO�j�����K�>�8�_�Q@Ap|�+�6n�\\�n�x�דA�,��Cw?���9w~0�F'�n�t���6
pfU�S�\�.�A�9��>�[�gJO�
@��R-������cT;j��ތ���`me�^c+G����?�3�z��J�>�;�V��0�3��!;ayӣ?bm,�ާIreL;bkg&���O	WU"0&������yi�[E���S�0Q��Tȁ'q�Ե�s��D(�^��L������p�Ùi����쉍�u<����S~$�����<W�8�z��#̹?J@��v�H�r:��&տ�r��2�]-vg8ߨd¯]���:O=W�(�֓埣r�X��	GU����^��������OQ��w�2t���h �W���nܧ�L͚��w�∂%�)\���"���
QC30�3�烦@fm~*/D�z���ՙ�NBC�J��8P�B�Q3����<��6�z��j�c�1�L-En��_��� �qo�c�j���|�!������p)��fԅR �9;��C�Afq&WW�<Y��<j�<M��ѱr#|��,Mz1�/��`	WޏR���l���8�:���
���Ʒ4�~!����Uf�����ݿ����J+�Z��P� ������&��P��<~j�J�z�|�7ӧ��>�$ʇ���ꤳj�r@��M=6��[�%��5E��u�M�|��	煈� ��EJaZ��{V��?��Sm��!������AQ7P����I�-�ׂ��mc{��(<�^���O�����l��;v�\�/Ǌr����0�T���_I1��1���<7�����s�@��M���@b;��N"zȷ�p���y �h7���� s��(h7�f
���M���Ln�RQ\�������f�Ϳ�F�홃�z-Y%4(n\��	)&��gh�(�����m�����hN�	J���GPg)���c�5��i��z�)�y�]:'����61C_�,]x�}�I�u�S���c�,�P��Ȗ9oZZC^-�^� ���װ8��@��f>e�"ˁ���:�������Y?���2�h&�����pg�h�6�����9X|�MhH��V�������+�k9ھ����vś�
����h�,�| ���	�����`l!���@2#�8��êL#�'�r�!T��`p(Ek�&)Qy�k^�cĚ�i+R�G�����
>q�#S��V!7���N,�gV�h��˩H'.���+�G��W#�����D�_�Sk�¾E-#5��܄Q������{r\t��5bWrQ�4x.�(//�1�C��n��1�VMӖ�>Y��V�[�<w�a�O�2�7E���ہ&ڈc��I�3"��G��iY־�!���,���tqp�Q�Z��\���Kc��~� UU�hq��I����6�/�iU ���=bt��]YIW�G\���/P��z-ף��\z�p&��<ƶ�����n �h�f_Q�7�t�u�8���;n|���{����WQ�Wn�L�UFg�n�E�⼯/^]7?xT� ���v��Ravu7W_�%���[}*6�Ҟ�Q��.͉t�!�QXuxT���()������l�d�_�g�U����@U�G��-�Lp7��0\���e�#�*C��\����Y#C2�%��c�l�˹0�SoAG�O��代������~��Z'k���R��|�j����I����
8�U�{ �JGX�~F�DDG�=K�/O�Mnd�:�,�n��;5F�9 ���7v�ރ'����8�q�W���!"��B���p����1b�m�\ߖ�`n+_}#+�rg���h�t�5���D�ث�ϲ�S3�'@��������07	����{Y�cM��Q��f'xU8[��w磇�a����f�p)\n�x����9�q�%*�?dI�. � W���T�7h��au�����2-�R��(����&�~$�.
�.a�Oa���b�][W��
����!C���1Ѐ�N�	��4�@�3��N��2��Z�W�qP������s:�� Irֹ���6�j
�)�r�ē�\����o٬;#��-�E*h�x� +�P��	�d�-��畚1���+k�
������J�Q�;�``������?8���=9Q�+���w<LԼU�ތ�G_)���0�|x�������Fz>����x��265�R�~���r8
y��!�K+�,އ��y\��T3�h���LJ� �@�<y�?���/�<�u+\'��c�IR1�g�j�fG�5���~��V#j��Qq�d�)���0�M�y^¢Alma�P��<S}�I�*��pz\��,��_������+����P�G%{�M[e�M`g�K�K5~�?���~S��<r��숿�kƻ���!O]���(���-U�W.�_(	�G]&�v���BdO��|�e������'���T�Ui�gƸ�!	:V8j3"���>#���m%��%'�p���)FWX�(� &O�B�"��"�(��1|��7#9�ʯ],�t%WH��i�#Y�},N���(�2ݲ^���X��G�o2+)x�J��)Y&A�����ݳ���v�Q���.<2
�;a�����mO�����kn��;�Űّ���C� ��,!xC"�x!��L1����T6{��ɑHAӊ��}5$��T����W ��d�	���3+_�����N�	&��!K�Z�s1�]�F)l�k^�љ�+,��SR-�{^\c�wl�0�Z��ʊ �'�b��U�����~����#E-�R�OK�abK༴�����W֫�`�P#{�1�w��v���� �Y��&�u���g.?]B��N�/��H����zLB-�Þjbo�Mu�!we������FEm;��~(�. j$�
S�K	WLղ����K��qD>�R5e\��ʔ�@In�,f�hd��lS�Ě�R��	s��5A;�N_?J��-^>�}��r<b0��%B�ʝu
�yŁ�V(�.')�mx��r�,6�ZF�z���R���)�����?n<^�D/)u��5

�c?z�$6l� }ٻ��'F�Jv�>���`���Lv��85_��Oz^6�9��e�A�'ΥgK�8J,�Y����Q�Ъqs�{�X�"��ڶ���"c�r��{�M��*d�ܶ�����U^9�/^arf�K�G�V�=� I�����b��-y��۪��`��[9O �s�C���(�1�]t���7��p��6e��|S���s����}���k�6M�ʗ�O
n� �*��n}�}M�T+�O"QJ�������?嘏-av]�������`h9�����\�H����	7�<Q|�B6�؁�Dwf�BQ(�xӃ9��@���?���y����>k@���O*
ߔ,�(���	1�WYH���6�0�,W�仞i�pr)~�N�T��)Zf�K���c�>Q܅e���»��N��t���Vq���.�w� �m��a_�vi�#�U�Z'���l��+>���j�L&f@H�\	6v�$v}ޒ��9���_�č���Q��ق��xכ�|�	05n�p9�p�V�~�&������"bD���`��m�`��8^��dT�7�*XHe�'~l1�$���r��B��U�AqE�]i<D�r�T��7 KU��29{4���x1+8<%�
7
y ��1� ��'�Ū��ަ�yy��)�Ȫ��7�����y�[���&��l���~���K�בKZV�� �`�M֙��U��:?���i�fz��&��љY�����k����Guθ0����������=��(��?!���m3��w?��^�悓��/��v�WYo#=+���ǌ�եQ��x5&K݅���N:׳E��IJ^]��kJ�|
>�[�H3�ޡI�Ͽ��]�M� ��nM1��hc&�G��r{c�|�U��V1���-"E�B���/ɰo:��W�40:���3IJ����oq��.�z�^�@�RF�<��/N��qGX(�,�������C�<�ʮq.�_�O��Ohpc<�$�T�L�(�wZn~����F��
3��x2}/�b�~�7�~52���Z���4������-+;O/ܑ�ߥcu �UM�˧vz-�j^`������Z��s����Ù֡���V@�ѕ:^�˽4�V�tl�J0�e�+ly*�� �0��M%�긋�I7��΀-��D�/h{�a���PO�a�����x[�Q�B�#o�y��r1�f���2��W�m�"��`�G����ȫޅ�1*�7ߧ־�m�0%�.`=e���3���h�s�}����d��>Ǳ*apK����?&�w�f����_X3�����BwkM8Z�-���`<�h& Ȱ�P�R��h|��\���ɛ��v�t�\��O�7,3��>�"�@�p���Gb�'����`�x"�mX�b��-��+�u�`�UF�x�ۂ^K��%�b�/#0c";(	������
єc�\��� �ń�U/��C�#ЧC������*�9*��lQ��h���t�-�	*��qz���#����'1Way܅-.���HP]=窽��|�3MIeQ?��P}��>��΃��T���@?	R[N���OTXe�l4������g(5�JD��Qy��~�P¸�=vо	s����(�[v�}���	6p�7����CITo"��O����-��2rm��6�!����i�Ģ�i����S½s�y�X���߼Y���;�g�1�����\4��T��*ڙ��.�JI�+���gj6w_������lƖ�zÙ��Qc�LX+�!rW�G���ٰ�HM�?��"'Ѩa�������aH����r��4�Z��c0vl���� >�օ��-p��[tܵ˺�9��O� �/Q�H�Z'78)�<sݟ�����tXW\�h����'�Y8><g���R�X����uW�1W�ZX�|`Jv��W�A��)x��ݷu#`����
�"��d{���M^@YA?-��èR���e0��B�uz	�w�i_1��2�I�l��}�?����l^&���zA\�F|!L`�đ^"�=��,���:�ۨM��p�2%BcO˺+Y(}�D5������$P5ߕ}�]����a��H����b�^��I��U�E�`��<����/���-��F���2T�_�nlj����%��1S��KT���jG�%��D*���ՍXh� �i��_nR�ӸR
�\�6T΂]#��9�.z�
~��ꅽs�j�"8]����B�+�}ni��~BQa�50B�v�?�����W��L9�	ta��-�P�YfI�@�ގ��ȁ�G\����ΐ���M�u��ED�x�<YL�)ǿ�[�оP7)30��v)��F^3̈�`���jV[h�F{d���uE6|���V��f�;V��(�,��W5W�E%̎�8k7OJ�����ټ7���`G_<aI>G&�DGn���~?��`��Q黇�;�#F�D��p��c���2ln�>��\�JY��g���'E�?�¬i(;�7"�}�c`�=�ε���e\t�����^�I�{��G��K|M/$�˵g4�!id�!�Ci��h�Y�^i<�E�S��;?�T��V���g�0���LS}����|�^�ɐ�n��n����9��C�2���t��{���!��Yw�Ƞ��՝�4o4�+�T�h| �,����F�1[o+����'�b(�,�<>Z.o�Q�BYV�N�g|^{t^r4�C��6Q�2vK�a�e1\/������٤E2,�P�,��x@�4���ᇵ�i/~B��;-�^����/jY�S SPR`Eؕ����qf�`��.���WnV��X��ן`����u�z��X��~����'�q��Ƨ~5��>��ڈ*��Py�}B��>YV�d]���$�5�-L��
w-�R��"5k*��q*�6|(�??
qT?`�Ľ!\�pYv	0�h���n;�,��Ve����>c�q]�� ��m.����'Zΐ��^w�܏�F�`�*��=]��/-�iQ����i�����C�W=#�e�F���e���O@������(��1�I��v��Z���W��i����7�m��,#�O/�x�D�Ա��\`�p+��Rcxq>�i�糧,����a%�e���G���=Kʲ�$���?;�X�B�Z%4�K��_�~�Bw��nW�1;�	�s�:����~�@}�v�m���{?;�"��@�y��[�c�7h�y4W��s9X�*�N��e�_��R�Eϩ$��p�|wK�ER�J+�'��!�$��Ś�0֠��� *�H�c�q��p�b�)Q����$�֤��^�r:]}��J�YE�t"��d���F�7�|�g��_/A��W "���U��� b��=��~X�h�����0#:*I��̔&���}۠W�A�C�ţ,��7�C���O�v@�H^�=��m�Q(֠�S�f���>�"��:X��$�a��L)��Oj��
D#;{6�١��� 9G$Q;�R��0N����c�4} DB��;n���yB�����J�\�Ǥ�UlƑ��Թ��\�s�u�5�n,q}9E#ڂ�Y��GQ�q�U5sT�;Zx����;��D����/�������Vض` �����6�H7���$�܆��&𙢣N��o���] Pe�9�!��92��
4��Ŭ��B�x���d��ȻzX#>�~��SB�	������0�Tr��E�-x}�-2�&�q��"�x|�@C�b�ZN��M\WC����_�ce4���j�}fͅ�]���盛=)��	����<΅��9�<,��8�Ϲ���~�;Ly�"]A,���!~���o�&�i- e����) +>��[y�x�{p]H��\�2�!2C�FGv�ł8�L-�G�2��>?F��Y0�}�Mmn���f�	�(������� KK�"1�p^�%�Qwv�2J
��[��f��q����C���u�	7�M�
��ħ�I�zL����1��ZL��T��(Q_��o�0�.(Sl%�G����UpЗdt�%`\��&߾~��!MF8 �}��i�I�����1c|-�y�w���|=�� �sA��Y��p Tā
����d(�*43�[c5���D%�= 3zޏ�G=��̒�8��ɔ#��^�H�S��$ރG&U�(��y,��I�.���0������7�vj�ļ��J��u�{���5�	)�^3�4ڄ^Na��9��K�|��bi+uIJ���0�*���������|�������d��ㅷ�kT��;�n�o�#�r5����m>�%?j����Ѿ��ا�!p�:tc�k]�dM��{<<2/|���]�j��'�
<{�<�0.'�f2e����!7'a𹊕�7����(qÝ���}7���g�$��w����%
X?��7�5ʹ�2҇�����&RN_9�'�2̚j����u$W�6�j�l�}k����1�q-L@h�����h2p�?�D**(y��;/��:h	�$��D����#���+8
<��֏��jV�<�[$w�h+ZJ@�5z�^:o��p��J�6�p�&'��a�GjT��Q� ���(�R�7��S��OX�����<8՜�I�)�YF�Z���]�J��;)@�N�br��$�|�eb��s��ۺ|�W�t;��#��kx��Ǧ��s�����ei>y������8�����*�� f����,�cckԼ�f���f�Ѽ���d�T��9�.��^vM�b��o��!����]�g^��B��"qS�&/��I�a�XfMɼ�Yu��̗Z{X"+'�7h�R!���̴r��U�enKD/-�ʊ�@�OX>w���(����'�l47@�w��SL�] �Tf��z�K��j�>"��i�]��gHz�s.xM�,[�)�!?ᭉ1宷/G��tbe�^��>ʖ�I�so�2�W'f,_鋳��˹D%Hm�ʘ���P��,��P���>�i��NL܊�=�TrKP�_r9CDgm[�&U8�i���g���f�� ��Y�z�"���}���]���������h_��
�g�D�Q���+���)a�����.˥��g�ٻ���_���Q�9���ŧ`Ny����z��)��p{ mI��ǒ��H'{�B���:� ��WW��ӟ�	��bM�?q�c�I%���H%�YawtD�����_�'t,m_d���dd,r'��D�,XP���p�� u�yT�0�y%J1N�>V��YAj٣0 Wh�����hh��<&�5��-�+��}b�^�EWa��ӄ�{��Mz|��c��%�XG�H��N��6�����>�Iy\s��ل����Q������ʳ����Y�T@7W�du�V:
V|zf�Fu�|{�r��l0�<�ʷ�����p�I�OO��
��d��o7�yA0�� OK#_V�噁�!tٮG��1���'�n���Rw�d�e>�O�/'�����P]i��EF�C_"�Q���ˢ�9�9���ܾ'���Z� i��J�-����K~Z�m�K�A�lEY�K�	���q[�Q��G�}�����La� �;��������mXoF�S�ǹ[ol������7k "��S�苛O���%�ԥ�Y��B,U�})5��?kk�����NXi��`�ݴ��%;��-FYL����+����/1�{�K��,Q'ޏf�1;��p�l�'�ӌrb]^%wEa؃���m�NJs2�|n���G�-�b4��o�s�����~�������m�׎��9��Y/y��1�[��R0�A���%���kx�Z�=u$�7�l�T(�zw��)��Y&؅ȯܨ��o��Vc��$w����w^DϲB:�F���f�O(�ĜC
�ϋo\�PdvG���&;�,�s�*���S�][�t����iӍ&J�Q���P�|`Ȓ�?�#S��>�E⌋'��+px)��R�6{�߀�j�R�2�/��d�kS����_��?ԯK�蟏gӵNt��1sV�@ Z5�$�b'&�!�f]�/p-��J�\.۷h�|,s��Ϗ�)p�e9OI7��ʦ���Cj��9|���:X�,O��!�������UY�]��ҸlN�dCMe�Sh����-� ��<�!3|l�����)�������>�￷�t�����e�׿�	���m�`�PXj��lS�\|���6)� d�ÂB��Ʋ�ͦ1�W|�`���PQ����W����!��A@x_��@*��Z�'=� ��<�� Sе�eɭC���I����,/��;��)~�Vu�;�t]ǩ`T�%	�'5�zxҙc'�P6g_"�h��~�k���VY�m��mSPh����y|�����DA������.A�|��V[GNi�X'�m���}���{o��TCce�*�.��T$�ޏ!�'��,��܌)�k��ʐ9�LB�+Jp'"<��͒��L/3�ɍ�h��}^~� ��	9�b�N�����(rܻ1���_>�$����iUI���z-9L}�QN�����tr���hN�z����%Z7�),b'
�q��i�i�����.G\�$*��Z�#U����\��[��db;.B�.k���R�n戤�ןڅ��(�j[˩��3\�x��^����e�E?Z7�e?ʋ`0*;���u2��SO7K�G(�iq�=�b��v*T�g\�"�\1��f�e�곶�V�MZb�����P�`��m��}|�G驖�x}��Ҏ
�~��v@�H���0j"�7��m�,���Dp7J�/{��_V�YͻZqs�М�é׋?�P�;	��aU�Q�<	�N�Px�E�[�]���5�%�[@9|Wr�B�ď������f��F�%P�:�Bw;T2G'H	��TKM��:t��#���Wk2�p*�鷜�6jh73?��d/�Bk}�/X��l�d��Y��HA8�=�K�	��c�S���rFHC��[�Z��0Ԩ�A�&�:�+��cCi/�(���i�m���e���_WҢf�~�WeNt�҂J����f����z2<(|I������o�f��g+��B)���('�4�_ݎ�7��7�^	��%�қuS��m�|�������c��ɿ��Rҽ��U�M
�{�ʚ�ޚ��/O�u�;��x��ɘ;�?s/���a�M�z��vf�!~
�����X�M�$U���[��l���X�'������r���'�"�llC����P���R�S-p�v������OXT8b» I�"��q��3_s{ .����[e�<���>ZwN�����Y~U�cp�=��ᒹ_�fk�0� &{<���� ȍM٘\?½!�lcӁ�)�H��X� ?�
e�4Ҳvͥt$&N����,��U�	sĘ.�\��\=:�}y'fQ��<��rI�������/�i�KU�Wc<mvTz���01�f+er����D��a!�u�(;����U�5 y�� a��E���W���ѯF�X�H������7N�3�6.H��qL�A5�]n��l�촼*� ��\yg����أo��:Ra���4���2=��s�����\hP�ܢ�r�fk8%��Y,
3���I�q[Cq���*W�Dk�����yŻ�USs�?��Z���~~�Gm!I����^*Tg;����ci'{�z_č� O��q����-hY�	B�oǁ��Іh�Z��Pblh�1b�<�A��Ԙ(��cZ�jb�(�8P�û�x����G��v�D�<q����Hа��˃�@�7���+� 8u���_֬ٶӘ�a�������,yq�|`�^�ا�J�x�Ej^�x�����M��	U9U{[����W�{�Abdx!I��ga�eH��;נ�u�]�����Eì?4�a�yP6�P�H
-���qi1���3t��u���B�nw�Î-\���]���Đ{���bgs�������=́Zn)���Pw?���5삳j���x1F�MT�a����;l�dE�������O.�-x������B�T`\�  "t��r $1�"d�(v�,̩�&�@=D�7����
�[u�v
҆���/�$�1*��U��e��]��}X���ݽ��|�P��U�P�A�X��F�!@ʽ"��y�q�/y8a#�W7_~޾�A5L�S�/ƃ�>�R �U��N<�<w����?�[nS�*���UD��XJ �ح���h'I�68�8`H�LU���E�(�8�·+�Iơ�A��9� �����$!ON�
�O��'���Vt�G���� �拗��]�!�7��>����םW)�q,��q G�j����'M�F�l��#[�z)o�;٫�*�-����9��gT����K�aIB���V4ӭ����b�8tcM��Os����eB��w�������w����D�v�P*ڱ��~	75��iyt�n��eF3y�Ds���H������"'׳��"�[�T�+�+��.c�����ޮf� ��L�Ƒ\���<�+l�������`��Gؼ�Mz��q�x��p��T�TA�҂�R�\gMӚ�a���1�"2�4�>H�9rYiɋ&��wz�|���o��pT�W������<�kN����~����+o<��Uk�c�֭/-%lO�LG\����'�4Q�FV��2H�+:��z�l_Vt �A_E�M���G"����)B&�]�:�C΂��g*�,��ǲo�)4���^�*�s��W �:��4�K�T���i����A�:� 9yJ$�ܘ���1~{>KaO�'AhA�jW��O����;�۳�Z�$a�O>��6��b�.�l�_�~�	�b��o�_����e�DE���U�饔���`�+�U��n���-m�H���(敨��ս@��g���9\�tCHS\��>@�x\2�7$�� 2[�?>�B�1�J���|p<%;�ܓ1��vc�l-	5;N����h��$Ş^+)���%��� ��!�g���BD�e*?��n�qm2�[�;~1th��E�&��W�ծ�nI~�\>���7Z���m|40�a�����
'�����l��N�7M���ι3��ta��0F|>����ߢ���\���&���2�}�����~�-c6h�$˖!��h��>.cGھ�Li!�M�o栕
�	<<���<&�9���X��y;�v"�swE��tr,5��bU�z��j{İ��#���a-,�z/M}��f�4� 6���J�.=87��m�3ZQM�0w-�&j	2���%]ԁ�#�z��&�[�3g6Mᭊ��� ��1v�	c���΃WB��5TP���S��$� .�.�1���
8��z=?zzUg���Nv�4��o���Sj]�I�*'I��b��	��U�DG����X0�={�����=����,IS�ԃ��~����K��c�!�<Y��ե�v����B�����#X��4L���7���j�aw�Ag�P�V�$���VC��*JWٜT`��� �<%����b�%N�k�#9�3���PI�9P�<�7�ᩡz׶���#�K��]������b��/������r�)�X�~�n���U�+�'�/��2��Z��`jgqM�#hozӽX	E�~�F�4
��I��4�r��]��g&� 0�=󚂾'l'Ð=7h���6�K�>e�R��$�*��\\-fZ��B�3�zwp�C��^շ��B�r�~�P�/������	S\S�6�c��XZ7�6�FZ��;i_2F1��aGa��P7�i7�4�+�(K��a��b�]t=lc��S=���]3YaNd�»����^U>k���
<%����Ψ��� �\�F�܁�v��l��[7k"��=s?�	�O���&��$����FPXst��^S(Q�2��gz&�i�R"|���Y}����c���u��C{#�,�Rj�A�|�Sm(8�5�X�]k��\�>����6s�#���Vl@�x
9�t*��z�Q���ʆ���<C� 1�&���6�O,�'<��'��U�WE�o,����]�>0��� ֛[��/�6���hdL��KLE��V�\�����,�Yz���S ��\�.�U�C�W4�����{���ҕ4X��a9�4l27����o��1Y�	O���w��ח����oP�2 1/ ��G#�{�~�g0���V�7����G|Ed���3�"�6��ƚ�SL�Ti��J���)=J�B���eָ���
����|�.�Ss��$]R��苤g�0I2T�q�{�N��̭���c_ߩ�鞙���	��=��E�j��r��Mb}9Y�i`���R�^,�+ɍ#̊s{;C�_�u��hB��S�M.������y����@.����o���'G�"��?h�8��XD5���h0}R�cL��(h����P~o�;�^h�����v���sd#p���фwl�wL/��F܈���4�W�j���{��?it�V'���ƃ�����ȍ�ڐ����̠��֝� �oC�י��)}��ש?�uj�JT4�&��13!���D�������3V ��,ow�_��Ʉ�|{���������ǟ��U�5Mxa�s�W�1ߒ�=�Y�5�`����ڹ��v�n:c��� ��$��G!F���Iߋ��������{�2x�U��.H/�&_n���}��≴T����s���ic��ۤ2 [Ř�[-q����������j�s�}��Q�Qp⿢V_���'HP������y�Ў��Y���\�D�n��!���g*��A���V��5��fu�@�{15�e��%F�ܿ��^;������/�f�EZ[�%����!�P�No��b����.�� ��V<%D�cK#����������=i0�`���/����j
�X�س���!h�?9?�"�_��l��IOSѫ�f8�R�/!_��6C��!�`g`.0�Lb~�7��ӽ]�Hj@AJ�. ~h7ߖ�UIM
Ϣ�s�� ڭG������T�E�O9nB�F�S�����V7,I��-�]Zf5�?O��%ce����l:O��]^q�;o�ۍ`V��z�Z��:�ƕU:��h|;Ѩ�뭱[Y�X��zE��Ͽq^Q1� I�W�L� ɏ/�+�!���0.<�AA����<���:�p(BY���9T
������T����ӡ>��$�b_�~���qk^��G��!�C?9Xsy�ux=����4�~O�1誡$h��B�J��΂'�&�]���&i��c����g����>*)˩?��!�κ��IК+Hc�`~G�pp
	s�����fL;,�t�T�Q�U��;�������!� �N�#i	H��|���f��v�Rn�M�m����Lt��'�d��[y؝�f�Ceq������F����9%���56��&�A�jƊ��Ns
��&n6#�J���+��y+fK�����	4�_4���]�xb������z�����C� �.$���:X�,g���N�bb�� Hv�ʈ�Th�o����6������sӔ��N}-Ȍ䴚�G��?�}�m��+�����-ߦ�f�Lg����+��1��@R��1P�OKNxd@���q�h�7��ű��q�¯�T���+��*�Y�T�����=���$n\�GKTy+�K���wB���̐X�}H���^f�ϙ\��Ļ7T��E�|�ltw�
=�6�8h�� 2���#��u�ώ���7i���Q���V�ҭo�R�����LFR%����$�d�j��D�����16a�i�'��D��Q�&�١�9M̷��؏��[�L_���%�����f03��u����PEi=��`iZ����=Q]˳��\�<V[�	AH�Y<�����q�h@ٴD½�V:�1���O�F��`����j5��f(�ZM��i
;t���
E�y��?�����G��M����-�~�cE�����5�D��r���������mt����O�{��j���g��r��z��޹G�*K�;1,ׅM	xAj㨊�����"I�{H`�'�/-�� �_bD�Yh�'\� YR�k��-���7ِ]x�ʃ�p�t䕊PS�.hOn�&(*J���Y�ԁ/��"��asaQȏ�X���w����H�L�N���Nu������)�-��9���֋o&1jUhc1���%I��s)=s��@�����(3�m�S���l[��B��|�0U%��b�M���X�h��n��,ey~7u~���s3�r��~�|9: X)a��E�+rx u"gЅ�E6&)����O}=t��/�R��5$3���D���{^i��Ʌ�43O��F����r-��EqFk����.A2fY`rr/N{l��f��/!�V��/t[*듁9%m@��a�=������X$���9Y��'�ݎ��Z|���M	��q��pk��.k�y��uH�׭�j�	բ==����<��4�B��';7�������̇�ے�w�`��3gY�!8,7��Z,6��:L�n���<W�x����:���͹�J][�"�y�x�V}��}�������:��f��Yݯ��=ݿ~�����q��1��#�<�z�OVm%�%H:��5B����O�4��YZ���l�E�����	�\�C���P�������:k�LW�B|�����>�@��`L��'�D�S-���ې���4�ւ�~�JCQCv�qk�����S뺑�50	 }ʾ��G�|s�jMo�� ��if�B}�6�R�w9>	�i�+j��(��<1/w��N�f��a��CS�'ӡ�Σ�i��D1�m������v;��[u�}ɳV�^񚮗D�p��DJ�48W*�pd}� �����wF�h�_Z(Gq$����i"��i�)�>�;d!L@�"��m�x��j*1�l�?`�D`����a�-�lO���O�_�d�0G5����]����H���I!h54)��+�s=���`��O�~�0I�(��J�2�PE�!����k{�a'�Q�6z侹���B���9E<�n� :��݋J��D5ga�d��a��ˣ�	��\�B.���������ʬ��W���ȹ�v�����_�eT���V��|!����h�*�3��>6�t���÷:S��͊X)č�0�1�n���;>g���nsx`�|׫\x��wF��?'�Ҷ�T餼Bv�:�<�K���3��瓞	�=6�!�\	z��ӌ�D�{Mx��:aۭr��J�d[���h9`�ئDp�Q0	l�,d@�ԫF5⼅�~9�N�:�o]d�(�B�5��Zɖ����w*��*�9�qH��»�?�t�K�d����a8�q��cL�4�7�0ih�����e$W���]'E�` ;��1�Q�`:iti�,�Tdx^T��<>%Rj�G_�����DK��
rlگs���;��[c��[S���"�%�:!N����Y��tgEn�����%��T�������	u���<��Ćzr�7B�j��|j��#��{��Q;:���`�x�a��](�~���1�l���]�Y�_��@9�>w�,���|Lܿ�KM2F2����kՍ��w���ܸ(3ȕw/�x=&tP u躎�ŷ7·^�2pq+.#n!�X����v mm�U���B�=dl_�� 1s7$a�h��F(���A�l��0v���D,A�.��M���/!q������i�+�t��{�sphk ,�cy�6]��4ȇr��f�����yt�Iߪ���YC	��f��*0��H��{�e�}�e+%<��h/Ypn����1�Gtm'�]�n[S��s+0 jiL����f�Z��}�\[B�ߎ���!b���Zcu�oņJ��$/1��ٓğ���d�t��֏F���"����&,Bx�-�ǲSf_"�{�񠼤Zo�`�>���(�4WW<^Vl N.�&���ԅh����ݡ�#�
]�j���3�N���Iy��>	05V'����w�p�JS[���{�Syovy��fD��,�������P=���Ѝ&PN�f��G+�j�Q�һ���+��v�7�s������Y��(	�SL�H|C�b,TB+���L}\!j�@I:.y�5&�h/��"�%�Y�7j����f�����i>:����B
YG�cC�j���uV_Q�V����| w����'����6#oM6���]��F7�~��{���Zv9)&v:"�ד���[�1^��
.\̘\�N��/���ް�͝F�R��&����9b.e�G�Z`�	폪!��U�E(��*r�����O�����!�=�L�'��pWMb-12�w`"j����|���i0��p[f�0�~Ә�F�4�0��Oڽ���=�~{K��2��w[���t��L��O ��tſ;�����/����&�K�+{�eL*fR/Pdf� �l���J�e;�A��?9!{4�aH=0Hb;��� G�F�©g|�	E}������4p�q�����0�?���mͽs8n�C�	�/߂�~��ԩ���Ʒ�nԏ�3���^	�����0�y�۾��)�����.�)�1�,�&�O48C���t��u�+pS��zL)��A��iVW�����X2����V�B)�9䗾�.Ê��݋���b��ܮ5��8�'��t�ܰ2�7}�J|vy����6��
G���Bv�q�3�ݨ�#P�xYy�k�)�?D5t�TX\e���o%[��P�1��=9퍈K��mB��i��#I秗�Js�70P�e�f��5%y�S�I�1�t�D�D.�zS�^�LA�����>dYY� f�*\y�!�����rf+1�\�}*ڮB!����B�>��E�����X�0^V�ɦ$�c�i�.�.�KЌ���p%���eq�:���\ƣ=����>��=���[��M�SŢ')�����ZfQ���Q?��ŏͶ9�3`��y"���K�!��h������1.1�ژ��6S+d�����Qڳ����޿u�m>N+��ͪ�fn	y
9xJr����#�4�I�MQHk�5,�~�/a#5�j�<=�B�a��r` �����8�%k�֦@�Nџ�O�d�����'���x����:Cэ���B�5>j�M �r�%�O�9��8��>mJj~�g*��rTw�^D1:qV��lX��B@Ey�?�B	@��z!�0-������	:ȎFכ�Dr�?O�w[�@��9�V��È#�=���G�m[l�b����v@IN�Ba��a���|�t��v�	�H��.�C��|�.'��5,�b��Ig3�u^=$���=���3j�`EDYUS���L,խFa4X��t�N_�|9�x��}�U��[Q�d�kjgH��Z��.~&8�t| ;��?bH�|���Fӄ��Ӻ�3�\x4�{��TZ��1w�i͉��\����d���ǁ��_pq�������b^d�Б�U�F�ي^�/��b�7,�x_: �� 
���S(O����ɂ<�`k�`e���Ez�T%X�����N89h��WӨcs8]u0'X]q��7�"�v������)�8��4u1��=� ���n_*��>;�L)�(�ծ�	��	��'' )��z��LޯW����.O�_����P4��m�.�B��p���$���
e�>j��$g�P!@�ô�xuwY�����j�3�f'N���E������3�a�!8�&�=�>�(�]*�ZЛ���n>٠8���4�YGs9{���|},��ʨ�=ُ<�27�A{I�N8�v��ZlV�ۂ.�~i�\�j���KoyF3����tג��_��<+��auu�Y@�j&��R�ȍ�}�@z3w��T��멌���\7�Zk6��hY>���4�kM�p�y�0	���[���Q�}n�=[��a�1�̿��������>�'҅Q�9���$�09ɓ+��jF�;���4�%7 ��[H<���-����ٿ`�
\���U0%�W��	��&��e�Ɩ��Ș6Na�{�bv�0�|�;�E�b�ߜ�C�3��t�޸�/�0�e)���(��Q*U_=�K7��U�+���e�P���x���;�b���?
#�S�r����P������T�Q"�y�%�1�`<��i�u���~v�[T6Ѧc��E��g�Ge�ȹg׌�̯B�� ��Q�¤���u�{���<�!��2������������͘9T~�l���:��>�O��zXz�K�L�c�#٥zꘒr�gwVV6��R��O��}��Si���>��R;���8�_������;{i��9�9������oX��T�&�z�
���{3*|xۋ#�z?����ǁF��j��:w_�-�2�Z�GHCl�*.䶐��Iխ�o��Pl�T<�ہb�jpt�_��DԘ�_xf��7:���G�@�H���ҫ�Ѥ��h-[z+���u�(ϙ<��ޠ�ZZ���cG-AI>��*���H�By��dqm_��|�t[3����,���E�-�I�m��vipn�c�F��������}�܁'�nT��g�o�W�$�j&�0��ӟ��  �(F�-��/��O�wr�lW&�)"��x�V\QM��e���&�o����Ql��������T;|���s�O���F����k��*Iͪ�q�a~��ty�������Zj����[�������3�/=�fjRlK0V��9�9qG���zGa��` ����d.΋Eth¾�@<��[����ė���'n�X�K�� ?���|���RU����}F�nO@�Of�W��j�gD�]?�eM�2\2����l|�)
���G��R�S�n�ԗ�ċ5�� ����l�+��k�����ׯ�x���=��O�U��U��J�5����Z�4��ND���3��o�$-�	m��A��Z��^� r"4��?.[�[�c�g�|��>��{�4�3{�y��� �@0�{ ^8���!�����G(u���8�9��1Oտ�h�>h⏒^��2�b5�+�R]!�*����	��$l&�з "y�%���+����qWU(k�\軘�.�v�-4W
���$��R�	�M�'h���C!l�(�X��xF��ǺB�
�8K�g2�W����pp%��m^M�����L؝�1`Br����[�V �P�yS��
(��2�Yr��p>(2%E�������}���@i�z=��\>��*��R׾4a�J���D-Ѫ�>��95�pH`��1��tbA,2�H[y�Ű��|}j]�&Z�����,$s7ߊ���?�MQ7u���uz�3��$RŨ�'V�!Z�V������@���9z�Y�	��Id�i0�6M�`/��!��T>h�0�g��r/%u�{2�^3�O�S��S������(�G_��ek:~�9�"J�ŏ�2��Ռ*ӕ;~��lA�����ȟ�.�<�3k-G����H������:����PJ���Vn���r/3�'�q�S6��N/�j�B�*���p�����n}^�M� v_()-�.d"��!���ώ�mI;�W�3|�(�#~v3>�O�sY�dۜZR� )��Lv˰��s�ʉ��*�VrH��hB�֬��[�7�嶁^}� �?�����Gok5���ט�F����L� @�Q=wݛ���%��>pa���Q����ZV�{9�M�Ѽ�W��xg���x�綱s�;�
ǰ&/��{��ʎ�Ak��聑�D� ��9���ĄO��N�q��U^�<�v?�^w���`��U�*��}O
7 ��R�����PV錒>�
G������8Em��ńĿ.���^$�f\gHN�=wGaa�Z��hB�k�⒇&��a���q�V�J�ϸ\u��E������#2۫H���'��ԕ�N�����P����"�55y?�^����<#c�5+o��L��Q`,�KKP���c@J��k���܁876�E����̾�޹�ۜ���\���3>%0bB�tN�Ph(����@;�Q�v�N]�ri�kX����<��;�U>�^VϹy]_$������\g��U��l��
wP�-��.�%�8�WXv�w% ��!�A£���m���PᖃZ�i3/����ƿ����Y�ӬX����n�N�DMn��������%���Ur��ٞ�76�47�[	��U�	D�1�ɳ/չ<��(��\��%8�.���3h����2���6�
����y��k)��[@�) �]N�d�w�Ǐ��@�Eb�%"���Zk��g:M?=�#�c��%��|,{lw��Cz�*���oe��y;3��/g�\�r����iK5|>?�2�C.誻M|��yv���-`�jM���hCdx�������� n�����&��GuY���������[���G��������	�E;!�m�8bG�1_8�q�/��L���K ʜ���.")Ŋro�����������VJ�hz����AT�\=�Sy��5I���IH��7Nl���/k��]��*C'�+(%�Ϝ@����/5kI� #� �o�Q�}��3�@1�������J��
nS�}��g�q2�/ �ۗ�g��A���-��X8e3��q�I����m��i��`�,-|{	��K�KkL���R�x
TO�Z�	ڵ
H.�u)h�2e8J�Y�8$�"	L?�x����L"ʜ'� n����[rv�Π
��� �J���ھ8i�=A���@����1�`zT����	B�	��b��i?mZ�iO�Da]��Kw�����oqζr/x�#
�	�{��n}H+\�a6zN�*�B����(�F� �:��p�����6��4�J*��&0�Y����_�!u��$���z	x*���� a`9��c|f��T�*-G<�Mx�d��Vՠ��G��!�ӯs�%����v����o�3�Y�3u�����/�j�� ka��!3����?:�����k����3T~m��_�4�Ϛg��2T�[���,Eb��]PM��Xc�-�{��5�@7�?h�5m�DT��r�&(ɮ�s�tuK�T�S*b�7�%��T(�ؒ�چ�m�1��H�H���v�zA�S4�v��"qߗ���W�uM˯ s����t��cA���	�� 0ʝH�?G�ڍ�Ki8�@�cC���zw�|� }������X��&>a�μc��WGhq]dS���),�?G�!(/7f�䯀��Z�fE������X�@Ղ�5Ʊ}�/@��Q���w��X�yD(��L���׳�Oes�C��`�k�� T�~_Ћت9��\�E��cM~���X�&��.��0mmp�òy��j���$c!�9J��Y��>�`�'Yb�pu_=7�:���fAT,$M�6�p��6%���N�p�ԭ����-��}�Jyȅ"�'���}�1E�uE�6�J�����;����W���J��~�}P�jr�L_�"`��>W@3��o%��Y�'@�,��\��rʂ��J�qX��n���F��p^�<��x<(p�[Ug��g������x0ЀV4��ڐR�����`�ٶr���?f!=� tuԒ�RY����z��4�Hj����c�3�c���eC�B��T�SƢ`�:{� �f�" ���2���C��-�˦�w/ʪ���q�$���9P�d hb���-2b���#�m〔���  摟�c j�Z��Σ��jG>���&�e���.�#�pdǍ�!뗵��A�4ˇt���7��e�Yϭ�&v��vΙ�s��vĨ�p>�j�&��a��A\�:ERc ��k�	uX�рܞ�8��r��L��wW�����T�6K�v,�|}+;f&b��H�5U|�4$ g��}���5�����y�-��b��1�2�Ai&W���r�'C��G�ԉ�A	M���?��M�]�k��~���"��2j˪�w^���ct��X��~UrN5 �nW�脞6t˔ �垒&Fj5/���s1걍A�I�k�n�{֘��,���� ��獺m�svǭI���3Av~��1��ʛ�|�.zYF��;`oI^�ȭ<�k�I��)B��ٖ���KK@J�s��N��*��8�0�_�`�}�c�u[������N��ٰ���9lc�<��)q�J���꺧d�����A�'1+�����#�SݤX����k'1W� ?��5Z��վ	�M���I��u���M�u�h�W:���L��%�h��`c+�_��MO1'3���3
֘ϴ�N���r$?1���;�9���?gh��8JK]�A�:˓�
\T
�Y�Π>��ǜ����ŋ+�����4�rj>�*�~�?UB_�U[��7�ְ�@�Do)���������51�%��g �-��.6`)m!#�ÔĈ��屦6��2��$���`�G���n��f���F��%�
k܀�Ӝ���d��$峗���9�ـ/#�݆���vB�� �**�~��Oo�oμ/��=��\��J��EM�p�SJ�`*��1�њٰRWGX*N�0�^��B�c�u>f"��{�F.��J�Qt~7?���`bi�#(�X+����׏M�Ibf������0�}���AEDW;Ҵ6���Ĭ��W�ʑ06�{��Ņ$ɻ^�A���*V�� :Zc�����`/Fp5��~?�-$�ik}q��� �����B��6�� ���Ou��븫D)!��pS<TAΦ�?ātމq�ӗ5ac��|Fme��7�ڸ2�^AV`�~%�R:t4_k+�Tԗ�#!M��qE� �W�����I��	�_2���1�����s���!k�]i0��2���5�T09�b�f!���؇_�&7���~Ƥ��4�kh�+������bl�Ҡ��'�- 
-��ѕg�<o1@ �\W>�dԛְI�#K�:�%tG�9g�h��
��[�YW�� �-rF���(x6�5�nݝ�� $��+_�
��=*3-��!�i�b30�^$AP��W�	��ԑ��ue
�";- ����ۻ�{�w^�[(ԈH��D5�v&+r[!��IK�(q��i|h�'F1_1��b��X*Xek��g�#��(�2[�����x�2���S[}R&貉AC_tL�زU��e#%P'1�r<`���8�P�]E�3t�Em?:�~wæ ��.�ܚ�_����ۑ��3�)�9�ӇM{����f����q�O������Y˗B����Gۋ��[���Q�|<&=����9�}kܮN�@J��>l��u}!{���>�"��_6&K�0>�9U�
Ʉ�� '��D�pN!e����w�����1hu�W奾\V����U�^�� �&h���`і��S��ߙ����O�����;5���Nd��T�5�g�q�R��B�4���Q;�H�F�i�N��O"��k�,���Ǿ"�eF<��HF�!�Ͷ�{��7vk�nJ>��LD�y�ף��^yI�5\[:h�e�&�A߉t���� ���>ti��^�;6n.�5ˌ=�p*W_�]��Col��SE9��Bp�l��Jc�8	�����)�FfP�Od9q����?��:�����8�����.z���m[������N��1���M�U�[	}O@oo�c��'IFg���T&k�#��>Dh����[�`�8�X?�
�-@@h��򃂰Fk��w�,"��≊;iTgLPL�g��ɍ��H���T���ID_�2�V��M��q@���c��<��ׇ	�iD'���f�r�vAI4A��3��Z�"�d��Z_���ͧ��*�So+��le�NI�|!�L�k��NO�f�q�Ǝ�t��qd��E�7A�:��)��D��u���������Q���y6�u)�ۙg�ioU��V#k8�j��^���J��`XwR�A�]t�e�H�Qppt�{�>f
�������^����6y�RO��Dy4%��qv-_h�o">�xf�e/�>�~��̍�qiTEs�c-=Zm�m(��F|� ��?�;=�?�V�#����ˬ���9�_̋�	�� �|K��r�|G�K`���?�����\��r��k{O��I�4� �y(hY���_՛Lv �Ql�b!��]��!�B�9?��S��?�~�\ ������+oW��h�r�A8Հ<F}َSK)��C��Mww5��Fв�]LbZl��G�;(��`v;�+F��.:=�%
K�%��5���^D��2�I#`�GS���x�#sgX�p3�#C޹�Dr�����/V���T��,�sr�栄��A\n7��&��l���� ��HF�QA��H�NV��_�����|�=t-$�����{�윁	����!�Eh��X�A�<Ǒi�ˡ�������	$�r>��L��(,b��7�Hum� f�к�[d�B'+j�$��Ʀ"ߗ�B9��D ���l��]�D���V�>��`F1C�}Y�o�bx���-���!ؔ�����ZԕcS�R�����J��qx�'ӔHѐ&{�c�K�:*Qo��6݌���j�]Lū�c����䨻W7��x3yb4qt�g7[N�g���5e���"�*�΢%9O��M��?z�/zz�@�KyzV�O���^{ݪ/F��	JK	�%"��K�$Z��{��(u��v���,<5�.�"��A��.z*�Rh�04�DeO8��h5H�f,��)�=�[�-W��r�F��:�׀��.rӸ9H��E�r{��w�!�`{5Ou����u-��)-�����i��(�q�c�!�6b�y�% ���] U?�����0��P�{e �8b57[�0��,Z�v�=ӨKu�d�v��A�ϝ�8�Ԇ{}L��A�*f�2�]��d���b6�C�N����/��]��:�	z+RELȯM�Wt���Tc�e74��- w+�i��q _`�6y��1l����f�N�?���y�'���@��X�r��$N��z��O���#�-N�S�v�n�wqt�g�z�&#3���К���I5řs^x<Ci�E7 ρH{��@(
@P�tv�0�&�Z~d'	�yK�b��(�4���W
jv�B&9�8R���~Z*`�LjmAh�Q,e[��Q's�����^�J1�&/��kf�?��������Q��\�U$+�#�w�Q�}k�S��:h�wpIJ���5_<�[�_�/�Fvl�9a�xX�oaT���8l�xͭ�rv��z��u.�pf�W�Z�5�❄6`���|n��@Y~5�>y�{��m�qϲU
� ��AO��Z�Y��Z��c��kG��Fy�^ȫ�؛4�v�6���!��:�I'=+ݬ	�=߆E�4
�lE'����W���=�i
~<A�S�� Qv9𺛣��[��G�����~?�D����Ż��ݳ���}x� AC�1:��nQZ�jB���`����@x��& }~�ҭ�:-ƭ:�a����}׽���/���2Tw����`W�Uv Š!��	X�b�:2fñf�էzw��xhjd�����3��|aUE��el��T�v���pmyB+M�����w��r��O��.��k�ǰv�D�� �<S�iԼ+���{#��C8|���j��ӧV�x��[���m�yƁ�.��L~�m�r���+y�5p
���r�w�Ԕ���e"� U� �l��]4�e��'�O}rt�g�Z��-k�M���l�z��2�b����$�>�Ɂ���� ��@�X�����n�S��Á伡k�O(�}c��_�z�VkGGεs�Ezkj�1�疦��]p����c͡�S{:Y|S�FX0���K;c��-��s��`�����T&<���#�	.�yz���.��a��^lBK.�k���;	)VTv�T�˄�kL�M�
��{倡����������%��j'�z(LMF�Q�jy{&���a:7鶇�7N�r�X5;���@6�I"�]���ƃ�dU�yqU�,�R	yR��=MO2�B�-�`����L�I�SɏQ(#��>k�w	`a��M0k��i�V4W�'�-��}��H��xI���	��y�4��aL��}�+E1�	Z��}bc�^~��|/�7�o�=� k�xF/iy�p�0{di���I[2��~|��,�)�fl���on�����4,�P�F_d虽�+,
�G5�S��������`��s�BK��fi9u��̌�[Z>,�*�㎌q�
4{���5'4���iw?H�(�xLc�z���x��Ո�)�v�������f���ı�Y�6��=�cwk
v[�����1C���ӻV��¹�S���E��9��C���vͨ���Z�χ��ҏ���S�F�+;?`e��8����}��[�m/"j��E�k~-��*����E;)����M�[k◶����� lY���t��Z �:6�L:�6���*���+�T���
�G=�.o^d�YVV��Qb���(�}o�/���a���) ����6�F'�23��!�~_����T��آd�ߚ���Л�`T�v/s�ܗ��ǯ!wՎpD)%�մ�UY�tV�<�X����X��^ã�@d��1YJ�;YIɼ*Y-&O�� �ňW��D�I�l���xF��o�sSg��Ev�e���x�,b�<)����E<�dO������o�=V��^LV���.76�ؔ"��A�$O�ƈ��]?gn�Y��Q'����jt`��ԘZ=�%�V� ј	�����(䱂��+�j��&��b���6�����W��g>jRl�7"����A�8�Q]���gX��k��o�xqTq�)�u(��)uB���`G���Ő+����20�)}���e���ƒ��m�ps-�J
�6�/����Bw���5��HGĔ�mʶx�<D�R(�0�L�a2�k�
���4ѩ��)��r�f�;W�B@tg�E<�6dm���4CRu���) ۚ�SN*xB�@�!Eվ�fw�� �o�6�ԥ�ǟ�?�#m�~I<{P'�-?L6��.YLi:?�Te��>W�9N Z�b�_�^�~Y�N��W����x��/$�P_�X��H$�J��&��Uޞ����ze&���hl&W؝�O@�nQ�ON��iU$C��!@0�gN!��d�-J�����$�v���2�
p�8��g�G��]V�wӹ?F�r�-k>�ﲯ|T�g�rǣp��D��ee1�HJ��R�lR���`���=Ë}�� �9v+9��lB��qi�k�����L����-��A���U8��܈������A�
�wvX�n�cP[��l���z�=���KS�����C��t�l\���6g %_�U+�{�^r0N��b�������R�p���=��7oER��.��+�{��+�rؓ�����^����+���L���;�[0�m�^&J��/¦$�(����6&`���Z�ڻ|�#�Y�&~[��xhݘ�Z޶��Z��d�s�����W���꟧�������P�9��2��sR3�<�ޮ��ێ?NBj�xq��96�_ ��X{�-Y����Go�N)#*����P���%��]c�m�%�D�3�Yh1�[ė�L�5O�s&��7��!oK^��l\g%Z̭���g�c�'�)�^��X۪���P^�����@���U���K&���Z�W�n���B[M��6��QQ�Ѿ+u�� ;Y`�.��A5V��ࢇ}��_�[n�<:O�)�2��a��h@�[����3�����R��G��;//�pq�4���mH,��*�qn�XP_������|��*r��k�(x�~�3�����e݌e�sXC�]+��>2��l�j��O�u>�T&z�W��]���lz!Yl�C-����r�i��j�7�)�&)8T��#�s�i�>�ň��m\Iv�� �j9��rp����ld�(4f㾒m�Tx�uW-��}��jA(��/q���[�;�Z��Y�����I:�����
�ohX��[+���0NPX�P�u�7)�cj:h	��t��Ddk�z$`�?�鄡&�m�`�._�ڒ�p�6��螬雡k�A���k�+8�E�;�.E���\̍IL�C���;Ź�VNo �ׯq�w�1��5s�4uK�;7�nz%ޭ�و��b'u�
�ckr��QQS�!�K&��.;.�g]܎u1ĸ���"�\U���Q�=��8E�
 �qaа0jU���ބ�`�p�UH> �$�_M|=&^?&�C�p����9E��q�d�؈%� B�4��������Y� 9���jk���-Ӆ.$ς7		ד���u1!t�%�C���]n-zK 1Ƞ` os8��D9
ҽ��uJp�X^�.1��}���f郙��F��N~{�)S�٭��qC�\9���hZ�~�I]�)�&T�R+�s�O�v�Ӷ	�J���o\��:��(���Ps��#z�濇��
_l͘z�y4�J�Sd��[���6���|#��4�~�T���K��*�`��������Q��v0\ȩ��']�]O�(������g?Ü��k�8������/r~�b���A/��i��������gX&D�,�����#Ey�,���W���NhAYui���Q��Ԑ�K1p�&��(��G�k"�t?�挘b���R*�t�6U��A��1�_��ډ�xD9���!��o��?�=��:�9z��M�Z�k<0�zoZ�O��A���Y���ۜ�#�� �k&���1ޢҊ ��?i'�����V�6&X@a�7>���Q+�2.��5_�ff[���MU)��X ���+h�&���5�z!:������3��y�t�I3����s�]\�a>
��Rx��1�	P��x S���p�cE!��1b֥#]�Դbl�_��6x�x�^���;�(�� ]n2A�<�_�X�s�K	�΅a�B����~J_�Y����"Q��r�1=٤����G����y�6�0k���֌}�݌b\V��I9)�]GL4��>�2���,/���,�A�XT)͝��Y��L +ݛ����Sl�?Z������6U_w�O�D"θYc?4�����q�B3��r��Bc��/..S�_l�L�Joߏ��F�}j��T��]6i�")�ؖ�b���Uf( �",C�Q;�y(���|?H� ���C��A;F��(���'�*L#�����K O`vg=�P�uĖ�X����X�"̘#]��P�@��V�d�!/`��T����f����_ܚ����r}/M��<� � �#v���D��߭�%RP�P6t&�T ������ �5H�5bR�m�>s���6RCY+�
������	��F���%45g�z�6'���̾q&����=�\`�[�H#v�`i�����S��\MYYq�gצ�G6*h2�%��l�����jz{=��,��_����kG��4�����	OR�&�ԉe·�<���f�L�ߗZƤ�܀�\�-^�FΦ	�e��X)V+WT�Иv�^��$c����r57Xm�.��*6��ο�V�j������	��c��lk�@z�xϑUYgLAc�Lr�S<�FaKP�����������U�0�x�i�I�����lB�tsh� u��x�O�Q�Eg���3)j��=���qPT�Y��d݇����^���!or�I���� �*��!|*"�Fi�p����=;1a�ߑ
�c���9	�\��x1���rK�W�8��{V���mh��;7l?k����H	M���W��	&O�#�L��9�,�2���c���$�ЌC���',��6�*Ϭ2&��\o�n�(�h���EQL�D����#1Z(;�B�kpʙL�|�����;E�&�h�%�P�u���J)���a6��й<t���8L:Y�e;	ͯ���Ez[�c���:�=���Zb/Y~v�d+e0:{a/�D�sOE���L�1i��+�rz	���J���l��s��8�#�� P���c����f�t
������~H(�6��ǰ{�S2���ҡ��s`kMS{�����cSc��k�M-4'����έ���w�ۂ���8�R�$�����cͱ;���[�?�(ͦ�Z�����G��7�<63�@�0��钡s�E࿛4��G>KG�Z�Q-%��¾�m�M�@#s"�˘��.��k�  n�u���1��V�梒�Gf���5^�1cCDʻ/�0�E�W���(�
s.@FH��j��m��b�-S�|6o$m�O�0�;�T�&��ƽے�� v����G|H��{ۯ��ǳ"�6Tc]����!�:����5��)*
z �O�P���!*�*�M�t17OR�VC��S�`[�d,7,�(�3@�x���n��m9T�Ph�^��'�<�Y�� ��hޣAXXo�m<2?����8�8n��휨�ѱ0잹�o���M�r�J���TT�5'�EP�����5�'U�,�Bb3W������(��-��-�<��a�	=�q�x� ��R�`�4� �<_�9-�|%=T����z�z��s`��x����� �׊7e�@Ot�k��KQG{Wb�q��o��!G� $�n;Ֆ�F�gb���Y�>9�������	��k0'���?�S��rg�[�-�ϯŤi%)Hg�^��]ʣ���p�;�v�b���`o����te��
��4�YݩrsY��x����|Y-���Q�N	��Ұ8+^���De�
���¾E��� ���`SnÅhfO��|"h�&��UI�y���-(�Q[�*r���n{z�l���zh�S:�B�V���Sg��!�;��Fr��!w�ώ1�}���v�VLe<�i�2N��#�y��领�-�O�oE�VG8�D$��T���w��O�����0PC7'q&�Ͷ>�q�N̷V�������Ι!�}u-���9��Ƒ�M�ĸ8�_���9!ݟ���ǣ8� F��t���?��4<��~�� �5�!�%��/d��~��·���to
��jb '\G��t8�j�w��J�*����#�|M,N�z��0��ņ����^I���t4Ee�D�;q��L=�L���I��A�Bƥ�?��;��z#��M��z�I�[���D_&9\7�p���B��fFt���c�(���������"�&�������[���H��s���.~�x�S����Ѣ⛲	B���=H�Z�i�򾸌k�NQ���+1-C4y�����چ(�FB]4��0��0.АA�6��ʻ�&���rٚ�?]�'����Tz(����{�'%��;�ȼ��xy������5���f/n$���F:F}N����������\��j�<����]8��a��S�r-��J	�&�{^+�I��������,jOԥ�/@�M��xdu{���I��)�o}��Ǹ�!(��Ń�i�1y$i_��B�æ�8����ë�+&2��;6���?g�j'��w�i�V���ƞ:�7^c�����G�_ةG���+��U�<\!�؇Vj�L,�/�_��<d���۬�,�������Qr6s��P��I�� .BJ-��A�YJ�_���ZO���ʏ���&'��C�������/���Xʠ~����,m#c�f�!P�w+�\#�f ��c����|}����0y�.��G�7�FhOv�C �L&�!����R�m �w ���p	��6BB�+�O�q_f�-tP}+��7U��~�N�G�i?�G�@B�O��ۻv�>����ꢺr�m�H��ȃ�T0>n�H3�W'9���W�3@m�7ćXqk�5�W���i����Zs�����*jv�m">f���XY'�DZ���]��Kp�����2���i3��CPɀ�j'G�9Z���2�	��zo�%^��ـ�Y}9^��S���O�5I�<��l�D� ;a�tb�5�;����,�T���g�	;�F�s��u#�i�/�����&n:�O�r��:})8\���Q�S��C�$0؂���g)��PL��j'g˸gԂ$)��&��R@��:J�U-�Z<��X��VhLgx�GJ�K�p��Lf;B���\8��3xK(��nR:�6%����vn<
�1�������L*�j�r9b=���ַcS��^8�k�@��7�a{����K��N��x%��{c��F�+��xu���_�$~� ��w��@ ��O(tOdͺ��Z�d�f̲�ťt��]���;�%TJ;���Cǖ#�ީF��}?�5�[��S��oN��!��P1�A?�2W�V���^��D!��in�������%`@v?HK�X�B=e9���6nD<�p�D��Ì��yP�a�P����Ĝ���\AU�o�?߅���*����+/�J������*�DK��8�$�ɠ�^o�ULg�f���w+8�T^�N���#�}�>E��~C�}Dۺ}�t���~ۨ�P{v�)R|' "�2+��=�?�\����D5n,?�p����O%�U�)_���z�{�0��a���$�cp�-�,Iڷ1rh�M�~��U��(�y�@������n���8k�R�S���!�B�_""{���	��tg������8K�%�Òf27�0G����A���+�:�W!!gn��Ү��q�AW�[^����!V] �t�2W�׫/��N����ح�7�G�� �˗Jʮ�1.��g���\�/��.�
R�z"؏D��r&
�l�@id���vN!~�8��TZ�v��?�IDV����"�PNBVs7 aAZ��+G(������ g| {��~�n\&2���oN���RF��pW� 3f��$�u+�P���рMv� ���QO]�{W'��I��,@V���r��������(�8�0S!���-RJ��6���C��w��rNn����*?��(!GP��b��P�Q�����?�G8w��..y�l@ 1ߦF�0��x�i6��.N�����Z��{	�y ����I��3��fj�6���!u����}��厌*�0���o�g{�e�7��D ���U�4��bD�Vm�2��ä�2���I�-"3ɕ��Wi�e�+���nͫp�30Hߘ��s7+P�{��S������ w:��/\���(���k�1!���	���t2����N ��I�"�T�6M��r�� ������1�ׂ~s�2ZZ�������	+�G_��i���<'��ZEᩭ!�hT�0�q��E[1�~&��\9�>����uŵ�ᝦ� ��
U�~�\J�d���8�X��m�ւ|���k�_�b����x=�3z�Ȧx[�B�R���2?bu�=Iu��Q��<�vs����Z�n�Ծ=�}����it8�P7�f�>�(ʞ>Х��i�u�;Yit}8rQ��{�Pp�e�Fs�.*�u��qD+�����Lt��UV�iJ�3�Y�w:���5&L.�R(�JL��ܚ�����%L{��\�����Nl���pJ��½����l��~�gKQ�&����())��Ij~f�q����H�����?о������|��2$�C�T����yP����e��N�z���}��J�Dh��dl��\�E˛��&�2xM�I~{�4x���ǽ�& ���f�.��Iߧ.��4@��E�O"�n�������>�໒�B=��Gƪ��z/���	�L�]���[������MR�u���Nn��ֶ[u�|;Ox���f��gC%Q<*M�X�
SJ��xS��=NrB����k�/��w?D�.�Gc�]iV�!:��c;TTA�� <�D)+�g?��(B>E�@��OS���"
�B��~gͧ$.�A��C��)��g7e�S�
�ْ�l��� 3�w9�����A"��N&�tFʤ+8�vW��}X�)]�����+W�����ʽZ3����K�xa��{a����a�d�t�mA��Ѝ����#2F?���/iH�w)�0����B~��$��s��i�w��z�	7�d��iC;�~�� �X�������XToH!ª,�P��r�s������j�Y�Ƴ�c]i���t,�J̳@G�>���@6:m����0@C��(��ߏ��,�v�� ��ϒ;i-*�����eǫ�:$��4~Fc�˜y�{)d�I�̦,�LT���($^�M�.�m��΍Uj!F\b�D͑oY���p�=�yS&�
c���P����q����T!����R~m��t�!�U��xU�u�j��ll6[��P�A٘&�<�IA��	]�K�M�g��q ���	�B�����F*4Z�͇o�'��<�̕��J�|�@*t���֊��s���g�0�����@assiC�Et�Z��A
Z"�(ŧڦctYj��[��$�l�|t��2�`�ǧ�s�r<P�%�9-�@���o2�����<C&��I\��Q�+\U)��w�Lruj����KC���cG$���$�Os�ԡ/~f׉�@�g�,��CȀ������NM�s��jk_�f�K�9Xe(\�5j��1eCǜ�-�Y��:~�{�ażE}7�S:��P�:�z����xz�������,;��޳��AX��H�%�X1�[ij�%�I�Z��8��\��'N��`�:: � }h50�ꛠ�E���ӓ��Q��Ě5̰j��R��^���Y�\ݴ�vE��=-*� �Ω-�=���'���^�5 0�u�&�Bx��nȔܧc��tl!9�s%T���Èɿ'�v����0A&���[�_���#��+#���A��t�ή:՚�a��a��28M�h��dG^h��[�|�ϳ�]�p_�?��J���0~
�������J���<�b�����Ʒ)�>��(��	=�a,e0E��`����ܮEK�(}쉛��b�M���M�uam�ws^LY�W+9D���6��\�P���c���\�ּd������ɵo�gp*��zL���ײ[�="�-eo��n
�ВoV>�5	rb�$�a��d�R��绤���K�1�]K�K����֎��G�Dp{3 a��"�@��M�|��Т!g�Q�3���&������5��ӝ�(�-�L�} b��d.�G�Gj|�c�����G��9�����-b�I�N����T�y�|��x���1ih-��WZ��rյ��Ѻ@N����Oc
��Ĕ���tgQf�Qқ����/v��
h�WTt�7��>LF�f����0T��r�i�q����@�v� m笖B�P^�AOBP\Ze��V�f�S�=��g�S���$B
�{Ǻ����W�*�l�Ee�Ʀ�[��?�Ќ�p���u�90�h� �1y����@Ϊ%*ϩ�+eR�r�cP~�-���7�U���:) ��td��j���j��Ơo(���C�C�z�M!CRP�bOZs�՝#y]���6�>UN�����>�-�Q����^\iv�RfbJ_�
��M��}�҄���H|*)���C�#���`�b<]
-�`:Ɠ�8�J��6�����uG��Pg�Y�zf�,��Q��\���1^��}��15�,��ƶ�?�(�<5�����G����e�1ypk»�W2��tu!�����Kh�����eV)�Ȇ7琾hǬ���nA��
�����z���s�M��qz�.���,#�8���(�Zs�93�2D��
�I��ÿUxxL�H�S}��=�����ɕ�&�~��PKH�tI�7�g��O6.8�+�3Gb9zjzڦ��y�F�X�'^�m�ê��G�����"�W8��|
JZ��Z������U�d���u�<B@����e6Ik:��qJ���S_�ϓOn�o`LQ�	1qˤ�ހ���U0�u�DYv�y��Zs��Z�11����諳�Sti����Yn8������Z�3���MY��՛9�k��j�=!��dC'E<A�3�({M�>��@Dvl�u�w;�;R�v�/]"~���>��P��.��I��9�&�8$e��Ea��J�m8���f�+%9��pɔ��_J�ph�\DJRKіQ"=�52��W�O�����΢N���(�@�����;n:H��:�%˯�3��f���M�9(�;��t���7IP�*N�Y{�l����*��I͐��<���h�l�k�&4Gr�̂7��Ԩ�|�����!$�O!۲h��-J��6�_J����1"�(���tt���������a�r�gYǫ�\��+�P+|���u1�ȔX����5[���I�8���@�"B���o.Y����j����Xء��N��b%T�7׎y�W�E6O�P����#^gVY��"�����v�l��$H�M�l��W��V/���LRD��? ��{8����c��U��L�&�a�?�������Fƌ�5&�ڙ����n��w�Β��\�Ùo��*q����<��DO��IJC����bDK�u��T��2�BT��֦{��а����]"�+if0|�K�j�	q�!���~�O��YO���I�YAYk�\��3�� ��BO��.�c��^Cw�tBN{m�'���E�$�q�:X5�3m�p$��<�r�������{���b썫"Ʌ��Y.���$�f�����$�M(�1n]UcTL�t�������p�?�ƣw�Wׯ��9�'p�=��.m�V��}��f`C�RC�ޓ�rdٛx@|e�ɹ�5�n��׫c��~�!,.�4��}��	��L	�%���F�,�p+8"ʁFR�l����詾�{���-TwPU� �.��O�zˈ�B<�� �鲉 |P����������$m�~��l�5 ��@g�"��GZM/��bGlg#qW�3'�x�`\0Ҡ��Ԇ�)_;�d���"�iiޑ�=�����&1�Ѵ�����3J�#v�o0�3�����^9Nvdy�f����\]�L{|?���T�1΀��OLv�� r4:!ˌ�h��($�l.�%�m)���(;�,a�s�G�g�K���{�!?����ꭩc����7�����23�'�2��f՝���)��F��p�"6�#�gf"(@P� E��Ic$"�ڄ-D���p'�]A�s7���� �=<�K���q]C���Ē���_Ȼ���xo�ĳn}CZ\�&�4�~rmf&jg�M��1�Ke�h�Y�&)��o�U�6�����J&	�{�FX#�rv�����5��q�e*� J��	�m��-�+n�2�A^!���H�"��&���oŌ����x�z��k�)B�ћ%i���P9�fj��](qOEgM��$���R|1`�Z ���]]�U���������͹˳�j<�[��8:�;�6h��!O��pՈ��|m�����&SIL�uH�0���V\6�ʿM{ek������⅐49�06?�����H�7_)�<
��,e2�٦��������Z����)��t��&�3q���7Z������-�>H���.P6+.��*�,Jl�)�o�s������/,Ag`�v��H�`7϶�7i��G������`n�
Hn���\^���|�,�v�=~���&����֘�]A��)�K�7�Qj�R����Xk�=�����#��Y�.ŰR^y�{^�������x����DZ[�dDpyB��AJ�����qN>�]3�۶.�}RM�l��Gd~���9V2�փ�?��~�Z�Q:��nt�I�V�s�	��'�7���O~���\Bx`�6`Bh���	�����L9i���?�t�#Y򌡧N�c��O��Yy�z����-.I�m6���M�e���r�L�[5km�!�;E�,�/��C�*�AI�p|{���7.��`]��ؚ!�%	����)N;����?������ݙQO������2$'���BLQ�f>Y�ó��Ш�����p �"�ค:���ʺxW��m�G1�r{�_��(+��r���W����trD
�e��Or��T�T�rC�ڠ�y3��:��c?�-cn����~������yW� ��(:D��/Tbk@�*���
�?�T˴�B��� R:�0�+�se�
�압�p8<��7޲>�y�B�[_��%� (]K�E����k�g����Z���ٺy��G0�Jo3�pO:���9����nJ�:�/���[�ʟg�?�eF���� �Z��@J'ՎjYzr���y���#�6����O܆�K��Md���d���*;�̥%���^�IԽ칣��k6*�X���~�����t��0wkT9�#��O����-_0��p7�N�uQƉ���);�[�b�@0�	��S���n���w�ҏ5tݵ-����}F.���@��ԭ���)����Smy�ʸ�k������?�%jT��/<�DW��^�'Wݼ�znJ݊	�x�v��r�4$��$�j
VJ�2\�#Ǐf?�m���6ﯚ������a���N�RyC�jS5g�2�w���v�_P��_��
������{�Z3X�%Vy%���L3��k�Z���wx�S��9�Fx<,�!QMO���!1�ٯf���%��E�6gS��Z6��*h�#���>�i
��_�L�Y�_,T��m���K�+u$�n{-Ǵ�j��|&B�4�](�ܚ��6���:,ykл	��,b�n��g/J�ݹ�	��&߿�ش*�rf�i�d�O��c�B)�����ݾ\�4��`���ׯ�R�i���~�?>�GZ�¿}��b�&�:��dM��5��8乞η9�o(6����Tٱ̌�_f��|��H���hD��L� |`�3�V��;���`�͞�4/�P�W�>"^а��q�^�Dpi�, ��A~�|+O(��@ǰ募��R����{-M�eRzѡi���8;����5>U�f�8� !��AԦ��J���y�`ʰhƷ��o?��}�k٭�<M\�g�����B 6e��"@F���%��i}�b y�DP�#���#�fUٜ���*�5$s��h�������U�:g�h�`c;�D����PUʙ�M��%n���ώ�&��U�Q�9P��@����H���q%[��,���9���kq�����@� �~�[��HF��-^��. (B�����0*�ƒU.�45Oebh��2�!��]`eȱ+��b����^S^F�V�򧷳.���R-p��"��c�H�nY@W�n��J��"�I�����F�Ju�V��yXf���6��#��A�k�'kՈ��^ȸ�7^���>�7og�ў9Z���T�s
_
��E�fq-�&��ݼ�:�i����ط&�\{�Q�$M��_�m���$8����'���s���R�� ���X�#f�P[��F?�1�tYDb�e���SۥRW�[���a���:�oǙ�:i:u�V_t22��˚��bݭ�2�~�����0o5��Oa���2��Zw��Fvt7fz�`χ��/4�������ݶ��<���U&�H��!{��دE Ԟ��Ej�Ⅎ�n��f�>u ��x�RK� �¼�M�ZJ��ٖma��:��#�D��>�$���:�xu��O�~�	����JYigc��)�&_z"�̨�ع���rz����q�y���� 6k��+c�X�i=�xN��ٰX��s�]Z�� M�^�%���b���F�x݂��z6&�*$�ѣ�zo��ՠ���4�L�����u�s�^��
�T��QK����Mqţ��ϸDӦY�L��_�s鿒�l}�)��tN�kS�0y*t��3?a��&�#%��-�PN�g��o$U�Ɂ�����D����XZ��QKQ�J��$+�X�ϰ�+�M�P�>?NPpe�w�d99wz�wi癭��A4���ؔ	,�O>Ô��fM[�/�cen0ѻ�b�o:���K�-FVx7����e
�dx:Hɡ%�|�VZ�0$�]��֫��!�� w��t5�[��J(���y㌊���?�*ŕ�ƥ�R9���;9}�Y����:仍�xҶǐ����V��
�K�A�l�B���tF� Vڿ[�£�W�Y�z'2[��N��ڪmi��aE�=D�a�W�2[ޝ��q���|$�NU���$��%�͙�6v�̴�m�0�L�Y�|�|괪���%x����/J���3�{�!���}hVm�#_�r��p�������B�	j�����r�T�#��Z��c��GSfM�P*]�-�F�3+��Α���Kh�:��H����bA��U2��^_��c�vZ䳞��nu��]��?Y�0ou1k��4E�܎�O>*U�g�R�#lC��sziN��Tɩĩ(w�f`���m�0�8Y�ye��%�[R%�W���rq�E�_����t(CG7��U��k��8!U�d�z��'=�C�����Lg�mJ̻;�U�٫���3��y�df�~�y��U%޶�"��XvP$� ���W��Q���5,��;\iؗ��g��qv��b���L9>.�|@��!Z��Pm�oE�;T�\����B�a0T�W~�m~�%0
�X���0n6��
��G݌ꈳi�2���xc�kP^9�,`p���6�v��P��;v��T���n�ZA�ei�/��(��S��:h�_x��nW�	���$r%-���eM��Go0��x�;Z����0�2)��[/���7�X� ���dƺ8����2](�ɭ$�� �w�ޟ��!
��@��B�?�Ċ�S��zԩ��TW\\�f��,3���=;#a9bE���Ё;�J8v.r�?t�Ax����,���E�����P<���C"c�מ�������&>��f"��4vi�?�02����#|���ҵ>A��ǣ�F�o>��Y#��t���6��<�!Ʀd&�Y�(�8[�U�J��P���8��B� #�K�%�^�~R!29d�U]{8�z�����+:��6!'�#�P�J�[
4I�Ѱz���0��c�5Y_�v�%T�C-D��8�@҄q@�+�&J���N�Y���a;�>�R X'���2�۵�$����<����mLǱ%hl�Հi�0��s�j$ʾ���̡����e�\#F�C
4�K�6�O���@���� �1Ӕ�[>�h��CP ����cGC�������*���=�B���I;լ ���ZeΈ��z���[1J�j�M�98�f*N�ޣW�
���a�}�
#�l���z����}��ėnY��]�2"���ԘX�z.z�>�f�q�-N^�s�;��ɷ��0y�Ri=]ǆa�Eu:�1b͖&�C/=X8>��uc�H�`�HzG]��Lڡ��L����uX�-y0���6SA�pyeg��?C�2���I���t{�v,۫����3��{JNG#/�6�p�B����xT:Sa��Hg���ӯ���F�6"&|0h����3n����}V�hkf�t�ZV��SD5?mu:|��7b.=
��y�����>4Z�����@�gc��	���>�⦪�J���2�~v���N�������ò��dt��\�S1��A_jO|����-1R� �l�m�ܾ�.�l�;�^g�y�aC ��]�&���6����ٲӪ���/���'�	��L��h$�`�L�k�d7q��]� 
���1�6��(zZ�K�]d�&�GA���Mg�C��'��>D���uC�Q���hc7��B��f/-U�ZKE݈9UbP�u�)�
Ç�C�n(u1�ο3�ػG(45u٪5�Ǖ������@מ�&���O�����8(��%���J��X���6bW�
>�l���:1}!���z�07��a��0,�F���$�A�L��-na��5�-E���8�d������SX#��mJ�D����/�w��\	�,�B~pCO�-n��}k�F���v�{	ܑ�ոY#�'�AA��L�2��ޙ��#oa���m�t�l�Q�����S;�����v�T/9Z\��ۈgr�U�M�WE���X��*Տ���f��<a�K�KbĒx���F�$ e�3G���u�;LaA������� ��= � ��}>�w�M�ח}�	��G5�M~5����m�p�{{@�n�'���I,�(��əY�D����?�i��A�QA����P��P����K]�W$	G%��Q9�y�`��g����~�O�p��D��<y5�:b��*��ُ��l���Z<��iGt����@pS>���b��&���&%g�\���~�t��	�<�0��Ӊ���Lq�[��VJ��e.���v�p���������.��ӹ!p�p_��4pJ:�004�7��6*XU�S����uȀ��RoF֠�$�1ڨhz�������*���k��y����#<>Ύ&�矩W���'�2��h�o�]Y����b�`f�Q���{�,����YB���;��SZ:�VG��p~M���>�~��g�� �������F�A'�g*��H ��T�HlE��_U�BJ�L�h�N�F�F��Δ�='F@�G��$�#$�4���\���e�g�j�EܤR{2S�R�������s�e��pۼ���i�Wy��^p��]��2�
�H@�eP�!��92� ����m���]斍k:�X*�&��C�O�.N�`7���	�	�Z?�E9K�r]��@4C��QŷMjОUr�+un.��n6�<5�؄�Q�I\"��<��'͙")1 ;P�2����,�[��M�R8�c�:b�O�^���pc`[Z�"�@ []���!}r�՜�,�:���	tӍ�h���Q��a8�Z�Me��{Z�?��h�L��vp��l���'߽���>D��}�����G��+��TChU��	��8Y���z<�j*�'̶5�����Ė�ޝT�q�|���+d�ﰥ05�n�)D˭Vyzf��w�>�:n{��I.L�&�&6N���Ш����9�܂�[�rՖ4)� �sŰY#6ns$�}�s�������b��%��5.���`ˣ�y��ܶ�v�C��]@W�r���B��jƖ�2ά����ؿ%iR���)k-�@n3�$�
�0)��c�[�iv0�9�Ow b���qb5�2�{GEH�ȡ {=����M�GnuϞ�xTH!j�H��Z������)"�G_3;���z��ǀ$�;�;ue�N��QF�����Z�L��1�Ǎ��8�M��\wF"y�_�1.pK2�Z�?�	���tx�GaW��qjvfhL%�/R��b���'�� ;%2����^��7ܻE��BYZn�<*�P��_VMU��|��"W�M%����*������RTAZo}A:>�G;r�N��f��5�A���?@��.�]��X���;MG��,5S���׮o��j�p�E$�a��D�>AĂ��Y.E�Y�I�޼�ആm�4��DcJX��xĽ�XwM���6BB�>��g:<�Ά�s�e8i^����*>U�	h�r��b �ϥ���,�����0��,	E.j�=��hk�x5ŝ�K���(�i���/[\�mz���F��KZ��f�����w[ޗ3"�p6������*S}뇄� [3b�u�IV�(0�1���A��ha��Jul�.$z�\Y n�i܃�2�h#�M���j#���dn��p�\��
f^�ǃ��@�O-1*}��-��ӿu�=';��\~�]G�b�2��]�����)!X�]R�ӟ"I}\T�z�ڟ�2-~F���P����	��E:L�1x]���������>CkQ�U%��f\/oƬ��w&��g�̽x�f��<�0��!�5���+��5��=�&��=zR�[JBV!����ݦT�=���՛��ب�󸙚�v���"�c���Ɲ��|�@����Y��`{��D�G���p+��>�;�����`9iU�z�?��H�_�QW��C�k����d�p��m���gS�В2���e
z۲%R��V�=E��W�Ag�yx�s����<4�W�gn�1+����H����źƸ�X��0���r�ɂ��%�y.�F���ܬ�6�����_��V@8~�E6o���P���4�PA���rSL��d����Y�7F�y(Z)9���+M�K�q^:T3����w����v˥M�uQ*�a	,J5� v;�|A*��dr+(���[q�|3������=g>�7�A�����H#���n���7�m���i�Z����ј\�n���kiHǕ����[����B�?)U}4:����'"�n�BGmBw�����<�/?�UL˙��̏>����ȫ>}��U���8����AU�
vP��j���DQ񥓵%t�*�+S��#��W��J��-�C�0�˶OSȽ΁�� T2�y�х�y�X��"�EKK��S� W��p@,)[�$x�t[��aP���xY�n�p������QT	�0V�	I���>>^��8��颮��n��}�W���}���Ґ�A�a_�?�La��|�k{�I�ίC�:�����J�w���.�5%����\4J_|,wD��(����v�z��xk TK>�ͬ����_=��������l�����-ː� z�nM��[��b�08�>q4�L@j��@�	)��0=�A�8�; ���&K�?�.�4WgN���)̕�M���jX��5�B"z� G߼��m���۝^���XĽ�,�rZ)����9g/�)�̃���R�%$;y��������E�
(GK@���~[C8������<���"���:Yv�d�,�O�8�H7�h̲�+-�=�6U�^��1��pBs���sh�<�!k�̀�ZL���dL�KEA����M�ƙ��|`^��6m�n�)o��j�=:����Ƹ�T�fnOY/[N�����v)��dj"J� �9���z��=#N�1��W ���~��X=�����U�����D6�����C`ş�e��Ƿ��뵭nj�vZK,�T��2��eWwm����FOΠ�`=lS���}����n˄�uP_�R��f2tiKFl�����\�#���S��$_��d�n��`�`�N����rgbc#Nl�T�q��O�ן?�BvW4BT�V27r43SuD.��ﹰI����[�(������� )�^�.[Rf����A�Ⱥ���A� /]2ڔ������&�d�(<�_�y7q���t��Օ�����3�D���ҙ��,���w4�\@U�Ƭe���'I;T�.��¢���<�4���6�ٌ} +�]�9Q��#Rj�C����u�_|��(=�E���Ě�"z��c�_����p���YN-���宊��h��c���R�́�,�f��]�I�x�C�%��y�� ��������ťL/���
���8��[H�g�Pm#�_��� �@l��o�$gQX���G!��R�Vْ����tf�$����������h)]=v��Ydvf^�b��H.�86�f{Q�"�8�T�~DC����� �~�{�3��&$�?�+�,6H�D Cu�� �ӣ�f ��rţ����ښ��S>�p a=IX/��L�[Н�ɜ=b/�8ɓ"�P�
b��
�d����1;t$��%�ur��+h�|����-��!V0jR�>��#��	������%x�&<���g�-vt2V�:�#�w~����$K�+,��,�nS�G
>�߽���O7x#�x�R������z
��$��ګ�@LxG������
!��������,2���d�"(��R��x.M����Ux��5m���O�E[�*�x4����Z:14���c�I�R����9;���3����g.i�`�I�1X��8z�|pa	te��4pޙe��kv�S8y#L3�����Jhs�$��o�
0|��01h{:�\���xjI�oe�Ȫ&V���H݃X���V}�"�o/�2r���Pc��:/�B��"�O�XoC���h���;(&E���`��L�t[���A�O���z��'8|R��+ Y �?	�{%��,����.��A$���*��[�\���E6�/���J =fN��̋��b�'S��²Q�"�#Դ_�豁
�b���>=�c��\f
�H��'9qŴ�+Ȳ�k*9Y��Mrk���Z$�8m�� �h�=�SP����⟤5O_3���"ˋ��^-�W.�=e����2�!��L�$nDg-D�_��h�Ɏz��zQ5�n��c�&�S5�}HBn���+����svH$n�5Z\�w�B������*�D�vta��B���14,��`S��g��g.� ��ӡA�c�oL��t/�����+�̆|<�op����o��6>�S1��}?=�j5#�{�������(w#�1�FBp�aF����!�OȎ������U�P�^eVh�n�R��ue��ᇰ�]WYƬ��l�J"�HA�%ز�a�b�Z�~ҞG28��|�(���QJ�^O���P�G�u���L��]���ɪ�K��N[#�9�+�1�g|ګ��=E�T!G(������	�eȃSȗ�_EtL^lc����bS�w�I�t����_���z_x4����'��gD+�sџl���`����m��_,=�T &I�R=}�w�t����@�	��kYe���z�߾S������B~\��=�F��(����}�	4�(�^��?׻A�Z�Ԡ�s��	H�}�����P�=A{Q�����(��XY;a�T�bN%0�l�9��Tu��3�*oa�p�����k���=&���oGݿɨC�|8
�¢3��WͰ�M}8��`� n�狞&2P��,�Ǟok��	�`�����Sb�M���?�(˕�M�{kf����{!ٷ*�*��C7_ ������XPQ�I�8͎�]gu�˓D�k`�~샔�s#�{����ʡ�}�~q�W��n<@�LקF����{ɝIc�{Cѯ���{�4��r��(���q�v����?l=e�u��n���ʕ������*���1IB[D���er��`��5��.ј�����?�CqL-k:2�d���i�Ƞ���Kh~�"%�i��� u���W�����޵]"�)lG{��`�p��Y_���=˱�o�0g�o,�q`� q�q%�����x�oV�{�������=��.W�)+�dܲ]���XD$JB�Gs��w�M�J�����w柜�ltyG(_i�KZ�튄	.�E��ǌD�l�&�ff��i�cNWݶM��k�ޝ��5���!%�A�� {�>i!H�y�8V�N�WFF�O'=G$t�����*~]+S��V�8P��-�6�i8j&���J���txQ) R����x�NE)��;�v�}���C�|����:=F��3[��8D%"La^G��U�Pz�:����b�B�J.
H�Ѽ]y�n��/R���zF��V~q�:���V20C��9i��� |V�E�-y��3�`���d��D�j49��t�mp�3Jzě�l��8-w�8�"�wo�v̪�zDߴ�.i��t�	�[����,��\���B���e[�}�G�.w��>
�x]g�n9�%�u��T�l�Mz�o��v�?�C"�6��K�s^�0y ��P����ԅ&�PFi����\�#���ZNƝ�ޅ��}��d�{�]��-�	�e������w����y�.�܍a�.�yf�=�l�s��ҝn��.j���|L�'٪$HvW2���>'!�w\,�U�^Bĝ�Y�Hz�e���n���6_p�Jpu��ޘ��*��d���*uE�S�O���p����F�BA�r�l:�������.�mU��P��O��N
������$��)_�6�25��U�%vj87C����SR<u.�]^Q���E���I�Nh˞��Σ�s�]��:����@$k({.U)u���ވ^
ȧ� ���Y.��g�NHL DP�K��`���X��×�N�jYd��"���4�sb��N>����θ��{¨�W�DD�A񯣅{Kҕ6cƸ��J�^j'a� �r������6|�ۈD��=��Vs;���H�++��*ou ���J>p:-�-*�E$}\������ԑ�-�r麉G����F�@ҿ�NT�C#�32e��}&�L'�3I)C���h���J��f7�ժu�Ų�������y�4��=�v��\gF��պBJD]�$�4�	�/�vZ3I��5��9�E����>�\�p!C=?��("�:tXXT��.ph�KX��F��^}�q��IUs��t��������o�OuY=�N�j���`�/ \�Q�f�K���~�$GG%"h�qZJ*���M��53e}"�M���_��k�k8��k{V�Le�3wn�
$ �3t!��T�36��]Fc��Ÿx���ݩ�.�iV�,F����7���)����_���vz��Tg�p���2a�8c�'c���T0��M�E���-kA2uق���u+iWC�nN �7�#����:/�B#�D��u�t�7~6�ɫ�Q���rW|�c�w�/��d��u3�|Һ5�7@1	�pO���-"�������^��x���O>t����Ў��U�z��H�OhKdE�Ɉ��ǕtZl���{�N�cj�)IP��R�d�Y�S5�X�u�s���RXlLݹ��|5�[�8��1��W��z]��y�:MUUe�6�_F�^,)�"�r(O��a�Q�]�h���C-��&.=\��$X�pm�P&��� I�h��~.!^����Q��٠E1zC��Iu1[��-r`zu�t�]A
��?�����:�X��^���>��1\H����w�W�cQ#���bJ��35���qIa��� B�����6J���=&.��X�h���U�v��%!SUy�\�s�8ON��z���RF3�'1c�Rg5�1��x\۝{AT�]����iL�|�m�c�B������c��ќ���@X�Ƴ�u��Q��:0Y�u��i<h�}9�w���a��=��i�{���蚋�I�4�����`��6'��[UQ��{F� g�+q`�H!2Qq_�]S|�<��t��2:�c�e@�Drk��+��g�?~9u!]�=.W:]݈�s8�:5X�rz�L�&��1_İ�y�$��H�XѷNl�&��l�oh�_�����]bbP(uڒs^�������d�_[�]5������0O��j\N�uV4��Km�t�x�x��2�B����p�[�㶙>�!�s���^i����D /����6�_#�H�h�s9���F�J}=QQ}�{���Z�����"sD�2�`/�\/�lQ��2N>��x<K�ڈU���(%2����������f�	E�"Rb*'Z>U7�ڈ �5O���K�s�3ah>���(�qh@-���v�s���HBn�5��>�RU1�G�!k�jڢ���a�h����A�c�H�vv\AUp8�	�!D�ʹ�Γ���n�?P��1��M	 ��
6V�h^1DmY'�y������7k���}t�5�B���ӱ�f�󣵂%�� 
6��YQL��o��>c����D��B�Fɳ,��<�z~C���f���,7��V�l��-v�T�-��O�I�8�E@z������4����p�v/8�0 �`$�|_@�~1�k!_���w�V���~��	�	���_��$'��O�b]��S�(��6���
Ed���W�]���<n�N��{\v��7Ie_�'*? l^؂���H��<3ք@U��/����	���I�W[��\�>���7��jc�:@�˾��%O����z�r"�e�T�����S�1e l(�z.�����~*{��i������H�1����᫭�"��j�@�wf��늈�A��W��|5݋��c�n���7^���օ��'%���v����i�`fTp��G�Ӊ�}ck]��V�^���ب����
t*0��*�����X��6ulM�"�;��7M0mjT�C��a�l)$8h� �0�C��#�!��K�π!IZ�T�62v����v�pf肺�{�߿EW�փ�ǌ��x�
���ji;�u�*�(�B�2{A0&@��D�&���Op��$�9<nWM`�>�Uֺ(��Ћ!�9���4����W9��پ�X���If���8)���W�h���,����i�B,�v<���M�Շ
���~
���8�֒�����)��d�m8�b]o�Ǡ [?��d�>�_+{ ׌�����dn$,�wj/2��r�ޞ� ��5z�	�>&M��n`ގ��,��Zzk�����f�Fo�A���.�b�oڒF\JZF�0�"P�zra QiC��b��4H|�9q�u����9CN@������[G���®�Q����S����k��`=��ek�Ok2ո�}�a����E�;�QA����.�.d#�B��G2�;�t�Tl_֘G��^���E�_|��<<20�	Mu6���І�z��V��M^��zF�?lW�N>9�9(L��Q**5�8��rJ�^ {�j?��B�����&]�X��׬�n;d��xq@�<��c�@�TɄ9�/@,�����ɜؚ����
=�K�<�������&g4��3�k��+ܗ�}�ح�V�mY���e�KyS�췹�$D�{Rnc�r�Gl�����	Y�#���OΒ�< Ђ���'��3|M���@�j�tzfLr�8?=��$|��=�X��<T
���'��LFO�9`�/d�i{e�mDB�)l�Y���������b��W��P5��P��˲J���a�4����8�t�R51L(�\��@��d�s;�:����}�D�U�C�NA15�f�;ױ��4ULD!��LP�+rS`;�Ί�u���)����RCIu��4�t��B3��_�%����p����u6��h�8]-U���w�An��<���f:�B�D�Nъ��?~�|,°���?#Yl����?.b�6��^�Ak)����YA��i��W���[�����'df[�����O��<�����C*�fe��&{��U�c�|.�Ra��x\�0^��I������r9�=n�����5���Y34ӽD3>�u���+)B֨}@I�}����1��p���Oo8+��पZ�K�q,�ִ��rN����'�����y͏��D���y$���QC�N�N�w[|9��e�I�#a�H�v��OB	l������^E��xBI��_�Z7����3�wV	�Pϊ�HDU�Q�4���h9��=�P%=��e���=�F8�0��HV���Ff�Kpj3L�-�>J:�
��t��!��'sʮ�G�u4��ӑ����r(��H���^�y�o*�Pz[�.O������)�h}����7����VC��|+�%��5�w��|P����Y�TT�>ʜF��ύjO�m m�M���<[�(^�̄vkU�%�S�P��m���w���P�y��H���Ҿ3k�V��u�$�G�;��	Q��Q�hӬ�'B ��y���9 0��}{F�ؽT�SHn-��V��r;+۞����$cr��G#�X#"(x38�C�9o8�\��}W��D��ƔAۘ��¢G����t���'a�)!�R��+,���w[b� �����Nm;��mm�����y@�	�����Sz<#:W����Sͪ����B=��)��_��=�̕�c�I���|	��X��;�v�\�K/��((q_P��tL���U�q-e��b�4�Ys�ގK��!�L�b.� q������]��7�j���鑟�D���O�**�}�S��N�H�F���>��/*y��~	T��Mռ.w���(����&���>*�W�j�Q��lL�����]�l�a���q��]qr:�z���N�py��J�rЇ��ؔ���^U���h70}d�u�\>:Q�~��*��[� ����#
���,�]�שc��0�wG��W�^�v�H��Z�(�����_�B*Y��ڃ�i�0 ��jy��#z�4�Wv$=ƪ��3��̼�+_ޡߟf�Ȕr�����=��S�RG��2M� �]Y�����ᰂ�$���s�@��q`����"S�%�������x�`�����A�[�i��/)�%ha�*s��-4{b��rA������0��lW|�5�f�,!�}A��N�36cT�ng&�(��&��=��)���$ܻ﷉�A�p}s|�+֔�gE�{o/`ƽ$��"�q�,3�(�l�_de%rb��������i�lN�K�l��&27	

���y� i�~.q��tk��)hV�z�z��g��H�(=U4�\���y@m*B�[���d0N���6��w��ʅM����m�`��J�QӤ�q� �Q��s��/o��b��gs�;_��-�-D&.!c��)yl=����u�D�����;_��q�pd� �RD���!=V&�*�]���.�������3��?��N�d4�Ȋlטݫ�ha^xO��r�s߸��p�&S`�bON�u�(}��,0
���]��4��oM��do�T�~��:���Xs�d��w�'�0ckkm��i�ۜ�`���*������؞�b�4���}��O�͢�Z�d!~ل6h �������V�'u�
R�� �?�ڍ`�d��xz}X�����]�QM4ǿ�ɍ���d��g�m��,լd������B�D�5\�1#�ްΝ̰x�^p��T-����Ҩ���b[�8	({^Lv.4��{�vIɣ��iH��Z�\�k�G�6����x�J��3Vdz�0�7ϤgơP`U�6�H�U����MU��d5N%�褉��;�oB������[����/��Lة��Fh����L���K(��P��ƭ=2�rW���E4�z�D���L��?��)��oI��O��a�5[v��<,��8��=trՔN�԰i2�Fd_v��#�F��E[�����퇦k�|��'\T�̓����>u�r����C ����,�摉���~K���Y�D�^za��� ؟:�G�@ U�H���Ǆ�XV�H<�Gv��(i̸q��tř��ךo�[�o8�~�P|uغe\�jiBUހ�BS=�{ܹ?�'���H=��4�m�B^bʎ����g7���s�d0��!Wק�{�ـ�n�:�b+�Q�)J
��0�Zh�Q�i`0�/pb�;c{Q��灮�K��&�[��+`޺RD�-��F��I�~�an/�01B˨͜��Բ���:�F�.�K�]#3�S�!�n��$��_�ڇ_Nk�.ٝ��v�DعIVr�1L�m�{w�ĉ�YG��J�~�C�����.	�^�)hm
�~���Մ�7N���`�Y7^���O}�c��<yK�e��^����7R�_{���=iWC�3�O�y�m3�z�fM��9һ]O�2jNE�}g#�_����ؓ�RQk/J��=���)������hZD-pZxG� O4���ng�z3<&
MtycC����E@q�~@�-��L��>���{�eb������m�n�V'x�F��
�Nդ�l�7M�g��,ƠLP��éB�+�f-#��Tw|Q�@������p eB���g8��LP�DX�,4�{FGޮ�����>���ť�Q��kB��
��j�˷uwg�:��i���� )�q=�b("�C˚5�E���hp�r�b(���~��0Q�w�����7+�b�:q1��2YD�+�IV9�(��U?�3�r�$T �� �/K&]3�C$��n@�$�ʰMߚi�"�]������#�VŒ�n��u"Bvz�w�J�5|H���H��=:�I6��ȗ��Δ@�鳔!�VC�>pD�����F���JЈH>Cæ�孾���w��O�&�}l�H��V�/�2_��:�AX�V?�f}��G���pB���+���?!�T(�5�,�$:���*Ns-�\�:�w�Tuk;mj#(���gֽ,�I�r]25O����E�`����d�| �� a׌��:�66�ׇ}��
��W"�;�t!Ƈf�Sb[T�Oے�޵*��o>fn�%AI�qMp��B0�3N2�M�R��$�*;�D�u�+�>����0��d�]/�����}u[e�j�k�=��mܸkc�M�/��(	�ǩ���9�ռ]��}�5ڎ�K�n��ѾX#Y1���Z��;�-�Q���R�� A���x�>Y��lu���я�~�SW�T���ܬ+��y��t@�����\OsxS�m�Q��C�;Ǆ4�y4q��Ck�`t�a��V��󕬥e�6�)q�cm�[~?�\����o ��*`r�O�K=EUL&�~�^�#��<�Iz�GA�a>�7Tn���.���Er����g�.b�����W`�-�@�-":O?��r�r��,mK /�AT�S�[V��Ige�T��/�P����d��q�f����d_��u{[�����H  rl�*0��/�܋\�2�7�9x�H/�{��v�CM�~Dڵ��=�3x�i��nx��Mm�U�֭�E�l.^�ro���u��PB7�ݥHoޖk���H01��GE�: x!���k�_�(m���bžN����4�n=��ۈZ7�뉠eEӌ�*�7X}��_�;IviN"��T�c~ݯ9��ڥ�^�9~6�vA� �����8
�o�4��q?�/M��le�}��xuS��d;�����;�4�⹅yُǛդ+�߿�6;�6P�����1�gUi�h��m�n����pV���ͥ(��)U����:*�g_��?�� AhmƁMK��q��8�
�g�ZGE+MI�{n��|.��3�5�� �<Uc�`�B��?�z���</�R��O�5�UX(X�7�����G��霒W_u����	�V�kH��� �A����*�؉�/�e\�h�����Vvj{�z|q�[U��߫;�=��`�h"�Xz�Jx�T�wLBݫK�	���4N��'R�����_�_�ܭφ�g[-B5fY��I�"��c�e�Pf�Ӳ��a�:�C�+�T���[�יi����`�6�66S����<�-6J����7�b�y���4��}��B��d�g��.Κ D��Y�����A�s�V'��ձBp�	�uf��p>�k�K6��q~,��^N���$�w(��ݰP����!��o��%�_.�|8��������;>�G� e��<�0J&�,1�`��<;�2J|7�E�O�
%sj��z7�(������a�Ĭ�G�;���o}����� 7�{��~)%���:� ���nX��|��r��NH@�q�v(�G=�V��d��4�]�v�6c�"��$(�Q"����tR�~~g�V��Yf-�|1��Ma�*f���T������\�;���z;$n��`��*Qr(���2���5:9�"fT��!N��F�o�O,UM�տ2�eg�ZOQ���t-��R"���*)�<� ��|�^8oXݝ�~�̫~y�_�zظ���E@Ô�o��O%B��F�:��w��9���f-ˮ����UA��,���51� ^1c,���=��c'��TwAh7P�-B��T��Ӄ���p�8}	�\��M��:c���B�
�$2s�C������A�)�bH�u��6��q<��p��W�O�>��	�}��ڵ�9���!�7��l�e<��>	����: ̓�b����`���*��m�avy���!�o�	 ����wn�H��?��x�)'����Ƙw@H������S)��	����d$��O���$B5�~[g�Lq��pq@��wS�s�F�GmK��2.�-��k��<�P��pj��(!��0���会 k�>�}ѫ���=��:��O��ض}�x}�c�d�[�$,��㳒��Eq���R0��D��C�)܇����>����?�B�йD�,}s�1�B��"�wC�It��V��s\g�w1��[��j#ci��4 Ç�,A����$z��!|�0���O	4�H�t�8L�BJ���|?/	���nj���.7/�iZ�$|������VJv��7�@�������vFn��L�1�:]T���o}�����}:ɬ�%���+�G�{�r�|w��M#u�/VA%���1����^Z�5����m���ģ4E��TV5�^��۫>�Z���Nd�@��L�n#$�6 P �h��=�:	�Lu\�^g�.�P���71�)W�ö`�~�z~7R���z��vL����Ѣ?V�!4I���صU��=;.,�ĴR2�s���+��)���9����-?���ȥr��w�=Q��P����Ei�b�߶���j}a�&�j�A�Ƕ�`���6�țU�ew nGJ��7ۓ��@�U��^k�[���$;3���w���C��_���#�t��u$���x����J�����N�o*�Q"��VQ8���
W�Nk��&�-r��zˡ�fUc�8��� ��?�
�_4|���ݦ��w��jJf:��V+&����[P����	�U7���T�%;�8�<�Y�٩F��I�c��qxbO��ġHk�;D�	B��-pE���HM]�hr�)r�i���k��o|EF�\b� [���*����
̨��"u�kF*Uߴr|G��+�o������b)Qy�*�I�ꟃ��3ó���I=��&A9?N�HR��+�ϰ�	�g4d��W�#1��d��I�cv�/8s�w�as���Cg孍��nwy|Pz�d�`Sg��4�������h�n��,�Nc��n��)||,X�t����8���x�W7NY����l� �/����u,-;`�M�e��"HŪ�ک|��"����z ,��^=&PKQ�wVv���R�Y�EEERX�����T���i��T��=P�֝YѶ���_v�~C�Q���N� {F}���>�d΋)F�ձ�O�EX��<�{J�����ޮY��B�Tz��FD��{�a0�4����vi���*M|�q�����t��OD���	���*��eZ�x�vC
���`�uE�
���{n��|�22Y;2���@��u3s_G!?���ښ��.[�+���`�1���+����s
!�7a����9¿V�����D�� ��x�}$.��L�wu�
��c�$}R��p���{$ƅ	��W��<g��_fx����\$>�s��a��9ኾ�x�:p|u��%�#Q�َ��+*�T�o���eO[�>}�ޏn�L��_NY��9,�QH��37���)O'Q�� �	�S��i
d�fг�s�W��n��M��H|���!���X"o��ĊW�8����o�	f]���ٿ���uc.�i:�q�B��#2��\��9�<WzE��.�����7�9���zy�\�5=w����ml^75��������x�と=�qo1��,��~ݽ1���ؕ��S�I���j��%��[V�C@�0�f���E��	?��Lb�k�l��y�Mທ��	���>G,��svVRT<y�9�����@���&f,�L�;�3������̏�5��c2��׬�wb1]����:DN�S���q���ﾪ���ɩ7#�M��>�'sQ�W���${h#��F_��Y!�ܹ�.��� A/���X�K��TT�n�#c*�ͼV]���{m�zI�����Eݬߐ��J����J�ĉ�SV&ֽ��7�a�)9�vS��Y���۰r���C�� ��/�k�ֹ�X��Q��l�r�y๞�q�������N@��L��@����6�rTi�I�\d��/��>��j0$I��!6��=ÖЎ,��"8=G�vC/sEq�L���:N~z���|�8�9��l��tjNz�"��4�RH��E�2n&y�����A�'P&��']LH�D���a9`�.�iHq'n�UZ"!�%2rҪb�$�7M�b����l�?��aX<=S�Y&~���"�/��`��r��dz�-�u:&[yHw�$�a�_���@{޹F�YSt�A٣�"�d����0��ʋ�����#��ׄ�
�P�6����"s�o��)͛�L_>��W�[���%u�e&],N�!��R3�ӻX^�W�LZ'Y31�	�>½I�e���v�,U|�{~�0�[&w�ص��+�9x���*�{H����i0Ŧ��ִE�i2ؤk.PJ��cq�@����IhYjN���!���Z�/��߰v��^*)��-\ь�h��rɅ���<�Lt�uJ�R��W.G��D���A�(5-��ܑt9�w�1�*8���[���M�N>�ݧ0ϥ_e��G�/3�P������k�%�>C��Z�AV윯s���+1W��+���Fb2����_��5,2��Ѓ�0�ݖa?O�yR��^+�.��$5X.���%B<ա/}�>�8�m�"�3�����}c���~+��҃��qW��C[�ɘ� �`���Y+[����5�:l���?4�b��y@��ԁ�!]�K{��ϵ)�ͩP�&zh�FF�K����aA���U^�#5{ڰ�n������c���U(�M�Q����>1!�&>�c0R+����'��ط��3F�P�N]Ŋ�,4�|��q�����.���J�P�-8�Ӊ�y���ojF5f��[0|���ʪ���\�5~C�%)t�
?l��2�w�@�B&lj� :ޠ���P�1�'*Z�TX
8����8I:���.�2�e�#w��R<8�?�IF�5�E,a2}���T��m�\5O���x�L[���P��:hf+:1�6��NU��mJ�֤���a��S���L=Г������p����ZI�Z��yh2-��X�,�?O������?�*�V��~-w��5� 	%&_�E$0'�g�NLdz�:��c�J9`9�� ���ib�w,��ia���"PHT3V�IR��	-��F�p�d\�
��-Ċg�����Re9�-�U�9ud{�Cv#{Q�DC���>�,I�7M)��
ba�`��H��T�.H�I��i���x��	gq�AD��K�]СI�	�B����w��z���L�,�G,�&��y��I�)C*��$��@�m��2r�)35��)kPX?g���x3.\#GW$D>��vro��m&tǣr�ľKd�_�֘��8z ]v���q ���s�C-9�ÿEa?	�|���$�����k�O(���G66���ا@�A(�x�0cUgK�b���k�.�&�uҰ�+K"�~��T�9"-���#z��"�*H�D����)�&dK<k/�p=�|�J��R�	M��=T��A����r���*�΂��Q���K)�ڞ$7 �d�P�ps�O�82����f�(.���ئE�6�-�g�{��<x��_��īp�Toʬ��0a9M���ir~0��0avM����(_s��GZ�� U�T�Y?��Y�,gL����,oŏ>#��$�V����7#��K�Dމ �j���M��30h�ď4i'w�����.��2|�Ƙئ:�J�>��&��Y�qTDߍb���%0��XJ�o�pq��o��ĭOm�^H��,����X}d��243�F:�#|�&n
P�SG6�C�4r��Y(��4MΧ���y����N�4���=L�>L�*��t/����s��������/8(�g0D޾�d�#ѩ��Y�Nh�=��3ƉW_�x�OF/�T#���,	��+H}�Lp��^-�����3�0O4[������HO�w�;�%�-����)!U�l�@��v�ɱP[�CG�l�Q����(�����c97䝎�W���J{�����6tLb�I[x�I�	?�P�M�ae�3`3�\CA5axRN$���htS�[;����6�����R��T���h�3�,��n:6h���=��K�I��$��8��W}���H>��z����Po����k�ׅe��5���-�2Lh#W�{��3��Ȥ�}[��ub6�E��5���u�+��q6�w���
Cq�_�¢ke�y�c�&U��K��S`CF�}u�p2��ΌP��K�uiw�25!���P��"�>�ҽ�6W�����+�_���%^��)�&��S�������Sm;}����E��ÏA]���"�x�T7;�,v�?
�9YҼ26�Ĩ7����-�MU�0�	mS-�cN�@�Ҏ*�8_�Ezc�B��}��(�JU�ĀY ��}[rl��ٷ�kNJ�m�������PGD��xM���2`�x�^9�]�y�U�<��H�~?�gJ\RwL�\���gjP"1'\�۸W1=Q:���Tyū��J.!^9�iQ��,��Jԡ���76@�nKߝ�u��%�c�f��E��8����R�[-�!�w7��7�JМ���RU��9�أ�NJ�h�#ϫZ*�	��NPf/XJ����T\�.�<0A�x�e�'�"T?X�i�RKn����K��E�!5w/�_;#葂�r��Ǩk��=l6�(�c���!�Gi��� RX�����6��XU*��TXs;" ��P��JW�� �wO�M��!갼&�`���٦��X��B�صZ�^�\x��C_�n7_VL��B.��RU9_�0�H�N+��d�����w�_;��1�`�@D_��w�ϖ�C����3�Kz|�&_͠�K3�`�!�G��Mw�0�X����=����(v��$�`��'>����ag���Q����G��:��h��nm��HSx�p��.Y�ŖS��đMܸ���?g��.��a���_�|bb�@�b�m��.a��g�)<4���D0�jC.��_H�w`���L��>��LK���Z&�.4������C$�W�'*���B��@��Ad�h���F�,i���m^q���}}�����F�������ϋ�@ԥ+��Sr�>�C����I��q^x��G̧��m\,�L#&Qq<��	�2X@��q�gv�߸�+-J�b7u*�+�P��{,�%�/��W��I�m��#��].� �;���/����%L>u��b�S�́�}��1�(oG�+�쑬�_1U��A�0S}��bu��`~BW^I��hd�~��>�Bހ�P������R��`�vA؜���.	��S�B��s��_�^|6���3������A" �d�l�0��檣��yX^fKԝ��"Kp�:��7����l^~^	�n�F�Dw�0-'r[�~�|�۾'��~��-��]6�!��8�0�H��1��X��RU\�"��g�|�<������A��c��C�)��"�WM9�R��̰�}�G-bZby��b�؅�H�{v��i�~�p����8N�	�:�)��k�a���fxNng�7�5�/ʚbۗ�B�7��o��~��z�n}ndb��h�X�jBɯ|��;|w/%���鎲э��:&)u��8@�ݩ�}�:oYҸ}�+JPD�}�3�r�����p7�ccgQ>e�Q��oVF�����O�![�&+�IF�k�3Ku�� �y��T���2 _��z���Pm���l����$�J��g����*�&����Y-�\�����$����Nmwc�(d�h�P�bj�h.1KP��J��QZ����!��y���y�����#8�`z!}�9����yL`��Ѣ�A�vȒ?���Vw���d��R��F*�X?�%;]���,
*�})�V�Nm�
f�a�٘�Ŧ��N�U	�L��+�"@&t���)�'��l���<Y�o�.��3��P�^����E�:��H]b��N�w~�5�+ �� y�/�kI��gV���*��ǯ=����˜�:�-T4ꐝfy�a�qs�-Ƒ�c��˜�W�V����*� ���
�6�[��Z��\
���/%~��H������V�[���6uPМ�9n�����^��콛��*�!M�n|M�� G�Ѥ�
*C����j.�vY ��<�*���s���/�∁P�D뎞T�Ł�'v�H��p�H<�������,�b=�y�ԉ,2!KZiq��p�K�:r�&��7m�����O���x��j�pd.c����������ɢe�!RUP�{ah�b�f����ͤM���.��5�u�e�*�'����1�M­y�]f�a9,���8�f0�y^ɕ�(2OʒK����8|X��XA��Bz.LU���Ǣ<A�w�B؟�H��uk�F�A=����$�$c뵝�4a�LR!^Qw�c�g$%��v����Z���;��c"y\;(�~�ȝ�zJ�Ď��W��ސ��;~ �J}N�{.�7�p���qS�;M:^a�)��u��<J��g�ӭ��v����IIi4P19�j�6'pO}/�]ngU�*>;v�?$�u=�� ���7�u)��eu�"�<f�] �sp��`5-ɔ��֥���k�P�8���o�*&Y�ad�i���w�B�%r[�Z�}��4*~�T�V �w�;���mS`#�5��	�yn�A�_L���~�s��ى����p:��2Z�R�bur}$!�:��>�bm��7�a��tЅv�ӧ�G��ք�j;SAƂ5z���tΞ�Ba���	��K� V�'� ��p�4� �c�+�6�5o��C��L8}k��z����1;5��jPPd�*VIp��{���N���LI?yG��]߂�]W�T��{�;݀n������v`i��4[���P��c��`ؑ`ٺ�}J���4o�$㷨�V��D`�5΃�y%���L�S��C�TzgR|[Xhi�j�
k�2��݁�w%�P�U�?Y�q't+'۳C>W8���I���i.�� ��y�^/���AU`�:>�4��n*�h�c�rF��ն_��E"4��+��pi ��u1F�u����.�H�$Xbjd��{�������@�	���D�\��]�E6�hX���as���ZV��6��[�W�8��DqL~��ߋ����H����x�l& on��(��EBg"��h^�������mz5�VMZk���>��0u��
�G���	 dU|�d��$ـ���J�Ҳ,�D^�3���Y���>�؉?dw�{�pt��*2�I��I�b5��):�����WnT	�B�����=��J�J��MX̊�q����2�z6]�R��G�>m
��X�I�<SNG�H�Nx��[�;&�e?�*W�[�Y�]͎bD�=��j��xM�nF��3&�����,d�h�/�2����b�p�"Q�����f%���e�Q�-����gf�(��rIX���M�ƽ��CH܏���q�a��B����;G*{���Y{���9�!��[pf_�걢���%��|e|
����U誰�-�60���Z�T`@�GbˇO'ɮ� A?�pQ=X����SE���O���BMA�����?���S�.
@(ie���W��Y��y��)I���nJ�]Py�%��d�9z�j�8�xԚ�yД\���U�����?2�|����G�9�Jj\F�r/��5XIi^�e
���\�[Dg�keh?g�=!QT/�)�ȷ�	k%��LKu�@ ~�q�}�w����4&�V���j�Y�c _ N�B�'DAĨ��t?S1�/X<@>�-v�\��Y�s�i����<S�����^><5�"K�ڵ:�Z�Υ8�&�T
��w3�����)�K��Ւ�h���ל��\t�vO�p/����(<$��3�ԉG����w����_����ŗ��d3���I��Z�{��om�+��j�s41�TB8�-��+�Y�O���G暎����Ԅ���D�n�yZ��4��d��u`���U��:�t�v�\1��1s�V��K�eej�e���,��P��Tm��6wa�#��%5�bY���*��^�?H�£?!��.Kۂ�Rl{C.��8D[�k���!�c����d�06Hτ����ĸ)�%�7#$̧�P+C��"[�sF�Z���)��^�ϝ˝��"Y(�Vj��}��L7�A�2��n��p[�:��!��|�!d��궷����o8mq�UZ�8E����	X�/�YR�M�k����������%`L!��0��k������?�K|��$]�hf�6ȗ�1�"dvWr���R�L��K^䉃�^��#g
�(����Z�v�4��.��"+�ѹ�~�ѧ@J���6��,����
;0:`<���4ϒ@�Z;�m�kt��|z�"#y E��n\�����{[2�48�_�>g���}̓�?T����6��7����ζ39����,��H��V_���u'�/�o��
��H�>}���ў\�&����0��Vf˶���+�J�OV�'����"_�q��Et���J��Gs���4��/�]T�Т�R�Rp�u>s�5^!������!G��;YT��+�uza[$�4N#g%D����"��Q ñ���?	)�G�4��uN%��o�̾�h�?D��Z��i�B]��=��
��BY���݀��kyW�����@ =�a.	T���-U�������gd�qNW�ЅV��B���Ҹ�^������q��w��sk�V�AYM��2L,�����Eg��n�k��Na]�T�\X��p焜&��iQb��\t���Ãe1�t�hИ��Nk���	� �Z�c?N�*�0v�,j
6]'DS��<� 6G}���_pMl�:��Q�L�W<Nh0��Q�b?C`�j�Y��ԑ(E�� ����o{�[�Oj����r�~t���̊=~���mU��a�}k컵`����e렽�("�Z���v���*���]�Ί���FJ cA ἵ�9���~.]1f(�N���t�Ii���7�āa)�6a�_cV��滸���g�:��@S���Can	�X(ޯ5��'p�o�kr���L��[gg[#,�>�&�1���(z�f�P��t[ȯ�72��3����Х�O>C��~��y��1�kA��8#�f�s�GT{�x�G�Ҩu���`uf�
�#V�~�ss�?7�7Q�"��� T��ٛ�Q���� �|��W'�W�C��Q �C���)����1����2c�B��iZ�]��%���CE�'w�^��7>�����w��Q��5��{�b�=\�i3?����mD�����n��P�l�V%�xx��]��T��J�UM�c��mT��Ns3e����_�1�3i���y����hE���Ϧ���-������d���"�_���\���F6ݠ0���Vŗ���(-�n*�x-���r:�)&d��+��÷���J):7�W���!�V�)."��)`��!���S��>�7�C\����?���Ώ ���oqʥ���S"Šh���vz:�r9��:҅kٜ�r�������
��i�e�M
���n��s�
mE���T40��)w��Xo�	���9���D3�V�	7�*�ż��E��^5��w^@5 �q�@�l��XTet;Ǚ��p�(�j~�ĩ30o�93l'���п�lPR+TxM���H"kiRy���O�����UQ{)�N�R��$>kZ�@�0���7n5��X���V	A���t)-���2�:W��\yCӅ,L�������%��=����<2�
�����b�w�8�+�a�H�b���ʉ=��W�bF��~��7\}�n��2�-*���~X>I��������d�G3U��3n�B�B�7�3m�]MG�s�E���:V�JwRg��f��]�adD��1��ˏ��ߵ��͗�J>���zl�U��9791�1����-�Mq}�? ��ǖ��ka�RK������٠:��w�  pA�/ ,];^nM@ݕ�u�n}UV�H�^>o�M|�O�H��ü.�L�����j}��I�v�K�~$5=��=��3"�I�J��І�d�}筕p�+U���6*���q��&�v;�6��S��)c�R��z-�^AQ�#d���i���ɬ�(L�3��~e����,�Y�Ed��Yj���5������H�5���0<�!�i�c���*�wJۤ��
�
ߋdVI8�ں�~W����h��E��������Z;'ŔpxI4�kg������xc>3���Н�x:�U��$��A�7���x����G9U�k�!���!m!��2S :����+�J��]�:��8-1g����P�����d�)����)��!
�kd��F� ��Oi?��>A���C/�@hc�L���-�v@�R�#^��j(�3���d��@�r�����6~>Ա��c�b#��r806�X�@�攎!���Cfm�H T2�#m:�h�C����J;�7.]�V���D�sbm���5���|�	w$	�Ϥ��v�@�2�|w�!�:�=�Й�����q��l�f��9��n�[���k��G�q��م��^�kv�zV��LU6�q�(T�ds���is�-��;'�C[�3S!	�i1�=��֥��g�GCG�*.�Ŵ��7�-ʏ[{�*^_�V�+m��L�m@�H��9�7�2K��d�Y��[��>j�=��#�$���~����io����p���Y�����	`#�&� �ӪSɵ�j	����ا�>���E��g^�v�gj^X"���S� ��"�:�&�cm�#�����{�4�k?�ڪ�F���e,`Ҩ����O^̨��9�7A�ԕ� �lJ��t���hcQo��.���g��Gb声�)�Fl*p�Κ�Mp��l���jb_���g,��?ϔS$u}�?�)	Lu��dv��C|�1I�w��ID��r4��,�gF-��2H_�a~�qZp�~C`��@r�C	�H\x9;��mͷ�VY�@��bL<ѝ�v=�`ړ����M��0�6���4gc^u���z>��5iA�*�N4ٶ�;	Q�0�OO>Y�.��+
� ��� w�B���Y��-��ny�d����b�6K%N0�_'���I�ƣ�=��/�+,o �q
���&��Z��*o�%W���
�M�Cs��!Q�(P܈�N96��]��t{�O�E ���ۛ[O.��0���
@�c����ސ �]x{m7�q��WP�j|�)���?Y
<S����'���A��´�1(��_F�t?޳�=�HnJJ��>V����[�t�VIO��|/p���id �0�*�OA��ݺi�觧��@� II3�V��rh�/�_?M��~EhZ J175U7�t�L%%��`�g:ү�$��ѕl��V��!F�$���vG{V��Qr5�5��n�T�{>�k�ױ������?��Hn[G��y�4��e9��Č�ՉP��7�.s�/܈��b�R�J�ZX
������\���:y#Q�.*����36�m�W{1U�6��YoK����D��H#��iGv��~��?�T��!��w@n>�25[`��a!����)�O���}����X�UҖ��E`r���tH�\�Q�0�flKnSHР��<�h�4;\�.�q /fdp�)�	���:�J�S�9�t�6���w>>� H�١�#�I,�G��k����ݣ
���5�̿`�	��Q���܏C�D�wA<Ffs������j�y�ܻ�kCc���b@%yo��Fnz3�j���
��d$�*d�_?���	���=�q@��k�\�l�|d	$�rWҵI�U�����`��q�'��i���
|tʙ����r!w��D1�l��wz�a���f�^{l��D��yCg���(P�����B�T�B"��w�f1v���a�{xZW˒o���9��o��ZDZW�)Ҷo+�7����ð���*��0���]"���v��\p�|&��GzS���D"}[�ȴ&r}��!�C��Y��v+���x���H�°�mxE;��bwvB��
Rf�%�2������'�*ݺ������v0).�W��΢scd��9���!�-�(�������������,�MQ�<�0ȗ�(=i�,��EA¬i����!�y�Ĝ
��Iծ����]]X��S��4���ͅ�9S�YD��jȻɧm��#��xl`��
�/�z�I�`o!�T��ĭ�'�\��*դ�/ZD@�۲�{������.�|��2����+I�?�F�#����K���Ѭ9�i�{n�_�W������Y�:�BMЎ���PM䊜<�@th���/%�6����V�d`�G�c��d��h��x)[2FW6��w03ɨ����&��IY�����2�(_$��7u�<�m;"����S�H�p�.*��\�vk���Ii����U��u� �Qp�M��R=i�ƚ��Zn3'֨$���Ah�����r���c��>.�y��D$t*sC/�$��a��K�^�=)���[X�C�|�V\�4=&�Dj���H���у��^�v�#����y�C������CuI�XtEG��|![�P�!^q�m�Rbf �6��������6��2R-	x� ��3�J��u��hp(s�L�7Q���ј]}~�rA�H�"�������*��`BZ�?? ����B�[+�.�K�
L4���Q?05p���cy=���Q�5���̈́.�Q
�ע+jJ�1Yک��蕫�]�b��;��������(�������]a >�L8�Gµ{�gu�Ǵ�Ɣ�~^U��Umxv��`Zy!�4�j[m����#���� �5�쇺Y/>��]�����%�|�&#K�^P6e��BNt�<ͺ�aMo�out���E�ϐ�0W�ٜ~��4��$gr�2De%�����+;Pe*h�����#��LTΗ��$�%�c=r���%�F3'�6��1n�f���W�#ƁAU@-m�.�K���)�N���b��`� �>��_��u���F�	8I��9������Vm5@1}%�'����Ӫ���P1<j�p���˪!̫�_�GE��LJ0�6�ms����"fr*S�b�d .J�M�8pC9��1��s��b���=�!p1KVs=�,���!`�`}O6[�5�T���[4c^��2�L����H�E��o�����_l�8R���P���R��Z�^�L�:��@U�\N�GX�;"�m��m3�Ƈ���K�6X�>��ء�ly�>'���tg��qP�{�uU7�ʸm�J
㣖+����V.[��ɝ����M�V�=	���zM'A�1�5����+?#	�Jy�ڊi�[�<ǫ��`s�2e#@ ����&$�����{�Ԥ����b<^?�4����7�}I�q�h�e�p�!�e|M�!؃�M�W�c�Ԗ��J���{/�Jn�&���Җ�%���~q�����M��>�͓�� � �MhtǏCi�>�-X ��$�T�De=��#��
2m_r6꣕��&��?����s��4U���7q���N��yvـO�Ja�i|xl�s|�+65�n�VT�W��I�O�-:?r^�X�%��1v}����&wqFE	i���us�uT�,e��� �9��m�NB�ƭ�z�Vp4S��M�;(���x�Zod�|g�Pd��N����}���L��-�5�I�țȠV}����L�R#�3���5R���o���g��,�a��UF����(�JY�ڔ	����/�n��䗎E%bVs�5�d�^R��X�ݙ6�;#�}UU�V@��v���iCbC�'��N����[d%��1����c��F�S���l��4����{�J��y���],�Q���F��?����2.�Tv �!�����E��C-&�I
\u��i�»Z`��z�8ity,�ڳQW.I�W�5{���jul�b`��M!��g�ռQ�2>�QY'����<��e���}p���N�j4fʅwǁ��n�eN՝ΐ<�<G@����Cv����O@'p&W$w�O���]�<��>�����<���V�aV��*jV�h��3&�1p����������Y�(����a�z/ۤ;�QhZ����
���*�X4J��L������F��N���~��S��bX�S#��?8�����H�u���$�����_~����r嶳[[�_A�@G��_D�Ģ�<Ѥ���'U�:Ԕ?.Xz��z��L83��Zs1z{|�綕���>�a7��%ck�l�ϗ�ʾ�� ����;�pb�1ၛ�H��q�;������f�X����	�#ύ#�ndPt���"��D��i�y����9;Y��X\{�4��(}b4��"�E�T0V�_���b|�!U)�)�&.�"̺^o2]��QS����?+�U�ȝ�|�����w	d�{�Tۭ����R�X{��@k��"�x%���q�=�1��÷z���a\ҷ�D������� t��$s�q21�y9^]B꽸!d�"��%^}o�Ԍ�f	-/�Q4�y�M���v�*i%�SN���ݵ��H�	3}"5�a����0
n@|7���V��R�l�[	��x2 �mgL�
!O���-��_Z ��`]2�0����S�ɉB�x�Y�OtC�u�P-!��T�������}�S�����(�GCNY6t�ƻ�W�����}K�^�!��W@܅&,��0�$�
a{O����Z5b��e��o���o3�t���<[U`'�X�����| �Y-�=��L�R�Q���l8�E2��:f����"��C� MU5��7)/pQ-�D�Jh?�3;�X�~��@��/���6�*+J����){��pc�����Q�
$��r�fq!Sc������m�Q��o��6��R�dh#��8:v�: �~�:�œ��O���3jU�F��sWKʯi7|hj�w~ncߺ������R�'C|������L��Ó��k��I�E@�m���ӵ�1f�vQ���5��CE����DC�%���jvɦm�2KZ�sf~a&�UJ�3O$����o�D����o���ѽ�p�Ǿ.L_E1���P�?<�C)��3�yף]	������j�B�)�= l�8���?~j%Ɠx�v��궪���
z�8�I��^m�=0V�{w�G��zxJ�]|�N�Hš�a�a9�}���-�5S�:
Ţ��IG#;�60)�M_'��&��z���4��c��6�g�@;ߜܱ�[�o�R�3y���~R@�5\/�.��[�B1�[�W�<9>�Pz0W[�G�<&��y�g����{XK�Ml%K�p���H�6-�ߌY�s�!�X7�����K��@�"�䎠n3|����@"k?���II!�ߟsULE�ȓ���B?;ܓ���i>��5�)��GT�es�f����*�Z7�21ǘ��(Oe��zpN����
���伩�8h�&!}��Ըвc�Vؒ�Q�
�|5ж�2"r��ݶ��
 ��B'�d�U�i��y�Na7Yi
�2m4"�$AI�1�)�c<�4Q"�8_���͎��/=}=����������B��t�2+�&�#R�k��n|���-nyb��e�{�`i�ߪ��S��0˯_K#�႒U`/�*� ���4r�$_n=��7/)F��h,��;��ݡ�8���\�� /��������>!���."�CK9E�,ݡG�3�=O8"?�hӥؑf�VhO�>��]�p�62m\87��74�uB�#d�å�R���E�Q�k�;��� ƺ�+���d+U�+j����d�M�Hf�=���/���zM�[���*�j3�/��z�g)��o���Ԁ���V�	�Y�����������Z�;�5���ea9;3&9u0�/˗�ɗ^[{b�<�A}H~ӟ��/Ҍ{�\��gi��azFX`��m�dxb	���(�.<*��<>7^Й�x�3��S?���5�C�D~5��Y�7�3��ܪn�.KQj
���˶]:�n�K̫R�F��8w#���ڤ��76�%���5b�c�l��m����dZ�����:z�ދ���+o�j�T�"�O�*��o]�볲|K=��z��:)�|�H�{�=�KZc	!4\��8�5���'�g)���a�}<�ua���}��We�o��]�$g_��K���	������z�\X�p0ܲdv��שژ$��IBt���
����&f��js�\Ա�(ի����zN"�-U+
�E�@�m���Lc���`��Z�YG�5�'���ܐ-_�ɓ��f,�<����
Х0�Ip��]b<�����~�F�D{�L9z.-�BvX��dE��f�-Ј��^�	L��1�R@T�It�j4���(Zi��귘D $%�D��|v���N��´ѲMK���T7�!���5�B���OZF.S� e	�Wl� �G�X�f
�f�*M�]Bˁ%�?�X��^���!*E��v�^���wz� t�����
 �t�絛|�d"�2"�5��J!�x�Rr�^T�-KZ �r�Q��*ٰ���"��y��e[�,_b1�����bŧ<��m���M��6��޾p�[t:������7���QTH�#��Hm
)%�>�,�uӸщ�OZ��� �M�W�7�诞�'u�{���r���+K�����-�J���W�ѿ�S���|�.�vϼ����Y��b�.Č4I/-�t�_(�G��5�~�+��.��#3 *�&�hG=Y���'N�Z,�������HG��a�?��{��o���Z��$#�z<ٳ'����f���\�t��H�j���M�X�1AɬY{���R	�oBvB��!%Y�@ T+�/]�`��Z
�%7[��~�a_4�K3���� e��n�!��)Kj��|O��R!�������m���\�0�S�%���3$C�L��hԤ� ��l�Xt7lz�ǉ��_�tW?���1��� �xF�:5�Wy�O^&��l�/n�緾Cy����!z��!�R�C��E���0�x�@w�9��Ah����)l9�CJ� �eZ�L��'ӯy%�j5M�?��;�H� #`�m�Q���2+�ż����J��E�Ɯ9q!Z��9���v_D��h9�N�w���Ud���\t/��w+��d�K��I`���K��A7�Y�Q���m���������z" "������o����c��S�Yw���hS��;.�Xٙ�VaЪ�r@����ҫ|�c�T1��H�qi����ͼcFL�O��h�M���W�r�%2�g�zj�"o9���UbV����:c2e�Ep�iA3��#������� ���ǯV૾0�.<���yޅ�
��`���n��J#��:��{����3\W����=o5�\Qw<�*2��Ox(��6�݇�����uA�?���&D��E}�<�w�H�HG��H~�J�G�����Q	'�����^�<8g7��Y�8��l/J�D�]F/�H'Фos��Ix�0����+�)SUn^�wDk۔��%r)?Z6:��O�EOr�k�B&����ʂ1ü/<��c��r������l�G�%��pA!d��gك�>=�h��:D�ccߍ�ς�ƍ�X��XЭ������T�}�O�]����N���QW:�Ս�^E�`V�Z�� �!�e;i<Xl;� N�Nr6Օ ĝ:ɽ�۹�LT��R^d�h�M\�W��iY�o�Cx��͋�r^dЧU;� �d�3	�K��;9�[/��p�f�?�{��!�`��=oͿ�����5H�9<��y��S�|���% L�f���α�s���U�2I7&�7-
e&�!�J6�d�ڐ�!`^
�C8ypŐ��� ���� �[��2�бW1�"-�?�;��3����4g� I(b;�q��%4� (�K��o���!��tD/�T��%'�듂Yp�}�Ld�u
�t),L?�>f��'��y�eDF�4�a��z_'�,~�zܓ�R�f�� �������h��B)w9fL�'`L@�W7Du��/Ad�=�G��kHq^�����	�!�7��kuq�����Wf��;�{'j}����zn�S`��7s%������aW L��DD��YN�3J:u�E
t+�=&zl��~ վ��	��ǎ��,ncBc\�e&7��Q�`��#�Q�~�y��L�|Gv�KtO�j�0_��شOP�j�D���+Lݩϕ~�I4��$�a{ACL���5�.Z�)�6��뛃ψS��f�	:d"+b� ��H"q�D���{�kq|!<���]Ír��������vWC�79���8`�}v|��N��a��r&��l�F��g��CH+��g'��m�~�â��?��ѕ]��=����K�g��6�sB�fp��;�������'����t�3��:g9S�B��,�z���!�]��,��,M>���o:��D��8��/���$.��!���3�+򏅮UR�!�+E�л�S���_)�"�S�Ŧ�H�&1�#�46sSj��/g��f�C(�2j�?����)��b���B�5�3]_�+�3�J�*(i��TJ�Ѐ�-�����Xf�v��^�g3_)]��x�����Efܗ��'.���P�5��"v���H������P��^L]��Yж'��\�C"uߓ��	ny���Y�u��C�`P��RJ�n,~��I��%_G�>��jb5I��u�5���t+���;�݀%�d@�tR��xںb��������H
��>(�CfQ�I���X�.�����*��\k�n~F��B?g5�%_��2�����3��&��˫U�W�K�6�c��1�=X�7h���hF��F4_!�^�N$ژ�c7V�G�47SB��_��1A�TΞ�L��q�I�*��Ka��5vyM�{2��}�m0ˮm
�G
Sܬh��
�g���	�&(�n!�`�fm�ӯ�	�!�P�އ��2u�?��+=0��c/KJ�o~���2/�jE��X��qt�4��HXOQj����~ꭵ���?w
OO��9B61��~ b�f���S����R�̃���ku3񧘬~���W��*��힯��$S�D�� �Te�@� ]7�*!�U�}���
N�Ľ73Hϵi��!>J�}c�*��tq��{깢R��m���ӺY	���;��(��Z���{��R�8�n�C�����z�&�,R��mD������ل����L}D�:!s�}-�(���;�+�+6D�$/W����D�Z�7Lo�&���}y�:w��y�\�B8�kw��J���UѢ�"�/���Z5@��'\~k'�0";��飮'�L�H#����?l��J�5E$O�h;������Ϲ�ǮF�\=���D;�8��jsJE�[(Ћ�?�S'�ĉPx���Ti��J���.V��VcsZ|� �@���5�Z�m,�$+�u�����wM�gm�"|l�Sl���+�{�7�7&�
�u����-[�e2R��%�H���;�-FA����Y�}%�xk�Vq�d�WZ��"�����E�}�Ky��ny��oK;�S������o䆑�R0ktۆW��}h;�Eɇ�h{UJ��i���%'�%Ӏچ���k`�S�7��`�����=�ٯHǼE����ko��0�<qI��grͰ�7�&�s��U��]�0RӠ�W�(��6�K��X�R�fÜ�c�T+B�������!����\��_�J����pS��]���u�/s�]V��L���Y���`\�P�.[B_�#���-����Ժ�1_#��ԡ1�y�P6�{���+*L���"��t/���0��5��rRO�|�0a�, ��?mY���J�Aj�N���)�����	[�jSs��s�����\�0�2�$�W5�cv���Ѝ�8�Y����D/0^"M �F~����칂yDlֺ���� =� �_�X��!<�ý�^�_�h��Ҕx��	2��	f�{��v�a��4v���ֹj*�6�T��~���1�����/V^��_�@d̺,���p��}�9I�Q����]��I��P*���ȮG9�I2r.����i�AӅWí�;�9�ý�FXGs
gޝN����G�� �8V^E�Y8���q��;�nf J	����=�~�ugTU:E�A}�ތ|��$�h5���=������+�Px���,˺H���!���#�t� ��ȗa�%��0N�t�h��l�h�J�����^W��K���t}8�ф��=��`y�������úG8��A���%ĵ^��N��w7�6�q�!颶e�H?��pVB��G�d��	�㍌	e�	T���^�S}��z����A���Bϖ�w�l�6�k�a7ؗy��4����9�,Z��6��������G��x�j|Z'���i�^T����x�b���Aˑ'v�] �'"����UƣQ��.�P%��愃��j�_�FY� ��v��A+�'�Q?������@��x:��ķ��0��Y��*�w�g�mi��-��G��P�
��XXep�"�
b���zy��|R(�)�d|�5h�zѵµ��j�I!�ز�&C���O�a�B<f��˾�v�K���c�	o��5�(~��l�R��Cs[h��L1Ķ�Q@����٥��y�Ь��\�@F�\��q�=�V��n.iŦ5ȹH��������f#��Vu�*@r�?�_ӎ�u��X2��}�Xu�,4z�f�)��#��9�/3Ĝ��k,h�g��zT����ƙ<Խ�Q�v�.���3�3�8�Ne�'���o���s|Nl��%]x�BJ�BK�ȹ��A�%#훷J�> ح��ލfgC��{L��#>y�*|K�+����� ��L�l���t��7��qǈ_C��˫r��9�6^�a%�xu�B�(�� 4�v�d !դg�r���'�,�y�����1�ݰi��S���2�Q��7`z��az���i�`z1u���
\��F郂������l(4��R0���W ��8!,��?FJf�	���8�2rM�Gx���3�~�F ���:�v+^Ս�G�$w�U��(,�+C����P�8!mμ��t��n�:�o�7`��VwkM�Q�
�@�bh�Uh�vE�//_UlD�ص� ��{_�O��n��lD,���r�$���a����5����	���q%���ƟLRJ�5C3n�I�=7:�Q�^aN ���Aa�bx6���Tk�OiA�-�9xn�7��4h�Ĕ|����gZ�DpYK�d!'���Q`��S�)0��Zt0��S��X��<U<	��(���|^D��j�0 ���)��|���5Ե�'��2���~ 1��W@���ϟ�̡���a� ��/n�3ga�o�f��fބ=*����Җ��V��Fq�V�v@;Q�p�r�;$��:�~�r���N�r�3���0V�r8r����s$�rӟ��dkIb�\��I��:z8%ٱ���-9M�7Q�r��Ne�P�̺�lS����Gg��~�Z�q�$�6&֥ǚ�7���?�.�r���押���ӏ(�G�</2�km�S��n#ہ]~��>��[4�ʦy�6T�� �S�^�]�G�%���(��]1����qT�$���Wo�I#��٤�%P���b�{��v�x�o���G.#�`/��_|���7��Y)#F�<��d|�a���`l�8���z��Ta�N��斤�z۪��{�ڑCF��y��֠��a�&n�Z�-.gη��#c4�z:�j��օ�O���]��hf@6�iz���;bCܬ
�qX֋YC��v�%j�dh;�=���U�z�*W]���U�����֗�I����1)f��y��
�%�N7ȫ���&��ڵ!�Âͧ]�YR~�([c.�#��V�='�`�	<�ZlT�S7�7n���Z��r�QJ�`ӤyΎ�1|�
��L�?�6�꧞F̗��m�`�A��@a�SI�P��I�7��.��\,B�%'��L|c75��ͷ]Q\�[7IA��T���Qd��i���b�n��hl��F	4����P�խ�b2�H��g��9�c�HO��ϝh ������ͅ�:�l����Mw��W��Ti$ A���l�=��R}����0Qd�#am�G���{<�˷FZ7t���N
&��+k��SԐz֑���G�0u9��e*W���͊���M���)�[�]��q�� j	�"�N^$��˞y��[ݑ3���E��f'@P���d�,�g{��e�j���@眴���07&��n�s+)��h��zc��w����߈n�I��ZCD �[����� 05􍥖�(�kL�a�$j���,
�Ⅷ8(�����Jԧ��,��V�i�G�s��p�S��G���culeg��7p��V��ـW��4�f���ŝ�aFR\�W'2�lgh�s\����T>�[IH�E\��D�l^W\VL�����r4��E��ͨ��Gt�^W0ͰTI�S���iۋ����.w�bL��z#m:���6�:C�2�'V��r1"��XK�yU:W?AC=�T���*�oQ�������V���zMmMGȺ(��b�@���ߏ]+k�'}߮P=g2�Š��,�k�)\?�ޣ'������%݊%��0�[@5Z`Ɠr��Rq�uhZv+c���k��jq��t�K�Y_�d��!� \�ü��B����N�#�)OX;���ڊ�܀[,ӳ�����I�MM��Z?�<��;x�5�[~$z2w��;�@���M|D��<����g,� ���7�o	R�mt-�i�O���ic8BR�.�"��R?�:�����kW �*�*`�P�3�s�H�:����N\��(\��b�i�G�:'f��~TJ�zA������ �@@/�VE��W��sO��Uկ�gR8'��T��U����{�E�Ʉtpΐ*;?�:��t�vY�&�gj�̐���S]>�Q�xC}R)�z�yJ�0�#xnDڡ��{�u���GT�Ė�A����r$�G_H�ԞL�3���Od$Z#�ykD4��~�J��"BvJ�,r���D����[ɉg��
�=M��kh^�_�?�br�A|���/Q����=Im�T�&m��?�!Ϳ$�T������ɷ����2MJ>)�ov��@��?�W6�$7���h�v�{�Ɖ��V�l��^�T��� ���eek��<^>�]D�����Σ?�~?]=����7��Wd�Z�B������k|ci��~�@�P���|�w9+�pd<1٫�І(���'�������lN+Q�}g�+��Rb��k�B
��U�����ㄪ��8tXcM���
����W +#��*�\GhcZ���l���hFU�7 )��%��)�HM�������x)4�������z=-�&� �+�f6Ⱦ�)/�|ɳ.��{k^EV뫺�d�������bHߟt���̩�c��8�So����"RזK���a������$��[��yA����m������A3S���1pb~T?t�xh�d~�*�r/LcZ���5�T������DJ-�=��M���M����8�j��,ng7�!F�B!"��#�t7����,���2ս{�\����rs���q'��j�՞ �c`.LbۙOA	ٸ!��O��x�/(��6�F�"�&zL7����L8޽|���j�V�(��:����Q=J��r�m�=!�:��7�7L��DJ ���x�	�x�?C��B������*}�Ur�a�����q�E@��ԭ�����|�c��������	���H�Du�y���k�D�cٯ�Ap{c�:$E�lZ�9��sq����g�#g2s%�@��||���,�<%}�.��%�� h4B�;J�I�UK`+�k����Z�֩��6�w� ����Ihj.ݚ ������Ǔ�Z��2,wL!�.�5��G�>l�P��G��]�k�?%ɿ��H���/�d�ny�2��+8M�}k8���M�p�8�����'�� e^��N�r�K��VkK<� �<�(3��;�f�z�QOao�kb�Yt-T�
(4�&`� ��`k`��2f�ҕYV�bS�әC)�)��}����ե8�a����*E�kV�G��:r�oV�V��9��A����7�\��{`g��s@�[��(9��T�0��쟛_[}7YqB�+%ۮ����̷����i��*�0�abW㫝��˥L-��o?��zH�=�L��+��D�#48��m/h�� u���jr�M�%�N�u��{qL�a+��1�n����Yֻ�a,�_v�� ]����]��鍠mz� �s��ջfQa�FV�T����&%o O���Z��|=9r�q�`�Z�[��(Ѵ�N��J�z��x����WkvA:����<�7ԫ��Ơ����4;����l��i�w��5�WL��b�,f��p��D�%�ж9Yc���o)�Ow(�-_�l��㔿��{�ff�����?9�85H��/��-������$>���g[D�KX���/�����vi�bz����	�0���S���!;��U"��[�WУf>{q�`�&�T6��+�p&Nz���A��>^� ��+xu��D���}h�f�����R�k����y�a�
*�=a7�/T����c��Rǭb�*?5 F¯\�{��0��a:,�w��+a�Z������ J���wa��Z������b�� �",�ƳFeA/\񝁓+sm��_P�5-t6� �H����%��3l:]��ng%W�S�I�2�K?.��>t���M�O�"�3���k��H�U�c�:D��-��� �-sIp�&��p�z1�V�Yr�p������*����TĤ�� d�e��c�x�KM�����J�	�Z#H��̠�6&1c����΋����wQCI�+v:��P4�4d�¾h�r�9�Z��+�4�y�J�����Ye�1
�'%�;xa6���,�K��oR�+���ac'�f� ��@�z��d�����MG2�OWЖ�=tԊ������;�PA��H�v��ޞ���D�i}�\v���X��_��P�Va����{�UP(a�Z����� J"-��I��W��B9K�����s�� :���ߘ��˪6��g���MM]X�����,�����T�%!/}F��<�ߛd��{M#��j^��u��IJJ ��j�2U3{�t���[�7�K8�(?�D��^zk��x�0
�@O��SBڶ`�5�����;ϋ.�I��â���P��r1Ƽ����W�Q���.M]φ��)�"EtL�5U�z%<K�р��'捕H�90��ܠ�n���R[�$�Z����	�@i���v��1��A��?0ŵ�Q���5�xR�=C��$2�W8u $��|{n1�y�:���K*֔��b7H��9��w��tZG���!:�)��N�݈�Z��x#!�9��
�2�Bv	 ـ��X�o��h˯(�u����0�=W� #��h�Q�/��Z�7#�)4�;��q;�^�N>(�+��"�63��l(�>��Ο��8,�ؿ��B�Qi���<A�����
��\~�q�{-��f�?{}f�cS����D&���T#B\GC{{�8�pX�u����]�M�Ƞ����=��7�%�f�%jYx[�r�g��^#k�Ȓ�{|�Zm2��I�kݟb�"�h��H�Ġ?����������h�ʰ�؞g3`�#�!`�"�5�j�����s�:���p����ߠ�'�!{�7��AMV��4ꥃ��i�s� �䙐�S�բ`����	�g��C"�e���*�Xo��4@��,("���g`���&��e���e��W%� �s ��Co�&�/��b�8�;�|�zb�Ig�3>��|2�dț/��i�ؙ��q��O�De "ɖ�������)C{����KJ�t���k�
�_6���0�d�:�#-?�`�Ha�q��@��K�x�z𗃺��z��=��v=yuCN{�/ u�,��/�.~�)J���)k!������~�H1��Y��z}�{���7�Pq�㼌Fn�'7��%�j�^ۓ�H�~��|���.a���w�d�uf�!ip�	+��_��?:�v������A
���Fz�`�<��D���4_�BV�ha~z
�_>XQ&�SQ�P�+ +����=��5�m��ڢ����s����k)��h�y��>m��&J�T�KСk�9�u��AΞ��2�72'�ƈ�1�b�q�����$ֆ��;*g  C<��A�`���}�|�ӃįJ�=>x�a�ڴ)&��%5��'L2��E�E��w��U],��s�2��㰭�hYu�b��Dx���d�����ӿ6��Zj$�8D�Z��* 'v�]t��"ܱ�6n�1Ŷ{�G������3��S��?>B䱒	�� +��$5r'�_K�u�F�hq!W�2�*�W�KI�f���r(�+[���Q��&L��,�b�!��h�z!�I-�����ȏ֧&�?�.T7�$'D�f���w�4|�D�!
����P��3�7���j Y�?���ҷ���';5�BB��2J���wȒ�����~0��LJu��2]�@F܃9·O��6WPȀż�mv=ri��{� 02��$K�i�'�Lh�sj~��7潚�#g��KC���-��ḋ��Bț�l�ħ[�}�#��鹔�a+?Q��L�^�W�[O��3���|���TM2h�*�����x;j|��e���v�PU�=W�YS� |���#M�X�)��%��\����Ȓ�}���G���g��9~���4�`J����Cfo&i������42寙�F�}��� ��qw������keN����2��!#�e����j��Ů3��)�s[����NF׫���TEN�\�Ѥ�v52��\
�p~�M�>N&(&vX��e�O�3w2]���C�`<�W`�_����!�I_���,�#�¶*�k�EN8�ݚ��C����(��-|�id�/�J�^�^Y�ˡ�?|P�bb���i6� �Ēu�i&:-��ѿs#4���(�Ne���'�[^-����8��3���..�)u\6�P�aἏ5��n��b��"�ٛ6ÓY����� �Ҧ^���W�c��J�=9c9�PP��D	�!
�ê���'�2�5D�)+Ztsà��K-�e�	(�� a�ڊ���2�3ݹ'�zcXK�0k!��"N���۵Gn�W��{
�l�Tv�;n�˔���k����LVu�72�V�M�v�G�N:Ħ�2�� �;�pL{A�����ĜjM%p��F��av1!ofCiJFS�fܦ�6Gt%Qe�����c�*��g�9#��䐆w\RʊJ!x���J9(Sk2;�#$!ԥ����$+�E�]�6�r��y
�v��H'�vKc�1*lwp����s��T��б�����$z�;<SP�^�A[��|ȉ��[Y N�XlUl�����R��bL����:A�;s�7�^%�A�##=�`��V�O|gɳdRވ�b#u��ӈ^(^����8�A�$S���M���[[�bJI2�"��Wa�U`��g�<�n�ӐYy�c~
;k�z��*�	�f����/�S�
�"��E�`�	-�t��|S�~�%=M�_� ":�<x��p�������ceF2@�[���w��be���ɲ���P�M&q:>s�d�^�����%�l�О�u�Z����e %��[�筣 -ڲ;��tQ�Ҍ��SE�^�	#���Hm�I�d��X���R�`9�f��Le6'����#m-�ۯf��v�k���k��t�M&3N��^���m9��q��%�C��ܔ-��:�;����/�����LR�߮Y�:��:��B��5,�	�"�;���Ew��E����lB�N����gDAJ­"?�&�L-L2��iېX��b���b����g��ɕR됮1��Hnw��6�R�9�f$�n����[D8ʴ/#q��f�Y����L���֠����2xqr���sc�w�V3W�A�Oxړx��@b���b�|���r�ȶ����)�w�<���Y��f�'\���1�i�x{�%��D��-�K(w�%�_�#�2	O	x/
���Z4%T�B�g�8����$���#��	��^���=88�5�g)3m�LQ>�� -��!���MIRg[�D�p��߸�q�!�e�'�aVB-~I_{���o�̈́������G\��h����+X����^��zw?"#�ͷ1���O�`�Q/aE�c_t�50τ�_�&�*1��4f�ʏ�$"�!�
��P��j��R��[��c��h��O�Kr_6�W/T����<9�%]��s����;2��?E�p�o����lŨ��[���rB��@=��I�'�a(�' ���Ȣ����޹w%��8v��QmQ��N��+���ڈ]U�	r*�ߎ��݁v�!F���,�0��ۋ�"�A>ݿ�j}�9�$P�ϧ��(�t]�(A��ᰊX<�c���J�)��|��*]o�d�)���rV�ɂ�	��R�U�f�_P_���+Z� Z�﨓"�e��|stI6���;o���=�:��!$y�D5�B$�s:��h�Aì蛄�G�ؕVу���F�m�*\
�Aq��P�s���Ȇc�A_�n}���(m���I1K�#����a �{�����c�!�	E"��]�\�Jѓ�U*��b��}��%H�U�&R8���m�6�F�{���6��6���� ���-/���%6L�Iݗ�[*~�[�*�fa��-cdV��毟�F�é�o��~��D��Qx��"hn.qn�����d�5~���;J��\A$��yO�'�4�O�R���$D����m9#U�BB~9�\�H=mdu�Ll%���gӉ��ίa�����/�J�k���g`�WF�?��	^7��Dy�YZ��=�>���G��L�-λ�&7Y�g�D���X͓�|}Չ���OKc�{��t�ZO��WWO�_���'�2��m]��
i��Y��{K+��?�J���ar�!F/*+C�&�0��ʌ�Sj-Ezw�0{+@�N�\u��G�쫘Ā�g�\�0Z���_?��I6�_雫u֠�wA�H��t��	��㣇d��D���\�߅���q@�.
��gTˬX@�ʰ�pn2��(�����V.�*�|��r��L����캐�]O��K��-7�|�Ԛ�%��1�7�3���R/��A�{���P]��<�I�B}�F<5_�W��օ7o��GUK��EYn�
B��O{�:kC�N}�SN	���6�%-W�^��R�y� N�'	m!y-�����SFa��h��nc��TWJEr��֛r����˟'��� ��r�j�PW�-��IJC8�w�4�#��{�2������?��� �f�`��5�:�0����aoAc��ʈ���q��|xAp�%�N�C�{�dȺgK����)(�E�p�i��FE�@/o�%�d�wb�x31����S��"!��ɨJ5���_�y:2����TOT�b4���ꀛ4��3#�9R������Oy�d^��p�������nu=g��h<?g�J��Q�_+����p�Ę�Q�mj�	��*��LqI�+�I��c�+��%�̈<�g�9D�>�qf���dAZW�zg�����Cp�y��U����T<M�#���|�Jo��\r��F�W�$�Y�p+l��!�)n�����6�ؐ�0s�{���oz3�u��9��y7��B�f��zU���LR�������"���J䑫�e#x3fF���8�f#6���4���Go�q�Zcf^d�eOF#e �Y��U���u[_EX��F��\�e��a�
��FJu6��?����om
m��� ��}I�U��y�h����^�AKN!;8���/�i�s�%x*�QS�k�[a��,Tը���m�6H��m���� �(a�iU>_�w�7^��]|�3
H���n�S���B9��.����1M����b���Y�5����M_�&�F�;EK�6U�C�@.c�p��O�o��%�"в����+\@�*Q�L{1l� p���G��z�ք˭Ɣ�%/�5�D�>�L�����h�N|;�3���RvR����Y��W(����\]r`�h��ZF�(ï?�ݳ@si�j�ہE��J7���>]6�R�b`ҩ~�M�=���ff�S	��g�x�pe�(di5l�Li�������2�ZR"��Pl$z@�nMe�r)D��z�y.���4��:��h�m_`�be��m�5�d����&T&H�T^q�G��_̡ci�B�`e����K��:9��u��ओs �$�2�QH_������i�N����z/���\�/GZy��b�u����Q�Rw=�mZ?���Zv/Wi�������N�픠�8րY�� �!�A��Y^��0R��BB&A#H(�h�SV��d^�R���_6`CM�H��ȣT�y�wL�Fb/sF�R��U�pʿ&�� m+Pu�v;I������W��D�l��?RY�lc�8ip�I)��4�
�����!�>�v�o
��8����Q0A�&����7J;��s.m	g��x��Xe�/I��ӷ���@��b)z���l<߄yd�dx6Ӈ: 6�დ1s�&����qk�D��¸]���<�% ���ͬf[R��^���H/ft��#���d�b8��Fe����rؗL���Jޏ� |`�nj��A�����l��Q� 3�U2\�!��ڝuꖣ��nl쵑�8P&|���@�o�yv����h$M��{;�V՛��P��z%�,l�rL�I��� ٿ��� ��V�9�ԍ�X#������sgeR�\���V��N��)��*} �v�a?��M�G���T��n2����T|��u��)O�&���Fr@�A��;w�)jQ��(�HSE�<�Lp�4v�5�f{M	Z���Q�FhW���c�Z�v��bLGE�b䏎�C9�-��%ÃkT��e;�]��#4�c>�[���6���>$�y��}'�F����/�7i�p���L;�x��DW�4�ӡ%����l}��.�9dӊ�nۀ�u�6 Qy��z@u�Bv=�'����a�C��"X�^����d?j+�c�Y��$����ϑ�TE&�% 5�2�a2(���;`
D�e�O�u\�~�[��{fu}�nO�����F������(��JP��(Z.[]ҧ@���i���a�ۃL�t�F���?�\N�v��K���.D_��}F�e��6[�EL42z�(ԫ�=:�J~Y����Y���*���Ϫ�b��J����0P�{�o��o�x����p����}�k7_{}$�X��qls��W3��I�K0�E):�R%2@^Ԣ�]�`���L��ęj�T�����P~s~�Լ��י�=���8{Y�����	<`�|�L����0'z�"��j)�զ�X�o_Q2��l���oZ���&=zq��%O���o����w�W�}�N��v�y}+Гg����tZ6�s�g
�1��_w�e�z�*�^�������1%��@-t��m��:]��&�o�,��������[�L�l:,g�,�\���8Qޘ�)2Y��Ͼ��Q��a�QbH_F&�ޚ_��M�F��	s+�g���!m�7)�V2���b(�-TP��\���x<���I�#S��(ij�ݩKOٸ�}�}�ם��m+��+2�$�BZZ�w��x}���j.�<0�Pc�r�z�N5?�ʴBION���N;��g��DoF6��O�2֞�ό��"sD6hE��#��`�n��E'T�L�U�����pv1��V��&X~�he�q:D*)1/(�PS�5�y���^�@�"������H#��r���&N�~غ�A�s�����pB�v��Bأ(_i���%�l��K�-��j(�۷��I��*7@�t��^�j~��\O�[Pt@�nv�A���5�/~Z��}�؉x"Y��E�����l��/����7NA�0��} v_�_�n�R�>Ҫ`V����ޗ���u���7�6F��+M�y����D�^D�c��5����P9�(G<t��vp�g������$����r�yM�Fw��6�R�Lpսu|��L���j�>b��	����~g>��)��e� �`4w"�D<���&�?��<�������*2}$UCJ�)���)l����.w�X��Hei��/�Nl�X1�e�2>��)Ǵ�����W��N	k���q��6�	zL2�	�n-u��v�-�`�t-��J��B���c*:���@P�̲�^��gl�%m��:��]���$�o�Uo�	H.�ǴZ�ӠS<�%����i��5�},�`�-�J��<Ф1Q����*.ph�e۳��j
 �kKe������A�C���F+.X�v(�tQ1Ek%#X����{!Q�v�
�?���x0B���M�{�~�xpG� �,���u?��	�Mj%��B?�p3e �mB�۽ơ\����RA+��1����S@�q��w?�1���iÀ�喙I�y�T��8@ƾ��T����]��M�P#��E���p���u��@i�#�	U<����_s�RK�u6H��?5���|�����}��+�Tm��u{��w��ɻ��D�>�����q��n
l�\��x�e��D["��)x���R�L<���*�����uߟ|h"��=�:>[�S��������������V��0]�[_�r�ɏ_0wU�Sԩ�-�ԃ��m����Q|5:�tP�ȍ�x���~#ߑ��i1��4r6� v?���f�/`ȚO����Q�v�2��Q; ����ۛ�nNX�d}�e�^$NZ��l@kΊQ#�g�\�zP������6QDP������k��Y� NO��`���SZ�1���>���wF�	�.=�҃�(q�^�1�BH�W�w��b[ؿCHu���\�P{��t����h?
;³�sR��/�_��)���[��='3J����.���� DդP�ڰ.Q�kH;��_;�C�����*��!Q����@����@gv��e�˃�߻��D�%F��**gP�;���ǵ�7��b�[f�^^3F����0��WOO�������m��8oպq s�/�S�a=-�������r{�of�m�}S��cֶgWx�垧��|Šק��+8ǚ��T��Ϧ��MX@ï�ȭ_e{�\t�c��>��f���W�o���� _������}>RR���x7�cuf旮�L3��W>R#E6ű�2+HJD�^�b!���#�:�*A"7�������F��"�h)���B�&:s�+ù���a�)C���,0S�V�4*�����_2gj�x�< ]�-|��Ku�R���$��v��<��'7h9+��;0��z?�P��?��zm2!%�:Z=��4�T-Qnt�y��������T�n����<�r��[��|]��
���#{�$E!�1�\��-����֊��)^M���kj��FVt���^|�`��[z�(+�`��Rω�z� 0��pr��2r˰�j>���(ͰCp�#��	(���emH�r;�ʤF�u�&�u�n��X�Z��:*]�¾��F��8���n��ݵ�aў^)��ƭQ��Ȟ|�18���D��2Q<�k+��9�r�c#�ꋷ��`I��O(�ڊ���������Zk�J�نxL������x�9aH¢V"��/���-��dA�Ϡ��4�A����ha��S�����s2�m��7i����˟�ɛ�<�m۫�+��X�Ώ�TM2�`S�=2V�[�MFxhI���߉����o����`��Cͣ��;��Y(ٞL�fƺ��+�N�4w�K�Bq`�LDW����JC�����oD�?Yri�I*���#��8�ѹV�:�3�k��9�������v��!�$�(���N��-�n���ς�L"N[9�њ��`��H)�"z5Yw2TlT�4P�z��5���[�еi��Շy鱵9�H[���0?�M~���9�L󏃷�$ç��j�+�3�SاȲY�ki���+��-�B����41Nu�� �T���)�e�'��c�������*���>��W��$f���͚����+b���Us��D(��y�I)���uH/�n�F����ua����C��~M���w�D=3��4����v�+��F�ؗ�Un�ٹ�ήnM��4����j�fk�t���-m�G3�!H��i���}+}�:�dlM�`�ӫF����/�R�d�hw�J+�>$Ոk� m���I�B�0��J�B���e��W5cKn�������G���T��L�
J:��ґ�2'Qۙ�r��So�ה�`i\,�=�-l��P��rx���5
��"�%�[R���N�n�ѹc��jpM;�/���{���A�C5����3���^���X�/U k�W�Il�9OJ��=V֐Xd�!��	�4@�f��N?%�RB[�W��1�é3�h�*.�꞊K���}�k�b���g~,�dR����Yfe��g۔`�k`t�b�v��X�5���:��d1�TB�o��*���2���ەD�8�iú�����8�m���Gu�{W����v����%6�P��%���w5%�4:�v��!?��'ȴ���h�~����Ř=|��U����ź�{�{�B�����I훧�x�����pV|��R�P�������q&�V\���4&��D�x����y���r,�� ���!,.�񂉎���0j�Y�����Op ��٤j��h�q\��yh|�/ɬ����n�n��1~v�#��U�+3\��8�d�$ؠJ*X1R�p��!�{�?�V=vW��f�}�$����L�h�T�V�g4f}=���7���w������hdU����v~����]3F�!,!.�	�֯eg=�VR�*��?3�C���v��u�@VM��r�'u�q�&܂/�w-�͐o�T}	[�p�s�cJ>m�p�ߦp��5(4����B{��>�a��]��j`�e1@���Y��a�6pۚG��2�G,FC��Ǫ�&pu�E��gs��s��`.�\5tm�U�r�x)N�Q�?�:�]���؏�)���Q�$�°���3a��0?��UŘ(a����>�|�ʙ�6π�Y�PP�Wy�)w�Mw��2^g?l�<��n��Ų��$(:-դ&�jmC�-�FM�9�[Mo�#��Q�V}e[��l@?Y���<�v;R�j�&z���ۡ9�>��;t�T����tת�+ן)�e������\}?d���2X�jt�[�S��~1���o
�#�L�B��V��b�Y���#��j�F.�k���.DQ�א�9����n�|-F�ch����rZ�8F�a�����-3X�(�*�@�F��LvC�: =�4[9�Iݘ�v:;.��=�������8f����;��'?�c��<��?��Y�E��)�)J4Uu+� �kQ)芶u"��Y�D��Q�H���ջ�i���g8�!B�= '1�@C7������[)o����⮚s<���9�+�)0x}S}�W�yz����1���{�_؂����g)��8�H2=��:��H6p���v/@{>7�.w�� 0��B�jճ�B��g�ت�py�g��yӲMt-��˨�U~1= �T��N�f������ɳ�"zv/���5-��ç
9�p,xI��{Q�T� åٹ2=-�F =�z'�\kی}q7��Y�%O�2�J+]U�:4��"���fܒ�s߬pf?c��Wgb�g���dy�:ؕ�;7z���n�ܾ:��Y^���;de��C9+�ş���ۘ��)%���md�}�Uz~�^�+i�0�!I��x+>.�������Xp���fPq��>V�re���q{�g��R�C���ۭ���N3��o b7�~叢�q-��=sԂ6������c���(��F��/=@�h�9Sp���|9r�IF?]�Y'mt}P?:E�)���Q{���&�o��@<&�����E[ i���\�ۢ�~��Yɀ�v���:�_��aw-S*�DtQmo͹�d���	��X�
,�~���R�m.ud��T!!�5�VǄ ��(?�쁟,�`���aP�>�꿡� k)�"�T����bqgT�NR�ů��(ٔ��۶Qo���:�r@63és9�B�mS�Tf��Դ��+��<<0@%��{�`PL9��
vY��h�Et6�<����>6�M,-V#շ���lZ�k�V��ʿB�o��	"E$.�ƨ�Cl�kک�A����o��G�t7 �kR��L��#47�" u��V$k��^�,]J�=�>�vT;\��_�M2��l��ki�`^���ɠ�o�g�g��}�' צ^���}�X���:��}��:c�~}bKP�Ke�l���<
a�ňk��~��㸱������D^�9xZ&Ë�����a�Y� ��h�E�dt��f��; �J~׸�6u:Vұ�--,�_Բ����OZrJ(}%QԣA�E�)��.Pol�u�qM�)��A�4ܠ@d������B����� �Ƞ����}�M�Z��G�2��^�R�`_˿��D[�3�x�)<��g��1B����Y(w��^Y���S�C��z�-%+�O��r[������N���j�y��M��^H�خuz<�:�D|YWr���k���+��!����j�Y���b��5�c�T����6o[��9�_�����f���:��}�g���v����6?h����q[SrtC@�cQC6���W��n����d�WA����}�\� ;�Nm���8� �a��Z
�\;���{�)Ȋ%�NR��
tW,�Q,���E�.	���3dO����ß��ДVC�%�#�
���B��G[���*8R����J��]��2����M~x���ΣwV���+J|wfb���o�k^[�\Z��3I��a�E�ޡ	W�Ϥ�nn��9d<{4�G�Y$��/<A<�_mf�U�Z^w���N��fә���J��L{�䬅h�B�R�h���������B��D<�B?� �dj6{<�?��˳Em�l�-
�3����ByobՔ�M�:����7p ���׉T�:����-�qj������x`>�b=�=�Nom�u��{D}w��j �R)������ �\�/D�s��B�{y)�
;.�qF��
ϭ��'���>lA�A�cTa��\U�����u�h=B5G�Q�);��dw�`U�T:�I5*-2��~���-r亾AQ�Ɵ� �����WS0�{p��.����c��[�#"Y��xqN*�$%�������D�i�`f�<�թG�4_�����,�@���.EjNx�-2��{��^����v凐�P�e,�,�<4���LT��ޚC��Qe���O(�E���.*�!��隮��PBX�Q[؂�1�UZ2
��<@�B���|m����Z���cU�{�In�3��]vf��Fk8)5��nR8�a�r�p`Ѹ�r�������X֔�y��}0�ۗ_98�ni$��d���ؼa�R�&S�e1(���L��_������`��@5���ռA��k4���� ���f���Xo��3$�5�ι����::2���gV���,���m�&�J�=���
�&�9��0z�iu�ܖU{�c;0�@�uN�d���ny����/���g���3)���e�]�q��a��(Y�G�lt�C�ZpVx��(�}��� ə��1L�r�g�_��o`E�E4ސ �OG�?1����)?֗�*n�V�mz��(6�A�P�51�]��ؽN�ͷ�q�.:I���m��w�赁g���_���u�_����O�@�h?v���G�:���w���r�`�y}�C�ajSʣ���E�}��O�8q[�&���#��d~��g�W�$�VUT��ճr�.)̶Qe��P�������l�v�!Q����{�lE����6�o��f�b"����Z.����^4��r�T�X	�8��~��� ��yi�����k����|�kM�%��v(�E�:P��w-����h�c<��OF�`�&l{��A9h��!�g ��i�G,���t�'���J?ǼM�0�@k��2c�z/�-��c�%9�Kmɟ��+���R ��E��WD�ShqGt�3�W�(�H�@��vo�09��0@n��mm�����1�|��m&���/��Hz�2�����A8%�q���ο3�2�\�G4v��h���Me?e,���G�m_]m�� x�F�bUo\���n�������",�Ģ�`�4�Ϧ�)ʲ��.�%C��z��t�'qRQMB�|@Y#^8�7�X%Dɭ1�#�^��3#��g�+D�Xr�������wU�72c�W2���I�IҮ��D��S	l�w� q�f�W���G���cI�������̚BQn��1�C 6q�.>�G�6g�c�ۉ1�Hh��m_�0�ؾ"	��B��Gkt7�8ѥ66�:ːr6��M��Ӧ�h����$Z��;����t"��$�V���%:o~�*x���B��p�R�!���K�fED�.���T�����O�T�#�R��� -�f��#@rŖKP�J��V_���5��T�3Ii����4��'<�"��4s%�#6�Zp�%��\vc}�!�H�!�j�v�Q��t�e3�!���Q�kίq�w95���QᏂ��L�Ct�����@���;�뒿i�C��1�2t���WDV�D��n���e��5�B�Ĥ��pA|���F=:Q� i������w�0M]�/��lg%��
^-s���T(�R^~�����B�6�e��0��x8V����"h���zH���� ���z�!�Q��Eƞ�A�p��9�7)�9L���"���H�O���P�����Y$	�fb��6A���INęH��C�W� �=}���jǙy�
��3=�U����P-ӱv���z���?K�d=��nuYL�~�o �}Üm(;�!��J6
��X
�`�@DT�IT�.W'R��pVy�(4�9�F�=G�ק_�M�1ϫ{���1�m����@�b�1�b�n4:Y�Yڤ1��}HI�n��N���w:Zj�L��e �IW} ��溛�~k^x��y<�B(��g����b���ٞuK��]�c��V�C�M�T�V�ԡP�^Q]�����ڨ�q�bN�{���q2���3n"��u��-3!�
����[^&�E�w~�jk���5�{�6V=㞋)L'ʆ��&x׉�z�'�K���E��3���]۵*<��b�!�&�5�����`�Gʽ�
�hy�O���ѥVm����_�Z��P�7s�#<��j�����s��
��|�����M�%g���gk������LT���G���!����B]02}�wu:� ��	b��C�7J�a����L���<"�3��[�5�i�[IwRZS��� ս�h7��D�]P�'��dZ���v_�p�r]m��}�C��/�5\�/��M���h@�����h~������]�3��B>(̦��זt�^r����tjc?`��A�,H��|�%�$�|a��&J
�w�YK,? żCf�Z����;�aJ�# ��GתP*�{��'�:S�p}��]��٪ģPl��!j���@R|r��I����^%�ӂ���E�Y���_0�{v���E�L���X7�3g'������@7�,p���d����E׃�9i�&�ރȒq���x_�C�?0?[�~^�Ι�����Ѩ �[�CzFt�BD����_@��-A>m��i�>���B9)�+h�Y7���0|̛)��L�{G��[qYT�L�4���y�d�y�	��:������m�K�C�o�3�/[]#�z�-��NÒr��o�椼I��+�c��ۢ4�G%�OC2�X2qT��7x� D˾T������e�,,B����ϥlS�-��:?9��xB�&x@��[��r���#�Lٝv�]�ue�A"|i������)�X��$�V��nUv�W-�)i0zD|��b�>�;���z}(1?/�Jŗ剻�� ���,Ck5��L�Īe�>���7�΋2Ҹ�7p�g��-�����"-AU�����kd��s�a�?�||� ��U���q���ѹ����w\��<��<���\(��e-�j��]k@�^�6�f��'����y-��5aq���%髍/��K�8�:�7���(��|B|�毳��z]����P�eV�qCb�_U��U4�l͹7@1&'}Jv%�w��{��al[�_3���3���#rd�z�YkͶ��+S?�D+˗
ߴi������pH��퉙�a��@�n|���c�����P�(+W[��,��)�ː���!F�{��.��hj&�7���&sS���ڧ�����|�&����̅�%���W��^<z!�ȏ��_�&�O��33������'���p^x$~4��c'^�N�&^S�]\ha�D�9h�&�0|$4���VpK0)Ǐ��.�U��s�S+f:��l���1`��n�8�!M�~��\'�~�o{�U\s.y��{��kiT�xRĜ`�Mh��zwH�
&h�����T�Y��G��k�Tg�F�OG�G�  Sdm^:I����5Qd��f�c	Ҿ�-��>���3��p��ae�"�_ϋG�%_pp��k�WL`�Ƚ/r8���p��qQV��H+�݋�"�����	�9�_>G����������*�(J��m�OuO�Ro����ɔ�!�ȋ������y��̌��\BŌ����ʽ2kTr��10�<����&y�.�(��D�߬D��:�[1u�G������i�i9RY"ԆB����	d������|N4��8��ьu�6��,1�N��.'wy�����%G�;�~��;���m��G"�[ȁ��/Em�����0>V+�㌿����l;vx|�A�K|�J��n�ƌ�1K�-���=W q����e�8@�#T�t<0�;�OrM�:�(��J�p���6�=~��Fi��M�6�$MM���Ʋs�T!%�݇��#�-��b-�9`�N�+���Y;��|��<��{F(�q�(��:�n� ���Q9�p�J� �E��W��D��fb�^	ՍRk��
�n���I�l#��f+F�"���ʾ4��G*�JV���%c1P�U�Pj��UB����n��a���`U�]#��~o{�vRK��C 1���ĨbB7�1Y���� LC/��e�?\h�k���w�5
Lu���v�U�y�/D̭i f��Î���'^���p3��lf�>c'o��c��Эi�~�Sdf�d�8�]�a�RC�:]-,^�{�� K��P�=h!D��`���!�X�r]�:���%I�A��%Ímt��'��\d�8[>|�h�� �^����y�T:�)d���"S���SGl-�K��P����Zb|����zY�-ڲ�;O� hv��rg1������2l՘I]�(&�<�0	����Η� �� +y�.��QѮ<~��N�	��}�Z<�f�P�x��&�<yN�ǚ�^ez��`�rG�9��w������S8��Sc���m,A�@��}��[��n�`�Uz�.K�2����2�
A�iNZ��Ȕ�ښ;�j�W�V q���0-�a���]d@'���d7y��v��]{�#/)�>�'?���aA���MR�l������oɌ�Y�Q�}�gq��'�]n�:�b��`��8�i�0�t�( -&:2�����7&h2�Aɓ�0��J _!O�-�paJhbB��7}a�j����d>֑tx�F����� ���"�P����e��� L����pN�vo '��Y�j�����ʹq@���{W~�r��_o'�B2(r������*���3*���)@�uH�����9��M�e��J;j��D�E(�ބ����-Bv� $2�.��%��9	V�I��O.,��ЁJK�� ,)�����	����%%���~�ܗt�m��
�Z|?�Ĥ���I9��	_��0�,h8ﬢ�ִ�s��kʏ�B�Mq�]�hd3�:�&�Ln�7���+	]�3���E�����N�Ԏrk�̈́[$�zsz���se�
����s��d���bi�;3� .��&��a� ���8�3VI�(�sy����i�N��>��67�T��WBy��G�+r�f���V�TMR��[M��XX2?�U��p��@X�����o���^m�����-_��)�f���}8c����~u�0���=��\����q�z�,�76א�y#9�V��[���N�O���d4������FVeJ	K�`�`�JD$�a�܁���ʱ��W4�P�Q�9J���Q�W�$��C2 kJ��E���mvdWbF"1���j��bN�4ՙk�	����������(���v����ʥ��4B��&��i&�NƼ���4V���Z1�gr������(�P���u���8�[L)���k��qH�m��f�3ε�ڇ+@���<v�W�5��bj�#P�j��q��}
�ε'f�!b�N��l\�)'��k�t�(V4?��!���;�����Av���]k��R4˛��:����v��+X.��Z-�ES�a�!�լ0~^���a]��_����-O^p��	����� e��cM=��\4�I)��sh� �����6�QW����� ����".�������-����������=���&��� ��^�E��>+ݮ�َ�;��q���*��G%]�pjI��4��Q�W���1!O%?D�V&�{p�a���ˤ�y�W��&=(��-d � id%����"�*+W�0
4*%kGd�����E+�hܫ�Ȣ�O�3���ֻέ|�6�le��[��0(i�
M�Y�Z[ԌrZ�F�߲͔����bm��A@�`���S6�yT�V��7$�F"4vS�bw�8�|��]Yat�BZ��K��g�m+��U0@n7��z<�F��{U�\-�.�;��	�t�$EP�J^�$˂�<�����Q��u�h~�����Ga��+����~���Z�� {�%Y��
�z�H|�C��^Q����(�N���*!�Δ�e���x}�?��n���D�,�"��Wͮ#QgZ$��ÏNC�
Jΐ�n���I�?n�MW��� ?%��bwe��ƞ��sI�����fy��vsj�¨��$���
��u�����#T}K4nNyW7�B�z�(RȦ�Ņ6��ߧ�D~��C����mq�C�;j�bg$��)ķ��k	�}3��l�d����!�ق��9���'r��?�gM���u0�C-��?�}��VW��C9\���Z�j��Mn��'.��+�t	a�t"��MYJ�{ ���Z?������vR�3�J���y苁�{ly�u;�<x��י��8��3��}1`.����@��"4S�]$��� �cQ~UB�t��nu�&?��,t�0r������}����u�����0��t�17�6�?'���YtN�%�7��q�@�.�o�k�nذS��'Kݠ���b�0I�{ f��U&W�4t��fH�R�&���J�Xr�eGK�]����/|���7+���wr-Ξ�~S>zN�<Z�>ɍ�IT�z<5]����N��S�cL/pq"�����=���	�_�`D�H���dX;��A�q�%�	��_�3��w��C�I�v@���j���
e��7��?ڭi��`��F*Eߦ �fVϣ�5��~��41ȺB�_	��b��#��������H&-����>c� 4 �m�9[��̜��j=�z�E-�W�ꬬCU���XI�8[��Jc�aJ�0���&��L��׸H�=6�����#S���T�Do�
��p�%����Ie~244��g�\�6ܻK`lv�0�;b�6�����6�> UsS�g�Q�J�9=ޙ�M�"��5L�W1f�x�{��o��/�x��։JY���kv�9���g�O�\���$+/���H�ov�i�	P�l������vE�kofl�˼�u�F$1�H_�B��j���B"r�H־��� ��k�Dd�<2Ѫ�YG<9��AO�j�l�I�á'5�oo5�X�T�c�CB�-zq�T4�8��M �gCRa��
�I�:���Z�ϗ�Z�z�D��59�����j�"��f\����XY���O���� ��!>�&*��';{��+�ѵh��"/r��(�/��X��P�+:d��ݎ���� �t;<G�%v�Bn�N�"C���#�)�]�D��33��6V=]����KXi�x��2].>
m�ϾkH�S�*�fo��Nj���נ]JYd�X'Ma����ERG���VS�sފ��	dyRP�q�[}.�줡̤C���	�c5�ŷ�[ox��t�+�:�p?ryG�%wu[����T����k�.о�n>��lv�c!�E_�۱ k�0�X���mR��g<�C��L�W�fyK���ڌ-T�ި�p�q���$�E��G����p�Bt�[T2;�EH�_����\��_�O.�����k����v_�
A�p�^;��n��}v��p�	]=����0T*�3_~�@�����N� �²eP����d,l� ��m�� ��-\ ��y�N��+A�7��GY~�X�74mq����t�E�$P�S�/]��T���1J�5a�4꿄�4�N���hA5G�wB��2��$O7�S�po��U^*�!�� j�d���2�&,�����6g�M0�.Xg�s43�Z�ڤ��I_��l`D�q%x'O +����V�?�4���<�?��0uS����&P��5t�R��(���܈'��f��Q�m!hp%���p���l��[����2�&�V��Nz��@�H��)?�a���QѲ��6{��t|�
����� ���ÁTr���g�p�`�@v��	�mz�
$B�"1��=ItoGjb�G6�0(Y�-���G��ꤋ�ڥ�ͫZ���q�8��K?Q�$1$Lm]��z4���m�����G�%�����3Wf:~R�����U��$��]M��'�D钯Ȧ��J���s!����E��4H�_J# 6���z|�ڴ����8��ܤ]$�]/��S�\���T����%��_}r�*)���y���NuC�,{a�����>�L�����eR�z�q6�9F_7U��$o��<Pr�9���v :a�3�X�3��]Z���
�'B�Au��Ӿ����E
��b=�֎(ML��/��{�r2XW���E%4��-�JL���7�O��9T��S!W�ܻ=O�v�S��k���h��%� 7�x�W|���G4��j�J�r1/B�u��eQ֧�ɟ���E��ugؘ/��ꭳn�ϙl�Y՗��#�4z��f���-�ɋ��� 
����mYݷ,�d-`0�wY�K��'ni�I�~[���\I�b�2�ϴ������sȤw$�����@��f^�̇��dB�ש?�;�q�k���y� ?ظ�A?t6��3��վ3��B�ښ@u�����WP ���h!�����/��?Ru��TP�%�G��j�d�5�V|۷BI�4�N�I���쟆������N�� j���C�R5�W.I�ܸHp���*+�q��^7����b�U�V�h�L��U~��`��s;��`"@cIZ���*s��%�ǉ �(ؙwD��$鰻�+��jV�jV����H��"��E����IZU]pش`ߊ\�d:w�+��r����WKHfN(m
�;�;&�u�k �9�ZZٹ�ڒtA��m�V����ٍ�8�/)Cབྷ��_�~��F�PvW^�k�l��b���z~�;*��|z�����d"�@���a�,Ӌ�I"Ejd��U �O7�8V�Le����Q��n�l���b��,w11�����"���i ޕo�Z���0(L���+q���ߘ�}�8���Z�(/r��2�+IL��x����R�d�Ђ��賹����u��`�u�HU{t��1>�֜I�A]��]�{"�{��6;��h{������&&���8�����(� �Jˑ�����;�V�l|�k�����Ac0���S�~�|�Ơ���اTM�q@yC�{���W�ݺ	#���	�����v��80Vk�mO�a��3�w�u O�3wȒ@�X�~�yX�;��C�G����c�K��e��+=�Uw��"5z�������Է4�=��dy� �&��J��4$d[��I��IC��x{��MY'���-�qYB't
W�y��R�zh��� [��9�l~!`%o`��7���� ��{	w�_��GZ̍�#��:�=��j��3��<;��U!�7�Kdl��i��ac�A�ZF�)�����fx?
9��f�,#ĭ_Ή��*K��6K������vK�̰n���֗�eQ��l�-�U"W�ci�)"�>������w.��{����O���+M������T��� @VT�阐n���4�(c�D�
Ҡ�]��R�.�\)|l�)���}�Y\([�6�E?��F�8���H�XA�!��Qڱ=$�EC�0�I�.�z��1&(5�(���1��T~��Ց6�/�Ki����O�ˏ���(��p�}ͯC�ɥ�����W�$)'��;Zh4Vu?���v����OC�0r��Mޡ�V��;�F�QDo����p#APqBGR�kfFjQ����"��3خ��C�4�+i�p�r���O�v܀�D,u ���6�Vb��p��[�Т�Bk�u�ֻ�1k�o�RĪh�K@�*�~ Q��M�Pmʞ�"�&�W�%he|wf8`��F��Z��	$a�����llD�-�@-�����\�5Kt$���Ps`��R�JX�g�[Pڍ��>�ѪE�v擥�D�V��s�g�a�	�nu���<��n�#�����.Ɵfd.!��4Q���bv]���U���R�dEE���V���y�B�Ze6�98�g&�H���MF<	���,ܢ�|k�9�Z�_�ʊ�٤f���\�Q:����۾�"{��v�t�@@�ZZ;���s@3�%�j5f�C�b/�PWW�~v�T����H��]II� ���wA�Iƺ����0��.�4���E�KtY��a+�K����d_�L���C����=ѕ�iW��9׳�$��QD�R� f6�����u��/�-O<�as��.�?�|o�-�V$E��\��Mq:��m��"nA	=�Lfm�m0@x� m�]���� �b�}؟Fc'`^���p/>�V�7:�ʛA2�9}��W��7�������͞��:{�C����l?�gj]�t&�P-Y �������Rg�kB)��Ls��w�o���)'��R%~V̲���g�;ج�	�o���6@�x�G�lC�o���L)���M�	��2������Y�	���]�ev�(��i��!�3��CD��K �F���8z�\� ��y&�ʩ@@�����س*J�$ӃڽN�b���#�FK���(��Htڶ�B]��y�����)	��)FJ���#P	�	>��K�*=����z��kh�O^f_�?	���� ��}ȋͯ:K�US4F���U��<F��h��dc�ԭ�y�B7oN�S�9��T��d�ݘ|)fx�:����\��lA�9`!	ѕW�5�O�
��Dy_q���}y���� 0��T��>��KU�nAY��nC�-�Z&�A����H)�ت�s	~3f��v�;V��V�'"��Ĺ����):��V�0�@�CW�Fɢ����>ٻ��MV;L$�B�>yFZ^Č}_Vи��15�quQς������_�_:ݕ����@QԹ��Z��7��|�&0{.��dE�}�˂G'y��^��vl����'T�8���<����o.JU$}�t�`{�'th�)�d�'n��FW�ٗ;~_ɥb?�sH]�5�x#�UV��J�k)����MR*�H�\���r�����p�P���ʌt=�h��FA
���8��Kv�E}Kz��f���3��}�w��Y}��/!��[��r�[�&����d�(c� �cx��!�;��f��9ʤF�q�0C�pkz?�EfJ�\�l��rVJ?U�s��
^�\Q�y�'ߖvC����u<^�j��a���A�̣:��)�[NX����������/��������E�O<�3�;g���2+�v�셼��ͫ�x��	��$L2߅��e"�U����i���kB���ϣE��<*���?|��b%�!o��9D4�x��������r�Y-ݪ�է_���'�NPc���>$uT������a�S��BghZc��bRI�X4�v6N�<0t��W�k��}t ���Am��S�ǀ5�s�����:��A�e}v�|��GXe8¼�w�@��k�[�Lv��v$�e}0c�Z�#/qG7$E;����u'�V����Pe+U��	J�`�k��R2Q�����{COࡋ\�Y<�&C��d8��t-<�	�'��JjD��Q B#��'vJ���a9\楙.x�<B��ф̽��ϨWd��X����a�G�q�2i:��F4T�����[C�)]�ٞ�Gr����o @��0����Sc=��� �N��*#���s��鋟��+A)>x,��'��2�zHQ��/��[�*e�ڈL&M���GC�Z}^V��4߰�R9ͷQ}�u�h�HZ�p�k�o�������G׳!a�}�H�_O?�q !��+nI�u\if���OTɻ�G&��`�^�S`)1�����z�I��A�)�7�WZ�j�R �y���Ќ�n燷�N%*��@,>,�z~�\P{���QO����X��J��|@o�=n�g�F_Bvre�|��c�"�y5XoT���-��;`����n_yDوlA��WD�U3݆�C���gT�L�Y}����Ց�$��]���cZ)v�Ɍ8����K٨���qɢJ�;j7��qMh���"�nk�ԑ�&:�x����~��pE�c_��`���_e����Y5��Ij�:hm�WY~ͤXT]l�*�Jq`��U
�w��D���d6A*-⇇��o-?%�-͘]�!�,u�w0W�"�	�@Ϳ�h��TA�>�\s77v�Z����������&t�C6�D�d�)32��I���/�qE�0E�y�AA�d��%����H�;�[��V�Z�	���,	�����X�b9�]Y��{�Z�����]~����?�}4޸_�	�-�����f%��Ï;a���.,4UX*Ռ˲� Y!	�RE-ң,!#g*�wC"�=���5g���䲺��1?b�a��o��c��?�g�9��; '�B^��ȽX��v���4��)���������BA���b����<3QH�|��~=�:�IV%Ai�E��Gn�T���/�ױ���v;#v9�%6��|��y�%,�E[��E��>�Sm=����tv�h��$Xf@ސ��7Ko�	a�B��e�:@ c�TP���}���je�4mv�L��d�Nj�+)C*�����L��#��G�03�N�}@�t�5��~���&J�wPr#1��g��]�0Ix��x�������t�ש[���)���־�An��fz�|h�*(^��ѝm�ts�j*q��3W8�N}}5��o"�#����(S���x�	X��߳:�b�ruUd�r������7#^lf�v�h>�E��GfKi,��;���8n����3�Fb�.��#�ڧ���=�3�_��SrEwH��վ�p=�D���QUFS�"L[p��U��Q����HNb�)؁) ��SC�7ƌ��g�K{�W4��5"	|��ZxR��R�Xà�&�VzA�Z��	��?Y���9��c��c�ѢYѴ��IuK�ȇS~]e"�=���
_C@]Ί�H՜sv�gԆ���T�U�M��jM�ӕ�XV��ZP�G��Q���XH��D�]W���j�����/\�%7�Ƭ���]����U��l[aJ���,�_K$�|J� ��!����<N��w���e�:�D[�H-|o�ֱ�I.tւ��������������+��o�i�����!�����{�#�q�.�k�Z�3:�6{��$�g��6; �Օᮝ�8��C;��1�x�� d�&w=s�����L����e2ɻClM��+��\�G�5I����Ʃ0�H�ڣ�^Ѻ���M��05�f�f�AC�T�� �w�A"Mp8>%>P�KkT�3�ձ�m 7�sdcx)y�i���Q�?o���$(���W.E�Q�xl�Ǖand�q�|�e��Oc�*�\�I��P
;\M!	׺t�y��ެ�qj�D�8���{��}8;��6?oqԐ��=�	�WZ<K�%����4��T���|pϞ[����w	m�<��L�l�߲K���~��v_�\���{��۪fB~��L��L�ӻ��P����v�'�\�Rt����Nx!zN��-�ۭ��߶����P @�� ]��w�T�Rz%�hӤ��sn�1���}.ް|ݩ�hJ�/	B/Nf&h�aӅ�y������;bO�Y��
DɓN6�*<l��g����@�ڴu����i���Oʪ/n��+��s4���hݧ���5�Y�kT9�d�b��6ot�L#��?�bw��&�� �f���������j뷠�`���6��ʓ�ɸfØ����AiM���|D7�^P2���c��K�er)�4�^YH��l�n��0vn��������a���@��S�h�&of�j�E�юP>¾Y�Rk!����> ��T����Kn��x*��}�ﻊ�~C�Oms/@0��xU��K<�0Xj1��w0�q^��n9����A�l����݊�b"m��o����r&��29������<c���H�3�Td,��3ͣ�F,�ʵ:�\:8������ �d�9�b���+��v��@� }+L�q�(�^�W��|��9|�P�Xh�풩E��"D�l��~�X���d�߰���R�a��SW@�m�؅n!��,98�o�_��IQudl����Tw�]X�F�
��w�Z���ek�@5����gk� Ӥe���j�����pq��"Q$K�����/M�g��1n4�>���ȹ͓�)us��Kݧ�c���tiT��U��5f��	��|������f�/�#uR�<>FH��bvlfr�E��X<k��NW�����T�BU=Qa�h�y�,2e���-�P�`Ǯ@�L>x���+uź����܁ξ@}� Rj+s��p�Ւي��1���Z�7%���S�DVS5
�t�����	���ໄ�N ��rT~�~1j6�-r���X�~KX���
�iu�2��q.�Zv���m��Q�fwz���G�m!��Ɖ`��Ť�lo'����מ�I{�f�"`��5�FE�k�F��K��Ct�+�	y��F�?��e��%��Ke���\��l0��>�-ɨ��ɟ��Q.�X'� ����	¯T.O!I��6M�#��*�9��o��k���%�%?u�PtL�y�A/{�h���5;Ӝz�L֗f >נI�49�5�'�����)�/z�^*Sݲ��2�p�U��)<=68�L���hv��,��Q�!U�*��J�E��
p����݉z'|*�R���c�j%��yTy��߄�st��t���yMc|�mk��))��)�0��4��Bh��>ٙ�A8�YgGo\�&�F�rx�H������:��C!�cM��p���*���m�.�r՚Ƣ�I=U]Aʉ�~	$�&���ni���	�)�����K���&���ozW��1��Q��m
�2ԝQe�Qֳ^"�'��LS���;�Im+V9p�CՅ;�rU��D(�a�T鋴ؔ�E��-S��Ԃ��h��cM���s��f�j�'��w[�W�q{ŭL�0l��� "�5�0�9�z-�ӸeI��;|�n���	�y�
�ۤK:p,�#�E��ԋU�jZ�Î�+y֨�h:hu7��Oqt��/�`��������o��|$��nn��{3�)C������Lߒd�P�^�ۈ1����:��u����c�XRӀ2u����? DG�~}����h��g���o�_�EV��آ�J�����J[��N[M���P��~v��}9ܨ�����ݫo� p��꾖Sý�u�m���U�ǚJ�����s}�.]�w�BPa��`�-�e�LkI"�ޚ���.q��V��j�u=y1�N�ֹ��̍�ZbXR�E�j�&;�v� ��ǿ/��>�)ib@j�֎[	�E"��"a���~ ��M�A�q�F�bu�jT~���x�ʟv|��U�pX�@*)7�]�/X�'��b���>v��(j*����)< ��NF��c�o�~'�,�I�ցT�:�%�� �j�k��+�C�ƚ)㻁�I��<#�� �b��Mm�0l�-�T�� Rٶ�kd�##���[=�*s��0nG�>�\0�!��-�X�z�>G��]N:��lSO�_r"��s�����~�s�r�k��^./����)2ɉ���f�����\�0y[\�M@?kf��y^�<wZ�0���4�i� �v`���1E�A��M���`g����֪,i������/�<�,dKx��C�}�wi�@��k�,�N�j��.@�*:�S����<��X+j�ɲ����e��o�F
�����[F��>|�MY��&~�TЂ`0�ْ��r�����Kt��XD���޶��.ѡ0=�����e�R�u�lP<��f�;8�Wؙ�ۣz����r=>z"��1!�<uu��|�t�c�9:�����:�V�Co�!����j�&��S���DLJe�K	M����#�V��l�0�ؐZK@ۙ��(�#MH�s�=�eM�t��H
�#�J�^-��>���<�_<���U�A�͖����IW{�s�.���-}Y-_q5�mHh5�g����(���"B����m�-ٓ8�*7%���Ք���$-�/$s:�)�_�棊,%�rE���)F�&bl�|�.6@?1��~�H��Ī΃�1���0��6�Q��A�9<��b���Q�u@K��k�m���{�HÉ��~���g�5P���7h���ҿ�U1�f&���O?ц��M�7W��t��[��s���T��`��%W���Wv&�X�<���cI>^#�O	��0�GZA������v�e����e*��D�����,�����SĪ����W���l7���lC	�Jk�I�S���t�i��uTԴd������fS�R�@�@.Y���>��a����g�>˝���$����P�mFhIg�W�	�?���W�� ������87��rK�i~�	P�� ���-� m�Ώ:�Crٮ����@�^��UZ�{�cYޮ�5��u��V~V���W�fZ��X���C��i�t�ޠ=6-l�\���\��ʹ��KEE~�	r��+H�E��¸��� ��`�	�f���&?-�N���67����%�gɸ.T&Qd�՝�]��,������s��q���z��lq'7�].cL+N��ʟ�c'͛��{յ�`�܃
�Ҽ|U�]zAUo�ä�JD]��A?�DcΆ�S���5L!�^,�b�z]����krʥr,��l�,f�(�)?�f��Ʃۋi����5��%l֌��(���V���
n!��L�F7�Ǻ�P�ڀ�	���#?/��&��1���a�׳3)�S�{��
�Oby͍t��Պ\�Hi	���9�Td#x�lE�,��
���-�[N��kC���vH��&7 �}|f(?Q|��X����Hغ� �R�;|�� ����l(F�r��$t]����H9�҈߀���_X�|��e뀋�J-w�t�nq��"t3�q�)�"�՛K��&�n+��r�=�O��C�%yVW
�34��ud(�*�
E�0�0���v�����MD��c9����jDKg�a��1�+=� K��)�+L �>�w#[sIϴ��$�^�Kw�K��Df}���/�����Z�#�����.�DP斋�*���h���7m��iy�VLU��j��7H4#R���3p,p�j��	���&Z�_���́�'��Y�'Hԍ4a�5���?%gC�fvO��dD��R���J�iܦ@|�!϶����-�0�����=W��vL�7�DG�	1Q���5���lī�T��s fũ�1��Pf�N�0�\��1�Ihω鲴��{�Bj�G|u"¼]ڠ�&1�k�菤��l��7F	���hVwv��倧Z����J��B�Ó���/��}���J[i@v��b٧��摁�i�Ug���˫����|�3�`�
c�}����F {�
~;�3����ao��(��:�x�~�&U��
���Vq��J��\���7q�� g  �������~�L��bt9��T�tK��hqZ�1l���?Zh����������[ �	��/�C�����8x�6!]�"���Yac}�}�ϥ�xhMx8Y�������J�Ϭ�>�L���I<�hoǘ,+�,e7�M�XfMS��w�&߄��UOD���:�%cC��"�8	st`�gjL*/��Pqs��u=Q/����q��̯*%�S8�ś�	G��O?�9��X���i˃P�>���:8�k����V�f[!��BR�0��rC��XP��-��B��h
H,�� ܌�MT�x�� �䲨�A�����ؚ�z՞��x֐�1�R;���������fJ�A�՚c��lE �?C4��c[*�2��g�_�K�Avl�S�U��h8�H���������G'K��-?ҳ[@?�r�H���ݓ7�F�3t�L/mQ#��hy�c�e���l}�It@8܇�m=E�Pj5<�+�\������������O�h
4YC�5��֜4o_�B�ce�n�Ѥʕ��:ǩ5q��V6�i*J���ݼ�ȷ���Y8��?��8\�2�:xMAfz�Z�@��'��vրؚ�1^�h-y��-�`k����DR�����g�η՜�欻�k
��

�3�S��y�~֦��#K��NM�ܙZa|�,X$N��Q�k���J�CTIi­yt�S�֘���/e��^l�7�t�r�-ɏ���eTh�Yi���3q�s��6�z���I9�g��V`�~����E�yc�Dƣ�ԟ�f=@Q��z� H����M�sp�p��E"Ҍ*�Th���^�"-�=�j�lC������/j4�2a��%Q������~#���A��0���\����&BНË{NmX�cB�$��~��
���8����t	o��̔�.p|�Ì��O��?��.N x�C��
����BWG�W��U+t�L��y� J�r����,Ms�h@y���AN[�)e��)��=入+Zҟnq�ɏ�������[o������е��3K�}o�
��h �2H?�2ƕe����F�o=��د�:w��c�EJ������thhYˬ\h�5�-tyH/�J%wAM�e*��ѽ�����}Tdsp>�w�[��ίB��������L=�c��\k�j�<[?�q��B���(�q֠L�
n@� BC��:H�F�v��:(IԟSy$Ԝ((l���ѬZ�7H��.�Ɍ�<�`���l�̵�钾�.qG3bW��%:�T��{><��/��f��#��Z�'�.�j�7L�J��R��*�
����4�Tj��yd��.������;��S��]��<�0�\_4ȩ��S�FCd<�l�um��ҏ�'�D���f/�C �Bl>`��N�V6�\��/��1�~]���^��?=C{��c\��Y@lK���o,�R�.��wi�
Ԭ|����r��G9?w+��,F:�\��ϡ��q�] q2���QD�u*��dW��[bg�U�;z��h/&��JO[�V���Q��"��H5,���k>�Î6�.P)��HJf	��*�}�ϙ|NCe����Z��	&��$�ܑB�D~�g�f�I�+K"�-�N#�uV���a���* �t�� �p�gj��n5R}��;Eq�� #��2�;`Q&�����p�� �SPV<c=���faA�]��!O�F��#�����B�c��ϫ|�6��W��+b#��poU�_;����Bby�0��J�ȶL۸N�����`�mcoDY����Sm�?�a=$�����Q[�����c=K�ˉ���q>N)�Ю��>�^z�H���N��H��V��ה�dV<�cI�P0����ף��'�8��knF4W{�	ͼ���~���K��ALgZ,�=J����B ���7qD��zP�UÃ!N$����f�W[��~��fk�;|�]���n�,��r3�>�=a͢Ș��$]����4Q�/痊`�}B9kp,a��C�?���oYu����o����rj{eh��T��`��P���Ț򻩬���R��l-��3�T�����b����>���h㰂�z �e�܁s��y�$����I�?��l�
�m�򱀀�]g��,0<!���W�@,�*�Ƅ���ð���T59�s��K���������j3�?>�'���BX!�D��]�&�1�q�]��3�ZB�)/��n<��ol�����s3�+��˲�h�wK�d�C/��eT��c�QI9sh@OH������k	�BK*m��GT��C*R��;&H��-˹
��41_��.�4�U��H���a?O�}1l)\Q���K���e�����K�M#t_�N�w��@�{����tĽ��8K��#!����?n(mUCo���[D��5/{�1�i�T�9C�I6�Ѐ�=} I�.��> �D8���ˣ#r�o�������f�.\�[1�.��( �ߝ6h3w�Cs��̍~%�� o��A�g/���艣8���p-p1Ma��W��j���#���� �u���eׅcK
�`��j�3�n�:�/��kԫ�����/�%������lűQ��#$��u�:��kYx�g%$���KwT�_4>i���[R�P���`���VԊ�*q��j�B���L�@?��k	N/�Q��ݐ��[�Dfp��]�a�Z��z��{e!����e3�M�do���bUچ�\��s�p�G���`��O��!�{��~?�� ��!@���J�^�Y}��9:�RUIK���ﴂ+�� !�z;��Ҩ�J=���@wP"�3��hR(���8���^c8e=yB��!ZW��ҶD(PUp`5�f
�ӢF!�>k�hX�E��s�n��LS��\��_!�G�li�>���| ��Α�#��y����	~�-�<n]ڨ�B��3��X�/9[�����M�Z{�|�.�	�7�."���P��Z)eOfCK���� ���8v�O�l����^��9�4EG�kx�F�fO���+�|%�6��Vwf���Y�f�T�.Ȟ2�%�7&�{Y����3c����+��K�{�����e�ܢU�����l�-E����_&o[=|��g�L�Ȯ��H��7Q�
|/ЪXG�8�]ԗ;����Iގ:��ؑ�+˼��O������8��˽*�����G��%�����6�)��@��*��0���Lp���r�paiz�h�n?e//kb0OA��u?B�φg��fP�/�\��s���~I��3�bꖨ�����j�d"o;>r�����C�������m�a��c^����2O�~�;�L��y���M��]BDl�q/��):
^�Aʽ�X�U��� hE�ɀ�i�*X�.���wĢ��Y��Ц����0m��":��*�`��|�|�h5:�~�(�oMO�D�㢶�ߐx؛�� "5u�\/5qЬr�2���{p��ڮ��L�֟W�3��Y���y�����ƻ��I������Cg�2ge�ةNb�V )pԚ��S�U<�����>�-����_��������� ��q���
e���If���|��	�
�-�vl����'��|�p$��YߖAB���U�i��~��Z�9�9�g1�+�Q<�u/G\��?����B�����N�%��c���↯�Ldѹ�jQ25���B���\��a ��S��� ;����"��Q��$>�L��{¾BV#ݦ��|�Q*c�e
8��!Зx���~��a�曌���KA�.�z	K���=�9�N��e"�� ?���ܸ��L�~��p6y��.#MY"��9�z����Y���l�
���(��8�����GlE�-p�zIk̪��d�;*�UFA��Zp:��1��q�s��*/��}ͪ���%�Cp.-�^8�Qn�7��l�b;8�v�Kic,1�!��� ފW�"\�~��Z�#;5yC?� M���b[�֤M�XH`�3}\I��Ɯ�{��GW�T�x�7$�P�.lmuH�O�"��q�*�o���%��]�MEY�����.HJtN`o�N _����� ����g��:7�S�׷7<#+/�V02�{s��S�:���Î���n���U��̘P�#Ξl��G���8�
�yq��Tq!v�t�<3���Wׅ�I�eZ<2���t�[�o,�v�s��0�1e<��b�ܡ)j���˺�3� �P!���h�V ��߹�:��8��b�k��(��c��Cѣ+J������0�t�w(ђ�lc%h����CқD����w�Փڟ�<rIgi$�F8�:�/~Ɩ�;Ej�H 
�%�z���g0`.�����P[ok�
ҽ�w�	^���h��c�a ������)f� �h#�XD�g�TON��=�7N���Y`C�1��vD���,�ƥ�a���Hd;u��l�d���Oe��*�SB��Aע�.�0��/���f�"�=(x:C���%�t��h6��y�i� =�F.qp�s�c-yu)u���Y�}k�f�TP���
�
N 4_ е�T�_K'9D��YА�`���<$�/m�pcI+����~)Sw�)9�L��ma��nmSDx�����c躔��*A��v���t�:1�A���p�F?��^C�a=�팔t9hE��ٖTƏ7!���We�ݲ	4,M�oA�U��'��B��KMs}�r�Y�N@L���2�x��(�}�
��S�S��r�H���<��c�w�x�P"An�m�m�.[k0������1?��G��&(5�F^!otQ���G:o\�o,^��������R�_.�K�P?�K��
���e�b�Z���n~z������&♟��p�q#ֵWNbd��N[`b����@$���؊"���(O��L�*!�u�?K�e��oZc�Yy��P!�~�8r�a�Y�'����~Ah���t;�E��;�6tI>a�(��v�$pA��zI��ۍ�� �߹�	T/%�~%n��a�u��Z���u�f/(ZB����V�U�G喙�+�6QZ (�]���x�JCUߊ��q�e�*f~�̅B .a Xɠ��b@��CtC0�{�Ӊp8:��q�my��F�A#-�����TZқ�ZL�KNTB���83��8硋�m��h(��ż7l��сOڹ�"u����&�Z �oo���528�m��e����q�uJ���!4��o}"h���q
s�����ʮ��^�%{�T��=�$R:�ۂ@}q���m=7���x������,J��)4��yQG���'i�v�/�.��N����)�9������:HlW�m�㗡�A{���Gw7�6Riֺ�2(+��
��H�U��ծUGH��h�p��AS�k2_�F#�P:;�c]��)h�}с �v�����̨���4?��⑚�T#�.��0��{��S�*Hy"��%��T�D$�>5�l~�S6�#T1���n���T��z,A"u7T?��-��G�?�\�;u�H��.`L�:�&*��k}�!���&����%��T�Ȓ�t�	��׶��wd�eԞ�Z-��wHș���
SAm�i���X�d{���jė�x)p'���U���!��ŷ���؆��1�
�b�1�r��(�C�� ���Ƙ�rI��M��e����O0L��LO�0glC�z&xD/��?zK�ǃ��_z8�tpvl�����;��<o�>b�V���Q�t�zr�(542�&�W����ҹ
�b�jÒ�������UI`G�ɣB��4�-��
���X�'>K�%ҚQb�'���Yw����nh=���`�pZJ��{��× ���,S�Kr(
��z�����
h�nS�����:���n�N���M�@=�>���$#��,��cʕ�I)yYP�����$=�gq�o1=�1�X�C�H~���[_P�����:���R��Ynj��d����jI���{%J҉Ⱥ���a-'� &�/��du�/y<}�(�J�"��V6�x]��h���FnI˽u/�Y���Ǵ�C�����V�BL�����;�e�	tD+��=ԯ�n��}��BpD;:�1A�? ��>U�a*:>�a�H�j�nX�".'.)���֕j��%w);.��l��Bv�i����Co���?C%i�kk~����C.��)2omGn}��!gY�<�("��[3P�bh��@
��p��`�\�?�`�j3K�[����~XW��jKqA~�䵸p?�p��I%̌��P�K��XT6��WR���t\�J��L<�?�LP]��s�k��B�x�x{�����2]b"��X�o}2�(zj��el>j�Ɯ0H�z��Ʌ
^���oBM���v\
,V?�ĥ�3�U%&��
ڰ�Y;Aq)e�8q��,��Rh�nm3�iS�4���XL%��p���x��1��9��HI�/��H��@I�eF���dNu��yE |�c��:y�.~J�t�X��9�UV�(��s7*Q��g�2Ed��`��~նI<� 9�x�40/�$��!�Z$H2p��Be���a���z����Vi�Vw���i����"����#%�6���.����>�N�jx�F�<���Z����;G�<���������s�d�o7�#:!�e@!��
��!Ck&]�V�F��k|' �?a[-����3H,H5����Vz1���7�G�o���1*=B�����au66T��\Hj��Gy�h�ZoѼO,�ɠ(������J�l������ٍ���Ȋ9t s��OS���ڄR��<
ZbF�0�pd��A�Ӳ�m�����dL$�w���K�Zy��lt�{��pD�ee�1���|���@@v�s^��F��~�׻7����[�d��oN��v����G���8���!��v�r���ݷ0�⢾�$Ǒ��;�y�	ö�Գe�JY��k��S�a�yR�~�Yq����Ur$�)�_��N/;��8�o`)D�	?����K-y��fgnA�?���X�-����p@h��C#	Ѷt��+���. aF'�gP�ch�@v�dܵ�EAbE��ҷ��ߩ��9����SԸGs	X|vF|g�9�j�����Dz��OoS=}�	UNl9A��s�O�蹌��!��[>�C+�u�#�#rKm���mf*^r]����ο�I��}{PeoB0+��jҽ�n& t=��1&��36*��7�!}+�Zr�+�!�?"N_���z����s����t���a�q1�7۞�Q�)�(��M��sG��݊[B�8�M,���9�;�^�ks�0��ӎcd�Qt��\��rG�I,iUI��Z0
��)�Jl���ƫ/�E�>���n@ �)��eB�5{���Z��p&�L�ŮW*�5�u( �/v���IІ��9��ske��I�-�V��@/M�Tb��(��Z@����p�J���7*��zy�,q�~2`W���N����c8ke�0��k�mV����F��__ rд<Nh\�`�:�Vևw&�Yc���V��vV�߼���?����3��'���	l+�zh.�j�E�)�#x"<�_`��_/O����'�'/{�lUyd���K�[/��8�[pj=Q�Xe8��ƒxd|���k�6c���Ĕ�Ĺoq`$�������w���	򳁪ZӾ������v��,:��Sf�n�%SnOQ�6a��Vg��q��X�dڞ����*�N��@�:~��a���V/DR�Ҷ�+i�{aM��c��"u�|q�+��@�����N8��5 �Ʒ��)�e�94�B U�T2O��9gx�����T�S�u1�B���^Y�=�m@Z�ܭ�N�֟P��\����Ѫ�7=��`�����#^�8�T��v|�}��㫤�{ R9���u<$#1�d1k]�g�����^��\	�Q��WLJO�����.�o�]5M���碵�v6"MA�,�;X�JK��b�{D>R�l��6L�jn���<6d�|��f�)�` D�+4]$Qx��
��Z;B�҆�ɴ۬��6�*]����Y�����hb@�]ij��B:Ԏ'-!D�%
�%�,�ADIon	�b\@YJ?ǆ?����n巊�^+y��q�q
�����j����k�85۫�]r��Iy� ���a�>�Q+��v����0�ӄ�A�bh�Xdޒ.�Җڽ�(@�p��S�q�3�k�N�B��׹�81ބZ"؃�Dd�YŬ`���2�jk���S��]�������Q�o���.	������c��`��oHG�²1gJ_u�	=Ad�<��w��[/_[H�D>��sxc�Fz_��3��}�Y�i�~e�0��AV�����K�@��GE�}gC;��=�Ab�?_k�.3�T��`i1CW�<���Ջs'uک{ɵ��ם. {�"
�]�̾J��[aV�qo9�)dn��֛u4��<�Yt��.U|E�-ZLXs﹁?����+'���)����s�[nAP&�r�b�	�q��n��5�� �0�J��>i��i�*�6�Br�!$	_������1��pX��l��n�3�^�T�[@�������{L6�~��"5�uj�"���r�8�W'�X]r[����M܀�H�?dc���������8��vF�QT��[P^��-��	x� @���㭪ٻwR����"�kG��§FL��	�&��ۻ��e�bK�~Vl���ԙY�'__�TJ�E�ŎY$���ċ*o�.�g�(Cڢ}���<���#<�16�+����iL ��0��N��"�V|�0N{�%��-��� �W)���_����� A��+��UH�ب��9;�ۊDKTW�5���	�WJ��ݭ�q��W�jR���d�)~����Q1�+Wa����� �U]`������Qq�M:�X�7Em#�.��j������+���S�!Z�pH#V���B���]����|q��E֍2�\����e.;�%7���Y6uP���+=��l���)�e�DT���Ig��C�Q�%EKU���
9׮LMw6vacc�F����뾸�G���ߜobOx�@Y'в��3�S�6ǹu�"�o2HBx:�8��L J�L�υ:����]o� �*dý�r$=o+�b/|���$J�rp��T���d�A�壭䠶�(5@H3/�djfC�<ݽ��l�1�Cd�~?���@4j|��*�
 ���u � ��JU�ly�>z[-�G�QB1��~j ��L�$),@���Y�'��9�*��i���C��Y�sl�8U}b���D���}~�koX�AA^�ܢGǗ��0$C�&7�`�؃=��u��S��\t��s���I�޻  ��6���հ(l�%#�Un��}��]�3ܮw�ٱ_>����-�xW�_�Z�����[�uyD������Avh�I�Ja��Fo�ƙ�:.�4���?��}���n���'t�[ա	��8��|�6
�'8�r�(����>�}��.)Q�Z����\?��p�0����hl������䏮�f����F���!��hr����_y��~�V��`�z�]�gmǅ�X�"�)29��o(Z�0;dz�@h�_g<��q�@�;�a��QpiyHNN֝V5���'.J�tΟ�o���$qX+� ���J�Y���Yu�������G�@*:Z��'@��z�s��
Ŭ�\��b�q�<�ɃKi��� �M���1U^��1#>�כ��:�<v��`I���J��{���1���:���./����={���W�
q�?��ݞ�K~�`�g���a� �/��Hn��䞳t�Dرs�ѐ��/��
��������:M/?������d��%�4jy/�3V70�?���2�ʥ�i�iߡ�dP����(۩��^��1�ě��y�J?}�E$7h	����zY ��*���Q������͍e��>daD#8�J��#4y�9Z�P�{�/�ʫ�c}g� �M�g,����SS���������w����-�r��1M�,��TV&��rYP���Vɸ��=y���I��.�M���� ��@}���m��>z����^�M<�J���qX_�azHp+#��	����j,�Bȕj�����d���,�ro�HGy�[���^�Ӌ���@Թ�|����48�5��c���8�ͥ�U�[|�n�LDu�x����k�٪N��Z��ȅ���5;��BL���S���S��M���sb�N�`�LE� �۠3f;]H�>�ڷ��|�M[�4��j��.�ڡ5gkY3���=u�4�m�����92���t	���J/Ԑb6�Oy�%����7�$K��K<�r/�hO���'����௑1�� ��}�	`���#��a&�t*�9rO��d7sl�Jaw]b�x �ڳYz�|��l����Г�f�4`���,��x��r�ˁd	�(?�E���J��\���gEjM���4. �>*���w�_U����%8�/=�2�+)���%�4��,��S��-BU�D3ns�4o����yAf�����N9a��� ���'u�`RÓt�J뮠����c��=���c��)��>�'z���q�3�J1�#T�*@�Y �zj��(?��*��|�g�8���QS6o_ `��Ŵ�A����˖llXqƘP~x��iSƳ��ͭ��A�-k
��?<��X�  
L�e5B��� ^�4�P!�+"�)��!�1+����FX _���:��4�%�
������h�mJ&��&���j��]�)ǲ�1h��������nd�08I��Q��ߖ���K���-�~�0��g\G�n��z��A-*�TVJ�,S��*m�k6�c�:��w|�"`�)�����<皿����p�d\��O	�3���f�Z�@�G����2����j����4�������c��0\z��b ��T6���<��/��G(�?I�����mNl��e\w{�-�@P�)	C���w��I��)��'ի���9�&7�6�(OV�AƂ"\�h(g����i�2:TW�%y�_�!䫢��+���f��-���]:>XY�l�.��@L�3�Ԑ���L��\��:��mM��0��9Ϡ�|	E��l��74�7�,�-vӵڂ )'9AH/��x	�A��������a�ha�kz�{_f��t��X��4%��S�/��h��*ƥGt%����X\�M)/[j=wH��fT����Q����t܎c���?Ñ��m<��(��t�o���K�@��X`ND�q���Љ=6K#��z/(��F��
�MZ"���������R~�W�\y���1���3>����(�Cq�%^h94&�(m����� �'��^9��@fޚ�:�g�Q
������M�}�����0��3�����<	�$��H@<�Ā
�-t)�%nI�$6�.26笀6M���Ա�����I�%8�G|��.�{Y2��;nD�>��@F�$b�J�~��߳=��S�ld��z��2��������d"��!���y�{�۠�>hu�ױ��y�Rv���T樳��*�")��cF��+�4�dx�,�3:�Z�������X�u�5�d͆P%#}ND��p�{ہ���
�E+���g��l93\�2ZCA������� T�-<��x0
�?��}�^}�/�$0����Oμ/[_�U�~�K�@a=����0��qR��)�a�~]��C$�:D��x!xy@�M(�\��p��J�_P��~����)2��މ�62��\�:HVE����%*؏S���WɅ���.o�ڜs$M�i�!�����pNqO	��
Ź�R}��AS�[%�&�R���.�d�b:0��Ҧ�.��RUl�W�d2n�%D�����hL'ⵁ�X�:J��|z��Y��0	��pl&���l� s���~����b/N�9g�ER�$��EH��K��'ऻX�[aΩ��-AR&O?��pd�_�p�T��)�#˸�Z���u����w�\�9�ag���235#7u�yD�7Q2U2���OJ��	%�A�"3,��-�JٴWKCg*f��A�Q������O����E�@���}�2hݘA��H`�!�b!D �U-�L�����(���|����n]uڙX�1Jߏ��[�Sl5�p*O���^Z���o��	B�'>g�d��k����	���(�6&���+��v�����A ��V�ӥ:NX���/}��Ӳÿ�í���Cք�#�(}�B>�#�{��5��K��@OL1:7�^�-���ƄMg_���b��'?������f�I�U����N|�	�~�Y���$�l��'h#|YN0E���jA�t0�2��#|e���\[GD��Z �\�mKe����(9|�/�G�<%0�����n��"��X�	���Ƨ�����ݒ��),Z��_�%ђ-�s�,����a�ɂնa3|��9���T��79��0�o�@��+��1�LK�1���-	I
׾X��T��":��Sh��S��3ME��܍D�xG���j��y�l�D��|H��+���	��o#�?�7
��951U|��N!����S��`�oËp����v�]V�>4��8�^(w��C�"~�=�4���u鱧��.�3f�M9-�;��z����<	<	s������S��9�j+K-��ʿ37V�C�s=RkL eM� ~s�C!o'����\�}U�!����*a��%e��k��o�R6T���|V��l^�s�s�ڄ��/AkJ��c�$��(�	k�s�O���[�qQ+�1J������{&Һ!BBw�,�
�嶘�-3��#�EB���d�fʢ�̪j˼-+�g�S�$:8g;M�����hJX)��t���P?(�Ʀ�U?�w��R�����h����ҁ6G�*����U�K��0+��-M`������ ��%7H6aY��v
�GC촎�s	l/ܪ�o;�<y��a>�(�P�ǩV�")Z�*)��-	\��]�gMe��t�1&2�nT8�`�^O-������q����Z{
����H|yi�0������aX��c���@s �6
=W�`4�N(d9hrMь�L�����.�aD��h�rW�[��6F�c_F�մ� ��[(f#�|Q!�OJ>I���MҠR�^�*˺�Pʗ6+DAy�V�`�yB���V�Z�����:�4��׃��]:�g��^I�g�~
�0XM�;�.O�I%5��:��hY���@0G�>(~�e줫��.�b�R�G����:���6���X�U���l,�sd��}��7���οˤA�\�vIn�Q!G���M��ʂ���ĵ5�z����/�/j��0a�ϰ��a���^U�^���4��֚�QE����ҩ>Y~��Q�K�>X��g���L.z>��m�w��n���{	��j�#%@�y��fZ?�pQq� y���Op�����-����dPyn0I��*x�%~���+s$A|#���.�����Q�ţ0�����DZ�t>A���������3�
e�9�`��#�A/��N�
٠���Sa��w���#︅\��Dz�a�6��m�����$�P�h���@n)K��,Oc��w��1tJr49א̈́o��~�c.b�U��Nmz���
���*Q�r�ks�A���p��8 ◁�Ը�(&�|W�v*Dər6OK��r��16;��N���ş�u�&����t�y��L�n�~7��P�Ď�u��d%���n�"��岎}�22t���LA ���	�V����+Q�:(�+^���	R1���|�_�i=�5�u��'?�5����-�{;�Xb���&�W �2%|8�e&�r���/�������5�E��O�:����L���4A q���w޲�V�I�5mP�j�a�csY�E��G9��]a���i]RX��`�<o��i��0U�+�-�7��$���oqj��J��$W���^J�MD����=WC���"W�@J�n���ͭ������}P�1]��V8؏�v�}��ȉ����Td'�˗�2��B�K[���� tKP�q���
��^,u��^3�h�Z��c��� 4�6��\{&.w����SG��\����՜B�c��T�
u��<$݆b�k� ��%���\D��d3�*/�wZF��_$��\r[���d�A����k���_MN�r�E�1���\�_�W�xA%����3v��%�Mq!��3��n�r�S�q��C�>̋�G)�5�&��pGP��hoѬ8�����QG1���'����Y�k�7t�M0��������� ��&���&z�(�Q�0~��?`�`�S�>��`n���dGT����Jw_c�kKk��;���_�=r`%�g����N��忆���?8y�R}.J=2�Ou�aZH��g����*fhؿ���ZV�2�6?�ol[��˸��>5s��5s�+�,|�v>&3oֱt���^�ʱȧ#�#�&:�r֌�-%�6��0��@�y���TJV]����`H��a�B�+GL)
s62�`��%{?�����F��4\����T��q9A��ff�B��G�����Q�����>�R�|�?�|�V�4�Ļ�����k��U�M�wpʬ���| �K.a���q�C`���|cC��&\c�������"�|u�	����]R�(KSЫ�U^N�@tl�R����[ �����O[GSX;�\R����W���|"��]�xNB�B�]�����֞��U����2m�ӿrLۡ�b�`����z0j ��{��yp�#)�FV�k�h��9,�(������C�w��(_!6�SE�aU��yH�=�\W&/;����;s���`���t�AJ�m�h���۫�HdU���v�oؐ,��j7����E(���E�Ő��Z��-_JC������.�����6�|}�5���$a�MoדT"�� ���w[
M6��h�LFM	�G�2y<�"�:�|�k�3.����;<w6���bMFf�Q�c�K+6��/��;�hb�,�� �<2��3U�H����b�� +j�j�%����ꨌ]7|d�����nY-j�td�Vm���z��x>Ȟcޛ��g�����P��y\Z>T���&�j�R�����O0�<�1��9�i���)�ěƆ��%���M4+w}�ȓ$�^��_�cK�����P�/���v`r �R����h�cj�ۈ�LSv��Z��j�G�HI��E+��;�` }�,�6$�`�h8�_]���>��� .���]!D��y� ����>���ߙߏ_ڋ��i+�e±�q	�,���g]LM(^�0���P��l���6oS��f����ג���O�#��ߴ658NA7'ș��6)��p�e��><��z��/F���M��� ����e����Ł�e}�f�R��������sw�5�����v����"%5#��P%��:��,^�/��Z@�apT�,,�43q!�ٿ�b���c�Vb2NE��va���P���!Jz�+~�om̜w�G=���V�$�i����܁v�C��)���GH�~�je���?����࿐̏�\'_��u��c=|g�=�.N�'z܆.fg10�)�05�(݁��{� �q��F��6	�vP�1�)ɰ�T�,�;v����9�󡿤��1dIJ�����皾�U���lz@nh�I��V�Ы�F�%.��v@���`3�(W�KZ�/ Nw��פH�L���Ն�����#GSPǙ�)n�>�������}�ګ?n����v�� ��ޒ�z?���`�Xq�U�""�#�2���k*E��Rx��j��#z����6�W����Y?���1p�Z	�k`L�,�Ҍ�͞]6YF�7|I�=�x{��<bRa��sƔ3��_5�yu�k��U(�7�:\�4��H�-����^[4^b��?I,Z�Y"��Zl�x��X%)/?��Ы�ϧA�ß�4e�
��c���5.򘿣�}hlQ|%#?��j�@#:�:���j��Y��-�Fjl,�A�A!��C`Nύ
�E��:Oup��}��VZ͡>7�%�Ӌ����y{�4g�wb&��ۡ�'`s��s�ϐ�d�34��u�]/xrЍ���k�b�%�5�{[㢶�F��ρ�o�2�E9�ī.���v��ytF|
��ijo�'�A_l�Q|ͱr7�;;E�>�8 ��M����]�Np�Ƽ���ۼ��S�#��t�v��gH�µ];x��n�͍��{ɨ���v��h3:v��?���v���bˢ_)�ېY��(	����>f���}��U���u������+�Bw�l�_�CJXP����eG@��Y��|�7��A��}Э=5�J贈�$a5�o��ݶ���~�q�!���$HOG�.���)�n,�-��v� :�Ԕ���cc�r&���̅�z�2	,�qR��M��~��mGT�~	�X�V�g���-uB)S�7��$��A:�t����Cӊ��/�O�Y_�Ѻ��bj�^p�d�^[)
��DĞ��4�0T$	�.M��Ds#�l�w]���鉱"�0�_�l"p���N���[��ާ�xCz�d�m��O�r��.�Y�t�4�el3'�W��9����W�B$�#B�@�!�U�8�oe���T"��3�*��^36�őt�3�a���-�E�Y
1���ᱣ�O��1�4�W��aQ�5�̮̎O��kw��Ԕ��7y ��)��� �Q�u�r�e'�b�.|� kCz�I�k�K�H��\(������FB@��bՎ헧O�Ib��q�k�h
W��I)	�Q����t�<_| �!
�A�9BԳ�
)�7�+`��]�׎ o`V�F�%�Xĳ�[Pm4No�4<�P����և��اP�Ua��c�!�"\0����k�{t`�D��͔�c��Gk%w�����P���xM-�73��k�<[�&:ЀL�'�����gffS�yI�R����/�$�#�Y������F��W�x���(_v��@k9��μؐ�
%ޔ�1����/Ȭd�V+�u��wlU�m[3=��wƀ���fΎ�fuf��������t:|.���P�P��nv��N7��joE����)�'�9�Z������I����5��<5���v�ho6�\�F0��2~��!3*()����C/���?��=���a��X��R!�-D���z����=�jB(���K-�17���^��j�R�Wo5ٷ�C�=�ǎ9ۊ��R �g�u����F��QK��J�<�����U�T�<�1��&�������7a��Fq8
|�̞eEK�z����bd�Et_\��:0����"7�1��.��>n�m+��fa3��p@4I����#��Ѫj`�ę��p�t��#���i��p>�b�C���x���)�l��6�h@\w8���;?�:��TV3�"�����Up_�5#8-�NC�$��Z���g�G�W	����	T&�]Zu��9MK��7z��"�ߦğhe�72Ǫ��$�W�@q�-~�o8^�(҇Q�PG[D�%�;Dk�y j�e)��_��<����N�}3�v����5�I�� '�)�H.��k̖@�:��h�v�_���|A��f9�]���22��I��;�:�[�O���E�z�Dɽ�q|eP1��%�Fk�K���j	��f��V��G�����9tj�̏�d�IJ���Cl!Eڄ+ݘ��D�,�7�IGzڢ�뽂��'�"5�hN�V<�xᏪ�.Ӝn� ����Kb����g*�_��M��}t��w>�(9����+�l��jA�	E���t��oK��M��¥�c:�H#�>c2C,�w�	�3���[�'�GVf؎��򹸃��?(�����t����<�*s�0��SH(�=�x�U_Ҽ�Չ��A�*����c�Ya燐��dAg���	�.�ۋ��h7ԼX�*�~U�1�M��*<�� ~۴��Z&�NT���ЧV[��U�S�d�{�j'���4�{:��_B��*E[�����az\-�?G�WM�E����q�-H7�&Y��`�s7Xl:��I�H�r��I6�1}A�q?��1_R�{�	AU�.ҫmH�Ty�7��h�k�?d\.�;Gwl�a��$V���徘��1՜$H�o9ý�&�=�EG�������M�uGGEl	�P��=x-��8G���415h����A6��E�CÝ��{ܟ6��cw
��4�l�\�P7G15�'��?�ñ����M5��_
[r�ҥ7���AE�RXzC)�<��%Sw�%Fd���!l3|��Ȱy����cu�E%�G��Ǣ)�W��Y�%�;��,ϗ5���0���z0XM�rRC+j�&`®/����-$�^g�+uk�xb֚{�� ���dToxkn�_�3�
��=�WZ���/hgA�cN�\��4�iFd�j`fiLf;ǥ\�I�<)�G�t��Yc'1B��Y��v'��JuUw���dcn�_��A�5���y����C�<��]��Ԁ�f4���@I�Y�q��i.�}S�>?�r�j�y������K�j��6C �Ԫ�R1ϻ�h��G�P嬈{�psӦ3�t}�(�6X�0�=Xύ���6��W�b�^�(ĽEg�o�V�jew��Sx��,7o}�DUS����X?�R7�"���X�q ~C��5A��d]m��R�G>r���1j��(s���XAr��,���3�z�d#4���K��6���:�p����&�&�>I�^i1�.ŝ��PܧV�6���K彆��*(зЪ�N\b���ړ�j��
�*]i6�OҮ�v*�X@
>\���Jh�i7���Ӱ�Ȅ)�`�a�-��B����b�岏{_Q�%&�%�G�Ȍ���z�=u�|!n����3�Tu"���34+���Oms������'Mb�X��7�<�W�ג����
�E&' ��げ�"�y|{cUg<�Z�����\���I��J-O�;k������FS�%��HL��Z�O�@��?��r`lN�ؘe�Xe,�׍?yVc+$ǂg�0B>�j��G�e.�=t��i�N�X'���'I$�I���*}�tuh������Hp�AcY��D<��,fH�Cx������Q��cC���ߤ|��ܫ\�����3lZ^����[N���5)�ц�%	��<  � Ft1�??h�$���E"��2�����.@��֖��{���@�n�;�*Vr��S:=���L��4���7]Vw]��� J.�Br�-���T�u�����NHB?���
���Y�W��gQ���>3�h&1��?�����Om.�L��	�x|%���L�t�[�?1�$��Yc���0�i����K1��:�L�?��*ƣ�o{n��Z�	�3_��Whb�,qc�Ģېi�e� �OJl�3지[X�����{S�U87�+>���U���&9������ V�6��͝���9�k����Ҫ���/P�e|���l�WE[%/��*U�#V�"g�ͬ�:c{�W3�>�\Œ�Np�е��,���XM�J���:� !x(-,�0����MM��t1[��_�G&U�t�T���	fR�_������҇+�=>Ƚu��H�g����z�2#�8,�]��#(Ͳ-���3���z*��"s���kJr#��\6_��y���L�_����̫�&�.�݊2o5m�:)LH\jK��$Sa��e� �o�-��l%���`1���."�}���۵��]旈bߦP�]�`Ӑ��jm�	V�3���?3�����8�CW����I�
8�c�rP�.Ki~��-`D�ZȚ[u&��r��%�����#y#�J��)�v�?@�7�'��L����Pl�Q�S�ǽcƄ�;i(����\� �Kҹ����h	��z+�l��ַ�}���-a��������$���?t��2t)���u�3	�^/=��I�h�N0�1Z�9����F��{iWJ͗�%�t#�0�n{D~<f���s��~��e��˗�!;�$7�BbFj��*H�$�}iO��&�&��>Vb��Z��,��V�)Lo����7K#���+�K��v���OD�Z��G��u�-�2F�N��Pz{�F¨ �3:r�����ħhB����u�c:Y��1b�+�_�9��j�����c�z5���.�F��NWW0(@�8��n^�2	��{��[�3)�u�Ś��KI����K�RC77o���(�ɮ�0(&&�z�H��z_��R֖S&��~g��99�w9�̚�
��GE]R��MJc~����;�N��p�v���R(�%O3ʁ:3�t��^y�W�_���'���؜c��b&�Ń�Li���?�5*���aϞq�4&��aI/vL���
x�I��m�jW��/b��L�&�uy�z��:���2�~SU�ɮ��1<MM�⺇����{A
�POzD�Ppx�42�6ށK��W�S|����!($oV��P����Uzi��ـ��W��3Zٛq��Ԝ0K3���г���i��-�`��)��u����z~*.�fk�	�w)^v���3���P�M`��(��e��(˖1�Y��;-:�׏PyYD��Ѝ�@��)܏c� }e��w���%VQ�����9Δy�Υ�!;k�[�eB@�N=R��R�����o�$�脵�2��H����������ТZ�	��/)T���_4'�+��(hb��ϕ� n/1�_qA������b{����ݭ\C�L_G���E��v�S
)����]R.��d�i�d<_#>�#P'�_@����@>���5�2�F�����$TwO\�c�=�K޵�&�0DŖ[{��|3m�=���g���M��@0�p�����m&Gy~�g��&�ex�Hs#���U���sT����C�p���5Mdn�I�<�ב{an�����T��6Cf@����e��)�+ܚ�a���HC�č&B�C#\�B��� �����e�k�,�O�"ι Po�@[.蜊�L��OQK�^k�M֘��������?�w|;���b�n7ւ�Yz�i��v��t���W�C)�H	�u1��Yp̈E�*���S�U�%�߁	m&xJj��0k���}nU�h
g.�����%O��8���`M������kZ��x���f��h�I�8|C���M�y��ݺ�q��\�Id�:ŎEŰܷ"���(��z)��t�׊����
QA��Z�3Y�.�yڱ v�X�J4��Al��������K�v# pfqe�)^2�୍\�[+rb�?�*C�f���2�n�v�jbrD���H���b�K�[qj"q�-��-�g9��V��њ��҂>��|�Zؽ!>�E��w�D���&|��R���*��cY<r�iֱ�-�-�+��p6\1F��L��^�1�� �6HBg}��x��d�*s����~�ZŎ��j��b�r��eЍ/���|�7��7�,1$���ʞ�Od^�y�@��)��dp��I([6.}�7�߸��ʂUDe�U���k�H���>*�[��&�iŜQM��"�q'��s�O9�̾8��0���]4�qs�y49�� �QC�CI�x��RƎ���܏��$}b�����lY�;BSB{d�d��Ua>Y�xGo�#)��Wʥ�Nl�!�1�}�̖"�DQ��E
�氭Su���}�(����E�<��,���&R���{[P��~�ȼ0����!�xљm�s�i�������Y@T��u�'	�aL���m@��P��<��wϞ�E�ߖY��� j�Xh2ϢQ���$뼈H�_A��	�Q��^E�G�Fڥ�6�ב,�㎠�ֲq�T5��oYHs�c҉�d�������,�� �m }BޛS �,��~~�	�<��*P���P3�-������!~栻�0�$l^h='����~p�^3��8��k���yQ�L(g�mC���9�ƷXA�R�����5�im�|�V������h���7A�����&1�jn�J�N9@�똽��Sx��+@"ݏ@��G���ÆbEʏ�m��q�|�H�7��G�~���R��l V�t��GN��R�a�A�'�AX[���~�<0���HVB�XV���`bO�`�/�c�cW�����S�YU�ےZ�s���I2m4���_0a�]&�k���'k��1��HL�bd����(k�A���
P���3
o����u��KAZt����^̛�Ӭ��O.)�gZ�Y(��č���s�h#bU ����͵W�̂6)b�s���i�b;��+��Ku���`��9��֞/��j}m��ѯp?!���т/*�͌�:	�+o^I��g'��(�N�V��^,~8`D.���%��R��������W�/QT�m+��.q5��M�����`�TK!�A�孫�J6�yO�ơzOU^r�Z7R�"Ct���sR�ÿn�g����(�df�<���b�k5J��~�gZ�wVo<��A���o���@v��:zʼ�k���:����sqb�@7R��l�+iCr�	��
s��;O�*�kJѭ!D�W,c� Fi�� ���ᚸ�T�:�=�0��\\�3��峢��M>�+ �x�m�<��	�P��=������\���6v�nĞ��9�}+K�3$�X����%���Z~n� �W�" ��'�8���+7̧� �_*A6a�w��?�c�[(ߧ��t��j�A7��Y�Ϊ��	��mo���WX`h"��]��ŗs_��y���dPn�J1��;��5&v�� ��0�7�ۄM�A �z,���T��\������#���9	������✏R�'��xJ,
�s3��۠W!������
�o��))3���	E�Q�z ��a���M\q�c�B��0ے@�-���ڃ5���p�R����G���5%�9|�]��"�n�yO�S���J�n��С�V��*�9s�h��v�Ýj}1X޾sQ����X�9�Yʣ�$���!b2kX�d�(v�D�b�d�
�p�?Bw?��wv��6dD_�6�?z�V��r���@3���?��jA�Zqú�Q��QE�s����k�|fO��5�u>>:�~1�C:<�E�Kt����AeP( ݮ��ټ$���T<�	[�|^��+�"٣�	��$P���!�d᤯��;z����v�$�����{$��-a'�>�I����A=���/?$j��$+5 !\��$2�HS��T�
�-8����o�(��5�{c,�n3T%�ܡ�.z�3(�k�j�ů�2�Y���Ey=r~vC�0<c�!� 8I�� p��s����g`0�v1	�*������DH�z�6�vH"�q����iw�/��8y�����W�ϙ�p_4^1Տ���&e߳������xڄX��lQ�(���v�b�Q��K��j	b#�8�?x���5��/���5�[!D�Cz����:A�D�=d!w��MsUWY��be<`�aZM�ם5�LTU�tZ���68
���C^E�ѣ���@&��;:w�t��,Y8�j��w���������#�|��V�_z�O�����h��6�-J�Sӵ�lK���+T��gYšT��Tg�;�çU-�6|H6�Q	F޳�腆!���Z����.��`����Gs����5�qQ�=����=XR(�	�U�
�p��m9��kެ�ElT���b�T�n������~���c�~-~Ww��w����-�кe�D��q���3O|3����	�og�زU}G��ΐX(��C��0�K}L�hi1`��#��dMy`k3D��{su��������n�3	�΁|Q���!G�/�r~�Pk{�ӝ_�H+��/~z	"I)�W�.*��
$��o�D�K�Э!d?���Npm�jR����%)�ؚ���t��IrҴS��/KJ���&��ɍ�E�P�Kr������\[���
�Θ�Ȫ�a*D���`�A9��H'^���zw=E��T���Z\t3A��zOlh���)wL�_�n# ��+\����f��MfqVє�ix��(�\���$x��a��\�Q���p/��Mxq�#�� P���g �#z�pV�����x�x㞒t�p&f�1U3�.Ļ��A��5�$t�3�'�M�g5R�.��Ԑ�d��|���	{����K�Ө�&�7y#��E���>b��2�j?P�r���X=�zŹ�$�p
���m�Լv �jfo��~BE��T�$���	R"�?�a�/�Q��F�ZDEʻ:�(��2�)��C�<!��FE�]����V�Oe�W\��׀d
p��.K�X�R%�Դ��6u�P�cocE�V�~�@j��Gȩ="�����'��mA@�<��&��lBSk��Yð���!^4Go�>=lf���7����v����l'����Dy�W<�jh��������/�ݨ�����H�K��]�����ܝ(z���ț<���}�}8ˍ4c@PbҔ1���8�:i]h?��I�p�)���@+��*)5"ͪ���D5�02�h�z��˦|[��C���O���NL��
�UW�����;�'S&���D�����HB	���ڱb��׺7��<fp]�����e��zg�����xϦ��J�>��=�{=��#�]�_]^Y��B^�ƹ�;C"Ӣ��"�Ӈ�E�3DZP���
�d�GK�
�+�f��}(���j��A��M͜b��y��6�8��;��4D�w��m|.�w�h�ˑ��{�ɧ_u�{d����?�hCJM��`|J�Hv���+��pں0)�Źc�:��ACh����wd���]��J�k�)�<���:�w���-CFÃ����/�B֦CF�f�'_�WZt	6<�'����i��9��!�����Q
��Lc����i�؛��v���d� �М_?4����VA��q�5�V�������Cl��÷����%p&B���M����8�N�B�v�W�X��� >����C�`�O��;���!���!�^rֺ��	�k�L6O.�A�Yi����~���$��P��᫐�q��~4���>@�S �8O�%���$UjT�����D.��U�V��wH�Q�93�,��KrC�s�ԅ�����.�1ec�d�iԯ1�0� �?��eV�̩���濉�� ���(�pV�(�6�c��N�Y#e�b�,�������2�Iu�?Z?Ւ��"��w�
_��|�4@D�JlU]��9�Gm8{���x.�*u&�B���f������-I��'��._����/?B�+���!��}�d�=��:Zd0u�+���?�r������
-B�/�?r�VU��'����!ޤ0��I�R��␼��c����2�>����~Y-��3����q`�+im�8و������mNݱoO��3�$�֮v??	�i<C�d]��)xy��^��g�0V��O���>~�3�0О���>�GB�D�/�G�һ�=����֎���zZgr�C����#���!��y(���LGޱ�p��Q���H��l�&�p��{�~�m�v��;T�q����}��I	خ"e���v�'=�f�o���uT�G3Υ�j�i�[�	�a ��i��lm��l�k7y�f�
6�f��^�ђ�<��̇�Ĥ�`mٯ�gV�5A�_�|�0w�|̣(�떾�"�ie-H���� 	a��4�D.�&��pS
���E�-�SE�U�*��cͷA�GT3��ܥlZ����ybv��;��~̞�h%��$� � GӣA�
�;���N��˸[9����]�4�*bJ����]�'���ȍ�-5�X��2w.�8:P��8�>����Q4I3?���Gt2�* R��������[�%#`�fi�n��9LX��7����=�J����	��!���k8�a.����察֎��;
b>��޶hGo��3�죊��w�.m�S��II ���
��E��#�{T�S�Q��K�Ű�K�8��S�]H�� �K*�i��r^Mj�:�~�D;94���u`~$�4��Z��kɲQ��}�o��8�l�}���O[R��A�Y���k!׆o���, ^k��e��*w������}�d�-К��[����"m��ț"´G�P%�:C�(����s�:��R�pJ���e��e��q ��[�	���Hb�OM9�a;E�C���nʃVԸI=Զ������==dmN$Y@v6��v<�^�K��<�b�f�p2�8f��0!��xZмv��Guٹ���Z��$��z�#Y���^M�?M%y��%o�&��$�$��H�J���E~p���ya����G�1� M�
,x*}oK}ƈp�5������>��F�ePpO�����n/�a�@���3��B�^yR?�z�V���LA#�E��9S*<�+��r��������U���㈜��f��rrI��\iPB�%nCt���5H�_|?ꀇ[,KcF+����5��{���
3�0m�-~���Zn��/K�ვ%#�~�$��">�fLA�cd��{�ήݷjs��
.ʂ�	�Z�+�nq���c�abO�S0���.�F n�oj���5+��k��w˛&�{߇1s*��e�1��fʾ�Ͼ@����W��FR���"[]�}`��f?%�|r�.N���Բ����E��Y1�!���ς&׳���j<άw��O���w����2*��ǮM��1E����f� 歙J�~Ki����JY��t�y<
�M=����HP��ƋcP��&��`
b~߅P�ՌI[�����������pv(�R���r�L។� K�=�<iG�t�����.995��|���~z��� �f���z�LA�W@�F��{1VB�p����'������)�����j�}��T}Pw��@N���� @#�{l�X�]���
!1;A��P�E���S7�>`������m���u��![�����<T5A�~*�������}���Ş���ó�B/�I���K�I��F���V�ߏ�2m�� ~�|�^��f����X.����R�Ӳ#A(Tq?6,�Y��#������S��AJ�w+ ���P�w�^!���`�}��K�K�]o��.�*�2�����7�yC���������4;dy8�^0x��U��;��j�Jm�ځg����9��R7�8h4V�fX�Y�t�l/G\��+�qr�R���e00��n�I�VQ�(ߝ�U���v����ݷ����zo��Ǚh�/s{m 4�D�9ʚv�7����_�<2�h���И��y�)�_��	Yc�����4)Ǻ������:{���,!�r1��bB�&�F��I�d������zz8�5`M��^E��|Oc�C֤{�oA���]v���Æ����lY�.�+J㱟�a.�}k�.�B���yۂC�ó��I�(A/b�w�)ז�mu�x^�H�%�����n���Ɣq/"�fI#;�^y,�Vw�(�9�k[������P�;��s����Zý}��I0w3ǯE��箦oM���#ܗm`��?<�����?X?m
'Bby
BW�׹�/a0���GiهC`�%m�M�q碠F-��$���Ї�%�
��נ����/��)�p��y������NSb(�����:�Y�ա�6�[���ba���+����Zt2�5b:��Nϛ�ҸK���y�t׊�n��-�ى���3�5�X"�l�N�1�Q������7߉ζv�+� �����ϛR��*�w����v�Wd�Ğ�4�ͳ���t��~}���O��L�����ʖ`�0���<������TSXfu����VuUՈ���srT5ђ�IZ�����H�g7o���\�X�a���1��g��G8�>�_V��ލXJ(!�?&�'�j�hq�7xR���,����d8s�6�N��~j�_'�3��εK�x��w#�	@5���+I�=���>`�G����j����Rz�F,I2.E5b��l}ٮcC]D�U$[
��@���g�=p�\'��%�,���:�k���&��/�À���$]�(.����4O��9�S�.2�z"��n��uy�z��+�x��E�� ���a�9W��U�a�*�9�o��.�|p�4 `��v��~��D��N↠Alӎ�㷚U܉gY���W[�"Ē_�^�����2#��(��]�ݹ�������Xh�2c����a���)*�k��߃��D�'چ����2W���:�jȀ�N8_dݢ� �N��.�#�v�lq���#��@O�e��՘in�4�)�J3f5��&/Yf����u_�(�	e�>ӹ֔�;YZĒ
�����`L-[_�~�P���x�'��o�{�����.)�:��Eٺ#�xL��s�$tauEؖ�MbRm<�8�7`�]���̟ŝݮ<�]C)O�S�-�:������X|#G͌L���T��!3�J*���vK��_�@�7���G�GAFF}S��I�b��~U+S�r�
�s��2Ҿ��N�O�o�$`R�,h������ d�4�u��rQ�����5V�Y<Z��_�l������5�u�_մ���Z|���WJ2kS�4���KlU�C��������Yb����BA.�����E$�ݕ��=��I�h��%�tމ r�}�A�ӱW��"������d@���B&@��~�}g�{���T��cC(�v����ʞ�vH�T��O��,�9-0]7/ڀ������e^������af;y��U�1n���ǲ��rh�j����{ua\�!֥p&��^PGǐ��T�������e�>�y�6{Ab~��[)B�߉��~� ���)]���&�q�{�0��J�v���v�����\���-Z�a!��9A	~L���/�J[ԕ,����+4_)Xy�Um��7�J�0=��:$>5�?�KF&�<o��i�}R���Vah�k����gylO
��g��]��4�E��/׌\���[���I����p����])�y��	�\uԦن8I�\j���ȕ[^�8��;[��$��Ҷ��  �r�>���Uɇ.�;�nn}I�����_����ՁU%��%R�{}�1�S��P3���F>7�����]��0ʟ���/UPi��j5l��f��H��aǒWC����;v�	>�(�Y|��}Y+�bL����.��#Yyj�N�����vi�B}0J�9j~ªP{�fa�9��z(X�c?���쎧�Z$ ��瘬�[h�����*�l�]��$�d����	h��Z�@:3ǖ�5�Hݬw�����a���E�@���j�&d�g�;�Wa~���~���a�<j�-i�����m��'�����������O��]�Ř�Mv*O�ӌYri������8 P�?�|��1�Yz�K�,��)\	�I���\�"��1����%��$=��a8�	!'�tN{����0ʹl��D�پ�^3[TG_7g���O��_����߲ٓ���X���˨v��B�~�.5�ZO|�7a�5%����㍹���F4����/1���Go�.\��Ƈ�Fڝ2Y�</5`�����Q6y��!��nv*��`�v�L�@2Ҿ������)�b� Z��cK���+��W��C�5tG���g4c��[|���`�Ln��U}���%����5X������f��Pm��d>[�z�#��.]9 o�ABGWYC�����Sr��9!~�-�o/祸�\y��o��& �	��2��j�>��h�j��q�q�>��-�+�3LQ-�>q\�	���J�(I�Fx��j:���\5B�Qus�����Y��քs.�B+n�YY+<�sĞ�U�?�oQ`6���!����'�U�@)}��cA��s����1O�Hn̙�)��\���&s6��n|ȏg���uVTUv�}YT����[$�g�\����K�3N�Eo��w�Q3����c�+s8���z�+�2u4E��a�$�d!jT{�}�5��S�����w�P��hC�
rJU��;.��Y�_8��z��F���I�^�J�y&٘�C��s��i�+Zs3�&@�^���܋��L��)����Z�Q�6JK���U�񑪻*c�1T���%�����3��VY�˅�Z\0BT���3M��-�;Z���-k _l�}��"��v>���5oUUӃ?��kH�w3��9־��	��V#nJкcz�Y���T�)�J� ��N��P���moa�fʖ>�G=m�q�hN=�<���\�u���l�/UC&~2�S��qkfC�G>}�b���y��ظ��3�ʝzF܀S森
Kbi��H�|;���~�`��������<Į8�I��q��;����C�9��a=�Z��9�C�\D`HT�8�~Gk��9����9C�}��*fB�:�S�-��� G��%Ց�S�o�y�����\ϕZy��>��0��X���ʞ�m@a?A�{p�w�����k���{�����D+3��1�	yY�g��Ff\$���{�4�`����0?�\x�%~uz�2ߺ	�fOi��7+V%�����o���@W��Gs;�����|_�g�$��1�J3{�դHy�m&��EG���f'��.^VQC� +j��>����F¢�g�ṱ�״�T����V���^�o������\{W`������s2���n_�;�"�WG��b��ꄴ�K�e�CO���{�hB����
)��,����[߻�tE�A�
}���u����ko�	����̂x�=.[��.�9���=��&(�������f����bZ��<���6���
�|�~�����T��@�����&�B_���7�P�����6pRE8�X?{��F�;��"J�J�|*�V���e�--�r�*�@�b��]��s��a���:�<�pA�2����(.�y�"Q+�UV~�jV�h�R��f�bwUs���=�n��7��ܑ�B��h�8P��2�=�Cc�FF@Swt�!}�v`�<`���*�s�����a�f�}�{J��M.��@�_����a^�՘�I�-&����@hR��I�K��5Y��%С�����Y�fq��\>�Ⱦua%_�b������GcJG��Uˇ���1'����(��ͻ49�3^��mP�d�L����((�WZ8nHk��^�Q3�tI�2ߐ��Լ���g�E6�3(���9����@����~ߣ���BR5��H����~���d��Ȑ���Ǻ�{A�P>�ޥ�Y7������Nk�P�?�#���D=W����ھEP��jR^�,�Z�^9:2$�H�G��ԯ
S�(�� ;�U�T0���K�F I��!B3�/�"Đ�٫$�L��ld%��@]����>9��X���_�m4@ˈ�ɦ�4�+@�Bb��]���:'�� Ǡ��s�f�ϐO���gm�y�ƴ7���4���a`<$��U�BT7��~�X���βR��i$�̀[���ݯ��"�]�O�&�VQ� �Idq
��G�K�<`vN��|�'C.=���2~��1ٝ�{V',:7���Ӏ�5Bs�Q��4���T��X�ӎ[ht�~���|=�G>]�"��)>�����@���i���"!c��:~�=E�Aا���j�uTz�//4� 9��3�,��F&�End4��,�䳲�k�R.��j��-��0�ܺ��[�r��C$m�zr
�ƈu�	y<�槡R �k��/s6J���x������n;Y)=p���ז�؎A�o_����7���5S���P��xY�#n��iE�e��}��ʘ��4&��J��W���,�̪��0f�.jmO�����C��&���� �7Y6��V}h��g錼P���?$I�Z�P<�	T�"��H4s�kp�'�]�s4I��$P����:���E
eG��I>K�����K�3Mu�c)b@��@CZB$����7�@6��5�A��\���Ͽ�����>H�*83?�������{�k��}���0���2Qf?�[:�p��x��*L,{"�H�����������J����B�_��Od6�#+��:�Sl��R�mԯA��}�v�.�b�$��v{@��U��^s�΍��.Ɓ3��ﲖ�����7K�	8�0y%|P��^jyu�D˓��{=��$��*�fa��f����[,"����wo�qћ�A���Q���[���g��]��&f���,�((xΞ�����+!����=���ٗ?��CB���/x;�����~��ی%��St�1���RC'%÷�._-��L�~�\U(`�)�� ��I`�"�Y�i��ju�'�C���������[M�BXh�F�y?�_E*!g��(�V�a��u�koAL�t�MnO�U�M�\�c"Y�N8�@?��u��������AT��d��sH�����q��}�޶�e<t&�د(!x6*�����l)���S�oG�)����u����8g.<�J #�r/��3�9f��ދy|�x{��I���K5�ES|�K)�w��U ��׃j���l�X]M���bj��At�4L����k�DO��G�I<3�om+���@��.��Ҳ��&s{9�X()�[�����,�d��8�bP�\�jf�r�>�R�^�hɳ�,��5l&��F|�܂Q(hV�kg�k�h2џ���z�5x�@�3ϴ�P�F��	]�To�����P����+ !52ꐪ�n��@�)w`��@%ɩp�T׈ĎT���є��+5���������T��<;c8�[�R�(XX���]u�p$���J[���Z�X4�[#8:u��H.Т���-�C��k�aƍ��B�>��:�;�n���T�N����#�u���ϵ�W��ΕK��ǂC��]5�W��D�9��5��$<���0-��.Ѫ��l�&ZFa��]m�C� v�i����纂4(a����n�4�w�tZ�r�J:gpp'%���+���)�E)��q��j +.�W�2W&������\%f@שS`�WD��X�NN:�����Yªv��=K�s�K�8	E����C�^���3�="q��H����ӂ�רKR%�_ �H\xt�)���6�q�����2��5�i��o��9+�Ԛ)�Ӿ�����`s�V��)_���������Sg�{*��f�[G�ߥ� �;n����n��,�H��N�tT5����¥���\^�&�9�{�|����K�\��I�ꥋ���F�7|V9c,,||�l0V�_4�;�TH*�a�M��W��P�)�V��QL��lI/��'sL$�qL�Z���6č�B(2i��V�ƹ)��j|�>7O��Ic�.N��<�}�$��W٥qZ�>e�r190��^O��L���������L K�m��6�����{������7@}�?K
f=���(���W���I�%�8�ȜƇ����.Q0��v>Gٱe�'?��\��S���Q��ᎊϻꆳE,��u�d\���!�vb`�=�
����%�F@�=%��S����28yb��IGq��JDP�Pj��^;?��NL)Y�{�k�����q�ǋv��vgyJ�a�+|�����{.�n0��		%t��GWtڸ�OC��-��[іU�f�s�Z�,7ɮ�w}S4��q�nF���� /���;r�7nI�I0�HB�磑�����!��!Z�{��-%n!��ѐ2y
���Z�=A����ܜ���?�R���ך�k�G!
D숙�1�
$�	�an��4���v�`�/���#q��ӕ2cђ�ې�~ٲ��<��Q�ﰝ�zjT�����ޝ����෣g���_m �P���B"����غypG�ڢ�ռ��ɨq.áf\[�2'ιَ���9�7�s����ǰ��	���.���y#~�M��>����{��|DD\L�q���,�jS��c'��y)H�	%[}�9 �=��q�jSx�)$eB�X�K�i��</��M�=��΂k��<����	v��A��^r<�	�u�0q��������f�]�ڍ��ʒ��w	�C�z7�2��a�5����gnЀ���RW�����H�>jZ��}8ڊ`o��v�7>��g�	#I�V�|�R$Ea9@�k�`�u������^�Z_+<H�ˀ,�"&,���� '�]1�B�\���G\�)��\4�ȿٷ��܏'A�h���po��b�
giZ��?�hx'n'?2�~���=�fI�ރ`�O8j�\���L2������a��c\�az�ah\��kGI�����UP��zx���.K}[�.�LV�x��
{�������d"��0��H�K��4:�M��KR!.��Om�].�`���t�%"��ɝ��'�f����
0�V�4NU���-̊h ���*�*�D��zb��Ȉ�Գ��仗���ٺ��zO
=����������:n���@�ac
Peum)lh|����;G����bb��h�M۞77V�1�: ���ĖA�Q
]�O���ƣ�%�E���}P��1�Nܸ����l 8D�g���I�=��NL!������� ��*�X#y��'2�V��!�1׏̃�����+�`֠Ɩv(��*��LPjmC�A������?̣�#2�דE�� �h�t��=F�%��Y���ߡԨUu�W��_����LH������ ���$�F�Êp�B\�e��6o�߅x��_���[K>�r�d~j��h$�ߪ�I�R��h$8=X�y,#m�jH�m>����� )����7C:���E,���]�@B	�ޥ�v&����V��m����U�@��e):��u
-�xĈ��S�E" �����OޔyΣ`&	�$=pK����BJbݥ�)�F�5�}km��O�8��k��8η��'�e��A���׼A�b�e������ �T5�+�i������*�\-����_U��a^�>�@⌘�M���@i�ue	���ҿO�t�l�w�n{�[�S ��I�%��GrJi��·���f�|v�Aye���1�p4����Ҋ���xKB+�H�d��C�Ӯt�E-9�P��{���s�v���Q>���\F#���A��D�|Ȍ���`��p8���� μ���Z?R�؝�8.�Q��×ㅽ� "�ܯmb���Ж�Ue�n�K�K>1�G� ��˰Y!��-
냸a�/7�K]�$��0)�����bm�ҟ*G�r|����?��)�%���㏳�ã���� ,R"�0��z��FAΟ�[��?q�d+��0����[��0�pW�٬�P;��*	�]�������/
M�˳і��P)���zX��jp��)�eum����x���ҙ�Q�+�ǖ��*�Pڄ�s�*��o�\c2H�v�M��7��yǐ�ZBK%N��4��;���T�*�"�yи�e���a�?bt�~��b��TC�F���<q3G%�?��Q|{FHm�A*��6�PwN�
cRm�Dl�&�E�!��+i�����t|��8�Tn�`Lʄ��������%�j%`$��(�:mFҪ a�h2w"��U��H��Ú-�^ŉ�>(�*6�D�����N��M��1k;���c�A���A�����d�	c�����:�A�1�5:��/M����_O�Cr���Wb�׾ ��g�^2�gK��V���m�-������em�E��^���Xet��O���;�Lkgd�,H(-���^-����'�P����,C0��Hsc��|�[OK�hT��Lk�v��u�m|{��k��n�i��^%咀f�(��ٴg��w4����]��"|����X��`�w����:����xR zv}Vo�n:��� ��H��"�7�!!��y���A$�$���_��X>s�w�Lj]t��������=y�;�h�X{�8��� �R[�`M]�`c���7�B�.�r��]T#�%nHk7�a�x�Dqq7o�����X��nß'X�3�Z�s?��HB�T��b�{8�J��l]�;�x�N�%��V>ex��h�a@��bEZeTR�fP�_7Z��_�1��bp�F^�-H:�M��	�X݋ڊ�5��c����w�)�	���RӖ֣�j�O��<�h�gO�ę	K��DCl��1u�xEڇ�0U^�E��D���,	d��>��J���n�c���(�L,� �"�� ��E���M��x���լ�\��6l�2>Zq�����	�S_e���3rғ�|22	�s*�
�%�F�	�	�Z(�2��_r��	 �uX�� g�z)i���|�����2���(i���0��]�#���S�׋z�
팝g_Ls��8�D�}q���-��Vu�.�h�k�5JW�Ē�|��ݪ{��r��e��7�|���p��r
�h9<>���h�!N�w��4�H0׻Ҿ-�f��:�<�4�{]�� ����Y��~C"��܉k\y�<Đ؎�����n���y��i\4���� _$3'���ιn�/`�mu�4$D�j�9�n�6�e.t��v:�R���(��l�*�-I�{� ��F5������$�,�u�9x��X�t�X��>Au��F�
�r"*F��O@S> d`56ՠ�ɖ��>�4�Jp��_�7���Ǳr�AӹN{�����?� mK��XBhf�[��<3R�gf��{������f
�[>�#��k�f�	�QS���ʗ p�5"��lt�[05}`���HšfY�_����UW����?�G�q�h��؋�N"A��?����t1��/^�<��'�l,��A��e�T�A�V>�C���u�Z�呂���m�>j�ZGF��7�$4I?�ލ;?�'���gc��~�[���i��* J�nm7�q~��5����Af2�<�G`��M�v�t���J�r�r�
*R^
J�s�E���%�[ Z�!C3p?.a�}�`S��ϕ���V�eA����	�j�!Uؤ�]����Rn�L����'��"&��>��J��+�Y_/ Cȵ��BH\Y��Kg�{y� N�5�����u'<���"��ϰL��︜���G��1`�ƫ�������WNDI��9��Za�n��+Ṥ�hD[:�c�xl�'��g��R�mD�UX��\ΐ��M2N�QW/�Ƨ����`
g�I���F� <��&�����	�'?ۋ�"��E]['�����Du�+��qx�A�h�Pʽ&0{`Ɋ��ʿv�(|oD��Qj�����ݯ����	Kl��-�����Fr�$��s�E��q����z�c���z����ZI�c}�.��8mW��ʰ/���s�r�{6��z�`n=��|K��#��`od�@��l���9�C�`��/��JA$?�b����d,xd��P�+7�6n.�)�.������,f;�+��v��%�|;���!R�4=��F������P\�9�ns��7�z eC7�Ѫ.֥%xP O)�cO��a�����fU��P�w�a�u��s��dLo�ji��sl�o�S���
%�>��a�n���� �Q���}�V��Y���z�	��f(6��M?�=����+�U�B��bu�#�=b4z��E�r��e�@��-�rx7uk'��د{S����Jd��m݃E��o�Y��.��{�������ĭ�<M�oٍ@�n�R2�!=����t�m f����ί/��P�^�}/^�9K�;�Q��2��d�`�v={�oM��+IzdF\ZA��m���%���Vg�R��G&�؂����f$ׅ�;��_��$d�o13uxx-�,�Bj����N��@L�|h�<5f^����� X�>�����v�_�a�@v����������w�Ǖ�	7�w��5=j<H#���?{�f]�d� �Z_5b�t3Os6^�]��(!�?���V�4�"�{��^�U��;J5��M�%!F%p�Z�p�u$���O
�]�f�YW2���f����DH��{�
�f��*\A���[�e���G���e.'��ŔR��w�}$׃P$��|�_T�_Ж��?v�[J��m���%�5��m����*��f��ao6�G���Y?��(�Ո�F��>��B�.�9\M�$2|/�pDӫ��������\�0�*i�S<B�9=E�-�ҿ�:'��-�)�'ǙEr�� �������d�<��Т =K�)ie~w���7|��Zy8�(z3>��p�f��x����j��y��3uq'
Y��!M�"�=��c�|�dB��2^p-,���T�4��z6�=���D���E.!���	]9:��ԝ'*���u^?
%!���&<ŬȎ�f�][�S`p*�d��y�&�dF]\\"�Ӿ��1����j	8Ќz��r��S�g���
#����U���9�@�Sݳ�=�y��5�Ι�^���,�������z�p�mC}c�S������g�\�8���┊��?��ψ����yI��}C*�����C"ML~!�\�C;�n�%�x�J[a��_"��,o�I��J��ڂ5l��c�҂Z+�<��pE����GHy�f��V��KN9V園㬍�(Ch�s�Ը��B�S7���qp�нoF�T�FQiW�!�B�r�����P"T��2Tj�J��)$(�!<}W�yO�w�7�W�Z��Գ4 e ��ǻ�9����:l�=]�]�h_ڪ�n�@~�d��tXRׅgI�^�(	���]�ɐ&�:Q���=�Iһ������kJ���?��2�K��b+�Gnv۶{y�\N���v�K~d:���#���Zل4l�[" 9�Z�Y�}I����/q-K���w�>������e�����M]���ɩ�|��V�3y�mN{�(wL�Ȝ�gpgU�f,H�����<��Ak�-�[[vl����WA֛/��� �ilR�Σ��P�"Y8�5_}�4��5�P@���m7@�i�r�h�m�$ڊ�Q<���ĩ6$�g�B��l���Vj��b�޻�a�-)+nՍ���֨
<�4Sʎ�]U�z��bW� �f����?E���i�o��6۷����+w�6+���L��~��U=��$q�\����Z�2׾�7�GW��=��l�>Ix����15�Д���n�f�?v�9�0��cL��,��$ahC
oId���*�}���G�z�>8Gq<�u�1_�;t��PH��eƒ�Aʑ�B��@��>EB7�b�����J���R`�`P�u��V.i�>M��T���(I�1�ԉ��$sVп��}�B{)��b��!d��p�8�a�<�O���됬�Z�*� :*�kπ���r���7"�V�j׽��=+8�Z�革*i���FṶ!>���L�����M�L��%�1�6�x����S����̈�=Tc���ܟߘn��tk}a���r7���4x��*��z��� �i����j��AEMM?|ݻK��j�H0��J�3̲UĎ*�H��璶�P�
\O@8B6�@p�ٰ��%�0c;x<AHYpD��ך��[�I�4��&�й���s����a<�m�E�]����_
����xFl̓?Ŭmo�Y+�A�51�8,xdj!x�A�B1��~	̍W�/M�T��v �5)��N��Ť�Z���&Rh�Qk_A[�r>�Q"z풊����H{6�pH7SN��s�!i��� �1,��n�aг	]Y�� �E+Igoψ���e����7-U��Z;k�,v �58�'�ڸ�<暛�Yx��8�>|I�� #[3�=�S�,��D8�W�~�ƥ(�q
娛��X����h���O�7�@������5��/-��6��#�F�{��7�b�o��jI\l��9�*�������H��^'*��R�.�c�wD�Z�j��x�TC`%3�b+a�n`����[�Ⱥ.�\0=o��',hhǟ�����q�d�Ku�V�<5\xy �T�[�ljl�ל2��)]z�	M`]�<!��;h�B�m+wo���B����S0�-�Q�c���$������d<S�x�ЋԚ���aOh�_�a+^���
^J��0$�y"S���UB_��wX^�H%�]G��Fr󬲇I䰵g�oY��Yڿ�Q��O�0N=�`W�+����,���m���p�j���Ca�EQd�F���$�a
��W&��v���"���:xhF�˺���Q��OaYf1|#`	R�"I�K,�(sn�'՜�T�eމ�,Wr�$�X�a�C(iv�F29t`3���o�Oi�{6}��`&I�x'}�Dh~����Z	Do��C\e�<��Zk�Ir�z�Jw�b���� �'�egX��Ύv>Ż� 3���]yڹ}o{�ٻ�? �45q���7A*�(��TP�H�dUJ�������;��j��X<�-ñ]�Cg�g�Kb�w��s���\7	Hf�sM��
ԫc���>P��i{�n⪤�-`��#�˛
&�_Pn�h�(�����4,PrV�2��-��n��F�<��a�E�'�UL�1c�}f߄(m�]`#���A��42<�e7���
����',5�Zv]�$����R��eZЯ��ӌ�/z=�HVJ>���,�l�րC�h�����ؠ��G���(��$Z%�q� 1�抟�	D�?5U��ώj=^������j����ћĩ���X��M6�N��&���q{���09�;��2�0I�{�=�Ԟ�����z�.�(����Y������~��NX�~�A�NV��W	F�,/
k��B�!�Ѿ+�+C�'^RV�tJE��W5xyݖ����
#*�~z�wd��1�ޚ��x�d�+��+�l���z(������~�"�-��LP;��DRҷ�zW��k�/X����յ��܊��v�U+T?��G�M*��8��;���C��y*1;#��Ah`�b�����ո�Ȥ��SA5˼���iݿ����n7��=��d�D�R���"d$�q�	��ʨ��vC�Q��3C<)��$R��K��ְ$����%�~�������ՌkO������}_��q��^�C�qr@}�-�3%�ٷӘ@�:]�O<S���T41zVSe<�N�p�o��@����#5,�����ة�BM����n��������<�r�),�U�Qu�����̍ia�p�� ������0���1��3|�h��g�_���:��æ?I�@ŏ'k�ߒO��Dũ�@AZ��ۿ\�xx�P�b��(p�:�e��2H����(,�TJ)I�����!����[��`�`�'�Ώ�{E��&��~o�1���VI7�)Q��2䅰c�y�mO�){����BAIP!�AK)�3@�C?�W'��w�S����D��[�+J�ʋ�C�W5?e��\b6���*)���_�'D}O:���[�Oi�p���5:T=�31�5iy~��GTԍ��8�B��h4B�:\@��.Lѓ1O<�k[�e���Ŏn��C r�e�B9�9�>�:�_܆�c�R�-"/l�9L<�=�;;�3��&����"K��^�;�rf)0�K�����t$R&�`Il����-��QFlI�K�lu*���)��\��[�ua�	�h5�GM��rr�"?{�@�����\�#:N��2�N�_ԋ�,C���=J�5������<υ�$��ѵ��S��JA��_M���
�^9CB�2ǣw�,"]}�v�s��Kb����,RZjU���,s��+���87>\{*�	��(��dEy�����e�N�m%⿥��*3n@�L�87I6�����oϒ���;�op��e�����r���C��N�9��MrCO(�|�wc��ѸRF���Xc6��Ϧ�֑�&v?����U6Tx�]̾D\h�/f=t7���@���R�ٍ�D�q߄�zM��y�w&��z.�#�|�x�����~������r5j�y��B�����U��c>�a�����@ Mi�,��V0p���¯�k�S*�u\�kouu�cq��D��D Da[�7�Ǔ�+y
G�D
��4�=@a���13��A�鍘8�o��Gf�t$\�s$`���-��T�Iuof,�̛��w�0Ee�`�jO� �������A�9�~˥G��"s��Kf�+7i��+��Y�z�6,�aPX�B)�d�qЄ\H�V�r�&�һ�<�b؇��:�m�����=�v�+��_��!}i�u�9Ƿn^���ƄV�9ꈟ6r�QWL�8��7�qc#��Ub��9T�,����x�T����r���(ᦗ��|�KۜXC�l &��}���"ʒUD�y�4�ӱ�.�rZ�/;`o��(�H
f�>�ٝ<y���8p���?���Ĭ�:.�?��^ɷy�|�OT�[�pH�RN��C}����(]<l�",�#���	��O���B��ȣ���?��U�oG���1r�%I�U�AHEBMЪ��W��Ҡ�jҏ�꬟Օ1O�S��pdWJL%�)���ONV�@Z�g�ۥ+F&��)�"��!݅%ߥׯ�a���+ ���)��a����\j�7)r��V/pH�EN��3U�a�Iq?�)͏�m���{�W	�e�!�Ž��6r{pX\��W�5�ܨs�G�8���Y�̄����6�M[����5G�j)a7V<c	4�+�RU�;���;���T�}j�>�k�B�#�����:{�~��%^���{�[+
C���w����0g�a:�^&�o!B�D|<�4�e�/#sb��y9׫��|]��R�%1���6>���=$g���p&Mz���OlR����w�}:^d��\�9|�}=]ݓh�N. S>�5�׸�/�h�O�-��	�2r	��t-��	CF�KB��s��P*�!,f�\�6(b�vj��F9��XWs���4�B5�J|�V�Q��Cȵ.�^L
���+�'�6rP���)�V��'up���E4��R9���*�o�Ry%d	cCJ3��*��T�`��
e��	����O��`�EC��c�n�����p����gKˏ�7��"8��h���_�\Y�������T��[K�pͨ؜�)^T<����@F��vq��a�o F���o��e�e\Uo�s� ��)}�xA6�˸��dMcR����T�
$$�ͤ�?#���vn��#P���$a1�sF������8\X�^^T\Yiw�|5˦s{�D��۵�lD!�:k N��b��&#��74�{�d��u����O��:�R�;ܜ�e9�	��d�G����a&Y)�נ�m�;�%<N�>��%l�!�[���Y��X�o癕Rjt��ܬ���j0�M��p�M�b��{�ܟLH���
3����z&bΥ�(�;3�S}@c��Ċ��D{�} =�v8�p �ݘ[�}hӤ�un�\���׃�Qϑ�)#Ї�'�Xe� �t�Nc������9:�@�Q�sgT����6��2w����H�������eb��l̟пP���92K�X�e�_����|��Fޕ�$l�̜�{(*�]�`�J�+*�cƗ���ʛcT��V�x�|��1��t�Dv��:�}��������?Pof� ��� ���$3�Ʈ���eDG��u�����&�rϑ�:ֽ���6�}�L��i��~t%�H�(x}T>�oHN���M:9堂�\���̉�ϟ��DttB)�}��}y��0��*d��K�yQMk���glƉ�Y9�1�`tL>��$"p(0* �K��M�֑�0��vp�L:���<�^�'U6h��n����A���֘��O��-��HJ���i��o0:$l��i�=2��ɴ�z�нN9��dˈH����9�5������˘_�d�7U�y�B��}~rr��Z�r'V�'�����s�A@�5vbb\����N/���G5�i�ֆ��'��Y=�"��ϖ���6���E�" Ɠ��
��]u���CD��r0�F����둁�F��k��27?)즍��[z�>�{vq��v�*iX�
� s��� �4ZY���WW���C�	���)V�.�*�����m��߽�i)cD���N�5=�gx����)��B&�?pe+�>���⥮����y�&����RZK�:g<ʡ�N+J��?���LV�j�x�SE��{ܚ�(���c�4���A�u�e�^~\�C}�#ȫ��a`��v@-l� 4�v|�m��+W��p��F�FRNQ$�	u\��y��o13�>�ۈ��_�!���rc�W���������� ��S1�������-2�r��31�� �`�о���}ܜ�޻�D�"r�ev3�EL�Ջ}��o��'���^@p}s:d�������ٔ!*�5h��ȯ�ժ:���f��:�v��]G���F��$}m�$[���ڇM_���DP��	�pJ�
3�r·f1�+t ޲�#�iI�t8L��]����Oҙ ?��L�@$�w���/
߉�i.��X wt��4� g�lN�Vm�\AY��/��
�»펄�]�+5�c�v춠��߸o3[-�3�{�uC�,SVP��O����Ǎp�/��V��ψF������"<�r)�d�a7�ひ���!i�d�����c��zk��to�9a�ށ���1\�! 3�kw��B�-�#B*\���tri�Qà��l�lsZ.c'�=p�Bn�5�7b�x�}(�b{-�~�?����,�5���C�2~�2�R�(x6�R�~���¼I���*x �a!���;���eZъ��ƸZ�/���Gb
F;��Z���kx��&�e�;KϘD�' :9�[$#^+Ч�Mz'׳�B�CO�ج�B�|d�#�� �������>HZ�.u����)4%��w1k��TM it]e�Sl���4ӭ����Y��/b4p�=��4fv����Q��#"U;��_&��MV��LȞ�l�끔�4�	��{Q%v)���~P����n(۽����H�wZ�X��6���5�&�G�g��'pCڶ�d��Xe��	�!Sm���s�ˑmuO3��Ck�!�ľ��~�F�2�)�a���v�Ē���y��&��7P�=�@�;\��g�s<���D`��g*?����Z/>�HHi��_94A��J,������'5#F΀��1:jKK�s��=F 7(N7'��g�g��B�.�O9���@��9�9�1tH�k?�>�6c��� ��F���8�0�ԖI�����&#���G"wQ˲k>�sF����d�r8��L�ݢ��׾K���|W��M���wu�(�{ů�����tI�YvgGm�|Z#����O��nF�xs���!�"5�I*�붙�K��m�5l�<;�� e�vLd~����[�\�AWxǀ�w!���ZH���1B�,��;�^-�^��7⭟8������f"�cT���v&bxX�Ú�CiO�������ǰX�<7v%ˬCka���'��!�4C��+#
mndM�;����kА���#|��kr%7	'sb�Mpe/��5Ee�����@��)\1�$�%kb\W�\-�,D���[�=�|�>Η �z�>��]0Z#���$�I���	Lb!am�M+|�'@�U�D����ɑ.Y{:M���k�ĝ�4�@�� �o�m��b�!a)��䎻�~P	�z8;� w���b�*�z�>Q�I��b\`	�n�]����t��'g��f��� nÜRΠ��8�:.5�y>�G�|\��W��-ݿ`�}͘����m_��q�y1S��'&�|����'��
Qm��"���?�n���s�m��$x��$ȓ�琌8䑴��,�{|>��#n����(+�;�/�Yk�[ٿ	UT2[�O�2�=\L7}��%n�vFkg�4�?� V�o�K�ʑ?Q��]�Ҕ�K%� �k'=_���XGB��]�29�M�� ��#�G��ut��;������n8}Uu�E`�:�U�Hgd'�ޣ����O�� �"_t���jb�j�o�f���̵��K{��n��X�&��\K�[}�Vz��)B��;S�C��!D\���zY�%#�!�����&[�a��jZ*�2S`#'ԣ�n⏒>�b/�lx4�����A����WPϯ��Ƭ..��Ew�S�ö��8#2�;�`�7�Gp��h:�K����g��w��xnu�f�똼S�y�=��5���N���}JX����
�h�{�q���-�tR�V%~�T �f󯱌�Ȗ�$�\fY�_���n�T�p�}�T�^X�ӿ���zL��@�����$w�*$ٞ$��f���)�ķF�qɋj6��"|���9x`�_��yQjO��
���v;�H���o��9��{V�������lw����*���1\�p�hyM�(h�m��0�H� �~I��|����7<�O*�t��ސD�M�:Q���Ǆ�B�vG��k��%��E�(i�o���e=��(Um>�Jx����i�?�`�����~,ތȻ���^I��٭�K`��o]���jR�F�n*%\,��!%U�2�t��Al��3�5�у�@���to�+��N���e�����x�B�R�b�[®E�+�'�^b:5�ێ���-�}taCG'��h2U���dr7"jm��Q�˅�U�S(����8Cv��6�A��yw��]K��١N�=����쑏/��V�L�ٿ:^^)(��؏
���̪���CPZ���k�?��h������ȮBIR���z�N!��)j�}��B��ﻙ��AO$��-�PT[�Ə��3,���� ����"~�{�FX�}Ω�ɫt�l�8��qG��lt �!�r�R��Ϻ.��zf|��gh��-��,�ڄ	z�z��SQ�����W*��2�TץQ��F���ug��cz	��N��;�~��~���$�+�s!μ&��B��u���G��j�7B�V\�<���_5�P`,�6Y��m��CS����+�����(X�m�*�����XJH1�D�VX1*i���?�����Vug<���P�DWq�k�����B,����ѽE� �C������D�|���)�j�c�Jb�I!v����NA^��A3���-wS>TzkC��N������%�lm!C#v��̮�Y�U��j-�J�a~p{��M�e勬7�D��T���^��ߴ����d���d�ղD�]*�K��r�g;��*[`4�#�=T5��ጹ�~�T�Q�4~啾�|�\M��}.R�-�CPLA�Ǝ_^o#��Ua�,(����#\W��C�Q|�ģ1OR�{�ɖjX����:�Τ=��'���@`��^�J��2.Q`��	���g�խ��
���4|�H��ĵ.>J�߼�$6��#�::�d���4�W$^i+�W��z��������5��b���g�HO4�-�iG�O&"��UuMR6_ ��c��LOtw(����oxDƷ[n�*���a!;��x;d���p)���v7�Ve�V��Q\�b�c"���fU�{���n��0-m�wl�&]�Mm4Q�n�}*$��*/a�#��3a�y�e�~>�Z3r ��#& �d˃zKL)�cCl�]yϏG�l��~�s��w[|67(8 D=�xEC�mo ��Rz��F�dM8�8�D1R������-�q�%d$�g!�Σ�f$ 9�
F����AP���Sdˢdl�c�;Q2oŬ��Zq�	T�Ld�P�`M]t�w�LSޗ�'�\g-B1hw%n�:T��ν3[&�A*����ss,@%Ԡ�Ң��(���o��	��=��	�ͽ��G�}�'�
2�@��HO����S������r ��ܬ���ZT�ު}�W�#�����f
�HZ	�9܍:-(1
`��$�\R�<��L%N����!�&|�wfu�x���]���L�G����R3g�����$ak�
&o��QhS�m2�5*�J<��@X/�A���_����G}D!��?�����bDU0��9�5���@�h�x�����c`�I{U9�c>��,�hoc�ۖ�
p�&������S��A���ء@|'� }C�������a�6���r a���_S���Y���)�ƚ~]��#��C6���q������b/2Ru#�ĝ?y²p7����g�R�O�%h�ߧ�f��u��M�ґ�-b�5�:��@譚��Җ��� g?��ąvKB� ��iܓPrDy����#���f�tw�� ����"�y�� *6�|1Pq�dsޢ]TR�y]hk�*m>�����h�-�3��/�G� ����q��	LJ�hh4/�L@֗3ܹإ\!��Cj�NO30[��vp`���K���ې]��|���n�&��pevz��L�2��zV?��"�'*�V[�Xռ��$O����xX�&+��*a��°wZ4���r�큇vY*��{'i@�qT�z������ǡ�6��G��;Z�PKN*��'H��`�{3�{uf�agk�+�	Y 2*[^$5'�]�%q�c��*���2�=��a�W�}�l�ֹ[�q����_M���q�Eۜ�il�P���d�n��(6Ӥx�+�e2xG	��p�Y6SM�ϋ-�E�A����X٫�2A�n �-����O�����~]N{�;|���j������o=�'rƦ�r��D�ns{�T�$ф��ӓ�\�i�.l�g�j�h5��Ep&P�l���}���f@!�qZ�]܂���!}�ms,����6K�@��}�:9�M���4Z���� ӫ5p�R�O�V��7L$���<�ΗƎ���'���G+���L�yrV�4�����I����{{�<��݋(T2�^���K�|��8��|}n>��]y��Ӊd(S��m�$D�z��K��+�;�잲7�r��"m��Q�Y���1Z�~"9�z���Ωs����l��:5`����|�B��yj"��U�������>��4lw�M��9[���ߠ쒽_z�%��Q�P��ucge�0�cf_�/�� A=�l2�'�&<uz�[�ّǁ..���N�Yst���L�t��h�%	���������S��j
9�2
T#~�G���Y�E\n�	&�iA_�0W������2ϱ+��>��h-�ȁ��7�'?XhX<j�豿�K>�B�=�Y�A*�}�I��z�B�.Qka������Q w0h�W�3���XK�[3�I�}���3����9��㜥	���;d�
��f'$j_�os2D�j��V�`�����W��R�jߋe��M����ab�� 
�sxތ�"����*�q��n�j�%{�8����	Iz�YA�0M��]Bϰ��u���P��Y�=�3�9E���6�����Vp@
���%�X�w�ұ�3�L�c�A�޳	m�������&x��n��&>J�*��4Bo�_W�^�VH~Vg#�,�b�>aIH�M7ŀ?ci�����&_ �<��u�4q�y�\�,��9}��VT�%lwk���?+hav��-���V*^�SbM"z��((p����a�R�:�x���`LA_��O�Ώ��q�=�����F�m�������C󋧝8"��A�ᄎ����A[+B�Xs��~��Ƃ�r�7l{u��81�H������ڣ�K�dwy/M�Q�
J��Z&�侁���ꈗS#�����R��l=`��w@++r/_Ͻ�7���3�a��=�E�)�~i0�~�K�Ki7&H�U��ߤ[M^�阑Hr�α�(aZ>�
�%��2��m.=!-I�� ��mN`�R�YF�czuS ��� r,����4/�*����X̫��{m�j������n�/�Ji¡�
<l��W��̮3��P�䊎u�w���`V��c��D��FƟ���º��v������x�F��O	��wD��I�i���(��Tz�d_��8t��;�,h߁Ai�O**?B]�(���gA�G�"��PK�J�}�G���%��h�f1"�jV]}-ͺ���ڷ��(�~o�ɇ/o�?,�*����c�3?0nU�a����G�N��ŏ����0l��g�3�M��*�E����C}���]�O��FK�'��٥��_�r��~@�6P?(�����Q"S�M���E�v�O���mc���^�t�)�Ճ~��/ri�-;�f3��
ӳ�}cx�s	��J$��Js�n
�~e��s)���IPm��[i�E�FX�Q��/c�F�I�2R��޺ҋr�2Bde��ei���3Qz4�>��tʶ��hkK)j�����Ђ���GH)��4=S�1�ɀljxP��ft&���_�[aG�i+zoA��(a�l��0`��2�18&��ʢ.��&�=@���w�Ǎ�m��[^��ŃE��W��)�O�n�2l=�����p�acbPc��o��칽��'�H"%&���oy�j�O�b�xv�0�����$]&5$��XiU��/Th�Ex���^����A���м�M�E�u�h�-?��0�@�}�s��9��[y���+���TqTPu]wC��Y}�@g���:�d̫w\�vi�k��^0�������j:[<>	s9�qQ3^L)F;cl����R$n8�����䥺0�ʢ�o�SP�)��&V�>�ߌܨ�n|��~v�ԗ�h�\�(�,�=���R\�ߺ��t�O���0lq��t�;}�E�8^r��-�}_�5v!�!��qHy�����lY��XI��S���I8}��r�3��T���^�������#�����+�v���b�Bn�H�?hS����Gp{l��{���� H����	\`[�.�!���#� �����-$LY&aX5����C7���� !C���_Ҙ?o�ݘ�%5�<k����9�G�]��բ�������Y1�Yt+B���A��k�1\ϫ�T`����Gb[U3]a��fG��AܶA������a/X�6-��^�ƶc�%N�g�r��/��Bv^ ��az3G"̅�ӥ�����)l1��'�華kt�~ب/�ce�9v]&���ӫϸ��h����!��E�rYK���4�#"b\% ��f�^�z銙�R��y�}�#����<r�kչ��5l����k�=��Q��V}*�p5�t�#�A@��e�*��������0�Z�;8"�vm%�u)ޓ�uOָ�Ĕ����TeT�+Ϲ�Xħ߿�]��B]q���Hb�+��B�� ��w�~���Us�[�cvj�)�i0��2���cxN�bP]+���x�Ze���ߠ7�O����l�6�����|��D��s�~�i�U+mr6�q��\~@���Eq��2ё�
8�o�iS~)*�<����%lC��s���B�{Ç�sb���$�2$C�Z�(�+*����:��Gc�: �=+䆚���� ���������q��㩃E��'o�6�L�1�ˡ�*���$/������K.�5E��$b1��M�{� �r���F�v2�A-�Q:�p08?Y���ln:펉�aѤ���@���8rꄓL��a����h�����3n&Sbs������v��8���	�NVmi��WG~��] ��e�EQy�F����vG���Vy��И��|/�9X�u,����
���d��q�D�͒�.�F����8�r}�1Ad��mL � �Y� [��s�p`{�R �'�m5vZ��<6=`T� 7?�k��WC�ӫ�6���?~�?�}�Rī����	!���]�
n����ܒ Ft�l0f�~5c�׭�Mc3Og�s�����������I̍ɲ���%ԵW{U!C���O[Z�b�;���߅fS�u�c�a8�޶r���I��8���öP3oaP���	�p���%�Э�%��Hq��l��p� E͙?��z��2E��:\��Eܩ��.�D9��"��@��_��E��X��쮬���N_�y3��P�DYD��I�A�OϺ����d�|������wc+�`c���UҀ0��S���P�
�.U����i���./t�����Kb�	�Qm��C�$-p w2��_�FE�;�?ڌB���Zd�h6Nw�h��tv+?���!����h2w�����N�PS�6�k�\W`ki��}���<<����5�6|�q4��Ƕ��8�#*:Ĭ3�j;�n݊�e���T D�
��d��s-]z%C���Mx�<Ć[�~C@�)����@^^Bo̰B�K�`��!�ק��oY�ӄ�������n^Q���~��/���\(q܄���Ҳ���u�d�Mİ�Z1u��0yPj�"�3r9`~����XP�J$���I\!J�.��/�����b��ya�W˳,g]�4�ݍ�yw �IV���$���O��C�\e��-��Ε��,��
 L|jT��®WEN��Ѳ���Jg�֒Es0BA�x�%B��5@w_�2O���f�Gg���5�I�i��`#k�;&sp�)C`��;����\��������]=�n�%�䶐۶���E���Fq�̚#ӷ"ղ�9M�툋v���b*��cDsS�H���	8��zsy���k�C�C���Fa6ɔ�)-r����H��]X43�O�*toc��U�1aѡC��l+Yݓ�%֮È��G��%|z&�������[��:���7W�W�З�4%b�Lvº�%��i��ϡu[H�I����f"��wVW���siV4��=�b���M	l�uE���۪j[!�|9�I0{+#�j;T�ۦ)�"��.��L$D.��ؤ.����w�%�O��~n������J4���WK�\�"�����ѻ/��t��>�[�XUj޳�V�[���tK9{�i܂�c��A�ܣ\��	~�����FHG.���8�uj38/+B��'}-6p8W�"K9���Z'��h�{�~�jp�~TB�S��Z�/�c�C�b�)���9�c �|A���˶��s렠/�2�,�+R�W>��!$DR��Y��:��Ou#p*��8�q��F$g��]>D�Z�T4�J���~}�^�	½]s�0�x} �ix��O	��D3�4:}�0�d��\D���	���3��"����AŢ��+�����o��Ivm
����o�w0}����אZ��/Y�C,�˞TZc�95�-���� z��ڟm~�J澾��Č��ː3���Q��x��;́�N�H�Lr�Z�R��į$��@�g,�0��DY&�a�m�ow3�
*I���<�8�|�s<n�%��)3,bF��/jv�w�LT��HLʋ�*��W�Y-�x��}[����xT!�c���	cv�>�y�KߜaB�V�������g�$~J���n�3��0-K��ceM�!���M?�N���cT��o4�02{��,�aⴸ�j��0]��`��}����K��18��"~{W�"14֏���T̝\`�Q	��Ic�Q7�a�����~`���#'����� �#A�Gexvɒg��o&>|�՟e�U��x�� #�x'�*X�s>M����p9���u�Z	n�P����Э�C���SFӷk}��gjǕ��ij?h��u1�����H��<�0
�	��|$�^��ܧQ�3�Ǵb�(Pf-�負Pn:��~fo�u�Jt1�"��w�T��4�J$��`����$�O��/�>�o�
���kI6�4�c�Ô��<��_KHZ��ܝWu%	-�ic����~h��S��N�K7�ۖ�cN:Fy!�E?��d�3�A̮)[�j�BC�#ݽ�d�@�8��[�|��i!�&��L�M�R������_��g�O��Db�2�����C���&���Ea��8:�	<1)|K?��!�[�N��|}k3E�w���+��"A�I).<�dM�6���N�,��sw�]l�-!zc�O�Jޒ�,�3���\�2��+X�bRP�Y��#3�w\+N<p���d�	j`���N5zĜ���6%˻àa�{7��½��sl����3m�<��$���SH�b�x@�I�Z s­|��Z$�fm[J�U�Э+BVOw۸O��)q��GxY��F1|���y�>, �����,��z[:�nb��)�g�K�K����#���(�#�[����oaX���)�ѿxw�������a�Q��4��t뗩IB��+!Rٍ�Wr�.�Q�sJ"	�^���P����I�_y{����b ��L-.�g.(�41��"nl�t�z"Y� ��G��WLOT.�/�6[K1z��Lt-�|����w�z��i�� =�uI��I6��n[+w��M&��ݬ��Ŕi�ND8�5+��Y]�~Hm����3�� ���z]��u����mXڏ~CI�?���븲��&�i�G/��|.5�}�����( /����Uv��E)�a�tT�4~"��O��g��@��䡄�g�z��K�}V��{�1����N8"襖�i�x�E��!�����jߤ7���o���^fI��km=�F��B�jo��q��S��1�'�y����?�� c�/y�l.yTI�������F�d�����x����1�J
���;�i;�����	}��НK�*��;�,�r�d�����Ax�r��%<T\����:s�a�2��pT	�MV������I�M��oRk�ȱqR����i���~�q������<b�O�Yr������%1Ml�&���-�}�V"���6o��v8n�G��Ұ65�W��d�G5ջ�ag��}.~ޮÓ��י�-ϭ�#j<�GY����LXc�?O���jv��dU�2lk5��0�^ $�7�5�aw'^���m����b)���:<!Tł!�j"��U���U�N'����Ј�ڣ�NOA�Y�Q2)�gv��4Z�x�JM bȴ� r,0��3e��uL��;��-���� p;�V_�s�&���3N�U}q&YiG�ꖻM��#���E�ן�8+h�R(��H�f��A�/=�������!�9���I ��>�� >	�H,U��h�fM�Xx�"+�>�G��w��'�N��&(�0�Q�
��p��V��C�x�s!�����g~��#E��<pӆ(�L�F��NdF�rky!`14u}!i����j����7�<�8�j���{Xto|�$�%��.�*L��w�M;	�N��w�5�A�Qć�e��.Y��D�рr�W�`���C"�p���1k������_�����M!l�>�*��ܙ3#�?���X8j�j!QS�U÷�p�gyY���DX���iI�=a>|`�uNA����&k�㈍�ֿ��k���U��9	�~ѥ,��4���?ˑ��� 4e5��+���9�ny the�̓�s
�%���c�BWQ9[&3��C/��7ah�f�K�����Ge�;خ�iS�BP_��F��Oɬ��o�>*{5�	��Cz��D�tMF���!!�J�Ă���tl�j����!��%���.�p7h�o1�U=�?�R7%�/���3���;`�U��hΟ���M����nP[�� -2^ �~W}��huJ����K�B��\
ŋ"�z
�kk��oo^��⃷�p�3���:�So�$�a�ǅ�V�vr�-�t�u˻���ga�lͿie�TRU��/� C�)w؈����T�[��$!�c`��9N����9�w��8;�#���L�ؖӐ�t�1N _�b���ti0
^����֭=���6/q��̵�;\S.�y}��&X�B�:�A�|<+Mκ���+��}o���a�j��Rh��"�{�&к���[���rt`���崕���m5Po���M�y�v��u[���q�.�t��&RaX��3bȺ%�z�);Ǘ��F4	���CXN�y���	K$�ń������Y�b�G��#,w���m��5�6u0dL�^��Ӗ�W2����I�03q)���A���b�q����j��M����b��_U���.,8ߚ��o�k�)r���B�o�x]`�ЎϜW��M>"L!QZ�L�&�k$Ϯ.����{�6�1���p�HZ�~�W>z����pVغh7�۞y�Qj?n&�Y%���	�	����_�E'�b^���n��&7f����r�G��"�9�]6Ɯx88�:Pdď�+��� ���1\8*qg�>ǖ��bfoS����E�ʶ���;�trx)mi%w�8�&y�O֥\��C׳[����/O\@4ee%��մ� ���o�6��r'�BD`�w�A��@I�G�R?�PrR�9��H��bD�&�d�����$?�/�z�5ڝ��A�� ����3��~��#��*@��ձ�;����Z�p��E�O�>���R�B����G�h���Cu!�D"7�t֗�HE6�k=U�m���4��=M䏝*�`��E�z;$�w�.����#2��X��f.;���$s�����2p���l��/N�;�:927ItRH
G�fIv|g�;?�d��1Q\�Ɗn,�M��o1X��h��
/�����Հgz{
t�,�i��[`j�!�g��n�Z�U��W�l��T����d��)_k�b��A�����-����֙�^h��T��>:`�4:���&uf�D࠴<4e;N��b��rq^6f��ܑ��l��<�h���:�8�2@Y��j���^m�� �։�o� 8�+H0�x�9)��f����	Z�e�ȇ���vqW�|����[��Dܠ�"�`zK�mv�=x4R�r���^���Zܯ\��ԣ(%����4���2�ܐ�0;�z�pk���]�~v7�$�ցƥ0k�n����D��܊`�Y����7�zי8��  2<=�):]�c.�.��EBHhe�{fr���Y��{��AfG�	�+M�5Ƌ&A�ҷ�CAKe��U�����Ύ�$�v�y���L�L:��}{W2ί������Dp9"j���j���
��-92(E	�x�$�l
�W�Z�u�S�m���j�GSYUtS܎�jRoPo�G���лF7��B]�9v��W��|h�/,�?����\S�OA~�{Y��{.�j[襞^aG>=!K����%N!k��댏_5&̾:K=���N�X����m}�N���)�Ա��&iV=��y5X�{^Z���BŦ�N�����%�h�����
����Kci�C̍tA�D̀�6ىZ6ۺ�nɦ
�����*���O�����j����g��n8�hrr���X�
Tj@�T�B�)��CW�:jC�}�/�m��`���I���ٳ�|���7n���:���H]B��>|�gS�>�
0ż��m�������䬀�y�f���p�!*�g\K�=�D�W�[!��|���������A��Ǉ��� ��]P���^�ж8�fK����FDz�z-��[����S�����f�*�|�ȼy�</��T�]��;z��ڜ=�c ���lGns��z�~��^�1�4=o�k��� a�fA�	{!{"`��`�<h�mt,���à����89؏>�ހ'<�6��|�����H��o�~�F5Z,�]�����9�RFsg����������eܑ�z; U�D�3%$fr�n�\�p��\Q��n�-h��:5�حg p�ՙ��C,F5��Hi㽎�©�T"H/;�!�����.��I����S:�"}ʠ��Rw�|��{a1ֲ����&bu���}����w9-�8�U�j�Y�&/ʵ����Up��v�N)���rKD2<��>^S\�e���gW(
�d��\�y��}�Q=��)F?PY���խM9�-����݉��N����f��;��C��Na!���
���Ш��<UXh<*(�|r��f�u�Dу5���~�3�u[uH��$4�����(�Ds�	,A�T��~��73�6&$�嫁�W�N40�ILi��O#���Љ��lO��
�)�	�S0Np��0o�Zl/���J�C��0�'k">]��h�G̚\��-EV��yw�`��*�s�Y��l��4�D�l�O[��5���5[�=�Ys�Tm�����g3�47���5{����o@w6-��F>���L��Ҝ(Ѧ3����q��e�.��f����"�&�4ۄ����zFl�i?���9��H��i�y��.���@��qP$�n:���ꜝo�*5�1�f1dO�؀�a� �� ���~�d��>/��ƚ�^#SG��'di���zM����/�}��%�q�S�ޫ�۟��64�QΞ0}�|1B�찊4U*��*��Ūu�� ��ذ�HjOF�Ϋ-<����E9��{u��mE��7��v.z{�?�COB@�O�e�m{ru���:f���*e�i�'ڞ�� ��XC�aȯX�;o�k��D2���5��420��h��]i�p�;W%�ul��*��
��K���Ol�8�c�kxc�(a`'�v,�j�!�y&�K��� 8�֝z���c�w-�\2I_ק�����0��t����"��N�y^�;�W�t�j'>A �.��/ZW\�iORΦ�u���;ᘻ8�����N4�Մh��_ǲ}6��Q����ณ�q�8n����+�QO�c�87���4;[�F{\�.�-�R	��g�<��؄�8|Ƣ������'����w�Tߡ�daܧ�75K2g:��Bf���R�qX�M����k��B�g9A��6���59���q,��)Ϭ�7�@��7�38A���c+��$�N,�ɫ=�1H4N�!6�H>@M�r���8�d��co����6�θ�����*t:,�EbMNu�P�J�6�±w���S�HQU 1P<9����X5���>��D��=v� ��2V?V��}���&d/����������u^�cr�&	;�!\�Ԑ^Ղ� � Z,{�[�d_��
VϜ�j���Qp/l쏝�8��"ἱ�7�4j�:���Č�%MWq��nLP����Zz�/=#�}h�2� �!���K��Q�s�=�WX[yx�}H��_ �j��>�*E2)k���������:f����9�Q�53�9�m�X3l�a�2mD�@r{VJ.��%�����	���ϰ������`�8i����"�;���)�G_�WՠJO�H�Є|S.�o�A�n�Ry&��)PF��r%���H2��旰� ȝ�+���x�F�L?�+r;*�\2��j?bfqALF�v����* ��F��V5���"��������.���©}j�>58F(o���({ĠE �S�6\S�a�2P�`jC��i��$��!�9��E֖��a=iz�j��1��I[�r�|���MI�<"��7F.#����/�ɫ"�[�+��:��>���4p�|c�61�����I� =�XS��"��]J�����mRZ�����^z�o�m�l�Q`�ǧ��'����)'Oѐ,����}�ηX�� �3��f�I�����AP�T%�Π�cocoz�o.���aYX�:N�ˇUy���ڞd�ظ���e�`��� �yV�{�j�	��/�E�;'��H�wI�)E���g���J�vR�< BQ��<w��|B��7p�}�}�b�~�E��d����)�]�R� 6%�$��*S�1��7>�9**_=p筭.fQ��=��E���3���$@����!{��-;8.o*�R�,?ċ�8��O)�Sī/�w��ۯ�j��,g��YF%<z{�eIt[�N&�~?�|�ES9v���(��I��Q�[U��b�+��كk�\`#�	��B��E�و��فe��@͟ �����CZ�z�"S�=ߒ�+�V����)-0��x�~�m� W	U�a����g�]��+�z��ʨ))�Q����;���X������iH�\D,��T�H�f=�Q�ߊD�Es�����"P�1Ua��YP���5�/8��\:�	�ɸ�A�K��Fi����ˮ}�����S+���_�{%�;���H�N����*�r���ql�����s>�W��{�oV{K�=
�?�$p?�c��62��V�\�D�<�0�����.��BMB�!E��ʦ��A%80l�0ʹ�S7<�ȄS�c��]��N��*��7�$TW�V'N�J�9���_��0L�i4�F��䚛��QW�!�-�~w��$=�C����V�R��ή�U��,M�vk$�/X�,c��r��u@bj
7&�﷕fO\.{�������kW{�=�k�t�B�������Ǘ �O�h���G�_0��,Z���ߝ!��2�,˾�W��@L��g	�Ŵ|����n��,:P��s;��M
��$���];�Fl�#���K�b��C�u����L�Pe�uh���Jb)D��ә's�s��[eX��8�6>��d.HF��s
��av��9DJ�Vc���T��L׷6J�k�+^�{�ʈ�7;���$<w��0<v��S�D&���:��\�B:�AK��]�+����]7@_������lQh���N�Md��y�f��؝��8NW�m���qo��=�������Q+��f�����U�e#��2����#ۭ�0RdG %��:0,3?��5-�������&���k��Z�*�9���b��H.p�6�/���FTW'�����{�nd���ըx�9/]`����-! ���.uy�@��5����w#C�u�i>n���I�C�Ri_`]WTe�+�zm���UI?����(_�"�pvsw'���f�� �v�1IT��	?M~N)<q������Js�
+7X����$jZ�y�K�X�kybA�c*ӝ���g�B�����鴔>������O��dA���c[���P���X�Q/Ю-O�������UA��1�\���Q����ɽA��������ͣ�������/�G�t=�J�~p+:W��}btU��_;
�,�Z�3k���E����X-�ql�������raj�s�-��o3VjT}�j"�e+9�{�ˌoLU	�˘���?������5ö�/fʞ�Ld�j�<]���f�fv6��{g���c,�p��ђ���@Adx��T�2p�LN]����x� �Co� f��on�K?�(�<ȯ��DؾrL��bfY����	T�`����[�i�<D��cW"O[�"��)����/��m<�J��E�s��G�������K=�W/���Ng^B
2ݱ4��.M�;uT���f��)��MA/��:U�`�-��5Y�X�ʲV�ZW���,$J��F'���&H�d�B}�_�qR���깾�6�M�Ü\�x���k��Y����V�C�w�Y��b�@Zj-�<+�)�d5�{�V������NUe���S�}+d�z`�ov.���a�Y����d���]Խq/���`��
���<�+��Ӝ�&L.���X��U��w%L?A�l9�'�Έ��>'�QP�z.x��B�&��&�ʬ#ik�O~!ً�l	J���D�����b��a�Y�j_��<æ�~a%�bq�� ѳA�}�M�҄��z};������LR�&yx�z]�kk�Re�w�ż�b|EC�F��9@X�C�q���{Z'0�LM�KOJcf
,�����<�,ӟ�����ѕ���]얯1��[�=��<,?[B)��y�<{�k`]pL]�xc�"c��`fa"��~f����i$=�3)�^�=Q�u(9G>	��㼭���1wR�$=��ݠg�z�3}ؿ�8h%�m+��7��F7� D�>l���᳕D�&1DB򴍙�����`^6�B��(*���O��V�M�Э���b�& ;�7�ZW�(����(�w�q8�Cw��B�^"o��t[�ky�@S�B�>�{؆�*7�˞��/$J�����KG��t.����Ia��6���a	q�jȆ86ٽ{����4�'\��C��2>�-X?݀����>r������l���}h�u��τ!X;|:1Ȅ�b!8���TK�v�U�9*��ܻ��nՋft�U�q��'u��:jQ���d�[�f�߉v��ꔏЖ{j����Ӽ�@J���-�1�4x�n�P�]�͉2[�o.&�	tL���ڔ�Xe�$]�����KJ��>7�"Iok��5�b���'�W( x	��P�*8�Mg�]��>���e�vⓆ����(��j��g�?wg��~��RP��Q�u�H�1c�B'C}`Ჿ�ʤ�6g6�E��?�S�me�g�c�Xb��"�����ˡ���4����0Lb&Y�Xt���z�b��Ĳ�!/:6�	��I?�r y��~�2bY���rҺ�����v�����l�нz��ɍ�:eje��~�p4��1�o�L�A--$�i��-M���O�U�T����3۸�U�T�G��y�pBŤ.o�볆��D�6��$|L��+�c&�[n:̓��'�� :�]�;A3�����expb_��s#YS;�e�ʬ�_JSE��y!U^;9=߽阮����Pi��II��I�v��:Jt�CwC��@<�����J�^�����ä� ;��kH`r�Z�y!��
=� ��(�hڑ��H
�鏅��T�7������Ե��/�!�&��APOw1�C��V|Ev�,!x�:�d���K���t#:����[s-��˽W�?a~��5��M҂����c/�ɿo5��r|�~��<�ғ Ϲ��\D��Im�3AB<���w�$v�N\	�z�����W���&2�XEM�?z�F,�#�+i���i@�\��':���.��O­�t��.ߏ�R]&�'a�\kH�m93C���3�yA̆���<�1t@�$&Z�ʫ����i����G��+�x딃o�N�<Pm�ު����1�	l�b�w�#{�=�j����*I&�p�Ft���k�u��fu:����^ ���AC�=n��-Kl��l}R���r��p\Ȱ���h5�|@r��?n�`C�{#uN�Pc�b�cb��g��+��_��_��^;�gC�+h�� �+d��6���d�4+bT�����n`ӡ˴�c�|]1�`�[k~R���mIKo��mb��>k	2���sIO
���n���~L��#�)��bb�=Ȯ����V�is��ݟ�8{1��w���b�b�u;��C��1�Cj���u�C���J.�L�\�������9�������B��a�p�K���֌q��}�K���J*jS1Ki����Y�� S��9������$Ls*��S'�$q_��)@p�)���X(Se��f��Z��?�G5���x4yǨ���FX�wuV�|L�3�$���*T�;��v��o�:A���F�J����w��F�$s��ӝ�}�ҍݡ؇��N'�TzkA�@���t��s�~#j6[
�o���*���K�L�g:zБz�n�PS�3�ټr���M�+�����xO���\,�á_�$��$#���܂	�lR�����t�����h�c���w�=�v���K����'RL��v~����A]R��/[~J/�5�yz&��<�)��j��o��+p�a)GM��l�z�$9�3��u�C���M�v�7%��?`�o��H�6Ol��|*Y���f��_�|p������'�\6�x((0H��;L�$�E(���s���o��Ԁ (��@����Y[���]��jH�3�$���HH"���e𱅔p�!�;��W�BZ[_�u�s
��ٗq���I'hBZ�(!ƚ�M�Hx0���J�ĻL�l��)�*~�<�:)Ŏ9s&�(%�iN��2�m_*_A��?tL����(�M�o�u�<bݗѿ��ab���&8mk
$�B;5�!�ǁY/,+��9�@[���굮�X�p���&	z�0�h���ޤ��2�{6�{eT���Tu������������RنՕ����Z[��Z\��ם0��EB����������t2�2�Y�?��:ؤ�d*�;�q�P,	�M�H���",)=k^���6���h���,�gc����[�� 4�����ᔪ\�Z%��
���9D
;�=�_��j�8�n��R;�=�{3�ع��Grg���	�w��+�Z]��ǼKK]�&�h��S̉6��Zc$�>��)<C�#�t]�S�dml�{%�p5�:�4Y|bfg������2gW��s� �F��ڝ���p$�m�lf�H"��ώ�T��� ��/�`q�S�L]�&^�b0��������B��5���@�J!7Ѷ�wn-�N���N.�u@�-B�hs1n6#i��� K,BZ3T�C0c��۽F"/���H���I�#aHՊ� �-Ck��	�/��=�!#'+j�� �*��=X���ʵ.�{\=�b"�~_v���'IJ"'����v�q׸�h��G8+1����)�f;IG2����_��!�bR�'6:�P���#����Xz��yE%�ܽ[��f�����鳘2�V<��Ӛj|���Э_��|h3��C����&�Y����`�ןSq	e�˞�/V?�T*_����h��\�G2��h�GŇ�:��w�O�wߪ���1!�De7
܊)Y:z{�࿵�y�UF4��z5t$��)�f���o�@�J�mgS}fVC���LN�ਖ਼���:��O+ؚ^cFr��L i� �̑���lIF��D��&�)X%gc��s'�೏װ��X��V�_�x�����T��Vu	/��o���u�Z�׹�=I\�>Ho�-\6���5�vE�����g,l؉۲�$s]_	m��2[b� 0B.���m��
���̉���	����� |Na�E��P/6���S����{�j�R�5���
�\E���ZQ��,N1�`�/=��;S�	ً;�u'�>�q��4E�hd	�o�O�_��Q����D�N�a��:[3�!��ډ�e���������nF���u@�AϥB/c�>�ܒV���kA��BI������ǉ����bs��J,�B��Cz�K��6)9�g=�/m�\�\��ψ���|�d��̟����΁��f��kcrR���9��'I�ǝ�Vf�JvZ�CWc��yD���r�}�h&�uxr�x�E���ZZ܅��yJ?���ߦ�fY�^ա��9=pׯV�كͮ �4}�L�����Ћщ7����w��i?�b�$5`)?��A�r{��_{:�V�;���ƶL�}��`j���/ں2+��W�������kق҅�_�8�j|��w��?k�S�����r��p�$������Ԛ��SFp3�-F�/7���
��¼���mlX�2�,N������'�������%d�*����#�#l�{OR�F1�)p���e|�ydȮ�PC�$�5�}pU<�N&�h�_i�ҌRσ�묜�#L��E�r�FΙ���	���_�%������rz���B*V�)�n'���9]�B|��3�&��ɭ��}ÏNE�>���^k����]��@�*�w���瘂g���B���W��k�dHM�V@#�}6q�w�`S�<7�!��	�sm���B_KŃ��<��l�7<��$W���4�}&�x�*�n����V��1ߑ'ܷU�T� \�~C���]Gc�!��5��&�-:#ُ�}��C��ϣ�&�b��F��sȞ�41��ti���*�dh�R�p��y�`zYp�Dy�zZ<�Zdw�м�����H?>�K>�D_���-Ч�D᫕��n\H���ɽ�QX·oE6-}���T@�,���c�N�h�1oA��n҂�w���{S|��`b�z9�
�b1VܥQ��4K25'��9�fR�4T�bhZ�;��>d����;�eR�'j	���}���}Kx�i���ޒ�F�- �#w^�N���IF���������7>��7�[w�Ŗn�J�%_�e�i��3/�9ٚ�Ŭw۹ۄz�t��'��&U���{���L�ت��p�a�H��z��?�D��DW�-�a�0!�t��}-ί�u[F���F���ȡ24,���SX�o�����O:$�;K|e����W�����r�t��Ԇ$Xm>�Â��nE���-�N��X��r6�D�(�&�>J��YE)�$D^�{��R6��&Ƴ|�������"�}�ok'���w�iZM���.%Gm0�r�{5Et	f�/�&ܱj�Q�0��`���5��oݬȃ��������I/�����3���h�&9��G�'�9z��"�N�~Wg�=lY��
/��x�����}�;�O�u^uDI��;�Eبcm=�Z\�)N��NW��f�{��X�{��$Xc�1U̴:��i�Vs`�xĕ��]�N��/XS�Wf�d���6�bD�SV����Ö�t(��b��� �\�"@��q��&����xZ,�3����]h��J���1+�n�P؆^ZZ,�|���	��Y���0x-N/��H�^�1F�X��~(�q"Q),��YGX����ƃ_�O��E{��O�(���b��"�����?�R�!*턊J���8N��@@q
���!%�ZϏ�n����K��CO����6�"aB�S�Z{K�YmߑF���?{)�U��P�>��\��o�P��-)N��eV���S�*�-AH�SҚ�lHO�� ��׹��҃�]=ͽq�:��)���!�����;�?/k,q�{a�����ib��P��#K�Ogw8���������K��;u�1��[da}P��%1�)f2�-z�R7��_�F)V8���%7<��Ө�� ��p�yd�ܚ#�1жo0d�}����ɥ=�Wզ�p?ٱJ,��O���:a�O�	���?�^L 0bf׃>ܯ@�� 1!�\��Z�Ί=��&~���Ɇ-=p�$�
��Ŋ���o�����
D�����D#^�L/����9�N(X����p�)%a�<��%Q�� ?�H��*��,Ԭ<���@|�
� Ȁ�t�F?}�4��_"姵�t��#!c��K�|ˊ�
>��H�G�PuuJ�G��1�8�����5{�?�1��@��1=]����I �U�Z�[M��W��0����!׻�Q.�b�$E�A�^�]��ocFH�*�&��=�c�2I�T�{;�%K[�׷�2�,�Ð|ui���f9_���K�r�LBR���<�>o-�f)�c�
F9�3�b%���CW���Xu�����=�$���MGr ��Rc��9s��xIK�@7�2��'��8�#D�Jn��n1��	�G��Op�[/V ��8�r@�0�!4���IP�l̺��U��d

�Pۀ�?������Kh���E�� ME����&H�J���I�I�}��G�v���������k,�/;'�M7&�1�n	jk��|A�]�j�I�zw)�+hVR* L�G����14��*Yѯ/��>O^3-2#�V�|����uM��<�L	�_��{jQ��n�j���d�	S^�poI*������$"j���A;������1�if����Vm��%w������ȵ�\�N@���#� �8�����u����WX�1c���4�	`�����_EwF���uV=|�|��Ӳ�&@�uq�k{��Y�%<Z�����`T�/��Fے�#�[w�av���RI+��L:9��p��dxE�ߊ5���%e]|���$�	VwS�t��&��Ć�JkM��-)ٱ�=���J��/�˓��ț��:�w�?tMI��]�Ba��f��yˤ7e!�RBw�OfCxq�C~�/��/�t�{��O^�v4��ne8w�.�w�;�gH+]<�/xx��ob�D�89N���3G���+ ���cfŁ����u*�r�H��h�k`7�c��]~nQ�b2֐j,qʱ�����R�g����h��gs�:��c��L_��N
6��g��q���F�λ������4jS�6��D=��=�!Р>�z>nnQ���OXG,��S�K��Z+@�!A��5��l�wQ���Gb8���ezR�t���j�4�Ֆw.W��26���JX��S��F|yn>lg�M��*�K��m�vB)��R)_*���pf����/�>+ 8��D7��/�<:c��(41WZ�&U7�_D�M1 ��ְQ��"���$΁h�1�|������r<_:�'����C����,a��M�
86�[w�';���is��!��zz/�l�ޢ�H��_������~��^�J� ��[ՂF��Y�N�:~%^�8ON�ؙV8��.�ׅ�^��LIi�Q�7G�k�;�ޣ�署�푲pB�+�QPR�ݖ��ׄ�1~<)[�+#�k[eϣ�{�i���|F���	�e�./*���(�2�N�0,�W�E��ǡ~�a/ml&9dVr1�R0�/᫝Q��3��[[�5�h�:����j����A��RH�v/�s�j�F0�����Q!r#nD��Z�3����K5����u�h�b�Rګ3N�fR�AJ<�x�l�!D���섂��kD&jZ���/שּ�)@4Xi�q��d��Bb=�A�y>����l�⑳�'\�)U�d��6`^�]M�A����(�n}v6���L�8�PWu-��	N�F�x��<���O���Hꁜ�� (I�<#�~,��,���u�3\�xȓ��[������|�`�5�_�t���G��  ib0~~�=n�뱣��D2w�do�����8��)G���U��b�R�����?���hG߫>�7ۥ&������rx88ji
^X���gc3�{l�	���4��U��։yתaCC����綪�3����Ɖ���+f�4|a�Gns���(k�#S�&��g>�M�����^E~i=V?���.#�_6R��Nʛޥ1j�Ց��l���g�Il����h
��eāi�u�9K��FK�I�*qY�5��f�{��P�J�k�_�'T� e0�䟹s`�w�&v�i������lm؃G��:�b�J��og7��b3R��s������z�(#���e%�"9���h�$ۓH���|�ٖ�$й��!�����d���A���ւF���ŋ�~v�ؿՠ5��?�a�jb�S$�ڶ�[�MR ����KXg\�Xs/�ʖ����ׂ`T���� Z���&E�a=��!֢�����3y�����\א/T�0{!���AK�����Ƙ��*���.���c�� ���N���"�x;߾�C��:��~��#�3#��R_��Ȍ���0!XFu2?�?s|�b4DZ��0h�*ѹ�\�������)럁��g�����x�_(���$��'�3i��5H7�� k�E����j�#Y\ӟx��V���0����VR�bN��;��6B�n��F�j�Ѽ�E����5�A�\r��bxR� l�;��т��ӝeݦ���c"q�(��S�=?�iEc�������s��"<(�ۛ���g���4��mϏd�zqU�r��yq#��B4��uSJd��s$dx��<k[�Ԧ�q\���NhpU��~�!9�y�l��;U���������)��pV��K�o��K@0��fx�eG�����<����"�.�����!ܐ�ԅ�j������J�X��<b�v�{���y��,n$_���w	��_�)��g�w�ê�3��|���b.�?��'Y���D�bQ[98�7Py��)�l*�-��wE��Dg�f�,z�O�{!���NjM4�1ŭ��!�����u�GZ�6�.�� D��`��_�[�C�������⑵�O�+����O��8���.��[B��H]a����T�`�9.@��n�or��8-�د�0b�}�Lܢ�E3i�Qν�,oI�o��c'^��m�;H��s�H���&̭r���=��P�l�<ʾ�Q�P��<��Z��0��eڣ^�0h�Ƃ]���CMB���M�G��e>p�un*QY�'�$�c�.-�����uvE�'g�����'VZ,��M;�x��}be��v�ꪙ'��s�D��Į����.�պ0�V\����}R��V��}Q�ɓ��1���োr��Y�.E�#X�wv��-Xz	���)z�::��3�����aɸ���ig�Co*h�f�}�[IN4�Y�y^�9���6�k9�����{��Aqu	��!L����FT�EU��d�8�a0�ⷃگl�x�m����m���!���d�c��nUS�{#o�=��<e� }?�<Hc�r'+ R� '�H��&���I
���:� ^��N�G��4��z�������ʨ�|�$.VS�Ny����	���}}얷�񣊫;���>�s�)����߇B4-_�V`��֙� &6'C,�e�O�{��P����z�G�:�P�ʙ>r	J9/F��jN���1��*�K�����l[	$aC^�lZU{�{�k�'��l�[��(K�U�;*�!�-%}�e�1\UKu26���0LA�3��w��E�{y��K:�[ě�e�iB}&<���<����Vn����&�UG8���a�uH>�Ͼ{dnp�`[��処W�@bNƆ�Hx�A�,7%�U7�U
� mw1���4|���mR/K7�u�Vb5��E K��^Q�I���ydC��0�l���J�$�ꌃĉ1E9/˄���A�z]������'� �s���y�kӧ_��⸿����rb�h�L$��|��jp+̈d"t(���#�������j>��b������cNB�FV�LT�����������w�-Z1
tē�wܯ_ĴjEJ���4����p�����p��[	�P���X����
�zO�9���Fǔ߿�bS0�%lUH>��M�5�MG���� ����>�c�4�"9��� ������8K��6d�4&h�~(�w��"�$T����IE��O���Z܁��fsa��oe�%3��Hz�����*' �Nǡ��U2%���E_ [�E���՘�����u���X��H��y�Z�`o�"���/_�*�kGq�f�G��Q��̰ה�G�gs,0ri��e�w!6���32��Q��&8��C��e�̅�>�zd9�VQWf[\��^�5���߮�
lI���'њ����Y/X,UI��P�|�<d�<���DG0<�6kmk�TUj~o���0�����N=P��o#I!@,5���E�u��@VzO�ڢ��]�Q� ����F�٪�>����<�Zۿnnj�g�H#ȝJ2%]�Ba�
�o����Ռ��9����0�#�\�~\��/��K�V��~'h���滃�i���4\県�����I[���:����g���MȐ�T�����<�k{Iߟ��>��'0��`?��oc�y���"���v�3G5$v�5v���U��ֵ�:b��lTJoG}�G&U�����z�����z�3��� �+���PC�uԒ{ ܟ-T������x�J^��g��f	�Yz)k�"���bƭ�!�x�ltEy���\>�k�_���H��
C`�XA��"�T9\d��%p$� ey�+��y��\����,��[%T�#^ǖrb���P&�PY(SjtmU��;refe1͡����fBG��r#t\�Bg�k�[��l�q��3 ����Z��,�.�@Ox�o=�m -2z��A���0�}]I�{�4c]����T���/7k�Ϯ)S?�ƽ���e�.}�*�8?NLg:�<ۏ��Jg�e@�fp��ނM�mV�R�1d��$�9���윌F���;9��y��C4	7G.�Q�b�uJ����,���;��@Z�ʵ$�V||)�$�_m��|U��՟ȷ��7����t8�]R�_y&ܱ�F���l��?
�1}Ґ��Y5�+y�^�*9��3N�)���$���J��w��!��c8��f|���YQ����ݙ4#��VT��!X!�����l���7组����ˠ���$��4lt<�'r��8���f��D7�p���ܯ���9{�;ߧ�c��CX��r�a��p�K)�Y�{Ή�+B� �w�r��}�����5<�Fe�O�څ���ˌW<�f+�}�|Lt��Jdd=-��Mb�� ��̓�=�2Y���B
�M{q�����Jx�(�o��K�~2��Sk2Zh���>x����,�{�+�;h<z�� �#�(?���Ĥ��_I�����^P�Gh?-�<1�DT*~�e/c���L��"���|��n�&��-��AöS������Y�*�t��*���:����f�<[Q鄶J���9�tl�PE�&F°�?Q������V���e��2��P���x��X8�+���r�X�=#��z"*Ʌ����rz�����sơ��-��$���)�� !?�0EX&�R�9<Ϧ�~"�BH����s���p'tH�S1-��M�co��j���)�İ�fr�"��ܥ ;�:@��n�F2�0C��[��<W�@6�ȏ?,�е�[Ș���u
nͱ�H�Qf��pb:����	"�-@��7�����e:o�o�p�޾�N��4�4�h(⬌4�x)uΆ�kL��;���f������L�Ɠ!���+�8u_t4v�d:��� ���4��ǺJ��#7�\"�>p������P�ӵ~�5#ﮌ{��9�U�C�Ʈ^���3��艢x�C"���v1Ȗ��у�"j~�Y���̺|����:�ݜ��{Lૢ�"�zLn����{Y�bh�*Tр���
է9��#���n\oJ�7(��0�
V�X�;Hԃ�9�Њ�A�ƻbHv��|��~�E����-"m����ݱaVF�8��=�K��?���lq�61�C+俎M�~+
y*��锐�Kd�������]6>��/Y>X>R^?}��f���=3<^AD��I
ڣR������ ��Hg�?���İ\*O�;��Q��'p�?�e�11�]� ˬk�ƫ��S�PxV�kz�[�����#���e��
��m˜���ľu�f��b
�����(��\f�:�d���/�o�~�t�Cn\�9_]��]tR�R�j��@v)*�ޗ����<n%�T�^"�%��ʜ+h����*�/���r�q:La�o�aZǆFm���Ԫf���C�HWԍ?q:�lP|B��,
�di���&C~�E{s����ξ�MC���`0�7��߹.��]z[�1���O+��9b�m-U?���7!c���Z$���o��2���-e���> ��������\i6��O#T|���NfeF��i�<H+��!���g�t�8�����5�������h܊H���CB��}д���w<pc�b�n=��%��a���j���Z���^�!��}6��S��C2��?r-S�����պ乭�����������sۭ�c����f������ZJUl渌� !��hD{�����߉��8gqI�%i(źP)�3�m�E(���7!��SW!Ia��XW��-	m͌�������R��
_�ʽ�Ƕ�����ݦ�Z��y	�^Q{WLf��C��bFm8�D�F�Be��ԃ��^�̲���E<?GAzf�dA��nC����,�|���Hw_ �x���N�����/�u�m�A����Y�}NZ����ț������O%%#�I�����2����ꎤ�M�O�;Ά�X��t�ʄ�ǚ��Om����`�e��W���>��!�*�8ܝy��!�(��,��yG^	O�v��lƒ�x4X��B����'��]�Nv�]V��\��j��=�A\:���-^�QF��<O�B����ԇ�-b��0M������$�a�-���wJ���������s�������l�w;��|�_g~�0dn/Dp����{Cޭ2<�A�c�4��3X�GюU��M27r@��^ބi�}c�/^ԋ��fF;��:����nǐ$n��KIT����m�;g�Tr�b.Om&E(�(f���G�$$�߈�L���h���G;S��6�&=�~�5�-�M	��DoաǛ>D[�]sYzZ����d�ta�����Y�Tůd2�U��i����m���j���Bτh�{�P ��G���{̗(0��o9!}�k���[x�nAZ�q.X^��ʞpw:�Ywc #M&��`� �l��^�`�ɛ Wa���_J�s(�MPS��q�P@�WX��XZoj>�VP�]�H�TS38�=�z���A�)����c�Jx����|G/�>�ε�����(�Et�0o��Qla݇{��t��Z\\��mBU�0Oc�*2�S�2���.�M:���a�r�d�	s5K����ʥElYW}*�c��C��YOy����Acsf&].�[��"��Z�l�K�*(���BBӕ7<��X@�%��ʹ?�?���f���y�y�Sv�Bݕ
-D�S��d�t0��#D>- od�L�itJl�.ɕN��m�8ܜ���N���oa����Jb��^5` ~;��&�Z����ekl�0_�A����f6�d-B�n5�5My�<��r�d0������>�FE�F�<%�LZ�H���zT`��������7�/������I
SFeF~�G�Uϼ;s0���D��N��B"Rd>���9R�u!��t�}+fO�A��;'���`�pR`�jO:�H�$���"�B��6�����J�z�k���>��g���+Ƹ���	,�,QU�6R$��k�*ή�N����m$A�.a����\`��RQ��Wy~ޘ�UϫЬ����_�6�e��ikh
��jo?q���l�P�����qt����Sfp:'��\f���C�5�=8�����	�L^D�c+hNw�}Dj+�z/�3#3��!}�tE^�1�=&)�!�]26q#jS�'�>(��@���;�.������?���8i��vH�r~��7E���汷{���ӵ'#�;�0�x|�Bl�6EV[��	E�J�KG���8�
�-ֻv&.}���y<�������.�W����;�,�EL�b�Y�Ĺ�u$�x�e	�RQCU��?�51�6d8�o<�O!̤��ܶ%��|�Y�F��"�h�3˂���mJi� ���P�r��1���*ehn�]�3���6�tP3h��,C88)��c?q?ȣL튯,Ӥ ,#��e��Aĺ�z	Rmex��؀����
�Ҏ�X/m�7�<
B���)�w�LN8zT��ZZk!���b���j�(��z�2f›T'z��q����BEU
��ZD'�VYF,��{Аr����r�g�c�yu��B6#�同�n,)��稅9�g�ZH&������C�Ԍ[8"�g-𸈎���o��ʠ�+�y�ԓ��US�R)_7H���j�9R�ß�>�#[Y�{�tÃڏ2��Ԣ�w���Н�i'�k���<$*�8��<qm �:i���zm0>Ir��[��ۛ8ɽ�d�gla1�5�y2�9ͷ��׵b!&�C� �� b�Z��4��N�)0s��v�-)[T-nF��5i&���c��AM��X�S����¶f�����]�����Jw�A
0�t嵱��b]Ї�G)C�ce�~���(��$ҾcZ�{4�����9�$l�FT]@ l�Lă_��%���40�@�{ҡ�g��3�|(��5�7#�,N� [�o��b�Z�_X�a����dDPuk(s��Я�%c��6\�������~<OPn�/#*�,���c��-^D�^���CO���1�Up��i@��8�S��?��A�J��"`7R� r��䂴Nry�W3Y&߿
�Nu��Ч �+��Ϻp"0�i�!��TyQdfKiƫA������]�ʵ�}�h�F��3��.eK9�u��;y��tz(�e)Qh���zt��=/����* ���D�/{��ux��	Gk:t_�L�������'�w����2s�@+Ё:O��M_��H�J;w�;Em#|��â����c��G~t���H��׺�������䬈��1ȒӞ����d����Fp��Q"'�zDIG�ܓ+'ӊ�i�� ����DC��J�m�Q�������M��V\�vb�6Em���&��d9/Bͯ�/s�!��jL�Vp���l�e-k�c��T��ǉ=cXN�T����ݡ������1��`�m5@�~���Vك+��jC����9���,x4��؅�E����<v�{w���-(��y6m/E0-��x��f!1����ӡ}l;m�E)~83�m:�]X��Ȅ{x�ȟn��ۘhK^�eT��e�95�wܻ�U��;K�o9��fXPB{�0 .����6�V�^��q�����o	/�ok��- �(}5����) 7�D�2 ����?;5'(qGZw��-Ȍin�c�Z;�ͩ��/r�ځD��ˤ��`6�h+����0ɇ�A}.{#����0 ��s�������A��aL���ݢo�m��n�>?�1EO����dWX����3n��!�s�I�C:��2y����S!�u��H�m�38�T�����o�?��&A5s �C��UD��3^L�BKx!x�+���)�,��0xl���-jV��?��(��9�)�C���k
��V_b�3� Ԓ�0�%ڣ���{�yF��FtF���f(���
Qi�m��4]�_)Y?,�\�`��+@�p�ξ�f�X��4Gh1��6�`���$Ι��Ҡ�ɕB��T���R�<С}�R���aÀPi��T�(��]bK+Ɓ��&t'y~�����<�_r@�wl��:����p��W�2\i�3s�o�7�A.�l :��I���Ҟ����Eg�^����d��S�wP��r���gE�.�%�?�(�Q��%�["��24�8)l���G���D�E:��,#�r����
Z�p�u�x~[�N.�oڠ�9k*�$���XxS�u���Ν�&V&��WW�GdX���.o�-�Y�7x
�?�мv�7�1�Nj�$p8Q>I���F߅E��x8��U����0�K*�.�c������������0ri�6�d�n�۪R��Jt��B���/רa��Mo��(yj��Պ�ԑƖNx6@ju�ف���S�~�L�B}��2�"p��q����-!�؉�ԓ4y��􉨪�����m쾀��:R^�9z�R��΍MN�Ce �$c�!��<��}]��Jx�]�a�-�C�eb���{=3��5&�%���d0�!��ȓ�,�7,�	n�!O�8��@5S��tǊ��iP�A��P4�T��V����(��(�}36���Sɝ�tD���1�1%*�����!���������L�?~��D����1ɪ�����(I��[_m�H7��PҦǘ}�$��kѿE0N_yڝ��f�$k�k�s�a�i�b���=����V��T����ȸN��>g|��OP&p?��|�/��~��]yٜ��&4OP�����j�ᮚMIÅ1�G��!c4g	��������ٳ'L~�$�R�D߰��� ��[WϽr
Cb��Ӏ�K��-�_0,�K�i�6
-�dT�Q%ۚ��m��7ኳ���Ι���[���%{���V7~���ODw/�Fɪ	�Oc���K��=M�-������O����f�IX4f�ZN��E}l�v)�ڗ�!;*:h=�O�*P���E!�C��赀)o9���}��ܽ�zuj@s�Y�a�ޥ	�� f�N�;�lL̓V����y=\v�6k�������]3H�	�Xv
y����)�I����l�x	�BV��6�ɮ��j<*� ~���5nT\vu1�Y7ms��Rvw������|�]9�{��)ԙ@������	(�ٽ3��,nh�YŻ-���3�a�@�iC��wV�E��[��P$)�ܭ�ּ��S�c��@mиۓ�BIp8�����culǽn^8(�N0��B�[��-��:����9b�g�B��&�`_H�	C���«���-��Jg�PJ���n^bF�"�G1
q��R���US�HN�pf�w���H��1�1�����ιa�\��'p{�s�^Pߋ�q�x&��$(~�[0ǣ5�d�"�Ť��I�)���e�ȴA�H�Ѝ�|{�B����3��g8-�B�I߈ ���]����ϴ�cn*��Ͽq�n����L�O��}a�jѭ`�� ��ڃ����ձ�nO�ot�[�a�������͞ͽ��}`S�{���>�a�͹E�D]vGP��K���h휨���]1�R�Nǳ���ǶA![/��Va_y�H�) ��rt��e�:� ;̇-�eR
S�]*�Ro��%8m@��ۋR�I���$�o?hq��녟lm��6G��?ڂ&��%G��N�s��k�_�	蹼���U�>$��+���XM�F$Xz�{)J��t#>*�=��<���{�����疐L��w@���}Y@X��6�^�1�&7�ۄ5�GY����äbs�%Dv�AZ"N�H���#�X��j���b#���`��Y�	��ȁ�9�'���AF���3
m*���mE���]���Eg���������=t��_<Nq-��b�&-M�ǚ�R)�W�#��v]x�0�vt�x�Y`�P���2����Âg�O>��@��m�F\I �ËYToi�τT��g?u�$�Җ��G2��t�~U�A��Õ��,e����M�[��Qa/ʶ�e.O;RO��]8?�s�&�mD�G���rq$-�Ұ&��k������)o���);����y���`����6�Je��k�؋<�/p0�
�P	L��H�K�j��9:�����;j{T��g�� b�:q��M�Ѓ%?;]{�k�19����_����0��P��[�X�Q� ��������g��.&`�'}wdM �1�^2i�����ު����<��j�3��T1�(�&�B�qXGq"�8>R�>�H�i��J�r��7+e��s|���	u���iMN�2d�?G*c��3� <f6�h B��r��n�z��R���i��-���x/%��@�+/a�I��4�`i7g�$�aS�c���[a
�F��	W��q�����i�#�"j�uf�D��f�6�74*X�%�R����" <@����My�
w}2�qZxOu�T�
ݭH��#(�Dt]��Ь��u^��I�,�Ш\�Sό�ںǺ�q�vH;�>����JAH�BA�9i�{����L�cw�J[� ���*��E� �0�z-��4�s��̯;ꂑ�@!A�#mj�nuc�+�2ƣo(�$Ҷ�S��b�B7:�竩@�%b#�y��z{G8��*�!�����_"���T[ 8חpV6�춻��m6�!߱ j~�\����Kx��P(	������i��D�
��!=�'F�������ƭ�p~q�i㵬)�q�M��"jt��©S1��b���P����cR��ki�)�v��dY����Z�Uڇ+�n�۶��ۦ�Vo���{��]3�t�Ԓ� ���ey�*�+���"��l�؆;g�!~Q~Lv�6*�v �E&j�u�k��w�D�����~�O&�]����u��b��ʩ)~�jV5]SOA�҄q3E�3(�H��5�,�l�/lrH�TǄ>�[�L�{E��E.B�p��?�Kˁ�u��M���\5zUd�෽I%"��O"��;��1pO+�%[[Q���V<�x���rWߒ�{�QDv�Z�qvS��$�o�o4"W���֡H�����A��`���l��]=�\�`�\��r��YIgK#vo�8��h+��>w�� ^�v���yN�ahԠ�U���By�?W-���8Z޽��<��� �']�؟-0�KOI�
�:�Ы�9zR8G ���	�K%#�6�?�{��+I��C��!��
gBI.���"������x9Z�FTP9;��A�lG���(k�6\2�&��n!;S!�������ឮ�Bl��+,chW#(���K�vܫ���S�}���	�2���[����i��!�J�w	?��'R��XYgo?�H9�f��Kd���y�V��Y������?�����hylv�>��q��9Uu05�����@b[�Z\�f���vD�Y͘����4�nRV�������0;5�c�g��b�0&��\V�d�@�i¢���S.xJ
�����)���E�*܍� ���J��eZ�a?8߬$�<TE�{?E�%�G�]�
�J�i��lc�s�+V���ETn���
��Au&	�)j[v��;�!�w6��r����GNf��޻��>69�%�h�z�,��¢ގ��V�����uc9�5}-��r��wf�Iw划�������h��f���n5���V�O@��*���+�Q@�ΒE��>��$�%zϿK��Gb���͟�u��'ټ��1I��C�����)�ݛ���vIϖ�=J�b��T��Ң<*z�(�������Z绻��A�с����
�P�r�����Z���c� �08��̼�"R�d�?z� �߫��)p���S?=�,�p�K�'�\L�p���q`-�Jâ��H|r,�� �����}��֯o_ךUrWBF�7�>�>�gˍ)�l�]����=�EA���FW�+�U6w�<��¨M���P\	K@?�O��M[!����ڌ�Bī�S�R�UiX�r��q!��b�� ��aH���A��Vj��Ӊ��o��x�
Љ�zx������F�$ ͕���g�c��1w���,F�ED�%�h?���t�-��A/�0�`k� �Fj�i�!���u��r	��s�.�����4+yW|#�S�)C�R�z��`{�1���
7�G)˓i�U%$/�U7;�@_��̻mź��b���!X2y�9�y����e�CƗ��df�#�"����y�0\���}1�u(��t�L����cД���c'>��F�v!ҧC��[X�T|OZ�K��
z��A���&��Ydnr��}�BGp4p:���jRtG
�D�*1l�T�2O�s��*H�]��E_l��)�ui�v?d�\���"W�rz�,q���M�����q���Z|��V�h ~�,� ��=��FO��Xݣ�#�����p`
fh���Ӓ���+�$�^@͑����h�m��`H���Wm��S1�M鮪���7y�̠8������lu���!� E�M�ih�oB�W��~	��NP���l�����.u��7���3ث�`�=aQ�į��������Zt���'�g�	�h��R��������R[�CBC�LT�~�U��g�������6��X���_'~)$�mn�fCb�1C(n���'�[Ȯᧇ(��f�u���z�b\(�K:2!w�N���V4��Y'��Y�]y�� ֫Ix�ч��RJ�T�2;A��F��Ds��Y`�"G��TZu9���x%��VgU�E+ue���Q��P�q�m*ۊ������t��/C&����h��7<l��d�����"ʕg�V�/�g9 ��{{�@�=����+�N��M�-XO��3��:S ���c���)����?X1"�ś���H�����"5I�����L�ߍ�ڎ��:���V؀)cס}����Kb���E��T�l�%m��!!b�����f�#�\�9?�����H�P���!��jP�R�������B�7!��us_Ơ��N�V�EՅ<q����j�-��t[l�2Yj)|\��#��p\��<��/�-�QG
}J<�9���u5��U0�mő ���G�k�-&wR�E��BK�Ԋ<o��O�?��J���ߔ��\k��4!Z�/��[��#��IHԂ	�L����޾,u�s�B1*��Y��F��/̳,��[��;cHw��A�|���.Κ��z�j�<q!9e�uQ���<
��U�.���=�m�9�Gb�{񉻊��U,ט�����к>���E��qKl�%����_��ͦ�YFb����[|�� %��TL��5gp~ 1��rtziǺ��АGR5/N��z͏��=���
`P1��v�Z\�d��ŊQ]��Ũ��Mk$�]Y�bf�n�j�w���;,�w�U���V���ī)�����#��>��@�>_��"1>�A��Ta��?~(��|�ڹ]�Sq��͔�&�,w�GO/�ļ�j8�\(~!j�#?J�vY4(�q-��j@�@�X����jqz|h��+�#I�r��2g;zՉl&K�/�dP�#��s�.�:�.o֔�;;����e����Ʃ�����P�8��%e���kh�,qNe;��glk�M�a�g;�)���7��|8��Ϥ�]oE�$-C��/���7Pi�`�ƔQ^y�(N��0y�:(Z/��P�  �`���Yd@��%j�3N�g�ٗڍ-跋R����:�sO�*����ǆ��c�rL��R�H딪�V�;tk�7<����FJ3ꊐ����`����� �*ĳl��t|����قk���9�	(2�D�h���<e'�����d��s'+j�v�C)M����$:��:�u�*ihފ�q��>|Ss�i�W~\h�;3��y[Kp�T
�mʈ�*�]�ޑ@��������!��Q٥�9�?�qYeƤ�٨Ě�-�yv�x�MF[�)P��!��G������|(:y��7ޝ���q�ڳ�U��T��l&B}��.�A��U*��Ѭ7��y%+k^�������=���ǁf2y��`�o\*3D�n�k�qn��}���F�`uc������Y�Y���G^������If��x���\��h����,���Y�.-�P���/�ޣm�m]s;X�P�~��.'I(��K�#��T���ԝ[�b�h ?��V��c���m�����6 )PRp�iwy>d����;K����?���"c���d0��s��c�Bw���V���-y�?�&C��i�^	R��#��� �J�4UjZ��y�4���C/D�O.gt��B�--Ә����Ki���;bEs�r�/ZG���H�G)�W���v���bw��:D;2�����k^�G�������`��������u��I�GJo��`P�0��6}ncG}`yKk�5�~T�~Ʌ&�%��ڐ$�?�!�\��3�=7얳��D͏�����i��p%�v��o�]"��`���KI�כ����x6M�hG~{�*^%�ӈ��T���n��~�fژ��P~�4}�
�0����Aj�[�M���4 �$�%^�>4���\�����+I���(�:�Cy˚����s���ث�R1ν���e����U'3b[�����:#/�G^[]�5aO�D9�O-ڂ�|'@�l���Gp�M(�13������
%�XTe����q��؛C��~�L�G�uaRJIo���;���4�RS5v�����@�}�"_ۙ�^�]o�."����]TeƱ:K6�G?��u�<��5X�5~,��W�n}o/�ߟa��n��dm"��S؏e��m�,PI�����"���դ�nyK��'����y�b�=c�J	���[���.�JKurvB��s*�L"�l���^/����x���7�%�َ��=����	�+� "T��0L�^����\��m+�\nA쐰��e�\#��L���y]�}�a�7:�D�V�{Nٔ.G��R��|��Z7h�����1�<\��j�PC|���Z�䕃d��������em( i��>����1�	�&^6��<4A�8�o�?'��O!���L�ɛ�6,
|�_?zM�6>�$ v<���X���ct�I_�����C��ހ��K\*Ȕ[�I^C�1�����J�-��*�Y�L���=c�a\�u��-nP���U�?߲pPx��qޛ���J�=,55�XؒD�����W�Ӊ��6l�ʋ]r�A��13���!*��T���p��2�U�?ܾ�ʓͼ��������K9
�3��׌�jA�������s���޳�%z�w��ɶ�N7��U��?e�y��#���Q�H�H��!ڌ=���K��=�O�ӽŉ�U�|�ͯ��ȼ�e�c�w���hF�\U����6{�ڙ�����m�x����|�@<��
�Y�z��#ZCqV'��X��n��;�ΘN�CabRf)?����k&�~��η�ꤑq�Ab�y�}/���6&��?'��ë����Q>/cM�,�x�`�e���Ԗ#f��nz��&�x��S��
`:��_�V,�d��I�ش~��W�|����99�h��O�������Etｏ]'k^������,�1:E�D�1t�Gư��c��w�����lu�y��88�U�A��ho���i��s_C4�K����FHGﺺ��U���^�BHoOK�2c�A�E��̃2�SՔuF{
?��^�؝�y��K�����P��QK���b�I<���Ё[i֟�[,m����&�9���J��G�m��*+����j��ځV�(�H�Tƞ��4���[�U��*��'<�c��#WP�����+�>�~!a���Ʉ��z�^��W�����*o��Ǜz*J�2�{E��?���I��1A"o�Y���OfXn��U`�l3�c���'�[!��O�C��(*�
b��}ȀW���w�h�s���؝E}�W�C����˶���g]/>����x�u��A�Tm�r,�Dti���S6��U�b�@3���T�˷�ȝ0nB�!ܪt��w�Y�Ɋ1+Х7��C�^|��$l�O�Z����a�+���S
�29��؛�|��a����^�vU]}��g� v�Φ�����<�"
9ُ��_kz\���r��2^,�����wd��^p��`�	i�0�/�r0���)N�el�]`RC��Y��2���������`�SF��v\A�2,�QN�DL~��C�)�@�%�s���<!�R�l�*�f��������/��KS��7- H���;�l�َyŮ��+R�Xs	f��v����'ۢ6��9S9��xJ��4�F�c�����/�����~J�',��E]���t���tc���#��|��G��pL�Q���=l.�A��?���0)���p]��k"�5U������:�;"�K�҆��i���	q��B�&rL�Q���m�ιf=A�NS��0]��1`�� ���K_r~J+���16`�?E��΅B��:⫻�&����S��W��x/;�c!MC��:,��>Y1�9ct��j_���sXճ�-|�W����e&�J#�n��T�'9T�
a�����%桇�ms����
�/K���I�� ��l�i����|�z0�'�O]|��Jm{�^4"��U�^��>�~"Y0��#<���6*�-O���t@́����0G�3�0�Z�	�Pْ{�B�4kS<]�����We�%U�3E�o<FQ��0��5:���� Zϛ�������[*���zv,x#gҸ�H�W����G4=Z�l��̶���v���۲�tq�Qnb��k�Sj�g�~�~��G�e����O���\)�/mL�7_�c�g��h�eV<�9߃4�,�h��[�͋��kM$�>�'�6@"�Ѹ@�BOL^)��%���� �ߚ�k���̍�s�0�Q���!氖��GS�1�p�MT*�22�$�PS7�oo�:�F&?�
���2�s��;�r�����3Z�Y>|��rb���)PZ�,�Sw��z��׿�Jj��&�
�^(PY}��uPe�*���?� �~ܱ3�h��R�"�V��0��4�Lu;g�\A����)�u/_r�k2�]'_%�tC75;+�;�oe��pF��c��R�c���|b�E)R,l�Oe䉵]���`�'���I�!�ëP\�O�R����"����dnR�C�_A*���qD@6sC��Wugo�f"l����$Q#xݫ$~/�����=�9-oΌ��(�aC�V�P�j��m��c�Am��'><��2��W>Ml��b=ӫ����4Jʎ�~�cWB����Wp�帻�������\#mvI3z@U��j,��CZD�֤��!�8�����۶6t��F�{�{s^�}��#���#�b����1|ܕR;ܕ�vW8,c���T���\,u�Z�o�)�v!)#$�%���� ����r2\$r�+!זn �B���z�\h��$��M ۠�4�$��Q��U�/�{�N�hfv�r�pq�� @l��OHF�x~�߇�E����&f(rb��؝�'4z%�M��J�_�I�gI(�{���+��L���X�+�ߎkK*�'�b��J;o2˭٪�S+���������b]�NT�橔���ն2bɉ����~#��F��EX�J�۴ �������n	�۟8��猗�)��ھ��U�^�dڸl�{�)=K-У6�UЂ����&w��<|��t���^��*3="��Q�3��qળg���R�X+�>He���-�S7h��p'�!�Q_��=$��i��OR@#8�W��Zt����:�#��b������}��&��d�)�U؝;�O%E?s�nշĲ���>�Le�$�X{��c��q�wъ�(����OQ~_\��w>`B�{f�e�a0@�p��zt��;���מૼ�J9����ֿ�	/�¿Ǌv���&^"��c��UA�x�|2ۓ��6���}��7�S*נҹ�Ċv�����[|����Q�Q��34y��>�l�Y*`�s`�s�+��hD���˞�{7�0?�5Չc1�Ũ����$��m�u���5�^W����Ǜ��Mӷ0���ʵM��#|�}��R�������a�[��lN�mUGaCv'S�{tݾa�VF��A���ɯ6�z�M�T���^i��|�a����A#�1VxD�Ћ��]LWt+�yͷ0��"֪[��O�N��o�bh��\PG�/r1C~��	���6 i�#Ή�?���7��i8�� T�f
L����#~�����,K챌Ĝ�*SS�x.�W�q[�8�-�Nz̆G`G��k{����#wy).p=��c�BN7�z�-"�B�ԏC�Ł�~w�c� g3�X��]��U��m�f�)�2�z?�<�Z-�[�^����%4���"�8�L�@Yz��B�E��k���a}ݤ�`f5�UV�n�4�E!�q$[���N\,V/P�y:���cj�\����|�g�&k�u �+����ٜk��v�_}8���}�7�_Cɂ����$8Ʀ���������1�'�AE��<��`c�	,^i_�Y�D뿧�T)@����,M��z
����A���(vO�#��c�/�4��D�Z#��/��iy]�g�;<!�J(��Kc��xآ�'�vCg���:2�nk,a������MP�3���Js)�ҕӉɵ+F�l�Ѡ��������JgB͸�XB���ȍ�&;�^WJ��ޓ��u�V�Zn6��)l?����Ć6/����C��h���6����p�w�o΁�����|(4���hƈ�w��B2�����!���3��H}@ix�H%�A��6ڗ^�˴���6ؔy�p�d�YM,���ߤ!B˜������z��g�����B�����^[�t�w�u2eQ��@̼�M
f��� �_+�`&d��ǥ
7�i�r~�^`|�GD$T��9;W:h��)��exV�9i4�ۗrP`6��ka,CjVJ[�k������v�2��y:�:['��~k�r��`˛6;*4C,;�ӯU&ϩ~��c�0����y,ǒ.�)����<�&2И��K�yV�.�ZlC��˳��J6�}*n��4+�/�i��y���
7=���v�X}�7�EmP���؂�E PHw�_�p&@Rf�k Hw�\NG�J�=����Xw�Ŗ+4�`�o-�UH�߽������n,��`({d���W�畭`���SȑL��Xc�|���c!\.��E�h���)������0����A}�]��D��)���O!6�\����{��2Fx-�V@\Z�w��q8o��mO�,���ܷ鍚-���}V� �5/����w���)��¨@ Z�w�m���͐��֤;��:�-�s� ��jħ�1�W��y�����_�fH��c�~u�(Ĉ_�|ʑ�&�7�tmqs�\+���vl����^��*!2y.Y
��Ou��1]��ں�Q��`}�ή�	Df�_�3Z���O=H�ok'O�sw�?�P+��$M����\����-�r����l��B��bRI[�����cзO�:���q5�k�sHD� 1���=r�]#>b��#���ӵo!��8Z�=�	8�/�zp�;`!(�~\�]K�v��M�.�����r
�1Jh���Մ���E�8���h���� ӈ�f�<���t�ùі���3�@�D�my�xS��dUpz����>��Q��QҮ@����x#5����ln�#��u��@!nJ����`n��'4?�]9)q���%�r�\\��E��)C�dG����A|:�����~@ok����Ɏ����K%FG�<�#}:�F���|6�<R�� |
� �7Ț%;y�]Sʵ�;+���!�GV�P����V��̢z��->���;&i3;��4%̣����.��C-*Z��1�V�����=�Ɯ�u�UfڸE��W^����g��������U^;�UF��RQ_�q>s��w[m ����Ȏ"*�}�Q�<�"Z�����N\%3�?e͙�?�?q�Ko�D^؂�"R�6QC�`����N����!]{k�*O�N�mKܳ�|��:b�DB�7lں�CQD�#����2�,O&��g$"�eo`�d}��lA��+:vd#�֣ 9*{.v��|`rf˱^�#h�e�g�sn %5�>,T�
�!'0d`�9=\B�^�����k��# ������m��{/%x�S5�nn��;�(�'$w���٦�����/#e-4n���"|[p�E�B��M�v��2,��m{l#܊s<���j��0c�T0��Kd�Ƈ����i���6��5��-�p2o���W��p�f�^ ���>�X���4:6�so��e�N�O�Mh0�����"�B�W��СP���I�jՋ�� >���w^<s�VRՖV�T��d��̹r�� �:��=6*(n�M�U�v{����Z�o�aq���J���7�bFO%���f�@���<f՝�$�)�����C�NL>'�朣 H�@B�E�lS?yOIg�H�<�+l(�|�`4SώWی����w��w<�(�w�ľ�ȝ�=W,N>�8�_{(��hײ�mċM�x0���t(�b>��ve9&��C�P!)���`�/�S����W����;�&��xc�d�,�r�3��Z�}�M������S��zh����$i�W�E�n�{�	�)i����H����5&JBCTN�:m)�{ۯ�me+����X�PXv�a��[��e��xK��v5g�-�d����W֚�)`]!���JTA�6$��=m5����t\�[�8
����g�q�q�k�DG�Z���R|�G��,Oa�}g��W	p�0�EOY���S���G�8��q�{`�\t*�D�F_�]�MB֢���+Q������� XO

i-0�m�3P����ak����K�J���O
��J�c�.E�������8�Hɇǲ��q@�'��>B��e�7j�����kU:YV6����1������i��z��U��q �N?j���p�0�F��+~6��W��5�׷]��?!�ƹ5 ����*U���I����d2sۋ9��b&Ӡ�G�7$r"��|�9���@c��^s����M@���6���³0mza����<�e���ܙ�:[O���fTt��ӡ�O�J{h.�T��s�@c!�M�a�������c+�B��� ��hjf�W���lZ�&��و���n)�w�<�P�	ߵ�}��]ȁ�ū���/Q�Q �jqVM�"��c��?@��G~ZPxby�XI��n����KA��]m��96ԔA�a7 B7X�#�B12������(Sq�E���^��~�Ԫ��~��9��lYjR���L��"#�@̾�Q3��&mR!zWqO�Tʖ@ȗy�P�q>�3�g�g�w�1��gIjj�;���v�ڂS�sR�|��q%��������-�w�!�y����#10�;���H���-�hK3�z#=R��^��@�g�1I���`�A� ��Q��4�R�o���*n�o�=���U �a'r~W����@G+2��欅w-�ݽ%�v�ɦ��_�O��G-/;>��m,�Le|�w���;��t���XJ`F�1�݇�lgu���9p�W[�
�%�aЩ�_�L��wIT��?��(Ě&|�����r�]|1<Vhy}
�Boo��hv5��g�pA��<�d�+���q	sp4�����O��OE���Rѷ� p��L���rwߨJG�Go�۶�7��.�ӻIb�e�A^S÷>1�&�ArIbC��х��`(��%���A]�����}6 �R����	HG�<�#d�#�IzR1m��
�gu��6gO�䎇$�b��Mc;���1�td�&�K�ĺ
�ŝ/ ؼ�Jp�g뾝�9(��U�r�Ypt=.!��a��{�-�3�)ʥ���8�^w��~�,�	�x"��$�h���ug�����>�0^��HA�M]p]o!�|����`� gx|�����Lѭ���?#m�r75J 0���$7�L~ �;�\�m{X��0\g^�o90�s�G�@,��`��t�j˻����Tˍ�NF�Z�� �P���<'|�ud�4��.����{�V�Ҙ|������M�oR�]nxX
8�����c?�yZ��i�+��i�<$W*Ʋ�����=�0˃��hp�6�)�~�{��|�����>9�8��	��&��\����5$!0�&,�͔`R� ]�ٖ�/$�U�Uu���d��;�S���<X�2J��9�a�͸��m:���I<8�> b9L[�K�]������@�Ck�%��C�($�yva��]�a:��F#�_K�	~�Ui�)�R�����&P������L?S��.T��4]�^qH��^�۟���J0��b`m*��k���A�C��Lf�V1�nz��x�%P�kƸ���@{��x�L �OXRH w�4~��kً���18ʵ�W���H���,��,�I�5��J��0j,��Z��ЀV�� 2#^�������[4'�EA�����{����7aBg�߿�L���7�6ȡ�3N�	H��$��&�I�$�L��z�I�������Mh6S|��zcsZ;��K"S���Bq6�ڸ�*#q��)�7W�?LS�<G)_�۲Pu[-��}�C��fg<k�"x҂LO�Ι/)I��{���
�OVƳ��P5�V����`�Q8��"j��Se�Z�ڷ.�F:�~�u�J�\`W��wWI��u�E��% M"���ը�o9ձ��9q�	���
	v�7��.������L�&0J8�g>�hB+5$�=7i%-�@��ŀu��b䨴R��l"E�O�o�O9М��G'F�b<  �����&�����=��i�J�h�ѰЬI޾�,�Dl��K���P[����j9W)!�?G��:�t^E2�
�?��]�u,7��iY6��U���5�#<�Y4a��HG��ʤ�������mՃk1�(h]��H,��ROM��F�	���47(�UQ��4�G��L4� �	��?�v�teB�WX�,�ᕏTN�v�4|�607cMW@��=��4�Y���c0.&Ѩr��&[�*uTq�P�B��<%�1��.�2x�QHT��x�O�x@X�8��^��~��i���m�U��j��k�b9{���As6\�u� �}��D� R�o��zՄ1Z3��ϏͥNI�=f2�Y�c ��a+D�1M�|1]��f��fPű*Ĵ�$����Ʋ�#ƼO��?^��vX�Ds�a�P7�8��@ �ɇ	N�HZ͛fAN�h
�
��c�T$����@r뺱(���_z����Y�e�A�<wW���>�l&���U����Å	Sퟢ�C|�JGQ�tI�8v�
,	H��J��k��V2�%B6u��ݍ��P[��B.��9��tɣ��`UjLP�n�t�>�9�b��Z]�Ӄ��|%�
\��^*߈���Je B<�ě��kcU��(K����1�7Χh}񤋏K1e}Ʈy�1�jo�������T�`�S��b��q��;����B(���CqC�jj:Lߴȵ��\6D��8G*4YC�Б�s� ߪ�չ���3w<O�ln����(+�����ݓ��w�����_L3y�eє2�l�X�Q_D�S��f��O��ˊ�
Ӊ^�=3'�D5�;�B�bN d��C� K_m���Z����3�S��)9�x��{��sz���г~��y�G�2$�f�>8M+m@ߵ�7�<d+���ӉޓG�K�,)�1Ż���C�xq��\�5�e~�i����ە���J���}�t>Nb��viP9��i<� ����b�B#��?t˺4��:���!y�ٺv�	>3��,mOiU���%���6���d�%J�t�1�1j?S�tDd~��p5��^�Ţm����Ĥ��,y�dvf������"�ɽ�q��e��8&M����O�H�?y���q�S�[R��u�迺���/���ӽڀ�QC�I,U8w��:F/��>3�L�Y��-p�y9�og �7�7�E3;P*a�}]������먜�\e���&���iپ����B�=� 8�;�X����b>��7���qհ)ҎPM�K?pc�mF�%�-��$\�� -���k}�kl�]��>e�Z��$M>섧ަv�i��]2���ֹ���R�c�������vx�;=�x�藬 )�2o1�{�ߒ@ز�UU��B���4M����n[[#/�����a��
���������5����|V��x���nvl�-��ۋ�A��i~�?2��o��߅�մ�u���4Ǌ�!+ቭ��̰g D��E��c�5�bU�����@�6C⒋���a5�V�����p��g?�g�� ~*����n)JI�B�1-�uC(�vhM��I�))���"�%5�'A��Fj� |o�]��8��������V�`%�B���uL6���8
	X{�$n��掾��V|o�S;u:�{s���OL ���c��a,�q��K�cvl�1
������1��H��/���(���>�8�����0a6�ª��$Ȟk]A�X�YAJ=J�a�!eQn�F\�RdU⑻;�h#���Ӈ�bs*�2���_=���{��<Z�{m�р��sA.e��m�Wj�����N��;i���R��7���$8�#����f�kk4áv�1�T�X/l���1U�����O�I���7���T�z\��A�^���iͨ��G�>�J��Gg���"�
$�cJjI���%����~JD�q/[_fG�"�����<��4�W��¿dY�SHY��YR��$'9���C��/�kt	�=Ù� Y�L�Sy��:F�����J�z��Yƒo}����T���w ���+�(����D!�jz�o�F4�#g�^�&�GZފ�z�]���xB�8�(oc�^o�7��>�O;%1��,3oޢU�B +d1O��o�c��^|��׭�A*�qH�1Ӳ�˙9�c�AJ���x<��ۃ�n[N��E�����7a��o����+� ��yw�D��S�b.�x��W�?�6����,Rx�f�`}�RR��=.]:��tݕ0�B�h�=,����	N�(鑄��]�6��⫨��7z�Λv����u����q��7Eo�IO@��)$Ғ��o]�sV�������&�\%T��9����N)���]��"V���-��V��8���{�+�i�0���\q���T�%��Z���B��x����a��5�wƾ�R�C�B��.A ��C���}r�T哐�
��,��%�4���o)~��!0�M�r�y��-��"=�����Å��趧���,���I���܍k�����pEr\��C�F��D�j���N B6��0�����j���H2��k��Ơܑ�.C���9K���B��c$R��#H"�M�~z��W�qeL��T�I��xγ��+XM�{����&��l�	[,�p���%�Na#;����Q��֙f� �=Hҡ��_Y��B�������1���M�V.P߱���Ҟ���k�HmtצּY�r�sc�R����_�;B���P/�xG#74b�H׆�D��<� ȭ@$�Xs56"�(���*^���W��Spˇ�*p�y+M���w=~!���P����� ���'�,R����vN�5$����Ο�v���ˑ�&\�T(�.�M�ἇen����j7�����ĽW�o_8��|V��x�?��w�{5��K��?�_>����f�ŋ��p�^�N��B�-�jjn|�~���߸"	y�)����)2yj��t ��¶�K�˗4QФ�ۺV��?PӮ����L�[�.�]� I�H\=/�f�41����Q*ڈ~����?��w~��n�MY|LԣW-Qz���[+�n�x���Q�0����?���ͭW@ Yn\{%�� ��r��o�/�A�(K��7C��oB�/W!I�ƍ`r���#�$B�S�!��_�6�qڬ�i��.E?����ϗs�$�6՘�q_&������w�ĳ��ڐ{�����259�(�k�U��;?���FSMhu};؅����h��_X� �";��&ґ n�/��k6Ћ�5�ا�w<�����ȰҮ���0����ؿֶ�6���� �%x��������G���Z�$��[��;�|\Aw��[�5Y��������{w8 �WD��a��� �V ��{k-X�$�́d�L����5�Gx[=QԘ�f�]�����;O�#�  �#�'�������$A��YV㩴�~>��ƕ"-�Y@��Z_=�?��A9-�rpZ�3�	Y�Dr�����(�D�(�� I�߁P>S�5�T\�D��#j�`�/l'=��(�"#���^F<|Ek �����q7q%��B;�V�1�wm�FFͅ8w����W-�Bv7�3/�=+�4���7L:B�v��Ѿ�Yub�bPZع4sA������S������:Yb��������!��'C$	-P���a�����hI�b��1.�ٯW���h�ꔐ8�'��k��ݾ�'[���k�s&�4j��;�S9h��
S��/'�(�"��!����*V��Ti�%Χ�9�7�3�~p� x	*��7�ܞdik�!I_� r;��eM��=�R?%-�T.O�ޢ~�VrM<B�"�j6 �=�4�>sjn������sD��~�珀��H/,ǈ�.ٶ�x�5�!�p-�Z��=��ۑ�3�ҭW( zp��T���v�O�����e��#��$| 	D���зjRkųЙ��*����K[ӣE��I�D�XSA͉�섐c�n��'Z��;x14X�N�p�k�8cّ���6��2nq�&��f].Fe}nj&��I�C0D�D��-��Ġ§��Mq%h�5xW� !�Ŋޏ6�*�:��J�ک0�:¢������L��Y��"�	�fџ|�諢>�,�(�)Ԍk��+���TH�H1�A#�3)�p�G�E��4M �N]�z��^�L��
��-յK+]�І��	�h��������E�=P�m��k�OXh�$�5�eU�&Y@Qe �W0���n��ۻpXM�2!�g�կ�ޙs���~���r&Y���,�yǘ�8R'ڷ3���N�/#�2Q���kü;���M�_�b����Ԁ���Z�e�.wģ��w�3�e��e��(&��ŝ���4~�a��`�(�>�X�	����: x�ُ�r[���}YB�x'��R9����b���+ɉ���c�D9Kz&aP ��Z����Պ�S��]t�����:����lS0-O|�7��q�����\��V������ɎRM���>�C���=8Ez7O�X��=�Py���,Ż6uF"b�����B�]U���:H�%�'�u�ha�9g[�p�衔۶��b�\6 �����oFÐ�\�QԛbZ�WJ�g�Aޱre�{
ט���n|��tЌ�>J����tK�����1�S^�7U�l�
o���uy����bK���C:��-�#Gp�d��Sk)f��l�Q	я�׼��f����d�䏟.$8H:�[�%(I^9?Π��R�5�*� �SO�M����):;��"vl*lZI��7f*"�4#���ɍ3%�uh�١������t����K7�=,��иKĞ�d@����Q�2K
-�e�[B2��r����UYZ&|�ދ�!��2�xbx��?�:���/���F���B0�慈�Q�e/���5�^�*
�"61��)�ͫ��7Sy���Ҝ�zG����}�+Gs���'����UC��~6�I"���j�L�UۺrN@^H�{�5�iM_^`]d%��GF�����oQ�Zԕt8�jIBs�q3�~�|t�`,lm�/Ks W��_���v�a�.lp��1����_�a4�رL�>r._EK���������Ϛ��H�(�NX����a�i�ټ��գS�����$�$��x¶�"ű/.6�))��ݔ{�����.}c�N��8d��O�6��x�U�r�i�SPX������ �����;�l��د�?�V�}-Ǵ�n׀�m=K��`A[�S��`v���\��k�l����Z�O�B�Ȼ��]�ee1��"��ˍɳ�uV~���B�d:��:���AF��p��{Ox�\9PK�a/�yɈ��ȃ��'��5v�f�іU�-�\9���o��%^�L`7�O��u����/ۉOQ�,�TEj�EGA�_FT���e-eګ��{���ԯԆ�o�
փ��3va�xF�f[�;w�=u�
�D&�q���cn��r>�mw�ŋ�<������Г<��G*^�XW;R�ID8�,�3��L�7�{�*�f��U1o��P�zG���d�p�rjB[�6/�<��{�w��>զ�:��9Z���%6'��
��� �!Ahi�H�Øn&�llɦ1��.��]��]�P�S���Z]̂T9VH坞q$�<�P�q��G��ḴH��HV���� 46|�	�����TԨ��x�R1^s�)��"�
��?�m���p'����0��6��]>*e5�jOݖ0Lw,��и)�
+Q%ZnI�FC� *�7��Pl(�|zJm�l �y�«�D7/���ܞnbbb�OB�m��T�ŰP.�U���]�o˼� �G��2����*	�A��>����SW���x	�X86B��⋈y��h㷟�d�0��=�?H�@�gnMƳi��+rĝ�[Ƚ1<���_�lF��1�D,�l@� �7m�_����K?�Gms��E��R�������?+�`�j�
��I��c�f#A���7��
,���F0��`I(}N?�=b�W�J�v�d���)�\�{�~�Z�D��c�����.O�p�q����w��`)W��Kq[8
+�̳۟��[�VT�S3��}47��3�f]�8���T$s�9��b��y	�C�{�(0��.Q�!��|�X�R�'��k���A��8��U��.�h�w+x�����|P�30��L�ʦ9���͎�q�{v�Ԣr������e`L�Ma��%D�}&D:s8G,�z�<����w3j@һ3���Y�����;3l�^p�K��*�����8N�g��|�8��;3���pm�J�A՚�I�4�É _��nF%��H�7���\ڦ��i�v���U'���`�fJ�#G�s0W�$���6@R�[,�Xn�l�"i0�u0��T<*w�:+|��^���Р����B�V���WD�.��[Co��mT��Ś<s|X�юvaDu��ExWq��f���G"g��e(�f��)Hcb���i��>B�����$$3/�t�F<��U+Ig�0��ntM��o�Xl���=��b�I H�4�mڷ$)>���ד\l<��r�|d`'B����y٬ߌ H7E	��
�[R��̩>
�*�YgV� 8���5��+u�R��;��E1^_?��{xm��z�ѽ�kx���7=��ى��#���FK���w�hJ_m�Ur[Y�s��y\{U =�O�s��nߢp�e6�!	��7�1��j�[���!�ݗe&��Gp���gq��0�mi�������</�Vǳ�E���F��AQ��������$�o+I{)��ٙ�KS�����&�r�a�|��6�<��ͧ	���D��Q�$���ѓ��N4O'�T�����X�������k;�<pYo�jb2��t��'����a��u�K�~�E�Noe�celʗ��fz����x�ng��]��$7���e644�IS0"��2=�z%�m;��{�s���
լ��3Me��v-��$�l=��Hx��&i��6�}������ɀ�K!�hu�9DS0�NFǶe z��B@��6��y	DA���w�c�����V���e��1Z���Q�T~w~��1�ӧ<Z�����b3��?��H��A/h���;t�����E�ct0�(3��@!n>Z��&�"�ʑe����s$��ZQ��v�f��������n�����3NG�EV��p�D�w��C_�Z`��ʐj�T����ذ~�vdA��):�gu���.5n�䈤k�O���ؼ�p稿��e�ܞ�� "�8"�8�ONe�E.AF�21�s�N�i�I��.�����6Y�U&��9|��f'��y�4Tr�hhH;!��#B/|�(U���0۴�w�I�{9Z�PnY���ϊ[Tި�Bi�(�b�P&����u�N���ӵ CT2C��Ȯ9JS�g����	��Ʒ���_U�w^dv��@||Df�p���<�����A%���������A��&\:k��?��N� �������O��(Xe8ێ,_u��p$����<v�m�G��%��Ψ������y�/�Xw��_5�.?��r�������5�Qݘ��q�[��]Bx�3"��9�=�G�2�5c��i���a}�7�^U�yѭ�Q	@�6�f4o���[|R� �"h��Χ:��H+"9�ߨ?�fu':c4�8��rZ$п�u�+�^��cV7��sv�o�>P�Q����o�7%�{t,NH�"6B���Y�8�ֆ]��)�� �15���`^�A0��$+k<�t��{U.$Yg�lE&9X�d̓�#����l��gX��M-/���%`\l���bTHG�ҷ�����T|�n)a���)�̓�L3�1X��X�BTr�߷Q��Gmye�,�Պ5�6�t�a�[=ym���\�l4�Ŕ24�O�R�������KT'@�k/xz��1���bmȰ`u:]i@�S^��j�nc!.�Pʰ#��-%��pj?�
/"\~	Gv���7�f�%�K�= {�L9���hIE��級���&�GE[�\	�yz:p�S����"�S뫋�U�Ok�Q��9p�,�ş$T0�_�o�d|�;ڪ1 ���
T}��_�'�ڇ�b}|f���8h�,��h��s����h2�X�J�ٖOMx�F|[.�@�h�Ѳ�^����I�_:���_�'$�|�5@��-9�be�lǺtx��`���n��X���M�ȉ�V(�-���c\a�~�ĭ3�͆���
�WA�=��7��&�=�G(IT�]���$����:��nc0{^�>5�c��19=��w�Q�N@8�+�O��<���U�8F����_6Ue���e��Y�鏪Z�E�#P}-�k�U�@w:�iXN����m>�CK�졭I�1QʫO��E����c/#iN�\�x`5]/d��	m�FGf8�VܕݾȀ�T��"��Ok�	,EQ\�.����A8�����ާߤu�&��I6AZ�o�X49�%`�c"XM��C΂=B��X<�kb����>��k�EshD��C��<K6�4�T��آMiU�J�'*F����W����nYU%?��B�y�2I�7fi���j'~a|g�8M<�L��t��|�-�����@ר<!��|�qr��:��XD(}�+g�y�TcY�MOf�m�	#�Y}�0�i��*��b �F�_���'_8���b(_x��Ɇz$�����v�I�*E��3��f�1�l�W�w�/�E=�n�a�]��o������d/��֩q��W[e^�9E��`�c�����O�Қ40�թ#��Sİ�c�䤽�V'=�!g����;0���3�iK��CH���s�@�2�lt��Jq�:^�obD)���T&HqEO�t�x�q���@�T&፴�'A��#��u��榗4���֧-k�U�ELE��V��Q�<V�Z����فr��e)T���#���}�\���U{����V!'!;�)���U@��P]l:��p��P,O��I���u�ԗǖ���aʏk������C�t vJ����$�T��<hd��/vDl������kT~y�5&�M:��&o�F�����,��UA�fz�c��t�у��Q]�߱�ÆQz���t��>]g���a��>^\q0D6`c%�I�tE9�Ё��{�̀g\����<5�3j&�}���� RK��D��=b�w��Y�U'�Jn���ר���e���7��� ���uu�q��2`2hd8�{�ҭA|G)��f)fB��]�(����qE?2�%E�]��EY"M��S��k��G�%���{5�L�b����=--����FY�I��ܤ����6�7�,D�1��'O���Ґ��VE�#И�WVk�׹�����Q��>8H���3��t���n�T,sOeE�bu���>�q�N�7ȏ�'{�Ju>�I0�K_��t��3�v͊d�BD���["3���`�%�j$ ����YoA�J�k�Ms�3Vʳ�<���P,]��v1�!t)/���J��o��U6�@�#�_�t.�"��Bَ��h�u�I��K�]4�Cc+-�)pI���cÐ1p$9K�\�U|申�n�C�쪸���49�mFQ��8j�8�#�qi(I�~!z�Ѳ0��+�(]�I��^�.��*m�fQJ ��������� (�F/i��/Ѥ+�{��<� jzG��yr4{��������ś�dl��W��܆���#�Q���A�g ]�x�n���*��pO~Ff9�v��Q�H�'�o��>�1|���h6I�*���}�*ƒ5���"�+�Fm�j�ZB�����V��r�*3T�-G8�}cj�n��>h�7��' w�h	9��ӎ�/m�h0͵Q!��k�`Y$H=�Kbn%^i��,-r8�$�,�T$#��C~�u��dG�"At�v�
����o��97A���@ߏu��aA�:|������Nv����7�|�N#v8�^ȯ�ɤxM�.���ճ��CP[�UEM����14w**��S-�!&=�gx��딏����0�pY�U��H���s��Zw�\��P&���˩�N���?���U�V�
��P����2��^��E���ea4��f���s*)����!!	��(f+ab^D�KU(7���>^�����w�_�a�i�kz��I�/���2`��P2��,��Y��P������˨����U�d�@ә�u,-��]hӔ��7����X	�;sղM�W������QW�6?���7�,�$WT���})�UN��p��Ů?�ew��6�Z�B����/���Vrq��Z�
�9{z(֋�
�킉�>6a��M��#�J-���_+�!+��g��ꚪ��^����߁�}8�����dK.Xw%�w[�R_�$ϛ����a-������r6�򩝂�����98��A�� �\M�"}�[�WR+�iR#�kr��-��: !�� �9��E�>�:Y��f�ԃ6K8~�0�{K��/�}�����.ش�"�Yd܊sC"��g����K޸�+��J��)x��k�5	^:u�$��e�E3��zp�p��Bt�����
�K^>]|���U�#ݾ�	��5f�v�0�63�M�Y�q[ ~ #���{�X��Iߔ�`ڝ%J
�پ�Fx�y.i�#c�/*���߷��O
KY~`���#4t��8v*�^�z%�1�* �b<]<�+�U��?�jU�⻊7�.���2XL;nc����b�Ea����n���C�p��
�1��쫖dW2(%3��@��\i�n����|9�*{d`�<鐧�E��&{@ ������{�凌�pZ�Ȱ��C_GMW��O�a���J2���j�y�ɦt��A�)��t�����9d�~���\�Z��!WI�_�d�L==�?�a
Y����m�#�}�\�Ao�\��;hrx/�y���3`�n�\�k��8�w��zK�MKcܦ�7EGZX��!�`�c��V�S�ˍ��E���'7�+�Fu��ˆ�b�\�a@�Y��V�{˰��f<���V���%�+*@R7D��:u�Ȇ�vQ�[z%��r���-���J�)G1�<ՑId�p0fh&������6�$�2�S|/�0m�*��KA�?-�/
czw'�'��T,F�;9�����L�X�4��y� 돣�OI�|�P��:��͌�6E��BŅl�S���ax�g]�#u3KWaL,�IWL|�\�v�\oJX��r�7L>� ��6'��6���r�� xT�[s�a<�X"B���*�Ko��8�N7f
���nO|�
��H7�f�������h�����gT �����1	�}�w�Q%=�:�&�{���#r�,�ꪞ$-��,�h��=$2Tc*�.L���n�s�� 86�;}1n��ǰ���B��[�%=��=�"��~iO����3gM�\ެ
�<V����^�M�P_����&f�|9��,���\�D��a6cN{{��db�tK�z�]��Z���$'9N�D5R3�#N��a4�N�ق(�X�*`��rm}�抛� �#t^�js��[*a�i�0�����#�bC/j�Q�0-�B3���r�̱����\"'�EaFp��t���%*�=�t6�j�� .W������y]/�N�'��R,����g�N��_�s��Z���e��o��+��l������;}��I�&.nF��R՘��e��*/{��B�Y��sQ�9\m�v�"'�.�y�mg�HV���G�ķf��Ɉ�fN-֜6�1A=v��=B�0m�
.�M���=��*���6���g�<��l����/3�}ۄ��=ݚ�,�m�OI���V�*PQ)�ڷ*��F�Vz��Uy qKM�T<N���ؚ)��p�T�MI>`�����J%����̀!R��X�~�n��̤�س����dio�Ϧ���گǲ8�p��e����[;{/A�M��h��
:�foPۃ����we�:���[A����AV��0*MH����|�i�m��n6u6��p*hq��4���`�)�����MR�dy���_f�椝(��C�YzG��Eߗ<�L)咥�L�48�E���F���@Z�S}&�	�|Fr�|�'!�����/��sߛ�J)3�.qX)P��a������O8��d�`e)C���n����h����OD@�GA���7�����q�ADQ#��bB��N<���n���.R�9�͕��B�.����?���|��a�����@Z�<�/���)G-f=
�
q롘�/�]�\\���|F��k��}Ь�i���
�D[Տ^{�X �Sik�ӳ�I-��V���D)/'��f�hK�_n6�v?s�����-�"�k��Yt���1/v�k>���#v��h�`=+��%&)�樕8��GϷf^6/����� jSBÌ_��R���o�.��pp͵��S�Z�~�lCH�;t��O}����
����s~��7��e�K?��X1�qG)��{r�C&S�g�t,�5�J�/灁�V�K��1c�*9��:����I���1{�@0�pRl�Tm��^��:�&�w6���9��|����	G��1J�)~N��z|����lt��y$���X
��Mdp�ڵ�O!l�*�b��A���/U�NV�:����/Ap鯦����.��pho�A<�^�{�Z)��f6������!Y��u��*(�q�[�Ȑ"j��6�yO�\um5ͮDF�"}V� o7r^Cr����e�4^8��@�}j�W���w�G>s(>��'�̊��Eɉ@�<M�4*�﫿Q�-Y�N���$���x��@,�6d�B�4ƈ�!��/�\w�-�"�	J����3 S�����д��4>�]}��z�G�Z�2����Ym��Ψ;�(��E��������4~r�M�'A��ݙ,���ı�Z�1B���Y��D#�@Rk�NQ���`�<@����9�gÓ񪤬eߛ
:�|��R\.=`�±��-p�1O��ߤ
�(���3u��,6�c��M`J�R�t��	��x�)�3^?�0�#��l�g�,�9���3��
����E�.HU&'��MZ��8�ҁI���K����Se��{j���I������&2'�m+0T)�6�M��xN�~X	�&�F���X�"��K�Uf3����K��4H4>
D���tO���C�;�S�8l<��`"J"%�R�*�O/=�����GO�o:���쯽��/e⟪(ӗ�s�Q����*���qP�`K�M֦�i�nS{Mp���������m3�;O�>�3�Dx�jm����h�ޞ 4,�����D�X请�M�ˎ��p�F�FN+����zf�P�Ar ��p@g�.B�H����b��qV64�"QL��]�ik.3HD����	�X��"�&t�c�EW U�mezԾ�L@y`���Cy]'O��,�'�5��joC���Cs��u��;s�n�z+�S�<-`/�k{0p�P���!я���ac\v����kb���6X\r�0��+�Ҏ���&����ʻB>h4����Į��Ihˠ�	��������@dE��͠�l]�a�!�c�%�*����w�}�?�������������J�J��1�й���;.b��z�Q�N�ca��&߀�^�]>�5 ��n��S{��u� �?����ܘ����zP�M������|_{�l���֛9|�$�YL�$^T����,0ы����S���F#��E�(q� k��c�hë��x	0as�e��'s��yݞ�n~��2	�ђ�w��\��<Tis�D�Y��x]L�ӌ��Fوf7������݀���S��r'����?�<��>����:�+�_g�.~��8�M�~��Q��i���d�nILw��"��t8䗿��ؤ]��yK	.(�v]b�hI.������� ����_�����_�5@
�0�+�F��t�1(�DCvt�4�)�RD��u�S~�jeN*�p��܄%���yf�&O=׵"������Rl�x?�R$\��ݟ1�i9�_P�L���u"<Z2_����r"�������t�[��$�?c���Q��pnM#��VG��)�H�yq!���6ާ2�v͏mW�ne4*�*׊�I��k���Y��u��;܌u�����\��h��M[�<��������{[���ڢ�:'�u�)�~X@��S��%^
hp��S��ȗݾz'�:�:���I��l<6Q@�Y�6#7!� �=�!Q�z�.�?X[��lq8�<2��9�7s*�i&����6�i�kn�A��@e�I���RO@
'�QQoOz����Fy~8U�)�ݯ]�F�#����z��[��ĭ"yc��7I��N٤*|tR�@Ԝ/};����!���Ц�EB]Rh�d���u�����% [��ʸ�g��O4��k��� +Q���i� )�n�R�j�5=������i�P��e`��,"ɱ@��	����@���4��m�g�"���̪������o�L{�o&�<�J�i��������k�@O8��2��K9����ؗW��f�Q�u�FbM��S�fYHr(��Sx�;�1���? 8�2��	���վ��y4�����œ}�E�@?�מ�Z2�
��>� %?�*��I����N'��^'LQZU���μ洼xQt���R�&�	�ÏB:�q��H�S>��ww���3�?��=��w��
�� h��(����U
]�%��Ux�!��З{tY�S(�X�I����mw�{l��{,Z�[|BٛG?�b��x�f|�b�Y�**�x�	�C2P'?e\���O��a(��A�\��T��_i6qXd�h�n*-�u�R+^9��\��ɵѥi܄37؂�^$�4e�C�ng�K��T#;��w��m'�\�@��`� 8�����	�z��k���^�\U-���%�Gz�A�����q}D�y.��+�"�v���{�b���"�ܦ������A��Dj{��ЂLSv����dl]۱�gR�,t,�_&��tI����@)�ݬ]���tؖ�ة6�S��`��:�>$�9F��F�R��v�� P�h��g�hRt����p~{i#ѳґ�<
#�_/n�Ш��9i���Zw�6�r�uES��:����d���J%NY��o)B3��Ƃb�}�ފ&z�4}z{Ɍz�9
m��/��U��j����Μ _܈���	�R� ^)1��2Yo_� �2s���(���r��� �	�VU���Ul��*qy�)�A��XB72���Z&8���q����|��vP�[X�F2�Sw�� !wx=@G"̫_���-\
##�f�.���ϴM��/5P��q�f6�4�C�KA��;�c�l�X	{:�闚e'�n8Q��ߚ}Pz��j���)���\���;
��(ʇ|%(�P�~i��w<�a�p��b�O���5�&Un\�	R��Ǿ����ͥGbB3����8��mVƨ&dlLf����@h��4r�&�Ny���B6k����]�� [i��Q���<�`d��F򁚎Qe�hy���x��طk*��"�Ɩ�>���O�����8�rOe8����g_��Ӳ����"���.�1�������4[��:�����N�4�)c�ڟLS��Z��Lt��}B��`�Yޡ����G����)��s�c��]Zo�N%kPz.Ns�W��!3�,����㑙�0F�����s��'J
r�%T������b"�`A-��X��U���G7X�K�ү��\jK>i�����-f9��~�k_,5��M�5贑��N��w�D��Y��tK�h9^[��?\'6�tgz
IT�\j�1��U�'�Nb�);!��e����Y�=�#������m9�)��iO�i?
ȏod��ߔO.ጘ�s8����~$ �qX��̽�q"�zQz��T�RϠ~�>x#F���=�Ý��8�������t9���]���\&Ȇ<\^\������B3��v�՛���J&|7ļ�4�#��Z}�,tDv��¶0]f���p�$z)�e���ΫSnHub|J��u��H���e�d	�<R�F.meI�!������B6�?����:Eb�������߅蜬�)9Nޙ���<���A;��$3���c`�X��s�D#1r�~���g�/bQܯ����,������8*�	��L*I!.�UD�!T��-�O��z������o�I�u���,`�3!R�&��fE+O��0��yA�p�b�:��e����� "়�o$L�t:��)�����ʛ' p����Ȃ9]�O)5J�~��s3���U�<Z�`�WwJ�p)���ِ��Dy�U�Ѕ�N��Wfߦ.�}-�z����e��^<<���a��^n�-��/��=��&�gR������j6�,�J�c�~B��ˌ�-�KXD+��.��auۅ`�?���ٵA
����p�H�˯�Wx��ܫ�L�I��H��R|�0X�4�QR�n,0�W�I��{{��!ڊ�‼�ʆ����\�^m>Z6PM�+�~��\џ0�M���k�N��:H5�Wݟ�>�g����K��^�W����0�FRh�A�Ti�Eºs�TL{r��,�\���E�}��E&�y�z�#"�&b�_,K�_7��^�����J���7�W֞g�)�iXRbN�g���6�4�W$��X�a9�r9v.��GL�T��!?��7e�&{�
�Q�K�ئw��v�Y�0�לn�v�H!]�5XC;�eW+��G�{I��ԊvE:���䴲Cme�O�C[�ak�x�;أ�S( +6ϱ!�!9��(��Q{��0\�cŜ_��=�̡�T�_��n���ob�$��(���5����G^`�9@���B~����]�����
Ii�7��ƌ�TX��( $�Kg5�_�	��K	Z�\�K���/�H
�NlI�);���ҕ(šV��/���t�G�Q��أ?�R7 ��2�9�@�?��"�ѳ �s��f�'`Wk�2�=2�"��ބ�\�;�8��6��Q;�q-g��C�K��s)�*�T�)ɦ��}�O�/\�kM������v�����WY����L�.J���.Rי���>���3��"
��������ރzV"�tF�KU{����-JY��w�I7�`�m��<߈=��ct�W*�<�1K� ��*�	��	8�1/0�M�Ւ����G\�|��Ok|�`w,Zc��-��������i������)y4��A��5B?Tv����zxr����'>���ͥWZT'��0_�Y.����>"��nu�.�Ԗ�j+��j���g)@�Bh�Ѷ��:��X$���+b��lU0������%��X�%%f,%���K�k{P��\�h�h��~\Orv6N���gu+�rm�WV@��Y��zh<ao��_��7:b�&BXq�Z��N�oy��aVΖc��j�C=,��c�Vw��?�N҂���ޢ�11Zl�"�V��5Z$ؙh�=-��9r���CًsM���Ml(��Z���cL�/@ oq�tQ+��T���jg ���_[Gc�a"�TN���<Ҷ���Y��@�.4R�/}^>����?&��� �{O5�'��)�<Lr�ִ<#�i���	b\91�Tt���B86���k�8���V�W*f@�=]Zq��#x����N������ʈ��:��n� [��/'������Å��I�HZ�b-@�MP��v��7�.���-u&f��H�4�:Kt�;�N�c*FT�Y�N-�vt7Q�t%�
E�W���7�
������0-�B����é�\��Zj]������V����L�S6ܥ��p�򉘳�y�7`���A��s�[Egaޔ_�̽��4(�~\�����ssa\����MLX�?�o��Y�n9X�`Û��p�e�s���@q�*���n%�p�-SP}���-��@2%�ͽ<'������Ӱ��kK�|vu��^{��@�Ҍ�Zv�H�1׷��vʪb/���"��S�'�ȝ��6$F	9�a	�U_�Z��-� 唄Պ�g�<h�T4���-�n���\4܁β���`��$�P~��AQp�U�/�7���+�p��W�����X� ��$D����	��(m:f,^�����/�e�e���B!�s�.j�ݜ-r��0ue�%ՇDh�����^����9G�?7���Ԫ"�C�&��?�������Ur��ł|�?p��+�Iqlðg7���Tf�(�3 \e�EKW7����C4�X�3�h�s����7.��reJ�Lqk�c�c?��.������&	�I�<.�&l����Fq*�`����e�6O�m)J�����Q�(�9q�����id���]�D`PH3΍��v���r7U�@R�VޤȈ��.U��uH��$�T�wcy��+�Q�q����v"�dtu����u��-7���V&�.9{��5��F��d!m�ĩ,�Nʭ�'@����F/�^gp������&ar2�&/Ì��Y�c��>�0ok���TL��!�F_{��P+���چva�^�U����p)m�o3�@��%d���U�IX�p̄"m�U�U8�]���o`BAK17mI�2�0Z1`�7�8O�~�jeP|���� �'5|�n�W�KL��p_�Lo�����d��\�d�d�=�W�_�j2_q���jt��ͪT�'��]á��C�����u��@c7+R�b�g2������aP��G�NG� �E�ڍ�aǯ�`o��߰�i��Q�Mt�R�%����Ӟ�R�S�*3��~���y�"0����;ѷ���=�TZ�~�G&�\�cy�����9nH���0h����!�|�������?��"1<Pa���{����s�$ζ���.���ӵ4��������:6���g��~(��TY��l���V���6nN3\Қx]vC>]���[8�'5v$5׏�>再��X�v��}A��Z���ZD
�q'\Y�=�\A�L�c&5%o�ˑOF�J�z�m�#��0lӉ�F�X�;(��y �d�	bʾP��� 	��n[/�tc���|I��v8h��B����t{=A��KC_�lgzm[�v;�ߐβ�~5���Y>�+������aUk^���n�H`=P�jK��5a��9>�Et��$}�YO�x����9��).�2������c�t����0��d\3t�R�W��9w3�1��k��#�m�RУ�XE$Hؘf�+��})m�[�#��a�� ױ@�yn�}j�.ZZ�a-�Pg2Q�B�/z����ej���I��#Ӿ<��������<r��u�c.�ƙ0�*�qM�Y��k� f�e*�1����øP�h�.����7-��H�OL:�bx��CD�r�\��t���-N�ɆhŨ8 d�ml�h�� ���W������Jb���]����S�U�dx��bBkq 0�- f��q*}��3)/;�n��Ɋ@J�6[XK�X�>9BgYj{�X\pqL$@@���>p�R�ZO�Xh;kM��U��Y��I�"8����u��)/�<'�jK�D0�����>;��U ���F1���[T����:����H�Z���r7/v=O���kz�-�]F.v�>OH�C#�Z����A��q����̫?ԇ&0�&R?�!�b���^���?;a2v�g;�#��8��ؙ~b��?��>��N��<.Y��q���9��`��f~���_4�7Y�
�q�H@�4e���H��q�4�r���|a�I"lT�G��c"��3��h��w�P�(���C���8���������j����}�D��R0�ό;������'�lf��S/�V�6�4�ԭ?-3>4b��tS�"�V��B�p�X0A���G*�����y�ej)��<��~�t���}	��K��@���pT3�^jfoa��ɼ�:s��������w���������ė��l����Z_ݶ����my�BS�(]`�_x��!�٘|4F:btk,O��`�$7���h�f/��Z��ȱR�+��@	�|���D���C�k8֎�[*�A\ó��\��0W���/��Խ3��G�J0��ҿ�#g��G^&ǋ�}�A�]��VN�~��3q���|�
��M�=O��
+�z:H纭����TC��[�����:#B�tO}0���إP�~t�ԯ���-	�C��B�!��\t
y�BkG]�N���00�a�z?o�+�>�"�y��"b;v��69�Z����O3����N<�4ؚ�m�
�3�%�3e�j����n�֍4�?������̩J/��C�e%�3�4ե�_������#�A��!��aa�nie�~�ͰZР��H�fr�J>�,
<Oy�?d�:%w�K-G9�<�0vH(Tw_@�ļ5h<o���cyvW�en'���!^�n���
D���8�}3���+㟶��n��s1�	.�Fɥ�d���taո(v&�Ф�"O�35ꎥ�����E�Ó�r�oD^��O�*�M�ݙ�瑚��� �������;�o��0���N.^���6�Rޜ��
8�QD-��}_l9�P�K!��E�tj2���@��ҏ[�#�R�ZA0J���ӧ�y̔��g7�=s�b�c���{�ݛ�)�C:#���aj����!v��Ȫ����PH��Z�r�>u~7�N���]`d��(r��G�?2(�A)%:��]�[��6���A�K���=A�&L�9w~�1�ӳ��V���>_E�/�[&J������sGQi�!	tDV��$e.�+��WK���'�>j�W��&k��mX�P?�|>��kj��?7�rm�P��N�̐/�qQm�8�{�n�������8��L�������}.׿9������G�*��#��H
 ��g),Yz�E��͸7�[I��'aJq+s���[�'�Ŷ�����&��%�8;�-H4vVK4��OJ��!���,DU]
��N�xy�&�0��k<��K�9�׿t_�q�>t�l�TH�c�Pɾb�c�{P̢Ö	��-�|U�js�11?ov m�w��ד�&�a�'&�9:����N�Q͟���M���5�UI��ԈB(B�2�获DK�M��8��HX]��������w���]���W���v)�6�<�h.=NLI�.���iO*�ַu�\�P���Е�$����Z����j)y�e�m�R��.���t��~���a�^*������eY�}���JZ�2��O}9����rXwл0?�	;�d�f}x�),n���&W�@�@���40���v�jpܯ��ަqˍn�9������񣞀zY��0{(�����v�o�vg.Dk�U��=�3Ŕ��67s�3+�v��2���m�{�3�Q�f&�̜�s�V������!,IMuɴo��Ł>u�[��3�Xz�lz��-��@���z5����8�z9��ug� �ڵ�B�>(/���j����~��@Ch '@z��1P@._}��u��z�t�s�趉T&�hn墑�
�yo����B�N�:~��$F�P���g��LO��������!c�N.�+ܤQC0�-���<�dg�x�����n-�鱶hY��
��fOK�S��>In#��3D ��1jlMM>*�`2Łt�h����V�I�6�S�&xN�E
sD�����o�5�(���[��������c�W��M��if�j�Yg�	'��>�,S�u3�j��Q�?�R0���@,Z�V#�������G&��O�L%[��{k�h����W/�~�����H��n#�/�?&jP�zN����d��ET�.��^�+T�Mx]n������5�HI6���Ɯ:\Fm��l^W����4�r�iyͼ��=�g\�WR+�LUrߒυ�QoC�W�S��ޅ~�et��\������0��nL�q<�%�Ґ8[0zo�NJ(��N,w��/��;���5�� X��O�V������7����sP���+MY�qU��Z���<�!�Yd	^&��h��+�e2��+��U��J��/�����X�*�X�8���r$��� n��������|�������E����#���ԔD��z�6����?�Fƃ�v!�/x�P� ���c����B�H�0�-��h߭��j��G`W�ܭMV./1�h��Dw?v_��2&3��޶���wk�����J]e�ķ���w�0a��h:��1��h�#�[|�B��1}�a�g�"�S5��eƖ�|r�m��^��S�BA(��Q P�oGU**H��}��o�Q\���}�>U�,���`HV,�yLeS��
�",�sP5�pd|1�@QH�,���Q����&we�0���<ʔ�n��5�����g1����``�*�1��Z��a�t��FRo	YG��>wd���+Y�҃��	���Rq��*����w-��|�x>+��d����'�;�w'��Q*9D�Ud ��1a_[Mń�Z:��/8j�
%�K��x5{�����^9N�t`�a���?���g������v�?��n>�B�ͪE���4D4[��Sm+�B��#�D��O�x�Jv�EW�q�'�� ����%ce��m�����DpQ�U��4AB?e�:@16�&z�ƅ�ޅ5��J����ka�!�LE��h��I��.�M��2�����1,�14���s
��5Z������<������2���Y�{12a*��κ�c���� �� �UP���Ѓ�ɭ��n���Մ�����D%d *����3�l�1��n���.'Xv�����|��ټ����fr�?�)���!�,��pl����`��Y�H��T����rH��� UU��C�� Q��JȔ!��X�W�S�����r�[��{)2T�=��c����`3żle���Y#ZG�V�Α:���<�ډ��&����<yb'����;�����,�7	�oC��a�L��,�7�i��,�"|�Л����3g�J�{p[(m�=��ݑ�l��DZ�j��2 �?�{Gu�}���#���% r��f>�ZE��0)��w�}S\�V�MI�����f��	|bت�
3�;TΈ��c��U8���c���"Y�`:a�k�\�Z�{ܠ�$�j��ڢ6dO�ަ���&|��O��i�}[A�2'������8IE,0X�`�Y*K�uF��^�Ay�ʘRɾOVh|rī������rM��1���J��5�àa^����YA����2M�G�p���w�0��0�N�V�*m�2QS{����d��F��i�(�OP��T(	��l�Yд�������+�U��:?ϫٴ�'�[�6H�U>p�$ۓ���z���Ξ�۹�,\y�2�E�0�C멆����RRʲ�!�G9���q�L�,y��)$C�d{�J������1�0N����W�ȓ�IDAu��I�Wh����&��W+G�z(�QX��~��7%fO��^]�C&�!3@:�� "�;z�_��d��K�j-�!|_	�����b�Bw��h��4
f��^�_X�j���KK$�]/$�ׯ�uICY�8!����5�zץȏ2�9s�d��pXL}T�pd������P	��=�Z�����}�|]N�|�7�h(ƇU�Y�K"F!W<ϐ� ������m��슩�\��ʊm�V ����H����th�`�����a���^㳚�s�eP���ȼ��ꀉk���8W����A5�D��&~�=�с�� ��ߝ��Ќv�^�#R��%e�1/h�6A���YKH˯��XL������\"�N�xa4�;F�i�b'{(tvȕ�]��jx���a%��i�I|���M�����c�$G�]}S$Vv����Z�E����Qr��VaM��[�֎�`^SC>*I�r7��[z��0رs�`��4K6�R���w���!�㍆Ա"Il0��pS�'�:l�<�0��*N�rA7�CM��i7�Ubz@����/�\h�+=�k6��Jqӝ;|�Nw����#B8Hrl:Q˶vJ��!�ہ��e��m=E7�Ϊv؏���uXƤV�?rJ�bd�̹K�S.-�yN'�5X��Q>Q�
< 3���j1;����\�TBc��%@�:.	�{#����z�������(n6�>^u,лN�r�j0)4��������@JJ��t(��QSm�&O�HC�t���j�4�hOR ��M��/��{��U��@m���
�Ї4�h�Ca�'�f1d�b�߽����'�1h'�]��^vyS����蓶"(���(-���ț��
�d���r�li���r�kHTߘ��ӋG\lΆcy\/,�܌[�]�A2��,�˾�QF����KKά�D6��ם�5,h�m6����*[7}��̀ӔT/9
[�یB��uX��6��J6-��[�����SG����~ 6�D��8��.�,���F=���p'�X��@đ�� 1�D_G�Sٜ��֡��"R�5e8��ȰnOM�S� �_]8�1�a�&�/'C�&!d����=�gL�ӆ���@(s�a�_���.��Jz�#��GZY��Q��7��������5�@�I,�|�I����
����|�����7�޻���W�նv��03J���H�eM�xg�yTs3]m�:[�L��US�;FΔ~���h��!¦T��b"�����3���`Bz��2�)rjfhhV�:g�������q$e�EJ�s�j��EY{ja���
�y>`r*��oYҶ愢l8�M�dĺ�jꞮ(�8�4����Tŧ��ݜ��S��7��Z�@�ͳ���I�O`ԑQ����{;�ϯ����񎄅�AG��2����j+�h�n瀌�}r	Y�l��M�|xB��W����2s,U"J�2�ʉ�i�������P��	�6q�M�e@P�R��Q6]�V�H�7@*C�to��-v��O�^ 4(����x�P&Y�A�"�Y�lY�|BR[�\�A�|Go�Xp
]U)�=���l��^@gm�?��Ċ�	�dj�S@E���j?�sZ�f/_Jt}�6��W'����>wZ��7��PG���<�po] �)�-�PZ�7����Uh�U�Z�$���W,�������E��c ���))>���t1L,~Fo(���x��ݧ,U��z��ٶ=�-1/>��P�m],�0@'�]T�W��Zs�M�}X�%�Y���_�;�� ���?�h�P@/��Z)�՜��?kԄ=IB8.Z�����ҏ���5:a��p��e'�Ѱ_Tt�Q����DZ�c�B�UC���
����\��aҧߟ�O�yL�;R���ˌM���~N9��S� �Y�g��.0���6��Wl�	n?C���b�/��>�B�ְ��=�ZiO�����	��|7��0�s�l�k�B��4�cacꛍ�1f�W�2f����p1� �[��h����aѽ�j�_�%��E_A��q�հ?�X� m�`�u(�A?���]��n���ӝ%�n?�y��6�~�hθN�U[w�WF���H^�H�zW��aN� � %�>ں�\���������B���g��F��kv��^���ιk�S���&3�x���.�]�a����O�3�n.j�gn�}9�ߌ�=`�U?w_BH����mo�`@�V!$O]��{�f��p��(���j�E��'8@������f+9��
�����"��4�������>u-���~Q̞�Ө��+���ɒ��*2��I��E�<FȪ�qcnH�ji�$͡ޢH����+?����F�w�_f�R8�Ἴ���R���I,��Z T�	��/ �!�����8��J1�C�����I����5��V9<�6��`�v�^���E�!X������7�\�j1^k�X�Lil�j����6\W�M����v?K9.�~ޛ�O�@I'�ᕚ����b�C����Sm�0���Y�ԊŦ�N�0<c�p�������~�o@���	�,d�PB2^���ɾbw�T9eA8-�m���`$�_]�hZ^�g���T�<¦c���{�����ȪL����(<���sg&�ӭ�d��ӹ)�!N��r�h\�U
���9uU�T;<��W+�}��u �>H���R
P�_��yVC�) �}J�ӂH�t���7BCp��Ӹ8�ۛb�a��^){��"ɯD2�J�l�(ݝA(�����^C�?�V����IG��>z��':qx&:
y�����~�$���\n=�v��� 2 ]]$�e����L��6��U擏�4\�%��"ᶜ���(�ï��I .���6F��\���"��m�����ߞ�+*����Q�U4�������4������.������'�^�ȋ��r�����Y�{����$�%	�t�G�A�2SgM�[�D��8��upż8�9LWX?�*q[@ᘦ��p��5������F��h��ա��\H�g(�Ѯ"�z�̆Cj�L[�o+��z�m�� �ȩ" �� �������(m����ޘe��&�\���,�BG�ͻR''*{"�Ң�7e�o#KGԻS����x��>zagq�H_��%�O���xp��fbI�ޣl�vv>P�� ��B���Y��;��
��P_������ �����~vnѝ�4(xs��y����K拮� ��e��h|��b[�Qu�zL.W�QA���=ev�Nr�q!z�?�����p��	DX�EzT����m�R�5��E�������Zń��-�׮}t���[��#�?f޶��{��G�AЉ�i-���D��@P��<��5% *��$�$o/X[���F� 	��� vqY�9�G�����7���{��cPjI�Q��_y�0I�Cwj͢��*�z���ܕ�2v�r���i�ƇO�PM�<k�{L�P��瓊�q�Ępf�Z�`�<�1K�C� #LV�_$�lz�A��dᗙӡ��gu�& �C�00���Jn������/��FҞL�}��I�?���qG�4��b
�OU,�mu�ä�4nH�>������LVƳ�Ab*�LQ	� �u�򿇇 {�T�j��SS�x���=g��T��:��,r՛�s{/��D1␎�o��oWo����o�;3�N� �'��bs��C=�wR_��G��<���J�+��%6��x�d����5&؅��њ�r�F�
�D27Q�z���	�`��v�"�4P���~��P48�� k|Z�8[
����ϫ�◿=L��4�۫��T6�O��C�z��.fV$��:�-�yÖ��	&oP$\��m����-�|)x��������� ݔ��4�z�e�
4[�z�]��ԃ슧$�}6�׳ Bpdyp��Jv��_��@[�H�)��N�j�-��:�ٔ�*��Ҽ��6Ҹ>��NY��G���o&/��-����1���]ak���EA�*������ �X�+<����R�Y/(mM?�N�����/���8'X��~,�'̻�)ъU�.�#�?�W���1g�MU��Zr���Jd��¹^nt��q�M��Xq��Bj�^�~��$M�h�MG��VQ ��+�������E���O�������u�����P���rj��I�!����4d��^���.6~��JĲ����eP�b(أ	��)�ׅ��^1����xق���H�M>.��U�Xf\}�����K�7]3�ߥO��i����_t��!�����.���5����:OVʬ��$�z14 @�;���=ẅ́��V��:�+���趄�$󫢦��g�Օ�Y��@�x�
/��U������ �u0� F�,@E��X��s��éw(���d�x�<m���I�kO�SR����>#�lĞ�ÿG�,ʵ쭩�A�^���5���!n@����aJ���������t�VD�b��q[��'�5�|�)؊���,m{�3a�X`Ft:��:�a�6��af��B���=�$0-�݊ٴ�Q��졣�*\mT�����F�rLѵ���j?ZK��Ùh
�QD��1��M�K�٦;,���N�`ʌW`
i-1&s~18#^�O��ƓS�)�!�K�za0�����Z�۳�rG��	$C�������A���~/�SXO.����kMpۀ'�����Q�n.Pi�öa���#*�<!n~#hl�����֔`e�]U�ח��E��(ú|���Ƥ�*u�r����ױѐ�o�ߓ�"��Y����9ȑ]6�D�6���E�Q %�N�,māDq�7����Ȫ�[��C��͌1���-`��\W��F#,sM��>M�� Ț��OQ*���p,�z�#��4S�z����V�T��P^W��r��P��[k%I��z�G��ɑ׳���Ŧ��)�܆���SY+�{u 9����*s���~(Ċ����Qd�$�Hm0w�p(I@e�(s���"�?�2��X:^�i��5a�(g=qZrW�a�1�{�����	7i�oN�P����&�ٴ������g/\�q�v̪ز�N���d
3���L��A�ݵ����ǜ?�O]t��׍�{X<�ǉ5e3]�GْctDpn}��]����yXz��U��������9���:�]��Z�-���:+3b���RnY��_t��?��ҭ���߰�V�z�b��R%�߄��^v����~�Q��LݓRbU�"�w���?/0՗�>� �hl���\�v3�H�����,e����gQ:eVZd���~��m�̄���Mӥz~�"��P��Ј-�糺s�V��/=�'�zT�쁯�`��䎟�
rn[�^OO�z7r�h��e3c%�_�4(CL�[�+Vʺ�g[j����͎�7GZ��|Ղ������͐H���K
x�ק�S�Y�!i���Y��a��\�+D�j�^s���ɬP�i	��7ཡ0�;\��^Bո�5{N������4�����	e��Ѹkֽ�0>uR��
S�}e�?y��lx����c�s��W��ĥ;� RDȨ�Qn7���Uǔ˷6/n�v��2���*Y�H7�=LS��^�X}h�{|:h�VV�>rK��M@�'l��,�N�����sŖ`m�/_W>�b.��
z�d� ?�R����C�e�1���Ҧ˩���)a��|x7P6(ԟ��?��bi� �?P[�Kc�t$��7&�YV>���{J��=^�$���v`���î���!�0�&���"�G��E�_�"{e��=�A��z��K{Xrb���2���xW���s�g<p�?�/Od��(`	d_jp5��i��q Z���� �}����m[#��d4����,d��(��hE76���J[߁
��1�H�%����P%
zϷ��9~�������� ��,(�K7FǒP��(jC��}\&7[��9&���*�����L��"n|���¼���F*��Ev	��Ӣ�X�B�5/Ţ�1�b.�"��1S��l����.7R�$KI8
Iz9w;��߉�x����?��P>�"c��qYO���Q��&O��d7����9�Lt��:�v�(Sk��?�K�d���r���s�X��"9�(��}�6����X-i�@�g��,{}��J��_�/6��1D"��J��q�[�����ujx��X� <񉉋F�΍��*J�KKm�G@�;t���v��jjt�~�xb+��m��&�ʏ�'//���b<�.p�L�F1���ʞ�9
��(Gi	�#���y�6��h�w.n��ɨ���sJ��x-eEi�0�Nw�����ض�6�u}T=+c�ݳ�t��h���:+Շ����U��d�������4	���ӒP���s�)�5"�A�O�s�=y�hǏ叁ۛ?C f�#]��M>+V��:���8���g�� L��g�2}U�ę��\���Oɓ�ɍ<$g��/���ՃF�
ۚ�B5n�B��(��8�l�U]�1N�+g�=+�X�����a#Ŵ2y��\���!iLl/�����F�&����bK�Y��_ҫ�&D�v���Cog�>�4Ƿ*�2�Ͻ�t�e	d��mN^W������(�?����0�#$;���K�Ee����88WR��VB�n�@�S�C����)D�>����;W\�k�ӔC�4H�'R
����A��#�SIAYU�F)õ�E=h��;���d�#3�u5"���5?Lk`�RF�؟�9��/ ?�6����>����e�t�;���{�bJ��Y����uF���N̂�	n$i��_u�
XF0S	�ר�}$ʹ�|ś��x��̔".)u.k��B��"\an�<-Y�"��r4>���D��G\0����n��&dџ��=�O�9�[�-�㲽��󖔪	�>x���$w}u��W�fp�C}� �y��r��,)|󔵜!�X6��h� �/h��iy?�xr������s��Aސ�֔�'�АY�ulM�<�[�#�:N��������g?��&�瀘�2tu�0 ���,�A_��pYU�a��y�~��;�[���|@6�I"Pv�ՊlX�a��Ȱ�g*]�2��ݔ�[�F8&#SU��:Uw�v\~���z�7�.#�� l�S��`&j��S����4s�O2)Nf֪�\\���_���'2�*��D�J7��� �;[y̠%�G@:�X(�;Ԁ�OK�U�tߑ����5��mB�NH��=5$a���A�p�'&���F�4���t_VC�%�;�"���9i��RS��Z�ؑ�"��hs���a�/h�c-��H�5$�b�#f���v�JW �h��$Bp�n��d'\���5 w���N<��Ka�M"�B��ǰ���o��C[��r��Qw�O�5�m�o�����&v�qi6����f��C�"m"4td�qyT�,7�@��ĩ�G�	��'�E!�hW"B�*+gu�E�o��c�)Cv�&�t��J���l���hR#x���K��.{��@Ggv���-�<(�^������X��&B�︅e �� �j�p}��\Eî2���n�G;tc$�G(b�S�q�~)�h�:ء�����s�ɜk�;��up�)�6�/_�?J�~k��J��������eѕ2�}ns�U���I�*�����߇�K� `k)흴�R��_5��2���������@hS�o�YL a��:o9x�M������?��\6�TԐ)72�0_7J{��# W٧~�b��Q#R3�a��c5�d��l&.�)?�*�_�~ /VJ�G}�1W�ÒF[���2��<��ԉyw�.���(�Z5r��;�������ZB����\IB���8Π�q��lٴ�}�0׹`�#�Y"u9��iP��q,�d�T�U����v���$g�����b��Z�uS�%�z�ߓm�V��'��V!�:���+�!�Y�r��Sb��⻛�9d�	���Eא3��p�pf9�댕��;�������Z&I$�[`P�y�k9'r �0E����$uL���#vтޕ������J�MCjB��07�At��z�����q�ӠG)�'>�}pz�&kLw��<���N
���� ���. �@�C(�qPT��� ���sf��{�BN���0'Utٻ-�!tYV���F���8DN�z�:���%�n����B^��a7� �t[�V���m�Cd���#���o"�B�p��'W+�fd��җo�I�_�Y��ێkGx�H�6C ղ���Oƾ;� %��&�|�7F�ݳ�X>��1��2Y�ֈ��� P�_�G&�|�����Q�O3�/z�QBw��8e��h��F@Qa��@���t�ZZt����]���6��pܴfq-ٚ �61���x�BȄ�5�
j���E
��̎�=wE��+�QqQ�j�(�ۂ@7X���}m��_��%픫�쩯��#ׅ��*։���7mx]q� C%��Eih�;G�xe�p
�����k���9�zr�SYM�rCM��qc��N� �v�+�Qa|ȗ��.\�s[8CTZ�IЅ�;�ee)NGw�>��7����>��D"��o��j�O��۩0������V�26>��aM�{��l�s��%QѨF��4)�T�ś���4ӸI{ e}� �j�����K nY�9,+|�a�%���7E�6Y|6�]=����WWe=�؞\HaT�{l�ҋ�f~��N�_��/���)$�k�1N��
�c���d��zZݙ�s��W���L�rc��S3����������v�[kcU��H��Щ|8����ο�jB�(��d�1��������2z2����P"'0�{�A�����J\�}��W?/o�'�f�W��95e�-�0R�
�/Y��@��Mz@��k�_��+�7hv��*5���O�]n�L�U�a�K��011�O����o��!��s=+���d�N��g� ��9���O^ȉjwp�e=$�`���o�]�-!+���M����~�"O�?���!�*Xgja��dK�W �mw���za��gHf�����-}���{��lU��v�5#�E��� �!�ԂǤK�>��i������P��t�ֳ)?ac�6G౵��I�[�'5H�
�}�Y�8|��e��dW���䡕�L�x� ��w5���I�s��(s�<XRMg�W�:	�+�Ό�F�k�ݴ�Q	
Jhh��283U3DH���9*bn���v�ث=|`ޅ�������Nf�^����ZЖ�P��!��!P�=)�	� w�gK�1��kY��B#-F)f��[s��⑌FL~0�v����Q��+�r�A�z�����J��}��˿ �¤���-k(S���^��AJ[��vdM�^XK4�v�2�qY1�tX�Y�U���\��Y��*�Ex~�BL��P\�1ۢg���-�1`e�Ê i2DW��E.�]�3T6�RN�qg�	�4�S�g�=`������1M�nq�GE��>�y0E-��*��.��~�H��5��<���P����z|e띣���(v[��W2%<�����UM-\�a(/����/�Ú:s����2�^&7�mb#�w��;�
�W|�3ͬ�"�]�wu��vjE���"�rkC�HV�k9����#�;G�7��n��S�_T$�U�"Qr�RXB3Rqŀ5ljNΘ��$GA,���"�wT�V�4��ͷ>O��T�_y����žFVڨ�_^���4l��eR@�%_��K6{�/*S2�%l�@�ϟu+�g��6�w;3hA7@��5�w���3������%�{v�]�����0S}�{��e�N9AJ@"�
�YARl52�Gy�㍎2�/K7�
QR6��t'nMP3wV�Y�8ӥ�ܧ:gS��VIH���b�)c�<�����(
��yZ�cQG}�Zz��6�	$hօLi�� N<
��>/�nhxmɘ��{)j���� ��-��w"��ߛy��D{`���sc��^��q����xפ�F��.�S z5�;�ZZN4n�1����Շcu"�U	����b!���� ��/M��6��u�ԏ�v�u��ەi�����)�:��R_�����@��2}�@E���-9��������G�t2��Y�ӼiRV�h���I	�l]g<f��D�*$}FBW:؍ąެ߿�,T!��K>K�?�Vr��n���|��[|��]�&��ͤ��k	Ks����4�^V���
�U=<�ĦfDp�8h�;�CQ�l��T�)�w�&��K�%�R�l)/��{�G��V%�)�$?��QYC�I�%9E }"��L�o��2[QM�u>�IJ�{��nc�4�v�X���'(��X���a=�Ls�46����]PO\z&]���y盅��������^s#��OF�����'	0���Ǡ%�������(��A�~�ci�:�>%eր�`�y���B�u�%�����*(�	O0fn���2��p�y��&˽��g��|V�1�����|�,�m�X���̔>0T��2M4�07"��0,�R�v�­_j)!���0�(d�;�o/�-���\=���=9��Da��Ξ��[Q�s#YBY�H���b��9���Q�l��~���Q��g�[J�-9r�8�)l��HGn�|����f��ćp5�,�b%�m$]��r�&H������i��[_�4��A_Qj�*�=4b }�����Ke�vI�X	塠��V��%������O�̈́���$UU���y΄�m.��D��Xp���3��6fo��9"<���.S�K%�B��C�z��y�6�7qF��ʯ�n�S�M���]����͚�o��j�X�Q"N��"\�C&��G�ݨ�*��_��VǺ���R%��t�!a�Pfi[�U_i$�#���Me���X��� ��;�iD����H��i5�^` �ۍ^VEQ�/Eb"�{�э����kĝ�� 0�/�Јh�oE\d�Us�6^��Q&�a�a�|#�eY�쟕�\%ș�r_��@�1'�7;����Ǵ�<?i�.�}�Ϊ���V�8^��Nvֹ���!�+��ɰ��ׁ]]<f��z~�J�w.�ka���Jb�!4,���gp7�S�=����әB[�G�k��[�p�lv��P�T���c�
���!�(M���*�Tn����S�M�����.��+�=="3iK��8 5F������Ê��Vzڈ�+�C��B�n�[}a`���Đ�|A7���`�-�p�j-4 ���n$ZR�kb����	�h.B��T5����ɫ�Kq��-�1�3x+�Wh.�<��u#�o�������Ӈ�����q������*� /�+�w������_�Nme��5��IY�Њ����]����bN[g�-}��3o�P*��UA�S���َz_ ��>�U��[�Zu.{?خ��˧��c��f�m�\�^;�6��������|�E�Ǽ�0����R蹰qe��ٖQ��j�}�Z��	�J�J�_LhU�-��>� �l���X�����Ԃ��E,�����Y�G�s�ٝvKq>� ��|�f�\+�9�$}S;�&��N���rb�l�mIh�	���!W��
����G=��~��-���jW��wh�du\�Y�)��A��0��L(��0X8�l�q&{6?d8���:D���i%�Ֆ�U�1i�j��ْV1*��#����֝�cp�|[�O�]d}�A�N�x��,W!ͧʌ�SZ'E��/�8���������E$8%���*EJnb���<����q��ZAKTy��]�����ů	�P:I��s�]�~0��fr������y��ƃ�-Wlu��k��mg^)H�Lq���bzr�R�������Q�t.����>���y�/7q�M�η3~�����Ðd�ze髰��������E��+�Q�����
�8��D+�X���U���y7w�#��x�>[VN��h�Hߺjl����y�$A'�o��Q_�oၵt2�i�Ȁ �q�}�}�ұ@o��n��M+�3Ft��ʾ���(9g))�5R��/��)~��<>�A-I��నM�1lf/�c>+et��?"#��!�Dy�}�X3��k5-�s\��p���&[�A����A��n�F��5�ID�yW
�^��)���i.�t�j��ǥG����A�ܵ�P�ٵt9��P@~�U�s	�d�i�߁�Q����X(w��q8԰��O���9qDZ�Wu�`c!�1f�o�#��lX�Y�����%��Y����߰��Ӵ#v�
_/tHCT��@�Pe}M
��&juHbC��f{����Ș�����T.����N���k���rJ�>/�P��������共VN��ϗF^epqr��pU��G�^�E���cA�L8���.-��,�?��Y}��G�m�d��+�
���1���*�>Zl���8���2R�	P����b�/ds"f���O��H��ʢ�*4& D����"�����9����c[���JR� �+&��i����r�BO����J*�u�RH����~2��N�����s)#�MZ;������z`+������_-�]��ݍ<6��S���oʖ�_+F��ou4�S儣�b�H�[p���[!Õ�S�R�@�sIUi5�ܐj�7�!Ǡ9ݟb�m)�(����O^�ץ�^vNO���PNO� ���!�b8��#RO��px�Z_)�*h6������GRM��Q�*��s� -�|Z^X.8�oG�lJ{�#�A��Ͳ^5��NԊ��m�N��0��������x���.(T{x��*�x�m���d*�u ��ݣe�3���ѕ��f��������ad��8f��2�C00a�h���=�U�[�P�!|hMl\h���:�����e���3>���o�l�d
⿷=F��`!G��|y��m����oS�V�/]k�;F�΃����a��}O;ޑ�_iW��{������I/�|d���a�+2i�f��'/=n�9��%�9��F�>����/���]��aݶ�ҹ�6��V�HNZ�5��'��tg�J�����]���� �Bep���1����	�A��2y�Mq��n��.�������(dC��M{�6ȍ��/w!��G���g7�)6�!����'����0�t~���Sk$���Dc��{�n)�|�?AA)<���@�y
����V� �s����zO����)���l���q�O����(ǖ�V�zP:'^�)��>�Ao�ϰj[��@��&o��R�) �,�5��6W����`�X<5�R����D���Ѯ��e�����e�O�A�=��T'�5sf���a�i���uG�O��G�k�_�ڰ�A,���n,��Ke�/R����p�B�9 qB�b���/'<ap�5�V>_�pk\�a͹�F�2h�G� �����ӋW��g{-j,Ϙj�e�2�EE�U| ~^� j���Q�AQ&+�`�X��$8�-.{�Z�1�c͂�\*q��%?�*b�D����C� �>"�,�.���/���fl2]B��:�^ �����Ho�\�5r��dܕ�8��ª��Y"�Py0X��=܉H��ˮ��\�1���Ld��~����9{��S��mD�~x��bi!��ƋE�ӕd�Bjm���y#���$�������B�P���7

V��g�������h�������#k˩��Ng�p�"R/��.v���u�h��⛗����ŢQ�����K9=��[�W� �Fz��]�&�C����d؝�i'9z�|VBH����2CIiF!C�
%���`'_H�f�CΉ2��D�f���v���:��7��~�q�8�TM��;��#�	q��^i~A|�K,�ٍ'�X�P�s;�� �Bm}�A����)�I#$U�Y�o�jn(�K��� ���O��@@�����Zon�R#=��rz����2�ͼ�| �"��൵��k�I(��R�V��>I�p|��,���D�m
������:��.&�����Jf�.Zj�a��fQY������FA�X��/kX>����K5C넉��..i��W�>�\D��b��-��o�����Յ��1?mf/S�فe��(���J�p+_ш����C]t21�c��\PK��q�.[��|�Qȧ��;_�~��l��R�AthU0�\%���<Ho�H��n��q��z����H�˗J��I�v~�̑�kF���I��5y�q��X�Ak��t
v������R���=�C哷�y^O#���/i����x�jF ��H�4�u�}!8� ��2��	b����]�������K�k�B#�8"�������mrW�s_Mo�tGx�d����h(�LR��؉� ��/��*a�e�o����C��fꞢDg܇|���s����5$.��_(r����B�9�O`���ʠ��ة�,�-߶)�I�$zuP/��P� ڦ���u{mp{w��=XC��% Cr�\�䳔����:J��'G�l���W%�$�z~�SBQ�d�.b���&����@Y�>��/R�A5�m��?�͖��ן��R�OX�	F�ȱ`N�j1����C����/�y'�����n��T-|�o�a����g���q_{� ����XJsL��|�{F�h�m��ޅ�4��(�(˞��4Q�v:XN�z����I�%X�~�����~��A�uC��8�u?G�sX�^ӯ��ajFG�7��O��y:���7���B�����z��g��j�����a\aJ]�ּ��*f���Ei�cb��ox�F=���l�٫:&�Ŀ*;I�iO�I�8x��ʔ��Dk�Dn�,�UA�!�5�ZN�엨� �s�ad���,�����g8ڛ���7,��^r],j��A��%�i�8�`�[���<��-ޗ���@ͭ����7��$}e���W�~��<9��6���(4e� �A��#oSl�$ѩ�\��:��(<G��_'x �H1����yҏ{;�Q�0lb"-<(�ZsA�s�y?ƺT�� �ٰ�X��[u<%!H�`J�܍9,�&���+:E9��yh+�Y�=���!7�zhO����K�J�߬>6�<���G�)yr(�9�)������b �>���Љ�fݚ�f�W�=zHȚ�a�@�ŵ�L��#�Rm'[�Z���nlN60ѿz�s�CД����<n�l�j�-����b1�����o� W�8�����pL
GL�����L���qn>���]b��(�+@�<�%�h�N�!�\'Km~����g)(C�*��J:+X�Z\&�fv)���SXt4&�ʟ�W�ǃ��4�\��VD��g*UR�)�_H����D'�g���}���6�<�ݱX%mD7�;�<�4Q�|f��F'���f)�s{h[)��㍮�����+>a���t�,���i�&��2�uEj�#.%�C<,�[+GhyS}U�F��Y/�V0s+������>�Xilq��a���3�.W��#:7�z㺢y��כ�p��{v��k��]w��ݻ����ːR��|"�(�^7�h���=��wxO�=3��� �@��Q�zeg���UwO ���Fj������Q��;��|p2i�&a鱪�n^sTF�?�n)�iAJÌ�Q�P4���g��Δ[�~Ҕ��^q�J��)� g��ש�]9A�s2E��w�������dܺ��x��y�I�>���['�К:�����qy&�F��"�SHQ��S_�1�
^p?v�� ����r���!���s
>Y<j��/�Rh۴u"����mKj���uR�ͳ�H���s�+��r;�Ĳ��pwK7�hc��N��߫>��h���;R���!.���mt�O!�j���༝x��dP�N�Xե��'��﹄�L���{�����S���F�b�q�`MH4)�OD���@�ֽؓ<��2�3��zܟ]M�γ<�,.ϑ[h�h����k �����s[[W�w�ɾ!#B��O�����F� m�s=d�y��	t���2�?�!Z�a�z7�g�Ω�5U�������l� W�N����RT����)����(z��ӑ� ��|������N��Řk�t	1ܷyѡ���wR���v�Y�7K�����♅F�]�ͦ� !���P��;$�9�'�z���A�#%"8�qW�$�v'��բ�����f�P��f��¿W���MK��H��ၳG�E3���~וՐ�O`���Hab��I��)�-0)�?��ܸ*�A
P�L>9g��)}�3a��}�Ыp��V�!+�d�B��:�t2�$�v�?D~w��ڊS'E�rsJ�ų��GW�>�&Y;E�� @�X�6��a�s֦+��H��7j�%����+�7kɒ�\��s֪�J�+
�k�J-�z�I�Y�P)�R�.��o�������*ELF���)@n
�Oz2�O�!ep󟩆ai�������z>�Ok�R�~�{G�>��YX�gy&����&��sϵI	~��m�"n�t�:���Lw��$���j�i�Ge������\.��
d�3���.6Kg�,�4�Y�F_[7ڟ�q��H-��R)�Ig \�4W�p�A^g_ݾ��F�ʷ��#�8��HU@�`�bQ_��	4'>�%e�_�(k����t��!z;<��$�cw���	�Lft��a��Kg�ۢ"bռ�}v__ ����������B� 63�.v����p�\ab����5�пI	$�22��k��[��A�,��t�ډ���y�fD˛�Jw$n�d��#^�M�<2)�
���L� :�)��F����c�M��'� ��ܻ�*�,�ɲ[����vuoD͜�0�停��F�Gt�=�^��ئ(t[�>�Re?D����(�����Y�đ����<q|��x{!C�W�.,�?f�G��΋25.���B�\�÷M�9^�h+�ԉ�;��E��X��m`U���̲?�
U�	��*
y]ɚ}h[��_)::m?���P��|�=u�s
,
�s�_W:�q�g�+5$\� R�^w��P��f��V�)+hE�,���-�.3�Bh@h�R9����M�Wa���<ЖĮ/��M�0�t��e���uu�H�PMn�]�R�#��Z9�H	+Xd�������Ɉ�uV.�`�-���k��r��P�����V����1NȮc<�-ľ
?�fZ����+��zk�BZ�~�P�i����@����oS�<�D@O[��pJ���̊��=�tiEV!{�$�/��O3�%ԙL��#
6h*%ًa5���sFK<+v�خ*m*a��j���}r�f^�I�h�I�ȉ/k�EXjd>�pϩ�$�}��b�T�}M���0O���B���`QP!JX�������?vHT+�T�c�n�B��P�F�'Z�ѥ����G���A�{DЩ9M)�s��(����ŐC�z�:j��������P�Y��nL[�/� �fu�oY�4�eu��d�#�,qù�~S�E��fT���Lx+�S&1D��AH�]���^�����	b2����SQQο�7IF����^s^Pf�0����v���:W��*���5t'9a�m3X�hc;pvJ����2[����,(�b	��z�zm;���
��ԅ�fsM��U�:�KG�� M�W�,'W���t�R���"��Ӌ�k���ȕֳ�H�ʲ!���g��Z헐	a�9o��q�(���
w��p�������=�LAVt�Z��$������)<+��vT	N?w2o�?�J����i���=(���x�����2,fA�]�%�U&�q�R�#ԔW�=�K���ksA�]G���EU)$3V��@D�z��!*��\�x��;�^�����b�+FY���T��җ��\�1� ����}�F3�zc�N��O�-��k�D�`@\(�d3V�L � Q�*C�A'�����Q`��.^�B	l�uy ��8��|�iH؄��⥫��Y���������߇��T�ƙ�D�i�A&v��Uu��
��Pӗ3>�B��.�:C���m���@2�K��nר����l�)�r7l��LB�2(�+n Wo��t�Ǉ+�E��g���InW#��������;K��,���[�f-���� Y�cʰ|l�Ɯ��q+�`�%Gxy�MQ�`�!���&�@���r&a �8��:�P}K��p��	�\�<9�,D�UZ�i�|?3#�v~%C�M+U�e5���2+x��}4�N#� ��D� ܃L!$��%3��b�M�C�pы<o O��� ���Gb ��N���ެ��`��S��Z�$�#����);PƼ����r�Ȳe�
�9�̂ ��<�m� ��;c��(�U�"��g�/h��qJFp߃A㯐��!��2�6�����{�46���e���Z.�����w%�Ww�?���N(1�w��yeS���YM�M]�9�N�M�.C8m]�����9U���T�DW� e��t0Pῧ�	�A%�(3*�(���C�Aѳ^��$�Z8Q#G�c�oV �����Vw0M��B.���^�gh�~��b�P� $��i` �l���@ 8o��8���ߴ��[�S���`צ+p�Se�F����[B�;ک��`BF�/�Yj�̿٨4'{ζ�z#4=T��ܴ����qMy:.����3����&}��>�w���`�x�@�;�+�U�q�dWwLr�'�D��1r��]ɖ)s�$4$��8��B�0�X�<�L�*0���X����N�Q�2�a4^��]� o��&;�IV��>�&(�}_���ً�S��^�c-}�;?+�֒!_��4|Oc�`J�Ѧ�z*�~?$��r��g}��`���\,A�sW<�V((�����N�3��BNv���[-���K���2H���09;�J�u։L�^�N��������5�b蟙f<�bd��^l4�k:�^\&�eh)�q�%�V�K�m�P�e��
p�J���(n���8�2K|<S�q%J��"�@4�Ic#w�5�e�71٭Q'�t���8�-��e& �~��@$�ȣH�iZ��2�Q����u�ZFB�UE��Ց�v.���V�H��U���$v)4Q��,�~quW�'�9<�&�G�B��"��˫�dk����\>&G�z߼j́�.�w|S|���2�Q���а�8����܀�����0�60�~NHB:�r�"�F�I^�wm�-���?)y������>� �2��XC��
-^��>�h$Sk]��
���{�#�=1�H�u��ۏ������t���s�?W���.D�Z3;D�x�7+G'��к�`GV��U�w�$�P<z*����zy�[�j˪O��t�W��X����k� "[�#�o?-ІW`Y��|��͜r�`z����]V��|��|��2s.��c[?4��4���;�NӋ
!��P;1Z7ֹ÷��2�{'88o8�����ͥ����Ef�1�*��fYa�%��9�xT꥜�J�{{�&uT�P�ov4e԰��az���+�]m:�&��!B�j��"��KN�C:�M�|oq�Uj�	����k\�M���w���ЇR/-2�~��Db��e1蜼�����5����G�5��Č�t�,AU���켼з��C����J^ӣ@-���51ȏ�3�bG�Ӊ�ik�����X�M;i��qҨ�;z���uMN���_N���p�M�����{�Rt&WWAgd��'�ѻ�=k���کu~l�����C?�p��;u�?�2�>˳B6� �Ӌ1��%VU�������AF����C?�"Y7�qj:�y��������3I�r�+�-���M-����(a�̋�J�fe��D��k��D}Y���S>āR��T"�#C'qo�=���{U�zy�%��:J�d�oS�ue������J��qy�]�X�C<��1Z��p�n՘*V0-��X���<�S����]\����e��[�g(HwVjc���}鰵e��m'�ե��ԧ<��h�޲�ж$�34�M-�8�C���&���{�G�3pMc#)��\n�9RBL����7o��"U�uH��"%y�bi��Ix�Q�aha�6��p�S)�Ke�.G���\>
�ry��7:�(��u�����+������v���X�]���=.�s��u�B�&�]J���Ua6��C���'��}˂K��=���u���14m��q�6�K0F�#%D<�' ��B3�Ub(�j:�9�zWhR���;kG�yy����(Va֌`0m�'��"å����M,��E�e�Tc%����7�F��N�s}�F��=�_���w�c����o��S1�4����-m���4%�c�S���+U��-B��/��=�z���O,����eB�Q��
��i|��ާ�u2E����lL�W��9��=m8{v
w���+�L13�ET�b�oZu���=����$�A���c�s�ѓÆ��W�ƛ���VF�&�_�P�^Ŗm��$��N��[b����.4��b�+�R�����s�s|J����a��f0����4ts�b*�T&FQ�;���M�}���y�裕�a� B���2��aOxR���4��d���x
	�_��׾��t���灎���ޣU�Z`����Z�(���!��rR�6~m��tZ�y�4<%69qۘP��	E��(5�/��|I�r5{�"���5�aa�E�n�擻*�_�> �GX��7����'4ɚ��r�I5����h�3��ջ{��TO$#q�\�_�Z.�����%�g�b^��ֆH��敱�Ë0�X=����"���?8���
F��0�v?b�e��p�'�ր �� hm��
T��`䰻:�`�1+G]1G&�+ɑ�� .�����,x��G��Vd���h�l��7��ձ���p�a-g�SpLk(�����۽�ia����*@�2ꌮ�e�,��r<;�ꇢ���4ה��d�Pw��dfg�4��w�&Ǌ�P_�lu������RG������A��B㘛0��t�:g�����;�V�Y.־����6�!0��j���/b����;I��,<�f]���%��m�:��p��_�0�J+� =%=��鹑 �u��nQ�ȏĢ���N1��oᛥ�ɡz�3j����][>�E�p��H�j��	F�'�2����C��S�2�4֭T��0>��h��������Cͧ�܋��4��o��1"_���xŃ0�W�%#�Q��^/�v����;�Sț�t�!L`�V徠	��n����a�ٸ���	�UQdA�y�k��x�'q٥#DGP�	��i ��a��%^0c���A�J�*d�U�tc��B�w;gn���� W��\���遚YJ����W-g�C�&��2��߄�cf=�r{cv����O���Y�l�`�W�~Q͞�"����31u���(�0~q�&�%�Ǹ������(�C��_�|�UW���Ԧ )Ӌ���AoLH��M���[V��r�|x�o��k����OXq1�6585J)��0R����+#�Ư�Xj��_��Q�J\��.%j��>�QZ@�NF�e\����Z���K�x��&�V�d����`Jf�"IL�Bgv��Ǖ%��{wHx���[���s���:��������spX�ai�n�٣5����K֏{�Oa��>��fvv�=Z*!�[_>W�9n�&��uy__��۵u�T�_������� a���K�Z~�����u�$/�yk�R�Y1p����Q�_�@Rc|���*;:bg�ɼ�������T3�f�^޷b�[wӭ`p������X֌ʧ�in^;+�Ďj�iY@������z�4	3�h�n�N�Y��Q2�1���k����Kč-���E{=�#q>P�2�����z�K��W�B��N	0����0�-�s�^N6���qb&2r����y�!�9B׽qؙ���@|���;*#9��H&x�$��mM���C6�� ��<)p��^Ǜe_W(�>�`]�~�s�n.���`NI�����s�fM(iU��j���~mEn�%�;ɋl^`�A���N�#��q.�g��
���� �ar��Lήzנ����vӔ���ڃ}�<�
���1���Mm�+Kg���CN�"^�������m���CT2����|��cZ�����'��ZXo��_/�h�c�	�sݏ�~���4>xA���v������|:v�&\G�������jV�[n��h�I0z��X�/!dk�K_�p��M1�� �SZ:�PR5���>�E�I6�^<-�j�F�(��'����T�d��8N~�Ð(���k'�v��[��vN�2�Cd��V��j�Pp�֓}/��H+֢�����e��vP]�F]�\~
i!9�A���o��(���|@}���^"���3%K�@��lr՝����:��Lؑ���x˹lG�-�e�2��sHj#�l�)�!��͙��6�~�Ȭ�F��5���;�&�b���@�׃7,_��k):��M������Y~�|N7��z���W����>�j��v��a"4���X*@�o�R]D2�Uk��+wE[�M#�
��p]��V���\��=���Aw��������{TM�giXxė�J@�;�}Xʜ󓂍ݴ@y�a������|g�ٯ ����	��J�;t������ya9�q]q���_/�ўDt�Bw�d�������K�GǎɑO��j�uk#���G�d�
�{�٘�wk�\:5!��4@3d���P=���5�4<�W��{���o�k]5»|?�p���>˖�7�9��R�!m��e������P�l�v;w��C@��N
sF_��@�s@�DG�߯	B�p)�S�0c���Pe���>'��.'x 6haY#.ob|7n��6�m�acT|���C�`Qa�3V���4��*�oD/�Vm:�[d�)��?\RV��slc6��26��v��̓�'��pSl}�N����E��AA�_x��_C2⤇=9d���¶�����#ς����e���W��M���qGl$�Q���%�.���?.`� ,V���Ӱx��gU
WcGRŸ���y���]��RɝN����v��0���SRDDYd�3�/*r�_ �Z�����;
q] Aʨ�l	Ƣ=ޠ����<�vތ��P�/<*�W�^�پ��	B��թ�K�&�F��Մ��-/b�K�
^a� ��,�5�W"ZJ*�G�(#0����1��*4�^��N��1�gE-얝�ib<>�P�kjP�Q�
ᆓ���*ړ���xH~���^����u)�D�! �[�4�8�{W�.�Ď�\]_({�{4zE���!�[H.,���ea;6m(D��������^r��Ĭ~���� ��5J"�SY96UvO����|��D����������:13-�Rh$z���4k� ���5�g_$-;˹�P\	H�N�7��/��2��2ne�}f+��)�}�c*V��XNK�$���=�oC�A;䇞���`���{��ǱL����v��(u/,Ͽ�g$ǡxBK�	�0��ș����/3��*>��)�n��Tl���R�IϠDY���*L��#�]Ƞ���3����e
���j��TN(\)���\�+�{���U ތ`���E�;��D3ma/P�;v5���	첔�4@���UQ=��!�u��9ā�P%���?�{�:D���7v�2.��L=x&��L�x{zu(��P&�5xV���1�_�ˎd��@�|�7���&�v�
�^a��d_'���:�"�J0(V߼k�1pR`W*�y>N1㕴/�!iU�nbh�d�,6���-���s��Hs���ΪC�β��	�kG~�C&��^Ȭkb����S�֑H�x8us� �z�e��i�y��3ex�ج�P7�d�眰���y�A����1��B�я�OFɸ��mC�<��Dje�W��ڈX��/�a��U\W�H�m����M�\V�W˄O�������D��_���Q���QX�e�9w,Ͱ�=�.��D;�F똣�rhň�ef������mPy�xl��Ĕ%vE���U�
$˲�羚��Ԁb���1����;\�_�q��d�=�K��):FWOy�j�3�*p���[��	$�#��ݕ;��_4�1:R9wcx��f	*��8	��̞������$��Q���0�G4­ �Qv	(�Nc�+����T����� �����F(!�Q��@��U�� ����޷�YG~��u��x#��aLɁ�����W"��AM�B���_���_�i��|n����jy8����m��]���01�8j�<�a�>س ��ba�z��I ��8��6���U��dg@�ep#6���ᒀ�ad��5ár��W��]�/_wsF��+�ho2N��=X;@%�#�e>Ԏ���=����<mV��'�wl�˃t)�����v���6���usf��2.8o��$_Ɓ�-/S�?��o�cIR�}��Ԛ����k�'�����Lk�)��L��C��������-J����D����Д�`�d���ߛ��4n���<�~A��&������|����������2n�ܩ6�+D����iTM��R�}<���;����C⁑�@P,��B��`�����+I~�78�з�3�	|«���=*˯?�$�a��u���^�X�.���ڷ������� �o-��C_�ȉ��s,�ݾp�W�>��	��R^�	�X���������ޒ%��"�&�/�2�.���IRާ�]��a![�*����7^�汤٬��+�x|c�v��&I�މﵡ�͠V� D�X�+�#�d�C��~�z�@7�A80$z�5�k76�>ԏ��O�;�=x��I����=���ax�v6��3�Oċ2y�,���B�p��!?X�u鋗>��"S������z�J������5:�-
W��;6�5�k�bv~΢G����"7����9%��p��ZC�cpe�X�ߘ@��TY���pK���������ƙd�ޯ���x)�uI�g��#�-��S�?�U��/���˗4�G�����h��Z�Z�����2Rz��
,���c�Y�3�0D�:{�bJ�`�Ģ�( &>�֗WH��Ӷ���	��(Mo�j�w��(��=oY\�i���M-J��z8�Ǎ�/�2��󭅘ɶ�8��筑��۹�|�I|[j���`��a4�+g�(�-I�_HF�}�ꍭ�̸�O����?h$�vy��K�Y&����ϝ�L�g����`%��1A�hT"KÙ�)K�M��5q*Gi�ds>!=y�ͧ�O6<gƤ�����3��o�ͨ�`�������TҼ[ށ��JT��|}�Q\`>1n�y����[�	���
{��6-]��5rl��L�/�OE�y���IOd� ���`�ˆx������6wh�%R��%��+-)��,b�t�Ok�x@�n;�3�i5����KQcs��z�$��Lw��H�E�U�0C�[~�"���!�.E|1^��!��v+�HtE%,B��$�Co���{K5��Y��ϩ��Y�l�G�m��1V��V�|zA3��~yA�I��V�X\��؟��$��qhr�B����ʱ�؉�p!� U�\b�|�J[���*z�	�i����׼�	��v�63�5�f=�@l�+٧�|v������d�^J{��_�`��r'�9�!*fWaB�?�+.W�M͡6�.k�k�q=��R�3��BͿ�XǶ��V��W�:|؆�������0ƣ���xG̚�$����pxjX7�/��p\e����ģ�(w'�(t��22@��M�W�p���Dթ���΃Mਫ਼~R�:��َ���uŢr<��E8���@c�ߚafYS�Yݩ�9�:��,P���v����x?.�?�f:Q�����Yj��7���N|�Y�c tQ�v��Wsn�3��V�O�^,�N�n�ƻ���Oq��9��_m�9�Z����N�#�-Ǟ�������{O�R�Z�y��cE�N�Q-��_���~�!��o*��B�O��f�_H���%N�۾�C?��+�ȟM�ei�ȁ��W@'rZ�FW��v��d��!�T�g�y7T<�lM���b�?Xӫ�R�g�����l+���y���w���8>[����ܛH<�;��]VQ��"�E%#�Ҳ��������H���n���7 �F�3=_��9/���pU���Z�6U5v�x,��I�+$ca{^�K�0�$��:�¡������'�˻z&?��{@\-��xZ�����S�e��_*Z�'��y��A�W�Z���$%��w΀�݊Ad�=9y_W���4i�)6r��Ҿ�pݯ2��p�S�1�lmu���mq���[ZFu�ẛ�����^C���(}��	�c���=�x9��0���&�K���hjq͢Lƕ%xA��lӯ���N���S� ����m�T�����6X`BП�zz�wk-���v�ld�ճ�)�?4Ӵ`�~���j/m']9��r� �*�еsa�_W=m	�Z��;�`5�,�OzR�T��'$KnMw.ӈ����S6\���e!^Q6�cC��%�Mst���5_�(k�ԔK��W��m�J��0b�L�˫��~l|CA2������|��B�7���65z�g֧��REKv��npQ� �H#�dKR'�V��]����d�	$�c��(�4�!��S�)�5�X��d������x(���X�u�n7��N�1р����䔡w�H��q��-�������w�� �8Q�I��l�cr�	�v��>����­*�@id��#���]�k��>�����<�]X7��!��[5�&IaqHe���D��(ѱ�a��4���F5sq��N���l>N7���Wjh����4|si���B*��,�mS}tn�~��췽r
�Qw ق�f�9�E��猥����Si#|&�jG��Gu��=
Tj;g����^�:e\}%2��هT��M�qA��d�+GGV?K�x��Y)�� )G�t|��#�8��.��y�Zm����&󲆻��-�vi�t7�9�A�ʨ����V�^RM�?�޳K&�yL���9 �2���u8ȏ���F���n�Co����.���oE2/���e�g�.�^���������/[����lBi���6��kZ��"~��P�f���7�2X�W~�UXP�%��Ľma�m�'A��"z0��	yM|կd\�gI
X��!�+���䮃T��>�:�&�X$�`}i��5����T�	أ�"�s�K Dv�3�b�0�n�vkg��0�,�S�Q��I#wJ\J|�������"V�mS(c��a�f���/�G_�HF�QW��Y�;�I��C�M��(�9I���['��΋��`)Y������a��:�ı��W�j;S�	���t����G?�ۧ������E&aLFH�fVI�]p�\���3�D���������a��[��A�O�Q��J4�&��>��"]�12E��d�(��ٿ>���Wx�V@s�z��yB����>�𔻟:
���ȧ��IY�φ��k���uY�A8�r<�B����`c�W��m��+�so��@-X���K3�,vJ���w
�6k�� i���̏�����K6,on���f�3�Q�u-G���$jq�5e7���G�2|UܸHշH��¸Bݧr!h��Gh������W*%���^�ύ<�'�	]��/�c
y�%��礛�(
۹���0��8�T}"^# ��z��F�d���o��,ϵ�P�?y�8T���
�q:�i��r,�a�Z�O����L{@��<e���!!Vk5c_����]8�G�����8�2���~m�d�y	lt8�N������򻅆�����F�x���9/��^N:�j�]���Z����9z�y�'���B���<�lb�Zne@?jSz��xF����6����yQa��+��o�H���)f�L�G�������Z�g|�����ͽ ��|,b���[��9�����`�5znL�6�*�:�����Ѐ�N�L|s��VW���K�-ڪے�p���y��{5iUH��,Z؛��u܍[�'"Ù�9(")����뮌
V�aI��]� ѴU��	[+4�{G���|�3"�XEL1~��#�d��ȓGw�G���w����5j�{���l��hb�����C-t /�CJ̍Y6�K(a���y_SN~��Es7�!��g���.����ގ�ޜ`�n�@PŹ�	I��m����?j���hA��G�t�v�[-�+H��,�:������8��l��\ܕ�
z_��`�)�I16c$:@-��f^���G�_~p`�f��i���1̴����\���{ٗ>|��2i [ѷޖ��#:v�'P�h�R��L\���HD.�ۋb�� ]��c[� <�J�p���HW�*�:7�i_��f,;�N�aѫQ��B�X��/�\(�"#�Z��r5f��N�,��V�����sI�,}^Ň;`�nS�U�.� ��|�Ɂ�`��lW�|��M�g;\��@ow�<���3�@���L��$�	�le������,��D\���5�5AL�.�ʟ�]?+M��KFh�N�ʑ䉁�ua�ɽ��L��=��%u��Y`WW[H��.O�ln�MU�ʖn�K��r����L�=�k/�]O��h2+�-O|��ë�B�j�* ���of��{�hm�k��|9�v�/J��a��gb瞋H|c������F�\ ��s�<�OsMɦ:x�g�s�[��B)�H�1\5��~������֣�鱩{ߑl��_���p��q�.���636��i��ֻ�����4=�qꄃ�{�6נK�[42��s{I~Ԫ��'dM��!���Q<�l��g���l�����5h3��.��Z�ӍJ5x���� �غm���A�rGcm��u�i+�A������H�DJ[�A�]��İ��1�������
Wi�؉PƸ�B��f�%\��1��. ]O�{Q���-�X������
Vt�I�K�(��Fd�%�gK��υ|^<Iz��0^�v�s�|� ��@���V�tp��N����)5����n���Fl�0Kj�5ӅNB�t����K�71��k��1p͞K�b�X�G��H���!�th�u���/�X΁�6}ap�����_׈�I��\0�O|����*
攮�Φ�bd�r�<��ZK�yWv��"r���숌���c�x��ϩm�R>�`A"��*u�����7�>'�L�I*��[�ռ�(7��S�=���0�XbMB�Ζ�B� ���������|��������d��w�k�>p�M�0���6�w���k�2:5^*��&��\��r?r��(W���L8���L�f7.���&��Q!���g�X�# ��ۣ��$e�r[�B�����%��|��tw��s�^�Ə������+Fי���T(�5N�����"ۻ�x>B�"ܾ�++!$ߍ+��@Q���;��9�YnDX|�4�L����/X�@t��T
�-����@�;��#SI�֌���,%� |�����Pa��r��`�q�������

�L�Br�m皛�ߞ�o�Vv����bg�D7h\�z��J���/�Eɠ��"��i+�.F;iSG�i��ї�ʦtzW���Fg(S��z'Q��΀������x�z��d���F�Y(�նaR��2�3Rlܓ𬌁r畃n�p0�g�к$<c��kk�-�[*-�x��Tk-�����#�ll�S�c�"�>��[�w/�M���+Y	� =��5�ȧUa>��x�㆐����]�Asv��U�Q���6�]%��Z�!Ņ*�e����/\��y�o8̑��h�v�ҹ%T�Z�[G{�J������3��:}���a2�to�K��M��il�x:�?��� ׂ��w�,4Z�*FN
���a+a��3�[��ǎ+rJ���:k�v,uU�ST���q�8h���o��>��hcn�Tۊ���M�#�W��u�:o���Ma9��>��*z��Ƶ�������Z��Bڿ����bl�5�L 4��pu9D�9�mqؒ�V�.��
���l���[I�K�vݕ%a@Ks��X �������܄�b���q��0�����2�2[��ħַ�*'4��#� W�dd��M{6Vx� ���Vp5/���V}OFqc�Y���n����O2����r�wkS��$YMsE#��x_~f���4v����*j��Q	��F3G���|O�m�@9��W����fws��� �����12t��L^C�SFX����b�?JQ�>�f�����WP��S�;΢V۟��.��*�DvE8e,hF���j�G�ׯ`Sx*.�T���N��ZH(��#���K�m�BЌ�8���!A�Î�WM���G��DS�(����@%{���$�|w������F��L��bm��Е)��<	%�2�$�s���+�7�e��w��Ö���7�-ѯ��K	;k>൮��)�E������N:�~�Y�g�~��=i�m�0\١�1��"_�u�yu�d��%;��/$<Q���N�O�#$5�\!�#D/�M5�/��6�{~Xy$acu2�p-f!7Ξ)��$hkʪ��j_����G'�/"=�˻����D�˝/�������d2X7���>�̀�5��+����
|�w �j�� ���f	.l&���z(���=��R��s��~�IeL�
x@��H�W:����آs?�(us�d7��#i�G�/H�J
��� ��m�$V��B)z|7��5:\_?ր�S�A�PQJ�H���b�lJ�L�?=3.�P�j�o��O��f�H���R���8��v��;QڡO�fB�׹ ������}��uka7�=F[��n���z�Puou�����!��3<���?d��AF+nK�H
4�����Ɗ�,��L&CQz7��?��U��O�6f�xPK>�|s�Y]3F�FE>���$����^�	��/h[н�.w�l���s\D�]��������������%���L�nխ�����_]6�Vv'��O�I$1�z@+	wЕ��IK�p:N�M���[�����LU�2�K%�
�sQ�NW�ﶿjlG���1[*z��C�=��`���g����C��q.�<��r�����A�"��l�@�O@9�!^O7�k�<�;��(�)�$�6;*�<`O�c���	0�"�={���x�%�����
� ��/�uF����0E��a�l��a���%��&[�����+�;\�}�]�mB��� )3���c��,��&8U�����-��'�ąs`�ٚ%)��X���7�e�/�=�`�K8�����{ʻ�=9ćcc+���i�B�Yj�T��mڝ϶�z�ܱ���0�Գ��w	&�)��|���M��{����y6����G��>	!op���ņb"ǀfw��l#ڥX;��I�<�������T�aeC((�����@�c�V/�	��,M��5�F��cm6N.)���c��\�A�M4�2�f�J�R�H�:��`gX�؎�oz%|y�<&�3�v���������~֒U��>��`�Eϊ��� "���f�Pz��d��?c����틋���Gh�RX�$Yu�~�� �N�G���,�a@�,��T�k=2�EZ��u���*u�5���7���7p�πH��S�ɧ�X�f��XY�7��q`�ue�>���dX��Rm�B��6}��w��B�_F�e���~R Ͱ�{zdal;tj�IaX-�"6��5psE�V\�,�O���+wB���9�eqČg�DF�������q�\��J��� >YyGB���r�\��T�Y��J��ٚO㲥�"��>�\6-w�
�$=���*�P�Z�%��ӹ�N-����۩��HP�e�٢m_������:9� Y}�:;���b ��"�SL�qX
�0I^B��Gtl�,�=�3�j�A����@=�w�4�Y%wo�̙d祝��D�V'�����?�����{�l\�3���<z��k6[�$���jtQήi��H��ݺL���Py���'U�b�]FY؂|������I�#�Fz��fg8�����+����4�Mɰ��%|��gbA����x)�|9b�z˒7���6}]�!��\��4����F5���/��sڙ�Ծ��9Ki�h�Ǩ�؁t�f�;kE� ���i�Ԛ'�[�v���%`��i(����3`����Q���_]�t�p�wH��1�j�}T��H	ZJ�����@"Q�"���0ip*a���J���k�&�*�� ����F�¨���/�B�0���ӎ�z�&������ ��u���Bf������1
�s4��|��e��Oy*Ij�fD��t�bW�gA��0��y��6�wd���!ծ{[�X+��;y$��(�V�4Dk�N�hw�F'�V���@�T�⊠��L�ț'͆GE3z�:g��6R��_z���y0\�n�58 ?\���,5u=W$m�̕#uP{\��C����4�$1��;˯wNf~���{�ܭ����M�=S&C ���3�jO�5eW��]곐�΂(<r뇞�M̫�EցTKSR^�ٸ�z��h�����%P�~!ɂ�Rl|g#�k��5sJ����=-�OW�D�� �e��Ɓ��N3m�@s��OJʿ5ʓg8L��T�\�;V��o�>��)�zÜ5�D�����X��E)�2�.E�9ΙSmb3Џ}�*0�p��mpz�˴e�U�F���T�V�.��E2�Jz�(����K�6���BD�U�b��n�!�U��hX];]/t(_M+:�^��&R��_W���h����u�՞$b�^4d��.R���eICR� �/)����I�����G^�Hu6p��X���9��+�Ń�J�i"	j�f�l")�.עe�gm��I���" :n4#!�!2~)r��ٕK���#ЏDpV��"ʉ�e�RG��R-+�����^���2��~�ݚ3�%QY���3����]�h��i�!S�g��3Lh
��1wP�3���#&ʔ�BݙC`���xSG٘�-�}8��-{�x4ZVӱ1{������q�`,skԫf�\;<����� O*k~��X��)vD#�r�p��
�.��(�e�&=-~-$s;&���'��%���b�o6!+fWl�����v�V�:���m��˻A�ѭ�Z�Sg*�~{����L$��,��P�]���Z��$�#�т�����D��!n0�W��*?ݧܶ�����b���������z��"�\��[�-��ڳ��<#���ikp��ȝY܇�1����a@Cv|\Ʀf/��^�b�C-��$�^>?�Sg�:B���K���}�3��=(�j��ߟ|�ݐǏ� +m�R������8WuT2�	��"�b,���w��:T���J����pL�C�_� 7d~�v8�wi�s霩1T�WK��X����w>H@U�ŝ *��c+�7��_45�ٝ�-�}�ie�~�O���H����1�-(m����v���׿)��Y����}E��|}�4$����a�r=�]W��ب�ޙY�]�����g6l�~��+��
�,Khf���z�����Z���٧�-y`L/#���PШY.�;R�E�A�Ь*�I$�)
�Mo.R���$��=�QӒX�˿n�Q	��>��̰y���_ԧS���<&�wE^R?������t�������g�M��	�~�/�׋SY.zVC�,�8$�E���*)㐋L)����H�G4k�v/tK���U��r�o�r�v�^��P�J8�H?�,����/"�?��fcE�]�fQ���ip�p��|�q�!+@�?��

cu�37[|�I�xC�2� %�7�@���1�-� X�aT<�y���KZ(5�S)��-�@5ɤ#��~�nR��Q�W�x�T�� o�fWcFr����o!G�u�" r�����V�<LS��)E� ���S�� L��~��E8�Ʒ*�w���1��<�[�3-�ڐ�@�<�T3&-����1fAr���J^�6�-��Y�N&a_�e�H
�pa��n�7;b�<���@��dc�Bw� )�RD�pɘߩ��ؼ]Q1�(�K@^P���F���=���9�á{-��QCK�ܨy�u�r����ek�Rl*�.��;���ox(k����eTL; >��$R��_��U�ƒ�*��'+��*��B�L��I���X�v&ƛ��s�����~j���xD��
F��ԣ�=n��GjY�1��٠��(À��H��r3_�H�&5L:�:���'��b����g)�q�|/�Y>(�������H�n��3�ħ��`U��9�3��S�����B�W��K�Sq0Z�[���8C2\�H/JB�nj91_��Tb~��G9(U��_Tk��J��"Z��\ρSn��v�Ѓ��/4d�T�C�(*a�2�u�B�c�W�x�X=� ������R!I��;;�.$vH�:����Tyj;���L"I=��rZ(-�P曇-�i�c�/�U�t��O���`:�Y.^Rg�f'o��Q�ǌ���f���.S��y� �Z��`K���Ϧ/m��Q�NRV�3�5�Pb�G��HI�iʦ�mH{_.�=G�$�Ÿ=�q#n�*s[M�6��(��|o��u�*T��I�^E"�f/Kb5�T����Ia���hp��>�6qrn�]��胃1�n��H�r���'���?2~U�KGw]w~���b�J��`�ߠʡ�F�"IW��r�"4q5��q�ɥU	[��dWV"��(�R���l��-��4�ב:?q�Q����Q��pL��E�+&���d/89��ʌ��~��-~S�������qv'�����GL����,jӹR/�t@�e.�MP<z�/я��˄�+@�OS��z�k�dz�l|����ک R�m�F�<.{ob��P��Y{	nP��dC�ޖѡ�Nv����d� ��jԦ8�~��@Z,���j�sVh��$�Ҽ��3؉7�%p~$�J��3��J5��_��d�n��B��Q��|3Մ�\�0$=?����O�l���B�E4��{I���,<s%jF��2����p%���Bş@�l@J)/]��#�����V*�B�mHs�y�E⫊/˴��^��h�[ǆ� !��v�{ƺ�+���AP���k׹è�%�ml��E/�
M1�����^ةgV�<zTz�캨'��!���"�����T`Ѻ,�a�3��-����)$���j�P���0��=\����2~�s��汤!AÄf�h�����J^�H�!�$8yO��A�B:K�s��P2��Ǣ{c Ƣf��ҽ��$�lR�ٖ��'�K�0ȡY����4ᅌ6���ѿB<G�l7-|�k��yv�U��8E�1�-� `�/�����F�ֹS�R`y<"��;Ҷ�@ G�"�
]��7��F�Y�z?ڒ���m�WT�)&?�Z�ە�p����zMp�6ݸn�{ə�*�A�p�!%�;�ż��=��x�xk�j:�#���@��b-�H���Lj�
LU��Tk��x5-��{L��t������ɔ[�(wy�w$�-���+r�$\tm�\}����_���e�N#"u_T9�;"�A�EBɽ�m퍑4�=[�m(ލJW-s�}/>��&�K�6��$��r���u�O�ō�h�`F �I�5�<����%-��9Y�:i�)���Ip � ���rB��D��7�v-3|����ړiX��T�|d�wV^i=�Y�����9C�m���D�����2�R�҅ߧ�7����.������.����Z����R�+6��a"š��`��r1�Z�)p+�â��I�L5�����U��r�^��Y3'����c�ĮR�+n͜��[gT�d���Q�Lh�.�2��}���x�1���6�~�$�������ɫ�	����+K�Q6��~��n�:��YK�H��6!GϯH�`$��	<�S5#�Av����5�IO��NIع8�����$�gz��JvUm��f���6: �-�uWe�ۍa\�>���¶�̿�{N�A��=(�!&cbOн� �idJq"�3_�8�sFr~��9FX��j��6��~�Z*�\"4iu�ָ�a��8T�`B�Wώ�j_�c5����\���ye�nla���T�>����RV4&���
H-���.Z`�X��]�d�^�.��V�R���|O��þ8�*e���cQ�����-CAV,�?<����k�#�����k2�l���gX�r}|�(?_�>���I�;��%�h�gHn]
�l-w��Y�6��ɪ�$�䌞����I
���O�l�9մ�֧�b��ts�D��V{2����Mx�"~�qO��5p�}��p?�¡��P!!��3�퓤�Ϛ<�'�YnI<��*x�H�TeV@9�|5��+�
*r�¨)��5Z%�0M��	1S�K�����l[��f�rzz���!!h&�Y
*탂�d � �O�Zb��y�!� &�-�j8����H �������V�ׇA�]�+ܸ��X�N-k�Gr$Ԍkn�@ſX�w�8X�}.�ҙ4��Ē���E�n(*4�1��%Bڹ�����3�D(��'`���0���zI��H�O���w����z7�p� ����)�}���J�\Y����d��O����;��s�x'ԴH{�	n�I��l� ~Z��^K���J���t��HR)�#�5ԙw�8l�g1h�/��Sjlz�-����*�PE���ZoK)[ACN��l�~u�Ѐg��/���q�c0��RԿafN5��$�r�=A��qM�:��Uc�����2�k��x��\"����Ƨɘ�s�97���u���bI\F��&O� ����#��ۢ�:ӾX�^F����;����џ<ѧ����(,\���񿘧�e�f 1w���y����]^	uF�D�$����4:�b����2V�t<�23�w�	����05�n��+02[������|�c��-}�����嚤��vfٺ�h�'T��w�	(ń��]�|cn�������!�p�$��9���ʋ��d-t�D���c�2��I����')�|-\���fy��`@��K�ٜ��+go��ĉ&��ST�lMX+�N݁�++-�L܇K����/l�F���u�eU.��2���w�;�*�FG�Y���PS�\�kTX%I<á��{�4;Yv�^����%Z�%�%HuI�W��r
a��OǊ< ]Q�H�6�����c)��p(�C;
ߊC���6��?��i
�?��~{V�mJA�?M��}Fk�^��+}o��rҀ�t�_�~nݺ������j��f��8p;�#,/DT���Q����F]^+�'I�!$�`4q�K�5Ǔ�����?0�������U;���N�2��UX~7-�B�7�~m���¡�zk�T��/��g`�x�6x�'+ҫp<i'2�n���2䞝V|���K�Ar�;��~�rΎ���^%����I8�7O[Jۚ�0H|�Y&jMK�W�������Iz�p�W�S�u�r�/V��AE�ڨ'�� μ�b�\��r�x}:���F��2PhhGQ澴�.���Y�Q�TL��d]���Rej�W���)g���p�xԋ���ZuXқ�e�פL��]وu�v��ᖀ�Ŕ�?Th�B��d��|�<T�l�P��w;�>`"T��Y3��8��ߵ`Jf�nE�5��D�	�=�d�����(X�˴�߷ӳ�Ɉ%��=�L���OM3i�(ː�	���� �L�������a3�D���9.B��B�j��)�K `�՘��u����ts�V ��9��y��Ƥէ���H���_�"�_Z
�82�%� 6���dK;�0����E>y�pT�s�!�22�j*��X���G�a�ٴ(��C_�5��������ӎ[Y�$L�@�3����J�.� h��.;,fV_��P+�%b����
���/�N�_�τ�X�5eu�Ӑ#v�!�^o�>�3K0=���Ty"����&�<��X�Ə��HZ*��R����!�_,QX��q�!Sh'%�EK�6Fݒ�(a�$�qDu
��}0��'�Q�=�m����Z��F��y��g���T�6��"�-*�z|`-M��k��+x�������	����7�To:���K#�06)x��Ƒ�e��T��iC����j��/曰��|	T1v?�����^pk(ef�O�qL���zO&q�oe	u�v���4�����ϷE� �+�ǒ=�"��򳿽���R\.�0#ȑ*�s��P�I0t��M#�M=�tr������jK���eF.Ҋl��x�@w�,�:��#YG��7G��G��49�;�:^D���c��i�Q9�ɓ�����}����|��,��W�[⃊"h���췄̌�j�-�ϴ�pC@��?)3�c//�Q��'�+<��6A#͢��Բ�*�e�cr�o+��z�S�˳=Ra����\��������>�c�Ue�S~tp7ԯ��W��L�_�������36��.i��P���Ue�5���3��:�BH��H����n�8N�R�[A1D#&pns�u��a���ԇ�,bG��֟����;�K`%�u��f�>����Pq?W�^���%&d
���F��΋~r�hQ ���G�[I�ջĹH� ,�U^�/&����6��:I�{��m�բV���
��7�Q��,�&Ny�|�R'E�c��߰��ε�@���+�`�g��)K:)��"�ݚW�j)nP�&���lu+Fл7"j&�����4W��n^&��qtn0�>�~M.�(��v�z�M�H �W1?^]��S��-vؔi��B�����#�Z�b<����[���о1�~���*\�8��#�T콠/H��^#�`䥒	"��ܸC�8����Pu_P>����Gs��B@��B��Q����5�}�p�ú��5��Ѫ*\T���{��+����Q^�@��|�A��~BQ���곀,c
��ݡ��'�!M9�#�3�Gc�͌��D�ą~���<�CZ��g�ś礒ʚ��s�{|�NP���L(��v������{XȨn���I�c����k��@S��z�1oԱ��_�<CD�C�	W��Z�3U�׮t�\2���ݧ7p��`�j��VX���T��%����G����6�����"�Q"yat]�桊��O��������v$O��"��Z��O!x�����'�
�2��B(0خ�?6{+Jy��X���ݔnY�M@��#�#��$	䪢�&��뤌@Q�����O�a����Y-��&�ګ�+'�Z�C��x�D#
yI���}exį7P*j�g�ϻ��xt�<�~�������[�NNy���6*��UQ�<�A���;uB[�)�Yǹ������Բ���<�O����X2A0g�{k��٤�����4eu��޸�؇�� C7_��p��eF�cGd��UU�G\<0�����
���ʍ%�%'�I�����2�lwݩ�s���Ko���Jh��J?�1��j-d�Av�,9r눑�/.!�+��c�ܱ�� ������o����W�-��q����o^[%Йa��P"�H�.�z/�4�x;3�o�:S˙����
{�Wp��s^\q�tL2�����h��O7�W}a�E(s ��d�+F~;�K�*2Ek�J�Z3+ʐ�`"w��N/�;�6�ʦ�kz^Y����x�"��C���S`	zw��.�ox9���ho��F�4$OL�#�x^�:�::��AD�F�V,p6!�!H e3 73�n]�����҃b�L?~���3��h���۽M�<��5\�n w>�1@��k`�|��)�6�^��z���c��!��'�a~�>��9>e�W�4x
�Q���:�h��v�b� L�����Q���X���s,�-�7�PՎ���J$Z�X"���:C�br����I�S�Ġ��-EK?y�M�O����lrk)������!ơV,1�Ov�
�S�2��Eo�_"�AX2��^���Z�ax�0A�����ϲa���vK����s�QQ��6i�M5<�2]�ӯ�{Y�	� u�+��i�}����e3FPj��l�:`2`[��7ѐ�V��z-VwXg����0|�p!#E	�ݩஂ�K|ׯ����}�g�p�fi�5+q'~-��<���ȑ��`��Fj�qQ'N�F��C0���=h��>�-웏���".���h�~rb<�ן�*����i���Q�yQj�����^�!��M��|����tûT_<W5yؕg b	 �Jk
yA��1u ��?��o	 p�W(?	�h�+��x��#��ob�����O��ԫ�9+Z�W⻙��6O��\��*��͊����	e�r��5]����jSB=�r�	3щrC>ܽ�]�Y�wv�{0P(�4@ �=�8�<w�{cC��6 �@�#:�qp����=,a�}j6�ntpM�]s�f��{8 �;���c�4�$��B7�5��D&�d3jr*L��E���i��7���X�'<���X"�]�_66�NRcuԞ��p[�Y��Q]��q�j-����K_�/m�M/�yGD��#σK�T#��axX���{|o�����3��Y�.G8tk�]9i�lB(��K�VCJ�$v�1���&Ffy�ބb�S�n��a��4��Y��+�JE~�g��Y�[�C%,%k�O��$��?� �0S���~�7�rfp����ֆ ��kʩvЧ2y�3�wJ\Ic�1�j7
R'����9]H7J������"���[V�t�B�EoZ��Z����0�5A�1���K���;%�P�
���l?hp(�g��'/E�9FFY���<�-硢̰�����7�m���
)�R!$05���C+�\�'�'��tf�{�U��0�h41��J94j[��Na��ԥH�fҎ'�V[QSj���^�M�|�Ϊ �����>���H���u
�<c����	�o� ����3]��c�L��xK�������b(�Y*�ŝ�Kx)��;��>��}�����/� �X�)L���3(�w
�����M�ϫ`��Ed�_��Nz�t��[۰���	�?[��RX������ZR����+�|��ya�I�U�����Ă<ʤ���_�4$�V�"}r=&��2ؼ��)g�ys�D���_�=� �,��G$DJ����5^���^3�G��^n�\P�P��7�Ѻ�����M��~�&tn͂�F~^T]�y%Q��C�
g	} ;��\A��"%��:�U! �г������9�v=�S_|����R�Q���ڤ1�)Qp�t�#s3P
D��Ȕt���L�lӮϺ�����t{<A޾"�okZ�XA����󚐢X��1��o\�����u��5�#QfP69m��VaY�g�f�����< �H���*�ԝ�'�P����g9K�pl7��q�%?jN��7y��D�9q����Ԋ�dc}/e$�S��'�
n�����b������&�I�.�Ю��M�+�A�8 �Z��4ms���t7I�X ׾�:`՟�YŘ1%i?�[$��z� n��Qs�� �Hi=���93'��T �w���R?)�xP,�HdC�ߌpO��[7�6��>QK�{P9sRS�aS-F�F�A ��墱�T{H��(�C�&����ږ�.���L���������5ar�s\�<�{���	��ly$#��$MҚs�-ݥ	�4�~�P�Z\�*.�?����i�!�� ��|C
���_�:�zY6o��eQ)L�#��їKV��魁��!4��Jdޏ HI�<�1���N˄�
ʈ��S	@��Eo��p�t�,��<�>鉟��z�=��w.uC�]	-�'�ц�"v��li����N[�4m~L�3!�b����)�9WEn��v�;ޖ��|��	O)N��?�.k��f�XN�(��w�~�:s�MV0x�l�N,�0��G"���l��p1ڲsPܚ>��Y�Ǘ�׉�a�����r����=��y+ъOG^���HV��:��d��:�t��3������l�@��gwo��؀�� �h<E��;F���8]ڭ�q��޷Rg��+���n<�ve�&�!�Q�<��e��0��O���a'h"x��b��Y"@ƦH�R��?%;���M�Hz{:c�`z�&gSs�h�g�g�2�4Ko��{�K��05H��f�;���^��}R��G�� ^9���S�ܕ��=ʷ��`蓟����*ⷙ����Y�-f+;�(`��_a�+=��Yr��B���K"L!�4����n����1��F��@C�~u����H)��rTmP1�	��oTD��L����I��S3�uG퀪��������[�HoK�����n��zRz4�Go��L\�I�(��/ �д%[�nԵ �!���2@3')'u�E '*(��[������ʆݦ��8�s������I��*���L�g�
mɹ>����l@s�5h5e4֠<fzaI�צ����pEˉ��K���nS�b�=9��d2�w�'ݭw,�T�0�����Jo��r/N5��ۏ��Fހ-y�_ѫ�;C��3_HFP�yE_+R�r�!Ta�b�N���ĖS�����#��׃q��B���Z��A����1�;UҒ��OY]Jp�X��_��v�����K��,E㱙�Q����Db�T���c!�Ƹ����I�P��}\�kP�C���I+ Q��ؗ�|+�j�р�e�Ę�4a�7e�EN����g�D��k�5�J�Юc���uT�!ӛ,ݞBC�܇Av�Y/'�]'�����N��I�cG`���e������Rl�pf�Yf��הY2�ʅ�9Fe�v��q=��Ϛ�[<�#eo1?2��9oV)y��q�����Ѓ�V��$d)�Mtf�����1���f~�|R�Ҟn4c��nW6B��p=���_�$
X+������dG�D�$���į�S���cN���U�1�#e���A�A�*z{\ڹ���P�"}�3�x1:�I���2����;�ފ��&��+�j#
��U�������zf6uOe[%������.�oWM+*��Z-�u�bF�ʹr{������0`������e:��A6$� ¾�}�z%�)��Yu�����;$��^W�LQ7���9H�b֥�2��̺K�$Ĕ�(���O�>�)�����'U�Z��ud4wa���Ub9�g&Ǥ53��4B�Fg�0���.��eT�5�{��U@�L�0t}���Q����E��I�5p��P��kOE�ɸ���}hNWi!8��,b&a�
��_A����o+���B0R��,�2_Y9#e ���G}/A]��닩d\?��~�]��fA���q�7�Ib����B6�A?Kt�O#�#����|��V�(w��U3 �Sƅ5M)>J��s%�%��Rx�Y�lY������2d�c��}���2ٮ���l�0G��T��y�2�I��+��r�Zs�,�3�Q}�A�>t�h�=@sr��_�R��8�������Ri��]>@^��qKTTܾ̕
=K�����������.Xn��F��*A%Q�g@1��}�:�/��l��M!}qXb�-S4�Q/���pn]���ұQ�=~lmGww�{��wvqi�� ���6���^e�߮���6�O{�-l�q�5+�@�F<�ӬDIfSWs����٧/��S��{N��W�R��	�PA4��:PРiH7��C>�q�*�����%��n"���5L(}�ع���x*�1�m��cif��O��(����<(�F�nR��-)��	&P[���ˠ95|H���>TM�&�*�%*�J�kLVp?7!�B^6�����c�_v���@؄j��7?7�U>�;Z&�D�nꖥ��$�"���}=L���6�h2H���~�Y����������A�kgj��󓇘��Z�� �>���]��[O�/2u@A8n%�av*�rώo3�b��˞�/d-�X(�F�y@`wZm��T������s���Wp�NV ��[�H��}f=��)��e�5+�6}kw]���9���qwNa�*Z,�YUʱ�e�;�wD�X��/����P�{$�\X���9�kԬ�SM��	��p�$[�ʒ��+�<�Nl^�L)�J��Y�oY�E@�j�P?ּ�x���1�HexMq��(H�3�ϧぴ�7Bʵf�2(�ϑl2�Gsb�%�^3?����G�I�vAܤu���+"�Z}w~�x�� �F�V'����#��@���Ƌ��R��a���򬥄.e�M755��H�屍�;���'L���s�rr��[�i��a���ܖ������W��,7�h����?��^:����87P"��cG�H�S'�|4R�X�KS�l��Z"l����M�I3ڪ����v���</�|u�����,n�H,��E��A�4��o�X</�KW�y�Te��D����9*�jСӶ�JV1�kI	�T�5�0�d��
4�Gz�8o��΂��S[���_K�/CJ��m�r]��ث?CF,f����
_�LB��� �<�x�"3���4�#����?j�ņ�l�j_����X
��v����vB���BRp�wGX�C)(��#X�A0@�����졹 �H���3E��!<B�΢�[�;�)*�#j5D�W�=0;�z�"�3��ea/8�h���@�0�m�~L��?.f��Ľ���L^�D:�I�1?}��RY�yk�Y=ߝg�wV����~H#�{��ynW���`;"b�*��u��;ɅF\��yC�����9Lg��"m%P�du��:��abp���`�7��"HS||�3���qb�P��r��|��O��>����;u���%�qz���IN�~laT_���tl��2��1u��D�wgE7����q��a� �f��W���V��726�k�=\��}��`�X����x�B6��'���ؒ���k���B�J�ʖ���5D�M(�_��i^�RxC�r�e��(8ݖ(d�W�|��s�����H�5$55��5l����ӎ�p�7��)
�3t�(H�m���T�歏Rm�m�>(^m�}�H��4�}F����@3I�$�רvd���u���Ƌ�;!��II���I�����qgh�ق~G=��v7F���<Y�c[:J��H+؝�M�K;�g���.���<m-%�S@��W���nT��Jw1r��~��9�g�$L�D ��0n�0S�ReU΍�e�J��=g"'��{U~}�eN�� ��Ї/���uG؁W�! }�#qW��c{ذ^���[0a��	{U�l�RaZ���)������W�>BJ �~E ��Q�.7ST�M
5�@��AV��
�U�!OR�%�'����ﵣO���8�s#+�<V����M@7�?^�ͨ��`�ײ����U��R��H��O��6��)!
ȺX@�0�7�]�?Q�����X(e�g�P�(����nU��(���tL�l�m�?~ץt�̦[Tm˪�.�YP�Z�6�
=Az�s�b%�{D�dR�@LO�'���$;���g�9��}�ݞ+G����퐿]��S�~��{f���!��]�k[�B�%6��7%�E���#c��0�ՠc�)8���36��h���܇��9t�tc���~�51 sP��Z~��f��#�Txn�"jֹ�"��P����A��TO<CIU��G�f"���L�E�.�/��>��822ߪ�Ű�C�����O�щ�5n6T��zV{���(j�E'ǏY��0��\<�BS]!v�&$NU��3�k���jJP0'|�k�I�q�v��&>] w��n���Ő+���"p
�>���,��F�|�عd2�B��D�>sp?x�����Y�n���9�V?x�Niʈ?�i��2N�E9�Y=�|�?+W�>�����G�v�[��;Pw|;�������Ei��#�[b�K��х���F�G��{��ГS|c@�$�ꦏ���L��{�a���7�)wҧs-�$J�@ ����J�Zj��H^��_s���x���v��R�J�c�j�J
�&z�^ˎ&cL��`��H�j�0oU*X�%�)��q�\�����s�,J�����B��Y���7'cyuA_?���I�Y��x�$��NH0x�X*��|IdhA=��1RN^�B	O�3A�)GD�e�:O��$�v���;C�Zꄣk��|qGÕ��PWk`
��V#8�CW?��GL��$��i�h��<(.<������)�A�,��!{��#�C���0?�Λ�k��Kv7�,�xR�8�_�$W61��6Di2���q�����,�+&�Z���cP��+{~����a_�u��ډmج�{\~��i�J�/�x kpa�I�nW�F͞#���C<r1��V���v�3��}���{��P�����	���o1cp� ���-�ԟ�����������.V_��o���4L2|��.מ��߼M���c#�_�����c�R&P9��/�캠�0&h ��g܊V�>\Z���n�>�	��n���mխ�ݏ����m4�bo�1�<��8BV"�VT(4�O��o�vˏ(|H?5�p�t�����C��XZ|��6IDp���r�GR�\Uo4QkP���hyR�����v��=�93~��� ���;� <?��{�N��&�;h2W��p�ی���{]�R�}L��񎋋�g?a�������m��^E-��N�uҍȼE�����D�)�]w�?��x��H��ɖ悥��UG:A�60��wb�`�*vbqBT�g�Q;*�>�cz\Vr����J�sas�v��p��Eގ�"T�����dF�?�#��y���;�I'�wc����F��v���.�y�t�4����c�bl�?�@�h�}�������*��L��
y���{��7H�������n'���� /�îwe����q�D�[��	�i��=G.�u��W@Z��V$e�Ϸ�"HbH���Qrq������<��٪��"4F�%�Z �O��<�h'�1�u�g(!�B4��~��U�3t4���r��U��+T��!CjpxF��n~����Wtc�=2c��.�ܣ��D%�1��Xe�=)�BﱫG2G�{ĩh'�����fp���86Q-ƺ�$����&X�&�Ѯ���oA����j���p�=X ��*QJ�K��/b�}%i�7U��,��}B�F���nkLd`�D�/�ڠ|����R߷,R�ھ�/���K0W����@��kc[���;�Qs
ϜO���9 �S�ÎR}���/��G���_r����3˕����~ܤ��r}�;3�f� s6-����5���E�[vZ��#��3����	��D�
���_�%+��t�u[�Ѱ�Oe8�vk��<E�E9�Q��_`ilȘk�N��|����15�q+�_�;AD��*����G�:�����:=����0 �H
P�^7�%��Խ�쟈V����j���B��;V�-��Y�Z0P�������%
ߞ�
[�9d�+9]�\x��J1�z�zMF4�.k�Aa?�+��48��1�3�~þ;�w@����~1�˪��8y�ĵ��g�q .4��5����Hc}zG����'�rٞ}&�seb���H�֌䧋ځ�{���y^�,�z,�u�@�ܺ��x\�#�d��Yj�g+B*`���4�m	G�`��^�Yo�A*ǸHر���-(4��g�B���a�)���hȏ	�6a����d��IJO���=�4k�#%Z�7��T0_�|�g�"�ٶf�ݯﮫ����k��N^�{\��*��y�k�ij΍�c��6�{$����vI�Qsx1�LT-�
`�x�yo�	��O�&��;EQH�	f�OaVH����!��覶�Ld7(����+4Ho�*�s�Qp3@�fkR�"����k�߮a��%U����a	!-����$ə����E�pu���C��gO�;-��`DS��~��������6c�Fo�*!m�o�B��c�՝�B��b2C��;g���C�M�_I�.�]Do���+�i2���4��7�"�����Ƕ�@fӶ�Al�aL�V�=Tdپ�{�e����`�r�x]�Lg��q(�Z[&rOf���޼D�]l4�?�9)�#a���L
{���5�ۂ0m~��A]A=��Q��V�ǌEu�Y��j�>� �A��"�ŝ�[��^҂^�P)�&p"�s0C��6���,�n�Z���&����`�=Zץ7u�� _K�h�w�٢�ܵ�5Op����3r�1����-<�]@m�����`�hüՈ��\���[��Εk��g��yA�#�Axi�ne���aI���%������"���BZ�'�7��_������4sp�!�P�f<M�C:�͞��)�P���w"l�m�%3"7g���p�JC'�����v\���-H��F9!S(f0V\ EY4�gc��v�g����w��m'Sݒ{���+7$�
Fq�����â���G[SJ��T7쨰�#H�����e:�X^�źϮ?��ڻ����Wɽ��2����F-��M��K���П�5Ҥ�������t[.n[�Dd^�>@W��d��sQ�����~i�4�R�z��"iR2��E�UT��`b�Mڙo\�J�a�3Z��|K�P����h��P�u�R�t�����kxFh�7�d��6�Yw�Q�Ĥ7�A��sm�u�(��#S؏��
	��z��nz]-] ��Y��`#0����O~���8�o�QDʒ�/�=BJ 1:��<]so����G�u��r�Hh/l|��R����]���u+��������8�S��eP������<��Y�x�P�_�ˌ׺lP>XQ�={�� �d*q�]�b<��#����s��6*;|RDi��|�:�;�G���О>�������-��5�_�'K/^jƃ⻅ط��^�n0S�0>��.�4��
� �/,��3(�;萪��V�d��3�+��Q6',��9n)~m��6�W���{�7������l<��U��@=b����R'��׏��1��쪝W�k�ca��q0G�$$F��q����!�JО���M,�fT��	�Mz3/���B�p�T@\��15���3f�i^o��Q�k��)ɯ ����Kr��[r�˄�=qHCFJ�I���"���Z�j�_y����VcN悪:q� ����`�'�N�����>#����'iE�5�Rj8�:�|�|��O�8~����i}�B)��K[2<�Ť3yd8�eW�ZOnQ9�����j��<�v��i֬3蠗����Ri�H�23��3ݧPF�^ޘ�s�b�D7�Y�,c5á�`��P\�!�>��OB�����RowL-��$S��S�f_���8f3X�2�5^�St�J�7#�H""�ftV�I��}b$q�h�W�B�:v�Ѫ�,�Os�g�C���}�M��J��x��I�M%��a>b�I����΃	�=��+&�N�%���m�Ĺ��ɺSL���`-GiE.I��T�I2�kK,��%9+,ݯai��V�F.�jf����G�/�/$�5#����l��� n#x��g><��u�U�2�/�oL�$�(ݕ��`h\Z��6�jF��g�~�/b�J+���H�:$U&��)�؝G�\nk�z_�����{|I ��Wdn�$L���ȧ*���h)ŵ�p��p��m�����d����:5����m�����������Z"u#,t��<uӪg�Gq?�@z�/)� �
űF�̩lr&j����n��>CO�_^\�E\*��������4�����2}�DX]><����i.甸kGMb�r�RH�N}�}�n4�k|�$8���S���d�z�^ؒY6��C#~��&�\p8�����Ŋ�N���?�ف� �٨h�ՙ;dt@�����I���1�pЃ�CqЩȈ�����em��h}�0{�fr�4���ݷ�8H��y��#�
2�z+{���!�U���4���Rt�z"�����ٱF6k:�5��.wk<����-�>'�;/���� �>I1�Bޤ���E-08(�	�������b�VEY��{H���<x�\�h�V��E�J�И��a�w�
��d����Q���6�}|��Lh�O��:gt9���Q4�t�y��"~��9��6.��|�4'���	��K!:8��t������7-��A��PI�_�T��Ć�P��}U����e$	�dNn�"�c.&.� =>�o�i�=Qc�:]y2ނ��˧���gi �
�ND]���-�\.�2r�;~t[h��HPA�4�ᾁP�5�[�D�!�=[|�C�	
-���[X��WYx����wd��	���B���|e�rl�ց�r�9�t^��i&Y=7��~_����w�O�8��FL�����`;��?kk;TųӞ�X���~�7��u��#�WT_tR>�~�c�:RÁ[�yg&���e'�{&��]�e�h"jN���ϴ�Ni�$s;��ot5�,\˴���8��홠�/���W��!��Sbn���V�?�D�H���{�]^�ߡ�0>�7��}x�}V�F�3b��L��©�M���1@��֛�/���A����zIuA{�s�=����,�X��FpZz͈Z�!�\�i�v�w��B����m�򓐙j��eV�U:��/ ��(��6l�L^��׌��J�"�Qo���(���-�,c����Px[ Q�C���2�:�?!;:FBO��+�b���$�3'EJ1I����
��yi����V���z�c�:O��W�Ha��L�}>Ki�s���;f�q�?���+����d�j*�i/�˹����"V+;Ðb�]���%d�eP����a��V�	���Jy��hޢ��X�&QQX_L��[M;� ����` p�3J�n�=����äqlq}�H���B�6�&�r�������OcڴX�R�r|�N��3��^yd~����K��3��\!����l
�p����5��<��+�c"}}x�y�t�ey�3�Y�(�Rr�l�*_L��>d�N��mACۘ~ݸCb�~ҮI�L`��6@�tkD���Znpꮼ`Ѕ�k�3�1X�4wD+[��/Cߋ݃ߋ�J���n�a
�4���A�#]�@�Gn��$����J��N�iV��!�N��6r��k��J^�n�m�E�e(.޴0��b����ؙ|�Ἆ���9�G	ժEC��~!��*jv�#���\��Zn�C-d9�~�N)[�
x׋�`������U O�J�Om�O�Ǭđ���*ԭ�sD�Յ�k���rD�a��`�O`7�֏��q��z¬��sc�4�E���t�A\r��N�G��)6�%d���h,Y�5/W�AԊ�OV�ؑS�;o܌���q+H����[G��|p8�RN��/�y�%C$��I�-�f�-���P�[�{,3�8����֕ć�N<Y�q}%���ި��$x>f��.����Bʢ�
��X�WV���P$	�R�_���Gz�X���� �a�^�50x(P�-Wڈ3��<*���սV�Q�{��؇2>F)0N�Y)<6;�Ӈ���,K�ze\5s��~A$r4���ɰϹ�Hp�FF�⵰x�?%�2�Y`�iF�m�(��+$4 lo�=�>Yu�H8[Zk_��J:���Z�� }%��b����×����L� lSWM-H�>�E���dݖ�1�i㼙!�ը6��������FO��'y����M␬a����nWm���"��Ɗ���xUCY,���^����w�
2+&p���ފ 73��'r�)�|��Q�è̶������"�12"�ƅ�*!$RsF�X6{�\��u�0����*���.|C��z�C�J�F�q����C�9���h˾<R� Ÿ�O�c�����$U�����&�j���~@jdUU���>�3#���ic�/'r8&ۡ�X�}UGS�-l���RA�cn����Y�N7�d�W��k�,���l�js~�Ú�hYK&��ّk���~?6��h��"<����V#��?J�M��#�H�5K��]Xo2���&����VM82�`�:�?�2��ι����d�4�Ÿ��;��h��#|q5�+�8U�ۄ�;�SL�V���>�vii(��w�ן�4(ʧ���9?�'/!�X�^�8�RU~��ZE:�����;�'��<�%�_f�?x���S��0��Z~ 5�LG-5�'��]��ު�m�`�,j��nW�������eiӏC7������n��&)pUZ���|�@�C^Ǆ��R۴B#�X���qV��]&�#�%�m��%9�@��۠V�'Q����������Z���_}>6P�q'��)Gz1��	�����yx������A�q?3�=�0R�>����2��Gݳ~����o��Z}��;0 ���[tH��}�a�8������cǮ ;~:���Jt\W�1:�{
I\ �QƱ7�~SX�^�F���k��՟P�sOt���{e��H�`W���8� Bd�.coc��s�z��ǃ6�@^L�7$�5���-�h��JP�/��r�a��c\����>0�d�����
.���Zs���>W@aI��Q_����X%��#S��Q={⑫�o�視*��A��lB�G���4�Ýc��L�+���͹鿁����}�,W��Nb����w�xi��Lh���8��!ϳ�iNզ��Z�eN��t,j���J���L����(���@1��C��w���m���3�yG{��{�U E�_3�D��iW�G׳P=鉺.A��x0����'3"E)N$I�}nc�<���Iųh��&���f��oӡ%�Wȭ1�bjrǖGW��09���2$�i��s!c��S�0��,Y;�A_�¥�Q�՞�f�!#!:R1 �j|�=d�f����3 W�r�"��ϒ0�H�Y�nt�Jk$m���T�L)>��X�}$V��=��Q�����3+��䷘^���`�<���.f.N�,�U�p����14���ԥ>yDΝ>��+��%�5�kL�0ON�Y3:��!D�LT�M�rX7��j���4#����N���\�9bӈ� ��,���,B�?��4�U�;(��[�l��4đ��TaL�k~����B�#R�I�l�4�x���R����\�o<1zA���|�C���.�OG�5Bc�K-o����'��Vt7�~fXP�#� ��y��e[���3��uT#�"���3��gQ|7g�,n�r���.������d����'�b�32=�.y]��}��{?��f�W�D����콶ڍf��Q�IP@jz�X�B�M=d��\�01m��L��d˱7Ph����i\x��#����K�R�
�t�XSWSRs�7ل�`����U2I(/���3�eP}R�v�rN�سO��񽌠@J�#�Z!Ę�3�c�uZ��9�.u�yt�X�!ǅ�n������N(���P܈�6p�]4�u8L�zA|�xs�S�|f|bûЍ��xo�U�0���X��ٜ騝���o�S�Å˵�2��Y.�-w�㗿� �}2���'?������r�߫���hV���_��R��JC@Cy�Hj������q:�����fz�|Äx�����陿��!ӣ��b���Y�b[���n7�.�x���'�,���R�v���`�	O�"h	tA
���؆IM
�'S9��qHҬ���+�rx7F�d��Ӯ�Y*�T"$�1)��q#���-�e�(��2�ğ���	wޖh��! 0J��b�Q��)���J�.,��&��9��W�B��$�����+��O �\��9zU؅<�Ǘjܦ�A%��n-Ё���v�:��(���_�p9�֔˱*�94��2�b"�T&w!���(}~���҆�#p�g����B.�N�.�k�!���D�T�����9ZG/�8r%��3qh3xL��#���%���$�Z�2�C��Ӄܩ�qQ��mdk������ �B���kU��q%)g#;j�ߩuGn��Xh����i>�9H�'9,U<{,����'	��VS��,{�i�y��_/�i��m�C }���%ǵ��~�
�݆�l����i^�ܱ	`���!���T����#�dWQ���5��}�B;�<ʮ(�1v�K&���tD�9����2Z�1�0�Mg�ʵ���2��:�;zk�i�+\��3J�P��}�h)Z��VVO������q��FC^�����_.�*�j�V�ír&��g�����'!N��V)ʽQ��b^�u�l=������}jr"]q~a�T���������[>z&����{
�;�ں<t�b]�s��漛�K���, ���w$�&ࡁ;)��gd��DjG��#9`r쿇a�5q8�lJ�	�w4�1I!zl�쌻��Z"N�xe;��NT�m���D���;�(=�7*ܚ�`�ٕkHt�o8Uc]G皻N�b��й9���,Ԃ�����}��&*�f0:a�.n*���Xs�6�XJ�U!�B��げy� A��v�	{�$5���$���v�8�k�_c^�c�G�:D]�uNJ}N�,3ݬ �) �������;<{�ǝ��>�_��9�aƏ�t2�I�iPL�8b��ރEc 2�2�\Pn�jauxOy��9��d]���	m.-���~��|?b���d\��$6Y%���*�?;JVԳֆ|�����hv�P:�^��[j�	�n�n�4�`,"���/�n��Ts�!K���i�]��OP<hXi[�qel'�;��s ���#_(�����5���OZ,�dǵ�[C�u5|IgAw�,�\�*u�tU�MPƄY,�c
p���^�mxT-����u
|y}���{a�UR����U����Ȉ'�]�#l�+t�}��[�lA���,��h~;�~#��r��	h{Z���$hV�'��FĚIFB�SN]g�?���,�e/��c̄j�{��� V3��s�+�ڪ�Gމ���I�BE�g��9�0u7���Ć�\��4�퇒�PL��5׃����p�#�HΒ����!����Q�[y>��Շ&�D��bq�{��EV�v^��y���U�d�>��CKxb�I��L5N$\��t5��;o������lg@/�T��'����XT/f��U�����g}}�rLG�х�Ŵ��� v��5��/Um״��1�!J�F)�r�ty��c���mX{X�z 
Oz�A��$������XP]}~O>ϐ
#����9Y9w��+�-�MdTƑ����۲�-�}�:�-:��Lc�L9�Q���܆&�1�GJ��Y��q������t6ed6��η�/Μ�t�|��~�8>I��2 X�P8k��Y7*�Ĭ熪����^�"S��U���c$�`�2�z���T��Ot�Ƹ�����-7UԒ�m��o�`�: ��Up� @ۻ�>C~�x�)�~��j�Vc�:J�:�7xAU�O{
w�޸�|O�]�cQ���Ҩ��}��KQ
f�-�3M�hC����m-W�q��}f�[�t��~R��*�ɷ7�7��'�;Q�����!l��uŕO�l�؃���EA�DZ����[��_�)�)j������o���R�����ʿ�Rf�#�;R�WO��Γ�0D���%��H+f$��ux��$�.�Jj(V³��(���Ax���P�
84�R8�N�/�1[��Kyj�X}�ȟA���Ө���Z�$<,C���?��Nz����=����[)��������L]�����OäA��
�J��y�Fa�:G�i���CT2�v��2{��n��`�Mί�sf*pcBr�����(��l��� O��{[>�{fv��4��J��������!���K����X�D�8w����$!5�w����$��M�m���t��� A�WlA��ͯ�M����

�+�vϕtrg~�X�p�&��B�Lj�f�ԽH��t��~�3���UMSK�������-�����V��P��e`��0X�@S맰�-�Oh�l@�MV?�!'Ynm!��Rt��PD�&]`흎[��C�Wd�˿jɜ�d]t6�2����9��('�l��q��ro}�g=��g�؅�� ��̻�ӛ�z��`�]t�Q���)�$w�,gw�t�a���6��J�D�!9�͕Vۖ�% �U�G���e�!�e50�^៝�4�i�ZĴ°�$�Kx�XC�uv��H ���a�YUW���h��ɘz �+�d{��vEob5���Sz�S?pzd�.r����֌l�[���	���P݇���j��#��Jjjk��P�0�ű��-'�蟥�]|y�( �s9jM�]�w�hL�Z��5L�5�C��%�ıUDA�[�͔��-�h|��ը18�0�W�}��<QP���,Z�����N����Z�g��$wU��R)�p�Zǆ"6�pֻ�9�d2�b�u�7лv0,����pީ�S�������v��1A,c�)�#D^ŖɲSl�^ӂhFUUMRkt��F{Ee�ǹ"|��0�,��jjN�>:9�9$N��Pj
���gjt./�"l�{�5����J��
�M���}%1{�3ڙ�p�nZ�	WH�]��l��˗��GTm�kƤl�O�@�֬oxD��p�JCc�%��+��B�:]�#���8
ue�JP�/ֈ��Ԫ�^ü��S��h�(]{J$p�`���Mx������`y�t���5t���UA��U�+�S��jp����7H����	&v��R��ɣL>_�C��h�>I~5V��˘����"HB�&$��K=�~�Qۆ ��N�[e�cnH����n�0��_}���@� ��a$ò��F�����VD x%�x�4"MM��(�F�]}i�J��6�h	�]qn������]>��a�|��o���%#2������~��B* 	�P�>�v_�]�����޶����������U�gA�>�}(����K��Y��p��fT,��մ.[O��q��zw�͍���&4̡��kP$�Ȳg4�*7�Y	�E�WWhD }��xI3�3�5<�m���G.%���?�������u3ջ�s��12�H7����^�Gxe����!BxYWl�D	�����ӂR�՟Z����ˑg��.��x@����C�.f������N��-D��Uܚ#J�����&'��ũ��rQ;�������++��R�"+���п":2������ņ������k�}�"8L����;92�`���w��R: d��e����Y���	�o�lJ��`�,�m�kN�� �^�B����ڎ���*��ӽ�|����E
�_,Q�N� \oѭA��l�}ᴼpC�Hb��'o����oF�X9f�"S9���ؒPjd�e�][�jڛ����<�x�f�&����>�����j���vV'��Z����A��7��e�R%^k��2(۱I�Pz��V{�4��B��u������̝[V�H$&P�ggQ�PC�w��|��̕�/@�;��7ݦμZ�H�<a�^�aN�+���rǌm�R0�b�k
?��� cS��)����/�d� {�+Z�s82�	����n(�]ψSD�ҥn�C=��ӾDv�'7�D��\��]L�*�X�~z#�
J��r`��Aw��m|CdC�Gm���o�n�o:z�
]��gI�j^]h�Aܭ����R�e</ϫ�����]��^�~�M4d��6E�)ˑ'�@8b�!���Y��� Cج��;3�R]f��jh#�2
穗`��2���>Q������ވ_j�\�����c��z/�y�ܰ��6�2�̘���l㘏{�+B�����|�FX�9��o��݁�
�ƾާ��i�eƾo�Ɔ�z�걖Px��ug�0�t�^h�v�~��n�@�ߟP*S*<�%Q�t��6r�	i�PG���e��R���*x�����+e�ͺ��y�u�#3�8a�Z�%��GFj��֬�X�*u�6\��.���?����OX���}�1^��`�L�Y�y5��@���K2:*�=�ݪ�}	|�W�TPQO,.�0z�!s��N���쎜V�X���R�7��r1�te��3��4H�hڏ��4�9�oA6O�߆b3r���8c1�R�#�(t����ē^Mi�FZ/��Y��Y�S���µ�V�Z>�7C�,�ˌS}����昅=,���I�D
�s�6n1�w��Å�L� `*H�C% �Q��ݫ*'קy�q���Vh��M�tf�QA��y!��KH�z��)	�`	/��;$���Ą�m��}�ď��*l�~��U��@�D'�O	�Iᘏe��&�X�i���;���w�0�?>�s #�b��pƴ%Gߧۻ�ot���\��c��[��?�pj�?�/J-fYd+��C���9V�b�@�ټ��?�� �nU�7N9�ICw��G5��8����R�X�\�� �7H�m���<!rAOhu��^x�j����S>�g��[���W��ϡ�ێ��0��yg r
k���:m�'�uX�Uh%�B,�`}�DEn��]Z�&����/�;�?	��mN��Q�j�b��1 !��g*�U�w mpX(�~'�1�%����I��vi�
a=��d��g���&gj����2�7eE9�m ��u`��<�v�{$�{/8?vu~lϱ�=�g0���=���w�B�d�Â���-�I��}t{���J;��\�@24t�	�1z#��J���n�ㄕz�J
,��RmӾ9�/�r�����2U��ɍ$�������S��-�
��jЋ��e�]�BO���t�j&-kpă�����֋���"HQbgE�������`5��7G�O�,�#�0p(W2YY��ǃi��T� g�Gj؏7 B�~6�1h~0Ș�W(xR2��1O��nY�����n�� jT>����S'�Ȃ�¸��QDV0]�	��rb�ML\�f�c f�6�BS�W&3���<ĕ��Ϻe����Y��o!�U,tG
e�S��/�%YYR��\ ���ؾ�Y��tbj���[6t8ᔇ�=�0�d�k����6�A����gγYo���|P"��q�]�[�!�Ԇ��\l�g'�O��e*�V��q��z)���P̌�T���j��I�p�5	
���
�J��^���`S��$Rt�m��h')a����N�CM�r���F6-��yŃr��T�.��w���ܚ"jV�nP8�?&�}�0�m��u��r+��R�<d#���=��Pɍq4:+���w��0�+x�R+�Dj��a����b��U���lN���3�O,@k�s����J��-b\b�KR�Z���Q�;~0�r������N�������i�u��>��Sak[��"��ٌQ���r+���g��G�p�`I���0�P��2mw�N�/�9=���9�F�	=����9f?��Y�A�a+������^8���6L��:2h������n��LN���c���t}M��L �j�h�N�i�B�����cZ�aK<88��ׅ�=�$���I�u��r氎��J��ĩ��
�S�_|�����0e��N�6ٿh02/�a�#�3�yd�=��i�!O�(=���}�s�x��Q����J>��vf�Bb���P���A�j�}	)n�JЩ���x_�ϣ�Ιc�D��KL:�ẃM����M|Ek�\���H��ܭ]O�	�q���%����l)uQ�Ȅ9T�����"%,CH2Kv����,o��T\��
9�P����|k��f�a@��Ga�F]��/>�rE�Z��K�_ ����*��#A�(bO] �6��6��M"���?z�u-S��H�at����(���R�����\�W %�`�!J��P�`�K�f繟:��#�HUër�p�
��<?a�r]��ി>_v�����z0ѩc-ô���C�璛���Ft���x��v� �PM4\pl�,%��:�c�L�<�)� �!O��l����#s6��I>!�fiA�P�z͌����C�W�]`a��Ũ;��:�c\n��E�!�1K�H����{yvw�}ظR@�ݱq���E�jj	5��N- ��m�q;NP,l���^e5��&=��h-
?ZB�b�P��cFG(���������ɢ�$D���Mƽ.�9�U��K�-�ٳ/�����LЋ�}n��&|3b�RM�$���������l`�.���N��P��*3}8� 5.��j�?\)tBdVϼ�bN�X��!���e4�Y6(Yۏ��6���4��34�S4�_n��͠��cy���6�����c�2�)�=e}��.�
z���b��V�^����Bk�?4fE�����Ő7�E��A£߄����O5x��J�k�ŵ8X��'C��]��Tɱ!�8. $Xk��aoD���ܾ=V�@��7]�t��R8�ۦd���K[y6�������uha5-��ް �B�B��~=��'��}81KŉSf����C���z.@�'�s�o�J�˰�!H�dڭ7���t���*�x�T�D�-��_���#��%�����X�j�ۊ��`�CN'qx��X0�Ps�n��J��E��o�Kif�i��$�g���(`h_�D��PR�]�c�f�'nx����-j��i>87�l�B�ܪ��v�����q�C�t�v�<����F��'b�9�채%��,��3�~����i�}SӌwH��4�Pɝ�m�L��碪;|d��-Aoe=��N�S��$���Ê����S�������f��:����_=�1�kA��	�<MH�����m�����<UŔcD���:�	
ú#UL��&���U~���V�|P�ܗ����;ƺc=!�yL�������vk,@��5\\N��vM��΢~qR����Js�c8ʱC���u��/9�w l��s��P��a��X��+�9?R	���?8�/ U�JLD*�.��i��M}��#e��Oڑ������U�59���K^8���̯�j�0�������P�i����^ӻ�z/F������L�'���������3S�#��M��#W9Ʈ+�t1��7H���jo��@�(	ǡO��s���Z�G����|�7�8x��p���v<B�������8���/!�����#ɣ�M=�|���L���
�`;��ס�F�(��=�v{X��h�Ś�zQ�m�hx�oR,_���e��ot-��:�ً�n[��M�>����3#���B�L9��p��H�a��3�V��1�37���r'սO��T��x�V��$�qOaF5��.r�V�a�+`�����x�-e�V3�Zv�o޹������0��~��������(�!B�
{4:��	����Tт�3-R��G������Cxә��·�(x]bF*� ����*@��\�dU�$�?�v���ޠ~��5�c��T�8�(ڃ��Gxw�r�;}��F�_�|��L����O"�3�4@�]D�<s�t��{9����@}�7^/�¥p ���}� +�ŤrR���O��H7 �*�|��L��h�� ���f��d������0���pnC9����z�Ob�zZ�� :fZ櫵�u�b�3�+�#���ٱVg�	'$�d����u̠k�ӊ|�I�Va��*�7L��#��_�ކ���b/����@���#%`�;��񲗂��v�^\-��h@~����r��q�'��Q�rq��}�uu��c�ߡ�/�S�<٠�N���K�u8����H�Z#�������,��S� ǧ7�[$#ټ�ҽ촜��!.�ӫ��&+�~���*��te�� �'D8ded�iڻg]���u�:��ǉ�k�7�>�}��
[�RX{t�W�A{�,�i�_�*f�`���⥟��g,�&��/�<�W��Y��$ٿ�G��Q!�ʗ�J�̑i�&�/�qM=���v����ؑx W����bz�؞�O�t9$�2�\�·�|M8��>߰�r�K
&j�t�|ʙT ���j�����d�,� �R���4o��I���)���4�����#< ��3�H�Q�8��be/ΊO�J��=���x9:�ٳ�0���i��q�6H� ���k��ú��q�)9�n��s�">�B�W`��GS�&�S����%����/	��?]+�����_8� LJ��3؅)�tۣ]x��N*�Ѡh������3܋�xK�8�?�E��<s5zE�+L��UF����\1�5�|V���ۯ��+�k٪$��2��&���Ǯ2�K�X	�6t��LE��Q��e�?<��?�WF<q�g�@e�W?�T�0�vh��⷏�����i���]�0ed/�6}z@ �Y��G}�9���@��P|�g�>aZ�=�@R�rr4��#T�x�S�Z�v����X���?��6��*f�@g��O��7�AY*�^�q�D}��C�e���~�(|��9�h:�ó�iٜ1����$�	�7
_!�������¡Ol�+o�038w�W��Y&�S�M�� 8���ن%��_�{�;|���� �ܔR�ح$�����F+|�͂5�"�%5�g.�TN���[��� ��j��i"鮍�6%����l�.�y{+�~�2ʪ�<A�Z�kx�'�@*'�1�2� iX�����w��U�$��;Ѷp{R q N���Y=h��@rO�������:�����kv~l�zU�3�A_9�^ranzGz��9��Zũj�0@���0�H����<�� �&��3te���R.�YΉQ7�߃dY��L�� ��� :�RI/�>ĪE^�[�m���|eU}'P��4�/�F#&m��d<jnK��˳��Y�g�>[>8$$u ��Uf���)���o�O�U���"��h=�!`�rru_Iy\}+p^�;SN���� ���V�Ɋb[䌢0}DD��ެI3d��ln���d!�/��`\C�3�����a���&ڦ2r�b>�a��k��a�6-;S�.��O�[N����ĕ��Pg�>��T7����B��Y���l7������2��^�*����ғ���]���'��#��F�A�g�"H�"�W���\��mrJBG C�����o��Dt��;��r�7���/B��~�ت�J���n�\�l������U��}���<��pA���P�+�i��=햷�vR�0q_�B'�\T�,�!R��A��#u�=^�8�n���:ə� �"a��s�������G��n�&	���.����Wz�=��T�cs���<4�T K�a��cz���s��'L�����e71.tCs#K��$��j U�F���#u����z�kr�{/?&8�?�:��6/
l����4={&�bCW�B�}���O�I4���0"�]T/3�
W��V|�k����(�i�T��k��j>LB��ew��h�{3<0�F�䰃�ϕ ��07��W���,S��PY@W9�4Kͫ/Se�ɝ���٢�zLus!x}B(sG�~$^N�����OfՊ%B���9�ut=��F��������F���;
�׃�˙����sz���=!�B��h�6�HQq��ʉ�̬i�-�`���8�|+��v������*�ք拉eZ����^H�9���n����9��W��2��a�� �_�GX�[�|r�}N�_���j�/ʠw&��%'㋅�Fy���������?����,1h�y��iɋ`RT�a���&GR�a��ھlzk="�E�{{�U��y����[��0Zr���܅G�h���b붗���e����z|&$�P�l��(�ܪB����N\���Xy|w������@�'��HvUIU�T���rPt՜e'�j��B���w��9��sI���ud�e$��N���jXC�\�-bC��Ӻ���TN���[~{4F��rw:d�w�^�^,)4�Fx�U����$l��AY/������"���U����(-1��,���L��/��x�@\��~%�I|���xB�mM�
3E''[u5�1^:8P!�d'i�3����D�R8��V�
�%0EMߠ�"t!��Os� G M#fɡV�	�r0.���Bu�dh[�T&��3�X�y�Od�4�?hk�h�V�O��?������Wx�1+G�R��� ��}W��qH�����g��օtCL�$Y�x�ZG��\�骭X��V��Gfֲ��\s?�6ਿ�vp
h��p1H!��ճ�G��R�	DSYkFp�9�S?��7���*c��H��b�
�*6��"�#�rg��&?��o���h�BTB�8�T�T�"��Z�jU��Q��ƅ������!5�j���
i��*ZO0�}���ǀ�8�ݵ��!����Ⴋ�.�-�������nZ�N-��Z���؀���A�KlJ�M��W�ƀ�ذ6��,/�[�ðR:PݩQM@�"��3���X�مuN�E�>*��a�^�Ss���p/|�T��0�Z��80m�$-p8D��Y�_��?��y�-<F�?ւs�R{�w\� �N_��A�H-F|�v!D�au~�c��Ή��r�}cx?C1%�-A����6s4�o�S�R�u�N��K�u��+��a?j�n4�����Ϣ�N�7%�f˧���JW��dGS��2Ap
8f $� %���8����}���&�x�
\��H�GA�u��&bU���)�[ý?�Z(W�:�m��`�Ljt��'m?v~��	7 �d���s��*9${s-�+�8��m�U9
��*
L�\7����G��Z��6�Bx�D�񵁦.|���S�T\�t�i0��=ӵ�Z���h����v{��UȔ(ZX���P�Ij���pRjw��P�~�l*6wq� %��kk��ǂ��c"u��TpDD7�c�w�t��õ��۩���@xm� f}�dۤe�Bh�3U"��*�V�<��6;���Q
K����j.��+���f�q)tQot���ek�@�jL����+0W��}�IWc�l�Q��b����V�d���(��/ℊ(�C]��(�>�(�����$e@�IB��J���)L�7��ngͪ��eu��V'"
�ݤ��'(�@�-��/�v���#��B�b��*k�Cc>����l"�E�Nﺻ����lg���Lh������lƘ�"h/���t	z�p�0�%=��gC��f�0�y"�Ñ�x�=��+nO����i����a{�u�J�rA����8���t-��m��ƭe��&�h��w�y��PE̎���1H I������������у����ߥ���.����E�!�*t����o莐�f�>�C�����c!�����}�Г������^S�|6��O=� 	'҉�8c�Ux���}9�w���Y��h��C�:�	I��t��������#ŧ%�tF�V�NAck��0��;;�����]�t�kfj��C]��,����0���m\��L�`0Έ��Z`!T��3~�Ɲ��ǬH��&
9�@���5~<�̳J��~�<,��wݘk��b�yo�3C�Iβ̶�_���r�8���3�p4҂"�0HO,��6F�R�"��X�R��{�.�R�D��p��Ѽ�sq��KMթ�==��4�����O����-��q\xP���dfG}t�+/I_n��_m��߀+9R�ˋ�Ĕ��X��egi���:���5ږ_,�߱��h���rR�����ŤX``��Y3p)�D�"Ч?�8~����M=}jJ�:~�-
ꕻ:niկo_
yñ�i���kn�"�:X@M+B����!��J�5��_S�o�{��HFK]��PRw$��1��{`=�<��:�#NY���e���!%Pf�त�Iq�~&��C1���̘�u�ྟi��
�_f5�
�>�۾˺�c\v7�%"�����c�oi��T@[В�l8��E�MX�Zy�r���D)�����DTxtF��(�
F3{����l�,en�~��R�Q�צ�[DL���h�R
J����w�͇���SW�ʷ7� � ��\�lp[�e	e���Y1�����A٥�#[�؀���1U���^pm�-c�����x��p�hL�wOV��D��?���ה��5K)f���m6():a.���'�Г sL�6w������N�c�xwkǘMI��P?��0�B8gi�7�j5Z��	�'O��x����CSmS�:_]I�'�=��=[A�!��y�� SRŹ<�&ܝo����� ����D�� i�p,f�șILՈC"5�A���^.��m�B6��M�(�Ծ�leI��yNK�<�W+�O}\w6�XP�@Yټ3��}�iHbBȋ��*�;hU7�+�����e˞�`������o	��0�U������-K���\&���yj�ف��cs�[HƜ�l
��w�#l��ʅ��BKf�NS��b9`�d�3�B�!sc,q^�r�o�|~��yq�w@��{��
��g{,":^Mf�D\�e�߶_0�°^��" �sĝ��E2N����1I3�p|Ş��*/� \��	�X8Iz�(S|k/y/�{����輙Kg��ǻI����t�Ͷ�3�o	]Y�E��kD��Py�&-�@��m�WʫP���̂5!A�т���"��R'�I&/T��c�H
�ޅ�%d�u7�Fo��@..��a�cm�v/�.~��Ɉ�m��7�+V͝�"ь�=�\rw��ęu5�G�>wq.�=�F� ���DO�_2��i��J�� ă�S�5��%A�(��5�%b�6&��)��sT��o��0+������m>�N����)��v��,�T��ear��+�+��<�S�-�w<�RSlu"���I(h��ɢzt�={�
^VI{�cͥ��	��z�Ƚ����
zZ��[��>cI1L6�@�ﾫe���(���70�SZ�-���$�(){�&w0@�K���5)���tb^8k�����W���H���Z62	g�ll(̹����:t��(śMܔ��N`�ʯ��$��.�W�j�[J��C��c؜b�
@�"�t|!�<��2o�p��ʔ9�����R0N�s|�q16��!�tC�,�{�]��tѐ����~���z;�A�'eTSa@p��>�!�& �V�+fOh�X7��3p��f��pZ�d�O��Ŏ_�5�_(��YMɲU���CkD�n�H9��2ё�Y^����4a!��4����S~N~Ѯ����S�.~��f�N{Ry��̠�[�׾���d"$�����K簻>�ꚧ6�4U��؉���X5X �|�&��(���f�nTA6c�f<0���3�������I�a�#�iT�#s�1�=8���Ť,':��!������9+��	5�;��M	�u���h�˻U���]4<��St�<����N	����vP'A8� 5���hY�:'���igP�E4���{�*�����e�)h�!T�l�j�:���SC�q�u�<i��QTf���^�xH�X�����ڧ�3�,rA
��4ޱad�W�΢�R��6י⁝�,_u�H貒�6�z��OO4@�.��Y�L5D�Y�L��72��-յ�q�G���ߏ�g�RP1�7��7���J�H��]Jy�/�-�ڤG�˴���X�	xT��<0��*�:�����$�>�F7�Hd�$߆��W��n��q�c�>q�<���#��;+�����(y�������[.�B�!-<짼"��B����ؙ[��˺5�0��N��Is�
�u��D�Xm�X ��Z �2���{���ټ4_�Eձ�=�+�G�W�ى]�������Y��5^Z���tMw�b$jJ�������PD��2���sĥ}����z$�f)4s�9^v�ҧ=S��4�P_�*$c0N��r�R��K�}/�8i|g���2�U��T����A\܇�	�T���n�3�=9������&5I:�ʐ�J ������4gu(I�@����UT�x��g��Ȳ8g�Qa}�O�_\E�G�\ڛ�B�x�8@_H��F| �91�<j�UM���s�"H-��ź�뗊�I8�!R��A��� h !}�Q����p��V���"��AЩ���.�A���6��\4���dg�h�D���TG��E�p�=�_V>"��y�{�.�N����!-J�@OH�fI�qz����uf������Y�2	��Kdg�'�69܏�c��,NrE%ڝԫ�QM�"�u�.�Z�z�y˗h��L0td��F�)����y��3���n��`Q�h1�(B�ɶ6�D���4Uf7@��Ͳ��x4�A�rX�d:%��i��Ȑ����!�L�
���>����&�V@�1�UJ�d=8����#�/�aYo.�I���&��I%nu����CV1�-^�I��1�([��Ҏ���4A��RB$ӢN�?j�\���*MU;�鳬� /+o��������.���e-�Xe�k*���Ulc태�����<9b�]}��nC��*�ޑ���Y_�>�GksF1���Ⱥ*N���������Ho��n��r~� ;u�f�U����$�����j�F <�0�,_]�
b)
�|ߨ����+�q�~	�u�x��!�R�S���j�7��4S�=��G�!�<:P�k�m;c��Ja�e��<���J�gJ6k�8x�䥁��@�� �7�Wq�2N*��hԐ�ĥ��]*����lr�Mu��pѪ�y���vc�l����@0"���SW����~��y�z��)�������~I�Ʊ4�j����X ����'� �ɬ��Y�d�F��Y�G���a�x��ڨ��|ш.K���u[��1F/�9��FM�撆��N�L�y^��P������K(��N�=P�M�O���(\���A� %���$�7ݳ����hP��i�Jy]3�:2Eޡ��	�nz��q��ͬ
x�fW�8*����5�g���:=Ms�)�k�l�~)��B�Q�1��h ,p�
���|2��M=�Ĥ[���-sᗼ�����9�k�%A���-�930KH��x��D�ڈD>>��-"�+N�~�J�12҅f�MF��6��u�^�l�^~ ����ʵ��u���䂫l�F�3� �:n�E��R�֖��������nM$@�7rt��ӓ�_v�h��Rb)-]OI�l ���V���yr�`]���;i�J#�����L�)��V����US?�U�4Z��?�%�0��_#���K$�MpaJ�o�g�+��hpx�W��S��C&Nj�A��+�B�R���F�� �<*X��w�� \�N"'����H���� '}�0[B!������uE�ي���7W��� �;��F��r�'�O�W32M����s�#d���z�=��������㼰CZ6�r�V�dH�	i�&�z��H~H���YW�A+����w�<vFG��yf���S(��X�)�7�x;i���A�n`�B��[�_����ܓ��W�l�>�%ѝ���m�$����;[M��P��xc%��ྞ�Ṷ�+�f�*<���}�S�:GC���[fKe?�VY!�w�9s���_t^��l����w��h6���?���u�y��dw� 3�D����3���-	�ތ 5��W���rh�"e�kz ����&�G6�xWIc��7�y\�g`^�{�<�u�n�`]����xd<K��@�E����$�u!�Լ�!��A�{�^�g.�x�?ff;�ʄ&���W�!w�c���(}Շ�y��9xY^h?=��֕��������r�UP����ի������Z�ݛ�f?�����8:Z�gjxq[v�R'^Q���c���Sk��ࢌ��h6�y��X%��v��D�C�f��;�M��\�0+K��l�l_i4>��6G�Pa�3X�k`!ؤ�?P�m�����+�)
�vAM�Ο%������G�YY���ؠS��H_���v�O\@�ڧ�Gh�i_K��?ח��-~,���\�L�b�}��kM�j�l�4�MHjXU[�R�F��''
�/��=EZؓ�e6�� _��˱c�/���k�A��&({�Y)o�%�����XI@�)i9�K�dY�Dnfy��9�����s�!��C��}z����AY���ӎ�g|�P�~���bl	]�%���(S��1T\���zx�Y�����]%�M.2�;S-��IA���k�(���H~,Y��L9�#)+#�r���	�.�����/�`Gů��E���:��mm�����<�Rc�-u��!��X9g�
u�:���J����&���ŏ<�F�X4~�x(X	�_���N���1��Tڸ�{�;4��^���U����u�܍�̷�4qx�����ǚ�aū"6����m�wg���rQiN]�P/w�����ό����?�����X&��g���gX��"����cL�$���*��;���=?E}m�Ӳ%�6NB��N��8�ŦyP�F��x��%� �]Um딨��#�g��9������˻�Θ�UT�e�h��8ӲˇB%�c֝�Lv]'�'�Aj���6��|V�CC�-6��-�#��gį]V3Խ�텚n��.쁮��6*���3 ̺�E�om�����s���n2z�z]�~������}�6.�k$���: o���!�(�U�>�wF��]�bO����pqO�V�c;�Y=b��{h9�\;6�N ���R�H�>ES�7�caV�I�峖���!�߽�f��X�����s4�7�3P����Q��4��t���N1�Ύm�4���2�]�!��a��v�)�=�4�J��U��8�B����@����s���S+�Oǭ�]��kn7 FC�9��n�#��jpr�񊻾�I���,7
 4T���N
��ͣ�@�ɱ-��;f�����[�3�j�o��K���>��_���=��u>���zT�u�K~��/Lq��|N���-�$�-�x|#��
�E&끪\��*�RR1��S�i�U+�!�XX�qN�QqB�!=# d>�T|)^�i&���v��2 ;�M�]�lч���28'�6�0��!���������3�ů���U]�n��/�y<�&3�>�*�Slg�lV�as�9�E�]���#&
�>�Ymd�	�N`{U\�I���+�$oi�ž,�������3��p �����Q�h�`�<Q��e]A�����TRGaF��� X������k�jY6oM��m�.Q����QA^{@��׷Tn��^�#��ҽ+�%A�_����ts=8IEc�3Ա��������3��Xzl�'�K��Mb��Sz�tw����[��8<��2��cZU���Iʗ��w�����g�Bv!"�i��u3i ��#��Ťp��ۼ�eCSF�`���5ȶ^׷(yZJ��-ǧe��iUt�g���7_���T�$k:N��/.��]��&2���`�۳�7\�� o��2�<�o�1g�7�X���d�3LK!B�@}	��s�ʯ{�e'{BS|�.�q��! P�7��U��p7a��{7���d'6��nئH�q���ߝ���`�+PX/����3��Xf  �.܃o���e&��*���H�>4��&�1�g�����z������m[Ǌ���}:ݾ��8�K{J�b�|3��rp
�|�")���A�/��	Lͩb���B~�BS�����nLn���E���n��Iז�"⣯�.8�#���q��
�&�� 9��M���tm4�h=�����,�ʏ���t2����jz�d�+���{5@<-j��&���q�7��2[��kwz�H��CǍhئ�~�(�R�ež������:��oWG�`�W���#~���yjl��F-~R�V��-$�y�q�U!+�b�*��e�o[B�#:_h7{��rt �Ҫ�%٢ʣ���SL�@���Z�&�Z���j7c��4N��w�f2�f���~�^�H��*��B���a�ݱ��� d��'4����v�"Yݼ�@��?2i���}S���R�����>�/\ �n�Mr�W�m>o�N��'����5@��Ġ��	�v״��A�s9C츄��Rb��$ғ�q�+0��aG0��-q�O��<��|Gsnr�<���p 9Ycm0+-�Վ~Q��<t�g�2�!��g~T��"P�� tg��)qJE�y0,�Y�Sك[Y���y/�œ��zЈ�(g���Z�	�\������-6�`H�K�C=4�+�A! �,d�áʌ��#�\��il*
���쌮�9����îӡ}�{�[�2�K�q5������]B�X ���*O�!�������ՓK���HP�@4��.rP�����f��r�]�6�wvMp������3��.#�Y*�A��y��w�bV0�/��M�,cp�oq֋u �Sx���HbV�L�����$��e��r0�d_���*2l�f�zCGĹI�2��ZB|Z�|^U�~N/��ƀ��
3J�>N�a*4"rAm�~{{/�n:T~τ\+cP��vu���[��푾��h� ��*�eb�A�dr^���!����/h���F�E�Sv\>mu=���G�X���.�|�O8p>�i�Cb
���e{������Ay�݌���>a��(\DZ����N+�$�+baW��r|g��D?����|Q����Q����� �~�	�Ó6@����l��~��Ӻ�nچ��|����� �Ȕ��&w6���cv���K)�Ӫj�� %"ں�v�$6b9B�ڳ�	�X��hӢ�0�P6
��BE�1�N=�����m4�Q}�3�zy%8��#���M�M��OA+�bQ���{4%v+��<���
'�m��R�{��ӧ�jZ�hn�cV4��ľ@`-
ù� %���@��4?q~5�*6��3Pѻ�7��%�0��[|��/#�!W�E>�GʪjΝ99��¦O/�����MP.����Ϊu!�hB�GW]2ԚiVP,�����aU��9 �Լ����-A��{#�P	:��Q�F�i���<�Q�ZQ����w	�I�rq!�ϔBSf37+$(泧�m"�pP�,Z�ع~���i07@S>���Ϥ�� �1�($���&��S c?�% ���Qv���D�k�gNVԕkK�v8����n�>e�p7�!�?/�vmǍ��n���7�"�p�3��/9�w���x��wG�
�ѐ@�=(p�č<�yW�}K�.��H6��*������l@�})�Z�8:���=O	�ڠy�"7���CSlri���>#����x�� {o�M�V�{�Y1�F%���s#:ރ�⩈������i&�E[b?K�T�狦�\r�1��^�k7[��%��/
��iB�F4��@�ō�������DҦu����bx���*��E�W�i [D�fηE��ܗAc����7�7����1��l!�Ѡ������co}Ơ~l��a�����Ʌ,>e-�q*aH	�Lɻ*q�,/����K�
x�\�ԧ��69�ퟅ�UJ��=�����2�1l"���,����1�~�B�Z�\���mٱ��˒kr��$���Ɛ���,"5BܬDt�v�~��ɠ9�����< �l[����K��N��Y)�#��͆�I�̤��2ϫD�1�x_�"Ȁ��6vx5� +�O�+���d��;(�T�����V������f�9�uH����V�}�ԥLP�6P_�(�{[�1���3��n�s�U�J���cJ��������`0/ۺm��p�7�;�Pe�<��������6ޡz(�2z�a{Vt̫d]c6\�I�W��tT>cW	5��R���<�G��+7�k�UoCᐵps�f�|_U&<�m�{��g'��������C����<un�!�
B��w���*���/��@b�����j�ڱ�rʧR�o/q�&<A�/�鶨����8@L�|gjѵ*Ф�A	�y�z��r��ETC0���{-XjuqԻq�]��P�q��'�J�-����#QC4��1CZ�x<�a��4r:v�^te>�je�($T{��"�q�@%�x���%��l�V}�c��7JM�	��AH�Ik�T��jyih���6W��0��9��0�H	g{,e��$n�Y���> �_�[�2ֶH0��v�Nf�f���|�nx�YQl���;�QnNx�n7�#�Sz�����Bx���K#�h(�ε�׎����3or�6�e N�[��t��N��V��i����i��F�%�n�R�r
���go��E���I�rL��n��넂��%0��O���������ĩ��WQ����n�{��=wh��J��C�ڐz��+��[:�%e�w¤�~̽�8��1�d�F�7�s�$=��ȵ��.f��P���="�DT��P[����Ǆ 
�ѽ�7��_z�Ĕ�l���|t�2��pRR���g+����;�k�D�!'��p�E�.�����aeqh�oy* l�E�&1�а8�9|��z��(ޗ��Ă�X�QlXx8v�=w�Has��N:m����H҇~ёU��p,D�8�+$I��ɘ��R��9��,��w�`����͚���yHaK��� ��;���.b��9D�I��bi�]�ߧˢ���~OL	|����K�\L�K���ʚop����G��EO����|w6Z��q�A��s���8B��j�G�4�����$5�yF�6�A��N�x�dX����4�9ڛ��%�D� )VC�DKgL�"��vD�⩀�@�s���v���)9�n�,LRC�ƴ}�?���d�˻AA1\�fN�_a�j�"�.� �����ҶGW��
})��7��0��=�t�;��9ok�zHۥ>������PzƩ�˲ ��{&�CӜ�����&�������h�Cu��y�b@�;9�<q&4k�S��������Ƃ� Ƨ���w��!%$�i���υ�k�́ǔ��s�T��@��ݫ�f���_�;�zS��w�h�T2�"W�#(m2_sr"tЁ���S|1�l6�._"�2���{;�����d��+3SÄN"%�G΀^��T�gS�na�"�"��/f��F0-:R���&+J����樇�ɱ����2�'��T��A��A�����9%�
�������?�����#�2@o��:��
��t[Gn�������C��������_��j�*�Yi�mķ��������~��#�x?�󳹨�b���۩�Sر��,)�)5���/���VHD��?���GR�C���8���Up����,�'�@qգ�+�&���:4��������ޮ���r��+�#��hwOƮ�p.M�¹��Q�ɋ� �M��Be�� -���˖��>�Q�ӫO������֯㤞�j�bd8R�99j�x�᷽6r���س��^asb�~��J'�`EN�&M���\z:uK�zɢ���qd>�%�L#^��$�";��Y}հ0�G�(�tN�4���)���|�T��ǰ��'�4��9d�o"/�
���}�E��9�ً�x��0�!��U0{%������VT�N�����b�ȡ������I2=��U�M.!��'���C'T�K8W�쇪������^א�$	���R
��,k�%�,��+���.��O�rG�
!���!���R]=��aД�0��`.d���lN��@{!�/���dI`���-F�v������E�o�7I?%	n��ޓ>�ICg�O?��§%��~�؄+�����6*�5y�f��BV ;��?�a��O�	4]�Y�N2��`$���M0���O��*Q�[3<�f�G��O������~�>G	9�r��N�	���m����p=-��D�K��E/v�;H��[Tt�n���4�3�E�7�p��]�|jtsH���O���&_�M߄�������\��Nz���d�p@#g�F�"2~�A�Rh1��&�*��}�%�6	���E�^x�b�|�ﯩ�0����*ގ-�� ���|�E��r)��M.s,����g�H�_4� q�;��j�d4���Q&俠��?���	�aK�PI�����6LN��2��WK��O�Q4kC��(��Z}�r+�]&������1��K�G����)>1���=�H�Y��`2�pRP��XL���&�ٱ\��pqDL��|�b"L�U�:E�G��Q3�W���q&#"�#>����������;#�I��א���$�@���;�a���-�����V�$�r���E_u�W�����p�i6UY~]��ɏG>�%� ���K�\�L�*��|P�*�+�?��[�i�>(t`#�db�d��2�`��_�"pc�~����&PU���v�e|�׏Q�c�%!�F��� �����3����U��hC��X��8���؂ҁ�<v��n0�	���*�u�A�	�J�4M�@�����:���kIX�b�3�v,��q=m�q��~[@k�<����Z@��\���NK�j�wޮUI���'�
��&	��7�l��G���ގ��'��!�8��g6��"��{�$DD�+4�����Z7U��*k�p�7�����O���NLy��"Qx6�C0ok����^ϟ�o�^�w���&xۖ洒/���Y����zPKC�26������;:u�d�F��p%9w�ͫMb������t��J��a0s���z���`Ɍ�^�b��FY�OD���S���|�����&�Jx=����6�zL���|�`�^�'з}�w5n� ������g���Y�P�g�īX���|�U��5�|�1���e�0�b�au��tr%��؇Z��R���$e�`���©�M�sW��Xt���s�ҝ��Z�&00�����&��|��gZ��Z>(����S�
)V�������[�[˨�BMC�O�B�+bp�2��n$��7�����k<A)[�`ߺ;����N�bߘef����d�&Z�0-�_���,�a��q�
�L� ��c�G���'"|1�����U�}���$�#��KH%����R6��8��;�~�h%��k��)�}ͫ!.����+�0��,��܉UgK^輦:��`�D��,�G�o�ʡ&zj򡭧P��H�U�1̥_̩k+[[.b@4M�y6�R����r�G�0; d�7����x��=�|�p)y
)�iخVh�
e�!��H#����`!�5v���\P�e�=�\��ĭ};��"�L̞�1�q�|��ի�W5G�*{9J��F���]�7q�s�����%'��u�z�1�ޖ&*�)>=!�b���w��Q�/�Bc{�[�N��5|�3������UU� /Z�'����_׾SɁ�����ק'�mRU�x�o������bR��k�N' ,_^�֮�BG�X���㴀lT0r���B�Ӈã��ze�oI�`�'*�ޢ O�m��x5�w�+�y�n|t�Q�����R����*�F�#XU�/%v��Lt�虓i����Ldy[��B7���!3��C�cw��[FBl�<�L��c����Н&,S��:؂g}���8��Ⱥ�}�~�en|����$ZZΠճ/��g]���y�'�O�7=f�&���w���Z`��Xt�\-`@A��e~�&��)�y+&7���TIE��,A�g�'�+���:JR�5��3:Y��F�:W�Xy����-��'��_�~*��.��ү�,���df�Ҫa�|���˓��M�(M�L�!t��LW������c��;ڃP$��u9��h�?����b^u-"�f��Oc�ߵ4I����w�>�2��l_�D��k�}�ԩ,J��kNy�,7��3����2�8Пo��T�u���*^a�(��ǚ��vx���D��g�9ݦϨE�J���:⧫WW�0��:jGn~�K�j&ǧ`�c˃� x$^����zR�'��n�8gTm#Jػ%9�]jp��e.9��K��<��φ��]���
O�`���ߵx���)(�^�/W��r��W��p�gEP��,]����>��T��-vm��l�_G[�{P#���u!��4�Y�;|@p�U�#�X��D�kr���b��k��}T�=W�M�H�џ��T��_K�cH\c��:Z]��Edz��������O�U�m7T�X�D�S,?�z�=���>a���iPZ��(k���x��ɩ�`\�0M�JM͠�>
r�_w^Jx�u ��ë�ۜ0x�����+�����Q1�=���\�����b(�psk>}�/�!���Cp�����i�"���x$]@~���	�A23 ƊN��/F�2����/�	3m	"'#&�����ԫTg����{��'��~��+Ԑx=�"�H+��A��:L��d!�q^�`�7?�377��Y���oe�^�f�T�I�!���^��H�_�뻢�n�Q����Ư�\�ΰ���VZ� �yd�ߗl�'._E�_xeQe��i��k�I��s=[����C<jH@����d�@r<�xMz��9�`ɽ-���I�t�<���O��b�#���e����aw�
�l��Q(��/���lnZ���dء����ʓ�N��1�h��-uZG�VM��G�<����+�7J|ƿO8L�/������j;��1 m�8�4�q~���1r�|�_Ԃ�h�	���V�Ø��b,�FS�	���T�J9�\�ؐ)���Y�f`$&'��2�w��Rc��3�Ҿ����M������}�,���w��{X�^nf��,�U�t��]p�@r��=|.��щ��1�B�X�k8~$�ׇ�S
%�L��{]1H�	��� ����7R��7;�l�.D�] 鰒�~��[��7\���?J-�ٗ�Z�o�M�?y�z��oϒ���s�7�`�r;ë�{�Z��t2<��%a�ϑP���A�R�:�s�OH�88o�O��։����7��
����_�&�C%~#��}�����8�U_��8:��p��6e=?��t���4	�u�Y]�-(,\GD���Bҽ�V <��\=�T%"�%��T��V�o�4����0�	�dx:M!S�=!L���T�����a���~������qU�������z{� 7*��~�
zL���O=�s;c�k�8OO�[�����O�a��Y�N�lt��
��Ym��d5��"��HI�0>��):��M�;$=[�4���4�)=�o��2Uއ��sg{m��6�2���a��ǐ�)N�?�)�E�h�~���R� ��vR�6�*�\)��L+}9[��U?R��������-ҭU�?�7CA�j��]�yy��u�5O�>
��p5r��(���HT7���pU�4u؄�I�G�K!R���ڭ��qĔ����͙�E���`�u�f�U?ưǲ�a�����L����;��̼�<���$�ܥX]H�(���=KA}A���ӥ}��1�~�u�~��%]�	�߅�0�X`4���&�}�C��;(�9!sc���5��U���ж]�Y]J�&[�o�q��t�/*���5�}ǵo����G�	t�c�X�� J0J�aЄ��<�?3VV3[?��L'`��0bd�S
��u��[�T^� �Y��x��~�G��)\��1垚ڿ�=,�nU3�/��*�2�/���vhh\9m��T��<B����6
p�B�I/�\��]>V�c#y>��(r��JjbYe��R����nkQ�	�$ ���il��skpO��UZwJW@s'�E�ݺ�N7����4�����C��������V��#M�%�
L�_�h�7KR�u��=Kh���A^�qEhƐ��~M�V���+��lo.Jqb_2��y��Z��B��C	J���Eq'�A��邛��,A.Q���9��
�6��c�h�y�+]i31�%%�E�:��j��9u��|�@�+ɾmYLty���㺙�� !�d��|ӊ��C�ȤZW��}�a�W7�����W���S�/W|g)[���qe=����	� <ؽfx�Qtah>}�#r�w�O�����p�Or��@?+�[�v���\�&���X�{���"�1v`'O�(S�Q8 �v��'�$�H���C�Ӡ_5�p�g�`�0�L���@����s�%�
L�wQ�3X���^̆f��S�;Um�1Ya���q�}�(�+=u�y��㌯����,-;��&��y/�E�@������aw2�<���������ʫ8�j�N�� �;�Y��T�"����e��%r��B3��L�Q�G`��y~����;X$i��s����K��'�A�7�����/`�Z�������ʹ�\i�sO.�����ݡ��WH��9Ѻy+[�J�(X�:y�o���YW9LdR/vS2�tpzUp֘�G	�4�
�t���%$���8�����MQ���|��}��pʖ���_I�=`{�m��z�s0j�||���Q���ɒ8eֈ��5�I���:�D%���ci��:�����b��d�?q�K�vp�#�X�Df�{�6�Z=�{��&c�������m�#��{�Ѝ�L�ޚ-ZPd���s0��,�� �F�6:_�8: ���VxMҷ�{
�|���vHX�Y@=@�3�ڊ�b�� �X��n��n�Db #xLI����p�Z��<T��8fa!e�L��A�&I�曕��+[�7l�dK�ʍ�����oKG�`���� ��KJ�Z�e_��I��ު�P�=�reyC.z���r)�}�O�f���A�g����S��j��5�9A���$���O�~ae�n������o�I"͜�M���'i1�0~�J~&g�u�S/@�
*��A���c�����pQ�̼�nٳ�%��^�x��"��^���_�N9��Ϭ̆�rԗ@g�#c�Y�A��+.�Y!K����g_
x�䱌�O`/7R�j*m���?�h�*��Y�p����5j�>L��{�c
��M����ٌ 8��FK', ��ہ�#�={��`�,6A��a0gn�]=˂�}�{��*�[�_�f�f�Ov~X��e���
Pt�R7c�2���z�C�ż<(�{�1Y��_�%�y�;s{��7���fi�Ǆ��P{��Ǭ扣�A��ё'\��%�G�тE���㜲	P��Co3'�:c��L	`�Oz�c��#������!-�^��a�~���g<���`n���M[ lC���{�ԝk]5��q�gNU�}������JLj�c��}���q��",9N�j�d���p�J��/3�K�� ̻+p��^V���+����
dW0$��8GlP��&f�X�tl`��x� ep�%�s5�}ȡX཰N�?`���,(=:q�Y�2v�����tLA�Q��R��,`&r����`8��jt���Ab�\�=��Hl?��d��Y�a��F׏c>���]�΅�H}���O��qZ�ռ��x��Aev���_��m� (F�mW�!�"��M���1��dm��e������ؗ�����?o���LXt>�O$�g"Gb8#�g��#&l���\�B,<j{�c(
W�|�c���?lT�o��{�7jЖ��fݤ8���漅�1�3��& ��!j��� }:Kۺ�ƕ/��-or�ʧ�$���R�E�0��ᆶV�^'�y�fG�G!Sb�n����x�9u��R�(e���M��OX����i�1�nڙ�d����hR��"�hɞt��J����!���߬�v\(�9�^r��l ��q�W	?�d�5�iWvp�-��~13s�����樆�)!,��g�(0�0<�J�HyC��W�=���a��|N(�K76\�	b��p@�o��Z��?3cC���	<��-+h�<���w�(2-AʎU%S������M<����v�A�sw�.����Dah)n�f��X@���kF&��� D3�X� =��Ӫ�1��U�h���Z>nR��C� �3+�]"����YHXbe{�K!X�DK���E��3f�.h0b"�����H��������;��?�"�7����x=��zS�����֊�/:
A֞�&�Q.|+S�>�X�ޖ�3f0�ٔ:��k�"sT_���Vr�8'����7}ORZ�~T�l%���Җ�Ç�==�r�����"�%�x�=�`�Dp S�I�T�^��_%+�������*Kk��Gw|,J9P'��V��F�awx;�M8X�`�7��,9����6"�GO{��V�5P��[;�۪v���w!}s�n�ݪr�uP�U;#։��R�����~z��d1f��|ǂ|�:^��	)w�9<�[5�@�b�$��`���V��v�Y�Z�U;�U����\]#@��8��m:�9D�t[��*�,�^`'�A���a��_i+�_-�8�MނB���Y#�k��LϷ޾�h��^�_��L�����`1|wf�e� ��|U2Jy���4�� ��G�8��Z`�����S�hF�Qq��p�bK��e�vγ���ek���-�Ү���P��