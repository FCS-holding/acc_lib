------------------------------------------------------------------------
----
---- This file has been generated the 2020/03/16 - 11:19:27.
---- This file can be used with intel tools.
---- This file is intended to target intel FPGAs.
---- DRM HDK VERSION 4.1.0.0.
---- DRM VERSION 4.1.0.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Intel Corporation", key_keyname="Intel-FPGA-Quartus-RSA-1", key_method="rsa"
`protect key_block
nB0nBdRI73jasHOGAbF6he/iwWCAiMFf19h8W2wDDWzmlKXxZtsp3l2YIopdjRw+v3aKRdZ0rHlx
CfM1bO2LIf8jhMfHZpIzsn7sVSc//m4ZpGb4ceH25HP8WnyBSb6UkEUM7uihXyjOEVsT/1cw6U09
g/HqS6rvsrCepGyz45cYARaecc6xnNd2wtvDq4WANRY2xvqVilgKG8KZMsPfk693Z+uT21ER7Do5
2Q99jSVohiduGs0DPu7h/jSjcaOWA5Wmy0wO7kWRdFbxDVSgTIsj8WeN7HsxjbIiq64J4zV4BcXG
ZgI1QS3qs0JVo0wm4nCO719VbrtxsLyrGisfCQ==

`protect encoding=(enctype="base64", line_length=76, bytes=834624)
`protect data_method="aes128-cbc"
`protect data_block
mQlB3xJYx+kdc+POJ+NNSWus05zLvyszjl7HvQLWqARBDQHfa3qGlhBTvcoV/9RWCZvBYauxaMj+
+pkLJQ9YElciCEPp5JfjTvqeLzkXG2XswUdKCSR+oomk4m6uV3Kbp6pAOfsykwhvh6kn//zoxX0d
Ww+kHLH7r6ejOxLAEG1LAlQn6IRuqvGceQ5xRH7Rr/gvWeKPH0/Bwz9nkVZTH4U5ZTUCYhPs41jB
qLyEB0Ss2v/A5DMROq4jdqYv5QKoEKsO1u8Cn2OXr1ag395fsz6jZOHI9wWgrLVou596H73/vzwr
L5K3guO5A6rwkk7/Y5TbmS8uRM/dWxgMWb0LjbDe025SyxPO74r3owCVO/IzAJhcYsAv1f/YMDf1
D9RnoZhq/Q2H6hBxI7PIJXmLLEiHxl70q2E/zBAF4AOwtiu9nH3Wg0fs/wwEeY45cZNnuoDxyX/N
SVSXsfnGaXtPsqrE4HR5Fg/iBNiHu6h/AcBsKwYgy9FQwk9cNOfxt9IMaUYtyyeQDbdnAMrmcuFi
Jd7MbGiO+UigKf9EIfSeixNR04oTyeuee+oVc/+Yt4jfTf+ibbwWHe2SofLijZKrwDVTRPs0Oa4N
b+aWCwoB2QHY0M41LUflQq8dKteCkRY25aFhHxVdhBbRY9zkdQ9c999ghVIDLdtHI0zZuaQ7brNg
fjKjmGQscVvz7ESLFiFNH+Vi5V6KzoAdz2OEDUEGX3y58HnCLd+yyG7ug4T0ILs2VPjPYzpRfamJ
od9kxLnJpelIWanmSIPIDD2EQXdAtIq4U9wFcbQAihjGvC09uXcfM8x+z0+edd6hn6Dsp7MDMJJt
KrclAe7gVlumUx8mirRiCf4mpao9HYDCV4GsK8tIH+q5EvvpWdVOKxIRPgSzAoxzuQrJv9synpOt
ESZj6zENsqLG9UCd3o5wB4VPHpAtZdRSx0Iv6ZFTWGfwUM2vpQKbTna+ros1U6efT5zJhKq8CfR6
hpGIVo9hlRpchlYdRrSSh9Q12CpxooChrOk7pUwpqKu4Q+Z1sRKqVMpb0ze7F/Xpv2HZv4XKQIHT
G3joRmE1IztcA8l/L+Ztdr0DkvE5VDrIv+EQJsZe2z9i/o7jJ4XGW5iX8+3UeWPMOE1zmpVXDOqE
ow5CwuftMHl9Tt8x0DRycDnzUJNl4gKzzIvej3ikqd0+8/pLK5Kno8S6Pf2R3pPzhvOCTgn4b8pg
sBDM3cXRTvDWptKm7DF9QV8TIjfojIi38eC/iEjx8V7xFaKPxE1M4apbYzC7dUJAkPZmM5lERp4n
yQ3Iu7T12xqlzTrpvyFk0ZwJFwq6HCLsc9JkpiuiGjb5fL+7N+F2UJLxT5iV/dxQPbQOlyQ8ignq
Xir1uWUd165TglHh8BoWZENiaftiediW12NuFy8YK/jrqdUoBBaxaM7irIq7RyhroJk8s57ign/e
z9LOFdiwGu5RU5GbFqUNSviy/oiO2Evssa9T+WpgpdjNlgkCPIT+bTBDbVsT6wLNTnn2AUkQBifs
FG1kVYB80Hu4bljkspXXSjvQ/pBcBTJc5tp4APvlBtyl0mAYdD757kBktPdGxQBHHpWbnNe9PZPz
Lt85PYyUA+jpcJPQxLEh6qKYitMyxvEeQ2Tad7C9T5f6+L6PFz8q4jgrtJ90G6vRNBRcwgOfU4jF
ToloGD5IVgRUQnpqgUfh/lYtoyrQOgHLRDYSCGdbbINYnBPSkiYUif+XcHFd9NlMbEAL2wwFH05H
igHKPFsPA4U+AxIZGQQaPYkLbW8RPI8cZ9oorKFZ08/q/xW/EkIyHgcNlMVAh0m6Hi0YlIy8gYpb
oRO4jIyVp3Gs4AHvz4oJYR7VPxOvOoQmhpta26kkD1OqAZtYmGLySUBP6XFRFWdGX06fp8pnxqau
4wGbecGqSE0CUWmM7TIYwHz0x+/M1kI6ZcBsS4w2lFz6UXUpBIkeLvakgkavPlIt+03TSrT0M/MX
WEx0cFDzybRZ1Rjb9g81t45+ledZEKzY22a4FVnkL4scwHEpCorBlmagujUAJltRCsgbLjcyaM92
wz+gcH1H49DIl6naebbiIlRQd71KjVOkdFMGlWODw2j520NDs6MSbg0jZFfPYv1OCLwNlyyZg1vc
9sJcvG/WO7ZlZ0z2fImV+mwDEdGDjTKlvP12ILfywDrJECacv/Iup55RZ/HE7eJLH53fYns5zxqs
LzoEjK6uxd6W6bEiVsXHE4zQwMyd1Q29lFmfj5oe5cjrNamcQHUMfFIJP+PvkiYIsEcWvDVrfcOw
Y1xVN0R3MhH/LTB4bCZnJ00NxnYQre7A3UdMEuNFsZoPN6SeEccHYpFL/lJLIHm2HZzVkyDU3dOT
Ilkqh2SVfwSEF5ge9xggmU9iEdvbjSb5yYsCWgP7NYfFyrMQjVUZdxrY89jhpuDFpegLjgo/KvmF
Qo6iLKQvLxKGkc9GHCA4eCNVejubDube1juguRHxSfds9kU1mN7/EDgV2wHeeW4JxNKhIzqdVT6T
o7F1fd4rXt54aHM+WR+Yr+b1OF3nUeh4e8yGepJC2i1P91A4HrzieC3TW7dDK90oFnJWKUy/588L
TtrCMmTPheXu+cF5Mn6ZoPqOS8N1gf4d15tN8SdXSQDWov54jtXvjtACbHVUx4kgb46pozplDtXu
fjVNnm50qALBwQxM7Y4B9shFNzEcgUf5ZmijDpnlLtLXRSa9uEDixdLvFB/sm2R0uT7/beQp3tka
4bFLyy6XbqAO+R12hj537J1Uy0UPA+A1UyG4RQNVeTLDUuBXktk0fEYsVTbHobliVSZAlxdAv4Qd
6NPtqgmXYceIbQ9WWvDLDeKXe0zQnaSPm85HOCZw3yhQzciZ/uozKFTaTUykrO45590qo7t2XDH2
EY+tT+uFD0LvUkhj+tOuhlfrz2JaxPRBFDaNw99Mg6n4WXAEqopOU2/1jVBclQgQA8R/Pb846/LT
he2IPDgqP36GM6nY6/dBXSyOWptBgSM76oMt2R6rkLE86WnDhpB2vqJJzqueBuLRNPrQrQGZ/iGh
m/qpyPY80d4a6Yjq6FsmRGAi7l1gyLgtjituCNanWeWR6MhihuexG+Ulff04f0I/uJLd3OonpIJg
rTO3h7kzlCDKL/BbtmH9+BJBNMESdgvytOleaNSOeTf+Z1vVPMHhe6nxUOxftNzmHxPRvCv8d1yq
QXUocidWL9I+XmMkHbLuoCl/Ll+45nWHP88fjfHWIYqQs/f51pZ8kSaJnz4woh6Gc5oU1Vxy+8ZW
915gNMfy0NHsy1r4QWpL0w67v01BrFYoOvGkJeF5Arat0XmN+83kLIFbSM4npe1ubq/N4ax4bAi4
tLv3ibDkzRody/DuB7VK9EBGubU7o7qwJtrRjZRv/6Sw/TfjQtBS0CglZkbSJn54QwWc/PdC1Qxz
MFWTI69HGvlTZryAMkbErt2KgnS029c9a5TbUaRK8ry8T61o4NDgZmvyH/e9vMJrqnGc9rE2Na3K
KcVptH0SkUsXzMYegY4raYVcOGKpNFchTwN/XmrWCe44MoQ1C4KvK+9lL8AEq0wBrlUMluE6ofto
2dHIqJdhiQt/JgEGN2KqE033w3XPdG7PhINHOimdMoNKWYxbR3ex4MV+66CSubD2M9vvCTynFfsb
SfA/eQEztjcSNF+81FjXSk5dWK9JyEhHZjGMaluCIf3jx/CzqgNIL2KHsy9lwDtnUSC01Ou8oF6I
KzLFgqu4HsOoOkzl8LO1A8tUsLskZfLWudcANPX7ZM/TbA4t1W7ju1pqpNqterQ4WBZEKxVCBFmB
61jGYteZpJvXVkzYW2MsM6zsmaRRnk+d8PgywjcbYUuF9tZBFSO7q/kiCDpNShqiBq41zOaRGsSF
UE3Rxq005z2Rd47vQOX0p7V4J1BcmXmrUfsaOytJswUo/5nkeRbJE/ft0aMl5PRMKoiJjd58OdHS
9mDClNq6DkLDosGhN18wSC2ykbdM3jTuKEJZks8MlfxzVRs1AINE8X7g9WBZApfF8Ri1qkxRXJKZ
aXuQzz8i5VjyPb1UbOglgobw0K0jtjIs1lxAtqek36lDEyfc58bWPwqnA/EW/8L4hAzXBzNATb1S
jj1IOtCej5sMe4IMM0IJbhqBjMAiZDXglNpDnpq3Vq7SKpDUeIWlX9tES3S05TGUp48Zl3p0wbSN
FNZF+HATZLCi4PfgERPEG1n/cCMrLvmBTBtwa0Hh/MKC11uqIYJngfzvcizETci64+lhPJhYKC/h
7xsbJ7ibrlqdd5XdR4ZA4mEfg/HtReyHcjd1IQgxhCqhMUdsoVtPGAfwqUPx7BR/Md641WIuO1x8
2Z9fEDsD4eWGBcQ8WDxIZ0RqqUWxhpe9n+jQkU91/8QzyIJBCuvJJ41R/EIPCKCEHHa+W2O9CbLc
jY55y1b6fWWpC/O8ARgpXMGcR0GYgvxicpGdhuhkbzkBK4zS1KnlKU+634U2bbktd/MBkhkPCsDv
JxuRFQrjWD+JqXJ/OCGTLG19451RV/RE7tKYLSrEGrKyTNgrvGxVo0XtpgbvWLNs6Fzlh+KdQdQl
Ze7pJv9EmWwigBl+m0KEQSZ6Q/+BfeQan5uatZSvYp35xrahzNWEr4/+F61yl0znjbbs023n8j+7
6QVEs8s6CIGxZF80qHFwAMFckMdx2FqFcntrH2wSxW3y2v28XSj9+7kKaef9SebGdm52GR23uaNE
hb5R9hiTwpDXOB5ckAeHBRUBEnlwt8es8PmsanWT5a1Rlft+/eM5X+bKUThGdCRMxnWSdqXFMA64
7FIQTx3eTTSgtvjYN/Z1w3bJgPFkPVwQUN5zLH5uYvT4eGWAduwjbedilICnJ9/OYA7Jj/Ie3qgJ
YRvUqOE6CiYKa2K5DTSwFEiKkl33LM50ZHYfIOAeV3nps5BS/oRCAfAcw4VH1cfHGiKKR5Prs3WK
eYpZlRiYQswa2IGX95Syi6/k+u4hc5iplUrKmJ9zwayxxgDupIvMN91zExgiLRmBsBgjcG+TcFxw
j7OHQ3Tk9eTbKd0XpqwkzTWxS5r0oqWkJOWBCWFHp1bFbR4aI4ie/50xnwJc4Y77OgO6ZDL51X3A
8zYbhKVHUJNV3QZoue5gqFI1ZH7JpRgCHEjqVIq75KjMLlVz2wVXKTr4PxGBTwYH5t6Uj2XRuNPn
9L79YzvKlhzftQ7UV5/jTlFtsJw3vt+Iszrs6ZsEVlQ9CV6a4ny1rW5oqmaUcEQ8GSqhZRzDT8r4
TtIa6I+V6fm3ORH/7wTPO37XIpc0AjPEeM9I1qo+JrMOV8AUy4LZ+4jvh/q/4EOllxS07a2HQ6ZL
joIosspYbl79QIxv7UiVkVUVyFCa4WOA5w69y7+YeHytog5kOPIfZVA6KbdqK0KdQW79vjYTBzRw
yhsGke/tL90DfUTYtIK1wLCmWsKB0dS42MwYfA4kgcC2CH0knmrc1Bbg1s0n88A1qKIjDxunwIYq
918S2eArxoOgTgKn5Bb2CtcaQUQSnTi3ejkID6n47zDdRLXi1sIlYHpmdGBe0O785HbK15ajClad
5+8Z7DU5qavPuxlYOGZF+vyXqihwLkccxZLJeEcUkTI9A0CfMDq1I6pDkGM/uNJpDCfC8/fe8WLR
g+r/WK8iveDY01KOUHL3/a0D1LAXtcwI38SXs5kCxcbhANm+QTPMp4NWI522QtpfdTqiXDzJvZet
KJR6QhuU89KZzfBGW7piNS3YK1t7Rlb8BiMykjyA3V45xFc2a4olmde0GbmLREYF1NYNYX15AfCA
fXx59Lm8ZUIhPtDoEVQJjIjLKC55CuNwOYK0jDfXMXaam+zd0bpa10zvkw8xo+IfkvXVzOq82dBs
d0Bxfwa547p2foT1PFJ5Dr7T4d5os4tUaOo1UUr9E4Z7rlxL4qhnzAAX7KnQ8l5KFWHW2ek2L/UT
RD4yYFa25mLM0saU5yioncMF3Cip/vVhNW1zKNdC6h24e8hEVfx0KWyY8zI7p2HEd9MqmZyheiw9
Aa9gxcxA66WWso8V8iP5Sgib1BojnK7gmn59Y8SnUMwZ/vwJ/Owt6hGxTCxgZL8W8wyfzBWUQcyY
d5m3UfU+zLcOtdz+h+Q6ZvbL4KDZSUNnxbajAE6bvSSvCuqFC16piCk//RCw6/FBAPYNsVBDj6wn
tKNxK1Ya6Z7635AClVeP1RT+tIJ379Y2UkUvjACkk7DvrFmXyecQNBeCJkylNDimxrbEu16PMjPu
CJTf2F0D4tfb4DXwq8jcQhTO7HYenPN4Tp19SYNxy2wflfTbdmVpiWexJiGaA1kkMQyRpsD3W2T9
6BXJZq9EOhiDBnVe2xuYbV5xrL6rEFZ1axu19x75in7GhxKat8um2L+MXhaOi4hNm4DOWmodQsdr
bG912+XS8YO2jJZ0ciagbyPK61zNG+Uerif7BPudp18nTKoOuuFnADBeDyfi6MIwMCAlGruYUxTC
J9M6dZp79Rbc4YNOSUllG5dZyYyEf5F+cS7JCuanmS7GPeWQZXcecxGJfziTlT5hC1nTiecUp/NF
YFHqV5CTWZ3J9cNHhWXe7UJCOM5YNFxc8Hh1aGBYg1Jrf+OLUH2DW1OnCvvWpbFcKKoyZJAaRNDp
wQ9P9Ma7TqscwBpb4V3nwSd1KO2+0HgwdYk2kIRAry38J889WO2O5m+ES8xbXx6GjDkdwyeA2C39
bSR1kUofGTMX5XCvzkPhXNMYfZ9okzZJyXCewhPHNrQWD9y3qh4v7cpvCyi88WH3R/s8stCgk6qs
mioJGv2Aeas1Xk4HB6kk2nn/343jlVWA7fiEdfU75I/fAxXEjS0zMsjQAmEQ2VpOmO+H/KuUo2Y0
eOIpFB2VtgvkdUH0vnet0EcbG8twKHWewaoUZYPjDkDLxIngCBj5og4wo7myUP9XV9d1xKv8IPkl
WcZlMOfW9F4RXMqpYf7XhPEPymKdog3zmtmqsqpng+OZqsi3++vLz5o9It31G9xs38PEe2txh814
zV9u1xgW1TuSl8Q653bNwNt1LTbCJEWaR2QQwZN27/pT9lIwaO779O1bGlQBlXag9lk/HFjHBpGz
fh1IN1R9k0ZkIkKFYQ2sadIlclZTZQOgAo9qNmvvPZkU80iVNbrA/2HcimBR7swJMgfcEWPNi1R4
MYP+nxSI+pfTEfYE8Mc+k1WL6KMu+d/OHmCEkde049Y+mJQQpPvcu1ovfC/VRfrgS1827tZWR+Lf
Amej9Qk4BqrHi7fnYrYLMYNcsUbqC9tX4/6fY9MY/XjoZW9bIPgH80McvStk2iPwVZrTxFxvsVBV
IO18nEEPNKdEqLqZtFIs7p/HM4pRi7FNtC82Tt4zJzsYOKnoIIe49PhaltVO4swFPBRpUgymIzdm
nkd+CfH6qUVucWFOGbPoqfHv00BhATnU+OdQgqqWuVXPAbEjtWJBiejuTPqIIloz0HK98j+C8n9l
kauc7YJzglqLyfNoCKm3NpQWi1GJ5pBJdO8lbO3XNg2kyZhG8QiF/oyKZ641tmKStQ3iUKg2GAp4
kqViCw2lkECou6equQqCPhCONe6fzOWWpySQiCyLbj2VtebcHLjANaxGXdzTKkdtPx6MCPJyRNPZ
yNldUfwMIMYx+bD52TxJWqqdyhU2BCrywmclmbUQ14BOPkxQw6Qa8thrtRmbgO7D77TeV1KKg1A5
6wCWuNdnXTRzt50COQPSYsdYi42KKKw1jHi+6aojA7elY1jioMfxmL9uI5YQ/3YCBbWtbqd80ymI
0aFXFheP+kocOeAY3LdvLUA5p5bBmxkgRTd1A3DK+nFYqYvZKmYAF/RHD94ap06ygp0M0pppb4UO
Ps/FxcXu0bXbukl5OGvxgsSEud5OaZBOvwsY0D8XScfHCopeAa89KqQ7B+bob6eQ5tnm9Ps8vM++
ykkBLc6yiYhaXYPUhVYdstTgycCLRqJUA+QVMdEEQAHevbsZ71yyjge0JlMtXmgd3lDL1nRDlrM5
jE4YikzxKy/5vwQUB7iJPZZBahWvbIUyqu5ZnZWGogCin3d2nSZ6CMGNlLYEVOlvR/aU1jkdSHdT
wq2lTsFovUCTep/gPKMUhwsCAfmK9bMpgOaHKAlGnTuYplU7dra3re6Wk5mXeS9D2YAcupYg9tCs
heEcz6XEULeXgi1CGceYxZTG4y8Iq4MiS3ns6FgFLNELaWJsZbbWRlo7q3AycECpcujxigaGj/Mq
u8WHV0PaZA1eFtm0oXUuWLlrEJ3ztg4UD14GlNFfQURhS4OmLBkldmIZv+Q5CwjqiuSmjHFp7Say
7oYVVugbf9QtSxk7iy1259ikYBorGZ6VoNeIhfjZW+3iX/skyUEbLJEO+L5Z0kAnNjSxjQ40Yw9V
iREON9PQbfRcKFiwPLTcbGPlNMv29DaMOxwBuSyoXeyC4NYVR4X/vaZq59IQs0zW1AG72pPAUZ7c
vxO1s98Uvhq3+2t6bWYcc4yclOf+9pOQD11+ImzekjovbPbIqpuT1KLtdARZn+v5UlD4AO4DItak
s8AfjMJBacHWI77oYZEgeQJEGv/a1998/uTxq6J94n2GNKL5TiEusoTpv3kq6qBSrIMi0d20w8tN
OSEFhDLkCW8YMN4RztAaGyxIIuWISiM6QANSUQ6mLenu9SiycxwWWg2Sm64zO0CpjnLahuL7HwpA
Pdekd4+EKZTSAmkbFM1U4tLaMFDFxKqotogBxT67HH/szrNuMUspDuZKYCj2WN6CaESjK2294XUK
D8zCBjkspfeZ06Pffefc7/ur2I1XVa6hpQOj+2Pzf7FtS5VZHa36i9LCcrMbHVS35f8Bv04lGY3y
AhuKfenXdSlKHI9aD+g4RhqOWc1/LOEn3ryu54dXWTgDLzRDGhnRl2vytMd8FhNLu6SXxusZ3eBm
Yu3sP/5LCRbdc52+0+dKCCxvzbBHsnXXpz9dFGcN0SSFnx3vLdDPe+9TPR/tSod7p8bsCCU+mpjV
r7iyL4y+ZFftMQ0J+PJFPv/IFa30/7HRXxhWKY3efK0wVWAv5qngyT/ZUd4PEYQ5OOQZOx22Iq52
Ol+6Yy2PNPVD8nXvymX+hIapo99oKeyHdPBFCwNyPy4i0bm7kHn8ydhabPLzRKO6xgiu2x8KbMiM
7VaSwogNqGOwQhylsoz4VNFGkU2u7YibSgBIGk4tTWUlYfIzGItHrz2FzYOBn+T3Ju8mZ8MpYqIG
1qtYPl7PAHpFx4t6zF1Oq6IVlWPDR2jRmNFFGBKCVjsZS4fSau7AkLc092vEdU7gtFAH87NAqx07
5AJFoVj61rAFMQ0dzVr6OW1bgBnC/9H0MpTxg1bfDue/Um0vYQZBV8U1If8afQTWCGTTwAwNG1Ys
brrf8ngWHNaqntDzsxOPYweWMH88T4gouA2IBQkS7nTJx9vTXWR3ii5ZEEiUMo1FwfnRnfFOz9X2
/p+o3TM7qv2NQxqow0/nH6FWkcPrHfWB2dJX/YmCCsfKtCAVj7VvytqxzqFxWfi4tateX0axVuao
iHyqbM38avJ9F7flFjbMVIxddapweqwBrsDRvHwghW1keH+hRTjePLcFuuzFsyBLiWrPpP3BLoU/
I9+pceG+dLg4isHJARQTYYFZzwJZNCCA0XXjjkvSam5IZe1cqhroYgOeNtU/GD0PH7unAFyEGbWq
5n4ClXRLulCozRcjUqTvRLNHO9i8CVATzLI/GpCB46gcf7kXK3qHgIbk5PdI60ffGK070nSSP2tQ
i6caq3MegSWSsJaRYXEoLoGbjmLMU5WWY2Pf46NloxdCfujt5+3IWytToaxqmF4+DO6QcU0kHyqh
9WMeySJ92WQ5DtZNkft+Oq863fdJ6WxXsSrtBU4wHsXUJTTIiqkKlu6LgdmgCB6YR2uJ98B1+Lz1
SN35slOdVxnCTTfmuGGBKZ9L+xr8QOzEQ/7VAu5MSJR6ce6AFVeSUl1YcZ/JV0Juat7qkaKNWeMH
N8VLJZ0NCqmVtkKRX9hdsLNUqRakVesTyAT87sbBLUBagLk6GnjILyDTAch62Uo9Jqm5brdh5Z29
GpVwfXboU4pKtDtk6csLlOXfa6SJOY4NGJxw92MSw15SNBmad9xwFxwfSouFvpzuQqHrr1mbA0no
xy0C0vjXqqmqK7gZQxP4kePvBaHFfxND9f56enz9fRBQUhzXGdm0hUUGmJEY28kkXhNuKBg6GMc5
rBYXSDqoK7sZbp4MmvLkZlf/ECkNlTzUVMuJ9WH2KqXdZWiJDtz1g5tPbg7FhwPvaIhHSMWNM98Y
aNA0VrokuHbMKADo8bGPXgTvYP3cj2shn1m3uQ+uz8tYa0tV4Z4tniYzJ4neHgYql3cdlrElaD37
rJNLpkCzhJZw4McoPgaMo1Y5nP0yjatmpXoIACSZzxOU9wK2/uyQ1cg9SQu/x/75W3HTsSeUMUWL
wo/EgDKa44olK6BkSgJXr1H/E0IF123DbrNjEMg+EP0dhTruMPnRJncHgLwTe8dpHU/J4B/6ptqU
rjJd3P+KIGPg7XEZfNwYuKk4Gxh9LnKTWdMYl5Bo3HkQtQSkU8JgDD6JZhY1CBDNynLEMKXQuStT
6tHA09rq3una+ftDxq+8YjpHmkHKNBTzwyuXkEA+7Hy0VEtmtXuP8K+782DjTa/591AvmLEEhAYY
/9GI7d8jWPFspY1vugTQbGa9L72xs56qYwyMKWybIyjx0IIJBbbFJmdzuvbjs6rntBnVdX/U7j5i
KstRtW9Rk7Qo4XEUPzkAESrV5ypTWgcPnRDzEluWjOP0P36GxzpAQmkZmK05oDCE3AmeNwGzfKPS
2AcSTHF/SKJprnHyJLBn/hCnkcDIAB/D0hyzsksTaQZpeJKa4+LDMcKjvtykdwH45YrqlH8TPBCC
zuCsV4abklrhJmVLgifgMFiL6y4HhxVTlop8fX9vYVsQ00LYXOJXG0w5w18rQH+z3jfNLmupd8eR
FC12AQcAUkTMxJ0yVQdKGsoq87zvymXjXA9hMaGRfpCgmiyAtRlGigIWRT/sc2wlY50d6h3a5ZeD
pk9zNi+4aW/i9i9P/cFUjQ0VoOopD4N1esglMHD+mPz/7Dw84+ZHzcq1JSeqbSZcedbTxD53IraL
zfssG3ytS48jAxVQS+iAgcTt+JqYjXb15pvUojtcWAK71EDjCQ0T5Nnm5AYEiX6SeUPqiqOJEjpf
bU8EIlKhaIYFS71frU3/YogWegGE11+mhNHxk5S9u+dpVPr9ZAqzA92+9awBRIyw95VuQyG9A6iJ
Xg7/O7z1ziOnkaNw+aOpDg78nLSn1nrHl5eMWEzvhYGPIG9UbFThdxm51yPRmGQKGfgfMAxftm67
2KnaLuBfzfsR97jDuhMkz6rR5jL1AN2D5p50kwLd2xf2UNiEYieaER0HYk+Sd9J00zDsyjk130g1
8Sc7wUx3rz/2qnAk9e7rAVB/qEY+miHmEpclMe7qnZN+6HaJGIqysNztmpkxtF5Yv9V9n4Nz/wen
oEuHAYJTIkB8RC0nzy/emEwAo9WNdimeDbeIdfaRFMME7Xe4CDZ3ZJhKP1lUMbG2AT9rHLg6rTQ3
SxcWT+5hes8BUAgjhNa55wSzm0Py7HKyOCAmtYRlb6wBzAs82SXueiyedD2+SwoS4cY0O5sinN/Q
koXt/atAQnVPgH5DCUPWLqZQi6durEpplsu70rvI8M1Cx+yimdzAcrInq3+V592HNFQYBlQGmq7N
6YhFShOKfdoSxuCs3IzZmyb5TvhKU7g5MHPnxBqfP+XJUTTbpkCL4bZQXsht3yHzbbjsApJ8+xMt
lYbbloifhF2dA3P+5KYg+/P7wqwjXdsUUpZViASHso7c8hivSSb6VCYzNGtMW2ivVaWoZoiIJrv4
Xvj+KynKcdFHLtsS60WPgyiqLhotIz6hN1pj2bAgIRfVMwtC1J6Vl+YQdXMk36tCra/BTUBphCfm
BbMXaQYv36uyHccwlcOsAiRPR1m13DPf0JHwKPHRrpntrVN6vStDegAgypUFF3PYlDB9tqO+xq2M
iErp5J2f85jlT8JONiTrstm92+CH7avNmrxbbycwKgmtQVtMpCuuB98DY4TflJQgXasLjXjhC7iM
QT+QSjmlUpFTcPTIDcpyLwavtFs/Q/QLDVA4yJHr60UN+00vMdpxw35/KD/8nlPXHbpjpyzlcQSq
6M7q02Jpt5lEZNDGDTvawVKx6TCzMfyI2EL+FI06u0Vr/QAeBqvxHEwMlcJPyTDLYKN9bHFWEHkf
ebiVPOKEwaHXsXbrP4RmMK6+k2ixDovP/oPvfWvfnwNsV0VARYIcDGkDp/VCfr6Tfypzb1k0YR+e
RJ/uFkOX4dlnLCfrrrpG0F2EIoj+uDbp6GZjSQTjhTgJwCQl2sWhaZcAfEeA/YfYSVNwJuYNdW10
PBY2GAFBiWlfNsF8Bsr5kwOXOYyFFhDOhtlPZWrQBglKaPCYAEaXdojN2FrRjm8yQyxixeTwxjsN
3FurKDuZTyby9bP7RN9fVi3BMbqw5kpOvE+FlQ3TtrpcXW9doFcvQWH0N6AFER9+Tpp+U1GMnDo/
2lLGYB2ONqQstJpf7tNOV7HRspZ4z1TLOMbuQvamGysMioYxYxFxaxi61SeDveQqM3OXw1RphMGr
F37Lud4cmYk0RJZpsxAibI8Ey+ekd6XEkztUdyZY13/IqjF0+PutwKvmxFI1MPRCoyh7I2EJScbj
q0Yogh0HXCf9iURB3dlQcENl9N7qoLby+CaMR5M5+mvHjktXCDL8C1YHVukZcRbPiZBOpNpXiVgI
oRwoTwBI+gbV/pJg0EJ5dVv6yMAtAKrRWE9oYLyLy6w+fI/hGTDQVUcbIgzFhrwwWjXlVyk0mPS5
4Y3zlJ/8Yz66Lx8EhbaBjUm2miv4Nd6ISRQaoBSjMzQcO3TFErbLjkbsHWy7bVOPpviVvfY47+pn
CuAwx6U8uGUG8zWVr7HGwxNhGxp3GXmkhr+j+yBaYcf8MatdfJyw9IjGQG4S4+tNjrTCrL+hAtBf
n0bVlAB1uZTUAPZT45PkPmlFHHv58zGIctau0LedMmcb2NkPtwJXFg8z2XcCeAKMBrEtawFgARwL
F1z2iYcjRtHGI08MJpaiCLEo6jT1WcI2EftZCbEO6/+DHpX9pLXmlL6zXXZ0rb3GbhHK2lhv95jV
ASTpVFRk7ycFuZgbOw5+0Df16lxCa8JsFwue9l4dtKBIAOunRXCYvzHH7BLSvqRbTeTqmbBgpUo3
2iQFRIB4Lmn0mkot11PzhH5bASo/VRcO4rRDwn4MtoncYihl4qyggKx7gxJV8Dbtlg88ey2wPYza
3A8H16D/LuPkokmMWe/xBzObGSRVTTBE79thiEGlFrzFUv5K5n6v69jcVZZua3iK39YRE71vodRR
5puhvlgtJy8bhmI7yVqjsoXouS53ERw3jEBNVaRMnF6AuQQeXwuT++Eq+/eZsFN7wQlOehZjZdEe
a9YZ1ugUUsZKZq21npaKfE4PHpOpLt2hkQ5XuuA7pUSh6xDTybv6/lwIKywNkDDX38iqdBRI27ng
EZCDY35/SpE7TCq/XeyI88yo2vQL4Vz28pShFkvzHd/cPfUzifig/yFWSPYox/kJPOg1wntFZKgX
M1+aiYc6MNvDZ6k6qlDgjFRa8mE+n5AL3vg9xHNNEUjMKhYR9hVyG6r1H7YCuriZM89YPyPZcYfo
VrK2AXXXuQJpduAdE55JvfVhVlWJxhCvcRr/WvN/XWByvrBARd2GrZ/cwiXvQcFFJqiD+OCWfUbq
m1WwHhvSJPskeIZ+ZvqO9m3muEGCdeu//xsfAG3OX3dEHnXQ2SnOz+IWlzohTAEGgyIxICLvAh7Z
FXjSd8n3J97PbSlUSj6vaEtvpUxLfdhk5kJCzHLcAoPOZqjmTaMQUVEQC/Gy7U5nOniasRIMCPMG
coo7ueSEkW+QcZnycUeJ4dvLzKdXLEtDtNFOQEuXXlWwRskTt/LdldvuNRlmvekMnKZNxwGpbGvf
qITeT5psu7qDUI+NHERrGtb+czAuVGWNAqqDajZmmYJFDHgKTpgHaQw7krqBBECWlkWGFZ3AGePk
25trF/ZZi/sjBX31YQTHFpz1SKug6mjaMg/yx+j8NxqyRO+8wAmhWW1Gprrj4ikXhxubmGHNxDKb
FWqtI2y3sa1mclJhZIRmkhuzIDoDao3t8ll4OW/nvjLm5ZpYz+UFz949fK3zcpRPCiXJmVD/q1hN
GKJY4P0bRW4sYLsWuQcT2JZaGGTq8yLuVzSzBVT4wSGvVNcPyU7tFSB2Y1dVesYdq9NoCGX5F+nj
LHKuze42kXWYOOuOL+WFXcGfGbUuPY0/oUyLr2hhlijOlEqTk6vza0F9NY/dUiKZNuGhJKJc3MxX
W56db3udyvK1uEPzFy5TImSyGMYnZw7lA4onXbIkC7B3bn6nTn5ko3tQV/uNoVBywmhUgyZXW/v3
6PH49SGo5HmP0fZKByCRE0aw+fTBbYBvFcGd6Fed8YK6t4heD3g0CydWXSMUifl+cIbL+G6y7N8f
FZmHUdo3io+dr4T3z+MJum4NcbJnmiSlP4cvrwYzeYDGh1J72P2GO3Xxijo9/FZIMIZfMquNDfXb
CA311oPBMzv6t4HjxAUsbJTJGnE3xlOjCil87czSQB8VDu9yiYoLXRCWPo9cmvF8nMBEUHDeHX2K
F/kiCV1JH47MofUIqj+zcEDW9MgtAYhVyFwL4aV0GOVZzZjtWQkp/0mEvLrWyiINqw22yVqQzVWg
B4k4Lh+qSgVsIi/yihfmnNxWImNBNcERHJolR8M2FeZ5KWz6lh9bp9qRwynHCxmSSJRX6BiCPQhA
k5fubq94Yo5YEOv5aeufz6NmbI+eKzrzSuyomGQPhw1l2jK96UePmwySRfVWV7fiaTbOGQ6goY0q
D8rzudifEk86K5hfcnF+dn4/SD4Ozo9tdqfS7xDsCYEG92UC6K45S5i3/4xWEdhzWvc8zjZqu990
qN6BD8tTgz5iCpZVWuD1ZDdgC/4YYe+MNaH/H4uLdTmcW8JMcw9kM3G7dmE0mIrEu63ORd4U/It0
f98xZKG7nAGIEMvA39cBpXi3j9EZxgj0bdM4VuFIquDpWnGGW/Z7RqDqM+m9KjX70NfCVdK38DIj
98GyTes7qssqaQQK6awXNP9UIG0U/adyq5K7u3d53AVxkAhVQMb59l75XWcf/GtVX4OBlSJ/2h3n
h153Zso0z7J+59aZsctF7v7qe4Tdk8QxTiaS5p/wZEkJ6Iuub7hTRvKGh9zG0iU5k+Bx4WG/6X+A
44IxbOdotwdYQlmLbuKgV4n/Tix5N+4O7OZKwYXHpfNqrLNl6MH+sfxzCcjS41wJDiPM23nz3d/8
9H2pNfsCHAZRh4L6evA6uBRx2roTL7DXVsjZq06SwQhUilmKX6GBL2TJDyWNYhLdPl7HkZyYnOT4
nT8QDhT+z539qcw7AQSq0pT6kXmpi74/ruUEEe7IaIJjzZtDSx8YIWwlVnb44Zlp0eTYcs3pPvGr
VNF2/vc78RNGMsmdH6xVCNJ2cPsH+O6wt+xz0vCcHfiaOotguFdxtjFzVk4R5HR51GcWQzDtXiDW
cuSkD2Ey49meBT9H8c1QmtGxIO5+DRhVJ/PTrbXg20hP039gOL5E6wah4z1/4FdaWHJ1p2IcVQBf
GO2tLaYCxgoI5+m89AMWqGyUjKeagKS1mWrWO+JwFsmFst0v3ANtUXACcGhd4aCKYia020K9T5J4
Z4jptYb2ENweuVzelU3gtQfJnwGLyJRNwkYz0zU48ra1wjz9h638JrNbAso4XEm13yznRbyR/KHe
m7+rhiNpj6/2iVOri6L86FpFuGoveR1PqKv/+tw+aSXqTj5io3iR0iWbO8XN+ZBQGKvpzgA9aY0u
DO9ryRcqFoliOl2q5RZkkyJAxjqwXrVB5lYq6MdU4fDP0I7Ba1RKRINgLNCXyLdFpVRTz0kTbeqE
7FQKXZwHszSwEPRiwXCQqIDgIzGQYSe3lBT0U2rb4NjfVNA2xbjpttXNbn/FFryB7RW0XDtUEahv
FqxKNblZZ3lyS6sV8I1cvx9DuXE69UXC7LB6Lo4YudOIWfRPHW9l9pkaNaPWiMCz2doc+NNon/P2
yuPBO9O5QoyHfbUHMjKGBXezIjm0to8yFDZ/0Uhe2qNr3xILNZ/wNtGPKyhBuH+xlT+ZSzoOo/Bs
WHPhRGWDiJd9jb7qB71KGPoLkqZ26+aaUKHsFLNYnUHfGlI9oUObPg9eSfdUHPIdxpZxbepiYHEn
eqNawItdj8XFvmaaXjkpPbpYAjrLfx148MGgDeqBBdUJInU8xsz0Rgex+HteaBnmQUhsiVFwKii0
FrShXqt8/fTEp1ibMbWMED5Dz8qeSGI5xicXmGo4gPCEMtRDPM3EWv5TkXufPJZjiVuAjmW8T1P8
e9UCRvsZF+1uJIYtf6cTZ/Nh/+3RwJUe9Kn2lgSG1DNGgfXn1VYiyiPYFWe2HWg/5ijeWU0Dk7PF
L3L5BmiYG01tKrB3a+xYxD/yARqpAZ2yMKjfJiDDtksETo30yAOEraFglA/KyWTm94H4uTb37REN
IisAWuJtAsPwQfqP2r3BLHb1IKSd6+xZjS4YejGO9AsvmUfC6xUjobkRGEnohHdw3tP4gAaZNB0/
RCsCsSG+4qzq8TLuVM9PfFafcVE+v+FJPa/BF5gqI9D4oHBTmma/oadRPbCjICmgmQ88E6rwvi6X
5ULxhy2szC55TDGwUw/l4prmkwqOswiJ/r6L7ZC9ZQr3El53aExMa8ENxK9KwCgBEJRXLTVr14vz
jJZJMMbdN9J46X4h8BYtBgcCVaJmktiVYxR45YLOGptp7H0P/NGAoh2yqCD0o/uWRAiC1E5kAGoY
jEhtS0PgFyhyNawjGSLFplkn+wBm4SMt/MegfrqdpUhNZsxmiDvkmXSVO1+BXFGH1CMLDBdxMaBW
/dr2+jGD0sD4LnhhINbDrFEb9Zi2hgRk8syUg4GcNcdnAQex+Rj1rTjX5NhdMYSnraZUUeLRaSnI
Bfae2Myi/RaAbejMz1UVAlovcjEXRsF6MX1TtkRoRIBiINKuOL2tjcBZAmaMGzUVUB3pl8zRzTLv
iEFV4wBl9rfLA7Wu4jwE63rznxZ2+Nhvf6V6nP2l1Nrd06lB1zP3Hl2KJiqoBoqYJj82CPGxRfeI
IukhobDc3DF3j99HexOQz9YB76XAWj0jaCXvlSKVyt/zLe/DcB0y6jRpDCAlc+WCiV4ucAW5k70y
zqbwdXOc7Kmz6AAkACxoIqkZxHxID36qdbCJpqcwkTd1Ncyp90hnNR0defIX4DTvUfY1nThXgB26
YxadJYqrqNsQVb8kwBBSnKC5LsC1TLCesT1otobiq3fpzSKLVwyNnswxZIxHYjnwY+dGnEWk+OGV
zlcjrdFcU+BXvmis2HwdlvfKqWFjANT0w/O9QhEiciq2OhE630U4ZNRHvzmUX6hRwJNTAbmG8Vrn
lWuKCNpTbwLkFwhZwB5qel2+XLglSOlrtHUPFVhlj4nN/PuOjk2ezAN13+0fPHvg5DDBufNPyJmz
qtu1Fd7QqsE/OnNn2ABL90v4NjEpoMgfdOaNf2TtioBNPJNJDyK3hEj5AZEjz8ECO2DwxYmBSWfk
PE5s8FDrFvrAhjJLl7j0qB5ZNeKiXcdKWcAbZ120Rw905DJlPj8mGAzseyF528XE1ZHLHnzOkQuY
vX2dO4rq8SRdB5x3hDa4+ouwHuxVkTJ+ssRr+ck12S3OfK4zC9LadsxV/6KNBirWfAf+JM+pLGSN
DD3xQUqxLWlNl09YhIewlwORvaldSpy7pFD3SWILbKf+qjixwjM+Re3mMpP9AjX0HZ7R7tN/xSEk
ZlobcEEUIOd7gDlSrUpVUaNw1VJfDQ8qO3KWM5AhrUpwIGwcqirbsgk6Il1v8ewA3HQLLSU70iUQ
8uQLAlT8mc4I/NKrSKEd53hwqBBpm5zOQziwE/tYWMlr83K2BCMfgSqG0AY3ULIL/p5qLLTANup0
3vpoy0l8JqPtSbYC0Td8CeXU+Qro2bHzu4SKhaCp/2N/aw2mmWuwPBMW/KeSZjI84n+pvUjBoiQU
S2bzdXFc8GPLpmK+FssMOt051fNHZXujvKl4sqfPnDG/CEv4K17JXew/5aMaiFbVtOI6NjyGBu2T
csUKVQX9t35rKIe2o5jnzp+gJ+CQ3B21mUWV0pfc4yVvOPlMiFFVmZO/EeUXcm+JOwy1F4LQ2p4Q
ysYdenWlg/qUIMnxlAo65VCJZlkPGtBCkWbFcjckTMQTt3gznR8yahfbjXpp2bZp6X2H7F7xoeJX
pfsT7NHi9aF6CMAVFfRZm+QKi8ImNaViRFojezALgwHFfno2m4JSbSiLrkBAfFuth+yq3BavCE3f
bGKRgpqb7OpMYQxAnzuVhPGGO3Qpt2r8VucMpMOMrV3+VdQO6FljHAk+WtwH0rGX2DRAWyk86b7x
thZO+CQt6iUfRr5ZZT/ffUenvFbO8UlQI/fsMopjNzvfwGyjLyhMJzDqC31ounTh6+/Awq8V5yP7
EoUM/n5OWBwpKGtgA0NqdO3C1B5nwoczNOk5Xn8WFs0ePIdgrNgFR9Lv2tBc5XEZmOiT9PbCx0Ju
N8bbA00VafumVDEwrHP5WVUqYN/1t6p4TFOtYguHSSTLx8v1OebPYM4WL2VgTcfuoAIk/YDjByJx
ivC/3DFyX5agAS1qTIXHITtZ0cM+CZ0YvyCd1wBGrB9JMCIWlrAOKM2Mtpr7thOLH7YaFXYh0U+h
O99i76Oh2qjU3ZHmWCywUV4zt46iFudGSVYrUNhD/IXVb5MWYVDClazvb6e6rbVm/jx+7vKtex+D
ZPHhEUmS7LuZmnmkKhb+N3sRQcbGpesL/bEmlO4TPZyUOR+e9VFtTiVqKgJQWhIywatGkteaZGLm
blTluSAVUrOOrews6WPEOE0e0yQ6JVzEqRR442n+1BZf53Hb/0WBTLCffKi34ttznYO7parYGhdN
DViS1LUzXLPWLWies2A0Cy8V973Q+uc+FkKMs5lDDUz7RI92Oe1/v6au4v94WhPH4KAEUFnrpRgV
Jc7fwR6ryr9PIbQnZHor7S7px8q4XO7SOdkggR/kiWt5g6gZzx+0HchjdDggI3u8OCC/PxFMP0Te
K/2bJ/j1gVCURlxkZqHUBo4vh6ff2IBXy9w8Z+US+shtbnBb1JRoNAKx15a2E6YIFo/EXe+IooFx
GDqbYXH5ZTPocU4CsCmPu2KEHj6rVerEs4WIsyTvhiOk6KwomgQ+hp3exz3tfROsTceYxbB+X/m6
trfRCM1vGiVbtbTCfZPWjjzjBspknuAtb7jMd8tKuH2dF0//dTwU3CR1I076dAD0VNV9C2eQvrU5
IAEyq2FwyMltxsjlqC3g9Lcl349lBNscVx64xLHNxHjL9CFXNQWh7dlUht9HzBN/U0YNEJLzMjhl
/S2jvBZ6HxNE1wJzokirIqq/kD0oiuZGc9IFhqB3bdYtFfzpkmvekLXIOGJjLzXAE7P56qqIwo0p
wQ/hHmkDiyBYP17WpOcToC4rLnfC3hNWz6oBagiWhAAVJrCxfobIxL1B6F9SdsNYdA26kxzPCpxd
QKVxvVS5tJBCoeAbrSTPnDzljV2ecOck4CqenINmrE3WDNr8+sEXtC4fZjJAn6NRDx3MrAJCd5pp
z3V5uEckN2UZBdmYeR7uFmt0XV8nEOD86iOKnJs0Qfpa2/h5Mci5RTW7bEfif6XhshwhXYW0MCow
HLMD4HbWu+QeRxQnBnNFO4ugdk8ZF1zkmXXDKK+S2CN/ZoumUe+d86Uccu8Fl1hFaf3pNpxCyv+Q
w5KtYQBAyYsKFquAFfn3MM9Sa7U8947R5Cq6jhlLfkPA+DeEBfIUoBJO0sujdESnoYsRNX5oHSr1
Oms3VYKNKNccsqBLp8XTiRPOWfsZQdWr9tdWF+xUQy+fzAKNL1HEKSlNaAFYYvYBS6pa3Je4KXd3
IoN7Hf2xym3evZZuzMVZBvEzxT+CJoeH0UGEBU6vy+OHB7tkBvQ67cU82dgww/qS7Co1iX1IMA90
bFalNbNpViB+ZnIoP+wqwwWGJA09GnkoxEdhYEDOFf24ldqzuUpG4zz0JcqTeuKdGEP1Kq6ETZ76
n5zrDGPwd5eYgrHxXaYdDACQtk6UQHMbXNK5wSwlhTNYHfdJf5LgWiIhbusGUpBiBCLqbh0tI8JT
Nr0MPmBoQjWszwz1nTwtTxxsIuDcyCxEF5Jpm1dxjvbTT5m6c+Th2SjHA0WjRRvgAMcCkM/ooneQ
dT73b/1KscEOLRL7c+2jEnKEP4Zb/Ox3ZxyfON3Vv/z1IfYNksoFUtRIIPpKTdVQzZEWzjetE+nl
taoIDjU3Hwkcm/gXwVpaE4FIncvwwJ+qJNIcjaANHJJDujHoXC+XlGIHLO+7CabE0DFSbKNbubNv
Mklz1b8ENYEXhrEHLhEygjbnnK68EYK8Dglm+t6xKB9iNaHaTf4ceIJVMRPjmhsSejyCMhNBmAJ4
CuQFcWYEghP8fz+1T88FS8HxwIcrJzyQJiv7sv1EnWs9GKDDs9t9zrw1nkvzwF6CVARsLhUptY2y
ATvtQumfBWlZYq5QGxeaG+/pdwc271yWxc/Rkktrqew5w90RiFwvaOTrDhY72wNS5z7QPv8C8/WS
gSJBvqOraC4dKtogFb/KCxVg5glo2sSKSSLSAycEATZlovvHwZ+h3FJFQkFep85dAEzIY+s+Oo7D
uzkWnyfMCIgUw1XRNOLc2NUSYwSVv3vfKJV9a+CVkwJzTXz26Un8ewsTD/su2WWpza2KXzncHYbL
fSmGv6kPbfR99LqCVPGhuvt+7m/VFaOrKQlQ/ejxjdNOlxKossh1vcbYtflYaxmB4dbSQCkYb8IE
PGGhSBHXLqor/M4fzAyj/hqvsJJCI9eGAqyBryRaogVR5pBht7S6bs/VKVTOxhgfy0QhDtKNKoJw
TQ3Pep57uwkxZ4OR1mQ2QgbWYDpi9a3S7D3slcojmygM6YUX/YRpZyneHEOKyNXGWPY6RvAoLRfD
hTBG+mZvTkrSXWhG77dwGP4WV+oV3bmGDpTvOLvwt4g+2bZi8oTAeAN3m9G477Vf/MbM5RbvHQ1+
0/bg41l8lZPHeTnHOf+GeYTllvuCkr+L2PukgUIXpdJ0GqjocSG8rAsI1+2pEx8+hKbJaM7zv9Zh
0f99QEsQjjKlLEYAovsBf2si9CMfgz0hzOzXUjXfHPOfqzaANQ/hePPQziRJ++Yd4h9eeCYLsZl+
nbTLYn3TL86eT6kCuzXPxfpaBQW6YkcaZBRC2Pi+YCTiPfVzyrBvy9cLMdaeGR/nO/K8oA4fvT04
l6TWTWPsWYKt1yd6CLEWg3qCK0WQFtiX1b5M2xs6/uRj6/VouuzgvpCLb5Zn7i6wRjf1NtFG4O2f
JhbsWZw/L03cbfq4iUZ/nAV9qYE1fQuRow5uuhl/km3LoNq7jgaJJCHcHIA2Uebmz0TjOuNqQOo+
tYNEtSQ5toQ7tMDPvinMCbTUhXH4tZB31w4aH4n+i3jL9EYj57bBXzGwll4hLxIoxYOE0SgGi6cU
LHvXC2MJ8zKofjDhiMfllmI2f8OBj9Gu4DCOscYlAGFo6CcYcB4LFnm9uliuVCIYApHKos8fLuxH
tx+xobIj23k2UvOnUSZx3BhBB8ahlN5LEJdmHcsjwdV5pz8YJytF1Bdk7nbt7xBXqmV2cjL4Zgku
9QDGyRD4msTVwL8zHC7bc96qEk+vjdzHu9f4J97t5hznsAsDLjtWn4iwSQP8K2kgk5WOW5cAlTVa
Uc1R2xzKTJZDUIabzPML8W2fVB6TzHtcFcvSL9ozwoKjq1H1HXusJauoGDra0cDh3TwcEeWuIzXa
ciPeepYxR8Wc4ntegwpARcueKboGIxz6Pt0bTmg/PTUz/XDvPiWDmhxz2aM4PlPBg6VuSCq7osgm
w7xUTNVSswkxMYB12swUWy9bXMD0kBI3tSJ+JScUnneIppGrMBVDoT9IhcPQVNMd2Qk2eKUQ3dFM
WCYM88pXIy8xldfmgtB3y373oBfTcc2xtAjdI91MFvQN0dhpRuVFgTcG3fNVyn4RQmxuBnO3Qwr3
P6+Es2ymJCoOy7wD+MewOUGdzRHijfQiXFaVtsFnUse5gBhiYhgdouzleK7RtBWZV26JLAYhopTg
7uumoLT0x+muLpCnIWiGsPWGXgkbF5KiQ+nSAq8dpENLJWPvxWZz/EujGqLMkz04FnoB+UcGPhNY
gzPIhmGWDy9QZORzFwqUro5QLNZlJVfzmecyEDCO8lYFKx3hbBa8/zfFt3X3fWF4S3KEk/3IG6kZ
7xnHQWXcXDpuqyRa7PhZ92PB5NTOoRSUDzaGTiULBiyWsYc8oF8gAt+y+jlVl87E8SRvLoiAcXo0
qxdYeEY4PdDkfLHC9PgKY4tSk5OeYE7YAQCS0zvPaEDbNwHHyi/9MLUBU1gOODFUbaTpPVcMaYdD
IBKEdT6i3WVBdELKZho1G0yBKkDru1rVVP1LA7kwUZ0gssUwIc7F+bYe437GLZcYTpVZMlVYxupx
6sKY02QKMkReXl1/incBsPJCAswrefmTFr919J9M6iFEr3wrc0W23DRvX09Zm3fwIyhPfZgTtsuY
KNOfoil87ZS8ZvKn+lMi6bjnpRtBn+ocSEk9UtzDXVnV2anb033Hxtv+sFE3rQkC+gSzDYpotPdX
NwtGNTJOG83+D/i2zg1TLdko9qebHcVi+Lo2f6cRqCIs95kn6uQdSrb/ZLuwTipg/QEslYN0HVH2
7dsihC6ZXz/Ren1oWPj51xHbbRafUGrwwJVTDS4rrW+sj2/DvYP5weVnXKquvyyzBnczv7xew0So
0suCsdqcAc3HHtnwEm9U200LPK58Eoqk1Rqd4QqcOvxmhN28zrImb0LtFd4pGGI+mvgi2HIg+EKq
jITLeVnmzmuU9QtrrM1h1Fi8NhtH2QCspwUMMXYVUTZamVexhi1//UFNCZGJWp53o1D0hbqURTwd
paSDPrI70oMSXw2Hb10Gc8UJKJtg/C+UNdIVdU2MsyPXx+WO/hDtb6X+RGFrGnggqNtIaBZ14OAw
MGSZ2we0Rafe6RRVGNT4R99fpCqt4U/TOw+HgQfORIjyG77clHcgt556MW+GZbis71EqAe872Lxj
citcpeRNL2h/2MgQ12vUqftJLADmHekcdPmj6134BNmsAxOsSYt/FMcyvd6jU6mUVqUGDRVmVy97
dPOoRSM0e2hNbJS0VoY59vkOxQR7YFY651YKgdxLoOQMnNpCY6EC97OEo/dVN92BJ1AhWmuVjxZ0
m8pHYaviiFt3u8RpsuV4PjpCxnA234FdeU/NEWolNl1Gd1jXQXlEnvgf8PXvS8/bVZZlg8jRYQvX
Skmix0GLFP3+wa4/ZWq93AzCCwNrcr0cRjTREZcyLf3PTCyYQaeE4bbUR/bzCtJfQnrmlmbVZPt7
G+/FENgmyWb04uchkSNoeyrYvV6j4I+UwkXezHlKgYc67SGwyc39yZgwdeaL7pqyeNUSBBSWznmI
HEEw/IYM+gi/icnZ+S4rL55RvKi2l7ZtWC+QUuSyWR/Z3ydzGUktC2liNE0X5NO3kW6Zu2+OmfpA
VOCU6C+TfuIOwcT5x6MwMXzqHgRbqBc24nBjkHZTLiSbF357lYIogT5EEo5hhPTP/DqAdrcvPkdy
wWvqDGi8Nape/3y8SaI1UVetWavPYFtuHq9boXSMMYksZN3Z+1lqSIhiqR1qXJF/oqwl62RZRrs7
PoNkjMWU0y6x+hC29LyEEEs7u9N8cXS4Q+NOl8ew7i8o3I4n1IfQgzEE8muEIv2eecKhQT1qeIq8
mq4nK40kr1nhq/xL2fTAIshOUgFlsro9HP5WkQRhEM459AmOgujqq6G9lWNXRAhLwb9K/zPVusRl
ohxW8rPcbFgTLEiF6VkyaFqbm3YIj8sTx9lzyxGOdGGpLRZteHdFdzk70skDcKXmW9xfzNiiL5HP
nzk0CeHl0llAcaDzf7Dlr6U5MsJEgt2AyAv6Le9n/W5uTiRrkT4q5j7F1oLCQ6KzRhqYaJvO95TJ
tw0bLFGoOCJQNxDqmBWcAzCUW4EcKtJCYYrZESVqaNUpW3A7yEuhlkkHY3SenSRiS2vRu6Y4YPeL
ukrYQElNRq5UpvU/d8X+nLmJhVZK5GQB2df6B7OGAp0F0YCP6ImZ7fCriZCTxbr8Nux4mqiiIta9
Sr1j1+lVKC68gf+R8VpgEZFTypwTXMJl8FcfPm7T3YarqxZrU9Sm/fmoYwWEmdG/dXqNGH9BT0px
RSX7Fo7cbtS6qlAt7s6ZVF0PvieeNXQYJIPym3P9xfXXLX9laQPBwluLSdJzH2tCu8FkX/FfUqYj
9Efr5Tr2d6IjQY7J7JahrfvhW81AfSZaWVAelrvgVLkO0hfdyKmynjTGJeaZW7ZiA8d7eRF2rIxn
YGYK64GSS2qVSjCm+CKxPMsi+zrUToND9epOo7JCjqbS1sZUxyf8jgHUsx/zfayOp5YUF+LBKWPm
YUnAptJCY5DOD2afnGFRDWRTnC5wZlzPAMAlNRbsNH+bt2xPlXwx1uaFb+oJeVe1zTlbro+E0d7T
DNHJ4/D+p3FczprLzk8VfmvWnQgFROJIZ6UtEgpeca20JxexwFLRMZWNhxUd6QxzZpNBuZGptz+A
cIaiNycSJo/Xi3QVOJmYdmxNVpAZ5sGoTtrxXl/qvOW53mkiaf/0CRVmZngL+KKeLng9CpMh8nF7
30s/RLsFqwrqRR36r1NPG5AvzwM4+DXHCNgJ8bCsDnQUqvl1WCs2Vsz+e/yimrFvall2GMIeR9i5
b1CVf/TvUFHmDO9ehqO5FmbG7lNmki/dpdYkO5LH9sh8SNpI4udO0eJhCN06PdPHMqv08zoKYDOu
FjQE2Ja/DCx7ciLSCfOYMBbG/1jv+8TsdXkbHYGErD29SIPr+dJpKs84Act75gpMx10FIbog2bVj
LOD+dkqRfT4oZNNzHJDrBXDux3/YFQ36VSJEkv4Bi3eJaOrmHweo7oRlSkEM6X0UJmlodJNVtj3x
hzV1tz632eMRr5THfmUgSa8CmaCmUKDgBui4iQ09FT69lOSwFlZV+Y1mgDenCV8pAlxEjTb2Arpp
iit0VD0i3qohD6FZfKBtAoCqlTHw+g/nf40ipwCgHy2BWC+uMCqpS00uzsKMJd4Xocb3zW+Tfi4S
2569yUBz0GV0uTlpJO8zzPcpuXM+Xd13cUkLWRiagnewVIzIY+KAJIn6rNmL0Co8P3p4Zj1nw0e1
O9wZX0QtCR7gQGSg3dVJVqdgPTHvG5IOHvReMIZfXp0kVDGFHrD2xVUaoyGieyPRo5+CwW/BMIWK
zeWNb0YW/UVBmLK0DkELyHNCeAkybaOlD5ghOl2E/CBQYmbk3KcCvI8+HuS5vKiSQb/yLYgWg9/6
mB4o91HnDfWMtHf6/EmBDrwhNT1qpWv4ztIwJgD3P3rthzwNO3GqId19E20xBEEDhyWPMel5/m5i
+ivO1Un+VvW/7Dl1hCOwesx+HOthbcU0f5VLDW6sasXeu/9qnPbGqmIq4tRPs4t+fkhtyEds1ZRz
hu+13SN1toNSdhxMaZazPWBr/NBAch1mNfzkw+5H93dEjLEgD19ej3N2NUmxKTF60GFlsx4U3Zji
VbLQ0CyFESYDqhgWI328K+Eje17HJdkBpVUP4imcyvz3rGEIZ025xkS3AvuZuxGbT8UH6swTdXMd
jJhc0YzQkyIuyWW/lxRamWnQ90ki6UVWfaMR1IuxzRDcpXqqcG7irNklye0B1KlWNpRm2Vc3W2te
FO+PyiMaised8OWwtVdaiMeStP5Cey+/fRwPsLOTjlDKjwCw6EUa0afrxCRpkEXVdUVrOGokw9OH
c7Fm8GS/aFqZLOBFmzMPRgMFOWbrSyopg+jFJfVqtR17oHxCgT1DBq2ml6qCH+Fh6ASAzxgdKswO
4yw6xehR9D1LxU4p7xjl8EdQlWIMaJWJ0ZArthM5b6aaQXIxyYabw+YIE8G9asW4QzWAHcpiE5Tw
/n4O4UdLtLu0bJ2jbvod0501mpv/hs+/Jof8e4nT1YQp6g1/kBGtszPqjthGhiMH1nCpjGFyElB9
w5VMZcNZAzwSUz16qMDkr9VJI9j7NBPQw2BZRA+Dw9oVJ9Rp1vQfFVaXu206+q7HYFGbpt/41pfC
fpPyAIOijwHyNvXqFs04VyAmIEUwNFOrfsr7vmUd3vgk4kfu+eHbjfczesnuRJuE/EBDvifGUPc4
7cIkhL3svJaBnKuiMX1S2RGoAanGDTjNYk/LlCKzgW7iybiRU648zl7bAKTlnXnQ/ppgMjgmIoQC
NjkTmbMJxcf75gm5oq4YyrAO65PLHO+IMwCPKmgtEbG1Bdv0m/iXF82ttF+EIsZFe7GD9tYbAdgu
50OxRGVN+rFHX6VRPaW2mo8iRnuB8c2YtBxmflpngFxBeYReKd9nDKWXHXTH+HY51w27ndqR8q6L
bpcHIiBzdCaVM6Hi0B3mNyxECDKURfEJekcufSpv1s3ACJO2tB6UNGdbGuybCBcyUWLzDUoh35r4
+FYgMJBkQuFOaQvpdTWGTvNoxqdwqzRqqQXmQFznYZhyGoz6031Xjo7Go9keGU/HhddxcIBf9zfr
Nr3Kk6Vl4GQ0Bi7KKVPCAnT5upCOciXalBA0JP/jSix264evZraymR9THowrNf/Ke5bid/vVZC8z
UdezQ3uG1KRAsZM0jlTs7iNNetWO0lhrI1VTasDImfLwnH8E++kMxxsslRIEZtVKTBl5vY0yfuIx
HgZ8JZK/czE4ZcLAVDCZLBP2LueXJcNuOeqkODDPCPXZIBmfkWkIrlmqO7qIkY+ASa0Ll1cePZi3
5o+g300ogkEOBpgjhSbbX39Lcmgzm73yPhavcLPtGViCKwPDp3gyqQi6gMoIapCm2mqqL4JeZC3l
uMvky2nhK8FigGmcDkl/nhCnAO+o+ue6v1W8YVv6BQi1mxRH/TWzO07ZxMkPmy8bzRLTxzAQUPFm
IsR5ILxJVvci8p4PqS1W9G5jq2+4jeIjH7wQx1DClj7Jsv2FWM/ReI1XTPflg7EeWnL+/CFj9zjO
52/LFwWuJMTMbCSY8tTttQn1vHE3p8uL8kmy6ff+CA7A5YVHh8sSu4HZGyjMNTEzmdO1YpEj4m73
5HdoemUoCW8QIPXWVUA89jj/vJwnRCzm8i10GRdGsYjBH0p/qWStEKfvNeVOQbAPTv2TM06N/YQ5
GbjGgYGEa9HyX0+XfB9AHaK67SF3u8+CrCfTTEmf95MiUJPPrIlFtczPLUvPfn6PWps7/HxphQVO
deSYnMDMAvNop+1zk+1HQYyCplrBl7YbQY3TH06uuzvNoFf/6js9cVg399wy5K7IHua9hGGxCaFy
2jd3MpBkw4dHPzqi/B6KakTaMnC7R4lvxzbzaSE+aIgoZdXG056G/0euENCQziNyLiwNr/WD8Jm8
O7fn+OAVCD9BmpuN/M5X/xR7GkY+3z8NQF6CI6Z+5W6areme3FT8iPcTy21agfcuzKjkjekGx6x0
wsMhYnLlwl6k/C+zXvKXMaRv4KxxNDdkbzORz6/avCkTCZOssEb230HEgLwXBXjYu44+8h8HijNf
LzXTMSpWXBXcj9zVBpjNa7iwInwQNKom3ldn6tQCK4IVKAjmYqshnspfkeQi6CirPpMqzY8QRvsd
9huxMoEh8db+MnzZZyTVsF800hG7Tr7aLtyf93zzYFzD6i23NCo1G3+weJ3goB0qjKsv9Hj12IGc
StxHG4hFpg3c1i4lkYMvm52Y79m1mQEKiQgt2+JOsgnArcckk5dXeZBQbwWDZaONWFcNmPZZ4pkH
FxKri6Ti/ogs9ij5PJFN7Bx7dzio72wXz+0qUTJfobZLTHV3xOe6k7BAtL/vpuBfnldcljnz+Zmg
RbFdvos1tu546TmCL5QRz6GjnX9LiNZnSQF8BNwfqUDU02mal9g5JFKo3W/og371fdv2E8Y6s9oJ
VBJa3SRW+wtxGQDGXTRjW8BcOb43KZYtfgkyxIEEVumhVfl8gXcknW8cufR2hHNKVmT9G2cdBr6d
HClkPKmsmYRzgP45sOFsYv5f5ptmjWjLlzeqHRrLxUedBIufDqcr4i/qXk5zER4zpTsDj9fZG1v2
CxP6jDYY/7zI9MTVcIo3Hfbt6Q324KNNlvua7I1+2r3EpQ+SsJXMILHY5s4QThJUKFmouvPz+s5p
1sOXV6aREsBkPPabtvNxDlJkiiCJlOftx4Zu9S8OyWIRFUmwp4/kebfsUUGGiSFboKLlbJSAzzpR
clbxzY/tAzv7Lb7hZdstiDLXp0tsh5ddIHEvLHBi70orZ2GpigG5Fg07d2DCZo6lBlJKWDCRD1U8
juPCtfiArzmsaymPcaXY8s1//Cotw9YHm9j+j3hCv/MLIBgOdMjphWuH1QCNFJH2HytFQJ2Q4jro
3Kq7OT99tAB0OU3oDwyI2g5H1sE6Wg4BDGAS2+3CmJZResWezh++hglBLLRrij2eQwvHnnh34H4t
VfiLPK/mGSL/37ynfBz2zVHdIwIVqXufjtO6vdSOw39bk23hQZM6EVwo5uWw8rq+Ee4X5+8m9ovP
K1o2UFnPXoCyPFLjYqihoiZhDR2Ws0s+Co3fKClxDgrRE6cIiNNN/1cVN4jyzWPnoaFBcJyE/s9z
W/ytulJyo+45ZkBeY7EutmGo0+LhHUGqchHkR2qw7cHt1OIECzthuUBDCO+l8J/m3tCnuT7Ohc6f
JxjIPQNu/r3ztjBgjIyxLcaSWI8Qy3jCAaWRsoK4Dot3DxdXu454ZMAP1UuG6930AEMjP+c73QA1
6dkjzIsThTcFlSbCkOM0g7DthjkGCgiU14opAAbwd0TLqi6xfswyxEKUig8IT06MLIQNm8RWYwXb
kXrBg11KtAVqg2cSfBjhiOSm+yWfEkQ06ypiedCN7rIgM8Y+PRDTOfgpvc2J5RtK6t2A4SKkgaV5
UziAkBUqR2zlc5U9PSiMq85PNMl5sArvpc4je7ZqjUN34IPQKw0GtyrARVZF6LGDgvffRbrQcy0Z
eMr2OLJn61zYjJo3CB93A4q0t49/TGCwL6oCCOweenA0I8JGE2WpDvUht///zpGCgFdYjpIM4uAq
zD72uLPM1mnlRCSu7tJPtean+zSUwczsxtkX9sBeZT8StkZxkbnedO2HCY0eXt9/yVXi6lCP6qNs
S3aqoHIaYODxLJ3euLDDpEzpm0BslDZQHuAy40KluHBL9g+15jfFHVF5DbkUb8lsjpPgFY5b9Rmi
ONrKOEjdknc9mPf6Y5miqgtua5pi29CVT/rKyBy/EHpTeIepbZu3InitvWIo7NpJszruTbiI0/+V
gUrOxxkdaN36CNWJzc4NyyHuUW3RbUdcbIYQlmZgoPxGUE+7qLwOlrhRPx8o6lgtfSGfysORt+6E
rtzexm9EEmzzSpy97nniLPn7ebl6/r8ANfuiNxuzB6PbAmvA5Rpa8ZjEaEJEZcb+7byQzGBadHBP
xRb67682216+ToI6o1vAH57x/IfWmop8tFU4hALi1sfSjGjjt537jPYD1mV+U11rNj/INYAlnAm3
3ZdWjlhklYvTbhzAfU3X41U+oK0C/FgtBss0/TooH4n5U48rHi6JPWne0xehK/SOetnk99tPskOC
FkqECkRszjTemLQ5RiQK01NCTNwQUEwqHJHW3Qy+sxkuYQc+hRLJtgnldUYfqAtMdIE1KFdFC6mC
XafkO/K4WuPuL+7An0W2PhbpVNu+62eYQXc+EK9t3krHBC7YdaSDIA3jcXg25Lg0Q0yLC+Bn2AM5
/fKMIyKfM/UNOIYuCvvLjWTIK1KoxKlE5SZLyhyz6ZvUz2C3l+jdb6jcj8DInkG2CEF/rX8tHcWh
xtxFAiLCBaM3cOV05qhdOhM/T5P2QYayMqDlbIVJvrgrXoUlAHODRDGn3Xu+yjalA/mCMyS4B0fq
pDVbxbUIJlGO3GPQ8R5T8sGx4lv0AMwaQMboID9wV+9rU/L1LM5AlFI3I5/O1l8KzgM0ZGVB5JWh
LHHdGmibjr3e9DgcopyFh0imavZ4STn2O884EkO3NbVZmsvZ9u8Nu0TNCAmmGlpMAAiCylGyzkS6
0pxmxnFXh4dJx3O4Ozg4Z9NLFUsz8TAd5OhMpH4IFtB2RynaoitGinzOwB9ljx8S7PwftPzaGpsL
uu56Y9tj686RqSYsl8COrs1KJeoPAFFu3ZEUvTZC1k1HJxvt14weAEga9hSo/7HRA0Awn5KbfEob
zJKYSAT9GFCeKjhQUS4Wju6B7YnqT4efhvK5iEm1x0DeVXHWTez+Hfe44Mvnke2jUDqe63/nR/Zw
LBzfQOc8RDKtpwklBQg2Dt3fxShEPWDw9uoOnsRm2yW/mFi58S8zVzWbbjhH+ghK1KYXqDIt1iMv
iR1AgKspqeVZC0BoeVM7/pZ3/2kQfPKHjuHg3yohQTAfae87s6SSCP2cftAaLmd7uv52SK6Wj2k0
fyZ9kmORk7/yOGPYjOnZRO1eAN+BpWnnSmb3Kbfp8itSfaaWdAkyoJBpruT1BGktPFBcpxWGXL65
c2cvLfUyBR5DuFYwMjNKJ7Z6OBD/V5KCindoOEKzsZoZeyKcj+W3yuieFKnWr40jKMOGJPJz2CWP
GbnknmY9RdcCL9uMBumnXmcTQPU3yMkZlZfSTfvZPkbxU4FJFwRzCq2tIphybdnL8nBxytIsfsGG
PZW/mt3mapA1AXfovIXSh0QVjsUzpb8jknu36wUcVfrHdUuVNpuhgQCfeH5K7OMaJUtQfKTKndSt
3T5L/Cp2yr8skQyiSKRlkteXHmsSonojmMuFj/rwCWc67QzSOBri0+iRA+S86nBtUD9xH8qcIbEX
/U6zV9ixJMsptVN4XipMqWJYh+AowszBjxFJ5uP5mIfVQ/h104iXmY+fSb33dRoq0DQKryNaM1li
nK7KB/Cua8zV00X1slL7XXyNupc/G8zihZ+1jHH2idqLSnKwT7aoLVAyKFGxBSBtjRYxrV+QeSqX
MBWxqpddQsYelyH9ODKt8BxuGJBddmy/kwuKF4VamEan+IWkhUYnp7ue2V34ca2OgqexP7h68t7M
aDM3VdADaH/cJP9g9KSN+eJJZ9vqZOMQIqyr2ug56cXiVXjjHHVtUIPiI/rl9I+WtkF5EVTcnoc1
RD4ez3wuAEvG9SSztm5S0BXndVB/NRnwpeElR9PXWMI/WA8AwrzUPbklr/9fz1E8f1MlTTKZGv+Y
ycxFOn/jXqFkoS+1RJc17LoKuExU5nonATtsnJl29uWfmE4xOPbsQIPAFS2TcX1MIMaS/deI0D55
3udqBKGJL6qEjqWnU70ZttY2IXD/BDGr7wOtVbpSwh8Q4UzEUeaUwZEAnyTVBUFEJlKtJWomcDBy
CTt+wcAzejbDEN4/FqpVScR9aU2fQYN6S4Kvoh/31KyQEb/h38wIbdSYze3Z3yq1tyWTdEEJTbJ8
lPQENruIW0px2hsmO4x9As/wP26if6G/IY4oW9kkC+vmAp2/hKCRlhvEHfKjGQAlbDHUJyFlA4jP
Xs09tm+tBGjOxbsYY48BgvMAnvudy3zw2e+2x3EWviVwuaVnPlXyNPbHChmaVeaRmBsw+PAfXUzA
RHYOjQJ0bf6BZUY2sWlt+AZbIOIU8nqgXzzBrCQ+k4Z5SA30uYa/x2DMxnHTPzqIeHlkJ2+4bOOI
UPcwem0mkJIVLQKmPJg/+PCBgaYXQvTSlfQ9pbQu0cUOCdCgEIkCeP6fhiQPZtisr2XGjC8qdl1Z
kn5obwrtGavwvU5xe9yC+FiQx7twbdGRWJM2nkP0LVUtPvVFbh4J8JrRw3Qxpx6qpiBLdPeMf8l/
GGhuCrbClyuhzQ/7fCZlMUbhIxivfZDHANymXWxJqvKQ4RJhW3pI+Dm+TCCmr47PZyq6VeonRbom
wpJJKI1pDIA7dOiEWGD5LvQ5iq3hmnG85rkYTH6ZTingvj+8YP8+g2LafeDNydQsK7IgKk+sCObQ
tEOC8PCzXynl290FcGGDfKhy63Mzp7gBDkAjtahzBd/qfvuf79aS5SN5tbg70f1JEIuzTnCc2EhG
g090w+SJnBvlacn02bN9n8lvpcB1nWIYjm5OM9y4h7oC6dL6WjEu3Ox90LB1WVPtZHHY/ahsyEgn
SO+6UuDIPyVP3PaUVtYPt+HQFAiWkwRqq8S1Ir29Tc8CkbGaODrcv99ib0q9jU/bYboSC74JB8jo
1X0w9kyzufEZx70ds7koQAhHO+ZJ7YRjyvhKRSjnY11DlrVng3lVtBgGFliblSIOeCEw18a1zRGN
cDAIL13JcFvFNXa1mSEAMCqGr1CzhLARcYC/V+mEjah/fgswC7nKQLyUuooCL9EsxF3kNE2/i5EV
qiW4Me8iZIm3TNXqKblWxgmRzfVYJ/Igk+0Yp5ddjlP0zGL8jyUNmlyHJRELiiHqc+WIaxIXeKDK
32/zTb8SI/zzRJQamuWKVIjRHfjjq9Ag+ohU+XU7QPwVA0TGho2WDbu0ji4Ciez/V+2UN+hExjtr
oxXVpj/YqTabCLDArY+QyGUZncgJ/P4NjIO+T0cMdIfx246Kj/sw6Oq+XPsC47k6lLe/ArToh/an
RS1b8URfhbrA4aYyiHwYMXh2yVvL2OIwUVY9i8y5PHmKQYxiBqp8iXy7tIlEj4SDQit89c+09DRD
/aZwJK/YPu8e6u67uW5mqTcvz1e/o/fWgtlceAeOs5LUJkkUI9aPF2mFq+mvF1Tkgew6J1oqYlzM
18XqxwObFH7WZmexzCxkZiE/+D+yjUoWR9Hf4UVAouKXMUFEz2gJ4ZS5KCo4UgGFWFeRQMitYqM+
qcTHgOdKRBYkSuXlDuAgco9WnAicYYZTlMGqc7UczO+u7paFW25MfjlyoC3jziy7aMVQ1DBD4ClP
PhUX8sN8U54XZnuvfEZoixy5UdAYWnVpnREX3Dxx3ur9vMNRtmTmvdO+bNXkeThbnJlDSKT3NMiN
/4TbjXf1GjAJi7DGobJWV5xmFJ3v+YjxKWWAkD7KDxMpcwrCIvbMY4mIvw9GTMDTMl0uo4sYbjad
iRp/sjOv7bvz9LOHd2UsslY4zcgssHeDcPTJMcy4K1VmKe8ysza+6aFyCVg1E3NVFn//Pi4K+eJi
1YkRbCxWem9vbG6fcXIir3gMsjz0+g5c0VLa+Or0UbhHqs1O7wfXfDKI1sYqWbZjNTSqxyC/Obt+
21yep1bWmCTM9I1r5PQaAYN8souh5FC94RraBCjZPRDinNZOG5gAu3afbICEa2KejSaWsS7sSGP6
YOUBzFIp0YwUPk9jIpXafv+6ukBdswdU7t6AktP6snImzL6J8+jg1sEqW8/Sr6Ae8RwIO9BAN2Sa
oPuf7K6B5Wu1uX/TjJoRimoOn4GMnHIPrblbhc3YiHr0RXUA3FM4IMGuLlOSOxs09pM9ogmCiRvv
X7BEXBTzOuu+TqYvHQ4XpWhS7PfQ5E/UGdu+bhE28By/H52EP3YQcsAGo8vvV694bUU1ENHUCnHL
va4yNVk3USOf71MPAP5y+vQlRyUO/MZ5Ik5x2gMoaQO123o2pmwa+9b8T/2tBExKCjRKnpNm1E8/
UHWA9n7H39IE63lVKxsZtSUkMke800J5QTXKBCkJkzOWLRpdh0NJlQUpYz9lp/TLgeLBxzglh56e
1R+4zFJJwWTmKm03uwOAcDXU7C8YpnPoZkf5+eKgevCEAMe7Ul8dvebae93VExdb6CqKdgcq0qnu
EY6xqlQfqY1gNSxMa7Bb4fbojhjzL6mcjyvxexT0rRpBvC4VvmM9m6dWycJS8qPkfWL7aTWF1TA4
BOHKauyey5fNEf4i9URFbugoIxm/3DZ9nWPPxNGMwykCXzldrlq0ZyzYuiQssmYm1lYLc31rwN67
zFfJDuN/1rjUiJMHP8Q6Cxpb7V3SwkKUiMvLXXfYyM3HzEOYfZSUjW6inFsPAVeCyG9u2ePBjneG
2bxVUd70j8CC6SI4vMZVb19AFiy0zNTpnurFObXkoqp9xytHGU2WSwWh+8lsBfWYu9H4G1ua1UE3
0IwPqGy6f8WdAM96/OlEBKmdmkRbpP0fiWrrkOJyC3du5Y2lxiw8H2SZaAwEaTTF6txKzIY5i2ql
PSonWqPefrUtYo6Z+qlCsIjkZaNGtt56w+Xctc1IiSQ4X8lT9eC0yFZb+yHLGQ+hJ7/lMP6iYAQ9
ZHG/IrXPTy2xKv/A5vME+u2ER5MWFnwK2uCn0Q9/yq2whlCrv1T2+kDXkzKamYaGtdKKpdYekvYF
5nnbf7x0EiqVEZmzSHGl8NbFTwfOM17VSWDbJFKJ4dSIGoq/Q24FlPa4ynsH1e50tsBl4iUPkBEf
P/Y7mEnn8CU92yrGAmLmYthz9LySwS5GKlGicUeF6f4Lfq/Oyvk7ZnQC0bYe/U96BkbCUtJwGCwL
EXgf2XNwQN/LTr5oXsrnwTU6u/5snPZ98lcRIr2sgZGMoV2lsqObIMDrKB4nKcwjHZ5waJ+7kyIC
u3oR1smc7dZvD1a5BoNHSTQSdE6O4zJ003+TukVMZXv0N7DymIvLJSM9gsjkWis33gjDsrI9lV+l
MuPbJXYq8xGp6LYmR0tDMUbTpRnAxfgCRikcm1R8jARcw9kixcPkGuKltO9yUd52cpT2q78HV5wn
n4wSk6LHKQL+W77PG+OMYoGDXIb9EZPfYapEmZ9bR6o36dJY7fa5imgMPFZum82B9P73sG/SUeLG
xCwX2Mq/y8fxXvc8AifavhD6m7nSShw4Q6IiUsQ5hcaKLSdg0IWKyJBptFO8luEMaZNObbCWWHYK
puGQ05KhAI6z9y82tsMu6nWngLCMoov1W+iQyppDZdeWFiJmTeRBgbuxt9bAnTvgmc3DrqYK0XuQ
ROVSeMMY9ttmMTp0a3kzeQJzoydXGHFjfjjMDeflw2yB/nEg8tNVD2YtBqryD++16X/S+Xjb0ZeM
Md+ClflqNelNop7nIgy8FMnM5vqZOa2TNZQaoSuxOGc1OMfoshqzmOqhcJ4NamOBPPMo85qTgL9/
ZevuJ1WsMr0t3Uec+zlFL5kvWNZ6tDhW5AgdlKoL5rH9G0RMEpL1hAEW1goq57Bo/OO+2sevLj5m
85zHAeS9xdDhdQ37Pp8LrUCqsPvOLadap6rzpoAmWLqBuGSAtjswRBLS73Tbc5b/vNVu5efWhQTc
GqzWiv7hHHLt9UE8kwxOsLxuz3BBHJBvi2G/cJcwhavzijKMI5qKJUsxDwiq3ecSIU69ctjl3G4G
j2WlAx57qHq+oIgUuDF4qu8rFMlJdIkC5GYR6tlM5KOJcIiokxM72J7Al9td49Rpq3GGrVTztk9x
X4YNGzzFUeLhy2UdrABEQZeKqpNDTFqzXrAyyp/zD7z/yq5McK3mnSsXtvwpkliaDUiAHDuhrHbf
RvVRqSCz3mhi7a6HIQP4BuzO1RX7WWmo+3JhQQx2SY3VZX1PxKQ9CSo57O0RlFk4vGWk3jxbjt3O
snORlUjf0sETzLal+xbS+mberi2nvprQhyh861LfZHrx2NIXT+td9Fc6x8PTeG7vNmD6OrRUxcUF
Ogp8FEuFduQtoZqpG3DS/nK5g8HO1kJGB44OHIaRN8v9PX9qo4zRImk0I6c8avijOtysHfMoixHO
gjv0GC0v5+bBbTKhATyFaJycKkpT2WRiRwh+hmIkEWsUcmJyDzTR15vKLPmNINJtMKl3zDyUVzg4
GK8ZBXq4e5I8CBzgHv0TNkgRraaWhfgDDc/8W/qbwLUwYdcBivIr/T+JZswFjrLBaFE3Jls+DG70
6nMYSmGKMqwL/qeenngoMlW/iGTZNapTcLfSoCHSJH6HaokKYaV742yJ4hZnyKbXXhG6YoYwH1C+
MwygZVZwlLeBIpu4x4xCsx27YMVfx1ON2QGUdRfCkGqXlT5xZ4AcNTRt2TVDbYSbpCwheUgb2ynq
BaIDP/C19vd7AoePok57Wv6sqH/FkDzAder3rlrEE+PLsGSCyCdi/yez/OVa1XdlujqCtocXObrj
hVi0kDdgdcFCxk+DvzOMl8a/pto8K2FSZgXy4oS5UVWUAZNeUcT4UMc3ItWpt6hF/vueK1I4Bdx9
NtAtBVpDtrswDphJwSOp+YHRUlAdBvOBXBF8hBTruTeKbyjmWV3c60w2Ap4EJkcdGs8RaSeMd8Ob
Xqf02jPWGn5sgAlHdYWGb2vHAslGrz1RVyeU6h4YStyYwZhRiMMDsHXPh1wLA/W2zwVJwye54S35
9pzixuJx5e60zYAmf6W5ZNbyF1cAZQXm4bRO35VgZodT3b/5vOiXmUMe5EFNA3fOIvdketi+30r5
EZMhA9agRWzBb8+DJFKk71UchskPDdnBwGU2HfnWgA9Q19FjthR6L7kM+AXa80mBHnAimVuS8Qpn
GAzJfEoGOkj8WSCqUzMRIiUr4+Dd3U2myejrRoMzdPsyEQloiOlyIQ7nrsaGOgftcsbIkuZ91TGE
GYpIZLt92PpUskc6hVluoXmIq5sSw9Sa6udSdoNWhdL69V/lUjNmq4wRp6MaCdsYCoMyb9LMmJu1
WqfeodDeQ9/LdQkr2I72JPGyLrp9g7y6YQCarEdyo8iPowFv2wgY5E+VwwSHqUzHjhUIySNK2Pht
q5YZ2r4N3wThKBO+Fi0pAtAUb4DsmOe6wm/lUxbHzWfVz6FpO6NKRBlPB+EF+DbNuRRd9JR/Y53t
zBmvVVswfAEykB5lHX506+CmP5EmiFRwkxb1XSkfldTrx25SEiPE3bi9DkPNnIp2l6NVJhqmc44G
Hwdqe0NbHVEhDmi+XFZwfQPbC1tsA6327519HjMphxsPYrrHF7X54hANnMAqmka4oVVSyP7nfpcs
OK79kJeT1lBH6I4muEV897rWVgLT/U0rN71aWrINZP5fVy4WQFOjfQrqY7ciUXJaY56RcXHEejWY
A3xKPCO1RRKtIGw+5+JBditiEOVoUC5YeeQkP94aqjB03HzB0dT6Wg5ksR6z+xqfEyHPt3CjblO0
Nvq4a2OFAFudqzVcdAu48C0CXvqCVTc5PBOuHku9kauzXR2mmIrnDUMgrF6vUMu5/WmWGY8KZLZx
j0xKfpUpSYIngDrwxZ5dcoNRayh8iAGGQM5WU3FgATRcOOm3jACOloKkx747gM/Npsb9Kn3Z3+NY
U11ngGwJeoJk+6wUhMZeC6PlEOWB/43/k/zDEfHXbxH74dYkqtCRy0xEnljMIB2gvNVLIu7okKFg
eSMyDXUw5DRV1G48/pAPxQOneWtm0elWoQDLPoKue/1DiyQKC46aXOzw0AGzPONP5XQl1YkKlrAW
gr4z5YRnUw7Vj9b4roOZNcOCReHQ511lFz62kMRrYX3VfmFqiDWpahLBX/GCs/1t79hAS0hO6Pju
TxqayBQOCfF2FS8XI0JvV1Tgl5BdI/11bbr6Bx42Fil9wwH8o8JvA5/1YyPYv4Dz7Blx+eujTS9S
IDplD+LEXtb+Hl71AnbHAAglIWN2jfIhSigZG4mwmFMAxr32aBRNjNvO8zqOxrENVLTAuu6bougJ
QjK5c6b+11fk9swggFNO+9eO2OGNS/1bxBm6xIlgoGv/b55e3QmJFMdLsZj7tujDgm/q+Nfj58vz
jvsNUS2yFgsvku+txWtnnLmYEBQuuA2dSjlq3P3AJORywERO2B6r/sJEcrKkWTYx7sGuUmr71F7e
39S9vSWbYqT2eaBLUEkWm5DUVFyJ2Rveh9tdvtbmbQG/Voc0RgfsMTt+AyCEOW5oLm143gGbvDwS
SZ6Xpz2Ry6Idq+ZQUz8RKoXydWV/13MofdwUU52XDwS7PrKb2fR1Moi3liJF98L9wmIVUEPq+o86
zwKsncZvy7ZhkLeg89d6BJY2+PtYtO7DQeEI5p/GUmbmLpXFXbGKVI6jJFdlQ5W7W1dkeNpOZXdQ
ee3SPSl+X0fE01ogPUpDYVHWxsJjUlIpCtYp4vnphu5iP24bltnRectco/sprcruvLQT37FacXl6
z4Vl8FaPtgXV9bEdMYwyfYe0HV3JOPrDUvTGu5WDuOs9W8f4xdHC9k38fbQdk9YLPLEvXAnS2FC2
oah1dD3TYmvA1cc1aQzJKWYUbBtnfLUn1nt3eDKkv9309VLX4e9IBx3egW1n3tKJrkkrLnuO0mdt
pUX+EDUlb2eJ2/FZmDWhFt4cMQrwlBDSAY/vgTYxE/6J4Z2D75EMJiDuakeDXUcChe8Fn8wBHVcU
0npRrJXxQKOvge5EKNMb9DoEEQCuOe631gaIdYTWVUfdqGUk3+1V361RgjfJaBXOy5smw0nn7r4N
bWOqNWpNg44aQaXK1Ldi0F1Qu8zoxB0ql8eckVVahlwM3Q+LhPQBY9/S7en3Lxg2zPDwB2rh9Q76
0Db6pK0+ssZvhlt3zWO/ipOhYXVLK5tIVbRB/S1HtDWpb2/t5OkRPBfh3/nGGu81Sy9ZMGFoNZux
fNX7FHAYLQYmTdqbZ5pBjTFj+hYrvIHzbz8QmaBn2/g8IMRIMPR0kuvSiwnGwuM6eTQKTRm3EV2u
5KXU6zd02U8p5a1Nyge0lpmEGq+GgjtDgpaj7NN1VnkZ8R76XzNqraUTWZpG83BDUMCjK3YQu8qq
66zYnT0oSLdAes0CYnxhQwCz0otyKpsYBH58/ochjleFv82HYzW6vJPcpyiSOMhowWU32nBrKdeZ
1tUGsO99N+Vm4wGajgTxghQgMcRgp/8xXBwffykntt6Bt9Omsl+1brZCSqKMstu1zwPZdThGWy8j
mJJ6tSd4vSLXWiA3VlYbLYAaVM39ZUVSPr9Z+mbYeSuVkxv1ejoq0g2i1OTGnmzF1GXrcNL3y5/W
HV9nTAJjhdmMLjd2s3Lv+IKrH2l5PtJb8Fgvr+14g3eG457E9Xm3Ae9if1HCBXv9Te1d25Yr6wX6
18d7rgENMiYQLZ/L3EsjdICCKqI/d5Lqh7pTgokVhwEpjlbZjl8bd2/Lr7DMxEfPIEkzB5P3uF8N
HyjjpathY5FRivHg+AkDW5H2YTWYPMpaa67tZx629GHAmmtDemUnzXTPe00HHDEUP34QvdFVRVPX
fZA0+WFt+b6stfZT7bRtC4kDpeAYwckjx9yZzVJ8eWzi5OnHc9Nm81Oe2YZ4S1qkJND9yLbNagQ+
utkXTUeWkWdATHQdnkUIOmLMHru9ZoUKWbCguUjM/vUlnQt8qXHPk7DXxLUAhLWnYw//4MoRdF64
iY56OOoHFmEDGxpICd960nvgiZnYwy9cHVKPvDhBatpH/1poXfz/AXEug6fTgNw5fY5HmGYRkmmO
fqE+nnjBdpdFruaWE6tOMhTrW+rSQw4bs2INh9QjmudavCD9mXG3gEpDjgr5WABpSaKDpvdjQJ32
p4esQjfhU2frLJBnHobkz+tkClKHt2rdwvFXzB2FrEJ+LI1ofNPG7xhRPFEzoeBPIh2uSNTP4e+6
kEXJRf+tkt7pYmq7Q1u3vKxUSUAnY5w4kAnWDalCLXFdKY4wKWjNIyi7uMsHue6kSNC8mskVt1eM
49t1uEPnOcKHjPOXPW5mkG+0A5kRM1+YcewqNhdXItH2HYLPFn6MHO6Nv4K0tcyDnib7XJJnYAoA
M/2H7raRc1wD/5c2TY03deW828riqP0qdfZThsVxmV6lVqNHG8vPIpazCMNKJ8Cca0q3+el6ZzCh
3oKI0MnD0DJ1nSPHjkJaJdFRd98EoWLZJ86KdA2MC9IemjwnZ22d5JNVyH7aDqovJ1bac/vB4Dtz
Mc+HRFgbOLDmatnYUpjPtMly3M19TZRXoh99pzwPOCcoHIvUD6anKaQZB5St0/6uovEH6xQOVQW7
9gB1Hp0Cn+CaA3CAcUgUczoSeK/WwwgwXH57h9YGNd/VxzW9DcCzb0EYDrHe98kmxHqLwkRDAV7w
JzLGap5KFIGQXM2/f3jtwjoVMq4WQmBcL+aDNNe/hOX9IFl9ZSVP8bXPzwKT8FC1aGXiSXqPNyCI
nqNfLg6WGKOB/+n5q4DvjierYLm6LLeAfLk/6J8kPOQhY9mYGvTxKPYvfNVBLxlbuDY9lsjSFXJZ
6UJFw2CgyUQhcZGMpDl6BLsU8sN1ahVIjqrP753iheA86gewisW3IGXkPuiAqlRzn8DoX9IFOTbP
yFPtQ5/Wy8X0zdFCH6b0FdNzlnawdE1WKpNFeu0F47ms2rx5npqm9EQiUmCcwLGw5J1gqFp9toMq
afwgTne1DpBCpCoErFcJhiZLd/K0T1hS+Emy99pqXFPTIvaZWRUtxXFyxez6HJ1TPphuUO/cF+GH
G338u49mCZXE3Dum+2TDzuZj3HkD2zE/nNGZoO5RS66Yijvu6h2apVc3nZkuqwsOjwKzcuENRUAU
jZti+Vq/5NbMQNBmLUBpuJC+B4e9vP0rkmYYjqAh0NpXm3eHG4VOP9ednAdubLyOhagace+KDwoe
zQJTbu1k9aiJ91XKglT2Ieiuad4MlQ6pgrNrJK+HLJQmZ67As+ZOeX45UJpOK0oLiMYlK1exfVMB
nvwfW7eQwUUDJ0z5vgLUPUil4QsQBVPb9RLc3HHk0pOQSEJFSo/G+xfePQ9LGDZf34W1laEpysHY
aZTo2mAKcPCv+CtKyrtfKKgXhjbRd1ikfuSJL3VhVtSMzEOhYaj5LrUaAwfLUC/GthaB4c+4wqL5
/mZ8Bl4/mJ7JFlgv22eUMbrf6stpdlmYGhz8z/5aKEKkMPzhGZbYJBp4GM/PBmhjPb3yfSmH+Wnr
9bPtgg9ikVHMULTrEcWqaaSW28y71xZmauOgbSuxTGgwIAFYRJypVweMmE/uSd0NTIP6ZqEiouGQ
VerqXCPcKDsU//64JINoM0C2NhLkpVpwtG9JXrdCCxq6GOBNvXsc3VEuunsHoYFoT/IkCOUyeGjI
6Wb4ykHO/Q3to0aftP9CF3v0XGDPBoQQ2rC+0CvLX6W6rTe2+vqREiWGd/anLTPZVl4z+/a4BtUf
bzmJPXCW6spW+AQKw+B3gq0qu7tNcX9LoO+mVcpZ+9DSWZ8tpoJk9rKpbMac1sVjgUvoxslNhDja
FNXhB4hG0+TuJmRa7/QvgjD2r0hf7A627g7ZFIFbb730Xb7FNS5k4Tv8+bvUNtbrZOBevT9/KDNe
c1SNpYI4EmHC+t+g/rf5+b5oVzaF88g9SX9qwhZCXvulkomKb4NCmqWxm6m70G0g3F9mE6njhZIn
1RaV3LMFPcVwkZatJudJ+CoB127D9jEjs+J5suRyAttC4iWODPhp4WKddRXw51Gv0DnCYJJstoZd
bKLMbABsEqrxLZHcbEqlqSjSC3RUw73ZwOA/pmA8FAL6RMi/0WSborJSXJNJKwOOr488yseS4iVP
nr9gSPeUleG7EL/8FloDdxRtAzVG6PvHt16/Ff+HsNWGfr4EDSh/P1UFdAIy5uVrj8MT1r8pVGeN
4bncsU1S6hHCEo8ZHKyu5v7cAuQAMSq8+2Y0yIgT6CAPOlQ1egWCirSBMrNfo3qk4mqr9cLy7D2b
EkaG6vkYHCMRT6MzOWAS8Os+bZVFcmZ4kUIoGwGE3bXFQityqWW59rb8aZN8sB1FaxZNKuU7uO2I
N2Ufrl/1Kphe9vdDENerpnMaAU9o9jKnfQOLmfKuf0w2dmnG/I42gBRLJcqWks5AGuGGB1w3pocM
PZsg7hL0sGriRjWIvYF+wBPexSCF021MtictrYzyshzxy5ldxGg+VHd8s5lKHzA1jdQNuLQVr5sd
d5MlzeScleyRijksPxXyWOrgSx/gkofiihRUrYgBzglFr+E2GqcXXvAN5n1zYIc3fOPwyAFQnXAG
/ToEIHI7E0XirDMBkvUfGJC0mD2k02N6ffJ2xDbmhLzmopd4NbwIOtZgy0vY9wKeKDI2GVJR9KOA
3rSewxMFel1jwwHyrT2nDkmGlTu39xy0ou/gKz4lJjQm/FU34NrFt1STpJGvdJMKlE0LXYW6UHSk
Js6Kjj9Eokta6w2ZH16tp6HlOFzefZEBZr7l+s0Xm0f09i6/hwjUCwSgyUlbq6TElJpuiKLTpamM
u4yAlV0U9U0vmY94H4IelXBhzM08XcRaDbNRZgKiDpVQfFJXn94XeuCub7i4HK+lvroguQxG9fjE
sE6zBb0HFbRYyNFu7jKZRbq7t7+EM5rgFO8ERWTdPpMUet8zH1UFVbm0UpVxqut0gPN6I80eAXTi
ZwiWT9ezl+SSYFka+jXMg8JSeZ3DLNItR60z3DDRQkYNr3PdVA/G9GCjK3D+7Zc4YaubJy9amRIX
1jBhSDjuNkBRib7Jqh/6LyaFnsUmSnIhM2dIFIarkqRRA8CJKSVXuSU1l3zw35MGnREVDrWTwLO6
bY8xagP3ytWaCKnzgNPc6W8wxUAwOCV0vvcyl0BLZb79VriubOqG5/EaC1vJSXBfGumaHe00YjSk
19pvoWuTu9qnQU+RYcyweAfjgyZ1kVYjn+ymjzIUFElFlngxh4H8N+rTUe+PL5wLU9fztwKrgBQn
LbwPYqD9tGETBk4CXdaGDnBasT7yd9xRbUsdfKVhj7B70mc/Kw4DpOjGoyoWA/HiR8oke6FBQUpr
TiDFHKs90UCfBwSFYn+GY5woQAQj7mq6y1LVoZsbAImpc4AKPaTvDiIRtUCeBJX6e+HqCuzx/mL/
SQnLUUuSM2240auQtEuWaCZmKEIS3PlRStVT+BrvR98tThiQkvFc+46atlogVk29SrS6XkOgOqeT
aCh2ocGfuh1ynekanI9fF0uCCKLtz48ywSLCqThREf6/2lyLveTbF79NSp3/iW0cpyXIMcryBud1
sVolESVGKm/BcEL21YTVvF1xebkQAtxC7XAD0AeUajTJ2yOKvP3Oxk+anTxQC2pj6H2innx6M2dP
vjlYnxnOB43+BIIzOHoHkFnMt8YtU8D+ec78UdeOgaOiMadWedkUocDoD2lqR8vWOgnrhNd2ZfUi
gvqUKoDoOoq8SiHSQByVmfipaE+eDUSbndenGHDCq7I0W2asiymzaS/yxe7mDaivtmOesc0FK7KR
cHRQEcMmutDM01JdDsYQTUYA8T3iczcDaSNMfz1M15VE+h4nRd++gW8SsYqIK+6QVMhuS8zGd6OI
dk/Ev6eMIs2l0Y8f9kCVY19rwcJlwYkV2AjkGNA+ejQWOWxEZKIYAR0szYXioPsxe/N/R4bcT7ih
EoKPcb/42WP0w/PcEkIfLNy8NN72voJwtF57YN0hUUvRBwEcwODdKc/NP4/14ZGgfOKuW2vGq2cf
AEfTWZCHoqLMjwpOHMX0oEelO6H3CxR2WWfSmAyMSeuMkcKYJdRsXK4kY6eLDQeFJ5Dei59YGai9
DuhNLuRjWsoZPFDMAt98Bo080/kGx9To1iBDkoZa7xdLANOtAB0Mmq9KfNaQJZ62CdcRMhmNk5Ke
WkLy+PKq/S28GUt2QfJDB7jKx+6ZGIazsIlFjkgRkl/O2uVzOe/3RlrjGCUbDf289U1za0LJhYg5
AG9azzylAcUbRWUDxCBp388bsu2EWrghaU4tUyvBfKhd5xus7pLeb6p1eN7RnGlwTghjBCYBqx5P
eBzLZHWHyCVaWMFgdsc2SLwSETOqyLkI5NSTarQCF6bs0ljz2D7DcCcPSHPx3lXGN4xmxwsXxW/3
9qrK4TDoFUqkzPPAo6nNC9nQcL/blU3vccxA29yAMMgP6SmjMvdrrIwfmFJsB1f8SJmnXnn3MNAj
nvc7/xtwswSjDiFLHCqygd0J6tw4ntsS5WGIJRnnp9QD5se8Yg6p8DJseb+aw04zk4u3MI1ATEih
39yiR9U/Przqj19xel7JIDVKNPa+pJrZLsVpL6c1T4ZUuDVsrxSJzueSq44f+yW6Xu1Oi80S1rKs
Lc6bmwwJKDKOmrgFrf/bu4xTg8p2LwCovUKXfLIZ3E7B4hgoFkJK92UgLaRo2+F1jgf9hXRfTcpL
6T9Qe4ig7liXbepH0yBAPJKq1TxCo2gUnMweuQdM6l7Otgfm0apytbjipll1KxXzXz5BKP88smm+
jnQF4HuyhgHlL9gjaem+dVSV5+ey/q5T5D1g6bAdMyWp3b20G0SoVcWd/W23fm01He39G/6wnkPM
Iazya/IxY2KAqJyZcf6aHFJnCP8XvtZ3tOCwlaNhlAdRrvojKVD9KhXSL464CPnKGxQpiwowP95K
I70WU+YAmG8FjggApLnB6qO6H7QcEk0aInQXUMJLXcV6matcFxAMQYyF6nsa5dCQULn6LHDctrGt
x/C1eABCVZ4q13Uj2MgZE582l5B8tfgOUJnP5kkc3u0HRhnUV6dPoqVZe7TRP+cNesu73gX+2DHr
sqzC9KUtRBJOeovx6M+Km4IRDVHMjkUODNPaYcPjIC9X53HPeOrHpRNH/aUQIu6OzP0ok8fV/O5B
yeuvPLtnWxXSvnleBvSnTBRPVXjJX/hX6173dH/N8/Ea0VhCIabFfD5KS64CXa08aGZMSVJmTK0j
TJHUJ7TN+v13K4cxZSEuJsSz5S/F16cFlBAmOv1teNQbcuZCNW/v2Z5yVQZsjmdd4ahg73+195b3
8d/lHgMO4qsJeCM8YTQ1yStpBd7/zCQjBfgHGwSjGwMnbKZmbgFOyxrAYDMJ64G1SsaazSRmomOF
uTgcUgDwpHa08YcClZykbNe6TaqCS59tgrcfwhDDEivfOqNVNYLBPmtDYm9MbMTW0fSPMQRkHA1S
HClymAbfyfnarHBEGN2zqP+/g54J6iFU+baqHuDveo9LB2ZkR76A73fps2H58MvjvUadFZvs1l2o
MhCXGVOaJgW1i5151zPKp8NXPCUgezFgIdk24dUsT0tmaegEZNtbdFXqMPIl5OaIIjbbkbnxvUjb
x0639KhvEe5DVsWabJmPnhSLvZ8cGcv1u0tthNEBqcd91G7rfZXlf2igC8O75qxKDyaTUrDTj8q1
p+vlVqGdY+NBKZZTextpdTpKDZCKJj0qLmBem5poo+hnOoeZ91Eofadz9Ajob+7MN+feCAFJuCdE
jC2St2FtBYwWCfhjRe7K1QvxTn68SYDr6ixzhpJQ69OOZ2i5fVHM3fLoC2ORb0/Fbchb0d1oE933
gtMDHqeH2X7IInYiJTFJTQ5Ev+1H7saBJSqlJppSZiQs62QkzJCDs78f9+1MwPRJ5bAwWK+2qv3w
1HaHxx7lKjO1jxYlolislcOLkLwyw8uQ8riVL3V/+UM8GrtyW3hwzs2hPpedxLCiRlE9oB57GZKY
/7FQDjpD7mJrElYiCHXKckwozdNerkVuKInp8lTm0c3pksPsKnD5bNucDeATwzN+S6kNe6pJUXdA
b0cjlq40oNUb3E4kVxNX+eQl9qdKG/6vXuHQKkVKZH8N4Ta5lnWiWp/E3cKBdUe/kn9TG+JBBrOa
NQdfd3wYXIc+gzV9PTqwFb5XZiIGYeN1aDlepSiSPrXwcEqb0Tq8NjyALe32Aih6to3ERg07rYwi
y3ECCfF/u4qt7vFlGm+eEyxE5JZEK4hokVYj2L7oXDRFCP3/giJfrwnQXH6OaEO+64l/PMgOSPaP
8ZBbpBX7eM+YGkOezKNwHuSOYw5poU7VkAmQYUTViEtmwvMBVVj7QCUMEIi1krUxRFNRixyTUQyI
bFPwR82tZ60MAz8GEdQ3F2EEFGVcSQ4GsixuDjQjz70hfk2ErqVb5qMb1pyBpJjjxmqxyijnP1xd
we4o5kU0Ytoiq1hjara2UXr81DDhIhnvn89s2RxlWPHbmD4MXVVOjqRcVKgtbuf9yFGA8InoQE0b
PXChips5y5RQE3na+FABBPWY0/Pbb7Hxb7rwDLTbBKVa2083KN+9mtfe85ITV/n+0Bn2fxnIHIET
j5/U4TV4+eTBBWEoxtGkjjWyvUJqq0ZwmeT4HBCIQ7ijIeyt1kguZUaekwiU7kZALo5ofI/KjCVC
DUlZzkA30V5yMf+32idXfiB5MdXxeHdY3xe8Y3jD/jhBtzgn7EXZgufNpSlS3S+/DD7lkLTbptTo
o08EIqP7zvK/w5S5rsLIfjAwrK6McHtd3a4/JME+lBWinCqhRiiHGg2fxTwdIJPa2g6JGdyRaRBp
qL6pqIBwShgNyzQymiiuKgoVXWYU3/do2CEcBtQmDgHpMNsm+gvrqPA6u80cU/oSjukL358KBON/
lEUhtzQkYm0Spv7IrdFlvhM26xQAFAxtXocorDPLZRMZMaoB0CZVLRIYaIgVtr5I3jVf4jUFhv/7
QGXO12Bq7uIM+AK0Do6QfJZiZ8+WFB9Ha7GopX2Blj3n57nhsrbnxUiOU8ydFX6pD/STyfpiBHs/
25+rN5FBergzyqOgc/vhN06EQXuPtqRdWGnQKPQExYDc436sqVHq+y0BrvJncimsDEgR2JfxqWXo
LS2RDzIDpkBLfy0nHzbi+1OTCA4Qm/Uh2aiZuoNiOAGjue+68kvzvKxCQV4G8tCCkr3RMRE59i2Z
VDhsDua3OB6ZzWutR/tcShkSlXEac6SbKPlXBP6g3pRI+dUQ6Xo52a41b9lmx0woQx0WaOLsAdNF
R8ZLcfVzR/0SDtQNrDMYnQavy/Mqb2+tS6BHkBAcFJkLsU9IP3fIEVPvNDSopZe9HfCi0FuHc30l
Yknz+enblTt7a+EgNBXv/blo9aj6giTPb/pmeUwkaFOfnxlY0887KpHKmA6bnBCwzvBwUZpsWIeW
LkDP6M8XQxxxhzwReRH7Fd6M/dH+toUh1GSTY7GGA40I67c8d/rpGJBNUWn8wUb//U1QlesvrIxN
hcropf4l97SPOrLxKNqms/y1OcLbBvIDghNwMFXeiCyOwabyrlpewCq+6uxqIU1byFXLSQ3CR5Hc
wFmybSt9eizxqQC+54goQvI4splEhF9p8DNdA+EMm7mIvZOSjxggobqgYyqWBjwn88HbxaeRWEFv
/I8JnzVjd8nCoUBN2LBdVi8FD7H3zPWtUs2kpMoWU+R5L56Sx5pYD+rJyYMWdqXt4xbW/MDMQab+
+J9j6lgo3fesOfTH3P75NgBNUKliBVByhwlbRsENiOyfLk3c4eNmd7eCyXnI95PrpDiTCf3fqJ89
r2Z6YibaQE4kA6R35CTYEJ4KegiMyetfuly0cND28Pm2/HvwrcFQA9wyPT33Fyw2oe8USSv/RhJH
HP9pSrlOepwyakmyz9NKB2FJmgjxQwwqkYRjmWoSIqlI5xLKXXvEcZoZxta8ldBeiSgYZcwEhvUm
LUDB9ukuZKYfv+6LubcUAGPkgDe/N5XXlgAp31yZu3/zNoZqqJz2iEtUIZ9cjB4uR/nSYTc9HEtW
KCULlVRfh5DbnqGyeq9jQ2qmKb74hUJ9/M0BzjYcSNKYNCY20mrPo/8kuRP7B9DeYckgFwVjggKP
gMg7740ekI4mnVFmX7z8dPY9k7aNRAMeFMOBZbUXVpIA+E9lEUDZKdpF01Vp9pt29ZlX6uamSvG0
7wqS3lhmztkpGEMpFBeBEVJjpq0cUafjuxBxIdGq8wQxAqXVEp3LI/FgPT1r6foh6+bzLDqw62hU
OBR5+ZSpip9NZnGdxfxvKYaY8inD9jYps8p0kCDf4r8oLxuPuEM9/WgtR6f+FVfoWX/T5lGYWAWY
lqTzgs5iHN8osF5u0GBcyHENDhvl80IPj7YUTCRjZxvJxWBfAl7MHeHTonV8+4x+MVJihh1jldAZ
5LAV4DTbKwfe2UaIWNqXbKoow595G02aMli8NTmqi82+1R/tLVOkP/xeOa0DVz4YBcR/Pc6dQglb
aQSwTzQnpjIeNrdMhXG5LIKvlkEnUim3UnV5bk1GsUvAqqZHzf7F3QqY4XDPz8c4J5rkSGDWzlMy
A8tWWHqjvTyAV+eijRKOuAIcOhdfMOxq7xnUWj6CC3/ZFmulImp07Yr9/Cxo8GzoWaTr5VH0CQMF
W2bm/j/SuVkXIQTtiSnUzpJ1AzmGSX4t3jH69Pak+539Zb+0xdgoYzNrZVm3UExbjo66Uz9aXYSr
7kmqGOnsjM0cIjdU9kebze+OLMzo7Jtc4X6RgxViamkm9Dp36dyS9bxQSo1qVN9/dmA1q3VWGU5H
pUroGOZ/6MNxgP5vVOPvVJA0JAkMiFSYTdUKU8phR0qI9o7WPFFHBemN3zJxBqGyEDX01eqQZGLe
G7MsnPZ7o5mjl7niipTHEoYQJ6l2Rk5LZYv85jn3PLMby5H8x8p8RNjAxzemesCvrR9eOJhmVY20
IOvvZzaJOzZP7Fm/wUng+vBH74rmcMdpObvvQClByUuOlWakDiARquB+64E5YzKEe42wwSyzDsGW
ZJPq7pnDqIaoW3alEFEfmDkG0sfZdyqyXgRIKIpoT1bGTt9cimk/TaVcxyO9AxtL19NbZs2d3Vcf
JtAFroIbwyB3Y1b4aGuR2uGES6Dlembz3BWwFaTFAHJR8xlJhjcL4PfzNQiA/JylgpV8yZYWQdCV
VKrPb1Vk2Ihs5PctIKK7lGOqq9qV9H+SzHTOLgU/9jIfCuL1mLXrPu6172pIZG05/lEKk6fUTat6
KzEzprxOGIXqMJiDMmgPO8WHa40i8EoNvJjLrbfPuSpViArIb+sqQrPjPb77phVBzRyKykgRUoNy
MsZK88rFZbSkHSRld7TVvD7EwZlLu8lJEzVOGDdvF7M+Z1CRd90FsAAZ8Hz4GANL4O5075YTHys7
8h6LioBwcGZG+QpUt5P1US91NYIysGD31FebdvJF4LQ7bU+tw0Vsx/1bJNsaVDGPj5X90rb2WeRO
6fjm2dDOUInLXANOL85a96eIgWR0l+sQpYiFli4OnS5jdR+v4n4prKrnpEqwWQzHR3UOCCsLEbX6
q7Z0wkKtQz0+2eq9yeESlBA6Geo4P/YsxG3R42+pB4oVu7t3xLgoaYeLGDz7Gw+TfuPsm1nztMsU
wdSVCcjy9iJdxGbWrixduswrexdX+hJJ+LCLA/gdvvOBQAEhVgyTniqZq5DkKal3Xg8GKrSzPcuZ
0k4kG1SRhUs10oqlfos/E/U4HIVxcx4dxBogg2Q9ia2ezD821kJwB/NPVSwMNyE16vk0clrEpk0y
XfNz7tP/CeLZgIsRK6LzdeX0MgFYDpH9pth6o1xXXj8ZpUhPB9RNURtCMo/mC4BxYdVYFUomC1zM
M/4Fs1FNo1QBFERBthMzilcrOIKr3yRre0RqeXEZrc3YL6SzbBOBa8lY7WeZu8CzvZEm0xPybOxl
BPI5Ac44/M1jFrqpolOhtnMWgu0VjaQWiZMVb43LS1HnN22IrP9fLtOO3wiBda/Acmrg3APJa+85
3I/kBYDVXWLOT+S1EEFCHYw7mtuVutm3+ILHQ3rFBxpRO2COwZRO7aLv8/+UFDvuisoTA31aUhQE
mnwwj8Qi6Dnpx3hGzfA7tNSW/+rQQ8yUhuOYr+3RoDEtE8/6ti0Vb51Is7MEjKGocCnsv3b7TC+l
cWfu3RIVkzPlLBVQR9V3jruQm4uykX+uN+3VTmfwqTx6SzVtLAFS4wKH0Yoebw7tUD35Y0tjmdYr
Ym5uY7Um2aSvyIjHV5F8uTcZ06EUw5t/Wl6QOpBs4TzdtJdFe4ueTFdQAlojklAAtHdMhMayYrhd
30Ghi6tPsHWBwwvWIu4C+4Z0kzOKvc66FNfOPChlGa6pzt7TY+6yLAwro4IBZjWaSx1oNC8RmBEX
Et6PyreqPEQx2uOG2ykHp8Yzdt1Jn8yw5NDWn44DmRq8MeeYQBec5O/LvUS2c3LsY3Ry4hqe2ma4
q4Os5kEOXIvMEbwEWXGw4zHZiRYh5D4pPJ7e60FnHS4JmieDd0hLfx80YZPJFRBnd8i1kj0/C94G
NbdGR7NM/qd7s2uwdIGBO94OgMGhO5sRK/fh0UEZRf8UPs+uZPSslWi9ktFqcYbLw/Pb7+P1bmRE
2XiiMYKQIw59xkEblv8Q4M7vEBQvuB6IuPUslhPP6zeQqBUF4N+y6KDlVu+lq7NChSSGWIIjZUoR
8L2UPGvybs+R+8JimopIhIt6aYAsTTZYX2iLeSo2lI7Th7l/lH+kiZ1r/ML5bINOGriMwP3pVaDZ
6WkgSTj5lujq2p3a1uWQkVr77vxGOAjMNYC2yFQgWQ1h7Ohu1b6MkgrhXQGOp7elKC/FYa+ycM3Z
AQEI2azqM5u9T40hngWAUCEV4SPMp7pVvrOSYQX7q4K1ekSWXZL1bMKQlZweh0DXbhia9Owm45P9
Z/HvnIv1xjdUF+MspX2NnEHoAIyRj6uRKBSTen7rY533XFgYbkTxmANrQZzSjwjbUOjcKHNGG1wE
v1HZAUFMWSM9mz1Dz1nn8EF9eo/Zk7hxnzQ6pwULLx2mp3iHbMSzT0baVND8mLqYK1N8zWRX7q6K
amOZ9YFp7cGH060VJ82ZTovhaTMJKFbB/TFnHRfIGo2sN2hsfbM3IlW+MJBBFi8z62SzH3Tp8Yoc
rBN6eOLGllqql4Cn6DRLQIlOvz4UtdDFVSAifAbluYnZIpoDiB8zyzt/Ic3WOHUqCxmmrbf0wHrk
pwuFvh5/n2t0MSNSSLb2y86vjCGzzo0AzkHS7Y7uiO8g7gUsWF4D5Jndj9KlWNxbCEJ3R1esqjug
VqeH9PODBaPyl4LIZt1fCpV/e/oet/CoCoYdxhYzoSbm+HK/GzVtKnhuWFMvllCGoeu87bu+vpeP
tQ1ZlF9+/KVF4R9FHB9dg69DkANDtlS5VSYJhGW1LaZAgNEAFCue7Yu6ML442oPvy8gVGrLVZSjy
D5TMXw2+78V8OoOcEy2rJd9q1yBX8wZS4uDnzAwWYtcYTnS3OAVXzBFKQDp85DKRLVDGKt+xFjv4
bhH3bcqh2mFzUXSoJWn08YrjxaGEggV3aRf6I+UljFmMQNCv04ch3GVBKtTjdXHxaBo26p3SYN0g
EoafS1v56rWFjyQq2WHzoUZSmBUYAej0ADDdYuEKJuilWu8S3VUwmVBaV9TaLkg1+DlsyzT5ckgy
YjFBjYVVFrWrRWDCIVcvq4OLZqbXQW9NLrbM1jBkYGxrhensC5UeZxy/xGKD4Exoi3Cj38xiaFQP
DYEx66ZJiXbMagIHC7AiKtCyYyh2INjZkTOThvgkx7pCiqLVEpvXPT0rxfnO52D/n2tOE24J53/2
/k5AJGhpvDG/KJG6auJCTreq198uYgEKL5Q+GjDO7yKWkcdmBdX9doZHrUdCiDqcGitbYyejt25E
2MxnDkiVnLEwi0s0RHCwztU8fED8V4zuqCozEHFjzGAOfqS28jq4BtvmtXp92AnNaluwaCJaQDrZ
xRgUKuKPpj9fS0IGqhYsShySq7HLttdy9zR81q4YaYzNLAUcneaQWpYYP3XsN0DUxXCtmKcq262u
7E3nVzCm+XPfmghN6E+Jpm9J/yIffvvnFc+ulVOmhOuQElqWkXZOeFTisZ4z5AlxjlmZnbUale3j
td6peJRZQIcvmvImhGeN2GovkYcJhSuCrC6FCGlsTXkIG/2vdAlx+HB0jgs8ufqudYdjRi997OSI
nLFwQWwOrXCjLakU3ZC+mGfXCg0gbhR0+B5l1u9IPk+cpgL1RjNxf6/+J46Q8CNz4OK4r3nM5k5m
p7Z7pZtSFyqwaGpE6DhVzJoOWM1s4WUFOSAPPtwtVPuHk3cui7k1lXtSuiPoyOUYdp8m5MXJTdXj
TkA6Zsr634B/Y0C80TfVD0b+5VCYzUG6vRgADxwnHdluiL1UHghcT7TmpARrv1L4nMLoXIZ2jXSl
lJTGu/R4QLchg4jGqhRtAUJDD6DVYs66DSHPxGQjMz5RsmhyMhewxKtuLRABSUKgABr0hwt86qtb
DhRYI4QWxl7SE9ujkHx1iLYbPNHL2P5bkIKfL0mN1KRV2MfXkwjRpolmHrbh7F96pipkuPbrfEOi
hQYd5eSsbDy2bvYE24/whtAYGuqk5SqaDGpx8okbqWowNYQKnkqmxmj1iY3vaqJbpaA+k50BtJTn
YSjG7R4nFu5jQQC5KhqYNYC88Z47LC+cvlAAmlkdzN9My2sI62IJ+1ihznn4tVx6Ru8Wu7f1ZAwX
ALXK2Ehrf9Pt0rsYhYMl7Zzn1wkqc7+WWet4uH1pLbiArUA81+k8qfxbavXgyM2YYokP7agL0kma
aEeRdylEesU+p9Yc1KjKqTrYbM3UIsRZ3sszR4dWOocKJJqBTBH+QGBa4UnWQLnjaTqbM9Di8v46
uJeoS4vwt9RD5PjiWJRKkb8CKdVHmx79h7NKsefyM0uQc153TfNpd7RQWINfWEKjyYo/aXcIXHCa
7zh+hJ7a9tIJQlHggcqMZ+JBmzxTO31zBS4ts41tNitXVVswnVejQsX1B4fMR4N8Wqj13NaCjKvS
V4jNNb26pp1U8t8WJDof4yws72hf7PPWdms4+KSlulANGxKI3iuWwrS/j1IoKg8Hdr5Z3BunXYnq
Ps65votERV0pEk3wshwMx2A1hLOdeo1k+I80j4Go/6WX9Z8KXsNnAfu1kXavSlB+3Oz5AsLN4cRr
tUI/Cc16YGFLwMX/WYNds6QFraO9CZL3BkCTjg6eT2zDbxCICykGJ5JRaaiZavRLwisE36wprwY3
EzCZuT+Py/DTdW+4m89Eqm+fxOfedoBqX4ubakqhHD99o0irwi/2gg/kBE8X2VJKB6m0XvC6sgyh
JfllAC39Kk+gI67h5BY80oH1xd//viTIKtbL1c/J+s4AmkysygZTJqcXFT3n4Zs4Mvc2ECRl5UZW
Gi4WOOZEHgH1g5o4dFt4bO8B9JKDakZgCS1Z/dnkE4+w0TZgs268NpJr9/EFj7DYxdOOhyPbjrSs
eWdVyfb3hdkHIydLIiucNA3dntyjQHF6uqSj4tI65qU+Lq+pBt1uyqVTJXi2cZHGy2WyHBbPU5uD
2C93h/kYFBhUJRDr2H6iHAwQlWw6KHjjpNLmjMV/T8MtsjD2Odmj9ffODpwncbn0+2WrDg1uA6v9
lyerabU7zrHP4wuf4F4A1Ebp3SD0irsIyr6rJ5LhMCAD1YRuDqjzCV3TJl2n33EWEaowqlOpT46T
kFIxGLNVz9rPkMVdNip46BNzm9cftGA/Xp4UatZ/EgLtAdPRaX/RJfW1baT+nDSU90wz1p+wW7Nz
a0vyakU4BUCRZcM0Hc2O3kEkehc4nG+TISZ9u6gg+1WTdb9xDh60DEmmVF1P6DJhOPoksTtqaZVR
3AukG4tKp1Ejf6ALE4q4HS3sjXhfIdBZLUUpNhcnEP8IQc0pcHDfRUJJMR0UgNSdormKiSrdl9rI
61ItyaENFRsfbpcyyfpx3suyJXxaU7bO2RPCbn3796/R6ABwd1Gqx4CzI8lHc51m+KcvQXyuOwur
h6OtNFi7XOaflIKSNR8AMRrc5tTBcn4lRtQjbTXIGn9kstPGzQA2JEYJkOuFpxWEfJPU1whb5k6g
ZDfU/2E7QqBDNmbH9wFZcOkO2e6kfz/fusydDmspqFc3Mtg/rqxh2KI2p3qzu/iUVgHDdYOaNRly
y8WGpGABhaVJRxDSXBSl/AXdKNcdi3dg2wJkwbWeJ7OFNAe/v3bcw8bz+NYMdtAfXaECJ2HWO+hf
MWyRrfZ6PAZRO/uVY/cCbrj9BGVdZ6orxrCWwWBpkbJWBsCz5w28XgK5JEpuLOSQ2+vTu39SpCJV
fJLjNLWpj4/Mj3X+ZMF8IdryAiq8sOIb0tiJBMS9rpPaj2LB4sYrLs02wfsQlsQ711KrR6eAV58Q
VZtzB5wmKcng+VXK9PNlZGrawndAAx91DiP2zinS42h3EmDpWoA3yJKquFvJAcbIi3rmDaTBdHE2
0If1bCAmC7oexZ4O8+JxRrRFp/OIUfmPghnYZ0PE62bwjucKFULZ5y7w2QJMiiDoHsnEVzGPl8W3
L2Ztw6U/qyv2DiaDoj9lIn4+EHFKE+PBTCqUGyzq99nSs6eMsKbDEBdgTyzxi1jHH6rqlTWcy8RI
dUtC7CWX47WYGc/owtntPzz/gTgXuDy1YuRVXYTpGDyiVV4S8CNwwayGd54skKVZPCUEOlVegSG0
rc7vn1GTbteknrOBWxcVua/O3XSBD3CbzMIAyO6YbbAFlhQVK2WqSRpWYGYsQhV1bYs1cVf4quMJ
A7Baf3eaUSQs5TKSh3wr2VstC/DZXhJPOe3jfM000UlL6FdbejjBYA+rBvqf8MIz1RVqgAn8eEMN
1FTl3ZQewIPlOYiZJ5Ol9F3YBS7ylaJKkPcX11OH9JjW9dJ7Rp8wFhh6wj7VAKZeEyiVQjsYYwr3
WaQ+XiryKIlh4/AI68MKdY6dWCQYI3XPSBr9QElrQ+QLMon4gO/thq7ok+rvh5/piM0IDFZgnApy
Q87iBOYcaPGCLm78wqutdvdaXpOZqwVdcqW5LaGgnIbsSbnOPovtFiqIQXordup8rArtmLO7EqHs
CpwLSGjpVzY9K5z8pJn4tGu+6ZzarYeiRQe9nuVqz6tCKerXXYYuUNIXrTXATAKk8OkDEHSUE/Jj
6vyvlMm+YAlDXb7aJTssbPm+0f/4GMaQxOQko/X2/Uz7Ih6zmphGvR6TdHFmTiIAJ/IsC4TfNyic
aOmBxPzNngpHTqku6XLyeeVS/6WW4FLbmTwCIQU1vzeIy2no5vJAISTYxi95TVmW0Ll8bO9wXjfd
SxvGDXXAIdS2SzeXoBTZiw7GTAc6MN5zOmwrjpGvwYhd6aTElhaPlH2KKNtrXK2tKunhuj7nUijm
S52eD/sZ8Bl5egOmS5kMUg6d3O5mxRn3SyZ+YYR1yH2Ja/kXopgWHHj8KvenYU3xKroEGZunaAY9
ND7oMgqmadzfLNcbKsnPSe5JQPwSa4QkVCUvRVDKJRBoZiOET2eo2ouLxPq/0l5vBd4SsrBfIh1C
5uCgymKm/5Fk8cNHaQFCxlaPPuT9a0DinHIo4ECvATPyIFQTHvHq17ncOyhwtT+SxmPqJ8bovzsZ
G1Ppto6vNAcoHnP5iGgEmAKH9ZzlmwX8Yr4hMoMVJ2EwMm5wvr07SOs3AiP/nRCN+3+Kqe705YVd
bnQZvaq2SZg/532oO5dqBnhA1GMEP1CXvQzltUqNtgUR8i0bs8CSIOCXySE7N8gMCLYutM6UO/Gw
JiS8fAm+oAmIm83NPlww2cmHGzdl8+zJP95q55b1rSOYjkVZYi6lgbidPkBslLuOyIhAL14ViPar
gqc1QPGTHBCrVWiFhlBIahQ2HiaBJTBoaRy2hMfNpfQH6MtM+CNSQwXU1FtC2ABhQlFhTtq3f0aQ
G7qvSCLDtPnShrBS/yatrl4B7HHd3cU72aXJljtTuRYs2+iqbHrh1bDxZRpNJDSSGLpHIqtSzAYY
H7KVZC0uA5cj+H3sovkogEM0QUYYQGsKnB3Gc5KLc5jlVzOEl0X3z9lghR4Wj58pZSsBlmV1+gF1
iG2AZ7EaNuqIQ/Du4nFWzddwzkQMPfr9lSEonUcA9cQ8hfy6SHjYV1IxlQNgoLk/pyr3GNMbmcVd
TyvYjQ+29fIlIxw4DkIUBfGwctlNgllPpWwoNATbzHqbPgXdL86weIbaXBp09Y8ITzZUjOkxvzIV
lD/nRojrY1C7AD1IiliWYefPGLptl2jK73yplzNKrA+vJSyykAOf7panX1MY1z0sHUnra8TRlXPw
L+O0kvkh6X3QlGRtukzy0VOrG2kj6qExHzpq3PCqmH3orbFs+6jg7Bq8Xu7ldR9QeSl5CUnxSClX
mDvGFI8D1vad4xRrfppWA7LtAiHgU4KUDttG7u5vLNqiDXlGWCtWfg7s3qNMGvBlVzhBc2Zkjl/n
WksZcza/P8MrlIKA4GUH/o1/U/QMBOImolFn8jQlTVERDd4BCUB2fDz9KiEbd9/B14+9d3QR7n/m
iO/TeQ9cY52YgjrUH0PN5agP4j/iKI3R+TDL9zfXd82NW+7vXfwf4wYNpwxHlAJlFeQZPfg26Hk5
nOGIVN430WWz87PQrPzeNWnqfbmp2WnrhFtyUl5GAOsPnDkuD/oEJds+7Yuy1OxJYAZnS0eEGH61
JpZQo3QAGHETacEBz8RCgkR7GGsnxNnWsODrFe2wPK2Bb2HPYidy4PR9o9wa8L6pLl/mBtNgfuQO
+xGKPkn9ZHhgBtmd1GbNTpPT5p6bRW61RqmwJnilsbch75znQMMe97TIalyXO3VTCDXB8yZD0b95
VPa9r0KI+QyNZYKjsAdFe4Cnds7aNz5Pj6iH04OVedj5mWB235kQFu5tsZIDmkQJ6D7/zcTHyryR
kS7HYfZUmXWBOlQ84PE0Kjx/5INrhjNXZIuXrED8WNuK61OVymk6/Gh1HDOSDxZtk/0bjnkTTaS7
71ciLGuTBrpMID9H02gAOqsEvQm33LYCb5eLe2hauxoHftWJOjP77KWnA7cFaVmT44JCi3tLwOAl
ORC0Xam/D6eM26C0aQhD7bMm+Sus3NUFUFQCsJUO9lk7Qe+bKTrzSULMKaagI6qDdSiPE/kI071e
QslGcSq5kzpAY7LWWBs7ZJO38ll/nYgzgT2SSpuiRz9B3xEkV6ncJsbPtwee1U/KCBNECgMWbIb0
SZewp7nn9op760GTUkHkeS3WSINAfUk0sKSae0JxC9RE0/5H2sK8Cgyvpx4WPqHKwH34OKIZHz7r
GOLDq4Q+bu4AWamOQAMZcsNEnD6O4r84u8JikyjCPMntfpnrJ/l3YBq40yCTLYdWAT3MWGge5fA7
pklP8lMUykxR598ueK38dP7bcL4KpZOLj00e3FCIQ9Ak7cDn2yPVpSXa/7pUjnmnq7yxGgM5Poga
lNo/KGAduHq4IPau4BDDoHGVZjFNucYTFmLBjTe+h+qSpjyi9bf52IiDlgGrt7BYHqK2jyU/rCbD
RIvtJnngYNkYnTm/zHdWe58z6rb7GpCEBQF43r3HvGH6YkCIRzgbWJl7/p6Ehk23nhpa2s3nfhgN
Dhw+rBlLRV68of0Dlj0NY1If+k3WBxcgdqYm6Qe2K+heJZQXdWVSRUHMTcoi5Bp2rVwjn/rfF8JZ
7Y7Pzl2MHCKIOd7KcdP1nTzFshq0e/3HqaE1xXsk7UwUzNtH5E1hfg6TgxN01BsMpzLxtDPxgW+F
xnSTkpyjMHX5vzfVQtXRqpnb7YfyZeZm+tocVWrQE2xNSa7bS+fCtHr0r//VEypPbHNHT1+L/dee
xyNoPGTDBSEHyPrFN6P7o2dzqla1zENWb4QHBrx699d+4YZOpbNlvqEs59yM9QNYKs3manh0ZHZa
MqTx4r9nyJwoF2/Ro5r4VaL6SVq3gKiH98YXwlGiIYO9WW/11mnH3ZyKCz4vYjPl+nltOXiCECMA
Hkic/0dJZYJTpJL/KhfurS5ZIiiVY2HVocUzQzW1DGQJDZkSlTcWZ2svmHm+CIPSrbHoGpr27tzI
vEUtZhi7/estUELuDPDg2rrgiuXNx7bbykKUoJdfJauZmnYK71rmp8JYBLoyU9QnbbkCZB6L6xGf
2zec/nYdDH0bCbiXnthjqALcPA4PslP6Sk19BQe/pcFWgNHV9QvF3YOYjBpOZEW7DZcuhes3M0vY
YyY3hXfgArcv1u9kQRMjkSgEp1LXxGiF0vaEnWumNmE5mqSU4JsfKyg+yddBYIXAqk/bxsigAMmx
8WdJTF5A+Q7rDvxt7UM6uTsqWaPlQh79O+qTfOT/BTwUj4v3wZWUWGalMnsg2eaTqKEvR3bM5nti
hU46Ps8rfyuvAwdftxWzwcsuO5+Y1aSkj4/4jwLF0jN7CG4n2gGZC2Q6QQjhjh3//AM9EHUv2Nc7
tQ2BB1tbXIz0AknKBVlEaBjuCVAz1NKXg8iu0zmxKZWLWQ6GKuyxXOTELcRauhYbcFa9G7QVYkWn
y9Y7NMiIWdUgP9/9saPiK6YNUlXAduzvQdxJp+iyk1DMPgPrLxi2TWbmgxODyTUqlwLijmoo2XTC
9MN8RhnVrdr53Ws5fim9iykPyGOA4dtM7lBDaVBQc4smqG4NhsHyetvjKM8LNFXSM6/tvGG+JC9U
fO/zdHQ1ptbgpxsoX4kinzueyNR5boh2j8U3n99QmevwQU79Z94wYUW6SCwz+T2/zD7xBPJBi0H8
iuATMcz9p75WPCdVQexaxiOdii3IdnSUO/tvU8/ex81+8wZJjdXkwgFRALcp0H7YQhjuBoubog4K
53U4flmH6twa5pSDIEILuWQ6iPChSJuK1aYO/cavJaKHeIljzuSo6j6wTpUijBotTcHoFrzmcb2p
jPoaw8kNM6CokprK9ShWh/Fd2+lj4PnE5cmFtuUjnbdoCeeDzrMhILGZfPzbztf+TOtyGZALgZ7w
o5W159ZXM284vO57xc9eseC2A6/Vfiqzfo/vX8xSVsv74QldVKkX9Ww0E+Gr6InhWond2yt6YK7g
bfs528rtPyLJ/esFDa1ndgBnn/ZU/gjIE3HMlvGxTmLoJfARSPnpPsoizWoFyE96no3AJ5RdsOPD
vfUEqimwuaM0xSg2j9NZn4eQfvkEcB/ScuZ3AqEdNLj9/++1ad27eSJO2dBCLAjUvG0IYH65E2to
aXz5w+FKGGf2CQYsV+z7zYCdLaQaXzbCZ4eu7LXGcuQed1ZQhVv/2bwMnxTo7DeJRlSfWNsNC7bZ
gvEXpfHXaJHWd4rvbrRceyF3HZ4XOjB0tx5BB+kFkSjNQTQE2wHX8fYvjc00dMtAmdKVxxnXJut+
6xdBW4Xy7aU2vW62I7UP6Oj7xfPkNRDhDQwJoQsvPQzjzPQNk+9o6ojt3jFrKFdVqSKK6EUOUaUC
KgeXOWQPD73+Ha9cqINvpe5CkkspyrTRIX3ZigsnYyOzu7DXIikFkyQQ6UMR2mNvntiKdgZ3ramt
irEZyKg+nA8XGiciIt3KBNOYFK3yfutq57/pC7BFIAfdOf/ijCEcOEnQSbB0u6SIPeR/VXHY7ogB
zW+k1lWT8Mh7I0bgXdkDNHV0olH9Z9Y69XNypQCtM/lmzYg8RyRaiJGXh6Wh13eD1macCcay4R4j
/CG1bxUAF0gNNO2DTgeX1p1Jyalzh8wFpRDIaapk6zn8Sfeni8LxsL7bMBI7GTZARjcham/xjzqV
keAM5qVZrhh8n1w+JDZof1QiJgOz1BNQAWYUZKg7WZVG87SUmmPvzcj4UjIsArjwpsoCfn7UqePI
tG1jW99jB8Eluc4KwkrOLqH9nH65qjSgq4BuDT/jnCdFU5ooq0nMMDkVrQ/OUt5nTNoSXR7KAnTS
bYHUPwoAQC/s0ijbVqsKzCVrYS2TsSeDlIyK/IQE11wF7xnkBLxuA/PDYYTpAb6681xrnUyTjFPh
W9vMbS/0Ah6q8nNfp7DvK72zbV9yXQ7R8EOm+bVDezdeePHQCbBnaXtcTfzlbObJwuyIWsA5pI++
RYCIFg4w3EKjLgWmvJm43vBaRNJUiEGnVZeIlUX3Q/s+8N8992kqHdnHoiP+2TaStRy6CG4+gA01
RgiRP8xmtmSrpbthPlhk0+Obd0GwiXXk/ZOi27xTdUzn9NxlGQpk6zO3k5X/qTWAROE9D6UTCxLs
NCbud4ALjcaT5tXB3bKyMvK4UaGOkAaM2n5GpjXfF+dYr8jsZP1ptu+wFuibyXi+7FThqD/dnZtJ
2mrlXetiM9FeDX5WHwXZ11cf5LyV9p51Cqir4yNTRQAV/Vatt5zT5mSQXwlL2RGDK+AxCGRINB5n
O1U/xW/ABZZBGvfsyFzu9zZNctWHSbEFSYbER/DwvH0hWXHc8pjGLPKp1t5ISdglxGm+knZJJfNy
J3FuE1JW5+hZb/9hUhmkOmVgsgjNexMuHyX/8jyKIJKZxBIgPC3lPycCYO6LZlfL6VAAicIcKzVB
jMbNBVyC24/9VBpncSTBx6mvnJhag5kKNcKsX6w2VrcwMtA8yJQqqhoj1jhxqnqAqz6Vg+HbWqgu
aDpNLo+6DhRCSIdlYUJ6wrDyFWBz4aehJPo0+rEzKPwKfWIWO7PGRYX2hOnuwJPw8ms9K+e4guR1
0QvEBzJDqctKaK7t3tOF1MFGm98ACN4jYB83Clu1Zs+i3BQvAeD7+2vDft94I61TP7ZX7vyQ9rBh
PnFRpOaCaIZJ/b9jj4bBNN67Z4ki+NI2g8UqQrPYjudOV5oVfmT0ZoPk5QLqYMINSdc1bGyJK0w9
eik6Y8BD/O94fu+vsGfhtpZAvFq1CyMQponYCNKZVAQc4eeTNGxmzFJtWdZIluBgaRpRe+mEFbiG
BH3hspcazsknLQIkE1+617Fdx1LLJRpXdUHtg8Z8boHv+GkAtbtRCVycoTubbP3bgUPIsT6f5Vd3
vOoUYPNv768zIUZvyqxivja9WNsCpwYkUYRnlBfwV1ku5t71/PJQXG89HE94pyiJt81Iy4862CN3
mBL7bhhbeIlSWWf9YxEE0Q74SG6Rymbdjn/vRT22P8gSmh+uAE4C3FjZM3VJt5Sbi7LJ50G43kJn
t096e7PnPyrkrYRus/CX+InWQu0YEL027rWmYisd7TWH8fr2YjZ7XeI2ykrUUhmi4FCAC3pJboah
UYGBm6FRhiYrX/h06mO88P0wOkdc/ykQSCLmhMOGa3FD2YdNoJFxub9SX7iSxXBel52UBaosYv26
bYMbibb7JOYaiIkKxYCqrqpyA5RaddJ1y69+oRfK5GYD8gTh5WRsugI7zQPUVrprVRnJ5bioaTz0
eeFm1+dhoevb9O7AFLWL3GDT+yq6KkrnFaAT9/sgoAI4dsd9dcrUbrPMC6zuXBSFC52pParf7San
tgVwqzAa522LbMlF3bjrqF2ucZACGvik9uca3LJvHhMKh6JH5t8DQHwk0uiW0uSVq1iat/I44Uum
izZR2j4NM3tyzeIiXcW7R5eEOQS2trThu6WPywfgMGXVTDlozIMlXRMq1vOcJ3vcDeT/MJSeOIJ0
se4wzBYN5oFUXSVoRnjj7NUojUM/Rqv9qEx4zF5ZXxEAeOAsVJWD0fhntGnb3KOaWwX19/3QpLMt
l72dkbKdbYPmpIaSdiM4ErY0EBLD11QbWYmZDRGN2h63EL5/k+3/8gVLFnbNreAAnTER0DmMibiz
f3wTyC2wIQJMu1lZKCmJ59OIgJUfW3ovFfuv7QB2L0o7XkKlPM62Pu29UWmEm/dopZBWPzH67k4R
wttFhQ5qkNjYz9MiF9BDbFPKYVHos/SYXQBw+6nXCXB6GNER841m/C28Xyoak8g68plyB4+dYNtQ
jX/+Mow+WZfcMIxwdIef2Gbs22MXWkUIdoLgmO7m/KdwnVYsN8cljDT+3BiEuoGYLa102L6KF0Ez
rQqnFnzg6HKmMF7gVO2QJ6rV/sICVKC23YbvklfCwqS+y1BGBaBIza3h/FYQzZa1OWTpycg6c11l
LTu4SPAodp4UmpGLZuufugdogpspglragkEchDUGvEHhkDxIBc4NMX7255efU6X4gaHdeDNPtOaD
dP5hFQZM66lUmtq5g0nlZlLmlp2E9SRvvwsNReoZebXDO2rtIkF5r2oJhetK6j5ifCOq18GyS4+O
xq+QhnJHR49m+pB8wJU0xpmgF7Dp1LPX36JZKPOwOiyiMYLoqELRHSFg68Wf5Jj3ASXUBIih8R9m
j5qLMIM7BVDSVa7LOD9lab0AWTwahXs12yRIkjgR5MWz22TACjVyweBwDNMKeGieJZ1HctkBI+25
v8SVl+qijk3cXO2Ff3Z85xTxPeu3tmCs8b6eg/wjnYfeXonZCa6ghAuOKVJS/oWIMrNCFk0MoSwM
b2SWNyeKJIomBdCrClQ8+CC3zbnHq7/r0gvBAFuC7RuYhXidGDx7mUv1KuGaMQ/hRDEpUF0GpFp+
SFBXTOiNTMoRNNovyVKzULk1RugyNrbDSKTK31UuPfnBsqDfg63fo7+Z4YQcsdNmqds41Zycx+0E
iB20MVMCl+4L6IzIPJ2Ni71JhPHdj8JgMru+2f9B+pFlylfuZcL10WMFHMO6e3ab7aHWprraz4a7
58RpvNFKbhJjkPM1QXi77OXUiJfxAuABP5OOkqlG7n8ditSXMlvZtnEbOmoBdsANmXOgtqagtedR
H21koc70npPzn/Vpwhx+dZR+Z2fTDyw6Q2ta+b5DOoIg7MPHiqs3zscP0ExhY+0zkHX/2nvOAkOJ
Nw15i1WvOrrHdInbYdEwCPe+2N09hCjQHYy1arzONp/pWQ/ryM7f7x2A6239hjyqEDYCxPS75n98
uX3zUZ2eiCC4VnuieoXRhZZpVHN7kexRDOiBxH8bBigpUo+m9eZrQ2tB8rtJLGXvtSf4Y7qWdfqR
FRUZaWSz7fylNVuaUaWiuEGenM6Cv4jrPe4L8DjgG1lWd0B5FFsbK2auM0a89/YkJYfFeIveYz96
R5GWqRb1HsZ6bnxuH2ACok44/VsoDOvKpKCFDzaxKBQiari98cGcUiXhnp3apj7huDLlf28vzCw6
ot/ppw5ss10UxxS+lhHh9txN9+qZwR7PPLKJVIG6wRecjlnQnMYY3qgv6CypovPRCyWsm6XrHyiZ
EyYktLVYLY7ysmg9X4EAFac6zHoWLvaMOr41sTz3b4nub5a/+zK4+nDC0VnS9odcoe+QRny34beI
ZS2+MggQeklC37dt6K6Oo0rkegyEqy2SOQCtFN2bYu6YLcML1QM9jLfbqHqWlzeEItZp7yMLa33o
A5j4QomVipnvjEBc11tZeg9KvzchzO3/EtItpxO3Zp0DtI0BeQ4dl3ecKO8kt1f4PO7gvGejSG6Q
8se8GMnZ6IzxCUTd2VEO18YFjg3guXM4eIDxvZeyO8v97g9c9lDIqspdCWQLkQ8nZOlL+5VFvf3A
Zb6mjkK2cHRGnpyqmS6LN8Jd2kYFjx1FpWl6M3pbxQrf68gNLjbxOo4wraaVDQvkUYsISGAzCIvw
xHIHykB1fhFa6BywprmKQKefIHY45rs1J5vOHDdNHVYZDbo3mQduXp61t0KsVvACQT2+4M7jjyJL
yU13Pl29Jpv9tOdkvFjoz3E++1ZZfU91/ZenHlEoe6K8gDUeYU8VoovYI+ZvqFh1R70QV6+4xrIt
GOycpUvkmjXjbkzudyecQDF5QzViNRhF7KledEdFxreZUKtEepBxWsGOjbBmRKJxUvSB4zLIKxJ4
ZSy62tBfXtyhZjplkXuD0PBu1p532978tbAXVa7hRfp4o3nkGY0V4mZ59Z7NcjqsZQOvi307rrBS
yXDmc3nurEB8WTq95Os+Bhos6PciwMmGnCQzk1/F7xmUiKcpfSqw7kGkAOSoWfp26P5y9zSRvjQ6
q+sKEqwh6h5WRlrtg3tCQ0NysKTJHdY6mWNxX85V5+6xWzohK21FPV8/rgd+FMVaomCx0ugRZaa7
srAnGFtOJM0WEE40bZt/hmaD/bsI9SwjZ6lKZD6Ba27W5EV8bCgd4hrIqdW84yER6N77ls2xAyuz
mZq5tI6XImqfkYwKr0NdG2mHEflpdqWQNSQS+b68t0vttF7xon387n5+IHo4S5oR5fXIolJEiB2o
2HXzv0oA5LmfbY7/aVeg4eecC04oaiB2IYjEfjQIhDB9Kk1+fQ/IaRBJFwrWgSkqWGpt0hE2VqmR
3Fj7a3whelpYIRyw69Om1d5BNVe8v5vv1lb92wir/kkEWFI7E/iSq9uMFlQhP5N6iOVvhr0C8Ty3
1xeXjmLGJUVXdPq995KUsxIgE2KqnO7n3N9mTnqMJ9NucJOwYddr4x2Lneu+DI/WUMdul2y2ibq6
+pmm4J/IkEZL+PJI+5qL0H9jwyFO0u3epKgZe+wU/tfTBWNIRp7PovQbF8xx454TqKA4768XCxq/
S0rdLWnaGfwFhHnDEOOH2UdJLZXk7c5MpISBuTVMKKRgxvMqZNPCXnMxiPXHh4rCVwZkGSmTOy/t
SAdUV8YGqtO9ciSeTZOmbbrnNYIRIXOBElaT6EvFYL6uUmixz/UFjunJGi7DRkNx5vp2AbWr0cHo
Ry9+pfE6dkB/0zzNU2XVp+ofdDeN+NGoHXepjKwonIi1FRsK/dHESfX1FdRToZrC5dNNif0Mmkct
dzDCn8x/cx0kU32F0KLyuecRwPsNKRdF0A4BI95/bf4gDe0JYKM4u43C8NJ7CsboZFC4e+1PHDwi
stEPMdgTw/yZEK3D3qjDSNHWE396oO9sCQiWEYtsxp3p3dPqH/HuwTpJSThXmJdiztSctIdvzr7y
aKb0XDgczeSh6eWzLTCpg2163xjHoFS0PMo/WeioUfDkCUNZjIOdJEoYaPhBsT5rGZNFvY5kYHsg
NksCSJxsiJEf6pGY3gdsX29yg6RafM6YIFyk3ZSbeidWfDpp+HI9Us1ucTZ7KuK+VVzgGG4UpB0k
2L5TTK5a2t3VvtEf440TConXxEY6oEEC7Iy2EKMPfByggOcxKps8zUCb+qVI05Ghjopiq9Ug2IPE
sAeG2gtSmzhY25HYlswityVfUxzVS7SRkq/RR1Kqfmv4yLqWrh+nWlNBNv+ja7HXQH8yMfTMoaUn
8Ayx8uwAWTjPwgRrqLO8yeHReWwLoNrui5KyjhsSF0tknDLwQeZ2ESMNAaImJOdxUs0d6fvKcc1a
2T8LnPQRgdKjt+a5RxmiYTUqIgagnyYRv9ev4nr8YlYaZNEJooxTPjV0nXoVY2JcHfpC+AMYzqiT
/niyb9PQwmOAm+62GUmxFfWq37KFSrC5UjGmkbJC4sHCawpLCs9YAioOAyR3yNLKzREJG/HKAX6j
sCKbd/FIV8cdRlaYwSrzr52uhQcj4NbAHLUeqLon4nHvJLMYnQEEkx8InyYhex9E4eDzEJJ5UUb4
0eKeXA70yRLO0t3FuIty60SLr+z6MWOYYEbB/luT6yfhCt6Ogv5aL09aq14nVHdsMzNme9qlhmfz
Di+9de1ZBqBqSXGB/zNkiewy9vBKK2EUu1BtUk36Ctm/m7u87m0kEoyjMDETnxDweQmPPeQ1KlFZ
Zb+RA6s9BDPiHzFuT5IzxgB4PI31dQVJyBFam12GaekoKOHw46E8ebPn/a75q1a2mzQDOmfHvWEO
Uh+7CBcdfK6IS9VKN5xddWjHARBDW0x/toWxpQiE0cd2C3QUz8RASaDvfYoiSPHXytqZHsX/+dVk
zbV6vAuHCNEmUCwFGz9SJbZU55dVcsbkEYcXknle2ht3Yt1MM0Y/fz/nEMtMbX8gLRFMOriPbTDt
jUK/LrZPNOzj/FYcDB7jZDaOvXGHulAs2CkV3cP1M7FaeOJ/Dmqcjou0iDj9EZPAab9hJ4jMuyEE
6TVWnFynF3D0JAOGls7ipMcKg0oc0cRbUfGpWSUWDgZTC9IZ9sbqEOtTt+/1Rfd/x/ZblHvoIz4R
ctXpNJ+u56JpScwvLn5UrWMvXj8hsvTrkCeO7Zw/95y7WW/tNGkRNoc46olwY5F4bd5SvLAPAFtU
b9tHqbqksiR2DyHiykrfq/L5YHGdD0K8mGuizTbmETXzKtyo0XDKsAQhxBub0TlRDEa5pgITiQ53
bJL34S0ggcFGzyIzUntg7NvRlPsEO2R5Y2k/eQprjtWzMy9zSSVZOZ8bBmqjPsoA+9Tr8EQIqn79
jm5nrNG0RH8Q5qK+c7VnR3048CXMhSCiw6FEtWc3fHIdkMwgImMCx/FUhwU9LgUFZw4Far93yN7g
ZLbyprapPt5hkseSvpZEUL5LLU8ysVocHmAYUvLlnvGV5fEr+J0gduXQp5GbYvQBW329LaOziKRi
BqSRuqv5T3kP3WWm8PSZv+PXgx5qTAOF9k0dBrdtb/PK48ffelyf/uQHcfOxjqP6JbFLhzItN3D6
mP5UXg/rFJ8x4fc1e5aoTWO3NwrEDQRJ/y3XHewAFzeu7Sr2DePa+PTuxd6c1qvVUC/sajnkktJo
K2QZZ3y48LJhG/HGa8MkOgz4j6PPwwlk/6+LvTbpBItnuyCXkYOGx5YPCssA30pP/cBmkVAjGr4U
aXE0r5tkmff3suqCY8UFgPukwixbziSEkAT/rFofS10LANITEwl9WeLpH2Cpuykmzeb/cIFn3cdK
G3wVuKzy81mhkkx+rAQJ7ELbHqI5OtiFPln8FdTtyoZ4gXEAcpyvWND4d89e0HYDwwmv6JcLYj4B
ZT7gRmMrLQBjlQDUVsCbWsoSqE3z963saeAkfxkrn7hEI5rjOb5x5wr9e9RxtO+ayJiYdNw2FrC9
DxLFQdMJ2xDRueTkzA0zf7pFIOiNnBZaKvXxAVxpwlnuTw1rMGAWcs2Fjk7j76ISVjQioYVqNPXN
SdS07Uj0uMDoqgczUQfRjp2lS+8gDUzjcsG/wB3yugIFhn8jK4kBJceK/zKGuH6Sq1L1TIhwpKjm
YfEfq/o5GDAuNEc+juRkmQp9vCeA2h25N+dxlHl6NJQW13gLwc+IVz5t0ei3h/d/DDkcj++xHunq
+txiHpwhbqkdWaQd65J3dRIArdNlnERHV6opWFsMV6O1Wswp/oUneQdv8FRYNGyMDOVPgVIsJ32E
AEuhcGzEqj0RGQy30TdkwvhQCTQw8Wy+fcDLuaqB4L98NhKaTSVhSwR2+Sbw5J+lNPM4M0CpgFJF
mvMQ7eL2ypXgf5ANhwxBrMnzannXn2P63W3ef6i0WmEK5gzJOxvC6zmDascVoZXshJ5gzizH9EQ7
qPRJxxDrUUkU3GzBH2XJ6/mDsIQ5+o+fLUMaWqos79Yaz8oWeiOQwdSqKLk8L27tassf/cHnzDBG
Q/gUYdzAE4GYLsfV2we5N9h/DxMW+EGXGUepB1UgER4nNL2AnP4n2nuKCp1ylFbZ582v9McgWiT+
V+yZByh4wqqzEnEVv8bQM+yjfDCPWFGAl9JTK/I5AnlKZPxzOYwzPB3QrhtvFaEB3FiChbab7Exl
jMZWXqHSXXW0NNa3QOyvAg7LLvxhd3BfAOd9ufst6QmuqMYA+OE91mc+p3gw/SZiVltZsET/qBx/
UseYG2SmqfAnVSCenW13H0BWZrk46B7hAx+A9zFVvGq1SBJJtQSyKuBmwCtFVgpzmm0UWlo/KVR2
L5B9Wg4NgVgIUX1HQ5eBCM+bkFGwnThEizfQhKcd6cfI0iC3j06gOtqI7Ash1W3pk5zn2pa+q4j2
dIWQEm1Bkpys1yWnceONYRpSeFx6jEBKj6vv4KiUrSqhltsEREcUkKnXEgKf0UDnMMHoJRNE2z7o
R743Ec/cw2aeixMV7qeJ/Isy1t74DXrFWrMdNZ2lve0sPNt1ahaeYlTrlUaHS1vJ8dNIuSOgKZvq
6ZUlFiuhZ4i0kpH7RE1MJaRA7SDUu0PRaSpXJUqYFnRiYfw3iyNZ2KiuuOKljPNzQpc8zZSOFfrt
+YYXkP3q39bTSWE5ss7nCg8na39oprm4AgRzuitseVPZkvni+yXzaIAPtmSpeSq3TXiKJJh1O0Qa
Y721bxIVsJjabncNlGdjGS3Y2Oyq0NHoPQC7tHS/ZwlPK7FMdIldgzsFKSeyoLRRIkYwS2cK1CA8
djekyKxldKDAPF9GWTLAbmZXUhBnQUuoTaGAPa+rF4JKS3NXVDW5rOK5u0JZKm+hfD5gbDNJc4HO
tEpdcGwbBvPHRj49+cuBKC9gBIVdF9vVlq8kvtZwDITr8lNWQfEvtrkjk6Tw7MluzvMoahvHFqnR
ygl932Q0vn9rpF/p5h6N7WmVB7S6llhVb5iDL1fy70Q6cJMryDCc02v24U8UJFDPVV78HcCOa3oi
L+SYWX8M9KcfQ2hKRwzqAXEbNst7Df5njI4NG8LiZhUVgK4zxPo1eXFhh25tJJL4ArCZSmn5sAkf
2/YYnEMir4KQvpLrN2iqciP+0o8sPur5LxG2H1pPKkj00LktwSwzRhgNsOI7k8Bhj5v9fQAK1uud
1/bFC79B6oeJ11Xr9lCURtJmESn1es4oHThQrBCJUOrIhh92Xs/83fRKXmAkVBeHPblTple9Qj19
m1eISMWVn4nqz05z3zFsnETQU4F8AuqnpUYU9wcRlspXD1v2D0GGVXuw6qPZc0TkHa/fNbOWUZmg
BwYwMxgN9sMiRNETLPfI4X1bBixNDP2fpIox1wYstvSMztE32yCS7Reyj56GuAjpt0s5p4/EekV4
AzGnb8xxY8wXV8IZ1hx8qplOi2bMLnpD67YUcoa0TxkpYYbY6/Tm6KW6GBC3/Yn1kKAaWumbiKRT
tRcIbX8Nw26y43MLoKQmS8BBU3Pjfw52sExOE5EIaDYV6hrQGhz7e0bJhUWpnqGNARA5cY9ISCfV
fXYMmeMcX2K2x/Ayryl0S2H4GOJwK1uRATmZT+iSI+ewFUTX1BQDWT3cuOtlRdtaqxrHnjCQrGK9
g219ww7RsvMxA+XbISXRBJCJeWrQIBiJ0/wt8MokpinMmFV8qKZkq6uwwjinRFDw4NgCrF6Q6/lW
SuvbCEFss/WYUsY80qisO72VWOsVoZ2aeK4UzOzBrhitTIVSiWGcXr2LhJlOwRtIpZp1Krb3mMqS
R0Sz7hHN2z6L3CijtAC5KGvmG8ZI9i+GT62gzgNqxBXMnl2OA7/zyYnOicO39YqznWFv/GrEK/+0
nlG09amL90FWtbL2bsae8C76I3KYwBTKS/quDMB9f3OP2oOAmpH989X6oGxpwln5GPMyMEW+qSBf
p546uMAfwnCgJvQk5GLJlKdl3V7bmJ5cpCjzsApwEVgGk9aEkOwasZ5K8FfVCBk5CxrV9NsISs+z
FFeKOptU2ivKxL1hwofMCZjRM88tcbv2MfrN2DZVe/5ZO5CPsj/DYv8yVcnJJFlVWsyGWWNm4A5g
9KxSGrdlkoqQeNhm6ezIyZV6Vi3fCVPPQMVUggufKAdqNepMIKpBC0pfVlHL3avnPJ7G/rMOBeep
YpFPdwUr0P918Dlbd+5fHAazyqBqpB5pUnzF8t94ZN/+kQa+iPGKDY/UcO1cKsXv3r8kTUF63H2t
B3KrbviVvJthgn97rsoqOptY8OZHwx3UglAbxw9Xh/RwVj6SLe8Q9iRyifXOv9cszuvXI8RHnz2y
RBo5n9kQVByvRhviZ69BG1LK5fo4YJdpvXH9rAyTU0z2MhqVZgSGZBd502Zf/DNyEvY50prEuDko
uwrMi3rRvLT0yXEcll5YbAzsuKD42t39j8GZF74atM9j7gXvlnxqxm/XhujBfHr8fsE0XAJDINM4
2vywX59QaLq9wIyKy3mHwYnS9MdLsNHk12yqBatVtHwbPIFRadqb9S7AXCKhmMrtg0fUwVhQlk2G
PeXVx2qkfHELoeOfYuo0dyTT+NR/Djt1/e8bquq85CUPvpsG0XkOt6NjiprmLYLoT60vIAC9ESXl
VIrhKfW6wJ+V6KzCqDnCCcwyIcT+1DktJqY9B0h/Hi30rlHwhegezZjN3oial4I5NOgu4FxQTImb
AnFn1TaLIgxOhErJuqHzYxriVYYpbXaoVRpT4sQXWGNOxaL/D6hByOraLgeyWk4EAwhwY9TX2fu5
EwciZ5xIbZ0Dl6pkzQDqV//FdwG9FkYd2W7c3Q5MEuGDATikbVzzyys8BnyRMoz8zYqMaWmXiQ2U
1ufeNfjihMYHVj5iDmH4phS8bLub+L3597vya0UkNMn1A9g1IqIGjLIPjExj2KksRGLbSxhYa1lM
BC6AROxbGzOj6IYiuEcPydQoMbBrHGDxTqYtxWZBu2JMCmpz1w4rUIW5tI0i5QiGydsFVkPMz3bB
I2AqR+g+yUUfvSycWL/BpWTq8x4Qx9Jw5tiKDQ9M1VmuY95xHsgcdqsqj4pxeieiN/mlQW3TICmR
WyCIHcAfCxe5ADLVTLrHIVQ/pwfhXvvJXcPYddPqJWmyyzzmMOVwxCyW3x7d/c8U+kqM2/S4QMLd
QtSYeOYcpTARwPbVkRnG9CyWQG19AvYjHDie0rzB2BQqxtE1CpTJ9DXR44o6PBgQasldoS2By7UO
0ZkuF9O9MdM/U2hfKMXWat9CDuVrOfNhBegOaAowuhiCmFPKlJ+jSLi+pRqYBCqd6NDjW4Aql/hd
HosVGWjHFtxQY28RaA+YxwNt5k4cL61AWSWX/+a89nVZofGZtkp3yJ28Op7iiZtsm+3zLPGxSip6
9yM60BVJJrJHZQveDOyNIpnJwrlEnuBDvHMpcsHcGHldBK63ZnctOCKicZkzg8LsQbpws3QlAGKp
69dnx0GxfRG2qB9/YkYx4FDHar4aTtTFwA+4USq7i+53t2RqLWRHl641QQWjzoRGBr0jNGtcMKkb
DeEcKbyELv7dELOjdbZl0wOY53ELZypg/Txwa1JXOcnY4FeguNcQGxY7BlX86EuOGdHq14CCBO41
xW1gj24aylUPeA3Cv5QNOa8ucWOT4eHKoH9tKVHMGXJAz73Y6IyibZbgZia00Cm/cfSh6VnAKRJY
nuyEcZ/If6ab1U+8uiDHobERbRkE2swrb+OSdl/2NtYZe7DXm2o4mI6S5107kqIrJnnyhQC0tYvY
Mg2txVY5EQ61rQ8rqUiD3TfPon8iyW9YYEjv8oubiD+93UY805iXx/ICUGQHUt4g5I/DWPs7ziGA
wKhRELpgKNrSwuXA5sGuXISqLCBhjfpH3CfPODFY5rz0pXN+CBLNW5kwXMC10Pz1KpXLrk1WZTYv
8yhwWGNjdYH6Ps9TQzoHyfFeVTIPofyLDn8TyxRtz/Iahiw6FJCxtQoPboV6JnKpfbx3p7IP5OAC
CfwY1EHBBpL4BIKci2fqG/eAkiAO8M1T8qino5lZnOPtJHk5WBRJB/cWtR7x+kvKKIneExjF9CmZ
jMcu97IabCAsWAz1SIF+fLs2KGjN59xB5+1T1Te9StF/FDMlV+ydYzuFWNeLKDlG/01bXjfgEKB7
+jrWkd4pKhVAQ2e/CCAgJq864TP+N3k1eiYv/uJ454OCInIpAXDUUnR8eqsTwmbnZOj4ZBiMcjNL
iZfXFUDYf5CFlamQnwcHmxCXPZGLNPUU2bT6sgMwc7oCGAWNjrV3HcD80OXHZK6mi31nJJWFNIjd
Ydf7PwvQdNK2ionOa7/yLfTbcJUvhDK7d1FrhWOFMT+Xlju8+4v4wwDLApRGuMxtdsfXKkhLErta
ehZDl+yBfKav8l3f/naejjpUNy2GR8QLhdIPK/T/HJatZEndXfS5K8eY+lV2Ya2L2EsWZrZsYx1T
+OKJSApI5iATkHm1iee6BkSZShugxI9XwQSRxWviPXUkq+ZfjAOkXEovC9am8U+Zqp+rSqJzm/zb
O8eGbSxc4jwRFGcjD5ibP/4jL/s7Ol8HZjBdAJFt0a2Rg+DxyH8vJpCiz3VtnOYEfRIUrgU2brN/
a4l9vuDV0xe5oIHgpe1kGGEUbd2NwftoLC0Xvob6+772yLUiPeUzQHDE0nCpqYVXKK0o+3ysJOUD
1IMbVos6FoM2wwB0oS7o+vyWhEo9qkNbrTYp6CTptcc8OdZhD1epO4eU07Y9KbvxBd1YCwNK9S3J
saeL2EVDAGucDHT4aecQIHNexEghXlYAepx20fkrcA4+THLee5oHd4L/yY8YB4YC7qBqC7OoBhWJ
JmLAjIpHkzwHptzm9370NrLGzleQ8TA1ygSqQjbeHScH84HoMul8PXuJD9T+AWR5kq/PEllRKGqP
o6LxD4UQmwK+c9KUJv6oJmMA8l0LI6MmHn+UtXuANKoWXmPV9d+cnB3VPOVCGzOa851JvyROSLed
WOl3dcOqRX/KaCoKpwMoJ4kcSatGxq3RYIePVRoFNgFPrDuROBqbIc8oVN234moKf1UBdRijG82C
Ovs+bNu6Hr4klVcv9vbtH5p0QbEv4VPQtDPO/r5i5xFWwEO1i9C6iQrsuUFslHhDAEEyFGZvvJED
ubZhim4x88MsK8opwPa5EoJB8SHsmmCVcTSrH5gh6z7no/BGVW175gwuS882hCUaouzfIl6JvxYy
BLD71EgTc0McFb6Q/9pg+ZOE64kCENM136KvJu7EK71KS6npA7Fsimqu+MUpGLB099w+ifGyjS1M
lybSpCI0hLOnvBj0f9GZMGMHoyMjqgacMQevM3HUzdcdv8FW2l5ADqiEygYbPUC9a1ytSTBvCykT
8irgHg9HGixGsyJB9K2Jk4i1S5wNzVdSbokdhGEO/y/MIwBl2L+2XJa6DiyHOtOHX/bQVN+aiMzl
6W12v8O/OqIkh4ONz1lFuGHNoY8BQPc7fOq4rGvxWKMxy4mu/HraFxpQK/V/VDKic4NR4DlI9Pz3
x2nsXO+CwhWHvOA3ck/JXXI+0wY2Mr38LP0pVG0KYXSWIVI92kvUR0xFttFxy8BrYRUw4Y1D4V9p
21WLm0vzeDUYV7tuqHxt9WMAZU6nGzXCYUl5/fV9Zd2zIYiwd6k1iRfoqO/qJ43LSZ1XzgEFsU9p
GrDFpGwWBfG/4PENukEZch79Vm6tMVpmESwOhucoLTRnfqXsFUkhxSOkmwcwg4Tsj8G/12IlIxcp
3dXU7d18fJLPEnLRN6fVu1bXZxBgaST7YvSM0brm5E0YiEqDoMfmbX8Ar8Y/Rz9zNcTmEKxt6f64
sPBP15DQf4+LScqsdG3pmonCT1u+m2icEoufjUMBdoqtVLF6uKeFQRS9W+DZFsmwW931YgTP4g6i
l9ivX0pl+D6kU1fuwnge4gX1vLmKkERGoiE17dwATO74Ra3V77jmOFtbO/GWsP7qSE/J7rLbQe6W
J6tPNfCR+W64caWJvlSzQ0zrWgQAHsQvGpsZH+jS8FKLIWaJZAfhacMA1idcv+JeXEiswlaso5Ac
gOESr1esEtze8ClyLRIaS8WDP0EPW1DeAm6IzdtjA/tiuRxgLegP8qFb5DR+sQ/NvOrgKKdqXgny
DMq+bsXTlZWz1lmHmfNpUMIZxCnpC1DrMYhHphzALRkF2bK6vEtXjHRIdWaSDczA6WaOlh8ckgX9
4IOzX6sRcLp8ajzAXuf/4J5AW3HZ/rE2+XRunifntPYZC9uTQIOnRgMxklVlBctVOFKsxUsD8EDa
OS9UxBUTVCgkUItZFYANbk7cKKhvzbwt4rn15MKed9BBfg9FzL4hzPCoQ2fVwgUw3QycRnSBpRnk
y0FJimoyhSdjz2bABP1MHonr7n+wUc4Llir1/2sHNVg6+rNAOK/3xABC3coqxOhD5UAdmrvlKSTz
mfFwLvTehamOsrn8krML9vqZ074HJDqGKt/Yn62tn+TLoYqnT+yh8xwAwFIyljuDAsrnWN2VLr0l
sIXGwIawGYT3PmoVPy0PEqwY9D1VA1Q/7fu8xJvrm1rug20tbx29L2pWXQCcJTSziGjIbfJo6O41
QgjJCE1mQi+UfSdI6VxjvV7RuXDDluK7pHv3Ee34dg8SjOWGJ0jcM/vlGxWrzYvsSVV67P1k8rRu
ZAWrp2Uze0fxyuvQzXX4aonMWwd92xy5eCxTl2vkvIXVIcWkXsJ3p/ORaCCzjhnIjDQXYRxdAIkG
BlkRz5bLfdumBUE7afwxFMCVgEwuv8oAqPzjtW8E8cBGJy89L9rBj5eOkdi7Ev5i+bE4rlIyCjXM
olwAFTksjhaVF4ush46eBqGw1bJVALolFn9gGyP1zPhF7qVS62OM+RqbDXvjc5dJQTgKNp8OlzuY
QWFSVrwril4ToJIg9NNl7z6oCLytsPN5BLoWAMhsTDZYr0UJDYc1635g4y8iuCS1guBtCYKnUQNb
yp3g8XWPUpuAp69cHn0PEIYCFxaZLDmqf5+e/4qw0r7x4uSlYUnHuJ0GQ7us0KD7Cg80EDGBhQaO
sXF7BWABKGpYKtNi59wg63ZM8xy5xN/oGSK4KpxoruI+xZZ6s7a5pVFoopk4dWT3iKNpZVyTbp4N
puay7pizERcVKf9kghBAGiDi1snM4xxfmWny1NNSdWR0UEiCYASTy9J3wNGHEMqJZfh/XgZs+kf7
coG96jMeq85WHgaRe1+h5mew7IyMUGZ4XpKk99tmlBpgcgE3bkmXUXRfdsu9JihxJzBjxE/6qnlt
xB347n0uEih05JzmO/dCty5ecRTCodLcdrueow3EVav6xsu79K8ddjQTmYselVPKb2K5RqSrhsQT
u6LWRKKN+ZHk2Y5azCd3EbeqDkpc76h+H9ZUdPaW9hY2CRn/jk8tJoveV8K3RvQThf/oMvYGKbTE
pAjItUKjLF0fU0e6gmxWRFjioLpRh2/oCz5suUOOXieTGQsGvJ8fR+OLIeDdpv+6Av7cffb0voYK
sWay9HvBx6T8A6QP2FVSyfT835OsqN1oEumy439NHjpJvGdMmPIOJLaZaPV+PvEomvKdC0wO2pwb
gNC+KyK/iwaNg3zYEFD1nIusnVv0vlnFSkPJKbJTB2RLdz/Kjbds8MqUnI3wFJ1BZthI1ayvrnd4
ephUCNF/jhCVfGP6HyioKeVWLT4IlFMZ+q0OBRxMt6ifmwgexoNYnvjxAHiQMTNMLD0aHRdP9rty
sO2i+Ra9o+jyXuZ+Hs5mlsV5sYj3Jou4JvuR8vTarKko1Gmd29+Fux4htFglTOupGC9qt4vwJMTU
7RwTW3y+VPnoifcmlr+N0NJoXz3lQ/Fn2XEHEsK5as7SkXHVWQIauK1AYm3kO8M7hHxal22LiGfP
k4g1DPf7XMzrK4mS1vYZyPrEgDvjV3P9whZxCauLp+FXE6qOxjiMpgO3LlYkyPQya1GwR5J/N6rZ
TVlhFuU3xYyarl6iB725cXbiomrIEbLc7CiWLT+VTy+6CuacD25nUSB5e6x4Dw5vhUwkwF5pNhlT
1Rb4k2n8bvtzpDtaLBJfp8MTIJAMm98MP7ZGYylwijN+9QhYgl0g7ZMdsYJBouWLQkS7CxDWbHjo
wRjp7OIxrgIMWyA9cT5Yd+M+9i/NIdITVLYZr6GHa+dwaegVeWiqwYC8Lul5dXGThs88kXbgMTN4
z0ccA2Y0w0bH7M/x9ZEJ/BXXhOuVEdxgZbLUP7juHL7fjBF8mJuQwcpSfusPFXmewSb5Gd1tZYQc
MV2dZInRgQTNJVry9B0B3saiu/33NiARE+RghqfOHcFHrcJAVjTtuRb8fAO8AY4c7iKBhSNi2dpV
pK0tPJ3Xb0clapikT5m7/3DrBaHnF26+OjbhW6IJqq/PO5TCDZg7c1hX170IMraqGv8a65+Jpxm8
wIkUtV6QMclI7VKdfxA0ekzC6O0H3qogdXtI7dDHQWviPoVTGoEzBw6/Q5MMsWsKHdWOV2Oi9pyq
0n1+yYrL+zu628DZXNF/wKPxNV3Kpp0lNWv/FxI/wWS0LLfo9ooPq8l/k6UBqd7zODD08W07/Dsy
itBYXWerb5z32Uf7jE2bp/ohncB7EgXs7xN22tmiEWPObvtmJL0+HtyRfSyWgil1jM3jgdJgGSOa
sRvNrCLO4m/CK6KW0iBdh7LeH4VbeL/I6h2hpxHEvCowyh6zIk7UgrsAznCCOGoEQYBA4nrm5KC8
bgpnkKpm5ZJpmGzXcOKapRYlxJFVqNvu4DKC2AdnkBLQiF+LPf7x49ICR95OWr73PgjVrmMQwPJx
BJtzEoKj6BvsJ3uFzx4AzOCPd95cw2oc4HaElhvHFFFIoqTrO98aJdKi4RMBEhQbZr8AkW9crdyy
T71/VZFWJl2URXBsZ9cAU/OHIRTugN3ChofJa3djGALv2vtVMx/3gX3W0vp/W/wo9Jegfgd/WShn
E2eR+haZNMyKoSyGN/VVMQwAI64t7N0NRGQ+NrwEB7NzD6zgJgYOTSaJA4VtvQvRvPEosQm57Kf2
dMqeFOMdDO04KtIT5TYEr7khcQRzS0Vf12pv8pWa69uf/4dwsYOz6MtRUQoKhlgCSdLNqbtRPCoN
+dX2fGEErp7H5XQlo9sOKarg9jlhLzbGLGl/EATXZR376idoEh92RnFPz6Y7zunwwbf36q+flV7c
PSknc1hFnq9ETjNBKg++8I1byIqZnlVEz7MokjZzwS/2EoNstGJZGQ30dawbmtNOBYaY9wQ+DNB4
LbXCMWG0upCtW9zURJT+8GCoX2CJ0thNjLT4g+hRnwIyl5Yge+Ilw0IUy9PqWfKLbhLbsPNmXi7m
A/+vNG54IfPqAfC34SPfpvOuhK9kDWcUcJnCmDyQ0tdFb5dJMSevnG6Nr0PQ+9IAOwLHvHlMwh9s
cT2tIR0w29Y4Ov9VZRfJQd1rb8Aa73QNCjVG+DCg/RMix9ymlkes+WP7Ht9l7pwip5m+3CgomMV7
yqdSpwRXmBbndGKjxJZd7PKd1NBwyEEyBxewVSr6avXxi7VlBw2XSaPMt9wJgtlBHOrdVt4aBcJ9
BfLuzIfuvFrQQd75Xd7d/aBZqAWngTbg1V1bA5H8v593ADez/gPHbm9PhaDUUfmr4HgXZrKp6ski
x1yMrUg/OaF+cFOLSHr/dnv3C80FlwPYGH5yml81lm7qjUIQe9z2BX/GG67jKnZcgbYeKKwvXmMV
dgRZY8/S2vS0XI2pbcjtNcHg1vIcPJ6IQ0KmbP4fvAiFjq1jAABSB4xFDXrC1O0TqrSKDaEr2JOw
4LiHGCG1AZUs2YeTklEQGwLM9NV1beWV0jPuea2FTNaFHzCvyyNZRASxGG04ekwUgHqMrj9vAF8g
eEXvjLh0+xFIUrZhO03cxnqb+R5zh/XiQAPorqMW0ZGxrzjFxhjRb7Xe74tM8nzyE56X6ShhiapZ
974Wi4KM+fH0CmGoYvozdWRWY5wEVluHckJ8mXpJOFvMSv98OtBowB2lBG0/rKdRIQOhfdKSs9uD
vyPvsOy1eDyp/87D+M2qZKRs8iPWxjhk80v5HMO+3JCOCKhDkgqs/CZuOIzE/sseFt/R1yiaLHwT
4Kl2o7bs7hoiUiNgO2kvxN/DLXxCQZ7REWr5GwpqjLYDHYbhPYn+ZpGKPjbBPmIoP8+6DGJ+Hy1X
49nUPNKq/BhTuaDwEP2N8aICqgAw0pLrKruiYTkuM7el40a0FoXfNgfbdstl9PUH5uOwOXCoubu9
WicLRMqPrdpJvGTA9I9pSflZtaOsFhJ3rtyU+4UuMtCwRCgBZOBegpJa+VIPCSnJ+zjYt/ZHaZd1
HVH+drGh1Ev5b7XbkoomiVqVLjz8jcLXPfxOTEB9Oo8T8KZEvckPkryBkwx+HkVlyQ6lCMTFBKQQ
I/CHjuf0t7Nf4XBsT82YezJeha0unPW55/BehvcNi2I/fP9Uh7wURkmKxiHVqRdVUx/CXHnfMDrl
DMG4DN3Fh/DK8F1h5Xkozp7hWbkOIFtnqECtmrDaAtHyJf1lzuMpRKpsBh8TBwlRbwY8cCh4DCTx
wy+jhnG9woC/3g19EBw1hAbmQ2oiZkJH10Iduia7Yl1e/Xjj9yIEgmskDa1VB1POllhtlipC2n0I
OSIiJN8thBw3r5uPy2v+gQgRfnF56MFWxmyaBJWjwGhKSjq8KGwOfY2lxSPvCtqaGJEOHsbqrA9J
p2oOIdcq1IyIFcoA4uUF+7ccczXLoxM5tFt6MPnvBx/pU+ryzj6jWVYbUXPl8vNj/6+b6E47JGJm
04d3vzRg5s/9jmuFN0pZGyo1arv+5XNGkbZIxup6PRXtGhtR1TImjbhN0Nx1TsJne/5Wp2mgs7/d
jKoY+2RHw9R7aIw/sQbfCd5phPD74Vu5Vw7cky0lp85onVvwH8I4WNmTDQidEkRlc4HDO2mXR5Yu
WqxkSYWpQMlXuw3Lr+xIvnBPho0KIvVgfqRe2CPsH3Vz0pfK5cVpgcSDNdV/MBPJRYAa1za1EAnt
9MiPbBEsJIYPpIQvJTjw+0Vs1G8Gk/koQqfjRpksQG4GrO2wXv6DUlp0CXAQSA5p4ld+lgO4CLl5
+NfMAJ1Lsw+EZ+9rx+BX3sBVrvZxCSdSmwc2A3VVm39p3mLGBO16CLJrJnRXBAmgq3DYm0UNqsdm
h70wtCjfZbw0OlogPC2fs4Owv27JUvmhaOuzqztA9cixdtksuAyOiGuhOIxVtvWkgvAbBKn9K2R9
mJMHiQylVz3Gb89k2Hg4tpzGAJR3LT6LovjMbdAMGbvnkE2SH7CMMs4RWer2NYSeQGa71sCFNUeH
0rjB6KPn/FpU8Zn1R5lMe+0hZXe/Siu8xX26BThFi9B4wz5NvozyRygUPMO5Gf1QlDApheCmW1yU
h79MILbwOiwwry7fpyvFNGV2lvFLLuPrvSK5e7LAqthc72X0zp80N/NV5kW6mD7WPmcN5hSaQc2D
OKMgISZKxVNmte0ZPnVn72z8EbZ1ddUhuMceb1l+Wb0fitKAxnoNoN8R39kSybPem0MVJcwGMmjQ
JQ2yMnLmjlKfkP/WHh+cjD4Neh5CQ9czFhD1MZf0RA/SXyoM0BxXsdoMihLP7krxNrBnfECL92AT
sMN6Z868wZF/bou9ARXMhWzFKweiTfev8X46/TE5Oond8uXS9IaEfUPQZL9s7w79tDi6lq3xZ3bl
BarDRYM0MtSe4ucSQ12CL+IyTjp0Ry1HLZ8K7+Yn1wd6Z+9hrwtU6C90B8oXfpeYXOTRG0x+Kd6z
+/lHMeP+9z9GYMdN6XY5zAKOTcIb0omWcfBOD7gIfWr3vRnDCZz17ngQfnYkk0A9Ync3MOj+IcWB
UGnMXCehayovJneguuOeZlbVBhtekD2VB9WR0yleOUfdDV5Du4WsulLruzb2Roob5N6K60aZXrwS
907JPoXPDzYhWuAHiweBi1Wi/a/wQzKf5Ixrz8ohwqX0Bxc13WDdIs4EDSSBCcsE7WopokNV1WfC
xygzbhWYy/Ofmb2dB8HhXfjwICHGhBQMxMaY6FRn/9lWxKdyPu8IigGOJXHsePKGtPlXAdZ0sBsM
ZpyCcoeZ5Ns9JOTpLRJzQoGltCgaFyC9lhdJvAbSL2q9SKmm3Wwp3QSbpl7lB6n5TEbEY0KLPmno
rMdjg+iPYDrIfRncrZK8S0T7KwuhazvhHnkW49mwa+cc2dCEpIIgoEByKHlNceTIvWX6Vmd1xMP+
/UECsNH69GJNAXSqVZNG3r4R2I+Aa4B2rtu03i1JgPZqZ43wcgy8nP4SPxo5ATrIUx3albAIBqkF
ICA2BZr/4ARBmz03UqeLsE2aZHidqejWIVCB6mUjThkX42NvFHDQw3gfbEVrVFKFQbNI8ZGQILCL
Ex3YZtqnus8EQIxueEFnhr1TcErfeZ+366b39PniFtvQPemsJUSwyaT2/K/NvehpFJYrPqVTWOed
Tz8nTCjlxJKjFyuGQbai/sN2lj3XxmVZf4W+A5ThOKWgb6pHb11JRQ5LRcWPFDI/dGm+udOiGnHb
Rzn0eNRF5V5liyPLvzH9EzNLbOa2x5/vFPiYp0bFLV/0kaIqhDgtaeFYH7cnO3SvnBcgRBhiDNXk
UgLe2quYhE+PcAqfyJnhLZErNkrrlr3zXzvxD++aqjRm57ZCkyTa+mmNEpg1KnUuzrapfkUsoxXL
YvXLAk4XC1qVv5KI0KDeZAF6b8ZVuXLwHK2Jj4xa/3Mw3HKBTLgMf48QLscLfM/GRAwiOOBXOcH2
KXA4b8hwJY8i+OkYFqfLzwkL2AT1Td0QjVnKuVjo0s9Kh95pq1evbaUuYuYbGuj7Kn5kYID4TFl2
SvEKBjKwICAQ73nNbG0OMs2lLnwG94/rym01ocBotcV9V7iM4DB5v//Ysl9w8xiyMa6WuyO7MFwV
6IgGAhcNcMxNUoQxaDcCVRILPdfKhNl9AXFpNJ+4f4djrr2QYZAV3bHfEpIxGoyFOG07T3RYU9GU
CkyTlXrdZPb5S+zZHz7qSuMjgQv+tIBpr2/K8VSZP+5/CIHDkE/Yenz1iaJRiknipr5oMmrhFeFk
uXRLXtVl1HDIGQD+dNTIYC7mVJ+eVKNMkFealMDt7mo5edIh/IfNh+4tVpsFpqRmfskR10a+A3y+
uaZZtXFhXmk/PX+QL3GrW70WzP0M2i/OiyvrY/7MFINnSA+3TZtNdqx3JaWNVICezmIXGUusf/Ht
GrN+URCVSaQPBHHj9orZuuRdU3/TSJgVZGr0BqVniwKEINgEDAY6XC2GmiTEcQLGHm0iUw1JKUPa
ukaBLw5TEP0RJkeXD9UjauP6LkdvffQhAkZmlu52tYWowHiRzfH0MvQlalp36Kqob2bq22R6LHVs
++W56cGIox8+UhoY1E1WuJO56wGgZ7qYBsZHIfJy2szXH0ktG9XNBWKRr4Y6+iPqdeOUeQUc+9fL
eW1HaGPYEOljxs8Yp5M/mLE9I45KdLOIVSlKlR3BUEHVwaTZB6suqiwJ6SMLOI/jDqXyfSz/Dech
ZjSTzEe2CQbXvjS2oIK+SYPKxWRNjhs/fx1rII0oOTDX+kYy5Iql/KCA51ldtb+up/3rbmyOSlqZ
Z1WTqDAFAO3wRscCePbENXOTKiulL7XWl465/uwg4TO0v6xmCkbyB+6lkhiTAWFwvNliAe0nD5JN
mmHNqHWgchyRvi7YTmksVxhXuhuNDIE/Xb9esj/ay+Wq1f/p3N5z1gyr3VWHnsM5RW56uAv5uvO1
6vJjaLWvLSKpxupYyvTz7X0wSEeYnST4WENyA0i4WNWBCkFIRu7OFHrvQ4yeTE8EIh7cLCZy71B5
QMiMhFQH4weNywXe81d/mNxWzwUktZDhyAr1NvYkBrI10hWni+1wXiwgGnNLra6G3g71v/vOi3gC
aXzRFTyGskYadU5KSTZOYUGpKaRFAg6LgzBT0Y46lAGkFYjI3RlPO6GNeBLdMb4W4u9mKlTlXP8S
AvIKmSthj0I98dYLL9xNoT1+5dLEVS6qyqPiu3uEvXf18osJBcqeDu529TEo1GJNiZ5XXyenftlJ
pfMuXO9oissQqnZrF46hREd0qHNdXFOewWCEhmURSlkU7sCIIZzMu88O1AnnqfBmn9RtGHwQSRn1
nQO8Pnw95XWEdlJhKOGZY619m4hXncCZ47T670FO+aWY19Bu44ggN6KF9GbVeQTK0U2mD7GoHB/R
FR8i+wXis09XEbgL5WdFQLeisy0jcwaTfi9/wCznVqlPO0GqH4Ze7kgXEgMjrg/iW2RwsdkqFjH3
d5SrvK9U0uc8IaM081BdyoZizMCb3upMQz7PXx0tkKWGMjU+iOo2aghzVEVKC2ISDMwnnWASLaUa
ej6rz8ZZdH7ujWsCsnNrt9GPP7r3lSw5B9kEGqXJBNXOvJvwsBs1156fjLxDajw3TDOvrIFu0s0y
Enyz7PTGHrkfvO1Uuum4Y4H4+KANOktmBmrQJLBHWuXB84AFzbEblnnG1nq2QIiLnmzZJeKm790U
BUeXR9H4poGNue+M56LUQpm8GdEjECqJzu3w9bTy7XtG5U5z8AalbIz/sTDlFkChkA0ITdF8I9pK
TtlXBzGEhO1IKRL1pjxJwVgGWVd8JjzKTWjWjo18bVYLH5f4eU6XWYJoPETiCRryWaXeqY+MhKzW
GNJKWtMsMIU8rAgoC+ZUQYNDHFLT/bW1ne3W44g1ZBtPtiI0aMNvL/QWYpK14xu92SUd13teciFg
bqtjJRgaJgjKYBJiqPKtxsxGSU4KlGn97oixFzJutFWoPxYhd7pBYMLlovuhYg9TZOpArSJV32vW
JQXX3mu+46LhnlvVlX7NicHO/vvhwe3vO6DYOe1pFPraxGz/rvKWoijDYitSk1YIBOfJhqAYkHOf
DOH9ie9EpXozt3WwwaTnzQuw0MndSBTo6WwrLq05wzwrsHYmtjdaJQfBUMQPDuxM/wi77+6wTpnb
7L0HQK8BQ1FYNZJ1OpOXI49iKDdip6rDrCZ47X3T9/0zI/YX0Iv9jFQYWrBM0NE7fjHqF3/COvJw
mNOzYEm3XULEDMrWJ38pJ12W8BpOclyElrojIwCkaLT6Jyf/VeIBDNEAKuoCGk9Q5brkcocld3h+
9BV/ixuWGO9p825zTLghZHvbYktWhfKLHveQiZ5t+uwLX/J4PwpcN6SeXz9K3TrxI/AVU3fPYPd4
9xYQdjs5Utz0hGAAaNLE9RXi2amRTjNC5uaHKFRgmcgmcqH632nh1ZUBc3DMAadzLz1TGpmlHkvh
nHDjlMZNhPjeBZtbYwBJiOyB5eswazZXjg/i088zo0K8zJDIkdrbOWc2QFoxRqmTW43zaP2g/ywe
feoddTNxbeY7VO10tecgnfQY+aK9wC0+kRLfIZyD7LQaP6gLovQt9YsKSX3RZ5etTIvw2Y1J75EV
7E2/Ri7++dOuPFHPzlnexmp6LryBF8YfRa+wK8YF/PbE3FJ+fb+IR/5vSk8a9zAHgoUBfu3EqofX
Z/oCloTVLB6j9KjlpDue7MS4xS45L+qhmXuECQRxfjq9cGZZ1AHCELMWrPVSCPPZfXWGa02ZyAUf
KhUIlD8wHGinQtLt1vrm33h+RrxfRSiRiHAVS+IHtMhFJgUnecZxsM/C/0qtfMeTjVkqhuAhfKgh
CYmmAEXrRnNdSMwFb7c4bH2of8ji6WV9VX0EgLwpI2eVjqPFwO/EJKlYeWOAtmqXyGW7yKhGPRWR
nsOFkrDx5IGuVgbqthtQQ2ZuVLfxJWLFdOc/sIE1CTiMvw3DfuWcxFCRfQBHCn5Se1RtbnjVNoov
YIctzewqrdp4SWfBU5qhWkaznAOV9s97MmFCWJ2SoDmREliIN/M1UYFelq8uyl8aVAKCaNpFRGvd
8S/40Zh6PQVKCZ3LurxY/JSuM7ZXXxO7e1hhnDJB6ykHyqA6zuKusqE9fwob0rvZ3apEPvnDNJdd
jWsf6zuTHc7OiSpjl7+fmsIvB9VG4giA7WmXx5YfIH6jB+B27nLX5xt2pxcQWrFxDIwATzWByzjy
I+N//GCzMjM+IVhq0Gz0gYsdpQ4SzqGIdYD/jUModX9g9Amg7secYuzg/gmfCVG3h5NaiaMS0oKN
VvZSu5O7luLNo8d0Qh7ie4XpcB+M+A1GzpCBfidAAPaXUWs0yRNSEJyJx1ceqzLfxjchHo8oi/j7
6Hutc0siaYiq5QmQrl1hAxiQXxgG4CoGRrT00Pz0p6CBTU/9uze2Ntcl5f6MyUhYMNKio5fs7cdh
9rygtoY0tu+Ce0p79/ShsiJHTXVXdU0Y8jWVf/wutr7RGoTdYRH4HkzmSap5c00xbikkYS2HsLzf
i+GbFAT98adNFEwoHe3mqzxFwpTmvx0lXV6lqjdirtO/Xin67qFHXJmrbVl7Pv4vEhvDA16oDKkK
oo/yp1beOtohDIib68y3Cvuw1mwd76Vxtb8jRf9yhnDRP3gwOSQXjq0EUnctmZQubccrfz2Dighd
AwsOf4CAScvBLynVHYLHayKlwnBqeeDETzD3esxEX5izXJASpbPcKwuBpgsdNwXdd4gXHmeGASWc
/6+edJSUa2pHDcPOd5vDhXrjPFP0kVm1+qHJKoHjLLy55hWOTWcr5kPq3rO+xVnjSWxMPjTN+jId
L5YuY8GgQ5sxtopF+YjvuMqZ3Mrpwjv01k+5+pBx+JmXZwyx3keOlH4njUF52ghwmRD6mz+FW1/Z
v16IMCk1VA87QuPmcPyVEJaljgDc7lwZ0oaq5dTKETS+Q4cxQVuNRtvoS8faDYfSGE2ygn3BloJk
PwAEyPQXygCnNTpCkR0ZZIEJ8yE7Bw8lWq+wesM3VcOhATZUfJQd+LnYnYBlo39pgX97tD/UdMv2
jrTt+BMm6KChe7OD24hWYZmwuTmoPFBf/8RtbFH6awv8pGDViEhtQsqDJDIgYTWkkfpC0fDHM0IN
Y4SuAo8mYVoOhGHTyznB2+5Hey4BgKYPKcZcckpKlmuUz5QucFHyhHcgQRf4Z7TToZy5/O8yXme7
OAoh9yKBugtVoeQailomi4nhDGw74hL5uJteQ32CSdmxukzqTh2nUc9f34a2hmEX3KqlJaUu8xtg
IqoaVLn8kGl/d8+d59JFoJ5yZLmH688futcjredPPkTyWqtDklLEE2bE1mMLg4V1iRXYkbVzHpFH
q/zwoiTUGqTR29Zr4m3ALAxiF4lCUrfOeuRubnNmoglnRidqz/7RHaymuavk1AwWwddg9LGMpAzD
Pm7emaxAMq0Fzrx9U/HdWhjcrtxggHJFjKNfhldC1g3XzozrOa/V/rnh9mVC8eK42RT/uoPpoZxq
fjKOzluW/5YbJdsImWQIJo4ogy31b3AzMU8fVea2W/6MPrCNUvpopHQiCLXtG/yWnZSFo3XtSr7c
v51LA3T368m8ea/Xyn5t0AS8RlV2j4epJOeC3MXs68afNV6BMglZM3WuUsBd9QWzNOvsZaXZRDau
85mIs0c3dwm5v9MY9etTJBqYa16KUwp0znVtH73nrGfVrL5b4H8QwIACz0W8FJYbhDWiK6YlUD5R
+D3qjokeaQqrpsp5w5uXFDRukPjpuqs4qK7fLz0JzY0LpZ1p70nu3f8ZlYPVcXpEDCm4mtd4Dpl0
tAILQwCPJ3iNrD7xqncre88lj0pYkpf+E9+dBpGQ7pRhZDA7vl9g4/xzk2JFmN+vFz4BLFif74im
IeSGNEJiKaXu+CpKj6QD1KaL0aKxEQYdY9yryEC5K/cevOnJxbQJmlt+guHf5MmsIQaoJzhrlnTI
5RFunqYuUw7cWEklcqKEiwDFLlMu80IMm+7GG3qIv5nPR5u3eAKi5FFQZzIkZ/tsnrMwMTDFKWAi
x7c3JEs6/yFsrFg7L00hrX4rk5PheXrQfRJNHyxpHAa1r71JhlXmG8t6Ntqq7wiELTR7/8eCBMvU
L6dHWu7/op5E7Db3hU3hLyGqGleIxr6ZLMD27fyYMKLTAOCdHRlGUeuBpwNDGX8GqPQIm5PELj6e
tWonGxHSmzM8SBe7vmmmDbDUDEdqCdNpx+IM6Jiscm51BqLUmwJLZR96+YtFrpcHMB5qucf4et8G
3i9lvFGeEvQyRPYLxD4Z8jz1KL/MT6xQogZJeimOYe3d0OY1tNHJN1evlRPfG3Q/fUsvJvliEJOI
hSAw8SR1W7BXsGfRwnEapccerRBYOzYOJFQoVlogO/jSG9hcX5//VQ+ytEwBQuYyKvA9ObVh6d9y
+Avix6tMUE9POy1zECEDalcfWZsBVOTZy26zXq4cwyDbxv1R8EGBdRbpjMRMgrwk6/2Wj8S2ZxYk
QvdJWQMOJjHj5evGcAKywNJziAbCcveRSWXQ1RJdkvGWKNMgvmtPmYgKwS05gV8MbI6rXO1EwT+A
gUXuTWlcXav42LPHg+P48mNBbXJ1yge+NpkmTv7qpMmw4h2CNWVSnWzWF/jH8tDFzcb9B43XJilw
zW/ufxcKMt31idyZ8MRy2lP9rXzYopETEn66WQHlnCMm4ulN/zIh+1V9yuubuGxdNr9Ai+qvpzXp
7YBHzLAJnzlK9JysOIaMdknscdLAuEjdzTJISuY8d3uXb1/EXq5+86mk9FbNnZjZ+NbK9IcOMYV5
xdzaDk37CoB+DiTuM/12NXB6CNlmimMYM90XnPO1PPMJVMSoG+MhPCyRKhGSav/G/uR2ikCTNsO0
njOKthw0q0VEkGDRuEvW/oia2Nggpd7gafUtZMMHdse+m28lxISgyyszLLUAM1WGbPT57nkY5b/F
LxLEC7+Ggm5FsWu1KiZVzyKLpPRPZh5QVoHh97NeOAwCDaPKJ6VPaTEtF5ZQV4yLhnuYQkKqyojX
F60RwNuwTXKeBHqns54Hq0Eg1xJyDlp80Cae9rJNelfbcb+dtdksxscB6EmKPNf6ysm90aFWUrzK
FKRDmO7r3Fnw7nzVYduQo7tncVomacEt2Y1Arcu42aTJISGAxNv8wUUmfFIENogNH72dGr+jQIhE
ETmhQ08TtPpnTqJ39yK+ew7riAMaJHS3BHwgO/M3uwvwBDY/I2pFAY+XxI3fwzgNSgA6gX7v7PxB
JJ6XYlaWnxC/o3Qb3Histe469VZ5yv2UzPsoajBArAyBdLLX1md9oPCGtLNAtB2nFNngT+siXpmH
a6dYwfjwXI9j+ffBAlSdWvKIy7rkG9iCVDZJebQszuSYu/wbwYwIMT7UUwly6u+djJMnXWB8e4s1
mjOYLLrxVMH5GQdCg6TgUMwriBwfYYQUTB7EFNkLcp86FSSNE8yV4uQXx2K4+558BJuonqgtYdkp
p7YcS2G99CjhnplMcoeHuVw8f1s8oPeRp3c6vnZGEV77k8cRwDQhYBagtprGQy012b9g6pUUc+Jv
Zx/+G2fVIprQuhrzA8hxOUirmBqD8bTut18XIHErcElYPSe/C8l1DwYKDw/UlJweagoMNK1O8zSi
XRg5p/DIxObfezT3yY2JmeUiS4xBHgBNfj7Ru9eeciJFjdP2ox/JnSBCrJbT3Srypot1X0SmP/28
44Y16EDdsWSxlorX+KyjsZWSiinyMbFwbqDrG0vU/bD4I+89xVJ01i/objC1fz3Xp3Ntn1h4nHW9
BCnBEF+0njGmbqnYvdKzU/qoGLI6iPMkuZpVpIFwQbI6CHAfvnXbd/0vquicDY8cj/or1mRvElcA
PCajs1rx1PiiBMsObj8QY2X8haaueF/Qhx0nirpK/YlReZnhr9Az5xog3fMlst/O0WUpBz1E2g0Q
rJYdvnWQ8LLnIneTn+R7TXcGNJoN/w9b1NBlkxWMdKZAitC2wUzJNzfNIhvlvloFJAHWKu5TmGzG
qIT/3Xa8GdSjMwo2NVJ1cwBYlPrfgvXWRatxIuZglPjwcee7ZDcmK0ivwd+Lp7dPiRQl6b+uXm6v
0hD9aOBi6C0AqbvhgQt6wEWLNf7uUr3Zuf9p6vaz2rAhyrxMSctEBMSyvvcKFkbl/vpxws/55k3k
z8UlAhPpvV5OSUGJx+gZke8VV/0lVXamL6Fga/Rdlnb+pAjkEPjMQk+7KHkG0Yz8GtjnqufoP2uk
NnDXDAl17j2aQoJ2BP5/KS573WKdqlHIw1ON2STzb3TB6/ZsDt/QpDC1VoMj0KL4tnkrINhfTPpz
L9++B76GPxpqfnefWlRsvcI1YRhokGgH/HYn1RQRzEhNdLOExJ/Gw9qqjz2A9n69t3N5ZCF3Xa+m
sEEgbqfQAOwog7Put+ZMOwrLxZeVt+leN3FRyJSEX9aUZ0cBlwlhze2wiYdehNK6dUHTUJCyzLh7
Al+SqtjqxRBq4JZ+hlihJBRdPodKDXQScXoXxb2YnD0VHdz0dg1wgeVqkZOS8AqXnX+PzAH6HF90
iDZp2vx8bUVMp1suX2xuqOxuHEzXusKn3rZzMQGi6B1bRB606JdxxF6L4Th2VN5rl9Z4dpuRbXpx
B6WVR3i310wMwUDVBRKZaeftoukZIgRNLSFT83RuwJiIiSg33jR95dKOr4YvsODWW78D7WAdHqyA
jxHdTjoPmvgdxx86rYyVMj4mdxZsds2HuMhaCQqkIxhx50Sz5BZ7ghcCI3xUnl/6V+SBTlrY7PCx
w1gKQhCf7guBHvnX00sIg7HyD1MAyYaUY977D6hWQtddn+pHArId5+QULmhxWJObwZtC+YwW6lKo
qeL7gHJ+oYjWi2+mqaGqnlLiFTSTUXRjTc6QZ1oBJOTnVq3VSKI+MJNal9xNqDLHl88WpUHmsgH3
FEKkuFmug8qm3fgvK1T12i3wtKmjTs1HkLm4PlZ2R3fQersPe9i80jkTkDRF/wIwEeM6h9WPGl0U
c1j72b4BMYwP8BU5xUM4PEi7vRXMB9F4GkPwrc1slU5rJsed/gB/+nLPnfecXK7gmYSBfZEFmLo2
0lwS6wloV9aPQXT/RMaJ3EHPIA2+Do+d7D7xwTXoHaoVx7OLdaE/yXrggu5ncOAyCVJpqFdDj1bb
ho8hM5Vz/z7uyJgR7SrOVI9lfsjpWOrl8DU2xbaU5aUDb172A6dnT2tICjEpNF8WyhNE0rJQRr1r
Xiz5vPL0sExTQq2tCAU8gbY7McO3do9mf7rYEiLx71K9YhyQGtMcA7mJ5UOFk1VgJZdZxRgoaX1r
+AnQV0Grr+l1iSIuf2Mx8j32lt78eRp7QDngZ83eJiFOofyxvxxjBvEZ8D9aHVvvuGvOfAw0sYJk
GoJ4VJZbh9Yu8VPuE/guPDXt+DDB6jTXEU++02U8r5rAOTQE4Vh/zxZZzr72EJTNkv/dWHJYE8QJ
W+pTGVYqgSWL3E/ADT7AwtMo5Yo032LJZjkqvrPH2sz0yg8rUny7ah3sUwhY5+LbtfOLknnOud0K
xBU69RQthMH26T/Lc2FkaXwYLfJOSMSAL0c5Yby8A7A+emPTm0Nu8e/T2sD21nKqC5X57H4AMJ/t
6Lkten3p2JTDJ3ZFtnDONqkK2ru3B9wkARLC0qgD6x5LoIKy1gdaH+hnm1woUXjbOSAJdGqm9+vt
zw4WzGYLjoIj8Cboj7/dHBx395rV8l7TFVuaDFMXJOghKA3AOtOB9SmIZKYMfdhKqLVIt39Z8gXa
7t8o1yzv2c54xHD683uxT9j1cYLOiZ13v88UoSJBiOYkrqR1QW5Da6b0u1mKCjoOunR4rOTNaH0/
Ddkr5c9Mz/T/oAk2r1qtQ6PobQhPh+k1yImUYgGEBbMvFccZ1YJN20OLkcBqgjRxchsN7XswkA4i
UVIaqjRjDhXXRrT8s/w7tmusDdIabr+RB46tcJ7QDt5ARC4+Zua2BvNmltUw/hxmlHWhHP8DCuC7
YosjuxcweILnCAliJ1G6t9rokx5JOeP9ItDPhFPY1i8KE1AAh9UBTFELISXvbHBOweheo+UgDNTc
nIKQo5rOHVqujVlb+Fo6a4dk0V5Nt8rNfrMUn5hR/Ju+5il1Gz1i0V/cfv4zY1pcTeN+c98ky43e
DvLI5CMHc5ySUfFXgS4cv+OZ7Iqxm/vTMQ7hOid0ybEWgYP2bglIwGzLQZmXgFVM67uarDA/9QnH
0FYbYbyyD+c0arusUKAM0uftzcu1V/W9cxztozhGGFf8R/E1pAbLdmpwLoC4GwZB/h5N4ZiQWRVd
A0MAGb8wtCOu6Cv2I5fX9Y5xMtmA/NTgbBnQSiGXPbGmF/EjGzZtg7CmquQPsNmVHXuLoqzAyzeg
j1V1GkJJvmhu3bm88HB8IxFqXdYKtDdG4snj/4RCBdk6xJSXNfyB9FL8G/4oDM5kqnc/D/s9ZbLh
QLl248wCJEu0ymDa4Xtd5xemThS7LbxJ7jBl14gmC/xZSxLuSnmIcOgEf1yqQGgDNuT6RvM/OktK
aQp0T1bqYNOI40y+DhfN7xTGfjUw+3ScN4MKM9/cD2esouzqHUJDRu6cC0eOhPT3wFjbONnnDERa
M036HAxl9VDLtiHv3nKs/QlNPtzNIXLvxWtgIZI5z6+oNVZsFOmKSCECs7uFyC+cOAu04KFkcmYf
xtrLqdoHwnW2oWydnw6+6uZ4G8iNnvyYqBCOIF4eTY0A89PxSRHaGkK1PpW+iENbNPLRvUec95Wh
CX6neJYRWIjddg19aGkqZ6VMlYemVgPecdZERSqdInsLUzqP883XaIiWlkXsTPldaj6KuaJ7TN1v
kWJx48wuVxGNqCcGzXxRUkarFoLpsWEetaGTXi25hXsVJonH13peujBcCUpubAObRdgzEWYUC5rR
ZDIYCsSWflMnqYzxT2VIS/za0QSGvWwPlm8ezPh4yJNJ1wxNuev9/HizrAz1DX2mpnxuHLW1u+js
8/1XJ30xcUYPgfdaK33jaOjuXyfNMlz3R5mrUVlHtu22/Jk0D7UCObnOxUDVsGVgxCJPyRTN99mo
6HD5hHSYCnkGTpqmGLq2DrCduUYM0ObYPG/buQ5yUAy7JsSjFBOMnE20Bah9CKYN1BhAir3Uav1e
GJS3TxaReuWRSMRRy5csN/P9fqNki5rNP8u/Ww5R1LvzBvtwA9bHxiFm3s5UP0l6hcRat5gV6BGD
K6D0zF2pueKDh8lU9iXd8XWpPAQpAA7QQn6xTWeEuBLr3bJBexm3ybAOGS32id0/BFIgNsIgjg/+
aXUQiyU7z8oa1mNp0aWidwD1jzfNqgsVJsurFWZrgsweFiYQL/zKN1mgqKCsAVTyw3iXC8d8GLEg
aAi+RxkJLUZI1z/Lg3+JMsUB5yoqEROwWEdKfXB11afhwiRo5x4rUae0Uns+I66yQOe/p2dL7Hxm
hbfkpALQMaDqYGDMTW4HOY3SzUAnCEvisqHao0o/NtPSRICVMffHG8I2OdHYalyKP6iFCiIXrhYk
e0xyIOVnQbvvztav+qQ/m6GQuQYwinp9BeoYTgzBB9zX20D3vnWdWHr6NS5L4MM10PHAkM6FQNc+
b4hOsCPEGg893o/kdPmLdCkNYrpLmufVZyhMXUjf4Orhn2pt4aiyYzl3hPrMrpsXv9aFjb4MY6V8
sxdUen6QMupUHbbjbYxTeBzRsPN0rDTi1Iy3+BSTr3PEgs+PnOTkCGfwpG/hyLXOxdmYippAavD8
YXZBZ0wGetRDJjZuV1ZDBorFKgZisqxBUdMk1uKuzuoaE4NR5rMLxIPm16zgU7aIPnyyj9qweUtg
PG5rhz1IOvtvzO5jPeniUjKDkWc+H4shO1xYsgH7naBLjgZ3Kopt03LBGdro0EZdVuWF3DdU40b8
Zq/OLP3DFk1HfAFB48Gg7hXXabxLgm7VPKihML4SMeJOtDjS0lmm54X6h5sWIa2EM2TAtlk4VcYB
ksh/88mTNIaHIomJlV7rqmNznh0kgtEEapLOY+1NViUbF4tC7ZUjNx1lZqirKYv5WWfe/G0tYx/v
+50WP/YxM9ykwvOluFXLUa+ZNt93tdPXFvA26Zx3LB7In9XOPHbwfd8rKXjzUjEIPoOwm+/P/Yem
imic0HoiU1+HkyGO31iVHHq+A4beDhS24yndewRvMiENoTjiUIEezU2tydA8zKFCSfpBma3jLBIw
sdggCj+vNKWOWtLb3HBd7ghSABRcsfWA4PGEXB0gvB4fzMjgHv6Sg6i2pYIwwDqnsDvLntaXAFAo
LFOdxR9GOMgcvt6Lbtmn6e7MyOA8QvIsO77AiD7Wgi4Iv+jqvWZp9tYUqOkts0jSb2Dy8jFTCdDr
Yzbf/JYcm8Or/bML8jSLF3hM1s0yfvQ1c4t9d7d0JyL6zhUYqTf0OlOlajMjB8ihm8xvKjEtkt/V
oCaYK/bfbv1KUqEcxHIYYZ+Ly88wKLdkqAI9PfgSZWY8oCYZB1swFCTPkpo9ubqdrVUoqf6ft/GQ
XmFgS8O58WwBMyM0dMKg9LMBUf0+WevLTzXpt4kQ/pvb8g/01PfjxjfB8etBwBIju1n3TRKsB6NL
VGcs4maVArYctifk5NinrMPo/5D97Qkh6AON7+ZEiuG07VBcHU3OrdO1ZVt9JDZp89/msbqSjkIO
wOYTIjWJeZcrYdnIklgac7luLAjDg4jv2g6Q7IRYI/aoGmiDtDV7oR5ASMU5O5ZLSrhBSi1ZrYjG
WwlC6+OSjN44Xo4ubBRMnwAQngQLFoRgng0PrfgESqL+uIjMmqIZ/xjNTRFOaa5hBrj1kGo6PSOP
UJ1PJppX8N5JXyPf3NoOvm22AgF9+9odkdevGY80S3oyDj9WjaQrngsbCB62uaSOVi/lIGc84ib6
LaFezOD5hqkZTqhCKlxW464TG5kOBcJ3SPZ/W5jy+tkcCM1R3O0DfPYrqkbgbl0DgF86aJo1Jk7F
98Wn63wgdwWKuCR3dthbmneIWTRbNTvMjg+WnIPW35zr5GbdNCBItTtVhcW87StAraJ17kwK6w8C
6QBMEItf14otYasgsbmutEmjzwfqWCWpZS5bnlo8pGUTi02P+h3I6dHv9yjc4DVs+pH6HO4MVmjc
JeJVWUop/akulnJuzWu8zXdzZ5MGjIdavG321KlD9KbT2/kRYTUAsoRuaD8qj0zlIXx29pW55NZz
Nnrsiw18f5+FyTxiZs7dEZOPO62512VSa63f6NlwwPY4d68b6ERf6etFspLX8nx4SB49lj9Zg3Vo
FABuxRLnm6hU7YNc7yI6ZSExpA4A6W2o0jVB8DJ0icOUv6luGY8m0vXk+B/UvAODrtRPzjFfV44J
lESoupbL4yH5CIqZIwyqgPQN+wSWvIH0uLeZanBdSltFH+v5/Af85ZdPevDEKnzeRozfC19uxKha
5RPZJYLk33eIHyjSnO+CxmK/heDrEZfYmsva6AiR5XK/nMbU9Hizz8G3FmK4xx7o3riFwtXjFu3M
rnA2xKEAOjijj2kVXK6XDWkr3bLIe0B5VOnfc1d/PAWK3GseYXRt0Wen/amyQzudHFIzJIioFgPG
fgDmY+FQac3tSn4z0o3+8+Gs86HpsDLnpuCQeN3nAKUOPBTpHJCDtDbmlpW2VE1Zn2ideMnshnRC
OSKIrP3NCoZWfDgO99u0fx20IkGd9liP8lJW6QlP5KBaFlNwr2ufsSLzHtpdoLjddeXFZ0bcRXFk
Hk5ksswDCq4H8IFYog1MCb+W6I4LjRv0F2aPLLsrtjgxf1oCMo+pY9Eaq2u7b6UWrBdDfcShyjl5
eGhDah8AOg4PsVUQtwcWCYP0LJvUj75vsZXKXoPjGrgpkBACqc5PB2roNaG1Bw1vtoRXRYLAE9Lr
Givwd/8WQIkywTLIjziYySvYazD7RPuH184XWavrFvC8h8Ub83VRst3+tQy2ZWHW/kQz6FjcBQow
Z5U1uEqpFUkvXXp8Xg6xIhuIysxBlyvEEEA37o222bktUDdZR5cNM6NaqDKcZ861vjKrjupqaYNl
0tc2oo9QIwPKDgAW85zTrsgJSRjEBC6nTpF2k/il6S3uCfKbW9sUUdTZZZ4UfHdUxQ6c/tIr8yJF
3TQZbWIGuHLg9fz7sGupaNktO6WDRM8vd4uLXRuvpxx89M9qg6w37GhcCsa4bsZtC8ZpwbdFvvox
itnYPlnnl7jD1g3TNXiJABSR5KT7fSOrnB7hrG1dFL8S1WhkZb2XcalcJITvDqLcFeeoSV9eCQoK
x9Yxg9jIh0dE9tXVkYikEVYvcz4XJ4iXCVtX22vUXcAoy10EJWFLYwPyijRYLo6BjCg0M9iVYYc0
hCf/XTMo2kFrsGFFDu7xETGErd7dKW/hGxKYxMZbZ6e5er90MSOs+OazIDy5W/F9BSRaXcrBQ+zu
XOjAoRv3aKAD2Kr4zSTecg+9T9nZfm5uidun7xR3NtFDC8Ix87KgfvBjTXv+tGRltLG/JllDgJsV
oW/j3+41B79IoQ8/RkRMT8y/7Lea/Ibq4lShlKixQfD2FA4DyKoFZ8EwkCFv5WOE0GGHPrcs2C3+
19NWtXymBwGUAtHP01WOih1+VF1uPL8I+5HDiAeboNlZFtxPzjfScQ/z6eA6uoKDFa26u4l52VFT
7+yOeM4gBd7DevNEL8fzMY5gzMQscoK809ZyvExt/rxdf9qx2xmvBSwlAqRP+ObFQAsGQe2yfpL9
nFkr5/fs6pfphimwdtw8N4sqdCUbrChCZp4RRmU77ZEvryJctEZQzcx5dyk+1pCaWY/S6W8nNdGp
1w+I/v+Nah6prgpKZ2cfnE/pmDk1Bc6+dPxl/fRM8abvK7a4NCa/iYmx0JhS01gxPFWcjGzenCMJ
0pjqDYuyvL2WO40oviUP5QJ0TNfYlgTUguo1wDPsS0Eg+m99epZxfw5ykorvRbCU9qqCZSGsDNVQ
lhpe5WpIE4nxs50sWrMPH/4fBzcEWBxg2Y7m4fnMu9zf4FQcpBghjGjej/CKvT9UpxIZVFnsVdQh
1ZHkdhY3tI0REHUmzzbuXYvZZR0oGKFChZ+KGiG53KP+sSLdci2bLRcTsutOgQ7ml1v2hRUwTI+9
aWol4mxMRzxQWGdKyBARJmqgIA1q5qVsiXRqn8g+1a9kWe7L07P1G1AAKOPjMQco7Iz+iy/JXVjg
cUPue4T9Lay97EMm8t7+T530iM8bMzbOqmXHHyKff/NGoBAHdt3S93nzF8jJfdLe9exJTnRsuEn6
ysDCNqBsn4FHNw6PPPwHKXGVrktO1buIMRhdjn4ZKRu00RlpnlNXcB2upezA/bpDyxJlq7H5UpGa
aaT78aa7Bjawq1bhis9dqU4qBr+gbbK7v+bU97kJBbzYz2Au3qYoTlx+E9nAzsPM+oka1sOKuYeZ
oyk8VSxhbzGOk74og2sGp8GLlDMiaufHIn+cBuuupH+ltI0xvPvAlNeiXavXU+rcG4IVI0JOOPg3
8JXnaydauES8kbl859v1XTT/NcLPxhakPY4x9h/0Pwj8sjB7T5Fgswj+sVwWVNtqE1KVTJ6EVWZW
ZEQx7jqpriEkLY7Elk8/TaEcLWV648TxwMu+1RTzciU9WQIVKl3RFCTxeYeiroLwz8W6vMgzahXX
Qg5y10bcNnEmHvavpQzUm3o+2Beza6hzFn6wFg50iFo62my0ZmlPKbxQwS+qrJnfXrG2k89nB+qn
jXIXnF3Cc6lPrB5CACi9KuhmmlQwM+azhtbBSVUGzAOBOVkq21p27wKbCNyc/OoBjn248VTEBQbI
kFS4vijZZsCUGgp5UAUA8Xa4Q3ZdKZnAbLM//fG+VGCB/z57eCZAE24eOvPciyHFArbXGvIkCRQs
b3fUHhOUlfaFZlAh61Y0Stxw+ftZDTJQpTEi4NTSFeLoGLUk6eK1ABwl8vXdWsFwdlHx2S4m9KNR
+tW3K0qDyW6VSNFe2FYPgPo2l5dc1peMzwb/KqX71usO/Y97fX2H1dG907dGFKpdTlL95rC9KXBm
swcxSJTqG1u/joyMoLlo6qmQxf1GJC0VP7IYPGCJxwzIXMoQJ3nudtxw3Ji2q3FRdzkIb2dwKWWK
oPxweJZV0eqkXG1X3iJN/yEhfGN/ptcwV+N8bRD3n011omgK+EifDkndN1sg8neY025EOMKPuUWK
AAVofyrjRw/0Bxk0zAHX1bT704SCRTol/Dey9pLXLxLw3AvXH+eI6T7w558eMkgPNxZfudUt+nlL
IiuRJwtRHivqnVWIpqAy0tR1ZUIkRuqSRiJrMTowgb9H/hVPuiFCYTOM+gkInG3OEF0IC4YW9aCB
RmY1XRX5efwzbZxnXLk2Kws+klRYSP7+erDYS9qOIleL8AsuacvIlfNmTxxRdUs7mDiz8FGYYb0i
sssr3E2+8hmZBqG6PJ2/GgJ+NB7XS88Ix0i93dkxyZXPk5vmetpXrj9krTICCw+hZfxiN5DKBaAt
uv+nfEbhPPbM6BrDUWZDHO0I5trZ93lGdV8VRMJJEEqzJJjzLlmBrqpdRp7jyzhcbToWB9gIgJpe
bMhjs0JLJVBgykGoLT510ZXQ9QFfV5aEm+ysTHYp5ouZHbuCDpyLKrhYaIWNN9Y/NW51y/Krq2zq
gpUbxRtkvk43nQn3LpvAsDdf+Sni6A+OYMIoCnOxAe8X50CcwJ1hcfI8Hgl0EJu14ffi4irqO9JT
9Yg70Ejnm6Cq2qhe2vTG1DioSVOGHUKvoHY3+xulw7OI3soDTQsFmog5vQLcAsIGaXDTqoREi+s2
A0jxMN1G31vFOSmlQqGiU1tKr53MeFvR6gcd8Fu3yD22LahRBsisxPLDAqGttYlOc7se9RLY943r
MWCw/k13KzgRPZKMuShvRYMiMEi//3KOkOZVXSUX6lCISA4mrmzELumXgTZwYk13M0WMOVFt+b2P
CpOPwMLPd+NDPIQ/TaCqBp42YrIkhNgRIumTAwAjAunKUEAn41CqZtRv4GQoZYwLv6gTN7fTfNeA
6VjorihRonIDfnsCEix8TwOEMDjCh3O5MJ6mmyvW1pkVpgA9RPi+rIvwIIlivGle6xN1zgDg4gPk
sbb0y5AHW0W3R0xhIT7zQv04UzwlRHO8uvLCypIGlfZ6qMjtr8HssBTAFZdg4uRcZVtUTY5Rpats
kFFfnrQ+Yr0XXwFIa57ybBKrR2UE1B2LsKjyZKoek6l7rMOTxQb8ZgLB/3ZSz5ptKw40RkZAl6EE
lOBfwG9Gti4OE/xR/m4cSwd0Tchj5JAcfMKBhfoi5r9Pdnr3xb5xqPJVE3/aGeSHZ0HvOIrHvkUj
Aui1xJka9Sj2JwXIo32V5aExK4ym2fNf44jfjQbbm2YB+DepjDLWWW0IExQutxATHk9mFCWVD4X8
dV2uCthMQBwuleRtJibeRmdFrZ9Wvvz3sJD0P9AM8ZuNwJtC/F1owqJuDX3eO9vd+OKKQFPMXOql
k66JIL94jYRf/mCcE2NIO+i+X7eyVvDRofcDSJwDUjBfMh2RcvjTgAaG+P6PHLW1JRvIwMnxT071
uHPifD+2+K7u1VoOwSpVAiFowuoye8DLjnfka88knkQlbp/7AKPXX8DlgQv3XW+Y4SjiUDBOSPMq
RVObJuvRjXrusjzUhicFVO+9fbjHsFJxEvuI+bDwyDfqLjf0N5r5JqQOGBTS+3D8xO1gtlAh0AYo
dTVWOImJ/bmUYzDqGdOXtmc8+j1W4vmcoENAtMKmXbaV4FKXGC+WZIlI/cU59d3IMsDMYSsl79df
NPqRoHTExVpC2KVxLeOOtRXgXFAiYjuC4j4zI4iQkDT9lW+3KbV6F/fZ9wvgB2QLF3RN+GZliqMk
yGmnt6WzRNxi0RYnneuolNs9lp8E0Ui7vk7Q8SJbOQBA3MDeqYjWnkcyClM/4mZ09Kq0i0V4SxVe
uaRwE586p9T7CwhvuefBmBIE27eLA1TdFJO+323QSY3lYC/2gV2j3GePAoHIG3eKV5aeBCYnNC8/
7oJ8vlpQHTc50QwhpVO6XW2rHhNFvXDRQ0GeNcFaqgp9r4gRwFGajwbXX71rTJtGCR1HfbdX3vi2
B+bKChsx4H5O7LMkqXUgs4tXjkzC7ZZIky+uZjdKQmQyyyKtAyRPdcRxuxJZ2kZimLfNHaN04fa0
E8X8H4RA/tj4l/kTG6TC/UAhgSeSyl/p1sPotGCMgFCME5pNj0aPsNGqpixrW9Pyq9oZR63lhbUZ
QQq6tgKrjvULj47dTRQhLHGimvrMIYY1Kh3MGsUmcpr8Ll/1tnTDdAH9WFyFpKBoKDWPOryhqlKa
5k2bK5St5JqAO6w6N39naihjvdg+onob6XS0PcGD3Oj35NdmZwJ8GbL/eFfuo91ukKKDRwrbczlq
4VjVgbXPiPm4Om3dOeAg4yJznylivhjaVRuFbKi+uUj7Q1HWoQYGK/isE6lLNv8ANFE8xugWJSBw
NcJRI9a9xWOu/dYXyKIr5NaLI7woEuYb+UJ6XSMYv4RKnKomQ/IrEDGLkefa5hfSE50PyESfLRRO
AknApPI98EF7aFZIA3qjWmowLpI5LPOgvZhSSWig8KToZ5yw2ho6cLK/zU/vitwOoVOq2ferG5SO
w8tCoYcElUoyIl74/Lv7Pc6FcYO4rbXUAbKwZnD1524pGjgfn1G9UgVWFmlw9hLDB57mBdVcHeTU
9OqByCBIL1j1KJgP3vE7OGvgdBrLUMDSyMHxeYiHwcHErIu4XRENSTSYVnWywdVJxt9ULw3GPp9L
pvFpBXmofQVzEQCUEYYh9bwL+X3SlLcLlKSVN/CsIOLNi0stV5u6nANUfvITWkU5JyXS7NU6y/6q
skiHJP0uT5yEv5xdk3PyOEyYNkDaBaqPfK8ygc5Z9LtDhht9NdwTZy2cfaI8VVQj95vSGkBjprzN
2Wz8mIfutZ85U83XU10QE0va2PGhPA0A031JbpP3f7ucQqa6lUnb4RnO35zV18JYGKzprdRzCXsI
MOuCxOnBQo6BiDU5jqMMjtpiRxYG2a6nyU/6LzSycPGfe5zmmM43TSQwrjf7oeoyipEmyyoC6n7R
rDODrB4H4AL5Teo5UtbIwlDPtHGQMiT2KLTTzrPRnP8JWqFvKmi0yfQrKLW34HtP9YYO4eO/ktaP
k29XX8RmA9hxt9AF/NZVAfzILd4HwijBiS8iohHFiUTtKX1lYnOIQ089CQK3gCQD08VscS2RT6nv
qilKjgUTYmfI3ViLs4W8H47grMMezP6PwqRtp6PfHPVOC8fxhjrn0QM+7HDi4Dtt03AhMM+qhZ29
Jp7/1mB2SOZXjznXE3cDszolx/tlTCJLQyFyPS7refnG98L3b21UIXVxJV31hHyHv7hYhA6DwJdR
N0LImlu5rF8/1xkL8c9t2clXbgNOfRWnEgESaGy4v8QaAvIQx1n7158JsiCD7wLeEfY8eSBGhAPi
N/Owm3P231n4U9lMisBlaMwy4Vz0Q+606tkQJnrcHErK8a1sXcBuxJcqpIm0Z+7SpCtBUPfQ10LU
e1xeahx9OwucgGwZ9mYl4nVTNperhU4v0Qt6rmLmeaLdtrKaCeqcy+geUTamIAQaA5ex6yza10wI
1lIbuQ3JfDi2CZJmp1JIAyN6a8pOoc5SkiF+de6XXUtxVB9kp5pQjuZ8CjqOVeIMxl/bT7n5AJgX
h0BE9AAOQcz6NvLPkaQ0EI5CHtRnWhpzGggxYE7rSWgIkSBCW2uamB7riF8tC0oLLxuqnAyssEu8
eo8fW2v5hISfovqjuFPiwpzTB+1+eom4uveTJBzmWEHn1PC3m1YqQXiwybkqpYgkF94awKk6nGVB
tqpWEQojpyon5np62JLx58v6S2zOXjFB0v7eLEPey8+P+CWyZjb2tBu1UXIjh7iGQKTwJoGktFOO
RrYbc75TC70NK4N/emEC3C/MgYxoIaQ6CxesczKmlVZfFvo0xZ53aS6fRDDeg0v2vNwojv22/J4O
1O4mz9xcfmyVpnJdqCfcEdz8BIReml3hIV/MSS6t2yzBHPnkzZ9cvN7xmgRpWyBg0K2FHTiItOYx
zEJlYURR/A+ETh4/5azWVOjrl5TUaFGOn40iGSr78/bbXWhyFLUzPlBeQ8nSpb0OuYudccnCgZth
srNClVjV8NS8fm2chKRsViMX0ZfeM+9Z2W66MzZJR1IX5t2CAMopPm4cN/P5mbTmAuwK4CxK8k1R
+5hqKrlVkRmrVHWhuS8hzy4f+fOi46QJnVg3I/CTsS9lgQvaY7Z6VTdDA9lzVoMX6K7Y9oZv18aQ
tne8hIHbVdCp4MpcYbrBUk03tUezEwI5P3bcI0EjbnydEdC9K49aYGQW/ZEM0cO+mLHUr669CJ/G
n4VSZxak4RFoCy1qsW7L9BAfOLZ3gsLG7svkViRqGrlyCv6EndjdbLu+ifpVkDuvd7Eyvjs5g1vz
DriBJU51UEyoHgiXFRlLu9KodvHJNiiRYozqqL+qhbaHzw2Py3dD7Reqsh3jlQBlffUXqzcM88vH
c7kPHeUJ+wncHifkxsQuQTVDXTnq2QcvoihR4Mwx/jgRTwosO+ZrTXD6qNc2gzKI7Ha66GQjVrZQ
nDS2I13NARD8shFklfYfckGUrY0QiZMQRX56l16CO4Wq14N6r/RTvBxsgnIAzfpbRapbV6kZfzXY
bn2V8cshio1PDQeXd24q6xw9Cfe3oYWr3c3WZliExAzwnn1fbVdt1RSuISFfyQZwVbrKAZnynu7O
aCBeFUpm3hdPCJ+sWRQNsJwEL1kWePWG9ZUUEJmxr1w7XDTWsL0Eat6zR9aexl3JjwsEfuEmjK3B
i0+MUZJEdF9VI5/DC0+YCUcFXzMzzXF+6JzH89SUYhchL/BS8hFPDAtg+qXpPal9geKTiN11x9fg
JbK6dZzRXc1FXcYzLtHflynZPXx1nbnVvA4BQrveg36ehP/8M9mTOxhPbh+B/ISGDwlE/+kCV4i3
hqgeibmubyO4iv0z9tLkVfPexzMA4NL15QQBWlJH50Q3gV/+a/j8WH1LPY+ESCn9di3ir3qWKbGj
L4tiIudWgUkekHUBnPnt6Z8Zrzt2W2FO/Y69oQdIqCTg500yTaSEN5cbYA25GQr8oVGAJZuzNJm6
dlAkYyCYqRFsXMYkYry3d+HujmLUZkBE+LJjaGDfE/9GYyHunN2BXKn9fJhAuL+dXFdnJ0zmXheL
eu6YtQZ1soM+WDLtcpTt4osun2HEo3sgEsX+IrstD9+TDSGLk0yJcldWPadX0bLE1TrS4J89UsOS
+EmLd5VRqFM9QWgyCsN0vXQW80guYIcDTjOHM2H9x4j3p3+NBC2fOyjZK0mtArg8XnP4gZVeh1Jp
ewUta28kQFx2RY3Tj8aqLiiQbCOiz9SV+TrxaYaN3/xFKwwyulyY5hTgS6+HExcYq8fOkMK3te9D
3r8tFWhRlPd/RiRbKfe0D1ldZgBqNhQ69NUR0EmH2u9HRk0npwr+bTYs23N5C885+1TAxpuqr/F8
kQwqX2qSl7xDoYijyxWq5RqVTRmzqiTBez1d/W3aYrbevoOchITeIxpNtdNpfcoDTUiIGkr7J/+j
RixKzKDYaU01JBT/6BX6KVOpxWZjdOemNSnF2ULjPM5IpEO081dd+ACmvwbX5/6QrZi33H8tE+11
j4oVRPtIkkB4e2cFZVl6oAo8IsT/cWJE3YHH/9XWjPVLnpPF+ImEnziLdWR7/F6uTCbktkaZEAmV
UdopdVA+9KwFnCrLNkXerAHamrqj0ouvprsBx0YhMDI1Tu/Z/FMXdq+kLHw1R44ZuV0yPRyIedOg
D99oSgJ1g5Xrkpb5LfDCdnTXcDAQ9pCL1Qh+rF6v1cnaCOOkEgCnBlu6OmfA0z9U/6Pba2nsro92
GJwey4XyqnauTGKYnE/GnSbVEdXRR701/YVFswSF1wiW4oaGRbu4FH1KLCTGlK5oSXMK1e7fTc7s
vwSJ1RV5HngtUAiPaZpFSnyeNsON1+gT+Rxw8hy0jPNmgJIu4rvx/vE8nZ5WTeA7QwxF1O5Xaw93
aK/TtRvpS7J5gdD3HPIBxaiZNXCXdfWd/8+Nypzu88HZCbdDf2bxYZu/6x4JiLJCqwv+mmb8fcBW
8tZl38WNCmeOuYTmU0IPo3nY1Y01aJsjOE7RzcKE6MVwUtQWz/afJFTAFR7Hr6s/wE3BhHeNTlDg
f/YV6sy/EK3BV2EuRF4o39VM574G1MacBX/WxrarhX5iqcLdcjx2ykkC+E9lukuIbiPsS699R3Gw
JuDPNTdPBV63r3H5tBN7hSdXsW54g8vCUKkdMv36BPfC7TerbU9KzKu5O2nzby3A5Pqc9nrdIKws
8TuPqkyhibzcKF3NxDYojfLeB3KVuwCp7De8QZzUvcIoGDoeZXoSvDECb4LGQCCtdHlXYVjhDSRA
JEcphUiD5w0BZ/lPVRZxP+vRMtkZdsFX4hi+jlmlDfcY1eYM8B37WCmjfdSjdGAJPm3FimuTzGcm
rwe2M6KUPv2AMXNXFfskeu0nkIaHnpo4g0+YCaqyp9XXrPBOVF9ZCsXXJp1pNbSmPgdilgT4hMSy
Un9dSqFAj/rgrctKVZSHqGgXV4Wl9TONCFF+jAuNgn7GYDKl0kN7x8pPz35ugH5OrdZfhwBd5zTw
T2+wAQ8VAU3P7kRD2LTRslBG4G544HNRAT13mYv2LC4aKsjHKku71fBK81KAq7CpmZ9JBb9n1HIb
mfYju1FnVOE1i0xG+2SAQeGs27HOnKBHO7HL7kmN2xZr9iHSICcS9UMXmRUm08bG3AEgR8q3oE4G
EJIbYLxNHbO4ra91B2dk2RhXeLOgaYd8lG8k6LRuvfqNhHXgjFw9uQmDniLizKf6i3WPkhcJh155
2Q3Mqk8Yg+VofE9/a59yadtntw+e5GEG3exrBZgdXe/YIFQD1hYEOuRAwstuU8mfL8frO2uHL06r
+a6X7yL+Q48U9JCQM6Fo5kTk+/IMV+c2AAE0CzuWSOom5KIzCuAntt5TapIPzfjMUqVm6TnOaNiw
M2PhPk+4C8ghcNH6wae1y8ajUDBKs5LlvYHopHT4kklu7S593Nvl6pow7Z/sXL9s9a5awC3+mhih
Vj/ztBLJV+4op9vkQArkezDqLAV2vZ64pgLNRBKyA6TZ30loGDoO27tZ0fAsLYvS/XsqZYjw7EBV
5kS8d40IoASPm9jzxUQ/EfKjkAfxpUnmxV1Kdhqm15xyuOYEiXo02Gj/+QvWZrPwHP5rbd9n3SW9
nCjkZP5JDKuUwnHbn837jUlA5NtBmXxBFbx2zKRz1yA+X46rz3IU5NZ/Ohs+rWBsvTREfwKAbtRM
gR/DMig2ufRSjg+m+MRQIGJ7ulCMToWc50Pko+V1aUos++hoJ6V6Tue5Wrq5Ua9g7E4FGd+/wZyj
B+fG9EkDrpw/unaflwzX0dBe8banV9iSZFDBXrtygvNNK7jx1wUKNFv9DlKhCSKccOLfdZif6Krf
sg0EBgoXY8QgU5VkBVXWZZgBOarb+DLQ1O0AWvcaMO7Y4bxFetNWyHDKcw4cry4aY/98wXELtky8
Wea299Rml0gHutQ2sSG5zpS/qk7LzoQbMRTknENb8pXX1TeDi5Dwp+bdIa2zC2xVr7ocHzuZ0o65
2OrxNPZn/9H0BldvFXm1Xoo+xH4/5rWZgU9q+uQJ/YNJIQ2fZsStq+8G7e2TpKekRk9dfpMbQ17l
ncYlh6t78znJe8F8Ce4PRgDGwpzId0HT7muLJTiAQuuV8gowWEoCdDy3WVnKphvwNZnz0i+Xjsh1
74Fv32XP+/8t4kzjURoqfwvkZwLBepFbRbuTKMK9MMMpmXp+x+dinj1JQALt9bDIsVidXJ30K282
/AFr2y6m09rtQNSGLeS6jETktza8KANs4EO0+nGbXTfzKA3ynHyVMbLodd1E/ZaGibTrQgUM7hGs
4a0suRSVl3eMMIL6PiIpF+LWGEb8GmDgkliY11M2xVpeJY4cnj8PxnF1m4dz4xo+0oEba0TJVRbP
zpYHWFyI8UQ2pQfGg6R1hnhUazv0GGApslFCGbTfZMBaFWBdJTKnZO1O1Qyh3K0v5rdSkjYTYqsf
+i0caLo0MWS3alS4cLrLtd1RIoSXsFdbo4vEgmsTqaBJMO/OX/TnJdn+/ABxrJXJp5SyZpLI4AaI
0QzUIhI02HZYx3CECpk9Xw5OHAjmXp5KWmTaksLurrMdzRTNF8K/l45JvuOmWQKpwv5M9jrylmGu
EGQdoGABlb5gjV8B1tVM/QqZ1Axbl4k9yJ2xbb0cfhwXQQXnMspc3E0FczaPMCFigktWFBFmt2J/
sLntIaYbUFdaqZVPndyBv8VA5XAvZpV8x4bxsz2CIfmwUxObtsWsvOnq98Dfn4Z4A/Zrl02LBl/G
iRkGAfaA2BUwqWrAaCpRzByNQ1y+Iwyg4AuQY4sUDww2uR5HWBMAk761vae3BcesFd6POxW07iXJ
Qr/SwmR1EZ6ovL5L18Xh/ii/kgOuPMwB7e9TEWl80cRlF2D6OEF3FAz/U+x2TW07pixMb36bAjKR
WZPB1z3kVh/kFbJK3C6QdZcoFkPbpZ56kwIgkGQmwsnokKCQ5iFFcdbHvPQtpJDm+tGSmrCAwwob
vfbFIKRXHlKe7ls13lQEZH47RUq2RhqKM83sc8GYgvzv2nQXhl9saXHJbAD7mEu/XdsMV/RijOuk
+yR4cUfbhJiRaJU7CcgEhXwxb+nWpyomqGPYTZTZBYcwc7NbQx/jg+clhT5voBzmH1maN+P2+1j8
EkVs7EG9Ee2tTrk42m1ZujrbjHlNpk39f7PDm9GOb4Ar8Sc9d1r/fDBS8f5lg3DLRl+t+r5c12Q/
AhJeu/Ih/HH2n8r5YmY0hlyni062PGMK8EoQXGyymHMXgvYHq7QS31RLnJ/5LGR08mFwUIUP+pux
u095UVoIsvYJMHurpMm5tOSE6F1zewUnMPwb4yBCzgorKi5l4hrWcwzV2sVCUqUPgBHSILhaJ9gq
uHa9oD1wJsP+eKTNDRKADcC1OhSLz6UQfwtP/ODNaWNWFI+g3SApUtJLRb/BkfM0G5w7AMTHJeJC
rHowp0BcqoiXbmL7tLEXJ3uZAtAjo9pB6fblvInVhPnE5EQfSsYdkTsxoj9GOd1IFgDc++J1KVEs
JUx0k3NQv3z5uCCm9vRdkB28B0HTbsKBSGFZNnKfO3JGHMfeV7NB7qXvEc53C/ChmKd1psFvqSxF
QP9wBtGeJFyz2NuCTFZIbHK3W8kuSpx2m08ujaDfZVaj6VF5HU5xClh4sOygi08bgdCKrxhPs548
3ezlt99PCH57EUGBZ2H4l/xDrtiGpOmDlPQGEEz85XqWEhjkkmrVg4YPo0o/YSg8ohZhcNV8hxNu
7IIBmBDKYjnXTxggWpGP5mCpx7IBt2LFvr2LjX6jw9Why7W6X2QNMJddZ0h6p6G4fxwB/o215F9H
UYnreCZ5ZSL/lqVM7MEsKh+i+7IEKvPczB014yoGMeTIHV4yz9PzjeOGwnuzwcfLE0c1sloyiBcM
mXkPrE81mOpZv5YCeSwtUltBnltoFm1aAa7dy5ldOsGCFX6mE1/g8PBZrfS1fesmjvQ6VDusFeFa
/M/PvKuSn/7uYGNQZE2UOV7WIvlU0ug1C99GHxqJWlS5jJxnBH3lt+Ue7IXVJK64344s9Adl1rlW
rPdqhFBAUgrr0LfqqUxPITVz30r9CoEe/VlHseuJwNgx8zz9bMprh2DDjxeKKdeyxZrt8D27lJnZ
qEsL1WAJjlPzQdroQkhE+aRCxkZ2Xj5uvlNzuUnDmjECFXVX5JISLlnACxAj4iMVNv+dOTUG4RWg
wOU7aHNViHrJl/259/8K+sMfUswuJ+vmZeAnBpM1kdBbf+PymbGKNFZ/B8fDmX7lremFH+vTriIC
UFW0Wjsl7xo5Ck4xVdulytBN305wTzK4Cpbi8859cozVxMTln0Zqa7OErmW5ov9+pY2MYF9lKpJx
H+53Io6QZVG7TdktnnkGzl7SxBem325yl/g3p4TFcU6hzUe9C9sH5XGMDBFV5XmFuBs7XiqDOVS9
9D9M6KO5gSryLT37v/N+usqTOS4c9rEi/MsUSfXkCTQ5vm7f76l5ea8FFaCfaFiAHemGv+CZgRVA
FRLRH0UYeFgB79215gn/i/Xn6nJ4Fa5bGJvvcc9D08YdCkU0WOpU/SNp/FPiTHI31gcxJ7x3/+xL
s4cIIcg2BMTxw+4Bu2Gul0N59OHDfrwLmRk+9Ig9BFw1npzmi9T+EalWvSyS2+iywuA4JSotZBL8
gqVpwfCFzWiEBwtLUDTZ7Kw0MS2h7pT6VJk+wP0grSWJTrzDcLk4xdizZx8zab73LlHNDtnAqwXh
LmFQVFibXbI+rDJ8/ABlENyJmoHN3uPvbAen8dS/ToU8enMDdiyOAfx/f7CB766sJdb5jbS0DR4t
FXg6IbnX5m17Welpm0JM6T7ibDEe+nG1sugUbJsC0MzcNEJB6hlcbuBxRDWMM711fynQIixRsjLK
vpPeOjjIV3z5s41dD3tACeE/KJ1nnMD8x/o2lBGwtctMayasVdxpRkDw440J7OaWilmxlboPxPj0
Rvor+kc41ksZjwtWiYkI40ZKyVnObRLB42a19UPsT5R0Vxs3PeImvi8ipCscngjWGr4CQqgkSYMA
hx2R9VwQP2E2+WcaH3QojlSXUCS7yR43g86QLYp090pgd+mRI5lIIYTxlbgVVgN07tdh4sA+fqjA
NWe1btwsuUF4dC/j+YuC7vYNjMWnP4Sv47tgzA/7FYRjtrm6qKMBSab4TKNpo9H4+OuYUpmBsEJJ
UfCKLfANzbQ9cvwEnJ35wuRh2LF/dYs1Jf+D5kC2ftp8rF+Vzmqwio3OG8klXLzHN/EicOLAnE0h
xwqVStY1MIfnTTrnE2TbaFbw2inK+MPcLjlmj0ocQLY4QorufWEFEeHILRuptzp+YMkYEfDnlzMA
5DeFk4TppGjKINm+t7mVgYvG47Cb12/F3qhXMu6d3udGuD7+XaXrs618ZCdpiAhqQ2mX0Y5uoM9D
f2Bu1GJxVTXDpYxDuPWpjLXGsfDB1CTHSSikbBUpdFcgf8A3LrrM7Uv0r9cP8+x9hqrmJUmagNbT
/LQX8tHFMXhKr6blxtkNoTA5Fd9B89e+JgrNuwtNpE+KIr9u+p4QhhdJekEfDWs+ZG6nZuORT2Ds
kTx4TPHLykPD8LH4XlRoX3qU3cT3uvuFhbA+5cEeBrFv/wkCKJ4XVlQoSLMts6SCtL9W5zO72O0u
RlA7xs7O4g8uywm0bIo7IGUjAHG7Wep0y4q48YCx8g0BlN8MwTpP+/pyoIv2rLf2qfJUn3iZ0RMc
Djusy81vGEDVlY+b/1naAW3ZLG84tFA1KQgVE8JuY5bI2y7E5a2oBqY2kpn7cjm9wSTMpZMAim/0
MmzSC3qUsiC4wOV/vMjSpSE254OpEafmLjSGOmJPgzO7y50Ja/jAzF1cGAmOZD8m7MAqzOFo1nPc
bZfOm9WflLiA0Gx+zCyqcnvq3pdKAJNgGCUUFZPzXPoHBBaN9nAaS8y3c+Lcs+jM/Iw3Bba7rE3u
eKmtOspzD48MsxzM9g5+8K5zix7G/W0JIL5Yq83LdcItDCTZr895VsMcsqBPTWCc+U8OBqtwGMOl
7I/7Q9H3TnAR9yBru5fG0aBgBo6PJxAipyoah6fuTZ5ec1fdKaG+tueYvt7f12qiV5OkNdOASiEK
GbjrtnIqESXkb7rliCOA3QNsqGIJRY1HfYWtPadNdduwhLiTxvabgkEO4Nwod6cKzNqq9+eJzZFi
+XY+lFuWOVQYsEkOwrLZRChjouoY0Xt6QDbMHX4NpFdHFtVxCgzKH9PBE1Afjbd8RxPOB+wlYM+I
oHOkBLCAZ9KVffeU3FgEHKDbWmktn7jFfvqENKPjwzBcLntqc5caIUURQrLJL98jtikzLFI3Ppv1
gcjPJa+VCn9anyKNY/Qg7bIZLT/yEPwzI/3SJhsCoCyOZqF26blNvecKo8eE9ZdaV0l42VtZXDhH
Jn4jLfXabUSgzQK4v/e5OkLesopFM8OvnjFWC9DSwHe7Z+jZx74nc9CDOyc7ZMN03PcaWb1VamYE
XTlWg26+BuyXIXwhibS2nHZa38uxSJVlcQdlUZ4g/E3JiDdqe1T29G5zu5RqpHtxQ2FdxYcc/ChI
nwlWwf3ZX2C88mwBFmhez2YVmuwN+3Un9ppQlkMqHRXbgG17I4ImOoO/Guu9mE+e+TkoiApGwm2X
7hRIHynwlTbemANUr9+8ZO/QIUq9eurKwjo5G1HFn5HImU5Kmc17D/FyEUF1VnIqeI0Bb60sSp8A
Hef1B/ovY3QhcfIZVn8uOh8yXpiHEexcbpF9iQSD4iqV6dC363YFL3U+3AbGrnO2AbugAU8PqjhM
mPIt+LW+YVjHX3dCWLdRXP6HGb120p0uEp4GMK78dLVD2dSmmj7YDGn/ygL+vT4bY9Pi4yDPyR2Y
MBYGwMeUMky027jAqgeYb9NADWebTXohf31dz4oVVoyowh75vKnxRU+RXh3lAUlrULWqi6Pc8nuT
0ba6E0G6kee0efWZevFqvPPpEQANW01DJ0ycP4b8YQsc4lf0hRtjAuW9fAMZRZtENF2WQ2SctPz2
iCyYP1aic96p+amscEnsmW7+zwiXSkGkPgzoz7wtm9MfCGMgAwVIUds1H/5wGe7OmkyjsMtDOjUn
R/fX4JhStDYGgZDr/imF7VsZ1nWhXssa8yDCEGq4p0RTTusAZ7tntq2DvUz7tmtOEqf1dwLNU5Gz
olQIgQIoppa7AuTfHiP6Jc8xaRKq5cV5ObyOHhhRLU9UKYCQkB1OFUGH6zdcmNujHoBTs85IAGC3
Sx8UykVWCqVUFyFEfiCj+sXr7DjvJLZezdZPB6W29P7XzlNJSg1IqKRgRF3uAmmbxiySOVoBYdNY
UDgADSuUUUdD0jH1Uep8lRicH5NvODVeXxLfoNfzXFP/NvFGnS3fKrU0jq+7Gr0Sc4mi8qew0nUe
KEMV/comjjGZBNHujQZB1yVpMNgcSKgBJQEfUmOAUSBKKrE9OKa2rLtI9pThHoEnnXrK9cYFQUge
ETTy+kaHZd5ilIcLHjiZosrCf87n5jpOL1xUO1GW+vjvrGngC3NLMlBKVc8wHp7y9F2Z0J9b0NoY
B7NxO4RKrnCCsnAJ4BQgoQdqrTEP7HAyKL9EJ5kUJ8vTJPR9EAYURAPcfUB+5toYDvSzgbSt3K+B
qbCub95GHhQPKOrUAmKb/pUjszyjkUeRN3bTY8az4qFoBXcuX/oRnL64j1yfAX1EFbLwljTwbvqU
a4hNcyCKSh7E7dO7VWvAouglYATstWo7jV6j8KcFO4k+71ExwPYu2cnjWbbfeWfrIpt+e8x4tx71
aRePtwZFMdsg+JfWokBuu5A6QEuseXlAAzg8ahbeReI8CmVa8OQMYQuJ4wreZ9R6nPwPnAYqg/lz
2Euz+X/e7K3U53WV5G+28nJpD90QlYJ4B7uoeS8xOuHuHp7F+R0ztdQ3Ta+D77DmT9EFb21orBcP
VRU7fBmHPnIKzweQeeWRc6XvhpSk7F/bOq5aeSe0icRVz07rEyzOrWneyvbNJAZsLeberprwLupe
bOXH+XqlEFziq9crBVIi8rF1BtV+K+7v9e+i1FiZSOPS+BfDKMemd+SReGGXtka5PQCVNqeBv/33
52xULYN+31VyL4MV4jXN72jr5jG3FgGV7f3TXgt6/Xohc1YKAO80uhPkykRPjJF7adMX+lgh5FI6
/TPk850sTnwiNzgA2HyFzrHjLliZu1fYkDrfkiDpG1DD4SYIeIrSukMjprBC9tEFUPBm1jMVqyHE
88uVfIrbWnz+BBpR+vqhAHipX5THDxvr9kH2BbdBeugXk2cak/ozQQgmBORyd4Kr1LghA71ZB4v/
WXyQMgbsa4shtKBJw18k2uswM8hGuPM5uncAcuIOhH6zGurWriJrPDnsAcTUt28oURgLy8wufOK7
0WLcd6xIAMj8a915Mmt9wX8EEC8CZoIx7Vk1WYXCqiBAo0PTdLtpQXKAZCq1kypnL4oSj7+Dg74A
p2WGpugAqbVETcUH/D+7PHHPrp97tZ32zP34oP0/OgmYw5nzE1FxivTX126okwS8QVUCUgvof9/p
6Ujm4RFzNgv9s3FsdVJ3dXsKyPSDlSMMcT/Th3My96w8MxguQKSuvXykMK0osP7KExsAPeHpEpVg
3BpahXaqRi4lvTNW+BSX9vQ3P3cg2sohd6Vy27Ji9w3Vd8H13ee/1j0pqblfEeEsJ+oo/DauyLhp
IXOl7f/G99fFzgAk92ICla7ReH1xaNCTHAxhnDT7LIRWW03h9ThQFPjAatt4Fkdu8k50gtWK62Do
ERG2LJc6BNOPjA7fwnSdXfrVLpSymFGtUTZcYHVkenaDgd6q9rmkHLgsoic9oaYY6Esnb/0j2TDk
WHZXNKCo1kuc1hnQx6+ZU4pSnvPQ+LZZjleQfn5FSiTpFkOqUievuuzjd0xV+yLVNNZz6kU7VO0F
r2wr1aOV/O+lfVxdJ+lXMYbntA6Iv0Yc1NEpPGwCAkNJhWTS7e9bJIMFA1KDcCFCzWm6gTpuYAdj
qkM+49X4LWRo0WOGRYzWLQF8FEEM0RKdkBoDDFlG95MclCJeFwYr67r0DdXgoHPp2jSeRg/9oHE0
rSi+hjRLboFiON5duvRLqMmrX5zh7WP0prgU1g0kiu2ijnkiPfV1hcPjGzNUoCCvc/iD/FQ9fpfA
IyhLp+laN0UcZPtPMWxQyqbMjb+oaeLycXBkS240HRV4kSRScMC/PsxZLpCqAica3hD5R2dMqrrb
9gzJXo6By7uOhY6YoyiH1CcnmCyBOeFaNjDG+qWjZIL4UFhYwAjljBEWSTSqXR422iqWa3C5S2VE
b32Vm/zaLODS+8Bp9NvIJzYOPZC22oEukFKQZWv0vN/xqYGquD/S6zqzaADges6hkP44+F9+R77o
H3MUDQgmRyiBtSTqLoNGQorwzLGxie0UosQ2EGj/ZiRRfFi8bN2yoh2LRMB986Yc2+Qe+wBVGAj3
BjJJ6LcV7AbI1KB2UNdFGNR7YxGRqzJ/xmysir4wIhYPMZFko33JChQ/u3CxdCCyk1PnwMcFdoQA
kRFe23Ni0MHkytg4EPuVAQs6jVnVZ2LBhphnYzNCz8+QfhCvRMwQHRDXmke7qvM4b7in6Ps8QTVe
E8UqZCxSmCygIkRfiKZw4a+I6ywlScIRhWsne5KXNDoZsnTggQrTxgopKPaaW2gSpzDV/L5m6YY1
WJ8vFNnKRlb/vaN/k9tBM/fx06odkmz7bzDS64PsLNKzWhuMxop3eqosPnBY1dDfztWi44S8RThW
lBgwM7ZYp/bH/t0wckMhctBLvQMxuiZn9H19g/zN9CAzCZbKi1hyCzSfg8K2OlpR+eph2IgnoBCx
nfmwQ5VapgND/7idYS6Jg6p8wh67I5/4awhZjAK0uap8oYwVesFt0XXagbC1Yu7Yh4+1ZrPfsLdp
cjLAITZBKSKCOnFGWP62j+Er6quyVkoVxCzvtq6saFWsteZIK/MUB1v2AZ38fZeiyFtX6pEzfW+/
l2XQ0OtaYqUjF0LYUoqA0XLNgVKv353R4ZGr2Xf5v4J/7oLgLwEBdbfu8wlTviotVpNiRqhZriFd
uxzsBNu1aG/KjQ/oVeZV9CoBibM7jcQ3oFiWIFncAeDWAFT8wlL4S9ObeTgjUWfyVQx7HOCWuLYz
AAdq+Ka2aJa3cSYDj9TGzPGtypvr9vPDXU5WKfXKyFZ7BkJW6L6r2GqTe1Ex84Y4pTwY1+r08Y0b
IR5Jv7EuPRKjaFBtufy1DoQuVC0xRGqI3D24vEh3vEqFQklY7YSUwofXIvZWX0ofPZ6AafIkml40
pEfyxTHNc7Eu10ibZPZtnkD2NG0SwAc+qmh4KQBNU7fYHQZqemHO8iExQbSj2CWQD2v7btdFtECm
MOZGPzzCZ8J5c+5Q3TcBUZUFhTnTDFiXp4I7g9ZpfFJ3EtsyoV4NxlJvXzGHzRW5pYG/GeJhiNtr
ZpM5YCeVzI0AJQo9aTsVQQ/JK5OkXiHXJr9sz2ghhw84VE+C9FhVx27wYmkZ/dLn8Xd4wKhmUwnL
JtLlq69hnAiM5LIwe+2+8fw1BOyn6KWukFGYgje/RACLA/D6sNqwaCq9xYq/dAJXoX9lpJ9seWP5
g+4Ur+W0Y0EuEj/hQqt9h5uengAZa9VpPIp80QzFbpkCxqZJdxSfgkl2jjlClH9uvGFlY6B5eIT0
hcTIxlzMZARLFzeNKvGJSUMr6ir7CgxrrGlWtwH8w8hHkQSEWNbdRcny4qEJvi3c+If3wKifJ+2d
zjoED6H49N1JMNhspGaUyW2R7eDxCDqPXIlZQvByuy/PXVzsIz3S31xwupNcC/hw86i/84OEKGY3
4vnPbPKkoQirpmr3bFLbtoTnGoWfZfedl+tS9XepSMka2+X4ThmPg572oUWFqPG7vsBZ4K6LwhnK
IXYW4iW/Z4RHf896g86o6xNdUX0nIauOt1wF7gbkwaxa7Ee4HkAD12uKusQlxsZjkgoBR/Uzntp7
MCJGpxqKcU9hr7xWU1+mUdwkhyuMPn0SFjfEGbtLV3Y2xrmyQpqmS2l7bGLdWg/7/Rb7nBxy1DME
tqyvqfjIq31csExKWroP4fna8ku+f9OYI/+8N3gU2OYXN88j34/sthUl7CrQNPc5AI1ZK6W4l9J7
od5a0xyurYTOCZ9bZzQsmPa9VAG1kAl6sZ+MveZpM9RNuOK80E1VSf197xQHTn5TMR2PePTJgVE9
oPY3ePOn0GEeNpZeVLBXSoY8WODYcohh64exHzngSltJbblX7ZNCutoBQt5JZa2NXVvBAs/i6+al
H3v6ujzE+/QhsVLfLOjk8hXM+15BJr8jhBH4UxnRg0SS81K852xcXnchrG0TBqDU/Up0YJc3f+VK
tgwJBIbTMMEZJfLNwyJpi2l5tzcqPQ/HOm9mizN1CGaup5hBXsqAGJHotbUO9Ba83XN2gCL5m+5+
EFlixy/uYoMj9cfedl6tV5V/d1WDPjdGnVeKCmta/DYDUecwg6fzsDd+OUI4YHE4bzIZntn4B/pt
8H/2W3mdJkri2EpGRBHqgvaS1q1mHqRUsdt1R9fQhJXvA5IG5cHuDTzPyB2IKLxclzKhvZuAjo0i
AumQeSdNHjTs3hfmPk9+ZZEDh/uE/Vs5IcrWOi8GF1MensprNV+Y1h3wcJ7hfNntm/PAMcxessYw
7KjR6C7VkwwlQJMQSG2kLdhRh1s5BM3RiBx/CFZZSrap33Q1yq9QHAxzbb5icJ/v+qT7zDYkgE0d
88ESOwU9fF0gXHbn9HFPppZxaLcUM95HPZ1A9IMzd+Oe4da+Rt2pNPADcchvCnywl7fS2G1dIPHO
V1rGxPIF52U+uFXZ3yDEkyjirUml+5UUxFeoXMk2Shi0C1zhkzfFcPLk1TwmV3IsFuD4Y7kDESMq
7yM1R5H8q0E+QCxLcUMtCF7B8XEgwl2JTlxjqRECxWvG+mLGtbd2w0uClaaaKozIS1Bk3HR3UU1V
EZPAUtPKjADFvpWvFO9/e43yUCmPyRF2yAtMn1r1dJ4AeLwmOPWzjDP08fhSVGIPq4te6Ra5S3Gt
UwDeibEFO8S3OadgCbLKgQHr9WQ2iJ1QvL3UIJMjB5WTzh08rl81fhl6IhwJUhcnDkXjnb5Q2OFS
EbKRt43zFW3FQ8zMi2K9hyNWvd1y9iOBenrA6ax7emunzaZH/0Y0vOuN2yDCTZVh2bA1oN0dtkWp
82g0f0tPuzLpd94bMPBDkhQTUkztdY997zNm1+j7+WzgWwYjTVR+cKK6F+xNAV6e7qC29wSMY6Si
cvaFgwCkORFUHX5yQGDFtxqD3f1ATK1vtml+KLvrzUATxb/dXeIruYxTwtAKMwPTnmmarkVunc2U
y6EbZ9e3u+q+CzLX93LMrIjZFdYUbxcxUelpQuQrJrrZsP9gebcAucvFGHAwvbCYGXq6TqWEGp1H
KIP/h1cAy4YgNPrNdTTiufYLgNNpPZCuVVn9S2LSLIv3DpHV6JqWjipwhexjD7fdoMxufp++qSRj
9ZDxpDY34kMaVmcY34hJ7mQ7DZIG+RKOyzeDWNEilsl+XHka3BmZK00E4bl9WhCyodAsJDb/M/C1
lfaylUYH2NP8GqrycYj3uQfnOCWtXpUEMjg9L321r5KqBhrS/6TZ3+Q66B4HuSAqm44uDZdbPOWu
qhzmA9IJB9SpwnPwqD5ap8DHC/JFamJlCrpH/GxLnC6uQglRdl/pnn1aF2lHp6ZVY8yrlWIOqyAm
sJIlf5U4n8Jo1F16T6ueL4cRxg4zaKDN1AG6cnaKLMekB+Eg54gBdraBM5CxNCCZV+8vfnd3W+da
ORuAngQfAX8Wl8hVEZRF5DtMf2d21/OJSDWYDEHr1WA9r1gCodWfYiCxB97RaeLSOIfrxEMYX5d6
Tp9gj56+EqUazbNOrdDCLgMQHehAf1WUfNTeUUltxvgw/lDbe7yxAttDqjNXl7JLRtugsZF1XPaB
PH8K7rxDK9yhQ7yLXlUUmTR1+Mh45i+azKpJ5CVZ1dcK58Bsp+6vw21PJAB/B1Ok0ZWXQFCTphfK
Z+/WiFCSMsA8raOPZb3kTaxli+v8+3CZd32uWv/oIh04VxTL63vWty4PKaTzcMn1hh5K3BmfiEaf
BvAy7jm1c7cRBa4EyWhnPkcWAhzAA38L1YCQu+BZCcz+HUfndprdqvB/rkT7z4DoWwrgTkpQcGNh
qxpftC8DAC06v69jrQE7Ve6FFDv3n78DR4ss+GkzsTdRhOq+hjkJk/czoujPLliVNixTVvS/yorB
jCqhRwdSiw71aRIxAZtCRCgPYdeGeznmCsd5vY7XcKwcizbGrtfcuEpoAzxgZLdaKXaqzjb6ZjbR
FJO7PYUNwgt7N6vnmOhLHfCyZyiR2E1AEylXduNTB58ZgYNmKlOjlwX/aGlnKOq99YuOD5Z7rWvV
LrHWwOBssXOLFW0TWYDKdz5XcrNii0kbvcYOtaVvr4DdOHwHz44eGZi7fOJPQTr5AXpPIeG0QhkG
QeGNkGeM1NB8ZrVaIPqXNj/qxFb++XcwiXehAehereSe6weFRiipffs1rjecbBWTBua8wz7DqxlE
ZkQOG3gR3wmllO+zfbtxdOQVlats9Y5LNrhlDYKwnk1vGL9t1dXN8257ouh5uNGY7yHRehXwWnAN
DzeHH7aTAqvAqWpstJdg59g8Q15TcZfpMnmpMMFOULZeneI+a8a8kOe9qdVSazRv+5takQrnyrmD
SJvFSj44FNfTNzk3bV3zLBysXpLtkvEm1+Cj5MfXgA4j9dFOxPujK48EPIdw05ngfKh9ZWwAPVgi
D1J4xeCHLilApn7p/WpJkBY9HhKtkkxO6Rc3/MTGvDdSyvf87J+jxDJ2o4OjQ2T9g+Qm1RcJhcJF
wKkNjaQw4zGk1Te4Kgdq2dmRZvcy56oAvi/tyfFyabvjG078wQb0EWSbKPsq6Eh2b3KbNrlGIeJv
DvFP5Mo5J5kMyXdbDhTeZOFcAdpsl7lzViWyUD46O6ySAdUqsFmIn822jE+sZazrcW8BnynDtxcO
0WvV/+Upwf+m71feKgnCdPnNaAsZOOdYC49MvJwJr+lT5p3XjmGn5jN++qts6Hl4ZXN6l31UtRiq
pNLRiEEp9nriK3t6Y6dRgDv3EZdahVv+HcFoAsjm+CrNgNQFHl3DV2d/rHTH3/s1OY4rNf3EDZ9R
031kSWQbQz52BIcm0s2LMqOK4EgyhucO01+uj960N8V+ydhfSC8wnaIrTt/H2v7KMxxjuE4Kiupa
JHyf92Nf3qDYQtIFhkTCaZEIjMLwGPhwCGFZpiml307y27z/Q2XJm4KBs7uW7TRkfm319K2bhl1F
DoHU3spIdmf+psffPyVVF453TO2BU8fx2zJV2FdHGYbz+Zr7UpU30VuNsg6vC+KJU6pzDozg0r5J
gkYe4m2eHaD9PzzVp8q+VhFtj3rmm+Gx8jVQzqnGoXMuviLEIWG6Tspe8g/KAt68Cgru5dQFBTLJ
n2bx2diYV9NxCYuxnmLwUDWf4/nT0wiI63ty7/iuGNSMdn3Gz1e8ov1HNOnIv3Yw7N9jyz6kjtRN
qDbVRKxlhmNw2vaPvtFDVZ/NgINla+6V1Vvl5PwNyDF6QgUB2oMmcQdH6QUotE5dIsYHhTC11Oq1
vm4VhIKr2LgNAI0ZcKID9KbMS/9Z6GqBudkphhdnr0ad0FHt86Y9MDXRmZ8DUKlAFHUAhtPJowsc
WABZgHtkrUtEcPy6uY3EZ/ISOLALTAiqoT7Y8QLvzfwGs2QhKK9MN7Ej5DBeAeVLowB6DUYjIW/4
T9eCiK/rxKszZjrP8q2T0gaZbCAqVKlnVCFii9MT9lLPAXbjJNnUjhNVmGGJ1hg/XKKOKDsxMxPR
ynuQ0eSfH26xHJ+l1bpYhswrwktE7RARePBBxRWD7+HUNDYCCeViFJZRKXAvfJ37jvph2kncDQ/I
WwbDmlN3sQLldrl8FUf+4vvmXLUo+GcuGpen2FheRKmrOhZDUR6SPPVT8gaA9KIJ+aL5he53Fyfu
GQzUrz2ggQoaU6YweGX/eghrS1d+yCrLE+46UA0fD8NmYAALpnwe+tjRTh118wWVM2+5QwzLO8cU
+WULzfHI01PfIrJPFZxtQUpiA39Vk2/VET/Dk5H5iS8uaIKKfb75hfT/ScE/gPx9vhYzPNMQwZpU
7WJ6LxdowCGVzBoZzM+ERIhc8hL7MelOcAK7qH4xU10gt9yh/9osl9vpfqzisL9AC50JyDm9puwa
PKH8FGsPeOqqUKwyHcY3z3GK1W3KMXh6ISmEebn9C6psaJ8R6sUON4eiSq6uNMQa9XD5WDH+f7xX
0lJGeFahlnguGW9tEWpK/lDE7KaZCxbv4+9p7nb0Es1uLAQo/kjLv5mE0aRaBu1sfxZ4qp3wlu5g
B6XtQQuqdaPuBPIPGhRuvEKnepdFIFreN23ipATkyi+FV1fXWafejIVbK1U4cO5qMQoJ1eQda4y8
DZa2WaE/Z5GrlRwHhBCmFUrE2cNDzzsDd6wKjj9fBOKAn/cc2C2C0w4BNdQsUcGgO+AX1SGuuxm+
D1HwrnyPKlmJvJJwbQ913tHrvuYXIlus1Xsf+nrQG/pnEUlt5unuMLUMNHTgJabzeXVyQLMnEqfh
6M0pgMSavI3RR5EvYSD01YNE3MdB77A5AP2jBVdqW3qBBfCU2V7ZWE1AyiuaL2KIbufaewZty0m9
wCC/+mY107+3Aof9OZlEbRdFsjsvBLYYcDKYUwVjv7CVP6GPtDcSW4G9Vxk1D3+JQfdIegDTPRBe
Dsm72qLLkqoe+6fo6Tv1kqD0T+CIrJdKYRpyR/vZ27H+nIXE425FdqE9PHvASJ1x18hnkV3xwb7t
v38k13unWXFv1ZEQDRlgXkFkGrI60vvYSP/F3ecFUkZs7r2QW4Cmi5MCrkHyFeLQUpCiZhIdwtqA
JYpaOszESCjJIedC96Xjtzj3e1pDXWEh+mvtOmYVM9j/mVPq0u53sAlpcUZM3bbkd+l3U1zs3lSd
RgG4ITqOR1PM6bVXhAbDRmO8c13TYbRwPJv5Ry57nNIUxUQBsxFE46VuasXolsVjqovqVV9l1XXy
ep4N6fulaWdXJhvyIdf7/NyrLuiUojddkV29C0F2Y7tczY8FiAJAVSqjPJ0mHKomD8dkeCn6XWmt
vn41pKaUJ1+YbZoQx3bwGaACdtYEVcMtd2SYNTlklobyBenkKg7VWMZjvAAPphekwVnmjq0xEVx9
0+376qLXl/vDiXYu9ZqpNHUyYlLndwlZ4qUzie/3IwQkTEIP2LIVKffdsLm4hx02tkzlFo3y+2dS
XNiHDgzB61Ru5p1oUcHLtfqdipfMTfxot1D3OuG7V2SJIEhM+i/1SMvV1ikikZfxUShJT8vZY2pf
Re0shhC6t4nuPGeFiQr3U483KlNvBh0XgNScAjJapmKThi4MlnxsqPCNvV42Or7sG46O+wuxHoj3
cs1/yD5lfveB756R8nghNeTGByw6N8OjF+crbeSuj8kd9/faIelxt8BI5Bao5mGHh18tUEA71Y0U
racVqz2zw1GWwkyhyMhg/dM1IYk325YGDMWNNPz0q4oTZAex6wFLVWnx/val1vhkyPSItKfpvWg3
NOyD/vh88+XSbK+Ebs7prR5M5F2c3fEOuD/Qmxf4RSrprKxIx2shrWmww9DEsXXiq6J6ILkUBoQf
eqOayK5etwggivRg4rgZjRFRUPupbOI9seDakWIPtq45ZZfFImwy+qOXh2zWvC/NYQ4+PUvhilhT
J6N//sQtkpghkwlBr/mvAOE7/gp1P768smSHPkOFWxcCSHhM6DxJ5tyIpQSv5qaFl8Nss2P3q5Ut
A7bLWFmyxCj8PrFH+Udi7YRInzEBiRnOhCRXAQUIIa2s1d4OPbJW65ECg5szRd9JpkLLs+OoeYJm
NEHcPPaaLoune4AU/R+ixFIStE+kK2etrbPY+v+g2h5NOUpNms1te5sQ+1hSSbz2XSZVzJ6K8j8C
H5kL5WTugS/9s6bSoKkDq9dz6lzbsZpSeFfyu3doMdgqnU9DQujCvSfoVyXdk+K3cudGSHrxjhX5
ahH/pKXo4O5kjF1jA+VT0BlyuVyPM1fixROtbt0LaoAI4VaMCmJFStSKb0AU3LIjiVwErQ7QiAN+
02hTvM8EaO38AfIAyxXUtIW/gSSqegh9L8l1Atw+vRyYtVs9sQ6UX/k350NmJ167xbG5dlf4k+Cl
RIyWgTemHq7jcIQjNIT/JFNLQitx/HIT5bO0ksjLN4/yeg64qewVy7IktXQGp5WntlvXY59KlGBo
zzx4JsOIECLRpSZ91qsd+eAwTp9k2k5rALxcWBbQRSgcW6m8XYmjrsFQAdzD+nRR+aYNHCXoktD+
jqr/ezRCIOkqqY22knThqBJQa2Y2d+K8ncoJ8y28jpx1jlxv4vc9yJJzO1P4wuvAWwzSftshY6p3
RFiwRt7K1zsbQujM/Cw1+CDerpQvWn5+PkX5+9wmj9o6jdyMs0Dp/CTd7n9Pdp9Pu9zZ78jjmkcT
N8UardIF/vWBcDnYyvLmdkp3IUXQuhiEML88zaR+qZx+Wno0LKGlziJ7haun+NAZQpEOt/5e+Cyo
N0aVjgChva79hU1PUG1+lvYmB+X+6jNB4gqbtESgG26a3YCCO+MWJxq+0D5FWfc+Nl3RbjU00r+Q
HvaVO3c6jFHmBl/qG2ZgqGrMgSdKbKLfnfq+7H7TNBrQ1PPXhaWGJtwNqMJAmQVK1e6Mpp4G3csP
2EzzKFN9cyte4YdV+NvT6u2iq+ur18Q+oUlYcFeCrxwmVmR5lc82mPtVBEz0ZLCfdtt4Bp9J/3Te
VC9BpmedYZ7ptN7ZNuP9UrwvLu8C5TY5bK2F5GyM2R4gLkIhGiwOTWukaPXOpoCkEtHYapmXTIx3
vwxoUeoXJvePbg9F3pxpyztmsczI2U/WgXjoQdnrV1ty7fHowo+fhwR0ytTYq91mYS0b50mvmzeL
spFEF1P5ohr8xsX5SqhnnXt6rb2Mc3XSLz7oV9iZnS+wtlJGO2lnoEeaB67OeR0CPOucNNTSSKVR
mrhbMtXuRtpRetCnStp6057WPuXRm73IdGdKK2kpfyWILfJrgEzQClD7WK3Uvv5YQ+DjrbTr+YEF
PeFqOSu1hQ+S4JbVkve0vy8ruTHn0QZUk6W63iOiq5bYsUzty/8vYP0X2GE8c6KQks9AmksmzSFW
AcmFI55lo5ESmN0YnHKG7LCJ/yvzJgjNC9K1x9qn0qLYAj56jqtTEjj3zALq5WnpDgCYsQZ3WD8F
Ksvl/CAzW8Qx7WMMRfSGPcZfaoBruGrZ9dUrbW43L1U8uQWwtGYc+SUw39XMMuAk/X9jJfbrrDFF
XYjDOwXb5+R2GoFPjZE6m9WySWlauz/C9CPN3Yrd1380JKLRjMSr/AqPB+cVVFQKXSt42RZ1SLht
0Qxm059KRX7+uvj7Gtq7rhI6WNc2XbzK4mPfRqhXhlAZuEBUjkPg0b4rMM1atzvQYZHN1RaCvZvX
ZtA9MLboIjGnK+GYH5XqIJDebuPS/7XMO6dWK0OTK9wDjY0inGv1vq+RO0vbr0Ae9ToY17lmCbHe
eY1azjarnrOiFCWEYjJFMA97TsqErYhDDK5ixO1IyMCxv8SJPH9Zyqg+57YsCoN80LwTImFhJJqx
V87PRhO62zfjwAVPZYYrEmEoB0X2Yjvy1L9dN4ZOYQD6waBQpW+vLSvOwK1+A9wGYSpSSJcQ0bNX
oD4XDPDkhwsPeEagSVlLX0Ib4MHCaHR4sAShGFL6PJhd49n7epBPwOwzIahKSzQxlEUtVru16qjx
3tuMBl5zhJ7FHw4KsxOuFVHN1Vlfk/J+e/JI87xlrNKtvcQrG95UrYpCpoTmUQqRBweQFoHtnHY4
+SHqE5Ww/7A17LUGjEdB63mp0ffToj+W0pIfN4OlHiK8qeV81rJ/lCgx6i5a2zQ1vKPLohhN0eID
9PNni9P3jsrgYeRDLH1XBf0uueTTwflShvEyqAL9kgWP13E8CbuAJPifRaZNuYgQ9vd6vgPb3BmK
Gy2RS5T5mqcfP2d3keSZKxr73hELjSSVhgIxiWRLfjAa5BxaWJcuuSUia8s1zhy5emknnQhLQ4iS
OYkDZFszl4QTjDPah/Eqy5RAV0olqs+pNrKs4Q1KyJrs8ISvHEiUpHMyA+NA89W261ank0l75NeH
jRKnIz3bV1RrrAbElaJMXYfHLD06fhRw744UNk2p/LpdmUrsoU+PoQ0Y3apjg3ddOCkhdSm38RfV
xq98tnsurxiIHrWw79zehrpfwf/z1uLwWqVncVm6dLjQyhBK+pH/FNBaboP2/sQo9g6AgnM5jBPM
sku0dfUSScVpcouSV4Ovy7cr7558PEIXmTwzEiMqFNWI/UDMA0OYMG+blA4Srx5ovFAE5zhRWe5Z
FfeNwWxDhSGEB8f9UqDb0d4m9C8KH/2N7ESjImGCxglaJkiOEZgZJBqFEHeKAfNLXu8meRuF5ZhZ
kT9AHGwJG8SMcpR/bDPc9N/bltirFpGgpL4kZP9D7lixx1aZQRhPCTKh/tr1w0nzadjvP9Fs7Rf8
j2eoLg7zfV6DlR9jkpsMfEMUHZnEPbsHmIiKM4xY/fYkMlXGDgBql3MRG8E4GS4RGn1WK0VFl2Vy
W86fSSEq17noTyMs/Rm1rIv3UgeOfrTMnJCQnioDJTifzroTNaweaS3HXuam1cpRmeziU8wh2+Cf
KN/D4hI5hokyx0AhGrDOF9CEUly0XC+NoeV53BN+YSVH3BSGy5xGsKkKJWSTA8iVTI2z7Umv2fVR
ZItBWmZ9tVxQKbnBm2+HJDZi0KX4y1Kvpv2D6COa2zqWcksObqu7KYUqOlf9pR59HkW5Ql3rWVQW
VB3s52lWbS5dQFo/5umcV+oopKSxnIhnNkg+lo65TcoaWHMHqOjg8vbkLx8sH8HIjU+l9xlm9Ny9
GU1ZDeNXD7F9XsXAXBToydn/xgZNnhuJ2l2lnVcACaNl0DwP/ENH/t7iecG+jQRQw/LWXkO/JSdd
m6IYMH2AsoKduZZwCcYIkLb6Ct2NKL+fpXS1xXSovBE69w3+p8eEoqX7yl25if28M4TslUDA1WAn
Evr8dAjrqf5z49o5MRNelaWP2uny+3r9Eq5em+xY4JpDjot3r0IuRWZV9c/Kl0uQjEk+z5BE/Xmk
3ZXObpWu4Msbodi7CTbxgQer1VPGuHH9CPz+PRPcxJIXAj8GpAI5zoC2XzZT2zcidt3iQemkY8Tu
jHG1vGVNuBk+HzTJbYK9h7F/lm3y8ehz8ftZ4kKxCElTINUcPALq1QRlNn96QOsBjAVVIurGphe+
jbUv1r5UTkAH0mHodvZHwIOfp1qzYIx5DiKE6UzucfASkfHSty4a3SHz+Cop+N67q2tkI0DQDZL/
LtiKaTiXfIqk/ApJFhKLXMQqwEyOjX9gWd/jXPArqUP461fkZkpgKZtiBG9q1ioR8RUcdg1X+gTs
3RmhxvzbTsGW/v31hS1Z8CUJn8G5Gk4oolp/u9SuWav7KDvXR0xGQgof1zwPhuCY07oQ/ThybY8G
h5vRztgL9D6BbQEJFH8+6aZJWdmj13G276e0L7oT+ZsA4AjtBwEhYrtWweOKzLZbh8ACumhE0fQ7
HOGSu5pSMg7RN47uqs9KMJTgc/G8rJz+yxanL2SRK4igAzJ+NwatHMYFkIkdIExMWqIaxaTrYe0i
YPFtLkdP9Kmpr07HnOQx6H+ha+4DjUpGP27t7nVBk66NLE3OI7xhjVt2htYme6uyeem8/9E/JLmc
qiIv14C057f4kwgyuvx3Ak6B+rgCizrnQ+VUHTjNw+PyNwTeziAer7TU6MRQgtAH29Pw8n6lcYIU
k2p8iSBxAm8DX8jFanp0dczSWO2t5sppPfova/hjEP7KrSA0QDcM/tudaUwLYyIfZgT4dWX1a5NP
fg3JVQWG2LYG4Zvk3vP+y/1vpUZ8qezuYJH54ZCu8lJVjAILEX5AUhghR9usH1DWiTAuZ2tbqgdp
6jIBVJyl1pJmVglyCE/OWWf7CGSGP8Cr0Z4qOB82PCb6eTyTsm60pNx+aX9cAGBI/kBq8cSLkCKC
NF6sh289Z56EvcZD2hbFoZHflCnjkPIXksaqmo+HKMqRHlbR+JCH0q3moY/QcApN2SeGxwCBDIZ5
4QPIbBjARelWMQFFmNXwF+g2EgrzqyynHpUrzpuEPGzxyGTM/2KIRFw6oHz2wqjCAQocv6yffVKu
rvRlJmWK4lrzbZoRL5CejNM9pBmnm0C0dlH4jBkAi7DGD99gxvwiJyA08kkBGbkgZvkkzEwCrUTP
MLpjmdvo4iz9dj4augvyhcoYS8NGjmARLRQOvzfkaMlvV8Y6cUwHGdMOjAKuSEIBu7V+JCrtcpav
R2sQ8RGe1c8ILhz7/AZfJivm1a7PWs1ag1BDDfpb4GjAGPGeoRAbL6itd8Id+HGL8P0aj/bcI/ZN
nvkSpg3Gge1y8MhHQGY6tj4M4ovlJAUS2qi6x41Vo0Zotr93ea13tVUpfh3iuMgWWpFuQaRS/t3k
bW/Qme31LAew4mCRpb5mfnMd7FZZ08gY6q5jGMSrQDTYcXvyiyCN00uK97w+pMXvpywab5foy0De
eTx6B6OkNAjqpgaDqlW6TGd59lrNrE5XMgOH8gKbpvUuOvx//beSNQ1Qrm21r8asKv4z/jreLbXN
22TsY3UfIw3bDP+9xJMacmBkIixSXM/+OooK/lqHnj/qaH2v+cAsMhS7PU9qbYAx93NtX7rySASw
y7BJZx/0HLUt2I8KMhXwVmaI6PBwt1ZeaIMWib26pFThC+s7LLZeWBwDWFLW0guGWZ+nnWbynf8m
plr6HKVrntfiZK9k/NMxSO+epRezfZkO3ey277lXLJfqFGyZrOXugSE8Jfjpkzsvfm4F8Wj3TQr1
lo92uBsDM47Pir7YCTOMynFNRKU22yVZ18BFH6uToAdfCK0pJee69QFNi+hQ3jDRwk4/vYBaWBMI
T6tq850mSAUdimJWERvP7Mqy6/kghHh7xpf2+6RAV2GOeUG5d6etFnQAbqir/0NlZLiq3I5/eXGe
7+pgYFLLUOlUTgxCt+ztltqx45NkhBpTdHhaJHk75wtmkXW04Xu6P69aOXgN8Fxt0A6CMA/Ebvhg
Tm0pHzoCikE4CX8bce8ryY5d/yRdjd3pxltqXs0gTmC8YXYgtxA4f6Z5R80ofB8a1k3ofljA0L6H
RcCwtFwNRMoEXsiqVzGQSThrBIUCk7RLNn8zJdKeHaG7ft1gfhEfK6E9RS8Qd2+oL9Vh3oZk5Oo2
ldGO8caewbzL3zPEhoo1Gxwk9zQPpXrP/E6nL5/IiLd0PMz+5ks0nnAlRnJCuo7MJU7UprgZ055n
hMAwoERQ0BuuYO+APA0kdh4L5DoTqqaI276fVY3jGOgcwSX2EmXkyz7C6xUAtQYADHnp3sYiYYOX
VynlYfFB+ebZsCmxEAW8tXeva4nKKk63ER8Qg2l7tOk5G0Z79xJpLa06kqqEeSbnWGFRZjljDR43
HKrQETey5h+EEu6Mcqg3DX+cfIJTgXLyhHHQW94ypYDwy5yjg8Ar8DWTfBNAPwn7nwPXTjuCLwNy
3xmlYabhwf4wdujC4qpQe/Woa34vZCZkN37aXMIF4eC2MWG6mszvIA0NVNHlTHCz+SV9hSZ3G6ko
+XIFf1i+xtdfJPBav6qD3p8ySpXrzDGRdGJbfD7Ngcr3jJfQkhI5xMTOGskWlZBSy7h/5mDvba6d
n2hv/7WHJdoOCDvuptPCatgc6rzw2njbIR0xPpdXfROkevltJ5UcX1B/At7GcIUpfekAU7/dbyZN
+Z51KMfJVbqarQc1CuDWFhAGofCa5RifQjcBxGlcpWQd3XPO7SbmVVRlyIdPBu7rX64oshw+olPF
5EE1w07hR3v3wbCaxWp3PukjNT0P5unb/46wUw4AUsPezHkVKz/aMeFHzCxxV+0LOE6E/KyQ1Vgo
zcGXjM2rtwN4o9qlGqE4S3n8muI1yzMe44R1DmGbMRC+eQrFYLwO7mKrk+NJF264BPDz2Y6Z/SJQ
JUpv5OOIvUulMiM7eOr2NDzbSG1F7kISN4KpxQSsglW+hRYx+VvPuVZg5uvFpYMHqZr7hBwbnmNv
V3C2umnN1Ahl0XOlt/CJqgqap3yDS4u6bX1AG+QIRu1KulJTXf28+Wa7JLyReW72dyySAUk1Kbsn
aq3wSGX9nXwSJ8TQcaGp4MLcLkwxFuD5PAvPhD+xh414vmzuQa91zLGxHfvxKf/jbznFyg6/SG3r
FgDGKCd95jqFBlaDuCfGJovO6kiilOPgf/QShsjxq4ONv1fM/9spM4Q0me0EybvNva7/AXgOQqyt
M28sK+rFxkgKP0B0M9erjyHW86qRHl4SDzDrsKbrLHEre3kE7VzVnJjaHTObwJlR2Z9+qBKjLLxU
rVIMwfR7tXZA+gWbL8wSdrPqJvEsALJqhswGQjq9bCtq4a2gWG9HzvvhW0UEvY5aCRkndV7OiK+c
P2HmvlBu0pD4nWZAp+5JzuNVq1S+hlLnIhyUZifinPk6ZND1lFSX3n90za5bhX8Agf0+ECDbE5PS
ep6LhwZtuZZCvLL/iOGNbzoMmkAvDVXZmuw2FSLqzl5JUGU5yJ/78Li5K/6+IfTCqYPfLrNfi+1B
jyNpxD4z3CLfHJdv7ZsfaDPMFCI2vM18/dZM9V8wCw7mRNNCutU8W6a1HHe3dp5oD1LsSpUrHJCP
W/L0nd5kcrr/zywMZFLeTtV+uH+et+hc7EBg0nFe6uINO3/5NmkdKQlWgIbH24olnSOqH42wEm7R
GYVTRU+dhbaFmJ1MEdD3rj16SrDUKU/XrTEzFbEChFbkrC3YFZRVKBl5FttWvml24I5mHdd9myss
RN5AEgZskTBt4ODozZtQT2vHZLGO16sg8YOM7/HvOwvuBQC/globFoxtL2eyRWgWxA3VFt6lVwC0
a+Ih5QrR6GRUDbzI39fHQknnXnCN9FgMVl2L4t/SvOWbJMu2j17gFgRUpyRNmHpu1F99h+ISD3Pp
FhZpNQbxkxcmi9Cjv80jV7lgbffGPfQ4TS+0TjOpzVZvOiP+LZn6rajC5RMeBWLR+9Oz0Uc8EBhV
b68RvDCm9vnQFwwzBaiMsbleWd9lELJCNAROboEl9VZ5ZGg12Jc7b2mNW8fFpnFHlvSiOrcM1Bln
TvEqZDvODsHFg/d5/hpRgehg1sdOpHosHR3m8rc5/2rUVKgUQvNlPOLT4aCc2k5wPrvF+dA56qO+
PCn+c/S1UjSuYGSxwrS2lO8Rf57UXfiQPGRyqnfYx+oC0+tCjMPZnn8/p+dCCl7zQQTOEeJ/DjoS
EWysyXal4XCAXo+VuSLzeuwQ3WY74d2IfdS95yy9moDOmbox3yQYOUPzVApL9qusJyoDyuspp3KG
n43WykvNbM7vm1ZSInUBKhOX83eTL0ZxO954NySZOeH1WjkOVusJaLc0TtybOa03mGjmyQPCJM1r
M7D54GbX5XTNhZUUBlCiPlDSMNeQGESPbUbZU0phA7VFNDUAA2mrC18xuLKoDtsArJZ8AKkOMusR
/iQx71XRB4+q+djYMEgoMwIX3ALkb36LEtnES8aVvjLlu4YZ+H/E714+qXJfnzQ8/txDqTiNa+Iy
s+LiHWSts/srUYEoohFsrkMxVnZRODW7szrn4YIZ+QAR5TsjabCDUWp8vGuHDUO0LWGfDLwQC2Q7
GYXFUiFVOVC8YjcBdGSRV6zVj0AHm1ob77zLmEnXQ796TQkceLyjS8EX4KjtzprSt5trvgBwWasZ
u8iFDjxXajn0t6UkC0g6tlC6iGlW0EAq4LLh5ijpMBSP7DRbbaEwqZ+MLHstJpdwQZacyWSCZVho
IEJeEJ5nrznUjqpdiADleF+1GtqtteuB1E2cp0UUys4MmJ7a07GvvU5qfOnrygZpnJMU0vT5kl8q
dBJCUMnIdcaQMm8i3NiVCgvT/YE8JsKWG/vk3fD4B3LQ9RqDWPlGHI/tlSS+yRRlCU4E3s5ERZIB
qJgYFX5zsUZz3yQqfX+GoNpOUd+FFFeiUoUX56pHeXkOk6TKcb2BkhOgVR/y3XtgW0OXrJPtZo0V
cv9hl1A4ucACldxGgzODVlO9wFEPdbL8KxvIZNCeR7/f9aclGOpiuMztbcIJ557UXyEijj4a3rTk
0D3tNbx2jkwNQVDXUffLwVIN20aHqeEz0aj0zSzlziDxLmOog59WWxpRyD0x6WU8pDUYxe9sdzfm
Tktu3JWqkuJrs8vzWxWPvK2AIeA67Zg7oECwmmtU8KizjnIq/K4HmxSTf/cIVuGvjxQIn5mWm3Ox
qRgdZ7Iq+cuJl8H5Kw2pXNMlME7vzr9E1KOix//9A4VP3e3m4JnzxK1+2cjA6BY2LVMQEiAGYWt3
XLTvXo8VzYrVm6NPnyaW94xt7LGzbGYpJ3xNbdeDmZXVPk8zlQZxtuYgpMdkfDChndkl3WP9x/iK
ln0453lE+U4EqaPru6AetSmdBV0chE4Zr9/oFF2ukt7ZTW/Eg/JlI0RmARmmFOSjD2xeD0HtMC2B
9W9ezIUYeTxN7nc8ln0tA1W1CbOmmJdTJjL3aYbP+8IRC9akn1BUSFgty6WkcZFuC4BEGOQgn1OP
ByaqMDjSohjlOoVMBsybDvFN/KUkvg95Yw0jWV7AazcAUoLngESl+fVqTyjRLTR7dlEPOpEuENCX
1SA6fphODvFfemIEpC3ml/RiN78JFh8PXktalMpA2w2Vfyw0a+VZ5+XNRd52YDxOFOthnXdCIB0d
ZXk0ZgvQY2KQ5Ahvb4W4o3yGBy8MCI4ToR9HPVcXMdSt2Mj5hnn1hUqBdPXe79IWDh89G0djKHA3
7+5agOV+sHmWaryfNYbd0oCCFv2H1d8nydVrI+Mc8urKshxgHvGakpxld3KYwN+6BRUAZhV3n9Fa
crYrrIcPh+MNePkkUjX/xRB9VK17cCEUH+WDHKmz2lJVhOdtP3PBa5Bx3vRPKaiVqtWt3+riyHzQ
UdY2iDx6cx+jq9Ha6Z6bbi+jIT3yfsipQ6X9DatUnwlBxAN8O+1Eygvm95+QfDruGlm3QFRZ4BRx
JC+IKubU+UkQ0UJQPBeSQf0LzxpXqoDkUQ8V/uPY6XaAEQ+NmZ3cX3icL9ewxhm1pRDOQYlBRZ7r
esHlZQpRC1CLgfq7yYpIM9od1QfX3OpA5+SNnrm32fNkvlUbLMWP1AJfrwu8ziUMURxYqzuKsPWJ
v0i4Y9/AHt4mTbgxCJcsM6TswAZu5eCnNXgfEGcM8SmkgBrmhGUnjGBzOyRQDVIkgG6RvZiiUwNv
bnE5qYmHdM4sB27gZwEBo1syKs+a6vGS7RerU/AAy9hM+vFcAXuOf3o+zVT76tknJOJ2QJyGQDxu
gFd5Ihgdl/kNyLGfmV00itxp4FMH6sVEaNhsLjWI75srzakNAHuNMz1115B3ETyHXjUI9NDPAJiw
lWc2Ejz5KM0F/sZaBOzrdP4DyhHFUD9TdmuCk2yFZgZWt8SQnh4+fUfw9U4QPps1u9U8EyrqADkO
rOD37kVJr9NJXBa4W80KJs1p1Zf6n4CS8cgd01T8ZB8XlLv2lKVu6pgIS7dFBR6Ok7OWr+HI/8X7
aNrqvPeImolD40FGznRHsyhUVE5yCDkG8DGYELjdGQOpJ8lBtwx2dzt4VI1zjFAwcKmWZKVUv3cR
pmROt07McRFG4D+0CzkwaE0YQpStgPqnFHcji8ZkodLNhsSAYhA5tIp0bVeT/L9Wg3sbaTqqx/2J
kJNbY8YMop/h/soBQ1MW5hnthA/Dhc3xa90yXaaR8T/H/votmxQLR196TjFRg6FtWh7lIaKC1DmI
xGO2oPsjcgozUZrEiRnimeCAmS1pelCYmet1WUGbOQ1+vNfcwwQhm4NIbioDdIIS0OdTKrKW28yd
0gyqoQVeB8Hivs/PEXiFM7lKN0xUr89P6MTkdxUz2kxRs7MNJ+tSY6wRN2FxIb5XcXDrLPtCI3x1
OKwhN9B4FF5tVjxMrehyZOQMViexvNToSbk6Hm34ECJ0ZbwU4NKUvDdY/wE+FwcWKNsck5wuvgwV
5eDdjzEQVnAE3KEXkkhqnAoVL+JA05a4N2XkR77y7jd+sL+2s2Ku1zvljNNWr0mfAod8HmbQ6gBR
T7owlI/nWu03Q1iv+EfTi0rktJV+i43bvqiAOZvIurwowmc+YxylsvXyT6mrDZfyz/NGj+FbQ5Lz
Pq5rrhXrviW3Q2nC8O8vMZRvECeRpS0UJRz9OlgtSZFiSy4GWwTxGjmjgwraexYsxpdk4+jgnII3
03smIivM0dxhwk+atnLlUq2NXtcNwu/RSnF1K0R3lj9wZAZCfXqCbVzYRfRcqt9n+r7gNBj33J4a
iLCwKtnxT8pU08XuADpXyJG3xJPazGhZxrXoMG88bWfUIZyhcgjVQivfW8hvXJ8eJ3MgmI+CJxi+
hG7+gHBLvkYKxk2ohWJ/5x4wIf2W3uFImWz8iZqk4uttq336p+9AQuueZCwHVtBXz87fW404O9ir
+tjfr5sUBJfYW/PyJc7kEyzCmdKSxBag1Hvw94gk9YXYpReYsOJLrDoXvvU4gnaCKo3cXhNGSCXf
EnSxvcX8HQnaSwwxrV45zK5/6pAtXG7JhYJzRbnNsGVYWruT0f51LWd0M9K9edWub0Mo/sJWwNxJ
oRG626G6Kh4icGWURVVa4stp5zfZfh/E6b1q7fXNVHwBhuvTZlDyVMNsVr1/5lqm3XVPLALSs41Y
WgBRol71VHm/jqmF3yJPJe+2sCDvwAlnFv98MmtCdsVSJ9mDLsDzrhOyYYlcWEnxlzweXRaxqQ1A
xxfypEcgFAbfeLxPrwyzKN+8B5nUpQbYWbbrWGVN+ZWkJdIS/M/SwveYiANWPInCdYC4OOLI6KEx
gDx7ZhBobYL0P+PX+wFHfRUO0FxoC+fR/bPkn77PhUoDzUdei3EEg7Xy9LPGnCD43RRwgeFSdf66
gHsdFTUYMRVT1xkioU4mhGjh8teTgYVq8e4wnU6g3JZSFcbg9OM6GSN/SIwLfyWIIduT+JCj9Tyk
lQFu2Ft68lQBtqu+PwPrETvoqPT0WAiPlarMa5U0GDFNgUs0ipdH+DiqTlURV7IIbm2aG/IAjwS9
nqZluO5jjOUa8kyY4SHUnQ/DZ7VAIy1WJVK0eAENWPAeyr4vIE0pJmJdztbQKJW2SG3AfOE/UA2h
N1YzWuMjVlco9imgMDAI2BY2+aUOqhW2eoxRg/VYcszho/sosmx77wrjMlVCwjrAr86Uyl5ncVAR
LCTZUwAvEn71BT4NL821KFeT4gT1OIglvzEAd5Q7koWo8yotheQUHG1ea2iDBPMBv1PyvI25CUUU
pwYXRLDNuk1Rp3rNtfr9FWD/BO+Nr146MzdMUSW9HSAgiBoeOJ7p3RGitYmZTJ1pYQk5v12nDF79
J23PkIGy6iS8b7pp8i3DdZdeH+eZkLeFgc/+0+bQovwWXaPmWzpDdXlVzN489iWtyASJDJ3T13hC
8updDmikBF/y0B/HgfasVokv01Jszk7+9BIMI+G6oBRNP/s3L9GsxTUOqn2lTEUrtL+zXMc1+gkB
LjWlXDTWlD+76IjyXijCLenY0/le7kgRoKUMqSTz5TMAjHGbY845yAbNMOD87/mTklXESnJqtccj
CYKSHqztEm6A2V7RHEzqof51BOTawZMAxxeMFjRT+AVJloSQ81U+dMLJEvtB0ykxdXLBK+qeVAqz
con1yxgfl8mE61gfMStQ2VasA/41vhlhbymkmmptZWusyVOTKLI7E4o/URm7f+tAU83kaLDW2TaS
zuVxUxMhe0Ag3X1+fGuCdlW+JG5vX0jAKtjP+vPxhv72QkloqwCJBCCMNC/ZdlEyHJ2yYe0qDmjX
QuIj431sb5vGUouH6cTGpt5wpWkhjTocitGJlWsyLsV3aJd7J9TfiBR2MX9vVRYVsmPXs5f69bhF
1xrHBHlvwV9qZjU+33nqOjp6JNSyyyNbOR9IiV4HzrP0yFLrm+UdMIUT0DtDYGx0QYNSZpUXDz+n
uMN8wn2hH1+LzL8Tk/HF4VASRnqbtBz09M3ycol3JCprfPUreUv0QUAn7SkXN5lacKfYt9gi2w81
9Bb1e3xWM57sHQAgpYROziRX5LO+btbn1IjAUcEAE/Ng7rTaGzj1a0ffDChUzl7qkaPeUIuue/di
4uSNCOqPpaFgueBnFRVrJqMle3Kfakavm4PUCXwb/buj8yb6UPlYgO40E+iewa1LlAEGc7fBIVcA
YkNVng1T9IkHe+9iYc89DIzMzMSRTqTRpkUyN9g9Nko+LPR9Rg+rtBfA0vOoTaXHJnjPEiLNzYaZ
KipuYSSyJb95DgsKKxq0a0wIJJEcmm0yc5ws3CL8XfBud1IMoj+H72rl63VZTUfjF1e5xSiYw8MU
4udi0LAQTuXE524lzjf21JMAybXoR5xlJCmOFM4u35k6rRFWhwBw0l0VG/Kaj4YlOLqKsWCZcRJb
PXnRMMdBJxqiA2vCkzX/LwquoJENb/kclTDxXa8wNckeRBa8bf5cPHmbJYbSHuEpJLfTNH+/Vf57
sQp6c/En108UoZCwg/zWb0eRQdAFRlQiy6Cuep5Fwwo3f9rWDsd5rE0rhh5nM4XRn6WtdolvY+Ee
M4PImyel1PPamfsOTu0P9zWjEpWMzkBIT1bO5qrT3KLXTrAWNNuiXZh9IGLmB0SGj/IfVa/DTx/c
+A0JyBXEghYuS7X1va34n8wxZug38qLswStZIEm9nNhMlgaLhKmvw3dxiIavb8VGylRWF9QzY6nu
4PPYgjoqlzlArW9Teo2m76xuqFJ+53zJUcOBg5PWoXWhboeGJ7jL37lIXs/TryQf8ojN8OhZrzTU
TLO63N4eWFMOCNTafozm6NIjCuAq5fNSvbmnNEdBJ0AFekKeXft7snb05ckXWJ6dO2DAD4q0xGXT
UL84ttOdV4hOwfqVWDP9KPkTZNYPSEXdM9WFiLZdxxZfQL4Pak3OfCIDKUgVU2DlKMNQNnBgviJY
5Rk85Y1DnyXJUc+GPfxhzYh26WywkCUOB5+Dz790ZYNzcn1ozXm+skDazhXq1JWSboZxZ0BJZx4a
U6c/iENZoQovFvZsrChyPwReXiteg8rmOF/L3+2/n5SUcm0KDndDlKmgeRCh0waRZOxU5X7c6hdT
1eoXRTRoyxjhc5cJ9kWlZx7/lRBorNgocyN2GWE12H/J/bd6wrg3pfnVSAwCDkm9N53C2ua11OT7
T2ubKaLfc+703GTGkupgIwX6ckoTacpfxS1+ZfdJJLmDeChjQl7jHx2uRYEUwsUloymfD93hszhB
2luCvU0VKVY0Na5aoCYsLbAPjD9i/pt5LIYIAUDo5d8nPmbVZV9oBB8DaCIjwowLjbMNaz3QDoTj
S238hXgHChGt4dQoJDo3TCSH1Aj7kVIpOFEY/LHdNKHdbrX0d3YuxEy6qYbXvR4eIQ4ApsYTc6j+
rjHJ7hAELwAztEZ5WkUIMQlY5cWc55m4W0hdfHgVxzzvu8GAlIMpvwpfcidAVmrEvj3rylYUL7mC
0mO3lWYj1EY3M/B/fm6zsu2p+Om8oXw9MVwIST7/GCBoAdAxobsUqWML9nLgfgaytSn4OJLm/bHW
zAh1nhnJNgrXuE/T/wTNuC2vS5UPeC1X4ftqgfXomzTi+pSJwngBw7Kg4iI6CwH0oeYmkVy9gpwn
8ssP9YExE3ASAUKpimsrzW/ANy+mz/jToeaFIl0I4r9JBL0HILDFV1UBlyzozXwGyw7u6qdvbfs8
HZ9A7R1sJxXpcgNFp1bkYooR+xH1OYL7uvaZvnPGDrzHQdvjJypv9OAmKxmVrRq4qSOjVmD33bzk
jkr6QKgW/+UAYLqO0u+7u5hAOSRuW/CTqHYkRf0DDcMhPL/uoEVICBbnsDbc3O5I9xgcdrW0/WlX
xTapBAyl2LEib0E21bxWDtv4LIR+gVL/XTRbAbj0HIeLfZO3g8T4M1Ulpm+afnRCqeYEziA+WZTS
IVrSG0ELp9EIjDP+mjfMk2UAn3lDd3mKp/eGDdF1kWk4rm6siCdTvlU5oXJNcsoiuGd+56ZTDWFf
tyOCnnsZtHnWflUh9XxLSMfH3NdroPmgor0Ipf28txfqUTTeUbIqhw5JzmxKiYdteEsL0JYoK7sq
tbu56ABmIl97f+vBH3qcBd1gkM5pDxK7nQJTxKC7garx0bHgjfClo4VIlNPJYhP10NvKJRzJAIj/
s2Vsb4aGus8CN5ATvNRAfceE6+4XlxCELaIaZIN5Tv18lT5e7u4MGNCrt2jznAo8az9HV7Y2EsY5
RcZrrPQflWqjk00RvMPMOYxUqGYQZf01ZwfG/2q3fgVaEPeyjsX9mlv7AxMrLCRGDYOSXE6KA2dc
xv01M9oHLerc6XOgrQsLOE/38heGNiHICQFtutiV2FrmYV6AaiWa5uYG4Qy/htJmy5JOIvTz2GYU
YXvNAd+uiZcsvHfaLltYrpHhI0nwg/8qrqex8UMMMaUnnLuaHqxTbzCxiUVsEG2DG+FAjQZc86At
bfQNWL3GyUzLb13/kT9tgI8lHbH0rpqNiwm4XRF+U1zsrVm4I5zgyLzaBqsyQVoL4QDkZu98qavG
kcJOaYeW+bxtoVEBGJ7EiDMaQ3Azm3gY0HKFUJDRVKzjyMD+ldnMkogcHCc9RNZN0q9zJ3hUN+PH
VVnUGKsuSxtxg3yCDMYh9LrWlhQiU3H8JSDKfg5h520VwGjDqTNcMhav3XqXi2oixbvpj0XUfJcK
1pyk5NyFNbe958Ynf7uix7wiwawe4x9xBKC8FB8zjXWGiwhC4rxU6xoCtjgGKjj8LYlpwUhUJDZN
rNz/oUdHxXY87XOyZ7W52+o8jEuwaVwJP74alp384JwcORv8ctluCYDqf8dJ/W6f6EnMyu0o7J2Y
7DXOMVSc0BZtivhrljwXXSf6bdCfD03yzZdduFEnqfOucbnWH/5rDEM40R41Lov+uu2DdQdJbp7P
HB1wmFe5z/JHmIw04TSL9akL5UJtVTcMqRIVHSkW09B5CloASorN26l3t26CqdOHldRLU2/PK9jQ
xN4QSW0fCqW89gxAeBLpbXUiKTYQxzpJdCD67mfacmZvV6A6/1HVzLXvm05ocU5Q428p8W+o7aYP
wM+f6T6dqf/EzBXH3V2eaZ5B4pVQFJN5OTSIi1rbGsEetQIp+CR84OmKTjcXn61r3iyrEwMHogfR
i+mPdFI8rzj0TUV+cfOCBraDQ58jMxS4kbKj0vyTtujnoGkVcB7/h78P78z0cGJ6z/BfSlmdc1jq
RPGw/BoR1MjfcEwWHkAlyDxJ2rmIMhptp+FyY4WH/45v5pVAtN/vyQWX+UzHAV6ZbepjsZ8ddNeF
kmQlUIydtgZytRcCrC64z40KXiDp3lw5CQYAhfYCqCRvint/fkn3qf+L+stylHU0AqCAr08o+2yJ
YBMQ2ypZzDfMolMQAkZYDC2LBjSajMzbtTMe1b2oUPmShT7LyXR4ShQ+VYl9n0LXOjcNVwIMG19h
Eu9YFZRidWeMsjL7wC4PmiEMBawFEY6lCIuSG9h9WlwQyRMa/vSt1sht2pNTEF8gH9Wn6DErFFeN
8AYqVTjgzUCgzYjT4tfwDB3dzwvCucbFAO/gcXKruBqPWP+uKDxp3MjJmntEBkfARI3JiVuBmNcu
HRPj2APb2NlPT6Jqda7iN3vIf4Mnj5+vfCE5b6lRpXWigCX2wWslfCBIQKGW6enKALw8FxNld1tq
rzgq5LWAUjgHi4VpP9RvUBQma2AkFg0lRpYPEG47ra4B7yS0jL/48nPsml2A4FWgAuatbklw92MV
OeYRN3ntkiQ5zNoU2QWjqLMCZz2FyUoBsJ4+l+mV3Ml5Vq/1DThr2liCCCsnXJ995O7MRnGsMtQS
hlxPGOdI+sQo1RJMJPPzLc3Y8F/QOS6I0Xhp9TNSeWIqgBWPk1hF5lz1QYjvO+0VSsHo2Dd7C2jk
5MZawYMX09HZVEiMUeV3GUnljXIfu6rKQhDuO2y9aCejKURScZKyquZEBnWqCChlPYshW+IH7S0T
+ZycCuu5I5ExMiyk0vscDJoe4Z9rbHZTyHv9u95DTXOOMqCheHwwB9rYTLj86ugkW0XUEJ3LegD5
02dZ/tnZIwuhVRHkbHURmig2JM7WhRyTRF0mypNaGuUky59L9wMRog8FoLf1kToREUMUFmlMO71a
hk/JH51fIsB1lHhrdZQlCvUag1LSLh7jeFJwKcIG0KNZ1TQO1aAr107g879rIDZaGH0zpNH6Lr8u
R4scVfi9y0qyKJjzGiqBrtriOJxiiy6lAPHNqwLXYCx4ugJlreZDqBXEfr1fe3154/1UGvhL50co
5ihC/syyEiVdfgRdx7BGYKM8kHce860QE274yA53LeaZCndzgTFnK9zGIp9TioWLe7aBiyHhOJJ+
vQ5SkydmrPJfxjcF4vRqaflllPUZB3dVpxAQmN1ut74CV/uAodg5wcsTGgsosbb5JBkYnVQwDNof
HxxdPaVnIOzJp08c1V/3IaqAJwtPJUjh3hI7E1SVHTg+C41CJCcJ1jkSAW24xZH7D4bMfCrrhuYv
39fBxQ4C6r0oa+h1+3U75G3kh36bR5jAcs7Hjx7q3kGw7Y31t8APj0n+hqvUQBMGQBd8t0O7nmhP
47BvYbk1xjXwH0rHz6JshgyYGMP1BhqRnz0qb/rdvxLOk/xuM6sJj2cHFMCh7opAwOmF+EBMt39c
y5tYxkk2apo2imqFQW7qbnuoK9rUftxSNma4poHqzysqw3GT8JhzDGRPLu0xztHidy1Zy5DsQkeH
sWhey8CM03z4S4/B/S5l7x8W4lCUR+y2+XP9VeeQE+2Yd2pCs8LZ1DzuAiKCA8nnsvMd7eJlVvxI
SCev6WoCbFFqkH3+tjMZh0JhCCUdYqwgDtJ6oTxbeVrTiVThrc0E9EWgsxuHPFFPqybtH5Agn+vF
aWGYENyn2EX2yRJxSBEiT2ITEDx6jJUW3+t66T5UY2LK2fYSOef8Ukzj/V70O+4H54iS0HrxET1E
Egti2nmZgTT06xIjx7+W8B9LBd4/JPe2o3ieTZbXOmClwudMftDPbmjaIYM8hWrPh5/HaTA0/ovf
YcTCcOnML3wuWptapocKRz065PlWauoNmRdZxgLL+CSWmunypTav1ChCW5du5gC0a5W/WMB4on1H
rW+d+g+GaFXsvDNOvpbFMm/x72EzxbXTDF3M7uSfQ8FQHKcTsii4OI7MMSrl8Fv+KtNHgVv2EyqP
x5tdI/W0FX5+L9paMm5Hfe9p+r6SIHIoTT2TiZCELfVPyYltXimh3mfpgp6a8Cws8mYit0BdJV4l
nZFdtfMMfewbjiNhabrLTM4It693IxwT28mUyM5rmb05+nOe4Y8EwZ/CJwgffSmw14dZp2M60LTp
PRnlGh5T/sZPXdPRgn2iEI2ILHdk4V59usMi25tCuyU/iaNl8FoPzf2NhxR863Vi2uNuv9UeSNYG
9J5XFsj5cW4ix4rHGjp9LSNEJEOtAaIc3sOhdCOOyIeBl3Jae9oQJxsI5PActpQ+sTkaZ52GAF/v
a94fj2gbYb1UHGBr75yY3iPDCn8v/tPTEb95kLTIvuUxMQbFk9DkFMLooqrs5+H1HnmvEw85+eAp
u0YXlEu2kIGa4Eb1AqFimEShA7PCarNf5lMdKPQ6ncMGaomueozoJJMyUYRtebGt63QSpCwpaHtA
FtU/71ACeqsOvVd+XfO+AVpriOBuudlq7v4cduQ7PTAPOS/jH9slle510wVz29r9kv7JUH3aElZH
IANCKZ0XDjGfPBV2xVeSTfi/JJcXp7wsL5NOOkK8P0BdqInADxyvmwSGTM3GDwEGKm0eiB1o2UwP
xulsAG0xBQRagltQ2LlnbVtga3mGPCtUpvHahTXJio3y1Jf48SMyEQGUuHexOQIIozDtjh63+cDP
bUvjHq03OS/3KXEUl7FCs45x6Dzmu2HhvM0xOdlpae9vP/fgSctdktP46vtJNVd9L0uyApERla/Q
XH/EbQ5k5xO6R8gK92XZj0MoffTz9EOXoSHxewDtndkaTGlaHLKDKKQhpRw6AzYwdjuXJTlBSj/n
O6AEZIrAPzLWDvJ8ylB1e1xWiBoLIPA3lf4UqjpEtjUj4ogDX+tyN+Kunr7LsT6k3NZCUxf8TYV5
h/24X5/qtVV+ckR61n35iBNrvI2Xa4VfEaFoY32+4t7wGBEQqvetit8xywmtaDyPwfjkD/Hnod5a
VypI3O+jzuct4YOf1Iu19NALgOGKBQe9IdMeS1vB8RnCNYfaPHHbNv3afuAV05RnqCnGwGiZUgcU
CO+GCulBxUGZawJf7K9W5wa13N5064bBPSpGhqnqsXVAMg+ap3n2103gGL+exbE1rJFgb6TfFmit
vmA5UxUUFuLKPKcVkSmMbMPkoWphQPyr3jb4cF1wderEUTGgvOhTUVmlkDcv50EWHiMy3kdmJ/fd
vfc3fv7DgYLh2H57eNxb/nsnqQ8n9ldH+0K8Oa1WgyE53BG8TVHPfRJtLY4GGQAd3osHTGVg4ls+
DmxKdqS7wx2O2JoOxCEqOj87HrL/j5btgbItdsuz2I44nwjXb+dBwVzNZhjbHo3aMDfuSpJUgJSo
hm/GBiqcZe/dfLaYRuQNshZixcDuIVLv5tGVboUiq/6Tz+G3Ix5Rry9viap2QhCv0Wsk67XGK3jM
kU6Ysn8xs2LZk1CEHBjE+vFr5a57CRYzsQj6HSOnVDrp+22kcqE3kX89rpKMQLqThghjlIG7Nfg4
iuKgBBkz9t/ZeSmnt+h8ZQeLaGC9QzXN+rqANq3kv8YYw5TjdRAFLxynOLI+ra+YYTBaC76pgPuZ
DwdpJKqOUNtZfqQoEOky1XVrgDINsoTfTpg/GOXafekFvbwmVk1w6rOiVeee+B3nWS2W1FkxFwTx
vZmdIDbGBkeZamG3E3YTwGd7xvlQ0n2XkaL5cCQBVJ3d7mfBF9e50p/F5p4+n2kW6WRl56PHK1L/
dK+AwCUXv3X9SB6avlc6X8aq0YHJjdOKTqfmhxf7aM56NhjRdi9BKQif3rLoBgdcJ0sjg606Rbbe
mlMmXYvk242qe/9/Ldw7WN3lzSun3VMS0Nom42XEiq5zr6O5aFo4FVaV08CgajLlau4YXglzcnnK
ADAkSFVcSy9wYLeujKa2ktVam22QChSuHs82c5/0cLjkUujAvHnAiUgddiekEM9kVBf7UwTA/nUV
q71/WFCxMUOjlqGWs3tHTdXX5MraNsuwOrCCC0QUmWyfbo63vVSU4NsHijsiw19gNKvsL0Nb0y10
UVtBx6ngji7Po0RDovxzYBaZgDaPNjqVS+WSozFsFljRGFRnsMizMEFEH5COO0powXeYVRBvDEn5
1wgNpjLtykjQEtogfMNAPO+sJqCvEzFR/vIAZKSRZBeooT0VQUJ7glf40bTEo+IqNCpAMlzmf7Nf
agvOe3QK14Lokw0uFqypI3hh3N9nqLUSiSQ++yNJVvS7AiFKCBvAb6HQmQ87m85JnVOnWjlOd4J1
Dz76rYAskI6auJSKxIVFC48+jbcZ3C5gI/1fAucHG/ayihq9DeR1XPbf4vFqYgCGxqgeFAsl/2BF
GCEba6bK+sy7/ZQSvjeJdNHJllBoFNb3qQKDDAg6+KexoE/3ZYtGAaoT8xi2cs9LKQUUc1DDFpNs
JUjXjQ85b4WUSdPb5PBu+sv13fXqvIcZ1o9hG5PycRNPBPaHatym4/hgAKuQLeuFMmHzbBetuYZe
2Jn/VXVp8bKl1fjKfskkYl1fhg/dYVUTUFqFN8XY4Fa4dqptp97PRX++0inbaKgJgVEZddQknNHE
SpaL3EXTG5BT7c/C8kAMTiRISKpsaEqmSXjf8QMm+tlg6z3g4fqhrY3HHrzakEfpUwpO6Mrv9sA1
UFzBxNejf1WYuzSzsLQ9IeGujqiFgz1uNso64iqdb6SavBod+cTGBXf6wHwUDCazhc0skU4meZTu
AAVxxFARuUWiRma1GZ8KQwUjreHoAVZ0bibdVUDGshqPQx/ZHPtEOhKLu9XV7H5D58K2932fEfUC
jThn0WvXue6YsUs5uznxmt684y6yWSXC2+9kO2j14EybRRgulBLO4XoD+P1bP4lk6pwt8Ulhq7wZ
6ItrY6h29rIcyr5nYImZDB519rgcin2OVoz/vIZgYD8u5zYm5IdsM8yy3TXERFESuLmtvdj+IB/h
geQVB0K5TwDDray7uFsN7jtjHWYuu+Vd95PL5zYVtBXwt2z0CVSgkbGLP8kh1GnDLzUPoYAnIxt2
tkSrBebh8ijhvJa9/k0WBoJjOUpcmIVaqrVpSK2JJ2k6Ey3ksQ8U8Sq+5lgjd9aXuYh4KBadwqxp
PU79YI4QYuQ+juab2Qxl5cIvpNNxAuhuhBbLGCHFv+iFunLQRkSj6oIeuwHU+dHj93PE9Vek7Acq
6sA4tMu/3FY87dWwoSLeoaIknGr2m90QdVGKF+OIih9Ecoy8PKvFPVR0j3pgCy5+y3zV69Ezx5tH
/+CFZQKrFPMCJp4rLkDvqABznjnrqj8U2hwSDNhuiCKouPF2IfApsvcvir5FZe0lCZrwocZmUQ0X
Svufn3EeyHB7V8t3+QQFzXdG75hFQ3wLRFt5fcpiepWly/+3lvVbofuPUfxIhvr8dJGOXuT8rOkq
JsPYqP/91Hk623rdCC7xXA6XDPQJMF5T7ZIfPKVP5dlUE1rPdyPL1S3hr1+wGbI5q6diK9exxOWZ
RD+RNNqz/AyYf3jS7s4VS8WavnFs58FWH0LtPVg0tQelf6EZ/J/xhU0z3hGR7bhH57uR9FBVeJFO
sEDFfT8MgQmoUByOOMMAF8qda9OlkhK9NYiUFzf9QlqkYmYNXr/WoPzgFJwKRLyaW5CFaIcaNass
lwcb0eNKi1JjqdwgeSZXFCfqFFWqQ+A6P5rXzbNgUQAostN3hewaRcit6rhYcD47YJD4IkVTYzE7
krqdPltt/dmjwrq/XLijaflR4mWiy9du95jcoZHfVXkbs2DxokbPBVoYXN+VYKxdHUCThwok9xmG
VbLYhqzpZa3bOSLbTHG3X3uYXl8jIkECOYeh+G2wnmUNk8Ytohtlk9o9gv0PvkH4kSjFTPNRePQZ
MfpnpVuTBE4cpaS5E/8mrgvbzE2EPKAbPOSSIUowoaejp54Ppl5HNZGoD98oGD1xk+MMoPcj2j0h
A6SS8vDfFT33watxjdXMLtW4WL3HLU+H8NgPEmwRC7FA1z3r48WahhD25CQ7CLA1O1zttDGbjtsM
FjPwfILejRYdJnhF4wiB5/5ryjGLiGleBb931xSXbguYmA7AP3/hqyLQQzp95Qmkqr5lGR5bg2BM
syyBUlqF6RtZWvhU90JYdRiH53bXRKDgiFlH9iCWRXC+oTtr1HRatmTsuAhFZdokaGHPKQuBMETJ
DQwNBfDPZr+KX3yIOw7frv86Sh38pKOoLu7pYFcmWtSFCCV4Nw+W/I7Ug+0SRJsRDZLqLzCAg5ZV
e8YuaH/ULGfMsChbfHW//18GMwrD1NLx3/BMJ0AD9UHagB1z4bW9h/ONBcLBamsjRyVYxUB1AjBD
NoP6o3k8pxwNFiuWqnFPZ5EiTR+ePApj+UVZ+hRCbugu4sIBjEVPvCKpcUOK2uKj4sCH23F5zdZ1
Fvi+w/fDsM251gJqbjO+HOXq4ET7SFmeAhw6HvNnb1n5njALo48Ekq7FAYt+iA8DNhAFRyntLXYU
4R570EG0WAudE2r9zPtHY7Tlx0P30jTZ7ZvC8Kf0N8eyf72q4MCnDoI3kNQTzv59IU80cU/w2x2J
j+BeyWRjylPQ94VRS86ENHobYKgEj1GTjN+g9K9bY/RV+0b+WOQxvuQXE9UiKaTOKNU6gQkBqpjf
n+dKAMS7FMMi+HEG9VpZ06wi3y42zTbalWDgCPYsHs9n5ZkkSf8I16Qltlh3BmT6c9q+w5ZUNNDm
FgjTFoTVs1C0dPpcOURfNrQODqfX9D79yy8nrtbUL6u0kCamBsdkaQqSrhBBRq1kyMNBRlaL98Ew
UaE9+tNkS/RMRh/aYZm9Oj1aMIGhvuW45yjlDLSmbY+uQjvXLSfWmfWsk9KLRKA+Dn+a/wTdGRHM
NpefjX+3heCwCRfDSWBi20rgLsAwRIushTypaIdDx9zbj6h9WzPa1rJifkEpGJn7nOje0qFpwLO9
0z0ys4k+P+ZPZmiz5vvunhY1AixuWMxJJyabJorTvcXls4GK04JJvnZ+0Z68GN0NaIdGp5eZevie
RI97HIZlOimEGINxd0EvFG1hwLLsZ1+MGBtymKZsew0DFO1k1d5qL0Ft+QvpOwx1RTYG0h1BV8kt
nIwrQzWkASEgFh412L/Bff5+rLG8pdXBiDXGTf79AURSx9QIpmDI50hAU0s9DmmPpkeUCm68PcNa
KGsstd5AySlNh8r8qqJgCcj3DvxYWZOo/UeyyoX6V9DQqUuzd6ZcofU73XdP0rPx1pqpmFcj8AaK
qfCxphowTj0vo9EodoLmq32PAkC2Xc7UNr8PaDtvmfPPwdkyQ82JqWQnBC07E63IR/Kfo+V2oZqi
0oXCKLyfUA7K35Xe6uqj0bEkzLur+kFgUI7adV0Vwl9KwT1K3Q+OCZsGfqa2NLlqZ0A0uEN7ZaTc
PkVdPzfEPGJbnLdZNLbgXb5gTpTdvcs0/EYbzhzjeQ+c2aJXDaIsHY+Uza9Y/lotCoPTzrf84CaP
f0smq5Gbz8cCd6sNwG854ueb/JS+SMvbwWLIbTUQ0FjBaoBk1OGjl7/r/vM2Vnb/iUvaz5KjAVgk
apdmy++ebP3Aw7j0KpvKpnesiIS/wbwg48GnRnvm+mXq2jKpEif37BarAreF9Ob3KQF5iJTOD2xi
uBb0sEQHSFfqzEZotXsTX42TMpGRrui3uvQ6aSKckrB8fm3jkEupNarQNO8r70Z7ovwgTvmS1o3b
QRP0J4VmLxBpC3/dCRR4o0xZ06111IiBl7K2SSDfkKNczVAZiXWrJxbPiD+nRK4IzvI6ATnKwPZT
SP5nZDUSlxadaxxm1PeATziBLg7csrz8iDXsNhsvpTYrX1AD/cQiGH2/Nhr6dIkBaMGFAaICN8MQ
YtACniGp/oNSJrWyXYFOh4OR1u4Zcqviyt8SkVjFKOQhcF/2m9KDlAVSWTs27e5JPhkP8yaOm9LR
PGT9Pbd7K3Ce3bhUasR841BmfLWsiJxeDYmHTakyn8x4Gqk1qodD02D7m4ndMCE4j2cZ0Ka7Ve5d
N/BaAPh0ztkXbSCuLNcvWryJVD00JC1ocCYcmkt9e9caidn5G4P8wPlOOApGYtEgS/XwiZ2IdHCP
ZDQ1q3OGDHLAoBsfHgWu8D/Uw2e/ByAyBTc7YOMN+9tkLuwzGwx9REfxTx9rjoy22428mJ4bs78o
jWpSWhOc7/E7E2X4r5qmety9xfBYvo/Vm8XxriIwCG9AxaXiWb0i254Wvduijdl4zS4Ze+4m42Xw
eorod95MO5HwBZUbpY7QCgF4q2jiOSQtfOONKGon8ePOTZ0lxl98WXAEOQfnFI2qMsMaiU1kLQG6
RSOlVzYfS3ZiO+vCEVBFEpDf+LYbJw0Dr5SP2XszxhZM0lVdrxXKAoGj3qdqMh045sDR8r/wuERh
DY2me8OS5EDmPdJPEP6QqJ1ccF3kLWKTG8Oyd0FfeM18eEjH9frbCUfOAhlNB50zNBlnbM6CL3Bv
a06kwAgCMNSPfhHyiTdAR7QO+nrC/BKCjLjbIP+4GruNbkSgdodYyr0uZGfQzL1N24vTyyHa94JO
+CkLeMxyUQ70i2kUby6ODCj1DZQvFw4q6bENcndmTKQV/SYDqiUzYE++ZZdz3Ui6kaFoWVxk6hsI
j7+/Wyj5XG2NjiqxcKa2sBt8z/05F0dIzr+Ba3CMf4NhHF8I8Zr+jT28llASVhDt+wzvbstWQUQV
3v9QvdsWSAt5Uhm9Y+F1Rw7iX61P7LKUH2L5heFyR3/YJglvRIxblc/9OhyeYOMfQNpxy1nh1BEd
Qmh/0y4MedaLFuOpfo5N06Dlo+0fNgqVfKM2r6h8FKHt7SEfcD4GMWpkmF3KxXDY1vzIoCtorcBC
UL8Y7zRqs6q2s4pxkXI6kD6cRkg78puI2tofN3fPmqZYJJvsgbpT72dAwMjCYIjAKW7VrPqIBxh7
Nry1bIsnOm6FZUbOvjbz3gHJd1YJjml8Hvhfo2QZX4PYEiV5NZU9uUAx61DkrI/a1n957ed15M+u
awygz1+opdWni9RniJ708YOiGJsHDVVnGj+3lvPw1wCbAoBJlvWc+27qshaXY+o2QbKVyjW4BOVw
MrVkGC8nfQFXXswPJXVBEwekBVsPr+uQKsj00hJGReS25GWmyivCRxnH79/6SaEr49Z/upEyXB19
Ra/LdgVoUFbU5SpsO7ydwtEJhZ1y2QJDMtVxmuqHuGMEio03x0g/2lDASODEhKaLbrH8TRLdnjyV
cISjVNGG0N4JOje7dbVEs4HQ1sNHmg/NosiYNdK++tW5NnOI3HgWqmFz/zqesLdHHCqlhklLFOZj
lKoqINumN3Bn7xbAGLa6oIXMjuOuJW5JW1ouCz1TbOX4o+Y4rqknILB+3yWZzgTBp5Ma4mnVQAuX
Zt/Y4pSuQ4k7Y6nPXv1hrjpowDrWihwTUJ1WvSkVi1O181SHOY9oZm02fyEN2N58WtdKiYIMwQez
xmQ8q5IvswwC1Djh0PYZPVSZ3ksbLTfPhFqpmjP/kabtJvkxN14KxJO5mmkaTVjoOWR8tD72tVos
bgO1oRqIOOpb04x5jhx306feXUsTaq3iE/ERgYKp4p8Msw+SY3Nyyh7Q1pWT/usWadEBXkAelxCP
vOPi8CiwH4W4ZdSYMMukz9ooFGgTSIDbUF2cZHY7vel2uGg16yszuNDHoRF+2Eg0PKlxn0E/0QeL
O/xpF6dma1vHwyZELO0tpL73fDfPv/9J430YKEWieCZfOGRGFVD9EWNPeee+B4EVVHuAks7eg91A
11obZ4qwrqhJ6ER+nCCetHseYS9m1VTqd3goaTL8qAlUEhcnNNXW1qJcdChlTttdBV2P29Z95hd8
JNPRpgCKjx1tRhryLyUW9gEadRtFKzTUppNSmMo+QKro7C2JdF23KL9CF0Ix4iNv1y3HWOst4hfv
yzPpT+6Rovvkw8eT73YxiToEUjH5H+x4kbqiwDzJLa8bSExNNUP4LKviRkFbDNB5xCvvs3C+t7M3
dAriuddKhCucT5UHRrBgqu1+H+ZuKcHcCuMrsqU2c8fRJM0aZ39u04Rz1WH5znqMme/DtkOaX1E2
rjVFN2t0dg8/SKfQ354EdBuXtBKaFwz9ApV4R8NNR+InssLKxOUe1XTp8s9/Vf8om/pDMQffNnso
nxOishbEpjYnAP77MUvbvEG6SSf/bchZjYN26hnSlzspg97SlpKqYRxzRp+s2g6E7DdGofYfFDdn
9V1ocYVe0N/DOAlshNFJAz7v3aLBKRqimo1PMzqoKgauHd2YyP/J7s5QORtIfhI7zwP6G4KeLdQN
44fXfYYzfgYGyS0eyIjpL3uaw6gMZIcBsf3jnGjMAxDO2XLSTagQFBE8BhXeX8gZB1aV+izTdD4i
aRqBHiCeh7SY+/dtNh245YYFHpw7KrUgfekjbfDovhDO5bCLoHaQAhfpNxfjw46h5P5klTO6kgF3
b0cyEr3qLSqNllv1sWKR9stkwZRMo8Y5Hqfc8EYdsqOakwotChNoK58Y0nhP62bu3kXtg388xbQj
i/Ur9LKojBaCMJFYeHQ+G7+KwaS9yxP2Cv5l2yOACFTid4rBv1/JMXJF19edtSFo9fGqkzR+CvWc
I3joA/4epMFvM0v4pBDVt9mNUf5l+oo79g3EToGmQptWPolFpH9a77w6geTC1o6McHNu6+51iyTq
b8CMTwXGnJ+R5J5K3Izxs5hbWQ1b+h6q1j20QeKIUko9AOsQcBd8izf+2ChGB92fP3ErPx8ZxWIW
j1obh9wN3jr84y8kfyd2mMsOOKHh9VF0IYhybCC7QL7Y0DNkJ6wx8cdu78irSiye64TxyrIZYQEa
M/8Osg3TiPgmRGHbQ04evDDnjHGjCGH0AIdEozLGqjiKf+RuFOzr8sDj3l/6uvBFmr7VA1GNX42D
80v8qrVfCWVWxbgqcZw1M7eURXFqtPHmSInczZ+z4Zfj3zuKULx4Tkrn1dl8oTp21Gx5XXhMsOhJ
gT00xbj7csMoHl7ish03dLJPaJTA0If6qEHy70MUxe2nqnmdGklxTCAogGRypgBHb8A3e9Ke0sc4
eGinCWBGskf1WwfJwzla+9++xcvClrxBkRkjDC1eyPCQHKZWGlnEwrHiY4RudUptoOgxfcvDNFum
V3vK4xor2Cy2+lNG1Kqmuh+xzsYNF48QGrUNwGgECTPHs402D5wDZ+Fc8cQqdtkFiKv4qvF7He+H
wU+rCavRS3DxkvljyXA37Bthvig0Ykv3ZGGBZgruatId+gNO2WATXtdF3jPF8JOn9y+cFQKaoGUL
j+MJzF+i60b/1uCluFMXR/fkW0TLSl8E0XTjr9IQeGD4NfHXU4ZzNdsJWwGuKMfA/JIT0AeQTL74
mIUHpWUzPaF2kCnZ62LDspMa+xmA1moTwzthBvBEK50qrCkiFB1gJIes8neYLf9MAV/cdMyDMCBL
IPWPq7x5L0PwOsAD7+Lg5Nx4urcs8GbCXyJuwj69e85EqWqbNb7qsU2IVyAOhGuuteQZFlcBG8AY
HzI1+E09Wse+GuGhLOGxi/ta8NP8nKDgdnH4KNIoQAsdWArmXGsFi+lDUDVfyCOCpEAw3XJW1NR/
zoNccgT+I6cpl2mABEBp9vhGuyF0v4V4MSoVk5TM+RiXjMeRsv/ofQHzv7ucTxSX8s7sGLXknPx1
iXkc1Cwuuu9BNnAlK0ewRNNTb2ivWYALm2vuwHflicaZ1iYBuvc06AIOIAZWK4k6ntDfpAwdhKI2
byBXtEg8L5OfoHpAGR4IUEueLE6nYzx4qimgGDjLsMxz1+j8J5bGZTNfTNUwrZE1rRwtLncjLA+8
9vutVcP+I/2AzwnhT6lHWOJ4GShp24P93+HG46LTdGo/b/PCRcama7qjmF8ZTBoEcevqtk5+p9jR
3rXtwMGy5BRCjGSjxju0Bh6XcuqMWy7oMbTGWFK5OUEtloQgDp6mmeqh5iz8dU5mwaesCey1Vrp/
ZMbqjPKdIUcBN5ujOCxcVQZXyBic3XEnZOnFhvqS0CGIiKmBrWYFh5S/6Wz2NB8hKABBi7e6XsT0
EQ9g3O/7MkmmIahUhviZ9+Z7MA9G3zy/0megMCqgiSshl9Exs+OcVJVVfuP3jIyQHHh66lZfahi1
p+ot6HbjHAVbJ+rUrI0BE/yW4StzZ9dElldxwWSL978g8SNEdQag1eL2caJ6BLKCrHzodURn4gKg
FOjCRxrB6drWZsSPPPqhBfOglbcvF14rhAO4omwGua2+FZ6bWHbmm071DY2ERJWGQN/hGGdLvEoo
yZtKFAc03jIDJoqzAiJ0gE2fZB/ns2TaoajmRElxonYjXKHnMCQBPrqG0zsLGzWZYBW2kaEFyzRK
L3Xn9p9/4jLKOycMczh0Z/rj3I7iIo+PdTDJ2ys7RmyszrxzfN5kG+2WnIjR424Wj/kdvxqo/fNT
aA1zB00VIV9lTDmXcT9US3cRMcoNIkXNSE8jii3f4r9Emrvx6ihIfAW3mDay9lTul0nstvtSmE1K
swATmbvJT/Gysgpa2b273dF5KX93SOVc2LukjH8gkhiIH1ITMQe3vFLlK6n+/ElFZ0uHjnTZFEhQ
LnJxVayrK4XoTu9VsP/XtjxMsnWS53JSp5ATmq9vquaQWlYjepbfr7l9Cfn9Nvvdt8k93csMCWU5
+UPRhlZLXbEe3OXGvkXz0oOg8/LCtgbrkcBPA8lN/p05jQ2rzeWpPcofWSV0oIZ5v1WKbjMzCDDT
yzvaKR4t7M7BXhO3YVlldbfWFVSYUyuKbMinavyqK8ULw467+XhH39+HFdC2mCJTk8kR14w85uWz
JMPeoVY9UIUcvme4ieTCtKC1AQMdPVM9m/lVC28adBSyWYATcogedrUC/qzVs7o3ZCfG5yXg9/oQ
yHMeD8Q7qEOkGm1bdLLCWPYyeDhbLQwS12ZHf3xpkJvbCjxKq3oljgbcJv8PqPwIO2yOPT7qzFKw
82/xbXlkFErfogFdDlrW2ycKOdLwkP4m4Bt3dNAaWl+VhHWXFRPKRw/tuWqu1PoYn4OfCSoUqt1w
DhqZJSRsZn6yYF0djJD7F4mX96txxDVZLxILFCDATTwyWxG+eIJsdopuQ0RyYgsb4v3BeahuKQys
DDry93il/PUBirgBI+xR6x8c61Hd+DAwka+WlBP2xynS76A7LJXK7hLlArFoBNbARshbaYjmPD/A
DVpEQj7nDe/f1f/dHWBixLtTC0JOgoFmg3TEh3db48wCyZknioI8ZqvMqHMe5ue6uaSY70jBYLjC
+2QYfaqqY8/Qg7hW8J50EZgVYDrYdsJtzCCMkEEstsymd9XXgFY64PaTSLyzH+NuWvLAwTBGEGAa
bMUe+axK4PQN2uhbcze1aSyUsG9vtU8YlfXOGfB09u18u3TL3yqHFNy399xRszPYtU6w7ib/+NjV
N05V6SHA5zQrPEwCPrFwUH3qWT2iTYCQUIQmEciotQvUzmBqWdPPEu4ufNJ6cw+Yy4YB1HVAEjQt
spq3oToJfdWJurY44h6O3EMIJye3e2/Wdrb8eKroRv0ImRpUQ+VKDtBfXYShzSVpBLT5pMSd+WLy
zVw+VTOpKU7gR0jAoVbyH0/hfpoi6EjsG9fb+oPZ1fU/+gd/g9eyYgOhHqveeQYWyPlvUDYdo9Jx
+D7FtnKN2F4DPez/0fN+7zk2TJRzf8lFcvce3lQH3VxzuOfejoXxeADdaXrEf1rPzKljAmzXsKQM
dUxl1zUplAdzhSQYmFI282ou9a5Y8hCLJITzzaCjswFU/uksEDbdf3Byz7WO2+AAsXB49s88x0fD
+ELQ2+mdlMceOWwUT9m5RFdQCQy2egnBj2p9xs2B9SwsiDWBnKePWb4/8dFXB9C+6niNTkFJFhAh
e5MvC16d46id90Uppo5goHDbLKLBCVi6SXFXU40kuJqR8o+bNbJnIuJART0bo9TfYNe+xZW5cfcj
ZKjP/Grol5r3AXAVI4JOuR64kLnFPAqHjFd5yLQ5vxWIrNKLJVYsG2lKCRWWTCIyUt4aYyIxpFZS
uS5/TPc59lX2Ow/Ga/+3r2Dc63j3MIMyfCqqf9AlZGr0jbzvVAQrN64b10NS1j8OdG/jDDjNJwkh
9Cf5ZnO+pE/7Liqagdy69rrdVQPJMd9abeS71ZwUngwbfTMQse650xekW5OSPdP7ECuSWw4IleKk
IQbw0uopP+z3Ti/F1qoUYWNIEAI3ib5IDl441IDrJnue8uIwjT6TI7f9ib3vPB61++Phgw+6oj+F
zR293eVvd9ryO//+tKRC8qO9jYnkkwT8I5tpLjnImZZpll8BWg+renDVxCE0KP/U5UP5KRo00s4m
K2uvyr8mR9HYwhyw6JM3IvMkRWdZQ9LczWeaftPW118Kn0Ca6leiVkjKDt2k4fQcPbriHmvKKq6O
Vxvn4LlL6jFpQVgmv1e1qsFpBkMJAotYobAfVRWN/X64CkHqjUWRDz7IsSnrFqZfOSseWd2YkjIL
t7iadubx+ht67f3n72yL4jTJ47csqGaAqSvyZ/Fd0s7VpS4KJ/D3FzaJA29rmLoeDwYrS1HNo9qX
pDH7LdDaONxh/Hs5Oe3epbsswrqPPig1tsistSI6HbyyfsNyH9vjxqYSz/fCLCPWSr7J7Lvu1RZK
E+MvKF4OcSc41o4409jQIqp7oiLNVGv7eWZ8134NtMkyEQt14but7B5N/THbLvAiQNrrXLUIkHri
SGpG3PR9yt/59F1ACmGr++B4BVFrXojvnn7PVI4GgHVeTr/qXNGnsJpKA30cu5IFmRS3+0GULdt/
b8PTX11H/w+rSZ800NWxQQrC/UEQqP5kqs1oPbXVHJlag118WuyyjLSZGzt6bHLSeHUJF7G5yfo5
IcN/jvpCyI5VbmWPoI7Em02ps/NlLwkcNjt7uS0/jE3PJB45Qjdj9/0xOMpbelIANCoWaT25TdrK
nviTBKHKI1A5PPIZz7YIBlYFYAlQ6M3Xed4rCDg9+Tyz8YE7Bn+pRWX0gmv6mRft5ZI1cvdF837R
ZdYhzUXiiFc2rNkBEBImRIKNeoccYFGGWFKma6AG8bjLf7ATG4DJWwRua//70/whM72WlJAQEfdI
ROz+ldhf0Vqbssnyj31t0aQ/6sFlD/qgJLFvdFjhx1bTdUmBeU5R9pF25dbNpMW6Q/7ju5HdxdJR
JJXJaHccS8CBoIOzeGQAY0qXP6x1wx1QapMtsQNG2NvHCE3gJjRs0umBEoJocKrQHLSqEQvXCT+7
dNDyDxr7r2vidt1/JiUd2cWKQG6ggvIhHDPORCR2SfaDAnJH8dpv6zTp2iiDH2KU6p/e1TKPgEBD
mTzLKDj/o0VxKZGv9PTOBN1K4s787/z6X0kPiL/jtdZQMJ1ywAlKz3dAH2eHsTeqv7TlM0gQsJY3
5EF8LpLRuTl0+G1gZ5TbnrY3lWBErd3BYqXAw60mooM5ZLCn0gxygSXCNYMI7cNfW5q4AVK+llV3
nl7lE8rIAzbU76DqAxcCRhDMuxiTdP/gKmAopAFgjeCXSALamBfyl8Vk/THzMbE6MZh3zMjXvKr1
UW2GVAUqkYhY05Uc5e3mCAK4VySY4XjEUjDm5YHSiGHAHgZGc2d7qdjg2nvWC6gF1dC7N4v90pYs
i+QEalhzj8xhJjgQ53QWEHc7+f4Z8nPaB4uNvj9RmhfTPHKFYMnXxjWFV3Nhw2elnde3tSMD64Yw
AVID2VKAtrKjWQTTyj9O+4eDb3fkA0v+UQ2EfU+mjU+Wr379M98mHyFpPnY7H0zduiP1jYMX20Lj
k5plvcCtGfJU9jPbyf/pEasz4L4m6mwrJRBog5r4LzAcsPQEA0g0qNngK/bQlUhvMQ8Z8YxV7sE4
TYyZnMtdXFrETZvdvBSHMlKGH1GHhYPaaAqxacvjz9lj9tlq5a5hRAPKgsIvOdOsVQknqhkRhonm
qivb1Oo+unrtpZJw9JDhzbzhJRWcOQoty8N8CPRvBs17IlrL2MGGH4w6un9CKJZu0QzFjkhP9poU
X2IHznqgsOtAHhIsQmFZ2gNqo1qf4WRvzV1fPQR3wE6FXq0FWmN3gsDJ7ruJtKf/Dr3yyWmgahdW
VRZ08OaqAxBWCTWh8+c6CS/uRR+aSb3gbdXfi4EZsbAvueVvhajY06j9JoNOeb2/Mz90UGxZhFpt
9JVGuYXzh/ElZiMXoJu/XNmhBNgShvWxUq8P8OdjTMUeMphKupOB8Vy0Ll1A7wXlgzWYA/kUjcXZ
2naroNZL+8BdU+uG+SQuM+Ia++Fpb43WQbvAzVlauDFVM3E1kVgUOKwkuAAfvBo4Z8tAokNSt1c2
hCR48CW4Q0mIYWilnKWEUHxU03858gWpzhGKh3jz64nw+S3OSuN3ttjBxviaH2xeyWaeuyLtPIFN
pZfQ0yPAbITCZrESlM14KmehQ9lHJuJpWOWaxjo+1fzfumREZ4gUEMhBN3Z3WOgxROWAdjencIy+
lxV6lUnSiIMnY6hmmeayW9fIL9f04FtIDXB2Axxhv4bq7wGHUDergfgn0rSfobJ0JH9Tr155/Wy7
iE3dK314ADV95rpmGc907fYwbY5LQDjAIam7XTlLyMUjBep+qntWZ/qxrFtr1qwZ7JyYSZ8z5/2K
7HlwdGOvAzwNmhnCl3vj7pc2T5IzDQLwHrcWh548D9KtksiGo05kKb/TiICU5vfv3I3psn7cXOwn
5w8mDD4BywlGHHsotyU51puzP1TXy3stLKwU9Y9x1hPustTJx2qTuUCti+SPyw5jT6eUX6Wsu+Bo
Yl38Mfh1o+mgbbBeeeIAXrjTTPxAZQK4dRuTRMWqBDweOQHT78JK6P9Bjv89aghFkf0V1LoIhr7P
7pUDITBk6L1HOP9abWpPRb1D3kfFFqtU0bygGtanKRsyl/hyfgsvxRkXxwRzZ0Esfdm0aXihzK6Z
0sX/cFDEJg1yQYMqyvIO+Z8atHQDfOQi8YX1D45ectVHLFYF2pnvGP0uKbu9fQSf+6QShfASFX9o
Fgv1cISREPPzaauan9sBDErJw5wYGPrCr6XbvpxhIr2RjUJg5IuGC1V6P6g3bePpLvyswAKMYzp2
RktY7Wr+yyiU9L2277CGYZVcQLd1IfJ2uO3YYmFxakQfM/SUgIRsDKwlRLhkZwxoREVaBbfX1HFj
ZmFuc5y9u8Lngw9zjTOeOSrlBOTAPgvK9gnABKnEC5t1b12q1Ne8kOl002I/6yT95gUwm81m2qcf
oHTfJ/W2DLbY2sIHrg2sj6WzPiqskJmR8bZwDIv/FBtdGfaI5D/dveaX1ULn1Jkrkrc/sWsEAuTe
Gtiz8TIM2MsgPE97avLVp9NQ2AB9/V47ZAGgJIACOBwOOCXa+jO9t/McwYQEqArwVDXaJOPmj9ni
6sa7+ITLvsFm+KtcGLmiw2+zSc7125+b6736OFyd9hVmyY6+YObNj2wwiTeF0yFt9fQNRy7K5NYL
WOJZYB0jDsLFfkwxvymNYJKu2A7jVKzkY7WjcF2PBJp0UD3+KAOLl04m+XeoWMkYDeKdY+Vw9OrG
7CgAS/5GmHJHulrt5NgrgN0oGN1W7hH0GeJJTiNqn2vfGbEnLUFxAucxW9dINicEFpQjd3/Uh7/t
HE0PKMcWtPlTUSg4wayZYQmQ/ZPD8IEl+F8YY/uZuVWyx+aCCaPCK+9QJT1bbqv/AcrcugSuxYXj
k854v0xQNMgYxd2nOzc3WPGvAGTCsx2PzyNz6fugahFaDhNZtDSt5ttL/beBFUgsqMnJcX8CNjmp
79Lmf9/jvqDsrtucjjVFNdVkHgisVoa2zCphnGdOxaHAw293UbGY2fcwn4WW6xOCkb/DWQeprxpQ
5UE+s5+Eorz/GmlUGvYE2QqLOjgsXoVwz/0PvDBaxvyrdYGt9vJpV7YqlAOsqpKUzrnHU/eEfQV/
eEZ/b9z9w1SWJymFKtTBanguhfybgSdXd4sE86ff7Jq8sjfeWBfSmIazh5Mc6Fr7kefc6DJMOHWq
UbI0cEoapMI+tU9O4lQnDFa2i9ORRlUThN+xqnlYpsuSsF91AQHgfXkvZuCgsSKF/ITOBLt4Bi63
oreOFWEuB/U/QhsKEdjqgZOkZPbWLPf6EVvq+EquhjPoQoEMykYBcPVnaHn5RjSO0/o5gPu4OQbY
LZMvn7TXHTXBwYS0UuP6tNkC/VJ5KdjfYyle1GsPOLlncAGrVxxttkV+HyMFLSib4oC/aTBgkfkL
1ik9c0O4vijW9hqaqQI6ggVAVPn0pg3VC9osc8uiQ/kJk0Th4vf7vzycIx3qAv+mMyYX+krm8Cd0
41Xa9eIsnBlKRJfRnoGpqx3/MDpK84nuZESVPBnfu3Xz1wLZ0eKqtU+3Io08e5oXKd740ClNUdS/
Pk85JR4OellT6QFRVj6ydVT4zIlN5+lZZJjn7M3w8muZg2oMylj0DOb0SRtmvpmAd+8qLpKxWDbB
mMKSIDZJfNuciDBUTWIue2r9l34OYK0SuNhBS/OvPWLad4/4Rc8g1URalvxkDIUzgKcbF8ecVzFB
hCrLfpIGCx0ZOMRFPIwpRgT/orT5/HYckXpNzRrNYUI08lfms4rNXrfLLxWzFvaUJn4tQawfifNm
5BTtrAv3anEZdkU5Qwdb3R2l7ZhcpcpTlYulYvWIF0fSjhLj+cSMu9CLhVGg9n1DYDq5TeHsJWoA
tdUUTV1WwvYYK+RTuQyAduowR/IJetH4sEV5Jk8pnkSf6GnR6VkfcS1womJjVmRvjNXGJY6V+Zhl
b9/a05rzH/EL7tCtDRecs9xU/zkhV+oysxxAc22eqGifZ3WsEeYJUkJhTKRr1J8LPOJ8Y/wYy+cE
c8sSmQAhZKNQDL6X3cy6WPZfaVwSGcqi6mbtsvJYET7vvA1IU37A+ws9v5NRKMhfI96mN3YtCD7/
4b+0IYjvCQ2RC+28PXTbZvE5AgNV2y9YT6goT3+F+rxq6QiVtVO4HoIfmG7ceeRwv1EgN2qnq2fc
WfOteie/ffSz7ZwO5mMqiKpyCQu9gW/tQ92ko4D/J8e3D6U1D1Og4nXofHjj+4MiDg6l4q6Rhl/D
Dg7tFmgzplFgePJrx2+GAZGrbfWBUZsUQJQlhgu76sFdrpt4usXJyLtE5+YkY3In3m+zXjsXVCpZ
iddAuZqE+Ij0HhfdFdpiV66TVzHFfEHH39UA8P1kyGSzsz7gbBS3DQbjF89dajxlav3+ar4bnN9l
RuGfvCinfuoE48TJqHR+nMKfV7KM2WnDjMLcXO2A70CRvjGywRtRAb6fjYalHYKkbNPunDHVjpT0
TCTWbgMHGcLUMlEpu1kpb9c4jET3ofhMEqr8SsvV3WfNrUBOeFV+EABWVT7/VUMr8R+Mj/yRUjWF
jqslXwKKlW4DhJjatdY8aJMyp+D+hmaPxKEouR+62rRCle0rrEr7v54jNp6/AEWCqR4nPQgC6WAG
EtJiy6fihsUIiyZ34Z1rGiYuOIDAXjLuXr9XnfTWkHoKulsM41wR7Djnxj4OnjAjVPh1i2YBUISN
5/kOqM5qeTiXG4PmNJp3RJ+Oj7XntBRWuxKoo4c1MRmFfVhJM0hrBpWPiNZ1pHLISyKNaR8gduGH
UwIWykLolpGfYrjE5YLBC3E1m5q/uY1aniUNXZHJ8jH4Pr4P0fbstUca8KVhioY9Axq3sc/IJPFv
BG5Z2QqJ53kdN/vrmILKOixvbXjPdD/e9wY2C5hz+Sv51QLiF8/vVGvsBSdrKO43LahSaZ8esUzn
AsdwQ6CEiWpxU2yvjom7m6OxUtjUsi/0sicP6s9sWfeLoM6460ehMtNmsFngdNiXLahjKr5jAItY
4JH0tdvzfeDI2Oy8EBF37cLvl4nVsQupdB4xpzRU3ubhfXZZ1m6IsnN6rQQ+Wxm1AX7BuMoeK4MU
pNzVmQALSmjIJT4JBM2ll7lOg6jF7xxOYgDlDW3vJMcuzuW9qSwJ2+dCLmf1zM5O9+XRZ8bB9q5L
uJ6990xSi6N4PfHTx3O0sA4hlZyj88lGQjoPM2UuR60aYEjuhXncdIU86odm1n0lo3/JzwIwigMA
rb5IdfVDTaYEXJj702ikc2vKWNbS0KnWkx4TmcEYk7QxynJDmre8O6a13+KXSKIZK+eTB3rIKUqR
I2iRV7XtDuSyARoANKi/nEbUxa8+fvUNppX+OGRVrkxjbJ8SNh7ETpvfu+cyv83fh0FdzfmG4e7Q
UPmG2WR4uhPJntmDb8tyO0tcrB8S/Je01yCXt+JIKH0zIAcXg5KFCVcr8kt4Pkcwe+ldKOofIwFk
hfJdncVmQ6btRgk/u6VsbU+xMFmQYuVtrLE0EMWddk5I6Fw3ofvcX5t5TirT+lXCXOWU9LiAJW0l
3KgEqisK6ElBnn4QPm1+0SvgZYNA1mzhW0ipoB4R7vK43PJy2U0HSPBmoYIN7cOStdwqIuIg6f0O
v2pOFU5dfR5Jtt+4ry6CCL6F1veKIIrbWh06nsE9oxoJJOkaAW7G26DlUtnyGZ2hWj0pnm/bCsMP
sx4TrTpZrBxAL0r7sm+Z3UIDk+mx3WRCQjbfKGpo6OjIwH4L7kdjh8eoKZb5TGx2qhkofe3vq1lD
W4nxQmgZH13z9gMmsqbfH+wU5lVUrOrIR+oLlpD4k+K/khpkgEHquEoepYQ+5reHLZYrCvcbfA2f
CBChMI1vyMxld7PDfkDy4z9/SdT2BX5k3CLHYBGwrTOGyBbNHqIJbJxrW6y0rScc/WEs1sZZP/lX
LIQx8NQFBqeVGlr23j91b/ZZ5DYTu5m1oW7AdKxy+1UHc/JCmHAPrig9xdn94exTLJ/zVk0andzL
cffP+GwmG5/xcZfpNt5KvWLtDx8zFvVF5RrW0MHFeh0wKJQBVkKQspl2xtJ03HVtYARqWOIylazr
z3VVFbsYjrcRNsQkpSD8YH1i06kKeD+7/nNB7RMeoc9tDaY54g23I/V4Ocn56pMCgSqXWfEUUbHj
BI4PQndcO1ijkBDFa/wIjmJPPLjIGr3MwqCj271HKvYfie2j+w6HPJ2O4eKETD7w388HVhAG7o83
M/oqNvuSLe5KHB27olICLMHCEuiDgsUoWAjMyhVr/jJPmPjgcV22VkU9YNv2IaZWNniVxSkZ9VH0
dJYq1T137peU4Ad7Yxh2B2gRLbEJK7p5qc6Rc572wVtsH5VKCKxLpUoOVO2aXNL5uL+4CpSoiBkd
C3PvclW8FLpYls4N9m4kzexV68zzqnOt9AIQLAxd3EHKH8uo8jncg+IH10AeQmVehtBnpbj33zmb
bcQyoAiYxjH7ui1Xts/SOQ+m5i5V4SwuLAqBovtoQ32hvkrZcpJhdh1CuTh/7C4PVbE32FlqiGgg
ryRK/oMulvIxBNuL8PSisNbjzhQxYKJCpUZqExX/3/vZKMcLJ+p608EDJs3E+WOBEVBXX0v3W+5P
OIF+X+OBx3Zl1E22K8S32C3XWVMpZxslqySmCUxBf0h6MWIR5sLL76JWuARa9kTcdWEpjiO9CJ+W
J5xqDsB335jhBvw/qCsGt/Ty6BRPfniS6nxJ8KQH0LXvefehwWcxEESprJl0bNtygH2NcPuxvKzD
YEJe5LwyoeGaAVyfcdOOv+BYsy9x9w/k5Waqpn/osTHuWDbPPi1g+1o0ouJNVurpotNVHVVgl+0P
uZEIHvIjM0Td7oaIS4csS628leErDtT+sYVQ89c1t9pagZVAZeABvI4wKdwiD0wVj5sAehuHKadw
RIRVwBMCsFF9GIyP2VyRTtxz14zdmsfRtEkJxuXvcDu/O/00tESWwNjfiY9gWzmaHZqym9yTVo4u
vZdusBYSZbcXGzTRVZ6h/hwTXkJTvkhEhos9i6vefGj3uwMLXRfzA4kS7D1NRx6Jr8y/ORHxmoRJ
1gtCHxWdgGcKXXYGrriz51SN82Bn/TRew1/Sz5Ic/a8Z8myV/QjJ7JsV3trRQUiHY2gWqzjgqFwe
1UihwL4XoUOW4lkH6NlWxSRRMotJ7Kbx3qXe1u5/pyxkSoG9a6yBhfpzNV/b3hNp3pZqG9XCoWE6
R3H4nEPFXgcyAJRWyuHoOpY1ZZjS4cSSkBIwtrSUn314Cd3/ZU5tQI8spAol0WE5oqWwOYrF5OAn
HF6T6KmkXbZfpME5j1VG5o5mTvZrLRuJInbTnkw/oT6rOlxM9DGh8kQcp90mdUbLL+fR2WEommn/
0HgD/4QSFPAuMWtdViqgyiiIa7EIERCVhNnLtimUH8BXTyS/aLJWJqT04TMkCBVFbI3D4vjyBYWP
Sri1/Vfw0aIroxGXBYr8Z99F24UaUo6KLDdF58IE6WnJflsHh4DKVY0LiPUJWTjYQ8VYOD1t7WoB
y5MLn60ueEsRckV4r2FrvdLboQkf2DQ+r26r34C2UrdE4/72dEpZlKDF1C/CQbyvey4jERkI9a+J
JFS8nJhVr/errI3Lk80ucykprzdzEiMeIbfFUuisBfZ8iN2bkkjw2snHe9cnc+t1PoaKxmKrBV9Z
Rj8AI9Kq7nPQkvwFcaHcnfwpzVbS+CziCf6TP91M2lr0VBnpEb0hSLC7lX5S5T51niZV+P6ANWOs
veZi1fMsa37w4FPWNrW3sxrImNFelKdgqV5+hSm/TmJntWVTHJb16EEdB83p9PLw8QLhBQTEf2RJ
yAWORPyah4nigQPY7xDzd0DWnCIgURGcLiyrL6OdYGQs+mm7yyHhhpHEogfQ487J2s7VrBRQn9qW
P9PWIREVt3jpN+gtEwRlkCceB7YX8dWV36RH1cVnyCYDTNKHBS4ZCxKLgCFADLXvKcz5Jv+vsi5I
wHqYIq82lCPWFR3N9+CxcLz+wXfkfXJ7BdXW+K1iCqOKIeeOI6OSSG4TGTGpJpbzGB8uZu7Q0XQC
HlTbPtksVF7lqeWFg/9/DzZnV8spqjhgL2DhqkQszzUbRHGJiG8lnwopTPkUUUsnL3Bf9KchElSM
mJdZp/5ygYMURwuRLBImHvsVRawhm+NuQ77433R4gNIhfeAUndswd5YL9NqYBCuURrkwvK+jNb8S
cr8aICvtA1K5Y5wHU3fd/ie8eFR96IstU0q6KqZIyY5IganXWJ3x+ohjG7ud9AOvAHKSHImwYH/h
5oY1px98WfiVfWrv3HMatyCQqFk+mqBviMDDwcc3g7UCAkxAnrjxS2AN1tBbDMhhXZHtTFQVhfp1
RfaLq1yv2ylYBmA9FQAXkB10aPoUTsP8ZGASTnj+phEQB28YIiUhkYjOgMKBXTp/dia4yHqjCXi+
5BWdKGVKdZ3yPJu2MqhsffOvYCBtXYEtg+AUsYGDTwANZ5/ady1XlgHtwxhNnY83UgdUO/Fxeehq
o149ANwXl4ofOweVvE15mpceqlrAejaMJbiUQtCdd3mooY++tDoPdfPNotc42MLmsq4GbA69tuHZ
Oopar3HByl7ji87SPwCxY546EtJGjkboKSfIcizpMUcR1tGjud/cvrK6/0t65UzuNtfy7HuYj+Do
TbE0i9nU47F0ukVVi+dhTAudiLUtA1xq6xnxUyEqOrtkiN5orYUkKZKjjtu31y2ccIYsCwRpwqHC
sKeeD59J5PG7ChPv8EziDnSyYBOLKyqaa2SWaqM2GGS0owhF+C7h4fDcqYiyWkKgN7EQz5k4Y20u
eCsXzK6yNTXoTkw7SuaGZhHeq2O4kcOzR0qLNtuslFxTirnGwy4/aN9e7+p+Ap9EaJfcw83Iql1L
hlg+ys7r2dIm9dkmuS9k+P42TqcSQlrYdbsJbuqKYG+rvOnw8QGQA4gP05EgBAUChHKHVZnAn4fI
tFd3kDntmXKHkoE4QbuNZjp/UMzIPFZxq1EIQ3im0E0lOdFISXb8CO/T2Djk2Yv34xOhaocgFrFj
PwP4QZL6xCgitBnzB7L6yi5iG8S0zm6JNwU8Qt/ZAG27guNlO768n2eb/zGINZTvihLkUPQTBDlZ
03jUE7TNAHig8ZJApR4zT1U55VKVOEitz+lor+tMgIZNpbri7ageO0LhDkYz338SJKZi1h6Iji3t
J7fK33f+307U/fh/H5Hfs7sr6jhhwTR0YSGuyuOK2oES0MLnufK2NaOYwaTHI4MnfRe0aiBkQJf0
bRnrjNurZVVoEPps/UAliWq88CAeIc6KNjZK7oxnkRE5AvOEtIHnSEOtNv76k3EMyskpW2mRfy0C
KYkIbYYcACgP4GmJt0b5gcFG37hDKqKB3cT8SyVbxyc8C4wGV+GPpi/cOHt41PrDMHMzHnw30g+Y
WuEhGJZeVLJ9sWkFvsxQOFOOdBUDACw/asTbnOR4+IULHpqOxjmxshchAwO8dv4e0YW9FTdFPcpz
C7DxGwT3yUsBrQobPEMHAiFb7duOGKbzVaz3KLPSLEmRDzcZjbss+CN3LZyUpjkI5Vk/VTb9wemZ
QyxoICJ3dftEv8pZCCx9+5YCcO9vHpAln5ExSkQqpBVOXlIzeWQ2WTsvX3u+mFOInCOgNknfwlY7
KXUrW1b4wrbsVAUMx2v8pU7ecMSaop1ENhl/zCnXloeyYZwLdq1dxRRLMKSXnQYkLWtkta8hB5Pb
8Q3qhaw8VIlTRKdaoc80pB+OFbUXq+k8dXz6oo1N4B+Mu0bAFN7eK4muBfU+FPxFow1bjfp+Jhc0
pMY8jmR6ytfYMPpMWTkaG3epS7/ZUoMFr8fld6KwxmYzljAXmyMyu3EGZsM9dmwJT1BzRCW/ksII
gKsND07rZc4KKBVjdGRaFkNNa6e4bBfFSscHyr1PXMZmWbNz0lcOd/RJXdvaPE0ZpSLakNuvs3qr
lEUtM5rnAyv5ytUA2St1whfKoZPonHV/u4pQq0dU8YfdwFl295HW/5Zfi8T5Yqcrq34+pEsFdrNd
pASXWWkBUIreGdUHzv2zsr+Zy2487Q0/abeE4Nr8qLWT90M/SGd7tjiFOd+nZt/zbRPHZtSD+NR1
NqO/+skPFoWF5/7wqDGwZBOc1DuFF+x9zQx9k5VqeS/5SOJfa+lTBTmCE1OW48pH9avus+ipRJea
atYe3w4kI/hIHbCGBNcM7WZBKe+R1icMHJu4ujoCMXAoBeWeknJuPu+l3dI10q8Oa2W2GI/H9h0i
3VAbsGlYgNwJK1bIwUEeKDFC8eKVXt3a7YIkB3QhuCmIyawOSEYBOaHt3lw8HZpRMIJouO27Thdh
tynAlGSJTeCOobhJ5uGmHqyWiQgLm9KPfmgLHvm/1SxtkwTkZPdfXAg1Kvifknn8GNZXLpdI3Ndr
gf4G6yVx8dSSCvxZFVybVeCGH9YSOnt+Bf0GOPA7HLnzL4XJ6odcZP8/ycbEZefOjh+ABxl3I6wa
9LupMSGt2qJHtxcuBwjM/riQjFWrFJywXlGysnBTQlLxTjzEbSX/chDHHPI5q6YnfuUSS7mZbiA/
BSPcnPjOIKXgagpx3Jsh5fcyRh0yINyCAZiyXvSq40y04Qqx46Rs1ftI3eCl3qvgjFsipjJ0GKZU
kAGClkvz+xOaI8MEUYdUFRB6RzxYJ7vb3fUeVI57QXyoyotcz/Dv8OsibJzWnhyjv2nJ4RRZWJuL
zAaqAivil7DXsqOlYxDQTQOA9iGpOJQIlsK8VhTseGpucgG0bgTl7vz+zdemPF2kIcx34LYqOc11
19Vx/8/y2gQumQupTaKkCs5PrT2B2YeF3N0RPa0qo7JD2YnGwnEXm20jSsUndlHOJScVlNqGa4cz
FKL7q1S63FrfPB3YhZ+LIHwDotvF9HYM2S9/Qb0OtovrCAPnt3cliv7vfDmSi9g0Oe015wxWB/YC
7idpMLx0EHT55oPa7DfKQJYSD6m2u2Qln04CUPIrVUgJ9XKMQZ+7UH3JdxRjiXpOSNso9gEHeRrE
7440EZur/CleU0rVZp3JY+gsSWKGoSXUz+MWUjFXzp5iichOaFzFk3Sjw5svjHKkrvvTw7LhFCBb
AkoDiBnkqijUqv1gJaOTx2Z/hKRLhM2/lp4zl2SntxaIoN7mFAlwI21JNftTQUD8CYn4iQoCXnfQ
ZE9Ig4oWJuDusDoPWW0HKZGV+zm60wULaypkCuDwLecfN0dXEihsu6zDxaKDHGjwOtG3vgciFltt
4IBh4r3DKDJu23zuPHjY/xB/5A2iEQ3IWBeug9PHtPZlBePaE4ggUeeen43t/KVuL8XGm/o+DHIN
lpuRgIGb0gwO3cc1Wy3crOE/lUo1K1zOnG/kvnuSMFCbqJb6Si3eG1WM5CYQGSwLxroSYNGB+JLb
lcW8vx54XjsQQWHyP7awa2MQcQsfH4z3ig5oKAceGTv8PnZw8DEmhvw+wwglF/6ULiR9EZ8UvcMj
dlKKqOa5BSx+xV0jlZFS4Fkw19jz/9+b7GDfaSnwI3OWF2xe99TCgvjAjk6oK8fAdC/NuVBH0p/H
eisrQB98armg0YDq2NCmWRGrSsTC2h8m6aDNxCVI1X9KIhU4N9U8DMIcvfGKtzoNWZcngVCs3EFf
15yVZbggGMjLSLxUy4ntIeZDWuD9lu28yTN5T/7Uunel3kbb6P5o32tuA9t9FPQ2men5W2E9amLg
wtt/phwPPccGMASRBY+B/nhDsB6CyhELDboCP2/Zf06jvpvXmZYtNdV2sCNDn40sTiQmW+leyGai
HzYxCAMQ5uTCESHMBjz02NfFKAgQ35iMTPcAoOQ0q1r8ltTLLYYNb63jGX+wJPPfPiICifRewoyl
u6sQcxgPXfe2lx+Z2eAC5LTyA6XZPVi1FQzGsGEX0z4FLUplGjASUxHIf6Z3/bpWRO8xZME3wSjN
fOkgLHDcm+Uc723gpZjnwdYV16eMqtBNAL/J3UlREF8Cj2hJT6dV04aNayobzxZgA1H1otTP+Oqz
jTVUxjIRQfcFBf6WcRuvwchMlTuz+bv/5SfJzKuTTczzYt2/BcrDmwU/8EBOQZlYikxxFMcUWpcg
UHOBpQMna0fNocjrQzAu/RoPtapzEnQTT7tEB8rX62jFsLnnycw06wFkHJd5zhUx7DfgmHTbGRsA
nrWpvke9zir0iL+XDeEnIZKJHsO93r73Tq/JetVZZuCwdJuAE7O1bop9DDZzNItsOU3DQiRRaI3J
VLJph/hNCrWXLm9GEMnF5inzExN/TBR5mo+794I7Osspvvc2MKXzKhc3PkJxX3NFJIPFFLKvZLYq
FpTF/4DOF6ORHO5OyBzp1+9gR0Ux0EyND2J15/YsIN5KKV3mS4tNNbxy7ghOXS60erQ2SV1l89wC
NGIO+D0GhHGOsK8pvWeq7uMZLzUl1tC95SyvIjrfA5geh8i1I5rL68Hh1koIVaKX5/lU7D+3cZiP
q09gjczwZ7cDFyf7fE4wCKtds6sRlYu7rkapr+B8bD5W8j3mQXFO8IV0LA0521A4MRlvzacde4Sp
4/Cp88+4E3qrjsYal50rSL5hAzsOoLTGGCtDKACW6AfzbW45F0RJoxFMUeJ2Pr+viyfJ0zgT+ZQb
R0HFXbjyG8pSH1WKZjoXj3Zb8x+aKkBXFxa+tRUqyLojQZqZWxMtjm1nmcdfYTUZr9ksTm9M+coC
HfviUcW0F1Phk7YfvnIPM2uLzEVyHotGxiCZMjLdntjJR27IFKeCrfvNXTL9lsBZ28NlAUqPq2q/
5U6WkeSL/ZAMXaS9KBS0IphKlrHZ8kyG8NL5yBZ+3UjMbO1BT9/ARhd25CNLNA4nXjcqq7KiZn6I
+jdaLrF//5PCiHfA4nzoiCl12fBsq/4nlPvsNEbeVNrJnZbm+PdqdfcKsbz8XWTMECiCoT8UsS7Q
ywmzOudTtHC6Z0ia3qVAqlmXYuhA2f6aj/4YwRsYTVazVPw+EzIEfgZdFrHhRguNvgeTcE9v5zkM
II/7fiUYRiBIFk3aSEf0OIPxobZ4xtTLkmVL8do9pUkKERyltqBTCI9cGPRbbmj+5AZxl0Jq9Y9R
4wpKWMDSpWANtoECnXY1SXpMGCDDnBOYL6tRbr2lFxMNBH6FWIGhfLsqGeRA68Hb2EguhghxOEhI
x1ewIyCXg3URniZDzHWyJelM7Cjy+Ax4lIRnp77pwp5IuuvzOSIA7a3ej4HqkCCp+L9Mkj0nwS68
2p/f2Re+qq7ni1a74je/JrN0YKRnAfdXJgKq1Tvum1JSlNx+xPf5ZrNjvMQ3mFB9zhZ8hUj544Io
sxx2ULlDa38qpgRCLF5OMJiC7Wy39o1FkT91qqxTmoZkYVZvkc4JMjt/ZU/Nbir5pbH0aMLO6e2I
kRZ1ddPdYp8TWLWHASSLsVjzyaH/om+zZuzImC8gWJTeOXlE7KJy0OlH0TYK5LWqkMXiMLU2fYtq
Evt1dw0lFI7ZTrAzj7SZgOJSDAZ+Wc2d+idJY9uIRxA1yzO9PkXmPOE/xzJR6wquDacGxx7OAoS8
tk9i96yvM4+peKhdnmL8q/NQHVJZrAgJH806aX5ntCcbHK/DIk8yKVMksr1vElgJ2KHnbYk91pp7
mMLmttggQpPzt1yMzkQCcgcn4TTQ/+UZGs9eX1NT4edm37B+k+9CZ9Sz31ZH77uN0rsLZ2yS7RTE
nPElFxFY5J/FmfIQjyZdm51d3Xod4F6oBkTOLFu9vBu6Dh6hFFJXmYRoht1Ss2qlyx13p8aL01WU
OSxoycLVXiPQdx+K8YRhmG4XTnKc7eRP8Y7uHZ9NWw6qcUX/GfTy3Udtbgmg/rleKpyQyhZFoVpc
jZ08lj0V6QGbymPXk03C4drem+m36P7YKjP3m4YgPsyfZ2ozLiDSSRDsOHYaY4692pcRjdY54Fqv
sAOQwncdz73bUp5nhl0UgcY9d7JjhhUqFLeAGZzM9k/EDQC82ETCSDFAF2SOX7two04IwC13DTFV
srp3vmb9qDZgR7Id6JgJTcvcyTOrhxBGQj81cjP4dSt/RHHuuqeA6tzlKE9eXiSWR/bQWa7oQrE/
AMEmMtSQ+6Oo3WW14rimq+0G4Rg4HdTgT985Idm8nmXndISHgOLyudlyyPwZPtY8qXXwPSlXkblS
tcgsXU3lTxtc+lSmDSmatgeyW1DAnvpC6fJVRaZ/aP2zIJ33mk/jFDdfyu2R4FkmSuctYq3xS81v
F3LA3fbAgqDJ7zk8B+bWVbZtcput/VUDshd1CL3TyWlIf+bJrxzrGdp0WoDj/vonok7P17uU+sOR
hQ4TSYK/Fg5Y54Lwrc6uR6cf0X0k4jiI25tlsbI3v0sns5KssGquxXHy/9gwqWmDnapqfqJqiArt
NmKebGCCZ+PJKVmYTNfkOPkBQd5F/6Dg0q5QeQjs5jwNUXmg7+rCMmszWSoCBYwmnuld0oCMI0R1
MJvTvNr5zYH3jfepGg/ySzefQAlF7QGTCJ8XgIVPh2m/1vA0AtBkYgRq4OelWwqlS++Y3xC5JhDf
2P3s05IZeOORw8n7y2O6LQwtMXB5Izy2sPkQhSUirA7L2m3NX4yTLCI/uC7LNZUEC0xMMq0kmF+X
r1Y+iKlJ05SBIV4gctYEdZJasQYNaEM+LxJ/n7f1rCyRYWjGygHv48+JwahwZfu6U9FgWwhtfZiu
h1PYriWNanDJFPbgLNzJCIxoJmPSFEDZ2gR8nN5XwQW+mTgu47TLK5EekzfGGMXzqLz9jXm0hsAW
cVv+68sctIY+LeuracX/HAYw0i4ls4C1xwyahm3xPXpwGm30v/NDdigRDMjhC9BJIDUx0lGWVWyR
nfwELU/qjnYZjMTv8fpybZTKnnzhxwiewWREO+V2MYvrAjjsQZhOqTiwDwdOEHFUnis4X3D2Trp1
1SAnA3m4yB0hyFBjXWb6lni5f/lCS2+PKjSIVkFSvTwGFBYU5NrKCrB2j1aohOMZWwFO885DOnT0
11RWmUf4n079e9PMTDIe4y4z7+w7hKjXDymVISzj24qX5sqqGDrRzUrfi0eKUcP/WqpWQf1Vx0Bs
m6cJezBzvslQ7AcLQ8RB/eHXcltBbxgLzELmKwEDs9VYTaLSIOM6ylAkAOCTo/tYm1rw1Ha459C5
iRFWPpr/5nk3gNtoMzV2qkh5ToZz/5LFPK3UipNZWb6+g1FNX7GGIBfKaKl8uFAcRSbU4I9DSy29
iyDwwXEUtmbr5U2RyQUj5cX5aVTPFJJO/w1QwD1ueqY76C+/pXG+Bp8IUGGOzDEJVujDGMS102Op
TOVujyVxwDWTSLIIQ8wNB+tjCVE6fvl8KHZOudjA1fcS6oVJA2chftE1GLzviS08jfpWWCb9na/3
FB2sglHtzzds1Mfa2Vgy51vu11VuAWsNZuN9+mFP/QIaAX8VRGb709gQzVRDmO8BaKTRIw//1gON
vS5rszR7HfIzACnmfNG7/fd6D37WYTwtVmR/7jY//rk79QGwM+DvZ1uevODxqTGSX5ZUaxKmC26R
9WupKobsGhTD8JNfgW14vGi/5JV7etmXS3UqTLQhji7vUvJW5sGVCzx2q6Z2Jyq4ToDkzXapH9AL
cW2qfiwqpCqaCMNLuE6xBrey/C+8yKEqLKtexmc8H1pANd8yjDzawsg6Oe6KVUCaVM4w4bhix28X
8zUnNjwvTymnGUK+cYjlpUhQlxZYKriGFXSI94pnyds+eOA7pHyrJrNYp0fCBQ5A7484jvKahDVF
TrQ4VJPG0J7nRdweVn9XwVdmFcrWBdCLYeP27wMBVvg2CgkxI0VHTy3udbMe6jxJWgtmzOXO0ZH8
ZgyT0B4lgqBn4QzT6jJ3XTlvMW3CQvWUdGcuE3nVd6NNuTmXOeFDNFhYFIDxd1LN2Goa4jccAMei
k5hNFNLERJm4uf3GEmDHs2S/bSSzSetiU+lqrgAE/aEn8cIl+5q6uwzxTtuluMD0rledz9mHjylb
irGVGtGq8iiMfAfWpR/xVY6g5TVAYqM8/YM+r3BkdxxUMsseZBzBDmZUO1OhgHlgK3yBNuieI66A
0wOvY2o7RUXy/VqDeIchFXljl5QFTVs541wi8JL51hQB1VazZ63n53yT93fQ2YwWwvjOYq7cICng
TNfv6oNkeMUuqQ0DRS6R/S/JTCT3SqldJUJZErN9Y3GPgYntPU6AegoGzkAzkRwtXpdvZL4JqgQx
J4lt5XcsYtNvnvb1nfOseoSP1mFlr2AlvdeLAjaEqHBBT2QSIwZMCNQhNDX1WWhGeOIkbGocvET7
suDycQjXG+xmgogdSGU7ZyZDELeMZfV9y2Ro91N4CoLom5O2/AsIuNLPqJ6648s61jav6QFlNUNX
a2/OJ5AY9CUHHE4cMnrP+8TfsVLfP2hWTM7429lGKFuX3gZQNBN5P9rZt7hbyi8fCrxCSb8oWgnk
cqAJPi6QUHkEQ1f2JouD/jxYSdRYJ5xzyZvCO7AJZKRjffod9/mCLMXQsK9YE8yUuTfOrYSkkTKa
QBONXw0LtYnHZ4sjsisF1emd21hl9dNyKMtuRCZ6LkGrqhsZpJt+JuVDsisftu0ivSiMnZSOEWFl
dV7vzfBTtchdstHvLY8SLaucQeQZMgb/Y+FtrJY7JYlGhVeV51g/O18f7VMDSkqSEnhuxSd2btOD
LD5db35F17y+84hxo+mHMyJbUgxLXAYd7/y7cGhsFqy76Dhk20DatjEeg3wsXhbO2OSUoAMGNSm3
hEGHaCHdLa9ZJUFz+TOnK+dKB8gIM4GZEV1cC6/znn0s2H5l7Q5Ar8pAiyONIDY10/kmZuBVWUX5
Mt9tIXjzLQ/U52wpUDdalRtJs5TbeOYd7WDDue8g+z7XXY49e4+NL+xxOXfZ2GKRcsL/nIPOdYkB
bBgEPLuMAwSynqDhUixT8vVY0A9aBvIoQHllkhqBOWgstNCJMNXzAypQP45VaQZn6Zt7oClduGeU
nLbVIHvz9tvllZ13UtZqaL5YliwQRixcrqrXYvKVyBCURYFqATp7VaVJr6Hj7F7Sx2xqj8DMJqAK
AqTHntDT40tmFX+pre3nssEHwob/9zrK2MVYcki3m84oWNwu9mjwbmATrBQux5vzuUl5DJvKpdFQ
Qw/6K3b8vimemTyNAHBQivPKmD7Xkpn56bBY1dSltS/yhnZdiTTHPlWaslZgWmnJL6ciQhJrexqz
+z+XtThWYfagxkEZLwyd79GVx3r0q8MOucKBRMuuwu2XGGPw5oVlcKZMEkv3IGgFZRw/3BV+uZjQ
GIX5phq5BaeOxiCiK8FhPR3oifeZOACsCQg0luSGowCx+I2Xg8ZDqHnhuL7SOW0MdFU9yj1Oe/6C
0b/ub1jKvvfbgmI1OonjDBQsQutkObPbDL/BPmK7WA32jKT6lmtyxHBrCQuzUDCqWB9L5gc++2wJ
AU/2/z50wZ83Abihsvr0dVUTpKJNpc2NK1wicJho3x80Su4oOyPlE0zThzYfidNtQ52fxi1GypIM
d7Qi0oAacvLWQ1q0q9GDSVgywGgbKI1j2Y/VHWYGJd6yL+aqeIPQLnj4lsC33rpnKQeq+JLJ5SjK
TdWfsfafEVQDjmWkg3NTDIXhjdh/1Oe2R+vO1EiU9ACrXtHgiGtB0EhK1x1VNzmdYledw18uEiRV
bFb7ygwRtzhSWIxgcTUPsuG1XHDWPcCLVHUBbqV+ebOaJSXnK85RWT6OY842pEaM+GovVUpNd0Ll
egZN5zM/tjbDrb0iwrmN9lfAY8ZIoQTeFKiYWy/nal6L14TgtQoOeEgjrzSmSMKRTbvimOMFR8l4
rlIlZCsHhP7as6QmbEuBg+zPYmRgdjbjF3Dt5ek+aS+41pbQXbVyktE52K0rWsXbLhK7FUrJg/63
O+3scEyS3qWPtpwmsBXuXSI8Hel0kGFckG7sDcWzDH5Holc5eD9uNzXPCIpSRWcZuOJVM4+kpDHp
pOGoxVpXnnvm4/LMlZ/OoaXT4V6jPvyoZcik1l83ShxrPiulBT2LVW9GK0ElBZ3EJpFUZfZRXPxC
G1iR0nTQe6hpp0cVyjkPOG+kCkpTt0C1RNE96NJPvW30sGXf5MrEZTo4AptHpITEHXJRNLrd6Slf
cqjLXc9bNLYeSDI+dUks8d8B8/pMOH5ejF2CcDQVqIDUlhZFb+Yq0m2eAfdPW2kcrmYK2wXEGBqe
jh0DQtwB8A0tPS6Z7vZ/8HlERQVzlHlptS5Bw0fzCaxFhYb/kBLiioZPWuWkXb7SvWivtjUSpeyJ
Ggs59uBs1Bg5aVeGVkBx4HzW6M2ZA1a0n9yvT/nVa4vb+fFF5mK0tIsHoTpzwtsKT/UybPJwLJbe
xiLuBoOFAhl2YVZ1mTOEdjKAv05PjP9TqiU5xThSCH5gcWuLC6ukcvU5Rq0cnVn9NOqBstTezBZ0
8SVk0VZr4WQlxzOvvjpsOsp6xJ4J8RRNUFc1nmstXMIgi2n/SA56thsaSls1xd4SKAUnJ3xtmByQ
T8W8omP4tIjTi6e0CsDSCtNKDE7Mn5tiwXw0udRE3xUf2u4fulW9hXfrK7lZC8gvMPlSmAnJdVYm
Vv+OJ7D2B2TeDWOqEz9M7CtFtBrp9jfEntQ4pupzOolWjyLGnCXNWR8Lf//FiRFasc0DToBu5pDo
Za8R3rkGRUB6kG4I0VOXCv0fB2+JTsHvVKzHE/ieT31SILhhWgzcPqJLyqypRaAv/R7LKG410i7u
Zh0bUwBHBmD72zw3f7c+ArRBiJ0jX0TnDaPgI5C4V9I5ZgGM4lIptvc8+sTajDGNpFM+48ap3lYE
Zlt9fLG/1ZJiSUhb7snk3CIfqjcAagz3jhYlbe1FkZA/usOc3rJbwt39x+H0ZEaR6IaliFha1YDa
q2S/upFfsDoTUwkB1vBPlELhWbXETmVdCVJbtQo69dcw/AZdr1Qnoe37J0lpBkuuivR9HtrpWvLB
ObkRe/diiJoJPjMuKAPH2/mvdOslmlVFelJ1aJirNPrLPFyJiXLn4+2G5Jfb0lZ5cwWyjpb2toQr
gNylAIPaqDMgGkEvBIbJm0rEixRW3GAnTMQ3o97PcyUTPEXkRgYuY43/hP9bMkvP3vGKM61XPmQV
D7Xl7vUhjutWJ1Ce6Q6qc+3NROCr5WNmsvYSKFEoC2yqdcKbUPMw0lkSSY1gBuzMDx5F+8Z3sQqo
75HIcuyZRFK7RKnKNlEccozQVQTeO6ql8e/0hOVA+wB3qeBaHsW7IvQ5YUepmlN3s206VL9Ldf2D
vS4RcrMA4uLbp3BzEP917QOnW2eeo8JZY/fBcj8UybC7p4KQnpYhUOLia6TfbQWRC/VS2nKaKg4h
ZQL3Cdx1wxBn4ppMPx8pRYm/EDjsEK9Bu/2IYEgFnNwWWGjGoa2WXlliOM9Sem3ARxkDIJQSFXN1
Tb2JEIzqG07crOQcEpZwHKfm/IvriTNXObwoclSquoE4Q+rT/Z4i8007EHVFJkXQ171Hf7TC/iGV
UR7JQzcsFz1qGAXcvXnTEOof4R7GnR+aE3LZ1eXj6pJMlhGgAscZa1HolrfpjXN8IyUpCDSwrgC/
nAoHWF5JXoHq3ap3/PHjuu/4hLfzBCAW5vptvxRgsKDCxNcvXbtLYFuLkTlqzMOZcC24uaDDI6US
vbU1GNvVwocPneC5nCffIKEJkAP1SLHiEHrVc6OyGojlp3JUEm/2EQx7PbNGZAlH6HCSc8ytLgqQ
xnbhqEQ/k05LqdImXVpytFfsQy0yxsCpYxOjlXWZixuPJ0PfKDMgHrITDA43CF/GO8nuzuHCKQ+5
PIRckOXIEvbuKrwRHZ5gzfjq2i0zL47puVjFKiCK09Hd+tPMPmAd9dNl7VMoHAZZKRX9PzLDConJ
74PEwnOg8h4ErDG+GkOBSVVo2SfgipYIUiX1Mixp4aWR9vlNo6xuws6q2HuKh9cW9bPrtxOiGqwU
zogiuW7c+zNwV3HTCnWnAw7aCxcWdALeIngtfzDBubyk33ktcmqRnwjhtmM1164m9ubXSxcbZC/i
HjU1LONgwzFv4BQKKuuUgzW0TXb6Dc+p/HBCA8y0qHa1rpgpa0QGx9FyjD2xHWGdwz/PXKOEScJy
udbG4r/VRAxcP76XAs38cGbgpYCOOdP+SzvwqXX/yzbS78VSrWaEqOgh0zLtocO2WkiuDwdlEBJD
oCYd25GuM4Kd5rdk/FFjqq9iGyB/LMj8oJ7QbEPnimEzhLa/RDRVlMDZRwNqdbZWfwtcDyzCabFo
GuTec/mQZQpnLg5T6uTe5JrDykbWF7EXLvIL8Y+4nqvW66SXn1vEg+WvSr61/tB0Gm6DuDk/KdPp
RPcp3uU9MCsHsPi3FAoLFt7lMHccOgOoVo2XKEyZJfc3GN3WlrdCACkQ4NrU1ebGyDeVdc/htg4i
a/JROl2LViWI+bRw92ZHq7tGtzjd7LvrzTk36R+K/d9xoTgq1jSr9yY1j/YVDitLR67UYblNiWa6
wvjN5AtLkSj561v0DXGFoqWsBlWirrkS8JW/O3xny7PyDacI0FgKF4lbWRBmXLik+j0u3MHM+Hve
Wc6abohtKBlAl5Cp5vWjtCuwKlLeBil3IPGByZznHUnFiID1J5v65rkb9kQ94+ZetU28+oEh78y/
oYIcRhDm9MlxumBvTqduFm/rjEm1VUaUIz5ojM8WomP5P/1C18frh0xDyxkNKqL5eCVnjv/cDVJF
a9SHjcGXQVoJShdKAEyGrlk2noK0zjJQ7cC0t5z71ngzj3PU3ky+KRsIsmeaaviSaP+7hITowjv9
wIijQvPrtH33AOuzXUWrsVT8GmBK1xnpFRkJx1GS5SNcetEO8m5Ke03W87HerfuOHDrcwzuFkQsE
/ThlSLyW97h/ipYGoozKL0wQWrQXb3vHOxXOjSO8cJAL4K6pXvdaBpcDIERnfeTzOBfLvxgSYm9f
kioHHyKV2Dunkg4jRUKTQSJmNRROT1+o4LmEc1+j6SmYj/q8QDXFhkZKw/GkuhLEHI2uln91HbQc
cphpdKM/S2/A4LvH3l0Yre+nig7bm5Mz3Egzu1bP8P7WH1QK+Cxk4p4wmmgUpJahUdRvfQkqLFe7
RJvNCpT5CdcfijWyNSFuO9SPer0quECaw9wvExW6492dxR0lB+ux8L2K6MasLQZ5/jn83g7TJwKx
zNK7fgLSF/q0J03Mb94rtAjGWsWJCYtc3bBaQE73Gu27lEiRpg2/BF02ki0f+K8KYwmbnyDTXlDB
oUQVSNwSFgSimiajrWDH4v1zDI5AsX1AluDuSnAqNEqo4iJN/b4ZeinjyK9fYhPqpbp/XYFzme36
vCNyaJAOrsy8l/QcruSRvFKITyjJDpsL83U60k511QJWlxLuM2ZT7Y4TMXQPFyJBVvQQwvL51L0f
SKqrrAuV+t65NssSypT/zvI9/SxbJhXq+sq/5vPeV/lSihffSgM07j9YycrnYQ5SC9GacbFIVvzN
TrmpLaq+nizUkM8yI0V+cHlb1egqxM32xchWIiXqNXvcH0zTU7ftsqeWHYmUft82ZrbiKx55IAv7
gtn1EXQlbMyZGDEf+SEHqoVnQX6LB2WEuH6FUhc7tOoNyveYdNXg/1HaQCw3XM7Vnl7xTw34r5TS
xfmVUOv7bYo65yKhCQYs5CAcVMQLLpur/mkS5JblVnKWbwgyPr+dQd7amEg3Srf3bI3dY8zqPiue
dV/fscVoR1PUGePDJpPwLEUZ5CEm3q7XUkKhcU0tDrPbX1/VC1W6nnO9qWqE48Uv5IxknIy1+h7/
SPcDeebX0Gs0smbSO1yDFeaVcer13LwWZridIi1bQtTfuzMekcBioiabk+Fib+MRCfylFZytaSOX
FLfqddwPvV2cMi/qeKZg094EFHlm+frNLcCljgTPU91uG9HQYJQ2LOqYysnJzWjd2fC+G0Mbzsbi
mP9ax6G/MVAgq8GHStxy7cdKGIy29NAObWncwsrv4o76FoNc1/F8Wh4/u8rWGCh96cBA611mGwUp
lW2FW0yOU/cJKHE26kk3UgufpMQZ9izonL9m2EA6nV9a+89Ovd5MLTni5pLJL2WZXTAUFgPeeDNQ
y0hmnmBUjDWcSprsDmBnoVGASScZ8pbpXFNGsYKDdViycyPtamieET30oYONmDpAxMFkYOWVjmO6
JBVkLZRYc4HgKO5r/WuLQOaHU4lIDYS5aV7NI9QdCCweMZlCp5PV4t/adD96xT2vSuR3/SwKbdN0
kQeRua5U+9+rwqJ4MuKAxrgNRhQbu6jF3n0mmgQWNuSaWQTbG+mCRcRkHmQbRKuyj9jSv8fWq+x9
+OIb6BidNJG4Zt7pbsKHT6vA+FB/z5TrwFjmIryxe13yrgyomIaKpA8o5K47NjMVFycClPwwRNKR
3aazrtnj7v91SjcI5bspurmLf7cFud+Kqr/bOgul/Byd3NVJnh32dofJJ6pK5i7sSBK7mamXbV/J
8DKhA7f8QX2Qbtahfby0cafXxQzhCkTWl4qT/TRO7ovpcqez6BvQrcRYHQ9A/IHahORKXWOItu2N
bsQQ1dFCd9/eRWVY1UvnCw320lGM1IcdkJ9/JPO/ti4XfRnoH0pW1eIiNoFnCoUh+GVs3cZK2Ayn
ZCRE73wH8DlY0z0LRDdqqAv8Cx1QuScVMfcs2MqUlH6kDNcHcfGTMKlmGT036bQvCYvdizyeFK/s
D0LHkseMrA2kj2HNxF0Jpx1mA6WcwdSuHFU8FHHRkAn+uBl2MmzbVIpssPmMlrPCE7RQdkjw52l8
trc/AKj+AHZeFjI5ZOzlBP6YDZFht4vVamZfBs6eG3GKXcZT1NdKwgsp7bcixuKlV4kc1l1nK5V2
7R44T0+I/+Tr6H1BjKO5TUN34Io7gNV+sZUF/+SZgXwL/bVynUbvrpmbKBkF2pm22xSuVrAdEVIv
zJlgXoLpCJe5GOWvNaLFXggCozwTP6xa+xL0ymEtKXSZbwWvFdfeeCT5GRqcKjtdx3lhq+BueOS4
gHqXeqmc5kTvVxzZB+w/bT8hEBSiPAN2TCxvDMdvrdWynfSC4tkgZrBKneAIrzk54BPMQMa1kw6f
x5DlP5OjX73OC4SYI2N+sMDA18/n8zHySW17ybGYXj6cyyPjD9hIuT/D6WJ7gg4Y7D5zhzXf4zxT
BZ35pMTISkM3P/IUzfGfueh77ojNEnTq5rUaM8ziIM7pP93+yof8zG7Z4RJbbnYZycOyPqAixFFd
nYCYRQB0TYeUrZiEOfJdjUd+K6kss3vl60jhEpr9f0a30gdUZRebjw0+eIuT4BLzKe2cL+fYYPHs
ncowXJHNoXuGxG3x5NxSJrBPvYVhI3yPW3UCbdp2v54I0hZXCXr/dMIWuvMUqJ7v9K/G1ctovoZj
N2D+TpQTpjRLxQ9a4niiQp4GgseIN/v0KxbVRV8cqysRV1EototeDl3a58Ig8K6xvUtx0dIH/Wyl
Jas3dynkrwOeuWDbS+d3stvgfl0vUZO+7giFTZsvowqCYL6fu6lyDbdOwlmwLBzrPQwZg1OHHuit
MuTpUQ3t9AMNQ0Q8FyntoMk0sKry2Z9W2xsmWXz+g0Yqmt7Yl4Rc5unwxDdpPKKvGAHv4YdcPaVS
uJRssIEBlVKCXnUsryfbtVYXer4dhYKEuLV52f4mIuCxJoYt0vXvsecu1TbX1SJf56SihFgAcAnw
m8ZCCvLlg+pKJQ0u9V1n+Jd0FfJCm0nsm8o3L8gWvPE9ZH35YWXtQ06fFXUkRDTmVrj5u+3nY04L
A5uRSElrnexAzutzOnW0zDhQJ6u+M15tlfGzPKJgQYhpibmtbH2ForNYk0KEREivqzvdB1RenmbQ
gnyj84M9GKeqKB2phkNxhYr/PK7dLM3HEp1QYjRJ6tNqPFIejd8vAP3TOBXRYH/6rxfMYb+0ziId
hpZJUFUUSnx0zOQcmncStwEUGSAVZlznDe4nqgdxe7meRzjBFauvBPVF6RhDR1VQaq6X8HJ+tRVN
qOz8/G0u1Zk+3FvCDxfrQaXHac46W+i+zwuiRfQa71otzzubt1oKVA7JmQIf9QymCW+YtGJSmBnW
5DffYFWAEsLqZgu0n4s6143ybrFKlh/UoclQGYMJOb/4Lo/LbZ/2SAoaxP0NHaVp5HKNvzv++XPG
VUUv996ceXrfFzgV1pOWNUbwFDFg957S0MncJ9r6KKECdyaOC3tL3Qrpm3JDO415foS7Uwc7A7Q7
UzocRP4Z0BVeLVH7MhJc7QkHvIfj5D1/VCJmoDXwRhO+rtleZUB+cnQOIehWAVNMazDUFbg7Ptcu
r4ChHcE7Tx7YVRvaaNZDjAjJNhJMxIouZBF5GGTfrloJQAk6hpzU8bkpXZj/qUiTExoUE/ieP3MM
DgsLgAZ/CKSlLxLdoy2MzYXS2XZDCsPONthAAfWHc9HFbd+lgJQQNHzEhLCAsv2HWAN2kGJjAmvs
rJFHfkBKboVoHh0EkxrXQw3W7XfhTvy3tXOqlDi0cuEfFyYiXFbCdnCCgPljy4Q7GV0v1rWa8OU5
UWEtxU64hyqOWL3iy989NjZyGU8Z3aKoGnp+gmw4TilliCRgCX9PrROBu/R/Ei7U/8XKu61tivFa
+AbhfaEanHU5n2PGkhSsNgamyzffH7xQt5X1qe2jXg988zOwGNTJq2TDACstnOv/wZMAGCfvMYjc
E6CISAUK7yvYsPblPReOesv1uC8R01LGEoGWXIQYzhvZIL10qNQU+fVyltMCvccG2Arz9LifTvKq
Y2io+a0nOHwgxT6n/mGdoxeF8Vb8IiAGvl9n4s+264woQ4mDIfx2AfrmT4yZmqVlEI1cPJR3kDL7
ej6Ee/8xmRHvKazWZn5eGiJvicsGWDF4SYifUxfnBdBOx5ghjmzZYJLv9xT8bvWVBiyoPaxsHP08
IOxN/CYHrcsjwYuhJ901EUTQUApTpgL4aLC/4/id9zyEsMdA8elpRxkuZN9eb1r4Yo/47P80apxA
m8KLmEWwPCfdcrGvYRJ7N4tio6TSaD4i+YI8xOA0D6CwFwsXjVXYcS34xUp6a59wBFCp0shtZpS8
wwYkmxVDc++RjHord2VhKzE7H7pp2JGfmYSzhWcCnDycHlv7g+iDC70CDSUJlQv60RALc1FMNbAc
+slJidiJwvLtAGHLMlGMwkBB9iJxs7lNje/hUlRKQUCLabmFGt608HpLEupUpY52BTmPZdy9EuCH
ZZmhjLnJipSxNk8aGhMcMI9aBMqHXLGdpHXMO7hab7LsJDV5euMWcD/TVfjhC9CLDuTkul6lDijL
rYIOb0ZJantq6gXKxvKiwz2HM2bTMmFJGypJ6STvPnDTTxOpKAXDw9BInwtauPyS/cCimpWicVxB
lOmqSYP2T626QmLNuMf/zwG182omC/flbhSSfaDgwvUhLT7iYsk9a/UWkb+yNGVQsRTdE1lZp4Uh
YuF++oMJRh/6Lj/fqizQXwepHoHNM0l4nIlkXhKuExaWIPl7iEO6UVL4IFjd9PP1ORJIfP2w1b0Q
kGOKTJoHWCGdi6WpKUTYBDx86C5Ehbfx7hrAavLXDbcjvUgysNMI/goW0jiFbPuAqx5FMjsJarx6
3mGpKV+FnjTkvdBr9r7l+x+4Y/qY4JpS06bm0am2DAxQtDDhXW0dAQ1lLGvgFXDAQDkq+3/WFHMI
PksToVER20U3XixfXtztC4UoTIJpo79P9wlwBY6AzKWhcGMU1JHKdab5z0VZwMqSiWDbJ0Gi6dhV
8z2rO91uYAdxyFO8pYxEGuHZwqP2YMUUiOYOwxNCQtW6kHMqTOen5l5VWQSKL3q+l+mKuM8WZyGj
6Ih0k1GyftmDvojzMhWccaMxgkqgUg1nFaK4y282oSV7fJOZBU0gkmdCokr0U+XJOYoIVI9jrEhB
f6FrtdnjARwbWQ/WrDvvz0vYpXnr/6bDjyqxbPDrFmiV0+E9izgPe+O6zmMr7MdKYt1TogOE6Kuk
8Ew6ozrozJFxdDyAtjtHhIYIQtBoOd1eQzFw8+NHArHh7E33PaO7/sL3vMQ6GhZThzNyBi3VZjAs
l4wygKFclT68vtEAXfPCnVCdPo8eRekQB8tnx7zd6/nZQX33He8bahd2NnoRz56cz5XjXSbruJoB
5073jRafmGcy4aoeZuAkkCB4eEw4V31uDMeBjWyy/09b6I1+kzrJdEmTJWAxc3xAJCG6iT1Tu1SP
niLsAKNiq/2r/ZC+dk/ctSoQbb8tIWfiEL6zJNGm3llvvqj+k9D1JB+8l+EdgVYkHKlsImC+FWSz
JUdSvrKLUJ63vSjlQ7gRDJwFcxv2ciSa5JK/jw8yt+4DSLWc5A/Geog3H59drQpPU+9e6bTT6aE1
xgzOh/VDucXfeFQ3/1h/v3Tx6awFhEcZk/+5Ix5qtEwm1ECPNXc/mYWSEVejEb8QlCKPRKRqZKWz
GfobS78593HQd3LTGSrmaAWjPuUhNuKVCatLqsflY6zJws5/9uXIZ7actGewBQOHlE7zpToNqcih
fTJMqFSPrUdB3kFT8PktG4B6PU+zO8Ltyo62jhwGzaVEwSScKzL1xQl7m0RHTGEwe0d6+meX6syD
gKgshd7yhOifdMEtiIfNHkJGiA70KkgjOR4p57/LjiVI+2KhkRpjlJBnRIBiJrynww5o9rcfS+WY
q1a80fQW0CmZcgkZxkYLD8mvXDeynPTCDMFAmeA2bAz9/dIaEoXDKDPKAgdZZt0TKtwFwbygh5LO
jsVgqBftj7SoINNnRjfRveY95mI2PHHIPBlKqo40nJl5IgVVrPh1TUChOeYAtzTHzV358IcfHTQ/
4AZz+4wucpp+SgN2uWPoDuTkJL/gw0BvpflsKeeJGR5q5d3wAJ1jA5cxu5vVfrLDC9i2wTwG57Ni
/FL6eEsME4jJjlzQzrfydk5K1o4EhXVciH1988SmH5RpZwY6PXUAVCNUKUNBHtsiphLdOMqddtjI
tfh+Bf4bTcdzSpjlmsUhpsdyHXNd/UF6+zp+/umYl6m4KiA7Uv1wFNUlCwwXNVeZ67HeYZSZcgDo
ovoCdbW4NNoBnw4TcJ6RzEoW9qOfoXs/Pq4RP5YTBOTmf27HTSo1zvChAEZPj+evbxit1WJ2NxXn
nw7CtBmTdSYsgAZAxCzi8n/Su1qAC1l/tSp6tNzggjsBjdjM1Dbf0bC8Taew/b0MblH4oLJxD9Wk
HjXpwQDhYEHT6uvLN50dTYYqoLsxkf8YGz2PjHXgFi9jQKaCNFC5P73a3TeW//9tV0e2PP85RYIr
I36YY9+T3XXMrmUE5g9WiEWmokhk0Ugy+ghpZqwDGxvuXU5+MO49mshQdwLKgIyEgR58g2nyswUy
vV/AbKXEPYELgHaRnAShoKcdwd7k7RZhKBZMRV9TMQgiL7VbzW1mFTLrJ8SdPW3t3/5quj/a31uT
3irq69z9M2kSaiov03WwYBoR/HOH0HPzpc7l5al1ctFfoKxcnBp7s90Jy+FAF9YsFM3RyPh982ce
YbikihlmduJjvusu4922+0DusEa+KSXIt5wV/5N5+L8PaCVTWvti3xfXiFnl10FWFiqKQMzVbo1p
5pe0VSRLLbJ6lAw80LkCq4StDqdl5gEF/kykvPEm8+0NRgJ8Z5pugbPTK4V9+DO4DzLCNcTGjzjy
b8j5TzHvC7w4dYnJZi4HFw1CMGRAxbn8RqdreVthqZaW6tOM79MSIsDKj7oeDiFq6LVFnJMtIYHK
yQe9m2lq+oGyv+P6Ctwa9yqRrrWEs6bj5R4HI5D7h1qcZAcG3MsAZ97SNy23mREcRLK7/2kQRXTy
1Cu+US7t5SNsUZoZTIhIVMQ/w3JgIF6keMDH5vsxkNAcCLJx7q4QoXWHBPAQJ5tX8Dtx4Y9upOmj
88/kdBxZ/7VJhHYKHezZSaWuhzVKJZAPgK+QGcMsl691Cpkl8bDtxSOfVF5gFu0D7n1Jno2THsdC
0E96gzMu8ZUa+3bza/QRyyuZeAVydEnUK0e/FF6yClwfAixmMiP/r/PrzjWcb90LLJ5I+jMRqWcB
q2MW2C+qcyXFv2/+C0Df5XPAdQxyGTH+k173PV+RrpO1vGOz9YtLxV7dJm7someLSxCb6mpGBj91
TBPXpnHOsWpCX4z6161twnFJj01Tvr/SQ3+3tJers3/VVcG9v4IW3J1xd2SZizB9MQA0nr1yNErV
qVYbj/d4/K8T6/vGGl18hUIJHPzLd7N+c8TnznjfKt2PIj2/vqGJdAZLi5OVznpAuXVpbP8I7XDb
2wGD7RfEd5zFlo9vr8XxP1PxncDIcAc08AxoOPmB91HZcjiQt8WKcZs3mSyjpD/uaRm/YJnh3bYy
JyW8Bm7Sa4tCGjldTOw/fHkbuMGKkOy3OHtw9/00QnjaRggmhHhhFzUnyfrGBdWym/2TVrgpUzAm
qR5U8R9oG0GwmSp63eo293Vv7b7fq2Fd5QffNkwjhYOtgdsdTrZ7ssFgpLiO6Gxw8RCR1WhcM60R
x0Jqjc+9qH2uGymDxboi6OkIXIvcKGxKG8r53C11C6iuYn49VUy7IKe9Y0/wOueK91HwWelcFFOz
jXy5zjS3WyXyJEncaI7bmn9OVLBWp0kDQEIAswpFkeu84rw/XTq5a1TsU6+I6ZzvAMifHtg//Etk
fXcA7YjLKD5yjCH8t4yHAaHAmByLl1qHUsts9+BZrM+J/VSMMl+nImLZb0kC15XB2jCmfhnHF3p6
gWWBSc62y3+UMGSWhprqaIGn1HJJluqvjO60muH0uZmGLJnEI5ORtnRp/xeS9/fad0wkNSgD6qHt
tdjJL+UKRf5lZvx5YDLU0AEJJjCEINudBYorhR0TQD+pMyEWQukUAzuPVJE+GOSPOo2nAALvDfcz
buU6oXcYZf7GVfqFEylNoPKUQ8F5foLxpF3kKquFF8lsGRaq/26Fa3lTWcLpKXmOvki4Xl93mZh7
ZO+kOE5O7fW8uihf6Izq2q5ohNBz3lRRIPFkFSIJVRnRgc5QJ72NThAP7nGIM2404FcRs8OVF7WN
VVCHkUb34DdSNygbEAcTX/NpRCuDbymbfD7OACjqS3AyOwk6qDcYB6y3U/xYl2scTEWUK3kdILC1
UPsQ0u7KOUDWfqGX5kd0/BqUk4GtHeRly2o9SU2hiL1VlbxNzs6DLRGHRn+EnKYa98fVSCpJd1c0
dpqVU1sSumP4Yn7/R6O7AbAK6TdYTzIfEhPNzHQapVpWHxyHn9RsRdYs8sInukXx1BgsGHy+NPOl
jloovsjkSuVCmcG845mhVG0mkLuKGWhOZjRwo6peh5kzwvydCqA/sd0XMq7fET8T+iCMUdn3sHro
k2ZulR5WoPbjp/oVB/7r3ZawT45OmV7FI0TdwFaMo3S/wMagvY7qI5KATZD/sAQ4qKVKBfHpEq4Q
Ckx4dMKn+/D5Y5RM6LJ2iA4U7WnQwj5waE/qshLbQlwRjlXnJha3sdRA4xHWtLBBNho9pfHaPegm
n6mIo/OX4512HlvK0Xeea7BRBVT/9E1v74G9b8R5IF0IODel6gmit+MKGZD/0fQK6ufuh7kxlITo
oNSp4JuzzeK2dWlXJxy/1dGZP1SXB/+8NgPX0IldlKq/PIZQT+XJj9ijHHxeEBQTSWnXhWcgiO4m
XDXgxEdgqwd4AQdOIS7dqiyM/r+5WXjg1Z2Bflmx30Xgk9N3+7c9v6R2N5kzigw8nj1LUkbxfzwg
w5z9jkd92DeGhoPY7xVw1zCXkx09kwPOY7BR2hF8EAlDfvHl2iyFsVBYWP3X42yL/AoD1eQbKSCQ
eBJ7fEiuoNc1Paxd1HfL2oRIlF9akr7+1CUmSAXxtQS4/UfLyWB5w98Q2VYlX6pO7x+IgFictzuH
Y6GDyTPb7NKlcZjhk1WvfPYHhjDNSiWh8ngmRfJxV3uKva2IOdEBPEyJHWtftm4go6wfo5uJgiRy
QBv+p3IdVOTLnKHFlqHvriskv7SpyDRyrmGoD6g1PyJvt83jVSomQ8KoCJ46uF3g8EIR+8g62bCL
yqYQJOf/t9Snci1vmW+yqr+grDl58TyxaCrtPDUdVSo2WBMC7Uy36dgaBCGyGKW0G6yQSAwx7RrE
rQ6tEfa9RmeXbgbE3TqvfYlGvQqxmhCmZabSN0AN5jFafwCIy4m0pu+u1InsZPgTmbxFTpOzEppi
iTjAOuQAyEtpkAXQEKv5fxjku4GFEuY8HLYL9s66f8xuMpUlTLMgXRj8voB/uAL2UgUztdweQ9xF
B0wuKrDqBZLlcVd1VtYID34wWkF/vb0MW+TH0XFjmlvUHx3GAVMHPE9PQAYY+aYKtw9iMhbIjHvp
99Xpv3Kp6iA/3ZfJGBZBPIcFUjfcWF2ILt8GqTfryhRZIzaYxb/3ZC7HZ5exKmuIL9F+L+GT4Kcw
3o9FBKXjuWpOxGhC/sxyBMTz56Cxe1U3ONeMD7OCklZpcuO1Oa6dDgBgfmN3tViUwOjjkuYdAUv6
Nv0ymWbD1UvfmTuqFenxkkcZxNchCj/gR6QEG2UCZiPY10i6Dg8j4qBCQreIa3E2GuYfU+yLgeYc
KIvPE15bKPtNUyCfz4k+Tzgs8pWhShdy10nSTAqIkPuqj0dgjt/fNY+Ar9dmAa+JGb2kZplZTGfw
fq1wT0lKVAnZ4iPXGEATFd/qytV0AESfdahFk5Az0Y8ko3l9IF4d0FEYc8Nu1uwiKMPHyAmVymSs
bahcYszg74dPypx82jJB8GD9zA/WBYK19AwI5SsPBjUJkso5FjBVIOth3tjVOevSxxj+Yxa5qn8T
woymBbkn2BnR+OGtBa0g3rZlSbDgKPG9oAZFVBr+PBTRaQs4o2dxo0zuJ2D9eJuX/a8W9A+kfBsT
lddtSeQcRqXD92G19H1Oqbd2bpQ3EDvvxy1O7rkGJCoK+CsDSWdj/M/3tAm5X8QLhUTFDIgYRWZu
vfGaH5m31YDvZUIr4z55a83fv1mm6VpD5qmlgmIrqGCG17xDl4XZ4iw1Eyd6Fm1DlUXkYsBU689+
Kd89rRr2Y9V5DzlNhffvMoAs6QpKbNQmJKWbfnCx5seV6U1lyPMu5z6JAlSN9IEp6oO7jJafHlvr
mk18SQ/Z/fp/i+/kv69gs0kaSnD/frLLNFUJIArgsNLeSr5ESSF5+QDYFfLdXeJZQyvIielBDkS0
UhP8tLziVloJ+xPWtwoLW8mgwY09qzAixzQ2DMGZAwbQlUtEBQzTqzYLpNBTWGogjV2h7o3i+SUG
j0Fpzk0B+tZNKgKZYK0x3S8T+0Ea5NTwYoY5zN9VEODsa96uOHMAChCfL0/jWhrcfH/aW/sJl+B/
WHE1x+pUJvUKAfv03Thu9u7QCi8ILw2kHsAp7aD5wU52dthm+eiUBM9eyRE0WmaXOxBpEhspYU71
Bq8NNfkNcPYIbOq6PyMnU0wjB3zxv4sqWmg5WxCO+C3yAgxqNaJ0zat4xJV+k5vYE9UvBtI1Q66Y
52o6i47eFp+ppQ4zAWl7MnOdObluIDw/WFZdy/DFv0qfNmm+qrjXDIgftETcw37oeDFgL1X8YSLY
Rfwi2bYIE99TCbrAvYe/jQAsFY2AFAxBrlPAQ/vv3SSFwiZ1FnRZtWBNw6c0xpSvjta21/uB+GnJ
pfi/+QHWyCCnb9PnizTAMclSB9MIAkxrlIZS5TIPRZGnjpCxtUKmmCQOknAetbBlK24S4dR+EjK6
VJDPN8QnOGhHHnzzgcdNQCxodfy7lMalyAXbGjVQ8mosVyFvnqEtHEgzAU0J5KN3xHuZvzvN/VT3
HDQTqXNgfSvLKOfb++5AGdkSkijA2G5Gd7WWd7H5UAQEc9mg7OaH1G7TDIlZDNkPjmFs4TKj39Yz
U425xrNgWjzdwqhb1Xbd+okb1mtZf+boQo1x+MHZcV9EJNSdJSyj26t0EEcGUW2zIJowMSlRVqQh
ZtL5InkFee3VgIroVXZx6NiufGZbwW8FnBmygaYHldlUzPkwsgJPBSuHEPI2FQb8XeaTOLOPHVJF
KBU7bTnW0mBG+KurIEcdziVQp54kM5LvZEiw3hIQ0ES++utf9535erLyb9pqbIsdSiVk0x5ia+Pe
DaePqPVnhiz7YZa5WVpSssa25EgRY3hekta+qyyiCLLYiSHQFNNx4OEPfWMA3kM2WbWtP9U2ebIf
Rs0kmsxnODOR8rrPcsamcH1uizKxf8+etoEZVJH4oojkc7+ohEXfsNq9K97y92axQL34hyV+UXl1
BtL5SUkXlJ0gr2gddW5KTyymao3f2gqhaOIzv7jNnzw4pLHh7HezoblKm1JTqg+NkrKlSfIcrmZl
b44IC7lFrp/EPHf+l7vfF2L2/3Ib/XfJO2Qetbr1Ui1Vu5SUKYLecyum9sSvFuO48RAIMCl0LPAu
GynOcraYb5wQJY7gGrrDN+PStnflMwsshfDx9gxT2V11o2zqYVl/4s7AtsQTyXhdnN/gv9pMkZf+
g1FeNQipeuq9ui4E4K60JFTz1ryVrnWP73CQ6nLB7ke7ezopv7StpLwpWpJa7uquAcx7H5H4Q/gP
OI+i4+cDGh/zGikvPD0RuhZjQNjOx5gmAGOT2LuHEOgH+JXgKxakcrY9SMUrtMejqs4XlFJPx3ZO
W1wOoo7LrsK8CROOWCKCCuo0FBB/OsdGkH0EN0ftyy9lqIcGBvwbJprBYesLzVzTLgeyoPRmbzZs
sPaolLXk2dqzxGHuArMwrel7nhyD4+gTeUC8M5/Jz6vnqpS3Hm182DHEaIZbXMSXNhHlUN5UdjIL
e3a1z8HNJeVVQRStBKgzUQ7Ci30fDLNs7VPmhqCygP9JcrPRdy6YbzHNu6J+1zQvJqaaUlCM3grE
k4cs+2rdRCcB99dNLAeowXaUovNhlyVQEs0/5pwX9m+zC3nBlCm1Z1aUhFDPhsoRs5JPqIjBiiiO
ceoGrxbmmKMnjoJGunAfwxnWRg3r9AWEnY+6PAkoX84Z04KtkX7y07+KMGxaBLrgyGJXfSd7IodF
ChJmF3vzIceWRfLAs9fNlV+l1E0WO1RDGPepuRbbNfvygz5GucIpCIf4KYD0ATem3I4vF5YqSm9a
TRgsyiqC4qdJFjDg1cNK6gBBkwxQhuag7E40ktqOA952kC8za++H+1pLGVkoCSbutZ/r5UG2PXcA
/QMklUEJbzq/0JPM63/gTBTIkNLInHZkQCyg62ACXiFSJZWtrSSpb/b2yiiGoUBraILCEiqfjKqw
siSzyDrPXgG1p0tlt6K+sh/d7ZPghk6/fNYnneMl1WqsCD4+MzK7XuzlhK+xs4SJpvg/p8xHU26C
DfXZo+IxpOpMIN+s9T7fXtqdqOaCacjWGeIzTzzcVO71Ezqnwr9rTfJaMmgtV3ZNJZ8NAZPMjm5b
YXkmjyPvic6+wxu1gCx18pEBr/YhVn++2IZ35ovs4YYAWzD0dQtfpSvDZYXX/cKPD4pIvlwLCRCz
6Phe5FbYQF2+HKkfT2oBcHgbB6UKdE8YOnXEG7WoMMpMmlKuCgP30gbDzCpIECKbNPIwnICikDyg
F/7cXA3luH+EDsHakQaebwOw9CYcNQth1TlHv+JxsHUk22jklwz1o4sJykE7fDyEKvS+zivRzSAy
FxepzDrIB/Z2Y1uvtiL/Oouh39Dvb0b74uTy3IYTPh4I8jcO6vwnJ8z+tUJVaxcol6Vukb/+Lzft
V4B3ZV5viOgWo4yKQrLRGrCtGuQ11vz+rKn6WENH+LF811Gt6AmzSl2mH8IxcX1GV8sChfc9f2gv
iyVrCftzzoIovLcHzUHqg2toC/Tj37kN2COuWWkcEJsnttWW7gaZctQwUh8eygQLkNCt3ETGZquB
JD3MKqP8kHp3I9qj1YL1aTYg5N8ko9VoueqABpntWseQYRPj03Y2TXctgjPWHONS9niNO5LX1hD5
eEXFxrEu6lwEEK5wTCt/Xjsxr9X/6Z0JsnamaZUc0q5Lk5Y2pF31gZ470SltPM2hXzQhAT+tHYjX
n1z4rVbeNOl3hDcYAVCUOUBCC615M7A4i2UpQkQR0c317Wtea72hGQGlWkyjYYsy2tgO3zWjodMl
xaw+19gspWQC1Un6zhBZlw041AQYhRRozGSASxs6M3ZzdiZ7V21jBcLFY03jIBcvQ7V1zNSuCHiY
diWWHIH4f5zkQULVis5PVMG77nABN3A8gWhsGRK8XM6Kw7B/Zm9ktT4sq7Fib3MSLxU+G2kSwK50
ICSbTHhipduwr81uUjef3ySnRRQ4m7ditUaCkKRufaPCxQ5TmL8sBpS65tMYry0hOoAQC8l04X/C
1/LRV/5nZaXk4dfajv8kLfPitCwVSEG9PVBTC0JTImKdHX39Lh8B65/gOdBRMAfqbnoAVc2NMc0Q
WyiqKUB5IDS0k0F4j/+p78pBgdM1Fjixvbu+WGqdOrovzfWAcH5I0bbrNMow4zdjfOXJhLX85fCo
o+6fcrK+Ca4iz7rxcubmPfbXryxDN6Z+u2X73kU+t+qZ0XKGBynj4IMqfA+tl3kaMYXJBa3a01Z7
uvrHzyBDrKkdhNvrQb3WSNGXFPpmBpbaegzAB7URDZCGDwcvZ5bUOv+liHyU1/HNppzoRiJXiV5S
eOKG/PHpVMhnR7EyKmyxHzPKSwJvVqKDymmbuwR0v7fH7Pw5mqMPW623KBhhnWrAi94Hjx/ck+Ne
mvyYSCJ8DbNtt03TE+rwVNZYe+ukBPFbVyNcBnpDwj8jmdU7O3TMFzYqPV2c8IKFwiGNCXogGJ3H
7I7/TrO0+V4ZLXUBJNR/cs5id4iVoj9nQevKfAwjRBQpDo6goSTTPzwGIWVRibve0ffZIxq3k4uA
pZ8wy1g4+KVBhzxifMR1j3gKhhb9qxlGiq4VbY7WileXwj5dMj1CFpjQtRrwMFrYnRqv86pJ9mNC
0/QmEbiE7kO+XT6e3szkbaMfvOkXH74lhP+wytVgmpbzOX+ZWXC0pB1TlIgYn1vIVEZ1t/tJoBKP
f2JBpRNPoRH6jEf2nyc+a4LV6hQWSZ6oozcJUAjeAR/4aau3G6MF92wws0qBKWxTkRAog8fh9sxq
eUSiGpmIptYTaFPWbwn/BDM6pyufhtfAu/7CJStMDtXJqFRqJD1C9uZ8H22yXAJGHBGadGHNFKi8
s7lFD9iFaXFTC5/dubuTKR3pVqQg0QgbqDHzEHKpsrStaRmnM0J3lw9V65f7mPS1G1LqYkGH6HSp
dIbsTbAHICA0H6CvFWLMDByu5T9D+S/UUE4SGMouWl3SKqag7EFrL/Bv+Bh8HbMlrq2Ntx6tpnv/
XLvURi/x8dURnBW9ZDW2oBeo4hkTbV74mJ6FWWMzUUh+DstHIsOzhxxrZwPvHHQDIb53OJN847hY
1EyQhEDvZaxJ7++zcuAEonRosGbef9We9gCtROsc4505bOwhvjQ88qw01jx3cmuF9695txiCJabY
cGjO+EDU0srtuBJh1Bp4GrNEY4rdGMHYgvE26FDXO5GgNgIVYmclzMBX8YYZOPlwrZfXSmgybFJi
nhbPieE5hSSmoU++/ru8//SFOdOeCzAMCRNKEIg2pxtH7+wPkuLadXYGXhOrdIF5+W2uyU67PIt0
vKg+t2R4huilHtMchJTfycfYxWXmxf5JFPm4Av4TJIzPufNl/CtdHlDuZEvfA4/G8kOgZ9Wqz33V
kYVS9AnT2LhCNfxaFGj9cf286zFDf6G0ZdHDxHnfyzX3It70L5n3nUmkidzgwxZUp32prDih2zKu
Xe/UrQUFNecYT/b/dQQH+YA7g0InP1htreHz9of+Lzab/dpbl1txqcRhhxZwenOAO+bmdCgpiuae
+VoiMjtaEIDmcoQSYEBzD53Tm7P4eCIfkjqyO0kPWu++hitChPUgyYnz5nuZ9vCJevwotvym0+XD
KmmUPP+gXmmsR1TCdgnh7YFxnjZ6j0WPrQASz7fczufDQqXXNWVqagcLSCH/eKiaW4/IKStMT9ka
SPEM326jNn6fpD9YkM0jn3MFx1Y37FVCZpkwdforsV28hPbXf6iRvdFho6ak5r/Oh4sJjz4nqVNu
pmf89Xz1tKcZa3dPyXDVdgpcS6DuAzSPdedR7Qd2bsJ/I5IypPYwB9rkMXNT7adNZ7D/qPOo19P3
tsN3N36uJ4gYKfvJWweTSrOCl9nnzrKByjFRgydpScLJYG1y5sj09cbYW1rjTwS4Sa/VlnUuLTP1
/qNSCko0tEc8j6Al7U6BhkgXaT+fRYf6p3Qz+/4R7Yx+SPzKnlpS84UFgI6XR7ESOc4TBgRpnpAV
7vdnguBTIeOvr//YdM5Mkp4cAoWhs6l+/Hykt9zJYSphpcziV5vPAIwqLpTcf6yL7uo78qoLQf2B
G4NKXYeVn6K5oYFncor0COo04jSWLNVgiYz/n32IRJEArZu7uA53IHo5OxXu4TWd9kJCr/LV2dMS
IsPyYVUCUapc9gvCXUr9Szh5G2nUbG4xwGg5Um9kYaO/eeh7roO48SXP/Su1kAyAst60Nh3Hlxp2
0W/mgmPghIWj0UmRPDpi3PPc2Vg9KQkbADzv3zfyO6tJ/ek6o5Wh1g1DAzritTR7dsGuqtDln9pn
/UwSYlLY330Sb1CLjj7a5tW2FbGRAteuJ1/jL2RFWGtpMgPu1T/BIsoPREDBIGV8uFupWpyK+2FV
avgPnLhY/onwJHYyg5msifZ5FW7GDWAEVB0cSQV0Iud69D4kwp4wjhz8IPSZxKW3Rf+z0gVAisd4
bjmjj1Lzdr52JtetwbZzcOuxZiszVUHQHk338HqCfq8pTSOt1UNwXVJBJ+Vezj7z+27qua452Uec
kYOOxP4cj5RLhYneI6hkivJfStbqO2pas0y2DExmHXIqK+Ryb5xgHGhVEx2kB4J50G+9gRAQTKS/
WISyjUP1Zb7qIBaTnkmdPmMlrUuOHpjBGO3106WSwJERsHnRjFlXvzL54Y68juh946uUzC0TFkme
N9Tq/SEuVuMEcoRqRl6QHZr9K3jbq1IW5pI8kUo8t5a7oGXVvjIM5+UVPXE8tasfFJUdhtVvyj+k
uUkqkkNOe3K+mlAka6bcRjTFjQsvCGiiRh5t2yqXQmMKN4l0h6lkgytFlnRsErtcbjMfS0tghsB5
rDPCVD9nYVb/PF7gvdvY/kiv56Lzvg/hdA3N+Y7/wRQu+vr4qRdGx1gtlxn1ufAQw/bMvfVw+iVh
6ySXP33m4auXhE5wVU279ZKIuZGccQFOvbPubzsZ7HfEbtnC4/kME6HXGetAnTavifKo/zvXA68T
jYYpVcKNLA82LAaH/vsoduueizRPVXor94T11nR/B06hrQPPuMR1RLSJZ08DFZZ/WxQk/61hnhCb
VW1il8V/eYc/Rp7Jq3zahfMpjQ29tc1g9D7Reno3vus+oc46nQP2OCvVUdapEVqe6Z4S4njUbVih
tFipp37affe62u6kmId3s7rSzCV79/S5vF3wYS9tQTPCGl+Z/xjJZtSotlvc7H8dM+WbrfZF/2Y0
ncHDVFwl2fDSk/3vEl7g/DPveotkCJ+s5SuTR7D1+goWEbqEXMukEKdIiYHsnfR3M3muPky52QF7
EHFr3H+WD+0qki9TMMCY4avAhmNqpiS0f497K8G670Ln1Mvm2hsycCDtp+obD6jZ+3Ki2fhUqeTF
aJdfGufa3xGMwHp8Rnj9LCUT2RJld7jua7x1j0JX98xuGNbLZ+Olkicp39kCFvbgq0ySpkrvSa3X
+ozzThxqfY0i89D1nL2NV99Qjdzofl8N/RhfAFOxlX9ssnnU9vhD/PBhCdV9KICD8Y/7tpRwLfB2
aAqipysW029pbbDxe5NhuAuHC4PQuxLADRmqNR1c30+WIjzOd8c832asDK8wICosVBdOd9Ew+klj
GpqwEbm7ragCsjD0jHQYz1f75EtDMDkYD5eTO2LS4JkT+RMKVEa99igiDN0XVMgZO2AoT9xFqOgZ
LnbYQ4pZssN1a/vrAvtVq6LchWGdpMAHK+RFeHLK2FgZFaoBD0kOnRHfEHyQrXPoIsqOHmGBbHGc
PtomZwBXM5ZEEYld4+gHX5+pEzoDjp5CYx1RWgJcr72sODzzk5PumI3jpjymDfUDi3Vx1OULxHXO
b+oVoifUG2GmkwJGyFMQbFyv9TkeVnTdJOpIwMT/aDA1vK+tCi3uGoVyF4zLLsSotU5J8WZR0szW
ZY4+/90qoQSa95YgixEEshix9c+UkM6GFs1T8+Jk2uMs4+9NbLzuvP6yTYAgxU1HwW/rjul5whFo
LyBx5dSeR/S61zE8Yrol3u58rjwao+Abz+n3ka6O93SrAb7vQwcco3/KFUpOzbtFPjXH9FSGxfx3
uG9IDqAF1SQnD2j+f0Jmok3MeHxG+uqgqG8cR6VoS+nD5PBKjt522xcS8ys4DfdVF9zfnK3AaNl0
M+k5ES3SEm2TEyoENu8/O1FDJao8XTrSdjRA3R3DklgkkgXuLegdhqsmvPapOQ6D7lSWQ5BslnSS
eXhiFrBRflhs5whL7z5uIepms566fajY8UpRW0t36Z+lH5yo930+haySuRnCF2j7IwgyO2sQY9/u
64Yr/mAMF2Pt6libpm00TxYtXxOYyV3AmBiX3OIOpHwV87gpEve9T6a/TtA8LSuPQBHMopEzrIwc
TkgY2lky0iHSm7kgI1RoVym+/V7DoAfVGm0E2vKWOa0k5f05aLSCm/nkESn0Eb0f7k2AyZ3c8lT2
+yesT1A2IyTpVXxJPW+XxKGdHhEMX+8ydGIdu8wDBUTGpLqv6+U3v/MU5rVGp9darCJcJcq7nH3g
+OxfieikAeEC2iWz+qTak06bY+oerbHi0Bu01DdvvUCoP7nAoYncT/x0WJzmwggjbib5PM35ofre
VhX73oI/jl9V7i1YPjlKXJOi/IFq1XlXwDVraxeU09WT+NPhTxlHlPDk3OXK5JSTJgEugyboUoIW
qEw+ltC6WMFffDwbrMuaFACsMW/otDnN4hLLK+Mc3rddD8N4x7qJ97LxICtezqWSdecnVUwpNbjx
v/0t+s04wwSreThXRsWaDUlaJwpkfUzcVXqa4oGFCjMDfTVBvzho5KOF+2Pl3dqT80XHVWBv3E3+
e7wdINWrSNuyFxn3tnfJ3uooW7jX/Iny6UgLbN4lRyds6r6NRCBzA6i+gn3yaLWwH7j8zODiR2co
qnlOQcAPz06ZW14Om/2ZtcGUJz5xgbyi+JY8R1vNhzZu4kXpudUkLd3moLXBarwIAZ2mqPCLJZ4P
TZ9t/q68T5y9Mkd6untvumAnYQ9egNIMVinLxov6BINRyg2iOte9Az2wd2hhFPOKTsszpRdkaseE
2JN0RQpXTkTki9ntWcmce/aNUh5VybEH5YF/NTov/FRrqQhmR1MzN/9GeMUGQfJ1HBSCokrM3aKB
1iIEUtg2Vg0iUiBUM21fy2+2e3bAV0yWnvbsntjqZNyZqwHVSGb30ikNNFgjO8jAgWSiL/iC+Zpv
SecQyzPnfr/ooisAezV3SJfX6tMvMeOIYtrnKBgwIbdJcDKzUUUZxt3qT5x/3rZYwC09vVK1Iuy2
scSc7mO26YGMYWBQxnYlRGHNG9w+crtw9SRgg3g81i2PUEpWiWMAwkFkmZmkL9N7lBSAxJrs6Od1
xPEhowION/8J3VtttBiWtVk/H337TgPmsMIrPYfglOvg9sWDjuRmGYSgR7Bkq3GYT5dntgAw9bhk
+7MO7z8w0wNe3zbBz4VJjEanQLYQDaz3qlHvu9OqDsvnVpNa2Dds9qxumQChDX1im+B/+kpT6/f/
myCFtPZkm2+NfCtJzioAeWzkm6P0ocY2OwhNz3EjBIoRBPzwj1lvfUtnAtWOFx358JFoAJ8f3URz
2PTeMvL1EI64VlsxCeXfo65E0ysN+OSh+1qb88ea+d4PtP9oILvjv8RCf7D6mqIxSu6doypxlDDB
FjilFUZVPqkdCI1QtGhNZT3Y4wceGad3pOyTCaa5anfGz4vrFoDWpdKPMHRgDpsWD93jVq0L7FwB
VCLmDaUfY/nZ34kPyi4GdOUMWlcGaM0a+vXRgL5R/LEJf2YuRcTDPj71CKZ5X7bXhJMUuDJC2cpP
dupb/T2N50EmacQiMuq8PXkKerWKnCCGvw4tcYeI3o4zDt0MByEVtdW/YNTxR24G8W80T7PYJyif
CSLVN9UA3ULvPOht2GPFTA8vTXeQ5Two3WKBGOx4SKngQpd3nMH/MVshh3X3NN57OX1q+8Hrf+eu
dUZ0vNHLYhFvbja3DGEnqTO3zXrh5ZmvTRs02jzSFP57i2B5lHz0TuyZ9JwN/Hd+PFvFOFpINPk2
EN35MLIFrS6zj9uguV95xwFSHsv3nCi7UEf9lokLDQXTvdBjYlswv0BQ2za1afW3pTdGK0J2SjQ5
cCwYpLt3PDeQ9px91cVxsFDZN29sOl/sOeuK7FYrI4nz1CUXcctDqK/TEyFfVR0qsb/CDMYamo9j
w5kuSEAXZyqrBHhUuujJY3DQspqwHr3mby2s27gCqSHlUzdUF67uygZfjr5po8G/8yVW1r4wMnMo
7VCYkdy0Ld78aNrhTbcjeZv+EoC8++ta9fpy8UOIU+izDNkk4ZiuwgKsBUax+lCw+8nBoPw9ZV7/
96Eg8cjniZX5gkXc2R4UV/mcwU9idQY7pqfI+86vTTOuiD/QpminnDQeb5S8UCBf44ICr4MbhAyw
oaFS4VNi+/ilap/JXZjdp36ETefqT1XGbC0dAPHl21WZAQREnzTpko13h7Njr4G7FTO8jeAVp9Xu
d2cMaJgRt3gYneur4pdznd17qNQWdlf7khhH/W8du89aYzugChSq0xI1daNjbXiEpJUP7K+UnK6m
ZcYCmKW2SxyKFUmRk0Z4Z6RWx3iu7/dqhGBVHFeeEzp6Nl3Q8FpTC2bqxHUxZYlM4MIKdlxsdG2n
eKslJodpbHHlyGQvWQGwSdbOi9dG19YkSisBRSTlKVuiV4XY9Kv3d4XX41f6lKsvBQa1xyXTpAHX
5Lz6Z7KLdRyYUGSNnB4RQ0hJtgWOKuYF9mT5/xftNxktMgSgxrknQxyCVYTCgiSD99J/VySvhvXL
QOar4N+kpPRkFJw432i/X98S7xcVwNlwAzoovZKemaWuj0u2x/w6pJHAWTyFILYtXdm1TN5R4OZi
mGyRDtB9foum/5/OKfWapDT/+J7u30BSJHAFUbt7+LhfYd9RGH5ZW9tZysX6y6zQW9cGEuU0suie
YHiuCKrQ5qDfSVO1g9bIbturpPbpogz4VqEPIhz5lKhOPabHZbgnO3gTeyoAnORALh/ECa3IaqmK
+J3kqlFU5L7rMNj03OpfsjNJqKqNEF4kU6pXORcfb9qbuH0CuPDrFx0bc446B97SCwkWGdKWhTBt
O56LomYIF+SqOG9cfISXko43Q+NFWp2/BfIckrUqwjyg6LG2FJQgbYTkYqGdTZ03VQKK3DqC5UWU
WW/f9i6hsXQyyz8dzvbGko3lm6r72pdvcG7go5RIHS8ZxKq22ZmYUrkyEfSAU9nmWTtCfHvu9NTZ
Zv/yEdleGWNZIlRJcbe1diuBE7t+DuIe3/g5aPnu8HEAlv0aD2VAU2SHXmURl8TwWkFfpn7URxY+
Qb07LBi61eiZBk3hRxXZlKgIUJ7Js6ARxXIoUs6oCqqGrMw52hG0SuEDzTOYts2wr9I/BCg45xLh
58OgzTAYehmMM7pLA7hMAZoRXTeLF/q17HTM+XaA/8C3DSXIDJqIM/aoQtgE9ZYJZ6Q7mkJ2L83K
nDBRE3mOq0LY9zCzCw7PhstqiXT+tmyyhlQCD1uvFCtsNYUQF2aXUGlIE4T81S+N+tg2ro4hVfYj
KAO8L6jTcWHbyAJ3T4CvtbgqsT9uP1aMnaMsBZgza4GnZbnl8u3Y9suk8x6SZPmQsG6yAZ7YlcDv
5Zu3NDVaQzqLAmMRL4G9lsNc0tHhOc166d+abkV+0LRezMWMF0uQJBMp/5WEi6imPbrrKJYVFk54
4rTn4e1O+EA5M/rC2h8NS5wFM9zlPxZiIgP7+77NO0Ngjpg1nOFIbwGMHK6UDObtehwtnzc7cIP0
58gySK4S/ewpNydxQO48WKp0mXeSWscaeh2HHI8e+6a77BDBaiONpNugJiCW/TlDkGgu0lA3A+gu
qdLUCTpDCPE1vN0x8OMvrOBoouxC62RnUa+OZ5CKIm5s3Wuq6RtunYxV/CMHd2bIqkpO7ghUlE/V
Br6pAPOK+4ozBW5miATa98mRbPfaeMByXkRdquP5MkLw+JR5A6aUHF5+zg7cVbiR+H4FyIYxna/Z
rFn7hbsntfVyQ8Ei8PqJFNX3k0gl2RV+uD956QwlwsM0oTyUokFJZ9C29U+fS5C2e7s5+pj9qJAn
rJ6dJeDPTFcJI1tKi4g57Tcz3nejcIOVCgTfj2SZQbZFGF9qwdcDbynVQb9x+J41Z0f7P5IcDJ+4
DQpfxwwySt84rXlomAiysn6AQ0ZGXpBq07ZOB36GL217d0UbthQFu+6neco5rl+MotuxxfYJrmuh
LYH0mBPIavdomrJBjVToDZeqGRSXYBjf1xhlsATtR0UPCTm80QdSdQ0JkNjEp9AAbuEkHBNDzne4
Hpas8sHFbLssc1H+n+RsTXGwvV5bfOW9PP2MvGN/GCcK11wLNxUTKhzHgcB7dLjHesS9XYLe8Pi4
3IGzM/zjymoH5O2/pzmhddIXft+eptV/TdgijOY4OQJjdQSE3TGqQu074vN0pJaRMFkf9BI7DQCi
LYfGK3qqb/ehk5Gk3jdFDcFbuGFmD8cPZ02YdbvrlcJhQ5lP7j/x97yc+RQ5vNUSNrmjvz5u4ybg
CJ7pTVKiXrvLF+swCAFotRNY+eRIwQ1kdkJ+2SUYvYVVhUhy4HcFf/3V1usHhvbabaJfwhGDnIzZ
5DSa8WFWdH1S4TVmWqXgJn58iqC6RHMqU+TtoFA5vH5uEMH0AP0bMBxeS/IkWtc0pNactuFycOnv
ducyvN4ra2hI8x0XAUG2hXLj3OAhxG97PTNJKj5kKo3sVK2eTDzY1Cj6MpDYaNdpzyy0m4m296qc
+xlPNNklPb4p5HKE16tL36y6RxJnd9uurFKSb+T0mz8V9SefOsh+wfCxdogAfwNIrmkJZs+Jyfe+
i1nuMttrYlQyaoxbLDzJ/6D8hXR9AyLrNW1a65lrYtKsbHHp0/o7MLjojybba3dzvmexHx6A87XQ
iZFdVa+zGYRR+FIaRFiSwqPCC9sJql6teD696rEr5ATbtXQwGzTP242O9ow/5Ryh9mAVD75iCDQI
r3X3yJNMLo6ZyW4226+GeP9qBiiCqACBmyAAaJs8Dewr5lfN7hnecnOFhaABMKBdQKrw2Ty0a94y
lo0y9qxybZLqgsjf1cRJdQna26Ebb7SGjfSGQjm5lsmS8QMC51h/h9SN51jbXc2Ux61UZdCcXinE
LHe3f6bxiU7wzT7pHp278XmftJ4FAeoi42p2IeqYCsrLh9g+qmwR1h26AymfVIg9WuCKDKtAIXDt
AS9LRrhA+dpB4CRWJ7SGvDskgOcnZ17ceniCod+Y+9jSETN3YU4fveKeEP4C0M7Krrq2cGYMS248
vna4DjLxLpcAi53bXHeXBWceqmi5pSaI2yOm2dsR8QtNSCuT8d4g5Myb7MciD8WuNj4vjxQKcHB0
GTfZUlC5iw6bUFhday+5g43VXiJjs5qxETRoWhUnsCyBPQTQ16inhbTUBzFHJOVaOuKS7LrwZGP4
c+nXhGM8QOCvmaq98gd0vtXifJEHijYll6K7DUmTCcOb6rL95SDx9XObAROB47/eAqIqLJlLiAtH
dOd3qSsYKYJOqMZsAjCv9rA5JZNgUK5wmDH3x2x8vJ5BTghYopL2em9D+gE0qrW0vbB8i98TK/3y
thpBWFILbYGvWaGxbSIBjYxvRzpgYezLw8ZuD+rhzFDPt22cFDDO5Fl0AlucCbgyP/Ap53VrN2xd
oLV1zg8TxblbvIa3uumGQk3qIbZ3bx1+J3G40KamWpzH016kLz5T9h3Hbk3m3JfBw4M/5KD1aKZX
vAYzZZn3zeptCr81hgzbYPLBQw6Gyp2niUqKMZ45zd/h3WY4TaDDWebf0Y7ikW03f67Pj25x4dZv
l1JGNxOBrGza2d96/G1qTOuyryfwaSncuLbdDqHPXG5JnYFwMQPXQiPzIZaa+Log/imrwn1N5hU2
7SRQaBRY5wYRExDfGP84niR9k4eikSuRuHJ/AoNKFO/fn9t1NJDVqFyKpZNmOAni6uWhDAeQZ4JC
3zMKuv81uZGNr2wf4Jp1rT4eDnyt3ecTeJZLLlpK8RiANT5zMpNC+SR0WcKGxMyag323byMctkkt
v13RdhBWuoyhFlKJTH9Eytw8BiDBRMzW2evQtYa7k3HxuhErsrQ3IV+R65B9bl5EiC23yqFMoQJV
/0Y9YB2usIKrr7TqLZVBb616waav+u3Ke5vASezj64YRyrp607ty2shQnZ5uOvm8FSiuDoA0mz2S
hJ5XGgcZX7l815BtwJ+LsKWrAP4Mr65GvEPOFlqRvsC5+4n8aMWrXXNtHi6XutSQzS78tPMW+f7d
YmlodsCgsdRjJAt7RVw0sm7Xq8skD0kzrP8EQ6wh7ezSCLM2KMs4tQjoLUSo1NKq+vgbJvjR6Ato
QBe4Oa6LjYtWE1o9bVsFZyNGAlzfFYq9nagQPUCaroglb9CeMa90ckg6dD17RHGxw9OnvrhVQ0bJ
obObK3M/Ic5ukZJbLiDDX3SsYyEWQaDzFTpglPnsizeojGIao9vOBVwnqOJobOsOqNzbmAMzaoUk
/uwd0oOQWdHra0d4U/dRMdSJ6VxNgyPCfEr4bIuk5RtpCPUmd6PBlrrBwmscawHA16HNrY8BlTj7
bzlHK5QdeJjBRrqBNBWuPYpbVTuMOCnBSa3t24wfq0CyvTpB8GCSsNokT4wfG5chYsZA4r04ua9K
hJAyldCpohpKxTorOAYCu8tjoiNB5qWsIcLTo5y4XHWD0Dx/d4FpDcQnjn6mtWCMQW0VCvLa90nR
tnjz8/Qe3xZubwdI7dn+QA/DlPQTzgU16WDYzIOZshfGL6Jatrg09y6N3oGyLqdLdEfbYOR4sLZ/
m63UJOPOAefKUXebCXkk4q/Qw+3SsTKH4ABcTb8vGQzNyPSC5xYz+EQHNIWiUdhJ1mynstjvMIZ0
jx4DAw/Pnqmn+Nj/bqfWHbvzRmclbi5/nN4co54/1VrwE1feyD5twLkulptEhe0myTQeTP/1twXV
QcD64eaSsGiNyPnuOtT2Cig/7wqd8yzYZKsCk8uinSgWP6ayMjh6MLWUD/V9jZbc7JyGVOMNhdXG
GyTMLFXlj8JRPN1eXphBbIe/kr4uejeStYmNNb3llZ3KZG6PskmrYvJA6kX3Tp1P4+gItBzbt6t8
NVRgFCx0OrYXUNHYbhYKvEy+EMORa759HWZ9Gv0Sukzv2ut/Iid55PI0pvhJ8VBmkAXKvVzVY533
+85oHR4X7PyDBcStXIqGwKPwe+ZTsEpcFYUZejYGdbWFCwkyj+Cd1AAmRWuXTPQxGvtr3iwUnmsd
LxHjGMyTfpvKPR1XYzEZVTTcdCrw72Pt5P5CDcjIsrnA66k717kI4zAHK0saRHVQ9BvWD9Q9H6jC
ecdYF3LXZczmXdxPfJxPqW4Kddk0IGlfkvSPO8RLG6E1eiizPR8s2klEhrAFiljPHevOFzN2qt6k
6Q6/v5GvBeUYgAd+JUy6JFbcK6AA2DcTA8XcsAP2JjRK8GMmZByUYxq3JJM7JixTbdUQASXKWIl1
i1zPhMEMjGQw0V+Pcf8biMh0r3kZA4hPrUkOn6aXas1NJKj3Zcr4zS5tTt1ZJMhOQN/zbSTGA7kq
b/7sasHAig0R1AbNFnndDsOdicz/YgeGwVTtn074JRR938/vQr+CQBqj15RuSGZsM5209u/SldJL
C2ukcZVwXA8J32NhI+eSU7qtdEX/tPxDHQq9dOTb5xsxW+oXBW/ixeC2BV97a1xq++PQ08a0aFoR
ulypqNHRrhwHse0pH1glRHC8a+NsZ17wLdgtokhxRz0Zvyv4SxW53p5rmHNIC56oLeB2IPpqEH60
lOJzs71kElRtbOce1rmmhDwdtWeDliGCiRPE5RkcVBrCgaH/Q3BGNwoRT5icS/3I+cZhVcj5nsDg
BU17EipIURLzQQuExb1z45KizB4fY2mhV4ySsYXt+5PxH/PSPjLzA85yZAa3397lqgkuzdvBdUmi
mfXYbas+FQcXWDs0zBinS16d7pQ82BOqypxpW79BQxFtiwxsmNYaLno/aa4h6Lj4MXl3yWSKNQaD
q4RVbq8Wskk2P3pGAnEIHToNXdR8V0/zTsvKO3x7bZB+8fFIVvBU4P3QriZ1jKdjToJvdyxKPNXk
9cC8snvEw7gPmN1FNFsipTvQ+1jPQceuLIrNQ+PeHgdtsrvuaq3xQ4osl48qd94DvuA5umiOpcie
ajdvAdbdD8waePyf65W34GJYI6LTJ3+qvSkfTnCq1ySZMFHqcPpQrG/51OxHk/gDAUQy3jIufqmv
d1Nrnly3/g+Mua6toSk9QbPul0d7w6mflDwrRQf2BxVgL20NoFwk4950bmXhkthBoSZhUA3+vOcO
RQm9/kSW3VCdlySFwNjkVeCHHfe1rAIPXPoBZYzh5NiFh/xRupKwFsB999E5pBCzUs07tGkrvThH
OA0LI7wYSsLEuMTNMfq8jvbCaroAcdwuaiSGe0HPGo+fWe/EaChy7ZXzpy2eMK8NbtbA1YDI/MVd
5P4cjMsT6P+pqBsBx5OJ0uND9z7OwercZtHfUrfFrqskNgGIsFTCiVdOKzi6Q6DCB96/KmhXVKL0
qdawczRYdCt1Hq4XHRwaH5OnfT9FcCLduCqLwO1CmEL0Xq+PhfkZ7LuDn8H7KMtnucYJ1iBVPJ33
KMmXPfV1z26vrDSgDc+Jfptqdx8wP6AOSL6ryU17U95JhICNoU8ALFs1v0RoNp9je0R8pUeoP2vo
qZI39vS5qzLl8wkfEym3EXYGzAOYOMvtQY9BmSLi3xC5fGpaKH1RhL9l/Pv5nuMerYDI/QrKgadI
uH0QR5fb16kXML4MbvEA1D+52a6orIZTEiQlA0G/z1hPXeG1NiY4YgQVNPq9dPMfv9mjpimfzWEL
Yiqlc4ra3vkgP90wMK+nIKcZmEprfo11YX6+HLFC8G4uxGyjiGEKVWI3OQyNvvxQVOR9xyz4LCbi
EOj+lFFwBFmlBm6cUNGCZGZXSA6eb5FUwQrVAiPeMF8ZAwykTCrmvHs3fFTH4734zccg5ik/oqqx
HdD4gtWaeNbKktoREeVwDVdhR/P4/KfC2pQrISt+PuokDEkHVFcp5ANCRZfyvq3cwFjzBE0qC8bU
KxGPxYYmS4C1CbeEGACNOw38YUxdIGDJINndBews4gZMSXlTz7heTwjfTsgiemY8T7kQEm6S+RsK
TmftYLDViM4qd/iE6Eccs8B2vCGHp2braiPhlzUrY+7h9LA/YQrN9r0ybVFvSC9tKu334LHL8C8u
uofdZfW2yi632ybtga2xSnpdbI9oYOdZsYFg3w3ug8laFhTe7gdWmmEutx4uZAh03SOdB2UFe442
w2aJMzgcPZrO3wP0Gt0G6jcPRrCenq7En8KrysJSXfkYgtQ0Io7ABOohTXWb59r88Svh+Xdrp/c4
GCUohkOGel/eA76M/3RD9f765Ty2lgLkaB8R7lQwsTNfz2KLouwZH1I+1Hh7dC4LFvEdMaEQgClw
QuWkCQRoe6SPCEUUmcxPlFMCLe1YjtYmgSvDtDir/SkNukx9/3AUdAu/idGhjaJ/uf2rvghCJ+J0
a3wndtvWAud81CbdhdLkFRG8GC3IO7ncjL8GtsKsgoG+lQy78DR8ZeTU13cZ4HCpxeAKX8JQlUdQ
AuGwcisK0+Il4Qffiv5pWnvi/N4+oGjb9DDRhGDDyktZ/2dIpwpd/E05Zf7OI2hK+ICafoi+cMja
LDc65fzQ/DWAf9gAU4F6dHMM0RC1xuNhDqa0ahBgfSEq3/FVGECrXYPg49+3p0dpOP3aOK3+XUVN
UbLKjbI6CH3JfyReK4+YrS1Mq5zh2Cs65tCxhO9+peaNSlFnUttsDTeOeQbALOMuAXzdTCUS/yi1
CvFl+H0QCxYA773OxsfbGhCcY5ySvgoeiKisjnILpEosU+cOYIIiDdYrpSTmsSjP1jG7Vx6gv0HN
ZHmhWhDyZ9Ak2an40IR58QIffg4YmFNMPGNHaix8cISqEdwbbDQi6hg9vJUrFKp4S8Kd+Q3kB84H
6qM43dgrDDEqv5aHSx7gaF5eQ8RAh7gPfddrlz/rEz6r5bob/2A71RQ0VkmHg4f9YMMAn3kz4+51
fnSCYuDrS6qhG4V45Onzy8EREIAJIf8BQz35Hc5xuJDI5ZJIVpwi42yxVwF45XxP6cqLG6t7SbPV
Vq3dkjxNj7GVBuhC7Vh7OpdJlnZZidlhpbU2usH9fprNg6Nr5OZ8ywMr+srmAbm5VN8qMuzoG2X5
hAd4Y33icMJ87yPr+HMNHI/RfyEV2tf75X+xB7bC3Y+kYgDrPm6F2mofWZmmQJx1mXO6fOcvEQeg
a5S5bcOrL6bK3FKNVaVw3uZ71tMceoeAEwZ/iN9gvLLGJSdN9eEGbRAsspMu6C6zlrr1DBmb8K7U
snGuHqjB5fEELr8Eld+lBV0McFjhdt8+99p3+8dDf12X6Vb2TOMfVhYCR8Ou1zrwzOE3KsY+tc3Y
tkN2fu3C7cawgKR7HWwj8oGvO9by7FfsADgpmg0dCcHWuUvbUzDxXrFJzFKCTa9/74Y0lPClSMk9
iHyfVFGczkIatmAADJkylHT232ygaaDuIGPXOVeLdagCZ+O+C3xJs2O6JLe58pY88V5O81aKvIeX
keZky6vdTj2DT/gKwceFSvjrIKYcPpbPsth72MTrYUssNo6ZMTCSRdo0OlmT3bgpNI3p3ptk6uYf
9Q6FGK4wpBq1uk4XA3/vRswC3gAYHJ5r2xy96hfryZ4a+/j851Ig2zXIA6OokLeBZpVSdyp45iV1
YRkCS8v9qMVaC+2xvIL/FgOOi/qEAZmjDnUxBUKYc4ssrZrM4F2EQknwCxmge1pu3GAvT3i1AYQP
XHG2VqSrnjnsjZuFhtf2J7URN1kD9xzHN1MYozfX3U/ZnMlMyuiheaOalCXPlsB3P8fIFeG4LEIJ
8AEm0I1LOlOiYsxMv76DNlo3dSjVhiTUcQm9YcJXVXl6siA4vuLy7eNPPpwbpdd73n93xWDNG0WP
T6XVCy9Z9Pwu1O7q5VmeEYRl3Gz/U1pDK9LXjKNe4bQnd25V7hJEMRaFqYipcsxWv+1o7E5MkaxK
OkXbQy+MeD9ObDlDFdosxHnDT66GeDTIj/6+0pb7ctcI0XE6gy+Cl0pM7gSpSo8W08hk16xkQ/JZ
IDPJLKIbh/Nqrlq4bb+7ORWuFReuNIKGxPT8ZVT/ooQqzDWt+qEOsbEdyAgH2SgbAHMdJxri9BQS
jio32Q2wFpjNNWvn8k+zOj6/aC3P2yDHTSQHhrawbZlVLKtW5JlOJL6GIt24pgrBl9w1FBjJEodl
cN8PfvVw7km4YuvaU+7hzavhMmCntt6tEaTFP8PDy6EwSPyrc600Iq5JvxhmxriQlS/xA3SRaUXl
x7IDpeBwDvqFtFGZgpthB9OBembJbPP2SGbKZ6YH26Gt70Fe/JnjOP2g/Uwg8KOHBEkc36lqd7Gi
rOffe6ttQa5AwL4BJ3qzPTNcYJlQmSa01rRc34KMP0lpFZmPAQoKG7MuSqwW8pXRaCCkVCOsptdJ
0qoYvC4JwUj+L7/xmY8Y37W+olxmFDWIHXXWCu8zlmgNc3EnrGolDvQxthopMw/nYT+dHrUw4gjk
SxFoZzAlsiglggYYbiyQICw39U3fDSPRCWLjnG2uxMuH8fDfcKtrl2Ing22jW3UkIz0yL2AL+87J
WGLHyUIKMFr0VIALY1h6FWecXRIvi+QVSceycfpNKEATgBnIRPaas53IdsAw4kH09qdbvxoklYdP
YZrBiX85ysBJO3aJL/AgSFZPqIM2CK6gORKLxAJ5kYhLjD8fxgvPgxJaQr5N6dD+vI5RZQ23kKcs
fo/CJZhe5N/dAdBSDYq8fKmF8V99gDW26ZeAtI1Yn+YylC7SfxPOKPFApNiPfLDTqJfz5vQQgzHs
Rao13igK0kHT0RWJaocxR+rVLOt79ijOzg7rlQ2codrxm0JpxNZoqsJnof45htcT1fCoGXFaDpoI
MO8jDQUi8t2vvKuoDoyIhZM9ijVTynk1iYcgsOZo+wdn8gF/KyUe+JgVzyISgiTjUKopXNPUPYWS
bGoSSKcM7dmiN4OTpfvMBcA5F5mHVJchi8I16uLXI2bb2GCV4OMKG590Y1B3KPprrorF/PVtIakU
BAOBw43BwGER+usjq/oY6sJDriKn4UJJc7p4CIv5EsBGmh+QRU0VmY1jkb3lmhr2D8/Y6Q9blJP5
QK1C/rvfEPE7elT7CxXf+lA1XhhjSMfcjqEl/rlOeaRSl2Jdu4cylv1UFdU+qWBuyG8419N54pj8
w6Qscc0LWBCchXQFGyOdtjnfKWbRi4FQBlDy8yHovXBSuf9ty67wABqO0PWOe9LxkHkflNK6HzYr
FbfJwi68l4AocMrhrKRD6nTSbhVOqhzYwiJDwsSDOnX107uHwA9v7vdwrWjBXL/bJCcjV17RWDX0
vXAsu/A7x0v4AXLT773wp3YinKc9MPDDLZbLFTBQgmZcgrGLQqpAxCCsmQIVD1VkUiN34f94dg6C
MeMGiqaOCwQqAQhGW+IQPQlh3ne8PMZj8HjTtClpkfENnzpM6RLl3A8FFqrTKm7N0nG+Cz2iPmYs
C9I/Bf4UR3kwFqyfR/tfwAYAkY+WzojgpsD9+WET2GnLiReFaRThT9tkHva48i9Y8FbNxkfZaOoy
UTJrP/EdjfNpb0vasCCBU41If8+C380OU8WHpTF+j4WEYvGT01Od3uKkft/VEwaBhlzV/xL+cZms
eBh78rd3Jm7ylUA59y39CHYU9c7IU8NmWIdDwHVOu5uIXc024lOJlclr1r672oeinyhEVs+qZOnB
Fp2jjUovlbaDKT2CySuHBrAl3Fb6bxvnNuLuokbfhW6AwZ/2wqkE6JjA63/UDpndkKevbY+LbgX0
FJDR6pmVv21hPtNSOMLWl6y9UhyGJHf2EZE0bIgZRgkptd5jk8dnKyCzCiVoyz5qBp38e+/lQaEd
SnGOuGqZezvN80xEXm7q28E5ay+HWwn9iI2oB4FFFz7RDQoutnUuHWQTOfng0ghg1FAovt776WtE
Z0F4+8nmAmIV+sLNIZzRBS1REa5kBYOzPqG6b43E2iDmbcScLvxZh3f998pio0ermbG15tGZ25fG
0JMSBkZ9iNNu/6z51hyNsIhycjTp9joAy7FIHVcRdFW/rkYZa87EghPO1T2zNkmxYENas/w56QgU
2VWvFpcMgOoXZRaRKK2IR/Z3wav3kHRxxhRjdovXs+StVNVExF9kkkDcDqgGKKTlFoL9va3uDOD8
/xt6y+7ZpcoRCMwAiayHjNeXjpo9IuJnxj4M0CT54yB+c3nqVirNBvJgIjteQ4u8SR5KKM4XN9HN
u/puEW3Lmh1UIYcEZ35GCuBxXPidtfsIPKKigJqXmlopE4rDFV0/45DwDp2oE4pvEOCsZdH66Cc8
rambuGHnbZlTCa8iF+OiQfxfX42kZ3QRo0qu2MAOYzP4ft1grJ821q20YuruX6smAOsU6Ru+HuJK
Ml6dHdghhxKKe4ufMeSmhGwApTpJn5uPWMiZg+07+yU/LQ8iVTBEecjssTIIl6cZ/ByOQg5IxQLf
XnpnYT1FDOOdtHfohEqw09vD36KQ1D0ehrXBsxlQxVyr4DtNlRjIFPhLcTsHyhs+5Mem8Gk5fHol
Jhh+rs0u2MecL66nn+NlbSdzIXMRykDJat5OyqAQXjkw7CfwBxYokwEjI035bOxBpIko2IAzsJx1
ku57rO3Ln89z0/tsD2X6BX+qG64D7yav3nQXExE5SxgG+yjrdVOQY7Dp+9ToyNFqUXlirad3vZj8
ebaunUaVhH5RuuQ1qn+xMM0g3I2vDp8kBsbuaHNwv1V7x03VkzgTa/HxDr8np1f9sfJiQ3UwECfP
r+exPvkye07jbznvDAYuMj0MX5n8gzEOX7MGU6nHnLmKwzmnqejR+AqYkcPGOA+kd72kKxipSWpE
r1GcoEKd+u4M8c51aH7fLv8VcbVtP0WgKLzCgQ9CEPYQHJFHzcxX3q0m0cbkjC/91B0iRxHH+IeT
mdHVG+F3xh264d6rL2a1/+MYUlrefVMtAikX8OMwxHiWsJ7UCrTL4SIT1kF/SY+NUBlqchofmX72
HvTb7+sCHQLLPxLXYActkeOo/j4ypv/BoQaiRexpXi4nZHngwurxu0qXoNUMAhOSX5Q4ZhxWsGJj
XA4v0TMm7W0ZLtpAz2vHj3/xt0tluDmZCVGiFEDsVBHBlYtdwTWA7RMU/BzQIaqALeQOuWmnBNd6
f1di/e7CLH5TqFzckB7FU5u+kxfW8z1j/kVLJqjy/++0Jh5KIjSAd+BtecuN4c0n4EGVjG0hOOBi
ob1P0qfPk7kBvGqekLxegODWm/fkdbLCTdQzXILqu36nUgUYYrUlZgrfWi1YkiIo4d8iQksnCbYI
otztTLw4QNaAzBHym50s+/Q4/nKNmCleZ67qKChxiejn1eN80puD4g3dbyzBUlpF4CgeLKM4D4Mi
tmuAlfXnpGFRYzn3HDSdUqXQUdKwuuKXMswYUJyie1VfEPrq4c6jlIYQml4/0iRnlqt4oBjeDzkV
CsJxlBuSxy6HthmfagNh+aGwD4qTy8nkJvpl4h+ivRKqga46Wuub8OofpaLm4KBifprxf4INiFFa
eq1gdFjQNdkEvKnL2qOyf1lDWd6jKdpmvvUZf7cRMMQzkj5MSSSw21pEIa84H/54gwCUb7nqZppy
axUAv4x+IpJxz+DDS1R9n6HW+gjeLBN3alAuRQyJeRz3QyzDHFPeBRgS4eP1zXFGvms80oQmQOAA
oxJl5l2FVEfWeSdHul2OHE7mmaR6EZfumsO4brZ4bo3ei4CAI07bsjPouMeYReRBGPxJeIKVOMxn
1OEt0zsRLDlSb/fFb4gOIs4gd/4y3VIjP9qp+z/SSxoAXsbqPTiCBvAML/Xq2CoYTlFbgHHLACl4
6VKytRdQK90jfurrwrKJtwYodI6/jWJMMjCWpTYwSQMU1NeWpixHWYq3+IXnloMoz5UAMHNVdKf3
AEGot+iqdavFyELdbIRc8cs39Eb1CVLGp9Pq1nrfh8FVWkWwfT06TyPJBI/UcqYjl651Vh6vcwdI
r7xiub1j99UXUCNsNPcMFUzhPB/+YWQLZJJgi19+CaRQAlZ2dUnHw/GN5sn0a5MvJAi1LmG1Cwvv
bntYMIKypoZi51yt5x6SStsXmtryuypySOorNYyxkC2e5Co2EZQ6o9L+qly3qnQbylP1ab3GxVtj
pwK7tmT4bvaa65KKbZSVB0dG5H4prgfKswBtepvEfEmCO3YukMRdGohaUbaYD7whLXNg8hLuc5RU
6o2XHVr/anSItxlDGnfWikE/YUfX65esiLZFP8AnHUko5k8/tQ6DUUwzuhXh3YkyqiTez33mM990
zoZp/41gGwgMp7o/QNcmQjrs3mFU1Msq10QOwb9qp839WzvOS83/Vvh+qfDrz6ALpPHwGwCFwWRT
SCnikebc/Papg/6gkQgGC03f78fEQF9Q6n8k0/UWMWzSrLgvNJLmfvmAw3lHLYrFio3L4fSGrCut
71nz75xsxi0tMDRTC7Oiq30lhjcAjZf/pPgi82pk509PsHayST0YmhZaHh5BWdv6juj8blGMiBBN
pNXiydG5bMHZKcot7wb+LHwktqtxMAaSlJk/BIrqqY0/i3wXjVlaaisOLMFF/lPdaasr2YXAAoQF
Y5UWE6LQ7v/pTSe9wioGiJ/gnqZNDWRxVoi+Ikw0fXwXysAyHepP318z1q2XyRJBreUSLte4nCqp
tN75f59YdDugPBmn34G2kGRfFBOYGo/Xyd0fZsNGawZEpdqjvtsysDO7PusDnuNmbxlq06jXf1dQ
O0UENPdA4B2gnx6H7LrtwM1SItLPZzDW4WPLs7V7lZD9r4k61YwqZjLjp+tmxCoX6UfgkbFylCa3
V0CYkIH9/OjM+bDyNiJ4FyssrvNDsN42hZK/jZmOvS8OhWvSFzVpAXNHo0oy+iZC3K9QjHp1wL4S
xrLSyA4RJ8B2JuJkVDRy5d2G3ci4hkGeGz2p3X86vqvcJK7QFqKcOZOAC/RtYLnkbeDQCylSF+zP
kwXByVDAKS/UdaO+X4YrH8DLCBxkei/kh/S8nxF/CfGC1HJG1echEqU/zBSySdYKO6JD1diJNaLL
xUJmeb5c1glTcN7l/ANy1cYnOMGGulAuMOHs9jDiQElsciwUNDF1KAEDZkIpRAsIA7sCGyzGbcrH
rWrhD2rksiXdtIKKm1Buc7O38VeMl8w33eOQj7V6GfaxJSHbjQN6vv4IeWIlLS9NoaNrn1QZxHJY
ACYSF+3jmkJxG5W8YRbgkTC1QHpEFrPCPQz89McpWwpDNByimr19zSzpzKPJbMvW4gjhtKIDFdBT
cOPhQg0bmkusOEy0MOFs+6Z9+fK9WS347/qTkOCvlRDM+H/+iPTSXtQpgKgk/Ej+4BSPePW0n6ab
Clyv6HVXK0T+sqJewpIrrtWrNeFx2Z2zPivD24uv83z/3EnXmdNj4H9O/d5yp56JgdpxwNaMw4oU
FTTJLjxGZoH3/At6jm7YEFOFrc67Sk9DezwNd8lebje62eaAq3LjRC6UhYZmcluybBhjhsx4qi2/
Dy7AATNDiEeT4awLsx2FkhlGh2s2BiCxSheam4YdwHlN5YAZXzmFhPbHcS1PEHXOWzGAkazYKr12
d3Ij5u9j+b83DMnZIgJrAqXJeGFhs7RK2H4yFYS46i5zXnEesAJ3tUfrvrKRLm71l0Ul7jRxXnZG
8TGCf8Xt18LsF81RERZ5dTcQBzAFC1Gy4SnYNWeYCT2VoSGBNFsyUj1+WA1ZCgl0MyftazMIPvkX
aAgj/WucSLaphD1RQluIER0ETM0X3uHl1G7qgN8E4cSa8aSIuNgv1hzEHrEV2qQUa2QKY7wbqJvF
FcIj78VGgvtPwmsaUOc5m6m2JMl5VcY5y0o2uLlVsKm8T9TMS8GK1cX6AAL0IeQYd2L82HKzkUXf
yNC3c+vLAFZzB2yinBeOaB8rXnUuP3PgeM1ia7hdOV///uYYZk3SyoWuIua+cEJ4K94Pco6yGNj2
qlZ33fk/1/G95YoWwqaWBXSGoddRUSHULgPl5mO3vqG39ZTQb5YsquvYCktspC96gqeReTrgIqUB
aXkFRBPbUjfzzI/DOhgtOGZR9R9zXuZmUaPK2BvCkLUuGkdPj1I/UbPZvW/KSIcnTyFOPc5r/2vN
jXJK7S4vJg6UQ2wacwViBHAl18UgiTamu062yw0gEXZIPMMAASdOPqRW+c31tVs4ZjbpDfrYYrO7
bLGqNQNLuXkeSSfBio8xGM0cBJ72qdr+N4gumXnlPIBpnsozim4ONGw2W9oVk3pEZ9FWRrTvXofk
VESN+m33E1tEw7b0PiPEFTDZyCyk9ShpzBMY45u4VdimLPVibxn0XpF4r/Q6vMgDkgXPEsQcjBef
b9S+rTxf7t8F7IIYlAQ3lDQLwFAe/q42RBCs/sj2rU/ZQiZyVrwIe1yX1Sc0Wr4nR6A7fE6OOVYQ
VoOFQCI0wlYgeRM3ibgGuU1JWVsUqe5v+22bv5VHlw1GjiNV6qikQl1JBorOuXlDEXVD9nbAP5KL
o1ZE14XLVRY11k8Bw4PIRQf7Hgsj7+WygkoqJwvVi0m1fh91K3Z5iEkTLk8DNOKHBdWFegZjAKlo
vFOcylHaWjzgo3HSp9axoxyt/ZRSRuY9yzkcWeNVwBSn8hpOkoJ37FvMFntF31yQaRe051K9L0DG
EHSgNMlDMbWEB9FYLrVX6EDIDOZCZld0K+tDGW+OfqdVtq3KVqtmTfFfC2+5glNHR5XGwVD4Tb9K
pBrXk3PXILUkHms9jw4SXt6Mk6uDaaYKD9iQvhfxnRA8ULWO9lTue4tJP/WVr1xdxbSGYYb/V7TC
scQUcmE6wEjlNAal3jDDV37Febk1zgDiMg3EspkWgVJ2T/zJcwUfSy94nV8oj0deoGCt+5B8iOcS
9yUcxF011PMpaJK10kyVPRk/1ALQZ4wRLFuHxdQCwvb4IBmenF/VrxIeTa0jb4hxT3J0EZ0fhlE8
Wh+hZAsSi10JbcWA0ifNQyaWsRWeTc6cVrZP/rruxQn0jJAJwXeLo8QBOCqNuW/gZLxUEK6JSG6o
zgKkh275u6miO/uD1AEySe3XgS4rntsmxUDKpvPQHiJWJX0SfYhsp5c2eRIYQwaMYez+YHQjnYFd
4cFVuTVz9ILSh+VwXdEf4Mm3UW3eSXxxhrQpy39d/7KescMYnSFKgf3prMmGxP6N/9kh8XN8NQ1K
eWCewCmVsENNwWA6pmmW21YoIgRRTbD03RNQ3q6NptX2Q+3J0QXZ1ps5Zj2k5C1DCEN+/Jjiu5C9
J5DfvSLDfmvXEjSEaTVAyQkBMj1o7F6+py/XtOujiTT1u9+Xq0SBBeSMsBAioxSUIf4FtT8ksRkm
ajLe0Yzv0udb7Dqg/rKSXM6Rvvi+LCDlYLyktVdPUbe1aSmAMJEqRBe8CtRbF8bF/kbhdCy7NOOX
XHY68VFCDszoUK50kHDroyNpQwCxFjn0zVD3ZGvgmauhJTV4t71Oh5arz/l4MvRrjajhuV2wDFL5
IzUX9A0t1MWMQFj8aCNbGmEHtLbbpSSjuNWAeG/QqfGRXhUwhN9H7WrATOXRJVVPEqyoG4M1VwQk
XTmHeaBKyxXZNCPP+u01fUEm0jbRWDKo0zkU6Wi7amdLo2nvzh6TRK1TlEoOgm5TW/vxhZbHBy9o
tp0DCbBQ1B50YYc41wc4Lwflah9MXFZ1osAmAI+g9Xxm61nd+YfIO21Bmn83B89y02a8xp7MQFsu
OR8fevXCtNQTSZQ8SqNEHuD5ffmhDRFfPRpQQfcTBc/CAQYPXuYGZ3A+HPrmIwAovd9fZBjLWTff
Uldk1Rd0yujfQ0L1k9Lz8XhPRI+wjLf/jXPNO40kynxdJqkIFdDRkANVMGEMFqkY9C1ji7w9f6Bq
o6PQGgJAndNH3GxV526/LdNc8wCdULWCm49xWk/3ghSG0LjWtflzpuBPUAgxhSjfT6ISwTYED8el
enugXg1TlkXj0RS/XpQTF3WekMZY6etJjYDozwy1aKSastB2b+FgRQDe+NNjd+w37/Ky7CsUyFq4
mSPeyLezlxRx/fTcVQGUCJQNQmS032NDlxtFVdFkTMZRGjVFinIAyylj78d20mm6EWnhYc59Wnfr
jASMFlFIsrbojmhVEZIq8hAcHwb3EdIP/OC1gT4i2OHl2MoGhPFXq5V91xkbrYkPqwEcLc/qdL7T
4OL6fdbVmFlyoJU2Yz01j2e57XLYB7IHgztzWydgHUfJwhNMWCL0oW1POzwbj+2HSQRkNO9NeE59
EL+BZMzFZ/iVZhEqfSlD9jLithHNcS4q3CYRKt0GRfD7e5PUBi995RUZmN5eVqdVJmq7Xi7IV6um
pBC6vqTEemISf+l5cnDCDen7QsxKmXQo6Wpu0Ezb5ZwxHA7T/7nsBjmfYhD5iA1JGPqs1yPLwEms
VSY9Y6HliNIaCf2egy+NdrMZd7yMBZzCBS2nwYTbr/U/TqGL+whO1vW86Xm6Md6owTcOwf2FqgHD
KJ0MfiA6DGQf9mAX1arjyAyK9Kvb/G15yd6pEoxasPIWy0ytU6OSyJoMHKrlaU90see2hBZ/NcpU
fLXkajODZM4u2w4x1JceLaaoPBcLc2iQljzgbsZPHclKD1KYsXIXsp1FjSOHAQdqhY5j1y8A304H
gaoMCN0jPl5zqEudUOnhzosBbgVwF6ygRpONTvRUzDNIIQQrDzgfRtG2J3z4ygLE9nBerH6I8VTD
msaTeYInNrAn8JxelSntSuP5CVnOpk42X8kbaYWLwu1dSKo1QQAhvytzp2T4jalIdABlJKctRqEi
9UAyWGeauqEDL+pBslrU3J0hHeznZJrovd1MYks3IMdYQosLEMOXrQMdMzIiYy5nPFN0xczPG73z
/eaHQZCyGOSmG/dVk2r4dvdtboGmVqEJu2jGwYZy7gBss2gejZ9iLmM9PdynbLIBnDeZq6ziIB2b
3rcNe1EIT+EdsS6+03BkO48AAQrCNKnjhczaqWYpmyY4qlew2PcEOj2iGbGCP0MZf2HMRsjg9SR8
cIuihpcs46epYNWsqWVojHMYwEzfGF1mz7yG6cY5V6ZyqHGTLM5a5uiadLHmpm7k9kYz3qiV+t2+
6HHa4XtT2oRXvHexYdZaK4/gqOy8g4zJfSGYRsXey2xmEN8CW2wgCmoKsxzYPPVunxGvuu3hpmfP
R6OyAXhOaBlNUspgh/BvKM6c3HlB+bGfQ48TbXc0y+XP3JR1qUCzahlrHhWw5g0+mIhnfPQpiSaq
aOrxO6BX2kCFgktS7vN0vQgdLVuXg0gvPtQKtCUQGqbztBXXSsWKv03C6G/JMWSERrSKARjD5VH1
Ro+EdmehTiFZamt9XIcDk5OEPR65lxNXLLQSw6jV8so8y87UMAc12S6vbE4HEmWke20fh075SvdA
vFPCQUqyKHfMQS9nsxEI1ACgrdxs6gB5THVPc3Srzs1mH0g8nWxAZImyBC9J7/aeO1kF/gMIaYLR
2LiTpwr3YhqnrQIUhs2pL6/QLvVp4UJdKPKgeQX+5ty7GEZPFjPwhFOF7i8FP96ovgyzWxSq73kN
f08xi8+lkWxIhjPR8YtHTBI68/cpcWA39oiArzXx0E727GO0wj2WSXZq33ZZY7+kQytLIrkLBlIF
9rqxjTS5MATjffuYhN9psCPqLl6UdBWrD4g8fXZ5Mo2RkcTWl/NaTIDX+66rGfbgLKkgR9veJgqW
KWZhlsJL/x7FdUNggqYBYiKa9/HN/B3NBQFzehlO1yLA9+MPXirDulY/eNwFXeCdAdL3kmk+j5Lo
h9cjElltbcDRqhYPubUPiSLpv8qx6ZSk/5fkqHqaUe0y+w69xmccM42zxSA/QjcHbKokvkRU1ohD
2tj5nDabE7Vvbo/d40ZQ1fW1d7nHZvtf0cQND9XcqJITn+GrX0BGeeZYwHRSS02BvsTq20dHZ2B2
ME2RNHT9rMsAiMMv7I63On+zfUZ/jxIcESFq67MHEU3ZK3ota0rN2odTahEUy/1M4QLJzxP3IzUc
WAUyO0M94qcqO55h5xtCZ5K6xwgj3HcYVJ9LJPPGez0OUmyhoQ3gzORYlbYHLbTgCLXLxcR8I+O6
wAac589EIlSAMlBkPVzhSjUDC4knYjWaFgg50xnscBiPAI6aNZjEmKYeyCqP5kVZPjg1XQB+NOyi
E/gsFiWECPpcAq4TZpcZudZyy/qnF/0GwmWnwrz16bI7BnmpJ/HmRjMch9115VZblGkbIK0Bq4aK
bIeIvc6kx+yQt9ASTHL6ijGF163Lo5YBE5wA7ws8qtfJ7vca98Bgi7CcNwmlr1/l+hCs/N/IRoCq
O/Kk5T6WCFW59Jr1Ywv3BuOvtNRMyWX4hx7rIXLQhwGJzUh5LNWBHDy11V5Asld3ws54DPTRfsiw
uciwkb7JX7tKuldESXtp7kKb5D4nvKZeS/KD26VwSPY+2BJBD3ggw0aYrdwdIt2xrQ7Pie1LB2UD
XZpkdAM2YRu21Ag/Qp1zBRWfDqTJX6r1ls0Z96Bbczn2b8rPTTIS++vbFIerlv95a2QxOODuhNKT
JfTlSAXO5ynveKYx3/MScXJm2k3cm30gi0i7XYdMsKWpI/pqIYGhAv8jra9lFDPXjDPFGUxoxKDs
JtuCpUXEqwTF/l9GW9Pq+QtENTjlvm61w2fRQpHw4u/m86YIkmq+Q0/5Kj589z6FPvkFO+JVZus7
AMIcFBrmSKCNyzk39C6QQxa34eHBxNeLtBML9J52yIfQoUMCHUT/7PMId6+E78eEjqZZhYxzC8My
YzYnaH3E9YkxTE+Z0GYEiTkFLJnMwOtqeIZSpq5s9N/suo4xNxRlICurbYGxD6ioTI28x+frPwCY
jra9QC27YmaREZCtIsX/3pz74SUrPNeV6HMBqWQrMlMpCzgI70XD9xasYOpGSA7MjzPe7OEw7gP0
4in/eZPIfRMDdA8fq0LSdbtN3SIkL6W8koiDIBTOhuBymHaRxca9fhgSPtZD0rRcLvz7GZ8YozZl
RcFRptZvmZPjiYYGsVZjUjhvvWKKB5SIuDb952oy8jdyehSyBH6Rlk/Hz5yE0zDB3pgdw3yHDBSB
YwV98Xx4a9DoL2TtfFx97X+yU/fZ08Ou4VnVJLhUWkpVr4Zop2XADVraXYNFPxMhHKA2gpXixErG
bElaEoo2Ewy9pTsrp7iWIOvat09zZknUHd+iZPblsgZ0H0KNCalAPsTWXmM/sUW01LFcrgzVgnrQ
DyFoBZQbpzYK1Fo4T9QRmFNiiYqwFG/jWOUEneuh0vocZ/5Mf4kjqUJFPQL189XRThiBWrQXgFJp
DI7zmxSduQfAUEIrNUDefVuIwbBpA7KEMCHenMw/7uJYcO8LqFx9ERkFXjclC2y+zD+5/ijF5kj/
EoIiTAOvR4kSgG8jn+4pfU9pPC/uHFh6tqVp0ZPce2FBN9pqKCm2NI7l9xfy+dRCSfcIUjWptuDm
V6IH27yvnFmXV7Tg+vZHop2tuWR+dGJKWbJh7sxpWiVGlqxy6bKatlLXWjMS7cjDVkcKyztt3RXO
OrbCE8wshXdr5II+siPADQpLsXYw4SrI3iERywqsyJ/PLVtlorDwBzPGHXKddEWXK8yZBWok+kd3
JuTFULV5tKJhoFZJajn38pV6Z5AVR+x6B8WD3PGz6GDDQdjrzxTJ2zs7OtADwQhc/8Od6kWiD6GW
tJSku8T1xZXCGYbe/uExlHl1F7wKHEi+qPenEKyNP1iquycgcVr1LmQO4Ape/O6HP4Ev6GW8MxsI
76XUd6EAn2w7tx6pX/2GagIqYVc4TGJR5pEWXbdswBlraxsJ7K+rxa2N5Y1qhLwziTqet7JQUvJk
ndl20BvegYDxXqA21+GGvMWFB+7JRWVxvyYiCSOqwSr9g2M3+cHaBnHB0PpGMSI+3XK+OfEf3kvo
DzeL+2szBwjw8EBC9bMq1RLd6hMUZqoYtoxPBQDRgHmD4FFXoLellpxiNNxni+jj2lGMyps6b0P7
2U3+Va3uMgjmVOcorwDEMnKHZe/M8hNryFzQOAJV1C9VSM9ghR/a06VzztWU6l6YrzqcGW9u8rNH
ecO0L9FZnF6htX/iKXIVks5efbMoKGftYVe1TCyvz0wPaJcLo5wTOUOGIGBNIy3hH4lMNCNqlDXf
glcu6wnUIvWYLWz2Uf9JtAiIh0JqLiJmkRTSPy+o0Zihdv2c4NCFUjqwDJ8Zn47TnkvBEEn/UH20
Nmpn3a8q8Qra2c+6hapBJkH89DOqMrtOI/8QKYzQFdPgJdzqa1D6b/xhY3NT/dC740aQqL7Vggje
1Rw0o0q2DRzKm6s8fZ6I0VUwEsPM5DuuYvoAZaW5l6UlAA8ovxf6/owHB4cWUP0FnnYoLgo5j3Gh
tGsgOdWdb2yaDPtBihK2tedAcLgHZYZoDFVL+mOSquJeKOrqDrX3qhklVpGL8L52dp/G0xHVqjNh
1J3UOflk9Y2X9h33/qs+U6GanYehavgpCTG/6kjZt2TxVJCiCSBSSPy5C7WONewOvLPe0Y58uz9d
HrMRznskzbmCpEhqWjkANS0Hctoh6H6x7f+NCvk9K0JpDuMGN2/KHRhrYUOGR48dUbmIrurOL8FX
b8Pa7XgPUsNrnnbA0eIV0MD1rHjg+UsL0FB8dJu/dJrZbmIP7ozeFjs6zEVMb1Zsdv1ps/uRND+q
OoxgLnLxYkNL8LAS/Tj8JbCS67opBHPSaEbiJBrunF1iIluGUgtFJj8ebCSVarDIZMnAsKrF5QTA
cPLCo85E/i46ChrRfg9Ll6HfYxTWOjvGOpR4egG8rpGWy1QnRgZZEZ+IicX9SGTliLRxmMCB0RgD
lYfOe0veE62gcSNSH+8/95CTG9wg9fWKJTRUN/c5MDsoXOmikcgESa4mqRWc1fF8RIbIHRVIcy34
UvoWCKKydcW0fYepFd227dwrITxX7ROVedoSwlOc9oA3Bm37TbB0GI1HbZBZrfmWRBqWa3uay3qd
f8bve1kjQZukAqnlj9zrmKie8eAlcvrgZ18sMcek/1Vr7a+9Z5FifmheR0EL83P4MHmvefuDydfL
n527a5uSQBLhS+jLWLp8o+fmHmMZaCGcgkhIocTNsJgeS1SsNgEtWEaOKBsGkcgFfOi6mwp4AQYP
TLzSPKKpM3UyYn4Ew65fPaD3T6p3nvPr0byTgul3IfQXSD4R4H3nWWEu5NLW4mkGYFVreGS+Mwrk
9kwQsN3vwlD8H2+P4t+/ZQw/HOZ4k457ZNiZTuPEjosi+9zVH5VTnnnrvo2xs26M1o2aXA/z+7q8
8kC2rmCX+2qRQ4J9Pjd5T8oagbykHJQkaoClVrvnTSVJW4fPGyea761vpJHm76ssPQ4S3KkdmoaT
UcCmMjA5I9gVL3cww055yu9wWS+EUI6EUf081kvQYD2Hs3p/scWbRwrY4jurRXUtmI/dLp5Fk3sp
PiU1ZXATdm+zEfzRXXyzEm07y4iP+2n/VWhNTZujrF8fzhRd3tYs7JoPkPStvREsi/SxIK54U8LV
QgCC1w+9pmqJMzqUt7CaGbTWkedJ+w6zixlCh3vtfVaps/Tk/yd8carh8IUWM32u3vipjwAKYEp6
AQaoaNX5ufN5LJOlNPl7p3fTgt32Pb4ESWFcPS+EumP+UJLfS9aZLg2YCg6kZ1D3GV71bszG/NLI
fM5AF9oj++EuefzpJa7icm26ZCBEjAoje1NRXy+6KdqwWw13o5GD/SjfvqW0REZshGsRzmcJjFyr
3eu5eJWxFp4mg0kZ8EZcv4fBCNYHYTuDxnC7euZ6kBk517lNwQ1iEabewpjve9xt12OaO9kYMs6M
eI1cmf/d0ufBuGnrxGhpkksQM3uvjZ7JzkWiQRLsQMGq5Pv+VSqPVlt3fpvZHvGUJ2hqOqDq+X5U
/L87qB14eaKTfxNlVcxrJlVf/F5XLj5S5Gmet/xLmZm8aknl17Im/gTz0SrmjRujxFch/zS5D/Cj
kCzgwUzpkt3RBF14KtnTLdWFVSf5/egGXpvP17+4Y6o2q6fogD5ZMBoUM+rAV+B3HwiKxErtSC29
Yoiz2iKELMFEdUagOBryJQs1twVYpu/lCUmIT6ZJklPs/yQuEizFw2CtXjQW0au6Ofp4dAyJlQPP
xFRK6yE/gP4i/KbLM3hR2KwOqSmFgGoYtE94ZzUrUwqPCmF2CQgYOkO1LFvdQ5JmMv0zTuIaINZ7
LJNYG4KQvR3fWc1RJakRY5tBI/Of4/EiV1bM1e7B/tXYKq2MYaxk/ERv3eGx2Oga0SoECjvg4pHe
Yxb6YKcs6EGHsUpnBMaA1YRXM4YPDDz5svdQp6+GjBnmk78bUdgor/URm4SB4NYAJjnU/CONjLQi
jSowZRCiRC4ER3ZJEVNNKCXInujYLYwBKVVndjpNNIKe/XzQfOW5W0fK+5BaYf0S6CO74BK069zm
GP714VCAPMz5ukPDoNsypR0DbIltdFHSwDapCTFaORtpSPrzFJIO8ZfSZcJtWSs/jJ3tjtPPNiy5
sTCpTZqKZFIbDzVxq0H7FeCgKZkvLB3tnCJopn4CGpeQjpCtYY8dQHHE1/u93+hE/SkZwMTBfkxL
Xg6bIbCXnX0+8OZtlfizmhul5pZg9BsWilmlmJTZJEnUX08NaMUcAhWRJt4Ws3Go+GXvnvncZJLs
eyMfQ/Yzm483jrudYDt9fyeYzpeQc4x8fh4NaRuvVs5aLdPGE9fjYV2YvSgg/4O5zPJIQz4h5Nd9
0ISAsymP2Smly2xqY4ma+ja/UcC9qIbw3ZNCZ6eFDeM78OnXNwiHDXvvot73F89eZEVvOmoHqZZA
79lXcEdfRnJMDa5U2t4ur3zrRv0N5bdBXCoEP7tQLlajaP0xE1GBxKshB/6Ve+RIXShPjnxep5+O
kE6DAajGDsCkXH0k0CKGYFx9ykiRGbWucSDaclcD+yVTjcV1Z4itujiBkJlyMBfEHaGAtNHg40o6
yleatMFDa8YvACk+T2P+D543jDenpr2rkEp18Jo6whAmroJwO81hqasIOYffQ6szys3xKchhOezy
jcdLMDZrTuaFvD2zW9+9RtZIJiDUnIxd6nf/Hafy56Lh1CM4wUzUGGmVSNIhY3aG2QXSsxuEu6UT
unhYr72P3s6K7aVFFUDkCShzmQdQf41oeh+nmu8n4YsvjggirvbBmK8KnSp4LrhC3vCWdFdT8IHH
PXfWYBLNd1ikKMhMJ73LPd8K+assS4Im7aBryz6FjgvrzLRxmN+XWASu9N3SZpKA63iopnB8NnFP
g0WU+3ijCBQVQ1oAY1Snfz+OA73IHj/4/RMqvYm7vJ7E5bCDTv4SkQMGE4DfpmWYFOQ8RkrR+gDH
Qak2Rvz6a9VPJ3btw5ICCmH+UOnN3pOG07GMh/pD2YpNcWFHF/ku0yTGkPacgi8ldzm5Qk6cDEXl
HSiiFOLuTW65qaADFcAghzkpP7us7ftW7XRwCtT/T0oIEoIIN2CwPvv9h+wkrVYLCLWFPOb+2pnC
DJwIqjZag5ojJG0L7MYN83miEqcfnRkclaQ/YtzPv/bOkhn8jZcd+KbQVp+Ua7XaQcrv5k7id3w8
znwvOOjb2/tDyRve5IE7QC9dVl/+YiQj2HlO7b+M1bRBNy40MJQphk6yHv02D4mKtvipv9PmrquS
jsX39a7tUZUrM6Ld014wZZKKPoONNgy0SAyNYPO787DW0cfdYt1eDnjlzxLb2pAYBmI9md/ZpvVp
lwgNzKHhuhndqH9Ob9Gn/AFXBwalcBvI7cGppw4e0C1a+1+cz0IF2LrpoGv8nU9egf0TE1hUfLFn
wCs8b1wgEarA8fKebDvGAQOKqe+Wt3UxpmYvAWKaWIly3v6+qBGbJOHqATot/b4826Jr24mZY5M7
9X28VOA8f0GHP1ZcGvUDpUXw4Hi9jINYiuVTPmM9JjmtGex9yuUHXKqQWP0d5FUDr9AJ6tSMv3ip
Kjd3BZV7/9yruryLYgUUUGmhjGx9DTkHZl9VePI2Kho5MpqUbmAcCH/6crS3VFj4V0/r+TIumaOp
8OO7wBwRRjOgppUdcgTmSw7zxcM9EcnNde10/AZ9IZ3qtVenh0C+qjj2/0VGbTJjLz3KTYpBLsC2
CawMeHMPYZHlbuN64OHw8MxN1b4X+wJzb4gLpYH7MvmDnOXPfsF5gumuVfKXl1XRgFFJp4ZOuxXQ
tafPGDUsy3kW6+s1gc+Pk/tDPFlVaBCtzT29hrUqwAyW0KCuxbhWZZ134DMjddjuEMRR9C8b/Rvh
8Aj/u7JL1u/FpB/OCoL0jHGcHA6jH1lklVXloDAg1e8vToESQw1pIBDMQUFOaOskjFUclantliAF
/zhNrlmKN2vngFfyCJFa2moVBtkAudl8wWOQbjTSOHsDYAlgoIzy5cuLdQy0OUVmv52h0mkj5z6L
JBKHPSKjc3gK4oHxBOzAhluozERkPebIWcntbEOFmaIpScNXwnI8UDJzvcUqTKfeg0aDOAU/Cs8O
v3huiNBv2NeO9VaAiKetHHh+cOkLQHYS2hoo4HFSrj7L4m+StZEILYmCd26TLq8YZhddU3lfDbgf
aa4px8U3kEdg70dXkA2doeoc3UcSAC2hPbiOKSE2bbRooCPP2J39xrR9VTDVrgNO9Oz8Kvtad44i
zBCSFnUckDLyj+2gO7Bk/jxEEM7FlxfE3SupDElgfgJw8bzLfLkeNEfZmNd+DM/hyhy8qL2jk/Hz
HlJoKaqOH0Xn1PVbAl2e1SINN/E3QCFniocqrZXuOWmVrH9xiYGRUIPMwXb9e+4m+uR06YXfLdpq
RYuugW2TKdr5MvHy3Nhj9VSa1J1r2weRjHcbciV5I+IZen4JVGjH5d/negrVArbNxv1mgD9ZzpVC
rBs5e9OoftUY5tAlLvz7CCKUuPaeHJWwT10LdJ7MY6PoOpjk1pZVaxqS3mbWX3jRipkKTbGkmFSe
ZntnjpCC9o+HSceMUH1mrYmPdr2CgzI7crxUlbUEzFEAK1nSx+RAEEbNxy4LwisoYdDWRsD4AYZq
K3LeHGi1QZtLXUWi0rzqpA8jVdM//Oq86t7Bc0G0pSY7w6xi24qZKYsYfykjelInyple1JPWF6ll
0uRo1dLhbD2mZFLXWmUrSCZll7FOrClrUX3Emf5Hg+SyLoghLE92nEH+tIhdD3POyL3O9iM6k04i
xiW7hThhcNz/IEBlurNkSdtSSxlWu2OYONi5K/vy0hN6qwihIXGBV6Arm54pagk2rxmpkBW4+i9X
xt0p7kxy3Dsg7a/Pk3b1IsnvvzfUwrd/jTR76TmofwRFrixUf8BLdC4/Nakt7BHKf/WKoVteQWV9
7ykxyj9pvZdo5xJQ8ScSIhB7JhSWN0cZuEkKElVP35hWjIA8RRF9soel9WkZ8cksRhsSUwN4aIrA
EN0Z3IPrB3npwNExvsHY0ZkJA8iNTVM/HUKjSYC8VvUHeJCMobMrtSZQxoNedlozkbpOqWX2+DC5
5YVjGYFgPlHK4hrCdufQGXFIAN+BHaB/4gFPIx8i+s2g6jscdQw3URzaOIZT1aj1wepOLmrWw/vW
HADPt5OmuHh32CRGpfGGqLNYP+EiNupMKsQpyLLPbP9qObn3HMCM4vzLRCeL4qrIZElusG0OJ8XK
CGYNdxPpcolMfXLBqibkFZ6M5QAoUKDp/sfY4hipFTcS1BA2W7GmSf2Z+j06Oio8lyOzZTmlhgMS
RWAYVeV5b7QdtXPB7Kbebsq9S+rBCpmvhkWv1nEVDQTOvcH9gAfINDNw7T0ylTOSAV1pJ6sranNb
1fkBAoshUOiLgbFOKLz+9UF20aMseFUIPBM5bBg6bzBaDWc5DTQS7NIPlq2RcrUb2P+ilZVhEJys
23CTnimoVoGYZrKVE4YrLHV15EmvFoGzt1bn1qrEM/CARvU7sH94F31WCaknWMYzaJ4oGtx9qi+0
G2fA0ICfct48pGl/24zfNvid5tOFivoVlNhRkND8uY1z5Ql38L0zwZw4QSgEKr8/zk8AmKYcjSrV
i9MMHtS3FeCtNECDqzpQbAf+EMqJZj2KRGxiHov8i4/utBibXlM2agCm9O3mMEBQkVtoj1wdzIAh
GrUYeEZZISU+8z8xbIn/pY/nFLcIlGpvsJTleRtE0sLlByDFBtFLYb8F7o7lCoCOke4Y63QWwHuf
G+ejJM+06J9S91AskGywRDkXokLMiiV0K3t6k/qcMTxnRbeRRW1xLswVGe1bShDmIHjC27zlRXhp
KFc1gI8U1g5qD+RTaLhBQ/QLxX8JUKwX2VGv1PnNfIE+tEKIBsilAo3WuPhgXFKCb/+5a+IQsV5W
SuLTSU2P1GeLKCYlE6h066Q2gaJGuU5zl2Io7HPxxB71x8YqEcDwCKIIM5vH8rMGaodvglp6oTSg
Qdk1+MjQ7yYsytFGNx4/76Ix4jSW8CyLF60AcYRN6VR3zr+jnOgA1QU3J3r8Vut4evvNKJ+c+uXd
pV8BsH1oYr5E/Yfe6yg4yUNCh6jJkvxjFeonsPMcpsjUu8Ptz8JiCSNo1Du0K+SCWbq6EPlBd8Do
lFTUJ0535pcOI3g8X2sGbIb9KhmiIE/jbGDu4sybDAT56k1ItmkQezUs47chsQmuWiMcsM3AU6MC
FnQoGKnUFdmnHfi9D4CdmUy83wwoZsPx8mKaaoqLmT+kL++0dvsdlZyDiUheP9i2fMLhD0tS7JK0
9VGtWQpzL86KI2rvXhZEd4y0PDuuwheMNFsiku+pauyKd1gBpJNPThCIyaiihqrFewAGbCVyY9Cb
fYkGD6INScINQxy99A3Tox6O/ixBdCXeNjJWEF/s7deDTDicLPyaIWmMdX+Yo6KzzTVzh3h89g37
mElDpgCEM005dL5L72ds4HNzUqEoRtZVnkcIOIDQgy8tfNPiUdnJbCvbm8uigQuop+0teS+yDGmY
KT4VXeQ37H2Ry4glCSdPSMS28FHE2yCiKt3LesCfRr8Fqxrhhjz570ge5yu0Mcuisxdr32V2pWQj
rzrr6mLDpIngwzM2a64cIkaClPlPwjeZ11vbpdE4xNr6R7yXGWm2REOXbeTwnoJcWG05/Vj850xx
V3QCC1PLexHnfl2e0g4Kn34iH/4ws5n/SkZ04QZMYjQRqM73S7e+VtVrYEPJKmLDXR8Rr8B9zjVC
1D+acugE9Gr5HAphDOg6V0BlKcz2MYHPB9xNuxehqoVJ8pndYUL/nju4gv0LpgHBUaCmhN8hld4x
MSbf/eXg/u1rwBWN2pGFv5Pm8I68ZCFX/adfOO4LuNaNcivRL+dLmuDuGCDKOLcBtEZt5V0AHxvO
+A2vrpdnrEhEoOljKbta1RfdGYhnWSxQ3I52Yl4RbUmWD3Nz6aF4sGrBUpGYNkzGcXrr+1xUKMti
Rs42opE4JQ+5fhxTM9k8BPkjUqjRjX3nzFuOdiUYY9SgpHv2GnbSiM8C71cAJZJXMd7atCzWw31e
cIypMcn7dav/QQZJ9hJexd6ncVc4QNss3rWZzg7+GpNB2mxeL+eORJfjeZPmSQV9ikJRcILfYc1Z
l4Rdp/iAm22NC06RSYBvRI47E84OgEUsVGtFmGqCroCyu8VrNAak3RDchhbnCVNCssohst8Na7SC
PFxaKQaAAkHXOHVr28+YoL859G3DnT5Y+RwNVsAJ3QS3UVJ2T/p2y2TGDlM9T/s2mm4Qh0wzykLd
7t4QcBQCZyA6JKx72N/x/7PW0On6tK1xWgVSOumxl1Km51LyU3MlAZ3x7m/qSrrsBU+mH7DZ36jB
IBMd6V+L58gSmwGNV5yOe89E+LHc+8i2GiFrBxFGjypvlIfZlDqCG3vNY9IkgzATsY1sh3h/9UuG
wtKBp7th1SEH8B2IHlHGYZQxqsMur42BjcbE9z2Mnim+xrh0NfmVKRAOGPTtRYtXP7t+S3m6fd1t
H50/Mb+u+Ol1/AtviVPCyfSE6tArFoj70RtVCojV0y9JCJuebZtM944MsVCRmqnUv5w+O5pbzZO1
FAfv1k/imNT9GmkkQbj4Vedl+ycd/wMZJzGYOCq2wAwGAHKGcged+IB8Nn0fohrJjcBiG8pruygQ
+nqM2l46GYqq0UlCH6IAj7xlJ2t7bHc33lWRKPH46utxVsb3xzcuYTmPbw5XwjF6U7pHxvmVGidf
2dJFeZJIORMD3s6cxNm7bfoWjX5gQxjl5gS5uERjiJl4qJVAps/P9sN8hTckL1l5ZRgPtXv9rlRo
WGleWtkmD/IEyzBc8y+Lchi7thGeJQeDLgyvi2FPqXj9eLyTTw6SaFHN2eUdKWtgnAR++NuRIAuz
Uu5Md285kDQhUx8zLv5ThtT2pTyI6FW/j0PySF07wLvndbZrP70a27EpBc2AMecDmkk4tbF9dSz8
06aa10hRptMNTx2n6n69mKb0GV4hHptJ3IXUuJF5MLz/MgSYtd4GLYbRfnR+nzHKNdgfvrNB0jSm
hR6hOfBmA+f6+Vy3NFIe2nSOUVPN+u4NPeduYBRs24ruxm5L2tFccEVSVUMZKR22+/SB6As8Y9pz
fVqJx3VwQ2fHQcBun/G0skGipFqXS6qflzCVCrcdCQoefczpEV+8vlov60Dku0QiXnruHX6xCEbb
9iR7Oun/TZiwqD08E2ixcE3PsSCsbR/RQpnWOIiphBur5+cRp4KHFm/rNYZikw/2ZuDm+wHVDGFD
MB3QuLTH3CWo832EFbXBiWDVHG8LZvlFBPQxfMr09Nmc0DInYL8Ld4tvY5T7uEFvxFpK60wJ7PUw
ncwXX+kxmgyGFe/jOqZMDS3Qyh50dYaqjxdmKSGCm4n4J9rgylBdyVpXWwgXSKcWSHFVmSFkfxNM
d4Hhq5jVbae6NaMmFkp1KUHIknoy+zIBgfZfMp0Ghu31h5IBHys1zlAOfPe1E01MsB/VI0rLC/jG
V/ZkA7D0rUGsLs6mdydVXrQEPC6ytYYRoBT3Silm3eGn1dXxSqL2BuMwXpVveatMzmhKiaoqZ8G5
iuy9h2QiG5FrUCsN1IOA/37dSIhNDxB7Enp/ZrnTF7nn7X1U/9I1UK+R7HhfDK6j74aEUAWQdfou
+f5gNFA3s9ebw2qkIhN/L+SQUOjShlTw6MLvf5Kde9/4/X4eAB/M/MIfQuJ/ee8tUqJVqP0WUUHf
8fTGLlZxMaxAl15XXThmgx2kFwHHn7J+iiIrjlCoOfcaFJwUywlN6TZVQg8t21zOU6DO/L/ry+gG
IkKJVhbiW7eC8endszpxjCo4JF8LhJjb7Ss78Xtk7y22x3FAAivEOxHMcyvXg8iwWSh3+5IrX0se
WftxFHsHC2ujBxnsafSgObDcexy5po0uW2EjwLt+1tf8PoCnBvaPTU6LB0Gasq4VY0rXQrN8/2EB
OKDSBQGN7t0sn8olO5g1tThqOeU5big6K1stIkFs/UG7Rqo/6L4KVjv+rM6mh0lMZANu42XSjwX4
1iFmoScX1wpbnolEWfo3cErlVY0gF59Acke0sRb0z7fWrbNGHcdz1tklewL5lq4hD5JGkJehqLCS
bi2Z9RtYqKJ59tlSITf363AU4u1H8buY/6PZAb97wWmtlsdv2fW9rH/f/AKPhwjuAlHuBHDGYixL
FiS17SXRO5JWAkfPvsISSQxKDCTdVcc+PB4V4OelY8+N++VYou33yoAGXx77qNqy1Wuo20SozAIb
nxlcey2Lsh8HFtl3UOOPl0C6GG40edmd3v0UDJflJNe4BGv4jw3rqwm8InYmC4uclVAlGr3jxxXk
DUm3eHxTJqV/sOkz2mFhQXaae+z8r5HjGfCZjLuGjZ3UXRTNIJbewj1/Ql0sbxBeXvpUawHFZsyW
X4JGg5eZ/6t1zQzv/eaUkiFnk/sq2L6cNarU7Hkcx2cz1hlMkLfWon4QSAVBlTacmA9ioSwNS6RO
/7im+RGTg1G6xgAf9EQr0Y6+G66DQLSSEyR32sYOBCnW8m0YIFdpfd1HLS/C4d49GvaFazf08z1a
izR/MJ3qK4qcI542WuDxLz+eLM7z1wZVS1d30uIo9EzrwfiARSevnDL60vGSh7Kw9aeQoFEKE0+S
d9ouYZKwCBW1U6lT+k2Q1SFmNtS+0Oer4Zyv6xocVkBcsMxPRmlZFMOSWn2f08ATSQNjF0h8vYln
dN37mRC/3elAL5+zObqjCnVekb8JZ/KtWDLXaUDnb8WD55WB3AbP+AHSUPrN9RtN5QSqxU/e41s5
V6oxskiXmhh9Y6ZpRK6fkcR9IIgxfun1nHRaoEI0Xhma8IR8wtGQHTFalvwOUE5UEKaX+MzYzVlv
iH074uXW8CDhnAKs1PYWqXPNx7PA4W9+8CMMM07Us6zWwK6Uel+aXa8vSJGHDcMtUiL/6jnb8GpW
m/M3HJ2WlrJfgIWq2FDna7Iw+wwhyL6vyULsrNIc1oMr84ae7sqQAPBl9bGKSbwQkxoekVgPH8T0
JHfwTlezwo+NzoyVS7e1DfWD+Rj7Ko9lyyJcAqtAUkeN7vDhMuM2uPJH3wD2TsYlwcg6qIOmlYcB
ozCq8phwKfg7MDT3UCbhEHcJBEOg4bEzzB04R1NwrC8sbHMcB0dCKCEKl71vjs4bAv9vu0t3yvzy
/a6/JS9yR/NyDoIDQFWLdHtS0c+b6Wte0iqLiUvQZijPChHHEBQJIf29/n8MVL6XiRVHEgQznzHQ
OY8lzZSKuGt224+aSXkBMSbZjG2+PI2OT7MiTkK76nG5fxPqzKe0GiyA33ODXfkZe/LqmH5Zh9KL
QIT+IgUQ5GlDTtXyVIbQVZKHRi4hxxGktzHi0R4U6Y1FvBEtSGLt6QIA4BkMbtIPbJ3rZ8KJBmFi
e8RLP+0+v0OO9b8fAXnb8oqv2Dr0pi5PYOlTHxaQVKm7ulKoEugLEVmOJiK3iq76Yi2SBKlqycgh
u7MxvyoXoJd0CoGpMjUefsHwwDXyElal7+HmugBllbF8OWn12AVzDYsSgWsPKxoJ5FrcPdVE8g32
gMh1wfOXSkalAJWWn7hJD555FavoRZ/DE4zEQH9nyzVn4XSCMMNjB9wjhbVe2D2tKu6dUL588kvR
X0cX/jK6zAP5wVbg4wOTAikzKYaOjgtBUmWR6i6m1FKZDRN9zoN/xdGYJvyUY/eTQ/cI8M/29buT
dIhznYvzDT2CDq0Uaj5Ld/hZ5StTeDJiewbmzl1+6QU6A4RidiymKvQMqEdO6cPM1boxEWkKJ8Z0
Mx+GfC9+lXTwnj6EW8M7fLWpIvUIJlGmf+Yh9msLqoH3d/RVBt8E1ludLWgQg+78Af78vzvMO4L/
zsrHQbk3+/Oelbcc533x0gsz2P96NjlaITomzJKizLeasOkmJBOe1gubWrX/VLNK5vVVz0dQcU6Y
vDNbzt/2cpjOpfl6ka2PWDpqzd5sSnHZy0PVy9AFO+pCbLIJ1nmexOn0WqZ3TZ8aOmi5OXfPzh/0
ylo+onMKMO61BrrN2PbuFusYBhzUnw4Ev0zeWogmFXCjvKCcoKRy2wm6C/b+qd4keGh2w6pxxPZu
3RprZEqqaYbk1Bok8omZToLcA8E0vKBXdwLd3aA9unTJUv3G9zbxr9o+ly3IrWLCeYOhKgu1JaUI
5wL4fLpQHxltF1jhn4O+ZhIBko+NEvs+Xh1gL3Uc6nSMrVYnIIa/cNIKaPBQF+CEsAyqcRB4XsmA
jFinNbte+BYmQaleCb7O77RrqvwA94TyDLUJd3q37vngiTMBnvW35lCuOFRIGKwdriS3YanUW3RI
zYty6Z8BPbVxmzPu9WmIMh5XigtIr1Dhh+UGNwKkQwlJ5O+RrMY2Sh/U4uhxTmy4liFsmTnTtS8h
3/b2nef48UHMxwBVaBqmYgRH0o0XnPFOR7J/AJ1MMh/W1doppy7Sq/TdxsDTUawJkNtqdtpQ6IHu
32EPMoB1Qg7GqqV+5Zts34ctyL8Pt3ae0/Gn9RBzPoCLtomJFuWZR8JcTxE7v1/wUjXPfxhSVib5
ADt5mjXp5n4cTXekVPYFdPw+NoxlCVF/rt6F4HAdua1VXslyWvwrlFVX82xZNKhtsmp4afMcDh2Q
YwJhz4P865UbWZSsE8i+k8ciAZNYKfZtWBWqafWciIf6y49bx8vhg19/9WOL6+HF77AGYTHZxT8g
asSUeNBxcdUr8jI8h5wJJEm+9XXzTedrk0S3O9Gr8Gu8e6eO96mcD4ztMGs0RJAnplBxxf+405mw
KUjFDKgZFI9wkz2V5rOoyD7ClU99/WTR5oXKjlEBxk1yXcvMKG1vn8YObWjDCzlFl6x1wa3dwtva
Y6W0nR5k/oAD4b9JzR04w7OUy76jdHsxsw+6U4r0HGGRPlzsFGJemSjlQ1K19scrfY7zePpsJkpj
Va0GyGiMKK9Jr2XrKOiIXnh/ZvMv3Zebx0u7DZiVKcij94gg1AXFCIB0ZpI5dEmjFfBtqfvaSe73
iC3VBgvtWoblugauYqR4YXZ1Mh02tl1QSNz2R14qxpTyqnV0hqk5WIsh2F0DYWkUPOEr1Ef00QLi
kovJBTt9eea+XduRgBidxpRS4gOig5CvIE+5vwUlw4ailZu/lDZAcDP/sQBSPf1N7Xz15Q8E3Y9X
kDOJsLI5kJ98WMw3CWmi2pwGODaAe+YfW7oLbgShH9hD2OIcoKfDCTUh7xB5Anf9/ZI2CMxDAuA4
2elmEmrMdoYy2Phcdt0pwkRDO0Rhq2Pef0AiYVmM1M550EZdytM2xWuQTcj/kyCxeFvGDaYMUTj8
qmPC1pJ6D1XjVZb4B8FgjPLl4SshglMoV5qaQ+Q+W+YSAVXkgYVFSsMs9rjEfbsv3oeOMnF0N4Zc
3OeO8EV/59nE+npsSOXbVpmQSufgnLgi4FKOUxYahDGlDCKdOxcDX2Ajp2rQSI24pI+m9av359+x
g7abSV657WxoyKavO2jGAXpThmwBCyXgaOsokRPySwIa+G/AurH1iKswMGg2UF3M3yCXyCF6A2O3
3dBi+FwlmjXOjDBra6NBy7OnMOzqG4F6gS45YLTYdyY8ScRgT1s8FnCEfH604RstkLev/1aoDX5H
k9T7euNvDutl2mUR1LP+dCdTQqgm3gVsPIxqobbF8t3TOUmVdf9H16tMe6GJH8vMT0jF1+jJUFU5
pTDSz/PgQ6Cz0clGsscWC52TSTbzeWJmEfAJJCdqxQ0y/tLZ4olA48o3sye01OjMHsMZn/nSVFpX
gjRGu/P6wHeP0DhFNrAXEpGVaJJZG1XBjLAfOEbBj0rRcgF+lhJWGIlsHGQFd5rbVkqaxJvq3Sos
6txGbJoyLrpgI23WT2/K8Tc1z2wb5xOU360Bp1AlEn5FNQIgbhrKQTXFxixEKLWDXJ9mFiqLm34g
tFDB4okLBCrgtEsGdQnSSjAaC88VKazfYdPsEK+2xxkMaXyYhokDxD231mbGHB1NMM2Zy7JewFpf
3u8rQXsQ4FMJnBKq0Ry2JFwufFho9+AlLrr46vWaE+0ExhknAh71LtSbO9E5ZEmPrCbc2WXojVnn
NqDlkXqRz1JJtov0XsQXvdoSKGDzUhJAYnNqD14THaMovJOsQwiGUM4hB/OqodoLUjSfuGTTXZuM
nY0yZ6Mg3EPfks2JGxq+wYTg5voEGTv+oRV6ydHBitHz7Ej+RmqKKhZtX9auy0DV6G2MnukkefdT
E5qJl3cV3eOIBrW6vdg2qNUZiX13C0Vj2EI5MCkCZF04xvvgqAgA3ne2CChXjaAM+ec4sSSxuUEL
gidKyng12rEVp1LAz6zZdPMLBH7x1sQBiccj1cV9fm9Wj20KSv/mo2V0lH5tY9ue7ufMZV0eOMl8
GdbKEkRYwpLHhfV+JnNJoe8g8XoHQbO289JR3/3Lev60UHA9tPdPf4IcIw9uZGFCuQILOIHQy79c
olUYx77f0+DKqdM9s1ot+3bRXqlc2U31bcUlBkXADqIHKth6rGcNurbrsdDqRe/OgW+vmB3euTqX
nztpKueWKNRyP12BNfRtaompfq9C54Xzwg4BSOFLW+axbg6qYiS/uo6cZNUvyKvPVyQuTbRRUVNZ
kFYSc7yj++kYpuXFYnTbaBYKxcNxvOfs2Ur3Br3oLrSuGMEtW/SxPi+FEOjYseVoJk65Tufelbid
2/0SoE2ZDAUSr1PlzNkbHu70mPai0mYQpFlz0UB/+oR2rhgn5JVmVXsv25oQowH/Q1VGRmIL5C1f
LKUJyyO017WnhA3GZP1k3PBX3Ax4EXTKLBAUrPEvj6dH+awwlfGiYXZKbEUjx7LweE14hwVQoS9L
cAPEs5by0FVCQZA+GTiybdwnAnIM7hwAlXfLwqngB7Jk7vmBBJZxBxOEFbJ0Bj+DvfH3hvyF1V6n
Yibl/DnS8/IGuBIlOBUdz99j49RUZPMw6cfEgx3iKGfLqX03G3Fsk3XO0JFr35Uu7pp1/e9gutdx
R5X5+eGCEYyNQ1urz3WeI+u6m9ZWwNiF+fBBLNaK+WRY4/uwwWqfuWFi7pLoq0hTFuhlUw1+z3+o
MZxsNq3MRn6wojpOPspkmWYFwaClUXBAKZM9ZTWQO0yvr+LwponYBg7lkAn4Lp2DoLZ/JqafyeDa
XZoTusAEBIBIbhoF+oqWOFPyNQhPTpkRH41mOZx2N5KDgADj/M14yX0dezjPSh9OUHigYf92fCGL
CWxfV8pb2DQycNN7tZ6rHxF3fcpGTlZZvm3UoGPSEpE7A08+2FlilNoXicWdcElQ+pK4CuV0eNNv
HMQ4P69C0KzUdJir7ytcASC5jmCvSCoaBMA9+VS9bW2oVWip1QxRZNUIuc25QflwYdlGSDwBVknU
vdB8bo2KB6rSrybT7croRlu82FAVibkL0OORhiN5kBkrkv6wDPbTQ0hZ2WzGICngOX+7nA2lxMGE
v9jf4Cv6TYmP61kG7Ivry+QglTgtN+5LkdwqwIKtWmK6Tk5qyKPw6XXPdUotq+2hEJqCJI007nVJ
xyIQvlWVrT9ncj5qk1Bdz9KCMcsrebwxMsnPb4VQkERYqaW4/UNkjZBDvEV90PEKScEjuuejdvZg
Eno9iyd3vmuWMxItN+42rCSdFQX7pdyHiznosYbCoZvhLuG5iFMP3/bZd8f1Z6lhxOiK3gXrwImb
cPJgxCKJT3iVSj8nIBw4k4wJbLRWmALkWLZ3Om1wPATaX5ziBwLtcn0b6WqBJgOON9pZhyDpZCMF
SnJOHZVQPB7Me+FoHqOWkEaF7Bt5DmpQo7onwtUYbt6KikNzLhUNRAX5o39OR2tEwNYXylHyov9h
5gbyLaee7KOLvGzdSmQ+AU52KMJwsjhfMxTIg84LizA5WoQItQ8cfzGwBcKibUc2jVwKH5Z/5oPK
eQBtfiCCe4ag/6is4UVJkCzabjW8inBmj0HsiuSPkCJXWN9vRkWpXPOkXSJ32Yt1YodWnAmje3zO
6M98vaoDQ17uaYRxjkmBEHoTbyKdM5Vk8Pe8+M0CXlmRV7/0DFa55MMM83ky+1GTsqZShKFbQTEu
cnaNNrfajo0g2IDR1NLJG1I250budbLUYVtg2l4BH6/W1WZv4XEMN6gyN6qCRi6A81JI8ONk+GfE
PA7mPWRuBLUySN2c+V7VPQaQb7hSHv0Q1zl0KkiVFd+kV4rsh2R7bHK4v4ISOV6QpIYXVckeEzRF
3Z+WukjUQKBkNsIde9CDdXHACE/c3kWiz2o/CNNCeVuy+Fh8wJidoMs9NniG1zDkasmswfWOEupw
5wqbowsB6JmK3pXpTruJcZIJT0g5mhXPZoUuyKSJtyK1Bow0NKvoUHwiaTN55iAq1q2Cn0Zdd2Eb
TdA1ChPdebVhQht8hxCUVP0S3ig4JN0FyP+8WSuYR5yOFlAC6upgHZ8gzFdka/y3Aqc+t0X67qQe
7X6NeuUMzE05z0at9gf+vOPF42aRu/mpokErw0DlRxRI2qpYbxea+LeQ0e6vLw4CUdandEufoJuU
ECyIeIeQBSbmz+b4OTWGAuKjdvz2GhwVMAy6xxqaCgPMGBHqubTEbso1snCML1NJ1dxZa90b8wjP
AKCre+Nh5r0RXxaKHyueM3HW0Oh6Kt5P50a1hs4BVI8+kFUilN5kDxT+ijKQwu+xIqx016X8GDUg
urs60df6q7I11pNt7akZCYEmj99p/II8DHZTTLE8TanibzrvhrdHHBSs+OZkZvk2LeJc0tx3Tkp8
6qYQbercLLFfLkLs/5WcCRU8K6T/UdiG2HwD5LJo0BWcztZfqz6JdY/Kd5tP4eTgwTtdgCn+CGf1
pcnUtwnkPwiv5KmnH4R4KV1HTyu6/CXIym4Ed/nmR4AgAIeBfk4Y7277JOk2MSXE2mBxVrsqFxhi
QsmAOth6k8h7GbqlhFDomUgp5RuPKGSBS5GSn8W8VluN8+FxC27zY1tadrumnjE/eXfN/QG3Xhm6
jCI/+j/EUE9h/Tht+/yYiil7kPHLHgEQs2EKC4VSC8K1Oij45jRs9AqQYyckF1c/2moxBHl/usb4
uVRKTZRmRCTDtFl7a5QZHDlk768XZ6jwcPv0bh8M2G6Yf3drps+Rq0N4iOWwkalpi1BH/MU98MAs
Rq/75QnIkLqGhulZjPb17HAvS3pV2IKfLtaKPdys9zjt0QVRmL/I4s42Fspc5GozI1W11d4u64WG
prA1oIiaUDM1IrHYDYf31fnG6eX8sWMRnOLWLk+vMuTdJ/IiFrTIzNHvRqR5t4Jeyxs0Q+krqfQk
+hge8TxfDbq7o6jfuE/7GCoV4LZATf//zUZCr8vWTTAcr1f4zg+mJLXcCKh+h393psTJWLHROeH6
L5dkl6v7NDwTT19E91bJT7/mTR0XlNg6YOSkSpa71AhgfYUnsfI3dzjJBjRH1aCW/lB98gt1jyw5
pyu8lGQxMJNXqvhYhuCX/wg8zOcp25omv4S3TpSbaVNURx1RcQDIVTjLsd+P04aWh+b7utsAqGjO
uI1N+ju5Wr48PZWQy1scsWjrv7FWwszcPaX38ByJbO0B0KCpwX/vzLQ8Hu1VPQ/Cwa37LiUr5+l9
4MTUKjaWtoLDuIJn+qC244sIr7bOm8EBPXINNVJUSqKPOZumA2eKc9hUKPmFNeA0emhs9w3jjJ2y
MCtujZSK87tOAG52tT4UWEHDu/xMab/6kjKgoipCcxvtqP1+01Nlm7MAFPbLrOjTrn9Cp3+OgHkU
bHdyuvGaxeOBNNFqZ5KYBW+zvpho6rAdqiSwJxp9/327bWRZEqqCyPfCqKsb8pvxHzWwZS56DAuY
6ylBige2oEKNiTe62ZVw4aCaNrSyESNIgu6hIBEc7RaXGJrGiAW8T/HAc48sXBXqmTspctru0jFh
vTg22D02xS/SEyZtMYjJuYIRAWUTYG/ak5dud2aiYr43OpNg6LNGTj/WM76OM66rkuByo5ekrfUn
tCtgCaoF7XcXU24u/PXq99WWDx1RPCW0uavj4S+DhIqXhAyRwy+zoPV8IBgQyexvQFOMf7vDGUSF
R0OLCu6A2uSNDXl1euZq9On3v7py01KWd1GNRrob7vXzkM8t+O48eo4S8LxzQEeFZZAfzK6lZAge
Q/duYbqWciUkaFugTYkzyIaw/Q+2JftsG0/+YgJLFya9mdd+++NdJ43NsKW4P8hIyvc9d1/kTRZM
XMP37S/avmIVo9r/ZaOwrJlRmK8e57lcjqOczKsqmQ2dVnhbVCmOoFzD6SJAdCXRlg11dSGTriVP
fZjV2vueIUK4m32cEDmkjJJ0Or+n+mvCtHYeuI9QkLGuZaOTTVMRlJA2IYBeKS7UUsfjUNldSYV7
xlR8Dmoa0EDQDcl6J7+entwgW9W1FdzrGKbYbjg5If/crE/a/3SODD5p5WNWbpsAMRrCxfBCn5M1
fMezh3ukWhzbZC2A90G75zQrm1U4LtM6cn34nmf1HMeGwsfzVBHcLayZGhnBGRUNfmTprWBJ1FKI
qjv6uXL+Fe/fmzSsZYbblbvlFFLlWFTFJ7+DaEdE0/I06dCkZgMSSOIQAskv6XlE/qlGmc7WHQu8
92vLFB5HZOX7g+s2LJ6wH83cJRcju5Rb7avGU+xoT4LcfKmUE5Wh9dZ4NTvfVmiOtvUheTDI2Mh0
HSg2AwRfmMquwzSF2wlKTsuw5RHmZm72XO6LrahjuXoquqqVIKySKMF0/hW0tvukM36uUWgSdo9h
7/AdTekjYkhl3Q21jbzHJDwOSThxAUv9Hcqeu+gzngDxYCRlkJjbyyaJn/MPTQ6tT8fkUx/mvDc2
7BEPungOgUH+QOkE4cJuZXfLcpcVNEudlOrl1m8cWldVmbzS2wINTyooZb/Xd2XeIk8Jq6hS1VYV
8+136HwgnRV8gsi/GDKq11DOMpBNtM8yTMD3u3M8m6Y77Me8huoXTiaDMgsLqpTSuDbfnvjVYIRs
+A/V+jgm0aa3awG18OA0oXMwZN8pyuM1qIizPA1Km7jTOtBdcIzQpSZsuI+OFgnTkFLXywGy3rIS
KtfdYJsBsBvE+Y+b9POBLhMErGJkrxRQU8qGyVA8Op7DvQPH3eUnTqBzLeAgL7HCvdk4vEovBK+9
JAxGNl9ia7zwliYtv6qd70yB4rexktCq8WIwTNjPI0+hQHqZUPBObdFkLQRbC4H/NJTk0dPmW7ke
5G4pi+LWGL6woaLf1P+6h8PoVRM6T/AML3Wl5iU5JxkfxpexmDncYqokDtyNVfGiOXjRvfHm56s8
FURTCeqB8OUwh733iUAzGPPW48F4mfKq8OocyAYErd36H6L4qaTF1VOQNueCGQKNbGGCA2HPSxLF
TjGYbb0UGpRy74DXpmj0HvZMl6zyRzdBy6a1OzF91yEIGlAnND2ZhPsAyp51+SWb+4daW2j32W0T
esEVXWVK2Gswm+o3WpvbRq+XwGKsW/+kUbqI9HPHhfC8rS4F4m3V0ULzSf/sMSY86E2hZjB8Rgoy
wCjJzVqZpSvNI6Vc/26TSHtYc50KGGd76CgXaOwvemUxF+HL+r9UUklEojpQGaYz1ez75sd42w97
fkskKGrUT58oyNGkWtvw0yx9GzhWA2jYiNmA7N+KQrCrPKFFtM3upf53sXhzeq2+/jRVdhoM6skW
vPCuMH4LvA71jfiQvr8Cnf8YzuqCZIWDmHG65jAG0sYP+F+qXLczc+SAlS2teWK19h0IEC0p285X
Tt7mls6cpLag31yENj4eXZRKuOmvXO5o55WXjkberfZ3tGrs7CSXbB0w6+puxTvT17BkO84/nrlx
a2KMZN+6/rFbl2GZR/EKZ4gV9q0M+CXV6VHkY9YBlHTqQ0Tr/+5L0/kSSfhzvHZTnK+F4aE2rawZ
zrnOSxdJL6pvMgyGcFnnMPxw0W9AyblFB28DlMdx+Qv0Ox1K+TVyT7lIfgYvLLR461OEhbsBOnli
o/zVR3pno9A8oEl9g2jtMyL4o5qgH5hqh/nHIUAqkayzqMuPgakx48/SbVBGOGoQqzRIC53vU0U7
7NkwKIFAnH5JlzkW2GRqsr/pGtCvagGgJZePIY4mn+gyHZujTcyoE9eMJk3gbfr8la54gPyNrgVo
PLxCEk+wnZcc82SwpdlSaJiiDOidENm+WPf0HPw+awgLPMgeRB2tpN/m/51C1xym5FarXFsXSCPo
ukdoe4L3SFKIeLqWw9EQUjFTYnUhebfnfMkNzMFjq5RgXpbhASOdzDR/sdEePtqas1bRlZ/C9L1X
KEXrj+tWjUBIIwdEBWA+VehidhDg7dzwOBRGA63ow793ILXi/379Tm6GOXQsJgveNv24CpI0h+bJ
cC/SuypM+Gs3nEIL88boSOV1OXoVDh8SN4pUPcAbUPL04Vh9Wcv3nPt9Fx1EsWPHiqGnn3h3jaiV
GSB3VQO71WJ5x8oYQ9T2y2ay/ejLPhxBVh4oQY31Rf1vqyGQ32Xziotu+Ohe15WNSiR9zWpUuyUD
dbYbecs7TVcE/K1KaIiLQRsf4noho86SvIeARz97wsR2wxlEv2i7CORy8bQNZPOwE1BoTIuW8TJT
9l88cBfHie1McVxiZlzV9PZ6Ia6BRO2e1KkXEJIjyER51OeMElH0FquPYvr7Z6RyAc4IV3/lUxHq
qH+sAR4rj4C4gxFdjm4DT6C6uGklUGd8ui0Xk98NzwCZ+yOF/QMTk3+1vuVRrCarXHkFWJT+9iFB
f2rDqa8FsZihpERxHQkVVleLXfEu3WUNAVvruAR2YSi+IadLTMBJmQ3GOfRwJKmdaeuYek12ydvD
T9T6yQxIHXJtGDbQ0QytFveolHWlB+9DFSNYSRjo0hT8AqQgIstTGDtF2ua1Ahj5zwGljXUm/mNR
22vNxlkBeRYuN1Of5gFQDXTOBetWcizL4LkJh0sIex1rqCvpAPPcBSHHjby5ciVkrak/q4AzcacD
psGk4Z5BXcWe0NAQSjkYmIIRz2dqrwomLeuJiSwVLALDAnUZM7zNj04zuwmgPbsxj/vqPzeuJedU
lqAzlTbinLIYRhenrhpyr2xvQPaNMOt8y9uF1rvfeXMH9YMwJWmHGCFsGJNjZbeN9WAZBOYPb0AS
AmZAM0ShSS09qxRVVjN3calPIq+sJMd56iujU9r0QD2nuo9tzDTBegfBlbpm5ny2Q7Y/U/k6c4yF
4/tpYu6gQFIsdCsJTmzAZDcPDC1awANDY/g63+/ZhasB2u51lM7noiPgUGpZCoGwjnkVeS49HzQ1
w455/0wUYw+qQ/KQAK8ZV1LwpujpTX8daMUM+AbjQEvzRF1Xgz/lLAAZBHbHzfSX5jOnD6jG6+Xb
WbxbU1yGJtaRR4K5h5s+HtOFbu/2SyFJ29t2Dugtmb3+7Ye5XK7RLbTmn5iWPSUzoHKy/id4s+or
nSYa6eg/P2laNm3SUxGrZ+NHFBDR9MoaYk0USadC+MYgszp6+cPMqSHwNIlCC9n+G4t3e197l/fU
qZr3qt2080THPhiw0Q/aBlNX7yG+OVJG101bHpeLEei7CAE721Ytf65pZcSiH4JDJIJfheEhjVSC
6/3FE2RdN3LSHbZ6+rb6QpybxF3DeJo9nB/ZfC4Prwu6FNojUC+xBss87FNksJ8atCZ87b6OWa3L
zAeG+Nl2tzbnk60LhPnKyMKOw38GrUZoVAWqEg/XUyMpaN/8a/FdEMVca9HxVpRk829ShnW7PMFP
bCZkAbEODUPN3pbsmopAt/avpnR+6iXRu2QsjPSfyzr7M8EyoDJ+gW1LIbRb+41EaoY5DX4/vzk5
A4w3yX43IifVJZVhinFi3ZYSE9xxR+ri5qkYsT76U4pSqTbrG4kekFHAH3CmFoaa549kNhtKrnd1
1RWcAlQ5spEPVlk7NeuHHISMzlXtviG1JgdxvQWiIpnDVKRCkdK8uM2kqYlaIc0Sn5LIIQ6/uhD5
ZNRuhwetx/nlHT4TvaRHBxCUV2/73xmd3mJQtcPZZNqCvyHc7LlkXCpv9c3xJaGfX/hj+4Tu4Kty
qXFTn7GQWQM2/mrU1uEbhOYoV4UHEP/p4RFUiJYpowhnWl/a2k8UWau+/TafQn/uniNqIkimCQKd
8JjbrmUFqeZRmDxQa2J/sE9+/pJLPi+dDC63mx1YQBrYOdEvSrB1d4JFghP2GBd+9wUw4VEu7F/F
nydlVY7jdUvRYUkUB2D9cD2n4l2iIN7K94dMN3c8actVl1jtb2vLU18pA5qRnFGVSBjThth6KgKF
EnIlTS+AhRm9JphDZnspcc78/f4Ff8bdw95opsfC4UCwr1b1KvKFt/iGUlRRMPOjc/aKGZxdvwj1
INUAuT2OpbFOnm/XyIp2znsCVMwy2lL63LPiKZB/6V2BwhSl0GuiShtgukPkY8wEo52GcSDx1fpY
NQ3lwCCKTmazyaTKQkDIAJXrwot+Gq3EYfnBVEt3AFSesPl4tyc/tssKB/tceZH9Y/A1bpSJjWHS
FnJC+zFxi4+Pd5xqp9RDg2Q0qsUArerdv4ktqWn9VSKlouCxv2d2KRGCnluVUyWHZW6knPHTDIOr
sagMi2FEuEPhkx7/VfcTezvSZu0B+38L+wrjY6fRwKhmu1FeUzz3ihH58d0JUd79PRKUKxXYJQ1T
jOlbu1D4PPWS8NCnP6o/sdOR3x2zeegk2Lw1rtn/r557CwJGv0VTeAAWU9QHGt+xW8/Wtr7S+nG+
TuwoUpp/QAMywRevJ2iYX9P/0ZxllLhuBdkrtRpMBS2qnRhS96ObvxZTXeItmDGQvMsm2AaXeNDD
wNJjMYPerRyCpPyY5iChv48eT0TWBIbpoGN5FmwxydfhlJ8C/VEKaE1cRUTOMnZ4R81bClQt4iU2
hawpUcr9MBDqbhgdWVcKxTUR0r/9kspuLWp/+ithbbKq9A9BKJJ6vYzcLSjBFJTvzsOn1P7RhGUr
+Una5p6YIDYbInOzR6ab6iJvGYsIcMjbe2aFyXiLJfS2kWlXBeSyUycWJnL+IZzJpZESupYprnBK
uTqtHtNDmvi0Mfj4eW/mOt/5PrWtAnM4XUS2BgN9YRkr8AhsAMmXlLsOTM5K3HbJu0TVoec6u7yI
33KS3T7ozU1068BETrXt1YNrdhjO53a50Z7fqIXVTi8Hdye2jK/hpTcp+XMkhGWHQZM88lRqTO9q
WDO5lwFnbEUJHgpvC5bCR5OKbLE9KWJ80iMYS0w8bP2ADHgbcCep6uh7C5dgeB4pv2oUl7PbPXlI
SNOL4CSqBObiNHJ3EMq3vm4jQImevadmqF7JfuAZcOFiz/KyEc5SOr54B5XXkGdSi68dfDyU3+ae
8nyqndA9KlJTuktnRwklbEZtur3M94AHTL51oXWZRpwuNl58VBtoKlivcaIyS3IFDjbIao1eI75o
y/XhaIuiIAHPzG9KlEJYV7iuWpl6dusGgmTKImUMwtzbnNDMAVRdPjHxSzsUFpDHzXUUcKIKH4Na
sH0Q7PCMMjKRb9lsnJk/2F4BqTUtS90Il3PFTiDZcCqDKe0OPwE1pQHrm97MrFOYzCcbYMa6DwUo
aGFyufRCpUHO8Pl7BhAwuLtP1OE59inq8dbi/dDrPcoHnlhVcJHe0UxfXfCFjnJheUfMq+KZO8sW
lbq3wbjTIP5wPE9YkK9HIuLV7vjos1FecDLqa9PSC+/M2AKunNWxXjiFgSGI52cD3fbMiGBpEd9o
k6fX2JGtKclO0PaaLKAH0KIEmyPCt9Scr/wofydkQvT1kjv4w56XGjmT8D+FnZaQVksiKuts3hFN
vWjVtGRw8mDo5/eGHIQPSIR20K20WFWnkrVv15XxQqPp0ry5LRZ2UgTKQ+5Z7ZQICH3em9ijswfM
FV9ji64KmzwBmeZQqrF6IGi+kgBU9WTNDg+YBK4k/ZiTs5LZZIq/0AZe478kx2AfFBoirQ/5lNNS
58lYT+7oda11Cv6e75/M+YhOWSyqSAC7mHrCaSB8Wi2OBul0AixAOK9+m0Fm2vXl/lVV8F9OGFSj
mQFnvlD+Q2Tc9hSOuy8OpgRg3kSLMHNHTmV/kiZk5WLqzy6UyPkecO2xuUalULBghYVyqGkDY527
fIxdoq+F8ofyigtql1OON9+ppghcprRKorLBoN6KlwCDevRldTUhTULp/y3Ba2azpCXNhvl7LTD9
dlI48yEe1bsGtpo8Pu1cLFXpuKt+pXCWTzFLAy7M+4L+5cUALDrFEeQnF6Lqlb/y0JJ22Zh5GkRv
9VLCXtHOzq4jX8OgxSjWD5fCDx7g8Gi6wU9OIH0c8J2Xrd7+FZFEMq3QkJk1l9aRy12G3CxT+R/i
k7e4WstSmKoJC4IEfJMcoqjdQtvbaot397JD0F0Wl0SYmVlGD9PTbWHqyCQXEXHw/DRanYDFCo7g
rX+DDJIcTOQP6dAXn2XwMkRBaBdh1grRCIUBfqgWYPea0r7Uje8LU7vsaME5LMb6VJtk2k0i+yKL
kSYz+pSM0ovhqU9GA/jU3twZ7pYi6jruwy7aQ5AUQazimPqU4u/WgcPpEWreJU5GLRekqzQQqxTq
ca3LfEmt/+rGcwrW72hFJUplCGB0nb8ttXPta3sqZcEzFEVlE2+7nvsn6MWISnbR/W9GWWnUNO63
yygLWzfTk7tIPqJBNEhUb7ZTD+Ikceq5ZLnwS8F4sioeg30K6oJtphCbxabp65M8E14Fey9tVndl
rpZ7zlLvtDsjgKgeRuHfC6XW4L2lKYfaS6Qdexqg8vg0Jdp/2HQoKr0FeMLO5r4xmTejPEXICcvU
N47eqKNSTg6YRyOe3WuDkWMAVoHKOQUsmVvf8qkhXzOLnI6Y6UIQ5IsPctkF8DE82Ns4mWMUhIHA
zvfrwZPqiPfm+VDDjosC7xDklebmn/llVUWymd1PSo2qlDwo9mZ44oBlLrKjTZOfWfSmxLV3dyG7
cJiYNgvvDMHikWPIK0HwYaJkz7sVd0p/WqaBlfizK5YBfau8UplA9lVkvWbdFspZUeM19aEisqKY
iYfJlTZyCpIGeJw39G6k4dH4KGSrBeG7SXgPqzfJ5p3KmIZkePJbu2N6qy23A4XMP27uOHp1aSQM
OLTQ2ph0OqE2pUbhbrngctfCVKEeehlPD94fU2SbwjTiILw6DHKLsBOwZ2C33HQuo2LsGWao8ZZu
Ws/cuAZc+Of1B9uzZgka58PyPx/YVeEpuJUUfFWyvbd/6ZFfAiP3mZ3YPYA1RD9dg3yyORmv2N63
hr1uB1WnKuB8vCI8hJ23Svrdk9YnCQ0/0D6eMcBEnJaA12PmTNInKjYSDC0axq6iyTkxyg8wifii
iVL42rTIJsoqKZvMFSlgz/Z1yIrW7iMSNSL29iybexKAkTwGDFilba1fb2GMdq3sSX5XBK2v94cC
eoSjxjUVfd5b396tXWSZz0mBF99GBjprFI7icZkHl9oyFJOJur97t5xh/QTKPuJkVhdZ3dpNdldd
zFSM7V9Ot07GMW1jnlln0VENrUYTM3Q31gd6KdP8f5CGu8QS4PR5e0LzMLAIaM8nTJSxiHjsMczH
IH3DNk729NL294nWqkgMW/ZB086dPLYQWajQVPzEAbc0g7ZLTKSEx5/GdgkgK46n6hC6gMIST4j1
B3TihWmTbJ3mO1Iql9xf65hxfrgYwoplgSk/Y+kpHQiKid6nyJ2aboGPzNz16LDe9zI0XQ9A4M3y
mgtomDr5zFQkM3gSu7RifMA9cYCekgtDYATKavRi+zYqhD4IP8SMTuvbGS2H8xk+njx9o68V5dsB
qJ1LjrsgY3FMg4YxCIQAAO8NuRRl99fWiFmXc+VkVv8UrcASdeLdS7UHvpIdlGLw/sweKrNTlBxc
a0oK9fHqtV7mDJorMDSCHUyd7pi4jxKGLc+RFY3jwqILMbk3EmsVNuCpwyL2YhNTU4la6V+3juPm
JHQY7ovf9CVo4Nq83id3/ngqLk00D9OUdt1iHjjrSD71E9pvj/MSf5DMrZLnK39jZD7oRVukg32O
ZGTIypLrqTeqBh76OuT245UOpLzg56lZFEiWq/Pm9VGaP3tnlgNA8/rRrfkNVfU/827JjcDX42Fk
gIaZgqFTzdVhO/Fj+kJjE0xy56wa4EyZ26ziTPD/k1bJILMwmOJH62b8UtkR6rM0xhBhoKTpUlkQ
qNrsTV1w+GHfeyDRfVvt0WB/mTAH91v/Wl1mX+tXXPGgea+/1wD6EpNBO+Kc390otP40qBr/OkM4
Cwnx4xkNrs5IhuREWA/hgMJpjlLGHE+wBl1anYt0EMrCA/2yJh7z6lEADoCy957kXd8lqbaH4+AB
KfWbyOVGjRbTYQnTBGPpXfWyAB2lMQNxezId8hqzQM9ZRio0VZ/2SiEQ/24a/WmIIczodj7jkEqq
rsQW3juuFkkAilZaBnroCzyoQUGUzZSWlu82Q72fSWNymPKjo9NTlukMBg2qzEenSuWEGdQ++pIF
fUjq4J7x/RDQAs4OdZzv0Hfyy6YUlWr3hDf+pagUgsfNZSUSO/2P0bE46AeVd73UKyqKaQcMhaTP
7B3l6Q/Kml2VEP2WwN3A9VZ0N//0wlOsia5JwDNvNzJ+FQ0+64kJEBang589eGwwn2g6QVkPm7H3
7nttUt+7GKLKOA3SjoD9Bb87IE2mehX56vAovUQ8MhdTkRS8ceMUujFOpMkxX44g9BpYnvZa893F
M9zjouw9mUvry44Y4MYaGQkEN7BH1Iv8/IpSx66paaNWX3rKilnb2CR2YS7t78Rqc/935yKYCcbF
R8f1qk6khf8mBnLTTSmyqvtAOf/HvZ6dfWh9HhlhHLrOmURY2rDKsRf0nt0+swuHus9PDA4pGi2n
E02Cnks11KoC9KSERL/9KsipjPaXjq7WSfNRh1j6Iwetj7wDW5QcTZlACl5HuVHUxRv2tDvglCJb
NiRXX13BpPYGBOggvS9/7dbSJFNy+H5tLx/DHLiJeQa3pYH7hNwqXAqJYWKl/gfbBDW0/v/uU+VZ
RKtEXaqHYTxSrrHQgpHg+ppHsmePTTs8OLmKT7Qc+mgEXSKlRjZnbjCzzpk0QX7CNRtom9D9aCKU
lfbqKkj3+5CcZQD2IPQ4HtM9irfXqYa/Qwf/y1EuNRf3ecMqX9AoYnAMY53jXdfHX/TgS2XT4O+U
86t+xcMao4THEzOxGnsL34oAy0huxqTkwhsLKAQQ9jdDVuM96P81625tSD3QtCoWCqG8jvzIscvw
DamKNiylsssmuxjiJzoWmVee51YR6RKmJ54XBxN4gvV7LMo7GomElll9E6Yrv9q1uOJdC0XXL91i
knVofmTqhVmP1TOvYEgnunSSCU27luJU+zutozsdUuCxK4RbW5qeaD8BnB4mCQi3+6fmtTS3VhBv
MyjfwAyHgMZt1we6av5MeYZTNqqVqqGxoFhH419UFXKDxP3+C53MQ7Oluakv2Y6gJuvRZ4PruPX9
LsCwY+vuq8AX2i38cmh0XfAN3pzM+QGxT6aOU7a4gkIQsamxOc5ZuHNvUVUIddAJMA6aeK21yl0j
ScnqHf3mDMhL2Qtbz8cxfId5D3o0FMtkutH5cdOP0GoYMo7/rgQDUM0X2yAELhGwCsRYRBZNK0S/
VUV0j+sSx4BBJcJ8iMJmbsGItn+1/IC2mzj47Gvz8FiOuaTggGitWwxGV94XhAXR543Jq6KWi8pX
Y3JjVNCLaJZSmGPp0f1U75yrsPW9QdA+k6aM8b6Bw3GUfFhEMNJzGj/Mf5QBC6N0Cn5dxrXiDJHM
qvPK6Jr9JIkZIdQZZcAmHOFvKX0xrmLVRYeMYxZPf/rUTi22lKpmzg6XIQYeIIuROjeYM00dHo+Y
XMtNgV9wGeec9Een5319H6aEBCWL/4FDFyAfqmi5/qkZqm2lI7mBgC9URXn3Cuj7l9hpTW5MMMYL
oDWvYAdNuHsvw3/+efvr9OtNuu9XJIdN6SVDqALCVO5H6465OLU0vn+cnM6nNy8TrybgeQ+bNsFZ
LdG9LM37U7176a1VX73DYH/Xflkp1zjO2wI8TTK8l+KgTSALhEvHrXJjOOYjKwbzZ0rhSzSR8pRl
JVpa75Koe6ylzzAPB8kh1mYrnrdkOcUfSzohs+yah9sZLGIylZLSWcmJ+RL6ask7k+wa2GJTJOqV
E07UHCvO0f2Tc6zt9/Di3ePJFZB/QrBZJyx7JgXv0xVMOOoiSzdlZlR/xSxUuouDMxaog8+e5Bcj
PIrC65ComqgYW2VRm7u1YlDqx9y/SaGcPtpeHGsZe/kiyeoz+yQsbprybLafBhUuFpFrO5wqEir1
f1wY7zR6AQ8ic393knxJtJbkqgeM+yYaPLevmTcGLXPgxTIhihjrTg0rTkDses2Nrji01xQeO/iu
cev9aaMwMeUm/1d/y2F23wi4Eai1HqqjpwiI3TE0nVGEN+UYcunbHsuDiuSeeG/a1LV05rQJpcax
cQlNyu/VKLuMrUoX9aJ4a21JlMbEby8dpQc8mZp5931lWnR3UD5GtFELhLMzANXSQ/ozA3wNzx/m
qJNqmXZ6FlNSZ9QY4wj28m0H0zYWgSgXka/UxJ240WtqV5rLBV8xuoxVB1dHQauA5PvvaG/ahde8
fAVZEKq/nR7RjIdmARPknVPvhiMitUpiJPxoKkM67RsZNa4qIBQNK9TF9RjjNbEb/qsWSjvmm5zi
hlrXFylhJqcHDF8X1lDuo8ZzNlDx0Pp+6lTtfzJlYOqpMcopazI7mzf9CfIxYAkvP+7sU8d2XD0M
OrwLAXRatuZYsrV3VKI9IfukD1dNA7mGbbRzOyB5h9i5bILSQss2/rMV/uQt6kDaGxKz7IliSi4C
67qz7nOYcLUR9TSgP7YoxlBH3o0sSUr2cqL7JvxrWrECGzNQ3yIBNmQgGVPqhDFeIiMIVVhfXzEH
NWYNJZ9Ge0J2eBTJ69hsvrsjOfONlmTzhvgoFBdTWPADnrWqSdHCokEs03nDlqm5zumhG9RvyBCE
3RSEVqLAE3flFSTEw9F/9sBzp1ntJTg10nagtvJNHNjjY9ar8e/jAOw1I5FltkY5aeN8kP9bQJMB
FZj+0iIgpuXzZtIq/jRnWbKSYKwHeZ0Lh+gsV0f9O5cY6AVOTxG3UY/HordYFAExab63jEJpELiE
h3WtMJM/i+fwERCoIogNZNPi3bgIStTlzg6X0+l0ljyt5eK1A5WPfiit7kAt5j1D9AdfLOjXRt63
aERyyUivUgLEU1oj8VOL3aJ1NtNEQhPzsodcwYocvPKLkqDQ4Y1nWqjldMaoP1/kjaED7BiaXHUM
+5tOoLCK2jj5LQUgpMh5k2T27rPI6jGMBMufQZmULgTDqvsdJDn1kbtNgC/0khPjfb0yeT86lbou
wKMK4wd0+r8lqIMpXBuN0slgVKYoU9EC5BVSRgYCDCRxfRytZ98b61Rw/gmgtyHz39mESnHi6BfS
uuzRyRvRmLsE+1szqlzPloHKSMI2yMjkaHb58hyzCv1X61Ovi6S1mwKABhiGcKb/Wtenhi176SA8
IpNcfzS/5jcDjLC30ar38fF9FPgvH2JMQJzxlviRGKA6bnlEmnOIXI2qY2AkdttTwPmTGwLe47pa
paecVR8RO20E/F/EOhojm2iqKRq1q30PExehuvbmdIX6afPVnPFdBHXMIIL43dbyQDwB45dBzTCY
/n+bEFY5TGAjcnPPnECX5Llz3ZMsdsTxrU8p74fr5+rssdMlD4d+mD5lOXbsAXHMZ52VDPpq9FWn
e//olDJo+s3Z8fHkbrGqur/97VxYA8vp3x+4R685wCikQY2iHSbk6zQCPNQVYByhmIMxgYtHiJpB
viid2JdVHwE7N1S/LI/6xH3kNbm51zYoeBlK6LEVXGDSIEUzyB7xUjbT4vdwJ1I9J5/A3/QZHS1T
C/LSDS0lyDqYzzEa6AEoaXTbY+K1luiEUjk4kXWX1e3d0pw36RDOfwfE5sZp1XjIcS/rFxK6f22z
/Wykit5ngVBylDUqERS0GzLY9ERLoqCQQYPbZurCOZwkCXDNBIe+8hj0XJU3z6+FUamI2JSaaQ7H
WiSiJEUp8j+mej5IEm/0Td+BeWR6py6UmGIFFJ7hvoKxHjxGAI+rR7SIuNWJIgdsZIQwe/TQQ4PI
4CPyJZPo/SI7493TvIckcfZp2tpcwvQAWhe5CS+8W7dGXbA3wP9y2E5ZcwxapEw0fG9U2dONzzPR
Ka3cGRBJDS2qXGkB0HZw9/kdHPHFT3wpNyqxbSqfUAIbyuIpjRDBDe8ByxGeSyS0f3rfAPJGsKQh
rOXXHAFmRu8Mclw7Hb42h3Vf5dxX9xh+6TiHO3D5a24kCXz2KtPR9nl27i11Pqqskmo/ZnVHLaz/
VrltNEftUG5pQf/EExtLmT6XQAieNQxR/HIl87miBRUEZao1Cu2tjf048CrwWsW+XvGt5gKcGeFO
0aYk9ow6sQ/Pzo1tAymA8LHqycf2oqIBva7pjvEg0/zHSZ5PviUhAjV4L5BEk1TM+ZsVuQ5Sq2Mw
UtBmUWVPBxZXaWhzx1bZBSCu2q+uoyxxa4CcQTUNam6kKJOybc3B74xr+5xURsgKN4g3JsSUwD18
51oYcEL5faKPTuOkzqq0qhfRh5oUtljC9vm0enyMKdvqdLALJNrFwejil3jRF76d8wd0ODvTSKHY
gMKaGbNFnSOI5DcKxrFHLjUl5YPevKecTSwcoLoMZsK0tp7z49bGpw3ni/I/eRoBQ4qKUX7IV4IQ
RSMUmVN/N5ZwwerfGYXq05yuHUYe0fLFiNgjB9oZvXd3KEAUqOVrR6+iyJgPI+9qw5I8IDzngmSr
fLP3vYca5UzGA7tBmVQcNWo8xTe35J2gURjApY48uftpc+xWB5VY+A61CRrzuOQyNdspegAYfPPs
aUZF+zXRJHzDv2wdJuGVMZqqKK+47BPYDxA8fEVKwQESRe+yLn6UDqMnPaI5Qcx8gN/NdgY975QU
IkvjifHXu5pJMOq4jIqRlQv98hU/4lyRKYq34BXKK0ODynD2Pee0OXC+ckTSKlcdXoQogeUJ8xFb
9XUIEKfHpnT7Tcb41vn+Nu6AZgc0PJELBLQOHyEvLHhnh92YwBjrk0QGHzpR7MRrwYX7Km9r0B7d
Cwl/T8yJIYZwj4EPZu5ALXveGOMrJLzPpkgeIoj2CMVdYSzSQMHjRRXvxZZG9jT3vYLh5uW6BlVJ
3j/M8C6C+X3mOmkCozfGYhJ79TfEM9otRlEp0yUSB2KaLKrdmRl0ByOmcYFDHALl0ZESVx3E9JR7
9ejyn85v4uywWodWIzf47BccjUxKcV4uj2tRzfH8JuVdBqqqQX97jbAPJsT+HCaV3vdrEPTlYUlO
hz8V3mKfkrGaZD8Jp/D3GIllGn6680ZOBXYw9Amlf76i9+brCv4BN4WERIFU4Pn3+/3jz3DT0EpL
9f1Wli6rSXGSE3CDt648xAv22lARILuChtVEdWHL+THbVHgw7Vuld4BfffgiL8rLPcLtXUXb0wHY
2l9j3GuOQp21bRe9zuYFx2eBDEOR4tLu8m2clT7Y2lJmf6YIwDIQZ3E+TXGC19GYj01SWjCpgjZy
BexMAeI1PvfswW/0lx6FFshGCFUZBvFN4jp+wRtEJLDUF86StzUvvrOdHb3mN1aF/BBGOHk3CmXZ
KYD8vfvZaqcTfdhi1tRKZgEZo/Ro49QpXzIb4N7u1eUPhf1bVDTnL7uxCWedVMlDUW5BwbuHGL46
d5qnjmXvWHZEcHVONi/owZjNMYWd7ywMIHj5IUoedt4HGkruUcRndxURQGhHQQgA+0i+N1mCJ5/Y
jOYHqIMX9ShXgKq4waKv3BbCslsyh9uEBhyf7fUy0zzlzYBlu6L8I6BgqMmT72npuIAluqgqzCjJ
F2ea8nkAi68Jy3n60Ey5eUon4SlMOcN2cx5BV0eiwDNfEOk5Xu9XQ0j+qv1jDAXwsXpH0eKazzZQ
krqloEKpEs4srplwDXepo9PY1twP0T7CYmRmLVws2sTozW750IqCezALVhahB65W4UXEIQ7WmPkb
0ahHR9RkD82FW2r5p+PsKCJ27sG25Ry1XrJ9KlgS9UBXrVncwB0lVRjVhRziSZ4AkVanKoahB8Jx
ULXs8xdbCMBSG6K8usbTOkyhXw0/YGfKAFcWf7OYfNhrx3g7A0AaGeNMvajX/gpxcjWSDxvMeuju
SSfS9dqVDqlKhl4DJyvjUNE/UUGYYoNCtQacK/rZHLiXHkcOKW33vvqz/n7YfXHtRfWfwINQazgb
6T4dzYVD98y07k/XPayCFCj8ieKJ6VB3ra1SuwhfS0PFzJX1AdVbwl+G5LpIsWKjVXgcFd1WZTzC
Y7c2BU2AnFPHC6z38jCuUiSUBGe+eLS6Wu+WOtfrJo3hghmiS+5XnQFQBdxkInHy7gCb9hYDxmq+
43sY0nLl3vWUoBFr7sUvB8nW/KtLRWEX7zKPhZgsQ26mtl4fEEW+gnEdbJj/teo9WSzIGE6Pecub
SEAol/j3mmplsoK7DcddQYU9dT2/5tazX5BPZ/q/zjvsCzQWEy062QPYERWRj/c8wnaFNoHbfopq
cTHK9iOnpWg0/tFAdV9WXeuaLi1BFxJocjwHwM3VM5dtmirLawR1MNK0rRr2CJs6dlSwHP//LGd6
3xYPm2X5D+ixJVvAk59fWvXsFklWWA2uEsW58J+VhpEsKBS+NjnyNF7T3sMQOw6doY/vUKEp3hnB
C4uTssmY3dy34y2VmhGpRBEHbQY+5GAXhwmGyntfqcEkg8wqZb0gdRLYZLJQcPTOnC2snXwyGAH1
k0hkb2UpbMVhdx2+L3GTtHqUIn88R2XV0i+QZnrNnhYMV7I7RLa+9Xsod9O/d7CPWwqDcn5QF4v6
9kAfF8Hk8uumG42cUKwvG3ydLVFHbDFY/W49TqUAhonFNRcxRUvl7M3SPvFiiRmeJoAj66pWFY3r
tGW1Lpy5AkABCZVB7byvORyTY/LCjMzINDK/b8OhUt2hnDKJqmmI8TRW/+VVV6P5niqpedSnUfgM
jMyT/yB/B/qo/5WjxvYs5x2kAWwdJI5Gu4ySu1vrkKpgiU56ttSSNVsiERMudslyZ6G4efQxCMID
lFAHXvKPsJRRm+C4WZqRuZv91Za2A3bXG5rAmPqNHBitBB5OdtBft8NHQUbSdtrq/OD7qdv+S1Nc
dEJzb9+qHB9FGGymLlZSEqqrqNUOqLT7vrpE2QhWwT/9Wd9Bfhv3ecCYuyWz9rNRSAo42fEdmGOA
GeXvh886OcDYSSNklVRh3YkEqeSE+9VeyOUhlD2dIFSQxL01mr/OhO0T/gOxZChvqSK2IlXLQYEu
ug6IihZqNYEIV9BEWM9dhBVM2w3wESYXz7n9Dk8F79TyeBbtg4HhiZUbxWsoBqyAhmrwagp+XyrA
Ttdg1CjvU2oimdazevVfdNxotWKx79wB/if8t++fNbciwtIv+rgMNtXvZtQDLcC0lqN6CmKRX+wZ
FaJJPsbu+SE1VtCPy6uO9m+TkLDgdi36N/glptArBJW/dER+Mb0E9itdv354zBexYeqtsjRLLtDt
HL4aqdJ0RppQbriK53Bx6cghta/TCBpEI8eAo6tuMzvkg1kqfllVBG2mR6yt5gHC8FCGrbvBKpRt
BGEJp3cZDG8XLVxzKrkIdPO+js/5Z14uHGUDVV198fDtyuMLtRZ3fcuTdA9ZeVsst3FAvMAIeZpE
+fOJd4wXjzBWbbTK8Wf+Cn2IJP52eFwj5tRfCCKHc8WAf7U2C2lxmABJYtVJiiq4S89Eks1WN68G
gO2C9b2M5fYI5+AZV7Pmh3T8rssR6UlxdMKHlteLKHHZvjQjqYLsQUWSSjbXN8y1gSb+Tvld6ILH
gBdeqdU6eq8qT21iVxBHstuQILCNbHQlfHsUK/CrUc6+80JlBZhjU/xHN40BG2cPtP3sHUiXrm7W
c5sCxYI9Ugu2hiHzWRYGhp8Y3iqMYlchBgAw4f7ln5JRBStBqSQJxSuvkR5MmZs5hxzXRKe7KXuG
bvJKw/dnAsbQI2Fp5Q0HEFYLVSTA6eJHWMM+ItjKwSW+xGPIFrhU4h2fsjUrTThHpEFoIUh/+E+k
RvYlZ2K8JYBfP6nNgcJ3CNZLL4+t9NhdfMoBF3vlC7VaHgFpYG+mEElNWhRZVQLQgvqUNdADpMl4
fLZjx6PLwFOAnHlRjtELHF8eItvs4JDNZ+LTRaGjoQbDdKc40davleYauMWop+G54ok9uKsCm2hz
0RTM8XJgCpHHNY+U6ViwE9zSfIoIhVCQiLFL+F8uuQIBFgCcvFr0w0JUwexG35PehnQlJjN7loZ3
HLSgsLJjpxyrGIWV86DEIWFKLdVH1lw9Epi79qPP2Pxfhn/fz3QXB7JUDoXfLinIvw4Ml+eCNI3O
HS013bJhJmBu3+ssPoVBTlq6zvtQ68lbxp6WhNHUUz12E1YaN+eJoMRoGp/yJQmeVnTuNpCz0Tor
Xe2HJ5FNgkYZdxa/8mHTJMmNriPo2qAroEIjjjZ2H+D2le0eoC1dYsTbHwhbyOh2ZjfY9H4TGbpQ
Xm4kGb4QJ8q8GufbfFGcXNiP8UQyqqKRBXB5bw/wmDTI6JSewB6ZhCPh6kJypxDpJKH8/y4SGEFi
rAEC498aCTNfwhxBG0r65GdL+nIpShIs9aYL6IH8UapS7rHlNHuV0ULE8QzL1yyoL5AyCN8Cf5eX
Rug7wnjpzdRE1Gh6yu1K/AUPLJ+JxCvSt4yiD06/0JXCRguxrBvNkzN3IdACG8Rxd4QkyDsxI1RP
xIXQteGpiUF1T5BlP7FTtFq6hzxTX5VcjQ2QPPakGb0sLhQeDWI4xC/3w/PEDaXlIpvMDlIpUps/
2ROPi3fwlx8Afa7hVf3J0kJz367Ye7tuYOqTHQxrq13jIG6OUZqNXN09AXA+ctC27fprsgq7CBx0
fyzRt07eYZX2hboTa9LCH+6m7l81fsqpanhUZDTH55zAEJ0+veutfDTJCBeMrfjNMlpb+5+Xcvzm
ixtEQtvp3JdNEWhTznY4RGrFNl664Rm3zDuG/P9aIYaHsG7JwNZ/bDtohJCW2E4ntGPpWkuyOpCF
ZfIlZsnfVjpe65ebxU9X/IJRcVmPbd3YPCEa/icrtrEupKwekV4tDMEkcLerp6vOalV2nE4hv4uO
+10RoFrjQJYunAyDJPhOtAxbdfDQjwz0getCfAElfzn/1Zk9Xz28yz9M28CFa3+YdQObs3PrSOAB
FjXz36kE13XZFy0vTtx1TNAQieZKHyNqzW98ovdgS8tpTyYwTcufttOaA6F8Zc/FV+i62VQPrcr5
dtCge6UPPxw+noUr3CiQExWL/HaROhWGDOQDU3BW6oIjD6A6yXqIhpqs9tplpMAso87GvG3/tN3L
x8x14xH/i7w8eKrssBTOlwa/PffxYZIS0iJc9PsmiwI2QfBxVkrTEoSCHhyd1S73Tsfkhv6C9iLz
g7c11191dE0XVA7/J72Wu+BKwEzMRGWm18zntJb3Qvb5I4OVxvuKg5GuK0e4pxJIzxh4ZTOn4zbs
/UDJkw085bJXMZvIzkASu+cOszxQbjamCSA52cxvubiwK8Trxhsc7d/CNC4b+hBoL9YpRyU9JZwx
zM19s/TiGNQKl20TaoAHx0+aux4ORg5UsBPz9oROFrdUCsoxOK1ZA3Sull3QqhK9+JZvZX9rFq+w
RqIsyjargFckP6fO7FaE+MWl5SAQtZYtkrONU/nQxHtSqbkg93Mj/lMKUQLZSjWHhlc5qlVE9aI6
wjrkWhM1MmHwtBRd0dhy1BoNslp8RupyrrToH/hzqFRmjKoombdgerFuxh1jH5AUP7PIwax6IaMt
2icz7M+zpH/ZpMVW43ArHWa4M6LJFSw7ZW1vVIQitrlVYHPvjGyG6l4h+z9a4/xDZfYdWv5BzHsf
YRKRSPBEX81M/gdnFeOTU46G3NqBAjbUyp75RJttzyVSjLE2N42MGM6zjj5GJQQxp3SiXomhbpAZ
P1R6WG7NJlGXXaPA3DYC15J37dnWf+Mq/hulpWP8IOxn4+OzZG0w6okWo5Vghb4iNy7xzqmkA698
vEkk6Day61WdPly7eoos/Opc9Ce0Prn28BAxlwm5c55/IT8uQrNtQq8zRoIrUrafEERlKq+3H+gJ
55Bngned28G7ObTxiNGJPl2rgK2Swa7Goqv/+q1lIJvQdBgpIUOeuZCSrMItQXqnW/WpOp43mSv+
oFgfMir/9VdvC9r8qvIg9QFxYh1SbPqWJNX43ka7RKfV/aBwyJ5mc/sFd9p86mANSkA0bKmwx/4h
XdHXRDMekNPTbaqRKJYx8dM1FA+awurNT05v70n+Ofpxt/I76g4MF9Ezy94Qu8t85i1SZCi0Mzla
BQ7Wyv6BPrmt+UKUWTY/YKxCF5YeZrdFBqRvuv1lO15IWCl842Pw/mzeV3UvOzs2Mdj5my0f4I+Z
YFq/vc8/isSJXxgcIf7br1FUizsVFdUcvrxBkdGJRCkQn3IugfvuCSJcylwItv5nU/1rrU8bLMKi
TscPCR3MfILm2e0kUTI3BLYYVeBBZA04eNyaDy9DMeYB5kFjzcTRmGI1wJ/G/V3LmVk8+NDQP1M7
X0tZ+ZpN867lBeydlPNvVA/qDQ88QmtrOvBoL6wt7nlYqqXSZw+bDlaXezCv+oVqxLHDUGt8/imc
W5umJoTciaCWKxT3uESwsHkfV9S2ob4DPMvoAWsTBs+OWHcd/kIrBZMohMXvpiE/Wcy2j4AnT4ua
MoqjmjAmf84TV5OFL/6rDlgZf5KXzMaqMyeEOf0CqeMgLiEra7aWhAIM9sQSP2kmTLT2wnMoA6TC
Y8WYP5/MaT6fniL+VEHZk37erqqfIYOOkAJfwP2OQXy+Nsj9w2MoLIEuRnoPhky1/EABTZmh4m6Z
xfV7eng034HHpvcfK9uM+HHViygITK+AvprNQ8P+zFUgczq6Zl3ixaLEaNM6YEDTQWwrmo0I8CnJ
pZ5qz9/zsbnEWqgmG7zCzAk5A07mXDE752zlm8PA5OvbtkQsI5WMP//lfcEhzVUjxm55lRjhzc9r
jgKd38T9h/NW69FyXuPOeZ94Zgy6wc+lbFUuieKG6xNCFD3XsVMI4diNkDY73bg+GW4wmT2rJ4Wj
7Krj0rj/1iyoabtuym9DcJCJh58DZsokdiBPKy/4LFl0bFXw9FDIjw9Dko1t34NmvnD5ugjp5J82
Hzg0PDSjaXumOLwEMoEcmgtXHnpefHH6ToyGbp/vUKU5kXPVWl1OFi2sd0Cg8Xrzy336MmnyfuRK
Lxk2URVR+z5b57J1uf4ctRiLot0apN4rXl/Bb0yOYmhgEio/tJae5kQHMnAsE02XoqF9zC5Kcu+l
aYRIoD1XOrpLYds7teekAI4yLLJ/Tr4Zc+5PDXOT8ni0QxQgD52Yb1524HzkUIqobuZ5AgeD7gky
Vjo9WZMhi1jx0lPYVsHTk2dI5g6SVSZxqWB5DLvKjmlzV2LvFFIBNDjrgnoznb7jkgKlTYCZaPFS
Bs3YUGI5SFcLPY9UYOTycz8MGngbVxY0ynK5FIL3DL0qKhaHm3uddv13eO8UG4J9AUPucomC5kAO
n1hG/oAIjoL+aFfRWFcnypIxcQU5a7su4PekmZTtdslbW3Y2fh3uB7pYqA5k3G0z+monxw9h63JP
SrjQuu9yjrd3JgfeSvGtktW+Z0C2yjOTVpgpziHoc+/ZYLCrq5UBC9hR3q3OuL/JBJ1n8Ua7LM1g
H326LWTnJGtn5zJ0grtaGBqfZzOn4IjAdcQI0NWorXx7Xr/lEZMn3JvGe0x0SpB+IG8B+PlsQcTf
fWWaeb+qDDqaMTko/UMQ6DClgpSV2yOx0ychPw6EzhV5G+DPDRdAWQ4RiOiLdduSv7s0iyKwsx5W
00Te/esPFW4j4WXYshd5A28R0NE8/OOFZ6KQG3VDkS1+ArTrXPw+arhXOMU6TSlIow704KCBPx9O
NFZ4kb0mZleiR1Gikr0umuD7rb2Xo2SARdIW0mneGVcqA30q24OI1xN4fB3YzXH8MLWJ5T2crfjY
hPygJVsp5HTkcRQ5costI3i5DafqUlYL1WBvPUYDnRfeBNxsMEiJWIgPRa1XSpvVrMk4eCjM1BKu
fFxcxI+F1ALUXLkwbdLyUgJWSGqj0PvkUDe2F3ZcDVrS63bDwkSikTvK+6FOe2wY/RHv61WPkJgz
EtdsYatgvcyVSkQSiy4h3W9IXBMogRkK5K/0aaK715UPU/VsSG5fyISyhDmlBWjlkBvy9UJQkZut
9ObUf7sLkloHpcNBxU44j3WFIEKg2ohWvmc2HYkYY12ormqcw+nO/pXb8YR9HRGzGdS3EQpzW3I/
C13ttS9AkutBR+cQHuS8EVSvQL7X1Tq2roPtZ6kFvzU3Cpq9nrGhSwgsUu9+eVtei9W7Spa3VzgU
Q8wwMP3VAxGSCQaaK9YokrgGQLZpLhpxgcSW8rOnGIQ2KJeutYbHocdQNmbEWNziSWo0tWJUfLpf
War6e0Nmmw3Zqb9wBq79ARKomb7FNuejy6FnuJ7otWCIJg3YmnVpQRhQZ4604m38xt6tXNMjkMrc
Ge2Y3W1Suwx8kPA5JVKguCwNZm8erEZJ3ZwXMfoIVAAOfvMr4+xnpus4rwvYCOR1RxnVsptPcRfD
O/go5pCf1Ky4r0wIWY09CnVb1SYQ3HyI8kgHjXLCjeoNG5ipJaWEXGHihxXFTa4rW0qVHXTWA8xj
MF3XekzsSFH63753KPoMoiB1Yy9jFnilzMScARjaT0t0zxoR8xa+Ebp2TOEJpZ270/DbQgYWVP3f
yRS3uUqpFdBaPubZ7Fz3vnboVjcXOWeEaeiVRVHqlpX2+PtcZDhSO7m7V7IW2JQ9J/BX2cH4J0ac
PYFmGRkqucyH7JY5StKUrkYMjEGj8lrj1G2cVXgo3D1JsC23FwO1fvcJ9dL5d69hQlFXYirYXQx1
HL3Y7rjnrlfk4ozZH+XejXosL05GHnHEWVxWeXlC5E1MwTw8Rj/PZEhIPe5wl1OsDxJiuqpq59EH
tDvEH0SYUlypJpbYZ+bdbUl0mBpSGLQ+NhiAoHSP5iCe6HkeaaA1vyBdbxLQBkjaslpICmwk+udL
GSYgQfZL9dGspt//f5yU/RIaEoPoZGQ+tfmBqJaz5AllUH+9DC6zWhhAfi3scdLW7ibwKryFMVYh
YJ6KbI4ajaKDt7EHO3B3c4FutbqBTOedsx4Lbuj3vDcIDREUDlFEWHMmO21p0Q+BiicG+F/3u9u1
hCptk7lizVuoK3iUhDfbLc3oT9TTRKwnaNJH1mfwIWGCnA4o9Zx65RopYni5QW/TmJrumlUD5MdH
Lm0t5Gjy84w5eajnc0MoU2Y0OeplqhLGFBMffZpc2+km36Vl7xQjF+/JXVRjO6USxsrEg3bNW0I+
Du7SmNlPeiL8QYyfpknAq4e45dXnTJdrT4tYWIfEp1uX6CTBAmBrFSlG65maIAKIhL5WJCnsm1LC
XD3JWKX1kuR84ll7mBGiNLtFhAZFY8Pd+6ab/s+mFbQTeW8cBYHarwE4YUZjKXpGLwklgBDRjt05
YpNBkLpuz/QsESHltMjVkcznBJq+IPuogWuzFOCj6jKd7O7ijMozUTisuw8MVVbnTfRxWXx6Ot7C
aQuB/WZiIbbA/6DZMAqZU48ZCxBYG4uv2AG3j/VjKZvqVIlnpjaAimWuRCPrGylSspH+78TX0rQd
EkPGGlowQO8upxwNyoOnveTDUHtG7+GYFyd1EXhWCpzRTGVdlXIruCmlcu/tt+hDYNXCVq3hgtmP
qDUtZkFF1g0mysvagiLsxy10nkepcqqp8QU2UoHPE+gaWz6bR979KAt/J5qJdXnLUNYHfxmHicI6
IYfyO+QQJw5suDrVlyt86fFcJQ1TqRHVLs3hMYLxBCtgy5dSAoqTRMhSvsXJO412FC7jiTGVe2+A
5X/8uyTIWSJnPZQp4NZE923hDgLdpFLJolIQPNGy9mLOuKi4NPENxbzhzUoJ3l15CqGIVxOe+11M
8qQaM4y9PFgJgh7VA9YRQq3jR29IY+L61Px3E+TolYfCu2uG5xZniPgSEgooYjrVe5/maKiQfWnt
YGPihDV5u6q8Gvf4QGizRyooLf7lh+b3+7qR8Q4m07wWkSHELwyKLcHjUK1EkTocn6DyCg3BEA9/
RG57tr7PbxDGdp3OsQohYeX1farYPPrQn7iXeh/706aRhVvI5oZj9Bq/21g69twLPbUtMRz+UmBf
YrvgvuEPChDoOi7md8faTM3Oqh7GrijBw7Fu5OiIYb2hEQq+5KG9w3atfj6DTaItq2I2DMY6B9qn
keKdUln0EjDN9GQNWmb1gyNKWsOwIe8BCs48t8HP8mgQh6TnvorHzkHyMCNqCkSOa2PfcUOkEG3G
vknUEmyZgRQwwjK+6NnWs3kG5DM1r+QOgRhz48PP3wWrebyJo/RaiTrZr78Ol+9SHcz5U6JqiHGO
IEue5XpxEJXdT9AbSrOvKau6k0pK0xemEF13v38Fl++x30DZCkFh02mALUyil22XQ5XbAEr6RYJT
oMQZgK/4ZEpr+JZMLh1+8hpnWmDOjQCqLILs5WJyaEPKiS1deoaol8QKYx6bNh6SHtyRTw+lWKAk
21WdqxFfLFnLPG2tkagzN/EPVs8B4t8FTlmkAZHCLFLpv18wsXCk2bMs+vt+0UgUHPDYDTKxoH+h
47ZuQ6j7RMSe3AFGuOavqDeHih6oaeiVoWpOIyDlTGemMWvLA+lPg6b+2JnV9QWfUy4LLCAwk9eH
27/V+dccDyAKsAAaEEC1XHlY7mtEN3v0No4IFW0Y2Wiqehk5I9HABujtAD81jeUeH3e8qsMFb5Zj
3rriLkIuQC24Vmn0z97PbE0sdcwIhrnCqZ/63HYo/AchQxMBEMNjERbupt40nBYSTn5LQOuwQuve
YHtcn/Zgj9zW/qAEqKI2FNgFnUysgXyBGmoWAuiVzqoYa8pMhcE1vJCwprZ4runN3CBfvftgQQ0v
rpSfO7eJcc5g4fGHa8n3sEOAgxWdVVdQOXaXmMq6bJTlw93RlW6pfcpxve2Cvqk7ZUeSTDZk+J4E
eqZp2by8AZEGbtcNFg5SjLPI6mXZX3YKUqxC6KeWpx+/8VCk/A/1z5C1WTeMLRsNMfuDUe2s9xuV
WLulefvQf/rHFmLig6RIimcf23U2hfWoe6oM3eJzgOuPARxuvtRJiMsWOVZk/GrHIGIomH4XIoBg
tdC2O1f81hk3eCvmPDhtRFJVeTPmSAbNBhJ8Uim3WcbKsDPiR8dSSeIpoQkX+ByMdrAyEr6usLF9
Gp325qDJhRfg85vD30ztj5RN1wilNYMQCxUtOR7Xkc37IgWxfCBXlJm++YTMIvBbqV97A/I0ADHo
/kCq2JNwhtagL5X9oepTWIH8USjwrLV/rIF/oEG+vqsayMh+gHza9jehnJGAKh+10EvrBn8PJwx3
4/b2BrV5ukQiAoffnUCl/OJucJFyp4k7prSWWEEfc0Crtlw8lc9fl9Np/lfxscbukuTncwgY5FPO
M/soYA2jFMfFot8bWPSu2Fr3CwuaGS2v2PfrwUevuVGaKx01itLF9bsb8cXTpL40CL6FqgVWJPOk
N5xwkQj87dJFMYhmGofmTjJR5XoYWFphSHC/gJtjkslUOUCk6EF/dPTudGBsQZj1JZo1bNzqlUOm
Yws1LRfOxMJ1jAsIqHCS5xuyYnGdhbp/ew68+Tu6g6jINy+FeQnH/RAw6CEgsPrE9Wt7LZXhw+bX
ZWSWn2RbQYTuNZf6r3ASI9RM0ZG5kaZpz9aY7Ilbq9WJ6QDvLBzC17Fgkxx8ZZgiZKn2qkcEOp5f
+vJaoFdaCiQprI2G3yhJ9r3e/Vjxtc6Ii+0l3n6KtYej+e97nRB8K8nvOhZ1T9hOpOi70dDUP1GW
NMB4wYpMoJeRPANyyyaabYQ4sPk+W3OGvxNzt6VqI+suhCMEkzzhtSlK8BhqcX7d+0YhG3rKFkm1
wAMueFjnD0/C6H/f8GYsn5/52kamf+mlvjHe0APTliJvEtVMiEgI01BMoLB+2IbKceumWH2GahnR
cOR33dpNqNuNoP8IszHuXbfdMmOFqxsCIwY3OSHJVdkc3H0+U+x3/J1WFsgp79pfyTe0guu973eu
vTx+HBYxYJr3rgKzLQq+EAO9h+TPH3/9MtYhKg1FZQbgum+snesqyiN7sIP4KcGH/Eu3sYgpe0sg
bAGFeh9I5E/3I16V+dbatljkXxrw0gE7iUJGUjjK7rBT7urBOEBS3eV6Cvlpq0lVRnDu1qQAg3mX
dlu+DW3QxeP1Erytn9ixQRTNwHWz6p8jD0Evq8AV3qhzy6T0WAqznyRqLs0l4RYaib4DJafXM1vc
aAhgbo31f8cs77VJel73FdSwm8pOpw23lSPxLUySru5ncicRDkzhjhh81HrMEBVWfHxNjSt0CIvN
q5AdZjF69kI/w6hNPi2JtlKaxnO9T2SQgkuUBRvgAiFtPw+i3IP7uXqodU5XGdlwvh6t5Qai7DQe
0G+hlBq8bs/g9xTHBUYeXHlWNLEfEKzLTyNPU312phnjromz9ES8+ZDAEhLjW8DhUCKUfxGHbaI5
xq3DNGMQ6i3hB6bUa3Q2iBGAz0qVtjseMp0ESsWoOuhHOvo4FdNgQtSVR92mcme1TJXlyTPWNZXX
if4KhRcnyUUvc+rypLEJW6aBXypvCvTRf/MwfS0VJr/DnDftFaBxQ2C3kiwjNSiSPKgZYpAWMLvy
tDQrUf4kpJQsKhvDN8h2UX7CQovPnV9CdcmZMvcpYmDUGN9JTwrrOrtj9BkyJL1o8imr3NXdS3Px
dQmZz4/K79VTJooKxvWdnHCm6IZFxlG+fulWfYNIKgevxKslnfkWVVUnwXUumh4FX0iawc6z+Gys
eUGLyqSG1O8MKWjQ6V2Dxj6AkHF34TXG54N7CK5CxT6q+8vKCYSxuj63aihIKQH0rHNtX3wLD2NE
PexKyKrhryU5L6YmKui9S55yk4oZ8Aq2noQp+7j2MFnLhMZT1HuIMz7xLGLRbR+Wk5LRKiq5XJxM
aPs/ilISBO/+MD2xs0jqrXk1LzCGFTMjql0kpd4WhLw9TuCP75C/qY28kI/5Q5F469AyuWaW/sY4
0R3nU2uK5S7NkIBHgC12jw8VkRb+RTWgmyaBAbq/dP0qDnaF60pVUzAlHrUyrGi0tatwJwp79GTG
Zojrkey7GLV1+pQtKMiUkig50eO5pa8EK4Pd9eVGh/8JCqjPyKCRVcc+N3qkWBPWBOVVu+QD8x38
Fh/rJSSepZ5xRD5afPzqIwX6xuVU0FPIO5ioo+DMCPMFl32sMiLzV7zoQtLyCJzt1BTEqfV0TKh9
vBV76TmiG9+iBr9uJYYR05UtC/VcjoR+eq0ZAYFG53oodq+UTokHlLX7q59XvQIRu4KAQmSyhBpc
YHGcy3X6t5UadkhS4G2mDa+w0ZeUPEFiRV1XLVpLbE3+AItjLZR3U6fSkTEWOgABQ5/2IaeiMofo
z3mjrYTJndiVbUTzKPT+Ub4gV+7Ll19XA72AqkHllFsWTlMzQDZy+kCwmz9QxyuZimp0ERedGxTZ
t3xesD+UOEPBh24+UsoefzEANNZ1MBrbonT9bc4vrTi7levzoGeV75gNYKrbjnP0OpeO2KeBxOKv
EPGxOnJHlRHCuqq7gQwL8MmvR0MJc1QP+lCB5FvcucgGk/UibarWtJeq6D1uB277M9WlTHagJzeY
8oZ4zc1RsujPImbbo0R9Sib7Gw4fkfdM9T0ffR73w/R92fQW6beFJS1qX312k899ydg1sqxxcdLz
zno26vi/4Ct/Gxr+Y34wqwHxMDbdWu25Ox1FrNO9jGEh2F758Fsimr0UVYfVBdm6Z4C1qMXsITwl
AGFq8SzHnP2liZtVuTQ+h5bNzoX/ZKsVSmAoj+hPA5IjNPE9p8oHMa9V7N3ITZWrjO/HvM/pDeS7
OLeN2ncI2R1r4TGl+Rxbg06GMlRPEpy1AKDPIxe0QT5s9DirBdFCKdaTTnSzUUYayA7PJbBxDqOd
jO3JBdNkmCU4CwbUWM68KH0pmatZDI/QtDrqzfUDOMmXfVd52+I+t2rEH/49JoUUM27Cx5RMuSor
JtsO4DcZWN0sIoq6yzB4gAEJ7P4OMNbaeVwcMVr8KyeifftWuUSN2rO03VQ2adXW1ImZL7mtr0po
QzLU7EJ3aYW8N6eiipY4fGdwKY/GXTSBPdLoQa9wPb+rS46MTlxnZ25pmHaMHCjlr7dO5uJ3qv1B
73vHLoOsv6DzS8Tkp+fnXGjjFpnqIlw1uhr80Q3iyBjEhTr5G7pUuP0XZi1gv1D4gaAY2+49SHQ/
+C4kr6LVjxNHFAfw6v42c1pzVHEbRTVJi6Nh/LBELBczmmLbSCc0D9WX+CENJ6L5+rsJX5ZOcilL
0NN0LHEzrAd0qb6jPqnNwClxWOYfpgbV2W4H+g9m+WtnTI5AS3yGUU0odLRR8U8e18N0YibxfIeh
hzRy1eWl4cCh9rd/j+t7PDKTf6RKDLqAxkrbKG9MDDhT1WWr+2W3CD4H7Gl/rAySCt0oi97jv753
ZmNe9zFo4jRPaVDxYvQ1RgjbpkW2yvd/g1D8WS83ENQJ8oXAKH/tCxF8+C3ByjMoLBSZvGBbpLGv
wu6Tt2ikyEu4j6lbS4pJA5gUWKcFdMWsAln5AN8VkJmpQV0M09+NERCZ7I7ow2jFdzgXkfxavl/z
FlpbShVwQzZ+IhfWzjHIhllvIwQIjFU+X6J4hjaJuAr3gx6siR/o5HEUaSpDcID49wrBvSv8z5qU
2wUckz1M/awVg/cUWzzygwpW8AS45nrTPvlTQlS1N/qWTxQTFotq2CBylp99KyYmmuYRjVVoNkiP
K1W53+JaQWZcHjxGqZNmLmBGEdbq7YGaFVdmcR0Hld8kSE1CgaVy066b2ec4Wg/94d+6mHbW97r/
gZADEAoIAQtIbyzM3Vvv9jBjvYfBtTjIGQw61wbdPq0/3+l5+sXRXTdCurymKm1ie01tRvLx9TtC
/bOtoqtoN2Uj6YSMxL9ggL4cfMoo87M9E1ej8ymgHnu0OSp1CUu+nvi0Eqb3un9t7oObgB1d+3Wr
U+UwqOQgJ2syUlpEkxPbEzVhMUcAld5NNwFwTT5RYXYeeuKj0R5ULRODhOqD7gAN0Lr53yMpGFKt
2c3RI6gjVdPFPxmMfgkI+2KxUNHR8uHfBowaBPtCUp0TSRgmarRyg0d3uvkJaOFH+8uPE2bFpUr8
MWwBt5cP1+jLx2R51NPOgwOtMlwUnJBbMK5MfDds02yCMho9Do7yDQUBTSJNefcSTzgY2BrTaZje
6eiC8OwKDeG4X9dXkV9O1wZB10w58z0s7oS7RCf6L4Rst2mpnYaDZu6wXlTzHi5nW970l+PXkLWP
H0nPyKu6mTlB1+wdXqkfr10HA4wxA8WE+fvQtPapuAcID0BQDrSu7MrYQhwqnv2opTuR9PgPV3xV
yh2wpVtSsbKXJJ6NatYvuAtwPmFdq5R1JSnfPmZSg20wFrkLGPmcZeeXuDoqgNjmdmqZLqFu9PG2
zUkxwW5ToSezOaNc0tv3gchyCjMibuEKj+BPALRUl8g9AIUglKreRnIaCygbz8bf9Fi8rO037P8b
/g4a9hOsCyDdf+RdYe3bPu8Gz2SJuvZvfn6dvkU/IlF/f0p7A3LfMcKBZWoKVi075Stwv/bjtif4
JhHxrpPp3SmgWFafhqtrufLwYCQZyasFx2cWOT1SEO+58Ag9kiNcNrY/h29hT/dB7s357HBG9xmD
oHRGEd7Aua7iyxlbM7BVJtzMoCtS/0+iteLkundPTekAlYdUXJp0f60QNYiN4U2PMXBhEQozmNwQ
MIru4l8A1RQlZQ6cKPW7J5P14Lc9oDfo4RD3avnN4HnJfVDTXl6gbsAXiGRGu6QjwcbbUuApNKc+
YCmFjXAAp+JApLSncFVwbp3qccUc6B929m/Hkn7uvSE3ntZhaKeF9vpkoUaEUc97or5j+NnuEzL0
B3Ek26pSmc8CbRTzHJa47ddC58pnsAFNYgxQsQLtFsBMXcfiPqpiC0jL9v7vlaLHqDCwD6cNzOxV
tJqZPTciSblr/EwXv6HWYK9IDW4MnLhyK3OojA85Zr7oAdPHdkBGW2bshNpFS4d2Ja36+N9FDVdT
UPPErru0PA9geKHLxeKvV+9gj6xDNTGQC4ylY7Xibc/Qys8V8d1PtxcbQvIETJ8sL2JM5Aby5E7O
5VE/9pYDNsa+pFMt84SH7ScZ6Gc3aSBmQkgE58Z1Pp4uT/XmpMgC/9AlTenlJt/qLNNc7x0KTESa
PqoAh4+nQiEkCwlpD3HcpHP/jSKO2wZdCoTXSS950Hd2SuXyx5elhgC1YX7N9QQ6NZnhhPqRinVN
WiKX7Uk1neUKjfI11JiHNzKQ2f19TQq535gZ3iUWGHgupcFYp+dJjd/XxVRxkfM0T68yCc1cVUNi
6VQtznxI/px3S2CjgmekOAcoCVHb5//dD5GV3i5b8Y7wmnfhYyJ2kmoa35IU9cD43SN+fvPadiVj
07v1xjQQp3EA+lHmnlpUpSom+PHVJcyFMQHv63e8Z+LVZy/CIjTIt6/fEIgvY6gcdOGO3XZ7lG39
oDX/FslBNoJuKrr7Zq3R7A9oXq3x0S1xZKKf2+yC4b1RMEO75xpxTKVrhdWJca/URfwfMWFUfmVJ
erswVCY+gD3n2ZPaHqiwYQaYnXKG7iWKWz8iHu/hpu+MftkjDWG8Zu/ebGd00YNValmT/v1XHpfG
1Qr6mAkPJcUDeIsQ7Y0eRg3YsU2MEGzs+0nKPbcgtS9gNuggoYR5GSgYjUqbMVAtqeVJaQ7+XIRb
4T0T2NiY6pkrsj/c299wEclbYBY82kq6gwMZsly4DvXSLJj/p8unmHoPgNSutrx/FnyqHI6YfoGW
r/ovjuYxyarMnQ0CvpVShOsHEvaw/5jY0FMS6jbRyJAd3oTgOGH2ZxaQI7OlGULweVN1CG4wmqad
ATMIi8l5+SEg80O7Fxe6/x3MGr4szYj0jeuNgpsr1waTQFp6vy5wX7/ahRSlkT0vhWcUvD0jJqpE
32+cADHsiinNsF0vXjUVSIcs3XJQTT8lFFO+/FMLWm08NAZHYAji6g2/32tIM5lm1mT71Iwd7aSH
RGfN7mDDeQ8JvCmK2nNAaXUiUZOgqIt52YfChe0sOkX3/YqUUkaGqjY2hB5XcvaNpnjEfeisbXbx
OlRISCnPtUvnZsGUJdQHSQf98cD86WEiksEyxkBk5u20Ez95ZVzpMTYAfWH2v/r0uHzOmjhm+S/y
1xY9vU0/4zbwAepSzNy/QAlOjPb1igqU07RTKWQg4ydfPrDWQjZ3H2ohVm1u0M6EuGu7P2Kj6Nlt
F8o1zrHtBG3hJ3Ma8Uy+/PA1jos4S2WieVjIAyuikmR9pleYFdFjDs3/8IKmeCYQLwOWntVLkuLL
85A9WgrchI5YbPINwxnR9k4uyewbRN/8BR3LTmFqDKhTXAJ1/uuMU77QfKdDYuFC2WRObwaLfzaj
1RgxtVvqY0OEDOE9MjK0txPjtfnqtKHVtwoco9kvCgZzKn3flw7kX3GreIimvT7g64DtjwyBmAkM
vW08ZicaPglmxyV3y3zXbvxFJsosSFb0bvEO2TJm/rfS0vUkEo8e5qvn+9ibxyq0l0w5FSzZ7r9i
D834MuiKYwzjQbNRJ1631Sngv46MX8vz6lUnZr4jM3DBGAMQyGP8l6AEvJPbwKbSfKv0XIfVkbxZ
ssBGRiPNDVJpoQgduW8Sttbog8G4GfNg47h4MdRSufiOjUGR+sqDMgThx/qSClkAAWl+ZMQ0y2ac
4X7XIOYt+4+hAFuDBDChHSEOY5w5OsgQAcEzCYaIIua8Y3w07hlxOX3IrdTmSp+jJsNdVfu0RK0r
EMgAiblCptwqKRVnxmShP5X0uH56ibJUnu02/+6Ou+HSTMf4IxJGCyCGF28Yb5nRlgZZ9iYS04J+
HTVs9pVtlsiI+4VQg5BtzO6Pv4G4fO7QCUgLK/1fkU0aTGmKpxkWMLejBCD6gQ3M2t+E3NXg+vIq
TsxRKrI+NbfgNuhfIr4/wvXZW2GVBBJabvxETrn8p//NA2ed0mOavd5IQVXONwHMF1SMrfPKqdAe
jNRokunavJ1qDbi7vNmkOX59Lo0VbDawrf+SDakhIKylDEeacsXIo1eLdeuv9tk1DUotnbRrJb8e
njSIsUPY8E20aLzgK7WBHs97TAW8Da9j6BR5ivjXdG69BBjZvRHjOmY5Cn5m92xAaPGxfAgQCmig
fF2CTXA84devJVcMYdvMTjnELHwyPBkEsnpsMpuCLgD33OQHOAmp0k0dtb3Fcq1s1yG5w+E9/qj2
caOBLjxHOPAObTxrnxDkVYvp+MoEG7pI9xw7hrbM9p0Vw3YdvOhrvaepCn7GIwkYGklj3BOypLm6
veokfwBCszthpXW03pK+OpFg3HUtPRJjMQ4rzbHV8J9IXPhO9735Aqod/rl1sGP/+VFOAHFvdezI
Q+GSzMun1X66EV1KoAEkD7+WzxkLj8pyQY4gjgBZG/88c3vJaVJjJkyKpTGMgJ6aD0Nh+OlBkVxI
xR4Wm5sJOTrrJSJd8d+HG6SRvxntENP8dKy1EuPVIvM6XjljGtXoiteuiv7XHOC3TPh7Z1GRZnIC
k/ykxrBE63wtPwBquMcDdlpnxdsWb6/PQxy89eJzdEV723JwNJFZUkj2A0XhIhnTYx2YspycPAVI
fJyA/X/odpTRgrDiSQ+yKOFwMlIxK5v32mQ/fqGvHpUxyRUCatiq/lkQev+iAN5g9hkWb6PVUM3V
BMepPPAfWAsvAqaLVyuO67ZrDEDde4JcqncArN6VJC9rMd8yQ/czRfyb9Ipdr+Yphm96wIjKkpxw
eSO1/1f2FJrZEGm3SJi04LK1GTvzGFhHosIq+8X3B/n39ATil37yn+Smk3y3PQj381kHNkY5CrlG
e3fnrCYZWXvfZELJtjWe/6M9hnEm3TpfQ4IgbS1Ie2XtWpC7DsVXnsf+M/XR8rc2+eCITjyXf/Le
MZiIhCAmAu3+rDIX70uJhPuA0txOn/DyG2ro0Xyix+Nh4pGCYwOqfc278rTTzhWSwd5NrKtUUt/u
IkFUWcyyZSEiC/KErtKXgWICynBgFnzcUiLt2yN4W3j0OTYGPr8Bng5ul+WMJhQuMrO8u6Wjy0AT
mxzM7PecWTHQnO9wzCuX5xciBN8HFLqUpT1AEcxErYjbvRpic/bChSCdDrnt1zPGr1cGvQXGxRAc
QEgTnR0+rMBX+oiD68Gg7R7Ji2rVjYTFQ4bACVn0GBg7FVLOGVxgRJFKkH5ZS54ScGigsjprVOKo
74VoalOxgRSU8liYhgAnLu/JVEUQfjvx7EXtzTIq3ZteXOQDaI3EZAuFqSLA7SBz2V3pyRgEi8Kb
YUhsmMJw722SZJSGb++ldkFEPOkdQ/Gy1WviZTPX4RhyQbxLECBOh7YAGJMhLkbhnWePMzZhRpCh
Z6nF0S09OLwUUKqEHikOgGI0IOlOjpKXA73PNs6nxZ4nqyuWyL8I4bPYqKAITGYTpBWHkZ7ildyG
PVDy7/o9VHH2K583H75+UndarDRuNEhqqbL42sCyiKK3lMLcuBSa/w+7WDwebyll6fOBMnJxAjKl
nC6eWV3nvzAhAkzSAqlN4nc3YW6C3d8H0RExWco/BRSgLAsA3KuQ2WHyNBgZ0yWMhSz3wbz11R8j
rX3joq+IWhlYN5vfpvNn9Q1AimKbr6ajl/asCYMqV3qH+pEsFbwncnASAhbGeQI2J33HPM2CHe++
6Kn4VHZuQItBKtSdp5qu6y7ITXLtilnLxdG47anpdkM4p6VKQVmcOp0TNReRywUmoT5RKS4GZN1i
Fj/fA3kUalQuwL0D62JVrkIHaKFroypZP8KWToyHGaUq6iEgL6Vgqxv82rQUWHC37YcgJM09QVdV
RGnvBoe9jY1kKJYrWiFIWLpLjZs1EH9wSCWTs3MoXQ3TDZB4depjbhaCjiiOLGYM5Om9cyNrSLm/
3iVdpLMmx96XCgLiDCVewLWix26xWaYQaQlWr1r29kgWVXMB7OaphHnE1x3WnwPX2G2BRJOWQ2TV
N0CFBg2Yf2QRMx+k7WqoXv5ghLsvsnPw9kwQxxz1B9kKICU6Wv1CZs2IgNndk2+9FZekAPrWlj8B
WaNg4l7VA0l9nasET2xkvcZqsTkimzDER8seXOJNIRSEcHSwFhrjly+zi6PWM/Zk10SNFR+6ZLFv
UE4VT3CV8tVniodVugsvIv16ieGv3QG8/KPnld2PGwEb9KoQboHlRszYorfiB7FZZQCSjHYFOglL
/GAKm8w363yhJ3XFbidaV5ZovNyS17qphEsFonh1rzbDH3XD/GWxcsdWEMUATExrpofKV3Lf/sfy
3pEX9Thf3DbgmJkEpDX6zZfLbbq6/uOzHxsV8JmmYwbkmweRq4wAlRg6Gg/J7B2oKmEuYb9n+WTM
zyyxR3HNPR44iGdo5rU6FvcfDRDArOSGAJICx1TSBkFnu8aUNUsgUSN8i/hACJwrogV3knoO1rnb
zln4Lch1VHXu1TFzOsD/Z7IFfhn+boVPRT5nYeBJZkF78CX686ImQTUsUgsINjYvG5Qkdk4oxI5c
FpFnYjfOVQ7I6q4RmaAgjZXulI5/CI+R2S3lxwKykDioTcuD1Yz9Ckq2WOjtPSU1pLwMUzWBmxQ1
JW18pc1iHij3ssMgExvpRwygV52ZyfSgvW9jWMY3DtNFVXr3/KSnHCSSIYR9f6t/Zbzt7YBgkduf
nRUYMzeCSwj0EWmtemXrLFh/amDEIBhRmLu+PattBc9vTvWbfd7cTaLpEyHM8v75kxpCXTWURODC
2Q+n1ecD3M59ZHQYOIXSWmnjDJFk+v0NWPgf/v7iLZvxYuXOVWaHvUzNwcndKAFIK2cKEfUt3Lnl
FDpVQv1p/FTgRlmH8eY9hAI+K/x3/4I3URUv0mru1EmVvOXvPscpaundRHu3ELv6/3mgjQoEKEcF
5CYJ6i5DNIWwCJTFPu2MMVhqME/VBj2EJsPyv3Ld0N5mC1bUgxoOy8+R1IOMYvVe/g/qduisxTO8
aSSunsRMhcsyD2HpZvD8FhKkxj9qVLFAHWVQdLQ4uFQ4PQN2T02WtnwtqIZElpTq8aZ5s7ZX0Rlv
gGGrv9SGyT4wuwRjjkGbn9M3FioPFpnqFZypH8CpziVU3+G/7pPcntKD4Sw2GTnEAYPRI2B4LG9M
wsTfQYO5Tov4G/3BmELBTLMI4NGhJ0x9dAjbZ6xFeOrlQTED1mxzZ2KfBKEPWsZNSoJnxX9R/VTq
hHHsKpgoSAkkPsk2Yo1QPNHj1t8E+xChdCaFM9LDiqCb/SZydJfe/cEYMkfxbxhM74cm+tWyNwx4
hRC4x03P3Z+tukDsWCgNHc0OYiSLtWpiQ5ngAOYzis0Bjf0AVh9aSlQ0c0roSQE3mkbVR0mu1+GL
mDKCfna2prMj6qyMJTn2y6Huh0Xw/YITTgtxKDIFaVb6waZerlkPsNW0ct0+jUmWiLr/o5ERpxx1
5taRojzvGXRIDsZwMfNoVJ0Ort+VtU2BWN+NalqRzMZJuMRPleSe7z7viEU141Q9D6DM8AA+rvpA
fmu8yP3XzMLxIrsxElDr2lYlou7EvRHMlzquGoZiqqW866+Icp7c+dZMowDYZ4PfQATEO0D/b9Pv
79HL4eL7Hx1BgUFWACrvqYc6XX4oV1HlyNkRxAmkN6edIOfY3ROj/nYyc3wEc7mR9q74Q1yN4FM+
aPiikcZD+4zgWGTCSQfibalDFzDkHrn6xH3M4eSqoO5N3zNXLoIOCeaSg677rAUJQ0Ncs448wzkL
ajpoN7QFdD9iYS660NA40HgRJZ80L1CDkcosNQ47VZRxdX5OcSbjOtp80tkxPY8OBUdgYzOTeYG/
9V3DU1AOJGbs2yI9Dot0Xk1vWikXqxDhnblUupWxW6Tqir6WuknEhU1x0c9F+cqbjqGwfU/BL4xv
ZQh9iEZIaS5VGJAtbU1MAUiriiz3oxe/7O8+vkLfp3mjLoysunmctIXEJLnyrqXRnZWIu0YZRgCR
vu25GQOUkUhf/jbgKei5w3Zn3Aa3c/E8sxj34CIttwoaY9rRPVqLtCTaXJHx9rMr3lE4shY5lMXW
0xEb9Ju6GXvc+MRca1bIP/zT3qP2eZcxvK3sVmfncpU6vfU0Zt1kqe66srhMThHGQWvwH3KHJfiG
Sf5e5rN4MIkj3NgUSVq42fmOthFvgUa6cw8q6SkoxAlfHIBgE8h5At4l6gm04hv/6xqw977eXr0H
ngnVCmAvmcMcpcJ3t/OxaoSyGwORSfqfAhgjXknAZSX+Toa9S6lB6xqL5pbXhh5k0RRPCfVAZ8yP
eGcLByq1sbyPRYB/G6XN43XrXqze0ikz3B068YY2V1oukCnkebEvxLyMKxsnXbu/tf1X64YPtgnS
V2EH+LIWiZnWQHs4ZESxfI2noXQjtxjoTvXb+msh29YCo3VXbe0RskCXMoPBjvLMvtmduAqvC6tI
aSYxrNwrBep5HIOX1uogv83qWh8ILAqaMlgX4r8tiUA4xCs5wQyGxtTjhb3yMlgz8LPmBbKQeLkg
JalCgoLWilf1xSNPN/WhnL/bhI2g+kYpgk+zrEfQg9XwH9Keivo9UySXCGktmnyOPGu+8rFugk9K
a0t4SwfxDWwDuIwv6k1nbjbgQyUUkHeh8yCWkixOLb/H0m/Q9l8H55LRIYiuTOGQ6RLToWMRLy+k
e7ENF7r8BeqMB7bfns5m0w2bDhBS8dHL8OBjdPYP5o/BjMjwVms8bY/rErpOU9ShYdpZoz1JCHr6
g3+4VZtsvXplks519WmTIXO1xFz8QjfI6rVBAxo0SBTx1kJAPnkOORrYZnAhF3EsRfyYDiU0M3FA
XDTSPqME7F3H2/P0/HAbf21qD274aSfacC+pasxNGle8QmQ/WZA4QpHYZimC0By1Jvw0kNTWKIdP
cTp2V2INcoTvF2b93rO1dcLa/7MoF0684KGjXLQB12d6vKP3Vr9rbE9/KuHXJb6R413nEDkE7dCw
Cbw53ecxuteJqi5vL3WO/dLI+fiM5TN5wNhsUHbzU1zk2CNAec5qdELJh8alH3oav9wGnomkTyeJ
LKjypeLpHm6EUoZyBovayOXDFKfq1XfGbWHdr8A5TLGKaCVAdxd0V0hES8btUdUGUEwjldYpArkr
Ie19AdQPPDLDtUnbX0eUwDXdy3CTisVvgYmZGletrbdmhik5pMNzaTMg/GH2euK9vcUg0EZt87E1
y+QATVyYvsTfxAG7OspgLnbqVqRtVCbGnbnM65EGmFBFcwukTN63fhClnhPjT7MMCHy2CN2YKPdi
NMLqv4QpZclkhNKez+mXBE5qrI5mf6xbvUwl+g3Fq9s8hY3+mzzkogPqIMpvx9MVDdXWgEcpQGTE
V1uuMANyB2Q+VAqDBuknf7hgpWFcGzykOJ79Xv3wmQfibgDNP+NC/aW8OToRXrrNz1lgDAZJkxZ2
ona7Uj1i4Ixzk/0JOej20m+GzDZmVZ3xBMsWUs1i30ku5xOHGk8zoXHjopAHTwfXYJPToTPAxeTH
UasVPrZlL7RtqhGu/jCxxr8VV8MfeT5ddrQhJ8ntvUMCNosYqhsnmd+Wqrn83w15fCalPwbrx5T+
NtqX+EHltji1IkrImI+H7a3Pbj7fgy/Zs3NUD0wDxiXQL3h8RB+H4Xmo+0Cwe2yaQ7/uiK0GsO+J
sT7oqrPZ1xgYZJ26q7RNx8p7At7zBdxeni1SnT5/2y/LRmfSRQuP/tr8IKe9xLIRPj0LkiTFseM0
KL9KhxzKD8hUhPZilH6yndmg99AqRtukgXlJwnVBUb2VObUcb3kzR5to/ImEfWLFWobsliEzxDvv
ufFihD9953SgLkI6v15aBBgs8GT6p99x2pv1GeP4EGogdic9PYHX8E+zPC2+BY6nqVoLzRQBkntZ
urAxwDIX9ptoSaorYhhWTUCxMxozJxfScl2u86QAC48Gv6abpawv4Hojmm5DSKVxoo9KLzywcWby
fZFZ83oBCImxDsszsjvZzqDX5MnTtPOTetAJ8LUChpUKYQjwboUucP+Iq37R66X7TlVMFtsDPZF0
jyix53NVr/aOrJs1G8tbjHS8hBYMxa7hUK9HcYHtiHNrdRWwfPeJ40uSn/NR4PUyzL5dxMqYU9AC
1Z81lnmhE8BUNr5WbDt5VlhMHyMcmXirNGJhK1kNQGGy+rYMIJ/Sw/wAMZ4qMV08BH9H3dv6Xtwx
BPU86++Ii3/SDbtIKvz331zvh9FprFk/MU5jt058Y6u/2GygXQYAakdT5nk8T2Xbq7w2HXvKysS0
ybVHlfzPTHMshQbVNBZeW0tuztTFDsBBH+mU6efaUO27uSeTjtzsj0MbUSjm/w6GvXdg9NoublNM
U7bYDmY0ygg/+OUerD2bi7hnAI06OpqOafcDr4n3vH0FE9nFhFr1tMRl9SzfrxfBBcCgMfarm4SC
En733UWMtVKxF62JcZPDulO0DeavCfBkH+Fl7QXMduEvgE/6sgweNSC6p3XyREvul+2TgWt7ZwHy
Ulo1ebYvCrAcL+8L5xg7nS7zA7FlTBxUZx4C+yxPHWgR5bTvvzlqBIEHspe5C88SYjkwbIJ/1eY5
TWg7fzieI3EvY5jYpamLU9w8W6ZrdiJuouhMWTjH3uP81wkwhVtP687pHkck5aIPWlo+I6psbTlC
dgJVRrtQNq+OaBAueRyvZMv2zKzHj+S3vNibIkwor21Fx5HXQn7Ebp8AFs3LfZeS4FTh6cYCb1nq
vPjpqpzFr9X2hNEpl3Git/ndk9ub/843sdKkCqz9s1iwJHgS7Z40soY50cRxgaHD6PJHItkZjZNE
K1wd7S1GfG6uL+gfVEekPubbcsvUudgMNwHfYzX5YzFo1NgHzYFGHuwmW5YHTs4vKUCkwB7iCEKP
OKtf0IxKm6/W+VrXRWIzwgT4PjMrO0xS2V1+xbgh1F0QIuE0SomXwwkWS+tVWCP1xZTEVie3JQ/f
GD1j2LtJc1hxYnUpgLYWDd0puok+3Us6FSgYo/WrOPp12JbyUB33LGXiJt6wz0Yp1zt4Y/LsOj/H
tuV3cqoG5r6Bjih0daIhHrdnAgvrNS+pvRXpfILjnAL5VWk5DsegXEaZMOkzSW+Ug3iK3y6CHzrw
f24+qQarejiQarAMXUAr3Vrmn2vjDBRQyWhyl6NN7KBPx5hqkuVGActV8EE0bGHId6SPI1lo+hdt
x55OUWbGIepu/Geus7izcP3/12j5hRdcd3IKUAREvbyEVYnQzGVBhXHuEVT8fgoMT5kPRcBCDsHw
QHrjUtRwVvFqMVyr6L/OOU0iuu7kf+mnI/KzavWOCNYX2OvRGFHyDBRUfR6/5ctAx94VG7eyNDnV
iIQznRQ+BXorHILysIrjvYmxOsWyz2sxzLRlAHPUJnQXWMBxTStAHjSMWWudllDyzBuzmKR349WQ
0rGYs7Os3vyn6EwxNziubz4c+6dkdR68o71aDEqh63fQL78FAHguRYW/TJl7u0Tfsa2wODObBI/L
Dopda5r3BnUI61utgBtcULj0bEgt4Nb6ZpKMGocCC7zSw0Su8Ts9wNOQ6bGPJvJhaVgvTczAaOFd
dggzI6UPNHPFSsvrRfQlgt6mhnhAkzHF7GwQUyN1+Vc9xEKF3fjttnsffyM+v+P8GRBFCYnpCrgs
tH6STyfZjvDmG3Xc0XawAEWxZcLy0Css1gANzdepkZF07iinpb7sz2cBvucIhPTV5gKEvVRpbV0i
RyMxqlCZRtrUoPZgjg0HakD+tNKi6C5IGEgeTjO32F8oiLoXA86TmuHMlrLSumUj7camQ+NLb1QP
WQnjPnZm9qUDpBcVEQc3OVkJzsKN0QcL5JU6iZv0Ux4XgpDVdk3dxITPYYhsaxeyAeDjQZH7ZvYh
5Wx5VLSDXR6EqM9hbaMU3lx5ZcSBqhpeU17MdT9teyDCQZUPx6t6XC/PCu7J/4zQBertzYlnyUQA
11SjdtHMQbA0ncM1f72Nm56v5/7TPuxb5lIC86acO0ncJMf7+PND2JSwC+zBkd2gvqLQVCAAITva
WHvgDMOf9k7Eg0hGkN57iyEXOUnJmsFnCtKduvTrbahQXO2xlVliWYES3pkI1ZQWa4ORUfAtxMJX
Q89+kx2kB8vSEw8E25J1bHbIjjNhebQ3vGyF9mdx97v5uJ5ve5K0op6GzYt8Oo9sSzeIkmn2cRpp
WRXPTU8DiN+EFkv15Kk643XRdFw2j8w/mfCtDyCDzUtDTilWYc3vhY91Jbo4+IetxnSIohDoti+d
Uaz/FTgYVm+NNEP1+DFLPVANdX7HX4b30gs5iRZwxJNucPr+D3K3pHF5U6QylUBu8hLachE/IHik
1MTQzTejYIf5xbK4HpDKgNVw9oyiAqMfY+cYtHasFvBvdkD14SnxTpIpxINc5NCcs5kC10kyBhPc
IeefX0dx+M5IKwAr78FodmV98GT/aeK95Fm+mPapMU9V4D42Db1usaNXQlU82ETtEuEBYKSoMfBx
3Pi8vna57AEbp/UcZWYK1mTxbXiCgW5jBAyy7TTcOgc0V5kwWUs5ei9Xo81/4aj5dwUIF4MkmNRu
+z45aXGf3aOFhFI+2wC8/Yg/PVPFSfPMZvlxRAjvZbxdozaONyDppNU9YSskcH67j1DfHKuKXkVE
jyDk7eGlIe259ntmpfvemm/DGILMjheB/H/Ophrus7wCzxLqCpTwqCi4jp/S997Awf2dBYvNPKyb
T80hwjpyIgMC8AllmKzHT24wqOvWuWoNbVHqljIFiRFSJGQt2pysAe6gRjzmre7v5qAAv7ba2CKy
2zIWzo40bNRJ2ZOE1B8Wv/dMiNHqu9VGTLpWfm1JcFFxvWYsnwJhhFnXHpHyr4aBZOj3aXcpKrp0
cLlC6r5VHgemIzOBajkix/qBbINVz2Lcc2nPbIQ2MniX8RSvzybyzjq/9uO7nRXz4Muw9VK6hqXr
8zK+gLNoHumUMOfBbipTrKZrFibLlGozdxILjGraSoPgFFgMEVGuAnTfQQuodhS7yVWUXep9+tkv
4FJL5hfhAnW4BF33fVnmsVVLrkxabUoDPHpyauvLnoQUf7vBejDmRpDTUrk2XEWX8B085XmNC5bF
aZf+S1H7J6CeHoVvPxwdQpduEu1O2ja4CnhOs5YF+ziXad8am/3yVm11z91SzP7g6fb7ISDZWij7
ZaCqF3FMW34NDhAdzjMBTv3eiPr6Qc4e6gdJqYDrSNNuM1Hiw1Cxhvhd/KWLZFc2hIrx6dPXCIXG
6FdkgX+uy7WwFaWU4z5AVNNTdWd4DqywnsKf9KVhBgFmi9euLOmt6SQVxDEmd9ORYJoizFTgfrbC
GcPHqkYuc9flJHHoLam8vGd8yMGJqiMT8w1dgpdTbo72fGg6fLnR31gox94Do2lR6vWLXJG/xqJ7
YK2Rhd1uWQRl2oASgUGhuqhR7QiZMv4Zw5+KFBAxcYg/wckqDlhXEsRHva6Q12OTcdqGTTQ1a7u9
dcRAQNuLVRAc8mSVTyYLmyeDr+6nKwEKzSbS2EkgxUl3HcE9zyqCUWBdI8ng9gMb5iuaTbUzdOHx
/+ZQD+5akqgJD6FF7KvSqMC05Yo8Ju80N8Au6zYhXM2hPnknvsJ1g+CHUvGFN7JIfr8Dt7poAAIS
cv0cX5yC3gZmE45ravFnQZGDdjXT7LVQ2O7cNpa5osj4dBAXnkmiSndCfCJuBOPx2ahmSDLVzb4Z
TTgKofGIIU7+y/j/wPpaW9KUrpCcddvz5A/OXVgaqfUePo/A7jXN6//JyBujOpvqZKYFK60Hh2Yn
TKdBY1GqK1ZALOqroHzyPmUcORpw3i+9ilD/YKngT7n4TaVRO/ATQAfOKVWC56F26v/ep6Ck1Zsd
BsvJkcbU8obwnJAUp/u5cVDGC2GzQRPpam5mAm/GijKmBQo63mNX3pjZhDriI//O+N2K3pNeovX+
ZEwiGc5ACjCiTIZ5R4izbzPCIm/o2kBuV+F+23IcCyGv7SIIQqXZ9P2NRlmwjrcYyLjkC8SsAhWJ
Cw5ThQWR652bW0rYlmGsBX+vCzQsIEwWWdesuiSkrWjdGYRJi9Zh3ZfDSU7Q2lgAP13xJ8EsOOiu
IX7HAeD6HHTZ1Ws9P9z5QTyXSiuv64DkjHNxxHDY5Aitf8mccWOAY63YbXT84OhQhwopxeo1xCnu
diJb5SEhcfhfMgnkBKGNilO4yOVnuxkGaMwHfKjID14BbWXmDefDYL/htsz1gbBbzPPHwhd7tXM7
0qGnVtPbL/p9V3pGADLem4/ZmwkpWIXN+jpKQCBpUTsjQfFErGDh0Ti0ZX3xy5R0hDaMmpCLAv0G
WyjUUkUyzzs03oNqhHlL2+p+JQ0fEUix3fUQCYu7eZ7C+Sqa8ziCG3cUiPWkd5JW106SJPJeogVa
4Q9NNb7bK7SMxmEe/GKlxS4cEzDiFBqG+eTiHHVBm5d7/2JlFEp5wPahLyMmtl88AzRkHjLUSR3g
znMEEz33KcYeH+v1qBDQERj0E5EUE7rYVR6SZBll/ycEbLadBnwQubqUwT08M4V5pZMT96gB6orB
YRtJv7YAs0F5hM3YNFFh2kovP6IkjX4SxVtZ5ZfIsFQWR1rB4rerZg/55aZE7gVLNpt62UCJ1A6O
XNwSPUtya21TFD2VgANKVy/VkeGyR+5DKNdKCqpt5x20mfGSUSvOGhmuX3NhM5+bpuu8nlr/cMNu
wO4ADrWW1NDf/bKqnikKxRJn7z0G+bFuOyrwvToopODUHUGvWSUCispKC6mHFraBRH+vgXjkFaB1
7L6wHf7vpZFWV51Xesuh3obSDu/WzTCFiBH8aPR6U77+U1i7v5v/Io5E2bBGeCOjRSjhApA26yTV
V7x+PpyVAaBtTMISVeSpVcS9E6aRn85CHuy+vtaPjlRUkNiD/X39tVkjZNaVqxvBptx5N8gOq69m
a40RdkxeqlJj1XV1Z936T75AO56aZB9HgTNsVZduN0QAxzMdUwKg7qFtnBRDT7+q+Fn9r3H4tZXv
KdPjOkT6jViZ272QVFDlKrU/h/bQDqfDLOIuoBp1OaK6XBq+pKt14GcfNkHRWJN7LeSIMoai+wks
wjy7v7MLBQtiDa7KnG2eqCrIeb3oYdmj9p9nisj8+HM5j5+dIMy0vvjc4BKEZy6N6NOqFgHh7AsM
hjss+++XVEZhfFKWJVhB/2RclZH6+JqF6WE3WsImFl27fwZmzwJ3PqNe20bVMe1PpERjKjDBObDg
119+6rDwIi2P/JYaEZ8sGneC7BenJIXuCgYPygoqR96+B2yIq35RMOAjWA6GIH0BkCqYC9TtdeSv
T+eVGxXPxuiCmuYMUOO7Jf7JTTkRBrmy2Jj6aUupMAPIOCSnH2Tn6cvtZhXeI6amd4uI+9ni0w0a
sgxzK6IG1clwEVGIASXyBR4ynf7T+vnL4pJJuPqduuJHDl3OBM2g57Y5U9teKjuFXUNqQeq7GOxx
EwxTwlCCnASV7RlU1OAfuTQ3vSZJFV/QJaaarFVW2H3kHqQF1y3rfjUSbp7R6bs7FqfCOQGWa5Kz
wdKDYieYAM7PA01rPGAa0EuA4ZXHDo/HNItAgHkEnDX3hZR1NzwYPy+R06+/w+yNFJ0ucnuYo1Vv
IT4jzn2DeKn7c+LHGCmCxss5Ym9rOcg4Pvc4s1sKWj9A/A4s8gWc9md4z5tdTMkQksvBfDkcj+VY
yytTcbW7LDEO7f4V2Cyp6b+M8xsJ2gPb0mbhkcwr03eibojUOLXD3lvjZE8yN4/bn4skwqgcpgL8
GRfRt7puUo0AQFqFeGUhb6uLbn5i0Njy5tmI/ZIu3c4NGooLLJptowXyWnLb+cY8ttdygpXW6xp8
EdS3nSo5Jc60oe3mXMHsOaSJZmuwqzn/Q5P+H4jZAWEo9sMbLYw2eDCW5SibiKW7y545CS/OUI7y
b1CcBSDHf5WawYYLsgXDFkVxH/jEwOk+P1VdYUZHzeeMzG+ca/9lmAYbvjMYvC1WvsPj48bT5pzt
2gfcmLpLdid4j65cz6IibuDAA7WLqM5sPDMYKI7gVjk80msxY94jHfYvbdAsJefEf3Usl9ntdVwo
RcT5aYxxpxImX95KykmY8Epm0wGz6vvYjujiqXj4H13vsRENesFmrAt8xTXlu+9haZtPonigS7/b
K6dl76bFMlvCqt1pUKKXHy7Jyi2eMxIlv7VgXwYjnO+amJH3HkglOLG6NkGzaUxUNMjMGW9IiuaR
IXFPllbO0TbVxpid+2WWRL3/ftnxs0arISOUGwS8CPBrlWvXdLdimMreGHYmMF1+0cxZeSQc/vou
jcyYdglARIfWaQgkUSWOe1cL+HVBLS9g9o36UnMA35MYuKdZVhfJFq9ROlQLIlLqeKvOWeHnFOid
IXFzyXvS5H/Jq1SuH0qX12u8wYpvM67jUYFvv+u15jUs0OoNmh8WrWymepa4P/9CR1TRcT9fov8w
j6dB0hlY79QP1p+WM5bidm4CJidkAfuFV3wNy2EltmBYgOiqvPVQb4AQd93x5WB6sh6GLKnDDLaD
H1dX5/UAAhxW1F8E0DIN6MarC0HOeqyNKVTve39X4EztXMCqoJGgmr9DCH8Qx8tRMmRrFrmnu8Dp
KVToeqNkJZT3wzwpeD/4E5QiOe+5Bz662UJLBrPTST6C+HxTC0PrTB6fUZZKrz73sl/YzEX+yga1
wNW69Y8f/JBprt1w+7ZuaOlAf+1m1FRVWIByKlzIfpbw4a7ZSDxGESUPNOT0vDLi40Fu/OzyfSkq
yVz06UFZm14x51xbUtsiMoSUPq4EBfBMJTBvLEVEH94x7/ZCmg/TE7IWRZZdodIMWPv6pjNxzQCM
YhCPtkJxXM09F2hFIRhj6hruH+/PV2DoCKtS/UxbueE3DG96Q84se9TtxuJH9pB6lXGN8zPeirs+
hscMYjVDZ/f/zBnDrqYlHrjOPZxaAYmMJTa9WN3P/D59MOk/RkLeJ5dpYbWmyJS13Nb2MV1DRqQe
A87bsZ/1Oqh7BrNEU0gGG91YnoEbkyZ9D3Gx0qPWPAkiLR85FsKmEhUuWbNjjX/UE9gMKKliy/0W
xrnKis+LfA0clrTRonKn9hog5fdb/bQnKT7qoYDBUuxcH1JCRl3s1i4vSGMvGmHYVDLs14fRGTlb
kVCi3/r4RAkNW9SsnhVPcx3cFQ639SQtuKlrMTjx645+IGfZzmpmD4+vY2LviX54oTkFpA9o6nmE
VqaDQ9LKd+wQrR+9mJrZ0BwziZ3+yaVhuFqngK512Tygb7ue5Mzy5RzHL4Q9tjmCt5Tshtjm+Y0p
4dqJGShMWEDmpbaBeQQiAFZes8Gx6N82dqfm1Q7TNtyYmNSByD7TjPe6vForpDuknd1ZiQJgMs+S
ZM+zkZCfz0T3lmd7FzhkF4Y0RlSS7f5c8L7Mrz6eLUVGDYVJjIVcyrGfZipvIcKt8626LI5OhFSG
i/C4kjEvE0vlCfRPiMZBjN0CMLRQ9X7VH+Qw0vu2fXjA1staxmZmztDZ7ImmV2Ie0kIaEMhldsUg
TGPZMyzq8SOQW70QEpILYVgw7pwnigfv/hgLvCgMgpAQ1Xzn9cgFD2880df3sEoKuHptwpxnWNnW
fxnQecoxGG/uF3V7pt9UZbpoNGo7auZUWDk6qTvBWKeMMBhXtY/FS6lvCDTavmx+3D0mRNgLFTkl
jCznq/tD22IzURLuw8IQSuwv/xeZBjDPrWlmRgu6ipaSz+D8cS7wYl0CwAQETHrAujFhRrbX+Azh
HkjK2YYyut/98lHpa1ZmJottoTqVwfbZ+9bvzNPN0R8DE5my/tp9o4LwvyqxPFrvpaKC+fsVr6Os
wnuzVXJuA33sNAp2dYHFPKEFTQd19w77Gr4hwyG/8Ojm2Uw5BPvP8NZ/MjlQvYxmHq8KMxJCHON6
m79gqHTt1NRduVTPBE5MuhhviLHA4Vy5zW+jzBnHDMu9Vd7DKVMlGU6wchykmKXXZ8v++3jS2nuv
BM7MQVedBHpJPNIdGT97S3AkAwoWLliPf0z8ArIlTpUgvEHPupln+lOP2NB2oMoxrY5+5Fovvyxk
G344CI95E1NIV3/FA8+Kj/wgMkiBw2bhczIvA7Qdqag6TP6xM02HfOPlZ2P1fNSEBndz6iCWJNz5
yd6YnPSmSwPAijfe/P6phd7JpdMLZmN6hMqMFX7O0f1v4rAiapS3CBtL3B+bw/wQeBBCYn77Qpbw
Y1sQ70k1lKV7RTodTaCMCFneejRDeMMYMcDiNESEqzWSwdhyMvYi0vLcgaQbmZQ9rqOOe6Fhep/X
68jfO902wQsDq/C/UXeD/ow/FoJnanYrrMtOWSkvR0gFt23su7PsYccBs6SwCpnFA8x6pzI7SzC5
+cEmi1Abok2kZmx7nVl6RhBVFYiouk4dEmzghNqtMs2PyIxJzI4Bjc+BdGwy4SHy9B3/kWlnRLIu
XqUpnjp/6wN5W978gmTzD0iA4gyZqdULbkPeljYiokbNs+y+H/O72f/l83Fp20mjo9uoddmxhq/8
ym/JZtdj5P3iMSHA46HaHmEA0bLqtsbHTrU4i56O/5cxdiy4xgRminnI1Vj18E2OxQRCnffk9gNk
tqULBVCbb9j8fEcSUeAw3hyFiJYR3lq8gGf594ZUZEVFpai7+EdQjE4Zfe5YtxBFVeBVCQlQfhqh
yaMhyGb93+eBv9siaE8JJxim0fNAsbO+QB2Pr4IlX9+SiVA7rH7BdKmPXL3u4WV85AS5eUkJ/QvH
i+gtOQpe0/4PIFAXsTvap3pQEPsJOyhMipgSznW0IhPXvWnclIAf3BA+R1XJ9pfVoYdnI8ydzMQ0
6TsmOOMhuQz842iSgbcyaCNQILOe1Z7lJZT9uB5jyBwYPVN/uryFHwlnFbvMHaGK40Bv81L0//u6
NEQfCTEh68dh/w99sV4K/2S4VqCwrVRoAyuw5vOBA2/bpjcuENfd+27swp0yIIdVI0alR6FY5HTL
SbryPWlXoJI+yKUSoNDH1UUsKyjrSbo6xLmHCpExHNroho3t/3MTlNnnMiXSHTr+RlPmFC87JCNj
I/QQTii9zkyRggkV9LojmlJbhRPjxjj8ldFKzlhHWiZH6xSFk9FLLdfiZuLK9YrtAd6WpAWbAz0t
H02urSTcBwjcIA0u7XyYNV+j+xOe24qn5ZMjD88Ar367Ra8JGxJSnrlX8mJmLl6E2KjISdxBIVAb
r79R+QcUdrkd0ErdPQew8DcS8g4Q/21Flx49K2tMbr81eGVUC+pE710z7JiUD8pI8zIAmrlNjbM2
QgxhPJK+vfSF4UkOTPKKRvaKGXtcuVt2IdSBbfVeqvqMEivXdZpUKQL2rjhHFiwivZ36TdtQlL+z
mKPO4OyuV4iutdOyszIhtjClRSuofDVz2/sGI0eN0VYI6yfbHZ2PNj7lUoud5uo89nl3Jr2WjSl+
HV0Yz+Dp6yPxfdtu2YfO9z21Z+xJAfZkZYNzkr0WHO17xGHVG+BHcu3qg7ZqbTh9exW9eYo4VgKn
2MK8Eg2saUiqqYn93RZl3KjwQCtAKJv/3YB/iy4GHEg290NZJDJjLeTQjdUYbjJmpmKFOLozbs8Y
dbqByA9vl6kzc2rG9mxxCJKJUI52xPAi5UVaC7N0bgiFJk/3WXCDw+Ouvdhsgg3XK6ylPYO43sc+
cWkpu4/a9w3eVGEHRA60ts09KI9312ka//zJJO5vecLH6hvxAePbJmIdddwyPDW2JJpDiozkWDHd
oqBIcRvXd7zyPnNWUftDxj34zce7rC0EjqiyCw1ZDyZn1iwSGjNNpmRxH2bUiqk+PHSDjdcctliz
mHHwewXbu7YGlxQTmZeZIudc2UxPsndjdQJzfp/KFsmTtcH/0oTHW0S4xzJs7OogNQtMImeA64ko
WOWpWrYokatGZ5GKvY/aoTmAzgNp2hnK9ZlXe1B7vxehGtzO+5WXU4E2nHzp6dMfisg9jiYixL0u
9qI30bVcHvDZ+U5Hl3/2b7dXDYD6DnCDOsHvfGp2TNg0dDgtJDxWP4Yp4y0Ms1DgS179lw/e2xM3
BGfsH32WnPn90Uwsdo6dc44YPeNfuo+b7Sy1EiQclrqKRI/uU1GBx6+nYROflR2wbbY1fP+mp0Yk
gac+mEznMkIZoxjmVWcGSmEPFwM/fJI2KaCt9h9KZ6y7fbp9TCDXhUMlPzMWGQ/LY+nyr0sfRvlQ
PG8BLtYgfjcnaVlRy6kY9rs3rbhOgr0urcupA8W9uYVQaTra9seP67Ri5SBG5GWvtllvIDQw4UMq
2fTNDTsyKcAxWiWvHiWGbFOxlJQ+eBOgkLXKMX9Hp3jv2CXdzv3dkCR44UdfebENJfEjA0Y9vVAM
Ms0d4nRl27g7/LuhC8QKVlEo+8+XjbUFUssZjGtv0xOdYuwDuV0Jo+W1GKQpA9ueEoPXNtIaCsjC
XWKBhdQemcTWDd9sGjrmzMBvKy2hx+zc2888yT9JjVmjEud3sJj4ocejCm7kZxlMjDAr0Gy34lKd
41lTHYG1XYkgXskD895gPY33xn96oCPtla7/iGbdfsoV66y59df8hVSRlvp16vsuZl8Gv+VOPcQ3
tEcl3NN7UeLsv9yb0jxhykAN51mUNJZbLfUDLsP2YESp84lRwdk6fgznzS64Xl4rKpa0UDFu7C5q
TMarDSsfTb3prkaZAwekTJW1FjGelWpiza9ygaEbEAf4bllHWCgRR4y+GYPKUIsS3Xb0y5pJDDB6
4vVUzMbm169MGMDzuTSb1hmaIuxHBTmX6I7W7BVhC4kMIrajD0WH0yWbyjHwGClFzrQha4XlfReC
6TUb0wLrTcoJHCidHHNqJXdvXBCdQ6hRWULjfrwx2tfdVULKRJEbajObMF2/SiPji9bfh2Vj5OEa
ONo6rntanzlL8lMCPAVeEIW8+Z/MldyUJVaq+2OrwC76pm+YUQcogxWiFN+V6CwGXzkF2wtPHpDs
hdQ3cYW7aL5v2l4Yd+fS6P+BEYYFW4dn9ih3m60yq8sDLKykPEI1ST6+bUWb1MTpRb5p7qXg2wAI
1EQM7PlWOpiOQO5SJk/VEfIHnAizvmgamL6P7Mj0ffplur2v3q7/MFp8FtTO6O66+XQgesucnbg7
QKVMoTkGsGp4pxAWPj0IbQoCWTR4SCXPFSY/2QDBHvETY6l9Wb9U/qr6xM1EgcC1v4iy6+6sYemA
FqRyAenL0fbu+wstW98Xsn0yNWFTwNfIkLgm3+PIWS5XOiLqDRAVOTUqeEIabDKLahmIEUOcedCR
puRY2+bMjjIcjnLPQiiwpFxxZXf5bYhKnUaTXUQTMyKTLEC1FzmDq6aDLTMMzkT87Hafsw7Why8H
D9BeZuYJXSgzK/uQrZ3szFpdMFzfMrJXbEUT0Z1zgnJeig55VOY31ZRnUbmjdsO/Cp1cu/jOWRFD
gGE9J5oue0N9msL6YO4JHvTyNLRt7nEy5kuPZ8Ye2CvfshJhysELF+B8R8oJPPDu17BCa0KfiGrj
447+PtAjMk+0cC84wHBTm8A0es9bRhmOA/vraYGWFsCY4LHkAz83JBjVm3VZD0eao3MDYisMFvip
KaG3kcAkvql6IPFWViwomSZDX6qMXCFIxymhwx5KHPJTbhE7oX884foJtlz8VOxenMO4sAQceN5z
Czxz90MBLjcORKV7lWcINHRgW8fmag6mNP3NzQa5vac+pvrtKCFLTDWOSp4VY5VajATJMP+/pLJD
hMjxTQC9WXR3AFePJYnKBVGvS+t0yJqWwLu19JgFeR/qQc9kvknCoDpmQtIxupnpwWHPTkBGZ+tA
PbKjxTO6c0WeHAipzsDEkWLlU2c+w/v2oagyDFWtXoyIQ9XkB6YBahcFRYiioGcB4axRRdeUqWfA
ISo40fwrQONKYUDrBeJZzib4G5lcdeLyM0roFnt9vphSy1RAIYTeQV0yQ7jiMcdlvvBFunAvn89U
9uCr9ZDbJKaxrW8Gpq46hHAbK9lzTFbyYodVQdNFdj0Qzm8BNZnXjq7UcxAKfgSrNsoP/WKgiWdm
tw+QgI0beHSiGSqM0s1Bo0um3Km6sOjqapSSOIT0OwB7dRyYm8LQ1dGuN/7yRF0M427byG7xl8AF
bv1Pc6G9v7ZD6dqR8ZOjdzb6xzUkX9rIpHlw/NxD6/YOuLWNQJo7ymqab7SrDlzbaCkp7VgTKBsY
tanN8Ej3DCAGllive+JrKGJsP3HoHk5fWKbPwmaXroMQ8umQU1xMhKI/0IO5L/A/vlCfqaGh5SA4
Qc4pE6nsc27aVAFnw/EAmmCcNevTm44acaByGyBwPW42GtVXMvg3rxdEFkckpijiF3np15adNwCD
rsycuIDHUGRircxXO1hECe4zPljOnE11o3IYM3nSsM8iGVH1yRwVgNr4A0v9u0qMD3KFO/lZ7X/0
f55wHrxhOAZx8Dxbn6vc4l3aiQZCUbtGXqeu7x+X0h1+kZk6kJBY9iVb3PxrBqUrKBzQYBGL33QA
GCshONDFKajTXUXGUTbUOkG6Bwg8B/Q1R0jEYV5eLJg3m/UG+nt7VGnLKwKjvRs7oC0Fa6ZaOP/0
bG9B60WxRtWtg6A6/JJAbF7eZFLOz+gvqMvVlmeoalXk78q8s0JlOxQGULI7cvlvp9AlxanNN/Ku
RdU27v/V1mW9sKrsZ7mPYPf/cjVlb3Xb5lt7EZPxCHnGYTZFGBrSYkl0/4yUaECrSrzSlzAccYR7
Gqkg6W7y119EMkJyr5+k3iKc6KGb7HIE0kH6GZRFIMXBStuzO4jIqjX+tiXCQrLxelNP5XvQoNCm
Jh2O+w5JKhkJfBXr1IWONuX4b3rQGglulUhgT432vVbkIgAvS+2rlQjitqYuox8hZ5X4K/bl/yqU
fSXjwL79jNU47f9A40zW3icIDj+96uUMp14g5Ger1ZdIyF2/WwTKvJypOa74p3zWB3TeHMmjS0h+
mHVJR+GGguMnVlzQEKqa4vhdRPQs2E7hrtL3c/eyvvMk5vKcnPdOUiy+J+I86Oyaeg6PlKriVnVB
+j72uvYqSZ+4JOZJlbXFf9YlGLRhj3IdX3ddA+JGqgdxddPceoX1YGtwMn31QS8KUxzPp2y+PhKB
3ZxNg8jeraHMdDdWNUg8pZiUzm7+wZgAdyKRLBzi5zLVerJ7lKNWXXcTxjSiS725T/UunSiXpn3C
sfWqfmsSbjCR3VJPnhVe5i+hVYi+JUk8KswX9UpYCRpvU+VGy9+h53krxpU9t2mfWYgRD/AIFMfJ
lWRz6jSziqrqMQESn7TJIyNIwO2VOjZEzBZYaVa1HjmLOlMQzGcFo4xOaXRYLoqs/H0IqgBt3bPH
0gSGvg+pOm6zhZRGwTOgdH45Nr1xG5NHSPwvbBM7J59BWEkUk5ooTTG1AYe7t8g9+LoW4exAoEsk
3x6eNPvbK1QJsJ0TaFWiEqkjgqfkLfok7HqRegVfqtInPcaow+Xy+BgVx/IL6KYFFK702p/TSY9n
B9oKdsLHCYLPNP9BZyNSh/f/MetELtGQo4UNV3UOn3Jaztc01EuGB++8/GkrrNM/RaVGAjJ5lI8D
0bANGreN8TIqSUVISR0M5bWSGWNaMho9Arvt1u/yPaiiqNc+Guwg4MLjOFfAE7hv6giyas+rNEkz
SU8Jhb6jvB9UqdzCzdER87HmZ6Jme8o2fQCxzCj4EslkE+VM+FGop/nXdRR7yOxRjhrdi3BShXAq
Uo4MORooxW747rPWnkyFonUpGPlptOBijF6U8UfIj4xKGmnm1CjSkLR0+oG5EoaeWj9U+wt4B81p
OinngYQ7fCMzaxMol6EldIPamIoUGOlfn1dAuRQTAiAcXRSIVbB/dZ1qWsFIfLmct5+jja9cNOd8
gHi4cgUMYJzob0yCCTyCLZ/BSw1TfkLz7TXd6rvuNqMTSnR3oacCt4Q/7mQKeWcOCYzcyDRm0i0E
+Rv5AoJUkSWA2oONCecZgU915ShVWxnJt62dU4/jPYUHeV1//m6HPW8Ict0y7wGWF3jDMa4Ws2Yp
xYDn4GgbUFupNqWuDkbqvLG6w4r+jK2iirjZ5PSjzHUmi3+RTI4rFNh+e1Lr74Cj9BKVfv2WW3rj
yG3It7H1l7Uu4xO9+d3xu7wI/BVSCpCuUBiMlmXB9x+jrx7X+QNhWvHhh0evW0rbXVUv9FjCyhce
r9xjyCTmL68JjEcFTAa4+FoWh44pwj4rOnKEPmmQgBlNy1eaCNpailDKqgo05uVaV3QzZwijVWOy
GDbzHn044KbLyIGILFD5oKYNlQ8Cbr15GDNtD5kOx6s65kMg00Lwiwk95g6eVTr/S7IEyn75uSqR
YFEIZMo7J89sgzINYA7frOtyVExAQE+0BTWNA6R8ENDQfU1t8TQ8ySbo6QiNMSTfdLy8O2YBNEm2
frTiGWRBnATeS69GX6NkuKlQnmgvN03KbzQn7MoTPpmp5SZa0Et3ul5IZx9WzbgO5uaMI7hpuPNp
NaT1AhBF391NaRNs/kK8tqdERZzbfXh83qUbzeqGmG51whn0ctqWgXSXHJ08trdmW6iYjTzxWk89
kpTjlCMlT9i5F5x4+xyPSgn5dAE0cnZc+qZMVRbLW/0aYfeUOi42ngUlzEuFDunD03eQ6sPzVIBC
ljSFSp3XL65iABFmZ+5c4df7boCvk2b9VL7Sd4Ln1zvaKyZz/hoK5ZBXEVr5gvxvJ/ubs1T7UjLP
diDXScr+KHGK7zhGa2sem9qt5xQwBsMb2cGWvMBpKrmn0nbKRxyLbh2anvFlxsdmIojSTxE6q8/X
ohEkVdDCJHYf286SuJ1SkLw2uRrKj88/kVLADwvf7pL4vr2u8ZVejwtskfLe6HanXT0GsJZkB1Rc
eFXK8V8r6Lc+VXUp7vwb3ORcVwyv0JtnEWbeXeBUkhhS9rrfuFm5TVISb1o207wyHATDqUPd3kJj
CrgHsydRCCcwVL4f25HMc75BFigAat7/G9Svxg/J3niGjL00Mgs0DMBi2GH0F2NbvGS4aRbOMqiS
Wy+40gvZr3VIZmJjwVGGpOeklijrUl43vJ1ruwoec+21YNdk0VGV2OtcNQkLfc9brtTaJBrY647C
UjoUVccRq23WW0JI9gfM+T8IGi6g0zru6P1FPbBgsLfh6k/EU/MbFn/irEi0YG0uE7vDKAD938fr
zZUnfv3aQc/cTmzZWkN47hG5uHKVvzvkNhTqsn31gBDijwBsrCH0cy7b4Y/VU3E6KisBRkLjyzl5
zOi2MDY1Pjwa8Fo9zmDDiwIuj26WHuCszspZupLKSzTIrzue2rSFFPpOMfl4OoCmOPTILmrQ9751
yCjiFV2sGzGEW20nA4CBRuIWGRB327qProMWbHk2gtDeqzs36et5pROOVTYM9FKIH0ra7gXftJBy
WwcwiMA9XEb970mCKcjGRc/E45PlqDKE4GnbRRTG9vQLQSrUQN3MnXB4IUrcwTJBPSm9SrMYIoYZ
O13eNh9XwaAohNHu3YlHr8U1pTLOkP/okuPbdaC3cz0bCCnGiVztmrlSh55Zzuzvt37drGqdS0ct
KBfOWUEsxzcJfg1yx48Gd8LHmSLi/zu1HHCSNvDfEnnc4SJk9Qn75HOxgAMfcQA+w1G0PQQ9XCOP
sRYdDnTOZNILvuIsIvU5irV7jauDaGr1bH4eu/sOyEd3085opCJRU1t2WKlCFxdlN9WRLbCbS+4o
jPovZeXuZxGkWLTqS2gNq2g9/S8BGDmff78bt/43x1r3wbm6PrKcrTHgngLX1OEnVxfTTsYs1Qrn
vgypIOIsOib+/Wbnim6Q03fbLlhL3SmttkLqm7JwhhL7Qae24ZXmsABshRB/d+D0A1L9o+7+eFrU
VQ3vcxk4rBKkl3ffn9AsyVeqesxwbciH3mQjsty4qwfOVc5C6Pz3p82B6iXLFw2qpBS/hjBlGSiD
2dv97LBz28BQQmhCHCSJoTB43CoR+2MVLzwalsxj/DBOiyNmsnvTTiih0MV43hhVqz+Au1OWdZU8
+SlqPG4aqdVVy8/VrDl+MwXIjKs77zzFJw4yhj6ALQnNI1dhWTI2BhmcSyXwiGxQtPfgkuoCVdY/
+swCdxLdPzzWBNyB8s7BXzhZYSgvW3ZrCwLg6bay9GbIJWAB1Jh1y6NlLRa4+kFwDCTEzAH9ilB5
W4fvEZkYJSRPwjGhCzQJqnPfu7gw9XCz9pCg4iUa7fpBHbpw3PVx9R2gC7h8bt9edtyv4a30YXTP
ONZpPHFZUkFfdPGaIsEj4hPRjgI9yP/bx2wM7JNxdSPq5CgSbm9eHU6hGFpII1/Ze0u/K1Nj7FeI
WoIFW+zYzydBXDUBjXRVZXqisL77OwdZRVQ1GTXNsfTACGxhWC+1WDzNfij3XyC4gUp9ELrFKdL+
sdIGZgOxySgxU2Af2AGlQJa1e+6u0KntZSguVxcGEVR26bEqNXqo0x0dHbAgQ3xOyf6CzU+w2uPU
EzP/cr67HCmmnV8gmMPcGb8eMwRl4V10klMiK2VISMlWMeb4PiUre9hkeaAfaC5rcA/TiDIihdGC
GHaW7lUui83HgCPUELJg53ZXXidJRbxgEhXxB7R2M9RarJmuQKAIYkDk6OsGzIYgaE8FPRwVUmM4
Wt27urUceTLquzNI1qhwocxBSzobqf10yDYWnTX8zUX4MhmMNyYgvtMwMjwj0Xp6po60ii7meU3t
U0oW5OQb75klAr7ZgORuLUvB6wi0mbK+PkzcHh0mI4oBC1CBuJCuxJ9Cgo5gHp0xFRIiqIQdn/1O
ITz67np4K6K9zUIDvj2KJwhOxLp0OzPbjg1tTl71Io/zXJE6pbeKW/vSTlELE+hs7CU1xzkB6MKU
ngzHB/T0RiO4phghJKet8MVZrRQrDRpto6cTsJZH9sY81BZAPx7VYdswvHWtDTLOm9KCti/Cz7LN
0T7qTpOIagNw+NWKHlW4gRDNgywSOPZ/uYjt8A3NChaTvnbasiWjsLnZ27Odp4xTxvfFWLqnSlmZ
MiYUX1F083OiwjF2b92Kq+EwwaLAVCK6Eyq7vTmvy+gkf5t7B3pED2QOuGfWBlEVvujcchTSOHfY
/kuxiz/445Saz3Ty5cdbPGZ9+oT7IrUB/1Xq+yXMkblqbdN1gvKeBQRj1loS7+lHmozqNxVy+egE
abxpQvmsyRuDGAC6dtiMYPdZKzKiUsrFOUVaZ/lnKiau3tJHS2soAKYWfVlw2bfsPUOAQOdt4vF8
7hraroEF4SJWoYgjRctznTg1ynhZYVfchRNFlQ472kg8Lr5H8G1iXFANc0Mum/U5avWZ4d1+2TND
3f6Imp0IolDOV0iyr6sQYBouX9FIMEDb+qGV3Vm3zvvgYRRtBwUwnFifL14aVbClHph+Wu1DRohV
vjPd/Mvnl2CrH3moHbFxp5cIBgGaQDGvMLusOo3lIU8USdw8hR01lI3poFdpwMtr5Ejciu8ZeTYj
A43GKZjnHtCx95RFg3CJ4OBZJaIJfwd3NsCSrEdVK92RRXrx/V5+QGGbQ9jQ/PnJcvr0TiQSQpqT
ySBBx0mVe9aoc01/3Hzayk2EVKBwgaBlCRvpmjk34PG6Q0p/cCGR6RAK1Li59TAGRHKzSJvG/FcX
KN283ySvI2BD13IkSzyczA9t0RKrJ0CZzxLA4ZCJBWISnQ+1dXDgGtjgMIjO9liTx7cDaaPRglJ5
HMJ2t6t37VAHIwcUtWl4+diVCS3lh6THuC4h51BZkQf0jNnN/PshU9I6YzZWcXdQNl8Yqwg+QZUr
85DSVebKRqU0SqPGszSJOIfA9Ul+gjv82onnDvuSfc7uK6rmhLZNxo6tfykuq54dbT98HyzR3XBp
6hQcEVOM6sEHROLTiPKTDgneQ/TgUxtqan9XuSNfeml8MplxaOO3/bGKi5va0RoeaRPMWOO3hneg
Tnl7ND5RIPLz8CKYVOL5JwIaBIINTYrz6N4E3IJ13gAcyozcaYujBC0rbarv6W4M4wpWkaAHyPRU
PGoHT8EIabIL7Rx5t3ACSHobc5ll03pIT1aHsdDD/kKO37hLm35j0rm2Z2gR6dXUX3+kuEip/d0M
dUbNyEb7r4lTjxnBB1VZF5Piu4BTNJf3zhOTfS9Ogxs3QSxucWYAfFzRzFCTIEMjCHD4VWI1fncY
hPSxtoWw23a4NddCcgFwQWODx6llTY21pTl0sGv7J2vOi3I/2ZpPC1V0E6U1cVf16vqfa6Yx+AhX
46n95U7sPwJc0kD9ERrqAe8RZXMHkiW8RHibS2kl6f11MH5mYLfy0c4ihfrfekao+rkuR7yNzgS0
3CHUISsgWkaxWMPir5YD0wnNO3b+wStuCpMvE9ZcBMBjbPy3kkcbt5plOp60pjYeYbKkKV9tF1/3
m1S5Ek5Sd61awwP9d8KaUTX1XjG+i9MeupO4x1vO6JKQMTpTJCDdVw8v+Zb2N3wWS1bMjAd+83EI
BbFP82hUkS4+tXJPybGUsvht5jUyG8L66t3f9NGKOHVPxRjZDDBT1vh/nMkzUeDqbZkWEqAI3iSM
a+q20/b9bz/8JnCk7vDi+0YD3lpMKChRgQen7SBorB/nYPgL6zaW99U65Smrl/cO6vROjFJ7CxjG
CBeraCD3WQgZ6czaDr8NY6lDHWdQhd1vIzhtgyh5LwGbHnrue3O0/lwYOZ855e7EfpP0bYcfISCX
d1sXVVoiiSPKM9WfC7rvy9UJ8FTv3iHVQCaO7DZ+CS7VGrkSRco/LM/YJvcUSF1GP2PtB79a1TlS
K/T3PJg8kD/pz6rLmC7rTrp9EdbxBDrsZL4KOU5S+fkdTl/mO42JWl2M2cTM02BaRN4SWlboovk/
QszjcXxXYfcU/vCfrkkjo+KNyiAZpdZt3Q/7hew4yZ6Z8nY0PvAMCz5KsVdJly/CEkAtwWiyNMSA
OoCHu2aEC4y3xT7wp3e/m2niOt2AEM66P7dxkb0ODvSe7VTFBwtHypUJEWgCpHJCxbx1Fv32WdZA
iIu0rRY07kpRL637yGlJ7TNSOd/iJg6XNpicqR9fumC5VN4zAAx87Ua8TTiTOggQrv7DD31qDtzJ
98cjaxlCaSWz6pC3Fd7x7SFQiNmAETitkKNlHcOTpJujVJWChiPhIamsqAd+e4tsGU/0NHoioMkw
O9kEO9GsDCZS5r/2I0JTHr8Gm6f1R1tJJGJyNw6Gn32LksC5W4XtTpEhD0fbniioZGRdRQpz6wYr
l07+9au/AT/bpcniowQ1XWT55EUVVY5A8W8uKne3vDRdYfrApswhcHUnGi6CY2PacW6U8nTK6BZ1
E95p/L/KphsurLZhAsBf0kiDdFccukN29QXOV9kPsxzA2g7qyc2fSu50ugP5EdRM1dyU5NRSHQeu
/kDvJFoi35yIwXYfZpdBPVqLPwfAhQ2eDqlp/xTETw/b7OEfi24ljUgg8xvxII7DR7nscWu5mr4x
4ABh97CQCaQm/0vdDMBur6MuB6uki1dpMhLeT8Ka38/9SgYOkfE+S2cTVZDLss+7WcQxwUjGxQfi
zEQ22Qf1e891x+BO4jpvo91t2P6jafiKmbqOf/pDVwFCpi6Kuk5lssTLD2MkkcF4RiziQCOiV1BP
G8QAe74PBmx4dvLH4IXALFP30wsv/XezMnJaFR5UozdbIkPZM+ZG97KT65FrCwdCav71tsFFKYzJ
N//8UwmuroFVBPUTUrSJHfijVK0N2ltKIUf3tm6vAaItu8NoDLGr5XkPZe8D9lXBxloGl6L7RMou
NtobZhlfHNPqwdbU8wJ99zKkmCGKsRrzxoUg9OK/wMJ87br5xy5E+7X9yJdibrXjLJfRNHlOpj2e
UgKMn1l0e5FhxluHoT/VPtefQSvxdOto0Y2SrG46BwcvxBsjJk4VUA2Ik9WoyFiX0oJfoUbmCqCw
pqHEs5lKm7JIXD0G0VxFYCgh1TOsPPJi1UVPWRuB9pd0ZxKRkXz7sFJxiq08glu+Wwn186jS2z/3
Qt9v7Nm7k5LwtAhpOA2ZlwKYryLl3/nqDFD+NveX7Z4+We7Qh2/Wu2Fg6H3apo40ntCVRrH7Jf+1
81vvzJAP516yM7tosdM+1uSdKKudSR+VRiE0u+KZz3XT6L+CamkV0UxkpDDs8wsf3wCHoJp3J/rV
0tMC/5oII1aWB8DeeeqwlWDV9bVJWIn7hdqZVIuOLXOsSogAgsl/Gd28qKH1UJ/c5/6Ve2nNefwa
LbDLb4QHw9UMrHNm9/H8+0AUtvzkOd8vmO+hKMD4KPw5RHBTXhm7aw9mjTO2Z/ryFyhNvxMxuI4Q
ted+WShRAlPo5JpmevDcypL0AwgKoh80DmYBu6gkaJd3WgKKYd5XiuRnXhwLcb1iI3ULq5NKfGdP
M3wEBwbkThR/2Yb9WOlc2m+GKKM7Kl2+sigKinUHGcA7bWeRlhRVNxr8sTDl5TTXk/upBQwyBdEJ
+/3jBELKJYmo7DuLHSwFLSOBWggma03EMX6v4TPWknzDmw/URDmrGexVHPoy6P6lbvjYJw26MtNx
JJ8WL5aUFKIeQlmmNtrl+6DmdvZGi42yhLd4SsGl3twkccrtDDxoBM3CDkWsSZLyZ+QS+JLaCWf7
3PZQoGHbJrVksXT6K86pujvtoYWB6fX+nPnRTjv9y5KJbOmBx7Qb1HlXKHIAGX093GvD5gG4LCt6
8H0+SddBf4N3FhnVqjV7+7j1n32yJeCvkbgITeZT1/llWd4slEXkaHEc2M2y6Dr910nV5bmuh0vp
EV0rrHsggHv5kfobE+kGNgSrsdl9CRTpCYoDAP+lCBUprjvOaby1NN0Q2B3E2aLU2DZVzMXDF48l
bJ5nB8D04GTbeCEjGYqcSF1g6zyMpC/hySj6cm0YoGDluzw7URDNRhXT39jE8LynDqkaXdmneJ9K
1GiTdEcBu1q0l3dlHuZnxJ9WKVpW9WUIrBIfxp7echNa6IG9OOmFADx3puc6aflYaMApiFHOp8cW
hJuS8dSSd8z1zbZG+8AIXF8AssbtvPeqTDR3Qqp7j2fZ6u0o++lbZ/BsD8tp4dqyWbQgOaxGHW7r
Wwt1FcrSp08vLGqXpWHfTqHyW6te7SGW+XrPvJsMEGhRQnNu8mqre7j8ebCb7d8xkEPUHB3vxADQ
nEEq6Agaf5o/4kb0j6AV1zm0WLBndp+zE3yVLMFoXqUHNewx1JUc/ojbHUNEP6JTadVyeDGCbbFg
B9UIb7AJSfSUQmSmEX3afyBxOcWBMHXAWBLUjJE00FKMBKsDLQVG7uKj0hVMXzN5kIwszxdcPxoG
4l7osi3eat5Lc5e/2I/stzxu62LLb9bvivZ+vL9359OBQq1NZX1y1i9z7H8jpymKV3PRLiOUzfip
wON7/icyWNDPfEumYErhqEnP+6UDdp/iN9rGSXHn3NwrxX+NBSqBa94Kn5flN1qKeg0OkHFnISBC
GUsVywuD2HI1MR2Abw4RSqYLXZWOIXBaesMn+utYt7PBHKDb0sdAyvz0TrWQEvZPnEzUCfmg+gOc
ZL60hRgW/QHfObBBZMdWLVXIm0SvPHVhP1EU+25sHiC1A4T1VwM1ZMPI2Pqayuzwvj8qZ27sXqVP
M4DmEIaIyD4IoSm8UX2eS3XPZFUnc73FybnJXUtcKMhAUTezxXq8jnr/KBMxBH5XylPuHHQvFPkA
WRLrgrUkAwQrze0cspEKu35srgGSZR9j76lALmx859bVdaykTvOErRIfMvoziuTZzZdBttWN4w9E
DRvzQ81mavVpiLPgiKx9NesLWWxaUR9tMymOSmD+PQCxmRcekIm64wkTuM5mV3GbmligWIBv9Ss3
nN1bx9AfpHLQ7Qzo5Kbtt8uCOn3Pfsh6CQAPOOoz7n2EJve6zDZ1dLbpLvKwR6lYBaF9rLd+DfD/
HtEalVp0gwSmc7oBUKGlErOktMTXPRzWp7JhE2WluHSLxMb2fGnmEVlnPpa8eGTqP/ZME4fCkWpZ
8f/PHAafOrWKEQxRrheL7Og/Ubjpj7AMqmnadsvyyz22yEk+mBs0s19YsD2gOkpFGwRTfSMiQK9T
8Pr5h+qXrZxpP31BdxaPelmBJfD1Eg7lKDl87BYeTuvAnhEWrSZnbTQgPJIT9f89TzYSYO9WAxum
QCe5TDMR4Kk6WYtp7MlCcoPUWKvuiVf1fXEQq43/BBAUol1w2K+a+CvmOz0znu1IMsc058KO1602
dptjvmCJdA+fBAeNn2SLcLXxeUAZvpAuT7tK6g7c/6sqhXrty52y7l1Gb+jghTLhiqRLgROuEuNX
Wd/R+Dzp2VojaJ/XEiFzIBYSz7glYkN+DDc/l+88E8zYOVVctIsQSwnA42+r6b8Zzy2uB3hGWUqz
OrAzlTL2LRZvusSxr4aI32ICLag7eL8XGwdFi3+D8Mo2fr/qfmAHTp3Pdmi2XKCfhPEZKS481xsu
ynyt+tpZc6A+x0Jtk91lBG6tW6SqrsOOzi0XOz/nx9Ws3szdB2W9tK3gRKhE1XJLAvFfVFNf++Pm
fmyELl5H0TTpb40x+WzC+d0DWbzKX8EtUa8CEyYhwZMXLAGF/JShygzHmOmk3sgjoaAioLrIm8cj
QdYuBe4RQ5fpKaRGJof9zGTqzIbXZ7M4glQApL81euIQ17q8BbPTISmqqj3dSvgz+/wnldXOtq6q
nzo6zV+hxA1ro+u3rukPNbWuq6DdsDDXoTPVEzmp4653UtmbM6CXug3yxx2tKrnNYDMc4D8bsS3U
DIMbkRWiPsE5u/Q4hmZZ8MVLAilhUFy40j9Yz+LPs7kGh2LmXzIH8HgrkP3bGK9JmsjA1IVvE9oY
9ntDKNJWfDqNBpRKUYdHHjP/7UcRpfIv+6D/k2z0GAzHYZDYlx8Saqd5UHQZ8X5KUF2SYFCCGUHg
KK9TqIF/ZU31kLIxmNruiQ0RMXerqs0irY/Ip/FefJtvjFLAObZjA1VcJJXxFvT+LAYVzhPaUPHc
K8PM66LuK50acZ/wzhKywNOKuYD22UIEwpQMA06wGIp9JZaqrjBLZP2lasbT/ER1oEMXvnNzDaqK
UjnQWFugrrBZjWa2tp+uoPHY5b1eT9ZHxl2y/V4hfufGL5kD9eaTlB+kCth+WcgJdHbwSfdlgk0J
RoQ+tyZYyr+p8Yy1cjsnSiOkrLZqYdTRQ7ezcsQ4pYTRa6s+5VcDWwslPlvnnUJW7lqMxOcN0Tm4
uWimliZS7ZSblwU/txO78+byLWrIMi9FYH1ZrgKUCEF0yc8xGEc0KdZl4fVyoIaem7fx/ATTDcAs
1Zu/ePfg+v7yaJPGJqIesrNJ4AMEFhuY24iNDpMPKzw+r+c41NRl1xInMkf59hhODU6iWvnWvFsp
a9etNJrcUG5phY9AbateiVXSFaXxh0vaiusctoO4JSOE1goQtbLuIds7wVXTeR5XPCeAZ+L4ojx4
huwK8nhVFWSMngkchQa6SD+ZdE8aXchM4XL/Qfoa+sTWZ/DgnRA0fS0xmDPd4XWC2oeg5gk0xYcN
TD/+Sbrdko7zuKdi7c9jpeZS76Q0ByWELk+2buz3Tojz3yDamyq3DUI6ldYRqOzrxuHT9mpNxOvL
G5iA1BqJou+Cm4Nk+ssP+31pY40YJld734ZXyqJVwI5vqx4bhF3vlvMdw4rzoSMoz+BN6DkGfKMd
z3ppqfquqsxrkUrTGwcPaR58bhpHh4zxsyaitTn/gfr84AGHbDdP0V/CFv8b0g4C/4vUDe7Sc0Ru
wvarHeb5r+b4mpCBs+ZDVWyoFv3xbaJt3ND7fv5FoQCtzVypez/uftcDfVMBtBD0fw0WQtah5baB
giyzIgu1uFSAGWLVrp0frQF/63CGZBj9wMuXEd4yLhS0G3BPei9CMlc8Msq2I9TkasiXpXQHoX4L
0jlRfBXhAQteQg/DK5xC7m8EGXmCNvGi5Rqkx/LrQYtYy/0qx/wFOCNPLDSv1MglefdNMO1AWqmq
54nU/pJd6v3hQJP/kcwHKEiBUJR4OsQIseJihR+CFJTV6y9kic0g5EM1v0fIOExVIedk0e/3j/NZ
BUe4pfoJ3IPnGGsLzWqY/sLdquFgyRiTzwIbo+mfmVw3pXaD1ZVJKuU8eH65t37TVfUSaki7UJO2
OYooqtNwzVezzXDI7F9279DLzX9ETi2HUx57TZA5+1uOKvm+Be9NWJPcufuSQJMItbOlirmIZpb7
djbPm1VkPDdyiu8JdaHxMfuj85P3O6vcQ461ntSO9tug99rgiWY432t73Ty+6OCXh+EbXGCxeA7n
tkuh9ya9DlYN4uQ9RWJbPF2xHilJG/lE/c077l9t5coApmMsPblBMXW5IJB/d9gKh44cuhiOYvz4
kLX0QbMQWqsgN7MZrKTfvIMfUv+V7iUPixSbdjbPV++FIFBiFWDpdEo3tKjwjOylrdbDpznmMYX0
+b3yPzsVGXFq+LgxAlaxaJ5xyNiUTEiDuBygO4N6/e9ddFT64URJoJh01Sq1C1+qZjZhDt1yPiKf
pTDaPJ/USp9avQFehwq9kr1Wen9CSi0ax25F8zVPpJtf8r3jh0H6G/csOpC+k9J8eUpnOi6V+3Lb
8eX2xGlkkJ9d0uWUF65LIDy3mHPzOS5nmI3adfgUCK2p+TI/rYCqrQuh3+G84xjkwgoWD9osTiYw
u/xwfLYk9+CQEK4VNvDDZWslLX6kqmu1AocvLgly8izYDabA7jCKlQ2gQ+JhMhez0QCjEjDukzHc
1OlY8LRTdp222i6XsRsengsI8UujdrhAboa2D9IrIqtUCzp0KAIYPm5BcsRSsJ9Ey7a7xGfjqlEb
Rd/q78ijZFhp6IjvbECW2FjPE/bUk6DbrqikfGmOchZVYL5dQsznRdi1dvKK7Wm9IENdoFNRu12M
10QUlhzsTmmWbdyStpbADgwALFsumMwSAbU6VqP0pMePFF1n5BgRJyPqMmC3nJhTKsNpq/GnyHb+
ZQVk2+xCsBVkyWaaiKS/NJL/YquEJOaYA+R7vKnqfl8czh2O+AZuRcdqkFNjU7Jm2w26kABm6n8+
Lb+41hBcR3D/WL2VESRq/jtp5Bv8w6mSvCklGCLBH709YnEnVexEGAuR/At9MJkEt06tOQjw3n4f
V9kDJti1b60+ejXO+tqcYUXvx3IlB95D855R9MH0mmTbV/TxOx8ib/Kt1ckyBWaBIcj7Vm+CdIQ4
wiB7Bo6QYSxtlW8DhkqJT9M15tjOsh4pUkHw6LeJaU6OzIgRMJtWZYDL+WXRAy8ZOSVW10dCmGFU
/baDiAeDbhfEdIC2Argh+LXZktA2cBLqZA0CxbUdzv8k1UTZWDQXZWCvMsp+ikKgok7QAtrP36ge
Rv40dMbh04oggGMJtVhgvOgECUWf4D3Zss+hV9EpEEgf6yRWXfNeuOc2MU2+FKGOz4LkjJIaeE6i
6FVegXpRyJ472YiRpntvplPhZ3AGflBtg03GcUZu/ZIwx8BoEFs26Sjp0A/oIgslUUXXWp4U325r
Gkgu3IishVgfxq8YJrmjCdm60ONCRexbYI7/4QUWL/r7NB4XjTvQPKGBc/qb8bq3MDusDNQ159x8
b2v+z0DBj0ppfsZ8j+HQQWIDof4HMg2od9YEpLFebFhVSzMO3M/QWTG5ZuyInrsoe+5861sAC+oF
Xbovvp/UZhGfeUSbSw1yl2Xl871kx8fFLHC8n/3QVaitPmUMcAmt6KArAZAuqDldKaLXfZlrfaum
PSuVHAHMC9XV3B/7GY/zMkVA9j1j1wBeA1DLdy/t5zdPAA/8XY+Im7hfXrvuoUTVNkHPw9aZ+PAq
MkJDKDgdb9tOachrZt/HAJNz9TAajSGpCxteXvZ6qkGSCERN2cP1r0VZhtWzpxkgR4lfPuqOM/+0
QLo3a2FapRjX5UKjHYvl3ogEHEW3GAGFFCynql1MqNEfC65XNELVrW0J1sNgYILnpBa0PN6o5A0+
E69XwS8mUJSy54uWeqz1BEbpH8Jgh0GA8XwNVEmhylksidzG2xcI4CmSdhDVAjuK27e2UpLqcUH5
Rf9eRIxcEkpNOmuiau05g8h7rzOWzlU44NjEyc+ux8eoIUOkaZzBZWkEphhiLoyZlKI2X+fb3FTF
1ap3M/kNxfItBOpXJ7zx4i3C9aZwqRhypxlU9aBYYSQna9t0WJH+7f8KcPb2tID5v2Y1YcFoV1Bk
zm3J5GwNNbnstfYikuJdLM3Cg5OL4EURSWSRRbpuDKZTxL4XyuvaxkpEeHXfVuW7ugYhdjPQz5Pc
gfKj2jqkq//dT9EmyAGGXy8Bindcmy6OVFySh1C/CdONR0qeSK6r6UrQrFKW3yWbmklRs9J5CkJr
HAcZ9BNAm+C6TRoanvvlvOenqSVQg0BwSSo6Kw/l7DafvKSPyTzCJMxj0ZDXB5V4Plind7Dh8veT
MZk/L1IlHQiaEGC/yc6MNhpfgwaJZqcqjUxUWddbUyJDoF/yTdET2eHm8N0eiDZt23stMlMgA44p
0VwI6Uti+yrMuQCEB1uucZOeipEjkSDzQMW/MeWbtZtwn7OMUwdKaUu8UBq6X5SpLyJYOwdwL4iR
Qs2eYRhpwYdO4xtqyt+Zj0ENc6ZTiOXtIoNQlT7bANdnvtiUpIwgLfm7RfX/RLNNuthW61ZbB4hv
BokoGVI2YDzEgcaMZ9JLeX1bDj4Z+GTUv7kcMLWZitWQIX2qhmkBkjb1K/WqxWbPVAszay3gArbg
FzlK4aLMQ5KGFlQuDxtsGYxafM0gVqZ8hk4WGir4XSMVqm74AnF0d4OKSFf/vH9AnFySKn0uKupo
Z398aRu6Gbg41ysRa7IudVNjp+cRnT0MjgHfn4no0w13vkEEUxCJBJygvEfYrvl8CuqHeJCuExeA
bkLQCQj3uj146A8vYI7eF3eM8fmtKOorL5e6w1zRucBhiEnmCWMbw0yLQB4d86a8llxtxxhl5kPk
FkXEunlvb9CoeFCgw5M/E/R5y4dOIdjGuXY6RNSg4rpY2yd2leLqIzu4szWl3x23QeKYCIOZ7WmN
7UC6BXKH65VNJskEOsZAhSWmfGq10PJ1m+NFQkq0/wQkEeBrRzgQSrEVJtOSGssSY8KzXIcfSek0
5dmsUJkb634DxknIUG1CaiAV13QxXkwQLwJ+XMJOwyRdp1pNVPRlduxUG6TAsUKLWZ1NMjg8mbqY
sOEpsi5TrUkPh1nFHBNUYNRTZZcNHI753fdl4Z6fTX+DVWuL6p28QpVmCmXomnDRWaMvhUAqrOBr
k2QK4sJ1yYTfh/94L5a/DoMWdsqkrqwpmk7itZYWiVxHiiGR4V/rburJ0H/AAnUT9pMe+ouzMvsM
XR72CJ8ZmQPZBdINXIJ7R2AHQ1AueTA0DW9J+d/sW5BBVvJUjQPcKC0ivj5nyohuIlpd54LFkH6x
WpSTIPygg7GOd6IBhjPBxRHYnQBQzh2QsfQBXC3QhON7uxveqFrGvruzlDrpFXSKQYfux800KepV
io8OWBVy7BEBE0n8NM/0waNnRBvCRcM2gHTgVVApnkO2gDtG2JW4yypFy6pIRcjgeZZvLHWz1aq8
Y5EX2HpjerZQb/da6qXe7EilXBYRY+57fyJ+fIl5N/K5GoDeY6Mja9QXbHZ5wrwvm7MgviN+ZOvG
s7sziHBywxrODqQRpF2Dld8uTTICKvGqSwM6i8s0koHtAE5JlCsvR3r/Abmw9bjlsLAtE4JpIbtf
HUHAxPe/O1EpvPKTbTgFWIubzSmWyFHG4Z/0E/joUvjBjnbsQvJ3tyOwmJ/CLeiVeTfMJ7N5d0ja
ABxzwiWMdgRVARfmIkkAlqWtUEcf6pP2P5SOv824HDgx724Bru33izadBFrbNuvBYPrvIKNqI+EP
6yBy97/tAT41LIy5JDQ7gTkKucmFbTkO+z4LdAGqgI6OnptrE6sd8apO+m19ZeXVcuX98xi0SiML
0eLcjaGbJTiU2QvsdPygHIBQcZD5yfhekHXbU94TE9Kel8Ktfo44RAkwF8VZEbzoRxESaVGqvJrO
xn7LJf+LBX58Xter1oCiT6+zWvAxLUNlXCIAdsZpzymfNFaq0jPD0n1vTe0kvzyRjHryLESL7Bkb
FuA+B8RCGOnUge/BfqStTzQE99V2AWtQIRbgQ343c+WbR6aX7B3ZWvM+bJQkuqlPhjrKr5eU26YS
y8vf1W7Uy3p3xCQ/NS31j2r/gdBVeiGD7gEEBBv76ElEYH9TFvrc4r9lso4Kq90LTTRYKv1LKDSV
7i2jmFvoGaMSkcIZeG5K35vVvV+L2Dv7RZIj92MjdzqkbVixc1GCcl636WuGPhteqPizMiOYscI9
l/vp46EoBcy8oA1XsvILbqUxyLYTRktN82t+XOd0xwtVxdcCtoRoIS3pBQ8ewPpStqPCmaXBr9nx
2LCy3N99Zcwv1KH/rv7acT3VKVGYNlEy8WQaY22zYtOQSQTZPSAR1ru+5nQqh0ZcLC/C4CTDDbmC
C8z8STh2/aSDwJwlsoerIggDe77Tv/6AG/0m3x08Jeh+CHn5Kiy0xC6fLazws+zar0WEHYpKXmRl
2Ny54On4DKQaAhBjGlGY3qe0mVl8bOTRM8n3qYPqHTneR6+48nZYSdWveaQ9vi8kuc9O7wABxKm7
7t6khP3mn7ZK6EdSHT4Jp7ezYg43ctZXI3SYCrUISQ9fEWdUgMHVTMajuqnd+6KdWIyx2NcjkVxW
jY5WFt4Z3wqcnGuGQrqmUjHYghIriklkGB1AuDKnxtjyOipBKkNyQoPzfKWBYKPtC6dhxcJdziDZ
uiZEJfdIx848z5YN6SLteRFzWj2+A827K6KdhOBeP6EvCz5seSQr1i7UNjeIQjxleAVySqo5/7D4
1kDJmMLnHaSFJEVHUB9o54+z9C63Wj+b9d5BlQ+2U5mXKqv7blVNnifd9ISJ0yjAiURdmySEvZMK
fNTtLFzJzzel112/GJaFAyvStP/W5vmL8+A1fWVaNHkgl5t2w9UN1Ag64LfTYkogXw1P91HZLRYs
2XlhF+uxY2n0N9dEHzgH/1OFdhkdAz9y0Ueh9SzXvgfMUSE5JvRjoJj4jUg6rKLWVeltD9mKTEaT
GhJcg+14qwTikO0wrpAthdGqtQbtjB9jaCFK7OtCSdcSqI62tZsvTLtj1nvKC125MeZYdb5BETO6
SjCyxpg0A2y0/nyGAgQ8ePr7HJ5GGYjxtxXsLuDxe/KJ37OZ0bOybvYpQ5W8duo1TI2NMd+cZFTJ
p44gk++UHtHCRpuOUvfrA0vfg3Dq9QsCEsLM1RcK8JANAN1ciWPNRH3VlHLUXOoDfenVNwcOkonU
NJbqMsySCjWQ269fwe/kwpCNxM3oCZjUnsPs+aiapSgg9wAZGHgp3rAMxgfyz7iLY0Qs9B2qBljq
/85W5bnJEK5mDhognaja0BDAI3p9oZcZnDJyrr9CnzhaYGYEoekHRMDcJXRq5UVotAPhTD8CZc+V
sKmC4l+UyJLmYXvu6YHAUkKfLbdR6ZtwcHb5rEmMN/BjZaaQjHJdxPjVyKdWWl0RkSxIWZrNrCgV
1h0rxRHdPC8zb8VdRUkkI8bHok7LtfCkWyXjtYF36lBX2mRa5x3sVTDPfm27IZDmds4CoG/kQO+h
e9kM8p2zbpT8h7SBzNQ1GFBsVVACxZ4DNaZ97DDDXzXKG0QXSjOqn8Ospqf+QlW6FYVNuAfIqzAm
GrJLsBpH3vhH6czNuQ5p+oyxQCtpzrKHKyWnMRb9gKcOgTLq4vZLEf7w7P5JrZ8f1/bkwH7RVmgp
zp2qImj0IH27V6ovKyDgm0sR3GOMKhECBRCETUh/tko97h+SDhV4/PPRyHu/8BOw1cqVqlk7cQ89
yaxCJkP7pAFPawpf9WYcm/bjpG6ybSkDy/X1G7bBzs8/mYqKkex6a8b01oyy/rDEsS5uVV0f44/p
BDV4U85kNg1b54sBCCw4F/6SeCdLGUozfbW1a8ciKX14swjZHLrQttyaDljytwn53D5L1PSn3/qt
s9sjka/45eKXgXnf4lFw9+j7hcUcele2HSKmcIksPb3eOrfH+PDDSqNNC7Dx0Fi+jCf7cPN6musz
tk+VZJcFPnx/yT3czEwZRZLU/3DEZfIqGnaTDnNQTxllfYvDdgtGUXdAl0kYcvlTqZEaP8j0yN5Q
/TccIxfT6x0bH82CYolUqtqn2TLdnNbXR6CCFA6aMsqYoUHum2e3uLofnCAxtmbPhbXeUD04Uxww
IxjMdpz1FN7JF5uZyzDa2ZssegpZPIePusDlFPqX3OCZYxdDpcwekbKZQKzG3OLDaVS3PLIYhuSB
6kj08WXKrNkl2qZvc8d0zK0imdX9PPyz93AWoLuyLVApwCW4uAFOMQ5ogmFtaQCXlLJasoD9cGT1
GHtCYAKSv2IGoK1anXzgqY7c1j7Y+y6bIEVrAf36iy7VRx3hHySTbuc/SfeN5GIHta2530ofvH1W
giD1zKdCpuI1jimknTKMa21Ld7Wc8xMFk6zWedVOK+RT+/Lu5zNpAQQ8j7HK04UMEv3n4IV0jC9W
Uh4Z6c6E5gHyuJX/+Pq/ZsyvfKEwbhvyKnoJe0wi6Claq1z2XIIQqr1lDazU1rthvsEqg3VONBxP
KfePz1CS4M8PSH+1vXuALf6GXBwyd6r1FfB49GYPcCggfJ4NvqSSnFK3jVbMOxMKiaPyyrRnSVJr
apJcma1FiOFACzy75aK5YLQRseZg04rbZei08THkn0U4eEaJEK3BKIfHS2ChSFgCXwdP28vhgv7+
lsmXJpKFpoHJZVcH3ySJWNlbfMAo3n0p8gBiURQvqVYHubwLXKfHw66HKu4W7eUpa+hNjhodYiq/
wFwfkXzWrjBoa4hlxEIgRbZ2v0rUd5k4dyBAaYXE6q2mJZx5YbWufh/WFiII6cxGujMsvmeOh46L
dWTlc8W7PvIIlGTCirKvg423hkyTtmOyZalRNkzSCiUld5YzeiSj0oxJihnXpkLb78d5Lpl2cn3e
2EQO/ZtHbLBxO4nql/FD3Tx0e45YsDvwodQMT9N7Ujcx0my/A31CzA4YzFyzyWZioCAZmUR4Tkk8
4c4derS3MNpQFVCQ2o+2y6K6/Hc9mX27xjtzw9uYyEdIUR7OeYqgjdCsKKmRWXWS59lDQ3jrG3ls
04NM2Ul6kYhJ4VVMyjqLAQBewIpaoJh/4OAoo/i/KSmYdZZHF3GhvYbLWRF+7pHgg8SpIpttnuD7
Sev3cujzJfKYAYj+7b9fA5z0zxfi6EVva3jR9p/DTqOO1YQxW99CHyv+hNiaOarOBvTf6sxnwq1n
l9Qp9k3TZXAmMk0oYbaF/bAxs5ogTJ5LHI1UQAep++39fAytzDaZ+AfpMYL4CkLDJI4LXvH2IT+H
u8yclf0W/zVr9mgiLVIBJ7PecJME6IthvffwWYVaX1LIIqfgYDuR/ypTHkgJxonltTj63yN0AW/j
uQcC7RLQJ76J3zlEB3H/jys5IeqkNj5YxsM5ZGdo+/Py6YwCQnrZkGSTrPKQLikqe1aEB7xXOFkb
eZbOVK24H3BRKz2mLH5lf771RF30nrbLvNE3jzvPxYjG1v8zyYoQfKuTg1J1L2SFg2eKpAE0Ykvt
4GqLD4WVq9s81uncBil8aSYEtB6EoZP7LVRMNxWMp2oVaFU0rllyiDvqg8qpVZF+BezIUB67Mh2V
+VYmZIHneZ6JhtLVKk+3CKosbHUpzgveLBBgIPFRWDdoFsTYb9WN9LDfkIIpJHErSHqwv0tKyfvw
LQANSTHIPch0VJ9bxdMVYDYACSTglwpwY6cNbviWZl3Aylslls/4UfiFUfySAAYfcduE3XFKnI4r
J2bdpQFP2hBLQwTlefRNbqPr3RHC09hacVoztUKzacm7D21uqdY19ldzkk/a4El9WeL0kFzoGSR9
2T79P+607dy8Uo8xeych+P0G89637r/xkPso8ruxl8QamFs2bmSSiM94Z6xuSTDJI4ah7QRTXQRZ
BZWZzBWFfuuGh3tFwZZcK/T0Oc3RLkJgXXZsa4Kj1h3usVng+OTAfVwRwVkow2cP/AemK5BVqalX
vEMkTgKnKL/qtZzI69mo+lxAYh1gsjyYUzIv3K3E42tJ+sre8KjIPE3SnIOH+H9JDFkg++CWps8+
J1BrdNZzyGwzZJ2wVT9oicaJFt42KhCzG9IPH1PXjLv9lIYDI1frBk1+GQITBRcjH19p3BUOU3sf
RlolWCAYiwesvX0gfdHfFA95NcTTWP8bw7UrRpJDgwxYtMrPP1/MmGLp3RhBIceFvHgHksfj6d3r
M28P+BKCwDqiS4L3oP4kbDhJxnfRESWxzGEH5qP4P/vDshWaKy3m+rDFzuBBN0yJGRkzjKL45bZ9
A0vPo09bBAjAf+ec30akNkmehaNO+3xbgspwpq74SRkf8wdiH5bPsyQQCv+abvtrE/LxHZjOPGGs
sRDMFmB3rMBIufhgmNiqnLyWTdT4syEdLp9CJgSYJ+KPQ6YTDOKiIbeX9WTFZrCcY/RCG4NHyWHp
+r/Jwi8l9mg4f6RW7d3my8SoY5+cPOnZOrgo1YevrscXq/rjDm3TKOGMEjnTg/U+Nj3nXSfI44Vp
EQZWcYEqaTgQ9VTMigschl0G2BjtJl4Hv/fbxZerhfsOWLm813lp91rYhVuKtGokg5rz7/uBDMKt
Hag/C08SKgy/LwZ3ZakebTMRL0twWsIhqRjUnPi6VYR4i+eVkTIsuGPafp3nWU2WnY4u5e4suEBz
bH9hv0y3aOSbhzdWEQ9JYIrJmjruJXm64Tq+rLD7yIZFr6Amva1F+EP8YDrXFOBuVBMqo4RIaCp8
T+N87SlTDhsznLHjLCSyIqbjggvovWZvVqncrnZnFCzgEKgmqHTNjJJJaI/j2tzgxi54vjGdqZWu
cCGiAHoQKrRVCIlmwBGeIKBaQrcr1ENTv2c1OvgrwyB6EzUu532Ix/bQTvcNnjuKW9OsZM+r6Xdk
oTgBYnDs7WHJy4aSvA5LS8nq7YvPNL+Nlo4d2OsI4hFGKHLHJoQ9M681RjdQHrUf/9pLLs9KbVBK
4E98gwN1qSm8TN7VGsKXug9HDdR9s4DpsnEzUWa3DW2gFu0kw1codNaJ4Zg9LYWGlhlcm8+4yfyR
PYznQbLf+M7iIHodx0DgUAF6iTrpQjjeUyYby+Bc0mjvF3JjarOR8C+TPRr/5se7mnQR8SO05jIn
W6sEvgrVaU2gf1GcPnj8HYSuKcrUnZTb/157bN+imiuuwPkUeMfFYNXz34O8VLzCF8JQrr/MNPMg
gNyHPINfT2LG154hiu1zBW29da8Dg1CJMEA+qrZtrjVIvBJAafp0eY92QuZjH+12eIEnNa+ieukM
Az7USXf/QC1oYhxIfQ7qtNfAWHMJDnykpSOFtZ+5rI+UINeIYZHF5NRnl+nnmFgmFXJFyfPpyWCI
uIFL7ZPR82Ef5/8Gw7AouKKRyOnYx8qbwGvwwi86YHzYeGxrwPI8JfkwacmJAD4OGFS7CYBZtwiK
HZMzqvLIPAi1k3FayX8O0MT7rPiEXAaMuC6JGaUvFWyEGdG3tusVnMMpUKwnzaCB2aIaxqM3vovp
AmxjufktqnGchweDsNSvrTGt5B/Xbs1r0bs3Yjl2p7I+yxC5r8LDZN6I8z8Y4t/T1daqmOwsN46q
atv9VrrrWEorVIHa5CYbYQIsn2wJZtolU25KGBx2bBRMbpUKHbiMoi//V36uURylqZQlPt3JK7GB
Hp1c6A9pvp+H9tLLdZlV8PR1nc2XSu0gLVagV15ojvSlcunsCfLFs6PiHT1RnhfxX+Ma8ux3F0ZK
VsCL8cpouNl1tsYKYCdjfY5raGrdG5cy5eyq3KN6DGh6FcaOJB0bOwNWHcX4MTk3zFkLo5NzeWSc
nAk4eeJ3vePmgXUFgpzd/Vbfm4r5iWPe9Kiow/GbyRMvS0EbjDsStqYM9iUlcpE+h1p44ddQRFck
5aeiafTGmoizvbX+9c/yunkMelLMBRwlkoU6QMyzPAFjM2Ld92P2riIoP3gaGYllciJiApJUcfbL
clvd7z7XZ1xZTi10YnSmlVEwADvaRgMW1unorJScLC8Njf6WBhOvw2zxgHx4dy1r9lf8XrhDkC0B
EOXjUGn0zNgpCxVJ+f8L9j5HRcXYZUCUTZ6PxBujECws4zGJX9X4VQxyCyF7qsHcjvqQaIQWZ2UH
B2HMMo3JE3lNKyvxSxXq6sXxKaGF63tLmdmDUo+bODaxRShj7TWCsmj7nu0nM2UCmBFn4eyva11Y
f9iXJCtUWy5aCVcJlsXlf52Xd2qh4iHvTD8yQvwIFqGDVBuboDGKQ6G//V96QF2gn6dgPs4xuF1P
Lr4TytPADN7wz89twozjVtyBEuMZnOv5xlZwuGm+QfInq3ic2QEaSvxxQ7SoMffzK15LZAshWl9O
p7IrOdhIOMSmgcHfikvG2lwX02F3YIBB7LmLQRWHlwwrsRn1ofJHsYWGKDReblSj76NFYnqDxfq5
yhqW4I5KAHrSAwDHMYg8Z1kJqVvHyPqI+oxIDWUDC1K7QMsEHZDQVCYNQVe5WPbfcz+pDeZJEvgH
6iIppzEj0TJ/tnMoUMH3otdfVXWozL/ooeg1h+wriR3siKFHjYiBcytjer+yxvTQRY0kZQn0hGwW
RiWttJyjiM1Y6b8nWsheub5cgXFsgDcnvMitJzMYVa78ILWhNRHb1g00t7K8Ne5eoXmf7ytLutLR
KhdKhe7zfg+P4ZlMvo8al6dFn2nv5JJ2mezD99V5WTAF1w6mT91zR0fMrSHfeWtaMXM0ju3sLMGr
o9tTosdyeTlRjapgqYyGHcznNYZbuRldw0JLmdsm/i+jiwPQSX/hKzu8b6sLsg08qV1S1Z2Tp+2g
4dewUalNLp8tAuu8M+zubv/tcICr/xopjOFQVXa+5XGtcZvzploqLy3evVhMIRggKme6QAadbWkN
XLll2r22vgp1g7DXoibZbeHSzQAwrMzWesCjMuEgbupl/1qABOpYLLT2sDvekC9yIZsZtAB/aeRM
bTynK28TtzZJzug7gd9Ys7kTJNIpcMGgJtDuSX+g1vm0f6ZBklc0BlQeBHUJon38itxPkmBvZ/9M
MWwgY45Qm/wrHhdbWJ0fH7ynHddIMs06IyqlqcWlbwWR5+5h5Bnm9y7FctMKI0lnVt69Yanil54u
0QMy4Xsvmry96j1iLCAWzlQXGE2Y6dnPwc2ysoK3bWkfuvMx6jjZxoB2lJhykw3OxWDKZRxYZSrf
08s2Xexz+5wFbzan91eaQi6RakrWLat1sXgL5CbptxBXgcck2CQ20d2MDv66vsPKj0wK3uRn16p1
0LxHTAnwFYVznGhYAFY/3+K1aNXTDzo93IfNlc/XE7Yq1PZY59rzyyQxtsLkUq1OfXCJAQ0/DGO0
HLf4kcH+J8yCpopi1Yzj+9rXe0WBnJuYiiM6lmhZLEgFt2ImRdvKcigLevrRGeObgUMGdhhjxW/r
B/VmAOzzwETdaI/mPv8px2KSDZG0GEgO6BjJfAtJMybQv/Ks7tp0vltov6H0OiFNvMIp2L8Fndpg
+xFf0ywDyhkPIdfXOg6ACZvRlaW41WuYNsOU14QDe7cuIIEuEZV46vwtVmOHCMFnd6+Lnd60itkE
lPhZTHTY86pv+mf4b+Gec/xsrIOicY3xdclLc+ynTT5RKzetMQeOMUb+DM+reWTWNm0EGaUiAgRd
hM+X8PkyV8rA8a5FKg3xE+Aqp90iol86My04nlAMAbmRjlpmnW/B6BfhW1/AQ21F/frdjD+aqlEp
Yxu1jTczd20b5uUb1BvCD0kakliueHQbVO1E0dfBYDeIYzXASkz+6LHZe6s734GFOHW8e1zh4RWG
BuxWNgKNdf3VKzDTv8Qzglt9mwHdnY+Da74lD/0GBN/1GdqyNECaLVjQVZoK4jCFJ6VBw6w+5+u9
9zZZi4AIxBIpkPrSvzaDpbVlBEtfUOWfpYNpdf2ZsTrnhxWcAgIgmjm1PPYwMigEQx0ZtOMnNhN8
wLj0RqudSnIi2jHOsGSQT3VDkIo2/MMXanhFHTykSwR55IZIKBbVYGTg8MPm7Renh3GcoMM3AHrU
i104sgK25+81MqGMfmkNOCYcXOmtEyk3BmJ+lcCTqoteobi8Y9lG3t7OzgNMVsFBTC/zwrrjtYAv
TCPLrWcaK9xYeq8mxPdHkHbzMVPfIarVCiIsuDUdc3y7EuQJx/ml3tiDGrByGMyI1QK/oyOW+R6V
vEGRuIQBnMf/WhH9AptF0/wi+OaP4jAAy+ctB5AVs/JzqEakeWATIh+FLGbBFkMynRI25pmRxIuc
AyGpW/+ajZGeuPR6leW5XW4GdUMVa81eYDmoicpwdPfldJuZEwA0Gmbd3jCIk+AkhBE/JD7oZ7Ex
av+hoFrTVgt12tTaZs4e/dGKr1LT6hDdCxCgTMaQCfLY2nMLq6Jak8N0gySb0pAdHDPqWjYWBoSb
7YphqGLyiPnIyRn1coQGBS9WOwkyRMQY5DWFyRZNw05EInu3cCJpY0Sroh5zuu5ywL7F4uddIRde
i9bRcBwSYzAlyFafvU4PbBm1hKNuMsJVTs21zPqVop2AV4hOpHLxygC2t3qENTADOeZdZPLpTjC7
eGCsLPl6MHrq17FmE6Yolga12nu3JuMLXUTM5LUAkcpfJEBSPv37yGvA/O2dU86GuIoMuAs6QIAd
xJm8satLAnyTNcPGD5rw85X1JAVFQlMzFKcUEv+4mNw3cBAPMhE689ahEHvs3wS+st+Qn2kAiAEF
L0jods8G8A8po35erl2Qz/36xHSre3RDUKTEfkQCYcfT2HniusnUcCODc4MsROMdRKbwPmmHym4j
xEgXnKt/YjNZHpJ8TJ/ACbRT8Iw9DXrwd5H06a6VZauB6Yrs8QzD2jgweJ5GU0jiQntA4aCltBpA
05VXTpm0ALv23GrRBjXkFYUnMCXeezvB9tQJd9485TVY3+L5ZqGigaI3g4GuH4j7RjtCDUT8JwHG
tbx+gz9y0jiPrU3RDrj1QJez8Wq2Acc4WDE3d2oqd8L4ryq4pzaAHkoes3qwJ8gpWCxSFD8dJEXd
s8zoVqNAvo9ZCxb3s93APVZMHlKUp9ZdWEWd82GvCs22hLEixvkl20xaqYPCN2eCANtRSVLN5zIo
N17kVONu0YK+LwqQAdJ9jN+9HfS0ygpf/INZEcYlVTWRETLQ0wasROvOxUse9S3okMdG8skP1QtP
qbTBqBwdPbuT8gKBG7YULKmejjSs4i/Zr7iq+P2lz8m50yP/K2vN1VfoG3FF29EoKOGKeuqDqsCf
1vxieQRUYBRUN1IpKrWB50kciBdoexyCosdEyiErrCIXx0ZsFwm1YpbD8nx2nMXf/yE3L4j7g+CV
Q6vogw7ylefqTYp/iS1dKbHD6q8qxUb+d1CESDT7ZHVS0Tdk8SN9zExNPMUw3u2AsjzQSqUM4wH5
9EttmsSBD+8G4/wDTNDJmyI9W8WAeiHymep55XYyYqirb398XWUA/99IxO9FB4OggglA8y9w68fl
CPB7iirGqN1hZsED25fKlS0dLx7peAyW5oAt8iDgz5byDm7WOJl1KKssROukPiisC7YM0K6EMVpK
asxczxlRbOktYiKVVHG9WY3JkLx5+F84Kxt0Jm0TJwh/wb5CoDdPnCshbRiT+Ot2IrANT37AR5sU
ijyiaXA0LkXFHe9RJydZCtD8S+3lZeHVFmK1ZQpdPmAiu32Be+mNSg2dH83ootC/gaVeEmMUeckb
894JbQtMBjUU83hFiyx1CEf37edm9Xt0FEkkrBFdaOgFi3Jmqmp61T8VkyKIAktZj1aOk+8xEOMU
s9citdOHciT7Oc27uzgXbnozALgZy59CtjGujX+du2JWguu4DO2Jwnd11JhAiwh2ayhVEtosXIax
NKkiuFmOEZuAfdlNS50N3PzGG3vDqsamMMVo08Us5ciyFFWEvqZBDxlUt4RnoqMHqVU+2bncTQZ8
tvZeqLApVYgAzus5R5K+6VrbV/Qp5c1TP+S3oh7zhxLXYyJwmOKotnDx6HK16vR/x1I6NLKB8fip
BjyQZjSATXQLSRlt8JiycNKz20rNjJOmr4vskW/YmJlgtjuumbq/qXuLCLxQOK+GAvbe+XZ95fqo
9hv+0u5/C2UBWEred1ew4MzAHK8Suhcg6K6B041rNpeW/el4f01FdacepTSgsY3Yvp8Q3MrN7rbK
JWoeohnA0bD3RDohIW1hy5+0Oct3hiQZ2kKOBB2MevkdjTtA+/QFy8iRPvKmlpuAROQHP1KcTgHg
rdzYL8TjifrFnh8POPdgSFj/pb8A99dVam+Jb51IFmn/dFmFppJq1S7DweKuvQ9lkzbz/oXxlIWJ
yywWB1sO2EgLMXHp5SCdQ/kwvGP5F/Sh8wPE6p3SYQQsBFhEHML6L78sLHDClA3FeTWBiSgKPwth
m5lHOUcTtNHpGa7DGTrpyzFId1k2xS5tt7x98CnOT6GhU1QHr8m5xFY6g8KoTIYPckN1fLI7eh+C
lVQWYt37HD2YO70wix37kRwx4NeOGbzwrQix2YcHHvHfiIDUMZJhP1N7TbmCAA0xQQfyGC8ge6Zw
xE5yUTXwAFwTg8FhQCrzqxgMfyYRbc1C0iBa9/arLhRQDWlrwdhMyEu/qkTKNLLlSriTMGGXImhA
3UeR32B+UOWNWP5U1MI5dt6ygkuDM3p2KV/X6aG5uwDvgIW73GalP2PK+b78gOelO09MeTTGxjtg
qzcpfxtpfUaffGfADQ8y9GMZPaKWtnjDJWyszinlW6ZLKQUpJM/w7lSnMOhWa1xIY8CpBkX7ylX1
P8jWEoD4prDCEVTiJizdAd0DVqCq1+QigEditAHMFGeourKtx4m6G5Eww0LcYVfvQ8pnwFZDfBXf
pAYBflS4TKfOWJdtwxeqCfQ8Z55ApwIgzIrCnxjznGLWh73xRvy9o5wzyQHn7CXwdUZrj3AM+glf
7weRAunSBd1flU/yYr41OwQ1OQdzz6RPFnufJgaediWlIlwrQhqoKH2tDjg/sDXuDJMw2dyFpb0P
8dP0dwuB2NI3ryQOsUExa4QPMAjG2lqzMztqxHDkV3+SWeBip5Gz3ZEwvpmGAvsDYOsq47YsOAIq
TP67G9Tvlv/zbJd5q2U9LCYI/QlnQe/j08s7ZMcj9vr+BihzxWAYSO/I4K4ZKVrd5rImEVQffZaY
bW2Bc40ynew9PlpfdBHdRyqrBeUzEVkStomlB7uVHWdvY2SqmBiEos1LP0v4GctsHKYNcAReNADM
7+/hTtdIjlv23YiA4wSpVbQ7ZKCQo9OaULyjYXSFEqTjTprf1lw+QUHpyAG38S6G3/RaeW+uZ9Xx
Z6DWs8MCvG0Jn+zHJkjE7RcPvo7hDpTORss2QaM7Za1jRAJkAFEg3Sa/4LDpoj7TBFgBfYLsppEU
3XrVj+Ch8XQIU0LNs0xnZ+dcLfJrUBzFN0fp9rotasEkXnAtbhHmUjsQfsPIq/5mv2LTA6O+GcyO
QXT5JpxbqJoGsiqj/W/auWy565RIIT1WYIGVxVDPIc/M9nJyvwpi2H7Z5rXC5UOO+hlKlBTUi/m3
a/yKz+uF0DcViASC2s5m5upOqe3WwF/vv3tdR9O7fl+8wCUjt9Z2nu+yGyWjF3LIumQMWsU0i1/B
El24fJXOf+Sp0ojXZFh/r0rKU7OymKZv6iaqh8seF8AL4DoPPYaYxI8LVzJJ9KIx7Q16l3zcA/A7
KzHkf4B0mbNvU1vvVaoAW16C+OdnayPo0l+9nWd6Rthoz05fYSOjki5IIf47gz5Wtqcq6YrCBE7p
HuZSdesgjK+izIZ9irty+Lt/tu1WtnX1VeienM897t+uDNJbxau9eVqlUAhc1heXYdO+7n5SVR0k
tfSCXUEfYfkXxzFkdoxhL4prMrkM4MUYAWj3GVDa9ZEotNHIRN/BYfQ5tqim+N5XhReyRYOs6cV0
+IS9nZo5CeaHGYVjOCFmPRxPyJRjGCuDVT0E1M94wSbunm69mbYJRc7Kp7tm9Re8Q1Gug6VzcazO
TK/wYtn6Fx/8pggCQgha3y66udiJwpmkv65xArBO7iZfZHeAHJQKn56hlEBJdrpxIgtVzHYQLJed
LRqELWNfIm5IsYwjMi0ldJEORCX4RIz+YYu3NGCF751YjlsVH5FYZI74CNhLtbftbou6E7h+bC8+
6EUBfsLyV/oPJSKogeYwrGsWbSUqtBTUQCKJ60L3MbYJ03kzzmGJWMkGaGBhTPGn6tpssEaB8Szw
YrfpWGhlLCVTSpiDDD9MRmE1mO2/OfBFFMh1Bse1efishzDiFZ6F+Lew89sqORY8kmc+zGF2DbOc
oQKsZjGn6I2i9xSozIs176i/oi7ODvPuJ5KaWbm/acEesV7l3xJcq4kPQyjN/2DAhvczUu3hQMAq
KbUgYrE6kc38XbMhb1vCxNKkN0Jma5dRr7ad4RMsOEGUHCc7oD3gMnNlsGKWGrJShBkbD7JEz1Tp
CYQ/aXr+eZTmS7Q9J5HoYeUx2vEZG4r6SAl12VLxVs/xXOLKhla3rUApn7ul4F/j1Zp7JZTOI8o+
D5wTtNum90ggwf0NS8aY+OuzDmeoi2Uz1NXtdWqRctVtBiKkVs08eElCMo8XD48/2KSMqgEROzVG
fKMarM2Knf9OJO+CUtxNpGqBnIdEQqsM3dI1AQmxkyfLPSBz/Hdit+BhqHRqY6BuXzQ+9RksKYvJ
wPL+/ttVBS4IfaKjIx5xDbPDwnzyJd/t7AyXItbcNlY31vvt/Dz9dee9pn4o3CZZKlhpXd9QIg5r
uW/pT7Dstir4ZyrbZxTV9NH0Sqex2yuSx93BSXEOzUc/A+LnI4K8O2ZEzQHl5nFHsjDKfNFpTVzL
RCMB1Ehuc35xBe4emjBOqC9ygLAmwdHT8/A3GfF4dzLYE9hZpF44Mb2GIU1JX27Y9po8jaKF2ku6
Mqs4XBYBm3unINLXAOv+Ic9m/Ufk+K0XIyd438d5LyDd7jTLpofvzdxex1ioTdQGRaC+j7OuLpTF
NbcAGYG9+vkHRrHsMZ1gNSmihZ2D08/NKjhuP8tKoBim49Bc+Lj1GXXoVa7ON0v+DEmd4mEC1c+y
B2nfWqGKFruCnGh4UH+YZ6gQGQmPVP/jV1vQqOls2yQDpf7YltHCdfPCk89ZsuQPBEPZjz5Wwv95
9A3OcQkv0i2xk/2BD6q/5KfAY/teEA354aK1PQGaQkcXM/RKdfF5QEyPeoYRgsk6xJ8kdA+GMdxn
RG/96tCgoRaSCm+ivGZh9VduVBwedMPzjG3MoTJ/s05CF6Y2Wwql8AlqgETNdwtsXNZLuhGwLvIv
VGi/2timfBshfNjBXUq0gabQv7VslWptH2v52naybVk0StYBSURPZ2vcoaxwA2w0IHC2/fXNUfQb
N1Neiwq/VrSSvxPH0ONgRdZDzDyoF8k72srQTAdEY8yrjyGHhR6y6/ECALW1dJyEzzGlVO+0OzY9
+/JN3C8sfS+XUqlGpN7wv3jvxZr6CbBL+CuLP+99YvEvT/7iaVHwdtH4inC4KnGx7q0JvcOB+DKH
+Afxsac9o1yTZwTf3m+/xlNLrsL1X962HBp1EOMrV1tRKzscaoGAkCRnzBnIJF38I5TN6/Ph77nf
1R78Ny4Eo+lqXv5gAlCd1ex1DJ3RQHeFeiQQJvaoy2CxcVcBP9PIfhH4KLmnzcH2Qw1Bc48H5uWG
dD3yBEoQjPRggoiqCD3HGxApZstK1c0bkyHwSqIubzAJ2rk1I5+UO2RQwwCzZcgPifDH/fbpW+o9
Cq9QMAF+2NTi9KV1brmqxEfMnlpvX9jTt1Jske4tQ83YQqdG5/3R/wx59lkOmqFCwpvKvGe/V7KM
PAHt0wkPEKODej29Ce02wfM1GUX6jf4eQilJQ0r79BuoTeoQa+LW+CUFS2O/mYbzdUkvTl3a8zuY
5Yg4whrm6S83Q/brd0v7Nyl3Ck+1a0A/bJ62XVevpxGxPM82+gz+KOTB/HEj+FzYfbQRyVmkmjh2
P0+MlEL1oL65VFBPxxIW7GimYB8U+R16oZF0AOFCfDc6sQxSgCGIOdJjaVe/r/J+v3sQP55C7udE
G7wOrGpQ24g2tnhHEFaQ6CoW3gxm65yJxp0ASk+K1d8nt2TozYLjjS3YMFoD6biqQV7oK7FIfovb
EpVDhNHe8ERmP4MWIDBcircrheUBSwSFnl4dDA8WV4NBQeImJ+mCCO7Ewus6+2MxJEpHuGZhn8k2
Q+HhJ5UhI4MQSS6IFqgiTms5WgsYsvqNDHccw2sB4z5x/4osndhycdkLwmShFfHdZX1R7I6s7ZWM
FCTf2AXzR+BtjJylGVTsqMLoGj70q2u5dXiwWODDWZzGrIXOcN8vFsmn6ZcXn7PHG9BxRLWyIUjH
zvaD5NgNwPDF1uIkSTqaNDIXgfh8fCeO+4tFsZ4Z+qsMeyqgL5A5vH4euyFEHidFTBhnhGtCY0Xd
NhK97GbZ7fvYeBKg5HitK8lww5PGb8sF7exS5Ie8daDirlIgT40HuJtel6p7tDeNRn/0ffWTqUmH
wg5rn6vYQx5haqBIF4uaGdVNPiEV5Loo4xtAWLZDqcs3JCRIRB5oNYa18c3wANTO2VpZIRkRZn2Z
WtK/BCAyxR099MC+hj/67UuktnlZRqdHg0F1YppUoqHBoYhy1nZTwm2gvpv49SrbMhE5VWLytB8R
3j75j0iDChiy3vSvavt1xOTijGvwpO9smX3JGjnLR5iHCJz1ttOGNcXoGrNfEdSSs/kXMhDRDdpr
We4X0ze5aqXJ7laz8th1LFqkJk2rdSI+xkNCdTGtUiPKiBkbbq6h7WnHM1kgIp5wqsk+T2u/1MJt
0CaXR+TyPNuqv3e/l2V9e0U4OAtbRGL6g4844FV/UNKLtOg7lIuA053BwystUzDvjiErIBLxPgA5
FbmOwfw+liFEwQ7FMUxq5iqC4Z4pVj3K1ViF7PI6xbvyZmTbpCYEB8CIL+y3Etn3b0uTKQJYDgEB
MO9kKU0jN7BQ31RK+9e8wGB2zsp4u0+G5/HCqxyJuw0jF2WlTdYbpSgVkfSxJJNq6+kS/2TZdNgd
c0U1jxIOuplAxE8BscQidMGW1LQ54V3slsd3lgNJQ56DlY9AgyYtjubKhMfZYr4EzBE5kS/YyJM4
TgQ5J5Zn//SVv+Ye01ooZ9NNOwabqCulNwYRBK33pDO1aXh1abUOQm8DoOSKVZx5PdPvxkby+sti
kylDykcThnWgTbcMZ27sA01Wlq6rgYffSt3ByAVoDsMjeIKjpNbjKdqjCDJZQy156XrxP5Ol+wpL
zgodfwItmWiwDrljf67TjkbNoJaNVqsLbWPmrofkS0KPsLH7EAtqnFBKj1YWEVa29fy+onZTMCR7
v/5MukOYW0uzRIiza9ClXcuXbmSudffxTdw50yFZ62H47swgGz3QOvMHRy5CuX662pC62BPize7i
d9ZVvn7JuIN1oAQxalRXzrz5a5KOmGzrKK6Dncs4Jak7Hw3cePTPDcC4hfZteTYiVmBxLNoUrhJ0
c07sjIEDRg5gWsVLRcmR/8yXTNCkZEEi6e5CE7q4e3aXA5Fkls0iz2q5RiZQgxrxbGr6H+MQ98Dd
ZK2xKTGMSPLKwssyFBb7IWAR2SpPXGIvyPnl7qAroWmlr52d6Vl79w3c63J9u6fQTCvsgWJpS+LK
FG9DAnfZxb7RY9Ga3homNXiQAqBEWfXW7raWlx0prl6WBuBrZdlLzbrqM3AVcXN4ACFtxa5o2Gyz
odbPBmYeALlswcWbO2eSv5IxzpD7dydgjvvq1B6fZq8JJjD6vdxnuw/TRsjkX7IExqychvhm5xWY
/XqMyZ7FGV68C4HzcrVIySsd3RLhAXJti5EfO/08+baE/bsgvAB6XoA9z3GoA2ZQXWTM1XlohRsD
jPSu2hCUiyFP0bwMkkB+S8AlVCcd7z+Ur0Z5tjT8dQpBhYroelkBYleva3Dz0PytqE9WYvMRFkGf
Kp4HVyZ+kB7AYI+qR+ucnFS+zkDnbTMTvvYyKlpLv/tsXcIxar6rpuGHIXtzGhu1oGmR3ufLzFRU
yrSAMldWUNr1i0evHY8bFBX9u2e5AFPxVTzEcuX2wQSOb0qqFxM3P4r7V1Kmf/g017gp0/2BtKls
YwM3d5f6HbZjR4szJSy9HT3a3r6wygSBOwUWVlULb/MR4e5kVyFdogOfEAjmoFRNmzrJVgsH1kNq
kQp4Z/4GdEAOiakKxKFDsRsjcuczgLz1vLCHUmYi3j/fDfYYeKM1oaqY7rqiJSCu62hNyikz3lu+
OOSUIlQpV1Howw7yi3PP6oUHgyAMkQXp+huF12GQIM3r2bk94lXrL1tLFA7tqsY4oxnV299+Xcnp
DnlDj3MVsyDhPcJPZFUPMXUKkycDrQEuJhA/zeaVgPDqh4JYKBiqyeQIeEOPrQfT0pEaF3Cjsk/q
34SsqCJNaBlOIIywNMhLIoqtcsanncPLsvvBheYtkqMtwLcJ/iuDXelvYi2tZTpvJ/Glf8LgyQZ5
8hVoDiBGT2/OmsfOmksHGc+INOWidpHstR30XHeigeZ3IQswzfASPixYA/ShLg/B7W5Js5Rp2bj3
RdTVj3GqnUoZac8Xe7TieByK7Xli/mOpgVj+lpiMuk0xFdxSBkFqkG8gkT655bAQZmlzmgl9ybaR
oHLz9Wwixv/Qjk+I43JfksUkzs57ZxuChRxmAy0CaVfyanLuKm5EXvb+IHasQB3X/+A1heqVbNyr
8r9Nl2JTGyRqAO7zvUfHw6RYPg5JHENE7boVXTmRaP3uZMi+krtONBolwCT9+2zWDaHNKbMFvWTT
8lTOohglnWYskhbag+koYyrORLY8LsoJ5yH3T7xapdayAs7d+KZHoIrMx6m2G7HGjz+SFmdM37hk
hV8jbJ111qNjxYufLXSLVWFBsv8TgCnhzdrTGx2qGQJp3nn2+32rgz6UB1s1OrPeEVpYKNNFh6ZH
1l0k7jPVpqpGt5aEw2P4tmnKa5NDwguDP0bNyY0c123wXvoPcXJly4/iaOyInUIfaVKf7Z3Tt5fp
G1mTEu86uJHOQ2jF5wGEBnTpWw7neK4577vL+1g+Yi1v2xhl/HyyorQ9hD5lDLCgV1v+TkYqB5nV
wifvVNOOzJk8ytAmvr+7ed7ZwXFGY9NDKMKGReX5+axFdeDJQBioDJz07aXubXdVNwGG8gNYfLIE
4z5LvyY2Y9VrKX9dleey592xg9cmeE+eqjsuSHuBFbKSEPvc/0IpbcGhxwHqizpEfmwHNhZvFYPL
g4+ucY/YZTvhJix3PKhWRspPVYEQQJ+ZzsFF/5E0cM30THOS3HxHsWfGlOXjeTOqXOz031GDhOsf
BPB1cDVFDx4OjyvqZitAHCxuwsus3wyYQB4evi79pGJRKZoHZNeVpeB/+9uf4kdUHN5bj0fxh2TR
GcKWnb9mTdJW1CJq1JhIkQDWWhmekIsVQH+fCJoZomUizI+usJm0yD09SvI5xo36CTZsyOUZeWOk
GxQNoT74cv/ipRF3Vx5QntTIYEe8NZJDMzNTXwo1nGAvWx1dKcSVUZIRUKNRvZT1/9KDkbgZsW/D
IdxBf+Nf309C8SqBFOVG1PFDgCNv2is2mw6+k/C9sjQMDkgloAG4G6cADNNHzd8bWoFIWyyIuab2
ZXeUTIkfJ4AHRkr50WBFFfSbErFGSU7BGzqyMGpWrNMZuKfeSqL7liWPFkrwqgNW2q/rIs4yKlvO
q9gOWf5SYusw5Z0A1xc1AjKqKccf6kaNbeevLA9zhGSUyVHuR99rss3XMb0vkg7vU1f2KQYIatd6
tWh6vST9u+S0zkNWNixcjcz/emBMozXtpv8SnUonROqw8RsRRNQmbX9ITUmr8O/KMNbcM6MqLQZz
hqNOip1bfZrTxG4JUo41J+HwDhL4gbSajHTM6uGIodDMFAd4xFh4zq8mcLWWtPaU//hmkruN+Gkh
Oj8SbfqMp036bAAeb1Dz/wnXV5FKvdkAOnb3XCgVKgOtIQXZ/KICnbgs0JK5iUoyl+j5XfdYtK+o
jfzUeRxcgKxWfUPHoQ5jtv4tikC56Mqu+BgAbpTCoAl/yh+vgIwuaVUxVEDnNgqpMMQ04QqpBlZG
KHuoHf8NkRuYmoHbAir/CwSJphMo9N17DXvONJTIWtR9t9NvzodRH87+1YcNCdP6a6oNBGO8tejN
ChlKSYYJYT1v+VMxA7UBzWg0LoE7/BAJsVS7Jy34LRA1+l7oFwpQLh62Ff8/YzQXpZb7DZKwa/Dm
DPDF2A3kQRY6q0uZVjTyfQ3ovvk8M5OOWjcXHQA6uhhuyUTg1D7Lhg+iR2oumNVKWgzLDd2HMMwL
YckBeu38RL8etRv5l/qhp42DQGVd1QayrtIgs2Oqs9VhMRPloUWWiguSzMOtSN6s1faRo/S+ftZo
WxtAm3UdiZ9MTLldBdpBQkVY3Vxg1hJw4kKTk0cWW8cfzwnkSqwC6QzJ8PXlMCAe476L8pLqQ268
yHOWAXr0PjOTGHkvZPC69ij4hOmzAhTNIgScwTqHkmZUp+KfmX7+mTTBtJtZByRCfxmNtPhSa8WC
a691kgP2p3j7YUKlfe66jNhN3Z34SQwt2yjhhfhdLUlOhgYI6+552XSDQ6KoFCE6jA5ms5NtPWVa
kcgQlHWtRtpqsCeEUbeLEQ5U6Giz0MDOUR79IBiZKHZ7hFoCsLn6BgD/GdchiYvud3iw7ATUN8Jb
ywg1yH/f/CreTmRFuem0m54NWg5VnTSi4NaLFPBHTMSEzdo5YdseL33zT9soBvh62DyrJDMNvg1q
wale+oYAyY+fq/xsFTuubJ4cJz32HlfZfj43hC19spCG5ghAyYvt+Jn3whSO0sP04RwSJHbC3IBp
88wfV1cCq2Uqp7Rqwk45c3GAJLza0Ug9Tdf7bVx8Y9H2xuC9bwR7uG0y6yZFI2tKBJxT4fWUC7di
cgx8P0gMzCyebl32fos1rp0xssW2xCTuuG1nemmrFFEpsDQfhM3Yx0ILEIY9Dz5OIAS+yhBjRIMu
8HcswuNDvEoaY6d2jPmPoa4NgrZUJCHVgFWtt9sWpE4mBQ21GT9sfqgrecIzejMi8NoN9vXxEnn1
B9zSTGXd6WN/qFkmHepZDDYyulyEmtcW0IXZuJ6iSiRyVQ8JAgitb4KcqWp71ZmOtwhiMP8lCs2m
bRMFwSgAFH4i/+PHiZeGb/Zdjo19sZCXSTOD1Tfx/LHNa7sy95n56N2oI+ds5lifAuSuUExEZ1uI
BrBspTYMTzl2NlKIRWRiPFytRkOAx3AZwMevWejk2yhXWPcnHZoB4g32EYyzaTqk2nqwTO12uP8/
Iz8tOeKz48Z67O5DiAoxCf68k1mvnXzZFHym+vAx3WfhQh3goMoam7VMHENuvtyE/Vg8j16LkWB8
cgIiLm1vP7klEUxSvbOqxtxIoosAXE3Igzc0s4Nvt8NRzAC87mDZ+Y/PzMQPUb7PBF9jrO0Q8xN2
YedA6gC1R+LQ0Hfffq/n2QJ5QJ4vffyqchyHE377hJ8wNRQUZLogXCECHpF9E6S3HEcMg7RZsuLG
RPUSO8IG0ga0Sdrzaq/UjqivfsjPjXYhflutx5jPPb1aVVzdO1RCu/bVSfddzAVOj2D4C2jqUrZu
dLwwnoUB2D72VHllFhxNv6dZLXAQT6tR+FZ/unBZBbNyUyxu5vXUntHnLAjMHtOHfm2whPeMyTPw
nJ92/7yIabvnhxQr0xTifs3Ps3fARsXMkNaq7ewFVV8ZV110AyWi8+0aqVZ3FdLgs4wnKiTTURhb
M3f8lCg/crYcGZTh7x26cZbsrH9aNB5oQrpSARiWb7ikC4v+yX4YSY8WusHml2MO+9zx6rBEjX7n
nYbf0814+sG0STawKFHpAJ1ymWpNqkEzokhOBH45wQ49D9IBFmAjQSIrf5B2gr6FcMKySupbu5xk
jDYJHCNMD2IJ0Z+CmfwoaCYN7o6+yV7I04T4x92x9qzNrdtjUsxStwChF/j7UC6ayZI5HHGmD1UT
Nx4388R4I96ymfTC3xxn6d4fm1VJ8kaTTnOKJVMzGZRF5cnRG3lY+DTICTXkyhmABkL4cusizsDY
IiGiTeQVnXIbRV/MNe1DZG7OcX/QdQFGfQqzEZEKTZWUNaEevTdow2MOILXBF0h1xxPyP6BMrNXD
1SkADYLb3DSPlhEZBWYIcKIe+APpCZUkCnJN3+9NrE1ApeU/XZ5YIbEZrDhaoGbf3zHNVrU3T9h8
3xifquOy4evXo2Z36drYKl9eFuqYUHm8MdWgNZMmbYOmMxeR1eqhAn1hV4+DgdNpIKQm6zftFOqs
3U9WYSzEhhb7t880LSsvqGRkvDtPZ7ykAx57g+2pnFmDClW0WxZfhLv+WNRq9FxLXfpXdpeBKaA1
VJZvA2TpaVQiBIG2yUpY62k2Eka1wFhBSctaeM1oCD35zQjaxwOfs0k/sy5ddoah5PlyIU0K4/nt
II8VFRdzpNdfQkU9OxiaZlschy97z1OVvZufQtpqzYgRMYCli/G2NRcAFQc8rE7tNXLeRtv+Z7tb
EGG7owxxbwnP0WHNmJn8jyA5wBfw0a7dFPOeYgsjCvpiSLU4IjeFz3cQJ6873Zbj0G6IoN054qkM
0HmWdpkvNV5dTy2wHWWMBP2zK48VVOaXvmzxX39ycyv8/BLOcshiL91jQnrNmYsdztEPVYfJdlZg
1Vlu7g53bFPspNjOnej+ECaH/tpDv5vjdkFUGWyfJh6sT4Fus+Z5u3Qg8w6iGDknzGwdxxq7kvEk
hv5c7ywpE1Rm7y9TjpJzWRixV/jaDNc3IpOBGXLNfHO3LtyKs4Pnohvf4vl7EQIuuqBMsRX0MFLi
mu3Jh2FDWmOaS1x8XRkC+OaDcMMQ8fF1b6xmPZXJMczrrvRUdPw/Cpmq8y1kJaC2KSFaIHccv2Vb
/DuLWFF5MJEtT1KHn+rwpfzGI1V1Kw83I2FaKlUP1h1PXd4ElQWkOZfbe66s/U1X0OoGyRQwh1iX
Dh/qzqZmxUz/71jz0j6oWQzYCFUHP315rn+7GHZ7VvVlYU7Tvvy1AD9YA2N8i6iqNB6UGXJae+OL
g/yvaJkKaP/ISvZJE2E4KlrkKVuLZbvtCUIx1rgGFOMYs04bybJXNaPdmiGv9Ncof+tNxkqetV4i
aUojeqczudzxkYOv2wHXrkZmeOtS6DT1bLyCrjeQosrLEgLekIY1uuAlIZ670UX4IoS8qrkIdEBn
06V9H5vEFs4KOEVnctR2oaSATBFIZv9KHJktcJaq8KQ0Bf7KKcOh+aGT2uYGDLHYDyKBL+Ikw1KS
ePlsEuAw3w6qIrwkZC5518/9i4tnT6sGJJRK2ipR75E0H58mnwaEf9wmyQwrtlNrY5/03MnJEeQs
YdqaCSnMm+xbaUn6zKY70irw8TTO1yH7ZCQp0dIDuuBb8I/bit84mHDmVxATGMbz24CHexs2XMG6
mMoptUFbapZcRK1i+kOIZzxeT97egmi0TSU2uMx4lRBy7me8p3iYTR5w5hSsH72Y8twRB1pVEv7Q
7I30W9k9sVyrRhQre8mvAQ81zqiR9th+AFuG9J+G8nwGMCOmkUJxQ67pYRE6pPhMZI0yqCtUUDRe
tO8VV1NcfBU2WkY6hpJBer4AwmFGsjJAAMS9CaV7+fOIyjHL8HmDOqWtPVJsDyfwwY4FX4nFYO4M
gMPPtxxxfpuW032OdPpUlcCJUJUSA+RvqK/gNnqSdDAToNMR94J1fD71HiS95tFGUkuwWdaGtI7u
/tH4pUkHl2ccPJ9e/pr1CcF3aavZOH+kxG7K7vqjqHfXPEd/F+HsGsW4IcHvN6VefeuY6plOlWgT
q6nhcOtivKacWb//TSG6SX49Tl2n0mJkwrj5TpwkCWQ2vVGs60UyiaIOGdltA0m7inkElIhmBjcv
2f5jS/B7ij+EXjnPkQ8CLN1YPiRqq83EguFBZ6+WINDp2562xNVz8477+mX79NxKFbKyUjEq5EzX
5PJTcZdA5yydIeg1JqeToebjvsO8z1USJZm03BK11TYgERHk5xwrn0xJL1/TXOz8stSxPqiOGesf
U5qjecbIejnXf6oqc3Byczv0BtXqzKuzIPqrPKqMHjwtNOYKS35q5fYIjxYEh9omoxFKVKXKcFx0
zgl+8BCxbIYsgSp2fxjQtQmIWb+fHDIlrglnuJ15fuFwi/OwDk28JFpQ6WeKBtbjaAH4Vaz6EQlo
Ia14cgPHqJZ9R8GqsD/JqyOc2z2rdm1usRZi+xi5/SgjVwjA1nPbDg82Yb+nV4TM85Yacr6ioaaT
ZL7vPrt8CS4a/orXjlXP1/3vMJZSRMzHgLOPZ+2fvR4xqN21wMEatv7AOKl4lE7i0j49TAZsGpfH
cG8VFH2v7vuTjmOMg+QacnA2OBqFvo9PA3or3R3uBlmJhHaHhkKXbKqyNvGrX6pdWtFLeBS00exo
nCr9PaDIe08fc1HBajdunTcqEhnHBFLvCv+VVbuEj2btRViRujZzpy9tkhnzK78yOq10JJu/X18x
u5Unc8yfvOEtx1rxGPoiGPJD0tMLGJZ6LTezqvbRF8JGmpP6ydrZUYIaGS1gGJzxx7Ax0iF59T8h
rWO8ed50epqSGXSQPGFayE17YapC6K2B1ocVLc0wEB4pfTjdlS6AukE3x6SUTocNnvjexzzzi5cF
qXLeP6JPq2czEbFcJ4346BBwt7hcGEl9auIANVT3EhLqqNUzRQIHQBwLi4y5LGCcJKspHa0fcRn/
UVrK56wv81Bbg+Qaxz/VYMxZC55zg/j/BEQXouzgUe5pXwn/DsiJj6GZX0DfEoJhG6Q7LIRh0IPP
LRiMcf2jBy/WyB9ZSvd0On61eI7OOpCpOTU1kEwjYsMFIeeaPU2QVaSyHqJZS1QGWa0fufl7bY7v
1unRb+hNfhbcYUKS+Y54hy2s+6rNenhIuneQfnuzEZseQjIWPf2Z1cc/lOvudq5AZa8dswAEUdcU
2l6h84A24HEFtgvb8kSpne2NuvCuKWyhJbeaQ2+aP/T3Mku9w7yyY5ruCyCvVk8Cg1UgZwusu72I
FQgaGDubJZ3u2LB+vnslRfVoe9yKrxawO5+qfsXlNd+yi9xMq0MTRgb1rXkeQTGagBu0RzCIClDJ
9tCrZcvzXD46MTToi+aVSVdsC7Z7w+sKerJQaF2VweP2WQVC72yalSesQKTd6zeB2I7/Lv4IRoi8
55V9iBn+YwjTLK8iRohl6K0jHnj0ZNr6Xz5TPac2NrLUV/7kk6N5fDzGCpGpxeDlIMVuozk6iGdS
1y98StU7rwy8Es+Pi2stf/3sfbC11CoF4ltPpgfx39Zmnzw7ukr9T/DDQdGtYln9Z8kUM8bVS4uI
qMB9gG9mHzhmHdptweez/N+TfqTqd/OuEq6i54UkZ8wTs1ajg9zNGlz1QOtp+6uc6EStba7I7ggy
/8NPb4ddhmdvPEnYVizinkYADV8I/YrpdV0iPIMgrpp4NzN3PhlQxjvTtLx0e+R8tJTuVqtUIM0g
wkucxAR2QSONC3bhyVCwCAi9Mo0hzBqdti7EEVYhcJnAeoWUbyEdIjAubqTKO7/pF7X9atyfeoWJ
mRo7BwdNOpAe9/qS9WyMiM8DiJbzM4AsHolUWrazbNXJPwNaz9nlXDqgpU64TbksTk5bwhwme9uo
II57n8ZWkZcNj6iR9aHz2VbfyTKFksnuN6AXYzEs0QWGoORE/1rEyHrNkqfPQy4DR34pbpp3TKN4
/hB2h3UnRjFWrlxEXPQWlnsdF/gezxef67qpRa7KcADUAm0UyazO/4gWveZaD2eSv5siFDdscMQI
ApfhKenWe4Zq/UU/TRrUBgYEAuYQyvK5N+NTTIpYW49LGEU1PFyZ6KyBVYP/TBayQp6Lrry7ne+8
yQHWqyZ7X5xRkuKkNcEx5Ab9A7oUz/vKUv1nSc48Kg9LG5zN9rj6SICxf3Z2ewlE58CUP074VE8g
qul6T+ooF8/RRHoQC8uu2hdjMIAOESknL1U01mYe/793qms+qJkzfP9bk/kc/60CZ/+nEjYA2xTK
enwlKWL28Jx7ukzVVkB0OJxhjgUfvY+DxtRGtxDTJomudURcrmDcH9nWJgpMDjQ2iC5dUz6fVTZ8
SVxE0yAlGLajutEmu0wMLr7ub7IrjwLshBETAFtD5F41TpQRGm4tStG+4JWYXYiwQX/79N7LgsQG
JoQjwe0x6mxvT0MSTpT/d5uz7j43cLib0BMqrqYoMQY/RYh9FqKakLRkbqtQgq/9BN9hfy+UKeEs
sIK7TAjN+lZgsknE2CTRnYfDNpj8eGB0iJcXIz8EXYdM44PaDlgNfOPpZCYiBKR8LT1oDZYUlNGI
FfJYqaH2bdZdmtxpIxEWgIc/Wd+mC4yFoESL8RwtH1pikmGqcLpeuZ3cEcbFndmHmqQ7V676kZ8Y
SFBjixqI/sXJs2+mz8Yd8sXv+NQhXPsiGTB0FlxfgJQLLEWwXeKN4OCUhPuIl09VHvrLVNAW1plz
7RJPmWkL7fZecSZ/NoS3lhLIEQlX07wVH0dgb7NVAxuBZ0z7VR61QbpSGOhDHI5hLphFKM2r3UmI
1IaA83tDNnIy/5FAGtuq2m4SA0tXE1QgdUYem/V3NeAb6CU66JV5o1lUOwZcxJXcZTkZ5J4pV2ws
19F+AlkDOTiUAfrDIsNLjOXBsx9uhreVoiZKrHuStx1XH9MrRP8t+KmT3ROwC/3QNxZ19/jpHQtd
+xiIhnzEHStejBPaZL+8VR8UYDlT9eDn62qzaeF42MeEQan5f0JEZnEArUO3cLwdDcGTD9wTUsVP
6+SroLLZX6uiYH4cZHboRFXGo8dmuypFvYDmBf8+yFvlgsznrzwgoRd8GbjVLcpI9rqP2WAgI/Pd
L5Nm88MYL03xfb15Dd7XkiKfK40+a2E4z8Z/qhXC+NyeO1YWR9Q+0X5rBWZL07wExdgL+RU7+KGv
w1DGOkPlvxJAZzmFYfC3Dpd8N3Qtdf+KDQEY5Qg8DJhd4r0F4729iVd3RSJgwcsazeC+RmenpBoJ
PNuuuwwgrXc051u9GBajbjsPKge2uC+92kdAoHHt8u6GCrFLm/63JSf6Qw5aHu7SngPOVr6fV0Ub
5QyoLxHT9IdAbKFPxxmyDAX83w0OLP7NQnaycI2qpNmeqxum2HpbFzFL2VG318lvMdtqe9tMoZ1m
b0GuzCIhlKivaNgQyawT/VB6kMAtHeJHgTtI6v/tTFrZenKH48/PsabVtUHGBhOmWzH2TS2vFf6d
kt3Zi4935YRNSLgpOCw9orEQZj5moX4oLQA7SOX8jzfKT3yw48dxShqDMFi/D80zwxOyE7ZesTQn
bvDsTIryV2M57M2ZrSPCvhUt2Govj/Sb+glC4KzSWSfEzlYtSPVdg3LW9024lMVgITwvuGhwiVKW
JADPAlbhSUT4y6TAH/5d//n/auxkdutDkibT6bpzNpcfXx2HQK+cqHkQ045eN1ZVVHaHEeGuNvZn
nqV6djkzrzaSbrw3fjFvW5vKHAU9pv2cNYVEHP1CrUUTt8NdepCL9BAFuWunV46ialkMZZN4JBT9
NDqoQhnwkD8VWsek2yb3os13lQKhPTrRblJIMHkmuY6rmdgmjzcq4aYhVuGC5+qams1YiHb5xp8K
kM06BMcCT0istkYvjMjCLaz5lACQLD0ugLTkF3VA0awoLsyHWejR/Mn8eEoOK1ZutN+2eutvrHnH
qj/MjTB+J0epfJ0wmYrc7sDnm4ma51gcVjLph8Ky8l/IJh/RchhThPG4jEI6OqDzfUMOVuO04iWc
+W9rONa2DphzuqxJrLP5pKI7omd6+QekaxHwg3UuKg6RqD/oupS/B6yeaRCaTEvoLws2R3aZPljv
GfO+HQfkJZM/mITzOjp3GXkqZGlKtR+xUrgb0a9xo+TZJWAD3Wh6DE5O/eiXXyfdneowqRyu5NYe
WSBH6CvnoounIz/iKtwQEpoZG2Kn5ttkknU5T02tc9xbcCzzs+Pt2mqMUjLcYcDy4fXDNGPfveWB
WsOO71t5kQjrO0iULGvzLqm1rtgGMTm9JZxFQmzDOZy922YLbuEcJo8aHlNtdryLY5UJ6n3385FD
g2gn9/fAFCo2Fu7uIVfMXCyLU+bi60jkHVP/FHyVnZjnsvp3pGuSZXZxa7zTSLmjWKHibSBTlFmz
7tagbnMcmU2dbsb3r2AEwoJj+wEl5gBS8yzJ665uINVgRrdZZc6Zg1HMoP6vhUCXOQjz1+zXMb1t
U7bH8Xk3Y/U8bjqKtMwrDvHqqL7S2ZYyJJROAUphHL216DxFB5rDNzVDk6BmuZg3GXwPG0nGWtnx
/55SUCh6GSdK6vDoawXK9gXz0xxh7RhFO9BFSdHMfFDV++fMcyJG/sZAOF5Zb7caIrumIDxEtvsl
Dhyxp1KtzP3LANUxc7szHdU1bsiCRHXoYTa86ro5DG4ddaKHF+fCoJC7Yny3zRULxiJcvBpGFE3L
ZMhIV4IrTnosGgPo1uWIzwdYjrhnw2olPAJZRaK9xIqJw0tymYoh9XN5HkRRNcG6NFfmkUri4Ti8
slgiKTuokkwzqS7Q3SV3lGd3b1th+26/A7hadACik0f62Jo1ADiotq68NEXd2Uo3S7NmIHrlfCsS
cCrzQKtBslDkUO18WlNytKETU2GlUbY8kgJIqP+fizsWF4NBumNUhafbEXyuNZjXuRYiB1Dx8dtw
BbxpcRwYSn9YHj6XnfbqILThC2FGZLY4TpNiKxH0XhZlHruhDtKFZHNN+2b5vPqOxhSSQtVPSCFk
drZKHHO+13r9p9AUi0ckW7Iw7Xqhumpc26/fMbhN2/3f4AL4N0OPuN+SJ8d1X4IoigRHIx9eWMe+
yp24SC8mvM7utBsyErrvxOdthL1AcMGuJ/FLqZu2853+yyVKqTt62wVQDUgJIRgjzkoaovU/xyFg
Y/MU1nGLOolfLXEpUIQrzFv3GnYcjxAKM/cdqVCKalSohzyRTvPZJAE8wgETWq0Sl9NrjPau5kmt
TZvUg5lUx7XtKrBUtx6L88pjTISxp1T0HDLLvQpMIx+prOrvmeD8WwOXK2Iu+TTjPx+yD4QDDO2/
UMZ4hxraSceRxhOdxIWUUFpAbSiX2PJfVItg90h6ntJ6yMukDxvBO8YoelLELlG2GPDXRwpLT1Zl
dxPMLZKuboZjO9bJj2R7iQ0J3mpCBG/38hR8o6Q9PziN9M/JR8n/HNvJsoCXC4gbLQyinl9Au6FQ
ffV03oiKDF35hiwWBYfk897Q3ASuGveIaczM2VaaJa9RRBzV5SDSdiUtnVbp3bizIk96Q1q5u5kT
tucnVUvYgt9ELBN3/bDM0MKb9OfIZPDUWFUPe6SSbIXWrY6n+KEKz4FFhpuHVD2mnyionVc/vAnl
/6N+OOniKlatXjL3WtUkCgFBEJ/sb9hMQ7Zqh7qDx1Y+9sjWYuvesVpB/YTWaTu8Egqa6XKIl4Hf
rvBcssGj3iGCB01tHo9wNB/jCChY9a5LYZdRu/COWusxVAdYz03M7jL0uyQjmaqQIwxBHHvsB16T
437eCh9bufmB2ce2RmcqJ6F+cusS+KJhq/76IEubEtR22goDN/XSCQWzXipeirJppNr2BddeqLwk
it71VPubfFqFVZsF6Hm0hDK+Bz7Ggx+fLziZBUfXB0ydUa43C0OXaK+PIzDUrlr4wQ47CuuFDQDg
Fskv6DyaP4y7XyoTBwFZ8OL+S049T4Dd6L16hG2TT6KM+vWUQPPA7igCLCUWfIXK0FKGvkIx/KXv
TiuMiDOHDaXgzPSMzXxaGxbWPyQntflo7O6gQ+yehi4wi7UBmfTE4UCu+iM3p8zY8ETBmjvoIMDT
yo6wJOT++uziXhKQfBeGHOzvZ438yqrIBc3LlV1gU6Goc2eusxtXfe25JePmQYCm8uXgCq7poITr
MCVaXr4RLKYcJdv8HDckMHuJTRTsjsZ+YkfMUNe9WpPGoXMSZB92FB29nSywq++YGalfu5wNAoiz
3JaspiXXmZUObac3njFZegxrTKDy6x7gxdo3e09N6fjJHVNNKvjWv6Xi/MV3Ub35DnUPzet6dei0
MJDdBCSnGH5n+ed/1M08BmrpRKNrt6XfRblTOOH78mx2C+djAWcLqWuCd/6BySluaLDy0jFO/eJq
PSHFOKOsDaJ/XCJIY3Jv21lPFb6f8mFXNHrFae0ottLYZ3VDOukDT07Qusqxef6TtZAekNlXELU7
QcLl4Su6ZnPcPn5ezkv8FXWJzNloD1HPnQsiAN/Pcry/kleby6UDR3p6ZgW7uTqdXIfGOgEIsLjD
dIw2btdJTWSG4vf6Z/HXHi2sG4HXYx7peq/2utaCGp9147w8M9mOeZe4vOVHOEx60dBmioXX4QWR
ChgGn7mb6cK+fTGdURz1hTcrxKpXTZCfTbFXQwwn5NtWt61OWYZLmfiy7QQlJztaFRBgG2F1m11U
wG1pl2n/E4Zv0tp8qxmtO7UjqLwk/gncnOfmS/Qxcj+fvYudQsJoI7ZoaUOTpBsusxbLQ3OrArpb
IZ/WCSFH/jKGYgolTUjcXVwt6KIXuhgIEktwU6RcrIiMzUVP87xbgfFJmnSywNMBbF3M15THu98o
uF2lExz4okQbfo6ayHDG17l02BGr6ZUcY8QdvatavJg7+0AzVznb/RKvrkev7VDNgDwlGu9MGzRX
J6HGDK098ZS6/raVAuAQsmZ33yoKNcRbyMpKdanRlsSP12ixwd/8pW6ZJ82kqmUZ7r+RHfF83Xyz
tFwVPkkhmKigu59SgelqnRdJf2hfncUJP9E+vYTKaEIjyY64Jf0SAfcpELyxsWiQdyaZK21mkcKT
ib1c2RubIyIy5fWUUe8nZP29vdLZJTdNlTvMPd0qjaZUhEF1r9tO6Gbd6RwlnMtynYxYgxGZOGzH
w5lwS2H69O6Hs3hxgI2tcoO4xifULaJLDHaQQIcrCUbJ7kyjN8ybEsryoEXLFI+b4+/eGwVDwj1u
Bpds60BYs19jJhN83cAHE5btnflcXB+OLS3rwziSNiuwsOcaVwLe56zMBOkFjN/WzYxsZGb/s0zq
xdquEEEvNJfdorRoi+1vrCC1eWM70gO17NVaFKxaRZazvXVCE0kyPEgSEE/tSFiskEynDxug+T29
zQwEcKiERWgBAjDCmicp8RZRFUyfyO33Gr6wBXBujHqlMG6yeEOIKrdKUAxqWWh8tDkW2Pfb/N0L
5IFOKcgrWVe6gbbMDST44dASv8EFqOXG4FsYajrCEjBXt2+FBSdPX8YrEADg1Ynm9dxfXyEtOw9M
0u7n+6G7vXpg12g9/e2SBa10HOueP0W9zThqYGNzvwmOD9kajJS7jcMDiJWB/mUzGhXB5ElpZul0
kMTC0M+VM5ts0XqwrOukbZuZjw3hXFhK0t0mToZCv/jaH//LI218AhGLskAfr8EFXu48fiZk+3tW
5r9iIb/6fcgIkkrHTyaT4/WrbyvtdzCj6jh3xU3jnM0Ezplpw7kiycd60nrtCRuf7FfB2GGEHeFO
dxnKyJJG8SqXsGUhPcBJKn3jI7N/XUzbLcy3LSWI3fUahp0ZjPo43LKJFwKAdpMEBnWNsW1oE9J9
QujSTWZRU6ZeHuzu1NKhPon3aQmwXzPBfrR324yLm3YYIF6tK0s5oqdQnM9LTazC8c2hTMiuWGl+
O1CeIYBKzFNWT2QX9QRogA4L8hD+7XOYuvu1FK4s31kNq8diDACwhh+8jw3odffqgBrQBtv7T6BR
N8UJnY45+Slx5O+4/K4xL6+t3GWJ4USYVAPN8lDgwq/bptBv1YaDM4WBLtUG2wfPNZ9ifYFTU1Dm
g3o6dz8bC/hW9Wc9Ta+/w4VAQyrC67GgBXQMgPo0LuWYSLk8cUiuLcmt0wRoRWrGuvR/XAkfVRIV
yYRlYf36DGCA0lLOjUiR27WEsj6kVJysWoqcrjmvvjB+NGMhEnzqRvZkPF1T3jkbAb+pVQ5n/20d
CXvv0zXo8eGbg/HqdyJp5/0tW1XAHsB6DC80k69tpMSIfgoe67fgO3dfAPHfEzwEhTlsXNz3EprR
rDAei66O2O2fUt5mlO3NDx7FsvYS/bl/HllwgoThnXVrWTUJJd+QeyEOqhxTdbZC5GGdjpWlvk/b
4uIh/tyZnRvXqk5ez+38KTQ9Npj7NgUmTdoPbxlygfdUBOCZySI4riB1vpbAlgqNVj6U8oSBpjfF
LTN1tvpSHyJI6hyev7GikiHt9FT1voBmdlt6VCM2Y0VadFyoSF9Qk0QPPdtG7VVV3vtPBMA7GtUi
9m8a2nHCt7CLM8JA1mX/QZInUsM9z0vHRVsIq98M+61AyodxeibrOmawFYwkdLxej4F+kK3t3zZp
H2TloBSvSg5kKj7qZTVd+N83un4+dJSlPVpi/lLowLa00hPZfu5r+fBmHt/o/F0j1OKVronfMj3Z
FABKCiOK2eDwXiBZ2IHfBtCBK8i4HePLa41izncvOMWnK34fnrDJOy88AU9FS/GWHj7g/i18MGwG
+udxq5T7ARJeDAAcpqHNuUrfNJAY0Hy+cJoDgaejbfQodKwQHHEUftiPzTNlWn8dxCVeH3gcy1I1
PCfcmk2Pm7+c0X26Pbur5O3ekKathy8Pznyn2GJTzAGpOMsZFlnM9FrynMX+qBobuXnsGDXgzF0p
aU8W/SnfejAUVImc/9y7Bazgsn7+kZ4OFkEQttNva4wZu0pyjsEM6Fvc0SNWeDidAlhRuGRdSrut
t0Emt3lYUr1oJhRwpd0gJALXhBnHQdL4F4xgnOhIvFBB3VInCYnsK1LcVdhbjD7DbViacGWT7Yff
Rfr65FjQTJGosGMhGcseo6WxH9bxfh1tykB/Lf32Mj9qkdoYZ0A5kRPqKd/yEu6II3/uh6iJ2nas
WaqG3dGvj/qcT5rzHt1sJ5fO3VMSlcbp1vPHuiw6vdRnb5Bt9IF/DLK0biewhJx9ZoXyM+3mVrkL
wg+Qsiz8kRCs1eFABKmcjHfo+Z6In28SXktbrM/YGYaBKgGw251CNjsTKWmb2S228zLUcJcGm6x0
yQVVQz7HvLZsXeMfPmDDTbr0PiOo7UNgFYVVdDjetldQEiLoYs80vF/Y5Hjx7R0m7OlJ77F+HZOh
vyCGNlDF4Yp+4e2s03L1fTT7NtBcgjoH0QOyaX5UuIeW17wvB1fGFoWeM4bLI/39zyai7VO7O13V
y3m2Lb4iZRvGbkaq4t4FD6OYasVo6BInoxhhxjYoCvTP7q6KgdeBy/dkN4Cis77e16XWxj5WtEuj
oUcD7WZg82ll1211IwUmh8m9X0+KU5Vc+GaKqJbs8jHOiYAB7Ov/duU+pt/ljsZUzn+aHLZrDIdt
mrklLWH2uDN7/xicdC4+coGpDJiYZgR895qzYMvLIGKLYIBLOSz7UucHcT1voJewVrF/mu/ZCtCE
IRb6dCMc2a/UqGNHn8s040Xa1lW9cluJa1FZgoezFkleGvBBojsKbdDAr/yzIatn/3KrNNJUZhgw
rHRHoawwmsgQRiccnW83ABWcvurcpcaIJSJ/DdwVRRNGBYVA7Mgd8EnlSgMEqmHIVsVqltPwO3aF
T7eSVi9UPPlhuoWH2Xk2POTtPFXiGWaIT7gJ6KUOzkQZ17RKKT6XEAU2EKhvajS/6FEiXGmIAHU6
63Cu4Sp9gFFgAy6RNFshkmVcXtwogkQqrOfHihUeePGUNs7DV1s+fB2JMB4oZy0YMvGhNG8MwZrV
JwAVzXMBai00kF0YmIf7BWfSb+doM/adaEN0axt2WmyRwgcJhK1hzWrfW8ma6ALtyQIQ045Fum6P
yShKwpuBtz1NJPi074sd4/AqCdOKENGBarlpXo95SDk4bO0xqKd7YtgbSzx842Dd/r8ZO9RTfax8
AKzdB4iWR5ca3xHI1gpiASNaeHUytLCReM1nP9YTfnuWdAP/RqnRXfubxlfXDridP4dxIHQDr+vT
sXW5ICQG/Nuzo8mCmZ+VEr3SuXzopC6NCDCz9xqaW45zRSvmDgByG4+5HRM0kLirMSURNkbx5KME
iQbmb4PmfJWaJr3oQyrYq5f8UKVbMXgDi2rglqTeAXqyE0OFXgKie/WiIhlyDSluitcKIzvcVnvU
znskXbDR8+9fhXG3Xq17E0HEUTbcgzaxnZ5+/snOpvugk3DVxAHSTyyIv3B30rIi0LU04XYx6KZM
DUZaU20LhIGJyWMncsU7R6/zGw4aw5PaUDa+CbhPyz4fm0kePN5XIJxyHT3OVrZqr2T038aPu8BA
yrtqliBxb4Vs1arrpmg2msY1Z3tat8NtMtk0lcBLIpE42PFJkgBBPfRbtGQ/rqkwKkfedp7gAE5U
q9buY4g0yCI7cmkNXIBrBo+5axa7dMpV6BC9C7vjv2IUejrFwhV8/COgiWpP1LAffNHkp00V9cn2
ow8bz4i2aMImpfhGhh1wa/xw8muM1Re3rc1p44SsL3858Q5zNI4q+0Z0YEE7yAJE86+sFeYtCKAA
/yktdOgvAYCVpMK3KOtM/ru/EcAdRTkCPgI0jAqNnmIYbYNkj4WYHx969I/SSIOzhP6SfypPcif8
RwvSYF8LYj1Tr0Dytdd0F59hvAiO8mjtqIOEsEV3H5OFuND1Lky7ZIAKq+U2x2F6bSN7b7Le6wCX
FDnG7eA+H5mMMKqvRcbyCiI7CdsqvoSZBz1ix8ivwM5ae6hNaC/Ht+o5cr6VC1l6/g0xcyMVui/Y
0gr0EzEiz0P8Q66oJuMZWif2C3feDAnExObfvSvXYIZ8utJ9xRCYzyeTUN53YfADIzq+Ha+EG5CC
hLTE+yQvw2XEDuVFn6tXjUVDXOJ3ZikVVP0dBM2y4MzajLAQyQPy5IU17rdv31H4GoCEFKOAWR0k
hnMnjnRc7OtfQzzWHNg8ODwmJAtmS0d2NSOrKKYn+Uhc68wPDJcgmJR2JaqanGpkh5eZJGQofFbp
EiLO2nBE2ndUd0ItWaDt8cGfCX2SnPtOZ8jt+UZ5E6OkPHfDJXlsHffI15qVSTTOaKdHQrU+HxFs
Y/FqYbbdixV4bnEkETqwKfWScX6qRZ9nFmUL/XhhZnoaL9Vysq31Fj2+75u74RR70MCIkdLkpnsv
Uy+15S1hr4G7sBElUq43SwVY/HcvyG/wNavdbdzEi/23DhTBJiWzFGABDsGkpRH2Jf+eDYcBXIeg
fOYACXrVaCuiyvfydn0k8vKRD+f1NMm9gCHJ1ZH7wtoKaMEpxyTl4GbiVql5pCM6WSdT1dpAMns8
YAgBNXulPuvYDWX5yIjIpqwX3lxakqW8J5qeRXaYBUN/6xF9HSxM1bKLU3DXOKy8ecEXyhcPgF02
HtX+0kBXR+i4FbqmlF0kJCfrU++kF+xT2O9tMNl4BhFlb3iOEF+d4VQWSYXlvxiy1wS8SZx095wf
QFlNyNLZkLsMsFSOIoavkqKMfGgZVL6IVLJSaIZ3F+RthuDsPkUW2ulCiU21enkTPHKA/PBdtnGS
BeSVXfUOL356GzMYuNEYFRQa07EWFVQldZ5SuYvfQ7AnBGaJvrHUko/SLdxzoXt3rNGBXydDtvgj
KbVfqrUae3T3Q7qozmyWU6tjZGerro3xp3UP98lcP5gvtkMMfKIyknyAOHkVLQAuuoqQXE7MAXNt
ZLiZEU+BGbA9RvFrZaaDkJD/vp4pii5PfiTlj45Av+1RML8G4i0w5MJBR4SXYolbZxp9WKFkaxsT
IDoPhXv3Z1QfDpJ69A1TXqYpgLnwlGzExITWP/Xg+qA8oJShrDK1VtMPNrobGbG1TSqksExpDgKf
NJDuK+pOQp1pVbkRwhUCCh1tEGey/wLCRRJ6Hxesmdla0jnMPStdeZOpk0Kjx/DT+qn5wDp9vPw8
ug/hv0XTlpHyLf7IxQIHaXcVZ+F+OkhT0XxBKtnvQty8s/UcSUhkGgS35mRjRlMEkO/rMBH643uo
PnrExNoAjEi+IrwOBv/WS/3UqpsXIUdu9rZ3XZpj9cc1DPN3+AijtJdprb8KbWUT8p9XBJOjMUoZ
Ao8PmF+pK2kIJ/8+f+/FX7BoaUcBJTwhzGkp+0R0QjSwsUukLf22r2jHlphT2UKNEVs0+yT+uaE1
wydSHxvMbQDLX3r06HgB/FvhUjQuoVFcNuEDVnMxwJxubiZAb4fWZNI55QiZvwuPaFSGjll3R7Lr
oXvTtgjys2CV8cfdYNTDAZEOHtZts2BdX0O4s6Tee34SHZE8lBsWR56Ro7Bcdc4owOrtWyFJBDc5
gLGfOU2c85oSkitwrQFUwmmslqQOrdsD/Ayn/mOdnFOEtl7GFQ7kZ2mRaJUPMUQ/0izIik9pF0OB
pHIAVQfDcbMAGUtqvPksqwzfUqpka54F8UQP3DTUWpxtSG/ZaSDfS2ZTUSh9julzU7UYk+EOvWHw
geu5ArfvJUnGQm7mAG8uLsblN64ollmMyARgBZmT6NSkIGzYr9XSvuUQ+MWPxGnRgRR6ZYnfO3He
rNVZ9sQLvEHXqWtG9II+0FwCp/vL7dnz0LHNNBofGtGVkQrpTNhTlk8s+jZYUy/UGaxIB1lRvlD/
UXMP5iRTbk30/yJDj0X+F3VS0JU8pqkGLqBwOswvCEarejxNumRGuyHi90SrFj80a78Tp70gCQ4T
ALZ3oazJfaEf2KnI5wVUpNNwrt40z8v1r5VMdZ+cWzvp6SvrfqW1re35Bwjtz1p0zmwmNCI1ZOvz
1lOs6nyKjHgbyliz6W7yIE/jjJe/XmFp6USAd1EuqkE+Ct7DQtb/TMafRrO+wINFCrj7hqr+AzO4
9adcKOvKUHQmld3OpKUF9zPhVT/cDMQA7UKvSAmN03Pr8jZiAGvAqMr/cDxpFUPyD0Se7e0S/LmE
GgkcM6rfOPAGVhB1Tc5cydnER2veBBEjdPCGvgFlzWYOvEP6XPHuikXlmW0riWgDqFtkN/stFx61
Mn/YstIbB5hMCXDFJUXRQdIjD4owZBE8AzeAg2ELi+zssPJBOgBJIwU/MTgi77VtFl2X/cU0YWew
g0nRjWTgvQx8UXEulf/jT4tP5cAY91Gsu1Qvc4a3gR9RXI6/gkXIafnSeedutrLHSFOpqD5rwyMz
eSMggwpckfKpTDv+SIB/g/kJPdb9Fzy8LiBzoIAj0HlPTNABD2X5JTQ4to6ogso6wvcZF60XlDL0
jRw7RHRbJkPaZxoyHkir+l2lmQIc5feKDHN2/U7EaaTx1BsYWBuV/wfN11ABkZ4VXE3eLOe+SuvV
thf7qLCU/+kXiC/lgd3mfKAw2o62KNV3pvOfTbVUUM4hVf8xwpmgxxCAjMoidqUQUwehbEsgYaA2
riREDzDTRi6ChrUwWG9gElfnoDlAr5ghKwxn7SQDJmGWEnqP/p9P7BlFfFebUezgMWk1z69lOJSx
bMquIqvP2N0g87zzi1ve5kF1lFbphSHIga8yKPpR2bgeQgVHtqw/KjgvWvcqkkH9zDp2Z1hdcaV6
ppzxz2YyoJp0kPIEuqY4NxI7dasHMNv1KuecZEgLK+qZUAqswoWAm7FXW3mDGl5IXX0LCEHxRsNh
EJ/bw+hTaa82p2u+gz5LxOZckNf8Xs4NIAHqV7mJu6zxV9VUUL+OEAvg8ewsZfxuh9eWqQC2bt0k
MmRYPT//RO4yck4wt56RbJcb0/fdh4AMPlSe8wLcIC66tSakLi2LXkFE0Oigzf1pGtF5jJrHcEmj
7d4v6xCMqM6E3TEuUEzWIaG3VAVA3Tr8PqQuEjd62dCgHgocr9tBP3sYb9rkTWVpSBWQ49L6i6XS
KXhu5ktYZQ8YIfAv8dwD9EtGYlmkZpOUOPqlq2l5mGSr4PpJsylpYTar1Gbf4sRh5j2ontDzXXt8
tcwWzvEQrW5ngJ5qW9gMO40RzdZoEtgqLtl7/kFsRLrGMpYCetTslTNadgva4aAG2+EBjdO8joPb
AE9X/ptnLzh9fc6Ml5F+yJctHYi9GuN5BH99lPYnEYsguoh9cYoFHd3V88RiX7AVdvNaUlDAyeP/
7BA7FY0Gx5GpINsFY1eFszh//q/LOmwFVh3DZoayYFk7lZdSACfsvD0vRypI2tlc6l79pUratDp4
g1iFPLNQhaRaoLUmMFfhUOHrLvRmU9ZIq6OdwKaaAfG1Zae7TGOD4eZ4O4hjTz3S/I1KhVqvxv48
2BBg5WJG2Ccv6LZlA6t1YdQx0K+nn4EFgSFD6aBohiI/m6EEIocSvLt+fpUMogTV5BIjdt3Mvw4a
wrO8ZFxDSDuz2LioJ3V3htpDTOzLK/nO/j5AfbSwwWPPhj7nfTdCYAxHmuiqKCeLIJENTtb8WrHD
VW+6PzW5BqQXJSdCQD00hzpeUFt8Q2KZxXdb/kCG8FsLQZsWpyjJLUWmVd0mNrRuZEurNcs3W8V1
qiHUC90zmv3cx/a6Nde07oAZsWFrz52ocTLuxWgnD7XIsOo3QwiUJ+5Gemx5fXwEPZ7Noa+I/fzQ
aInEJGzC7oR9OZHhPIS2ksjLtcdHwWYayY/m1rAangccGmP9bA7/NohbPuertfIoUqCxAMkpgbkV
sNPj6E3ErULj2DWBOlQTU2KArnTMHZZ3eUvWdkETHtnqoASvEkZXe0ZssNf1XCM5QmafBMO/CzoI
ojEfFGXgF+hZvOFvMgIyiRvUk/HhQl6uLjKqCte62UnKdJoRd9i1UNZu0gHA6+En1BKrALmgQJxD
W45t0QAbDTwPu0olD5doxlSrKFndiZEgET+a3glR49oQBd5hDPSThKwOkKO9sPkfxah8QWbmoXEv
TLE7yiro44GN/OCdmcyE4vVGhb2674ktkuT5+tYX7A3iaLZT8fnNAbpvA3M/s4xAi68++EiUCJhp
7ZV70uTdT0NGezWemVSqzBaIruDjY5bIemHKjSkmdz0CJMY0DCC+ayyIXjV93qKv+wjNAdRKam3E
2NUxZ4oxHJi4lNet5C9hY+bzriu+TxVGIJQo74eplhGD/QXWTTNWC2P3OSYszjSmqV419/BtgfDD
DQlEHcLRJoCrIJGkfQnJwTxV+EZsIg0P6MeR3fR4parnweA1A1OFBS9W7f40Cq48oGCeP6mhwf1E
U3+iAQDa3m+u4H3EFGU/lyHS0IfMTfWYxlt1fZl6t4JeDRkFITY695VDvfQr6GXqrPLVMk5kJzxl
kKoKvQyKbzm1FpEvA3pc9N9vCjylUMrLN2Ey4DWsLT3EGrsucSr1KfP4DKUdF/kfMmXAgKJJ2MF4
nwezsbZfdpAEXtUT2GC7ph7uXPV99rkrBfpwSdNf0wPIcUc9VN3F21G/AngvtSss/4dP3MLsc2NJ
cznUCnovK+sMvPaSbP1jVBEF5v1ViEYHMq75aYbWlL7AnqFR4nwa7Fc8WJr+ZdCW1CY/S3UQd7Yx
mLGEqu9a6JMCD4kdn8Fmn7rzNFTNXMwCwBF59JJYKbnHGjIYFJoWE02yT9PXf/s4MrmydqVWEcJx
e4Ia9n1wgqSdkSMsXH9v7vZWdd0kDuNshhTg0KrshIG5+w8UMI3CJdJYkxvylN3hgXF79havv+/m
r4wNwD07tGHmKTi8e/b6O/E5YDScyWpH/4BKeJEq+yu+pGf0zi5XFANHssa5wf1MrHZzmKys+ftI
Fw3C4bnNsh2ci6BldBQnSPYzIOst8gewDhrvGvUwY2nHxNp17O26efsslwEqTNZiucoQCpmu9nnO
+27ypfOZ7pCJKvWhvCwqIkJY67UhxmwUB7Ug7Mre0khEqW7uRGt4PYfVRMp1fg6Wzay8ncHCcRyR
x8HU2JTjutbTV3G7+AT7P9v0T+RuZnscCguDpFm9sC2GOn0REEkc8AX1RBjS/tGclRFNos5XR72a
ZL5a+5hzXbepJvFTLQ3Fvpg+3Nv+IXo6I7U2VLtyKJip6YsZ+b3G/rx6CbPOqHwaiRlcs76UNnvO
sXVPwI3KjzpG/E8C78WdqtpHQ5OtJ7Tc/IBeG18PXmBd/offo8MSMyqBoI0uJ65Yc7bjEOtI6ID0
/6xbYkN8LJSkQX81yIjzb8DnYKVGQI2uULoQuMUIt12ob7tIoK/LjYvgjom8gDhA4eTlzp0fT3vF
RpjIB5mbGiikJt+SS7JcwFzNm/jpjvt1+eTutIkIp/ZarrZtTCjQ9lb+PaLxzwtx5pLALWEn7jK2
Z000rElSODY4U+nbslaYqDQTwWV/8yY6NWWPu4+3sfLBLxUr9CvL3LyCb2Pe66S56b+5G8K0Ah4i
lLwG5NmsErHLMYRub/h0rWR1gbcsw7poUCE82nfpH1xA///GOwXzW4QfKtybjXTn5SQPCtJmrOhM
4JuiJKEiDF5zpoNf5Er+eR9q5XOxLGWlpniHvA0uhK3Lf1idwAPT3jq07eCn/4WbjF2inRSEE207
IPocZrkwXQhWn0DVHb8ZusN3Y9LkZgvIHAoqUjkcZS6TT9Vren8fzArb43GK9O7bnmmKAhizD16E
ngGvhEGr3WU/4n0i85cNd1xhfpnvyu/zl0bn3yyTe51aKvdfsKmZ2Qk1KmEcdAbkSxt7wc/F3/iE
t+Vpv3bzDHnzUJ2Tnxo26fXz5LSENDVG92jYx3EIuMvmjZ9/ubX9bJ7UIG9b3wYAxGRptWNDd/yL
u339d57+jz5OGcTq6X7h9/b8D0ZSJvQ6kUqFDV8kxz0bidya5g2HfvyarOyoJsJnUpvGFtDG2L8f
H+phY6gnP7mtdoren/UzXPK1Ttbdn2FNTftPysYxpJ5V2QxvBOpAN3MNca1Pwyp904CRs2OKbdgi
EXMNoNgVJ75N0MDRSDedOwvk3Rxrre0NxKu4LYnEHKwoYyRDd8k3lCnOwrXP0mhyM9vYORqYOniT
+5PSQs3wnKejIuVBVxM3ll0yJ9rvmGtFraI/JZ0QzY/OlJyzB/PFydJvDghmw5TOTrx3WjNb9PZ+
MW8/bwjb4CcsFnp0A4LNwC5lmv+j2dcLL3GYRb89nJljrt/bDdI8hPVi/6WzzSCgG4DKsDCDrJZe
X+uN/umRmFwFRr7TL3hl/48rqbM5E21SpdQ6w+cSPVR1HoF4oceC/P/DqpzROGt6wn2OV/3zDOig
zOaHar0HWh1I9FsRSnL8+iNF3h+AYLY7LPmrJcZjpF2Je6pcI4h1qtMr8vUM4X5vS2s9kisgCS0+
Qip/KZvpJxUFjrWmwCcUk771IDlCePTkjzvG9MKEzDvhOhPvONNITA2yeJOwDz8LqdBjHrR8vj6s
Yz13fheCYOT38NWL2Plp1V62EL2P6WxBswTev13q1vsRMF8yoqInQNWxxOB9f3JDWEju5Qp4TioF
zGsYylniDZf5oDRSGQGTfdSbJheWq6+YVQbGbzPX8Y06xovStDgvXV8Zh8bqLOLvq8zPV9EWCYhH
R1bQkbqxj+2AjoZmtsANMKjuBN3iFwErK0Pvjdg/ghY7H8kuTO5lRJd0niGBtxEDxRaXoHlsdzV8
s5C6sia0AqQJ1bTkjRjAuSXoUPIgChe8mtZb8HGpq4RRQxokngycJjLBFpIh9TIcJxX4soG6dtPe
9+cE3c9jlpNUAOVbDqS1ph84CUcUyBJd5XjUYV4UR+p0hKNaKLuANDSemjugcgHvODCK/91Z8eR5
O/ycyCxRdE0zQ41zojJkvRO+UPpIKlSkwIzmyi8drgy5Rx+rNdsHJCl1Snude5OMNhpgNPmF931c
Iardx/y2MpzqcXM3G1wK6xtLdLb4LgRip0egeIHLMOsd3ytuIj2Nx9FtWb7HYpgm7cXAXkAoc1X+
n5zj6V/Iq6NxzNBGRYtjGeQU9cZXfTMc7KCmcZRaD3rCgC2atY6TYa2HrNOEI5gSDxIppoiPJKVg
sUjHuoyXl5zuSpfFmTnpenLrVd45eNykd0tIbPPVhh8wnM6PEuWd9IZ2kt5nRVaZIV3sYTv4E7U7
TeOZBe2dz5vBlaRA7Xoqk2pw9SNRVGKllT8xz/IQJjdch3pkDknteNUpkI4/8RlY8y3wmJ3EKLQM
C31xK627nYo2JM96qdGQRYEBPTp1btpjXR/mWS01NtbjmdkmmFNUy+AkvQcbS88inyFHuix6NXqj
nPIsKiTTcL1IDAnv9I3AWs/YGOu/pbrJyi/Y5ka9dldUc87xxe0F7T+0hmqf0ypZVLsRGNw/HTz0
F8KY9TRoIuQ6Ed0BOZT1IN8nfO9xu6k1y3nJtxYBrsmn6KDTacQVo03ErY4Ts1+6WrnHM9XHCM9o
S/YGke5lOGuhsD8RfwjudYsYp3JP1eNZnGu5YEe++jGezDS1eHfE8AObj05wTVY/C9zufJaGnhbn
Gl276TYcjACU+oBKJ2/Uky9ye82K+lufSqeQ2lzWMyOd15tw9jhmzl1I3we/eBIShAgtJixrgqD8
x/HXJ+nilR7pM2B9QsyhoPGEWHX/RGKTiCwNDjzhpbfaHVHe/h3Y9Q+H0zwWVHq0SEYuYuQMToM8
YmimLe/p4bEav8evuEaqefZ8qbbpBbD63KJfZ54RrneawEFYHmUjXPVDrKxCuD6UJZ4DsjmOq8Rd
8iDhaRrkR4tkB7iO9blCxF/jBGwPJHa7Gm9aac8y2Zyfqt7KA57QvS6lCZRi4pTMRYwvvICTQxc7
6gvXoDSuJUCE8bCH9Y/AWRLw1rRHDNb+BEjUGMYAbmEOquJVUp5kRWEYS56ZE9AwPvfjPgaahtyU
Z62xqHSxpYhoFG1g29MEY5BnVo5AXSzVkRTUh+V+u1VgJbp5F00Nnuyr3ajJi/4CUFtBu/BHa/Yk
+CmI5WoTNSf6p4TI31E+Kq61+a1aPSyJwrpKqmUxRGcbqx3uKwCMqhDsmsEsjLI77B6wqX3nBvp/
tnTz8E61aMCWohurLcOtBMXH3nXZkqGCL9CR8uQGPSbT7YdQtCHkWkWln6Y+phewcJFrV9XfaE08
slLbU+048FoFNv4hOOLsR6rDY9wLLzttOljkXJHYBUR61BXef8svstpPfqEUMczxp79261HShP0n
5UgzkoqObbjW0y445MmRUIQH4d9pijOsJmEXcbYqUygNxm2Oqv+qDNoNcNf/1an2qoqA2lWiwhJy
OrjNfjgt/St4ACjorLYDMFsm6GJHUys7tojzpz+AX+RZx79ARw4S0lWIC4fqT+BUM/LyBXdZmc7b
VKIGn3B4yjA3KXVYd3h/qVKFKn/F8AxLpmZki+A+Aqy7/6gMnL/gD+C0OdbefTwZpqp7P4VrsbKK
AwYq8bZNdfR15a9PEgFp4U5R6x5UmPiDmTTVCaS4kryNr9IPV5vXElXCvGHUG23E1xYDf0CPKoSe
QxwvVUQYVZHLmTubQGAfaZAXCRKncXjV/Vqfj0IDGYLgRPrrQWeTb+1X7k/5132MAb+bR9rdIysX
G86UWCcpWjQc/MWBCsfi+23Dte/LPSf1wHrPF2iEoDqMf/qFeahmYCv+aDgh5BOmrvd+T01UY5T1
K9DqqvtEykDtbjSmeENtKuJnCqHkPzFj0+QnMi7b9BVXOyvDjHi1g3b1TJV5bcH2OS+6wumZ2KtR
5pXh1EO95ge1cBb9LcLBBGoV8GU1YEtxqDZUiIX2ilPFdW5ju9x+dpwPXmaEqv+YoWbRJpz7W3tm
TGbdJFfMulwyyyqA7A7z7AY5P/M/PmA3gyKlsnD9b9n0iRzejwV+2sAKetHjIFwOFpI2Ly08kbOk
YatJ/x29hhZ6JcoMF9cRZ3/g9Gehsrv+S78KpTnKxWc1sFogE2IgNOGHmSDBBmNyLNqsLgQKneds
WmpGZHUZYdEkpDebYg2DjAnhqUE7t+4JIdFA1LoreiTelMugicol+zHnYP5yq4f/MYiOgJtEzLLg
g4fpy7wrJeD9VpGZ/G0XFVSHuhVD/o2ntgvOBHXaAz1uBOsAunsqYyALrZnIpCajwobVNtz1YP6q
eMtm9ij4V9l2f+Wr72g7sc4pohlQQiPcmumg36rRLthVx9IPf68Q6h5Cq9Sklo7xDvRMXo14M+g4
x9F1KxJ68wMwtg1f/hvswp6kIJPsEqvU81a3FPTJIlyYX0TM73TDsH4Ej4Q+1ZnJX4yFvae+aB5G
mO+p/QKI588mppS4UdmFETF0VSyw6mYWK9M1R+AnCfT3bn7VwgLTaHofGTwYtGLxGpylS2KTGIer
5FME038paybQb8cbvCNn5/CNsy5sp7wXdn7KYaV7NaX7lFL9dsxX1GUEfOQzCQBfQKR5Zjzv0XDW
6xpBY4XgAZcs+ToHVpy1Ag2V3QUfoAkwZgQmshs+b0NX3c9YllglhsLZO/31wkEhg2n7jdgAC3Qp
D7TF1R8F9O90CJGtapMeVuVSTYbMo3ILM/Nh21/f2j/v9TW7IJzoZz6TBNtXvdvRFm7gp0MYoMdw
XSMYOLyBzBlTPaQSsahvqt9AM8k1eAaPDRIvhzIv4e/nAKObJO7hWpCjN//d7wTT9RhbYgJZxLpe
zmQUHCM2ujY+J4ROVg1xrX2XAkNKaBcZ/3Hv7SLdITZRdmHeUzLPAc0TRIa6wphNjQ3lMozQqxGM
gYiMKZpbL4PjVJZVWhctZ3OzbzW43Bo9MVzHrMIx4A1U6p8XXmgbBrRksK3gJpqHIGmxSPEgJHpP
FERuNlYddrDB5TVAeDKfTyPxwGD+2VJzEpBbrCLebvumWCRWQiHn41LorASlll2U9LsyiG5q1lRT
N/aNQyTC27M6i94QANYks+z8Ei/Kiq8jAwtgLYLyU4MCXmQSPERGwbbNB/Odgw2lA5Mrj20ycN8U
rLtMTyctn7YMT09jrNaNP1A4/dyMq+iK41+X8iLZdfHcT8n7kxnU+eMyV8NH4FtO4PITZXE0MB+N
bnU87UeIqKRVgY85OE/a+BLS3mUOVrHZo+MTnvfUI6UXNH0HghvuEbHMtfkddOHo3EazLvyo+/H0
1CgdsVmuc09LWpPoZZX1c6jatvZKdb5VCg7ILUi1IlWwrCDrMKlWaOjIeeQSfLO4jrQNRs2RG+Zj
KgZVRkUMpqMWUIDVgr+Ze79BAQogogspM0UDtkILAM2Ef2sS8JdjX5mxLCO8+Cy9Ghj/hGDEeX83
MNGZKHkaogKHCs+paIlmmOaMTxZ0YKnGJYHzwMS5uulWbww+gykeZ9RgUiG8aLOT8NzeNqtdjFe1
RrotDAVB6TmoGDjnsOBdm6Ya22FuGBq4EODnNjt+GBJbQdMp+8IPhJZnDkG80vduh87mv/AvEpI7
4OgUnNYt1azoPqLYIbawZmjytUIuq2Cl/C1Ugxf5rJbaCjX3GPeojTHDcCpv6kXPqP+qJ9Py31uH
/qBpUz04Pb1N6ApzzU3keRwUGVh+H7GDR7hehVhrQkUuhjPxswAbhvjDjQeM9yx44TPVL4MnD9ch
wO3EWifjZZI7/Gy0KIfBs/Xa3MMVmuKhD0fVk4nIpdeys/9UvIsjxCiUTD3LbdDaUXZq5Hsm++0/
dUiZ6VEZ7ZwJExgD2361BFYHSEOOD1PBzroMo+1U71GVdqBgD7jBNtOWr1gj2XAu2+VQf2EdIyAZ
xUL4FKyJqeuKvd1npwU+W3kZNt9DFaEEhYAeMC94Ghw6XCcgPCKxNQstW+tCVJpqAi3qjgJ+AiSJ
F/iF/0sV9bmtn1E4jHAUryJOs+eYfKUTTsA4rf9vdtmFGi1k7bPMh03C7NbE2OgUZVN4/NYDWYxy
qgAbk1jQ9xuBGVCXHGQoSkEcAwO0+sfwqDEJQ+vyeuVvWomRcMIWxqMCDQCv3E+Jne1KdO8qpVoa
Z4QQadjVI4TTshWAAx7Ef2tyb9kdOZ06Yoe8+ti0rbhkPPvjCDwiXUjpI/ivU+7uCPT7b62xcsGW
237UiSMjRNBRpiBp8TZIc5DinYGXgBQ7/cm+L+W99HufyktvId4fDKIV89zgzggT7dgLq9HJxpDT
sIUlcpYJ2JzgyL15pdgqZeQulxNecQpNq9hbEvti1MSB01qKdlqHMBhiSFzgXBKYWyNy74tQtYJA
/BCCKfuBVOUcYhYrrQKoyS5XJYbYAdLeWoym9OOv74uqaCm+f5QDLemGLB3yUmYy1d1VqcRez6ED
a/BlkH/qoUPmpg9+pVDTPRY3SNuIbR5I7s70jeHO2g4vb5VKsXZY311ga+fnR31tm6pVGOFNDkSj
xx7eB75BCsegvtSamPyx5zhFo5OycTFe9u0+N1AHVhMlXj80m2LfwKVVMCalC8d8vC44iZPouNvY
GVyictU0MWM/Uuh8nBgKU1J/hftyYTgKSboR5DPvOZevYeExda8bdIgs2aibkWn6vOE0MyGGWZgv
xl/TFOnvtjJkItxdDygwMoCku3jdiuYbzjtEjMRuNVWag/nM2ri2eWIHOWF9jcEoOQFvkE4jmyyl
5/KQutvFMqsazCnalq9Lov+XgKy90BPRHrUY0OtMCtx7/xbsjLO9KyhCyvjPxojV6Nco9htMnh7C
o57FLhFHzEm5IopL7+jvnA/H3lEfzt7Bz+tiypXR0lXxHW8UTn1TlL7m6dVC7GAUSGP3v9H++UhZ
0fEvaxNuGVsLK4oALXyyu7oUGtgKZRZQ7+g0yLh63KrasztILl/WHSle7hjoa1tdaUBEISCHsWto
dEVaOR9gNJAW8WuAYhAwJJHHvyeha7w17Bc88ZFf5muO+zjffCjIkjUVf2PAAmvi0tLF1bqtJfgA
er5sdbM5EBSZkW0QXd2ijrwQXgfYe7WRTT1CZXceI7bvYLQ8eD2d595HNgRtb9afc7LRbL6G5w+g
3WmwjjUCxZg59g+u3jqUHVQivcUM4vRErZNWykTVrTrY7MaUx3jTCu1EKSx4QkBhYs8fGlI8+Lt7
p5q5ffeCV+SOCkxtQrl7+r3iuRPeOK8xo+V32p68/64P7p0TzlQsX2Ejgr6tvWGJjzbZNr4LjiCK
/cXCpJdZ/XI51aEuEmGZ2z186ODc1VX4/qdyyxlc+E9PWJDBnEl8dWuocGIfv//SZXTSqp7PDBXU
lYRaeU0HFZBIDNSwhzZOb+gR0esLYY9N8lPKUGltPlP92P2eYsDpmyFdGFfF+6G23f69IjxEwLCF
/io63Ens/0ctleD/cbOmH6vbxjEiNZtPIJ9sES1WZCYkqsSDUIDWFQ/7kYtcz3hHIewvAnjRIw/Y
1KTpT7rDXoF2SJ8S4pRycj7vRcjme2veQPZNKO9j3QQOFcxWNHb9XweSC1i29dVwFYZrxCnPL15r
Vk4xE5L90rXO3G14qe5/dGXzgfme2ROwUG97pr+L1cEiBIPNCFsStI0qCXDTZzKo8M4/29eYtekI
hyAPgiAnc0znwSGCljT4qnwf4vNkRQwACyJDMuix3srv4D7o8rAcbWvT8X5UZuVAuF4GaNCTbulE
poMRAuqe+m3pagKdQw48dzN9Gxteb5+0y4xZlLG/Xp+IYRGM/PO7QL1HZSmjK18BSAOIid8/EWyD
DJXSvXp9Tf4U3cWI4ZDFYjbAOueasGXwRE+EvsPsFfxiLnfx5G68pvLBFo0Wr/eKjkYWkxOig/oN
86wUbbHXI8f8u3pnHDT55GpfGVXlt/Ts9lcwGVOY0YxDhEPe2A4WjjI+qwf+Bmt9gdV0N7z8tvUv
rgtqevUT+7Y6oRD8WRI0RRMoeu/aQl//lkQ7fKAfaLCB/QcPTT37IQXoSJshZwodQl5Y6r8VR+Xo
ftEbdwEI7CLFjYBDp3KCwbF0d2fP/gqHCry8RVMLTqjsGrPtBEEZOxbK+OO7Y/BwyKFMGo7DQQfr
ExbUt/84hswbzIz9nlonthYoBAQyYlk+PF0AcATRgkAhQPLogZg49CNeX6qB04g+TOGgatN+4Pw3
npyggQ1A8BUGiDI3Ddk7TxOe6Ada56n/ttE0eARS78VlhUbjESaI+QGc+B+Fl0N6Lfbh7h4D4kxK
kLzAflhVq6OUZD3px9btxFncIJle/Yhq4afJ5i6EEmD1PCXJmvw4NdGKIjGQr25S5oE+CuefWyul
fSmoaV7Z3efId51s1rLFGN/+fmVZmWOkMf21Oppbu1ep9AX5JY1aurWZyW9aXaNy2O9jk8nNJdS/
vSrlMCn3NWrO5HtVuAvsUCB2xN8EGiNN7V1aF0aswilg2Ey3ckG2CWhNK9r6xg/Vg6/ECEeQxzP6
3jNWroREQ0cSVpEoDaFXzA4S2ctlsFUOVfnU+5Ytp7ArVb+YHnkN8r+x36dK6MKcJUFr/fbos/5F
1Wn2wi7UCg3XQOXfaIW0YFSGXHKmPepDt2GzDpZ4Fd7L9fEjICm/HQzswpI64Z5F8BGe85q3ovJ7
X68T1RgyywYahJT6mvrV5NCu8XvuyIBgL5sRubTdbf0HrpaLgjHy+Cq2MXVsraF3GUL+N3VKEhfv
KGgqLS+kYehy8R9cnAo/vnS2C9EaSUlPmlDe9H5u2hPuhtppT9gY+MUlKrkUswfAlojR24+2Mutd
piGOqRSma4LKrCtGA0AzhPFS7sy+KsXGZ8muCtiaJiK++uA+H9hUAhqchHb1C3xps+Urx6vxOiwz
TGtNf4AJp4CpkHFJHOLMclsb50zdFuCieQSsk374LbRYKX3Yb8/yVxUvjLgl1/5k7/NIH4fwnOkR
UnKlAejawlKAXBf8C/vzqVi4IeZUeCGotej8iACWybrEefkppinYa8wrQIWocMmOuTOL5phTpS8z
6yMFyXCg/t+wRsQ4XKsw1lGLrfA1+HwlEyNRUQKaRJNX+xq8ivazo7P6OijGWUcxbjdreZsYCh3c
C+4AvRWnwOy2dQudrknyN6HWRANCtaqFbFsoEauMwZwZWewMyrCA4aEk2dr0yIL/yp53B4gtRh5t
H1dcx2TgEmqNPQNz6iYjfVpXjwgbus8ycyPfnnBkaifcqGdsdspt4ly2JFqHS8IlQjLfLmNYHbPC
bPqK/BiH/LDBzIcWWhDI6Ick1aE1FkTaAD+Bhr8SVRZmNGzK2Pe0pGxEvtwvNQNBfr6eAOAnSo7q
bg0pz7hFQ+wLmJcyTSEq91Yk2WdfNxzD9inHjeiLVPJVxqTz0BkaJKM1tfNwgRGLmNFP+PC3//1T
+I1o1JMvRjPu6I9DDIfl/DRe8WV7NlgzT9hV57dD74dgZzutmKrNVe0PvvjSqifghU1mCXhOCRkJ
2s/5jat7abKnuGQ6WQs/Zm0YHeZ8WfXbPHVbWzxA0b0ZXVJsdDagD/STBNaNkel8QsLZS84UBItI
St+EXJcyY77d3Koqx5+CjNDnfnBgIAt+T6FIioSN54Ax7GPqIk1eArXZCrvY3jwtg2+Aym/nMNiV
UYBPSUQjTO33kYQY/W8Qu22pfcVEtNx+d+PCUGiadFhAUJW32tpqU4MG6afZ8F3t6LE7dMP58wXL
rwj8WddPhjZ0FzSvm7o8SF6McksusTNlfZJVgr8CHuLNXd1U4hpLLp1bSCJwFkc6EXusTpUr+0X1
xUSRVsx4LJb7nFxZmnlqE1hrMdYyNPc1+/76uQXxd+9qLEcAjYKY4Ab5upmVydbzLE/+PZEoQEJP
yTUor9dT6hhqpHqAK429C4IB+Jv8Noi7EqA5fRnZtaSzV446xLd9rkhDXowcQ071ec8/XsYPlA0R
t+nnTpIHpDEzPyo9uk9j0VXefWVfSkB8nFcx/WTKezWJdIB/lHIJPmPE2dY9+7hWsuG1m7dSN8m1
4jBi9reRrBIcBDrDoHFP4IKhlQKUkBQ4xdwAF6tYmD39EGpQ2s6CTiJHgokgmzh40xrfmJXHg/9b
n28PqUZkf6YVD0pJlRSIEAkqhJ+U4OybfyNe6RLR6JTmzVDxW4tYhy80pTQr1WiP6C0PpOh8sKG6
QeGYLQ2T2Vyg3FpJioKCDBKfvevLyQs3xUZkm4VUVR0tbtgmdcJmSq52Xt0tZrLxep7YaKo3Escb
5ZAvAQJa8h1HPKpJFDIhl/wu/VwXLIiNJqGvjpYYAT946QMyiB/j03qqWQfR6Y7eV7x4boNk9Fk9
0JtFn65Dlaq2S3CEOLeB3xC2mwXRvQEpSuecm9M4HaXegchjDu4QXMdJ4LRUXn1VetvnvJFtdRF0
V8a4zkUaY51+m53I9olb6mMiD0LlpgabiHDc/4eAf/58nBiE56oueNtwAvAoJbkLXbgncnIDUcaB
PvVjPPpZNJBeY5uFYDY3GA3CxH9fa8Bn0rzqINQCEhJrYdxYGyaFwnsuqjDkojDMYOcCBGI7QhsE
mFw2AHVWSXQOvu114/OFhwm7s6qBYhTHB1Yy+6rk9ZJFLnRWYj5I/qJ87adGN6taCiRWY5eYesix
adqQnjUvOwC4xqAP7XnuWHg4Vjfbqf+0e8Uq8lbj8iyUHJbipfmYGgAGqq1V8c4BsH2qo8rwBfEV
guyg0K7SQ2+W4sFYYWxv2R2gEJtZRLmxpgu4sukEgn0x4a20AyU/G38enxL1io/OT/N4K7yMo0HX
s6i/7X65sA9Hgf4OxTn1bpWu1E+s38IyRE9zI0SythYJe4V9XkjvQ+z1+FMcBCbrVKS+iaqVTEQT
aXJxDssAaxvhtcGtdT9oXbunDcxJ7iEqjpe+YqC4Nii6ldKvT40JTJTOnrFfHk6+5mcKRwzl/w1R
TAbDBeGJUFOXCaLft7DJXgWs0MBcb/0YiCrTj+Hlpby87QcNvnfqWhYu0hhAqf5mIcDDTIeyPEJe
jVbZYP9nS78PvkeRG0mfRD0Zj8VVl9zFtpoy2bjZPLsfQKhV8JJvID+CPnOBTVAvAUNCaHZ7BlSk
LG+O3IebvVA/54s49lniaIjTdRCJwbu9biqCW3SZTUifiRTSTj1GGQiINvuy+tZpCzT/UkKuFO55
+NaStVDMkFCliypy+zOqA6eY3F1mIQI06rjQjqDZazml+e5rVgxEm98u0Y4XEBijL1MtnAOIvYCA
2iY4TPQq+G6xLRmwk7ARVUhl2o1m3z0HePIX/26vjOb1DEVdFSskHYrzLx2bQmOHlD+2MbBzLFxq
3YAVDmpmriFkTDZsQP3lkCAasERas2ykdRYfkTLBKycQHhKacYaSBOT9TEZ4k3/XkwsNFEa+VY09
PZI+cHUeEn3PKznz2VaLM7ra3KLSiCMO2OzvL2ZADqiOxXsDz1+AIQ1cXGk1iiM6eYPPZUT1gbn2
89SKV8MDDH3Kn9kDm5C6oEypWr2IsbKp6B8PpqdH9BYJ0Z6y7iV3mn6/4Nj7jJWn1AeUOGU2jSGL
fkRx9rGSC3pKlC2mWpRmpxd2lmFKv3NNCuYu83h8yLnBy/0/VvQfZay07/SaQvjCWSXhssa0MbgQ
WZiGYL1VDEgejhsJr+VnXx0D2If7j7q9296TQY2XFJICQk9c0EFV8KyL0YFH2N7CNAhANglmvvGo
vnieAE6/QppDM5wYz3QuqEQ9HcYCWDfD9HbxNu9xa7nCjwApDNpVaxzMX2nE1mfzxHVjuksbIodO
0KCpBz/ME153n9k42pdTAmuTa59yqKnIsse7H3P9H7VqLKGNa4q2Bm9XPIpHoXk26JZvAtxjlagz
Xn+lLCqPzeA+2SWzg8Kc2Lh+C7R8j9/C5BDQXVwc9LSvPR0RHrXuMJZtrlkhjgJ7WSS1iDFkw7SL
FWCy0kc5dXAEiA7G1I3YIzGmvTfqBxUNkXEMs9CnIrAZgtjYejUWiUAVZK+hphNhcpw/qWZz+sHL
+jQf4QLTfO/6J+Q48W4IGfKRlv/Tc+s32AM74nc+hLCG0GT0Nz6zVIzkdEHtCSxhkTMP+qfLGZMh
FZrpeeeHLt1mgSib1wtRZMu/z0H3RzdKJiM7JeM7zqPbbYG5SCo4y5Izqft66+Y/OG6Dz4YpgXPn
6sct4Sy9fJG2gJDs/Azg4I350MM8Qx9a0lY5Sm7i+6Q6Rmmu4Bwm2LsNp5PP971EgWhILBI4Q5ZJ
ltPL31qso8IuAklJagBHxwMEkL76sgmc9qZixUAPS+bXV1eMp0Ml+1DFlIiuhahnyheZee2kJZSo
C3/dWybY2J9ix54Y+TYZo2FKkN8b+7rtJarFMyBFWIccUP621LjiFTCS929i/LC9A3J9m0UQkAgd
0DxuCgQA/XAnhHGWYwbUc/9+PgOmGCNSLR3bdCVK5Txgl014W0Fa0A7hMtzixXS1Pib6MQOtvugM
zYBYFjA6x9GJ/ol2CSFbWsD9c4IiM3l43xF5jUjLcvmqDKwm3HkVKLEZDdLCfra4mRmIAzrIICtw
66cF6+xJBnFrby8OmVDzrKglFxoEJAHGnQQB9T+6mfzd8ugomrsLigoQIlnbD7to9Etb+DK0u6JW
3bl/EVgVMPLyPcQqZDuec8xono52Wwkl05Gsx+cDH7PvCr1di7YqPrGKQyLcEP5Rrs7uaXODQZ6b
ICPbHzI8MoCIPG/30SFxH2rzN2IsVpClNQaHH07qw+jUbZmheh7sw7sIDUt6BwF/w/S4x9UQWFf9
sbP1KOK3wwGHyCj8xo03/9YoOrV6kJdLYA+wjNi7G05XCTwM5+/GJf+BEPdxeKpaw2B4opKNI5iB
Sl6/jdseVdv14XEpJaBtKb95VYlhLrM+J7KrITu2SKru+UTUrHEurxNSprz8LI8yxtAK5HlbW5Jz
43xLB8N86ncS+WnyrKn1VEjADUzaIWfW9BeP2srvdbf9J3z+ps1nh8TVq2aYtBubm+4vhADk0i4G
8KMz9/Wp5m7my7mEl8dZt6qEnM9cqXnkhJNuk8J1J5BstPzsefoELe+HZEbcW/yxpx2xCx9HE3w8
0n/SHcDaie2bcaHt6x2NcXKQJJOykYafH3+rQStrr33L+0YFb7Gn1/5unX7AgoXeOsarNqXrjTFE
L5mRBYnxwF9jXeFiBpRWegy0JpO5GO6uYlSai2SO1iq1Fwx8unvdIrox+zCOaduXyPoU7JmWhZWZ
+ixahUoTrJ6yRBNMCBs4vEklHK5j6IPw1gVsMhujBFQuw+qupMvTkzkDvjtT9XkVaYG41DtlHjMH
xiInqGHF2usr1p4NyRhsWYY7OllC67cEIrUphv4YTwn6p721KNoM/4ycG/F+3cxHfDOlIwPUZXAb
h0Yo67RPaiDo6ZwJJTONlJtHdbcjdGW4lEKdDg8XeN0isJbdyiYjFr27ecQplQPjJ24Y5vW8t2Rr
9bC9pNdGGzABwryoihvkl7bsG+7uOzNH0CP0qIV1iwpL0EagKkPNSzW+JcdrxBup7V1GQW7q0CvE
lx+WieC7f45xiQZW+oRlC0ndMPAX2FlJTzTG7/MZ1rQulXcGlZJnN8vONUVwf7U9xFmfoHaDUyHN
7YXtaNWKaWw9DkJWEXX5BgROTCUsXX/N87rxGBwFaiAMFtgEK/esNs7I4ymV1NW83komm41WJ6KY
RokB4T+KZjbAW5CTR2TBhjnuQcteLXlslB0gQcjLUd6gz2t22wgT/VruJR3MWRMtwVZG1MKFZ6m4
3Ynl87ajzRqgkgK9sGap1vz1iYeo2wCQP1mv1eGxvHdF1g7oDUVFbbFrdLD3WShy6fkGeZRakXmj
DzmvLH6WZq6Q0OBV5k854WVWae6I6SOUp9PBYBMmM4Y61oouIrumcNVjCF/7D/34wsLP/ShiqliL
B/DflsccwhyXBkAtFkothB/SUvY0vZkNDVQDo5p7/CVYAGl0P0eBNPkJHGmOAidrOsmIYAhxbzQb
sg39QpvZ1UmEGyHzvutS630XQMaQCNCL+oj//u9QEqvMuFuE2qUXRMrxk6W/BJPLijQR4ooMbQc9
wKb2H/ClDomiqBb36HhUkfudhkBnbRpdZO2Q8gGOO/4YrIcXIe+2OBMFNpq5GdeUsXzlXZwA/oUx
8ElmdW71tVzotPecFFl4RcDYGxO6nay9b32qVHRlCvzN3qO+t3v87FvcFH3Uy8ehgQam0RBTa7PB
nVqIv+AhcT/ves8LT8abpgmRI9Y4Qarz+mqQHTj9cSRbSmf2MgF9iZ5NFiyo+XifXstz08ZhA25o
Mv4BZxY/mNv/3INQWEvfHsTzeIwAtAomr2OtRxa1ceC91+5ixE9sJG5MAbyziVt9c13xcmBMPyR6
GT5B2FyzaaisR/NdxEbR5qgVOp4KSeYRSQWmeGfUPT0FO0Bvh3E5vUtelgbZaVNY+wCGM4BemNEI
6Nb/h91CUJiekg2LmUuVpsOkAIVnKhSaZp8tqMMwiiR7ZS4WxAz0qQjVcJBn7fs60itgi+o49uFC
BPv0iOPVvByvL8f4OyK/bueKsD/eQMyxecV28XLovQG4MDED2CVgJmbwBI2JWMhC6G0LnUUnsW9R
uJL56kmrzgu0AOTdiV+VvzEIxJ0pfgQAUGmE4Bi9QCkEXLgvKEcORN1rdXLbez1klJZUZkIIsT5i
C9IU+Toqtm8Q+6kUOyl5UKD1GKrE0M1j2wl1UJT2UpjFyD937JTLBvbyLHZ1fa1jvePywOQ7EBRR
rNev4Pl3UTSwv5XAIdxPnCh+TeWaXfUajyGXADKl4b8SDB6PID3PY9VhrreM3rDJYXW4hLT8Rt0I
rT28zN4hrkkRlRIYnhOKmlV71mdg7akrEc8FpJuPZXoQE0NRSEZfEK9pbfuw23UqgMFFq3ZfvJ3s
Gy8eeBh1Vaa6JVkYd8BP2qzR5zIaaigzaw0lcvmzODu2Llr+6qjNiloLyBVhFXB3ODtrVKt6PHTQ
+cdM+kY0K1dGkKgZfIjR/vrMcSjGOtmjcsYX5Tmg3SqRIdkczqZbbi03MWKY49Zp0QIpUopaeYdT
kCami1fiNBk1bWlWg9sqo0G89kMs3tFzrEjRwx/BYnUnd8lnpOzThtCjTFezZXwDAaw6QjVX7IFA
b4jE46jyD4OIffgBqpv+9rqn7GHrAsgEiU9KXNm5TlfrNHrSLqVeM8vTOpUOh+SesPxl6xGENsdP
ywu5OchLY4uWfiCg4FHmYaCjPAuNyAlmo74GGRpwcdV6vcKtIBfA/ozXT40WfIddkep9AUMsI+d1
Po7PrTEOUyHbb+KVjCwcBTKO8y4vI9uhuV0g9smjVeAxcpJ/DpXizOyaeRsAXaIssi3H2sB43vyn
0MHL1Tdgrg2lKzxRaTsJ921uJmK74tzvCedcRPsGQRIvscPL4SDc2rgORj7O/bNPLwzcJfshupFF
YTFVVugEnCHWFONQDRLuGMJBk68bib3vYUtHXtSrwgNLaIx8KUs01Zy/RwgHSrl5UG5aS+CJ2uyd
g87BkDPGDouO2u/gmJEjNJQ6PxDOJAUi4OzOCWYaT7w65c8Xw6482mMEVYg6SE89tQwIlw6xkdsA
3cVkBkVb33T1RXxb2XGu2f2MxPZuKuyiDC4LMKwM7Cu4MWIVPy7onQxlHK+95ENg27tCw86xagrN
a9Xi8dOSvEsDqmpQrmcvnXj9PAavo7QYQUh2NqaIZC4SHHJMGM76EwH2st7bCvT2EhbfXrEPrikp
8+76RT6f+ML7eca6lkOP3fpsUIMe5Y0PF9fz9JBI3fVglsVRIpY8JxZWpbi91hRqQRj9cx3huaK+
QhTGolst353dazdAQd9btfd+Q+kMbWx6kPL2AZV1wvP8Fa6GFbvuSNH6nwOugdiPxjSMhn/qWf0D
RrcV9bGVQxzKcgLKwQ6XTUESP6xDj8B7oVK1TzUkfsV8kACrkPxSH7ykcn2YvbkqF2f2IrK09gao
gwojbPfrRHL1Nnw+p1ei5oar2FMJmVsveo4RFBDkss5F7yk7Q/Dc6txyGErPIdshPcmzgMBLL4Vc
C98fnWIdr93euCRGu1+EoPoi8lSFYJCo+NQzKcdbAr/2rHjKnCbZVCq5Crz8XPnEd3872gTTHb6o
uNwU6N8aBQyelP5677Sv9VNNjvlpGyTRhyChrVSit1Go2Y3J4ruV98m185FvRsHdBx3SmuonWKsB
npJZOALnaf+MySU64cxwcv4LHGtE//gDN2d6C6RWwm+nPQS26oe+GuG/Wq09iQEV1mIcW+uo14LO
hTprr8sOBMqc3a6iVlNI8L9WSkwr894M9fV9lpwn8rylSbAjKtPlvr1sar/L48jJ2nWEoRuG+pSs
VxkTpKdVKpadg/jiOz+R7Vd9RhF12/ywg6gqXJWubScV+pIQ2w90/kIZBlgPPBWrMdPIScAiQaIe
pe6q91SQJ2AcG5FQNqZIJurHr6EgByFT6mh8Cr53stgXf+WVRu0Rh6FIJnLF4bdlGpMZwiV8OXU9
w5t56OVVgdUwhFx7oyPdYwVpZMXpdJk93gHNRAxqHC+vX7Bk9mWydyzGwUOtp+ug2+lBZjEi2O/1
Mg30xkWumGLIs9OwHfJCIbGQDNhuZmOPBP761LLpClDsr6l9KhllY223njhQfK0SxbnTcmw3Hjbb
ZeL+zNn9PojInIR53GyyVfqoNyPrVtGw1QP+RAoC2eZIagSwirgDQKKTjMiTnrWnfYVIWKyandEv
6qPQTGRCHNlNPuB1nWcBnBok57PE6vqrhpZAff6UYNxXsmjOYZukKOuS+xOyar2OrfhIxwa9HR/I
iyqKqEfsvYf6qNk5XdYu1DGFPzW0xi4navH3FzS0zBDKdk0ykH5qccv8QZFiJVi+uyknRqXCILjJ
AYRBVrfzuYf5/6B/qATxujFYifB4plBg5Yv3lmGxNGIhWY1atOESuxSVZnh4W8K5ESERL0YULrhK
1BRykoYqvHKVOkiQBGYPHglrART/xrbXC/C5CpktXibJA002utuieSe9XN8V/S6piMGfqGQ3OQq3
aurM/ptYhAhS+vaf5twoYiHF9ZYcMOhxYe87AFwRhSezN4FQ9I/zem3kGUCDcC2DhUBIiQXlSyQC
xtoeM4y0uKWSkiGu4zD+E6zMwsEuKtcm1+Lu8d5rGyg9wIcFapxhmmMLGW9Nko1NdbVBACz/kB/k
bDqXK3m6t15meLfUuN6E0uzm2TlbBGmdbP85sxEnDXxbePUEZDsyFmDYxrmnY/rB/bUOLbpc8M1/
Djeztoi8PlbSvcb36xcdvXDP3ON42lVcopboZw+sGGVmHgJhpyaY4uG+mHDnRAVbma/LDyUXGDKY
OFgHMYpNqKKr4Vnu0u1R43WiqZckb5icmkb2elZgNBqA5yyznlNXrqf2nha+nFh8YobWPmclf0Gs
cC7PV+2MmUzT8Yl9DJAlG3ZiGUWGLl8OtPEg18rRMqdjus80cU75eswUWMPVa891eEgaxX9Pl6wo
STt1JMzgvcXm7h/h9L0MAtUn9eqCU1B3k87TCyv9mfi3OHpnqVqy/bVQXS3gT1yKooF+bzTOoMS8
9c1CZopIoirfNjzg+hVc2DUSP5+PMGCPfqaEWYf1mvLQl/q+MpE8f9CUkWBxV1mCU1AU4TPcQtcA
VbbWPMyJotf8GvLNTJXcDi9gdwTw2xwmQSJQVZVVncZqVW9ewjuGjWxzkcUAaCcRnGy+RUx0rfAN
4TQ3OKCNQ8+FMuNwe74XuoCZiMVjHT3XlGAvSjhTgrcI7db0exILz9J2FYow+NE8QmEkoXneG0nC
H+WtQD7uf/5MRGmBa4vXUAi0zNFr/LObvP24ettve2PIdhw8n+0VQGaQNXV7OwsH97SYt9xFhZZg
yfGhDjFX8Std0PlsX7cqiQEyn2aIhAFB84MeQcseRcMMCpz34NWQe4FsN28TZtcZZh7O52qR/e0j
AxO4HJcsBNau039BRmNOOAAZ3tKQ3IGVDcwbEv/jS+Q8CEoNsQW2YvjQ2XzteScqHXwuj+DOjwnN
MQrMX0ZXkOskrZVxj2gZnRpR+k93lSrAs2QkDi1PWDo3UW48tAV06Yp23m8DsOMzHKVY6zBfh0G1
OoAZNZxpTJa9JuKKX1FRTh/PdwjpSNFc6XRES1VdEmyi08sV2lgxwilCga8uO2FPE88TrdMbomES
mn4lkFCN8lpti/+AHvHjgFrCPAicQZrsmgTYHtZI4QXl4ukQ7csZsPHC3ZKFGzlFpVhHfQrh5CWw
N5lPUNep3I0IFzL1VYZFUpA3K21hY0k9bhG5vsqfs5rWczbblR1r3WmM/bOqnFItKBmwm5HRii/u
URK9jbDhnk2/Mz42TXqczzy4w3ehfGaiAojTyOJkEaIifjMPGfg56oTnqUUmN84qWxF35O38BZxm
xN06nzY+sYp7fwTbkrbOdSKtc34f3TDiHZdP9YTPw5zfvyQ1kiYIdwTRKcFI54Nn+1gmoGMbRESr
r0YxjS89qmlaYtGupAdBH0/nMCZT0tx93F2+M3KsHGSt6dGaXwYjVBVJH3RRYVJWEqrUdTPSine6
HsXLCaWa7jdzUBN4//vL0OXpo6DalZAxzaY3N4+bIKyWCdcsbPec4gWZgBsqYkO1TH3cafMJNFS0
9QESRna9oS1YwRQM4OqUP0jTBuQnpEyks2q23oxRRcpLSLOjItKHab2Ks4dwPgzn815TvA1Ot5k4
PtaXh/14XxQrkwhsPArics5Yhk/gKkRRVrby5gz3hiEQ4x89W3h9NOlIct9Q7Aw6WotXM2m4MFvp
xSp6Ku11KQ0p11nIISoWV1DiOMYPPUa5t6+t3Zng7WnbXxeB9oWJF1R0fWRnL4obKWRPaZb3f2GV
HPMLUw1FgJ/L8rX7Va4W8UtERIEV30F4Xi1QU+BLdstZ0lKN5P+zfaQaxvdZOhT5UN4JqTW6GVr3
iW1t15/ccyaeAZhAQ7S0zNxav23b62wUmEx95SKi48vpfTxU3QnRWDdS9Pd2D+/6doWmG7q8gYWW
aprM3SJ9tttqL6xgkOCOSRS74XAEFd4EFRc5rl5kWvLCo7WvP4Ag0e0eTxZtroCiWyb58kU0+y0B
Ksfs5Ig733HmAmzwbJMGD7ZSzUG2nVoRYK95oX/vRPkXtmOxcEWeg9exZ7n+4HAOqA45Mn91j+ev
OjRAsBVwfQFif1RgZm1/6bJPy67BNPhYeXuESXeT1CmKH1lPywnZ0evDw53/aSv/GM7lKvushal0
1RRaCsBtWOWqpWgLmjnZUrlmHIQRGBBv86cZ7qIFNEpftLkFTR+egQ2t3CZ/gwdz1YQtf4fCETwh
ajZXiwjb1SOapYxpi6Q4/tVwKiUqJPUAeEzcwMMjCjMs2GNYb/8zt1vpZhgAwmPDeyPoorrkBPPG
BETvVGuz5koOBDAp029W9MVM93XCpX+ksyFvFxKZXXUwS0QvSGSKd0wt5+/Fy8HAmHFrGK/xaqlc
bROYfw1u3x9NXMFGPGBFsRBGiuoilK4yCRn611n/2/o86Ib6+HMKGngmueyZRjifBN5AYFNare8q
J++vy7XjP3GX1iB4t5gpAMhw3tfmKmufBW0oNljgFkAlPyk99QJyUw3XWsAsZbVpi+MUE86jy31Q
RoKNGSUyic7etJjUEfn8bxs1ta3X6gyFJTG7VFI0vv8oNsPtaDWaJgnxbU3GoxxWHJ3cOoUdzTP3
ld6ISOFx2wubVwRD/3VsSytN2wE7MuTz0Sz44K64KEE+96ibP1GiXKwUEaiK4J6pGl8oRTmYqH2Z
9g2wynS+NYRC3CnOZfJrbduR0wfcOCb2+kxf6BgkbDRKiyJ7f7wbiT2gxdkhHg+cqhC7GlpHXPr8
Wq25KNW7M+g2BeX9oHbDqa6S3I+F0aWm+iXmporh07/w/MEfRQcPZyGXodxnFnTsCgkK02G6AKwL
+Q8PvlvL9trVBIUVqSpb9/i/7KKS4QucBJ10exITJGgmgFWjbh50MTpH14g3O99wOTpO7T7BIZWJ
jNeEbxen9o1TzhAAR+nWhEsEQEKoICgjOnk+90IqgI7qdCB1DTjv3Ud1GL1UK9URlNeMpz9qUqBk
J1VzPiBOERFNvmlY6ZeJ/96WQy98J3NZfwPKJf5jz/YFuoNO1Nbhy6mSmQ4LfEafy7CGJbxsK5Mc
K6hzg0hQeQ0sp1u4UyDsC3GTBezSFMmtnGgoEd3e9BUkQJv55C7MQ5t+n6Vghk+eTQaOx3UEDnKR
4hBmCd5S0kV5QkXTqN7tJ1k+L418v+LaVfJgtp8BFWBCQ9w/ocQ+xEV0LahPymV9u/roKwSQvAZW
oHH10eJy7GFiX+xIEg9I93daTusk4tQI63A7X5rddaGShx53Oot/5/8zV36xMLDO3nlP76XByXmy
UOT5RSqRfb04+/ywkkMHfTMiQ+y6FIR18SQ0+P0ATRXHy+JDhy5/d11oBa161nV956LyekS+iT9d
r5ggcP8yf5boVTsjtcwMLkRF4QW4N5mkjoNBqBFnK8oAz2yLcsR+A+EtYcq9TebMsWfspBjm3sM1
feTmm3Az6LuwTMOxt/KP++hAGOz10R2T8WS2ZypvT52MS42RLEpQCwsgj+O8TEdcMd2rX6XEzCZ+
nRp4PkalihQWNmidAZVigzT0r5w51KedFtreVN0Gg5KTE7E4MsR9T/9aOJtZPv6NaSzfMfrR8UJ0
kl0v3DDvhGbe3E3AxeVrecD7p6SM9qgNVPuv2NsgF4HqfDilz77s9uwZ9TMIKGTHFhntfsA0f7fC
HDw21WsL7J7IBKR2Y3LXwSKxi0NSomFemIhoBXQk7zsoTWaYuciRl8c1lhme/8nw2AKMOG9OX1+v
ZLWUNkn3zmFEaCrPtpZLfL7wB/vuHWsbVo/o/fYEiFG/evm5tckRFFt+4BQ+PfHpg2vxpSpzTPdJ
1quSA/i8KqtySRJz991dV0fG+jpfObd0zvMlgkzpCNTSwpR8l3CzPIWi6gg4etmWiTYPkzoM1jAb
Ozcp0I9PYjQ46ZAGzJHFcRavYH6sde3TdAN9ec62Qud+P0n3uWEXyITUjn7zF9z41g4zbK5swe5y
7iw72a9JopuXUzbKQjCymlJuMMIzmlsmPa6UBp9m7g9Rz5qq/j7BdBkwIbgz1FotQ/DT/kqO0EE7
Ni/WEL8j7EP48vpsRztbzTL+a01pbK0UB3Y6GmjiLl7tina2iK2Bf3XkO7Qz62Zt1Fb67n/W6Ejo
k6Nbn+9I6vEI/5KJhnQ3XBziF0faSyVrqSLJk9JlvrkPWD4/x973XKibOCHnK69AbtVAbgHaBi3f
QHsX5J7Q4nrExA4GIQMLBGGoJTU+Skz2km1/KobmvS7mnpiW7R56s/lFkjzQpcIZ+XSTGwjlup/M
OREU3ewl5fhi/AGJbIIOC5fSQ4t5Tbp7Axa15yaVtAUq051lQgAWnud6ZLT/pkrKw7UcUJkg3AHM
zEVgfHHwYot21WzlXdlGTagAqA1AkTRrEyf7WmiNHCE1GRqz/JtCaDUOq2Zei4p+fdAqHEbJehrA
3tLlUikePZ0clgMqGdjnojip44pcGn7YYDlQPW9H5NNHnDM7vrVV8VvKV3YmujJhArC/BjnNY7zp
OcYiH1AlBWMPEBfWuGmikDD8NTPkU1hX6gyyXA6qT/cvF+EjXVT/Y1UaBjU5PHxoqk+oD06xoCuL
G2KGo5rknUF6pBkYi7v6IvHWAwDB0JbHC9QVyk3t+R/GVBjLJ3uWqApdGbaK2/vlm6+SxcKDpOc9
nLPZUlV0lOQ0P4Vuzkz6QCzXFD20ZTdiW3b97JIJs7TTkL9BTFvhlhaYzumr1r4njHsxCTvd0g/+
9JPsQuDfgHLoYJp2K0k9aQSfuYzxQ1vSjtC5J42yDUt+TX+GoTxfymH7B2qeWZsIoHNnFTombfgg
pz63P2MP8WL+tB2Zy7QXBqV42Cairokk1ijNIq3u28RWGvosiAJrV5pVt4/9Wr/r4Ow1UMUCdDj1
YKAUGJjhLZ1tl/W/kiYDNTyhMuHQ0VtiIgTfkRZe3JfuOjDqxk+f/ysZCbmGG87HQOyKAAKFuQ5U
4KU4rmPxa7JnSEcKB01EVwMUyY91MIVFZ/SpYpjNOllNtAFGTnYLHr58fjytIqq15nmpEVwHVtuw
J0UKnKkRVc+k5vSGGjIzQHYRAraAWaB7bEHXIzN5T0+FP5Pa3+7kYTySSxPKw3sj/27TM6uXC0Cf
5wzMbMTxYh8bKiiNhcaLtGtoVahY+1cW8QXJJlduz+tkVZ2xb2LMFtiXMRxLE7QVR8HhGfA6e/6c
Np8meeNWYr9TEkf8YnozKhQd1KKiXDIxKGQrDvbxxWApYk/7zmWVOA+d3KM1JQLZyas41+XEl9Hp
evcVrDA5hqmSvCL98jdZGN9ZiKyoJrEURboPmgcJizR3aDcpnkFPbcQ99jAbj8oJFlbakzn9xFQp
0mwIbr19OaF4anHPkWiI6ZKesdvpilaWHX6ZYGfQK+fDDx7rUkBrzu7K3KBnortN1rw1tUzhe37L
TLiaxE3OS2pOaPgizUhsV6axbnUrB4XY/nCxvBqkV997qiIxaBpdPSa5Awi05lhax8ofp/8ekjEF
rFcscl7BDC3UbU9mibF5n7e5vKPqnAQt212XTFlcErsAMoSWoj9S83w8yG5y8Q9f/uOKc5aF2Fzg
KopXfoBcLRpaE4EpJveOI/UiN/C0xeFk4KeiP5GoWhr1J+baYzzSIBL/t3xpmovwupCVUh6QV7HA
PS3IFBCJZHvGVA2Uzf4tIQ71FXPtwZNwAFvi1gJ4CwbSc8Crf/YbmNlj8RIAe8fm78DexM9w8jzn
+JKbDDdXRxaQucJG5Pebvd+GQQwS7gaR69z8AaAhMrh4DGcIyvNBanQA6D0yLzz6tmpaxhYra9QK
Cn1py5GfNsjqt0vJsVuTFxVM7c9blAfifPZdNOvngi8rbMBFi0U8y86hsMCdgKsWD5mK5dAvahyp
APS3hfvkUVyhhwk+ejWVgv7PXgMW/c+wI9sUZkzneF4ggYTWz9T3r6Cn8k87qi6nkApLxI74Q3kx
55pyi7e1jxNa6E4O/Ac7nN6cJdxBqgBpawMorE2kVRGPbDdAbzqCVTQNqvkuocAaAkxHOcu1Lopy
O9qHs84aj+3WyRXRk3lnWrBWnr7KSHYMXxMxyvQ8T/72TMA6KFTB0j/mjkMOfQSW4GXJurCBMLgq
KOW2TLCJsz1iFkxqJAQbQTNYxLzP+GG51NvcoPxW2cqcnCsIxx5wr6ScQydPhwjN95fHl7MOpvRt
m6pXRgtN3u38gwlAtHFiqIFu56nyESUye+JPIVX8Dfg4dQj7L/lTS6wlxWjRqwsBsGGxzc3QF2Lf
PqyljLLBPzl9ujdmB+XV4aeT60Ug3sp7ugFYMO/QxdjIRcneNaK0LDI23viECu3ZX9kUqQ/3c/EN
+sJReBy9LNOZK/xr369Q9srKYnlOr2LpVhhiuIZ3zFfXDo83P+RQFL6WEwXNHtnmMYXaF2tETzvw
wSA0zYMuVygB7FwM4wQNvfRoTAQo2gDdKJ4tO3Cj32rxDIMqOFywUbdv3CDp2e5+O4UpQq385ZG/
wrMHkacTCbCi13IJVOQvf0v8z93G6ILt6l0jlbQFvNnxoSwnvVHshSQH2ZYgNejnF2U2jkgfVU08
+pKT5x8f1pXlD+wYiUg2vXQhekFCp48959LIrG82PmTRvqZFJPNb1FDhyGXLA2UqdXZnSaxc8ndm
YB635iuqKersZ6MFMQF/3w+BuYb4175AOg1B/h4EdgZhTu3n7aJlNUTIClPI2RpGyJQS2nOuGS3h
0C+MO/fjpfhTQQiXQCck3XyXRdHrOslP/cRWmMV+iwlhA40bcwBsETkvrcquQJCEhDTZJ/6I6qnb
DHOsMOCPTLXUb8OoI9reQ2Bu66mU3I1TxDcs8kfFkbG7KK/q9H2DHOrzQbKg9g4D080CheU5Xpc4
V86H3wAZYzZwiN2RrHEUzkA7mlkViVZ4RZh7rtw+EuUpbr8WSsUJs4JHTbVIPC0koRCKgYNHHavf
L5uK+KdEe8Aehwiw5SQuqzG3NNMzsJNFLek781tnmcQfE2ex9WQmOnTibWDhQEvlBnfkDHASoeA1
E15l9tUapaSl/c2+AGfIRhRUmCUpB9rTTAMdexgYR8SyziwLCFRFu0dIOu4v8PpNsYL9f3gnLxDx
sRiXg8xPo5Kd/UnH6XmRSxpT8ieF+HmSIXgjLho5OhgfqOYsROWRddhdGRlyUSAM7twi9wy0ouhT
EVMxmFJdxqC9U9UXAhZ2KToxfjYCJoVbNZRexsD6JJH3VqMSVGK35DP1+B3yEWezWW5JU/QbOzGZ
+u37ceU5DX0gfXNQ7ycikhRcIiTe565UC+pvp/Olpo047FI5W/YkkmzMG5Qzwv4A5qO8sJnTIoUo
ESmPQHzAo/HWh6Zpy603B3sllFPYIbB/SpUbUpUS0MIxG1XY9cbl2i9kQnjFmvude6OKV5b0avv1
WZtXAd+pI+gZfL2eTgpsk/vfEy6HiOoKBPnhQ4ODOJ4LuPTNfGLpAl8Z7XDY/1oMrenpTFYJF6PI
79Pg0ta22AwC7RFeUNdtA2uT5PBgLn+2GkBwH+ufhIiFJ84ys7zWet80qBHO2mAzanBB5IxZmrDU
z872zALK1JLqxqEyM6orhj63chqB96yekTBv9XGG6EMoIGbmDv2PMVUpFC1fRV0fCK0vTnXgbFaH
RugU5ok5CENTdcd95jQTuXgb+2xJXJa2iaU1wJmGR6zwcXuun4wt8A6O9pnetEchJnfeihu7k+xB
0xRqexR+4Zro2hhFRBENT5y9HctzFriHRwHM5ngkCl+8w6czQRilgIFijgYyP2Ctj8NIvnePwEpm
iJfhqPiItxRoanjVxD4IIEeujlckXTc+Y1DN2pvPA8s1nhpchvDvAoC48Fu7DMlHnUgUyxFBSJap
pqqeOfi0nIabnVkG7rEV0i6xHVWnRfqISpepFRKXlUSjqWBMlDzAWlPnMqmtqSD4nTnyDxCaQrou
izJVtfbfrKXxUqP29/AWCEiJc+f9lCmoG0bLcItOFbfXg3RR6axiXheQyJRw8MnPJr1ZHiCw8OcB
nghsgMtY8je/IVJNGdw9L7E//zdQN+NWlNjk8cr2pJ0U3jHG5lPdwzE0/BQ2Gl85BSSP5ABsBhkn
vhv8jxjWPCTrTPse7C0tzpqXkAYXeUdPFIEYIDtlfBLCeFAECqgkr4pBcfC1X9Uo1NoDxEYFEif7
ORCCUC8pF8NFBDZeRjj5a76awTaAQ7OCakUQ6YMpgApDWyv9sc8sOctm+wfqq0w2uT4KLN2zPQn0
0JDNNnZNqrboWXBaVf/66u2/iNO8hDYv7YVbCOxfzENy+TiQezPkwAsMqGIomrI36EHzonpiYBud
WBOgjNgXY4lbLxtieskEgVrmFK+3N42iCUV+n/g/YtqMKaO5eOxR4Hgzf5vwt7ivsfDAnBoen08p
dW5ySwJ0DirCHUPrPr/QPcycxdYWAqEvlJa9sxHMY7Ze330DnRYELATGZzL/E6IczrSDYDg1QbJG
nbD6XlhLZ765PgmHp7APi1l9lxo6NjGkjZBb8o1IlfNvonBSGfSpUHMD9EEr0lLpuwegQBgGGs/u
48G5/TMBv+MnSu+hA/dvYfgPIIh3Ot2D+DQnYOF8Sr8s0HKrTQqOQN070yIgVa6AB47pXqlO3Mk8
ynC3TmAMilAFPcCLWESsRMhCPnVwofQgfeKuLIinf1HWUfP5pLcTrsVf7JEj75PLIzPb6/rKdGNb
ALPIshbupIN+2raEhOr2ax98QMeX8GuG593t9AC5xmQkXfhf3ZvPeOCxL17bJPMt3P7v4rt3lXvO
THCn8MtNWOVaJ95eg0dGFKCWUk6bAbB+KU1icQEwk1VVhrstRQ5keEGid12MKddx1X/ojt4GI/pY
J6c1bxrDKkvtX54JY+w/2LSdjVan+jjfXrYuLLVzjw5ENX23jp0W7pwe+tQ4osE4g8YO+t0VKlJX
KnOp4driXfzlB+zNA+THIrwxUntv1nrmrWiVeR8EKBimhhaFPZxJsBARqBoymsfUd+8s6gu/Cgr7
5DVxFsmSAmpaMGPluaSP+R1RNjNa9hnbnCAwdANNSTdxEZmp6NcMTLBAuTe00aa1lf26LRZV1F+5
ZQUGsTubQpUhBUWtsRTh5O1gUcnoOBC/QtL9ATPzDFpRMmj20PMaYb514Dge3/5SnK1j0Eek3XXS
hfAymy/wgd2q2q1a35BFZkJb1AQLTkEYI83yDuVP2GHmefhWALWaZHMEUBgcgWJGBNvF+XhM7mNy
eaYTpaC9oz9OhE8i5pnmnZgtXYwyxnC83aO0uo6+BbxySXri+N9Rj+Qghi+OMxWl6yCAQddr5ZMs
pI+pgXihtC9kn4dfDNXarNYSzn3fuWByJCvyYOsv8VgjVY+kRG4Zyxvys8p1Tpt7NfTu0ILu3ity
EODIWZG06Y1SkNPJEcG+/2TVAfUlh9+FVF9Yzy4iLa1Ngmpope+dpkxsbelJojv5Y5lEUMyl84n3
hOpSDSgieypSoLREziM5jpfb+G5Ndp1vrQzEM9AA+WVQIlgZ11JVnBj+sCveoujuW8+D0HErou/7
7VZCVNYLJS0NTw2I7bcAXkH5qlWeHVxhIh7fwSVdA+aPCDx9rMMNtfvYwHXPOmxycnHYp5H+YE2z
KYwc6g0qIN8VEBsBxIR2+SKOrv6kKSrf1P3uLtI04UscA+Ir9OKqVuvulIFeQgYSm+XPqqG8wPtu
QEsQfOgI+eWoUz9eKw4CwXFIznVab7IOaUY8lST+zJX/bDB4VFlWPN8d0+v5ab6cWIXuteatIMu8
luweP2ZIbKryozZyaPOsRFXOpMNY+lVbHPRUuUnNWdpuBGP/Jpu1qAzgLyS5shG5I9HxNw0DEeoo
LGj8TEhOYaXwo6+JgCO1H0GQkUR1YQQw19xtE9spNS2uWCMQkxe3bRIfRDTC5imYcMaHYy0dBobG
/bmDBZpgRmYJ83/S/iMDeMDq8j6cGwHk1qPu3moXPLtK5DYmIkVvB4vSkwJ31Jkr9a806+wPMbOD
507E6SOLuDi456QO8qZ7m2PRE35Dtb0yH+FsQV9FEl78MdvuTiPGjQDW/gSrsVtv4M+H6wyOS4pR
MlCFDMsS7NLuXhZueOXapOXkn1Xlfk3HpLwL35RPjiiOqgbBZTSml1Ry4DwuC7oxgNzNarUk4Wa1
mPyC3KheDzK9AzyO6cu7gNEN6Ya5BsFNFcwiZkqq3IHdngURAS7TE22nqdu0v05YTyU0cTw3M3OB
yIjacpnOm8az6R7FvnLLarYAXC1aTC5aHowMMWMIbaRpOGhf4+Rq+8b5ACdMAfDERYYBNYlnckO1
47BCmiP8/5a0tN3dG2CuqLyT9xGWCBi6vqhao8sgTV87J3NUM/hREQfSWQ8CRJScFUiVjBlC6XE0
fJUO35gmBeVhnLJG2LMlswfYx3DSASwf26Gy23u45uyxiXat4XBaK6gRy6Giq6jDMN569Wq/Oqw+
EqzR8+Tyw1gtT8Mc2rpb9NWRgdFRYK0mpBlcwfxdvDDP3efxzCS8pNR+jgFHRv5sa4v3bDC1z8I5
FTrgMa/n+qZxBwoZRYsiZMUxiucItP1FO0kjaV4hBN2eWu8PySY/2hm9a0EmNJ9dvEPC2Xo72sYz
XCtVjp21+64MVnRkgRiEDSCYNCuobgObmrm0QjFSjSKvWHlHae8NgbHDS1oW054bJ9fSJulbYE6O
iBh0k8SipyjlJUL3a/h4+Fp32w0GQS1edPjSfkqu397B0Bv33/Ig6sV1I2JhGedQfT7ylrOu6weT
NK455PRYf9KhUk7p7MucaUtdI4/+SMOjpbd3euY8pTmC7ykw/CkWf7aUotQMteMA3SlZjy/Mj4Qm
4gt82c3x7hE3EbQlMEV00S+h+cE2KnJgykDzJKzY0nn0R5EZOdGP1Jyx/A4sfXTLL7/jk/yoSnAI
UmD3yYIaBUttvSichON/TqR3WTz5QyJ+lScH7MkCzXVZJ3hRT1ruAXKp6rZ+wKiBYj2MJApmGlin
WvmURu5Qvo3Qg3njkfzz1OeE44HO4NZkTbhcewnDEToAZhueEAc8y/O6l+M+BD/uLxSPn6898oaT
kvbX8CMbJ7cheTObm4zOygLXhoxYUt/PxxRdgAKLJMi3eLxu7so/LGHKryRt+ZHqXpTHqJmpXES0
fMgTLbgywOPPt4PelLhTaf9lqG2p+BCiOybiPb+zXkHPUIPT19+Ddh+MUzejrzcnusCroQWSHbAO
AJ1+GTzSEYYwes/52gRff8g01kM8qWgtUISVC+L+VPOKErOSZS1oK/zOk9wv8VvJYWcvmOYgN/zW
Z7ctOweJKoiYT/kxdwKeMzA9y6r1fpELyzvlbOzenwbEKS+cGKFAg6cFvkU8kFVEE5WPcZeVXqWk
D+q/BtZqzbOk8f0uH2/zgqGEg3AgzS4/r5s/wfGq1zw1DQW135WOl/E2J/4c5RXJr/dtav1yq8O8
N++9YHD25i3zNj71Gl06JHQTB8SJb6jVc01g4LMO7PS6LzOhJ5LdWU65wWmb297QVcbsb1+Dsy/U
ocDPQ9HF8fKr0nKOvse7xfcEHuWlL1zuwqMYT/eFmLD754MRtcFi8coY4cJc2X7xlLG4BfqNkoj8
dXxEiDyCbFgT5h7q0gOUV/Nia/K+8/5olqr4dTvKQiY43eYawRkp9yhLNExWy8P2/UkmiLmyZKyj
H+pEHlLAlzFmPDd8+bcLtCAX5jiH+euf3Sek1cCL4GWIltzg8lB/TORuLD/jpijSvw8zPUGOy3GH
3TireoNPYwrprOmql/vVPrB9sp+bZKj1m3dzRO3htuJIoQTjINRR9kwfrbfBpAaAC2kBP64L7DlA
ElkWRfdLeoZ4AkH4k/dil1JT08qmjsV5nRZQFHxa5iokUBJS46ZMx2B5FRteic2iXhNnwC/r8ZgG
WdlL9nUuDivQVOPK1YrdoQOic3cb2Ke4qyVw4IKAr77fwqsdg199Nv+5ZoVeBwREAhSBu1/ZRHhz
l2K03QisKD2K8IQwqummB2I4rWUXK4iFf1ZiwG8DUuRFx7XrqjFVnXwDHKA/ZsnB+Ll4bX1a9xt4
SXsKswWZknyI6gh05su+bwEKC8R2YSoklojwd/eD69mIbFjhA8HVnQY3OyEhbTEPg7HZ6aL1ZCwQ
HkFCDyi1B2JEmPKkbJMJpyKncPWRvP1Xe69C2uFP9FG4H0oLJM/aWvlSqrldELLwts6QETZ6uenN
llTswrzDTeGsqwd7OXY0Z/dpCq1elcD1iuBQ9+992JQDRzA9C6AegYY2ktySlNnXhuRxTdp1VNvr
BJabe0ZuV9+W3LSU9sguzLQS7C1zw/jEyHaLc9DY7rnthuFow4r5dFdzmEbK5q3TrrhSx/A42ey3
5SWbNorGa6trvy1OHWqd3Cah+1YCocO5AvijyLAisvVGMBPyIuIfnBLJLHpV03ORcpM8QTiGjC/x
BIXAI7hqDxvbHtcDDsZgNmNo2Aomst5l6XYoJMU6wK1q3zMFCyRfFs9UILNdLrNmIw24eLjoOW+r
LJQ7EYu1wDzWKYc+Tn0sATCIwPY9cDNAYv2FQNOPELN788uW5zLXJQgaXLz8z28A7HtTghxEqu1y
87pqZT+9D/QJEQ1SUmAtaZAhj/ciJ886f/ebgvPCw3SeAaJEYhxglL74EUCGAjLcZvafgOsoH8ZB
6GvvTNAGwDuUzW35PnV1krBz0ebG/FFV1h48oiKN0cqB9v4I86xs4J5ADVcLvTIA6HltfMeKxlta
laP1Gp11EMf2XpjoXPVTSYgfJE34t/zWYCJjTbweANTM82I40agfPhT8FdYc8kZqmf7JiFKdfy5Y
z9TUel2rEXv8gY8uiy4XnR0UzuMVKJ+n9HS2dyMcgsFl/xKNQygjEc84+fTvtISv35mhM7G068j8
XCOOIUlbBKeB39qQ31vXvL/MoNiRudmXFfCLMTurnjXi1k7A37Cpb0TjvDh9aTOd9Fg/KcY6sYST
Qbtd/ofNh7HmU2jY9TpQDyrzsiNYmVtJfOEAbPSefKNlGUzxlfwjQfYBXPvIi3b5IRQcIrGD5zLR
EcOF4mCldxrezxyGRvrduIgZumJ3JR4sDB0X0AWQMT8lnJeMlVz9BoJ8iVCHnVyq2iCSB6/CkuAa
yJIb8ynx3khb264MbIHO46vzthI63mzYxdqpLyKfaWnd1nckJe2/fvOJqv3l8RGzRXA7U4ySjhvV
oYxkQ21jeF/uxV0lHBPdmGvX4jDN5eQvVg9PwK7d6tj+wvgDm9OfGBv83VLSxcbByHfbs+gbnyS0
vHZwufrdsYHdvoJZH6MVnS56Eq2I3lZydBJ92jbt5nUYsp1H5Wy6jMRzCSgwSTdMzE4WO/lhM419
BdXnQcaOJL+oi3oxK4tiCVZk2OCdMY6T2Vf+Mkzkq5guQIDUaN5I/xKJBKsFv57xKxkflpQQsmVn
fAJOzx0KdYVpCItwS8JSg57yfsW5R4T+sSbqI97KEKZrQ6oT/YLR1N5QigQJNfqWsZVcIGOyZSzD
kBbBXENssh1PCNKEF2pW9ieYFImeS8qavfxx69bwFr1ejfV7Is7n9oSgOWGc7+xS9YTKA3KT7N8N
28KI2grYdrR4C3MBqVuaaTfGgyw3JSmmxs/lYPMWTYmcFsKtXId1lhcpB5U8C3D7dDSU/j4iqM87
ItnIHgqKbWf7nrTGvXXhY9j1eAbWC+XOd7+WMvoQZPMWcC+QjFwkpVGvpEmi4MCTTQ0kz1zg3b6w
v7VDli3PEZken3UpZtsMxc5TK8SHd8jDkJdAouYYGRIpY7WumUCBm/+ZcHUEpdSqRefydGoLmDsH
lDpOovzyRw2KodC+ptyC4cW/FkaLq9mRPlVS4mDBG7gktsSZ1YhLiq6ncH/5v07DO8UNCqq2rbvM
x44AKXeoKMAPtX8EKdAb2CdZgj/f40O3+pjn7G1cCm1/tN4zbhfI/XBPBtUKRbNVHXqivbJZnl9w
9QbzGymevqvNd2lvpzHZ3rYIcRSYi+sdzgLZSNYhzXbexCk1TwK1ablpcXDqt45kL7/ezPPc4vGd
OoZVoEvSn81Ys9ic+OpJA83L/NBxi4ZOWvp2z1vhrsN5aJC4mcVES9kYbzcSP2WDdqri1ISZrbut
fsrtAYQMXMl60OhNwQLtjiTzgfNpgqiNDPZxdPdZhpl0SdwAjt3hO7vueOf8GyqGIZuFD0grJzT9
P6slVZo2Wcs7yUippPgb7ZQ6Gx5df/0Txp27IYSv1xriqEsqfnhzcQbldI7WVkB6Eni8cbRhZ3CC
Su84dYitdyKvc+FaNIWE2Wnzv1J1et5/LCW/s8+5R0FiYK/bwqpzj6b7JAbnXp5hbEOqNYECAUbq
x48l2L6M0svp2BhAy4N6xAL5YhA9MfgKMUUY5BODRHTwhejKtMgErSn3ygVRcp28sEnqIuuPcJIN
dVdHLm5Cj8yOk4gN/UDh3gtYUDFStHaEC6Q6yM150ivHBcDZHecm1Iv/9SxrBV0TTAqQ6fyrfRJE
PGQYbNEtJ3O86emfV2L6+Q7CCfjvMUh7sypIujfHlz5eWXwZgEsMwqsU7cSb3ypeMURndwFTgXzd
qfJ/YmnN6b77yLQvf83k5YoZuFT6BxeFoa7vxzC1LFOMniOWMCjpSsFnITtTS64DxW6CtXYxnmRt
daH13qG4Qv11+tR50vR2SeN9JGWLnSGZMdLabpgoe6bEIrE0Vbv8bH4HuI+fGvht4FUOExDtTRSG
Xi+jZI2DVN1jBmhnyjHOqeqcqClluDtbTMntwUY0ah7uNQt6HnkpNjzprHCZLNQLmRJ/oEAzie1t
SSu5SopDQT0xholGqNevrgZfUvF6M4fM5ELYDejtmnZAnsIM5QvC5kyFMxnimBdcuf2RebRkFJl0
ZzB+eq7FuYzY1ftzcD2dZl5K8kJytyF/5RxMedg6xRQWPaCsCbtAQSVb7minHWKxPLiSdbPZhJ1x
igCXHvILzAmiNfUMUBWD3BB48Y96QiK4igXHKhnWJS2274et0T2aih7IxyKgWVU50022zzOOqbog
btbsuRnOFAYpOcn3oI3JeSD78UB4G3p964F2nKuzs/Jj94ov+cmyGMxif06J7Hfcz1YrFrTa9SUe
YXpgBJdjvxJ4JhoPQBKvjpR0Qk9DwTW8BAunhtl5Rqocebe2hsm2Oxa6lWKuyCBVIOOX4wyHHJJ6
BPMSQ4kqFDfqgiXghS9j4jWbIK8NQtZL6GFau4wGRGorWU9MPirezv0TE2Q653qB+vpMEK6monfQ
6UGjGfOFCQh3AUYeV5zGtd7vWCuMnTRfq/p0tYyUleyr19r1/zS9+kChm7XMqbodjIcQ9pob8ueB
0Mr7W8bvarF0frB15jzSNw47RFcFAcId3MR3ONVhA5DqJcdO03j+YurZRPn5jP/5NVOPfV2ZLzht
mykMOtHPztpwm4D9GdH704fDm143yAGqKaaABZDyZQJaFD+Cy7TpC/inqlJYIszSxdIjtR1V/BbJ
Vw5D3WSflO71xwcgaoI7pe0ApIEjDF4f83+1duOleVnCm+/j1cHKAR2TXNrdbkzilSBho7PEDJ/n
1H2wVYVjB47UmrnbRKIpmpaqxhZWHGLoYW2NZKtGStBuj+alfgT452LOECDPlOy30jF1ALiiale6
r0QziyH7FgjaJQ7NGbrQc5CHxufuTPhNeNKQVJwOtg6Vp6Pvg04XDUyVmEaeZhKcY0jnicWfhPsy
iGzmjBPu6okuzE3C41YhbLdV8GlclBVZs4tAd6LlokwUIjSYnMunfiMohoC1iYpdscKm0n5n7Tn2
j6L/8lim4rh05bWP3ZUljmTSEfX6//Gc2D+O1759YosrxizQbpKFUFsivW/eo3o+zTIpRBNyU9lV
DBBPFbgCRsEnTiSF3tEGWfvc2ZxamPgmnFyknHzxDfVkDeFCuaTqWdj2wFAVuDjZe6A8zxnbxw8x
U74olWA2wpJ9WPwGEFu2lJlqjN/LfkBJcZqM/GLmrm3zz9OSAvyoERQ/oPejUDyc1Awybd0MQGwm
Sc8QFcyT7shCUbkvVb1cRt0OD6WpMGqctAWA+79ZppAXSut+JeC3KLd4ug6vneMExiOk0AQ6eycW
ub7HvrysO+fD62vRvS0/nKvEkO6JJZxb1Alo/tBKwCYk6suVW6n1PNVelJtdyIwgpFwd/ry26jen
rIXseyAzrfbjNNXbOzJSv+FlBGcyNJpLmHoPy+17E5CBxnAs6gubsJcSIog+UdcdZGZ1WWY4ux+K
lKKVkPfgiN9mC7jhGnXkDq1O1YXLKbvLIgu4TghZIWL913KbJjGhON2owSI3hBGC38IIT1UIcfbY
ghCTzXNEe9GnjgJaS9criQtcgs196CoSniGX/D8thnDZjCkNOKOZe9O9B0iJSgIs2L6pUZ3mbGyq
Kc07ZutSHnTSrTjXBXtA2pDJzvrGYHRZdon5knsyOPaFujx8VwUt7E2W9iEdnzaaDvmR1vtfn5K0
YFGCskp2Mb+eYJs2U4QeAC3u8BE0NWU7HwWDizfyzaf8m87ytrGrqdtuHO8yRdbj1F5Ab7TBsI7y
czWU+ppQz78rPzADuKuLTFb8BWfaLxkhUL8od7HclRPuDzH1o0M9BvnT/iTRxYJ0A+PB3/dYVc8V
x5dx1r3NG7EsK2/+NnuyDjxabIymf7nc2gnvyPgkpItpm7M8lii0AcaemvV2GkihODmOXwCRE8AN
xC1Aa699kjLWDlgHEi54qH3iXIfHyv6MxPBVVGUDIgAcp2OZwQBFlwZeQVayx99ixNWlk2SD6qAS
neyA4dYLIPY+dPFzrjcHhyrVwxtHmjsJGZq7uTCyTI6lZlISlQt5QKbQ6W2tpvVF1OwuoVXvq5q5
HPTuQjiu4vmaJTzzdD6E7ryRmeFaUYmg5JSZ00MdShl6pm49gEp0+rV94ZY7HwwmM369dl1SNsvq
aB9iSLe7bh8HUU7rm29ei5g/4tzM9Idt3zpgCwNJ24XiqlPHEKSkdNHEHNdPUjaKIY7Ae7opAaBD
Af9JRNzC/uTUVhvEnGlu44z9w8UgCYmlwIzfZmDfF5nA3SuPL+ipbCwHdmjtoRdMw9c3PdJ93A2D
0s0zrpT9gsjjFNzJax1oRFV1tTwmRjDW5bKHnp71m1Dq+OcQnFyIO3N99euvAE4Y1GuWVKjRB5IU
TY3XzjgkADB+pQerH4iKUFSJ0Vri78ts5dYOI4ZF2GDNrgxS1qvD1D2vhxsPaV4+QIzsp5MPUIe4
meVksbyHj054lic+KT1+jtyqtzDpyM8e/qV7Gyc8Z3KVOAuI9dr267VH0icqU+x5+h7Rn94LEsU1
EO+gobQAPi5BNayQ0XYwk+ZYso79f3u/BF/JfvITrqGcO60Khmhfvntuy4TxT105LTHKRxQ0uX5f
8haMKdl4MJ9jFJH05gu5fAYF2sD8KyVVGdsF5kUiAEievIvf+z1u+uybxx842ZYrNlbZ9rcRoQSh
Hlio+KWDZkExJsP7vU2IhTxvj77H7kwsNFigECofQbcNkYaX0vzdDOnE5DG2vqWTwptQfUNLckDq
5z4ZMqIB4LSytF5bZZ+Z0Ha51PBnToMcSUAnS6mb7b1jUnFnDoqvQYo/CrBgUCQpn0mzSpMAVvJ0
ruiylwLuzBID4fwTfD+iP0EYZD54d2RTaEuLYkz57cDPmhZfQyr7xbxOlNltg/C4Cop+BedPvS9r
tCZR8rxo9J/G1LWgI3Gk1wdaI/AY2Ya2cXByDXyMwzWYRgEsKTYtQEClgDUxipzlUwWQ/M39jKag
i8ZmjdsaHhSGjuva95eDoBnRqmZdGuoFtXaKr2h3DuI9YFB8X89MkjLD53Zx2so0rtiINL5zaOZy
CyATB+dHdxUAfEmsaVim1Ikbh3om0R6O1PsHAr+HyZoP9PkQyl40lzBahNUUjjRzHvtxabfbW3UT
QFvF9SmM43x8yTXix2Qh+NlAB+xJN45hiXgvky4pB8TVjzhCnBiiVH9Gt3ltIFoWtn0FzuLS/mvr
dQBiSJHpO/CKyUGP19SzmYi6wzcXaUuB5XHpGU9F0FF4SSqg25qk14YXYg379n00VNd4H1wLdVA4
kDBq6gPrhofeqh8vofCdIQBFOoHxbMPtZYVQCGhGj5XA4fdri7+f84jEO2oj1ch06m0JmQTqu29b
1fN7AcP2dqwkObZtLj0BjEe+nFYSRNvywU/m3HBi6T6Nybl0qfqj5tQPdRrBfxDvU1EgkgdlkDuB
2d3xGHEmagYDkDj4vKmYpgTV8XRYoLQmPQBPfA9f3550gO6ehdm1La1NovwOfX0UMr1ZnUcU9apI
8aa2PUb2V47U3PJZmRXEmlAo2Qun0CxfXAaCS59ccSEkS7dXbUizmQ2UKXKfB6Doc6BW+6HHVo+L
m/XR3U3tq5PKtydwPpeTsM5T2MWtbr4echVSWVilkkM7+F/Wth3eRge+UVALq0E3WKvrP/GHQVfU
zvBqNTMg0rNlKfMf39t/4Xl9e/IEjVJwYk3WBESjbZQ6vuW5a7Wlbx13GmIz/UcjgALwFQPqHoxP
8O+p9g9l3sfiXBYi3oYzXADSKW0PvyQ9B8ic5siTjDUtTeLF8jj3buiGsz/FWtb2BQ3WyoTEbmUX
7JnfXTlOiKopyzywdXBfydJwM3j1leuJQ3f2cw3pIDUYmUgDbtGA5exBjlUzF9PhHsOmsf069NNx
vm+iWHfVdHiulPG20CmKzInoMyMMldz05i00E+4L7NokCjiqUsz7c+n3Lt8xScwqC91/Dv2QNDv/
KH7tXqJyufV3Ez5qtV//DxpYwIWKcwowsVdgbScxfq2cQNrdFsw9v1bSvtxxiLZj+Z9o7Ls3h5G+
aOUNWbyeTkHIw6V4w2GbA6AQg5/FZLG5YDmwOMZsukijY7P3y/wSd/RZfkZRT0z9dTtTN+kAxKkK
KxRd6xlvmrr6hI7I94mJZBw8RTIvhMVYFv+mWrCmKq70h9B2BiywUQRVsBH+z0PP+wqvEV+ReyYs
epgrs5iyyHXJppUDHrqQeQ+ZL3j99e5G8R91Ez7Ifrg6unqXXuy498fraoYfkryvlkAWoML425Dp
s5127o4VR4ELVRHDV4uxYBZvNDSxEct/iRpOg4pVGqdl/XPz34O/buMJoRa8bSSvWPU3mvqdT1dT
pyUMpwO8sQJhzOf+oCjn/EUzNhY7Vemy+kH9zdyt/nl/+bPxF2VZcRvzcO+1E99KKHxeN9Zu3Fts
tXQSJmFd6s+mh2VJpdlpqySqk3wXTDrZTYDVcXhf7hl5XDzGj/wPVaWz6Q+Yy0geG6c9PtIPfs6o
/TE9eOuWtmZ4N3fuZ3O9QWsFe3twaHE9mjDG4+6zOxLMqacH6K/I1xGXcgnENVOCrQxkpNuZUk2O
971abpFGwqSEf3atj7xmlSzJ3nOMeyni96NcJ8g5ziTukg1M7Im1Kw2rSg2+5DBqFb0E5dtHRv0f
dM42iOHzEThLolkjKPNOEkND3b0jJ1kCd2DeqF9+ZwemE8p8+tVX3fAaUfYXZ5Tku9OENsC4Ce6z
0KJNtevJ6ME/1T2AdzX9DwB87h0nuxBuukwUu+u1/+dSQKB6r1XHxFx09lYJ5oJA8G95vy118Xti
d0EkKwzqCko1rvrIC3pY+8dcA4rIyya9PtB0H2VIO/a4JmmB7z0Xh0TIucgPthYBNV+lxuv/32KE
DPQQCFOCy3iwBCqP+Q3dS6iNi7grLgN2YWVgeLsDn9S72PA0JWT10+JYmYXsZ6V4cdvxhUxKp4WX
xbRfKtONrIgKZTsCXVrISnQds3k4CkL1FX0t0v/reN9kXks/9ZecG8epD2rN7NcvWmLI7OuIHBF3
uuui6aHZVdN8mJj8IzODCtZJZ3Y5/+5QC3hMEsbleLgQb6lw0PQ9SvWOxmoXaYcC9XJWkHBKDIWK
EO5+dZ1M7TD6oi54h4MpzEgs6arzu1e3SShGq9NkeDjQJykezSXxv91DTpne1cfe55/Hfn1PQUl6
rRjTCCz7Elzr9UWa27xDe8BsMQOefX8H6SwI/ntOTAbbju4jQhnEDLgJsGf3TsaWAR5lxosnQVfZ
anIxg4W/FY5xTmKowHd1s7U4Opmhrd/b3jw79QKs94OIsKuQ9X0ozbPfpN0D6S6hsQW8oD9AcyFS
zQI0ONWVpUp22nws6RbpN54PaAFzsUdlVpgvy1/BRpNp2IAEAKVueB9eNo7BID9ckmLgUJL42x/z
xukdxCi1pLK65zTs1UqTxlLDg3x70eC8Co7928AmietlMQbl95ZrA+x9yblh0Cw0hs9uNVe/6BRT
WZgTQEcz+DqloXSPQO3UB4fD+sEYM2TtcXh7GC/YxoWawCPcektuqXVe640jAVd0ZwkLvCJk2Z7u
DRq5nOvjGZojlCXdYa5cEphB7uwTDwEgjI6tC7gCWUkuLNhFco88h1qVbn9PTOyBXefvc8q0+Y3U
zZgKPf4vWb1TABf6T0x365nZL/l8u2b+B0UYwVmFUJz+aS51Jslf1a8pOM1iGQ/ZJEPG5zZZTCE7
6apvmZdgs/aQOiIH5NV+THxVbyYysa5wkoIl/MxZo3w8qL+4rloTgQCxiolkGYGGSK9dCpbPvd+Q
QuloNr2vHi5Yl/0dVa0pmZH0HGm9ZJ2qNC3ZcWJZy1cv9Nevcyrphugb3BXygBmnHljN0qRWW6QL
YRSpU9sp0NQ6u5uQA5rEK1vM7JiR9VCROmTqHkwmm1NIIdnq4HAVQiqWgHk/DQV7q0MIvyBtkTpT
VCy+RM9Ao151z9t8RiXu/coRer/rfspIxNxnoluKHuxJvqC4g68lddAwN5vjyPN1HHtwULbZrBuj
Jmmxf4Jerw4qyYWQuILHzO6Civlg8bURlkWmr3n28sq60hUsmcNvq4md7j3h/uDW7ibddiTjhU+T
dRZ5iZf3YxYinAeSAj9bWtQlcd7+05MHFPJNveZhUMHjAm/Zr81iZumbYGOJYS4DJ97FHXy3bcUa
vNb577q8n7swZXHZbxtkmyHDCutaKklkRUpW5Wyuuq6kL10bOozdIhAfzE+6qaZvmFJutOCxzWMx
iP/6clImOhPTIJ18ptFIWXg3o7RoaDO9ItqZY9dXO7aouzlFj8h2Lkej8jPUfsCpMQ70oFaFLfFj
qT/7/wwGeZUE0Ef4mfRXsfI6T3PfyE4XmiIK7IK1lEPo7CADXaWhhxMZCxE8QPR+zN81IqON9Tu7
eeJ3AHt9jPGIRGgC8v9KP7/N1odMu0e/GMKhyYaFA1RE8M6tOjN/oj1O1AC5hJ/6EXP0fD1y2bCi
VAhFlq9Rbt2rEu0GLZ7qJzRFLdu4pB5QUM/UDpcv3N3ZROp0UvI2Dxfumi3qbZOjRDTYc16oCHE7
VQjxlrC71b1PXVVEWM2pO2VBF9xnsqHM27fqzeA0r7x7oyW+A7DD4wCpKRmdEeF9yIiHQr2jikHl
ifiQLSo+Wc6vNrC0P7ZgVZJF3hr/xAoiM0PXvEbytsOlRZ9Iwq+E6NSj6fIHrFgkKNRbsW96wdEK
xYqZV/MaG2GGpIDyeMAe+EPtButL3S/wnLpzMJqKoa3dM4mndYqu275MzSNdlFFaie1nS/eO9fa/
4xpsYNQWKtvIIseFRdHs0XEJ6DwJ6mvuN5IbIQBjLi+fLqA0AuFMANjmyg2bdOcKsJA8rLTSSnz0
GkfC1Y62i3VYSUZBx+1QsOfnm+bXNgubKDjhRK1sZcpaFSHzgCRLEzUz20OuOhLQrV9hs1cPdK2Y
UY8zv1syViehhsuB1MJQKkYtQInN5s33XhAda9IeIUI80sR72NLurXP1AVg5LmXOlSUzPd82xRRa
WcG2pQ6aTC0J4nFuh/FWWzj7rB6fWEhfP2UU9YROwPccICNNR5T2kkyTU9mgUlOW0QR4jgIT2FcX
OwYnrQ5u1g2BO3F5qxtcrxzeZxekCmcnzdXh0T3ewtlExjF4QThmcNiP4hRv3Gvux2tx4Y6RsP7H
HNQuOw+LmvUCCzjxuy1pJfVv/KYO7ZssLDhlk/+IJlX5/diVDr950FFYXK6QYKiL92M5ztjcbeIG
hivHP1e7z8fMmN/oTPc72A4T302xgoF4R/pOI9+3D0O5U47E2Tds9/pDMPI7k8VMSePJBEWhZelm
KxL7TECzYfQA239JCg+B9CR1DrxxUTD9ZM2N9VoxOMWM4/T+I1CtYjOEsA8wQXrH3VffwBycKONr
vB9M9pul5y7/Zd4hCbzWjUDaqGPAumf3N6cPDW57wiuBTveVCZN+pgFeM9cOwUu6Rn8DMT3Iixw0
Swr02YoDIJkLNVekTOMTs35gSDOMKxBTcrsyrH55S+ULlz+RY1MbJ3vUqW/KfBIP5CK/DMqLN3Nt
1DyQBPDhktU4VuniSMe//8k8ffP7l5a9o9GldO/0eGkf2n97LcmTW48OUJS4vJFWuQBowTJyVl+H
f4XSxcSJNK0wLD4p2omYQRvVjr/jzJ4ihZkXu/5FY8k+MJ0ENQd10p2EeIASz+9PE/LTBlEUrJFG
nN3gyk6P0rxqrE1/k+HeDkkyLxVSnXYtD6GlQkFNKaXfZvB2GFHMwgNDB9xL69yekr2er+ZWxxbh
9YHjg+1p1Fkt2R/bcKZuKPNkKyLNR84SlUEweUVO6Yz3AORsdcGWFKwnXxUbDd9OgrW4i6KVXJEH
BvZnO/jfsMWHw5vIlGVniXddiHgvgzrZNzDP7PwnG8Fooz9p0s5cHWcsv5iyRICeGlVOGxFCWXL5
XK236YkRXvtaXB+GUGUnZnbOwigKXV4pnmVdrGfGq7I0so/7oOheN3B6k++2R9LL6JlDZhlk0PbL
Yqdfox7qhRhiMxvZiQniODfEyhGL0tQOn66PMUONehmRNMLLLw+k0sxxUCGzDcUOQO+awH9gYHdK
u376SGu1EW++2OmA2ZFtfJWhGd7Z+2vkAbY4DmvObgoxvdhHV0dvHwVkNAZzOk4978Q8idm6s1T7
fqIIgYM+d8cU2SW4n9PHbfbzHcuBOh35al9NX5WONuS03+XG7zjcLWCqGJcUy9m0+qki3DACxl+9
2QThLB/gNOsBQR2mUTPiv7+rg11kUrtcAl0Y22+3fLuQxqZmTTt5OQVGkKUEVFL9I1rBv6cfAcZZ
VdKCBXepzyMsKhUrliaP8li0uW4Ik6c3GJygGciStvZ1iq7nKBYz1+fesbavfK4cCXVn3X0/DUhN
SaXvTo2VdPBPI8tXCZkLwIWE8CBFaeTLnIx207LY6xiwCSG/cn5YtxZAhcbNvPIzohLTeGw9uce9
gO7YigtiFIA4zMK3EIIpWYyOo7Is50Hi8mvdTYZbPFIuElWw3+qPwb9/n557BSvUrk8/gTEUOaSm
zcXzDrkOjrQESqyoeZ0s9NpCecKBaxa4IzRhHDQD5RJrIManql5MkXFpxxFEgPFfYIKynwtDTJOB
I70QH1lyJrZnSjs2nHUk4FA7GXwKGIZiSaVvI9l4GeNPH8vJsCZ4S+sWg5LdN9tgyOUELCeTcI5Y
rFPxp5+0umSp+2G3uJK2HVLkdV+hD/WjMebkyurdw8tPjQdbQ7zTs3/ys+UOOkawIeiNLdWiMarF
Wj46bpC2SlcFwLVbr3sHbUq2GC2c3RDFeOnIjkgObDErAoJuks+f/jd95lJxeiWh7PxiTvH5FXR5
hChMj0PP0G9sIlc6MP31xqthIkwUV0De7/7SHxSv9kCzTNpHme+oMcHXwXBkrhlKS+Guuq3OS96N
wGFKVF+tASJj1aqIsDLnp2UE9s6bRTipoMeG77/ij+xy+soq8dGccLEq/0QI2POpsW/T/OoBw31o
Y3AtiWyoVvXSyjRX8KcldOpsg0/iWEdRJxocVIme+F9B5kcNAoboM6i9k+aNxPXz3HBsh97kLlfa
qblvZZ1mlMUJCe/d9WXckJZftUrJoB0EZaC+XZgRe2bdlJeH/u6o8Dhihru1Gk0jhFLtXlgiQQoY
7yJRwk3PBWe5upHHWEXs+/g+TtIm5ZbryBhhIbaMvdXiZu1gnSVf8nbz8f7yULTBuKC+kYTt44F3
vO3tvs/JpUc2mOJ2Pgh3EtdEltZvIAgduFNPEDT21cI86kf2MlENNJ0TZtNTqPir0x2KaOmUJVnk
BAgjwk0Kpx4jvhfPaQhiU0P7p4pHEutYcG6LYS3u+0On0WKoSxN1ZnHR/jqU4SZW3GXF/FeC2Hiv
Jbf4duqzFF7iNHtt1Bo1SMbn3b0GbWM6Yi66s8it5J90Ue5jNmnVw0XjvxjksMAbZLcc7AseZcV6
Yp9vv7RY3jSv/G4Mu1x00XYtcTxgbzvQ48E/FIZJ8xTLw/dlGHJ34BnBfLac2mdzuclbpFoWik/8
P71eZhja71dLYJ0OehTZqy16LG88Rl8Nkyy/uEd7WY48oY8rZTIhUfLUaiXb/h3xBQEYe761V3Xc
cxUYnRcbInOgru8Pj+SkV135OLMei2TeOzAGn2M687dTBra/fuof5kATAEwynm/sDoumOanFkRwo
8Wnv8x0OlT9y3s9RY+m5Xyh43TZCjVM18Urny9iV2GUawLT4DV7RCMjdQpZwHAo+G1Ow/uXQC+ne
9XXDYZ64mKewfIy5L1oBD4CkbGv4dddUDmbDFoHYuPDWbJknzknNhJOBBNjZTYry0vh2J/QTcmLT
01DilxLbSXvPhDFwaBIm8zRW2azkkMbWbpT83zFJCMJDj3ztHhopsAeh2Gu1599lnqU6iuJh7KcJ
vsDzExzCgprTxlksDyDQsFYzX0oSFh/quAUXkitCHGnfMRLfeJ+dWToS6hADiWLLU39z/ojjtahQ
tbQSoaJmVpZ736NRZfMSaBSut3xkAlcHzBThJxIE+3+8Zc4ACOHgy1em7upwl7OOGHhdE+RQCtv6
+IeD7enPOcseyTAq5azXphvfqxZjdzkIAVOQvnxFvKVjXeoimWLJ7fRqdGrRuP60QBpVw+MC7jp2
bGJtfz50ZMqaJ1Xkd0bjZbj6ly9w7RVQRVpX4nu2Q/LmZBzT5VOSy7KBccVNEk3RdMCLeJExZTyY
hbD/TrwP96OhL9/AlG57fDZrp3miYlQY6gDBOXCJHNSPBljd4Pv3UAMxwsFalQ70WS5j4MNyoWuN
AtS9G/NCHvgxkxJ52vbsREh9RSWxG/Wx9dpoclYsNwjxruzu5fydo63rtCUCnrp2CaDavyIPo96m
5C3mOBmj3iLJw7zjMM+6tlZ6BpOG0YgS8uTnzAmox7g8oHSLACRYJuD2mO85liOJUKnJNy82rVpn
3vAIMFLnbO+aJO3XYB3/2z/wKc53YUus5aHww7RBmE9cYC1jWsewWZIYc0aeT/ocvLaWKDbLZizw
26Ys1PGOiltfXJ2GvvhBJhNa1bxgX8dolJrmX/qwqYqwYN06l7h0kNJH09yoNeBT1Z0y3yTg6QHa
xLzyjyQA1JGrYRvrhkLf7IGJdzgT6z0T2q6Py4U5Ka56eVwBkfuSqCFRiGt71S6riOomA4gWD97U
DAqtkJryjqprVQYZ01Tq/HweHJa71UDPwuB8GqKmpS45Q7ep8huQghPfy7demk/L+ZpENlcoXzgH
V5zyyJkCqF39hXUhMwPefPSbTBwMZpLoinJqdABFe6pK+WHWc60PamFPIuWTPkC8fNgyth4Ru2lQ
hhfdccHdm5onyjTxrggnq024IlYNWA9jhAJYWDxoHJFmTwzS0c7AgpAbvujIDlggeCwrJB4xpRkf
C9BC2ZMwvUJETh3gif8VfxP6pmEpNMKwEHEnNyVQ/ae4fppjUO/+MfODipQMYd+2j2hqAXcsYan1
tENyesar2uca2rfh+/xeIitZgWpMOFX+tPaUt54jIcL+LuAY9AVTsK6ta+0ZTcmIPMaNCwyIPRF6
6juD+o2jIz9sILlD4Lr4syhRlbrto3rDC98JuHsqb5CjEn5Go1TgOVC49f8PuF/0TrfH+RnDXzFc
NwICEGhqo2FKZLdzLl/qcx3j3WJR5GMk4qdyBOvIYh/Y/Jru3ZzsTtA7Y7XeBhaBbA1hOpnMwELa
tVL3TYsDjCJZjzNKz6oqSOEE+cVchrueC7BlYz8/d3jzDQ0KyN9t+nkiP0hZUOLi5B6DeeECOh8s
YJ7dH98HoAycO4K32v2yUrWzDhtnoJUbFKY6BVpA7aV/W5Ei9AbSfO9ZppGu2m2RlYop+aAe9I5l
fttQJrJguFoXF/PfJmrg82G/JHian+xVHKdjVfDX8qKE3YslUFemFF+ebvJabZFGg+tnrLL/Ej5L
pZ84EnWWkrukAMt6VsRmZ6q4elqWklxscrbJ2JQLlP8v+HubJ3DZQf2Dnw5/Ea4VZeTEJB1XUQLu
OqHrZR6265/VPqkGeIR/HEkzTH63BtZ0fYV8lNwfyMvxJZnYNhknCVncz/75i64sBSww/q9w3Z+o
XzcY9IMbYXUF6s5SHKk0xVdWqik+9StXl9KfgR1OFFd/oYLhAAHOcUkW5UyJwB5TWMbSsZ1JNan5
qgNSaDvkEefvoCbrhlKYKagfWgZ8Uv3ZkyEfZEN7lnMHOlppAp63kIA+8RLbp1Np0BUI0QtmrQPA
SJ2EBAXoaGsMAydRojBVA5bTeWtiCVfbXSdFX3kaauchoL02bka3xPiqyti1XaNMAV60QK8oJuCW
kfz3VNm+0+utCeyAykBToqRIVRLTg3NFr5dcxxr/sAuqjQpchfcMBvyxZosV/ZHilYjuOkOPopSS
UpWr4fjiDqCjVvUO/7o6NrpDaC308wttbEHu5cVRqzXIEdGUxMmZM6xjmHA9o20AzlhDKVCCv6En
FDenXBNMaXijzRp2TOQDY4P212Bq1skuhzv0Kb7DgXsG6FYAN8Cl7KAPQx1QNeHKTWtFSv6pPaPN
uqdIlcobCFHTg5DGSqqCbdUgfEhc53XjkRTNU1/PSqHpZ75AOxz4GlWAH9EUKrXyZALhx0D6476b
FW5eJy9/zUiqhaVI1Dz3ZcOK3woON1JOv3O7lo9TJBnGfgzvRQ07JjG0IL0p65F+ZL2Eh5+PPIU/
HmonQjObXTOS1IIuqhK9FDwwbAsA2r1FUyohqk3zxzSeAX8eoyXLUUDLitbJN85/jCtDjXrSMUOR
bpS3/qeJLNCsDr+ilaZRXpngulidqXAsf2Rqv3aOxZHqJtIlr3u7GvpjDftrGEDrVI1rk+zJzxNz
LeCVHX5FWzbWCieQNtRtT76lYVSGOgzzbK2m49+1FXy8J1D3GSRbWVUw2n1KW3ccZQq+dv2q+1yY
jT6qLmHsie3YDskZnAFsjb0q/4YQbv2MGO15nVMZdRT+wSBOFVTih96v+6IpbJcdjrWmYsZhlQiT
ZFbpaL/mteA1WCi1SzDZoRqMo9YMzqtylaknVspngGo7cko8MLIjfc5guRqTIrifDsT3dVsNZBaG
OYfJ6ZJkBNZIEDoiY1fYzHEsEQJub4PtvJtFlXlVmoh+tey/BU+azq0HCU4qlX/P1GPvB3oynsQL
XM/p9iHGgmFkjr+YSbGs0kzmwK7UYye+1O/DK3Mtg2sbTq3doMXIvLyMMc95R544sr8H8l4VH7XR
fOyXtx4z6/tCNqnNSwVgO9XmO+bdlfXci64NQ2eJSkVN55IRot8eCqi4URivz/Sqw4AnePrfAhxO
RoDA1+LrhKYu35TzojfSgvI0tOPXRB9y6nKuhjSFnosUED46ejdDollXvp8JlgNp87VbTFRGvqQw
qFKSlIWERa+G2g9mvujBUe0zrdajKqw636ajeLOhr9pXJbOaiwK4VUqV3+2KJbRGPQETkSUEO7+Y
zCdE/fJHLNlZPHkQtOF/s9X+aYbsIqQ6vqi6i9RLWCMEuzLwd34opWp6+CdTyVA1FfBEJh1xnimH
MpeM0VumVVYxcwILNzza2ol7YWj8MUhsgOx9xLKcx9EWoSrJ09y0tw6CCSNJ3JrA6EDXwB/deyLq
1OKvfpnx21mHgTAc5Zs/SpC/7tkF3VbIcb0v8RdnOsCrQCgILKhI2Pr24baoMW0Ru5EFILbx/cur
UWu+uf3LuzYrEb44K9xsQONQpjbPBzZt5qO95dkYG7unt8Y+mmwV+VvnMhHiVHvfb3gYghBRqL5C
uV9OZ3GkB+Ac1Ffoh+bDI+OJwDas2OJ6l08hFofMqjIOwitivjWlvmQkSSiLPBOEOVOFAUWrwHTL
jMz1zU4lgrHi4k045qO1eYOSW1mOzqlvU7no72+ryynuh9YvFT1ZjhXTCS1l2FJvv5bkXRtFp/Fz
HZmJfo1Uyfmjf7ODYnX9McYpKS7Ofw295RI14TLMoDNSy2x7qvBK/y5bkpwRh2BHk/iv7OEyF9iC
j6li6lBBOIM+eOH1CdGMumYmYBPb5ThVlznYqBwUIwFCV1lwK504+lZmXHK9McqTDCZFUorr71m8
8oAC6D7u74ofxcfWSsj2kX/0sLPSmq5WX2LFf2ma6n+5TAWhvIguxRahEtXH7y5DAHQuVzLTgTQP
2N7ke3FzuUUniI7YxMM+5qj/u30WUIbMNjreX9Vqndj/F2iq3gB92vW3XHaZOivh9X/DrqCdXNdj
2WWtdDc2hl8HJI9X7+3eE6ENjz95eklsrtDTn1ZcNL9bUzb2uAMjKalVwAa1lRUkx8eAW3L2LkZ+
hpQt3TSWs5VFp3Ma4m5TGMuf6ejYJ0F4YZhng2wtteXBKWRMle1w7UjZNRtylCzverctW1Xci64u
6LExGMiT//s1suPcttCxiIs4v1TEzeu3gufNqR6gIM0d61Eifc9L+n8Wuuolifi+nrMFDSxRwMWz
tlMnEkaFL0B2OlNX9QTohnyOy+HIXTcOHn0sJVN5N1TIfNDqRtXrFQZV9KpKTsLj8NBjwk0nwLO1
kzfg+k35fa4VtdHGQlj8U5ukHf2jNY6k9hzQ49AXi7h3RbHPYwoBJA7qBvdKjdC17UuFJrpv7a+o
OdEY4eTcvYNPn5DZimv/xwQKJkJzU+thMfro4yjmm5YumM55gyyZw/3M8z1asV1QkLDGKipNOHdC
UCxnVglaDOjDiNA7/9BeYTJcvn7vDSKPmL2hpZTwMCS5Lf3eXwhFy4juEcMEO/rx0AX7Lrtx7U8L
m809OmZn1/ip2iHPdmEFVy+T2rmOc36mHeR93tXlfuwEd2MqBLifyM9s6HITM5znwH4q+dEungnJ
i8ayy9Rt278nrIiV885bNm8vnVIw8ZO7KsaevOdnPIoU0DsBsp/AOJI2Plv5hSITlWhwdixp7LYx
e98PHZbCk6RRFACtak8XNty743SwthE7KNIiM0qJU8q18mpSngq2a/j3S4lPkYpvO8BfumIftIOc
T3q0qLv86mIyHQrbUZP/XypkBA/I6OS8x0BpNqdItkKFhqEzDPuDuv4e+CDniFt94o/ub0cz/9EE
UTMOoyBXIpjJLotYwlgGrS9BaUepUweLgV+42zHhJepqMlcKsda25aPKqAfbSphkOEn/wz/p3kvv
QN0e+QvEvKVHy4H4+xgjCn3+K32OSiJn52ZAm4Wru6P8Aa+u9trqBAuWtjwDmoVl0oHxo0VtLK3m
uJf5s9jexs1gxqIZQvN4CF1HOAcE5HwsHKmW6dl6tF3DZnNHUPLcA19PFI9Fpt8q6GPnvyYmodsw
aUzrUtjgjuLpg3pRyhAxCjJq0UOR2LAjVijvpA4TmKr/6TkWzM5MrgSbH75W4RnvGAGD3EFB909U
noB7auv2UVo9WGQtIniLtDXVYv6iTuf9sIcPnxgYZZwbALDIeKAypx9pR098HKDYC8H9phXSa4Iy
X60blz21h4EpIA5i05JGuOdXN5nxE7CvFPs9tVM1x0shW4zyoWa33Xee/m1DSrUUmM/u2tyyIAXH
7DyeraVI7/RIWhZ7XcE7hOsyPJQ5nlp7gpz+WqHFTt4msQWHrGqfk/INJ2sAVdvbosXupsnNim3s
bImfFAGHg1iIeejTukPWUaBazyt8+D0R55dIW5TAGaRSzOw9Op8G5l0FONcf0n91ajC49pPo6bUG
59uM80GrF+Fa5PI8GKg+opLM4HO8w9Z4LJbSGACuRcW9yNCTsSRpgmd3HUzTGMB+pE/oyrPmFMHh
MVfY0a9pPxkiDm5J3N+bOX9J4WiHtplRGEjDhjygpJO9FvdXU99bldhX04J8Blaf61UW/3bxufgH
QBsTOHRqVem82QNXGjuTVAr3Wgr7YRpFw+og8Rj9AM07GbPSVvFe/ktU0wsLwj6m7g4GPvOq8/H8
1uVXYLUMTYLRHIpew5EIZzg6pc3oVxAXApluZcRpQOlbZqp38xC6GOvPdfHhlUFrkrN3BIcMObrb
C/S1OjjpMhD2TjNghnswsmDdMfP3XnJIjmvj9/IcmS1qCvCP8GvfF6v1GZJBBNwlzImm7mPRV7UE
jFa4ST8xUB4N/il3/my+ZigL4qScDAeivQPo6z/97YC55lf4ytc3Qx4KHMzHXYdwmdlJRAgDV7u+
eEaS1OYDiuzcf1fvTZb1V2q7yao9hLhiDupP6Q/vdp7L/iGi74MC5OeyIe7IsshEk0yEsNIrYVMG
I5sCq7Dh+1p2EYVE4F63y+rXEIdUa2xRrJpNBSq8LBBhlWadVnppAWTElBMDXI477Tv/DYLZRlbB
cuxsnHji262DN0pkCI7p0p1Z3na1HIIOICqPydDPXf9PUgpJKkQxCAIOR2h7Etu+zCViP48S/DZV
p+BrRlsQXzREcWj4BpONhblFGVPbpdEv6wy0vD+U+SYcOR4mBFsfj5sf2ZtplZCgI/FUdVOI/uE1
wLe9v4fkghd4JL1a/QduYTWHO4eJiQeerz1OSwQImglOSjN+KnXJ5t0okb1Fn1+H8eWk6pN1cuQm
h7Uuzarq4xxpul6DJh2nOfgq/G0ZohUUHw9KChWXQyErLKHrKNLMf6ksH5s1DWSOpcku4VWLFnT/
0nLQt/LCQ/By2bJxkJWtUVKQHgmjpc30RJXne/IAeClUuSRHBJW4Z1QmL3IU7hiO85B2v1cq1oQF
B0H7RdwzIwJnNainHbar0ElDXH1zUQY9VUkERGPXiV05qyiYEtlF1U7GGXqrnwiEGzKx6S5aZHay
eaezrMe2pDsJcH0usbAfiBvvdM3wKRAMTp32RlgdaSE5UwpV82aqEO9eLgHyigFHvrWgroZ079iy
F/LREicT2seE6Itu6sNrTQ0pnlu0ZfsfdjVXaGMCb4zwZbRkzmTsz/1mE4Ft6cPM8K2qkrdfpPF7
qCcHhFpzqcmM3D7DRR5uuBjBK08dJOaziE2dycq0uM8Pk04c8yo94LNwABzeuCXxk3usppz2wnGk
v8JZVrX5AkRq6/IgM/DDo+N68lE/BLk2JpL2njihPs7kjyt3IRiMmSaSQETQ3cZ3v5uzNZNpGZBz
QAq8mNVwJghKQNfelgG4bF0Ddmiv9w9t0drzs10GJZsot1zrOSSbjt+nHTPF86gcX1/Mb9dZIS/b
LBCYLp2td8cERAXl3rzeIFJw0G+64cA+RqhoN56rOE+100as2+yPPfHfg1aRamcNcprKn6hCwu1c
JL1bd3oSEtnf052zdSpXgmNCKOu3VThxrM29o72HN7emO9Na9bTAaA5KtAaz9MPS5ateKlZk6KB0
u9iRuDFjjhSOZwbOSYqNyNz5bn9kX3FKlYM9SNFCe2QujOomxLuXXpzLwdjLXWgRvui4aNqFlGZ2
wUcl11CR5cEBGr1Lof94izOA6LTpnyZ1SL9nmBme9U4w9GGv0y6tp8Mou0oD3CxzpC1pw6kFqMo7
9LeYIhr9vaF3KMJuZ+cwSGpRIdTdeLyWWnyD9/BLf9Eh0zJvb2WB9QLUm5yHpbldZxgAwrFFQSPO
0T/8uwTWtrGTApAfBlBmRygFj1ohvc1UY9f+x+8ArimRXXUwUcxlkZGdZcGBQIno80UC+Nnt996E
MJXa1wGp61sP96ZeAfJSz2e19as5pYjOkPUYojBzhugTH6kEAyjToDelIu+PhhsmwZ7inUvGWCBn
nqBwS1ddYuT1rbYXoZkE5H1ugz7aOkuoO8YBchn+dzMMu4TfI+2aS3P/iYg3IeGN/pqLWdV/H3Vo
6vj4L8T79BdyAEphZipv8eqkSfkwCCHCCI8laE1XX2r+yIUTyItVYrrrcSl7DkUJ2KROjALF/kGn
3gxx3FydQSjyQ7OSQ8UxI/BJKTWqAiMkQWO6tNTncXoWZVFWI5XdAKRCnMjbDs9lPfwmFw9rmZLl
R062c/fWh51cPA1FIPOOQTd13gTkCAkBCv1oQdJbOguuAq+ljT7MTYHE2IBYlNra9O+zMemWvLGZ
CpXiBklAD8q7TKCf9FElWRVK4ett3YEb08X4FD/kbEpl2Z0njSeVbSoJPgR+O6jMDi3D4IH1JTYv
tV84p2rf1ZvSdfweKhA6IvkF1W+2t0T0uR6J+N+cCfPogYva15yfkE2XyLfOJJhj83p51vHdpweX
EYdm75HM4Umi7VxCYzGKZ0Top9YZ55DsfYUNQ21eLORRfO2Bi3DcnwrXJz6y5OeCq4nKYZRPNbYK
ppHN0IzxNa+w1E06UW+ECpjhE2BXMIJhGzJYkUevlMN6Khkl6a2PoPEpIrQFIl5pTpCsSrrwCodO
o65AN92t334FuDyadss/YPKp9n346CsoWnYxd3+Vn3w3xDD51q3N4zWUuH7WL7y1bKCmFZ0hOEpd
hDFJcVwIetyijO5hvtanreTnkakCqGXBewXOIq1xqjJDkNvPidIUO3HhUBkPIZaolhfb+AcOtdGX
Rpait+naE9WwVRKi6Z6CqcDAN9nCJXflRhypJCgbA7fGaeFbf5UBX03N9NK0MS1QodNP7+Q5jixw
sZq3OlY5fV2Ca1cpxKfT2Qe66hZrR2wwoC8NFiYS15iDbOWbW/Zzrnk0eVaOspmk80HSqRvKZSnj
GnK00QOO4XMz5O0s4q7FRJCw02EA9ZJ4oft/Rx38pyjdyGVUEINCo9swb37XZVPTC8kttqtzcH4Z
igshpHxupi5Ul/fhLW+OA/AVXcJw2/J1cUEaNDgUvCz9+GQ0fkNbiSoOtJnWUPd0NnWWn6eF5yM0
JfAXXM7b9CSfRhLiBSC/R78NHGxwPv27JywoEhcpSc27KKzpV7fqv5Ne7sbaThKYCB4yAYjW4dkY
xS20vucAiNSwCnCK+W0Eh4q78DuNHKgrfC+v3EFOKsnuEJzhNAFj9Qr+9eeoV3AkX7aKGYty5PBq
0tZub+ix/Vt9IKGguv82jaa3oXaJZM9br8cvBm84dDx5bMf6ItREuSG5zowQCUbU9mpfN+4DJ4mX
sb4XghpxvS6EvlhLJ65LI7XNTARPUw5TclfmMdftSWxpVMXJMgJ8wPdJ+iP3J2Sc3irJJvheRUnl
DS2YxTDWPkpF3mCfLZCuGeVmbWLnW8X0S50OomqKVbeMFWOWzVHk17x/Qxjs4BMjLx6yIQkuH9Rs
h4pYo8IROi2LsrMaida6t3TLMOXINfUfuzjFk/OKWRlG7Rf9Z4waNKluo09zsdDvwW3h8/XvI0KA
DR9hRWAvDeLte6tZVrew+awCs0Vq92ErJ0nlZ68L3Wbch/cUyWkbQQJ9VRuZpvJlwvOt4XY899UK
+5rbtahK9NqHeMjQBeQRK5/MXtktt67HF76U+ALbCMStQgmwFy/M9W6g5OFtGRMBfSFwaWFSw8M5
BWnMzNNkMy8RYx3MYTngPcjAJU8STUDUWXkEIGdnuy4FKZrmpCqqhVlN3QPx2e8TKpq9HV9XgPPC
6dkuqckNAS+OTMVEeE2x3ojyC3BXZUnkjYogyXAg5RBVZXqpZ2Fo0rtLx4n2UL4thIo2RDSwIaHc
Px6ngF9o/x4D3xTAS94+G+cGx+hcj/F7aGN+9J0q6QjywI183pENmfuecDL5Bzwhj367QJrht+WI
wUnqiBIpvMcjnM/FD3abXOUmbBfYXgsUfpTWmF4kMBH1Bjk3roRHKhSnG2EZXC3eMwwjfCiot7bE
yRX9O4I+w+yIhl5qUt/a12d+moqUx1AU/QwLpk6yXhfEcP06W1Tmm1BT6M+M9JeDidxO21wii36a
RjFUdIw4rdh5Zi4COGQkJkc155JPNLzx7jMjqWXIrCF8ABPEWipcRatGZs+85KyRwsjEyRBoT+Wu
6lbW2ViZtWBh4k8lOfo5wDr/ckGPq87HzN9iKRw12F3mQhQ8ImHWMp0v9eWU33kjPlD4bn7xZX2A
qycfRKb+wXJgJlLWNgElpK76Nw+pfA9a5UHI/l3nzSCwpNnmBBIk+jLYY+39m7l30OORk40yy0en
ysW4Qgu5J3Cd9eOOjLfJyhX1EW35/wLd2Rlt/tsdtHMzwXTPDVvj/936Nkla/QQKsXcSKSFFT8+R
9/lUqf9+DfweA30PbVOlFaQmUG9SkzkkFBTmValVt2NbVr1E22UKWsC10ZBTHGyL0m3vlC54YxWj
Xrjvo6wkd+vTnSXmG//OLpG6hmTykNfQjr5914PHyHoNhfCsHBkJkUynw9J1Uk5r0ii10WvqJLri
WJX8CNi4hjqwctUDSfDeZoSatsMpg9HcKU0hIWHEe76sQNkShRRohVroXQO0UyC7xQEa6R5Uv2i9
mO6Nrha5qsgSQkHicES4g6ceDScp9sqC5LRxRTU3jp0dFf+StgXg2eR8fMNbGlwqTetoh2iRjTue
tASyoT/uw6Jqa8vQsiw7VnyaNYZ2D1nX02/GC/k4fnDbSv1T+mPxil0O9ihEo6BB9tYTnq+S5QWP
fhe93jozYEJmhPo09vSY+nya6wJBDCfYGdX6yEkCkKgpOcyoXoN8K8w7PqcBtQMDzGerNwRsbwU6
JUPpWCaYpceAtkMonGENBrTFdPGrH68FrQZNORvrDr/cgWMG+WCUIUmEUWgYM6SH1ky7GlIuhHWk
Tt2qB5achpr76rZ2hs8sppEFiIDW+I4CsOxaxKyGYlCmQEA31/I7bJjY6QdNrbbebxxIaffu/8hs
naL+/oAx+n41fqJXuEdABzSL/ZnlpLVe9r5R8dKl8iP5ktiuuspq4auF81SygQLF2QqeJRDLQ0HG
IXcK6hnp89W5XUy4IKqOtfvjpu9WrImC+1JBAsHck+jsB0TrzmO2Wd03VCgb92rtfp0irVb5iEn9
Pw0Nt+SMzLVL5TCs4b6fDPZjtZSID64+45YUGnQjnXASpPhuO3Ll26sGZYZPpeiubdRi1ke+TfA6
Zr8Z7ntaLSwPkJiJYZ3HQgnbFYh81H6HfXxRrOfeOvOXD0Jubp9bxKKXkU7292MZKUeXbra2wYDv
q1JEOzIxT0UKm3vZ/OvfgQmKKMgnQNbL28Q44/8l+uFpAJo+SxKrgIO5Ja/wjzzA7cU+ApB05hD1
rl0azzxEfkTdG33gPi9a2eIyrtndLBlT4A4JyeLQ3riowaEdBXNraA9uy1zJ9N37KsUK+KNSLrxk
Cv1LKZMWq58yGaE+iyTWBLJDPeCIIxerHPWMseKhEOHXKUk+lkYL7rjX7d6Irm80HoLeMeeZAOhm
2njj9Bvaed1fGojHDypN0zJcDWzYne7otUUIM1zIXjkpWrSJXeHG01DswN6Lqt4K186RPgwqnjRy
6wR3WT1Bkd80WiDgq+9QDuz65Ebq0K/1xlDVlPN4jT+HwjR4sBI3Jq8vG8C/L2qKn+gIvSgHOvkF
2WArnX26sPyJzQtNLEMzAKZf7rZGhDMltQWtcgtdjQxJCYTg5Lv1RtD/Vd9apiMraA2i/PCt2gbm
ZRx24h8CzdNerf33Th313ZNuoTs8D0xAOug8ZRXBKbFy/KWc8TTRFZ/YjUvnumgjR36+Q9I1ssi4
QaPfWwuAw4J1kt3iang4e4gHfZxFpBxWJuZOLwqdb8tbdRia3MG6LNQafT9V5m8u26npIGQySL8+
hiNycomNne3rpxMGetDuMMrv8RZjIZPzL34KHAO2Hfd8lVUfIH9ipSmYy57HhoXa/+JpHq7yDXm/
ECMHO3dsNe3owARJp0YYIQaIvbSFl3NE2CVlZg56aVfVeI2AHRia3asSaZQ9hiTAj2QXTI1bbS35
C8mAUZHf/SW1skRCG6WTLkPa+1NG/g+rjZV450Uv2l6GDbolDkK/6EO9ZIE4+hLv183zoToa7e29
B7ZfqW1/Q6oNOLilZ4WiABo43qneWept+WHchdbLgtSDSPU9hhpfF2S2auVF77UKPBDpNfXZi+Zn
fBeAyS+19jtGGYtMc5iFe5eHtPCzm6T95M22M18x0gJk+iLabtvZHTvUB0YWL+7EPadJ72XrjUPm
7QKqm59ikqQDkoTg9CI1QS5ivGAZ4bSlP5Oi13LbXDRz50jw6YJ0AtptcBpUEwTmPw2SlFdoFZeV
3b8OosNi2G6TgZls9eWlvvAAT715nEX8dVc8NigfP7BPf6QLa0FeBizuIqSNrnqyoyKSMdfST7pr
ffTogAGaGMQCClomnPDiwlCbtd6CWyw3XOL1xrHMeRFPTsZ9ldC4A5EVzjHrOpW9hch5kkZp5aMS
HRVFF1VJulfufeqAcqqUuruO8DnaLFzB7Co9kAgxp/pAJIXlYbEmdRGoF6D3/tHPne+YqP4CUQ5K
MjeyW3NOU3nQM1BaVlJ1JxZPXLOfuxrv5LEx3UXc/CSzSKAnCpYmk/GXVoLNv27rOvLUvg+7TdwE
K0bKevOoloKIf/a7PNMlOsLUfRQ+wArkYGYtukMT4bB42X9/G8y6spAf/8DDiiczk/8LOIvK5OZb
CVts4XWaBxmMvNJbuLglnfOW1EgzExAzBfRkrvYwCwGnZeDzPc5RRndVQka6FCQM9UT7H5mr1XZr
/11pfrEWya5LlduNtQk/JiZY/BdvDW9ClOlmZUPR4ymRKlVDOWHdOeaAQ7UQimpjttFBJUlMU2M0
kJblQNS5Ay/+AjGQbjy1pTCZara6+dGwIYa4KBgS55A4gm5Yh/O+iDPbaWvhaL8rcGVuCqKS1HUo
687sbURHQ+rWiW1eGUhWMsSmv07lhq+lA2zuM4oP70O45btAVaDTBXInBrZb4r9jdK4jxnndhvtH
eJZx/OSt6FSmOHeuRjmTUAk050GHHwLS2DnzioMTy2gxjwNUEpeiExwsQ9G2R18izQtfAkxPaACb
pqXID9Q+v0BCxTqE7cjcmhQo9FQ4QZfxeTpI83/W7d9tRGDsmsdFAtWKBQ7EtUwupqz+1aST5vbE
dayN1kI33/6IyJtqebjZB5Ua1x8bRsIdQosMy56zaTsciBcx+lID8S9HR8Yu6XDxNKWo0NMsRr+/
75MSGgcfYIOgbB7IN5WMok84LolLImiIm6kRQ+38EuDPRyOoOl1dn9QtmN1Xbdiarzu6bhYLIZgz
foskofP5woTFWbKZKUcyErQ4ydSv9d0LRkRJnvKJhr3AitfLoaUvXaqwHRHCiQmLWcgUSn+6yyWY
bgkMLxHPWzL/EVkG1jUyG+eryO6KWzTIlBgijU0H2nd52ekkOERlfScBigYNezi+gEskRe2Oj9/A
fqVISkmpnWJd0iYf6UlqrGRhHE1IVYO2VGZGaoynV9+NnLh8mMP0qjVQxbSwHPNwoCsVuXfRwpXc
YV5mXXu+pEyJfgMQy3g/1n9YqftMdl0+vICKqM355/77I2H+Yupc6IEcZ7xToWYJaDxnmvNrls6i
z8+A8eRhCcSHvixYCdTbOsp5Ao3F/sYQGNBOF17QUp64Hxlq3+h6dZh7ESM2uS2ROJBwZrtx9FlR
BOy3gipQf1E8XEFWtzXp7evBRzOAnF2EzD5224NaNQMD7Xu2pJu9P9bLLXsamaS1LfhPvK5fez1p
QH478ZUkhycb+RI1EjqhIFVhyV2GGzx1bKC2CqA6vQqEIFwJPgR20YS2jDFYvrQ/xncGApOANgIk
06g5ls3TJQlnLPWOZk8nP41bO/lQ5BTyVQ5euwGyCItEJdXM0U2mZGqx8tdUDHH8UNb3VdRPr02i
MGXAIBXKEyhJBOFy3GSFj0XX+ckjqU37u5WYK6bZE1J4kFtqpRzURxCuZMwytlzqomHql3qIz/Tz
TELaDLogtzrjDiBHfcFv7yawcfTUXwcCVFAwbHy3wJ35dlHEdu9m9/WvLnAJS7pDqOYtBR3K5PnK
ikC8yTyAT+WEaFkA8J/mIKEXjL00xJy8dJ1KTDFNf//zL8tbneIji7FqTUJDArkOn1Ml9COmQBU4
6XZkuy1DaTBI5tMj0Y1E6dQ9MFyNugtSKgCP39InuxgpTB9JtlbqZ0cI8YQ5QW+5TiwjrN/d1wyU
SHYR4DbwdDC4pLvfEIYrSQsPPxfy6H1zs4IJaoaLy/CtnhZPRh0D/JwV9K/KSgrwVhEBar6Owy/w
rWRjbVpaXF6hj0N1BaCB6Hu8bWRy0gi3lgVh2JwJihqcRz6bnDLdQkjiw4a/KMmgWcmb2vOEUMd9
lYRQWu6lclepqgV6WvQzL02Vrr0NlxXlpVJztpPgthgabM54ZcvdXDuNE1+HCStiJQTRfNHVsJ37
EFFtzgTRaCw3/VLLs4VGo1EKKRndi9J+2BytNoWW3kvUfyhjVxaZGXvgYimguo5XsxTn8zXWIQsf
JC/AZy6PfMW+uYp2LuaY+M6mvS3B0WgUebhQAB/Lme27RBY+QT/T+vOMQgcABNAL9DU2Xe96mSpz
hye9sE0F0Y3++uM27JzRZv1IqjOK5G0XRLZ4I8LWhA2CF1CHEMDGT1lRsvbF4wCj+vipFb55Yqp6
5d8XzDw3Eu8LpzN0d6VB+OHDSFPwIoD417iTQx4ydoRm75ZOcHTN/ku7mezDAV+QX2UWFIJRXj/U
AJ9G3hMSH0lCCoLWCDDpItAwNvEp1GjUZdSYWm/8yjvAWdhDJieZYJcDxa2IwSQyuJnz8uZeoEXN
AK6w+bD4eEarZxgCI09ZW9892xaHsQadAsc0R7mr9gVgNSd2RzKNSpuPaEDJ20agxxlBAgihJw5/
jerhwwGIe+h6x/Ghkp6NjkKtAeCSbiYHM5MCrwNTma04a4NAV5A8hB+xZ2uuo3K7tWjQwVGWQDqb
wkYQM++Di0nV9s8A6TZE0rKz1NwRChTS/pju0FQKOk7ikL/ozsEqeSPa/ihbde+jMEqNcoLYMUCZ
vZADYyd0HJ8h75gzJNJoXfkPISMwaGt1jYMv08TZr7dYe77t/sILpI44gufsw35JgWho0gaBgPHT
S9rLl2RcSRXm9wnGmLokjViAhzULdKDEYC+XI3IdbZA1Zvzh3DNfEQWoUUU4V+c1Yf0Kj/gb2/dY
XMiUG6HmWLm4FobtCijMv1A9tGvBhLZeSojCDDpThuC+Tl02xBDwu8QbyCH6tFEUvTy5ang3xrHz
jCRQHCC5ihRDCSFGmRiXT9EwkRF0nsEcxO4o68OmtWoljYdf2ymYHWsTD1UutADIkyB/cHk2q0SD
RSi5X6wzGZLMYGnMW/pSy+PNAjTbcKmngbX37Lm6E08KA+l6DRY/oTk9lVTwXtXB0EyUvjVRkQkx
HBTjPra9Pu/VLh/0AvXOIhvn50Y0uYeOtCX4MMmu/Jfdl6E4MPnix6ZZWNM6bHVZ6HGzX7cbp1fs
vC3TdmA5cneIL9FcYroqgRWVR+ehUQregQbUTMjYGoTT7DUc9OITs68dMNMtEdKJXPIkmuMOJewt
WcEL6Y9A3aPavkK4LZCBLHGkoy8WPHPFCDIb34alNXtobHmVDOmTSU1vhboKCTwTCpeNuwEnFoLG
hm0APH5fSK7BQ2tP4R2SbNiQuMB9yy9E08arVbJXw5EyEWRlIyS0mtbk30oupHVodD5KutT1gTlB
32blmjNIllU7mv7LRDKHnfGWbXlvn1u0o0NfKoqeWrYveZnLacaycpLSPSWSCpwcY7gN6KqSu6V4
ST720V5RzYR0p0uZbR23G67TjSn2SctPkUIw1ud7e+3TgQz6cRJICEZjBwdXVhxVmLNrVkVEUCdi
3r/7qva9SF8TRrT8RweEMkU9dojxU3d63kEt7N5NjBjS17urs7tqP3Q4bDFOEf6PLUqfEdXo0ZuT
eJ/B9ICJdNdHsAT0Jw9BrdC15v6qSnlvGiZ+xZRFmHA9tXEMjsZRLK9CjAk0kbG4a/c9/pxifRWG
3NNtS1i/Owp61tmIeLR5JHgIXLDvqkEC7xHpQPGIdHzjrKEK92gcLc253uFJhIDW/6OTx5PkHW4d
0v6J3B73nkib7640T3tOVxKaYlODBNiWKgW3LPiCE3hhhkUvDQOXUck8w8SbcXCuVOJQnA1JYQQ1
kZ5AVmXIvcxVUoWWfbz+J8qU7hmMYdL0lcl9POIDB76Nz3BgV0yIWJSQtMlW2AMSKDdyEiTmmFIm
gc6lTBWZx2YG7daTE4qo7WgSirP9D3YacvzVMxQC2X3cDCM3wvhEEByM7GJDrG4yzGbwU3Iq7+c/
e7ICSX3YwklzdVoUYETBM5E695tIUxMITW0Ip5MwlngXB0oOn1D3YNqYi+cBmQFc15oYvbnpERuj
wNS6SWYjX07gunkvqD8y3aXPxaDkGR65tyYOUjnjPI0HGSPMrshoq0jA5CKhdpRFAeV3N9qEie4t
ty4WTSWP3u63N1RuUlB+jhdzROCE1tKyanqZVaseMNLi5QbXCfeT9sM0AyGhH+Xp1aA7HIylNkxA
u8OV3D2TEHhmgsv9/eicyP4loDhyhx1Ld50H0IXGqyuLMfZSbY7+DCEXnJA7KdJnBmgBrDHwenkL
XL25uUVCPu7B6ziNmixXyFdNLgM0pOe6+7Kzcyi7qXKR0TZQ2KoUS3TnxLOCrkSIfeNIBAgZmK6j
/9r7uyQmgxC+WYkyu3rIUSwVJktgQqg8F8xfgvBpqjs5mMAdXeHwmLRRJfHzzjrmNwGz5IL7vpuo
SANR2Acvvmt8a6LgC7mOv18WisNTQOItrbbRARQlx0FUt1wL8NaV7sDEpkkbD2VxX2XTZsDl8Bs3
mvJ4Dlot3rgXD1svMoZDvLzuHO0ydr1QVeixgC6MAapIjP2kGfxhWUFzCGODp/Ddvxg6zkgp2O2r
0gAARwIB1mgud2rN0JV9vjBVtRmTg0UtnJBmD13HjTw3sjetPaktGcbRHV0+IY9di6UCGtMdMtHG
gm4o8AOkQDJNlPxrg0h2AQVN0As9HleMjzDZ6+dtTDa/CnelEIB0qOa4nnT5qVj/97tDtHLbg42u
7UYqMfdS/vn/8L4xZyLeQZNaWeo8WolgUGk1P15GKWfBmELTGMVx+Sc6SOuEAlFhIxYLnzecYBiW
v/t2gVjSP/0aaEA4X/j9spTRfbE3vMOBEoEsFqZEXUt5dz15ME9N8/4fpGnM8zKB6nSmYiGepKRW
ZYwcDRgmqeDRNI8Ou1svKnMxd0Lmk8Xq/GlFzhMNNA4RQt90hgXkhRdyNjOQXHJXDXNP7SF69y6Q
XES6JJL8A9sTjUa5hUOH3B7fTDDCT/EHwU/dh3LkEITH4zpDEHqYWNtLwCsEsu1mMK3fNXV7PKTt
yj11i82yt6VYMxltAAqxcblLoaOibcXK9B31vMaz1O1wkCfmOvSepeQG7CL5+EjpXQbYG7pq0k4G
xNLRYgLT1Av/FytMqOPTyuih+Yrb60atIohVeV0e/q8biCuUZluqCD2y0PmzWHIXx/LMPYKuuhMJ
YhCh8zIyOIQ+TNSBnE0IQMhNYwaQQNoZ4aqZRIhD8d3HB4K3pFaw8UJnj5pQux7oe9maO7kPWgIy
QnRWeczcMZBJOFj9+L1e9r1nptr8pwcNkh3VZG6iD45hG3j47WYKDzj8CXVHbNhcTqgC3zQ3gorV
U3wFeT56m8bDDcZrkhoaDsSPdUaSSCfeVZ5z/6TCqeoj2UX0EELQRyspbB6UlhfMGA3l0VeLf4aU
T8VaYTou6PA0UKstP9Cj3O2WxS1z3XWLUoBXJuhBc4n3TQ7wcwMhhCCXLTgj5mtW30hsqlIrdxcO
OwiC/VOIO8/i2I3NKg1WPbAgWxtEW5D7ylk3DCN2yylgBTf0UotYl+mIQzC5Jx5Ujb+k9bCzzmJQ
I9elzxxEAAb1ZL2VHhZQjm6QXesAiJjTNcSj5c382Mj1OmCLXMgSWPAk6mObQ2SieINF9dtJn5NW
A/OwgbkEh7hqoNlLZ4ROpD60R8LV+a8SU87wx+nQfDCGsMmtkqP99YnCh1ZPSJxf4FyQxYJqz9ZB
XzMTBrIKGB5WbVhQ+X5VgUgYRRUo2fXyW4IbY1v5airIIffgRkz+4udgndyaLpL6lkVB0F4oAdRa
ASgViQtYrcRhrNcVJmxgHD4Mw52D0ggqZTF5TgeFz7D+b4L8s5iD0k2LP/UCgTFfIetEs0Xd1lvY
dbWf+7Je6uX7S6xQXrqws9hjYwjZkbv4E1CEL/xLx1QSsS/2uvC8r0lcrdRNrSqCyD9O3jAJWxYc
HSXpwEeGie7aM9WdDFYhqcz40rlhEVKtDwA4OH4hNTHEeS62RWRM31ysxkvh6DoAEEl518DeLenc
gfbiHdqUneTKI6DV4ggenwEWhT1dy/n+48OoxavtmWC/3FNvwqXFC3CoF7jdz55YD/x7w0bYh1X7
uBYf+1X62b9p3Lb3fsC6epsozBj23dyLHvcNLeeCtUV9pDwhsCgRU3hTNrMscRjXKC1qtTNVlMFs
VACAI1evfSYJTkX1/KQgfZ4x8Ttr9xk7n2MIvG0sPqX/HVzT4yuILnY7iCfg5oktc7jNUt5CSyuQ
RIlPX15pF124d6o/jiHiu0zUowZsK+kj16JsPKD8w7LliH4sxNuWsUSiFRSBWDJb/nbclOdRMVDN
vBaBknH1shh1SJPvOBgycnanVKC7fwDUkpK7fS8BJP78bQ6cJUi9WzJl0hqoqdIu63KoJd3Ji8hv
D3Xm8x9q+jIymxGjhT/oT56wcSUODZ/SEtRU2pNr8VJLarEjmiAAuyL7G2+2zoo2nrbCxC480mqa
TLZyHg47Uj9k0wCG2+5ERV3VVW/r6mqdJ77XOelZZ6SbafPd0eoNKFSIcjbDu5I+6uHCWqE+SALK
5Z7szOVuIry7a7rslzU5sBJlT7TZ0YqgbYzBWh7x7j0qPXJ45cRTVOf1JLJIgGTo8rm1Yzrv1bQz
yDXM1CsduK+mb2P9d5wwoEBkmZRas2irYkI2Rkt3NlLdPkilFnJ/OVJO9qKWmuf8r1Q+0B605qgL
k7NfDHFbxu4r5JkxJMveZKfwT1h2baA8OLRi9jyUD0jZOrESTTGN84BQPaxGXov9oQ+Q1yrt8p83
1p82LkuyR+kKlv196jWKFhHtboPihcyGPaXxVQA2cfasSL1Gc+7lbPaXMm9rFKiGTVA5aY3zblgs
e5NJJP00XKX8oHrOzehscwsGWGQZlQ2qVMAXGNEM9Mv9vGmRX8kDvHhClDRdQwlhuZBAgHhpVqcp
2r2dtPehxJiFWbBZErkGTvIImT6XkSqOIDgsp2FAnpqgq5k2FktUW75rj0efjr60ddRc/ZQkSAEK
LkUATn2mhp2FYFpnbBpao17n9X6t+3HPV73kC7O9uVjyveCG6CkvYzWzLKL4eB2902Li4Hxz+jXO
n9uYKnDQ15sTIgVE8WIfNmzGWh5lorqY4x/RH6TA1fiWb/Gq6GnKb2Ic2mBrR3VcZZz/wy8VeqV5
TFtdJmAVjphZ2dCHyy5t5CkQ1siitnxUfqp8bEDw7uLyRbYh2tgwwtNEYCXSMuo4wZXD3O0IOdtw
1PrSKg/r+pg37ktoAx3RAFexhVrX3/rd3vKVSVzb1w0TMko5LdZvjVN47TXH6TjJ8TGywDO23tFe
ws3xuSkUmdGyCiTcpy5dffj4UOC241iweOVQn0OU3nAtPjaAhoILFlPjSxlwfHUgm/g4/t7kpDLn
LT3ugBc5YjMgq932NyVrhI/48SPz4jd8VpWdAUaVOSh7rJ73bBwBhq0Z6MwGtkvoF6jWAYHbgFJ0
NuAiB1nUGR6qjE9HnyrWPQUqIu8rXN2Z6V28A/5Z0LG83mkIqvl9G/BmyRLeGkgQzvbDGGQazhxP
PJ+iVT8hruUUTsHdpP8LEuf37rmU70Pjp7PodSBYTZhCOvuoAyCONkOyaxMh16HMPdDRABVWOTI2
f6sjtj93buvfM0m48tUNwlr94AaOuQF6FVvO1rKAI8QnAEa3uQWlY57oyAZzQRJVKi3ySmRNZ014
4iTGcIRzebmfpr+Q6/hl8CuqOb1hl0zSa9UhSJE/mIyjo7wUmn1BVM+oPkeiOkwjcc/5gNgOapVK
N+nNAPf4HSGkBe6t0BRcZTsnEMwF9J1PzObxeFc9Hed3y7/+o6wrieHhGUdq6ALJfDwR8Lz1bQxX
hQEY5M8ijLaa0T8QZwHXNWn6BAjYJES01gxSJG0OPT0FO0Vie+ah04g/FWi3e7o4RT2aDVRU4GM8
mEX8rlBEIXNOTTMDVN90ETqc9OBvFVK80lBkcH5RLt65YdPpgO8HR7SsDrazdmJW8vQkU3wnGiJ8
NdS/XvVTOfXpmN/V8os3Wn5xxukgu62UEiip+xRrgn81MJAr7Av3nI3fGSPZe3N0sZVlK3aKQhEu
rm3CEuA6um5cT2Wnh6xl1QMZMbYs70bIAUmRQZn6PgSFb3HngThaAZSunyc6mc8UNlYrx/v5HtJA
u5qgTa6NczqwHSzs4zVD8Dr2YoD09Q++IVGccWtzjk7tJWms0tVkwZ8W5Pf3d2DrDRdQqhk0npi5
vkERefS6g1Uw9B6up6JRMC5wtQm3qPBQ+gsIYmgOJRxjiWKgdxG1Yd5oj/k7Xa6gk4Q7Fph6/Vlc
saxRN9T3QwOiQmNwCu6uSo/0MnH0PCeTtk/lhUdqOVB1QUtw6iKwKRvCpIIKFOs+zY557caR2cxA
Y0BJI9am8dx7kEZV/s/UBUw0CEjBK8AHp3eRP4LIWiP6iFCg8CPOrtfJDo6/udFEfCCiLxj1WbBy
CFj0gOO2ZvkHA9yXEKWTvOlvEMiGa9+cCjRDJvtS4sWIAFcJhJwTuIiYVHw5ok5TQ7ESM5pO6P6M
cl9YQ1Uqbl/owNjNaP6FP/IUdETQsEuL9UpS4CAGPrpXB6GBFp1KU/ZMBO+mOJB6nuh84k4Zc7zU
41njr8VHUIq/AZJTb2sFDtMybyZ4xEofnulaee+YwssqGuxrcahqew3NBfR30tfOYQBx4vThSnXq
KR0Play+6IJ5KUMs4zZ5H7kLHeUkZAWDKLVB8RyazF53h3K9DhIUjW4HSr8kpYYTdzUoa1vN+rut
lmRh86r7NtJcc+xHGYFLH95Y3Nz2GDog0Qn6MO8Pr1mzgmX6+nOc/3d4jZTcJ3fmM9NW/LM4IcLg
RD5YpUEX+raJ0778X+ytY6oL7p+cfuAu4okhO5Cntoq1LSS6METnrtOccIO9hKZ4MbGGbAL+xF3k
3Q05nsOMN87MQkAf7qD1mrdzDTT4Tkke2X9FPTSy+CAO+4LFpVWLk2XPQd+d+R2Qc12RwVOkd3O5
wK0u5Oo9+gF6BlWjyjG621AMY/z97jhyWeqsVBYhsYjYI+3udPbQkLVtpVg+GqEHrrsv4SE8gNlP
1tRnT1V2FMSZ8S/rZekYnB9x4qziAGw/7P0lDjTgewgFXTR7mv+HkwyhX8JVUQ+/ra0vpyX+8pRi
TK6t+VBUSmG4YTWg2Vr0Vq0QjnQI5S2WNBUrfAuKHLzGAGTu8/uw/GxqIk2u09tx2vxIvPkCEdev
9eS7j7JX2TYd7e3SyPREsm8Jo3QQcU42+4GKg4pOY46RryqNl4WmgzUO9RBUysYRLGJq7T55T5TL
7IVNcdRAMclyLDBgZEuT9jeG22yK8hmi79pvgTPrVpTvA+uofFFh3Ejci0oR8G4pzsen+yD7Xu/X
tMkurEU6xxut2Z430GOnvTv96n8xoIJUnCSjvZilNoeuMfwDIt5e30fJ3Yhowp7CoOlviETvjetT
7CrzLUwTFdJR13XPQlCTPWX8XVUXN3lcvro9f4SObd086CPVISbRynZCuBBr+Tmh6Tir7RZXtUF/
gmkkdEMgheYac8SbFqr1I5v1HeaAgJGe5CoPcfhWS3vBBGJ4vfJpQh5Fv8J4gRgQ1ireK5pPLuPT
N7CqF6EiouLJM+jr1KXarJvMZcoArBy8NRAblUTl5sV+jZU1kqLKLzUgwBz5G20l13M2JMedCy4C
3soVvP15cnwCpaSAlRajzOHBdTZrpntvC+Ol9gU4GfVsswHW1xsGQbDQsTY1+axxY6qqAxucAAH/
U/ltxWExAwIOqvlkjwuUG+QQ/V4UJN0k/uvT7WWnKquiF0BSFTboAjKc5e4x4GVdJh8aPEwce4PX
VQwi/7DvHSFUgEYUMzvo9Q2NwNPtbqy5NbDjyU/MMuvIZWC+ib6tIK3cptiCsJCry5/+bls+X6L9
pi6n3pe4R/UTybOiq196m0MU4tUNq05o1p0b0f7UHJhb2k6224btFpqEZXT8CQH2P6lJawJmpDNX
WY50RO0Lqye26Hm7SYzhQb0bw2OWiv5KuwIN0TFkxMtqXHoguQb2jfEc7bFNSSj60Vdi0IRG1a22
wXtOWsnEmamgWBAtGUJjqwwOQubYaUyurtzbdM5VTLRmNijMmkDWmb5Ob1M12B4qU5Ta2bxLlSUS
jGQW9pjwQNKxb2WfkCQqhLkdb/CJi6DE62KthmN795nXmP2iq6E4HHlCafiwfisSYgEiIkBdWiB4
N5LFUmbhztk8wRO2Vc+7+Bf+TEYr0D5XYy26TfPlBGdcAdwOYDgf0oLRnD1s5gLxT7AzbeRhayRf
QVJM7M69f88byNUZynYWVG6TxS/zN4zhW/wJxGPHCKfhZ8C+6GDIvdK8WC5d6t8jZvstd9a80Srk
pBugrGowm3+egH2YGBi01ucMesMoEQswOUGef5hWOKf2MYzcYL4msX8eW/JJ6Ng1VAp3Ew8QKeEG
ltI/nGji8naCw+g5TCNPM/27jXobiJJdAty8Ey+gy/9LZzseLmCS+9VYsq222byaTx/UklaMnG4U
GPVl8yv1apLS47FLr1+D2w0f3Pe6rXWTVqLzic0afjsGAug97TmypoclCKdujC3vGppiYD7HZsMY
llZv4VvXK3clZ44qfxkY0+4tdUy/XvJcaTlGed2+Eh3cBd3NJub9FV0sqtNa6yP6NiEi77IfqZEy
aiCVVXollLP/ETfPSlgbHBNpKQSR2unSGrqtQNgHGDGS3EGaExvyFt0kOD+s/AhELCiz4IUMha7/
35FpXasm6yLsW/oZYhB07SgeAEklI65fLAlXRRD9Yk7BHLvbDx8uWezaVXR68QZMBdfoLaKmMtpN
9FU1ouMmoGeFKBL/fve2vZ23Dk0GfAe3wi5qlnAd0x5SxpkAGTTRMDHz1afzAyZcScXQ01k6Fr/r
7Y0uo3P0sVTUYJHRWjhtRawtVgMuaoTZEyU06TMnVffY9VIBliQhkDzyI0VJ2khnV2ZuTaAF7aUJ
+c78/gv90ziNU/XSJH34T7ZEpehK3J4un4yp8ywCdoUF00Aw+i1E48MPAUfeVbptLFOUmknpBDYs
ol0lHGX75r0DdqecqnbJ93UgDBClNne33Ix5Ij6Cf2vMsKmjHVsuMJivEPvfXNzK4CEa3Pe1VV18
4i1iFc8p/ubYz7L/nYmdg94ZwmmbCJ+GAOKFNh3tSjs3LbRTcF0fFimVFxfXwm9sMhkb1Ux9yApY
Dbt3/OrSfQx79DflIKe1EAPgaJ45qyjayAFXIK5OwyxEnLNiIDf+zfqDsRmnDKM+X57qEOyPNuMX
eFG2DwtVzvgVUHRQFv0iidsktqAVU4Tc2JfpmXyRF0UQ0+s+sC32R/4Q2SZ1l3iDdk5StKzo+Onc
Lel94J5I9ze7Nbb/1Fxs/UstPFwYsnliYO5yb/ssf++TLUibE7TYH7+F6BGjGXG3cd5L77nGWvrm
Uj69fdbM4d443rL44F1advwWxqOtKOoZKePRVkQUz+XrUqz1G9+ZGI8pfhqeOCYNttoDH3AKprxr
5jDdL2Wm3KSpB/ZKpeuZBIYjFecSNrm35d/GfDeQu3Yb3e200/3GvVdrp7T8zU10xjYM5V7m9nfn
/BxcKrRIyr0VV6LWfh4QyhFkWaRiZTu33nS1qb2HeT9t8GUvLXlRRR7J572WhsLnelBKfcMBmj0f
/8N3sTqZ3zqoDgN27OjYgNE0eTZh4K8T3enS5+cmv05IbiZn2Vyd2VFDhcDZEFCzxXRAUL+g6F7H
M2U6K7IjDQOIwmMM2QynNqrsBReIRUjPBq9EhSwj6cnBE0hiQRKNVkJCmTiO0L27uFVyVX19/2w3
w8gf8NKSCaSq/UeYswwjlIofCOSRfBprULSe7zwX03k39s+T9z6RM4Y0tkO7LrXxZSj3v3C6XWgg
9r0t5dZLFRKKjZPY2S9kktC9KNY9jxDalcHbli2UhgeX5F8HPCcwNA2Ke2f6axS+XRkNjVTUkmzx
sfMPHRJIWMjFgbOw3z4xpGA3kB6AMC5QSRtBGUt8yU+K1DepyPyVzxIZmmGGe7mVxRWo9HqL1mWt
lAGFyX/Eq+EU4/urGWRS9Xkf3tP3Q/P5pbvRY7m8Bus0/vh2Uk7XE3ya89DlzjTGhjA0wIeVbNJQ
26JzdRHbU586uQhVqaWudm5D8oaPWoNmhjYPxXH7IdK9kJwTBnd3s0OaKjuZcRcf+nf8VglCXbOR
27sS3AVvP6AZCZ88Dw3LIbfyRCC62tBmQcq9vbh+yIQ7eOxPLFHF1IiMRTCpdWD/9XUqWrW9rXhG
wg7IWQmwrHnI/A+TT4oJ2PT7eTq24Xeh6noSeFjeioIj2PiepcyHEpGy9Nq2ckHiOElgrNhgKaWi
OvGQiIUcfI27re8ok9YGQPhyKZo0xqH0HpAHPWLBkMmsvs+SuuWY4XWrjUbpIWPqd4+h30SHQAXQ
dWFS2ACncp+hvbQTTw0nr+yfcbH/4kPCkWXY+/0C/KsZ9PtJgcfz1LaeTxVw/hSKO8uvqNq1UV9l
6Lksug6v+RMWtHmGIpYwgv9bWyOsmtmbqdf2nHE+I3cWt5o34kFovFU3IVSy5FnDOwXOo90gKP8s
tov33OdXoQa58o3lXL1jSkA/5FT9AehXOVuTK7fGsu0hVm53holdKFspHMJbNB3tQIkKH0d1ffJK
CR4LME/CMLxtPKr3wnseXEI2bH5kSKvaZSB/cTlqUklRfXgshq0M20lKOpUcw+OGdETbDOIV3OBk
8EfDwevJ77u1POyHvZAtncqbAJVikQD2j2/mpY96r8E4Ou1PS0CYLNosOveMxjicCiWMVY8/4HgW
ix1a3LWnzpPwIfnbmukyVzAyz8579LC9mEm0oCixtY9sVHWqPshmNQDAtvhZZkZps3YnwtsOrKJo
dr5Rlue/swJeTmf4DMUKj5mPjIdnU+HoOqcV6RrsrQkS7xBTHwz7JeReFnTteFK5Da5dxAxzF61B
UpTwrtPsLhfa67oOw7ljZKXHb3qVJTEAYSBKi8bihy2fyoggvzz1PfDZ2GNJquO31JMr8OJ8kPGk
DQGsGoom7mar325OPS9ohORC41p3dxWpwyY3mK4j48qxG3A3hO49qPOMBPvjb+Wd/W9DyLRmknz9
EPdh1CpHkbcxO2Y3Vbu92R9NR9TO54XjnpXFk0c29I7WMQ8NgHVt53ZlWrP4r/P5c2XawvToQrBx
C/o3mNSWzUahnprifH5sUh6vjU50eccpjfqA9+TZmL3+MP7LpqgKfUMtJCTugQtNd3/A63fUr81c
oJE2AtLRIBRa0B2XST+N5CjUHQmkwd2wdfZU+hhAJYfjKUgiawafj9bF0noqL7OEswIyeb/PwAne
LG1S2+dWDcBqoLADxSwnKN+/ExWnCSZbHZwuOhjgBOt5x01fQpxJBvDl9zSTir+J+a1YKf8ghLe/
pozPlzzc+KZxyUIf/5BXvO8Lw6sIM/d3FF+2QXsu1wDkEs1TTG9XZsQSHDuwbA2/64tv3cMCJ0Q8
hMwZpk0bEA0T6MgDN6NUj5FH10C2TXDwdeJoZuqJ8xtMd1r4pwE9irKvpq2wcLPrSr/gaINmmJFI
aUDvV+Vw3HNjU8PZY/9wnXBtyYwfS+SK7AANYaFHww/KPEZim3ZeB4BqkLpVj+sccBXVFh8b9VY3
fA/txwzIU0snvnZCi8Z+m11nFODjzqjnekwZXSxygvkpxBVM//tvh8CmUU7sWb/1KJPBp2GnWhhL
WA5UeF0KuHcuK9pPVHMMyK5qXhkFJkhNhV1OCastuMdc0aReKWbDWX10bDVUcp+Zew78gW7B4Hak
B7szQ8NdgayeDorWAaQlR55SY3icn6WPT24m9+HN7H4GGwu8ecly/TH551229SWGPMeRYJ8BA80k
VePve2bPeKJm+RX1zdhNqYLxXUMZ7UcIBAnhnmeRfaMGkw3kvcChSnW7xg0qaSgQ2scspk371ahp
AnzAGUhszyT7Mgv2wPjQs0loby7bTNEIT7jKk0rE4SHvp2ndaJNDZY6jr1hL1KK1SCy7J4RLbZTb
PH2XRvFhwGpL3UGBW1Dao6x+6I82T1/a2cuuisDVx0nxLtir6M/PDW2fU0jWMaST0yQUUF2RXauv
cHLeJCqF9caCrm3bo6E5PwUINduSIpnBPgjsOr+GIb7nLzH6y+cj9IctwBZrrLovDvivYwJUIBv0
IoRI7+LMWCPw3HApzSfiLB1LwdAN3Wf/6baEk3Z5MpRv9OZPaJbkavJ6pipLFLa4jMPmgb1R63vr
WL35fBf9pEkvAdHEd00ZSl2+MSIS1jizXjbftAGSidWwhaKgB0BeZTKKEw87h9x7zXjiAS3zFRwI
cbJ/mAQ7ge8edJJqHx8wEj4DwNYO9sEFnCyqZQp/YMjqeOSCnb6I6LHS4K9LS80f1Ppb5fSBfubq
mxu6Kk8+Z/yipLgjupOC/KZKZq6KVlsY+NFcTFOXOfghzbfc2ikA21SnRUr9kdzrbcWeQeVq/hZR
lFoeihZMJzw7JPo2tGOr/hq49mjtOgKeG0ibjDV6jLevmEc0Ivw+zryK23sDIIyVq210wxDa4XSu
JMY8PN85TpBNsz1zEpqkBdbqGcuO/cJQTqrW7wb+sXuqeEmbXfUbMpBFizYjBfFhti6NPuLpSROZ
cDP5Hut4JV4etNH9J/ETcpahfSm/4jXNlZ715JFGVyxNavGikQ3yTMqtE+SeaFeVmLPcA2mZhTR+
MoLJkIlZJxAB6SU/RqNIOfKDgC4hDhFcDIseS/ieuPs/04zrSNUzOvIPgZRc3DYlVuFcyxNcQPEi
mAKyHdKvzPEIfUXqRk1rCKjqPp/7oVEGtGM4huoVWCkX2W2tsW4dGv4dFWJnDQv5r23aU+2DfDNK
0PfYns8P8xG4IwXrxwJsyyV1T12wiLS+cr2dxVrJmZdkuMPXeRQd5PhKFfVFW886zT8LUmaK4YNB
RDvAutYdaewzJaCWd+ps4biCF5V5gmjppSIinDkTPA+4OFzsbiwTMxyflDvxmUZr/nLsWqqYGDEt
7lbR5I9R7aLwArVmdISJ6OGXhZ6cD9zObPHkqVJ8P8fNN5+P5LQYHa/X4DB13tsqa/cnk+cF0ZS8
1ftVRNmTsfxs6kDLqGlxAx2ZIMVzh5LwCLKPeEBjs0Jm4WRo0PvKL37UZwfQ1/J1qFvmIu+LwuYa
8GtITayD9h4+XvS9ojEaly3fy9Xn+FKaLno383YQPWaiqZwA69Gya8xzjqzHs1m3qbMGq0sWsL6Q
cc+lYz8e7FioTSsuznbALEZ1N8CQgePtohdRUqsNAAafYZGC5dKU2poYeS6MOf1NI3akKg1IKHDh
3dqjulqUWE8bihbatiDOsYNS4Ttik7eavdx5179vFutaf4OCDSV3+RgfvEr7zHGS+Ioaw6BqnVk9
lUS9LjPkq8dGjKtkEm3UrPLrK7S/OTctDfDK/Y0oxpymDZmp+dSKqSAvcpePVqgJ1NWgpYp3Uf3L
KluxlVs5ftCMUcMHBWY+CUPVFvJc6nJWYseAGqj+AJsKrxyt2UQCLRKa3gril2xImYf6n54ahVpb
0sDqnf/uhuw8akIhJns9GSJaNyUhFT8klxO11Te0LB9MRdDaK5t1ha8xZwDiIASJTSq6tR46FQWA
4OKUfZcWLfAq1WB0TULyAO3tyGPNDPrHOGsT3aJYQ4Axo0jTY4lmWrL8d9rGsPGdBVIbRt9lRz39
acOrd0mdv1jCxoR/5AJ5oUDBmumIADZE9Tp8QNZzyNNKfHxfZdoo5HtP/0BriFXFyw6QvXLmo4aj
xFXXwzRplU+zpMJ0jKSk4l6K4O8MnKRt4MjkROAmbDcDHIR3NaT6JiE9kNEL7BfHs0rKd4FH8Eng
xKSaiSUbpjxo5W/XM/icr3k6waXnJUboIIks/s8UtdY+izWAQPoVUXGBIonXO8K4rhp2zCZkGtoT
FmNL9Nv3SWZERaA1A801JWuP2CKBnA+0v6KYIPqBs6wJJBqcJx628Cff1HVKDkcE5thtAqHggAf7
jdVux5DDnTgwSPWxh6jVbgygMXqEGiyCjgHn1KLiYT7qc025hhLGwa1LDdzEKnOxT0+bF9Dif2cc
KnRT8qeF50ksc+MWkh1l4VFydXFw8CPOJg5V6oi7Eme021IYqXIshnZ7JEJtsQUVrnpmlinXog1z
TMQ+THvMuLipuSAhSZAJcq0j3Sg9IuWbU3ldEqKisasg4Hx3xxQFVIkbTZn/Wr8m25zPAXXPgtk5
3WTK8NvxPWeSwq3aw+ILjZ6efzd65K5zgkGt2BDHq2ATWQ1YdK/ohgA6ZbvDp+AZYzNhrV3/8+Kw
h5GAoLYAhYzb3oMQFuwdTzyeN7o2XlnS43OjdkIx5pUiQL663gNPB58YNUKJJAizsH7YnFeIBD9r
Kbgx1qJwUBO9T4FADZpQUiswcjLtJz3lYJ5lBaqX9kLCTM5oR+mBTcn6jHLaUBpvdWoiYJLZqLvG
4lQLm6KC+jDy95ED4tI552asA/XOhSLr+Ax8FH08PW6j53OOiFhbqR2pnOXGnSKCO1kz7YvucUtG
VIwaibMK7eJis7/w/VPS+UyNAQQ4W1kknAvDUxG6izxSUiyHRFpBzS4OE8YcTsaRy6Oj21fUmgx+
pW++Lvx0MnSspfAUtZDeLZan6Wv1qIscBbSqro/tOnir46rUEHzA0YcV6GomRi5EkDdd/Hb04kfu
mltYh7m8w1X3f/aut6Am3w3BW5p1dUhYog8sHNvoZSBcDtXAPHr3L2OyhKenyIcHKeDLo6Dho/Lm
Yb2vtgzWE+NtIV8w3cpa8YZu2D1c4gczmXMVIFF3pD2GWlg5FSpT74jH5zGlI6PoLJj9IsDzaH+B
4aFhbzVx29P6VW9uDRNOjV4rmnt2ax7EeZ5dNn7tnzrDXauxS/trQ5zGV/Vv1gz/wPYKpfW1WX9S
4N20Cx5fyDyiFgnL3JayoBonpCmkemGaKOPxXYFeBQnqVBPCChTvKbEAfJXNGxSL6Tf9FnGhleq+
FfqLcmivZ6A59HXrYoukmc4rot3vkoOAljuEMzw5VeHvMBXsQ9zBwTTgvE2tKuAqfYDiSbJuAX0T
ZflyiW4g+xJQYfnUpSVIe8JXpRjm+8GDiRDT9Km6dUPeAD272NpF+bZxGzvYpZd5wOWkNvN5Q6Zd
3tv3yrHiBhIcUwxkb+r9kk/BI+ZohNl9oQQw/1zm/vqt91yGiPoLzZTsIwPE7wSCSkDlWzO3jbr0
g+OPmhVYXXndV6uzzJ6PriciIaU76rnHXcyahDIhCHdhd0UzMG0Iq96mEtwEKM6emX/0kviOnMLZ
DdlOVy4GPrwrSKkVT7fSHnjyNxQJNy/kAsbh+2+pWGLpbwJszlpvLu8BsK8vNF7Pto6O90WtbYYy
FSaQQB2hpMvx3npfcaNbrBR4YHUw+Gv8TALT1JkV98++UozwMqCvY9Uh4wjYZ5hTodp1qHFHSngA
249ES8MlogwmfhuHVcYTGGdrA3oy0DkDiVKmFw+fkcP08ErxoDakPCh7w0Hi7zfU17+n2/7WYnaw
+rzApjVVTj5ndNQ0cTQ2/DktQvRh1ZE7AZZmXApa8mq7X/MHr+O9gP3jCSACBxs6tvEMgVq4eLRa
+n7YMHKEf7xRyzef/SImiL2vVWW0GTtL5uQiO8iawbIp64UvgEDp82Dd65zTmba2Qfk2yAYM/prO
YB+fDEQEWqKd6gLSpLkamdS9Vkspypt2PCcyDWIjroEOf6WQh84KXt+1BkAFR3J33bREPdF4Ag4j
ooTgQT+G1/U3/6QISi8j6dTcWcODmmFQjRVhieOEEDgBRBj//gM1ckM2SQfElh4HA/9RGq5Kiew+
a7hZrChrqA1J46Zai7/QrI3R85farHjQCIZEXrtbMNAi719ypNhlyGqk4j2R/OaHYeZiMyFtLkkL
L0yeqtdbJZ6iND3u7sb8kvNiPUZ2RVRSLyS3KLFIrFydxbBQXwgi05qUHt0s7uzqYO/gzOdudZkU
VZpcny3GQSk8yBPUzgU7JMYQdRQn2TD4WAgV3CpfB6yMh21flon8XK0pt4Xk5aenG/A22uKJmSkK
QHYs36TdgtASo1qpRUYCgiALP9/TYPWFOJPJyEQxiMNPqjhT/pnFc97uVU8AbxXamrRRutNTuqeT
48bnymfPocT1oi+S1aLZ96LT9twIzg3qHSx3maaD6SLLNdz058m+bY4rJydscMCRQimkDeWRkkEN
5xn9PHdnFK0EGayf+AuidH/coILVBT67sfW1in1kUwMy52+X0jGiwiqo76AtoGz+VaKb4rSlvEf+
BsMCkGGT/VbrEP2V+le+Kx6d2trTccA8EQhVOzXNN2sToEE0iO10lbtpRgbTyIGKyHyNuEBvP9XM
V45bkAW6YOomshtiKY9Z/GcAuCeJn2rdczHkstS1vb75fRJtGknH/q7ly/KhGP05dEU2tYuTYIEj
IfmWdHtIzS1WmVutYwe6VEu7d06vTpZxk6bosf0gYzrPgQHDtgBvW1rka4W8K/hZ3cT6sYKMgSwf
J2q7CQmmnHjuKEkAFlPJTAAwjklUvSnlJp6UK6GPMzPS9GMQz5PC8kVuGB9Hc4keZm6RNC3CyFoJ
4T212VWzBxdYn0DqvzSrpej8tqH/WB+NX7ZA0vZ7R8qwvsg8lgy43WarxQng9c2cJfZXa/1aLw+l
HjvOJOpZU6P7TsXxVJcGK4qQ/DijHpwRP3db+XbICS3Y7pRsQNuNVWIO5EkmqIt+6UoTokUFoO/g
/svkv8aD4HuhMGYhSWQDUrNH/5A53CWecnhgMx2zpNvPob05PTvjWGz2Z/RRADy3kaeSq7eh/dQ1
XUR0P4GB3XhiKva6z8xbl+UJbiWuYP/L1NXnQz+qZTngxfS7OnPT69v4Pn0uJCsjtx4gIsZ4zj9f
TNGvakAE8/krwKQNpc1t5XZEfLM8TBca8YqdZPbMABuJABrcx+oshQyXFmzSY83+8bp8f2UHpAAK
ZcYsTCU/a92ZeewEAjCFhkmBwtyijVRn+TAQUbS/W6WwFFclib+v5hQPPIeBOSWVgjM/UrUMh/h3
zcT1walWv1TUj3pPz9PPuptlLV4vrN/UuzRfVNGYwVoL5OiTdog14M0yOS9QdXxfZ2blzQom3PIb
IyLH/0k4nOHIl/HacTVCp6RYOrVjcCPuWt+ie5AuXFh6aG3CXBkYIIUYX7NhhxgzRjgiITBwQzfh
QXW0zuARmySgp1ahF+WxrVkg/qR4jBP2wn58PGRl5H14O9F8j+nimHSiz4ZjOYtmf4whUTafm7v3
R4XwghQ2WbjFuirlZXy2t168nKRezzFMO9z55R/8uij0oMGkdhUCNosXnTs1jC3JwjoQA/Pr7tol
yljSf3K2n+j/gpm65iKVWyDuFMc0p69q4V5inIvL1HNKyjQx7+vUOG/L/vKDK590wQyALYgTcWhi
7IJdLkNpftHipM0sUwsKDl6R7CwdswRDfSbaWcjr31mtqN0gsrlzmnpw348aB7p0tw4D43Sx/BpD
bOBNvxS5MUGlfojCDyJHfu1pNAEqqqoxJR6itaZ/mif4YruN4RsH4acuoNrFEy28NTAiFNhsBYcs
Rviuk+ZTTlCPyrTBTx1LXwIZ17VhGUV6I4mA4GupwWpCtwJP/f1azfZ16CuI2d7FigPMsb0LSyhe
NW7MLxFzvPBXznfV0v4NU3tZ9aEKIFQHBYisub/VuUmJhLQqYmdu7nkM9mU3K4zFNbuzElBM3+8F
x44uc58QLZBJOSvSi0oDbSf3siBiBloIY+AlGnPbCV45BapZCKlTIETQzbktt/lnX7hYqWY4FHf/
W/funNbAI6cZZ6CsEY1n+Y2X/B99ReRfjk6vWostDdvSCidua5c7r4JtlEXmeuVrE2gXe9tHMe1r
IrPgIpC1iEh9jxTxLIR9omYbFFmKCB/FBcPtPophCwx4sIEXq10QMY40R0Rtj1DaNevVZxR4KOkv
9YKM1KLBPC8krYWAdweUqusf1cS9UqK1Iv9okFCKAvqNjDdFmBpr7l3i+ng7zA4dQURL5rWSuKt1
V0b5G9YH5C30JT9iuFGSFMAmjA04aJJuX9v95j+DSau6yCiz0tiyhb5bfxqltrihCrMzshJnlAi+
yC/ctisL6fl1Ie4npeDmjn/vShuPRiNgeYjke3DTkBmRWkVioRSELTy5PAXeUc2Ha3FXY6fWJza4
pYEut6okcWL8alnOphS8J5LJwdRXsbVDdMN1qsAJbBFCgjriSL1gTFPxXFT0TTl99iVaGiQpwcCJ
fPsqBj2UNwkdT12ris8SBohKEtyzU9FUptl34PhOjm9JkiNpaULwUddAxdxjlYdirKj2i+W+cSc9
z1OurGx3fzsND+ySK7i37PjU6lviieLLkUCZ6Ba33Zi/ccBWJ1Ry2yzzhalyTKEu1ZhciveE49Vn
GnUMPraqQOMj5MUyr/3eELGFiWx6+AOjIsTax6f1q6GEt6Yd0hXcxJZnjftIArnb7EbfPW3Dr+PV
aSy1J0PFiZBWaKX5wemra6umXiGJOolxwq/wamuGkMCxu5Y/iyXJxJzHAtemGVSCdZKyJ2+OUp2a
SK51WsyMWWLleHom4lBMCwpoHP8GqXREP8IYwMTopMU+7AZgiSDX47t0A1Xj+U96rPvgEJd3UKlX
iwomxibdpLZIOX52IShItSp8UcP4FGKcldCuUqVXJeCvqMR/iMrqFyiAFXchdktwWp/l/UL8jFWr
dh/yphheJJB6nIbu0yx3HkkGIaNd3HE6kl4CMYZTPfKugulGzZzGZIrZwaNsvE37JfE5MpVl7+Sl
xck5CVGwRpKpQHWhmYIBvY6N4jjtL2TE50h41dAyA1LxvsxnXYd0w2Sv1GjjJgJzJXS7XPOAWKDi
sivUFFXMtjPS+J/lU17r7ZXhvYcM19ZWPHXEkd2UXGNdnyeYt+b7RwVWWdhUfGV0o9wcX1Y4jbIE
Z2vB4uWv39rsVKYw83mK+8PN7oPqNZOMDvgbh3wn0qGUCVBoA2vHh7XsLXpnWhfbZiFDJL8RQJnm
iS2ell1Dg9Etzj2r7FY/kwPgGIr1HRqAhDTb5QbUzPU/7a7iGmIkw1ewZnJgPH/LUi4LW4f4vcnh
9M7QYIpz21AfNTgXdzbkruzxqnd6DfmpyoY0vBbVKiTv+4uKeFNemlIG9y171yAjW/QMeUhzg19B
4SKkhNcolzywZjGUFaMZGxziwiWSDLZwBPIWAbGrHzB6GM46oXrPC1Dpe1I0BTV3t8XLS3qd01tG
ioAdUjgwNZWFo9OrNuNqsMatBH1SHez95cBb0+haSrO1g+iiZDp5D/SSorG1qdVUi/ZQB49EayWY
in5mINkq8djztZ0EBjfQtC1ftQ+jusRuP+nSC6qmz4zPUDiNM4SKepoA7JD56+fhoHrhDBkgmlAc
arG9EpBqGraweOVnFirpdfUkE5h9Jvr/1CP1ZSJ/JuFQkNrSSipPU5x6J9MHBVX60DnBkU3X1AsJ
ZlM1mgUMhxjC+tTWj9gxYJsMCo9YMSGEFO4+Njrwz6LCgilgr7CaGm+reOdjyZOFKlmf5/1X8Rtb
HTqxDpORD7fBYpLaGbRvN9QD/SuD1ZaY8az63SMvR+aZujHb/y9BooPsVWAKrOVflKp/c7HAGAoH
0OVwDuabtIjdjpfzu9dcdVsx//rRaNPeQ+TMo6eV+HVLaP9/EmLQjvpChVChI9Z5ahgn6hC+vpom
OBTw+k1+M8Tpm9NTTdp/jZe1HhRu7ZQaN549iHxfZRBMrfTaZGODABdCpzPARIjIM0QDrWfbVYbx
gxjEM1Hk2EEuUkGKTg9AsuwRjnsQUY4q95aaHyTuMikT2QKSndeO+XWzlR5O1LH8z0nKNTNPSBG8
AMENS9kndf0+6x7M14p6VkFaPsE2TNsoquOrlskddmFT3RhdSdvieqbdRP+NMX2zfAaSadZiN3Ce
zFgVsBLL6sBtN46Barl+OnY2g2plRU8Vki4clc9L4W2whydBpW4Tx05WAL4IoogdpFfjZh3/+20p
ekA6sX6bMpRfwMYMLFkg42CSMVbbpY3hghP7FhX6+DunElujPVvIfjSJJfQWPgsKphSosKK+heeS
aOW3DHCWo7YMeztJ9hAF5L0E7FuVZ/Xjp3qCt0cRm2znfgM8oM8hz5472n5nI0ik7ZI2OAR/rU6Y
4v1dVFRuRvvdxR6cLIkNOo8lqaq6+P9kc5cLcD3NdjscbqM3gC/raO6+ufXLJGS4cMXM2TXwIV7Y
MBzF2izIaaRvfrmSmaiwSdtnyFQAPvhrJsyM0VdDdKTNpYHtro4RdnuD7bRp54gd+v2UgVc9i8VL
OXjDog8I4nnJ2mKUJfzpW1D0WER9z6AmND6BfyaPd71jksaRDTJpr+UxuswkKkuKj9cyRbX08APE
gcEXmLO6bUmwvfw8k9U/cawrweLnze+iz3Oh3uDsrNDstYKVeamD3+W0MLZBw4jKr7mGeTIbsRRo
Od3bB9Z3rX78gavXR6g5+ZJ1nCR0lkfBO8wk0F1P6zCJNM8bEepgAhFushv8vXCDVLrepjGfUhY6
DKVahmFdjeMdMuMLeolpdPVskJWUEjUV6nHVS73of3qjFW13rZsC1C42LH+M3nA6bCVze4/ZkeAx
UTPU6Zb6G60VW5g5wFI8k3NiSbxGarrumTTspvJU2yX4TN/vOh8dWXGzWcjCI1ObhcOko8wHfmtD
GoOz+TItsR4kYoeAzI1G4eT4+u5h8V+qpjI3P9qx4ma/t9TOR/YXk5E1qSJk/X+yWToJgV23RmLD
WB4OHXNMmkF2jWVe7sCS5YoMx/rqqInU7YHDr/AYeipya8t95JHgxOkwIVEUwx8DixcQv6SJysxc
bFMk4dWiO8cFWV33WA+e0sUVon1c96WkTGIZFxqK6hgzdagVp0LGd1T45U5u3Z0Vyiv6I3BORRiy
f6oNJh4SXV/6awuwnHm0yEfWmyHxRn9SrHR8hTUUegdq4dOOczngd+qrSDeT6MjEnFLynbiiYN+1
P2sWnzjKAAMixzXMMtfnaBedqCoI40qd253mmycfibqGTQgUZnGYDel3HMID0wDVg0sT39n48bVc
YiuMuuV7EuoZz++tZdKYaLKdvQzurE7q8Eb5qCNnOJ98NvfDu4NlRt9CNBTLvOMAxfJWh/Hb1MIp
6xT/bw7pM7Mv2NSW3vyihScLQXXbZKpT+9BbeQ1WFiip9JxGQoBwNOZkL3zcilpdn6n4B7Kh167Z
MFkEKW/EWwEH22yKWlQC3pDDYuHLNISB7oq+LtSPQq5ieIF+/8JjbQCyqWaAFLEEuM4SHcRQEQ98
r4CDmwYkeqKC/QnqcwB4MVR25GcUm9/IlL+abBfGwzt8fzptHbZsAqGNuGCV/MtX/b+EmQZcfMCn
YVICSzULmXkSjvSMeDEebSKmYR+/CXJhUUyjuSpJaHpQ+xxa3NaMkA3Ez8gIt6n705EHBlcbFU8i
fZodtoETkBRhic0Gh6riQFKc9yJ9saxOcIRRnsrLRg5tYSDr/vimo+C9o102EPecNLSpevgQ8V6L
ig1jTjk4pAVKG3+G7JpFlunwldM9+1C3xNUEZPpVX3kK0y6MqS+7IhJ2U5cG+MB75kTiAMQVvEFq
13JFwOVXRin1/xUUZmY5Zd/wma0o6EXPnJna1+H6i1ZPvF+1l02tSRJEg6RoRwuaNGpQ+LhqZVSj
cIAQneYBE0zy/DUZsslGGBIO7UHyw/P32TIAxlOR6DIFOhUeTVCp6evo9G6gbtjx5tBmaDdgoe8W
FaMWMlCI+WSgcOHbr0297WFM0IoqctXHdRsQx+buUicLZYxxVrY/jknZ2/JkNlUZz7C6ZoypfMlk
4jcP7DxHxo95QMgtnYNbfL7Qv3rafett8XX85ZZ04FLJh+SX2j/tFM7RbT9rSijIvDkt1kZgKh+t
HrVpJMV8dBE6f+PrkWY09t2O5VY49t4Dzk9Ll+8Yo4AoMiSvv8LeCd/zKRBC7+6AAM5s+KhL9E1z
aGQuoJLZmrlVq6B/S66n9CPl9YxRaheHFpf/oHq0gyP1jE92e+rU6jsB6t7wUYwGhXA97zS5MWDd
ugz7rT9amNImxqiZ2WbwuiyVrvtZ6h0Zd9v9UnCWEngXI3Z27VqI5V7CRfo9wrXqGQupOZAuL0Kk
7TDutoFlPazPmLxP1hz3KPr1EhUt5J60ADOiEig5Rd5J8NkmtavZzhjcCEczqZJFcJuYb4ojlcBM
665l2djqzge52clKd/llJ12wFO3YaRnmIXCQnUXlN2DQ2+fKNnWk12g+3WKJ9h1dl5Vgl7z0Z3Jy
e/WyuEmtZYlQQfcVMncHxZ2vhqPuTHHyO8ffG8K72YwlytfWSiZNcR/UXHfMIjs3olDhe59ueBxw
Fr4clOyzRsIUEHubXweOMzJDdT4ONA8cXe1RBdnlJuIcV/tVZiEDqicthnTxo0xGuFd5nXnXqXIe
ca17BMzK7Vpq2/6ksrCjDeeMdtSa4Fmn67t8MtmW4hkA+lPlnpaNysVtqj8VYZ8RcYyHXZ4ctZfH
5tox4jmIjz0kcWHaFFpwV6P02np3y2Gcxo+KllSfvGnsGcoGmOUhl4Zyar2Z+yFP5bk3hCYSxCSq
UJmLKIrsQWqmoyY46d4sM2hlRNsxeTeoLpa3m2haF3LqFH6NRi9Y79Wv8rewp7V/iZq0KBteLNGM
LfAOfyWI2B/UF4yc7Ac/9ndhihUkouwbxKCBfGpsk5EH3vRHMqiQZmb9qoYPGOyZE2mAQkRKhanr
FfNvjFYSKRjmoyazbqCrQCzpni/by2kwilydjFcJaAQis6FmZK8PxK2MmWsswtj7TLIL6rXFaTTA
cef8mD2zkigW6B9M5Rf5NuUa/JeB91IuglL1j9EkiowzcOFzzYu8h1w/WY3TTwl6qBwU4OnIoirP
ck0dDswh8mStQEILkPAaV6s4GEQ5O314TvArYmFjBfBkLm6ybyt3tCqEXPp+eIL/3wGVAt7pRZgv
tP5ikOVdKs+o9l+ICVYWFDDW7CeejoVKmncP76IMIqGQDTw6zx9W88oFodi56VEJyX8gjfNnXbZ7
27wQv76EYDA9XXUmMaEwFh8VLRQzlQZCeNt5sirqq6lv21Z0i53IBdAWZAl5JBRF6Px7pO2Uqcc7
3ks+kcACqr2tzGp7OD5oQ8i1hEMOv5H1lrbw2XKu9DryxdGwUqB6+7qayamEf0R8Ge80Aj8KlOfO
BV9oNE54SS3AjyfX4gAxVAmIi0uyg3UuiUelf8D/2Am5Xxz9zN3TptR3LxWv9gKs3NJpgpnbCCTx
dLPSWXrM43z5uATEWsR1fG+od35wxcGbQI77g3KubwwZ/VhUhlQkkexrC2xIAp8iUZk18C9xqUmH
Q5+J/q7GNlIvuyQ5+oPhCEVO+6HpX0zrzEy/cGnYbxwRjOv0cZxEDJ/XWo9B3bl6Zh9YCnqN8zD9
AiXS1W22iVHOr3MBmsu0K9no7Q4/7dwFkRZ8Y4k1sP8BfSazq9m7YR3J6ITZR4uOK6MSmUe6MXrt
odnH5WTbdsRuUVB5fK304nc6en0KaoPvxMpT/181RR4TqJDZzP3un57cWzvuJ0bxbmedjP5SYB49
cw239LtAOGbPb95GxQF1YxZDBNxb7grENLIuI5zrS1vj2Cc6H4jgEU9uOw9Dz8sWeGfk0UcGfXuo
Qtc/UcMQEXNXX0xgziHLJmo0jkKKaGjGZ243irUEn5x9bXTP6Uko+5pD9heyZCP+k/JHgyYsS8w+
umsShrgwgis0k00+6WyvhjOSGBEvQuskLU0x/K8PxKTnTEDOGFyToij8Gi6J/jbg8/7+EjNejP83
t3IkhAf/68wluNwBFNaF50wfvqz8mhs2poCgPrjI2Z4+rzUCvZX8GoSSxlWCGwSkQYoOabyE3FyF
g/+77wDtb49cS5GEsvFbGdkmNUyg+IjCs2fsHM70UTKikEw/xoSRiVUkfYOspN2TP16AI+9HK/Vh
LrBcoL2Vp5zSP6w0kjY3WpqMh4IrrHoECOiCJ/aykb6UmbKYw3wIl+k/X4bDcwCqvBoJOCPuNo3r
IsERwB53MeNsZpqYkxIDQH7q/EAZjlEVIVzvPNoqNuCYUUIFp9LP7UVunlmZr693SYMYNQ50DLf6
GcZgAqOIo9STSTYZ6HBkI6L9isDFc9K00Ch3SbCIRaL7bhdAv2pASAQGujozs/Pb/r/q4ZfeKsst
VYw6t/4WKyEk+LLzJLP2Hr3EXFPEMw7/6e/7OZQdKiPtmzqbHPUaVuo/VaFpduSbAygF2y5Mbwae
X/TRWFXnf3LPmjzvlKZ/HaqAMViRTkIUKwaocHeltE6usLsNj1q2s+4JUM6OwUIjhGHxUryFm49u
2oHhN1NO1IqahJTah3xM28ok+4arFygPFr8y5j3VKXgSJvaY6lyzkrBY98ASSU+BAorVzfGicGEn
iivoDjhlILmuhHOcfX6M9VXYXvvAJeN3BsKo7gTWtY/vOdpBj/bKkQhOSOhezviOk47YTmw3QbuT
SmzcH1+E7HPGJbnJmKKtNLSdTlP9p9ZcliDV8zOPaRI4be0EPKdTWEYpO57xYdKzZZWD2eN6C4SG
b65qw4JoJ6LsCyngYYZpgkC0kIZ2wdckewCE5PEY3BSWapUVUoHUn/um2Hn5w0SWqsQFUbQRBL4m
plF2VJGd0AMLu/UcVX/zihiBNUfpDlujAW6+0euBCR5wS8ZFEut/95A+xD2cD1f/KqoXmeozgdZW
0G57UVZv7LmLBlM+OMv3Z9bih/GommOU7Va3neyL8W89iU6IygWoNFeM3EXnFJGrnB11I8aEEqOZ
XIFefM2yRtGw+Km+umNf0LaVM7d1ZsnSO5pfl1QhwcMDZFRm4vQNg+i3ncA+i7TXCy9gSdLT+7Tv
RbETiwKLM+p3UasW1OjkX5u2JSnU5I3zxtmZ55dnDfOjTg70+E1ancc3kJpHt+f7ZjLMmhXLRL9B
QKQI1GyyqW52F3aQl4hz05g2teCKLK4pzypsNKGqTdfyJ07mpl+HsJiaUnT7AKugVGQBOa+7snZs
0sPX5Oe1p8HFRIHF9CJvvHz5XY7Pu0KwjKHfBsY9mzQugi1Eas2ZARAeCi6s1ThUVXNpfQlxNQ0a
6egtZFvN/i5QfNrXFazfXnu/qgk+fW26TXJdBKXTABkC3hrN4YtP+WUcWAobknB+++yCl9Owu8tJ
GHgap9G/GVgTkTAt/fQpcHRFI/c4yLXkW6n0vVchU/kJA4g5njSbOowQ0KOLo3tfEPr3joNGmrjZ
rjTdTPU38T2oQZddVajar0kqBPMpjZLMO5cncDAsGvtSGvbrH9i8++iP1rtPROloZEF/WeuiA7e2
Wa0PqltO4XO0Gs8HnwIIzmCvszC/guJkcQ4rGRRFPMnruqKbR76NdQIP7OcaQh5kXW/YPXKASr+i
45SsoyNMdTP7IWY/O010QgduiFH+uUcOEtr5Hcpi9l3BWxccNXYNjfX+/yBHZIWHBx3RqH2bU4df
KT2u0KVnoA/ApKjSG2cMCdfu68bRlSMHARRhgg8p6PX17Ub4k9wgvCon45W2CCV7qEoaBiuA+581
W36yM4/sRuZctkp54+v4BQomEnk98o2JuP9MbYzmr4OEqTJkP2NIoNtYQ/rQ8OiMNg6cw7ULB5V7
+yG5w06N+oCyclrRmXn79OPVWw3g+ZFVHVALnh6Iovbbm50pEiOzur3DlIs8YmP2LdEzgt0x/m3j
oVP/GFcNpKD1t4bl+ib/wzwq8UGeMn/zSuMxQGYTWFM9qWCUCBVuTLOrOK7E2D3cKVW8eTSujggG
TLyHalf66M2J4jgeANhGbgoto7ipYXsVzCTtgRtXl5Zbswmim30QmF6oWSvhdErITAMAITd1+7Vt
E0uszyKSfrfh3c9ieoK/0W4ugOMmIgtRrliG+unPyk8F+SEgK6awAWnpBTgTxjhdokxZzYsjLexR
2zGJIj03aTGM5YYhS8v5yV3bdLjsRMdO6STu7+o1TNe8VoW68JY5BysmrcZKtnlhbiJgyQsGHElu
y8V20kULEJYvEozid3raPJdyqhqssOrDlhqzVe0yfKCILFt9Uxp59cNtt9Nn0w/wL8sIB+UDQixC
JOQ93LrP43fWh1xeYrlZdthJJKB3BcgYe9gdHn94sT/KXYgzxQ3b87UQWZhOtMBNkEXZPkJpMl/0
BIt7DuMx0U8iZfzwDbHWRdoszkatl9+m8UmJjJffOWhM1iXeWIStF22img0UXHhkNASkXlz1ASVm
K8ZUXhXD3J9ifnv+GfcuYJPISvmu/LvH8bkpdDP7XitZ352Uc3bYCIvQMYgNd9EBMmvCL17eTcPM
WEZVhe0/Oy7WD3Lmnn7E58EnlIag2Sz/SI9AgIHHRVg4ZkzyD9fH16udW9jgAfOzKXXvxTM0gBMv
eTL7OWoNcP8HeH8KFjkL+bYY/M057yInXjLfELSAtyOvNTt5gjwAzobQrl5n1+Dt8Sr5DImkV369
J01LrQl/JCIxFGCuyd19EwdWxI6Z46PWBBpKC9y2BBTUvcPVKvZcNZlqXD6W3wm9X9PLCRNNovHp
JtjAPEESvF2spP2RZZtcjoUn7Iv8bPNu8WnMM6s7pY/KUU1X3VFMW6NrNoVbtsoAYO+fFD+g4sRs
OjsMZzxsWuNnF7txNRT/s0e4R/2dOjOAIPcDMa8KmGAy+oNXuotoFbkS6co1RtNUVjm+Ym9VQOiH
Mck3nIgs2bjSkevbS/UVIyV7c6lpDXDuDtkm/5V6LvGzSqyBlAXvlHPWrvb3sevYgRgMb2jz3nhR
9+OZCOhvWhVSZ4dKhfPW0BMIfWBKHHtCJmkNsKLIS/Z3FGfqPyJmdRgY5/CAZcVAKxnE9g+mdkSa
T+M9jEAkCkXf8PO3ODc3mlMnLpJk15g+NCfTjyUoasnHUR6bTdv0BTBGQONXV4V6QD1WBEKeGLsa
DHSAXvbIGt4qVCBL1zNe/H5HPxDGl4tI+//yCWLeibJfnN7mTAMRgMXAYH0oDldJjCbFwGs4Utn6
cSH10D+D+f5n/YINS6cbWLfgu5BuehHMm3dxcnbGZcXg3VfSSBj/iZyvGuFZ6Ot7X1qKoaIGh7kB
fe/HVUqh9ozEMXxB0zrZCf8Zsvx3vreh3AG9q8xIRKJFvEKmPmbzkEHhYFMPevZ/Q6OPzP279Ir8
K+0PxhSXrMK4OsUF5Jq8gF41NO/xed5n2IaLLwl4NRLhB7uRfJj6x82LS8iG6k56VAXCgPeoEcbB
AfSRs1ueBFGWjGX+jig+i1TTEC+/ZVEFwzrQC+8GYysRKraz07JFeGNZrPNMD3QWLQx4oz3YqYoe
25EOuxalz9k8zU/DhwWGc8HFogSjWBnYk/h+j4c7wg7asuIqYnZVDXvHKfE9Hgwcb+Kka6vT7MNU
cxVmwlSx5mj+Jbl02FKlGmrOp436g/1LP7HmJCtNTBSGwjDv9bvaaepViZn2+o4pi4cRClTBULFh
OaiYSj1k37hwyVxqAE+6IWRN+Hf4ewG5eF587LOBW/55MMxEfNIKzBEcAdnH5Fgb7z7XTS1hRBeO
wghxG0MwWwKgWKLhZ7bRfbcyNiTAmkprPP6glJjIflqGEoP6y5/oBJ63sO1t9urkjBiZ2J2cwRjU
DARABT+PCpO/qRZYEH0Rk752oaCkuNBvaQj+wHhf7d1jiNTtPMN9gTcHrf9NvAje7L94a+3No5IB
g4PjGyCPmiPuoR3kUq0ERHpvvBZXzLQQRMUiUcZZD4PpYbmSg4vJ3g98uhjmryc4QL2cgGHyU/iM
DiD/JPsoNO2RVnDs/kRHONbHOG4NSDxIIy8RQRmJH2d9/ZiqdV1ktAjJgGqcHkZpZ6VhWSoidZIg
PPf++IF83PN8kyKnoiKwlWsSdb6qNdlgOmgNndpW1XYvGnttoJwZZ3EyDFTTyUIvZQSky3bXhVGy
5Kbu1N2HYjUg0bJpro7XGevlkKQfYpeuTB/MO3TnJKnRKASxUxy7VrL7z61wMqJd6isvbnGhrPrN
q/fBTAsiqDMktqQVcD8617b4YQMg7XO+ICOdIjDiRfG2B6q8kj1UMjcozquCvtnoU3wqgHvdRodd
60rEQgBjJK0J6jOkMkaPdNYz4Hxy+Dq5803ix5Q/dMQOtMMe93J7YYk3PFmiSETPKTShBEHgS7SF
apcBNSyuDTajyOgVNKwnkHhchEF+Bnaqj0dBbaMXjUxGpg+h0cWK2zs426h4dbPmHRryEi2ksyp1
iigKfnW6PvbwWfL9m9NxermmH+hfrDKj3xva7nZcZaDYwIt9Zi2JtzS0CV3V/gwkD5evbnz4B5Kw
tPWnBXXULB2GayXYFgem7tkT1EYi84lhDRss1YYEXT/cY5TbVM62rtanvnguZ2BF99+FkPZTXlkW
E9C4UBQAu1APbOsiN+KhQLxYaYoyb418I8KhotnUy6Ia4haR+Vb+xJDe7/F4zL1VTT4eKqNVVy70
eWO+5Azx/UhsOGx+tJok/NFvVuVu0yrW/Q8TEAdNW/JzPnf4cZs0Nkorpr1BKkf2gkoEtRHVFkg8
DsNh9uLu8kv+mk+ZWzrm4+qC+XX+Gdm5aXeZRJ/85XfuIji93De8sLJoQC0O8AOUTf4E3RGuGzbU
d59EcOMiwxN6gHFeVSAjaJVO65zGl4X66eD+Hpm5gHn8xmDIyqeWFlA1znN8o9FZmJirYi/znx46
vbvlHFpj9rV8adM71w2TuUxgznmCL8B2SmqPmh3vhElCOCk+xKqOpsWmueQYxdx0wRYNMP4E6wy6
wdBaSzE61/MeTKsJMpkLTBBlIR626PKgn2mnWWSL8EOdAMkPeXndiWOPDhPQzLBwhnMu/dFA7FOU
zd3VZwYHli7YyFigrCnI58pxDCuOPsbchlU1om6EwnLdFnUW6eEyf3wiLr3zzPNiBVjObjOEsJ1t
wagQMSjE6PtN9uDOnFMbfNZqysOnutVg6p2my7DValwdiHJG3FUCWVUp7NqBrfodP1ibx9pDFScp
D4yvbv4hKpFpdh2WwTO1TIsxdxS4X0tzmQ3rU48E7zlthPJ3jzC4MMBVOLpbj4VeBPYrp5Ln1tyD
s6NYebqk3Xl4U2FMjdW3vTCkEVbHLsZ925dirHCEKTdYEWdKSJyn09902t/dNlWddCi7NhEtyx0h
oeMneYwvLUNu6KpaNXcaiVZebQocaELzA4AD52e4khsSHj4w97qyWTez3X5D9RA3VmH5SzKKr1LW
codgeF9wX1CFNTL1lOgDKBU6gBVKbfizZg+hdKdWiAiYPr8kqU8exviyxmpEFjsZGAliboc+B07S
JJu8a8ROD0E/fAbMq/e/59Rpn/qpCpI0p1NBWfP5ehhQZ4l6jG/oUGtzIA6Y4ekeq8VTTs/nx4Te
p3nHGxriYrKCUTPlHcsRkg1ti6LYV+L/OnBhZK6pYe7013zhIzjVRvUG1D7bv/QtGiKXOuPsOUFA
yGXJr5imQ3K39UlwflHmKGphFJcZl12D606aJH0Uh2khf04ycI2ABZj9JogfWtXqPzfQkSQX2GN+
EZRNfjmXc3VrAoh9jQ7N5xGJm6SApPzfhHOT+1u2j3PT8TMoG8pDlSsGFUUbjuyBsYThnbVrNvU9
43xiwm6BObmYTSfxaceVDAQyhhJkfZqHxzziJu8zSaIXxlwLaVo0+4p8g5secDdkliIfVbch2QBC
4YSmhfqj3PaOMFtlgCtYo8OkzbUBLAJY389C3OA+yf/rd/grtYVzVmDnHK8I4VdbNfpF3jJh2Vy3
nTgt0nBXn8iQeen2G0H0TrH3rINSOxOdz1gKFEr1Urhlqr2b1S8P1XJcW0osBp+E/UA2AH5xfx+8
q21ZEWX1kk2VTydDjlY+FMTFiJOF4CTq1gZLvIq+ehdC6d60EnNWnO8CrY1wS1DzGg/0zM8GO98d
CqcJjQD5Loolir3HHDIgQjyaQWy+MP/dYo1ezk0mTrkxiUlDuuUNBOp8NyxKo/rLk02kCv5i+m86
OMuaeUBytCukgkEXFf7y6BI2lFh0ZRMFOsNXDJZYJG5kakS2b00gvq9Oh/a91iJTaljkXiVzVXKl
uQtu0ybaEmWXzDXlBTyS7o9/cZcTi7bdQDZHYR0ilLf1/w5n9jIdVrMurBzwcHD2pev81ixS7dM1
+DVudSVKIPncNyt+GVrORtSOZ6UZ6EuBdtVW45YR9h+fNDoOCerN+EdIem2L6+6ZA8EJMLoRJyZC
r+WVTsIFFq0btnSl8XMmF976b7obobIrITQAXHXfVK1HL4ra9xROrMWvhb1ibnjs1+9Zmv51vK5R
CrCDPRgkMHjgwyrep1ZB7CAIA+9JPfLB1WXcEY70IhMdN3yCg11nOwRfMwj3i72r5v7NQ6W9HA+i
R8GGdMK6uv2mhmE2qEqJW/67H36SWhPHWFLwXZJynH7Aca0+JcDWPNtoLxMyiEKkxegsbdExVVNr
ZhnDhjkRlmfPxp2YGQILgCpZMgpKIg6OKxkJRNfV/o5JNiLMi9jkzGdL7oY44xEfIWo9Apo2FXVF
RD6SMlslDxsjpllycMPKfvLvkWp97G3Ajpk8ux3nxvas2or5PU21Vi9WAczTWx64rcmFYgO/9WmY
veKf3BadF1TwPQI64+AYzr3t7gxjSFS455gTUVfgqRAZ8nM54robcG9meDEKAZrKulMA0l2kwpKE
DkVgv75YHyzjxQbw9QkQeFjECtABrQIVeaz/V/pUOEXUHdUWaYg2PfsjfYXmSUHwLFuCsRYQnVJZ
ELBQwZ1Ys35bVPuW5ZwwxOzLEB5zpdej9Pf7StpED8XloerN4mgL+rvw5pvjH1Bb1OLTVjSKuuo2
8w7EaezdVOsyJzmCrfuCpCBvpmOyHOf+h/ZnLys+4KldrVF3YKjGl6Q/4f0Nkp0ZqmopNz8Swjvk
8h7SRksALt/5Jhw8EfPGIqLHLEZpMNXNF90yhfh/nhP1rr9I2unB+A40n1EaSQHpa7B8/XfhTMaa
7scIMYZ9W5Lh+FIlb6G8ag7uzZfSrHBxUpXE4HwY1zEyViY9P1x/gqVXtzKZQh1uj0Gp3EqFqjnh
OxOaEpUE+bt3TyONvTSMM/xdyWA3G7ijTic/ySS4r1/nN9U6K1/8zFMu0dbI/Ggd6MUlF3iTsYKH
UsDlveHswNVrVyXJYnp2bCDtewz9sr7W/3Efd04UJch1KbD7TEW8qrHYddrN+8NM2/xB8Ewy6vxP
uRGAmT/OEOyvvuVWgfUxYaSFskqbPoNkg0x+Khk6VRNwHbOFpBbF/OSATtXgmi6J+A/trIn1Wdtx
RZul9Wmou4ADTLLPSV2npQt7N3Q1gx3dKDE3YnAY7NfJm0+ceR5HKu2gKC6foktTWMhDe/mzsltW
pOZgreIy3QSiV4RGLZmw22wXn8M7u6+bcj2Ia3OG6FMVGwEAg7nAoLx8VP/c+kAIfTNZOtoLrWAs
B19fDHDtkOLIX6TLuqy7fsL0xjg+6YSByQGIpvNDHwBS5TU/OkrHg6cAgovpIn1RO7pg7jbyMaId
jsq4h/Ww0+cVDrwKs2VvA6NTLrSuB3HIVLwKS7KK2CNvRHCaiT77sSUbOTqYRtYkwl47dFBO2Ou7
VuV5YYKLNtDNpikq7fsdpYKzZd4OkJked0JMjpLgO/T1aAOo58KKD6O2nCifvWklvvpun6IHVyVU
mU9yJOtSTUMekzlmDWqS1ulEdKKJNjwoUwZD7hoUjkjkJ2rqEIZYiXxuc1TedJEJSMh5GHFbt8Bi
FSlWCCUUqQEqDr5jm/uQNmseEgpKPZDA6M9MhrX0ior41x0fZL/KvqxYVHHQ2VRuDMTiA8g4LvHG
F7UBQu4u+sLB7e6BI/IkZoNtG1YknycCAmz0P4J1ALlCfwFtQEQxwy0c0IL8otYWRQrErQohhADT
lXYWqwvBkuKWQGlhXNbeIKyxckTh3pthNhWL8EZF5T83bygj5JDqt137tbfAFmAo1VfEvUK3O3ZG
rxVFkriztq6XB4W0UDaErc29oyk/0W+vvKuyVoh2T5FRLucDSB5SnZ6WqKguGAluU0dAuFxVIb1U
5qMg696+ejzfo8CQeMAvLnFoUIFWcuHa2VlCY2CFWQkP9GM2MsZ4rHcwkTu4O1Vl5aMFBob8kr//
SN6Oh8FVrJZdh7Mu8XN5RDW3fSpr4DjPri4Y7/TCnj56xMb8tKmgwchDMexMfxTJ29/Cq6QAJwDg
D9qVYsfqwWVJsqHQyEnsI/+9ocYo1DT++nkBMt5hOkk8Y9TjgV8pBl4hYdW53o1dXbpQiMw3Gboy
Qa7DOmL84n/bI+OjMbsLo5EQ0/oHWTIAna8hB/QGd3BE3lYDIW9SPutDT9QAydZCI0OoqPrXN3nf
CqfsCvWEpsSl4w2Y5bN7WVlVw4b7vfC+aWZTqmAtY7UVabHhOQQ2FXkm6OA7n14bI+yw20uVHgJ8
G1cshQTbCQ7ml78GKq8itMos/hdW96LrJu/Bdb3FGUaRK+WARPHlWqS26f3UF5qHAq+De8mmrmc6
K+gZZp+Au00Vr+0OKY+ja+DXIkSpUw0a/FAiEn+/VjNGZs9Eu1zm4nMJPHrbO6WvrOQKzRsZDsaS
zeBo8VpXGWZwglBVS89xFN0l8FPVAuyj/pXk9iZrtLkG00gBTsHbFMw9tYevDmDu+/ffw3HAK8TK
MkRkuzPa+65Wwiw5NWGXvZPVctZz3xmMzrtke3hs7f7sn35U7KqSwuiHse0avxo4kB6HroO6YlhX
5JBhyjm7rlSLvAkSnpvbjof7CRIvRepqec43j2q0aRUGeIAqq0zqeevB7YRJm4Suhe7OcUrnPfsc
x0b6TH+sssXPmsdadFm1i/7XG57eHopWpTUXqqRTauuUYK6S5uWpyRj+VtRZ8GR0yK5pSdCa1ig4
DcrYosuL9WCP/LvhFkZfe2dmYXTMbSEg9puKI0wuTkkg7nemCRrdL4azE2OWdLpe56RsYn9068Eo
U751DVo9KJdRK9FkmlFhGSdyX5okTcZSRvjwHj4Iz7XF7KVnKzNWkNl5VsGd74DBlDDnkY4orTMr
GWzzGDnszUuSLCcBwGODQE2ArNRVJpxQ2UtnNkjkQCntkq9uEA27eNyr8dEMcopTtKr4NnaT4tB7
gZFAKLY9NUi6bhOSPf9f+XsvyOSIeyI1nBAXO4ElioHs094i+gn7EPCacR/bnP+J9MI3wOLtwfEv
j+7+644S0SsfrXA2jHVXt62r+Fm+ERXDbaeF0fGXKUk4zZFo24Grka4RIHokGwmRV/wDwIq34oxa
hq+sZI0NLjTuDaZ5ZpuwAgF/ORiK33IHfexqhtrQmXBPJRZNWmvq+hxlyvrZuCq4K6UU30/ih8Vf
fIMyqxUoBfZsKisagWMtYXF3lUDSQCmMjtlISORY4CakeigX7PrrDQUCtV9J8kurEIK+3HgJJIiG
rsNvlfR095NtMgW8imSkzc3Q9syAodiEbYOQczPCXluPRr3IpSvSLWrlbVMAbqhA3NJMV4IKi5zZ
uJsM1cBbKsqR5RPn5rinJmN1rOaqNdaLHPB1npRjjUjWhAawIe8s8FXfa+eS2GNNlZhK7AuMXudI
+ud7mmZxzZ/EB4oPXb4XS3U44G2Ogpp6/VDa9+5TTuhttZ65Dl7ot2kWD6lNwzK29rtPgy7pMF+O
+9UpomlaHnWp/md3RdyQU7Upq67sqIHj3gaYVWXiXUDtSxaV6kWzus9bgRjRz+Pv0MAZFBkppH5e
bAcmLOM1xYrDQYoFqaWRoXgeOujd/oZY0p8/tjDtu3iKIdnUclMfmH2ySb/PWwTX+Zt53OQDNfnU
SRMwm2Lyn+XMd5ro4buOlAZE7CZzaN+va+AFX02msE46jn08zhsyfi4daQfew7KRal3Pxram3Wd/
7n3Hc0ziruTnpNeExPs2frPVhcYgibillFECUy+HHoYY58qV2XFG3AIyZK+ps8rFOD6uR11sn4fT
AViqwZ/HwWfnI8sj28U8LPZbq3O67HCdVl7GmDz2wKXkYaaI1tmP4BFqxamx0T7xYPcbUs6wiUaJ
uZ2oNoqlVCSkTv5VGv5HEKbrTVuCzafKmXDpX+i3+Ijc90lkn82Gqu1SnSSxqETYE9rSAvWssByC
YFN/TueGtXRgWIVV5kwyLb+A6AmxFFYcI9tQLGtOIOz1yxxocb7tQOmR1H/S6d/0ghtRZ+QtKT9S
XQsAD1EVU3TIfhYsvRlN5a1r4q+IZVead2VjhCKilU+PU7fTO8lIEIhsLFa/4MvLy5nYxcClxYl8
dBOeTQcW79mSLXTbDhH8pLdhYuCmJlcK6IRDshl6ht+1uBvrLetbM8MrE8fb8VrAgtfqxdAwKg4c
JMaG5b1OjZztu8HEuf+1jcXEAGWNTNXQRDHzrSHD5RPn726h5QmbxvGW3dy/FwXBRn5lJOX9HMlg
elgE/WJtimPnYrZRJbgNlWR3pU2AYsPkU6zM/2nIcow5BjRTLwN4ehWoVN+zA8jfQ8bfn2OEB2iO
i49LTaxa+jiF3mMcGgmcKaCqrwqcIngB3R9cH9YVr9g5ESZnu4WRdIKw+GTOlFYPyOd1Ie2B6O4L
x0xhVLAlKgfW2X4AyHglilQdcfYs6le153q6PuTXWhuFzO18Zcp4Z/DfCMIPKUEv/sXpf21EF07+
ukFRPyWX1lCOowb0Wqxiyz08+fa+Jznkr7oC0ZzTneAabmhTRH7AuTkYACfgkmJrjB+dfQOH1hE1
p5ah4j9YMipiATW7GD1CmiLek69baKetWBBIs2djjg9WH+MKytXi0wTfjSdtMswsqw9mMimDKeph
sBX67RBwOlD4HzBdaf/cKUe2iEoPBEjZzKjdGz98WosyYypOsVtY6ZCPS3/gogR0NEyzgqm6jpPz
3P1ud0J1Rex0rAX2S22v7a4Qx7RKFzfI8zsHiVgVF2tSzfu2aXjdNKGhoRgYShz7zYo/ZgVKkQl6
5bcBPjM8SkPlqfE+QBnNqPWNwZj65q7sRiJPIssn6aw+GiUuZQhOEvxlcrx6vMA3BdmMi5jjNvRZ
asgX7sBRnhNM+uAjo5V2NX5cvMlGDBS8I/4fG3qCPswee0v9o5OzEgUW9JTlbgnp9o6SRMeERWdK
nZJHTNQTiQ3EvbSGELEJ/H2eiBEAUQjEYhMz80Iwt5L3njHv4jnK6lbTo/y/6i8MjahAqVd86lnX
JrZrmDwCVmLfs3+rowrULNXpcPiHG9MitEMMYJTHysyydQmxq4L4TfGgPyxHvuLujkPFYeB0elWo
sU9BJ7EESMbxf+O5UhEeRtQ3nLxw5PYvTgo3wuM9qYzd+1Vbk9dkvHKg8t/e0bq1Ck0jCvPVeS9f
damU2v6EKli+DmSGP5j0gginzf/kNLSOhhGVg/qPaY0aOdIfJdyJVMMVXbjyWHp/QZKsaLCwbs9D
mG55B8WJBf1sxXcujDFR2MXs0d0sjV5LPLK6kJo4cQ8ZsIwdrynBsc4EDiL9kLFVWrrMopRvd+zM
jgvSjSj0MS/FMPSpPZzgTBixKZUkJQ366fW54jOeoeScBo6QZCZjBizDZ92YMMmqeT/ZXX7ZTNBH
j9cN5zZUJ0WP78+YKVNDOf7OImYdkwOKkLBRcsIFrI5kxyd0uCMRlj01sCrZanmwgcVVOM/hIGdY
HreYdexsLI/NeBUTCHQPyLRbZX0ynoa1Dm7ncCcOsoNAFookjixcrAfQp0iiRVKs9g9fs+ku7Urn
6akwAUOmBrTYWmDsX3eOpS3kzixKFKKwRvHfI+5yce9jk/aRCJcSs9Xj5g7xQ077W1nADTX9XGis
5e4FiWDz2ChUYHCX522isEcYntX8mSNcsDy3Ux77DeMoL97wdhufab0bBuiBDXCMQ3xkPrW77kOl
hkXSOIHsy5EnQTRK0xg5IDtTHDQjE0CZhrP0bifE9OQIvo6a0W3oahNNfxRxzkB0LuPD1u79BIf4
gdac9vyBh3BNhRcxpjVpVlGBEqe1KNzRNu+Qsdhj7DcNzDj/iAN/iZU6EkIuroseHfUp8J2rtCbk
YEAlyKz10gHjmTmPXbOIlZN11yCXD+lRn6TD82Kh2sINOpLHd6/fftuYH5YxAZ5KIRHFmhE1sYxp
VIdvACxsI96k3SdKfiubLd9x7ILzq6Y094xGEv2yUiCNkhmhUkZ6fQy413ZzeZoEFBTkGDyA1PkQ
yV9qvZb0DFYGIQzOs1LpT9g4KkulcuSUvKrqfRIBikxg1OyRCt/ojjMPSKhkR5DAyziRrlmUrZ50
3HBuGMoJtlgsss5xTa/CTYj0lqm+oiTgjWJfEPwVkr7sx6/z0Dk3imCo4D6gIhtiG3KWSotYregK
nwDqUldryp9PDRZfONppT7axKIi7KT6MavnrxpCL2kTOweq7bEytin3eycwyF2G04hvDC2V2Tobo
1QGwnmWqU/LujMvpEtVB3KejLWe3/p9FYad3SsAquxDYTxocn7MGyZmadB0jMut+1RYJC2f8VKGT
t9SU8lJzytHXoOzI/J4581GAT0R9sr0MKEY/zbIKwey+pC8sCMcZb33MRU0D32uNZxJopbHM0w/k
cPwhd4kBINRHHDPtYUEVFIJ02ajJLU1sdpzOubuvW2S5iVf8JoKxrEQh0yPKzWNhCqLqcz5q2IuC
iNPWrdayJWpo2COqwB6NepBC3qLVTz1b9XdWhFjOxu4eGuGwcSboNIRufsd9nt+xlOayOl8xKv8X
3tY3jbQeN2cH6pFHAHfxdDOvflWHY4n0kPfrDUjDu6XGoIzpsmQ8gJyyGp5mln+x1mcGU8vPwDYj
AbMAouduhIWnO+vmr7O0J8tC5UZIVb0wpi9GhssAnQXJjg+onro4ZSQD3cVHQp69t5V9IM4UUBV5
ouQK3D4HqBEOhwqvVALKS5HAueaMYLtGAobCjQesmGXyPYJpWmm3rxEEh7NA7Dta7lU9IPVrqSug
n9J7ClkHQgVZuHJWOAcC71fJ8sbOt3wE561oabsYU6yYc8BnH03cKaGyxOtzQTM4B4Ju61Di2L0l
5AARHDZGQG84aSOLfEBhxPhonKImQurwo18m3OtTMsS1CXzKeOpj3WrCu3Oprx++bDtFoYK1ZRps
pGcFEU9IPJEfPanNRRjDB56eLDpag2ZkmdKy8Dm1aqTUU5vAFi+0ahIvXkN50MnOgw8rG0KoG21u
xkx8YSU3pB7YQb8FXPGR8KrBAa1cdkvyZkE79qxtu3GhsW8CANvEcFyjFKBvsebTA+r/w4xH0BoW
ea0M9FhZqcI0FNOztFdJwvCeyeWJCXs3GzvzlcglhW0e0vlG8Cfy6f7BsRecvdAFncvuPgOjvV2C
yXZVumyautFIK9rVrvOOq+3jQV12jCe6Sh0K58WJfHhCiS/uLiiAZ5RP4z1SKy4/2Bj/oBcGqyQ1
O0JaJzAEbGbYs1900Xm+TGHAvAEbas+xVUeiRsjgvqYAl2Brw+rMuTvoeBuXIQhY8P8a+Lx5rx47
7o66Oa0o9imCEChlTEKzxRu3+XLcpyq+nkZe8PaRd3CKEHljWlL0i5XfjPStqy4qYkccyMCyR/sC
HStKB7Ivic5vbtu9955dIB/aeIlDcn2WoLjHwr+s9DGHHTwojaontN0CFFuILIzz1ELBHkk/IWk5
TL2lyXKat4ltsd7kps1f6Htaav0Ve/KId7SrM4CN9bSbhMF34wYCUqb8X8nXHrK62RdamzuDYJwy
SpoOC5KLAFbF94evt+5fvf/ARnZN71prRkSaf+UxrmZ7cPVCc6wu11CnjXtqLj7+6CaZEMfQ1T+1
vKoF6sdftWq/UFkHW1HFA+A8Td67QAZf8IpNmkn8RgC64joqiE3DRGADIfPdmL2jEBpmzMVQbVdZ
CkwWnCBPSqs+3zLG+zq7SU5dWJ4IaL1EcICu1syfytEhlCl5DKdGD1S42KqjiukFU/VzaxF+qG3c
sv8hBeMom88lIX07hlEL2vbTa+gGtJhgdHoUs6ZL5nbY8YA0B8O+IB59STor1wJs+knaWdWAhm7w
ukbkPetv9aWVue7Opa6LJiB3A5FxtIqj/APKHYTJ//xnLv1LjLm0iN7A4jPo8kcvRZN4Oj+b0MRk
+NipSW4RZywhuWWxzC3Py9O6WoVC5JJP5Y8axV7fwX3JBTqMohD5FkP8yzFTXyoelawb8ZPxot9n
wzX79qT1LpkJm1GnQf80ZgU79mkZdv+Vt6tBUYMZjvqOhhAvBkX7mURXg/1Blmm22czasDuhdRtE
Wjdp1oeayRj37v9qh7Tj2F+EbfOBMbgbZq0JJM6TXhV+Pi2NpzPvZkf3VyFJxNnH9NDSZB8XWL4C
d3xaieH9dglIt9PBfcIxR65Mv99FuFAcM5DB8WyQ9JWSnoiy9LvFNt+aJ8OjNYxtdVL91bPz9nN9
MNbQeYpvDTFiYkUtEghh0EQZaujHUdwGc0wgovlPek4aTugGpZ9oten9UPA3qR3rxeEwR0fyTdM2
TUBOUoAYSVN1E9+1e0TuQZi5VAB7CPv3DV2r4TAU4xVDbmIZ837DN0xNzGBlHvEm7lioEKRdiU/P
EMaLcWnD1tkcgTuOAtUA/LMiW+jxok5JNEziLC2JM6cmq9u2F0tdSXY8cF3WAFdLqQogQ/jyE3Bm
ydB1ZiTbidU9RICYphkPUDxNtyRkzLwCpVnw7Ka+TWHGgN73sy/kFlgh35sop7wjgYYaU0XsnUPM
8wQZLHa77Jb8AXZJU6hhhF5JkdygTuiYeffpC4VAFCI1Tk8L5Pfo/Gg7GVuVmeyd8WNqMwKVGnHW
UjAi9CEMwtwv2KYrgt3a+Eux5XxOzWgzd88zWA7uZf2CeBUzzj6eVzbEwdi/F5q/mFnz+nyyBbhd
qhl9oRYj6S/ObVZxn4w2jdXyTUwGoNMIW2rRJrbjHsfWFOtIO73CM/hyTLCDspL7FSw+ZDxWBcrM
A20aMEP8/UspzM8o3nPscoikRYCbcpunCyuXf6+dmyF5BHphWsNKtigIi3jH8SWkYO8H7J4p6fgU
W3E1y8K1LuN9w2Abpb4O7W74GAPRVZpauDgNgUlSUTJs25IiZL0xgnB1D7YCaF2jjZG5WtWfFhm6
s5oeuNt2+O496gP7r+5kfTS74pDj2xDbF8Prh0B6r3/wUNex1qbmt7QPC61gPdsWaKu0dnMWmalo
5LHGSkWEcA+KKJWbcFtSm2UPTgph3xO/Q5pnw1QKN7g6yG2ddX22OZ0isngeKzjNvSERBvGAkCuL
HbkGPf371iFyyzy6YRo2ZKebQI57b/mhvv5qq3FmVK7AnMn9803rwv8eSFL/Dxs2F8lHkMsOeCR7
uyldoLFbAWr9yTd58IU6QGnQHZ9wUZknhQ+p2sDWrf0WMoDGxjdEPw0XbuRVFYvNpsgiqefPh/Sy
cbUN7sTMeSP6Vsa+yeXh3+ZbRMvdikHG8y1Xbdi7p6S0HENzvR9jxhSKA3sDzQMPdNDUKvTNLRvF
5aoBCDcwtO7YPmnnTZ1bfAAaGBJC0Na0wnM9uXptHBrkv2VBOn/8TXtrnl2lDyEPfPDoRo7wHocJ
zeI3N2ZCFmxjMIRBZ5wfajRjSvWrumnjuYHytjTX+vEsFeqM2W5PD7YApeRmb3pUZCHHawFNerOf
0HF57qEdFR1qVImgV1LkR6yMwYv8hQBOrncigBynM3knGVIy++VatGcUQJ/nLCaqjUihZrNwHPoR
V7p4dvt1vHmUG3z8bEhxh0lEuOiL9e7lgBi1uD/0MScVQ4JFf+GhiE07YbvirSH6HJoVSfrPdPJ8
Z7PuWDGC0SWtRndsIAv+Vnt/VLEX8hSMOLBEpmfUjg+ezrjg/ZPG4vv2YMlWf4vvMaBV/rezAiRJ
gJw/udfvwEz3CqEYQsF7CfA1wABEhpUXTz8nUrJmXHCAvnwtYeZU4Ibsbv3zxj5kFRbq6Vc7/7Zr
n8Te/V9RkBHHTd6lGWG5+lW9JNFZ8tn/GK4biyeqR1EH/Pf8spy68/iFtoq9cLOnmz+yr/UWdzHx
OGZzRWi9rqYuaMZXyUaJ6K3s7ShI5M9fPAjA+oJgwQgG0uC3H7d9P3MawwYNbCqVSzuvrDDBdTr8
dAKmmdnAhXbQB71vdPf7K/1/X19MFZX1VZu9vMYlB3AzCiktxz1NFW1G3jBXDFdv9Zpzihr56Vpk
Ok61CQmzuMPWoBc9oyvV8zU/Swo9LhtYXf43abj8QW4Rac2AWuVAB7Xzsd2ry7xGFC4BuIlcjj/9
7AOpF/0iubzCTMf71VdZSVUlSJ7GcG2OjKkpmH7jTELG6cUZXsasqLdeXNFvMbre6BTjEzsSiUoi
9IRIhFq82u0/xtZuyGGkMZdnmQBm5r0PG9fiKZLdtSwsS4MBTFAyWM+6ARvUQk32qLOb1wowTv6g
HlIAa4I9gxda8YaZvhgPwblw5M8wAB5bGaRf88LLz83fQvmFWC3pY1aT6HvfhOrpVS8qhKkZ3ny2
N6bKuHLN46KXkYKoUtX8JO4yumks+pzBRJ4c28FMxm0zG9j4tHTArFfww/57z2P5yO5CZBBBpC89
kutq++QqRd9izYAVDmUVfchDsus9J6sjjlPusvMh/fIRKiAmbcwKoSUHLn/S8Ew3gB+IvIHaopjK
YUu76miwschTnKF6/dK7lJrgWcYFd1Ki1fNeIbn3MeUnaFB/VlzX2m++160Q/afQrHX0L048k1PU
ovmf6HO32JA83jQRXV3+oCxuUUm+R89QOLWz2A7mg6N7uf9I+BVCGn1VoFEJz+qYlJqmNhOkof3e
xWIoheUDVRDuDsYJ1+gnr3umMrAOlhfA44AQ1YoazONiUcy9zQBqBqbezpGCjs6P7U8fweGP+J3d
OfA3KrYbB/dUMLWHN708qNnak6mmA6ImMTNvMJ+FdvpZzSFhKY8ldMy6JLJR3XEcheT8capb7fsE
FvMZi0Xjvc3P1k7x3iCdXS6obp+pV/+8JjBwX482nra18aOIaa4k0Yxs85MFmmE9+ClQETLoHgoE
+duzBjvZqQ3ugCvSiQQ7SqaV3NT0Au53/x+7vRyE5RIvGCPOMrHf5bEKLNSRptNMcHz3UV4zhyAV
lRH5jFPtEpckyFnn765ZLV1mlRtzBtcT1yaIE/O9m802hdwlc7eBgfMriIUCad008yCjGFNPkwV1
tusvLBLjSDLJiS7cvYB1A1wo2WIpLyUmqKbwrz+/lbksKjfloGECOH2uL0+Mv8hZ9DWVu4G2x9F/
BGFo2a5OYzi22MTd5qxkrI662ZIterMBo5XmZghRwc6A39S1URSV6qvd3YyA5o7JsD3lLqyHMYRn
Ks5EiZLDOP4dOHfsA2RKKCo3FMltVoTNguY/+ofxgNgrAVsatgZLwtgjPGtrQeLiV1KW2PUbcdne
ws7nRZJKNA9DEdjO/hwdw0VZumqYVnK8MXRbbGjircEm+2J/c7eO8a9UoQkmOS9+dnA17JHbWzB1
iaQAZdlTPG3xGCoUiPbffeCRi7uMjYS2X/pTFz4CE4cqYCs6wQ4nPLEQdXS+HkVDnlA6WAObkGiJ
SOTmX60TEqK1jTu0hBS/eWISJhmqne+E3fn0vn8rlJjdgAKtFhtvYFlabXz7wuQTImOmYz5547mi
OIHlwyKH0fKaYyUXWMq3PjxhskTNTO+NQxuLlQddU7Wc3V0kbAJYBnDR7E39pToMI4FGKdi8Xmcc
yqQB79s+60Z/7zY0vr7sQ1TndGRCcMbi/Y5acLN0SdkAEGCnI+redtf0wPI0iaez/sg02XEh/Inc
O+9XyJDkTNeIOThtgRoCEn8dyBUAOKhTJbX5Zr717RP2hKUUrFU7qqbeVg3ULTF11iTPVY4hQjOY
6oWF1TVYtBBQDDcDT06ZDUBDg9k4vIkaRuEXH906Z1AfFmIdkLFZ0K7h+jt/hVWgypH8Jie5amPn
jOgHGUbLOcKLPSjk+4QhekOd2g9kFlgPdzmF12ALIeSIwCxZctBU0qkvF1hQUI6s79d8PnIX5/DS
RS6kJA0p9TiQReUhUNhYfyX6H0EGNVGGrno7lOLHkKxRkxonYPFggBR0a4fkuevhrpyuZormS2nZ
vpuvG43F4YNA+1zG1aTWy31OEJTQRs/bW3HI7nV13FN6yvGz+eZ73h5UX+B5TE6A7db2AcieKCcx
4QhRsK2aYhilSDUYjsZ6+fSG3pvS0ke1H9DCPwt3lRhiezbovPsWwJOVpEXbB8bsln/b9xu66tH6
sMvvHkE/RxaNG01Or0eNQXxRO93sVDu1MD25cTsL9/hEIjyUvfEDjSnyTobp13DAXoVpoDiRIB0W
D4gDVUBEYQBzOdt0wA2SjYKQjZk4TSPDLbPKQUxTH+sDpsnHBq6QUMH2h0AcZAN6/b4/4kPBhYB6
MUKD+JxJfDpwCU7yFBkCmx9mJknQ60uot7Q7aJETmB+TPzA9I/jTMANew9fCC0cQJOTXun6kyluY
62Hp7P/zAoaS8K6MY5U3fG3ypMAYq/ABHqFpceso/kRuTT/7ssPrH0tnL/U7oBm6AQeOFO3Mbx7k
k89C3UIBeV9X1q9yEq/gmS00iJOLfPHW3KQ2q5coz+yUBgUAUvlhtXVa0mcZAi3TWIbeHESLsV+v
7TL0MkganaRrVjBZMZi999wi/Wvvq0u4OoUSQnGKXJRe1kTZdmofs9mrqosfXHXUf8TS0aImgXBg
aVVvay+3JvWjWfi1tYRL34J6Kvehv31tQNFLB4ebEGbUnVbCrqyl2yjDxFt1YrVCTuJPIf9+sCVo
DhGA9JCqJF2Jrm9K1mdita5w69CTtJZiSjlva6yUmYn8EYNgIgCkbvyH8kdUzjzni59kDggekUM1
obLf95DOWxQluRX8IpfDubAHCRZ321uWuaGmDcLpUT/zaVJ9EEfl0ibT1ytSzccrtyL5WM9rNa/P
w4VL942Z4zq4cqR1si5BFhFFUEDLInWIfzaoskLHtEVsmZ4HNBBgUcf4NCp0Brs35sui6kfYxuPL
qvWZS8g0GMV2UTXxo2wsREhySMW2lNDDct4+WzcKUSvjM1U8k33TO/xvu/RRzYsBpMrNtye83rsH
rurMO8rTA0rPX+25tFMxt89sOYcz1sXftkHWzAlSFgGVSvMVemrZ8x/9a5htr15ZJOgzv49OTo9I
cb6fJ0BL3FpxV+zkJa5h/yoa4Dt3qiIGBn5MZFRiR2OeR59nLvoXebKdNsFyw+mVzPuXTUickuv4
fQwLvYDYONbdX2pVEwXCUlgZWbH67lShlDAT0oFjx8roOt4xFT+Z5p7QvbHM0hyKSS0LfOaqa5lW
L1OELfNyZIw7mrULynL+2paDm4nmX5VorNWhkiX9ZfYrNo0DqWT2mlJnD3Y/qlsqvfaIYn1emGVS
LLyLqKKe809Dtz9phbdxPg/HwHCN+owB9154agl62WnJsja6Or2i/sVxHlRqC8nBkYbl5NaRYNKV
rwYJjX+1bwvEiTMf/wXgnf5wQI3vqdI6oYuC4MGFRMlh3795JgvBN/Xnie5+duuq4+f0jQpefY6u
sLmoEZ9Da4W5NS9eL+zpoOu1317Mj7hOdCG6fijsKAUnHcrMWY1gVwImUc286HxK9Gr9FRs5BZSc
jHyeRzL26DDU9KeUfXEaMdgyTXiDrlthkeKJctoRRPQ8CUUcG4IItroFK9NO1dS9BUgCo9gOYqS4
svOQ+ZdRtnj+V+j4mBmB9eQeQsqWG7xy1W4Xu9B2ePckat4tPO5c/zOIQ7IlyT6L9aOFbMMf9FsF
isCeKJXDVReDMKOJUBX0xzGlOaz9UA+WTAmnZYwgXOaG0Z7N3VqQPZozsIJs9IgFvCJ6H/2rUXI0
sV4Hunbha4t4OkQgrPN2KSvnTWvJ3odbpdOKXtmfw2EhnFhj9kl5K4I+X+12TKstHbXYBSmoACrn
Jb1VX37YiolXiwROJNcVuG9UOB9yNrK5dOC4mzVCRLfyHiw5X37ssjBitfRT9T6wLkznkMW3HW+T
V640Hn8NHhf8V96YMURKm33L1FLGOYzLyP0I4AfxBwxVuXL9ZkiwhYYlMY/YsaZ/e1SdoknPWneG
0ptVAXzpJMjICmJF4EcHjbKPErxkA6dJq8/lhNn0sMNt2LUTIIWRVWVxYLGGJAwOdRVnpMJR0Wl9
AbiDtaIA8CmHWnFgIuUq39XpV79KGFaCF6jgWa1tU1sR5Zchulxw9ifuFbUkgUT4n25xmyTPQ9Jx
NU43CT/0jWobrCSQV9Mw25TtEFowrZa1r04pL9uQIY7I6V3z9ioUHqbAyNN6s989XDJqxwZiRdlP
Bd/w8pdI7lI4Bx0Ecyj/ZBO2NPZPSYovxU4unvXRlsDMtPgnHsooz6cvEOJGoxJwuuKrU5lmY/ng
rewT32gwOCZ1t6rBEHcUHRhyX37eTRjhVhGjTO0CNU3lmPGx0xYymYJn7qDaRgJzvX2x7UgjnUxd
vG2EL20FvBazdA6DyCBU7z15M6dbH/MevR5wV0V+4U6ZOPOR531YvpbKsbq5BfAPq2AtQd7jIBbO
t9+wLEYCiJVKKcIdyvq/P8yAHbi0yryPvHKIfGa1ZbY85Oap/aIKKomOmGik6xtVXYI7LMN+2YiG
4MxzuGvlvdbEKMwzuoJRsCf3EzUDxGlCLRkeTDns2uOrsdfDQG1KX7m0tgN7di6cE92K6DXu5+cV
Qo13le4XtA0gMLi2D9B/QpO2m6UQpjJ1MAGI4aKe0DqdS5tOZqib16MynFmcdDpnlEsAh0ao8Yx8
UVV6OyKZQM4h7gquvci6pj53Cv5D9rmhKDotEwEkfgZ71MCyA0UYeQGQx75mIU59hw/4kmXmAJea
KECJtSeG4lwrlKPR+eCFsEjU3kvZN4dCWDfqJCUPajtus36D793kJmK6ugqwYGW+RDbT/esW8RYH
jbN7KbFD569nlNtos1z3sxKRDJcqxbL6dfe16i/Sefn86TWWJR8NNlUyKd88kOQ7lsCWnw+z9A1Z
FKURRuwnL15mOFdyLJfXsteCyX2fuEMxAeINWSZmCb3Q6wJ+YMHoSMFDYJ9q50XfLi7EMtW4P/lL
h1lyJhHjiSfnNkl9ztMJMQHkz76uGKxL1jX2DaqBprTsAARdCmQAJtDAsTKyHKdxKTOXmoQF/ZH8
5i7wY1Zi3meh52kBqWJsvYIAA9rn0tk53/FYicvuf5rpqww1OBV0Vi9+YrkNNMdB5e9hQvHVaISX
a9J7uP0Fp5gSXuYVQIjeaYViZlpa7Yzur5UNEFwGUaWCgiDy08lRc5JdriRJuHE0NGjc9XMqj/yt
XSD168uIkMA1xy2cYmrVFosClLkaUm5+jJmxJrvX1toMXHzj+quSNAdswdzWeO0ehCPnKmoURL3q
0uziInIFK0tkhrFztF1EdigDkvLhzFCMmb0BzKeXEjOpHbd/5kNwFMx/ghv4PRjs7nNUmwMduwik
ApzlNiySVawtk3ZX9/97FoTfK4joY46EmhyeB5vNg4GEFPyqONxkWP/4Fl97lbHm3BgNXMFbVCyX
AvsopXPNUG+VoboyggY8QBA1TTg6sMGZyuOEdx5Io8lnq0+iuJ7g8gxAaPg7V7nQ94ugfqCg0s34
Z0ry2DtGuOuY1ZpovKb9l3JPwe5I1XDDsbcO3wctDh52IaUoO2Hjt9Ene4qF+IE2mD+WPZawcD2H
wV3sCrksSq2lDJ4SXLgfYmdpr2oVuWp0Sqij03lNcwv6XQUjNV5Sk4UlTPgRZnqwnT61nn+8GaZu
d8GA02rPFDZVM/I4wmApug/je9yqRPtk9olqwIxc21lEWJy2nrwHrW/vfQwDEuut7chgsSTIqAie
G9dEPkxQwWUD+cn/7JClKOvNcPx/6VVUCCqPJ7dDsl1X+mvpRQo52a3XxdhH+DNXDdFHSxyxFevb
hE/xSpoZIQYYKAxtC6CehQ17JsDX+cqtsVYeLyBWhow8A5iUAJMMbNbvafGK05hxWe9Wg9zIqpkw
klDLm0tIP9WDnT6ls2Gg424l+LJihzahIGZB4nO8zvJyHCBybX3aYiYIKtbxF36P/bsVyLU8xga6
1PGnz5N5u7K9aDiB1yUsOAbeIGWnuvYhvu/ehIwJ70bJNWpvUrfUcuVF/XDiPUBKJF4ekA63Eovt
MmAqUvb3IyKrDelEu6OmiaFtw21KKIg6NVSiVl7H49P+5TsYVzeB0/z2eIzzVim2SDrGUjB04z7E
Hj5vNSn9bs/18krfiM/YligCQtP26XApFJ0a43HP2Jjyu2VD2LbcZuDur0L7eBw8FeIZG13/gits
y+hxKdHUBu2K3eGp70SqIfyqiVmwJwB1hsFIOYocCTUp2UcvVbG/ueEYQYuh8SfJpJeY+PDBrBs8
bZFAdovVa3B8nvBYJ43psxKxSLeNUT1mGZVVdfhzTlFzILlXqRc0AwWo5jECwo8Nr8Yy3JENc7tE
IuVt0webeBXCVwi/qUilwhF0o/8+L7tv9GKH9CDafQlhgahye7lQrWTQtoNLInzf+OFlfeqqr9x6
3/VbR27MF/iSzsGNFFTB8Yk+2AzQs9lI5founIN440aM7+bSjpnzCEi0ufhwVgnvQVEMd5SibPbu
PVECRXbUkbiqC11tjJ63wZmWS1F9cyK2opp7Wu/IvkiZ3Dv1Et/gI4/Wr6hgkPzIf6jty5yrVd6T
jwmvGLUNjqZuWcdLVuwuow3ZocVvwZJ04I/2vgRLo30zR1zzFY+UNNFqRKDl7pckXk0SnchZaczM
SSzmbui/aNKG5jK5SuM5wJs/5GglxUsWHIUE6hzI5Ibm1b8Jr/1kCcpCqr+s2zCyD4akGgBh8+ag
H0Hy8IeDlS05Ar/2yV7IFOvgkfuxU/ykiWFiqF0He7AyR9c+rOqEaIr69vuR3t60DhfqLrUUMTKG
mWTCChKKZKwA5fiFFnqjFsq1yTuj3f5jPB6F/xELiZiVv8vDOeY862XrTUI1Defh+F+4rKp/WYKY
+pa/gIaucube6BWh+2LQGMJpI+u4Ywv/RcdnMMxDUq0Lw8Sg4LmUfqnTnwV+Y4i6GlY5FjQCiSyD
8rrAhbvRQa7EuAs/59z19z5E1y7RlaPUZs5+PrAOS+cSm3L2wNKakQod0yLjT1TVGPeBb9tgsUYe
FmY6B3qCB75ZlJwk8VjRHcoJUAcQr/dNR3qVjYL2GaBygDZvWZbG2mfLzsQcmytviFxhRbycLl2q
0kq39+Tzl1fxStmdI5EhgHzEY5mf68xRs2YnUqQeO2yqRXBMJzqdNlRaIoX2kmfiQC5DpeSZTUnj
BpVzh2FI0ZrBMX5VhdOFp2/tkvzp8rl+df2HnUwiY6LGAnal+Gn0lyDNPrmQM4ajTdqPA3l70EKM
uPxfNf+T/3Gb5vvX36zp0E+BoFjGlEJLo6EIdd0M76Uq6+gAcMUHBkIs/p4lDjqZupwzCgL/FWRm
18lN92zmqBJZI+1Lzn6ExszWZ7X1GxsPA0VDg5GnYhKQFhQ5h5QC6OeuuJHTZ3JO+G58liXP2ulX
vEFdEl3voa68xTg4PE6AcanCK4jxHDDQJnZYyjpjvk0Rs9PUp6hLD6wzU5ao2v5KopywtgpHmL2x
VthPoNCed7rAaK3ji0LMx0i1pvU51EFsCBgHEhJJ/2T3F6DrqcmJJneuf4zrR6QQQhFbCrYEGbTK
f130H6KphbUJpS/CjSCTCOcEbAgzUzJPdnrTG6zzUzW58eYCgpvs43TttNTZ87NWElvpQPqnY+DO
2ONmJ5/TTcwdHKnvR8kpPFFUKaUBrnntkh+deRUdO0XvFhAB7HOrR5eCAoVREnsKkGZrIm1ZkU2W
weoz75PqqX1PFrtQkZhsKzPD2GStYj5HMdRf9Pp7A80UnZ4P5X1OVygfUK3jtQXWZPg9Ch3rAkPj
6VtcjxA2vonDDIgm/U2HX0O0+fEaHWZ5BlTUF+l/aAHt9ijPKFB9MhpxONa16iOfWMnqTk39CFWP
wpu93SbbxRoZ8YMlc5z0keTcWPeNor+uq7JeDkNGnJzhlgLaMfrScK3UYqbYTTURVS4XEQs2575D
PPLQOa2D8MAdfYg3AlzmEmI9aNO5DmCj7D+g5/DyB9vnlIKASuxnR/InX3ZBPszTBUBS2IBXuMBL
/qAfVjCpnxIkAAQ0VyzPJ0FeBm48mCSPR5JGzJOyiKffHYt3RxVYlTZNpnXI/TwV9q5bX+jyIswo
IsznEj3W6R+c3NogZ4lTiSIYawTDwXqkMIFLxZc/c8GhvZw6RddhNkWnzS2MwGiGilA2JsqjxRPt
uqubRLzENeg13nVdCN1yUDKbefO+HqyWokeUhEd5KxXU1YKZyRMj929PxQycykqszeJp1y2PFf03
WIT+Yu3Q9nOLUwwPh2TEJxFO57A28OS6w8Z8mnQJXbiYkqXGIpXloNDLLBevTkXiMb8WP08fxe+E
h0XdHRXGP7mTFPUlCnDCLyq/N8sFpOWaWDvjEzYbnr3F+RtmRnaZ+XJpUHzg8AGfcsGHFZZvkvLH
9M1NcnIXhm6VX0ZFHdH8qZvbQfIVg4zgAzao8SICz8hKAOS7twxPSG1NDXxAt84B9wsn7HeZm/pH
H6SXhdXLTjIT+is9R1yQZK5gWjuUYAaxXfNMrVuVb56K8w4/evdzUmo7UHg5PEGAuEBnHkIN4pWO
ha6Ojwmhsr42hziQjWV2OutdTf+LwnzO5TIe8+JfiXEX6SeG/c+5jLaxy9MIUj5AQgNgNXU+en2l
hAvLXJz46iLu2tc1zYOkP+M1djJvTyWp7zTgOutRXMeM6eNWYuL59Xmo/NMjZlWGKewt4474D1sS
kosntrPL/YQckR47QCU/4eGEKPV0MdSyqb6SoG7NH0zhhgo+FM71te7OL2VRrg8c/d1t60njWtpX
V8mOxnvf1CZYVEZsLj423v4m1RXIUMgnFy3QaFJxiY2ooQPmK22VNfXvEymr/+QVSRH76sNNnmw8
upXWc85tGVrvDkfK9t5B78RPQuIKQJU9ht8qCGsF/cLcJ+s/Av++020dcsuRo0Ca5HjC5Aclo12T
KNyNwL0UB3TrNB1S5lJFLeO78nxc3w4SqhOUVn8wqwPLTfDpB7C7kyNTQv/n6pR9CswVwKX+tGxx
09TysaG91Ad8xh66KHJR2sj+IJbGO2w1JllDg/fmXpP5CIIiYlgvUbrfJXBPkIJ+yqIk56XHrvTO
1C6Ed+7XnVxwhD+OFrExbMp7FBMcpUSiPwmlfjIuNCyrWUSE+HCRjO3zIQggDxNQDi3NizS0z/CF
oRnsTNVhqH6lIitsMd0/U88qm0IHg573mWsXKyYbNFYG5ieOaW8NNSnR9BSkVE3uTQqSR1XC/eYm
qm7x1ylcliRTlmy7QIjCKVSJF46fOG30NN1bBWr+VpudB4DZMAZ1JiYpjwhUI/DWhP/m0pBOGwh+
Zgq6hnndZ/TIC1JbezeA/qp89JrNpgBFsiciPtClaOAezeN/P1Lmw+W4yZxKmkudWO5mPhNbgCO3
x6MkWVM/kBAESlBJvYtMZC4UuG1hb1agKqZt7pfqEx5GMdCZPUux0RcT03TwZ7at0XfR9PnyZGoP
3YQ8wDgztQA0zH9gFx8cZjivYYHMsYbv9UrGPzNRmnbZFuJI1Z2Y1Xn/fVF/rhRax7bFryXRh0cF
ckCMvCiwFtW3jsTzZ5q+j3Rxb4TisDUKz4EJtYuO6oY3yr+4t6Yei6PsjTLMsD/5Bc4CWX8RpvcS
UcwCDAQEpu5kkddMWw10z0j7UGf/LSE1LlH9dKc3wlnOzyH6wQo1FUNiZ6cKWDMQiqxf3xTggtft
BOfhRRgCWVR/Xv4pIzyFnzm1ySU/3UVLmvVn8e2Wv4ql2Wq4B4fCF0aDW84/KLA+WdGqKDHMLa2Q
5jVk7CouQlcCQ9SpqGbk445f6F19xJe2p2NvaGcJiQ4b1pEkSuG/dLtz3zxq/52miukPnRQp4rcE
A0mNzKo52+uSpeIA46yu+oK2a3Hz8ZJ5K33py/bMGOGAaRvEpGrruenuGOH3mFzUDFJDmkee92Vl
RsSF6YTbH9wjN7hyGmarIAHknUptqcwnORMHAWr/mMvWGjrkkM+pZZ9RAR0iWKNVIb6ARRhPMsgI
TtjAtivUzQOJbZtg/E6rAeCLtrCmM/ScX66RWukxEC5oN9quOZEQTsDWAbtg0DPEBm3098lXI2Ml
X5NyQI5Zi7P1ZI0QDRma6l+CWXRAv8DCQRIXxeB1tNPJcA1Ao2N8Wgl7dHEln3YU3zaL7O8MP+BU
d22IG5hfa9PyCnwDFaraFs3S1kowvtvB6phblcaxJ41wq50B1dz7V5sooDpPcXIvlWm/abYK+4In
whJnfMd0KVk2Q/8hu8IQ+OiUptC5l8uzCxWU762uS7kijyMnqg1HC3+aaWfIZRZdhxPk6PAC0s7l
P0gmNhVpmxPuSdmyVjB7sxWowe5mzBqRw5fF6S22VQCXyekX34ZCq0EzLXfXWnPXM+KetH+fIb8+
enZXr4zzBOqug54L6+j9UYM1aQUUm/2bxgQ6dUE6BoZcX0BsT5vUV2FgC3LxIHTV5ecDA0xvWmrj
qHSLIimWknrKyk/sZSYGyMJxg6LVbj9BLYYbaksM4iaaq4mOWUW8h67EJVohGdNXAaLQKtHHLb3v
UgFWh6Ng2zbgLDdAuJGYZh8E2ju2QSweyqUW5Uoq+NnogwbrjxtYgPJ1lAqvuSwbKSONgn2RiMcs
8iJjArrRVH6XZPGJS2xhuRLDHy7SqkZvpF8ITBLuLHjhUHVGw3tWHsWQ2JP/yyP5FtiIjtvUZRRa
ltOGyALjJpvOI8g4JJQDBUB6AKj9ejr7RPKMvs2BPc3VOb+LGwfaXt6MXGCQBednRoCmYYwnyMJB
7R0thsWyyybdILWw4zBDqFXLyNGqAxQ69Eorp1uD0ZJQ8Xwuk6C84dKQncDhRiqAdqpIUq5XFBj4
dk/MMs8mmCqjFxXDTf5viiIb6oQo4MD9VAM27yQdoL2PtVyQvS8u/QPdDTh0I9H/4s6n/RXRxiDH
I4vv+CM2SK6w3H9y8Zw4vOWOVFIWMMrHRCIwU3Y+AOrWX1n0WWYZOm0M5EfshCki1hZULGBa81/B
s1Y3+pU8UZEjffBCFfRZ//xqNESJuPt+rGIurSXmeVpY8sh+WcdzVuXEr1IqSF29AlLmvOwvQQhk
FxwsEZvCqgm38KsFJAJYfXyOeu4Nh3p48EL9KGqrIzopX/YTTDFG84/UANgY413kqbA+8mNCdda4
NHMBB+JzvjaBJtzwROHsD2q4ubnjMwafHLbhXMatjs2DMqR3z8qNGHK3PRDbAzp1qqmdXl52Ii2F
/Kk5kNsvsi0sSlG0xGmpTbD3qAcaxb+ImMhkdIoKJmeRFOdkR4gMN8wnqDrO96nfEHtrKgfJpvQw
LqsllaZHATPe6M2ACsczn/L3kroD4pFcGVQkMubzsHcTSbGflnwWwzWUXKh1byyNaOh39mamY1+r
ZWnQUy80T+SPXpwcBcxpQ8zZT8CpEstBBwm04y24NMmxDRHaGazKwgmaLYdsAnWbqjJtd6/4gICv
mqR6a56psvhWmHvqkVyzgdQuf7nczzd9AtRF/feh/JesoR+inx8Q8jT2rCzRuJ26+uuyruD90fCR
MOYFgfTE2AYdTdB+jpMryhHVuO+otpxrvtHgFYDXN/HdRt7nVpzGVB5+di+2kmQ1gvzlqKiRsA3r
zOl77zBmmuQcLs37aGzdIuKl4VCYjasEG39RDGUod26pcVpfMUkOQVW79dAI8NNOBnYUuWwfysMi
DavFZq0Jg227AFfqDIA5Pqqo5NSTauVBjCzMBod8Zlh9XmH9cr7sDB8jfGJtU9LLp1Cu2WE3zlsY
WEcxfvhlNWW7/lTNvfxZCq7eJggXUbxNfPvfb7UW2X5hbJ57NWht3CDZ0/2cyjHFe5gGfid4guWy
35U/UPj9wPhPFrVO+4hg8tXsA/zwasDlYGULDWZBx5vpB8E2hupbkEQmlY2jiKRG5+Zg9L9xY93Y
5blirunz75Tn639mJELMOwNcRVE/D/ydBj/C0q2Au5f9/7/B5ahyMR3Fk6ViE344NPvMnp+s8tQG
A9B2qhUdX0+3vQo9zLgtjkoK8PqKKVtPDF9xFYvJyGRels3vFtuXGfEDFq1QKDgQdyLCijGyPz3W
hVCk213rtDuaX4XJ6Oh0q0JvFx1oF2D5z8dMTp27i/1MuDn203zNL2LF8cpDv7+ubdBwRgLIzyec
5dlMnH+Ixq6mUeFD34aJEAPu+gA5jcRVU+HHMP/uRar7+Yth4LLmJEomTLtRALYysrJwTkyj2Fu+
y/pH+6r1XeDkFrzetD00A9WpH7EypOdMjMAd8bs5d1/aEY58j8QkIq8Z5iPAEhSPzcond/GrmvO2
jyJaLLRyCru5U6HndCmuMgoyUT9cnAln/CYIV6bjCa8tcrXRA53C/CkpSR7SrktWeZdtOhTW/iPR
3QzGLwSCaWRgHLq/QZLIcSd3DxOIdpdviant0HqAqm/eifMb4ywHTXVuSRh07yIWc828QyP2Aob4
Qz4eEa4AaMelbCzNbug3IlksSIJ39doYGaiRnAFsOV3FJaA91lT8NFo38rd//rF5MA41pwOzsjbq
ok90V49/iVaRuG1UVjt2eLqU3hui1rh+GCfxtgA5PvvWN+xAhqjJxn0jYA+dC/ZSeOVkhYLa9BNc
gDBjK2cHZv5ermGu3OuqQj06AaHFrvFWnf76zmGbXLv8d/XP2XK5w+SFxxCQKog6oIsfYFmMQHzi
5oU/amc4tez6Q/3bc4NdoXOUcLPNBCz3klDwQJJwQ5bjD4qsIq2RwxWK8NxqoQJ3umeI4cW0tQh8
fPEPApzBa5QhKgXqQeXyXUaUi0EK8SgwXPALpKDIjN9DPpg1Z3W/SAobfhbsn200x5l2WdnhCexd
zD7V3mSgMC5QcAZMgwrVlNiTAY+wMk8k0M2tY7MmXtIENTfu4AtNaxURpkWMKCPAbCg4SnY/N2dz
c0tJ1+vof53eXhdxJv7fEmcTIZnjKB4qAv/9lM5W0cR1DwKD8WAH77UKGgFBEy5h3RciA4WWMfOP
EIWHPO/UagEJ1YLhqRm6M4+w6T/B9wqR36w+H2fRoJITBJunayqT9Ekrf50gZNZnq5VvLlwxlUoE
tD6ttnj/RYPJXLj8bvFtZ7ijq81jlhUmYQ9o9B1oOnf7TvX/h/K++WR6Sn55PUlp1byQzEgZxgtr
TJMLpx7Hh6GQRWVeiAVELpTqGlHNmVIuQSv98BK9IN65aRuqzt81L+mX9DBnhdNlTbjZkZ93xdEM
Cc1tQ8l0pvLKBbvxr6bQqGdjisQvHVrUzJfv3W8+KXFhYjROmliKu2uFvbdXLWsj83dV+P6PrllF
TrVPdv0PrjDu4ZDe8ZzXAcyx9mb7UyIn91pP6VrRsKX0POmQcX4UcFzFbi420PslI1LJGvQHfz2V
KgTAkOcCl5+EZfGNsu58DAAjyc6Bk1aqkqm4/X3gJIKueQr1xD2eSiXVpixeGz+RaUiowT8KS7XX
zm1LlfOh+mZ+A/xN56kSPWf2lxPgz0hYJhVG2YrWkA0KUXTVobwjGvWoG/g4ihybTDzFlQaUCbPU
z5DQ52m1QxwTceI+MfdKsIG6aYxWcpJpitOWvKsb6Z0M60ABmowLzcLXqJK+H9bmE72M/at0T0IN
8CSeOUPiEToQ3KYAEtJdhbWRg63ehCxTA+cL6evoDu5xCkY6hevqL8HIs7xTHmSkqEY6QQGz88Ym
TIzL4A4yZbpcSwPjEeubCfMatyyyVDnTzkZ1/X7UfcV5ILgEMlbbJ4KxbGGr/9UqD7ukKkiqUScB
/XGHBSYzK0AVnfrbTuNFo+dhyfA+PSxQmZa+im7azTBrOpaA4IoLIOO8fePleZhn+h3sSYupsLXc
Skx7m0ZaiqQgiS0+8P+weA96d3NchwhHH06FAHBPhQfQprSuV9M88u233+QgQaAzuC/yidUUXDX+
Oa1GmyQ1pSWXhmVGsUsDYKM3vuvwUfGULoSkt1KOQLRLEMZNnSuyvhBvIY5iY2lBymAnvAZSgJTz
YyBz0/GXsAodndVVut0L6eCmhXggc/4XICMZDLpz5tofErfA2sSlkxYXykLOYfGCHqoX6MLPH7KU
obzmnegFAhn2pkgctVnA5EVbmjWNL/TBxclr+sbyTLxdGchlLh/VXLQbg4hLfN1phSib2vLf0fsA
zaJhyl2iJ6E2GKe74mN5iQe4O3Akyr7FtpRorOt1rkHDLZCSeOuLQLt4/PvtmS+TOsm+41FITZXR
HTh5kjURQQDy9mBW8IrJoVeNkoPVNvFDOKcAC+cWMblsJBje4RplcyeI5iYEdqieAF53FK59JAj3
hN/enAMz7RK9PK0ch7yCNxPMQ6w2oKTxBlVBcWycrNDdlG01+Rgcz2SbvnnkbYfInVlQdWISo3L4
pRTE6JCbwar8QitnaKH/IYKZlU+R3EwSZrbIhPdjGPSwu9/2JRRpJKwcu8LvuVOKMhZTfUZMYpQA
HlKIqNt073KZgvOlpDyvrZdCW+uXMUopHcRG3jsOspKM7JxlorA2brlvmxoPjmB2DJqQBM4LoYmN
zCKSuSUwQuUlPDRtZlQiWABmDz4R1OKi5C13kVLQBmAcTFpaRp2yKM/6CnF+OOfuVDLmDk+LJDCG
7IINfAOhjzgmNaetPMcJf1kKHO78ayvJO86UpmKudyH9REEZbbIEmO/D6jOqlwKkh6PN77qonZg/
b8tmDQ2U+YHxvb1jthZQYkfJwfu1V6d8BIsAInRiB8dIFBMGVoRGKQktkbsOwm2BIacN0RxwWsiF
3dUW6pqlr6dOs/DYws2j6Cb4/qZXuTB5DmmfzepFSLxajbx4vNx7ngLvguIDLJC5L6MsVirekSwD
ivCiMHTQjcu3IoZI5uLAMbkO/5CaKHnSPkOS607mNk/pqa1sl9nx+UsQ7jqW1rX/wHegvpaYnz7l
8vVR3yWu0+hwt1Eg9qeQGbdT0z0WiY1F9Nmvy3mXzv534Ghmw4kCfhQyRUOMAguff/Z98HG9j8nW
HOmPcPI3zlPP/3fUghfCoKvx2YJAVlYRLHF/xVQ48cOaissffcSMTu0c3EN9mu/GoUvUMJQksg3d
4tA90kKj0RPNCUVwncUkpo9bi4clJyWfU9R3wvZhS/bL7E3qJOSh3nXzBXQwFNS42DF8k8RQde/T
aywzNKaWTbaTStxpeMApk/Dhvj7Ci2Eu5VYod6QGKoyX9XvaSxs9nudY2dtI5yQz3wgkXKfOeFHr
xjCAa/KHf1hPqsO3nJKB+sveagkNQfzAk/JsGTypmdmhY3nMnHd8aLCr52qquEE/1xUrIncY7Jru
zzT2JW3rdS/OnWyIwDFv2eClyriBz4zrXJtTGQvAFLlb8I9AZGpl7Ox5/7BsX0aVot+umaEVIaxb
dgxRhnYlNwqOCjCJGJCdAqVKV6wcMO4rj+gRXvGV8zVJmbiFLSe6hq68rrmIrIFUoIKSllBHl4s4
ew4fy1gaUZf1APip4XnGH1Hk9O0kMeF6hexLCS3CSi06iS4VbYNVpPstlue6AKzhKj2Csf/TurDO
8iKM9bkLm+1W9OP1J4zRZ+NWzEPRmk8AXGDcLHCQ0kKm+fSxduXAzdmxWl+Sk3/909bysfnm7871
4OoKEpAKilZMUaeroN15sc5yj5IxRbCnfhpRVhypBBiE4+bX8j7kHu1EJUtv9UFmh60nKkTa1pzz
rC4RNQ7/oFoK7Qj3UtIAFs1A8QdcyUVpKP47p1ZOUZGHEbxbHFfkS6uf99yy+scSampN8rKTYSt0
GWnK5mV7eWKy5fQ5UBNyVtEwIseNOR2mbJmNv2mQ7IJVR1g4MSWNTdgZ7yNEn8PhLMA+VqOPWjyI
UnEFw4v22A8GC6gAvGCgiVArK3PdAOGBHh8Ci92dddfeTGob/Nomx24KXCFtFyzOxDUfj0MhXNXH
fAQVVk30cHTeS1koPmv2RASjUC/Xx+JQwkk6c9J16cbH0t9I1zwLeS/rh2HPY5aOgD6Pe3oLKYIB
dSUNcn53FP8DDlZjXvOQc4lWvKt08STBNmY57CL5KZHdrYJD3EOoIlMR/Nu618xK9UugNu3jRcHw
sAgTIhEXOGkw1hTQ54kLQKwEJlcmnercaT8PW14+1x0uRAL5ISYh2fhKzBTdKp+dhGyN4NXxSvIG
sQl8XveEQJ9wZRnLGgr9jCVzeg9Ui02W9af0+bL2nBIUk5MTUkMFIhHLHF1MmF8Q4Xo8SmxPzDpb
8PlLGdzvvkxikeJ0hr0pJnqL3yZeOjIcPzJu5Imf1BHapXsja9RPSe7sZpcmeC5MeDMkTCyvaezi
iPmX5JAlS1WvwZgOwupmM5r716FPFIjwQd92d8VJscPqc+djhJZjjoQwPXMTwG2Q5LE9nSjd0Q47
0KdVhXpbbjhqWnyOwdgXzpe/GnsEtcFHatfi3MuN2QlN+TTJMomNU2atVhRoZTVSN+5qM2/eH7d/
nkWt1jpHtm0xWSd3W070RA3RPj0aKAhA8eYIm8KG9nb26nLrDMoNGCJfYlM0UhuYo3kDnwJAt/y5
S4UnoA0+LdW/1oEG5dhFCKFItgl2vipkc4g86oFW/plHW+jf5In5k+1gnoslfT1mX9iP37Que4R2
hCiOqTC3paCSTzK0Fz5HkVtchAGeiqffkUCgFlhbEgUEgEJt5GB0QL45tFL9Q+uIcFrySQksioXU
3QfOajvJGAec6YI/7rkz4rGWTAhy+zDWrGEtMOkY6Ohx2RYaRYZEjHmSntOOLLhkyF1rm9SEJlYO
aNbWQv+FRHL3Gi24ubCHDG/f3hFbS5qodvKXiW4smoY7wUoxoY+zYKNoe26WwhunmmKSS3ynIBdJ
qSudYfwBCwZV5kN22HBKENoIncn/jlqHrRWxIAsVpEQlUOfC8mPYdm3EN4qFN3H8eWOkxmA9bqTh
HyqlJZefmg+w//5H9Qc+xxdbcAH56L2khWlHgElJVXL5EwaqNKylfVgbrluY1nsB63skZL5YWPAA
qLQYerwBwm3pVb55eH1VcFdLWcjGyLTdS+wmkm9YKCr2UPUoif4p/+EC/ZgU267qHHaangvq4INX
HKjQK58DwZ9/mleixnpsQvsvuobIKLhaq4Xh7hYP51tPwTIB5q3d6RDlEWNmqDg24rMEcG0xI7Me
HzdVsqf4EKu4Ah/zocd4c79fXUUDN1OdTbmDIWUmoCs70fHZ5Rr3MyrtsbKL5Hnw2QosAXDmo8jt
x3ZNeRqbwZxVnl2+mfhAEYoyXau24ixTiW4BsWYgGFdtKGX9DLkcaLk/Z8/0sJ/+Jwm3TdbByPni
fribzw42bDqcLteOFfk8kAQJXdDQtiPVWpE8ErABd5hHMrjUydDmNQMuNKSzvFUnkprxCIJbfufM
ReNQoeieRlGcIUBB9ZkkXOYtsIvAFVq9/PZ57nfsLzgiw895jV8ZQqnT3VgYBhnfMcnpInjnNncE
YY/TCRxmeEFRwHX9OzUM0XJbS+apmtxYMKo9YdmKMr+9vPohIT5VQld5yQ09Zc3c2q32/NoG1K/S
CJeqYvyr/+fzcspqwu2qKhs0vwk4f4RcEYpRlp5AuraN8dnw6IIC+lLOuMZWYrHlQTgbdVCp+L7k
KBcoIYs+c+C+rERZkqMEbNaffKxZPmqxglG9oIAoEas9Vxf71kiJQkkD9uDNB0hViu2gk7Xn9BAz
M3qxBxcH/1fKz6ASxou7DjTVrkisqx3TgNsCAhRn0OyKiA4A5fMirZYE26PjD75VyryvlrFqcTlc
dBr6AIQDdhIWLAvkLAxK3LYuByaOlp5siWZ6yijL4E6tkcWnr+gAuzWddOkjeaQkZtxuy64hQmcR
zQkLiwrafggQODvNYLEhajxbticWfQtQ+DOlgLBmH0U2jA5vs/Onu4/qOKEpxHqJD3KLnRgOpCAP
yD7Q4oCc9kqb9j/oNSQsiBQDHodVtRDYajiugsyo73HaATDoOIZRGKrOWujHORVY795TA8tLI7Uc
FD+OZJII9vilj8C6lYgQGiLYKO6pVbS082GYyn1doDxQN3QNuoIoXPBs094X95HDVxrCoCvhZ0O4
hKGsnzrIiz5JLuJY/dmqKJ+c/zLCIqiQWMV3brcb9cpcfhd0tX/t6+rzEpAYGRBRKTJpWozBZg6Q
ZU1PRv05x67j3j+r0v8jElJMdvE+nlM0oH5aFd/3vkja4Z24CCH8PSG1bJCgqWo2Ilt0q5rRndRY
Ae2sJeJi9nf4jMMol9WwV80XouzpdKu/UgKh78pSObnNlS5bEgJFDLD+KkxwVHDa3wLqRZIUTF4N
w15bzZJgLzhM0WzGQvvLyi5vhI0w/UrLJ76GPEMCXKYe8BMt9f4CYLqe1xL4DRKW25vzz7CHitde
SuhspZaYqqP2SoyS95FMl/Jg7j8+Kx2Tq2hdKPj8j6NVr3CGdpk7d6dLFmJjGa9xyFnX2PkG2QMB
XH4TSyAVE/nee7k1FNcY0P0h50pVhMF+NOmeQNvFfUAiBLswBSTj/3eq+il94yqQK+BGbw153pD4
zrdn6mqP4vsU8Rs68GjDnI+bZvZdKe3G/jdAILcW3QNcJB0udqACLVv0eULgpgPi+XBwh56ZNqGO
kfK6Pxi/4/Runx0w1xS1JrNdeLh6X0cjf/8k8sTggRqyZH6mCtmFvZhbkvkxG7MyRqQVS78ByAB/
k0bNSNWxbMWTz6cdQi2fVpp7FFZoJ7hqA+/x11cBLKWZ5/Eoah1WzDJEovy5PX5kXqZ1/BRodCHZ
wLUYqS2oFc2puNDQ2isbQdigYoBGOzuma7e4J06vGW6tHs4sbx5t8aiqV8zSgeV4xaTriayqQ6ZQ
ewp3Sifdyklq/zxfvk3v4elNfgfGFYAmjCuvELQ0x/sO/1jqrMJBQo2L6n/gsCRyHauCWX1d7/Yh
pqzxFJeyWGkFSqXVGsHFwDh/Gy0+D5gErj0jtAUreN1BuWKyqgHDRm7xm5NehbFCXsw8MQ2J+NeH
dAM6AxGEVHg/avxmg4LKUfdQ1Ch1UfpCEdta2HemtEnWZsBzDPlD2lm9QkiZLCtQ0R1Nv3G6+bXT
o4Cu8KHQT2GFxMoXJ17tEYe3dg6MztpV7Z6/BUAprGCBSAuYS8nhfZZSk6nrqX25yAAffmdO60um
5eCIA1auuiBq2jlnH/+CBfKUMKasd34ZyuftPtgncBIoz81K1R/wKcxs8JKcB/8xAg2MqpJHHzM8
s6BcLyjKddp1EUY0jZP9kVK339NfmOHhXg+uGNdETu5DswJuxx6oL7ugEOyQS2Wbe2xwLx3JCq1K
l15q5tjsd1F6qO50fdehKLbMnTnyNsPE442DJOEjjE+NPPcZwMR1q2F+ZPhdN4/xQ1gWPsGKah3x
WUQBNjbyNPmBNG1FKeb+eNHz8TwVU9fUqk/sh9EFRmxLG6Xtq+GHZ2uDvM+XN39WLlyazIswVQ4T
nk1CMqmealBtF2OFCibiZGpQTT197bOd/KBupji/HBuHY2GPjKcbt92GBUFVDIiQB4Cej5yjosVO
Queial6abdFgNx0Lq9bUFaYtXn74R//aT9M/U9OXsona0iNazOLnUUcW1obZPyuaA5OxKfqj2Rh5
T6FK5/b1hNYiAlbNUVS7ObYnpW+P5aIHNtsZ/kN04zeA/hAVAkZOBQ5Oow3dNsfhxaCRhV4JT/WE
3iK+2vZjBH/E1V7u1UiQvbQJqVafnWLm539Xl0qsLJo2GozzDJxwYn9B22yEW6QgzuR5ExUwPBfj
2TXy6Ju6uvksb8LjyZS9tS7gO8+Bz7B1gb08GKH+jrzTXDoEPzudC3GrrJQrw0vtwycJtycs/dSZ
EZqaD/S8qyj+CgCnmIrqZzJs/DsC2NOt2/gsgKC82n/wY9jrwSu4/fXkJZa9b/8PEANRBqipfkNS
oD0GnzPBXxGIGd/GR+AvawspNTKM37iFCIEiXmTdnabd0WHQ4WKIfN5ys4MMMP/KzeG7zYLN0Vej
yH7CxjGGyhIiojMigopFt8MRewoAZIc0PKdVnJzNVMWui8hS8UWtIEjSViUTCnimTbj0OCCNtJqJ
94Fhj7zCklhky2MuEXzbsNmVOJhOyYSSv5b/X3qRPpBg+JnQuLK/xq1yIWn1vWdhpVPg1pKSKTUX
9nzSs7qnAqnia1hicYUdR2ffjVcAaQfapyO377q7ympkiBgS5VlVMpYIpf7Hre7shzSWj4/FUl3n
dhgYIhu4NTztgUwkkhGGogI2oRwhzamNeSNZF9b/4p0oSxclydEyImBqc6jsUTGnmnvJVKuFOGP1
illSuQjBrhZvB7X56IIhEJWdepOf28UR3f6CkYfeKdmF4eH9CJiFzE48BY6m9/8HFriLvqut3UUO
ijEx11eqlyk8pX/6buj4zW0Dgn6hgH8r1ibIvOVxULNrukcQIHzz7+HwwLixRwHE1UeQicHIA2G7
HH2kOadPu0HcgF6LSot3g4jNeHCjJmyIPkKXVW5Ynau1QPRDjEb5QQx6Za1JCXu4DVtZIa8WcIVG
Ob986MdNgkDJ8Y4yM4xfNDlvZa5AMA4qZs08N01XFgjiWjxZW9xViFtbfxH9nGZBiRk3wOMDqw2w
arZ/pAOlCnpSlCZ62y5CEk9ZmQ8hH5bKoBkeywSC0YfpQrA0FK0g3s76iGhkQ1faTOpfV/M3WdY2
/7c9kceHGeYHP7S63lez0vSJM6lnlH4wAyH5eBpP9WbrNTOHkmJjKOIHy2BlnvgeUs/LzrrFq1ne
s4IsAnj6cuMY6bLr0cTtg/1JDGomPorBqMhw0f6/QOUHHoo6z4WQx0g3CTvEhsiz/s021Brm5GPE
8Rmsyg5lIenQLECCHHtRvkXOYBH9vqvkk0z5f3MwJcCtJt1SPItiyB28WbLL3mrWhHil2Kh3xG5X
21DBKz1bidlBRkx/zsCkhvymNZHxxvb16vwvcFZy+HcjkYuRHwnJmOnBAL3tILkntCyj1nlSJnNC
xRLQU/IrtxyDFaMBSl3TCKFdyOdbJGP63jVTPPbHFcwqo2mIkJFhvtKBu/W6OLtLI6OP2mAKeBXU
9Gf3HV762wwp1q4boSYRnIgLxEcf4WIE6lQDfWl9PCAo37TRrV4p7NewVCy//7m9EewBhb9PON6m
rvYkkEBmjXd5QVQLeSqtjj/farfilktYcVMwU3RCMmVQyePyJqB8BCFTAY8ShuEieNgRmdVVqSE3
ZrFdOVTMFnEYTvXR0y0nwNmih/JFsjKeGxxq7BHYKwqqLAmLDc24TtlZOJVUkrnYkQhmphwvz1pa
iR0anGPToKnVO2SFHneJ3mm65EJgddElYusZosit4xl38NNCrl/KDrinOgMqz97j4nz22e+6ZLCY
dnqJXvXa1aRGksF9JeRt89GVBm5HmBil5c3gwcthf79ygSC2dUwk8xDtjQN4M/Mah8om7Mt6GrWf
AhUpbAzuTA+E40EM2KF+H1KlZTGxb2e0qAUL/CKrMrnS4LKNOgdcZQAU6wjKo9dU3SfeZCyWEfeQ
Kgw0CKfrPSg6PsGu5yGVUupu57SI3QLK2k6OU3x2lJsoTjjPbSY1H7JOSZYAVOMvDIY4QYTDvr7p
4S+WxLdCr2XjfMuCW1SaD4oSvMzhScx3bbYvgH6svXyFfRf5ARvRy+JG/nbJ855DFZUvqmY52Gcb
5Qz/HHNnI5P2blArLs5oRE8hbq8i1AJm/2a700HDE6w2DNddYMTA4O9D5PM2lgOLDWoRAseL59xs
0Dm5qaJf8EkHy7eYML0d0mfvrgc1DUbHFh2QJ74aS/U5R5E6wx23vNa7s3/ih9SoNY5VUHHUS+t2
YYGxRdK2yEu41gj7f7PDqyu7jtnBR7UU63PqsNOQjgv7vXKkW/pgZwzlBSU/lAfer9JM7nOUH6lL
dopvSuLOc5NFJaPuVfRrc272UjgJXRGQoKX4nv3SKMV2SMxqcZRcHkOZ3PfuPQs5/d/o0/2HwZRM
EDDWfk1SSBJdvYjxCL9vhcMziTOFgLDnJTp5jmE7ATtoo5Nz7NJbQJPunDxCdJppNPngEsxSbYn2
O7YceBQNR4ToiMyKZpidv3dsZ9+d0dZS1fzAQZJBZaex0Y61EZx/w1QB9VdToGMmJoPAhdjGjuo1
QukLxPnL8594qj6ORts2/hx7p9Gk0pFEkvm7zl3xCPclb0VyZWsMwiAZzT/Pm665fkm28Tfq1d+C
GNwjsJTR/gZuLItXM52/X9QPWcDhZnx0+2utj6//Li7q57RG2qRaatS5wRqbv2IOnExKtObvWHiQ
918Kp5LRxe2mR33X7AngaT14aejeHVx4xi3SpKAq8qTpyUbVUkfHgaZvhZ1KfCLKZNPrTxkJzQG4
SEgSJJIJyzh6PL6RN0kRSyirkwRFOMk3sG3MPELG2REiA/2hzMx0cx99Kch69I8yoySTf15CdXMi
j3fFON3LfjtCkJYWSmRXgWJbTVw+aKzEwiMEF1dtaTuFKyMdKaPC47SQXOHRx60AMiSn/1UBNu0O
DxS/HueVySPD5jA5AOhFQmpMIMr2VSnZE+cS1O8G6WDlmeMvLFOaNVXEQI117YcCdz5Va0VGvkRX
x7DPxCuHtxc+bnKVkNiugpyB5Lkpz1pW0GJb4t0bMHre2nNjhSraFgmw2GG8YX32LGuZMCzd1XmU
SBQCrwEkeoilT6jWy7tejKnFYj+7gXVv7aMpOaNP+GpcniHSeeg3QFIOcm7GuAgOAgBfD6YVMo6o
pP4Ggcvj9t1Oy7F8oUJjUhXuwUf/1gPm4+QM4ewRjol2tUuBXfSROLSnjSF9XKRKIOydcWogI+RC
rEEBo3h0zVOu8CzDUJ+58j5iHWw7hoD4jxDQ4hY8mkki+beoVHWMjeUgf2LgzenNPgdWyuagjsQX
V6Pr4A0CqJfpFqDzJI0H9CMGSqX18Si7c4SCUjl3fIKOqz1hNOHWpgREMtAEEm5eIqa9KpsBlLFR
Tk2lNHcOmzcvq+r6lCjhnYJEazi1pzEbBGxVdzUV+LIMvxN2zAr1ak2jJKx+dAAKL0yOJZPoBSvE
7aTP/lzw/Dwy8B7tzs1Zn5kp+1ZyVG2QXPQ7pDzJTgV7X3cbC9dhwkBk3HDge5gb/6XRlyy5XrBR
zyip2BAn7npaNuJap2F7WnayOQB+ouRb+Mn4ii0QQs+JaLo5M6NUKfdU1XGg+zev6aCo1S9l+XuO
QtApIDLUex9UK9BzLkOvW3X2gPHtRV16Kwrm6JqqWsOGTW7Tqe9MdJQqnCpR+pUMyFLxPAbAzPwT
X+elNPwylK5BtIQOvi5NOy62/tLnNfByB0bX8KBWIEwSrU69e9LaYUMtjdB5sotltuW4kjo5XYRO
4nhFBdcZnjglTwWkeWIpot+RfSKR5snJDG4V9PWXWjz3tx4as52AOYiUyZ4YhQK4lvOkVPIygqo5
bPL5wvhHKXg5ew/ey21yK0UgvtuPzJEFIjyY4Kw4mROKHPOIZsXqkqdJ5Ul9P1hrVePJlNwRd7U9
tJcGwjreOUdr2uvrAL2PRzqGUDgippfRxqDXb3G+BeyD70KEJs0KrjwNbMzHfOhvoj4lvDZPM/95
VveOHR3oFyCYY3dqae4PIvNwkg68OwzZ88OO+KiBfl/vh3bw/A3BYR/4mjbady07Bp6GFHbG7PU8
4rerTwcqGs5Uqg9Rdte21P7zp/O85vs/dSvyWX9ETZ6mHhgrpBsN+Oty/uYGqatQTTtF97uljlDk
2+lwf+nAP0QDcMoAhpTFD2x30SgsBqnNmBm2DVBd9Lss9IRmNyNtaPf373wG8cy1gEVoS1Utehi0
6ggiDz/K960nkmiDlOy5k/5iP2oOrAce6ZJSVKrU+gE9trPIxbbo9RJGTXR9rZm160wg3OkQ8cMm
kkiaTNh3lN38u3aQX4jKXVb2YXohXZHxu77WjxZEXZhmQ6US1mXk2Z25m8yD0zhecwtOpEnVXR0S
KlEMsQSzqaXWZi+hRIJ3IfuRwpkTZqb1m334tHM4p3BCxz6oDD1pKXCMVOlecKt2DdAlzxFX9pDv
wCab9D1sQVVRMqDBplKk2WVR5ONCyZh7fdtz9jfOEPb2ZNBJ37kpOI1lX8xirc39dtjLLHuzjqbW
nTuJNuYclMSuuiT1sUGDZJwu56V4gXa+zobw3ayTFe6Rht910gQoBhL+fGo8PrXop9nLYM2as3yZ
w7Oz8ywAynQ29RBSYm2yGdg3azifM6vnmaAd4XPxSC/vjPccFlnp4mbP1ShfvwDCDcn5nrYssnbE
2cGQfpeRSGYQ2WWbWnr/624vZQhMmqv0GuZYwWXkFVD5IP4fenbM5U11e9i9XQC0g1H4DfRFWlly
AU2chpl4ApM8u2+YbrFSx2jabQuCDfqvb8wNIILhhCwcSCulN4LOd6dQyn/9XeWebkOdrr/T0fGB
bpLF7dIYoRhAyrsZ+JWfzpJGg8iMgNQ6ObBhVPcEI8QHLYZkQZK9/DLPhWOWBFD4kwXdbfgPb5+m
LyleVPyM144PhiI6fW6h1wu/StL1j89WsPMzbN55rXAHvnOtoiC6DCaAfqs5UTgOrt/nDObcDMWr
Eqio61zEGUxHh42WgE+0lOA2ZYSpYugiopp3uccUkR/md2Uhb5Gfmgk3w+7XRue2/0CDgbKz4qc+
so6KhuFby+ENiYhB5bLw+tJ9rrdV4DY4pXC+25s+RcOA8YlR+u9LAooXmWeZJhN+eoYe0t9vXWbm
5I6uHtAjhXvieziyJldKOsQ5CY6zzHDDcrkiVL64z6+y5IhThtHzqR2yVNeFIqjIFQL3jqnUDzTq
WVxOhsQrEiPp/G1JSZuIdiQmXrfds+EB/vzHEOU+VP9hFAcxvFatnQ1gCpp9KdGrss0gwmJhgYip
QSD3kYOLB3nbHAwb9IBmr/7YA08+oHjOF2Trg9baft3bUXLMIzNF9tpe6a6mxT5b+nTeKgC40x13
Mrh/RJvqiN2JT3cFymMNa268ox3VsH/q9mY/mkHm4Qf4nHTXxE/XkCJZ28jamIHJMJYzMcO8X23D
XYMeOP/Jncr2rcfSZc1PvZahLVqoPV4vYKQ2s/Zy/xa8UMN9MpIty0qIE4vHDZTwrh4dHw0z3/E0
TJSiRTf4+15VuITG67l6GTz3BWIc2a8C0lcb1RojkYiqjKo06BRtylTO/3kI+jCfUX0a9uBPAmkg
n0gtndSeDW0uRwuGkh+4as0sge79nTsjbTKpe0x+qmmaH1it2YBhj4abBuhNE8slZ9HJcqB08xXD
tOYOOuhMXceANgYeTPER4GNxsL4nHpc2kkCjmTu65QvOYYn1sTu+YaT6Wgw32w5S0lu5QnLalSbj
Gb2XU3BpAFucp+Ee55p51/1EHpYPgT624JxorXa5Hu7fsuXIZrSS3R/UzWWXECkoZLeY+tXjGwdL
7TcCmtylSj0PULykqqnT4PbFmfi2dH0vjmgELO07FXDX7EfUIKmOXK2ykHrE7bLkJuqCSID9mDL1
XIdpimjuInqI4Zp+Z7NzkcWAD29LRp9aeMrbonEaTP9EHHu6ZoDDookRRNygrmqrWt9uVRtZevl6
Pja4R/6LklyAymbnZg2z2P4qv0QME+LDtB2AbWkoa67kYTKADPgU9n5zPMqxKNT/3VG4FNT8rHQY
Dyh4y3EbWflm2AIHJU1g5LrckOlocFPI0lVAraUsOrNuVZhZUfr3CMdDXM3pDILMTN+9IaWPYM/r
UwFKj80rwlh5e9BljaFuy5kQ6MVHFhI5jMBofpriJrE058pL+UB7TVU5/qmKmJug++R1kT9v+LfW
GG6tFRDMg2e5zi35Uekbnu6whE9moj1AXnBMTl0Kct8pdjl5CH2SvOOGK6ahWP6OQWN/OY/PMk3H
tWB9iC8cY/qFU/T+lqkrERRWzZaK6HlWc2RFyOljCqwDoLZ3Yse38btx8qXhAroIoY8V1XzNENf8
g410hgBPkbhvvG99ASevnnHGd2gE5U+cQ2/RxkqJTTlUZvbb+q+GiOxDT1iQT3YfN0h+NthXeUh3
k1526IpuOvzBh/M8EeD+lhMLmzceMEduVSSKDQzQ2E1LTscun39vaAFoilwz4vAWR+17G7BiUBJ+
/dgOd+HGPiu0KZ5ySyDS1WlmVio7ErrHFWyjWjxzGMad/8EnTXnhhlfT21aPsP8p2PRWUG/ZKmX1
k0/q+u0poqJj+tD9swvocRk9e/Buo7Z8KkrEC27h0Pqyi6Tl3pOIx2l828r8DUqpana2Ifssygh4
9NwK8QXDbhFFf/g6GM4MN4f0rjUG/KTKyL3ub4ZrEOogACo7eOpfDYikHzrcpz9zSKd2K9pXk1wd
d+FtjTfNFj7K8XU/0Tg8I8GsQ34s+yJYHQmqul8TjVktN06bj5IiDhsvJDn7VW1dpPXCbn2cjCNZ
+iTOt4X5Fog+RQsIZYTdYB6+koT9wVkQFBXNsqJMmNXXyaUSyG8KMJrUylwSkE4JAKYO9Osj2nT0
n7sRBcOorlOpyCX1E6VfkWfFNyjed2jGBgXNLxnWCyS0Db0/gCEjRH6nrcMo/8oePigqlmAgElfw
iNKm/geQNP3MQicOvenRIi6W+QB+v7AxiY0wj2s5otHbn5EPLq2IcRajqwjWl+zmQOPc/TsXcwDO
95zI8w5+ULULUDsQ9lFyHQhWq+cD+orermQ3jjjKd9Dsi0lWO39M1CGf5XilIGM8GY1i6hJC61ZH
zSbV3u2cHDQdn3yTS2VlCShiAjqULp1Ta9KySekiXfXNLPy0Y9mJKxzVKcBKFXWtG3IAVGbgsHT+
QPMuZbQGkKVSoKPDhKn1UPB3NTF0gFHiZ9TJUf8qfD0u77v+otbgnfvkSb70KcU2FFHeTncGYS1S
6vp+UULHG+G3xVd1YNOJFngmtI8wAXU8W2xgbAe5h5FzjtxE6f2KwJxsjg0cDJwrggT9Sjfu8GS0
vtt2slRedrr+o/pmJBS2iIcEJbKQ4h/sTm5GOserVlgmN8GQDxg1oxdn+yXfSwyWQ7LJShyFfPV/
ZuvtszV78FyTJO7w5edtjzPm+8BqpgpYHgUE3eWHkiacGzfRzKCVMf5lvNOWBBGMYXvr1wLLjG1Q
VUC1wQVZxS4V2eY1gIdJkcePOAQjY6R4P8VbzNRf7M7Jux+FkbLpNJhI/jrKtsaqJSJayH9wSFPj
TAHN+QP5BdQ3dFjyAyTU27uZ5EFh4f+Xi5ZMVR5YaVJhqxjTlV1SF1Us9dzlc2Id91mdy6LOntbB
Gzdqbhj07CBm5NgvWMFsEvZAXuTs/RrUq3GcxCxGCIknJQmyIncO7KhLEVv0ChZcjZqxtCWU15gS
29ibdIMoUk7+7CKck+95vwI9bpoFC5T5w+DzZRD0Ga4lr8v3cAtOkpOL1ReLK751zmf5ak6263KL
BA2jziESACaMmECtPKbGI7CxeOYhAa+slutQfcAEKMJUgr3vvhAV+FIbFMkhJ1G/FmnMHoR4T2kp
oXMSREWJkJyeIAb1jQwM9KjeWecz0IIpw7vV2Ud/y5xSG+0wkdHzWzTR4fFPxAjmZ1aDEQKEgahJ
02LrPh9n/fde2ZHmuXXLi9/PrJwNdz8b0OvniqW/KCD2KbSnrN0qAGzseeFZQbSjHqkPJGHW5efI
DRzKonZHKKydn6Dz1S/4g5NOR/KlGDekhhTao0eSPjuegJZSOpJVLfm6LSNvnZFM5v6B0rL57Umd
/i535+Rv03kYzNda5ijFQMk6D2P9uH2dLRyxj2DxM93oGWQJbHaL9Smi03Xj2le/3WmaShTip5Wg
j+F4fgQcERFeFp8ViIiDFbc56UlqlJvsOrjKykAT4C/qvtKwoMsu/JyOui0a/qeh8owcsNmsU7d+
qSdt2napLHClvspRSPhpjaeORkYzGO4/x9f9Iu+7j/oA0nnZb1dPfJZqhaZJQvNmOFDkaLMM01X0
o5dKvOaStbBLOtlOzyPiA6EQ9GcLafnBwHtYj2aOtFl2OLXmSRywH+OgWZSrMYPCe3kY0u81argd
M+IHZ1nyaz9Rvh5C+B6oj8sZIaTNbIwAb290G++DMUNpl37zzm6vKL+Vokl4r+X+zt/dwDzaS7+K
7r8znQQyW9SraJGtKBQpMRhCpeLaTTFkdwj0pImmGNhx/lAgDpVmj3yaVyyNVgx38mDkIzFZdLwP
nfHLU999gj70KIGmjJL7yy6o2RYaEBNJaluvxjji35Q4Ag5IZDHebyq260KoIh4uMflvA2Sqch/+
O/GULIk46UqXKa+TUk6kOVkeQmDY2qEY16V/+sfj8J/3zgbdSCTcBcerneNCjj5NYlOK+F7hlF3L
NgUu7x4KaaxKEnmLt6Ejj9EIU3MmCk99Gx42fp1hnqzGqkbnxGYTOT+XoWKw6LOp7pGyAlw8w9Gn
FmiQC7iDwe8rkVYoKYd4uE+1Gs9ww5mGS+SpynPrrYrGKWh2n9ePPblARBlrFLhAbsyEOneHarb/
6Nd85RCp7JxoYxRDcm2EDkEHiadG/O03GzZUS7CPDGSGrf+18ESkrden4qfMfQpUZND5UFV0E/D5
6Qs3VzQOjOeMqBVllyjDod6/R46+sMCfDdmbVC8SvhWBUoQtAjkMd7085jenF9uVJIn4ioks2cnl
RjhznHqeYsTsm+S6u4hLm9dKuVj5bOj88lM/e/PawZ1LHeZARnxMNdMOX7QFjTk+MfA0M2nyAMvp
Z3KtkOS6LvWQRdID6xEfydBFfz9mLD4cocniO0ka+FYmpW8CtFN8AxVOFfd8iGyAiy4JDaO2izcM
8Q2LQZupknUWL/nXUD8nighJYUP6xzEf31p/ci6m5Y7kWjotKHASDgTGAz6jmYvzXx5F31pyiVRV
IJb07WTU8ia78yoM87XJXTiwLmrSCPQHqH9rqu8tCxsjuEhEP95+j1hHQQNAPXY1hsggHBttFjDE
KKotu/vsX0vrOcr+mlllr8u6vmaV/iANXVbT7R62t76UYSc37EtKasLY4gbEaVBBwMtFIqt/fULF
e3TOJtBpfvmVMO1GuvzVKcKpH6MUu1ImqwfbwRJOPTQnqTXPK3812WXwCWcvXz8p/jhuvZa3u9Hg
ek45uyKJmkgpnoDFItvRCe0QhP4+HQr2Ry1FpUkN9WMVDFXHboeIUIh/dmzdHOnMd6FVZZIoJzl/
BNDe5XtE6app2Mjr1klyNDOTbhuHqrbRcIh9dIbmEN28tczwiYNWZmnd4Vzk+qzJzZfteIz0+gfv
idlRGk8vCxmnLJvvS8uMfhaof08Eb0XJCfhJF7HtECN2F3gWTve9Sm1mlT06woHrLpRXDn1rk4qt
H5Dw8VQ2UTAFc8NmGbSpMytJSdwfOnOSS4EWVWgzC76ETxGPSXSLOEqqPpZXEww2LCRcWt/zVlmF
/ElPdjAwIgGgLwGqTpmlRAEayvSv/N3fGhhDW19HVQC3YNKhW7iSDVW0sf5BGLuMt14n0RqpYi09
ZLNxVSvh3B1zkomIIHqkoAOY3IFA5BWljAm8BfbO7q3EPwVUaX0DZ9MBDIBjq+J/N90GOjYf6BK4
n/HOHSNHkeqrc4w49Zy3/z98xLvZxt0k28u4eACxszPvGDch0AYMvJik3ImhdBzQMzbMly7IQSeV
ngi+bTaKa79VHJs+KOGVleizfpffCFf9c4ROmCF2GEEf2yfp1FtXTAYbc3z4+84AJkHcfCm0DaOD
HTP9qxODBBQxhU+ouDAtkoMuIKxfY4cyd+qK7PuJ6HW81F7qCMvxhvN3U3Vt2d2/0YBA8N6i7nP4
5Q1NcenQWAdnMp6niaKZTpGHdQq5Zh2jB58oaBJWPD5b2/VsxDh3xyGJ+ZmdqJvcP0uO/12d+kKH
JEiIE4vngfpmxaJvOgoKlw0wQOK63xtLf2Xcy6stUc1K4/cyx/m+HLTtfzCtwbyKw30qM0d3wt6h
u1kHHxagMOui6aABrB67FjtXSxalL1scy/cNsUdHkHpaUSFwDARgA7g3NnyB7PEWLxaBw0tLV/Er
++MU9OBAvLHrOfT2JybR6/9poW+b4asScbxDjhO+RwUlgDoy0WbV0DzEFLSXoo+HoAiZL0Z3IziM
P1FYV+LEkd7eJQAQ07E0Kg7gs1yhXqLSTJZdFEXBcTvD7LukqcCX4dNce1/V1EcvBGjJMjrbMDlI
mnhyUrjZL7k+H3WYDn2aqUvUjOZx88iRFuQs2AJD4QtGMuP6wwtrhV1h7PDh0mrbwhdMcqzHQxjy
WFSs4gcPwknIKHwt8lslBhZFMGeolQPzjcnY4Q12NU7Cac+We6hlWJjnrEP/+wP3y4cyh/PweTuM
gBs0EHHTdwh7gvuafYzmKtSNQUTz/JkzMdAAFzhypjOJXldM3ULdMyg0ZHvNYZbWTse015Js9PYh
2W5zfgzcMrBOtvgQTKkxdsEAP/hHA/4EK2UdehVxr/RB7q55OrwC6+OabVkzHu9OCjwz+10ZYuVS
vJW/vx6905/kNKkeMrwPG9litd5uUqEDT/RJnC/jesd8c9xvyQ5zIGsmnAsNPp58Jg8qTaYQflmY
mIsGGTFz/1d5oH0kbmBc2wwBxs5gu02sEDIQrDxhBn2ch9kVVyHMCcit14G+7+mV9xT8UJ/zt7VA
WMgZNuAhNlDM7xfhY0oe0v5r1HZTPLfLWwSS87+pfwQ56cnAiff5NYwt3RbcooOno0Lcj37vrEgA
L6TfbaGSCIKtSG6skQaqtnAOhSzeYPLLCelOiwE9HQvdYRAu9pTZUW2RO3Ra9HeGdNlakY4r0eBc
9VTOOgOW6FtQu36QLkIbjQub3jnPN5/rDY+mbD+gtMp4zrFKHa0I1KCPwaFnepMGOX3gg54YDxKC
qElXu7RALZdLPSyi2lfpXoHUp/KodlvU3YfcwioBERZ2n1syTF0fm6FSpPqGygJmUNpUcMMJMSQG
O4MJx0f9d4P33ryBMfFfgOw9YLZUVdY9x2OVC15Stw1n7TkD2fNaEBUszvGztU3ylrxJwQx7I8yv
UXo0NlqvwOF5ojMtckEfKim8HZlq8qjMzfCDci35KlF7ND0x97Bq7/6NWUsQ0WKGSAwtTStIwkRw
pjiQ6TueWWJXhpnlyFrFY5pkUbv9/4zAqx8oYlpOnBCGqqdN4AsOKiwPr4gkO/6A66J0bKI0bXKC
uluA6chz0QrSpGK9IeXxt0OREpGZzLvz8OAz0KcO/rp8JCJtiUGm5MKUFL/MJePv90R/PryxIWzI
QyMQnWWV+jENTPC8xwy6iUwXHA9bJTE5hcupGCdlmRQJuXrNiCyLF8Aps/1ih+cqleOByzHp0qEV
ASC3h7S6baCsl0nZF8GAvNRbkFB6On5Oe7sn0dNvPb/kyaxahJZ731d4/j9riAXONevH2u6Sw93I
xV9MjmGwQNWg5NgXFrwunEaeR4+Ydrloet2k+lK3JWGejnHeA4gmLexWwS/VKzadLom/0g+0qSd5
c8X+6ljJekzuNDPVB8z6AZpW9txarfeonrhRfHTy/Hn7Lsh+KuNzT7JnAPB3QTbyAfWdQI8q4/9y
ssyGt2/4CxqNV4JMdcKqRrmAebDO7a/aXTwvbjg43swjS9O66aZEolqSp9LVZq5kZF3CxquxdjAN
05dnwk7VY1A/DG4csVvjbZHryAMTXPH+ityVs4r2t3/+aeU47JwXrhNxOwcp3UIaJZ39Ye3wAqTb
4NIcvl64bevj67LzMjYHJowcuV4xnnB12d9ev+D1IfX1v1JvLBml/x2V7fLTmHDaKshpsqer19ba
tRECLqQw9vAq4Gnu542FfzJiU1+XbqMhsi4ZU79MotJezqKt1k9Fcq7I2EUL/8Ln7HUDSEzKU//+
zuaNwJ7nOFiVcpgW5LCSxdOViAo10oHHd89OQImE+bdnb74VpUdRNTxTQ1u5SqEk+xRLoQEJoqpb
vVpvnDBKu/Qz0o53GNzWX5rHrg6Ul1X2/CZJO1PRi7MzhsYYe895Hmhv2VEaraA4ERoJC9ydxVrp
BcRZB4ayJifyIUCyEjS92eBn+8XhOOl9BRoyhEcjJUXT3krBgx6uQROxuX/JNtaLm47y1OOIOGTY
Jrz6V/dsaXRcvzz0iY26h0AtqUO8bUs7zQkoeM+ysJa0UsI28h5b1W5LoMNENj8Dlyw7dic6TFJ6
u/byslKOxZnmbQmi0KiH8O97ZZsGgmhqx1FaVncBCvp5VZ90iZit9skOH6OeQnxh4TCVN5S+ii5i
KKY8LblIpdQR1LKtaiOTQKpqC7nKhAgsytoK3WQtfth7E+R57mmzHFw27I5V1pYeN9hZSGvRnw/A
RVrA/jxkfWAPfnKkvYvDqMEpjDaM4VdM+Kt3c729HkV3q5plZsqpwXHJVkBrIXpBJfvDKhqcSB8j
Go/IUnjbjqKdFrOS/FNsjjzP+88vEGIrytWqwovj/p2BhnpKCWhyP9NzVXyBHdbmUIV1taK+K81p
ubwfB/l+pzSduudM2Sxr7voN85t91eSypQkTL/NwSxwaIHDZhUmEjOaJ87IwvwZRfcuAhKbZI/jl
cdIRyvIlJYeD4xYmOz0gxD1wDRcue+LBinwD0nXsbrj89CfFoMGjpMFzSr5BUUotrOt4o0ad0Za1
VHabPAJia2+MyBuRUwbVVQHK8vl0Zc2v0YsChN4Td8afuQyUjBhlkoqCj++Kw0AqcddS1UCSgTEe
ir07ConUrBzLGE5Nl0C/KOuj5ZPj3dXmIxSgJHl6mkZw6kEShZuQ8Mfjy26O6yxPQP+Ql3vx9qvR
qPBISFe/KIaQxJPxtpmO8cRvX1HLlnoJCSSqTH4d7EZS7OOLQ+RwWHvSI1JzZrdCbhqKRL0Kjlhu
OHCqEdrPfyFADgagouiG2Me4XkIPuXidVEPuYI4iKwHbyznEhuWBhjOc/G+yobwvjEVAWKYamd8k
KBuhUqN+40fsO8seLMnQdgJTK/ErP+1eZc9ulaSZPfsJw74RHm8WfdKR5gBhk7DsQT7usc9FgvLK
j96+U5dcfUR0aWSTTC2ukWg/zB3zqrCpm4xp3HKgYqdiNUSD0XcUuiW1gFdvo5dJYnz5DR6nU83L
I+6jVVctTL/sO11lQB912YsQMV5SxraYfB55X0rLkjcyCt9qm4o874b170/5PmjUQGHmASzgutq7
udPWKETdmfP/p0lOX72uWWQxRHwdZsRkOcDPAaCXDtqP0H09eTPZA53F9z6TEu4hHnOVpDnXzx9K
dRXQKk0GPVsrTQ85P7kanGW8wAZ1r7KmyHJNppJAToKAGHIAceKoXEBLcU9uVHViMP6x6r2jgJhO
t9gYTH1+iyAIkQCS/ZQbhgLr0OzjyxuX32LyEORNyrIusiFLTTZYm/l24C7lyDfpo1BYEuO2rT4g
XY1VIoP3o30+zzy+2N0UMldjo+NZviHmSKn5q7bqtaXUoWICKhPGQuSEP5fTEVqfZt6izRmUzbj9
RQh9cDYpTViscA3r5EzQ9iK0QUPKd2pj6fSfH1My2RpzoBxJNKnINibJ+c7e0BGFpBs7fqcKjeLH
vtrHv9QnnGgby7GMz1/48yVQvVhEveF0djoxY022RdbNCp33d+P4EpefI2XH4ri7app75Whuz92D
EASzpuO0cxDNfkcgUaPEOScNBm60bUCY3Y1xBlH6W63rGP/Sdgzb8SFX79AHE/gsXddZoMnJinBr
s8Oi4VqTPEZbTBM/bZCEKyPu3DYha3CCkkcRP0k7LNd3eip65mVZFb47ifBuBMb83Uk6Qh6P0hBc
r7wq7mpB/0Tu4sEQNG41h06Y/cCWEuKUKiSp2nOq+zWxp9wH/1E6d4rwHyG6ikepVotEeF/y8OVy
zbe8234v/8N6HxX5TZ7Cw6beheI3djFwigsYi59rMgKFyGpyc4Yyo5CFKrGMlZiYSEQ0elUy0mZC
B5LhCH1bcsNVGXo5c3V9gOP/dBNYt0GoP7pG4K2HfhAp7/xbuqYjMTfdu03SYr46TRX+LDbTCGWb
9rHIz563OR1WsCgD4SBzfc0RikwxOcSlX6UZBwg1omDvmzqL3BBM2sPbR2NTSw4ENYVhMLAKY1CX
NEIi3NNxNHpCuLApW4uvK0YvRonU7I9f0FlbPfC56bm5OXZM35zjaOTIqio9PjffRVr21i3rD/7I
C/sgkW/pMrDtV6xeKkGTZsuJ0Ge51q8uhXVN6MdkDHqoA3bCyosvWN3WXJBqfrhXve/accvM2PUl
PgIVZfRXNVGrAEOy56K23O80In7L/iH9voq7xD7HyILGDfkyUVQepDiehbiIAS7lZupDSpZ3f9Wq
e+VGNDFdZPfw8rse8OLhL1JVlQUX4dTZxMj8yt67X8k8L9jDHseJBEii1t8JijaP0HgDQNdtOC/V
FhDzpEyqQurqWUqIKkKISuzCIZDcouYIE1OG2+zzvPm8a59/kO96RRwcTolXk5wvhDYGinMje1Fe
N5RuN/2T0anuc0Yhbq7d0qSa95Lc3KBN0nQw/B1T8PUYla99uvJCIT2K5sTI7ncti9mf/n47hzvr
EEG5F5WM/eEc4aOxBQ2xDMhINQEAaY7+LNQzg+8VUvlfOXBVdZ4J+rvNgHC76BW6lshufmBdjvAA
g5r6dPz0jO9pwUALTDtbAJcCEqyxgE5dgKaCMkKHncxr9hU77Q6PbuS/nIoVdmNx1uWrBKn41D+e
B329L8wmL3+uEQ3nrfvHDKZA8gCYEjlNnTHRGuoAbsBLihOcsYlUOfhymVRvU6BY4D8FNXde0sZI
WdSri4Cl9gpswKFB9Zrb4I+u85FGVKpH/X7EtYUlOH24mIvsDymh/SbNoLAAXzchb17e8NL7HigM
v+EyYbNVYzxXzwlW8c82mkZ4scn100q+POrBpmzmaWkBieulkFwkQionNayTL6jXkJMeM9BeHtRQ
DJ4DJEXIDLrY2FomboGPxK0MUVXFz9Um39qvCmx4vAjG9sZ6wYyAGlkD+m7kjDancAD730EqZ0k9
4fq5iVEq426ifp+6eSsfZVwmriFKSVtBcv+4wIoFi4bAyxd1H4t645JuC6yVHLXv6xOKbUnAWyhq
tvotzfpGGo8qinvzVwTYCmmg13VC5EZkJ1AgLD3Mta2wrOq5exmg0w9gkDBF22nV4SgwF0FHzsVM
0uFPv6hsYZNtGwRJaWPHZeAHWIezEnakqO3h7Q77T6gxV0jITZ26eVF/at5m8xpJMm8I3XOvwUeT
LtBMWwS4zxMOdAFUOUZEk9J2/s6LJ999xa8HlYSblzBnsH5qXKNeNC6XprOhpPy8Gtrvpk+4Tj/u
cXOwaSL1McO4STVMHmjgX5j3519qrvNPhgK9FJlRKcNS/L3VVdHjrwXv3ZaPy+P9B0IITY32ylkw
tZ6nLYT8D2xyV/i1IPFqqSzTvJAUe19/XMqGyQArMkf1gQqpmHkTgEVi7V6sFhHg8Enuhw2hug6f
bdNAlK77DpE4PJRBBlsracIhR09RQUdxTdzZda66s0XiFFAdJPxM/tBBnlMKl8OkvZuB1pwtZJar
G3PbzcdJ+OzLl6UNGiuloSP3TUxI1Yw4MTA5dnEriCaEcESwQ654/W6ddXWAFNNKaojfXBGLbYb0
pVu48J8bpFudKcqWYOwIatu7JT+I4Cc1PV8bGw7hQe4eDJAOSixmpqj8al9kz9+G+cQvC9p1v5kX
UvbTFvdxo7bkKIixQCJ1m97RdMkMFdozIppN+S2fB24mVfVrUcNFLHZD5tc0S+9FqS9DZPGGIyro
n4Tjfk2xs10kSiXxang+8NhS/45w5wUwiG5IsNH94jOxdIWNbrdap2cBU1wgWGbxzWyPR+GRe+2e
oPkDPYiE9S/5SyJcZtYf8slefMXSeYCSK9Wp7olurl9cIVE1vOhrWbLpoVGfljd/HmMXIx+S8D/N
f/ctVLdJtSNvKtGVSS/mt2vJkB9FMSAd5mf0S7RE8xsLh8xcrWwrL3uqBZwVgCDm4a8W5UG6rjJw
FRPTzVA6bfdKekoXKJjhY+pq4BiTywE8SFgHphIbY8esw5jYlMs1YAY+AXJm6OZcrC8cuM4K6nYB
ab5mO1k+VIxKMwyr9BsOES3gRCxPgmjdnpGzzvO5j0YYQSXQj7AbWxKI7UngrJGuc59Ws82i+KQb
e6IVd/cm+t+8Myn24E+uSsYoo6xBXzM/3NFWAxiOuqAaUdCq0wlflqxLsdnTosTLsl+l5df0AOx2
2gK8bCurJQ7UsF9OwUX4yOPwfnez1Roc0iD2svmgY//8oA4kmqOKBZcK7mGhYDKJRYTDbnRIcLLa
k1ZkPaUzE4jZFB4NU1DX3LQeKv6fmdS9QNwytzUYyXEdOMkLN5PmxcxUoQNEOP8lo3UNJLZrGRH/
hFo6VEcMI8roxRMDvrZ5VP3ldCnLCKHmur3uGhODzU5+h3/l/QCs3WeVLMJYXUyiZ5TAMw1mJRhG
oaZ/sua+wegQi/Kw+iwIbn5/DGiPe/vbHfT5qdHXfonJKUdzD9OFnQgs3rciPeu2/EnVoqkbXJGS
EMNDXKpHfAphKuXTR99ZbvWGn7tMaeuS4iSmwLej4dnAeOydZhbnNZLhX0DKpI4AcO0b4huM1Ko7
J2Ik1jUK0wSL2RuyAw1URpn/u41nJaMUzgS1maq/XlAAaMYg4yjjMcnMF88kA1MgKghbcWxO57If
BOrFu7IxmSJ52Uc+UOHKMLdmARjNJq2gDAQaxQ3kxf2DhiDFd3hzVy+WKweul0vdFWkr8vW25/JF
/Zr6b53QQN4B9cMQLRBTFcBoFgSPQ2nYvfi3NHSP/Xk7W1mE8QpVOlKTrKczcBXa68zGjxCuETn6
T+OzITQ5t/0c2ZAa5tKK/ytP680laaODtiH11ykybBKSvg5DQveg6rSp1a4XAcrLJZ/nHnoHPnAI
zyrYd7RABWNmpeBxf6FOnecimDQmrXiJXd1PiyRRKqgiaJ4A0LNiDnu50SoijDjv+FbOgQAULyES
7zGxK+laDgQLr+cnOn4ZSHQvYuAlK9O/YQu0PgPSxOSuODN92k6eR0PNpfImmImFt49REtp/3a6J
CVhxfBEIDWDd7Ujx9dSop69u287b9yRRV6bwbiIyXlXCIHx5vHxWq23Q92ojq+z+AzZ7MsILhJUd
rEf4C6rtJVxd1EY84/huywuieU5Ekml+YtGQFV1dreGGw1a9Du9NBUu9R9e7iYGwnIU15BI1A5ml
dPALpHdq33np9j1QxM3q6QaDmdQ4dy9nLaBRJho8aSLwGe0RP8s3ufbAHAkibr2jO9gObpFzAsNR
VEGD8lb5lzCBvKwiwvq85DKtPuJ3VK6BjzKQpIECoHtqo43kVWM3daUIqfnBJfl3nPfdlBgjqL0u
th3WYp4Awnsv5+vx1zEF1JR+4XHozRIqX7dVRwvyJhVjzNM81W/6Z8RCiFEfeLlwbd4FeIL/B3Pv
IRP4y8ygnyBC/EsqhZ92Nso1/lrnvXO4alWawXjC1/PI6PwWt8oQmCB8d4jXM8bFgr632Gfkioo/
mP16CTs/xgOh/ysGJlYqNXmHyAM7h/0VJ1RpeOa7/XagLPLWL1Ja4IGcnZdiLMQR9kkLFb1zK4Bk
LENE4/tisJWjarKOMX/aExeLeS672QP78YLO8Es5UbdAdBMYgPaVgQFN7cr1NlMcVZlDC8ZFii9B
ze/OJ0oimd36HoE3rIWm2Ky9DTMLXSBjhLZ58XgQZ/l36fLMGOcGZqK3yZvE4EoiGtNa2pitNsIg
lNr0BuY+NVGQfGenv4l+mGW0tQXGcHqAmJeG1sKohO/XvqGbpWyhUct0TWWbpYjsO2O6FsF+2AFl
66Bi3FOSKT0oLeZTop3PxxHiXYqSqn1G+C8p7wLAqbDuE5pOd3MG8nAIeGVztL4AhLM4Dbc9OO+m
Chf/hqkBwrzSQQtQeb73ygjyvPEAY85et6FkvUR3oMoDE9Ct8lIp5m3VLlvQdLNXOz0h0q9I4ee0
Of4bRLfQA8zafSiJ1HZprGyUWordT24N2jbdH9W4Amn4gBxVpB6eqf+qtLXwcUv7I/I+ERwicJtW
a11k2Ek1EVwOVoF6/GhOZg2PNtlUoiLyyl1OTGmGJs2pXfiKnNL6nbXvFFYJTIFgmiMH7Z0txb8N
78BshyBf/Tm2m9xjYKAKnGtZGrao7wWC3bcUeAGT47dZ8Vsbe8Fq7vIy1d68v7LVU/FPmNOsnXPa
yoRbaw4qJ/BAeEjxnCxuq5rNfsNx4d4blS3PjBe0eakcpLX6T7WAjk+pSb2CBPdYc/oLvrJwRlNw
5r8arP5TO7wpm1RsZjud2CSy8pMSws4NTQcYFwEBAh0xitePqlvJyrWUveojGEv9CX7R/5DhHjbk
lywFW4QvNOGYDKT2U4KPfrpBZZnG6CI3g0fvIQe5BwXNjdTn+xg0Nm94WhX/plJYCYOtyyDmf8iv
ki58MvMvogumA9XXEAdV695knNL4Qmpmpamw8/Yn7xMscWgsdPy83OfG5mkPQvCx7Tnu0raJnfX0
ZxkvNx+KVUpuF7eMaUst6m0P+QrE+Lhn4sjvi8uGOq0SE8vHwxlLC+pKqdcOB/vXQqLn6eXjg38Y
2oOKEOlXm5ReRyshsLpfZvv1vhoByaSl2EMIXXafDPGF1RmPPJvwVpbKtiNYidIvXFkOw5Xm3AVc
r/a0TvdLaHmrdNDA5PvWCuzgR2F5nbYg160X43NkDe9VyvepJznZW9MaY4O0NnmquAffKksHwwze
TxBcaCNbn3hdfy39Z+CeDCEwc0EmC+FqAS7YS/sOo38PI/zkmwhe+TWsTUp8+66I5ucOeD9NVbJ+
Gn6dcqYmDfTGy8xvlRcA2vynipo8/L5ZoAaukgNDMS5gKnjtrdGI0KO3bBAijNjiROB5D7C6XwLp
g8PqxFsrsXxcHjwdYzMkTkKIVkGlffzVYMnBCr6TeVnE2zo+n2qvbzbZ2vS/kIJhhwEIyp3H5HS4
rAmfvgfrgV/rv1CP07EkpuvuFE6oEe5SnnOjnZGLZ5L7ZxK0dseKSbXzgI7Jd0NyY9ZzTH/AfToC
shcQQPuRBI6lkTxVBssd1CB2buta60Wcd6kR7d2ozBAQbdKwmKx7ZiXh7+XZkiSIln4Ao1fyG/XC
jLgwafR69TUb/2wodrkgCKYEypyDpKvDw6hwrmD72DxrDnVMjcQJ+ARq+A+Etz2BoSWK7Hxa3cl/
Pg1ndscB+qdbltt6mH6qSjzt009C2rjgJoO9hbG4A4CRcAjPJXJ7MT+VV/eeAHv+iyzf6PuqrJ/h
QSCuVaCFqaTR4VE28G4lsRi1KcCStPeZyaVOE1FEM5uXfhwzC6tS59f7rRCRxj2bR/gQSsJDImOj
g4+AnX9zh++7qPTw2XP7wz6b9/WSgPxgfAL5zOnnVlw0tDCQo9tudrU2DqhPlH5K0IltWyp9POkw
xBJDofkQ3uwoQOY5ANVSpLKzr9+eIDSVJ06jly9OQwGZJSk3a8uUk6yoJkHWQm4yWeqmJb2YntdK
d8XLXJoHfAuGP34vjqoaKBe1UonNBsSU08ZJbayHm3B2yPymv5rqPUHSXME8gW0rr8l+WKtcHq4Q
dZyUHS+XJMHaVzm0IUPdk+TzhF37ElAS8wB1N4TGWbtOIXluFeOmP4QrEnvv5c+MEfq2q1PEZ6Kn
vZ5cAzNMM4qQ7E0fD0I24/datSzpi/3ZjZNyfTa6eY9iRfhsi8VJZSI10bPqiinYs/OfIrZt6LR5
oOKYbN9RXkPamCicYo1doALom0OWLY3XW38/IqzRd4M7FQw+rWJ/RzGUuL3WmradUBVg1xKvnA4U
YA8kCzoOMycLTMN4xQcUJyC2+6H51/HcHf6wZU3o6aOe2ePxEJzcLa3T4/rkTNQjxTMYnXAPCl31
Cluc/ggDEluIGpXxUK729uRxxxSlK0uWYKoWNZPEMR41UfP6+MzyoiVACO9QoD9JrNZQptIhyat+
gcXJNr62/EfjK2GNIpL8hWkTPtPSDVs0P5fUV2vRJioQReDI+fBLM24NjTC78aLczILWn6W6nKeX
MDj72XZdgw3k3YDtDsscU9fLT40BbsPsaZZAHdVNDl+mW24Q+PAa7cn2jBlMBcUL97+bQynaLeJe
Yd76yeYaeiiipN5Lws0ozv4Nivabk6BGZfohW7Ni3q0Cf79JFjndSYwyS85fsGPz377lRXy/gfxD
jGdPD1JBOdz59L+thlfLf2ewDCwZwEIo/cpTnL2YlIhPEbOqAsHKQv0HagR11nbj3VPWgrwUR0dN
nwIzCQtlW/UBRdNd+F5brgGHeIXACVCVKbAnCz+H1FlbhIWClhnU3Fa7q2EM2yLMvmDHHfop5IcY
gtDzSzv07lx/KdTA/K6nVplYLKTYu9dcQOmUwmiUgJnC0rZZ8yweLaHe/ma5+pxIZyjYMa6d89HQ
4MkenZRE6JxyjiHWKB+VYBl+66PHcEcKxcfHUspktsegaGQtbHh6N/jng3DtTqmEFriFYKg70dk9
wqUi0injOp2pe4kaGV+HJgz1SloPlhMXRO5N8S4VFq0SM1XLiESUZvrm89WNdvGuHBKG3LCEmCIH
O5u/wzH3b2D5/g3kInvdS8elLeekGvvdeJ+jEdR4mkAZjdHZK9MypX2NaR5a/xxqqAAKhrLIBNJj
2gzV5qwvTx2OISh8tKZO2p4HGnsD2azfk+rEMD4TLc94JANqz2KA9A64piBujO20MrIUGLY8xhMi
rRa6fseBPtvo+DkGxrORekg9tMETGmspLCvyFt4KX/2dp2zcnHl68TOga+LZPbvplbjcw8zEqySZ
CM/5WlrYW0m7bb/H0JPH5hnwj5UI2+V+iS9VPJjQTgv6uC+E4+JYeUPLk6Q09Ct5igOs8Idzt6zu
IYybJthoJa0bF1w0YxpbgB/KnlbGod//630Sw5yj9uW6EAjJA019MQr8uQpbYYL5IG9IHi9NFbmR
5JR5WNJKjH8OxmC5cevC5EFA6sRKtuVUsuTZZBC6HuOnda3NN94Ge+e4tvD6vfX/Ktv7A6ax+Dnm
m+4UO2y4jxBupL1l5cgtr3pDl0UYK884dVhCT52RESLZtRjpocjIVs8hoDQDOr9WvbwyLhvbIJy2
mDrpe6oXtxCiO0csEd8RcMHwHQnXX002VPAZN4uN7UlU05dXjyGMq8uHejKBHKzg3fsf78gaGVJw
GV7ae9PisYMBoi0NtmQvyeujtYccYJZSKYDn2To9mdCh2EE4YwjIeqcyP2EtFXbzRiRsEK+0NI2x
PEh3qPUmg+T1qrBYMYJiUVqyQ2aODA0HB9d07Nz+1T7fz9jQWCvBLt4/pJzGIXz0ZGw/QYKDP92r
hIC9WYkFbW9z9qjZnlw3oXSKsFQQ+0IyBLe5jq07KGW374zP+BC6VxVzXsMwVeu/+AOF5NmcvUio
YMj1k51LpR5NuvzXvCUTBTkhMf6fH3GkdgVb+jrYeeEP3luy49ZM5OressMWjNElB6B8OWAcEAOD
zFn6WrvY2XlY08DjwHHe8H8AXWix9XIwn9GKdwYgvEKL4qUOJ6THAOTviBhHEUMDlPwk7zwt3dBG
HbnHer3o9Q2GAdrpxBK+GN4saiRYJQ8JGXiwUo6YQeI70ISqVW+66pP5PCkJyO+hno7F3XcZpmSh
w0+N9lP1Wue/4HzrCq+HCAwzyyVULw1rLlgo+YBA5hb46S+Rl9hW97mwAd6ZrsWlRZa157F4ypWh
CRfjahA9KpakINiNFsnP5BXRkIZSwWpS3r3rqyT1n4UfmVQRMNJHkAXsPLkbWnY2j3RDM42kWRM0
5oMQ43nSO0IV/wXaRab1nMbe62FilKkGfoU/DVsj0wtOUx0+VJGreBpCXlIl79gfjknsltcPz+k+
BPMVfzUD4JPxafryZDd9l1hVQINHLsEYhhB0BfpuH1dRP9faKOsoZnjNiSYy/S+8ujtbV5Q7V0KH
BfgdjIhtVTQJ1KdqpzeTP9RHaxipqkTXImHLV4ET1Zj2Ea2INeG+e31mVQRArzJjl4ff5Sj2fSC+
ab/e5bQN8BAOmnh0BO058NHQrMQTPqHEjrDjruF6WO2/85B5zzN6jrcdTUCCp3kAVlaY0vJjg0sJ
/COy/H2LGAD6erUoUqpPHkVNnwVPQ2w9qR5MISHh3pMa/gck6o2O1pWgSy7GyT68gWDWP+VSeysC
EZKjTvrqzbA7wbgtPmr59fssqPsKjHs8lobcZXOj0J82pQ3bHNH4UY/HKw2Yiab3vw7R937CTwi1
pO5hEQ39ShjNl4zxj5bM6RYoSoFJu3YaqfjKoKRj4jYoNAVgZf6JWxwbVAezyEryMXpD6EmhTdwb
+fVcn7ekfPFxtB4YeuBfFUotqcwVrKf08o4OTmL1Jw/T5CkXKJlzToPkkt0rNrIN6M4FgTpgbZUg
QDoDcznQLPoCGcUNNPCuNE/xxD2UADAzRGCwgs9Eui42UvdhYe6bqee5SfJ0VQYxsfcA1R/1zYRJ
bsU4DhzUOYkQOCbKp/FKPbR1kYVpd03UlQADKJtZlYbiYKriyVbw4hxjcQko9RkwqGPv0Jo+Ssq5
PqF8o01slzQOGZynEcwBSafURaU7qSrvjK9+MSYHaRQnIC+l9P3gNPj7t8TDEwnwZnd9ux2/OeJ3
wg7d5poNlCyuW2CcJpA4UEepAicIYpfpZF/kOAKaEdHAb6kN8WNVw8lj31F6DFWKQV5mtpyPdQEF
Z8dkLhfU1eX8clmZuopinx1OBApUvB9tCF1gKnCMAYlEx2mqK74K0zORpdN8C+ujKGnBSb3JIpND
fZL8LljY3NBPLiA9FWZpnCBWKh6WZkH4j+dOBvOpZqgKilzGFfpTVFu0cSgVAKXd22s73u4swEnH
iOFymzzMLYEEie7dHtBh7AiIsj7vR4x/Bmv9UauXGdmmeRacMA+zjVMT2Ox/XsyDykZOHll+b/tt
r1eHAdYUXiggRNzVTNLDAvWblHQLD8jUiwhHlRg1yHas+IftzSzZTI/T8niFuDjvsj1G50Khj73q
DuJV8yGzlcCwzBmU9EiKjmA2LQ7i3d4gFn2/ObRg4Vcn6YNkCd8IYfpr+22uGCQJGZjOgFeYip97
jP08BEwIxdFURp2694vNMpwpZ4l/nnR2Y80yiHTVgH/zl8WxjdcwYgmyWfRGQlqXPUtUxDA+ZSTQ
dRLDRre8lXE2izz8N4jA/TJT7b+gnsAai6baoXJ6BIcDkSUT1e/akoDIKX+MvfByoC6VS5IetzGP
DyiISrUzo73miFvoN1XB2ae2PQ4niaw47O0BLnlolK/WWTb5WJt2w5sOlRoruzB//OSTesqSDI30
bpYHMAbQfimQHZcBTVF52PbxNINMhbDJvke+uHTMYDoktPf9DucNOphVWovgH6IPx6BK0gWTMp31
wAlaeP7xvuknZRac83ug7zr2IH4U0chScqcxBgAjvJ641tzfH8SFpAQhUmJBOHA/DPm3eac5oTlX
N1yKxAa4Irm895BHBT+XRPcv4F3uaOhM1nnjUfkWswJC1NuNa3kagl9wIJPBFG7i++rHHscVT+Tn
QAWkagg2PrMnieN7SiHxBxjeaJsiYv3PmJt3/NpDsu+eILhJ5Tu96VVvZVnejIETFUc8fgxrB8Jq
kkNvycVdmwwECuMF2f6mOZnMsLXZ7ErOm3vuFPfuQmlGUNRvZ2EgK8iVGdgBcHuHUmaas0NIaq9E
L/W+spv0zWVAvm8IzEB7jSkByFK4cZOVTizuk6Qslk7lQtXQAqYvuK1CVgq4IsV5j/cL3C0TLzac
L9Jh9+h2S6FiUFNHZPOR4i6QZG7eu3i+/EiqdCefxWLiMIjgsqayBiYbs/zgK7sdQe1cgez/SBDt
79hAezpOMHUv4cVPrQiQ5k0dNV9DG1vQFOHhaWM1O14Un5R6JC1L9swfLdQ5C7spCrfkNvls1R7P
Y2KvzoB4ORoc0SHG1avg6NxFS6ja6SFbnurvRDYgzdmww+/ttWI/KcFBqLDW5hv5bjFR0XVbLCKv
2BTfwoGaDFP8obv+5It9rrayGNOAq8GrsT0QsjbtJ8YLgPL6MGzaTULH1HQYDKu6ZMfwrF4+Tafc
kgkIl6YbCj4nqSXyGRQV7r5OUWr7JYt/IqIqOlWqBM8xwj/8R7ej3r1wjqDUr7fWpUjRgwGqC4Yx
Bs+EIrEsFYak2ILL0xXUNl+E7aoj7aRXsQVHlMJFSGs8Qqlg/+Lgkrt54izXhtEbSkdvPfaCyGNa
30b//pAOcVS/74SO2NJkz+57I5VG+4Zm1OwffuP6uPn40CJohipFUJuWU1yK2xgTE480nmRk5OEi
wXg+j+akexKHrNj761PuuHiwGOK3aCkVe5C9G/rrHWgE/mzkP5keeWUXXZPwHnmi7RBEFtFEI/1m
IQildNdHK7FDHNI9A9eLNXNsST3TZOhqGuXioDc2TFz+1u5x1BhJU+52swERMzZbL0Oh3hL5bCSs
j63z+Vr8TNBn8LR5rBdN5JC1kffN7/JjhqDADqsLm4FkxnXJNskmgUEKYY4UyykUaXEgfOgk+0BD
wzg4C7e03ji6PbJLbwD4/04Ma22niE2tfFbpIFJ62aopjN2byOzWTq2WJl1HfWX6eaghtjxrzjkC
eDwn5WIaXXZLU7q3K1pC023PUhCLAdPxR9XwlU6czWV7ruL14q40AiQz6k3O5Q9ZlT+Sp9VJCSGT
WTX2h5g4qlbcuy7eta5J2giUE5gLVcMlrc1y2vvAmd6RuZSXUkW95qDIp9LVtxKVtIMjUou0ax3W
o10cj7RRodIxd0asK6p3N8BmhQv2MoFPautPmSz6swdBCqlUREpZ+ebf1pLgpp/jgT7y3y7aYQIx
r1YklHjW+LhZHuY8p7Y4YPN4aMf1FtiF+XRKAnc83NGJDuLsLOiEryn8VUe6FpHg5rCnWnC4CZoZ
7dtUQZPeDTAjI7UN4lGitl0M8HpUlvLgINwY2rxyd96b6R8bf3oM57Pif0yKHp2lwGrCfdLP/JXy
jHJyal9ZC3Qp+s2QwDYs0sPt1HihvVu3ZlxD8Gpi8mhLBAA3F3jW73aljuXd7ET3e3MjxsZBfaS6
wqL+o/D6T4aWHn0xXysXyR98hrfhaz9kW2BCnkkVXFcfoFctrPyKdY0Fezhvr+uGysH1gl9kNfRC
hwR5EMrAS+yeQiAOjjtY3Oir8g1zLPjQ6x0Hr0zLpivANNWld6Z5DeTHjAkwhmhgZhqnj6xbwrMj
dlYDPCEHgXF5kEpzkHge5pUzl0yXXIf+d3XuPS0Px3j+BnTTjlTm50KzQfQfblRXF1WpzIFnIZsg
NiImkLOdkaAvNZbc6BjFJVDec4Je4PQZh/de7IU2jZafaawNyOTNs8muSMx3Y7727543tokRtH6v
c7aEyyd7XyUSUcw43L9FwIRXbv6etf/5lwNsjJc3i+YPJiYdaMO16CqZPxWEZV8JtQqZhqBLKwUQ
GFKYjY0hFzDoaij0gMquG0enHQPrGSrdF/0224cnJyI1ctV5tStvC+UROsfWw/bnfktXksdAXPnr
i+P1pt1uPUKndzFb4B3Vy3wzKFGlEX2dwn0PaZFWVgIQ1wHqEkJ/MdGvnmmacOMmB8NWCniUfZAs
25Iz9oS1BMGV41SW3NXnXlHeiR1smP6wSKSMq3PLVGgSAnMCyulN4ui2AaGQ8HLjwAuwm7ZgyS/e
3WUxd3FXsO+ZJbkfsrWWQSCUg7ph5V9Ydrlvry9b1wzcZzMM2W3gj+O3QLNHWo5zS/E/EgYs3Axc
Moj8AkOgYlSAGiTetBhXVCcnNkfQIFZ2qym4CPb+yOEnxgnNQdAWDpTIpdmdd243CeStnqpceApp
9/fCS3+f5koY240edpgnIHnNghYawZVPBqYYaXGprNA1PnCHXufrht5b9lbJ7sbV8K0Ud2OfU7QP
fEKa5NUQCsVOk32PpHjprCNj3HE/Ltdp7EG8sRhGUlC9jCUcmSjZgsm3Uyc/GKKbN5PuXbiJq3Tp
bfVcuJ8yYP1vxaRdy9rI+kSwdf7U6AG+GN6Qxk12zAty9I9n2dCMbN8pG63CrTcApxBIFgPqvXRM
l3VrdK/ktAh48032wN4e6XJ7/gmT7cdDuo2YXtruWGSZcL7DrQPYjG6kE9OxCHe3eGTcJnhwzJ3v
3HtgWZWi1lJE1sE9IPQ/fPK+CTW6gVBrH4Npa8AHnmfa8PI57HMEEYLWhpHjm6HcneFlWztW4EuP
tKU+c0c/Iyz1jXUAFNK98V2/02GvVHgt/vnKPkIZeYiHvfeKQCv5+yFgDoqLCOq8dCJz8xtiyc9o
Y3Mc4J6wAtERp3Dc+94KhGlb3Z+lWp7IzuSFC/xxJB+ebad3n8FYAB16img5wxY8hWUozzbQc4NZ
+49YyfrW3vF+uoXkHRaGAwMmlevqgwg/hrl9Qm0503k93/wBNl95I2o2s33eXcYPSrXmPV62d1dP
CgaDfJqdmivUixWcwR6auRUTV4j0am9Y0ZMpJm0zoJX4UMV/OFmM/Zjd7s/ZxbtTiLjhZ1pqMIdw
2Nv+xVjQEwd+G/9bLoqgghn/Tra4Y6sbmkXrGW09TDborT85sALmpFL9hMg7UVLVq0X7dnpFoUYx
qLwmz5Z3OV8BdBnQWoPBD94Fyrc8dDLbi49PFwgedxbX9YNeDvwl/nqA2bbXcUK3NdWiPiqFJ1jv
CtfXOIG6q+i+MXEGU+UGjf3jSmb15E9rQZAz5HiTXuh2Jv5k5de2/pruN+gbG4kdwWpJWB0mflOQ
7suWc6p05sqT7dc5bozySKZb5g3zOxPpdfYaa/gwPmhKi0fZGrX80pz/I2I1PFsHFBln7l+oIuxr
tSUM0C2x0xNOLtXIg+1baW6cpALq4EuGRMxwx9ZyQOT8A5MhCNPzKrqSBbSBBvuX3DvoNJuGRiuu
tFd7fBQB0Rr+HfwTTabSqD964foAKtPMkedX6ludhmiFQUfwuotMFQli04o39ld+A2HdDG8rcDrE
nmb8cV1x7r6wW3d5knENDyL6nmal227w9MHhJJ3yF/ZefIKL3weoHTPhCIh6PXlsS8DgquSfxXxl
ZDpOYxtYUvr79avB4mBNgZg42to1nx/j5GsGiMTvRJ2WhSl5yg+2Vlfp9+MRKWsrYA9n/yJqPtbs
tsh1z7xlI5o+minqu65B/13E9m2qnUF7fRehu4luH8mpJgL9jfP5pjJeVBYQe19jXX/RR4zmk2mT
h6pO9lHuHhzTwGRE0pXxm4/wsI7f6tSa2Zw/9i/2PqDeif1HKbNK/X+JZc35btrBlvc9hsWUY7+H
6R83wIvyolRReoYPzlujIEcT/sVJ/4/pDkiKTL5RahgbCuXTv+SvJH5AKEjNZnsnLvIo+aT4E8GT
Dh+4fQqqgNbsE58pWKuFoaaiNRBGFzrg3Rl7arpW9hy71z5Io/KQ3jpMcNhN3jTXZ1l2UBnQKHPG
XDX3bsRgiZ6Mf2nvHMRpeP1lg97lmzwNKzz7KGiJfHMeOI7cE/LTT2lu7znCjAxURwu7FsP437RF
Qf/0foB3X27tvNI/Qzct8L3UfFrr9OVnDwnKvM2DkFw79nXM9arHiYH4+IExO/+olowO2m5t6MRV
iAqLfGW2AYkhbjUU9eAxtIKO8fma9Z6bXavwugRTMEjDOh3p115En7yEqA1fi6XmF+opIFGLfF83
3o66q6O2JsQhc2o/SS3L/ajBRkKudgPZyzItUn0EZBYFRBFsn7JuzGFx48V6xPMcIg/io67YLgv5
RlYDiEGoUUaNa7zUWLn5/IbQbhJD/BMJpPztOzR+J3ZaWGPLFzth9GDTgzy8sVUAmFS6WkZaW94/
OBaNsetBGsmVVXrgu6oMo8x07FL08PHP8x3iU51nD66XwNPUdu5LMobyl/n8nnGzYGXEJeP3La0y
vxWPLafLWsdakM4SZP2FT7LC1Xcp2HzFbiPLrIRdcYAUkOj9+pMD4KcR0JmTk/sg0SA6FjlY9BiR
5OJeE6AbgDi5NMx80x1wMUnVEXHh6kylWqSd2wqHyBDbKSDBdOB0K2IwNMX3vD3s2XGR29dJevOh
jVjPz3fPerfJ7SqDmv13fLXVFH9WLv6UM5DHFAl9SVno8jtolSaXm9zmfM5kJRUm6dTNyTuGxJNY
r+3VUftKaIQSFiQxhVfTCzCRYbpNTOxtgocBBve2dTW3//96oVmvUrJL456P0RirSTyxdQKIg+uI
gR+QmYZ1PkWbZU/0wluWo9qemdAHe+/+WCSqnP9F/wM8lEuQVK0aTFTfYySB8wkEyrbZqFInsIyj
h3zWxvON0rSWfNIp1RqcJIMyDt1PS2DPdoxErLWDuJMiCNJpl6wAUZB93u0XcnD5r07LsTAE9TBH
SOf3pBC3Qd6d2Hrg40iRu+1LTldt3awPu5TFfuPnKb8eljn8Tf3HEEi7fOqHqzOLBL2/fjGF90eD
JvawAwuhoMC3pfI/+4InskZpLw4UItX7wA65m30U0MX01YM2wAiz4XU0HgfdAKqxuOjQ0fCA09De
/fuF1tTZD60oVX5CmuI+t5apnhn/99Etbay2Hun/27LxyUH/iIN4zxCM3ycLYdnq36l8dQCc8LgX
owt+6fNgzFiAzke8/Fptltr4AqC1aHe9SjGBe6u/NL+aQygiQU6yMg2DNK8vKscS+lhxTjSNAlwj
EeUf8IA5lUOw57QA3EoqQaGuxmKgXjVEyKEn2Lg81u5mjFgb6GPzl3grO93gD7M6KknN4+fzacu0
ETIk98gepGRqDqMDrGZM2za8TMSK35AP3X+1UnnyXlPaq96At9hdXcMsb3PsbFjjhcGhmCrD14co
nC4KR1dr9csDYauvtj9r6prEQflU1T2mb7x22HINMKJaEpvEhjK/2pQDT7cU7KPG2kosQl5m3cxg
ZqP3O0IUgBOAGFt1QvZCuhm2psTJw3fy5Nf17N9O/q9IHICRcfl3UUP7EExdEMzvS2CMKRdFsZth
DVMyAoQUhWF5hCpjNdq5aJ6SawdIoTUr1mU6O9ZHj87LWgxTg4xIXhWke8PgQPH66mxatjnvHvjv
72dK43oxB7gh1GL2xWbB9tS16L9c1+JMa5dPOORy2Q0X1Eq6Msl7PZcpCoBvgSNyBNcNEvoPPO8o
7kdwWCrfhPK2hjPTjGj+sWa0wOmGDfrHEXYDbeufOR6986Ky1o2cBpWJBvSYrsB8qEdWpmx9V/l4
DEPv/iqaCPPEAx180oFsXZ1OhiBBZ+WHOYwDHuvQrntkcE6AJkqfzvYsjAvv/gDynOdPFJgjIBIk
BVJ65ykyTybCWvEZOT1lYkD26OtkT7luvzMagmtw1iJ5R1Mf5uCQ+Ux6EgH0E+AFtUkOv/sRaRjj
vfcEURzEaMFc77H0lORz8s3WGJGrw7v5ditfHPzbEGDR4NZBevyAD2X5JsC3jonHjub/vC5v8EHC
+zRz35PfnEeVDdCwSpWa8sPkfPAtuJ2Za9TN/QXe5KCT6w7ruQiBWygBN45uAkhIqi6bnABAPnqw
SoAWxu1AEBGlSJid5tB7WbdfUBSh/nJG1k6qBAPWVlGxqJTKjJGQTcNUHXlO8e6IDpKkyWf0sIG5
c8tgQLIy+WvMQ8PrFUUZKLCzR1fbUhTHjGDiC/h2G5B0lZywTLRSBwkAnh0UxbmwkSylm9stEZyj
goNtqLq1tlIMgYJ5ORkLuY3PNnmQfP7G4zBHFiiRa55xiTe6CcYYGSS1f7bkhckeIiVWcgt8E6uh
cV6abKjg9WLPWtX7bixF+lJ13o4n1c+fpavVTgcgLAquO6d2vEMoJNz1owioIlmvTyA/sTbP+Dhf
sQ/SSISido45qFr4y/0B0mth1vOsaR/oL5V+oGxhQLKhbFQ9GN6bumVvvlq8NVrdjHA0QJlnzTza
3p43ufPFSGATmqW30X2kG+3DhA6R7R20JqlvBEk/q7Q2HN6+EwvL2S6eV1G4Iz/SwklQcLYF+ysg
b/3R2BOK1cet61TZsGrqmsRjBUmyiYyKpP7GgN+xd/e6xbpuDRdZ3DCZNJsaepMkFGajjWSd+RUS
WAcKyog+SP4jHi8agdcu6bzTKDWsj/746VBzq2SHM1OLmslJ+b4kKAXN1OTC7VcgXd/uTKEyBLvy
1WEr0INsn8apzKJTzscKjOq9la158A4cTXIDheutMNGyCQbxJgonqphVVQAUpHO0opAuvFIuDJ8R
vBL8ooFheEkf7xsbtebz4gV/9VUqWK2d6RXbcyC5HAEBzvUqm1LSscLVY/TFEkrLb+NlVXZJa4um
6gMRVEBp3EnrFz8mpw3AWPVeP0Nv1e4nf9lrsfNonKHuYZDurUsPgMV95y6mSCXqo0Infxixl9V7
hfn3vfOmeUnoqOKhMP093NprEbMF20V+8/x4SUpD146uqXgfqifBW/N0U0SQUrKZIP9itarDvngP
2xIAxh5Kb8KUe0LZCdKsWZttrbSYe2DSfVIZ6RFJdaqgWhtLKpTj5kopFOfmUUtyXUlBEBETVNpF
L5DclBw30AsBoqmlkIyy9zqlHQB/irp5jfFL4ZcH9SO3/6Yt1WAMHJWEwy67lt/zAA1TEFx+GuXf
ki7ChzfVuW/uWK99SddH9IynkkWJMEuoaz+KJxBaBAQ9CZO6KQAJ58jH3g8VH9QnJmCUb8i9R07i
pVgCfXpmIVeNbvfIe/KCTcp7FJkhtwm4mYffpO8s8Nq43I3weAW0Y/UArMDQXa0pmEarUi51UyS2
59/djKiHpg8zQ9pOICq74VCi5hz/BtKuWOWJ/3PQWw5LfmtsQl0qQmyH+CiuKDOpXcomYvDg5XDH
94pcSZUB8tUtSqwSljmSQsRdOsvbOatTIcZCB/y0HK2e1a98yWSmYutYiuCAWj7U5D2haxreiD+o
0E+bu45wH8UtNNlKtEsAWZWHl+drfZeM70oLSVSfZBcVF3f9QUxM3TIgxzrcNwtrYoenl0o/O5I6
VoAoJZiT4+nUaYtLjqeNOhZ4qKavodAnuEDSqvXON+L1GavrbBIok3LygzVYX/YWiLwOOBB2a+ZR
3e+Ku7RoxdXU8ZIemnluPtQSrr9wAYs87lz8+or2HJanimuPqYTbqOoRO0OUOKITZ1y9NAPLQrUa
J0J1R7YS4oxUhHMQ9tvBlVaZ2tmuXIRw9UtIOoQHI4u7NrYPuOLuNN49D5qmJBiOsHQohi9yT5kI
OBXpFGRI8i389FdJqEPWp5fK4Lr8d6oEWJTfW1Mqdt2UGt7xeqVz85JysfvDV0tWRW04MyLrbY92
h2aN/U3jVehUtplNwE9kVL3J57Z8UulEocbEO6/P4JOKVvjvn/SGgiN8qP3TrWI/fak6cg1fIO5t
U3sbMwHpJXND0/6cY5l59drTWotDwLxLlr6m7VzkEkEJN6StzUEmUAh3N2tch2rTnR5n3aN/SkWb
0pVcdhgx/GTz4Z3Xjau57OMQ/jtwDt7fiaFreZ2wBlq1qX5VUTXRVgeuiJZBb732XolUqr7bP2DG
cIDX3CmXV/XVLSmXCabpf8IsNV18ZhqJu56A+vl2i9eCpknG/DJXITj/Ug60Bd2jo1d5JnSVQenz
cLKZl5FGve7N8uGEgxeOTxNSukz/PznKKXAMu8r9aWoKcPfsaid44Wsd/38UjfdZ49QZn4xEwQIA
UPZ8zbhLWUYlEIrqs8mZOoxqp0/BHW7XNmnayndDaCwc/pDUvxwhaDpj73VQZDcNnshB6jRSPM5a
y5lfAmEusBPKM7sqgwlM3rvbh34RWERNMgeEJ1ZgoXglipS7BoIO11ANebzggYKTLz2Y3uznwxv5
7abB1Z1BPMmgU1h2/Q8Ce55xhCZvxAlfFjrctxkq8dbKm3oBVRYRBIyL/c+AQp5bSE80LSfbbTnM
sKSyr+K2KIW+EFuZAREcp0irQqXGOQ3pF2aNp9X2y75eBeHb4292WxwQteQQ2Iv0iBQ0+ALS8ltH
lGfcGL8N8Xdahgul+fW/mMLVftuQIOiwPUhNO9zfl+d7e1X+StEyhmAlDL1uLYGeSgtwQvvd2r+m
mB3f7wVc0xxgh44To+BTIryuWJRt374HLPcwqOilsvlBLgqPf3mEiWSId/2U0zN8C0yMPMuzBkoQ
DgMsqLPQTu8sK6g68Z6BXGDLcRchg6eox7AoiRv9h8/JYzzP96FqpAMKgu6H8MlBuOLM0r3CvEKS
5hqZzwjSgZyA1tMdPIU81mdHnvpL+dJB8PVHAKL5tJ3V7hnO3wMZfcdixaAMyB8fTmzEO9Ml5bsP
TIyQxPlxzeSXOsElaP+pC4iAYbUPbMng9y1kWZ2wH6Tliikwdo7Hgk8q1/qzzNatxUhZjgNcUmyv
YRxn78HmNrnlWpFo9n+kvesydD8dz+Wh5VntsRb18BErvVhU2hmjzVM4khC8ShDZxgMGZJMF+b0l
dBKHfIpCclXmduuBhSB/c2Q1CyYIRQWXueWe5C12l026ZVP4H3pNdzMEDur7V7dG0HbnUYE0Niyh
tjz6gQGW5NmJ4XcZQUS6f0TDqYvqbjM/WtFbxd1000Q+nkuKW2yIQD4OzwK1bUXamggK4Ovkx/09
uwjoBFWRWPNwwDtKQxm0G0gXSxxHe3zT+YNZb60Ir1Z95jX9keSJfe2ENngI7p8mjF0iWJjpj0d3
lw8pdpYzsTAW5jF1QzUKRGh95pKEzx8d7UR0CFKwJkn0GWuBR6p897lFJEk9yUtMSulE1KcfAZSA
QVgZtQU5Km4dElJptwzlLZuq4QDGFePBO2qM8QWkPkdWH+KVFJo9dTo51q+SHXPKBhlcX/q+jqqi
K7utjCDq2P8Q5SHlqcl9LVxOj2nzjRR88eePaC/asB7efr/tHFvsk8OiHIaHwNogOXZPglVRPI91
qEyElMbsON9+Ryr53gh6MlNtG5wE38X/4ror45Goy04ABF95fAoYrKrV5Bt+dMM3xeHCm7+/IwUz
l55hbwwqsdDASAsaGRhi8PXEm+r1JzcVSbsbI5Upx33A6jzSLgXTjQsySRJanjFd+VubRxRbbWJN
etBkWVEWkmP+dbaK95VMEHMvN5LsLx4NKuNt07JLifhhnG07TWKhgWWWv4kXLLyS9M9ufI7wiDND
RRqGvyopQJUbyr1K52Xexxap4m3llkPtbP0p80dAbofH0JR54cTt4WS3hELprNGdVBxyJBHXPDuO
uCA0/FDDVGpb85sR7x24h95ORTRyR8lg9ogYS3uxgeN0G4g0cUgXVTpx1UGyOYsiWQJ4pNbjmpzo
iK5qZ19Tn47YWXaegE+BfcL8LMQ+YwRASEuudedJ9T8J2ihPYjvQi3zBfcaEcB1YphlQ1sruV92u
gC74w9Ci4059er77mrIggc5XGQIg0p2L6XXUGlYvsRi0t7bdt2yTol9uixYKdUdEbdIMOTBcah84
g+LkZt84WHPrp3J2W9Vhc4pBMA8h2TfJtIr+Ya5CR5ghbcBOBdGF9yI6KUH0FTS8c85NTxDLZqe2
If1HQlCBmMCJCWtLHLbRmKmQ04GZ6AE3+gL9PpTYCl1vNIcX7x4HYpaNZF6FeYzTx9FOH7BX9L/g
otw7EPFvHazXFvD2Mee8Vfxc7BlbOIqZSuqXf5UVGdX5DxfSk7EGviQnr36VpXytQbzAJMUssaXf
/sdXOUxH4DtNfj5+YHau2V9u+3xv214IBpXeEb1xWR/zRtKBDHX/G+x+DKwoDye1WpwHEfnwEyBt
WHasBcBf/9uPQDLFt96t0b3BX53JBu/ByXVhF4wpIAsIMTG86TFJNawsb2ueJW4vUXvVzcXaxZmE
4LyVWus3fcrkLEE3qGJhQtvSoZ9CTbgsAS4DK/TVdL6gCVQRZUqtaIyARnOrhEagK+4vSvqaGrfv
KQj2nU+74G2O2z5P7F7ia3MkMnlCk19MFc6OS6+nqt9Gn/t20pQtnnWgCeU/tUOB8PnaPHx+Vcai
ssz1cpjqbTw+Ersvy6+I61RSCaaQQ9pZUT5rXG/v0b9ubHcd9tzh3RTdV7DDm31QixT3JHEwaoZx
6Nh6Ur+cxmB5IRk0D/q2+Z5IWmzfyRipZlY+SES+OLBX30nvjftdmephakEVl9MCV8ksRZ5a+jKd
frn/x56zZj3YjY68otE74taTScwizUqv3zwb2pYEr69D9LKxM2lz0cpsapEl6w49j4Of1BVX0DDE
lrddFZ+LlbX2sn1JJxD7J48jMNqq6BxQzrMgj0QGAZLaUbM0dfdV4ktT/SLyAgicVZXiNXHfZhrU
15thfMb2OWfTfPcke+Szf4y1yZiKxVLIadg6+NC3yQGrZUtQOfI1NUN5IAVEJQPkLUN88k7Jr+Gx
Rlpvy57VnDdDez/8WhIWuHv1v9TjNFZTEv2hYFAglsX2H6upzbLjIJeoOva5sCtDuHuVAFatwO54
mSb1HYrfG7sCZ2/0gBY/j3Ckz8HUnWvIWmrCWfySsZnu5XbU5pcEB5l3Z7ygN4nwH66SJvzk/TQA
VBfE2d3K11uaCMoar8GRJw1xNFfSH4ftoyn4tChgXYGixQ8H0swD8hZXG4ryA00cRctOtlBgZFM8
9A7sKP7aLnc0Gzkx4rdLpc0BMkpUkg7cuPchU/fjlYWs/JCyFdchYEcwqeF3ZMaEliQRqPxbBNU6
8Ad/sQOLpwEsNmzCUmOaCq6q2qL1SwlsK2lq5R75/ZFhKzJYAy6mh8coRehuZBrMgTij3U+H1DiC
CLdh8Z7kuoTWYfcIrNzzCxDDlgOyzdndeJq80/K8zhlN5Zdu10/g0u5gk+RhnwZdDfW0qSV3jBY1
bClQ+wXP65NJjz5enTilY0o52N+Fs3WMqkPhSuJcyt10cdcZH61LSYtOCbjzgxx9cZtKwWRdUnos
8r0D4E0W/fU5N9hMq4b/lkZRO1X/vPOLlSOJh/1X4aanfW7/cRhGYkuynqNgMDRxxbb3gSygoYOX
cEoOkpkCemYgjuoYQbsI49zFMC7O6/VyPefSiwjTUP0a6zfhHpKUmoBb64BPHpu7gs8hcFckmeTW
tVG5pZ3HyRIYeDT88Y7VMFe6ohMmQrRxSGAdIk0Th8JydPro2LBmITLwAMx3x2Zu0CPbMAEEaGn4
TcBGS8t05J9M2/GE22XLj+TIDctnts2994CucPRG0qqUJskVKIQz4b9E9SleIsJObDhkbayYquE1
V9RKpGWzBARZftXhsZq8PyxPZHSpxlpqYbsDIeuuq9kci6Xwdaw0visSZSfsixlxO1xe8YbxEyEA
+ITpy4ifuHyTe5K53937KbeVOULyjw21DVMTxY6BJFEdJWooTK0q3pNHvpPNMtPvo3uq1iRLS4HN
K/ZrL48Xa4My8Sa9bKMNc31irk/plsE6xTY0Ym8aougYUMociqGVzMZvVJ4VmjrJWaPB5y/3Yb0S
zrcjIU3xPEZ9hupvzJmD58N8miA7yofiYEDXSExzdRzuZUjsIlWHSyda+gfuX7LXWTu2SwMTNLKb
PqYRV2KfyJlhrR/D2V4ife9LdjWvKELU7M4nYEi21R8hYuQoVxZ+RJPhb7Ela/b/sMjmQY0Bo5+x
XgfG2Sa4Bm/xkh+KNUjFcYWNsBu4MIK+1CucOLGxW/yVR8Mmd8NisDQ/rLqJNrd22Ik2Sn+vuAvI
U8+4nVK88dDgjRrScMVx22Mrobut5ONpGU8b0xoSe1AaQuMDRXFPCHTnj/iRtYvsbadktqjG/nyv
6klfnOFeMOLMnrU1pSpDRkLH0ZLv1Zokh8BFPGYE8bXD+/ji9AQTTEhW1iVlaWd1Ipv1YncbC1PQ
ZL3Yv02n+wgQ9gJw0JFGplkiNPbBLh+8SeWWHHfjEfKdW+M9PhGWHod9mYLGiyQ0Sli4HBZmFTcj
yrISsd3FnfgNLfbBeidj8+Pun7Xf2Z3MwyNbKx64agQmLpOD3YuOUczh9AavkXiFYP254a1fRmhO
Kd8yaRNtTm/nFf1j5O1Rbn6Fv5jWvEBYsVZ12BD/AREPlI+vzhKxSc9FKEXvlSA4dxBzwx+z9VN6
SOReQ4U///q8ezEuDbddBqd9EDE9777xUGkZcw8SHOgApYWcUoUlIT4+7sCVkPEjzH+6GxlkJTL+
/nbFNAOrmD0NY3XKLMG7hm2Tg6Q0agnejnlmCSBDj677h9ulcjKYcnAUlSQ5KXlO09/lKENplYtV
1DgRalroPAz+Y+uD+kZbNCkOadzbWf3KovYddrbgH29mH12nFrN8fpAjeAV9jq2WU/TaXMsmwam0
3XWY7y91/12D7BbOotFKgmJOR1n7Vt8OZ2i+qY6e3WlpP8tk68ukJaOxRSRGpWwwQ8ruvGuiUzsF
NQ29FgQkU57/PzEoJ9xch23996Jkr0NhI54TgSvYeo4rAjGqfKaUYZumAHwwzAlazOJNxXcM6Rgy
hO+A832T+FEnPVkUB5/qEGZdMfnQA/+dHi5cA9Ex3SJq2ZMgTWjFQzTGHpRWA6QYRoHKL14XsvhJ
YJvrcQhbN5QSWcAgrUWobB700PX+k3krcIO3IM1aCox/3T0mlgrYR/f9SJxezZSqUdsnKH9AlBC3
ep0XfWplQazCMvgYMxqUP8zaz/zGriz1rke4SqTdzYRE27xdtUEPkD/40P+qwSaDfVRGUwr+Rn6c
TWt7uErSCGm+mKytKrbP2OvPjLVMF4hkg8+mRVFIsiHWqsMPizyTZgKA1RyG+8DSsWNdxAX8Z6YC
uK/f0PgUMG2cdTd11zRY/TR1XKI+2Zv+RCTBaM4pOZR+SOPCSuavCrifvlDbJGtgnKsMimYbD8Xx
g8dQusSSW/RI9LFUPYUCCvNyeFDTJiuvomeK2vVu51E72cBjtMN1+nAi1EVpy//jcP7onGgspFcn
tPoSI1ahYyo/huVUCPQz3BnUxx56kWn+PnXuTSf8ckP6r00C6K76QiKE0cW9n9zFFNEzqdpk0MFv
wekgX953aWF8sfj1vw3i1HxlVBRSgv9W0vaA4sroPMMtaic+WNzzQNBIJUHlttD+yydAYOKwsb3p
0Ti5oKcUIyDQmi3eSuTGMr81xG5V3WFhNa6UcINJFhwt+E216u4x52I+Kc4SVDgKODSfeWeka6ul
XSZzOdXetNzWosVu5a9GZSeosDwl1pNi7CXC6nXF/QhRiGJify4SzkvK2FeEq4qn4RExGWLucoEA
2us32b7Ny6VJ/gu6/hKypdB70vNXe5BtPuwiCwuHrJ2OZlDPt9uT6Rp6ngHMOPUaZbiUTIuki24o
Wrn43yzpOogAUCV/V43V/oRzxO3ubYggdGOqionRzfCkho6ZwwEZafKGBWyYbQaMWeGlXg1cxFkh
W535bveZt5SBUn7SXVUQtrPk8Ts+BoOyhYOw8WnjlOlBiAYOL+qYkHHQwEYHiWLzprjwlfDzEyU3
tU0OOYzgoDF3vEwzxnN6yc8Wqexdqh1tFyA7lqLWvzEC335fliNU0FRb9Z4Fpficl8u4K1wI6gJO
GawAdJfv7m++gYHVUXkb92WXmtA/Kv/bIxheEaylHTzqkqiLKYsuFl/pEptZ+fDloAAE0//pnm9p
cl/akq6xVN2SpEA+Qt5kZIHyzey9+hjYia6crfBmfnxnFJ7hMb/oskg7xfHtZAGX5OP1nMHQfuFe
mOFX1e6LKipKng/aEk6oBTjXkvyT1ybHK07bWDr3oXRWwdHvf7+9L1ou+ovxXEUw/Cu6TCjnGxD4
FyjclO/uBctv0pXRfhmv7dvHBrmPjw8vLh41t8oAcksxVoAFdb4F5OTZ7Zd/fNHD8EYaebBiJn8d
tN/gyGIyJAudGO5FtKLmLjh2ut/FH5YF20/b1bzQzgFETDV1K2bQ+spmctHd+Ji/+vmTkj7c9/wz
PM6vfzpqaF/1dXf70zVvIqThEDc9DcgX2F/XHaGVy0HT1tEjHf47+PRekqtd7+AXZvogWnQyuUCq
irxhYy6rNCeJSrzThSYw/xvmG4v90c3X9YYlQHzREOz2x9BhLIJnBOB2a/RDW3HUyy/JI/kKT34/
EWJUMuMOoVmtnBfaSapE5rsmIF7v/Ziabii4wozpZOemPWRQynwT5LpLTADpA1vAiVQfB5whY4xA
XlDjyN35tmEfeiWruu3r5sP6O9sYLwvRKn4pwcgGCNLX2D3gvcSd4qZaX9nTf1aYevtlwtx87rh8
INv+RG0DvRjDNY7dAGNX6mYpboJuhJQN7c9ZdApp+0v/QWrbDXw93FFMQwmraRekLBgEWb9SeHTW
VRqwiV2ukHcxSvruzgsW2DZ6m1IggIWSSj2y5qs0+guouRJmTCPdk/tR1OSF3cDAIBoN1kjY9Xr0
jaDBlLjhqfNOKvWLy8N8mDdebghnMXbXubJDRLnFTo7mG5j78wMHSDmukgJ3bDYlPegIcuBQ8Rx1
Ub2JjoncKVLSKM/s4KcRn6DqpyOc23NY6WrdAol93YzyFS17sv4ozFzdaRFhdK6OBh3Q8BUKr9SB
BngFspQvkRkz+WqCaX3LFvYkkBD4bEwEimBB5k3+bdIa+MLg+3jy2trAUywR44bZOqUOwtZWR5Y8
ig3uyKNHk/1/WQ+yKOoHi+RjnXdK4TJ6APJlz7yKUxxmh6xN71ei89XChZbD1veWf4QC7/UC3cTB
zIg7KbX+kjwHXJUE7qiIelxvbkKXDTcXo/gLr2o9G9/7+CuG4IYZSs0NekzkU4UnW3h/fMu0a776
Zt0UXFRc3q7cKuCE4ENPUEQhFqQn0ULuwn3Fpjy/1QuYqj02fZptV6j9i5SBZXfNSLPGe+g1IAoT
OBCMC06muTP1CMY/sRaUc15UuzOonzBqAu1YOG+cleZY8mDyI7Hmt9zaOIrIiDXoJFGmGUBIuPJg
30Mv+7gz70hYQXq2qqx0Sfzg4peFLHQSPl9xffTyw6RsjVS9fAiNRIEA/Trb49jQTlAANGbjPJpt
MJZPeTcj/lXrpaGUa6NSxoO9siKbaFW0UbbjiJ/PnpNEQsaMtCXPGM51sttHA1RIuFjLFf0NmvSy
7ZYL0gBBJdWpuaL9qdSFvt9A1kBXrIl6fCvZ11GTgxjIjGNjWVc+3Q0i5DfAKpSDkjSMjNp0uMr4
CAEVdL4AjQKWIoIt5NYhIB32uvBeiR5930xN1hEOyk9p2NsPDv3oPJ5EKp3ncV5o0IDvDpfaL89l
6KIM1UhPCAvOeTXT6lQ3BvZcLqbJGABK6e9e18Bxpn/dSasrFYyBxRRnUfASP6wKzqK+nd+5ruYp
AUszwa9OXUBJgC6ICnaGc6cpwKgJ9UcqNj9ZFHGUi8PrAWcA82EkaYEheuEN9LufRveqUMI/PcAI
Dv9dFSbeooeNCUDD/7+GwNfYvC7QUpIQuAo2S6hbnr1Id4xogYKP4re3Unltbu8d+niACIuhxgDq
bm++tdmL+XC/alZ8fRP1xs2jUPIRVSBty78x6rfYJykb+F/3LfSzpThIqTOerX5Oui7F8appKBqN
it4AuFG+cq8xSgV8kyzWzPF0//M4YXioNpRQnqWoMYP3xum0AXG8ycUlfGIrAWODhZdo5armERKU
uqO41u/Yc3Gfs/N2x9XnqgGNwedjxE0LK7OlDRPwavc38t6ZDPs0BS/sATrErzWH8eKh44AZCrWU
bneIwwIyv5uUapFXYFaif/+E+QbEJu6plOGn5/ffkwxGSVDnClNY+S3977AyhZpDvwRq7t/aTt0D
n4q7nkpM8Yps4RAputcW0FUuto6SBfiqNykSaaZNnVTTxkSwVYXVpWjT76iaob5hnQt1d3qXeBlL
VurjyfiVSQ4SVqVmjKClB8cjkZ6g0+RtML/0dtauOOGdPtI3LhRfSOmhNdeUj+7wloujeQ7ISFUX
fbQAQUxN/7N+8OoRN0D441SCcSrSc9Wxu4A0UE539yRyKou3GWte96zb7HMvi/kzURKXUqQBrG/L
2oVfMQ2rvVORX74kLVGIDrrWQNQ370JtQnrUlXnsgsIGA8chzimzuCo6BbXIdsDZStDoD5yOZ4IP
vBmtPEg/PSERuGrydqC8Ci55NrojhkPaqN+H4hYWon3eLmdUbyWWNDBuQ2rHBLdiTU+YKnlH3xIA
LnmcVXzH9FatqTnJwbP/fD57LzaPDc9Ok5gyFQba0wjkNEjpRlhR22dosAb0og37ce12CGNDnbMV
wC3B0+Mhfkyb49l2phk1Pa7LOq3ZCxdsm7pKZA88JTQNGWsDVDf1c4IShAHmUYviclE3c7ux/vrF
o2EznQltNIkD1fglsy1N6ItftUhwgSAccqQmLZXfn/ncijeW3YdkKtsygjrUpadqEUS+rlhscFUP
DILl5AxjU8cmzEw/4q2PPe5Bts4eRDT0J/vFRYFZH4pd7wvf1cruzEvdciub5Sef6IAGhhei3Yf3
zgG0U5AdnnedxVEQ2/ebgduKHVw+q26eYnC0+gVMjYkSbvVco1J/NQ5wZ61TNemTiFPEkS4+UP+R
CqCJosGwjZkRcgskkR0gNoE4rGJ9CElCxzr6VAN1KU/YiPZ+PyNp40hQEZDYBkvm4/oPOYn9LiUm
WXqy3rzsA2b+HrdOs4QKXJ2jUKGmwY18D5OmP0kf548vzLQzLKvHwM23b6MRvhU4mWW6Lo3HSLGU
Fkl1WDkmFxr+uZOaXEjpDTYS6hKeZtP2tc7Iq2arGv+5YJzLLLnXtLVJbU4U/MojpMGWt2eSX/pF
gG+EOZd2sozN0YbZ7L0s/p3BPOAFGYyQo+zVxiQ1kQGVDiiFV19TJlrjUcfJj8qEYBVyFolb47qG
8Yc2IjE0hda2Yl3LfGTX7lPifNWw+lOufdyeAjJPZetrWboytHZmMotApGAm3XsFQRF/yi4PK0RS
LWuGxv3cT4E2Xqq4T1RM2Py0GCduaiXTYQGdmdPknJSxvDTwxFQdyVV/oHg0j0zm3HYPRR8FhTOj
l4fQEW9JHvMs6fdEIZfwN2pc12/2YdC5wuMDfmCf98OgL0SfAxcXIYvvKJm+yNqKqL67z+Ljr/H/
d5FCfFskwbFH8HZLQIRB5bCC+U3/QFUJH7/L7rXMc0+Mm9rtN7mSDygOXQ4CPiOdw9Tn0gJw5MHj
yNc29m2OCxBd+ErWG+CK7gacB7CQdVcoxTAjxaXH8amAEv9YekArcOd98Zb6InZMnVdoTFORUxaY
qZKhfJqcYEb35Fj1p5vPGOuyRe6QaWZpnz+7Zrq5PfYIUBHYYJ4yE0rctqW2bteDVLVT/8R7BYFc
9m93rPHsy/79tcMyZL2d9hdt+gj4zWtJ3MXH84Nh2CNiegECrjS9OLZrHaN+XSVOgRHmmPfN1Mta
BZijocVNy/23tV6v7gyO9+jV5U6J7COlW+RAOE+2WjS5w7xuONWGXe87iNFWGm8m5KfPzybF6TA5
k6mjdp9lRSnKn0inmR84RkkJHt5QQEScgywfFxBVXIsBbaa+HvGtYYJK2XJFu+W6HJOuTdM2WtUC
UiSZoRHlqgVjmLyK0Z64TKlwGRHhzVw4+VtRepuQZnqZOeNrMvO/6OeD45msiw0VAj/btJ5o6riL
3oEw52hlbW6ppJeQqjYsw7WG3CmlcwGydqWCuNq2wi2ofq0Sub7xvxzGt7H7fF8XLnuGTN4RPuPK
ylq1d+4FVohehynxxv90KPCvcC4cr0yjQm7Dqm8QhYBshpsBqJFoXhjPQ5/1n2fhWX1vFX8D3vSe
iXq7PnBemFBSBgfB4Q/QfxVw+y4uwxrKq718Hlo1VNtTgwU6wpV7k9rKnRarYLS/bArpRno/B3sS
qVDU0nYTyp7eV+VLGLPyyT34+2b8dj2PgGdNZ9ertWch9YYAJxB87pkLgjbYYXJMURuh47TlBG8E
rSOOSDcEgRxtilLqNrDl0rAXF5I8tq56X/YsH017ntaluO9kxwPRldRiLhEaztPzjsPjVpxXkCXQ
m+xdTkFuuvZON8x/uupY7tF9PAGEfDjJ0ScT8PiWiAuOK7tPh6AkG0gO3pmSv1s6YVh8cx/SSqbT
06YU0FhwfC7E/aiGehOPKR40PgxmUd1ifCiJRV/hvIH6sEMhTg/DZcldjo0sqWd+7T/RbHNmLyyN
pI3cLIdX9d1MIhErcQAeYNtkYKLIX83fiMASR4i5kPszjCNwJd0vUO2Gk4QQGXM1ad3aHXLsd1CB
vvlz5U1leZIHPii6VhY5FKfBluHHKaDxcyZCG51SLFJ6zii/7CLB+QcOB0QE+gnzTSYUvy8+aTxJ
nmJHwNAkwHQYuNd6xWc65nq1otsbS3ZtHvTHJBLFFGX6i0u2xQ/tQv6xaV8N1BrwPKXSjmXSLQwD
DN5hnErJ/9DlLgJd7WbG4/iDnxj3yIdoIwc92AyS6mmxXlrwZYgoEF+il/2JRjquaWaurJecOB81
/bWLoqZ/Wz1GoBpLGggEPt91pYJ15cpu1NxLg5OLEEONER5f58QkCoz8YWE/qVPkCBY5iIwInuOQ
BA/vQ/DTq4sXV5G7AZLxWcQSrIQi0f8XpgOMJQn29thDenDMhBlYJy/QKjiMR/gqyoxbkispiBTJ
RMHVoH1TXbze0CUNnpCywtSxyp+MRZEoO7YzyKTq7QQwwvKupcOVYFFA2MCkffT7BYHCEhCe3Apt
hjMf3nVGEpRBE0WibOG2B73Yfmg4bxgawTH2hQuzpuuUlmuQnwkzj9T4cF7C1W3hg/5tJNrsSIlo
o3sTlAbonTmxA6MQEAct+BDKYy4A611y5Prc8BLtCoG0MUrwtN1ljdkSKyzDunAwSbgbnAk5ZeCD
RPb5Kmd0+pzEGzBtJC8sTz+MLAJl6cnP2Wc7TnUX/iIYthfap7cBa5NTU+wD+nfoAQQ0heu5W9tC
5dHUBEWb60fKViifdt1UXKPW1W95D1qa8xlNAbCf2kQ+wsA7vfntfO3M+IUeyrcX9xXNsmtPHkd1
H/6RPJE9ijNBmBLPYchqhTfRACz/SeBBw1DcbXcK4Bi+XWuwXrf6N9JwBZzUYI4Ka3Ac7l7M9sGY
McOtlijC+5uYyuPdTwvt9dBwglM3NsVBqKBRl7VTeAQJE/Go7C5Dj3w23pbJAmAZjCBnH8/CE49w
J3AMj6P4jWLTRLMc50KXYOtePErfeAY2fv4z1Pdsle7dFfdEbUGJUhDGIaWYmB1L6nEIkf0BMfE4
Wktm/KMql8C4dLpovfpHBrA5+ShAcmyhu2t0LJltbV6ETViKX+eZtukZ3Ab2sdgrhfp1J/fLf4JA
VlP9zAxE9FCbj8KzjRZ5v1MLR8LZXe1m9lnvGDh2qHAzLfGmzgceIXx2BTk3sl/n+6trl5sYzSSN
a0henIv57gxqMpemCUm1ros8hn45asRmmTHNHnqLbFPa17WkftSDYIG9zptia0DC+AZ5wZriWwdo
ZWeFO/ls30FS3rXF5GzvKiuL4CFXL4N9s0gCNQI5HVW6WyJBWKz8FPnB+Xk+Ebmt7uoQFC5eTkcy
qSnfljfWhtJXFpWn/K+VPZyybz7Z6hQNUDXXEpn6pe090Npqys/AP/yMq6kritoFaT0kKtzg/xvv
t1vEj25N3DPgv/IQeTnrbgBEuqX3Fp3bRRi9nN35QqKz3RcgfwHIOJ/ijpjq9s+AlfcCQOMGKaw5
V+XuV4zg2lTBS236a3ErI7LDSQAqDwsZX53iKaJk/3bEuiw4MidBRZIPrSjttmkptSVeuE8zGqlW
5Vf0VLgc3USNdbyJAGByHLMFvZ58umAu54OMLOnePbSNFZtKN+xjdyNMIAgKVskdV3SX4mwvNzFm
7N6O1chEIvoToxwCzW4totY9DGojwsiFvzK5dFGS3H1T3ykcdh6LeFJmlLg1a1po5JbzVnq5pERL
pRswL8+zKwPj9R/3l5HoZ6kO1xoffT07Fs3e1FahP8VxzWkUERMlnFzi9PRzc7622mob00PNblYm
+PBvPuFu+i/lvHc7XxOyuXnHsCISKmP5e9I8k4RCeHyMfkF2NNH58CIPRyPL3YhsuYMWIv9yx/Qx
XI0WJTVf/FTDcwGtgbTxtYOUfHl86IM35PQ0nqfG7iWD7Xn3pYXNwJ4QdBmclrY6mckTqOmEHbl/
Heqh/XaJ9D3EKNHHT+DB7aX/G3qXGLnFQsON4MBjOlOAMSvW8/QeUcWBRVbygWz7AvQMXKNcrpLX
DbFcwqzBvqQ0wpLDjRZuEuuqltn0SyN+a1Q4/qI2L/XUzXW0shNMvT+GbDEQW/Xa7jL5h5FBsJc1
GMPHcWO/s3F5URtlFle23kIAGxJ81ehM7cWAnE3mb+CHYv0Hk4y7YlcJcjPq1UJDbq8W2s+8LzPR
qM8es3skD8kfEsGsnRUmzHbECvxwx7IoBJWNLyC4Fd+xSDeHEqYlmXqRDfcL63JN+IquhNXG2Aac
tKbOfRD9PBBPjyXuvEQIA7d0rstWn/R2fvkjJpw5SsFETfrB3YM8etEkYwACAde8cuLzFYZusRYL
OmrN3z/NwCUUecCD2i0pTAq9XE+CtFrvyDvU+euWXgvzLfK7Gtxtj2GMgFPMDUCvoTMRhnE3ISfK
6XWcOQh38osPNWuqL2TgTMw1G3mztPW9LXQyu8O6LJp4cQDzzuWZVVjsnfzyhQmf35t10zIf+NjP
la62fzbjd6oJDZHA6Ec2M/D8vgPsS7P4QoNjzi5NNqSSUHff6VxNE426f8v6D6wx2OaAGtAqkgg9
4E4K6r6lsj7GWp9wzfOZl232QlVArL7GWYxlG2eHVWzvjiyQS4fvocPltaEdTvEMjaECybdBAede
IYikWfQaksNM0O3gQ8NR9MUe8YK0bxDLtl89V4JP+qDejUUY7f4mx730F5Czsg+tUbpkl9kSB6+X
IVBOInQ+U5xgBX8tXQ9vOarNOtrta4+miZf1WUAq5y72TmPs52QKZsfJYGAW6M0WWk3Nma2ySIWN
OFh6ZnRV88oSfnyVXE7jk023Isb+Jw1yc1ZOMfrNyxWMGTZUSR4tDz2K8OAVTxyjsotQfBqH1AgN
LAxuzFTxN4PDJMyP4o7d4B7oWCbMUPOIF05k3/sN9umxSrYZTGWw9JXqThia4rZd7PSBOnSHwyfc
Xf15mWDke+P5f8A/Xft9qHPLEqMON2DqP/eRaXfB3+CkI1yHWcG1gClYW8wSJ250Xzrku2Y8SuIt
4jplUlbMUZzqvnVsxtc2G6mPI+x6DQXEwI6WmKdpLZE9cAstlfyVMk5Nnxomum/iSVGGKElUIwdV
ZVHG0mZ8wDpIsNJYGZ1sso1xy0rZjGysRsrrhiLUmjM9oohzcIaQDuO6LP+IqyixPWMR7LvtoETm
K0sacNUnwuW6k8a3KVg/PZWt9XV3UpBriqbD3PXJLIymfWuomIaGbfL2aecMqQsEAcRcca4h56eW
SOx0fRWaAluiPdHRftTG5IqfydOZ5E3roCsPraDWxktggOUa78xyZftrP1dxuGinwNMVmKUspeoR
8riTXC3l/lWRxmJ/pIMpNRYgBIbJXoYxfyfEJ0rLOlrL2qhPd8VdpDsPwzL7yaIosHBfoU/F+H7+
1asN6Mkii8tRytU939Qv90mA0Hj+MkZQ2ObFv99BCpkgj3JlArDhQT8qPdivFITf8LLU2SHCIoH5
N5KUY/aPMuezcGYABKXdcpUTbS6lMzOJOcxfa/fzzql/yKYioqYrx7ghSPU+76KNiD1j57OpFCl1
HLLl2kbMAtPMCLvybAaGcn4O8IWK0Wm+lor10qZjzo/diQhajBB1A/XI1XuZ0tLORgejrtLZJ9aE
rRvA5+roZLA28c/Y6x0QlRxKCcLYBrKYvrCs3mhUdebhHBL7kWQ2w8TsoleY5pHewNl8DYuuEuv9
n0vjKGhYQqrbLUZ9t7ZN5moacPLMRDfZ4VrO9m+FYMfKYBCv/tr7t7E8RL9VjqH+ETfrsGvm9Mdi
tTSzog3i3uWwJGKfVpAhbL+5k3jbZc95PYWMeRx4+yZl5Xbj4Tprb30OUXzmrX+OOVOdy6hcFkGy
yGBot6cuSrBm2/jsrtOLyrO5vI+hLnfzS0s7pE88oHpNK0c0XbGxj+ot71dwPdaqBOuqBDylro3w
qNWMTyEfkKH0doEaQ/h1pFi1BOuuhqSxm253v7lbUWVtuEwhrNoo7INnPrXqTKabMLIZ+Xxym50F
d/Han0VUenmpdej7ypDx7tDjea28d4bEtcxBhY9EpePYZMixKnFeO/UWgrTtRWgHVmCXI/UgWpPX
0sGT8NlQpNtY4mPRe9+g/2LGKReegRTcdOVOCB5SFFXPHZQnLn8wWihGKk88Dwq7rXnOVg+/CIrs
1pPfaHGiBUv+K4T6sN4oFqd4OwlV4oEUAEjh0sg62Ih9aLNf5H5crxXbPWVeow+qSTc4gIDaBOCG
/oR1fhG00aD/YqxO9z2KD4AejmBZsFbf3DdpS+CQewFLEorslyjhvN///OGccS7WfLlTCPewng3W
9tzOd2NVVDM3mjco++Vgf+4WD9QDrTxZ7F7igjKCTblcFVfbJSOJHf+hQA4HKYTKFeBKQAkCNho9
K1M6bTPGXUoAvjLN7UU534vSw9KsYBWx6AutdxPVpirP8qHI5JRNTXUh7XeX/hx2iG1JpIwnFkJC
P9YqJn3i9fGbnrByY0ip/BJsSnGG6+dXzChE7+uMgPvZPQPqfA860Awyaw//00ZRkdzLP7T4u2H6
iMr9ohE569l+jIZs48+26l5ViPSHZgs/rXND5nqjAjTcgD1/0Xz4iu1W/kkQOvkINt4wvm/y+fC7
SEN2CU+ZHdF/FCNU47luvWrGBdjgheFeByE3BMxVWQfKd/1DoUhB1wtaQo22Oog13UAGYATjWBn4
Sv9rKVLlKhz3VoVPI8AG/WzdRO31ydHgtYCgCJWdEmCf5ykXbHlOSadBksIDSHCZH0eeYDZoA+MP
LcCz0OJj269eAGPZBNTZ//cnbunAHj6bElQO3tHuwZ+N9NGP8Ir3nVGAEHrCOupY1QLRbGInjjqf
SoWERR4A4XeBzrlVawPDB24TMrIZmdSP1GsnMufipcDsu8TnVInXniIMWzXcmNbNx4xf6N5l779o
zjjYqmyBF1bTRTT7akuxSwESIfbVpY8SacjhjMRwT+YaxFrEXEeTjDP9ovVJ9yYj+t4OO8hCwrBD
ZVNFPSMIKfTGU3Ar2/ezTnnfb2SNWb0Ygi7TCaY2CtbMegzGawg3xMVj6CB5/fzFzrqPBsmvdfOV
cL63qdkRCgAie/iS2/6UV16ThKRqK4iAo16fk1J6wy27441afeVr955x7lHMKIi71FOqdjHiGu6h
W3MKludRfRa9QrZhH9jxe4fWyTrCDPk3tmMQCfaWXEYoUhVO5r7jTGNhKVZofL5yYorIYkEwaQtF
o7RbCOQPxgUgLFjb3JA2Djemb1ekat+TKlizujYpf4YuiugW/djUqBUa9nJwDR6C3K1UW9f5pzg1
9Coslj1yp2XHC++raswoGMhUBaofIT8S3QnBMYRIoB4k68Xr6gbrLR/ySQEPPmUkrPL+qRGb5ijL
9h0GV41mKOO6cJErl0AmXOmnkl92L6wc72Asg/bg89bUuJmVucMNJ1sLQfJPcbnjmvNy+nWGn2Vu
6hsk9x1mYNYVBNQViu5LGPV5vYgMyp5i+r6r8nNVjHz0OIryfOOuxjpJMDEIryFmgfuu19LZdsEB
R6lGrm8a8fVzt+DhzvahesD6KMQ5BiunF8WsGxXZB1xE4cXUxJdQy4+MwVuvG80CM9HLFXZ7gBVa
MTJZoc/7GBr4xNhDI0BQPbe0ervE1KcXJYo4zfcqZMQam5uodaTDaSH9FVdflUlB/NNzpI854Jjl
C5iahWgkct6KNW/6E7yyhZc8KuEAoGJTWF9Pk1UMws4rcarECfjqeVqfxl6H0nm3HpsOqP5HrDDI
3+KfDslV52TnkE4xUpE/QecXFTb2R2vrsx+25TECb7PIXOpD6vQfab9Ak5Ccxash18MekWxd2FAu
JJDVwZrn2dg+9mPo9kRkU2jIffXJt+PjEXNmP7lZE6FjjbzF9+Sp5OO/KIk2XHZB2q2MSxAd/Sok
X+nWOP2dKFt3n71mfpylxn9deTt+vYhRUrumV3oBCM3q+h31qvyN5w60KG6iJFI5SQ+KZKERGQvj
UzQRsc35VEAoTSYuCeGqOoIy/fHFggsH+bECb3Zs7Yd/DTPxur34gCpqczturNBSg1K2U5KFRhcx
yd/v+nc9u5tjXc5ifPJG2wYMFyuB7ajVTktb8pjPedGNq4N32A5mb67HX52QaoWe8P6ZBSJL8AfZ
DJzBATaAOKP0gug7IOX5B+4U9NEnQPrg7Bzw/+vH5z0GWST+cyVTaVdU/xI36kvB49vmUkjaeuwV
rwZBs30E2+mdyBk6BIO5eCHjRt9jLcRlw3XsPSr45OcfnG0lTViGTThXEu0K4efsxeop7iawYSH5
ZWZ32AfEq/gKhuSEDSpRo90Fbnon/BgqPzeqxXi88pUnwPSRUZ/GApHuMO4OuSAZRz9LedH6r4qO
CBIFvlnzQUSmVGMFKZ/I/nYlAhWptvY7rTDik6RCELURsYepe7ky3DRILb3v2nuQX69NVWgyEhxG
zEs6PBCXwrVt4fRY4MYhqXlTOywWL8Cx9lTK52zblOPVBj0XI9+8Vo/kQ+og8oSeiqnM7omrYstz
liJSzFTxcU5DQhgdJ3hVUNA2xyTEp9JTn0EDcA9KpDoisv2HOnXyki3fqb/REkyHPjaSniH2fwlP
sYjY0XdGk4VUQg4KpgA8DdJTdyQvu1UstqGDULQhRmX+nCXN6GIy2L+gcmvE7pKLS7462ulDL8RB
iY8FNUqHYvYlFGaJlQqrCMlRSvB1/AtVesSM9w1/DBs9HUrWbHycesVt0OM/FlE5fAqbBhiCE/Yl
m2hA9ZUj3exoG05Vve7YVBbK1gXDO8W9AaP+Fvf2n9oU/CmIFxNEcttFZHu5N7abX4dyOUzb6g4t
fM+KrenrBZo17/rk5RBeVolwIpKZ8dHrGW+QoR3VSDhMgT7RdEsU5xwAwssszPYdYrwKiekwzzIi
Diu863yZMdMDsjk/jWY5hHoFBSNhmJVD8wMEgsacS6fCFpFv5mCRJpMq4Yq2FBwyIEQnyrWccOM6
OuZDfQCc++st+EnZNNXmLfQHhDCTRR3GvAcW5HWhO5F2W/kE36ZbFnfQH7NeqIkgyLPeDrIgrgA7
5C/d3L/JatHyIEp6zAUEiaaloVq+JWqNbNbgc3TqxBU6QxJOL5wwUtFNePJcQe+5H7cpHQaGzXDx
30jjUbEKn8KDAlo6SajqWdsR0T++Gzb5MJ94dIyp0jqrBIKh4naWl8QRnE/ydPEw91ai4OwkD8u2
meOpwjM4oQeSABj4ZNcvk4jyn2tTtZIf4cvgyL2icT7FyR2tkRcXIpFmTpKnDNd1F69s6NyszaIk
mLnObPZhNpX/n5MffX0Z3ouyd1PHudBPySn1wwh59RZlmuUy/pi+Iz3zRMJLo1j8bC9ZPca3oiEi
ZAgsx2oux1+jZ0HtPA+higwZuUXTKP3Dz3gei2YHfwUWX0bTIEgtV31PPRoe3OKO+qWbMmYIpFOR
G2nO3/seMTc/6T2ROJ/Q2VgcxeYHPj/lSjzr5RWRw5I4cFn+wv2NU8dSRMqumzGaYsBaT7i+5i0l
+/lyG2c9mh1Kank94OxcwdeIW/ZE+wMJTXjtBR8Mpu1wZgXmX9PtUaBVI3HA3S0I67P65M9aeCmW
V/hN+W1/4BF7T6Dl98nol5ZpgEz1sAkC/Z6xlJRRJEYcYqJrfCveqcbekxT78JZwdztccbQCG1sf
ARDTmT0IYmYSiLzTiI39KRgg53C2yF29vKVGegnH97qSLbcVeeUC2ZOKP7EUIQxxY5HmleXx1VA5
izU7oHHamAIORd+TKEtEOCw4PZ7q/hdVhiSY2aIMg0evkg23AADa5N1s/K/z2chG1uVlm6vv6SvM
89UdOqFIQ5bNG48T3wJGCl6bMi2qBtBmYZsiexPMFPkH7DtxqExLAUDY545Sto690TksJjjNzl+b
hGXbkuFAijmD+vhgs1DJhn+mBV/pOaJ75Ji53anHYSVecpYHGj91/eCXr55UioLVJ6Shad3ttKnI
cxA1wTR57fvaHEH+caATIM3v4jHBWBbwrGp0u7JkxaC6CbgjeKi8pKXU+5PbexGG0YeIvDnkYvaV
WYD9NDzBuXxKURK+M3SOva1fYRwajsJto6uX1drJTbsLHIAkcIOZlDcXgk2DDE15symPYbUPO/+V
bv8/hgvr0yGXw0sw4ADExV7AKyEpE13Lb+d69nZiOLi6et2Sk/pefconKelrUfnTNkPV/P+PEnJw
QUN6YickCDShtT17VEkSRPfnx2dQfpgXzqT7K5kx6KGEBm/NLth3jj/PiCEhvsCXcQpSRTlcpekS
6Ewa71NZoCyoGTVbPaI4ZhzArknaMMX84ggW1YqN2bJ0KDY3oRmZjboNMPcUgxbZJ4IEOKqRs1TU
caHpcg+pWMDJA181JadKstDc9ZDpFpdhgKWmjSZ4vhjpgjlyfxC7mR82OWBHcYF/0IUOz3KmOEGg
zdahEosHNoadi1lvGSJ3wRq+NI4ecdG9Mpxr4o9NnwH9HgDtXSjgqJ8hyReBgD692fXgBe+41Jad
ZsL0INajFHuWPJV5ntaG2uO5LR6x072v1LrTUHBdkRs8tLHQRzazKPcmXhrZCXOr7xi7PjFQwSGc
N3XKLqll3Zyygn3QJ6KpFNoLjq2Z7lbxCPzDMccMQgWAoIjA5JZ1BGM6fjtMf2mtyMujZltzuHkR
12X+TQpiGH7Aw5eLGr69WA0eO9+EsgXJe1WVu0U3f9sOJSVMdJa5yL6k1+JEw3AieTRtZe9vNCuF
61iVx1hOFwR5FkIFJRRwK6Ta+cLPIROEU8tGY7TVz5ElPIyW9GCmpNTNExxVwbgjSxnBavA57hHt
yzyi59wIUlZuvpa0JaAmsUs2uaJhIyb3XDun1Pay5h+e4L77BY4QQ1mqJw8meFYBcEQYVF7HRc8N
ZkLWRjt2Czz5UNsW8MjoNoFlPgZ7jRC/rJNASfmHPCPK+BEXvUKrwKMoRzsP+bYtC6mdX3gCybf9
nPkaPFvHaBim5fsCXPswgmQFLinqhuO2+jUrx9H9gXAZMQAiC0UMxy+tsZFKHEjvwyX9EQTgDy05
2AKuTjzoMZ9CpaupcLx7ipcJMvkMzi0Q1CIk10VdxKFbsmnvhS965aqIzrO4con55CA6dnQuZS1q
QIcj+yD/uprbNA7TZ1+w8B8Ii5V3i7eJ1kaQXeqrudJCOtRp6hn60PocFhk84WvdVxpdSiG1lTOV
Y0gpwKrDPeXaCanz6veARLgJXypO31Bja0Vxmn4hzSgEuuafmP49uN4Fbv3ZX4DPz/2DNfLzHiqx
H+KuJcGIE3ZD4bSkbHKwYnWRW92erjGAx1h+4Y0gFnfacAmtUE/r0QYI1KfkXMVS74xHY2l3r5hj
x25P5fayb+nVXpsvHtsSzGBP6WBKKdHtWMnL77uDdeyQ9JHXR+Am2LfqJbWZd481rrY7/cONiGGQ
4BnkmGFkMLocubImx49y1uE422wYIb14vefEntuLwWCRQJV8dTlRANa74D4MecgSz4SBN5ZoaO1X
Zh4+1ceK0advunyOjf8S8UpZnKiFrMdDMTgBqgWoWo6MwjKyw+UgqDJnIA3P95mQ3BDMxdJ/Oc63
cniWnYS1BV+u1IVir3YA1fK4cHTjicd7XFU2d+AEFjEHqSnzB499iUWTQZFxTBKa+BpOltm1ZN1j
2oWfRtHvMdVFEfp35xaXhJlOKe/ga5UYwv1TLjCmwF0/ZJyXsuRRq/lT4WYN+R89+Qt77s5kFC+X
B8J59HSxrXKu7gsMsS9oQ/wDJHu8AxfkMJRH4Ht4AOCZpBsnTnFLyHt7TFmzYRFz5MijOxWZ7PgN
4wB1Ji8xh7/GOAvng4dKm1KCH3aOP9abSzM670HBb7iIlGmSJwLqqOb6SLGT9FKN7Jj7aV6/MVVl
HonnLS6qOyNbmOFzSnZerfoxJqeF62XS/Jp3gV8gZjaZLwgEhVIAEiJKgmN3+v2GW/eb36IJsswv
4levRY4IVRQCf5qRbTQEgz7m/JLcNCRnlHuSjD3NQv734AizrmGcWNYBplkqs/4ugwzm+UGTndWi
CJowiLGfBtd99NOHo9yJmtp/uTVoQ7U67WrFWT/vM5VBQfiAe0oo2GZxG2xvIkpWLcHZqVwgUVGj
i+L4t0tDId4S9lBqCkyIrmY4wkNtQInN1T5emt6e9SQiOUzGrumJph9faHVIKqtiGB6Sx2uG2YGD
HBeCRseaowGEYmdNLagdaSamzyUPmb19WQCwcWi1TFaNIriUGp9xhcjcf1kyITfaBC/AJ0CC9QkG
5PXNm+WCdr9yTv87MHDmwpvh6W7Qpgt8kaxhqrxYEC5rRg9LRpChH0HDM76vZVhQtZm0h+jKJZNR
GjY+9UMsG70/qknm2aUGxWQumONCgc+5hF8hrXAt7UcLHXQabeilRBRuMIcCXt+yNRwlKjuWkC+U
Sc+L22QD6G2vWAp2WolrZiLNUDOakzl2oeYlWey1bi2cOxgiejK2cDH+We/mIhA/qMWEaw6GcWss
yNHMI1VokIAVpAwRQxyHQrt2amwE7a2f5va+S3xVkWSfx75AZjYbvYZk4k4PfhI7Tdx8ZomymhYz
0VcJQ/TWcbpBJtuzLg2wPOaTuK41qD9KLHOkb2Xw6LtfYzFokDAs5NVFHp2m3ksZevvHrG6hOa00
LQQTfqaffQwbaukvaQcoXFdTIQSlVJTx0Tju+bVpRnSr2ejat1DrCLc4CH4fiT4jgCNLJ5zTHEQ8
WL1g0peUQUwb/qbe0FLp7rafCz3zMa0TuE00mC2XgDufJ0c2sqC5xMPsy+4W4GEojkqHaNa57a+c
WLmZPOWQ3RAiVaPpZSfCn7cW7G1Q+sSXGE0p75My+BeVYOtTx1Jc2XwKJHPYZ3OdxRgpYfzMrUiV
XnfBrNMlLO+e054ExbXsOo32kyyckxrl8s+eV4sVdJSsh+DR1BYiJcKGvGft2BokyrktQVs1pKXM
ZnvLMgme/TDwXf6m3DVnsRHDuXt/UqEhlwdDt3V4zp5P7bqBlTE2U6OWWfyn9xzZZvzLsoZctOyu
ZCisybSRhzAoh/s7jcGvrLQU8evi/NqJlG9pX8NMSMeCzys8Mgs+S94XlvWEvtvm7TUjAoyk0c7e
bpNy50ZOsb+cqmlyDpoWe5ar2463t+fkbJejAVBElBUvcXekyyLBpPkVwjuixpDw9G6IzS7w/Jxw
6WY7Rbu3ebK56Ed0IAtTtu16I7+qkjDQXVBMJGob4SDo0Vf2NWzEI7OEL9tm48d/Fuh3XVCzWgkG
IlMbjxyXZWcvf0sBhF+1ejBfXnnzGkSptlV8oRim0jm6NE6f+8dKUMW974XVmNXAS1qSkjFcguIh
EbNvLc16KqVNJ/LfUdVZlADzjF4W2MQ1WrY0X79fZrOXd86vty2G4znu/W3WZfNlcSP9l+L4qCso
eRpfqyxXxG2APK5TgTVGc9S0FmVit3etbUPFwWFzkxG6IuRqqzQsMSNANPnwvOq0BFI+Z7Eb9fEl
bN/Kmv7cGwEiyNl5AesOaljoLnfbvnS/Clp7MjDFSUbscDcVZpt5WQioepTlbOwTXGaMUoZ/cdAN
qKF+tf74r1wNU2wsL+GwvdSjWLa2QlFo/riseGXWVcbQv7+gW6EDIsQ7CvrOuoOTAM2Fd5gWXak5
KfBCHZAhw+0PkCw+q5eBUF0fXyvitUpMOGKRlR5hRd7jD+54QeLfD23vYZyVKB5KPwV7FuR5DKpY
m0cg9ckQbQ8X/qL9CouRwu/27icAQu+ZB4Y23WHTSxuHGMZetoJUn0/l9bktrDk5FsUpvmu873mT
/f4t/rHMLpuM88EpGMX099Cz4F6Bvtiv9Qzhnba9on6FsAEL9XgpN3RlMXssJRp9M9EUxM+4ov8L
YWLOVU8KQwaiL+ZWUnePo3to4sAZkW67qKTSxjGpusJp44LRzTmzcziKl9Ulvy7W1uWHTQZRhbXT
hxYV4UfZkA5rB3EcmJDMxxsgfMXJyF/aKzgKS7XTJs/wPrT4iR8U9RwKXYJFLXN2CMwRA73ifIiL
VD5OboIvUC0bhMpkgfrullkEvssaI92VbsEjKYh5eC+ecR6gdF/YKMTMn/3i+CxsksXEGryIRybO
t9UlVEihcAo3v2faWzrqCPW3dDeAOfVnXJEEGeqvMKF7qrME+yGnowm9e+TiiaR7RL8Ci5PvmBLY
GEDI6rRe701oA4/9WnSf5kaxANesnDIfGw86yWJdNA4G2GIK9FVEGYnPqCnhMLYNTYtYWid5fyoW
XsZkvTHUCczeQ24vKRfyIkOWWBXu4+/R9bj7ZEwsf2AKJqOiMEwmG7awhnrdGtbTeGVwf0DzR5qM
YnW31VC+1Rl/o0RSSrsDmJ3EzucUVcTvTUoYDtZQcBVZ8z8ezyNA1R6HlwAmProQqYoo82OIdqRm
8TjP/7CJOJMIi/1PIGXHM/SwNGeAyIPlL/CIVRwN6zAbYv6ak4cyCmTys6zYDWOtRRHuq5OWV5nI
4cFmnsofww5HRBqddmo6qYPrSmqRmQukB8vGwp/g5ECMpH7P9qzkv0kEOhebd2ifNGdYnJw2N5Uq
GHsEbGWOoAEn0S365E1Jd6xim8qDJ2ozNvhbtStJvP0OspNLgi0fVi/ebg+zkOXDnHmvLc+4Tp/D
8ihn1xwSjl5YPF61TBnizI/vio00VfEox1yWhC+ySJz0E34xnX0tHYPGOvjLdvm14qH7b1cj++yk
GcjS1HP1PTgEcbTi/4auIiF7f2lZHseHVrRztiU8T9f0N2qFMoopx6VTOMjwwDHxEpkdiTEsp4HX
2ZS/1zVwwxBXkYSpJLSd/gT0B2XWFFb2f2BZQVwD1d29CgkwVOzuCArvubB+qivuMQDcLapkJQxT
e7BD3Zmif9yesK2cZAWJ7eGgv64gWYKiD+jD93jg6Ila0nssole4yo+bUkgLMzWyK/1LSVHkQl2g
ynq9OIUYfVNjTHanP/PD6AHvBwFnTBXO7qXjZEM0VTRi0Jw3vbdr/umY8xMuuWPQVFNuERgQt5Hd
twxwtIdQAU/OoL0J8+Zfotks2vEVdGYMYt3fhDvF88TkzFTy2g99CD9RCw+F+Z+ULYh6f/HKk16i
7WwCRR854ph0yC82lkN+boR+ek5xhWwd2iDTHlhAv8qj+ey9nJhq+/NJQiUvBGfLDpCcb7G5mImE
01tEFo6AFhDgOTD0MLRBRkRy1Grtr5cHFJC50GU1G5dfAFCbBKywpkDXqhlSbWnnDatjGPB66h4W
OQY1Mam21HrvwdYWisBD7J4QpdkyZ4M10YPzWorkk1mORwz3Z1IxaWehcUfzcWS0ERPa+EsoFi8M
stZ9EW6KsVtX5iwz4X6euBLbDZ5hcoGo2DycIrdyYYfSvN7qbzukts+YzlfnxtCyD/hjQ3ljTiXL
FHXNrOSZr6IHPjYOwj1OolK/cprt4W7lh0s1GAmqJl2qnPSk7qL+YaMce8sHJOjfy/hFZCohNN4p
E0CDHSEktAL1+aN2MymF2DaSKz2u4ledHkJGKohs9a/V6ZKy0wVf6OMLC8QVmephh8TprdzU8FIJ
f7XWJ1YF15Q0u0GdS4Awn6FhSpAeglPa2HaNVFHAyo13l04WcFkWEjUbYb7DrMMORFO0SMjfkLuq
LgzxsmLaAJKBjdCJutfbMuRDw90uYYnOAHTDLuzW/nUJRpgNOnBaZBIThbgvVt0Hfdzp+nVZkgQM
IlO0xG5AxhGBNCh1ENI78yFDM1ALbc8TgPeDm4eXkH75fsxL4f9LtNdaNrsQo1fkyvTZ+RSOWeex
hE+ChA04yDSSnkWhtWaS3zFGtLy05rlR5A5LPZkvo/tL7hy3CWhlanRf/meZ+D8LOzwTbDTEMwIv
z8dnisP+G7CrfbH+4wBKfpuAXZnwVA8hwkk0wm9E7L95HvQy54zbE0goW1JwdB8z5vez11EaqhRL
UsC6P5WOi6ScEZ4lYEMoAlEEELIKG97ckpWIcWCp21bau4hvWl6UeWuErliz5Uzq3zd7064l7esS
gyRzm9vyBRm0c4MFfGomNKBIWR0Z443d3b62UryuTOKvv2/gjGlliHXB5NRnxxkAywzY3H5katz1
S2TSh4FDk+2jQqgdtfqWIjkttkkTHKKT1jOvdfcq+pwDLtmzu+5Z00kFrwvbwfoJEh/2zBb9v7K9
JfM/5XCgLE6o9AZDcW2Io4EGvNGhlixQUinDYye4QKc54XYhPJbM18IiNDwQgYs/mIhwi686lpuX
zbxgHRtpJM5Aq76g8o9AT0yCLPYNH+8YVLFh0RwSTPpQfJWVeNf+67mGtIkXaQarJOjehxneo6G7
vYDlodwRP7Q/fPwZvtjXv5/OC4UMnFkxPDbzaU1ztqTMV8oz8w/2odtwPQlqj10+JoXroGxXz7tL
/Oqos7aByok3YGInqukmBU3YnHgqkOUjGWC4OCzbY7oCUmQpfKKPLrkK5T8XEBcuqJXzAQSHG9AC
lKKS0I5tLvZ2SKoeHko9Oxv7F4hwtj0iMJJlt2hZkDoKSUCW/87NCy2GR5yc15ymbLgaZjTe2rKK
YeKWlONnF7ftGpdCSH4dCClZyotZHf4gHBMZPWxUq6xd0Qu0HCpGLr1YaDInRffAPQtLS3RQG8m2
vwpYAEvDUCvCAqxal+cOcGNe92qrnylcgAqrceGQBEVlrr/9KCQpOdTmGu2jCEBLiYvk6/tdMuw6
9BcsAspweMdhyLp4jZCIm59haG0c9ZP/snaVXkl/4UsT/vnuRBPHYb63aa7iqTHrJ8dsczDBqrYc
DzJDMMKDHrJEhKMi4u8oUP/6e17MhtTcMQmVYgWAYs4dOI9OqcT73m4Dmj+nDBP4n0mMEJqheyJC
dZjec/82Q3b9R2vAzwMQIGa0s98CF78kDbldUeal5pWO2lbIHX9uTxHQGt2MKDCHLB7hXee5hWCZ
yLTOIEHSvMLLMFjISHHgUK2Vb5QyPXZ2YbMY79KgYo7MNX/Yf032yNNUAwxJfg3jt1hr8EBDPogv
AMjuwCwpoL8rBFxZzsAdD3zqY4MgdlMGhaPhvOEGkZv3LXhiWo9BZ0YFUfQMUdwnWXSGDZ1nL/W7
nZXkKMGmmUGgANYt507WszS15YLYyKYegpH33EvGBocQgptQ91ZHlIdqOVnbwB7gNlSrCzoZMtKV
wEmh2CZRSGdNpGe/oWCe2jak2cYXyxCkKVDgm2YUpyxG/imSb6bzEre9PKx2WDhMpwLh+i0VdLvM
Hq7pdsJGBWy6s34VvNJLoY39flMYaSDuzsswBEYTE9RsWCwqvKgh71iYjsV/wtUpBP1NvOR30i9/
z4+6j8ePq2QCMQFTz81qX9WmFelHbnpB/aV/eNFvwDwbUT2z/KjZ5livbLk05DhshUymFZp1m5L6
xZy5IXtSJS3eO/yWkeoZADWACpiOCddukek9F++xzGnWleubjBnxx/wkZ+2sp/E9wnuIF+lOg5Y0
fheYTecqhIoHEp1v/5Cfyhx9zEhN4Pm/0DUY/hhm+nzFmkeUsF8GaWfRYgPxTd5le+WArNMz7s4a
kOAAvcuxIw0t6orKp5bUfFcPszmUBZGvVwsXlhronBK8ACp133SVlPA8mvuxqCxiCI+vNG9q3lwQ
YEv2+amO6fu5jSIbjJ2nCSXflGjgHUR1dM2Djl538x2jRHV8PY4Hh/L9C21K2omNDt5AfNTdwwsf
hF+SNGVPhFSWHic/Z7y+dkMQGKru5TbI+lqrer6u7erZ1MJsqMh112adrM/pTTnZLFq7I6kAxqqv
G4Ge2QKzqri53jqa8cf5I0+qXoutbElQCWwCAa0ejXFvwi4XnIL/oQI9/KXUlI9GOob0744f77Bn
kLIOh2VN4EByb0c4r2SPyRK5KXMCI48yQsmf3n5Ewwkg9oSxpMlRru8B0Etsprc9obWU0MiM6ay5
FKYzt2HqjC+a3+7CXlWxi0J1gF3mux5p614NDKRohxL1xKPpgzWmUodUUNN0kyDIbt+1sv3zyL+B
xIDvJTXEWrosc2yc5tl35qhe9kixSX5nKQT31hFUTEdeFXSLA6bcwLIg96Ec4gVPXN0YJVAO1Y5C
RPuDPDYEq3eOfsowHCo9uOzUQuQUB3PVvENjgMfxHi5qbEJwuw1P47fgBPML3DJdEhpLJCDaSL/3
jSwWtw48iO9qc/LsswBy/gU5dqxnFiNBjoG3AjhQhpFB+OKkmFvybiHxhbDWK8yxZFLpv1r6SJ6n
iDVfcVAw6rTWHEEdkZU8s867AZ+ElxV6KN7L+0VroY8y3R6Tn7QEhXLlZrnnUB42oKi5WnDaF6ni
3Ip+BwvkLmov3w/4G5mc7GOguiy1rhUOtLNC4OQALUPlBl0x4vqUE2mENznxfQAsoqRTJ9TXzm5t
UnTMFR89BYH/M//4D9PplfHNVcPls/rc6vuoGqcwAg79uVDBLzJr9TrQ3JR0qI/IZpbfoiGc7L2L
5YiHsa3oJE5tuMFvADyY2kqiGo4LykPgAPL1mwt3wNY3/eTr/zkaDLWg6D/rpL/Dvx+EIjBFzmkK
dwSWd4C8rDfrLiyxXGRVkYI8xO4syiw6c0lGTLqtXzDWZJltX8cHVOeqZ5XbBLm4dmRJtMHHFo8O
zlned5ehAO1KHDtZUVg6nUEti4kmxvUSjXB6/GFTlQFe+ar6TIQh5oDCaTPebPigExKZYV/u5SVY
dg+/JhSYHTy0sbqSaYcLTVXZDrmz49DMs58ziS+jX89uU6qlMFUJVVrThiYsSU4HDG28k7thakjL
Mcc9nPNbalnPU7JEB1QlHlHeSl/n2a/WJ7QK+x1Cv2Rmvr+ZiUj9m6NaA3Iewi4zIrJEvjy17lji
0n5bW3hvt+E9krp0fRBpGBNswuQt9nIXLv96khhd18bfNhiqHhv3A+ltBFY1R/ULMHoK1qw48QE3
LOxkaIVza2sTK9KC0AdKkIglPFuqNl6JawEFmVPZjRzsyoCuys+uGacJL5Xcmu8C9hFTSgFOg/TC
E1wkHXHXTSRPcagnC7T8OIZc6f6OAeHbN8VkeNpnpAW5PE83tWa26m3rRGfByKFUu3kHEvraiasX
7ZrayyeCiIEAaG5Yng+JlXlR0gk4hrO1TF1mQ0dehWcrtOiuxObfl8Itn4lI8of1dEjrKJcpGEYh
4GxxU8D7Ciwe5gCOHaA1SbxIGVtjLCIQUWVIXimhqZ4YAzTLI+c80Ixj2gqo9ytAXxXco46scuvY
T/RAzPzp5wzlSTimFesAb8K2OvYrsSnbo7Hs9a8cNRlsDynUm6SQRv1xJxzKxXOlt04+uZ4j0kYW
BOFEz4J1CUnfcNzPJFDwghUa8YpNY9dGf4dx3DMElOq4JXIoAvw3hNXFAbCIteoYkg50dVQsEki/
H9OGnJzov7yV3VSQmjfjcMTFCtEDePmWBkIqu6SFcuWJvWy2nTTBuT74kb5tsMPJi4rbwi23yPQ9
g24Pux+BGHyZf/zYxUID9NQ6085dgfNu7TI3hMucHX2ssmJtTvi3PXtksbML/PzrS7sJP8Y6LPO4
8eXz4ucNxLb1gbQz15nTNetahRmS5a4odo+ZdcIROPMVYxKFhH6+x5BiYTxHkqLW4QYJki9o3o/A
B9Wmec4dYAg5QisDCnnhJCWZ0U6NjSDtlnHguBxWM/trr9PP0IEiswbj8aO2JXT+hFEb6pprSemC
3UzKqV4L/xfi6OD306PGUiCmzvfzyZ4zfAevdfmxQxJs1KMQ2sdWgMJ0AoN1ln6ltrkWcxD8lmyo
6giq40lZ63zxmskZ3ZoicpOjeyn1scXYS+cv5rIm4yRGnxiFWeVHNHw/fpzmaY2Vx8sVd1pyaIsi
3ZFf6jTb4EHs7HN7YKBQHQiba3BFoLKpRTU4/GnqaXOuM5Lw+q28rfFG+NTKsm31DixfTgIc7rrS
sJCJUM8+lozLjHpN2hEcCvpRuUGRCbL9shjZiZx2U2yjSTM/OLqxO/0jpvPkpwJk1uHIzyDPcjPi
79VNw+JDhOSkPAjcu0ZXb2lLzTI3uRvw7rZMHKuJIQMzwiGQyuBCT3zce5NV4HWifxDc7VXfoeN4
+zo7HkL6znvjl/2UO+lcdGgU9iDObnvoYaFB1IOs5w9QeHjV4oEAmZFXDkUvh66XTjBDBufPqW6m
jFJL0kpylowcQgNZiqtd2pwwNqpVO8bjwQElMYmv8VaoWeZhKnbvi+dc8ONgQKUMdKmcunadrQdV
2tRgLCyI+h7mW9Xoe4UQfoSeh3e7MM1+tEj8Bfd5q5mV6KSFuCC73Bt104xabNUOnkbuw0VKF6tq
33qyPEZwFAMwqqhI+8Lux+Bb6nesC9q/7VII/xmzPz4984KfomRgECgRywwPqhWBokPi7OQMp8ZO
bBT1ZagKcXNg0IbWwEML6hJGb94tlSrzpXin2HTzcQpjnwZoFoiKz1zYZqtk9hUT78zaRDnFhvUK
h9BQ+Ufheoqu25Te864aS61uBFAdrPI60Od9MGaWqjYEhTZHx6n1Cv2c3g4OHIHVQinmEaUGKn55
q6xYVpOyfN9PB1FEKT+mKmXctjLRhnUIIzio00NtPg81GAz2zxP5degiyHMFXYYlb086bptzn71S
iJKHNfmnm7vxXrJjbhyvg3AfBh6ogg6e58C32T6kzSXlT1Yhp2GMegpFA5LLMsQ0PzAWbxtj5ce/
tsPTu8j820FyVAXUQNp0YLW4y3n2yH4OKwgnlAsv+z8VlUnDYatcyR7H1IIPsUmknxQPrqlEb82v
OCKvsioW7Wz8Fg553AIiDDJG81U1P3f4+bqma/kDcVU5XHRyPJjS+o2LGW8JRh6cuBQJDkEz4URu
pw2PARJ/CkyorJ4TXBYCreOGfDtof5QrXN9zRSHm9uV6ush2/Eo5r4PCtAecTnUZeOg31hb57k+x
6Oe4izLNL8GqaoBr67Ml5Xp+rKoDKqd7hNWuFbZXna7GY+hLm4O3eZFeHeXxTNfvPLwS9ZBu6mas
vbawwSQhW0ZRFmh42eww5Xdh58mO+9a9sXUTGNwe3auZsn8Ep26mhlik7YKiElVzAa13pNr+6fya
wHoD5+6RfuLCu6cpTg6OA8u6VeivsUu8CWjUWJylZeLaSHqE3KTlC4Ubx6wgHaDeHn6t0G74akSB
4z7PaACKcHS2HFjMHKRyzfubNdxYwckw5W3uTUh1N1Er3IWFy2ohMh4CgmZ65fNByV436X8eaQDJ
kJQZyLgGWtfbyvgIpV9l27nNaGNsXNz12pz1r4yv0pUw35gZcFRN7O8JgPZ1A/skapBVOgtkVJ9Y
dIy+Vo+Fts7Ts4d0XYtrz7ziyuHRU75b/QTyW82s1F3gz2dWNzTEnGPd+0JNpkyHTfeNvk4674M7
d3rQYtLG0msmDgneRK+jw/n4vI9zrSQQ+JQJuu2ReOehrbSmNEUpj7fLAyp19+0gLYt1zvhd5Fjm
/cu0NsygmGlp0j2INO/Unqrtc3zjaIo2vl5ipRLS3bV8u6uMYksfwAYZ8O5mE46bKXYtaKAV6Xfy
9/fFfi3v48YycS/Io6VqR0E5+tLK6FYgXdqbNrbQhkLnVBDmq4ggDsnKoZ59MGOG5SQ1MOYkmF6s
xkPUUjI4Ilr7g3EuPDteh4ukj/hWkOpy1YECooqjSffFY6JbC3Z2jw61z9wzgE6wYkqBOTgNXIkP
CxrplMNvGjJBse0VXNhKB+hIMUbp5f6n6ruWTAKM6tMM3bGolsG7ZoBHNXpzD0lIYARkoCzGl+yY
ZquTP1Pc40q3A6Xkc2uB/o8vd9Ha9Y8EJmMZOqy2TJ2APzqnjv4JWko83BjfqyjDHFZk71og96mG
GocYgkYo40yh16wRT3enTSkUCw5aC6VA8EXKSIGxgyHusKwuhyP6wgWy61MO3Geh1BM55HtH17YE
MRD/AIWYsU6V0zAH72FM5M2KbBr3780pQd9fD4goso7jG9OlrUkOnsd7Z+utU3savKcrobshWKdI
8ZiyoudXuXYEFHZCJikiCMxAOYdwWXsw0stx/fi7TZTXWv1+TKe0yCrDQGI1eBC/dgCLoJNlrcis
kEkbZTD6bVJuqDHrRjxBsCzFfytgF8ixHBfvCo5YmzNfnZdoujaKiUiaW8gBfTIqxe47yT6H7Mtc
mvl/fm564S51uTDPNJvDLPRTYotV/YuCCLNARp8b368YVINhf1zrZMo3aLamSXHj7unsw0DupBuL
vCyjj60cWRIfhfbVODHSHXF21dGnGgZjTfs6crfYlCPf+VHE/ZS5LO5FSFzeGU+bOzHXWKuhXQoa
XSYWpLodkwCtp0aK31mcHsdyeDbZK1LIpyI7+d654MBMorRxUFG2jnJU/aSDmMYJYQbjKUenOJPl
NwjtkRshIEJzhgcDZv31/fRJMoejE5G9cnMLpsPxXq0aVaOxFOXwbaUHtvSRaqTNTm3mTa/txVPe
rtIWTrZey3u+mZisvpsfFXxEu1eowjzsmq7bfIYKTXunFNhCEtL4TtIAGWDuVnz3v+QJJBoA9tbD
6fLhppjZbdnaTx9RjMniUcpDcXf00zrHk+/11s94t5Ky86zUnOG06wx/rzWi9Kx5J88Rnb5mnk9w
uKHHvd9XsAFSB/LNYXZS08u2B2wDzf0hTsAvbfZmYG9MMbtaz7hkr27MCKS5dQQ/chSWZk9Zu4Ie
9oTmaVyq5Lky0LHr2agZB/59ORKk1HJuC+KJT6DtD5bH+C1jSr2h9ahYZUF5tyeti4HA/1h7sF39
D29rTqB6zi50f3bx/1qEjgqGe9VHAufQJEBiB0iuRcJgjWNCXlEh3ybH//23SHYcDM924bv3AjCG
MJfcUWC30/ygs6NSfxtacXxxITrAFtQkRaF/twJHxpIt6VnkPIGh3kC2ZpW3d7ls+0Fvo/v38tgA
JaJK861MnMuazFKOfOFVgIDAIl6EeDGkpGWV/DvSy2i2cLRsBmjRxG0i+l9zmxFLt1EWWScH3AF1
5NZUfRuOM1fFC5I2ZXeFH2+0+90ogCFHj3KiqPUdExUC0U+MEl4uL+/UJg+agnwDPE7E03gqZ3Ft
0W26MLlHg8StbRvSxUeNihSDPbgYZqPLhQNboVexDA+QuE2EURnlqdlQYUSM6tpezbVxdjpL+kLn
74VGT/Ox9WMOM0Xwu2j0K41Xbm8Fl6uTTG1nImhS/vA+CYdXrEXyN5Ymz/qVZfZ8eP+fH8JCKxCl
e+Seyr2DbB3v99y99J4y6cKr6BuZdCdesaMV6wf7h9gSPT9g3gLZUxtWiIvf/IEy/7C212bbl+xW
68iIALK5Nc+bagEcciMETZUPn/rNShpZY+qDCgjnQ9muqW6hUCdfCqSGPmSH7l9t38ybPBIW6U+F
vgfJ1Os8F412WbntrSDMBVHu/zAjuNnG+o2pXxfkjD/BRnxZjd6aeuy09ntYuNn6ovudw3rWM+mv
fvflLyGlpYt1T8Yykfd5IKkRvaxXgyBk6eCx2sIPg1hxN3Hti1GN5+2sbSKES4UQeV4hSJKOSBST
JMr7/B4dj/e93TcIuxzCwKnFSYXbfrMn/fZh0S3lVIbBpPZgwojfKfwkUE+powIgoE4jUvoDX19n
jNWIOXgJ5SBr1zDxXVHFXIAMpAGuBBziJMND4ffnImpGNATs7ZxLhKSB9wAnmzNbdjGxrocKNOFL
9KZy8vdPMMr1u0K/2PLnhZAOf4jDAc8+l77NhGNILqWhr8EkgmR0/YQvNriDlwTGAo4TFvsReSIR
lcM/xg6bJDTX9pBzu2Skc3LzmBm84+agKr142nzmDfFInAvbJd6Dz/SMgsGEhAKxdqbnl/h0r7eM
R7I9BQBuRF8ubnBYxV7KxmsKlpfUUm8IO9k2PzmlD6/mg2MnnzreZgV293yl3rqyp6RNI+rqXe0V
oNsMa1hPmWRxou0dTHhrZM1TPBUaZ7VBYqAjnDmv3+RxDe7wNPRx6TowaqsyQPFYpZBj6z2HRdiD
vSe4gaFgk8EAAWtML1LOJ90YPif2lz1AMWq4M2LYI8fNUL95awq7csX6iMs43TRZbacReYlB1ghq
snz6VVYE0339jSvA1Ezg4dNfVYO8CSQsjQYtVRpPzCoCCxmYZdgSH9N8z2bvUBbTxEBjr6P+RCmf
CD7l7DfD787QdnyiBqKcm+cayhFQnga4GfjOXacEm4itRpo5nScPSoInf+2Nh5eeLpY9nK84Xvz0
C1DOhiETV9XNJWCh3LVbZnUbY+6gKU1PPT7E+SuMW3Kq1vWSFqNUUxdzDOtMFE1HQfpzjWeZZrOj
g+KRmBcGgi4whTW73oKO71u4Jf5pKiQcmY7sTgU0XXhS2Zm07AWrb5Jce6azYDgwtdfjiD6vkhwc
O5G7oo7xTBu1t9GTvUVKJk7kGSjnI4ft78ypXeImcEg+I3HwKqjkY+KPuceOrTq7OqXsz7vMSWa1
k5tOW2/9f69WQM+ztj6bALjAsuiR5nyrE/RhllxWxfBh5qjYnGFtVJSz+HrrYXLMINAwMTnUFyIc
2Va+juOjwWadeX77jlnujMZJwKv9Pc+nJGcKsoyElkMv1l6SUGs21uAPMzmKwsJwcllV0szKozLr
pD8/JFoZ+qmVFYYmYOX6q3aMFeto9jXjjfQgr7N8LCnLT2Q7LYaawJb9pe0z65GAqQxiR4hOg2wa
nk1ThjJQtuXrIX07k3MhdEddfIGm357zxqTsyZQ8uc83+fnLOzMbQNKNGMfwN81G9gJ4tzp7OoXv
3CJ3UiuudI3DEpL87i03GaaYUFYhN+E/Ldy3xbvtNawosJrXUvz7XnQ12ZRqxtmsqT5trDatfSL3
jjvL8HhIt8Nx2BEiC39OT/+XMsIY2mS9lgWXkzI+ja3q98EmxHUgJbRPxKf6KXxzsNtUYBTM2FQG
wG3zBIopHTZ5W13DL9I0u1ra4s3tE/RdAfZ8PLf9XNXmgIv4BIOOHr0TQ7Wh6ajnduKA2E0GCGB1
C0lfUeYfjRPsaOImHripXSAJ3LjkRXVgx4fGnNqROK8aHtxQnPZO4x8EI9gY9AzeeEHSC5TJDsER
anLZApcH1p2HlPaGGYvKlBDARxWmxkkBSNdj0UdH/qknyrnZFXEmW/hBoSpgqGc8SzDK5f3n3Edo
UL8KuCb5agIMQHiyp9qm/DVqOCnpdcl/EWnDhfM4AP6O+spepU9Ood4CYpEys+LlkudGxffkDtQB
9n32Fl5Ug15Oi4VvLsbXYX/5YxB7PcYt1DWxH9DXZducdAxZ/xRMLYLGmyOnWHCX9bBsduMLJqxX
JZbYdhjOdNuahgzfxEH5vk+Zo2H2WYDo2Kk5lglL8k4/miIFf7mZe7epcsUzzDFBUlygqku42p6T
GyGTKEE1G07J5FOy0IEMwETwJUkGNEsWv2d5iKcyAQK2wPrYzYA+00q2zoFsW+SBNxCeV5d6cR59
B9A6rAOyyh+EonZYxxcbgLS4e4ld21TkxEkyp4SLeZ9Jzu4PhbEzETwnUGQfz7qhnBtatF17XKET
zoIRNj1OCOYVfm1z+rMFbnbeEc5mdCW1pn0sEkxYjpfJCXCUq1KI0VXJchKq+0axwcUIwCbC1XaX
Cf5WZyReB1VtxOr3AD3hiCu19RaBCCy2OAdXwqCEhL4dQB99jOGM6J5Co5D8zs8qWRonnGr6nM0e
3jIfh0Jkvt/pvNp5yUcORJRzSHQ7s5fIgrxxAplCPvtvd8VP/e+BjqARrz+VetCt6R0l+I/jf4dy
uOS1Twi75IwdxnhwCAkkfz9nGOW9t+GJFSfAm6I0tAvR4faHX6lJbZK1O1Rbi2Uf+/c8Gz/Mz+Ob
lQ446bLfiLek9KCMAaqf6IjFZx9PFDva5MkepNz8Z4PbCZkvxbH8yYjMEJK9rRHIzDApmNo3qixD
m3Y/2c90zeLO8Zi5sGZwDPKJDwXm38vdKettNgoeS18w/v53vCvWs86dsCPIr7GX4+ZrojF5SYgI
2q26xjI6LVAjA+M0Fhd0G8PXlghJ/7vfGPwQndBPuq4Lw2eegJFEpGnu45JZ2qvvUp9gEkhXDBI/
Gv6gcUVf5JSpsyxtRSOsKM/0q///SM1AsDgoowgzqlhXZ1OGqGyjVXHQUJU0KLG04Ls7Osn1FA9L
3K20++Sj3gy51IK1EddPyr6E2FGK0mgrWNB9vEtYSw4WAUhsM+Zc26po06aL+wTUNSrYpiMsD3F/
iF25cbht6VPDncdyzf1+AzXx4FclI2+ejf4US1sjXY4NMAknJVavyA8EGptlv20cDA3Rzb1sHETk
rx9jNdVQmytlYogUWj4QGaGWWD3KJEL4C2ny0GYcC7hWbl7LYTm1Y+M7L43/NEQn3hDGgbQ7md1+
/yTKLQH3yIaso09OoqBreRM4eTXW+/pFH9s9n+cThdjU7I492PsIAr49ZEWp/2LUnvwpyLl6yOZx
OdE5KHYFPRkbSxslIQLwycKa4V+DGQGtDhlG/E1IzqWieV3NiPqaM80Q4Xs2mhM13ZFdXrJytKMA
HMLM+GxReH5YwcKF0YQIkrQNOgzrQc/NbpBy99FErH8SPLxGPaABbP9ACwTrVF4g3S+mvOO5oHMv
QUfrO/8gboJlBMrMLZXAst2GsngzlOI351VtouNT6GZbxM15S5epQ2AwEmhoSpcm+otjtJv9aDzK
obBqLuEhRlo5EoOll2OrGiRD6+LZfrwWJKRyyYqGY6FQT7wlDKtqOREdIW1iExnvrECTQOoGG1qe
3lwGFfaZOYX/PRKVmqsKGY3b1fbLi8L4Q68v8qvO2Yy1QbrOTPP8yuBN2TuCGr38kwaS3v70707K
CHYr/930HLzBnwqMVktG3n5PiG3xX5DZj9Ri6kFFIgwDz5tlAgNJlj4kGfeTp3UbnkP3+Xy0Kc/a
vSkoWekRWnC5xUpSX/Ue5FZGHc+qKvGOgzFu07IM6DnnCeHYaFa/O0/2NcqxhudPoy79F5RoLgbH
D704nNuyurp1807zq8y2WnP/Ip+ypuQGDXnZ5bw28FbGuiTyx4Rl0uyONh3Z/z4a+hrwpwt8NqMi
WBYqvSB0VT0bFx9GKFBF6pren5BSDOrDsmLnn9WpZdkweoE+1Y+qzxFHi/ucdfFTGUD9E0XZE6fw
GZe3WukRAl6JbFhzwA2bRkja9L2sqG9v1BRBECIfTBfaPuyq5I4oFsDqqK2H2v7dejlH4VrUDu8Z
MC6kmskVDwpNEoH1rN3Lc4vsXAhNwnCVxaCUzZiashp77c6AMcofkJtqAlKUMJO6O9Dyam/BBthk
TWcJyr2jTWjn4zhpawFLrKrpFW3g8hMPWR8+OaMwF0DKwToMCT7kM1m2nia+GxYVMIC7QPWPC/MO
1yaoYR7xbidPEzdufubnTW7w3SIuH9ctkm5rXcondEi8x5qihgRdg4UBJWMz/AkLtOEjsg6nYixL
IuoxElIXyB+y1iRwVDOJwfTrBa/b2CGoc+p8lzXUPSukcl3RyxOjRbYtZa17jnH4ggQHhZm73Hg3
AFaHQSQoJAHVCnkPbi6WSqN5pJrdXd87+AVKZOgO/tENlm/Zl4LX7dxcXuc81kQwtvg6oO9ajE0m
DuQTF2YW4yUC3CA9kyFp/tcs0L1Y1bL0EY55GyR6BY3sj1NGEmHwTUVsGQt8+T58jJwh0K+xIJ1u
lEKnRR6pyBjsvbGV+vPIe4eEk+eTjiYcijaVehgOtXV3rmPeR/N5VPDFHHesKbxsw5MJm6ZPmhmC
7KHzbmZcqPW70KkEBL693Xype8KduKFC92OtfC8UPs6pqGhmSBQiOTzX42j0eTwnGCSZSYfWggvn
wNECH3ziexec6JC7+Kob4U74oUwIBkunCiwk/r3c0xjsvS3QEJdzIlH7MBUSjKsnm3ibm3RybbKI
HKdnznrkB45pByxGQcONhQyepNyQwn9gk+Sd1b9l9GmwZpae24PSA+v/2Qsh9FYPiRCv2ULWOCNN
c55Dyuv39JLdcDEC7rHA3rZ775AKCQZBrwiMuq+QURF/AirdMBh8uxtQ2WhHzji7g9tlF/ZBCTVR
TXi+DJO4v2wI5ABIDUBfx4b8GLreDPTymLbLTxuytr2P+MwlJmL8ZainmejkMULt1253+Q+06O43
1+J56EUITym9V49ziIgJmXCbNozqWOR9g3yuvhJ4Yh0T+NkzFXA391zHV7cBQm2bdzjoqA/VQo9m
rZWuUdmsJie4yVe31o3kxB/vc59i9dsL5tXShGlTO+JI9WLwOTvMbHyY6RFpPn7Ojwq3joLmaR0l
72jyIflDB8oA+MpjmmNPHRTsOaah0PdUqrwri03MVOcPHJhT5dUDvZQa21H4NJlnfekilIEjDQT8
3ZXI5AaX6JlD8ca/f2BgKOe8Uoi0cAjYlV2NgLeYfLC9Pd3dmVuCXNvkF1++YP4sejAVU3wP4LYd
XLWNvAeB0fhxlFYbNjj27DBPbTyYNeY2WoFfTceeO4Ckv0CrDgvDnJt5AiUpQaO2w11YOVxAA8Ei
r0iSYSjJyLXwjWcC3bySWA2aurpNQBs4sPZ3+45W31zBbQM/y4arWFKxr6vA20mz1W7Zl5TQOSew
f0MnrN5dOjJmcS50oa8xrMZLgWw4wXI9xZ9SohVStetWw2ITS1IPZSPRm4xYpn0YjUyAlF0twGqg
VawK3qyHdNXgqWPLGA5lf6fXRgde1yTbDrX5Q1xa88u8PlxDtDfT+wDD8RCam8oSdGCt7ihAy9WH
gCYCTpQVr7TVPpbmYlysZBBk5YaltZijVeZRTl9lw3olduG8yoHNz8ZzyOe57XxLDf4D2telqTFh
b4Rym/Vx9WHW/YknQdymwH5E0YamSGwJ9h+EVO1WIaLQRHlvUYIzzHiUQ/YBgISh+ccU1ff4DyDZ
mc5xUWpW+jGsiHuaKXsOc61+7v9aK4QUx+HZGHP7EEadF84MIv71SowqY+Xp18iPuZvSXKGpGC5w
bq+qWAJCrttaaKJhrTL8o8lexmQpMuuxQOjozD19gmWlZGsmoRmLUaDeMU7vmJoR3AuMPZz+mKu+
EzCvVmgwBE2zDvI2eCUOWqaDYCkX6knty2ylMm2RsTnVB0ct0dbzLHUo6H0v8nlw57s6qOPghfUU
G6AOl87J1CDe7hLraRM0Kc/H/DpR//YiRTu0HVjx3VD1z0YjDO4SghDZUP+D2o9Iw8r+WUBa6qFC
6M+K6WTzHnFcEL+TS09+bhUX4kgzJDyhaFDLrNsxqKnG7Qm0aKI0FAxc0TJ6Bgth0XnWwmEv53le
apPa8HuXnA2ki8k+6o2hB3CEuAPjD2PLyc12h/gLsgX1w2LSz8ZZmfwTZ5SwzOIzYbhE7/2ZBIET
pBgMBkHregzWgR7+zvLyvfEwQLz0yehuPI+4ICCBEnzvczeJwdWiCVlzCA0JdC8s5MtWrwecYIC6
zahFf7Zvdn/u2G10PWYgEIk9HdpnvlYbqvAV2fZ6mN1rDxsS0NAoApSVXjh31HgFOc4RBm73d2G+
/UdChVZs/wtkjLTYv992y3PdXxk4ZowkK24AdY83TN0eIMzRwFa27j1sslfrEcxMIyEsLyoJmSyx
BXJaYN6glGO1dsZY7zrrzXOF9mFTNzTkmYvj1Z1AifJ9Txq6K60WbYam8UkT+84ZCrMsI7RrfOtG
AakwtZ+Onq/f8SdEMrYoOfIw97mdoVGIcy5k1A3Dxn9Sp+S1JK433XEViNWfbpZXBO7QJxTvelk2
SKFSQ9InadHVmqjcWI90NVwXoCMANk8wKLlNPPdxlr2EcuVP+RxZD1JPO1ynGmsBnRPxyrpJK4wn
SFp6ruxGuC7FUGw++KQbR8zNM38Ed99ypzGv3HzZtH5l1Co/DHbN89AWc/3QCnODb/HJe2dE6NwH
HLs/zoupxpY+LRKtPAv9wrHiwi06crpkEXrBFqJuIU8vEsSX6wXAKF6hZ2N4OZndZc/YRW3Dh1P0
79kr15u8rDwtx1hYhaHKopeYa7jb1fNy5gSLOKClNHBeZtFqxETrQIx+/j90cmhCyqaUNNEaeIo5
574QWHgN4wR9nZFXilTVIxg8zqPZJzlucqfydxGC5Q7gvoiPEKvHEAB6BNo3/LDpPprr4nA7H8O1
c4Jguxa4OJVjH9evaHnkv/J3h7f1aOwJgWqjcnTYP5tvK7YmNJ9GJEp0Vmb1zAws1DMzWT7cQ+6x
wwsTwxLYN5Hd0HG9o90mRzEleX3MiZcX58A69sd9z39j3UTYDIiJDH0YpExTtH2D6mZ3exqBxsR+
MCQ33HxDoDKQjsdbk3pFo+RObbZsz9maHtxSKQ0WoBYKCe+9Mh1rSU2Yztm2CrtYO0C7lpKFlZoX
mtEEFAX4anH6QN65r0wuEKUu5E4SyKX0B42VOOYv7708FY0PufG5maz0xs1PHr8LgwD6mNVqu8LY
k0Uep7dBaqnxX+pIRIlrdeivDQ3j+rsSFB1rZZ+2sTsVTh93xZ/h7yfd8dc9VEXQAhGAmeS3euWG
ZoQL9hh84EJ96mROn5EIU9iD11Wdr7qbZmYL2jpCOzm1MvBbB0YpgyXevJBenZ1m99VK2G5gD6cl
ozueGBkgq3tTYuIGSn899X/8tBhvtGzbGKzfdolBAMe7Ew/RAjrBVPLCnKudpSyuylidvKulYDHl
c41qUmi75wR0R+BfNN9ZX7jSFR95A+2Wo3fe1KySiDgIhpP4gem8wCR/dATDsLNqL0Xuvu7bu0oe
HLYrl6IX+SyhsUGD3mi24N8GsL2ocqnDcLFVeBqzDVA7cM83TMqAkLoGUccZboXp1qHDWufWbydW
nsqoDzQjFm/7jwk7OpQo+GpE2vMy0ulUs+tdkaqNbQpxDgnaKL6+trWNq8+vbHLbVLH7vOS8+dw2
xe0kTr/87qg4lW2kUG1OcOrYglOgmfM2rpVWVXoD9dtj/GcC+1jQ+gN8o+yF5GsrCcCRsGGBS8Jz
9pakOeOrRtedbE/yvVo49sVlfCe4KRRoAkcBHE8CfymdTOhWkq+Tzjxkd9rIPHq6cRH2tzjjtlFZ
vc5QTvH/Mj3Yii1jR2V1hxAG5oubwo3Qv6C2P/2B/rWrG2311UgHbULXjX5pD1BFPUjh8R/aiMqh
X30qu2MtDxvLXGFpoeRNjpwXZnnl2MaEzHyazm5+7micUO41c4pLkwviUFj6/04ti3FB+OsjIMu4
ZZif7tKKyXoS2LmcN1Ytjyug2PybLrmsWKylZd+v2FyRv+RrCRH//Rqa1qX6V3a1Oh2sBKsAd7Dm
IQdc+M9ddj9tWJTPChQUOCA/NcLV69i2rXYpsENaoPcQW6ibaGsbaS4OcXobGQ036Ct2x42f0f0W
fQDS+zgPAGEBfaY57FT7vLHw0esqFKbCtO+/fi6+hONnEAQPCF21gcG6TFl0UzqBqf2Wuxx+ttkp
fMsSa74zFBKZEKTj6pOO7Z2QhdccettLH6f/efCcqrj1ap4068ba2vN10wbwk12h2ICD76hmSL7K
4KB1v6h1VSqsMs11rlDlE50vurjzpZK2w6gQDAhQp1I9DFWSm45R3VPlREffk/OlK/yu1ELrwYe2
gi2GDyMjv4a2mdE4jQtYDP516jkpcTX8p8OjYdrNoHmqZ25EgeeaUccnC44kL8qmytGZVFHB7JCT
DfPhrZ1wuS6kUp1rXvHp9DDbGElScQydsn3L+7mPbYGUpdYDOi19rkdE9qKsu+YTytD7Lc/uYbNs
W+uSX/dv+0cALvbrPWTgD2eITmodlSyRyS/LcznjXiU6lIDXawvGNtdI29yT09virUxo6PmSFNVt
Brb+o4CIIgkSTvGE0rvWO/avc+u7KUsOMh0H5lwNvZnVaBgnHjlu51uV5LvlL9Vksey6cDWyJlTZ
UZY5HgpyQydzH6kUwWHW7NsC/vATVVWbYWUya3tvVK0dfac0rxhFgwrrcGaG+JRa8P1ytpHpPD22
eWnJT31GO7xOYCWcJbc3ByOvfoL2485JNWvrPfyyTkqS/lxZxP04qvxxHac6OElIPNN+gk5us7j5
vMvuydIGedLnZIqeFmrhHSlCH5XAGBmlpRLNlbyZo3snAPeHqCRWDYZvlDIh6n7mknJulIq9XA6I
zbSq88Jl2WkP1zEWaHKHk9ZsVSYRD+qLRr1OHrHJRU38Sh1Op01KkUxAmPZUbGH8+ApZmqZl72Tr
hG5EF56EmgJ3rUS2/DYmEFnVtnK4n8NPqxqGLkNnbkFYRtrHXvvyFEg41tdf5v6UmrRmMPr1ujsq
8CbO4aSyfdcPPcm2xdKzb/qeX++TaOZatRc9FUGA0lelvieToPAGZcZ6A15wG1bgpcSgyUJPn1Uj
Li8S4CYz0oaADXJoZv7PI5DTo3F22T1Lzs9dDmD/L5uGIyY24v1L3nwn6XXv1JO/f6mYpBSumJAG
dWHNNfYXMZO8bAJxK9PJwEnvBYsMWiXSN/z+rxcJulUAjr73IlVtxCL3s7vTEdgkl277RW/hr5I4
dXSOfNU+40KIehKxJyqW0LvdatrJHRgpQJsxX4j+e1PZ0Kk1EYzzp8McN0+Tb44i7FC+LbmTaMhj
zzwZp2hRX+3kAcZHE43QehN3I0udz6937Yc/TSVbujxpfdF3GwbcAp8XWINF3Aa4lwdrRbOZmYID
xdBJDzAs4CvCCUqw/NKFayBc1kDKhcNubevtvVv/hxYuAbel0NzMfisT2zjpaljtqr/SgvGsr63Z
LLL7tE2irUfvIHTFss9AaxoMmgXKZW56cgqWEPcAO9BqX6csJkE/4zWDbGHvy6hYe+uwTf/O+3eq
j1fVVwJ8azKgTopLHsu8ZztuYKpqsERZ2nrY0gwUi7kbzd+94b9gCWunPCiGBLQHVJdsf15K3ufS
aKIVOpgqErLl3kYISYY+tgWuj8/e1VUS//fjiUxyvBErjad2iU0ZNSx26gfgEY0zDbqHzt6XYkYP
3+4A9Y6pEpVsV9xsTFRO2FNjGZJiXyhtVd6VQ/vWTQG6sXwKAUeyg4aA4grCJGOUo0YPT92pO/po
ehG7LPQByGG6ayiH0upSLKZ0FMAyANlqbyVFPhOZtCumyoYfrgeD0MrkYv7ihrNkvJXWcaV4V/OO
PjvnGOr2OiG1sVv7EDLzjwZmthMR+QXDsVt37Wc9C5wGWf90QeDCM/F2jYc3NZR8EsO7EKfAbgdS
3hsj25uFChz/zS5MbR+dFyczRWngsfaOyQ1tnFblL/yy58ZzninTWkbq6j+5ZKqBp6LLStQQpW1c
Eu7U18uYZUcOw3MC/Zyvzusx0yXZTPKmZJJFLgYqalGpqKi98sDhADLo2QlhEbu5OSXFvSQmrHex
oBY9ExE4lSR2WQGM0IWznTM4ECfgLDVhqpr4X6ZePPJSnsMFcbbF9sNN/QvtYiLTH5Sta/UNEldh
RdMclKTlabHQUc0tNFxzaFDkQSDtkz3m3hNa52kuLJG3TaCJjZVjDJYnrYFyT0dpvOKmttKKicH5
9e5z/Ub5Qfhmk0saEQJ8g7+FN0mQJDtLH0jECWu4ixHehCWXhd+UnOkX1xfcq/PowWooX9x+HO4J
SSTdVzgKcVY6d+3gfUsRAu04FbR3iJJ/D8+eNMBbhJ1A17dhREEKtObbF4YlkfFJY0Sp8oEAoIwL
hBFYDN3D1+GtP6uVOkxd8pQYBsliwA2AAytc9mBLkm9kfOloRBFXRM5w44SH1jb1gXcaixYYvAbC
hYFV/wPv72yLWu3W9SPN4vvrvHlEphK707CYZZedWk8S4C5RBnWEzk/PU1wAkvf+tEySdu8s8hLO
N8QuELCyPESi7tGKptumNYGU12vaJUsbd8SzOpJZZPfy1aPLPpjpywet8uzkuDxKueYXxLgOu8Jy
0e2eskj9xN2FgmfQ8W71DS9MwcpPuEt/WH71RSQ9H/4Ru+/qenZj/jGW/fphLwqOrTMqbqHhWIN+
wA7kEfvSftQndtZRWmjRIU16Ae/66JKrdAULNetE0Pei0TIN0726Uyyt8+rdl8rdNGBu6RMJtdE9
XdewACWTy8kHt/V3SSpaP4BOoBESxFWOaP7hJ1JaWdPbMikied0fxqapc1Y60Mt8ufjDOiUkBVRM
bVKQj4mXPSkmYXr7jVjDn2DKB/zhmzD4Jt2jAR0GHe9qw9Ii6rGzH//fXbcAwQ4n85+QtVe7fHPI
ce+FyApI+utu/1iltyQH5GZHcVArCPCzomeBlWq7RSRO7jtQw9UI7yMM8qz4XB3b06bCyuyZkzko
P8r0RiLSN13QEmrM881oqn29aNQcxZJdjmipnFaHPugcaObrB6GIhHBLZ2ATmmE8QbiVlEmFhHrf
TPRKxEEyEq2Tn1uSEgxlyI+KJsXewgt2NhmYt9kKh9InnMHQ4YxZ8r3nFemTf0bvBZpq9Up4i6EL
NHgB9IPF6WYRGPME+KQ4xEZurOscCHqEzHdbAAR/wNsY0WsWBTAZPLGc/XD6+hXmsqRZo63Ecfoo
ZAw6EnkM0Cro7FrRhYnAqOLXE6qWn9lLHEkXbo13HvfiLy5KCCX6qk3ckxBmy/w27l1HZT/hr0Yx
BXyZuoXzz971iORerHTtfyJp8p4gQUdb5TqJ/ZVDPmEUr+ulejRdptsy0s+hhRdBSithWvh5DXQ7
sDTvio3pPdr1unrgMrbwVGNb2qAXiWoDabFXhcCk2FR7Ls5vpSt980i+sMFd8kOVee55r+xU5nB9
UOVezeCrcga7qKd15il2i585pMReUbu0BbJU7UxKkFw79Ra4rlGx3zT5X1aIJPcLOWHeZ4Su0GtD
kSQIp3RQW/ViIKoEtt6i1uQ5G33WJfkGSDrjxmYgIEmuw8p6LGidtStOGx2mjP5SDip95rcxzeIl
Xwl41KtlwwAMit5kCH/Qm3fNHgUWiqjv2iPHrNi1OlpJdy5lKyynwTOhAufe3BYorNelfjrR/9Sx
JoMTT71h/A33JU1HPuNC6ZkxpxH7ijxfl4f4eBQrM0oYnQG5a2jC52itq2Yr2UYVwuhX3WloVWkC
cx6/G5gd4LmIwJ/LFn9mTjcdYUScU59UDsRG0MwHKZYZr+jtBCRAjAPoo/cjP/AE1eLlqLI8HXNN
h4r0cVa9fJFjnq8JQiGmKtIOYEkbvSQwnE4wo4G9LHth7YHZ+unwi4FxWZyLj98CrtyOogfYgCAW
Ys4Cs17cwOWG4D+lCDofIElf/WT+04tBllHe1Vxy9NJ2q9DnOS5RZ2nsWOC6YHucs/VHv9rqzSJk
myKv/9Jco8l3M8lyo4R/2YtBqQkJTa6FAeFMqz99Dg4YfxVL7E6onDpjdV/6XLRa4MzW6sG+42Mk
f2aCBwvr/KdrpJy+UbN6OS9aRVlXHpB/CDwc+ZlQqIexHXB3GNg0fTxlJy55qW4SO50mgsMnNffE
WAt5qgmhLHFbeNpD9EivuV/dX8wRS1xMjiz/vRtxiR47yslqDy/0pILDPJ6nLZdv+PGloWLT/qPH
JYrpEgqsh7xI5t/UovXwb2If7bNQnqjr4m0fKTEqF3MCThVGX+vMwYtlWA+Fb47/dIKGTCDfxwBt
tBl3KE/0a2dj4HS7KEu2OifpGbuyLmVjiE36EtJvlXDQdsHLdn5sxat/jluH+DL8rfqkPTrH8JQ3
EL0akTOJZdBbYuQBIRsVGdhOg9vyqk3OPw+ckRwA17UxpreIJ2APRXci5LD2y++LWw4owWnxQKAr
nCA1RVe/b1DS4BtAOh0SWPrf08Muu8VkACIZPmhHq6Vpqjp6sUs+aMHTvz6QxTzWQBbk5wGUPxCu
sgBM5q5iuE1BhLKoGhQjHMrDP/7K7Ig1UsizAAjiGcJzOb9tOno4rS66i+C78y+9uRn4FUmvJuJC
+I7v5uovJdMNnhsfW3RWv0Xgne/HO6af0iN0bRgFvelQZoeTkL/peNrrjy72CPkmeCtkgpPjeKoh
UK9YA/aaP/0Y8LrZ1eX4guKTtqfqLWFTYewSj1w6hKykTNIrQqADLEgEL2B0oygxAHp+pG3T/nzb
w2SqzD3PJHOoXdwhj4+IK//O39PViyQi+qJXQOgCqH45lTcnQTgATeaZ64svbiFvSvWiTBbLeys8
lv2JpXyAclJrlXgwyfLb55FnpxQ/8lo3l+SSoq3mhEckiKV9OH4BpQ2+z+qxvhvhKLlZOyjN/UsS
HJwJF8ZmEpyzOfCkG+l5y5gXtoiuzQ6JEe0MxiH5CyISwDygrBqf4LZ6285H55+cgnz11PqJcauk
TVzLOREpYlCy9Dyc/bmpMaMFpt/VhbgJE6QDyVbICFdf9OJnr3u8XAEInLvJwyd3SMgQNimUfooB
BlvTc+htRNNsonQSq9c5C0hpjBXsDoWR6UnGvXWm5CY8XWP+gt3ysku+lmzVz3IDxDRJ8pnS5TD7
SgVzaZdE7XzXJjVXoMj1Av2F11f7xO+sOGZiXTYsmAYu7N/59QUXMHU93qECP8gIFuWaLAHr96RH
x4FqO+Hk5NYen3+lnpCRjnaMsW66D3VryxWA7RXEOxY4I4uuTknAdRsawH05y5RxdlZg5Jdbmgp4
qBvUcvLstAaNFE0k+JcR6ysjn1ao6h7bsOoYAB6cL3964NvrAUynPF8ktokYbH1oUdG95CqUwdfq
v04kDMbuEsvQcYDa711tjwxMUIc0Mz2wa6D2GmFXbptH8EMwUsPyA36KprE0hZRPJo/5jsysP/T7
r2ZBQnOl7xMrRakOBTM/vT+clyKwD75kbGF17TzBlkw0mtHYTr/ORKK7QDwlJMs7opAFWDgOGm0x
jwYvl2UTd67l6ObANyrbIluraVCoa/lSVyON8zCe0CJkdeNmG8y4yTnG3Eq3eOENVONdNWVCWOsU
xWFoaG6HRX+qFZubUzLyfjCtepuWDss3SsUILPn1sJZio4wQG7eTk6d3zVWHcPOgpsyjoaMXtlUP
Zm3gp2j3fiG20bVyISnVa8LaNW6CQticd7/Z+EJtYpEES6+tPY1YuxrCwfmYNbGrkzmLsiXKg/Ac
HEDFtLIvMY6bg2tEM3te8dvHQygV8ZWE1v/jpylHPETJ6VtQzhokSDXeOnyi0LDql7rV+oP77ip+
Ce3Ow7zolFbHn4oh25tFkC00xs6mdD6FZMfsKc/a+rRbrPN9/zEsipeyKN+yon4s3ZhZKT/O2LFc
uDoocuAbNu82D4T7Qgm7oDxBDtm671TBPsbjLJmgBBUaQ0ztcfUNsptsT750GmUKru983d63K1wk
Npf3QFq8j4QbNFcI6UJE6vKfit9EcurkGWUVSR6VoUeoe1AyvZuT2oAwPtYfI5mRwUF/1NM4zaPx
nUUHhuz8p1mYA9QDNaNoo4b2U5H6r+7V+LFpVd0FXhZVZtCKS+rjSi9CHXg3oEZMvnwxqiliEifa
MDCdTVyqhG/7aLGcbbbk0GEU6BVWUmhF5J3vT1jBPNuI2ImUvOawPVI10+qvVSzb1TTUfP+wmgVs
2Dr99VJJZUyYweLKX/HNbcXiH1WzluECYCWg1SNMaKnNM6DhmieeK4VL6gTauwUHlv01HBPJUaVT
qXI6IcJ6xIxImHk1Rn0XaQ6K+CaoWLx2YDYrlZjipigKiXCsqz7HwzvZvhsRuuW/Fb5oCDwwwZIk
7uGDwUnGmrzTLk+IU4jnHWjbsjQFck/oSyk4Iw2BRmFaBlk/lKONnObD8MqpW2PwXUF6l/FEm8QB
iViR2m8uioPTf0+rJ8SKaABL9ZsFu8sM6ewY423y4jEPOONHr8gCx2jPkrFfmsxRW/5hhJ0he76Q
b+LPE2rmDbdXiFN8jcyT08XaYSiZGB0QtPbvhsWa4UZe7rHKNe/Pv951c3v1Cp6VedHA1AGQPata
4X/PImuTrxEdF/pJ5MhRAt+1EGGM+GtxB1CnFNdGpU+xBLXPkScs4JlLiI5buNPwssebycZ8Xgv/
E4zCCHusxGZf9ReOO6NgJMIwDfEf4h8lfJMFFChZk3TAtyaVK/iKZlIOelJGqnohw5QsC57UucEy
MFtbRLzTfZ7t98BrLM4Sht+uZh2KqQEgpgCQHhzt3/OWKUmXJKRl3R/IhXyB3NJkMCacPYdCpah4
tGVLTdqZrevXgAz2r8Qv3UfH+wmfNqSKcQkbGzj8rYfffqIw2RbJiXRn8x37DTbcVJGGl5s9u6LE
R4h3/RewKwHeAm25cWUYfsM3FTl6jnG2C/w6c+W+w4I9ch/cJ5LD12qXx8K/h1/86tFa58oGDVo0
hIIA2bAIMJOyJB/3qrsy6K8MVVag4vQ5eX3LOD0gvUP75mL38+K540ry7A/dn6ts5Rc+7U4PulFC
0yuPmePZbCLHHkC9E4IbVqE3lb4CWD9Qh6V2kQHjgZzmNH+SMe6weNMb7VO+av2WG1F6yX+f9XEr
sFCJB33YkvfXIHG2f3CO6UtwKt4JrFW8TP2w3AVxok8oLR2lpV7FWjj90J6MnD3t1Sg2++efd8Kw
HQpEntuyKuR0bfaZ+aabt2YsStFSc6GFvzaiI/pupo4IWCDAKNZC9r+dvea062K5fyYFHkBhE+DQ
E6mDPck2j+HpvnFJL1VH4PsO1K68ficEPNZGCDy17Xvlt2bMUd8UE5TvH2oPYHeRh8h04la1lkzY
z4iHFXFAw7J18oyD/nv+JC9z97FOoYjesO5HEEsFhDzp4RyvUVopZt8uxtInScpd9plnYRTRh4r9
ZLEYDu139qs9AMcRtdwyYgZDkVFnwHdwg0I0iw5QIHdeB7jgBNn4qjOGgFkkfQfco5ZrWH6YWTBu
q6HXQFUre/5Qhn3IZw6wxVj1vU52MU8YaV68Xdjv6IlvxhCiKaE7uBl+WlF3AwMW4k3+BbyRtIRP
vRiwyXNJGsabBRLtZHdJXvVzWxpYr6DoWXs9N0DeTScjQdQl1RwUYpyNJSSVh3zHCDfrFHrPQzoe
lXcUbegaZtgOaRg7knF/Zrjj5cMN/ShLF408ZtG01+BE4YRiz9mfBtSOIlruCi+EyOkRSKrgVy45
CTZGtvXwWExH4MgoSp9MY9a6vOAJpEses7M43q4OhQ+K4yunhIKPfmtnlfxA32G8Y7qD74qDmT6X
LcUEk8xP1GuISAvuvYJhAPWL/Smpv0K3D1+aM+F4ZVvak9N8Sfxi3w06T/ePZdox8yrk8iQxvz7I
ZHZkR3CCroA25WnSdufYTR0gxPOeS9n3l2XiQfGSIacAzDqy1kL5Q4+cRo6gJpZunKxg3KaDBN6H
hCFDzXpZEUXflNtKF66JX7jKL62ytZoZcWSs+Dwz7WY7r0kRfBx4TyEsu2oYT4Q6F/k4y82KSyeh
tlNg/bFR6x1vuf3Punc53Tnwosw31zefRTZBVWmwocwYFwMNIhObuKh55mpKqFKXxlFA0OMBNAeQ
IkHcF87RU4fDkQ9KbOw1kv1Ps6SsCl43mRFqpgJzCJrFA7VQesOPONLlIQ9umcHLK3zAex5jUdmM
EWDPYMJ7Zsd+B/I9RN+xAxHE1imrcaknnt8cJH/aZdt7Sy06Aqt2FHA9JQm36fH7AWpxk0xDRP0Z
9Ze/YULjQQ3+/soEI5IqIi8m8jAL3LeUl+wo4jnyFh/p/gz0wz5B1SBnELTWOwmpX0aKOyFNyX1c
GlHgPZWBlBb/Z8Z28GxaprDMRuUP5nQ3GFKNF9VoL6vce+oX0X3gt+/c3ILWnYj+caRxWWShcHRh
s9EhKA/lR142DLRHxliDRUyAiCjikNCgyz3x2XMBKFlfLOTr+o75gT0rem++Z58c9GbyByhGgSWH
thgGLKSruZvkYCRBHLaDRAMVX48iJk9igKEYsAEEAoED27JRPYoJ5iEZOlI/s2ZOfJWx/ZC9/v8z
kHtSRcnV6qK7kiyeCwRdHSexDCp93vhDulp9CRpn+JIAIO6VimgsLLl2UH1x1xJN+st35hCLsxW0
+N7QWAv7WL9FGntz4StFl73YMP1Om9wbVt3KgLLznJu1ptSCE6RpToQaJY7nHB5QD/j8D2yeqj1+
SM0xcPeRs/f7WIHUrMkPBEiSJKbjPMA8XVtbs/GzSXSX3u+Y7vAxb5Fe7jROYwL4riWM8owx8B/2
fRmjCFxT89UtMW2JpIDrQ2M+kVkGJ66aRTZ8pODnRjpSZZ0/VgUxqrI9JbbgUo0EZq4fGs7zD/U4
RQRL6SEfdrp+jBqx1xUs42hkgyHyrzKV0x2O2lKZpwYpFLH9QmBk2xJndUm9aSnJeLTKZtGOS8Py
gye963risQy193AImC7ZOBIFlhY297pfEawIleg2a84J/VQ7ZSglgjNFaIdDzvhcPHFtoaAfuELx
LTzEt5Qy7gwczwr9RfFSPyDYXPCsy1Yctv/+h+XRFw9142Z1LrdnVdpw6+p2JGNsn0gcFg/TGw7k
n2Rhc3uDVflQ8erOsm6EhoOsjycmeRabEhOpy8jf6XZGIRaHIo494k4kR+4AB+DtjJDVBl8OukHF
soNXSiOW2S9vy7DWPnfCkIl55oWgzj90r9HuCKS4RR500EkDigJgahWesbhY6y3uOatc0wPoxQax
p4NQcNBhSIrfJg1a/QYK6B5tkwm1/LBU0t1fWHXGA7U97iJjKt28hmzxId1o3xA0uDHGwPwN/7Zl
Nv+Z7TbGljTmDv9vWjGC0KQ1Ph4WNm3+rUrkYoiTzzXn/MacZ32r94iKFVy+zk99bhGv4KGUVqnC
JiIbtv1qZYuGGyl/HRvEg2UYHgVrvfzArriZ0I334J+McAgUlJ6Va+m6ZpfU44atcDh0W/PN+88l
HXteeoLhPvIEwtB6jt9k4ob3Eb8BIoYUVelOQNQWHMVLSunl2JRZT5pJm6BgWXiOF4IIj0v8A4hT
4xk9oAGMiXdz55yNB59F59TXz9sUTW5ldJO86shSP14sB3DjGMcEsZ4pTMpKfS/NDC8NpFRJuEbG
xfKZ6WXgYhNE68DkHphXnmY98pH1rad/Slvlnls1wgXVAsCLWZKNDgS9ZdCXiAKDgXyHWVCECSYw
0BO8LryH2HaezmAONQHEUOpTPfB/YAxe384Bs09xTqc9dYP0dHbv/CXbkeNP2AJfbPeM/ahxwZ/b
aarbarCHoB2bKBIza9JxTAJCzl4IHDCoFWaVtVPelnNaIhv4DQ94DyWf0psri5rAOuZNWZakmOKF
GjC0w0RUOg3Etj2QL/VGuMXuQdXCCg9oJb1GjU78kD34SMynWADvkyydzwIHPHR1djjHGFo2HcPg
nUmTpTkgoppmzMNNh9cV17GwQ9Af7ib8CY07rwecAbFmY/E+HLevk7MYPwq2x3H9Cx5iCBCr/CXN
vVw2ec9z6GRSgrHGLLb9Er8m3Z3Yr4pvo1pSlZC2s0vniJ3ahJgVEgbqrlYnnatB/apGGfQyRzkR
sFwFUiT0Ri/ed/Zz1Se5I7C2cAFh6ngQZDuuSQyLJphagndiUKiOnA4FsP0vsdrmFOo9KlGKdW6Y
Ba6cl3dvC2Sq4fei2yfP3SsjZL+OjTbQjHYOcdWRTcWun3c3Wcv6FLl8o+UCUj5pKK5g/ZXmoqXH
1WSKa6DcpEouxILw4UFDdt24fQy8zsok+MOeIj1Xa+cB+btfPFkxlbhZni8rQCHx4iZoQUgaND17
7E+I2XVU0IJiPrVGrXhiHsck5B4euytiB3yVxsm3WplDJM2JZWePPglFk8k5FzbIhz4KGL04+LXe
JW0sFmrplcHalKSQ8vDhY7pZbh3H9GX5Hz8ixveNxcME9KhcTzmwlW2VSDphC4oe4mCSnA3qHRhL
JyHDelo2x1aon9oj2IVk7j/885HvoO6JfgH+TA1Af2meOODuWUtk0q8OFs/WbRStLyzStgqs/KVV
p/+kvYttkIVEB712UmjVDSAoLDNpYsMmeHPZZHNi5B6rJhTS/6zVxVcyFq0H6wUh7B4Q6ozySCYW
IFrxlaZC/3JOO7pvzDtwKyiZkjT3Hp7urZjSFhhHtNjAdo5dLKK5EnqtVLitplIVcdnbPoNJC4IL
gkJIW6c7w5PT4n/PRNzuwBnejDuFWQfDB30VBIbIWh6m4u5ngfZhEfzdS+2I+oV2S5LzOUp9HAEF
KlcRlVMTKeCc6HCPeXEDzSQjxkfpfDyHwDAQ++Fxww5kzDbR49nLqDgLN5Cqc2B0Zsvn7F0RwjUs
1AUhW0RU5TTo+WMEdRgA4NiVPWXIQ92zM4dWPMA2bZt2jcdBtggxBftp1v/nJsmoRrGiQoshJdJL
VgSsmJTIaKq/xPLUG8Dmc1yZ6Ku3bHI+e2b3wm0vBil0ASuN5vOJLEWH5MjOFKZIC3J9kEEreUAT
1lJjcG7trpl6GKhBDpSnzp+fOWC7cIQzfT4hgn4hd0rxYIFrqsdQM8ijONqPgGSWuWPiW/mZr2//
SFgEDc1n12B+AH0s+DrqlDH4s3jwUWhS+aj8rqzmS6LyUKglu5rsYEKoABRpMWMuFTOgHt5YtU9E
pCJM0ppr8DWtsrDKSU/42mhXd0CcdldSnubBGEcyjmXmQ3G1XMSEWc+se5FZwF8y4HuGUp5FoQLc
oGYmHJhQaWD3AiEYn47SLEXyL4o6KO78m7wzn7zZSTSdR3UqAJXRn/lApg0zSfradEyhSZCZB6rm
afE7cFJx8MSSpOQ4UlkLFZYMxuXvMVaA378arz0VPuplHxIVsxVCTYwvPdv+3QCPbl5aF/K+MId4
9pJGRKn4G65KnwLwOf0F0cq/mMR+MoSszY2n+hDmVICIb9cAK4htYeRZOmFywO2CXivDx2/gfQ8j
t5LKHo+Z+Jl7pNhSecddgfhu8EsgEp4EBIsxa4q0bRzBbfn+tN4NU7dRdBdary5FbgGKe+KyNbBz
G/5JL0HWM/UOpIbrhGkBQ0nycvnR9ax5Xpczh7b/cO7DhAygK1OBtbzCMpGycV2G13/BaAWoGQMQ
Ky+6ty+dzWhTl69FqswwqCGf3gVXUfDDlS7MgbdV2Gm6D+i3qSrummBkgIKTy3Ph9EfPjdOxGu1U
VkWo0xc7ZhoITEu+9BkPeoUSFOP/3r5T9efqdQDIg5AjKxtuZAyZKg78pFbugPHBmxqVw8Zr2Gau
MDE6MF7M4eQpADiOAQxoS6N/DPGGzGGupMZrF33pCr5OKzrTbwSTQwBX1UUwB8QeAx0D4QWHzsXO
BKLeABvSPWnRfTgtgfE3zQseL8O/BtDYy9NQ6ZmbCDefUo3Bse7qdX/HPYGzhQNrRs5QWC949YQr
z45A5Vu7nh1pyt83MLgclL/DH3OUv0R1imG/uQohLJVZqiWxLHSeJGrkHoSDqlS3UBghrLnCIMGJ
7Zv2NqlTmhDDeOODm69zqSy0SEwvc2DWT4V/L8pTGEG7uu2D/9LacXwNUZywmEo6Of5HXj1Ut42P
OaAfo7Blj90HHaeNglSaKwuab6k14sL184udltxllxBc9l1wHdeSy2394t5wtHJdudv7fZwx5sqy
fRef00M8P8NM72EmsGjqeyKqqG19G/bSW1CLxHb0bWE/aFyzvFg7F71a47pnW1L+buDJ8Uw0Zas4
/FE/RmgaT8uxDYeJHw8lZak/4bq9Ys6WZ74HFSo/022dRE+lj1+VyojHwTxTOgl5KYaQbPtEeQDP
UKHJAnO9V5jtaSfjvX091uZnAMzPat+e3lJJ7n6XIxlu//KvQplajGmv7xVfJ6Dticre7JUQ704O
SszSNIcPkSUxYEjxugq2zo41UZU/cuo4Q6e7Sc+2BjoH6gF8VWGEMkzwG1df2IOkmCHwr6plPi9U
EXqmcRROXUwkF4zTkzqap4H+rm/iW3KKybi5d8qJq2Xbu9QlAzwmBMDIzM7Vm0OQyX/dCz2FBE2P
pLiFdy05z+YsvZ7owv2JhelHTb4JLlIJcM3eP5v9ECUV+1WKvY8nJjwbE9ItMcwNIUR0rMRPBQmi
e1YrVLNUImlNIsBQkyrZGL+x0s+qX1VZObM0LUC6xxdEwYCWeXexUfXWYCvNCrk+WM8dBxlWC1q9
zNOy69LhTHuewffeUZazK7mCbhqab8I1W7DZDZiCaYUvDJ8vM2Yvc3ribVHKvzFcOY/Ti1PqLR0z
EkPIb3rovDkuqKtU9lp9YqyX5IVBU0xgZ7QhYETaFJ0+5p+pbNlMjf54O6/UaZ7GYww8IfRl+OYa
i++WRYE8jQIkwNiyjIOz46qnfiz718pmlRQLBRmwin9qOojOXLXzB5aOF1TBhURs72JfyYboZj8K
/M9i73bu5PnoHxeBs2GOLSwnEbuwz7mQv3cIjP6LUamKeCdLS1M5I7w8Us547ATL2H6GrucjvPT+
4jSchfRIiXeNVDeQK8xcspYzrND9Yo4L66n5SUThPPPSHTD5O5Aw+HXEzveLbl/fII/2WcYYB+3M
8bRto+VrjCoD/HfrkDp91RDWconua2wUl0Rot8DXLVB+2WxCgUZ24rcxtsETZj7GV2C9ciFQLXGH
guSSkxw/g+q1jHw+a07NUJqYZTpXmfK1VkbK2e/lJudGeHk4S21/PoAWjp00bdflVkkY5Ad2eKto
fpjVqqkdc2MaxkZ4dyuvfWTr+UagM2jAQP3gWI2kItzvRrx3wNQeaWC4WHNrKFICTEs6rIpr6/pQ
9gkh9Sx6Gp2aCKOLnlW/QCa1gH7W0EhyFzMl77LuXzwYzDUDalnHWkaKEFv4ASxU0Dn6aLhrP6Rt
FZY6ggaSoJ2LReTFhHkE2A7vr8GgI2kLhM0r8szw7Miw7QOi4s9a0SCK2TLH2QOVRVt8fKQ+5iE5
4x0/0OzcRV7eR+8nciOXE+94TneQN4DctVh4sY0i3WMQuwnVZAmOdQgKNqCuV4IvESxV62P5SZNK
we4KiZWX9YVXyCyzQB7dmpqFHa6bgmVaQS8RkCZ1SappNfSA/4N35fJOEicr58dviO7kvRzxukat
zH2aztuqrMUQ+c9uVw5l06QcqQN0ycTWwW+U335+Gk1q/OBTFAF5F1TLsdFYwXesdhDbZGEjnGUF
yC/7VUTU9knIrLj+b4tkXwMp1RFR/eCh+SMrcKWp+p/PGP8t+yfAaAgDHrsDfAo+CBZqaY2QCcQq
AIV0ixp/JgvoUh4izV6ZwkvmgGHFKGm/bSstc6MktOAztIHigkSIPSgqjms5HjOIwIDNFF5LpSsW
s+ZPkTIjFMiPBZr/EIfHguSxUgAFff5ZVfCNjHjiUeCXhIXPZM7EkhPdYJBTpzbsu/z+3RKiPHp+
em0Nk2i94PyLJyN+0w27GVneG/jqYFw4zm3/KUwQLlPkPkiiOoFe33alCAxFzGPZ3spJXx+MCixG
X/SB3V7s7zGkRUv0rPGUWmsszg+cEmm6JZRuI/aXmiSUMCtOpoV1ovSVgQXz2C8z6NeedCzXu3on
KHVLfvM8/Sem4Rj0WpHXKYwsTgBVuroW/ubsvxfijJ8BjyTo+bVFuFdogo9pbCCeFOpZ0JwEcbqW
0ztpiopMbHveoPUXuI2R5JjkmtOfkcOvKhwS8fomTvKR529azObAMp4l7ySjYa/d7fCikMJ8p97p
OpVimIe1CKm9qZZz87ChdBEhu305K6RNE0l2mOn7e9+6E6h0E077hIxr+Z0orWgToLZqvaJpeJNx
N8r5BxeGfu36uxHK6vC2fAs9tfxeXf12votBAEc7cPGs8d1IiHMcLkp48lOxlhQy7P6mhTO7DTVf
XftYq8hvToH46WWZFwfQij8lUZlxPkc1DZhfs39R+6UymvrsG5U8C3kzJm5BTGjGzU8qfQGyTIGY
NJxVEEdeZySimOhb+iYK1lRomirSgecQML89/eUBPwtVGHMjk2w2UHOthHRB33fyAKqBCHpkIO+P
79cvmoorSN33FrIA3fBYpdy3IHuu80i/iBS/hhDKoyO/CF7yaHoXh5BfXvzzmQjYMH/lVc9/K8jr
8SvPOnCmItJJPkDE6imcHmUKRETEn5x0MRIHfnz8MI38YmSBWtRPjV4xlGL6LsbF2tyql/EaMJ/C
JQLG6HCmgL8Xcv9gcF1+AIqDRftO/PJzNhKtF4Jv7O0Gd1B81XQm/uITk/jpN/MEan2L8QxxWpRT
n7Hwq4ajGuaet61+VBEeeB0QK/T9mQtTyjEvWvpgV25zKSpwDAw1QT447BIe1woHAvn/KdDqw4UE
5pbGmLGw5TZUvPis/XOXGhEXN3QoAPqtOwpuQUj6HnRNLsbu9DzyD3XUTG+cZge5xCmAToFjlERL
4pIlmS3SwsnR7Pbzw5GITGGrjrAjemOlB6h/ZohPW/qWr6HhLrnw+XsAMsBRPM8lBjKvSRL+kFId
utysV4dRYMQvNbBJJdc53DBsatNyIryyBOoujYg5pLTCrMD23BI+WAqCqdgLwnsdpbcdoUpGO0P3
XUVQvnsceGVDZUkefxsBtRcVfu825WINTN2WC/xiaEpNcbRDN5u8YnOmfvDSMtRlT9Da/823riTJ
9/FP/GPxSjrjhYe3ndGpSFTid9+KnHt66WRXQVLz2e3HjAKlGIsFBdEnYHkP9L1fhdSYgDtO3tv5
r35Td/nNTKOqnIWtQ1JBYU3vwJiFF0obxkIEl84jodmIIG9T6AzdI9M/JWXE81d1iN10lOgziXO6
2xiQ+OmWpjppIiYGf9TmvOiOp22PDXD855JqofGMchobEZSe3BpRoiXW39f0VmqT5LJvag6TZA29
Hn3kpl8ZDvuZgqmMPtg44+2XYY39rkA5JiW+F/7VbH483DXmudKBpfW/i56Cb0gErEe6IptBbfIw
kO3Ip8+o+v/eSLfeCC1mJvljONRdlztUhekKilVvG65+c4kKOW/RTdr9ziEXGzpa7iBoD+FDgmJN
I6HRkXicH6Rj+NwfTuAuSOAyWc3X/3+jW+c/JpveEe4hjW0a0DTjw7y59HfjhmFDtawt+VSRivjh
NNZ7ijmhgXD4VkkNWC+eRnjxiFKR9G7PpouHyIQq57phM4QWXqXG+bPK1Z42TmKeYfQPQ/pXKhKB
9FQwBIKMzjns5e2Bxy1N/SYJqnBm81TsQhbxU2E6ja5wHnwRUtaHFZjsOv39i8H03dezGLJGAiAQ
/uMFh0MKMNt2VD8tXceNQNtxi5G8yywn30azKdXpFkShpH2y2I9GPEIed4JJsnoMoG2u0UGBOmb2
C3oIURU5jJkB5BnEaxNyc6PlEomsIfqSrxH+sOt+xyy2zb+4I8sti5M3h5ehE3ZFinTAhFgIr7yB
jXvQB44oJdleBjYb9IuD+4M9a1dpnDJ3VkYPnbMIRH+U3Ed4qDJe+YuDcP2ijvqLwK3eTSpxswnf
1p02wJJGvYKDQylishN8ScQSNxpsGdNdHynU6reQxd83LxF8kFnSyftSWei898qIqGnTfzCe2HCJ
fjC4nO+NNxrdfjtg4jboHCKxGzJkq69xv23fm7D3Uy6jdjAMc4+1IQCyrOmf+sOS/7axS4tAWVcS
wlY9w/mHC6E/ewbgNUn2dTsG0jvdYUalQdPc/J8KpfJvRhfl/LMBscAqN2FQxTiR2tE8jU/0XpYs
I+B/FyIJC8tFi8kLMSk8hPHzC0g1PeJr52u9H5TZK3L/dlirVgzv40n7yyLPKfvizU4JRHU1TnWu
owfuIHboYTD3hqvTMZxB8AuRL/aVz8LTyozz1uld0kuJ3Vp64Fc/X2qHJPCS3F+wbH06HP/nVZQ2
Q+uFDNryvNpu684z1K64twSOmBS9rmHFEfPXy/CIoVQADtAALOFwyYFKsMYuodpmYsP3rL9rSH9L
BYrdURVwjGiwcVsmVPVbvto39ghNSh0RZ82r3DtM9nhuX8vz8SxYIJcgFdngxqcw42Nh/XNj3l4v
1m7lFdSkSGT4wMdYrRolXyyhqyPgOtkeq/B2lKjI8DuEf9v2HMNkOX8u53TWPb26WF1W3AxRHX36
ZUntoE3bml1UkFTknn9vrF6jHIRkRubP3pkrFOWY1P4oyODqbjTamQaiKfZxSg9Ct00R3NR5Ocej
4cz7MHWnPF+UQnhGeEERQIbEXA2iDYKMOavTGENBJqCi2DmpYbn/BmnlgXknuhm/6RsN2Y6OcORt
fxf5plfwp/RntQI1hM5nAspYrx+7KJZthTlluyqxZPgM8tuz2qmCuq/hHvg5f0keiBPyMKlYS110
iyO5k+1tP2YRQwS/Wk+ZtA6JMnEaAVRDlNyzCIRzWNcE2fzZtPVvEqd5B/2FjdYEbvCu+2OJXVSn
4o+9C5nJWl3H+f/3HayaOTsbnDrOh+Eu5enfzFt2wuPU0jgYD6ALiL2igBUJfs+MT4QgaPK3WetG
/t9GoCiAIJPR7wy4AbQTczp7SGCnDLbTldFDWPMkH5G6u3eomL1O0aTzsxIgTr6kpkhhGGNPTkvY
b0G3kMQCfCDbLo6dy+k50HooXQpBUjKClEUcgeVLsweIWlv2rB1N1VMNeDHOrMtaNjpXxsk5Gpbu
mmqeS/q0zXZihK854CogAcAQ5DUD5ImmpHw90lZTr5C6K9xp6AlunUS41mn391+3Lk2I95/AHz6h
lLBlORzzkGTNDuaHFcmUfV1YpnolTXTj3saikVHtVKZ7cwZOzzV3SEfKDxFN68DmWlf8zbxYr0GE
0zwtKm3Q6yo4GcrwkOqR0MO+qEU8NLz2/OxQ3iSukzqnIiDxH3nW+pT75JripPxHITlcBPPeFfiV
38nPWayV1rqwUXriDWVY3ao2tDpGW7QWEDt+eos15RjmTdXo2jK5YpTzaLmHgHhOYxvm5zg4tKE4
1SpyfpD7kFBRWhbfRXtDjzLnCCJDi/KHn33aXilh6PzDr35yC6v6fAmP8i1v6ltEmm9xHnAdfCw3
HauTK2iavkPiryF3eIa85YqG08Ay7dFOb/YnqlZsooFW0pa9PiMyL9uGVtFs6FPT65m38YWDLLy0
eNAbKAj83UJs5XZAVAouhTiq+v2m2dGjtcQKUQ9OO22LRfjbzI70TmJ2NFImz1Xb1wb+WSO9thUV
qkTeRqYfMXAB1ydfsUCd3bQzIVWL9b5+P5g/Y9RSlcmTJZ4vFEvEkTYgXvpGm10Y3VVv4aKDpitu
5eP+2oIkJ7Ncu/VFxwHamZZTk17qGeM65tUV3yUHjZKVzuhR4AOAySdqSZqDLcX4PipCU3pHwSxg
GWhZpGwjxHg1Vh68kVrfDnBW3smEuASSevxrPusvA7MCrcCEkXZBMMK6InzZb/bQV4mwYJsCC5TQ
0WhwDrHe7XwgT4JlBszHXB/ALDZ+7gqvQvtXSSU1OvjMWGDMlYsl/4QtrJ/F2Cy4rgZhwQMCoApB
WvzuJpZI0T4XEXWJzQavuqnng6sBMqd0dspMFKWVwDYA+uNmS2+akHIMLSrLGrUk7eHBcjnt+8eg
KQn7Q5dXzUoIjNVTpL3iyDqAr0TYX5PI61KYuelReIxaw/8U3rpyIBxGGARG+pdLGsMxjecLHdBn
N+dQgia/VVRBZkejM+CaMdgvdVuxC69ATJZDobI0tum7hKEAUIzwEeINOs1PUaeUPCc79x2YmACD
kIbqjfO8fyA6Edkpi1gOA7E3Q9WXE3PX6DKbQ2lPjxUiyihOW/gRyHaeUsQGAmO9bTI054gFuTfm
qdV1e4jCwk9vGgPDSc3Jqs04a7e/+FSHNKEAg9IdjNedz1flMIDq/f8Mgmr10fblxTeYKGLE20FY
MhtrtUzP1cphnd83eTwxuPtk5FqB60V/iV9ELdO9BI1G1INFivohKJ4fTCI+elGHZVEr2pDAs0Bm
vF5Ob7k7rt42tuJKDFO0FeLMSaA46gmS2RzKnl2rf+gWjfiW5JZuk2fgHev4KWB6w3wlezPvdiHG
JkKJlLaOoeJHHXxdyDLIOdR4QpWJudwBIIF6r5fgwOedsQrtqXQJH7Le2+fQd/DA0DrXQeqUmiLj
c4wiHkDBO/XSPXxMGwe+CoQ6OzFhD3bwNo3roCokJkTgLmJUu3xvHUNuXAIMHIHl8zn8YkvWNIZb
D11fBQCrDq7ox4VB/FKefwKF+GhznVDHaII9MVJnaZq+I685fgYd7uU8Fw8znK3Cik+CWMDMZdOe
WKBAgw7ZGrsNW+DgpgrL7JDmW1RijysH7KzelUjS/ic4nkO965TYLvhUyE0OueNfszSrS6bIZoF/
Levn/7BjJR9CF7WBeRiRrW+FklBGJFyGccckb52aPxA5GvtkeEhNwiFT5lXQKORx4SCMXmxwQ+i2
nA4VHr8+ztT9t/BYpaED0kGnZUcH18lZJTLU4vUYDhAyMEHYlNGgkD90aDFMtcBYWkCS/wiAFTRs
hkH7Ql5htTOR4OnSBKbFb6ksRlqbbvWJ8V8onEwzzmefk4H4a1k0I7FdWhl9uTvM5X4qZQkSeoi7
oh+kdD+wILkCSqdk4ejIopors1gayhevsT9B0ipp/3HRrSJ8OIo3JT4k2U3jWVMU1IGKSqGzTi3b
tONRz3nOeQ00PUxlWLZzoaAiAlxDoeyvZeCzyQOuAIS7bq4cyr4R+WeuXs757jV+WAtp/6xutYb5
/hoW0s8eblM5bc+Wdajzx+kULkoQkV1eilJneRTa0KWJqn6tO+el4JVk9aEp/E1HmJd8VakJjBed
6OH21BIcPvtKgD8xYCOLaP/tK6XexyXDf/excs9Dx90+p5NyjId2G+zm7iBIvT/v+umqhVxJwwYK
fQmUE6kdgQp1O78xy8nbXI4on8Jo9do9a58sWZsQfxwFrA52zKGl11YQghOk3XRTXK1joUTdUvot
QBNhVUuPZCvDbsf8sUwotH+j0iZ+P2AQFGhFZYXmFP1O+2vMozpSkQhTBnwCt7aVSv2LcC4U3YD8
oxVgExc0hIKaXXRYvkq5dOUhiiieI4FmAp4BkYjd7/9qcFPoQWCeVqoNdrJjxFkLOZsnUuChIqsQ
frP1bnCbIZ21vPdxYPJlMWy320bjj6l2gmOmpWM5tpGmuvyYQitNyRKjiZI7F0AJQHZLzvHl1a6/
4KTWDPyFFYDlABqWKpSgZ6ccO+6p5gxjY2Q721qgiivbOlzVZD0FvjzS2GzhlT4I4tGKP1/YlytQ
FwiELkieaFIlW6x32lG/6RP1CupKAACp/2Pqkpx4WGZ4fFFEaCjCKIHLqbKy0Yxi15kkx6X4A8s4
IrWfSHYTvwrroemKPWwZq4mxYqgnd/7lfDmkx1VDYih7Wc48rh6mg5h4mrtJOiLSUDDqMyqMAQkI
3jZpMIXn0rtDPYz3BjFYcwPml77rBSti8B11U7+QDB90R77e2ls3A243NMxS3g5YnFhi5Rk22iKh
4Jn7bBwHQmUVdBbRlPuJmIksRCIM3waiPkKjpmVwW5EpzX0hgK+WqTsICWiHqXumAiTRDAlu8FGZ
aNXx/uO6WC8wv6mDHMVciAwX9h8Z1JR1/X2buKV2WBRuHR+nCLwFpWyIgE4ClYEoGCioSe4KhaY7
uCRyUA2qvss3AplzO0sYqnVQj04qFCSxiiHj7Eo0wWvzqrLXPZisuByx44Qoq0Kc6osbuLFICuu8
UuMDMtQTtzr3OJLFyBtuut/EwTwcYRsoUkVW9ODg42FN8WFYa9b+Wxes0tAzDFtZLtUxKDNjN8lM
xpoE75Zsc6Q7ZJuvaSnj+kTwkKEMyNQmWhuBLEsdN1jWUtB3QCXcAwLqqOf/diQByj7ZaO/n/Squ
gF7TTbagZBCELfz4G8msIk+eqtsItsKZG3Xi7luY+JPfYOFgJHQrUd2yb3ArHVdzfyM3xYRnyeGx
lQex0oq+vVp6WDysbxA1w+IufGjwYv+gkHLbeRS10B5ajpNgMErKllTpu9JV8hQW5t3jgCjTFmdb
/2N9tskuWvjMP9FGtASPnjCHjpFLjmR03/bN1hGdrw2T7sJGqec9jRL8TV4P00LLKY/DI0VFiARC
2tQCKjNgRNkDd22tPAy61aOgK2GzDrzVl94f8GXf2nXkz7uww7tpEK7BDkgl7JalpDDZAnp/sx7u
ZblDENMbag0xeJCfs8xh4IIHb37Ib7yYvWVRdvxW3e1yABYZ2MjtB5i6umjOL+0bwu54BtDtqaIf
dRtT75TDAKFns+Nhn57BKuzpziLEI7+Gpkt3rEWtnyLQJdVzC3v72z2z5BAYuAszUVMBh/x0Q0GM
GfBdKPB3sL/nJdVobnx8SRkzdqCwDGb89xwKhzGF9tH6nvFGzdDcfjRENLAU4z+hxLgznycICUIr
+oQYASjew4PFASHFm/CO0ZoSEoe/3fOiKYhOtfoZUrtriKBo77ot6QjSJfHzGZ8HMxqkMdhKqmia
sYKlXBEEUBAkNby1DiPijhF3F0skU7KD3vr1BIUny/vW06bRhIbTF29858WWXhPPaSO0208uFPiX
Rcwue8cp4IffWdXFsTFFOvXM2dogFqK7Z20dqYmrMe6nVRxVH1J4UBC7N0zQ14UhPoV4AWS8F3K5
kdqEWp4GJt3aCg2Ic+xmn/lPW41ApoiB9fjoV7ubp3BoSpFogleASQvSQyPeX4zEzyDLIQTHVr0B
jV5pwWYeUVqqAtYizg0YfqlMTSRJZs2r2psQCp/LhiMHj9jRsPkiz8jRhr9mHyycFdI2LsA1sJga
3FaUj3w3BFu53zmREF/UJJmaLkBa1CuwYuTPul3TqmTjzBsSq0siNbfym1PhIw9obiUQJIxYyBsy
fiQFZOi7Y5nzfZ1lqnaPVZtXGq8q7j/9NB68Uefo5gU9BqZxYqNyGM8qddt1EewpPqaWkZjr7zpi
yr85g4YaKu5oJSGRlbNE1LYmCRbCL9tnh4kUZCwfIifj2TJOkmsvhN2/FHQGoheNI5b/GVmX9/rB
aImJ32ghmspD7duAkdJ+QwCHb2O+iZX+gAjpco2A4GiwJv9h755wti7KkukwT0k861RLktYqZYvo
YtpByO0HmiJfGZDF0PU6laQj93zB9C6zWiwm1jYndTXyOV0UqSOA5FZYBhxrWuAEFdnAzu46tl7s
zQcc851MCb2+efChMr/+FCKL334D9OIFmThLdbRvjlRmPSeu3K6wTl8K78PksdjdYVzFdw2j+FnV
M7RhGxJvkSqV43XewfFV72eMqLzjabfGlxsgVaAz+YJqRnkFx5rEtmtzA8YmpJJNHdaAcu1WyAKb
KXpDHOXB/iyWWbka6lCRdjevGatY4Fe1V+dNwqM+qdmK1t3AfAHl0rKflrdqr+XC7UXWC+ZUU7Dl
VAnVsomj5/fdBkXh1OIfNiiP18vkXNWOgwzWzmph2xRBaDFIdta0dZfXSv6HGjDUheozaeSvhuqA
1aB5R/vgP0oie3Zqj6lhXk1h08b1Qgpvg8Pb/0SwKm2SzOYVqHXIqsLHh8X4OI05pgSSbsNIb9pF
lpsQmtFLAr4cL+XMihJFycx98gyFcmgCoq24ZJ1Xx2g9nSPvUResNrZF3gajPsGHn17uM4WalIq6
0EUfH+DmY8yWY5qAx4/Qb1Z0N8e2hd+KCV7XeMJWjbWNPwKvGZaeTilFEXp8GpGlBP8UrVLbfJS/
LDNmfZxvfP4AdkFi3gFE8ATVIF0MDf9tbb5ttPnpbBfUB37SXY6Dlsbx8M7Ith59Q2SPk8kjzEAw
5sK0EBMn56sYgGjAWn+UUTwrPUDupLhXwt1v0JiObEj0K/kFjnF+MY09mm7FPYCYfUBHjvotxxrI
2UnXuo4LaMyuEgy4Y3O97FIMPyqrBA4OtocS3+5vbDMNUZJve2QMsQV+y6wIH4m+RF4WqSbexxRs
EOhJF+IaJzZkxkx/UaXOAV0Z+kYQ/n4zN5VEdObOqd6MhnzMzvB0Nm6zt9gmEry2IWSKFyVgNIO8
PunKzdEM5yBeuMCq3PghUP+9YZ4Ct3RoP4cgLAuwxQ7050OLuKjoODGmAdYzAC9uhhe/VKssjRqx
3yNrj+BzxmmWeY5xQhz70fZ4gTOBCtMsCxcO0nnQht5M1LKk4e6GSBptslMfy3vO19dmolFT4wga
xVpVD6ArR1huIyMMIXKeDMZ58JrHvbvVF80Nmgj5dgOYGHA5I951dR7gE9nuuBWKja/ZUPRzFb8T
9v6CAvZa96xynHyesFuasBwsMaa7ezR9t+O/OtvoY38nZQdszB9ASArd4bY0s7FTNmfMsRjYRruc
V7v4uH86eh3grOIW1No720Z+n2RrL1BxaZgtIPD1+ZqFkj4h122kkskmF54dZ/uy2Uj9W2/KdcYv
AChH6A4GBE5PjeO3gxRezadFLvOSN9VHA3FqHzoMObggkQ/oFHS5MgT19z7fgd2+eAULym+u5p8o
DbDlD/pohEdJLVlkEbBwyn7W8o8hpR24vlG+7+6/H6kOxEsF3EFZJWt3wNYloDf+p2oVPp1cSpnl
n23TVRZ+lEBqB0al29g4+M+TaWACwUcK/77iIPurakQmvLeRY9YQB+3xvCavenyXHx2pIDFBG+mx
kZhiVZOWf1yOB8PnK1n74Bb6yc2+mfQDdAoQit1WXLgo9iZI+0sd4S9UGrIGM9AZ6HFKQNSvZDFi
miBmjApUuYH70uG1htroRQ2ADg69tAS81lJcDZk+6/Wn8oCKSoZcDZhxdqkf8v9bWxlQhGNMxMF0
znyI3G9uGuzqHmsnIUuHQje+PG9EdigdGsiHMCWP/AH4Ct2bcQXXrmmGglTWfHbQh4WyQA8JttiL
+nqCqnVwercKGadk3HneyUr4lX3jVedSeGcpvs9hHEOVAWlXoIdLYER/biQAai5nxF7HVtURg1Md
2OQz/SiUckPU339LVvf5pIx5kKjTXc5oWncVWH96LmtQkDQna0zkUCSjDMWbQhC1XCBL2t6RBEdJ
GJQltR+zZYVLnr/96Qw2Sbi/ecIZ8eTpYcoMT6ARPV27x0HzaD7Qin2D6vU2WGj+FISJHmfsBEwU
5+1e2Xwazrx+U9lxMmQVrmEj35I1vxKhm5RC23rlqCkxYEKAOhatjqjPaA8FSJ6gbRdg5S45BpJ/
XvLYNr7eglWzrdDa2FPLZGrKHVJYReSrROZWLO3zk65in5WzPhFOulT6RnOQrrMW+kCawIrm7ewk
yFyM2SGehJa3ktRBc8xpTub93jA9HK2wSO+6D3dUo63MmsmVODoXyl9f6EWNWEDfVWoMmqv77NFi
I2w7KhCKpi7H32TXhsFl9ST0R5e2b3mRCE6kfGI6jzUaoXO2yVZxpVMLzaJLI2fUH6Fd5Qy8zJcv
S64NVF7P83tNCJMxCnw6y9VCLEk5PocA6o5CmM+KdFUq1vylNrJ+me33KxOCo1oEtLi5Q9Rad1Pg
NEphCAh1RWjPsUVbnrQis2Q7TTlfguzrn8zFE2aMovgf02Nz7s2atAvzwd/ojic1ME8rzwFbe4V7
SXYv2qM7NHDETZPTp3s0e+PvuajCjnOkA78uZLtEsoANyOAQC1ck9blFjHPSma6LfI3sWmuYIURi
mHMwqx6SVW8gJWVcw8crWuGTfchAPic+I187AB9cQffnWbxnXzmNuvCIxTVWVp+wUqthRdRZV2Fa
S9Ih9FTOVDjT7/C2sVnsm7503X09JW+48wzBrDAcjtNdd9DBvoDV80oRc3ePcnqF9kXvoAOS1wS+
3XYw1ZbI9cmWzOraba9X/cNE0GqnoLP5tPMjY2u3z0CMKHnb8ODSzCfNF6eD52q9+OyqpaMTjlbm
TiqMKQ0kK/Bng3oxq5PFXbojqY6ZFvPKAC2CY4GArl9I2QMbSktpBBd6X7BGYJxGstVb2J3UxnI1
/sCe16ZgBhjfnHAO/iW705EQpSbYlx6BAGVr92yAdpZCgsmiYlCzVeQOx7+xWBdRXxwhcMhAOfIJ
Bq/KKbq2kC14zjOim+2czvPa4GH0PyVAoZqH70NB5vJQgGFOsUSWkEtEU6CerilMs5uYZ7qBn/Wv
KDsKpQwgyVskz4eqNJolFDjF5G9eC/7izzxES7iCO29qhCcpxA2c5EZVuaaRY6BD9BQ7RHA2fmxe
33Ry0ZQr+2tVnHKIDIDxnc6PiEJO25jdOTK795nKRrbti33lqPTiKQdIBv7yWazuUT3LnFIhA5Fg
qd+MoIrN2Na0AoJHYsWhKaDkJEvl46erkmlRM+rqSOcKnETHFlpdbpqZu6XF611c2Ib/k0vK2Ptn
rJ5Wp5WpJvehkmBYbuBSdyHHXk8KUvvLgodS27QJL87Hv++R3ElqyMZ2MkmBjpB6Qk8BLVvp2o57
oIkpFCjGBo5wZaagt80q9mugTaM4zX5A01px7kISE+15qxTjrp5yv+F5oAWmp6xYIw/XI7SGevmI
vRRmqqy9RTu3gzSmu8pjNTADd6Sj434YTqVldR568B4ykbadzMqHdQB0rCXk7Zw5b+BI3ZGoXdu0
uULCt0l00Y29CZus6DvJl8fYM8yVWyfnnJpWq3AlAWPk1prxCwWYkLOVcI4WAF5VbeafFKkbP36e
dd9c4K6irRegavBQbBUHLM93In9ADaM2xKFtFkgavVGOqWkPaY2LpIhaf/aK4EVPg9lSE/E9MaEO
r3Yv9QLQwFQxCiei9/KIf2Hmn/lgkjvsmySYfnMK0c64e0xfxNO1xn2Err8emZlPTVjlXWG/19Sa
KoDp6CkiI/JI3FEmt4y8agpov4i849GJpcdBOoY+Cx6iWJyoLisSWgNheQQa6V8SgVMsGGTPHf2I
R5D3GTLbybpdBD6QDuMqM0UFtpBeMlzMJboyqzVy2jHQqtS0XYCIVlpKb38f8G7UaCC7FiuSRNhO
0meXRChtYPp/4qs9NqdFL8DKqP3egghdYLqF1yEmHkWuaG+VqoOndORaHp07HdV6MOmNspHOwBsT
RhPhbH+dPLdD0aw7sRl2rK8pvMGX1Pn7UVpAzv1Snrdz1c9CvZzolgOCzvtbZdcurV/19r2uFWW+
+XtzGdGw3sE/PuAyGytQNdD8WnkXDEowfSYZFLTmhXgp0J02dLK0Nc34EwR9m3YcHqbQ+kMB2X4R
h62Vf1YacAQhsiiKB7poMY7v2YN/6avsyML4dgBUsHhPm5HF7KFUhTc2ndtfCjaV9tUFDz6KX58g
YcNYZURZxWrC1JD4sWKdj8LeIGxXupk0OsUjjosXFtHRO33TQoEdNM7qL2hERWPYpz3HIdEXQa+U
KCkUwSElIlW8oQtzJIYoNqP3r6850hzYqTW5JQbZxNxR90uqN4EDMR3Tjht9m8IfPKS/Hy3gjrkj
vSeKU3mUNfEhq6mB5SAKTQ3rI5JdkeCfArPvPBlLAAzxEUSTuPeALlw0eLSQowvwmsYxD/Mn3lXf
cq0PoGc2yHKzc3TNK1uY9U+S58ooWahkBjFzuVMR0m61JDjxH3E2ohNJpBXIQWbN+FT9u+oWvbk3
8b1m2e1Jygl0kgNjtVvsZyjvTj51bp7FbyDyIkog5Qy/r0cmckt3Qitxaosgds2BldxoOPNgJNmx
7nFtUQG/04y02kFNWq6Bv6Ezdx6lHw27WMI0XeqbC7nUtJye3sOIifA0ilp5TQA3B3mCjcy/ufpa
I45oLuUGEiatmOZsYpBjUqz2G/59xu8s2P8zRYMfoGhHMpbQOS53i6eEyJso4x+MAo2ku2O0FmWM
6B6yCLLcqcFkkpsOhn9vt4HMWe2bi7cYvyS6z8kNYKLCEH2TQcmJFYy4rf+lIw+lCsLNOZlY90kR
UKB3d7nmh0kGD553tUhQE1Cr8ac2dT1Ks6pXCXQW/PVY/eOvBNDqdwH01rSkzzGFi92IAKCGZ1RP
Skg0BNvnwVAJJAbrhvmp6h/5dJx8TCSU65eT6c/lSjx6/alzguMx46gwHy+aKs5nHBr+oSZ32yP3
iHrlWDFIWWM9LGZpbKQ6tRB5Ke/v/Pj3C6HfVsGKGU4nPbKrR7cK+3oU3RWQ53vCEs449Qt4o2mU
s9oAo1UYpS/7eiO4s8xW0E9FQqbyrlklwfDD1a4VRBHnQpKL/EmQZKZbhMksTy9xiun5MPir3MM3
Ez1Kewvo8E1eNVVvtzG0WJIWqNX2DlkhsoCU9jPQSKzI7sJozra5ZLUgRJb4h7+6ihCoihwkOpYC
oYET6TUNnoT8VsQHmvLNzUzZhSsf7PEW6h9cDpxI8vPQAT0ljVeVQtoSMxNJj+TFWmwbRlitM5Jr
E7JA994fpqQWks5Y7cgZ5aU1ExAdb9lUYORqjYrkQHUkOO8etAtRwPYqdV9jgk+883UWbokrxN+h
NOzydaturT8epVNkXakh47hOsbVvlxdIrosOMe1YAtdyrEf0hV45yKhNMBbNmTG+ZR+sFnHiaXgs
VnSvkK2tJF+75AzTyXLi2lz23I7+ZKem1LvdVJjYzW4qqOzYQcwktUQocLxppavZxlFiUxDf+f8Z
SeR7hhQghW3E8v1tBGF4jcMLRPTjFPOyZFmv8RgdDTf+5xRJMbN5RVCGNrISXUfpIS6iY+b6HVxJ
yTiyKMtD4XXPsQWYvpCOcqfvGSUGdGaKxUoDy8IWYE5BBHivujKpznX4CIScjKQR0uL7WQb9DKYT
sqQ8kUrmqYj26ljkc2itgJbUr7PCFgnR/0wOKnFJylCPI4gUMUL72SVQ4fvrOm7Bt/UTz8tSF7Y2
R7qkAfFuZ7aoVjg4Ad4gEx2bpY1uc3xp0OR16GFmBkzfCTYC061PcWrAJGfIgfIN/4vWb9BwnNRn
1XDhmbi+mSGmhLVsfem73XXn1O7t8SIfPtI1OO3rb2psPLgI3I7gXwrPuPHscCfSaN5hLqKQ05le
c0irVcH7MpMSiXRabB1NPMXvWGuuIA/Zl6naz/WpRnR/GsI0440ipl72rB2j0fsJSMs1NusSX/1z
/JQ4ERNnpVf+QFlGIz6bKobjDycst8By94WIN3zxWI6l5inF93U8ACzgVCqthMsjKTtFJI2yA6Kh
1gberewXLoeqR0VSRIWt8lOZ+T8NprHrUn6Ziqta4hf53CSfhKNhvrr2NxE0DjGMdyZ48hFK8lmd
iPZ5NS7JWV8dhhYWmrqqSijX7Kv1aX4foTt2UCFI7P+nxZyvYJhiefDaPl+VXPoYLtOxN0Q3g8OG
E+gC4J8NAs5diAOvPBO0HAETt/bE3DPvFdWZ7VAK4RW1VULi6AWL2ds8emRY/+o2hrJ7Ub3mjh+2
n/6d/QdEal/fABJ7f+TGbyieQOojK7U82XCHNIr5I6ZIS0/1t4N4JRLclTnonGxeJUqzr9MmRADP
OqRKdNDgyswZ7Y5ZYRmR4p+MmBEj0XTxfNnBXibdH8dVk6FLsm/KlYkZC9xarIknL5K77W+wOSo7
z43dJKToscow9VRJnRyXIA5PtJObqGOZOYehMYuTgJzgsVFadpOi5iVyNTBpOfIlT2dydrOYhwY0
4PHQ5eVV5LH9MKv7xfg+bRMAvLnoQYtMH2udl4YdhsxR4wfOEoEoUOTvIfeCVZc0+CFbpfF8um63
l54lZIoLcZRbmRFcluK+FK5StxyQraX9/W+lSfZtO7bKX4psD2qLAm2WjATPRdauZZTw6D/4D/ct
4bypv/rlPzUXyroC+ihBqbnAsVmbZDF6IN9daU1ocYpldw9DOaNQODysESomBExlL17V4570JnXb
VAuq1InxGzuBTn7xqwMY9tFhuuBloqYJmdZ7R6Z9cavsaxHJ6cGWc8sOLelcufBlJT5ysIO2J/mp
vFwbUwHfJl4QGCYcLf9EUsWPWED/QKbrfItz+gTqEoXRVTNjz+Mj9kzAnVh9emBzeM4YTeyRel6K
rYJ+wN3EddsDn5Ts7/oL3x5plHC+IS6RTXTPnUSk1/d3WsiC2+JrvGH8Kw+H9e2ew37JA8jvY2R6
UbwbXD6oH72Hmnw7kWKTI2bA5YtwaLpPitQI+F2w0A8/8CYwIVZH3rq1MdZHEm6b/CCsL3Ig4fef
F/op726m7mNcqCl43CkuR4kWgfq3Ifd4w5tGR6SuB1zV1L13lzAJJEZZmDsIFbzT4I5Sncsfj2bP
twaYUuWxSdhX30kRgYCdtTzcahR9aBjW6vP5w1lTkfa2d2c16wK+NXgjhEjpACMPp2Wrel2JC94Z
S+kaemRhzlQn4jFvdDhTuLBnPQHyMRfbnEyzbYc9rbOQXrCbNiwTok5BE8vju6x6pgPvaEQMkgK4
4J8s6uyj8tJ2YF20rW/1ZG0PzdRoKWzjO6kQTuuxoNx61QENjsuWJ64jlEKfQ60rIwWfy+IrBAgU
k7qUK8z4h1oiPSmXzU/RzBijD4iE7f0jzkMaG3FEZH8bfwtvac8pjtWw1bmMXMdx3E9tbvPMIi4I
gFp/NeQh7+gfxUdOggX/ndbhflcOTIuNN0WucYW2ah5lD4MiWBh1Mk02+t4sU6lHzbg8ti9+2lNA
3Lyx0EACYAumU0OXtViVtd59D3FQCGVhlDvfAUJnmwgjI7JKO/biSv/AX3KYpjbFC1ngtMld+oxK
Shjfivl+XjLMdxuMdy8sLFbaKR2cbG5GcO/RKq0JenbYdyfI2VqcgMDUjN7C0kNO3SvdtyJHEzoL
1NdttzG+rku/PAyVUmvn8MUjJO/61tJ9r99pWEZw8wz2nePvtg04htAjB5Y1d0FF7zEQFWK4YCXz
kzJ0kDCdaoK/4XEJowaYqigEbMywGMnwL1S0OuRzIUGmHIwk3lgF5mbAfibGD0DgqfCkNXhBkwoS
5nrwc3NEYFkba1No1/K8JxEgYzayWRxjt2XLQL16Djzv0NOm5cjQxcwVAB9rW9yqU9ByMsZCY6NT
gO0I/fMqU0jGNLqwXXlbxylM7IVtnjsgmUAaeLdh6YveDfSHVDJC+BuMF1C7eWtJ70KUmcjUgWqf
0AwOrySKHQWfdssoAf+IvD9jwrhgOzN6SAA9MLOQYBxoMlN/hrJCbT9pulr1zPij7cbeEYEAWi1P
fIWLB+Rixih21HqWX2CV/Ju/8X7433K1KffW62OxmhcXyR0rwoLDMx6Omw1RdWZzN3a8aVWskQL+
eXgj6LAtA1piIbm4ftexUX4O2dcwtZkje0Jy+ia9oA7ggc9+QGvCM4vfWvrf3MNbbduK4gBOuYQg
dTBwfq/TIRxkryDB1pkyZHouDySda3p+C0i3Tj9iw37SdM2O0hECUQJwO15g7nWTkMU4c02hu5AO
iA+a7YwVybnp7rXZntDdJ1d2g3G+SH/+Toia1u3wZlctUVaymtA9VsQFs3RhtpBUE51oRkyjVfH2
XdgtxzAuu6nOtqXzw4shCWZ5n0F4RqVipj0x+WjVPPeRd1kacm46QbKjU4fiTsGS77WZvVBnwBeG
ZZ4RV8bcUczX3KWhprJz8/CtbevOBrUL+O1UF8qdlQ/V/GfEYlEuZ3kQvixbKxnop2YmEzhdoC2x
xlTEHsxEv9TvybBz+7pcpDASz1lfduk21PNg5Q9KNwZpREbV5BJEFxJdendOtvTvxKYCTsg/0O1J
CWDcJaulHjSuCROfHBlut81wHgn7fbQraOhfUuX7EkWHp+6PrSosfXONpSVJsu26M8qGKob94VsP
hiPqIfCcXTZKTHoFo+APC4kalJYQyHjJraFAe2mWXsWkVs64Zyw1m5/BrzxbjBPHQby4YnJwBLUn
rBXOzl7+HJHPSggR4FtTlZoqAn2Ztin1itPhBVs97mClgDx05I7WJqONS5f8QbvJRZ52cEgNOwzh
wFr5MUXazzLfSW9uBwsNSp49UpWRMDbMW0QuDlEBq+IpaTpYv52CZ764LzyLinm54drnaKFNiFyx
IvAsbnb9yXKBUdAQ56HYltyY0m0LpXQ96wowsKZLrFRHT+xNTc0KLQzwprHArb1hsO75q4qfEHJ+
LBC3JMvPX0Fz+G7615kYUwT0IUH2jet0J9fKSLzBSUql/E90u8C5aMNZ/kHsUsxEBQgTYjtqK7ow
AeCDUiqQHPeUwWYVKaYbidj6YixBLFfQRMTGCQDloxglsY3CBULfPbJuYpjRV9LewpQwqOVA9Js1
1B5kpYbCW4gQblkmJMq1F/tieCH5bhKbp3qDpyHKouI9JkTEVbKAEDgY3+HcrjhQIc+u5v6v8Cm8
5VhhfK4IeazySLl4JZoQqV6pNsmKaOPATdcQ5M9dglBGzh9EygM2ybjOYzUIXvv8WYg+1NEXur3Q
MC90ZpOL7PYHyfjTH9rVRBaCdivKcfeYs7EKJUbC+E2dQw3Xfcf+5IidG5PM3kP4iBoYrmsaQHTR
yHhnwl22Fxh2lmi9X889v13K5LUyn47UxL02rFhQBf5jRw8XTi5H33e8sWSj/VFoTrSPEQqaQ2ma
KhborpXFZG8keB5Ipkm+/wYXW72ilJ686VDJEIIDhOYUKlHQJvCqde1E1U1CitEDHrIRuk8zbhbh
SfZg+DfYCPtMKYHIh6YRIKFHeeCMQyIMTxpqqAIdHWyUzPxMyca3BMe+ruR2C4KaKYnTH/iQaomn
Jg3RLrEaDVQtWTYKcKRj2Wo78zi6cCBYn3ITr6pSs/OjSxhodE5bxSxrZ8kyPkxgmH5kIsde4GMU
5xK0YXPzT+ga8hXs/vRA3MpVCE6eUwJWvSqlD1ZPnfFii8KDEZQxxC96YILv5hCqmYgy7UV2O6Ht
4Bqm8q2kxuGbl+sItUkSYK40/WJ2RfYkM1cvwj2sVU+dwHUEpLM5j1tMfbJXjpBXscrdefJl8eYI
q12dDBtEDnW16EyFg87G4Sdrrkaq3BDJR/Zy9dkPaVqlypend+TdlLZQSyHue3DOFVFt+ILVY7W0
GSYaH9o32LoXJUGXudeBmutF6BX8CEIBMOw9TODDW/rFCqh8BSZUF1X7ImlMqxZ4nYBFetjPAwnf
pY1ioaJg34hd+THmRnUwiqRGsAlLWGUffS6hnV8RxnIe0SWsFMsoN8bCpIa3w+IPvYjnpjOsRFfV
yLajtmqKNWdBXOxzph9M3VTsMKJxw5/0Gcx7YYzO6TsH6UikL7dcZ8PWtdVuRvdxqvFOAIKQDp1i
FvbF0xX6ZsgsxKQ0c2PhYvOM8gj2JwQ0RD1kEkKX9x3bG8yntBAOcJonttP5Ta9uLNkOnjRbFCUR
TTXYYCuL1WFMcLtLqIXRmRrSMfCRchcE/q3chILnoLgzq/crxOK3G/Ds6mWIQeFTyBWmI1+O3ntc
Ie972VV7sXvM5j0hM2YbgIDyaL62eztzVp3Mq+suLI1/K1+uSSGgi+lbt67S68h6X7lzUQvVd9xf
lyF+vOvrcB3U2qchKrOb+xctHg12eWMeeHJizcMIJI5oq3LkbezLevFw5tkUtbqeS6P0tY5e5i97
worNtyfxKYwNqok4PXuY4lkfhMjkbdBwjfx93sp5t3x4cL7NzsilQNdgt/2s5dUZjC+wS9i2VZza
rd6OdI6DlQ+/ITBPPFvX6EvWRp7igTTLhpHBpagz53mx5+qb/BTqnyiWfAls2AgVvvYgX9kkpu3G
OjwRMiGPyEZn+0qbI73C7npDVcn+FRW6ISMBwQa84Ks4ieCAFJu57st+CSU/awiFULqUpNywJn+C
EafuW1VCWDtzWxP7gWYM5pb2P7qmrxXy5BesMlQDnwN68wnBCX6HswiBjShZuIeCjQoI6b3e7qqW
TI9xc6FkVwewJo5AD4xl4t3U9R009KtkhkXuIQa/0rX8g9YjxE6GY00F9/Rdh6v6z1zgBHCWCwXY
rOTEeJ4mP3blb8veH32KpGGKNOEk91LUlOR3MRLJLt/CsqGiR1V+agU/VNijf/qjWYi3H1eNLWdC
M6SNxkbLNM3NYwsG3sSeob6X11pDLtxOoGB5PMpXejWOg/EN/fhwU2rvHZg/cHEG82XMyaK8dufX
2n/PHdGQs+hOgBg5MWEy++m4huWyEFbPtGgLLkzsertRbcChXIlpjiSIw0by7Vc6GCgZomOtuTSx
yUDthWGx+Do81gZm2Sh7MumsV5+um7WCMm/jy1TrL3xHKlIKf+kTFJExNwA6UwXW36opQ0T7/M9H
KWbdr+kupKf145G5kXI+8jum4NUBnVK0CXxS1iMZmmpy1G0FzcHFkTmDGG76JcG8PL25YgYxOIKF
+MaOpXHl4l2Ho4POxAoO20hurk8FSHySkmFztf8O2UAj/klanMmw/vqgwCfGVNCG19g+aTqXa18k
RVGyaI7VhAkBZ2Tpq7dc9BaapIkcAAlOIjmiMaEM2/p7tntvpPo+6tR11o6Wrsz+9CyV6BeaHo+H
LSB1+cE27d5TvcdTaqTDPHPy8zODYsLs4AJfVi44ml0sfClu0IDA8VP6AXct5mmECa7F316Ng+Bm
R5iLTg47iiGB/reIJ5ZRWkkvkjd88aSX4qfg3vRDJ89THwEFK/ecPu35RDe3iYMaO9VEh4WGcbkc
/s681Z3Dq6btD7rO9X1R2qgX5BYG7ZyIksabMRerL8toEjjv7ulCAm6MLp0SuYBch+mSoqJACGq7
lOuWC9ROPiiQYOEkWtHu6iT5dh9mP6d3zSeHFGDJc8ZAaaEHqIBWH6mHzFcNn5PToa/laMF5PNzQ
UITTq5OLGHTurW5bMWcIrQ9hG2HmZggoqVWXDY1dBzmttUen8DeApYEtK9xKLhNi0bhNDHqkeT27
O189ROkcYLj9c5wxLu8x8D+7WJkD56Hc+3eW00LPrehRlF9LshEeGGwe+gpivV4qIPkgEF0ALU11
ksHvrI0RhIOSB7swhTvfM9o6HLOsNzA3hBuI4sycDRpuPKZdR/A94a6+rM2Ds41vcN3OMi9DczmL
SJUm/7UI3YcZpxPk4BrK2xLJgg7PBtf7UFQSBBCnPXIjsvf8i1Y+BDBTo1rfR6KuL19b9AzRIrp4
JYV65Z4CZNGj4Z/NNKVSiuq7FSQzVV1h52NlqYLQK7RWBfxbwltp1g5RaEOnb9JepzmAnh5WyFGp
ARa+2wAXdQizrSshIDmMEhOKGnlW5HHZ3UgyXFwnif2PXH4SVMOfnpMwIcq0Hb6RoF9NP1JJYLmK
I8HBUYthGvPcHl0HIVUcv78ehYQvNjUgkGDHQqX5zgdEq78mdjFTL4RrSJcGCMBrvvma/5SdYdFz
kjF1QV4ZtgaYP1Q42xHG53UCoxSjRlypFHs52p+47cyN5o5qmxyx7iIEMz0ddTDpJYANAjwaLlgC
F1p6xeF3kj5aSvsx59Dbw3GnVM6hfCCIotIGpgf4KydhWF9UQjIKSjaKDe1cxja91g2g5BQtAUNH
ca0gxnMhUONP/ECYxBuT8zwW4BwrqaknTLv++J081NKEpgCGo64tXPpm6WhW6BHyvrmpDjyzVLi1
pOWQEfuQed/Ug4CUJWM9Xby/I69zV+mWdwgyQu8xYj8G3z4lRTp/QS+mzYaIdjCrgIGEFMJKTAHl
BOx490GcF3Bi47IZDfIKLE+UNLQiF/5f9ZK7/BLrC2QV0L1UXQx9frdbx0j67d0zuP8eo0NvO1ts
Jp1B4aY9oEgpZmdyysagELyVR/x/2MlPd1axx+G9rXp9NWHkGE5na/njfh1f3J+6Wpe3pNEWWWz3
IF83NjncN8x9rsNoDVu1Qkv5qjhFg94/1T1eSil7YIlKSrAmjkz1z9NKssJQHmToTDDsujxkp6V1
vUZ8FUoGEDLdW1/0WiWEyzvrwo6SwlXD7X4oAFE4pxWzSOAk6nn7ZtnQB/D74CPZMLYC7Oj85q12
lqowawoXPXYdJuvjP/pCIyfAOyi3WEZIiU76+/dE3z4pb3n4RAOH+KmsHk8hTB42tIlBWcp1QaZX
ExX5Cew/0cBIfBRTU1fBPhU/s6PVp2Dgv3GYuMXgQo5yR+FyLSQgwD51q8Fzd4Hv8bh6HVUG/Lio
9Q0YjMcKgNTUcjt6VIl+Eb7G0NFjzTW6xhcmmBoh/x+6YJWHHXNNuYUpCGwx7jVeddpxvded9n0e
mOV8kveY9ZgXvibD1qLf5toXCtEnwrc5Dp6dc1dLVC9Zh34FY7AeUF4jT+L0TaK/ZrdSvKnmWXsn
GzFkYiSKqQfkYiZKAHoieYi9C1nO29tTl8YIIRd83HdI46YFyXk3PdPzDFJH+p6cflBszunBXXYJ
P3vHyt3hfFPEMAhKLihZx4kcu+Htn+fhJvY8eTKZ6vFvqwiPZgRMyqTZG+mrMiDC58WlKTSMztwq
UUEOOP/THxNsXayj8wQWwwbibi9iAVx9HZgBL62NiKd/RL5cLJCKAYTkC9JzSWtYo/XbAHXxjUN+
9cjQF7TDRT+MCNtmL9BXqQZR4SOr+wyoa35EO0s7tIUj9lyLEPutUDTlRZYVBz7plA2ILoLfu2M7
IEcapLUiFbTSMPWl9M7uteHS80aik3OQ9g4ibQxRIUjR5Fu0/ZUf3YQJ07qkZATRva8KFtIa/7oH
Aw9cxUCaj3Bgkuliy3AebFRyIsp7ucAEiokv6CbDVsfjY87j6Q+h56IX1e7iXGRuwCsossGbeoNA
qbpyHbg/WK4pUZhl/NxHWYAt3WFybFCQkgsI9TbVm1/NEEooDuQOiGC9EIKqqHuNy7FfJuOkvsi1
Z/TputNZbQedhUO65sHICniFui4HK5bRYlfE8Err5gDOVhIPHJGjHeE6rwA2VMn3PnUICG673WJm
236zPj4nKHmtU1vQ7/a1bRlROQiflVEHTODibIsvy9RwmDN7fz1aILo8Q/z61aUdqDJOF+MEt4Kp
g9CDUrOKO27FmTqj0LWicp/s3Wk+CBppgR+eOmZh/CGRImT8dw7MaAPBsCHA0Ul7CjHQ13xyxR/x
JdGV7ECInlgnn32d3oiklJ6XccmoLAjg66yr3WAS6Oy/kUcD2zROETsFof/eyWqyL8B7ZeBwUJK6
CTDkgRczxsTtT+6BFMK5MII/g0J76a+dIddt3LSbj8xNO2TQa3YCsn5ILBGakX/LSXzuRrHiKZZ2
pAbQkCeGmCGAguCN0gb2ACru2Ctms1+szkYECNsE81c+XN3Qpm9KEHE/V0xBSlpP9pUQzHhWMyG5
oSvljtfpVCpL2pWKoQVr3NYCczZFZ4EarVsTdevY9hyESo2V5362RXccJOW5noZcs++gA89yFO2r
/PkcuKuWNcLMIiMeDv4WhmiUjJGiMT2UFOuNDQnEC4aCEJRQQfhgLLJGkv8P28Wn5L+iPEDSE0HL
IOwB2KozIv+hPVgdIM5DVo3uvpIUBkkw7GOGXz1VK9Go+pbrfpUnicrM8tRylwbWjAS9qpEnoGwZ
3JV7Do8K0AyaEFF+XwddGQK5yR9EU3HYQWBOTBa3L96rosZfwZUyVzKqpm9cOPQdKhH/UWIVx831
GuLxOuTn8eQ2YdiQ7Essama0xNuYhh5Qbk+nZA7Og8mZtZrP4ZQfMXuiiGS6FxzRoGn6SOFW6Sl0
YIR2bx3AJ+1CXOtuLJbYhv118t5tx9esGFU0qH8jL75CGJAMPsFidXDBX0cnk8RmAYuS6lBFr1U3
vr3Dwc8/mlkJIz5VarKhUOvkYfzfM/GLgKQ5EkdasyTqjnUsV9Xv2oHglkFnuWGU3APPZnmc0lZ/
7xbnKJg8A5V66cRJkvuFt/w60CXet5C3A1Vyz7PlIXKFxRJEXTYm3xr/5XNeoIE6BUMeLqyqTOzK
cURf+OhAotDjWIeRlcwF6sT85EjilrkZNXp1CoM0St6jlhFqSDgul6nTV9OZA2wvhfqkE9XBt2xe
dMizKR20rFkWZz/wB+7jS4CrO7eXSghRGKV2qZ/KoN/X7Dk2SqUjhipBFousScjWP9NAQWNpBWdW
16h1AB1alDNRVWGkJsPKPCBB/UfuJvDrhaCZMECaf4gOEk3Q5XCEZ3haPryJLSQFp+TsSwcW0w31
QaDebVgw9ydMolakMloqkvbODbrig56fPSAw8uI/0zBrKKfvUmUqRV8BufUU/ZS4xvdxAj5Go0op
1UPNah8qNDWzYvLxwVXPXG0XYvuEUfPxZy9Yb+e7ECvkkfmD89jbbn77tptJtQhc64H9LxXPI1Os
DLNKvq7OCySV2Ws8hq8VxHghEy/dicyz9kY2dVth6yihmQfBbZpvdAhhT0EHPvix9v6FXIus3EBU
6TCE3vDSZ3IJa2JidnkLFM6dQXDxX9Qcs3kJ2FgkOYUHBzAP1riW52E2noFCT1A+/bDda/vJu9MG
KkkVOG+69BObZmghJuK62cQlGKOhbiNhffwpLYmQVP4UGHtLGZraWA3UyqWj8IIsmre9dlapTANL
YLxOFpw9su6C00IJJoASXRbIgsUqCryLzsunxJEze6W47Ow6bzUT2h589BMex8aUOVCndb0/M3N/
dR24DA806OmOGW+hK2/8cH0s4wk6x6WwSTz5sVV3aBtfjW2yv0wTC8ENnQK2+8Ocpqpm4RTWX9tJ
i2boaVvl9byy0Ul8tw+qE4XKo0M3Isp4fA5aOW64Ax9Qp6U+BTzzxDpMm4HyMxnqgCf1YOdvO8s1
l9ZCR4ICsFwW/uGM9v7wtJ9IcKUy3eQpA5HnhA9+xC9j4kVPEC6MbZBJ7Y/RkqPseQ7g7lAJZyc7
sZ7oqxoL7VQQrGCK89KkroqT9kxIFzb0lbBKM1W4bBYTQ541C2dYHcvqvZMgyr6IdK7nJ2O4y+Ry
0fzv9Mh0qNzX5Z8Q4SlKtFSmmulJHFsVQx1CTz8CdPCiDQ1W0r7c6cDHPL0hlGOS7Tf+chfvJ4zr
CJaBpAdGEIzMOjujHYFFlWXOQN2wLVJhjHW7iUb2blZVcLx/tbPoyIwsZIxIDBhd1V3bKO0lwCfK
hf8tG5a+mdFMG+ml2K3WZ1r/QGf6M6L07kCq7X+9rEc5uMu7g/tqgkQLvBrbomki2jUwtDEZ9WuY
TubCqtIDqs1Lfldiff94mDBj8VEw8/LKPMcKCdffCr1ObkSaMIhlv7eq8HGclrRrpcS83qCfNTeF
xkNwo5bFKUIR9gNQxaeM0D7qIN/V0M3KcsLU46YkUZkzoZahSJLPlAmvMBSABOZv9Asad24Vtug+
+OxbTPSiHEKeF6F+0fCZObCItDOA+K3RIT1DouFqFMLG9dKKS9XvyW9tpltVG/vWTjD5PhbidsFI
BEEJ38hwrCHF814tPv8X7sz8iNOX/c8yDaxpJI2Y0fYeoXRd/MhzsYEPcrg2Y04Zi3ELn61RmQV7
URKZNo9Vc80MQFh3beYR7HJ5n0GOWFb7mn+x6cVMGDadFP2AO7/UfusWQYWLEFdIou1m2y0g+hKj
wfG4dv0ICA0apzCs5G925Ut1s1/jzb0rWeI/p7YkgkLRAYSpK7nAAENq/axYXRDBIpk1S+UIEt+B
HY5m3e3iyW3Rf7YorDNYU9dts5xCk94NCTaHVFRERfJCrWAeDiW7PwqZSzawk1A5s7MQBYzEHIVK
alNwn1UCLlZg4twFvB94O3NKwYvKUiSWKvxpcyubrbpHQENrPlOY8gMH//alICLxFH/dhUdG86MK
V2aKE9DsgSZYlZBb7q3ej0fx4rpH+hHEYzQrMy/VsAB9oSVS76iru4+LB7r0l1/D8Ay50VNYmzUw
ORV1ebylsF04ymGyN4JXR/AHAdSJpOWiS55PY70FTJw2hC5GEg3E9IDZPkBvWFGYLh7sWEKz5ARW
U70FkCMoGbn4u//uVkq8wjTo/ci4gXKAuawXY7TUyajyHCCKyezM4SsS+RAthqNBcHP+PTq3ftA1
/dwoYz/3S+OjVfsczEI+XaWEa6FmcG0nUIFo+8MNQyp5HycC2jbKMQf2LFPixsHlJOx9ODB42MxR
bKCcYlsTCGX7lrAqHKiXZpHw6Bm2pEh0hmRI/ZQYclLwa6OKHL98jmFOzN8Bg4y2mH2CBGFxaoU7
ncbh7ZZgKq+rc8xb7GqwoupcKtVAceE0n1Ke8Hz86obSg8iAsVUtjotI3itI20Ellub768TNeJug
JS+vzKxgsVNniGn+eGB+WNxHY73b/HIXVzneG4Ny/Ipr3jrv3DG9EZrEjw+qbQuWZComRv3I880H
U2X7ILIn4Y6tjZHttVUk1N/Cr39N55ZMW8dPvCdL60hrkI2aGYgu/f98+8fZv+oT1OQHxHL1dO9j
Zr3Me9WJzIsfSm/+65PNJSQr3XIwwlYLY7GGAOY5H/7DxDOjDfCmXfFrkkMJJVWTWXL1cHjbW14v
l4HkDF/ZzHuHVBUDaQdXsqaXnlcA28cARz3p31xw8EM6qBrBl3CoZFB9uCHuQWg93BJcvBgVfYeI
4ZhCqKtlXw9Ck74vXyuvk1gZkIa6P033gwHVK8Ytq9v9boDGexvWl5Y7mXunP384KnTu9geK5Nlw
8HI4OggL/P3/GLvK4kvgnW3CGsm5cSSkgrOqpVFXmQWk6DbqlPTS/7Z/ZrD5pZad33vK4d2PzTeO
uOpiTJmXS6t84T6vTnIgoH5PvBvjA3mS04TXBBop9/CpJa2+WWbaMl2skmSrL8BRSXNHa4SWJvv/
yD2HL/i8DRzRE4Jlfrhuht5qOMuKJbLkpYjmcTqz91QUWWzfXdj/Z3I34u0jDp2apGjhLBuK4qdq
TqbUUle2aW2pv6fH0uo05+kEuB8ipeqhZbECwtJgYoKDyRscKW6HNCdrHAQSFVY/kpPio9u9Fru3
8q3ThK/wgdON7Xv6iXus2mAERkJG3FygPPOTx05L+YpkrDo9l7Fz1en0BMYtkbAxzzwIZYmRIhEg
l8nQzTvi3meM4mqc73qtHAlaze4fg4qT6vOCSY631N2ASdQ7CvDUP4WuzlwiMEPEkeQquaZTD7O/
aUodpmXhN9qNhWPiFLFy4AhcNBVhPk811wqRS4B7z+6VUzF78WEcrtu54ropJlxW8IKIQUDfYgE/
Ra1k1BMu9J6fkYmdGC96OPMm6NKAbB27HBkv1ziIkgguWESUlQjjk0ZSBDP5J+MpaFSniIrQSoev
3auBCkn3cr6C9CQGat447YON2j0QOOjaUWrmTz6xjzO3WbNynWI/Gl07Aq9bnkIJONT2SS8oEZny
6oX5GnZaiSQik7RhgFtyxbYa9DnTkBGeC0Op7n09WwrDwr9hqL9d5M6KbReqmYy+WVE2L01xY/7M
Z3IuhPvSqN0pkmVfDj23ldVGLmaimTKJdu6p/XP+ZGeyKYHOTlK8/Lo5WkS7rsOwHKWcceZuCWyQ
M4hMctRmEJOxP5zBk6u2XL++lsW35mE95gT6QGirTpIJo+htFR3+pFa7UM3Iy3ZSguHLvBTAMwL9
NK4cF1vgxO4CjWsSZFw4mfsd80Kut1NaYExZzvcY+BZgShL4XN8B1qg7M1Ra8BUbJ9u9LRXw9A5e
zivGcuBTk93Hw5auhCLAHK/3S5btDbxMj5qO+vhl1jombtpXOOPBJXjwg1q+yOgLwOSOVyiPs+jM
SpaNeBlBv4N7/TA4nNWkneHt/wZq9Dta+c7aC/tgQzIakxsVjh3TYo893NDzwFmF3S00vHOLrUjh
57TdYNexYESjrF+PXRvYVk+akw//I4wfU1EFTCU+FvG4XDt+18yDGXBL4eL5pA63FaLqsKKgE0V7
/feyxZNrhVlxrA0TBmg6kGbr6wbJxB275BguNCI2QaXCzXqNntH8xJeRCcC6vV6wAaYOYCU87beL
ZlF8Qb1CS8kzMSaRQDFF2BmXfbubix+enw4vV+k6ZnbruH/tagdWDp7e3qmdaeV09koFGV29iabx
cHU+7Z8JFFdbz/T5eTAWKFzLk6OT7uQqGHM1TbuRivC3hd2Yd9Iq0C2ifwWS3A5PmxgFx8X6QSci
qvkr+jvzwJhWFIVagNEctGWWB5TbYOsvF/JosAEyK+eyVaIIkXNWAuvgyq2zN/K7HKTfv/CZxNY6
E97KoqL/7VGAnDTzNr5yCxdGAiLSUSY5y9ERVDEJYymh+z2BFl5A7yanZ5hQaPqHHTH0UPydvQgE
/d8OjneGvRsn9i4p5191WzbOVOpjYqKZS1y3jiy/zcfC02Wk7kVXOe31Nor6yz87FYG0ykAn5Ta1
Em8tjj2TnHWbyUfPARJM/n4Mm4ApyXYVRxiEN9D4kkdFiWO0sunM808GBEk3qJD+9vP5U4WiOzeF
O6BUK9OCxNPXQw1NJcTxccvUPjAeD74LWsf0GOcAT0dSHEYa30ucRJOYBJYomKPxVR9rkVcy/XIo
KrCAH9rfx2CIEFKzp/hbM/8s+xP1KiI/huEPEdZ3VyiafG/X+hgzwo9skv18qX+M1Q0gSduZWyZY
70hvXTJllxFZb7FcmdyS9tB2b0RobcgrdHKV/hYEqfbGw7G19juq29zSGrYo1TrFEU5udgit+ULd
bHahYET/eKc6uCC1LXnV5OITwqJEgI7/kLaMhIj7I17Fb9d3Sg/T588+x/ZwqCAW7lVaFbB08hDz
FjAnxNVRUZN0HZYmdirp6S2EU7g8itzEbXZrSnXvTn3zIDmt1UJR83FNAEbmjcA6Im9jZuKXyRbV
RDTyKp6PlMUxoRL+DiDY7BTiC0jLxv3aCcMPcrBHkSIMuRTDA7/VumHIvPyjY3po46F8QrVqF8bB
ETuH/e+EFzq9ugOoqySX/X6Nrad72nCR6ldZe79Gq+NV1ONCuaRVEy39708MssupDFx1g/7ZxyMj
3JafEaCm3I220dIpunwRtemtJdLPKlbW4O+1HWudGVV0TSc099PKel/dSt8rk9fXMECKdXBmBNtw
TlqOeXOyRGjvOONOI9mpgjtEhMxkkysedQcD9VMy9HUG5nFm0QI5yUtGn9oXfuo+BnTS3u0u8rO2
AuqxlRqGePyQxtugdrVxFKySUzMUVhf5gpOJOyfz1zgCXaRrocGPQdZSaF2ahYPVlGvUZo0ScT+3
l9bdIMIyrGuC7TsJhR0I5uoKZiY+7MbhLjDbx+u7x/8jCKXcJgzTJRNTLdlva6rlcRI0dMey+AXb
Df0tUmn7PPWUlsS4MxNfP2rp3dhpUXVre0q6ULyB2qKpgRXkWoBw6SsMNDGv4hnSwZzCj/Up77c/
dIAfAR7Jfg0I8bEiYi14WGqYZ8DyvQznOHpUaVubmGcR+6V8iuTWdif3KLfZvO3rQqqk1jiu8sJz
A5er+1S92x6a68vXIvnaQx8sGJbrfz6ik2A6G9EGeKuTMfUrg7S3RDcfxw3LaMviOXggkXNwSqgi
AG0XZ9sfMikD2EutyHuqnTU94VFnHobZmN4C04ZjzR+WYASSTxZ04bjbc9GSV2APPisM114Ef/Zl
3UNX5w7vJxRcR3K4jO6ysaqckzirorjdDcmoYGA5BdBNhKufoev8JOOsOuxcVESCRaCakBf3RH6H
Rv2HXZ5EypdGh2uEI54RMqb4AA+RMVqqBDx7ATBlYxB7SqZ3aYt4YmE65lYfMGOABS0AEIeREIlN
XW8RXVg6Lapir2olEGXPLptD25pAV58jbDVmaE82wlK143oEfNrJ8gXDief+QXfhnb+LsluSdCID
qc1dlSS2bOWyAQX2RmXrR9wYKwk8FP/uRD2J3fW59UvMqZG72YchIidkCYYz6rZRJC6xr0NSPtJc
9laf16mYL3mcp+b9CbHCN1xIU3hsGduNoy+ar6lotRUeqTNxcDkyh4FCMsWTCZSq7aOpdpR/a722
6WT49dYshIGMCQLZmGJFDJtq3mRstsqWrwRpJY0yl8aeA8DUAcv30km7rRsBiTZNHvB06UeVIDKj
5LKQL5CTEkQ4nz9AOX+K6fUa3cHA+LJGigNWxIaXVqLD/3tr/sXdTbYrQI/1+BQy/53LuV6rsAk3
7828hepDqPBragwmaJOOOGqse0809OBI4NoDNGLLbF0t7oRs2frMzLC1oQwUAtrJJgtXl4dBpW4t
BWmeIOZvQm7rba2/znJqRyJuS/WqDJ4uqTyWEjjbyB42WLCQHesfwErfeNCN9ebl1/UWa75K9zS+
+gtAJvz/Cd/svnM9r+xd4UAlqrCtkHVkQmy7mBAOc2mS1WguvbrIdDgEHR6qSzYk55AbVFCDaX3B
PEhaBkNTrjvAtGlI/udfEWDevTYYLx9KReJjzV3bVm2wO/8lGhrTo0NKzjgmKxUmfTMSjab3rUAG
/isCPHLymfn2J9+WpkH8OkJp4Jeiep1d/9TfdY+yXn0pv0i8ai07/KcfPlfrU/6ofynlAD8kQogL
xg8YgSl1jk+sg4xWSnTkFRCLL+Us8PLSrnKc0XM0Tg0oKrAjTn7/DlyFPbn1Xo59mpIBLtNwdz7J
zLdZEV9PESBRvzBhuK0OgxuVT4UBEDWEOQMVvDKhPAan1V7ZpXogJLdxBY9zUaaa+EpjPlbent9R
zluVIXMOz5nAr3JT5qwZurQu1ru9i42MZ8yTJssta+f3ZeKdoYDrPvcasYgoQvAGxpkn9FuoC+Bi
zvL6fKcwqD8Ed499TG5MjtHFeghudjXKxkUjD8drL0Yuqns7AIjKtCVhxiIkfYXHsmu+MzGfZnro
JU9WAsS8E5zrjdup5Z/VLZcWZuDAScG2eBc7eI3wUeVJkos8CXlCA7bqA93Lz2bz1+Xoa/2Ep7x3
/pfYjlwsmArtLhN8Dz2euz1ubzYhv3T3adsKy3Rx16n1nGxzu2z6hjshqXyJyxjXeFOzWyDm6E+h
eYmYwYSRFIt8YVGNbje5YGWVRiQV3w6AejWe3CnrLM8wGuP7zS2bwkUGyrydVGFwMcLIhyhL6d3u
6sUgvAu148oBOCiAG69mtt4rswIf0pQG6cMI4+LUyIemAXqTVX2Kqgsb0Hi/Vu4eCHHuDL2qjMvZ
D8uc2dXC/LLMNY5FGn7ie6VqXOvpaJ0g/BNEp3+2BQ5MKlUtqk460hGuRyv64THHl0W/2vfqadZU
yogWmnXx25/kV0Urgmfpoi8zfAY/tijFMsc0FLrTyQGT6l6C5B9HbK4ipH6hxIn3QKMOIc3ec/EX
0jmuhk6mHVGZWA3IjYqf8yI4LbSySaFKwsRne7rbLpxqzuFy5aGU8Qq8If3/z/ztQWbchuG1FgpM
N7wMve2lKiOaDhKCThaFumv1tlk9XGYD3mqmC3sF8t+LVVabFcJRoQti9k2/9kuo0c7hlM9u1IyV
GyS1FzxZZXXABWRJxeGa873+aXhAuSI1LbO8AsyOWPV9Kp7dhgx26xeLIvF13lFjHgGTgVFl/E9Q
u8tWhdwoXM9WWjEbm5pj6Y3F1scXThb+MRP5Ny36ZDOTTANvMB3FU+CryjqDen3GvXVbYUlP19eX
YBz0bmWayIh1kNjTS44a4ycZBwIi8o20loG5YD5F8k4w5M7J8y0yQiP41k99Nb0NLVEqWeaYP2tF
W99FH7N4+zkQBXMQ3EVTyq8uzu+1XJVdxkQ2WFGkwdCPXWF52+3bCRVcBHE/KwqD6dWzqmw+7t9n
83hu0znBqS5pfZmmS/CnoZZAdSwEm5elUuW3u6vZ3irKB07yjmWsk34Z/GKY4NiI8A6XsWA/DnMT
tgX38kfWDiGj3g7Vx3ARt/S14x4jixIKxOHXAN+EChnLAHqpADjBFEV9lTOk55cYWDJGj8wOuzO0
1MHRZZdY1SvWC+o5124E0wviheQ59nFBOErigzIw5mPW3rDne553L0njcMviixyCRhA6lKTdbrOW
OqzKgncgy9WJK+fNHA/tv6Onp44jIBMQfahL4CWn8FoOe7Rw4I8HoPXV5n+iat+8rkKHdNOzSad4
0rY/Y3BcZW8qnlyZ3KLxiOGlnMzKg1ewTdWIvaboWBt0pXBLYdriKoYOPM702eC5CviTtnV/8zDu
TApw1rmRJUNBN4pMzg28dTDSic+TRqRJ6FfFisWDIGIFUoYirpTMoOm2sWewT27X8Lunt3FVAifu
0moVnGS26LsHLmhwgBbEYyNFZGVwa2DYMeAWGz5k+2VgILlsGRjiHvfPZHb0ipJT4tWGqHDoMYpQ
0aBfkNIIWBLS1aSQlj2TE+tcnlqKRPKO7HZYU2oh59KE1H9sunk5XdXruwBWPFTUG1aXD7zxbBUh
Tzp2ZUANmC3cxCpV8w+tsgJT32/0OgPgx5XYvvqLP5fTePvwF6u9ntGLPY7rWxydkAQC8975P0rw
Qu0AMtJe240/SP4RRJ5LBChHMjhRF3xB4EoOFztNMjLFXogI3fKlV5y85R1oc7uquklDZNIiDXnI
3NbMElcmq4o2UuMDCTv5k8QgtV39L96xzUAd+tnmNzE71tjY7A3+2Ht/ku/ji0DtckzdbIncolpp
eeQ/X32+1D1mDyzdIFJrxb6Pc5iVlvjtcP5EF0m+8gRXh9nDQq3hT+XC5czsJHBQXyt04PcwhE2X
+8NLqjr6NmKbRGmC1sarYr4Y864ix0en79w+qixDPE4kpVL3KYeEbK5s2h7QlhenTBHVw3c83I0G
ox0vKCh+juS8qLkBBWZrWdMM2bGRXs6XjA7Tys7rdzGYDjgFopDH+7HYkECT1mSKEIgg8TH0hOrr
nTa1BRj/4qtKieCS8hDDBTriWlfX51+1ns3BMxYQJs6Eu3e43FzbJAJwdtWcYaf1FMpzlvBVCapO
xU541Vet92bqJxLdjNaDWX/Oo7HJfsJcIJhThf//s8tKcHnFSHwDGEp55t0+oPB6vt6VXmNMumFA
1vuR2ZdlUkEwz+KstxclCykQ8QgtWzLx9D2LUBOCD3+TjYS6ezTSxBJxWbUjJXkdGXQRPmh99bzf
5BV2YLQtRBuC5vDZvGMBYC2cVgrV0ACwrJRv8MZn64Za8h+5ZI+ofTytQt0zmXIYtNvDK7SVrweZ
qA3+6HkFR3eTXqlBWn5LREaaz4vdY98AcsllxH0pBPXi8AfbBP/fpojBlIzcc5VyRS0y1D0bHf6J
JZPvetjIdghhHCZV6RQ/rp2Wy1bRlvN2IJuPy/odGXYSXdlE1tnIkg6lMHJnOTMGCb8Bgjrcs/9i
H3IPq15EGmMVHUaOAvWOtE7AqgAEd7WFxEbybA3UCSszPOUYCpsnu43k/WdjmL1P/t/KPYYibGFz
VNl7y5YWNt3gsn0pg+aH7S3jD5LoJUrxaCJtGEq3+rKwGdsswoShqDivfpCjKPD5Y+PfTfnfnBfj
KWJm7E7LN7HYAcJZHYbncnpHIKPC91EnxWHfVr6WxxJJB3XDTf3lmlWlTKYGkSffdmf09zNphw3T
iDRFdsiayPL+7BkFQ849HYsYkE18gmLpJV4Q5yGa8gSnlUZQi1I/XtezIdLmZId/qkZdA6/fMyRI
JC1xbyZuPPtgg15srmGqctm31kluPRij7SVxHlbkEBLRkQW+AxoHUzJNLZak8HJPnxdu6r4FzvAj
BqEfDzkJl3nkxaM85grIXgoNmTgnuhiosdbZgK7x3jw3KX8vUbe97C3L7Rf2aI1/fuX7Ba6rKmbg
pLepxI45hGSdc5pftlrbAGOe0yFRbIyQHzaOCcm6oMk3IEUNILpxl3MgnsNVqqpb+/CfZikUuwYM
W6k2FFGKyGZZMEfTevct6DLOoL9yJQm+fWC25T73YYbWzL1Xhg+BfTYmP+dlBfKEXktnImH8he/9
d2GD4/YryEQKmLJyS5Fp/H0mlosVUEdB2wUxIh/qnsVw4fVN7aCfygXsxNpE31hWaHg9BaY3TXYg
I5H1B4U04qL1x3m0FtD0PFyGeIXoJp74RYAbZ1hOO0OLOMJAFMEFM6gHf0u9MFjGDC2WzRehEjKU
fTnaUt6J0D1xEUTTTG28GMekH98CqEN5s6acm8U+Fn6mzjZspKlGvn7RCAoin7QAAxyTuzFtFarQ
xFnzAeIJlCbx2C7dTOja+jKZ6Xrio4LgaAJacaFKO+imIiN+fNEdlt/MS3E7PGKq5CxlupFkwdEZ
AeQqdH/zxZw2V9qYuCKucJxXbBsIkXnkd6OSt34t3py76pFwqUSY5Hs2TYby3O/V2QaSwZzpnzNq
xDvSojkpHuChJ/ytPGAeesFQ6y7Rg+tIKUQqE1Ba4rdHjLWdxUldb9NGTEBA2DOJQgf4+F2MpcLN
8WBfGGubGafESjOp3uaZz5iXdHk7kMS4+YU8SSbH+nyA8HHcyTi+OOuRA5GGY5kcR0KgPNvyD81k
v14cPY4U8bsu0U5Aks3vaQFdJAG2tKG4iGEXYMEG6AK6roJmTErKM0gEqGV+dKxQalI8qFl9rOTZ
6wzxCReeXTg8QbMnge6cu67BsJjToFidgrg2ESFBgh7b/vfCpi0fuJP6IzWFYqQMp09OiMz7YOy6
QfM2G7foKEY9vKwsu4oOkRqEkfKci6G2O67OOWWYEUjIJiTEzLoZmzzopVRUtLMG99Z5AHyx3ER4
gYOgJ7Ev9Q85pRLZmTQFf25twCce8w6ftp90uiwGlVARWAhUMiTdWv4kY3EG1xDe9/Ko2vcVenkV
jc5UXIO2ipUyDI3puwEzbeXkCsE48mTFAQq19biLgGmEaiVScLVq770OoKzUmDwf75hsc/n97cjc
OGq55a/jh9B+WcfYmevJQyJ9sp8BLZz6h7G7kYIu+V2XZRHs5w1TYPKcxyVz2LSDyoqBALAUjyCm
1EXsLusyIYdG1KKGQ4yqER5taDtjDwSUba7SzRYGepXXWT0t73uROZ+nbGLuCBfYCGGHwmT2gCXC
3AM6T8XnYR8h6afQNkFdPw8Qwl3Y3zJryhJ+yTsNTyoxL34y+NJyoZWutvOsw6UyIGkrCaIP48Jy
ahJQSal0mth/7Ndk/RlwgOyc6MeZso/b8GxyH6ZE69bV6EG8WI/6cKpjP1k1QduN14ZbvAOQz0HM
wb3OkGWnP6hnFh/pswYtx7MbqCeRUX8ykLekbT4uAKRO2ZdfmBlb5aVtRpUQBbpHLxtPMVauoBWK
BA5IV1aiwrY4+18N1hxOvOCcG71tg+TnUjGCBTbSVUc6pYiHYJ/mnEffvLOD3QPMbWBxGMm3EiTi
0WBrEOT3QkIUFsPu1C04grnhr7YifcP18tC+YsXTR8P7loMW1W+WtdNVGCYIIloTFDfHK1B6oTEi
QvnJ2qbXmkhSM6564N6cxpZ/ElZb7f4RD75E7iSKrLeHtknfzRky/edy4nTNu5SdpA+hBuGE6QAY
LZNCUuCuRx7xs3vaPhf4J/5LUOyqqqKdjzn2liK20IYL5/+fdLaE6JRp0mirWd8F18Bp0wzIM+10
w06FJKiDrId799KipDGwztSS9IL7oa9Isyedw32VSOk+8BIAq76RWp5P6yJeeKzOdCdQ69nw6y7V
MZoZSLWUXT4X1hbjlE8voK8XAkyDNjKQ7tEVaAFULpyyOu8UcuT+8Flj+vhKHUX2rvLxnqSMXW7H
VdAKmLxrRIHIEUeK/x30xdwnWbDQu1EZ0YB8vYPX6/QLWuG9llzAjre9wmuiwn4FZgw/8tqtdWCf
jUCUKSSOYazsVj2JQRVMawTgDSOVl0bGbwP6RyKowK8FfjJhGUeZyTvsfySPMtjvlT7E38dpZ408
SrxDAQ8MOfDUKzNT/wfLqXboHloU6ar90nmBD+M1lyV3Kq2UItW54wnOkIJO0OG+kahD3rCp0QqV
ttT1KCWFrSwiliOuyGKRs5CAwXpuT7VZD/2ScRVuqRoh6E/K66LyQvL1KRgyFIVga9dhw7LKjUw5
MH0fuAoDFmlhs0Z9EJxUQuScLpfY2GXSII0rMbSYCDrNLP+uHZAW1tllwu7U7+b1SEN9ytisjxFt
NJN2EItMr+79VCupCdkgI+Lxw5nVOY/52aarjdc9CPAxqrXnBKjkwlk/PqA441/0CG7Eah0neMEG
Ui1Q+h6VfpjHr7ngfR9/kHvNRCDD/J6+iNXFGYdUufg2/OUBCVYxLO1dxkkw7FKoC1tXCKM2dycE
qUZaxZMIt8gcK/qqS1tHoDtQbSErHEDL4CehJ435FiqG0tjbJij1wiX6AO3LXAZjyS/4s47g063F
3WAnpi3nJZdDsccqvmK1dQHoF/xNmtMBPXKIbcij6bXckMa/G/Im/VoeTuqTrh09SB9+lta15Tvf
i7AQMiSkK/93HwZVQAzjWjTYLZJ8NwYnJO+zq5F/VOhuoTIaykmeLQJ8iih4GNwouBmywH4Rqwsb
XFxYV8Yo3kXcUi4wstqHkFtxa1TbkEfjOxjktYIrVq0XNPK0UbNZZ9wv17Gr+xEFJ2MDUIOZ/dM5
jsVaOfeg4G1YmMWFIf1Or1cq0+3UHAKhNXR4Sungpf6ybPoregxNSn8gd0EIjDyxB4J4RFNn5dhk
aLJlHDLAnmDO70extzN+a4BWY9ey7lJLTNBl6VfOQbRffSgpZEEVpFztipKngfGW5qAK/9mS/dbE
/Lki7blF1qCCAt7Hv9/DBKcT5G0S8mTpDe/SYP/N2lMO6/ZyBXAat3Meg4CGnmj7ED4IZXJnWb7h
mjY9+0nflByS3QLeFKuI1P6jK+DWX8jJgMsKCzLZs1PUzEtbDHqsSuo52tppcJ0METlno5SOr7he
fNtyadpYdqacANHsvJD0Rqu7hQTPMO1M1SZ9XZlWonPXUB2ieMnjY547KUDRrjqGsYZXpnjCyst7
QMwcuOl5dQDJrMQCXp9+AvanPA6/Uq76NpjCWtCnX/Lrw/Qzktxnouj5YpeYzWCMmUd4OE1YnJNr
vyeFV43lBzouo4euWkNZOck4A07GyOcY3f4L8Pmkp0ioi7dOMseLStMdU2RgPDbrWkbjN4J59/vh
26fR47YyoypCKznIF2Pw7EgltkBbbX9KIfZXz3dmDxGQeHsLsxdK4P9SGfm4pNhScS4Y0ImY220R
hCAKoL4b4iefuC+n1mgwz1AUHSdAV2cqhTzsD+lW3hyy8nT6k8IHA4h5VKG0ukCln1WsYnbp9dYZ
RbTCveUkQHuW6raxhBvXCu03SX7ALk7bmO8hPjd0V+wcBJUJ9tqj+3dEHMw5z1a5SWK+SxCgCgSm
FGza3/RqLFPzG3Ct5MTaGyOHq5QO5MFde0NjG7WihyR3oh2GVvmMt1Dx7g5Mx/e53GjGgEl3zPVB
PUgXYe5/kzM9codWek49wVANzWuUxiB+gIT6UvIxu0I+ivDYg+vJiSkq2pkP1bCMpOVdCxVm+MEM
GIbr4jwQrQc29StncpNeqiYxnLgijykM9q6ClxPNsZTQZSb+KBN/MsTXp6d0UTtJxn7N3TseLj7z
omQn4orswy/eEuLyFo9KLzpQwOe5LNZZj662snYjffCTbc/PN39iiQf4HtJbXtRi+UBwSxqUP+7F
+j3VjGA+Y//dlnzN8O8TeQsYG3P0Sfom1kA1eeODhxwaJhHVQcgL7ps8PEEotNtaByZLDf3RhKlM
yZ3WyB66uDiSDuy2vmsG1qJQn5QxQzDji7Ay2QNt4gMDwZWzwExE04PV5TbuL05kM+Lg5NDiC/DM
rCsQObzjof6SEnl13hfIOaMZvmviAEyTGXZi6VAI5nNUhmjGD++hk4ndBii+/0ZqpclLZzEcMVld
IN8b1dAX56cOEmsjHJUtIWa1vpDkROx3iFEepZL7pkgUA45l9Y7IE/KGhut2BKbeYw7/iJDmJ7dN
+Ium3fS14jcK08t3anrA0pdnsZSMX7NFpjqR9Lq3yMonEiRhN2h4/yAhFu9WoqmaEhwaLr9lPQSM
o0L1UQ1qbcOFApwkdIc2lU8NeF12OxTlJUFay7v5TSsJh+jAES3xqcIHNOV+KQpZ+ekpvVx3W5aK
/GIauNJYHsJBssaS1yq1KzfgAKbTQMStKXXCfq7V0smqNtflvBG+5rEYN8h2c3ciRoOMrg5Vk2ZI
qr3ULLg9Sy8SxI/2CMFzeV6myf4R9IeLLMfAHAZMj1vccecCPVM7qsB/M6mF1LQ0esql50HhzARQ
ReMzmM7+IGdldHYw+BdMSa91VsGwIZV4GcMmXU5EyG4HmcWjPmSowjurbJEQo3A6mflsPDoQIWlm
mFGQoznXX1tpAFNRkUmYgUjSU5rdtzF5kyib06jsZJISYKdHl/iJdzIoORqTIV9g1y81iy2vfGSL
4oNq0/vcaXNNL54NIlsCfwMSgI2sEuH7uLq0Oad2dOYGMEI9hPI3DrjchU4k6+z+OSUOBdFrFCve
b5T6gl4Ss4Eegutoly0dbdWsMR1FoTfa9QP9BMDBECQm2BPjDRC0PS+A5kaki4S8j9xD87keTEkD
wcNzgU3IvztURAMAFOy/JXSPEZxqVMWdbWclVQASjOG7VrvdXTOy2pY6eNqRAWCMF63zRyAjcRlK
XZqtAS2n6b0tG5ybjhUyrzzi/B2qA6zIFXhJkWSkDr/cF6dZ4sUNnpyBfK43gy1ExA9JKhWG7qKO
6MLJkZ82PHnekUkzQgdiFPgKujY8SILuMmURlNtotiDMwD0C8bIwt9r4kvlL/zhhkkMJ6J+WuXgA
LlEcaUmadQ5S+tRMi08LnTOh7tsKDXYNq/X+Q13Yd2Stgnik3s49F7wk00Mdh7ZgeRaiSY2LeeP1
IUo6yRWxFSGmY1rzxVNWk7a831u6iX2bfVMtoVrNJHpWIzeyNY9CuLcjvnT36+yvPYUvI8PqimV4
JiHLSQcbO3kJIEZeqLZt92AEVlta2xKW/sgKDmNKqhaxE3wH6kmoUju25TSHjFKyZE7I0IVA3vQb
3Cwch0Tac8V0S7eeR3Y/lEo6WLZb2OuVPWX/M4DbYjQm6vbCEZZhU5LKPM+Op/lLdtKLhhIOy5oL
+InyAQMicCt7Uqf2pJFp8jvTHALH0RDs3IxFuLs4DBpjg0eqdcSJHpmXzBhI/DKRuDj0EwxQcVAG
lXXxiULhISTxzst1fyDie/dbO62y2t4BoYKGkZrtYbceSsJnvio+uqNRbTa7pMqgcyp5fHXDVJUa
ZABXoeS1w91Efdq+8mJUpFN45rSrVjgiE/LWyu7JqGVoiY7JmXQdaMbnzUEw5NZpjdtHemepw2zv
aJi+xQyemXwpvWkNKUbtVUbGibkICDw72VSRp8eqK2229H7gpT9BD6H6290GI4YF8hGulM8+r91s
tkwD/W0n6RgVp5ZPupqtifGdYbt4WQ17X6IZLGznk0v/wOT3N447kU/XmaXH0f1LoyNfD8SgX2/m
Hm4s20u6a9C93bwzB7uq9SChohPC7mSoAvLhP3VDfkdNu79rs6F0/9hFNPtAoZy+VhKMs3eMv/xs
qyTe0m6iyBqgnTxOxpgX/VBc8aqYAkTwiYDWkqjvpLhvmdpOvodv37TH42Taoh5bG2EMiOxMb5pT
FO0fRXEox0cIY3xZmmRIL46o9+Oq/hSNLbMLSe6IH9x4eMktOhfVdVIolXs72YPISFDhjnhZh6E+
tK9mJuW9Gan6i6/cww9dEWjkQqAxXqWfhIeJoAa9nbw7/rC/wmEhZE1XqBTCJCVdr4Suezo9be5K
ivXcOwTBUtJI6AGTkdRz5RQnD2vvdK5NsQHj6OcOo6v6/YdfdW8WgYkv137Qq7JSh+rRub369Wna
wZeqcyqiW2PlqGBkvAnSTggcSkYN2+jGeXMpRl9l/h8KidRlLTc6wNS1bQ6m0hjWtC9tVXbGU+pZ
ThU4F0HT4AyejAMmVzp0hih54+W2PSfWgLtWg3rP2vTV0jFM9LtjSEd6EPyA21C5JOHr5eWjWCX1
WzllbPNmMGfgP6sDgWF6iSgRr2C2ofoP/qjvx5w0LTiZI7mrvnv6AwdSGXFaR8H/goJsYF4zKby2
8Wd8BBvVNiHvP1gYX4GAiDwn3gAAmP746l02Cbtl0EzMz7x8xx0rXVVkNm5/sCNWgdlXJMBJLbD5
EwO05iwv0pC0tsWM/ZxLp9EdTlJzVNn5qB1vAqhnl1U8V539oDDgvRc0/y0CweF/Hn+oN40eSYKt
iRQYM+2zii7ttxHKK4b+cdkr5NgQCLCsi/b5Ne4jgQCEwo3eM7LTYB+P3xz5yR0TGdJp81NHtpqw
dOnzksZiWxOEGlGKcbDQ3N5wMe5K/LGeG+AxpJ+uLsH/DDgqRbbwE/U0qMU1vhQ9IEKPmT6VX0OC
HRMfp/E3pPaEjLFTpwG42GqfCjrBFUKqYNliS/YkmeJFoJvEwzLRv+hVZ6x08NZqL9RjD8EGFg+p
DKVB1B2U4rVHBkFWNS6Rg7fxqi3EH1HmyQOSApe7RZbRLB2ewXdkmV1wLZhJmGUQlUrPvGxdzM2G
VbRzZyYE0pXj4CsSN0XGbmHec05Amjk/AYwJeetxRNk+t/o5BUEDJOixpbBqi/gXUzYQ55UgDvd1
ORht934KOoRs3if6Jr+Ds3z7wSkyPfBb6laI0M+sPcWG2sOe2X9u4bDmaN4OjgDTBuZ95b1e5OBS
ZUzBB/ZINkSbWTSuzezxmeXq1SwK71Dyc+yfdhsFQrZ+gV3KQfHVmy4m0PvRZcL0UMsXU/Y/KreB
LPGO3WWppkD6WPSLvSvhiVx8q8m+uUQ8OvLBrKXuvcArX8oi6tFovIhiIQQkmg6IfeGKCzK6Q+Rj
yaDmY+f5Z+DUimUQXlRBRCju2KCVuwPOnfZJ/7LJiBdYNwTqSfCZfjYuuMmPV2DDPATl07vCGfEF
7SJN082IHZjJfHBt6ljj5iy3C520l0JSDfZl3pCa87JXJB75PSwvHMNYI1taVKzo9Y59PdYjbaWX
qmB9f0Hsi87W1Rsa64XpTrM+3amSinQEel2IEIj+fc83OduNlsHyi33LRGQPnzX/WNv1kOdv+w3j
Oke0UieBnZJ7S8i2YTCsQEuKcKIEjpU2JkZpVY1lT+ulioiB+f/hsk2BE+mg28NvoLw5lViNFxOB
//SjZ5Mapgk8bblL3u/XS/NyiLhc0mgpkclZoqKasH9Y1QLca9+gFZaKHKFy/ihR9VWzoAvNZ4uV
ZW1ZrKhNsOOG+TyyVQPdnyn+KTTrsh+LoeMG6TgyG7J7otEdgJrYGz2NFLeqSzGvnha5cAvT2esi
3xRSp1hYqKWiDr13rdY8QSpy9fx7AtwTSNZ5wO5dHAuuOvFdLFuXgDJNlhQWmxze5UfBEGtESpIE
QRHnehbQEd5vt2ox25sDw9/0qAxWTNdDGvM6jgTVWTcbZ0spbMEyl/XoijG1gV0K9LIX7qN0ZWUc
CVTetzWkXI7V5+QDapB76g7JMC3clMFsja+CvdHlULEclb7gadbx1qyF0KyQxTA6rw3n/qYgx064
NHJsQN0NtLKyMis8SguoYWQJZywfF3IlmasWk9/uti/LDNT19UozYuZQ6AQLCNXBoP+PFMjouITx
ymeBHg9qwN6Sl9uRP5eRRhRHITkPgGAyvDRXGfac3dfan9zZ3rKkOmzUiKg75D2+pQgPHv5cJh2D
wkPc1DULAiHB9zBVDJ9NSPjbWH8JNrOQBQNmhpzNLdULxAiP8znNY6LGNgUC++DQftVa6xJ5orO1
Mvv9ALr2DSw24YnGgmOfB2pMBGxm69jxI4aWdneIn8S42XLhL8HXbfgFoeXRypavS9TSgvOWHTZd
V/9Uv7h98lBTqojUJw4637LJSNNhl/yp2NQMFJZtOIAqMX+jnpTLiPL+r3+2f2aRw5AFh4JoTxJJ
DZO2Sqn0RmypcPs8acxcz9DIL9w17IvdiVP9pjRV06QIUuSiir1Q5+cQIX08sO8Vz07n8nUy1bvb
MxOOeoRw9tvnqDZZ3ZUD6hEazuCiuWJpRwMH+x3BaIp/Gk4mPJYYBqujoNg2sKeaQknwQDd9+U2b
WjHRnP+P3N3EyeBQ7tqISVqxye53ztRix/Von0o82fFp7hAvvGsrollkikwUJdZB/wSKTRVNWhau
hARLyqmMpEM97XcdDr5EoEpmSXGE0U2dfrkZl/qQGeszpFQvVuU0tAyyTSdRBKW6ykya5EVEDjLi
kAe6OQpD5icY25ZODyes4dnfuxglHITX8llynejTU1YC8ZmZKlNBoaMUm5vsh3rzUL7hOpGm/XBm
uP3rtVGkXEV9lub3NvAtAuesHKU+s5AasPflIerlcXD5y1fJ1l+tWZijLGpTMLztWK/x1ef8g0XD
tzbrFS8Ri/RRsnFEx7WhYS4esJzjte02coo0JlqQovgQUiuiOWjzayWCY1eIJcts+I7xUUayORdN
4ZCHJPF59oGX8xYdteZCGlrf83lEIbnl/WfDV50k2bXxtVokgknCWbptl6veoJHoMb2sbnUo+/r8
WBhw4YkNXI7S820dGuguIiPdc4ZIQ/9LBv6Y/Di2MvF0UpUUgV+VXV7M7XL6P2vmh7heWgKeofD1
AdX7DWYv/eLGL1FV/v+jDkTp0Y0JV6Le3HD2GZj5LzNjXHHz5hQf/oD6De4VYuPB+etljSMuJssj
F8d1HTagBihuuA2eBNIiNUpccLMp/kCr6ktn4igNsN2NB/cVQ8wOzaGjLcRQO2GGzx2l6a98TvHj
Q5lCNYOyQ+NirGFlVt0qknNFWMclloEqWljpTJlHkNODEDWcQ4xpoG3HRgiIZbWnYzgxAxUFCl/X
VS7g6HxtUY08QhP78oX449U0y4q7bkOPUBwvRJ87J5MRC/I7r6xMn8yEv0us1ATfZXO++/xsBBnk
6mmmEugr6PV4gcR5F6PCe3JA6zOwq6mOxdeS2bCehtduaTSBvTPvSUmTM4r/0X7EO0H6xyOGI/tG
E04sqHL6h9/EaKNLVCq8SAPGKd4YKuhuDRwZpMW1e+U5AU2r0Fy840QppRB+BT2qtBWVE4LNqOFo
3vSBdfg9ktN4hmg0CNFWk8+vHvH7NOstjzm5Ew9FZU0Rt/0D6s9udv0ECsk3FqkFD31/+uQEu1Qq
wqmdDd5GEr/C6zFVuwabTnjYXZE5Dh+7lCy02YMo6EXY+7N45UJuHDQThjG9KQ1uIKokzY2cw4aG
NQ17hAWce7i2kCWpygicBML/aI5GwklyMIjwirtvTCTwi6gO3N5bxJhxbKvZpLirtQgk0IMHG2BO
3to6psHbCkpWPCVa+Jcj6B3NINc/9UEqlGDnIqQGdTJWQwZu2Z13psnTrYt2cm0mBOuw8n95g19O
LRBWKT4/LFofu47+ylMiX8300kc5JPkmX5jLKORmmbvTpQmSG+4D04P/QTlPLP7BzjITxczMl2vf
5xW01JFJd/2k9c+YxeMNYQlgjl8gnP9LLtQ6aKh+srVcgqVtf+LBpXTBKinL9NMsDmKSTRGO4Lpc
PZrcb/jC04LASzGTBLhe2wCsDPgzaKxpPV+06Yp+1qgbbqdBzmCg7oqHICXQf0hu5RnytgTPT270
dV1lz0rR5XWa+nNTiTVCAU7x+hnoPpwvUhVZQRYCEVxSP/OGbPTwBpNN9WyC311GofJxK1HBnk0f
VOydbVc0Uo2bzH3p9HsdItZXtx84jeO2NM7jVGv5HWLFEk6B6Y3OITrEbIxQTnCngnbTwLQwqfsd
rM5LO6FHOhldpUxhdOMulkgaxto5cBt5tXmDAIZo/6jZmhturi0dCDPl5wj13K1s/wXnTEHo4VO4
0q0wWdaRJGqcn96w1aKKdQ1DYLuXdPq4bWb18Q2f/D8KG59t5JHcsirFpIA/e9FhFzUamJE+gq31
i6iA+VNUscrpKCRgFtE0MwnLHGJHdQhLr1bVvS1CLZqLpoFRABVDx2cyYfgGA0XczfFdMMcTA4Rh
W5UBZ1tmLXR5NZLb38i+61qlMntVl7QFRemBzcYmo4gGgeqjc0/VBzNNxQrf/YO9CZBecJqKsvwE
6+RdtG/a6Uvsof3XXzsrZsmxkAo+gyBm1I6u3mRZlR2hACqzqNhQfXSHN9UqAXf9C0dBKA+VcIz5
1R4rvwKccy+R3nZGSB3eyaWvNHkM2KfGLZwx3NuBHaO2Va7L719WPxhiCyyrnoZCFjq44rEXzMcl
8gTc4aOsyFxLHJVPSHER4evdcGUPu6YXZ5XtPdERKLeNrHv7Qg7owCovtj83aWXQ3IM0k/qhDDK8
/BlBk+95QMAvxLqTRszifrcTNmSij4cvJYXKNSuvqwdCCtZmnsn9LpvFpcbdCOL7QK9eb+UJT7zO
x74UI0E1OwiG6ve2v9DajI16kPA9uKgi9zURiJ1+r2l8Rh8VmrHOSd/ap6Y6BdXMh6ncv+Bny9BH
YN2EL8YweUWB3heVhfQQSvtNVdqygfr6R0kyvrE1bwDrsBhmMBw200TgYCoWODmiYhyfTwwemgsO
cBICPcPsIe14vKsXU+QNR21dp+L+H8tGkxLoaVQ4A86atimoSoSP6GLWwTJO7r0Qhvnm94pmYpo3
ZwUu+HADJIV9QJH8Tc9qtyuBkCLQXaQM9YIY1KNqW5g9WT7VaI1FhKRZCgIia+zeb9zlGpMQnHd7
iVopZuB2kscmg0a1sxm1WrHF1pwsgouIFMAAhJ0ThfLqMqjj9t3Tb496YTlzgLq6t2NLJSznz2WK
bvpNm2J6j7mAEaDOfMn4cr+RO0YRNB+gDByx7Fo8CBpmtNijUvWgh2/7sB1a1IrhyKLYp4C6X09L
OnrgHMMVObgNI1o7yMengt4DvLYA03mF5DKKjOb8SAyiwgPggUjA5TfXphhVWeAVnDAGMpj/BP7a
WT4QJyW7pVRSNQB+9YSRyBpZuwDW9ziaOKYjlKsz2kSB8p7+eZr2hOzD8NMNzx0QKp7oFi3UeaO/
TK+XfNp1LuQLHb0aThssGh3leqm0Cwpq3k7gVJ00S+PhbispGZbUmn8wGMkuaM+mQiIPcc5McX4h
SIG6JoLcWTM4KWC5xirODiQ2R1unkikL+c3XsrRE1Apo+53dXPatwqATYTCFaUDr+x7qM8LeTJpU
jIMzx9PiugT6Yix/K9oiVAGMGvF810Ql98A4L877t/8P7xRSNhE5EqSdvPMZ1Wk7+x4Ws7MR2P7H
NbCRgeU0T/1wwl7PsmH6Qkq1HmXL+EmadJxYSaGJxESxzR/Qu6ELtNm0pY9E7hXcxjUrfx4D/4DY
gBOIy4hhrr+Yd9QjIUy4RxOVJQK9nGd/jIqN/mxL4Ql6Y/uD4rXstvEkYni4DpghOBdnAMvvGOq/
wAqm/W1mg2l7cPIjA3r9rS0oJZDwFv+5Lyi90f5whrd6hpmerP5XeUzXsxxIOzq1rVmYh68W/+qH
QcLoAjpTYmQqhWFyqfshhf2LnhfDcZs12ahwdzGokVuUSaU5Ity3BjmuBq0SjXry+nb+M36WRPCA
wt8Qhw7A/yqnANQQ1+vAeQVLn2ynfepWexSPzq/xhUpUJQDnyuuW+HB1hWcKocq1WHdXZK3hJ9pC
rXj2k+eZKyJ0j8v5aeFE5jgbpy4dNXwFP9HywdC+2WdxFb6qeAkU0b5aMMXCOE1bjzO/SbCyu+42
FKYNzWXzocZlB+vDXy03cKMIvFlwQLDm5S5NSeEjXxy5YDEdPNUtOKGD7kjcCQ2pOhsW7E2UKUi8
RT1qEmF+YdPNKFWPxdyyB9AfniJSmQUwCaAA3xSytPFcoYGP86yehnZR+R9kWdmg3GhgV1yx/SA5
+EFD29HO4ZDo8EfI19bA/zJiQ5XANn2YQsFsNLZml7nECxmd42XckxcrdgrJOt93/IB0tlcV34aG
8vUq24lg9M4Qo+HC5h8FkKm3MXeTunf67Bfp8Ddd9ruoy4r57B9b58vT+8n3PeYIwnaiT2A4duY9
n7x1QabUdDuF0kq1iDemyqigtVw75CnnN+FsurSsDekFUkcRuoKLACXXQZA/ztdcLKs01//Zzg06
6DzZMDJdcqxzGXdz7KOCclluWr1k5P4pA9JW1k+prynfXBfqPFXCifR0b+SMrOVEFL6KEAioZUUs
wD6NMveWBpLxCq6hJKSjcWRYi5Vgfp9hhEi8D0CsqKjMnh0sFUtKy7mu6fMhzrpOA0GoLfdyhazW
IV1pYQL6gkt5+Enp2VrsdR78Y96Zs/mF8r0zK7g0qBGhPATjf/lZnQPu1d8j4Y8bTO28BkzpmUyM
m9QOMTIMNGGnV8FeYyUE2j759xXNuVJTB0BvTDS03LHA0J+UIAd4BzVuCT2Q7i9qa2nbHXs+Clcd
LvBfSuigX/zQe0EVugcsZCo8j56zQd9dyF0tDTPJwyipzjZ1imBY5vurlFfDO2nLyxXR3GOwjsBt
cEiNEwi0CSwAhtckPRA8yBlmbFOaLKwgwBM1+2MNL/sKJUTOQJdtrk3H1Y5yk8TvmswYze1aaIlD
uLO8/CdhEy4lL22XyASNjGhsZaBRYeAUbDa99BJiyo/JbJpuuO8R8lj5y/8aGqIGdgSf82sMNXcn
OJw0Mzv5iB4Uyh8Fok5zalfxRaytMIlbFoXlWM22OOCwGi7r9EidGBinNeoX9soUxsTe6lcpyS7m
Oip5WsN9eIdm2rqrgqrcHpFKXql5QWnjgkaCp2DSO84G77T5NsFFkNqQhvZeXuRVq6qbuPe4P1ZX
NBc5XVrViwP71vhGw3fJEAkzc2N8Ejhcp3388O/Ic2plLMih13mblh6TQJqIZO7MYOx0RoENlC3W
tS89hGM5GPuSVAsoFyvdg4Uy4YFLp3A16OEtIeCE4SWwMkf3yPFhFUT5btqhS56uUPt6aq4Ln429
SW8+vdpBQzR/Q/cuboSSTaZr44zCrakeB5nYYIzO/KZHTa3yCYwpXDgmSKMHQxTEqYDfb48aEjXR
WnEDUFisOiogzOF+GueW4r6k16Cxre3JiQDj2NDLANmNlhXjPFyS+61LES47A2pYzYc90fVrgw0E
qqaalDwGa8fYfMdEF2ZlOnkubpPDl2yKu5Xa0YBmgAGuofZCHioiM/cMEPukZJoIUjhP7bPmBhEh
cMETzU4vEpbekG/j7jz4oVIgDIzB84bhG1/3JGukloRCxtFtvoOtYLbPGbL9cH+RLYiojbAp7/YH
dNiQbRyw9AhEimLE9H8MFwCPVs5LUGEa0eCeDY5fCs99bEPHnZcb6zEPpOgqmNbTtKqmzo3OQBD6
06oQMKcC2j4n0n3ownMCjH0pWYTw8XeER7HbJ5kGKtuUM1W//hIQaUN1dkyzVCOeeItXUleLMrTr
GU2pZzycxfrEJzLuJ+9E7TnrjJ3YXrIXfjnjVGNiGSW1RWNiQBnFJU8QvtZRgl/JbGBpXBfayW93
RSVEAKejJ2we1cD2Kc740VBsz2prF0lQNhHe5Ldklx8HtRq1veoYxqdZ/quGN/TYFrayiULh7u4i
kFC+v+DvsVcW/zZmma2hQsYv3Xw9iG7PuLBSIuOJaLMiNrMGwY4KACu+1vL5SfWQr4zkDHTlORDY
jk185F1Li/xJjgHYUroeDHAd4LJziCpxe5goRqP/I1mNe5lX2H5XNmnAe6YlNIUxkHzGAGWotels
LBiKVLyvvLJUP7sm0hLy4SKVaRRcpsHgORDBk2c2TmrRg10t+GlA7WzEieesZVrUa/ExrXkARtBb
IhPzA/cv55YSiNfBC/+dgd4AmN3/8O7+TxGpRMPWY/XEfr/hBRPsop1aar5Ze5QuGCxWBybIXzFV
EzmZ0HHvA56y5Lc0Y29ESau5KsPLpDYTnD2BpmRXAt0pZFLUvJvs00n/Yio+8agc+47BeZ1uKbFd
2zXhH+yI/IU6lCyQrxqkin5tQX6doTG9fLwjyoie4lStk9mvAYvpicoiybI7Yg3WbhlJ/8FuXnOF
TE5wVdFIwjGxZzBnGqQe/GIVOV83AiGUmh80cy1eOO8Njm1Dsd2Wn/X6bwihvJTKuVXI/nzJ0W2t
sXEKmWSg8EfGJSWjv22xeXVldHrHa5LxpweYsHEJzuasTFSmDY0ljYN51nPCwc1YgJW4v+XFSv3y
osFa1geQFEMsRHRrC5rpCuegcmKbC1IqHTmOUvKPDsD/T5nBlUzx7w5KZo14YVcvl2HMgtdjoy5r
dLIYG8z+aojEjfSlOIGo1n2m2GbpZaH/KB/J3YlGkE8WwrH5WyIILZZFhAt9eLR2rKROJRPcy85+
JwTcLIHC5SF+JtjJzX9Ci27V8U6bo0Pnf67njsK4XOXQ8ZWRWTvIss1ZSmVw/OQQ2WPbId+yCdvE
lpMjjAk3hlMkG0FmuNb9/qK76jthA27PEANUfjL/MysAsPKaY82bLKGpPYv92U5uvAAslwNBLDDU
+EqJhmPuXnFTfMQkkhW+W5XCSYSSeIPvBs9UbegPXdjs7ET1ndIzW/aW9W6R7yNjhhzpsHEkE805
Jjnhe8Sjek2U6YwvAUbk42hhJSnHbGve1u8lGq7gnERGeHRXMBRJRLvqEjDWq22vkBqZa7Ovjng8
ZCanY+xW3z3hsqBVJ7Cf3zu6z8a3iq7SO96eVLRDsqvr9NpwDTURkTUg9GWXOHy4V9aQKw0YVp2W
wdC2bY5QeZJQigxjruXi7nsmo/2htRnuZ7RiTnf1mFsDQBVFeBOYBGhdlovKDYHeP4/MgpKj/EXh
XS0XqNp1HAbiWTV1pGbi7aH8WtSfstH7b19ejep0tBmOiC98DSzFfCmaBXY6oKIFUlG/UaGebI1x
5vFak/8MnOM/pseheogdnPoXp4+JBbQ6PjppUQip66WgLdAJnkFTEFNTmMJGkYt49L2Gu3bd1fAX
a0wLhV6QKcsuq5vlXZTSf5nP4y+YNn96H6P1Tbk4R00k8ZT5+iBDSPEtS98d4StBVmuYVur3CCfb
b2Ziafjp600IbJMsr+gnMJc5oG5krhP5kOwzaPUKIXePHJ0EZUiW8lagz31NG+/W4nvv7ZAQjHIS
q7jNxFnSnOWzApQQK6MG4829+tcEBL0/mGHg4RJngL8tv4yGlgiLEslHQYAQ7HxPLmdd8BcNznDk
50PLlSSLkZvPA9e/xxaOKCNY3f5PSPt5DJU9tTnJRwMldAvONxWlKFXvRdV9djbsVIJg3YEmpfnj
p6HADpIvI1tcQTNRYANNtIGcZpKtTWV+dZGE/6t7uEgaCSgKMWgHmz8oS88A8I/Jj3ySTgu5a94+
PWbkUlcp4m+iHyVWSOrP+fcq/Mwmg4OjBMAWepbCZ6azGQobBn7LiMNGO66P3ifaR2ThsCOYwZ+M
09/79C3ovpME1AQMylHAYN4766Vb7pIS1tUQFLMXhelDChi6XykAMzM6G6CeSr/QA6n5DbV1mC1Q
60eBxUxA8JCZ5EFT8NCokuIr/gZy4qsX4+WEtjcxsWz97IYZnA1aL2UhjTU43o8ljSOJYuHAvEN9
sP48977JDpSpD60AJ52Eps1FK63ed88gJ1dDZNoAvrxxRG3XZWUG99MI9issgnsKLJebAKSQnTlU
TVQecATWOTIbu2qBoSIa0JkKwjUVpmgjtV0sDAod5sey5UsyhoOIMLbacayltT4T2Jbb68rHfWHq
DCVrKeWLfgoB+JB09wn/Wu7/doJDsR4a3zH8+tKr/fl7tdaEL8t+0TvGCvq7wPXmebm00/AInq3h
rdexELls2y04KfNrc8uNuMriymK5JkwQHb+/0QK4avRTbGE1PHXQMsYK80U0g/GKGeyrfQ9bA3jw
KIWOOlz+MWYZ9TLRCHJMHN5kbZcameZpgrmna/TUQp7VsmKHdRkbNImfzkRdzghP/ekPRAHAQgm3
EZfuG+FUP7VecRICXqeeqrOq/Ge7Caa1Dm/wWcZDDT76vavM2DWH4JZ76WlUi6fw3cthuIw/Pbqf
LSSxMM2t4FJTgjYx3oRNVm2A6V7DM637DUkoMgPFRAHmV4sH0pvoGNfsq9E5POout7DVsJ1i2hYr
eTaZA2tJ4Uurr8FaJvkI/DBoS1bcZjTUnoh1K8bHOABZd0lQlYgLzIczpzVMOlzeGuKCnknfASJO
yUChB8YLHOpTUQPJggcqlyTq8rGgla8MHrocp0RiJ3nE0eZvmtVxYTYLyIVdJF1M/z1AvMM1t/iy
J3aDkgX81ZgCj2IWTm0jYAVDbeJguy8uwvqHjypEvKfpsCYJuHAX3HCoEPVtvRnuje8xwuLnpxZe
3KNZkufmzXZspZr5DgBhQTiM7n5nE5acFy2DZUYuGBH0/suWMbzPKkYfMoLDs6Ak5iQNWG5trWr1
cbbdPkDR07Ol31OcUh2xjOhTh48tGSSQ54oenF8VXqlUMwMBcWTEgQEtyO5g87mmuW3mG0BV5U5x
sS4NDSnmZ1a6/ri3u4iYHHC7YYsxwr01EPgr2vMiC0dCGDDz5e94770MJg6Xk+miOHrYMEuiujHF
0ETwBY0j8KYemLKC5V9JVM76wf9jXQLmOsNy5myUycgAsNPTE1yKRZuvkVyuU88TEUCOqqb9c3f1
dwGi+mg+crLz67AcCVQDvaBqBQb+NpCh2inCs4B51ihcpV5y+ot3iAerJvRvKaiwtlB7UUlSWxxi
/mzo/nG7BpZywdab9jF8TJh8pJW/nVFFpTTgrIBNGadeRrE4QC7khCLTXf6kPlcBrUTkPaIu0aVQ
e4DZHm6lWkN7wWDdqSFmY+zev7gMOULiu+RNSs0ritQy+QLw7x+8sdr78L+e3K8jY9X/V3+Lw0D8
OlNhlTIhFFH+GqhrnLepluHT8YTx09YvL09LZCuYKCbtQ3qctfqoDrX7XyySr2x26tOaBDrRNKwj
y0qAYjPR2+XRyXLJA6uJ5qrIevH19BwXogJxVSvNqV3bTrHbbLeKc7WHnxc7TngVRWiig5wjrh0M
eIDSp/DHOQHs51vA+N/wshSnhsHBeNVwf56h6O18LMB2X3QEwsnzAbIJEe7B4THwtYcjaPozfXw+
MVaWROSjbEnehXTimYUbiG6yJ7CdDx4n4xmULynry7GoeW5XUIS03VFGB/OtzjtRX76pa9iBaU7I
QN6ASZA7SSD6doTe6pypD80WBg5xzh9ZvffuYmgPJHtSdGuLTCSrCYl3MYMRuLUjc7Y0jF0/IYwd
rSJpP8QYef9dczDcIH+mrKtsCi4qNnfMArZxrcU2WE2euhLSqhyn2AVfYejewYYOG2tEoLtnmyUL
UNuiDm87JWJnhgxRXXic5VaeDoQ/GFHJvXbh8T+1uR6MpAloWQ/apT2CehQArANkrF4KeFmNaESS
LC7vffBOIXofGsCSVtpMbp8BTa1LStWsDMFKICqlwsnQrhVsNyxX6CZOA8nfFT3gBUlV1qteb5Q0
vXVB2yl6p7LscVh65si29xEOx+CSxNzVs8ruyWF3nsuLv8lYuWIq726K5J98EAc2qGiP7gy4ADXA
+FFn3/ToNv19BnL48XmG146KTjp+B8QaELgyf1Us5yPpSSZZKzOb+2SEIgZwmsdbKmf4muoA0zCK
8nGrHp7SBFH4P7sJBgCJTAbQ+nwF4d0uQBppGSmZxvSrdOOSrLJaSVev34OLFeOqkXUHlMpex4p+
hmfwgxzru/cF69c9AOH45eUwIgb73kDxLJ6Q628J+5RDlD6K9lRb3OVfG8n95cWHos5faHXVGrI+
X3KJ47qaOZdpQL6NwOovs+qk40EiWP7pA4gME9VgZbDBQ7QVOraXAD5c3xqXcld/F4XDonVThcis
8c+ok8CRDP6DIrFOcJEWSEm0NA4BnHH8mge1UYJttu0wtzfPTb5EnnktrzuAc8wfZGTh7mrFNRcH
rgQpGFvX0paKigfg/gm+IECkLMxPgLx8tvUMIcRcBhi5lCP7CKk/OTHbc/srn/Zpckt6dCNlZB7F
oOQvoU5JQHxyWdtWIoe9HyoyOckzF0dm+XssUMuNmSzEGEMUs3w92QN9DTONudrH3Msb6+rV0rfx
ORPFladGA7SxsdOKQNIbqRgAMT//eWLcm+eW+TpkKR6VhWlAhV2yCvjizWJLU0BwvHdvzFJkIHiy
lh1o0aBmM3ZwAUUwL4QzKYV3TnKJYVeTS+ZpmGkK4JTMW4M0FOYufekfLJbCFyv1cdjW/zjDLpum
bPDcsa0hpoKbkB+n8o7kLndzPcdIcphBPzjvwknUZfcLEx9hlpkqTovd7TLmJIv9rM8eW5v/IpNI
9RfpHisO0biw1GK9QoN9yj2blXtUb7eHhmaTpZiSkD3t89GUAbN4E9AERmo+0fir56aBS1YNmcbA
YV0VU9JqrUa21eAm/eNC+Z3qluwcVmyaRG4WYWeZWzrNCk5FE0lyuAke7Gcyum0t15561RJsKavw
X/x5sTJCwU1jH/NM6OwryvkDUXDHUl0vYQR62o7Q8WU3sGbbgd1ENE5GTsCcylnl8AxlUxw0z69S
FSlw/f5HM0cWSV+K/FiWljleITZHWS4r+eWEifiTLhaObcqFxYetogOajmP9tWTqOrv6R8rJDNk+
sF+2ga4SZTr6JWQHQD8KDqnv9Hfj4eQzv3VtQV/RuH+N1eujekZHAeOXCPV2U4mc9QZgo/72u94j
YqGF+F28EGeLMmkydMIykWQI9cGb5O8YzmSAIUs4eG8oeVjQ+QvCrRlEJ21bpvHXz5H/6itQ6t9o
g4LRuSn+edwRZhdpbYoUERNUJXcn+Y5nZqHUBm7llzI+s0HBnSY32gJW2ThLzOQew1joqum/7Ssn
svaVj8sYoCbGV4xFMrDv7H4iklO/sHIPiuYypVGfiSQBANQAY5Ojr1G7+Z/9KkqRTS/C3f6UXZJl
1TcT5q6svTexcCUgxCjZMO065GiR+IY+JgYAELfZyZN/SLSXukr8E78Nly7+q9my7ncq37uVCIO6
aAssZ62CR5gsS55JJTHGm/iEfO6fXBTcbwbvyRCA9U4M0iNpHiM+uxn/kOL7NGx33+IcIUCCthKX
UTSM/NHT7fvk/Hkp5c6b7QGzUF9clCYq9Bb1YEE3ItA/TEdupqVVRy/ACbPVO/uKLEIjGNOaB4wv
97TS4X6TsGmeIiCJSI/uZ74z0joYGMvjmw5Yq3YN4Mx2mLFu1bpWItFolJLXpDC+tRYuDfawandL
Nvnpfpa9pqZLaRzCRR7hDJBV7cvUIW/o9y/Mswhilze2183td1rZ7DEmzYHPhTrEJ1wruKCGXKmh
zjPjHTv9AKMsCvIoMyBNWuuBtHZQrWGLGR4RWrCGA3dmp2Q5DCYA3PLL3ZIsXcfNDVRGV2H+yb2M
kujp2GFvDHKUZYhZ83gTspuyeVy7Cm06zUx0GicA4+Sgsqu+5o7MnRbUdQNuqxE0AL++AAYLg70K
IMsFgKW7P1VwXtom4C9SSorMAmCHIbbjYtQ0STh6g0F8qE38oTbblPsoti/HA+FB1s/OrKD1YOeZ
t65mLMBEMqo9EhW5swnoKDb+f/rf6I40tMxv5vSidbGBuBdaJ7c3L+cKlBlfVu8HaKtexWbdNWs4
+AAgvtv3DBjuJCFw56T0l4udwaxELj42Ta/yd3/3MvJoKGZXDWtj6sWCuC0OJPsm86FOCK2IenyB
VOGMBPdUcMOGdzXRPJ6YdYISR3wRx9h8+X7OFrjePPYLYdfwHSKs4yCZI0K6nicgiIsQ9ZuW7BsB
R054dyUaO2HZgJoezVlYoli0XQwrKoLhwdUAkCXN8pq+yhKgipECLQPvVm2C0BMkW6K8B29OfLaG
5VsIVGQWwfuTaB/GC29rng6qnTDmu4DF8F+WhB0CQkdYrIvHKJJ3iYI8T1jL0rnTq0OMbxno/BtY
MNQyHWFq8QpvHoFr/3jRUF5I9gt+JOA7lcbO6sbarPOn1ZiIJW5DoHkQ6Qharyv5WoXh8Sq9TYCz
3MH7vm/rYGq+xqJlcRudUZC6iLmyRfKuuUYH4GUjKGmfxGMTsQgjXzfOwjYUH7RTrhDhXXqWCW6j
dyzGsZuQiRyXSIPm2dbV+aWUtFVwCZi0dZVFMy7LwKsbXyY2rPZR2NrxPkMqtbmbTXekoBg5UqK5
ZUCdIVPHx0x7hED9vQTxJJ7AvAu7ivOpVsKBtsf348RdZkUenfITe3pBev776/a1/dkJ+B/LpNXT
3KcLGanC5GNTF9oIovGUgRF7/xSvLDy55FvUveyXj+BDrnLb7gb5irSmATrkSkIBS5DkASUnEOzA
iMFr4IzX2ZjDLlLVAX+BQVDG7MNx/O9WOPK7TT3FqZmMye9J1q573+t7Jzaj/XihIL5cDQmRZtg/
B/SpdA8KkG193SXJpJ0pctxGsnio1k0/8IIgp8bMVq444T7UtqLol2XDnaQFyM3OKSzaIf47khoS
SSDxcQOPotsEMqw73uW570nlMNn4zmcqvYxwAz5xzU914/+fx08te6dt2YRhBQ2kV4GVA7POEq7j
4S6hNRLAwfXhLO3IZ1V899vJEqOHW+HbOFJGAyhm8ERryhZcTjUNjPj6kaYJBObjuzSNFs9N8vBS
yuPyJjIYonAbeQ8/zLPb9V0xGTcu/zE9H7SoDpIniyZIlAk4DX9SVZZzGB+6OU4Ji1cG582qW84X
6PGNkEJH5t+QMiCs/lMIxrb+hMdM4D2oGDvPF0QqwR28O/67p3nDzRSPfAciSSBnUzq41NnmC33k
QKLaSB5qnMG6pNH3WZJiRyElE7ShAPg6tPGVbV6pvjqwwgrYv/dzxhM7MValhtQM8zPn+bxuKT96
dnhJ5WWP17VEgjS/kPA35TRcd2V8UsiYVop3FryrJpR7/4X4eVb+6BGrzi/C9kbklXds1BPQ2KC1
nnVOhRgADpKoYHs/fiSpWQc0D9g6nZYGhVhq7ZeBQS++0Dzigz0bPHI/Ormofs43Xx8mCZhXkyZF
ZFDdEnaPVaEIQTHAlRLyuXwEKRSRweLVJRu3D7P++cd3Vp59wk6WDPVAS07/1H8uUA4L39IbP2UP
2XrLkxehcxSFN9NfzgmEHo64ojxmSE70d6k4AmbXfxn7qQ5U21GeMY72oFot3aI2vECXo8GPoys7
vTuHcg8jTYsByLs8axqN7kZj/H/dahrNJrbYmW4dFTKzk2xRkTJCZeTv0iUTLqTPTsYhVSOuyfRQ
FzpXhJVcS8EFQWm7Q5XHBCbCtQfUDJq1QHHz1/o+5IckEJ53sdBq/7mEa9158tkMaVikt5yi5wLp
FRmTeOq/8nVSlC4wLBAOVRu1dUF2LbRM3S1KA/HaCI2a8MDnghB+ZzGaWm4LqpD9dAibgB8DC+Dq
YI3bsdZ4kIL4jR0NcZfO4RU+6SQwWC2COVWazsdiPiUaHBEEoCkPlgSRPo42q2/rckmGrKcnRoDf
S9q4F4zjfgbyNsF7K5EllIPmBkVcScg2+rkQyrrXWmOxY7eM6HfoKNiX3fB6yQv0JISvS+/+LdHj
SYuJsnpe9xmgcLlrxIKJ5bxhMC7ObF9cI/Dl4UyJ0lC9VSLwY7ySfvlElJWEHZPtdWdIbDz3uSFW
6J5d28fMYLpsEV/PmldNOS+bKAiULrg1Mb8OlX++gKutSsFiv77EYdpZuIKXVGBgAQJCPmuNUcLN
TBCqnZ04W9mX06kNuemUv9zCxY8Ge7fhyuAqv8G/chTpOX1ybnfMD5MEZQGdhq8i0x0Ogws3CTwl
q8i42I4L/SC9qc5CP71ewhe1Xfh51q/cjnzGh8273dIlZZ29KQloP1GRhwd7KCT0bSQn/6e5TycE
D1OQxS0h2N44Gvjr6338o1mePpuj6ZdDZ4qdUTHbAwD5YZiC/jL63fbHn3bkb5ZfUJsmNz5+zpk4
VVHsvd5+uQyuwebdoTRyJmh8quYKNSSpgs8k0eDHyLtqUj/nwvar8cnS+PwM0oXIgOBk9ZI3N9rM
i/cLw5OyAkCh+CrAOvwbQlj36kEz3RcBSoI5Uxie9IyDX9e8JjLj5d/zbzYsObwhMVzEBlvOk1oX
EqJi8tlPLsYXrbZArZ/DLGSgTTcgbIDm093Pi7fYO657ZEIqNt3Nal7S3qSxmuDFpcET8cjrgS93
Zh3zSJ24+0qrbr/0uJWocMd/naGoux5RkxIqsGLNjpN+sRGRlQ9C1/6p18dD+Ug6yvLdJrW+UjuQ
lRu4O62VuYpKtxT4Hghvz3CiL5vSy5ntn+wDQM4rG6YiXO6Wm1dy1iTFM9qHIWEc78YDyXfD4aI1
9W90743f0wKph4g6TSYqhHswIdjnP+eNxw8aJ5m34JlEWvEsBhn6ZkIvKkQpezYgSRUz6kER+6k+
Z1yhp0alOAKCfdDa4yc4nnKD2XHM9LPam9cWih4g40XAz+aoEx+RiIE8CY1mKskbXsxGB4zwh0sS
9mohT/b90lzhZGVFU1ywov2GmuIHmxd8s4+W1HABjx8V2D4WwaPN+9+YGq3jzXHuA1gGFepM6UA+
ARxfNIRoRPLG7aRrDZrZH6fWsWxPYaOai6pMFWph2uAnpYlb+KphxU+aUD50bS2xMsBo9UD1s5RQ
K4fvjsdk604gxiyfvWZouCx0m9lb+QcfCggMVUJvgAuOfo2Wem3kU/8dGxT78CbxK2cHnOkJe+T1
5xNiDHvQOUy/sOmZkhZxmmar96pnnZ6BznfkkIT0+l7B7GV1QwoCZ2yNTuDHq+atFZB0EKlHvXSV
5B8ihjNiGfNuObMMxbeYLxUwVQ9p8gXqOMh970RTsrotEsu3L9096EDkAFfhYg8xXvSomFcU7dt2
zUgcuiLmwCtFk9/rR3yuF0etY3GWzxvNZRuiNwKtXcHfEw9kNIv8GVJOoo1Px2A+gCPti+cSHvrb
eZusEKh1cuNYhT8NyKoC/LQGlUidlO4mMtwJ17k6TR34rrUM2Yr9Yl6Z70NYXJvxit3geastDWLS
IIc7E7RwH2UM0wyyd3nFOj0Vwu6X1xhdxUhixpp4GvbV3zojQpzNJUeGoBx6h79TsU+1o4ZlpeoN
VAhQLBGWeo7pibCLgxxPpi6w40FwABmBiGK/01PgrnYRw5xmTHAWxEjeIWwZ/2i/IE2VD5NWIFnO
tRiYqHl+iYCyi2vFcm6IK44QYuSogP69OzPmNS1w1fV+sncnUv3XZ85oVBqfqldWTlT9qsS4KNBT
f5ryAY37SBxyp/hok3qLYez7kfxZ/tmihWg666qUOzlr9/06DZtjePGCCppNhDD1sqSqrCPNiAdc
yC5fmNul191vXgFwL7I34J353oZYldyOspmg1/GVHs4khLDAFTgFTkYBlDdQT1tnKkM9/+fAc88c
l4tdnmC4AYChE1kkcge7xlwrN/An8xeuHDXtz4e3LBKu5Ylhz7M1DpuS9CG/8mWC8RSxUXYgYwor
rvRJEZm6sWEk8gz+TGkTauHv3toGkz+yMspyMUr5E+e/CxQZMnrd6ArwrZv3GWqhA6Jj49QqcwRD
pqQGBxNn2GZofaJpc3+4fb2oUm0ab5xD35t/YlaK0G+s/UlaCTt4+xZFJNX/swCcL66/XGi6ao+N
IYoLDHAB4cyHw9+agCldFeTtkh4W7JTeWm+wEzejmpPetQkYNLCFVIAxLBldZ4xrqF1cezj0YXW9
axj7jJeoEjJgfKCHRRZfIpIjxjbGIdangtSHYTnWxbzByyVw/WohmqGoFK0saYE/ZvtwKMoYhbGA
BTcfbG8HPDJ0J4IFfW9Ulc0X3LjjEv+ElW/GKcR/kotXcNKE8OG9CNjMEIeXnR+5iqUvARxk+pr0
iWDPjEcMaTgBVN/zPGo179HBGxBaxmnOKiqLJUnE9rV7/xxtsqgbawlecWxRnjuXEugDreA7uAak
sFt0xFmmnTQBEuczoCaM+fVsg5KOXJRlMOPslTZ5X3hp12G18VQ8FVu6QxrBHLrPSe2OvdjqpkAk
fWs7iKwe6JgBQBWLjgJWRxQeuWl3iL1UNBCD4qj1gLVE+OMdWGUuUi301PbEPCWY78XnF0HRgmzp
d+BHjD+9VaVV1AgvO8IMA4h3GR2kOqswKX4PoMhSWgQRy3MyGutiMSPDIJ5G8TUK80C9ciGp4tl4
rMHZ4THh3VSmEx9+m4IsiL7P3XH7kJ0Sv7JUw1bljXqdFuWK6h9f9vNZX70CKxUgEptALG0ozE9c
aYeCaifrJPZphMgl07bT37I9OSAIeweX2jaGC/4/SeamiHnXj8xWfKJZpa/e3vhwlw931YTRETW/
CoTmipH369u6gojj4Cma+xMlGiIf7FOHsfM8lLA5jLvJoJes7je2eL1ReB9osyXzFSuYIU3iply2
Fhk0nZhQLO8bqMh9d7DnHX3sx4nLxjiSQGZilKVKPOQu0C7Xpngo47G5Q8retA/lF7/jNnxSB9yX
O8jU9mGcJ18DEU4wl8TUgznA0fq4Qvz9NmhOCcnESiU0GgOR3Vn/mxo0Xqxj8vZRzUOIVfs1WbSw
dgna5CuY6lqHfusJzw3cSeArlfm52qmXmow6cJ5SiEM6XbFJdXWEjcMOfUoHbzyE3T7dzEw3aA4W
/b6ME7gPpZWWV+QHYfeMsepLjZ01ncjkmpT6vlFoyYfTIGxV+yG6Fv7CdY5kgGMUJTUPE9RKqgjZ
WlAMAo7GX2AIAT77twODSomfmGzrWdw0koRjYbbx/ZpjU9ULeD4/60nsOunnCqNqkz6q3t0YoZfn
E0OXWlicHXoXsJa0JxMU4aU50kq4o8ssZ5pR/b/Vr4KVKJIlR/YxUEKOvwbQL0/rNiiFAoG8DlE6
Zqwfbrtpv957JfEyRqn/xkeK9Tc9Tl0rgO8Mp5bWzLXf2bGrrEIwmNQm/17WAD0A5La34OgC0+cj
h/P7V1Pgj1LGFpGv269YDlNW7ww+MR6h+rL/g7ts+1SC5b99eohothFZm1Fpsi0Xpjm7HIEvSNNz
gQ+zeGGvI+lQ+2KDXylVheHzas/KTYpZEd3/j6bnlouej6rmAL6b4qH7Y56ieipSPWjVJWb6/r8l
lZZ5fucqMRgfc1Q/DWkXxWqL3xPtP+17exsS4StkZGOkeLPowQjd0vcOn53h7gYXXVkAlwKRH4N/
sU7KdXngZqr8KkxBJAxNvy1Cv0ZovRyxVPBr8WZGxIQr9JdF+/t0/56fftnNb2LcuMSfUH++sbjb
fnYKr0d7Ibm5O31GwUfn1AIE3FyJGEa8qH040QxOo0qVbZm1/4W4Zm+3tCMY0Zv1TRopq18GdkVK
bd1yKeEaTD3KSrWIKi9QetwEvisLvsTd993girRv18hN8QAEVODjeVkgbOXcvh3BsGQe/FJ86dk3
c8LSUJImDIipJvWTCx60Y2IP/QOeC1OCs4dDA6OGpAaMGbCa/u+XtFRMDniayIh4CUI0u0bzpfkC
w+DPuAC35Jnsf2HupZ3nDCSSE0CAKGLJaq4+ou18IEgOa5r586kAi3wmPDtmAb/tiTYaU7Yq0GWi
PJ8+khq4tTgk3xZIoNeapoclzCUuXE/dC9rS4K52hKODQZm9e6Er+p1nWQm1r3HaKyk8DwqgBIOp
tIfQHCAZzTrPQEV81qgqDbBhTxA24JSbgk8zpAvvUvAquJ0hIOJJpca6rpqKwyPYdGKYkva7xH24
wUas7bSa/0fZ5DZXjtKvv1rEPVismkfEEXVWXRby9BzSYrjoqbR0S4v+WJQKqVqdqqBeknLi5dqj
Kqbleh2z9qXs3hZTbRNkRumXR1blT5KzgSU7qiXiW3xXvt7C4WYFiMIaagFObGqjcEWWA3YEqZ+C
9n52IJCkpp8+tYDYVdj0vQW3/viUzBFZH6Yg6fY6EXOIWcD7wF5/7DGnCy56VjVwpCX1h4X8yP2k
5F6QzgAGTe9q3TZjsGfi2RQX4MekqXDkSeyScOSdpJHtfIzFSCA37T+sJxvHVqI4YjaoF5mo4O2O
q6XCftKRMl4BWhcmTlk5e+rpKG4LRwOgW99WomLVQX7ku1Gjx0GLBYegrtayMbcIRc6XO6S21XCw
EPRPeR11rmv5SeYUzzSrn8sTRmBtyk/ccIhUdW5kGce0ZO90Uk9YJ7/4dtGczCLm6TXwc3APvYNJ
SFMzGk+1qibJI9TGKWieZRiAcXNKC+0vGNmvEzcOEy6Jk/+eHGwzCh24KRoIdaOSHR4jC1IMnYgy
O7Z63+a5s1cjXglA3oYrjoDrcxVOdYSBV7eK8mtrcpskAb2QQjEvVeiKXe9YpoEsHNMSG6lApByQ
0Ui6z/YFaZ86/U4bN3IBmU62siO0s3GtLhBio+cNUz+/oBopOluo2c+XB4HA3IoepDMB+Qtag45o
zzNvai62r2w9DeLcSpnNGUo3dC2CTC+qpOPEKX0qqPqd4v0qrHi4nej2B7a+dCFEV4403mhPCg3K
8Y8wyXxtcQsW95qjYlGm7dQRDTXaV2uc/lSXRewb0l7etRF9CqCf6XAZCZoSPZPZkBFWTFP38ZRN
rAbv0tjgNdvAbtvU3RefVI+4o7utVnkanfiCt+udF/hwKTLhvA9aKG52AfJzr7ji37B395UcfYbP
1YUGMWtESyazn29Z9kg4L42XXa1q9Mea4eDNHHqu1tfPsLk4JAIlnLoQ7Lp+kDnUWRH0CN5bFVdl
v9GNzBkkW/m8KVxoCyhWhoO/xFwaU5C1DwvfMa8FwoFhcZLeV9b63w7ysJSZShZRVyDD+XMNEqDl
eL/pwT4nTRBUhCxpX0Io83hHeyffK49xKSGo9EDe7BIIkalTccSvIg3hIykb8Uz71CIAszY2XZ/X
eqnKpOMpukusCwNQdyyZ2SN1mI7nHBHbeUFJyF/qSQlI7WlvoNUSvWpfsdMulzpK++wEoz1M3ZrH
Jw5tWz3ApadVG+Topit9Cc42AswIQbwoCRd6ZzoSyiYiNP0TsUvueiUgmCEjgMZN9vrwIH+o2J/4
5WBZNqpoBMWnDXTeUZFfFDffQI66uYcqM07/oevljyirmR1fI0pcL9ehsLoq54tC4mksZBNu52+s
mmOzqxYvdTx+C6npafczhWb0wdCL9uo2C6Tk4GjmfEStF4KDEGJK7tfdG8yHrbmzlVIxXoYO9JWR
bABUnD+hMA+0hEU2WTpmb65FH1CanTxjiykr5T1c4soQGS1PpUX/RDHYM+TJWgCy6YTuHAWYXulP
wv6M93JY2VP6JOLqkGOMro2QSakJPB3NxD7tL8VVnKFsuPQEYoj/p7EfmzFvfJPEtqSI8oxWECY3
1t6U2PESdbqzM+DLiw+gUWyTy7qeF/LkPSgcNold4vDXbVNa9dJE2SFNGUWLdcrMgRLHEFw0iXBH
mtihBZClt8GLHm8mu8dpaL8VRgt6yoob46NOdPUPqsXoOd6NMgDFMzg+HYnTAv4iQ598ne3ICWZ8
FsytwEtECT/usHJs87FByMWrUALruT3qBm/snDUmT9UEkYy1qM6xs2z0z+3zJ0QJrKmuvZSM6gyo
NNtjJtjOa30vLi5KgOKShCOGr9ye462omnSAHmvRs1ilryVUtZ3M+bxXMpBDYluD+uWX4QGxqL4f
O2gX1ZzYB6ENFDKUgY8t9g2uvn+48FLTsnwL/vQIDVwmAUJ+onuuSu3RkHROeFxON2GEuLnGjaPV
Dw1sOxkVILdzbURV8urgS+wS/0QYDHKjLYROupQnxUItMR7wRSTPNEX98GywovS8nnJZFnPNGbS+
xxed29+wiH4Pejr/0tSWHuoTAq7bmsU/DkfjsG9q0p1xxOrUcTrc7UUTQrN0hKSmhvHk/fSRiHpZ
cNOBXc3qvlmudaAkmAEs+EwVBZ0euPmm+Z+54ixMfcWJFYohV6+c64FYASu1wGoPndFV+OCSJOyJ
/UfvegU2p6Se8astFBnFqJE0NSpOGixaLmvGXm8/ts+/bItEuq0kr9Yn+whmm/vvKz97yi1AWodP
qTbfxWKSrFQPuYsJWbATgw8X0zkarD7cIWl0gTOGajQlhk7Lz0HUVwPwBUS450aAdFuCKgZhPoFG
Shz5QYCX/IaAZWSqqEBkdYpjyHrrE7lwf8XYWIzKV6Pw2ZTDdJTDd5gd7/GCjphpXUp2PliPsEXn
rJlKvWWpasHLVJUbutBZRltRKinn+AVRly0rJNjBXd8OqawtnVNNywEV/sTAUhr3nan+JutWxEc+
fZeEU+8NrEbb21emQImxGWpEMji1NjyDsM1oeEyFp9BvF858yzXLgmnEz4CfZH0KwhmaqoA6rL55
t9KuQF+ob5zhQ//9DWzIsU7NvKT2NVgssDgmpM9R2d9dpl56gUzLsLdJejlpZasYIyr5/e07UhSF
/8Qj/AiUgBwTwEwacjphm+jL92fdgfNWf/qw/ytIylufD+lXvtLxXoFm8PWy2hUTA6oREJn9YoKg
ftMyIZUC3sECwKVpFlI2FsRcaVYgw6YuHm8KbMtgjOs6l1CJp4XmXRYerrTsWvMOtCPu0EVjus3I
SR3xFJjmv22+CH9PVmPO9uMLLsV4FR2oX6dlpzym2gzRCY2MeiMhMIDfMkn7AmypVmX6o38yz2wj
X/vsqMPVjFiV/3YGKIK1MemUmE4nfXWvbOkS8Ia0xTGEwLFSw5WKIj6bRdDoATRRVEfMRUKBH7R+
7A5DMTKaqDEqCOAg1kvcia7vCiwf1I4qoqHlsj1KK2r523uSHepV7R1VYn4khZkThJ/u5vxTJYy4
pk0YoOgrZpbw93TYQS3hI3m8eC5GcdazAa36tNW7Ib7k6Q0HAJXSG1hkdr86omiFThLuGE02xidh
k2w0MSz5J+cl4zBBtYYvjf+lPjBoFN+LW2fXmDp17dnNMl8g7cGkxGNqTckzjGnd752sZbapmAUh
xrEWrkJyxnEQa+hj6MYkQ2tF9c9h9WUnUiQeZM+qW1ZMEH3eeOjUt/8DVZtbKsm8IY2iirtro8Gv
HwoNg1DgPQYmCZ28xFSndocW93MU2DXoIfVDFSp9RBqSqaMdrVMMZngJRVGw9xPCYVzHPwfhf7Ww
fr9dJar4iZeMLUUDBchBV1CVniELXPqp6ZbnIWWphTs5gi/mH39tKobYlSlcqvlsavWOzIKfpexw
z0Xmy0K1zNwaCmEDKWhzJpb5c6LYFp2JBpZSrgywi/46uTCJIqPMEf54lyJvGtB4cRfBKf6GzykV
r+mYquOypw4xQpEwn+lswjRS0MJo8OTmerB3J+RFh11Lk0OJD9sWA2NGY8RHa1QUyD+9qlX9/rn0
fhxeIxHmVR7DffA8hZlmohSmUqD1/YbBMYDZVPivlnJHVoGHQDRtPxrykvR8+3yQ1awnKFb5XnbC
0d0jEXMf1NYb62j2iCj5krwFjhkLB22bburTh/x2cmutNVAeEc8TTMFifgyslkeIQYm0yJC95nMs
Ub3CCZzgacVrL2I0cDNq5DP9pEKoYLDffugyN9moLXdj4FNc7xdMXpU7Gyl2JpT4djDHmjyiJzUV
1GB6UGkbQP10D8Z1+DhtTzXxYqjBUVBY7NOsw/o/zUa1OvadbUYMgc5Fh64x+PWVRMty9zbuZIt5
DBtKAKIXM9fxi/6EsfHYgXByR7WYTxBcsUYWwp8H2sUPWPmCb7ZAEhjdS/ihDU3N/nuYPu5U0S5k
wuzejrjju4hin97TshD1+fUiZoS5R62Q8QQaHI656I+AjyjXA5LzxTFjicwb/+ahsQaRbEeckTKa
Edl9UZBwSF2Avo9Gw7ae8rpDkPY3YlWYwomoUg6476kYMTUunpjL6jaZlkV2wd1NpHA+eP+9sUgT
d4c/CYyx5f9GY8dOw7P4DAO8BDQZWJ5RdabSlQBZ5QIzM1rsIsNAgrfCDOK/RQfkb6ECxBtRhEB8
PIoHxvGCBdyh8UEO81S7tgi/QzXL6yRfF1OIAPF4oU4C5JJJG8O4imiw5VkujYZFMafv/ZSLNiGP
AUuF0ys7hMxLl34BDV11Kp7lFDu3h0qFUY76yTlSw6fr8JdoA285oPw5ublr7cekEGP1g22ysf07
t56rAWznzEd+fSQQIli1jd/9UWNluGJBHU4t1oi3gBl2BGnfW6BOdt1paOR1xwxKsvVJzILn0vHa
+IcxyvfeJzisfW8Z/NvPiPGm2HbJZnx1usGav3kzdnZ7yNAYLweYPcvAQHJTRmkTqbcyeHB+bY6G
IAi6z00ASD68UXe5CRFVA7edkXjpadQATOnxU0u7z4hiwmAWY1JxczXXjlOny/IPsT7uZeSNCPh9
cbKzlRtcf1Q6HEKhmHtCXCm4MFOIIbupUTQiRY3vEjAV25eTOECMFxsewN8uyge3/KPS40Hq/rYb
g718Sx9tHGIXGSGEgYE5y0Qsn+sF5rqInKf8bsZ2gQWTYjLbELC7n1ZAbc/5XtxT2hbqCqtIXJuh
zxJp8M/+0nn+yja2boFC+9YxUigmllXgq8lmRvoKCfXBZAfS39wcFIoZO+fTJpk1PdoVQhYWUXnQ
fdGOyZpLfunMaMd4b2w6m29YvuJVVFDOuZ0+UktsLTZTkZjomIwdD+MyiySeD6VrgyPkjvvQEN7a
zU87PdWU5kjS0eauHrGMTNEmwV45ARz7xiLpzeUKrb/IWEPAce34FTScdAkfklwVF7R3i6MWZK0q
5CGp1taupVA6pkkYV62cm6rDnJ/p+D3D5/wHYwZhPjN7bLXe0pXh4LUEqQWQBBR02r/iysm5c+JH
FQQRAD1aOn8Ds2d93EUz26rH0LrwzPSSzO2cW/kGwz+HQNiqhF3gfMKqhTfx84i2Po1WONnsnEOR
ZIbAXWTwuOcfCifRz11erEO3lqXgeAxOM5Wg9TjbxKM/n8CsVMNI2d+xZUB0DK427v2vaSACb6UY
PFTY0S7UjgBb7jjIf8RhjDlYn078xw6GINCGPLQTqo/IHmcNDwtOf+KOQ7JrFT/VS9IaGTlsibfZ
L5utKV5I6dfLGYImYMwr5MLwgGQ92tW1ozVPCERo/9+61XU1PBXn/rivwc8hsFGcmko69qrNEK6h
vA8XrYUBV/xZ71EF4scpMRTHlKLK5oT8rBehqtYazvYO9DjyDY8wvanEBblwowNwuBQ6oBrfO/IH
YDgkNCKJy/t94AbaRZddDriRMPv0jJ8eSfJAH/l5p3P/8RP0zAUVBxPwxi0njz5lSdjqzmI18120
NOZY4FrkSjEEeOUJ0a6mRJoLMigqg79R80JTrRF5C0v4KLWStgAYEZZYcfllsf7AGvXgPEBzhIlr
YmGeL8SVBEPXNhaM3xdNyW4UFfisqHgHjMCwEIIsXJv/PNxxwxqaG0/aO4ztQZirM88j+0ypFfgV
PPmm7/JihZDQFgDJDiCKxLlPmZNCFoaZr6fOs8y4BQtCG3Gvl2xTm5GbBpEYcGK+GFZ31RclEm9j
skbb37dGWjUB8JzrzO30RCvuo8PjJDNeBXK7el3jETjc02dSII+BiAvQpxle7l9sM4QMvIbVhX9Y
FYvl2Lq3CFFmzcZNZaTOy643u7Xsq/L8U4e1ZGOi7nRqKnrxhCKLEJ6NYapKZ0ckiNveabo3pCMY
byb7733mRw/6a6Qyo3/5YfTQ07sx5d6CqZ5tmajKr+dk44HUpPodHOqiw0NIqazkgwFnpXKWsIbf
CQwBijcbjiZepC6y772Nc5qqhQaLLe2tjDsrTC09oOj6nQkjoWPglUHHpieo4WFHzTEqfcmwZi2y
dutpXeUgvbgNkfnbiEFMEu5Kz9yLDVyaITAgpHdFNBKzMNFdYWbWei3cdwCcYRDkMfRlgQXzk8pQ
QrJ2DHq3OHkrBq8Do52/LSld/oreCcyXqv4HXlk0esz8VSLJUuJz99tJNyRzu7uqgjUxTqILP3Bp
KLJPzHBRZ8dlRufd0usVRlCBY1N3GP60SXuv5/ItPvUp0ibAifibt5PwjbOy//AA010gQgD8brel
e4wZlZpbE7pgc5yMFFVFa6DVrj4bwMBjo+P2sYLvzHTf8FpPZuwDPDJxpmZIB1z2uDglyEhgU919
oP3BE8/QKtytEbCGzaXSFeZxdIkEFgDffnkcgjdAFiAdspWzBJ8MuKDrmlTFRj5cqr26wCmy28rK
uRHO0Sn5x3WgVzUfG1JxHLNE05rHN5+vCIl0U+GC0ujnci5Njpbim1gu0r25i+XHWiBBzc17eboq
RNvRXldEGkvCNzi+7J//yVetDqv91eItGQwFqLMtt+kpRyYpzvWkjQ0zDmSg7Dw+JA3KGYv0gBP9
mHnxumNK7sr4z5/uYwZJEHyCV/KwI/FPqf99P1RMU2E/hbyulzkfASnUpcgoCf89/cIbLGH4G3Ns
2zFtSV+ubbnNoBCkj6EX/kENK21aiR2logEIE8oEm1Xv94dy+oi2oAvJsAsSD/ImeWXN+L+cKJLr
CMhfNfEhwEUhh1iseMtUNiehlDlLGL8R2pfjhhHd6em/kWg3bHhagF6REybQ+PPE+UgFo8DtZorK
4uQlK7RTHLn7mlRqJOXuegBhznORdb0+mruTj6KDyHEi2q76I7C5SssQoq6MlG4NUMW4DYHwcghB
VPt0giATQQ6CZeJMWeSYMk6LkZ5FrSppTyI47Bf4MMVxxCMML+m+z8ep7wUBLi5/oLqfm4RksYJo
7GinMLyuxFsGKUDpDz6PgeidNCUvxba8By4moUQQNb52rKuyrpJSpdQl1zwlH7cr4p9Guq5yrl6b
z3Irr9Aa9GPJ4sYmv68jYV1ERa4pQm73kbXCaM1MTmIOUKEQuYOfKd50N0IfEGh3x8HGwfgad5Xa
6QIvep9RiJ5ePFwAqq6rOeXHJeFzNnNANOnqtXVCXMnO8ymWMuKPk9zMzgfXcTmzAEH4s4kx5qgq
kkZkJ2ZT+ih3y5+5ZVBds49C6mQcKzILrqqsxO6v2cSxBPe/GlhS+pvdBNGYD0gKZmWcWJmUILom
NYaSNYOJWkYQlU8F0WdX22vZHQ5EzQ2N3Xa8f9b6AF9L4B5lw4TV1PqI47iCP5N4LdJqaLC66jtm
mpEZKxgeHGsQLllH7FvVoXaPOu0wEuPrhWAboKglT1CTBs8mOBrZkORZfSG6agTpdPHG+sIJrdbw
2sfZaZ4u0KFFMHc3t7Hp+BCTX/ztb4B8/sze1bbPlW9gWAxjPFp+JzKy26Xgc8LiGv2PH6x/q6mT
KQCCevGndA/7K0iPGtMtYpj5lD0xiVG7FsJL24DaV2zK3exFRbM0cJ3s8nQPhfUO3uR2h4vUm/tw
+jeCOjL68PQPe2G8HiW6zK1cVbTJHDFRNi0wqeCRKcEbZUrDNfw/ntv3kbyb2knPb7Mf5Ub10h99
5wvLxXUgRoJU8AXcMU/k9F1qbK0he+dmVAFHZrclYFGgZbqHHjINhhWi0KvyQlSGpF0KaVdzNnNO
QiFMRzpqkKpYODhJOhzhBm+HhAm+Z1gWixEZov2mbc5E0WESx1qKXrTvYydk+AjK1GOm0r1ERQkx
bV1Tj1UxCFtenkjgI4b8C0tQkyWc8TWuDkDa6jVujxXifTkG8H3L9zLU1tOCzfQpzYrCtARy2eiU
Ps9iJITM2pSQV+/9vvFET0rLqKCGrgALYI8gwlCqhg+TGSugtxNb8irJl8RbMEVE/FmLn4Ap80SL
9hSF8HAmJD2nyArclG1snMGp2xjWk+ufr6jZxVwMAazM/JF08joM50p2FxQi8jbtB7MuKRldkzBb
NigtoMK4Z72h00sHDIGeen1/9yt26vuwGmk4G6FeW1VU8TlcoPdfF65OlxmflRFw84R8hZHc5Nb7
o2/N47guJGsx7IUjcaZJusxL3XGsQuxtqn5YBVBcrH++F4kbPWzFSiT4fqzbNjerk1B3nVYFYoDv
KNs3arDjaWZBZqNlVtntsZJy1odSKdwm4c6LqJYaARI6q6pXeoYWg0PGdL+zpCTQ4Sndlt+xOQ4Y
JVxNbME3+hZ+MDYhO1JfKaycvtqzoJPL4G8r7AUrNZ7cLjgtrFaWas+3xmUbHtDuoSreNUmbiT4c
xrKIC6R0zbb3Pgp1xBuI431s3pzTDDciCbAYMR31ihZaFE/2F/OidDHjlcAwDz+NBBX7yXjcjfbm
OukcJ2k8GFC941ngFOYFR58LhZhWzHjF+tJr948Bu+YvPJC4V1tCGyY9rsOPpFOqyKZpG0cPCi05
qZ2uxYj+E1pqwf2+lq3L1UGbMDyNWSJbd9ccmJipTTvIesbZfEsyjCOGx20hMairZh683SiptfwN
CMSEci+kMSg0ozxLWXdsXFENEBgeNj+TwKMtrdAzLYHITVXiAzrTCCjy2lIAm82jOgAzV8dY527E
SKSHeRFV9tQguzk3YEWo2DnbdlonMtKIxbBVG8AsqTH2UKvj2uXSCF5cczZEor04n0TleVq46wf5
VTDbJWfPfFvIlPfjSDH4heuFyVLJdDbcpHW9gP/sZWnmsiiwDjAcWQok1wsmsMq998oFIazoZZyX
R2DMztIAl3mqG0tyZGVxljZ6yvvoF//usDBSmLOQXR6qP5swh9+f3JyG+JXtabiQ9ov5qcWd8+Of
Hrp5OUHNB6nU4eNQQ04uDtPb4kKBsCPZsrtcWHAtIDobBST7acFb7NNAQNS9LCqpTp5rp/v5GwMC
aAjSsY4U6HFeopoDO/fP8NNip9QJZdxWZoKkGEge88/yPbQUwKDRY5BS9svdUGXWlhu72kcqrR2s
S52y8xMzspJTlu6f11pbCkDTUFeNfRvw0uiEBse619KIoAPfd6aC5eSkCIZQposGUoNZknaOu+qn
EGLlKiAx8IqMn0B+fPZRpRDowMwbE/B+4Htoi5S/hhNupbdvBf4qvvJouGwBpUjsl52RrU43zskk
s31+/+Nm4K8cB3RM0KUdylvvEt4G4ypiXQ3j/1sB/cbG1iOsMbghphFH0PgdglDo12dfDZebxQlR
lx67wfY7LvIGXpnwwa+SBX3tDPslANgN99su9JC7ywcW7ucnoN0XwdvonCZK5OQeUl0M4eMbdubB
LZaaI7h/RWirIG5kVBvbeTUI0EZn4f5QFqYRYVsPzOwtf1docJEJKeu2zhZfHa4UrvydbWtjDFld
7PoZhF85HI2004DF4DqkC7WDA82hRBUflc3B5gmouKr2LPQ9Fytc8hyRhxpGbBdpdFr6eQoaaiH4
pNkrmYOOJWs84QeNlXCAObRki/hEIt8D4n1X/9qWexnKHZHmWjLIfqcWnnd6+t/m9lRLKA9Ml3Dz
alsspFdVzlSHds/aY03lluG4Jpo0fH0A2LZ2CCNPVAlA6OHY7v6EpdWtdD93sT0msHZM4AjpbZe5
Bc5tgZ9CrLhz1i5w2aP6NVbizYePcUDLLtSQb1QA23LpUsACVkrZrJUfhBPvBg+8swCri7vX2L6D
YDZE5S9UrHNY+Fx05Xm+xqHTANdYg31mBYTrNrRXQh0Ms7hipxooJldkRkqLd7lwSjA6fAR3xkDv
Z0AQ9HrU7Miw6Aiq7KUDeMaijeUGXg5a0p5LyKeZg3QVZlmUmVpZFn4AVVnQupLgmwyuN4dNjnjR
P3+wVfP2zxAmGfdbSa77/YizAkvW+jIhiSxCQPygIGsidJ5dAzrOKZr3EszgPQ2n+XWTSySWc4rG
l71nygr1qwRZhkgMAihzm6RDTDNED1jPDepXuIy+gaOY/Bte6Dpwx7NTDgnjpFpQc3Vbg5d7umyf
nHTR9/Fc/TZKgTswN+2gx2tWH+EKzvh8B68nFLjnEJ+pdxKRIyPkaaUJn+zFstTa725ElS4opPxz
JaA946ghWoBnyb6axt5bNCM2GGbOmjO6BusDVJou4D2xDhwkbhE+KQ8mpGgbxRCI7JZSaxcyY4AQ
rqkswQdt8Z4xdraTbUOHUwqcco9lIvky38icP09TFrDVnhgiBLKK4/69TIqJDiBDcuH91fH6+tn8
cj5t9jKyomZzFWZrR+giPefHUBN95N9lQkTlCDgZF0UBKMwCbarXQ8932ypibMYYz9g2mhY7p1RN
zM6eElP79vNtSN08tebIK7b/HCFEXtJyy85Fugad0faVrQOGrxLTaQR9ZrEf5yrbG2Fce4LsUT7h
Wt9ovVJGM2POqEfCLRthGUjziETO0DcL973HsbJyTwRDLDpVZ8Az8O+P6Lt01alRgUHJculmzcJ4
UznBRIjZcl0MCbJKxY6q0RKPA4Mr2xrR1spjbY7wtoxKNqAoG/HKsH622Ln6YbuqBzmEolAI2XjU
Pdg1N9qEpqwhE2wy7Xyz9oXkANlUJf52WaBGefM0+ZZKTKSQgdQgRM2L7TPHekiI/y3tar/R7yar
j3G2pO1EJPSNII7cnBQ705w0BDW8vqz8QYwYdEAJOtEomciccadIFjCPR7aLFbd+T2XXhIvS66Ds
S3B/bNfv+Hc76hwTbp9cVZwIq3ETjGe2mrm2Hxd8Wf7Mk4lYW/S/GxOgQPL3JrJsiStz+OCkj6wm
K8zJASHTwbDEidNga9uPisg7HqWFaankRDrATGvEm0PgeBhx3+AxHie0Hhogl2CSVmKNMJKDb10m
HEFiZqtmy7YKJgFf2FGmU1tSGBgNL3yciaAgZDoBo8YHFwKCMzzHDe+g1CkUiamWd1OH6YGU3WFQ
QeFqxmkC+H7W3vnHlHPZEWFL1a444pX/y0gJZoXKatBVYUQv6o5GY9eovUPvH47TrmmXQCc0ZOH4
AeC19zy76YjGtgiG6C6Vnn1EupM3KeuOzj6q/wLKD4aM2gpD6POg0aaqQOE8WiWbbGUTOvkx+9Co
sJIuMr7CV7qXXkezH3C1aJyeALzXJyY9S9Hk7VPp5kOMqZWlcV8EUm+xZM74pArmY4vunrMEoZQm
CMPmqCU+LM0hETOaWzDiR23RO8sqUsfvImGyH76WASjZUm280B/DMIS4zOnHJnvTStnClmybCvCw
iQeUSeRhxIpVQ72tz9R5KHq7lgGo8kWI7VkWgLiRhWu/UkQkQNBsxU7jllUhX0rC6wssxn2mcwZj
wwIagpb8+vGZc2LuYBPqbkQYtcWFNVQyfRv7ClEXLnd7Wz1/D83m++9rF2Fg1kvMOHIcDIKg3R1i
SPGIa1ZFbhoKjhAV0JZjJgueZW62LypfTlcn9Jl+V+j6ybaPIgUp7/HDPpCHAN3evSydJPtqzUP2
LRspV6JYjKkhORMvaC/JYwTBQ06WsSFTNhL9ME8xHJ1kXWsAgGsl3fbntwYfm0pJQpgK6659gJ7u
o27s4nOL082BT+jaydscFy/150Nj0GoNFiXxJuod2zCABinPvgL45hFQY3uHqDl08kgH2Oz5pbEp
f30zjb+OfkcTDWIxQ8WMXY6Ak0cm9NhG4UrPHu52yhz9jGtb6JZlq5qxxhKzRewtE8Iun4ZSsgV9
m9DxbpAJAzpNEEC3iL2hi+VGZjf1PQ5ZcUQKaYvMj/ZCtQFBIH+dmL4LDnVYr8fSE4/Z4Fxm2nVD
oxjSunON3bOderAs2IJYcotPZLhJLOm3fZ9J8NBO+drSJBlt4mOdHTxWAnXjJUpY02OhEChrtzD2
/eUv1TgJ4pc0F5JhAN3AHDe8xtnDldH86BhL8lqhwNyKSiK5EZ0YdQswhX5zngJ22J+O7GBO5j+H
Xycw0V4NUWKdQ1zvvXeTejjPT/wD4wurkgKMqPSC8+p24zkR2iFV1yIgL4J8NBiBPkK6erBXG2VF
t0ndL/w3mFaliF+WWeMkryGA+e/QoifNQlcqSPuy330MAjblYKHD+9Kf8m4jFGQP+19FZgRZmZjf
0spHWiaHWDI1r+aI6TxbAKeroV451vKtxOZlfhB4RsePYq+8n+IjowgsCHo/Z+ANlNt9YTp140qb
2aXLp79HiL0hE08HrfBG0OtdWtaPDkgX4ePGQsHFWbgbC8Seh2EIJ3O9G5Z71IeSJp/gMHbFfrBr
2QsI8n3LVluzrr2RvkQs3vIG8Vym2Y7ST/2aZCN8VMfhXreg9hrZBgMW49c/Y82Ekrty4XpvhQDy
vGcksqz/2tSujrYkmuMMZeefJ+4+jK1ZnfP6wWb3USAnk1ULhUW71fL8GPlgz4FzAp9xrAJq4wt+
mlXTnIs0ldJ/6lP3ongiC/r0/BLkO4mksf0GE49V1TuAs1nEjoEYfZSGbbWqTmHNh4rZUz260cJb
X2aSQYo8L5X2iMYc9kRyaO1R9X0RVkaEIpBXyzqVSAXFMGhmQWUNm0It2AHJzBEj0WK4UVNnapSD
5MNYdrEj0+e7d7YhvVzyauaM6BkB3gk8OrtftoLMKUhnKkRMG9ULEAG3gy5dkFJlTSe/sIICZf1Y
HLYrO3iFDmmIVdlDtcy7L2SvUn0wZZ92BG9BEQb916jMANjGEb1/8F63JuTz4UnBVX1FFDicrV89
MixPviG2QkngYKFZ2GYGXFoc0mluXqq/vXbu0a0UG5Q2Eb7UmEhAclteSqgeQGPgpuzbiMYU9XoJ
qAlR/HC+SPNJGJN6I6RzDNDLxmYlW7UFOPHAycP3Et9GYwALIvomKSVqEihmJ294eT0tr+1V6yh7
xpgYSE3fbiViEpCGEaTMvh4AyQOTsQ7vHV/QwVWdkGvJ8Sf71PWzO3/1HeDOl48ocbHyxQV8u+Zk
GjZDOraUjNCl7HwBXN7jHjIOWSIvbdFTaITMIfSilnilAvKZZ5zoKHbUKjTL4RpZj4MM3XCFMAta
8drDF0vuJyCb2Av5IeRyt0Cxxou2IlnJQSlo9Zxfmpv4YaisO19/bXqV6VrAIt72NLD7ORckgkWx
nKM8vOApJG/HLc0NuPhJunz4gJc5w9g+jycIAdfDp6fpqMRSlulCzlG6mAJSXfkH7Q4QXcyoOYXN
s9ITisJ/IHRQ2l6+hRNQaClVOE6TuQbYPu93hlIs8I0vgFduZ2aIJ+VDXMQa6e7Zi1BLCs5kG9sA
HtMijW084DU/7CCFTEgfBT8P1pVpYFLdS2ts+ltX+WSqIf1EcTNKFbcsbG0SmkwOLJuOQ9TfqV6O
08lSS/xJXovVxkKP5H4wxMnRqRYV03xU8VSC6RgMOIYceDyG9jZPdHiSVtsNLxtRXe4Uu6JRuzsh
ZiU6K8K3Djilfh6cMcoBcaGY0LxqUO+pulK7R6b6TF7cmZ5eJOL9KnbMhEu1IlmV053hbDVG+6yz
5GcDj5RHfA1UZDEX2hTwCHc9EtPJUD1+rVmWgvZjAWF9/oN6gMoCdEOStVtFRfCZe1ci99fWkyIU
+D7Zbcjh6LEJ1+AFCGmZHQM6QFmerYatPGnARmBvwy6ggoO+18Nr/5tznTSIrWNjKclH95wm755a
KFWgDia3OluH4POXkUthoB0JJNgz7MRFIH5RSF7rUwpUD/YBOO145PuM4027nCfZrB8aCn5TTWSe
DPTSC3lYVKfrBdhnvrK0HQerSfzaknQmsyfUY4vi9dvi4czdZvfDMvMKAFPcMVNdt49sltcxrUJu
SUu1aZCsHj3ijIK3DSePvzobzvViAzZCfD6ppv7bTWrY3OWb9WkTyHrRoO3ctE/RUzMfr+DqEgos
a28Jxy529b6xJ8CM5dWhq2pc4WIU7D8TmU5ryASOG4+qJ5GSQ/1w9Dwkjk9LdL3UgNctqbwxFyKs
f5e8Y8pf9RfBSW3ihxNb2VYx0Fv7bvHz7UW3O+i9S9K+kwMKSZnoXS/02TYUDek4mB2N22E3UaF3
6SU6MnT773hjcY3TXh3DQ26For8wixt5ko55RQVKFCHVQUU7RYT/ZDTLLpQ64tMxmSJJT3TKE56A
mjKy0VwFXwVNc/1KP59f9GltsdfXZ0+A79BTPNff5dL0Bdcw59yMUOVxXiijGuMV90wUO+GvBSbk
agN/AcouDyfFDFPFeZLKfM0Y/d5Ac6sRnWmnTV52GQvlVa80hL3v9NdWkOskw23q2aR7zZ+S/Fdd
z7KaqOPeZEdzm4bmQlFS+S6w00M4/9kUUrgDDv9QMVfca3sarsOFP77UMbBhTrpfNgU/Xc/aHzQy
tS+FXEn/AXb1BqLibW991yCdB2VUSATFH5PRIroeXUzy1Wo+8xSZXZBCysnxD1AeUZxNUw1HF9Gl
ksZt2Z5y6AcGtgE3+uDAfQ+bkiTZDEG3IPtqMmPTMyV+JC+zctqYW4Ext6FlgztZIBxuU09/cgwA
pQqjcKNZva9xAwd1sQQp6r/DZywXKS7YB/AdbfgkNmWehuMtwgjNou5lQ9+diXzgiDCoSMd6YK1D
GhnTML5n4GFonqXANBpSGUim2iV8ns4+eDAIoHMZ9AwXA2H7pWCYLw7yP/KyZyp+os6vyBM26X8B
5Lqm5jwk2d1GmWcXKUOvIjcwfHo8P6bErH6+ND5KtAk4DYOhCyP+a/WG0NcOqkRPFo7CaYynhfcV
WJeKrK8Ozqa6xmEfGX7cVR45N5NREJYoSwPOe3Ue9TWYcHcn/9tsDExoakZ+3dWvM4i+vxqXy31N
MzVEqJhKxxxboAjGZnnEEC+AkLo3L2eMDeVgMs6BR2Dc0QyfOVs+JC3UMz5D2QhoJXmKzTOLM9S4
/0Ah5t1fr+NR3CNm5ST6FH0564hDDbz9y3qFcw7U0Yvqhm9FXN6gzoWvFPlEfMf+yoyzmiMMW284
qQc8vCFivyAf0+hfggN7Dcl06KmmExpP5wMutCESbHEDd0zTzRJxUR0aAWJGm18X/jzSki+lPx0y
WLqtS4KWXWxzagZNAYBQ9qnVQgRPUxavkLXT8wm9pqilgzwt3IY4ozdGEt7ZDjxq5bOUvonALO0r
G7WN5HTiqVKYv+r3KpQV47xhSHyuTbPGMbRic3Gx531hOcyWVtkkMMbmEjlaTLW675b3fxsnEXaZ
kl1uqLQFvDyvH4R2ijMNZ/zpdU887VNouUQNCOBJLje4YZXoAtkRlZm3Ru5v6vX1WPBGm7N7qRw9
sZjnU98j9rMrzWq8JBtOlS12ty1YYqhSk0lUDoWffcVbTnl9c0X+oukIYHrjDKCDaKKTi42RYPaU
Fk/8tGdbP0GBVPDCGdS48pOFe70VtXKBpyJDgo5GZc1gNZq5+mQtO1CPnu0rd/MjxCO4bAu4qQJt
HQDI7eY6KObuPN8HENrw9M5S97ZSlda1E2PBMG7xV6uZDuFhvQdpiQlw+366HO677nw5CoKTlSPR
P1XCbEiqho33V7uQafbfBLm3KbzbAUxMNJTVyJSEqvgYIFVluw6Fvuw3JzOWgAkQLlyEcNkFXhh1
aVhERVzlm5BgLksZC7QdiNvNmaA8gDjOSAbSnt7OSmRu502rlC14iRepky4txY1UKAq83MGGcfey
5rx3UQv/94TCr5F3WTCo9DNIPwohZbhl936YWGotK66CSb5Jg1+7cFFJQpQzQcU/VRBJpQrPa5aI
h1ov7nar7+cbxXdhfuc1dC/nNdVx+1FYXmodrsIsuaFRrW0xfeK5+dQrz1syu/3qKxxv04Lag7RW
Cqc0wRdE3oHwAgNZ5Lc3UXwO5qX6OAAdbNMbEP9JTWqskZf7jCRt6AKMaQo7TMWoDlc70b4dDWEq
ff3EUTOP6cSFrdOeQbnY1n/77GaH2FWAlJV9c/WBaFbhVgO7RWH8iVuR22pjXXszSHt6kZnmhMtx
W8Cvi5+057qDmCptEEWDSJrznDgLlCBArK2Zzhea7lL24DwiUS47vvL/yRcfShJYkya0S51B4LEU
JT1TG1cm/yS6WIL4CFqLxr9AU0ZjpqROW2ms3qexdITSNyZLIjPQ5uS/bcd66S6xio2qlv+CiDR2
3dDfeaeNb3v4YmEPJSsB7xNC1h4xaLRxFyyyq4qOxHoiKI2JTr+qUumnRLa5UWMOlpBAMii/GlAY
kzZQ1YvEEfOB75T/CVylxZtRVThnK3hUtMPOXa9bIAPoViwZxSRZd89PX1iBA4kKdhxQLRH5HdHQ
WGXktB5zM5OgQVQrqZvrm6q9LQcr9/gbcAznukLxJsg4v/DTDGqbs9Dvy9MOUYcQO/TGa94z+yQY
yGeQDr/nyRvTiS5X028FtvQlGbyBKsGaqoOkaJS9Hzzqa8A8ExI4bYlGcMMT4MVmwHCIC2NP6Zqf
icMdKXA60/66B007dlD3knnU+3i9Io0woGMtsNUurrF5Jr3fBxDkhSeFdiDm42iMfl9q3ybemNsH
6ULI+CCrT7NdWh8mD7kTjnV75Usqp0TO1vSW/Dds+3lJXEAUvWDqaav9ZsLWjolAWkPrd37lYkdm
KLxOhMhcJ22O1vBcjru/nu2VnCbnq3EYOCrznyZDU/jhQTBvTXMxoPQw8LQEpDjg1voMYBxyQsl/
cqrs+K536fZhVMzDBaecD06VtuDuQ5k10wP+IAar9MJODcoh9V9gj+iIsWN6Qx+bQT27+5DdtmeS
N4gYzvkZdyEBtnCzqp5YsmvsvcLZ0OcpcDNtCYrral9YipKB+CpD+8YpOGmdqPBogxFXPUUL/Yjx
sJoP6BH3kBvC7XBewYvlog5frIz58VP3wwgdIB0mSy4JzBfLRX4Wnu+FkJ9rshI8HBZiYeB9K8WS
oB+UiY36aAVaBuEELlp39e75Ry5n1pnoAfyeqc9WzzU871X82mjltGDujoZuUDia034yVXhONJ3R
KV2VZUPSmRSeBP8ovWn+fCgW+GYMYv+IpoPSezaamefYW7Bgl8JEPSHcE7E7CrW6dRGrwY4cEJd8
K3343m0qosDNq8b0UU1bfp3NANME1Bss9zeytHmWDzSfiEyFNNrAYkR+6Sx9s6pH71n4qqcBMNJ7
abXw65J6DqCSsEBEF/ENnO/90ADdg/6mS8YGpS2/Kbwt3QMUU5nzk8KzzYWJR4gsuJyD8XWNUUAu
09MoZLGpyJmkXTG40M+/g1gTOyxbBXsM6sH5uh6Ee6cMIWsvz++m1TnbcLP4XqQu+yxh5pwxgkJG
OGeG1aGMXsFUDb2t1fssvwrFEn5aBGwPQJrig7Fzf2ltKwV7N4R0waa6z8diFRTDrOfUOjeNOaHj
hZzo1AYX5eGzxcGMtYHHWnob559w/Eu3k3xStSp8nJWFDLR4C8/SvcmMPxUmmpyplaZIJQ07Nlkl
uLOzhujFAYR/p9IRZhCnYDlTBpBvs+v/RP8h1QifHjWv3/kUj07kG8FAMRMK0xoQVxk9XB1cuSFm
ibPFKIa1rTaF5LxVbs4Vuk5Klf695Ec/8DirBQngHXtRoYQQB7z5jd9vRFZAMJuYtjZv/ZBRWG1M
+CkvkEUTg9L1J1TcX9ZAImXExTzCTBzb6i/gkz7pE4Aoyf6zWtTpv4CK1o6EOAr55wQVSCDHrtPK
uwpplUEM+LSLRvSzQJwJkbRyJRgO4YjBE1K4HDnhvVnfSn2wkb3XM3j7TNq8yjA2faZQP6ufxLwW
ISIjbdVLq30YabYpnXSBE3VsZ8ub7ws2yNcgPnwr0oWRVnzfEibAtsBgQmiMANsUByAFMj7ISRzc
amTbc5DV6QLBmNHnpMiZn1myTXFofPItoP6xSi8XkV5D1ugYLkhezg+PFYzF4J1mo5z3/vRCPljS
xMIAnq2DkUUUYdYVtW8V2K7nHE+pr+/zFh4enafDzFGBQN6AFz8jLzz6gFSFTETURTtkbqF3viHW
2yBLYIKfgF3zOX8qh2CW0SGvk3AXEkbjvNiTwJbnVpYhP7kQnkoyqYTfMmxOlGAdkI7o3aLdb9bW
HXnoH0pdTct73YQLpGBu44p/zUVETU2IbB5rWlXUQdTONWTsNRfrX/+TWSKGKyBcI1Z7z334SkhG
hJQW/G+7QgZThPqcd0/kYbFE3GsoT3ohEDckN2uYpfV2hZ5z8Ukrm82jTR0VvtbHYFL4OPaQGbqW
qfsuFLvyKyUYCKLd7zh06A7ZV2nZyMI+zl1oFjwUijsODNEbL2ua+IkUcuQQTKTi6dF3i0V0NQQm
n86ApCMYJqKwmGl/qI7isuB4NOOcj3YXTY6YcmZXwetstwxEsp4m67AHli+IURwVy3anc0wo9HRe
K/BIpaGbEJckc1UyvndWy9lhbYcseHdAh8fiVBPJllOoeO0emo4MEi2F68o6kCoZiTLyNH50UBOi
p0MLL1XdrsjFAyn30cn9d1Wq3qg1zWc6UMO1CBhAs+1z9TDBgBJR0dc6eQsfgJkSrTSpM5rlj6vC
AIRJ/Jq3IAByfburJLDmQFKbj565RgnW8b+WRczKusUT4tuegAYxwGmQzEIkMYTsBnln7V/Ub4L8
+1Rvp29+ZbFYvHsKfA0rDbZAY10cdEuFDfI8oanTj/vz10BotDCjes7JdD0fo5PyzOoRcwDSsUX6
Za2WOp6ukA9XBWangupK7i2Xz34p1lBQGukvMnzbM2KiIeKl/Ial88F7AvDa9Bhxe92e56muqYqu
uuXkfi2R4n+ogTd1sQk/gSobCPw67lXmMmE9uanBXhphQktI4xsIPhR5FuB6EllBzhxqYkbaYk3v
2jqat9qWjwr4WtRbgfFQWNDkjYdWaSTmK41ef/RYET2zbueRJvj3hTpVCaaPfPsx4ovPdYguJuzP
35bJjNNgypuue9EADB9A4/zig9kexnYGQjQ1QVdZ4wXzclft4NOIM4mMXkHrp99qebZ1Rmphw7+t
AmYQAFhquCSw9YGxrud3HTyNMuK+AqShaTGm8NQgAUZYqbOEVA7udHWZ7MQtsIjoAlP9OZNwg/6d
px685OoETSw30BqqgjScB0L5ZB28hmeHDOwQs2hE5WmzUYZSTWeedVew4TPB0cSHJx1xo6Fw9Q//
iMZz90Ephu/DYfQw/3Ztgl/J8H3l3gFt/lysy7JHuVpfzccFS6ltrcZ9CsW/H9aVgeWoSwKxhXYE
DcK7eo9TS5ccOI/4kVNoS5aN5nh0YB5kkeJ95IiCPP8EwUoHh7FawVvCQiTKg+WsCVURZ+1NS8Ip
xER0Ls1QAD0lP1CjM4kOPxBY3xZIpUZy9TW/angvG4UzkuRUZ29Rs8g1YrcZ2AMor1lqNHqivCP1
spR5tlV0JmMwtP17QxgfgYBbVWeTpS6ygNIUQYWoDAtKs5Ce16M1fQHO/z2jxjiY/cXRCpSx3Cso
wU6PQWpPwoeYk409HtVvBP5aD7HdH4DIoNZ9RuK4QePaf/LSf5RX+aakyB4PUb5PrkeQbvlaSZ5I
7yr422DBFftuNBkIz13JeIhIT7iQds0VJ79YfHp3giyIov1E9C9Wu96ztMwf72WTEY0HodOThrp4
RCQtLYhmDBwkdqdkJ19Ugka+/Ytb3KBY7YammgVl02fwwDlOkZqXQ8t2kKGWgLm+upblWe4wjXXK
e7iF0yqsBDepdj7XvcWWinHOXa4c6q866/LG73p/Q92wK+1aO2oG8xhIFnmlvCFWJLFB+0ao8I5k
3k0rxKeSbxhyydfMlqZP1TLAV01KWhYP0wimxVOxADz7HqZJ9/mK+kBWkjDrTbQqM6HaZ6aofAJz
k+i2BnVLepCE5R4V9j/IPjppDv8Y4+SVs4ky9H3+tJhAgZcTGgHQuv2KC55xxiptq9aXQ7ubdruq
t8667RUxt247rxRpe8MuMRR+ANtngrh5UEXL0WZxIRHnK8/mz9K+jQAiQAXaZqTZhs75KYjNpJR3
xK9VCkIqbhGnPV2VXLxMyrorzOYvKRvoIP4bxghxofELVlqHyWnK3tEWyKzfC9qMfm+iXcujVcv2
zItjxvqeoS2c0c5SaTssG8HBjYGzMW7mp9D9nfjRrQSjW7fSvnt43PEGeY45ofZ0BKLVbVh7K23p
sgX6RMbDI3Z0NcVJDOfixlmoyeVdEbiojswkx6s06kb0nATDWjfrh7l+9B/U/B+7u7GYmrxmTqQB
m2adK/pvmuJmo6/lOu7i3FxUFd6x0EXSYtUZnyhGGAZbIfoX6tBgEW2YLoQiVQOgmNYc4itvOdpU
yqMhU/ulcUzWjdcJQeSZMLMmYNCDiKNCGPUC9Dn8DokyT5d93N5q87bC0GshKhDHku21T5dJ6o5N
Xm+DiPe/gqBop5wb5kHaFKZVORDy7eZ6lP2XndyTt97NF//pgw95jVDcIt+kgIoA102nAQ+Q6zwY
TixnvoyxRxQHjo2V3ZNzIzrdW4VW3vqrC3PMIS90gH4l+RE++zkuSmDmk2w6+gBsQv6AnOudEuED
RlN5AgVHyPm9OwsHGnZcffewEoqBRdLn2fP2bv027EU9eog2CwXqurVx/XZXO3K4jUvTNgeyPcGB
Po/6s5Q/lZT56Ej4Wckv6EtqlaJ+mlyZQShHPFQR049Adq1ue8z21E0tlzWHb/9OmN+GA1+4P+8W
hsIPoTHXkYizZ75Dn2Hml+VYWhPnHiTsOU31IvwVFzIFx80BdKn+Uq7PkrSz5VnMn3UBqXcnhJhT
DGgoKVa+uzNmNGR+0Mn65Cxo+QLuD08/FuaMDNDdEVBCOKXHwrCwChomMPluaNR7FjXz6wVf3cOp
/rz5VW9nKiPcZFi6AWjo9YcYQliUfbZjYV/rAvEHwYIrDcjgDy9P1mIsixnXIwYr8X2jKxd39ukK
w9GNnvPe0bRg5jAAepUURpF91jBZe3ixbKnWE8EHyU4BW61LVE0r26X4jtxkc7a2Mswe1eM7yfXV
5CkDoCdFhA+RDivPg4wzTjJBvVgTIe84Udcig3Ax6tC8DZBfy79IeU7gt5cAtIpXVtyySRiPNs/J
0ZGehmhls9kUb+UbqVqWV8PsW24+R8A2PtDmPHVsAKcsa+Rjx7qsLgD/LbM2xJdbvmxG6GaTOJjS
Kka7UDpeoRoGQBa5fk3Y/6do5cSQ0AuPriJzpTPPtjmZMIBKjzkqXWmKKFuyk87NSsU8bdQ2vGEx
HLqMUjAmdO+1B5+0bk2ScLO1Xoj0KfcAOhg5zKWntfrc5CHwniPPvJok5HvldDSGVRF2f/kmTC8/
WtnsdDiBq30hrShdCff/l+MjQT38I+C8/HN/AO0d4wZutYGV65a7gV1hjekOKNj1Epcm6qXboaGn
L/4/5JrJ2qN6DJLyUFQZRQtKl47AgRFpo55XzzkwBoVFVHqYUABu8K9nVti6n3d44+fUMlYE13x9
VvqhAltPrnPZfptm9t3mX1pMgqeVXzs95UJYEQChCzpv0/SIW/vtfmi4WHpHfGZPBC9ubRAecgnD
r4e9x/8nGwNv8QCMS4yqgoJNu/cxF7q0dycQ78vE1PCWCdK43D0QB3nwjC6E9Xj6WKMqZPZTDx/a
p7CAj9FsNiEDhMRIXotiwXDyquRdKaI+c74nbBUkFJTIUBg0YZNM9KXXu1XEBs/5oCPe0MBnUkZq
jzSaupm8OerdF8Jwh98xh6tf9AdyN4N8IhIFJYoNqzyr7cIJqobc/GdbOKwKCZpLh+M2Fk7COC0c
562XJd0QUpMtxfnY9Yi6WFMhpKN8+s7j0h5AhkkDUdWEhFB6sqK4UKlUglm17svgp5XsM2a8vmDK
08+jQ6pNpRLvhWMCEPDsPGQeJJeKv0Gbh49Mz2OiqoyfD1yhIggjz7c7Z7q+ZSxo6Don9ayxe8SE
bN9Vl2qKd4htcIMhwJZnl46+cx65JWps6Ch9xRcuRl5NAs9oi06vjl8G+b6+WO2goh2DPNnFQB3u
Od85HoJh/KVQ7eGzY+1e5jYWV4hJFhI8GJXeza7MfV9LGk7ACHoiQUPLJapMZNqkUFKEn6bSUVf6
qRUY8kw4ZdnR1xgxm4n7nScuse0Snp+qnXd/iSsdLa+JZ0DYPXXrrDuXmnEuawnfypRr9rlQSHYO
NpM6UozugAWG6fskshkj6d6XpZkKIUa6S5uPDLSH0Q29x2IbsK4QQ+w9XKyWMD5pSOqC82rISGPM
ZI0TNdbXNgBDjnJNt3mypE9Vl8gtiDAGzs0nDfDuRxECoalpPli+S3ltsoGgODlHCH3mphZh9stu
rGCQ3UbJ7Mv2tEn+JVwHMqAYGWHQ8OcPEhzKeTPs0q0uaY++jp/UURhvaDN/0n7VwKRmGS6/wkg4
BhKmTj/Ir59d2DqBZcxLSW39kPSKmhp3/AUrVwh/858BqLzb17rK5zjtU/SAt0/g6eK33ZOOPgT1
rjYmDqmKSH+S0Na0SnNYrS27TdP7Oo1L1sAXZ5P7eRULbm1oKHV7CJ0mXlQtg9obXwlTJjLpLQw2
k3gGO+hgPdas5iVu7bFTNAU61QaeTrOlfTZhtX5FBmEsr27ULD9oJ4iP5/qJ8F82sjk8oS9H2cI6
n65o8V4LUTJ2EG+TzRl/Ps/XGil/saZIAE4TQDzV8Gjmy2tJFV1i+pgPTjW30g8GtQofiYA+I0o0
+zgYHBa9tmpraWvYyvZdtodkXMnENtWsZwcenFOgD+p0Xo7UxmtcsA+JGgpIQ19YCahrZx3Ixc6l
Dxx5fzKTELL8qu0jLxbihQTCyS6/vv7JEiu4DYt+9kBRorbul2/bgzqmbDutdM3QdYe3Hz94tiGF
hDIoE+2ajiNxsQj9uosHp3g1trSEcijszmTHe7m4Yq+diP0VQdcFf3g6kNlrExLcEz0ZlzaaudLr
OieEkWtW2cCMCeY7A44+dwQLnPIm/H/IqSXUG83eG6mZr8VA71ZXmcjMvX4Y6hYwdn43vc2zT5E4
/wpPdVZUXEuPdbR1Wxjyr0GbuiL2jQZiJz2G8ze4JfuWczFDtr4sh8orJA7G/0JOjHS2XpRnM1Dn
h4dE4er6U0yciVKzzcCOcZTHVQ57nzYhFM4ZO9eHeNZMFIfBA1n7AmndWgr+4757d7Wzs0PS/nKK
3QrgYvCDSsKj4/3caz1qzzQYU3VDUIYYAU8OrCXb4QjQ1UlSXfcYCYVu3k4p2EOsxa4gunFqVtH0
OX2I/txn3SY9o1pqKdToAh1Cg8Idlzo4aWUeKjNN1x40Ju058hAcc6oI69Firv6aCtq9EcSWDi2E
Twb7fo1irZez9GdeGNIsyeI6DeS5xdIUFP3SeaLUb+Pv+eybPwhJpqxJi120gcIW0ZZQlUbv2OPM
FYmIdafEBIo19KZ/79lww/eICQ3LliVqx7kvvpDl2Xg9hUbpydY7QcgNAUW7r2vr0j+qa6q87oFh
IjzybNqmtcpmPuG4noZmwv8sVWJR8AD5HqxaDbXxDgd8OYFeOsYRYhb2mQTzdXcLsdkQzBXRuBYX
MeU2DcZjBbD5ZqFkbSRtbR4JMtXwCbFhvqiJxA5/jQxAL3AO2zhnEUCHvbHxZ1HY5JdPDCesAntZ
cfXkvc8pTuCS5xzhLLe8dzDs7hhBLPJtvaKEnMgflujIgwFFruGMf3XsjdambbYNcnQtSr75cUVB
JtcLDdKB9DZz/o5xQuUzeOAkGtNzz7qPJfRi34S5uFQHIX6dMenDxpi4R7pslGWIFPO6h04ngDS9
/eX0k6RmF3DrS/EaGrkqB2wIDnK0nu5b64lfd4knV7y9TbK3OC7hll+cxYlSseTN5iWS2CDrSvrX
W1xN0UC8ccnot3v10+kS9e30VDj9W+GNcEHejoZtqnYKQJlBeaeS7biu/2wn2gOiaA4i+GUL4jIk
Lr4ylGZDSKRdXA+RxpajdDkEAsW8QNq8VKN66F0p+kBZXZJwo4NPHw5ALy4wt2VoJWpUaan0Y511
4g7g2uQDDHM1p8S1vn3miFin6UDfmfrK9iSniEpx0qxaZHjbbywevZsot2VSDtJoBbrUW/VAPuKO
y+jp3ql1BLqqR12I4aEzVfZjzlaOlYkNcxYEnhShbquSiQ10nj+4G9aED4nW2VNbTcLtYD4+2wHN
+U5/gbATjeWf8boyfKBN/20iqC+5p77XKcFIe8MZVOGA6RvEbjst/0gQNQaRfjgmgAEvYO7AZsVJ
au9BTxTXWixzoQ29TZB2E/HclolGOswRtuv9omFMwPf2pbd+BS0knaVjmhhrauLYFE9Ur8z/WzQi
H2uIHTvDDD+REkp0nhV3pqVYfaADFsTsx+ym5DQfb9iuyI1AbHo8kliYyruM+9Uoh+ANLTEFYEuW
ILfaNb0Njfy2t/mz45XnTIYdDhROF8lv60gzZmJoi6pN/QWG0EKznAjqLJ6Pnydd9iFcdaPasxo9
K85j/faFUzaIV2sYcy17KxSK7hiB1TFYZRXBUedkMotAUVkEeKg301kLAiAC0w38Wmnu6XSXx1ga
61Wt6elWPq5tJ50XPpQqQiYgMTtWb8ipVmdLswMYJqWGw8dFLBJKnXa6w6/t9QZ0tJ2iWrlq1z4H
YT6IGvQGWFZaEU6p5Nl8POp+gM145Jg8c4sjzXYFA5qFCNCuToRo4HCMiRHx8M/NzVUNG/1gdkX2
H/pGKYxuzObyu0+uEUtfNu5U3o4zmTgGcRTBIE+Yw1bewvN4p6nvFItTF65KP6Xqf0rb1OWdh5NE
dJqJGkPR4Ajh2jRW9NuZuCoo+0lve+FaXiTzLzjSH4Cua0ErhMtTjxoxgrLBkuycGdDkioJk6yvd
ldp5/Wwf9ziGV4wlpKnXjnb7D6mw3Yy3V05+o3v0TN5d2muG9ldkTHG8hJAw7SRCXQN6ircGn0e0
fggWiGeKNLYFtwX+jT/TUFQqIcTFeIWKZdBh6xDomW2Q7kphDjiLTuh54fLfD75T7jpym4etJEr4
ryQSwcESGUlJ30xXtTgvxpMKSyHlkqCnbadIa4jMGqO6E7x0thITrnV/Zs2GweCEv0HbTlwDRQBV
vrMRH5V7/WT7rNl/Y+yIPgawvufMPYObLgXo8U/T+qJzzgW8560RP/ctPFmTkDtP4CsppRxTzYBV
HYprEqMXTeDuofbQWXXCnSj6fsF2l61bcaqqXzsQjIzH02awUMy+MoR7S9a+zjTwdsylKiFBaT/E
ce6/Oc5PTLMvare98GOQsEC3oKxmvO8lFWOwPDloJXHFyP0MIpKJLl+WqUEiuX4atMoR3ggipzz0
wc4iPokQ0WsiDgbuF2H03Km8+piOCtWDEp1Fzk/GvbbHmMNMmht3h1/8CAL9ASRtAf+e1vtpm4U/
eTR22HmnT6ZR9N1l9mQ4SYUaxNIp1Rl2hTI1xLwDS4LytbSPDXubFqKBa1iZoj42oYbe7TTtoqWF
awIrZUsYoR3rR7/igeLUbeC/omTsE6uP0gD/jL3Ul+kD8YLJUJGksEje4PF9VuXPx+lMZCLLsTvE
VjzYR9NIKexYt1Kp6wW5nWdX0d0QOdN1E21A4H+iVf4epwi6n02SEus+Gv8dUFKSP7b2Vgj7bCFf
kyGD/sIxu0NDiWbrk95RWPCPBFptcdvqghHmp+k0eU0iamGpiCkM1Z81Kqnx+YM4eYR8FgXmvkPS
5JukppZ7+xOHa+wyTlOUQPDm5snQZU9XHgOyjVg0PzfLgA8DmiBiXUrhWZnVIMwfd1qfmHolcQoR
OZJkJjz9EB/3h6GsKRZfZuGyNW2ebsqzv4RZa0nbX6J2gtUsxxV38cEiQdyrHry/ANF7bf1CN0CB
XT7H4j+e+BHnS+kS1vRQpatMWzsQSkipwI4HRZ33Oyjlk67BZjvQtjPQZu7sIf6g46B28RhvHO5N
tHmbEkb7NhCvxBJpCaEYBYdGX81tKpWTEUD6gpyRXnvV7mvrSI7NIIG2lWhi2JEQr+Hv4WUG7lbj
iF/eAD3caHaQ6nBOrXYGRciJ6GXEXYWUV+QHelZ6nc0HZXHBoBFIpqp9E8Y0LnMCS5xJatpO8EEf
HK0PG5en1hAOvkCWOdqHhrLzi9QUsWvt1ZxWj9DPNA9nDUC9RsEdsPJPvrMHgb+v/Z0Ni3HRNE7t
YW0E/tdGjBsKQJNtmHqs6vxUrgUag/LaAb8HfGRORRBYAXN1ikaHXpYAfhnPLotnGMRWjOoTaUR7
ivLP9i7FdNRXq+T3HExAgWWlTlPSZ0cNssIHa0xaPPsuKrA3oXtdx2wz2T4Zrib+v7VwsvFcNtmo
xsk7/iHEPb2Uk+B/+OgrVJCjAKzH1GnNgqYcdf0BSR7rnGiWnOxqRKVaNSyRf0jiNbj+I8QT7G7C
teTIzmqjuX9GibjSke0KW/q4oAzhb0ka+4+3FY6JaEMSZc+Dca4JJoYMQX+xaO2mSB23yBe1plv/
QebEn2KLWYxiG2inbmu8umWPd9VvdFYMNpxMBjO0JiukNSdGWIRzl/WXcFIMJC0hXZA2sCF8Zaqb
6/vZ2tpNJ4FmFIVqPJmE/pOXwAV0LZvMgcqYQEVGvSVRdLYS6ksDYi1wks8ugoZAKVf89X/PC6Pa
kivxKONUEDZS+5ZYGz7owA9o5VlAr8BXfWz1ygWPIFClUHqM24qljY43sebKnFp5ZwLp3mOos5Rj
7Qr7p8CaYw0oeDInvVZTgoYYDo4QficZXo2DlU4ZqaQDckzo6aNG+nNAY5rNtu6ZOcY1ZyqsHKhx
O1/voUGY1np82VpfLKCQq3RwxOjyZj8HopoCTVT0jZyVzajJ1dqWKsNwbkMPblrNMuXq+YRf3Su+
kFIWVh20iqcKGluZTkMCjdk+awVM+8TTzqkkNxVbX6ZvQXHEYDxxa2vDHWtnpWqE8lCdOvkgrWBd
2p+dQiSUTKfMzwHjLMzkw6AKfXsVUEMavs/pPBNSMtXd5QcHnGFb4FTCBT06ny8Xf8ks9I2Mdmtf
uejm8ZEcYY8OWJkNXqPBGcyu993qZMo292QjOtXiUOMHAbd68RR1SZPzLeSu3ThO5/VlJvcUViSe
kBClSVhef/VxHMLcVRpnqvHkStWrQ2B0I7A4Pk0lS+AOGaWhujQpBkjd77vmVilkw138FGDhE3tk
r9pkbFyi80hnoNh5Qd7slXxau0ZS41mhxT7qdyaye4PAchPSCKI66n+UBRyt7H0fOACZPPclC19G
8a7ljmlFsx/K2Wb9M2c+t6DrFcTNuBspcog6XCtKiOahK+kMX1a/1HfBaQ8p1USGUVgCKHaUq/ho
QK3/3ij+H28SzFaFqzYhL9sXgcK5iibRDsYw/GuMnDnNv5Gg61pf4SfeROAyAyAIbwcrGJIhZlBS
z8oPZqOuUA1W4CNN9FDqESSQCPEE/0fHk3MYx9nce3ZKGa5OhMnaqJcEXnvtb+kz6UcdpkyTrxkj
hTU0Q4jAVsbTt8RXY377p15TG4BrHofeDZx3XpSeyUdzl9ILyxpPKkn26Iibpo6xzb1e2rQfwi7u
lSRl2LHptqCfucYKstE8bL3a6rzBoFnA/OOz7ZvfSgZhDADCzAWmF8P8rcL7L88bakMFH+c3Lam/
Jra25pCB+t2JUrgvz8bC+C1djpSqhSaUpGCvrjRsTmzrbxhtuP87MvPlfSUgtHYnZNAP0EmEyIzw
Bl245RwyhqVMOUbjxqkDJGIyRQJhKGsH9f7Ov1D3AnGXhCZUysOUVceRHssiU/xFzFGBgc1PeCmp
kefgWARVN/Dtf8yL2zphVl3Lrwm1pRaAdhIQV0intZ9gBkvTwfxhu12UgEdqA0DwhXCbz4a2CG/5
6hTuQwWAH9zxyUg0jYyOgT3HDK6WazzvtpFulypjbIX+ZFrU/DIGFdNbmjFLuTR0v0Ne2HM7rkqX
D95n38mbudZOop5UIgD+9KZrNg6hQH7C9tEEBY4pvnEcXSfbexPZksYV+N/AZZw8zVaujCmGhOUq
dr5zRXvG3iLHbZcfgHqoLspUaL+anN8gwMvCP7x1E8x4kOKFO6x9V6Ue+QdGhGRlrcmg5Y5kmFCv
dToBZBK/SyCEWjy9z6kQ0r9ClwweAETLLv61ux+U3S63vXvzA000InJ1jC7K3JVPeoKb7SR//wpW
WG1RcrMYDoqXnh3/PDAszGyGE8XGZJQ/CPLpt0vm+JqlER3TNqKrViUQEP64nnMjNqOMwHeTOXc3
S1bPkOmpFU7mrxBpbJSo5FP0kJ0SeFDJjyguh026QKaVL3mMyfHViq1FYZUlsdqU2qvdHdO4W5Qy
uUZGXRnOhWni4qG4yKoXaiYDsrjMIfoyuNRIEOVHJbv+an6Ryz4UUtp6BeaXlcZIkAPqc/2y78eI
dZxXP7nu2LSfsNIKDoSo0q76gdKwKXKvgsm79M+XitlQLgz4hQ1SiJU3IBHhW0AlWHY7c8hlCqPW
4VhSm8lHdX74yl45OhNEqBFZ83xZlsBSYjnguK4JFgRsZYT9DE/BlqJNwe5t9USJ0cm+YpOVjkgZ
3njK4PsDF6U8RAZJ2nh8OVpiVI7dVJoP+8tUBo4NNzjPurMD9l8LSMVcCJq3bVl326UqSwunqFJG
4hiWl8T24OOt/x5pqzVzXVR/vP9uUXYe72sSUNKwhn0KYdkS3bqU6m6hZRMDW9D2gfWmj8yIffIA
h3oEvC7kvBmEBsGd9UvrUrEWh1t88O+wngDMtGdz4k2Uumb9FZuOQ6QHZ45YpgTOuacftsrBFYrX
DhiQzmpOaL945IoWyF3/fSY9L7m+Mc5cRt4lvqoShKCLjGnv4HKRBMM2PaNtUPnkrRstTrIKLB5O
D8TLZuZEj4Zc0wdx7PeOsdQ6tJr8/WA6kExzqCc9JM+SesMg/PptfY3yxS5wo6MCUMaHXB8DHpZs
a8lhY6A/5dDm07yoAGje+JPeSf2NlivDdVkx/ZZ03Xmbi/kbnbIJxka4MY4xLOCfIMirdHFq70Cz
ZRCf4ayiKaD1FbgI3jDqEdLGbeX7lgqbZfXSWAVqWeAOGLLbyl0gtZi3zCU8gXkSpeG8wXb70dwz
GCGqHWwCvAvIPMQj8SVLvjbNawkFlf0Rht3GzC5kmjEmwe/U9LoWqDKQ40DE66aeZH6pnzDC7/Ef
plxg4j6XX8d+CN72/+0tYnnV7MoyqH18+vw407kxhyXxMxvtDHt+WERP3m7afccARDLFqFcQIgXo
/zjL4hiOVVYY4oSFuncF6hpIKLgA5lqF1BOrCwAabIhqlYowccL31Q0ME604LXv920O+nFzB9WgP
Unkvq88KWRWdWPjYywNlUo0PoPMe85NID6mn3/+opKaJUEIQ9MGyjPresKKs6rzInp4g+w67iqFJ
Y3+W7xoKsXSZhATVm4h42g7zuf/ypOsPvlF2YCfXaBCdNe4Vzylzli55VUjLRxifUC/dfZtfJAnw
aqU4RcbFUjoJKQsOwe3yTD7YJqoyJjlABkIvkeMntP8sDKHRLZJ8Waa5dMtInKgQhutpE3LFU95L
CfkLEvaImB3DcQikWO4099M3iQ7a+SSO0lLO4AIBcaMuE7FjtGRD7WXg8pA7bRmjp/SElMfpJVVO
VHAKuwBqQPd5jvHN5FnD8ItfgjexUXW8+KEuvRcztaTu5sscFte4o4bubZR9+W9yIdAbM+N4SJK6
+P8lUwW6zw8/0a7MK4gRvwHEr4YI9VI19cbu7V84PGVB6cxPcCqcssol3bl9uzjcwmIKJ4S7u0dt
7fOeqcjS9ytFB2qB39JeSpAtUKJDrSV0KuG8/3S5rT38VHB5b8Ab/6N5X+r7hR3Dvu18MvE3EEWn
61TAPM1an0nV8XCHyMuIRGVPG3JXXBvhAUUTGSn9OwWWdBO4rSv43Latyu0++AEm7bmPzW1A2+7V
RS3P4OAguxr8FKlvTDrNsDyP1iRIdgvZJti3iRB40GEiOGcQ6s2vjY3KZJPyn0QLJQgGwG9OenmF
AC8t8wt+7XfZyDvwhKkhm7zLqNl5/OiQTigT/CYz1vDC/l5Sde8BdM1jWq3UGSpFE2bXSVE1wZMj
NU9rh6t/CUnkjCQzYLc4rC/RwIgWK1j6coMpzxXFV7sdPFHFwtQlkx9tjt/TkvcbL/MaEhYr+MoM
Txc2vOyhj5Hl4FewcPjEGaPaullb6Qm45U8MOREq5PMkIrdQHdMg7KkrT5h+kBGugMMweT9f4uAr
x60HSR2m4e8/K3nnFqiRBxs7I7iCwYfgLQzt4mqexar9Q1t+zF3MOuodGz9spebsavL5N++TxFJZ
91JRPbiHc/sLOxh9I7CHEUK6JGo2TQ5I74K34f5sVXZ6DAH57Y4f6Clhpl3rHX111/E0T6s/69PT
Uf1qa6V/FRoZTx68XHLBtlEZs+tISRzYuyVLAU37R+nOImsL2LYUgmIwvvPQCtVH2rKcCxpLqrco
dgyhz4QHb169ryyVDXz4pDxlxQQQc229+X1+DyZs79hFnYe03lTeqC2n+nhY0e8vkpnaJC/qB2uG
daK6LKhuXXPb6SOK1kPCo9VuFCXDD00alWfSDgNyvvNrYhFMxqsvqtXHnZXoprLIvnoSmDOwOVYn
oBqRkEQrDKd08Fd1Yi90zOEQroYqCqndBmemBxzdD2F9JDaU6D/nK1CWlWtbJ1yFg16YZ2wNoHXP
3ck0teZ9Fd1snTHX905NCn05Z8T2HknLmWAD3ixKLeCm7Dgec2Sat7vkL8yo6w514Hs6TQs8c5b7
itQyGcK5Jxrga2xv8rsuxDeGPh76EA4MGFM2yzZtENasE2LbiZVM0Zn2jZBCSckuY4lHQ3exu6ZZ
7Z0QXOC6IikeprnO7neaX949kFrQyah24aF7yytytpCwBxBHOljgiIl+dWVd/hB4/h3h71ftEHiY
HuEeSYGlykL95SUkesTbg2uUu2fOGS58Ttj4k4jCGYvVf8AhhCocLo1rizTAaEkDNPOjjbjkQFS7
kSNa+GChpoxYmPymk16hDnKSFTi6Sheprll1/ciSiHyC9Nl09uF+w8sEaslYtaLJjnkd5EJheLrY
WhDx76ytScy5ORK4iqoUCvpQmtOFjSYCPtZ2gONZSHmVtQGIFLG7JOFFJ/g16+arkXpUkFxi+0S3
xS9QW4LnKiOBDLP/IixQvnUsGG39w9yCJtMdhHzEOhuGmGKRrZs5sKXMFOEKjSKpfeOV7QkbIwNE
yc6XusgufATUdHhoXEf6DZZ6v6bsE02XacpeIuctObhIWema1nV+cdI62a8ZIXGsYO9ybeR+nYXR
faLHPLlaVZ1fTStq7bYwoeo3uDxDc3RHJn8HWfQ7jss30DQTSqUOK3xZhCdHPdLFwyd1YUNSoS8z
wD8hGn6yjT1qVeBAL3RjgaGmRx3b254B2lfiryBrbb3Dc7v5+claFUYR0gjxK1B3+jZ1wagjtb8S
dyg5LTs5fbqFkU8DAqBLzm3OY7yf9C11PBElnBNjDoL6yKdnl8Bdp/Q+OlPCmxbvhZNxsX2/IdPI
hnPIbj2BPIWcKI76d0No1KO8+bMkXqLqPAvqna7HTLHQwRf0PS3SJRr7P+Ai0iIGBpfgMu7Hi4Ik
nEJx33aWorv9eY7U+R5UG/XXLAzDqW3c8Dtn3OjtUjgqw2SLVF05bq4trFblLoVKgmxyfooI9Oqe
kU85fztB3quWPn6Zew9FRvckjzAhxRXwbSr4vl/ly3kinLgS70imwZGnyLBKQ1OwojjVfPNseMFj
pjMUrEkLkelCHKlsVhG1h2KZM8v2hEf4fdshlNT/gSzKfTPpdKA879tNL1Aqf6MfV6r+dJ25UjkH
9d9aRPqwAZWEhQefRa6Df85nie/+R+WjvsjoFzwei7dCPEnKi/S/Nib/L6NFn2bTDmySnhElTyKt
jRLWCZcRvIR5kFVldBuAFlWWzj8Vpp6hnFTi7cRpkWlTDZLCoPb2ECPefMqWD8nPQ95cD5W7oQHq
qubFBVNRAd2SW2wAmSn7kuxxt8/PqScl4HcaVGGUp+AfqaxTq1zc2vol7gxkzMCMmaeLqOAE9bkI
yQRmzaS9VBTgoCgSY68sn+DW/kZc20xF9qAJuvLfLZF6QE2vRZdFHepSPWW7wd+G1YxSaZ3A4XyI
Zj0tNE+2bFJZp7Dr9Aw7Oxs7WHQ+WgJ1oKMkbocrgNwDwbNp2xQvKToAK9Sufu41I/HzMxcvmpNX
x+w2D1EX37K8Sh0bit7AJoOpJovGQr3KQ6Cg9Sqt8KuDFEviQd4dPw8AdszLFv474TOPHJzbOxeW
TmOUreXWrPjVuuSzSbPrJ0m/B+IGCLxb3YJ3z45HRoX68qNOez+X0z+hKC69Kv6o8ipZ7mInQQ1r
E0pWPbI5UkMo86lI0ds+DGC/4oPsUfbIoBg1vYxeKUkVaKPL7F8/ArUzWqjXVX9hLWnI4SobAfZG
82lxJhz435jVzAIsmfzJMaZtJNwv4wknZnFRH8FqHJaV3RxB/t7xVCKI39yDlgRa2naGOWbX1WE1
VX98cCbYcuSqkvxARkIvcn7tYAhmHq0uwRigC7I2ZFS63LwKxjmrRB+toek8x7IsqCv7qZGHFLao
ubc5C4pcE0a28djPDfU+NmVYhfYqiGcJ3Lnrq74Wcra+6b4xf6VWbJuqZRP+9RNbr/4I043XQ8mh
79cr60spPU50Q3k55DUgeXyixV/JI7Z/NfyI4vpvRf/wM4DozZlHKZX+12WJq/sQEOChLslSba0X
2HfAQVF5yDJWI1y1lSKj0h9Iu6HfHO0VUkF5Y0BHdqRiJ8Wu0e8cZ3IahDORuLknZdMl+ZWnvXZB
CplBJO+LqnIjrMbqRb18Ve4AUr5j+a1w5wAD4q1UGl4VF5sfrJgzSMu4SA0EKFd0w+5jcb0VhPal
H4V9F3P9wtZVU/J+YEwM+kIf1OX5vRBNiVXg9gmq2evIcpofiYhZKHW+FL7jax4qFEj6oFkwZJP4
46fCkDM16RhJU69QsETICubo7jNjESqiRqw/Dieg/unHiyTtGPvQ9C2iPj0c8aOsq7kf9DyM44yF
v+vOR9dK5mI4pNSUNjW5GycweFcx6SFer4GL+2Tqj+qfe+YS5fOfWI+xU9SMIuDTIeO9jNCKh/eq
jCniipbOmf3ufAuThosYhbmZVZyETc5Gta3leYN9cRZon4rAg8RsLS11I+/OgHe5wXtxkNNkafF8
hVPMPq9GCXTbgEbCK5NWUGkm+yo9K70ixAWssLYCrg9eU8v6Xhqtrz6Us75X+NSTmQbfSP7tBZDm
5tNkpc9u9qbDokgLoccKY5P59U5nEKPzB3wYqqBWOAzIGNnwxZ3chHcv0FueM/7Ha9sbyYp4blMr
fF4mZZLOm/Ottr7IKJ1SS0nlnNkQRBgrawbc7bXysokZ1kaFEQRbyepTFUjmv9ALdm3PTiOUohUP
SN4JJARcM0vU34jEfd8QrVOiLmkUgmNVPXWoNdh/hsJrNvZXrziBK0kTGMpT5CiiGvg2NNYzA9Wz
MgDEuBrqMt34lwIQ6n4oNSqpvGvAsO3G5WECjJciFuJBiRjPuD8TAHkfhR688ZyQJFkXc6cvc7YV
Gpxu6/Ru5vgktBIZ0rAQlhyxevufUWybZsL1UK9UKOi4JfBiNF3mBuGkM87uW0rb9Tprf3t8ZJbB
g3Ak6PqcB/VN+/Bp16YZKNY4FLHHM18HXSoI8flurAENxXj3ZUqSe6DEV0egFaBddgOkE8cmmg8b
bVsQkcZbqD24/emE25cSKSowVG8+9v/iL5nBGXhbSN6RPmrdiKzkatarTWzMosx9HzEGbbc+x2HT
H9lSNIYnPsFsQP4cPP6DdwQ5y9mo1RCEVMG4AWltZ3tqSNiRd0DLdRPGDLAgpQN+aE8c1hhtunhm
P3b6vzX+LJjzeo8/JT6MQM15a+p+TLAJJYr+BzAvPojfCRFSiYstR6V9aPyj7BENSIxM98LBh5Ok
q2htvGutMhjue+F7OmtNNx7i0uME8jGpk4MAJHm5KOt4kx7b+vjDfE90HsKFnRrb8p0PQFCMyZ6o
zDkD5d8YNlLQ5B7qsMacsnSVfe3oGNN++DEJ0QmapWxafbBFS3eEku4OxE19+qCqWTdOy7VXgQXz
/tBU0an58kbhzsgxoKr1MwKg/VKTYbaeQmNMc7x6D0gofuMqGy3uKk9kfwg8v5yC2q6NMsacTqDC
FRHTuYnx5aIroU21sendlyANHPYj8+aOAI0WRxO81C/MF8NLgxzv8to6/thYy6UesO506dlvYwFp
1MFdxb8Q5yrbao+2qbn9LlYUbqXHi/wIOunCvJJtvZ0cIlRVjfCyRIgakUEXTbIyFb+7rdMWBg1D
/zY20bcxaoyBWaLDiwzP2d2Dawx+yertiQGfVnWpuETFXufbHoahX4YxPxmQ6Kcq5+Q1WeOWqQO9
EJGFrIseluuC+njxXYGUCWLMP1qmq5gfjYRP4S+YzjBQkCx+X7L4VCnzpw90/Rxhc1VkiOkFlLPP
zley6Dorl5eDtTnVd/t1ETI/L4g9/KEaxNfY15xkx9gzoHNM42XD0wMRbAxEpsqKFUQuBoJL58rT
12D5KlUOamiAK5c1dK6ZGFZPawXy4c4pRni+OjF5cZy4Cd8fXmppKAbgfi4pozi96vX7Tn/QMMeQ
/rHIpa6FZIWyObf/OiCnwPWEt8syhriikeSZFdFEAFPUzY32mJTRdTO5VxvBx9GsnMZyHNghVKop
K1g2k4heeq86lJHsb1jRR0HeSxiUFtK1dnx7yHJ0CXcuuI0bNXF5eG0MmK3xYNKeMdTk0t0aZJRy
OlUz7NK+nxcbXvqmpxM4EtQDWJZ+HukI5Mdv+3MVdl4ylAC1xB19UVG9kO9VxCyiHXEDOeSQ7oI8
s9d1LUPJjlAn6tQnc6Dpp5/YCLHHBcdTX9gfY9Iv2jlMCGBkQH79l2frV2p3RXrD66VJA20nbev1
aNDO7bsPDiJc1DNzw9BRyg2vhYPG4+3zdwRxVuGH69LgtOW4AthSTgx475O//1Hc5eDgzun8PoSw
9B1MnyJLVzNmzdmPI71Frh07sK3NWmAFS+r33jNvTVePQ8d/3NxaAjkugOJlsQPAxr6uJfvTC9kT
IpIzZuc6RHLmTaOf+GC7/zv1T35xCpBYvSxm5Cq5F7NQ6Joz0hCqlxQ1q8dyeTgIAZx7vqO4HjDs
T97qFEBuoZGDkuiOP4D1IiJccnje6AfNfN8XEPAyP8InHtMNygz1QnjLOhN2FW3OTCcjZUrzhUV+
QrloOzNqGmzvjiB+6TmObSzh663j+lu1zVUCclM4GiGFWcMUyiqGzUIIhmw5dyWIWt+jgyM5Av0Q
36iueseGwhj4PW8fIYMzP4OMStym6kIOWfxZWtp4xDHB4iD+CqCbvRXCRNcrO8HdY0YZP1CYRrVB
n+4BaSQ+Vyqac3UX5Y2rmBBUp9DsEVaqR4po1uH9+qInrZBcwO+M4c4006a5xYsqjunmuDsx+raM
evIWxC+0dV5GZ5EWl8/2SYaHU/24nhv26yEnaygr7zxaM/mG6tvSCzVE3TXk/btZ3/7PxtbMK69T
pfSQM19WyRqnR16tn9uJGDrpsWAJjtaKcBMryfqk1BtWaLAcFwv9Sosco5QHmgY+1s9CoPAbR9fb
8eyATn3ql2tohITAB/mbFtEP9b1iybpmcvxSVO5P2vEbhoVsVivDIO9moF5u/oK6H1JsP0vgyHmu
Kg+MCXRLwT/GYV0nvH5zevChBbWObMNguvYsT569P/Xg3TPs1nkc6AfuBNjsGKpLgwSzOCGy3Zu6
CdJVZRiX6DQsOk8zcIK8AsNDUJgLmjA3F/SScbiwDXlZSGdk+8Aj6kfwmefh8+SUqzAGjw5qWgNy
nx1XJT0yH/ytIMoUqHy0Ao/dfxTjCu1W1/oqWvevud3+d9sQDRiCB/XNxwWrQVzRxW11AVPdzeDM
XJ7ejE0lI/eksdt1xAGhDP6HtnWC323/pF4V3gO0S0jk7OZSmjsK2G0RGgCB1/nX++IrOJh6ZX5G
pHFZ/m7016a0MZ8tmjNUAg1xPOWX+F59Y2gugPfm5TKMdH3Ba14b9aC+BwLUu9cP3JM7k+RY/9v7
MrqZXjqguSQqS2PM57AaYtV/+HlaHhR0dTI4jHw81sTvPrH3LvaZsGechbR15Gf8xNV7nfz7Rj2L
f9Zkd/xLChJPC5l8HY31XrFkSQVs8j+yMUfy5JD93JnEHvj2DR+/SrQM2W2Qvri+IiYASq++K3vr
hlJHcFg65aUnD5cA7pp6+CK1wowMf0E2HMq2h+HJ06NGzN/6YuBqBwqaOeBwD0WV2Btw6k8WZEyo
HWK5FgRKo1ybsPHGlZlneZtv7KzVnsOHIq1t7e7w+oWEkl0ILs4hM6fPqIyIhX8mtbV8sGMaAXP9
/5x8D5cb2BmWPfh15wnLoWEuNf9WAdSD3I+U4mahe2w+zK8CPzQmfmPnXHgXitMQdwOYS5n/HtoZ
fMTVViTUKUZkR12yQg47OCMwmBhlvgFHtwXv7XXkToVV4UE32A3fgBF72POpg0bNME9GLZLmdTUm
r3bM4YRga7lRAcGrslwkfEwRsdSJNH101e/h0g1wAhL/IhRLg2nCYEi5nqY6TuJeQdJ3tqfoonPM
lmc25c306xCpfsiDFkNGkYufxlextsOc7mInYITywk/fBFTuB3zdXhgg8K4+q12aP+1C72JrpFK9
GQjB7ykCNkMu30BnnCXme6wsmOZi/qYdc1/Vcz/2TmDprxRuLP1fs++ahKU+J4W5XAr7So1BzN2H
W55eCvMbOfEaVXGZP9Fh56BXOQdmpAM8GAH6opXp6VQwMvvSxpbq9wvHg7bKW9/BLRviL38LkHMF
UY7x9aAD/9OZOzByUc3FD5p7vjeY2d5ZaGHfE5N+LKcHTTLG08IsImxzzM0446c/83iWuDPU27d+
HzS2rw3QJ/mrxXQLvs3FeCtrUuzdoQ1e1aZ9QWI4x9DcZFEDYY9RUFqybtXwh1e6Z48bWnW8Xzro
d91CDUoAEVCziW9GTXNUs4EoLBs2GHWWH6M7B8y4uBEAhPUhKQuFdRXi9sa7hDVFGMdbIgu7bA/b
cfLvnUZ2J/Kqsrn0JSNuEpEhsnkaCwjd0eFM7pmCcGl3qYQk2QXX9lzGmQPma8DAXTE2JnO9n8pf
3jylYn4kbtErAWh9PBAnPkld55cyzJywO9Z1CHnOEtQhnnOzf0yOVmSmtvcq9h/FvSESpLv1ee9V
AivMXexwe+2hTf78BsCqa1ulYqBgBdrqQr/eK0OcwMtT+V/Tyi6PqrqB418dy3qsWdE+xLYg5OLr
PWchwxInXjN1tYrxjWtfhSRVs/2WvFV+5FwSSKtiwARQ9qznDQZLGNWceGW46yteXEyY1XCQxPC+
3Kb3D3FBMIYxROAZ480FN0guedjAHkarMa0iWLvCJy2x2PoPGMwpY9Klrv/ICzoLrPv+jTNNdinu
9aa5Al0UGj01nf+iCcDAawGHU6+DNLzNnpQ0O8R9gJixuE36Z0oUojEm0uHLjhEhYlfYbzG8VqPE
TAW1uHezw5I91yyI5mg8e0AQxacwZa99zyADLT4nrLVmaipagsoeKI5yPy6c5dH90T+lUlp1bT8p
LH4hZGCMdICk00U/98qJWnpmaZz7WUIdFHf2ejEgdvJ3swy8koanJSpOfuev5OdvyatkDed4fsX/
327oGCju0E8OrnjZC3lJstlj9VMdTPd22lDIGFN6IAt5/HlFGCxNRi4eyepltMg+7AxDZrOZStmr
3seDOdhp9kqs8gz8kIqsdkZr9msMO30K3c/UHyPZgfhHkZyMZmliGCX0w/S2QLMckT0eWm6CEJji
CpOeKFK0aFLgL/ydJVzrbUsp4P86nDNNJ9+IoiF5xP+y4+nkLre5huSEEohZbXHDCDHCOoTmRmSa
mhKx2ZsPwrZmKV4jpo1x14G3aYYmz5zhIIkSU/wmWzIRhcwsbBir77pba/wLnwcbW7DfbSRUFkT5
6BHP/C+6d6fdJs0pnkUw2qT1mx0Ucvifz4j2Kndk38f0aZSrroewKpm0u4k/Xq2QFZdBO+jOhyHF
9KB2txhyOoBCHZ8Kv9A9+UqJwmJQTT3jsI+Qwz6PL6KKenVYaOnTs02qXirLFI1/ZlEI5OsNPZ8o
7ERKlCDjRbkRZSIDNURJfPpzbKaVMtY4pkQd7tXbm40J7hMXHRQ4diAj/95nz+txslxQ8k19Y6DA
g676V7xOcMWwZTiYhDtXvdETTAQIvXWzPlcU7ULMJkzUK5R8LUPE7s/1Vjyaw6zeHIZvHLHxK0X1
v9fI92KRv3/3MqHxU3M66fR4H3iaLfC0PApsDCwHWbg2xg3Ws6l93cwWL4YrIdCDJZYJp6V4iHfl
MOAwoNHI+u0mH87CrZNQyDUtciPEU7LSNrDncTvQfh18JF/IaczV2OtkCcJs8M5ImAeUXmc+1DRI
3vj22fBA2QYu6hjOlJ5Aprk0dVc4vljbbxRsZjS6mTfh2TCyebpAklLJsjvqYpxSFG//sVbap3hi
eBrJPLWFTiwDsN+vdCUQelY1VkCQ6owPiUN66Cf7Kv5Nxeb0KGLd+XgfyNred6TCWAthWKDFMIhB
U+GCpzh7W+f29ui/g16B6sBsB+6CgLDfynwVwohmtjntxrCam8HTOvMnV9dCYbWc4VpYMZBgjohP
d/MIIMPCoS9dh9HIKQfAEcXgX11e8jv8grONgO+M9X+I6Dbv2WTccS+tWTfJNEp+PLJJsvZCTwmS
JrLI00hQH5AchrZY1Xskn6N0dN5VwcynsZOMgE9lIVb4yfi2SM8T2eT3bCXly7VhVc1QDD/I6Nvk
qObZ2Xsi1QP1/tQi4Jz5EtYe0Ebf1msyNJlvYstVzv+QN6irOIOx0zSOA95XYrxfkPaRKI1DvXys
o0MkK7JPM8E51VrS5Lzhaot+ZwqNP5+cQNuAQ+wHsupiYKGz6GzCuIS04BQdEtJzd5LEPyXYIc7j
J68Apv5FOG44gc9bLDtbI8Z3nMR7lBxOM4LRbqs/WCPf8jGuhZaHT1Wxq560XPFPmHqjuMS64eDX
dg/WeXHRnYgTcs/RmzyI5Wf3Ig/4AdTY6vsm/zVGjQBRvXlzCbTdRO4LGuEO8DWNeipFmXEIoJtf
cCYQ3SO/w044k75Q1nP0Pwe2qH1rPh3T1xUd/1961IDyFrjKb/386HynXMADFQySzos3Ft7dpAop
7tuMtLMygJBKhNBWJ7SuB4d3V22dSTdkDk995t8bF+dLxXRFyXEfSuK2OJVFbRbxupqQ0QojzTE0
WmOhqmh/tBJmWH2M/xNr/QRiQ47zA9C0QKaQx/z3rtnI0QATonsIAxNTpjXg+QzlqecCGGxVmjXw
syl1H4Ta9NbCHR0iVADGZxV7xcoN6bFP/MeBX9nmKMW7ngi6xx8vJXtRdgGs2hBZQffhgm9SIhN2
XN+5VhXpgtpP/61JJXL6HS/STMsObHYUF3ZgWpFOCplh7eNW3oPy/5WND8MEjJryUfJbs/rq9ugv
k9oZJuHSaiFz545SdAga7z92ne45yXgSFVUUUyCI1SMvMxt/Qh7s8+0Qzlz6pZTBUCGJ7uPfYPbc
444gKRs8Di13v5XDvAG98CxjTN3G8OERDTDoA2plroA4Tt7WABHuDuf0FUzgwqbx4kJZO47lzajq
KFznxoR9hevxdSyd3fg/nhawmfxUxO0OBhkZVEUvmEkwP0Od5OUX05McBd6NmiHkrchyY+Q4nd59
D61Nw5HOcFmdTJCOWox1ceEoMjodv+o5g8JvyjN+L2iOYVFhx2RICcfVgt7lv0LDtuhC8o9jjWzC
LMCoB5XS/E6UVBJ3WxWkXdxb91RGzxtYf4QvJhIUlE3cv+pIVtw5fHWvmMwtwJ7Ibh2eLpZqyZRg
qFb0rVpmqJrWLCIUgFMX8pgc5We/HGiBq4fUfO5s3sFDwtiBYy7U/1PVrW82afol5bUBQuz+txLD
9bHmxHdh+WFT13Emd/fiW9Ae6j1LG8BdDxIX37c96gn9Yu/ATjNAh41bmpv9IrnrnlNDD+o/43cQ
FjCwjYg1bUKt4BQpdsbqRDNgwcgCVRBliRvXXhqm4i7/BgcADM3A4EdWCBQlDNDLctG25OQd4Tvz
n82HxSq81GCPK4caU+sgwpj+NyuL/SXJl7GgDxuBjMq+lpY6tbCpkvttK9dBR43epWl9kq6rwGM0
Rewu1D7rSz3Cu9OJy9Tv2or5n7sE5sgDdiwZobjMYSPxlgtK8tREoPz86ONhXDJhcXSjNLVJJUle
Cvv7KFytRtwl7NvwIciOqlHP4Uv+xyMHfFMIKH/IYXZ5ihgY02w1IZCs957dfI5DVQdRVAC0+vKp
Nic0D79dYEm+mlUX5+ietpdbESYGyjjgBy6251fTEOKu6SHST3+0GbvwNuW179cXY7e3XYPcAYm7
wAOBDFXuZqc/QMniKfMEOaaYUX0DwVajMEHWftf4A3v6fkWwILZn96ieqygAiU1/9dFjHVdaUj4n
7OKPZnz3pKczk5d3k/zBcTCZg19oJQyp6wxqoDQ9cVMODYAMwSbOMRKCQWyuzUosPzPnyO+qEvP0
Pspr2BNZPskYK2MP26wu1BO+blo0/0TnDMhp+YHjuL1oeAY8lJYInUYRRskJPxQYzYJ3rgQ3jtdR
BKyuyw3pF++aJO6k30fouc1USb3cs+8Ddw25yOm/6K/O5tKRoQJ9j+wzX+KK/8aavywnxWZ70EHU
zGXQcs75i3XxOlTGX9SRTjZHT7yzmuL54xBgBvNejf8cwvsOUxPyg16UBNl87c3TBWDF2pcy8+zy
JJ3pVlA09AaCTTBuOsz2Zr/Fa4CQEwjKkOiSslgR7jEHnLo9uVEiInpwH3mRN/rAr3pI4d1ARbBf
QOxmcCxpnF0VLVoPs67Mi5ArVWvn4wF83rJEN096Rzfp7mvs5r8KHRS2JpbDCxQO6zA6i+q7voB3
cddSwF87C5zGWjSbCFYF7PmXZ6eTemUAgJ2V3fJmUvnwTXavU3dj7Q4Y4/JWlD7lRCW+p1hMSwYJ
6/yHZJlDfk7bBbltpB6J1HS0cTBDSkwmcRAhZEkEQF2BIGnYhwin2EANPeH8BUSs/X+Oy8ZLPq22
FQmx+SwTacyq9BSn12QO41GmI6qmBDS7PpBP4aBSaGBuyd8iXvwt6KSsIiqeWQetuBdDkjyTrHOD
zk55grT52XFLAcHbt4uvMkK+7c2LGbpo4wX/ClhsyFSodPXO3ZNeXrC0SPVraeajSOacoylCRfDm
jYTrhdlH4sUspwfPKaV1sRm08zOrNEj9lMcCybLRtj4tggIvXoqovUgXz4n+yPn5URag0zK/pdV5
cEtAjUjzPqsoLBGARMkbEOthgV/yFnTKP6eQh0n9WTVbj+Jyla4ykeVQVJj/4YjsKjji3R7GDNo1
nTXLBde7NGTjdUrXdOfj8skIgXZ64wdClqog/lLchT+LHyjLMIPW4ryZ/OqMe/vw3ArhRpY1dkj4
DV7cBSfzcGFQrxamVSEP4bNbq2z4S8+OHpjRHPITlZ90BRKa005XQjEDBX9qyfn1o+F0TYPUqSAa
SuB3o3euY1MZHJJeYzPndrtQqAXRXfcsl7G72OVVXeJxqO1vOQd5TdPD4rEmHicMWzxqtNNte9lh
NBecKoJ+5cuo6rX3nIuymJMZU7tvwa0yUkUtSoHKHvzL/JlWZXQhGTGFYBq6VBRkPxzriJkCIaD+
UDGeqRX8rUd9eXtYIw00jwEaJHqNHzche0/DZl/QSYIVslqEVl+Df8Iv57gy7DgIsT8llFzeM5xO
HTPwqKLiZPx3xC5npcLyJRip0Zdt8RLDdpPaSaERLIB9wo4SJ+g3UPV3+J5zco2XO+48RVnga7Wo
CE4KCbPqosJLEn9QM2hJmnZ8C8FvonGqNMEDJYHF3+KT6YKIIcQNfF9DqNrdPXugdvufovxBCM6z
p7cvsXJqE7Pxzyl+l8Ra7zLHOBoQND7hqdlMVMfO5QnC6Sld1cFouaWGEzEoB+3yyjIYGFRfe/Fd
k1lG6pJQwgi38VpfV5NuicCcSsfjDsitahFtLbX4YuKBlhuOxux03ZaIrjlvrOZCmMvfea4gWIxX
8exHJtMaYY1N2ce07vGsRpJ6CgJLXzKxNCcNx1Tx+oJb7wuqjnMMW6gwOPt/3vUftbrE+N/I8Z58
Ft8q0W02MbBZmNf4ddxGRFiH3ma8+iMGcfK1Zg8FzVU+8vC2cYAgjAOwOMjG5Udl2j9leVSZ6uix
amKceyOrFaAxqtjp/Qy77EdN05NsfTZA8xTYHFcfMvY7oJhLU5RIiy41FH3upuIYDnV1UIbWdxWb
A/n7wLOuK0po6CjQ+JrG03c8J49v7Zw50le9KEMQb52TN9NNXslDw2yL23k6h+SCuONnYWsEp6jz
GHSH7p2HnDri/EC9TuWzcjN+1JOwnHxre0i96UoQgxioURh2khttWFXf+d1riEP4yl9q9YRIXugi
bJ2BawOO3l7Xe7IHQ4EPgQWHrmlkzLMBcvKtQDE+R+BiR+SYbDV4S0VHJ45m6gGEPfFr2MvFgumO
grfca4bxazHmV1V3d9Jjj8HtHIF9ETHXhDdf+wn494yNxWgrhy0bbQoqEI3sVd19Viy0p4eV2NTK
lydv1C+1zsjWACU3Dnvviy9Y4DonEYGTygC73KbgR7uUKtl9oEeCijRRE0dGzw0p54kX3ryitr11
NOMW0q1nlQzx7m3q6dnXyfV5ybcW6jeP4/SaIdtrKP6lMKZMJERVBMsRfPZvvSg+tqplE5tjc9R9
lqxEm3QfdXfmnLKlTHwBzb5adQc7DkWuqa+zteXB5Blw0292C2FE1HcNuECVt+oyphF9eWsQUpYS
3LrNG3/nt0xzzjXAosHWrdOOXUT0SU5ssRVQEbt4sKtaKSX+a250AJU8F6XVxfBMWQ5OZLrsLPEx
/gneyJb9/RZxQxrmtsDXU6ds9OrAM5kOs08h+Wczp5bjZLM577Y5tFbQMyDWLaRfroUZdtdNmX2F
9FdF+oyJq+F3vBqH3bXiBgBLLvqFEw24AZtq7IvFDwwUnRNSbVEEtXM9oZ5pgKBWvHHgQKW3fpyT
lPnzW3/cZt2+3YdjQZh/IY7iyq0jgSLVJBTQ3602bFZmWheN6QYbrD6S5pwly2OHJNEyVo7bwGL3
m7pDIt/T3yIuL9CNj6+B9caK3RBjp0E8DvVhdDDdaMtenNERmJ+DKtI4rF852NBd2Eq7GAnWGAly
ctFji3BhbgsAnnpo19/YcPnPU2DB8livFlG3em7Yv1BR2ZzfZo0VEh4D0Qrfom1LB3MSPYFRVrb7
62i+nzLpAtrMCoPWXImAZlxKp3v48hH6XiySJ4v0GG7p+ogR78LCL0Wo3bcwFFkOQYHPo8BbKPPs
VCK0WOmfuUWYWOIbmzfe9SCQ8C9rwBKQT6rKy0dC+myBv+eR/Eg6Vjh7JFXTrqxfmkBF+OQA7V0U
QgM1ZY8iY4JWQGgJFxHwbsePDKsiaoDU67UyaxKXEswPLJ7wQULnpdOPGjFCBegvon/5TqzVHdud
I0ama2YePhGEAAhRGrzjvkwe+UXk4aIPglTG5F+ihNNjg17r1d/1jAaf6V22Sy5/CnseyFwzmSdE
7LKEN+aAEyZRNcabrxJ5Tme5oeIWGWwTLIaO2bTBsHjMG7yc+zIUIAy6wfTc/ZiEvAY23agNVx9G
AhaYPMgNvRSS/mQCyjuGaxhY2q4y27vbaYf53BBskkWuNoVxZvt9nJ4ZnqfmCF8675pSMJdNnz5v
SgWkDZVhd/8xfI/yyKgnYrh44e4ZAH02wawvyhV6jB1OcFe1NGxO6jn+VxU2JbjL1ZC9unMXXzgC
TiL207l4PZg6LX9qwMvmxl6887FzpRb7WTpwr8qEqNBcmVMFC8dtgvieiyV5owe8DqCCdy8utlA5
vPaRBdbaeQNX5H8KUZdbNrdlmjWR+lBvN4oLxabyetNjeYaC1yru/wOfwejGwdx+xBLgzcmd1pLa
QKyJjEvRMUfud/aTNZUjC4p2BKVYEBFxg8x2UrraFvXP5QIFXVpWo92Q3yImhnB/X3AT/rPuJ/Ph
4LFREyplbfy8pIhQ36oJLdveHJ+ie6YmwwErEA6OG8L8TOpkc7JqNRs8quJINmleUnQVgp15hc9h
3FNurTFClsyN2JuKy/D1WrRzC+UV8bcTMPYrjkPnSt3lDjxboTNRp+AdgY6OdrBJUXxDDFqvWgX7
le6PHyKjjJdgO48TillC839JiNTjUKpNgqTuWjTPNhQK4Vdl1j754fq2kgxFWKWLe4AKh0WNnWdH
LBHFIh0NUs+aZEAFFCvXAwr5evuoi2fLeksYBvzzc1Mj1fGUus7BJsyG8f4HkwKToRXGRrZuARmt
tpSTieV6NEf5VyG/xH/irrDmshwuvSlGsvsNcH1Skr35HuJj8+SO/oncNBWIT8uFe13qGMzohGHL
yb1MM3c7pWXfpiZMUg9ouWq0AtbPgRFN93bhnL/BrW1VcU38ker2GYl3U+90vGu7bTFBc5V9Hn1G
AY+K63ND2y1TsRjZndIK9f33lSxQdZ/kQCZo1/Vj0Fk3NzIpVsfbXKYiLuCIfqV3mM17gBhHhgEj
wQCZoNrPOQIjkA5RS74Bu2unSFOkeVR8x5oovGSoCZay4r6Sk2wWilhYkD/HdOkauSd+rcUez3id
6MdhYAsf1IbU4EDZLytOVzsOTeKt8cp7viIUyJWz4vT/4QG9/Bc+GX1uc1JxyOf8vFSDEokg5zUx
SF1iju8Q4FFfKwm2B53O+V6YQNvbvsCWUYyrLLSz9trhniWD4mEz/rEogQLkCOIwjGPT7P4QenVZ
ubeOP6joEvSNu9vEknpkyMBqaMZ4zjLssmw7oBVRIyulwhydBAPxl6OdlQP5uLIk2cGy1FTLrGGh
+hoHaSLs4+agWn29Jck+HLHqu8ZUeSKH818/BvQWh4meQkWvtzcrYijSML7WUsmWnbwZVxiFrZaQ
gKX3AJKaAJmRvAA1IRnrj703kKN6dGO/uZRKSJomXzwLt+H7e9kjmn5ez1fh1DckAZ+qcuPIB6Qh
wmASGJICYNL2SGRbN04+0YGtaF3Teohk9kuSKEyqV6WuZmg3J489jUMqBE/rHJjAOUs48CRZXiwU
oFbyv2kwj3sqH3QkCUvjcm4ZEZc/j4ipjeIe3tTGkRppbPN2bb0HxKz7sU8X/jzJjUPmYkmkLpbH
3abhKJBPTHYegJFYA8ojOJ9Og0tTycS0PPSOgw2cw2ffmrwvV0xsTVn5ztidyLy4n5GBWLkU3RvS
scTJh7NDHkqfaGvxEeg4wxSKu6C4ZlEEvMuDEPM3VvdMf0lOgWMAUh3042j3mzzJJ6N/FnET5KRj
2zimDrudVUm/r0O/LTlmo5HkUstHszoJOX5maN8AL/COjJsaQEJdARFsaZRFzYB5QEvjKa2C74zG
I75hQYGZZkq1Sw1NyJdh7SJZTBIgdDQGHS4e2hBTILSdSG9LyTK8H2g+tk4njaN/fRHp+68xgTfR
JyXeekM2pIZ2/HZ/W3ngMocZ+3Wkl5OayKczNf1y9MpEmsff9Q8NgL2xGR70MTglY1lt0UbS3D01
BkkhLU1e1erEmCHVYtwegSIpSkX2HhQrGbIzpRwXzDl7bS54rrZMq0e90GEh5S9cqN4dkAUSrLzI
+FMzr1weN0MROpATJ1FEIic8YXkuqO24C5At4IM6y7+mAkPU87GHNgnFbozEzD4r/lYpGHEgMyOQ
OiQFOFlsVVRTxjCPSKNWnAeLGzLgA9iV3hv++jQDhxoSZrnNR9bk1ffGOYaxV6Z9diJbTPSpZojX
am5gHnu5ADQGtcBxa42ikS46Kejyn5RtpBABA+WCTdoqXU4oUXxDbvQuhqgx9sau1YdNOIMxeJoy
pqI2gVWGrx4UE71OsmAoNrM3enfU/0hehmOesgs6Sn0sEUX2wrvrHNnR9qwEoGG/flcoXBVBLy/+
zIiBXDkqSK5/0daZVh79ZLrkos23+puJLAlor6sKYljGJhftkRqoekohPIGxc2l7R6l5+7bC//X6
IdLEYug0D0NfqO+UGGy9ClouoGZekTcTFL5DKGVVsYdwpc1lJwqRBO5ykC09a1eEkX+SZrB2X8Yr
OhXyMKXhzNMWerv7A9a5QuMgg75w2v6D9bX4suSQwhUsOdD8gI+/Upxk+kkzxYLJ30+lJ1954xJ7
YXQ3KOVomgTWavp+yMWiG+H3EsDJDmh3oYriR6vECaayrJxCNT84AVA+HYa0+HphI3Ytdu0UJCn3
EqwYSvu1B6BThEedTPBE28oKYjTRlPGzBmhwO9NL6tTtwzeziv/YPfCuaGJY4PTZRpY1lQwsbjTh
Dq1KvOspC9bQ7Pc229jrNbxi+7tyPJWWWINv+s9CUlqCRMOHbamJjdrHpQQVSZrUriNBXspySsK2
y7Igoq3OSRKru+t1UUdBGuwKoSDyF7c0qj/xbvw28IK2Yxvw5rODmAsoOo/gQAfU8Cs29TrhbDDN
jezR3X8qi46yvNw5wEkh5Woiwfw380UQwpXsmKH4Z2DwYE66spe9JdprNrGu7fh6CZZ6L1Mvwpll
ZzBvsGhM8DU+kU3lU3S57IyQHvAgZpBZch6ssPdtx02k1WsQ4AYqR42MMYEexrECanhRKpDHSPnI
0OhU5HjlOSHGdkot2gvNI0cFj4p55KV9LRsa80zTA+LUzn5tv88lBQjIijnXy0U8V4vVU8KN1hr2
2d1Q8PQWVh+yCaKwV4ChgE1ft1OopDT0r6nYSv+/0Q1j1ZiqJ912kU0k/DF8/DsUhap+L6pzhWoR
0W6gwy0HgmIsS/DKO9cTYh09nd5yZbuatMksibSlALegEBTFsv0t4/M29L3AqQWPyS/fsL4mS4bl
FsT/pQUUQVFvbPhcg+vYvOjFRz2lZ/HyPMGvYf495z5qHN03DJfEs7JBux6KauPZguiRbXVy7Ob5
MuSkmhTf4hhvXClk6W4BR1zqJc6aropE/G+sx2yFCe4xbLES/lYHYrQ/rw+hudH7jA5fcp1TpD7p
v9yuoHLlJiMJHHbRPZskTWi36+SNWmci60HFyIt8Jg9Yc5ee8A6iwJ6qMPVJisY1PfRNMf8/sQRy
2sXtiOsxOREJO9sgDeu61I0uutaxA/iFkU0/KrAAIvOYUWh/AaP1AQXK4Bxd9NGhyIo0qmsEmn1V
ANYz/wlvTNh7NiBxw+opBiF16clIojkDKmd+fvup2jU0I4D3sWGWLU5RxI5HbG+7bTUAHKUFzS9C
xumJr6tWndvxCOzDXAdsENVUSRsWIEprhkFihnGhJKB+LQhNYEaQy88JGgD0RIVajy8nTxei4p/3
y8UJ5co3qzhFg37qvYXFqwF2OlpuZ7vbT1UsxTo7ykaJLe2hpUU+ya5z0g8MP7g/RPf3fA6zmwBL
kwhHXbUiupf4VBuQhHbtMWfwzgVxygmJJecVaDH62UbNrO00YjD09oX3TqQGcn9KVeNtiGGp8vjL
2yuIwIcYej5xNRW4NM/6f7xaDX97IgeH+v8QX8Wbcu9P8bBXCMUSCbKVVi/RbIBxIaf9mZldZTAE
I503WlqFlpVA8rQw9QH2ZVz3BlSMHjW2wvYKAbhAvHV+SRCLy7TO9sCRDu3rxXDoTWIROCholxb3
ksry4u4L0aUWDWt3y3R0TRN/2g6rioa/a8wB4cOFHy1mbBa2srDb2y78M6KNEdZ4fxeAukAuiK2J
CF2dMQZJ9geS87U/2OyhCwCH+hIaw/6HoJnUnbgKK4/4eS84l/n4UlhHBk8KMIL92jDo5pjSQ33h
5+d9WZ+5SNBzxUO4y2Nt5FthwyihLos+zZSvq952pKBpxpq9Ozahmuwx8rnVDD4X4LqeBln2wAwd
9Nq1qSTmQWzwMkViovRgaYmDjEb8jeTDlqqvwXc8Ov1i/PBLbUtEIweESihl2Zvb7md+dAxYbNJH
jS/smfpoc785x1A2lheZnhqPwG1e9dpJYMilpEcUmT4NzE7Z38MIXxwUjIocO36DbX7vaH74PNOQ
i6E0kiqF9h2BO/cdMjBrzRTtRGRllSyjmpIQZRxlQVI2QyjYz9gpEmWBjiyQmhjqEcEfsA8VcrNU
lsDyqRqd4s5t8HMkgZwTYNXHvfbACe3TBl4n9qCIG2di9rqhCm7it/plnboZ47r66M1hheCmsZdT
VuKu3qTjCon/xcgXsx+rjz3IS0OPIhvUcafVGeNWRDdh2506b19thyZkWlb2bT0YRsPBTOgw28+k
nFShfmYRat3L+x9l6/yIBhPN3tIYos4P+lCrnU4AMJ6z5aEmoS1UQrD58nJLpsU4YYQVR0/pn1/s
upGywonjvQwHmUMaz30/vcquskpI7bFVZa+0A1q/taW8aSL6PAQsJrFlIpdTcsufBDN+dP2H61cy
tBXa8Xvz1xqni3SI/z8L967wIFUM0B0kJJDoy01sD+/lXZtSVRqZc+NAeOWsHiifb+Mw6yLm4Psr
sA3JLiPBjXmUMW45adEbzoIFJbWF4vwKDxPG2rABPZVW7RChgx6YHRq1rDW6CjjnZJG8b7j3RYJV
85+86vbhUCIyasdiGpEK7EZwponA4yLlMRsCyYxkoCrmM9+nxbnwlHDtXigmYlNhu3fYF6CO1HcR
ievh7czk9vhrmGTWqNdVIFVFpzynO3Qr8Nnq5rNvArV5ykZEGK8fECnAyM3SFnQ288Dq7s1gu1lG
l99VmBIcwAduJEERlQ2un9fSxdyI4VhZM4MivhD9hD7pOS02gfxyg6marYnSNJr0RsYeKciofQqk
h1UiWETJIGdLkH3UgeAwAkfXBESC+mEaiXquA5AilW9Jp7lWq3VIBIdp1sn6EPpQDv2seudaXf8w
v7623y7q4seeKX5lXrObnMzKap+GfjzmN4BTvIDj+hhhk40XnNTZU9ri3s+dU/33yBnoritlyhwc
0O4gQRoqPELSOLnnl3LqLjGZwAij+eGN/BD2sXmGfTbw8HRcJYMy4zGquSW6Q+laD/Yp0TQGMI2g
9tR2srRrgpa7AuAjeJJ3vV0fD/ZtWKtsWfkf+wcZaYwjSG4qv7DLkeL1VI40PWigWULalTKzzo4m
o3wrITyW/18srcAqKBZAfSFJ31IR5irX9n8T8RDqEOmHc6pKD2Ie3tynY/f8S4aQmPokwayKwIcX
1X9B3dDN+HQ1wSkNHjPyqLryyj+xXgKxHB891wZdmtXjY37u4CaBuXhj3em99Qf/3vfS8SWMjkPU
T9Qe5uA0V+dPWQJ6Sdqp+3HRIgcXNDiRfKdkOK40gEOtFayKp5MEhU8Vdqxy7+futh8kgHqglobU
nUQXQxSUT5UdIWMMjIWugBKa0ktTZMCP4rhK8kLS3wlaYvTLBOLT3a34BS3+toKoYwBuQ1bGuPo1
5c5d47YKR4aLxNtA55+0ZYxaSYB2xcE/cRO5ieEWhv/djYD0vTiJQMcMVTFof7T+xJkixaO3haGC
SQxvdeVlGO8FawnbCNTmbtaeBRV7rWfYULefoPM09TtQnmY9NA5+8ElVMTJSgitKse5KpEmScJV1
yU4NpkYdIhN8B/LTnzngfsO4+jGPGR9seTVYNB26YSdxhze0Ka/BbpZ6nCMFRrUnq+Gbfjw/wfO9
mU2uUlvDTLh8LqiaqqLGbpRvvZo0jddoxphH7kdEfkuu6pOTVXRPgys2gQm4geSUJTgdcL8NruBo
5knr8WtU5HSJJnJ/WsWq/PBE+b2/IEot5A1MSJjcoABlmaAuDsRC20qT603q8E4qi8HpvHuqFo1K
/Z/rbx63gJj605Uuvzi2DOc/8bAdNfzuB4Jbuv6Kw7+4e7a662W8JYwQgBcBHArj7YUUyF9m2hqJ
UVu2zT4Rrt6wCAj2C08OC6vZyZEvN0l9GfY0a+uyV7dv1duxP3pMRg4Y3Ha5XLwVzDi+CoGnpn5/
m0nmk/+oC6pY68TnyW7eC9+izFH/sn0rwcXko2ZWFCYHJazqCoTmj1PMTFKrDnI6l7BBmjSE9iBH
scurds+J1q/wlBxqxXrntml1dTgyevW3yis3tsZDXouQT9wseSqk1sT0Sl/z8HYeCIDP9NdGpkhg
ZfktCVv4hlTBqA2X+AywQl/h8b2tC+OMnKEszrvuTSRcR4taVSj7Veobk6eXZDSIgh2A/p+i6wVN
rRRskldDpcmFENOfExKMe6Ln82p9CY0TibyUqrJXjiVR6dP1bJLqWV4j25D+vtSbWC2B9wXZT1IC
mh7KeEtP7kbaCcY+9pjduCKf9Zw+VyWIhCla4uxGCMYlXU/JlnJjn25PRiIkVgZfexEBtGdMZG/r
YiPcx+VVHxkH0V/WSHPrvZaQac1axmKG62Ggnk+SUQLksvDtvjweGZS7s+AKcBUIY1u425u/enyY
AAks/+p1dgJx7WrfU05Unf2mh5v3dbH7G4uDWQlkvbY4H3/1XLUi56r2zNoK7Kvk915ycLqkp4gK
GoEp5LsTPC1tJsCID8x5SDr/UPnwSP37KXNs35KQ8z9GSsC3tINQlliQQgPzW+JuHe64pyZ6V2fr
AJ04IYMIade6TGCMRxUKdStYWMKDvRgZE5aQIGp0rQqb7r7Hql1x+msdxxaGA49FF6WRc/RLQWzR
VJLPod5ahG0tiFOeuU5GuLFj6/d+2Gv+BkH7wNH06D7NsHuq8CQdwIVO8eyqhVSfm1fHZMVcl8d9
rji6fqq9KCQk81bMY39WwkU/H9guPijFuhg1D01N7XqYdRevsomrG/6fXqdBXMi2ZivZbrruwOFp
diR6PZajH/k9vWM9BxONGjb+sW2K60GBQK12sOzIjbjuwh2TlHV8GYYi8Tp1IGNYlHKG4K4gTgoU
k0OKuhPEgNKGjLyTDp+301pHFGJIT9Ca4MKouVuZ3dOmG8Q7FLXdE93/xuTv+WonTthqMHgfsltL
5MhEDwN3fKgNK3qfTQv52ilJL31dutqJ0IRLYV84IZnU06yj64BI07T426i+pGMxkK1BpTnDUJT5
fQnJwoQKd0VUXAotr+A4VePLAvvj0jdfXD4NzAI2tAs8Doi7CNQA8tpJleL84km39Luasr4F8tgX
EyDsmz+CaFT39pgcvHVjwBDce1YW0qxE4V8vXriv64CyEPaGfqiVsNS00iyeQKH7DjrrouK1bEHy
L1VXv1YcdyMd8+t8E0hP1QpCLo+xzxaqiwSu3284FUUOstry52VDmJq7PupaNgJw20a7yPUZj6OM
KQQBn+V468frnW9U5hR4yYf3w4Sh08ooFOSdx8CIKm9D1Pj+DhFucIw8NlRvC1alXDre92Z61h86
JwX5H85X3eywVaUE6m8MUiBtO8sJ4mDqUXg80d0M3Opd85jLjvC6GN1kefavZ88RRbOuLFV7AhJW
Bh40zOcr+/7OVuS0vniz4LJcCDUQrOEbp8ZXqZ6+oS1h3vHhL2sSdqXsrhTehB+aoBJxAxMvti5u
SMTbrDnaqGSyp6XGoDftTsFIWXgQDk/wjf/iXElHjpnHF+Vy1+8Ng4MAliYh/aSgpjwQvUQw4MLX
woVhLDVvaO+M0DYSDkhL3MA3TIGCAdiqhl6bGkYaMVMtJM44TYdyzRsjkKtPl+vClk6oLxHJ6Ana
UQQQiZDelubUuzUWRDNs07DnnFaP1lcahQNZHoKj+IfLQd/xbGcUqgHViY8/JdpjQE0Ne+MTzrOO
yZKnFY/0m2W9jVii+1041OzKeIpECF4wru7b++Xa27Fa3NixqY/WRHB86yvf1lVUq7LRITzys+m3
n0ySstPusGm+WkMeWztnJWTNa7kc5pT8gionUn48zr6OTdGKaHVDYzE8rfzEHjUXCZIsrDPce3lF
MH1zmkHobLJY7G6Bu6dgwd5VXl01Czxh9t9zG+STN7wdZg4puW3ecbYkYk1EAtOqEh5sGnkSQk4H
bEVY0wkvmhuUolMGyjFqLqTGzGGe24p851n8M0sIV3lDietMjeyZ0Vl2KDSvRCZzB+Db6CgNBpgm
qelAsUzXIQ1VL0uYVHW0FnnCRtkPkWIl3pzBWhax+rydW+l+gRClpRyeAWGnpeSstKe40MKBgIQJ
DQDZQBYFRtOS8MrzqvzDabqSdb3/kXQ6IVkcZu7dkqvUTbDizw5g1HprNWKuOc0bLXjLokl/qegl
REyF0S3sAAAxp8jkQD47BXtr5hE8znaYEMdvGfwseSeWycLY/sW5OG25JBY4yKDUVlTC1xKb0f7+
KJe08kCqeVltoXE1p/fn/FriVZ5E8j6tsEVswexUwmcGkQ38CuGu1dSyxilfdarc85JnwVizCCMg
XCJbtCkg0IxSmCR5g22S3f/TPx88keWalhxy/jlXab5hUfbEEaH3W0UvTTuxPvFNGqiCYOMR9ku/
Hl0s8jKpL8bvsbilTOWPI8AI7/PWS5cmu0TzqICLSUVoXWW7SIrg1rRc7CK+fSuRbVLBONPRGlf+
ojCxZ6aQJXXOyLsR747D56AtfhezaN08xmD6sy4dOzFYTconX8ALlp46rX84zp6hOuHRrEMFHfhO
r3hrZ6KkPlyWkvkgJ8w92bov0H9NB00iuRYIe92dckVxzrtSDrrVuc2upowsYXGcuLzocRDvOPen
/a3nRR6X/BkPZ+aXLpqa7oPpsV5c1vgdc+cMdtYwtQrpDzeE9JqhRvQ1ler+sKvf7VricNbXe6U4
9KQUoMHoY2PygQ4d4bQM3d2Z3/PboqU6mg7v1uLHOyk3EUmN6hQnLwdymGSH+v5CiU1VziqEoRJ+
TUnV2TM3oujVFS45zeKel3bD9+4tOQKlpER7hzmtLkk+htZGe+PU2tdoiU1xJtk7I+zgQ3DLyi+9
iPI0f9xgq3EQMtNttRj+cJlaR2Ukuz2uSaX8L9MkT6HRJv2c9CTDOi0HBIYchJbZyJI1s1LvKwdx
gWgNLcABjBGShodaAtsvQJCwrKbAUY8r+isHQUOM4HClT6j0oPF7S3NPRtCLNP/4frTYe2M70cU9
bkWKG3pbcbqPnRBVOKjH1l6nxy6Fzya9TwyqnsrGd4KqiXqwdpe7AMurZwthu3D7ON5PCYYfVHI8
tuVcpp93hj9Mp+U7PuzbC281mlOmWRiVwA+XYx8E9/cg1hKoASiW7S2svwgYSnnJgH+qwOg7N5SQ
BFJamMEGn5IunIJIA0GUVkKoNsmcezWmrI2ffs/huJUGwxZUBYxDFcFpax8BtTdLWStgw0q2UP98
hmltDCvdKHa24f2r9DMunRAythxOeLiqOCwJBM/styNBF506zdbW9VrsDaDveefmaoc1Fd13YPa9
jUMNXmvnJHzbBb3ZgpsNoezOZEHNTNxlFpBfmWoY0CSvJL9nMA6Gu3eKgBvrX608ZNe9C+WXBjkj
jO0Fd+F4j88JESZNhpFKQ//uTKy7Y8oo1zAxJaqSncsJkyE9TLZPW0yfP4MbcsJRgSzMopeISaKU
mp4u9JZUwRAzQtGN9lqvHAusNRwh4k2vpQ9bKD+s6cofjLv4e3s5ItKcfZp7NvsDtbVQAOA82rjk
H/Zkzj+6Q8fjUSkaYBsWD8e/QZBHksAhyut5skjiu2juSZ0GSGdMl3VIZP2NAR/958r887Q7lPQB
Fro9wrS//LQDujbkYmTjyuxSEtJ0oNiYpw8JlTHFMBXIWbdtgocySysd6sFoD1gkDmmPIZGO2K2z
NkN/wf932RQVwH7xrlIHPhrgw0atYmGpG/Xo8YMs95APRxD2y6YL+sLPjggEY7SSPkRxRVsExzz+
lEII08EaqBfzPQ/qzz1v1neVzn39X3D6D5pKf+qcYIuPKRyHP4gtDkEi93NLw8nQNNi9CO8ftMJ7
0DPvlxsNfe6yyTdkz/bJawbMWQrinh37bDg78zbJ1OlYHEv6WCdIrgzJp50iUhbOLm/gke4v1VSM
mzTPOfjKmo9xqkMQmoBqRo76WdiiNYZ7Ios18ElJyYkoApjdgAfJ9GyrSvdNwcCPM8yNW6rSLaAB
nz1HSvXkvzajR5Ptm7KvyGL6g9zKV9bFIJRM5CIyEI5++YunuKcN0ep0j3Plv97O+EVeQjepIEpx
vFer+P3eFG2okd1bentewxShU2gjJrJMOChc/LnO+tv4pFhMRhx26SkdaZ6SQHaYDQM4hwThKcCD
tCyRdkKvsEkViK4sErvIJ5vBI7HCvcrg9SL944EKXjJvJwZ7QvKf9m4ehWzUjXvJ9XpZeeaA2UAo
w9DDt59cSwHV27Xmr8ruEjiQJVJ1DlKu7lIp/okTm6vL9m1beW9ULZYFiKt81jHhloFJUr/x3tMP
c9OnVsn7T4O3VlWPdShvkgepVyqmQCJxjL7l3Cs+VK2bK6mT9XHBW/FkE+qw7EM3r9C5+oLTMRID
PD9kxnBuKyjaygoQupofcrMrGCduDBhbh75vMF5zRaZJDi5oBVK3kgDJeuP06su15tAW21RmJgMQ
mqP+Y1eGyBo0fi3TyWWfrTFtvT5TwBo1PgnWOK8kOXC6KHqE/eEHpBcQUlV4KjvsgPhsothcGwVi
buC/R3ZWYFM85U0QvRlmJngeDT6s70UpxcoEHtmJWQqdNera4/9YASnIVhOUWo3dkp4F2N301Q39
U12JR1rkcX5ZlRCQWoyelCRl0p7JdCjax7NrD/DgEMA2qKkmI6JvADdYM+B0nOLV/MM1JB9/ABn4
I7mFH3Pi8b1YgW41aykY3+OAlfD+KcAV42CX+IREhcOl9caFIxB9KHjqk3KXQ9Dfh4yzhtIM9WFP
ovoKYLhNJ63ZRmcLYJ08NURU+54T4vHBkc30nINS0+tngADsPiSsAiTk9LjmrsVpjFJIVqc38VDp
i2q/Qak1X7NL2u9/1QGzv80DKFOHAlm06/bVO+iGRTOV7Cv7kzWUW02F34CgM7IFCZ5hyU7pr2a7
thbfUJacYQ6njFaEKCGBSsp761mSSiWqACtHh0OxNej6K7qfXoKgQLNFzJAu3xyH3NcW1Uqs3MS8
JC9gn6I9jvvwr4ZfQl6mZDSxSyZX62aZVzTTcEOXPkvBrLwvcF+EVHrzEoemjDihZZ4Jw5AqjgDl
s8J8Xxl4+fzodqYVg9xn8vq2sQ1Qgv6X5U2FieFhRqwx0LMl8duSg3als8eAW4tdo/96sZaTIr95
4RAzNq6qTKDh71rVKrgdUpPlni7XHn98dNlQasi7eAMmgKlqKfRT526TrFwd/IPXJSst70Edd3By
hsU5E8IHrurRfogQ/V1bX3JGZHWrkayXUNnqyrnG1Ju6hw+9tEvp5Lz2xA3LAOZ3eOf/B5kvZ7S/
wxAbQwMI/3CTgZUVFsRt119e27Nn3U+umEzzOWEkuJDHoRAWmpZELil1PFzxuc+L3FaJyy8WEeYU
9SuxKpJg/Sox6hdhJNpEwqqg/3TYF5aFEBE1QOaaj5BHqWZir+JVMMmQ1jMnVqJ86LccKVovfPJp
Yf2rwfq3YvvLglcqSsqv+p9k2mMbK+QeDsXJqV7ajc78hFhhMgLdE0bJSVB/NuLqUL+kNzXnu3j6
ZomhOUGq1T7j5Y5QVH0sGc2Q7JAZowUhi5YKIlfAlGTacDpKQzT8jampNQ30K/4cV/M1kjWRsmYK
/T9kMqoNRLfeOmLoctrdGQcFRPD5nn/vdt5/JadF6RcZLE4htry5eFq6ZThsrg7SxHF3t7IL5FKE
cFJ/gGBx+x9Wxou4+2GT/f5VqeKZuocLSGj9bz0S7bhN2zTcOIymGgXvOZFalKfNS5pCKxFGZKAS
mmghyHPh0UaxT+BfCSWQ0ljimX6P3H0rUZnHYki3VCX4dJ8EScLJg7T7M3u1URBJeGCiKEGEfCfF
O+tDxMIq5eqBzESHt2YfI9d4UTUid2WwNtpj6i9uPHwhB4Yd2tIVVcBGY9I74jK+0JNxCyhUmmok
appk+yFxO+BF0kVHKOo66G5yhHKmiGDs3vseuO+RMit+cOUdhfVvpaPjQdpydW5kugfxPVPFw6MK
OWx8iTxzR529TwuoP2QLOnq+kPc2ceuIby3f3UTXJMd3D5ccXqcW3AwkmDhnCtgKWKLxfSPCP7g9
fuALMAmazNZ6IbSZrfbOVsn5Ywt4LVv8r4E+1skp6qsFdZsRQR33YL3m9u7oUMMVXFqBZwPjnY6z
qprxBXCJYkmNX67LxQPnrDPN7gSu71kSZWSFeeiUmQ9aKsJPQijN8eT/gnp5RyWdaK6E1HB75uWB
MfizKyJVIjlubW2mjFel6RxahdRtmOVGFeczTAS2aozyColFNI2o1IFEXDtQCJJxoWTAtEitYAvw
uOgC/x82K0qW28Sz6ab5sQ9wuUJ2aFMnA1/iwQiU42nRSfKJGc31tyeh2v2w3/XTiQT4WBU3ExNP
EqOHxqHAHKc2mtQKj6p0XO0cLjQxT3uwtWnJ2fkEXNnSDHZotCknEj8f1GKAbEVM/Gvi72zdC1mP
b6xWLQDosPyK0YdjotTyThz9+mR8+Mk2pTnpk7SnSxyB5KY9I4BMOZ4Bo/OgYlOkezhWCSZlr2mp
hzZ/Pj3N0c8OSxj3NTzGluDc0gB4JhINm7k0C3mvcbzk4ZiSpOl0Zd9gOgaJwRxUCFn88tqp2s6J
F+dxxU29ee3/69J1uyWHfmr6lE9GUIYJ0+HP0G5vGsL5Kf0srVIx3SIryZ+y+qTjKRKd/BgglRVH
ZdkPCS8Q3mSzUM/WuHNiMRAOrekevnjWbiY+ZWnHn3jGt5yDD0EbL6uFM4h16JpLz9szbZTD0fPS
6vlweUW8J12CeMRlUoMM4y+7yOJSKIGlK0mI8pPh+BsdeDRstSeACDNSH7y/O8uHVbUgJNXRi2R3
PEAGEIMi4fRvEHsnRuSEa2Z7qBMr9rWU/ytn1vgPMtCl3m/bqkfidINkQxgKmzduUDAb51c053IN
9NuYiecbJVUTCcpxmOv8lKoP8CKVxVPhE1kXMvC922hnn2w8t+SwWXK30LqEoIXg7gsp51nCQUc0
7gcuGlBSBi95qU6YuDf/l8q3lXThKBvUfxx52v+A02EMHbgF2gk0EyNqcG5e/+dK2gtsEQDQIHkv
r2BOEr9ia2Aow3SVhkldr8rTmQjvq7dZR9tb/AQLeF8EIQtQe7kd3uQgqxKjj6OuELpzUvE6FiPM
anVcdQXDQFQZB/rpy+IXlWAQeUzjyI/VLL6sFHv0Tiyvs8mTLCxmCcJ+WnyVC3/Y/1Mnqdg/Tajp
S6tC8EZy34hCzciFhdfjFm5Fra1zz/UpSRAESk6n53Z3F3n9Kdn6zvTZ2FB2+bAojcsjSBJMwcIL
R9QrhIiNvCg4ui2bqFqnW7o4+CRJ6m0k5YvUArAvSbeLWbM3aGZGkybBiuL7rFduH47lNq7Q5JLM
BlvcIacaaZqxTSqx2LebH9vtTTAA93FAKO/Q+hP+8At6QUfzY81+BFGNtXd21S12uZxVfHRKTYkj
REGezsMcDXKPaCvFhBvF/dFOPXtdKqkzwPPqDwR1q7yCfMvdYDmUeVT3xTfRG1seSEQW986NZ4L6
LkVoC282rQZlzxImARyw0oFSi9ZAKXedXeeZ9FCWvuqomYNQZ9QWNs+wCtwt82dbsou2uxlv10u8
n/m6bQUoqPxuWnYYBgX5kC+H8yIceMMAAisa1kn9qKsX+4odF/lLar2tdqiWXTCOEzsC2GpcPZtd
GZb4FfHNQzQNmO3lw0E1kFocB5bFYWvU57r1icN6K1kRh1PGwivMGoZp7iO9xyNWijwdpm+PMQyT
aj6uNmzIkshB6pQIDqB98pn1gC7Nxy7lo45rDzd5amAbwqA9dNZ8/WYQZ69tp33F8g9QGe9AU+rx
7wdRmPCMdslbme8h5P47leu8kJt3a54zeD9Z9NDICHeVaiwsQuQJ/+bbIAusc/+V2hGyS4rjox5d
DHaQLA9VC1bBCo+Ccne6vxCLRwdtqBeOU4617FeX70Ahm9iUtpq9v/GLCGgarSVfvAG+ubLOEjAI
BIeRIFt+zzgPsrz9OcFB1vxLzxYRsN2g9e4jd0BvPW0Me7Y3jP9WLPWGsyqa/zdMPm/o5GQJ9xy1
X40uLpQ/sF4OzYlz5XWYQ7NH22UbbJZO7JB4ktqd1HfjHCa/HGiCLNzMqKUdLIrxIjbBnViG6hj4
R/pWrL1Vfm4Po/GUeIpcPujSsT2DDdDPW5nBJZouGRUQEEZCEPYKhfPKozS3C2Db73Ra3nJQO5SU
Q1iAQN5Uqc1UMBXzkXAsA463LhrBs80gBee4w16/AZYl96SQvn5LkFZfwej8IgtHxyphnPl+YSoy
efgFpk03M1AIYynt3Rw1p5cG3QPUMBGLlhAtWDfMOlUjP5OXu6t42IBgJCpi89Q7W0MiKM0/dV/2
s0snEak4ZDr/KAYGFrfhi02IH5NRzeBu7sw/ISdjJS9S3Gp7pnIYc3ge3UjHE+SclVEyBejy2/D5
v6D7QH3pGe+PC4m4GyvmkZIVIoLvbST/WxnIJt+LF9mQmsar625Arcco1CYs/pBA/XoBMPRfLhDA
bdY8qlkHwMfsPtjqFq+yUWlw2zd9J2ZabwtT8JSIGlvHdb6Q4IZ/WcOughH9dDhjKSrl29rhFokW
ZnLi2uSCuG3MbmnJmX7BnnS/zTRZKhJFilhPwNs8QR30Qa66aSKeq7K0f+ZM6PlxoWeyWBUfvt52
Awv4VbZ0DjB4kYEO8jeTyLsoavFuFEjqaWCC4HDK6a3ar+WmviLnOegcsO7zghyRB4+A6ADPPFmQ
bFUUoqJnrgjnP+gtXSaSxuZ/jDL9/JG4qBbNI0ZJiPnHHLl+T8jHrxzA8yj5mq7CpwY6N29mveAn
T2L8EZIb4swF29C1tBMoHZn527JQkNqhfd+cYadwFyp+VVah7zO7t7t/88Nlek6xDspCtZ+9q7u4
x6F6KlQavRW9B54moA0D2eU4fjWW26TeHdTOOvJaaK3fzq2+VKcFYmiOyfuyV/UsULlwqYZeyE8g
K+q1qjZosOW62HPfan6BKunfLy8x6HXRCDuhfEhOapllBSa4RmSmxjE2Bj+k+kpY1/BZoG05dBlz
48wwfYlY3AfU1/JyPCJuE3JzlFVV2uRiviQm5Cyat1kMOr9jzblohosQyPgBcmCjBKDDfxWvgh0r
+9iZpjoRUAh3xZPOzVRpLGUqSjVJLlAG5lje3oLv4QIXQRvNrVAl2MygF1z9wsBE1M8H2Pc/KaPp
a4bnw6VlqSwM0jwAGGcXc9BDL8OqEVVFB72dCsWeaKyNcb3ailRBbdDXAX0MJasczHZo/gr1ELxd
siRlIZKemozDEgtSwS+IsIVPxg+5ZtCGISDWm/PDmYGGP8HE7GgDdriK3edwPaxB2OR1UtNkDf9c
r3kJrjfZvuRbkc0wPV1poz/QQS7fWpsyCzg1x69hQg2NmfOoE/lICH8Hqa2iwYwV5QQrHc1AEODs
rebfziLOPGqkI9eZdIKK73JRJsZ3bZOfr716u7tRkjXTpqhCJuMRTMTje7nKFSzpS1qmtUWoyDss
2C9NX/gKLEgZravFsH9dTUFRuosG+1Aj28VGQPUXKpTejRgYEF4WJx+gJ/VASuW8aaIR+Z6w18RP
5HUUhDrXka+WC5+WIyIv01hwL7sW99z8kNFUob0af4EkTRXUlFSyfGih2NRIBsfDjWbtToTmCd+j
/NotsRm02FevAMT48ffBxi3c9uhro+QquU5JHpbUTMW1uGCop0DfWlW/kJ4XxiDGiviVTtLus7M/
+NhX4PNzxULgODZR+lCRFyrEEfuo8MJv9SoOviNWAkzf07QLGKYUkSjtj0ljgPwYhbg44X3htBgx
c1laYl/wycsbB4g8x/iBuMNAaadLHjkrkE7WlfpuyydtZNi1nCB/vL0T7ITuqSxICd13R3TcdYS7
LTWMPk6hSW6ZruleQUP8Ra+2xzeBbzuof+7AAUa+NbhCbj9k/wJXtkgmpzS74qwzaUAkZP+jQjcI
lB5mAa73UMkpk1wo7gVLk7rBFh1MUdXTyOM+SO3e1CxriexES5yfvRh3awqRLaJmb8mNmQ2haUZI
TD2ZvHsCQw6ejsDK+sn1gD4lD5YJSXUr+OehvlnKlg9itu86ob1aPqZIGZ+zQagVW96AJcJYDYZK
EOafdgQ9cUZs6VQrNQY50hCPWes2Piy7BPkjcF9KqAjx9/gGFl2T1Th2W0LJ9e6ic1hRTy1m3EJE
NfJThUZARGfJ88EHmYm3VBosa67z2KZm2fPJyGEw4YiSgAVxD6M+VqP+BGJ16GhetqNUQo/ik3T9
+82uyVaTNF5gf/ZyHFs1ucOBjPbi6IDFsKE4cXAloFwh99/dcXiwqnG0XAtjeHDle5NLSlkTdwFo
05KuMQqDT+QTBukB1fkcjrZ8CVc0ceBZTfkyUQd2jKAnb724PDdcFqc67QTXYq7vSzGBZY78pryJ
bZS0/+Jis1rpAC8MCRxvwKbAaY3YQJDEvaAK8XSNUfDUt9tC7lh/cOc2a+ssGMCSZlcl/b7nYZNG
zjuisEu0tNGcfgs1PgFG6hPJQVN2lXpJ1vOWJimZYWcGmOxgWTr9yEY0yt7vbs1U/8xVrFEfDlvv
aVCcVZ3ND0BhUX1IRoYxC7JmmrVDwSI3PlyDe/nbrf+rIehPZe+Dz4URlf2EAsyhhpBxOS5hamTi
0I7aTeZfaYwhqEGv9gOxhIX4iISWBvMvSmmkOJ8mld/H75KGvfw3GWKjRScQlmG+pjME3dD40Zjh
aNj080lq4HMc70L9TfHR/BBh6vwOYxI3/CazkVSGScMAfTXN65bohiwCnHqNAbg5mrPyq/UV+Pa2
B61W9PV/EfrpV6FCusMbzDHXjDnpjq4J96OY4m5uAu2vAJktq8PPQHUPa5xNMWRgzkvcRbt7j675
OAfqEDqZETqIrO0LVKoavyHWQN8tgfwHoMSb+pCXeLeeN46haaL7bKhZIO7e94WsKs8WQpDvTdIE
NXq9ROkAyUWxOL1s9bAMEx/s0w52GUA52rGyGsvMqkub98Tmjb7eY2rmwD+43fYRudJDHnf+Jxa8
3CyQPpOK5Oxf4AqFYdJ7LmKXKrSzg8mngcyrwG4VWAtcrmxNuhTYtbm4QnGvBtCx+dninjBtzhxo
bljhfcjStWKWyN7GKzCq7xJ1OmKZZdTwXHsEO6Aup6bGiRo0JcmCXUojMzNDKJxaXOVSBz4/fD7J
YIYpSpUGX00kekpHYrYc4zeNIY9y2owckdduCbGtnOQoXu06etPxwx3rzscIkYq+C5MRBABxAd5r
sa+sJrbiVtrA7YdUnMl4RAYMy0dbAxdjPCsEV3fTlbsy27XocieSynASjSNe4jINf8rNHW70IFDZ
pkNmiTRIzo59nbdnydoP3Sk5J+LijQ+KbOWOz6XpVqbLu3PFFNzCU5f5p4S6llr8U9IG3AwH+tAc
g68CKJLD+LiNO/Q4PBnGWwSXr8uPMaCsrpUvIOlE4w5UKvTYw/AjaE8Hm0WhQ8RiNMoZoLMFg9x7
UOmnZAmxI6d5j+DQ+CIw8jPezbGyhDc/Z7XvK0nAGlSGj0Oyk4ef0jX2L1gP0Vi364JtN2riX/lO
JgvyoiQq6d65ghgp6PzkJIkKVWku+gDgknuseWCXGV7YL0eK3GDRLoZIRdvKf5mh3i04GLMDClCn
Fm2Mix5MaqaT+0BSl04xG9nOM08/fUQqQeYGOBBQz7ByJc1ioQ3xubDax0GQgosFie3uhOV73kvI
S32Qjp4Sh+Gz1iw1XfjmUa5cOlv2OnwoKUR+13YFpgsjsi/dngGZUR9VM2Y7x1HgZWcyPuSOpeCa
HIo1Vx3h6WDCrH7QUOwWn5TksKLZEcj1duDYEd+p2Pd1h+JBESMvq1O7NLeN6kWW/1+iGRWalZ4P
PEuRK0YCBPbyC9bHl0rfg35BYKZR4EmC2aHAipk26BuWbUv83EqH59yRPClNOp3i+yh+/xU7AJVV
a2fWuGfXsxOrlCw0GouK8nAiLVP4GnpyWrH6V1dhBbQyaaCfZ1R7EL/BIECvRW9xs//NV60kkSc+
2sx5v0O88XoEo8zBCxGm3QJL5BfQCkmYxbMY13TQkltWqx+jivuVuzgljsMN3veT2vm7FXz52X/d
za5h8J291DG53Kvbs+u4K6PQxzLxmcq//uKEoUTZGCP+UmK1JmH6RxFhug1PMA0h7PwfA3GrEGLg
ancIte+GSvC5orUvAXlHte2+7KUZQHZ8VMRiUuVIYKu/fjAFYNuCrb/1T9XP03aKFzP2gZDLgwsG
+DybujDkW25h280IAnx/3iRf4pXWYO0HvLp6mNzhuQcVwW1OCTfgC5PVfQEmPfEiJrEP4HzEjREN
eFS3nvAsWL70eKMcNSt4pYtOe/M7zKouWLNGWz7jRQpbQLqtmjT8Gsu6+k2Re+tJEvXaVVo9c/la
tlmVsSz/XArdzZApCofs8bkiUMM/jFyhHfuhmuFdpCXy6Rtp+app1kZzCcM5GVPJtTL1DVy5dzED
s7ualzivoItBXNjPvp1uNnMKtLX7oktFVJJhyJ0fpi+S35PiKbfPDG5SLlJ4vB4E7zoVFGkCK1yp
SXCGDvQCRJvUNrNyk+FgUX3w+b6cuREumKrilmIYyPD68hiN/4DEPTxFCIYgimRZtvgXHFVjKvfL
SQeP1nwOTzuYpnWnd5k5pf3vxY96oF3iouh1UrDdeve68g51qd7dBjbqSwxYWcNKbhHoR7k78QXM
3CxLVwIwDsmi/He7Zqd1sbWwlP6SgZNGu+tNxT4s20wGJLFoq8S2dk7QAK22MpoAZyIBpWLLQCkn
Rrk92bzidMy9CEi+GWxT+16ARssHyny5SDrLjWsPfS98BZqsq7w5+Yzf/f2woCWYYmYBX9JSHObn
LOg0OcmUb72LAyqClyVGBHbbWzdPJ+sm+oJtNLAcmHTJ3gLcDSRlkkvJJbZIoHEhOw7Qr0EC40z2
UuTZrTqfNUDL4k3to6XU7nRngbxMlfTiTG1Bt8nKp8WJ6J5nAtYLRUV2jdrbBOLPGhwBh+0J6jya
BUoBRbLE84vbEhHhBdIgMwaNW9p/xvsUkGWqCerupw03yrRNDrHN4uWYELc8/yCtS9rEy5htg7bt
R7rzxtZnsAHsUUG34H/Se2bE14FbWsLQxCmxhSETWtnZjFZsyhEcn9CetDgE0udNVXQ0V6vi8CFe
BRA3eoQlKwWN/mfVDIN6ArsmacV/hw4UNVgj202c1kLJHEnodk+bms6vaBrn/7SteJPrInx/f1Zc
yJ7bzA/9/tmXZ/0qvmx44Wnv6IFdj61d6V3Yo+grPeAyySS1DTD7JmTdSMbd8rtvN4ikZnqle87p
pW4TW2IAZHiakeZpVH2QcdnaykNL9CGAS1X3o7I4oJ0GVqHnqSYA78U+Ye6qxba68+dOwm7gbVKN
BeQvnxPDO2KSBQ5czLpniwgDUugqlrZzej6PqybXDFeGfQDZhIbJas4W4W/EUV4gkX3oE2RI4yis
99cYWv651piU/FhuGOSUEcoMu6ysGvp+rUmbVX97Lc37qZpqm3BT5iwHYEfQpk2KEnvAVy9dpQ6X
HY1RM59hiSXLG06R6sfi4OkQBdjtfnY9MHniV9rBo9h+Nyon6S8MiBv22wmGq7ND7hO4Ad1ii+e0
WDfQI9mrFl1CaXMILMJyurqA4xC/KQPFaJ90CnO8h6+F7P2BRW/G3Xc/wGN6WT/X49LN/GCI05DN
P9cVguwsd4iSltBBzbku0wDq0ORqZBVKDRvhYzmgH4UU4uHuaCyieUK9HLJ56sRYlG0R8FkEVdPx
G8atSaoXaCf5fenASWXX9ILsxbh+Ilvwl+ubbsmU4C48ovbd2f2Cai9n35ahejY7T3SmQwrG9SV0
kAGFLIVwxCfytbESUHlUjf+Kntq+Jiwi9Egwv44PFGzIFBVqvhpkiczZxcla4D5l3Q62PEZqh2r3
SlGbEJC+1+xU1wdU2jtkK/b1O3C+iheTLmACFYDSW7773gcm9dArdx3EYrfi9IltBafOYjrlPkLG
kOJDbaPuWVpEUGHTg+AU/ObnlCTSSJuQavp+5Wxvjtlalu1IW1LudtRjGGoFbjruyUkhFwGHoeGg
CNJAT3jAaN4VOdVaofgW2xRsCISLeb3kO5PwhRQ0MIAg1djS8F2Coww3G8Ji/hrAfvUE18ANNQeb
W17SaSKTlBYy21eVqFMUXmVjRYnvFu7CKi+67hU9hHryb9tWErpeJTU5UHxne+Ai+NywmigFG2ux
QURUmXe+hLxD2rUt5sBMSUyaZ0B/SDIaUe2H+bjb4qBqE3NytIxSfpca7n3e79CIHOE7y86PCjld
X9hyFGM99YjqKEqK1kBHzP2uZDF4XdTj789YOKVFbeprQ+EVkCNeV1ST5GAW1t3VLXxP+8B9c3i7
BBcZQZrIpeVQv7BYpdwP3ARZO8uiGFjhI3SRxX8XhtrZQCqoo8TwbDQ0cxzmZZ7kLOCNJYi/cnvD
dFVHikJePcyzGiHC5iEgcSFinHsUdZ3UwO73adZ/s5BRWUNPRBePP1V51hAYZF+IhUV8qQ2u+Zwc
igz5c34TuN1mS83dJpeDa7OJtBkA0sOU3fi/WqgeSiTjuwnRsml3IcW5LlrQ/ipc2VqpPpqpVkrt
yiahFgaIyMIzaV0Wqhnxa6pQ7ot8hFd24Ab94uq3OW7pb3fnO06IQ36KH+G12mRyQHj/voM1dE/+
lZ1uQps9c65r4HE7gXWSsl9how+6s5GJXlHSNV4Luekm0ZPXsLCop1Y6CAfJsV8PXl4KPWWGqi73
IXWT90Yv+qyZbl08c5/FqmdVSZkuBkfq+VCyQ3Bg9WYABpsx3mqKCAWVLr2yXfXHQh7CDozhbrXu
FQ6R3VF8VZDcmXGG54gndz30MBIqArMiHvnUgXz6j2Ij3g0wAZLiZ83HKKkBXQSziLmv4dMP27Jn
GmKhAH+O29xW/sNzMNE1vjHXZt73IlEhGEUBVsB/AUKI4syORjoQTbRyosBJRxFT3kPl7Q046paQ
Wp6kRJT0pWjJZIrHhH0Ntel7WcYquu+w08f2C6Q24x+o0WAsqUoXc+C5qx2oqLNSMaFYqpFMWRZS
+XBGJF2Ls2qizvRlTD7yHJuw6I2LVlXVAL93nu4SGdU1KJNiwuwos2mvsfO0lVILtL83qIhrSQqJ
8ftOYE9KZtW/Ke3N9kbM+H0OxT9Nvo0E+iDMhgeEYs9z6NjtF/hSLa9engno8fZ3RQC06nKM6RqA
MGn5ID7QWRadvDMeeaa1d6kCcRFC2oBmGxgAx2UnXUbKYGVoAASFTonyoaEkL5ZvMsijGVyJPcud
vVe4hjRvXP9KTKK9C2PjUmr2Sf+Wbd3AG+S0qOQR7jxc6rej4CuRcEgTxwKVA2DIx9B5U7wC96XA
WkGjjabBH2VCNI54DtpbJF5teExgWZcrs1GYKGY5QVmJk1xhppDLyIAiVcdxLk90Mxepde356zra
C2kwTei/lugrllDxA2cGhT/EmcNgtToIIH1+TFporZYG3WQz3gBaS8jqa5tC6crrhrMwNpzZt+s5
UZn0eKGTFTMnkcT0Szky7L9wWKZEQ79wskLqWNTPxtHLlCqMnD/W6bt2yvcNkHXtIiDvzt6fxHSd
ykSTe+0aFAADPSkwWeZ2cGfsgWh2pwGaq1H1QaODgyocb9Bxinrwn3xspysObpw4LUTiew94vwvT
iZyg7i8OT5JX6ymEgm1opAoZdorJXpGxnoD9OH91IbxmASIliKF1wJFgqgJbmWZp90PMaTVrnwux
6b+9eGIVBKM73EM9/wtxLp9+cYAWsJs9/gKtceLh0Y1u2tRq48Fnh7wEWF1euUT+DHHkJ4z8WUum
OElrK5NaOIl2ojpjDlfYvKDtYgP83fCHhPLDtWQesns98x4HUibw69BA6SIW9YsidSLuyuEP+P+U
7KMbVcxIJ9UV/aWYaoK+G5zTDKGm3kkxlCh3uMd8tP5XS0Apx8gzcCTlAU/SW5ZZpTKFhVA6fGW6
sMN9TMJ2t1arLjr2gOWmVa/NMZrz4BGzKMSwSiPRAjlyxvShtlDsWG5RNRbgSnmNnsuoXfxtaOp8
zItyopoIvwRuWxfzH+ugk5+CbZoHtlHsjR1qYvs5MWxNOsDlT0PnTJoHfjYw4ryj2Tn6HkUM+x9A
ZF50zUi8L5BoeXDu0loomM5et7cFJKiJNM3+AvY52d2vK4iQ53bsyZpIInJTE7nT4mrxp8StrTQU
sn/bwtVj85QXSFZjdMYgyS/ylki6V3EF2W8SQ/ylQcAs2/g/Iolwxiy4FMrS0nwjryVzdEPiHXEG
fe9uk7+Uals3McTfiTNBLtlKtV5Yya2Vo/FLgPC+mepiZpdiHUsRZRHLm2wvUWAcE15VUgHFl2rV
kTVK62SJqhdF7Ue3Evs4h0e2unHHsGrJdp39e0+/kKMCqGMdlXYAJkBWE7ZjhA+4TxvR01Lpjpqk
57nBAutRS/tfET5cUymW+IsDMduYycb+4hP+zK+/1OBhk6GsiaDoeLU92SS7HZBneS2I9PKDpIYC
EyWtl+4nkr2k0vqMxtWNOS99cYmoqifedcA75WMpCekzkzKfML2wHGO7HHOXym6GHCFopoC8Zeal
M7oCJGuyT4vnd7UI+qaA3m8nEv0ivrlysTdRpXVbz+fcBmhFZPwF/1pW84HUI8bWqVW7kns7rVXM
aN1T3z9aGPKag/hmv0pgvcPs0f3rU/lPybdRI+jRoQccA4yjZeLokqbL1j4PA0Zo2YTnfwwmlj3l
38iNgj9IQYcF0gX8MP4/y8nLrPDs1VZqQCnOe0wAP3qXG3owwbf9N8iAPBZClMz9DAdL3kYXnFFQ
/1+P9Sr+XOk/QXkV2fMnHrCtLi8GnDc5fMsa8ZbOun+biPK/YrTjEC6cEAegDstLlvnUV3TUvMjc
Lk5xi45ksJgR6D8RQy2Qz2POlVfu3jMvz8TWa5b0RVlEo9zxvFveSulP24nGYvM6I1zWJvYVnmh+
lrrfZX92190vilfH0dQJf4xdZs2q4B0/DiLuDx+ffsKma0XxTFxn6V6xFsf/qF3up1wStXZojHUY
KRTR60qtImEQbf2ElkTp1Ok+wkZkNYYjYaxJpyFhfONhFbLDfN45MCtmZS6cRsXGb9HpMnMbAHIQ
Q6F2qQfpDaPXuh8gawDS9nB4vu9BiLIo4fGl7aQARW1utJ3xhd45j0UyuLyYrv+zBYFXYEsnGnJs
om5zK6QwVsagBSeFJ/dbYJ3hEc36ZpUQalfbcW2K0zRL0TiLkG8VRxlqTmK+FzTFEDE3J4kvEi9A
TppWaHevAKUWn8munA8npUg2GMqjRT0svnbVkmPfKp7DK1JwC75egGaQ+SUvOPf8iQUuSP/42Mv5
UCQ2vZ2Fg+NXy4vuiPYvDk2bFdA/3xDkTeqDdmzQrhuI91En9kRxWka+IYNpdczkVbW1uISwm7XI
1goTON8qXoAbq2J4/s7zPkqK54edBkwY910ykCBsspiL/kMK+0jnnVADwzWhEvWr3ueQEylEmDdz
0hQXKIt5zMqZibGKMWt9/kkHRpxAOQ9Npdm1CJZkX8fgiEhq+o2ePfruPIPAeIHntahbKEhBmeHV
aT4voQVDKImshZKvxiYzQ0cZ4cM7r1+C+XBxfK9TcfFXQo8ONU0QjR4QzhYhy32rrd2Uos0scJMf
1xXy+Bx4HU2xbHfyZIWyZ/eOMAKkngQt7sxSDAADllnXnS4sdodx01qfZkp080cJJui50PbK1NZA
RaO59cNyM+zEArDQqZPXGL2rYUlMRpQHRfwnf5hlaI19Wej4efAztndlVJCfrMPRI/NnOPpd0Aeq
O+7NPpcTmThQnp/DKAK3vjWhLj6f2i+Wbv3n2UcQBFpxXzJbUUzefRYLjkrr0Qr58+FLCZIxC3cH
1kmkAWDA7ZzM1Y3FTouWmEhnStFW1mq/u0O5v5X1QeQrGYxqY5Zqot0deZJyEvNsfdro5p9ty9Sp
iukDX9DtOdN/2dGSKuxPVFVtOiG4XOEjSfwTEPlYPDgsoCwSpXlG2jJPvET45J7E8MD2uNVzXJnQ
US4wT1wQ3ZceTE9JvDVQj/E4RZDkbYeMpoS1HfsJIRcLYiAQqFHLC6AI4ZttYe2wseLJMwf1FMqM
lFMJnRcvEiJIQDuvG//Gt+7F20bS7Hf3HixkwGnWHylFEdZl39lD+YFUAzWGT9aBY0+7/2IygNQ9
y9VEgPAY+icttZJ4dO2TEyEcd22o6jYexDhlkTgHJtTanw+PG2ROrGjq5/cCvZJt1WusjcAAcNKF
I2MzHmchoTL/cEDbjdsITk7cTSgOZaiqMerNrSlq8ixUM8qCi+FZLd/nd+YkFa/nEu3YysVqBgGg
pGWxB8uw2Edzqq9OZ7kSznPEBnS5/AbCHQyrsIdzkD4Zakj5kxYkcD+ta+JLRFCGEXZG0GB7rssF
4EwszqwVXugBnh47vEy1XyfVkBnbKcCE4ykjWM6l/tvaCAwV6BebMesCgIW1obDDtdd458bfq1Ah
effRUVerQu6dYSFfbSJvnclfBF3uckt80V3yMF/B2w/ULNkKgxRx4WxJjIsWday/qqviYRNiP/ho
Zl/9ZflQlzyZtbz7fOWebKCnGhhEDWzG4XmHNN26rFBLzO6+foz+UxGf28XLQBFhks1p89SWCcRv
+hdcAk+OhRZxp3JX+Ws6ZPdEVZU23k/jZwHOb8P7eqHtJW/N4ElRiQOaOczohfDgwzUSLZT5b3iI
IxXeRWUCQf7VK09fyPNLRX3MvPUSYGBsAB2WLu83TWBZPtIFokW6o8UyCnMc84iWX9TglUGgj4Na
ENW5bT2aUn1xB9bp/4TLuMUaR6S7ZlVfHBv/uOJCINGoF0+kP0YkOp8C+ZYNFdk/WpSCeEgKJpJo
vY0S8HrJSpD4JZnIlF/+yynokAowOy1pY3xSr5BAnVkHndxrsNsYBCb9UR5/FaBZJCsr5AfSHjl4
ptkIwirqb+dAjNjdqrSFynbHfD/s2GYUBXeGLJiGREQm3drBTfodXAi+wpXjMoSO0lFIdKtDWSQ0
CdDU06wtCIIUREqQdrBc1XMiDP10YW99vxhUOQkkRa2nl7HnxBaDg7fW+TQ0WuHX5f1EWlT1p5o8
vk1U3T9Hm5WKFV+u/LH63Qoss2IV/Z5DkJYIsZpR6NYlDHnFfmxfQrXekPd1a8kPQRAHMtgSs+lc
8hLYGe+ANvCGEKWbCJFI7um9d7QBnmohajwUlo3pLCMeGqN34FWTcwMYboQaQi28WJkWRYp0mW1C
x5xKjG1gzjCQhd5vaqtLUCjsmfba/wHVN84VQ32n8qV1W+uQ5Ree4APdCSk/WzijTBq19vF8HJYH
WB2lR4EGC8M2u++M1LMRYxDZNnSUGqnMI8O8eqwEMr5rNJc8Q7TqvVUPgOy9RYfuuoLp3baJQidI
X9zzVu372PXukhB4PMgVeG8obdCgTLiBqDkYYDn9mXnk5d8so75CwYNhhFg2vH39bdl/AxVdw0bg
YPjC4Nt7XXT8j59HZPd1JWTZtmO1D4G/iDGuNpqtV8ijLF4LQj1OFlQSt8YJvKGI2zZsWp4dj4bH
0gQg/qVTRW/5Js9ttYL9/UKicjqeqSa1SAsGHRi5NZCDmFe+qLL5XM5kqVkaEZfj5AeqwS/gTmPm
4tzvbsLDneeutt3jXFjKDVQZVi6v++JYMGP2l5okbEM7yA9VfhYivqiUqh6tJmfPXsgxMOHZMUsI
OQjj9L3X/b2/PoVwtwzSo5/YMUS/A/Wx9d1QoIgC0VMNbeMw1MTzqfk7PAhVdk61UrH+MT//q0zH
FU1Puf9NHvnneu8JJQVFwMPiU094Hvc19Qh0LN6idz5L8kaPGErAxupKNHcEKgrPxXUNp6/PDU7g
g8SZn+TD6dylkzdNj2kTEi4aZtTjLd4oKra6uNfmgIUotS/5FsF1XgZM6XrD3MVhYQD6CgBjapHn
eIW7/73XVmOQO1ju6+OMfMRpLjDBiJuqQ7USOr5kOGVtPiQfCxIDiK24JjEnAxy4GZoQTr33J2nl
IiF16+UBPi4DPOr2YbQZigO1y4h5kuCaGgjOn35epI7pSqbSkIocnOGvKvwtFHNJfAa8kQ9AwyyV
GXhNXUO84YtBBGD0epfNmNK+JevKsxPWN8rmQQul2dhioztdt74ic5rdQWuEAUNiedaacbnIRVQz
NAECeR8jnLMnZnPd+B7YXMJeBJtQkT4bRM65hFX+YXrelSuQNpCLtJu3ID1I8kj9okKpKEk7GJi+
IRjTHgyc9YkHlwJ/WC8Dnkt4WMv2Wc2aNTMYRrogOkRe6RSf3WNvQ1nfoinTM2sMqPjfBC9qehow
kvEU7qKjt/C8cwlp7PpbJV1qhOVl+5G4+8MIlFDP6sWUGEOWUHKwgSXR0hyRqKg5rcpuw/Zo7Lu+
D7c+n8R3VZsMEMjjmTE/QrTpUz9i4u5oAZjR03QIl8IH8dPgti76IspA27LMVdoTY+TkwY7+TNPf
rn8pibwbtG+cyvOMuzNAuD4Kisbq3EAmiYbxS0zTGgJ11JkzDCkwDg8OYpZ8Y9eH4yTgEaPfFzIc
0yPEDTZsxyFh5tTii50lRINRkroD7cakRgr0R8lI1V4E6Z9PzCAVPjD/JPA3jWfQecQekq5kxpwM
jbkOn8atVBD6QcmqlTLMGcnLqvS0tOS/DxqrLEpySgeCz3YqAaKFHbFVClRJusIFsIECZ0a0aIXt
O3Orzoh0iXo9iVNPJZzXBH1Z/7NDbtFYYhjiX/TbT7qsOj1ia4lWro59+f/HCHdxrgCifdtYMiHs
gCfmnA5ByH9PG7SurzEc0RNkE5KemuWtwGcJZeTq+rzNfAQO/m4lw1xsLShEmHmxqgONUIYAMrjW
bnx/YHLJac13xpKXSW4LJSM+sz9NJZ2MGkDuEi5N3I6FjwzyjgZaNcR7ye45ihQlDYjeUzuom3U9
JsW39WbHT6rDCcWvkcQ+d6mV4mlraraW1czEb3uMA/EfOVYXT81kGm2JtpoI+q0fBCvTt6LfqjsL
4Pa/Z7vpcuFwIMZbj/cu/Uuuziijw7RyvhLvKNjAZ8wQ+zuBZ/J7mrgOYSJeoIsYYr1fr+hjhAdX
uAwI3DXy2AzdOfsIvI3YSiyue6q66hr12YSqxdN4Pbhyekh4UJt/YMIufsaK9DRQMvWHkfYhKlXV
noTpIsBjC0mzgdXf3Z5q0Ii7tFzYy+WRpM4guNeRsyxShatRuytsoRZHMLlO+JA1E+Ockq9FtDlN
17BIHY5BSn9/RvFOnVLFxxV19rYPxzCRUdC3hbjnmdTABLO8+69FKGnaSop7wK9//7SwB/M4xUs0
V58KUisNB6gtSh/kjLpsOGK9Acydbv41P+SbHyYW+BmnyaKmGkuqsZMcTMt0GfHiREtaW18BDAhc
wW6GIi9G/X/5jvaq414IxbKNj5g9gV3OQa5ItRHHu3iiicpOpk3tfm6OrSgDd7zdiFPBDnLN2OwR
OL/VxkBJR7nkjpsvJbsrMIJkbZoS794ll+REC+2QDH5/t0BMOMdUzQHV9Ebk2Bvr/A+gFASX/sse
ba7F3pt0TjkVh7pNVkAACsqBTVXSox+MglVgPE21CFPiq/f6o9GEOvV9ewe9Vr6L8gQgMNq/UWis
fCflVFovCJ9ZlO+00uwdSpCW1nWyRbN0EM3CEWwvVXtI9U3Fw/FD+RUolW3GfktmSCF/CxgTOtU7
Ur79HZ/NkrXSkrc5ajckXjFGbH7T9guzp22Sc7hQltxF22h1tMHdqwp+H7nKhe0CMNvHyDtK32xx
hDeXahkx+xiCuQbzBk86YqbTWUPDdI2aApSEWM4gDbTuAkGNhKRAPG7C2L9fDiXsLi3WBfIMxTFt
SCdwEn9S+WwBFIDq/86ue8U65y3l5952zOqCy0NW6KH0LI4fvGubn6GcpJHMuHCaezMRX+aMgHqq
0rQm6nad+wzO0xgbUml9FWC5T+o0f3Bse79Sgz4jjmgY81Cux/XLsdwQm2RR+hHm9bzNydUDEim+
9T6SoRx6bFH47o3vKUP0OXmN7ECEXoSD1GACCJPQ0HhFLkNzwIQf36ucMHyN1xu6ak8ebHPnddfZ
NpL/PXA6aat92M4OsXMfD5ZfwffpzaHDeBC1e19DiaXMI46dXk/YdorUhCq2/0Yz57WqFJgog7vR
4lXul4dT9Vzs+HPG2BL2tn75hIK1tV7ClqDyHaheOUyFio4jY7UPdu9RH6dTT89/Baub4nYsUGbn
iDOn3Nd5dXa8d0GRtLgGq5xEeaRZUYBxMZmxRV/+zl/qaLQ6L4CwRUKCT2EJGCb94qZxNpBQKpn9
RXQj613L2WvjTy8lLI+FGtGzG8SLGJ75R/sgDUy5USuQec62UT7cgsp9mBjUlWVS+4Mzm/RRLhl1
UBQ5ikoD8HRKFgwa1XArrd41b/TySe40f/WyqLoqbv8ziGCnkD0S1YDvzeIKt4idcCpDScoN6YHv
WsfBisS5byVsMNKYkdwwybIfafjs4mBQxQnczbm/9vfFU0LIV5IiQsBghLQGLLLoEBogTpcfJKJM
e8dVmaRs1KquyreJmcqdS4qVMmksLD7akpSp5xR4I2RUqUHuEQE+0nPynFbDi5YtVNxTEw5ZhsUZ
CBoO8gz862zcVQc1x9W2EbrK9Jsgx0YpWx9Xrxnpl6z+4RGqme45bKxzSNlfI7GjXe58wL6S1pz4
d7Gk0E6ZVDCdCZQk6KyBfm1UFwGQqPYhi1qdL9pMR/hYJQEgKomfx5OOd4/SRqklLqTfjKYWdBQ3
Gbivu1kX3dngo/gFyl+E+uDC8+XUezHwm0Ta42GCzLJ/OMidLJFMLGK6pZfuWel4gQ4fQYKtJTOo
3oB0LuAaC/b08lnr9680uxW+ZeW1tyQU9caKLMEi8WgYZ+ziTrp1/a165udATU99fLfLCboraG+K
398aLFSea6P2oDO+6bg5eODOff2fF7XkKXyFEsfJ1QbcRpCJR9co9TCxQI6BpT2rKUf9jn7XH2Ba
O5JmSAK7ETM9FIbvkz3m4NzkP722BDHiKn6EpwavuM6u9FCIRPYu7YCpDFaw5MwdaAg6MGhqXC83
sCpKI2ehqUmW9HkqlfRtp8ukKo2QqwHOToOu9z4fkdnVCMpdlFe/waasoOyuTJSsbrCPxRsMQD+C
CseyN7tLFWsPqZtAH2FtmMVLM8J2skwn1noeORyGws3e3zXyth9+J376Z8eBihTfgxr2NE2fVhU+
jfYSWHzQNIH3houwXUA2xTLWfYGSWQfuvI7wP2aHsbcXcG/6t9RveFMXh+vUVOwRTDgv314D9q+D
mt8li7sHWucMYVTSticOhL2pBP58ZzjX4JOcuyQQJsdC91OCCWiEr8vjJVUsAHe8LBSrMcWw5NCH
ESnb0pkLa9a0/QgoLZIxyK3fM/2CyBfidvU3gUYInNMM6aKLnwYkODxmRxIHmgvxVJsR5pOMXt0y
GW3HXvoB2RRXrK0qtELgrbTeidiwBom60i2DrD4sEinlL9n/5FSHj/S5kb7mdQsvLjiqXsdinfWE
WIw4irL/+15Og+ydR/oNr5m6sLh/1j68cl7aRwDtALzf7dGLHe9wYDH+nAcF7EmfXh7DEuYsFElu
XBFh1sm7n2Av7HFVoDdN3OJww3oEsizldCdLivneRy/kYN1d3puvAbxFi0vvYKTUNJHuyLdj3xvs
jXKk8zf5a8SqSok03xwj9s7QfiAXgfe037Rcg3DTV+VlASvRwCJR6TJOlk+ekSu971OgZpBmauWm
WRIMKz68SCqzjb5f7VgfQKu3OjvYoByILMbm6lXIVncJx9YEw/7K3jGpO5XVw9r/9cLPVycX0vU2
EBQ15xI38So0+Md3hnKAySQNb/0/3Syuff/gWd6b96wt2HzWIVhDLUe1HuX9L1q6zhGW8WKWB8Bs
Jt7dSeHDWQTsikjqQTverxNxU+5RDj423fCXheX69FaHu7M1utBboK3vQyBtk45QUTAqerqdIj5u
NDRAhOpwNUzGrCO2paeEzgq4jF61ZjXr9ufNNZgS4Ji+dPcNX0VaLtiKLLCRXftAxXds46r3aPud
FIXLfQ6+2CfTlWI7RwpR0OAikQc0bizJphT/Cvz4MEaxCsGcXkGV86hvcCfjtgUx4SIUQIWQtdOR
EnOTBoYtYCVwso21KgylZf+IDSJeLtI5PBhK1iYjfpFjmURxKfqlKDb5Yd+BXU7sffjC3XeX9PnY
e2oZEPGAezroQ71q4UjrBpAAy4bsqCqQtlxSdidSuWbJzv68q/mm2UDxbpdNqLNEZQue46dwrKay
RurKRhguYnjjxSYmCCx27/f5twPYBtuE6REJCzhdubDz0AW1sECNURUKYopCjafs74/25o6wVZYf
aNV27oV7DH0Ay6tpIMFbe7vUFBCM+ji7yCQl9qvi7ROhqwB/oSg+6mmY8ssc5tESWMkyKMRfVXPD
YYQSg0FykF7ULAu8ou2kxXKQ78QDzzlCb5aDfK49QndlSxSDPoVFA4Cjl8quwSOdkOPelt+qoUKS
Ka2WwJ6BmpdxyLwKCx6LgA92p0cDb8MzfobxWsNiHfmf2lPO5K++xqqmbF62+s8iQfzG3+mzbPZS
jFZI4zGknFURX+5AZEIOJqhYj8KOCbCEXifT+gAMBKm7gE7iH5CnxXTvZprwNXR3EeFNlfVyk6NQ
PmzK6NZmItKN/D5i+Hn5AEdKXYolnx1KEVlgt3YTInDTck36cvpS5Vldtar6yFY9wHzaQ/wJ0uV+
VWz7+szNnOnR2kNZz7PQiKV3z2uQMU48wkP+7H1fTF+VuAJ61Bty0NlMVIrv33i9bNObI21/RpbF
VSKCPM1WwML69hTedyUPRcFAbqwISTibkFjw5p2aJH4W/8CT/r8KLAj4WxvYOzlPZvyMkCVRQ04z
ghxEvAnFQtZ/rx4IGvNkJVNMXDP87cwit99O8xn2+Zxtn1wlPoRq3BqTzhAKtWPDl8TB78h5f3s2
JUU/t3TNd8Wzc1a0/6MNlyTLAoPv0/R6G3ivnbJEjZC8vU18oIpSwyTAmeiBel3PYrAkiGvAUugN
CtcfWdNcsziaV91fYybbE+xqtbVbFIEfnPUAqTkDPQZkQA+TatsPh9riPveCVcdErDPxq+QgKiT6
xkk5MURq3bTNWQSEO/Pk6sYsOGPPs6zuMhs2c5U+KecnoS2Man/U0D9SU/3mEk1dqDHEhiXNeGlF
X9Sga8aRONyTVupXqIk9g/dsqeijHVCGjGRYauepZYKozfU7D3tJio91MbFEPZFlEWPXTau9Lopq
lPSSLVPlXcvjBMqeTr/aEG4HMDAptaIKiAAH8ZOFwVrWUIrTBat3yORPCPnujWWylYvmARpf1f/f
9iVacOFk+z38p5t9jeqpH7xBjG9GlmOEXZx04yWE3ScWHdxHxKXSgpV+Z5GI4TTNTl24stKlZ3GP
soL/GCkCKrWn6u6tdQFZFgA5wTff+l5jeEnH8pNafXbon1nnxNl+xuwlIOXnFrNeBlPdbgj5fdkm
d7QKsCG9cJENPNxQyL4bOaGGGjsW3z/swEHTkKSscidSczG8oSFC+2f2oW5jNyC/FWjHD/Af2tZI
EwblrKYpf/EUEa3QGkQxlw1cuyk2JQl8UHj5+SzwacckgVPkm0smTh+oGIM+JTeyZtbwIAL1ajk8
vRow4PRkklEkLS3GvxB7fjdiilRd4Ynu/mVB31nf9VeBLBORkG2bYL5/fHVsOEYrWZGAWjPOnZpd
lD8dHXF2wiUmbCeAB9guNt0tvkUCLvVs+bEiT4YNNJZ8H64EnCPArtdWymWkPpLnEwMaWrSq5cah
n3nN62kEYT99K+pOGr020p25QBC3ChGf03CUT0VG9uXhnGf2+ftmvzyeREmF+fJRJSP15/tChQSc
3gSvHBv6OMkOA1qbcdh6KTrpHXiclh6NKLWFIglcYmNzFjXWekO/JPkO29Gezcg7Zc5f4XawxLGf
W5e+u1fiM9I7TiCPNovUTOVAy0qbqZq3bkL011SFPfckNlnyhuVN0Q8i3i6UIEhVyLgoNMughHU8
YjMTl0rk3qDALsvVId3hyqy2pdmzYOWwfhBp8jXSJ20a132Y2XyP/pv5v1/rEJp9OIKZc+Nf5YvQ
ElpJpMzbE/FHUWoo0PhSOZJf/AkFuPKG2g7WWblplJaTaABM7IrN4UP+1EbljaVG7b4As9WWmrEx
lYcVdkRnQTTCmX5pIBhj9BOqnJm8LXFXkksOL6kYESE5iIA796qDlVIR8zmC824SdmONxK6+M5U4
zl5G4PHfA0lnF+crhOS5V10vQsjjuX6sDZ3quYt5MniFpSm/lGWcST9vrenxQYfo42cPcwpra7oB
kpJdhPJHWA6aeThyz/ypj0/2xeT441sxcpp+HjzT1p5xcqs2Ad2DazivnA9pHGUtIs9Q5y8yQH77
rpVV9IwvVCSKvSfci+QVf8QpniFHYLZ8vGJM91e7+Kbd8RrNPt44BHkSnTm9BW/ydYNYMs4BbAww
qQXGEM8vVcaiPC4wRpqbqDL1+yXa4yQsnuC8Kamwr55W9UZSQvSkL9X2rEd+3wWKWJuTTEF9g8jB
1ExbAnPyxLNJwe/lz0SYbFQH2bBYTUBfpPDS3XQtxkoIAFcrrNRtEYufMORrHlrBrD5DyxHh00gg
2IygSf7HM+ulubKbDcL+XbrnL7yer7bHloNwBp6QIP7aRBKua8YaEQBW6ZZl8KOAhtAVcuHqFXY/
BkCNscPcaBe8MtJz8L9e33cv/XDmD/n8HdES81BDEaW7FRmNci6jYspETaLABzWvjHonzbUvCdAn
AXyhiCDFow2LBqcth54iRxtR1VGh3iDyf1gqx3tGCL2grUgiKdCgpKYqEFGKof64VxPsTU3Ev8M0
iNhKOut9wGNWR1D1EZj8stz4FQFseAfj6gGSENGFT1h405VcWCgl+uFpPFxeuVyPTxygU4RSrxjr
5xj5ty5vfN0GOMpPay0IR5TrrselZeBFV2v6CkDlUkz8K3IJptKfYyiDTjhDodqxT6tPqMHsDhig
GWliTimITi9Z20gdw7xoiZkLbcTovgYmP8KHDK3Kx9lqYgdJckbCd/bFXvszLmlTR2HNa7qNPE21
51+bMcUD+/RfF9uf737BrVhiye76C9iEdCvoKsvTMKlkBPBQPiqOIbf8K3zGTgA3/NnbDXAX2MIM
c4aYPGJypXBbbRYvE9eowG1slvfTMKiaVc1G9D6sqXdsK5KFralSIvo5G4fsklHQEEG8sNwyrBvY
3KIgR1WUxEVaPYMq8McIlENbJ9iAhYwFON4zi36C10ALPwXgkraCwWEV80QGKbOHU+Gp5UVq+bPj
dhVNshdriaQCyP5DSr69KIgqFlaQBl6CS0YVAF3urFd+YGUJBskvS+mXzDkvcP3TWQ5M6Ho3bMEj
RBONStg+jNT11Ok+XARg9BQF4x5DfMblGnnpK4bmKCNdXSJFAffDN2wkVego5uP6LedCcreZ4CPV
R4k6xBU+JhBUZxExk1JnKNNGUAWx9HOrMh5lAa2j/sl0NkCJL8bN7dIgCUe02rZB/DmEYxsnJywk
U+0im7iykqCKE4KruVRuz58HeunVulXTiHWqXXZH5AVFKSw+Z3Rtwyh+vYE+zYebVcwuhrwQv1eY
wiqxahrWbdBDbiahJVsL66CBU9k1bF46F7U5KoIxAbmJwiYkpE9poQni2ZJi9fLWocsLtxM07FmG
/omdv6/rb9jXzYtpin5nelftFqR8/xA3uWBWo2Tq98vdb+AocnOqyM4uP7IuQ1eYQ39P/HJN2+PW
qWpGiqh25FmzRUojvGfy4Y3BuIDSTwfQfsXMflvFfwZzP/nnBtSVnHlHZaaFS9iZq5HvalZCo0gN
j5XdDUC8k4XAOJ18LqFHR6CDJIhU5JIMMXA7+LNiSfRE4rmjZEUBkW/2PFwC6kj18zbazZzdfVvR
3MDh5KdH0MQEpV97aBKzyls7bE+Dkgbz0tJOHA2hVBuQdHSDdpy/SMCoRnjN8Xvffg6N6oLDFjaR
e35KjykJzIeKAEN6xFlIU+9iQUZAFwvxUCZ3Pob1Wqwf+4frj3TJBtWGiHAIt9ErmZOUCNA1NmTA
d2ujD2UVZdZtzwtbFRpk515EjtRypv3PIbLNo9UWsymG3bfTgyxLhlRJc4ffcpE2T4Lb2FSy8xdi
4YSqylxIEB/TUMx4jjWEgOzBvRclXi+fVWMp4cARdOCCGG5wpGgzgUFzHHPnJnhrdCGdwvUyaVIH
GEMTDvZqhra92z5WQv5jDHCFUGVv+KBSRORilhuUo7K/FebUBvHLyInRR3qnmU/eH4O2d0BB1tYV
JLrhkee/msmqyFY8lV1I1aM3T0HqnySoYUe6xViF8M9hRp3huQzvohGiXBDVjG27ajEuv9er22yH
2FRH1TbOi/M+RIpC0pjhpkRUhGIuy9WQOEi87TauGwyXYG42lRzVBIxzhUrRowa3RMp317Y64+dw
P+mdwM+hds88DBgfIhNJiism9AnxPA91tcjLwbwi/V+fyH0LuUkjGSL6yW6Juv+lKNwbEpJF0Tp0
HpISf6WgAT5ozIlFp3w+9/Ag/uA99R8vBYilYZsklBWR+qgS8Vm71DI5W0ja8zrSxrUkROnbj/8H
4zb9PS5rQobeT8dOXw0vzw5CsO8ns4POdD+/OQSbQHY2VrAMixp732ziaIC8oCiM1gBo/b77kXpi
kpFmnIQ8SMA6Hj5Qf2AfAbkYHJ1Z8Eyvuj7POOqL/O482g+q+HT4CbrXPBOa7sri53j2ZE29p7jV
rSyq8Lf4Yt/XF332Dk6Bs697uEK5LpS5elEBY9h0zfDRhmODBmnwh/rYrihXEKSGI5V5UsNXzMzX
m0yNJ/CTuazYnZthht4Y+WIAM58WhYQSEqErioJi97DU0Gj/ccsAaNBCeCMknaWBoDBZ4b0OIAbv
9viOzJRlVTuHJIgCiQrG1K0lPIcgeHl1j7MylxmeHHQZ+dzULUaT9OtVBRzqSRxzi+yJ4vFs82qb
NZCpTnbuMdWh1uadv5wilplE1OnZTrOJLyb91LD2QpMe2sv1N4U48fpqfUtPb4CKPRPzyaskYJcx
8xJaqlIdRgvcXvVGzNlrlGrDzxfWEqM7DwMXNnsdm6SRdgvVcHkWFr9gU4yyp1EW7886lDYsDXXv
6YUAvL/VYgSILTSdAtUBZ5Y1lGjrjktjXZXeeiijJ03AMUbCcaBv9FF5w1lb+dCI1//yK1AvTBg/
VbJfVRMOHwjgQtUp6d7tur2xaIZRujAfiEeU2iKb+Rx2kHlRIEDmAHwm7pPeopryjFQcL4K0OJC+
jaoPY0+16hME3FMGmSNwVE6kYQmFGY2hDVYr1NXrzvGiIgb8vU0t6+pHSfu3uihYR0wIo8SD4KMN
aho4OUYz2gdId6scfmz8mb3NGkAA/jCZSysv7z68s1y5cFcJyn1JzcGQ5hzubCmMYnuVKOjiDVkk
/HcaHC98A8a/E4w/WT758sUB50+MKvFd+trvwLWnVVYFDQ6meRrzS5Be1ei3413OG141oXeD6m/8
+nrzHAvcXW4FoR/42si66gwmNXgcO7bVHTrmxvg1eowGDUF2t6JcLYNY9K1oAaBTll3aomoOyJtz
4iuGQ/LanQ32XMC31Mrdp2DRkfl9KtMIU30WnjNvJNM2E0lljq5KJx1OpDOMnGBRQUWT+e+Ltfvh
7/iFs7gmC90QRAWzgrVQegl96VPuly9/vO9mjrk+VHIPDsGggeqBMJDwsXLoOAi49ycC1z5pa3Dn
8LbDpLXUvhLeSIlDmBNcT5rxkO4s8tUtZuEhbEAFFGEFGC4GqR1+wBKwCEDwGC3ZmKlkkkTKF3SE
7InJaNEukQdiLyI2HjJulop7LFq1sH3+1I84e7o/rO2zNhf0KRYjDhaVQgAwxTxyX0uOVz2yH6Sw
5zrSDx7QloiA/jPMzgQZtTlCXIleR2qqK3uLZv9mLhB9kw+I6DmyMkvw/fzVLV1SdNdBzY9Dckpg
sFyVZsYyp+e/NFMmx7FpWVRdgYsJY/HPb6F73IfUc/l6jeFmJjukDBlhOMrgmGRKpAXrZ8GNwQlT
jQ7dXfeRX3A3kxxXs5RjjJkWE7RyHVsfnGviopP/+QtQSJ1fT14nNlNSe34dtYoZQN9WN9FGTrsm
2OcB4YlqgH9vRvbW8RcMdFjtLMOOvD/19HDhL5GxZi9beZ8IixGswOSIsUURrdGj0zFXnZbrMqvK
jYi88ZpgpkVK0xQFQy1vaSYe99hevILq3j4JvSu7eGBbvsp0luGuswPELiEkZ0BQDldegSDgz9vP
MZDIQmnaisr+U3Vs0EW11iVKu4sRNoE0r0etbqz6W6ctNH6B9o/gGjuH9a7lVwYG5nhwzeQwXjaL
kJ/ZRG3xLB7XoyBdQEL34eXBlvg6LLEdnHwBeiFStXhV6urrdTsLECYO2MvUMT6KB/0+zwXs8uwt
wnGRzvnAC5Oli9AT80gH5AXOffD84p8aDJj84dTJY9C1aB3B6Sl/a4KgRXzEA0mHK9wQA4aLNHFm
/4ogagLkhYZT5fXTgq0XOPCgtReNP+23NuWjWF4rts2PPrjOM8WKVFrg4l3XZlDRNuAVhrxGX+ZZ
SY+R9M09XN3E9Th6szGlRtRngdVGk5ZfU3tkGbDwPw4EejkeMKfhKW7j/DPI11QHZKvIo4NZJdNH
xmsTeYQbEH1i+04mUk6dTJEuc8P9/JiArsyuVCwQ8QcDNO6MV6iY4Sh6wlfuJVzORlcsfA3hNcIC
iHKISdk8kQ34Ylbvagkr+CSpy2yquhIxRnl5JZUL9a5EQpxL3Yf0y6n00eEc4Bstf8AjJQ4D4XuK
87cumJvpdGPKoRd1ysMQuJ9pX5YX6IOUi5ztY54kp02diODLZp0GthvG0D7D+U4P6BOqERW73eM1
xttfDoxASWFA0GM/RIuvrQBxAJomhdrvUmtDm+rVzT6XM+2SJ/sW8R3rScNCZkDon8t2VNrReQVs
iui7tdpB1wgMUw4fS2U5lEBEge/7MOVgh06Ne9QmUaM9aEIJSdv6g+aA86FPbiUevLHQ3yhbfI8a
QSpd1b3yJ0PO5CqouUyUG+z+1/IT2sDHSeIzOLVj19JoyhEjGJPA8rzD+z829D2U+n821XwbZiLb
BK5/y6UXJbDWKn0WKekdg9k1KuuqrpRxy2WCR9rg8WhLFd8tIaBDR26bSgctvOzy5EUVmPLB6ZBw
7ZMxUvOQMl8H/Mk+xDy2mxJY+UROoSNe2b1jm6W5ttH4otnBYTFTlurBdGPs7XIAtrScAANAMKdo
2PhGzpSUecMTgp+yOSTjO8rAmaADx7ghZbqApxZ43u6DImgOg4jyz0kitcjm7qeqt+w8MlAC/lg2
mhtG/4+dJ75kjOUXH/FVB5Ri9yXBWfcAqYUH36wRinnRTWvAlCpEh9GsAI7YH6Wgmyp6ExTbfJk3
k246r5VjG4MpkhQxpPl717F5YXIqK4M44B/9PJD1Z9Je063Abkd5G+o4QgnbLhNGgKXCTlAjzPYL
Hjlp1BB3Xnw9dpD3kPC+8V6190ZJPM+WMMhlFpmHc4/smh54bDbwAnddgNJe9iKV1V/EKLVYFmXa
I11hitCXvisPWmvGtc3+YfO/rvrcfjjiAdPt0myvNgbxvVbmH/F7TUY7hmOxoXlCDgx6Fiw8DwSQ
7O4D5Khj9WTDInNrz2ycb1ifCE+t9S8M0ZXwXQyDQyUlW2DLoPF3J3BU62N92MhMZTwpX1R8kmFt
UgLL1iUGkq095bElG8twrMBfWk6SUvcV4FwiaanSz1VdO+o13K3qgnYXdgQRZPrB7JH+wZhk1UNx
oXWo6YUn03jUMmrih8TnieAnvtyGKtqYS60QbKQYjbXbBh5IdpZjofS+0MlOSO/tstmYwq9w2eU1
ExUbGLyX2N527stS+rPVZe6SYZHOS9Xph2X73QeFicTpN0zyP9l06JvFpsAs/y2fjoOLBnz4TGdQ
yXAzNXzv0VFcU8QFFId7J1bqEDPy40bnaCx6X1M/eeU5izsL027bsTweAAIF2hakw7KI/KhRZL/P
nQmSDg5Esn+Stnqk3XvcnRzi6u7mdZHpk9g6kJfIyQgn5Xx8O2GYMP3FwVX+hWoxGwRNxrf8/Haq
pEMViqzxYTX+Q62wxmQB4RBlvM3KwkYq/bNtgCppTWQ8ILyTFLxE/ufL5QDRTGWAdhB+LHTa4134
ZSVNw4Rpe3DLxa3S9ZwnHjmx5Du2k+x1/fuIiapbeK4M3TaMWPHE0jIp7hD39nyUnjlI+SonIwMY
RyhB9Z+WRsk8wPrvsbx/MJYmDh6eJi0/7cPcBa8Ipeahsfc9iOd7dmv3jfdYtQjEb9riQ/1V2D67
nlxi9wo6GpU6n6EbkV7SoS7t5HCRe2CnvklzpR+d1ucAHq7JVApbDrqc5QV7Xmi7CWf4KyZU67zD
mHbMNFq/WwnJoL0YKVHooRO6d/WjYFTeNvCmZQaOUtHD0mh1lRUAzowh6yGkfoA5PrV9616mhMgK
Oo5DY2w/MrPjJxKfI/uc1eYnvLGl0HjqAdBtL67HSUVBsucLSy8ASTPK+Q2iJbDiuHhKf3LwfZ9A
LMtgx+M3hDNJmYV4S2LwkEdLjfKPPLgqolaFrdunE/BJ7V/F6KMHAMz3cY2vRy5qyhYhpk6kbuJJ
++pEMGxG3zlqY+69PinUNcIsGI6n/jr5MKhj2QcvH/IrnMk/5QB+ByfGCnbwZKfrCTOzCyneGrAQ
GsBCLhZ8c9WkBmVfjSwcfvCG0J9LvNX6bqziA6ZRGf3VJXcG/ByPuc8MF8lPbF0HrQCS17feRuzs
cDflKj53sG/QqpHbPziNW3CenPgBQg/q/+CinYQUrEzOnjOZHU3OjXXk3vNvKk2+S4hWSZwV1yru
Sb73c4MsblO/EFZU8Xy++BNpHvtqm8+U1MoJp8f0SY4IwRZBBkC1DvMgIPvp8E0eoq+QE2JGfD6T
lYDvzAD8BF+pLaIqEkO7S60z9UpmoIsxsvBUIlotfGc+36TedeE2T59Mo+MypAR3urEZEphlN3/d
uv9Kk/egte2j5PAvpVoosDc5Bh5IrNj0meRT01Hu47NkXLR5EI4g1RnAU2ipqq+QxXJYoHceY3LZ
lOCwPYHh/hX828QOvChijJDVKbOIb2/nVNfLAR137vEpt9IpVzaerhArTr4sUhc8W4pq46UpECF7
qqHvk5EDo5JVdfA6mUzeO0AJmMhjZCV6RByhxYFQZJKuZj5uzYAVygFs4VSUwdz7iPpkNSl+s94n
MXL6zIL2HfK9LN5gJVoxpMevj3eR5Qkbwd07QxiD+VG4NqncLTG/M+hukHMxYja98sDJ3+sd+ov2
pCuIrddnZJEJMgZdAzOg0Kurn9ezPACRjzFn2A9zAoMTYXnzuoBO0xgX9IWwzRlTorVxjuUz4tLU
Rg/jzvrrJCP+EQp/tLNVD1c+unlrtNISSCslxskCCUkO37+SfLuslYVpSLcsIrlMHcOSEso0nuST
DN7apsYFAN6ze436K+jF6GaYmlMoQRACzWUUJDwEtmI0Aq/WZEvhs/YliVNtU+73yCO9WpFlQf6a
HbKtdAOtEgB9maH5aYhM0g6L97WUEp1VtnL3Rc9rQ+QEik63XMS7AUgKy4+BsiEUU4rMAoCo6dWF
AGC4Ycla/JWQeQNvugX9Ad+GHlSnvAA5BnzMo11BzBtFXNTFWQjqSX4R3+1i2tofIuVHzrnLol6I
NpkySIeAmOV7kjq5UvKrbygC/un1pLHZq6ArWlTaub1M6R/o/iGSbtUdqjKOm9pcdM9RfJoRb5ni
9IRUrPMTQH39ocFH98SZwRs5GXBv8EV6pFag3VnXBKXNgd8nV2LjP+L3l2vCOqrcMcTy/2Z7mZyr
oSQS4SuQlNJLNuGvb4Ru8DAjpM4ZjIvc0gwSCnQ4XnoJh8N1h3bYpOPlVDBNKQh2uVMG5AAol+CR
/1szZ/x8ct/aq7WJ275nXD/tINxu0PNDPAzh0aXiF+sXE1MI+dDtpXX1YoZHju4V+jbt0anJENmj
5Jb5IfIk1mRuLn915uVMMn9GyAJL8sJDeYx0wBj1TQRJhjOq5eGlKHTamTCbtqv9PhEcsoQ6JME4
35pdTQMN4bQScqJoJH9HPx0qCsy0x1sl08eIG9QJB3lJAfd/H8TPFnvMAxOoPFxzQtTz1KHuaRfh
VrceP3fQnKow3hUQUr2VmlyHw0NuJINV/an2d+qRA7Chnbrw0FxgYOjU6/9zJYYtdInCfFFEMxmA
qnzcLMsgrHt/SJBqUVu04SM8uTrydqJTPXsiVHaEFegj6GEPzNX0BqWZ3Z4lI1ZV6Udt+q20dlJh
D2bL2vxp0bUx8xa7J12ckfgbuHuPHMDonrWSoBshhGvTUpL6SpMv/ZWfZr/tLitXNgk485V5Xc2c
hwJRNVOebx4BPVeXuS1hOwzbQNtSb605PHPbu/hh85Y4sdOs/KpnJ8X+mdSPHGATvGda6p7vtFuC
t43Ojkh0CKZJ6lNWYcFCPqZHyvkReE9cXy/g136JoB7zNQuamzIXyY8gAgjWZmzRNYrW7rXfRBv2
CVnck6tJDWF32RaRpUD+NPhfcpLQPljhrB0dLwuYWVTxm22+t11wmjfG50/BfDwh+r+FMGBjo/ZG
E3KyCs8kSPJaMBHBLprTwBjpI5Iuhzn0k8b/y2KkW86y2BI5Cl+xElayLeBqy7CVVs0LrUNCF7+t
Cw6HizDXk0dgmP2fkXRtU44rbWZNUVg05dwncND3hOQth0IyZbG5hBOJrUV876/UiB7W+hfSOHYW
Ke7bvHdGBjoYIOjZLQ5UKWS0vCI9Tu5mIyGE6LdDGTCMtE+JHjYRRF41hVvBYAOXVaqWURf1rz84
t80PeOu4O9s2ba3ptCkVH4X9NSCQquGufx3ftYe20SBtVh4KY6kvo2EdtMMZqAo27HgtYIcjBb6B
OfgXwBpP41psTzFs5h3IFvipwoPLyFvyhc2w+GzPvM9iLlmtm57GNkDxyA0orFd0xb/pFH6TSuWz
1+cXlwcyGEw1SRIj4GqiBbAA6Z0FkK/RHjONYNYvEoVNiTyXrmW9kyBs+T047cYjoedTkv4Y5YeV
u2RdyiHvWNBxk6dos84wjf806c7APiUN5F8pWBXH1fRQm4mkrQIZFBnAbSN4JV7ftIDZRuhyi/+9
qwlfNKKlsDNJ0rVewbLMwyEBKxD9BkRUQ2edex08YQn8LA7AlcMhxgTPrbZTmKJXLvWnZ76FuvO1
LJSUiO7dL3jVanB+ml2n0B4hLy5gDWcGEC8ekM+2NMVml9CDYAzOfpU62hplCjyPCyNwfbbpWEPW
PssN9Ncc3qnrg9zXY+OpKAZ08nkCmGQAQIXYkDpJhK9PD6bD8QjOosQ0j3W4KESnseKhBHA8Lcsb
Qhm4cLgJoXSVxyhIADUKiMetPEeKWuvs9G79E/0cpig9uM1adkUH7bYMsUBlJoAUQmMnM8kQj/2e
nPD+OMq2VCwcgUn0B3/9fsnhIivk1PyP1H01QoJn+l+9zlmdyyuF/j1sH+fEgUp+8+dlQQzujg+5
dPM1cAFfiR2zjSZLtrc9s/vTwiHVQKsKpheR2CN1PajIY60VrdLrLKI4dPZRAaCynliV5H0UcLpK
3pT69/HUKlc5RthIsp3owtbunwbGbJS5ljfiIaf2jpwFLtCkXXpTUCK/wdYqdkXvyhr+XRjaFxTg
rbO5DQ8lQAWPrB51sz8Nz5FwBsOdlqA8hZVuJ+TKeSmREOP13hsHWm7LYxRBm1fKopiRUYZEOy5R
eALGQOGXiVugrY8BlTdB3f80jrWRILIFqnrU+VskoInbHMq3LQGb0lVx4WUVi05cwWPakGx8WxDK
W93hENPqzLyrUcT8dk+cMs4m2CQNqa91dTMqVg5PKPHm/+GWZz3D4f75qJ5emgh4Bu8io8/8/lXv
JK+GwF8v1GQv1HF/6uqh0fVIEICt2VOQqHqbH9IY7YpQD33hN/DqLxe5GZZhjifvCEOK/mysKtYU
qWH0EaS+/l1U/EHDqvunxz6qR4liC8R0caisQfVPAfQlmGIQTCmD+oQurRxkzbyUcRpPgGX5WUi/
Ig9xy3l1g1UbURA76RpPeErvR9Mihmx5RvjilAHQEZ/TYSG5hwbTze6FPjjuAwwI5P6MkKE5fAj+
X6cRWQrDJGg+s2sRZQy9UsDxM7AlUrynchqFkVYO1Jud19HKgoZxKIOt6DZH1/892KcMhbluo2xY
+MpD6SAfkiIeSSDqZCGM4cjvd7V25qsgcbVQfW0BTdFWh8RlJzYi7rNiaZQDMjYQ+ZjjWK1BN1MU
DflMI0b/X+E6/kF8nj9wdl2nvxhPLdFr+SBEXH07uzx3jVkAcHQwj1GtFeWxanrbZP72IcurU+4S
vWsV9LV2FYW7H56D7ogi9V5MeMVprZMSdzgswaOJiyxCYAADCfm2F/kXmB8BSbX5gFqXcT4UPAmk
ZLCoCe/xASWh6f/8lpTNvAEHoxzMpHMc2I1mP1Y/onBhfnTSt05lawMZEGEfdpeUZThGCMigwjBt
AztI2cktCvkHmaLCn3VfbxHj5sYJft3JDivGfPPSEi7FGSuKPRObTmz+x83Ci5zsmzqP4K49MleJ
Is/FS+0IrP6GyVGeBSwQLroJMZphXA3F9+QArSSLFGQy5fpKjO7rpRbZKUT9P2ou3tred2BAHlpK
TGor5q0/I5O4lUuhtWYneAQOY+Cqe7mFJDTPH3d5wTBlz5y9ycc4mzKSUVQpJyTGs3N3AvcusPys
8qiE5efyHzR/30ZrxOvotYZsGP2pt6D/GphS1Jyo649nvJroZAQJE+txMQca1XYeipxu4by0auyZ
fyq99Syn282cEDfzaHj3P8JWkqDA1bq0paAYnKIyCZUfCisdBKUubd7iitzsDzxbvYFuV4HOxasu
jJRxm2ytDMG9t5xXsgYcuIc5oguJP+nJ2OoLUlFbF7jSZyhlgQAzHd1q6uTjKhElxTObFksiS68O
qyftexpcP4D30zNIu15UaGf4+dDuTVji+/8rdCHWI6yhKvGLLk81mdkXcwBfJUPRxXqH2udUuneE
4SuVS1xc3id28cZzGDShfkAw/0W4zVax8+RnClwc15S6CSl0Bj3+q9USfGf5l02hv8sEQIQ++gb4
gNa3V/qr4HLhREWlxA/bMtgg1ov0lmPhy3iOpPq8akUuTOG9jmUiULOhiyUFfY6a286CR10+a2aL
FvBRBgyIC1GJ27iNRednlmANqZyQLzfaXWH/27tdTEN6BdCSKD4CbEC0tbve+z49YkxKvHqurlpU
C/NpXlsAYLPWWDtd4c78xf1ZjDBaq0sz5pEf7LpF8UMRJl92/7iPywDI8Q1l8IZS3Ddrpczm3igY
UwFEmNKT00Ii5FyWtR7ALZpbniXm5+bJAYF9cW7DX9T4nku14cZd1xibjQmYchAeAXKHqP5LQZGG
Fp3jlAXYt2vX/d6CgYMYEtnFPuuzIZh0FzC8rSUXWRL/JGZsbxsey6v1cvIO5yaSdlbiUj8mk7ZG
TcBbSni/H6uwIyKGpa9uCLd1QPwfmoo6jATsRmBdF7lZpzXxqCNXt8A759Co85jnswKdq7xYf35V
dHJZqBjISSfwPjAIbUwAslv/xbFg4AU1mm7Ej3TJtaFUZKEDvEwcAnqsmkDsPMto1z4C9Ak0p9FG
luQ67QbswNDAjUvOjA2yhpuYlYBtxUDZmx28AdTQEjsYgZ20eB7jLFKi/e6g35g1HvJsz3/HwKX4
lY2s3mTwUVxTwYoPir/YbspeUazlyIC3HbYO9rVCFSWFY68bvhim1N0kI8S5qBc8AGDWu4AW9U4f
whqOXRlOodcJqN/KuP4l4Vl4qC0I+PMifc4n6Gbopp7REuM0eAiNmx+WmCj64MrctpkqQ3CuwpyU
cogiH9EaLpVKT26S1S9gP1yn/fRU2wQaLlvA4VmSoVc0QymUQ9hBpdMWi6CFBb/HCrG9V3ZQTA3A
x3QbjByJCg6OKUfvsZKP39mnvBa232LHTFxqZuV5g8Sta1gqPEOHo17oMqqdZ/JfiM1Tley4a2st
2VtQhNkN+s2ZWTUmPHsDfPWvmHBbODuxOlxO5Ki4xXb/2CY4U94RHNvBe9WaeC5yMNc+PkX0/iTr
3ggTRcAqt8EftpslbNx0QHSmRlgxeguM4/gWI0+V/faBl1dgqV7iexQRHUAFbEnh505bxHF9vnLH
pqsZHP/MX1f1o828DmzcPe4KaOu+Z5TgynKzruCPIKFEDyTnbsdn1Ju7W85F3gvPluwPGqVd5rH5
aNlofPSFLKMM7x9kjVMRW/dGEUUO5rvBAlfXDyjqee2PeXzPXTMDjxbprIOIRR2wYlqUKc/OaYek
mZ9WCTcR78xdsT5/GGgxPmAJt84kCYBISA1yVD3KGqGMooPoNq4CFLNuCuxj/pUlKn78H+oDM8eD
PJvxGEfgxi9bob4euCY7NZKISNHvnan6pTAn9igBKy6at34fUVaaOPxHt8aU45+pVhfdRJKlUIXc
B0iEgI0zB2JkphNs1NI8Xgv00FVttQxRRkjGSD8bMJx2X9zjoUSp2bStY9UB0gw+fzs6YyILD9cg
XCTLWV3NEy6o40Awq9FO1jxQa1FsDMBHC3g+mDXRK+SRXrudwpn5RRfA4w1A1D3txGANQ//UEFXy
jm9tunmpB8uIv0q4WIu9fxC9n0kdnAopmDIYPipTqTz8jkyPB/3N5HC492mlZbIh+kxNQQrHbsYE
z+FT2kNFwnKeyCGI3jpGOuskh/2hgRCP/I8erUa4AVJrP2L2Xik/6iKmiSQE2cVqMC710GN9B150
WQIUvkuVe4tUZtIJWfDQto7iMXSCwSJDrRhF7R6s9UWGXw1Kkhd11C+3s6ySWV/wqDDzGeg9zOvM
Egzp2NTs0hWRYgEjdTQvSUaZWmBlsIqbgZ4I80nCgdXgThfFbRwhGwiD8n4EmZMEF7YqTwj81LvT
eL1S/1iloD/Ce9bmBSrukdXmUFpRobTph4Z9Za13z4Rg1Dv3r8Vw4Hh99o/c6mij7MY00N3JFRnf
6GsNgKceumSaCcMiavTLQIeHQPf68eqxbPHOr8mdg20968vdX6ILJNsG2G23qRixMgjbcQCo+V32
ptWAddvK1zvogfz7O/34j1ZAx4BrttOAIaVYrTOk/VJanyL9TdlOFK3MzXDSgbs/LSQQ7DrvdsWY
crny5zKoFxahumpc5ARLJrlv1kyvShtZ19bJCsMOTdMay0fa2c/A0AOGNtpKE4ciT0/+ScohgxUp
nZIntbdUDglVieS3vm35WciUiPZM38l+8dzDkqm8ftGvrCyIeF5hbShHpupToRczZa8IBZVQBWDg
IOj5Ni6UGGnaCeDijdfgB+8bw3n2KALPcV1c+8c7qSKUmNgjoY9kJmRW3KSGflRexnofYWQeFplx
VGUP7vlQf+C0Y7qKI1Yx/W0l5wljnaJ/nm4BEBD/XEOcrrZZbi0kyK9g0OkV4IvfWCXXVY7ba63V
OAvpZqjViwr60nwiYmwPOZnIYEOXsHGyGDuiq2b69JZ9RnCaKlLJE67nMaadF/1C4ey2nmPfC5UY
h7VCOEYmjuzIVhJn+axc925Fd3AG8Y4TFk5JmBkZqWOuyMdSiRidamIQOFn//xhaiumhqPNFA4y5
hpRNymEiio0U3Lvf++ZA1ddFodEN4hkMYqGEoACkVY0vVbU00SdI/GyWb0/nnWZPZKUrBWFFmfp6
4qyaSgTPHvhErhcBMzmuQXxuD/2uqe6fVPgrUSVcz72TwXLQcF1Ukc+LJP2cKw2vBSc7fpL6TlxM
ZLit92s5XRjMiLgwpqx48ioxe5jeULgKotw4HJgz5GvC5uozuR2hO2jQqgZcAgRU4X/hErTBSNLS
uImFJrG8LOfXHp1aPV4W6N/JSN5ZOUfwrl1W+E/mYtsAgRBxX27FXYvPwCPl4Jw0z5oyISOPnmkt
TMwt8C++YDZmXDNfWGorrKpZ5NQTQxS0XrJEgvfJbTCx+klxB8PT2rvSm2tiY1DatSLiMFlfBDEs
ZKKIvzLL2jPCNmMmTD9aYHEiuKAwpPNpSVxIjLPSupM96XzFuyZN3U5WBF8m2mLcm7STvJF2Zc99
uJOj5a98WTv6JwI82HxNNrNauL/Uf4SR0/ohBagMcf4JDo6o6rfDcKDK3g6XPJfYsCzWQ3b0FtB0
/heAOC9rMhJH5wJIGDDnJMM3oAa65Mb4Xb7CM5WjLJxdSwVfrBRcS0v/BW6bvF43vMR7tba6tEZ/
kQJ1vZSPooBAREKx3V3zZ2HQD3z34WcJWNOlrjc3NdgevPkSSVTdLT1DKHubS6Xr2cP8oWPya8ev
ocJrwE1kYDIqXrccTGhhspybtvU0Fa4Qo4IJ641zpwqERcYKmRDR0Dx99T3GIwwVIVihIgZRbXx4
FDPdnuAF3ZwlMg2ZEv4IsNPA2cRgTitlCZjuZXcYqQZxn44idkTdlLp7tBzCXx/KI8M+5JcxYn7m
eav1v8lBKSGmvgOzwkdn95N62+xL3U+aCSn/tA69rRnZriXs4Uadmaio0ZOaE4QvzRIOKMui3yTZ
czCnxhLAzyUIzZOKjL6ARIft8XeNfhezQLmG+fdgIH/nf5iu20D1jjvOJB4eeRw35HG2zYIKaZ/E
IPDtohBDQ4VBN5iPvk7e6QYxp0PskrN+5zJ+pjDsexx3sCjmXZEL8t7B7hnai40XsACtez5+jawU
oejzv4xasuARx+Poa672sL4nnGF1NaWvRfTJXEr7Rslba2EuZ1MmxBvSJIEOnD9/PDW4TWdggtkD
Jv8d+StmaEVhU9zcsjrt65RtZMw7HWfwzC/dsQJbcIXCDKzr8vsun5p/jZ8ZAZqgojDjeGQQBgeJ
BmLXzg/hiCC8VNF4VRlV0525lfOkubKubM2o37NIuNt39NDoC/AL9TVrRjxfRSkxUugUNu2Mrexd
agFcoUYQTZa0/c2civ05TY4xD2FtlvaYsZiXYANcrMbAKiSArE+nyLz0s9Q1XfUArlX7FRWXR7fh
+9OCVsnKEAYWvyOXp6T4STVoI7OieESegQAp3otmxoLJ1uf3jzmHNa9AUaBevNtax3pvq0Kl61mC
84eq5zElschM9j5+dZIkSifGtOeVJ3oq5psqt6QC9d95nacvGjyqmxXoi4/oIdveJ8Tkl2rs/j0A
0DZq6GSZ4wS8TJqDCm2YdWTP+wLQ3e9IeWrvEGjSyeyzF+D6uOOpqjyTawxk0On5BFQ0h9CbJuRr
JbRFp/PCogT2U63Wt87FWLJrSfYD9uPyV62KlWw7bDKXR0EXri38ziQiQnxM3nN/qKTgRvYEoX8s
6JoCpIetWJGkJpg5vxerwzOceUYIkcN2N8Cqiv7Men3HNKhn6GV5x4Depf4j+Sa8PcqN6bVOe0Fg
peIYMPAMN0sI1QDYjepnJVBkbuCpZ8NP65mh5kiJiYMuDotTNkO/LyYajCHFp09tBTjRSzsLJ4Dk
s7Uyg8sCpSMZoDYzH7BpIMkuXRk/7xEAshrYfIxoQnzaPghFaY6NtSQkRXYZg8DqFbzakkzd8l/c
7Ik2w+Is3Lun31oSEy1RALdDboHBnewrXO+Zqihdif0tz2UESUy32a/p4YJC20HYVsZc+OwMQ2qR
lI9jpBNl0ybxfeEwG6JS565bsWn2MxjQ1xFeI7ViLionfYgMrX3r/02qCfOBqcLuT6b/kuT3a9gO
hwK6Ya6pWjEz1c4xKUb64kfm6n862Y+Wmt00Ad03ZpJFRbbE9YzTWOa0o9rhLVqGoW2kr4k2wXD8
sNaY/D3SYNRFD7aWTTxjHdVkFfiqLMOxzL4xWWPFk9f885Vkq440pC5wH48GIFIZNREgM+G4BjHM
Cl4pZgYgFfOflIQtwRTeRLA6u2yiqAUHjdlcGv7mE5LZoaBIQJcinAuie9QcY9xDWjWejCl6m1o5
dWMGH7gBJvPxotsK6Vwf8NJEy8vgVCYRb0lDsrYLeZGr/IPIZ35VJlha3sxAmYazrZ7KNSdG9hsw
6lk92QoPgi87M42a+sYyvqGUcVfGgW+W+5YSvljW+BGGP0d6RsSZ463FcmLSRNWDkZVyNK9aVj1s
iduK6UXNTgYZtg6rM+ua9M/j1i1fWUfgRdZKVHWdwGmAWd8uFuM/Q80SsBjh0en0v5bdyBY8CfeG
7Qog7rWcw1Ikke4XkZweMMndqsEfhNXQIm9H27T+Wxwx72sskeEJYNXAzEVVFf5TiVYhZyT/dYnL
CT9ywPke8c0Pvnr6adnOyw/VHBgej8i2P3QPRvbquf/Wh4pelT9GYN50QiM4VlIg3V6Xj7LZkeXw
TQafxa9GsgmMcTeATZfVgWbpmz0BtdoeZeGPK+BMogkOCxTTw7Pa61FY32uU3nDUgsCYFBTyayx5
hswlo/2H/SfDi4Hdzb3lejhgpImXeakgFGzqZXTJ0Kmfi6XemZCVpFxFWGYKRnU2jJfcgU9q5jDG
lo0lUUOkhqWz0dbIJ/FtzITu5cBSzdGj9wO1fyDLtSsKJUzUwIhop+GhVczs61BaRd77IIql+RGL
bmAc/IS3nTJHfEPQ2TBwk4ZVE+OESdnWEj9orMQA12oXjoX8NbZItCVQYy0xATgfeA9Z03Aii18q
ulVRANfSjUEAldvCkumL5vjgZC+1dHbcUeKALwgFdmcEJXATBPwLK0kcR0B2dtCFs5yeobmVBsat
EZbZAWTUppUPf14uP6soXFQ65gBC3TsDaFlL5UJkyiH9Qd87GCuiwrPOzloliK0fiCCSUFeiTC6V
bCNYd55e+oWjA65+G26XRESUIY3YxVL7YHu26IOUxh8rvoiH9ZaMo+9UV5nEXcq3HWFI4zeI3s69
KTuiPm3myv7pXD5Feh3szADpN83ZRqvukgH7bEYcUJZ9htOWjlDxTaVoMYeEZrZzWFrErj9rmCRR
uMSgFXOkzX+6xmB+jO3qJfF8AYCZNFT8qHVxumBbedEhr0uTfyGpdXGj+ZaS5Yc6jX0NvTmy7C57
VOI2miUjkaYrdrNqt4Z0YGpJi7vViJzBRmHpcFffS7bTiSan371qCLX7Dym0pJnkNQr4+9xKkhs2
AMU6O7D9EzEPyoop7VLx8vJOiJiX9SWq97Pnkl065SZwCnNXPpDwKXSFnQhjEncafv1TuEJaKHF3
TuVDsSigjoIgKPu7KQNLyTAHgSDnUvJgLwLI7bOcQUBYTxxHSyYDEmWpiYtkk+IF1u10heOiCfbm
M/CnANZWfjSDYo9cOq+/atoecHMJ2qaOx0VySOg9P5yx9SAQuh8h2rJJo8UHSn6WprINV16fqQSv
VtqyrABqY6/qH5Ek8N9Bp1ND/y2fAmkON0mg59A5EIpKowzUxnJi9vI6BhQZ9M9s0LxRAkRrslw5
w2f3A6+B6St+8/kneQOWG9hqxMh1eMPYD+etdwpSq1QNpFMweRdaMTRlJGD6rbwMbxfN7drz+ThS
MXr5JHffeNRldE1FomJQbf1SqaGPWl/0LtDgH8Z8rYW+PwXutGIZH9ZBNYZiFIQm+Jb6t2tGPX1a
xJ6G0IE2yMRS5gbXBs6/5g0eDwRwLDTjqK7ec+N4QrPR+2FtiICXiS5wyMrVPB9s/3I/ZLWXyhOU
rzjXpswHv++kxbAaCe74V0xa2HP7PAZbNnz4ELsuR9coNnMV8/gVYDNNy2faVFlYK6a5GHwQrBbf
bC8+zb+9xFmc7Ck3oFjNpeO1cYONmvu4oYAdKrxokric8zTtjXLv2nM6tA5rCkJtLlKmOmfn9oc9
4Lm+UkC3dkDHzlGNvPEvg0lcccYYQMqpDMa6zJ1DRyLudhXjF8wgnZHbSADDCMwK1+Jmzj4ELS0/
4s8dk7bWTfs2If1PojD6K6mAfD1b0eGksU5rRctPAhxGqFyioa/wzbtsB3oGxzoEhGTIOPcKgzMp
KdyoZZvftCgXgxmRbrJfLNdX434oyCHqST0GTwUlGq2yQW8J6/m4XEzFOJEQ9bffCDzwYeHwDTuK
p3rbIKt3yuBWsEqZF3RyrSL6jdfctdRTIdSbsQ3mqgG2CIJcLyI6Pd8dJRMYq0hSJig5vzXws/lR
0GhmY+oaZFnS8RjaZMGqzVBJeQY/DGnIorLPzT87GBnLxToj8GfyT6Kpi1SEGofXpJv4Coo5fP9d
cQ4Eoco59TWwcbF49ctzd1UnqVHo/FNNkdApibPz5bnRNhl8umq2kEEs/hBsHdIZdzhWYwd+2VC+
2Wewk4JTaFLyqkCYmW5HUMctI5u6My8KjuzowdNeTuNBxflc0KVSJCsOP4DKVq5h2hsi7P1Lv80T
B7NjyA8hQxzsu/CvJPMsXRn4clnBp4jqSqb4uTH00OERfON98fO2CYIXt9r2qX5t73UZlNTrtmQI
1ZyrJ4mqcwkrF8e3qVfagrf2SYHOKcZODNikPlFlT4s1zx9H54m7B7n6mVAp/LcuAj+K0+0/CWR/
LzwsI7ujSLgpyJmjPh6QJw+nYs6lNb9ztW4pbNlIsDEkZDJ+1bhQv3woS82v6OhxswGLE8qcdKkF
5c+A8pHLlLgfNot65OnaAl8U7FI263jnn1/lfuEAnY99VXu0m4q3/ltOVw+uTTtxKXO9PSkjp4Kc
FRh1jAcc1w2NmfNrQ91jZLE0QFg4Q4jiiOZABMLn4O/1vVs6WNDl9C5pMkv2ftdQQzl1PHgnSO19
WsrBMtVN/x8bMXYanJ+ufeNdSkBjbo3+vTplLyUQYyEXrtyMRrSX4DMZv+VO044BZwjIUVyGb/c7
vXENEek46tzYjYZr3qn5JWHnkaEJDrzvDiEGgB0N104gHPatasYfOdXAj9WReQBLP5Ff9rllxqFr
zzvfz6YqgUwMaqiUtd73vxCjMJ7/0yZudAryLU81/BVn2j+8iRlIWOWy3TyxRFbAbAvgSKhRBZeE
dIJq52tviJnxJQAl/sVD7kJnxQRFupO3rNno6Fvcmfb9XuunIau2jyVg0EbWppb5rcU7FWRScMEv
zh403WhNwZz1VOwuMSwvyGTzp+o34lTxmgoPqgw9Z8Iet26lZ7pKjWiyuy1D2lu0to3hvfN1NtDu
VeZ/bTVwW2m4qDgDEWG0IShP8hJJwQWnKYL1whTqWRBfrX/n8ZUcd/ahF0m0z9REwMVaXzlEev5B
wU0+xOLsoj0GXPqHZ38XtHgifl5M402F0xeuwO7Jdce4kSm3R9SG/tDhHRPEXDiRaR+6+wT9/HmF
zQTbhlGcAFmfgRFw5sPA6l5H0EMJrjpdwTp7A+2DJi0Vg/sZU3di8H2ivYpSX0wOUNqOva/55cK7
6LCH0rEJFEoa/W44UVkCWsnRQAQ8XJJ5AK08W7Wy2KypWc5hiVE+19loqucC7IKt8O8wto8HtOU4
8axGdU70ulj1IT+ROHofouMFQVX1WooHTUs83XXM/xZrG8W7jI2Llqupo1AXeQI/af5MKqtrZZcr
FO27J75WEJ0Bjosjy9yLoCeI0iFXkuHzsaIib98IMT3Xj5S5rzJTC6xy4HBd1HY5x4aWW3FGEmH9
kXMJm3H+zWShJUTlDw9Vs4v905qiUgrSTbR7AxWSERrDtsksCeYw5dXCVIOx8S6AtcE7Wr0uL9J3
qkR5iBGApeUwlsTmrMl2ZTW7ZKlpoGcmyQZNHNZI0wbLk+AQXSQ5ZaNeIxuEAnCJUzMlyD/m/eNx
Ven4BR+5DnjWX3VMR2FFMujplkMBg03JwlvJLCd86KLs0wh8uHDzM/3tw+lI/TWy5Rfp5LkGi/Ru
7zd50ensWaEJ1nGXkRQfr3Qb4hmAO5/pv+zjPvfehg1m8kXzPHZE1Zp/ccLoqJO3fgNliIxwQEE1
oMM6q+VreizvYQJ+ldGgg9N30N42B7z5crOE2Wj52ne2ym9bc+wLSxMGWwFoa9kYJ5mcMr4LIkSC
O90Rd1r5XzO8lenFHc4enl7Bu/WWH7rWDWxTkHFFOLT7+zdWdPDrVaU65gdtjLyM0JOqK0O1k78F
BfoOFX17yV5dzAPp1MjDqujCi8WEagTCmjcVjYLTKAggpI9YeXRLa5JCwnYAmyIZv0qUzgb/bhKE
kgvj2N1OvlfnAWwhBzcz/JeLvqGQxgTVvuTtIFNud2WZl2pl7nEQIHGIL9zwpVI2txe/EjRFuk+V
rFDpj4vuHbJtVrqamfimI0MMVmXh/h8g8GtcIB8O2qWhJvJgzTFZ8DWEEinoFvlxhml2EwT+bcRe
jRDptwvhQiVvk29Au06XZMwo5VRfOXSVxxKh+E0uVJ/NQFvB4Ap9gEwjxbCicsZDI5bBfvMnrF0c
TzJiJxExIF2jnmbaZeOiKSC3p8Zkht1TNJGTZTTGE1LDaZRkQoemdqwwbL1QNzaNUKtI4RkNYgb9
R8lfTsm0OqJqFNMpsI4Tvclprlje4pLgF5Cn+m2N/xxzjNfABNzx+rZpRBkE3fa5DXJaQEeKIx3K
/8b5VsADcnYgZgMOP6Ql5OTeus/tdzGfqDwaL/0TgrA5Vwwy0GDChE2pJ7imYA+BpKWs+L4HWyFC
yZCWnX4gD5gDcSbS2wmOWNWkcdSDCrQES4IDmK4j2Yez2+IxTaewCUxm6vNY3nKFZMFfm1PaHLWW
E8IXsft06TO2R3zwLWGhjrKQHNGR5MLRNOb6muavPC10q9AWStX7zgej5djjyBdYRmhwVLOlk1pm
dTl+F8KSwV1xX0djASg2P5O8jtxkl5sB6dba+ThBta7nvAOiJ5+XFipyVt01x9wfAAm/idlLX3gZ
3/ml+XvBv5UkD16GmNPi7XU64uCF4bXuvYs4MTh1rinoeqcd6xasui2LlG+IdzIvsWb3Sx2WbaBw
4Xso9SYoAaoIhg+aouxAuSiPq3wdCcPA0BcFr4+3T7p+x06Nr/DfwhiGOW0jjpyNaPQX2iHvtOQS
V2shfSY7uc9zEY75duWB25No5cU+b6ogRQPZu5GJf88ZJZj7e9ZzGrz7mXjaLtzVN/i4MLIK+ejm
hnIizP1JwEK9ogwKAVsSRLmsAim2PdOSoxSDWNbBgbt3fswQNapLgqYT4bcnf9tPA0dUWSbYZRxs
Vw2Ax6UMJlPklbUB0mGGBfOGuNPF6IcI3QHPLrUxr2zfGEb2amCBT2t3o1W1SFrEBtlrt4LDFJq3
zGdRjCtwB/X8arEn3Vxbqfgga/yA3cdsDgievDLt1azjjM64zVCwEjBgSkraBGK8j44mtK7fHDb8
7okQoiUA310/Lus616FpzYyutZQCnBf3rb0VcCJqbkA8kn4fHmNFyl+FCFLkmzJp1rc5dkeZMYOg
VFUnidl3b42NaPj5gid1pz4UNr1EAQwkt01KX3PKUfL8fONBh58kL9bVLFPO9QL9/wh7GuoO7Wvx
9LgBtumKD3GH0Sw8fs4XcAbp6UbSzGot7XQHwZ1bRfS8WXjbziUrc8h6H3kMvTqeK1zvTdTMPmms
MB9tPqxRJqiclcpoQrhASkmIjKnCS4Vlzs9LtMv/SuXT33zphanDpY5bx1qrhrEihmIApnhNyiSy
BQ0Oc0WvxlDe55/JUZ14IYpAjbtPpWp2h7maw2TpQhMWt7W1LTPQI8rZYPmmj5TK6X6pDPMB8cC5
P3AyHp63KHBwHR3T0qZ/6PDNiEMJWZ7Ah6xw9eyn6ttNSu9K80n5+yeVT/WUoWW9eUJ+kus8j9Eq
JifTuiq8mg+7dTmGEvuzBsff8//era6yjTgn9930JbxTyvPklErN8yS36tpxAdi/O9wjtwtZcI5z
4V5uBnbzZvdMvDIi6LUztlzhI74hJF/tLiFHoYe/B/gPaKB1sbvID+ga9LLOPeF4KhKEscWv6V6h
KLtRok4BiDVBL1FISikfW672VMdGJXeEDDt6TSB33hL70PJNDTL/6+2eK2v25EvtRzLtMuymxJw5
kNi8nz0MISNSlSLqkLZOEtKjyyCUu5f5GOahTiOOOJrqBi7CFOSgV9khCOFZaVi6Z4g1EoDb5uNK
vPdesIImlzJO7abiwVF279Hg9q4tCiIam+4RSZjM1kitS+BnNJgFn3a6J5eTMym33kWdoFyndiMt
wQAkoVwlXJhK7ylzdtOWKIzET1Y4Z06s9mMPrjuwBaeD2i0TPbN5Re6hFAFGgoSxiIwMPeZi8oNQ
fByI8N+SrblGEBhryknSbHEDR0kPb6Vq3mN22JdowRS+FGTNRxYfJmdKnpUQXy3C1u1lheJ3+Ukb
clCZWVimmeoqGqDWyo8SQjo2g9Dd/50CyoPJlfb1z/xqCqAB0W6Hr/i1tHa4d3lVJ/PW6YSL+5ud
z3xvfiYZUvXXi/3cb1rZb+g5agrWE4UuAnFNoBh0hOe5TDIZ0rM1cDsibHY4xxRsTh6pqoMBGtp9
0nv+lp6vgvN7yI69Qa7AdAZJYDGdRD+vMSRsevfkG6Xorkv0HDAnAMuCwX04xHZR/EQAcmXk86Gl
/U8DKasyUqw0vRoIhVMhoU5t37T0wSkbFT0OEwG0DMMvU6VDQu/1HI5oYzRzTrvWyr62pj0Vlw75
dnGy6QykcpMz3DrQpoHm9AHiZLzeRi9OufR2am33+csuWHojZ5qI6R6tF2BBavXweyyDdD9UVf0j
3NZ7EbdDcTHxceoeZtI43L82boyvKpmIReXnChUOrsV4YNcQDs5CNislxLgelYcyCvhzKoQawgTJ
Zzu62vrFUqOl5wCNWYTnBi++JUfGF9RD0KtmsoHmJJK2EOoefsBKgANwhi2oG9Aj3IQBp3fOzL/l
5GozOXOa0QecUwVc/yP53uEBM789shcYi6/wZu0hCdI7w7Zokw8eSpkZojz1BYlsYxWBG5hjCvSy
9IlJ/dTzXtWwRW4ZD7LCvJ0dWsDqlDVXX/0VVhWn18lDU3K0uH2x9Yg5r4Kj7xDrsj2cCVrMeuWm
At3qtzlGgQ5F26JilG2QFKkYQTYH8+XMlsGsb+0QAVv9m5Z+eU+LLBfKunwIhFAGWUacDdW28Hbk
l/eNBee0taKtveYg2Zvmq0omeOamFRn8zqV58WecZoCF+4b5rlYHyhW3N/POu5ZvyByE4EG9E06O
5LiqF/yyS0bTxeq1GDcGc0of5isJ15j1oDsfpot5oKz7lNrgBxht91yEctieRhYtHbqlrmf4DuoX
S/6hJnn1ZqPk45ThTYH95BwMnBycmvRqL9sjzY6fmio8SXdYOInX2e5VzXXRG7QnZxTgsYymQ0KW
DiISKxdIO11FC5D/2k6GZrXCdpOSiNc76Ac5L8XO7MRr5ETu6TL+GAlpXovx5xnTsR+mRfYT/c2w
5b9cIcTWAr2o0AOWrOgkg92VQVQVNj0TGUhp8SzvvqnD66ua3yGPhlZbCsNw7K9WnE+pSEgqUtZo
YEf8bhDxDA77e7o0c64XhH9GBhRJkOYw7KqAHbY9tyq9EhL1d8Z4M3x2yLd/f3mjIivJ9Fl0mhQ4
OLW+yaEkE2SRsaDNifmjBMpAX5Ysc/+ulqr+n7pJdYM0fWLjaISqurvm/kKfMJkzkjyCv5Kg4+5W
sOLqfyZDyh+J71SyOSBlgKAn0CfNn0nRt01CNvoNJ1vtuJHl3gz4dI3QKzwlrsDM6r5q63/ZXsME
gRA0Lx1Wkp2MKTo/uTjShy4rFVT75XtmC1dVA4ToMfQQrnvcZdaxsAOkxQMTQwYsTau2djAMxQ82
4DvA5MtzKUl7VXjhtsrlcezcw3l1FFMpzFJEAkfEsMJjlAfCsbBi14iCzcisGwHv55titSvDEc3h
GAZsUUHZ5kgYcgkXj83V68ys0phOvvvzf2d49cgGkcj6I2ebvxSWuGoDSaRsdn9JFpsGQcKbVU5m
s0yfbxIdGyrL/It55NnkTfOQcIsayFQP8t6pCegWBptGQ3OOnFsnPLN1Q40+8aFtsH/ytIfdKoG2
r5BmXmY0MFQx7E7s52K6u4fP0mbWJOOlcj+6o5/Q2fs4Q5kV4Z3UQESFzkLB4eCP35D9kVh4DsPQ
fcH3o+0wMnQlS/oZHHzh1N80xeKlOWfA/+NS5IkX7l4wAhCWDceMAqg1tzcLIU+t+5s81jmvMscf
u02tFNYAv84ljbVpuoy8WTO+0Cyn554i4KX7dsKwlrUsgjuADHDTafJOZAo3WMtX5LKwpjJKC1sW
+YZQtujloWMi8n11SKyAUuHm03Wt5H3os+H5RDXpcRp4tILvveiw4UXfQ986lw9UkeMbAufX6Jrs
LZl4fV2uNHOxtiY2xa7/Z+ZZbtzH+LdMprMnmQ5T16T8ciwiKQZu+IGynQ2i6O2pecFV4PkSdZKi
FLNZYi4Vl00C5CB/zBmETZyKQ8kzH4HBxwpf7vNRQTxhUwxalWSRLr6vJ7LoxKEzkbILZIol1dAg
8//xg18m9scbsPlOF8sWc0rYr7tJQk09Ojh5QvqHofIGxW8SWfSs3x1jGdjffmnZYHTXp8yr9CXS
9sHup4L1jtJ+LQcKTzLwSAzL0LhtxJAhevEGS3bkpA/tCSpLMwVoT2A5r1PuyySiS5/uwik+xa4/
Lc1L5E2nVrWnzj3aA/qwzENmDcR+nL2nwDYRaU8zYwE975f5NmM0+WAbJX+/9UufxNZ8GzfMXarz
VRAcyv0RH5Nn+9nQLo4AnRDgRX3Y37RWlIT0yvnR1vJ+MPsEoS+PSHpLzZef5jOmtymHebtQxfaV
+6ZsH3t3nHR5appiPlBQlQVLw1tCExQNDSezEbc+yCTDO0j2Lyy4wjGLkgagXevqkymt8x4hHPJX
feRY9VHm6uGpOsKe5K4Cz4PJ5AVOxRNP8vfYaZpuzu9golHVoHX8fLN3NI6oKn7xVz94tM49Wbi7
MUVrwfnQvl+xx+DQNq+A0WcFidSqZc/ijEzYt88N3uf5WmKAL04UUcwghyNKdAL+fQahInGeCCTd
FmcpLUNDfyrrqUgIalSk93IFveqerA9FKKjVPQgXlm/giD42yB64DkvDxylKjYmbYJi0WfjgFHu9
5S9jj9yummVkCwKFN6mQ/1BaaTq68euaFDFy9aKpSJW5zd1rkVU606x9VRXB6kiUGwtrAlhC0UW+
dOxZlNkyVAYSD4sMAaedfWpExjDzO6SH56fkuIr/hhos4zHqN9ifdKc6/6b9XFtcvFeLwQKda2nf
b2CrXjgempdybWWbtDBCiOac+y5CFbxjHtIEFjRqaySoeJo5Zq4XjECnSoX7oQbNgQEk2uBk5Ds/
OPU7cCa+RokZObmXME6j2efB06uXKCwN3QagyKN9/y/BD40Ub2fXgMoS0Wn9YPp198O//unNPDZ8
4Md8qUGNASIsoRxAIXpA/wAx8QmtcTZc7cZaY+43idDShx2CP5dQorQkjGizjidSRAyqndTVxkdM
hJ90TQD+ce2cm6i4n78xea6NbstSTQCvNjzRpc2/zJ1JzDmz45h/t8xGlUn2yvIKSM4Koczurecp
hNEyAJNtiEZIfjql8HbL6MEfiopNrlXdDMAqX4HKSYv41JZZpN7R7i7FbiQWVO+qgR7Gq5upzdpM
Y092xioYLeXmYuQnSh6JT9pjTjCMoyIulLEUcUO9CnfWQhGUMgnTZer8mFG8OCracH8XRsUAqv3E
5Hz3oSG4WG9iQM3tD9R/lTI/J8bF1unI/dgJybGID9W6JSjhxv5Ia1yVh8CY89MZd4xKpy9AqvXR
V9PbKUVSFRg7BKMC1+xBTJeJUziXweZogFwlpuD3fHzRFeoQETqdzT1qRC7bLmVEdF8sAN+sivHp
oYWRJjta3AHPJIs9FcuRVSb1JIFVeBilcqJ+2R0EuFLL2HKA9+LNhQIxqkjD+HlUy1MrAF8NHnSN
qW0ly9h0pVp5ATtqV3aJeyAjezFmVElHN8kQh1yhrwWSaM5RDh05hPx6exG+DTRtUL84x+UH+Ew8
UGKsQzqZvO/C4SSs0/Oa2u2ZF3bMNkBhdK3IpNyqXvMVnwfaFTrgaeFChf6qw4MuM/3Q2E1ICw+g
AbTWHjjzCNyiXn4Up/2UR1nFSzcv/QXfjmhBe/XXowmkcbn8I2q39Wp8jfz1Iuv7BhAZnG0KG+Sx
mlnk1pk03cda+QidCvPsT27uhihf9bPCDu4Or9p4jlwDm4oSj3+xme5Ets3b4GjPGM4DbvwOrWrs
B7UUKemajXZNcZjdbOHfCX5v2pZjgt0ZX7InPtsdCs240eaJdtI74kExq4zCdsqXWwoA87n7hI+8
wvnOy2ElaJlEtNEEjNqihIm6TejtZ9VciQfEuocUbCNrG+2zhgtMjqTYDbDXEvZ+jWOVwr21QZSS
WrlbZKeFDNvc/ruBJSLuQtk6ELhNQRNSDKmCXZHpSmtWsedbanpR8jbZVLe7jflQX0hb+JreDt2Z
LfKVmJ93cJWke4UNTc3t63Q1iIH7opsFzZ7SdVI3Av4OEYluB4MFpO9IYLthNFxs/cpZ5InnBKaa
H+HJCMTSACa9ebB/2rjdnpuh/r6vOBuSJo++NppAEfkCMKXRbXabqevXPisLyTuLrTbAbkadfrYv
maa1slCLR6MQySlNqZOg54uqBIcdzSlg7iCK+NmQWCrb2Tv/kvOUqJLdlnxigcTRNo4S811RK9fj
rAUOHx5LOv0raZfE8u7DTwAfRbjbQVG6ynk8pbdRmFqnEi1BHwpPOSrJaQsgQpxkMCKyMC6xLaxI
Wu6qg9dmsscVUpLRDtXhRF6Ec0Kk5L2Sq4JtXss4aQ0OSbV2X6ed0C6RcxIdJAdNUCmhJVyQ1TwO
G/D2wmMk1jMT/Vgfpx4EqbwI2M/zHg7s6kR+HtZyo4wX3y59QHqAGnolHzyy09bPBPHo9d1BFBFS
SMYx3Hc3Jc3472F41QTlj1ynaxOWQIWlMInWmcjZU4jV1mXGHdWiezArxSNXq7yhavlys2xsh9c4
6Uoir7uc+iBjI1poiEXS7k5u3QoqNGkBre89jdMRP6DurhxnXbXbrF1UZFWzrzUW0qkOJMEMle1M
cZThm4Z/9GCxVOdQhGsilmPsjKM3iCWemC8u4gnLflFCE5yXNkqsjRWdajF5hAX3hwKZtojRxmdr
efAIyuy0zZ1cEjQyNoNOvzinVEbffhXY0TLA1G4UWGsRcJ6ZC4oPPnXFq513B+hZLxnHp8rLQ+ST
5IDV4Q3GddMG5kc4yDwgKCo3iU9xqFPZGU15PHDlaRfeA2KxXmaDogPiwagKnMY6sdzFyzfeyO0y
2CdzqRIPe1SifyHpTqHuewmS06gdTSUEcLFG/lfQ8sMGcu7pINCpx9eSzQiW8q1Y1YT6tvtmZa3p
v7gehbOtyLsTK+puebsJDQ8gciUvqB8D3NTbF9x0JzKNGutroNZC5oFVK6/NRxIPFyNCrq2jmEsq
DdbGYkeokBQcAdMPY90BJCt2/FiDbQoy1kr8OhIWFeU/qcbTC6jUaFsNshsaAzKGC/7q2d+PK5AP
b5v5JLo/ZL8MeNpCVPUqqil3MQnjwVPB9VZM0MxMsFz0Kx5UCYsQ21AStE3buCA2lIuo5KZYYIGb
VkiYY5l+sxzUME+bZHZbQ1aOoaE8nnkyH3dE8SEZ4h+Uwb8YkvG/LR5Fjrb8eX/iE1L98frVgGJh
nM7FFvFjagSlwdcLAJa1haoxHOpMql5WlknSWLZWlhbjM/ZJTLYtaSUfy9/QXlPaYATKRgIgJ3kR
PB1y8ePvF/AhT1pb5RlvQywKWz5uHncjFSyWAQNqPQ1TkE6nbjXlMCBym68SqE+JC6B79boOpu3o
Jk8gVxzyL5t7W7qLiLHiqmK3HTXisdgU0S7V/UAcF54fVUwJyulFWJ01aG+gyCOH+TvlZwaweDWQ
HTHNPk8u0DW8e+qZRm1aJ5pE1Wqlm5SBnQI1uziztfQiJrYiHnlF+hYst92JIaZ+EJnyKJR7jc1e
5qGgAm9TOZlOwcFr9EHVb1qOPWVO1l3nhIqrFL80sfd4jYJoUB8nevYkOWSz7wfXf6rEi/Ed9261
SOc85ndwS3v5CvL28wClQPPpWnhyRBzmt99awQD0KfSdwpCUOFK2p+shBvFxZnN5mLhCCQXHU0Ge
0cDtuC8T4LNMsCggovOhv0oUxg0uwuozng/wLaqVdy9aTloNAUSnL75CG7bIPgTOzn8sWukCxvJK
RS457npHs7IiybC22wmyjKVFulB1q2VtRmkYEUjrZnc3evrDbYWIGh8p2jdS/PbiUVf8he0tGZSa
iYb1W/gE9ebxOslsniAVJSs7Sxo8xXnuZJoxddqJCl9FWm47BemnwKKVqHJdSN2f/vyOY1QeeByw
Bq2nkJe+kRoR/8WGL/+yQtr0s1vxYjE3K96bx6obRsCKMEzvIFbA/28k1YPlWYXTvErrReoqRskv
uDshA0c7JkddJU6m3CzGh2cJM7ZbrgnqFOuyQ+CoKym8XqmjdmFQW8wRc+erVmhWM85XYERSoQAY
8qay8O5bdwwAWHuyliKItB3v14ECRmyJ/xKxqGSER3DIA/dvC9oAY5mutM2pzAwsdDbzLkPwplTn
MC0fIB4sFKwuviCkYy0w79MJSGPw/jF1VcjgufON0fSdKw7xL61nKYdwiKM2wlxl4FUgU0wTx3GN
DT/5DhbCEvU3VU7wEk4EkD1FKGmAFMUvT3stn8ZnJPnADKOhGGxNFsBD1sHQdp5n71+1yKFU39zS
nkDaslfmKB+MjyWDroKh7DThM39m/Pu6CyulQgGVuu/FR2bH3YX9LYrJCUXgCDpVAaGqk9czBDN1
W9QL0MNLnm9dLOgEZznuleiUEXsYKXSj3rPrD6rrO2PJq+fcVmhaXzYR9Z9X8J9xJx7gsVbSXsB+
CT2jbQgbG3ear0PrZV4osoa3JEti/M0NW6Q244EwVwfCxFI/J6elEwBO9rsjB/2wPn4uBmCfFqYV
e9r36mwKxdBeT0UEnL+QkmxgvYdDB9VuY1LBiHdCjK3Am1alNome6/ziujJofCwW+1CED/ZyuNQH
Y/HMn/l/AyjkN63QaQw/jGksxj/uc9Uwvu9IamWFgUcuHyVY81lFGMI/+cCtTAL25ZrdLe6dX5T1
NpaXwIVTNDcYFwza2Sl5tGD/kHIv/3zdxJsnxwxSerSTZZN8PExkddf0OLXFsflEwxmvogjt7s/e
mmOgFQOkGBjRZCHAGwuxj7L3WbkPa22h9yPsTa1nS/hF0LAtx/YDSve6s9wrf9zjyujzL0YX6PKg
zUZmB27sfw6pj59e5vBppSPXlqyYXD0F2Y20irUwGOt2HPD+x9C2ifGxW383JOwZHxSVVaxjY4Y/
oBWvqhzGzM/L2qUZNWkCiim0X6z2jSPc3+uCnjs+cuFdy77uLF4H2shX1dziWly3P+SBzx1rO/6d
G4YHRkZuhq2c/bgVp2hsyBzEamikP8uDEt6TXcoWlAQcBMNsSvAfOhzJptK/jH88DztV9V/+sGnC
ZbhsouXpWYuufvhM95v0AP73BluUYSXn/PhFW4xbjHSn9c6qX4ZiwxHWIFu1rYcRh/X00lfip2fq
3KpiCDkjN+ynIdyWVW274r7FUappX3oAbzMqUzDfYXZKDzbT8XZQRVhZdTtw2pOCDxo9A0r8Zo3w
L8myx7cE+FeeakjCSELUMeR0Oqdod7ZexR5oi782lOpY3Wi+k7TROrGGqKzwvbEecJ/VuXtwS5Uu
wexrSTF2nnYYdJDIyKBEsnUr4DONgZPhJUXLeAl2zigr9lrpY3x6ma9gE8EqIiwKsMPQfT5V85KQ
Xw2VdgVvISuGjn3D/YUctNC8g6OAnO0eEca/zdqNOMGevy16j92dMUXK96nD0YOYoxqeNPTtsQBn
Q2771ttDScH1bMk3k1ULpXoWimUW0TVi92UclmuLqMbQ8JhEj3kPOYecgUqOZ6nWLRjVrB8irgUL
BcoAKYsYtXwEYWHptbI03vweluezCLrLEo1CrYOPZLBVrNFlQtQvI/p5/J4Os2ttyD6Iqap0AdNA
Wh6puiYP7TafyQC9XeHw9mdrdA8R/7+eoRFcMaEBqWCLDlVZwUKi9FIwPjH0ezxPhZvHBKrS4Pq5
JRsrKz+AWAoOTq+wDzZTOhcBirW5XiiOBEMNGq8YAaFmM41ayFeZYthk7lX7dUjSnKgTs3SCtCz3
C3nzjJo9hnl68u22uOuetMSBybEPwghOkH3bLdrg6HvzWO/feZCM2vSv9hLbWTvuBjPNfkjxv6lH
FTjVgQsisCXty1RDwhXS04t+/abUS5o/7/PCgBWUt6gfPQNov1LguUO08cG0SBoO9z+ghwijZX/G
+uJNHClSSMX8d7/J3dwjfa/MuLC/l1wFxAmXdXG2ZaKVLYMmzeRjc0bX3v2OJcDodsvrM3/9PZJ0
biSNF3S8FQMNFhaD5H08m0eB9B1gbtPpdUaDqVpU5XlmymaSY+iRgzMmFCyp1OD9H6Owbdso3VpJ
VBGhKE4byxtn6/AA3wPOBa0TYKPM7Ywq6jTxzoS9FfmSqIAgKQE9GiNk1/OguNjRY/EhLOlvGjeN
Gjf15xUMTJda3PxJzpc+zxx6YGxcfWXTtvqXCm3l/VY8Gj9bUHwKZ33NG2cFDSM1ieCthHlSxNYd
eCS8tCvZvD12QcTOGb0glqsG43vBnGXihl/Y212tIn14G7yB5I0lLGxvaB7EpHpIvdUx+C2K4jhf
bZ5R/UouVg8ll7uWme02Do8T2F7hceTkl3GAWw0b637LKPJxLwWzUY7Ur1a+bD85Y5wiMb2cZL0c
0ZvKeLAmkWETnosww5/RuqDIHPoGxpMHvrv/SmuCbCmZmZedrw0fxaXNIUWYWuPLe36xYO9bY25c
urNnlWaQOqAS3ovqbWbyz48sTPgZOVC3gPQpVg/caA939uDO7BVT1Ny7SmkYAnNO3dLoYhbceQ17
QxsJQ960HTdZnrH6GVP1PVqtzWeLosQZQg7kAuK7LFgXCTIEFnfJ0onuS8FCondn0Lfk4EWUbLd3
gCkUFSAE5cKbBeXLcgTZ42vs9lrHfZcvLiuizPXj+CwNB1bzYxekJqYkIJJFwhgCl0RNUPRx7lED
Dx834dFsLfhKqouULO7RDFxWLE6OkfaKuf/RHu/d1YPQ4/m/+m5xZvzgd2HvDsV5vbRyR/shis5x
ZVy0kpZ5zPahbeicgVEtNv/6XS05fs1nS9gNQjtq3AczbR4yCiQ9yj+6tbm8vyD/meZu5U2Ud5AL
YEKosgrXWbhEe5c8FuAdaX9sMUDF7Cy0900vNj9Js67swU1/znpOgzC2f2Y8afOoVPhJPAbOPD/1
PnGnuMTEXJdLK1Dwd9OtkS/Kz0rv9TwlHTzYb20s+VO/bydI4rGCFf4t8PM+bHkWmFahzYFsb39Y
0IOa7sl4LWLW64jn70s+HXkpcO2e19hkEqiSq1cOJYfPT8AMs8gF5AmCEqvU1XDSzAup/q/UG5Sg
Gx/6fHqpfgi6qxxbA/xcMj8+Gcaull49sCz2q+5jDgiyFYhu5iAGYNjSuDdiPjxfOOt1ggKrlq/Q
qG7wAcm6U7cx3OtjmbFShyXcgRp6R2SFdR/jueZEAivQecjYatNOdYJnZZEAdiBF4WfcSSkVd24K
jZTL3F4MuapT28PLE2gtBVxwnkT0wFWuedTgG1hdWkUl6gtYDWl5LMDhmVgK2n9Y4ID1KNkgA20D
rfCKc0XQ9qt0n8I/XExW5R9wHl50xFlFrrfKlCbLSWHpfjS4Zc/5f4zedQGNpdJqF/oiQaWvnEyM
qHG2N5pkmXxpqPfsiebP0ZNPmu34jd0FLtF28AWEXN+u22N2Zvi+4Ju79HRVc6nhJfaNzQIu2AEN
/1kREqzMu06OEKsHBgM/s3ItCUVh/wnsrh9W4LSyuwQqR1M7RO6DUFjzDUXW6rq5eS6fVfBkVB6Y
L6Smq7eNkDw7KgBAflerNR8oSlMT0gV8G2kpv/GqnnPJOYdI2LqR3nHJ1j+hpSUJc/jAtj/cq4yx
+zmCoa1DMS+IPTVOM/EAbJeE/v43B3qf0mQw3Cc8fV3irBQwFmTkzcuVptmwq6WvSUUebGuKXnKp
wNqySZEv4bZ3EVqgI0ykbxsdAiBw79rOY0V6n8W64MQzZH/x9oEnNlOA/2uYlxBfV79Pez2ndZH6
a5hEUa/ybvPb4TCXQr0T9qzpNY6hAsRd6LyQwyWziTRbgBTPCyNKTtgAl4/hIPi7FpyFLvMHXlw3
eJwmzYWJwV5EUDDnhLcQ/3E1pcOy+3xqtVJFGBKhSghFvSEHN4aU8ErKz5MVCid7Waf3jRnvRjfP
drj+kIpncCiYUuyrNvO8R9Jl15z4YAMQXtn8szl3EQjsBnPcy2GwVlOK6TSaC133g2h2TBz8JXUg
i8oukh+QFAbNjijny56gW6UGxxf9lvPCtBC6B1PtAv5pCxxuCONtJO8MstEeT+wD8rO3DhbWEbME
EJD051VscgoXU2NKQwEVIYcOgqVorOhZ9f8c3+B7LpxcjRAbcP2Kvie688EhbTgvwoAASnCMU6cr
kGjdMpLvmKNTSiYwNuRjxJZJX1CCmLCHQSIsVTHlwtvpXmN2SThbAyENUwBzOeBlQPgi2xl/DWbm
W4k/6L+Fq44bRLixJY7gjcMm3SBx5Pah6UOR3b2PEUwQ4rZgjrbuGcM1k+d1tAE1HjS91p7ThUo1
CGpkf9T1rSGmbYaRLGPoI57hdzG2xjC8dBtlOQGZ0LbqlHz+1iIl/JDKIrLVZVgzTEipJER2FBDT
dlsv+o7OXzXh65V1UlURS13FKdYGI7mx9xOKdLURDS8leEDJZZGmvIx1bNfytbfMcUAppZli4DCi
RGM+NfFtjAUBpZMVSu0PhqimJuOBNW1nYCbP2JMKD5jGMn8waqP0o0n2tcIdGffjVIWFWK3hUAbT
slNQTOnzAki105wgQ4TkM6zpGPDh+8aprnpcliEvF8pZOHrcFrB5RJbckHy+O8J+UmmVyysFrD6G
fyIYbs870DfJl2zljDPHn2Ig4lWp7yAUjp5WFYw09WeSoN9g4zvdb8oX8YKzlCIWDUKG0Cn1+1gj
2iwOeHZ+AxitwnRqX5g7QBHcOKPkZL963iNGbz9JE+0B8ZvfwXJTpscTPJNEmLd5ZIyXIHo1vUxH
mFb+W8hUuw+uXFyyYiH4YeTiNQlXOMaORD/NtUk3fMZtR8OZgptfOm11kE/+8cUfKg/2+L3CAVlp
YcpwrEC2Qmvy/8TU4tbqg19TsD18PKXZx1tOqRofrAQX4JIOUiK9u0+/JtWy3eWw3KMvFJWiN9Im
ABKfYKddpcvfmd5rsFSWVElpQbRHKwYtBOSf9uQn2gHc0rkRTBIQnL+HUwehF2KVwFVrNgFCjO/M
imQnRpKgqX+q8J7T1abKbPlTf47xnrGrv/1yifg1Kket5gpM/b+Io5/WKbHfLvL/dPk5JwCthcIy
JpdJvhssfQ3vzLIB4k9l/EaOkKpdKIxVnsANI+5xx4Vipa8VGCj4a1YWwvbwmncir2gFWQga3OPg
5mFPVM78Xt9Zn/WC6+wvHF7WyGTPdYuzyDZmRlSrLLolweEP5bOwej3v2sgF/5T3h8uAeyMSCfzW
G+1iUTjwLW5cAFh3wPCdFKpYiDW+zHWiqXNVXA/wHSSNDKLD5LCmK08SyB9+xzWfaxYCurwZONEp
d8FwbjteXB7pHPJiG08CI5JFb+7wevw20AfQZ5cvnu5CWSn9FtRb4/K9nrheONeee8HV97bHaDSq
oxWq4xo0ICSVqCNa0iqvPekiFXKe+j4AGzUjSMlhBl/46r+LXsNoNqCDKOclMA8z9JgP5NHWaQkS
dpAiI+nbTbX/36JORs4n9FMmkB2VEnIu77RJEjut9nlJk2048cXvWgsbyfs6bSIMbc4ANvkdTu4k
7ow4F4YNpSBGsCxRuZOVCr2N0m878w7aoFVP8SZgcuCEMDvzFz0xPLaMxjLafygNRdw8TOJ5tNbh
GXZNFw1OZGNMzKDssvNuVTx95jnLfPNq86l+REq1/fSriWUB7K+qM4lbCiZEXqulKNTPvbv00Pl6
OSRw1lLY2EFz4f5ZsKNZpMNMGqk4u3jqiUOanhqedf93c+8sij1Ny6gQrgHtc2D/Ba/iNduVPtKT
kgEmU+j2sa2Qiqg9O9uDYmQaD+dPF3i2br4WkH3SXpKNl5sy6ZYoDjR6v87801UEoJOEiIsiejac
ehTGznD7t3sZ1C+DPdYfqOMyfQpIp5MIt4Aj4FsNgytxan2xwbpwxFKT4AsYVcXzLXYNQVxHeZAZ
fjdY5dRuSRgFsTqrnPj/3qe3K4haXX3Apldov4/fJhEwa/4oZxJY0e4+GMkngQSCc7eTfBZknyzw
dBhLQ/z6lrwqerr7BZgjTqiM3Qf6g07K6c8HeLLDn7tbGfVsDZhtVxWMRlCDHN5BJ+NHub/X6NNR
V/FMoql/XF1qwygJU84QPIyMH54m0zVVIaMs636468uz3PwJ/OtJ16bDnJd9oJwXEZ5FYm5pG4yN
pp9MmcHhKCasZ2OPWf7NUdEHEkeYK1pZqQphjh4UEE2SsIiqfIEPSNO1KbdqpezRQOwTZbCsssAP
eDp6fP+zW5KiLE3jZ8ifl8UsEF1eLbbYKTgIckvuERH6FGrsiLbjAP8qTORtyExQrPvZPIuPslV6
zDH/WJbUtQNtUEQm1XL0P8FH6OBNFoUsMdu1p5k2Xk3P1qm5ujBdhnigUeoUwxM636+pB5Xi/PUJ
XwRGGy3fDJEe/zyvS2DgitBqx4VQ90nGcvylpWmGqU52NTZ3PG77AK616B/F+jd6AlC4DL/WQjZg
sWonsH7xHHdmAXeXXotaxxIw+bE+Pg0RlsZZ4C6rX0/oyLlkJQMzNiCpiusQ2vnVBbSg+JW7w/m9
4YAc7uG3Lw0EL4jo92cKiUIVkVu1gpVyS3QgX0/Ile8EzOYYm0hga+v76m1ohxvAoldgsVqgzArw
fXOicU3IbULp2nUj6OlEo7XDY2xTjTTe/PVTm+S0QZ3DOoQcgiweWzycFln3N3TBC4wCHcO7ffyN
bYeZF2JqDBfJJF/MWyDrESSQkhzT0bQc0d2xFlWweu3woXa5zVpb8utlqjwwemkUroUSM+VBvUPS
sPOd+c1FBiuJZuDkW/GUJf7GqVEuRlrZSFktQWihR1A6wd6Ivmo1oxO4wJ8OIhWSVR08r9IYiNcc
pSqWQYz3yn/XgnRdLG2cUw1P2LdKcF+5l2wMQRdTW+emqchV1rsxnR3DU1XyGWxWTm3tOOttgl6S
Y0T+xWpQWS70sVi66ci0WIKZOHC5itxj36vKqxr9rAQRUh+hnEYB9f1DBeOfEPWVwwVnHSA1EZm+
hTzLmSYltAvVuW4vDfVSHH6+MX9TDMlW5DzZXyecvLtpBJ31+0p5bIzVhp//W3vBYE9bLXWE/IUc
Pad9yBBGvYuSXSODoKQjTiKDpq0oEIFLYNfUMPZbjohOgC3kgsw5i+C6Ve69KW62b1Iu2MDSxZmA
tFVWZX8knp8YHhkKpH2DCgXYCA8GtiZ2wN8Q+MiAsdj1J+0wJZuqo/ms4p5PycNWPhyws4MAoA1e
tVepIT70HYqtbu9B4uTpHGoCPXyQr5vYzamyV4oiO3mw3X921tjTsAQ81cd7eCO18InY3bisEyPV
P4AnOedEIEbdf+c/TFHJlfd5j3tUFkTRo2RrFU+WFWq5j6+VGZcGM/owhZ7f2hg3O/17s4eUuSfX
97qs+xkNcjzSJ7iKs3+kJQp2ReGZyK+LCsPSKKwgBH2QaGLdjvNnyLwkiOlZa+0BRI/lW+CczydF
+b0MSCPQNtXxDrhND78VtHtxlYQH6raWdRTchUnxzK2Z8lbRLVYGOkdMJi0juEv+jJW7Bf821amH
m1zlUTKRvacXQhBbauTE78QknkGdZfF35WuPPaba2eBceJK6o3SiHjhoPJ1kAjDgO0+wxyv1q5p2
u1bEgYu/SBqZFPkZctIH3+9UuL0VLMjnVkSNtE4HdMamvZg4V2/niHV0dOR0YHejN8CJtsl0i4pa
+tYYUeis9RiLe4z8ousB45ZWPx1Vd5bKj7ZOcA40pFuVb5DbDtiEy/GxAa3U0ulTPeIAOAaiOL0Z
lM/wdZWLpPf7d2iiOhSvd3PapsTYqbHMgJn2Du90hUHMbfUbiistP9rozvgUE898QDHdPsXTpWlt
EX7k5BmVYsjF2DsPKKzstc2g1IeIReXhMLwe+zDOtSjfeLr5jvRFCbXpWHNE8g1/k1talsYZwBHV
av8BsAslLfeUT6eP7O3hT5ZxzdUib6ff9MIoINB1wf37nih/QhKftw48WDrbuBVzUBHIKxEcuLxa
PYAW7VC3InKmF8Lh5I9sn1ya96ghvDFxZ5kd9lZmdPupAyRT2cBEi0UtAAx8dBO8KJlfEmOt8ugE
2Mu7B/puvp6WSyn5/oUx2DJE5HqlYcAJHxngwXPbxcbbvMC7JeBZY4GydqQk1rFPNM3nLIwObeWJ
GsEKElev8KQ8grhk6rUCTLN2xxw1DvFjIFTCcEVEX/mMiYr+EmxQhRJKUmlZiuXKrLKlChRHBnSK
P7cqVIjb7t2V9A3Ve9GxZXDSx/yWwGF9zL74+1L/RZq4GwWnlrPIi8Nt1OQ0pC39CfChjHkJdlq0
MUSfueXj1QrW+tf/YcvUsmBkX48C0MbulFEzUMHLsVudK/K24pi+euko4yokyOsv4jHYxgPTJ+Ls
4HlHB6hRAxvk4DniTq/nANZA/PnHX5OP+3odIjYQrEaTSmRnRTnP6ltqpYIOGcAY3rJid//+Ca6S
Ji/kKPffFH5x8lzVYh+9WTQZ2U3PTgeTMEzQULJrNOlO/j4w+fB3WP4zqbFwKrcAMpLxvR18yjhf
d3b3CtDQtx1+sjSBzPHkC15V/pnpiUDeK0GsYeurdYcfrk8oex8g959opwuSp9ZrFijcasiXGv4K
xOmdKWu9FivfBRrQj1l2cVEKXhFURFxtO/zppg6yPakH7AFHS1nN5v4oVkuemCPvUqW4+emXwihR
jowmWWJohAx60o3I78L114vCEMYgzPdoFxB/M3b2Q/NxXYFSYe3IJz0Ax6WzaBO0wYfpLd+hV8wt
bwl75ik162orxozVhkhEwUEW8zQnMFUk90HdWB66OEITiyCJRw6Or2xWUXUWJB4uZw+Is3PnVkD5
S8iDlBm4ZARXZ4hI9zHF3gc+d1d1k/QUkPPsltAVZhVolw/R9QCeWxwl+GNtbL0E8fettt6bqGLU
/J9JlyHjszEpIlQz+2CjIf1eVZYRJouDd+h7J2bnPFS4zveLjjugUmbHoXy8QiI69dT4AGOvXd/w
FLred6ALKUHf5q5vZy/0xE+J+0FTlSpGZKAo/1gsCUf7xON4IpFyhbOs0oF6BzJdtLpTHyU5cuMn
K2zVsmLPSyV667Ky2Sjgp68gflH2wipTCklHLkBEdHEP4LmQW3VZoukfa0+v9PKrgqiBMi9Kf5TR
a9cs031SGPbUHtNDeUCXh9gniwwlgHp3ry7n89hiaOLufGkktpxUTAYs6Ru5TbCcvRHqxorcfnq3
WWqSA0DiBxgOKBUaQpYnh8SE2Sp2uQClPpdwH2TGj2ZTjuzqU2H4mb9OQmJSkyCvcvw1g1s5aNwV
g58TO5lo9StIvTkTXnBrUoYv8kAh71/kivhyNYpbg1+j54kstsIKxwlT8M400QyCTPUsqvVdGDN3
7Fawp61F8AtW3rH8JnDlpou6/Gfr7BzqsB+s9/iIwFPANVMuEGFm8uLvXNjsiZYCHIep1eYm7lFk
pGjGaZTjYnPO+3LPIs+9f+KmsTiaqZsXKet1gnFmsOCh+oKAvrfTIfMFVGxGjCisXfrNtH4qeqt3
wTCkg76Bu0QIVO3yhVMyJvLo+J10xmFYZPo7IABty/S4TxwdWzfCmWOqFFcEcTNnlw13GkH/pZBH
vQcuR06xQNoZIJc995UujXEqQ8PahuAJcpsMZv8A/PtiIfy9d/gIwkQYTx8g8sJ5XLqW95D2YgXb
gwFw1tipZDDS93fB+4P4rKSEeNCxy8faq65SWeKG/+ZzwZq3PT/5iibgNXPZwbHe8FWcHo5JMREe
seob4aHAek49TtVq2ia2nyaTvQT0k7maGoKviYs/CrlT4RWC5jjgcQTRhB2jYZ17i2BKmo/lu4Yr
IOM8gX8tXFsa+X9QNwp/vLw+NR28ENX2YYu/Lz2y+tQ9LyTbmkqXFbrPwqIoZMynqo2bLOqIRNZY
/gyGIuswzTXrMqHk73Wz5YBxw5e2mDnKkuh98ilrK1jfU6AvV/OguZkb0l/EyGP8j/u9HlkAP4uV
6DjEu8ffEulc9+ujh5UGKXIBjf3DTcGdQygP2c+ffKnxhZXipeaRKeaMDWiyOLje1RtxJRyAnp0B
ySPPMgsLWxEq8f9XjUk7Sgll5dXnlcWvO1kZEHWorvH2EiusYaiZP+12cgAWVHHY+Mzo8oi6XLEE
jeeXOm0bZxx6iz5DPYqOTYlS+96vsl7GS6kaz7yJ/wK7HdF96XO1UWXY9wiOcMgcLYjblz/jtc7Q
jmqZCfPcq/EBYt/aedSuCuhXvhVLr+55NA3M73FHN8g9YPlO5TAzg8t9qWbIBfjS28BwnEBxtnbA
sMNNOg9Y/6SJHZOXJuun5hEnrCv0C/X6I5paEvu8oJskxeM+kRme5NE85ac3G4SUNTvF6jUPuAqL
iQLKDdJm9uRR4tAZXcSQGZWSjNq9tNCZ8Z1h4EkCB53EXLSlXSH9QUyb2aXdsscl28oYs7sUXPlM
Tic8l7k4xgZaFIHQHpcktzobViN07EbyNOtmDObjqxCu7e75gTZMpE5UYtYJjhJm/RK1UFuojV3H
4g9mG7WKezT9QNamqOyaRdIA/7a0RNUN7qDc3/BpLYYtTA/J/bCmr61P/r1Qk/excSo+0Bva0OzI
Bnqpf7NJGIGAMjQJyuofwRE96cL8/UD4TrR+D5e3ItQmSN2abB6OyLGkIM4cGqZMDN6zBbSUP8ad
k4M8XVRY2nrn1/6ICMD7nsQzWzPWDm6BM8S27z0MwYrcq0z/DjtU/lPi90a6o5o2ABY/lsMnJDfU
J3hTYWMxquqVAQ+dgkPqSxdE34NKRlowX1aF/Abj0g08VQA0B7RL6Y7SM1/ITkB16YQalcpVfGqx
XM7X5S5nVWwWbo4GGlvlAFXuTIV3ACBEvRAC2LL5zVQz1aTvATBtW81FCgSkMNaO3qw7Uw/h6Thi
smcQtWVFtiMb4/9bMkMLqk90rDXhx63ebVRUnartIyJVDweZ89CAzeaDjR7jxtzwtcxuTTzRSEkP
g+1cZJQmBgNilRBKq0DC8OoydYwXTFiWLlIQ/egFT9hYCHgeYWc8tctRqgvniblnDb6pbjJSGCxb
gfXUpqeXMyAIHqQBebHkQpWgJ98C1ledvaLzam0K31S/SFNhgfnrCWwvhyjLSjY4mhD1kbpsFh2e
jx3ozOz6uyRqA6osGM82Bf2aDLDq2BuBs9XbYOkWvW3bsvm4pDwkGVllscGEzCpzkLCSolES4j8J
mhbYSN65yfTDb8G72jZ/GCWnH1Ug6IWLjxPfFub3WcDkTusiWOQK32mcb52+dZZ9XNK/ocxd/geu
/dyyecsBySCj7JgR5/K+ZSHug69EUWVItm308SdDNQsBDLzFXt/gUi2pODMkWmvNxHxOcoVp8DwU
BRmDwXAOCcb7vqEkvVi9UujqT9wvKDqYvVAhyZDO1okGKnnO9TA1glI9njkf3kuK65VP05tPc2Q+
iP0EgxdcFIoIrb6X1TuxFpEX3dYwbUUJ0uJZtXG+oShAYX+s1OLZjAFG20vEtw1mocejfytyrUBo
qtV5zhjQyzqk8CeTogA2aHOcBBIYV6QghslVXV/GPpnXbyzHvUCzd4BWS+l3JgFyola/jGCmMfb0
NNzlk2pG8ynwtWfHyBj8hl7VoaSlFmQHQpSj+j1/tOtuwRAfb5ygmeAVObckWol2WKNcgauQ6kCs
Liy8laz1bFtYLjJqnKQEcXs1L/ySlZwNcFLzLCR9hEeAV2DmuNa4bPi/Byj5ZEZ8uYPJxT2mu5HS
heQrdluS2syhDFWSKHYddAKWqYRCjkIDVGfKcVFtBA43aZXScFvBGgj6MJOQgPD/ny25giTMeqI0
llNxcN9dahePqLy/p1NA/PoNgBy54p7YEFSrKmwkxkGP/M88GtTvMawhkwVlYYmHnbLNLVGOxABW
aQgyrUIiggn3cfaksePvzCO0rNN7BT1dvncYoi95JThuIyHf6RKx0n5S4oH4ieF733D2NGk/3xIB
KKfj7Gtg6PIUU6ymx6bWorU5BmdNX9mdp1XoGAfA/tMPHhpZDAlmt5sprh97dVSO5bSF7CCu/9Wb
/mzbf7MO/JvS/8DlLhxk2BZMXZ9wcXMsQsvHxIMh4wQIqQkuUXwfxYZ6FPsIvt+ioIojgWQc3Yrv
Q2Hftjbkom16uwf9SU+vAvhv6ZslDyXKxLW0a/c9gM9CzLHLkbsDRjhEd9HjS2Il7fokNSmRW6cv
9jl6DdNZDV9LA9EZHe6xDOdDMDI/aofW0fnveuyO9AfnmCsu7ujzC8c4P7LmMFSNatfAbHpgL0e1
pv+Isczley6rKcYzDdlPliqeuMssriMAyM51Y6thuD+6BjjbY7ZHFNGZ/9WsFgqQCgiwTaXkqfpb
7Ry155YX9ReBfik3Ph/4vqAxMCAEuo35I4iup08sbVCbEN0DgDQshFMeA1IsvuCWqCEgqMd0bDTj
EFrySj5RxVhdA6vA2IvGRDl59J3ws3E50/Vw7J2P9sEikF7WVrFiMKa/oGtlWTDn1gTC2spOhkyz
Bw1tBZgZC2ODNha0jRBMd93zuKWUPRdPBcx99gicYWdzRH6aHMR7i9NiJfPcxpeMnixZ4nsT3Nzd
AuUZ+v9b241ukL1fciEuQtcup4cumIUTc+fSUN5KDqEgZHx8H7+ZFTbBu8Cm9XwcGtGFe291++MB
2O7WBjfbPdICgxUghUjAJDTtQbHGgm8qX+SnMwrAbsC4cbxCwPWOLzeMlrtklulqtx3PR4vJTspD
XcAVHLQhJWOWwhe5U0eAlOC7PW77JJBbaeSeFVJe/JeFH+GGqy34kHZDBxo7Jw+eD7RqMwHvn3Fk
PBDBu2fo9ZdUgiKNpbnyyMnRFtD0U/KlJLl2JXaXjK6N3WohiV/7NJF4jyC19QBBJQhGSB+6nSuA
ZnAuWIdjFOaLmG23gH8cEl2LIruNBwRJjMa0SUIwVMY8aRrwS15kfHoh+jIggTc+hW8X0LDs+wK+
PCgxk6rvfAu15vXG2mQo5hNgQS3Xe6tfU9h0VhMiHZ5PeMGR0lR62aU6YURI5ykM3rT028uatpoY
WiF8avZ8VzdcGczH5zHDY+UXTS7+R3ekp5LWQm71KuwwoyKoOmXn3lRN3ruoP1mSkWg/lwdfFWC0
JUjh/JEZx++r4crSKM8fzE/Le9dU8S4Fj9wzHmy83UB/vnBR5U4EmQ+H0uTnuUoeFvzIMmWWiS3q
vGKj6nri0RAHzf/p0s0Y/eVS9DBMYTr2WvTybgr2ieYaGbfXWhXc0AmO3fNYAez7A1dWJ2GSbd03
DhrJukSykZS7K6crJAjS2U6D0TZApxMLKo7/BeMWxxOt0lhIn8o3sH4+uJw0VhJgI6XuWGYYFr9A
L1+83AUspLv2gDWo1CsM0TDS1jN3lyMLf+XRLvxEnfgvYXSI/j4w0StBvy23QdERUS2o0Cr8AczB
6RHp6MqNVmu9sPM8o45ImHR76Sauy4I4bLznDDVcHctls6NOJCRDMKj0C4PRbPLaE8nYSOLzeu9U
+/ar5XqPSFsTB3c+0c4VVD0w3sk5HexwSWyuafxhIAmvyyB9tD5tUyx/+KMyZufFt97eKyyxlOml
nDEgMvZGOvsA1zGLyUZ+v2NB0A82dRNYAZttDhAc73bjaK1SC2juv8woa+TVBMNPjyS4+wmmDU6B
1EoegED/CmPBkgbXYyrNpexmCUfMkb5lLHoEUO8hHrtUIN7WwYBd4taKU1/48pqyzhBsB3ScV9W8
8L/l6Ile69IqdJx+T6e4GXF7+vqDBVnjQgdNWtrpsinGBenHYRGXk8ym0KVmHcRX61aChApP4s+c
ySGaa9GocGnULziYBYmRjU+hTcmHEU2iuba1iAh214254mtnoBZ+eroaIRRcTgUxbslTaW7VXxm8
O3/AGAmdmR8Ff7gd6r+iOszBQa8Ji7Aku4Aa0OilMV2D0WsGHOpMrneJuKSMg6PJlDagJ6ehWSOt
l99YHlg6EsF7Zq5MRM0wOfcwddmyYULb6QVb5Zeo0IFTZSMMP6qBFggs9XKEMju5RKWH3j374v5W
bxJVK1wnHThjbxXerI9jTaYVQqxIIzvZFBA73LW3lFEpst0HEcCxbUsyp6siZxO5sjqawm7lVpgY
ntNS21jnDuzP0jxDt8vsUA3wOg+M+kSJvvr8ye5nurH0djQY6/eCzAbGA59SkMKDZgdyfNEzwftF
htUXZyCvf0fp9K0o65Hunzg3iD9AcewUZL3O4StcWPAfXjpuIP/7u9UbMyIcGj7LhtV4alebE+f7
u0N/uqUxZdiO6AgUQsurdNruXMgiDlKZCtdlFdg365ywAU6EO3l5uakr0PC5brNHVXYVdcTIfS6E
1C5TvjFA4Dtxq7bAoimqeE5UXSkXtHnf6lJrzywv/a6ZC0OLUN0IjGBRT/8rT+MwrcUj3Sh7JLhr
XtnIxP8/57HxV02UikY9/RmeztlUDMsQGicHQuaYF8cEGnflOJCNkiVBTbgf4Pu1yYOCBHPom3vb
9NgAKGakHhnDHT+ZJPmYJkcSB9GTg5dZh7fi1KlwV1Ak1hSLVIXu18Lv+aa8c2wW45YD6BR2/y4p
dgxRe9E8yxCS1rruQ7bj/NAaYldhuBpac5lap/mZj8odjhwVxVgE5x5SLC4rx6mA3rpBtk0TcdG0
+DMych2TpFk4wheY1j4QYZSe2eoYYkeXg4ItEWM1/x54AldcwKSHWlB0kHhbgryufwRAqrPeDWgX
cXxDeL1q+l1OzcCJSXry6t585jU809eBiQ1+DQ7bMurlpn2H7VxG0arIYBKiorfklHEtfYz0pvgB
lDRpCw4gr4zPwhp4ojPHrS1g0X6sJdEnc2aFO8diXFPt5k4Ni5eo5mQ3veCJvK0lDxEy15+OpSy6
HJOTdRrqJmJ7U+8e2IoxouEi3vdWQKe9tFVeVdnqruPcaDejo0r2VDGdvP5NKiugULkffGbxb81u
R/TdLGuZgGwzJf4nZDDtV9RLLraRrjIjQ8/SmjrQGIprfbXVSay4LOvDLzgnJTeMfWP6Og8RLIJG
fKCqICwoeP8UnyqAdomfaL4XAaBd/CZb+bdn7nnHdOuf9kWaAWHwnqTi6lwhKTt0f6AKJVPCIi/P
hXUmjfadHULBp4348tSwG8yah6MxqcJ1oHHmPsNpw/AOEthUYaOPvzwvfggqTHfAd7m4doY5Zm1o
f7zEFzKtuuZKCD0aAnm9mDxGeD9hAwDvlZs5qNAaIx9IDvBQTnwu0E7unGI4+qSL/73wvMOr72RT
mzLNYRclMpADjvOwuXw/URpfKq9NSMW05J+qTicJa2agabv9xeXld8d3sTYAt4Z6LCYaEB8w8xCh
B0lKnr4CqQf0tPFOKAz1BUZZl1kocWLHrnVdMJSizG0+pcU+AhdQbMOxPC1Ekp+e2/dnipB49Dwx
P9YaRtQ4ZwySQyiAJlL1mrE/c3yz4hocRT1oWbr21MPcahe7jf88R6kRz03jOmtkFj3VR3f/evY6
uH6vjFhAEkvanhYdSye/TlPfAJkux8Z/f4bCCwW4gHCEEaLLmqwFY6i1MBiczfV+IEqN73yTvJHo
T3VwX8bMzbLTADLVMc6jRiY83rNcCOkmOWq8nOeB1J2CUTyE8xf7vMtWYFDWwJoiIVYTghMbFlen
q6NND9mwzUoFy6/ArMfZjpd5BnMqkST3VmA3+qeYBuMfTnPcGOAfpbvPUJlBE1Dp9iYVpctBSJrg
JFasB7Sd5Di/GFVVyiRCRRuVLf6Bwe+1PLCMrxHJp52Dwr/53iLayEI9NhcfSyxhhbDHJjqXszhi
mof7mSLVd9Q3C+5fgDXtIg/jcMaKjAS6GxUHKB3maMjwMN7OKuYwOzS5pUQZ/qq46bxcQze6YfcT
CvTJTyzshgnmmk2aN9DwN5uoPOpYnym0k2XTGnkmC8y9xotwXEiyW8UmKYFx8ByZIfH8jqTXJoty
Aiv12w9+wxVJ+9Wjf8Ktfa50RoAAQq+D9DWWRnLs6HU5a3mVpixoxitVrd/SXEzcyJ9TMf3dTBJD
h7USg9W/koimimPm4nYydq/90AS8V/bvRFZ+8/j+IEDWZvtZQ39Ldhcg3uWmzkmrSULbBHHvFzDj
+iMm026Y5ZMB1mQ9ytfkyrSyRjK+AQsN6rJZHYTwZrzhswD30oC0R5/G/h9QJ1TlSb+vyI7qt/n5
ArAnJr+C0QV1kFuti4Xi9G2s1mL5RUViqHiGsGmpFRwlOG+bKSsf+kA0ea4GR2zA3tSVq9U4HlsF
0g+UJpQtOHSvBq0CTahCRqv7Vj0Zakx0QRSH+vYkvaAATjMsZRPqzqfk4QNEmAZkwdh6Xvi999iF
wfHK+bgGmk4+gFvvCogrwmNB/pyM305ZDkHcLP0T4UKusWP+2eIyhQkvfc0DJVjaaDP2XXbOovYL
/Nls3bn4Ge4zpiVH3+IddDN/gKyldW1VRJFTaBJY5uOS+af2Ccn/8udmCjFAojsoqU0A7Da3WNtT
me7miLYizNEHpKeE6ThDA0yCiCXNvPo5xy+jL32CeG5sKueCrOZDGtgAQfAaKWSGxZ6ocMc9+vFz
SZRlDqtjd6K+dt2vzUJupsVsY5/ORCo4aJsQTvlOqzDRDcUhSVuMiqzL9tJaF8J1YNWCnsOH/WOz
sN4j7Zb1ukPAILNOzOHMgAfUFoRGHW6YrXeSoW7EWvjWPndX2bwx8d19raXZJkZ8VG1Itic68EQf
ty4AzACw4lqgd8xWtuZDGpYk7nnFW3Xy4/yTM7cjvXVWK5O5f3z76JkYSKhPiLBuEJZZqFOpoEZ+
tswo3VOO09QG6EotCprlzDptB2Y4QStdH81cbKPH9pfa+0yUE+C0jkU5/AnZbBoLkeKzzQ1sGr64
3OnRlgy98W7mT76t919CEapa04hS/in4WRMjO63jU0jJx4juVVONi6zK04er6k36tYQUkHnR/Y9a
mf9WdIz853M1wdjjbVURTZKXR5bCBIaJbW9vp3DOHrSj3JA1HM7NLTms8HLy/sZ9YPL0q3+F89+I
AJ+kbhmcEd1aAwRXcFnXtdlM9Kcl3h0hXzj5ZoHATFLY1WBRMuByg3bRLi1+H2TdGFSswdEeUSDl
gtlBjAanBqk/SbLR7/LCGfV7adTdR6wSEkKjxp2njUFx5L9+UfE4NI8fKvaWKjSDJP8MEl05ssi8
hN4QNvLlWzHMtNrtI8XkqNFoKrBOecNvh27W2Wp9sk9H+h9hEerRiGn2d6HXSUS1tE4qyW8f6z+4
hC16qqoUPojSTHHVZnlXF+TMmqlbB6MLzBuiBSN1X2lBtZsB7X65Sy1w+aCk0PfzgWWpRw9NOMTS
n7QowFwcE8F5oqLE7onj5gyGZqtyucv5ul3q9M7CAdlps8DKi0SeKANqkqDF16pRmfvQtbFzkgUS
YVaHqPWn8SExYRmE1P/jj7Yri3Q0neMyX6DtZdEgBuU1AaDI0M/7EDda9bpSVyz1839RjR2RAJuc
LhrqiwF0VUsII7gofoRi7+Lu6DHv0YLextiU6nSoPLyuAbo9OcUkIk44KvqQeC8QNGDwoSe54fDp
wNRGCGy1yRL3bakozRMHildNoJ06s/a7FdeVI7s0hr90oGsUFxkeGMhTDvUNR8o/brpGn+8S7d8C
iuWuRZK0TrP/7B7VEtakMG9hvr9aO5Cdjh/g/WXAIKc6qsbuHf8JbiJ9NKVCULC8/aF8kUEQxjyh
J5Ec7P4kudyfkRoZsoN5RfYXMvUysVDgXmBWOxWCOzg7pI6JyMtnAiH7GyHIpSN7hsVKn42d7f9h
Ad4yn6hoRI2RvXiqHsz4XTwDx+WniBAx6WmykKBpRN+Q1WAJu19xJN0Xj4TVoHWmbe4IyPZsinT/
xX8V/tjZ9B7wq+iRAZfwat7rZeh4C6phvJLiEHrHZKEszF4Mm76YRnLUSgQb7CuH+6+5k2xw6ARc
L5K4l8O+xQ4NdgP+oGk4i6njXJFmSQkJwprwp36W95xU8/Ej1qKJXKhwDSrLnaUIe2psVjwA8+IV
dkY0wF69agZ6ayNR3URzgV/15DCexkkz7V2ep8SyU+JG7slWdy687rM0CU8BHn2TNh7+yTwlfIQt
5WvJ5w6sN/1sNML38WVmp222xLK73Xxg2QmQSJEYZgm9vAt/2XMUBjkWqT/HKu8mshCDu15lDD/d
ZkUFkKwu9d1GfH170uP/gbmknZz+zPQQoHUi0j9Evy6jaPvWKoamH+2jhhnunKYotvOLqS9qciuS
Yx/HPDaiaLqlS4pvaKpjFbc2iDz+MG680GgDG3Xfpm/TQ/kSI4XkZDosqUktSh17TVNfFcT8tHAq
i2RRecw5PcKYN5Z/NTGwmoClIZiVuOrHMF5XeurHlkdbtIE9Wvgmxf6sq55nYw5N+19o1zZbAfNO
K0xnty28puei0X1RRvirR3b97CFrNCuJmjBdpurg4vl52tLpDd/YZCCguKWWfYNBK6gY1kXLM3HR
MUQhHzemYcW/x3Vp2ErbN7vx1YiaZ7RrOE59Tau4sRdcBmypihs1RD2Hp2kkW/LFMp5EuMrpJTe7
vBCC8JH2I/bXx7ybIzwA0Okvk6Dx5xFrEGbFhd2hM7vX4Rj4pvCbMGzG/LDSRixbnofxajmYyXxk
6tWm8v1UHJt/fq640FxHk6FqZ2r7ay/lB1k8Tq0pQuYB3QG9MNYYA+lV8UQyJCTjJ5enZ+cj9YbH
0TmzcanktBd6+1cj+Qq+I+06kM9fEbEwKyOIsohAu1KMpx5cHmsV1KhvCaM748/u8rQrTXfYiCmr
O71tSrSa9aLfFklbHl8Yo9WEz5wAmudbyjqyQxRnK7/AXFNMqzv93Dk1xzBR646+fgwFnsERAwZL
kaG2+AivGbbZV//Y4LyUTVKbBBSlY2ehsZXC+gNdqP735aqsiS0Lap6tQD8DdOdFdNFRBG3++tKX
VMNuUR9D4BosuP25WgkpG/+dquPf2PXtbysPdj4yc5Fdhos9EFpVZj3xqntVOUPW2/IIgNODKSvV
kiQ4hqlyOJS1LTapgKqFDR+c5ZJWBvlulpMvHtKFx52VABUSEIOCigXrQCoN3TH4i4Ba2mhqwVwb
Aw8C7BxkEMy8bbxLyQ9109q1tL7cys3Sf3E+CTe4sOGAniiwFrEb9cBQN8XcxExJlXnI6sh8EDTk
SsOnkUUV2IjqaEt90Nit9662TO5ZaDcnPr4GTWQUJpFK3GkhlcxpRWVQBkTLD+co+6RIA5aOYsxi
qzA3VFyOcLS7mT0SIG7+YNQxZ8fWmmiNHbx9SebXua+tbpCI8wK8uZHI++rhBKYDFBUT+zaYbQRg
b/FY7kXwnpqrrO3WJBi3wOnI/xSBLBIi3aejUqqVhdXZ8N3rHLe7vUtK3xKQaKVF7kfqGMvQaQc3
i9wf2INx2C1j8bCH/sNxoXbbiCYFjx6y1Nmj0FL5cLvVzZjoQkE3HwPEAPKznXuM3oGNZtj5xslV
FVNeK2TlMAIs41swt1hpWt+g0Q7cILpjFOtk3TmcVFihLPViLQX3910Vw3iTTOj7CYLfzYqVw6Rf
9IpTDgagRjos9iwp/h0rE0pJSrMALmqOPbDPOJmZZ+NXcu1AhNynzO2mnchveSv72BXG876phWb3
VeEYw9m7s74SbpBnabjIZoxD6vawiA3UUwpcrFTrtTc3tovA0N7c2eHot8zgO0q9eNZv99i2poFt
w9WkC2dZWydI2qOtNtuxm3Zjdg9DeBcouyp4tW8VrE7zX9TS/YKQlxAf8m76tH7IEWOYo3xazJOI
7w2oLfxL2rLJd6M+kad2lBfmrUlQTDiZtIlXpIrw4pIOhsLnM2BPzsCPG7GDoDNvXQfB9DxkEA9J
2eSFz4s/xDk7ghAHHk3/0s8K40VJaptHkuGBj+gq1+9htJt+GfjL+xJwZOlVuNVHOERaia3Vg/aj
63G+7ljwFrdmofWvR9Ds3ZFUUGFTU4yHQHWoqd849K6uqilS7LamhOEe91e64Uxr+pULkjEUsQPd
IxzdwCxPfkePOyihWrbeUYtgBaYtKEOOhyqoqoNIvKhLENPtCQT/3xJ1JOiaEYhagSxgSyWFvHu7
GOKKPN6Bbm30nVfHAJlD9IyJvWUI4AhBUHQn2/l61iq4EUag0rw7k7q5drD7qCEXAmGXkZmlhvJO
13hCUFC6fGZptKJrs/x/IazUnIT972nTXeF81jXtA+2Kw1JWdm7VBpM0g4zKEMVZJjBohFxvv+Jg
+gqc9Yfx/iN3XLHUOemOBxeH7vlu7OT3nH7wKNlGahzutzPkywuKNj73QPWnnGZ661V4Ep2OOfVV
of65b2ymNk1IsWZFSt25lSMYu/8ENg1eimZvc30FA6RlIaElo8vTQV1t+ReMCYd8FYaCVfFtf9VO
p0XKUfzvZlx7MMMdfGqU9BtMm+YHL1LLBEMHxDG0dkFm5/2w7m/WdLmktMI2rcNpPY4FYrVfu5pp
7heyNIOy9fDJRikiz2Leym1hWNpGtOrYKsMciRYU3tTdPjEHAg+5r7kPahMAxqbTB6HKGkmUpWqD
mMHC9NSjlOtb9dWm1dkaqUveIcq6RjbGMvwjgvVw+FhEUBFl21IRznmqgJfpjx4NZH7IQDZYBK7R
mKClYlf0d1jtB4GKsh/GgCvfL720CE8mYhGLne7oRX/xrhYqPMB+nIbfVlosSnqYGNJasRZsV9pD
uqEm7zRwjjqStBd/qiEB+Tl7071mvbU5WJZlzI9zaeHfTEy3Ox9zJfFhofQQhPmh5jC+TrKmSMsv
GcSyDM9EV1oTJM6FIVJAGvapjvNLqa1LwcaV5WgxwiOMxrKbDkpu5d6sYwkz0NlbFDu+hV+RG5y9
MqQw6pfe7DladnBXr05qolKKnSEZTB5kI65T47UPes9J5Tf/Y/YGCe+c2U7yBs+4CKNQkYSFFlSu
mVhdrKrU8pBjnsBvIJzV6zvthBAK7LnREgagA4SU4ttgggOkpmoa7qfNIvuxhqDS81MdVKJ3ybKs
MT6fZlRJVrldk2MupWcm98qef3DYxcYqIRH+vQm1C0q5sO+t5EYAExl2KK112kSPQJ1CKtVAbMzf
5KIuERNqmIO6NFouq7se46CUywPuUjPzKSF+gI2BswRKF3ajYobs6sC8Y7SigzobnrWUeWseZDtP
PzjtEfy//cXcVn/VL1tkJoIfVHkZUL52nS7IhnIXz3vmttq8V3zaglZsMpcjh/lxwD7KRcHJHp8j
nwW7EFiUgtePUYtaUu/uL+rWoLE9yGKXcXoOZIO0w4RM0lDm6ZtFo3m7j+7Rykyot36ISsn/yUbZ
qPI5BpSomzcrmdOfWGoztQfbGyXEDFx6ntSliPYd19bQYuIzsmQe0FUg0FOU/MaBdP0F99AD/FUm
IyfuspYuMFc2tIyUIb9jrIRkzxcRbhk/5qOp6VWfhhqSpnWgOyA1siZ1+K4LiO24SqGHMF7uJ9N/
sapzrwBktUfPe9NXUKJ32UFlisnIKH6HUv4uRJ+6TY5MPNx5Y3zV61nBRTPlY9Jd7+l2fkz81Yvi
n2xJJxQXBkW1ZL+5ukK581spc4K8U6HyiUu4Q+uYhiGVcg8nBQj/EBAUe00AdQa1/pPvvG0OkR49
CyfSa7ZJwszhmAR4J1Eg9medWO4LwQC6SkuP/Nu+211ofPefntfmiMNlMn5hMUy3wjQ83XAPlRBT
BiZkzdyDsUwWChsrw79j+qWuzvktRyhfk1UVnDGObBXlkem+bb/UmQ96ZgY94mgV+R+BicNRS7hL
5u8ZkYATXa07z9o4MdWIkIjHKbAnZ7do9dnMDmB4kwCzawIxoyhUWBEZ9F+7XsfzhGNKPvLGIXZH
UgQ70ToimFfJXwuoUysvC/QRSeF/NOhcMBkBlbx8YFz8czaniFL/lwkf0sTBD2JEHZrEDsFbPFWX
7BmtUsKVsbF3w3FfprktOXKMPMMDYbPeU2zAFRIV7V42yzvphPWUt1W0gHUcdPMBFzCB6xNOjWmW
xN2ZnEwAeTnuiC0PObHqkCn6vY0e8VUMYvuArYcIfzBxlrIpXo1rSP2ME2/mdpUlMfk/woC2wqj0
t5iwGZCpLoGhOettR9JK9Vm5HsEHNhRp1zSwg0EuM+NWhJlC4xLOxeuir+JbUIkAO8e5AqYqfJtA
P4U450KXVyVz0vo+Pwps3Nxc5NNYxf551P8c/tZUCKtaxug5vxA1AKuoWNjkMCssLzZhm5SZ9A4q
UoUPNIWWU8ICoLwMZHoSt/Du5lFJG2CSs1Bz34nlboV8Tg+O4rFYpbyx2nv38Vs67KNQMq3oQEBr
7tcqQ9HccCnxMJhccH8Ezb6+sbrJ4wOXL8wEi8KZKh9Wj96Hql3GUe/AwSA66SjUQgu5owF4rva8
YS8xxaiXqcewcx1FC0+GBipk1cMbLHftzM1N5TzUWP65oZfd85EAEi1Z5nIB8+PH3FY92orC7h8Y
yoOxfR7ThCoYcq4KfeBPAya+glVcjJntLynDKnu2NHpvPNIDfzmvJVM6Gb8pRDfARF79KjV0KV2W
ObG+k1mIXotGcRzNKdAuDu7fO34uAVefdX/4LB6BrQDgy1lKySsp1lT8MhRPth4aw7jQyOP+uTzz
8zYIPJvo9SvoSnxjNIS8dHRW7D0y5Gf9EAPluouPzuhwtF2UxDuOvkjgU2dDmvvyfFd5yiLffAfu
r0Kh7CxkMMZrm2E47qH/eb9CaIKMhQvG+AlYyGaOIzoE8u/LJMu/9fXsiWBG6qeVXjKWQRirNBoL
V9/yCDS5+YVRG4DikQda5/NGZ3U84mthRHi3o0c6xyHEcK5Np8Btxrjb5bPAwVcRCWlSXxUzGM0P
jcx3zQeKkuMpxbWkqkKdrSCrnfefECncK4yizUIvHPB8A5qXI8PI1tfC51d/ufIpB8azmXlirqGe
DMrCuJp53l6K/e/8rvOHqRQ82kreVORuCsVfDRsmN2mpnTriCc6Ixhcz80u+nTURxDGbFaO9lFn8
cprUwO1/7Slzoh9qUxpRxp+sIuZTe4I+nfpPZ2WepRekPyckydJI4UrceoLfNDDbPKnIOr4GGzcn
4+NhfjpTvcmF/1C7E5vnnBeDW3HPEabJ9/jE86FOMcgXLUVOoy9GmSuQvJm2O82VLPL46LI5snev
YoJRk2ZySlxM2TmUGt30hqQwkaZ803DaGqerZDVMcN/oF5e83mHtfidLhKpwZolu7iGhFgubK84Q
qGbXTkpImbPyBL8VkG6whWVfwEXhqf7TbC3CWpB2bmbdd80PeXGY1L0yzJunJw8zvQB4X17d555n
TGm9Qlh9IVE+QxrOaVmpqL6Y8aRkI57K5VKjKwDKwQyKmOtI2nrFD+O5Z5bAt85/9s3pHmDHAV4U
LRkqpoKGwq4tIoyFxGHFR5Lc1n3dvDk7OU+i0RnSzdbns76Rk5FGMVPClj6Qa6kRzabmi+nq6jvA
0p8NfdchBspJt/nEOwpQ/IuMHIfjvA6h1VQ1YlAJ5Ton9TsirV6kZy2NmiXx2+PXf3bwnZ+3tGZe
eeFh3oTJViiUUXlgiSYOPIdyRvyASweKe6KADIiKv+c3WZxQcvFbAXSo1WYTQqZCjYdZDZUb2EUe
mKvfbvLHSVZ58qbr/u88dQukNfCySwiPdddbXiEopuHc4mBFkVwR2PH4uqfwCmZvCM+5GIwZQoS2
sJwqqtTwueV+jco0g6N2jzumNvHI3kuRpRJsuNPHvzAaxeOhY0YWx+CeQQSRvoMNSN5kPTAaE50a
TCuNehM0f3SJBLLZai1YZR8BLmwXwm/tN3Wn/ghNGLqeBI5yGFh/NrDHmo5o6AaP2Gwnkwqy0ypc
9EK/ynp1ox0UhoRZ1+nZt6giTXIE0wQw5B5/v2U5Zo6Um5hG9mfKsH8HWRK479GKSaU7bPHB1CQt
EwKaj7LGhk5LjBrYnILxcVyObQtL7Sa1Pb9VedXupvqxr7bc0LgsJlsli9vfOvpEOUmSFmAiKHoC
bB8FS6WqktYqUB419O/2PBrhIMG4r7fKHsxdw0vpuDNX+eAs3WsLKuEho6M9y1cTWsvMOa52BOsS
BqcvtD92ZtJy3d3iMaYoHL5sdlj3/wrzvvf3X9xPVfAXwyvzxI8UT8Ptusm8IXDNo8/sTbevQh/5
l5zJFbWA0rRMXlzmBBAT7S7i9PUhUjy9yZBxvPm/LuDrmej8Gr9ww9MUELcgs87cWWWMcr3uYT5X
sU2CiHgyz4aiEBb35IuGiYmQalJGDL9THOWmpqnd7Jsb6UWHmdPVMP2Q1VurrdWYI9OMDGwO5SJL
a1ll5b0YzSsjDEkOaMOWl5hPDbQdpHD5YAw+1mAXsZXeaodWka4ooX1GMxeDejbhv3K2S+IUrmqv
cKlwIKMVdRsjXfmWzEiSa9qHDePlsvCRKx2xro0K08k3OLPo0k4UGk1XHrqzgfpNELSoxhIFkSpZ
ZARMFzBMbkzMpgJwsrcdTeQiKB4mkI0m05RGDurRy55mrOFrt2+eoSyULVCL9gvb/OsoSZ10Ai4e
F3SztoBACkq1glmEESFVPgHoFclZJvtXvBXVzHQj+v4EAsoXP6FHaWV7CQoJvc+9Li1K/+WC8kER
zcI28YWEjRpZnDXScOnrbRhJ4S3rSuWAADFJ5/sTmRbXbHV2Ad9MnTmkciYEycEPUx97YZjr0XYj
wusNHBkBJU6rxB4YfO6YFSf0p1hgBjS/lvS0JjVSbF0s2EJydJVtO6i47AncRvQdB+G74yy7TlFb
tNmO9DkL+0PIN6KgdAiCWU+Pg3FI1dIzfSZJHIjX5QybcVxyYBku69zn7ugeQ6HZdWncFGAYD/jx
CLPkh4WQLHMuUYABFlCovrdz3+KaUxBV+jumQlVj2QUL4Kc4AU9YcUeMgSQjf1o5HEvn/B1ZGKiK
HI5SjRfMWSOyQs9WMecYzU9dQ5xMw+uCxrpmqa3QWHfu1G0Csg5jqU/CP6VS8kM7jEQjXQgf/I1f
QVfnRzfWRNC+plW23Awla8ZNdB/i0YR1KYv0n9COQQBIkiTO2CdD8SQJqhi/hFL6LHgyM6JqkHL5
TFsQsnCdeiELO6X6tJI+s7t8qNkXBYJ68swezZRPQGJGUnGCa578+WUPFSl41exePYfKYDTn5ian
kueUSYbLhlNAAJ+9RNh3txtjLF1ePnLfThYVgxf8aX66sF86T5PFMObcNxLZY1FxdSeD29NJOmUT
HuLnnhctCpQYtOp97lLzDOZ9j76O9fM+VgYb8HwPgf0YKjEORqS2kE8qRCkL4ufQGGx4bU0+r1Z2
Ozir+GfZCeQSGgAXSOUomdFtSSfqCLO+hZMW4WfRNzfqjBzQMCOzGYjK19HwAv4oVFqDo28sezpD
s865mOxEryBKL15H6NbR1AZShiKni7Tu8iz55y/dip3XTA59sKw6BZWYk2/slk88cOBe1nblbKIS
KbjaSj9qEX4FAwZzt1fCF53R19cNroAXJ7DpW1KEexmEBIIKvERVjkCmqXpORi9giiqJAhOSsnTj
adLgNkXBbViLD62UDS8GslZqpRYacgbi46w7hKe60Zi3hx1MFB7NrzPogiGF4GslUXKCjmeiM9kk
Tq34pcLRbd3hRCJW05WVRqykoideedN7viRQyMUp2yEPrMCeeHI9DFNcqR/qPdlHXjnD5xMo99dE
3ERDdDWrxkUfwdfxbGcy9VrkzPBKpFs3ENt8rJIk8ODAnbc2UYGgzu5YEsuwfCr/PW8algfmjf9c
HUZeo/ne5j5EJEIuWkdrRsl1/t2CAB9Lf5LbCwutbpa4Q5TI7kFQabiKn5mXAyD1xRmpiP++PZuf
Qe3AWtNpON11j3Aj4WJvdhhgULv6Immn8snXX/HavYCFRxR44XkpKYNooi142ld2PmBiffwfi92G
1BUS9YVKkACgB95hSIY3jtZ4Hd50ZXLcokCWYhZa0PLlxLzgorLNWAntPN5AOW3W+kiqaDY7qV6r
+A+k12yVP6ID8aD4ey/J5hs8IRsJJrtlHEB8X2AiW8Sro8XbOk7tzmwYKoEkOM3y0QuH01EBF6bv
EVkbk8doI497/vkcOhAHqaqdpkz7hyxRarNLf3TGELOP2iG7OyDQoCl+RRshacU43GAJnc2AOGHA
uagwliywIS/LC4EUIWfjNxs0+yXN3J1H2yTaZxqkRVNtwmtlQc2Gyn8exYwhx6B4PFw2NFsK9m1n
pNh2EA+xhRWWkBVwxnx0IFRmihz7i6mORK14NXYU42C54sm4aaOLuzGRAx1D7sod+Xuhh24e2tfK
B47OuI39OOG5vluhHN5efTZvmWade/XG7CNXh7ndghB7R/Op14mpDCteWOBDkr5B61RofEs8jqXK
WbXrQXMBiQdr/ozBcCPgi7D0Ej2uQN2+rtmsu7v+FzQOsNcBJJ9LFWvGLLzIcpfZ9kDgLxyZUGFX
V8kF6l/a6sw+n/rlZTJdVTcRhECpZL3LpkegEZmTtxxqrMKRwVrBLvLlLWYINaKmk5ltmAaPvhuB
fRO+n9FbVQkNZRlSHkHYn9rd9WcMKOs0LJkaU2FjAt7DA/vRtJHT0t/SsfkIx4hRI8X2Pc9XF5Nt
A8Lw39QGQYPo5vT0+8huAmwoyhzCrktParQEABz865NSdjEXwovD9w2f80e5bJINuhnhrKCDymGF
Atsy82soMpZ/9X0nv/ge1l2oZXfW/UmdsalYdmySBfWwcATqEoQZ63VKzrhF2K8pXcFg+W0dr8rK
ZC+Y43tyWIE/vNexsQ5tRCtuMrLI8ds3sfvVLuiUC3eGjVSM0+mYOFPBaeflDy3X/R0WA139eNjX
MYiV5GYEQDHWlmEq24GKKcM8GuS3Beql62241oWnQmRDlQpwDa9e3zN/fTXi5F7ECb+VNmJphFUG
Jo89ufxK8BNbUMYpb2VWltSSyjyPDHvygC8EgpstGuqnzbNw7DOrNmLl6+gkzjyoAibfyu9Hhjya
d0PStYpFOGDY6gKkc2Kd0FGtgUVeeU0bVmRtRVOpxX7FLcg/BHCJqtjfFcVBgvKZhIf0LTmYdgci
+evy94s90txvM9+P/zQOoWKiGB42UifWJujWmMjOF2YedAxwi+6fwImxk7uRGaOQak/2WW8jBTk/
NmndIiR3KShmt39Vy8IKSszU+XZwpFyjmUrDRARWWc87nQsV3sdIzfvx1V5Xq7YlIlcuv8Th1Grk
PqlFyRRgnegY+33VObLMSy3NNbJgJV4RfUT9V3VrYlhsYX6B8yGHw2iRfTzvfi7AwAgI1YfyE/5/
kOQmn+ykVoPdm227owjlhz24D/RQLxaulON+Jv9SZynt/w/RUbUf5g94zeib9Uj8UFG/gkCtG5WW
c129EVqaBIC/EtY0BvRPTlz36qtyoJYPHwR02a8yGbVaNBeGNkBmSPTA9stk5PY5vhp20pt615ap
IV7eUCDlrKYU9U9s09XOi+qzKo5WoNeb/rQQ8NZMerRWyGAPOGFaYz4PZn6TDwNDY73+Lj6gt3ay
7CzGiJvAWPYwMhXitoZ4Js7yVEysBNLD5EbiKxiZqUjA3POgMiJC6bFNXsmHU9E2qpY2Bh/Ahi+M
D9/KdnljskcZoXXKU7VP8jw5I84w/FmPvFHBlFKrJbHBVYuMuS1P5kicY0uQZ3yoEOJeYcgFWH2z
SD9abhOEfREHxWSJiiS7OroH0Z9pwh3c2fTHuEkd1ACQXa9WQPiB+o2+gFrsc5lnloHroIwVOP/I
5d9MdLzcu54D60Hcx9OLpDSl0JOqy6YUza8n+1nX4m4eXkWiXhBgRJTh8NBcG30ABToTUKk23uR6
OQFEp9HL5OAlxfQ+uHxeudm7Jrk1P/ZUEpM3O3zo/PTDJ3KCg67sjed0x//KApVD737/JjwF0jYg
bwRGmU087t9POoT8PSIHwnPrZFPP6Ioi6YmJ6HkP92o2PJfcTRMg5Nh9Vb8v4HwDbSf3qASVbxrl
B8VJ3KIzS9D3N+np2n7xBE91DEVhs1zppa0X/ao/Df21YacFPbsRwCyT8Jm7RHrTBbzdWB1aYNay
p713EiIsTu/fI9eTw+bKCnuIdELUDmcqQ0EcvowpJMRejshz48VKxoqO372oyYdnEat6I0DkiexR
xCEbMzJP+UAEuap6MLW7MYN/zVGb8fOHKRzi7mSBi5I1tpRjcwRaqcgKizqkhOkyeGFaRPT3NuIx
2X2C1Chsn+9V+PVT5xRhLlZD6+/nDwFNhAesqGFCzAYrGP7kMzoJdcx2/55wKixZ5amoSczFqvs/
1Kckr40B1urUdvjI+otzSSFjcDDPiLxxePHdaXl6habQf2uIj99pzLPoqcwN5LeQHWC3rqdar1ca
P800LX/NEoOWJgCRbOpVzviXdkWUn8XUiUnhlf9uyRgJdYNufkd994blPvbWNBpoZPjxX/EcXoJj
QxsjX4SxDWXB64MDKIpDBYkY2YrVARYwPkFIhzJiDKIM7WUH+GUGyE6Vz+bI2Djlxy6z5K3a2tH5
p4HXhMY7PDCduQOuHsX+IqeM6cxn8hGl6dWSXPey5ZENLkywBz+1rbkwdgpuhtD77tezlyErKVlU
hQh3Uwpynnwenlj9+VIrjuOITx2gL2cRd0MJmvPjS5UVOZ9wkf5/eCgs0Th+19DmlwHqm/khSBF/
S+mZtG7U88bRTvA/b+tAePboar5zEUvgvhRIzt7fmmvQcFrYXsT8ndxsSLPd+knZzUwRC4jjdT8A
uObkzLgIjGzkxF/OmY6tLYOsKRm9yu2O9028byJIINSTtVH1XVrqceQWrmpMwZjmrK3msebsdED6
jvtjBhAz/05/o4CHT7FeGQmtnVmj95e39Y8/L6AuPCCCCA5D6Uh+1711GKQWZ1RmOzAANu+OPN3i
PufxaWduKCZjjaUxwDHnUQ8v0l2FJftM9Wj/fpSb2F7vBUYn2PHxjtBHvUWUoW5J2bWMnJVcK13q
Iljoo/wM4ZFw0ss66AyXKuqaIcJZATeBobANk6R8zmdkcpL3YByloCIk1hpFqCx13B+1+l6Qrguk
mbojG83mxi2EiWWFdUHOg3UFAAjkMFQA9bCUmGIIjWoECyXbYcH75cTYnMJz4+PSghJc4usfUheX
+g6t3L7DMCS0LmysPlF4KFHOjLG7LaGp7yR030EltmD3HHhCVrKbKjh3+8favwO/9y70lp52sOX4
xFN8zASn/kerAg3j/bGxoTmdgJNnZYVVruSnt8Jf1+nb7Zi+rlrvRtwUjG/B5lr3C+TFUJeHa0MX
z2MOsgKC0elNBd5Ygym6J9bVC9NBgUNKK33R4CbhwN3rHMPdbA5Hvi/IT6W0ekp68NBouED+G2jc
TOO8dKi6FMrEY9IQ1SmKnaNY+weYCWs4QnRHsuZp0S6xfEP/BEhzy7q32dRgmrya6IgKB3uc/Iqb
WrMo8rvZPUlB5IfehBEeTmIc86Hg7M8VOR8++LeSKe+Cz33lnuabSokAMfhkaMkID1RX3T+lWKBX
49txYnwBnjyaOuBjr4TZNr/CBEwnqtpfGyYcJTvsu32EQMppjEU4BqOclTGjrg0OHw5f5CqQqpmZ
GjBWTXzwOGKcEiYuzBvXYj9gVbafDJ8OKDpOrOgJf3zQCrKPqcB08SlfCMCwOEVzPbhi+UouHOhs
hE1KgaMoHqg9TkuxWuYvm5CzyLR7gpAaJ0cH8/ZZwgJQwsptdwM461DILOgdT1hDXx/XKRL7Irqp
L25WdRQJQ/zq70tSnMzhl7ZHM9uzkhJdSffVqyrgiM8CW6yLVCCA5IVEAjX42y2PRXsBZ0/deyID
BVrF/8XrfUgw3kUbX9QYyB9qKijmIyPsrO7l9YwI4dh+F1Jk/r1Fhv9fOtw3nGzAyE+KB16kXB2u
w4jG/1wnzPy4MLmpbxJ4V+1DPuHwddmQtRhuXTQhmSVLPr0ELLaFf5OSaUEvhW0WztfDaQ/vH1xm
l60H5cV5xM5jxoKCmCBPngrWTEOSdsM6U5BNUtS4Qz1JXu1lMMCL3m125NfBGBWNYBBTTSwU1uP6
HkI/RfJuSmVZikXo8b4epxxQsFSR0rGF7mzpvHMno6qRB2cLAfupBQl1A6f3AbWmSeHidN71dxXh
TEtxvZY8cWwHASRcgbCQgTcZ5czAcNGLD2tLMa4m35bDPxw7JZC384yuaypGPG4DMQSpe00A19JJ
Qj1dyDbjDg4r/kaj4hVNR63xFjl4U4Rwnx92k/mZgNO1V55gcu56MpaFRU1zsCrtlGNzezy7aNvH
7QL8a6XshnNBBepQZ8SN9LTPKpzFpRcEH/S3Jkf8G6yyVO+29AcE/UQa2lDeJHQwmyE0eXFPtn0D
hjn/vnNpoJDEYlbvIVpVYSjl6ByiQVQnraAeYlyOgpYWofNjurA/NowNzJNCwoipHkTfIsuEW7qf
bW2lPsS71UlWVpFYWNO9mtiqSYJKNll2p8BrtT69pZtb5py86cFuN5tEW2P4pVkVFQXcy8TpA+rB
a5Qh8gdead1Yk/GnMCDclfK0QfFdeMkY6MdD6r2bz+Q2DD6wZ/HO6g0UZlt0Sg/cqG1NH8oi3HnA
niuxQShiWPLbwv0Pwi+X/mR4diit0McMBBQiTtS/975E5Bp8jxk6T6ze1bA9rCMksA5o8p/yfe3e
W7g/97dx9ojA3NXWXm/BH8JziDqwxfmdzvDU/sABDd55EfrWMjmw5FzQacSWEDOp2/eyeZJ0ziZ2
Z9fKE+MwLP5VUuG1rt+nS4u7qW0wnrZV1CufgKzUPG+IW4h/MKOsMpUjoil9ZgWp2+qIp/CMj0Wr
0dS1o2lQlcF4nAxzzT69NnJ24jBMXmDAIrCG1nZ7XY6B2hKZivpMeuWPUmZPQeL6RRq27/jGRH9z
VWWEGwvm3l4YQbJ+bNk3yuOYaIbf4HW+zNfdrVFdr6/ORfgFBjjs1GfvZTlRP/WJprVm6o1i2YEb
jhJCC0NQ5YLFgHqTftWmi2NZEMdhQymQIye/VhuE/xnZADZXNmLUA2UoBB4Yx4jrqYpcSxlObZIk
2FDslRlR2AspV5SmT6hYJ+FiOvTbOLt5NKANfWrLc0s07ztrJTKTYbGlllCa3RCiTefpmNodJ1xc
Hl1Puw4R49u8fac/O4EabDEgi4/DSF0Pz7es+VBlneRU/G0pPvSO9AMdz2b+ZhJjhx9QoQR9HNDb
w8mWC/p9oMZVJ0k3GW3GDMFg43lGqnzLZy9tdOSFSD8G+1esEQ82qHHGRWbi74d5AUJRVqNYiGtG
gQvN4keQJq6mSCbus5QT6Ar9E2fr+pYtBsTGSZQlm3JxUUy23JLRzAXql8sgnhPggZ8CL2FZCmwM
m5DYCpcORVu3Mi1bs8v+2KzSXMegoncCWAyi1T5E8pghZ9F402PdRGUNvOhol+AT2I8tQFsAIxP6
JBmZgAQUAwG8hgws2Fzc4K7Ws/xkY4BkZFFJKHir4R7LBXlL8CXD1UFoFDdYLrVNu0mrSk//k3QE
l6QoL+ioBP/xR+8xHnV2TlHYCwPHpvDGNbs7wpsisHj+9Hf6YH5tUxScEy85StycLNtvagSRkMAb
Iw8LwTUNVbvkkPweqFmqHK2264AJZbG+FAZh60IGsxWbRSKv/xhA3JofxhlOzTHlGDmj1GuVPGRi
5MtL7pxlsTTwHKv1++AuJYNex1eFVPY/wMv04yy9LRTahETPXaRgcbqmX8cI1+z2Ja/g3EpQqAHy
IZ3NrxGqE7o0OfCh9Ah5BjfRkBpiF8pH3Yn/ldlQFVhtXzkNgdkr7nt8bnf0O3b9gbe2V2rfaTjQ
4mKO4lnWplLl1xibIC76SML23IekeQxf80pYXVfRDZwoE2aP7gQXJc44jsBQGoHznNUbzW/rIvod
9OrplfM44UTkdVqOB+/DaiJhMp0/KfGAXvcDF6yu+PDTgFQJo1c5wD8vIKvtJVa4dQWkrACqxKje
wKFk8fXIOJ7J5Krz6OYFhXwccmvvhIah+v6kxMmCbhgwpbdC75IFaTUtmAuaJ7HGIL4PPRbZqRx5
4CW6NheKZVOIObmh62HIhhLGA3uBfJ9mDE12gGLqNtsbJSD1rTyUeY5RryQTGIjVGmMGUIpMEHTD
JXlPBPO+2uvSV/tMhh055ufxreHzX+OXN9hgP2WWmf4A6JIc8BFn5FnTT0NIb/XQ3g9aFq/8whjO
e5fA9KIGQ22tM4jgHFgPteHOwczhJ4z5JMfoklyhL/1qTyyJUGxOC+fxi30D/UXww0ZF39ZaSh/p
HMdycl1YWfjjkrzL+eowV8ailFuzjm3qrldifbSFaUPYrFnnMe620OPjv7v1JRedpNG6RDjfZwoW
eRrDTAhAFIUsJiEXBgzliwWwd0MQdSav4uHYEsFtrYHN4U9z9gB1OImY5jxxir3T12pugkZrlNNW
C7TO/NcA8nhVWbgNt+vOtdhX4iXeXh41oXOz0RBqQcrvXYRqxnWZQOjKeE5wWqcP5OkwP3sj2k4B
GK3W9VjHSOi1G62KJQtXdfZEUuvqasoBHtuv0J2jx5BN0n2yvQhDYQK2soLUEKg0ye4dSx7jNuru
XypHiGRdL7Q0Zat+B77WSrgMboMujWF/J8gYu3vIfdtNLXqmeicSRR4lohRe/cgkddlMYWjxgC5E
0bGxZ+whqN0O/DvhXNnCDK0Rz1cTQ/z4W+evUi6c20eTBGc4UQkn0yjtSNdi8Pe0Uo6s80q7Yav1
tyCdtFX9607Q/BbpuFL92EJ4uFFHzBsboKf9DDbvm4y3NRAl59y9rCXVYCR+Mm+E9ko8Kp5wwzoL
t3zmW5F3QVZGVmRAf8EfB7fPAJ6z0AtLpZ3Msmwgok0GWoaV4233FOH7WJRGxvOwX8g/HJB2umyU
pr0JhEJcvKkko8rTiw05uSPf7qWIpZwGx3teKfdaBhAXUT2OKURavv/GZSwTXC1VApn8HxGjkq9U
lNjcaLFJJRtXNPLhWodo4DxqONyFbvVoVg/QpBfcYFGfnL6gteBvWv+HuaBDBReU6oNhb8egrUFf
zy2E6r8U+eagFWh7DZReFjRi8h8iZu3Ek4dey/0uJjBTxqxN6l9DdwkYvexSrWfnsrsUsTwHzjwb
SJ2KXHm7VYaX9XMZGRGuP/+hW8DyMmLPpCyxTDBfqO5bpbzvgjpdq5oX56bhy6sMr6aN3nhD/l6R
gN0YmEA8EtvsV8Gepm3XRC452VfvhEyPs95EwfGlRGSY3s21uGJsUtrmvHCI/k4j9HDiHt9kLUjw
ra1hyXyDe91a7lV/to5T1xf6c+Zh7OSkafLFv50eV6QDbCpPUoaBiNxOAIlMjj44Nwrj4FgXcu7g
ZfroKWOCQ1059s91sgjQuEVxIuTMWp6IHq7B1ditUVm5WeQU6JMbYVBEm+/seHXGXl0DGlcUiRce
4cHPeZV/9oFli3zOmUWtOPXJGTxV5insDwnX+AZ4jlcz9+IEHBlzrR8UEgazWUc5g1yDX5QhxAsD
rGQGsxLpG5ULYx4alGLx/+HHHRxoUoti3IY4zcCgSwwC3nxp2ptC8zz2cdo1YkOLLSDuPsTEF8Py
9AeleCkHyayRCwUz7hFs2GW6cmiCLBXHT3GsMsIzlmBrir7DO0E/yymZ1gQ0WOwpIQzQsEvaSfvr
GjMpsJP2S2j5lpNaVcqm8cClRwrmvmfRoxZiNQcdE+IESSFTUZmoM8cT6WNbivuiIwgu77wa/bYU
0sZ7wgqcJz56iYjThxDzUfcO2Kv624l1dRKbKnHkATRpVonk3RbtWm0TDOsOTsheZNjQuZ8GzmZK
rDLGGI+jxK8EuyvhqDZErNPh4fUXWsy9N/hxnP7uhnm/2VcwRbfIsCNWLbjwLpR+OcR38qYEbUPY
GIhlSNBbndKh0h9G/MHVsWdZIVNY3olKk5+ykQ55qQ3DjK9QRhJue5LBRri/okXagSmyi0HRDDyG
IkQXETauuGmsSs44thUlF2kbn4psvfuiResVHysvSDTRfctPrxRXPsiQodVImXJS3JUXbFeA4Hwi
Oqu+DCtkDp7ylUHL15Hm+83yD3YJpLGPn1Z61SjQLjN4Yu8NIqDwNhCUQsEtpsqQz88+tK1bie7R
rgRNK/5zGRKm5Cl/pCCy2ZlAN32zzVr2a/b8Or5NSgB8tvabT5eaI1h0LXD33OjMWYO9PzCXgvnM
1Ip0GOIy/ipP3+oTCgDIkQyYkGdbBB1cpPdGYjw6Bl2nDBv0wCAdS6WTjwfMTFn0Pv/cY+SYkIuY
HKtbjgRMwTs/4uNFQ0cxGoIRu83zsSXPSxu84VxHXWE8TuuVTZHqahQqtqol2c50UX+Q4tF4B4nj
EOeQmn0MOkbt4HRdbsoaoVE/4iIDgzkArS20BfiF04xFmFMH4udzPTZM/YVp+gqJ2aU+L1Z8/oFm
RRNl+BCEdAn9DPQ7oam2yzchivorAmPysiApcdTjlNfHC7+NFoxOli3SMR9Pc+MqoxyOeoJds1dJ
5ruvOUWueDbWHlwMZXYXW5dSY69meFctLe7g2qJIueS4Ph15RrKAUDfnSe6u92WSsiu05NAl+861
z+0kduQRjucPY3A+l93Fyei3D1cnHYyRi7I0d7ExjnH9SoDKr/2G3FT5u1LiFM63jvCJ5HtFpmhg
avJS47H2eK1FRuARFFq/h4ef9qLs3CpjTg8ZgtSzMqBkDM7zY2i9bAh62gEsEMG/Wn2NJEGSBct/
KBDiy0mGzYxFR4Hl4ZCJ/kVIA2UOAr0C7XuU9Ka6KhRMxnAVHBlBtbR6aHwmEAXaKbQhGdQGnQuU
4XInP5XeRRteMaxlGW9/5l4XIYRXktovxToqtjukaJ/n9rYYjJAYn+U/XqkX4o3zpAZFt/Oh9bvk
yAGaoG8+lhidyp94XfXI0sXr7YuTl9J6hJgUv2y0PwkQHGLS6DWuY7KBGiA/SmTlkUM3TbVJfI5l
UlrouzwQlIek1MrmsYw7ttVGCL1NCyZt6kJK3bN9zbvY6eZshKI3fl6DsCBlr8vA9BXGRDtH+5ba
e6C7D6m+iHd+DznmNsNJqKaafYmP2ggLGLbzFanByi1pqd0SkiZbzFNfZ08uzAQOzySiH5O+adyU
l46aEutHjo+itld8q8HbJYkYIwbAypt5d2ueswhUQyz4dp93JNjp1nLT2EPwaw9wFEcO+uhfqPAP
qfQtjnfGU0CFVKUQTUQ3m2Ro2JQTKIQkFle5ITVTp2kFpPtoXGXD933W3zqEHVkPCdDmIFuX3U8A
dy8cWWplAg8CFYj88vQacLUziFHm6FpO6hYm1lkYR05sJfRM7ks+o0Xe82itWoSaJhXQdFhIOgkn
AuNXctMOO05vXCKg5wCu4QHGcKpmZs6M9Ob1xenm4JQT+jQT09DfmpFpJC1VhUScG9IOllZUoKd4
pmcaEoN6gkzTBap9gsL+3OeT834TrknYF9ff1X+Q/ZsnxcDBgwHcJ7568x6RzEkR4VSmikXAMRLZ
FQ31EJFlKOwAeMBA9qYe1jRlg3+e3DNUx8Yt7gGbhJjrsj+H6kAEyyDjzyNMJClavKedLuyUxMka
S2PnWrg2VmxN/MlKrCo8wEnAPgSXjmg94g104s2qnBVqDzMA98KH45ZLjtKaH6v6ozihYxz0FegE
3YNHWkSRsH+p3o3NhUFx0ImeiBTdlTy6T7eRGHgs9yyFxg7ytVTi9xr0jchP79U4At/J1vQITOTf
PVSK5KGar3sv48byHPac/FxupceB76yi2I/QER94WJZ4DAwtQfpFfV+o74mOr5L+bgiDVaZ0NLyI
tFxqU0E+5vhU74xNdW8gO0G0lZm1IOcqEU7SdxS1tauWeHeC9VNg7bgeWZfiRc8JI9pu9iEDvn5C
iWByggWiff0kb+iwCw2WcoYuURFyKAAEjA/D9YPcOsHz8LluGyzC0Lp5Y+fsE7DWB8MWgGq2SDJ1
oORtNUilzbVambC3wmeL0pF+PKV3M7oLp8w3awZygUfuR+ciiPgAV+Vlm+YyrNpzJf9LflqLgHvN
JjdjKg2Iv2hFmHxbeiDtbVYFy3W9gZnwkdVPRt+9Kx0goOb6w392eKEp1dNtYXDspdAW4S+vcw60
IUzCeTBiqaN4uoXy8dclYSW6UJ4ZRNdbLgpS+QNZ9gP9E5PvNko8vDk7BXMe3+NXU1u//8te+gSb
Sv3MusEuOG2OCKwNLlUZV6fGO4oYktQtxbEIIuZWLuR7bVksHlzAegC/nx4WKWYWLslf1DfaOyVd
4DUxJoMb5ucjVJiLoYduhKdc/D5HypUdPTbx+Hb2kiJ8+FD2KtvdT99J0uVn43VCcD8BJGLpdG+8
TzZI9KCndTi/C0B4Wmv99iIwG1j87o4aEAJh1XQhwOsnFYK8n5O5GpmI11rmZI+MXyFbLWibOSaF
WGnCT8wqgqPDlGKYnJBzFhq5/Sc+98YS65E77/yq/9ehhwbdL+tdIpSGd1ylDBh0xXXe28+1g2zr
ZQmqPzFHOAZpcL93OP7djsvd/Cmxl+55F8juZWQ1TMHZU8r21PRCpDe4FxMidHqwS1PjcO1pzL/r
qc4v/O3sHAZnrMvVdiHqSPKHEi9yq9muwLEgkAfqlez1QhwNwBd+cRSymRblPVcUWxkcs1xhl+7l
PkVBp/B94X7XkYzVMM1IYTuhws6K+za9InG8AbhSZhIjYHNpxlcexBSej65/QfMjJ8pqpceC3+WE
nnupWL48TMj6Cuvaw1hGRN5kbAP/+wBlpOxcLWAFM8dVblH9yE6nQlSUNCiAYZV59CdYYhw/2XDn
CvHryUWh3MrJ65YtdT0JvI7uyGv35la/kFEgCIFOsVh87IUpIqlB/FBDtKJtR6oXhhclrtXZd4NB
8xy3pLTXAOTxSo82E25EJa084+ikHvHJW3omn9R2eYd5qmXntodNafN+WKxUaQFZ0zxPcBRRf+m4
UCVGh/ZUU2vqgkqlovvrxk6Hu5OtQ/EHLDDtTcXgFKedghm9O/acXb/X2utOqh0aT4w9UTUgxe4X
+REqLOkkWih5u3TVClANalbBU3CYijxRIdF+qW9XJEmyC/v1vbD1JZ0b0jhRYXplYrtLFvJJpQbZ
FRcI8u3xUSmU1T6Ngo7NrLPLNiZK/2wz3O6qEnsPLBKZDeqHEytnJ5sXihSa/iERCToVTmasSj8C
TbpEuDH3HNTiC7ArKXrvEuAvk4U46Iu1c+PrbJWXpANrmJen6ppPgM3Koa/yyuA0/DhSyyc/qlxx
m+rkcnDOSGXBbCkPVH37OmlnHF4aviA0kNzGaDpfmDhfduwqby55l2YjYNpmu2MRFdDcsVAEYpqB
u9hhUv8y4X7tkfa6QVzr0lVSh+Ter/QJd8URQTBGPuB/GS6WaI/2sqAC2+DC09l9KMFhVuZXKO7C
3xlqkhKLa5xSPCf0ax7Jku7yM+p7oN8n/krWXoqRVVWH6ydRJ0RAwiFT0xhLYtCCkhAG9KdEU8jE
VTvACuKF2i6lB8a/0wzqusbCOXDwsdxPPtS3StmJZ0aPba65QTRMwN6XgeVxSSGhkkaJTmb4cg8F
9E8Tmbezgxv3fcQrvRE3At91NcIGuH4kiXMplBEAvWWedF6I5cvM2bDdvjg2Z29w+B8FL0Wj0C02
34kpuO8XsCxiyu6b/UoOwyidm9aXwaBhusGipCGDTyqGwMDyBSMIMHdkPJKmb9wdCSurjbh290ik
fpC7oy+xbsASLf2MJICIzV3unp7AhvdVqsVYI3y8z+0R4jb6vpt5qeRV7yusmy4uynGpCaO6ALxj
xYNV7xbEsKrsyNGtnLcS75rLVVJvcsL7VeqDMJxq1GD2BFMxURUqXPBExGI/flnQ1ce3sOtvPCOV
a1QzHULf7ornhJAPNoIP+GhowR3seVP1n9kaWYZFr1L2T/v1CsyTHWtzseQ/0WPe7omFnmkJUDeo
VnGrtdNdJKmC8uGxU/t9xvsWTl20d/ymuECsKugz/uFOMhpyat1xcXdDJl6Y/VJDwvjEgQF5p9zL
fPf15y3qFRCQ9xgGVOgOvANJcza4QdcMJK24Sy2ckyqCuDh0T1a99eo0ZSwC64PyJtjdoNuxwBIh
6oNi6O0aiMa20WY9GcSIanq+tYgLzp5IF2hni2rYsB5+jzfPqlOY2MekWXS0VAST6KcYFOzgMoGI
n4Hbo6PZE+EbMGyycDKfq3nmO0+AGM33bPB+g/sZHylskTGmfwZyyd3bBtE2R3cftmz9/7SQD83s
5cEk+I3mIVLZ66FG6+c4jOl6uF2ixge37ZQBNSp1kSMK6O5xJj6gnh4wJDqpMR1LIHqDxfeCadQb
xqvVpKgAjxcDqRMkubgm2i2Vwh2+LStCH5G3t7lZMhJJSbkdFZf7JaV/Nh7651U8RPtQMKzXlYdz
Y7aekayPjExC/54BrDCyNYHwlFlfvM7LmofO+jlR/BLHVt052dwiJYvYBMO0dgowl9v+MkHVVFUj
JO6sZSFQvCrWIllDBOFXqQX8sw+q8/yLLq3XRQnUvbOqhmAU5ZTqSjGwQ//6pycBscsLaTcxOhI6
2+lih+NEeT2txD3kkuzMIS4GM8QsefAa7oXDAYTYQ/54UzJMDzgO6xW0VXCxYiZ6aklbD2k6gBVP
fzy/l5ynfdfwYguuV2CRXswhoZjbh8w1SU1QwWAWpXLI4Mb7PikJAkGfE80ev4p9Tdlpk9iFVpmN
hoAdylmHE3AEEfirj9ISUmoluBCs4geGcyDANGFfeQWoyq7LFaEhNGhU+ZUocirCnrgg8GuqGSXI
i1kaTBnm0UG0EvMBBK6R5nT/5xNCT0ZBXCzgTNb4yKmjE43MShgtGtQd+px9hGtyUF4NSyLPoxpP
lfv3N+AQ/knhZ5IAI5Ax2DBGR5fepMTWUUkDLojBx7rvVa7qZm3M4Giy5BM9S2Q2x4bNAEZys9Xg
+U6P0YmK0SOWBkGpJ5z7tB7lfDJVe6HcrJX1hIvcdSrFrWDsn4qe+vh0wFnrut4YNtHEdiP0sctK
aujrCG+AbLNdIodhjOKAaNn8hTc5E8OAiaHVPe1Id8/2q+Se3z/b899YGESMVrRz/frHpCcdTMm+
1lJRSI1Bv9Ma9eTVPS1ZCH+Ksa76/wFkmfTL1bq7QiXHkGt/UXoxXbheALQU3vI8giZGeS0MdPCh
iV0hW/emAkQ5fRsVGjVMT+ok1SDmiwID+59kUZuj3byB5cx+i75FzJyGgq3xa8yfsqKTl6Nj2aeu
WkkHt6+I8Rv0R0Gm1poPyv9R27rg5E1BxMxXaTjoq3nrsWbXwNd5t94NuEubLVeTHdymxhX2XBBu
nfCh5FBlbBnfIZmPsuVCfF81mSIeccECEC4z8pkkDlNDlf7piPjDijRnCoi/ywzy80zcnUf2eeVd
LX8OvFT7dNKbupVA1mLhO5uuxA59DMXWVeRSeJz6xFPv9RZtlqKZAFLl7NYc2AuXpqK0NFaSqCFJ
XACtnxbP30zEMra68oMemE7BHQNPtrz67AuVq15alM2WYBKFDT4woj1V5Hl80tpjkOQAJt3WUGLb
mDck6JEAYItCPQUDTCM1UrAPYKvMv2ji2ioLbHPieZloB45gyJHyjrIESaIzV1P6ZruOfJS3Sh2X
6R+zMML3eK42fsjE10Ggw0t2GbhOVRW2pWDAkIdtCnyru6+XT7+yzQhKA3baZh9neNUU6lS7da2T
JYgmPpuhacOizkqWzN9ZX56FhLh67YAk7EB3hoTTaItIqgTW/tYyYpOxKX9EtJFClRXxz9RZYdA4
+kpRJuO/VSel6xm4nn1vIYcdXqvfoEIB5C8/9lXgkJgjEtlp19HIhjqW/r48HGuh25w1c6Fdynsp
tLy3MlVTegxwryvp+FvDZvzWXer2aRDnFEmE3aekXsfnFjP+rGnQ10kE4r+LHRNzXhLsnQT+pKTS
DgGgNER5x+4V+y9OVQpqMTvK7/7MWjI36jZFIpuVnlBPeaEZrIyjibkLYQAc7ulG9LjekeQ8un0L
T3Is8yS2g4UE2kqH67VU56w8wp6atChO8MGQlD0Ci2H0PyPU7RgWJo5upUogFDgce4u/Tm3NnYdk
5/CTnvLlaFYsJR8fEbq7G4eGQpx8RAFQvHtMiylKUrLb/fKEZFcMMvVFpJ+EhRhJfos65Z8XDf5w
MhRg8asn9bz3hVhFmoJmVx2/v3+bK6FsTXcW6WW/sPug1qaver3XMpmm7AOuXHs1Z6jQ1FH3ktSt
t8eBNLGyiV5zAGaW1MmOeUM7dpiZIjpwAuaxoZtd146Rf+z3jdwn7Udo5+gU85HghTAu75SIafXM
OqQC0YCtObZrA5LjoPhs/CCErNVlDbVW+wNrBSDkh91/nZMkYzUgA6EFMuzUD00FeVlFPRsfoYcV
b9/Y0EGEbDGQwpwVNABFHR8bicKjFDnRr92agjQHM3gBb8jigH/A/kky61krsh6hIAMRVJPsFUWb
tKeKs3tmFFpUbZoyoZiaj7BQy+YeuLPuQkaKJD1YLR1gHeTYSs8a7OoBFAwfyIBUEcyVKAUT95v5
rC8gkl0kgIHwo1bc5K8mNk05dtqT0a6Od8tUSqxGtxrKRlmsb2WdS2B7LWP3kexXc7pK5UbERagm
tNLqyncjYl6q5vSOhaz7hXiIuXsMinWFnXz2a+9c7E8diaoSJ68g48dGpvL9tmrGtB4mf0yQNJgx
8syzWgdf73pbkUHreVzi+QNOLAll57Oq+mgaAKv6lXPz+Ywvu1cAMQZ37OTSqal5Brry2WL7G5XO
u/LeKb6l7U8mAXIyrj+aPVpexfo5QMZfjSdRQxT8MwuMU36HvOx9SXPKypwkWnt+WeJn476Q1bKL
gGO3VcxVICCtwgwI8pa8mS75Cy2RXtJr+KoYCyhy61+2tJVDFsmIsQzaWESQl2aQ0W4o53fFnOyO
qmRqXdr7OFOFYR320w17chc7ItkLuvoyD3CQX/42zOgkhjxHokr4xVhm4GVAAVoDHp61CS7bA7H0
MnC5s5Fn0MJsY+zcljncfDu1H5p5NNBrNThgloan+vjPj5nXjaaYT1lOV+2++7Ee5QDxWrxis9i0
GF1txo2qxWHcWbcaVyyx59WUanUCQlcqM+TcD3YCyE53keQVMWaAkk6AY18e1oTycffEyr7DmigX
ExM+smfMn1jP2C6KSx4b0M38cwzCKfkpxWhq5EWLBqSKj+aMK4X/69O32P3LJRQLEDPhUe8NFR7D
P/j3Y+Caw0okYkS/8nStMRpEl80PM/2YNdEuKSl6+dpXtpoj15gDazKjTyHceWUr75T26NChpgCf
aU120xdT6DP6flXQhcGl7gnSTjBsbr9HJlP1YxsxMuHVdM+1lTzkGodQDafNnDQJs1m8VLd/10Sq
hykYTM30fljgkL4b5gO0J0T9dRMXu5KURWF/GV3+4WKwNnYOL3v2ToecFiHwkvC+Njiddu77FuJK
nxsNKhKYsYmlA3JvkYkS01Iywj+lfN7SCxddBiJ5XSH+TMU3rso7jrQ6xVW8F+rz/8zHfHdvfOR0
GomFudsiXpGbHKE4embfno5AdiWF10JelohRCUjHN5+5u8xSHWTqss+oZ1RCZEaE06tHpuDMLvc+
OmNeHak6stFwVev2tMiW9FNd/1twEFDIeQOIFFpS6xeGlL02TGiL6ojIeqNbsvNDRZFlQNGQD/zq
PMFNKlEq8DyQtK/2ufqP9iawC6WR4zrNumgZ+bE6Ni8zTT3uWNSyzE7WiG+iX0cM7Z+l4CmZ0UPz
tZ+zUsqaEFcBV5oEN2AEFfyRhfJ6VHW28oUCa4sYLXPAcYn4p4s92xrobChn5X6lS7OAKx1QCqoK
CJIcZqoIsenFYrBI3sK/AcNAFFjjZ/rsi7by+DltULklZa9C3iK6q1GfHDnZ+rZtvR715csJuM15
h4DyHguiQc7sCG6dqE4tEqnNMqUFGxz26pd1sF2GtG0hC614SVO5hKINIryRNrGMPO6yitrKSDeP
m4o1Z9iEVU/kmmT+Ny1dzqCTY57Qyhvq33oCERXoRuVWPT63JIlyDcpgJWb3960iCa+8vqd12QcT
tvA/ieTtSfO5hZ6G/GnA2ytbrAx6Hu4ilVpLGZ7vnh0U61gJCR7dlFlDSknhprfKELzNgUjw9dyp
a3M5ie5jUwsWFSeVB2wUncsyznSxhiGYjvhiQUzE+Lj0zs3yB/Emzb4emal9E9AsBhvuvp2Hi8AQ
GnS1WZxk76sIRJ5T3wA18g9t9hXByviklWtdZXyP8UcYhOZ7FEr3J5UNWS8Afkn9Df0a6mpzB7B6
P/Sx0kE3kD5B45RHQWBbRzI0SAC1xkOh9qVHvhV7r6biAdRe/qBVrhVmg6d7gFTrmoTYDezlzVaK
866aH1kvkzCeKH6iDdh8HuPqDtY+X0+Xm9BC5Z+RP5aB6yHL4FWDWqFFDs/WyB1U1waKmoxUP+d3
jW5yfBcU5j+y8shHAzpT04ZHsd/9E2Hs8luXKdpW2JNiZB0DZtWTOf/PatFoAllGIOnTkq5ZcXfP
GKRYO/c5yWxHHRunEgNYx/C2tmP4IQPdw8bC3OuCI6twhUQGhfU4D/2MhQZNMK9ty8L+KhdKDQIj
5NkL2qagLQw/C6Goa5ahDY6N4U623yYAusbH1+//Y+JLGCBZmQGBGZqcfcoQHnfJjJ66AD5hvfIg
IJnUTipOoLFR4bQLU7ow09LG0gMwbmJa7iXHBB5kcQ3jzQCEW0SaJ9/AaPNzjQdGoVglemnh59r7
vXU78t/kk/dywCDaoCcGn1H6CgbTmp3R0vK5QAt/Un0NcuRpX0hFIFHa1gDWe30t2thVXbfP6V0h
F24hFH3ra31RqU9q0//R8nZfGFCg32uYwsLhSl2XhqQJQZg8gCqYxy5La3jysF9/VpqHyMBRQaZw
P85kSMWJAihO/a5EOWIHawwdpG0ba8ls/SnjGcgMgt7ibMLXVnnbK/1kkEMCuklMqeWwdy/usAzk
mHH1SkREqi8JBCowSdCCIwvtHleQ3lxVoG2OBpUAIv0t5RsqogauCwmVJ4tHaI61SzkPFvIqctti
hUwW8XbCKHHOabWvIGUZjMbf1qcsDwFtohMkEnGs0uHdZ/uZQpxYu8MoyQ3r1cBDHT+gnrCE8q/B
Mw+5DX7mr+zmCc6f+bJ3yuYAWrRlu6LU6cGJgV2/nDteSkcAFQJcarM7SX5pNCn6Cyd1neAVK4E8
Gr0vrAUIQ20MgIqgGLQcYThUlb4SP+jWP8HUeuVZRhQuIYPJs5mvnqi16xWvGYBwgvvfQAjRCm9k
RBbFnrRirGJHqkQvpK8/OWU6jwY28rfWaDY/CdVewINwEOQxd2MNn5E8d8vxpBI1qjJlET3kJ+53
dk4kbEKeFqcN3HNzcFRH1QhlqEYg91lyH74XkWE/aWhTMHbPpi1OZArDDKnjMkA3zi805twkA9vm
+W302K+ZpYXi88Up66xIshBxlKXCOifwOn/QJI7NppZK0A5vBLFv6tisclCHa2cUZhHPeYTMxem2
9VMo3z+CQJflJlC+z6Ld15Zm6COnBsbrxSe/6ZYGp1S+ocikGgOURqzsxIz/iHAve8s6iWMrn3R0
z4SkkEBjBfUuc5hJCatZLviM5dT6vc1pgyb5cMQBGxVmW7rA1wylcTBWb/NOgG8wu5Dn8kRsyZKJ
p9/GweFgPyu4tFI7nMyyBDgbzKOVfkrQE3VgB0i9Lc/8ID0r53Y55hLHMDf/sy07tnSz0jduEQEh
Wgjnzclx4hxK3Jp7AE3GEmJsJnKQOu39AF63w/ys/sugJEckaFgglk2MI7b46n99WmLzLC6I5+hf
alq6FCfprmEavpoulMvpeUBRwr1Zk+AowiNtK1P04GNGaeMBeU1Qat1ON8M85eD9yzndYQG+Oivd
3rzYLJick3OV306F6PaFlltnmC83jFzH7WL8Y16akntxWM5mE27TJWkB1KlQiuS25zMEuXpdGIJB
sv2dtGCiqtS/Ksd67R4SLSduW76xhF3x4kAmUeldaLWsKnZlzQNq0mtp9QPYc/+rEUjiKio0BOYr
VG1f0mwwxz7zWW8c9xivuPAe9Q3E4XWbjRWaWA4OnNwDfl9m0JpOjq1Yo7l9irqPt5V1YiJ/j2Gu
wAG+ioiikBvGXmvSDNS+lk97noV+t4TKso+wcxD5X5h/9tzG+R1/kNV/VNEhd7meYd+QVwLN139c
p1nWcIR86W4bjlY3Yh8UxT1elRZjsfMmLSUFilTw4liEEsghSV4l1BcSb/3kGt9F7uYM3RqVQ1H+
jPKhJVCGyOdF6Hi54n/kWtVunE8pFyecPxV/kNA0SHFxt/PeArANL6xabyPcvYjw2g9J8/RCnucQ
U1ZP3Erl5ljMErdvURFRLDuNTgYGhFE1sngI/taN9bb3EovInTNnvoye9qWJETTd0GSeHn2hU/Vf
TAz4WAKwrTXh3jnfwFayu1ADqeNjVXctlKuD+n8xmLIhKJIayjkQ4SjF9KtjVzQYZ6f2sKO5Emxg
lSY23Wql6uPl2bb2s1nmahBIHtJoflKO5UUpg7sSBC62ga9z/iuZbDoNzK9WfJVBcq3syhdms2SE
PuqrE2byD07lkRj+gbN/LxVA8aEibpfINNgyG7WYXmobwPRAd3LJw3WbQN6HDm3iRJLTfzi73HX6
PUbW6ADX99beQjjuemrg1MYgWma8B/d54RZnHNow5tT0FUxYxp4sHlZZYoA6reFRouqhgq1gGh7I
lkwtqBDgdeaTt+MjXWKQFfHMFIT9g6oj5hT8sDKW1XuWwxaw/ppKzhyPKzcd2SC0QIX9TISUxePS
NyraKQjjOAjpXxfWt58zKXw7p/9R2dU/l+iK6vujJlcapUQRRVWlJNMQajoTMO6o6VYWMB6PxF5H
66PdpNLwdnc7x39PeYPmqSwrhnL+tiYR92kBfJzNIOzAVovnBlV53GvFKSJZayhAyFp3rpP7TJtN
dS1OGdqRmqBtagI23nAGG/VIu6gGkQwleXAPrBfsjKIp+u3mNVWi9ULUvnRF56RYUgsWzS6Mx9eU
Z1EZaezhmyI/1XDXQazWAgi4dWlExj8SUzDsUCPflua4RDjhiiee3ho5Ape7l/PcibMgE2b/CeL4
/Q6tr2T+JKsvU/JR5SgSnf7iNbuR6oJnSNHFqW3f2Nf0sjNxOQ87UqqR590UKGUROQQLkyPKQHR+
PhpCpgnCAqeV+ZQIUimc/tTWIvcgnLJbu88CXh2VwsWQ9m3BwVNGpm+bhmjNhZAIMjIlKPbbyMjO
nQAqiLCMQk1qn+PiOwxgluNp96WI0ndfiqYLEuG4kJ4rvaUgm34xua0stIDvSLOey4+i+XnT9gvw
C1jl18VEVqPWPP8ZmRm4+jg9RVCYYFnQVSDQrtTjaeQpEgsrxRQt/61nRgFm29IjbO9LHv3NtpcS
qdZkBc8d6iTGdHjPI6XVcDShnHiYS42yBeqcfwN7rlQoIOb1Duo3bCE0UwZNfsCzz+xtTY7Va5Iv
urh+aWr/8eubvbvgeP12tiLVfGFVvRND6JnejpHuTFAv0rDSY2DG5LADGb6ZqvdM94VomJaUQvx6
5X3MpgZuiUpHxGqpWNbfqluNxLVwwfC4XQC87wioBH9Y8140HHfCrPWiY0TbhGOTOlqryTK4Fdlu
ad6BqvqSaRtBEPv9AaGM/i3S0hw5qk+uPjDNNWkSYjgx7tb+dzemt9aEyoe0FYh2XUJT8R67Fxag
DkUfzVdwHSwh/suVl6tXlNUayzjpMN/ENKsKzzpSb0WkJ8gf8Srd34LZUTIwKykjUuflDls3Cbn4
BobsIPoA4+CIi9quFEOyi8lnTmb+WCeI3VDtmcZkGFYhYzqb4V/u81ti6q/bkaif19DkmiCaep9O
7016KiRcrhk2mSGKgCQgzlN66IY7O6Fg9JhTJ6RBLTbgENfY8zl+qZCtDPGtcPGLbcuM7P7JiSRW
6wXo+7MZFRGJTk0rYrX9a6B2nTkIvUcnXDxPxXhWndYzBQ4MJK3QdRrZyRIoP9AMGu0wt28ccQQk
DnRWSTOqc847pUobO7Nkwr0+jJy5S+7/0hLiY3cAQOQgzGQLCOa4e5Ac9/RFA2eIV+ME8bBnQW6B
7wItSAtr8TJvOvVACRhhUMa6bRUq6oZECtnAWTtr+bZA1v4SDm5BxaSrq1AQp34g0DMp9In7V3uw
ISr32ibOIPg5jyO3CldT6uEePmZsLx2e5EuKqQowAf4pMBBi5S+Gnkx5J/YwvuzTgsJKu8w7cQKY
Woz4d6zAmC+apjs9AHop/wRz+ToAlTkSKiD7sZ9rk91h0YlDN/puAhKEj6o8aXSBlhumABu9ael1
lD9JCQ+S+waTEePXX5VRlEUuPfeTNSZWI69dHc/8Ag7BWx9FjxE3uQlGbKXNAHPfCXtvxLmXjimL
bM4OwCmDT7OnUlNk+0EXUiNhqswrokfWTh0dQG8W61VqSsOnaYaEA4g4PshMedCw3du/olAvS/tk
HIlPp7ezyF2MVWQCD1aZkBR7EKCKxNjEcECFgc0XnpL0IFtscwh8xMeU7Ul/lKW8IlFl/9l4Cx2m
8Vcvo/A+TF3NWtlrnLLrZU1OMo4HHl6eh3/oRVF4MpntsPH7F9CTxz1Fp0JABw+/f2TeD8maWrBj
bwvcV1ZWsrKLPZN7oVxY4GlioC3mnAjARX3cICrGx0ApXW6rySd4Ke06KFv2GGtYkuaSDVgUxES5
OKCwJI7G+5Cuu0PZzgl7g6CW0RwXj8GmHE98c96V+AsGxdW/LR2IaO6Z49EJQ7mTWf0k8YN/V+yg
qcNo/7PotSbKWf9tRnFyo8YuQlscqlRGO7rieLoo+a6iuTJvhEchQ8vNS3/sfEdUVeoIGGV7mPbk
eiF0sdufwO7mJ+kAVLGptkiMkdA7wKqg15xhrY3ByUw6Be8O/dWqSKApSnmlmR77bBNMwnc0yh88
uB1S6tAhJoPFaha7/f3eGbKSDEq19VMuijg0hUB/jUJdFpxD7tmACgV89huUm39x570LVfTqA20n
+LrmpgNYjJ0rn0tKgPuRpPC6wjAkMRoZeU3Sh7jdUgOQI5X4gcbDJ2uvzWLpy7JdHFDaoa+tsRBM
gvtP7Zzr+XCBItI1iAxnkBZt4InJz+4KrHhloTH2FMma+T0grkFBEZTbA1oBTBB25mw2Rx8OAQjz
EzYy5jWfJXHtC5xGyNZqd3bwDHQ7mkQe5kYOVMnSHLKD1/cpjm0R0AauN/EHQucuzGqkeU4aZF8U
xaShMEwjP4Y1sG4Z1EXnbjBuQ58eS99Z2vdVNe4upxAMq8TTV+jv7g3CMgy1OMX1r9Cv80AMoGl7
b0buMVQqBXDfzAm0t3Pczg6E+TfUWsS6ZjM3Qj2kkXIPrwuHZBP2oS2Oyhy3z9o51xBvS3eUXhXF
DJQ6Ye5V1hkckTeIRsqaZ4ZqVJcdddRPLejJcKLzEMQGcJKogXnM+2OkIwlWr8JHZHiTz35r6x85
Y/QQO3UUF9sIO4P2vgDReWcxM4IGLTR0vse9ZDka7x97l6vh+IrTQUylbq+zBNbyPszuyaHTwuwc
hQq8jN/g+QISBS33eTald/3ih8in/1tpl0PB8zJW5zgJHtImbcGt3ygj+b362ktc+ogSw1IncE+I
mlFNFuVwCDAySYA8suJT2rTu7Op6jObrf76fCkdsECEYICc3pYOEqbTkrfqK+Pal/FH0ylZtcj47
PxCjecRWKEmt95x0pjYuGXc1xK+t9edcwe8E36/jekgqRKfsk2YCqBxUImAnuem0UPvJGiI7xNY+
dWzoq4b7zGTIp0ODN2C+ad4+brlKMIT3fgL3tj/tOQ2MNZuFlcizjvCe3Vs/YavGSwUv6Go5NrRI
EC6W0rpk7yvNLOy3i6ZeEvl9eKyJEgUJ3zsnbi1yOTnqvX86ArMbHYNMZxe351PP9PYdpwp0OaqN
00j8Hg0GxeKxay7//8f3Adl3Vwzhmo68tro+NEDYleLtHCT8qoex42djYp2jRNiTa2hPC4o2+CPL
KzF9IbiKAJpEG+0O4HE5uv4/m3GSeP8srDnL3fZcXk+t9MzciMuFt8SkO4qzJUpFLy4KmkGPsAR2
SH46wkE50jdxgUXnVcCx9qiPkk2rLUsh0L6NLtIba4av9E97TT+DNOL0ief5AEOZWs8elokCx2jf
1FrsXh8ucc2IJA5r3hhusAIq5tGKS1x8BlEpEYzNzVwz+Pr2m8a3Aw0KGdtz4fqRnYIg5CYaYzUA
fcpG1KaJyze2CoLjWsZkteFZRNwoF3lCZD0xVbkZZYUPpx2sVru2M7ASJr+MEA+ME8Vrmcyt2zMZ
bbHObeTyWTcAGskEmBS1pHpdlk1MItMfd6BUnhjr7pQiYFhT7eABnlrFLahIkEawHBQRPeGnn7fQ
k7MrXRfIuEC3A8xkQ7M45gwOBN3iMdsH/bZqd8Xwc2+DYoURO5LZx1MqeSNPA8wLTIl/l4s13b4Q
LHZAVPrQbKSHil0cqgIpXmPEfGOR8VxF2dtCvisAvNTF7pzHwIImA4Jb8h+tQBGySqRmqqqK+bYg
afd9AeHYHygDNlyL1HaLoAn4u6PFKU82WElOYnMwTJ47Y9ahpl6vZFF4UMTdvO1Ddt/liipu2KIi
nNbQfiMdhqRzif1ioLu38TT5mgMAwRUy8toBBZgSf8Fj0gNYvJQo75HDlsdTkbK+5zCnEMizlmbh
ribjOPfSJK9119aFvPbXU8+N4qD9YYM8jNQH+UGL/frBreqWTu/P9HiJd261o1UBkVLU0yHlbH4A
hW4yDaxKrgpcDX6Vj8thn4qu9pPzI6A+uk7NY5pglCQw1rO5MKb3JNUv1aZ95uBGz6GcRvxrXweD
BtuL86pPW3nzJT0lJbaYL2fWATc2RaIoHDsqy3H4SAkndyXsPtVw35gy+l75jlLEmSdmutgeJlpf
u05Obv424EJTgfu0Czbxr0TDg92YfYKelC1rDtY5+XI2T401lYnwWy/TF5WeomIqpadO9XK3TwHr
Y79X2/B+4B7XlZ++NnXOcKiOZQt3ooNMIeD9WsYmnYQrDsrvNJXePdZK1JR7sfHEyWx1IDwNrD8u
XYzqpAi6CUDZrHWgAHqNpsgmltTthZ9kbVW2s4AA5fkWPjx6b3XUTkzJh9q7eqsRhfucuxBo5bbO
qhGBeK02kMBaF5PGeJvwBNKF1KGd5+v9N1tWWe9+A01YCVecpdkr9cDtaVEoA0d2OQH3lj7szHFW
LSQ9HIUVanfXlD6mxlQxiKxixgNrX0qNuyHTj/eJcdFy8QTFxKBWKZSwXCND0vqRK62nicmTEZv1
LahzWRFtg+Mdczo5JQxTRTW1SMbD40H9+4Yu7GFIABhPEW5bJmVXDsnrWdfWDiHGdAsPgxrJpM6T
cXl+CJSkhE6D0svfgK++6ceitkQY/QIkckS2yunRqhsR8QUx8KBkBIa9s6KG79+BdVxvOglnDx83
vrRfAorkcdyg4Uv6mGspc9omB+nYyVNcV/kBjdD8wvdSIIkrQN6/I2A4lYgLDUxP+xqDOAUdJNGd
CRb3VwsAD5GjXDCaVM2Ejc2qI7Pxav2Mc27gKsEoYOi0A7dckIRjlwoUWzBsYnWY0WvLVhZ/GNkP
DczqNiY8PnOtCFSFplQePuAjjMXPBEqxvotSSdGM+ZKFJ4bHIjMgAVN0635lsGylIF7jHZzam7DW
7If0l7nZ1knmpTVOjw7QQBnZcdqESvI40X2ZHaeESudg2H89Y9GzPoldlOU6VuAFaqbPBAjLxFBl
DhM0KzSlyXP7lEasU6rDUFzfL8HuiPchKnwnLOzZ/A7Kv1ni5Qeu2aR1jE0wUbEkrz5tgVmROpTr
BkvOG9JVAtT5+kzPlb++sVktvDi8EpIE5Yd3DpcTdZkszBVhHWkSWHlJ6llLftaQ3n8VKkUFiztl
8EeZDAnMyPTod76ZlrOrf46rIGUxXpS90Dyt/mI1ihvfLIWjAO+52zWRsEmVhyrsN9c947F9zSSv
I4UVt7ZdSdJI5lWzsvnwH7Yoadg20skFo7c001nqLEbrFMCKhCK2JjYJNV/+C8sJK+27LmrCVBZg
xx8qngq6aR+FcaMQIfqXJ9vHfWnQQawY1+RxvYlSNJrhnr8THOAALkEIFBg4n/nzxsHfFWR/w60i
6NBPKss2zaKBLoEC5ztYBqbncALmbut3jTHTSFiOB7nuTP61bSyGRV7s7W4h+uFjddJaZtxJRMoV
nrdzu0iJ5ASoBL/TyodVQb//kprb1ikaxiZ//2mBO3sZYGNNfczTJR1++VN6kaojxR/U0hL92gyr
2RA5RxEghJOCJL2NyCZKXZ3UIb65qgilKGGiVLmlgIvT4mkl6U8Mijt0sw7rD8Qa5juaNFpIk8nX
eZQqNlacxPuA13UXSfYIF07S6Gih+8jmpQuRUsUkAaVAF0ZKBEw6bETDUcNpr+nPo+e3RgxGrz2M
2hMPcanQj6r2MHYP52eAw58qfT+8R7Nbbj8WIbg3rE0F0pSJ+3r2sHQTcIT78d6WlPNsdi1h/mM4
eFs4tPBH6NPG3L8PjUSRVc3Cl/3uD7ruEhS/ksETP4XuJ7/W5UEOF4k4IXUNyX5u2hPCKt0bItGE
3oKil681LyPAHyyCUrNytuHrLJkG2xnS949snYmKKJ7LQdcSoPSJ5I/1sMHVRoBHyDbL82t70phm
YRJj2ocO7iZNc5TNgMkA7Kr9MtDBknZSV5+vWu4iTUQJ+F9d1ZVPSkKu3Z+Vf+H69f/sVziFaA5+
b4zTy955m6/Qyo7pouqM3T4zQDWv4/0tabeHdS4OyrkO1fNDkBJuEelP/Kbz+o7J5EwTf8Sl9PBK
8yZ8A9ObWScI3o6Fy3B2rXrpN9+Mw7YBBueYdrVl/uiotBfZl3pNw0fAYnOQ9YA3x9k7IEeQ5m79
RP0JZtQQnLJ0UDuu2XZyOGzaKJkxiPP2BDHoJS4rHRdWzAwVeQR/GsMjEjkxKpKvHgv6SG9APDfj
Yi4BrQc/M5NSDxm+etIB+tZHK0lpfbeKqR1qs2urncjyHXGOk9cyMYZkzS/wKJkpOPolQymoPpA1
5tHZvfIULzKcWw68DacpUcZmmK+YKKCxPjCHjc5rUzwSVLjNLIv2mgED8CZjf/029PjtpNK3fYFc
dwCdy+2jXCugjfzIFe+EpW27rYzL4sAC1CpFjPf82wU01fRIuu+RgF8N+IGOTB3Ne94iH2tuAJYK
kp1X/wkrNV9khfERWu4GebRN4c0B4dbdEDM/Tvk76rTf/T2I/1RhkmO1qzWU8C7c3UE87wQBJ3rG
V3T5e+nrDbfzr5GuzzxwGkYbLKxT38GQ0sIGj7qDEqSzFRtl7K5fMesUNdgCFwhcZnPSPetENa77
FeVoCC5DpsHZUmeHKFK6UjadQ9KOVrDFCBGAzumZDxpylsO/SftebBpGOBEQmH/e4JZWXBWjnHeC
GecFsM9jVD2erK8NnxmelXEZAKousf9IBXIHXtYHp5tyRsRc0rBbOJHpCqYp87wI7Q8zBNXARZtB
vKpaxipmSjm7HyXvFjwUySgUHMPZfYshcueAqzOyOtCxLv+EhqQGshRtdJ0OwPTlZc4Edxrf+QGo
6u5QJyxzBpxQvm9FIzBFMT4VMjWIk9ByZdawcVNw2bOddjXb4ErpwD6p+Pv7IIhYDZf8WAdC9hx0
EWB/63HsFBmOoCzbtJiYPU7hJbssNm3oocuZjhYUlQGwbFgOL6vxqbG9OY02Otz3MBu2hLkRQilv
76LDbBi9FQOn74f6JoZvNPRxF6+IwPTv75Hj2opVMPRhb3BxS2GjRBcFpo1YQvzxly6t58cjPRxl
ZZ+SESlZrlIKoqhN5iOJCgyT+n9vsfyw1TkNL3QyY4zAimrFA6leAVa7GX4myyiMCDNEG26a1J12
Bcq2m9r8d0ZZHEbAmarR+PJANR0mcOyAUaC3zT+Sz/oS3v2U49TM2Y5QyKVpN0xiuhBIhkUrgDQ+
786Bw4Z84cqyjfGr4waCIPO1q1bqR1wMQ8XTvbQyvtYj4yYECTuL8xbl2kCkAbLnQp3uNOdgHVoX
Ex51HAjAw2LQr1xRZ+B5mOAE/cEXZl+srPVlZjAiTIt2bo5O8+fVsJ4JULosNIjKXcTcDjJFsThS
XVk1tl257AzM3bQ7Uo+SZoPJnp5rnZF1t1X6StQbAqnSJ9Xmcuia34165FQ6FfNCO/BMj26QjadO
opquQnMED/GYKxthVrhZb2ZPSNM7alftkFfD5PHYI4F9dEHZDqr6G5uyk3S4vN4xLBCVw448N+8s
pbMqwB0LSmHFic4j0EpjO+GogjGJiwwAHqVFNdBFrm9YyaScipJlflbkH3tuoTrDG/HEW3qiUqqi
Zk3n+CPCswVHaWJEKViu+PAvEJoEEzs5s9+QvM9jVbj+XMRmosvyGRQkBb5MFjE2oCbf2+Zpv6sN
FuXMGenEdzUd+RyNxprj6Dhlo668xJPeIhGj2v5GjmgU29j3LKyBCqPXtnLzUcdITBQyE8cPuHhG
FlwMO+11/HestqVNugu/MhUhaRupOu56JEeeBk9VIhyILKLm3AS5OWXMdqMgazv+FaC/TjCpViDo
fAg/kANTELReicaCwEciaXKlCN+EilGU+LyHSyh/goS8zmJWzMpGA+Uig5zWmBbmY5pU3nE+BwrP
apEEtleVINRfbEtnQ3OWA+kHygKh+LJRNuEXDiQz5o/VYVXYwqRfdCD/x68JDvXsAHVULcH4wHx+
HXC3Gcuoc/GMI8je6uFxGiMN/t9JtIkpB0gQ8smfnVO+fVsY5+uG74qXqtu06esMRMazbQXJ1FsN
J5FZ/EsyPFafnb1cTpwX2Cv0tFxuQWHddDheFk34rsWDn0+AVfrEQ0N8G+WyEfugYfe1aJKjGjdk
CdffOxQ5eTnX4MFyOr0U5H90YIfX5uXS9pWo4hAvV1VhvpHqYOykbkC+C20Mg4P7Uy53RBqZy3Jf
mH8PWv+tnL/W5nZnoomrk2d4jpogVzhG0TF8xQjb31gH/O6l1K1rh5OMKwvAyvFvjanyW3PU1qHA
mbh7bgehblUJcdEux5gMtWqL4cApF5Vb8XjHD/ruFW5fSf798Wx6VNVWYWGUTRMuZdjPucxLqlF8
RJ+6HCXIq8rDyAkIYDOWlwrcIP03O4I/kGOYi+rBtm+go59vEBBG30h0RrHpra3KBIOAP+TriqKP
vxRFYRWsIXsadjnUw0MYMVvOQId8cZO/3o9t+5Y1fupDsh28/1+BhQeJYp69zMlyrDTYUaU5OGLH
c+fuMrR0mJ5vDHIWnCe/WqsGAAzNOWHGqVFzVT+VgeI9QPimQeahZ1f0RQF4+GUCtzGxkzMp2UAf
QZtbRP9kzYjQvNvs0lG1rFfgXVw4M25tmjCy3AOi5a79KyfVQjB/odoLCpk3C4ZlCtiKcvd/bHdg
jA4k94+sw1ufDZraR4G3ksA45NKD7dnU58/3OzG6VAX01OBc23NJuV1HaoMoHbuTueDkkAXa6xbP
vbzDUGoRvH4z0EA4sxQvDA9n9+Qy8JwCU5s8pFLVFjRDARQhRApv0Uhw6hohqeYKaFA0aFVSzHOj
FKo5opa1WvYFyXpi4kMeX2ZfXr5XZ7tNmuXpj7q5LoqIAZAsNtrXiPCfRBV2E10gtMdgD2IotevI
z2mzednY8AVhqz1bRK8UKrb47nab2t0dDnmpwNEYwxvz1QKz+Fe6E5Zur7dE1eOn7h3Otwr9A3cp
xCbIOJCL7E9RPaeo9flf+AHKcAbV2pUc6FK46VoEUgbu6N2tejdrledDm7ib1ihr9QWyAlN6ygdx
e3Te99I7HIHIeDuV4RVpyHXye5GsVM7tZitEKKZ2to+ZCjbhfcYuXEdhVk53bD2rrSRT+tSWlOHj
g87QZ9uwxHW0BSBiM6+Y5sm1/MYPi0QDT96mtjjVpOtEiJwyi9LHyiA0yPPvt3lMW0MeQTodNXJ4
yvZ40Dz1zetVZBMZsU0VR5ufGEMx2hfW+oxFV3htofz3iGnhkxCn6sfcfA0OE9Y1PhGsHNto40mm
cK7uHHV7fmXmzdx/zI3M7f/UUDHEgHgF5Tjjv0G8Sz5ADttb3SgDtrMONP+AXLnmYHQuLNp/beUv
DRDg2V0PGaystN//YVRg1tqYwrSmjyj7U0R/1IZLXsQ3X/kSv6WlwyJQgB3OHFsg1HupnjIMwc2d
24kjNDmMi9rDO55hQDd9qN9oVbkQYSsdzdzpnEbUfhBbzFjMoPmiG8LNBS/5L6E/w5P+y3MNX9d0
ZFF/9Mb0YP7bca6gXhjGRY47PGH+S/b5pixBEEavMooN1K/c9BxN2bf6dkUGxu8TMbTGxhXz0t8J
gJp96Oa/xLfLzqQeRHn2J9p4IPkIMl+XUklRyNIn984la78a5VveYXef+TkSIKrecAGy5eHJJGp5
jhLm6/jfj1CslaOM7a0OIe150t74EUo15+FAmQhdmUlv1JiMB7YOhl4C44JL+o44/pAc8YHupSWH
TWSgTx7ETe9eSPRcs7kYUHmaLk9cMs91lSC3tkmkbdtdER44LIvNPlFlNUM+SwdNFewQ7o3xeU7s
0w7KiM5BhjGcn2TYBzMpgqiwnQvulpDDoKw1JHwuFr7eobm2iv26p6G+M/0AlFRxznv44a7JjKuw
Jzq6vd6RtwTzG6vB861wIDkdDHb8LssFWPVPhcKKB9gdnqCMVeLSIdkPZjXn+HECuwfx5uqGOZ0U
w1NiPrMbSQto7M2d9RrTJMmgCc9tjxGqZLgAhFOZB1rbGI5p0ySXutjliiw8YnRdHpFVa2PP5S5g
54fHRVDd/NaQEya2D/uui7SwZxGtt0yY6OlIcYY6Leg0sMliTkT8GM62trLs0w2gwkgc7wN8A0s7
lg19tLphas2l18iM1WScZf/Xt46V7KvVkDWgmtoDf5Eagmy9X5TwqjoJ1hWiBYwkvWUUmMGlvmLH
x8Iy40s65Izs/emVwtzl7zECbcZt/Az1NHS5fCDbXDg6MqwKwj5D5aURc+kj1+yqjwqUbFjB8h84
b2eo++F0RMXjb84TDS+W6Rq1a98NeMBTZV9yT9Tp/DX1DXcSUS+N42BPi5jjFwbVkH9FopC0/6K2
d2LEFOeAm/iCcXZx2/LoaCqmYxr0p/9kYxIqiLlrOdFmKLWJxuCWOPVlh1PQjLpurdELj/pSbA+f
c/GmWgb3h+dhQIFzZ+CcSG7oro4ENYd6OcsykHmHC+malhBqjo3ZiiTb/6Gt1AFkNMU+vvegCLmu
41jRwrU4lUQXKVA3BqKWo9RSpMxbCCdK6woF1HoSq/QGNrGXzjKi0dBU4vPlxhOg+XTox9RiSGYy
wHOXKtdNNYp3drR32/Il5MrlwNTsm1I6gKdWJQbxhafX638GfcH4bX1nJiaDVUme62BpG3pRSt5H
EUp7o7QpXErqHEkqptK3HBCUZc9ZTFjgjYRyCzLr2vJrhNsxw0xkflArZHxpJQYqKEFv7HSBnFei
PFhIutcqtMnTsGzt34RKBVJUosil5lyX8CTuibbgp39TdLtaHi2X05EBuvQCYs00xlruh9vwznNO
VcxCs091vkNqarGU/0ipBhi06vOvTj3UFxQxJSdvNuaZvk+CkZzVcWcMK8XlKNuImgLLRxUTyrSz
Us3dDgmH1Drt89lO6KnJJXRvxfW0xsH2Z0POjPBLzyDW5voRYWAyelhha+zPiSeNiDKuww2+HsZQ
doYFdVrqZoqT6fKA5n9ZIWF8RlbNByJJFTrgNW1kZiqarGcvrkSzKuGZbHB5W0njMnlMcKiceb4i
7D/qqvcX0rMj2PB0/fzXHpx3TOAGteOzlc2pquTLI/pbhr6sF9KmqgKy1kYjZWwyAMmXFdJPOrdn
4L19aSE3s4pgOWzWZJVRAhEuW1Gop0S4SKBYIgcPT9dWWNkxCHNuzQVdvRQAGb2fpgeXH/RU/GIP
uGbkns7iQNLQzDqaBVT07mNzEWdFisxlO6tsXPaqhMCbYVyUw4TqCADSRKE4JjbjOAfzOobnt6Y+
V5+zCifJCL/lHUoNkF86IHzdYM2Ikqpi+IT77kLQrOf3aXxIEEulOFrucgv/bmDlXIwFezexenCS
dmWFP1nqAcZVKgAFmSqkADjtt307ludpn9DGG/nQKXzQgHYBe2frBusJHJBr1RsJZYTH49GzOu8E
7dDq4TsxvT07R14X/m0PuCmZ45P2CvFQe/TOywtqzHXZ9x1heI6vZMzp+XshX+/aLVm/oe0CaFEp
UkBo5SYXXBdRl/NuNLNgZOaKimqv9JgoGnaPU5q1rqUow1XVIZ8FynwREFgVuFc4hQQXM74iIlfR
8Hxq/ZGYs93UVDEc/BYk8iB9ZLqpVQUokQdUgz4aZjjY8N0pd8vLmH7fCHqNpxcTuPNVaeNJOV2J
nxYlzcZOYDNYBkBHlAQ1lf7Lh3jUeizHnm+PcGEMyfcsb1qhCC3XFqXXpZrBGkSBApTRppv2Bpx0
pS6opIkvQI7cpPUSarisjDDX2D19zjXvxPfyTkwiMRXX/SKoUDAevCEpN9tOLsTxcq3xBpnyXL7l
TW3KAjk/neDtSc0ecXBBCM2L/HsS/glkeYmB5DjjkxPzfvvn4cDB+/aQJN4cngEGJ0ILNW2zF5sp
NVe7omGSlOHK4eGc1gxtuFFcRWrUOdd7XcmjzKAMiCltIm03xVwEUoKN7DogPXeB285Qr57pXnwn
G/chBFDq1IDwg0GfpFdp3iCFONt9qcnwJaN/vGfKozBQ6f4OXywOifCjuR+IE+mw0nC74oJHO6Sh
/+MKyExpC+zWhCSRdHDrOxTr61/qt9mVAVZuwTdDK5vAMXwv08o/eVmAGUr2yxNJkODc3Vcl94vm
wYN1YGeW2zKmc1225fXYVSvXcIhs7gNgvdc6ydLlJjkkJ2kjTjdARKWqzrBDJkl4mUuVWUqC6cI/
XGDRWC7Fs4g7c/zsSARrea16mZEZ04H47UtBHf4m3Ov3XIVpg27zNR792AZh1E0g+F7xpBdP+shR
d6xDbi7HbzoFURWDZXwxP0keSQ4SnNOns5IaHuH2NA+z/NzNX1NFTwW35ZF3CAp2BZjfcaCp+yPd
ZNxVuuYeB/duz33QUlu4+VYB7+Ez4phK7kMlA2LhntbGz+yTYkd8pvw0HaECoUtcyBRM/npTdtlV
v2s0u++NpYxJijUH/V06wAWTpRdBxZUzhzYwOQGWdfrrxdxPOn0m/pcKzGYQLlnu3cULTm7QaF3T
DC6wJGWtyM/pHSqG/Soi4GbIxHVeAI+qEVVceWcxnSWdyekdrDTg4hUdM8uZ2Kv9WaGq7hS1X3yI
Lnqj5XMqxVCGNGyUWQD8LlCis7AQW11Ej5eZ6ijItXkbVj1Naxgxd6LNJ5AzvzNKwa6a22SW/etH
3ORwLOCSDkI4//JG28SxRk+coY7V6nfp/NKg94CGR/evZf+IPHssxnlvjaqH4x0Kv2hAhwBorW8A
VEwCBXzBC3id5E+tSUmtgMLEFlOKGhT/4x7Auc2fMC3fPnu30wHpZGrwHHKieGOCoCJK/tWGsnk7
mzlDHYRRyJHNlk9Lza4LXIqErGy++Hi6OqTnEEA31eLWPYaFhzx+F7F20pGWKswO7Tr6EHZQTmqy
m66bQmlN0IOxBwPlbJA6jU+jHNbNoXYYZRbkk7LfH+8b1UUooeRgmKqRq5CymNzyHn8Za/ykU/EH
JlYdO026VUfgNQwXSMUFWcG/cXZ3znYiEUh8L/LxirQhuxgF6b1SlTEA9b9XXN/y0EMckmY22HYq
QUwKknv99xvK/uZnFJwxB7V3WNRJUc6wXTke9GXZ9Czvr9+aVnvQDmmIyw9DFegOx0kZQSmQEdkI
Sz7tWJQc2Yl8lSoJsqVJ0FlmVk6W6jiKBD3C7sRoZEcZBsX2sz6NYtSnop2Di4VnZ7UZi6y83phd
VhSKat9r7qyGaTLfeSPRk7r7sSuw8NaSPpN44/mFVIXyuhfVwThrG4UuJjzWhI2NXTImUqNiqUh9
4xQYo05M7lWWfX/B0HrZLV15Mwe9OSNW35UNE6ddGFr2h0Y/FG8KucL2JgRfxgHXptgSCY4VSu0R
C+qx8Y3EAb83znVLRv0hB5SJMnhDlaRVISVRhv4LrNyKYTp2xY29g1FconJczaIxALuOsnr/RllY
+TYjpFKhnikgG0nVQ83KpP1IJf0w6Xq2de6kH8gVLaA15EA/3yzgVyvPYT7FuHvjGVKxAcrGPoIA
tsygLNvWYyUNz1xEX0XjOFCvzslN/kW/Pa+X/QnFB1gg644vBItsroF58Gq/mFo1sv2Df9T2f/5R
BzlnJR0g3oKQnb6UktBRzqVFCjPQdaTVuz02JB5o3GhArXCgV+Q7Y6tcfTgchP6Pm2mXKGWuebt6
emCeSP/9OhmyGESUKWdxUiVUz5XtTEvGB72PRF0jUWNEKrRX0mWe6sQPoLgojF8LHZpgGiCHpFV3
RK1HPaKll8beM5VWEGbRHR+J7fbVKT0zWmNjZbvT4QWq6XgvymGt0ONsDQHk9UBbX2RHhD2Ak+FO
YPCVBKN2RxR0riUg4pOWWqVtwKVza9GvsVt7CMGzVHwoQCHVZfmo0Rc5sZlfK13vp57hur7M78SR
bbW68MzPlKQ2kUJJYKcVLlnivYvKH8eMuud5QbILeCZcwZFwMURHDCrRZi6J3VWNPIUJtU6vuVbC
2tvSbGofLErnplhRQKYPWqiQHbjpfEe48PjGFosL+mkQRRWtG2j2zVISbjpH7Sk7kUBMxbj1Mfqb
CIPdoKLRYzUWoieS5eOSMk3imln5ahGLcofRMORnuOkmqZKtvHtuYlsnn90JrnstHAoqPgMKUN4A
OU1e4gDz/kQgx0Mh1KcC/wuE6wfX0R+88++dZjUmwUa8ucdCToOj/NDRjQ/KgrieFmv9XU2ubuze
+G3t2BBq4Uheh8et5CreINV7wV9JAaOJPBmg2D0KDjVwDTH9oaWPMTAGo8bXDICukf+juAT27Dr5
Bnvm+IA0ued3xvqQoX/4K3jGNXZeqh2z5VlyP5qbxKixHGdefg3k7eTipext1Aqc/Yeci3zTIMB2
WVZahHRWNekKw7hHLVOGljmIRaRanthcAOnY07TyOX3v5mZI3Ch1eb2+7f8fIz7DT5g8+s86f+yR
zC5zIcQN+mtYpTsCJDEcmyBRZ4HqAcufTzhFwleLC6nPZUGeJr9vLFqlLvEq4AQsAGcSPfAVHDVY
NZZXXx4u0YReuElqmFaAYjM6YuNzKnf2nbz2P7f7IhLcbvX2YNoVJfPfXE09xIgMF5CDAiL27plh
ZaxJrSqmBD1Y9oP6+2gtOddnwtNKtj7IgY9EWNu8KnOsJAc4L0gxDEXsMyyjaazOyqJAHOsJnFXy
rejb33UVr3TiWjh8EiUDfP9f4byWjtTINwdG0PYl0hEWdKK1g4+3B6Rc8SWEAM25998UefJLMnT6
97zVhw6Ypip/HRVMFBMD/MO6Y/B5gFXNIdZluA865OscUs9jQ1QCO8j8EDUc5OPfOgzttT1OlkN3
rtk9hKOp+uoWebIMp3Ut4SsRHAmSUYUM/9ZF2JCP+lsrZtZ7xo4a99SUJjUrgzMvJI5MXiF8Twjg
wBx+WrHOdh64TWIwsaxSbrTUYxPmP8Dp5Ss14RiZlCn6Oax3atL0Dxo19YU/8KbGN9YH3fGyQFSG
YH6kDlwMUmMFGKbBr/8u9Fj9D2nMIV/aRUoAN3RvjP76UbzMkyMC6JBScQppUr0y0rhUoEk7/vlk
YsHA5S+lAfKgR/MLk+SwxW4qQmOJ999EqzhECR8vDVaeuozjllZaD/szMBP+wQtdYUNNY/0AQ7Z5
wBrZTjUYq+EOdKX0zr3mKS7ceqdGdXl5/4KzjsZsVXjV4+jv/dbVYw+pB3YOx3nzunEEs4N2RvW7
fYEl0i6CiiTAokO1l8IpydlZmWr+pJI4lLQAEgxomWNN0JoYHRgvr3qoi6R6P4Go3atA414Shont
tP1Txak7W91nZwHd5fDpqrMlsqpAbkHh2o7Ffaw/2YjAnw+UPyjkMJnM9jNzbkCr/tfw6EdmejTZ
+2ZQStyGI72arq7Iuji6bpZOMGwZtMmv4YjqRtR5Y4/g1lPq/ZICeDecCR93fDPVL8Ztm2v5ThYz
YwAggb5cj9RToKrdU9xcS32dKQju0bKco08jxofe/qvGpqN93CJPTjotoJbOgOBQJb46gdQoo21c
Bq5iRcSJEeIdSGD9OYt59lYE8xDOW/RmkYaXdoLyZQQ9ua+JFLpzv0EFavGizTcfQnRe2C87b4LP
FKv5rlw979QbhLdMYqXlA7RKmM9wxlRpWFhHQhoah5fGejZmSnqK5unPPMWJbWIUCZAOAcN279jM
uYU7ST3fA683UdwseqgE9N0/4XXg/B6OuQX+1fJ34AC+GLiG0ieLaQJgc4FySeqGkS+mgeQGbqbv
q9Ti0hO4KzuiTnN+eK5ReGAXOETsA3JbmGfXqUHlMhCpzxl/dUa/h0mIUF1aAllGq01mIlHi+guC
d0JOruAumnqEhwZAbCChkX30DIFE0vm5UqRFsZRaQG+rz+w1400dtpfQxM1fBG9TT5INOh4uqFML
FL1HgLcpQYecmshhfredMjbLY/wpzWXBWAetcMwS17Qeawf+ao7jL4JymB+K57/rCCt7qQ1d0PdJ
xuEhCvS3fFHLPal7VA+mLRsVUKpCeyb0MOd+luG/e9sqWsMBcTVeAGClK2wSm4BcjW6ix05aV3uu
PKfY9rbvoSdl1EM78siFc12/AoQ+YoWQwdGeCNPyhVc35UHsH1FxDJjPEhecLOmElIUDuveCQqoB
s/b6LwYkgPtyYww+zNgPfJL9f8I29i3hkye1ug2G7OC3VdSTir/A4IpH1GwjGvNwPMlxlyDSYG+D
Zi1LtS4e/Y/uM1L1YA3UOjDj2zcsj+PfNSvxZRzk2u6eY4YIzlWdrwNm70H5RkOJyr0v1HJy6x1z
4AJPMbk3Q+hC3fbGVNSXm9phHT1jjoWEpaHyoswgbZ1nUsT4hgfIGKN7mzqKHMeJfEoQtFQgP66I
+5KWDi/psijulrHvHbg6JEaYG8FmoIrpCsXDlbqv5prT5XSCTOWQ8oYmUJUS/qApD5B2PGQcRqb/
thdm64Ud4uWClLVbIjB817kSFlsYfC+u3Idy4nfFLb5uUg0yn0y5lyQ0nabNCHUmnfk0cIMpeXhU
6+AVmoGRLENXuHaQrprHiLb751TtxsrLow0Ich8VqrZPakBo2/V5/UYAE8JODYlMlLqTd5vIHGXB
iSQ+AA0cu/5joJ0BRyDjc88tnrI1f58TGyorOUsLCbF3liqm5aK7ZEMUc+14dZSnzaQ4ZKrSCrIQ
l/Y9d3fEbbZBuLK8AZU1i5PRYp6DgqlDaAQygYQkn5wBfmZ5bbHaw7dqc8I5rU3pR5FxzCILyL34
hfbJS5EGzYvv9B2bWkm66wO5hUZfN2uhsEE1ap0diZbP3/gVNmz9aP61smKAg+lAVIilKOAFBrmg
XoaRT9SZC6ZRdO4QVsAFfYmpHZJG4ankyF+2sJc9PDV7hGV3/3oEgH2sreZ0w711sdT61fwWtJxP
jNCxFwonQperOJGrNDzQ7iTQGn4AAoZCLnaslrcXLSyt/w9EW41z56e1hvcDUvF/pai/fdg9hYts
17siAcgqBLDQOKfuRosM/K6d4AFuoP8mJMBlTwNxnj59HiS/fAdWSECKB+S8JoQouIrov4Qauka5
hxuVYgcM06w8FOebBGaiXMN3Z8h+kWGWoypGypwmwZCPrCRgp26dzPsPU/yU9zj9UhlZdLPegBPC
+qZhuD3cDI0iMrKMN7tjb6JdhbMh92Ky9P/TVZdyf1giLBhr9z0ntSrev/3BKP/u7PmyJpi91rx+
F7X78vkCkKnrsdZow45eeKKHyasL9C5T/JMs6r2GL2nCxygVzhzv0YvmfwgoUX02nmIBUROjvnce
Ooho/npAtO/psFtN1KG/9T1mPdegjiRGCwHNf11ev6FQ4TST8mraJB89+gDgvz+YZOQbwEPy4UFN
IzczZ/OPF2rODzfEJau2c/e0iMuXTmamTKb6B93DJyGa4BW8owWEutNp1o4BdMBjKPUfFaTRPoQ+
dMnTFXt7Ro+qWIJq5oT/cbIg+sKplu1gpzY4idtxzGprNk0BXQAro/6NZ8zCDmUSMQD4rRiea/lR
u5mzs2kZgTRrAbH55xIb7ZbpahZ7WPO78SmN3qlhki2sF7VnwCD6aTCL/ooQ2jYp6O14qxpHPwl+
+GkVAiktJnoX90+3WpUcGibiSm3CYKab3BpnjMEw5KSgireNhBdj6Sg36H0gy5gp/6zthKFV2X69
UVtPkW79qXiXuzMabK2DAL3gqAPEMDKGjIdpDNFbeI72ALBFZzgkZeCmYVgzuX3CMEf9zSdqXtEk
RfW++P9O1Z1rLNMVPYW16UjCeZ2QVLkFcb+nhkaaMrG8TMwi1J6RIL9Mau6PnWbUVvJNTMH9TdjG
ccjYfXznfv7K00AuHwL+9PpJC2xAq2T620ZgywJHQ0UWy5pZVJu3mmonZdTA1gOW8r5chV/+v7Y3
Rb9iBilaEW3drrWi6H3JKaAl1LT8fNd7byjA31wMb0vti4V1zn77wNv4263KktKyEp5jHauOLCFR
Mv8a8JO7I26WU8aLkMov91bJDqoB8nxYuWRN6pFVwkSDCenLOTuZVg0UF6ivAiUznimvVxbzkmkT
HR6FoHysahzakjb8EGOQdVSq1erzSX7o5uNxP+96h6AXgnFHOixy4DXaZYVd9kCz6lCevz3Yn5iP
8PeiKxDco4es5WXaPSPvjU31u7vGnF5Qq/Dn66EymlA+G3Y8TsgQw0vbTFa4qr6c9oaLO4OB6+dv
ziyW3Tdh0B+R+oChC1b9y4t+pGmHFJXg9VsaQDROmsJcSaZErZDgMGCdrzq1hqx5TvOE9Ex6u1vC
edy77CNqBjNJunPc5H4TlmKHT4W2eIZnxuIO6cXRKjUYCFCCdFnEdk7BwIdf9BLT2asTlfh38v/j
m49hJW6sZTSBJfAk7mfeoLsOeMtYL04l3q1uyOjJbkO+Srz0fQa69I9ZBKVNYi+z6lwBp4EU6kcE
gbI0NOi/MYd0D56Wwd90KWKuGCSOtRtrJYyctdbD9WPmvOLWDZCU7imuKXeNwm1Ajz+a3SP+a0HJ
LKz/RMd7CVJ4Wij6i1sBr6ObjvNJn5WX29vlbepmd0uikAex6JRwmdrfUdVaUSM1kPUwnkF2fYj2
n0J2Kdp4lTk+sm9pfyaxv5sQ1C7ePonKa2dJkQyOvBxcghg6hS6t4NxAoI9rVoJodKhBnOjKqUI5
nMhre/qU3dCXv5qhFcxau78M0va+U7QMVs7fJtRFIWhF05P78Q5+hxxLhU7thEOEnaKNPhxslHxB
xoi+XkeBec/rzFYla+kivneDac9E2E9k62rs9FCvqlB8QCpJ1wrIW4b/xwoSTf8HTnElAacQM59O
fJLuhJ+utUMo2/BFr7v1dngkuUZXIWL5E7L/K1nQWups/EiyVvxzZ2E+tI6/y4GLVOKC+mi8GbWY
bxAQ2yhn4nNBHZeHG8WoTt565Xmr0yLgOeg+r1HeNaFR3JTaKgB7vayM3GoK4+WLJf3D5THgNyLp
EfzlQT0JnsRFQO6Bc5W5amatDEr0oHfPhCD3P/YesBWhwYX6CMnnQhnfD9r7j4GaUvNupyzExnH3
7vM4afz8SmUWHlbxHYRySl3T/+oJsYpNpRUIeklWgAIBkYBuO8n6JncQhb0S96txVa5jIhSI5OdF
/BDgqJsOarYmnkA1+JIzw6ijrCNJIrzHjOQW/vkiqttaf5i4HdLchY57dNF8Ca8HWVF+1BQ2OPRz
kiZl7+BllwGD+0g39oO42DzBKR9nuUl0JzFxbu1uvkUKRTDeGoEt4z5Xnh4bSNBrLM7Ikmr2Vjau
IjCIjTQb+EkOkvFF2yYFimk4jd3UkETZVaL8ga25YcMw8DeO5i65JiOVta4WjqzlnmIYMaXvwpFO
Q4L5+GlqQWE6tg2hFfyMhuUMnBv72bBoF0rgB04B4T57nbNZNq7h7ylm6K0Ne73xJwsYTsj4rLG9
HQTPbh5ink+c7xrlRHFkAZA4X6KABvbg0kOJVmW0fIG6A7Mg8zERmJ4yqf9AC5/aRldqV2jTcm8N
+zet1//+caGghNw/P/ARLbGguIatXOLPpfS4kHKuTSgZUSKynD7xkpqgsak2fxiDhkRXn10wx+Er
I1j5EYQp2+cYcPYyvoPFsFVpJtziYzvb+cruL2l+JXYj2kY0N8LcovpMcvN0PqfU8sjq9dFCE4Su
VWUK1DiDzTXjdUq4lHKGC8I+zn+ve1rdbYIp55u6E/SWzsj6gboJzfjCxJsBPj1F+wVBrLxfwtwp
elIqGYGwUHfbwzgx8xfkN+1wgiQXJanuHOsH4kETVWzYRWWFGUXwspdHSB3+AQWOkWWVtiPpnpkP
LIIJFdu4BwSZjEAcwddcTj0KBw2fIp4tetk78ox1Pare85fOgI/RmklKaV23/3hk0USyNmfjBQvc
llFiAnxhj++dsJaw7OwLhKTh8IfpDCjZ5CvFlr5NUf7vn3Ja7WpRIXsJPCue6OBB1is45C+vT2Je
ktSSuyWHad8FbKTk0NA6nmxjRzEDP3Yzwb43/KqPftFQjaynwgHd2cTRlx9RUEBRahQ5trCzHY6g
xhyu/t1ArqOnl2fD9qriSlAI5oI137MM6rzP9N+LuM1fUMumK6/fOQhieJ45ORqEin+tn0SlpeiC
vI3pxUGAKcM+Hi6+0PhRwmIH0HPYxcnhJDFzmpXtauyea0u8CWB4v9hob83gugacSG0L1em681fX
ZrZiuqJOJle+t4+WnUqQaHfKHSIhp/jyzDAs2/miL7yvpj65i3e7s6Iq4fssm5ZBCGnjh5FKgp9x
2stGDI0gm5Cce9x29HXJhyFUuSX12TJR4ixTzk+d9pIbsKrQjJsN8fWiV6IqvgBhptUxTtuvCuS+
w+ZfOhDtgh0WV4XtEj4gaAWe7m7flngUDPfoBVbEBpFX2LvkjqkK+HMi+Upz1U6VLgwJWH5mTm82
2TBQ+4DdqgOOQ28HdTHBySaNu0zr8x4qaHTfGQHywTk8mL29V29QD7f/gm67tlQD0GlA6pUr2NeY
JJ2s4F4sQ8tmz/iMMwTYR90qUloZ8UtJqSZ+N11nz8LxVqJGhFV3hIruI5x1y/X8BWHOalOjcazo
58DyZtqwCwg6IlUAwiwmYxkhD3KhsOOFBHgUFQ2HhXSAdPDbXnNtUvd7X2FLReJqvPcusw4qD4iX
d9Q9k7vHXoEBUNrmBcvqExVhjSwq/dDpAxfybs63XtUqHBv3vOrw8dVkQKFK+MtVrUdaxmptWGp4
Nf6rOw/wRuzenNq1a4EHBCB25grx/KfXG71dsozb7oeSLs94YLlh7wBbqfVZVxrpujWLSLuKAmqH
rnEj0x8VSVFAujjrHZxij6bIh8eEaPwW6JG0ETkaiMe4m/knwOZV5pNUo8mp55yVwlPIl+hcIpwH
R6KqyIryDgmwaSSPyDzkl577g/5g7p4uDx7nQ50lHt1oIuWz58OQ8lflemwHjrDLLR7H9ZOr5/Ee
619EQ9wb9s5I/y8NfzRCOaXVd8UkXL0/jtd+p2vgSj9eV4YcdGyiav6bdNbnKwJzFEijis9EJHnl
mHW5yTO1BVIklBF05JMHV1XqMvfsXN89KdoSZ78A87TmSwaHOyPkZGYw86bN0nPdIAuP1D+HAzSk
DU5zGkJGIRq1kPqEIJavwAfad6Wy70S34h7pPDqqbM1AbShUB6ES8saIgZZksdFruDDarukbjjb/
KWNu9nJKMWCinpBzZ6WZvOgslnKH2Cy1+fcc3l4u3yCQDyw5Wh0X2QWxMRsgq+GnhaKTOaxd2Yx5
x29TV0iLFhNGRbHDDBOTnT4+n7iTpohjclrMEuLxOAVv6SfNoWOnHGJ+9NJmOwJIkn6dl0HFQ60s
vQhtOA2XraqRGlwx+l8yFUjNiIvnnkTTwbe1HQ2Y9QtFgQrDkNUki4KAQCM+PdeJtrSIDD1foX77
AXXzO+AR1GAsia07OgsoxZCqjT4ECxl06MiyiWqypJVhBfduElN88GtmjQbi+iCajVXjhe73Gk3P
htNObP7dRiZ6VjQfZX08wt+4JSRvVV9b6hf+IAaOZq/PLiMvOPX8HQ6g7inhPk6PIQkFIp53UPRx
JesLGAt0Pyv70w8y9EX/gfsJrVKukC89d1oP3nJ/A7vM6ZFqc11yzw9OheHV9i52bvClFNibEhU4
OIBHNRpS6XNdp5MVMswESQFuqj+doz+nH1khMOUx7y9WgUG62AFrJEe7OQPj2dYzxp5rNypzU/BH
VkbWzI+9I9cgoZTghjFQftadZBQ79KYBV2O78ZIojUOrPWG3RBhp2d9GRMQnPioyex6leFlz4f5o
hjWxyn9+UeHm7LaCOxAmme8TqOOFEkXKIRpTEo5TfMqyp3hTCuukN2lejwK5WH9u8IHdHqA6u64n
VfU7+Zr5soXMloUEqupPYocPoDygc9gZ4zlkOT1EA6MQto80aZiRKHLIqEK2jg8kAUrO0w5AaonT
r80p0Pcop+RQmlklCSN0PjDSuY4LxOgzZPcfNsmLfvSf3Wil3P4poRMYFX/cndUycmlyI68lCHQ9
NkGvXAHb1pmBz/WmoyLovozPrTVNx1zGbPM1ViNQLpLxe2Pg4Ulu/G9j8T/frnHILPLahfJxhbCC
37XnNQLi6P39+tKU+/PAIcAJKxBkUPRWC3lGCilWAbue3rAMOaY0Yui+TH9u7COZ2gVz9XlHuob8
JSH0sg06Jsxnl2K5XnmFMqFhjUZBup0gdxWwjAP4PoBw3tpkHCscQQiOlgZJSkiXJbJAqnMWQImq
OSQKFNO1X4IDUFnq8iGtHXFfF7FJReOY70sVkcBdJ6EigEenzGmuE6MgZNHV2cBwijnfxD1tBlbk
Yux5ihptVhyP91scGIEIyNstSSWQtw94WnU96fXGoAtbqKQkGXbq4y+y4yWJfskuDrePIJ1f7Qk+
UVSQxB3xZkeqkt3X++DRZdkI+NQJflZFfl2X7Mv8NqDRPTxs0KdsRlhV3wM/0kr2a3BZ1TJGWPfF
9FF+D1rMFG9sDqBWFTwTPF9TfqiWdDitywSRZqzWT9j0lUzePivFFJrMTmVWDoQpeZp40NgKcvHB
U8qyqI5OCcy6s/3KLJmgKOsnSSa2Y1x1Zo7p1Gt4aiIAbKnwXH1OuXjIKbvH+tSm6HYj5694wFtL
aV+5+wb1jI7FGvZsy0Z9gTsY6XXQpyv+BDKPaM1unS6QS0/AF06w0KSLWqXxoStreSK4LnHENYMU
pKd7J41O66kCQUfKoieB0c/UHfMuMedoi7tR2i/Qabz+b0uDuGqxDps67TDBQQQQgzrNC1mHO/Zx
RqNWVMN2wUH+K06i6x6L8pzRbIUqvjxu9gwmP74niSvOrMtyFHxTVBb4dM0vfs/Mhn/ktH6ThlrU
fP9nH49ES0K3EPTTpIVRHR16sWwBS3s548TREEl/H42H+vEZePaDOLBv+iE4+HgKV7vVumZiL7mY
uC1NdljMbTnNbHcVQ+RCo0+/mUfDWjUKerq/BqMRqNqaxjTuAOeQT/TdCLyYaT+aLPGmO77X2JYf
73mxtOy0gCbMaowO9+hiaUtU6+t8xOedgP8bff4yzO9zSL71AkQOtcX8nkipjAd2tUqZ/hB6+uua
wYs/H73X6KCTGHn1io+tQkAKJvUe5Fi24w/6WEthkEsG53UmwbQ5vmH66Zdd8KIhzw6PllrfILAF
/ZFZ32BNbPlJGR0aCEgOUTMDy8minPZPvL5lkhZtNr0klYxop9gu+6i2ke9BdWvDTSIHMBurrvJZ
JxT5UUwUCjfYMg7EC2cfWEgmPDI53oS2r8/DU1QqtmQhCFnoJwToV9wK8mVy0C7Ulc2qC0C1zwxt
DI0FA9R49COYugvBPiDKdchUNyzvThEzvIF5TEfQvhqNIS0W7/87G1WdfMI7ImTjYiIQGrmW6XZK
GeOmTwSKppwXgYj2aj/C269HSqtxA49E0WNNCC8zy4WPxJfoWwN3uKmzJE8QZtbUSob2LBHtGbKD
j/eheumXR9y5e1YHpnSbNA/XivMDCYglhnW5tnEFNxu23px+2BAJMFdgqob8KSon/alBL6IIBGoo
DDP1jlqnJnrJMZrS/KL6LcnByds2pLVbMtxJL3KVZWz/D6nNvtGX1HakAiPzdYe+AJOhQUqEE+dr
0ARnleFWK8vvrtANpwA1UIaLVjBKo1vhbDzAWHlK5KcChpe9YXMKMdKzZDCX9ybAa/iKiV8kvxrh
CgBaa/0RlpZYYpWDdADf/rPmzXobomPsNs6CkGin0kNyIo0pTsEyRnjNuGYPzhI+FrMiu4LNbyno
tiA0hFRJPW8werp4buwWv4GLhZ/QmPY9yCXKZs6q/kE2LqNM8NHc4fQEjd1fXDJSMDI0Ogzi5l0p
Rdu1cWeTWnQmq5JtImDJoET4UTMqEfZUAOPI0IZWS9nuL4o5DsXSqLKFKx8EQzTvNGVmWaIIeUn5
/rP5Ltw7D68Aw38uC6VuRhlvugAaPlPtaZRlTCg7t8pF569hsHP+SoqhSnJbCqdqQP8jAmfvuT+p
rZcYhHykVYsutVJdiUPQNe4tb9L8F/CKsm1ZuYrLG2uxi09/u0XG/QXAG56dCglendP0++ZoM5Lz
dsNMLVwyV7il66SvJaL0v6ZLl7dZr34dQFA03T3IYpXncrbbYJWpzOAsTgMzhV3pKrNugNVE83uw
Pjh8/HRMfEyc+ROjh61/C5p9KxCvMCNZCGsGu+70C0F9TGp2Ws9hgGHD/1CFkwmKGjzsEn9j6Kvq
nnM0ihHDU+WfSB4hUEVIsG918R6YsXJLqpFHtRR2YG3B/Vq7mJbBXIEstGPIvhpIZS28desC0cT3
BG8/lTj8Yl54H+dfRcNjk6JxxSIzsO7Z36QJaUykoWIYAksCxJb9D7tLxP42CRjje2g81Nveh+S7
3uWfOHyttCtFALlTKGlytAqb8+F65tRGsT5Cxm2OUpJyDQ9cZlsCnZiKlnA/1awDA7HH2q/YAu98
EBFpXHmL2H41KhErLuDtwcLNzGKvB5avTmBsry2pmnSGY0v6yc0LCfK5k119W+GsKdjRleI2lPYm
9uw9bwX2yeT9SzAa1leWahgDh56XwujbmcoaIK/8H9NbeTQ+JBhL4/HTqzgK8nGVCsRc2qhMBqx2
eBjqJeUj4fIE+nNTvRfAptwDq1aViHmg0L/2XDHhKUWaHDWhc09Pa3PtNSgrgZox8qv/dNPVrLje
ElRTsJgI4XX6f/R6bb1mQDu/1xrHAy9HSfV8zSFmC0f4YaI2IPbKmptioUdVkgQSsrxE3z62Dt84
KUK8upFfkEPs9FcPzYhYvll3Su8T4RiOgKJ9gQgP92HulwSgr7wnpi6RVtchLSBe5+4Ah6TWYbBl
fDeb/rPcHhKPKHS3GyxhwqtjDxelgeIkbH+3Pu8yVg90WrKfPm4+9css4btVRc4jVPToev3Y5uI4
jIROtLxftijjsmjS91J5xn/zoiFG37fO1nFiF9t9tXHZF4o/ZCniktDgvFnacSCSJb7I/SRm2BBA
CxuXKr/BAXCaJQSt53vam0BzGTAj/Dlf5YGJCYMUb4xizBipGwv95lCBmVVimcHScka4Jnjk51Il
3MsmkZCaYp/4j9/WiNT+9TYbTfjnJaQIqpw9qBTo3zJZOvzoe28eWkEIBIvBaNx8qUItjn/yKd74
k5j7j9PBqMt37KMkoCzLhmbxmWV2bq+DyHT94NYAqPzAPyvgOtZstopbVgZMs6FrS7/ghsf4Kg+E
vnN67NGjKmRK/J2DORq9cwU1HoewlquCI4Sr7Y61E45cJvrCfKm95bMemxB5bAD/m6El/XuckI6c
Os3KZ4y4lstIQ8BuRLEigzVvbR1pjHgNDWNAXztYptWd0bU2xcji3YP+rC6n6k4nTRuTmS0hjYby
rUhRDEU8X0GbkGdd2kJdlPiu1gta6XJHDZhOscuiYb8A/SBHEH7DVagmFRqMIWTMCFHJ6GhK39zv
McqSd0LnLoOi+U9ua2Jj7XcN03CI3MXUgdjEMfW+UfXBTmjmqu0gVN8GkF7v9CaFmXragSMoIMjZ
EkQUggnPvBBa7uv7lD23wOcgnQftaigdc0zcrUO/1IzxCPL7j9QHpoxO2jBxCGIFKnlhwEGcLcl5
mtsj9pOr2GctDn2hyAINpsRfwdTpOfNH6txa87dnpfA6iYJvUABLumFfPwVtjNKwlnAQecnZfwOh
Ee7m5uogdE9NZU7Vi6VcpRAfdYrO6kV2sXO75tfvv6/gWaf5PWxZrTwkOHrgFv3adl2tVhb29hTb
Uit+DWlHMYHPjBzVTkV+uSeNJ0oZnodOq1hKgr4PITTmSf5eKIlUBp/b8nI/dcE2LVWjuLkMC8Ka
1RNwPErkFETsHyTsesRwMKQZ2vXAA/mBTXi0IKbSprDCRN1Fi9ESoGP8Pi43uALubnB8eCQge48V
q0Rh6Z44NvBAVtO4yX0TJ+5L+gC2gxNojd1eRUV2IHpE6izKiRqF2DbKmqSVGSpfiBjnIWMwLdvP
8Q8mrHs/RSs/W/KZIzWplrffljOFx1OSdRUUhsNquFg2/vpNHzq7vvCNGTu4Y0qQ1xPvPlotNjAQ
BeAJPwORyDLyH/XD6NZUUT+5ICImp8yVV0z0BUBb8J2B/qol2lTx4xhVe9iNOJ+BkUOPBC7udDn+
sfD6JnDChx2ugRDjcnyTrueptEWoDkrwyoOCODtBg2xleKU+jy/2BXgl4+XVN1rH5DJFeVr4YU3X
creeY4x67dxZFlm7vMuNA91VoTWHnpoUClJcRhniKtohgThT1nefmbxon8sas2bpZpUNcxqGJXGX
Q05idD5m+D3aQss18p6KjKOesjF/66M6ZYECu7PMH1ZsvPd3BZwG6J64bYPmXWU1/yU7hs33ESVh
507wq3ACuBjuZMACMIO+72bke1zJ5LzoV0C9+Ve97Yh4YUyVtQohTHOq1wG4hl6VvwQV3e+Ld4Et
3f5GHLH03cPfj1Qx16ZsPY8/X58mOVl3ap31WmiOTu3livw0heqGVO/8ZezF/ELWnFKtcFDCdmm1
JXd57QWVw3zsAdYo2l0IVJ+/0UPjxOnjAmDu9jgr8T1lila0WAWhSJyC/gb+tm9ZB/0uEgoSz+SO
UU+nETIc6BcfIogdqi0SKYLbv5IcSKLBy8KDqAAgGRN/HYPKbF4+JPwXI8oYntvQcOzycriJqfgW
GB4SIDspg4s1CkTrALRgK554xc7EGynEOOqHnG2XxbywhcLtFyZryiAq88OzEvkG+wxIhwsdSG6l
EyI/3DsWl0/FPvS1q5ND4t2BJOW/NQJ3xIgbVjyDFioWt3/epFpVHjD3zoSOBSYMwGRWCxnWdn00
3jm6Ca+8joTtW5FOuUZ312j6xY2QBl2xadcNvYz/WtXXpHlIgg2wdwCspTWJxBBHoenVzM/FlFu5
Gy4d/gk0RxixFlApVbPHlWMJ9OUpP/4D1h3OSIrbclthgy+GAtecaceV3FhlV0ctOE0ZCcAQnn/I
0flh3d3jEKLz8/xIwQNVwtuPXcTGqvYZZPKzN9I7ZhShq+I8/bzjcLkEKxt9wK83V3TWwGXQ+7D0
QSZJp+pMfhxUaSnn79m3wM6+UJ+V6be/OZ0AI5AZl3SgxCrwUNZuvkj1neHt/c40czdtKfdKhLXe
r+ozbU/kVuz1NNLMK71pK3FR68nRcY9heJAxTC/fRZQi4/Ae2wOVysaAYlNS6l+Y89CMDnjQH+NK
yWdNvEs9QpgSsCn9v1riTQ6jX2G02UWiyzOMXn+sQLaT3VElzDQmO8In+wLw+vdt+sRPMI5tD904
InpQgR9sv3GK5g45hJx5jAA5IXnTBVyFYKMpq+eM4iONOdCoioaHAlC0ScDGY+9m40/AVixanMcY
t85YNjbZ+gIcITdYhGUcsdNpm7opuWXedDebf08oBpT4Z/wZ3lO4ixsWgpe+u1H1D3X60YwFj3fY
/PLjjFLTl9YHoLtMrkCrs7h4jbUpw4G/dPGJ43aPf0+MR2tsGwa7+uHlr4DLsqfSc+kvFyeMimau
sEzaMMW9131ppptcuQtBVa47qLjoPZS2q0QPVjPosx8kPwaS5iUgwFQpb7itBPCdQpoGz/lJVTbM
5UZfkM8L0lf+mORoN/HYyT4srBIKv6GKBtvnJJpmBkBe0veHU+2OTQY/pYjlYO78fOqIKrF8vA5M
Y0KPgqRDaXPgg+LJTYb5EcLQsRnNYxAx1vWbEcVd3HvDvRdNwFo5QkxIUNrqRs4+r/6sUbJG0SrT
LFQsn6sqMGPi+hCXgBoHBeA5ks5LjfHRfGoOTKgGQoZVr6BzzjUpFJR5AgTPAFyOf8S+8cg2aS+h
xFv9NCjkFqe1nKB3uGlYYWah8AECR8KU+SesdYgA/+nOepR8sL0KsGGoboNqYtoCynjQof0yVqln
rTvK8smz/rb+fUwLfIt6MxwFE6NS1N1kAx1MjsJU5otpC5RS4NWLHA7yu6i7ii9Ou8CVPExxGcRN
XSZNISqpxs5gJyDflPf/rxQUSZzvtKiTUn1BQHri+IQUmTXX3khct/+hgn0eUsX/b2yet0xZ6QZ1
Uwg0vvMx4Qo3+2LsWPz8U8DEsCmWqwgsTZ/+cwDa9NE1KkH+caXVvy+atSPyXiq5mktOLRoLwEZZ
UTIBP74qi5bJFdZAKXUUCpzLj5h3ErQnn5Wr3K+TcfCL63H8G+DtQSEYbZAFN2+y26MkHCm0/lnh
oVYcPXSuNfnmlTmnrCn0Dm1UcTD/+bc2crEyv/BJeEtQ6C5/v2NPkBMuj5XLOIKhNT91IGc+hHMQ
MhJOLbjYvpMFxPbz+Rd5Jgj1oQ+mly97WDj4mm774tdTc1FnopzwLvOfESn7kpIgSASioYoAiSOM
CZbQv4nUF7Ly5J8U31YSQnW1gVGLq/R5C4p9tuD8hnZmjzG1Toz/QhS92OB4lGV63TzjkZ0FrtP0
LK/TeyygNiVtDNSZV29hadIUOb8UdBmoNzfc2EMCPs+FbSb8NUYhGD4qCT5W1ATAaqbd5YRdyW1i
/ucSq4SackXmWC6NWlx4HyHKsMBjpGtrA4qLW3N8/c20z7QxTdx8NP4oJyIrLAxOC8By3lrs3Fvd
WVQopRyxK7Vjw2dVXzL2xzxyPmRY3DcILU6uPNw74jwVTr67uI54+qWg0ZXyIy5zqdFBNM9bwo3x
WcjQ4mB6BvXbD9WR0K1dcUH2Mlos+y2VJK8gQHQQjmvi/zAaCpRWalZT4Ej21NBeENg2/7otEG39
3FRbAZ7cFTXXLQtcPjSgKs0iSC3sbM5FMzCRh9my/dwj8Lq4V/1cam3PRTmF0aB0Dbt8iDSa2e/H
HlU0v4mao2MXTda7LluDS/2Q1hQtUgEcydPeXfO0MKFLHrylInyJSEfYS7PzfBI2c4YkS6nTwBOg
DbUE6YvGhWmwSi106poM3288Yayirx9n0Do3SvAw3pXfHFgk0kdMGtVWxkpg8kzLz28dR6JqL9ii
YOZcm9bVJA/tBfiQrA0o0HWRgrl0ktr9OhJaYxNLKVSPFCFVuqRiJbYjutl2Zrc/66k/m0cY6B/W
ZOjQDywwFxFFvQWmqx5NBG0U8UYxQztRd8Mfz9w2sHQyb3SX6iCcxBakT/B1clkuGrh97+jQFuC4
CfVGda6PtOCawugHOj6gNobSU1rflrx1vV9p4WEswilw1D0Hw702sVahHFbjKxy0PVRgPjiXG9wP
2OFazkUmgYrGwBSNHBBrgEchol0jUioJ+Q9VvmzpJEHVGOTXVnfhyWXVJrtu98toav+GO/pbHFVI
J0Tc6d0q24Y4Loet497EOLQAOsuOLginY01csTraqRkFhEzw3A8cRjPRZQjMW8dnT099q+X1Sng4
+bw1433ys2JV8XDIk5/BGgH3MDHaPQpNKesMve0Fkakt6m5LwJYkmxhYoL06Th4HCs92Rv4MA+6x
GZsL5l3ZaRMVSBVP4Tdmerf6oVZNWuhn6FG2gRRbJnZnAcTPqCHrMSb63Kljv++shBG75FpaWMNo
bCBrsL2+4fG8/gXQi1fhWnHMDMzh7YJpkLD0UpwurZ4OYwVXgWYfu6sI+li7kZXXx8A9+ourqR2g
n8a4L7eGZ8gzrRnGe+5U9BwQazZ/WoNOIUIfY6ztnsgCDAIO1MuzJShdNxmodKMKpyKSThW5q/Ks
pFc6uC/8DY3BwcBTzsu6HUsadCCzjqUjE1uTdWnOQEEcSlrnPMJRKvCGG08QTF+zUbs399s/HQ6y
VUXR2iLtHthJ//ZFpctwlQOsByeq1mPIIZH6HPUJ6VVtxu5IsgU+9Ikm8/QQL8dC9wgPbVba1vzt
9+ADRc8njnG0n+H4kgkhWX7KFlypqKfqnuaYsw/cWESaz85GgkJjVDrNBRsAwLmTaRWtxPP8C0m6
a6wyDi3csNqPyaeX//uf9LmbsVZIK7xrU+Ci9l5OkD+pLifUISN9i3+pRT1Yxrj4mMXMpFDAE/64
oqAqirZOGVdKbzmdoRHwKoBhMGcZ90Ayy99TbLvNPvZGTobxA8cVW7oZE2Qec2PbKUOSDsYjZhcB
fYLFkziX3IqHNalhPUE6zjlkjNIBhXA5pBGKHvg8UVX3iSXa74l0hFQZiWGAiKAMkqfCpQsaMHZB
auw/7K+QVJwheM62vaV0nxX7gWDJQYEYLtXS/2fJCMOhtBS0Y2Qw8Obd3T5Kq1ymupYcpNXDAgqj
JRSiOHGPP0q82eDJgQ+OjvvErPwfnpulF62KuLr3DsTHLwWQw3pVtZ2KHOYik2CXbRW0dfxmW25J
REcmvTJS1wdngCBGHXy1xA/DL8UkjItwoUejRyDwtzigvZ2Y7xtm8i7+Odp12U+IM925rxKlpa1a
kIc8qLMfC7VEzjPZyYPRLC0Z6hpYNq1pkZ9dgaaAJRSIABJ9RegKSgLTjc1JGL7ZTA5GQdJSgMbb
f4igIighiBr7SQV8FYnfiwZyBegElFFcVnVm+6ZOcS5ohnPrO9/BMMJRVtYAs0mmcDW+ylFH8fim
uOh58PTnETTKSqUdFJkfjbZlV/4vmhCGziRPiRQ+KrtaDML6e6GjKQAju1eoQNtEZd5hT9DZKThN
1q7zGzIUtyQCpzPTYSQL5yAsDW0rdS7/TnywJrIlBRhyc71FSWeNrIGly6J6i5CW9NsORnCL3tZs
k422ujR3/7ABHaJ06HZ9t80XLMqruhQ87QtIQJyk15OfbJUmWHiq6OAHluWY18FwOL4+TnYlyW6U
PkcWNgpObc4kY76hSxlJSS+Yx9l5MSWVv7ofJCgQOq3F6ECDhze0qCX/4Dl1i5uMHJVSHntr7hnw
aAkJ1o3A8x7GAr2HlSnq0jVfyNX6VswolDA0Wqp6MreCCroXzVr/l+wdwCx3GhOkibe6G9pRTQ7y
oVvMWXjIpT/TNMLCz+GMYC9IP/D/r9x92ci1xZq6qXjDueKcy+H25rdWOai6SGDnqaw52WGziyKH
eArYo+9D4hkcoVbWorH/t51xZWGrr3o13EJVxFdTxsWLpux6iieiyRQMP4wdsCwsBLXUlsbjxTAz
D6Ey2zTkWpvCwLU5A+Zhy9O3p7tdSiiZkppxRm5M2c9RUDw3KEJZzlfDWx24M3V3VD8iTs15Z+jD
aLHs5jwUx02vZFd0bbYlLZqcD1AvZEp7VCBzIbsF+rXw4sgRWGO/eYNSyVYsW00BVAqesdf1Amho
pUBA2NVCZN6w3D0e0WeYptIqGvdkFNlxI7Cdi9YIh11sQqbzt+EuL6MRaIblWGImdpfMDqeTehOQ
o6lTU8z786qLHxYJjctbxsfFlc0QbnSwBhy/H4JjK4UrR7F9A6rEoBQfDSfgDVIaHIewmISmKDxt
nXODlVGYT45ve4CiH2Pg7mUdmTgZ8EFgY0pjurVRR5mVZJDNDzFF/gMVwG/tcjhX8ByH1I4nVx6p
xMvv+2cyCwP8l4wbugmk2MTHBQ6mA7qAocV4GtAhH3iVWT9PyriV0YV4DZoy9c5xXdbGYwF5Xqdu
HOHlpUsUAmIVUgj8MA4d1nBPmUfOmGnW21KIqwb2Ug/ev9JcVqzJDuf1WxwhalJByKFxoojmIDRk
7QzEdHKUnA3K5el5GWWNXm8mgYQ4bYaxbsNH5A/W5h5ubHjUQfzKzfFdfwJcM5A7Dupi9uAm3fUs
avpqENM+DoVCFCfe6hUB9w1uu0NTOMsvUq3Vxtdk6DfA2pO8XjRPfxfTuSCPzNRxbl8rjxZALprh
psoXPvP/OF4D1w70z8HjFY+liSFyPIuKkknPZFZt+wo5aRSWYckOd42zqabN5ONNedhwiRmxW3kt
zBqvRpQRUAtb36yxBf16ozP9S3T2dqVahXKe/LdVqS7uxjCpdEYG5RGm7fATE1tL/cs0LSMHfHbJ
ie199NHEgxoGtGbj6/kwWKUy7Y3lQJ6DZDnSS+1oYOuyHw5YHoFJya6s6MxFsh2XH4FVIApefPF9
Sv+iEXeuiVj/Z+NiVShMmaw3Tah3+XY0aIoKsRhyYaZgHEEF3OLbTLCfv4rtgIXlNKIBl6WOzMZG
YDEaxJ9d8bHp4jdyJpUVtAz9EhmD20cZJ/369T/LbGul9fLa9GnJOWhx2IlzHF6Az9WWzPMpJf0c
+2mPX4sLE9Y0s39iLDzOYEzGXRCPZ3QVXwaEQ3Prn68MlA40PhAtyuslRWNCg1X8ZmAJyfUYuLb7
qEaozIucMMnUYj0Ghv0DHWQI9dgXdlN/YAcsDZ3ygtmSQPn2O66+RtHWuAIFG7nqMPAKwdXXMoBU
RUE5OyOBLzTHLVSyGibvac7OLetEoxqr8ljmGwMgdk2LUlstrkTdl41UOdte+jzQ4B8J6H0yaYZZ
DMnzHCb5TyhF3hNvDuNIgjxaZ8RxKuLymNF+p7U/WSmOXNvHChBZQzwn7zghDSmrhZW2zVT+T5Vy
zyil9oLLlKhSzgPF5WpzYiBlQIxoDLFNmJD4Qtyy4WyN7Srz0xKCeGG2hw1yVOJa7fsHkHzmeVmj
ho/56czUYx97MYO/txDke1J1q8natM2SXHMgGIPTz2OIkUnHNNodbScO7k6m1CoTkAr3d7CqHlj+
VclMkPAYwxtgmvDL+t0tOdObxCHW4zyf++Rdzy8dn+Zs5BmRXvLujD5lIeAsCXU5coDmcqyznEas
J7hVlUojlm7yfX0dB+xjpY6TB2F0Tt4fCBkO3XyBYMmlgALWj7/qBsX4aVyIIXxHtzmqHAfPaiwP
HSBc03pItHgPcAUH4UyYysCePkPU4QtDzZU84pG73hqgQw0XBVf7e3RcDITnPu7NB9AEB2jt6j/f
0LBA/w1FGBZNEp8Q3hbXk9Lu5M+CpAd8Flnv8cZYfpphKt7gyn548uWPbp7W/8kYY8Dvn0ylAyg0
zLHBNNWcNsMCtSN28TugA2mr3VvywVtStT1CmPo9ZRQfQGqUHm2gtVHfmD96uRDM2uVki3O0x46w
2bD37KB3qTjMZN8zDga9NWRRvcXqNN3ehsm9XLuy725yBF4rBnBJ/kLvP/wVx8J9682DFBRg2qxD
8QRLRxDaLR44nagbblzBkJWr9btiDJrSMHzmkVxnfmM3C1v926EB+YXUv1c9hnICU4Xj0iSuMmhv
pk0ESq10lbpYBJEIU/KRBjXwz64ABkx09WWEDuXcJUqums2YO3SaRlqFdQIixL6SPxmmHfMo6Ckh
R0/qme0/tSNNy4D1foXnUfEGuDgusDAm/EN3ishkSVKQ1n4qMyJjZA7xSU8G0r4kxmXMYWyflg1n
mXcXPAH7fs4gZEIHfanDRnwfPIKpM41sHC7SRpJaqMzOm90Utmm2fDDhjdtgyzsgfKz588YkPA2g
o3CT44NnGYjaIDnGejiEx6PvFkSV7sPuBBuTxLgNhfyQOZLa8wi4xMdLSfD8GBH/K5acr/8LYnc5
nlamOTmZ/Jwm0OEqhbH0zIXg0Uv54vaF954EBbwhfQPC0HUAIGKS5s7mKHA/xqPD/ZSYE+SGONOp
XlfsjB4/40gNvqvja3BXOITf2zUrtArou5wkeVO90FuXQMLighel2BNp/IbN7e/vwCQNehBx+7nZ
reOyELUihXopwpga05JRFpDa1nLXF5ffJSI1eJ86Hp5DmKdjExZMNQD90m0R999WRTuH6szoktTa
kxqc2ubLSqekQXETc7EB0JKHDVoOJxQisoFg0N8MDOZKd1BOMYzFJCWTD2AGNELyXAtnTrEYq+6M
EUtfzlmgABWKN4hKCtkTJ7LmAX/OMC2EyU2SRgl4r5/wj07jp5rHEU5VWMt4MGcUTmnC3z/jnf9S
rBWvGO8wV5e4Ty7SWGxGUsJBTYCnRcB/qpYY3ourEPNYzTyGPAIRUQzPrgVNlMBVB8vKQvEXwaLw
9UE1MNcQwKR8D5vZOOXdERv26/Ckf8DdtTTzJoq5sH12DGNA/gwvWE+kAotXcusOetsgGjiItlr6
vYTqO7jtj7+axwd/2HIXTUb7gRpSikV1y4i1pdAg7QWWXwO6n6i9GU7lqZJKFC2JJAWAyXtXJzex
hWrRANSaQPnXi98GeN76F7BRsSySAcLUgy4GyM39Aj7VnnC1SeHtOPRORprb2oCQ7Uj6zX3XmVnw
GLtvUPXdSHM46RJXqcVV12b0MVWhtPsymq80uQ7GShrPZR7OwGmqamiALdRHYZ6KHrjJfpABUFux
31gZlZCLQTdzTGL1a8KwQzD1QlB2FwClpPEsVwXfKobhKfkfmCQp6WDL+VKoX84GIgYrvCeeFF30
xsfsyflMPZSdoPWclw9kquPCnDUAiB9QLJX2VXQbfFGduTuSESpUuUAEnS9PZZX4i4LPOEOCkaVR
6Xt/jGfqNgTrKA7W24Rge/hWVa73E+RyoK0ykRkwlrFgm2JDuoBqBmJIVoeL06sKcBZqJ8iuQTab
eDAD5DLNbCbpaRt+No4/4dL+u6KS6Z0D84Qo70tTsMZpGKdbH5NGCfkjNrY9f66Hsh0UrLXLnT86
A+8O4Iw8+qrzSTLpcHpU64Prcb5DrYT1V/SWgeI6DtQdQIDuKaXtEPQtYhzszHlrxzEBkQa8Hnzc
KwhZTrq4XH36xGUzZEKCOUK73LZDZp6OgWa4votQkrbXbTOSn7GNwmsSejIXV3Znu3n9MSXjqVxv
Qo+AOlr4FXmrvZ6dFd3IOhiLjlHmt+bFpPMFiyTBB7zp3U0K8AxJknjhccN0K4eU1jY0aOUcvZes
4fT7dwG92FHyZBpcIjpPAlGVRAMp/Ggb7LdtF3MCv643HBJ0beucYL2ZewLXMB31YKTF3c+J/pvE
biVKMc2OKBeTMZH/V3EWVd8bopGcCb5eeU6NLmup2cFlSL7CLG8Xr364A3KEliSCT0GII5BnbpaD
AVWcdu+IHPPCCak0bHIRWtBgfPuCvYFsfNDiGYCTAdE59Gzg72ym25jjrYApiYEA1A0NkYlGg43s
js+P6EFs9c8MEdgxpxmeR8j5r+XwO4nPZqE8JdLlnc3c4dTiakyJeOZU2JbUosPiF85BF/pXRXWZ
Lxkv/Jpml2fBYuZl+dVm6AJ1J5oRBgBxXGTPf+7vw6za16pGwOBQUBGb0fbgy+JYt/vg4eZe2Z/A
6hLVQxHJc4zAgBkarrYeMDOh5lssk39rr4rr46tGO1H9H4A8lyDilwdpb9N6JWdJfzqA2EG7+LMl
708fQmmFsd8qR5C7DmHOZ2AMUr69sKlLpZxMyRsWAh7F8YP3XTZJ2T7TtLZD3dtLqhT+zOjmhWRN
6n83u7Jbwns5EckbEIJ0l91wAFWz8jX3nTiPA+qHKs3Svwoqfid82h41Vvkn2aDvu0aUeObImYRh
kD1zRTTCtrRIxrgSZwAbdohOBJ/sSIfeHvedR5lAmeGVqlp9DDABJk4LMPNh2qyRgc6xjzEAahQV
aypcBAK18bH69/GM/wyCCgsPDWMXhRJfk5hoiwkTPSHpGvoxNTIyZMo2iDGh95j5LSZEyIzxqb3z
bYVmptFO2ErzLtVAEpHRvye7L+LVatlh8rmkY5hzpXIEDkne0vBBUL8lH84lXtCBp62q+Nrr6Fpa
OK3htFha9pnMaYT7U5BtE1Cfd4iY9xHHph65gl3qJVr19whvcCwImM+lRYSIRL5gzKUVAsI2uHqN
uiWvCG6ne5yKg/jj+r14BMO1gBmFl7ytl41iC6kHF5M8qXb5mTUt0rBZ5N58jaql79+2bd6++koc
Q2yTy+kvE+OSwysG/cwbLPHESxkkmpQE28g1ac5/SCh8eDF/sFAlR4VwGvU6XzX2I8FsKyNbfDPt
tsB359a0kMcgl/rHPEE82Q4NpG4gZNzp6gchVypsU3GMJuBkVnY4Sj2Sf+rVh8ouMbXBISoq2TNJ
gE6dvBe1mEpRy4Eqrvi90xKHUzFKx6UbQoxRafZUigUohvs9sZBzsTyavzGZLl6ZUHBlx7gYA2BJ
SRKjo7Cz2vlZ2iya3T8YgbOig7fR5B7DE9TdZzB8uCCzod/k+ZGqrmD75alvNfpTHoHJqLQFLz+2
Uo5SHJof9aQRHKSiKoR3KrFzFIWDSjntAQU/Fu540U715rmk3FJT53pjYBBNh8FzEMI1Y9dcAlay
mx4nMqyiCUPEjR6fKZi/m3U19u6kquO4+x1jilgVgnXZ2aey/Mb1obbB8YY0e9prnKtAtj66eT1I
KKA1j0HL77Clz2MFq+zNzsj61zbYNeh5/41ZFhYt12lGvuLF44NeuaI7TmMSu8Z70biz9buOhfL9
XQ976k9M7FGiJH8LtrTrde6/r7kmX2VCF4yWlIjP9ECsa0q6iI/9OB09QXmJ26WreavX8ht+A2eR
UEDCHuU+L8dEem/IzZEnRqEL1YcE24X1bDy6dKL51Z6QxbrlFEBA2iE8maUSWdBt3X69EoLBdVIV
s7AodQ48o5ilcmrQUwhavoWMbuTjNXek5Y7o6SkBkAXYN33ys6aanf5IC5os9cLODO6jhSCQgBJ/
wX5oW50KMvO3UJKrdBpDwrciN5IWhu7wi9vSwDMYaYkok8P83TdvjzgCdVY6vH76ULy6yBTStpjM
kJ3i2WhNyr81cRGJKXO1P0R9ZllQKuX1wYc3KVoPKZeIS5zcOyFlYnXFsp+1g8QvMcvKfJltJPd0
AiuDR29nG4MEgTR5N8WxCyJGyznKt2eXbUW8Sf3P3TozGdH1GNU9Tn4tzawfZuOJBiBk57+cBcYz
LEK6Ump+iOTxG1JKm2RjBmHQEDfolC5ZOndI1dK/gxZleVwpnj2DzQqhFuZTWfl6vPHawdh9gDSI
/tRhtlt+7y+4AknhqxPTRy5p+Lrwt8lRzkJ3mvEzQcCpKvhgW1SO+qEfNoM3s7AZ/5UdFZMdzAnM
QRSkRJLXv3hpycUbNrWt/Su+AvLQh5AlyUYM9kMZ/UPHazqfMRjmlHkcTH19swel1mRy6STY38DV
tkM3UwnWP6SnZ8uqMz/ePq8a4RUxC8VTQ58ocsF6yc4OBu9Wnr1VN2Bcp/ttfa9h6mgBwukpwNPN
fn34M3VobZLPAlziyDXuTS6YODFwG03Kxe+lh8ms5swxT7wvy94BbsD23ELddRCrIycurxMJ2cz9
rZpm44HFyvTDNzgnELNwAkNTZ5rhd32vlwgSf/OkgrFBE18zRbE3yTmmbgwhNQinlUxarewfJACz
DUc4PNUOWGRmRZTjX9ubqNSda+A3dybRcrpuo52BmIOp4aSxp0aTg9Qee+PI4ZPrli8jiVGza4za
ddeQCfZrz/Ht/chIQ8dqQl0Yydh0pki6YySfwXgEjLaUqRBM2yFrBfjeKPdyjJHRLkxHeNBEfDET
tMQ5PAEiDYTSlSzSuuQxnHnE9UnC+nLsBTttqJvtELcGVnkPQh/mJqNr5kuMguj5dEwhBPnDUifH
aVyqJn60QrmSa/06VXreL9ifMh/udko4zUA5XZfX5FpuKa3OdjYiG9Tapm9HoKzIsmpLsn2i/rBu
NQFJcdcGVN4XJCwPhFXxyF5l7NO2J31LF67QTccjU+XaRVSIUuZKxhFHesVRcklgpJD32qj0jct9
Q+uVzaek1Nn4986D/aZ7u/iOWH27YTjBnnziLkBOp7wd8BBM591+bdCa2GKz53cbSkhbafl9+w1U
o0vL9eRegdE3AGPQPKXdbktAjeNQ9fzAnWOvnTfFlhVJExia4ikTzBi4/Bw1w/LZ4xobJC/1DFiu
gT+GLMmLHAlG7jRs9OoK/s4S3Ik1EvTeiYOq2ZpCvw1tYB+CJuQYBYIWYksfED7BdLF/+jwTZJFk
x8DYpanv2tfOx8D2Y/ECZQ2huv9iz9WPKIPhgowM7VLhpd0tG+NFYknXs3xNt2jYT05vJuhzsUnf
mO2FW1nHqKTElJAERFNZgPNXwaEYBDfWfdrhfysJtUzmCyD93AZ0j0wMS9ERvg2z4QTsDSDnDDYP
+WPq5YOHSX1XAxpWUk9r7NEmdl3lqEj4z75gW6gq8hzAEO9RMp7jir8TxNSUWguSzJfsl6xL1nE3
wjqSkqGt9S03cmNLjmKuUIU3a2r0DsMPb0fi/YKe1LnYijZrx4UeLuHXWxsMzjUC3Gjk7pjZMzKH
T+yVVLmJQ4xs1PXtk3S/F/lYlbiX+nRY9q2hCVEhE5VfMRudae/QQZTjkB25DHSGbxSxxWSgPwc7
VjO+cn4MPqBvDHkzm4loJIsa+nIVHoTOLfNMyAzN782Q9QFfPz4dX9dI40CzhLfaXFmzkFQ3nC0X
lwfBuxS1wDtA4ptqFDwM9pqieZAucoQ7p0cMTonBP/eBgKmw6baWV4RMqLzegLjvonQr3DJo8Bhy
951cRh7vk35PRO09JkjHqsmhoKqIF98EmjTDV7eorChS5AFGfOItVbyI6cIQ/YJagy65nUKAmsJi
b8F7tpidvYPQkuholTnPSAYowdHnau2zGJg6YIDGvu4kAVauuPu4uWHu24wgjPn1KlCe8Irwtzy8
MSnKN/lXBU8lsWTeWCY5bwseOes0+R5cKSMpSU2vszXrjNRaFXeDYzGq5enlIGKfNGSZ0ktcBYXP
cWe/7C6X7P2KjKaXLK/c5BEEqpwk01wTOdlOoC2AT6kag1ldJgj5aFJESwA+3ZKnNtbz5GzZLl7W
GULTIb9dZ7+Vm7vSEEl7WmcrOO2bceeUF7/MjmGTTAxvAY5taBCuADA32+QsrLHCqJDcOteFEVpU
sRtkek6dqYz9IDLxPVZz336x9qCmL0T+Ysj5uQStge/aDyXCfAu53qgytXtU1mosCfu64ub2/wUX
UBUfjWm1OTvnOt7OxBXZRzzuNlHh5XG0/8WCkRy9eWZnpaQM8KevPlZLBzy1iNngxvd692ERdxeb
jWCmm0HPjGGy7nNgrhdwb7tnmP5YkP6rYxyoyqyVMouBkAt4ZGPxqD6WrUTVYtAmFaIbJ4mvjPHa
Kenob6oz0DmpjA3kNKqnFRQYWDA6+0NEWc56BW4lVVVMmEivviOtkS7s1zW61MyPa/n9xHPBcLxv
vBfJsCy+ACOr9WK4OMinosUbtvr0IUlOHQQa6yfuicxDzp1s7vAS9w6FevGwFyJZEpDQgHtr1iba
i7q8WjdXLF91jEXskzrOmCjxLlO4nCfueeoHSmHOeC1XXE5PrhydOZVGGfK5Yd1fgwQSVHAX4RRS
SYoSQaiJ4a3TbrqWxXbdGoLEaanE1UyvHS7ppzYYl2ku3F6I5UAZUdeA5IjO9BN4w1ynnTQb3F3R
B0xVn9M0uO5rwyMj3KUOQRRu+uHkmk1/ClFHc7HegpB538OL2uryN3cU2m4gpxQqSaLRhbW/rKo3
v5LCfOmAIoz1u+5ELap8qwcfZeyFPf7K3J4+Ub46vrdExsUjRF5KHACeopIhbFUYYKW7vs2bnKyW
p0a288n3YIGBKmoJQhm0YGFfZsqMXz5+9sWJeVz/Mp3denxQIjzbPc7V6Dr3SCvLmBxzCsyDr0fv
JE3gOid4S5lC4hoqwss6o7FE6R4hWgOvfwa53wF5upLt3j0dEXO1Ep4jEQ9pUzyo21M5D8s+aDWE
+nFVCPlX0qD4mfes46aQrkqyd2VHS+fjsOpbucb+AyuXWSGZcsy5k3bBsAsIk0pVxlEVPUu2Mu5z
XQQkq/Dlx65Xg3is0nX8dKR5oe9mzoOEKnNqx4z8rv4pmOLT2R1hMinuNbciYjkzHn/xRXNzl5lR
xQ41JWWblS28geCZGr7SXz1ksoaFKkk8uJqDUapvnUr5wHdeGLwgLGdQLeR7mQ++OoJrqYVs1z6o
cPpoKh0p5OtklhZsmQVFqv2LrfCI8RCS9SrO892yg3avq9d7b1Lpc/oXHN0MlvuHNTXPgCrUQIAd
yLRyJrWUEYu6DxISM6BxBKILAUEav2Y+mC0iZwFWtHjoE0NykVWeI8p5S53atX4SVgiLX7pGksQG
MBFJ1t+pH5gdq/Qd6x5IVrYHAZCZ2AGzrNg9LkmqmtzzE5NnhoJWFtvC9xMEIgzRbxlJ+aeQ16TD
9pw6IRxTvdZlLPtExPw2fUnYPsEM3wruvH9FFhtfHn91LEW5PZKYUAfWikevB6YLXamfE/00uiDf
ew/uktB6KXzp5j1/sZuA/MiF2eXlRJh2inpBwZRcfoQMw0LWkF8oMdI2KU+uMSBoYZTWMDIvXxRP
KQchwUwRnnxw5ePvKXayynG0As99SKwJVXMinZORwXpFH+3ponk0P8c4E9H9oe9B+OZDhVbpUZRR
gqbnZeafwa/8uZvP5ZaHNxucSMiDl6bRR+yq4jYckS5wMvJl+/i715lAcatPJuP3J3EItBUwBxOL
hZ0ZtpX2WoOxpGb2wU+7F5wDjb0uXMAyOiPqFx7m+NESvx68sSNVMJvJlCo7YeZqaWa3Ve4QSDQb
HMuveF6Mwka7ASOC4M8DIPAZYsojQN/H4J6r8JzbMIV31MfvmqZXPvNYrTzrS3sKHn51V+GP4hVd
X7w7r+pl1ALlnALFo5KBZxGUKI+FuDDX6V6J3P+A7gX5a8/kHIK3wvhUjV+mSJdEAFw088MKacYJ
Nby9HvLSpg2HHQ9JfJBor3TcAClomf1BHXGXms+HBnGYP45VxcCESCv7TJiWo3GtPHIFc9pg0Kvn
BqQCuOwHWn7VlaUPGMiPCsuCyu5w2TbTWcROxPiHf8ZaO81/y1egkj5eqSGsBbiAJyvOz4p6PSVh
/GWG16nwVJSEPLBTBefN8v46YtfJKxa4g7NbocWaWuBNBEmiUIu5YFnRQ+ufGxQXAnYUVg16HZHC
5/2lRXe528y7ECiTQjwcWeLpIdyJ7pm+JPs0zLNTI5aclKqs9yIYtuAObR8YWfY/k9Ip0su/Q1Zm
Hfyad4iIiNoGvO0/tCUKW2BjOR/YeXryUtcHXyRe5DpmJnzTr4/0Km+8BmuBfmIqcqTO0D7pj0EQ
aS1pmypASDbHtJHKkE0QqTmtCZWXS6jUWlc+LgXSTTJLajSechlms7EzvbF39FIbPk3HvmOifBtS
HgOtQm2dBVYmjJ+zu4Z8wliEMNDoO+rUpabnwpHjkH8lvoQ41vYstetcSVJUcIu4eK3Oy7Jil0YW
CSLVlPzmKScoZ9HkLJ/W2k/RIRCNuYgUk6OKFwgWSh2H5B3TilOPYzdH3yxYitaqHJ+AGWjFpMlt
Q0P1qt1fxWTwSGFUBfsAcemEK1JLt0Kl2izzgmKTm8Z8vw0J5cg1vRG2bfWaHP41G4VQpECvuqLw
NTZ32MuHDS0T3Ls9tMMsh1m6kYoEF671RS0LoeR7UOvC4Iiha3qjNbW+JQlcaE9mC1wdx/SIbNu7
8BJkyo5clOWDfs79esI+rwAbsObV+c/Jk05pDWMmKGBU5hu8eyRP/pJCtqwU4N+H9rulb1e0u5BQ
TeUSSDJfJpt7RnXpKi9vV797kBPOK/V3Rze1kdv+Z8r6pa0uC09Ko6ZGFPWLjwe09asAUV6Lta3s
mRlqGW98SEKJKeMHqNKdPEDS8UKyriiZa9aikiRT25cOuikuRqa1YdNUMbmcj/oA6zpu3ZKcZuS2
Igff21QlF+LVKsDJ4ICZrqbvKaeCdkI6gYXfeNL0XZA2L53cy+aVXK1YdGzdaL7YR4q4g2x2VGNS
3wY10vIuekLhLZrjsp4yMF7/KWkbHt1JOatvCBl0b7pVvuoLUePzXD7g410Vo2GO/kKJnv1vczy6
I8lpUKnonwssUfRkWvr5FqqeGe8w3OEjWv+zoKgSUws2trjBqNWoSnkMEoMsdUQVdj+nPmQrXdE8
t/lDZytDs4Dlshlj2FaMUf7mmMyNd/tv7lwqcpOlMj4m8lOoop7Skia79rPtkAtACTCoKVE8b4oM
lT7QvZ9ts65xnKXEfEyFr/B4FpQvcemjlMvTriD94Htx8g831J+xj2Orx1qsh0QI8Fr2tVElW+bl
bxhVW2O0pgLuoIX1vGIEotr6sEN2076hfY+Mhh+Qr4boZAHHA/e8LwJeQBf6uGJbIUo26DZey7C+
9nLMoHXoWcdm2G0yaLVJpzPGLD6C0/oGaFpcNAxZ8wFNWk15+dQK1+WwrChlQ3SrhY6gr1wOrcTR
7xBYoGSs3FryqOIbnoJ1d7ZpTQw7Y02XOFQlKTEuDDNiaw+xzzPCjtV3vPBPkq7JUwRd3+aPm32p
QFUensx8rSyu5rcIkBkfRLi6kZyB6Fr8lz581GpmBgYnQreI7PQJzM/vWzRnMvntHrZ2E1Xm84Zc
qOEpq5HiTLvCZ3yBBrrdeNqXYUYbsF1e+Dh0KBSPbpk5PTs4RZ++dnO7zsUmm5YcQP6cHF3JA22O
5G0+s5PzJ9G0ZDMKWI8vobq8+WWvBzffLp949asPzSd63EGCnR5DiSebmmd291Gq4/SzX4q//nL5
L3T72kmS3G2gTy+CiNElAMRrp6RoWKLvqUu7otRVV9WEb6MwOlVyTujxT9pl6WrVA0NvXd6bMGqm
bfbfqsyMN5JOsy6jUZdmVBvl5Femugvw43SNE/XeVk5lv2ZGh/RF2Aidg7HdzXvmBUpmaQB+GIdC
K17UJ4r1crUIxP8eY3IMntnkHSPpiAvHJXBm5VWgzhcp2QLYvt8sJy+XXzSphtFh5+SI3KAfGiRq
Wx1OYgSf/fuL7Pl79UvThZO8s4rR/Mu+G3Gnqq4elYaIOyKpK7KybugdOBI+rZkoJTRmgSzoF9co
C9BnaTJLFEtnXaIk3dKlroKgaXiGOqI3wYnuOve1v8kHCL02NxecJ4akUTbLSff0UwYs9voqSTJe
c4/weL2RF8o4S/1BBrPlScDcAxpGwW2AkfK4VDqJeMkM5+katfP1fqs+Sm9mMbNm9laCp8AC3ho2
VS391MrRyu9CpBmnUL9oZiIZGzm0mf80mV6mV6Y+Z6UteG+uzixnoQybOIUKNXLnOnDLj25PeA/M
zLBjZE6AilCZ/mAj4LsyiqH/8BVVOAzT/cAL4a4wtFSO9J6OM/x+yuZuvHutXfE5aNyt86thufEU
0SoaDR/6VAVW6SvUHCBNQdfPzPa6r01ihhNrjfC8xEg/GVzp/352nvhd7LCl7UiGFOPAy+w0a7Zi
O+zcIeS3ybVuf26LamJU1doFyHBeMX4oa3synvOA65ioNnD3TcI/nPr96LrTd1DkdbCj1EOiGiRU
GEVBTYJiG8Kwfl8bPfmaC8f8SvZMZrI0tDJCmIZn9pA1FjkyDwtpfsBmi0wCoPWoDlrfhcMRS8J+
3lmXj55yN5RhLokzTulzSSokcOAg8WgnnegLGZgiKq4F8y6RKjlohNYfMDGkWkv7VyVQOUaak3y0
3b2TV74XH3Vdrgss/oX1BolZRwrZJQADV6T5XdwIJ5j6TtnJpVavJJx5rVETIAgugw9lNlbFvBeO
eqW3VVp6W1PSWDWzNXdsKaBSeqq1On3xhEHuo1l2VWI9vAcboB6vOiCiqeHcBwPD8/J2M+CgGuB7
cbRfdiJZ1yG2Jk5X7rWRRLplJvZXXSKlnytITsaYrI+f5xr7Rkx1cm8jm6MmcLft+7eF7ZzAJWFY
qzKAA2Uy3suAJwBu/MUyGOhDEYY1z1qT+Thkim0nLsd8fjklKyHdKNLc+6G7nG1Qo1pzzZqtkKJk
Mh2hh+1LU8/W3I8dqnsXcIkflILim9zl5nYRpVYmxszkqh3HkaQ1rhYEmqh1hFhI09TGPs841pRh
UhlKFvo7Fu7REI8jKeQpDoOmJalTzkUVcNzoqPMnIS14TzMBNbLHCTpbtzdA5CyAnlfax9V3Xl/2
VSDA2Vgdo3FKVkyCIss+chQop5enPOv6pUNBK7vRcWlmRy+ahCvTiw0j/X5OIupeblDOGn0pYEq8
PpEBCFL1qBFx5838jJ9BY4TlGW8YvuZb9cVmc2KyzWONi+ZCKnd1DZ1jigfYQ8DtftSKkSOOkXgi
bxrIY4md+xfynCqEtq90fbf3kedJ6qxKtxNWVRSmuxeZjvpK7fHMawcy5h9MGJgRcdo/oKrvYI4b
WHZKTuZhepX8/TDNh+6pcaRiqBwmt7p2JfQFZ+td+IwL8JDFO0FVcgsoTpy6rWZmw/cNMrG/BfYr
yrQ7nYLvkaNPhK1dNCNdJrx6IWGF3Bcr71mMF9z1cBRmN+gbrE4PuOlS0beBQYW3KkpiieulljpV
uI+wRMRoCKZQSAALywwPmtoL+B7A9A+yPPjK/h8/SrSu7LEPyB+FxbFpv6NDQ8v+BDiJ5n4fjtoJ
reBgMcJOc3ik9TMaK0jqgu/EB+cJr365t/RYj7QyuO8B0LmZOiukyZzN8DgIlx0tOhhmrvP5T+K8
JS6qI3hOxsp5YVyaaMMP7umvujIyjz90gWqqJ8Q7r1+KJLs8iavixuw/hCP+sw+DuY2jU074CWAL
9VOD+0iTbcSv3M4PT+EELG05vRUkIpUEI9WNER1JPJZdPIaWjvZK2i1C/cKpwtZDNmoHPahlDv9t
FlPUspWSv95wZQA4y6AMf/R8MMoHAa4x7F+5Kx5gr2ORNvWAgsxbcC77AKYDlhpxM3Qh8BmQdG1l
hcvzQi7oEHr0OU6X+ZqjsupyDl6aj8EFn36TFa4DX1yN+T8eMw7h54yEhzbHhlMLjuh+GIIDcGa3
ie4lbEBcyX4SrrmYxgY7qSvJIAUVuwXWd5Y7keTZU3LFx9CNvQpcnLNbYbYLBBSBUOnEqsAtgL4R
vDRnked2Lrr+OgL0yCcFkpH/1OP21EJLaYiejoFsc26O0dlTt5nGPYKG3S/R09knK+/bIiWqMi5x
2HquXfdIsPJbwT1VyhMZrvx/1LstsjNGfB4FtC0ehNOvOAx6ZMFHAMEnpyPrD8/sGzcfBUNxVNoy
XjU2VBxje7DcWQD8wBgTND+qpHdXVDBK+ayS669KGtLrM1x3bP6K4pM4aljIXJP2sv4A9jOU3VU4
Bowp9INIsQ9+ZFmE9kutObjLZq8eoiAr7Twf4LdAsyZmmfywZrEVR7sQv1xMuOBwvyVpfAx3VQjx
mmvVK4Oz3NqmTFsVb9Hl4Ucw5NmKXQvSdZZpmsGb1gaUojN5nZIwZn8AVhzjcY0y7OIo/0hB8gju
JsqJjkiSWBCXgNkQ2Dk0Y65nONinY/wxJKQV6pTsukc49kxyDN3Gyz/7w4fUsCdPWmFTSffUG+zw
6sHnnWI+7mWBne4exlh9xAH7WJKs6lPC7wjC6G+ZcPhQmd1+Y7fBUtFqRmIPyzrOhCLEGoNgJR8D
9/EQVvK3/1kJfhmyyem2XrlxztZnay3avUP7g+t8JrYN2H9Lpnmx1SWq8IoUkAXbnRAtDbv0MB4c
L7MkIg0KT0sxmbYUI7gAgy8YHi1rTLJZragX5ObAO6REilegNN+/JKHc25iBv2aUBTsqzF1JFh+x
ud/R1XBtUjN+zStGleI1JyPtiaZL4MNaYwshZ0U0JGcQI1+651FpK+Ev4EDVqGM2UJ5F9SE8IdFe
+0J55PlpcRjfK7XCg9SpIwANh+5mrs494gbP7SHH52ECM1QA5OwWXFS/uLtF+auUNXBEEA+w6KqQ
VcvlRTDx5fVW3RzI7obfdJh8Y005GE67TuMermRi8BOVBrDNNw0hrbSfk2L5wWMs6aJ1BtEfp9Hb
vhr/W/LAp4ahz7ZrV23Gqsxr6DH+HsA7CH7UJ6ML5y+76vni9IK7OJIEKPa4rbibY1odSNlrztnN
b6mehR+9b1wD31WCLRseuY6rDvfs4Ix2wHACPEkUeBCiz7xOUq1JUHt+pBxncgbjKlI3ael3Onwc
0cbiknT1LZWsi4EtbZB/eI0de+lgVt3XHUJR7wStdjPej4k0Zxw3zWkeRuzajLGXg5V28mqQHC8k
uqdJ0FqGDd4vdHPo/YpCWzS/C0khcbq/ravgNT3mWNCaIxYgY95+9whWZmkIOai/o4urkeTMxDjx
FYaaxjNchd/F/o4CLVY7Af8tzJiqyn9JayqC0mXWjI0TmJ2L2f8zKdVeMlOdOO4KYbTyvumnobx5
AfEae3/sx+EvTFg/M6rU944L3l1u0fE/N/DsGYx1RmzFl6PN46CTycTZGjAvisqSPSB6b0TNKDSR
EsE+5ykTNs4XtwnJ2CufXAIxzgqLgOgZjKbFigBjc3oZDPcQSGZ+C2CMvvGjw5wR3TxyD222m3ic
2fvTD8GnTflbTXCwqge6yr+JlWUVIVN62AnJdezvJDO6AOWP2a2B4uZbt+WplnCWvL/hdzesE+R3
vO2vSGZvgM9ANuDlGG2FAG9PrXGurRcQTD6X9/c37y2P7rRqXpWIzqi/BNzEEymziIUKBnsQnRQw
hJni7qrjDcOIg/X4+Ok3rijiceeRDyIu6TntuvY5Bk3pvQuGE10wQ3fU9VpWpxrUrleQuEzHsSpF
gBvI+dd2LA28j3Qvurzgm5bUp42yjPARiB0sfUvg55bE6cAUHeTbrUopqRSt7HSzcEyj7ncOAWaH
rgSTA1qVZ82a7y5+dPDhCEozZFnvZnVql20YFTCfZvVivm7JWQmwsZH2i86qhyABkfhas6vNUDH7
8c41XF089e5B1/8BjskVB/kjXUN01JVPNBVOOXuWnI/w+h3rHGN29jDYsfEWA8zIApBRinP7Qhbw
jDkfIAX40VWckI18HFpy5FzORonq65382y1iRtFayjSdXyCl9WnRjTaopeASawm/Qv5ItsbeZ4gD
L4C+LveuKjGSCepJwx2TL0XdQooYw2zp/aKRZVi+DjcwjhiOOW0bPeWGLoVRTauqmddMTji5pSDr
pGXoITBvxZOB1vZhp4Hwpwxb0YG4SPM6lDl+qpNEf18OeURnGCgIPOYZx7blgNI2e27kXI9jesPq
k7jxc4uBXshJwLV8NMKoxJ8U4lKXZonAc1s/34vi0Tme4mw7JeqUf+dRwZxkrWQ1COJx3GMo39BS
e0+iwQH9E2e5HKznNw0FfwpEGwF35GywWt/L+rLfKMZy5clpe3Zz1CFjHHPrWIYNSPbthgJPM1lr
abagEn2ufxZMfy0tolkL4B4Vo3SWC5dA8qItRl+R61kGk/Y+6X5LnxTilf5lmKpiCb3x5iHpddfd
Q5y2ML5KWlX6wpqfnNtsa9jAjIwiLZvAdvWcUywhX7SwTDlzNtD3WghqwoEDO9IYiTVFLZWLcP4a
XU0uQxLnRPVtnq3jURGMwkpctvpdb9xRUgiDLup5jCha2i7LdYrtqZs73sMkLvtmrOxfgwkbs8tm
qw4o95uEMqzWnNy15nNjgzNd/ou6nWTC9KS5Y/XzRW3V4TBinAHaZSTlg+0i0ZcL4VHEVsO/BIgy
qPy48iBx8lWIZPExSDCC8yPjoMXKv8wgb5WyAUcaENdLbb4yrNp/Yj0OjEU21x4f4qD0DAK9pcFP
1dfrSLJUVCYBKdln+ZQxgFSkBq2DL/bE4Kgw0TqIWVyF8Pv9LVmCl3hS45n6uBlOyUHprGMYkj1C
b2tTmDT5zmZbwn3P441v/yclNZATGap8hetrmXVMxZe9A2WGymsXDJenkMdzVx14WPSz9CDdN/sh
sF2Ng2duutfsCNiKS7eXW1df35zFQQElggFjHreBZu1B2v7apQglrtD1PgxErvmxZwIur5X6TFA+
jZ0iE+oWyTCZw60pQRkuFsH0tmaJ0FE3V4OYA6FofG52sfCjfYIUfC7DqjFyAzSp2ni3JvvZj6A+
79xAlcnj9yQNoXgAWHOnSA/kOQ6IlN5gOIUUvQJYS0v6BAN2qDQHLJIjbeL55r1lSb+z8tHxglai
KFeKRHx3/QqMxMZbgpvJ6G9WT8BI5fXNY1ZncyiDmSbIwHlsIGb9mP4ggYMYHYWO1Bnc4LqGvXNJ
h0xnoqzhj3IwI3CzWB5nmKPkYDoKgZK8YEsxn6pqEfJ31ThN3yVDqdpTAe8DesgtMWMjq9fQh0CR
2m+SlfeeK6HIj3XZTm8fE+0t+/CsblN3niyTnDFlyJNga8s/XW0ieFGIxDtFQNFkQFzwfkrY/JHU
FjqDPuVT/dTg3EGrudkp90V1OEw0GaYqGOooeyWtvzzTkvxaauPx46cSdvp8wH5Z2s3hud6k9n55
Z9vOX/hvm4kZp5bIbI5ho1LNd6WuJXhs52Bsougp200Z45dhqYvTvwSCv3qooMDnuKruqyfrvaGx
A/aS042zXpF59sEZ3sKPLR4L33wVVwawCeCmJvV9GTvMjoOXOx/Anoghg8pnTAivmAYUcvFhCNdi
gW7M4ba1F1tGkudW21JcWhWBm1x8nlze/oa+Gc+gDvzp7aGgbrhGP/yn/mHxCWAJRkYeubz24d5P
yud/oRjJF9RxVZxSBxPItnCgHdSmoEOlvlMjIYX4Wh+P4r6ctyPMuiNrwYTPBp5mAPqiTzOD3pw9
Hez9zjX5W+v2e+u6OhtTQKPZeAx4Zm2urkiF1I6LKAhS9107N1Nq7+rJ66h+RrR6MCqJbu+ztjJG
VECVB8xIo90Qq6Hbdb5Utk42RNuV0ZnfTBcR+M0+YIQUxOYI7D22ZQw4u7Ywo+I+cGz793a6yI3b
qckR8YlWuaM+da6MHL5oPhJkVFouQq0CodZ6QZi+T5P94sGLEBcDKMFBx5Tcs+MI+dnJ7lQuFlfa
1xTsa9RHNP7gncyrkrjqxFDev/eE8jPpJQXRoV6qWiOpCR11aMyn5+iLbwyapx4XHiZr5FL4/NEm
IMTq4Is0mxbo2+12/ZZePN80W0DFDdOIindA0pwH1qrrqq2JboZEoYldWbjisjRbXnWQjJzYxMSm
eAlz76QRI7BzLe/pEBukKtusXj7iedDsg6HD0Vc8Hmstm6bGKFxsu0JeHSEuEC+pr8c2DrrSbbaq
pPmug3gc0iJnFHf3vDTsDm/+4+eRiJ2cY51U0DsrDEzlkOQBfpgilWr7UZ/g9iDEMbEy9NZWf0wt
P4/r+GKh0U30umAaMuQ3u0SRm4h7seeNxIugS2eDRltiWX/6zNGEQ6opm3NKHxQVm9MKUesvpFR+
C93vJolJCDC8MsqKOJe1eGBmad+u0rMr87VQyOOOzniiHZLpxqOO1GCBzQfqg/nEnREVcM0BGFnx
tDvvGzttz4sDMLzwoWgt/f/XgLtwpc4wIFSnxRsiFwl21qtskkiKFF0n5cIqaK2lsy86X96L9YwA
ELig+RIZPbjBhIAVfQUGslJYNZ6KErrlPp98ECk0poTNnGUFflmjs4EKm+/EP9kZR5Nmbe86U4qv
eYGBIO4/3NECKN+J1rmgp9qkkg4Cw2S6hTDwgBUlcBRZQKLaLVTcFWRaAXIryK4ylgliVwC5XDxx
V6kyBEMMpohVY3bV9uUI/Zhe9ECiN9WgAVCchmiVHmKDn/gRp00n1h9yt7A61N3LtMtHIrdryQB8
Vxyfk23jOLluYMKbUPnHdkRoviaW0qfeE5So5fxdBu4s6qDm3/c871MNpvdz4yY+PBkELedrdrFG
qdELi5m+Sc6JiW4t4b9Ec9QETCZrMakna2nGx8lotuqeEuO7LYexYTFmP7oPsJ9Ba3IGbopqiADk
oNS9NG5vOGLD5xGHmn8TfefnxLmWFcrc5KoZvA3ea1Fg5O2AnEReMOy36ACUMVHV9TUsMl2y0yyt
YhtZBS37agCSTCCOjraEeFpf0VOvfcPpidx/MI/Nn70wj8vfOcnNzzfKwq6DrlOpc3a2DSiEGTvO
EQFGNuPgNaD4oOJfSArcir3rqI92YwOM3UNO03m3WZGZfDcdGFK4z6z2N18BAm4klZdpys4PUAcM
NDPARyV70yAXoct/CmjEJuLlK30P8IHUwIeOdCNYC0LQ2soRu0bY9BnjLd13e+8eI0P594hCWX0j
bONaj707Ylq9TB6OS9nv+yi2QRj7Bw/QUGMUxo2OyZ8KS8c29hUGSM4pTmzTfOLPMFGEImcpi01G
kiRUKN3jPCfPyut+Xd12CYV3kcVzr62S6nfWPsbSVUcRjpbUsTSmawNoVkh8V+tge6Y655+ZoSTQ
Ey2BlCZ9SvHPEuuYSjqSR1ZKHRaZ6t6akv1Q181FhL8fG2q0mZYmhzJgnEvPpO+/8XqYQDCD9N1a
hZAlqh6RVMVFFXzQulJKisV5zFNLpIb0Z9foKJVjm/GjAJbWgMLwkfcRI0vamS3ecaLPmAIHHvpA
6Q19jjPmj6sJ7k0XeT1cKi2xsJai+aPpY4qKnG339RMrXt001D7V6dscBhfdUT3yQyvtxHpXrylN
9I73NQDR9cFO31y6Nt17YkDfWqUc+sNIZ3SUFnrVNBXhXoNLe4Jh7xRMWSv6Aj3Jn9f8fLwIgpI8
uCrwPlSws6IDp5n4KxDxBKEemcEdSVUSuuhWMMAOiJ9Xw0//5zbQLQzfMhP35XuTUbxPmT6MS8Qx
huWFqF52cljDUCo8uMX+/Y4lJ6/EqCSaMxrebhmyE/XoCX4YuVDdOZcN7UdnFmO7AVqW00adWl+P
0/kUYysxJhVuGCiDytCK0Hsjdak18spmSD2pP0WnZbIKQIEoA9etrU75iiVE9AD6Q24aGGKcy5e0
xH1ProEXU+KyQd5zUdN2fH1l8EFuluS4ge6avEJ+/wJkJAjVdB6Geen0PDJp5Anhsb/5G8oqN2QB
XGoyXh0b9Piv1THzY5/S/xg2hlpinabXEf2qJ4oONK6TCIV7iLgqnZnHuVQ/SNI4jD0m8VCJIrCd
Bfz6Awa87CCcIp9Lz8TL0o9C0w3Wimh365wEYiC0dYCdiWFbcr3HcMXXJ9gnpupYl4AmcRiI5vrX
99hhMwGLZVcmGmVv2sbA2o07cob+QEq+zaORcCxy8NA0yBekHnYobAwTzNMwTL/ANdYhZAGnIMF6
e5z/NcGh/NK5yuz51SU3DBVdkwc0DlgK6ivTUlVO9qn1JSErUv6GaM0YFbPP4Y7Muk5NpkeWY6dZ
g8iEVYlSdPT4TpwgDFw+QORouSOSBZEguz/6esBMTNmmoRtbu2QFh4lDm1A0o/w5fvU6yx2qvmrE
+hCDCZ3sPUrM+xDot5X3jYLVWadJXC1BRNZdliUJkpjb8aYeelFTEI84n/ChiAPkvRobZykED86s
9b0rAHdqmwTBXLrImpmphinsW+uJJZCFecYCczvqykvLWDo7wAfAEjMuw98yoo4XGjJJNlNVEeA4
9GC8SXKYqT0ZWCqgJneHLWSBOzYdiyePoeQqHRqu/EXzVmMSwS0PXlILjlazMVfHGLcO/Eiw55HP
uS2PXRplV6IlH4qm5BpTbSC+MhL1e9ESZ78okdqrb5fJd5XQBw5pFX3lLZG9CsraQaVaQpkHW1/9
VYdNy4AOCrGaNA9K1qlqwbWGXaJku+mPZ8VCHOXZdRY/iba4STNtQRHHfZmV0xaA/rT8wUzdT0Ks
GdQDkaZ8sq8GrCn0bAHwJIyrbnpQ1AAJp1WG7U/Jn0JrCd6Ml+z+rUPV3ysQoIkaE8PeGgVZv/jn
qq6YJSwUam+LaT4BaRv7jQyNNfMN/c2RZSjDgb4GP/I8UOPkMssENGjDqm9oVvVwm/slljcWt0YL
FG9Pe5cLd9UdPzoZl980Seic6ikR3mabmWihwJ7c5yrM8LTQFAXcqs2G0WIlA08UUSyZWQBsv3Rh
w9CwRj7Ld+8dRxFH2tx3//5CHa7GuERqThq1KL3P9Aff9XL5wFwr8wMwJRStKvdv7Z+TwYqlUd0J
7eh/h3K1CylVuRm8vj9rDgosisxaTMmSeu10fYQUuphxHUXF+MtsgoJ5RCjp2/wloBO5nhhm0Okb
wgYp0zUjucrqXfbbmKLbDI5V++efcWC61QObxkkaGXDs1tAuiaVSDwrx9Dao/q8Lu7wqrw7yAcYe
bWC3fzYeqRq5UeJMZp6+kIErXJFJWtisA7TlFBMRQdFPgtTs3fPzM6qhADO72LgKJLqN8GQLcVnc
ph5vEj54lZ6BFYLFrMDmnt0NFChWvF6ES8OOTjBUQMYJ/ILEBGYSY2Y6vENux6V4WrDSZuuAMxLd
YoRUEFlH9kfQbcNtojhcz8X85NsZZrNP5wW67Xy9LmtS3roQF2qD2zz+ZBpAzp4QmPdUr8M83V/Q
wKYpr44HC8jKyHguPX2mftP9zHfY9eIu8ZrCtBgBKQccFNxtgZu1IvXEo4KXipOhjffTUaboJhOm
R0APwZ+IhZoNia39TxQVNhnGfyvX4qQ/O1z59dMwhW2qz3E5cf/qJL+ADYru6DPdBdWeNocKoGQ0
CfEQoY1/g81mTtVqGZSFxVeIuSf99MWjNqBcvCfmM/aP0ArpzkJcFv2YF0Zk+VvI4GbzxLPV7hwP
q4+bGrO6IpRlBYIWKllJp/pP8obSC/EqDPT7l4puvzeAZNfqt4eBcUkMPm4REFjo8GjrUbJZ+skO
r0FiRuTeGls02dWVF3gOi0ZoS/h5Bv2axZWUNRzl1uIiTu9fovAkHWkJPFtb5LjDgDK3SuG675DQ
FG/Mm3soqv2iNAQLYxf7DePsZl5SUddJhNl3BzTxyrFEwbLZx4BIKw6LDAcyK8VDjjYV2gVZNswc
FFjNsGkGKT2iQ4IqfGwoiqsRZYnfUSgpIT72d+0mdWhi6xEHfLEShyjO9Hpspqm67rZHFYZrMuzg
uBvZLDWHe1F5IYXzYylAhpLlkf2ANrhYQui9VJ1QWWUQJMGAe7CjH2WllY11zqPPkLMTnZQGbyT3
Ag8QKIUJfaI0qRq+74IR/G5eweiXJwcX3zBnGSauIRvcm3E7pWYGqFiM5Ptyb9GwVcWhbFDnWcT0
kqLFkxWUjv3v41cuPTVacvP83qHJ/unxyJ3g7+BaQcUV4NrlYhXkOfTd+snhg2G29JRjt4cIsaCJ
55G9YH211A8Mq7h4hmZkSOmna5oOV7yr6MgxBMSsD4j5x+M2Qfu4P4wCF9311E6tNbQTqiFWlFkY
UHPFB5PCojsB+HnUVQzMTRSkqYcJAxYabZ0UnGD1DsF2OQcHqEmR609XPoXBZeJYQK7u1wdBivZe
LNNfObXw2tH8dugHFOCPTiYP3FPrV8uU7gqfdoaFLbPFuY9gKJ384wyt9SYctZZT0/+14aLZXp5k
2vhC17rOJLPOd7SXvrojjJIACDqXTapUEjdzn0CG4h5MDgiNmXI00uJwkbZGpOsrMV78jPxLHAK6
2SnUn2kPx8qTUmEB5MVsugKnJJN4mcvhYGtj0PZ+K9YECVHfjWIzEBGRqRptChYOjpwrr/8UR5nP
mrIKtNbk4c3CjKDPTOApjk4VoHGrIsTyoVtID3V1lCV10Gg//Ip0XA03HIMY7e3mnuhqUUoOj5fO
vuoL6HDkCMwKXlfHgaXgLL8ve+puuRK8CQsxX9ci6k0W+WY9LE0zEOB/ZElQm/50dtnv1MihY/qA
BGCly/Qimm8/eeiPoG8Wv6UShu9EQYCdUN4cdhWAsWes1/xNbERnFwkbAad0C+6ttWrMTKYAaIPo
DO1XISPM0rC+Pd/bJNsBS3tHKzlYfzoROjLki1j8gTUHdEO7/U+3eIpeOeXBsR21+zAIFxtsH86I
+mqv5f3PS5xLYsaY7kMZg948cLIHE53P97Ni6Bl/3vruJ+bOWCZjYyNXUYjhGSXGC5upZ+fvHYPS
Q3S2LjqzLN7HJLdPkfZoXTtQnk9zqiS85MRhz79HNIiPJRVLpWaw8HH7PhNOXFqUx3WP9Ls+1tIn
EHCUfAMWgAkXoX+R3ucJWvyUuwD407iaB6TqWxrdd4QBMLljR83k8XECnAgIkgz8DhSe+vePfkBn
4qMDZ3FA+1DyQ2jBH8oaKsgNwGOgyMKDAGBwrkfkio1M6/LSmTVaMlyhsf4dhztTKoPCIsxJ5Slr
toMA0ovMHBypfMheU26+OGtu8xevmBjEAzxQcGXggtHkFYhAolOavpt+nUSjzwgVvZc9P209sfmi
WrqnA/J1+F3q/EWNgT+53nzvznMI+B9kbSY4x2cetePf8SocosvlNhF9HpyZewGYJ+h2ezx8Yswh
XeH6KKCsDgnOL6QNU3VJNS6hkOO2DrE76aG5uzEoj0VG4ckEWh+qLd/q/fWHuZjcLqr9a0xgfkeU
mdQtH0yJwu8AGz018TzkxTqu/P70TVfwhjjRUZIom6WeQpXHpeDSBP1bRswHCO1FHCmRqyqVJ19q
EbDkDRyp8iX1W9gBgUYi0mUlFTdnQBTUqjGy+XzKKyLjiD6IV42AqdKYWyvmJPMgzueBRfZBV6SA
HYzbAaasdFs/sEKKw2BAEe9OsAWzK6Y3B+3SlTY3kjlRoGDDbQZs9rRGjDHIH+eEax6dEnHZaI40
i/VuVDnEWpMSTwjecYMld0bZypz36NFDmfAVfPID4b3y6TeNpDaF5bZGdWm+mM1pVfMVWsWO1Y5P
IMdLVqATq4WCmto5W5W63qwjFe55o8S8xbhWuSVh5nDZKwZ0fKQkzYP6Q0q6+nD+4Yu3/ZQlIX/b
+eODNZ5LeoWZiBklww2+pQdvF091LzOdiZFJnp4wt6OV2mmxY33rde2tSBHahCJg/WlmOlnuK+yn
SkALDLxeHMQIo/VvswQ+EApcpQNYMrQhhYg7cb5cSMHiT+XqCYF96lDGbFNfN73cePpLDqVy+c5q
moIye8h3nDu8ESQF2eOIdHwaHyjeGEZNAH18gzYtxW/85wXMwCi8ElDmWHbxQQa4ypGNtcbg6lC5
Rwdv1LcD4OwdS+gaDDL2zNPpjgfIEQRUp8VUMBOh04DuHETBI/NO4xmXfXCJ9HZbHRZD93NPkLXN
58clHPDk8IzpGD9MgdBtwYzENTbKOmVV4M8Y+USyqhABnHFPfZtGZuxy91tskQUitMvW/TRncgv7
AJ9uob0CbTFzrKikuwtuM4uBcEY21DtSx0SjhskmUDctCXPs1+4csqiFCqL4pQkr6/ePb0BHOa/d
d+LZhxsjXMzzCnZCQ91uH468pZxJ9XLDYgNn5No9UJyN2sgMfA6/1oMwpG5uOc7mJMXGFVj24cHg
aDmK20HUdEX7QvbCNh/7DKFgnKA0qatbQrm0y9h/EjYgc4ofJkiXZvSnKA+QsXZLpcw5qQ976UUr
VWh7UdadBX8v6ZvDaW+z3tAgb3OziMpPvaS5WNi4LeFYcFLADwZ9gZAT88Kb1USSxd/caH3ZyCe3
LuWsQHvAw7MTiadcOZxot+eYKiiu7wiRq65SetxsvmTNC6x5ioq2pkiApb7LsveTEgLf6R/pFsym
JRESqSs62cfV1tAjiuNLfLXZsHzQBtnnYUKTk1mj+E8N6MQHH9m0i+UNxjKnpifm7nE6bFhNICVC
TrQx+p6T156tL+mxwxACTbqX2EKvRvxcfJjQgpsp37wikkD/1cdFPBPid7l6y/jnpQ61hlYVrzkt
W3If0LUHutFxTR6u7EoIs3vzfTNgG7B3x9a9s4DBEPnsgW+e7QJDmTlHGQ1QOS0+3pm64ifjAIDS
qkhu9iPEMkh9qG5N23psHj/zNIpSEABS2f68kUJDdyOmKRAWgoQf4KK1igg7/GbuGemXGTVbIgjt
NgB61P+rvV+JjbtMluJzrkRRUC2GDnBSRgV6gSE5G7NoxkA82QqB/4dcjoJcL9fwMZYUbJ9Zp9LZ
iHp/hjiBv391i8vHfjxY1RAp0TcIE19FPZFtbVcObZhq9Rf9XUOUF+PG9oVM/uVcvUZN0Us+dKM4
freov+iB7I/prsWIV7b+q2GuCpnfB36V9XsixsfW30cR+OhwVNwRie0hRiojm/nwUIjn6YJ37G4l
nml4TVEiIEJwKBwBgXzV0vvyA2SGOaL3ZC3jXumH37xikrGjzWi2c/EXRMQLdEYpgm23W1nyUHvk
pjVXipN+BSmN31uYrjFBmO6TJU499bqiPxjZ4oj3BMK95s9w3cKkpB98lV+/OSXjXd7SCLSMJi4O
WcCiVhec/5LdR4tuuJklEUZZX3TED9ElFPzcy++VLur9MwHUH1LRGm7kVfjRmke5JCIDO9s4JYZt
cvlk2D9Ou5/yoSSVxmJkPtPBuo9C1iNEckOLy15a7ICyZGoYIaM43NgcCUKl4Y7Y84OL4kUOxe5+
ay/ebbLDHojdn9LJhXfH4a3GGBUQ6COl9N7XwhaHRhHsS6jTCuxI1unVowTXaeJqUvo0pKMJphVN
a41oZ+iGWJ6UHh7+VMm4upt/6T6/SsSUqAOBHqNw9E+vnLBjWMRc8hL0JNhMgBq5VTLn9bKVdI3V
IeUpd0Dgtk/b75x0pxZaYNcgV0GbG3AStrXT8RxVjeZuZfFRLR6ipT0/z60MBjIBaK62y3Q1PmMP
w5cQ8qTNDT1NfteiJUtjTYBpalRvif3Yasbe3wmxocB97eTBIJeRneMhGqRLi8lfmVU49bJQV4cG
2aDyrdLKTM0ybp+n8NMt0GenU2tw3mF3bgvpjM8RQHEkOb5OHmY/vhxLPgJS+CqmIHngXcvpfKDm
SW5GzxBcYZSvQh/qQZ9nyThu24D5qz4ALb5SVexeu6AbDL7dUDkdhLk8aMy/Cl5DXfDI8qWf54vP
6qlrTTSyUZGdsBkmhXxTc2FQ5CGUyhRTenZkEiBlRsuGfhf41J5fk0Z3nDJ234itRwhunV8DZztT
DopSKvxDRQTkjON56xuh1+w6L4bKt3eN5m2fIgDa2u44RP17C5CpLyTiyzYnGbr8BdEa/LinPxNa
V0MpjKI/JooXyHs8v37iMcT0VSHp7QxUsR+JXFs/Mk/WoCyhicjoyVHzVVLmrx4P6H/N+V1FoPT3
YteYlld7kf48GvU1OmVrkozHFrEQkNcN/nDi7JeVZEMFfXElXv+AflmibLdVHUqdMkrACSd8eCLO
PTsaofy6N7fMravIKwAkQowZoG19ivGfSG/kQKQo/fH6PozcakzMRTPkJM2Yzwz4A25Sf7/582OM
SnUgHpDAacgbirZC9eAG0uj5c2PhkoFIafJ7S6FdUGkSjolsZkvhN7+ICzk31MfKV1CQec0Zus6s
VGVohW1ZRA2pP4ydEoC6s63skUrS5SFf4OL5TVsRkS5TVbZqPiOK6cPVikHN0fI8bOX1eYAPw8ke
panHHaN0FrIdShHtA6VPMLSKgv9SSnYMLTzOQog+A8RLJ15jRJ7QTMIa//giAzRnc2K+0X3CiP1Q
Yxlea5W4SsqbySmM14MvngrHRwZaBdM5CY2FAVZnVCQ7HivNohU2t01eele9SLVO8sU+YtsoJidm
MsnObhH6qysASp5TuhQD2mFD+6Jdrb04vseq3MS/eaFejxGFeUMguxoRXUWp3UOHtWAE6+qyNXcc
CRjsYMsNwXJ5ST2vsUZGe/mPZkCBunG7fwqyk9pTcL0vgZcEvpT1ZlQz56+LjKaxfbwObqvBrVPJ
iheKst5nM6UbPh81NYdJrQuSwSgraqJUftcEn8N1CBtVPjLpt75VK7CaBL7LgmwlLPZVjJuJSihw
zhbXQqXhXwRj24VqDJEL5vF3yz26LLn3sDuSPhZWQq9T1ZDO8Jg8VDB1Rg0Gzm6GVQSRx4m/o9J1
gO0Vq+Z7xPNZs9QrJv2LRZtPoY+cN6EffRbjJkuWdD2IHQAhWvph/tqgI8TihT1DDnkSo2Mbf9hj
9JOxBfYX5lbnd7/XauW0FDHlrPvQbEoS8PCcdx6+M9pkDk/Tidh/WasArK0Z4ft0pD6vJOSzBvy+
Xh8r9e+lDnCYQNKa08xxXommfW02SuZZrWmpmd/N22NFFIrVB4VSyLUHt3Vk8Y5UKQ9we1FmmM/n
uVlctkgNEmzy/cE50o/iVGqv3kKIrO0Bu1zLXmrYab36/YGa0AuC+GSOhpZaDLC81tamHwAINR0O
pe2zbW+5ZKIpd0l1qwkBTRwVygF2VCqVVmNr5v/G1harnypDS0DrQKntQY5YFd4+gMPcnRNB6Jjy
dlwfJjnb0PcZ+NreFB2KGy9JlNepejQv1tZfofBm7H+kekMTks90oi20h8lpYvqUzdNWK5seDJbC
P5QO/j3SA0/WmhR0EWv1NQgBedo7TMjxaF+GBbQMAN7Sc+0r0EIah72f+F33dF/N/0vC9D1GK/lq
NkKyyklVeac6kSkrBj3N21GPev3hBgx+oZ9bn+z2YDJFInavh27/SfkYWj2QLaaT/volXvnaEC5b
lLtF0dnw1sF4zf8+gE/Hq+N4zWEPIN6auFCuWUZb4VnEsV5u6VSagGJ1qIZAzZ5+VwVmNrXNrKjN
MRM0z/GLk3cc7QZIdKuKHEh8dPhWkudBChBuLDp9v4AHPWXY3brdsfonAmwJiuMiUrjalrqKBZSF
Ft3S4UqmxRYgu2VuKHEBlKtZzNVk6vo38vmV7OnaFmA95WsprqHEEYaDfXHA3WM7IJkeoUnoJU9b
J7aMv8RZ1wbmiNbpqYxVHInH3Y6PYvv/PdJphBxRmatAyEylog5F86GIGdjPLSLJSSOCVhv7/Ycu
C0r4QjrqdW2FrWAXB2CkMvCgdPZKLDEiKPZMWhvVyvSPWbF9pY8GkPC4RivOuhYGe/UChShsX0OU
pzD8qnEzh/ZpRtYRfRk4QJYnzuh7FlWKLg3sqkZRG0iomQ3tzgbRHmwI9LeXwfWFVq9R7Dh0qk87
6BlXi7pCUK7YVaujtTYFROYTSGzobEj1r0OZTos866L2qAD/DxItdHHVhhPLKtP37iYXomU8rzTb
PPup7LfHdZ54ptt7sLJUFBx9ZNiXf/jRV82rfBR5ZnD7Gp5W+UuIJt/PRsdp1UqUtM4Uc1aYNSCE
sPTBZ+0jXHGd+gGoq+Q3WtkxaHFvFDShLIe6YOqXp3bYh+DjdXdAwsbDVjBGgGjstjFFFxDmdIFV
JY1ZBg+D9SgnkR+5xtG3wGJWGdqhPdJsbTizc0p4NGpzTmuMk5+RG/4zEQbVzw7y7KBLyHzJ4B2e
KQWcRVIAAWBFzNkCREq4bt5r0gqex8awNgu9EBpnyyAnjf1wwy97exLJMABiSs5rCtEZwwSThq3A
+HEYEnAe8yFxSFChkD3BcYaMqVHVgwrgxyZBx9po82xGL52xuMWKbjOe9SWKn5XedA90gv2uTPgh
1km2gf/1Wv0Da6A5sRdhzt1x1vevJ6HFEndG0/XsGw078QQnrLhG1752Lp+GQhqPSx206yuMCjfv
RjpbMKGsC6cv+RGnbcymRMb82lN7WEn3DdIm4I6WXLaS/RvUY24277MzJnHGq6srCZ5QbXJInCTy
1uKj1iAT/R7xNVsWoWjqC9uq7c6OvbLTtgMLvVVU/anXB5zu00Ip/wcluI3omPA7YDrV3VHjjw/A
RVMgrx69wKsrDRZPlc4ATspQDY2qQV3W46t3KeU0FYN00JueS6fwsgfosD8oeDHQgYhRXNi5XjQI
a3P9IettpWLvCu4PFvBznWbg5qsfFxqIz/FHH7bwOdasP9FFmKusxlpbLuuEvvDCaEhpHdG30tqW
XFym3A9APErrz8Xjn+nQN793+jR6xJ/Dr1wpn/v/iGWp5uMvG8aNXqA5QesrLzXkPgZQ6DzLzxhf
aEJEL7tB0iYsVePYNN6I8MK/BokSrQ8QYQQTjEX5ppwCqgNTBowdgeA1HS3e5DzZ6tZxXr/HUj8T
QTm5XGEBlZsLXDeRf+eIHC7pIYZ+RsCSamFvBD4+W49tJB4Qqc8DIOy0Cad5S4KZOUbXdfNpD3xv
FDz+D6Rq50SRpp53GCJQ7R+hIcdlPYYl2ImjGaEwylbgGcjXOWSIuIcNYrRJ8YGydxzXfLl9+JWi
KQPXQrqkSaW7bvSIKgv/u4vmmQX5tjJrJafgmGYznWoDaEEFNBwC/fx3hC3Lu4D9nibsSeBlCT99
QeszF/MBek8IpC6e+RRJkA3lNscqFcgoVpOypigRKyL0zVSU2Q7HYHeG0U2JljHnuBHtiqAjfhBz
VtzMAEa5oiYi6x3PJG0Mu3XVCGWM6SeGVATrwAnZR3IdGi+4ngAcVcL9SoEKeoWKhh8xtZIUaEKn
NLv20l0TXdAFmNMInoicZLEo1vWAtMEwIGNY6OHecPZYRR38Hn+rpnu/vOCKjYsR/zy6auqenKxe
GaI8r0rGUp1pB1ukOrP+MnGNf994VU6hsKF+cr/8glkskloNFtbEGJpVNhXuuf7QLx0aecAZVfL8
odBni80UtVGLzOt9SKTNB2gbNNrlRGWWhmbbeVtMaQFsQvmLVsM047hbB01qNPsxPTsaDU7K0WQs
0WkZdnhA0rIXkRsyP+65lpykM4Y8FURnfdFYdQpdRhN2nLP2GeSIEtI06ugOtuJ8++B8iRMf7kgO
wuZ++dQ8KW54uBi1Q9zOZ2YcnV+53CFxH+Gu8x1/R3Q2UzcUiVjfe9GMs3XYzJrNskFm2V5rMRq4
cncq/wTPU2hhHTuGvcl1D9h0NdWDaYjCCxu1L6RnGQKJVtf0to18Ff3gPWqnHfQLR9h/9PoNQ5Gp
VooF12WZ23hkp1I4CZ/i6R7l2tTr3f2nMVGyFbMOXTZCDjRhsqQ5vDgnnJ8hhKkb8kBFnGPnwkkm
gZbZjrL0KK2PYwQMbUw244AphIX3gRAjHzOcuD47212F9/VGSFXPjxL79Q78Jv5PUGjkvHn4rO7j
wDm6gmzrTqlTMG7JCQMKnQfLjMboD6m1SDKX2zFyD3MgkkXEMQbqDQWsg/LKkgMYDEE4D0raFvLt
UxCzHeqBp5BuZ+I9ZV/O8jTwFzrJw3GDNfOC0luIkc8EoeoMwnfsIo1wS3KVsxyg6nr5NT1RUvFL
a/6Uj+342N1t3LRSvhFI2uRhPYEqOVTAtgc0JLT1NfWh3CYPvMVq8cxUQCTkoELjk2Z6Rl2Io17W
N855kp3D/FLpv4DIQD92FKdnneSInpbYG5xoZa4jedkb1x0cS9m9W+Sxq0ID+/Y85l57eUcuiNA6
Da9Y+LnQd4YYLID/yZYWDSJS347bBcNyWR5/MB6BdPN3VTev1KNyyubPBx3df6Ky4CdKDsBwK7dQ
ahsesBbEhGpNxtRLOZLwvIpebAVd8ycmkB8lXXmkNOpS6itZSxK4K4/JIEGYdqGgZxYtDjV0T/Ak
Iz1pfE3OJ1uTJUyAL+1rL1eJcIvF+yKgKZYeqpHJlo51WNbi+TflSakIMtHGL5+HyG3d3uOqEoEJ
Aqgnzrb6EyD8yuA3SylwUxrH1R/YCmW7gDACjtF++23ETaSR9NxC6tRpwuXhuaKeZYoBkP05qHXM
A9TuKxEszh3Cn/9xMbl1Ktghg9k2Lhkh/ZRdy2v5Z+qvW6u+w8P0ICbaiq0RkxKo4933p+T6Lq7y
nL8MkguuD5WA/VBJk10tRgz26u3QsJ6dCgVvBZlZw7vdo+gT99x7p33SnhZg7u3LKQPFWFeYZl9j
4L/5PgFrv2+Rrr6lzUhOvJw0p1dgMtGood1rqdrYcStmciBo28wUJpKj6rpdpQvVGyNBf5m1s8Pt
D/HLwqcMH7ejfZru/PuzlmIRDZBoR5/djPq+E/srJyXLpd3FwBjIluarGNSzb563STenkuOfaaPL
nAh6xbFpaCDSSLuv03bLJn2yYJtsFAeynFuBPgNgaKrCqnqZtQ5NRZ+h7BTZZDFORr0fw0mtmvjs
u8FEYqy3BYim6SoGlo2YWTHIPF5f4JKpHKcT6SChWITz6U0tPJ70qBh5FL6HuX7JcVwav2rBkXfn
K+zqldlrgAIW8F1h7W8G55BA7B9bfPsc3gebS/G5Uhb7tuHEMksYM9dzp7uafWQ6s5zn8BMrRewn
ftaj1RNuyJlhFyft8fv87NfbObO6J2+kb+LdZ3dU2JEvGsvf/23a3j34FlXzeyjIn8S1uRuKXonL
U++Z2X+afSHsJaWqf3UaWswHKGq/U+HqK9yBXJuF3qCGuFprtpEFdFgLG0qJp658WEgO1/TuFJal
UhH2FefJ9DJbzYgTiLZx8tHK94dSqWqpCB/bRATwCf+I4QjEivvWPA5Ac+GhGdx7pVksDpvlJLBv
WlkNBsnlfdTsC16UYB+frtF0OC9+9akYzP8MKJN4EXYx5wZWeB/hOBl+kk6PSYGrHCISm0X8d284
MDbxiB6I0EcH0FBhfFhYFbhYttp+bzEAivkCdaIgaRqN+la/5t2/X1Y84WqD2+H0SqzPBbsS24bU
I+8lCxAe9TvjQ/mStzdVALuqDs1cOo+XHJVDEB9WJDehrfCn3AYwkTmYa97pfEG3M/SQyJOrsh+C
tGtnGUBAMRxzuUHVEUyZd4TouGHkq5OL21MBHScpzH8LizRLftQ/Co1JNBEjCHicQp0s0oNwpslh
ULUNZDXiHaP2SDXpsd/851rwdhdCff4sA43JTiuKpqG9Rq5rkmdZu2GmsK4Anpugxd+6keDxHyJv
SoNXfDLclJDMGDfGnWcW8efYcMKrjutY3Dsj0xWdD7o6fdp3OfpH/n4xu5pIfODBXECU5PAEcpjU
Sqi8kf5aXFcCNzzl0yDw6tes2iYP9FzL4Gi0ceFscRVegLHTSSgqv85NbfpJwP+2SM3j8xEECJ6w
pfK63L7E4R2PGQsVwmfpgVb/sCiUIuhIu8M30Z5O5ptzLtlPycL3rjxzgyB0jSeuKC/qcO3AmeV8
ejAC6BIPGXRULnAiIpImRBeRIB4orU5AVtHLCMJ0f/+SdN0SJ14su8N37qnTAHV+aIW9eZRAp4oq
TOJUDFcHZk9LwqOqOx79UmKdiqD5pfgS8kkR1OwOVrxd4ATHXrLdRDaoCso1pFixwSdOO213+sFg
B7IzLEpllZ/dsR3M4qQxGWa5mvdL1Lv89EPTx5BE7pYmK+KcGh0uu7FYqM0+koZtvlUS4th4nzK7
bxX+WzzJj1yxMCpOFrdFaxjkDxOMmyixyFwcqa6pYl+nxNlYkbBlTHwrm6D9E7NQHBvR4/UNkfR+
4FeR6tfTnbNoJmPw18joBl6ODhHq9i3kB9I9B1OeS9iF8v/Rl8SXFg/8s+iRaUw2aEfXuSESf2bM
+HXxoPJ6zDGZiRCyZ7MRoUlOYYEIb3kv2YZj+SfK+Jhy3y3V2yYw4Z3fHWLHHxh2RW65aZ+NIaOB
xLWL9IEfJo9mDDV3ShdY16DeBYquR6pkuaITvEHwM9+i6i1Dqaf8ZfvBXBhsDLB2ZOBvlBmuEv3t
CdYDUQJHvsWoVYr6rCgUYSP7HxiIEbc9Ce6qW2Ueu8B8AFTK3Y3vUdMKsmXU9cp3jU5jpuiyX9UK
x/h+gkDJ+xnK50zuFprgEW4QjOYlIH/pIWdiSAHeTxa9XdMJ/gLTGma9s3+8hVC0QyqtEESiMZ7P
NeKDFYl5QKDDNzInb2VDihIfMEC7UhejePTXHdpv9HX1SDCAiPZiTx309X+2SmKonn8jcI7cyCs2
imkPlbhiPADfgmJCr6Vmr4gfrtOl0fmNIFL3yDyfXp/VZwtldg1RWfX8MBlsypgq+2pJZVu8k8Nw
CFRC5lwT5TaD0wFgA7Q4OhO0OMAtsRvrWxPWz2pSnXMyD2LjXvxQHg9umXhW7JSQFN80waZRWttM
eSdL8AvmhLbw5CN3RcUTNyA3n8EMRsp5YGdQhN6/DhH8VQHMUYfNhQNnwwVeGPtTt91MviLrkR/t
YBcnU+0fkuKu62HHMd3tyckXszy6AfLCA57p9hCGFZjOyaSHondcnY1KJqyP5HjRPP0mOREO3ug5
HSpsNkPZM2QXbT6ztxANS10t5ZwKKEHefjQv/BI/oFamOxmHrhasXqjDX1PjAxb+xx/x1u0Ww/Jq
F+qFp7MX5uyTnme8ky1TkvtcgTC+1KAPmgXTSwvv0JBbUgR0rmZkl6zWKfA/MsMEN9+yfGCBfZB1
MuY8TuU1FVgV12VmYFKOGmrZKi++AcipxfS70k78GJz2gKk56B+NuclRnmCcEkfo9rh/EJJ8TdRD
NJPqwL/xAfgo2JfGmvGJ5RVmL46TJtTwxRvCK28kHne6J2l5RakAj95eeCQyuVBPpeLb49GRODLd
3cadkrXJhIweRmEgjRxWHx8pSgLsLkBhWOjJTK3vqp+Wu7oMWWA2pCbcCwGAptV7mKwnvY6Dx6wt
XQgTvBOSGXNB6Hk74FLTMQmprZMxLkCh7s/ZxxaKjBrIESUT3O1s+ba5aTT08jyH7mKzjM5PmsM2
/9njac0TMXyhuVCb6pBrnb9NCTFWjGOekSTLiW4KWDwfa+tMeEwWJdwha5MQ8J4VdJZvrmNwt3Lc
ymwWdjKWQ6Y/BQ1U1Wo/MCVhmAzp2qg0J+rqOU+MHL4PjIu6ZEaRou+EIWIpkgEQlbSN7odmJh+l
APdxmU04Pm46yHWMc2DiVALcTU5V8t5SLrPpFqE1n0GUuC0IL/VBgdtJzuCtuDLivlesgYoCPOEc
X3CrLdEv62q6eZ6Bwie59wEKmFOyJHr2K4YhM/0CngyO7vRv1lGZkGCjUeBxH8ukVZapPHrCZFvC
a8SRsHdo3pMCWibHCv64G/67PjoYFzxhadTNooHnWuTO+M+VseMfDM2EsopAz1zuks2Fjy7WtuAl
N52E/lP5qtow3oKVq/+n5XcHC4XrUcqdzz1fgybiJzUw/01yuX8rkC9aN1ADfy5qF2+Eh5rQ0o8h
1jdxHU+zFRFAdM/NPtD26fkHmiTaIV2LDKGm6GQ9wtCLd7cwb/RtZWfC1GFEw/7UJVe4gd6OEJt4
lyumGN+ZQ0Sq3tquGWl+FAzHd4GLCpGcZFAYKOKUIXJG+6P/kow/C862NPUwQqRbHta4G+xE4HvZ
GzulY3lnHT3Uc0NL+o9ginaVd61nvyhFWeQ5y4J6eNCYP+toJBp38BoSwxJRk+llL/8NMxEcJPir
8JrbXCgx6n/qTEKuvidBe40REuZiIqmdlCpXJKeCL+VC9ajaoacMAhKlxatuqeD40oX6Fe0GX40t
1oD4uF2EpYtz88FpK+0c8dpzjpuSKTU5lDGR6ge85XDpzwdzPhZGktSMc3Un7BjlnKzxiExcg+FC
5KN1ASWVeDs+T8GoRY/5jHeISjLuFjzspFI9WtOLHtowtO3mx1I2Jwk7F13OvMpWGTWu+dYD98Bw
FfehAma6N3KM1yPIlOcKX6P5geISC4lkgmqPdLdERjr2eFkqP1qmx+tBQGy7bLIFMsvgR/zW2yTa
6mLcrf8d4RRSYISVgqnJduryZ+ApZU/r7RsCapOOQ0BHWTUUoE6GqK0dmwp4f8nbRJd+knTfAY9M
bd45Mtjyuz9fQwxS3FLlHWkO2OFqM7m8yfWRbepi4aMKyMmTqC63smWWQ5PgYyD+k600zzhSBYbP
gcM0yuxAiDRyXlYbAP0/Hsbua6Y/q/KjoILHoejj05GpOEQmhDqDGXcVBJTF3uCarG0gHaiDFbvi
z0lnWpuyknspc1Q3CYOzN8oeXUizZhnvtaUytqo0AcWvtM44/WM/aM8MYJ3kHLjcZXw4clkcUYxt
nQ9/CABTxwR6lzTe8EqFob3z0MnZSVpeCN/dQNq8aV9MtchJ4jquK++LO5O447aYfKKP40zAn50q
WpI3Yuxe34v3B587FCy8Ppzv9u6R01f5ZFtrgEcwY1ITtJ1MLH6qKvbHmBIvj1Ls6JQAo8jh14YR
tQCjY8mVE90qv7/bm+ZZGbyRrg9tBfTHBDSuG36UuWB8Y4OTHI6LuGuH48YfUcmwvwlLfVgY5rtI
EmhlGvudWlQeM8vUdCKzTCCr7D+gSBErddx2B7/6TPQVO7cH6J8dMN/Hl+Y+ziEVH8zX3ci2WE2/
L+Mrk6aCp3RSwk007bj3/3Ep8vEKZ+2Ym5m4gtSF9Nxpy26cUpzCiQku09Gzjy+TydezMmo6SKIb
B2x9GSgMibQ12BGyGYmvb9pxPjbLkw743PHllypoGSCKMoImtQvWjzeiNAhFPO8HEAv4aqd3MQoN
I1kmc+UOYZQS+sQCNbCBD+dqkMPPHZqkSJtkzsgY3VJOSHfEC2mvc/G0AQL/hfHr2mhRUMBiIAxt
AxcquGBK1H6dk86jOCtyP8NAc/OK+AOrpx9ufGqr4BVdWTBaGUjHxNocS4UFVKHVaKq63lnkPdr5
uzmgogJxGqVAKgodoOpltWnxyr2f60VvSI71w4xLn8c2qRzrGEIQSYKLXfZqpo8Q9zYCMZ+kXNe4
HAFYuGyldZH9Oc+/FoWtcGgBXiGRu6MYsSjilYwI8segV1tN4Bw23g6pgvczZHuF+Fw7AuUangGM
jgokuHpr+ChlpSYoeaVvJz7l9H79nw6cfmy6gm0y6C/xakxLoEtqNRvwOPlN1w9EQ/KZSUVmhq4j
XFrDyPBaz+5gZFGN9LmRQ/VAkJKYTRcqlRqpJDNVwixKZZIY49y/j0uucFToYDYxIg/uU+sKKnz5
5VUH6IaFSD0/7aBfLvUWsh/OfFzPSD2ZwvT2bg4m/9EYE7DsJ2W/JWqkuMnyFTMVFxF5qHwpyQCD
zLjag031LGLkmMPpExI78XcRbTHpbaXqaal3SmJG40nqCTNZoPNf2f05Q3YzSL+gI2trRyRBGkC5
anfIaQBoCvYxt6bczLg/UP3r7ufcUB7PfAtc1yP7atG3/tsJA9f4V228i0dGTmADFcQ1hy8lqhHL
1f/9BR+8fC3o3ZwksXfYFP8AjvzzqgDDI97keviJZnn9bvZNwcqqG8fypTfDWE4cUCElUu+6HH+n
T9+A3HlpEchwlk/B/T09nqcPRIszIbdFxH5LO9KjEGJNZSwtzkTKRXJP+m+5CsLwPA8uVCx5gmVD
5Bjo6mt8X4zcHrOod0XTWGTT9CHuYgx2kZ6xUxSSjWfb+kx2cQgSjvmMVKAKojLNNRL5PclJEs2w
znB7uOiEAaThNrsiBp/K7YPZ0RSQGO+mJjNB1ZW1gMb1IHcY279OSJQ1JZXLlTdivaI9wDIPVCPl
71QuUrEutd6IvH0Uy7LJDJIrX5FJmmujMQ+kBStfao619waw+QPTOaEeR5xz/+M2vfdrOXZomChN
tl4fr5kV3tDortAPwYOgzETc+CS2IYbmKvCVIjOaVm3bqMYrGHI0cX78hFK3yUNaGGF99KfTmIiE
RRvSPwCrBLms5+dfUR8dqWQWXJypnaB8xQhw/SUwSPffx0qrE3u/fZqMY9KM/SI0Ehzbcy+CSzCp
QMxRvtip+/S7DyjHeU7mV/fbbBArWP6jvnRNkaP/XxRb0maKAzprWGOXyQIX6Fxap9MhWm9+w5HU
anhJA39XF3W1dVeZZs0TvbOUy0ffjJaRJ32fKSF6esna8yBRXra/zU+cODU9PB8tXuJQZnf/ogGR
SV5ck+AGdRZOe0JOC0qP6oHt+mw+u/tCpjrUOc0XUcbIs6WoJ4MVIhjj5ksxWWLT2SUab2jYJdvp
bGhkkkHI4H87XAfXvJykvrUi3sIpRbqGZZAtpn5xoHDbBd/gb2DUPdAyRhIL3IynAesT5PQUTqCn
TMuUlM8g8dLpzkCO66tvY2iMUY9Sh5jBn7x24WeFyEDmaKaRwkTST9wXdSZE+m7O9yHsnwSNx1Qu
LRtBSo4EhOZDPf3yYXDLgcWTSBexaZDePsjkV+64eFSV98eGo9oQW+7Z9Yj8NTR+pJyzt3ClJgEm
pGrhoj7C7E/7xSkrwUlNnJ8DvKfIee5JoNL5OgmM9H7Os4u0y5I1XqG2UDFSeFr3bSFil0nuDzxG
lOwWZUrUsYkz9hk5r8NLqTVLurRjRbAvQ5OVcg6KcxKGZNBun4AWzV/3IqqmmmVCq0UqiN4A1wPU
bNEEu49HC7ZJoFqWNpLfOhVjlAMHxyJINt52/nkx7uuTnqbLQUJlC7cumoq9VuRb7GrJlo3dttv5
wuSLGiPRHe+zlzUR0zkbuE7fmUwbXIDtnHsf00JxehwoNRTMv7agN70gOIYjsp2fkTzgQnJk7nro
z44qKZVYPM8+EM9Q8Kbo1xnfMiHAgl5KKHUaLqgta6RIepE8mgFaosrFdeD37zyr4mAvJRCb4879
oNQpHxb6ITZWpi4PPYWAcJrV+X0LbA8TBYpIm8+4PGFxXlUR46b05D5djMmPU01Bjq4T2MfDx/rv
twu6QaiQWqqJPZYQnjCKz2RVnhh4Lzk1RNdZhjnzHC/woq3mJFfzAWpDGbb8fnaQruE7q9sOmpUU
g5Gp3t3owJCcJZRYQyGBS2BE9GRhvnaTPyQiNhD6jorxmqRKx85bH36L3/hMSpNZXcRXnM0xF5Uy
6gNK/h5mr6o5kKR03OFYoufREAI3XWUJZFXQbqT4g8KBg249+cl8X+DZb5aGoe3gwNKPpgswgmxp
MGRLG8cxqwh159zrJOyFrqNKa2zASHQKxN7dSkmASB4v7R3aP+hbAuAbZ7zPL1fBpEVmx/6aKmQ7
VEqid5wi5Y69JKGDSM9FlqKN4Q3iMVyABpKNEqbpNhY1UUJTZjq/eSEmWF7gI6zU/RZqPz+pgovU
WE9a3YMUVCKqhhx7Fo4+PF+F4cYp8Uc1JskpUQebjaGih8p2kb/KVud7B69mAI2/oa91YYOJaYut
Gtvxes1JA47Olzi7y9H3t1rZcL+pj9vU7BFBzITmbDLK0op4CI60XPCt2ZIQ80VfEI7mVemiThKV
uD887aCCgNvo+hYZK0TG8j52wEW0A0+DcQ3o+F5UpPZJ2sbpuoWXzB4u1UARrr8d9xctKVjshMk9
ZSgOkuZrLcK2q1ZLakERAXGXjfaOm3/LCjhM0F0v6Mb8v3R6+diXQiTqrB+CBUYPOCPFdYomJP2X
NAFpJ1RbYo8hG3+2P/HGM6E5qwLRpA7C+vfrwIfl1tMsntnskyQoiUpV/lZtl2o7HjXeaMzFMAOh
bPpmddfWvP1B7YGzVtN8PAjluMeoG/nmRobDI+XJ/iyfs0yKaQbcHEYXNbbk5zw63RA7MqTfLKvp
+ikP/OYbgAH1Xi//N9rvJM4T4oNqz6LeWxc8hk4a9eOnk9pECyAHh25C3A98H4clB1kIJHfW1SxR
v+wM/EWqTm8fA+5QTr6c+ZWwmLA7CU1vnUg02qFyFCzuEy5GMlgSUAyKQYVY3YYqwGUW8VsS+m1E
AsYSdJiMR9DKBd3Ysdrz6HO+Je9l3zasfzaHXDh+tnj2g7p2z0l9tQlytnpRr+Hq0fpPlv0+YXy8
AVgSqSGH8PZhn9lObvynNdnmrjf+UsiH8AQ334wXW/mGIWgWAgIDFLUeW97NU+VRarb/xTSe5lQn
CluXEZwqCtcs0I2Q+EJs3LiXol0iQypndWHFOV/oUXV+S2IjqHJ/zRB9Xk0SS592ZB+C+k5L1YwS
AQYdpLMNLGRMnWqeo9XcYRCw3ef52FVuUEYZ1ww4vYhRZO8tLTfRpWCXtSGBtXk3m4xnHA/KEA5z
iGYCSS11LyFC7tH8b4MIYI8ZZ1Fjb2Pkja4HqD6Z8BP0eRyXWH21zNfkjKbovtwpV3LctuFsudGd
hDBYHiXfGlCsrzY0nmXSYSG1B+aqMgNg4YYwVZqnUNzSMlK+r0OwMSpbpJj1R7BjX4EKkSZIDnNj
NLDtjtFybNn5zdwVB5c4kV/P0DejW2mJ0rgb8zsdbGUKh0bJSMVv4El9bHLsxHR82lYk/tJWhPEO
bE/vrVUu/EqpLHdMv1YQNl6TjjIMk3nN/8hm4Y90J/MJXQ6XcSgCPoavfoE9VJJsscKwx/ysup6b
fN13BQ2FDU3GeyxTIDMAVjsT6HBZDyW98yBHUyUnfoqmTXwuIzZcWHPC9ub8rcm87N8/RlkdsaYc
3WPAoh5AMRg3mjoexJekGUJxu1KmGmRp2mzyC3ipC5wIt38Yu711mEuyiHyRDa9dBkNXsauwoYcM
eNovnhO/mvBnWecOm0zaQEm7snK7906NfqOGlT0AyximYwKDt/QoTZDeO07G6izGqJ8DMZ5fnGAS
jppcxI18WybxOFeirxo51gz2d12iaqzR3QUCJGZiEtqra3cvrxJRydaes/0d0/IwBY5LRieKHRqo
5DASMXWM6alhlRZ5+os6HbQe7pWdjecRzaulnAPKy23yVyfqEtAm2NGrJUcQ41LGdiB69mxEf3hh
LOHo8yPxRUm14wkWApDWjSjoeWts0VKcvU2osr4cVo5uMIXw3yjMQxUURDMD442qyTTDvlysoPi6
UWQkURpMsu1QXwiFA3hQSQmeqeAsxeNbeBA14md7Hl0hS95TGyIkxjdaebeU8Cl8HYchG6zL5yZk
LIGBMcalccYiVg1uDK+U9hS6maYFAyp2kNTHFmaUNBqw8zY/JrkmSu8aPRBtr2Zd1Y+RgvXKg83u
kzo9cj83tT/YQTqYHdkD/pG/y+qET4b9xNnqRq1l9sxTk5gmcxPMxzYrqZmnm1kQa7g9RFZbX9LC
R0IiQTvRSRRFzrNkp+1PNnGPYLtAxkv9LGC9ejVxMGDmZqJTrvxZoMAifeSZjWDPb13R3TagsE2c
+LNe/q/xKp9g+MJXpW6ksfLVzxDn2hxArL3eLGdzDi0HdbJLy1ycpkaudU+OI7f5F6i3wMLHZDMi
REo33aI1eYrF0A1RVEdc0OnlKSG5jg4a+8VVHhQu18Qrr2NWhXpEsb6pWsBpyNNII/H0+yVmaVkc
RejRZ3Dmlped6wBx4PtAOLqVpuzjP9xjDUi0Z/6BxZQICavsCVhT6/rDOXLWXoF+1rv0yRqZz2Wz
ze5hGcuDgKmIj3BvpEheChRPKAD5MzhCl5JlFT5sXJ3VEEaZPPfArnAN3AibmJa0fEa383C70b2k
kc/bMBJ+Yq8k5R9EEoCPv5Lm/EgxZsNpcgUfeze5xGheQtJFtQ+nCRud27uJ6wXQIT/Q4b5mNWW1
XH7TXFT65DztcVvwd2qvE4mD+VmDZHZCzCyZvNhKNyfFvhKgInLDkJcjiyHQSDDo6cf0yVYo1Ryn
W/bDc3Hq7yE6ICgHgsYaofi6COaUuyWIbUDpX5l0P2lnXL56O7GpCvIhw7Yljt8e/e4NN2B4iU9h
a4np4hCnWJScPxSsx8pqQE9JGxDmiyhQZ5motER8tP5/uw/+MAgdV3CbFYP9LigEyZS8UmZPWlQ7
rTFNVeyNKh0x/Uoik167pD7lk2L2l0dFtuRUEI1l/gcfB6p3vR4Q3WGoa32jS1bwFmwtDQi10ke0
wso/Fi8MXtdc5JCFiXV1lWj3jNVnStQGJE7+JEKT1rlELkSTAZYOOXOMXNKNFDe8tQngg0xeTiCC
Z796Zeccx0ad052MmLJ0oD4NbzPw1U3RQY8uJ0L3HJQsXD3pZDL5hOTlb/TgMVABBTYO9L1MxZFH
wIl2g90dUoDQd13/oSIIwd1Mpf4PXef9IyNStu/ST60dPgLroVMJewoUGe+AU3qSP+tkT3dcU8Ii
G3c2a6pwlyY0apDxa/nt1yDftcyYl/F0ZxqPeBduhnzvVomC5m1LEjaqm8Duga5dh1IpBm2HJyv9
MjkJQjnaYY2iK2s8hYJZZH/bntDLKr8ryOS32BiFk5Adx/67qxbYvAoNac2aS/wS7O1FQn1HGbDZ
Sq+VusbO4WWPrrAjC1gMeyK40K6fdzw5a97Tpp3GHV/C/gYXJDprNeY5gqlRONjeW5set7a+Zg7r
cBj7L4DFwC12nzLtnicZqyKnp6rT8xy895Qs71J30eOIeMr66U9o5OVk+UbDXIWv+2gV8mXyGj5F
QS5UnlCB3S1W7U2KHGPrDEVyuFcoyVUW6L6Em03MRW6inngn5zWaOQ/HfcG09QEIpIfSr3g09G03
BmuofCCZmrti7iSyQI1+dkUP0jjkyfx7Y+QqsuRQbcPbXnpCCHdDYdE/kVypz4eF2EZFoDfVXTfn
7rJY4siEQ+mlFAxh+kYx1ZTUiJE2YI4hD7MenazJcE6vt/sQblzUF9Eb89j0pJJE3kVKs7sr4ECL
rVsAzLElEJmz6thVuNeGVjTK6kcgsPfOaTOFrOVVz72O0YEVwJSQhFQEzxhE7IrJ9Q5a7kX8E8UN
2wRR5OKA6RzoqR66zC7QkWt7yXM64Mg9+KJIHLdCRn750FhagpJN+WRgoplxS/mCfYRm/boLWJt/
2UXcsuHuZXCIcNNvFdRD8E4Ivs/5i0itza/vvbWlQdr4s3bpdycHBM3XFHsJY05sxXWXD02S1Dm2
5/4S2odQmNjJyvqLKkhoQg1X2efUpCsTDvYl7mD2zb/ozTloTQQSP+EvLb18Gdxrf18uh2a3msjQ
7e68t0OT7CU0FSa7Re9szGlKomWEU+WCKZxPLKAmsoUeoM1FvvNrwt+V4bFevLUVmK7kMismg0ps
9PQokDSv84nUs9NyqOdEvAaAvhHpSb93EN1cVPATuKFhaD523IRfOqEupzWOLiF6PIjTgISlev35
fHrdnsH8bOG/rWz8NzEqz8osZPPHj9DA7xuuF4afanBcsAu6OSvUPrgwSnDzrirFeUf6Wl6zqsp5
qVJDinx5Dmj+dYsGSgUtU6aFS+FE7Gm2PKsZmIChq4jH8cSOF5iHnLvBpmqlC9JFCPNmTtDP2xVv
nagZng59BkPNxt89Q675x+EOFX9QVHV+O+KbATYVMh0KXcmFaGUPAUW9yQmFF2QTLV3gwgz8Lf0I
Q5nZnjI6PdKMIeJR6RNm7EMzPpqZA17Xr8HAPxs17HWebFzWTjG/Bo/jGaDztizVHBoT06fjFdkF
vQDr/mXSpZ2yq5D2e2dsVhkuKEKF7YhhUM4IvWVxAIIe5UGFRtefth6JDuJJjGEEURzGG+lHV3am
AVqhTYfTn2QwiPzN/vz+ot17vXyw87d2tzuOipvzjyvz9ZAhIZI8oNS2y6RskQ4Fj5bU3zLZbuEA
6ASk7n5Pw34Taz9lkamRYt/56q/r9veoNzffiM197pXRMuXSL43gOcIHqpaPnpxQll6IVAyjwOQc
r6fzsdtwMVoNoHtRxg6nlMVOHYo5fCIzKJR1985eQoedCvpVyrephQBvPfdwBfDKXWkVOFbaqxTi
zd7pFw1F39yDx2hkdVMkjuIjPYODmPdJZc2ejvLKXMo6Us3VKunCmZRdm7Q77iCGUH3ypmxMRa1J
Qcl9ZgX9ambNnNuChHX5ugqFL2JRV3fipg0nZhWRS7EY/JLzvPThzXzjfFLHBnraTul2Rv8ySQtB
IJIT96N8W3tNla8u/W/7NZuLlZPOKmNttj+QPWp4eGXfLAU4SBu4fcnSM4FbR7uq4EUAthTDhUzJ
xM/1dOamZHx2lRVuVOASE+LaPaS+Tb5iv75gaSDhD4Qk6TZL0X0fmPxZscbMZtc6eMNVN7PZj746
q0qjgofS4NYY3ASui2ZuAERfTnI+KhVfNRib+XYvr2etfN201WFgJiCVvwtQ5lAImMaqbbPtC84E
qf8jHXME4RbUWVgZhcyyrSftxfxd81vWZyJS6RTkYqabHGkPqqLCmBCm1up05RqdtOsBGpu0rc6j
6hHz4VhfIZ1QmxDb4sUQS3nSvBiEd6wpEuDAVEbDAx95P7PVgnnp1kTMfc29+XeweIiz9rehhrLT
MdSn0KEomqRlY7W6ETkBAXNhoS+hWb9W9S++e0B4hvCoVpnFwJVuhJgA3SK8+UJaKk6abojkqaf8
kjuQ4sAcUiFMAk2q2zS3atgiBp8raPBSk5nubfcFekDyELNgAu9QPCMSm9qtEkBUHaF9skdyHE2w
5NpV4rvHDyGFybdU76SVPVGhRYiGC6rZud73iuNdJqMGh/8cgulC//XZT1khCHczy16aNABgT0iA
MC7fVVQAdSKcvmAvC/A+mCHrvbf5zQCn70LtLicJ7ykCIDdBuX5aKdS0wbsBRFwPrTJml2Fe6J17
qj1eBg3MsaEWe0Z3Ai2ygq0EXU5Fa9vD7ps5Pb80An15WRTSplD2JyektHw5+TAcJlZ7Zidf3WwW
j8Tt6WgoLnZNSJxzV3gBBqgwOatpfK8uSefEcH5MRXRBtIi/DT4Pk2cxkxj8IJdJkp2STJSios7I
rqiIptqbAmtx8FSaQavZm8XBrhYDdQW/2Tnc7FtMKn/Z20jPrCAw75PPyuTMkb0d67pncxSdMjxW
X28KDUF7JuFLEdlT9Hmg3k8F5fzcp3VmHAJ3rQuu26P+Oj4rkx9YQ0iDnEC/sjoMeKKkYE89q+G8
WZNkvEczTtIueFzu/gRd76bKefHmrmnXaCpskbwUN+RRU2ZscbVZZnYW9gXpqkzcOHWgtf4a6nfY
p8KjT376Xmoh9vtIbWWUTipZvcDaM4zlI/fiBINVSdbDhznRhbJpRC4Mq+HXRUjUv45W1GRCh/fH
HU+Bke+NoMKc2RK1hw7o/3rgYC0k/MN7QG4VOEAL+391hNmLy+fByr3eRTfQyuuol2NeuNiPNQiJ
ng3mbAxj0BwziNfz/oVg/2SZGz8nBXOrS+lLH9ZyMLiM6Tsta/wUa9gYEPDkHIEVcsPCKrvf1O70
ct/LihrEyQIt0ZgQK4eRucPyvOcroUFUoqjQ7vtlx9iXogAdP7H2d8dMcEuD5ePfzQvd7uBYl9qa
/LfnVWXlRH3WLt1Brgdirp1qiHOX0wb7rxv3Pbc9bOnPxzVNCH+diRm+9NQTxcYBirtkjXwcwOha
vhUQs4Murlu9pPXgSAHLTZuGNrnCzhWLldGputv4OD7jVOzXD0as/5pXw98IdxoEaesvVyzciWTt
IXk3UdgMMqjdOOQOeUmIRMf8PM47sUAf5gYpXKW2lbdJ8OgfDQADokjN2Nb0vI7NF/bOkvAit3wV
k5zfpUaeEtAnHfyshUUg/HWa7Y/QbSAtEeHUewq94H89APDC+BVMCc4pWxx+xwqcfkOO35mDaN4z
oQdJsjhGoL0ipVvYfFAudCisARy0J6gype+f29LcMnoZ4zL8uxk1YgGq+PgsKCVXUXaGZURa0djV
PusJFaiXsHM6Sc3Yhh7m9wIZCyqowopz2tHTNNo3vNi0ypF71LkPG/nYgbWUOpx1DEeYIZVa3uBT
5LKIFbpKc5+T5HqYoP6YCra6wQ/7HMj44DoKv6KFApBkAkix+PyD88gBWw867Gt3FGwcklxsUbnH
JGb9F2XpSIw8x64/PyNDS5WCB/effLemKA66AhkbF4DTymwy6T3IJqtWerEv7DZNVUmOc/hs9cMm
/J3KlvXih8Lgjs/gnhRTxxdAbh+IcT0W6nwnC0GLYCfombUussIDlU3pyNTpcvatW+vm/QDpUnC+
OSZIKXzMHKafjaXrswMzAf60unTNEIVrCsYjzf7fU/NHcpKxJEI7bncGYj5kbUsClThi17WDpP6V
huVeB6+4dLhdR/aaETfZxWeVMatksAWiCufMJCPklGMJ072bg5K0DBipqz5AM+8qSPAGJdWWapbR
pkifRuPOVlwst5REQN4Agfzb6ZJhshMQrA/hgVu3W3s5nGmbVAOpwQJnozu5uRtO2Ul87hITWu3l
op48xywac6tBGeoed/ZoSo5UUlcBN3GN5Mnbu3u+fdNQ55w4xdGY3Xn4KxYHVzaLkfDCmgppVtQb
zSk87HDr1AHjr6/hD5YzS5I8N8HlV29U+ObpRneX4QdMDss5sTcMTiJE6aQ5zj7pi0fSwmEOiq02
qWPVcw9PW/ESmf9GbR0KHhcyploqcYLewaBdUAED/uOu5Pi8D03UkCCNsdLfaef339RbxffUu1sc
2hOFP1JU45NC7SQWrpRMvIhNF6l8A38xNVF7rW5W5T9/S52o+6djkp1+9pWk1I+uMeo/bfERq8cX
QfkppCXHA1AXY/+ShIffntaSwXkgBX6xh/lv+vVZPardGjknPRsflzE9APzjPfuVAK+im/AwwCF9
FO81rNnSrh9ba/CqWZ2nQjcGwJTfV/iHKf+4X3kMZxNlBALygb4leG1NDR6cyIXd+0AvEXx0rwJt
C0pn1Pm9RGAgyGiIsX2q3Btua0BqzC55QZizJ6AESmAJ1BmwplYVBc4STf/9O1QhgmkyB0dZcZQN
BFHzHVW/5ezAlz+XpBj/nBqzW6p6oHhnzve1EuhIQo1HJqS8anSG1NVVZtPB1QDs9UGao+yei0cn
BbuVedpBc1Ml5X2ex7duxmwQbBmRpvmXrBoyFiiA1T9Stdd0Iyz7h8R+Y4CvpoSc0Cdpqu/iL3xj
FxNdiVKy/zsbb5X4TggxvoeQrTxVu7BvF3adf0EWv2doLPS1LFxzGyUR3U/QfjbQEz08UpRZJRr1
HXIjwtB9yMOxz1Xw4k9EMrgqnd1XjB/4iLRGAYnvsrUhTz4gyCM3cJYQQzGr09tx1MxGBaGtZ77R
LW0/ExHbvG0Kelltlfhm8jrXixOprrAXVaMXA11smbTnC4SnD8BfQARA6wB5TZ+LonhsEtFDaOKE
j/zteeA4pqgsQbTJeu2gp79rm9ZVhpwDB/wR3otxzlMVgWQqSBSLghljRcTcWTef5/SAXGa04deV
bOgRsQwqVuqZg0luAt5fOXsY610bCBj/o6b49Ioo9fl878wEf++c+o4EduwP0UITwmLCQyKUTBHN
CQjFOQSQ7sU7+sjJGwLepODKUW/kvemDRkT0Xx91ooVxSwyzLAgcqxckKX+dh0w+W62+w0ljsMM7
k9GqENxEaiutSOfMxPjws8UFYACDrUjkxPCgwNyurw0/qOKxoxV3hTEDViKNmU689ZK+GijAWliF
W/HJ9dxc+upgYHCyZa1BnN/6b40TDksu8m22Kyl2bMB8RtVeC9dvZ7C1AQQaYyo++uijH8hVM2ky
lQG36lY+O7nEabU00ni/EdQ4el4vI8boHa/ur9TwFHErmk73CP+uqe3q4NyzKk7K2gZsidNhW6GB
jeR7Lzf2NVa6ivZdx2XnEVR5Kl97NNuUu0FHNSxJsfBe0SPJE8+aopDuBXUQCx2ka52PMJ597WAb
c8n1wlUuMLsVb/fRx5ErMkl+bBXAWBUV2IC8LXtimf4bIDhbqaqSqca/fpskfAplKomqA9lyqj7j
23/ltdbyF6lLmeQzSa3YBZL3qZkGjRBMlAruhxAXV1hluCckXU2mPx1uwjelECnSUhNHXfo25U3U
c93OPaz+zufx3GZTB9K4QwzTREYgvtOvAmGt3i5bKSXtiD1k/37a4aUtxVUVThJccfXsvCHkaLNR
qCe759MYFoXgsMjRJ9VRiDJadq52JyoEoIBgJjvoFWhiQLLY7/yY+1km48LnyVVDFY6b1wkkaj7I
IHgmQUl9hNUG3WK6pCA+a+cz5ZC45NMYdtiSvnMRBOgaYhdtEaRjxao9rk/e5XbgZE/9bTYN7a9d
1rytN53TfOIh36KQNklLaK9qUPKVJ3OvSMn5F4Y5AXXYfjpmUgeoaUt6G54EGgwFZ2g+tSuwFrl/
//YCtDx7xQqpQRjBgIxaPjiruqU4WvbWk7l+mfUD6oN4oiqQGzCSHoxNf8eMzOX6vPSW4uo/QXLR
IMNhSw1EI0GxHtiYiXdFKzMg1QTcbs1qgx3yBdQXmBQDCeYSZCCfh2rzhX1fn43cRH8C5zr19ecX
2PwLhbsBtdDgmO61j1cqk+1l7/5i1pPE54ryjuC0C9i9lVUQmT/zlF/kwIW80QWFtYtGelsIOGxp
eZ+IhyqDpn7uZYgcPg/pi6760Vy7kIndBolTjQOU0o0x73HWXIr/9HF8VgA8t3qjCnDFUmgEqZEL
50NeLK1FY5uCLXBWVHHsCbxNCw4d1fYKu/b92REFuSOHEWFBW80Z17zY6rOyf55bJNbzGkWIBCv8
Wz1EU/zLinJxUvyWDuzCxXuNaXrdrmubkaZpAddUPyO8QgZ3QiLYcyGJ9JKSZeoqQubO4qgQFMK0
k7n4t/dCrzb+zLxTqRNTiyNsZBc8jGniSUQuRi2LoVHn2HQjpdk/CSn6J4EUsbEYfIRwQ3/vPked
J4XpyARx/YwXQzLVgthXa0aXMDzDyP90h3uSxUPRe48nv1xJTJwKe1jNbv3StkUXRZRHRHzHWHa9
YBVbt7+/Sk3yAiZaE/lF+D06D9q8p6YLAi1mw/z8QPfpb8DhoX0taq13pSSjaCoIbYk44qTKoUS7
H8OoPXJF8q5UGDoVaD54XJX3LRWOYnZfKibpDRUYYOHzthAizwfDo7m144GqolEhAhYb/oHRiJgC
fTvUVdKanm6O150mutCNZNBdtwopbmAbjDahwVJ8jfIas2iu+z6IjoiROg/J3JmjJ1WwkE1+YRQk
voGwzSsY7VoJmj751yRoCdhLmIfhV6vN9xoP78bYMLUd/8yboQxHYtvLPxetep1XCIcSwy7+36aa
mnNa4S0aUXYrnsKJUCl2by8hY2+PW6Q+rTSiaizhtB03MIa4h7AmNg9IKL10yyh1QGQKPt8+5paN
Flb8kFG4lzkmplrTNq1Q2SuebF+pZfEDC25ZDSDDZTeh628rufocmqwXof1XgH7fvJ6/R1POhykM
NqfoO9pU0F267Nr0Y9UOx/hKKJb1AIuXp2ZUdiNDsACw5D0MQNHqUiqJ6zvvVw+itSAhv+kC4xHx
yKNa+vhk9Yx/NOmWV989Y3T+S560p5dbeYVoFvux+Eu3wPfAejNYTlJzI7RzebFJx4P78/IrWM74
r/ZiAuCrCs8sc4/y3VIFvKPyH3LNtdEIWa071Lg22zXoPgxxy/v2L/Gq6el0F0q4WDANJ7UgjLuE
ZDcm9Mu+uMqrAsT9w45oBViTmkPA/jgMft6stFx++QzM3krDddcRWReNN4TVOAg0vZbyug0TTM+H
pp15KJd4cF+7e9w0O/w0sAltDdccNDsjb5xOVm7zZmqWXphCw6QUyru/eOqJIuQ1XpIhjJJCEXZH
amP+hV38ZJSA2021TbD8MvlbNlspsgph4SiOZuD0WmsxjyXgiBUfei+Mfuq84/5wxu+YvFKoq5cy
c2+/miCK4HKP01pCZthXTyCgNW5hbvqZBYIZD3JB5Uk3hwdS/ykVXpW6OYPqv8QsC/B8a/5mDs4t
UyPYcEC/TSH766pcTIKshtZ8yC9/CpT9Jg5OxZxH7W/rS0+FEJBv/atv0BiG472s9/2TwWA607fj
StnO0UjjcZMmwRqnA3QtluHRBOk5gwzTl52ELcTf/F7rX8o67MZkoRoDZllkZhhk3G5givC22Owp
0tWjWT1qtbTLaldvqAt0FgKAEU0FKYTPH5KbdP5EiXXlT+AHvEQXV/4waAYkxKu3SUJD+wR/EcCe
ZO1zTgxor9qkR+EmdLgpKhzhFzmVniZ2P0dRFDR/lzU/u/U6nqdECOZdO6rPpTQhxdVv3T09sBhi
Ow9esy7lGeKoBGB6ZNAR7cr3o3HGUSQmo0bGcza7BQgh9gTHwNqbE1KL3FRYFsgViemlMoiMsjJK
bxX27O89scXbAz1ge0fen1YuYf96vgQ9QYTRCHLKtRqS2J0M56qGXANnJM481CIhDQzOg5h6UL8z
v3IfaChY2sDS3zQw7V7jHpEvX3Rksq529bqThBBJXGwQioorVQukY1VTMm1hIBhSVUEsaq74e3uO
3TH/pYcNHTaT1ED9ZDPeLurc8zFqlTJ49G3ehBULpZtAZd+HnlFw0cFxcICnT3VdlCLsWvl4MZbK
HZoCqNSrcPfCxOhMcBaFUEBUdwtkz58iKv0xOg/JbOWIaMX6SZUoY2Xk2C2gwLpPZrGhtIkqtWJK
V3bP71sQofOPwdSXfW5dAEChJto8EZ/DLQlypfN0C8y2T7TmSAxvHqeDV6HA5eAhvAIAVRlWodM3
ZhNDG64NoK0KyPIS12j5HKIxW3wUA6dXRseU404BAT38a/inBcCpYsMmDEMmzCer2zTf07r1uWaF
iLoG2zzUZ3mF2C37Yt5ahmt3aWudFIAuTeHz3qWKUez41c5zTfRh2IWCaKhrbTINH22Mj5D9qvkm
SooeZ1lcmLfL4+AfqVPh/LAvNl/QvusC8vGLiBoi8vJgXG/ZKYW6362zrmmOZ2YTGfnpDWcqmh5t
6WMHiwm+l/oFuua3BWFk/4Hj1ho3z6ZV1KXbU5ODPwMmYTPeuobos6XwJQKXASceIT3D6x1x3seC
3y4Ceq8H2yMO76ZCUIyEgFSHODDAmZouLayU6KhNko62Kzk41NR2SBQxEhQ4yGe8wP5FEMH2tbkd
wzi+VwYgSTZHn5rql7TRAAGodGSnowexyktYW5E3oI1RoFm1u7m+r+8etIR1XyHwVQKafYvvuwNp
KWA6z+jtnotpo78+mRHWjuPxdpws0FwtJtUTQ/So3ZKz7Jx19ZNz46cBozN8M4U2suOTDQL5+mKi
oK0BUuYhD7j1fKHwyICqZVC+bv3hSsSm7G15w/D3eCMKlYhMON9tA6gGFspnh0od4AYGomLKOfe0
tv+0TEVivFLhWGz0y3yUkv/Wx5/ZQ8ZZgkdNwiwo+HSJHyYmWxLquUgRmRZWGqiLTXVw5iMaGdmh
cWsw9qt6OEInqG0FOclO1QprWaZdixJs60PMg6G+f1koth+bG+AdWyXYhbVjKTufTdC9ppwPfY9n
8TKlooldhlEUKT+TO+Rhyrb0AffVAOmCizLkPJd1X8M0pEDWlhMXxI92t5LG1mRR+oCcFhSvHomb
zcJA1bzJbuiIqinDdxLr5CU+RV0Oxm5xdLcFtRJsOAS/xGF75oPvDKktX+5YhJwNnwmiJteF0q57
Lvako98/YU1xcRA//nZTNfc6LGXvHwdSNTPet9I5Wrw5R08R9s25+TYwmD0T+cF+u8o/HrRMs/fp
98f0VVUrqSuRHDEZpgTvnKkOfXrqcy0up18mEdB37uF44WhvJopRS7l8yrRP5+5UHNf7O9Fj55Xj
diNrRYk+00Kkt5Rb/ZfluUVQkIoeN4DiTVs1TxPYHEpg13FAo1dDOtG7Lr91uH8CHhlMXdbSwVjD
JIYXqbgvzXfDsBFixUJ0Aygz+8yJeJr+IBk1Gxv0foYu1ryebfU4BvwGrujn6niTh9O8T594FqxK
0zrjlPRT0QnhnQpQgnRBY8OTlR1caFI0vUIwNN0KHv+sq64sOhx/jibuE3h4Ox28svYoQs+TVF1w
R91yMjlYLMdbYuxyMmuukxxISMeAr/il9PD0XaEhGwnzXaPcvzdtfeW7panBq+RErR3Uxnawu8GK
iMs9deSf1cJvUfqvNM/Uh89k0a/lbSqT1lEex31K8/f1sn0d7Lsfd/pJ8vsT1F/BJy1+qd7QdQu9
Xt61AqPVq0og8q8EU2MyO4wS3r5sNzrZKs1gEXrtEbptZMpBWPoNvpcYz3cQ78+SUoGTmmyK9wMM
s4Gj16KnhF+zh9otMs+017Gc3UI1iPIpy1K/+3k2uXxMpeFN8pbJWImLW93vSTBN/whJXju+HfkT
Qs/9Nn8q6A5ARV9xIMGQfeCOT3Pzc06ch6bJcHbjPiPm6EAnMUmZUD7Kz80ZvdrIWrsEBFcCF3E7
bDZJPqOJCK3pAg4+ZMVzJzGzOMKJR+fmREOtePby2wKLyaPgyMAXn5j9xuhSQi+scOy1sVa5P3dK
kW8M8EMu+axycPAAGdtXAJItwVE8sXRpSFgLXZ9j7SBnua8m0Zo9d8WJivDV2bevqwKFzQVt+baQ
4JlKxPveSglDkiCRM4CGYMjGEqZHgc1hTPrITzV9DoqRe+akzw2eAkFcjzHdotxcEkiPpAAl2iTM
RdXNM4TNoFsoRj50yj/WTJI/AECQ+6l5JfNOEul72mmJlsunfEt5zSUIqOPW/dbLiNOvsRMviMNv
wqGYNAKrKQEUKtfI2ZBgW4Gxjp0DrC46oaCyJDlmBLMPfQEYmk4DQH6oQzX5q3jrYk35D8yX+geg
/3UCgZS73ra8ZTPvWYpxl9DbgEtNoDuDJPjbkT8mAVBZyd3IdWs+JiC3xfdTu8XUOtXVhrfaWcfO
V+PLmT58U2CMoNPGS2qKGWg5w1cp/oOCeahOtafB2G6Gc0yUESqlzkaynoizCBEQKhSzUJRVeKDS
ntH9HHYI6qEE1onWkjp6ee6WNAeEKE6B2q0mFj1Cq6K41Dr2diVHUxW1ql7JOnwj06URK+u5VFqL
WBbpbeCQA2Gv3kZBGNkmcUCWILaEFDimufZGihTeCtVn3/T7Jm/UJA3mem/YRU07tDPcpVZG3in3
fbIOtNalGIRheJR/cnxoOuT7N8oqSIhQE6zRtuoskJSOy8Zea254866boLtTTjfqA8E5NdVtFPC2
MPPNN1pwxxdfYWLe7RThIgznXHLjmBrc4/katuAZlAVNuZUM56fB9LgfCcWspGzksnfzUib03/Si
x+tRgFOYByO1TW7719IyXOjz7JeCvhBXJGufwOKFXaSw11Yv8/yVUq8iUDtF+faunxAjItlMCJwj
GqYalAmLj8JEJ9YwMeNZQdLhxOy1DkNeNxxi6KL8YqaOajxzGym4vwsWbnAeRxa1mDYx0gmqes3b
Tw29tMHasLs0WOOF+uqFUdFCsnx9ZETaSwKLq8ZjrOLqKFaV/UoqzxDFpvTB25IC/L5fKdexiCM+
fc8dSVRRV54/33q6rOgTFtcTHP+dSky93i8NaSWY0RjyWwcHH/XlimpgSjQKLwYhnuD+ZWnR9DBJ
rd+OX72NvifhHTSR3UZ4GL07TtU76oqjQeyO8DoxapUxfA+a5YDIzYqHHQl7u1YmZIPjpvF8fuCe
fNncuYNXKVqRNXeED1z0jJkHrJ2LAqMbDv6gefHyP+EYjEHlkt5cFzVY+RJkDJh+0Ut634h58mAT
UDKunVYXXtYJq3S3tI0LvsrYEUZZPOaO4ZAB2rIFTHKj9V2O/yGnoliNm7U27yjXmTy/o+qdtfOb
SEW/BwFqhgQU5BkIColuI8LPxKCEwkQAZuE/zaeZmjd6WHgp4tqd3fOzma/yRMrp3Pd2apLByphA
SQh8Um4DjOkL0mpmyj/ArJF7D1BvB+EtNy04hK7Tqq7Dt4EUmpOKNguji47OT0DzEURite8Lghy8
N39U9U1nJ7coLryhvHx6XkG7ItCPn9K0YV5w9lIztP63/13O2E6CLdhe6xWJ/DHczEf2PgwLqUyY
jtUu5YG3w26GF2kz/ZugwPDiHc+wlS7xeKxCydnB8cFjAo72REu1qAdtuXyHXBkBPtiSZeuIIwFs
vJBTDD3DP0H7ko/Ho8YKrL7pADeieKMp1DhZkVkduP6XDNcyRuXnSEZx8455cDv7vsu3gevRak4V
VTy9oEAfM0U+SsNbo/Prr4IsEf9w2UpDWgBxp5q4etvV6Joe4PAZe+2v6WutSjn79V6BwbnEvG7d
F7sJGtRLW0R28atlnCWyMO0W4+OjdggqFSEsmAPgLj9+GACnLsvxoExAyzE6OvkhxhEMhLFtC8i7
jo7vr6dE6Cfc+mmgIv6i64ecn4h3rgUg3T7Qed3GjDbE+wvse2P0u1cy4cjPQfBeCI/3BWrIXaEV
XOjxgq90ub7qzISp+/IZIuuPW18wZShKIzMbCByQQcLzmrYJCyw9I5feAquo8B09Gb7qAVMKDG6l
wGjDQocV/wKvYxVu4hL/BuuMyItKyZXcqDfFMn7JS0I+R9/JeKIJjy9I1txXClUPC+EsI+VI3Iie
3wJxl+p8EwiVIHyrXY0jYkQu8XG+2wH1OqkSUPFh9IVny7n8nqAu/R4o5DiXHyLtTflW8/XbnRiH
LO3uOMsnXN0Wg/fFqRr234zGsD6fInABxmrrFwnBNspAnxaaMryS4wKPJwMySFogz82ST6W0B2gW
8rupsHyTcu2ZtyeVHVWJ42QTWQU6zXkSjLwwXNgYvGSr7IeE0cCFzxKjeF398gor2ra0u2034mOX
Z3c6mxGBXuJQBnsectAoZ8hGwgcDqKrF3zE4gi+LlIeRAPFw6+oEJ1a/esKobbyFDNAWt6t+RsRX
IbFm3CP6o4XLDHOaFfx+BnRyxcWDFHr2oOhFVANfxQVEubpIyrSuAQU0yw06u23iGWwBk6P+hEO3
gFU7BF3OBPDI8bjmst9LFbqyoEU6Kcydb+VciJ5757zo4Y0rLRobvTUbkT6kWa4CXLMjlqkZPNDC
qfes/eUKvmN7c6IRQios5khrAwgUxB1ovlV8k1aQ/FHKitNU2tNpzJYm1iMdyTtj4MVdtKkH/M0Q
ff2kw/aIn6xi/q6tuxpPXYmPJIOL4gukFyTNn2dX4yugTa0ER92ZHNN31pr9OOOu45CwXDGEuRo2
T5wNdPobelG4bV5lcGk5Yhxv5U/sdRuvr+mbkdLxSjYUHW0ufVu4IqkRhAsGgzMjN+OmBHsrbLN/
tNSh2CLK4Xxao7XmPn1fMBJdDH4QRriY8k3jooZCz8Ee9adeJr0eu41GXaoOxEJYK07Ol2s9xD/k
UwWxGEOFcSt6pWUOR8XffnCfeZQAPrtEqsWkSGMlQg03oOwwap34IFJTnahTj4uU8fCO7dq3qRZo
tYytkC34bsQwGh36y6LZHx6hxrTj4ih5EUw1eiln5auVtiuUrtYNRO9FtfygsGhT3b3P7mkBJbI1
/weTZOmE7L2dRKM7KqYTRd0RxzQ8ctLJs2mIPeAUHtOAtQE42s8H5k0kKkDMHNoP/IzDg0fwoLtQ
OJ+Nq0jJOButmyUZxxQ2Lx7z3hhBENiODJhlzLROzRWoaLDiLp48Sw2fmPwJ7Wsjpg7Z00amJa8/
hBz8QnlHDu1jzufHsIvzGl5pRP4FZsN6RXEHYbzeN1wk5PdeIbInQKb6HOnlpVJz9p8tlb5wpG4v
831ELqJVMjCw9KGhEDtQmiC+vhgqDU1RfSp5m773C7iL5DfrgC+JwpBm/9AXAM/F66YUomxsm+CC
4v4Vi2xiBA5EIJtIdgyS0/jJJY0I42T+Kr49/mbWpZgQoo2/KTFtr3WMhD2AzX2xUgBs1nhGBMtw
kBs5maNGh3dBZg2LHqfImGsEjkF6u45Hz16VhKd45jbDfRs2bnxJElOy76GuLaoWfBdj9NnALvGd
5KVKvQj8hi0Szy8R/etM0SXSDeitILyat+pq1YEsDOiJaOEjXLdZgHBPQNNRiuBLwcGtP28Fu8pK
P6VeTS/AZwFOPwFDm/QMvn0aDbIYw5zFTHGLlUy6pWqZDQj+nYTL/4dmWv54O2XlzZapfw6OsZ0T
l8U6v+qI1me6afK3zSrbSXADecl03OLKJ2W4ImgVRIWyX7/L+vmL5psmdRlwrVtIRPuSUvqWGOlU
yfa95H9JvnGNP12Bz4YvHehAxjGT8crZuRkpuUxvj6qwpoAep0PxIwSn7exNiwZekbz243q6c4Dq
klQVyLWCiN6KFiFeCwgTjzW2JrVexoA1HmmJeqE+HqcBmOlQvzpFONo+TuVxcmOVqgSmKtHE0Zw9
I/ju4kRIGezREtJD8xrxGclFagTLOizgj0eUGM2mq+yIE9sPx03Jt3WW77OWFv/tLCSiOKRpxc8f
RRV1pNTdgsYphkAYNG4e9FgSucFKXTHES97d/eubMJCI/JwEkUpdCf0HLDex/+YzVZM2GTDlEPud
Nk3QJvuE4+QqU5GhD8L64pIzrAGmpX0FP86kLJmC7hW0iwLvNFa06FK1AqVPvnHYNAcrBdDdVVj+
g2F52aSAPwpLBQ8ntF1MgVJMc0sIjTNJkmGUgky/cthcUrXgBoouqm3quRjaknkIHlFmsAhwLqbZ
q8CZTsSs/kfWrXztvg80TfHceCjVdt7e7g0CZHjo+NbjhkWNNL4kMh5r7/pm5HKS/O4q9kVmV54x
QMhFUPuVEAAjoW4wgw1N2F22EYxreha7bzDAvOqrqdTmxFsaK5ehGAPrQwPhjZKSlQdMSzIXKL87
GTk0QuM2k7u3XmJV62OrGROAigJn6UsTSqMfR7bs1JGZlTW35v8PoTPaPrLpKAjiyHMlwzoU0itA
XKYbfh/yCKbOLLyW94yZfPxG+nrIL5FGGzZTEkhwjUNzr0197w1YbycMGqmOhFkYPVaYkJuai6v8
nMe6UA2BmQ+3lNY0hWbXgN2ZDMDKOkKmtbjSB84h9dRpUfnNrLX9dUTqSlS5JrEz51ZDA0H5d9v2
9u0kPy6u1EWNM3a+BGUR64h59XrdWA5OSB3uOa1LqMNtM+OIMBMXKwgk+nnT3UiPm5TbhKon62NR
0vsoHV7BuoHNEyMgJB7hPUcT9H7tuopxZR8qbNY9pezboDb+OXMUFbBUfeBmAyoyD81G4ezLbUOs
57EK4xxYMDaYx09r9Leu6Kbf6tRDaO48BoT+XdCrfNZfF7hBHVuKUvZqKenM/TAMH+hWrrM5k0S+
o4xQnII88cXxbJARAraijrDMbi03NXpPZOahaXvrsik1kYfvDTOX24vGBqdOLYD4yKFv0wqIxwuk
a84vOcC1mOJfiAkO0It1AeKBn8aqnEx9U43Ja9zDdxXvmCKOQAaGXxBDGbdeihpWoJ+6FI321LZ6
gAK8IkBnSHGup+1KRg4NYdKa/TnjLQhFK88fPE3F2Nmt162czPUC2RcsNU3StdMaIXcMPSpyznDh
IaA9RcGFhpR9syIi61Tn0TZdMe5Sx6leQJs8GvDHoJiJHBtSxXj5O9jkq1go5VqDT3uyFKvTtUo/
WqRDZUW0N2nVyQPP+bW/82/oCTUem2dyAg6ju1kRMPnJL756cu/1mu82KK6Tgm7y0IE8WimeJvsY
7uQzxNXH/S9+MsOH7nUWviyb2uHSSWVg9NUM+bG9ZfWs2BjVJorO13QXlcQUluUwqH9uKSb9CyN0
vQnyuafRye8hSIv/mRA19GKPiFki3J5AZYofRnseNNux8X1ZsJHx3PSWS2lyrmo+ZQpb3eBQNap9
O0j0VPV51uKPfkDFKESyg1zMv1MPKaxJ3pTGeeyw9gvWec48WEM+YCFMKyUeTYUgg8MN21eEQEjh
UMjobTGW8FSOP2hjPGAq9hlwi90uFI5Zm+WWfd+0/laB0Zfk+K+o8UxlBeEHDbHtUa17E5jEB9zu
kDt/49zvDReagvwE7tFJyUjBUtmKSbkNJRgJX8a6aIyukoVWr9kloUloaTbI6kwbwrD6G9hT1vkD
CZCVLuKw0U4/Sc4uG9gfVbb98/Tm7qZbcz0N6qxa+vf5LPfu3hnH8jMgXppxf4X987H/71iAKsfK
6RJLjlO4se5gofnuh26xttficU7nJy5AQPvXRwvRovnEN0bcsOpbfblx+zWhWBls8T4gH1SZxIaT
4Xa4r9P7Fi2f2Nt3CgzqDGzHRL+akCsSoVKGX0sjFJcmR00ky5dZP+6XkG7wJ/oAJDQ4QRDfApzM
tu5pZ869rYQ9/m1DMf6u+Py47vTXpm0rUVQF6fQEZ2bNkozTOs7IwaOuIYOq5jrHcMOtpN2jDy6R
9xSGBFgjgC8/hYVfiIvQEk8e4CN0SEQgIfSAv14RavRTLN/nE7t1TQpc91StnCLg4MQHyjqEHbl7
8shGCw+whdspVHuKL3JnNJSLvxp9/38CTpy0+lR9BVPD1T6A0t1jiSU4sKXondrdLwsOferyfU5Q
UU2EGqY5aI+TN7/UJfxiz+5VVPSUaoYDIUeU2TQFUiJDUv98PC3XKX/faJviDJr/SEXrz3nfWRK3
5csUReBS7oS2RohkvAXXHIpanM9psq8nKH9b0Cf2ouwc8LzQREsrGPNlpCwx98WBCde8qFhW6VK0
nc8cTzB4qRtfGQr2BeWRtuHEt3o4cb3QCFKVyAXO1S77DWzqG/lbfUag3ZIxwF5hLAkBhv7EcbxK
MyX1WH2LSvGtbXMMqCNU0Gsr7QkTtkKjAlgTDKk1y28wAIf2oViHWNGkfw21d5232t4BgF5DI1no
L0O+JCJhnuA2rHVfOkY+dCUMSvkowT3So6BwScBNXUECYY/wAWifrcDJWPG7Jwm311adOReatvo4
NMhVRzEBFse1/V2EawCIKZqf5HkpGs4C7c8hTzls6Ou6uzyti0NlYmlXStDgKchtzYD5ghykVNi0
gm2Am5zyFY1M4xI/fRWQeT29Xjh/ADufSGKm5h2Jgqeui3AmFvf32MDHlcuFc/JOPjJWtbfqwCbv
l4Ecz/IeyoKhrlwsCAEtdCOe8CUeOcUpGY1UPsA0VB0dFqv68c5Hcb5hiF5daihkf0PbQ3+sZR3c
MfTXl1zli0NzjrDIrfsNmIWkeFTB2d+BlLPrD4xhzfmQTwsTFPT1ios0GIKvl0HfDgtaoPZT7QIH
XcHuqmNdy/u90BcW0rRYlg0LtswfjfgE1bZc0lmA978sF8yyOyYaV8fqsJxWfTS8Uc+8KeJdxhlL
IrXVjxPS0pxl9DYjClzD2cgoXXjJX4806iGmZ7zddPe48x9SKExkH7WpaOzce+JctQqCZgakYqIB
mWqMIOV6zrlMbZKATqZOHVmicbkvST3arvw7Wqc7gXxjOyqD8/5K4VsCh0+HPsvL20HLNi4bolGU
x1z6rESm/IknlowUk9rCWMq4ITKSHqNN5A0GG1RMQA5F0fFGPBdnDvrA2KVOvDKE3bNh569ASUIf
mVWlYlc/h/qgxJOotWkBQTc4uLbW5sMwB9esPOdNUTuz4nuaxV5bQUOVaH/V3iD/fHMSyoh9AcWG
2iu1bbwQUdxRKQKL8awSnws92P9JNKJjBu8AgsqMA2PmlcwLtQl/0o0CSPPEJmefp5wH8WcdIX2N
npAz/pVcAjGUkc77A6i7zFbU9jLwDQFFWAmS/07NyfYv0ZXDA7qyOmTruygjOAOlcJID4fzR2MRJ
SNr7DOd365AiCNOE7or8jM3xP6sSSJk/24aL9pwjyoQARmpmbo8CeJ9Jd3JO+8pmc9+OncdKeSVL
vTLRwqVzJHsgT0m89N67SxTTXMYF3VTdj/6CC5p91xOH0HbmsoHfkIq+dOWWe34q19taRR3uQpZk
ofNtF/O0C0cJc+eSEbls7/N5CjB1XBIEx+l2XDnZ+7J1S+OyjtSwTlZlPojydXtSfXyUzi6D1j7L
WoH9ACbcCPnLsqE30M13XIy6NLLaV5BdOgLrikizLnEGtkRZGMlBnnb2Qjiu+NnI2xZeMaQn9viH
7sVNuU5UQ9ZFVU/U7AiE3PcKJgcBv+/zQpuZswnF1Lgmn7w55m5bQAzT5CKJ56073VrqKyx5XrzD
XKOVUEB/IOyTNw55sDJxxI1VvM9I7a2R4QE3ec1/2vYfe7WtqseAIdVLr5IoM76D42ZcBxVAEbD9
8iXjLAhq5z+lp0P1qSLJjQhwftYevTFPTR30MQ7VXdqKPF87ZLeCN3nfTWIblItLqDNBXmMYpgXe
g5MyOQXUA2vX2exDJtV4JpMTnVeyMt5A8Mx0XQD1MX+h/kDxOBog1tOqDSBTtkkK8qLXKJvoPlaZ
WytHamcv/uwZNFmWLZ//aIBnwYVF0ToWWwBwhZ9r1WUYJs+lZeFYkCCDtM8gYJzuhJBfpB4P4Np9
z9z+toY31hb9iUbrDyuI/h5q0H27t9r50l2PWSbGqlzA9lM64z4UQ29QlvVW3cG+ylUFkzMvY575
9Vk2k445Q4mqr1jQ2E8cA1rpMiPwSmalSSn3c6nU0GiajWsFiS8x7aPU0lY70wWcR8jLMF4auS1w
CCfvM6pb+/p9tl0+IQqjWwDq+ugk3MdnDhKyb7c4H8CiZU1YJHl4x/r7t0KwTnYMIicBisQqEBSt
T58F3oIu862fbCNueXhZEj3a3FlG6McFNioU5oQVO83CXkcbnT2rL5qr50slhNp25R/CKWiKR5jy
XK+tCnTo2WJgG30yJHaQxF/LuzEOg+xYs+Z77NKBJl+wYR1SjEJ0nO5ssrJdGPwNz7MJ2owmgbkV
FvZQToY9SQyScA2gqBl6a7+SsYIfTw66DcCFnaoRbdwPXSooh6Lcjg+bFpcRLDFLfESRrpnN9KGu
cAjUXToulsrvAH4tnY6H8sbjDOtoXq+kFQsLfmtPhcse6F6Aq1PoTtCGIN/d9NGMdKoSfMIvPKSj
R3ColMkBCHXkthKCdMJ12PaaUcVpqXcc1QAG/ob0l7kHXUotaM6gwhHU6NZvtgyp8gwHRSbS8zsv
sS/04qgprA1ceUS50C1locX2QPBCxm95YWGscmhVJu65XQ+pVQ9nz7TXXJaoweoGOd2t1c0zDz1s
87YTjEFUf8sFFhJIIN6XJ1bYKv5czwjLj2BjcnMvImOV30YRIUpa18x6cbgFu5X4myVUmloLBZL1
PpMRxY1PZXrQUSBVw3kVX1ZZczaBO9FTNekoYJK0yaAYGvFdv0jS0fWEma/bQ7PXcY8JsJRNaSx7
xmrM87x5G9lrUUNBDK5FsM9quP5ou9Nwur3fxqqJ09Uaims89l1giZtU4qW/4Iaw9kgw09CyN+87
r7p7kytUMfXioSdWH/wjGbGYXI++F3yAP3A3xmGkyRddArrJI1gKGFc5Bj7QD/04fWCNdLnI4pcL
4ZSfz4bEE2cAufgxwRDdGQw8+gg+4Tf3tn02afr5NdyuV3ofdTyZEmWdgs5Dsdp70L0znAfvYpGW
FcQmQx28LpR+NtyoGsc4CRC2kqUZ2wJpzPVwiZyEBckLAImYQM/ruXprvjKQNzbrvEw4Apn3Fw2L
pKIDlthzE1YRXOeOzDZ5EEPOz+U+YETG5LP7y6HCpy0a2ix+1HiStX65Z9iff/B5OQI2UEKGpDBH
OJdG3Ioaww6imwYvUbWLILcYklX8EwbR9jv0XnASJbGHqP2QH2EzIXr0lnl04bmGShHA7AKPaox7
NlkZRoUrcgD6Bk2IgIE26wnrMo2zzPc0HBm/0azoUp80rgInC94Qj3u8aLoGx+Mh2muXLHzEWUT9
iRmDVsOvcp7pP+KCntCxP+NvU4gqxCVS6Dg93cbyf+kWJapluQZ5HUA037rHB1Uw5Vd+alb/3RDs
Q1+Ul+Iirglr7h6ei3ifHrqviVElsMEQb9quc0K7CCIE7UWvIUX+utoUReHQ0nAYghlCrpx6PnBz
A39lKlQuLJj15Cufo6Ite7+3XBV8PbMNJNOT9QXdo9yJCwToondRkm9rgu/vqsMuQ8aus5nMq/n5
aLMItCmJNCb0sJEd5VU2MzBeXC2zi2TJMBsL+I096lCdxB7nsfhEqKTyHVUj/2DEa6pbYOr7sUcn
o9j3dC3TDShOBYSHByO1zMSJJFqaCrRotwHusMvS9WtwM7tp6IOm5numGexS/0Cpuscms9m2dcgz
4tcxMN8rw1a+G+krCwwV0/IxtpleSiZFRIkSi2jlxX/ajGAAbVLlPVC3qH/yxq5txPuDY9LCJjT0
hNKvSrbPE+qzDjw2/ZDdtZ1dMo3IttGjZAwrcKgaIoy3FJbAqAbEvCmT/9tNhXwzifVhIQ30WW3P
ILXJ1j/ifT1UcvejJCxPNfCqOzA0MDD3rnK4pucQkspCiSQbInIg8OR2k6eFpC4zhxu4yBd6qlCd
GcrwrRxIG5rzZycPuIPBduM/XuVdb75WfLNmILSIEk4OAhEkgN6U4Cmi4ys6X7bPM9OzXKY2e9hW
XKyhSMxjr2I145ywcdQUjq47kE8wNEpKhsBKbpBFYHf0E4zYvMnrrch1WGkXhmH3w1/plv6wSsvE
eeTsHpw3SqyGr9ZLN2koYv40bIDTn9h8lB0lPwdxNlagWmS30FlW9DLpX8U5gYZbhnsaqe+KJV6a
KY3TWhiS1L7/MOGdWllM1rBdF+RXr7qDjjL9KO0Vzbrens87P9nXBnMWRtLmFX4koOxJISVD1cHB
8svfiiWB+ieutETxop4YQVEywC/Ly3It9yWSbcvoB3zdEnmnEPYIM9jw40lUo21YOweYh+Woaw+8
EBj5dSYUexuZ6J5HSiIUvIpKh/e6b6CLjR/etb28V4hVu0iRUzx7j17Kdz/scok3i1c8bM7toASQ
ru27G9OSRMvyrhiOHVbw0D82NaEply1d4rOSVi1t8gqpOYFFA085kcs5cTgXFR1JgYWMzgSRJHQu
1xA/6oJ7kyh25t/m8ujBgmKIweBBZaUEX8uHa7CDnCzYAV8OuUDm/IBg5KS/Ve/DdkMq8iH5LnI0
66MDUEKpjq/JshcEc9MDjyz7/curCHtIIbhJLM0VwLNONUfBSDDeH1cWPeippB2ARKt1Q3Oqevpz
g6bSUlz3p5E4Hk28KusAdBL0KPCiK0oFHRB8fBYM/yWXgjCOhlLQ5MkrNKel6D0/6i679z9dJK6u
GhHWjkNIPNeCi+FuooLXu2yKz3n1jlfYBZOjNkq9Tm/fakNgH+VEGwUtWmOVGlFBgvfuThQjbX6E
rX2m3npiKhiqBeiDZsSbLCkaROKpv7B8brDzspJPj76dIY3fHpfzcOlsDw3gGVuHjnBh5EM+Y4N2
xBt94PM2AoVLNbq53ww/eY8r6cU/Id8lI6iH+tYaF0OxdDkPJniZsBWsC3Aph0r691TSJJ4RK8uh
DQuiicNTEljtuK7gqKw/tz/wHvfVwvmVZ6O9QsYn13X3j9/KImrNJtzrsCzGMF/uB32+zXzxukJU
jExXnKx/tlonkIfpgb+t/yndgpq+oeJGd86aJ21kNCU5qEfM3fjySgOVJ6hBTxY/BLJNb6d497y4
dwmNJliIMq7SiIeHRvJJBv+C+9qj8xtSiQgorIECKMI1t084UaFtlJ1RuSNAwnhXBOkY/fCx005P
faVLbIQjS0Mw6PePYj46U0BGLAZG8fr1/+O+KuBSbFaOopibhvi7r35m29a1ciTq5sZk9O1amQtw
ZT3bIJQgXetsBNLW4/jbKhjNRjAmO0mb29rEsaavcu6zGcMlxhljhC3nwr3lANhl6qznE1/lI7cb
y7BYWQG1IPmhQG489wssn2r33mhsoyb+LRP7R9Ve0t/aH9PupDW47wBCP+qGblsDF4DO0ZnsLOdg
OrrsO0PBuuMPZsfNoTezZN8rzflNvzO760In7YK9OaqUYdJ4w9micUyPYLOC8N9FZ1ngviSG8X9l
+ok4k8hC1F36+g9oVHBrc5XFpaMUvie/Pf1/rHuS0PG4X7GeKdQjQmdfPI0aqBIkbh3PdNueUGBX
TZCN+ncm9fYDw5vCwo/rClbUEZMAt9s6NCaNU+cnCnDPAkPSvYcCejL5xDysTWxYodKcmXYBYPBk
/wvWTpKRVsQjosat+CEyzqPTXnt9Q54rU6XUTsFK4r3EBnPT0zgz0vy/kJPAWOBGjl7xChuvF48k
wLzVbjeRoHkSCE96MfbwVERnY94XrnkmRSBo/FsN5e4iI4jcOYxLozyKZ9I9oa7+IpnudOnJ3JKJ
5zQRw/AZFIIbTvxKJ8Jsq8M24LiinU64DzmmzIvpzdhnKLD+7dPnXu/MTIyzp1yEPcFvu3erDdYL
l6Te4AQr8YNVNfvC+WKrXV9WXS+ye6Rx82fBs9M0Ilqo19xaXNrV3+MqoDzHdfoFoK2GOPj2Q09X
8tGUsTyACsTIY3iWqpdQVxa+09IGzQOFjuaZIGtE4rKZvJfvNEms8wb3m+k27IE2g35JqI/E9Rv7
Y1O1Cd8x+qBRIH55OJd3ARoiuZRjkDKhQFwF1pgY1KDPC+5oAiu6kc1MxigqfIkKQXUK1jkN/dCX
IK31yIfbx7VkNnd81kChmq5cii9X/h1muylvWQymgUK1FDNx0FJhVdgYCTGktytyQ4qNJB1GvgxF
x2blu/fUMKJkBpUQ6CFIEnyjBPWHrfrZ7xhRqxnIs1RlTEljatMziU1zxyqfHehYR/2MlV7xkEZF
upULNjkykzxuCuQcR26U9YXJ99OcQI5lk4ypyBVCpmsr4VtjtDF3LZn4/d7wT/ICghAfhyOh/k1i
Tsya2YgOWPg61GEK/BqfKyDTzuoiisYTubkUNb89pNGeJpAZ1xM3xnKHDgv0/2hGXqI66snjZ4+y
A229j/6+OsmiiZ0uJcvyk42wcVmLAHQ7cKs9VaE7Hfsgm0JY9Fkyp0W56Q00wvAo93pPpUYNxyLB
hmtIkyykihIiI1Bn2jHh3tiHqlbn1+X94GMvyxQWpyWiB5En8Cgeuz5WiX8x8wOsZprN2FefAy4M
vdDd53BwXcVrNfnPiVFawYH2uroSBD2pYRbONjBV0/RAGzZh/jOxb9J8dE4bpCwSRLyCHIUvcNG/
QbM68ldMT4xHLjwZMnSwGwri9RDfrFWsUzoyPYr6rPU2QQs2TSOn4ltYszXJPM8tAQH6y5v/QMOz
/FnUJGKpX+Ysx5oqRVCK/nfwo+ZQJMfwlSDo2CTqEbgxX7/TJuvzlJe2J5I+UUYD0YxgIFjUgquf
XW6zhmZfHDnXro/VKK7N8sgSG5nPcpUY6ow0GWaauFYiHGlbjTBd/CL0EC69bfDX+xoWuKYM1CdI
TPGQ2L9QKGukptykOd0EjIhOJXdEWEqdSFxIAuKMMsAdKw3j00qiLBVW+3chcTXBiZPln4Y94Yoc
+W640GsAItXDjZ3DwewDKcc2qfVT7FkUHsHrhP+quBIIIvxHwnB6Y1lLOS0CqwDcZ7xWM/RuK8tL
3Iv1BVaIk2blzO6O4bPAQGD6poTG9k1YjhQpqWzesYQ+EKuGrTRkbWS5Jxfpec1ohAqip/TDiCwD
UE3OTPj9lh3+dVC/x/15VRRxJTk55SvPciVatjDOQPlTyA6tB5LLco61P6HETCGPvIJCy/rFzUjl
J5pf2izUil3i/fKbhAADEm2ligzjr7g/YsYLosWEdtlEgf07XW0sc7HGciK6QxqqfeiqYGqeeifO
RCCbmx2fTlCINU0QI+6jyEe0SSlciVf6Wbk9Ht5zm45wUrMgIjGat3BIDLYGdcFpnEaF+anQ4W3R
n2kuVXmo28mY7Ha2u1TywibgtetdDXGV6X7viTOLQGnm4JkwSDTMXJg5KlGk4JYg5DhGAkRb1vrJ
ZJxdBKbAWRkatHKRbC1RYXuZcAiCic1+Ralqj/N08FBPUd49w8A24NhwGPdtCZs9HpnqrQRtmOFX
VlLcrEjPzyxi02shqfFX8HV9CdFxdbgssXnpQ0wViquIH8VTngOyeksjnSI2jDLdHKRaUOIunSph
2QTZLNRX9TKnyWvy2hnIVPgjUcyU+UFdwOGayiy5/sNmUSd6d8y6MkuUWCeE+GbRTOZN6t8y/5cL
rBdXXJux9Hy71GS8l7TJEO9vsVQicf8aNy6GXFDtGI8g+Hp0uqwWYAi6z4Gevdc2t0jaIVcqxEIj
Xrkrhcx9E/1dzWdyp/P9b8jHtEgrxShBtyUOa4zJVZnpd7h3as3FpBCspHb6VFUKIDDlmzRYa0H9
gCOquLHvxGpNbCwn+c6g64mLlfXyMRdxV3TIP6jBLq9r/7nbnnorg0Ly30JN7FxgU8KJoiTQdCbY
adlwr/W4QDaWVaD3YSsYxEof+Gro8/s0dPA2mtmUsaIGS1zwjGwae7InRhBtaIJvsVHvZFU7ao9N
pEO5vO3sh5g60kKw21pp8uWgD6sk+Pd8uORJ0j2qanTGWkr490kgMN4P6dUtCxFL70YxB6FOBHqS
hXwvUDUANCVPK3PurCmYHgwBTQkujyOJyF5LtXprOIxtgMouudavpT1t048ZWUMOu+5lPSZHmaqh
gVZDdOO+6+T870a1L69hW82zyVGUK9W95ox+dnd9Z/vTNWBMorczeLX1gVJPVB6TA/JC5nZ0jG0/
NYgRwOJANvisn9fyEVyJCaEmY01Jhj4y6UdyrrCc1uTaBLcEJHCjAu3ZUSGpEE185CLxDfJpCS+L
XAalCvICYI55a5pVXFqVXC7OSfOIqeoTjob7KbQJ6HyrbuiTUp8p928WOzYG+efF5joBoyxM1yMF
1+Qe+F6Th9YQ5dyeB1EzK7Iag3wOO8kwyPMS1vbhyv8cn1ZvyfVEIaqKmt5s1f6iv9mQOPtiS/cq
mrdmHSX26+6QfrRdmHFxlUQXXMG9shCgHIKyqjg3of2CfuA6eTYvV109Ae6mTEZjU3wf03WAxsZH
ZoZZxdlcjbKN2RKWmKmDkb0BxeHDlPtxvHm1scKWEFaoTRHdXRwuKoq9FL5O86jR7ENjyLIIeLJa
R0ZhpyBfKycfIDurinJEvjOdqxhUBAzEgblg0X045vBpbBruL2KEpsDW7Ttu1GH7Zo1QRcENWMz9
UmJRg0KiwAbQA0QjTXTCMM83E37E0tUpAYf0JZawyPpf7xmXcyn2mnKJjH1LtRB6RK4fTIRbLP8r
Hb2fB9zYv4xqS/ecXhX4nvg+NUw/LooDyA3Ds7HOPT0BkSuB+fBmR+3FIUOVk3eG82RMnx/tg3X5
vds1hIGJwhvvI82hLt7MFHxpGbWJ6cuQ59ekVVnFH14MXnnwRsw8oYcBKEEMOCEJRAo++bYUVWCb
W0JWAM0KxXatDT5v2JyFSjc0pYVzNXdEQnIPtUWOGKXZokJPdh+XsPyep1fwgtkY4y7gG/90rG+y
L76YYASoSVl9lWNaVUyXQr98yGRrWVTXJ0RKxWviMiinXZZrlcpRpI76EcgXN1nW/4GrOBvMlprL
I4eai/pdGsamPAxVAwyRKjl5Bh2f7gtUtWrJ+GX+i4A02WxUsuvdcx5pvCogHcSlVdWFZfUcYkko
C4wQKs1Zc730rVaGsnx9yof5b320XMpR0kdIL2GxMOZlMZck6DIB6TYm/Le0apd9Wirbm6CP2X/7
1g881F3LjMTfQEyhswO5BY3xrKLxqmjoqWxuCBLW4SbseUJtOtOoEj+BjK+A8apRLqbbPI4yqwMP
Kn+QfmBANL0hbN41Yt4k350uJ4ohk/IjTec++YBgYQKO5ZeMEmUfzsqqPtqrGlRc4BdnTlcd+E+x
PzqxvWdWKGSTpqusMTa2eZF5e7eGzMb7zD5KijH1QD/qxTzmNj3MB5lxaBlmHqRpHcTpSGuXS+VQ
Eob+ZrQC/NeM6gDt2WTQZHQnSzjOKlt1quQZj2QQSuYjyhlm372TtsvZ227GHHi+4zF2iOw8F7rs
QWQHrYbwKZdTPejCNeHDBhErx1yeea7BPiewnJ1aWkfwzlhzPub/VJzmjbz4mM2NNWy1KMgnEA21
H1FqFho/7fiJHh7D/EGk/sYn1ocWG5xNDBlgkX83bHvQiti7Ws08BqyI1+/2pb0YG68+HlXA4nzu
NxjRhr2JcowUE2Y81kXUo5nckQ5fpCwJssxmcIvXP1B9xsuBKd4aU6d66mTiX+0hdOw+6batzIvr
JkaNb9B4zbgBCy9O/fO6lVAr0TsehXE0mA8MW389DswbCO9FuWubiSZBL4Gne+WhGDFTeSVjiDjL
tCWDL8w9R3vNfHtKRHlzFRPQKa29dlJ+kOd6G49ix3LWFZViECXulBKsH7mhd9tm6UKkh3k+ZV/2
tP8tMH3O6++Swig/aF4V9VZDJYGtvlgGlYw6DWcp3drK5jADwMesaA0V/XXpaYzu/+wblb4XIqGq
38G2FpwtYc0cecMyyOwkXmHUfjDTWlInudUXmGgfuYLvjLw351ROEE9EN4FFLbiQE4kvPoNXxwMP
BF2mHPAGyS34+qDqsB/hwGm+KWeeDboEcignb6v8zp4WoyMcM3IENLrsWMk8FR4OSQCd/KYqSv/f
bvvAbwqPEYJcX6r9Y5XFT8Tevm0pOJB4Yac+Qo51JUU0k8xkyv1HSfQ7w7p8LbVLF9M5Jo3GDd5N
Eapn+KbpyiD6ssIzpjmktJxuuVXHdm3stoJrFYB2jnKHpYtFpBdDGExMuexZGTgAlDTS3HWgWvBb
bKRsoQ6RdL65LkrsajZFJ7Y7YFZ/oitLfQs0Yd5TktTJm2TyVwO1PTiYXP9004XimDATgcOjIrN0
z/CIr5at5kFmoQa/EhhfogvrO5XJ1zotGWeKCQOEeoSw/jSsbTjlha87afIaeE0Vf16PvUk0j9kA
m8E7c5FNGiPF6tdit8lH8qfhSW209oRAWP1oznGueSK6BXtkTtZwBjOU7Gw5QeNx6bIMDwxdmqxp
GgG8ekIojf/3f672XV0JfTdj2FeeOtpw+60uvQXU6vPf0jqpK+d3Apb+Yt2VTDoOSO6Mir1F4eSw
dNYUyeRgt5Uk/QVoa8nZdHf+SRt/KDJI7dmkDYKsVTC1W+j21Xlsc1B0WfPPe5OU53h3wFVrp0Oc
nleUJP2RZHALTWCpftQKMXFXme2W7rIasBpWp8iBff8woYX0O5nBAwBbskUJIz5ob2nUmtVIYOgy
fhhLaw+tPA6r8GeQWZ3hwMUAp85acdiJcgFHTtudxRyIcNhx0r+YKcJzCcSdy53/zlpv+SCK1gq1
I+ZpCoElAea2SDw53oXJ+l6gGrzlsRV8cmPp259UXqT4RD0kfZguJucHr06dpZIPmsE1dM+c6W8f
/6xjNcBzWn46FKfhbYab0aE9G39nF0iWwKihC4DMGVR6yrdC0b8q1ztwHAfWXJfulJ+7GqbiDHfN
2lZI8rloOjHS/sAPz5PZdHFDnI16GBMMeIMuZWB7I16jRN5UON0X3hzk1Pq+/O62hJiUalR8JhNf
Jvxyvitpnra1cvXvqTwZuwTXouj/OUt8MlkvZsAk6R5t7Er30oDj9GUM7sM0RLSpQCwNkj7ezx1J
cPXtxRGIonNdAY9Z9WaChS+RpmdyduqPGjXLzBWPCiMtEDD0Z48UjjlwJnHozKmCN0RJh1cw6D2q
7f0aGht5yFbG4Apy7NIxwrQgz+luSVvr+J0smFL/FHm9ektMnsTLFDFHpVwCn+Xkeb3JVEhTtr9/
4Xb2gAzs7uERG/FqzA08UYSTCbfBIwM1P/dknGzrRscGSYpGLA56Dj2+oacfVtIWc/5Ly5Os8fvm
Vcd8nEBxI9XH6gMCjeywVrqltFNSa0eD9Xlhhhc7+1SDAw0mhC44AlK5J3PdiIn6laL49rlIBrWY
cyQHWx85GQi3uDN18q7etEO8mH6WaqZVjVQUL/SmIMQBW1ji8rof6Yx6bHXBnmHNzLo2TKgb4zGJ
xqjIwMlANVD5snwhg1Kt5BjpIfV0t44vebHjBYKVUVCCzZmknMftdnpDs+vTkC4kLCupk0QOyuY4
eUnkSbwLk+o0HcUp4UYibY+t5EKJThgxCDtk3LAERar/6My/cJisMi5ABhl74ZIU48Jy3JlnLus0
ewLb6lAp2Bbnk+3MIgwibqdaAEwwITnHcZsmc5pdg6/PuPH7DcoKA1sN0W9LW7DgKhXZ2BMXfJog
HoCFWc1T4Zmp6PWR1suP1T05ksRi4CLmaSdooKJWccBlbk+8b+AwNR3S8M8ALEHtZluohztZUO8U
IQAhGV5viQbm0e/JUQn2W0dDcUYeGQ6UNZaSs+eEOXBlxhSfiTD4srskf9tyQZXUtjwa6Cqkg+Zv
tg8EbBsMS5c6ZUPQS7GWPbUAyfdoualrlvwz42iwsGULY0sIhTxd3R8aRwReUZy8DatNtzaxOc4y
btuhalnvR+vhS/IRsucxoqEJrk8R3j+qZyr40pG3oMq8W9v+1CbWrlVzHF3Z1/MW0EXZu31RcMPa
vuzd0H+rSv8FgpU52G52jOSzU0e83wm85PH0mRwcZyZs83ChcQvMGj7ko+Wk86aSMIh36CrnUmJy
soWjJ3aYbCMwXcLk5ZHcJfMqnC2GWCyNz8JUxkyHBlB2bHjs/e/XaSOVumB7wY7dVc3LHhpWtX71
AnN0v+DCPWOHzH3vRLeUMRv0sI1SILkV3fwZO9mRDgQzPnweU1r/CBLF05QLNIOUy9Nm5sfICOSI
Sw4/QSKtVJTPhYIWl6srnec+mcw0jNSSinx2IAbhmD4jSiWdkaRmBE8auVD9SEJ0eKQbfzmXNXMx
nSKHSXVClN6PbAtz4ukYRQonfOd1IdCwOtYvBUTkH/d6vGm7qxVCkqalQVso5NBfC8hEeGYCUFmK
U+PVV84jJ+lPaYYecQtVbzucegvJvKP2Aw8dbzjuQ/BoiTR9FXAIhRw/a5xGg3MaKJB930uIMM//
sWxQbty3y7R9IrLE1/cUEa+R7RgfgEwVO6Kfdv0hsZH+wGZQ7vJgN+Dtk7EXi9b4H88phWF1gXC9
6V3oCib9A+R1kphsp/ZaDXRhErvii9KiOdCs0YTjiolbgGzXxVZ22K1KcedoHjW9IvCt2rWEpZE6
oH6rekH42t3Xsi03Q19AXsFn7puHnksXSrBhCU1LmJAXft2IYQ33NWc1nWUkL42UXflmBzwplFFy
nyKVN4OT5ASqG0CFC2YnmEVXONXV8NNnjEkUf10QLUXPE6lQUDURi0v+A71xpJ3x+RF8vjZmO58D
PGtdN0sZhpytz+Pnc8Srsoloab9bc5KpYkoT/apyIMU4mFhbgPZWcgegvYZILRU/GVM6ZFj4olHn
qEHtOGy+iN6LJ8TZMiCdyBUf8ltHPegxaqLFmysXXx5iopxnhCBRAYmGpyuOkSCS1iMpkvXgvbCY
EIxIkUtBzC8snU87LIVen8n+Xj1Pw8jtLvCHyFhw0l4RizDFp2TZyRufJF2/HTmukg5MyURg/5bE
ytTT05mgD2g044GJx663t4+cZHioOkzgOn2EQL55kj5sDYwvQ9k/ZjZ2OzldvfF8M8Zui/Kmr3Lr
xuI/xBUXPNr3w0DpKgzXhYXxm9ozhswzC6vVpJzeNNIFJZszuJIkkKfURPAtkCgjiv61b9yOVeY7
5WSSqT+SGJUvy4oBCAatgWbp+DTCSSx/I3WzNIF/VFGP8MiPlnpQFWPIfK3mbb4xDrq7oyErcssJ
1icX2ArfHIVoVQBMkxOOXp/ZjRBIVRQ7hGDARt1K7PZNWGOcUbrPhvIF7s2JrVBlm3HrTrB1jAgj
DJFnW7Z+Ycj8QohWM7vJ2JPAxEIRpw66+FcU46ctW5PhJ53216loIvB3YGkWynqkaiUZatZXTqmw
ZXhtKdtj1VE7F2zGNy618j4GBQlNJfwTQQlochdqqXM5XGvZoCBkgnf4I7gZ6EdNiU4oVPBd8wrd
5i7i2ly3ctG7qL+E4JBA/7L2leZ8Ir7QrmIKjBsQzLtSBosOwtjmBE0d1oUb9wWCcLVME8gBmFKm
VNWsv43PzCiW5x+hwcvn/nf5sRW02buAo8F0/FIl3jeEU1KSKGcG693E0Sewx3lesf81rN0nIiN9
33lXVTJlnkbnfHvd7MhYi4bLIccirf0efbVUzb/BUtr8zhFknt+62EHPPB2rgpN+JPbhs1vrDDW2
/dPLFuQAzH7Q2H90h8h7zmj+dBCl4TH7340pUDxgrvmLZkXxfMk/rHpSiNxwTyK41egnhmoIPr40
LBG+Q28xKhTfu5oJZhVJWYLRlDBRbtixGhBS3tRruuSLXqWY8VqN8bCzBxRpPaytHUrPfZKl+mdh
sE+M0HvOYEY4WInry9TvFmuldpcGPSidIAWFeusheNHjjRtJ92PAZXz1E/Vd4TjL/dMvq6NsmhOu
jCErVab7mzf5ZMWhi450c9kVknVkJPzAFUwiPeyuOMOX4p6TY8tdbtGB4sWUgN4gi2jihoxWY3e9
gxrDlHELMeHYl0OMgRlIb5FgVfr37pTKuh60DF4pAFFJ4GKT3dyeYX6jNxukygW6IfwdGDkdfr6z
Jih/hBIwJ+0eIk1YtcQMu7G2BoFhcP+8f3PEGs0/dmkxaGffxmFuo1nHzoUSLQ+1I8q5CSwMiaue
dSinueGvmOu8lqbwG7cUqRauPxAj35xHeesTnJEBVvNyca4ZRF3dERkrbzJv/i2S67J34ufSMVUK
3BDRel5AA6C9//S8WepoICkVf01k6eA1MzlqvgvhduFfi25/UnxnmDoLq+GkQ7NB9PhbO+sprBH0
Qz2x2itmIaK4rR/rycnNKBsJKPSPCq7R1aIvEn34INzRwWO+JmI8X82edz/IRbFBhcKUY1zzrr19
MifFkxh6p4rwgA+ldZpKJ+kNfbZVn2wBi1LB+LKlpedFPgyuENv2+0NJnHGj8ZdwErpSksqrnzBN
AMRQ9iYy2hYTrg6XTi8WuP2RnVUkEnkxd5H0Zft0JCe+5wnnQ5Oo5GkKhDzNYpYATQqrUEr93UP2
NognCeAlvrWdjzx3RhMgNCAvzZG7CO78CUP8KCqjBrztqA3NhiFcoxEbzUqHUxiCoYjSZk6XCBJO
pmbpNie/BHXDFzHkTh7F1ypvJK+KOWor2swTO4/SokEOws0qDtySin8SBBb6Qd/VYMgU1RaKwHAF
9eUhXdGmOgnJQIvxFnSezqV/8W025QAco/OdK6TtiQVMVubKcesag4OUN/Y0PK38o54HM2jPt+iu
M2kDDdsrwskrmQNYSmUszbUfOLtS28PFbnHNIhSwiGQu6jSLeth/a/ILdRgN0/2LrOVbezoEAgxd
jdcSx++mPbjBIo4VTh+bayBfa4Fs9EB8bSi7GyCIpxLSV/tQrMDbTVocuQO5il1Nxq54Ymb/64XX
GggZHhWnYhwig/WGNsR6cNvsn/QC0U/KoVpnNzXK0p8qj2D73VDvgmN7XrAjHzRJpGldkrJ2Uisn
Jol/9fgRzxG7YTVjm/3YbETHYwplAOrFzsz5aU1qan9JlU+hf9eyHF9HzUAB5s4mPMj7afzqCV/y
mt6gRrXo6iQkTA8nZ3csU0A02OLqjNAOhxMgNKU4lnwEzp75zIFvkt8Y6qahtMRNaDLmyXsJKhQG
5hBEGI3qWqiLr9RVXoUgcX55y5q6+1ChodgCHbGqp3rRkvu564sFpKKQpCtLw4C0DIJ+1wLNjY0I
Zv1aZh3ix1CxUfbnoSy3Yvh2eV0XeHfPj/EEgvbMRDeuH5/xchqWrK2ChlHz4Zh9tczc9ZM4Nro7
sHl4fyDNsV1Aj+fVjk9X5LivuefB85xwgJ6lGWbvDkIjf+FFfBBMTANdsCeM0PaV95R5bYV1+H0n
NmSlmY49+prUVLzJmG64aKgCQL5KL9hsGS4eVbFXxWAjXkq3jcxrndlScn0sy5eAmg+y6NGzVVM0
TOBubSb0WYPtyCbHLWeIx3NuFSHL2vwpjwMPNcMbE7pYUWwqZ8pWq7cdRWkOKq6k5kI4ZrUepcxl
wWlcA/jcYutUHrJiaG3WmUMlGA1QTOCmrDRoxhwSHHDnQVb5XhWCd8/9F+STKT+uxAIoOxPNPtWD
+zwEe9bBSQHshiD8k7xvB02jH6TZfkvgdGyWPvkXXU7FnxuydAhec1D4NfVqf6p3wupBmXMSnCnZ
5jcGa0fmXvFDaaa+6DBhtBZH6pnxp49k0vzYEhVgzOtc0zR8zWSYvaMl5qEB39geOgPQMk8NS34N
jfIAlZIBJ+eu4LU+PqUFeR9uH9qBmr2b9WBFXCw8v6STnd5+YlcOwBz07GHDDayag4eu6BnWXRoS
uddchqpG/nMyON+kIaH67iEoPStaamj2hxECvvohvJ2SiiQZunjYe7MPegtiiBYl4K++v3BK5J1Y
ko4pcqO/y+rYxngzAsljoF9ZI8MtzvNh7wsHHJ6JgTwA3jo8ko/fAV0KQqY4Qm1xnrn24r23cF7z
pXrp9zpic07ShGtog5RrhK+xCjN91Jjg1ryzkWx9GgsPrWd1OehSOX4EvMYshcmS02aoqjxKiUO5
PwWoxJXfO4lKEqeVlDAeN+MlQ/kGe6g51rZMsPw8KvGJDFkY0Q3jvz2014A2TOVkTYQNcbAWwaaj
XPxfGTdUZ/d3O7LhMuTND1+rEbmgyO8pY2JoIE5Wec2WLiKBAcehIU8gZpd6EFQ9iaEYy9SV1w7V
GKhKC9w/EGA2JeZPWLN8VOj/eREUZL7FkwwI7Sqc09qT+diQCq+uQWJxX8ZREGedn+ZTypU3BA5s
E6JgjEs+qpBkJUcmPWrl0frjCeEoouWTz+bkPfNSLs6iLmWWtjj9/6CJTk3uiSsHYq8ioVxva+yO
NvzFUd2GoL1s1nJXenpKSj94GnYb1hlvVVO+uZ5du7qsWkUWttxCxztF9zfVCwi4sLdZL+z672jf
FnqQY+GsMjBABe7v9xvoXZHCsfIv20do3GydRklLkUjbM7cbW2dcK6vbEYDRxKPYDxpstBYErtSI
gNnhNqkqNVoxeHoikAFP0guhdw81g2pbLDCpvoKtiZaGObX57rVObdBP89X4CVIG7cV6eYg9F7yW
jB7lDTWZk6Ij6Sb3NOh8l+0i3lu0qPfPMUxpgXuoQMtUhSH8nDx4KbemLOEnJsH+rpk5rDo9Huvx
Am2awLqd2UFZZg/fswF778JGO3zlBOiytlWU7SS+YtDUGXOozJUk5KjTZ6bpBbcQOlyVUUuwMxYb
s7cQOuYYqwSiHmERjavEWZAcxoTCxhmc/iPk5HXmAtlIay/sVWu1Q76U8ZePaD8vzRC/DmLHoD0T
dVqKPCBXg+LWA9KM/tCUWEmy9WpXvdS3lBFhSdvgQq5XNXevXeCFqYfQpdUGCb5zVL/l3zz7A2sK
OBXh6O2lMPnxVw3MYwM2suDuZvEU1+YcbG7f02n6dMlqMAY3Xh5ggezUZn3dLcRkfgQ+ofSfGCk0
oSYjHI77FOOtLBYhQzjgT6OttcP97ZCN48q+4qc8Lw928R1vcISBY1mSZtiNCfSUonpVdfUm3Y7F
YwxJCberIT0dxI9x9iTAeLrVXg3uHexdy8/QshOkJFAQ2QRv4wn94XHgLAa/oaTx7c0x3Cxa9Z3x
p+cHNDLgSmhUfCRrPqDHo24rUH6J07AGAZM8Nw/a9A6RKKqw6p9P7O3cvod1Jo3VLze8Hpp+SwwY
uuIk5xeujkVvHW3rgf8klkv/cIr04UI82nGS/Y3sQuoPzcVY+Jq06CmxyhiuN0twiq8IxGWq7oqE
gCiAKNO/z7a4GhKvaWuLeJd2vce0FuvWBJXfLOEh77Ayjn4UYm/380VuBoVg0LfIEzoWzW5vwMAB
k/4s2/znRVBxEXdG1cBEWz1lp232wfpxpxkNBxBjzCiKIUJz6RRYoBJ0MaEnS4bDqe8KK56ROJwv
oFS/gMU1X+9ZuYZ7LCzZf+zby7L/CqHPN+ii5X0HMTICXo5YJJU1dog4xxSG/8wx0Vt1OK6oCDXI
BuouTvum0EWP6Mx/prar4XK21PiE1aY3IpsiCFStISpCADg5aJxYqDmTRnyAzfiX8ehvfIXErFnA
Hjkq3ROrWSoptCIRHvkZ0Dhxkym901ehWcB9uCbUvUZExBa7OWKFYkljYfqqohIGopQU4ehcT9+3
70dLqqbq/PjQypyUkNlMbaF0YT2iFuTTMndUhdPvR9TsR9mZKfZ787j3uju6gsPEtj02h60Edehy
f2nxoV/1mSV8KGUYpG4pucUolX+qsWA1XXVMPjy9SL41XojMeuNf6CsaOHkF03U4/2P3KR8BQVhU
2xxQCoDSpYxto/hDOPvU9IKlDiRjRF5Ous4oG+3mAeeo9lL1fJIH5JDkxfw6cBJ6C9/icS6r30i+
SfbAvJQ1he2GM9+j9HO4X5cQ40zJkUOpZTwCx5zC+zHp1n3nLyTDHG3S5AMI44XmEjwUVq6aUK4l
uzsQfTpQaURYz5RdQuyB03Au+RTzjTovOjSXafEUEdkSYoLkYt9pjyl7vTQzCo6yVxEpr1q5afBp
icRSYHqgOQDc8uaMBBV1SObXbSm1ORF2ajv9MVaJMZCRxXc+GOapjjEHrnX6rU6UUfp2WFT4zdNk
Mt6Elecb73fTPeNe/ni65XRKmfP0MzzxoWUqjnjZJPfZbWhdxa+oznTDqUHTKXaI1Bnj+Uv1rUGn
O+WfnbSkVtQWHnA190uG5rznsuu77YYLEyTapUzWFE0e11L+iTSImQjFCeAWX79V6tLRN4n5Kllo
jMlHeGyny0kZhu0TYu+JnLI4w/2T5sgyjjGE+LR1EQ2Kz657rYT6ZE2rPfZnKNaEVMMe+++15eEi
kvM/8au2++ok98xCYBX5RyOjUvLeEW18Ww3UvXi+wkQrrA0IdaDI6NFxYiQ7sLL2NoIMV8e8IwZh
JH2eZTUQHElKS+5jyoUgt5x9Z5hUp+Bu1Bdg1yGUqAn+WgQh6Taxm7Ek4INNBjJ8EGuQz77tklec
KtiA/tDk3qRgy5vHz+J1KFX3SVku4y1nlzay/Xz+/9qdc+T4Tgzli2a3kNm+YMpGGz+yGpyqGAKV
5IlY48M3wm3YZPjwvK0mst9ztQ2FOSppeI7YFtFPcGfwDOip/PBtHeVvZXYuTV5gzJ2zSNcLFLtM
TAO7syee8sGDFFVuAe3FNjnJd8or0FBE9XtaST33Xw8QzWAO1dzDT4wAFvsmZFDd3ti0tQjJAqVD
tRQXAI/oY2jmLkR2rMtVRnHBHfkNMioQbQSfIzi+t0kwPoZMlPMd2Sa3owdAeQqZykF+xRKo39lX
nJdbc1bNI6+vHOj8IJ7KcxZ5mHBt1eQKX0CemrT4WwtzpgX+6L0EXbBNb3fCwBOSjxJbaTfFaPGM
0ypYbWFr8hDuRshM8qpdrzWKNvAsGKHgkJ1UOdn12niw4bEhGvXmyf6SWkZb+KeO0HRPpe4r9t4R
c+lDYwO0gYgWgDOBMyUa5n2qyyjJQFvvIvzZJgeSvWhy/NfcsjTu3sbZmQMS1JTFJuV+phEOKrrP
kBlMbknjeIbFBwIz4UvwKvMQTKn2FKLcWbtWnkqLvEdjk8oVksX4jqEo3h/nW6x/xFFMRZDUuj/L
+hWo3k892VppIO9qEhR9CwZf8ogV27wOqcxNY+9HecwvZ1GAHOXeFukSRP3KoR+h+AjCb2QkWW2W
we+lnBVQnrQhCiR8Lr18M1u+OLlNPEkfFLI9rXFGvBgVCPwzzmpTXiVL/5XoUyP05FxNOsXD2zJR
DwO6LdmS6EEuuz7PZFWImaJom9R/XxCJlR0NFtTkdx0Su+LI7KVMbnN1mhsGOfORC+M1B1avXfjo
NRi5RdsaIL9O5s0BpR0uPzR73cUsvVK8+uRLN3B6sO2crB5sYIlLY1CRjuqQQWCLE/1zDPKMAaNG
95drPDp7wU4fZ17EHYqBrxuh1kijmPGcHJiidC8dPmNOCl7GkFbxgP2JArXkxl7VQWuxBWUqAmZY
jXWIkV/LJ9M99vdZdE0/SNf1bESJFroABNv9j0fi0bfBhvVbBxdkJ2U1SIG5SqrFHmOnQh37ZeSf
/kg8nCxPP89bvB81+qLKKboyfWJhd9U0lBSDqHxBxQEYVkgmVRsbh/4uKt//BaUKPHjGhnN7iGW9
MOjtpM/7w+V3e703hIoxSzhzOAB7nqZOTL4pjIpKYtYAgsb++LOLaBjKpxESuJXXj26XdCj6VYso
9dZkvPMqj0AuNO2GbQPgBLrFFKSE0ZH2YWZGHpmSiIZiuFn8uIBdo2kfO0fLA+3drEFXuPIurQLc
mwVm36lWVXxvJSfu6/xCyhRuLZyv9tXvFgamvg3UKD6MADSqnLiy/I80p8Ka8Niy3kq+xmD/6KnH
3fU2auEASXScBepfw2IlkzgohGFiiKyfsgmvPGGfa82ID42BNTODasJs2L3G5N75pgCth7nCs5fr
q9eQEtbqug95ZVBgPcggvJAbC+ABW6LuHt6H95ZHvJudMUwAa7U+UcLT+ZrviquvtezYUykf8q3O
yM0an5TZBWQxOKlZva2TvvhqlC658sd8hGaoVPqqnUu4b4GViuB8XlAMq6Th9PiXGc9tC2xJOrO6
lhEAJtAP+XeY8P36MkSyKcxiiRms26DK1uq54GnIEaS12P6FEVo0ILDso5RyiXboDzX0d+r7N8gC
HOtrBXC/I0tl0H/k5G1D0WK8ZjBknJxkA7TpL/PIYNsS7tTTUcEDzDhAuY8YrfukrsY0B7P2sWej
S89hOat+meOp+Y0dPKiq1bISfDvnPw18drAbzTLPDxgCG298m+yHM0UyE0B5Q0X8NMYDMdCiXSDK
nezMKA0kkEtYARjxrrOUiiXgXpWto0hJ2r6+tebykddr3mZpaOfMWQfxbGsWPpoE5DFp2PktQQsV
3fmFytbwow6CZJrL+0inEJNbBbz72XDnGSeUbrJnw93dQ0AMuZ9x08mmgfC/M7vOO1N8L85XIOvl
m5EdzDnx4cXw39KuKsLmT+J9wNX3njA5RVROdyyxZ/o/LyqRKeZyB5UOtc+K0ggy1Fv2FT5jT/+w
HF5lMwGgzrG3gEbyZnLNZyWS02iUVPuxMGw+tYUbbhGsiZyfv+PT9SohOucn3waMZli0bCnUM6th
S2W6sVxpxc88lvkW7b3Mx9n6tSpLnJO+S2tqDyVE3JW4JOLJrtqtgHcAdIhwqSh+/Dgj2M8NEh2b
PnHYBuDUsp71eIxSDPerx0YsrWhNvC6xcs2dKwINsnen5P0rK2vHx0JnY66ijzZ+h00zbCeCyC5O
WUX5+b21fFAR9dE2QRANoNjobgwFLtK957Vy4UgjVCnK0+pwHUNJE+8LYh5aa3Z2CgN1EK5q2PXJ
IPLEGFnoMQJWb4JPCMp2jdRVjeZaAS/TSl9kv2dvgctgIpEqpD6aUqxWnrweZ8JUgtpxwNk11pMC
Q8qp6om3Yfce/orMAkS3u+P/YAzwp2/KMECv4ruBuh1CpYbTtwFxfWo5+fME5yhxwIBuvFI7vm4R
kYUdaPDnS8aqzoKCxZCEq5TkJrmGzujcws84NYlebfzI7cCzS4KM7Ic9peZnjsfcu93A1i0OGpKo
k6qDVg/2qiXGcU2Uz37Och0nDr2rsAjCyDaVcpYYZtSjcMLk97N0HlNOczrng8E1OEQUFnrE2Sck
uodmBod8Bs64KRyxUk/SRqSavVu8EOl3h/MXFGSqssFXnLLCcvk9t037ywR0NYfjh/RnAypmACTT
Jpopk5+5zI3JS8YF391UjTu4jlapB8Nvb1xrCARKGo5/BIOBAbnHkBa4XXutzkXUp28XB5uQbGaI
ansh2d6f0UmXlKMw6Gutq/Pa7CmiguN+UnAvCCUEsiolGBIIDN7qx0TrZlI+TFj9ZZKxQ62wLJc/
lugqg21H+sIZ5qfVGrIhg2XkuxfvNR21CQbJ+IgUnjF8YWI45hnhBQHxd7B0NvN8IT0TlzysO/HD
h1tJCGbN8BBLvaIFbuXl4VxbKyxx9gfvuPxKMqLf6/MPwdUu3RAJsHgCVmSEI1oe4FiLI+3ursQM
RKJUVP0LZUK8EbidMGsIlYVNfQmL0hFH88KUCkJW5g7GkS/kLLqBevuhjz2w2MeuWYrIj0zHCkDE
4IJsv+3wzFK2gwkWOVpdXjwX+7WXF+0yDvbq1k+Q3zuDymvvzIi8QiMjXYWzatqsKtZ5chfAvFqO
0plnP9cB0pkXwAJkq3hNAUUBfT8o8mNTa+6RUTKdwxj7TG7csjx5puSUlPBx6CSfDHqifwaj+051
PLFEKkiZKKcjcqweTa+gJZ0d27LKQXEsn0x6hFW1z14WNlvTLrSTkC/OPvJVX4LWJ3YLTjuhfNcm
0TyYyNYiGzptNY4HUl2Q5oKyxe3R+mT4GNPpokTxDIN7GHuEY6s+JmO+DWwHS8R444h9hDQL5kcZ
9xnkfbLJEToAH9LNvZF1sce4eTNu8V8Ap8v6ivQSkc66tpBUae7swLYw59OZZA+EtN4D8zuSK8Aw
pFI+chczYAEwqCv3P/lMTg7sIgvtPMZjgdZsYWBX4w1fB3kIAv76QOxBpYzA/9dW5KDpqptdGewJ
vkbCwducc9WHEgsXJy69HTLNoOf2H06z1FbVJwkUPghTOXz9iG+oAX1kzndgjtZaHS4nspe5QF6k
KmQECoNDaN5A4/59z3zioYWybLnUbec41yO0qOzHAth1EQTJBpMfz+aqN2UFJiy11SG/ImV+qD8/
J/tl4afIdxE7uPdCxHcrvIrI3CF0oncQT6yVT6pd7r9w98yjZsBVC0z6brsTYdTJBTjShF9+PGDt
ytNrLr6kiIB6iWwPEsW31LI63JeRHVGgubXNLtXb9uGhxBMlQ0WWuCUEs8vWHyLfseTtvZNoKuGZ
7T1tEgFZNbJbQiV4/X57WWHZ5buMBK5B2DqXCw1k70VNG73PFvvh4kbYw3XU1J8mFWNscwS1C0hH
3Q50jvKp9nacZ5WggOmRbd9t98IibtqR7l4lCvYeylOrdapmlshmvaky1BhrZ55AOZTmAzLF4HGQ
3icGgcxJfMuwkV/eeQyuL+XPz1kNY1CdmPwZhH15bqc6iEIDNBvdQoP+wKTXL4t0k+pKVlpm9HLG
H6OTUhkBSR/rPtpP4N5SdQ/y9Rc8kVH0xv7/zth3xz4WOylOX3WZgnzkBz9ErO3O81dYj4ivMdgh
XCxW+Be5jdRAVxh0HslmW9lfZSMhPB7qk2HYX7bHsF8cR/iJpYjUqnaageXoF8ATeqiTMBpEk5He
eYqGU+mNdL66V5+OdsqZwF/O7t07ZqhhfVU16UGN0fqz5OQ6XK/9G97Za+djUqgnGpQACZdnWeT/
AIovjC4wQXdnzSNUBUlgmbi82SChdGGfcOJYTgNCsWT7RVp1xwjvsGCDBpNCVhLC991vAoOLHdwK
4kDHgm0WUUk6l8c5IiNWzow84Vl4rv0W1RfNCZWEUR/eWBB0VQHXqBbB6+L9e322OgmA5+ZWkmGF
jdY/kOyMVHEa6h7ZIRGAY8NQXPjfu2HEBA4d/zFqQBjEIPn4Pl1YhoaRwJjzwqNJEMiDOsbgNOPu
+v0lBVh7HD2vQcGCap69zEb/VjrLeS5Xl5U+9t6TS1ikY1oIacPlY9WWJOqQ1xacEyX/Phsj8D2J
VgCg13TDGQ/9PHLW92Myi+j+LmRb4g7lphWCSWlY7oF5FonAlD6G4bo+uJ3c6q3S4JjAfrMRmjmN
8E97AJDhonieZ9NpX8f+i9qq/Rcfx5VFI+66Cuf5OOD1jzmF4t/Sc251f9DGkASKs6yhHIyNtZXx
2h0gVjje8vhy/gmwkHV9bMImTuD6Rkwu+/fewybjY1hF07h96ujXByp2CH8dMDCtNLPu0sT9fgvc
/IyAGooqQtpkNq1xaYnyYmb+5GMwg6Wm56gYzLJC9sUhb/IpmecH3Ms7fIWFFtAwIt7gohUjXmud
ms2XdcZzv5npNvXddSl4R66x04IWkAB1F+hOBi3majiLrWsrGBjjeg7m7fKbGtYlWzcT5bTbNd2u
ITQcQYK0lENNvay3MUY8ZLtxWiWQ++Inu8qYPORKncmezj11T4YZUYEK17bHxKQGZmuPHxag/yfM
isAg9bF9L2vF5I9tiK5w1IxCeuCq6P5kDp6aOjf3dR95MCEzTmP5a2s6ToaLhnkoZdeogo06lJEI
TnL0TTI4Z/PvjgXmDKUoYT0GWGkRlJTJWNDMaf7MIzp57Cvoxo/ab0TvlBEKfwNB/km9h/nmqCoT
EAj1vCBhWjjnLOdiO2mXBq7F4B638gerK0XdO3sxvri9xrhmUeaBAYqrV2tHBo3v+0lf+Nqf7mKK
GAVkakQX7rnh5R8PtTGDbke3+9p0r9wT6X1/XtWX/YC5WPV22aQqI2trG+MzZ7wNrA1rwhE2F6We
BAifK1sSxDMfmV0NqzXs1yMPzWJ6k+PjIZtmYIYgaplxn+LeuFupfJuNfyoUR/9K4ifjNnhyrqqk
YxYntIgjVUQVxdmfK8vwBhet/eHiXaxfi4/sqTzN1FMUrUyf/igyBN70XgxiMXB/bXVi1cN33UMm
FRRoIxPCnqJ7eCLkpvRb8oJMW5Z456wBBZc28Et6g8HLp02Cr9VpUc8SGibnFGVACvDoMS7Xa1Ro
jvUS1gmMmssmdshszGYcA1Yfn1bg//21Qvi7xg4oR6QZfYOTcBz0jnQs3qWa0N+4eBL+XwBu70DM
v/g21yOevBqirYP8K/MYsw1clJ6qZotD5InPXBx+0eADYpsf57ZjyxIQCiG5zl29MPjSuDzXSJtR
QD8suLB6qxAC3B7mVJw9/fRaPb+EXfA+LmlUhgXNSQl+BkwYVHNci5A/TlQqj9/m342kNhVR8Osc
GfjvqUHg3OSWfsjra5fvL+rjcZXMZse2NStE64Qyc/2RjwQ4OLXlqdbgUfOZB4Xx/yumjSQ30bEY
cIsZEJPM9isCzWPrG1nbXjNqVl13V9ee0Biz+6TJNkNyq7vPePhpw9XF/2ssY2Y1HZiBVZmGeNqU
DS0hT6tXbu7KZw6mTFJwvfGJgNpgSV3g3iasv5d1CsJbX2fY0QTUiOYo6etPEaTuD0V3ImcURl12
sjmT8WWxbB+Bkw8uVgHRkXPKfVb2EqCpXde6WNxS0nprMqGnriM9v1CIWFFMN8krZ4NC1iIwUDKD
qGAoCwljmkHT1Ux+VeEMejeQLWKw3q/kJpaDfBRJaYRuPpE0Bwxhq6GKpWBpkuJ7b/f1HZCs4n7P
d19OgFAy7MFn1lwibAkqb91yBX9XyzpBwKcA274T3MnJkdQS+LEuwZJ/s6efOvkICpLwIWpbvz48
UL6GZImA4A789TEi7CBnpJuBpJZ7m3WzlKA17OjOcH1RHXq7rPzVD/W6L/ODffhgvgvZ2XLXYUx5
tRUz8tUEkIiZ/3I9pZg5rD4CtNvYpNMR624qzqCjbUWeXbLtqxXF4y8mdm8wH1Q6h2tu3PNpzLoS
g1j3pPvrBVMF5hSfk82I0sm/W9flPm+VdIxZdT8PD9+mzzzykMH+Vrxsjc8kZqkUhgiTCJlkGUHM
kQKkLRzoEtT2e85VgBMLM+q8rSuc5vilFa2b+u+X49NFvZzTQfyzKKK4pJaY5Zn62/gEoBna5I1a
AqHdmwHLaJbRK3yPXUwvU/zteTl/aJUS+IfB7pnHfJnwKQfOVRP/SkClb05h3TKmAE7+5roPqT6r
wqRAnyjQcZnDY/wp+MODivDg6fTzGx32Eeqf2ClrWXWtVYa939zaHeIJFK/e5eJ5Jc+Uq2pFf3zj
uoJjjGhXeVLPhLpL7fVrWlxxWg0fVGnFxQE2gZof2JGmljlB/AUhDPgBGR51ZvQ4/TEjM2QDPuOX
VZ8AyTJvM3wDV4PEh0tJw9h2bN+qz7Kjpj9JWW4wX/SN/sYELlzBDhIfJ9nnnSIHRAxyYhE5OgbG
fhgwuZqJtT4pcxVgp82R/o5fgcYzZrDV2BZ72W+BCWsqjBXlRw8nYuoZF9bsgf27qUuoXKpzqkKh
EL8gGtqadRQTHu+Hod5diSoknlejaUs2KyRD5lgrRC8L3ibDf1k1adkhEPpAXXaqMpl3yMt/hXSy
izfUilMY/reEywjj2oxCFxyGKcKunGb+2Sd9xqTvJ3mX0i4BmA3aoYH3SHzzcRa8OD9g6dTUYFME
rKfuG+PQcueZWo6o0m7MB7rhIm/6mxxbgCZFdZeMCmnx4YbA5EkneoZ2J3v6sfQXr9LokS5PTIuu
jO8d2HYKH0EE68y11GYiPGdTJas/s+A/EvhtultI6RTzY8GbWTlsd4dHyaZhUJSjqgoLk82VkWEl
Vwz+Sa9GBkV2cj4Mie31FX4hXHwBX78H041/Jmcw48YKcvLK4NXo6x0Y+50eBO1SAbfOraE0kKnG
qj3MwVSP+Q2IvHhw03Ux31oeyIrgiv58L2qxjbbdt0+XFr6YD4Ar03xht5ErVzNuBWxecyn6L9ba
tL8UFuNQbgVNS+8NNbOd/Q66mPXgWRwifUvn0H+V5JbuGSZp15afIKkKB7pbrRcTevR3Ln7M+HwK
SY9m+UtFeUlaQPJjNYVZgVH2L/YbenGy1HrHAaZ+XKrEUtJu5fPRyrztGS9WWYe5voHif5bGdbvB
7M6gdWsKWgYwBxhzebf7a2OxUJ6DZqXBjbkWPwQtjlLgKzQ5QIirzZFq/g0WTGlW9fxpQfAiDHP+
xuzM5yyP7krm/irJSFdaZGiSLt/KvYI6zkmVZcZPnBY4H7X6C6aRSBMoexk1/Zz/uxTWg/SarR+I
5GqO+Ooxh/TtRH0LuMsFkPRm70iNf8qKjv7ftcEXlftQpeVeWOMpi09BWLfOb11adtiHeQijZ4US
+a/w2BLfbJDac4QQSGrhNlA2NFV3JzU/jO5ZHONU3r4WdFQ96abHP8zjVGdB+nepeu7TxpXIdSnU
h+nXby72syGQl94PFhZhLHvHHLA/vKiW033bLqFKwempekBBNDlohzuyfPDCilGSSQ2Uo2wPr7EC
7hqfm/lWhNdLe1/tPt2onkX93h8c3crvClIM0SwDON4uOzE7cwFXChuI9ywwf6QJQrepYCiPZr6U
+wIcMMLJQteuLdvNnrgh5KU3CaQuRQjL/2qQ2jHvOkdsFkYdNoWeLVNLGMylK/vq+3xLheQVledZ
OVv6OfDdMKEcMfKIWUWRWKoLRgypi4nQVfIfpCpkUrEfZJcDxS0m+Ti6EayQrL//dLgrElaxfPjH
ZeYzIItqLScelgx+Bq2qX6XDjc0YPAB9Jc6+90Ck2tdqObmQfs3+ccRc/VPxuK2FKCw5QyXenCke
QJqqC2tBUny9iqztrs2U37P3YurTpvhBU2aJ7BSegDjun+ykMr/pTNdZmBdVdH55YjguyULHt4uk
NmQZ4huuPAlg6WIgBvAi8tIf9L023qK9Bzp7/QGvwqdhkwmld7HfmQKoGWfrleYzRA38FicTmBa9
g23tlDRgcCIeVD5/3qYolawCRQ4XPtXOkX5UsbiFuiPBqih/v6/wnfIf/53sJYUU3tXN7yyBo735
mXzFj6vYrQbIMEssQvzEtsKnyuwAMpBSIZuJrEZfRvVmk/GY7QT12JRuMkLuZHaZQGcOhOi3AJnX
XjvULcZ6Z+zs75Rqz11zaHiXP2A8xtGYs9jv5BRhYm+wrjTS6B/n6pV2mv6AwGZ3oZfTGbr4Tqn0
Z0xwhCPNEYtSeF3zXkY50DX7Se0kEEAsx7NYlVOJw1ecUiVfUjQrTrfWfHzeSXPR+PlByQKJX/Tt
kgidglJqnLgdxgsuTH+ic3N9Nb5EyLgiYv1V+kDO3dDa1lotUViGVl7WqxaY5rPpoPPWuBIKXBO6
F5zVpx359JAwzl11BUdacPnO3P2DQmPQUVw8MjIlNJafnXm/nzg9ly7z6AZvb0luLfyqLlnn/4BW
0n4l0awMI0dNCZH76N4ezWdI0uOIhohyo274AgDmqgoLawLj8OhFuhpEb/VnzYkRdJASSGGNcj/O
qXWSc/I/WZlU2gCK/VJHulsye8a9r8AqswnsCSjvWTILhPqxLTqkDEDJ6d/QG8vYxaLJWNa9C/eF
0DRW2OZtStv1+9QDyrnhdWrhJEBi1nE0oJ5ewE/L6ueYo1yEWTMI9JkfFVCyQurtQdQMPGn56XZ/
c+JH/plCZ9fEkPyXi1ZJPgpLBd9BZUWtNk5abHM3IbCo9mvVZy7O6gPYrACUWah2Cqe8DcABJygC
iCA2F3RORUlzc1ygk5YbjkPgqLt7QXpS0FG5DXI1/OovK/swrOMgDq217S6y352YqRCQ0y/ckPEF
+yzUamRCFu1v3fCwm36YpRhyj/ah+PzSHCGZZWZrluT6DPfl2csYNd8aCRy/BxixBgZb3muol/QG
9/odf6oQcoS+xIhfJDbGefEO+wKu2cyOElinKN5Euwh+sHfR0q8U5lbv7uLlSMq7eCKHRw7ZScoP
OmeZsGaOR1hmmb6/ZxFY8Idt9TASwwhaSsoTpLHVhJZRUnEL3DxrGqO4jf9cky4QuulPDhiGHc+J
sc/5hwyK42WYNzCmeYWCm0qElhAtXZZX8hrHz4rzYdVoD39nLDUZ95iFARoNyL/ntb+xJ/Y59r+S
DsnJSu/PK769nZRSl1FwgqDAq07J5sx9awDoLO5cSp+EbaxdnPXWadFHCFI2M7XtkDlR+ooQFc2C
XbbdO8qEoZrNQTz7qWyWuIuIVIZVUlsc60Ka2+LuYSXf2wikrMQais6AxiUah157WCEhJP8EyhMV
hUcSCJD6x/51NFz7u5J7nsyiDyMEgoNaLCFx+nJUdcJIwoLIh14UPEEDYGL3OciOEb4jwxtyicPI
OmhIfO+7Kx4KDrI/C+8M28ejAiZKykpFcipKNXr9cXVyi2m+QvbSjyH/9fvWAtVxyR3jWoRGYfaI
JPAz6QcrF70sUGe9bz/C71uEXRA5c3aT233unj+VVbhmsgqNaXUzsTMbnPzI1zyMrai5vhhI+TGi
7CsQAywpM2T5SI9Z/E8cWq37pymis81T6ev3PW1y0DOz5fTVXsIAWlvdP2EYAqXCqAYfg7QMsFLX
G2KwRIzHjm7XbZKEl/y2lqiBqS+Chbh4lA389Zkd22eXjUBnSq8EJdsLaUOrrHDCXI50JEvZGa4S
U/UNBpEUZ6VRBW8pDNRGzjn6rrVs+9rNAP3ZeYpueySZL6bWbYcpb599sNNps6MAsr8wqWPY43Z2
mOhCWTK4DjwbBvOVVtXysJXc3frLiXhQtZu+HZob4fxGAc4DsWxippl3LVpBFgItZLybNUtDcbV5
SMRzycry7E7/aCHL1QLn6/MwruLDYGcyzI642rEWN+QKIE2YBLLig++0i4X59plE1FTyK9shAOTV
Ih/EGwkZtKNVJzzvq4JEuvegPntbBZw6aaRe9gbAscviqVUOS0bTbX0kS0HTnbsB67eFyzF0tPTJ
zpP3MWb9HeItiXTGcJcFlt8mkxMgHcbbz3bR3RfM1h3GbAYusXOeUNqJY8ku4D4WiNwnGlAcDpop
2Rm/tn7WkbKLj2mDTB/QXPwrzBOyXTY4YjB0YSqo2KBeVLLbGt19BRQPRhaETMoYqK8d9RfVNwCH
XatQz1QbJa6aNxY8ipA0eh212KMqtvqRFvc5aykgFOpHVyrRVcSi6m1TjyHB4PL7bT3HtsgdBwrG
67ntZZBQek2CF0GBXczQPBUIkXZrGnD1IAaQlr2gFSG97Y3g6Yb3WK51L0vVeL1MiNNwGCdtj3xf
faJDA6YUJdM6MmzU5GPPo9Jh6D7SS/SpFqg6Tszpv4F77dU2ES+m2aNrLSoX+RDYqfV2VEIQ551m
QdFuNCl6dTOcZVznh4Y6XfESxIZDTi685hjSbl3IkQ9ptKBP3NQpw0MPViz30ckTQ/uXDOwL2TV3
5jt209CHev4KWOHZ/gP5eZ807mnJrRZlTlKjsFMfa6ujfb1+3X0YB30EF1p4CapCutJLQZ2ylqwi
R/OBcFYJozi35WlwAFb6Pkt2wJz9WdIcr1YyZcis+iIGIqtBwnB3Uqf3X9ezHamVJoDg5/goMn0Q
We2laqnOUpkS+AScTt9QD6BIpwcAGQhNEJuuuqOhh+TwC0jngLh15zxV3/AozqTkcULZqdIE3Mm+
NW6zHreaDjUril3hWMp467JNFK7lnjrSmrDDg6t9TiVTRLKAR8wLqpehnd7G10LHTGAzcB03YiHm
TGC0F/s+69QqaCL6wUX2tDb7n6+4ODhFs8sE0Ma/lTwPaHjF5WVy0pMXEeRMY1yoj42Jly3ncT+7
RaKlt2b6acJHmTADdzIpVzI/iPe8m/kkIXdCk52I0LxM6wvI/N8NnPSKatmq4XSVQ0rz8yZQ2qQm
3tYztpmo86re1OSAZCJrWFRYt7y3jNcNKOMK6JsFyW+hJcDIf9W73UxCGiuDrcz2u8VPtpCAXH6q
ncd7Cs3JoesFJvk4txHxzfHgijcZ8femfuwO812coVp/1Vs3efNU/KVKq/FjAjsOPxtRIn4QxMI/
UcE3Wj+VRhRaqpdpxxdhjcO69T/fAyWp6OmbK8LQPxDSJDv/QnBMfEQRCncJqSAs/C0fcePAP6DE
kBmWL1/lyDhEGFCE++a0PTQz/gnK+rh/KzxHhLUWSy1cJxrp4zPpCw5vNz4IdI1ejhvv2YaYU1Ay
/JwtrYqRzVa4MYwwDdJ73/eiRtbtILLNcl8o6z9RaWOxlgKtJZ6bC1SUf+YB7GHFTacTYciGVw6H
vf9ktJvpWSMtlGrH9KJkHsL//tV5t3QpURXuPkbRBIC5Pxz64wgHGGyCUyLk8L7iu1BMREzIbYcU
N8Zg1ycHjQS50PBzaTJn0PxXyp8A5xHcE56vnQTSIUvZCKFNIXNrBJGQCW85Ur7Uwai1QmQfpQr3
yVdg6X7afX1HlWZsOZkRvYqwG+xV1QlViWdRybByMtWu2Gi26/AzjgtOCgWBYHhOChRBtiI0k5c0
ciUs3bkKosoIf+nU8Z5lVY8of6NHqNa2FdsoIuccTqODq13kn3wDZwzFPANwOCFqUY6AWw2EzPbD
86WHX5iJfVjYysf1qHekCOWLlIG4NiUI9fD/7aZL3paNflCu67cdm7ty374VHumvXbUpFE5dNiSd
U6kTRJ5ONd9mP3QiWyBXBfcqsClJVxcckml8HMB4DyT+jPxVxtZv4SArfRLFS2EeWqa2nxeDGeAM
lF6H6oR1OcqSLeYboDtfE3Tv9+CApPNaLy0kiGN+ov9V+8rxVIS6hRk5VyMtv/qHcZJdu7rJ+RLN
g1p/Mfxy8ljrAwGeEK1xvoHFyCueFGNSCTOx/dtLU653daHnE687mfiQ3XW2fO1uU7Wk8Eic36WM
rjOBN8tX3ZMTv5/5DhYhw7NyPYqsxYvNMJrtrlkzOeIuqsrg6XRTSBgu9KUgyvnzhCWLmFJtq0nc
eC5zTqCHfY+nGShCnzxMry8WF0hJT/jb2ziihtoDs+aDj2dbmTHD9tihSR4fX+9hj5ECzLq97rt7
/X5Jsrgx+hk+kkl4wav+JRfKtbBw8FbC6nDwN9dp1nJzkRCu6cY38OiAws0CIKgrn9QYU75olQe2
GvHrQb46TREqg/Q1SRh8OUb/u4w04El1dJL28PTP1f2AnU2Xj/0s2RcVnWklhslE3qukyUvo4lFG
5q64sZ8b3VHUxpNXrSTFf8JopIO6cT3GWjhBRPOa/GsATtmA4PYq4R9DwmA/bCsPK8AWPA4JhrZG
DzrYZv+U2zoypGzST5/znpp3b9zbToUjbDKWz3z734wDPSh7MPcv2VNR3ZcVgMbh4ckCtDmKPMKl
25/ihCNUTKLN0/mvzC4dgfMQGr+yYJOomcCTL+5sGXs91wr8aFMiw6R9mR8xspIQ+RjdXLD0/rer
Zf7kX/YoIMbkc7r58QodDs776Du4txtTGV+WIbBg2F0CHXOqb6+AlbwItPmtXjqdwDcGFuMb65Wt
d7j4KIRc/h6XMfgjGqWPV8Twl1Jjt4X4bwg2l1rsQn1p/x/bUgPnjzYB1m5iBKptubt8gs8JVZQu
rsXZg/NHHYi7Fqd6Db/TkD1B86Sd5dZHq/WsVXIbWyJx3psx/rmkSeFG7yMlgFUaazqMDTY9tldp
Jbx+IvzK0EoKRwiUjX/BWxEjLLQUX3U4T6eLmCuI77muQbMKm9F2hRNCOU9yAg2UBwB4YDjJilGt
AO6ZAHryywuv2SXiipvl+xbbiU6quL7phyuAs3I4Cg98D4brb0TmhzYQJYIvshYt1FKn5mTi+Dzv
J+qdL+DeXZ8EcjY/ZbsLFAsQF/xcEfYBM/Cs2RtC+MmHWcYs0TfTN4x4RIIwpaOL8CVAyAQoyh0J
qEwwvCe/Y+XLdGGW+TUrQmaYhSq4X52Fsgwn6nOQqXiXbmCIptZJaKDqgXDSWno3mTSx0iCzmiE4
KFBa3g2cTfd9Be0CdfAE95jvm0GNfuU1RQIrkbwS9cLWbiKYNtgHVCyAi2aBZwgtJPehBD+bzKfl
X+438jf+ILoIgPFVVC56Yw/S1cS8znITyOisvXHSPY5gz9/V4WK+IBm31t9XXCdhjMqiM9p2/EsW
mmTeqVO40I6Kywatz8/3P5bgTc4b8ub35zgP31osHVjmxmN7n9MbBven3kTnp2+bcrcfagPixta6
mbIdx0Tkml17rD0F48wgeYH1NySrXwtZOjAVWeDeQPV8PoBDya8mOSXPtCcu9tUnqqo3TDnAzHGZ
KGZTWrhvY1i4R/l9kwjWgtlCKxnrLEtNNRUCTqARFqPf4Fkg/kZwYbLI5WNW+OkZBS3l6pQ89BsG
dxlji2kFBEUubL4d8zMxbfpTDtg0Vj69omwrcbyl0N69yWkuZbg4sTCRtp1igkhjtnqSodT42pHt
m1TdBqidVnqZSMlhpdvfnnv+Ni29iHD4Vhc9b/CLmriJIIBob3Qg6SeTiPMmkFxJUGdspjnvA9s8
VaEuwQ9W5/3EuNuIxhh2Z19jAAXWKdLdzOWzfVHM4uHgqg4ys9rZb1bdJQlAFIxsXYMoPGs6IYfc
7ncELACNI97XEVHCHyabByQRIWPoKSH+PiXkNLyuvBHTPcxvuNfsWCjshL6gIL493n0luGUtN/aB
b48OBhIV5jk+1vdREwoBVlj4I9B0nuWDYGVr5h0JoK6wA3xZ8+7/o4sLHgBb8GhClI5Ggt4w1O2m
qIUyXcH8YCHy1Q5TgIyStvWtSr0UZMuvdNlrdkJ7Glx26w98hXZnkBywbB+qzVXtKVqiWS63BIdi
BIhdaNcZy9Lz/k4OpfC8MD0jc0mS5kS1AXmL5Zdr8IrWVWOnrvpK+O4Kg21q93e6FuShzTAWYuBQ
avupEhZXkB1+NCbtOhfHakuvv5HTg1evLLmsI3zW+H3WsWZu/Kpr+rv5GeGJ2ScFqmBkjVIpHgFF
8gFugRD5BQ/lHJWf/SCqZSWDgbvNJG3WG/kRLd4OJYffTX/jz1B8aSnn1jDQiIjNBzOGbkp9SQMJ
zbqcmw8+8sBIBpNIqH0eMJN1liwNvjX4vYVhm2coSVO5YLH7iVoKCWaqgXnk6bZMtDnEUJ/iCQRt
eWuWrPYdD0R5E6CLYRx3vVbUf9t+UaGI6OwaArQNpQS9+Fg0hW4OYIsO2kgxR8fqMJsIJvq2+e6K
ZjssX3eZmJ2+rrmkMdxC67a1ZIbfxP/GwTEJngauevqiFP1beTQBSFFrFAkKXk6uWkpdW4PEmLjt
/m2q1ydLvbReP3lgbHgE0LcOe9fYF8IUCLNqx5uCTGSwIq/9pcZHS+CprYBoKtXP165KtMujOJ/Q
wthiU41qwBKykQ1KKaEVZF0s9Slp7E6TCV8piWj8Hq3ufhunqRCQpYbpX77ujpt9OI2IgXX8sBla
IbOIA+k09VfBMoPUquaR5ZjK9QzdIGwfN/KNgBZUjNz+vIfIha3xhhl9Ji2lp6wehJ9l75qbJCLC
1IZlLmoANDde4s2UQUFYu8Y+VM4mzpkEI+ycUUdwAph0oftYnN5wFtjd6YeH4swBOBom9A85uGZ7
nro7QzQEUVjv0kDV9WSMgsRAdbIKXcuNG0JN/Ec9F7D1/6Rt5BivNvA1DgZVlhHabF/wFs62XDLx
/faBAXnRLBi3d27n4/Mk1yd9RHgpqbQLtzWMqd6nm+Y6y+NbwImF8YQnlhP/PyeloZxZCbZXr6Nr
9dG264/TXpZqJFH/ZOv7TBnHYC57ZdFuYxYtODeiX2AQifJT660FyC0/KyOda+hn5aIaFrv0qNtY
OQP0EdCGxp4sss6aGqglugwpnTQXAdaKv4S5TX8SIKoLXh1+aDa9Y7CHDawoXridg8B0vTF4CYOP
bSEw05CfdoyuCFMmMBUjJfa/MIXE44Si9yd2gJlDi4SCzPNBpze4np1Kwj71KjzaH4pKY4DDxitB
JhAvYxBDgIFp6K9IevFxECSb8vJ7nistzO7JC96kEqGwukQNbP69F8UaXPU2SRyTxWC2SmHFZc/F
zAkEUKjNafgAnFPkYtsxVujoFqei3/FF0IDXHFKkAA93w3YsTEQW6VLl+G1SLOKs2ilLeWJJELpU
egSNAVFfI6lywhSTUJ3boU23b7/AEEatkE3qOna3Qv3hSzKVQqctUeSOPqnliaQLXikyT8GBM6CY
GQV6sIindCu+JFC60iRG2W7Gx7WOrh9rxMU67LLuiiIgRs2Sg6Dn7UqLbul2eFJHaK7VXc/0n6st
w0uo1ZaHFQrYJ2Ns9BBVe7jf2C8zTQ0B6TF/LdY2RvS8dQYcbPOtgSRupkYuFMYIXE3wXqxCsIhs
iwkejspzE7dpuEzIGQsTb5cb26ZNe9exGTX7myY8PJ9mx5CWL66XQJQHvKYGG+pRKZynG9KhKWHs
9fItgNt7DWFwc92PYv+4kQpOOZ2ik+NvI1BtX/mfENUbuFbMGh9xbahXQR1XcH/TODiGSoQQETaV
TgAbgSnSL5A4n/uWJLR2gdeJipaZZvB09KuHhrFniE6woruoaV9GnjBGNB8mUo3EnWpPzWMl6JeX
as+nntEyKhwvF81+yVI1ZZD8d2bQxqpRORmAfjIPBVKa1iP1/mAzbEF0NheBn4sMTpn+mvHHr7w4
64qUjz/wkKwO/+PSoXFkn9CBhlr+xUB90kzgl18lwT97ctbZ/jhkatOIq4aNvaH3UjINFiqA/UaK
l5BAxgczXibiI048hJDCuDhYjm+I6AGJT+dMCr5VphK7HfX3+NVYMqiDs9s9+HOtCtaizjVoX8H0
kNmSo3O3NcPpXWifIojr6+ma4DSK7NrOMrk0iaPUA6sdRODpAzKhqh3+nfz8ue4C5WeQKOa/9SwH
xjrCnsK9jGVfev5EZBQu3vFjAd1KzY2LJxmnSBuyiD40Nl/wMBUL7LVy6SazV994Tljp7OSACIS+
/YtVd6T7nHkSWbnpO/iGOJAvYdzk+Kb71ApqpjOqANReYdwsGRJFqkMrCvQdLxSYJD3U5ESJmOr2
CwbDDVBBhJrZe+cWD2xatoiEeAhPgQmrkdaKnGoCbqakyi7t2ubT7HqPq+avtHhkdb30N/3uNZvT
h561nAZI/ebhAa/M8ehnlL+4AG7R/VUsho9383moz0fhGw8Z2q/r8aSUK/C4Me/UXwj+ENkjv8+K
m2Rpuc96lT6yrGdSO7IBMpgs7AjHs1cdN9/ClLltWkXZlsI79pi93Nxo4x4WVePCybAlNG6x21Pv
QVQUPHQkbNTVMUxLZjXf2ezn2TwGPNuHuVTJFUHxIuvDGzRBTiwJ8JD3GiBjNsJkYtdnQcKqgEbw
Nz7yo3244D2dDQTIvzIMKqB48053WB8DC262xQe+4z7s59PSvkqIjgC6XHiyRoYwdNE/lRANOcTE
eC/xPh8voa0aGCP1mslKGAQVSV6z+8ztQJwrtBZ0v15RuARb+Ht/0JpiXZZn9BVuyfdU2LeYbEgM
JlAIWZNBSEK4L88MVgzq1NF5HJfvIgU8d1gqNkA9PCT3WCNCUaNcZZblrniNjoKLk5ETlT7W8QwE
qkeD3oHortAuMMDpcivLcRzlmBmP7NZMPVhYpZ2UbV/1wbqpSaaeo4usn+CNR0+goF4E6pkoM8Ez
361Gy6XKoKLosOR5S0l68RnZOozS6oKFyNo4ReFjQHTP8X5Twxw/nofGgOWP9iPElVMw1tR76Q+3
p07igcMotq7UbH2dFrex1d8VfQDyEh/RPd8rZpamPbpzB2z/0TUQp+m83AwwmZUHQoV5k/VTY7y9
Aehzjx0BEsUY0dPr7xsOULRC86U00Gx1JNwGjVkZCPdniaRuQLVbWkvVQCT9anstHkqUf2FYgIZs
+xRiY3zdkHQxg6cIeEO+30yFh2Lxx0nz4NbHqoHL0KNOhj8W/ineX1jRR6NdX0T1Am9VLcjlLBfN
WbrtztS89zrYoCPKGIVUUFDmamiz0JRdUfYX18YWS4RSDAjKAHhvJkjMulFM7SgX6D7+Jqehi3UW
3kXK27xgYC3pHhgHnKNDFRMjIgNB8WMUJorDLJKEyak5CumUEGWop9q2CcbGFw0fnHnd7lLKtVNr
qssTQj9kGoy9F3Av2Pfijpps8+IgRqCKRn4lwXZK6nkotAYqoMEaD6NGcTyXesDNgsk3OmJKQB21
LgqRUOcBYjvAgKmRswADoi4EcxDfmHhdR10wiBGKEM5LAW/EeVqYL6vjtwPpohtw3f6Wdou+LZam
L+2YWZAt15cAD877KXSBwVO4bIO8ymhe+891GGby4G4KxgGih0M2VfA24GN71QGtaQPZbSTOfI2l
xUqteWP/8O3KzVP7VojCGk4I+d4eCE+IyHD8BcBgjn3CSVXliEeoSWl7pXmFsHokTJ/Q50rR9lOn
qVb+/g1XDlyxPAeWo2QK9JgWZ5uEg4ilB8FHpLp5XCktGj1V+EQJioYANho2C+unGjt4+9mz595z
rNgJ7FchTdeal/Y1p5P24EN9l/zChJMTl0a0EICJwMbPddzd+oHzdDyCdw/LB2FmM7QyW+NCj5oM
DR9CAof8AQWjT43PF86BmLilCVsgAU1jmBTWjggRSm+E5LVbgoOJut4tHZhV7kXo6UWHO35qlZr4
tIVM9EhuB6fYL2GGZ4Hc8+mlSTH9iqMrD3uej5bqxttEvxQWl1szDblGMFu1VMSHQt+27yVRT1jl
i3zjNFAxFhmjF0CnPmgswFftR7NN9R8XdYMGd3t8Th1R7nnDZAWSb5vkGqONaMm9qwlY+67CYl9X
Y71UvxXlhCJRlEguGWagAImzV+CXTi1QnhWM7udn0mEa3tmAomsVgbNO0wDxZ9i1nWsA2nz3USjj
au1893PiEceZjYW703VwXJfOTMBWeBxxfX/Ew0APaCFZWplV4Yx7lYcC9cw7FZuZpUyskoU8/WOD
phsbvpdlZf3FTgIXfFgnSaExG7Il/tLFZmVQ3n0Uf/SHFA7vWm986awv817giTFyE1rsXZVDQWT3
RYFZe+kvZnXgF+TjnFYIrVXjUMo4z683iEUK8CMmniutfUXE/XZFCojInrdzvGepyCN3E+pPhYRF
FwCQfH2dT3uMLI4jJKYabH6pO1KEg/r+5M6cxx3C8oH4x0f75fztIjrxKS+MQtSzYSZAeAlY/fgH
8k5oWn8dbdc6kFCsq0iSWnrgB2afpF4j24lf/O6JTMIuCDRLU1qHpPBHxuITgxBAwpxMtUOv02Od
1O+0QmiOuF+yOU1OCZX/YTJMKOCEsEDeDSULCLpOaBljF5CbrB+ITo6o34th22pEz/LuroBykxxV
Qe3c/GQR5gUltq7B9Q5rNAQHU3HW/54+TPVCWWKZlrJ9Zrx+ujON9W738Nlvzy++qnQWxvreTSjx
C5+panedRyiYb32npeiRz82mtikrF3p8tmyWP7cVgBZ1rBc7d600sF6NbcmV/nk2uU0eNxxREyXy
aIusAowHUvCXgyJccO5BmuPmN4OmlOtwFwMzp1VqQYncgdLMbPni/8RMZqbngIHQ5630ea9nFnWt
2gBvDdRH4NDJvA60wCmB3gi2LVc6Y5QuPKYKDfgXP5jjuwgcAQ7GfhNsCO31TJ6Hs+M1VxamoJbb
8XLCyvNowjVHmG/AgtW/nW8fiVVIds36d3tCc/jsaBQcx6r0bTZBguY15Msl41YomFaZtsWZS+DT
bt6/URuUmn5u14ZBPFTdSLAG2RKzv2mAgvyKa22NX31IlJCrlm6jOwlcgy7YJoXM6DVuC+yPqTA8
2T+1/OKSdK7drwp1JALK5WAsEdXXNKvS8AisnxkXsh3rvJ6jS6E3PUdDWdfX+vomln3yWfQEzB/B
SzH0du7ZazV86wUIx19STR6f7/2YL6zhTZtaQOM5rUzOcyZBzJdtnV5Jtf6ROlchLPV5gVsAJ0yD
qSj5yfkUi8XXQ5NFfSU18NH0itHUWfb3hDBa4AghDv3GN306ysbvyasryOCkUDnxwDGbM2sbYN+R
Im9sL7wqBLXK/8RGEshpdsdl0Mm1mcJkHoXqApB/nrjZ5a1exNrppoi/anNm2DHgDSAqeM+SKZiM
9srwdKAoSvYxyRJLaa0AXGvLu8mGL0r6EB7wBZP0wS1DWqEKsF7diTUYsls0Pv/+/168eAPGw4eI
aitGDFfoblvwrUAYuVBAEBCcNma27M+L/h9mK7PZr2wWTZK6geTvwK8kaKrjqb4RPiJLtKaL9oAB
gywYqNe6tk+cIeZl+8VBdHObz3NIoztprzgyp4CaPObPzyJNdBHgJgTJqYXzmaUFF37/F8wMApvJ
+Bg4crAkfjAlNv+EdsbsKoj6Dc2H0szlRFb/O77s+W6yU0jxIXiT/75dUKsbIvLPSq4M5trBbvrW
ILBVe/M4QnFA7cixzZL10CLoVTejmLG6OdeLdSdT3dCsfFvR/rWGWxUVEHNw9Ovnkuzhtg03Lk6y
JEVZLsO3hiaGYPaLyubsZf1EXchixJQ54w+AHIDuHITXGE22jBeaoluQgoKxmcZJ2OiLsU8CBxRo
//U6uDh7ql35MfnnXymrlPol44GmNX8+5tQZe6hQ+noLunSWK3mriM9ZTbvODGnF7Ama/9CyYqHJ
Y64SAp1PXpj8JucZZ0pywo6cs0SYNNHA6oGkQe5wFbMYJ13cC/pZW9AO11+EYopzO9MkCdxnz87t
qKCM14F4v2T3YY34rk+tuqkqtdvXs17bW7vINXvjlrLs4krwHdvjZy6Fr2VWxnQXu4XPeoGin/PW
Pjl+HT7NbICkRG+YTwSiJqPzCkgXT7B3kZAscmqxRQ+WNs5Nhbl4EopHJt8CiUxt9+09pzaf149y
qnWj6j6+5RAdNUezZfCPF08QceLPm2TtAhUdbryh1l0iCDR+Sk3bPNL264bmmFaMroVCHFvC/10t
8sLiQuRH6qNfPM1eMUQVaM1Uf7/ETagn96s4xiPcru/MuCVzGHvSEr6wSrRE2PxwiP10LygBsbKA
Z+2H3bbD3k2EP2cgiI9AoXjHN30FGCwr4d1goVnl9bsvqcx0g1OTZ8QufxKltDVTrzlpqgfbrRfI
kBYkSHHV/R7CtaSU/qX49Xb69ZxjPtdsQh1aM3wN41eqCzQ6dIbq+OTBHR12sCKRR/mEZqzC08Ys
iGhVuawwr2Zg3Yxd22E2Skjy5cTdoY6mcGS7KnEjMGGtxeMzwVwddQgI+E5/WcoQmS4OhxpqvAAx
TblNDmX0StWDkzhBtakzkw97FjhUpMCt+h7oyhZt+Z3IdoeeOjnmbe1I5Z4hqO1DeWJ9Wq37wo+T
FjO2ijE1HWRdTiGN9galTEGMVdeQYbRP31LUcpdGisGcf7cik2mrFoB3Y5zfKfFXNfwxZUDBavv4
2QXNRse7iNAWP+3zP1Sa8JCrCxQ/Kve4Y6Il2lQPjaCihvfib2RYLqWBVRlP6vCVAuX9dxGE48DS
Cu5O+SzAQrCXZtlXa5QjTbWgdU2DKWnR4jNi2AttJadBap8EdBsCmbdnvli+BjG9vW1y9+++Ng4t
e73WpV42HWEt/Jim6okcY7Vt2FPbgtJ5jXWeaNjO9pFLbBLHLVI7XXkYB4vMybuv81ewgBFGJiGj
5xW/AXhfGDjbWl5VxzcXDu/xSOt6Fb4GYpDKfmLblxMw2Bhm3kzhSk5xpgmdFdKzaqmAuQnVYiFJ
Xl2ZJ6Cz4mkoq7t3gLk7cdGeh7iRamnm8AiFlLETRnCDe6izZZz3JCMF1SicT/i0d7esXWLBFWmP
a54+7L46aeQeHN2hwMappnwzX5PTBip1EkG7G0PIOzJq1G2UoByxde2Vmnc0JZq8f3NZQ2Dvw38C
EIiuqC6dA8cbip9bJ4sAJcbcaZGSwD7Qz/tpfkzDBPNvGF9S3MpaKtd+vpNXIW6hlOHcvmxQA8gF
LrAn+yNcolLkiJ8dcd8VIAeOv8Ytd7idI4tGIathOMrbAxUwWS/nBFuet1h+j6iu+q3WXa4rHiCJ
cQCJxUwTJqqJZvnUZBvoQ7qWajYgieuPEAyjeGFfncKCRBweD2ZT5ANLw1YWTRiDmGbXmgDdcn4C
/wP4O6FauiG8YIpc2mHUX7p4Eg3JPTnNj+kjBZhasMv87z76ARE31oBky0HozZRrlTMlaB+l1c/h
h6Lki5zKSI7kXDzr0Gc6L+XHynjZ7Sn8Y0QRo/6R/GNQgPaszH4EgJ02oI8b6+aeg6/p1fPkimnI
W9jSH/0fPuYV+yDyJa8zJirLTgAxBp+hAADHB5Yyv9+aj9s4ALxItELGK8SjMHlwCjfiRdmn2wNG
DOkole9qIPi5fbdL1pNpC9OmxbC7b0qGo0hSAzZ+IpaATfetn3GplsWGWkl41+//22Fq6MzBPXND
Zx29293zWs5RExUbc1YnpuqLKuneJGhcqWtMC/aDjy/3bHgB1UC2kcZuDXGtwsKJc6Dt7SR8Yr/N
P9NImSCmQkVSf8LqPyCVmVN7o2nQNHYpLptDcwbrx59t43M0yqDnsbEe3+gBQutt3btTsMO/KhSf
B/mzp3eufCXjU49Siw+tA7qbBrU0Zx29CtRP6+RZpajcupYA5sH6pcXozD+2Sw2G7JAFFYvYOTpt
Alw31KZZ6MbUSiIJR84aeiUe9ltvst3jpHFQFi/LP7iwgsUGjqXVXVxw0kKFGPnG2SSVn7oiBPOG
ale2fA1q0X8IcwdM6qPC5QG9namXKFZZdU0AaIc6M3cywIBa3tKDXyf2fOH0quik7mAWQyDo7LKp
obVE43l7L3Ceo0c4PBiMYGLpEP6xL2hMABoFXSW17HN6FTjNuKtj8HqIOj3eBsjQpPpUOt8g/3cz
/ThCdKijAm+Lmkc4iw6wo5q0x0xnerISQSn67DqeCPpiMhiZtlJB4LrSfh6RORToDGWNuvnSgv/W
Q1yrzy1PvfojG0XybtmM5momdpggbmNCRSDIyKA1i0/iTUwHZliYUGdkaBTD41DG62AUR3jrRkK4
Zlh46wQZlD9KtzZowUdDbBGYYbT/A+4DGGQQeQQiwmc2CIMBPiYzNwu8Dw+51pwPpv7gI491dBYK
eQOlKAYfGQSZrQ4MQslLj6l0xBjoppPh2Tl05JkTHvW9shTRqDDlTEv/mUAHxlPmIBQwC3fJ3azG
oWXLeXbTzko1IpmuLdce/+ahIYQimwQpx03jM4WGpTsLK6jumvjuwH9O8Si7aVz70axj82W7gg2Q
74I3zghaF92IhA1GTnnDHGHhTjWHm2YPeGEBJ4EQEim+HksWLUzw21D3ew9c1iP+880Mx/b+R044
5xcqGjjylroPDNjn0OgHR+KGOMe949kCKzFlJmUHi2V8VKIrxLGF/jw64d6CuExM0zqZ3aD/Welz
MWIeumKnARk2nrDk8aQgp5SmQNpgSBAVc16SMEvksGokbEoW1zRee5rvzcbCk4rvQz27zzsNMbsW
rBh97Ldxe4RYCG4pAhSrtl7wwWuw6eo6qXlM2T6JBLeWLOImRbgfxjEBVk3XpwNgoeuvVgAEfDgn
f1l3yexf8gszOBxmOsy0yy5zXYTC8ldmdON9pF3sglzHNw5jG89mm4j6x6+ZgNfVIgc9ziOlWF/a
Ubc6XfFq/f0W9klt1b2RDLc3NLyMd3cCJ7EhrdUgg3/UBReNVPqqaQ4cSOJosswZykBtjfz9wjLf
+JI0eT5tKXshYCh+uVLdufuvInZeJzsC5OccISpJQB9mT3SyB6P3QtBzY+TGYpWl6ArHmUF5/9vp
X35jT1kxTexmPtByUCnn7QI94PCd+m3XzmM7A0CVPW7Axd86QavwDv1AB9waZcycLhVe4lbM8cf7
ZNywyfLcCuoF96dSymYuSoz4qywVSLsDeeey3cAVds166iAtJzPd28zqwhFjsfinzHl+iKocrxGc
3yq2nHJVCOg/SYuiBCvl+67ziBo7gHXSVBHXvGbm+0lMcUgLSkwagezDBVskcQydpc9G8PrfGQ0/
Qa3o5XCfpZBTjA0qeo+BEoScWK88eqwa/lCM/wzaqd0tGrae85/XSNHUFqHWK/QfoWOBpfgeIbmp
6r5F6u7dqfPncwTyOMJjz1SyEfrMTwnGpWaqb0XVN3oqF/g1WmbT8d3eEWmzEYbhxt9hCTBJhPpY
6HgV7RGE8ehDWwcMKhXx15x33zkHFLoyCA7xyt16PuExIR+MxSQuwZaETRD8LT7q3/CRpzn2J8jI
gq7zit1TwBygB7xSEH4oJlsYaXh8Ee5JvuSfa8GsgdEymGuaZbT/CP0pIiu/I9qCKW25fWBUnCGv
19Ig8XXy9c9CnsI1mHXt2cPsnr4MDxvYyPAGZp79S+TlvTb89YYj3WtukUTyhsS9o2kfRsxm3PjM
D8EE1YZtZJzQUb3uywuFC0+3bjTVEihFz9X7LKC82vvB9a1L99a5McXd06tQ2K+nvjxk9p9Qyw6T
cvOKppNHYoaogI28zUnVGGix5cunSx6g83eLPzqe2ZWxhtT2s5B5nHe681qbqG4m9Oe6uXf0meGI
eEut2fm69dYHi0Wd1V8QM9byiL9ntQzyw0nRVgxaxRVRBONHSJTw30apcXRyRGrs3zQPAVQL7+UD
aJ43Iw2wsnNfDh+L/EzMHpT4XuhAyxVwuBORCEZvrMNSIBRK8sbiWQX4cy+kPrby27mxQ4lRSsH6
8rIcO7c6cKxKWxZW6qU98PCSbDw6Bs11y7KJNloKRMiDcnh+/+/RSjod9gGocPAkorZSg0i6OZOl
Ap+jA1e+wYAHANqW9dcFceYzOjC2ipgTjdWrmK0Dd9VmMxoReBUsvmcz+cSm+bnIxsDulaKUTVjQ
OSzc74jcMWfnEjlEu0Iv7tRl3W7jOROoa2bKl1ecUaHxBAUaLFOP8iKIWYiplIfsHqlUP9MqcRFA
pHSIlU4IRYurelKNwGpQZzQQ9ZxOaR/Ldlw/w+92Pk3ccJEpd0BKhbB1lWNbEZonR5YONZ9399ma
3iiHzcksTReFwEFqX6bo5DEki9E5yjN6Y8xQrKRMWPDYQNNrVJ5DkwFzlh9cjQdsLe46WLzYsIN/
0szRBO+k+yIFtfSphzCTZOlxix418a5eFJdGZKGqiLQMKJunRdvejanuYb4XQD7QjfdJHTfNtZln
DsNxuRUegXeRa3JR5tv9RVvTBlZITPOU4Ma2AeDaW42waLXDoI3rLdvgc6s34qlyiu3kHkt+3REO
fAGEt1Wfn1kdCrjHFkGq3dwPYo9mYXjB55ZmH94w1tXT6JeTvt0H4c6srrrt3JOxuEP0LenVv0yy
Xa9mxpXKOneguf7pEA/oCZ2oNBo1XSQaX5m9CjNFKeYxcOPc7eZDi6Ww68a0U/5PtDTAAmHVtv/Q
d9jmzxXLl7Y9RSKuOlmtrc0o/kD0RcDKaJ7UV/x172FvLO+B6COB2MO56bAF0CY0DQV2XQJCPh11
mUaVwgZ9NUVLYwzE0mAXSzuuUh11qLenZv3zryRQVc8aRD2Kspk5TDBZZYdn/vhV9JYw8V6gwAsH
I11auVTi5NhnposQBaBRpLOOi9ozakOAcyizQKAI02R4oBxR8WICvJ0K4INn2iz8biwUlTLv0uSj
26ykdFb7k8JFGMJyvzIuyUGKKjjL/nSfoCmCurhLCf4FheYkfXL6McgV52gI4WaZl+XTzQUiY/RU
a7ELrKz+HZo2PnsXdDrybZAoo/g4ZRUG4OSad/4yUp4ef7/5UZSXMtV2p2EYGM5lkS7hookS7uCH
D32TZyOJgszZURL5RgZCdafYS+GQZmuUzOqGZ4L87ZyGw8Jsd/71/Tqbz+9Ju2W4JFay3ZZA+o7J
yMCyrTOHv+HbP6VyNbyE1Slm11vxN4E6Xh43+1LawfHgYHmZxMBHix0UCIIBztlouSamRzysofGL
O91ManYhl6bSZY3/PFLf0vYWCvQdJ+xfkIOy5J2OTCPBYEMFKtECjem2xljwg6DM9GlDpzDyvIM1
NKhALINDyvIHU5CGeDxtbN8jiQ+J6wwpkN5ilNUHqBz3AmECyKvnJDgY/umJRv9CuNb9hBOXRfu9
sGt4YDqZ8OPSio64KjnMApsztb2QZe8cOSMofbqIXgvKz4QiQGS0/r1KOzXpvLfOy2bqQKABwOja
v60Nwzse4w1h4o1GXAsx/WShNbENKWPoss1oybM/Z/WqdKgBCYJWIBzMnGubnC2cig1y2BOmC8d3
vRl0GMbHgWLQcFGtVMUlNBriqg3KixOBUloOhmxxnDwTubw8A4QCTpJOTpCPw7rSMmPDDwczVSlO
5xFdTo/bn6dvcBmcR7r49kqIeRarKaE5KXSQPQQVHzyJdyXF4DEkuHJ7A9ja/LVZSLOG47Pla7Wp
e/asomr8xizS9/VBHHlshzbVghXhOINDK3xMCVH+zGFDitcDunWlKZvjHZyl3p6XNG1yysLz4wCy
o9WLL6zy/Flen4NnXfH2EdGUDgJDOUf79eUlGtKGmoE+qTZWfZgfi+vqrPnLNmshIJJcYAD5HYJt
3H9/NyWdUAnUG9B9gKOSE+NC+z/iSMKpuYVWI32K4JH83w3fqXewHFi/fXbzWbOO/cqIKNrMf8D6
upoR5aWYUEw7eoyIecdSc2cIZVXPUd0GqVuctOIb82XaTFuAr8fvNnruF3zLd3IXTkYsyQcqa6Dn
UpruOMyBbHG10SlfHPqFXs2M4wy3WeFc5iPwRrA/okjw7wwiX5SizYRuenPY68ByWsbStx5zkpjq
T3jzHdavZXm8htqWhVGcLA/zA8A8ijo+pErpu9gzJ9pqmzDLaAVrdPY5oKXi9wFOo5wzQEDOIXjh
iJzO8YEm7xo5RZ+9m4OJ1OX+eOYSg6TZ1Bd6x5si3UejJkLudXufSPk9krOFNqo8+n1FbvHzCW6w
GGgeDaHVlYc+3n40woIbCt1VYkTDIGqwOtE1SveGYl9wFds+D9nt5vwQxYSSM+mUWCdWmaqIniDJ
Pxz+tbd5Uztgztl319lmycvuU5NrekCd3NE+00ttpIZ0RJ8Azoc86GjnTi33gTscyCnCzCbF5YlL
zHyyadxCm8nUImXOfFXdt4oI8EPaqFn4HY0jIJXUIwetFP3/hMH+tt+Kd9GW+nXbydrkcjgrJnk6
Qb28yR4MyUpaHOR7s8cpd0mNEP9hgU6S/m7jgrC82nOFp/WQ6pVRHf+kF3JccnucA/znHR+tWmvQ
E9T3hOFfEa5fj5FrEaacRe3EhyAZnaUAB1fMMoQ/jVuixQjZA/xkBV9PvD5ojL6I2RsfkWi/tzaa
yLmmgAyiVT56JwqBHwutJeptbRx0fWP90kxMGgvwOc/9erq6vGV96pqr4YMM4em4eDkgGn5aPPKf
b5btS8ZasGQvQykYpI0j42oQJFbdMYa183UUwyyhr2w78NRKu0tUNfLJh91/f3PF3ut92I6v+mjJ
XNwp19EeD84AZRgYZnSNVba25RoIM1t//ZG2fUac/u7atandjgH0AaS1G1cdDGseJqOjxK9mB2tc
5tb6vN4/VZ1J6ZiGlIMzJNkMk7DMMMdr4q4uVlqWJQbVz1kxkHY9kazg0odAKGRc3FzQ/YFdBNA2
nfCoKY9Q0O/zKMiSEkBiJvk6QsFXDq3LJyXgrXl+cMqmqkxhK8Cx66Y/1NJ9nPpQUEaNtE6JrKUP
acV2N9rbdZsFCxKDPgbbUaSGse9SoVqSTvTSGzimyGTZo+S7p98Xsi5dRPIoO6Uo2YXImrXyLw1/
j2pxPOmqz6SnJbGKh4tRd1PGHnAR0eVsnDPP527J3VW1lL2B4Bl406J/deTd0li16clA7/AdvYe+
mmWe+VZCWUJj4rmvt4GEU4jIcEriJ4MJY3Mv8l6nMAub0+FGZrQZj4Npw7wMqlXuxX4vIcMmhdGq
OgKh7bN2SrVBOcTFyNhKTju4VsI652v/gdr3TuFH6aoKVBGt+etAqiRjmAjt2Go8EnmToAF6Gj2O
zZi5zAWttqnrH0oCH+aH8afRMsP6aZTyAkTaG+TXlOrLeJy5mJ0v6eFmnfIHYafxIaJNSDea7uNE
hFxxMoupVDT7X1tDMMQJgT0T/yIJP3YiRaNZ5+6xP5g2z+RslfkVH2CUtIUzE9lSRtbzHyo9gx5x
Z4ZeHM1hgc7n9lnI6s3yCYyICAQo+bU4lwvvLtYLT4r5DiPsaRzVdwWGxZKmL3GXwmWv++h/actR
ua9crAwiXEk3i4M6/dA6IMxWRHqshulFVngjt09t4Lutsfl84xRMEyFFxYkJUFCHLpEu2i5B3yLZ
dcTTtBsQvtCIIbQtsLl3h5YcH5winoesCHhgunq4Rf3HiSS2KZtpDGovW3z/eN8CmZQf4WPu9n1o
3st8GJrbfvTNGC/qyLeZGrboS7w89XRJoeSdOoug23EKe6oc7OZpJjr/t249zw42x2e6iMs0MLfE
8Xc/PpKD40l3+lq4DOsoef3t1NQ4ytIFOKBNYiLwtjVNOwnr2opF3F0Mb/Qspvh32ogdDvpeV0JE
vloqIcmPipZkHGZrBnPwd0H+Xo+tmnsBTcN8ivocpEwMsKClUZQ6wP1Jjdfs5VSBD+hCLcNzCbJT
AYT1+RkNuVUBfggLswlZaRqKMHpVLEbkGI3GAbsp/8tFQrVIxX2p8j1i3oVZenkLK4hjAyFWE4yQ
TsQF4qGNHbJpjDAywNgLhtwjrz0IPhYWjrEIUFCrTRFUUwc3g0HIqNYuuKOFlH3zz36s51xiZBZW
NJ5xAB1YA8ObI+JzCcLbrfrE0tM2nkNZHh3hRhpEPOCeoPuL9XvBRUwf/5hMYKSvRFL6G4+ZFbip
QK9xK2/1poYsOTpoMoj7HmVJIj6uD3+oToqudSUxE2LFmIep1LmWKtldlAmn7keMWtK97ON2y4MM
0MynazQmideMLtSxd0GYrEjJuFKC95dMdDYsA0bumlCrEMruvfW9/iZBTf35VtBGAl8RuJnFuf2s
5uvKIadRMmU9Uyltx7AkHDNbLTVvh1sL4NtwDb5wlhpNAVXDO96a9/27ShNuGwVdbL+o6whyFIgf
609gyiTTf33VcBBWK8+8PDrPzr80BmIUYtfvTe+qAhML7bVyEHmBNN41UzHxGcRGYOtPYgjWo2w5
b8ATyHwTpl0zIfJ6QbeYXR9nSYZHYvtwhoUw3LCIWMxPFXkKsMkMa4l6cc/Etgi3+2jSHXTbHdMc
omOHrTvIaM/x6ruxBoU9c3x0viJXCKSCbpII+lFXG8nuiMCMx9TilgzwGjd7FwSyeAwsL8eF5Jnz
D+SyyDZbDNA1g8Jh/lvjUyDFSz4WvvNKxvD34CZJa3NRaBNXsPzUHtDih6AuHLa7C006Zs7Qc7VT
FfuQwGkium/087jiw3MnFL0csF3v9Udcw+YvrJMZbmgmX8bvKjHPifs9dLLZGBlUxQGklLfN8Tzj
TXxam8wQHQJR/R5+Q2zTb8//dWWWD2D9FOLa5p7+8FVjCam/7knPX0PyH5tx53GWKyaG9EgcFagg
lmECcSPtaGdzcjTrdWIwLuGtawFILnSHGP26ZrcTMOo6QZUlyGgXkMk4c+rRlEC9FQajGBF5ksgO
R/xxJcv3dNlgNZShg+08Z6TR4Wppd+VWYRxKwqZqdzoiIn+zT7mst3zMl+NBnDShGfku1Dz5RFh8
ZYl0wHOfU/mb7u+haLdDY/l4GzBkvGJT+2x5OQbknq2bM7orL0yYvOxTMGVGwRWqUwifbZHmkX5O
HxfeMssm3p7fdhGZUQFCGxsIVDzQ19F/549EZjcUh8DMU9vuw0ezqaoBk52OVwY+FKH2NA+fCD4t
Yclu0EdGinqw8XYHao9kRGd1Biab7fE4FTik6y9XK72NCF3YEVqPYn3qEdDTa0i/oLdIR829nRb9
ucEmkK/dIm8/v33KfxOVE/JRtFbNz/ql/t+uzXmjdYpIkq65GShUe7OI0a8m29mj/pKAKovbDjhO
XaJ7LwDxyLYgT22tJYQwFa8RGyDsEcCZy7Z0zJNj++b2AHj+RUUKz4jKqLEiAaFosBOdch+eMZZB
igz6iAnS3Exsw+qDOAJ9mVeKuNleiW7JjDoniHbEE8g8RyHCUUP76YYgm2ac5qXZywID4tiEnpz5
b8HobORxzdYTm5GBX6xi5Nmk831nG0tFc2ltVcvrDuSb1XJCCviLCQmUj+1uGpuhUC2ajvM09Slj
aUEZh02h7vnddz4JS7mAU4z8+rmmhyzAsIu4LlIHF531ur73ON26M9I0bTsK/+WtK/prN8jjtLnZ
jG0hMc+FtNmSNxVybl3KXq4DzrJjLweplcDHihSjxIvGbViBz5VpRrQGBVLbiiCzCmVRQnMdN/ae
jWRga1CGJKMW+QIrSZwpzSej4g70BG/n0bSy95/FZWLSlC6E3zkMVYfQqQdJoTUxe1eyF6o0Ihv4
glyysG6nem4ZKB1CptZcUt0QAKBDVWnwA/uo+BZ3EtVlTzAzPa/NrRdFOitYMsdPxMDtfLjApFiF
Vxq3oeUXsk/hL4AS8j2iVXRp6liFA37VK78x3cZ/sNF+4jvnX2NlnJBKuSr6Xdi39umy7CdMyFg5
mOv0t9es04iZedfqqFsCn8AFT97qJqWvpecTTA5aYokYYmNe3/3WkvlNIX8SizY1l7XgucRGUDvY
MoOWPq2XPfJ9VmSysMPKFSOg45Yj4WvWnyL1gTdYXebG/Z9bJScYPukHAlD7GQJQiej804QJNkNS
iyqTvNUUmpFSu/yeOjq2ZN2+HlLCtTiaJxY8G/3XiXVWMlokXUyvu8Ui3LkifPdO5iMMjGglq9oy
b4wvfeTD9z1/GaVhX5YiWvGyJB3a30nLyVHiD8v6xWRnfiI4LW7EW7614vYEYRseNPWdvni8vfnh
fdBVE/hEm8QmROYLFxB9MCT16r84OEtLCDruGRsC91IW2AGw88FwDizgALp7bj3a6s5JbGyQAMEU
Diwwx/UHJ7BnQ3U4Op9+186Dd9gBQKG6xWj3hgMnJGSPP7qNJlCQydMbbkSJvo8HTJLLrIhdHoT/
Gtlkz5XsFnqrgVTaUWErSj3obvH1+ik8UQRlrsXFMHHKHgqm6bZV0VgQYorf03cGAF4DlWa6R3Oc
dhaYXtQH5B4766XrU4o+PXU5Xy11aIn+KgmMLcG6kiiykAqGqR99jBuCS+8RQVyl/T/I3D5yr4ek
eQnQzRUrm2B2I79XgYAB6Y9vELBgxXklUr7KM9yDI/TqyNygT5zLwFeHrKpQ/s8IMZeZdfM7LeFi
GBm7nCTkkwgqrm7D6COaC701O2VT1coIg1SESjc7YlHMUjDtZ1ZD54A0M/x/ueDpfD7rKlU8vr+B
YJCiE8dYev1qmj6VEDPgF9pcMdTKa85Zsm4msLii/vl/bugTsHjR31mHyVxM+g3QPZn1kqk/kvy/
cFHUvXsjX5tdjITFsjdROt5qE5Qc7oUCi/v/XhxpqO549p3WzW4igiJCN8bF2600feBq9Qsw/qyI
lI6jXifjBVFRyFFlXfB+q/jc4SwIq9TnkcgL6zOuj7W1yjyM/i2Xg6uJhRbLCXdo86WT2Y1jFDGi
izrg3FJ3NZLLlR+x2b2mv4jPm0w125DLE8oVu2bNM0OgUgps3pP0NLoQAncgH+8A54o+lFnfOlzL
r9r3o4Zh4xdrFgQaqnxuxpIIHBp5fph0sx0hT1+8ujdCMrjiXv0+mte3Y2ZxuGqSy78NgXCMDWYK
R9bv5eAkF9XIJa0uEDoHxaCjfnHYt6zfXqCBMmPRvAkbYFK/t2mzWmLHsCTLEgFROmJoA4C44Ka/
ZEny+wjyQKHFtMDy8k6O2enWIFFRLYhhAAkrysTgXTPl1yeewhugJLQl9VJwJAgsp8RqDgIIm7xZ
M73k2loSk3WnB7UL9VYn70SmGhC6DuKPliQPAeUJMoRmtw7zdvA/SMKAcO0+iBMMcEMLqIaKxW1A
4mD3bl3j4l4B9i0GRy8ndFSqVngvQzeghnmqx/TEpnMaF/lhpEIWHurouCyNJbulXv56l+IbdCTI
tUvnTR//06BF7EBJtTuG65WhuaM1nXF5VUy7JKV10YibYLhMkpeoTd6pFDsdLke7Enn/+bOeB/fS
jKRFHP6nud3Di92MusoEg1Z23Osx8jGtB2y8Ht4L9mxw8XJqIrTHWzWUmoWgkwjHLNmCRAEF7QRk
rDeNy3FQh5Ef6g7AMUkSC2cKt2HdR+dp/dwOo9XIuoG3YMXomR5DRyETev7uRDiX09mvjVLRWm3d
7FsaRc/YWmI0ONMVW5KXLVm+ZAsrt7CvtEN3CpyCfrkpy5VIhFGj4hCCq6ceIt/wLVuJ9/mpziwp
kv8ZigL3UTRk8hmPH3B3ddwr02mesG3v/DkIGVsGI4GOOuJExhetOgP2DsjUz0+/Q82n4ZRb/kzr
ikZsPPY6mT5iTX4eG7GFjstqvqiZcpuLeda41zrs4MV9LgGrZ7Nvl959FTQ4UIRxj2uhESfkWesQ
TZd2lTkkiodkLCI9Cky3ifrxpZVbgnrNPGkaqVftUD3b3N5r4D0UCzbFaF07Tc6+bwD6MOyqTkNl
CneFWPFiZ/M8iQOBTyBs9NO19JRZxHn1tnCLJE9Lyu7zDbrJQxHp2VEHGHHxKNw1YgQ37wWG2D5d
c7165PNlqz6BGRRk2m4t1VmXG7eDbf2VsqVEexCiy5Ygwn0vMRGXlle3UCZJl3R6+ktbf+ioDYtf
68YSM2ChgPh6dZiQvKN9zAsz7nXsygl6SoFQ3GXxVdN63+60/rkINtgx1RUHaiv370orn65FErak
KcmgzFwRMnkPWwegyoztqgBycdnO+/jdEGO/q4roPPEHd3rI6lbomSNgoKhi79x0SbFOwqjrAPhS
+qcGawbk5wjRTrKZjn8Di26c0oz+DYlBn7wz0MsPsFCQWtd6FWYP0P4pZlOuvH5ox50Xl5RUFaUD
17yfJjp/vQLCiJlKl0UJdQWpEEPbPPLak6BXXR/gsm4XVCqgEOsC/8YGy2VKmoXVALyxY0DCdZ9p
UjeR0ltCuCeoAg1gf1qAwRbemvZpSiK2C19VsYhM6xn/Qq7D9A8nmQYNLccz8Z9H8BALwJtVon4I
qLAVKh5pzYFdhYgIaHxNPpSSjaiKHyOttl4gegVRhfo7iDKoEckKxGQw+7BWkXVN0MXtQseNOost
VwjXE4F/g7w7vWop+spCflqLro5X1rqnaYTwUL8RE5KpQzs39CYf1FZ9Oy/YtBWm4y0ldPNfMNPw
r6f4HtOtGM7jPWB8qi/CfLOsLC0LptitkFA7FoRdeE+Gx3ICvL2eezGUyc3fmo/uM7MJTyb3Qk/I
Fb6fcJsSMZVgNctFGTQ/qGkfrAF7J1P8mYExzcZt4ba5fLGai30hb8yWxnI9j+d2O8kiyAq6rFk+
2YpmxvJefDKQ4r/p9UtZ6SJ3ATp9KBNRhtLFoOV8M57lPy3ceYomQHKR+BmR1lm6s8cewpVrqwSk
I7fWhQCO7foORfF+j2GfMex5WQM302D4yjH7u6bD+ADw5QAMu8SXAfElLkz5YpmSZ0YErid6GsQ2
1E3d/3kP6Pzljp/8wsAyaJvsuqssR7p2cCVvt/aFk1XZD/+GfZUcILeEhmHIE3NBGHfLIA3oLyZV
WeveSvCk6oey/gBEGvlz4cH3tKE5IIngeu1v7Jl55lWdnpuYgdQlN9F1LrUl5vjPK5RppYdWifSf
ZRzeckmv8WwgLRzazgPMov1rACALrml2S5dpgM27KAaT6hvJaZZYwIvAshMvxbc41oaa4yxOMctS
VA6Ti9rjaci9MajrfPqtaVj/3eFcgj9ynFqgn0peRpSBm+VG6tArE31Fdsnx3ddLafLDhlz5/qD5
q09QA1p64xepUboOTzqNJfv7RWB07nYHCME638BA00Q2veHKlMuFUcTFSmaQAvWwLva5lIXe29km
o5vyzUjY0BGVd9QreVOZr8UN0UpYiLK4wxKYukjq4TtdpnxQapZ7x3FpLgDMCNWhahrK+ECAuMm7
7QwwdPRaYS9+xEBWjY15BW7AAkb+nbKCvASl+6UYwZpnwWprACCXUmnavG29GySDbxfwqBK5wRo5
EO30dOWnFJKB0MCwBEIAonFJ5NxAT99tY3FICqcC2FUl/SA8tMaOmTQqjeyitrxyPWaphNdUfB1B
/XDn68X5MtJ5++1Bj6MkPaw/dmBfcczO8ecGf+bfHVNDsx26yUAMZapoeycR5Vl5dBbrczJi1zFo
/XlVrCN4KErBDiEcd/lWDMSzT80xfuTbf4RKucAx2afxFNz29FS0E/O93ywfj10uxbSAhpEWKROd
3A0EL/LJuzlI1eABpYsJ8pc5E5XgCA66KeYLpil8M8QDuEwq5VKUuaWybF/7yslxhc/+0qWE3ehI
/ZvQnIPC6L1QdEkmzZ3Fs99kfa0PN9WoAMTYlNDuucRFyDDUtqkrSJndLNWHdUuhE7cxm/L2rG8G
K7aqt7zlsIooGDXI+eDS8/rQJ61YlFfit+jJHZR0Lt64fcG4fEutLfkGXbqg+C/6oSvYaOiBF6GG
tk+rGIAv71P74qm1LmocLJVsSjq53XFpGp+h075riCPYH608jWQ/I8OZkWbJxo5I5wzZPLk5ijSY
NRQXL5EoX7W0oRoP2GmVF1ujpEOcPXiCg5mvG1aqsY3Qj8seCbosRIiAKPgDB5cL/N5E5w2MD/+F
QscOWGjOQwvjwlKsQqFdP0aylyVOqqdVPU5e0peyGIyEl1jXyJSJJrwws4pj3pZy7vpEYdo72fzF
newUMAWWKCNNWabuSoVkH0FUeIJP2qeOOqQmVz0dVjjDhVR7Jjo2Y5F8pAIus/a3M0DmuOu8zdYM
gRfeyvUWjOMMT4gEdmkoLvr3gT1aUSVPYIcIM6mo1hg4M56hYjC/2kkXJ7LylaU19LWoLVX5jUHy
fSB+grPW/FvVqSJAk5JtIVjDhLUhTqusm5PsWhswXNMxajUpbxJaP3kuP+IyjaSPTOkWvF5/CNAk
CTUQkFOVT36zU9OEVAxWeGol6FFqPftdn+PSigmCV54SZV62HBDbX66Fn3MTBejQyrFsEjOntaEA
M5Kpc8/QXESlGJnP5BFAhNvxgi0PPk6KdjueBY6XB/Bi+eArPtXEkJHlDX7csKdjmS6GsYZM3Xvt
uznpzQAqcTqc69g/SzdLkGekZs2wQ/tYYnt/FiZHQJyuNclTkW77BHC55YOcx1T0gsA907IoUXue
9qfWC9j/R+JPTRnrXC4CxEcKiHE7xCIcx95PejPaByvbfXAx4axIWEPw1V7tWrAf52Bwl5t5wxUK
+zp4brKAJxKrLWXM3NDQxZYrN4IfLwggvLlkNlYtFMlFALYhfUv/6OHqdqy0DxfdcLhDv1CpF/vb
br+kW23Wsw5RC15NIfucSFg/iBR3eRAPh71eiD6rrhB5cVoD9B1xhDNirjXEA4RAOTxxLwziVrkw
E5FnzB2mZopVk+a8FfznI1Z/J2w37jE2RogNnU3LdUeOroaB6Vkyv1c1XJHsWu97pbAyM9xYPP2s
YjpfcFUjv/8MLWdo374Q/05zA4iPqA6ZO47eP7OomZEbdDyapULumTUrDlGfOdfoJ0h8Edso+nP9
zUXESDr3Ke9vnCNLu18KvRGI5GdLilUqpprVSZpCYSLWyUrXMeCoKxIsq7bE2p2GYVDyOBHEesC8
ZvqIDXnPc65llNSAtj7HvtATZVrG+JLqB+WeUfv9MVihoj+fpEoS1drmCNrm7sCYXDD0ejn0xqni
3Hm1h8Q9w0k/PFCGinqqIrWqC1OYfy1GtOkyDSSRI4mczzBWKXNS6Y7nBVZQkkeUBIADrxXrJghw
LABSnjlgwpw3oSn2i5R87bvCWmVo7zRqP4kKhZf07ZBhzuZxAQNWPKAunQLLpoYWFjngNNyWf5hL
xh9U+JHrjdrDQJYybaGUvBp0wBAJracF7nEkQcgBZeN5rHWeqbdx6kqJJeF+Su/yKLRqDkEGSRio
n2gJel4HwJcoYmZ+FFnM209SPfZhLFQUuHIZZewYd5Wmp0cpZqAC5BtXXiq4pSY/AqlRE3rF24+k
VbeM30uO0fqWOKUEE2s4KS2pOQ/4J0dqO8LD3m8z8RqUwS/EwNUHrgLytElyksq/XAiRtlpDqj3v
M8XB0ldaRDhBk759thIoRyCDwoIWvzydEvdyl2DB8VAU0idqzYIz36/UDssU0qoHBdC2Ice613H/
TAN6tGed5dnI2ss2q3RSFt9YZNd3AR30KMzVTBPfJYol9qJvSsQaK6FN1e+kWTaUoMV1preE1TpE
SRCBcJbEt09q2wRfIXcZmiAu7cOkcdie3ABq1DNfKWB2l38K7mVGqPBzRptd/uxrzzFJytiDcM1L
e7SMuhjoayl0NKv89Y08kJQZ+rDPiblCRxNScBjPc1cJC6xELP+NcDCufDibfHPOWYMLBKmm+18g
3zKGH0qN4TCD3hB8RKsrOMeNe4oANmTBZERZ0+UCIwCYtNv9w/b927ZkmVbij0oHCNgxpM4jJo8q
aXtIXH0f6N1MuekjKn5dUV/9vYw+Z27dT+eibW2YZZxS0v5d+62HJabizBi8ZlDY5Op5UoOiR+1m
Ckf71swqam6Jf5EKuXbxvutGfKFTQwMZn3mUr6U9p85KdnGvKvog6w+VQv0PaItzWcNW8bIQ6qDY
mUX5ChcKEv3kehoSjSOLKtN8qPpKzdY2FxlwpMhe75dGJ603YiL8AtAYnP7IV/zU8jGeLsZZAT0G
FoolnJs6qCVYokkRtieHz7h6f2xA4kVEbs/VTZj3xoACAvgwBbo48JkwqTkZ/YF5VXTJRiKPAyEU
EqAk2tqUebc4TeqfHDDu/A8dMOtjAkt7B2SpHX6IBlWehsRBEwU4BP5+57nqjT3j9KZKtT5tIpsK
zxNOWw1fk4lXIxswWq+Kfr6l+/e0/vGNlcM5rjJKiOdrr/5N+z+ScH6psLm6FM+b3QG5DYvMwxd+
xu7rBZCxmF1XL7iCiuu13uFFyuZrUq7AjZqbAX5MDbv/35JoIdwgNK0KeX2Kx3WkAyExHwSr//t3
ToIhJz0Q9tjQ1DvTADy8A0yUR4BKAPjug0kAHzHNY4sgZpTOhf/l7wYlhidzZiiwWRJ/r0RUX1MK
0qsG9s4pntz8T4XVq2hZLhsHDthJGHjTdOa+dTh5aK4NhAJAUD97RaQ3UB6r94ey22yuwP0Pn9L+
3NX+a2iA63baD9KRerh62IUzbSJvwrA31WGJ0GB/xFpB1Y1R7V1jUdHgBiKutqGX6kygNerwOAKW
3SFZbT3u/FMjfLzk+RtH+bQ51nsVniQtMekBo7J5s8yx7d+ny/AhoJ9AXlvcVR++NAoAHYfMx9XN
SGToNONsTEbfpqwtfnYHMqwc7xi+g/MzJfibc1fRoxT3eyea+Mh52JbqEXyDjT/pIrB6wxEYi3SO
MxKlpR2OLSyaGCLBU8pQS/AXSJBrpovVg0r3pFlG1xR5lqhzhkmRUUKUAfvN4lVepnrG7c0Cen81
fCGhCEtjztvyiW9Jfa01L0aaQmmmBbW3qlE91apUPLLtttppXIh5gcCLTyWkdEsbnxZat1UTs7c7
5z2TG5YQFslpeNO+GmjX0gDzr6roPQhw1QYfo6Mcno2z8vcIp95MrtIVa8+bfCXBOejcmG+fi7/k
thxRtY9gLKJs5QHJ3I/XLRpnINPCSdjehiBl9ovLO3+Mr8VM5DcF/ZLuL6gmz888ODWefzJ52CBP
ksbaMU2QfvZkUoN8sFfEySuiLfhBH+tW8kRj029P5la83CGBpJkpCg0cvi6qJ+g8kvzbJSwhVIE5
U7DsjU3MD9VI+CRk2uKIw0AY0bc+FsHJaAHxt9oVpP5SqocrWkzg9FKGeQpWd4rAQ1R3VLNhLsie
SkiqVCIJ5YAYyl73Y7zerxhfQMf/RfwPAGYh8+Ledim0/Yg9Xf9vi1/nVBLFuQdLlgR1JccTp8vP
RcPp8TSq0xvVoPxqRJ1F+tMZeanMmQ+xT2evpwDm0agDxCJBDa6lD0EKbjs8o9pNk8DOP+qR4D69
4YPDUo7BT2NR8XdUa5JbTXl0USLQmL41jpWUfCIQDPKUQVsYgBDUxCulOCMryNL03AraMK6M14wU
ehriiFBCnEaL79WBReu8iZGsStM9ywgKs2aAI5wUh8BH2x2PVL8S2xqGi+WWpbCJ4Vtf3EuyCW6H
XBbRs92chIpjo5EsqjN0OS7ra8jq4/9t8dc8Hl9s4TvSloYyXHZrm0Va7yY7M9n12xr5kozZsm/S
4EuTtB+W3MR0Ur0/oL36O5ZB+RZSKhMfIKjEcr7T29+cN9obd5Y7OVT96VNZldHEi3gtBsMSmwIt
OmEKSBqM4nlQNkujJRqnJVJTmiWyTDkyhafhm3SddPdCMIQ7ogGN5z01DAc9eBqfyExeu5m+OY/9
h+ygT5yfvTWS3xUQBnD0hoTcrd0EgJDO56FEXtxa0MgtLDXfSWGuk/331XkaxEFvz/9geYrTgLvR
R5DEbCAWkkGVKcro/2/TK1FuloMbEDoPm1vPzvQUCKvOPkKP7mMecvYe8jG+SFGqIw6Lei9yoGJ4
oHnafurErB+mMChTuGzMbpmsVxFBhq0U+kPBCJNIjuNAgHRZzmGwP3mzL97rRfR6ZTEEkJ15LNlN
cAyWAblqKWve76K1EMuTLI58nJgUVh8ngL4E5VV4q/SlhLDU2EGP0Cq3W4A0//cp9io570cbR9mn
algS73jLp5QQyUQaNp4Pa8LnU6V3V+enBRal+zKHJuhYJOS92mZHvUSXCo465UIDWHet7yCAKc+h
fuXEITLUv/GD7JiZw5e6g+I9exrqajcHAbg6Q0Irqif5IebbNbnMJGKTctSDXi92sc06lU569SsF
dq3CpJYTG0Pw4NxicFzCF7nyN4W8mitQGBygoX6sZbUSGqZ6Njiq/L9w8WCwc3VnhVTSbNngjlV4
YvB2FqF2nCDlRzPY6TotYY5iGUFfe8z1cEi56uafZEDFVQmduiP1/EKi5yRdXkGGf6YPpq0J8ruz
KYC48dJlJ23YT97JyoTQ+UglNxBwmQZEodqD+i/Fpb/AeRx7QqhtWNelaLFaEMST7QpnwI/pBbYz
mY2+eRWueSd4i7Dm8aMe5qST+FkRFXRAC0d9d5n+hO7zpqe9I+LgDlC2aOraQ4ZT94qJTqCrBZru
tsFR53thN6bRPhmFaZiaRbvm+I8s5V9BNXIJ36UHnAI6nId4lN3Kxf0big0omoGMCjSmrj8njAw2
q+Z7yttVlPgwR1DbeC+Qida4aSGUIB+TnbxlCY1qT+xVHD4H2deiWnPQz7LXO8FjwUiKicNO+WW5
BR/n8rT2pXelot0lP5yNZrsvfpXnCB7kNNhMlKL9BDX/YgAON5Pupp9xdXAkNKjQLTNdQBP8EUZF
JaU3Zlj+tEcfXzsiIGCS0PH2Lb9tGaKWREHwpZH72sPd+Jkj5kgI65XKzPDmvZZzib7efMMQvI95
xfTr2dOiQRmB95FMluPuKe+NFiauW8ugZXf/wk0L7/lHfwTONQVwiZiR4roLDia48RBfhf3UUNvk
MgHpD8cdyqN4PTxBJgCWSQcdfTZmDgvyDoXf0II+HGHDvXj+CBM9cmy6rbF8OBFV9mnVSLJX3omP
CzyVOWAiLjcpiypxYHW4ylILft+5pJeJk8ikZOxlTtS/htRf4RSFoWjxa/CysWXfB6+p8T+9OxWB
wzfP3Qc5C2cTdb3EOxf5SVIBIimU5vFUKJob8EgpS+v4E2FLSXapWr/ORJ1/8tXCQfjaQQZHxuCy
jGq8NFOVDqTtm/IdTkkHgkAi90NMCs4Hi9F+QQgGr9UbMH1Jn6gJ80HWG84upvcE9s2qLoiNJYvu
BwRTN496H6hjyS27xh+CTK3VhdYIu8GpEPnscYfl23PdCXG//fzxSz7Gcq6p5Vr3LNp5vWHFiKrw
95wdhmX/UW+9JtCpfiCLWYttzkbT/MPcnVkiHi/nhERDz87iZwuzypcFugBZi5omd6dOOI87A+oU
cDkyFA23W9TLkfRiVF8GQlUT+lhpwaFdGU8NidOolX8pbI7p62PnaQlENef9sSlkzZlUZcLZRtmU
2Obs5r2uyd4qofr18EWbjMD8uBGeFz8FJEucqNm4O07fxqVCLuvGfvSCqvSa5KKJwsic2hBzfLhQ
YdFU/lPvQUXkxTHieCEBhw+mbv7qYWtawTLYOuWgqy95qxSZ2vKBCQpLKX//2eLzMWQuYBYv5MjV
I5SvTlRV7Y/4EZl9evfqTjaacis2r7vbifnhndzzxfFPwRGMhNPcjqBHJBdbAjuu+yPjbkHxenbs
67u4QevTNxyX+k9u5tgxH11CoMbdYVttHCi0RM7P/4KTHFwMsTYgMoNgGJwvsjw5cxqov7w9tqr4
B0seAg74FTxydAUrtaR5PhJXROng0/qMOcYJ9WCmrRqkr0Mt69Ze46ykb+ZfZ3Rydoh4FnR0PH+e
N4JGcfNLo/rJGRIFYgVgraFPwyYFQpx1R8/riL9Nf+Ckq2kdolwhvYNFBBpYzVjV5dB9bygXEL05
vMoaRWiNQ+sBjGj+qwcEciPoL+0P8Xq6M7BOr6ZF20EA5Vxd3F1+w6hZmdkAxzRU77ZAyJFddUs6
spnsfb0eTQwPjU1FQgUwqyyW9JNgA5IUDvgjA0ZPB5LVS9/ZkXHaIkj2dmaKDp17TPijsUHEOBDP
1XfYJj9BwYYnuOZQRl9zZR+UHRRlwgTBDsoSZDbmVRbj6O873/B5WmuUevR+v2rKhBdZtlEJmaKp
SSMSgxseD4c+wmFh/q9udi5TP7mXUxuG+1VGheBBiqnmHIqGdrxiZE6q+P2QlRNjJnWtjiy/3mnD
KkQE73F9JQHh5Mjshkb/6PC6yYHAw+JLbBpeTKK9aMv/kGr2gwtX+5t8BPO1v3zt5TSe06bOLaKm
q2PY4R3zWU8gRhZQpHQPd8e9G7gPEsun2+MzVhDl0uTBp/GJexAG8UaWxHlYxNdjyKDXIod+qOm5
T6FuMfhnL5YszYp/iMCEsPxwR8F+n3bVmCfWFTLVvOB0sWqfq/JpX0iTwQ2GuGX9g3h0tJ6v767U
+i66TnyhWZ/7nmnX+fos5SL9NO5BuFl0vlntil2S0r8gzqai6NnvvrFjQucL3BeM29v0bg2l3BL3
QTr5nuiklVxmPLdbfeDHcuKoI5JAzjrZbGvh5CIU87Pl2QgVqwVm/NCfDVN1FoIDYLC/03Fz1DJz
bWqdfBag1wBIRF2Yv3WlG8eJ/GOn/KOyrQXdNorgxvRL2RXlyuKLtnnma1aONTpKQx4eTGxKCB0h
YxiSkfu/SATRKVw8S6adnmB2/oMKgVbORaitwDdleZbJ+2RKw2XmLvc8fp74ynaUCas5Yq/4KySp
34OKtdG5Cbq1CS9TuWevd5QOwtmHdTTtiZk88cru3kfC64CCkLq+I6NzLwdNPmYy5Y2cV6J5T/X6
+K86FFL/UcYq0L8B//TcoYioHJVhT+EiBZuPuJ2FMaO/IxkQfS4ZpCvzsljgFV+MB/BiGdxjsxr/
sVebIUzhN+1Mw/zCHUnyiop+uqswgFwxBul/M2gFeXvRTN/54db0u0yoeX4HIN4VKCF+ZPVbah8f
W7jpClUL0hyVs1LKfDQ9Jyu9+j9M52b2vv7rtlBs875YViUng7Xuu+V3CzoKdTqGFyvaXvZnSP5W
7szHhVwYE3hSlbu7Uy0GZRgDj9YhqAnY2YPaknwGk8WmVsqV0x1VLhS4/jVAWuwgvZVFWOC/zoem
Sd9Fvm5FDFMDU3TA1Gak+cE0LCW9liFl9v4Ni9Mivc+CzW1z5HOOV8koCYVCDn+S/k9FvHRydX6d
dDP0er52B+cCKTYmnYzGhhxHALXIQ1tSi9NxtgpchcblX+mnGxvIditr53bW2muyOF2h6hznDm5K
dUNpTgM1+dOgP2pV3iOkxcQ9qsM24AUKsaJv/wePKz4sJLGNaez4VumntGzFyP4ALoTz6+yxJ/L8
uveUwP5m7KcLlMDjTCSMUtSSuNWdLH8ndPdPh04fDDy0QlPSuIenN6kyFemG5mNVNh+Y2jDTL7R4
lHDe5m7FFAtkHhachNqtJqJmBwJ2w0HwQeqrvbzFI+HeLuzyCJJPQDK5iP6WTxGmPYV+IJeHrEUa
IIIvTKW2dYcwSEXbFsrLD43I3ogREXbfzR+3HordjDtkYwIZgcDa3HEzicf5UdH1+4WcMAwuaqhT
X0WeyEB3PhmBPVBXGPiL4BZpQ7f/vybr4q4Tcdu5QwIMrQ72jQisrsqdatz98/PUKgXRrZwXFJ1a
9iTel1fpQIxAl/r9kyxB1qAqBeMuHM9yVRZRDtnwS7rcFTMpFUMl4WVag/01O1zv8vWAhVvS8XUT
3V7i/uPJcg6YWu75uWklZwhikHI6rRF3EvKIAi0oaVBZGz5pEgxJfAHxNRy5k2r0Sw2OoGJ8YluI
YwHJWOY78f/Za5VvoKNkkJWlJYz1RC0VeJhZR0yx8b578chFd3kn3eL4ZTMJ8ZRTkxglcjX9NBqW
1bakGXz10dtjErxZtE4h1/08D12y1V/cTvugjeCkNyjK4d1ZIeOVPYYfe5A6RgnrEecOmIvdz60i
T6GrcRsQhWlAwdBZ8s/V1KLEYemH92HXS1hkpIDRQdWW6SH2ih4LnMM0Ux+hYNPP26VD3eMTvhdY
cBxlWDixRHA3XB4cES64etty62SUu9anWdXsEbhWEKF/TUki3X2ooFjwpaOTW2c4xUqPBqF3B6jv
rj7oLRcTTdl6jp+MKA0cXXgK0ycdZH888cDMfdoDzcv9trpKIei91shIc87P87QXViEMnX6XUjgV
MaO9yzWpT4+wBvMrV0uDQFKBHikCKXxgG9e88LYLnqXAgbnnNMSmCPlNUfQogNe6/7ILBBKL5gHx
2Qmjpa+fNnRrHQQpLjVXDeEOYOlqLT3e701jpQq6OSLv0Ybzztbpp/SoIn/Epvp5PmSXsNk9L3oC
s9MNAXEWiRQzygrAXWJS1HV7ER8nkgqPeoF6UiaC0qSJooU2R8x0pJ+J4rqkbDdTovc7cWmAZKlz
cluxPrjy/CG+vASU0i+dhcO8f0XAbMktzBGoJ0DNwb0sodyn0HTfSeJuQuxtqmd7L1cjENZKQdvI
8FxZyhrwfNxR2PqZ5S3ilFCBWJxfFSvqUPFmOIeoumXqAaog8rVbaMMK/mZEBOdPVa+V1hv4C3zw
3n+yuC5WpZbRNtP6Wbw9zNHKtKhhNj6/rvwdXmNL/3eoSXaS9vZAnB00gJXbkKuanIXk5cwP7Vg6
iCx52Bw1KczUGbfzhEA2WfMC/C+I671r9VVPtepwEwAyWa7UaHsJ8NG0sCDU5K2dl4SfVpk+7l2k
T5A8LWpDQkxFF5mTVdOpatV8F3Yw5pV96KwN3fwrr2XEaTkvfN/gtOgcVHZ7tccn418/iYUVFdUX
M54w0VWjk2oeu06vtRPumS8TgI2XZtIy0amBeQtIhK7AZhZ/h2cyuUCteobW1iVHOk+vTPCODdl/
BVuNpLhpSy1mxcrBuly6WtsWrpShOzRGJ9SjQ3aWGoFynfzLw184/92hNJTuUmr2BKaSYhQbkh1X
vrwjkskhEm0HcKNk7jS8YNG0dp3b+aStfbY9+PHYMZkarOPueneqasTElghC6SxrGLRD8H3Rh9MZ
ms0bheKZXWqVkFdiQ2h0JTYgVe/iCfeywCsUuyFrTUFtJV894yKUZt1kqSpR6x+HTtKyr5a38jpF
Kbby4EoOINvFO9z/4RyNIPg2GdDY4+E1NmPWARiwf2MGWZEyDpNRYAdmP7c88XbESPYkJJLS1BKp
DlKvsq3khFoZcP0rO+7tRl+y2x2gL/siJNVEDQIY6WLJEbTvjY63FsZCRB6P3j9JxH+Z04gcL9N3
JZCUKOYYRSlKUOek685Jz89Ky4canVKtSNkdpSC7iTmBAcpxiUc18tdWOS2EtdQaMi4Oe/7zFajX
EDv50uIKY4CNbKJ1RooU8AvqRZoGtBNs93ewWM4syP7VXGlh4t6D3XqkRgbkG7GyGYr3isqhURk2
eOqgXycMoGwuK4pCyKgo+c431HYIH5N+t1LamkWZCTqjeN/U1dFsCjycCiqHy0Rvj4C0FJtgRP94
wKChziTEFkaHImPkwAZdQ20lOETCdAHQ5qowyQQtOvC5gKN07KzHf6JcpnxWZnGUpYM9wju1d7Eo
PhOhAw0+F+vWnSd85y+wFWvQKUfwKg/xcf77EEObS+0Hy5rChL7YyX2hp1Jay1JYJPQI9L3OkAXW
TBn5bL1eZFnewu+gZZetEIaknOLwp0GbiDxVro0kuXT80zB0pysRXi2eJ16iQF4Y9OVzeKhDltWi
S1rY2IMbrIpgwHQ+IaH6XfxvDQMF0WZRsMCTwAn3odMOCktEHbYZLnzcVxne0dfJQwP2Du+6VgCK
CUcw/sTL3XyRWq4FR31r/baK/11k2feRRpNjCb+zYnoshDNyDB6pLlCBlcFRKm0zJaDY5wDKUBLN
2o3vgN2exq5LZr56Szmt6Z6WAvv6BTjhVRpt87Uu7EGLpZnVpV+oDA70u5DsAz23vpA4suGZM4yt
mAKEwIwwwc/o3zjUwRRNV0gAPDinlvq0AFI+EW3dKZTjmjMrbiaXqBV1dltE+zBVMC9VckKR5CmY
heooYFdMBq1tBKGnWm73uVmEvH6civQq+LxHfWMXySRDqF6W+2hnwHPNkuGCm1hPC0QApznOs7Wy
WvEa3ssqOLSXHNLQecxC4PmMr6lpbN8ApCL7+N3bWhzmMHs5i0SBbUK8NGWca0+OUuzJm8+qCsym
wM9pnpeZ0AEB6r/EAlKtXbrDsA6M+FoF7o5J0iNt320r9ROWlhySRhoWq2nvFngv73bi27jzqV6m
ExeqNGrqJiGMODehvT8LpinXh6k2XTf+fwWxkDEvjxn+dl6yJ6LRryR8pev14E5SmWO0C3GLwQ1Q
aPjJ3/Kk0HWk4qBSZHkY9R66Wa3KyOtlyBWMvBCwcmPvfwGNByk2ygPQkDmcWJ5jRNf55jqSHFq4
yKEheEm24yvmnoe0HjvVe0xa+A3exSzjkJlDq7LAck1pHSlvYDDSIOPXxLIKYmJRdcJ7HjvHbR6Y
vj4ZKBg0bVWRWKNYfl6/AIEH9Ck8BRpybV9PTO9PLpHqQ80EY8b+YiuSrIpDQn47xm7pzp0qT1Md
NTUHbsXsm/hIFyvZ4dVklMj9uPaCo5986CUeTSPUbJ6zoz9kGHw1+6yn4LXYtymD+3FHcOHgcm7f
ul/9gxYGuUOp2D27LwGo1c0VXjikls7OhZt8pqVnUy+8wMpPjDOFbTwdg16C0ElvYBAZGhK9io8w
KMEfKmkagZa0OHoPfjzywwMHtQ3QsKpR0JwQBGqefn6zAb8NAooFoE9wXo2+YuNgZqXfbBbS29yM
VFIJ8kwWv/f1+xkEE7ETQxOB+cTXM6BVinluo6PppSmy1J6iKgtvZewnCTSy925pg12qmpUfUBFa
cMyyC0m77H0d8nB7kcs5wyximT0Si8/VHjRdB6h/2+zfF51iFFk6j/JgAohCrQjblONqgGYkPyCn
eHvuC22FqGb0th9lfra6rZJYGZ+1LY/n+a1KPRuV2PNVjdch0RXYbimOZagsKrzByRW20pYtwIOL
j0yxR2RRc5H8zPDarywjjJPwYjTCgGRg5pSmGf7KlYKL2nS3ozSfph1H3ymcvZyDunwTzwNmhyzb
3KS7GLhyjxAk66q2aNlvg/pybfn+s+O7i0amUBXBaR/dxnunOslS0JHmrrLuUtz6FDPUNKVJgyOy
XyNc0w3vMRucLRKNiZGUTxItmlpA96lhnIve+mJlIfIf6yyb4KbZSMSKrzjgjQRucRm59i2Erc95
4aK6epWCO35zRpQydeq4a1lDPmhuEVXZDtN03D2zKCqeGOyVOcOCU2DzcfGJcLqExWxuTXw3R6Tk
mpLmAyhCqfELeWp/nze1ulb0QKwKmNwz9SenVNWJfoOa1hg6ni1WN9b7k/td9FhYqsHULZJNW0bU
3RwlzuFtKL161wmCK6xGU1UCkeLEopNMENT0ITWumA8l0zGGeePL6z9pabIFSxaFK5OG70ZokNre
hmoNk+H/itrsjfwbpHfduAQ+T6Zauiq8XnmMJKoSlZYrUFq1dONPKyAvMW9goEiMTPjnkBc+jFmC
Mgb9aXG0KxgSHV3E+8MrcMtwcWPPsQuh0URbbYxHOflMse/dsM1yB4UbSkAKRxf+sKowN4HO+wVv
TtyUHl/Mak8CBOO6tpIqrK1DPutGt6jTs+3grvQYMWaAcNZsSojQ2CBpW92nYRb6+FZlr0/KZO4L
s9uSCdY6ZoyfZL9wNqZ5/Qu1f0McM+W6+gm7Xy89uY/pRbr4qPMo84B1CF0ltp/fTgXW8VZIkwPp
/fipXDCUvcmE0W/eBNqLnza4IGZ1549uwtDWaSDGraypwZtsWbelDKW8FZ8jVcTTIm+S9g9Q3/dc
mHmQ2UaHDHzOcxmkKz2/1OeiHBM9PxMXonj6x3lHCIuyoJrUUTCaAFV2XEKejf6lFS/FTl7tc/73
vpVFUkQqRkaOyS/sjIb2/ThBi4D6Y0QlripQzN0KQ6snbh0UbMMFEjERzMuGY7jriAyZxj6AhZkn
yP3GdePOKHIkPLJo2tSxZ6U24LS/UUTatwEzQsm9eIrwciYayYUVgOSwxCc+Xz2uMfSEDpf4AIkL
uL3lvJ7qetCvegBWRRlrriGEd8vfmp2KLB1QMK+vm5uElwNrGbm3fA8nd5A3Mxo4mFrka2OSESU7
50yJS/1hpVdUlpJtzsJIkT7AA535+LMcInPwrAreFhlibb6tKTGQl34KV8jx/zxHZilU1MT0M69Y
S5zPjWG9mJtziQbbzcklnWV2elF97WqVBUarpbeJ4JQ8fOdaiHLkzK8ZUrP+5ij94Tr4V53YFVLL
0sKCz2WJJsoavMxhuf0G2YkSY7ZllFrqqSHesnNWuYNyDCx9QZdv3olRmGIf+wChdBlA4Mb30o6L
5Ekqp+I461H8e8inSMhEyrRVLNsHfbdOz1Ve1VNAARByWx26Hh7iV5AEZxE5nvIAt+f/Bmy/bK3b
GCRIhVu0iLTbgCvCaTuYAL5toJZ6klVdekhR/X1Ro/Jtg31ZpKxPhd7q14H1i4txy11IMGbmrpJ6
aIxDQ2DtXqiRSE6WEmOsm2IEbWLdCDRoV6u4fK0iEAV0X3JJmYT9qVY6GAFSZLvqs7/nuRoQCWTv
1CwvWQkFRtNjG2zSwli6CMyPJkXPup07utiuM/SpUZBSBEJXLDSPGpmELcCJXhN8BC+5DfQj3Cm+
8Y4lqMuA7Jbk4FqaAz7ZJZGwSIKeYgUAhXTgY2M8YybD14Pgakas9xl18871dObCeTuxjNFiJNgU
iTUQ231Izwbitga62Vb6xQa6vIaHX9Ee6fOpIHtbU/9L2dZK/kfm/tYzIFiMXeSeB72wwkr9q8I9
dPvM/cjeACz0fHfDuohUQqVbCno+CJSkoS0hyqMRTpMq6nqefLn/rqnHZu3dj4ntlBY3jVBN/mie
zED9SXWkejEcXDX5OqzOfJJeBwXWy4wRb8e5AMELZamJPahyUwQ3gG9OClG8gc97O0MaIiZ2s2er
lrWP87sFzmcvSU2oR/yVrG4+N3/WyBxyhEd/U7dE1TJOjFQHW7uOgZKeGoetfgjyaoPRMhc5y59b
pGNn5fqwSttIKJtHUwvaXKAZwlFwSj2Llrrli3wy082eV+Kybdw2Gmu9AXlGYmNuPntt04JdQWYY
wq/8P1kdEQFrfxJg/SWE8u38HWU5RdbfFbMJDg3ehn0SUm8oT+BB19eq1bo9a94TFliNqSi4oplg
9aqCy0ZPbdfciubSdc55Hj6X+9ALu1C/agpvLDgA1tuRbHf/2FsGNLSr5GBP3VRaA9ld/8ilqJ9j
0M2r57/C+Z1PxBz0sQzVIgFfSwNT1cVnnbPRHwAl893rHfBIok6nQ/BVWlSV1yjFWZCUoYKaDXR8
Xzmp0xfxGDMeTxYsvHT+bpqJ4mUpiZQXlySY8gXIFtrFf2GP6bhgB6muPgaASbtMe/EU9UkSnNH2
ZpnO+SjqJbRyXzmGP7YaZM77wk/9rYYQAC+cHiWAbWgWxSzmKtEAcotjjXrbHK+4kNLfiNYvxuGh
JYIHF0Vob06Rm+EwxTUpqO5Tr9fANbF7Z/Y6s9KTwIEESnqtVbFC6JewuJ+RjdjkYaopjU4Pp970
Vb3D5qRXhXUIuGJpGfrr1CSYNZe56htspAU9H+UuffRpd5i+mZYBybLPQrzui2YTQ15CwE/sC8Rk
epUemGjmjUtIpYgXThQ1rfgbQH85hdxL27PIzea8FXrcXGGb/7UsfbaOSbuPIlTKXlfh9+5nzTwU
tqWetxfuJFbaUE/oh/GKl3qtkN/60uCIlfmJs+0Qna6hiii7wlhSee/f2Q+2XRKFzs8rBdvJz3bg
HqFPX5skUxxtbLkQA8aBx8ambNWpYduKBcSdlZ1yZX/A2aS2GgPAqCxiT6a7yYKOJF8gamSwe0xG
aXJ9yTy93iI3NtqAtnB185KFoBvJqkwWYaMH2eA6GoFF5QXpGA/u1DgkWkbnMnNNVuj4ub5Z5Zqx
u0Ge64f5fYSu+qucB3dzDMKpB1xfMqi8ZbwuPftvdNJjZyP61pH2X1GnUDsodQ0o/4ZF8nJgti9i
y3w06Dk/6eWRbGjBaUPcPI0MfVUepF3DbblcmYcV8fcw0Fi91swqTqkIwr6isDlhooTqls42C5EK
iy6KSvDPKpRkO+OoUzVs7YBZoiSeBYVkcs5BG1mg3b5RCCJmkGCQ5XknljUjZEtepERjSBzOYyRP
qykbZrffkGHDZyW/DDccgoashQxTuzs+Yqkh7gq/ojj76Z3kPXupA2TXtgCZ1oEmOp+EQja4KHgU
RxW5t2jndwnN1LrZiccCJeLvbc5oMH4iwnHpchNuoWv3XUKbIqR7a0xhjaV+icb0kT66DZbUsiFZ
gCq0mduVimhMIef0N4f3V/KovLxe049AM5B5rZNSZuUH1LBCMVjuBMSF2F2k5VVruoDcdHZMJtHh
z1Kq8Nj++CKADArWbAUWPcuTpbh3cPh72CP8mZmv8bHnPfWeP1uB6/7s+ehObEWO2OdsgDrzOy8d
Jw8b3YgOuSGES4qkYI1ngY3Xph9S/Vrg2dQYIIXeVdFT/NewixXpQPTI1g/WxGxhfeJejg7Qu4Zf
CbBZosOF1ZjC3mgyqW7iT6fCyU+RYMR1dhZ7jf/f7Kq201jqvZjXlXhxHXO3FW9AqzFievHFOdd3
hO/zSwJoH3/1BzGiVt/JJKcVciviHS0g2TtJqE+kiiyt8SnDggyCfo5amobfGR0m9fGs+5sTizMt
c9YAXg2j5rZXCGslKy6xSO3G26h/l8CVfl5NTk+IU2qiWy0KLxHB4pvDjy8R40KXTxSgKat1HC+k
CzCTa9YdPpvFJnJ6XAux+C0NHs7li7ZlmyQqkWnPulNQMkiqXziNrKBzf4LYjqBfKuy3ibtZ14iB
TMJh+Day+efs5ZAjYmTdlFCDK493DmfHX3yFCiH3k4KIvTWuoOVB7+guHkCSqI7UyUAP39Zo1C7F
y3lvKcB9iAh8O01GGpLEWvmJFYeeJ++ZFlNBOwihg7g5kVlSYgYvLefKq4Tx9Cvon04/XkBa4j2Q
fI/V+LXc1yTB5fZXIn6vcgMRAOZqX6rSMmiF8RNO4p8OZt6O/zAHnJ+6sVd7vjR/j/0hiHrlGqr7
ozNMxphTrbV9KGOBQ8z1bJJw1yTW4eZtVzsGYcQuprNfo8+l/28LVPNDnvZPHniIUb7nEAN7llzZ
hbybI2OzHYfYraI0aGaYNbywfAk5LEIo8vRdV//We3Xz5+jeRHN/xGCcJ5HHwYJXGKE55bkDannk
t7ABdjvh8pqPLrg8nNuAXv0mtbjAkijG3mbzK3NExgRaGCBUqm5O11VE5s33JEfijZb13ESDJ9Pg
lE57unbR0a+mQLdBKL04j9+x9Bnx4P7ekLKU+h+oi5L/IHbFql4rEjQ2WN3TfpVl/r+ZBlrH04nS
wMUoqW0So0hLH50k7P6pikH6PIdOg2vd4Jzds+VNqPrUuQeqK8YO4cEiYRfZbNq/0PnCOl22lTWx
zUEuZm8AQtGQ8MYwTuYvJm44F01sRf38mpGOoxK1i24FODRxs5GKDz21aXDTiRyh8ZaEVV4A0QPy
iFZ5TRVbtSlax+2H8w6M36KVYbD4b4Uueo+jGonTvaNkklcMUTVbbbL5tI9mnnzR+lc4qkTOxBvM
AH04hBGmWla8e0uJBAgvPDjYyenpTyBW3iv6WhIGeC54UUmDHWwInn9uNiohlKo8qBdlCjF55zMu
pkJ/Pf7y20sIJqUPJiniaJfjr5yI12Xet5IaY7x4jmmZgQ1L9en8JLO7+5KUujkR1tEL2U+LGoL5
lrvmJUqbOcAJmyjsDJSjR4hJoHY8gssIwTxx+7eyFsVD/5NsDn9wTRmINnrEn/Lhhx5J/UOrFUQJ
93GOKxOAg3b7Q805Us6IgwYAx48dKB7n//n2TU0vbi8VkX9RBHg3OvyU6ktsvMDv62eTk+heWOCX
GTQQhRg2HwWWX5/pKttfrIYnUfU+wW92MJuzDelQDXXIGyV5/l/TkxHjbTdY7WIriRTRIK9/XOLC
zWEtuKAbLOI29Q762ZJ+nyyxTlpRj9+vwzTJY5fdJ9BCgK4UoVr6wqKwVkevlau0DdgNiSPlXqd+
dcydHLRWhZR0zWez26sxnqwtjrh/pQihsZph8vut5lEtGwl2lvpyjVo8UtaLpmjRGxuAOi+xj3B3
jQ0/aVwYlv7OsBp7SnQQZBR/nCRNWHUOUhAKLpRsUJWHXSTk5w1fxld4quzzp6hk3Ffi/PpYKtW+
adpt158L4ZtXwVlOArO15iO1bPYZhhoIvj8yNi/R+FlxR7FMsV5crGJCnIg2UEdxZhMnPV8pOKop
yT6uKmOAPwtGPJpgIMaaUDJbtFga8VTIegA3heSkNJckJhyAwuAt3MgGQYlrDuYaotOievVqueBJ
0aihNv6K5xFh+ouLqXh7Ii+n/8xDgNKleDUwhtsGwf1vSje9SacmqQuL36NTK7Avb+fiWU52Na7Q
S36fDy/Ip3rw7AD9sKcQX8/gffLsAQWlxYoDMZYmnX7EdgrkzAWraHCYLTyB04O2JC3Oj178IXrM
FZ6HDo2rmrTJmbHhlHMXrXGJ0KFd6GvgjHCtTnuvj60UiGYlAjhFtVb6y5QyloHP8ZNjXyZLfuvJ
V+wO5z003Euok/9YNa2WuwgOEHQ4+Do8jJboNsJKKT849mmw4EnMEi6l8w1och35EcsOYHQaO7px
G10fJu6vqU45mEaH0h6y3YZJJVyn+o9CKnNLhF/Zg5SC9Km/uGAB51ZXhQvSZgyPrl8kfr6ZAwH+
Ap78qr9iaMXwrrKI3l/QlHMC5rzdFDGt+enEQjBrU+3LWJHTJKQKWbH31CPnxK6EZx3SGuqfufUP
ReIEjhUNXSy6nTXlQXH8jm+g2giLcqLHMhSsYDImLjTxmUk3hrg5pk2L2go2ghjPyMW5jfP0cQt+
OpWxARvMVVpiyRoARjl2q12LdU9hOtNLD3b4S6XWDpAMUfDvgT+O5ZkktsWUO9sGoNUwTMlX8FJy
9ajSLC69UQ5lxkNL7NxnVKwYIOF9173Yo2QeER1CuzL+YvZez06TUqiUvc/EzAt2A2Y16d5AJBbg
ofc9Zmyb7/e7Uqc3zF1eB7aS6Y9FHh7yuRgEflG7i1tHDzMNA5/3tAwE13z+oejEubrECKVkp1ma
LksQVjzyEt0SLC9YHGo6prX6zVXRrCLHpN/ytUn28Z6g1IAAEnVUvSSImI/u+D1gKppKqtVdbI4V
pNxaal57M4+NzaJScTUDiuFohl8hvISeldwnr3cW4MSn2lgPDg39Tq+h6zzveC0li6mV5rAhCxSj
q1OUJqvf/QczzD4Sxc0vbU/LbPpdAzUsgBNbWTA+6p8ugy9b8VOQ0fY2G51XOavEnw6B4ijQtCZU
C/7a70LPNpfqEpaKA3p4TmyY4JNfjRwOwmZx+DsKdb5hNc887yxyMcK5f2PaSQFhoiAkZn7o6/KZ
y2HG6vDLZODCF81fjJPnqjJ5m4Tod0b5CpcPD879E1OT9+CfDTkZYRAoJAEsgssIiirH9MY4dYUs
OpbJDuUjhBbOQMfDfS/0Fs+7O8ub5GVZ/8nDupjZZQinSLLQfMHX8uIm8wLZHsibAh/5EhNB/gLl
DL7KcEX2jd0rzBgQO0lPHpGD3QCLTMkx1Cn1T11tAjkQnCCne9xVe6NPCGYqBv4FWmuf07OkLyA4
c9Z3dbQHyHo8MHUs4Hbarj53btlTiSdzkCKEQpwobYGH5Bpao+FeSGvyFIpPZaNPh/Gg2fnvvzZX
1Z7BetEDwxxF5dJnVz56bTCjumrbwdV0a03u1z8/OtT+Zpm1xAUWp8DtYImxmY+0uQEymcG7VklP
gjr2NlG1aFnEBTh2Jn3k8Piq19hFoH0BvmeMemwfvFMB+n3BkfFHpC950lR/astDo7/1I2hkb7x8
FOk+bntaIVUCcyiBOYXCokM3Ym0JSk/JNWVvlAQU11EQ+iA/ocqueSFj4SWNgMdjCGhXBbQ20wiW
KWJU6B5JgGdJOAvN/ayTXd+oSxuHqzlCPbp5BXblg3qEvvxiEcep6bdLLPWMNT4WQpd/JVpLrvSN
W5NpgmzmrpbU/Pn3QeDpR344ykTnXVxOX/6UHyOcPg9uLAlw8PSZGoMZI9RdIi30coylKd8b84Mc
TxakE/m36jUXf342fgE8yUiyMMmaqRl1W6pr5oPZoUEMX4t+yMdle63IfNZGCv3hTECMLbWYcfXq
vYBYh0DmoNJ4FaLba2F2W0qOwBlwL6ITCC6XsNYfaqh199zfnUnFaypSkHTTzHUwYbUWGOaAFceg
vKfkhY64GHHGFdRGqQOvB4ZL9xk3osMCUrImdlYfw93Wdz/R1ckCO1GJIMjI1jRxxTMzk2HUs0qw
YjFO/gtUmsLiO7rlLCMjeIn2ftl0LlEj2uS8hW7UGmxDLDG7UK68bquM2YVHVyG6NoHvVGFHDi5x
BK+uS+p/Uab1kgr/69AbMfS+5+hdQfbdjHNMQgQ4edjPPV38UvH/ivWTgAFuqfXPkEMxp/SDZLeV
e35NVBQnT8wkoE5MTjWLEtbZdEBHaU547yxm58zZC1FGynKrqswuGvWym//WqFJerKNy9lrE7LRH
/0Diyn0a6u3kC2WLC7GUaTZ+PPg0085AurVRPRiUjewkbcG5lK38X85iGYdl/nqYIxn7qfawSR27
JiCLj+qav0av4Ia8FAr4/j8G5DHWrgLzP/sq/axGiUhpHbPrBV24UYGccFf/wTXq0qVT+sRENvFj
V23SGzgY/lobMFttPe+Xnefc/ltXK/K5idM5As7/erCt/Oa/GtOLY4yz2H1T5OySyYnEo6RULbOA
Ine4W8McELlyNQRL41Jy6q7xdCVCHY3esskHuZpNvbD4/OSsnw8V5gZtzY23m2cbY98QivbD0F6w
DMxk9Op8AHg2/4mzaFJIAGLDOyrEjVUM9fVCRxyCv9ysXoPmIaE6oyMTPZc4CTLoovumZouEKT6V
n3QTw4EHLNqHQMB57Y6Zbu2t9ggh/OKl7sv2mC+6isSAkeE/pIKXHDlCJUK+rVuaYE9+4xc0ZY4f
F21stFIR7ThVxu9UpVk07oAGbl6nOsFqyUychx0TZ+WZUHXJ06GMci7b8o9zNwI6Zv2O7o9wg5NR
riZ4GzPJ+ozcoBQYqHVtodEJaQPuZedxpxVduNeIZiSew+WmG2zMUtxT43czL4NBcezYxKDFO7LX
Q/qkAMIpKsmHXI54kdYh7SHH3OtN/EgjX+F19v+Dsphd+5lmb+janpN+jdrQb9A51IEVrkHYVRrY
GAGg9beVK38dyrZWM2PcvEg28j6Welj9eZq6uJcWdt8tqlOcaX2RI6WGx/hN3SNPLpDlViIr4Xjr
waGxg+j8b4ICiQB8kXXAoi9+NUdRld9O6ktaPr1jBaCkelKSOldjYi6fZMR8/8LXbQhYya6/pIoU
1oXK/LiQasOQGrnoGMd2LSQhVBodzUsrc++8FQJB2f4y5iK4RL1cjFfc7DBFgBvDvmmkTMSMzGKn
HhvbuwYTRe3oxsiIoyAgCa2BdrTbdUsvy5jWVrCnriIsf95P93PfGwYSwY1zuw3yK8PXjDRofJmh
E0b4FYlQQo+gr1Le8XcJROenRzsLP1Gn5Wdpmn5lJFTBNP72g5BfCgulS+9AmvhzxqspMB71h2q7
KL+KzSLAYyxquADxAxYKztPyZo6njr/HsWtMB1a8hyPf+Jni+hFVfYTWsP6KUtTZBEN439lIZZoF
PRPDo5iHEFlxWtvA7f9NGnA/gbFORAer0+Y4x3TmOUmRfOQpXzKyHjtMy/XTvgHOumO2iVx8fm7I
MAGwSJ+K1H4yQu8sBxPYaS3Eq9Q2Gp+TjCrYW33A/SuppkSd0AonTerQhZ+9BUU8SVAorPk0t6RH
mGdb6CLsCr0Ga7ao9PmEvTctqTbslRr4ftfbILJBfXw/ef03OwndpHsEdK2emXzVBdhEt8lzBnaK
0We5DoaxTftSANSvZRdug/OdChdedsaFGEbA/rXObvSPzgPbaUw6BCaC1O0jFcHo/o7D5ovF/aJN
IR+L1wIX8qAPWSQM1okQEO9F+pOdcU3ybN658ft+vxo5pKHFPJhluteKm1Sp1ZuA5sS3CziTCeJM
wXso9nkKJOGNvBN7jr6LYQxOryDYU5LggC1HFmsbWzGF1R0wViyxPSSMeaq/sRRgCbE7eQWeQe5G
H7VwdcxMH18cKc7yHFvhxqzIHFB6mCKGNFRbvP5OxigMMptU0LpHL8oXJEneSNgcr7UniijzWcPh
8HKR6cVkh2fmKIjqY2kfVhxxQf33MpasVKvmqpbpfx7FphS4hvz7CNoNHezyQXp0MBqQ4aIB81k3
8tZ4vsjG9pp0yAFtLyfBVsUW3L8F0dbuHQHG+l1m3/btgtevnsfrk16GOvnKw+9ghnAPcoXL3OrB
gShHfBKPMc8pb3MlUlJ/cWRLzcXav9nPOeJghPl0S3PSpuAoYqo6/cMwTjG/tFpoyfH1BCJ5GMG1
fX77y9byPsW1VCl3cGgZWdp9gmvhy+uvv1hueXBk/TFLDyJtMIhuigAbv3pjalwO/tzzABVR4Dxy
lkIrG+PoITaVeMwCHJU7PHgmVgoZK8q6UOeVbPHYzbH9Gj4OoLjZVCPhYeirSZLrzaID6BzWGaqO
I8FC2q2kzmptjKRMEZuNJLBZ1umoLb5K9HJG5EHU3oEL710FHugkGXl9tydWEaXDl3jNakRVSkFm
sfXPYOpmFCncPbu256jJxdzHnngJxKR8DF969NTeclPKuYt0Jl6mmjJDT5MoW9rNg8P0iKC5NdQl
6zmYK3BTkeKxuG7W3vhaYQTE1OixrxIYZDYsFdiJ5ahn7wNkZLxvwjUfKz7PNWRucwzUSyw7Ob/m
kpEPcms9JC5dAfExUAbO+C6kujM4N4rjAtHZpGZ/SVvFAVeN4OTZX2lWXsuXMRnFvUj8v2nro4wE
yBhtOn4veiHWjX1+CqnEpqsJufPy7smjkSL08qjKRi7UPuHejmtDwfujASPZL8rQ/gm6pg3WDGSN
6yMZJhbZGP+g8fQiiJuYd3E9VntbkRHsWOXhNV9OMxcB/pswGbaVkQbnKn70akugKto05N7OkboJ
OppYSQz0Zb6XXt1SrTOgA63UEafg+tt3Pmv/04wcq6C6aMr/hQa5/rJtfOsT1/TxAWqrc9Xoi1BO
bCpx/lE11CVwtm3nIQzG2nhpPwnJGNKtdzeiHqJrUs7NeAEJbR14YxA1kTHmrRIywaB514gxGJJZ
jWYBX+PiMJrbJo5M24JdDTNPvmEmxY/F2jpDuqC+YCx2BeKkLNKz8lKuRsO3rBVAGlVu610dt7Bj
MouyDntVVDLOtlPoCnBNTqD3v5oEKl9wqrK4ArIwsQYxEe/gG2Hr77tT1EZ/KcyiY3sWLbYGJTdB
iZs8mWiI4N6/oO44gunLAW3cPqRvxbcyMhrdG9MwPs0VssA8dtch1VCqhr74+/4DrtGuq4Eexaq7
A+bakKIQxrKQJ0QysiKoY939P9S+atZpgq3qEskNxDmGMFZtsSpceeyGJgtVz2EgHRD1J6mhM825
aeZepyLnyt5Naz1a5XbelNZkQ1APAEa+z4k5puWV83whRsQbHXVUWbEwZ9s6OYQTJhCjcfV83ZyG
c7DKdU+62ayfuW+Vaaxmxb8oaNKK/EDATqwzFR/ZYOqua3QMsbxALEkwpPlNuxqqp5EipG/G/JOD
Kg03ellmMWpzCaLPoYZ9dCHdc40vqZCN9IO2wCrdIogBDs4pmj0McbF2gEVPljAHi+q5xPJ1EM/F
rafKHJI7hq3E/tbqDbIF5sf7YIBPj01oL8I4/1fH48H4f7F98DEmRDKr2g1iFujyxNSVRBCoZS/w
01NBK8oDwUJ7MlRUDMGgvsHTYJfj2KYe3ojOmXS9V/Y7zFZuk99STYQOIYjbauB4UZpp9qouuRip
hvsdKIaifFNFxobjBmsX1gmnwD7TGEepJMQdb+UBxvdOy3skA+EmFx8w9SHeWnupEEr4J20vpVd7
DSsNetHsNxQb+nhfF9DjudMmIK2iw2IBaaS5mzw+oxRQrCjrW5TEUpUzIBAlgFqE3OtOga1GuyDR
iEzgRYkR+3sg9DeWPD87IA5KItQ3ziauUpmOvxaNq7t7hs+0RL/ETivUhbDECcljO1o8NJARHqL1
KJgB3irH6VQQVXvDDHvj5bhZtVSeTcW+VBTvtEY738YRkrxJTifZb0CPlRPIHSzVEJsWZCDhBLtT
VZBZ/cktNSkHNP9E0EYR0dHKHY1SX36h2Xf9kRwk1N8RpEUVJjR0Qg6mxbiMa9UZJItEK6lEuMT+
+AJWQaSYa0O3rq0nQTIIEqAsbqFPkXEvDFX+rAsA2/LUvbu2qYFAiUN/FP0HRD7e2U16xiiQp7YK
akXaoaOf75xMwoFICcRolLKC6/cJwwijlR4U86V9R0wFpha8oz/09BeTH96rvvZHQK+DQiFeelo9
0QmZ0P25UoSZWTiYiM1LR8QF1REtw13GZ1SjBTybiYBp+VlgFMqptSgfiE4npeW/AilUoN+LUY4p
dw9vGFEtF6woVB3z5v9471wewn94365BiVvEdDgC3V+o8sB9jCQMc6mcTDPb1gRGmyg+faPpsAte
8mlnrgO5qs33ctFOz/jXHJ7FNb/hXGQDwCbtzMGo1OetEh9spnNNLy1YqqdujhKCm1nfs2Lky+AN
ycfy/j2v8fxXudA3Kqh1xdj9PAWqssRIHkLZ1wTF7+d5XrzfxdPnDYZQohqtlcDsSq3RwFdKPA7n
FppLEKL2GQwn6HilN1wODeb4AnmATP5/QGns1KquteXmtQBJAECedBDtH0s+ZAvO/8oY5Nh75e1x
BCh5v/XcYx9PWuzJjHPAkVcttnvP9x9GtuhBZQz2U30adUGYgVoaURCqHXJ8kiHXMkgX32sA2z8f
BVsFzQuGnsYn8USqyLxULHAP/yTmyjwaO5h9ks1zdq4gkZRGPBwVDxL59Zj38xlcjr+GPxK0Fl75
ymv9KO1AwM7x9pptxg4LkceqVw87Tz2+lvKPlKeWRVG7dCFeM2yr8XC1OTISexXuMikCthhw9lGG
bAcVW7kDGsfMs8ZX2W9xNiayBDIwiy3jiAsw5TmFX4Sq1orlqoKCE1QPROtZasIhy+5P4g6HFJmI
bS0gCiwinisGOJ4rKp9OK8YRetiNl9rcCBHqBg/EIK/VC2oiIu5fycwnf9PcU7MvKnWYgykRkZr+
4zbDEhR2xZMR2zKeUlLoL9hFXF6hyw1hRnqHZqHbVv25FhTcvYWOPehJtplWxnQZNaclSz0JVrYl
7zcTl0tZXhTMLO5rACsce8FzUvpXICNeOCFG5PTTLyEG87WIDhDWIa21Sce5kYVL7DymJVfgfap9
ioV82iGuu3syLLoquuHhlZtUbqrHTq8e171D7tc00loVuapQKX1wOdFvOSutOoURSY+48gV1lZZ5
bKhf8UiiUYmU0ArWAD575WRkkZ5ikjixK96qUPF8geQV94kPGvAc2zlh0deNgm4t44WPt8VvU6gK
xyHSM9rjGPkHIIqnl92ac6ku+QBWmQblJyfXIRq0FA2BzQFc1GVLwDl0u+uT/QHr1a1nNmrnfq48
JvVBs/NcsHHblzJ8NFPqGgSayEY/zVBKcUELX2Xat6eC1I5eJLnw3aoGnKuujXNcphYAmg1mucnh
QvKes/gg4QhdIczy2DRY4sad5OBxez/JKQ2BXLYfGIKBeXCTN4ZkF0C5kvm8VNAFZExrrjbQ2bw6
2HS9TMNpS3Zk4kuDtWTBL4eXVb/oQ8ZsJmtpuVzEUihnPZQCKJ2wc2IzKqlabqFod+hRC65df1HR
kZpzrJ1yAQbRTJDcZpUSA7k6QgYs/E4gWnAUroUm1kWwPK9n8tq+t3f060U7s7Gp0H4KDdIYmFY5
P52RZPYEb2rAtEKe9jOskTvNHP9QwysObltpjSkGbx0NT+DAm0vOcpRCer0NMMIp1qovq1JaYSTM
8WpnAT6VoOg9Bw0QRPbILWyOp8+hdv44z2LL92DnAHIH9bea3cP4mE/xS0hQRJzyT3us/JB11pa6
RTF5poPEmGTsYwA9vXW6o00s5Pa9fgfiBAaMCBHRG+nmLCL1nF8nzknIXP994NepLWjSkWAnPwBe
Ou6rJ6fYDAcgh3LyCH46aEm2WOkMXfT0TRpb0ybeVvtRl+oPYMZa3ez59I/5+S97lj/ZfgdWu6Cy
BR0rqD6iaXCeflxVjG56pk+AVtF3hQwgC2GuXcerj7hSSf6KX0wNJPxqeGCCxoVft/Q5St9rVJXi
6n1D5T0ZqRL4qO4hiRZ3pvyaC+zqtzukpcJxq6EG3BBCGEsvBuRUObXn+6yOq5BD1Eok8KzW7Ghb
pUf+xcH0qBiVlu0yM4eMmDZkBm+FY8B6Mbicp+4ilY38mGId+sQ1h4bOWOrmy1BAGAoV6wiwjT26
viJEaKNlVd8JNaiGna9TfOC9kpgjQml+mPS5ichpmeo8YOjuAXIA3jhkrqryifL3s2PByzYrtKUT
MY21g/XApzZ/xnQXb3B4b3zUas9PvhredPF0SSoaoGYqvE4hwDUPQg3vQ3YWcq5PXHWWaSlG/rfl
xA6K3lIQnEBOlEnYjIJOPGpP4vOM9rItMaoywXixmIN813SMLrMXWIni2dlSgM33YnwQ1YplIWgg
DO8cJSIybtJVxqm9FLq3TfwTnkVH+sRIMcwmlYCiY9aFxf1wnbnDrjuSzmnVpgRg5T3AnwTQlQke
QA391bBpOTbNmj6w1VSmPcucaMzqGP+Gh36Gi+fE3Gqw6hade9zc2teqim7l+wv3+EyHFNlsAsTy
mXlvIdUjQiOFU/FVdldPM6NSlEx3q3ARg1JRfxvzkFb/2hPJgJPSd98f9JzIlOJCS+FSBdpLu3AX
3nkmvKimhOYbnlzaTMlzwSnqixeBF8sELNS2tDJISxAiCg5oPUqvzhn3cBX/D0+Sjvhc4ZOCg4Jd
nzrH5Z0O3D97inmSDPvNPfl09ThDWQO3330Ru9DFicuCKYSet2bt86+oCEFOZH3ztgTXVG6HFjW1
4+vxtsqlO8vFbLeDhx1fB3Me4ofqZ+apTfQxGRRqRR7q+IDHltoeI3iSZTmvYQcSLgYCz5BCybAd
YlNCxQyPMERVfj0zIVXA11gM3pE7zcVTrChUrTe0nMPKDlER36Mvar05ADtfwMmTxVuYFRZi5/1z
Aflk7JDak7zb4GIZ5QNQGdtq2jvz+6LdjMK423FiwumXqnMOnw3vhQ82DBVLWES16djobp6glUUc
nWEulDuv08c8LvpG8SoundHIQefCLRaHuYcPNjcVf3RDeW80mgTAEWWPDglTsphO1xoUZX1sxmD2
k5OLi8lBCesbQdjMCPfrE3Zc4rrfVI0T8gjCmI88Sl4POqgyKgIXxqaRn4lhwz2P7kT12azkP690
JBPA5Y5BoY9/JMJZqpFc4iOzxJV1ll9Nbz5ttwsLu7sggczx28bcOwHfjxitEk5073lU7Pd8rzzE
DF7W/0OIS8Bb4bEY53I4Q/eLTpwqhoGBy6MTRkU66VmYNnVYPHd6v3Po6OVqJKrgubxfQ0h1kPxC
fu0CHHnsDoV7BxT15qFH0qw1olWxoiqh6X2n08fBno4PYTr3IAOAouvp3Kt+ZzlYXyRIC3h0OgGQ
BjTny2wMCdGa3znLeMqgAd2nbz4MOVJ599ujCfYFbZBlk3sKSL9ZoxMhIXcBhnKaViu00UMJkpZl
g3hT1gSxnKd3Voyx4ZzA4k8UKbKDXvHsvBBwMKhay1yGTJtdkvlBAlYmY1p64pw7vAMvP6XfXDUx
HXDPd5EylhDA8A4bQGYx7NdNJ6jF4mOsHzKMtsFvSJbOb7irxhoWEtrd43zfFC8O06JUpPUiNmyZ
hZg9NeuE9eK75wGTsb2ROXfkkYbPMApmI9OV05irEsTdU39c4ZsLDTsi8L9oXyQync8mMKrgAu/H
8B2i0wI8PAin64MdUfKCyDsfnYoCawKcwBbPpAXXrOF5oXpkKm/Tb10fhdEykAVftBoZAZPrYqF4
qiTLVOPZUISV/DexjQoWmpBsoOVaomSHUR6cYLj3D1RyIBZu9LuLCDg56NcfHueHnJO4VXGePIy/
PCjTowolz+hJHVUgSP+ksbD+w9v0BrX+iQ+zMXwTeWv8RUXLZnmjQFc2QlrnTLJ4EA3yj+NKRtnv
/kZcvEEbuZGDJYcZ6qlgR2lDBmWuBy024o8IEzegliwioZ4VzEiS4oGbcgM1IX6lV4F0IKoCXgns
1m1gbHN9AL4tJFOLFNBDGiguC0MogVrUghfUPuiv2MdIBsqpbGnzCOTfHln66MKuDg0LEBELcIcz
Ffksbc+qW16mn1KYOrYRXV6ZI7Wry8MPJVuhgwQLEoaAFnwcJyoWXxlwZz4b1F60ef5hYBR3mzMx
EBRnojRypy0TsttzxVAJ1Q4pQ2SADTQ+iE43bNZt+m/3BidhUkCC666fd2THgc5vjg+vJ01hfoGj
c5B6AcFx2AVqLMknLL7IqCMcd5UIJ0umgEUIGUsrzgrpUB/iYdYEykI3j5yYNVhFkhnpZkeUAavT
wSXjMBp1gJ/0aLMXbFtxdRlprf4clmk2ZrTXRF+5SPr9KvABgNIF6GblGk+npPaBqY9fJyvXYEs1
YHjJlICYDz5Dr+qoRKhNAiDhAzrbS9YF6qspQ09BdCwGsuoKBvisBA7x+EYZomSrphM8ahh3uMsa
7vbmiigmIv89tnzxo6AYKAqNPAWiQPtigdt2iZXZ+5fclNqEKp4UTF4Lu/VKxYQmX1psydSYcYiK
S6N2zEf8MNZBNANHKmlxWS71RoEA6/dmqYSvOWKuN8bjBl3EzStehkEWnaR9gPpK0ZQS5AOp9hEb
7PuzwdaronlgzM2ujBV26yE7C5uO82OJwWc9hZ/p+xxUTGauf7xWNOOn+EAEbuRKfIxGqFfC/7jJ
eWOXeOio6c8yt4aPpJRtXHUKUkNS+dbfC/bEC6UCRqZplmpIhHfCJZiDNRZd2Zd6i6Y6FziIT1TQ
adjMk7l4wv7dNvAbi0fNZjdZBCk/ZccfWQE26N0yVat5pD2spiQcugS6A27M4+UUk3sM2XUxWqPF
PvDpfUyyrv3vvlakEJym0G1FdMaG+XDBDDfmoF0m26BQPYq/Db1j/iVc4Rjx0Vq0qG2y5jnVDYRP
QnuTbdFHfAEbreHeeSHlG9YlmeArsdtOFs/mhDSUS+y9bzAWCooI9oYIJcr7H9GSMF+Jl0mARF8A
VqdsgQWCmcxw0Wgz/fyYaTf+3Q/zS36RYqJHSrAmMnpfvAbECvtm4YpvUEx9+OCWHf6eN1MsnC9+
TEN8ziO2WxWbDRvvDG6DR6HxpPHaTzaObfWAvX22LPF6ccrMJbjJsOXd/+yupDHFQAQl3c51ymOI
GSFarPcnzSJ+SUBTmfnzZol4JCwKZqxKcyuwKT3H5WsBT5gXBbLrTfg6d13Loy83s+KFkK4MaWpo
AevB1J1CWYv0DgmEGo570EAkfKn1sZeDt7Y5xirkwnj8Wqyu7jO32mV+0IUKhwj59N7Z8+5cYl/U
oNLym6kipnIQ8Qv9XDkERpHzSYUuI5cHuaiKjsrfSr8CKQG9Z/2Q2AL+dO/ATwQYHkFm9yv4rkhq
KP22v5at/jylB1JMAZqaabcJFDA2DHpis9zoGtovD3a0MeNAy/Synugvb8FnIKxvclwn9OWFmT52
2+h/Wz8WJ0jdJb7WNVN0SFL+XPIFWwht2cisdDjZmQu5MBwfG5XN3whImjF9Rze3Bl7bytksGBKW
sopOyhTu5HhNIgjybItzjhN5fxuY30FMdACtnoMiJPPZiFIdst3Cm+M2eNXX/swKELbsru0MIF6l
bNsV3wDxWOgN0ZAsImZNKC/fbQriBX+v297JOsybPyJTf0XU+FUVMAfuTKXoUREjIMLcWlaU8KZr
t0P6SYryBAjUxE4MuHqemEQadEhxBBtP5wv4RZ8cCP/TYHfw9H6pk6ZOon+ooT2YUqXG72Y6hMO/
OCMkec2QIEN8y6kRLEdbFNErfWzXyzf3HtenWdrg/tUO1lXGlU4oh0kARuGDGR00T8DV8aycQJnP
1CncZiDj2xBK2DVN5PkrCjZ0Jl/CqFnMtfqjhIAkdxIzuL2eP6NVu56qHAQTsMBbvXBjOGcgY2X9
melzG5p1GAxWtmAY2x0dPLR5+xWR6UoNh/agtI8grwKPsaZphaFaZXm5h7UE53oLmm55dRXNp2a+
5Oi3FQiS/8pvnRbtIMb97Gj4QX0gXjN1fvPPYt3/qkg/PSmCIQe2xNGh4mqLaGPTq0qF6d/BzWb8
lVo9/CwEGXw+Sgi3EkN3WNTEuwDlz9eZ/GIIWwIjT/PCz7KWCh/BzLgUxrZRlPbmzZ/ddntGp+De
ktz9CPoU2kbWBCLdojH4sK7Ffi7I+RIUewdkvQ72+Txf8wqfEcDZtgSqzWcN1kXYiSjPddfRNszO
RGVVB2KPV9CsVru2zeI+RePI/1SWi20BcLMPbBQROzlghd3Ou9roTlyfJ+sq0jAwbP2gJiJFdJR6
p65iyziX8znuo1K4mPXW9fYfj4sANjvK9lw9nsj3d++OJYgfj4Yl+8b9b+v6UoXD8ZxpaJJJ5qyL
UprdqRa9iqRt8T0H+Jn7n2DeqnqJEFETb+23BnLxf2jL9w6ovBNaa26I1eVPkW01W6vTJOCTuhxC
TeCaiO4s5I2+dZEdwZYYGGG79/vBq1Atq12luNt8pF75nzpo2n3Yb5wMHkf7e3yUwserZd35QkP6
l+MQGY+rOUFYpcWfPxb9EQxeHA+qL688A6k6MhRmNxNLznnYOyxWnTwD8kG8o4ywynKPfVb7VO8D
QxWiKc538KOKSsDIwcTGEHtu4K9UxF7+dC4BDL6H4XuTGhmXn8+P1XlZp20zkxcUnqVrVRc24mYY
UJH5VXBzFlQJqvbhwEOlk9anyxjxsnuvVJD5bgKKTvpGXLkP5rY/idZg2tJThaABWdDcrhUcyRMq
/CaS/FSNCUD7/tuKqRuuJQUfLLY0KG1S3eiWYiJFb9KiCKSFZRqskT1mBBHtgCSFhgLyHj60cRxO
qGRkoSVhFdymRkWxU+lwa7DLROKrUvTC9jpH91+JOeQtHyFS2EhSigOAvBDiJb1yCxx7yyjkbaWF
oFkfQYYOPlPd/+fSAqp6uWoDKA9thruD3FE2Yg2bnr9BnNT2ocwU8/Fllf4aT1wFQpsa0Cxmp4ZG
H2F8aU/Fm0ca0vC/JW0AIWK4IYTD03trNTzcsJ5T6omEIjNsm0/hY2cu1fQGeC5A0KkVSzY+d5xn
W6gXJnDwBisKRvdNZWUhOMJTbQuPfKbw71G5ncF7WxgFkD93EUELziFmld2CPQUXBdHT59DBR495
Y6XWrPpsPL7Bbse9rD1WEXHiuAVT1tuB2kiWCPza19DNlavKLqkMtFeaPPJmK57PNutJhULMgc0x
ZjfEKQsyVqEjGwrF4Zh37Hvh/ddjOow09xhvLljWEgiqn9FCzi+TcXsqb0XvQ2yAjz93XjFkK5WT
9g6ZzsjhphfMVeRDeluT4LjJxfMGSMaP9rexzxiBOU7EFrUcDrAqtgicD3T6m2HECkEOwoP85mPe
b+vqq7bsO2ZKIfQAhL5B+nXlxqs+i7Of2WyyMknVCOQUouPPmE2SZ0nMjJQGrmyhoNA87gnPydyQ
UtakG9txfcMviGSUtSKJx6fx+4tU0B1BAbfSDfsgPHv3Qorh/LHpiwpy45VtIC9/QLDKdfHcrOlS
vYlvxG7ZTqxEHnhM2DCqEulEVJQmBwmw8ZNrsvsMowZ7DFdewHACVhzu5CeCnugkbPMi4Or+AsvK
U0DzVsDFRkcX8wiUTs6ZDKSX3ptf5QZ5pKV8sTSvWVpEehhafvEWXILqmkV8ILncygfCBvDclaII
nGlJhWDmnFBFxZ8t3+79ImKfKiyj+SEpHMFWmt2lEWipoJN/p9ATv2WWEDY0bzI+svArPB7hbajo
tiyIDk2D68jAKBcNoWO9y/skcaMvdXmX1DKvGhN2E7/pCICpCrypvQwOGwhNyQvT3cLHVZBeypGW
6l1sH7L87HTjcyVx2Jg/t4eRJbz+zoze7n51LA+vOevbZOw0hSGf4RAMjLER9rMqxuf91XQ1sK9q
bQjxrxxjw1OKCTLolI7xCWvDLwD/CplqNt8HpGsuzwUjLz1VUjcRTpLbmMuFKz41JjEizD+GY5c4
VfKgZxofUIoFyVHf9anKBsI2mB3YUpgL7k3WRRe208WEXZyjHMG9NILrePK13V7U8WOVLgP39+GY
lHrTRYzikSon2R9Et3NxeV4HY9NNgArKzOFGSKfxgKvoJbi/mC5uKKw7/67LdfG8GEQaapo85PNM
mOtJA2fJofhZiRbNwVTi5DOAuggeXHFYG5TKvJ8+DAv8PQGl+DvpnGE1vBOYot4Y1YpGHUB1BwTO
/TyhKDJ75eybVXEe49pC3FgrttAsxYPEQGJtxelaQrbIB7U5K0fUiWrJYwOKvatOTizDXh8qZeK9
uWDjkHSVJlCWiucc2/XLG9nvBUVXIGYvxAbvDgFiSjg7n7ZYT4sH2pQfV/PISM+CqqvCip0/LFPI
fxhRZGyt7PxWwpQTBBgOdCYmZzuyNb9H19ZzQ/F/RogCj9yEYBI1EdOX65OkaAy7MxtlgtJwjaZT
UUUVebOh/HUNtugnSgSecx+EXv+bBQ1RbFlh7tqIH9jlwF3kryxVaIKHpc8P7AWiJu979Rs+Ocfs
dQwA8rd/ywKw3lurbYnTzUChuFT0ipsUBFuhv9hG4H35kYb6IFWciezV+98HTWikEVkvXuK7hCvS
NbLTMNkhsKfp9rXdn/wN7CJwVct2kdewsZVGpn0hWYWLkaXACTbQudebMfnKuC7/GUupfpnyKwOI
ju3LlW6cFgBCAXaRdDt+lzV+EChSkdu3OR3OgGzwSi35e+cO4baKYY/xj1zI2gzd7RAJktLEDpiI
pDZSC9XCF59Kh5q93M3nCuWUm0dBObJU/2zO7OBJoi3iNUQ7sLJR81bu7yXWIhUam1GmX1VtcNTf
i1I0j0EYE/tj0sHptdo5UFm3qoYJLjKvHZnfYi+6oZ7WWOPZbjjNA67ynhww6GnA65YG+Y1SUhpB
KywlpYo7z+dm8xGOZw8pZwwVa0TMIrUmfsyV9VWYHAyuJZL6/CdxtFGgkywt5VBUE7XGN4WIvUaU
o8VhkfY9+uqXlejWxNiP09dz8+mI/I1dCeLE8XaFrhnZ7ArTS370Q+HpKrhxDjj4ERIW18nxB53z
thDSHwJccUuPSezhofLSyvS8y1NfnXoyq4+cllVw5WYrnQMEsMFzsX8MSu49nLnrkEM2Nf0nzlO3
bMK3ffDTWZFTrZFTG2DRQZrQuk0n++Ql5WEzTNt3DUgvJfUp73fOd06meQICssuUSg1Z9KXxuPQ1
5dpo5vDHH9yFP8k1CEruhi0jFLeH4fLUwltQXNdEnWyLCLyeQCNaKwdHQrcX1D/QQhLGZIkp/LzB
QwlUWoW5ztmin7lul7o/lR++We5S2SszJ0i25qLMI2oxv1sIIa/yHyAxnN+Pqa6VOW14QU02ELnI
X2PjvrLnD1qu107oRisrGbdtZByyiD1YcsDttsC2qd6dRySuIkdUuT1DY6x9ZDnPg9AcbZSw5z+N
CHpIwm1YbxGlIxTgL49Mywb/qAOmPX8pICjYiqmQWVdFGjgi7dWrw4rKWsVu+eTJIyMzsyVujUN3
udHEooU86dgxcJI1A+lwrv8ATJJ3L/7BvJO7XsZwmLU9IOEnA+XdViwsUXLkmumtNE83Ee1ugO6v
RJhzsoMqlYQFz2//VEL9U+OdYaijs/8ZDNCxgAKnlRDN9lG+F0pGAhR9ejRjBTJNm0dJ8X1X6Hdj
HDzCqK5OG9r+R2LWzkiGCU12+ueu3ruFvN1bWcoGzcu1XJCePtx+MTl8zKvgBN24hey7UFX3OpP3
YwacgT4WqXMgxgZYLhB62m80iZPFs/FA5cBzrt+BJuAIS6CAmR7jb939aZ74lr/rC7zPh4RC2ukV
VmIXgahoi+aPaqVE6hCGpYW0/1+5X9Bpwwl6tnehl1r8hDBYYb1UKGRD4OHMx8p4bEUUeGpQ13eO
pYlWvHKSMC3ROV6YIoipGbd41HNHaQJJ/zxOvOYVlI2+K3DbSHXRHFWrIA1J3VGQeJeSFIzdnwnZ
errOuxtfqKkS6Uq03cAInhclEAHk/egQVWTPmFoOQwu8ScKr8bRBBeGLWb0OAA7lhfSCfMnPiRo+
Qq84gYoRwwqUiRlKhjic1WikCO9/A1tTfpfjvlFqHHwg7/5QzSXn8MOfF50s13yhzIIVzX5yWlKq
OsagWlkF5/FDqN3p5XxZdkwedMx08UIEBF3Q1pwFP0XBlBTfQNkjuXudW5XkVr5Ci3F7hKnA2vkR
OVuYlzEy1OOuoaNHiJRzYnnE2ryqRggRQoGchAmAn3hvh2zTxmfN0eJlB+YKw8HHsMPyKIulAcEm
mv4dkjgTiCH+90cOT9M/73W5ce+ttYmFFgfVEYNnqhxemXZLMnAZNo0FQLQwb9Ey6S4zMjkTSzzk
DtEsO0Ppiphh2Yntu+dwv9jjwdmdXwv3wCkHXFq4EE74tw5SNlHfD7oVxQ3PeobnE8d3u7RWj4Yh
oCFGAbTvsG7DSLg/JV6QxIsB87IR+NpmWDY6t/OxUreGMqSp1R/LdEJqpazWt4O/PQh2La+NAdMa
qqg4x1z3GT8A6dqTi2g9IEuxaQihPSMM3kkHYj0zb1PPz69D8zsdzg3BZzoBivsBZb75AyfTy1y2
WrbklKSC9x49+YcPXetM3Dl3n19HMzcJ3KM0RCIeqLLXkyqfUv0RYBtk1iasNq1oHLmOCJ/ZQHcn
f4FZkaKo7qJGl8391B7AHiUn8Ah0xOcq00Ho7V931Lfeti4SQ/N2IhEpt8yEJQs7p3A4cvCuuiYj
m4YGBd+WSjRtr2oQPe1crIqepqmMU+CzQNaCC0Z7wBVh6drXRn+AuDMCiAzZdbgQ/jJ93nbA3U2C
OSknpwzI1r5ygEgg73moDjwjHy+WN26MzHLMCSCQFj0j4baOXnblcvsOXXeHiteodif0ycUlwLVN
BnZZZz6KyQsGKbkRM4eDCEv7nBpLV8w4lJCBBx24r9AUOAUjr/4riLQcKs6LppWAyZnDTlv32UIL
M33VETegSpVjliTEpD5eOZVuXlhw9xXT7qg5xzYHJ4y9FRVPciz9JrbgZdP7d4fvSbYucyCCXU7y
3xWOYKS1fM6PS0TtJhzY4VRNI8iNzNpEevhw7t3Vd+jY8Ey8mDVOg9LjveSHSSU/NEx2QyBT/Nt9
G0xXVDlRIE1xuSHYl2VBFSg1WvrrvOc6oNlmOqdpR7vs4BSYAeODbiBRkfRmIRD4rmDb/RWNAAzV
oxG3cjsrnfqwr8ylswX3EWG2FBNVJNdMTGFxzIKf2LzjjZPlvsIOD5oOXpeVKrPFRYgtj1bimdux
Url6Qg6wE8QWV8HU3BQxZb54TSVRfuneyuwOKuEM1MdQm/dvW8TJ4FgOxg+d+hacNWXx1kA8ot23
7Wu0h0hkbO4G5ROZhFZiWyHSN9Zal64Ay4x6vqNWH0FSsp9GfmxZ2sPvHalEUzLZDb3ib1U/uLSt
V55NVq63Smj4S3T4CFbBxjnbxgHXc2gbAMJX2Fov3ArZeg5Q8vLWXthXgC4GMmAEZNdApJUw14r1
baKX4tCp5cp1gx/KLh9QcCuquotHBpMFtE3Lyrr/QQLy9biltXT2877eQRlOAwji9nz2757K+jnt
CDkPKJ20nekHc06YpSlFpsi3OWMHRhm9iFiMwHHF4tw1GIOTl3E3nDRvXJ6B+g+DzbCsmfSybyL9
1R/4DUwRheAzk7BcyjnjqPya55uTq9FykZbx/7UlLx0qWjguCNGpS4tyza7efeT6536B4vaBr0/S
DXOFwsc1GPCb0Se8WsE3ZytgxyZ9Sls5AqhHmt+GyQpePBq08OvH5owZzfqHzJSJXIYXmrUkDmnS
ybU72X/g+Um1nlEg9ttgL/H1op0pECWX4z6nJRG97nNLsv/RRGxecN+UdajW9bZjUr7oWdL6WAHC
jM4sQiLgZB+9ktoqB5Tku5EJQZxRp5xMvJbhaXM+Ox3dLUrS1HDb+/cKLjUQuhUiGKOOnrzXE+if
azdo5P3Pv1RjU8igJAq6hDoY2YgDN+FLyVJEfVDIYN4YfrVg7ebHnBmJsMP+hY8l8yyiTYU5Ej/t
SlZ05JJpkfX6Khe7g8tFfOjKEef2ElOLcFHUreM9+QROippQG73sNV7bipmQSr/AQAIc1GxJlVFr
x55Y2XFWlOcW7jihhffTSkLLY3ps3BSWq75nCOYUcVoqO2QKPQe2cAPHIH821ruzqKyvUvqovv7a
K8zeGXwNUjAwAmjefsfxJ/QAlXN7Ncc+yv1U+h1lVZ3FojVsgI6I8NHoGhVDbed21B/QNvjO6w+J
yt7B8OHhu7QiGIZDX+SUVIKILqUWBCgtlpIfsrADSJ0Xw7OMf7iJn2bshigjsv6jIBCWVk5t/zYd
Ex63xAxNUqW5t/C0AD8L4aYI3Y8fqeASoPhv98DuP0jNT464WmjQCFZxWZBFnGN1Slsu/BuY6E+x
LaRCSUH9Oqp9KfSeLzuz9pu26SVdmSmBzbuW6rkj92K5kqXzuXZ7CUV3DWojSgrn/9Q0yl4TRPX7
CLclVpqD1iwVwEHjlAS1LDlYniLnegCGncyNYqpHvIMSNxQlK0oWEddbgCrUtL8VQeEMhf7U6Vyp
+wVZr2GY5HV2/OeqiODwB0iFdpH+rsvJ+ATXAWfQ0nuepneqTvtDz8UVBURr6ld6b87Bz8MRFA8I
OvVvoB7G5KU1rH1RQukfLHYfqInP0DD3zBJreVqvNntPCycONFDOYsg14JC/uwKddg7nFklgOpWJ
BR6hA/UzO8+vlo26vWFhQY6hpgBALHGaKA25T9dHbQvIZJD/mfSzc9fhdsnR6ij+0hAvCnXu0emM
BoFjDif+DIAN4IrO0X9nnR87OScH6TAkDd5kBtk/HeRITa+V2IRWUslr0FDJEpQzGfZGEiMjYhOO
1cdIhsu7B9o9FyNQESyE7afCVKglo2bcVh+/L893u1s2CMEayGLptARhbZB0CbWYfv/qNtcWBTAC
aGF9++m7EDX8ZGTnDyx+pNmsIq/uFVW3zHqkDN+NRXieTzBcg3hMVyiBpqMTIImkCRWvokCezdp3
OFS4pyIhqhw5ZhLthGy+Rzlkqcve167Dox2rBcbrT1hL5+CrsNPk3Tht5SXtVwTrfe/zS4zn54hA
VIN1FKxo6h1W1ir8sLBwpIZto6MaPT0uX3wIXhn0vUnkcBDt32M8ejBKDgofOGTykLmBV7kNCP8L
Ed8CeN4+muDAOKbaqfLk0WgS1hNpKRC/ynTu0zAj29HM1OnOONYCC8E5o96x/3H2c3gyQFPcau1x
/Qfh1Mg2pbuOedrIeHjENbw+IY/O7ZHlqe/N/FSWoI7S7nRQCuW4/Q38Cnq6ePyhx2mHRpd3BkVf
GpMXlS9mQq6EfplRk9AFZ+I5hF70oqPW+n5dszEhzccqaElXH+ggS/nxOzq6MZSnRFl6UyqvAxW4
gawQpIs7MZNsVv0UiKx8emAYM4EiL4Up4Mr6RjMV1/M71nzgDi+wEnkKUh0lhpbOsgwiGkaRVp/+
4mWuyCStz5ikVzlqXAOKgVxE3nNrD4j/pn8f9NJJS7nndmvQvUQiZ8xcDNWUREBsMr5nS4lX+PFN
QuF6S6C5sTyDYIkNOt7QEchVX1lg8lXwjwetK+4YrH+TucYNmvEg/+CVs1vyk/nJVursPNE0gvvq
zCC69D9ZCs88R8OJG4+br3wFRwU6pmgsv9KbEykFI+bQgiokyWIrDjVidswZ52KAm+qSClBBBFKl
E70YVbSgMx4BOM4BdwdomH304MnhS8SZynKpFYDyJyd8800MJfN/rq82NqGFyIqj2MPwzGXPPYQn
xIkgqBEloaL2VCn+fMXly20HprzcUb9ZGOOCOq3GMdx+T/QRCnLRs7Lul1MPG+/Vs5qWzbkuqzIF
w9r+nfqGOrjxV6clDhIFoKiuCPrF9/8aV2mgUT0/Dt+fn9fYhn4DsNVb3F91C5JVd0WMVLxPTza3
2mZL10CiJG0H88Q3EAXfGjcn1bxINMBi8hVFFxBmylOthDkC7Ku1smM4YllY8+SXDTx1s2+HB/gW
ddyX8NZjTpEHZApkdGqCKVWVgk6zV9j45xff6qf9yMw9IIOpBjeV909vrTWzheTGnjPd/4fhskoK
mIBHl5w4LZDTlGejCTMG5axwpit5v6BX+OfL9tuhEXfNy4sj1Hv/E7zF9nI8dVnlztMszGX0ZxBE
tLpD9cToe7FxvQUllVq7IwFEAz/ogdTidMn4Ysw/UenrWYp75GV7lbsL/9xZmfWxuUxjtsXiWjF7
iEZpwZzAL3JfjM47ECBTBjhHK8+UZkj0yZ4eH6byDEPQSNLKBvJJU8a5b+bfkjGYdRpDrZ2k62H+
gluyb8pcEnM1b6Z3gKTjASlCnfptKNoXUHiIAEUz4NZx0Ozfm7/EE9Q1gURZKE9UdkOOM8NXRyU3
Jq1pMMnBUTxnQQlSbICUUVh3Z7LHyrAbKysyDYPKLICzhNK0L7dH22cm4T0o8EM7swcvh4LU8TMy
lCximJRQe+NGMYGMb04tRrfMZFExORhr26tR8ccW40ipQ312So6/Hd701NPQwvSFPg+05lEWbfMe
oy1Z4a5JOloA6z20T/B3wBcRHGvz7EhAhy0TwPKYHfK8chrEaG1PScDblwfoHy76JqfERpJ+toes
YHR+Ur0/fsRD1cUV9HpfUQd5EFZORGgfNp2qk235SjDIxqogCbQI783f1G45X6Q97Iau/JfLQmSr
wcyJ6n3+umKVv9IPGAC4UzY9jC5vjU5ZtCNWBugeEg74cBgXkD3jYYAM7z1j0Kr62sWr8tjSQgMi
KC0WLdlgdigWTA9SqL6ofoLsS0c9V+wkHs/q9uOS9HZY79ALTujzeiPI4oJw4gqfSJp9RaQgCXim
4Ws0XE+E4AGPJaeAcuK2fIGjqq9rC1E5j7PV54F59W5K5Pded6R4ktVe0yie0yL3PG+0fkE0wgD9
/8bgQ0gy80TV9Svqrjz76l3xksYQk945FOYiOzkPZUOjIdVCYkHNBezNjFauCrQ9H/6leMX3XrXl
nV9u09BK6Shq29Z3cLt9km9Sy4p/9aOPgqOfCmowNNBZpKFGqZSuPxlRO1uQCYmjVFjYEwEZ7/X7
wU7quUWgEwzUb1tIrGPz20/rdATH4CTSEtIzWv2Vm96rKRE3PfBW3TezqoeO8sBql1VK7elhqVxV
fI3RaVVyEtSM9NmPUM6f/GQq6WvVS8vN1G55SvrWVr/MbS8M+GV07QXIEly7M8+MgH80eq12/Fhu
9Bh79PBrh1L9G8ErJ/fMPae3x6otzWV3wcypu4WBrhVN4skbIoTs+joKY9AOC5bVRc+paPd0T8D5
d1TfpkwthludjCYcR/s4+5b5dlp7qz7CYc9dMhOTZQxw9wqI+pN7iYE/+MO/RJ0pu6xLVLmIOwdc
yiJ0JeE4+76HULTW7cPfGRLmcW8UqapBowbxHo1p8lt8rcmpTDnn9gyRg/bLmnq0hcY1RKVIXC9v
AEIXzR3cuTgOQ6asyzBvZ7t/kRPjgP1cdDFRtOx0U7BtojDApbyf0hW8hLN4hicDhsD99be6ahEm
QThN2+BGYV7D2AMa2jxds04vd0YQjtHOB+6pZyBhUHyLlHIqQk20DzrfeRX0/J3cgSIoWVC2pcyy
645gM3nBgaUAXzQwwvODlZquTfGZ+gmLwxI7CQLX2DyFu6tDrqSCMaQpAySvsvUxvQR6iBEEHLzo
j95nX4yY7zKMZuGcUMtJNFN7W0z3xLnomvUiawNrh+oTcwQlVWv8y20iWiPs4QFj/1W1glsvKkED
zwIMpIGRa9rWJw6Es/9eDLcNnC5rX/0mc1w6Qh2DxDn10a6kkcrb0KxdzO4hf8N7wfC8Uw1pQ8Ja
NS+vJPJCBTVxNoNMwLDmqGRYVi2vwNApBOX3zeUHUnU1vTFrNNeQbXf/4qZ3Ze18dQfe7E0Duwe2
z+Bm6uxF9FRc5HTJ767c5Nq469iUJa1LKVbUUyAzsD4qQmTqXv5bs0VwI0792QEbtXJGJ5yZb4DZ
lb6vWPjSYweR5pNXzslzo9xpoIfWK8d1P8s2f4SHMpKl1nG0M/TLzHwPJMCUntlQ7Kxp+nrJbg1+
za5O3cFCRyZgWRxFz6aeQJ4mYPDCfyFuwPhTchdTNzeYCDXezjufWERWRPiNrj3B4qyhM1Yhd1Uy
PdDKKStG58Sxser9WH8tjONG/Outx5+ta1oHcWxXwrB9cXE8YwwjTaj9CH8MENRXT9EnLpnjfeW7
QMsDAMD9XjhoBjJKJWEPTtXOqcoA3T4uEe6lpm6eQIBeTWNMjVfxCvsEcnddEWl1gvtp+erwcMYF
nnR816iwJ75evvdPcIJ/V4mSuAUpk97/uABnJ7N9zz3+w6U8Dfd7Iy9yaLNy3hvmS2vNcJs+CThg
+szqC+5Uea3vOS5x1T8euAa5m/QiDr5Sq1aAmlf8FeF7LocZgy+YP1R1x0YHQ8P2BSez9iMS7JjF
YAoDkDoi87Ma2o9PWY2femYN55wnxzut6kQANlQsCZR4CbsJQ7rWwI25bKDABfFo6SXM7iDH2VtW
m3QWznOlOvjfjjp2pAsLogaIReEJwS+9yO5SRNCYJlGZ+iRlkFtoZHMyJar5GNDM53rXEo/0niD2
JcYc2ZOh0WB4QGaQrkGgHzRI6cm5rJ598GxpJ/fcijGMuqXnJOp5U1+7E+Q8fcGlewxQ9MYwDXoo
hCZLDT6kkyGYAl8Ta7j+9jkvbW2Xi1gQKvEG6gTxBasCeNjle7U7bXCEfRvaCEDYeMZKrexUsAOi
sKoEf+ebOxE9XWdk2cD1EIN4MoJZ1HYRkvg+52yvl/3WOZJiBTG1UPXdLtXYfhJM1o2jsbWGlyDG
u370j34uofbARTjJS1sEqmCVVnE+it3dxxhF98lt2FqUTOBoKrlOIU6Zg5BJaE/M7QfFViSAOVsq
xKYVXoYh4Lw0B9nyd21ZJRG8DSRyPgQVrcWmt6P4+Ax/kUM0m5cUprL97x5R8sbyY64+s/57rKWV
0hNF8fY53TmYy18JQL9B09LImTwasNJTXaFT9yrQsjH3xA0HsSDwN7uBgbGYg+0YBIL8Uc9ckPPO
n9wclvwijh+X5hhw1Q01zb8F7n1jp7ZJrByktlplnAvW1IWKJepV1beRYPSBu3yNclBViYzWwyIN
km29uzp9hkJX9iqxkwCYk7McUmMcAu9cdrUAlGQwQr6+MAfBha81Olb1FrHlzkBbuTJbmuKI2gg3
0tA4WyQZ6oyO3fhDoXrv9zr3zu0sV07o/k538JnDM2cjxyNKLoV9hW/m/KKUCpN+FtNZD7kOFPcv
8CeCe9hjW9KowFDq+Yr1qDhHP06nUn6tB8J66tB4DKcm+A+wZksoIJTH0LH7eavSdDS96W28VbEU
TkhZjB0GGqLr7jiep+bPFweVUruMsUA/A4HwWXNtbngHfV/+QvQ0GoZPcnJFnzOPi+/3TtmeO5BV
RK2AdMHzEBqql6UJTO4qffWd//vRy70zLwr+pR64Q7XHBJXWesodV3tD0roUCN1UYKW7w5Ph9WXu
sOG5D6AUuhCyRNsfI0v+y9wfZUdXAtERa0J7fYfzbTc9nVezc+1K9whWVrVWFFVzgLxpdsKsxbGe
6nBmswvEF1BW6TOFqM8+1OExQeHi0Og1osNUDJAbRRqQQH4DryHa74wLJGz6mPm+SgUkDbllJbTa
Y15R9x78M9O3gZAjZvkn9aEQ4TNtX+YAOfqkHjN3C1e2ES1rBRmcWtkx+WHeIqbeSZOsr5rUWPeY
eOHs8ka+NZ2Xz0yfGkCdtgkUxpYZan1KD0tcW9IZCTuiurHd3F6pr4QNYNTmXUU74kbWc2oNf0wI
HPeqatHm4caXRymZ+GL7BK9n+Dt8sknwaxs/CU47o+1rXtLGQFJy8J9eEYNER4es81fN5qk9c9kT
wzv/imRpZ8+Zaa1haA6VJwIqLihmTvHZKSXo64ypCn7CHeK2LRiPbMRIMmF+HcqLjPd4j8bhgzcU
wWfC7ud/AFYW3EUqa3x24X04ChTgvCWax1SKuSe12OLvN6BzMjo0g/0mwAht/KlKlB3FyrbBd/s8
ydbAtG8a6UTrU1Lg+Hug8pErADOQ/D3AEUYpKRcC7KwL06mTzkbqRKq4tYfl2rQRmIrZbdxFfN6q
Ttk3rQNsD9S6r1YQoc+2hVvGMMq8ZfUSSHrUVqYq2dTOg+vdQn7qXshNZGVHLKl57WQ8Vs+Cj3tq
KiozAhwTWMu52fTYx1V5uZDMR6rXWiOPK7aJPjePRFl4qnLB2M8I7CJriy898BOhz5gS9Htsnq7z
XFB08Be57flgbgDuWqUlsDQGw22a3p6RJR72yT6nzvMxbAZMhM/qxNk+wP7JSmsMvSjg3jBkctj8
gJrHh0qVRDybNh94H4WrBlDF9FXOP/Mw3QCcbeN0QDSfOpbqUHbftcdksuKD6UgHbfzEPF5m+AMZ
Jr2Boafm2mKN5onKnDetD8uMCwot/kWrtHByaj4J5Tb/vJzQeK3EQgCtPHAO+aWe7ImG9/hjZaSS
TVLNXivAA867vtgoc+JGE3G8tBuA9ttQcbXGdX0ncJT9i2w1EPMgDaQtix/QpjCYTAQvArZWlXK/
n9q1mcOnfkHeA7lZEfDqSk6DR390usjPTJjA99uPfgxSOKT4P2oSzGBI9vAVHWXvEou5bH/aMgcC
I7GOWsWYyRlZwGchAht5JcFdw2EJTpDuR7RXNwRe3WNmLYe/r6Ra588PYo5sqg+zkv7KlV2pYX+G
+xSzO6bfOI4Md+b5UzsKthBezv7KhRrRdGkV/rbVXntJIvrXDW2ss3sAO3ZjPfmV1FYBh4vl4sOp
6DvpcJ1LMEAF93GIMxXobUTR6K5TbuO+y2H35LpWbAPiRqViMs3twgeHbFegI1RmKbNua6cmMRGw
BwgmAF+uJHr8f44CV25jeP1vi2zHW5/XkGhe5HC0AuAFY2vlZpXT+Uc1mqjq/K28/JkqILvgqh/p
9o2fpxT4j1ONVZsdHV+BDHOghQvg4neDTDr+iQNl9LjgwZlz6v+hATWF1VERmXvxXlHRnQpEeMnQ
v+AE3mZhRMCSMmS9Fe98F8ZtZuQLVLzaHJHp1bB61XpyTLP0NzvUkM1LnTBwO23SUP7JeWaq7Yy5
Pn9qF4Ft/MAjOeS2udt+BrhHhCB2La9DwUHPxYMZX0PKbvcZEMyh1mQ6CAs5gpQWf4LED+pBSxV8
zK9Fqj1hxqP5zZJMIVC3BNcwaqvDnLp0b5XUSTf3ry+T0M0M6u4+JZD0DHzMifW3CFB11wksVsj3
GVWM0t7HmF9Uxze2WqQvEtx6XwxRtjWnjLslm4MEzZJ9I4SHs2FVh6tW4Rim2j9j4uFyI5OjTw5x
q35HNGumxguiJrPo8V0PB7TutJ/lENt4VTJVGgp0aUEDCJKjcFZpsr7EE9f6eec2jhf6VWIimhUR
aGgqh35wZ1RGSt7vLTZI3BdJKMp7+qHLrJHpxYaRVM2DydB6vI2nVu78S4LyXsMCRIqlVAbg3klN
nUcLYb0gBpft2WWOmBbATNy4NAr8ZQQ4s5a214Shf0FhveS7nYCYjKPgjT69JZTyxZzwjSw8WoMF
RgeMnCi1+VqnuVKhOrw871rlfbhq9KwnXdwHsIhOEjJ1mH6fNyyrTGv7lTFRqw0V5HOrmnKpYDU2
WUxcC8c2QaxoNYY7PjgQrmoOr3LKO2fujDVaOblRjxMUJiVDecPFcn/17SnLEsxu8Bvkqu5KdGJl
6RiLhZr7hJfXMcaV2IE7ygHFmq7jiZYz/++/c1ZccwSb9IU7MGrIvj652VOkZtB8DUXpdQbHbKFr
RoMvc1Ky23SOm1POFu6No4J8ZnkwtcM3QPO3GEl54RtgCc6h1QIPWMu4Upf80B7fHMaY7ASjUASm
T8/qp4iLpzoXNu/vKHzOGOAl2C1A7Vl17TB2G8VmXee5jm/s1YpGhqk95TB454RvhshV5RrENcfP
1Y4VhFbzvxNiDePB8Vrtbokc1JNdaQYKVoFf2e8NIwzwc2TOBWTwLnYeJGBpagR5gX59CmVBodPn
plvg5keYrpFgqevW6SMXirDwwCbomnTsrDUVCmCKgStEcaS1TcSajwb21TfIRaKssk5YBjo23PHN
dolGEBxXshUQIs50xok7TB+x1izZbCd/j4/Xtzg2ICocULZ45s9huzSiOSV6za7sljXsDdpMKmax
n4q/DSS8uLdnEVRw28g0t8p+gKf+McL2PC8+MXS09yLSYL/mW04BiPdB8keGlMWGwoDm0AK61Ocs
rHn8w13k+6kxBVgF8JXRi3IiLc6lVAM4VD0ITUTGfvRLwdp5VATxOMxJeUc6d/kcZqWPjDP+AfF3
WGqc/d1kTc3WQkQ3U+ZsR+1tYxXlKbJFTiOhsE/gATxfBfi/Cypaf17gl9Bi/c+619spu4cQO7DE
yP6V3CgWS5Cr+ghtOdwA1imoxXeqPsCDzxUgXWxjwXSulYFrqqMkTfbdsMw/Gqklsnfn70zN9o9R
Ib/DacYWTKvFx8yHqX0IXe0JmZi3zC3PtMFzYVXTFPapwGANmJ08y36Bm4svtumIoMU+Z1qwvwLa
2c0RM7NdKjuOG2a0Sv/a2bjO3TgVerVKk/IhA/XtCSTN8l0ifZrXB3bDR4kQOG7VTJJusPPWC0vr
7N6gXFuQAWWUekfNCjvP+9Xy8g/AsjgZJQg3MCxKTVltZgqBYruxGcTx2MlvhNlLIDIwYHScbN7i
jJV4OUZmHHof39ezBUG7VBuCCjvQV+RQ7sg0k6kobc5KHOlJIpAGA8c4YvdgCgOsU7QHV38oWTZi
fSNmiaaizT56H7LnaeIq0GD8X/kciYd0a83eHiDqrWmcHxzTffnREikrKMScHe4HrKluFFFBAAb0
69krYyjD6GvGZSIBtwL7Lqxe59mXJWgaM3/ZCCa3KwY6jXOY/HLzbuG7xEHO0Je0cw9TJEU9xLU+
7MWbVUnT+frI31DDcEFIZdoQgVHSChNBFSaoxqOimqls7mHTIQdyh+eTcPuY/3A8kI8yfgzxIjuL
W7JEg+9OsSdU4bv9prE1vFhtU8OxsdHAjv2q2W5Oj2u1hVub62k3nhW9d4rMOQbHCbo3N0OeTXFC
GrKyXSDl+mVa/RXmL7VYm9KrlZWAQIvXTggPIpfChLJ85EQdCcCncQW8UV2VLP6dgosxg9t9b4BW
TqAyOhWktGMTHi3FFAFYaAeu1V81vw10GelAO9c5qP/Efpiwa/D1IOiwgFsm4+ibEf9YcpDxOn7P
9sfFzlwiWiHxfw9g3t+zjs6B0KH+sBRtAKHFTLPVOJmbd4Y4rqaMDXzA1LOenuMbKFhGCUrmxlzs
Eu5mhh4xqPkmYH7jNllB6N36LFCdGblxCAi1vRNBEaILIm2f8/1N0SvaNVt6vGXQQ2W2dLw5of8n
awydsN4jz0wU3AGmJGqHY+r0AnN3cCBC0s2UqeS8bUaWOnBBvc/1ERpLtKNUAF1hXzoPjQ/RIovl
GTODOF3LEV0pUQ/DB4oG6rAYagle5pGFWPbgeHC0SExlt1u20fLcwUL1byjNNrgVpP5C9oRrCTHo
DYTVzlO4I8NhFb4QfgauO3zrhbHqblp+U+4rWA2As6+jbXq+DnBF8X2N2Ljz2PQ4aAIRAgog5sMy
21gjcu+KHiKB1CcjBAzqn+dktc45pdyogJQk7cv4icDDbQeoFybKS5d3rgC28WtMIStOe3oDi0HI
UhI0/zX6SEBEbEWz1llXXjt0vNMCmzYV/v8WeRAKWylGb/AZ0G1Xlww9JRjdleCfpIMOZCR7uZfS
FwUL7SudSNfR1D8MrV4MWzjArZr7eGxY/JryrzZT9LBi8/KiQLyUcwecx9yCI1daKKKio7BehhiH
chBIq2Namt/uf3Ck1u8iu2+RVj5eK8sML6NYb3Lr47nWAUCsUkncfBPQHv+AmFUIg9A3+lO08tmI
m+IfOYVym7CDBOsrDfLra4dzcC2MiA2IjpTr7P83TTlarVQzvI/PtzTrKFWw6aCy/jBd9VBKBmcC
3wbRh+ATCNBDGr1NSQ7PEUg9IUgevjOi6mgoxGRWkR7VcY/uT4qbNC414vJdTYrV9DdMIqAvk12b
orKSmly3e7Einw8YOoc9DmTj6Xq4U8oMqnpgfL7W5hO7/vFPeCXr5Op2R+QaigFxWcXy3taBgIZ+
A83Cp6pPq+iYuFJD6Pl7g+kOSla/mb/5dmrohQxzxq1isgMpo9HscTbBRPjdqju1pi9WRWVDqbFn
FYXxhtDFaQ1hU4XoGKNfb4Yrh84njS4Wc3qIdmtyca3OLnyQpZ3PYmDNzLragkshRb/FKVwuOXra
XdNmEM4pMSYizVYaG8pfPapJsYveN/0LEVBqC21bEVwb+umD34p5qIHUGNb2usVMq5Y65dD3SXlp
NLyaGIfjT628RVz1CdQLRaSasqLJ0njhjUQhDiXR4YFtJeAfO6qf2uBrxPsM1nPed1XryLSHZuao
g3xADml6kkR4TV7nyY46RFHL4a2jkjPh0Ivi5V5dL8tqTYrLZJ08+Bb1FL9IUfx4PFx0K/5zdFr/
gPbrW+rwc1aw+GVPew2ScRZvpc1MEnQEi3gjbBJ8D9qTgztfrZl3xL0FAQQqN3cBJ6sA3epm3mNp
eB8yjR8mbUR8yYhn+mm63IzaNZuJlilNZOjL4p4FZhkxxhLVzG9zclQMEiwU16F+8QcXpqCU9Cm4
s7v1otsAEkt8WdtzNDWGc2aRA6RTJ80J0mvBz2xV1dnXAN4mSNB4T1IcYCUxAm9g0PuSLdP6esjY
sERHmfLYboBQt5oxbdfr0/e0/AgD1lGOPYJ3VtnMbM15GeIxqB41PCUhI2a2OJVPyWFLV8R0haG+
EWLEtC3fwTdeqieNGxLH0B6UViu7RcM6+WRUGEW0rWV7h5tR8j7QkLA26z3LkYaB3xucUiA7cSN8
EFbn1MN71SJ+CfJQ/NlQIewzbWyFOCeO+8YYJawYZm5alo3jFFV9TqgvtkvRYahw44MsyLf7EcAw
yrFtdzLYSAPGqaMKkdZTH4qRdo2i/7fYUXCmGf+XYUf3JHvyxKYHk/hWltGrS/dmYViyvYG0n1lv
f33iDLgHV1xns+7YrjUMZy4TDC1OphHp4SdbAaRfTAzs5zxL54UEGXx4eLj1qO8uQ4r7AFR7BgSC
4tcm86KHxpg0q6u8YqUGXWuE19335d1Cajtxo6H/KKlzwPJcyfBW3WOo/UPzBrposhzKnlMHqvNf
XoEfja/vVHrlQtK1ppvOrluuBf/Es6Ysj6ymF96skkC5vuAft9JulBCNgOhS3ApViqHZfuGCel2z
i8yu1Ig93ziRAqHDnJFB1BP25ZFojYJKk9Gu2qYTPzINcpuNCQgw02OblDA028GGKNaeg974i9B3
iJf9CMapnu4VlK+l4vm8a7pRXz7UQK0HwpyFj7zoH+Kt3h8og9hgEmJjyjHtkG49YQ6D2vRBD2q5
H4qwwvbkT9jC9UoHHA+9t1E9XOj0ioFRSPw9UCWC1GR9yBLb6SbZyMs6mMbrnyj1/iR1qYt3aFmZ
7NdTgGH9TDlaqfvue5rlGd9m7mEffH3JkUbmqh3RbYrLfhEkJX3qXHW7+/ex/PXsZG2VCTIk761F
RAZZykCEyRipStnzgzXFNynZIwYRjW7gyvEe7qy4e8XiEPsghd78MG7rOVivTBswGf/CSrn3Fqnn
rga1j5V1cgVG88sr+ui+j5PdjLlDMsQTU88ilKZHaxjoPVgUg+BT4VfXAdQ4pqs+KZUuD8AwpBL9
321tK+CyaFF+oe7qhtuIWUmqdzDP/ReoY4k6yFVEzRU77FfUJEPPg2VfbR2BAapvkedvy2B11ep9
slvk0QcHvsKORc8IhqdrS7gJMO8gOdB7Dm+WetUcT/hKohL1HwCd9MDMXndR4+j6aVZBcBLPOguB
r9GDskglThBM4+05lEft+0AM4Jv389wVsoZwjWa2RZST5zNJU/bDm8sne5ewF+WWbjTFjSCNq/Eg
1KU6RHNcmpavp/bVX2YoKEczePIIvi4SE4mQ4VprhHn7emv5fqsJ6VUwnR82YtQlioDYzDWxlGWG
5ivUBf+EYpM5sIOUFgdU8u60rMMmwH8EzmwLHnyQLntfjMV8hOMQBu1In4RmKa7V/CfV1ZCdxnQM
cOa7PKnTozzQEXIGoLrSnigUKugYP1PrWPsaDUidh7OlKKiuNIrDneQQBq5mH1N3iqdQDIrM3qh4
jzyvHs4/sUrpZ4mEt2GzLTExHMVSTaBJjYa93lOW6v/fdvrOR4jIedVjVef+zKyvwSS5HLCiwLZd
pIjr+OEuRmA4cMzOKIX14rv9MGTRbTZlh9V0jy4L9pIoikCjV3pa7hB3CQMoLut+EDyBVOR4TMKY
XqGL/wbxbOQ9BD83FUR2tkHOvwlnYHDgMdgpH4UIKKdG0ujzIVDlWoU4IXj83MLtXJQVx1oXTpYp
vzwZhv4Uvq2EVRzHjSrSLG8Pd7ppITYDRcJKUQPdUYHrnQTVX29ISjcKKj3HFlP5KtG3FYTC3YqG
vw5SZJtvcBtYgHfLRME+T8ZWDxMPGaGQM3PQvmyOZSaAqo5HvF4ain6wKphET3yW9RnI5NoXZK+7
DVoOQs7JAPrtxpRzFeiY0TlcJKl49KOmh56H/H8H9W6MNtvB9qtMxkUcrWpn7Qgx0na0fkR/t8J8
G3GaeWQhl+eSfQx3FS4/hrWgvD5xTrWTX1WdqnkTtL0ytVF4WkiImpeO8njZKYoHH7yM/+sEmpN9
gqxN7EjA+MhQFA5Mgmecro/wh2Ij4RI+j1t4D2wzWCK7/6pYVcM3dqkeOnueRkzf7NDb/qOKOFQj
6G4Cl+rhkCb3Zohm0mZ+a9LMD46+a2tkimdS+pbMzswCYc64Ppt6UtpNFeu7y9uXq4590qdt5PIu
J8KA89Kyh4QmxrM54LC+KXY0TQkdCpjqcbqGBCsZyUgljKk3+MeX7m+z8oFhpFPFNyzR/GFCDy+w
NE00tJHpUytrUV40TC9oXfz04HSFM1w1dD605IG8QXXP3o103C+CFb/bZ0I8OC7A6Dme7Gx3RXKX
mlrfnp8ikPkkBEvCvcejsNKW/d5zZSzx9yB2OFFZYO05/qsKnGdAQJJ0k3YYc5ZqPIO1PT+l+Kn6
6zyNgI3CY9c+HjQxgIifgRFElHP5ZGGmUInfJB/o/6nD08UdokBTEEI23ylYP9L7wE9ONoZVaySe
ycSZfYdlOsRm2sYY3XwyTlq1M8I/qj3oFzKzhxAPdBc8XPoRB7CuXsRuYheaZK/mf/nRzKL2Jp6l
9KwPHSIQY6KyJJXT8zD1F4XTKOB+IbLtAECBbaVA0CdYCIAMhSxFYH1l9MvZF/BQFeuyAKlRj69O
rc9YpcFS6MOB55Gcsb8OCRDbXgnYv2xJmd7GRqS997E9X7zlwFJwRaSOxDWELuFuJewDqkz4u7k+
lqarFN20mGEJhoidum7XMfZ/x6Jl30iPlNBYTDwA7SG/XutZQ5PqhDqS5/h1keAhi7lKWbOkcfM5
ocI66uwV6hLkPgbWjJrFLRRVku+3lIslYnBgisU543R3u3GWXwieAuVtldc8LuPRy66FET85pGuK
UlVEF9mHDI5JtwwjU3j+SVau6SnPhx+O2MoZAFOhLJ4aVvEyOs4bY9l8BoThZdFxuLMErjTSPMmy
DB7CeDkJKsB+xp1m7dUWHrBPH0pbsSnoXhmxNgK/LoF0HfzyHK/vcLLWDdykMicynMdOpjC6zepD
AmOvZXhW73SKl2pWj9tFHF5ngKLJbhhfssvmiL2RZAJAhoyQi6ZJpRnxJhf9JeQVVVh8Hzk5NlH9
h8JtPq1bQZ5xd1+SawiVeucGlLs9WThOsUlXxQ7+WGpBYspniMzcZvEIZrN1BT5nWXnyG5Xl/gwl
ynN5zx08CPB0KwBxGcCxnHxLQmw0OqQhThfJ4hgoljxwOsoTNPIaQ19IwWRHmA73qFsLozTBwuVx
Xf6T4T8LGjpJ/OYQxyDi4XnxdEQnFKiSWkCMzkgAdxLWf9kpTEkC7O732yH9XYFsGBP4AG9gUT/b
V9pCNbSKNRhq1gaGfeW8E+uV3MMJ9QfLMt/xG/yvoIogyqO/dwcLMOHRbansRYGa9izHG0sE5Qay
D/SaIgW9gGFKdfC/moZj9WH41swb7NDX7yTBVkBHgSSVk/da+EmikPTADffGEVyGwI28UpzJq6zd
6otnw7ua6oZrcxLRYFaB9cGfMoy8L6iGFlfBB06Dz2vztNPTmwMdK29BvXyLVKqSA1nK8BaBPxyk
ah0RVqjgbMYudQpUSBSQ2bc6hwQq2ifin8scOLjYIO4bmw1WAU958w26L+Y63HEGO7fVy7EPMmlY
zEnef9SwAFmwvBUanmKKkzCR/epj+s1r/utWpyWccMEUeqRAEV2hGC3fC3ywWZYozaw1cTWyp4Me
RZ24IRM4hz65Yg8e1rA+WpzHV0myPypI9sV7PZBbe2MFCb5uokP1Tx8+q7FI1N0/81tzr47UEiq6
8eIQpbADiou2qk2IM0GNrCf3Qx3xh/KLUrY4iDuB+wB2XE4+JzF4O27Q0YeC+1mEGdivXgYAAEt9
0J4LUx/q4480FsO2g1IgJA2ABB+lW4iOD/GQGQLrWafsuBKWzN+/pgzhIIOwv306PUL76bA1sF0p
WQF90p0OPcBOp4tQCrX+HPau6I5jDOcBRuSzELhzdJVqZzGWIoOznbRO/klTSRx/Y1zCK9d+TpQb
lGrjscyDk+JZAsaCWNHzwALkp5cS9ODNZir6WBXnTIwe+xsdl5zWczGOAu9f1cWE5t2wwi52D4td
rj3qgHVw7cRlhQR1OZ1X0Mb6/yu0hw0Bn95AJCqWZZgdtGLojhgjhmgwZ9eFtXBVFhLd1ozLFU5L
waOL86Bx0ZZVzhJuU4P74EACn6fV5uIPguQLea+itCj3MhEpjy6qkVb1x2ToUYyc2t1hfs3y9Gnk
VYF8av/fKGZ5AaEpLVnp88+v+56anTwy7/aoweoy7S8rCLWONq0q1y44t0rw6sx/SVBB4pzlhnua
qXOJKv2nxXcXyeRX2lBdq3V+L3CA+ySiJ/ZZQFKVCrXMXg0GGjAYvo7zt7EJVaSESl83GWCwM4zC
VYR995a0IQCyDrpafAmOwSUeFp2utWjYO90dAAYd4XaTB6lVYUrBVG4VItaCCn/pUkq99cy8GMt4
R4T18A0Z4STc+FY1McpDjHiJ9iqs6SJFpe4QlGG2VvOi2ZDqOi7NbdmX7oOBHGUU2G51tC7YiFoc
kPxr7HlVsa8UPjT1HOSqw4Cd5BMvUVLluBighzlxnS/d5Q99sloC7z0f+pc000HYmmQoByX4s5eT
6dAsvC9sa7RXv+3TgHF05IhdZ3hNNHg3qfKZwoIo8Ksgg7ffRxyZroTH17Nb5A/lx7xCpg2fjfKF
iWRUjyLKm41mmNFw7ZtTyWYkqCrapWd6l2lFzRkFjFiS5lnXDSdsqKGbh/nYMuRmIru49TRd+nTU
tYN0DoHPXKhEpVU+HDz4oPMSqsWrQNpMq8FPnkjxvpS+UwCrr3tlKvLBUL69ePtvDpo/hPoh6KJ9
jeD23Te3lMQkA50CfyiohCQFTfwMjN9h0mTjRcYyA2fTisTwD2n6+Dwkru+S+sPv1UDyLObQCdjO
OGaXqle0357yE43yV9SfxohmnOyGgXDo2FuA6szIJX/VIkLfWQ9CAVo82AGto1Cb63tUmPAWJ0ww
KKhYmjXL40Sizico6DeyMBjq+pfjElb8V2JFqcazXJJCvd65fK8HFWSszdNpkCP0m0dwGMnW9Jza
xDnejZnqOpHbs3EEE4ik9+elQErH0PixuzBvqBsnYTrDDnD7CIKRQQscIowXdzLKiscDkjbH/f7R
ZbNv4dVM9gJzXz/LYcF9IrgXO0Oio24F8WNOlsa+cPm/ugXm9V12MUUJ15csv3llH/jbhjjOnNkD
whytQlr+SywR/AvcH27+uXGrhENvTdtCE3x7h++73yoI43481QQOF9J3B+ATzY02fGMM9xwipR6k
cWKzrBvCROBArCYHT39eQlvCzJDMuM5h+2x7e7qW2R8oASxPsNWMUbAoKAyV9UjzO+2UQ2X5Zvwx
J/EtY/KiMwTuTpeKbAt3SfeOlosnhjFyrmFXqQ3ja3EkY5jccQdhL+r0ZLs2zQmKgb+fRuPoDFD9
KqNlw/ixNC82UV6uGgvrJjSCgacjpWa2vhkD4GzTtagbZ/ulwt+EOobCNp554zV1Ip9ROynobbdO
uTR0M7Sqtup1t7lbiILFn4Vuh9Y2LEAATN4U6+XoEujMAm9uW6luJk3csu6jdszyqlZ5GWl55+9+
JD2vDWX2Vl6cNA+JDUxsKqUdO4T2wzJQgXuh213eBe51+v037ffQspiAyJrwpgZYsqM2TFl9Ij1L
lNrpvCbCuH+HC49/N6xSDHv8bnzmftKLtCt/IWummhgZoeAMua18pUTQ4HnsaPNSqTmkR0Fm64fx
VuALCWtoZAde23UurqxBTwfdPaPpOIXxzLZe+8KkhN8SpoCzajH7KAi4l2NL/f0zaqWodrWtLDqy
En/d7VxJ7rDMMz2sXDvujlvA6CBKrayV5qf70ILaLLPUVl8pn+jYG7YbR9cq4msWnLsqGm7UULx5
AyQnNK8rk0LKuTYbpL64aXChTvfEx9D1X1r1hVPlFTok1oHOi0DzaIc2KNX18qqC0OrKb/ZVvs66
kkq52Y1TLwiBjHcgOVCHZeH40YYtD7sqX2oLcUePOPRFb6LEI/XR1hcK37u3/tGfDjCYqoUAeapv
9ZV31B7hcfG8vmK3D0+ibjOA8xoJFQ21aZvgE9IvALh8h5xvNIhw0SsPsWJKNpb+Ak9BgnY6ZZMn
4FN6wV6dXrTIkhmsfAopznkj0ErKVOn3HDfi6xiUB3QZq29UMwp8dlpZH0KEDL9OW5yw74E2Cp2I
+VYs7uwOOzokp3BJtRNwL0tV13W9JhF7CyIMfay0ob8TDKL99opztv9WPYR9G9Ju4+orUw4WW1ju
JRu3SpJHazxM9u2R+TR6npCBZT7fjFxfdKn8607xGOg5SGxAmdV5UzCvrwdhLDOJ9Dlv4fC4CtCl
eGmLihVEixOIXJjPMASN3Nnv2JGbDxVmYCJbsMjBI9mo6H+X6HXWxw+3oFNFw5v9RrIn9rglrDYk
fMnaBEXxFaMeKp+jfJvMLzmNAcqY32nG/reaEvHAK2LLAuS+iKIYFPEKu/cq4OGIyx7QhAg7HRcM
JPfZIdufjTuMVloi4J+fBRE48kEIqVRSQG1t3qLX3xxf+3EZ76Yq2Lo3dNyQiLG2vESghcTS1AiC
zrLAradcGx2re3k/XQAcuE5ERW6XnrB/I2hCVSWn1TqA+dElto7cgGm09pLJy93VSlbDMNY1NW1j
DC5dIqlp462ac9SasYp6Kwll/Tw6BTpk5KLUfFGTEzRTkqhfhNRXndKo8LwVoQq3NOz64do7trOY
t66bwqdvj2fF5t8673aBrNmX33tJ61JIu56r9Q1Y6th6ti2hXMubqI9F87T2Pigdvp5RmVTkD03Z
4RGqNNZPFpzB7nEaqIqCC9VJB7RUgUAt1YBwW1/eDp//djgRUNMPmKUufcjMhrwcmYFJc4oNbfAF
VLf8P0i+FMutSiy00REwkmLBDfeYiPqx0IcJ1WsONyHowStN9gjMMssFbfLG6uuDlgmjIx/AI5QQ
c5e6ryzSwK2IlMcbzNe0SnnE6BQSqeUEz01098Cueqy+q9BfwaAxmDLcY8Qgrv0XMbqsiPQOy+1e
Anj+FgUGNJi2eM5NnWAOI1Vc+KXXS1RZyva0utZL+Dwau2z9UdV7hmUIwCjeiA2+bEjigOj00raG
641dKL71J9yka0v+P7SP5Zxe7Cz9qbToRcxDKqcI1VF2oudNiaIh1cMqK27iIhTdmVHbfTF5EFYG
QWNvvve3V45TAN0TUYKssl0lyNjgeBjYhrEfPKg7LlXs4ewufWbQzScO7yY84gXmGeA31Plc4DD8
ncfQ5VQ2EgBvgR0Tf9bT/MEEXmUd7fgPVRyLiSmraHcUESp25yaJV/HaI9W37/7bKZa+dJMKrpw2
NMkN3YLsjyjIzdwlovF4jqkIyvTfYemFAFNb9LWy8WmFoqgqbcK3qE4J5STdn+itPO/lzT/o6po3
vMcuIVcY4UkZbxGe7UVF9a8roErgc6IWTbWdxrkZLQGuaT9w21hcHUc9wA60h99ChTQMcKl8GELh
g5kA3SbNM/u48I5Y+LHpaTmX2isvQ1mFuhIMSfVynostbDk6yGITV8LTo78H6ZKjg/D1uVx4BwVA
g4+ty/WJbW3IXn1y/khE76Pr0SE7McpjTbYDXLNUga9mQ8y2bPv4O+N8RV0e5HPEnSte3/U9QZy9
6isy0FljssBsrebRgXbNZubd9V1To+o2qQcoRogGpGoH3HiL68RhXKY8AZkCAk9a785Q3VNJ707W
OF0HZN+8WQMhKPrahto5BhjZHxGT7LIaKWAHjay5DtkKcE6peoomugqeG04mbGRLML5APzqYl5+6
oD3Vgn2SLrGRoviB4vaDnflHXvPEZQCYxE953PQyMpLKbIkfmfcApVY4yy3kSHlYMzOdRZgtICt9
O7tRkvmjJ/35PruTgPXmTY9I8bAoXckWowpUB88iG7j6bf97Kwz1nDhviKwhh0iMi/a+2kA/bKqA
Rnj7VFl4YhlXlQc9hn0Xsr32HZ/rV9Z8jY8MQUoGZ0trHLqZTNU+vocp5GEkwc4JTi4+pq4znQEA
U3JikErT6d8FACsKyTOLim6bYYjdm/LAMjwI2pAfEGR4F0B+KDvyiehpiKteP5Ls/VyUxfo4b14l
NPlXeuPtZUHV87JIlO3UaIl9sO5P8Lo65yMI9QmQbfQwU/7JDXQiE0bLAyJazOeUL+04z/3CF/1w
4Zd2NsETH70SODPaMGXqT87TPISzi4LtSMOQ3yi9DaiYecED7QihUG+TnNRKAku+IQYUbMb3Bepq
QpP9DoroU3s08QPG/fH5YW5mDSvjT/N72hn5wag2Og5//ulg4sT7B/Y0EwuGbkspGOYIdvpxQjAk
G48e2Kjry8XSrSRIX4fw1UGLxnrNua75myRUbDp88ar3UCgTtOZFGGMGSXEoSl+vxn46ce7NrnHn
AkYZ0kMCQwgpvrCmLoziEOxjqG7iUwbZa+9rCUqR4rmunSKLZrYySjUOvkmVh2dSHt01pIRZSx03
fkAn1U4IyiGS+MNVQc+m6aYRFUhI4QOQOURMj00t0lH2SwO/kZ8gm7FNbkCYhlOM/cylPEHiiG93
rciyCir+xVhwlsDasUetlmDQ/TrYRdfACrWDDHiPEoh119V9Ku1uCKpgYYi4mHdEM5kbOrFhx/aG
liTNgfu7vLG+1hzGH7CLsduuLCZunuLQ4XMTcpx/0KYsaJ/IF47DjRmaVJSnHBdwh+jergVvniPI
m/VBgswV5Xts58PpBWI6wO/2J/vi6bQrIJt5EfmO1gfMDX/X3TXQOh0yfehhxpn5gUWwVnyofktu
ppmhASQyABHCBwbdbL2b72tLw+Yk9DEQEd/91Vp8QnbW2XeHGi1G/q+w1MEEp6xBFszpQaUXKaC9
/4awzca9tIqeQPvR3LJ6ss1OY/fT2AOI+Ks0RxiDipvoG2+Vx3eh4FVbTKlzjPI7Bqjm6twoe1nq
Mhu1N/uhSF62vsXSwhY/zHHgUS1NbXgx0qAvI6VgjhrknqA2GZ/kekjqToxhYXmwFKmz0WDy5+wb
xPscaQG/agSrG7qH1awrsjupwqnOrAPsPG7PXRjgZHumDJRkHCDGEzO36Yf5OHMXFYYJKRqQkbs1
eSx751dGmXT/weH82r9P9OdLAVd8PYcDtPlhqSMiW2AasEL1lYbQQHqTt7Zs4xk22Y3mjCw+07Dw
UdBh9sJ9QhyfBwzXA6oCCmXRCOC8Y0g2ouCyXczeXGlPL2PB6Xc9FpNTY5T4VASmtnr0gvd0CEBv
/3PfwiLZ/Di0dGoHO51cxHG5R4hXYmK1UBXqHATo9A8iOataGcMYB/oX3PuDxnoIm/4VMQ3lq3i1
k3BFQ9+hdKgLYXDjvO2MwuGmhZTqHWyzmd4kRnSEHZIHmtZTCZziB7PuQanqlNAMsoKd5EotRFA5
R/3FW4RAxvb9taoYbEU80ABpOB3G20wpVu5si8cOegrzO9OfNDlZ3To9XSdEWvhvQQ5dbdpvLrU2
EIRKuUvrxb4e3U18polh69O8QtZXakBWV2obgzKI0+/NwakZBCExiURfJRjpTuyC6uzPZ67ePD6k
3sFq5MTEU3sQQ5PsFyo3o2GezcUKfONUdEcb4mK9CbMNtBsY+rQcyljMdQ+4ub9HDVjBgB2I7Dqw
bnMgQoqRiKYY4dNJXhrFahw7k6puaIjepiPKtQj1fM5ToAEN5wXM3M1QoXoV7/syffWcOBHzxzZl
Z55ib3yNFBynPscVQBxkj3x1vVX9YYoLU6r7K8KpgR+xcjE19vj9WIPoBk0lHLprAt77MEMxJ7ii
/VfxHSolhFmwXYftUL4et+OtOpVEvCHieibuwiFKyGvvUd34OHuS7HIQcEDFcMpNs7FP4Q8OYa+y
Haly1NPdLyNo8AKKG6JMj53M/PNtRa6WWj3Kd6CSvvWMo9/dpdKc0wLNQh3BKFWcPbZfNQXExa5h
VC3HX5WoFZTibP7h0Q9YpHAJXUi8eXakPyxlSrZvFRiPysdVB4mCqblPwq+qEkXkkRgLBC3AMYP6
BjWDUeU6QcU9/SS7jxGqqXL2qOps8/UZU0pd02qKQhX1FNcjjYbpcrDuMfFu7Sna7tGDGbuqprDQ
yKXMVfqBK16WTnkkrVltWv7HGCKL3WF5GHrurewXD/nwAhcd0VD8dbaIgnPYA6+NoqEqP3zX2qIz
WmmPCbc3JCr9nLYwWUrEfKTnsyUkeHpjH5MtQBND2USZc9EVkESYK2SASz6XjiswyOLeeiVtFERa
6bT+9qhfhyhpWeA8yTHCcW7oyhoIHdBgwa6jCuS5DI1NzGPC+9bc7ykEkGdVHRFY8wnF9vVaQU4B
20sO4CiKosLaSDxfdF47C4EfQanY7kYBXopSRGX6M9c9xGuG+n+YeYA7PFfsEoCXeSQtvYLGovQl
etx/hkgZQog/OseuicMvCVpJft3Z6W3okkaauK2WFuY74BZYo79KGCk43W3QHrLxZscrbCegCrzQ
yjBsMCdB0VfiaXIe6hvRJqWuBXlAiykpKKJ8laThsFn+N9T9dSbujX29msnP9bdddWJ0ELK+ZC1z
kYmUejxpakN3r7GTHI8sAtL9S2tL2QHyPeLmYwLcbPNdwHLAJqww12LgblHhrbgRBZwfR/Yj53uq
e7hmoCir2TSU9shodeijf7ZLScEQzl2oxpQ4MCQ8oKIz+4FeEZHJr7+l1kl0axvwOtiDD5hcssxF
tF38AyziVbwx2UnqtJppwIII0YCL2DCOdtIoJfREzZ0MHMMt0GM6qnTYBoxNRcijAcRJrU1zzfjt
ds36rNP252eobX1sVTiBKhCInLRB86PlBkjSSyh9o9uKPQWaRf7ETDkcAGOkYcY402qG/l9QJBBA
rJnUtZDUtgUfm0zSuWY8us3cr/R47iqGgE1xpX/MOanGZ6/wBvqtsAqYpto1b3v23+fwEL2GfOME
6ZjkPnUn45J+r6xgC5oGXXw6CK49iB2q69/we1by7QCbXVfA4fcBohBkTTkorO3BYRUINxthDwBH
80aWpd1n5oS5//TCc+5Bi86LYWFaLZ2Ke9L5IBXU1qUb/vWx3RLNFBg+SbEkWLwDt1d7+fvpHLgS
lJiFGi5xYlqAh9xWYp3p+vuWQuxBoYitOx3W9GZmchKdifJm2zgS9UHuBS+GlSwRnFTVvwmKsaIP
BP3e3jkJ6UoJiYrTP39A9xe6/jZJ0HnZ+oR/C3envVZiLNk6U/BnAoQL5BZnGs3whVbkLfdDVcp+
Xvf6lVIAw64C0Hsb7OQ7AyPqxyYU0qsYVfYP8hY3M3vw6pwYj07VJXBIUwUhHcp97nO6BaeEAvzM
sV1EUsIv62R2VIcqlpxIkyWzTUqTt0NSXCmMesY5oYprgXAvCZutyw+7HG5uFDi2b9NH6OZ2T4Cb
4mfZqckCwBF1AklN3g13qUBu7ZUd9Zgod0N06qtfdUMSIuZVLI6am78GQW5kWNliR3VsovoCXu6p
KpVrrSENhEj133JQyvhmOTFCU5SVUwDnLcdaC1GWuP9mpugyh4ef3D9WsRLloeD4w2ryg1LX3t7Z
VRLmta8Cnq/9O2pBAiYkYkPpF73NgAk6hfsQka67haAtNMeutbK5C7B+vwg8avhHQnZ+9GSe8wn5
1Kzv7/hH7mSi6tGwSz5RdCwQS5JMRYt6HQnwBV8wOOjpQeCXcC3r2f4yfky7az+Sj8R8pIdsP59i
J6awa/TSulT6KYo2Q244szUeYM//+ZnbUwMsP9UPcUwoKaoUA1RimNXQ6w3JsH7MBvkbYcj50f8G
dGHKTacyxlOFKPxMs/Gd2mWEzJk0RiDgUw9zbzieZ2MJ03QUF5HkYXsY9YRJc0N1/Rxl+/7FK2n+
/xekmlqFB/HRketaSsmX7PXkQ4e/LoREGpwavdUiFhzSGcpa6hp3IbrWhrEQ9v2u+u8/gDsG8+tZ
4s/YA7XddWMU4y4vU0QBO89sTOroOmAEYe5yg+FeX5d25C4helXyfwzs+PigPC8qcIWlyHSismZ0
8fZKr4/SrH6CFxY69epwwOCvLVWgQH9MkXgmsA3OoV3+uVzVOA1dyNKDVSrW0RaVSRv6WxeOwmVR
pJ1yN8F5GlPHOhAIWHs67n3P1E+qJQrgoHuB3phFNJrgmFJiZ+mzAKy0bCwPFOr9lGaoSMqjIUat
EwV/L4LZvFkiAMSz34iZeL5pysDognFYXydeqnT5H5uJYD/sbhuRH9MAg3+fIYg1EuJVSw5qza/P
ovQo9Bw1H445Bfi061UdNIzZo6glwFMApiQuoi8h/hGtrN8d37VyHj702B4elncoT+1idl7il1OQ
xLKgbv9b7XjLnEalf/YmQ3Iq+T8Tf2gz2R7A8xlWVSuzNAI3mF7V3kh5I8aQ2P7bXxKYsGOJ7aD6
LjDLQDKCmzhZ2Lye3jHsNVLI4IDmcw/yRs3XQCyFUVfHlBv5iCHObf/4KJcLisxAyX6BcY8BWg6N
KghTNqtAxYKh56mj+E5Xnldd9YBhchaSitZDiE5vAdmLXt1YRcoEZGEbQs8SsceNNH/mqoHNXbOD
ELqNaAtFmSnHa9knf9YYFH4pIijX0sqKXQ3Mlddomxrs7bSgg+XAnHFIRQjMYJ1RVCJ1AUxDT7mo
X0YwQLuuQ4dQ3crNHtc5omR718ujFJqAPk+H70IRPUU9oMHF0y/g2ZVdVo1sJ0dO+/xX61d6YTgg
cjydRa+NI2P0sL2vD9Zupg3y87VtN9X1V8gJSU1lz55lnPjLAYvBgo+gSOxE7nxxrzcX5yMmPKOy
KWnle0TNy4kHft3JBzZG8ryKPrgIObu4sNmNc09wLGmXXBXL2V41Fp2128MoUVAaILyoZgQZ2z69
TxVUYrlHfTwjFC1lXbf7C6jEc78nEm/WOSg6ToK91hshaRDjlUg4gPg8H7cqnH4tnwyUsLMJfjkr
3tvSbBH+45nZzQhsKYvX54sG1EV2vGyhBNYMOKq7wttsco1zoTNT5mhcCdfBTxRa5Q9okvOFB/Dh
TCYU2UQ4CdjX/PZHIha7ZEUJnaxjSaPm4juhrCUX9t13TQpLE5Yn0ciYx4E88m++0VpYDGs/4M6Y
OJx7+fQ6TBKTpPUbGCMEr9rpc4vw7p8IBbo81ARXT6S/81lc2oP5zSz6pbHkoA3B3M+r6Vz5bGtq
9Uu2JuAKdN2ETTAKLh9YGGEyK2aB/pNUKh/XbhvL9B74a6xAFfG5NCMwMo3JrZ5KtIpbEPil48Dz
Q0XQVFJ4g/EeY0szm5jg9JVCbpzbAIgFStONhSKfXxQwTDKhpbWVkmI86mG2sx8hlqwyKJLM7IQR
7alVp2hzJ/jRrYwajGnw0cSHpH2T3ypsdBbmPwzUyhkRxobNvbHi7vS7e29orm7UlH5aXgh4DQaO
pvrBKJeRTSQ5xmchdijoaSK6WrbGuPmOSWGdXptXIvzdRed0lXHeO5vQjLC4jVS15D7sZFqfOTiM
ggLhoim/u5Nj05uPHdVkSnbZ+yKidET9KE4X9I5AgOeOR5jBOP5trHugk6awbSDmoPyM/PAqcYMG
AuzPhzQUXl/00p1PzLv3cedw1GPeZLCKbW8/0/EQ+8VmMRvmxuHTLowMyG5zS6wYrTFd8UysL7By
/i2BpfqT+Pg0N4iJGh3XJ9XasrqY5LlfOHDlR0aPQZNlvTSIs1pWaqY36wEZmTumuiKcEnLQOzdO
6zUzJwcuU0zeCON9wiSqeoWn27e+zxBy2v6yxLr/obyEbbjaGFC2b7hAG0cyIpD3j/JZo1rKus/M
07Zzig1CtJPzJjzbv2S/llvAHOyRziS8DaDSl9L0+JaOhXrBydhVeeIEIQpjdRWK884cweAishGD
TO5x+lyzDXg4AE8nIgZ/Drd/+kRsgh2pvA5tS/QvCYwIjPZaA6B8f7La4c1igltxk7TwpXLukXKA
lJJt2ipcC2jXvfyrtLMaH/baS8tOIs1VkG2OL0g0C80GBtuI578Q4j5FtBMWoUJMGY/Q39cwZHFl
onXwbogugJEPI1TYa9Z6FQeVEjSLBjHe7pcsfD7w0UwDf74M1AlZOQ+6M+SMltn1aw5/nDsKjuYH
RttsKgkc3UiJOjD9G8ClnF+F0OVsaQkoMZHcmDWgQv90Zy5th/oVnzERITACJIDwwtO5KtuIwxkB
i5ZVeONcUcTFuWf66jW5BsDddr5LlrFQcwinP6V05h6EGtGdI3Jp/c0KXn5NSBPcqulljwpfquJI
jCAueAaem5ljMIVYf3vzFTpN0LtNXCiZSH2N/FDwp+Gz1n1h6is1KBwW82ifs3w9ApHF5n1Ma6+d
5yqCZg8dfaReu7c8a3d4M6OMdsSK4YiPUEbwT2/o2c1PCyU3i5Kuh3vA/vicqDZFLh0L3VuwvPfb
UWmLrZEEFoLZQTmmHgydwtfZc0oUHuqk1j6Zz6SrWmeLpSoiboPgfaBqScKxH76Ch5szi+lDezqY
uKokbbYQldChYyShDVjUoq3ZqsDVg+rsTa1V9Zahn4v0nBCuh1aHRpWg/LzDMTX27YMmrpedxUMZ
ZJIu2GUJJuLYRmx2DKqLaGgI42BaveyFc8Np1UhWJwEg6mcY2EOuc/4e9oQIX9CXzQBcBhWU11cn
SzMphjGbwKoIuJtisYjC17Y1LVCDhtc02Ns9YaTcl5WX1bE6F7JM1P0X8zb4fTvvjKPD0MhUBco7
JXQuk01h2RtK9JGwGKN4HX/Tb+rN6V/KTWvBcgyxpvpC9lv7WGmOtL3+QgttWU9uk19cDc3PH+W3
8EHW5PQzsYBdz1v8lZm1uK2Gyn1DQxDyIb9YUFMZW03yunqlQpTk2m5ya9fovQ3d+avvs2Gxsh7K
Dm+E8l+jTykIakLkybF07hc19cDQb1xw0yihuus6KR8WzycEXIylHdHSpRVFGFZrFQxm/tEfmz9b
YBq3LG0RVFP51nZ6u/J2uwIWG5OYqEOW1d0MicRQS0Lp6BRDrIET0arasD7i6iCjvvC2ezDmASCG
88gEnTWopzebLYL6gyo9nKppFnMXh6RtrafnYtv/vuHvv3Z6sIJr/r3nVzejioBhIP0ZD/WWjE4z
0N123bdObUPFTHMFohw/HcePVhK/LS2tEhk4V2piOOT/gTalK5HK0iDmuBysHigTEZKMsbWydcFK
fyGCSo1O7tcGyM2saQUOmIvdgyKHiUP+3K6CdIZHDLUB/J+XTdHA1o64w0hhdI7I2Szc5ju7YW7c
7wU5ILp4yXpgLs1843lNoHqtp4ObuAZ3EK16IwZRRP4DBmcRr5sswwNOly+0iIf42S7NUR/KkuMg
6hyOT77stWMUOR7e4M/794sW9oHXJvyqBOgL6zSkaZjBTPLDtJCnw/ZLvPGOcO3qJVpztFP+q/2U
dzy3ThcbzuLqU7Dam7r1DtdpamuuhaCThkU/ExLbtTOIDqR+ItxEwteUJZQmRhkNUWkeZ+c74dui
qBLCogenHmPnto57uwQe62enFd2hiY4KAAWyfbgEuqvl1sEahotn8voxZvPvynJeWhHfoHfoATws
5H7W/3xPGofLi6RWEbNOZ6ismbHkRi3cVoR4w4B/xJVHSVEzb8wGFyy3LmesDNb2puQ2IOsYiWJ4
RtfRv6CQBf/2o2JduwQVy8RLAcVZU4MyhO0WayonuF9zrsNoOyfWrx+a+S36dhAbjYDnRf4S/WMZ
49xoHCG5dAT9o8p4dzuA71iw5Xz8b15GdwtIMCpoH73y3hEqHQGfgUhQyfUh92UDW4d2Q724CwYf
zMnwxVhxB8fu6Jcze/eRtzHwmRDGIi4eYy4Ukof32q0K9p4MNFq6HZ52N1dR1a3SbNBXQi6GTc5a
yk+bPiFdj91px/dCAbvIkUGDLuPAnZpTqwplCmdqK0FV7nUbuXS/JltOh1QDk3CvZPmjG4JXP9Fk
j7nQBKYphUmHN6wRImFpiT41MSnwXy41AQyvIq8byjaASCQDWmlzWEZKNhHN/A2PddrwHwLaEJap
X428g7cfQmdwMFr5/GwjC2XP4ZtXYNnO3pRj1QfSRIQrNoa/Hg/aNjAKIDuUgxzBqN3gm6qUceuI
CrqhOYv5GbLEHRTP4mHyZbW+J+QWpbc78j4+P2qhtnOxcJd0lbCfGuj9ukbpms3XhziViG41qXfX
kpWfdb5FAyb7ka8HbuPgnFvSOwefTR7tJwNWJqfh8ryDM6mWqQLT5UWWdHfonG4Jq6MkiTiIE2+t
WNKu2K9Q24aIhc2w4wt4P7TzovULH8t2Vwo9SP6RR6tpiLbHEOuqZCrDSeYCWdXs+Y8OvUHPQ9uS
5dtEKM3+N+sznxtBOROe+urFN+JiW6JwJ4oh02bsq/RPBHfvpE1o7Y/hIplgcmamkSbCFhXuDwdO
Tcg/hXegnExy7XU529qNDbBYI5Mxd73o9Rbhp5sxm5Z9NRCO4Xl46lS4ziRh27bQrf0kqZmZ/hYr
E1D+3YAZd3OgWOFfhlrNrT0AM+GFv5V1wrkdhsXs/s7iTCP8qex2ga4w7GCMhtmQ/GlzlcNfOIPd
K3lZj0KaFHpn5y8VlSfhf3EXygw74G9h193MONG2VQhLlrDfwK/OVZN2fEm332hDD/sT3MKl3q7h
LnMNiklx2fKC9GYT/XizjHqNq8TmQNCPw250xpbFMBiTFxdRdjY2Bm81ef7tpQq0VSIkrKLscuwU
D5YyVepL9FkbZpiB8A04CWWF+lLWCaRH1ePkLVgM8CZNhKXFh9cNAUTWbGVre0hb3OhIS/VZJF5P
usJKSaDjiqp7Wxt60szkeTxYOjY7uXiPp9rtUd4wPp6d107UxtmPFJHOOxEHOVWfsKZ0LYa/Dhqr
mOfSl3T8Ey3qWjBymKR7CPiIM+elJSuTWI03GrxAIOBn833dLU0JhALBx48l2nU7oc6uKLhfIg20
PGkEZUdYmZxwtVWpuRCT0ba9ZVCWAYZSo0V/pNLunYjx9FDVzTGHPUsmBGg6lJ6/RhvvJUAZkW6p
t71yEZGUCpBuuEE9yBftHWv9mzC6YpvGDx2kJonX6dAJnfSzWJNuP2t7P5OU4/ouS3gDH1WjM3bB
oi9QwD9TINtAGOT+cbO8FOx2IK5j1xX/tD0yeuSTrMkRrYI5vicS7pOk29VSxmmaUdADxQP1dN2b
uKodQNjugrmts+qTeVkX3OT2d+IgQXTbcQQKVbrYqQw3NMRmlgHaYSjdAoVQLiBzaqSV5Ej/5fq6
262dYqDpgYPp68F/7rEypqBAr+RfSGVjUieMmByi49QQzSgd6Xr1u0QqPVuwdOJKTYnRoEM6gDfq
Z1JaSwU2/2JUfTU6FmK2s01Bnkjl0pyUib85882wZZHdcpMtOe0x31WL3VDaKkSu6wpkR2CsbDX4
w3ZkKdTIUpW/LIkfDb5s4x45TiisCGXBpn1+fWbBwWDER4zMKFwvH7yzcdhtJXJ51GwKUf18Mr7z
486BpHJ1lkV/zxXbSfW8yN1XV2obZ3XOirBESiz1EzQuSO8xkKRjiwsEExF4TN1gOl2xPvybe1W/
VyJlX+GfeoJ+/z3jLgtqw9ARkm49qcMiDowkAtJcF4Jq8egm+ffgKH+zg++PUdh+wxRuEFai5hPl
udP9QSvFrHDSLFPUeXKcrrUzek5S3ef5tQuKsFoOe/go6UIkAJ9Wl22spYlE58uM+kGHYAqzvdWS
VxOKXJc+n7nNsAr1s0vi2vEe/Ofx3/+5TVuZl1XxR6KrNufcuGAlvpACBGMBpDf8ikQm3H8/Rfc1
yxblK44drtrzYM98GmUWScP0NBV4s0mZ4ldTjwAYjgRuIUbWAKyPAsorpNwe8eBbjbKC/TQLN3H1
/YH8zSB8QA46K8ZoaOFGalqgcE7XY3Vug2uuaqJUDAPlNTtSXGEu1CSAbNdNTUkm03NcJP2Kw7wz
W25yH7TaKsVD9I2uCWnIac6zdUWDkp1nqrwKPpbL/l0r9RJdyPiF/62OXNh5zZFn8+tou6mmHL7r
LOo2l1/ZxXzamsFnfoS15D++pF1EiXPaIcPFGwnGHajB228pnhwYT8tTOGm2nAhHJM0fRrDHFyOL
W5U6MuPW93smkT/C/KVQez5tkLCo5JGxoDK1Jv3xa8zfL+BXkq8BwlGXw3aE90AntAuYGXC8hFXz
lGF/QSNQ7DUlM7uf9l/RHbkRpgCKPgw6krHu279LJpNlDH+O5XXY5XyDnYySs1lO3pbq01QNFEgR
JnwGvqMKRyQRwp3Fzipz/kAJz8TdW9Ok6ng2NEGz21kOC4J8IYFol/W1+94bwVe5dzL9qsRWbB48
MFCieNjer+spUE+5mqCdxeREm4KfFXQigYb5n0r//kM4T7WN3XzMQv0J2E+jPIGAXtXMAPfQlGHg
TJSwBRYD7Kd/c0WJ54THxyh62jbJoQhpzc1j+4dlVRPLsxs/zxWQ3DZl81YgmiAgpKXLkgA/uUho
nX4y4PWDmoknUhp0/ULZGmnX65KmMKWmrchq1fZ0vLumSmNHXByDjinkrdXGzmtuFfE6F2D5kuoo
iCCIb43aEDMPvaSkU+HPvfeHRG3Cm4DkkgxF9vNl0teKOjQ8EQIk/nzcLLjiJk2/LXt4/UG+KRJv
HkMtYtVdFtmp3cJiashQbfCbpO5BxaY5no6B2dn2IBO8xH9RCSiOpJ/FwzA9qbC0BvojxUD34Jis
M1N6U7LMpgMvLvDCXZjGPteGaumreenSBkq7KWGHE51lctif8iw5ib1asQ7efmB6ViNNV0GSggMm
YcOScmljOmVZBPajuWDRWQgyXScQnKuTrX6LCmmHtnpc4DmePcoOVNwF1ssrUsLB/AETFScdYT0T
l3SRmLhOxWI9hnWV43wvkc8VcHQ/vnxC6d6mjI88mvAro3ZTT89zFFeqSUr8Xm8m16W9OSwJFtaA
8J/JJuXFwj//ln1pIbsdH0cvfEzT7ObAwoHjndqkJ3rXxEDJf4tcq72gY4kYCADOXpixpc067LAc
DCh/geKbwZp78t+kT0+fP7AM49ijOsX+i1Yk9iGlaNhyXSuMzZYsxcsRR+LN78RKj8ydKC6ZUXYW
/z4+jH5khxkx/Q+TJUfdVk81+22UFKs1MOObfXtoP+SOAnVd6PSuHQfxuMQDOYlg0Y4JU2Y1aWTI
H46Rug6TI4RJKb5rm+JEoya977wdaKN2fwMYsc6M2TCsxRwt2TgzrOF0yz/JHejcTyOfvA3o7Gpm
3gLbIuv8ZCj3xWTEL9G7mIGVb6efij5KprMtcewZwG31yLJegS5RL6vJ14T/Qc7A6QRyhzS9CPIb
00Q3RQ3Dhscr1vbkfumDy141ydoYC2dnb1fe7LqVvm9wZ2g7K1b50YIgvYsMnk06GKJ/SNfVUI6x
E7RvRZUdFpLaAIzjJLOetVMaG7L45F+EvxCvs18b3kJ6sxueU9KdjXEA0K0TufajCpi758pHO6f/
azLD2RAzPU9DM9v1XXyx1rufN6c5Ux8icE7Fdepst1BG329ZRtV/oqRBkjoz/xL8XA5dD91U3+0y
kOMe99M4Foo2QPZIL6WzjOBli00rzxpc0sZawbtlDAVg9aRQ1UMqFHurD9jRnHKqV8Jtm6YIxPqn
SH/lm4nhSj3ze021cYrrhaprEC/O+GIG7+oXcXVMqjyD4jac41WtaYAxIPfHboQzSfRDaX+KfOn2
T7Bpb1QtS/qtALC2l4OrlTALTQ7WZ06zTWWmZMqVkP1AvcT6JEd+3qfRZ+sK9D83kJfdrIo4WceO
gCDkl1g3V2N6dlcep+cXCT6/o6e0O6T0eIFPbqhVwRSbWGacXGCB+TsvfzrIdCK7n2YSEtsk0w5J
ZIK74Kfd9YnTT/zyEG+2sHuLd6mXcWZSGtt66uLLTCppzCEqbBCTsdzTKA3RA/ezdQxnvmcoOnwS
oR7gj/kCFA4oYNd6lZ4Ua0ReYcbjq8jtfxfuO82PVBQr4gsy8PpPxgbz6p4lBMMwRc+S5d8Ml4/L
b3N8vS+qLBTGPWW4fzO57EOyVQyYgCsjPkSQMuftbFxOVf/tL9ie+gbICK9YzToFl8LMjWMe7juU
oOngtpeMKewoekU4ivH6/zvctHT4riGulFtt2iWzDpPttXA0OwV2ZjVH9GC2sps4a8LiJbjGS7FQ
O4X1GMyhQVxiCbo8NntBQk2HGIzOzfsWhQ4xcSDRABN1gOP9UF8xuMg9YT1aRuRG2fyUE7CbGMtr
TySyCEZmjA3IsPfzWcwMfkgREFgBd1MVBOztOVttuo/h9lI9TolXvErIzY3hYnyexia3IhqPW559
xIEjiZGz+M8EA7lFyiB0HQ8ubRp28FsfolyfV+GcdCiItBSaQ9F1V4jIUw6uaqe5+v7U/gZ3JNfd
ZlJfT9V3Lw/FLMpaH49gcgsIVdJzRfQbzu7TIHCETjwqasR3GhIMofmmYcUrCxKhK2M2u517rXdc
NIWkTquMnmTlhJE9AhAB/vwpOAuwKYVe7vPb/6OyFuMXV7kiibL9GFxHEOWw0Gbsq2ospCisZGnE
BrwT3I9Wj01jv98JUN4WLyWhzXuGNiyWmn2mzqAuEs1bqJj42bLHNsufPRCRd5JWcCKadC7Da3cY
+XULTxlozXXkR0rKLZJM8gflJi5LXYMRhNuX7g556m4SLxClqN0K8sQfkWcWkW3OKn26zajCwqdr
q+LGkAFNSGtJdfEWvUxHXF0f8liV7Jjq9o4OGGpEjgy3DxYjwaPm3lLm/RgOLtvC/BBNbzqJ68Hb
xjOdscsA3OIfM4XDvPi8QmwP5jOmbRRbT7K1hHB06cpIuAoYYHYSQ0wnnjzTiE2KslQ/eTeeRJRU
x48SHGYP1boxGwoKETaZCbxIGy06PrCnaqlC1FX8Q3UUjDu48ZLqdGxb38GxSFNlJahQKtyPHp/l
9gvKK7AycdFkDyoL1djM9K20/D+9E0OU50fBy5XRCdbLRls7oEA514NNuYEco8AG7DhHMD0rk47g
TiC5FMppyQU3V6ZkuNB547YjQk8BtrjZmlx/DHdiI++7EaBHfV8HxxtFcsHPn1lCGexylfcv/jnt
3D104fPdTi4m4rrM94H9M+HPNKTMhobeLghs5P+Nvcl+rbqFtkj97Iheun07/eTzwijU2/29PTXO
TYv5t4fttpAE1CopYA2lgNBBPKpIM/yjn6X9ni2TFb8Ls3sCJGjr6YngIvcRDc9tOMjVYDWM1gkt
b2rwERL2Nf4U/fOiOcp0Hx2FnXAHJcLUR+cwbtioqdYkFlohPWtOoe/V1xBM0fnamY80Mu535aLw
tiFTwSsfTpxMtEDl1bgnUObX/qU2WofnvIkoyJQ7Z0tAVHlo9FD5Efr3t58nLhHl4X7AMWW+pU5r
2Tn7+78EcuA1JvGLGGR1pNohMZed28xNExIXw7XtUKurIjO1LzJxGa9Rm+Dniu0gPYxsMwcGWxRX
5QObGCWtG6GvDIxsbv7UjBSiVZ5iBqJghHRXW22bTZT4Swfxf2OGuplgSU1EvaAG/6QUCIc0FhYb
6IJH6dYClJMnfJb4cdA1HtOYojY1dhvl2nZmZEGttypwjdpD4eB0TWj7R4tReFN0Hefx656mc0Xs
cEgXJY4TOdQuSl9Y9ZY1HLlz01mWo/0FUBIbi9nHl5ddxnB0p8nk95Kgr+TD77tTAwr//hdnjYC0
E+8UC5FYdffWYTSEDg7pG/B14Fr3wYyzqGKCQ8C370vAnIO/1LOZX223Scg/Qq1ENWGEzrknFeyH
MRbLp+/KAhiQtkKMoAaQCU/w0LjfNpkYqIxksqniuQM96/FzseHr07bwROflGVCvJn74DCOSf+1K
O48Qkgo2SOlx0jI7/gYfs/eqrs7Oivp04VyTMI94fzjL9RMH2bYpaj9zr5867a60LjD9qI8Gqi5X
ia83RhQvIF/2y0kc4LSLlKUyqq6VNHm6yKZu+8R9BgEtM8sTksGhTB4Enasrs3t+8c8j0PIyZyO5
gJ5Sbg86ECcXrp6OLyf0rprH6SlWmXSfmpkxur/Q7QnyYNcFfufyN67/i3gm7p/igNP1h6czCC/l
FR0mOKdHMTBhpnMkCnlVI5LDS3nKYhyW7Z3upojbGmy+KRWYqp8vB9mO1HkVvhBRAU7JgZgfkqjB
rOiYQ9oTGsQLxEbgnbrnOSbalIfhtUgYcC+6kCUH5VR8PxMKG+llI3GXMvwomxqOm9n/nS54xvhG
p5dSO2cg13Te8b+8nevdt94lhFncw7Z/Mz9mmG3k+qYS1LCd6KCROeNwu0Lgzh+yPw3r2kuhJ2FH
EKeuJWkjD70HXBQsvrvF4vvJOT8JknhFDYVGPK57c4/fUEAuXyIPg1v3fyoHOqyvUgBN2Lvt1yZJ
nwyHiwhvB2nz7g8KaQPGMh4R4YDdyoIlnDExw6ih4JKq/4k/HBNoYkaKYAGdRe7zti0tEjZ4+Q/q
8T5QP0LAPzu3GsE9sniP/N6ddzg85yE4SyCmUAKoL4n2ij9/GQQqKjZaCLafuwoLOTNRJ/LTP4Zu
Vc9FYx5XB+J4srLKEc5Sq/3TcuJ3+dW41pF8zaWTCUeXlmPDh1z0uCWV0UE9qtltum7FWi1q3524
Iqp1a1t9HjnFAju4LaobcKWzagNr+KYcm05Bq1BSmlO3+jS8sdmjIUFgRuR1+LxH7DltsgI1DO4h
B/8kTCkz7PEnsv+/G4LQo0tX9LmOOkeOTJDCP6gg8WPAyud2MhE8r5olaG/xW17F0U3CIaUQeG49
nkJe5AlYzFLLTwk4JitDX4PWF1TSH07v/lBCpJ7YhG+hjp+tsI5FUOsPVucv57ywj7Vr/3sap7c4
xg1ad6z3hYrzdYLaU8nZ1fi+dCUkLCnvnEAjFPICfcNuNASjL5QeyNNCRb0GWCenQfo6I+x+OL5Z
hUwFZuCsh8JQ0fjzcB2n00W0cBMPQ2/JqFTGDwszAtgNigd2ZM6GKpHnPKzTFMR1PyO2hTMDkWbg
GwyUAN5ppZNDdRPgZ8g9ih5Qz1FGshIanFikXgK1h318YDEcRe7dmRCinm8ROHb9xuQDOKNUUuLA
1gbFJ/Xa/V7GIdK8uw5IAjfJ5cCKlWWoOz83XqXQ6cv0cTTORVbrww5SilU3spl4qpwxGLLpbvpA
OoCVXfkD96M4YrAgwsw/YZa+P7SIFjQSiW2ConIVg+t3TE+Bbk1MntS4fy3riGHTrBFZOfuYRit+
7PDI5gX+XUhE+0Sesd0yrHYROWenPWEuCQjZyaXoF+4lhG9gct6WPHLTFt7v+DRiP/rOkejHOW00
CLKtvGdMj8zl+I0SHFWQRSUgRbqqx+d1K4AJSxNvF5KRG5+zDcAg+OErHOo2U+UgVtLWIDr6P9vO
ul4yjZ01f+xsnCbePxJxq3/jN0iOy2llA0tye8WQ3bU9FEm1CoABzeGwbBON25A4YVqAEkab6BPA
FG1jk/49TVPbT/iEXV3BGnzzwen5b4MbJpmgnUr96bO1qQGbyEx/17pn6Y+EM2rLfwLlzln3UK7T
zfwrJB11X91FJkFw70JvbvRWRKYUMoBcXFwoHSIJ/UqeRY9CEwEvP1u3Dk7uy7KaTnTLHIvZTvF0
r1QbYorGkR++OhgiDiFuPkw2r4EsdwnfI0rnxSrEthQSqnaptyfwj+aj92vpoOH33yFnsrA+x3xE
6UbCxO+3huvs4P8FdCmOk3aJL1lsk0qlNeQuxRpOY1ToPn4qd2gxvce9Y5/H0NReV6bJ/vnZpySm
0490n4aLZB9ONnHWH+Olq7nQoKdDzti9dbCjytT6rsvlS92nWCmFyQSLH88vo1LCSlwHnqwANot6
pQj38No4PsvM7oky516QgCYg4/u132VvVrTY3GAGgYxKKKBkJ5OYkbXrEhs3LPkuv24xjAhfBaR2
NcguQbXqVzYlqYrCj6CA0ERyRICSTvT56TCUW8QjOzuS9KaXEdD+4ksd+CssANcFbdqTsi/+wHPD
su8B29cJ53bW6HcNUf2ImBeF3cjDiKu3gV9f7Vh8jjPJRW3qnvLbcWB2SV8YjV2XYg6Nb8S9A5Qa
Cs00chRgguNfhY/EgKhAU9LqW68LncdjKp5aBhmpSuhbTL/UuuHI8ugZX9KTWPgVz1r6RpG4q4k4
soblFDj1kV5fdt9/hP/q9LFLtIWWLA0D7KtcYLoJqLBYECyzVGDFPz1eaB00YN1/cv/8Rd9y/Bdd
Y+WCPMZaGWeDwbtEdJmFyXUlSEGvXDlkVYhNG8vqqz+9NT+lgLbQlaoz8c8gccXR+NHl3PsiE0UH
IZoqAyoF7Jaeq++GkTpcZTQXeNXZLfdyOPS9BuNJPk/LBpTMPQ4yYHpRJ0jNOxxJrpBSxig5cslY
T7TjubCCH8bcOeGvq3cvcZ0TG37Or3RSLPm5ob3z2WxchNG0z3/IlYeM7RpzEQYXku+Ldhg0SS2d
k3JpIgBh0D4yuhVjIgTwKo6PkUdSVr8vhlGoYNWD1lgzjnbcmKJmCqrq+hwnB+zvS43nqcCCLmb0
NUc2UPBq5RnkRFj7hK3nG6xwe06tMr/9UFrbxyijtL7YLr2GrinNmZchi7vpuX/hKKSpJ5AFDtn/
nbK4IpttI+kceMu7asT71i0weyYRgP6tMKaIml5nbDCGvntnJSaqnkWcpYMpIbngAYavT7XvnYma
RTNqCOlgzueVgUfUD9nMKJwg2Ym7SGVF/4wx3RcrldO8+0rcKiQN/5yGoiex34KcdRm+eBAmNxwq
b88g6drzsA6Ajdp/gP0mc+IvljFI939t2DFpW321UwCMVuriTmPXkfrnGQb5GEb2uZOiYQ4QEX7l
dpretU0rHUJT4FLcL6kaJmN5a6GEktqTONCe/Qn5Y2S2BqMJDki48OmkcgkWbp09lQwnIBQ4FTS8
T04hRVXiU9jbwT1QgYOHURDo6dG/62kV4cn2omnf4a5OkxqhgBv04PeDHZ8EH6HITvWnsF/uaAoe
I6N1yFYigCPVkK0SOAVcQubCWgAoo7/0C9lVdk+l1NLaq99c+F3B9y12GhanxRiV/wObTlBAeCPP
1gcfq+D109BlMEy346jur6uyOlGATDhJTpYYjTgDf/VWpBj+2m2+QRQ/Ag7qwAEmWg/fu+mDC9rU
jeGAiua7bMchvHa5741mQ/btrpFzPt8q4Hd23hIppJ87UJgD9gBj3FurDbgp9DbX9Og4jxQ+qR06
h0w6ucPGifu1bnXIBtXQWhtjJcQaKN91AQx9hptwb5wKsIEaiLeWJGGtbDIVQVJKkUsg4rW5qSKI
smfYOTbEE9klbyjkG9BgUU1SwEEe4bBa3UXGeerAhVcc4QHU4NKx2bWmJTXH1RwXjw3PSTDMHuTo
HEWAdp9ZDPyco08D7qmEB5/nVbLy+VuW2mjqGcPiX6JXqxtdGIY996No09haBw262zrM8+jLv15p
aqDvTn5e/VbXxPLeosgGvymn42shzNk7y/rwfjaTkwJH5e2iOUKuUztBwLNdeNToDE1Bw85mfhU7
Gk/gWG0lszgntWxkFXmcDRTlK+EzsW0NnO6zGZx5kLYY4lc/Ygc/1A2bad5z02HI9xLvW7AQQh8t
HymOzMmw0ksupHRzi+LGgsu2BulwQEzEs2q1+kFqEG9aWPmoDHKrB8LNdGGBxCLS3Yz2y5liVdhN
yvFFs+/BjVmqjLZjvEmDMp/xC3SgusPoinedcurt8igPHr0GxQxVsmom2YtgUc2NQEN0yv8oLAZa
PYPDlAc38c5XzSUTpr4PO5SUFSVLYXIdnriFyP8k7E4ikvxQ6duKKDny2goJDikQghle9cMkUGzt
2166DlYX7a6AuYwygViDmjoAEX0FviKaqW5ZusFckT86s5+96YXje9CcumCI0BERtNHbvVDxLw0z
8QWG4GjnpVl48RHXAX/4QJUxPLfc4ied40p1935WgN4WQ2n3B4sQu/VxZ9qMG+honG0w20Gk0xLR
nYNClHfTBj9kYQqjYoTArDfr94vJoyaNskNqBH5FyJkwabwtOaNuhHGl9kOj0s0vCTa7VtPDMFyx
M9dU2HAtKLvzOt+dT3DYfTewqHvEiXd5EKsjPW+tSPI7MmXTUEHhs10RV7OF7P4v+78/IyKKBWW9
e1htrQoSeYZGBljrFebIiLWDAsCoojM9O1v335sb0A7urmgDHQw6u1gp1TiNbH/ga3KBk27ZD9eJ
e9tO2rpJ9ipf+ayZ9NGiNJ76UZM4SRCatXe4ZLIdhaF/HuYGrC+P2KgV2irQuCG+9OE4EE65J23t
OJtncGfd7vLcaq+zmCqlaKjH6g/eUOJ/F0gKS1RsgBRKEQrD0khwlJbzahTNOVeJA/4l9gzKzWeU
B7DXXF6mBPhnzUoKPiWu5OMKYMcMccjK4mp/7lelOS5aTg4ktXOTKxEtwitHBCRqeWoJOyWsRDV3
0ATDSFgqzqNDP38I5pzV2jEM3vUqM4OKPZNiwYpgzH9G+7BSnJTJyYG4xSIpgmJ5EVjXFh1BPS8S
4acy2eEc8W3zRAAXtLHm748aeX5dpaJ6TG5r2tj39+rHlATTpngaTQIiglk/xLx6PEldNHkfNuLz
d1l3fIakyGQNjjo2ct5OG25UnmW3KIWrona7WgNl5gshHUI6veHREbAIxpHDcnuhzLh1nKWMxfqW
Jne4nPOrgH6P4M2yFmkRpgqZe8BZ/rltTdsRoeXrBXvGOgBzflersey6Pxqw6BrxqrH+2rdn/QvN
pZldCpvU320KZQFiMgZmX6T362yvCkrgaqKLZ/zPxxY6axAyRsSVPtOfrSNlFNi02fBMQsD1VLj6
UxUYLQKXHRbmw+YObvcgC6FhxEkWp9oRJaHhx9bFq1xNOdjt8nrn6ruI+I3il4dBfBHkRQmP3iMU
/Z/edtIcTaLeVFaOyQ59ibhOSK0o5S2scVMv0ubmttHgJgm72jykUdMlFIAx/7aOXJNyOpLV7nTj
MECrvBT+3ZGK2juh5Y5pX5vmGC4pEKHGYA5lQrEb0PwPtR/jGQ74CTHzwmN39SMhvDg7oPDjeSXE
2QJ25UpEIYnv7GWhXfW+6LegKg1yzVk+KtO94z7nitK4y/YPk1Atchpl5qybscwdOaydGKc2EGzg
w4u5dlGjl9OWOwSp7oohn1T10UNCmxy3M2uJzccnVcdnVI9qlBAT6PcCDPIbyzWWyFwT06jLVfQQ
WN266r90X0CA7lEDpA10aLCvmY7uvQsfvNkJW0ZXYYrxs0XqKV7hgI6nW4xul7RfhA8/vFtpIzPL
idw/JeFgTj43G7XGTntFFWBxQmd5apNFL3aQ5sPwmNlhgP5hCSX9qhwyTz3yJM4B7TyyPcAFDecl
9F7JV78RU2zVoyXUHK2hD2LV4TG/jbNgU8BfUODXY/BIq0HQUcgtCvlFjkPvQo8Lg5Ejnyk0GRzZ
0PxMhFWfEDZNNYmhKezZhhftbVe6VWO6Q2QvPSctL9kGOQXcB7NzNYp0jOL3DVh0BF+Hxc19PQv2
2kkILFjS9Y3z2pyMuiM1UbPhKr5WtWdoWc7WUZ7RQLlTtn0xgKhSXuPfqyDRb1kQblevT/pGojle
1qMYOAfY3a356T72OGT0lqAEHFCFc1iaQ5EE2U+1S52pGWirh8H/KG6oqN5YdFxNkqopYjdVWWvU
/oRGThkKcvCfenEwCq97wZOZiCdmkNQxcm8FGlmC86rXCGw+jldIxT6ifgoofB8Zdba1L+9X4oUM
swoNXCnqUvT6llA8ToSWtxjUjRPl38kduaaJy0J0lt2d6TplVuqCZDoc1Z36zAQUwua/j3zBWM2v
QVL6O99vGZbIdFRTpGmk6poqEiVOgqYDvuGDNtClUZCfN8F3PEivYGu+gn3198+r6F4SnNWivZoF
2t7IbMCToG7Ebdg8qy7nUHrDCXjB/9lSoTfKhmMJShWBCgNj+PloF8Az9qeIJIFkSizINqCGVyX4
2HJLyosWt8Hld2jkj+5hRBphtX7WFLtTIioZG+cDtN//0iFtooP9AAKNA9f0m5DK8eZcbvPSfCIV
tEBz7vd82GExr24qay3rWp+KDdzfcgiCZWfaHYtLEROML6AmVLOd4/rZHfyLJYUeS58WGRTiT2s9
u4DU/HaxQLQ5L0KQlgt7X7CJApsDtmcIHCowL4FuXHH25gnGB+Tm9VbUqnvDLYo2otAq3On/VNuq
93EzHkSoB9VgUsO0MxIEfKeesRp0Y0qH/d6QXqbslsw9g+V4QzPeuslWLnOJZ1MgcyBoQp10C4mh
aHZGYPDxyLaj5W5vdbCQYrIuul4BiiQpFzzcUH/5jghbA78BG0MHaSgpKwlhtbBpFzDqTZgYwrFd
2MvSMigI+9lMB3jHvdpkgZHJ8TMWqwUnsBeTiDmfAhFAjHaR3lDEGiccWu3zCKLw6MCS543LYAcD
xdhrvC2oEhdUT8kTwIzQwkyOa6TpRs/xpdZXGlbrODjqY1vVQ2uIyWJ6WiBoPBlvHmdG6XtB80OY
zAoQCY56FwvclZCIIEH8jNUvB+PwRr616dQfsxGOG34W9W6l7gRtsEiaDJbTEb33JRKOONuiVaMd
VhPTXNjMFk0cp245puvFytQjb2CwrT9w5yWX1LCtoDvWfa6330XjgalwAKf6nasV+/Ng/n2/t4cu
gokLUx716VqXGugKLs4Dzl3QjtnhjkNiXVeI//C8vDP8kL+0f47BzCuHC0DdOZYBUvcoc+9TZxeb
2WCS363Vu/Mmokf2VWM7ugVgSkGUjhzUKQMil9S7j3mYvcQVRvJ7gPCAlcWSLfpy+4XLspfO8nSz
NC9xFxGT6Vne/mqdV2GeqL7D2nfaCM18Ng+WveWx+FUfhVacCSX5k2l9wnppsgCcfXKRsqSFwSAC
kOmEtRKC38s8kQ0aUciR+RehA1zha6CBuRQ5BpTI2l9wxyWKPUbyDx1qqxsisLkj9Tby7gIbORU4
ciTbew2/q7NwAV9jvee5mLvjAvUY2qJPlCcBMeEgjKB05UQi3ETTM8G/O/y8OS20Ppkz1EXqYxK2
TtFBL0ccORno2y1lqcLuj5+j8jGeaSR+pFT5qVy8lAngPSScALNSj/7nN5a6TA2V820pGM2cROeG
mQcIr1jxZQR2imWmW4kRl711kP1Kc8s5Z8AdZUPkZ58brfCV3VXwMRV6rp9yD7vw1iXMvrAYhrLj
o7NMpiBNEC5dhIzQllKHCCppXuITlosFYCN34QmWD0RKlGOwtXfnFbcVFa6z/c2YCYGnN/gwVJdX
34V1KYn3UvwUTpSrBoNikveqUaarG6tDsQUBa3eOAf8pna1A4Xbf3OJgAFTB+IkR/4gALLacljl7
xj47qG2gV0zjllt0BWMzQMH3MeoS0EjLFemZYtzwVsiYyfc094V8MWfJyYAoSSQKhKhdmdaWmZxR
9CakIQk84X1aZWOnBTLP7vnGfuFRRqy7vOJKdxJhMCUibzt+VmWmVHh/oEWf3tk8SA7brh213ngT
xhCGtav6o+86MHRVGD2RnIP5HT956at2BeV7zSRn/DME9oZ92l20XtFDCeQZL+x77bW4TotY9hoz
MDgprzKuR3n2mlGG+DfJoLa0Mbsf0eUig7mzlKrwGP5s/Vb6ICWzXlbyOOWV4997OFZRcPZ7SoyH
3wZDefSj5R5l4qCte3VbDnFn3qSC9oTYxLPZ9Jouo/cMdgd/M+ALcUKJ29yroMeHOdNvs4HSafg0
C85AW/67x3gVNqKrVBRaNWGxua5CLnRV2sObOVhrWydLtYQyJcv25JCjwbQ+oLarUHZpjNvDMzao
ETDfCyEkR446mQZpIzsU0hYXwlBpJ45M2v/IK3bWXI9SDaNtYcTQDHFplPt7tGJls7zsjxI0gGDF
c5yc7IG8RURIEyGcVCT1hn3e+VDw3R+0jkXfvZa+xOmeLQoZaEl5Xmb2szmG4rlAZeU9E0I9sRHk
u1xUUA2u/06v2XDia4m8RuG6RoujmPyDAiKV8wB7jIydgpgRNyhiMOPf0eAwVfqjOVs5f3GtOfEA
BCNGwj06Il66Wm6dZ64YHC8HsE/Sn/2hstzLr42CtgaEA/xh60ZUaZtRsEx9B1FODFNa4vWPfdgv
ZDf2dgvtI8r7fNAzF9qqrycIY2TpQS+sknmVUdTRbB2U8KCjXfHbzieJ+qIzMt9TVkeVgpPCKnbg
eyY4XH92imTfsnYmdXTAyiO1OQ7imf1U2CYkkDnVArE9ZAKZSFGy4UFdPKzSNn99h3FfgD08Afhd
vtf+SbNRf68fqoXeb3mv4j/vNdNj5KUWd4c9ratOEHLfHR/K108uYvL5cycRxY9MxySEL4DAB99p
rnD8DZmHJ0J7231Tk0jRPqAbXSfmUb+ti8r/abjo41ussyAWOigZrukhVe1j7gIPSSB8Lgc8J4pf
z6lLmEB2N5JhjDzycTYjhZVfhgkAaIl0AQLkWfMmL9/vBMWxp7/M2wRRPOpzMn8bB8deAC4dhRzS
+csUhh/VGTt2a5lEX2D1SDdz5kujeJvfGRIP2zU7oclyRPrj6PA6ggY2CwxUs3VNl+QUMYelIoCz
Qv+Gh24spfbbLy7y16PtrjvIGu5YW9scPNvnijnjulODdx06Fa/+jes8DG4Eb38V8MiQ8NNhGGl5
3dmFrdFi8wHgFwXYG9pVoBBH9jFdxXTjBgwwWTSzhbJxPG1uHCDEkKSdVDHYAGta3vkHYS1PipR0
sW0A8E56CwO+2qUehnKV7dJjAArizE1WTPa1dqp6r7mMq1wJfUJEqnXLLxSFMuodgb50QEuIy0LQ
tc/N7hgEN7SJff1cZ/jRzZFuQ5GNbYcNKEpyYmQmXUPAChUbbQP6ggUO6Vo2/tuxU/+RNhXKjtOe
1hBgaxBtuNM48RuSihOVrmMM7jj6vITkc6fuJ9YgprazTSuY8XZDeP0zfnCp2OEDphTXXYUF28rl
Ty07iJPY3jbIKg+T8wSD83+5nprvYcGDMA3T1R+rQnsxgF3hYEaT4EQf0nt0uRevJ5yvqEflsO0z
SLjobs70DI0tCCmcpvbJ1rN0Lj7RP8vxCdG6Yz7QiTyq4n3kBN6Q3qJ7H05mwn5R4jGXgHSdGqF+
v17o8OXgbHYImRVXUZbG6wpvLS7BWzlA729RJ8z0igRvM7q9u28xwhjsfMsYy0IaViW1k1QUPvXe
8G9+kYFNrNriydsTBUJBLUZLwrUJYQLFci62uEJikytPVb0Hx+ZyVmvSVQ3kn5VBb8fWzUFq9sXV
IADrcv0eprrxCQ1WkalEOSnZN3x3IQZMoV1kSi6oUoQZpRDBSs1qad0hzXxhnu8L7TGEZEYAFntb
ljyj/6Co2VxtHFBDzH//bdNJU7o67agVtkKXtkeLNWe3YQe0pFM9avPg0mxdvI7Gfu235lMgCFa6
3jYV/g+9qrDUc5ujqdwMJ0wgaADkECJ2G/t1gTLLD3VCeDZwsyrxLooORPrnZnFLsQAuFQtK5kAw
iS3IxeUEkrCeQ0tTxVTmV61rho9sOna5ezPtYoVJATNJfKn8IrjnaOcPPEPEiolsKoI24EeE/L8u
dHQSn1l+LeiUAz6KyyirLDXl9/rnkcc3PBX8sHBxtPjfDz+2y+7tq+tmJ7HsxMRHB5pN/r8uRSMq
NgwGauw5CxBVZAr6dnaKrunh3un2RW8axFLOM/dJtd0YiCmDJZLxJjHLj3WJyhGWdOI7GpPMfd4j
PzgJywxg/qItDgQzGxMfQOIPUbMVHn8SpM3r2s5wVMa9pA8dJU/l2xPS3WpWXcLeA+kAUbv9iv5P
tPqdLx5xkvc/lFEFJqz71Z86zd5hVdqPd/N3PCd7N+8MdhNGhn2OmKU/q+NSQGkRAaL6r8+0JsSa
O1BuW3YqxP4ntaaKzzmCHx+GyGbhOTZkv6e+J57stHal2aBUNkqQuD1zhlV2R5k3+k0fPIhJ8Ms/
eXUAc7eNPfaA0FdMDArfKrNFBbDG/P0Ehz3bS6STqoK+pSec4MoQdv2kqvBjHTRHB4kGUBrqrzKh
X8rN2wR99RwY1JsgcdLxzbMkw/LiXO0ZKXLbzNSK2yNlXnKI2XzfzyaCyX8jIQW+SPLEMP03rWjq
wpCaQB+4AEcGCX5fR/8JUx76zvyF2d8MNrLz+hbNcjPWOoI4cuRNKF14gQh6UC2ugZmPMDiSdXCw
tW3kfOfzun6RpiZKddof+r24jKM2oQyo4O8mXQCG7UuttBYTxVIaV5G8L0SN6UsQX/LQeYXidFrS
J8aLhFUMBRK0cQSaROqqn3y7V6MOHGNyRMZltLzKblFrPrSyXYE3D8yocCgiSYYtPh2khvNN6PKF
ykimx7SxvuLOpevPsNGSiDhFDeH1S0cA9SRDq/lxqMVNkvHuQI8OQv7YHvkBG7YBcR1zeBbtSq1n
jceml/dujmT2ZXCxr2qm69tRvogubqYOFa4gZVymtP7/ds7CgW5NZ3qY7ah2lnO4sem+Da1pqYSS
dgCUjS70YAO52UdfAxkJCDEAQJFMG5Qt0uN3Fj/1k4VS7nxWPoqW3KDTzhZEDA6wjsESqtYHsesQ
SLQ6zzUQia0fxgH7/SBj4k2M+eUYwmCfKJDhTyW2mCVFKumrwq0WGP0OOmBwHLf77ZZvBOwJuaTn
Z4VkdY0tp+1r0R41+QwIYkntuMPkqWwPnltNu4Iw7GAUt5k2z+fLCxpgevE8TGEdrG646+c8y8Rf
pSY8I/H7VVDqSJ3kvay8FhPWQGn4BEUe/ADSQMjqx3jV1Ra853EE7ItP0ECIJdUeW9OlZHoCtKdO
/8ezKlMS6Kf9DLYC9Iolhkpp8EnlV/veBaNHBwrHE8ycujSwcumfW0+tojGCo0e6xf4n250OpIz7
A5Dz2j7jrQT8y9X+QA0fHWJX7tS3F8qSHgvNOqnz37A2DE9zVG0f2XwXt/lzK0hNq5maXJ0gy9Pf
6sWHTSK8Ff7VyxFQ4/t59uOt7WXJU6WtB8JHsWHl+qCG0tNbFsk94+Aa1ndeviYxdai/V4mnyB/j
+yXoT88BxCVHE+vG0flhFaq6wioIz5qy3B5F0OMismwP65RljRUfofD1eZSi8L7zaPjlsk5iwi4x
4vQb3qod8CD7KjI2o6E2o2tdEXeRL2A3QtXwpOv3O2ecfhwL57D7G2jcYZTTSRlpkLKxJfOtWQy/
vrFKVc3M43Nr4hR6p6Q61DJEUPke8AdWPnNPHb7yCAvIiBKjORBAaWHcM2kMPH0f07YsD0+ST0m3
CYYxbf3XJvXjy6zi3ldd7bdnomYYPlHtXWVyilZslJ3D/+Pu/c+ErIGn+OLWznuGeMOgHJEZFNv1
so2NbwdPfqPUl1h1AJkIw3X5HaugFQiL6jStNRC8XVrdaSYFJhEpedTwQoT6dcYeAqft14eu0pwm
nrFmZi3q233QDpbBYUUfj8RNk7EqxvFzokZ5iNbf+hlSkJqTzu58ghUctlzdfcoAeJcUokaiopAw
0+Vk+wfsot35/RVgvTRB3kwA8wLTGcO7C2URSyChpKIbGWPp+ABTT02hGWYm5r4MooITcbtQKx+x
S304bO1trCkY+51liRquodkQmh5vyOuP8gYfyILZjVrCZgMySbnM+bR1bJpZpz1FbAApxkyzlD2d
ogyyDnWyJjj992DSsOkSjxv7rbnQIDLSWzkY2YmHdi6gxpsa0sQo5DERo+0b09RcK5n13tYtBiuS
NgCYChso9nyTjTc4E/8LcMRey4WRZlbw0DeNx9SDVrA4JSvKlStw13dxlYU4kuurK1fjNRVbPAIV
se6WwocaJcuSAACBMr4IYz/ZitKLIAVo2PJqsWIojD5RkP/axHAqbUI/h5iQCt0DcbSGnNJo3S2p
4xoUdhBuHBCx57MzYqTNNatnnmIXOQ9msfRvmHO2iH6AytE9fNmfKNi/5kKDE6S62fAQXnYldZYX
rvKXUafqlkngjf31wKnXyl9kkUaqZrmBRTAX/cBteN1xAF7vUMuMBylWccNI4jIDw1FtK71JuB0k
lQjBRqmbC2Y3iyzjITK0tQOhERC/nyhhbi3oG34TefiGuEiVvrhl9r9dDOTpv9PTucSD+61AaDZg
Q3l5aTxQo6UnbkPDJlMyPTljgaWhLB3ytTItaoip5pZfooseNjQ5OSKVZnvL0qoIoBjiHgPPBSzD
AM5ixuhH3ZYpcmo0eby4eHgV6akCsNisHL10YNp5tjemlx25SxOJSgCxY/EbVt/rM7LLStyYHqMU
EnuqQ888pBYccmX70Ef5gEPK4IE9nKhrgx9eYFK7sZIA21N1SdDZjiS8GPVz8qAm4nG0I5kgCw9X
el0SdHc/t827zwSZsHP8/tHpxieI0dB6hCchbqIfliHtROBkYYUEGCEFuI50gRBEHsvcZViC7nBG
xeuiHFlrY5Wjb3cyhuf9DmRPYlE2R7KrYKLou7NF+H/glk1Rr3SlidtNvneGcnwvWWAbR2Oyokcj
OD4y6OpDAeCCl6YQL8lfhyQYHDm62yu/7oFcwIXmUORmmFgy/bNUeMLV4poWSSdvKQc9geYs1hQg
kbzkVcizOAgb/FZHxSMgC1ika8zWHK39lrRDQygYdh23IC+WIleb+M9HrPWezfYvRUlCZijhN+jx
UkIAPSwiE3CPHECffzKOd9sHc9GGmdtzBskmc0GHSudgubnkWpaPX/+L4qqS97LYTExs4AzKq5E4
bKh8LKgpXOFpeA9OisBQ6Tjl5UPNBlVkIGDOCKsJcZWqMmLQlc32UliiOvXvg/z44MlrPapboltN
bM2jatgcbbaO8lLXgj7WvatKpiojw/U8k+txk6w+G1w/x1Zjw95oc+4jf/qBmpYEj2QOjw+a/CIm
TZ7h+EBs4NxgNjIl3nSUZTlVpXsKaLQJ691X/ILvevu3zOjL0Kmqj7hOlDz6BXCruR492et+00rL
KfUKOmcUb9avP13cCykYxcdJFFP2UmopZev2AjmHkEV4Y6NGxGM0XGlM4uLxyNDMduJw3CLzzqDL
2G+kwecPCjJXmbeLiNqUMiHdTIDwTpIMN3BlJS5lV31F25OzyeUQEmX9BdbdC+eH9q+adphb5lnV
jHjXpmKYQqhzlNKQGq6mojcTzqI1SpDut25spwlZIzNyb+2yd5mWupqdEczFWOuD9310aa06iPt/
du8LP+rhUHOIycfv76yroOc8mQJ1n++Pk3BEvbRjDgf+vsMXj9iBqDsRXtNTeOXBuGCK2/Pol3Jo
lVgfrKEzlxNJK61M3rLe7AgTwC9NojVMMn53H1+7MXEe6OvUeSd7z3L2lq6PedmDrCz+vrds02Aa
SZRiZwFoKW49Cd8ylMNvw5g7qxXCdRA7m3kFTb4IVFXmfMG+bqiZQr2z9Pv0456OPoZ7YlawU7yE
/LPgxdKSxORbqoU/lm696FuWKSTDiWFpDhqv9pbsmhxtueK1fsM9vOji5OvtXpnC7HrcgD1p/46D
3z8mgUI4KSghjE6+1NcLJItfBjdupnRaSRUSJIWxpdTThAbRxX7Xbh7CA7XBDchcSGgd/JEC2sSs
/wD8UeDCMLSk+DanH2NH2Rk+DU8Tp328+TKp4/0KfpC+YFPlzvci5DQIE8bcPMWvLfE2S+t1S4Zz
C1vXfbkFd0R9aUiyYkKPA/b1HwDKiEEUqrGxhy0ox6ONHRLOLaAJEqSTZJYar7Nn/yN781iDCTSU
ZzDtSdbaVRHHwI4G7MTkT9B2C2DRqeFJywAWZL/Vz+UqU9Raa+Ol4PWZACUsI5ecWM6jzxWh5Azj
MFNnBEXyOMZJHu1k3UtyQmFHUrmfiVe4s/xEX41UpptlEgQ232cWGWs3SYwmRv6F6gmrh2XiYc89
RmvqkMa/pYKWPlhcyFxhsHPFxk0+/N5q5KsphZcVetiA1dt6doGLRhvG1MfHq3FGoyOThp3fLLzb
jG29XMGyGW54dwm3V3u+OVZpnZv+so8umzBcIy3h/GMiR5YbBwhQN+Ozr01Un0qswoKmmoal4PiL
kzTIpxEOIMinizoJWH51kLC284+1m/vEqzWz6V95M3xsU0NPPxITHVl250vmhtishC4im16hT13W
hY3M0dWH7VrJ0ZWMxr4sDdNv4TZFluShhSEdV4GJUiU55cYBPvd2H8KsHzHf5/syvI1dFDyUCIXf
+sZEpJnmFf2GKtYk8owIYN+02Q03LTPJJjCB9NUAjq7v/qxKyMyPmp5/xd9XpkaSrLSKvRA93wqg
hNjE6LAjJyXcJpbmU9YrqP2XM8bHX75DY7gOZILxjWFy4jZiSohad2GdC60VRzflynF+W18cThI7
ZsmD070j14xjlXOVtfrL6pN6J6YOpiE2za/WBsyFrDgNt0xDoWrd0RAt6y7kHvFLhSqQS+ifk0wI
PV4999+DwhXYFybls1v9ZLZ6K2qTjk8/hlYDg9W7oQ+nx9SBXDakKtHqgLWKZZhNE1P4bY+YRb4m
4xbYH+ZR/5SFNPl0D039Qk4JLFuo5JYfIdBtMRd5M8Xek/nhJAwaUqlsNLwz92lMiY5mkpt2HWFg
EHgm7B2fRHdSf6CDU6jXbqrjoxMoMh59Jo+Us/SvEJiiQ3eH6HfTVxODL+A3uh0ziKWZfmRrpOb9
rn+/cdTIHnJU36L+JooIv++scd/yZPjL21KtIivuKjQ8B2XdR6X6g+L/v8wRDO6/OIqbI+ZunIYM
8mfN1Ah3WLm7DuLrKT6cxK137jbBbqbrlraZ6jF4wiam5cvI/P/CrshGV+cfADCikFR8SI3fPzdp
RVDEGY3CHhIgMVweZkoTslV5HxBNnQjL7V+Rpx724bh/atTIPTwI0JZyJ/mYXlwIdBdTA96pO5KA
xIOevyrt4sk12LvoR+XYY9vgkDR/ayr+F5/uzeMOx5TdHjxe3Xc9A0nXAJhG9NG69mkxbmlKZ952
yY95SSiDd4+b9Q9RpELScZH8nHlGvu0k2RNO6fAsa9zGnjfZlMTcaIppQwJe/4Eh0MBS9ggzZDvF
RzqUb7QxkCO3oXtSiskwVOQZYTy7Yd5VGiOBUc+drrzpDPwCkFG0P09269qgZWSf3fNemp3cb5rC
Txa0wHyO733iDY+jTx8t1XWGrziiiXWA2ESs03C7mkMf8ob5n8crhVyQiCRTtUL5hUc2Fuzpl9uN
WEYwWnpFg9TYScM0deKpxp/yVcOb3k4Hwc8GMyC9hh+eDql5qMmaSpdEmeBFbkcOrEU+sp2rChV/
fboGVqnu3XqK3n+MxB7hCqSJroAP9hN/RTXdg1yITe3KC802eKRzwFQnOvT0CPmLJcIthhSEol8T
fl/N2AbMafrUY26gvp21IaGa33xAr9O9sUW4zOJ76cNSb1p1u80JQveYb/TsfE45Jh0l1i9STQoj
OBFZqGxirOa99Z5no97FjOv63AWtuUxyGBiplFQw/Nlg2rnNivFbltSZ5FG9emNGRXOKv7b08xnS
ccPZLOBF6XH26SRmV060bhegLyGgoJaq9ebXRUrFkIX3G2qOmdq5+LmxQ30g4LNuzOmgEGDjAH+B
HYLQEHebyUQoiNFlB5/TLSd+LbHBAp9aMjViPAtC8TtiiIBt+5r/mpP6GzizSIlVjw06gy+BZDtI
TUDHDI+eMfbvBepUIhtQH8EpGZJgAvZm0x/4cwtiR7ucEucw1Mz+MGqGXPIBPQdKrMoxvo0Nkv9m
/JhdGEq7BoIp+TFICqIJd7QIkqvaFzWZX/D0BEeOKh2waLlMszPEXxDm4R8BtdLElRNeUE1YTBEg
mTs5LYezdyaWLvqXiQXhGIRFxRwM45GZqBOoYefIbBcGGw0A1oxsbhcCC7GjO2khhYFoWl5un+4N
ozlT1Po7DSxTXvDRus3pDlLFdycUmwXnN2RGcdDVBVDCIuK81531f64JvvUBSrsqDe2C1Q7TJoyR
a+H5y+Mf50FrQ4MyY7Kbpnp70v9zyioxez7bv3f5i1pZl9YTvLHj7uhQbOcuSmUpB0idvQpNFoQe
v3WiQSB9HYbD7pMgB82+8rcd94OcZWKm3M7CW0JEXNZ4Aqv4ghmzbEodpW6OMMbWLMkBw8oBCVnd
JyHyRVPJawLqVWXW8cyPuThCK0Wm7IjayL7nDjHVUqLfGdRBcZy/TQsC4VMXk/4Mbk4+DEqUJpJ6
vleMjfvxdQfwirLXt32aCi5/UJS/ciOC0a/hhL5bPz7BYQQtT+cbfKtLgVNG2KLfEeqm30ZKqJeS
S5BGLGvqgnqp0FG7KjNpQZM8llVw5kNTnwwFGvwnbMFL8tjDApAT4qSTL7nkUBERI8qzk8/b6OhE
vogsXwO2S9vgohplewXcqNFTrPaTi+lWKUfzFNl+LKco4iY/R9twEOL4HxQ+upMMaEgsvlBA1g0W
trSRZ19uhoWfgp2B0R3OTSwn0UvlAe4BMdOnSIb9GxXLOSYbDDURtwPa2PmUvg4wFxbTHdf4/100
9qwAhhEmEfPwxjzCdvTLhxUt0RFMVzChqQ7nLQb1XiuSEPzbLNaNJqankPPaw0RTukwBj4rw5fS7
YcsMOc3u7zI5HS/wNC6o2O3uePVcp/WNzBdxF2+EzJ1csDS+1XoaDRg/PQWwNnFeScNVnn6uXgU3
6BujgMrstgmyrhYjl3ly/wu1E/hsrauzyVYViUFfj0H1Bus9ZuWA89F9hczxuNIe7WeyVxnwq3u9
RYKj4DhPv8uCysFKxQHhjQt8+RyuS0pG6nHMhZiXv5dzvimYIShJwEP/GWojxToPJ3veVujIddhP
EvFkmkBTBLlM3lj9a/INDQ4Hzgy8LvglOqaIakLp5g9QA44S6T5+aiZc51+QbFLNjR9WpkSG/0rQ
eKyAiPHyGVkq3jfs2XhjgnIug8UGY4ECCej3CRQL8KqCBeWFHEL53dqgYM3tHF2tJ6oR7l++2GCy
MuYxB7B24PVl5t/rD2RzHZnYyPHAMp1WJlPfArCBTgL3ffdNLhZinnFSoFnEsDDvyYXBvDDr0Qjs
3XaEW4YlBHlksa75F8u6zBMqoGNkNeUJb6lr0xpXcL2ReB++hhHtkQ4unirbTJjaM3LYtYy3noaF
zpztn3PZ6DRYr5hvGXL4h7xVOYY4w2diIGUqWdzxqw2ObA8unbd4zt3TfgE88mZNpE1PrXjva+XK
yhz4RujApYQEwG5O074yQpqPRRr3Q2YdbToUyx0xz6w0DgHU+yx3EMe7+pdssB96/HwgEr3jhEwm
bNc8C0qCOBTTzVqQH+qBrd61tyjST6mP8DEET2WrR3zNWAKqgGpjrgaQAiYlTX83rD1MrMHwXXWI
mgckZiMa07caoktjzBiN68xM3t1xKTTx1L0JuRR8kN/uvEyz/8HPz/HheeUR9jGUuvvkiLGNIhX+
GFXlSPG/0LmJWPG5ENLUhSqHtc7F1tTp4iWxG1TNGGN7Yf0H6QJEiFMfgBC4zOJy2h2bj+BXD9/p
A1q16uJY73HHhdu6U5mIQm1ZlfP66GAlGQOo/SFPqK/a/QsSE8YZ2VEZvXbB0OvlwMiHvbp58o0/
t+LNwQO9hHrLcTlYU2RrZAtlyBizYTNjIXovUbWnqqm+ZZVB6ZH1I9sNc9QoWe646qOandbxrQIT
jQ7u5IMtKZYtsjlb6qyLh0PKEzfXQa0DwuDD0v3CBFqEwMIia69I9Gn3uKAMfthhRfEH2FqjYv2u
oW8/mrOLEyCtkt0q5Y8fHPuYkRavuKF1/nT8x3pR2zZpZILOzVk8nXdkEXRLV1Mbzycr0H3zN3KM
tizuuwEKvM80J6XgnRTiS1o5xu9/7bWJUFhmkDhzhkX1xsp9RAZTBKlDdE8fI4bIwAvgpLkYM6vo
HDH7cOoXGwEHilbqoZbn9qBVBV+sZRQKlmkxL4yW2iQr58bnjNp/y65eIHJjazaiEFJKhFSOWdnk
RyKsCooeRN/eJ2ddY9ZJTESlYcuRTcOHhEzEifAnYid2jOt5KV037R3uUgK5bPb3LczgvRvBX1D8
q84yqShmK5qZ/z7xshYtzmqda5dEmVaxZBB3U0vjxLuujF2PbbTdPmpFxVis0SkD8BO8OZyrAzYm
mAjoHOUl2lx4ZccQ7+86sn8MdWK4WS/vcHf3Cmsw1hukq47saCXS7NagIp6FBIsmznxBjfng08kh
d4i0bi3eSjMu62C7vCdmSNGzu4PonOetLNuX0Wcsrngeb0/r36HwVwM9oH0eViaZ7MMBwDuw744T
munwoditNH54jKkV9WOI76nnCVVdqnMZAl48+aRA5IInLv8x3ajNrwe0DMVrYacXF0MNzQOqoU71
8NipQlG4O2/E4eQHHP8AIyAAEdtpcuP5xsVNGFmUu6cWGX2vDdZ7ofDeFwHyZvXKLSEfiypwwNTw
2yhXtTXUH6GkaRmuicJ2sbCeIfno0xSFNgRQYaSLDbEDtkFXJT7iXyQhTCtRpItGWv2Y315GPaUP
T3J+DuKYM8bH7qINLG5+rrC4keDFmUC3eQIu+GhZQLX3lTWsSSvZZxel4l+UMUNemNKwElLEjoXS
xOMyPsYiSD3gYe591MjvVe7adPTwaby+Mo5+j5q1gn6/oxVBN3Rqx/iEdx8eirVdEd3iYXdCX0g7
Ft7pdox24olTX6a5fjSseFIPBk5RMxVWuuRtPILtjvApZB48dVHdwDa5gBwoT860cXhYkFuUC6Bj
KhrxGkgyNLJsir9NWFSQKepbtwUyEwoPCM0M+ZmSus+Ebl6pbRYUfj5jjzi0JdFUjF2DyJ8vvfVq
xvhPzDbTqxxvIdL5y7vegcc4dK/oLB6GOLJsJGii/tADq0mv2F72KfHoLBRjMttIN4km1nFHCHGp
CS6bS26XBBwfjcye8yGDbwKaHtxthYH9AzlX9icqDac8mcY17NtCc/bvxT6D7IdP3Wuu/bZ8jS+G
7kxk2xjWUqlkuIl+puSaD+xhKyuFdV0X1RKvlNHj7oQTah2ZhFQZDmygdEeTS0HmnWCa0WOQGpZ7
0YEQSYHExU1aeiQ+0/qBZJ0AaGTuWGKRBKGD1Whzax3Spw/h8fY0PYAgSclMDyiLDOG7GhW1lN/R
4A21zHHwAel7Xv2e08f6sUnY3OGPYP3urqR914uungCXoFarCBsRjv2S/57Pp1XF5UboCnUBPyAu
ns2h1chyZ9kO9lSf6DPMP+8eoV2GKz9v1WSiXJ5KbHVHlTwDD/Ey09ivXtTQGcgOwPlF0LA+jZvK
gpCGJ6PIOUYdr9BIJjPkgy941teDHCVSYXv/u7vrs7OKmA8ydp68TidIqlv8cQ1IzAP4MjLWZ6Y/
wP/exl0IUCYB5US1RNbozg9yae6bHoH4fiQL00+SYBeK4LdMZ1gnKoPVrtd17i4OAwu1C323wDIM
fTidNdG/yUs7Yqb8FHjp9eWs1sG2s/Kkb2yhj1wK3q+Rusd3byv3LlwqPESwgYZEMd/zI6XpTpy6
rP8ewBie2DtYbHrwJ7jC0JVImegKF2UVcsrsdoQz773eKVHOuGn+T2GQ8a/GiIUlMPfB5pID3v9+
EV1WKxMtuqUxd50vYFXmyVWuqIvUB4pbsZrkv9LizXJNL5qvhcL5oBpoV3FuRk/A3QLAYQxxYIgq
3gJxLfS52GmuCmKH0TfOp+BwEZGA6Le5C1LSRKGPlEL9BVxvLMTfyjhsjm2YHvBN7/FrYw//NV7g
IcDldwMi1OiMz1pX8SjFeCsdDnbWLGRHiMLfQL5hX7ESot0oj9gUbYMMUdowzP0+2gSEQeg5KKzh
xq2Tuek5/61nC2SotuVH8/XT9duMmD7HJaLvH1x8i6HLQ81l1u9Mj8F7OmpLern+q3CNmKpTyWNF
a5c7RCw8Oanb7TTNOnqqLCPiR9HKQKg0z0hkB3bHqN+kUnoEIO7Rt6lGG++53lydIXAUqnWl8NAA
VDIqyErXedjPfqJeE7+quWqS2qiBbWvgyKy9aFJuFUzXh7MoW3RJNEDUEInjOCVaZ01j/b6m/Lj+
vLEshAuHWhSk19hvX+g1eSfqDOZDmKFBBGRFJIixuy3QqSNnUSm7a/X2gmy6cwKsHAKUbHTM3nQp
KsWbiOEDC9YrEZBSUtpxp2sDMG4nNQAm0t6U8JoWMGwzR7FmKS1o1bNxrQ2OUG0iBGgMZ5llAlPB
Vg11BH+X3cR0cHsYJUwzmhCBi4KYHhMVy/wTJb8DSfr6vNbpWsWL99tpk7Mg7nODR5Yz5T0XqcQk
hc3NeJxhOZ8WDTFlsM4wsEsJnz5TCsAaZKIr9kV38DdaeTbqmfUHRblk8fqntm+GoEbYea+Nrnqw
acZ6uaVA6kOc+e5iKe1hwxN/fHdoVBkDu8DBBjZEuPfCXdkDk1VkB8Qq6HoWIDU8hqoSxKaV4xsA
GEggY3n4zzc0pWR95wqo8uVmknmi4zIQnVEvrfKMoewq+Qo071I7kvrJuUsDANKXBD0BZRHMC5/O
GtlXdL20ggGp6Z8hUssbPt/lMj73kIkFab/1MhoRxwTCD23bjRX97taYZlsFCBYDI6oD01yADBVC
v3mzQn3q66wDvGw7XuIc86ruxamPLcAkWA/fyik0uWD+iCF+x5hCtJCs4zSlLhzX4SjamxGDza9z
YJGX1obyZBk44CH8AFamLpsyU+IENy9n7DHk3lUw8ItU9LAU/w6+iYpNPMNH3qAWm9IksjItxYlS
5eQe2Ac38g1uOOpMn7/QdUdkT/x5yu5VieDLPdfi1e5PsKm82PrK9joyz96kA2AlUWBLtgw/gNnE
ZQhAR4mRp7xbqj+844tJG5XN+j4YE+acJNrGI3ZNaVi5YAgrr1L8atu52ThqSt3MYXWlbsyDp9G6
rjAZkb58LhZnifBna8yihqUMQQ5eV3yCaPvDg6LN15XoXzKXpdkxTvddjVwlay/qQSF9Cc2XnSPC
q65qL2aE392ktGfZObWemueMXcADj4YfnYYKHhIq0uWRBVMTvdCbICj2PzoRDzuIQGQrDyiyylDE
DI28bUYpLCc48SwiZS8cdEXfWmxjOxP5jjesgyewTvjSC4+JflKa0+8W3CYAJImnzTdGGg0z9F08
AOGEss21z4Hts91qrSz0RDU2vwoCnOMvLNnO+VMKNgHsY09Jn4qq4yMuJ2NUL5glu5S4oI/vwDTm
66WElCT+5lFon2tgbqGkILBnm5KYisv/Giz39tHLT8UEPldGvA7rIBK04PU+R8OtAbvlUjSe5ESg
wibZOmSDYXJsFpgjiGM6/ZsryI4Jm5pM2+RZNJlK4FYjNxCxHtMTK9CrO27rjaedcIvd9WHSnSwU
dwJO6+t3hZbMOWGXxqljmOcJVV9aHaKR4jKkDoJOVBzf5/ccKItTGTx9B/KWugpA5eA0FStonJ8F
30eZ2/VZByiDyCRCNPPWX3J2XSEyW/1NLt5CeqLI38BtDqOEW4R7SKWPcIzuwuq5y7G1Ix3XIVZS
LjdMP3Hcz6ms4i/vxHND4/VVvZublYyYtKu3YzrllTIu1kx4bGzBcSNPGv0Gqh7nzzuJ+c1xGyeR
JVFVy+97aiwYskE0k3VdwDgUxweEq0fMTNIP2eeaObZ1oXDIxlwo9H8JFqhbACdtVnc2Fz+UA/T0
uiwUCbG51ophClWEsWbXaABGy6CIMqsdug/4hXMqoJ8biiDhTkd9LCiIt09FNWmKuL9kNW7Lk1DU
kL4Xu7ksjGYcaH676fjtW5hWN+3MUA4iDnMaIfi9TVFzybzGPRjFBaxpaV9OVMw1N5JVwIKEGzrR
S9ekgjtBPYDiUEnV0A0h0wpA2EcJ1WdVGM1lNdrNsa+Ek1mfNKjqMatquim6dhZ+WCTyr/iB5dgR
Dl7PYn0GNtFehYHeFBIUcM6h0Lf27PTHPoccNxCqylV1jHxBDN20YfcjnrDqNedB5HvdH7VYe60Q
48liSv5gUCvQdwOivs8RASKExFTRMDbFsxCdpfxhe7jbdunQ7Mk+veOwXOXUwKwHbmRMcSOGbsql
HS6atZAY+olM2z35v97Fvx3nLW+Q2WRb9t+FgV9IbdvxMYW1lSZnrTKYe+e73yKPkuOfSErLkVo8
Cc8jEh+Ek+uxJky2h2mYLjWNeqE1myrs20Om880rfp34HCvWEULsktRuIRU/YSQNCP5QKqoW3pop
nkb5IsyAhUVz6WsqZ8GlrDa+5ASkuUog4s8umeoVkSTTXSWXkMd2r7TSyjcW8DtSobIgDLlDiI9x
Hh8T9SsDTgVa2mSRGDTws1DETKpfSqz2oyPpsHAZneA5ZdQReYi/0pIlFfo5XXIajDkPR4RmKRXN
LSWoNeP9uwyTsXJVbZlqorx/wQd8gmZ4JtcWgCWqKFGdvcXeke/G9G3itNpYoqD/1Vb/U1VM768l
HIwuSj5Locp1QDLt0EMqsdZPYbMyVqN/XKvHSD36B6s3yqnpjzVruRCIjY5FH7l9qjQHCV4AEgi9
ADraWmUr8su60fsrORkyIc4ae0QD5Pg8C0tx5dQPIryaIYl6TicNNRX5vFD0BGcdamOVg3lz2wUX
aTI0R+8iGKYVY1WmycMU6c/HqSjn9yNQ7ikTXMT03FZuVXOqWPWxwbrLp9p/PSTXbWK/pCrzNwne
5flQh7m2PM987/lLEYTYVW8Hnqog+Qs9ElPOdCGHlgCHJivrwOsgR989T3uHGd/P7gJ8da2m0N+V
MzGbiwy8IASBKJ43k4OHkhZNysDQH8bZNwMIy62PT1tmz09/jqNjkaPCK7a0XbNsS5fRIVsnBMMR
yC7jucK4BryBYR8DU/djcVqUVkxsSohGUqX97f7Eja+Z08Gwd0u3crgRXHoE5HrkoxGTMwYxUtq4
6gMTzOd5FEPqsVuPTROp5A9lBWE6fC5XnPmaF68verJCO56OmhNKe16f3tineSNa1GpdNyZFU0ZR
XWMy8TXWp5dmzwFZY3qWLdTlPa/l7C/1KSOGuwqNr/IMqUCo+nLQOaGiQt0gIIwTqDTnJAE6RoHY
sBOcnTayN0a95tLCG1V9x9H/NTcI0T5f0d3GIxcvSaZO1drlx7d5y6xrn076pO9M3i6C9cb/kicw
lR694kyJ7aTNxlRnf5+Ksp+4pxNVBVCoN6OPsYsd2OrdmfuVgWwLL76dBGMKdxV3YR8ziH/hLrmm
0UxtS6eP1c5aJ3csGekwy9ncVHc6a2H19MdfsIw5KxTYTcTXB/Q/mnJwN7xoDwUBx9ZXabHlGjoN
WERyCDUGSottxaFBwmVHkRzKeecqQY026xsvIFfXvadeOIIKSm3bfec/mFcpVOydMnZfye23y3iM
Z5rjkMVRo5W7+Ws//P1vNU+OEFxqqSuyTKjDi3wl5H0w950nQg8Dyr7yUUBQOn7bB6b8iVxAlM6K
N9TNSbLCsmKUbQ7vw+XOH7+9MV7IbTHpdILR3m3V0Wh99biBYY2Ecoi0R4L9UXzXKKetMBvs6Ug1
onxwC+28a7rWKRN0eGxH9MB58dHVHTppnLAyypPbt3bcblSESl6APT/fFd10JZV62W7WrmuV+9bb
2b64uJwHOeHKyeJEoD6+1e6RqGLJZ5PmKF/S+Ou8/HycDf4pV9CTMpF1o++BKHhFLqAn2GQrU5GM
NqS+mMQlb46CU7LEQUc7e1f6GHhAWQTRvaRIW0Ux5/UIp9PkUfofRg7JqteBEEFHoB3/tuqt4iKO
nDFoOQ+xm4seVGCXDXatBohuHZXVj1JK4WIfyK/AoRFCWRe2fA7ddFgSP/H8s67y11y41zF5YrvN
6K8qgwCUlVyEqPR/UhyPgaaDrmlzizco9nqcLYbGPP2HeR8oPFGSfHOTDhP93/B5DZV91odxISli
aaSX3+fnnprd1KaZaWmoUrjDXtDvH/RsgPhR3i9x9Mu/3iVhXLEVfyZDz6FrDv04XRGNYPxi34He
H7NnqTPtBCUx0/IEtPRl25wEqzQkZVIuI03egORQHkC0M3wiRwgVQQv/lKNLjDGZr3p8/9cUxEoF
oJM1cEGWvrvX9VJW6S6DSC8IQCdW2zlvhkguxo6MxTCYVc7ijbjgrc31kovUlbwYc9T73eR5/QU6
/HxatYiehut+GVywdYpXNQPK8i6Wju9ECjhWJhSnpKH+9VCVSE99oqOc1pXhEaxjmXvPfpINWKa5
WyvI8kpIjYIlC5oXO1KH8fGHd2Y2DJi8gQNVmidpLbCUS7QH9Jd2UpZIGE2GHntCHQsjG8Dh2ggy
V3colQoagQK0BjSMzJ8lPW0TkE5DZObjcQ5QgWsFYqSPfL71F3zAqFZLMa8Tz24+6tBXK0OeBuRN
HVo1YaH6xYluOZqgoh1TdMR+O2QrVIwV87ak1dTVFDr35kt0HzrL2u0lcFJ1Z1YhXMAKrU33XR44
rND38VQJU13r91nPDPtwZUUnHOhFKJn3g1NbaRm9fkvoRFelzH9gt+slnxutdlCg4bmbUpQn4292
mQ4841kP9755mGVKvqspmx0XoAcvfxbuWEoWiREqmVn7+tuvWPu7UHu1gw7E6EDs31Zo7VrXz/4l
foc+36QA7HRRYFv8VVsJ8FMbC3sy3uMPQuQH6L1CSMNzW7/WKt6Cul2WPFvGfOuqrJrVvXiHjpxP
K0QSDHBb2X6kIJpxKrmbdD9VUpcs0ydTYx16VaKBW9kvzNgIlglgTUt88EO/wfTJHVWnrI18McE1
NCWY9HoPXXC99vhBD0HjRQ5BdWfrBBT+vD8Md7MUFoFZRjdK3kwBC3dsavq60H5aL7mMl2Ia0TEs
wPWko/W0A5dKHHDLILLbTxTlOBfQqmwLA170UCr0N+2p2kegdNiYFmA7Nv+gNvO9QCELqQCEeLY0
FrrXWlPiWHzSL6T133pJEsZcC+uAUV2KEkwonVSXt/TsuVIzdj54ffv9q2MEO48hUHfuXq3LI0+A
M8IXS9UqcrpCvQadGsOAfeSTIefVUnRx7O5S+3WWUrzB17u6McIFtj671W6vtuBJyHUPyY0+JbR3
dBn1BEvLsoH08+poahoVQjRGjft7+Yenam0qUo1Dt75HgN6QUSOiGRq2mgI9dOMQM9wh/E8JS2r4
eAi9VjFPCj2/RDqNhoCI75ji9H6uweAh4wkG/Mz1lTwc/LA2+uuuNf8fmZJOZimKt9X+O6k1OJ4l
pQHyJy4K4eMpxHFmmi4PUQAHuoXqKCee12xKAt7O+P3X3uvIppodHDPn0A6JuQT1USoUmSgSzFOL
1n6WkuIeQb0SB4Z7hSVKd+ly1iB5l9cwVIK6pBQYXYRe1xHPoewjbSkWqWMqac3xC2WR8uxBo7zL
MihGvgSex7qP6s9ANu0a0czGUubRQzZrBGAivCVCS3PfWu6iFv9EM5FKTEIzdzemF24RmOjnjcTs
EIzEpPoThtYaklW3D2lXjqqsb1JUUV+UqNlsdFmK1ByR+sRGC4Wb+hwOGAC16YS/kUtane1DscEq
Ep1x9gW5DiamyboAHgal3WQ2NK+L1iKxdAvZZLmB0QFxENx+hxzm5Dlx9ET8SdzuB+HsQatE4O3h
/8t3sgCIfvCpPvcsl/hAV2MEpkGuOvB8eAbwtAJmlzt1BjD+xwhwegKilR4yhWRnpovKWQIZtDGY
LwSVL671WZARGfy9ZtKgzOTrv7KvNMB/j0FI2/tQDemd7QWfSRfG1vQmSa90PErXjnGIwzI53k3K
ckhmyKuBJzeSe0TEVR+nateFJihXnjuXkgNeRvjVcjQ/V8pkC4fBE/TMZO0Hag9EOcvwYERhbKNE
I+uo8xmBn86TWITgSnGnZVaXnyMgHOe9DDS4lL3cTNDQtuT/0x+LROGxJOZiNOV50lyQHqneDeQA
Bi5Su8GwNHI/u6JVIebrtAyeTLDB4PzVC62aO0YKAVhHiAFejsDpuCipFQT6p2C56AJqvPrZlY97
nri0n3y9RWjISe/bop1Es9igjIHkeCq/GI2GiBRGx4He8nOy0piNtzIBNqs/ptQMpzGI3meO6jUi
OFR5g5pnNuKEjXfrFAq1ipPE/aGSfVQ8v3JrMCAkd1gN/1pCzK21ht3ZVAZ0ZgiV/CiwUBSnoxiU
42rIfOlBbp48GVoOEDXDDf+x/GzVepULOJvg9F70uW6IcMb4sLnY59AC4erx2ZgkFUQvodHrCFP1
YvHykzMufAIdS+b8X7R6G2QA+EEEZF6xdnzSZWBzKAjODAVbdrZVJpEWjnk8c/W+zJKY4K/7nlzn
cZ34TB3JUOfgZABZoVVXPhCcT1XHlgrQaBnBvr0qjIqQH7olc60kp/x52rM853zipRnXzve58Pa1
mUaYO6fMRibLP9y3oF5hMTvxav+WwztDDBaEPFfvJLQSvBH8BkNokN6QHWLuBKH3hylCTbmCngUZ
OmynI8drllNO46Dh0LezEIfkB9fqdEdsbL11eXkeKyKTmS6eNZfXKQTRuMYGOgDRhsa9fbjAtotQ
dMFWTAFeEo5gRShuLKGxGtx0NI0/8fja5j2lF1r8mK9mBjPy3box5lE7gTC2xkhgDBM8AbqX9PcA
OsGdnNYtjqlMjM4exy5wOeJM2BThYq9uJOpgaf7PRbWaBx/gKq4lfh7GeBsFSkpLP7HSsL+Cxn9a
ENzLm/Z5a9QpV0UgtlwESBFtvVXmP8wBXsZ2ZEMITZcIQf0scc7JRyRnIEDsoFwHg5gRA8GDwXzW
nxVRgufGOme2EeZDjjuljOstg7iSHniWCoVSkGLXUr8YXHGVCMXdubLOWTRjbTF5G5G13jBySy/r
oPTmkqNHXmmII5nnLzfdzbCI/pQJ/u5LY14KDJs48iAX+tMhKwfvkLeI1aSLTDr+g64FCed8NBLt
3LQX1PtIIAeFI2Iga6E0zHjCAbRKHGKMwr8UcJGW+CDbgjvzIg7vD9vsZTRHN6U2v+72iiX18Dt7
vdfl6IRJ3imM9mcstuBqsz+fHbAtwo+z9sC78QXjkHQdKgBuUmqoVWSkH9JvXHwJ63QFicH+Y8ph
iHAacJBWLfCS2N1s/D3BjJypnbd+yvdacKiVU7zBg7Gx06Ynbf63todhcnjwy3V7AhzE7OXQw8pB
qx1ntByMPTJscjesKZqlhLdfFahoZy0c7gqgfMEtSf4o5lgYJeDy3KrMq1yJYsMqS4AJdpOkYjjV
yUrFEuIhZT9gWDSUHQl9NUlg2ilyHCM/adPpQIwYSNaVt3vz+2fycJSGOhs8z7Jnwd4nXSwjjKev
80pnfoPSWG+B2AlFOuRkoACFfxmi/hc9VHgJdOawxy83/v2jvLnMaXdbjm2L56K8kindWFRil4TW
E1CqB5sr+P/0ef25Zyri+2FfFv0SDX4CzdwQvhvSSWiNdJUlRdQlgAUXiyyBYgfHrW5e1PX2Kzgb
m8xlsuWG+udH3Y8NfP7gkGCAHxyXtbXyq//n2EIz4+7QGMUDoC0puIrgITKRQn+JGeO3luc3Xbqg
sBufqlEVH7jqfQ3oM+kW/ixS9RqyBAosVZsiOqqxbhF03vXhNZ9BzRoDtF1tZ9PSRWWonde3THjW
BbkZzMTLeaO+YBLDzlXkX3ZMIs0NVRt/EFvxI0/ISTfOyPwb3P02h1pBr7YaJbI0R+c8j7LRYjgF
Afonwj2P9CZOqh1UlPjgV2NqCoMhhNxtVZN85WKaxfHlaEVHluQSBqzxfJNkICcW/YYEXRTs1vgo
4cxmwbxEFo/aJPR7QdiQIO2anSDUuYCpXLuAcBNb7ufuX9NKdAq7BoAqwxyV3PUutiZVvJRu9Yi4
pkP10CJbHnv8Oe3UjANO6LqixeE7NJbdQv6lS2QVFgv+AWHEy8/Ytg2v26C79zekPTiNkwQM9a5A
BgbiWzkqK/4B6nWcAd1IlfFsW6aG8pwJp4QamcLSUYl2VdoYYvbGPP06RGhOy3VyF8T2uN3rQK1A
dAkhL1A5ljN4mrTFdIVNoEKU3bwc7OQ4u0gAbJ1PBNdHW6oaazm/GnRe5RwkmPgu1AqA8jzvfbBv
cvzJG/ZG0HIodvymudxoXNknfM92B/2XRC4nT3QEAysBo5r8gO9ZUaF81p1cBPexyj5ON8ZrBG6V
Jar3zA5U5a/UjD07RH6GwEYeLAZmnJ8X3Map+cbPK6+l/R5RChXURayCdXdfUFjpb6M5IM3MzAMi
Lpruan3KR6nHXbv3RPmt8rsaeH+SLoMuWbhgjh3a0AF/dut/QZXwzz/fDxUQ/9yyQeaow5Mx26YB
pWSm6ViZjhtvztJ+FODRUYcU6MhwDv+48V+bXjUWWp3my4fzrXE1LLZ0qgH/ziKoV9Cj8Ki2TdEZ
8n7ay4qz5qe+GTV6BHWZt9km9BKFt7523aO3rbmjE1LQnJuD/buX+W9+WruJCo4b3m4UyY1KJ8Pi
vwIP/tV7yMHoFBfAU/iwpKfyQ3rYTd6eBAfjerO3pH957NEOWmRjklWSLuiEuoA6rBDVpTL21hop
f5yZbLAvFYwP1JhloHIZBqhd06puZp1VkMx820wMgA/XDSBg1U8n/3Kmj9dJOFpqrDhZBte2gqpH
r4dZoObBf1WW1L0v62KXqJx1n+EEN5cYX1w+PlpcQUfcg3u4/cewK4YzEdo8XXmMDxaSf24X9z2I
aqrg+LGZAdmTl8t+aigwcvSqWCQRX1Wz+3XAfJujc9rpQqNtWVtGNP9xFHuCP+tKnSibWh/qfprX
zOPZT9A7Jrtve/8epshnxEzBPMpKeOIFNzmzzssnrm47M+O14suG+GtJ1hO0kFKQZxiiPO0dWD98
VkDGxevv7EEM9Y3AEOakZbokQz5GkCFu6avHSkf1h/2uBZGYjoaaYWs4An8lHBUqHOjTSGOW8oRT
ysqMQmcla7wrE0fSZ/VXyaEwVYapB/eS860AMW7nzNAWER2xABKQBCa64kux4jltjqI4o0vJhBcz
Vyfxf6mwcTBDZPpCeev3D1fF/h8Kwm3Z+KKcknrN7RZ3iOm37c1y9HqEXqJnFIzRAyOl2JXRL2t+
BvH0AojN/3+/JQH16ZX95rIHybig1cgEdqMoOuHVV4eh+O8g7UyUkCRDzjch0/awRQClTgRwDTWY
e192g1u13ua/9fgrOFKUyTYDCHftdF06z40M32eLmtowJYf7U6ug/5OEMFHAMSg0fIFt9SUEQrcu
YJ4tXnsGkxZnAbxN0OWHzHSQ8oakI8MtIVy563/+wq3LD2GPiS5E3y9+tmEooOXak2R1zxTqu5Zi
PzR/opFj8pZRQt6IYkqsYpYxXSJ2u88i6jgy46ZiS7auosMs3GcFUNRWG2ARut7rx/TeO3qS3yCl
82SBhXMuy+GA9pHG388DqwkoBdOztrZLFCTqrrnS1+07EPuo7JK6qAGODE46KrnjS4YquPkEv37w
AnOkEE4NKVdOv1u0Xi5Ufq39MKUJ7VnYAeIbwHtKNuWRUhKk6cu8Aw2RXlMSTqa6uPhMz4O68itU
G8uZVRH/k4dWNv9Tq/kFBNDQqCfvJysbbsQ9DATDjF6YRfgSETyvR9xlmMjYOnswAwiuCqy9haJn
5DCtYA3NUV1FaOcd6vAuLGvx3S7Ui7t5Tb7GGaClzggO47XfFODGclZ+gtSNE/9vgKgdm+VTdfwB
4kGpEarIWdLwfhRjKqEaobxhI0GZLVsP1+gPCSoRl2QUirYMP6LWTy8l5WKhwng07oENSnphqwht
WWJizYXBLSow9cdes/stAmKjERYw2rUYbfAeX9Ors/BGPsS/8qoVVYvY7o6PuI2AojkXQjo5fAA6
KiOjyN7uMt/AS/nZg3ltGmozaZTRi+sq3ooR1a95yWBXBlvTPKci87/ztmnftB0Aw+kplbNRZtq3
tQE04Ej9J5sujREyphFmeJvnw4TSFbUyq8GM/6Bvi7Q4mmwSIWzQ7Ur8u8i502wfQ4O8TFUCocNK
qvqvIil9fxcy3rvDSFRxhU4ZleJBWjbzK++ym0LoQHFKZ864A0alC9CrBWWptfGBqPfh38cUW13Z
f2jyLCEst2YWhFEGzt7bicWvtA/Y+V9jMwAR00dyXlyZIoDfdKun+Ihjx+y0e2qNpkcHGKbiyzTd
OVF7ofAFkyk2Y8gT34W8pmIky0DvliOg/qa9mFWcdFiGFA1+IMq4CENvadhT6c+8p+UNUMNKnGHo
UEmJtk/n4FoTPQhs6FjbjKxW30mLvnWpM+LFZ2NqUsoHayZSWJJUpk6X0QQCAUwXrCvblKVl+Cs2
2VyP2FmylTdpSFXpqX+djGIVUe0Fms6RACY22vBqVS1f2M9XEtb0RZMrdxOIczoAIGbCWtjC4bz1
vzX3xVT+N9HwpvJSloi9vAu22vS3yW7dy1VWOJTxhT1SHZoxCzW/64Kgw747Gn+KTF7HJufYC6Bf
GLq8RXrjo5US60SgVC4tGOFYXkopcmDnAcobI7y6zS91jueLbHJz8yQWsFacN2326AqwM/ZBtOw3
CRVlVpTcT0QKgLsutQqCnUXKcaPlEqsbIO/UUWuj/exRwSVI7xoXEnJ3F/sCF4NPfn7tmd9REEY9
3a62I0LhrgXEnxyUDDV1SnzO8Ce/ZoyaroDEYnfcFsplatdDM8jeku2xVe6f8DblaApYsSSLtmQd
wDydPhmd4vkapq6EhQ74XUt8b8vj/2WRRIb8JeNDO5HVKhAIsYRprHMQEE1HcdtNTQrGsKu7pZYk
43sp1NML3Vkxszx/YNdkeoALgajLqNOVHvban5VaWmR3M2tTvLedRPsdM1JNnYdZdzrZ1gHe+J2F
idE4aqjqmQVmKMwIn4dsCueDKzWIh0uYJNR9XKNuN/wfRwFvUhM6lHlmMN62Y5N66Pfcyc05jyZG
/Tn/jf8UQSE28LLzr+A0pzs9gOfb/wlTjdrmyfjY9fB1+B3BHSThm0Dm3PJv/xsWiEXyKhdJq5DR
8EORVQ26F/SGWSlPROVsNknkymanzKMhv1mlJhT9HY6882vIGFS0iJVuQzayP65t6KyYctzcJyws
WZ69NxnZua5xOoqX5IvFg+XathDvgZE6U1fw8okYqe2fmyBtQCeXDb5vF0d1UL0Ez1QJld/0vCTC
XGD8VFuxYbN56ymyESb6zQHKSO72F8XRrQ/QjxkxryEiDNc8Ehqz3vtPV84261itYRTwPQnq3Wz2
l53BK3e///kigH+kSZvbS4dMM5APeVnehd8t9TQPE+bviuWjfzipf4f3O278JqsfjJOy7uamQ61u
mQc1n38aX4oxqRZzkegmzgueYAVGwzvXIcQUbrvSeYjhS3GiHd/v1jE20wb1zDbX1yc85Xw7k2HD
clb8bU4EBhrpkC0W6cCj4KuGKJUTixJ8wxTyYikgQsMlel40tMyqcdqCidHFH6y1VWDm54gV/NBb
6h/sAF2pyhDEJtu9xkBA1OaKvl7aX63Ur9vMC5F9o6nbdKn64ffbdWLkxxyOsVU6yWd3CJnvOb2h
523+9AcoW5Y7DN/uDpydIFNX6UQ7RZ1j/aX60uS5PGEWAZhGp/OiCnEkWdmOi1YExdAz05/75xJe
ej6ZxBCy2RWffC3DtZzoJeGVG4t0JrGlSk94sjTNHjY4ovGan4WtcP0qlzYZCmU6JbufzIF7+bJL
J07Z4DAOPINBuAFzMm2EPhtm8AjtYJBPNSv4ceb+QlO1JZ3QaNAAP59F2kArxRMtcOjJVbq9Lm/Y
9CIhM4hjPr8aY8At/QYKxOy1T5KgBwHbaB1VTH2kTm53U0Icdx3lRit6x4yc+ELox8SyGzvmzSYj
rhgR+h+rVQHyH0i8I2/SywTFX67/dj0O1vewUYF+vomfwooHNvEpSU11Gp9gRrKFjQJX0GRzmsuS
XpFVSc774WnxBCmxt090HeD7c3v/BKZ5ooilKqpg3Xv1GoDYUdT8oxsig3egWqfP4CErsSyOnTSL
bmZit82io5aPwpDBS0P11IP0ri7cVLfT+DkQPueTvZ+rcCDxF9XLdZQBF2o6edrPEuG4DpttqF+g
cYTLZb+BBOctGSOvDy12VJyKapVzenZUL950p8PHvWxDvwtorPask7+/UQdgC2qlz6PI159CkhA3
Mf6hxHGC/0anX8CUmvPwBodUutn71ollQBNtjOQCUtYBqlMBFl49a77kqeG2rxXwRWxvinF9j/V8
NgroF02iPAjVhXjUmVLlHFXqsqyhIe9rBCMwLLE/vI27/1E7RDfCaQqdhgfeEacs616nobHXT95z
e2jZ20zBveyVaAGdFKDa6jNaaOeo4NGXfkPmIxg0L6ZjrwEvk1pjCzu2ZXsirNfj33CvNMBaqFvP
tKma1aZo9IRbqk6FAtBbt8KhRf5NgzC/Qt+PSgCjfbpBx9RHtDxlAiTIaXSaaxMA6SaLeLJYgavG
OZB7Em6O3rofj1p0kzaNDmsNrskIBSYblaeO+J7DtA6bhBd0KW/NorPay1dg2yOsSvr7AVbH4WBk
VehuuGZMVY68DHg3jIoZVIWGccsZhDVEzbvWWDVfU7Ib6JhoPBUa3GQhaluauAjH03WzmW8Nk4zF
LvGDWpMkUBdTDmTckpEXkrto+h/eJpJfaEVfVZ0bfGG3HVVv7ifWGcRnICN85FWdm44zaGMs+tIo
fAuFA/7WNp4CI22iZGZw9n8xdYAqZ565BZ9VlYhFbYVjNDG6FN43uc+TE3CQSYyJQsu+9gjxjwxd
doRSgrWsZZNC9V0S+WNckpI9AJOyTALGTnb4z2KOBx0gYTy3S22/irv1DHvyzBpOP3h86hDLaatX
VDyFPeSa0WsbzcxaiL3wNmfTroc/IzC5hy489cXZo3VTh6xXOqAMM95LzxhleFhBs29C9QWiCnYO
rWy/VBywHUUKKuuZZH/5IB33n97lQDeMK6TmQ4aMju+aZm4xeu5FwNcz8QfZONdrQ6nOZQnsm2gG
xHDQE1eQFiKnIOHuqGDJ/8EOHle4wrqrUQMrbhg8U3qM7iWWnv4b6wPgeOW/4g0pTBG8jyekWRc4
fg7512zvdAtzH+jtSNpyCy8+X5ihECE4+Z8KDRo961nLT7sUSqiw39Qd1kDI+TJJ8BxI5ivPkK34
OYRBncIc2KeWtcISBgcvlPtV/Cqji/on+/yMzZIhUQrkAzvYcWREu697qQjQjijvP56SRr+DVGE8
t6n3imdJ9NqXen7AvhUYfnmCUAq+fvc+tb9xYrgXuuK0/u1/pSW+hTGIkpDd6qm3xHdnOsAkr0AA
/rPV9WzbAxhHY1gDfVRGRvilE0uT3JcM4rVQsl1Pjd2HgBX/OF5SbuYaw21ejOLkImEWr3kYTvxC
ih6VBW8g6fcoMMyGURSWVU2IlO0IKszF8+t1juxFHjtKBv3UhSoUYNmBfNkYofKcA2q183EKSokm
39yoertRLTSONjgQ/1OPJCrLCDB8o6YkLWrBQgANT82I+/bieNvw/l/W0luIWvnv6/45W8xtQzbV
+QRdtmief1f1aZz8kiWi411uCrtmIb1DvMGdeGTxAe8YiYXWZ7L3A531p/sDRZsaCD4VCn/f5gJh
dClvNgX5gkiqi6Ote7UmU8XGq0CWHkXzwOCKqZpgMPFaPIQUCDOFzGqeUyy/JEL3YUJnrQRQJXrl
08Wc5QlrKWgsysu9fHnoNEwGJhVtFPc9mvzOvY1nDeicSWAlSIEdxmDlEOzJ5HGTAB8O/+oLHsai
32P3/wDkBKGuVwLeDJeomUTPVFwnK9KyQkoj//wqEyHqOobC1lVPDKnhBo2XkVQ6B2JUpHmpuHwp
sHRoQYMCzEmUerQ4/np5SfhMKEtkclAnIBRRbIBkYkmPwvnddJb0sTRsIcsEgLObtYkvb3Vp/Nxj
mfqpIAYh5hxUN1aDu4oP96jEgFBiffUqmaDwXMJQtQN9zyx4mahjUEgRbL+YF3QjAUw314GhU7js
Z+yALnz45OA9oI0vIPXJ139S8OVo40oE3lzqmo5WEItLWL3dpVrwExaylCgNrTLiOa+YmcOqkKdd
hv3Qy1yRnjx6W6e3yDxPCxuhA+BWp7zXD3wOkHcTGKXWcwVd9JEr5dB/DFq1m/yXxiG3JF0N41Cb
z30fy1Ocr6qZt2KXc9vvdGeKMBcDRuya/QA6ZBKaHXiK4ATRuv4RlLAJv9U+3OnAE8sf2r6wrmMM
MqAuHm0r4bhkV3b1f38TS7MhUbU/LafxuYVjwEADCdByB1A4nAiOOsLgEsgqj1072UNthnMW822s
DgfCeAFDO9TJZ8EhijBWiq9/Cbbip6nbpsX0SfTb1W2dTMkbSa2ePcX1v8/kGm0GsF4v549SkUuZ
J/NLtqU6jpXs3t5R4VM+Hn09BxHfEWRN6lL/Gw/ELFUdF2PDtasnDIy8swCZEMLBWqOxP9dRkPPc
Zh1EEaQHgtY+ToahX2O+VXUx8rdEhFMCy5aqcvjluHzFQXJGF9fi/lNHtUX5FbOOu7Wtu7n7HP/j
UyEIpHagL/GIval3qysATOi50ZysNet/WSPldlb64KouWBgrrupZ21vpMEDKWnhV4+jgJwMYjgco
dXjLPGy4WZ4uY7Zv8TnF7dpML2nhoyEKDk0UjcvMkdNMRPR9lSqQWEZn6zoTWlNYFbrGWVJIrr3d
rKV8PSzAXhtilq7BteRKnasid/9MVhmAAAXqKqefXton5LABMtpm2mN+9yZYgULYzi4j7sGeGE2U
cPA8O3X5J5bogTD+CpCAaIwnQBFbNzzjfg36X66FFDrHsHDxJvbjNo1TGVWB+r2zk80bqkTVZhOJ
xVn8d/SQkG8thHDDpDr7LM9CCwHdTq4bzRrLkjOv5N/DbZTWaJOh/IaTMRHZ9mIpAm0xGv0iyoNt
4WviVK/8E83cmMLtz/VS1+Mw4fqPCMDArYhfEiWJwNzfpdqrtvmPrcXozUmA0KguIQvtocoRfAeN
a3ar8syHj1DStdoYCye83kbJ8cC2UqiTvoFXFlJIsnqqK2D2Q/Upn//c8vtQJfBOWym8S7GLBWWb
S1fV5yAgH2w/2VosnumibD0Pgw2Xo14wz4LG5xgstROijNaGmCOrRkQ5DzRJ4Aw3H2+ahJgy1m2a
1CdRs/dnUQWhh2ixw/8LYmpLFE8aqIC0ZF38jXI6v7InevUk6kQlektDE9/VxC5FVefEIk5b9P7R
VIfn+CfaovafluwPp3uH4k32mLKrqBWHx6FqXeVcKuua2RBggnCmgp8yFxLCh6yvji8Yfk0AE94p
n+sND2/jV4lGn2gKCuI9KKz/gVjW9JnBj9robNhhiZ7ONxXiJu17a+q1vKh80GsLKv777PLQfeSl
3YcAAHiBNFu4/qy9EWbV9oimSutaRacyqcYKcweKwU54f9xdyBP1BwFoUMPlAoC+HMGlgCWCvCPg
7+9JeNozMs1eiy5314IzL8JW8brQKUTXoreTmSl0LWtd1/VzoUNPhR1zuLPFrgPCp/p9L3r4fDbA
nKXOA0LgdaKN/KI9i84rHCoF6fMqjUhAATYNNeZ3puZ4NnRzjDInpBpMB9qhHCVebAjxTjIn+oAt
NbBtSbdLF22M5alL1cWc8os17eq41Swq2aETzyslBBqXaipzlmFWNx7SOH/w+VKUErms2CrAInC1
SO4lTFU0fVyFxgfA35h42s1KGWsqi+rRUtZAaOuBeupqVKvFCwi3KZAqNcpUa7ivxJItrs05nnMk
n5K4B+QkgnBl0Lma9tstI0n3GGU//rx2s3jhhQ//L9Ni7vMCm0y/sf9fDUvunhzQ0CIo9bnNRTzM
LBoMKKUrHkU55HT1H/lVlBpDozhE7YAF85+To4J1ATqPvCiXZArbhzR/KCPS/tmviDo/+S8d7ex9
D/sXIIhU0XQcSlSu0+CBvPW2IAuV/lr1x7fjokgqoSMSvgkcFZIKwK8fgAuBN+uxwJMUeyKIFHWQ
9Qarv16bk+ArhCTtwdZtkLH7cfDaj/cztGDlmh+FQIOEAyfDTHgv/a82CXWV41nY+oPHysZ3Wd/+
IAKoGePkd4qHiQDVDzP6sN6FKRl6ul553lPlgG5IwpCBnmC4bAQnL3ioQhprS9X3etZYXAvW+sQM
08kekTUEWahOAVaaosuRwKFT4QJWb6Vnd6sEllqIpK8CueGE15ZZvqju4dsDSlTW+03Jc7bzWQYD
pSqCzOT11NDPAitqJQDWFStRyTQRyBbF68aVsLBUxhaZv1JIe2Kb8CiAXYlrztEkMseII0zmjYeM
XlKLw4m2qlL1WEs9n4V38+NGukHYSmKqL/mxKqP/lHlfKKgKaF+sD+D9tmkeMRYrKdAjXNsETdna
bRYqKMBfJF7cZkH5lndPB6wNtTGbZ4vp7ZpHh4JDG/T2GsRm5CiYlwjEP1U4cBJ14baukovZNQfO
WhMLo8MA5O0al9D26H7i8oPjiZngCcG0qbpqKyggUEPpSDAzlmFkAC650wyZexBifA48Zr5lephJ
ADIboz5n0BgMKjAM6ZuO6p1AA4ydfMlsGjKKfGgOU1tllXFi9bOssacg+sR4nxYYlJSw/RtDpviZ
r9qXu3gRssCHPVnFuIypbxhIiXieo6DtoyRZTGhMjR76ROn4m4KGPLIMIxHZu+LiOdVx/+dNtHtt
+UpPNQSZxDmzYFw4bl0exFc0ysQUPxZgY3psuXLzy5t1Z9VZCp96Q2KeZOl8k80Bc1jBKYw/LYB8
GC3IkLjIz7z1Rd+qDHV7t0s0Szm8ZOj62tUEvDXibKoTZycG4YphdCCc3axwX9vnINs3QcDRFRvs
+cwt8uzFAKdXNRqozJzT1him9Ohbh5uBWVCa4dHBvCsvdKvSfiig1GRlMOVzbJJJ2VizaI/k5vDJ
MkCCo9NxbCq8lSCWLnb+4LoRxgDibB+BW9P2bKP22GgT+3g90YM4w6hSapkGKTq1oOo1lqaxqp3i
+jh3WioG5fSzHz9NOLJ5oMQ6dVxsa06w3KPLcDG45VMm3EXIxvu/cEo2Di7Co+d+7dKRrH4KYv5a
OJWi4ELOJ9L5WdUok3gN6ql9ivIDG3+VaJhMGJICywucsABugxwn+pNYLD6OuKx5TKtvgwPqLaUT
4KTNg6jAjLHkGEBgh9nhVZNn4YroOtUvRA7pbfDaYzACq3+IRE/PFiLF08Jzn1yGugRSifpKWUaG
fR/ojXxjd/5IVzQQFtIE5JfkOsnrouRkqPeU1FdxzoyStZRx32fu7nvPTlRfAKpOiFPla76+krGo
cwHfjAtTyVjIKTMe/Gy1TD64cKA1t8hEH8SRUW62yfMUTClTzZb2rjORNGzvrI61rKgaQfOaaBEC
8yFvbWIJ6ke6ipOJdvSaqDfqpawraZPl3p63Ez/vK44H6hXeKGJWS+z/sckvVBBZeVBg5NAtvmeG
KcZ1oV6ry2IIF/MHbMjQQCGUg4EI+5ooEspXCUwyA/kfQRGCiEFQT4lSTxd2ILZNuSuKUMeeUCxg
QAEAlSqj7WBgsG38ENDViqdGx2PhsDCHqeXOUplBw233titqbVTurhAASaJvtkr7WtHUGQMK9mjz
6B3Z2sfZe0Xfkjqf2CRlatOP9ridYrfDKgISzRrWA6RvnRbTclPWsgt7RJXIzNgE8ed6ZjKGmNio
/8m+bEID5UsemqbHx7QEc+/vGfsdgD3Rb8sPOaNqnTRBeu+7EHPSuBG9ZdDZuwm2n3aM1HdkT0Ta
X4tBGvT/QMpCyrrx6of2nuYP9ZjAdNr7tgWgvop1LmeSTit79ErGdBbYjpjPHEXd2pPgrR+7rSRR
q2OhNDcggjVK4OcbPMbB30RkFdJ+z1KB9HwAjTyQ7/9jNH3hLBYOC5SzDiGraJfuO9mJgkZ/4qRF
+N5SMOsxUPcqX3YMYTD6Da7rd1EJxVK86c0W6ER+MfqJmiBm3emGjdCftKVElEB3PbCPvnXIXIyC
rtSMx2ld8OzuAzJNaL3vpIilF+Qr+tJtLtwYY040zBeOGNi46rLfYXyO234FaEItmdJiRPEfj8UU
68XbUn7G/9bfaFrv6EGJGcWFFSXX8EkRn9jvuEUURUmXeESVCoXiMqPERjUZ4yaNByFHLzfYyRoZ
A+1cxkiNHvcQHGjVtacvZl2+4YOiCrZPHj3QPQjzueBMjVN3/q9zy9Hb9Lixp4+Qtporw1Ga0wDa
tvEehUPPjlI9JGe9Zg4h1Of9xNCKJIWb9RIo7lo6m6tKBckyyxsrRIlJvPUID7bpuwzpfWo0i+Ox
P4ncfzga86KiorZf4R0ilu2V0hSP+HHZqoxEcW+VEsuAOS9q4jNeP3oI41FvheipyFL3gWB6Co5t
7ajn8jGqhPcigz1fHyFtlv5pD0lNX4xopTHwnQ/GyWLCS6RfMvAOn1N9biiz8QwFpL8FX0R6vZDm
s3YjkEMfTnMUifg8/G7YczKSpnZoqtRO3C1yIoc/v0xW11gxfoulbIQHM+wpTo69etqO0qiAvkLI
R2nNn36Rx7i8HALNyWyiIbwg+7q5Uo/Dg0fYuzULBz4IamjlQ4cEk27Ul6eHqHjD4AHDcowH8nLH
mP4bjGBIUi9JfhgFFjX+WW3BaN0+5rA0vqi3VmyQJjywluS2VFlsWc/AmBHUyQXlFay2JmIYnYXM
8zAo7TpZKREBPix7JAAiJjx+9Canm4+j26ctOl6YcudwKPJeY29Ywb4VNUixSofQuCmOITJc0Pq+
KRuH3OV8faVX4GZZO53NoAGvS8rreViMXP1AB9AiLr0BnreX+MA7FHijyXsT+UPV0YUWwZn2IlMe
U60Lbnl2HcOHuLWfNO8BByFnHuanf2yG1G6DmqrT9H732yizp285t+GzCT/LdT6ZwHVwEEYwlqMU
//AXHy2clCPMN+IUKArf5vVRzWFxszmhPinlJmCkE+vEtLJ5s8ReB5DFdRFrPeXm1PaxgZ/45Fks
AH2jV9OptZG7h2uAl4ZI+2bUzyr4EvdFEjnpX0L/OH3AeApv2BXLNcy+sV8ISMlM8+yku8XAyim8
vRmUnOpqxbhMTZ4p4Vt46HCfJZHcmXnA+MASe5L48xbpNYBeHaOS/FqE4Pg/Igs08+4/Fh0j78zb
ClAjNb7oC8qqPdKW3GoEVl9DEzBYyo1b6BrtHU1uFLX7KaeDUwu4k7H92kBgipg4FrIj8y72nvrk
zAskSC/WIcQrmJMacu7TGAzZdPEdg8iOIjqL2i/ZcDm+bYGt/vWXBdiUu1fcsAPvaLaJSCBAO/uw
GmxT+AHWnixRGrdXLjXYS6NelY9uf9YL7ssIIfD6YzQL961A7ivZF+iOdtKxBi9Dyq9Lg95bHXkK
mNUdSk3Mf01NfUTH8laZIE34q54+dgQ4LaVSZksOLSShVTK9gNtemeDO02+zPgZtDsaLE3EV42Gd
0NMmqQCks7I/MCzq4OurxHmTOgxpwVkyWfhkFBI8bU8JbHTonOEM7YSns3Kl6UQ8u+Vg5H6zjRXO
LJIpbHM3XzrW5VAYvfJMuZz+VWwQloVH3dfIiltWdHWHMPqQENHPVwIhuXL76ycUmHrhCCZfyfuo
nkJefvZercxBum5CPuSkym4viT2+ILDFZSgPjd1g8zGXH6aH4i/487ToNoz22pMOXb3sJZjFzwOr
QJugWDlkKMq1iq0t9DBjChzDoVash2vFoUH7+lkVBLrEn8XRwbAZExYWeyOitZnsPMfBOVK39Ft0
jL01LbLNBFiy9dGfOMfeAee5NPFl7+0XR46ebqREKBfwgxJZLuPIc0z6SCeN28iJCif+Xfn/Xd8k
um32zwMEwgg2ZNN0cg8y5MoGMeAd3r4XclRYiOgkCsl7AcwEW5trGFAYP8hDjKlDqfJotEjz2KtU
meKAbo2lCGeh1sHqp7xxGt8+Rn3wcnZrw7vtGStee0E036/mxZTnshuoyiYopORpBc1+K1/ytJWF
JGg4uwNFhMzGfVrxR2fdFNxdans8NBefnIlZtwY1nzXPCgC1gdVCKnct3g41qUbR0sqn45hIH0gi
1J6fyKfOnjTcC6kezpLZjfgX3Y8QGRgVfkULeDfvYPaQTLSOoqievlQ4VNUL3UJ7/9+dUpZIqpaP
udvhJ3mSTKkZv3mec44jb5232C+HTXRDKb6HSZEjt+EXaeGEu6ujvdv+A8/SA2uWOM83Rusx+BYZ
d1NwwTUEzpbl64blLW7Vk9R8PpCVAHoUzGSf+giVRr2eFuOfJr44v6rwYxx2FOu8kUXEC0h8zSQh
V3Zdalp9sOnXkNblk3JMfWPaLHO4tgtHJaNcwqr4UWrws5E/zxmpv7pCyzNy2aIVFm3CRtVPqN8G
q/YpSoiYWoByU0k2oKAGk/mA6drCYC2eR4rD73lLYAfkGoToGxGHGDGwceDRhOnaPs84P8hXurfo
4w8BsxK6jXRJaxcvY8v2GegIqavr2V/DYCFJy22VEDWaeWR4CF153OeSl8ssS2Xy7QYpBe8rCmay
aE1QfrMifx0mcv/3kC2o1S1rBoV1sQbBHEU1ekFWQ5JFblupujah6Cr33Jf891jMZSi+mIC8Xbom
ATseKDju2yvR648/VfRJbOeYM5emuMi425hbawvGGXTX2++oKHd8C3UcibFbIW+MDtIw3kMsimqV
197+NROccupRiEVtE7uMbuENkJyG833AM4CdOUeSxPxOuPLwnhVRVC5afWcIa65G8fn4jmVjN8gh
R10EWukmw3bWWhLo/ZG/Oqn1CCiZ+Z4cK9OFvgpV52OkPOOt3RQ3OdujK/dl2tRfsmtG+AXNuhA7
g7TT2oMIHt6U6zD7kjq40+J67QNKuZ2fzGhEuk6WxnXKULrij3ZEkY9UzUAoFJGqiS8+1fXe+MGr
H07Y9vhNTz/X5AZ22XyBB5A3gN1R99O9AQ/r+dKbU6fuULe2wIj53ClIeXfX19ava0ZuOXN6jdTU
XVjcj/+h/vhnm8NbHITqR4/UE7D8MBPCXeLmmSIJ1yFqI/HuM9aeCiDwTX/KOqYkorL24sX1IF/M
eyPwvSWfxmQqDfI8+N1D7vcffQTwgmALViwu4GmZLTzAI4irLNTrbKwz3gr+VnvVCn+W1A10VXpL
KUC8+wi1DhSkHXhFfh9nDUxrDyBjzUUVwTGtT5y0P6rUufRR/bxL3RUOcTGx+44vKzbcA9QvdLH4
HxR+lnqCBjqncNeRkKEcEr2gokKm3OCetWWWcZXa1ARzLhIDnUsFd8jg0KlDRVwXPuo4sGHG+ZEd
V9tCA66uNQrazGVHiUDuU1z83Epe+S+7+9LB733+UjQZc0v3S1bmjsgxiamK7rdf7q3oIF0l288q
A0uhhQsbTRQaTQUaNUNX7j84imvJII/v69qhT53aWJlXWRoOBDfc0OdtI92E5NvUZFrDLuft3YP/
WPeEG2BZTpFGSe3b/AmZMwVS7y6qXO5ynX4parz+/V4I+jxx3fqxREVy7Qh3FhbpiShpJcAnhMDb
Z1x+og73AuQhTf/HdaKU89Q6a76TUXm5FqLgbwyYHqCCveAVCf8RxiVY4NMWu6lfjBQn22PHL/HH
YqtGKH+kt032kuVB/tY0NuSu92qIarn32YKcdy8C/DDaPwz2EPZAu49mAZA112Cp7UHGvx/t3iTE
Yd5UWGxb5k4iDh+7JxMA5s42qru9BtgMIXnvqOoVQC9F4udJYVw5tJgqbKMrwlIKD4iy6lByObHU
CoJvOr3d5tu4iLjtpZJnP8YzYdFFQq5T7CALcu51YZ9eGwXl/9RyrMqJtxTVAvDULP/DxqDNuVCX
Ez6bfE+6V+Fiv9GZONyGX7HpGq3lgenwJysoVPLEi26dtpDZePGHSiLY/51oQxsJiYx9LbB2ZchP
y2N8PzfHXpjnV8SAMkhZjeXXOJe5eStPDyJBZGj7UZSd/4nKgYa0DNsEpEekcKSCrCqDcVZUW0Vg
SjBXkyenu0vTc3/2DLy7Krs03vbENonMWXkFSI+Sn57VZgnUkIAdIbldsq84eRAhRTDf/jtxZ2pG
x2ImUG5YWl/T1kRTc0ma2rM7zPxsdN6KNbgmlyakLhJn6nPT9aTe/hPbogxs/niig5dPNmBBGB+g
osmXZcgnmJbTcrjRmLfInVvgvBksz+c0Q/gLzhd5b7K5r1ixEpJ40StT63yXZwD3Wf69iJHSEMbR
3qpA3/zHCK6BBhB5LnFiMgZ7hUbdBlY3GXcuex4wjvzCq0wC0DhrXSTzb25qstmGJ+JDO6G7FV1B
r36nmcOvo43a2S1Aei5lFAmj0DEHAFXOG9easdgnjaF5LkkS8OQsSiia2ELMmC+su+DGnKZKUcU7
dTz7Cx6X20l+mPQNrwhDopiG8EtIIzbtD0e4tCpPozfFwMXvXlrjz67tS2gJiWG1fLs2ozXMbaYy
UrHrD6Hk01ndeP8fozEYdAh+Be1a1bnHBoas236UClhjfN/rdYaClaDPFcaNFzTvtVm8SvyS3QZ9
MIGSofgpF1rEELyzYNIpoV2ETR/2PgcqNVq35miA6NWJwLNoFnmnnDhNSBw4DhR0TCzYfr7P/c6F
Q9DcHwxeG9A0LhlKzbSLAV+NOgj3vQzuDW9uPcsmNf2PpdUjAF5ZFMnKqdU3aIcFkJlPlph5F0zR
MzP2fs4o9QS+ea3N9wkKrKtjjvpusXKMUyp5DGk8G5KMqu0HYrEq1IDyRNfj6bS0Ji2+T55y5SZh
W/Hb/QT5DD9xIOBu6BOy4BF3hPQ5zTfHwXRM3tAwVwm8RIeJjrJ6e383Q0ZMcOudig/ZRMVhs3pQ
Axu+mH4IgCELEQtbLWjWL8ZKt9vXp8o7VS+IsYUw0+aSnMe2+mxplIgzXqRe/IyfluCxGgZXBDNC
CSmsoV/WRbksur7nl4ISwTyL4v3hjIek2kHrbcuA9IeogFvlAyV2JZHSzqiAClkP0aMqM5Cwya04
XnetPTDm8V1SmxlSTpRAhOCjGSFziK6qMaD8R2zoH4XSJlCkFSFXFBFEUM0SBTW/NsjqrKAf0ZSs
ls8tD3BQZM9uUAets+8Py3yA4Dc8DMMSXWyohcrzxW5mRlBNnBE4LkBSm9owl50PWmWikC6PmGa2
3CjWOSUXxnvPMPi3V3YCfJCW1g9lYcEzsD3AlQED9sSn2DJnqTCNsSSDwDhISvJWSJjpV9C2ttOZ
QmK6GMCsSZkXeSNOi1+tb1nxjOSemX4DDGEYrX6jg7aeGgMQc/xly1Lc6w47/g7ZIU52dWFjdBeb
xUb8f+hExL0KkFwZAaHBxCeK++UbWbHMc1UqNpB/lsbo4W5Icko9EB4T3RPP16Woq4WqgNevCLzQ
3Qwfclh+dpfzV19aWWZSWfuUVeXNN4gbrEeRj6Cf5/SZVuedU9X5hKGbpRqNQm6lOO3G+ftAieJ/
DrBCW5lZ+OGoC7lj/l3p5hLK4HJYbLAi8wlPFr2i4u02R455DOsPvzfIg2CgHZLNNBPZXdhw+RAN
+jvA7pv1BdUOE9/I2+T4mvVeaWNadJ8HxpOsS9zK7XvW1iHrUZDd2uS+13tjiuQkK97lZyTWdhjF
Sdu9vSe7wIjxNUT3nlc0p7PeyYgIyGZHhMbD4y1OevdiK52awC9oRMmgibJI436GGX3K/KKX9bpd
TOmx7Gs7RcC3SycK2xneCWeyzTqc4rgcPjezPuAXYEYhUMc9hV5o07gjhzj73njdbFmhsPBhHRZe
2zp7YI60soF61zb/0EQcvezb3OHn5QJ1yQDl/DQBGz6OJyni4utvwMV5830/lA0/p5rvJsSkSYi6
8QqzY/mPWADL6hfgBspE/I5LD8S0gFgKrL3EzO2K4B4nKpJ9m5ZLUDf8IxBPd2uYrZYfqq/DD0X7
BLqkK4B+WC4MqTr2Wj55xnuYUkM4MgfweBhg88wHqidXKjc4niYIC78T9IjdGSfbDD+/9rJAgiae
o+9MAEbRoHnK3rEJMqrvui8ylj5hJ0nmv6d+P07RzC3/FxxMh7QOmIM21fOBFCCCyGDhLD2t/IxJ
PQpIdrQjXh09zPDe/ebLTCL9km8jO5ZQntQ8cJcjPhVzxsJOhKYgwfAC7ij3dWMD8RFkminxI1JW
hSuOc0pAUl75/Y6c6aTFeQFy6sFGoVVmbmi1jU3x/H5cqz+FhR0FUBAwkEVgbddDoaxRZcSMbMUP
kMTILBPE5j2V36yp+4M3pn8mhUA2d5qCt6QY1Fc55a2YY0GlwgxPciExjxIIazc7KdJiEKdFGzhC
pln6uZuhzN1NMBqNiILlPvQ5bLplz7UJpRa43lVGpDTnVCPauAclPrDkhBnnifhbWeg8ELlSLUBj
9sK+hBYMeEyNUnVAoUDSdJfKOM3ol9h8lbnwKKEx7okV6DysnF7lHhD87dbZ75pTOe+iQsuWgGhs
ldyXk7wplTaR64LrPjn8qjGs78Z4t02dHLx7nBT7N/x+usMogR3HDzWvbxck5g1xWLzFo1zo2dUq
JmdCEDOCPixXrREf0p4jYSfou1RMxBeZUbuO/5HJ9aADhAx8W5qd1t8Aj9NJswZiYlVizSTtHR6d
6nGYE0liJWft5QRHCvciJQh4t+YteVj9fvSpgi7Bg64M+bSulXwGWcxlQtGB0GJxWPInebhJgbFm
0myhE7p/ciwdoT5PJwHEpHSWROZEAKDy7+aic2fo2PrRqi7g2ubeHRJl+A+Qcl+yXI0ebwtVHcgY
ZnM+1GQQRN3hpHF3tbjZSScOYUYf3KAP515+r7CF7iKFHAEd8Lx4E3JwkEIkJrllUEywibV05Tep
bN6veNNt2K+91/Mt+ZheqAGqSEJT95P0Fe1yp+7UZ6qAlY7eQE58p6N5oVA3IIavJCdgZZx3hqzw
h1GxTBPx9/kcx/qj/mQ/hFM+6rH8gZ51WqK6pbBR8rW2Fk2/6BwmtjqbuWokYv6yXjbAw1kyUVnm
L0+HkJ+QGdpLLrQTzkxXPHMxjEw7ejLmGuDnpvgPOi+plyiwT3+elE3LabKSs28ccSo/E9b3/Xme
4F1toUw32m5D1FxGYECKbjQLge35U5OimVDfLq5bUmFIA1WgOvTBz0LYxG5s4NPunL6m6WHX9Pey
drpYoF7yF7nHGUw+bYz5iDmDt5+IqeuygTm7A03SSa0TpqRRupnwpkGZzhMr16X9h32WxKWSb+/x
YYoZ94kuEM1sAmhkkJHcJLFPhOgNR0LynyFAT4+VN0ViiguPj7URLkg+s8Kq6/kESmBcULEZE+0m
51ENlzhw4Z6uujYcEyUw5ckLDih7rCzStTW3lCsYEjZ7IG4SfQcb19lnPTzMNtJnwXwR1Q186ctl
vzmbheP2Wq+CoY2eFUd4dygNMhaG80kx5Gi2u9ThgImOQsXSyaYmthRyvixLvCwtNRS3Rl0HqYR7
/f78czxE1F9Ifvdcup3QXzDg7abbXNXM0if4/92ZYksTV0WllzJzHuRE8s93K79q6/Bpx6rAbJf2
V8h3Q0r1PBumh29YFbzINI+eOpKChGGYd6wfO7mH2ewl1hFzgQG7j7mGF43g05PLH0n1L5TqzaiU
fl2moXJQsIcQyBXIF6b59NUpTj/b8un7e5NjybVvbUTNGZF9MhrdBfADTviTdh+kpK9CPHUw7o3t
pUJ+06ZFaWbO/kJ0dxZ4mVtfHsHd/Iupesg8wRNCP/bN0JRoDA9TxgwHh47+xLkOIMpZTtcyonfs
RSL9RKiUTTsioOygmVta57/AL0B09LcX7keXjlo3OEEuTdtk8qorLcIXkFRlo2SW1quAs53MepAl
nHydZ40z7Oyi5KAVFIncocLH3hpmd12uSPXLIuaOf4K06yZSNj5R/py9Pyd9jgc8OTRnxgGdvBfd
8Q0bJjUHn+u0iU8Y0QZyZ5ckXX0PaKr+EECzvESQYomMtw3Z52/Wa4maQIzuRGObynHWLu7LaUfd
U+er0B6/YVB+hMjgaNNkk7XTfxqw4JdgogHxN878ejEs+6bLfHsABn7+iCTRLn0pQBS38qkUYDgZ
Impxg2HQE11r5rdwMtGpwEPq3FBsBgSIkCj2FFWErKi1DXNiX5eVBrtrd94b1+55cFCzqzTpFV2P
SKGVfwUFgk1/Qcc0n/7tEPG22MfztS565ls9CghegmIe11fw26WEot7x6UcMbX8D6y7Dy4dIHjAr
le8APPS6AosjB2iRGjkxrrfoupq61eTGr+bf7Oyim7WBfWquVhhpFrWSDqgI9mq+DRZVzjedPPyA
9TFno5M9OX3fj8HlNnP7bilrzFyds8tJAjXq68CXNhjzbQi0JaBloKrNJU4tMdm9gSucEyXSd2TU
w/J7UAXWtiblBwKVeJ4eQlNIS55ps/29l74ZN8OXzupOn4s9rzZbdzc7mR0vX+s2ceEyMuBVXzkg
O8pAG29vhOf6V+VJJNZMZgTACY7NDIwNEie4RaW8g/0Nn66g9u4GHYDTot64xBRZaEAYwaTWYnTV
/BPhy0kN02sC+09FmwBfLyzykvFi3pXVakRAuGjyvCZetpq+o7F32pK4pH8rDM9MKKePfoiG27UA
690taC3op1cEK5IfR6cJe/0204EZqhvgt4EgncT/WJzvij3K3DnZix02qAtlumANxw4O+ZalTUmP
FQi52dprapQZRTXlClZ081UtZaVGuW1HOVV+eZBLx3HMymcoXdH19UooDN7P9Xrv+PsaRS234uSA
p+jpNEv8ckeQ59iiF7X3Qw4QgwlS9xd7jSfpQRT759I1fmjs2y7UUQfmDBBDrIOmeL6r1g1vIosJ
bYzjtRtxtvPIbzWs2XULAOZPS4EubzIqxpf2fEV9MhgFNhOF5yg0q2s61u+bPxTLSeUctVPh5z1O
0CzjQjdJUHj1SsuAl5B5VSRrGgPG3QXVOBLQ1pWKmprERDFkEmT7LkHYFl+W0jKpbQKNQ6b1sgi5
X88ou2Uugnnm8hLi2SPpntUm0JEi9LM0TxT//BX9cL6ctz0o5pzSRqiniE5eB+bWhGp2b0gWS6lu
1c5QM8a4C8Oj9i0o/9VvipIQkEyts/DTZJYJEBya/M1a+0RCA7UbuZ/T/4N6cuTjTe1otsc+qEuV
6sYTvtInRNeT1OKSRPB9Q63x4tFEZ8jtQT6Jb70By04l6CY82JW0UiBU62eYaSAqU0UvcnrGgmO4
xt46bJPa0dmtwgIbdmvyrld2cTTJZGxVGBPgXAH4Lv/EmFg+Mqr7HMCAOzJth/kY21UUCurDSldr
dRGAiNGp3utnVwTho/kQL3Bo42luZIL/9v1f+XQDmO60OkXVzL22vB3Y5pbGhBwtNiPW3R3+09mt
KxzyamfeoXEAJaIwxdvPHvfP2TtZ8Gf3aTalZ3ktAeSnNIiWO80vhSzjP7g9qrJsEKj9vbl9Y+iM
jFscLGT2Ze1X0TtN7cf4PBo7CpD3C6i2axIZQEuf9dFnppP+8pnV5KbGwmB5taam1prYn4SvHpr8
auHorEwFFYb7XPcOaq2hsPgS64U6k7bva4H4URtjUrO3YRxchrsHyanemCMPrf/sVwY7xuwx6ybD
ikTOy5euFgXPkOwlCLPSavTPL24AniI4qT1R+dORf2345Gyg3sVKmfx2iTvXMldUtqCsKrbb+BFC
DNsyVQGD1mmagJb1Qly/S13sANz9ELafHIoZQ5qwUZNc8NErip8nU+7Ao3OnynjxhmsrvvnxjDTq
qMnyRCmwNbDQXZgimnjfY3snX/pWP0iUoexh1J8wlf2byM0XzwuYTZ6dWDwIIl5F16yGUE2SdBfO
Rrgv68oEe3p+Z+STOZEFep8Ks1bRmPGXLzUnrPM7w1wxpEIF4ZvxLwc39vB2hDVhkkXJjaz3LQy6
duG2C2EFN9jtURiN5Rg5KIizCZIAI6KN7K9duECXWcABSymDPwcfgX6Hodcb2WSupuEls/ZxqjF3
To02yxp6pH86X+87ND88rCYjPzzC9C3oirkOBVCouUp26+wK+7XU34ZQ5oXed9TL983tyCXNOoPa
Z9rr+omLJe+xixVHUHnIbM+y5ctuV7OzifygloI/OLcwsrGSQv9+ybCLEddhIa6OYYIiXINcP6HU
ZiH8snsfRK5kjmrKlWRRQxGyVfRRFbQWjUWKL/MXS2D8E+4bUbHaviaa5qs0C6NSo7fEjLIiZSLl
2LJfm7ai6WUZgmvHSWUCgysY8zL0p73X5hYtC3nD8Ifs0MvrjjNzb4/jA4dBNOaqmGP3Yzr2bYV9
EwdzjGSPPuX3KwOA58bbEW9wIk0s7cpcu6zECxKyd4izutFj9iKBuxWmRd0DqqZFpzyCST5vG9Xs
FhtXYPkxZn2Ci8zGSDi455Wja6qKdCEheSo1SEOeRCaB7Z0hC4WGfaPAI/6xIUcWGNKDaV0TYZr6
kV0+qTK2FenHonJudIO9o50S7Nff/f2aKT2Da6Wl50HpJ/w1c/rzXRVREmp0uovyYl+tsuIKNr2H
efKHR+qi64w6AZvNG1GfnGmzvHMVF5C3RuseNE3O0f+yuitDXwxZ3K/K8bgD8s8hG5StHOgaqRfA
k7U7E0irqi1vl4ksrnepdEHmsifYLL+7V3beetXDzSf3s9Vlht3ajmFFzce2j27n/ywZhzQZe8OQ
qkrtqBnAqIBTeq1r6exIAxYtsQd4nTommeHgATAhpXfgvPa+pX62iinA3imFMjru6Dq+mCrGMXf7
wCcmZfgyKV+wU2qTEw3MBNQRQQQrKO3SzGHXPfg7HG8YTsSwUa6AyEug1JIOtYM6qRcvnLfZLgXA
mgnQ+4TIsnxdfdcFxvxGge8glMDdNyiUcLSjKoSpOxgDxCj2zQB5ndggvGkWkL+Y61wfVyhzzkPT
8VDlf2WYR+H3s5UTvEKBM8FSFJJ/De/LxUaoizcBtUnLXWh9PW33MGkxcuhu2FqhGURNbrwChnpr
Ipy22ypUpcdQK83s8AFeLyGPNWY+h4VBYKgmpvzDUK69/WC6WEAmsI/D799uFv3BO98RUWyJCwKG
XdGIDGP6QU4tmJsSgdNeMCV2k/20M6ENc9v8u17Hf1ZS0BJKiJ0eAiuQDgQz6EFI/qjkx/K3jwc6
2ogDtR490TpkhifEAf9GSjIDtbo7GvK+tNZ11Gw+DYQPHJAwBhj5lNSNULapLoaZJcK1eysH1M/t
Xs/XoD+BKTm7yvqXRlao4/WhM2dxN6IVW9UI8Ut82Li9nb7/+CECrgWqh5WPubjWfqFRsT9Nh72U
My8WrkZGxdU+XsjVPuS383Y0MZj0xblvWWcIhStohSXr8+2oraluM2CNcwhfuPG02LPbavvcr7lc
/h9CnPsE65P3PRn6zlcjw6/BOiGXfe7YBRS4yBT+ivceCb7PnyUaceKZjY0Fxq1KCm0fsNwRGD9w
LkRUrlzFi/s1sfObcKBGLSzXp5rA4mFoQBe4pruT52DRGBp6RRiocSRFaNuypYJAqOWiERBJIb8f
HTJuHbhU00yskedUuYlQJEHTQk5yptUifbubUOLXRHkyUAo9fEVRBTQd8SDm3BuTBKKta3qQdjQu
04WM2iCMdG+acI/X0AELmbU12+yeCQsMgLVGtgR9xzzF0jUiKN8jFCkisasneYGKmaQDNBO6QoOT
q/Uwxr9azxRMSbcG7exQuhNGKb0E2OyIVRv3u4s3RBFzbcetdeDtoRghh1pbvpT0192eXAw55eol
oNxyna6lbCoROHWKC7o2CZufJzN49VMk7SQdz5G1ctvoxuYNE+xe6JGGdahnQl+GclL/nLdKCmHU
OqZSDHYvPTQs1wOAPXrAS0WspsN5P1QtZZnsgsC8bz0ByRHxD4mZVH0ERhDXwtg/loKRxOhkstv/
svDhFgNaJRF3IHGxxNz61CEbu2x2TFIgMoYH24ge7VclYTE+Fc5LbMIuMYafcXckocGM4a4rmKDv
TP1TsBCWNMG9rWWPOaixKQTj/4PgnTVCJpupiivLNbFC9ukYEY+d0OHSmLoAnyGS5gNdNlWlS9vR
jELpiezm3LgvrVsEvFW8PeGhfmb04vjYRioRfd5hHDup3y4aHtUlVu97AvOMLD37pur5iEbq8lb7
3b9DNHwdgkkW6le0CxVkCNpEiJKN8Vr39fVM/b/oHPcyk6DpxLEyriF9vss1RtGfxOhuSNbj5PlQ
sZSnF4sTI5JYTEmyW+iNBD95T/BweUYFYEg1OJ8fL1UjDwhuHoD6kEnMJkGg60uDTqfz2yLkf0kT
wGyqXPPPcpnDi2aQa087nOv09sQ1oUkeS7m6uyOTc+HP/4dfFZg8ie33FXjEVoWruK+PXwF++YqO
jdlq5O/dAi8ckkx1T3hBdTXcrTlVjBnzrVpu/QTio85t4Sd3afmEPDWJ1vnSNceqw2L3pLs5XYju
ql3nmt+Z1udXNCvnRR5WHtTLs788NykxKT+i0QHeyS8VuiWhIVEZ2a6KfcMakz/a75mHO2zYamC3
X5JGd/VWnyPd+udxoAHs0S1ndfCFy6dmdl07TW+fDopOICYcC+YdO9DiQ9pj7udOsOjU5lUNqJUm
JN6dwoAz9ud38EAN5HPgS9OJ8clsf3gyicrW6zxSzAwwcnThsREjwE614bqLFbujoXKSGnUxDznk
KPwnfLMB7OnJBd2gPeYRXlAtAn/dH0hBr5cyiggJIW/nb+OXf6MZTVg4coCAWSBVnCD48Xyh6vMF
IwCiUfyhaOtJTqNWgYCdCqrPvmSzLJAJtz0TnDShwdKvQWU+ikUTQ9JyPl8dofRMnpMr2MgUvFFD
2casLnureV/suqEAFCKnjhiWDvMKU4y8arIUlb1YS6ki3T66T0yM+Nd2HHBHiSPzDhfiEH1dN1Fc
pYtBqRQs/UK/u5zi80Ct4lP5k2q8STAuZcpBv0MzF+wRAvIwJJuxCR8q5dgZwRrVV+Hvz/6k6ZKi
hVYwCwDpXokD2JoUst9rNZk3Aud7jGJ1GhZbmN7bI9t8RqWPoRRweks+PXiCcUW+Ifsr0lNTx6tc
tfmD9a/yeXZEsbAR3sJToroOLseduEZuOU8Q53uv8FZNUVOOvet9z5TlHRDKQuSYIotCN0Bh+mFR
bDVRewEvFLlDQWDlGS5fnlA615DijnjJrjMZxQo7Ob2Q41yp3Lz/8Zjn/6YWU1YRfrj/v2PiRTQG
SXl0EIel8zdllCt9Hy0lMzaqm7O8AGL7yEmEzoeIG6XJN8cAaZOgiSrJu5JV/ZzH47yNMyUhK4we
nmH26mBMPz6zkxi1EkUNDkaKCBy5jUkT9DCWzK1wgU49S/uWFp4/HThzWysvAzml+/3lBslXnGm4
fMLGlCSn0rthAtwjgYITf3HfeLPvv0cO3nwrD2wN5J7HkLkFsPFcLnr9PVLg7Xb5kfvTlhS6WJIK
YsBIDVddPBwHA507UNMExtoWe+QgIVD3bVSX7XUBf+K12I276ylH41Lrvzs46+0eEhDM+GAenfHK
jKr7h8VObG4a8Ga7jeVRl5jjbSELH3d6uKOQfJl1zeO/zIeo4PTkNOnM3NFHTMjQ1J92vHCLjEsP
Bkir8ecZIyyu5IC3BH3YJ5vQ9yE1CLoUpHo7qjHPCSPwEVQZlAh0tYt+OS8RAAcPY+NVe2jwrk0u
cbXZ5z1g+xiQ0rgqSYnQObQmVcdHUd52cRkZCPbE5meSEi5au9+pGf0iR/6f/tX4vjl1YNjTwREW
8XIoIwbsmNJIpP4gankcQGeoKaS8s1dQryz1TAyuRqcRzo18VTeufIaK3Gnzv0vW/eE6LbdDbIIN
E/i/yFNOJ+8nbLxBLf30TQ28LzUr+bFTlJELtJUvRkk4RPGaKwW8I+niDGr3VxynLPkyJJMmFDak
sLvW3iTD9XhN28rlGyCUUjVclUqH0nts5NsZ9EgyAaGVA5rW/DlUyuzw/B9SBDBJCypHCjr9xRms
PmCXx9xAIVDLjHH44QUq6srpye1b7UNMqrO8hLgkzfUJ/IFzHjI9gM8xFgeLadqFkM9Ztrf17akE
Qm5gYwwbc0AAPbZ3ehddA6HQdqiSaQjgENbl8DnNK1iJ65iuzzaunf+gnmTHNpAXky7vC1bfY4gL
yPN8hVb22tHdTMucSfElNTAWLYLgiUBEn/GzriarUj6wCoPN2aeogYpmoEljZhUDmQMksy2lskyx
xm9pSj6qe7HN4Da+kgS/voRdEpXzUIA0xZ/uhuxb6X5A8jMVkuTLypB8enakgy88dDy8yGxQl3aK
/cBYR55r8US6edu2B4pAcIKrAqJeU6rDVSgOXE2tRSz0ozxalAdRbxEfiqQupiz+dDF8ni2my51c
px+zX/ikTDzhbQUtSnNc35EG21P7ZeuGnP/kWT43qh38s2h21jRrlJOvZ+DzxVccmOHUcrVOzd/4
c+Yx3RirDkFKBiRPHPgINklK0J/n71KN6HfvKqcbKxIVP9wFcvXC8iy9E63q8nZSIfDbHKfMdru+
fCVHeLudpIuNx3LI4iqzpWJI7DSZNfc65+I8DozuwFw6M7/R3hIEbjyHdaD1gR9Ip0Pfz63eiwIa
XgDDWWGcfFDhl5COhNtsIaBcWuPFV2JBeL+n25vTL6x4oKkbkVQjuowJlrJhMQuKjo8W2R4PPfyZ
fBmj60t+oJr55hueWtMBoSefV4ZwNIWuUx0/r2OimumBQhURQiNOA+4XPVzmL22lRE90LIbLhE81
uGKEURRWmpiKg15MCClvNunHzgtOgRGVgJbcPOR2BQG7XQCfoTQsFKnKspC16KdcpjCZEvCV2Drg
uoy9dAEC3S7ZCDELd731xrrWmEn7nWIwjHM89UW2V+OXZZfFwM5Kz2i7e+3xrKK3FG4/0Hn1yAAS
YYiaBzYSUgBLSO1We+6cNwNc1Led7bWATegY3Rad2Vs9gPGvBgdhGTg9nuqQR2eeg9xxO+kzCRmU
nfQsMhavHPIw8mmqXIFi8dPWzMw7SEYHCklqz2rMY77JOe7vZJF/Q/LPJJUOpxMzXn8l3+Uy2/mZ
tmfy0H+Lwrf8ePh3KgUPXnJ2mmqk3Q2EeZ6MTbEUeAd7QJP8empUDWnz8clZEzJatQwiUG847upr
3fV80SXKmF0Lw1yH9vD8OjCookt5CJHRT7V4EVk5Mfs0EYnJA4HdS9j4i284YWTxDoUl2FnC4wMZ
0fosMBXFHW2RmMOnCGJkxRUHsVZcvJzAiyxBzSLZ8t9teHDoY7wSDJCCSs4ni6WUxSWBE/bQC6RX
1OFzTC5KUGoDx6zcqUPGaio9vfUkjYXJNZ5OZ1s9Rq/xICeK1yLy5hwTNPsVSKIOPXjpBuX/9H5T
KO19SBR7P3I3asnB4AtvtREBjLq0Q6VB9C5RN776lFQGRpOqLu5Z/fzwwI+cLXJ/4+EDUX8T/cVX
hB/Z49fMnMXqJZRn9gxInPwJli9b2Yxr9q3sz2nfyeBw2ny4gf5NvaRyRqlLoBRGBhvhdYA+eP6k
17RkZ6xsE/3THp0vkE0CndfLZc4pqbgllQkLsnbQPP0PaBfPbL33p8koJisa3AuxyPgAf+fCQB8c
niQ3Ozj3Vo9J1AyZyobb0aUwiouUbK/LJ+9slZ6vze2cmyyImJIbyy7Nauclf50jvsrZnuJ07Ree
MwASDgeuKPwjcmBsOVn7eyikQIwLDiFffY3V90eeUKTgpear98o83OXB1/WOBmuHVD71GkCeNVht
obE7PcHe3BxY2rxJo0oevkhy9RzggP+LPqneXSZXKQjuO1ruyiE8B6feTkGMROFoqdGQL2PtqVd1
cDjsPe4V5Yh0fUuTKASum+ANAowRbYgtk8fxDAwGiBshsAFi/XAqN5F1lJ/mQ3dEmADSLZGH1gDD
7TyJchzWBYkYo4FiqsgDbiuiZcBF9sYYfWQUWihux4fXn6Pe2gWQaKfwNp6PxCr5BvwRmsCEOfhR
/HWAxlV2yEyfo+Hs5V+cfOEXGGpI3SAGELiSbD9S7ImwDlvFZaxeQCH86h3TpR+e24gQhrMzriqK
VFU/n5DryPWUzmpDklS0JDF1dCXxVXIVOdf+V7S0yl2u1gCvhYK60yOEiYOA8KRf2TkcCF8q3EoD
Z4EhNqQDkKXhnYGKeEVTHKHasSMJXj4vtC0gAM7GaB5FDViszPGUDkIDRNSo6JOEMxSqOjc0E/c8
q2MZxM/nKMFdcbSR89OBKRZf9fZTEZnaPpS1gHqFO/myPELyVMggWDlGnZ8EDjVWN4euz8zXeDae
1ubIAkArLTtAOmQOhGTCc/kn209rTuovnDrztK9zbjCwOOjSR5cFSJE/tyTxqYm00XY3T25FqRlz
BHv7UFiF2HwJUByGtv1ElPKsVEdnvoZF4vPmjUdGztYUwJMkGxcKn1jEqJgb8/AZy33I75xMq31o
f9NeQX+DtBjDtz4T+DB85I7ErX256HBWRVriDMR2o7LFjvnGrhBjEPYjeLgJMgy29IxNheyCjBkh
ozz2vI9UW37JNMuHyiwrnWIl6bYctzFCxKwZtatpsr9fTgewKEWj19lRn5Zpn/pB2IRzWanDwbKl
b45w9RnIteJ3dEKwHUx5t691GKM9uBQ2RyucaLBo9mWeE+EsP4OhqQ7kxA/mt1M21HAalGBSEswo
REoCY59S9DRTsH6wlrKbQXUP9J3pMrhUECIommIG+WMpbs9+Svuiw9+bewEPpK8RHGMyC1NazkbL
ByljE69mikkUf0COuMKmdUbHapPv7zRPvRsXZI93VJ+lewIShG4dNJ5Egd7RkUk45TI1EFk5N96Y
yNPrRTaks/XOb+QXKHnFqTVKf2LYD/Uyoeois+QZB1t2bCPRE/PvWoHTc56dAl0z7nlRSYrPMzjc
J5cuo8bTZc08L0XZeCk20zxvnTCIuYenFVXuW9z9Xw9tMkgu2eo+zj4FQtTLxBNT9fLVwrx9VvJm
ZUydBcQykENlJbn1gq4wt3qyEZXZXJIAkS/8fgS4ZTIxdxqMR7Vw0GVoHfAgglc29cZk5VaSYpU1
K73uwj29ElB5PdtCv/45e3vQE0a9t8C8K9lpk0R/bpy1mLahdbBFDFi0fHgmsrJTRoh0Qd1Qb8Fi
NZlCWbg2uRm3cb0cPsCboCxhPX55S+AzXBbWY/fdDL305cNdvvkEa4V+PhRywsdUFPxm+ZhbR0GV
6e4z1RHAIbpeh0OFplTFswyRPc/6fiw8dE71WCEKc/xA/E2Wmk8edCEW5j+hX1535EO98SgbYSAX
P0X2ZFHI5SspqgdVli+Cm/C0Pd6wqvFPDeTDMCqlQ6bbsHwDIJRCQV0mVrHg2nco9ZrS1BCOguWJ
cXyJb0hk6DJAAMsEKNl6wnc7Q8TKjnuj0pL/wRwFz0I3p3TtfwCHEWxRwcPJbExcNEiqgqJdjH7L
H+zQuQiWVpplj44+uYoeGiq2gyPnaSlLqeZpdQlqF2SJXe9LPpPhlfUHQxwtWotu2GT0W3/X1+yW
CAens1sFGy5lFE0WsyLDwsJR1zBUJhPLPoi2BTW93WKc590Bj6wCYQQVipBkkCrTshqkOp8OI7m8
cryoSCHEFvLqgJjXJ3yxnlI7CZuL97thV7A/unCRtpKBzunOtZKCH1V6LgxVZcnp6WCTBpVMxOHr
78BbHZ5z458kL96Gefwe6tfeSjRcvKI+RWHtTwVI7fT+U6TJEzs15E8sGkI5QmA7bSu8QEqCosyf
mYulZnQQZeBU8xz7ozj2beS6nrWTYi6W6JJ9emd4TNj5WYLcQkZBTgH7RdwxXNiT7GPCsPoGi8x3
kZzxraSF1so/Whzhjir4PRRevnXODI0PXcyqLNWwAaGTtPG5kGBzMVuOepa3GvmDJimJCvqwoBl5
Q1Zbx1K5PIiS113ZhKBci0POFyGbEzRC7vGkqooyAEzidE8zj8u9RpDyT6pnq5ZJG0ZMsWAxWYVA
3UqBinj/TyIavumu16Moqz83DczncZZ97XcmwXYNyaZaBr/Z5Zn97oh8BKBS6RKoq4f51+oyMCNs
cVnSSgip/Vgji54+Oibwm3wQkLvF2knboOebzqUTno/tocE4cWyLVYrEHgtEBiUgWR0ulzwEsLuy
i+XQxn/N5hpDzj04KrqlCfNKf7Jkblxw+EhjKaJWnDsXkdtu0HPe+Ty2bqzyZAK5Hx+QPB/1Dxr4
O6OkRpn/KXUyAJMHvHWr1YDaHkKdYiPhuhXKXKBAVLQj1P/Ijugl9/FqXrJAldnSYNczEVyH0ZnX
Wsgu14Mqcttjs29X8nCvxJogUKOUf6uXXj5/dAFbAozdhUZYCWX1pwgQVLx/gJIFYqdFzeclCMcC
5eAx5N5Dp8lieh5AZ/PxHI50cfm0jXsUAV4/cdRT6fujA0rd2TcZ7DS3LOvlHWTRy93ZhneRppJp
tNFl/POUvOzy8FErNmprrt4VNFoK8qwS9xNmqXntEvXg3N5+aPDbKtGoRt1Lq6E9bgYtuqXYZu8O
rUJbVN3HClQA6z3r6opJoQCYl/263IiPJt8/uzdNph2fl3bMC+5F6GtmarqYL1kWkjGajRIz08cs
XtuKRBfYNhg6454t94/WMRz83n4oDLHEhTOaGGVNvpCygUocQ6XMHMJnYi0Xu+HbYObh4nsmSZ1U
jnzGLBLwNYfL+P8XQ4ZywRLdDOmdjhaxW/ODYJrTjiJ3VVx6ms2yZCUjZhYnQ5wtMuaaDmWlvK4B
HGAdlXVe9F2IXZI7i937Ub3aqZvICZKAS/O61La3rt0yNTOekE+DyqTDWx0ryFKelyxgF6nu0++y
YV8iqNBNExUtcMZziu6z3VoDTgzCMzkxFK0Tjc0ToorIgwiMh/FNzmQQqoxVozYA2KduEizcVtGz
hdmSNfuwURC7NLlfFL5wLIubETlKkDu5UM7goBPTeyfdL9ijRlCMWfOKP7l67t7YmqjxJmzO6Gi5
q3ezeCEwZQ4/7TTgM/GXWUwEgeyLhDykOYrRL9oalBPBqAhg9XBf6UJiXyFyBH2W501+uHDBR9gX
HEuzuzSwkousxlG+ModciU9UzBiN4NMyDKOm8xWOOym5OxtF9Aut1+yO4KJr/IZSUGL/t5Lx8rtC
jh5Me2kYYDfmAXPlL3ztWqSfzX/iliy3o1uKBzT4Ppg//V/2SF+ZXz1bYdwgeIWixU5gsR9qn/PG
6BlzqrlTa1OQJXnBnx2MWRLaDVcI5TUCEPrLO7XCJqsfWDhlmvwdgUru6rTkSqT1PQM6h0mzpEQm
CHVNJb06Uoq4VA0dKV6a7Yp4bIVPqFWqnXAhcMbDWBuyfrYpluO2ngyNjYZmOx0ZVb6rQzK/0Udk
EV9Zcls8E5k2Is/qgVq1m9EumSE8SnFa4zS3Yf9lbziyUq7co0q+d1ZZNc/9kqrBnzGVtCeTuhlz
98MqkCsg3vYsTtnzHC41NV7GTit/Xl6qE+89kk4jSTAjFcu0fJ55XgplaDokHNTyZbmv86b9mrP3
s2ygQiHTJnEZX2CDb+Y5EhhG9POMmtT8pyFr7meH7E+34/kZ7Y3f/4vsLWz1XKMVvBsmQ0Sy+GnA
cmSbrcmor33J6S5qZxuzE/I+UuyfnMxhfyKr44sTbKl4v1rTu+hE0gret+fG7offMksQAfU7TNqv
dYfR68yNFBvgZfCYx9tVyA4+BmB5CMBE5cX8sGFbwycshBHIKrXo7IlULS2THQoWOoBvdQoXQwvY
g9xBDkdmoCjWYglMvzKFbr+5YHqrLZbs6WMTEtNiDBuA/sYYmzXMjMcDoo3apMlBl2hnRIAqya7A
KVm1qu5EjQulHlFMl64OIBnvBZBaZIov/os1W80p69/GLE+04J/Ahq1Zz7EHm6bWil/5H7YmQtmJ
vznHXkiLuiWrb3v2cMlzSIzU2Y7s79qi+HBNLsp0u37uv3rquxHhUsplSZ+HfbFZkPQI0lGqL+yq
u6AB9CoG0nRf4Hjw36yOH83Cn6gT4GPCeI+gla+7zrMEf3PGr6+sYJnj3mKCW23YDQbvfRLWDIj+
U6CQQlXgaGu8qdnFnqscdqF7t27SqvcNfc3ybBmQrK7Pco3MCLRuzTYs44FSh2jUELOVgCfygidD
+MRUZHRg2JlTB4IWXye/ccgJrzEFPkZZ2HoyQysHE/ftKNtL2vtpkdt1AEHLiZEVIsYtA/vrZyI3
6UxgQWgMFq2A2lkv2vpXOl/yRp/N+w4pNbT5JyNG4NsDXdbaTIw4EeTav9t40LgoFpVYe6eD1YtS
a1zEtmYs+ebsGTaWy9WUjIDv5N+g8h2/DmJ7aW50LE9rBKp+uhiEOggck6gPJ+C7qr6nYOO8S5iL
IKhn+2lm/i8c8skpJIlw2+mDj9WL6xy9WDDkkIkePXQ+SvJOHIVt+mcQeYB9nFp06QRLydVMV8jV
Hs6fDj1HjUKGm82GbszBg2RyTK7aBHzWcLs63fLEaj2JldUaNTt1n0zYfazusDvxJ9J+gxx1J7rB
SKfIaQmHO/Cy2ubR/GMi8elXY2xzxJqYEXrlrqjE42p+QgMu0JIdjJ8vKdxK75JP14tgaJI+PV9N
RA1fYbSEv+JFyys16/cywoQfdygnIRDK/5KQFt1QUYDSZ9wFMixXmopzoO7m92qZ8mvPpnJMq6BP
p76n9aHz5t4CiXkrOA4QwyHWOl9BpRMeyPBK6sCQcWuiwoD/uwAZH/p2jCri6xMM3FXgYMSfAe7K
WqXSlbBCrsOeOEf2ZWL86QW8bYVbAFV38yDWHFfosL6RhMjpTxaMFacEpSi5/PrK7xMHaZHY+YYK
E1SOZB4zl6ge3GnEeNIbINxadp913ayA3iHxcCGty5i3PTJD9N2QQGqE+SROwoAr/ukg3y7INPNx
bqjLveTxSY8/qjCQO0gHFT3tVLcGxJBfhULHf5Y41S29Vc8V5N4bLT3P+MymejLF8YcklO74fVhQ
nwgKyztEfQatTYdJl6A8MoD8UmaVPDT1P5lmbzBHiJrbZBRVo+QPQEalxsqUMe1pF4hE98kmIVtu
uAfRWy7jlidJn181vVWz4PiCARRiouA8JXjQz4EFeQ25dnURnnL9lR9um2Gc1njMEuz3GrEyCVTa
PTSWYlDEyp/BujN/AbQnleMmIlfIpZIlpA3JDMPJ6HlJfySd18cEfe0NV0fRm9o+8aCfxaI1n3w/
UblbtM8UvL7TvoFBOPhglkiMfJ8/sK/zFub3zCH5ZiQ9j+/LwZWfGHAkHyIwyGGLawqUS9VpNAt5
ILKNQHv2fLjOM5A+zV3davEUdiCFqHMdYQ2rSOGm2s3u9zzJESXRrFpcD/lUdrixP26V4rG19ePs
6Kt/g0uAZwgODe5YEOLXUo0QTue0fmmkzjZzSJY0JY8dDosKYM004o6O8Yy6l/3oELvw5WcOixaT
9E342epgKtE0b8kI+IyuKEOiT3WzIEWkNdlOFu7l0V8d6hXMBDFyBmsImJrd6xu10b3JfbFh9LZa
iiTwPWL3PU4da8tt3ND4K8F3YG+gr7teZikFy73kd/Kva6symzim4CBVoXj6tHlcGN9mKQ38X3sM
yOxEPEIZkpzQoDFxr1dhHtzZnVSOtFcur6UUQexSlH6UruLFoPCRMnpJMh2bg+OuH4GAygKoJtQo
26ZIQDrXdrwh/9irjPockG75aunU13PV/ynKeeGeaSDmQZAr/hUz+beW/Tda8HuHy1TqPgw/yN2Y
iANOh18e1un2cr6ASge9OC2XFoYHEpfgFbtxlj/Z2OULh3e8UFn0wl8dXE+MzNM37Izc5AdxKf/c
ovtMx1xSQBsmec9t6MaMfwtHF3NpXj5RhGB9e4mdb1rd2FFua2rhIkpRcf+XwMIpngr5kyWcshPs
O1WsScwxgR3X6iQCkYLrWthR1HDDoO4QaTrAWR+OX89iHSwCm/EaOtq84ZDE0GgatF3Nd6nqB+D0
/4OyD62y4kz6GEGMKyME8/XB60RFnJeMlR2SV4B7wtuKjl8VC2K9IVJenMk4y+K8iWHmIOs3ubvm
vAcnBZ+FT0t3ZVr/by0gHsYG+Dt7/3NtgrTswordH0WfDfmVeTtrj4B+aRrJ210YE5j2kAiciDHq
9MOp03HIVoqi7dEiHGWYASGW/2Si7shhDkZSto9W8yhzggHOz7Zq06fVFEOq/lMTNDz/uDucD6yL
dyq8VuxZ0hhrlmC4F+2AgSuPRrTGRBW+qSZxx0olr4zOKzuM+09hxM3mZHeRuChh35p4T0LV3cBk
ZxoXm3A9F0c5Oufhgqqpoz4F8lpORnFyS2gfrcjyVbVLTBDzyRalwhrdOwxY6UQ3WyNyTGyN894d
o21SX57KdRQx/EIiYY6/W9UjQ8XYv7Jr+fBGOtoTVeSkz4HhkVjKRD6AC5DQSPSrZl0EbTyZ42e4
xMdpZU3SrvshmMuPHO6CemVTT4zCQmaN+T+Ehfv7jNGb9CrhKhiYm3geEVpb9tAlWgm532xNwjzy
h/cjEj4EHaBF+bsdM04RZGssjEGQTYUF+NjaO0g9mF8WVzcmVLY7PmrzCDQrY6K9KQx+SwOuLb2W
7vDTnqsuG7z614Q0mJlB9mnVYUbPUbikxZ6hR031aupHJGsd7d1nQ+zFevxynk2rpv+g5x5c/qzM
J0UgzI8Vm0KUfeyt2RuLIzlyVLfvkobfPrN8USgvmFGQt4KfYKIugCwN2wF8HNjV3sbAweEqquWv
MxZg7bt0nK1lxlqNwa3W8PGdrliqDI9rXex1Pin2T/Cazn3TWtus3nRfOqBWYPX4i/DyDGoNE+LU
IPUCkOc4QufKxQmKglkpGJx6oonOYRN33RUlXE2zXawxLmo3FBr78ztitg31GQ6p1ZcErVITv+wK
CIORefpHagRDptlBR9gxOsDwsE2E4jfps1/m81BFb+vN5HyUxaPovBSGFyCp7CcAqUgE+eNldH+c
BeZPwDPxmzeJr2WNKUxt47SNT2p40QJ1y5u0KhGXD1APFryqqRjytgEuPd6doLhlcyyFsqOqp7VF
ki+L+qwPweGoWkYbDPo0+QG+cfemt+aPbygZD/EIBK6ttCmo3hQr7qLyYj8BvZNuv+UW2UOhPswc
PSB6hr/SYw2FsO2+adYesqANQUuh2abUcj6sY5duacL+oSWIgG08Bu98NMK8x6x/y1NNpq/X9uz7
hc8qrk0DkfztGOUPJKsGEtlO93B5t5hJPdSNv+L8g9LwrQ6/E2EYVLCHi19W6/0QwIS4rHlIwb7T
3pEfOCG1B3K3wKEi3isG+wJ7ldlTLsUbj41ugJ/8V1Hz3CGaZbMrh2/D9nhHEiC8EHiOFAYB9ct3
ObU/7me2kgoupJqnqfYLX7i02lOCp23rQIT/wbrtW3+XKfn4lgnJqTuYlttIlChsRXMmBRZ8dQHR
iPRtEJf6QFyscEwqZ6BYTprMi6Le8/SNdm34xe/vWGeGJ9PWJsjVOqaLogdStdywLIaHW7iacZlb
PybONTRw0g5NVL6fOLGGV+RTooT4QpxjeEfht/Qt96HSn0reEI3NIYMPPYwaF+adqVbTtCKv44Xp
ocZdPL2SYnP+1TrCTDnj96LFM+JjhzNVvgJ/aN1/LuQVScU4LAb8b7hz1Q5zhueskgKmQblUakrR
xYSnP3KLaI6eykbATx84G95/p0+PDctxvLT3/LRkIaFSnI3fDiV/lQPDpZZNEbm9eP6FmsI3H2ln
l4MJl3oqoR8dmvoB6rQdRCEQRJYmrCbb2BTkLB0VvZ9BEppKZ0cXR6mYyGKuwKVYWercdMKODKmj
Jnae6yXTSOE/maz+oNn0+CioiVc6+MOLR9/kOutQRNoK7K1hNt2wEJmk6dtJORGR56hOCSJKbvQB
cHiW7SUtF/9re8Kd52CyKmSJSWgeP0u1u+tH6sQqIFoogg1wFXrCYOXz+R/G/P7ZaoJQlZNekzBw
SuqL4qEu4KfvsAF259GjbYqtuImXTf6NX37sk3xPjaP/KZrUdVQ0KFec9F3Rmyn2AzaDmXg57SKC
zYqomvZISvR5Qd/ciL7iLKU3ow+iZhQMII/3UpUvPD8tsUpd92TUAIagCzT4n9hVhIOfebveAPFS
8g9UwTIVymheeGdCe11cJqF5XpJCifGQgKemsDL8u8Gk5lhhbznlJtWjlKW75PXju05Z8nmuxsGu
+0OElLjfGsLUdF64ThHx80DFuU0NOHFyv5wGDwwVI1VIbunjBdRdGKY2Rh8oZLHKRmlkUiyuca+P
QPv8Qyz6o1EilGhKnFmiu0Sl1aO6W+PrfkmiCF4WiltQpIwqbW/IQhVqK4OeXMoY6lv3HeuEYeV2
kSpKrwjCcN6lqmDp+pEX7nM3P4dxrbIdawQyVk+6w3QsDW99CrdWeHRSJLS+Cmk/99ibFlerGPtr
27wfM16I4GIK548wvi3PyFwBOtvpzan9GPnDPeu7sVnu0vHR+M54BR0W4WPsg7PHejsPcmp66cr9
GK/6WYWftLJRE0HnXAVXSRlXFPbTQfm80GGlBaDT/91efzGhk97YPRHOvS8OftfA/mh3BGIq9wIP
BmgM7DEilENZhgIw0ldYxL5QPp+VqE1b4JzHMUy/91D7/r3MRskFnNqQed9hXBIoZorYSbdHz6yc
QkMLnA579k24PLyHfb3I+RaKcv1OvyfI8qLN9emD7yVSftI6N42l7ALLiT1DHJK3jvj/sgeDmFHC
fmN8oRl29br0kKcY2pHFMyq/8J/mQ/iaw4i5cAbFMB9nqVKxpP4h7jsg0LsHeDw2bWoVSZ8I5NNu
84aftCI4flsa2hPpcvR7Pb8sC38kbLFkg3muJcLyi3m3FfePsDgdFnVkY1i0OCdLUio5xNnwW5nW
qDDmTn8OfO862UlCvzhvlylZuPcsJ9mquRtUUJ7/X3+fhPMPzOaO5LqzoBj5pyc9BDX0unL008Bm
0EgkH/zahZpL+2UXbPtqzBiBN54Hsj4bROngJhdeJRHwlqvPfcVwkU4L8N1+9liUihjzPd7TKP8e
HnqgF2/BAm1C/Dfex7FX7jtOKDLheMKZDnMXoIu+W3RFHtoXKdWy4NaZmtYSFXvAeJtSvQtRCTx2
PyRnxnNgThI0Qbiafnjz8c0GKBaHwNXpeVIyQZioE1y8rm/1306fbD24o7cO1zub9qxSpYXsLvfG
FU4JRF63ImuE9QrNTtISP6FasfqBk08LZr7aF2ko6c6EXed/w8PiZ54klyVbPADYAoHaF87DfVRX
TG44nCx3UpX8pJk0ZM4ulv8Jdh9IA1jVFza27NTv2Y7T2rHui1jw33KvZaxdV6oKoXlcDM2CEdt8
A4urP8VkVVa87PcC/IgHyH4fzDdUBSf8ec4661kcHpwIk0/FUOivkxwb1/QA6xyUmKJfbV/yk+EN
rt6XfHTaaBlqzSZb9aUAwspUGXz7c/IWTF4X8QBiZcs35NhsAGtcnwYR/KW30ayf6/w/WHwLyGxc
cQ5aWRLG3fwcMAG4LOjthLz90IEsazPnEIsKLB7EbjTouXxGyuB99Xfpxv7jrpIhq43mMmb0yWoB
epRCyOjeRj7/QZZwDIvA5yqUNYLqWFgEPI9A565+Nyb6KuaswrJQcqmoum1Z/+IOrwB7Ad753pBY
yhi0fU2Z9u004EaoZvIX6VgjtLU13m7CBG+zDmS3kG4Q632TlMIpVkj4RyICjGOW+TYsyxbXoNK+
AVQtgWzA1VgsP4al91zPyEKahRkBaDkhHTgBGKHdTFsetA6+4uPMBx9smVNlGmLTqAAj1Ybwr8y8
xTBXjQh5mxdEhX45wb4J0mK4URq5ALFqIb4QowxsBzus+24/dNRg1Xj5BcGL5y79TG7bJd8XfJsM
Y2PEocxQIIwdWizgDDGk9oqKJyNpw1waXk7yYehzgw3nf7lX/gPInpiQ2/56IdyQYzfpKOeAiImD
X/kYx3ZoS8plyGCYPqdgYfxdwx8Qs+eGQfCcu5sYT4eRLsv9IYQOCoLochFxnJjDfjnSIHSnPsVY
sqLyDPvG1UuasbhYjY1GzUA1NLtkAeoOERJzXu1xqrpPASXWIr/+WDXWBCI+JDAzWQrZL+wjt6fa
AhPTjwHDnB3Vr9ZkWb+R6VwSKQwxsWAZ+KaEH1+i6XfwnyIctHUoWy5GYgb22CEr6dAgErmQdfit
MjoLF3dae3n+lyEZKVkpF0vXRysPsANk3eglFSpTXyL0n2RmvUf9kSZQAr+hNytn/QmpwndzZeRl
akjP0GHy5uNE27pGpUhqAAv2fnCYv/Gwg/f8S2MxSN5VH9dl/KA8lNHxFHiOY8vuKGeQ2oqlCNl6
mU/QMDYETtmnVWRAu9YTm6YXFpk0zmT+lhocPXTvko3WpkP3l8R1gnLSIW1q/a7oIxSAR4Nn/3j1
3g0hYFTe0XYfWeSNZAnb+6p0kfOE8gdbyMiQOgSUeSiZXC+VLkxooX4EHC5LydiCRQY9bU6BPPh1
EYAF9QRYqpSnwNShAyeWFiP1P/UTDcosq5jqqRYE1Aqd66EVayLEfgP0POsmMvxB9KjYIjg/+URm
TbGmvqaKx2ri61YIE9oRYbqLCRG5EX/ByEqzrgYrv4Er3wnMrf8aN7END+K0mkzsLfp3T+TD6L2z
GrhV6AO7lPBpyQ8K1u1UT3aQdHIvwwb8JKtZlDZGCCFIBGGxfwN4sBHU652pzVHsme3lVwUVuqHd
v6dSrAdAzVNFUWh6sCCc+cs44apXKdzZ6Ed8JHd6Q9UZ0TaCcYqKbF3d6Peynl13jU698SIVfPyQ
rt2kAeKhqLLzba7hGHyTvcU+jorVFmNcW1U4fYouQg28b9MxuxoJrPEJjvrdqlQzQmeeW6SRIbhP
kZEGw8cKV+MQE2O8qSUIl6KuM3q7YLhBgChJBVDVoRjMfm2acKJpqgnRVul13k7Y9oshRP8adP/W
sKNxbgs4EOBWSb3xU/kBPAu7KUmrBbkbAfA4ZYGnwQ9LFCfrG6Z5dCTQGNSGlU1rFnDRQ1X5BEJx
R+OjuhbJ1pwUi6F/RQt+D1U+0SOifB05CF70h3dsqS/QakmRGSL/cJihJnyixrhVUAAlNavsKjKG
A3Eo1xnqcNY61hXE3bn0XEe/ZSLtg4it/UxthQjGZI3nXYtGLK6N+jC8QVnDxfmziCwkR9LcubFf
fRv1GdLMGDhmM+gUbxS13/I1m+0w1x+Dd1lUpfIdvIbLEv55fJHPXZKbSMImwYiqejTD3fWP4GFS
dtFeI/kSe0Kl2MQUerYLDxDgo7WWVr38roGIiDZl2NioghGV+lNpgRYPzVndsSno96u0sAOFBrvX
I+Tg3E1uXmSPHmlnJts4GwHUomN93dNPnC6RyvWNeWSINJt9Afl+5p1IigQ33riWFIapbH99SDWh
JdXNa/4ihavxlKB0kTN3OcAYhQ1FQkOk+IqTMSbG+v9J3A2+9bf9WAHUlHV0ooMwLco1YvJCaI7A
i9lgGB+e3zO0MAjUcYFNJchevd/17AQUbqTIAxHPXk2DIJxM7Bua45gomJeqqzR6CgLta1bMvzsq
DHxStd/AJVCyIUD7Lk9yK1WBh7bmtNjoGXUrT9WihQYIUS89BjLzJJ0+UjJS87LEp2eqlB/Yuajz
v//gfnVI1uvs8tKPatzgWd8lzjcKFaUiQ1G7i2RHgV4ayNl5NVuimNv7sQsS3+A+iAv29qpGBJsF
vsOAAOGrbjoVBs9DLTZw+EfH3QIfjcDy3pDLo7DR2SjJxm+WsH0fp3LEtxx4ZP7vn9maasZbOguE
+Y5KPPJ+PSrD3vgZ9sfR5p7VSF3x/WQbXXRCikgNG+2FkWfz/SEbI+QkksMY512MmJIp3KTFu9VT
kF/JCtiHrP7NETI98BsNK9/lyJppWTma7X1W25vxwhGhPCKLzIyTwkx/2C+3FRtiq7nrE/qSVUL9
u3mM0fdYzNsk0CftcjsvMCIWgjjprBCKW4gcPQYJTYF5+k5DXvZ4KQev3Qs3R4RYEpa7cF0U23ov
z8ZXKiKQRnZIrGYE+7vDL/Z9/iesrorn+6M2tjMVUcTPYFcfvo8J3Z6estJsR1Blo8AdjnAryYui
iBjZsVTB0oBeq75Bz5qb6JxjWAUoUuGNEojto/4gocjQGrTvxplEEd4WVpLSTGueWkt4t7xaDIA6
FfJ25264LEPqEjSd4lq4xXIBb0y5lmEtTweyp4iPgZ88NSIjZz3WXXqOd8NWtPrzlcD2CrgM65VR
LT3wkcWde7iUeDrgS7yKEF755yEJQ2+LEkVHCyz+ApYT+JiRzggYnP+SuHYbBapxPjyTFZLxvj2f
I16tVn6hWORaN311wUTFErQoMGDimV4WIvigBDwrXN1Bfz8sRqsowgKmcg63B/h1hXCpr2zL8sr0
CxycnzqWaSBh5Su00GnfiW9kiiWjS616/JU5eN3oG3TmN97HEE4kDOJKEztNWJF/7nGOKfRNvBco
EcQdsW5ep3eyTBhbJo7VuCMzuboJ/TNvI5mDvW8jywRgYvxklhNlC/q5X3UMfy/+i+Cb5M7dtLRt
sE8ao7m9FdRyYfzRH7M3qelhr9iBnTClvALvNLZBupu1NpsNZP9rXuhcU61DKZglA2vvKCHF7Uea
wtjVWNjKmZualaeZaRN4J2K+j0KPwap5SpVNmBgJilwdX/C8qRIfjBe3niF6ruHk4ko8yQyxhufr
Ay8MA9xiUkQVUuxW8NERKu+J/+r477I0Q+6UJolvLE9koo6E+gjbd3V/72D9cSvq0Ska0bTaoADE
DUL5wceW21tmZTlMfYaoNlRUonpoELeJJZC7OhHCoddMP/GXYAab197nbpVhyKdXC3y+uFcw0qNR
NF8N+H2z7dKFXs32KSTjlvF8j0D5lmmWGEE8A9obo4MhwqaNlI1f/AYPVxt6Jh1riV2wRmASDECn
Dd0mvKl1cRXf2xjVZ7W8xV7CBLV/Py2iYFfeSbxCLtjdVAl3efL9GJPZK+jVvCxAP9mVq6tX9tV7
hi2WgkGIwnX3FUR5YuJyyAousObdzDARSEfEyBoLNeqqaefsPsUtZI0Ki54knDLI10Lyb9rgEZJ4
p+72U3OvRqZd1W1cZx305aiaEaCts71gpDYz3+yrGTLzoX0nYgk8m5sBNtD9y5b2AU50mGS0kLa0
3kKNcGvZYTKgtc7Tif/nB57SuI7CIBpc0aKcF0/2GIG1awUnUxAj9Mo1JJDEu4KMhcxcUh4BwSsJ
fhaTg6VTI3zsKxXwi+ZPAYFDWTzfOfIZFIiQ96h28lHW4SdbixixpupmVIRF5R8wZ0H+DN4I4UHa
j6sDKjiP/0ggSflkquSTYo9OA324HKRtweiBJvC3lQkxc05GkQcZmgOhP6vzTYAOTi/RYpDybksY
bl0eRSRQcFUyR2gU+rSHo4QesCODnt5gvr39sqeRWJ1356OO/GcBdMvpSzB8cRrcriestS5cv57t
pLWHHFPsspdG9mY/5wwRoMOzWRHSMf4W3vM9MEG4/Nr8jpt/J4NHtOFyFC+suhMVDtZ8pJCULCxo
hb6Rp7S1PL43n9kQ9Cuy8XKdgmDSOxk+tdivCy11D7+wZjJOaRp5mBWK0l/88TSEvQyk3Ma4P30K
YsL+Bky8NiAVjanUSnhow6jspdFhIqKqPp/0oIoChAIlQ+1w4HHCPiU66AlDB2O9/nyJm/BBKS4c
4zJ0h76SISCl61RgZ6V9gGf6gWZ/J8Sfye+Z351A8Xc7XHd/Vb9cQP7RedCSrB5lbNBiQWMna0+D
KoS50ZWPn2R3RskT1fOID1JEJ6PxtfDThDWw8LHGbnWButtEWC9a1+3qrv84YjBr2ISIbicV78Pi
qQqp9yAduH9+3CeNCMRAPnrlgF4tw/c4kNMsckCJHSeK9LvuMWEPAb/F5fqkESQZ+7KcLccnASaF
PL0OZYUgYhVyNwiCI8DTaW8JHF81f9o/VfPZAoud9SGhAJuJCLV4AwL8Up8f6fx6SJeNLpskBoEs
8q4zmajOv9u9pj/GJiNlQgxFUDBXIlxH79X+Z69TJuH0yoZS/0TxdObKQ/UiWN3OURTtqo+fXtjY
k/I42pnkX/zP7wGfgC90r5XjLQt4O1M90Fw/oANBo7nFQ6TUYD9j1QOSe2+Iqrbnu+KKcP1l42gd
UoRY3GuJ8JYPf63Qci1xwG2FE3yJeTiEmd3TsIt6/hkmDESeotcKzxIbZVKusQDIdF/dgF40+QJ/
Uuey2DeegPK3u81/+91AQtZUj0lK3dV1MV/wi2vZw2YiuqUhheT4e9556dR2VAC5U5GtqXMQV5ao
3yI6J2DBKfpXsKImGhhzeLwRJSYJ1zRgeilQN8rMnvyAEVRYYxRAHy55eAA8zTSg6XPwV0lIisia
+zNHgSje75vsxE9kKCTO78htyyXtnghSdXvUfNJgirq9/1lqTN/qmIL7tfQPauFJ8i/XdlqtrXD5
v+Y6tGrt+BcZhod359vXO1Fm66tSj5AbXSlA5BjCBgo67603OnyY+guP6u9TzQPae+F3l5juv8HY
7eLQB/Rc2uoEgTrAkyHifccEl81nDLimAa86QwyPREipj3l5DXaLkjBFpVARuLOK0dBsD10p5kfs
cOAzCz9bWPLq/ISjsWMD1RATmlqK46hrygTb9XRe4drMROSup0RS1Ezpe3+stuQbCwd8w0QR9Xyw
ZEsRL1TyZJsDpeK8F+FpuBXfteRrBlbN7Aqvibg+IOa103Ffxvj2fsO7+RJC1RIB2f6rG5m26D1z
Uap7LyHIBHd5jYwblawYG4JFudlURYAtQhrhm/S5j6H2OJQ4IrpswzaaTxh+4mocxJ02Lv6DmDeZ
w88F5tUPbYMugV2kZ+5sEw+BRzPNJqCQToH+nWpl2OrHMc8OMQA8zGR+zx0OFdyrX2d2O0tsdWL6
Ap6a3Y4EmeI/+ZlodQs0lcIEidXUm3QSrJCz425M3V6gN1mryOCQ7WbJaPDMR+2+S6ZzbPNlEX27
RzRnX4KOg7GrqG36QdHBqeZjnwiUuAbHYsxWWU7Y+uV6G7rneXkrx2QWeIuWV8IEQCo03UBCshi8
B7xhmuYwviApllM3vl4pO0cK/TLhfVfsMMdmK56VTKTFOH5dfQ/U66nMzJYB5XzqcIsK58DDxyiK
6WbcN3Wq0z4PNuoQTe8URD8JAQQxN3fnE9wO+9kieVAUTt7Zm/7eaRhFwxsb2nRgsltZfvsbfi7w
XbqHo4xNQs1G1iEjdBKnNIDzedRjv2fq4Y/GJX4GR2tvjrfugKbkXBPKisJsmeurxpGXpKgwd8wO
CS4nJvSSSo6r33iayqmmkHxDy5C0pdBnv8aCUUq00qyZjcuMDgL+AT8S2qQRbrZEOotkxXuCb0LX
6oaVjIyHNn57PGFqxSwKgFb4OWbqzHiCxXTzf59Upolv9pglZxqwtsKoC7uoetrKlui6z4N+ln35
8bQ3XI8Fo7lwWoHvSyMUw1sROLFrh4ZKc4c6SYsZCzpzfMJH6gAcmED+/iK3NmARzQ2BVEFCHXSn
gXS7MrgQPFl0FkoK4bQjzn7aqywWhycQA4MDS2Eqqb5NOqKVX/lrBrgvVkXB4+Q40NWW9uTXSS9F
L+a6undM8Q2r9aq7HY8CxOdoO/2nmttkqmiYqRnD+8fiDTNU82QYy5v3M3dkAEmCftD6Xeod5/tx
7cD6z0Rl8yS7SPDb5NtqnyDGHqCzGxG4NJ8j9Z6rxDL8W42NMBOh7CEfmuy9RnzOYt5RSeNQIMTH
1tqF8riRuQJ6i5xI9Pn5j5nilehoYtDNKsC2ycSAHorFz/UgEk165jlg2awDT25yiZm+aJftgnYC
pbetXWp56PfcGgPmBk6Qf+SvyAzKCWKJ6YX8h2XawAIEMR+W9I+GBE9Z1/kyt3HZrT8mUszSkFpg
l0BosEDIyYiHgDBHOyJGOk33DpRv2RH4ag5rrnOrcvkfsJvowjtcUpubbbiuOgwSCHMTGRU3DJBf
d0d0ASHXTJNWlbSxgFS1V0IOq22xRhmi04QI2CcZWPYcUhol1TgVzZFxXmI6sMefADZMWPdynaup
vnBiUkcwCtAjrHf4ahHEs1wX46e6sBLGRWpFwB24sqfOLQt3UmDgEE7DmWHD4Wg4NwaicFZXJTZz
xsyXs5GMalXKIAKg2PGb2cvA/yAhx85ztGhKV4KuwGMYAPA44PVM35N3OxkY6Wnzmklg6wMDPU2L
TsI+etPDZb+yFKv/vGZfTkI7NkCKQrqVS1Ou4D5Bm3RjPFF3kkpGddj2JT25ks3DPvYbaVDiWXgR
6Xot1lRzZBmwkjuH7N9AZK4zKyG4O7oaJTk1U6Nze66VjgDtdYXLPf/FaiC7iAmRXOVh+BrrzDfU
ufahtpbeUT3mmA6Tb22TbYtQRrpc5Vc9C7VFzidF3PUkdPl4M2RG+kb+v/jFdmZJIu/IqiPT+9vh
lUImI2JxOyUXpY89Bn+21q9t4JlPFt9l2uoHStRj0g0p8In27x4tNkZ3G1vCKFrmbQeHz9AnBunv
X4g2g95bWsbJ/i2v/iX5iE9PPC+DvYCNLm2rMEyAJYvQnCpGZv0c54O7x1TARe/8fcdnMOogdqCR
q2D8qLiTfkGmJ5MgB5iA4D7iRewdubboQoCVV8iZKTaL9EzJFbPEH2csunooM3y1Y/2PImZuXoot
EWVg0xjVDTTa9aE+RYhd/I+ej9zPM/YxVudDOhrtx7SmQSsgAEhbZMPK7Sh2onDSs90lvc/CSuqf
sOnPes/yx+rxx+1rVPw7gk2VWehE51fd8ny1gsn/yHdAu0fIRWHc7dV9nliqNj/hKp7CsLuOAH2/
dmtg3g9lkYFjY5qCm4VkvGV9f8n6MVZqnpIu2CsRecvRfOgO3wQAq3UUVuwPMiASPri8XHJ+Zh1N
4+qubqvAQW2fLWILS3R4JIN3cxt771n8sDrjyF87timhpWt7U82Z8RLf/qjdqXTLd4SN5hDSxRlz
cFJ70ESrlKD8tJ54+Q9UFB82DhNthU4HH8LOzoSasfyxfbWz5NhcpijB6Prm/LKEVvfAdkRw62Ek
fNvi9JC1QFCAO/PeqEwaslsrpYnNJHZ6Sq1XRWxOArWO2A8amYHp3da04csgdtPbp+RVLRR0I5JQ
Qm7y16+u63M/f5ryenBWoNLGbH2P/3a+69V6ydhjX8QEYJdZwRjVimryWGfMMo9v2LlzmHLjw4BW
zQfVcHU4hm4ES2tJXp//rgMCv2kTgxsriABH9Dz20oxWmxS0MaXPoihwcwf3P9COu3SKnyzJVyg9
IF5OvLCgbIs7mYqMfzDGCOwrYnElvWslb+0GbcHBAMQ+Q9GiRszzG2iV68tiyc9DZ/Ve0AkoL553
4G3kjtEPbL9AJImdhcmO1vdwF9H4m9nayWs86ZvXpK+0dGB16zdKTIGo+aRA0VSNsEkb4Ow1/nis
LJgD3pkyz8M+rbAIMomU9z7wbSKBVySSaxj+d/aMRsXDWiGq/9MAKimGqI+rjE5EGR98n5fn4ruE
eS0QXPpXCY1apy1MKFazyU0bRfG0XnggtOdCb3nBXISiOq5OzV3mK8pJXpEfhoFQ/FRJGS3esaTG
ccor41+DJDjukOHVIMTL4AMJcEyGiyhXwx8OOQTfsKDBMMPR2Xa21iMmI26zUwWdZS7D7jsO0/b5
WMbioZH1p2Pg8/f4XDSMEh15A5yQuI688hhR+y3eLy15tR/EjnwQIlgng2ameYH7x6F1kAypKZzh
FLWvr9RXkeuSw/YcC1xiqMYpRi5eiC0FlbGdUkF2PJXQal7ZwwfR8ec3g3y0OzymwTSwhtz4s2L7
DkNUT+RvcxR/qFGHRp7JyLfWRUaj6+LZr4lZzsYqG8Mpk51oXV91R05zcozZ2cWnx0E7Wwdgr/cq
VEN4lGzZp3lG3bC2FldPs0A5YwcvVx0c26nU+qsDuV6OEz+a54Osfl6Z719M/KzbPGQUDFfRxqHh
Dt7rMdzhm4LAKEJnsQk6cdhBJF5cNuoFYbqpGiDckcQxj2IYpMAmfAmcytTHo1d7jddwCiyjFc2R
MTYRFJNn80yShW1JTCx5x+kBJaLXh764OzX8T+g6KK2NoTBBrWI5xeSYBoGqApN7dUO8fNyIF3KM
9SxYOk8Q6EnGK0teLca7Y0nkfVbtL75+DAPKhOOu/RQJIpwItvijvJSuE97uNj83QjgzjP/zM7lw
clEQ2HPAAT57ErLIbMT5l41spvQcJJS8WrT1bvmjC4LUbtxMU+4bEwSxTvlPvyFam2ANhCmNBwHH
hSDHfELc/bVjnGqJSfrE94MdNvg3PKNrQhKWdxcdBgmFwkdu4nOrA9xmbURWS6nJl2ulsZ/EiIiv
MNdMUMhJ5j4SNknAwjUJ8917QxVcnW38+d5If8qYPVDyPccdLjdWh2mBSvJVukfqj7gcUUpJ3NxG
bKpy3GwX3WG72VNGxsCbIGXy8xUF5ZC5gHifLKGYKdvgXVCqKflR2uH2dHIj5UuFqzYnM80MAQWF
dxCHKCQE35AU0+HtvXZg0EW2STpVf05T1OelEgQqD0HlTKBJ0Ii5Vl4XDcExAA7wZGviWDcTMGa/
5IV48UgL38jye1b47K1crw1RUXuqyWiFRvyCLuL2jL0/SlN2BzDdWCljuFa0h4+wzDvTO/6SaFWt
oRudswDo9uDwyUOzM39RYykRJf2TNmu9iNmXByBxAiG2EOmB8B70WMBOKcwJqfU0/WyQj7Os0UzM
MqrbP6lYkSyQyMOQyJSVaQasYIXEh4T1DY4bSG/2wQVCigU6hsQKUdAuvP8EWesRPp1XVWOjRMdr
FviylDn2wqCkGJ4UVl6ykpVuw8rC0pNO+sJ/75QKpw+RPr4bjRuVyAfmrWHxfK/z4ySpg4+9rD4z
bH5K7ShsxuqiPhTALZmpFDFqh7xcMCRBFkyxL2qUYVi8xqnNbUJX2SaWSCOB9UPVC3NL0MxkBDKp
kS7pSJsaKvlkVUhHzCbIPvSf+3w/k1lQmQGR5AbSeWU3fmzOL8A3o1wDrmFvSCtXTbXMNq+VRxXu
qJ7A1siS5F3AZ6sFQrgRsAAHdihjMaIUr2tZAJ6b0smql86zge8AXjcDNd+rKAY9B0UbQ6v9iuIX
oDFc84oKrmYpVAB0f3PtnMSpSdyehQcIKEdZeuVRTYM8hyBJnkb+SoAcJ3kHo1kQx5QsK4sefPtO
E1FlFRIheNiO7RcLlsSFvuUsJIeOu3oAWDmKZNcPjMVCeeEK3B0iYZr2OFA7e9z0xcMb1ZdmCx7N
PtFt2rQgDSKKVDvCa0UDhLcgtS0a2HOlheNJ02j1FrlE21TNMQR1vacQnJOYFCAP107CyYQaMU/h
Mewdye/UtWHRCj7jdsHcWTY0rV2nNVWQFTFMy5Cgw6cxkveqZJ0qhlTmgucPrzIfsqlmLxUD4oyo
uoQEnW3dM2glqh+NriE4uWW1VOTSNM2ujq1UmLHtuU28Torrhcburni1KPC7tmEE3+p5OxoNbXD0
n8Q2r053tTcJCD/7H8t6N8bKaf2jK2rwXLys94FzTWbOKhPIeEd7X8b25yKpDF0RAyHX5QpFNNzX
WKDNHeZ6uevFvZxCQANLvQN9rrFj74vSg8CQSx7S+0BTiqp0EHPMzUWzLpKCE+SxNnxlkszbRZW2
LzoXqFsBz+qpgcrb1ND0NExuZJcx96/GU0/gQThzuy67n4YV3lCavgcMc5ZozoDao9BvSwWSXuSH
+HN0qLaPsOWSIxcLdsoeY4FAsNPXuhy628rHHqiAwUjYL6XmwycJC9MM1O7qTcPTbPH5p7O+N0J6
/PRj5GnvZTstx1dogIUltmWE7LG44TQERn0bYJmD5c6Qj3UNCohE/vapY5uvXJDpxaIXXkllDsFw
8h/Dl6ofBbjZuVOe9Zi0n6vWyjLoyARikRF8CjtL9g1dEPUAZKwycNOM9oDnrYm8g2ijmO9Q5Pce
Rz4yIKXLKXPdR5TaJwdBLWUYDZ04/qOhfClzWLkRjsh6P31l5ffeiB2wrFGYAlJT/c5dZm2wffPb
LJIbYhRkTC0H9Xau6KhFQYeURRvlsswD7X5HTkHwg8P7/Fk3Yun186YwArG18Lg3TQ/03YrHz5Qr
k3M3NDnS8rEJB8OpLIjLxz8akAG5HhzyzwrfBcPAdsTs41KRTuyz3zr5GrTD6bNh1du3aYwBK6qa
JA/Um8tF1OMJK4m9hCNHZ90axnWPv4me75j5UZ1/p8Gh8D8KaOPDW0TopiVn1WHpA+kcImJ+LaeV
zwE2t3xUuJADXoBuI+tWPH4bJYR09Cg0q90S0AkIOPll8aCFmrL19cxlUT9xdVeUEEpoYPjp+EHY
AkVI4dVsdCSzbOYyh9SGv4LhmJMBTGFcDmQK84hMdCOgegE9UKiztjOR/01eLYQANVESLxnoQkJd
LzdEq9SGhUeZY8yQfwXDBhbL5b7MZhar4VVxVbvmiL6bK857L8pc9hkpws2uVPOSBSBUWrnVHS5x
6YzfcKxxXGqDeXkDuui8n/3WZ9/loZIpKXnYWhNSH/ogdHVG9o6/U4gZeP1k55hUu4kuP2DvDiIw
rlFzSXLOQxYCtOVHgovMHigrm98C36navozeuZ4+AnDph1WO5+nCAs4//vOOSXFeOewMNedCuav+
1Fb1/y4673psTvyNfLII+nBk2FPquxvd97tD5Me22C6XOQ2V1r7phUTSyNk4TWnTIsh/J8cvySG9
z5hu9MsCMwFsCPxkrejBy/kRj1158hVzf8SK6ivUSjqu1VtIpUCX6WuqlqDtlZ0ATECk3nSMbcg0
AopLqQfolwthbBs6ySdXTvov9g993T33S+c3HBT7nB3UMg1MkZQR4jeudpttdqlkhLXZccNxUVmh
kwqbS6uN1jT2RML3K+8KJssp7Yxrzc3E30ukdY2ZFCZa9sALA/py1gyrC1dlgP1698FhNpkKXJgT
yYaKg6TR0fOHbYGBRJZQisU2AC0Ym8n8dz4W9GMkgY0JuksOgdkMR9/FI48IKZWEZA/AW9skZCKx
LytrhzPj4Ft7iUkxZjEEB/iWTCIEDB31AkQcRxl+MvYv4Jsto30OiNE+0X7unasaZXOBNzaarb0u
fEPsP9Oz2e/0aApW0O3gH0R/R+oQaU2S77E2AfZI+2djKjK55rGAiLX+Takz+ANGs9sYMNPIgDOe
AUCpPhzA4kwb2myfR1tPzD4wbukgBaQavG92HlS5gP43aWMwcQ9fekydMx4vV3gkcB9HAzs+JSlZ
+1OJzBA0L5VQfx8msET/2ULWc6Q5K7ztuvuzziVqtc/ZBl4KOQ6R6VTSRV6FSYbBBzglZQyyAZyt
9t8MWe1iurXkxJrGorvw0JFEDAGihCWLzpj/yPMu/dua8FctaHS+LNuAmdpblUy872qaLbTo8wDx
JliDNIsQJzv2sdAQm9KFXHGMiDHdThiQemBUOHzoNNdt7TrVZCVsGZdiY8M8VFafxKYKIhsrtdX9
yLK6FUJcC6m5ZHgdMWmf8qbTM4XDT0GzRfdtXvCFkFcQFaYEXfnpCO3TLlJmzcasxYcXxB1gQ/3R
8HikBbBWAphu4Ab3Rrqo5alXMJkks6q2r131dP5QgRfbrdBNyHesFD1udjQ3vo/2umRZbdF9LjyB
3qzc/lRFq9cbWvlonH34G8I+slZv9CnSXKq4e1dW0pa44FfYyioGux9wFxYURmLDKoCZzScUwe/F
/I7aTICkku2YRFCWTcDDGoDrf6BkBOQu1rnDJTNMmAU8NxCz8vssb8zoskwAyWjHy691xsebXzsJ
/JXgsDR8DfBoDMn8HgekUaMNQjwoPseI+ycRdX2m56qh9ziqIaBDsVeNBpzmNg/vphtOD0eABaMU
RjpurlibjmtJxEI3Sb2Eq0zUEebco/CJ6ODmjum7c/M08RxjGiHougTf/1v/DEWzL0jVd0iqZxDq
TT6NxZ9aUaK2+1EzHNOrZToLbhw1mRtXpoRqUBDwPWtNCkhRsyfj6wiZ/OgLLEK+srds0J1h2AX+
Km/nd45XEAeQgbqC+qzVioYIy0d1BGy8GHSAVuUG7krdgjLfLtTOx+gIzhGhmQsLLhlt68qP81ri
AbjUBhU4YFO6dWcb/5muI/tf161QpHWURJJdUXcH33w9fS10ZvUuUsY5OPc1OAXQ2QhFl9zzza5t
4dAHv+IOEUvxQIn0351OzbJNJRX7HuVzLOGDL6vKRmfdD/HMd9/+59cbi4yAKpAYD3Zsd7fSXjkt
OqXI/jSatM/ys3wr77x1RDb/f+kk1O/eUDhF0EbvDQ9lkvz9OmWDg1SqdhN753/MnnnLJHllIUOU
1Nf8vHDPNwzAKT/wExLZSY3OCtKMRZf3Op3JCpIlMJL02kC8iuae+Z8okOpYaiSwMow2ATm0WRsb
Hp/lGWjPYRBEkIDJyPGSzGkCtuxvyjFeogrmiMDbPj0ZSyvv7lC4q3WfJAp3kSVXMEdo/2m/j/Ao
u7Wg5EUXA1nroX7GKkgIyZrzDoGEV/bEtojGTtDDGlJ9fqABQM4WyFQ6NiNL63f/eQp7dsluuV7L
avSgg5hZxUM9lfNdiEiwkQaEqyUJa9iXNHoxkXiwj7LYZsXqu9UJJw41UzJQew8oYkCwrOC1jPg+
XjLo/+rS70LSYtv2BYFSYYgDWADYFRb/egBk6kKYNn6jvvLK62JTkjwMGp85L4dJOcQMSih0UdYC
RZyFH4wbV3rQxRl23/KslVR+GQfVTTktPugQLGCoiUgkdUx7mUM5xbx10Mgx5HVd9zdc4emxcVpT
+pqA0Dnfl5dRDFAHMAxQTJX0Rpj+V4BasRtsI4yVWdHBXa9dmz5IieCvo4k+Qha0LKWcoo4C1Ez9
UyLtd/HjFB/7JK9qrmKzb6N0GPWd7xxgMI4uchCDE+XxMwtN5OqFyqrp0O2gW/uTm9hw1rEuLV9b
3FIjG9SviVko/Fs2Fh1RE98Ds8ssGs4p05SqS8obk3WuFPN66JUrZSkQHsQoTXWv90DNUhQ4lajD
3YAjArOh8QQAaY4J4XKpfRH4dg+9ZbAgSs2NBJ9NaI9kI8MgK/xTsqGD5UGuV3lp/fqvzBftoPES
YigSHHRTY1FFE+afvlzEgKuoJm049iZwkzd59BpBLimqxoJJCWOlQmLCbV22c8fxeCsOS9xzIQnI
8X9FG//0uEJZYhaJg26cwl2MbOz3AXRqo7w2eRUpYvReWgm8IWPKfajln2hlhLxrT8HNuVsUpB4N
ysmzRw/i4ep0VClvAYNvmgOYsiLNhaNptWLg57CpnKrdZwW4Pmu8LgnF+8Cc1aNFqCmFDgMVLcO9
3EdC21tsQaBVep4YRJKQ1U0+A6YHTr3TqA1yb7EyId1SswbpoAEyJQMdFkPIdOW9ZflNlEmyaGzf
zA23Yi4ka+Dejc5ZqMpcYU6z36IyLn3RcdctMshc7QmCTtdSjJEdi8LE+zpCtdK+d87liLIaqjFN
WCfbIfyB37YMcJtkr5QS34dtE9KaR4pR0aJUdxgz5AjT19IvY7puID28klABVjE5cC1yuuL4Gkvs
30J6qlI8sCwK9cmXhEprBscK+dvG7Qj3zvlG+RJMdp1HKgFRYUvkRKRmuwHdtCJBN/YZiKgNO1mT
Hegtyqzx1BZ8MWJTFiD1+RMUEIGqTSvrejivjenTFyVM0GTRDlf8m96ks2YJ/UWEnwMt8Et/jXwv
4MjKRhz7p4AEb5kNQ3oqJttD5OWrdzuHdam1wY2JO4ujsw1JG7vs/XPIyNJWmi8yIUaPdZM4Yuv0
PLUK6snficMLFOYBTc5754KyDk28v8fTw48EuWCJTrW5Oo4+hhPmD83NwXXdITaQtHkcepuM63jI
mAw4u3Ppma++G3sK1r1+kVRaWKtDZCec+6I48uSg+4RMJb6VXrFSSfdY0B2U7pbcNqnZytU5s9Of
K+Qi3gZ5vn7dsI/VyVyyXLP8jkOM5ycnF3LrbFhgXrjYatFw8V/v16KDIx0QfeqLXw12nADpYevB
M3KuwekIM6e//Edbrzdq5LHtbeGGzxoWvMzL14AIXWhdiA3iuPkru7FUAsVCFII0/Y0SMgSBb70X
FmFanfrb1M6/uiM69+sBK/M4VEIvEn7d8IzAYEhpm1BENdsnSVHjpFsmDlnOdDjx0ywCQv+n1cVH
tcpwVsHPn0UoOjwo8vMUN5auqrJEWioDD04P1SvsQbTvSRagIpNNIKbDFke4StDB2Ei97fY3Mne6
oWwtNCIWkHI7yY3crYYrtrcg99abZNs0wgQQZefTxWWIEvksIe8MD+sx46i052r2x30GcUzDdxbY
X+4pbDELVn/FBbPST3/V3vgNfSLQKaZmJHr5v8N1yTrbW9OOVgg0q3dsYPs8Ggw3Cg+bf4fPMJPI
23uqEYZRtN7nWkTlasoynT1PNV2SShjI3pyTobamlRwCp54q3JJakZQOtV+Ke5doukqBZK7Q4CJ7
zDzaMTwtacR83A0fAb4eLVlalNdwwOhdIYwV5DmyyvwQHVkk8pJsItK2Z60iU4MYkIZ5fcTr4n+Q
v4LYU0XnkdjPOO+D9LvWlZ9KoCrkRbucoijQqhSYPrF7wywaLJas0Zx8Wfxl+ft63ccS8TRZn2Wb
C7bR/xnLOcg1aW+xy/6O5k7Mgkz3RAVTgn6wwhWYtkLP+jmoJLtrZNkZZ2MTy1DAEQ/1Oee6HZ0T
qwaskiM6pjfbl5OQZTE0Idwq3Dac74hZmU5jhLuJtzPOys4Bg23T5mQeykOY3WLT5o9bHj0vhNTJ
WEDYy0PGIvdingxtaRYYaNoVxv64TPHd4r4Kl05r3kMMCUt6+nsIwzID2sG50yLEb2D6h4ZG2nXO
u/YPRu5vO2HnMw2A8BDyOuKDFflG5C60lqTOA3bvXoFf027gLN0GhVeV4kksKMnmcdOGjeVqQUEV
4Fh3DULrjvgAKX4ZWcfVjJQLDo7sJNLKseFxcuWe+nNpwPuEOfskXXDj1PUZ5LU/U5PAR1S6CQWj
5/3nsvFnu3IslrGqskIjrMs5N7X8o65uhMuOIqntpokcHRQGXtZbKqE0Ef1S/Yv4G9IxZScQOQvI
PmMLLRPO/6u4Y1YLLL8lx07QlRIfjIrnZkw/Z2JfkbaEXh4ppOWfAPe0MQBN/qlutp6WN+1CYVMx
lXl/EgAXUQ0fM6BVnOFKmDyaJ46f8DMK5I2SbYgqRwujjYDilXcSjpiloyiLiNrdCkuOtH0Buxjd
KqS8aeY6egLcEi8LQsfHyb0Ln6lzkbzUSkReeFxPqjHQ/YrG2UcDGGEFcRxtjt0D/b0Kv4EYGzXC
zmgDTimSdUA99Vvk6W2xrO964pzrNIrthkyubcWn9l9Wq2pYiDHq/Cqy0LSg65ES+qahgXa8UH+a
M7yFC34rmlBZumCUQ3EaF6dut4ZCbT/9/fICSlu3uEm01jcoQtCJ2jXlUTWQTckDg+FRcVoy78PV
aB3GUKUgS7E5XTKtVFiwG12KIxyf2P2hqcUm2ASCwtxUThFkdfB/zrQrDB/o69mOdTL/IUsQ3tkD
2YQYQrSS5c0Y5LbywJ3oORkLC+fhTh3y9ehnd/AxLgDD5z2gegAgMviRuTdXbW0RH694sDThoHeQ
Rvl8kGg0U83Oo8S+APSoVjVbUtX48qyOcjiBra7ACpmf2R6Norw3DLbzv8JBQIJBzogaMV5SRR1g
79C2IeuyKDTAJMbY4ok5rr4jhCpJ/RrruwAMa3PTR8fT/sb4W6eXwxLzoPOmD2y2Yo5FCuJ51f70
KCenoQaymgb0ykovun3pSH7AKzyZjx20+WxgFSuoYyU5kyYk0S1J7nV8LJQiEascfN/BEZirw+0z
JcAxbeRF3VdWRi+Do+KyjhzBPk/vygEIxCEiP2NmYNam2ThMPHMs55oMBv8oezHXRUHdXBgQDqXc
IhkSdqgSr/x+xEdWLVKVcp+hJn18xXAiukqGCV6ob0PKUPsfojnG7nJYjxUbbnPnUXEojTwo/RAc
ZjxOA5528VXUyXbAUviWgYTirHNhQIIGc84v6Sdg/J5LUXF75M4WIVSRL/vnghJFN870PmpoxziY
TFlq1tWFGhqR7Cnlaolqr07xXhjMTbV58l6Z0yaP4YO3VTKS5N6RtjZEN/tOhi8MCfUafpu5h893
UuoVfgx32nCitBTlzCeZG7OqHNynUWJb+B4A/APEePELCpjMNTg1sKvqV2azzzxsU6st+f76gdko
+dqR5FD6AVbdZsdBqd4SUMzPYMj16mx+aZe8HAs2oceHQ7igpUm22zFDCIA0y6AyLHcxsT9By5vb
qSYFhbi2HjU519UANPq9LqtU6zo+G5SeXummdyjjBHTAULgbOO1vly1BUVUAGFg3pFYQXXURLuk5
caHrHJ2KWFth7IyC6TmtKmumHawQ+uKebmJCzCL7FezbKgz9o+htwWhxpcTs7VQ4SGmMr2Of7m6/
wZZLhEZPCsUhMr+PFKx90kRTXwXsOwL3MOtYVh2dxC4eiG0qUlokvcQjVbPfTyjL1s3ekKluMkw+
QZtBaHKPmEsPChIucDLnyYn1wKvzj+r5Kcb8mZNU2xKe/xgrV6bM4RfCJItrZYz8E87vLCUjv5Em
onCn7LYm/JbM5dvHcDaW6XWeknYELM3W6YLS1SO2Kxyid2ZNqveyKkyb7hRdPKhxZyKyXOdwgOR0
nwsSPjQqi4ydyRCu5nPiQZEbdVoMNmXFyHriUStTbfTQv36V0st6WUr63eZvP89AEfoLwPTDJrhg
tuYq2DWc5g/Uh2zMm5XYo1wEcb4LzZ5NZwpjDhw5hZoxl6pnT+yCzv9aA/hUOsG16imanJen6wBr
1E8ThnUWnU0wo6LVMuKZ2yDqSOzTZ2w8L7T+tZQZePacbkMgx45SjQx74oywc4lKxRaZ1GeFaVNW
UwbwU32OlPqqXmtVst+wWX3dTcO/cQjYUShN59lp1G59WjQhpYwsyWZzR/0ijQKiyYfsJ6qwVA/2
sO5h4GkE0QQssI2q2UOrTRiIlcYlbob3fM44v/iF3h3Ot2HYWcsykMltMMVagV2tYo/uDdE8ATND
0EUrQl7Ytis2Z5oRQmyGgyiYN+dE+OLgZyLQGXRoGWtWRCwLyej5w08W5MAihT6XY+qQMLdOscly
DHQGzNKwm7s9o/LN3kmhPpP4VG3ubBe+boWmrv9n8o2zkizuGVULjHjgafCbdGIteP/ko0b3nQtT
IqFh5puM5fHtYylFcVFlyy0LSFb5hb24RUfdrJ53ftOTmplGHudpxL9AIgjrubRMyr4AFD/Frkdc
6wSPSEqOqlGTJMvZMt6ZacRt9MdiSRpkj7jj/MxuMSswbX/I6CWsaTYqOR2tOpypzNAuimyqP7hL
2nweEH2POIgK7TU/BaXVIbR4gptQoopJ0PIgMHw1n/4xrd+ngu6y2dM9fgPbc9GWqI6s/1hz4AVQ
NrIsRgOTEW6oMGoS33z3ggeo+6QVs+HuepkZKE0uqEBh/VIxJueD5JxM1b0LdiYzfAUHCjSrbGj3
EEUVWFPB1FxJeYAvnkPG3gBZqDkikk2XpaU1U0xncTR7k3jkhlkOEMb6KFFz5fp4h0kgtgS3ctAA
B43QjowoYk98UBfzaUxnmrNozX6LQ3TNhLIjiE1w2elWlWoxrc1NMOU9j44+acmDIEfk2boLauA2
9U7TEDhn/pimLOgf7YDMARCrXELMXbmadgK2tIjogiVkBdO/3iqRw2hcbjNKdkJVGiWYAoDByqFT
5CYjlQzHu+CKZRMa7HZk+tOdQ+QQK+dRts+GN2v1t2RywD9Lpf+j4QfUu+CQiEE/Ughd3/CtFryc
Zmn4Xy7N1lMRWDVYV1eXT5GRzDHC75S0oKvDQP+k1QF2Hy52lnTycPjuAVY6GNs6Mxkaai/YoNYJ
n5Zljm75WwD35FGiWGwElY3ZmBzurSa2Jl4k8YKPkGzOwLWbr75r7f5336Y36gynzwfPcboI9nmb
dn8WPUa76aHP3bBNeqKsGgFKP2fRthel8R1bgsbkloXBkDjYDtjNBhCRNalQKmUsFyoxs8K0Yprw
w1r38dymr/35dyShvOhSFfKcBjsR4ziEk+/qT6xexkz54tqYLYuJIBXUSt+sZwYOc8CWttKH4C6j
qnIdnpfYo5n68OcdbeZFEmeFKfHXAlkVULRl6O/CVkWtUXlnVgFITMxTNRheuaHTsJ9elFzGx+WZ
edIhO7qT80itY9MNph45lqoS1QlUg8RX3Xb7xVEOcZ7HYMpOUk5uv+Mi4GIDidMMqlhtPEe1e8oT
l1W4sfOFycnraRIfDyvMXRDOE46O/mE4PPvmPhzJVsUIIFSAPFKLSGb4R5nlM7Xwz3w0oUOfWzUp
76RyJA/hmlmha/NkYB/fNeGlSA3gKvasNFqibLmxdttQwaiZppVYveTT4Xaa4ksWXXlQstFQjI4M
kLvTue7gd/iSbkxVqFPdmhT0b4lUCBb/N1O/CKgCp3wkhqTSlDJXh6mGXivhhuRJqfASuPhV5fDv
PlShqyAeAKuYhnoyne9lPJm8QzeRISaMRH+xudsfO2Pg7o/hiTx2pS2gHo19dPELwGwKJhMaMLFM
LIW//NO+E/p6+0xIggAvSuYg89hEhNt1xEoH8VQfKqVz+jyvY/VvdbfFf+52MPSzRw94BWS2Shwa
ZfkB1SelrjwTEyTb1nuwGnf2H9qmymdOpaYGQLlCuZ8Agt3aj3mT5+US1rhi3BHHyZedJK5FZ5IH
Oc72p7Npy4DZb2w3koym0EQa9SE8UxeBkbdExUijYLd+sWCpQpXrbhOWoMBsJDONXnL5BVR7nfAU
LElPB5nrPo2arzDtPVZGDOborPBj2AJiAW94T7vbMpl9ubsiGgF8BuvF7PJ/jbXHKO9ITw+SgVzw
NB0x27IWoBdQ3vcw4LhT6Q+ImydoDSc58lSJ/z/1hk6ILhVchPeKov9fmO83UshByVOdgvKie2dM
NntNJZVs8K10eVw38f88q8mvFlz5cYDL7Z4T6M7qdcExyC3v/OWzVT0y1BPcS2A+hmNhvXCbC2mR
OpiY6QkrtLZ8xHFH4RQRRq+34jd10/6iVTJuch6Gm9zjA+Lwh9pXrXKFuPUx9kBzQKGdeqf4tc8J
MkKfC+eIFRg83BUTJiSvhHo5vq81/O/n+CYeRH68qpE5Usokz3Uq00Kl4v3PcK+rdvDRL0FeRkXA
vEGoh1hGfC2Mglpxt6GJy+YkAg9mUOXm5Lt8YtCbB4HMeAzqZv4DwfRkBg7lEhOTfP3q7omfQ2Bv
0uu0nDcvk0QRE4e2rEOy5lC8fIyU5CGCTmv6noBFQde1wV2kIyYhJ+KxFNdpHU0XBSi1InRCYSVv
Aekr+HJhbfS43tSyfNurdNJzWyZDUamR7lhxNMBX55nSUew9Fmq0Jvy4gSLGXU4ov6rBpeTGgojy
+LLp3g4FIOPtOK3/C6s2kC+sUeDerXko4U8OYx60hsx5kfv8FFKhCwTQ53Y3C8PWZNDO1EINHk2p
jnWgG4tjheeqmBkR/v2juc9CQSvfnNifHFb5Qg+xw6s0ws8jDWuuuipF6qApIPGN2YnM0BYDB7Ei
j6fBvP2oc/CdmsMZD8lg+RYj+fIgpDP2YRy06BqKfIRuYJ/g5+64Ga9hDLI2xo3Nhw5IZNlUK8Bi
VcfrvHAOQWwuo395GxKPEcMS1781qyI1cdZh3XL1apG6unywC5NC3E7FvbE2QI7cbb6af1hfb9dz
Om+BFvdvmBTcMb/kX/A176hHfClhQh3EvjTxkyYi1g96vlZBsRoRWPFBCEK4y8mT9VmFXuWBL7Jm
KetlhZgUXfRDv46s9pCsCFZy6w/Hn/Shj2jm5DAe1XUAz9k6uZje2GPmH6EXsK5k0SKSAS3GtO3e
G/Gu4ndlFFdN49L2ljenY3zyq0pbaNqnx4zKKdYoj9x5yVZjFdl64z40r48dMql0rWBXktegd1iH
a0X4JktKzZaaYwfPigr4O1cqH/fzsganLnASJpYTWLG5xz8hzY9bgxKFe5ehkgNpgrDHA35LKPt4
RhmkhHdGiZdqLgccn5rx4wWrImRmZHxZLo5hcaMKljAUHOG29KS9p0Hjt0A9dZtJbTAtR2eYYUVm
LhHaT24Thym3Slb/1D0bLvTtI5t1pYA2mISQormaOznd1SCeb7Cnki/K3hFKWDz8tuHOd2VKSmJG
+AwMf171nUfalY+AW5sWX3HqzNEq0SBNwgiUDUh7OhF2gs0y57sSJFZm4wl2k6NgTPfo/GjFcDA+
ZABDv7Q+c8KgpOYfU++DF9ebMTbriCdywguGgtu86CINYDh+xo6feRZDAFzBbuhNnsBGOmRXRygn
6Aas1OisV40YC60+qkxSUsy2wJ19z3UOdtPqTAwYYWj71YwCcupWqmI0RufHPS/kCCFmiaA4AIj1
AemfRrtYlK/l9C7zepGEsRCGsAzQin/NBiyfICSPIcpvxadXmwi0QRX6OIWvty/NsZP5hLEti2Q1
/p3z4htxHXcrg4vQqWjPdNahRRY1+g7WjkGePJbooTFcIaZmdYpUsIoqLgrfRYg11y2vTxwJrlAS
Oo5USUrXWmI4pZpfko+Oygu6ONhB6Ka1fpIejkwC0+t+IRKkqy6nl+UGz5YIUhsb4LOdqw5lVlmX
LVYZxP02gACFOoDmL9BGiqA6vYrvXW9p10O8lZPk3yF6JPEyB7syHSYKQlhrCBoxwDX1yzBguHeB
Nyz1Uz8a3pz33y8bfHQW+cHhFrEBpLKQB0ERac44L55O67eVG+CZAfJtQVN3Szs7hvVNxXo0+Jim
vgIQ9GvS3HhDMRzU2RwgTsEXgyldfTu9oN1WqO6omgNVZX501abAKYRst1UeUeFg37jKsLvSpbqe
TKVMxEWJXwlpn06+Jn3UcXo9E61wv8sIKMYLnWAkdnyMuaMDB/xPdwNfsfMYZb1iCdgUu3KUIr7y
JDBpwCK3NIZx+Lfu0k4wYF7qTE29GBuD6L9zNENiobAtfbNe8/TJKWNNanPOEjTcIcF1fkN5rUjO
QafcN5X/u3aMvljvlqp+fMu1WZ0frAa0jm0J+4KkDZ6kFWTfNGFpEu/nJsNal1WrbGAT1SWHpaun
8EbbWK+OaxTd1Mn9f7/axj2ELS/MM7ZxW0IiFFMolQMU8tg+jzZsAPvhwG7HuTIOxpguLkdxylX+
aaxafXgkPh12ERRWnmo30+VC8V+wEQwxrXAc1aK/kIM27KzMuygOdD7skhyuplpK2HKWsnO1awZ5
HENJTOkXkFQUxNELSDV9Zr7mrd+FY6REWDWB5uagaEB2/GF6kcaLzZ3dwteLPxtERtMAkRCsRjIL
Klk1ulSc348BBXNOy0GhubXPQRjMuMom6G8SiV1GltKCKjGBvg4oB7VZ0Us3DOKRU08udxsYZnd9
PDP3nN9neZ8bzwYrb/oyyYRKxpwMrXRfh/JwL56kex+YQIg1koQBoB7Oo+XwAcgImZLPZAAhS0TG
sFGoonIFoDvEzejep+d7TxnmG33JCv/bg7ZtANyviKSkrrBALyva/zSJVtsalRLQ8RaTlqro/bMq
wTAoY+gJnaHtbOMLxqfjoEpY/RGzi7zGKZrQ2kZkyO/cZjKc/s79TPY59Z56yWcovL2qTZwXGFuG
OXnEGmJqXFJjMQtKfyKvxQYR3w+NYy49cOeIiElB3A8JeIVuxZX5Ia5YQ7Tj+HAuTmdFBeIEEw+S
583oP618Wkw9m3wGd69+GHhexW2vqA6L4m3aGGb4I4uUxkd1F23gm2IChN/ztZ1f1c0N5WUIuMB3
NCpMHWZMjGZzmop91kGB2HSA/xcrBkb0tf3UwrJGrIkfF3MJA4qxXFqre7GXnOam4W5lnGLx5zCC
sd8JXJqaBCEtoY2sg5s2bA3jc3EOpqWXoa5UQkSangUP8Zyu2nPbIVQpyekgFDIQ3xY3ZQEbYOHk
IjDhKMJslGLIWePFkJXWalo8TDrI1AIaDLqldQXsO4nt422ChJrDHBa3yr6nu72QUEwusBlKvY1C
C1yY+IiWIsC0ZWt9LKc0aVWCuygQShlQ66CGqJliiXHKibWSAkYzMzor6UqhgoK1VjvD+S6oATlw
mDjmxp6IME/x1BcSO2rWL6ElVFTOgs8qh3pr4YTcBIJeGh6YlPC4TdGb7VmJNxXMnf7JAObiO3CY
5jyxkGvxJXUHZtAENtAcSrThlKJCDSbyiiHG02w+vKfwbceCw1j5c18vz2K6gQ/sol1T75qEhpo0
JwOhelrNQK07TYQPwqH9pEYrhA8ULEzlUV9EmIDXltcO8ModEL+HCR7MGikPv+RL2vOKho+Cb/V8
PQPwMD4WayneWCMH6lxKnpQIu16Co5Waq/ubw6n9Saer8Rja/lwprgGgWDRXcfKXREdtaQrh21N9
63U/8Rxo/1GBzQhktEHR8E/9eh1zpxD3Jtq1m7pjoP4Ik5rWF9wxZXjL+m9JIGJ5YVtmKTyaRgGz
K9on5OGeaxUaYOG9DlJiqsYn/Q/ZhGGwxwQyBNnwIfo2hh7c3RNEok28pIbk+1r6ibjNOSUoog2Z
kJSnobLiDUyleOuV8U1xpUNLZmng2m4aHHXxYOOeAi/LTa3UmLOeXMh8Ois0+BbzYLqPl1hbEa54
fcutHnpJakNrA2u4x3NgLGEQ3WCjOG2fFsRwsB70ca7fBjj+s46fU30ez4FGC+aNDe0QbdjznIgy
mmUrWBvdiyZvb4UEqmagrVdjGhmG5OAGeqfGSf13i/rmt2enVjzX95PLMs5xFfmoaiSnP3jeRQzF
P37QO3cUUqS8vjn3IjCp5AwhIrGzHXELAi51TRNuHDU4wSorsGJMyMllMS4coK/UXpZwc1nUWwV2
CUxTKIsTqoPtfxxp7xzP240t5KnBPHayLb0hepp6VCc8pALAsHmW8uGGk0s5EMRy0LdTA+NNrHRP
PDJpNsz0gbg06gDqmu7EYS0zUFS7P1s2QOhQF02wF+ylcIBeFnUPQyx1Q0xIEwWnKERJdyogimj2
y09bbQnUXPG7oX06y5h/SyFwVm68wa0IJ87XSV9EMDtbJPPz8ss7+udHeqwFqYr4+jeph5FyiBmC
zg+GpfBswedo378BIM8wFJI7IAM8v+sPQkayuzQAXTHX1iltDBysJ7WrdCDG+MK1EDd9MhMVZ+hE
kDGZLsQA9ilYpk+rGeUqPNClqcGv3ia5GML0JL4Oqw9cczz6EtERSBcNBdz2+c7g9CKa08IjbwFJ
IF5hbp1jAKXv2rilyrpsFN/uLUapjTQp6aNkUoUIRnlg+WNVt96+PZlXxciMM8EXitJC4u3XgypK
knn5BrhjahNQ2TJrw1FXVcg+2jawvL40oi3CbFj7/k0kgO3GElU9rn3Zgd3A16Q0yzjCqgackG31
in9qXPYYmoTcY/5rKV6sq0VJm0vpz13htln8pPOmppzRsCZXeW0eIg326qj6dWx5mP18yWL2QasM
sTsv8UnGVIYQPaDHvHisQXex1D+MKXZlaZihlazZP5O0U0L2XLAcgr1mRu2zI2xhCYewVO6Jnssi
aFiSxUwh0AmXUd48Cw+wbWCVUlj1rIgxGNyHF/1RPUiuAFEV9vEMrnBrD3IRQkWRakXxY21Gruv+
fJJBefhYOhhkTmkll4aGOwcO1JzhkqaWUisc2HYTD8k8KxuafQZiCzU3wZyEgbzur22SrZJGodYB
pE3vqR7oAFNroGpQJSl8l9+I0cd88UJQX2B6Q8tvrWfmbpYy0J0gcE3qfWYqR+w4NVIVTgHVDh8W
xHppW40ggDdTP9HSq60VUFT11WZNTE+G45chrbqf/rBmyK5ex7lQXeauXOjqVEs6DIqzpzEM9Skh
Yyt4jG3SreCDGaQdsKxkNWyGgeBpmidCQ0dIA9jhj5zhWTYs2xt2RsX4LK7mvWeo3aFWPEujTK0w
0TBeqUCiTkgFFNtYGFq/Kym0+VHPVhpD4NuAym80ppegMUpmp99MdU+zBW9MPv+T+pd05Sxz8ChD
YW98TVXOEDMlDqm4zbdjz5mDyx1qBy0bjipDKMgFsi9P4byN3nWQBYh49G3m+aX71NVj4NrklZYX
CEBuFlVxZHrbO0xNLnXB+BXZeq+5OIyNBWZXwzkcVlILGm6x+CDtmbya2FYQaTASJdQLTj9m66n7
t9aOX78NsxYGHc/+TKRLOe5YmYA8XBBkxjSDb/NY5k3kCwRBGX+of5Et/q49kZ7mI5XguRZDFCtF
zPRQODlXKm4W0g1lXWiSh9puUiD1bUYag+D0ZQ3kxn0c5p/moIUyfwPUr4Q/Ui75LRZ6YzIkTMIy
7BqKbLV63f3hGK+k/GGOB22lrwIL65+G6KUQCGbW/ZVCaQSj01voSrqIa4g2c5malIUscK5jo5el
7mpSSPrZWohctC+1zizpga1f1OX3AYqccolu5lx5jn2rBPpB2Qoxvlq81Th2ACisNRuXJVS+rG8o
JlruImse520I/Yy7c/1snL3r1pIAexJjcEbNeLv5gwMoazcsM3J0qs1+vdRn23hxGIheIAAT6zx9
/Sfh4WslnwRBJXXbKztgj83XTemQWhPkv20btOq8T2kCddIwx856T84YSEw+F7/SDjZ3BSroYBT+
JZh7nD+5v85mFllR6QmVaIu7LaCs5mTgf6VjfYX/7uAjJ8ooHFuIGA8k5dxc1VR/chVKTo6cyoMn
6Jz/fkEY4T+NIpsdhD7/xioGg6bZc9ioDQHFC4WsMlO1q/OCpUnoFqMlt4ZJ/udJ/JzmGk8B9quk
mrF4sMUdnopDVhoiUbU/Rx1C44WmDohMRm9jej+gjlqatUzR0mgcpD4wOVSXDllOXh1AUca/ZKUu
zn9kY9PAdHpopMlkq5BYa9IyytDFeD+6vdfka82V0Yekeha2B6RdMYvGJt+ACJ+VviEIhP7EneIT
g9emvPLFqmY0TI8MWb5XL/1xjDO7/7iEl0Zv+LnA+hoCiYyhgjvAKSM3QSVKejLlcE7O1iWoI+7d
1KLxERUU3PCgwYR9lnFrOPbn7IyH2kS5Y2AwfKniJqLGKT9M0w96CKOZ5zV8vJavxnfNSrsrNiWg
z1tKw88aRRcKPO8t8vPNCBhLpc+BdlqtpbwR1gAEcUV/YPXD7mEZXs+0W41WxFdHvlXg0rssK5Hf
DbBBbMd75yGxCg9ushOGea9p2PnDawRsMnEhvq9nUs30QWbhzoOVsE1NJRmP2qN+1IrT0y9iDi5U
By0LXL5nrryZcBL7776jCWxLcIU6a4dBw5/+Vz9gxSKSVUULjgfNBRombyVF3hf5uBsyGwB2+w83
WjN5KLkX8ZqUGgoh9q+AC2qWP42wlPuxw/F327Zx1N0qex1HfeA07QAX6VFizpZhZlpSuGjsXF7M
TU+eoJ1YLoffqaOkHdJf+t39G1Sq5gOqI2pEC6/2sKVPLKhWbJ+w9QfeU7AWe8Y4rqcogcBcwkVC
sQymVi8gN5sXgJpI80+3EfMAQKODKhub9qJ7da/yZtdf/8whd0keoVwKQ8PM/vQ5PhahfgDeG8hT
cm5PWSaY23z/p/5lUjA2Awt7R/VqKm4jawfIeH65CYeEgtZtfMBoIKqlsdWyzYUrNIHY31BfqDdx
5zcR1qWzViA9gOznA0J0US++yTBkeEDUo9xES9Sbc+KribEcoMbZR9fYau/y/vZ4J/n4T5TWta5Z
cMmBUEeRQ9GsVOnjv7PqJcJNWAxWrNFKp/gGgO85CP2nG/SZW9oDV+PzCHWwivJIOqungeILvTKb
wzEzDFXY6WUPFBPYEItAQt7Fxf2DNSLP47Tr/T8y8RdgnwEbbB4uFnRTruj6asf5g9Ip45aW4SjQ
oSArP/eaaTZQ4TN5wPq2eNgOEUEIn5tK0dl5wSTvipH74x2ISZd08xp4acxozmZXt7ZXVNN1oyG1
TYEXVNq64QRGR6Bt5hsHZ77P0k8PGvP4626CUgPwtsp8t68JTaLktUZ/LF+YatZVfOKLFaEkklxb
N5MgnK5p+EpkpFIlQLBW4WaOymU24aBvsXGEzhHIDxsHIfVVbcrnnLWHGigkfPs8uS83j/SOrbLU
OqjPg4OVns3KUaZZzvbM1GQ6BXWnIrz4RFCxfuVcf043BKWvJWuzSVRj2tfccOMrKwiMgqPJlCL5
ULQcneZKvEQIfmzAHxQQ1SD+omVT9TZgqlMaTb1f/yc2muRi4cMIQslJ+g9jv0nXhvCucmPTPB4T
bcZS0uCyXdWd8ozkXkOxw9ZLUEYo1A5Q+TV2FOWV8FvgjDvNk95D2yD+Ca63ZedPedrDYMifQ9e4
bN4+W1tDKHKEorPYVu+4JPMsFbUK6WNE29NtIVsWgoiVd+RU580ZLtvE4L2crxrRBFMKESZQFc+m
NlmQe2Ncx9aPL2Z8CWyUy2Ot49hUg+Lcv6VqDpqwcFVkZW+RFP9/dSSzm1Ds50Q3zxY6IrKl5v2Q
f5Nd9HJGhwRV95mmxgkhLtLbd+uy/9oarOXPek+2czeJVouVn9gq4Tp32Oip8SMoKwMbXX+pZQn7
MWZqj1FlMKEyeWkpqZK/zGFSdCnLWTBdmFH6oPECJy5jSkIk5GLuUMS6gfLCAssU461v1DkdzuBq
G6u7YQCeiS5DRlK27zuwURXd4li1595+EkK63u1MSruQjFrqq7z0K9wlJPUtL4AxFBdbvOG4jBr5
c1MMU8+Sk8CnSrxhcRVidRNt9zrB3bOYvWL9EIUC7Y8F3icJ3EIipIwiCtpFEdfxXJ5FjBgkRAC4
P9D7OSt5swI6W66oRI0fAixGM1Xpix3/ANhRCJ7MHBP1cN0mT7fLwVXyGnpNPt2Rk7xMDHoV82TL
L6DpY8Q3x8yg5w0inUrWHPJnnUTM0axHjyZzbGUGn0g64fAm1JzbsZv+E8RjI5gMGa5wfI1jU9i8
VN5AckI3/t4R5ynVORXS9UtMW4J7k38TmZxjM58MWADCEhB8KTNDeUdgRFVDhv1CPWcjCNds0Kmr
B/GUMzPek/55Kkk15yUyzbx0GzRl+aQnII+IuQREKZkVInSb6Im+62CrCjc7aTntxjyOJzYRfXux
e03R25YwmoZ0esfvRktlFQTnHlimhRnljwwZxck9MQL2C6AG5NsDToyi8DYTmNb6KoipOBcn3CiH
9GlyyFxjThe6nMx0bphWzNOTMZd3+z55gFXGx9eClgMNlacSSJf4l7rCRw5VVXCj4fkMlgdeYO9J
L+U4qiDY3ljYc4NA2tdmS+6PhVAwL7c8zqiuEFxsZl0EjxXGMFLwB/lp76CQ1JFRCtIcB0ugl1fq
8skvsp2tGpLnS3TfzSZefslYRvoEyh5ZWOFtlZDNs7QZH1vA0FFtPo6nbs/dJ9dZ3h2eXlh5kHrc
n4M0YRHXS8rYIVxNF78JWYmymdAdBNdEUftKdKiUTKyFtI02YYpvX6qIdygVgi7aAL6WnJP+BKp8
ZALyUx5uP2V3pxk7/7yofTpxTcl+UQKVIjanL+rgsTZRjNkQ1iNoAJ5zZeOqtcmcRXD2YvWmGmnC
oOJFF71Mg1yEWyAjqa3sMB296RkuVNCy5uKSuJxi1qfN/Cpqg4Q8+gL87oo2Pf9BtFsJPBdR3OGd
Hs1+zdjRBVs3hMxeYTmW5KgGrhnD0SAw5khj85h0H1DNp+y3EfUiI5Z6laKiUEKN1kmbCNRCghq4
6qxFz2+vOyyOb3rbH8nGav4D9DO3mqPuSswVjb14FDi0P/wwuKZVU8y4Y62vhVBdsM8Shq1mgiXf
xod25TLHIjUJDGpoVRS2NGZT0FVFU5LmFpoP+qc7IA6K29+rVJPc9sjT86N+ItDwGYPk7o4bQ3zi
gBLFkDXy6a3/d7B27DNNVKbSKl83Dfl03VzCGCsQQoFt7K3AUPdOlxMQXiMNxTdQCSGiEwnhSWXN
cj8iWP393BgUKGIB56KyyRbWtuInzk0wH5oG7ejuMaA+nBBFwOCXcUEVFbJ6YYNDgUgeVNJi+fhS
neGR9YUFtWSBiyjVl0lD0YA/Nl4MnZ3g5wpFzakO66nh71ylqe6fWI8C8khaac+7GorwEV9icnbf
byZ6eQhFPIOWFA0DmJaKJUhOK7n2uN319TntIc/4jZwe7CUWGIs3D2UCCjz6WZv51ah3iiDaF3Fi
Cho1OQrwUXH5XEC03no62gmFY7NEWa5JgwEnpC9ohpULPsorcOq8Ac1lTNWYfYp5DPDxKyESbSnP
a2wPDwKyALOUJx1eInhU0j82Wrm0pz75CrcDmhm11vXjVmGIIbGtIGcSA6o1WFALps3VMgVs+bvn
OxG9i+IRPBSyBIdf1c5n3GPi6iSkupmDi1gV1YN8PL2XrhIg0ndT/6nTDzIQZ/dpyx4EP/hF6iHh
DlfsOVqCKDA8KSusAtjZkXWdgH5Q2zac/ivbVHkOoE1bEdgFTKGFwAUTy09jEQwnb2keVBFZ9bu1
bxgeC2hd/Nng6+cTYjNfAC3i2jDujOsiHwzb78aX29HCi1I/dupj5TeM5yrbhNCSQUmZr5agyxfA
68kkKG38TqYRkjpJbyT6xQOu4IOTPEpNQmBnuq/i2b6EIVFLF/m/ymzNrHJ1SiyjIMaqhnMR5Czo
e21gq/YdaJlikGnisupwNlYDxWPBWoHn16ajCwo6r6JuzrnF9T2BXe5EVnfFpxt56sbpc/BRcT28
9mm4ZnIkf6AsklkgwMFvaRmxmWzPqQnS9Njxc/iu2o3oADxNgvO+tdl0Ixcao2hShJYQS7UgwvXW
qN5HtzfP8h99b4ijF+yY+gQvHNoyOyBcfp99baTaH+7WP9OyMIbLVM9I/iDbNohsR82w94Fv3/+X
vdGt4Y+9UpoR8ano7ausHny3LnqW9yzF/wqKTpseOfqCLNEkj+ZsppR0ghdhhuqWA9RQihAbGve4
F2xTFchga7qWg06YzPT4Rj6RKrp6we3q3uXvehDClnHJZF4PiNucvYRFUFC9sXuYLs/XyJEOKRY2
AP/RuNsDoy82xwhlDN3G/TJ5UE09EHlWaNXSz/BfjXqrz3PMUa4O5VlZW/lxdLJBzqLPZ0EqqXDF
InMz4FIngLi7vNaEZ3uciOvXt34mxRQ/QKD/ykSw4QezbbUfExhPbNWmw4Dr6iOg9xqZdePNowRN
PmYwXkdD06+78sQP7PwnQmvRL3Ez5mMK2C0wC6TVxqZrRr56lOFLz0qmDeagewUzYKcj6+c8AjVg
A+MY+KI1T4kBEGecEL74zfHydY6qiKNPVJ306obXS8fF0g/6kranA5TaHg0P0FdfuRUeXCOh9ets
OD1IvF5jMyfozDfVWw+2aLovL2EsjCECo1eHDn73gDn5F5xlZCP5wsKUPlXrvNV7/CuynefM6bD4
izpAVC5LiXVMRX90K/OXCsWxX/Q5RgrFKaLAQjQI/C3mylri7D6x8rvdv03Oy5Q2C6MCt8hw7ktg
DJwuFUxmxDGX+dDWTfECSPC7qnTfm6ttiQsMO+cW3/CfMM7yM2qhLWOSgPIVKF1rOEZmyF5Q3BEi
Gqx7v4OdA9x+OydslFj6BwEYURccT8NzRqbM2d4ZtAyKT3fv5rFNgPkHYISHawwDFjn1H7wyWltx
9XYimmlXJycEySJ54Ac7vmTyXxHQZXhhcaQd4Ar9Zh/OU6cCQtAED6BYjlvep/Oc+d5vfH6VPygt
EWc31NcGfV2XjylGP40/JoRbR/vqh4k1i8tj4+0WWvl/sHIWWoSIe0F4JbdiOQCoES9KOt2p8E/U
jcEDdKSjfhHzTMkCCnvqhHk5EFO4582/FVYOCKXyjQiKtCqAnFdA0cflq00/+6redPTO66XRZw8r
sKq+yQZFneUA7DMnlaKE7MvMfhs6YDwZYzD8V+HJnyaipy433oiubezvH04wj0Zr5KnOC0b4Z4BN
UmR2ux4wGo1E4ibLXxN5Tiqd6fWgiMFWeTMtPK4Fxu0Siqw2hAPwnSUG+Kl0AICLjM/jsHlda6K5
c2XNYXljXAD/hQGDaa/JxfC5zyMLQyHwB7oEHwVn9OLLsYjMSDJ/6dH+eJDovZ5i533sxErjdT+K
yh4dUwMIGZhzR/O4DnHe2LbDb4kU+H/VyNsr/KEEo0UstrIeqB8c7gPyJIbybTtpBKhrU18myARI
XkGPa6c7PdAynVSAYge7TpNLUUbEu/10hyxH5zvq7KEDITTnzODE0EHGamzK+rVeuqGiJlOIqUSd
JKZRfHq+63x2yaBadS4vhYOBvInxHX+dQXjK13dU7vLtPJkqmCKe7u9AIl24/cPvXau5TRunFpim
3vN/6aRMGfAEsZOJf8/6N7r/Dt4SigibL76jNLweO38wED+T6Ulqet737Be+BUUogNErO3ZgrNfR
3c9trzqJdGV4VFzRxfiQGeLMhKzvL2lJIDpgg7LL8SJ52quoN2s/5hrYt5OlgCRNdy7t9AuuGa2l
olMelfBErW9YhM7iPa+ymui9Td34MxP+W/FCz3KrZcBrvA+0SIUnSOI3rhx7nh4hgYR54Gt+NyaY
hPBr2GTiGpGmGWa/Xwkh3PC5O0Z4k3Lsqkh6vxWzWLz2ui04DqRjlfRmgpby8o/G7Pl04Hj2d/oJ
aUbs9TAtmFmvJKvLpbWToprm20zd1LgmcSuOm3Isk8rqWs0hncmZMqOEQhVow0EWALm0pELaxF5z
tOoEGtp5H9WKRIsO4EAsKJMcXrwyizVcoitCoQhorFXJE9aB2GXsbu4aC66/RODt7pCTfWdTNS5l
hrsuVzrKiFqcsrUbz9H0syYKauiGZkvt02Q/VAJlEIPc20cBWRoBA8Ox8vUdt5ZpdLU/FlIikiQ3
clIQedtg5cnRDigMpr/hSqiuhdZK6gAei4Xe6apfX4COIHFxT6910+oqZRclHtCzq85GHSgD1WIB
lUCqIWljhSvGo79wA2ye0x9G9LHPFQn9gOvK8FJxeyJTU8e7tbbdxoFFhVFAEhHrRmjpKcqEOFtR
ohexCwF/ElKkHX7M2I8hRahqCHRPyITJDXLDf7OJCBPTJTjJbGOfHBkgNnCfaxmSLRzEh2cBGISX
3bmU8WrHutMODEXUQ2KrF1CneudMp7kUMm/Yi3gicZdPu8BeVZUX//gRW3B0ZaLWl2cVugoVlFmm
am7jlXbE9lNz5MzzX5Pw7Pqx1Q9KOrgOoW0TUf9ZR5DPPSD5G6Cw/RRb84N9rS4qtNBp5B7c1igD
V5BzUSZ3qOecnmS3PH0SlFfLXCRR1JxN+d4SINxvZpG//H5rsbENCriFRMSoDlwiECxeqkWVeBeR
EToRQDVRjAT0FpxZJxyDQelwblKvXRvarm+0GryaGknwyfg5TviXZkvGFswhZ8uq7h19SxCv+pn7
B8po05FrL+29Z6vtIMcl4FkXXeGNy3IhqCFKvhASv8hHWgVTAPlPjpchWHwjCsKa0aiHa4ozmvC6
POI9uLHl7DNDZ0Peq1LIB5DOZ9LhK4EcSfGpH4hRf6kEZHNS45NRonUdqX4B+jdxwAeE1gTercCr
7LkNi8A1kKPyAWSayPLZ5VHgU1GQWrXgs1r7+W+Zu8XEsoSAlo1quiRr690TZK6kAEiE4WSYccEB
iVidvlvg1Qddseb9NyjRwiZs2FMMbuTfVOQkDgUaMnTUj55GmqD977Mo3NoCEdUHNO6BO0/HwL35
+qKc6Qtz29NhWmbii2eWsIwMe69n88lIljMp6NB5a6LU2sCkw83k3nu7vsielOmb8ZzN2VZjfNqj
SWjD2oYgycRRKZqoG5KZ8xWTgq8SpdhLx8iRsArw0OfoBsNlrVfzAjwcf29Wn+sgBPzKoGF1tI9x
YgR9OJXmN0sAUn4uHxKt9PNGplicM8UN7iIr5hiaRc6i96C4kX+v511/iMDrxIpKmnunMlwzYJ0p
oac7y/igGI2T757Ew8t5rf93phdd1N7H0ePQsFNKPI0FKp1UnE50aElYfPV9zloddTSlUJWPBbDb
liNHloe9Ss5gXQ00s83B9JGPULf1bRddddCwqD3Q+3e2uD9XK8HDH/VJwfK5PoouCmBzHjPZjk3U
v+IsQ71ub+NBTSl85KNLJTGgrFwbrdHjdkHAPfI4Vv/kXR8JVUYqknM3EiyPJMjdNDL+BYOVS2uk
QMVjdmofnhmDTh52VfBH6gWLJaB4Zeca46+IQf0r7QyIZd3K5Cm+EaMIg2TacOjt/I7RJq7If/DS
TlBSHDS0+AWSFfQ2lcOsbPelH3d+yPx4rjmdBYHjg2beolgH5xVPOHQuJrFE4RcsIRa3MGHN8dfn
MdW0JHjQ+Vc7NHFM3WkGF/44HDfSibNiLlAB+k7vIcGhvLrL7XOagQi+TftC9vijgUdwfYaF4zpp
KwY3pJEbLa8SwK4XeBVgW9gjaZl4NkWgR5sFGqdoZicSvdiYPLJ2Kj3N/tBjl0bVg8qlU36AIX/e
Qp2Gw4QV8JUeSgHhPbabsDF0FWPyLQGrpLl+FZ9DgnRBGWs/TGTtF4uu2I3hjNpLr6+GiOfmeZK2
rKEyjAXrE4S1mc1zN40dHR7iwz0zRthMCWgagYy4WeajAA9Cs1l6CSxwcS1lXkGoHbvIW/iPSyPg
Ea3eSeHlKWeRO+c1+C7mQs5dmUcHtYp7lJjB0oEkW82Y+0WOhni2zPpKQDU1RX5pJQCsJZD+uDlC
nD8KKyxvXT+mG7jJKZwJNHwbAQDrhVQTSHybjsZR9jYksTPpcJjtMT83Zl9E09Qo8+FwZQ46qmK8
DMta8/tY3EgszHnuIkvUk6qH4r6VhfODdZUWMinUOZsd4NdyWRbtCH4WT84SzE1PskfCnNFmaw4n
fBJB+jZ4NeRtJeECl8nS3v6ADKxlxnb1ebkz/TsB6SfAqlPHEZlfoW8QkyUlM6h0XLNFGd6Wr8/t
f/c00mHqacs7zwSrVpmlM/MbdP2hiQugq8r782hb7we/ronJn7sZkbCy5EeIJ+OPOl75LJ4apJ1I
g3udCud4qmYjliwx+1MHwfEcHxPobkDDqjHW3WGteUfRcZtAvR2gmB8hXbjCpCMmM+0np3oUGw6o
JscZ97tbQgAojwbG4y1AIN/Sf2GGzANyacDtbm9anE4/49JP9LBJHAsUeOhLWeFlBhWpBkKiYpqB
WQiid0cv/Fxi7+Haf+IDv4VIYOh2HKmQ+FO+ZSVh/vlt12Na//Afg68bSsk0B2oF0dczKGCittCg
wU8X6ZF/60QEjM0UoURSKdpA6q+6IKdGKMfVPGgyYd5twYHrCdCatSmCsC3wc1rwtWCCY2j8sU45
MLt3vqXAe25dsvFU7n9L9sEqmvx/TFbm6ao77eE1EOq3cxJDtYlJ+/esSWGi/hfI5m/3jcMEcmUt
43fCL2apmb53if8TJN1sXPDnLA+oBSCMv7bJzHFL/bGkB78tsQaGkaGR24HHqBsasxHVgOa3ea4g
bDUCytzYQSV3/1x9lyRLmFaogOdvv7OLi3G5opyzDhXzqDjQkQyYF7zMuuJL0j3QkmEjOnzc+1rf
QtXUygfxAYTNyHB1PlLWhiDzWWH9YKK/JOCWjAUXMTTx/DT8fB/+PyuzXhYks4kBgYnBT3WYKsKc
qaf/iP47wGOWD6wcZDAMEW9DdO4kITQD17Gu51LnnwYv90FGuNMn0YdnCyVbeIDgUvxkRuY+l6H/
O85q9q0Ofd4gibQphIJZ0p1R4gAcct7/GdEP0jC+xs0KK34TaTa/ib5cbNK26q9R5LO66FNsKPcD
6mk1KLTCxkIQpMUEjyLsDy+CSiRJCRZnXKSNulAEBjo+sSqmqhoXL9GylnzNvEOGCKiJ3+ZSErop
2aS5JnNSjQ9Rvem3kijpo1qsswHzo4WVgrrFCANpo6KNeA3++2dDujs+KYzt/86IuqqFSbD6cth9
UURrz3/BHqYvvQYpVGhDHJcvWhPgE7P2nDsFGaTbwN7fkVXrb8LuzncsVa1KG8cvle0FNGiqPw7v
Jy72J2+gma9HT+bT/79WqGCqkKIIam8TR8SaTzMzp2Uf8QyVogOTXWWJCzP/nyvySLUB/ODCanJu
hm4o09ipLOYPadbVPeD7EF43JTUFXS+Zzse7kNU78djS7IWwFGUCdBzl3vIb5Ekp0AuwnufiPrP1
tqALMScJghBHqtSXy84cFHqZtR/DnBH4z33qsfv8lG5OEIaHFGGu61UAHFGgTT/sUngaCbK8ks1M
vugAKjbmqxQdZa07zWiSSiBYl2FJ0ifz2l9y578lUz0f0nnOwOi/RsKQuDcZW/csVCKVntuCOmOZ
+CcpY3eHf3FgJXEUB6M1kIamowuLdbPaoTVGRbgYVOMQYKnRTQ84xktRz6EkMY4TOmxW6Xh3k7Al
YfKBVx/9ftPztsdmOTHe0OAda5lVo+a+0e0Sk7b2aLRxmkc5MELgI4cX2T6IW1nx1yDwqbHepdpo
ZWo35Q3injbjSzNNOIPGl4xUm9dkJTNWtMX8hxBqhFswlbdgCVNGs1s42xKZQRQodzL82W8SThK7
Rj5CZcTJ6UJh+8VMyyKUeL1a9AhbwJILCdl6TbouUtVFMumQ8vXq7l3HAtnLOKCpBJW5UriYj+QB
Aw9fNqlrb2MnhJV8DwBYrrvr1eWIt3EfApVDqqI563NJ6itd82tT4yaD5ScL83h09Bl+wXLssmhg
ocExV8j+y6h9npD2Wjscp5dkiOaVWGxvLQyQgR2Z5zDFw8yV9otLFTmapV+TLDTLb+OAAQviD3v1
MeP6Fvdrkt4zBAP6o0YuLS2zK37d+oV6Bt0aWXZJM5Eue9oGmUFczfW3ENNhnYYfrv+iLN963wDE
XMWX+6oSWW0pcEuBBitr33rs0o7a9K6LUwQVOnB4DnT0y00jkD8p0jXGtyxSEDbAGjVg84PVuCnI
0+cXcss4lUSCFXz83SWxsI2pev/0pWiTGsukjaMEyhR/SRVQyYx3mBlQlmQ3zY28fOGDPyg007Dm
CWPe/8HWQt9iqxT1VhRGuHcTOZL4QM1YPnibA+RVsIJaLfLMs49gtE6D9FLMIrw16qy6Z9j6wCB2
xh3itbvnut/M8p03p/H5nA2C4E0uBjG3oB2VqKEI07Vx0YVe7c6gchRIqg/W7Vq+tx6JvaXx56hL
B3H+Z385He+thHtlxWqAnsfochE9uvURJPSy0Bd8Ip4InbynuMOrl4qtEHjGEXmg9qREVCUvBa9L
GhF4XRHf/ikowRTEpafIaz70Pyo64VlPK7g+hUqIDFXy4NaOWVyLiLSaT11k1JTdjssLXywJxThx
lV3bd07wK7jmHYg0h5uHDxyAknB1OlequEfyN2jtzA9IfCAuiE7b/ImyDpySClF5erKqv2wu5J6U
BnFCgKChP/OJ2YNJksx1QoFMWK2o1cGiyQbxLPiyWTTt82PGw7xbKjcjdAtdkgKaAEHmgsj5Nz+x
YWszoIrA4QhTnq+3bk3yJVwdv4tR+VWvWF5Rxx0qyjCp7Y4tcfirXLN+Gi1mLosKQgY4AV9UqH2w
WeFmX48C89s5SlMoQcy+LhT0z/sPx544EYMRSnR5KefTPPA7h3+ws5cse3cvoBz3tWZDTYtJxoR1
STRsJ3UfpEcaMKvVgyN2Jjf6QpKry77WJfgPCeB15rJsASaU67E5cXkMfq+7bhoy/xaxybdfg0sp
XRUVBY7GEJVaU9t2h/hzwruTrcf4HOBVLYEXXYlKOkl5BadUYlv94uZbGbHDTisnvy6Vf37ib7gW
+gdDTeEJxyipjf4I2VSSlwGLE6FDPabTQ9amssGxB1laKLV7TuM60oQrJ1pudMereII1HztnZEfQ
iEjk1cJk/bNqYj6FjG2J4So1cntuUvwnyD5tHSofNeD4cC6RVIYForsiIIu7sul9kVBGpNp6hf4T
80mvUygIc+AcgFg0qqJUjnoetYJaS4YT6AMrRV9ftQgOoBzuFNP5Jj8A25Ufn081f3JO58xxY2+u
tHgVcjzX0c1oPKaW6COe6zRitov6KZv6y4uhiM71/G3yCcnmQdOARwlXCu10E5m4HIi8O7X5BOGx
9DTf3ZPtu8KXDYEcdmY3k237OXBm0/pHTedpqZwcFUoyD+JZqxbHv6QN8UEngNE0nn6x0JROK/WB
1vyccFbHqqMjKD1aa8krCFDQEUOcuXw3Ks9kyKdTrpAfX0VEUbHo/eKvqHAia9W6CitTabYi8r6C
EVaODvZc+ccrkm11ek4KaqC4+8h/4VeXJ64comv1M/kZPIqbYzxaOXqb5Ji8fPFoXty6hUgQJbPd
NEqST1TwNxvymidXtwQKLD0uVO+nM8ALfPUkt119gypwSqt5yMBUbpt6PkTSoEZ3ed+f7BegRmMG
ipE3o44K5g8XqgLknVYJ+RKakZ3R6QwgUuLFjQ97kvdYsHBpzPXHUs/MDkw9lREGomE4F1Wm4L0c
FysYdaVJepuv6dDQ4rigFELyfCeopaRAMqXfTYNwrnZWacYN6b0iNmyBs7FBvYtYCaNVmjxPzv66
8+3Q3OrwOgw83gC/rKvx9G9L5hNydT6nhw55BE6xH1qot9uri4ZpaeiVnZWIwSpL1EpA6hKtBkvW
tfejNbxxMULqJtMFwc6aK+iZbwFFX8BUKUHThYOOtR1LsVitQChq44I+wSyMDaEpJiyxVDsS2DRP
evrFets0uev/1vs/5npI6r3F+BqrtZ2U1io3GKiBlMY2s5GwL0bXbquFdiWWEQOq/28trjS/h7l/
PAqbOXE1q9UVg59zYI1OeYqVvAwWnfEfqz8fekPUPwwKt8Y3+xbLbdAzNJ9Xf2P61C2W8tU1T5eW
3a20wxidj0vma2Fqm+5UhvGa6/YAJuTRLNU08U8wtPwarO73IKmA1x4PvE8LPAwTK9KiPKOHThEf
VfdSEaAePVT+jFr+bsdUyHdaIY//6z0FrvFJzf4c7PJJMRxaOD1d+Rvf6mlnsTio1inmcXmV4hlu
FcadYDDig60kR/p0nB/u5p3Uf6ISbXj63JbI5+C9/GsH74WrpTGYqbRC1RkVD3nCEbtA/+r/vRST
zkglXJp0xSmzPGgwGXAMm8PR972BNwjdOyLUL+lr1L/WJs8zdVGIdUiueaotRdvRbOktX3ldQoVH
XtyLRla6mi8zg/IQ6Mev5zULyfu+GQlSUCFQKPcOQ25t6VfESvExwLbcQ4hDxNZRXCEaCAnRVQBy
VBvoVQMng2syFBISOY9TwJV1RPBaXqPmReFPE37vx3e8jWWhFYetCHrhmDFJb4kgndIpVNoZhlKX
PluA/t0MK8YWB6EUvNIZxXtV4ZBxYJkgDzzj3q2MPM+gVgf17fzrAjqi097+q89RKX5Iy0XCXjId
NCsC8xsaLs0cpf1gFU2cdHNGWGva/0vZg9ix+Sa92SvgvPpeQpv3Mdgg1NS3bhEuiaDA8jSjKf6W
iK5TKKOzHqrZei9q1ZHKl4keUxVuyyNZi0u2iDz+4QWgw/qk7nMIsNc1cnseEoEBdCDPCmB19Cuo
7ckOyGX92YRivltXAlL5Ank3ubAbiqAROnftmO4znY4EdYZKviNXrKYsgL7vVBsqIv+EEe72y7fS
vGdcvBFuqjOg11FNl3Qc3g8U8a4iyRvRcxZwQcGmovGx/IY2pQMywBm+UiWZygah61c2jtwiQ00J
j4vjcJxoECZNcs11MajmCmcn7dF8lOTkIoIn9N3skBd4Y0SRY+MHX2krw/aZKp2K4YF4ALPdN8/j
Wu4x7Uvqevjd7tcTF6pdeJmmlQ+PG0wfmD8P9fvv7RezchpVjTkCzx8yOJbXFLrb56PmI7h9UHRa
B/oLG+wTdqtnHHIdhA5a8lNkgdYPRgn8K0ikRRO/IjomncXcGAh+8L21ngg/yR8ukQHNSigm33Zl
uyqABknKH+9GZP9j6T1j5n/JMnUcSsXYkKpth8Gd2kgS4wWS7jurFM5SJB43JVlHF89TH6u95q8V
Pr6h+eXZCStQsjMELHvFZYyCh8JVpKUahKTZ/jwif9MPAISOkFATlaQLLIVSfM0XExqe1WGtiUUD
H2c1aqbTvBZVr2b4kmDKs9nfpeSHh/C2Hswv1Otj/Du24Ag/TXYqY9yvWJLDtm2seaMtTXTVTC9q
yoYmY5pJDwl9NWt52x93DuCkZFefKXE12Iledg/yY6zDTCd3fN2eVC98UMC9zb4KE0RcWWFwgn5B
WdQRHeX+edXkeNNzKREQLNM+/GrAxF4asYLc027NRjSlDHlHzBAm/IUkeKqDDcVAQ1n0ADI5I17L
th5Rj/CEBoca7/SVKGsdXDhZgwsHlKdtsUnY4Mx8o6ylCFCP6Fd7YaKkrFUUUaONiWuNs2dHYwmh
riWtGshJAgvrfPabI6lXK2x5sDWLqtHRGqkeeVMxKDrf3+UXBxqE6bHF4NP81BnBSliCanLV9tDX
OQ9kepPV4Lcm22kX+0IRHoPYmyHPp5a8MZIOodabHHXx58T/acIVRTmuLQVXy1mhkWlZ1+SpPjkv
QAC6ptxq8U3WXd2+Dm3lLDRigvgXHUiKix5CWZLfYPypM/kaTPQx2iMczAKoazORFrYGjaH3CkYM
OO7Pnlh/VFRIhKtP2bm564XnoHdB2jYhPwlSFYizIL2e9vGGF1YsHsuakRcDAyNC0vmTnT0qCiOm
V5/YmWem+0j1Q/HydhuSPw6pfwd2jyUJtF0AT39aRHRyNk4VsojfRrzIwoWlucxTNFpHj4F7lpeF
mavGI2o7bP9PLwPER8AjH6WUdoLSr3/8rj2ZXjGLD2QaSZxQ7KuYse1lprkxr8vJtGKVBIbkMLSd
K9cTXfFgbruoZMBaxEVQXxG3cyCbxxnJ5yBhDA2pkpTbmTQgPdJodTwC1rPTGdiHz5qXXLloKIju
1OUKaT7xvoJnbA+zv4VGQ+JGQg4tV6OBNr7DlcGHLCA46RE4acAuYC3TP2PFraJIwNhQdkT4ql5k
MhBumgSRX8N1piKy1pjVOvfz3kkdu1zKK4qblMbH4CVY5ghmic5FoXPY/blIY6tpxv94ZwNvvlJf
R1YAaOjvFXHnSXLNC/HMWWfH3e30R7sLI0daR6hQz1f2PqVl+GYbqvGXWPwyd8vRNFdMuKzJa485
2yEPTsRxX6p66ChcAqZSepr6B56tjdGMXVQs/Lzel5LNAsSvkga36e85qPQ53w6lNhDq8jRz2yHV
16u0SazYtzgAYthsOira1YBdTWjF0d61kQiEWRtikwr6RtdOReX1/lsHmdXFN2mZoVB62g2NwE+q
gy7DQ69mnAnW3EcLhDmoWNu6XIp12eWcKlLQ1717Cpcg8OVLgMmzMqGezF2BXIgrpYkb6HRM/PB/
8beElbU9V+8vMzxw+rQl8ECdl4zzxiEPlFZJ600qe98D3/c13j1r8VvbVgtVkJfJlw8yxVMYdV1m
+d4+HJY4NUT/GOyjBFRhfk1MmEylr1K8b7zQX99YHQKZlMxLn+POA2B6yNoG718gQJOntD93Klb6
U+T4IYvgr47ZzpluIlVdFBzs7tKNpqRJSHdow/H4H0pqx38PIz7rxTDnZ0MLUOSShZLC93W32R6O
IV4bEff/k+QqBV7J36D29ZO2pge+x023VX1UEcifp+997oR89eTaAMqzzLduToAzY2Pw8D8ZNOjS
g6/jj/hea3yirpKf8BhViaHONdGyk2g9yj9KKVLvyiM77MIFCc+kST7RWRU2uZiag0fItvshBBzm
l2R5mgGhkcw3VAKri34ORdOkhv3sEzYZD0oDhJcRxODJ8G6h8bBycXGu/hlEd94uxlOA9InZviM7
j0clN1YQGSYWMl3DF2aTj+EAgNljVfJJ0N3FMQAKa7goC3B6h8Xhphq6WNpE70TRKah+vrGLaTJV
V7eCUDHTm1w+NPpdMppqTAZLB9yT/eUsjc/FgBMDLhvc4KmQWDZV6KrHutwKBOapLQGRqiJzJG0i
vxQAFqXnpJjjvudc3PM3dKk8e98KKitHNQQ331uiPNjKfTNkU367guBEB7rjXBRWgcf4x7RP54hY
JO07jZiiAetnKOLEVTPfFIIsOW45VVFbT/Zm13Sy190jfwjm6g2KCdiA09Nw8qTYNqqbC64hMdsM
auopV7/9caCjSx2/HNXP3/83BoVfZSrkj02qpiwvUtNu9wWU+taqRxZSo00ykrUPLoeOdOPNQJV2
0pltw93FamkQ7N2IBvClsic3bpROjMYjCupHAvpVkbUlJWldtlYPruX+8mJOxtbupZn3wmOhUCyH
wXxmeYm8zIZHq9rHQBEcSahsf/Ys6jyqQNIX+qdidxbRhskzKN4kVRjYNgI1vqDObhLkgVppU8bV
AW8tKe3S+qVvOiq2IdB98YQ80wW3Vv/xdGXZzCgISQ6UikxLKQUrpTAQhXqr4SWgSqgDWpLKg3VO
myirXcYvOaL5/tltiKdu5X6sz+raCv9RNFSMMMsi4+dsCez/jqH/pRUfu64eAYh5/Q9NuIYlN0Z7
aY6vBq0KRY32jWVOACkX7WDdz33ZQHbeb1GxJfCcJtE5Hyv6mbf6F92b49OZ1ymFGJs9t+iweHpl
Gtcy5DNxxqFFdKwKeA4ezBoOPQpPi6wmGrmnbYOA4wbSnzu18ajRrUgetTRyw+MbIKmR5oIyTX4k
7t5WYI1ARauVfa5f2cgLFE99HJLBoPBxliOIHMgnv4tjxgtR5Zrgk79BMwhuhbD6EiFhYl9KR6/K
92ns0ptfgF30ZdUOoDuTmgZ6cY78kUWbW/lKfVqyXitXyGKn1EB9XmMZWGzcoVKFo7QROThn+5iZ
VmzEYDoear3w6HJCa38QJImgarDzCav5WqRlhQhHPj8tOHWhv1QaGHrQy47quhGeGHKEy8Pz3RGW
R9PKrvWuhFlNgacbi6mHyX+sN30pOV7+Z2tuxIp/a1aynTPJ9DUuOPDZCGAni5VCJaKN/jdlw4SZ
CMy/YXlRqTcIXAPDb+WwSawJihWPFY77BesS2JKN7eTYmox16GCqli/Ail/pAeBHFua6WwnEbsHi
rgZ7bu7wPpQrVZBMkdsHU3x073eEPX0L3MK+FfnVU+vh3Q26nfRctTHDaUtDulfgJfU6kYXGKAYb
C+qkFvCyHMAQi2iO4aG4zoYW9LdU0rh51jxaexzeREEwe8AjZcPAOdwbocccCxwjSc57GK8BMgC1
ZFP32d51xWNI6xnsp8aaK6yEFuAtX+o5DozJAPkPZ1fYF29nSAyvmF2KoHhuNcgZRAuqztK+kHpE
YCOXRCLWGxzI+BiK0tuC05F2uVRUFgxrhc3RzItvqjOTj7LQon9ASqB6ifbNt4X4W/u1eez8pldS
M9OAU0RpDYg+gOPdB55xARkGjsJaZHvcuCII84TOXbCrnyqu8rOJieVTUBr2U9eCqAx07jXhWfJ+
FYPt488mXHOtxc+J7DgNtV1tcZiqo7J49zit/M7DA8mkHDrRgjTgT4LdSw1q3PckE3e9Rvk2qyma
LkEmlyasLcKE4yI6mhogIKkmzZeVFp3A5TQERetp7TVgVHaosOXb1iKD9Rt6Kau1MfsR4c8JzWQz
wLefYM+3X/EptJUGF+erIk2qPCJLRqFSJNAFm4WfkgbBVv6edShEqNbah90/+Hvut6fy9F8Z4Aq8
tKAlOrQdj+GkDAPMmj4hLa2dJIoymfGAR9JU30D+cdo+AOtSB0gdgIP7FGPTpUVaamCr9IhsqozY
jV+ZoPHv9eoJoNPhNPsDwFn3V3DOHSQ1eRWZVZ42H7Vewfdf+2pFSNogoM0ToyfrvvU0SwNgI3Yp
x9D1SmyUVQboAsMsPmnUkmExE6OiOetyWIhwaDu2svrWiLtrMAS/muocqYeu32taNLOMikxyFfKI
21qVKsfaucmnhoHSv0rYmtg5kfOByGXwCTKeZ/v4uLKF6RvyNvoFlqXuwu1X+kEhVUUp6IrSqivI
JLVIofsgO1TXCqJCvthD6cLrF64ekgy5BYHBBFye6ltYYeDvppolhLfaPwwSy8w1ohR45ZWcxStv
SGygNcCFNB7NW8iZEpEzkhL7bSrwVm/fqv4JwOQtFik4WUczZpE5Bizju5xLUigScZm4QJz7ZxYz
9f+y5mlLt8rLPzD39eS7alzxaMvpE1Bh3IwNnvu57+K7SgWmDVWcCRQDghkqA8FqRZiVKBTm6Rc3
tdiMUu1yZDAnar5yDH/yDbq9AGeVPidq6IkcoDMgsAOYkuCracWFyKLAb1RocaanNoozBCnlwja5
sO6jlXA/IexuNqyWqOPO3LGpphnvWnhW1gP2UFQ2+KT1xNE9L0SEdP0224CiBdzJ2emc2lVOXoJg
ITq5CN92WZJSOqGSR4CSnEteIpDg2i9fyFrU4yZwYbLuqgbzjeJ+R6KcHircJpf4wfvClkgbsLpx
/Ahc7vifwz+CrzTodn5zezaU4rfqIsUz644feae8NBo2Ou/hIpeJIKn2646fZL5wm5W+Cug6p47D
0PEckJgP/Qr7Vbmu4LcibrGYU86plZorrKjXnPYZ2oM/IcNSirav1JKV71ywvntl0cVG4QA6Aubk
szFtvP7oK+oY0gPo6ydpqmFNEcCPlaWJYs6507OZMM4CsdRDP1u6iQmzyvz6HI+lsv5IqOBYvhEt
bik38Nj9lCHQM9Fi7WNM8E8jz+j7cwvZoGEtLEGxMNp5lc5EZI/QOk86+1/+Z0gB5iYFK3J2mz1Q
PIg1jcWbZ1XfSidvgcJaGY9wJCUeqNhD7cNp5AzGrKF4EZRpGbMpZNHrCd7nQnBRN3mkiEzg6FI+
mxITUWV4thjoM4kOcpl0elC2ntTd+uAAFyaet1Ei0KM+fHdELgKjxPT9XSKIQCG7f1QeZHKfu70U
E127zl5KweZhIGjb6UIeNwMrfe48eP6rieOxlO2yeLBYnfBdwGeM4GyF39Gp6IWkRdmFljATG45E
6FtlTOFq/UndCVJd7/3Q1JPPHKNC9cjnAfiILUsGfBdydE+FwXyvQTvhuAMyFEHh7tA/jsoS33zM
+xrY1R1KO84UVGFHaMPSkTm2PzFpHeWc9XklgcvWfyDgHeSo9sCdk1dOphwQSv++dbtDPxTKS8WM
8Nze6XUrD4ezAUiLXNJAtqtNh7UV6nrFapX9cHoYKOsj/pyQg7k1HJ5jitijYk1QeAIEuhgYqXoC
bVWJ+g+S8IMq6ctIPWHrmWdhPlHYz3/tIjvwceUL0P+et9NsEGoYy/8mtBKqujDzDT88CEFA5a2H
5JCSr+oYa95XctJGjhpyd/F5CbZ+lDVbT7NwHhPgCwoBxUg5NHKSYPhK/dogA/KUGar5My6PeOEp
hosgx5GNXRpOcftl1RkPSkkda636bDrAf1cxknPQcWz8i5QCeHRn7q3kPH66US3bv5x6cdbCdC1z
erUMRdDF6+Ba+ADa9AvP615Jfwq3wH6l0bVILUVwYw2KJAl+Xgd0N/4dvd1TF1Pk2Uz+vUkFV5Ty
sAyCqEovH0Ch9zsIhjJdcWsA4TjaMN41VkSXCPV7n7kvxYTekRkqxo1h0lTq0HXCUxpc43RO+GhA
VTYV4P1qM9dfJb5fBsgzkNGv014PloEqfNWHpCmqigFmxN9ENXr7BFezqlS6iMEs0zAMZK8nGzDF
Dlnzl5SsrD/8RG/fNeLh0U8nEjem1gurih3bmovTE7feyAuAWSadS7FRbcKFAPXxKdA2qdR7ThH2
BQZIMJzJF9xkm1cXpK+bhxxGpvwjg6Y9//IUjFhTKcV8u0KRcdIZyaogCK1lGhI/DofOCZPkJBCa
foRGinlo+VkW7Xrn1SXZS6iLwejqxqONq/bb860dHVtdNM3OeY1SptzZD2GfeQ3eAUstZf9XhIFu
QUnAHflh4WJHPti9ngx3d92oNZD0P0c2rwDKjxcFKtiW1GMhIQA4rpD52F7v1Et7GyLf7KwSjv0E
wFpkAeYbOUQZfTBCphQT/G8Lc/+i0jtJ88EH5MU+CzwVYAYE0X41AqCYgbP1NkF6TyEopAHO/Pgc
7vA+mcN7eIfVqrZ4y/lY8YeBXdLWizo2A6aBTg+MEtTGn0v2fox99cZcK3CPtXfUQUUHWmTu09m2
R/joO7qX7fqNIxXm+JaRBbwzBYJ9hdgTgQSxa+8SnDIHBXs0+nonpsMRb8KvYE4A7TyeoWpNUYrz
3/IGFHnUmNi41jIvJS3mwscw+s3ynjc2LAc5qpiaHiyG2mu/uKQyJiigbfrL30F/LHYwWQ257pzR
jRoxL7QnNqWqmIQBMYo6Tg/b8CSirLJ7sqaS0Fu7vUcJyBdA5oJHhQFwrg3IQjeN6iVqRISu1E4/
11NkIl3UseY9+aqcpORXGxF0rc8s2cbBtNkfDrzA11q/lIZ9YFr4tINpf6qx+skTHrNHA5sDJiQW
OimYMbxsZM5r37fcJ09sTv/Kluxstt4TxlvqvNt/RVFu8kbXjnbQUbyWJK+Sa8x1grMKsOCcATbx
gbEMdCV8cNJKo9Ec1psino6bbyTf6wzdRljmOBuQfZaRDF4PYmPVPYsZx9K8ijxKYSjkNEhBhyC3
wM/YAO2LDPdVtrH2EPUWCdd/FU+tNdTITRNh9zXvKK63gFPiIUk1FM/ClTsPf3cRYyQx8c2Mukn4
H2z7sShXhpUjDttCx88XtB1/oFoMuCbFwsesD8IaaSt5kmKD8W1cwMOg1XsNcCWSKq+bz+ugFsF2
cBk1K9vdg2PHVlwtOsg+yZ8rrIMJ1fPh8DaTI6rOBkn+0wyWtYLRdjgXAr0zt00wG2/rT3r6F/4Q
hyUJiE8PsVMnt8DyQwM48ZH4D8daflMntyp0GrSgZyB7lWO7cbqRKSQKSRbr+gRl1EvpHpIXEDCd
msbuSWQa98DyDOU1nEKLcCC4c8AWgV0xGqqRnQ4ausclAOLe5dV5sPJF3ygJfqiucHmjkI79XhFf
pFSQF5Z6TH/9zZ3xZpSOxaKxB+4/eDF/GEbU0FP8HN/FQ/7SAvABCH1WqVEoTZReUH2STr/IITpv
DB/77l7Fooquw9Q+gtHqk7yQVItY/Ww/5/UpJiFzMplMmHmRNU59RqdUoIY0ZZ78/DEHxuJnJnlI
2JoqiI5w93KlXcimBGrBZjtNfZhtFd9EGw4mhYeCINL/JpCTIlsddmDl+Qtk/1lKDlTG6H8WPk0d
qsXNPys5ZVBYZTA8Hq7LyBq5vtcZ2f70fwnwzR28dafs4ROhxk7Ckt2pboLn2sgf8/9KsqqpWoem
uBjaUcMs0EMBZMtzZ053Ury8/sdtrCI5yOsaaanSvcFzQ1UlEUwFeKf6k/RtE6BHxiTp4elHnCUe
EWFN7Jlv6oZTPb2POIE0837LNntRIVlszNnhpmArV/Dse3SPsXpZj225weqxb7eIXQnc2qdNTKWw
4A/xPcveT+ABJF47WzFYw/1jekzqTFYx2eI9DHVHJWbQ/8IDTsxcN/cddcYueO6Wnzo/8Ouj1LOY
GWVOFTtKnSmOHVzfyljehqYXuMyE6OAEC1/bFXbd9Z4BfpsYN1C+3rPMk3sYgetMV4sPrZs8+jPV
sKThVCDsQtUOmI3DiedClX73qc4LkmwHGtJsg4S/LrvppF35zx5F3QdJX2UH8+R42HmYVCt3oflN
jM7iHoskx43j4QE8GecYvLF7IUPgmptDQGODLA5x9DHFu/Qa2PHgGINmItZIAPma69wSc9fwHGxQ
kM6/7qYbX6/6Y2YAvVskmlrJLS2Nm8HxrS/Rd6v4k/NSdQi6CSM/KriuT6/IfPcWofpXOb2y3Xot
jKPRdhYQCl3lWp4VSh1ttFzaculSPsBbFYrT9Pb9FAns5yPtG7/7RWxoH0YTxxC7+err2hjxFZlc
qgrw/czwNywAQ9qyX2xO+EneTH2DyQtoTolVrrml9tTgNEO8HG/G0qxRneiM+3SdVS1KZFeXCsi6
NXP8VHK5Z97tI2e6aQAbe2b/tUSkDCgCmHYi6lgKBha+dSGrkF+GuEweMYXF/No9NFnN0rzvoAGo
ImznW5qtmYp8Z0gF5Er3aw0egibJpQHOt8WUvmjRWru22Y3ib/SXi+zkGnQcC7ayD4UrDaRmLIIQ
mYtD+sZbYlsqncUQRLsoh3FA5uHmKbdNGbz0R4zr0ldu3rgPZE0p8nnQOCLWVK9ALinRSqPOL3uy
SWtbygK+zAqm+lQVx9h+a3VPsyoHCvHY2ggiQ1kHi9xUmu68t1dYu8q9Avc/C0PR7lj+u4mXnAZm
R64rxY3X0zs49k6ExYruSG8Kw0gON/5FZeQZRQhJ2+Z7GevJuK3Gcn3NpEQl7Vu/vu4mXMqERJ9J
gKRd2pU6daZfbv/XYvnTO3lSarY40LQ++gCpAE+o/I76qQVx2q4JN7YVqYVmBdrepCf5v7KM/Ahq
LZVAsaxN5doG5ZIRe2pbz5yEDyMirQXakNwe1tcet2vKnxf1OA9pG8EVHCDWdBc2X2PRfKEx7dbK
rnUms4MZwMtRg/NxD6XBQyRL5E3RjWKR9zKOjyb41KnyIUbMEMhN4xtEHmj5Gu12qv0Zjf9KdERO
5Wx1PQp7GsMRss+KRnilqYHr5LLcrRmypu5ptnXNC+imEd711sM5eBN6pp8CoP9tZc4ebFm+/Q5T
6rep6GJgT6OaZiFLvcplNrod7CWOG+eekhOhAGzLjVmSDqww3K7oTdYIhFLOIHG/0hW65oYAbdj0
VxENQonL8hikCwtGanG+RZfi9AMIO3f/V6QFy6yytyP6O5ofyLS2ulUQ/3iRzlwBG2yku7aK/D3/
s9kIJTUURDotC4QgTHl7faTvEEToiFdXyLJvUAG2vCiHJbGVWR9sXxCk8m9lnWwbmDdNAdr5egV5
vhoGmB3sFVfo0nf84NSwCtxuDNV4sMLzzURZCJ7EmN0Xz1mqTqxBmmCaFXRLnHt/k9RG2W1/ylUL
d0X7LUD8ugvqFl0MMg6IHn3EFxp7vxTb0BuqLVLwwXzReHgEP36Mu6kCUmC+n1R9TTcUZ5PSwwvO
p+Dvf+1xxk8w7GXw8y79YefGtGTQAyTva63a29zjbHrzY2gxFVrR1947E9P1ULqvrukHSYYPKmXn
ZHC9uKtNKWazcNqpLrPs6dCicvELlYL7Fuz0YgnOegyA78k6kEmnaAk3lgfchUuyhj3vq0rcYcX8
5w0ho66N2vqrlzv3+X+IVeVHm0U2puSS2a/3/evZ8ognMwQHVqeyrv5A+bJalOVHSKZSzj+HdPZG
5cqBPoaCNtSIzTjq/JPx48TCcfyey1ni0kwQeTZXUSUovc9S4+9+wewuEp0n+TiNk5c1XlRWhIcO
QK4Yj1S0PFLEX2XHFzUH5vyhZs5NAGjzAhR1RouL5McUbFvFdMuEfGEL9/sWIG2k5Pk3cMN4knc0
FEHmgAFC8XOXab8liEztAK/laJU9U5czPtV7IdCTHq6qMwppAVLowjVjO64B5JhGTGy3SUVUZWYK
y3sNVnOfFRCbZH6hR4gDEW8HuiQHU5hFyR5Xwqrb5st7QbonGz8nSIHUh3GfEwGhS9nD8evAfYHY
rHUmKZGIuAJ21Z0AJnLe7XS/j1pFNj7Ldb6geMDm61Hmgm8arDxNg5D3iW4Dahk4ZBIbywlCsS8j
8gd+UeaB439IKy3bT0AEp3uPumR3BJC7ACNiiYVopCtsWMDLPU6w96+PgUVF376SOBYcpcHV3rza
uLGp7WmQR3xKgUWmSs44zWdwFMUK9cJ6UjX1FFUzTNDT4v9k3NESXRrGIj2GRd/bd4AvwYDoQvPf
oBeEXISzkfRZ4DStpaTrrQ2jTT+YC7ROi8Z4cP9bXXCCuIautONYvQbjaj/Se0ijyli59YBMmVne
jcgIOCMs/7WmxeKcNLoj62HnB9eYM0ThOZ8sCwhHX8YLZXudMQgBLohi9UICS5dXjYGKwMZRGLk+
/JKdM0qvW7Q/XN+PEDjeMyHFP1kJTA79+rUrOGCL0gbFRoQkbjmPlCEoG8P4rB9uqSlL4GI/TOcM
3NoEA8KOD68L4/pY5yhBfZGsmnTSOYfyavm4olfYWDZDev2culYOrU8c834qqxLqKaIquiInUPdW
Y8U5q1S68icMyYpOLPzif19A4yqV5ietmDFdHtTqO10HIgn1f/CE5UXKvjHYkAB80a6iBo8W2INg
QxF/V5weXCC1GKRd/RKojkXcSfMxu3wKxeVMHlkijqtG5LUckudAlrzXm0881U31hKLpGivyyem/
x9YhvmBNeT7CMHNUJJ/GMo6TH9lVpVK3eV0J4ltiSaTb4PYDhCyHcPoHAvjOfZ2V3Vc7/TFzITiV
Ft6KIBuF8fgW9Sd0wdHDio7XLdakzFVJ1bT5Kirw3XwO/CjZi6viFCQWjT0GPO4A+edVSDQfzkCp
4XRwOVJfNIxEOQUT3BHwOw+CM3NINF0LfK9x9PSxdrpFuSxsPgyZN3eP65dME7cNlsmPQfKLh+JM
vVscKSkjkK/fbfdTV1StND+oXKfuEwyDotTfcYfbhj1gf4vQlgdaizpFBCsivNt/vbfvBXUk7ClI
eDq4iJHBT616cpOLG1UaLOutv32nw4jIzMb1fJnoZEOPLoTIyRPh0Bt3F19YtWB6s3wxy4t4je01
Dfr4uRZ8Pm9kXL9sxFOQy0Yvr8ltgBR9Y99f4rVu7rrqCeQWxy/G4pBdvY6JK8cudNPnyxq0SE1Q
WwJxTOVPnqjOprJErtsw4XjzxNYfom2DXTtOQhDAwW3LFrWwZy7R/xco+2jxnRN0SSxt+mFz5QsE
1gyphZXjnljkpScwbU4mwj8h2bdhuDm1vtzZum9i3t3Qkc0/1VnUv+VD2HtNRfY7iJZh/iDX3e30
NH+UvdR/MluZyPF8zqLqrZYx3uRVYfNTa9Kdng/tf2x2VWmw5PY4W743VnvN7Vsa7qqs7ckjA/VI
6kYfsaxfElR9uuOwlckjMdWOp1eFwUd+x+1ucpfAY8kKSuHS6Ibg2SU7fqQ75fkcKSSeM4Xb0e8Z
tntD+XJBAX+QhLPW9/B93oLbiW1gJe9cPbPCH/Qd6hg0NP/FINJ/Gk2Lt6whQ5G8FanLU2o3D4MC
khG4kXKdc2kOxPd+YUpwN42BDHTWDtrHvoSwfeFORiNBUEIXXBxlPL9AjskT/VNNgOgZ8Mk7+Fcb
pON1HZkQyBgEswJG7jrOzlBzJw/YAHmEbhBZNHTJMihk6hWCv0ipF9LMBodFG/ABbHxdhvjicKpo
W4bYcKhYG1CzoXOioAOHQ3GRP/rkHvGDPhJZ/SwtiU/YbQfywZo+8M1JUAokwKz377RHf6ureTDI
Y6tDdVtsXwnPe123L1mIMoHu9FwT7V++FVEv2NEQsLSD9/KErR62ZMJG/AP7UrhxyakCXqQFyYGj
UxfID7h9Q4Fmw9mz9fKEml1+MXjhN2QAJmaMuPFoYjtXT6keJsGzDrWZGt2N4kP6A708hM6y3M42
jzeLxG4gxVPb4GmuDtoZ76KSXWCWET/lVlYVSaD/Yy09CLaYaqwKP92YkpTqPmjVtgYFAekPV9fz
lir07zo9WT/m1co0T9UAdd8KDuIrAlH9gqws6M7rVDwj6m/RsQJGBQuCg1X5dJ26Vc111EmxOjqW
GPwhE7BJjDmj5Mq/ws0LDyR8xKovk1zQI8q/IwofOudd1T6Zq1sloHpJTrPyk3LObF9dvwLbsRtq
bRbzu+E30BFVcuZcg38r2QqTEhw4UP+eZt6L1kEEeZZIQOH/UVGMXVJEhnlXTEU8FYABbupyrMFo
aiDGdpiXpzQNzdfGGNLXn3gNqBNLIg6TzI1TYR0Bi/ORUy1DBlWSBe3t/YIWzSbgKumZR2DapJ6r
r+ZGBwbSKsRQjJ4pBk+nqfI1XCluIEAASwmkSdIU8Hbb4WrdG4ow/IaM8gpFuEGhK4OLiXXfyStX
G3CaYDEUE7Y62YIchsJ7janGdCQqKtULlEyGuCkiWn8HiHUSuCxWB0hO8Sanidnph81SRcPE4OqN
bu9iG73zNvVEtzSCy8LrbtvbtryoGPQ3hryiAUwMj1lKYtEHUUmuAkxLQxnL9yh1cx0eGmaIshwJ
Oe/mkYeLTo0/ahZ6ODkhWcpaNW15ZMs7niIwI4WK9vYo/dZMr6RaXHvHgrMACNkvnoJqvBbbW/F4
XXo3VtFCbQ8ImCDcis9lMWFeEn1bOnsCaflL03ZLMdZGJ0xBRCrbPzx4K51qR5DjKhU72x9np887
qDdN9B7TR7UEzr5cQVNHwNDr+0sFi61Vc/NVQOZvI7iLkGIjg/y4PSEORoQ2K1Fl9FNhiyodpWO2
JXZo54C3KI43W0+QKdca7LOqzkR/IxV2GSs7iPZP3kkZR1YZYZ3gTVJtAvI8DkBJJNmC/OAkf37z
PTsrjnTiv1rNgX6G4T3QMO1MLj+Irg+3vE9c/qo6TN3zkSDLqc/HT6l8W9HI62K5hFy66dzYR8Fu
BUIqrRDqzsYAoTiGyZpHrZr53YkgS3w58eIL7RzTB/TMkSkzk5YwsY6PhPeao8+PzcT9+aKoOiyx
sl4v6xlnUHiq/pOCkHD7G4yITTItPWLeAueTqDq6ZqHlmRBXhhdN+LfYOVVXkfHA0URYPUncXSRd
7XNaZ0wCoCHjCmQjvmWIMeMG20jYMxntJS0x2725pRC90ZCys1pLWo2jFVVWTkYJ7mTEvyd2v7Z7
764ZQSR1jp1oe5kJXTLHRrQMipqrvpM0pQWkN/H5RecEnVKaWzyEC+nzBvc9pYaipW03wD4t1hBy
e15LgVnP1TZq8a3SatCQHQAjbuBVSQnRJiVoQdfYn48t3T6j/csJ6OoVVscyGHled/yMWw2fVa1y
tWINwOHv5aTVea6+NryXLYzgSyUTXsvQdjJPO9DpBIC+iEiahqlIZ8lDDOdSK/UN4FpadJ/96nBU
fuZpkEjZoxlPjFXSOXGhQHrF2km9i7G07kkuJjodvt8QK3OS9kEAv2sChUpyuaHvoiqgclLNGGGz
4ancaI1ZqLCDoVAe3nctiI30ypDmp0Y7eXA6dGq4h044lvAy3jkMP4OpixE8yg9ahS0vNkSEgYbP
Gb0tticxo9nHFpea4upYP4FR+SQgiNxrksth9cGm6Iu59jUY9sjqkpAisfWoJW8J392dQM651RVA
zgUlLNkeD3tmZ9wy8IXgxcw74jQR3Ako++oNJyua5HjztBgVVgzeObhjosdeZrXhQSZTV22xG6TO
A4AobLuGiv1RzrOKMSnvOA0Zh2bL/gO78mtDnfE5yDwMV1NhYcKAA8l9yNAwnEWRsJi17c69wS7C
g89rXqRtPcxC8vuK2iSvuFrtPyr2FFgNOsrE7OvjYFSm9KYXkC6k+AkQSc1UdmFXUCO8+zzdc3za
vzj5/ZVKHqkoX0Y9ZIWdQW+kCx9gejRKL1GWKrzVQNLo9DXCyv6pRiIttxJpNVreAfiwwM4CuOBo
Mu4xrFPTkcYEBnflTrUG7VdL2K93A4OilOVTAdBw/nh8jsPDLZjBTt6tlH2sNG+oP71kqaNV4N/e
tmgV6gBmnioRbngi6ZXnhm9iL2S1CLKIDHZjDpPyeEefa8xm/XJYm34rxiw2DdoTj3dln+Xvp+fQ
WHZhzs4XxWYyol91p4F5HEeb2AIFBJGB+maYW/x7E9ceJqnggR88Cf5aTZhYoB/Hl37eoU1LbYaB
xY0GYm3wDREPEQ307udJ1ycfAeHX/3fOwRbmf0w6zl+fT/ZmFVp+KPEptcGG8KGnUI0v7PV0vrN3
W62r9Uy21ZVeVY6f284gDqQES2yaNjBC0dLTwesDT0dK4rLnS6bD2J+Vwgjtl7C84fffq9zQ52TZ
M1Renw976p27YnIj4BQ2kC6Y74fOIz2ixvQlCYFtudssaVU/8wurqF3exUk74Kk1Lgkkwp3UCBUQ
6ulSWYoZdlWFlKD++YTpGpxDqqAZV70PHUmD+VIzCngl3wyfjF/6NAFNvJA5m4rtiXg9VTIjH6Pk
glgPX4nZkSWdngEi4uAOkAnfHqvLqCjYyps6sAA0kx5eLtUrYiQ6LOJPfO7hWXtyYP53rKRhQrDJ
D8AcuiwPKUhxsGJlVc4jDAY0Ylgb+y0jnFk7RevlQkjU8Y56dLbl1SxGFZvLjOFl/06K4pGY3Oqd
24CF9prYjqQyVHGE5nQVNm3bMpIbYUobM8W0fERIYG31BHEt5Tw1l/Rw+tIuF3maVKCHwzz3C4r+
eTInvLae2QmnYEWNjORpi88Me2m+91kuwlBrNXvXsr7FxzFYcpEgqgQPpG82CrKQW5lW6iGOVDex
v5BE4zQy/J9DnpTGroKbPc5VVKisk6qwpVaVWkqr0U2UP97LDPkv/RDPsQQn0498l0a3PM76K/V0
IfrctmKCtVdBiDMoxqI5qkQJXRLj5l3wyPPVybomuXY3/nSK8dWj7wj1FX2uao0HpsYILFE5AdA7
5luoZriHZRPXIoDfnLSPBUNEm/BYTxyRWgT6QdjZlwgI9PIhurjTPZBjncWEc0xCMuVtBpeimatY
n+Yjl+462nmy+NSW+6zUlpCKZm8RhGXXp1zOs8MOckdZbrKQgIvm+b+KNpGYL5ymQnBt3Pf+xzr6
hf8L+l2GlbOGfIXs5SzHCTv8g/i6wgj71MrxDh9m2umz+uWoja2CisePiPQcAIvD0O8THPeqXkYg
vaGX0abMqjhZMRx6ypfS5AEThDT2TKfdBe91Rm80aBbMkDHSqFaj90cIYahDIraw69NB9yStHl/G
8rYLkdcWuPjlZ7GCznTJ5KpiEXVSUfVltUkYU3iDVpytxDJbcQ3awYJQMLSSnHdobi//jAx/YeV7
DFHw7BU5J8mMGJegpm7ehTlkDNnlSNLjxyomwFw+wQ2tRgLOcjys2t5Ep1UYMn0mCF/N6igOr6JC
P4eLSublt74toeCEpDl/T5PjIR/054CBiYH/4ICTzBW5bgZyGcKed/Ac8qHqs5edaMz9eHH2zZrE
oZTduitSslMvnZEKweY5QxQgnoTqGn6DywiydnGTPxIquLkMeUF0d4i1h8LFtpHrm8sS8TAcMq/5
6VQBIwJYuSrMGXtfRNe8Gc+wj97zsNMUYA1sqWLvDEK0wH7rxwhgaQScwzs+vCpIjb9YTZJ+Ava9
/2ngySXk3xWvlemdz3DxspeKuFBuAijh217mdiksgARr5+BRr5sOOpaQ5jtP+Ots2TydUBpTaNOm
nDcXLZdo0N3bv7noWZ/Ko4BqQCFi5KQgOesM11UKHh0SWe82ngwlcvmN1YRKgHbJKHNgvMDDjIsF
MleOWcYxodnynWxDpeomhyhYSqcmC1s4oD6M3ekJ63xKZ0taQOxywJmqeIUZ5CNmPyr/YdfbRBY7
48NBJU+Ex4ZciCDO/RUTH18+QHzGZitHo2ZA00xNhJDS7azr/LcM2zz5mVx7rTAD7EjZTjixh//X
6SkGEN+r5JwIyYDyuCak/1bkHBYpfmu5Ls0GZnAMI2i4LVUZM0nLg0fWEUPBscIV6BZD6+mARqlD
419uLQF3FNfw4WZ/3eVFS5JiABPURNlroSfxoF6KOjmbCo2RfjQmkW3kxPS4rNTKu/vH7WVs7J2W
p8KHFHlPMnV6x5AoIwgSi8QWoAmQo0+Gva5nnHon+fC9sR78fh5G+lbt1H30g0ka3oDz9YFjrBvT
GzRr4JZh+2/9wIQeAmC+bZXGp5Np91ox5IlvtVV/66qchwsoCKRTk+mzp4rlJvb1B/NI3fzGcSDN
ihqgRfRQpd++idR72HKK+Oa1m2foNRUWm3YIX5174pSfeOr1I8sDGmH0+/c0WH/mvn5Gchy7Qv1P
SujZZ2BpYTXWuJCp0P5856WZl+lv6zYltB2F+N969pKYigDrHdRjsV+TrDPaeCiThOZE2qn6QWsg
XNokaY0UNhEcUttPfR1Ke/sKnIstwgW1i2Sxa5DdQ8eiWubABZtWYdRPytrXfLbDU+/jfTw/cN1+
+Qpx0mLJFULDLxa9yzSEu1kdFLdjuLzLCDp7Z902dHGp203Zuuh1AvMkF0QMTSvXDSV2MKc+3pUK
DsbLbhoTK+3WeCpkG9Z3IlJ3wfrbtf5bUrp6i9G1Lfd9BFW09J89ft8ee5eCRy/NqZvDfgp323ew
UnvQuAUOJnyzh3wwjlAD25m2Drp/rxChekoomazjUY/J3BZwnKbEMMBR3NdtVA+56p6KyY2glb4E
ag2aqRN5sjyrg3p2vamz7GyH3Pdb/NCFigJ5AI9aMAQAb0m+ofeYR01GW3SCcELA1A/2Tfgkbwgj
rJ0xUaRMy9Fopyb729yyNShyuWklH/X9tOyde4O5mu3HsQ7xwV+GnS68QvTI/XovGX6UQXHp1iko
eMLygRq1I8dL44FA5Q/2ubn8SdnXrItNmnlOHCKRDSE1CXb7b55jEVxa2KGUYVf6WNoI4oYOROoJ
5W4lJgkJ4v1TfvXMkEWqcJewoVKFpI7ZyMPC801FA56PZ0b8DQh4nqXKb+7Ih0Q3MBy6/QS9aUFP
eguSa3UvJhIxOJdJwpPNLhZMoEg4jPtTfrCD/69QHQhLwl2RBw4gAJz3VL04x/Z4n2ZZlDjauMgK
JjqykHZONhAxoMy5YKitJHwf6xbD/WTjDKzbsugV+DAHiHMcryLb+cxM/o4nPKWDWKePNUtTDpYc
Q0z2Fskglptpi9dpYbzH4O3mkNvVQUHm9CLlahKjGw7XE5vobPuPyVUqmAEu8ukPsMoYQbPyrgvV
xegRsVE5qDdxt5tt1RDCxPsNzFP0rH8qHeVKZDAxtadGgbkDrENGNt+Fw0Pfg6VnA/Slmm4TjFo8
PbOT6t1UsUISr2jNWe1z1KrhUSyXWz1aB/D/hBRdZR86szAuYVNZwt01cywWv95sRPiBoQsrlnOf
ZHnQ4JenKVkiYud8QMDphT40Iq8Na8maaU5qgEfiT9ZPMhgTIG6PH3MR8bmoyDh0Bjrtsl2Cixg8
3bqRRsvrhav/gJSI9SdLKzfbMWDpZ6L0PtqsN5EhKBsZqFNuyf+W2VPaJmUbdAInAx3LsBEwusfI
Dd1mqIaIemc8HFF36Yw+K5LXc6PQ+XtEzjqd/+F90XbArAyvSAxPry39h9EC8Psf7OPwXt26iqfV
JI/1bdQqygagyNeg59kXdBVHv6xi6TPpsb2wE39lLOPrkd5BQgm9Kkflik6RNQnBxgiMiSxcCmV1
2KS+7rorNaPHZaHqk15lWLTgVi8ANurXTTOZ8yP6NWOmQQSN/lKzKi4qiPkvKhOxN6a2eT/IoKlP
JQVNQvH1EEgCmLwrNQ6ze5jQp89NSCG97GFMS1n1nZdIkIDhV9bnngwrPLaKgF0WZQO8Z6pkVzKq
zvLT8M0+WShJcIGK4dlScgAhyBHMnvIBsEkjN3dXNix9VIT2xHOThog5ySUX3ulyaSRqC5Un/Pq6
JXW/qFbEFUGf5aEd2VlCTI4wsjWJdSjn1qkv61fNLvt26NOA8NnXI58QwqTVl5s+7fc+i0lOdj7T
GzR//Dik0ihopQeIjGu+RFoHgpphG61sptHZWFnuGQpk0GSbaUn7BdaicFXE8Sk06sJRVr5Aemq0
gB7Sm7NM8zFvKk3nzq6ZjuDb1GIfJHiT/Uj+EZOMNWYVqOFQBsNqUVR13nVe3LhlOOsiybrF9ZGV
M3+ZtysC4LixXgDS/aBR6Fd8prsWKIY3EEGKr85U/wwuZgj5iQA7wrDpw6+uvgHjzD17UUkS4Mul
REUAdmKYRfmKJR5RaiUwNT0PGh4Uez8x7+exyYPhj6Tx9mWdvFmTi0oSM97inoaAyw3CnZ4sPYGz
NOwgZq4zqnB20j+VP0LySzHtGpGwAy+/1oDteS7sLmR1NfYI1Rtp7rjWyZDC2JdJfD75DSMRJ71Z
5MIZIHy2ELQeHZQfoxBCsHbUg8TMn+NWaDw5tnWff+QO2K4+Q+kmVLrld2MUy0Rb5dSu4vNgnLPq
FXxRSKFJ9r1N+46sxIgId3Ej4KjueyHk3FPjpjKGFFp646OygfGpsq6ArDuzcTYkLm5JCBe8gpmz
p0cZoosTjaO5JaYV0JLLRVbhOeR1bQSjSHntUv3wJ6rFg10TNWnDrUD1fKRMFsDmJryrNzu2zbLE
zTFWD7VxVW5xUWZ73Hfx//pkq6ZtIFVUXGg0Y8rE0O+PKMDllcKMDNO8bkG2d4pwbQhKLZ7QvPD/
yCEmxuclj0yqpWSonY1KWq3ktahlqxdedeRofBJx1MoXqeXmwB+zLiqoq2dik+nraK+FIuhAlwPj
SyRgt6pr/toIehhh7nSAKSPi4bIw05QJ+7MXo0r8v6jemsV+PwmW8Id7ft6wKf1ANZVgy8AIt4V3
mUZRfcGoX4f7DXfBSBlDzf1I+yM5JPmT30EWs9XPL4n7N0ISpPFj4BFktdEp88qBh+m0lsZVJAe5
FrPJAkB+lBw3MOw1dh7YzFDJ00dcZbbRtmozZBlFAAWMdhp9l3g2ThY1tIGa99mh0xEsXXIz0wRK
IspjVlThAmBClelwi66/JiA5377xCx2uaBJJKECpyIcrQSKt/ClCLuU0jmfgUB8Jsx4U/cIupSe2
bYBIOfCNSELESWgnRaq13kFJX43s/v9qYkuG0HqdszqDfv0ngz8WA+hT8ja8SCbZ1pyWB+EAXnlp
VRZVs9n8wEKZ07RI1S7h4X/RZS2712lTnRcGHM08N+1X3WfsSYslj1RhYmAYa7D+4huYyyGQjg08
liPYNWE46y+mfdYNXgYuJi66PnZDl9Kd/i4kTLXxYFBPXZx5MTapoSB+E5EbyIDDGy839Gcahk4u
MZLOqCDH5qKU772+3ew6miR3qJKlAh3S2h30A5CEUE0bMhwTbg6vX+ZueGJ4ZV8pFAwt3JkFUeoR
zlKVQ/zTOtQA5uUKjBeTMUlCJrR/zDNw4moqIWFUQ6eStZkXxB5TM/w0ZDq02kgAnBdUdR1HPGBK
1bRSSIn/iJC3lEdDQe/UG0FyA1reezKaeArHupgR6N4d84rYoOnmKgkSFD8wcP84XtHnsgaTGv5H
mkkJELwaW50Ifc3o0Xs46NLOu+xcJB9OhjOUBwKoAXWwYbRjdyeQOloe+OKjjgfGbEMc2adBeAV8
e311GWDqCMC7s/DbuOQ61K8Ad4HBK5hbSwl6G8x5Ee0yz5g4Evua+jJYqV4yIRph80Molx31K095
D5H4yfdaTb3cUK/m2UXiLpQ3qyVRXW5gGExx57B1SWaZ2mcM2sIcZZ3pv7NfmQgSRb591OKmYgkm
7zaJC1XJCrrBfljPWMvZqsM1s8mcA2ODbaDnK8lvUnZblV1m/jnG0R0qwBa9Tb3qdlouxekN2WMB
Yg7D46C1xqEF0lTXpuHjmIpMtt5fB8RPrc5SputlSqUqSE6cOz0A2S1yR+krI+gf7XeQhlHnYRd3
+3V3CGW5qMkymRJ2ZkSy7vUOHtiPNzHKZOGCOfAiJOdWOlG91fWTiUS//BqqQJGuoorYTlDMncZS
GZAiS+gb7lLEzz190vrP2PlbLm63SB9x6G8CLuGQUgs18EFJ1s1RBhm72hsnm+S2qzeb7TURf6G9
+Bu4bSPeV0l7dFNks2p0hbyX9hi2v55AdENBmjxV+M/wtD/L6/en+XzKGgP5RZRs/d/F/1GgOsED
CBbT++GbkjRq/5ZcImpLOOcsbw6MjUGVzm0uHL/OJbcC4pBUb5oQKNoPoNTwA9fO8pzxvw0WsVL3
ka/XXuPmMnKwQVAfE2TvJJU9rdJHwpBLMastD/HLdP2MATFW3+9zN4B0N75G5FpNP/sfyzdeAreE
8MIkxaNou6Je9NdMReseeneQrPaefRgyFk2LuIeAlJpAf/pNG5I+KYeqTnzxx0JB9yB0e/1vpJI9
y+sQsW2OPRfTOoCKEw0DfbngR3RBhbe4ICmrML4hBsOiNoqZrr399umgIlEGYT3KXl6KxquGv6LQ
rZTVggj4ySJ65JNF5K7wjNxqNgPHMBc6Dljy8U4OC76jMQNmPeNEVQHZ+7jja3NEjCqSHubz+W9P
JM+ecOPFu9v6AHqNdI3gNN/3EN4wXKTmH74OkpZsdIlxyFFYPFJN1EFPCzOCzXeMsIYAaLJ2Ku0s
qka2L9fA3iIAKoWBtQql+d/zI7z6mflxd7IsTCZUFKeHC9Pl3kwurhJ1ViCNxtMxJFeuTxXje3C0
E2c9E6UqgS1MbORkmlXYsxrBY+sDlR+33YHI2fYaifBLvcbCNgihinCnMB/u0xG3KB5rfxV9ZvXt
REsfD9ve2QKtMGd0XwFEFNF3I7fW60suVlkgKU81Y5Pv7OHx53FUp7yhc984VANOs+LR1XKBB5PS
CFNqWWgTCPo6XlfG2bq3vACBwfevH5hwDxyDJGjxzwADfVqt73AdMY5X9wbD2SdK7Vko6Htsk1Wo
ja04Tx1htytCbP81LnQ7HU34j4RPpkU7beXx5zJ0AFQh2fKa541n9MrOlKQefVtlFmHznQ9HmZo4
/25o/evD5qVBvMJ42eCq4CGEIPzgQdCw9z2DkCu2ZPv4KimuSvedIceeTnYA3uTlvJwfbZOJSE4F
3yQXSqpLH0NZaeYD/DMBYrzePji/NJSvEZdpu7uRBE3t2jfow2DuWYukcXNPyuKS2ByPzuUvRCAk
Lq3f2fbazaiYcqYvmA2emguWY0eataX/C3ei8jOeOKGRgbAx4lEWhpe5yPWQwbU0awIVnoK6NRiU
BGYxqSGRLdrnZajRg5cpJ8tBrLqjdmcwRpKhTQcng/KuP3T3IZi3UrkJeBJZXeek+VQLe9Qd5se0
PkB0q5NtYF5oWGA5qts69xLAv6qFh9t1rnKhwix1A2C9030inRVr8Le0PP840Q5AwC7+3BvB59u2
k71ECnKxeT1WnMskJPY3ua/Ckx5lGFbfnlZPdiU5GSdIpf7dRC2kxIEIKYf9myHjn9077PVNQCLt
hhkukjTIdLFDNkjv34CSAENLmcc2cCKlE/gvesE7jUvFN29akOHoFR8SYaKjCgIhU8pAP4eBG5LV
GsuOZeI9UVbLk+Z3BVC5nmR41Yqg+p9jOLnpuwdbs+slu3QJ7EQkOSZFYHmv/bUnuBVvUuRF6SwP
a1ELdixFPSmErihPPLUw6yrj4LZYqJduFIMKvDkXkHe2ov6IllySFuh9WAFlo6nZHfTExk9TOO0/
Fq+KKbl0U0rLZSeqJTvqhnPtmnYiIqEz0Bc3RqSFP4O1K0+m+UHEEHR5/2vBvx/NQzIpRu/O6VxD
q0VstynOCojSHgLdmm8sZGAedMjF16vE2jah90Me/1iAUWNL6sZ78MCoFc+JUav3i0iRzZvkgli8
YrUrhWeUvvhx+ROpuzK5IJogeXM3IneKRQ+Q73W0bcFvsUjHO4pQ/3SZMwoAJqlKaaIVFIOC8CXj
L0EYCJU9FGk01FEwf5nBSCcVWEGbpqID0/VKbk+b96fRPIGK7rcxW31MjjWFOEaxqR00JX6b4kSe
xywcRnZCAUALvJlG2fpx+VcxqVzTkYZSN8ZmMllmiPD3iY8Mmz16uirc/yhX1HKA9v+3gOxrJ47U
MGEgunDWGLzXf+l0yAncahVf5cNMKKFQ50tTb8cDFR4aPY5hlfpupjOF0Pn9uSU3KFX6j4b1/8Yi
3moAK93hfJMg8jUq8tfoANJlFABg9SGt52nYFUYZf7htmoTIANam2SBKNnR21yCQCN9fnkVdlzv6
cugJtOgb/zxrLp3DTRSpxtloQ8pdwAA+1z11s2c23Saj1sle7iB6GTXuRgd44djz91QpHzZTQ7++
5zOUDc47fF3nLKfMfWCuj9Ok/XRiKn367g5OswCBU/9RAxCS/chkbpctIU2Y8w+tY715NgHB8++L
0D0irsdUwiLECYAtecy9LdVwpKRt42BjLXvIkjhQPUNp73bRANuNTsFg8Czmrz171kDzIvLNEFnQ
zz0qYZePHP4aGCGzRxdoF8YZEBC4u93zoXL5FLKysUJJRp2exz3Lz2GmMU80Uw4MHyIlRUG5ZAWT
3GYr3SC+jOjtBboZiYWE/CIBci16ijTnN9R1UhSoCzSe9VXSC5wmZ06ySUZ9oIlQwGIirh4QIhxk
Q3m+/iK1pstzI8JtAPJQS1j0qgJkSBUBglG0yBElrXBM1WwuOeRATqz419nhSkOM/pqDbl1IPcOf
cdZUd7oqtN4b9ZgAJvvxMcR03cWaY1lJjQZQw18XNObbm+ei4oJYvLv3QhXJvP41wryf2p8doeVf
TOfBLq+6vLEl2XIoQLyGnWDyImMuZnVIyCmZYQiKj+ggLnlIZXgCEnSXY9wG9Z/ou0ShRUECmvbq
01xIeAmS4cuSicdvx5UDzbJZdauIDc+GXfO9UsaXWvNGs0vkBuf6YBbdkByoaDzpIe2+rzmbtFS/
9ux0Rop3ifn+0zCF+ZQHJIXfGr5sxxAJwj6UzgXx2Rlh1BMYTkNkscc6z8afJyHKkd5fgPGS+WOE
Thvqob67WCslrLozk3XwIm8slc298YgieVeLv26zJG4YYKvcAV3KCXNnax9qrrPOKJsb9/3vzEtT
Vu1qMPGmgyjfVXpCu6ubI4LhLOzDcqK29FdE1HKjOqhW63c5/c8MlORMJyoEp9gr/fNwhg+kGooB
sqsFSgJAVIFmQD2ck5D7trF2oFCSQ1ikIo5Uh1rIs8AUpHVoCI5plHiUkmbreq4HF8tma5SG7VjF
/5bN9h5Q8yNs5mcbqqdQEieUZzREhtlK1gM5JYMn65sedUaNIOYw4fIIIQbpis2+Vpac8TdEUPru
fYJt6St7ZX4mQeaQbHLaiV/QhkYMCT6IJidLXU+wg/7xge63T2xk7iTL0eSJpxWLfs/e+vFiYGth
BFMecwaKpI8OrvJSIIIzuq9k03v1+tjpBJKccihClkdFJwfVXR12fcQiyGZhPH+UCJN5IJU5KS05
QjmD11zoKOmcO+XP381gI7J3HPGZZ7tERzyxvxY09if9VCzJJpoxuNTY9WSM/BrpqtJTt92T0Aov
9rL/W3sUt+b/2kqTIP4KN6IB1CLKP6aJY+YH1YvGjdx7f5drIPApW/qNnS8CWTA4LdlQPn5ONJsG
C/zbNn8vsHaC+K7aNS0ivqqRstFzOqea7dA5N5Z5XNIuUXSgUs1IjpbR80j52lhHfJcRaddDyhTJ
XLuWMTxX7KuPMpBTO3TBTOodaeCqKf3kU88VNPx3Q5LPnmKi+x+6kiCduqIVmJz8JoNJB+aP2LDV
1z7U8fcUXIEJoyts3AIEMZvXUa2eQxsAiYNcyznmz0z38yFVO7lTd5+ggsMlMIFDvwoCM/dhdgU3
SmlER42EdcjqDe1B0wuyJCSZhiJvxafDDNCbo8rZJ8shFvxswFpT0echH3YgMJ3A9SIwFMLpSw+i
qux2qkt32do9TQP0eSF4tblN3JKsTcS9Lpzzsuk5TjM+RgeZjAX613d23PBfqbSNucQbwuRbc5O5
O7l4kfh2JENsh+QCD7bLKpKaPoAmukMKTpR4ScV/Ok00RcDi1W6exG7kn1e/1y8owyhvyhp8aoQk
dBM2CBZVQxA93/MN1CNthYdlqqHtXNAXSdYRoCet5EDZXG+hOBOaz376CsIc+T5yL7yQpNSfhHV9
EPB8mgcH7RUqC+rvEVi3Tm91joNl2mD4PyC967CpqaWLApMNNrrThs7xDH5lDqqE+YsucvKb3Y51
g64pF6AW0McLmCEWCzEX0yajA3e97HMP77kewbsdUa5z6ElBTeA4HD0gI3mnPbKINg7VYuUKvpte
UzrsIC47jMSYUN3KkRlIZszvAyQEHeemW/MsW6NjHVq+J6Y0/YIc3dMUujgGFsMxALN0NJfMO/S9
qHNfFLIfVVI3TWoSVCJI7R5j7ISz9/HLYiZIbpQabxLvAnHbg8NPWVS7QElA+Tjm/UFqv3qyrOaN
fEhojJO1jNp4FqAFtnbS57DPg9bTgWy9x4LcwM2uUwkDLzVyOutfrOsmvS9UD/1v9zedv+KywA5u
PYEXCEvo+XirSsDC0nD2sv+f85NeFuz5OrN2U4vmYL8QXoDZAVIJUW9+AIYBa81rfMfzA9wYb8Y8
scZY1tLDoYq64fejt8k8rmXIMRIUCEZpmSVoVOb8SgytgDcInQ48ygpvEkiuOz6xCMid+vx82FVC
LecJg43eOABHDHB1E9zr7dxDYf32Ez3y+PqD5IYcP+VXyxakEglqoozLXJ5oJYKXkfLmfGnHCR5C
R47DNPd/Vl//ht2MbDddum8CNWLqe5tXN4J+jchYRA48f67fe+CNwfVWmHrz1Bh7B6uWzRow8JGo
sfE/afizvFAKAMpaR0OMndtWZ/jOaevIfkUyj3dE7+0UNkV8wuFSUZIOC6hsU0wkCdubll1keBgg
54p/ddZwMGfNOoz7pxhq36jIH2F+Bxutxtnpi79IhQfMwws/7nSMlnMlgZUPv5rmZYw8vbPUMNmK
mLAynF0AGojTOAr2p5KoOGtGcBfGPayV0MzwjYt3NDnZziDJJ5ACxsXsLomg4m+wKVwmCtKZ7xYL
zj18ucq074gxPnifLEJbKD1BDioEB47xwo3u00R2HY9oa1euEq+YmlEaGVHYNX0dSu8h5Y2j+Scl
2sBp3mIXp/HB0T7HV5nR5kmDgfbtS5f2MGwmX3v3mwkKO/WKqa6Ww+xyMyRLMG3hinPiJt79Vs5I
jvTuCV25SMUt0VCPcxZq2fHdNRySBZ94b6yjuPDfwc31xSBE2D2woayvXWBMe3nJAuZnlKdr+YCe
SPXW3txA2D3GLFTI+lDwobp3bSCcA3Ay1VvpxoNbhzkZbMFtVF66VmYf2K6YNNwV/hQ6r+J6NKux
fJaK1EcAv34WXYvB1/V69B/D8c8ILj59AedG+lT8ihvLNVvkNVtey+2ZJxm4vjDkB++KmGMXjtcM
GZMBPQSkg0dJkAB1vWHvlDpbWEyiitoyE4dbmoXTXivecXw020CLTFAPfrkdi92xoZO0w1+G8BuV
6lbNZEyXaEYmT9fUV+ghV/zJIVDt4gph7xHdwfHjew/xKpea4PEwUFKou2bHGHZ23plMYUljuIfu
spN1EKmbBoWskXozWFaq6w+e0mUEs8N9ueLD5yvOWo4Qq7Guo1vmMU/v3vyFFAT3vYGzcLnTGkgi
lNXZasFmkVQHs/NAaH+k//kfWPi8VceZHgObfz4iuYVNUzXMpu4F4wDdy9kK8Z59AWc/kgRoBa4z
adw6d2J+waZ6DAtYt6R9dIhpMkVl0yE+FZP8efxwbdgEZy/jkLepfJvmtM3N/JAC57IlVbMJhnEJ
yXGY38/LvjgOuk58F2LV1WRjZw+rVO+V+U31Vf/G7cqSKC6llhDWmXRPp+nnxtnsnbNPs+rauM6u
pX7oV2/XmWCSWPBIVNaBgDN6kt8H5xxCz7lG0QOJXqTa1klO6t62S3rTSPZfRNGcRYybNCw9hRew
N9KTSNWSplM3GZAxKjv+TqstyVHWthPdgfX2fkxhZ7o/tFuYmEd9ZLydXEc2D0aP6Nf61UNmhByY
rrS95tCCjG2JJ5ZzzIIV94Mn1lAfsO2oP45P+qvYDiUAb9QvcLQP81IZZNI4olo2G7kwJjVyv483
YBAY1ghwzy/2uug9xD1GhkE0uKFIHXb3qbLBSzuNdzYbJSB1hr3yY7Rfx7/osugUE0G+LzhSglZw
lwkZVFob8JGFv4vOdx1Idyq0gqroFldf2vOUjaHOj4knx9/zjWDxTtU64A7ubWbeMndxmOEPHjLs
Ns1D5MXdI5qN6jU10DSRY8RLTmK7YeUO7p15GjMIL95Tdfl76tDfOPiZKLnG17ddq2rPjs1Ue8RR
VBpFY9Gi7Q/9+5j8j+Bqrgh5t7ThpuOXWHsFoOYehY20WamqB93VO6YUoORu+YIIlsr4eWOuz4yN
KSjs+RLepDXZf5df1+JmgRA66f2POKPVFXF1DKWuq7DpC9wwgM3A94KJmop/vRYBS08jAeaPUaGc
U/hNvahtSuyYZfQZsH4vEcTYVLAVD4hSH1/JW3W9QgY+ufkxURtnhtCfusw87N7kcbHEUx9wxuHA
lqiyM6dqRMkP/aO3CMpHLFRtDmDPT8RCm7NflKarqsU4JcD2ZcBz5iTYbEjeifaYMmZnqVct0LAy
ozGkSDLY8xeXwZJ8vEDB5VRYJCbKV1iNZJ/ZvaqVFyAbXCZI/Ag0QhpVmKPEXWjVpw22pWoqut5C
AuDubuw+qmrpmR3hN9GPqf5g2W9XxRgtaVkwS8PmdmA6kJ4tNxSNMWAQv+cMWg1U7ByXxQ8grX30
a1hTyJW5HuyZqCIJ6AdNFYIm9TJHR9TCtCWX4HD6V8xKn3BJ0SICX4Ab1iC68c70msUsTDya4Gdz
mYhS0qOatjaDEoKnpF+wvjTHtMmx7pefVF9qgSBpdz3/CFsNNRudtR4VfGxwlzZMMVSAEp5ZDN3F
9drlFuwVQqcLuWLVyB2ZhHHcmnzWLgCHgWBSVzHkTHg4usyoM7t2JzUlggBHwNkDYT3EIe23rgvF
PkjH0Z21pv9+p8Pyi4QL/Q0S3h3SL6SySzC6hoiLihEx/3/qGIe2PIUG8JU7u1CcekiJUy9hzCJ8
vqZPS246jRANR+oM8bBuRLHz4XceZdaHyppJ+ii2z0jDfeXzTjt36VCHR9i98iGP5rFfn+ljO63n
3Tzt+LO7yqrs9ObUU35jmnKpwTaecxeGgglIwI6Qu89Xhs89r5jLZyRu4yhOr4HPgSJFFcrGQPJy
y+c8Kt7/ildKN3FzZMVhBSyd2Ko28Ex1rlLPcz3pongarFcO1kFnT/UWJD0rbWJnOsaVW31TVaXz
7bLVws1maN3YH9HOVfRqYij7JKzUXrjJK1UpSKcmoeB07BmNWcqb0JeryzSUb+/nb4KWBZHE19xc
qsTkU0+kPSmBbr4KMX0M/JwFO5leQIoWhMKX2oH5UBIBIlCgnqhd1ofXO/9AjS0bynE/Ad8l086C
dTU3yjIeCizT5oXWs+/+VDgHpxDx0e7W4zuWCGtJjTn//rDfWYtW/WcHZ5aErWW6khxJjvg/kj8w
E67oSOP4e4Fd/DO3rWDQfdJcRVlzH/gHlBfPnFZzNeilR798BLEAKAU499nRVVeA3+RBshWVRaiu
uWxheLIHqkjCvekSOwjETQNXjAs93Zms94bGD9hLgteqvhUYft4NY6Fid41DkyQvAXNDmxI6gX+N
Es6eGBSa7BJuCnxFYUnjbj/4VI/KPdfATa1hJlaw3y1Kv914cTjtxkPQ+R3iynXECd8lHWUGuWRx
rRoVBarwomxsmTBVPhyC6XzPlJ/fg5hsrp0R6viUSi+IPLWuR9pr7n8tmI2xgT5xpZFga9w+UQKB
Q1XlO/MgR2hiQZ9yX9ixnEF0rEldAlu2svlewC8syCR9GIJ8kytfyBLeznqF9J/qeff43dVP3ML9
fInRWEl39bjNBuI9u7IktW4eA10qSGLznv6md2oFLnGjAzRuVitBd6D1nqoPbFrverJG99MdDrmt
cLr5+zD0+mZFm1YPMaAUQGCWO7IZUw+E50phbP0IGOY/9A49Lj/1wHmXdLeCvTq6WSNKDHTWPlMN
XuQyFdjttHCrYwhqd40N/H6MdSxJzM0IM1QxWaPq+TqI2n0yPaNzOCIuU2f6+oEgfasDLWaOD1OZ
FJYVkvb796bAk7xjs/VmSkDKzPC57iLa/gN03f0OOO3WibkOPtQ/xFGigsPRFncwfAbtK2MX+2pC
I9bdscCmz0YLr70yiN7Aykst6bWEx/fnrXLpicz3rQ9sHYsZ2XH20JmUNSOrWCPGz87nDzzd4Sbz
qdR8qCCq/n1nD/HCPLayV/J79W0qbFWu3fpui/E0yLD3IB5ouOQ87PlN/c7IaK8fmnVSARP0LPv9
20Y4WfdZUVEuk5zl/Kj/fQNms2OPK8eDR7OVfSfgBRVXgsolZACRFioIHnXGbFudnNs9ZvuCLABW
0+WqrkJTBdJxBqVOGIBGiUwRypKOPJ0AlFZ0p6nw92CGsqGSqzcL/DI4Q7z78CrpK7LPfVdr20n2
QG8lF+0glmvWJlMaQby4I3BvIqugosihSOWRvFDp9wyvtMOzhJ89XQ2x+pXbB3XHM0M1KMh1BzPD
CdkQI8iHE8+FgXrtgKrEsq9Jo/ewW1am8gWuRGEZIEIkJ7tyv7nMM0bm2yA7hY6LQrES5p4Uhz+n
5sDlybMGb3vOP6ejKJ3bC8ZqKFfMnC7xXloDPjmLt+vrx8S3gpOPwmh/psICxFu91tug/qY6veoF
psdXkuqkZl4flhzWCmJu95I9414pF3w7UFrHJ06jZkW9DT+xApA2u5U+IxxG+Mr8I6FpCOVezmnr
s6ZiuoSMUy3Jna92ROjoYJ4ZfYqzTIUYTUsXDmVO4FQ9NUXXYSOmQ10lx/hyN3iIw5erx1ycdDF5
kRtx3t71dCWO6e/aV/b/2pxNWwiksTAXDjTkM/EMM6S3pn13vkuow2iIpuFEX4e3KKj6eCEkkdxs
rRAhuSvgh8gB+D/agc6wUYc2qt+znkPLWbZS5Ny+dJpUsKyqtEnVDdR1EnMfTKovZBnS3+NtSSPF
sjxt09niPHv9+HRq9rzGoOq3J25yE/yEaIUYjW3I/dAR1ycqnwQz6djzA7u+yZDrWRDHuNg35+lm
hYKIRRUOTtfDb7iayDKt+RdapFB+JYuhwdV8+2kw010kvieAA4/OGurWiUOYggqKwDUUpnMBVj4G
mGeauUatBGw0xtSCLNuFkiv+EQA04ZhBYVG1fxvX4eMtDio9DJiG8Z1kbNuETdjvo9FTpXU2Ga/l
+Gc3+ATS/k7O1gdz4SIz90zYUwFsALws+8bpjAIwAIBtsebkR1+tj0JhV1JA6g0sBLsoPX6fJaf8
zQZPXarRnsvXjLTKSdQ2ThayRYLI3tvKaywJJL8JF75uz7P2pIc4xn28Q0Uuk47de8+W5H1ai6pY
etju/tgiemuAbr/nylp2/btaXdqesYX0bHwc8uJGKEYvk/KtsswwDHNedVwyDslYGCEA8tEhMxRV
cUPWWMzJtbMv0PsidDsLozMQDdZeL+PLLB4kqsQH+rmjgWktGr/cNMsA99bTmys4a8f4/87to/QS
PCSO9c0IxqWssJ4ExZOBfJBtx2RSg6OrCnsMzbkrd/NuciaPitexXWw4657yIKRnCHnoNMXRcB0O
rmXwks/wLKWChRS4LjLxCqSp4pyUYOU8izZKUPmCo5pxz4GoMF8u2M80LrGW4bmiiL762sUyk0de
j/DowJ7pNla8tmzfDWJafsSvz1K8LSN4uqXtbBh1DZAaAVZk4OOHUrRp7zLUjFEv0q6WRmLpb+rE
rVYXQs5GcmcOkr+sqoRLjIqkby6OFqSA7wVWeYr+9+h0mRif08/AXJ1OnayrbBBdaG6zpNs74P1Q
neYN74hn5mMrmFft5bdLlFXmCxGJ+SHjG9wuSWIiYhhVDmybGjsDhsElo/AigQ8lLBuhakNa/KrP
34gttbfCJWoSIpZ41x04Ep0CSWct1KOJd3nYMpk2KbOcK1xtHfduHzNtx2LKxyr33MTzwHfytcYO
9ypAB0+9BuJ/RKSD/kPBbBuxrM/IX0CBvn3iIpjKhqW80qwx5fy5yXFUT9AD0w7NnyjnOQc5PCMB
yoaBchZFRAoPs6moOy8PGDO5DNkTU3foqTvZeIxOA429rkPa03CZOfb3r/WT/Z4c+/qaMR/LRT2P
VFuufKqL9Qdbh2tpfofV+DKUr+/4ftEzLhOBy4KKJZ+mVhAPBxLEfxLQQYrVxNF4DV7dQpzH6zq2
rCduZI0uREQFOqBpyt0fpz3nzQJoyklKLTJe4C4WqQ1PhTVP9JDjgTl1yGb2KvBQ1ps63BQ8Z2+x
BPvr7PJzxEUHKDizhnUcvV9x70rrkL/O33VbRFz9vYSSgXcxkguPo+cFz5FpQbF6LCs9bYxWTag/
rASugsBpHSssWsLlOEw9Ily50FmwrILNa72MnWTg2EzAhK3J2sFa5mC5ocYmJzJ1+1OGcfw7jYOn
+sD2v0f99iL6j/PDHFBkkAz4qMlMxQ8+m/eEBQ5Fj0Q+ZlUxUanyLF/sM1zOpmbwoEl6X1QaIasj
caqyYc+ELsBNYPctwvw6A/mmVxxG+o7+8R6qeNtJG56wucU/X5qwLdWOm5xkHhtnTCNrdF15ZzH7
G1eetZPzrjiv5Nd/yvA7yrQ02n16bCTU9AVT3ed4+lao1I4QaGdt8a0FYKySm283iL69QvgOZzBy
I4vzoGyZVx7+sV6ovQlGR/k/AIVsl1SWNsOMLoS7n96kP2fAvLyOod8rP5+WSXP6zA0qu490ku6r
S8N6dYWS5teXNSsUajojDQq8hjkZ703Z/rs8H9Z0nCEnGKhjbU/OJcnluIQQGtWvairfJlxABazy
L3yc2hOmOczjIr9sTqMPZPIwG5bqO5jszBjCzEn7y+RvvDgcDSva75L5lcXDr9ETOCJw5GOBWp+W
cUM798yBYawymfvmX3X686AxtN4j0mXQQoyjV5E/E4KgNUyrinxtY9fl45WfoQsSKJIzJgxLHrpC
RSF8+MCz/RBgdSXO7doYvAjc+OcGrwkM5LXKGPwOM4mHiAzn3oW2G9/kOdhe7U57HabSbmAYOnIx
hXrenLl4HCrfFmEPJrRAupTk5pZufzqB6duM+t0K+wYQY9av5x0YsCIuCHGUZvOWwVD1rOmSbuNK
fh3RcEDFPsajvmLcxEMpnUnTuKnbBtzFTp6uEeeWY8JsrCZC2aR3GeMOLsoYUy3EUzJpunZOkxxL
hEuBiL1wjtj9iR+EQ+MIrZKgt3RjOe55MZzcCLSd82P79Kis4HE/l0OtQR/yGORqG9LEGdfBco3J
g6iC6lr3y3ITfneZimCQyZ5y9e6oRF4NjYWPCxylio9VZgPe+MAXOveCjSMhIL+L5DF747sS7a6k
WKsAxDYshnLAGiS+Rgn0SxjHqfozp1PqD/0Exy/cKvaKNFcHWIzqLb9Ve0xG6O9MqmPJZVj6Sz99
3c1fjJOdFjA9mddISuTBAr4DyMdpLNvLlI1CcCYmk00xfroBZ+ZjP/SB0MBd80LrgqDDrWWzqiph
NNVyNUB22SAkfF6clrXiCRwHEkOfnFWYDLE112uNp5jVcBGtYHy558xnbDfmw+2SnwHLa08YBign
rmrtOhq9LOuhcyTnJ2hakgfMMdT3bup4YoXhJEebzQRcuF67v5e/fReoc/aKVpx2emg/0xgGbipM
YWbZuzadlmn4AEg1pqtQgHeiDFi3FHgzcdDiVGU4Z7l1DPkjnQ7ASwIltauhMfC9iXtk2+50SYeK
zZhgyBr7/liUBs3YShltabHrcCvZIUBuQl+YNYY49YlSfS5cEoGV/n+x0DLiuyAVHr6rHAChJamQ
bHXPiCJHG2QowCnE/3ptH5HqZYuwvgQ+6k8+0ECjICzvn3RR0zSlxMHEcPyWSvfv+6Atjk6vdYgX
Xp5eb6RLvWBbTJN0xxBJfEw7p9s7bpIzJmL4sEesjTZnP4TPp3N8hfTTUP1K2nJWNw2yMGgqeIsL
/mROy6PMAyhwpv3OVF+Nq00aAt8zWMEsfSad276J20UdewEQAx7pPPpJwJr7OiBRAQAuArD4Mhif
dL8O4Cmy3FkZZ6EEjl2KIOJopb/Y7bgB6YFR40UxMw3ufWObXpMQVGnW2TIZvF+PeE+KBL7GFIt/
cYjG8ZRRTk8WUSwl9c+Ss3pu8YHLicyHW8S904nhHduuWFO1Ez1vp1QkxBvrFSyKR+8brUviebSy
igtTjuWL9X2Z4idfdP5YFpJBOE/8PB0zv0mrqDJP+/A5m40ClcsVexrcvRmK2OmdfGE0HDvL09HY
KvLU2Cd+bAJ3bfbUdFppwHYR4VJiQBTXWVeyKwnA6GbeZixCwdrIGQxuYdbWvajx90Iz7+02e98y
RLybVtG39OE+HuM8bvBem9VdFjp/kmzZAaYJk362ZMjRSG3fg7bPdwjcT/bz57Hgc0R+/ycCQFQ6
xlv8I06jeDqKmlLtMIKPIdXNIunlUeMG/DOCwZiYvH222qnw8PU/HEXyFHgDyid4PzBhXSuXxdt9
XC521BkUzbBMT1U8bAIRnEAXqdB5Hz5WHSxOUk7W5ROwzR+KBF3l/ixrylbE+CT1gLkpULnbez3a
nHjnUuGDVV/E2B91hSoYK1tTqIgPk03xcZlHDI7hJzNwQC1B34q6gT7NCjSUIovRkYYAHmF6HoH9
FkK2+/RKezBgORhC57QkxHk1sgAW8oWkUv7MQViu1pNbZ1dYR7HEQK7D4jRHS6XVPrsQXA72h4ms
oEvx8i4v1z/op1k6jzWWB1hlNyN1P056/ox+tWWlSmY6fpWzG1z2RskkVsY0PdMobdogAH523Yoi
WlF2B3bSGVF9N3gGthi4zSFZzBaSG3MqrEEE64kC/th/3JA2YXaztZRSS0kUP3phcsvrs4MxjioQ
2FO8LpWgcUjlx2e7Z4slBL6Ut2menqp/QHgM+CJUH93wRwX0uS6eR8Sn2EVxb0IfGSpYegZdT1ZO
gwSgJK45eQJKKsy7pCQ8IzsjTjvG3FnerFG+EEZ3iv+ZB6s2kYeIxBz3nrkB4n7zD+6HSgY0JzOD
DTBqb7CtDX6f87+syM0jlxJNNDnZ2km3qQyumM6n3DOOQPqe5rfGcIfmNaso1/IsKM7Npsf+UPpS
344Tw14dzBJFrKNgdwV/QzgtP44Hhz87a7RFTRP1+GdzdAq11+KZLuEZf+uUKFfWID0vlknK6OKl
RgwhJWVCVQHcOA2ztVjd/BHJDSgd2wnVp6Wed714DAkCLH82gDc5H+UB6WiX9YlDUqJ+d5RFsYzU
P4cfcX2dxDZMtAWOveG5p0dsOGna/04OVivzIbt3YPwHDQkj40XimD1Tad+lovdTXlMKYuF728u1
buePfJZmTxQXG7KKXwF3FYkIIrGBoc7BDckz5gMWbDTrpEoxBw5NtGfLzb88Xp0Q1uP0WsBeRS16
HfPZis3tpSxB3xSArUU+elJUB7KsMW0YsOBXYwPFn0a3SreARUWz2rdv0keAJfCgeSTHHAopeXs9
wS0aRw2gvEeZvDkWLU876+TNFV+impc79YSO7yMgzmcT+XEwN/EGtqNDcJO24rkJoRAo9ISQchdh
nmUWeg/2NkyhSjrGcW2X1BuF0SX3uVbuaAfQ/UKuURFgfNag9kfgi9z5Ls2czZ55jMO8bdnX31hy
PLiCHxKlXoGkpZpLfCxukHJd4100Svw1pWY6n3U8G9jOBCss8DVO5e/Q5svQead2y3Njv8SZvmCP
IvBraAGVNXwu7m/dlf3bilqsJPTjruksfNqrpGMhGOH0xTZIQoqyUYteKAq+V547DTBaHBH1ylhu
X30NQmo/rmhDirJp2US0IpAiKKBKTpcm9CaJMl/WN6JKPmrz0H0Ur2ndvYjmJIqEtycu2CPFu9GQ
zFfgI9ExRvBrckwp5mPPD/VbS02NBnS84r5ucCstlJ9fKXXCwzkUGLOtIfxEF79raPZttIjmPRpY
KgplwYdQFt+2bQbmonV+yTc1XDk2/GaEpvZcx/DbMNzW3EaBzxNpOrAS7/VTpC49v2pEYUhipBP5
3etBNZyyKQ0jcYxX4UolrSDh81OquGxYGteMahdSMx8acVUxEXdaDjrpZvQRKdKTElMvAmwpEEb3
nKQ+TFIZJzLZh7/ZkbCbwW6XNc5Pe0Aw9Xytg91Y/McDGIPmjF+mGhQ0M+qI5AnBfOU1N8oaSlG5
BIKLuW0mK4++cmETcymFwQjvZdtXvQJYHb9Z+u74oy79nM6a/CQmtCRm7iOp7LP301Hp26ikwChz
NoO0xGopEggfoQ/Ly5Rk+/ifFHEzzw6IQP+TX1fyaDV1v0/DABpIA3P1eBNFJnOumg9p2SJwnWZ0
3YXnF84WcgHr44K/FGKjlfhdjawnj5RMH/OLm8BN5ncNNToVqNtvv/CBZTetlnSe6ORIj0IPSPqa
ZLer9yg8vUop9wHAAZwioYBG7uueLEyeb2Am0/dtUB3abbvijY6RbescCihlMIajGG76QqqHeBSx
/zDZYPyW6n5BRBalxYWHtb2+0Qw9glQaUZS+/s3cQ/K+QMIKlAZ921IMszKLb7/Vm15ySq1CGSZe
2XHzvIWMmL7Kh9GiFp13Dd/C1JyvNFJxn09rd0vRpisbL8OhLInSw5aQCqtTLIzE0/yWQHfcTTu0
wjbzt7SQjGGkK9zHENa2bI6Z3wYO3LfJmFrNBIWoygZRnRiatTKxDQcNg6BdKaFn1WOi+5gBIdMH
RcGXoQqQpIrTBVjy9r9/73blpyU7TgJJukCxNfm53cHjPOsMqeVF2rWbpYXujZFHnkW7nWfVQvHP
MNLMkNNE12h2/2htt92oUTpbrD2AjAJ42gCeLbJ7R+ZepUL41QhhAzbA8eNV/9fOx4kKrF606wD/
Q48Twcx8Y47Z2cygaYgv8okC/K9lbq7n16kFGx7pWnBXRP9V3S+cmG4hAqTTTE+5i0QRXeo83ZXf
TrjqOp/SPrtBwkGvcVGZ5T9qTRMLVIOaGbzsTPsfbd5w2tqGdEmcopW91Hn1HQ5PeEt5hPvINLB3
/wCEBPhVxLKfc2WTmE/eha2c5lV/DOqgs0qt0qF8CFC/URh2N61xXqR00oar1PURTromZQEMrfaT
k/Hz3poIncIJuU8vSBq/6DWKKispPgejgWIykcnGWugGKnHpaEZq2lo8l11UDwsCU8zal9wnbA+6
4b/YHYrJEmOwmGA6zZFzXg08W0i6dHxtKhQiZ62iAXARkg3sfr3bB6/UVRYHThcMObCSv8U7pYsi
eRZM/RjNF8FYZhiYbIIUNOMVqjytAZBhKng+KTNW4+c72mJrrWcQpG2K4fesO4ciNEno+1hfWXmT
zA5yC72lYD+q9UbUWQ6yL6aRqnv3x3303h295w43yycyrp/il2UHm/xlMRX2YcxjXz7/MMi/rpVr
osMKX/HRM3qpliImVwAEGEzZtlHGujxt06P1qjrNTWI4b1Bgl2CX1IBKli7jhHMFMLsh1Bn8gIL9
5QGqDetQ34eoBU3fU3qlkyTF01oBId1O6Fo05CBA0PDb0DOKfjJ845mtBwjacdsjuYFRHL6tpUv9
22GhDR9mC5XPoT93800W11fi8p9CxLN8B2zST/tYfz8P6lKNvYK7tj1d04XZt41LFKHIRxG9YdME
nMczaedPoCzjc6Kz+zY+C/lcHt+Q0szxmZKJdJRw5ZORJ6ZsEs6Pc3Qy2vqwdItWDzwr5Jfp530+
QV7k4nuctY2w4d9Pet+IeVq/0FVka9u6Yd0PgAB/+EJoPWv5ondxUEJMFpO85bqJdQbGM96FBKKW
U6tRAFeWLTEa1EGlrFCaUvz43mUoZtYnSzJF1Cl2l2SJWuGH77p44hMWht7k5LHCErxJBq53jEe2
1w0IEF0H7yhCz2dHD1obp1ENQ7slhJE8XWkzFMzKP2ypns0Qp6LQzmiB+JpM7EjenaK7NA4U7POM
qnFY1/vzUxnplmNdwlyR2QQbep2mV0Q9IsKU0vheBvvlLtO+AwxtN6DbopfsGzLyCf8EanqrYBtX
abahQliTwLJrBAs0Iwbmxi+I7RnnfVEHzSx3tq5+BEyMoqfUU2wDv6SJVh4X86C+gTTXE3qgm4el
epjNnXGIegTz3NmUTyyr/GYNyNVpDUeo+Jx4GZcZmnwtd0lGUvs0/7FWlsgL6Ix/EYm/i22PCc2d
WuK7AsL0SCbwwXQ3O+QS/vh8FSzksZITA/DGkmnB9+/loCZ7nS4ih6w3GEoa9IAM2+kJKeoFi4Vs
YDPg1XkdTRKufyvf5+IhTYsjHB+5ZGQelnfeigdyE+0d05yMGPCr8Rw5RNYVQTGZgSGkT+VzU751
mPoxbZNEmIqd076HU6d0k5k2fFQ0INRy4ZUbvDshHfubsmafJsYVtl8Sh1Ii40nNzFWOHcBQQmV3
w9ogMbcQ+U5SdRG4QcRIkGzL/THxEp0JZP2/oJL/eKWlxmYZTj2NhvIXahPabRvvhtWwI6RWv2V4
sO+gppUUEWU4Ohcryz3q7GnASmjffDpnBsDHbS4C8Fxkfs9o24MmRZoZcyeHSUy1iic5k6yghHZ3
kWu7xmlm/qRlwIqcgTjLeO6XCOjYwLZwy27kg9tZe559OsnhgvdHhw6gkZCg5q8nrbYdYB4wkv03
aiFdHqSGb+1FEnPJ8MSYEkhFcu4/IDofwYTPRot2ij40rmhl/vZP8XK90NOq/z1d2WHjxtJPnNBc
TL/Ggxvq6O2zcbAQrSraUsCtCiXEFaWd9Oh9uY0JZ59sgdud51hO/Y+WxudKo989/H6kdjCIlVJu
/KqyCCuniR7ZNU/q6+lCaig12d7DBUFBR4qkQyapJ3DdsSeYIpkZ29JKP0obLxvdSMr0zn2VmwZL
YjrPJLo/EnnFpdy3MRd+46mUZ5rdz6TpaM9gINGpKGFNdrcHTkQW9t3zuXQ3PPHkXuAcup7Jb4jp
pCTJc59keUndZDoUGpa4YZr/yi8iH2yOOz2XmuolhzOcMPBrgXVLDMYiAycCc6JrTcHDwG8rpu4b
jHtA2/tQP5TLgqn0zZd29eKAtlSywo/vwhlipgUeriaMtzx23H1ZIUJhQEzCOTjk80QjH5YTnh5u
JzKiq1b10axyaOfO7QzZrCJZS5O78R5ijq3/e4nqc0zDRb4nCDKTddV/Hu+ioV+FGrpuf8o0d2ua
gIq/XfzOwM0xZYZGKxFCuff9xCMnxSOGW6Frxhrsxf+5PJXjeYJtq0eZkOjCE50uNwmhkPLa/b0q
7wShVMCqbNBkjOrvPq4Yd7ou96jdi22yeoaMMa8TpkgHeIP12ciyClSr+Qf1zlIsY4TNkbVE8h7c
XbLnFoXG9ynv2vRbdjRlepwDDlUdzhFvTvx0dLfkXPtlWuPap7txM0RFPG6bgvXJ3QXvK+1W6ShC
ExH3+SaQPsZds4wQofAQ45U64McgXn8fq0sMbslxA9o6CHQ2ceYyuKgFAKBVDQC7l3B88u7DskNU
6MksXwx/r8vPfCS4p5hSt0O10Wh6I4W4pp83iy0mcoRSPXkd8kAtF5WXWmaDN8/XdQZ/O6ljF+bp
sj3J0YTd3kKapUMHocA9VG9qWjzN0xvgkDRwC0PXAcg50vbHAMdHb5MZsPFWsXCU0lriYMHHb2rA
GCgDcs1pZBZUHXozwskg1HKZHZ6TBPNk6ZkAO9Jw/hdWurXBg9LONdOngDsiBdslBY32TPqNsc+y
ssG8X7dn6L44joVzNmU03isdlMJO+6PsH108YWbzX1dnY9Ht3L8R/G6+duBpqYlaEeGtsXtKuaYR
RbMdMjyi+Bh84hFPUOmPeLCWoLMvlhC7PvbXB48lrN/4PaSr8RfceOxgdXTP53Do/3svzFlg8IFw
wB/UUTVBBXjYHeL7WjKfYw908tFuKJ4YEhV7c51W91Bd32K9kQMl7IPMrAf8RaCmfpxf/s3IWdcw
zOKp8pHXUxq0vWOZGHbJC40+ewuSavN3J0p6pxAOayZbYulCcYsdMLNQSPutEKk5W/l+V7WF1vuc
qii2Mjrxjd8aCBP67+lGMjzDVoqZ+KQHarh9kRzAOQiJsRdQaxJjSALcT2tm86ZKdZb3C2UqnQJL
aOptJlmBCQr6LwjTTHkGdvtrFXGB/YQHiHQEDdSCKuK27pWd8iDDw0gwipy4rllbSZf37oTy5S6E
efG1DJ6/XGPDcSSllNAhlVp2Az0lpyF3zS1k2k+O6ZbY4McIGOOZqb9mR/QAEsq8eTZigL5yH6Nb
c0zdIMxd87OkKmObZzLwEkhPf2MxK5TiNn7kehfStEey0ta92gT0701iaBBJdB7d0Z2HtDZIRxcP
TMubyOblUKDjg5Qro+6RaGY1UsX0W3maZ3AL0bNuVSaaajYhB/VLrOFexmYydY3oEW3bQE5QgooY
7glWnErwF+XCuP6W60keYEUgZFXjw/ZO/jEdup+iHA35oMsMTag9NtZ1b5TgcdjTdnviXtpjVgmu
Rd56ufELnyp8MfHScA+6IHbQk1Mzl9kkFENHTK/3A0oukSo/O6J2T7YTaJLi2nwMkMTuRrAIsxMH
GiIwC4vo55hnKk6p1YIsXfRItLi0uxZ4eYKz6h4FP504U6VDUGThs8OB3ySxc/lAgwMjpaxJPclR
F5bAERKVf6laT3N9tVRxIMO4E+oxcqKAYXAdjpti5nykkVDL6PVKQLB8G+P8cuM1hkCpHjGCaU/G
ci6XgYOG99d1MdXxPviAFNiylKW4cgc1F6inrtzFEyB3n6Q8OOLyruMgwhCn7oP8ayNKdGchALQz
AtUpNsu3vcXTPClWvWcR2xBV5WYNjAQrUHxog3m8zHi6jSZ45tVHeRTugNeVPm2C/y4bHsFiEtRj
MR4Em5qFQk5LfG0NxYRIdcbKdW+OzPXflD5j+cFjyIWGq4q7VuFA7mHzmz362QNy1iWNiCG+dwN2
uR1QsuPPi5tT9htMW72k0RVyi4c8D+iAprTeLTU13KdwSO9kS8fLZAY5kTaDrTX/geUodmP0a7l0
W2oA9dHx5Z/gk8JQpMph9KwxVeunGyUqP8sLqWiRqsgcWwSL8haCij/LayU5njOew75dre+Ipgdz
Cdxiaxz+Mci97bdY/2oQu2msoZpMhjIWvcS/ykpSFwPzonCRG0LcsfqnGqdT1x8F7tCJtsWhGsjp
TfxUNcXwDSJvwrPc2vu5DNwEmaM5F8bG/B5MVFBsSZkERJwTu6cZd5S9KzQUxt9grU+VjPdi3tPH
YZLCGKPTK3A/piBTpkihSYN2tlWlOnVzUxtbsBt9wYV/zRZtF3KLnZCdQQfSp8vp77bBOPcJ+3q0
corNvz4XW6wHJoiySBLHlgpP3pv4Ta+PpUlz3EfZ5l39pEma2fb1X0apn4riN6Tph4ip39Ka1MoG
BTpcAaapinjS05vwB0Vx8eMO2T34E37aJwHriyACtROfRdud5rg+HIbhsCdPrOEbvQzVDP72R1SC
P7lD3lJPNJ3jBRG4BOVuCmnWokoxxbG0WAma8Y5UavmyQW/d7i7zs/VrmoMun1wC0rDfuPLeBl/M
PiQwg9hRPNaBZJMv20Driyvq+ZwT7WYJKxyD/jK3t8DndEYZLLsDmsGfnmMgZCXrrr0RYciUuWbF
sOloVYxL4iL40PGhrHQwq7W5M1StzirzRb6U8mwQuHtOAJsDT0PiBsriOZ3OpfZ0RrbLlXz84UES
6J9NFOUM2LcX1O9m0jgCu6S+rW/BGTHyMa+bT9XAriXrSdah+Al5anO64RrPvtJHnAUzb1N8yOTw
kZvvJj0ryOTISw6QtePQkXjBoJ4LCp2o/dhGklkValKt88CXE8wzzp3o+2ihR6PqWfykqHR3UyeA
BnWIdIBMIULShsmpM7gly4YBxzwjuw674ZabDHPF//TAst8uR4zM3JXk5dx3wAdZh4Zz2COa0gNF
VM3Xj4pfPXFsc1hewxzEIMZTPP4igvFqXYv+JuSMM+gQjociCRQ8OvowxBN6H2awCNALLo19o7Tf
eTa/Lk+ueVfgKf/GrRWp0xc4flzIi9l886Nnfhs1UR6ukJs/IsZZnPyrZupjitBGDmBlbcTqZglQ
tDqY13VofrOUx/ZITUZyaAjYlDPhN7iftwcRvd8oG6PgHb9MnSu94rvKZlgD5oP3BXX7cmRoDvDl
LMBbkOgVknrA7wcAflLna8aCGYv6qrkVAss8eMGHOupLUJdep+1a4135lQPhn4V3Y317NNoTVEfp
VeVejGGLjRi36Ncnldb86WyWQRW6+14c5hyYMeN5iXioh9ESk/CiLnCfpWWfIXM7zR3dy5KlEQQg
HCzLL9FZglCXtOlme9ifh+b+a1yEkgeyBGs53JLwMhWIVOHRo9CUKd2ZSmzSJnR56Kb0B7aXUCEa
ApbWNhSmVAETseT/84i8LycErxwx8NcgRpDncSTlcdadj/2s1fUGWQSftiUuDsU8gKHz9ldYBw0i
v5OdgDhM0YedFijtHaghhhvRBpy+9u72wvUxlLnJk5wozWUGq03N/SyohnfQgBciQ1rTPjBgu109
MObJWJYBt/zFlI9ZS2tz1ZsDBog7PasSlCkuL6Bu5jxtjEf2OTaJUQg3YMgK5fV633ilJrKnLEQx
ctC+qtE4H1FYZ7SECVrBNhM5x5J7gg5hvs65562klzCTaDAtQMWnoJuanzGmQvldPqWcCF5Gz/0d
AAqV69WMHP3BAlrY4v7Ska7jEmXXWLqe3Vft4ZdULjfoI6kV2DRZV7ULWLWWccqQnVsQ3pTbwb3z
2LZ+IAD5fi0UQBfecEKaLFwJMZq6pkjZ/S8MWO4ChG7XbFEeLeU8LKmX2uOFvcU5Us8sSAjEN7kL
POoi/7tl1D97aLrg6+SzCB+4N3J9/XWur/X04fVYFa1qe+9ShtL/3viSUs4xyjeMBtWG/nqD2IOS
Sl8MuvUvvpXT1bvRXqmU92Woq/uQvMrV6wxbyd8FTSthsjxa10SGGg6uZKzCGNSgKQVZv0PSZ3sK
9AzPEMZoXEOby9cBXeWHIPz6yyQ+dphzvgVLjBcyA+M3EsMxNJAGUlj+XHN0xdg8zEUgSOhR9YAq
zd6+/a7XAWudWJWqh9IPMXodLR1zrhTBuV+KFuKHyA6gcxpcZkWDoe9p6hvCVkJSWPd9aWnIg114
zGvs0b0yZKk9jm0MaRYzUDHOb4RH5rUU24EeSEdxCgyr8PdidUuyV3GVTCSiFk43zf+lh7WYwQUK
9Y5CZzipuYlPOv6cm8oOy79m/EjF+TKrF9DNZzFEUmIPuHcr4dfhxCi7WwYqIHUHK3RmxCwIZG30
R9b0n/6R6LO617gll9IZnXnWvuYQHMe0ZGdGcCfrkTqmjh4fMTT6snoeQPiCMNjzQDCjA2+z/eup
UNNCIvQ6G2pRksRnk9gWSQndhr7qPjSHmwI+1YyQqImkqOvVyaSCiIdAaHC50WerJ9KfxvCdMwVS
b/fuxC6KjZ77I6ZAufonCFtCP635LF0ArokF8e/N1KVMeS8e+yNB9t1rglXzHZOiLcD0AvO0I/sB
D6orYj4gcJUjZlQ0kAwuRjw26wXVJcnnILJf4SvNz0pG0g1WeequJE0gSXin3La+cA7ePCg46tmA
AutclQdU+yWhhKtMZrCAQWs70R4MVIng9JwTDjVWY5RCBbj2SX6vQfml9rrK7x1hjKuf2fif/ioQ
ReyrVsJQE/F56q66gQOGYYFFwv4HG5Eu9HQcM2cFuC606DhkdQTiMB8E+w6oFAfJ2vNl8HrYe79n
Zs13vvAzsnQx9N6p8RQZ3FoiWFHb5k7axqj+uezh3IymsuC/XxVoicwBdR498/auXNTzPM00YCDw
DiaB2dts7Nv1GEf/shIMQpB/6Us9etPwaEyaj9LLpeSfYZ0tEU6JNL+cX2c0nZj4Wn6R9SIDAdeK
Z4d911ZboQn0KleGx7lt8qWHxVewGz4/sk96IeAx7xPAGJY4BqKaTOzcquHoMEwcwK8gHhZDVEFM
BYuue12Zp4R6g5VBXtyXdVFtE7ErAPeV9Fp48dvDf7zTMuaShLdm0qhweSkpOlRwvZA6ziCKDipA
4mZL1m2sKH4r3kM2mBM/TMewFu7AUsW6++XycNghTsRmwktjP/ZevpfzWG5MP51plgyY06uGv8In
iV3CPKDdES1RFbclOftAqkEWQDd6pXczgE8gpcN8HgTXqvxPpQDYFxI8l0a+Y2jqkljH5LgorloA
SrwN/2L/4wjr7a6sD/X+d0I15VmwcMjF6OZ6CoJjPG9E8zz9uoxKEXG0vKvxLOeQRoFkXesM98zq
sR75DwwWYN442VBai7dJ4BzmzDoynzafqZnO1trRD3XWvUwv6FEJ8hVJkF8q2xWleNbCRuf5EKGn
lIy9VNqZzjdKd4304f2LtPj7WiW41FkcfG/Y6AAD6cu8E7WfPecDvk+Hka32xFDzu64V9J6v9I+f
F4EKc4t+5yiRbE80X7RSIwCZ2IFss58L/nQtaR92sAbyGNMGHi6TFVbluBBDZR2jdDygE7DWRFDb
5ybIPIqWcbysvkIz68lyvMP2zWQ4nQP1RekUPDgCJyYNx7sQ52CNv9esDsV7n7ykh6UFS+bMIJiV
FbVkPfPqEpYxStaJCMYfABTGJkbo2aP7a9IHtMU+KYVWeRt9uNpIqa5pdKsluZJzqR3f44Fnroc0
Rewlzt8cx+SXMqJS3NvZNO0WWxuPDFmQFBbawwpyxu5dScK2LIzn5TiKzg1SyLL7OHekMFfcoINT
MnYhJEbN8rM4dbfw0HRHZ41ffAtr0zfCLfqOkfK7sH7WUv2cV3Z9eUNX68feJp0KfEQhdhZGdpzN
yzOPNwxFw0z9uShg9B4w4OuofjJjciEZiYApvydvPc3UFLbRVVTDtoK8Hz8EWhKl1WmpQ4qyNRTv
78uV8xz8CvB0jIRqfgAxfhCCEjiCKg4vUghnuUJiR25OdRGbmx+RKehHIRfSjbPrVsNWl4UPOkvj
R6whH5VxJsvQ7+v82HeWq28aybhH1XfKQ8RNotPQ8T/wCYmvaTRBZNHk387+2bfd80ofdjvdIdB2
oFczqiFeiBzl/dRFF1v4gnz9sWvZaw5JuNjjG27VTWDvU+DxXlFiQGaOXdwpXTpLT2aDD05uXeKl
YPckZ/xbsar6qK4pO0u/spg3PUycPOVUcDIMRT5GVFif8OibVleOUi2wV7iw1e2Ysdxtwojmykdx
nOJvov/KnDq0PUNmZgvL9/40TXGrIznmQNrQgAmz4RCDb9r+Pw6fHOIorLUR/f7ud/5jkLcXH6pX
s73k1/pBI1H4KbGHRMg6TNY+70tlWArdySRAdMCGHLK/qwsUHD1WEqhSSCZu77fOyCJlhJiLY2Lv
fE15o7533M1wggXMRoYcNfgt7wdMVNju9KDYf0klIDvJR4no6cnCaWXuPlM/qsH3lVChBt4Ow10X
j8WXGRdhwHtcVfYGM6RfQqPrs/S7LEITUlHWC8XK2o/qrslu1tBm2ukIEE96rG7NPqfgfcwib1wB
Z1eysSjXfcI4JK2sgGIRPy7ElA1vfOZ3eG1z6CmyYayU9zLY88gULYkh2lgpyCmuJMOJeieQXbn9
I2hVH6/iXWRaVIwCXhwTYawEPbNN0H7/5NxpYjir7O/UzTKGn+EXXIzFqbhLrMwIsNeiw0j6KCwR
4UFGi7XCROndAk40gfIo+dlfkS4Nqf4nvNgfg2Bz6ER0yxy8r7a/tiA6dhTq/7+Tn2mpSsBHa493
62XL3KQyGqZD3YRg87y9X3OjDv0klSItNbvHPwhEVyhOvfI4t/9VZ1NUhWoVp2rCrYLCqxjj0H1q
LPh7n04LLXqK71SJ235EzNpGmENSwaVXBgsYqJZ2VFxiBtgbnClqpO89pvBeGSZk2zdodDYGbabz
e2RwDUKOH6JetPVA48GoczQzusMuLEhw/WFd5naak7svN+IA/xQlVz6uaJ1hOuUGymfzbR6moPP8
N9+n2ln3lvca/dxJNNFB6yaO+ZnUTZg/kydK3LU6f7+Q6qYTYT2NIm+s37ReHRhGSz6lkN9aIp4f
KEgBpQA06mHojfeeq3Mv9OHd1uobrKzGWltbndEPNVnWaF0mpCU8x0rrKprZ1zhJ54qOz/YanG9L
NRFpfBkW84vYQA3sWcWEA1Z+c0dx7Z6emQoFa+/pUsVpaP8M3aYgr58VanU2jcaGXkB7bv7W+nrc
lc4NOdFwQDo3zmsr3sgDtJkr50+hDyMBxutwR4OCrqfo+4ijiRaYTF6GKtdUcvUKhrmEs8nD1WVx
HdkwEJCtYwOzCMoRn9/gqPJXTyDaL44d1HOWVgpTCdcByOy7axQL4Q8LLrRNtTIlVdWi6YVl46Vy
n7EXCqc7jDoswk5rbIMJIYNdncth/PG0lqIAfdrAeueTzyzzlqsN4R+e0qqRW+aTwqkpMF596x0Q
5GgfFLqDwjQHw333Oac+vEhlvGiHxfUPIUzhOgZkJtfJxExLKuEI7F9ujNqBU9NQTvwK6iAd9qm6
M4TqB+Je5ZGZiT35Vhq8Xzwyv4K434aaIbIaisLDo7mtE1ighB/jS/WvVaUQIdlFlpKLojwYY23h
7ezHVQ1y23m67pTloaZ3Aqr9VJWsRu+I3uuqU7dRhqoUfu0YyMtTOvZmefXM6mcaebJQ9DfOtGiV
aUz0pl0TTXyKfwaV0NmcY6w72+d11730Jv2QyF5pHUvPOimfqRrxdSRu5/7ixQ45JvIHbq24FBw0
HmomOgZfQiiD51qMRBYoBhrYS63Ny57uph8MIM43qBeag+u/aYPB0oVxRdU3B2+SKA0s65lEVoUM
ehP6XqVsZZnNnGZv25GNFQH8os+2B/lX+SiBZT8gO71Gq0AP0ZPsuQHhJ/MdT4dzgiI0GM8YjB1B
Q2GVHPJOBes9k21/pMarhZ2mCaazkXdj8ZSpUO7v4KnWQPpkjc5yzDRD/Aa3OMCEn/pRyVVvBhPB
Jjl6l3CVIjzj2ziJ8S00TDwTP5lVntjBPzNS0gcD0g/cih6sETiztj2gWA8JNe/3cI52fku+e0ow
Uc2y0Dp+rkUfDKJIosp97mH7gWBG7ocNV4K/VpSH9HE7KyK/ojXtu8XM1KUyyq9hBONQEW54vXSi
6u7QlUzawSNpEsL1DZp6JSpKBnQXhovlIdszk+WTK+6AqSSqjyglcnYNqxi0Q+FC4agqtq6PTVWJ
ieq5qXfr2mbZbh1wgrF6UE27f8HPRLqHvqIejfj0aL1YF9d0lm7U9xx5HIj2y1VfU/TlTLh3yR/j
hwtS5Rz7uXn05eBFiZK/R7W+t/D8DXImLlxhPlxW85rZRWAxkS90fKFH6+fy2dgkTqgRs0UgXO3d
rAUf5423lP5izwwVET8VwNOJT4f96KUIJEo2v39T/XLDP1Ercd0sba6lCOGEzlRLRicvZ9QyMSuo
30aQT0SZqE0K+5nSqRGKUoBBYsDW515I91q0sTIIKILmvL8R0VFGhyilL3IKJJPNOJt18jioyhJJ
m20ldQHwSpdW+AG9HCkkSI4WZHmSXZbEgJ07PU9efj9iJEJ92ZK85lqLd1NcJJqTpS2TUJ4xRxAY
kKEpVsDkigsh/HyjC1VnH7jK0h45ImUUnZ5v3ySxGXnSJ3a9YBtjngXugbc7/g2P59hti31ra4Yw
CFAtXJgAdCPqwmRHloSPsGK5tnoR1SeRlUvnpC/XFbT522u91QRSkRuC3/tbWtteXWHwxgraptKI
KQVjKbFUSq20/r+F7sBJIYvoIb1eYGdkNh7kHHi6SOyqQeUo1BeW/Vm8SVweYx/kUZz7VXH+YUzZ
+BNJFrD9LDWe0S2jS6B3GfxKQiZIMSN+qQlRwL0kmUIfbnTXqPs4Mg7O3LyvWrQiIMIt4ggFjZMX
XcbcKK4ynxbcCpn5yR++mFE1P5naXYcW4HC7jF2ERW37IRqHP+dkyRKGF1fb1XeQWyM5YloKRulX
LP80d3eiiozXtNpDUYnK+/QaqehuWJxR4fTbGbfpkYvybsZvfPi8mUQoR5lZu05I6jDmURz+1Ewa
3A53qNyRd3r7tTLBaCwk7H7PgnB1EhPDiIVTOcrPhf2jJbr860TPN4ZFyNgwzbXj11vv7XwG3Ey8
hi5G7rpoFOAzQlPup0YKDx3syBsbnW8fIYOLd+/dokHJxXLQKFpjlMwNzp/xPbsxnOJZsuP39pU2
ECd4QD6nvXjelZIBuHWDwLQplRC0c3TkZKDHih3rEZYf0Cw/DukEShaN0s3OuPsEglPfMpOAYpD8
cIcPzGsqP4MfZ867OmVd8o2jr6WOpznvn126/7Dc5JvYa36G6UD/gZCUeeOmEW52PGSyqU144yvN
AgByP5oo6U5XCH4DB0F2OIYlGy/k6/8/sLolizgKe5/KvRu+j9xikJlf3Ti6iCJ6tGbbExOi17uK
jtK0CX7hA6EIZhVW02Ixbf558XsPEJJXMyy3tMqCU8L172i81oWZYCt5sX7TQ/4kuRAqC/2zteDe
b/bIc4kOODwRN/x4dUAq60NF/iO+yeMLQ1JfHFKKKD5fFJftGYKSBkBSzuJGe7/7JrSYfzlJk066
ptnAh2uEr8ar5DAlfJ159kaBfLesznXjymDO4TBWuXmvtBQ/ZTv6MDQQwvk54sfOLUKQ+3xTUMxS
Lu5NHi2JTtBI1G2Fr0sBCiM8iAtTPgkr7nT2NXStMiFLdg/rsON7rShTQwRko2ZjPWIxkx0ZkfcY
VY6grT48DL3lqVFyM3qbT2L3mxVbb5DtTYkiSz1tDl9+dZOeemquhTXum+QsjxtCg6RqXTrGXHWM
7OOrHLFQpy8rIJedL3GktIK0XA0jZOKREoazrZH7oIlKTaanrBvuiMxReexTUXlVw2/wwGT0CaaH
3surU5tsCTrIFeyXCmKx+IWtGswdf8UDp7cfgJ7fk5Yo2ZHSeyuTxwJVwIl7kLF017FI6oiMM9fI
NjIkPpalReuFRzjvcOaQ/yoyccTPDRvszuc134PkRZ/za4MWExBkqvSIpu5tSe4n4QKouD1Vlgm5
0S/cckg8VZWnAflau5FISZoSGEYNVmWEXebz6guQ2lf2flr31Wp2JAVPlBJfcRNRUX75E2mvTUic
bRc6n2S5yHUTNiIXpgdPXLbW3UZzI0TdRRsxslU7nnvpS6rxTil87WaFDgq0XFUagc0L46b+SHmm
AxB2gWvZDvlCJIDu3iWra0VLwpqoOYKK0I8J66DAs1xYmolKk0XzG9wYxsOtlA1fl3gW4ISK4U21
w8BSlPnjhccqb8FujueeBa2WF3jtypUVKMAmTQClNHY9E/mn7yc5+Mg/PAk3ze1fQmlM2aA0SJFA
Q3FAPI1gbz+vNVgEWQYwxYUpaT/X1WPNq/qny1GetEgULC5NhIrVtY9McDOQ5b6f5GjLYxR4947F
PPRWhbIxvyCKIANjuWw/dvk9bWRdTZoJiaiuqqnPr5futT8CVH1wLiTp84iHWRjsT6/jrMa0rzSS
T6TID+lHtFDEqHkMWqIGPajXxwfHzf5ricM4z+6OqIuIKVwlSFX7I/xgS0C9MljMcVaS0+2pKxXB
qWnMqsjlQg2e8C6h/3niUxQSF3E+hTifXV4nmJVmd3V5Tjo2o1RBssLe51pGTbkpUEF4jz+cJ9AT
z3Q+5Oswz4CPWJgj2YeVpSOI5gVq/D2fm2SyogOSdWl/MfukEReBfnb/9Z+hiPAGp3LSmp6lnJwU
8dyr48Bl6OzheAIGx1CvY6IHcwzQjPT8R3n6Rx1ERv6Pn2ZRKSRl1n1NtjroN3mjkANVab6NUSaT
2GifI3HbTMjqaaeFcnhKDL/X8Jf9TRN0BPE5pnKFCxsK23zY1DfSS5B4RydO41YMBq1wK0BgAGdD
hmZgVANHInM9YC9dH4tEfrrYpD8cpL3AnTTSWU2drn8BY3bxGjDiORKbaQDq3GbpuIOTvD0EIdRv
Yf62LB77UqT3bPEzQ6jUwZ3wnn66JCvf0f5YFilZqEWHMMT85dIl0fXq6cgTUmvZzh020u7vVmPp
RhB8Y0klrPeFPEK8oyFTecfVMj0hWpAidWI3fqkg2iRPVFdpHnxDMTkYuc5e5lOWGE5EtciZMs8f
J0OYCfCvLmoKUrXv1qMZvIg7hjBzACviLqDDyHkrDDrBAfH4wtyChfMOJGPLk+GObLMS3Lp8Xe1I
NW9KYPMdazP88X0G+quqThVn5GBgZA6CqyU5sRrloufys1iNFdA8MnhBgNQEfrC/9v4UDe/bLeID
UFqNAjfLSNv6mnx+itaDJZi+jVLSsLJOiZ+J5aMwSpILy3Ie5AHPxY4f6unq0eV9Fl7+p5De3Zs0
0fNb8KY5rJhp2odZs6XoxnR8Voo8hoxiR/3L7IJUPkxnehI7oJ8C2oX8DnuirPbQc2UTvZHiYZjR
h4/h9nnthBEhVSLPQ8Z7EFh9n0yDNZcE7M2k+wKzDUQaHlhU9xOYMBIkspXCnaO165AGNAeZ24xi
uvPRoDL2cdvUe3n4cHT0Kvd6vTv47i0TGWRUOx/2N+kRNitGRJOeOQ5b0IgyHAwc4Qr1mEVh7P8K
mZXUta07bWbXcVL0V8oz7vSbeNUKEN/0fWzmsmONbSlESlOMKYDL6O1M/T9SqAyEcjxnFF1F0DM+
FJMgQ05PVLM/tJ6TgDC0zpsRRUYLL5onDBFTuS/FrvmNh3MnvNHtEyWXy39/vA46km90v3ZDDBPQ
XMcSklSU6sb9/9wN9gheFIR+ax9CNGJviF8Kqpcn5+1pQiJiEhDJjjlqC1rQ5EjO+X8R1hswYvHJ
g2/0/VFz+we5LyFclkTsmUhCdPu6USXRGzXqf5w3wDqHIE4EitM6MINE04CjrNrJhvGPsyy3o2zv
1ZfZYT5I5spSZ4yvkWihk8KaNHJ4m3hTaBDlDhKI2uQqNwIIy1vxRdUkOah6x5/Jwm3FhO92bGAt
mntf9rzFgfs2NsQcCN/HvJRvm0Dg2zETz9FlCAAhqOWoyLzR1feAHZckRNy30icOhvrR8oscppQC
kj7x0xSMItP/Ptfmy4HZMqjgj71TIRdo0qlQu/81HGLwbuLSZKzWshNupUUylQQcfHj9+uzzmcFW
oBWuQqwzeAgJPGAatbF3bA834csWFNLC3oUoC2ws4U4b+dxjZyJYAR5iDzqA7DVJBvxSHNXzojH1
YgPd0DNVWhbsxrDaHH4jXmyqDmzXO6+yRMbdJ4bl+WOOc5xwrs6rt2BnVs2nEL2ZsXir/ruLFiBu
Rkdzk8Qsc0wX25DTAeT3sEAVRhK8iJMkuqQ9OPo5g2epFqo+nXsKLOWG/YWNJzAZE8FNVuWikoWY
Bx0Fhz/KovXM/EX9/B2iu9AKY0fjBcFIJ8rVS4Kj7d9ZjgaPsqXoULmqp7uzJGQd+c81YAWT/B/q
9Pm2ByO+QhZ+Pi74GenoYvhbk1ce8hd2yNsvrkQCtxDlPCihto845zHTHQ+0gLDrAEtqnEYh8QtB
e8g4suFLzTXMeRlu0Y+7hChHnhLTB53fhlBX2V0sRRCcHYypO644RX1ouU7kiIsTGseSKfrncJPA
Ql/7z7HDKAH+3ro+r0r2Fdp7dtqrie1WXzOA5D+oXFt2clWXU+6G+YugtC0g9f99H4paUVPQfkl9
hFFDulrRrtqASGkHsJf45dbH8MJ6dyHrq36prRLNxF8zsYpTHrGlpgHcT/sicLcK6QTHwWFAAZsr
4lAaE6V2VlC4zSA2n/IMxuBptZT06NJia7SJNlo3tInOnww/a+ZIw0wR8yoHsz2A6UPMUAqusJM0
EWOsd04k1c/8ci5AqHvIPIX8MzYYhn+tFQz52991LOD4W1Rfs0g0m/ZoVCxmSRK55uoAgx5m6p9q
hAm6SbDvFyAExc4dWYra+VxUmZTiy2g53TIX7vKQLTod/BSQTV34CpESM+ItsuSVgj/fA/YrAknw
YwoddU2B+VgBEbxiS+Ws0EQdNLyKEIVLaWTMCubcvZ+QtPVNs/7AT3URbGGJEQNofGuavW4GAqGy
RAttneFhNM0mODq0rvDQjlnBzWoKCBjfRAZRrt2u9dWlbHOz1Ct4by25qQc4BwL98XFkBsBFJ1Zt
+AlQJ1p/W8I7Zl5baGk9/84F1JRIiLvazNrzoPFiMRYw66NKkNbaU7Zuk9SHD7YqSzHTSI5MX4lc
quuQDpZXuDYAUBnC31rF1GCETOXY6cmhBtnnIbWsTNjCkxx2qlmDiME8T1Y/ovWhLoskQOA50WIm
v1/j3LRl46cmFDIDZAYWTzZBnf4ond4a9TXPtv5ssIIZaQvRRT1+oid0T/WXzMulzKCUOViHzGwL
upYMaHFV+As7Ga6zzpQSt734GZm2YYrwclkjBd0QiEHetPJaVPF8VCdSUqmdkdMOb8Psov3rDLgL
V6iLyi4fh930/oKvbSYT6ZR65k95bzApdH40lA7n6pLIdIFiRNaO5MazG/f2+x6fKFEnxzcdcLgA
4WbW1TjoV695V3IsdqzDpPhQK/CmNa7oCmj+oKu3WvqSIiIaKlDGLSC0KUc5E+XVuXGVKBI65fsW
rvxIPNnx4iPx1eIr45GVbDkYIsj7SQL0NFoyTG9dTaPQyFuOdLdG2MEPS5Z7fevTnitECgtdVpOQ
Me38Ps14R3zz6wRKfwtCDYjDnWlGEmQUBjAR+17iv8Zu6mtfCM078vsuWd/LXCqlHRcMJi+TLCnx
BHFPEDthRFtuoxVrnpfwLFqEQCY2qsOq86Yu/mEEXlor8jFqWtixz0k/6hD36YKjclEQ/XEnfwO4
mYvefboBkkSQTcWPF8f4T7AbXqZleDhYoWANXC0NIYOhSjFKGizLr1tPpKR/+DOH6oBKsMBQR1+k
XCUvxsTTm2HnOTmVXgYbxigSrJJgHMf2BLBV0QIYe3ga6Z7KAIXCATonBfTd0lWWwbGsCQ16QF+k
KfM37ZBDk/eYBcxy0nyA+v6IEnysENlY42lLNiQi9gms/6QtIx6wFmqkffBgnTyGTIPO4pjV+eQd
SOQMF1UZWBdJtN5mi5Qa/kV2tGjjQ+88HxM7gnfBmzjFjQsAxHth7OgSudx5IUZ6kbpsKYklxJfk
lNeeufnt1oAhGUHnrRvfGc7LSkt5jVTc4qs3gsTz+zmZ7gPpHpTQSwi/1Sv65BN/O2jwHE/7vJGE
XhS44ZvTc5pHq2859oGNOFd2UpVDNApUwIHRxSoWu3VAkCbQUW62EaMRnwn5ua7BObuvqJOgPNRR
+x5yzWjzhIO5d5XHD2CZPi/ZTHaB8jTpBZxVmcdD38U10AvkrWeGAFWJG/qO+2xaJlcZzPZf00CV
SpumM0kGElPq++AADsyeWHuSirlge1hiBWZETF13uzJMCJNemy54yzvivPmEWDHdq7mF242/1nBL
eRD7sBlWaTaYcyUbzL4ttybfSp9zlD3cvdlmx7yja9kQV0YR8ZMM4Fes/bcmc27L2qBB3q92GRZF
ZMUsWERF0FORC1DZyq+2xHbtnxS6rSYsW+kOkae4/kVvX2AQtdlytiDm+2ZRWRTAicu1RIe9SbHo
kG0SXlAQhpG6b8E54wBXhCBvA/HR75bue94DsDxEY1oqLwwqyPbKTA/GBpEPl31CvJJhyW9jsNBm
plawWJ/SDzL0Ic6l/KLoaVO+J395ViCwORKeAOGtk/rB+b2ABYXeOyoiZKg707lOBdSVR3NFZbZR
ZbJ/yWhEQUdfasV/6gg//0XaEydxft9FdrWTvdY6A8Hx3XG8WC1gXMMacT2rx1H5vvVbY92YV7NM
yRn1lt09nLUboBpCQhEY2MEZ4U+VFFzJMVjVSfR9NqzIPK5U7WM/Cs5JBCLrrw+FVD7+ngHYkHVS
u2Um1wsopGyqCsa6Uc4DsX2I6V+Rs03+6r9KT49M83/jBs1BAnEoz9W93eGjZ8E59vF46zSODZO9
7tvkKnbD2S2LFWoR/KaMnwm9wn+RHcD9lkIULfbkfEbCLpRLhgxVSSH8jFVPDXENLfCJ9nG2xHB7
wAzJEbAnwEH+lY7g7ztUaIrkgxk0CSlDLToyZIgf0wP4+u5OEN8nflz6TdNdMoFnfTMSlc0jrxFO
nC3qq/3aXQNIoXB3D1pNvtI8/SMAS+9RQbd1CslFq/ZQPxs0eYrN0Ay0E1nzTaO8We6v0h7ZJDCY
h6Mg38+quDKXemTG7eSgD4T4ATyoqcdk3miAxwqYJSiYqk+2J0IXgphgMciZJ7OwP9n34k5pyZQk
vSpOBY0VYwt6TRqau5NXvN/xMdr682tURIddkMOTS1kFMQXhU5bArVnVPbgwh+2lZPbAZgifhWg0
qP4WagAiRFZslB2u22ztuL4JxOfPzoztnSAYwcN0k2dl6ymyCbPVVjX4vPNh9xL3dfwVU4BfcD/i
8tfuT/SIRn+E2WkHHRepcmYxQBJHx16aElvr/OKdfiitKBXSreFR3AGhTnu9Zx5oO25nm/kpPY7G
kJeHd1WOrZNqOpPvtZGnpuoSllUqKjv6BR8rIChe+G++YS+BADEUqCE83//Xgmskn8K6m1Oevpkd
A5tN22XzTR48rUK6DYc3k5Q/RP2lIedDPq7hhxuHyTCxb477G+iHIypAJjlgahvXgKmj3KjvzDqF
prnWGRGPUHV+yp8LTtHE6FRWR0g7KADv7KZYyFbr6wbWBl7aRTUlw+b+rz7E5N69afgRwcMmBvvf
9NstEeS8lwEMMIwyO3ffeh4dkaXSW08GIYlwWr/d0FewFsC5h0gEp6x1hlkVw0PUiAMOnYxbNvOQ
mYaQMO5kGJHLwLbQmZAoRzyG0vctZTaPiR8CnyWqrqHgkg9kecD6ppZImE5rNhF84/Mm/UdgBcjL
f34FGoyGowbUdItScXQDdH55Ac+7axzSgk6G/zrqQz63yLKGQa0eloCOteqppnJhXUM2UtQZwD7d
qJEdpof2vAssdX/IaEZ9LL1aZgg6KIJvrNDcNvy0pYHnzzWXxJUSHa7Azl56KJHDIOZnKWKer6zQ
HDM4gfeQRnVovpmix+/kaY50pIrTHnKj8se+YYyuoUnWibFREXRWeurTxYiutHCyQ9z4KLGE7l/0
lJVHwnqJEXSny6D7LtTEUrtuIjE3WatI3nYk15MT62BdDbklap+Yy9+Q4BN2/VFHRLARTrINaDes
1aeQf85EioAVFjvpfiDIeldE2ZlUvsUz3m9qZmAufS5MDrqAJlqBLtzTdlGizE0Vd3k0kBiKMBjf
iGk/N0qv+/t556OYjeq3qm+j2cCQ9vNo1qJ4B8xcvsqqbDHHzySehDD6CMrzjmC5ZSynVoXZxOh4
Oj5ng5ZtBcaLVouRk/y0J2C1MavY/YYWR73pOPoC6rpu32ylw9dn7iwsT5DSYb8rlL/pvGdr1z1s
nihtBMStITomrASR/thAuV3bZihkLN6pokwf/MpaVbkx7ioYfVH8rsGxKY2Xltwwf/XG7vPasfSp
T3MfkAqWofnycFv8whQNVrpOj1Vpuzc6mU5u9C+RfjRNccdCiN0r0Vb413P3FLSr0dt/tuyafoN0
RbgsDhm3ZemBSOmPcLUn3SlctEUXkHW56xjoejPsD83EK/BZdyQCPxqygBWioP1XuRvAI/sOEW0o
lSTBQ6EaNUGkewOq/yMm8A4ZgKVGJ8sxv+H1fzJDcqYB8gCs7IbzOeKtKY6neIdXjkHkD9M1YOqj
PEXat7/leZXtfrhoC5Xtu1oY2VVmOwskOx3DTcg6gO/htOEqrTTIxnIOaMKy6/72wmxBiq8xuJmI
2xV5YPUJzNn3AW4ak8GVaCgb6mGRyYYBxn+/xFG0yjfMeQQDr8hy5xo5K5mBh4K9qqsmGmuD67OR
5m9j8a0fbkHiNlNzLp1BI4ZvXIaTr5T46c7o3xJcrnp1EpxOhPwkyO4MO5OVFJxQXqxTD2QheUsH
LNZHeUgnHcCWn6OgkvgR3d8g3ETGnFEoqdVy4R1KFHl78lJOra8We0M7wTG2Es01VcfXZ/AHl/7y
Jkl+LuHLsdpGE5IvTT0yFQdElr0uI/pqh6yuRHP/bX3oloHqH3RXpFMFU0E20QYJj2tPWajLRICt
GYC2bcjknsIh6scWNSUfctXE8YKrKz8KdkGELLPT3NFNsdlc+GhX1L2bHAM+S8JUwzqNw+K6WMel
TELaByV2jNd0Js7x6+dJRSl96fV58/NjzkAoS6Ksvjr4RkcjKsxgUZQkmE9wO01YE/nbFxt4reWb
YaY6RpB1Y8TesF58KMI9mZCEzVs94mOtrFZaWiaFzwLYekhgO1V42b+Xk73VfAzpVmEywzdE8McF
sZAfRHRoF5YtLQHU0vd8d9kqbKPB9ZFc/haJP9EStWHy2g35fa/uNM2YhN4KP5Zvh7S0ldHXKx2h
WG3NdJuuwE2iJ/hirj4tjTAUtBIukvncRCVOHH781vQwpsvMsItCcy1ryrrUGefXcESlOtGYxxsm
6CH8nuL9vePsI0SR5G6gqtH67o4yiXQYK9xtJ/VVvr64qoKXPgIsznHvQfhaU7HOMReLAi/fJW/Q
7q029gBVgh3PkE1iPUlwRUoBb1mXYulA3TCUxco2x9ReW9Zan/d1ppaposYqk+SpCmPL/kDQ8Y+h
wRPZC69kODWvV3YTNtE5xJNRJJrSZ0JIe1v5Xg/vroaXwYa9Fo+bG6ZMVG9HW/ytHnpPaJuJrg5k
RdRZEjOho1OcQD1ILZ1O2ACCMI+/4z+VYugniBQBpud0ijH9UG5kqOdRpSk/G+Eqdta7+Z2wKeoA
1Rf89M5cZQii7QSQBcTl6PZU+tMN4ksKbsE2M57tw67F19vaReKQnSev+6YmQWUxA2g+/YxV+YmV
Hwrhtwdb8pp/JVSnnMwsZ85VNhu63EF8TrwLeAbf9DUekkuiMqp3trGSoUfGDNyj3aJvlpIX+Vks
BrsqTZ/bm7cy9/X1+cb5N0PHHn3OPqb3z3akoqmof51t8dkFDre4q1h2j0VX1G7yuNKddxiUzZte
tSY1W7Ht5Tx2NjIgo1KVSnYhk/stCeJDexrlYTerCFhrvrY+UmWdIBVfdwm5sLz5GQWZR0zytbsU
2x3kzvczyy/JZUWGjbr2FVYbNp4X4PjQ1sXkCLxGDVrfuC58R/ZZahK5SQTP2+8l2dnrqS9PEkWL
FI3jCdzJcSDm2kOy9JwrjMNXOwoJRj5JemTbarZiip2ac9hAPZFhFdEd8W6ZRH381ttiVe3PzcyP
7H6YbPAVlgqqYd4BcHw71GLE3RkpJYYAg55MqB5EWrfDyFsssSQSTWCkbrYEWY0/yZ/RHqZOClbY
vwoKrk0J9gDAi6o2Tg8k4AsU2u03+f/dva1ZU3iJtGjxzkMta/74ZPvVOhwg6Lx4iTQOVatruAFO
baB++wsWWmbjDUdWm6FJUiacE1awX25iDc3O4bcGdFAbxBf03vgredVIxdkM5SzRiiLuja1wW3lO
NSvCVqP6Jy/tGlCzQ6AAeVAquB6yhF24883bytQd1HPYHoU1d0IO+ZmhEqUL+BAs5rnynglozE1W
ppdobQC/3rMJqgljMdpbQgfiI4BAGvFfo2UIATgRa8EDW53TGTYDnlpODMQPvcfKtKIRB9KubU+I
nuW1lWLpbetTEPjgJooq8/ZiYbD0+FenEnFkN+4tZC9x2gvUVfwYLdNibaTXdfL8qvzfYiWkXOjV
hbZWz23oSvfNCFjKO5ezOoby+/MNFzdB4YAh+HX1O1QSLVi767t07zSU35Ry52rFP1uh2R0/hkRW
zoUre4KyDrKhHphi+fzYOoGOeClebftFFNw59a961hidcp0Y6U3PN0ImIRjmZFU88/o4EbYDLs5n
UUvNMGxIOPLDsSwwMQoPlzxAuP39NT/9vwd0WH03pFt+sKu6htLsx19OQpLVVwge0Q6nEAuJ4a4B
OWZ4gEjRGqoFqYeNS0hzwmaS/WkKk3fSQAFYwMTP97nZ0R9SKwHGDhI5rFwHLsn2BTKYzg0cpjxk
iBEPvTHOhWYT5l9w7aRJgpOc1aBnnrFn5LKmkNYfx6qTkhcLu9GMMJ/Ir5cEBQ+4IuZld/ZwuTvr
TX1AD66ALRKsgHAIFSdo66sAuD2RyeP0iU6csb7cKZTIUIzaRzrMZ/q4RqUY2PzOE5+GIWWAZdp+
oxqVXu1y+P+jiYQ2RYpudTFb566NEZs1HlO0qAIEzWRgwq7TABgGtOPhlM3aX/WYapTZLPC6iIAJ
wOzMHPJE9ZAo7TJvZb+BCSQ5dVXqAssdZ9tfVLG+0zcECfFEi0+2UDHHv4VUZ0JTH9StPdcAGhwW
Y85rS9q3Cc38WiglLA76KFioeOjIXtT9+eyjy7o/Pk2R4T0D8xgYwYecVHC9VYuXaeA+56qDLnGC
IfOtYEw0iLlxSJgDVINdJ/wMsxNAvliTYxYrMCR8Dgd5JDhWM/5U5iOMGMWs8fbB83KJmqfdPEMO
HQGmyUMyjQ9hyQ9KwZmqWbKx+wEnD9qyokTV9hUDMNSvywXwUAkHcXXyavVNZmEM2w3aCE+UHVdy
7jeL8Jafcw1Vdo27VjQSh+AV8FZWy98aFGJPlt2jK5F3BExIgBA0sj2lqKEDSzcLZYTPXrNz0aRh
h4Z8/hmjhAUXS930HtRasFlt0M/2oRcbwk0Rxp9OShQOcO57Io4Kvv6FiDArY3CLVRePtRo7svLW
ABRBIA7JAMppqGYUquREU2jI943ngXgXuW5ijQSOZbLdmPvNghibiGI0tpuF0P8YtAnbl/tDzI6j
HPmC7oYg6vcxZY26P9bxUDlJ25lO1tU7y9UamM9KAEIcLb1Qj+pYP6Abt2waUtSgt7Z0+nOVyDJS
zg964zrIdwi0Aqzx7M+W5zqhTqC9UZuKGbYTnNo5NlYNXdC+uy+zP6q01gV9IErEujouV+xQ5I7a
d+2thg/M0DkTgEBGyMEdCjOeGqddV9whKT7BG3dW0V2VzhbczpxJ1Y9dkABZjzXJSZhZRitjrb3W
SoOL5pEdl+ZaCqyAdg1vCgo4PFH86TqjHHBkv0ITPc+2zICQIZD7hHZ6d7s1GcXu1mzoxq1ExPZU
IMPY+QQT8qPn0VegKObOxZEBQ/lZRRjwU4E8Rciz0bMYkPm/osRehAKA7Ubl50TwEgqK6sYmKd95
+zrASnqA+lTCKWrLUw4l1Y6/EENZ2DZ/LoP0qJfXYdFkSdn66PwXEhyw71YJS5lM2Tmn0qhzSqi3
Fw5iESc2QiEzgQGsH5v7A4YIt0wNUPytQAUU/dfhdR0H/odW6FfgTgqKh5bS2HB6gVzo3gYw8YOi
vKPXHcnXCBXa4OoIRygh+1PDIon0pbaCnHoRVUGC92vgkR0ytZp3OsDgwUJtDUHPPl2EvBfpoRri
XWZsQSBf0jxibE3ogfmkpj1Qb8lMD4AEl18y5cucOPDCUc76Sukx5VPZRk89BpeeD0UQj2GWPpSP
JYk4Lc5Uu5yuj4F4RanBLmMmY58X6d/nA6Fy6jopd8tYyXMcBDo7usJUR+xqnYijm/Gb8ZlBrE5W
3kKJBGU3yYjzZmzlgHERXzO1vNnUj9MYeKyTiQm8MyOX22CgIz6WOSlaVmQ4vAusuXQ/Qh5tqczJ
gcX7noN8IflrXxm7UmSDkupfTd5Y6idaoae3rK4+Gg56t3Dey5d64cDfG3z+6kOvXRi0t/SnF0j7
E7nbv7FbL4UKP+qDfEdIxXTTff0mKNpbbT9eCKNwqYJPOZEFh506dU0kR84MZuLjG8K4j3UIttBy
E2MqcFLQdG1y8Dr2UHTPI3po8rLDiH63qrKIe0dcdTNHD3HHPMo5jWCXafZ0zFhUZHy9FXlMYpMS
uoUgv7Qb0jDbfydBtzUq/Ivdk0M0GXYHYmiT/CRuCFuOCWMyr0EqF6M3AeF9AP5qdnqyAxq0Deem
Jr6uAdTXMrnihvKfBQ5RHa5mRkOkluh1n7fm7oLFPlntB6jHJGm3gLtI4vyB+GuIYiqTq1y6jWeo
Yke/GqYKSUyNzzPMNQqIcP/hCgEJ11nGC6LAFA70gjpz6XizfUo4qOARQji57v+fracj/t92bSMJ
5iLcGNIRMYBHemdE8z5sWdY3gxTASj1hhmkc1pVU+PwBJ+0gbYIC8stt2uYPpifYEhLGjcl7RKPE
4TKvX/37OvIvPy3521J474mU13474KEzs5ZVPZM7JG3xbnPlfr9P/5Vw0vKugJIJzEC184BnRpl3
6614CF20NNLMO/3uheSqh4DgxdopzVz0xz2IK6osjwL7zs5g6DuZhVvPydPPblIKZ3siYYQhJ3VS
ZmLvtyPjP/lj2NjrR0zlWVU8qk6GsZXEQbi25hIEHW6kW0aHy+2JJixYEmiT3VbMbdag0SkK4C8+
Rf828bYHiCU4IjLcJk18AQluWHo7sEndZX43Cc8Oka1QBKXFUB49F6ti3uBs7c+xcmC4nv4Nn5/b
qJToDxHecA5mdhFYFgZUX5UsSQ6VnpEhXIrEb1nnr04kN3mxHRfpBR72aNuaizawU66wABp8I3H6
IXs88jAEMlRWPegG548/AYdPOFL6B2eFppGcrepd+9IeRMkC/h11zmTXGveiZT61yb2yNNR27kie
RQaDbxdufOP00JzRaR9pQdy8EhG5nY/fxi5VFlUAxoyOoSJh2otTDUanatzl06YUFvz8+Gy9B6Yw
OkfJxv6CMCSx9wo/ouK7KxmboE1svbZowf7uAJUu1NslrbA4EXxpJ6mAJExt7Jh6A1nCRnjrA7dU
ayVnuP/IGG8IBzSMzJzI7yFGPcBcZs/mpPt70iFErZtWdFLKTjbplg0URrFEnwIOiu2cMHtH9Qfi
0zz1o/gk3sIz42c7xaVRIFWpiQklyHZUThla8U6U9XS1uGd5cftGIaWCS1ZBoaurUQWo5jKucrzC
wKkh33/DsdKr4sdOBtVA7OUaKVni6EMXMdwaJypqGF4TaDfUH12Z1CH4ketTp39p/l+eRWpHG76F
ZWnBCB1vkdFyd1w79e0g4MhMxIKFlyFb4LjeO8qysNk6Zlmwe1/krDpJAToVIjmsbqOqyEpInIpz
zgCwZTX8gS0W/24bsoeYKXrzfx6uL/MldwS4DldXXo724szzG8jB60xUx1utw6X8g9j9AQIg8GHe
OnpUiR1WbvfTDP3hjPtC+Q3lh7tl4VPavISVchDWQderRMyEp6G1NjoSun64OYpLz0qpI81S5si3
r3Wo7Lhc5OWDrWgDfWJrnKH3J3PbgGBN2cYFQYrl+GedpMB2giIVxvnXzrtob1PjizUln+0EcAKv
80zaMKFEQvT1jrRCbAukC6ICFqxTINzt/EZl3V/AKPh/T8jkbBZfZyW+Q5kkRQ0cWU57t/Vni3xN
j+z8qIqo1ep3qj7mZIIyqK2fEFHMx18YJDStnnP85APYIRIF2/gOQl8sQH/BcrCE5hSBBQRGY+5b
hzrqJyt3RqC07k0HNWKo9RdnzLtRcVAV9zdY65M96XG/Gj9nUZudYSdmKqlDfrMom2LsZGfrG82o
FNHX36uQTfFfspxEB27LW8nvzCGvcHFd082pDvkBd8/RsjM1RcII05OkbVf/7KUSjykkGmmXNZES
wu3e6/ki+Az/6y0rmVusJjkpIJPg60I63+nifjjyw/W26+Dkl2xydKJou+hFtUdw63dhLnDE1F+b
XqRAkgJT6YSZVPQocBKxdhOHpvIht/4Dqh1qfbpbJcku5JCfO7V29m7lQK+Ajn8RnuwERp0xQBsz
eePX9iLhg+U4hw7xM+gEo1BIidVbRDy1shGgjmm3Ofmq4xUH6/yZb6ZPrMbNmjf8fjwkRFNme9VA
rRaRE2z90AAlKdK6/dFxCvjenZzZXWeyXLjkrYI73VN6xp9ZNUE01A1kaEf4BoYum2RQQvXgJQdN
TEgpgF0P3at2bxKyR5sCmI4xn9ByyURQ5gIsOrbOeJUCnjTzli59Blr/l2WGSgJC0vScutlX8GiM
3QFxt/Hyb7Ug6TVEdGgKSDcRig7B863DUY8bq1BgpgaM3C9eTB2HQyL1a5R6NOAnaLQ2f8cdqswi
43rvdfMcc0ddAtQ6Kdz/sCTlfIcybRVDGSwXthNGk8LCKN0HMOvja0+Ky7EEUJbrWv0i0zwbgce1
T3/EuU4xR3m1479p3d7Zo6sKdAvOR7sg6XenBOMqMHGTAi+K5JQAq9CgA1fP9L2PmsG2mDuwsby7
1yhysJMbIEoyqFkBHjzXjKLTzMQbOb5rXnW1a5SoVln/bPOpdGLLQlvQYSBT5Sn6PNSFa//smZI9
tGejaafXR+7n2lqmwb5f3e4R+9Xj1vdkW/1FR1FILIrY7XNL5qbLOWJ2EWUc63mUbW+7s8NKb5Cc
354MilDIXkEDL563FEuXgrPqqAJr7zZ9hRCa/EYPuQIXsAw8bXBDsGqtQ96lcRJA8D1L+F4zJRT2
vTjAmc0Zx9dVThAo+MvDpC+w3ofdejHMu0BM/Eew/My2pAWKpZTJCWY0KPgp2iD6MDXwzsX++Dm6
r2Eqz/zO2+42dSQxQ+lX1GHczGPYX/yFLZWgE16nbqUpEF7ifAQ6UsnYO6HwIdSe1HpjWjSQVVDi
Q0g6OrYq6LIVb+8z7q6UwbH0LtIznccbtMbDMKZkkTA5g/TGgXUqYEq8eJWIhDI9yspCzdCt41Qd
HGV/caWHLzE36IWdMn2Xt9Ty5nTOk935bj1eIhd8omRv7G2bgnLinfOF5M7I2sotGwoRO9NmjzQI
huMXH0FzLxxkD75PHl2yXKTjOATqMxWTsgCA/jAx+H00UwyvtWYQNokxB+i2KXDH+1+fo2G5Y55G
TVZFqyWSdkHBUu0c050K3zpkvNm6g3Amj0T+NeJGISCQhEv+or7tAj1UVoNak0Q8ffVHxy+gmxkM
2QBmqH5NQyS2J1NFy5Ycob8xydM6yJ9/ltEvkoE8VDS67a7f1KlDyG+YJc5sGgoS3ZirG8q8NNR3
IO2+2EIVGmw/KgsGO0Zg08et9RtCBjqIJ9FEHAd30aHAnCPEENnbQvpomISOT/F+/rZ9U/t3F1Ds
9vWKl46QdBcfkdrKADp+azfI3W4EapHfCeL0SH5v52Kza5Az71WFmPsrU6zvZ7mBqfw9tgu256z+
HZaCd1k2BkWbf9QUGTAJI6LPBJ5+VCkIvB+IFhqpMJ+SKfGrcWUak8E2aFkcjyHExekoXWkTM7xZ
DCOvSAaH1+Vd38N9+DFEJw0z8vccL5EqG83AePo+Hf2p6DwARqJGtQZ32tmj/jlRhU+SeNYMyJK4
QV+THBD2PzzTL/56RkBLczGoLQVHA6u5vDiZRIlGCHJJrOZVAPwFVG9f1BAqss9pidFEUz6o4Udq
UgpYwwqAsr10UKCd7qA+vxvb4uaHAhXuczuG1gQtv717V9jAXLpJR2Qwd4RrfvKHjTEbISkFBVWr
wOXmRX0ntrXlF3USc1BnHFf0tQcSxM1WZqOLyGPSAMUTYOKAwrZepZomNY0ZNfsyN1HgAAdPbuIU
BsD7YmCuEkWbNBFf5/9tgKUEWf2j3eiRZtuk5MaXqwVVgtm2E6XOqV/tvNsd2feaNSkDtDBSfvnH
q7Upnuw0lj9noixkXcWuB4gYjr7q3DoZ4OEcwOSf3CwSZ7chegJ84kqEX8v/r01qz6IiqcqHPpEu
N585Qu0BTWO9yTJpXQYpp7eBkF9o1bQ4Hx2mXb/v5saN86r9Vwfx3XD1OU3A8tMHeHMPmOPofUYg
vMjxd8LaH84sArZBpw814tQetJcsyYnkLW9Uxxr2LnGXBNZeA+y8xpc06UN4qtN3MkSc2R4IZMTb
q5dQLmGrws989h8BfTvzPiTUFsZ1KKMH7gfFlA9e/iNXUImxHCCtQJn/6KIVw2axzcB5nD9qqUb/
f87jUacihujhKqhbLPnkiwgk44CrTXbcNxRQ3YPREN+su3U1vYaWIgELoPtc9pbRMr47jlpaX7LN
qF70LosQE5GujNRC2k8TgxlyVyLsTVXCP/moyMAYSHfYoMUMXb8T9sBVoyXn+mfXLxD0Bzr8kyT7
sXwGAOZJs77fG4c9/HpGhbKqxpIybjBd2RMy4fv6egYJ8vGimabKSm+Y20grlX/SiHZiD6or93ta
fqgHMEliDelGE6M66wqnD//AvAyp2KrEG+f4uwivDMOrpu55F/foWIYCoA8juX9nU5VnSldvgj+0
YvE0tVNxKk90YwaJKrfwZ/n9FFvm4yTmYwBk7RlgiT8XDjL2QsG4CxHAywkUsS/wpg7x79xhPe8R
np0ERaBg1g+mQrXUZifh1yd//nvDHOHVUR3cG4VVNyyLwoiz0TdCDLrfY/W3+G8O8QtudVFm3ISE
ThwqSWyZHzhNgcrxhL0yvT0streesun71GT1L6j8Zx1RFa+EoJeuVOlxQJ3jyMcZqCoP2MpeX5gy
955KtchIFaYswFyxR2ZWFVBu6CRyeAUlJeYAKmz67s4P9VNY3gP3Z3snO/g9XN2uUJyZ5+1+8P/s
x37jvICTNpyqdMNn2UedvxQ9Juz8ZlD7HAmbKz4E9PD19E2CQCfQI5jqnzmBQ2jpNQFg2HDAr8mM
yCu5TjX8Hbe25Szykl0xUiNxF2gwJelUpA4W4lAkBEcb8zRJOkrdtHLVvSOFW5eS3e5+3WmuO2GP
PyCQ8vgwiUF7fPls71oO1IVxw9vm8sKTeomu+53FzEeFVPqGpvpHTLD77rs/4GvVMWHVaP6N4g4H
flqQcnT4H8G4M7gQVPDL5FxRZbZ7IrgdQrcx6ERosLg5zVOpJ0R2j0OGx8TaSiDCutLbRMiUpnLI
MMgTTa2X+OTJ8X3C7QwsF+pEHdAXlFabXLWFZBYvB2Q8Lz5aiawPMGQ7Lh3NP0jyY5E7JnbIdWAj
QzdtQ1U21+5Xk5ZMVfYGVJVDiBw4Jwf8NVQ0m57Cx7Jus85+Igt2p942yerd3HkYmh1/k3/NO8Ji
YWuDvOmWYiWE1/+D29JjdmlX1op5HFWp5liU0+FObYeWOtyy3Y0dczmiXJjN0Py3dXq5ouvU+ZnY
dc7yvSkYA22TE6oxTQJq0tpD28Re1pBoOu/JNpZ9mXfV3RYpGKh6FI8i9OuIip+7nPmgLIznsjQJ
HeORp2g5KRA5WSqUyPX57OH42MKB93K0jSRlAEx9LM64YSxAjXts3zqduOCQcOcKut9Tms9xY1hL
N03mqgionbYBleA84CAnKYunWmiK9rfSAqlI1CRyEzsDRmCXEVGXURL/QWlSvMta92HZhR51Fp70
VV9Cx/oTesNI+yKvfxhX9mLt6jhXoWvj+dqmIG+cV3rtPLOeltLtGrNUmnaMusYkZC0CGET3DGBB
ewF/cQaiRQ5H0KNqmQLn4KSdbQ7NbbzHPvs1Q4ZFtEEf6j3C/zJ5v5t4VsqrXWBgxcH4tikwT3Hj
BivfYK2BgWKDpC74LW5USwcx3XDRdhXNIx9StwzheEEbOehldRTKWbcAC3Dw2UuGqt4xKPAbaK/s
sEjsQBgH6MSzN3dohEZ8F0bjdkkqRZ2URduO9BKSm/Tm0eVqpZRR5LMey2PqG+kr26uh43Vv7H3V
F5di2U/M9+t+qe94Dcwbjkh8ESHHF8a7euBYxsE8Y0kSuf0OuOEfRPa+9falEy5Qe16ILRr+Uf6Z
nIVlL59zXM2TOYlaPX/wLLUbFwgrwuaa8ZMiYclZy52wZy+ebE3jY9yXfs/owc0EDYnzYdM3xigy
zNQE7fyrDb/hbW/IzhxGXt2lLZVgubII70WOc/4xmwOvqhTt11VcdiV56+O1fkOGiQXFqx7uGQZe
POnw/9KsfEHOnNeaxkHQGI9nSXwi1TtK9yq5bhn6H3rI18HNDGDny5TAQweN7ZE9G0MR+zXAOtAG
b7edveFFLCz3PjW1MTv/SHabdgojGTOPLpDZxMNoPKmwV5IaWBIm4tl6IXzMMeVaWP8TIHi8QA1O
acrD8jks1GgRSv2nA7IJZwk3b0xWtLtcgbIF5FP5WD1vSzo1unr5Vs8GZZekvp4zivcpAkvBQIDg
dknwt3AD8joRiExhX3ASEWnwvCRs/Pm8M5X04BXSAEw5J1AtNZjCC8SlgL4ZP8WajT9umU1d7y+z
z5rG00a6+Zbbu13AKIVLmt1OOizHIyUpSWnjQeP/Heb9VcmBWrWFoQ5jXoOqY7WRKfizlLFeCnLW
XU9KWCCHzmVBRu5vrcyruEIt/4CMuaek97U8u8p3BOnH9k+1FiYaivdPDYlm5sf5spgfKupNovHk
pD8FyPaLtWSbDwNmCVdoOnVHOVW5A/40y4tTLkePFnpCqYJA1Snjb0y4p+AWQcTClE06TPB7aiNT
w2956GxiTknPWFZLLTuQAk1SoaLTTXTBYJhSwmIbfzD/alyrsAlqwgt3KvbHixqB+P7bB+fusPBO
5zfSiC/SdelwSRRAIVTGBoRkJDXS1wDWlmlQg9oEK+TI1iKbiC0FaDVA6fb0vMBVBerKsiijmElV
nrE9dHqjxc2BYueVETvIANdbL449uZ6IhYHRiNLlGSYMs9A0gKFBgDUfX1Gp2i/JmU8sRRwYHRcq
7You8W44WwuP2pF6mb1AQaXZ37i6m7MNCbSV35TVkqrRR3iDoH1ugVnzv+wgMRGApb+WwjDBxRmu
9mZt0BPA3z6eRMLCNAUOkCG9IrGoQ9y0WKUQhbeyaEPFQWXMzr05B+OD3Wm2LThnPiIupmh3+Sg4
JFnpTZGAH4Cpl10e7zXpTN491uqABSq5/Eec6fvFL5JaZf3qpVc6YkYCZ5uSR3ZYvu3dt6kjk2G1
FfZ9TWYHV8CGts5US6w1ypNoqb4A83wO/CpbmfSGFvg/HBDylcObtaAnxj9j1twB2TJkvusrOmW7
XdDLd9FYls8aM0Ys5qGSho1Wq40szB/JgKfzdSS+4u5J4CV6vMEP9TP2Hzoab9ViNZ1Tr55w22QK
Q5Al7t29GC+cQy1w7hBAQSbHdGkiihAyIoaxaeQu/PVNuw77vx/kHhN4Bwth1NjT9b7a3Yo477kF
0viyFVBAen8ezc8554P1l/m40Z/sElJG0hJJe9rwoRPFge+Nz98jPPurCYHlWoMdUjIAWUzG/+dF
SUsqGbZ8SURF5afZaye6cdGuIgL+GOlnuDsyJXnnAsxa4GTcBBzRkBMTLGkcSAPM2OSeJmqtJMOQ
s9ebSKYJc1K2c73WW2A3rTtNYjzEVLaEJZTmknz7Qhzw9aDKazPdbjksWcb1EbcfJdr0NgXlAdox
Ad3ax5Q0DFAADY4GF4WYHGpcle7fZGK5sw+QI9BNK2mY4KxSXXM78ljk1Ehw7VcgMfcWUf1rxtvC
s3tzmJtlG6sKuXKFaVKCxEqf1vfB3OX9lVF/kOTnXwtgZ3oySB26kwTjF/KboWx4OtkQ0JxehiuC
FTq5NR9QNaMY2UB1nOfEUdF9E5r8FhVzCLNhhBz13P74te9iBVY6pMntwwv2FUCfER9I1oWMh39f
xiFTEU4JrNnZMqbE/K+LQk1twjAyv/XLoL/tq8h2uIrdtyXWqam7Hk4+N7poo9Ui63ko8z1z1a/k
7h0MJd3EbZAw3C6QGQjG3bpEioH4L5KgjmmCBy+BR84qQf48s2bo1/l13/KjD+dx9IQ8n6BWhLIQ
O6+qZ77D0URrDMiwzeCkMDPIwi3LAEIs3UffrHKE0i0xtW/insLZNXII1KZHTqg47qM3Rrm5Vp4D
k8Hfne3l7ppu/FRzy/A7oRJ1s2HegFpcyaGTyi4OJ9bf69so/9nOB0bxwdjmAaIe7vOWZV3Q85H2
M0hHYBzf7L29VTHB4sXHOjHIroGdhRRToSqQ4SgNkLMBqmqqMNQT/HMjYvQegofKLmhvitRbkPBi
pKJini9pPyMZcTReYjN/g5vrMXCj57SHzV8kltTN7M+GsXIojN/rpBIc1ZKsqSciIHOUNowM1oZt
JRMBkAoYAH5O0PCgyLalN94FfkPVBbUtEdjYIEk909OPlFTIyhzGYVGKCgveG03sPg/o3yw24a/H
jOGPJBEo4kLPp9mOTx2t2UwtUn7c4u9tKgZM4HVRV1MawczQl4LMaXJ8y6EZqnDAlJsBKdK952rz
a5a9WEdkXvUBD7Anne21ZuI19VR0s8b2kDlOMzJ4tTpy6MmRGM5SUaz4OUU6c87b+ZkOaveFHqcS
FwSikaNAvUGj+LIIYIqhF+WTA/uJCNMhV3KKrfFH/sUByd/kZ8+T6vkXaHC9itAnSFx9OyfeqJzn
Mw+w88H1xR9mbw7SDKvRuyT/FxvmGZODGqDmwE5mCOZQnuctzem1VDfi3SB4xZlmUKkCNm77Foa2
eOD5zxTuK0fDtNewgMo+jmx2IvVP/1yaf2p1s/lU5vc0u2NvFkIvmKVEoVldberBzsKATsp5leoW
q2sNralkXObolNwiojtO0Wc6LgoOhEZDtIUOj1juG74p0DTg/YLsyQxmYwsajULpriFkwMOW13kQ
yqeIICvxYK8uuvqNGYeR4P4YmhJShZ00e+YZZNSFx4beLWliaU66OOgAEkbIGIY52HozESOyeZjU
r452/cjYVNHqIP7Jzd8773FAnuc0+42rHwAroAmAyj2Nd5xFY6qXUnvpFKe7sIrtsZrq1j3CUu6i
ScnUySyNwD7sZS/atedWNvlK7ySc60sAkmYaO6Eu3fcYiT4AtWQUrKo5QG82b7upTUGYUGzRlAhv
7/PVFK743Q89YxKf6R/GFXqNR6/j/DqjhMCYcKGjmFbNmGgzF52ZsiMJisW8bxctLl+4I9nKOe8t
e8wc1Ylrqiw3/JRnvKJS/NA5ktKEWpcUWcaWl9eGzP7KTkCzGO5y/1wAWJoIWFVsPX4DZzqeXZmF
QbR2vVGtMPNCiCITaKe8a9IQqn1b0DllRTcOtGAu/vu2RVnjDbxKEqxZIxD1xrfhqyCuEit0lgmL
IU5EbnJMLBpciJh24XvlkFGb/U7iY6ePhrdTuKTsw0uLwTIj9KKrddx0jKYGhT7dQ7UxvahgV14a
e6uyV8hYuU0rJWlwYUjP+wTQ5sD85W7YqK9gv29tLcyRyQBcBRimXEz7Fbalqi3D42EURqLe5mbV
PEsjLRPnOYZT9K1TYdJ1alsShRoP1GeuNQCXDoHIKerewN3ZOaBlDhAzZpMRGbPZsqyAgOr2uhxL
SKRMwQgzRWvaieC12PbuSRWdj9UO0F64tqsd94TMdzJ6WTYyropAVE8xYPY4541nIjFi/d9YAPgS
3DGfSYLdF+/tsHWmC5d8FWh/xnLPepyiB+kvuDafUskBBgQKs86rYhgIQoCGrStv1WLdRKDpARVn
GiELCzugw2HY6FN19TZLiT0TG+HfXfoIH/sI9dgGYgu30gActhnSxz3G+iYDfnWcc7KVd8jQhZFV
KZcYmjszQF5OndPP2JkUZa/kuNCacCxrm/WIDwyQsHbnddVq8K8n7UIDwiFwkAACyTDUS5otC41G
AEYx0GcXouweW7ylcTbip818POahVFlxpSjlSm2kPWE85Q7ZVA4ipoQTcw8Arvq2wGIvzQgAYnDx
FL9P47TR2/BH7M0ZcvB+iGMVA1AaxBIiobuMK11926+fZ/WWwkSssY/A6+rICH2eteGuoCaePEki
94SZTB8P+wuMMTHv+HpyiC5VKjY5wTmhvZKgisuTwFIN2H6G9m1vfgVfW6gNm3beEEFxzTnLwcyB
EsyRbwxUAU3vEXRv2F7tXiAhrsaQP0bdG2OAdlhM61+6GQE3bmn+Vog8+XjFKlChqFbwGNRIwgAu
EnIKcx2i8YDogG+UlMKhANHitAa6PIeIFvnimu3E9MKve+74TSWIb9VMw3Cj2QZU4V0NV7zVxzb2
c1pv7YxnPkTWzMX4DI3tizNVMSESG6los6OCq4HLg49afaEjYKmu/2ddlGWfc+7Ct/eVn6xZGrqz
dRVxbSUDPAntcgo+/kKr4rFuuhaJW7VuJZ8zO8GEgqs+qRgITm9Akn11IjXJizXABl8GRd8le1+v
9ii1Sz6i4+5MO/wTkykpwall+xSKszC862tQQgsZgJhCkGGtRIZMjzmCHQBWguN4JJFJIIHe++ty
iUzLjQdkyxwPxCptIllgMOB3zV+J4NtExyqiDF4f6syUDhxmv9JvG0OMENqg/J1NzHZI1gPBBhU1
BN/UCetEm6pV3xgfHysu/PiMsRNuze8LZys02XiBnfoWeeajBFyqOXwkHFrpzQIueOLeEB0kRLmX
ECnUEIWfU1G1bLS0y/W5h6PaEFcPOvAcGy/i9WvbRmsA84V4UeTN7fUoWe2snO7GAtS/MJTrVAHt
4CdhW1U/uXgt4y4I8T+pGh/LEm4ROrL4G324+ovZ3J0iiG/bmepaqdMSG508END6HabFIRUh/DQK
RCpQ3b5tKjXgkgKb/bkJKnLLPM7PwZnJe9UVxykL1cxMLalS588j+2bU4f9QMsrB+MldUgJL6gVA
6g27DOTGMiLDOWoiwDFzEvsr03bEoBsa1FrbHlvVl6PBUFbPT27d2XqhoI80tIEi4+AH8KX3HAEt
cHQBLzVvH2v1j6Y4NABU8g629moFgh5DyojQ+Rce4Yp23809zwnm2QWkS/mHOlJkU3rloOLQ7RVO
VHUeoXTlasp2Cgfx9ADbwLbrc3tDvSA4QiSuv6+sCGdA5Nvj5oDNoSb0PGorGBH+s+cpTrcT453L
ayKqjGsIj8T/mE40ZO1weaVgT/BsjxifTezNzQ5KHPT5cdwnPemsbYuGVK3ybGRDuTpuYPROiQqA
t0msh1nXKdYvUVbMq0xgEDRMY/JabZrQGQkGGanwJo5WjLPoht6zMQs8c2p/v55EM6b/dsYCkn0+
rF56so7k2PjzHFvFjvoviQRXbx6aDSNyQqZ/ZXYdy6OvJPRhEokVg7gKq6F49Fx7ejQiYIRz9KJA
mCN/vryTF6sC2pIB+fQwR4rDUcJq8hVrp352WBghbW6PXy5e9Nrs/oifzn2+Q690fpKlL9TYEBGc
nvB5aXArqxo5GMm13rXzABOjsv/ezOoIb4v82agzJu5rFl6nHvNkjg0Q+Fwmg9whrAumpmFuV9Gp
juNoVJ0HymM60UNf0ytGjmSnTn7Ddq11kF1s8jtUA8+ZTyjgJRWNR8YsIuiACamkwpTu52p+hHFE
L2UdiLZkqvT3sxp9GEdUqBSeRrSbbMbcKJCkPsXJUArDHu40824GUGubbcWYhV33/V/KKec2q9xz
cA8dt30c8hAC1uRzO7r8JLiVfmj9SlgtE11M4SRTavbrTzc/h1WOcyShqes2CxAj5vxRJ+XwoIWJ
Lqy8XslQkRNneXO6PeTgN0do4AL96CcJHaKpWYr6Op7m+zo5BMkhHZSj/VfKf4Yttb7VdbuQZEgQ
cmhhV5y8zEdgV8UZNBI1luszIzxQtxFsrIZH9d8fzluh0mHxS4yGqqKEmIikwDA7F0f6dtp8ynin
EhTphv2aK8jU4P3L+rxChxk5M6EkWYmw43rXf9ZqDViW1mIg5DEWbx21/7gBQKn8CeDdQeuFDR7S
2VoIh7RPDXT+8k8g4x65fQrypINd11WMkkkM+bnW3tLs2T7y/Tm1zCShFEGVxeMAPd+/SCBbnNoe
9bGonPBiU8ZI7OQLDxpOKOY8YNuOrUV+Q3DtUbi7lQS6/WlUX+LNppnx8EynC+NihVDqU4azpdl2
HGaWHl96Z1uAzh3eC2QY5AfCAQrdAMIm+bFugQrvzHLPxMVeWkVfldxvHbJof+ldOG/6z6/ErYno
guBSY6KJm+KfIcq25tFPjUjl0RYYW0TI6dtRUNPGc/tpr1iu+x3HAKM2lH5WkAo4iULavVu1x7JM
ThBHYvt7AMfI+EBt5RyJLpvkzuB2F/X7Vy8oglmesvj+3KmEAP/JK0gwQE0WPMFiJZx3Nla8xKzB
IleT7RYMAZK0ID1NhyA1yf5BkuSHEA3wjpBkKQlbF4Cf/flba87XQIxpoiChpNlujQX+Z4o7JM54
2pRaY4wN/qGg22+Qv7GFycMNgJk9elQLsgyKTjVkqLrXurplYrOn4zuwz6q6NtKc1ySTpLDXNqHU
mG6ZDtMh+JgC/64WVGO+t2Ro4G28hB0fSl1QXz5J3d/uoWwRIqPtLSF1LBm2Px0q/qx3kLXWErif
U8npcGv4ew1VYy+XoLxdIZfyhN/VVM1iJcxxqOh/4fUHzeWHuej/V2xVVJun0Y/QZnYfqFdF/KHy
tZsLIgYA4VRxj97H7C7TBttmi3W7ay8bkDvFJ4DrvdoFDydaqSNGXHj/3c2YNj3voIPpnR9w+hbn
bQze1b9qFJDRG1aU1SMHRTYDhMXc8099PCg1nciUQRal1Erh+MyehWmK+I0Ejv8V642KkcLUYZS7
qzB8CO0aaX+pF3g7blqMOa8CWUb5wAqNaRh7o9Fgxx7A8x0RUxWV9+g8Gxd1QeA3oeKiQSYpKucU
4uL8qUlA3dmRb+P4IQYPmltoWITLg4bnr97RHexOsvsSSMJ+6od3FjD2V95EyKzdl9frh+SqKZJn
gHoojsy/H50Pk9AgGWYOoeA3OVYmoj1E80jqWCheoJGPqxcyafME4LHPJFbOBlEp6EThlUry5Ld2
2NjAzT9ar3h9mfgDTXZM/s78lGvig4DNO1P3VoEXTcgDDwfAIf7t4lj1CWs2J4/62p2ZE+ygLwiW
13l/QfnOwUMUmv53y04PRVs2yOjcWswCQ54V8TtYdHUCfcUelPnfyg6uh7QDY+KDXJDhuVZLiZVT
AbZJQJcFGL39F1MX1E2SajlP/Bz0DzkyQr7u0JKOeMMzcTciLhTQ+Z0BIYCx8f1AY9pVKCWVLlt5
o1hV4GhexaxMLiL+UNxZEHTmiOPq9o7tcArQCAsSpinhCtILh9GbOr/qfGo68skLJa5op74WRdp0
tyJx4YNaZ7y/3k9z4wCsibWa08m/7FNTVp7pDMpZylBhCgLAaw+9bR+GsgTU5bmY9w3xEi8snT0/
pO3IlZLNwGx1dQbb9eVZmutMNpR4Knf3JRBt3+Jv71CAFOk56I0Bm6OdqjUcNFq6OCPAc9XHhG6t
Xtf2EvfWmhx2EiaRU8sdn3dysWFDWeVZBYFU2MHFqbrq1srFBybk6AJjgK2BdyJ8IxsJV4FArRn9
AAFMGG56mKNf88qCOEdRogz0N/p8Lk3M4Y3RRhTidGTFL5hvt152hbFIJBMA5BkxPuCO9/3VjP7Y
E+c9fFioGtc2Cf6OX4UzTPHjDu0zTLnX6e/v1pGf8T2vs+6uT3zNYI1qoAJWz3jEBIM2OEgxd7h2
dyJvX8sqFv2WnJX875Y99svyq0X+a9MF2Kh8QbswsJwpkfOxPNd+deCQQ09Y+3muygWQPPBCVDzL
UMM5SIIxwNHZIQE8Hx7kDfgYjh7aEdz/PSV7z9CRpqTnqdG4NtT5YWkrpwe5O2DwBBZrFHDur1DG
bQ/QcoraLxxtdD4VvLKFY3T231m0NqslffnV2Q7Ek/DUtSJ4tIy8SHRoIk5Igb2dv3GQ3iYuCLB/
Q5tQqsoLuVDEeDHdPaoJ6rNis94qXNCJXwHtwX0JtnrhPxIvhKKuspqImG3nGGGTD386vrr9ZqG8
fKDIfFjQ6y3p/cK4f1pKTiiMsgfNjKufaS9syFXSldDAJXNdCtLxslQils7pgJXSEMdob7Ki4xMv
+21wnJWsXQxN2TYbLzp2ViHtR/JMzIz+WT0YQpCqlyRJA4BrAsMhV9whEOMmis8259UdA1vijHyV
jwrr+kx8fFlAQX9VX1Wd94OrhMGEfSfyRHqExB6Fm9zYddsRtp2I3RlUkjKnLONto7asmVDosCMv
G0hwTPbjZxDeO8SWFpbYiSrECnkN6kG/NyjwHESyeNinmm52yreq+A6AfBsCV/fIxHCLAKf7ubm4
6ABhhWr7AGDo3KO/xmSI9FCUi33Ycxsxooq5Owbv1+LuUbpMeVY0rPaxlbfVsFH14JOVgnszdKpB
cwMZmXQ///Pz2mH/4HThIsSFUDqh4l0Pl5nl23jkFsCxFI6ZXC/c+8X7QDlDk+5DU94hebBgJ+v2
dSV5Sdli6RSTXEXD1Ui1iS/LlvGw56Xk6J5ERuXhTDrs3hpFyCy9PKos0Hm7l8eIoboWLNeQZc+q
igE00TWPuwihOlckrG4p63Vk0bmREolAUak4cicCuYFsY/LU5ENI8psVhvgGPU5YFvxMQ0C02VLK
Tr+FkuyvAdCEGps4wzs1rWCuC4fjaSmx9oRjPo72KHJOjDSWR3PuGtVO77oXcFQ6b+zOsePQl+uZ
c0dPMepL5tZ3v2eMGPuvDDed/Nv7w8pErY8X7GA2sHDoEe/cJaPzHqFk+Nm2kwHhkUeeRuIj1NJd
M+9ftLFAOGgrQ8QVhDMcFdE6i6DxEolwWs1ZLXu8Z32NnYnh68r9DbwaR9KFgE7/9ZM3qLxnJMU1
sB23J5CCVku+4YvB7zEcvtYQM2HbA+mgyu+TF2vCDQwCW/iFwYzdds4sbLb2ggFt0OvUu5izpYyk
69Emzw6/2CAugS23GnPkHS6wJ8zKVDoq9fkFMywiMvpsyb7kW4WIh5t6Y2vMRMeOOI5QOhTNBd0d
t8CvN4q2zxykxkicvvjO42YKBdvMzpvPcynfxbhwM0oJMMfVwvOukcTfSSe9KqtMpeLU3d9ad9xz
A2MiGTXrGyBZx84qro8hWVqd8e2zB+Tb+OwJQrWx8SKOIBPsrPWajTQRW2iroo7yQnhC7I9ZxD5J
yovem6zh951Fyrlqrz8iRB3WeQ9AtXkL0PmEdHDCaUh/W4MSnafGmmY+i3LB9k2XrgQlJ9e+7V+B
jxNQfAkEVB/2VK6qJBOwUe8C3BF4dPZV1tV3oi0vV3tq+lFE6cO4oyEjSTMe7Z9jrIPNKhRBPMOx
ozuqIchlXuyPaGSm80rX/lp+cLAr4hXw15uVCDxHMSTBKm2yO7zVBkQzK3hznzjpJwJSyccKB1fj
S0favhVTAaK2E/ygnPUwBQh3BTBvDzbZcQlg77TlXcig43nqTbLauvxetR6JTSJxx+y1d3ki0SU4
EQ3RRkB5dOm0VkAtvDNzKDzaNopvK0L8OsRjOzbiLEjhrv5EPvF5BRK4DKLj8D8xPOCE3+aXq1I1
mP3mSRPAcTkIoiKUIoSTf75EvLrbfw3X7hFwKGpJ1FjHIAPr36vC9wzbUkC7T2HK/L565r9GcSof
uV8uHeU7mbAv2U2hallhKHtx5/XfPCd5tWq4QfwqWnxLV5RXvrkxshwIwMv3dlJzIfX7XKZQNAjF
eTRKcn3uq7i7DPj2dd1rNQ3ftMxt+o68cOggDH3b9U84KyAZmRJmwVnXNQACMf3vVxqNetvxk0Xl
56TDhjzuR2VjiPCIdqiq4HMAieGBy30EW0YmxGXg8dboK2a2KvR+/aXc1Qdzv+6F1f9gYFL/qgY3
BUYlGyxopBO/+ZRgxf1eYxSB0Pa+u8XUzZmdgSdPDF687t/giTQbIjiibfc6teFk3mFYIma+rS+p
OL5gPRM83MCt58o5K0g7o57MB0cQ/QJq+B4WJQIIHhCsqZSBzA3nKsdMAWmkwQAO4enr9oqx0M6I
9YykrHf0X/5/sQZekqgYK6St/op6JVbUgGmypSUH8U8k9UwcGckHH7chp+bYM0eC21aDKjU3HLnr
pcBDvSZ7AMWqyYBoCyKEjuiUjSt8p6ETJbdVQE6esfp5nFmxv1tiodzQch8nhjJYWwSY5g0UYht7
GJ6rzQhfXkdP1C92j566OtpPp3PbhnDP21SDuCgVfSyaOxcXA9v1gV753xd+y7VUMhHku73dRnPo
xsTSGW8H7EEfLLgrprjxJ4+QNITaGpV8R56ML/oByhx8UQHFyFJfwC4ECylb5gDOke+Skv/0Iw3s
K5ZzuUyOuIrF5m/HLG7yO18Njs+F5FQvHOW+y7BJSib8Z6bbehhxsSALHwfENBwI9EjAdTegSp9i
FZZuVQu3wcuqoYBw4d2qTwnHWsqiPH763pitgnPlaoJYTdG6O+61o3FHPP4fElqNp0uyl9C0lLup
2Vif+g0Md8922JGm1vv1MnqtaPhiAa32ynJ0c2X4BDOZQ2ShlOF594+ZuBHzT08WNaa84MmJAqC7
Sgd1suHItHOZhRkmAXm6HsCoM4mOk2Uj6xRDo9M9ksU7Wr8RyOWRfyHKLcsuZWH/+JGxOB54oG6u
KdLTZctxkB6IhXhey98M3z3IwfABo/lHtJCnvg6hsTxUSV5f2H+20qRKff3ms7ZBl3rtmkA6Z/MX
TiAd0FReKULHqC9EBcz3nBCWXa9ZKw3hhpl5sOnJr17zrDZRzTrnuli5hiMzNmx/Z34pVRE/+DMv
6mDrz7S/nKZz5+g88CjuogZ3n7Ts4HLn3Uv5ld/u5O4iL5KO7qPvZdVMq2W1i8dkV8WdWt3OcD9F
oobM21ZUphg1L7KOy5R34/ZIHxw79f18S0tMxUyNyYgMdSfEybRY1EHIY4bJxBl1iOOCrezC83E3
vUwGKUrGi44V+Zj6qNywKIi3GyU2ni9VDoPNlnQh

`protect end_protected

