��/  H�u�2<�k�pY��iI��1��E]u=�݄�8��J�59�I�c�����Y���	�����o�X�� ��F�xa����u(+E�kbM��&"z�~L]��ç�%�V3��:������Cj�b�A�U�O���I [ �-��]�*�: w��[� b���q�����֒7�k~���p2|JWFӮ��ĕhU���+<��x��S���T��`Hw����������7B�S8��ul�2|���*�!w����V[Nc��������kJS�z�t�$$ӊl�us�7�d{��t�,�f��9� |�y���!��=M$��J�����x��d#s7���>CNzI��r[��Lg?j�a��������,!A�偏���m���s��fs���x!�Sw8�>Q.�!T�%̪C�I'sɷ�-,D��KkO�e�%J����e9��}T��GQӸ땆i�%��U#�%*Nu�F�a�(G�?�!���(«=�~ 3M����Y�-Dgke�x�@��c��QL~s�$8��9@ l3�|�`ZX�Z&��l��Љ5���MP .v@S��Q�'��>}�P�g��>�Fe|R&:'�Y�^�Ɗ� w����Zm���蔠)�{��Pv+������㐢f��\�B$;(T�����Tjϼ�~ׇ�g����4��QX'��N�B*�����ʢ����U�����&��}oZ4l�#}���ϣ��$�B�Ʒd���rf茶~��t,r�y`�A��[:V�įB�Ȗ���[�Ws��~�~_�q6V����o��B�̟�fF�/%��X#�[3=�41�U����H�ץ�f��,Z�ʿ��N����b���*]]�����G����u�(�! YU���G��n�u~�&{ �]��O)�˗���~��w� IÓ]��+Dlhtf��Ƞ��SX�b6��vŵ�g�y�V`�.x����E���M��ֈ��9i�)A1q���������Y�i�o0�)��Q��l�I�sE`�sC��H�V����S�C\��W��43L��`?��	v��O}C�^���@���?�n��o;>˅��n�|p?h�@-O��Sdm���9�_�D�(�tφ	zp0J}�����4ɋ�;�IG��'΍���D�*���t�� ��	�U5��ˁ��4���պ�N��O!��H���.��'j�Ͳ$����Ҋh3���;��>��T�8(J|�[p�}�1�Wo�=�0y��:�Eg��2+���ZP6�����gy�t/�flK~sk"�S]&AG�-1roB�K���a�|����T��A��,+U�{�%�)C��3nTf���'~��Y�\x��B�:/x��iA�S�8�1�(C�5��xX��a��ߺ�������ܦ� M���A�-���rg�����������c��\�V��N)C�R���H��͛�f��.ؙi7�޸�Y�_:�|(��p"��%�+7nf��"b��A���O�6'6�����a	V��6r��ݞ��Yi��'�#��Z!uAWޝ?�?\�m��mvfZli���[-���*�����
�Ise�	N�%�G���g��7�-.^��5��d?����E�L�����"R%��K���o��-6彿�ƴ̏BeʮS�ݘ�I�j?��TPP($�N˙a�3���F�� $D�+�)>c/O�؈���r����rcFQ�B��� ���it7�@6.�1���:��4�{P^+�0w��L���#MgI�m�LBjMeK �%��F�@ɒ��ƥ�.gK�z[3"wQ����b�-6��j����g��a���`'T�=@�G:�4���];ͷСV���}ӏ�!k���
�_' ��*R���j�p;�%Y֏%�T���jDL6��s� ��	�c� y�3.��f�W��Ԍ}�r�Y�>Z/��^ z���15&?%@�u:T��d��l[Ka�����"��>=��5��+	+Uu�ŀ���큧�)�H��_�*��� pK�f��}��8����삛N��~��j)G��d$韉ۗQf2�X�76�r��� v;j,�*\��D1F�}[ߒ�=	����z�-<�U�-#�&�mZƺ�k��b���Z��ԝ-\�o���U�|�>��j=�_�ub4�,nt�%Tٛ�b�_��l��]���V�٥�#�nAf � ��{�`C9E�S��B�q�N6��6ve�Z�(@�C��p�ʔ�J� �J���U~�{ܙ��#��ZI@E�z�t�+�
����̲.��`0Y�����}��Ǻ��^�yp����
�����6�T�ڜ�G[ɺ�����s����i�6X%�e�.0��Ӿ(Kgea���.�UNR�J �85߉�6�����ď~��- 褴8�(]�d-o�4���~I�l������c��n�2&�È���}}��T�S�5_����c��ԍ�S��}eQ�4��&��s�(�^[u��~����|��K�2�Vh��V C��E:͂�z�߬�%������m6��v��[��:��$�+e6���i`��M��x�����u�;@9e���[�Q&~�Lp�	U��,kp�#vZ3�v���K��P�d1��s|W}<(�d+�sΜ,����E3���'���!#@:��ˈ��|�eK���Z[f)E~'�4�^����f�]X*��t�MT&1߀��-tW��X�/�Q��&�g�/��OX�������20Zu�`�3���}t$���J�J�ό�|�~0�ZXkl�3�E [[���{�&U����Q2�L����j����E�>��1�̋���z�מr?+X��+p+���T~���<+t� W��嫤�&���8xg(j-�T���a�����xz��ч�u��b���ƷQ��{�-$���z������և���c� Zuj��.��ژE���ع�9=���?X�ӎXK@����^|K�z�$���E��cɹ����I�������G�R�se�lwB����q�YYV������_;U9j��j[��|��S������|e�Vz�!x~8��y�m�:ǎ~� �l����_^f�q��ly�*PI8J�F�0k�Ju}��#��w̖]= T�3<�����M�7T#������q7�^V�A�!����􀏚+���������	�ML���T7���mz?����!�O7��~�k����q*v�N�`[P���o� 3��tQ$��D���c�JDf^�.���N�'X�ѭ~��q�ȥƪzSē1	�
�U�g��O�/r�*��C��0�� jzWάUuƆ��y|m/�I~��P��Z�3?�ڡ��bO��_�<!�����0��Ԗ��Ȇ��j��s�TF�XU�z<M0��&���޼��Ȩ�d� (�(�{M8�@^e�6��x~�n�@���2ち��^E��U�����tQ�Rv*Uf%ܐ��5K~���2��\dӇ��;�H�KЌ��W�|rcK�<Ad-91�{�1��(e�Ct���)wd2��3 7�D�%��5�n��1�9����KJv���.���:w�*��� ������
_�s��	p�vx%2�H��s&4�����y/�A0��r��K8�b8zH���K"����*)�<�Jz� ���b'�~�r
�ٽA!O�zw�g��˖�ߖl�r���X�ܔߛ;}���qy�c�ފqHĥ#��e{}�H��π0�u��(t��uoك�R�Y�і�^z5S(�g>f�n4F��\k�Y�W%�Ej�j�e��'�/�W��;AqҦ��|6���*�P{p���ڨ�ۅ�g�b�:�Ҟ�y�p��p�8$��K�!�4�vt�)��$��"w�b�w�E�d^�ڤŪ!��#$�R�0~�J���jAG�Z�bh�\�x�K>:<$�s���/���[c�"����^�/�<��.!9rN��B4�Pœ��^��<�d;jɖ�=���@�CW�o�ࢷ�b싫i(���g���^/~ȅ�'mz��:H4��;����P(6�M"w�S�{�OF5/���q��.o$��$倭,�L�E�ݥ��n�S�}%x�U�,��� Ʊ	V�p����c��H��GV�|XF%� �u���{�H໛dΣ��;CpPc��n�*��H�{mk�	SiPF��Y�}��*��p)�ih�a��.����
t�y+@��_��%��{Qg�}��f�>Ȕ|�'2%����Ց��%�>5���ۿ&Ϻih�)\tSΥТ2�dI_*���h��Wõm�F�?����t�Z����g]Ԑ�<��'^�ʇcJ��ꋑ��bB;ל���~D�WQK����o�w��7��7;UL�ӽF�Rb@���0,L��u�
���,|�	#��,�Ҿ|��\�j�� �Lߥ�h����)�|�&C��t}}wW*l�lP�u�{q%����Iۨ��}�q��󤖼��#%���;�q@C@�/U����-�N<���}m� K��.y] ]�'��A1,/֮I�U���b���H����	b����M�)��'�/̗ܳB�ĕ���	���j��'Q�l� ���0�HT���Q`���?}���"�r��P�O��5�ڎ�4i�����qO��8�-` k��43��t��'!l�m�t)��|����:��+X/�1��ߛ�	�GT����ZK����������ӟ���>�%Gy��<V�4�Zd�	�v��/���7�,~�K$���@G~�P�qEwn�e���Ai�Ơ=��h�SΓ�<���Fٹ\�r�0�������_>d�W�[�^/BU:�
�$ tJ����
�!"k�>8�4g���3FM�?�8+����5SV�K�*A���1��P�+]!�B9�m"y�Y��*�U
&i�}Ի2o@� ��Y���:��"�G�i!��4��M�T�Ӗyi���X	�������P�ȞȎ� W�.#_п��V�)�y�G�$Kdr�dCZw4a��ƣ�63�>iP�:��?m�뵴����Z�J[Q�oHS�rM�BS�'�WA�Āl/���<�/��K��w�0�4�#�h�\�%:f�D�-/��=�CS.�[�����g��
hH���W�y��s�c?�B^��Ao𷨝�����D�����i��D+5���4���ھJr�/j�[��{�R�59p���Ud���q�L��}&��ԦD���"ð��x)�����G{y�,V�'$��tW�D��\�UA�}\��u��*�~�c|5@��5;ʲgń{�?%�(��M*���L��OO_�L	ݐ� +a��V��n�{\ |?��;�ɀ��U���6}���糜æ�T\�A�8\�v_���B�6?�V���
m�a���:ؕ�	<�ye��Ҡ�_��hN�«^�,I��V���)��o�3r-^�O��t����Vd�����-�lnQ�AVH=��^r�$ŉI�1� ���\~A^	�?)΄d���MF���X
ۥ!79�����hX���Ǻ'}�J�uD�d��VG	����j�kY6�J5� ��`�YX:|C��\�N��t&��6:(�C���C<v?rgo/*,�9��a��VI����߉rX�6<"���	Zے����ƹ:�q����H��Fo������[���˽hو�b�}*=Z�Ѧ\9^ꗡ��mn�ǆ���lσf';�]?�
"X2�x04�\��<�8�o�`����`�{Vr��$�۱ү���I����Ȣ�����J�,�85j����YC�T��	#�_w5�&��c�b$5�bG9Ә�+e8�"kÎ���&ǛY���Uu5��8
�^N�OƷv��6�
G:����5)� ��ơ.��aO�5\�v�=ڰ@c��/A�|w �p[vp����HY�b�8φgʒ:����ٺ�	�8s�������^Q��~�l{)'�ɔ���q��)� w�Ȱ������r*��A
��M8����+�[�1G�K� ����5[�Qoi|a��V)Z�ǻ.�j$�D��u�h�T������NQ���<4FX�u��KG=-"
��T��־��:K�Y�Gb��S�Lʯ�$�m�[:��m�q#��}�fDa��G+����\���QJr(��)���5Bյ����LkcYL©��&pJu|����s!BB��\1�'�'�y���d�k1Q(�k�U�Z�2��}	B4)�c�pG��e��9�z*��[w�5����eV�>�b;>�[������Yi�İ�(���C�{��m�c��!W�K
������¿0��Y�V�<Y0\P���#Ŕ�Y�O���gK
da����̋7����!eW��ߐ��}v���j�`@��L����Q�A`\���������g������J{~�̙-6/�ɃdI�����h�>^ҭּ�72H�Y5�`�}��>�X����l�Xl�'�R��^E�|��ux���Q�a=������u�|��gq�G��>�؝D�VsT��2�X0�V�H@��ڦ�ɚVO4 �h \���H��	]�'���;�9Y��o�є5i�QD�k��.Z��C;�޸Ź�]�.�1{q�d�����.&o8�����܆qdA��V:j	�Lڠ<�./KQ?����7Í-�G� #߮M-	}���o�(��?"K�>n�$T"Kɒ�IT�����BI��,�����BT>���R�諍"�͜�������m�㨴�,=O�_��I�c�V�~$���[�.˹}���8��-���0̇�YzA��/���[�{�o�� ��ıNu���2�Łϧ2/�,�����,�[6Z��Q�K��mW�d��Y�
���`�-�W�5{���j�^̠����F��gH�B��L����q��i��ķ�MIf/W^7���kJu���t��ْ)E��: 3إuDNE�����2Q�!7��K�,��Ă�?]EY�*�=W�ݛ�I�i��l2����Ҹ����+��b����%���/�f z$���)�B�l�?�Y[�f�ZԀZ*I�PLI۽B?��\수�{m2��t���H"�1"
���>��S�[K,�B���J,(X�w������t[3�R�R�h>�w�����5��;,/k"v���ٙ��AAI�Ga���=�+�֢'�S��8��?�r㪟K�����u�CT���#r$��"������1?|����i!�T� 	�^��[��*O���3��AG�e��V��؅͝�7�>�~y�F�H�-���v
�_�$�k���iP/]%ڃ� �Edԁ�@A�o:��m�u��AG��.3`��q�W/x�F���8p3�ąS�3��A�h�:o��8��X�Jq��lF��̔�0j�:� ���o뼢�;�MϨx	�\e�����s����)�y������,A�N҈�@��XU�a\Gw�D�,F�C�x�1��	H���C��`�f��]W�3��!!r��'���ОU�$�G�����~U�����as�|��w,HR�=
�%�!�	����?y �]S�����\��7e+�tG��+�����k�|�p9O�B`ȃ����ٻ3O�8���q����y��r ��C��nIE����c0/ą�R~�2��w�Ԧ:+y��� �O���"��ZY�P�Xb�,��l��������a_��b�w��"&�����h>��'-/��`X��N�[s�&l9��eܱA_�kA�eGVS+�O����#x:z�rI;LH�O+��ѝ��w���ok*^=~� �~�3 .74XF�f.�~j�я�&��#�����&��ш�1t������A)��$�!Sd8��	�j;�N�?�栗`d�s�.X��W|��:�yX*乷աPNZ�W(�0��Cc��S�6����[��{&��~�!9`�|ڙ�k����%N�cR�K?^����;���'�]���j���%��ꨡ�ADN`=��f����Õov�Ǹ�� �y5��D>F����`��۱_�~n`,/:�d�9�k�ӄ�q�mkR�EA��~B����s�j�6�L�*�鴉f��9�%���,����e���"l��=�׳�ڂ8pq C*����i�
4z$B�N��8��D�z|4Q���x��$,u}7��th� �����!{�uS�N����:�9�{�V����4�Mqa���S�0(T!�l�UGMnmf8С|TW�H��">P��`�ǈ���Ȱ�ܶ���k��}�a�^�M����
��_���z�z�cҴ�-)���� %~x�P|��^�s��k��ֱ2~(CW��l�}᭪F*u-�ʽM:>�âTO ]>��7zq5�7fŘ/2�)���H�b�*�C��t��j�[V�2a���:���h[?^?�
^��
�L@��.� ̐���'D��:Zë��d���k6���}ق���x�!LF,j�w?�Iax��Y���8 ���+�.�0ۣ�V�~r���J��G�_A}�wHʍj����i���O�:��� �~�5��+��	 ��컗�@T ��ӊ4v���Y`'���*���p���)�G��
���6HXƃ=?�E�>�
t�
��FB�Hf�g/��.0t�q�*���r�8��.�i�梿ġ��Uk�X�<]$��Qg,�n�� �+���g���~�A	���{8�Xd�D�Y�}��%Mc���:j����,8(�k����~�}�(ϥ]٠A�v1gBo��Z����iZ���-��G�iE�=�6V�4�9�a.�'�A%i/�jk�f�\��s��'�����PYFĆ�(��2����~$|" !�Y��饢x�ߖ>���+��הi�����D�!���4��"����d�|jC�5&��v��P������7�YRp����pkj�[����9�c;S>�㊿O�Ad(�'�G�{�8|Or.3$����M�팿�X}#����n%dV9�<��<�St�iM)f���QJ�bt�U_�?T�2X������C�����'���`����Ff�C�A�e�bY�L
EZΫ5p�dȀgt���>hٮw��g<Ĩ�;O���դ�]g;�c}=��A��lK�M��wpCFDy�f_�E�����+��s�*X�oB�'�؋��n 8wED�\���j �?(Ed��Tz�#x�a�[$�d�F��2z9HN(D �H�4G/4���� Y$p�&?`6߭V%>71����>x�lbf�����b���(���A���u���a�HJ5��� ��O���l�r������� ��#�m�����4jؘ}C�5U�Q-�^`���+|6a�eW��P�����NV�h
Z��^�Q+�� ���� �L�T)����iqS�8�����nt=�(��w� �h��3�d�]1ԯ"�^�q!
pG�(������5ڊ�ȌKR\�E�ua;6(lQq�{�mF�Q1Cҍxa%�n��������U������pЫHw͹��K`Lc�Ⱦ�w��4���<�p�U�'�`N.�&~��[j^ԳX]���_\a&�n�Kq�T����YW�� 6�\�����Ƶ�0*�گ��@������(��d��K���c�GF,U�� ӼD�J}
�\U�,e���j	m[�%w���,��$�s��ό"|\�b�:5l�A	-�e�*���2%��&a�s��I��R��P +�H|�����[�◠&�N�� ��}����q;za��$�H�0�f@��Ϗz�N�����ov9���>g��/��dׅr#���������M��k\1��F���G���9|�s@ ql7���FB6�"n0A�;J�����ͤ�:�yQi��Nt{E	z:�����᩾;�|63�p�v�̻�Y���� Û�<	�L�N��x��������ʡ
:�F��c\��O����1sy�ѻ�Д�1�:6�}zE�`c�D���	֝g7�)�3W�O��A�T��&*�����L��P�!����������t߅�{�:tI���~;r鬦�Ӱ���ߍ�����X��qn��;aI���h���h�dx�R�!.���Xks�ܺzi{�YGm}�|�8P���@-Pݽ{�k��*� (R��1�-�G�����t�q�p�p|����~cP���{�i��7X&q=E&��)K�R�RF��Wq4��������ʢ�K��z��euJC=*>N��Ii���1�x��;@X�;�>d�rfy;sD��{R*@ 1�;��K��r��(��,ﳄ�wA�,��/:B-%�kO~�nJ��ڌe�f?)@_���RL�]����ј�&�,����"��[�A���O.�E�ߵ#Ɓ�Y8�X�_3�Yw��Ձ��n�w��^�H���5��!��tЎ�h��蒽#Zk#�a��򪃷��K��<�<V�)<���Q(Wr_��-wkr�{mH�4�����;o`�5�#{(���+7�{��9T<�B����:wy عKĞƒ���!��gk�UҐ`أ�}�4R�W�l�%f�^j��r��4����sLM�6�d^�f@���7��%0�1>��T��E���'�|�EQ��!��(���Â��2�s�ԱȈ~f�lb?����O���[n��i��+�.�~~����'}�/�^�ﷲ��$�[R�!�{~B}7.��ϯ�ʱ�4���nf{1�~Ê/�r�g[�~���($Ƌ���lr�_�{�R�H"xA����1M�g(qq6 :]��(�7�<@��҉��$�b�1��g`FEI�v�m���Hٳ�rt���R�����/OoW<��դ(���H�ud�(kJ��F˕�[���x.kP���w"�i�ǧ��.�Z��t��ծ��7�ڲ|-[ڳ���@��	��7�d���m��	�e�=���f�����>?{���m��!��d��}X�OJ�tEί<$s�3�ڂ�{#M��-B�bD�uΌ�6!��[�O�A��rz?'a�e}�����2	0��zl�vq���;"'����Mwj�U2Nݤ���YLD-��ƺɢ`�m"$<X$/0�b���]_%%�VE�1|�ls�0:,���bJS�}�����ؒ�*�M�@�@E�C�Nf59�� ��8��J�<��Xi�*�CTi�fl�ф�W���֔E[�Q�D�g�G�U_�u�Ǆ�B��ri��-����&���1�B�?|��	������u</ؓ9�Nn/%m�͑�Dc�T룉T���Xit��5G�2�[��.;�W�i3I���7��mNw�b��!�չ���,6py�n�A���
r��F�Qd K�t9���Ƹ"�a1P�gN�T���j�6µ��f=��[��kԕ���qn�-�]pG`��4(5M�R-���(���t�NR	�e����HA鏛�&tE����jr!����b�VD6�R�ꯐ�"��mkE��m6rW�S;-�������Á9�@F3~�D;�O�>Q�����B��;m����`��k�9�����ìS��I`���Sw�Z��
��:ܘ��~���"�;t����o�*w�#	hԿi�2�����4�>��s��t�Nu(�د������@䪗,ۖ������Qa��w��of�����H�dc����d�����z?��8���-j��P� �s�๕��{^�{�j��qΣ2"f��''�a�m�?3�a�^(�{�{���D>3�M;�!��<ᣬr_h�(��T4Ա1<������#t�L�n��*��.��d�>������� nD#�D'-��5(S/�s��J�e����	e9/�B͢D~�7^��<�6�3n?�V�q-
� �66���*,�H9�"nY�W�{�h]I�����)��?�]�2��� ���ב1���\
��i���)?[��A~\�6,�#w~9��w�q>������a�3�m�`4Ny_�CO�$"��Y��S�
q�\	P�B`˨fP�(����7Ef)gݶ��!�%�/�݀�w ��(���=u����w�zJ:�]���Ye>
\�hW��*���8��CHP�h�K��m��v(݃Ӽ�(MS<�Q��M�����3�c;7�v�Ss��v,���#�*��zi���j�5p�tf�����ȵ�W>�����0�q�Vz"d��a4'҂�E�9��s�R!���z*=�rJ�AB���^��/����M{ a��)��D�BY� C�P���R�
KV�!�w��܎;���6�}S�=gJ�{��ey:�[ˡ]L�K8��H��)�ϸC�:��n����׈�'/!Շyf\
ÂQ^ۅ�E
��qpi�U���U1�!��qͦ�ۃU�\$W��>�����n���o�2��o��7z8��&�����c��)	�(,��ѣ�%�4�K���졨�"������Sz�Mz.��i��W�jl�$va����Rè@���=ͅ�~�,�5tV_*Z7�lDp�{L}3�����8��1��1	+:8����5i��qWJ?��dy;{j¶7/��	�	��m��-(�|�V'�ڏ=�J�u�{�!1�z:肕	�n8t[��?�f�nֿݕj �]��0�7h�-�#�r�[�;<8|���V?��g�(�iaY3�9�S>���������QXd�}�Q���{��cǝ���+�f��N���qi��Sk��(W��o^�t:ĪܚI�G�7؄d�<0��2r�\�^��d"��i�%����ɴ�B�I���=Q�1i��z��Hei����+t���ߵ+�h�r�HaC�:�2��O�&s�Sr�ey�C!eߝ{�_�H-�c��ٲ�T�;)؉�y��Ș�T� �]�_�����?��U��RI���7�ɞ��b!�u��Y����ъ���Ȼ��Եg!��W��<|``8�m]���u�D�̄��J��J)�OCcc"�NK��ҩ0Jۄ��4�c��[m������!z��I�U;���3�lm�@�O�A�!U��3"$�|[��Q�T����>�Da�-b��wg 99M�|x:TF\8$E@k�{.n�:�5�����]θ��yi��ӝ���_Ҥj���O���6���[T�I�T�Lj:q��IZ@}Y�g������a�ocÓi~{!qBGPT�VKߋ�
�(���1~�Qe}U�k�l��_�bڱt��tzz��͵%������v��-=m��D���&���򘉒�"k�b^/�)�:�PV�d��0�T�uIJ^�T��.�>ΰ�2�� ���4?
��"�`>�����:۽y}s�(,�u'n��7.c3h�Q�g��tY,XMt�W�#�Og�rh?�:={��O5�9�m8 ��͢������c�2)49_{����r��+(�q�u�8�$�����<%��Z7/��j�"��r9�+�w7�T���A�pw�׉v�6oϓ��>�N�>��C|�,���'*J1m�=\Wg@K�1�=q�&|a��ީ4	� ��[���9��ɹ����Bt3iŕ������g��6W�[��H�p=���e�(��c�tG���$����:������R^�7��`{ p�P���-�s-+�6VMN�+��>Ş\7 G}��П���ا��&���Z�Vh��DwsqmC��%��������+r�\'w��Y�bP�����wK�N�LI�uM��.��Խ ���g�m4�g묗v��K�V�V���b�i�0�DV"���1�����:�k�t5׬�S�(v7)'
�T��;5�h���łi�%!,�yb¡?�B�t`(ۀM�
���e�xn�aèeݔ�G���i=�fF��^II%u�W�"]tF´䋗�=8�}��ltw�6��B��ګ��Y��=N ����2[�#�|k.����r�D�E����S��[�x�aN^�����ךeP}�<y_]��j.�l�pXq
Aĸ=���ߞ��V��T�����R��@���!�Ƅ/�)�Vp��;�M[��!?~��x17��l��T�����)�X8~�����%�@^C3�b���V���ҁX��b|���[ǔ��-2�I�{�و
2���X�3p# Í��͛M��ł$���G����$a�#:����t��������	��)4����Fxn��k�2� �_�j�c��J�h�96�bh��DO���+'ܣC"�qG2�5")�@뻳�\�5�l�K�R�:ć8����2R�Svn�w�a &e�g�>SK�J��v����lT����G��t�S'�c:���XS�"4�̓�8I/��%���	���:Y�вŒ��a��������$�e��G7c�Qm�9P1�^|��2��'K,�F�E�R���I�F�3����L�kҸ"�㿒U'B�'�O�)3�E2�GE��4�B��:�� #q5�w�c%���l��~��5tS�Ư�'6��<��
��쏮ʢ)J�����Li�����	�����@����+ܷ��:׋�Rr�;��{�æ/��8�zH>�)���@�.	��F�]a�J:S�E�\�Ǒ���g�A�ZW��;�J�<�6���x��3�S�]=��yܜ`R�1�옢��uWa�]~n^Y��\��Zk�Pb�R��׸<���lP*�@/���w��B�E�x��V粻�_��ti�v��7���){���BB�P�,)��]^K���᪗�n��m��7��g�{8@��&�P���u��0֮4܈JD���v��n��F�B�<��#&&�v�\���M
�*%��ctʐq��쯞�3��D'7��`5q�
����[�ؕE��쑊?)��&�U�m���*�gR��OG5�M��J�@fU�ӢBO�^���u\mY�n�|"�'wL���:�fDO<����F��͔>!�y���סb�Vrd�Ae3Rp��HlwqF{�?r�V]�>akWf��Q�8�kv��;�������RJ�:Sh������<�� ��e4P���С��ɷ�nON����q���=c:�tY棚'B%��|g_�J�y�a#��3��2aY^F尺&����L�LQJ=v���	��١��D�Dn�]@b�{�~�M���N��>��C��3uc�����<T�j�UX4�Z�M��RU%I���k[Q�Z\3V!R*��>0���]>�[�G��N����<�~�g�eI��K��Bϖ�K=j�e:8?�p�j���DXL��=ȵ�b�H�^�j�B�oCj�����tO�uZ&��]%y	Y��;�Ed�2A�S������S1�%g*ݷk�%v4�f�ps!⼺[�.�����3$b�ҾAoz$��K0��l��qd#KN�CD�^PTO�:�p�~C��1���v�|�L�R���이G�2��?��<z�@��(��-��<������钨Kӝ��U��R�_��l�x��P",;D�+�b9�P�Cʶ��c�J>c�@��L�|�c���[��{P"K�Pޫ�,nU'،}ÜW�@��!���kq{�*%���W���\�����F����,�}�f�7�(��0
F�����{�Bޘ@��hV�R��oa3D�}���	�FP��֝x�7Y|v�J��C"�VW�[�*&y�}��l�<lIYٹ�ބ�|@��%2k����N��Ѿ ��V�8O!X�L_®e�Q=����@�ȝ����S.b�jH=k��k^!�4��ӌ����d������)�H����٤sG5��!U��%��J|�8��)�1�P����$���}ߢ1��~�F�������&�/[�W�A�یxe�;y?�Xr0������[笟S��؝���R�h�b�9�&Z�^�"�9�k(��ʓ�}��d^�Rw���q�ɝ��#B*m9�f�]�]�� �����䇭��da:���xU�N;�7�q�#*7�޻�C�T�~�3�S xϮ62o�ҍ���l�@�h�Z�HO�#9�@�m��+ڗ|.�[<�6z~���A�'ɗ��┄䐺K �h`+-d��L����L�j�*ۨ��B�@���a�]<,!0��)#J����5��m�L�dR�O�9ۼ��}��-��vH��~"!׮=5ݴ8�<c�'HP�o��=VV�g�������4+�������֥��K̐�9;I�yx���wgb��\���X���5��rM����u���5t�]i*`=��u�O�e���5���N�N�J������vh�F^�� �~R�jT_S/)�p�wa��A8�����bk8�%#������<2�-�l��9�4�`�Y���x $��O�vB��a�
����"!�/�-u�ۚ����ʳ6��]Us�x�#}��j]��Oŀz�G����<R7�Յ�&O#���v����9?'7�Vk�)9Q��]��~V����V9.{����EW�dÀRȝ�j�,���舥X��輞�� �.9s��_v�k��.�"b3E�L#�S#�ͨM���"�%�>Q�� \9�:�=��$�A���h
�t+���Ɲ/�~�yO�L�2�j��4������R����_Aq�&EȺ��AQbZ�un�zu�"ȃ�'H��[S�X�FMPsOk6"��ʥ$����^�BY�6ےL�"͡^���`�6"T߇���Q<���U���o���̦^],�$��]\�b;t�@ߺ|��Mr+Ρ����Qś�ZWV4׵��t�,�ʧ��[�q�2��UË�q��H"@l|,��\ū-�Ԑ�i��W��0/��Q8�{�ӹ�!M �y��eI�~�������^�{�PI��{n�4/o����Q	�h��q�!Fr��A�Ծ�ʎpﯵ<����Kx�!���Bەk�Q ��wrG�H��WS�n��"Em���j
�Ai䅥]�\Q��?���	�S���$�����=�pB՜�G�rc��tr�<��Y;6��Vi8hw����C��c+���d�/ao��O]@I��s�M�и�4�]#C�n����2Rk����F�т�0��~�'�?�M��;�Q��g���ea���;�Y��t& rH�N � �����ۀ>�������0�v,.�e(k%�^��P�X���t�Srl��m"�k�͹�Jc�������%u� �\�!~�P|9��7�xaH�C�� ��կ�@(/�'6`O7�~V [�[-T�^N<XDin/����l�d��ح:�h��*�&���zMH(ܷKm����q,��飑���S��J� 13=.6�FX%��[��(�@��P�j�"L��+'7rc�����W�E�:d��`�f(ृ%{8��#Y[��ů��=���m~G� �R�m*��p�mCq��2\����Z�<��{jN,L���A��m�)����r�@�P���x�'q����`�QN�K�5,����"Ra \-4ё����\�ky�6�+b�+�KkǍ>S$��0Wb{P�&�t�@�|�S���EjXE� @��Y:��V��ågdĬ�K���l*�7^���I2K�����[K���̝t��|<ҟa�-p�ۼ�t	t �U7�$�M^��n���tO)�P�.��L�<�0ܱ:|����ܟ� /	�G�#�p�U����ֱfh�$|�=s�$D��`���K��E��{���&$�>�����4�l?�/@�=��BҦ{�d��}��ޕ;f�f�F�V�
�~��?�K�������$�*�+���g�t��C��c��}���.��AM�H)"�k;�,���"� wK�Y	����X�O��x�o~C�-#*��}�(Yb%.5#e�-��*_VS�~}���npj���z�7����oN��F<����A����Qr'�Y1��q]�����|H� I�6S�6�h9!7/\7|�?�( y���z�[����-QU9gI1h��Q��;::�){غk1��l��Q�e��هd[��z|GSH��lƩ֮��
բxN[w%�7�M�Zp3�Ȳ�I��ݠ�R~	��o�^�F�ߔ�w�E�1]+�� 6,��������=�U�C,��S	�z��&ԉ��:9���y4U�B�;}��i9�vH�j��e�Ezi�ɉ��}��F(.�*V_f8�҆��ߔ����O�"�o&�E�eh��;�ʐ��u;*���V��9o��c����#�\'�T�A+p�&��
K<��z��P��tTW��s��N�	1�^�0M|��w ��`�~zX�=�'.���+������.���=w\?�r$��ly��Y*!��\I���	�A7���$u�Q������Y�:>���2 ���+�+`�&�G��m��m�>O랯'���Є��{��@�s	"p��Z�����U]w�&�}j��\�Z�7kv&)*	�~�5;\?��X���^%>K_����nZ2���RH�xX�|<��������g�dN�a�:���=,��lY�f���Y��\�#E���ϵ11ig|Z����h�vo"���Ccr(�Li�aEV����?�j���� hA�ܺ5`ݒs�'�k�9�B���ݴ�~���:,��^Ρ�ɲ��������2i�Y�2 ���!�2����M�u?WJ�%QdN���eF��xK:	���_yͤ樎g,�i���#^
����éqZ�Ӫ"r���P-�d���� �ƫ�c�F��H�Yw}^�v�3�B:q�^����F��9��,���](e��q=�eÞ�	�9���n��l�{���{�d��C"��T���N<a�}��~Y=�f~�=^�H���7.Z��a�@��N�6��@��@M�T��f�r<^�����zF��yW�Uě=�}�˅z�#���L����:$j[I�0�v��y�ȳ���y�Ӗ����$FT ��Y~�ވ�'���b��Ԋ�j�����Ƞ�k��#��+K�H���=W�������j�l,>~��ۿ�����'�G��ԍ�Z� |�L���=@��5>�܂�}D҆�ܷ�7۠z�#�ul7��S���?ꓰ�����f�.���v�?	��*�	b�U}��V�� =;��y�&;]���F�>A/�{��pg����_zV)��J�a�ޑ�֑g����V�S&���#�Y����X�E>�:3VQ�Hh���a`³���/�i%��#ojE���&F���Y������	9����b�2vvū0��nf[�`4d��nQЛ3صJ���Ǯ"s3�d�/0	H�k���Avrx���n���+J�k���"�Nb��_
 8��a���	[�`�E\�i%x�ڮ»�x`ǁw�{�$'P'٣@�Ν?&��~����a��'�	ʹC
��V�N��>����cP�1_'h`R�
��n�|��'�N�Ov�M\.���4)+y956ձ�{6�J!���ъ@�B�KM�QqcM���۩|���IV[�5a�81���Q2�������7�y�Ǹ�n���WQ�����,��"�T۟ϼx�UɗC�����n��R��d�8BK��U���[ͧd��6�<�����D;�O����{��� !��[ Թ�9ￕ_(�t��԰�ȝ�����xT$�(kɩ�y����om*�J�a̞������}:�E��߰><��Tw�~�]��/���nC���_Ӆ�Y_<���r����Z]3�E�A��U���*�t����U�[ղz���r��V��)��N��Ε��_@�KOp��e�iRF-#��$ւ�?x�;�+�s�ҹ-�%�e�!4B��U#�����[������T	��_6�(������Ϋ�4~���VH8Al;�X�~fQ��S��m���W���f-w�:l�	���m�3��]�M�G�-{�*d�Z�0a��^I�)#]N+����9M�}��t���0����yo@�QWd�۬�"q�)ln����jRS�z��y��Φso^�Ѻ7�	2����׼���(4*���M4�S����a���0�:k�Q6���=��2/�f�� ,�Ww���@��4b"c�6Q�V��Q-�o�7!=k7�� C+ڞ�+��s��L-�<t
�3��%�t�~ZEX�A��<(E\;I��)QX��_jO��Y��ˁ���l��0c���<:���`y��f�ԱH6V���"a@�����逜3���fR<5�&:�4H���u����4�j���w>�7\ �..�df/7�����G���V�����t�iF����r+ĭ���tdP�!��)&��� J�u]OI_��|#TZ[r��#+ҫf�f��{�X�����x��u ��k��f'�y�W��*A8�qX�C��ؽ4R�����H����f����6iy!����T|��,x؉ ��g�\�"�����8��rjPh:�A����Z=��	K�k�H�P_�k'��X�����!Ģ�yZ��[��}ИcY�$k��/��PER�q��xk!�`���zpl��HM�?ِ�֟T�J	��x����xE ���c	 iIB��:Z5M���Mz'^4��-�����dLk�.�%��S�R^
�qж�;�ڎ��Gr$w9pߜ������c(����)c���|Thj8)	#�9� _G��8��y�a�u>'��]I��e��X���dk����*�7~��/_�L�z �Y��S�R�c����R�N1��%�]r�Gb�e�͢HBj���y�_I��Q��_J#�Q���ƪ^d�<lRٯ&�~%�%M�R�'��і1�hgђ���9�>iS��y'���ՊC�\- ࿳������#Y4$�w��G5e��^=mt)�a͝t��A:�yPz���Q����Ą�s���v�C#�:�r,��&۠e4^g��1|���-��r�^�yF�������Đ��!T���^��
B�1k�9���0٭Q��[� V#�zCJ{sC���r>s�,�	����T��Nb�����<�{&b����ٮ�Ɩ�my�>�8Z��7���>J����
s�6��k�G�>8?�$�n�Nj��ڼ�"���MF:��wu����%�L��L��a�ht�i�W��C>۳��9k�%�$��!���֜�a�h��]V���D���f#t-{�*�)!^]�j�0%Qz΢���R��zX*Z�mxZ�e�u��m芙�h���h���C�K�V��~ͷX/�5�4��Ed����ʀ!�;����YW)qT��`�<�(ctA	�6���>[TYD���D0RM�cqܳ%�\~|��vq$��w��fCl��`b3�o\9Ǭ��|-T��z�V	@�g N	QO�O����t*�@��=���<��0~�x�d�ͳ׷ه�f�+;��>�P#VS8.��>��ٷd_W��^�Jo��`�r���lreF g�"�Ï
�0��MѴ�c�� ߭My��C/���]1�܁��K�s��(�#_u*�Ȯ��Vѝy���'ˠd���?��,aw����f�Rɵ�/I� `�+~�:���u^m���vy�D���|���?�jũ�F�/SP��Wp�β�����6/���Q&�M�j�:�<��h�9`J�����<��՛_Z�-� �5?���Z����C���u�C��I��jG����7���N��2Q�gnu���p�ƙ)�'��ط<��kE��7Cn�Ձ�\X�f��8�NU,I3I_�o?WMO:�����j9q�
ف/�QJA���Y�o��Z�s�߻&uCTEE ���w������eq�ZB�+]C��+�����F�ϒե�ؒ�M�	�X��np��Uܹt��e:����b^�@X�D`pN�*o ���F��b�:�O��J|Flv93����xjU�8�m�����f���~�B������!Oo�a�t���㨬��#r9,A({2��(�1	�l�5wm���7�M!����mu�������zH`�L�'����Å��\6���Ё��W�P�i�s$���Ubr|V�s�-�G�r�U�|�t~�ֹ�#������ˡ�(�V�V�W�+U
A�̳xI#S���\|��=���&R�h����&�jQ�mB���5=T�B�Ěk2�`²�/���(d���d�]U�Q�=�F+u4s��{Ƒ.sY����� ����~�6r�N�Z���u��k��ҁC�%���Duc�)��g]݃*�30�'�&��Ӫ�P���i����*��m�������lt|ş��=��\��ȉ޺UxԵ8��݃:����{;�r\!WsO��22��6
�������I�<h��t6sZA<���	!�VQ�U.��B�؋��S�Ut�:DL��n�8��/�~��@�q#	�!UАc៊Σ���4yB5��T[���W��e�`�
 �{^���}�	��Q���a���G���V�{]��e�Ъ��c�Os��_9M�h�Bp/.�%�ɺ^� ����|��-�˚�B\�k$K�������̄@�˞>^�ϰ�MŢ;�g6سQw�;V����#qnJm_r"����+�Ģ��H�{�F~�k�������G�]�t8f�>J%�6�7�%k<	D�0AH��V��� �h�$�G��٬�"���d�E�{S��-�gD��OM��M;-6Ch����B ����B�O��]��/�{� Z���I�����2 ����t@Iް=��M$Ix�̷����:2U�d��b�j4:Lw��������j0Mִ����J�ܷ"�eRw߾�y$ϝ	��_��wY���ic�_���FxRD���X���\��CiZ��j����z:Y8W�+rZr6B�XR)�}*�A<��죰�-���vteT$b��4T�y�������I$��*īf��|�M���}���V��r�|�e>����/+�D�~
�p��Mx_s0�����	(3��:g(�峌�8�W���������(�^��WƘW��n�D%��U�٩�pCJ6*[����~#��t|�W�oB��z��m@�4�?��2����s���Y����i��(c|����9tL��� �BӦP�"}q�N[g�'2v�������9�G����B�zˣ9����m��u_A�2��{~��u��9f2�3��B��k�	�����'v�:D�o�(%���d��	p$و϶�\ּ�/0u��$w���2�8�g����>�`ݭ��::Yj.sh��`�mj��0'���1�M�E�M���D�kT@�'�����du��F��Z��%��5nS�<���FU#���<�]�T1�:������ʙ�;��ev8�; �}(a���KS�o��w���ԁ/vG��4
"m��/��n��Dg��L#�t"�A9A���T:EÀP���j�]��B¯�gܾ��+{�47sm�Ve2��f���x�h\/if!��?�8�#6�;������-[�3�q��,��0|#\��n������`�h��pHkB�����r��);�B|�j�	��d�qw���Sx����Թ�^j�ٌ�K��g�NƩ"=��
K�O�X[���,t �s���m�h���bU�(8#5����Ŋ�}K&��yX}Y��I�gA����/����"d���ú�M��������u P�F�{�"x2_��f���#+0�rη�ϩ������1�j"@a�k�$"\]�t�ت
��+VY���|��G.��w�����~ζ��x������֥h��NXΑ�쿅�o��¸yЀ��ȋ7�t�����
��ိk�`6�@���vj����=_6��\p��0)�z1�k�~rżuE/X؟�O`}���*���g�1S�Qi�^°�Բ~�
b�����<"J, q���m��;�֙�}<����T#t�
X��^Xpܺ����%n�<1�(%Y4n��Hb#v&��7A����2\'|u�� ���y�jB�X���d<#v+^���F�IS�QZ{	$�w�-���k���fY�ߠ^*!$� ��Β��ԷFb^E�{QJ�u�`�&�;5�kO�ǵ�4�%�����>��0�ε�.��#5�i۴�Zmr݅e����QjKi�(�[�,�V<8:���w�+Y�F�s�%��OL�MsJU���Z֟K��'�J^�y��^Do�A"�H�*�uS��$�5z��i��w?����Vm_U ������u�ArYLkO\�"��&�q� P����K�7m�d�j�E��4Fb��Y�1�z[��b�_M���e(6���F��"��tR� ��BD�#�#��!�t�\g��}"0`Y�x�Ѻ�p�:����dOg����>�REPj���[x���h2?�ګ�.Ԗf��j���;�v$���}��ć�@�GQN�k)_Ws�ѹ�omT�6�	�'������MH��3�?u/�Vt<�\�ɳl��6��p[�{���lث��C�齯* �PGn��K��∢����,�iWj0�oǆ�N0?��eI�o!S[�~Z��@c��K�~��mv���dǇmΒ�C�-�bm֐�$�zd?|�g6:�ևc�6�]��t�X��
 z�iP���+
���`�b��)�g�Z,���6I��1t�E�������-�N���\zJ�n�@�4/�iV)���#�B����o�c��Z��h[m��1���wl2�����^�@цx�������X�dL6������K�$��O��i9ɶ�I�̛@�2bQ/�]� ,������,&�41#�o��TB}��4W	�5��Q$���l&e��6��[�$�w�@�!�_{���*r"j�Aӂ6W��hvE=/4�˂���h8�+��"�1�O�_�N�0����S����>�!����v�Q(�;����K���le���C�Qj���2���=<?�K�i��z��k��H�6dh���蹯A��O�Ϝ�����%��`�����O��H��D~>t�߃q.�υ �/n�n#�2���d��]��7p����L�'?�E(>�oi7$A �MPL�VFfy����6\��c57|���6�I��;Xbz�9+ �߁DF�H,��[7P��t���a�H�7s��_2]�e�9�9���Vht���P	,9-���k[�-�/��A����Y��mB����m�j0c��w���[��U�o&Q�I�����u@q��Kgкgz��Ȁ⻾e�Z8z�5/Q���|�\�E�'tT�E�_���LWۖ�Ŝ^7�MP-	Ӗ�d؀H Т9�w�F��X|�hI�<�ކ��pu�	�PD/^�a�۠a��9г?ӱ\�&���oM��^k��uhE#J�{��|�2��9�㷞�#R~c9nf�C��DR'�0�ٯ�w���1Oۉ�&��P`*i5��̱����|���§�[�i��)`��� a_!Q���/�
7�hq.aX��d$� �Ro�M$ '�uO0G�9�WEI��QW/�Y� +j �c1�e�!����Fr0��\o0B��������5R�,�\��S���vk�7�2vh���G������
I��o)���)��ұR<�8	��鱹p���ú��c���&�F#�!.;�T�S�J����T���4�,@^�t׀a���Z�UV3�l�7{�a>�G�K<��vWHą<�sx��q ��A�@r]�S�5�;�_��ē$}�X�Zg���L�p��o�|;���w�L�|T7�H:�e�+�Ҍ�S��xR�-�
�=�����~t+�(Lt~}N$�U;l �FQ���?�Nۑ��c���[�����_AwR�U�Fp��sԳ|��f���H��k�+��O�t3�u v�;%�8I��9Z]y79�R$�}W�U�5���=u+J�����(z&�Z�w1*�O�Xo0���vo��B|;�(�����#^2e'P�y�2+b����8"�'.rl�'1�.��l�a׎�K��T�����O���>1u����ll��Pxu�O�&i�W�N��R+�̙4�D��d�k\��"��)U}��F`�ܲe���.�߃섹��;�%E�_�K(�p�`�����!�Ȫm�U���2�}Q�e��b+U���ýU�qR���Mt(�s+�A��Z�����q(:.n��_8��.�)��L.��?�AC�X^�@P��U�uZ���r����E��{a���,��r�����;dQaR�
��l���%��Cò���9�=m9�y�4���ْ�T'u����'8Ra�h���҅�=;U��R&ȓA/=��lY���$���K��˧�Y�;&g�2��g��xD<�������Mw>���M��@�����h+%O�F{��t��	���;�R��a�ؙ�Կ�ħ�W��:l�'�*J�P5ï������I����I@`��u'y�Υ�������8��K����Z\�YV{g�U]y���
<�7n�/*C��$[X����=�8�!{�� �oEVx[��o�q�$��V #�5Uݑ6��f�/�w�nQ;`�>d��
����4�mE�;�)Mib����ADh�m$C4���[u�Y�\`��|_��3�SV��C^���[k3���-kT'�/� ̡�kR��sx98)��*�[V�_�s<���1!��G��Y=b/Q��2�W��-$�'u���?�jތ&m\�ΊC$3X*{F�����%��h��D����� g�2���n�{*�n9�����͟��R_�~c���b�r��xTΥK��G�0 �&\*ԞX�^�!��#��,r?|�h����<яcsx̷��.m�"&l��B����<�o�m��I�_Ks����j��<���7�{k{ �9R��In"�l�."�B�R-�dLm���ˤ^&.���ɱ����'��o��m2hf(���9���c�ͬ�k��: 㯨�H���H�B��د�j#�����*�6�5��ԣ�Ǌ�<��Bc�%p蝾�?�����N8-Z��{|��A�7C���;_=�i��M2���T��z�@�.~�y#'3��s�%f�;_ '�$�+��ʣT���<�]��`V�UCn�u�엞
Z�"i�
F��m��>Xʛ�\���׀�p�s��n0�pQ WƑz��Z=("԰��㧅PW<J�x��o:\�ר�!T�M�CĦ��!ߦ������Q��&Y�94��~7��8����N"�>�_��.��z1����ET�v.koa��0�ŵF����g�]��S�/H�(�IdQ�ǔ����Q,G �7�y����&.���zƫ�XT��.2���>�1l�ϒѯu�1���Bn��ʩaL��h���Jg�������S�~�j��A<��ŗ��!�DϪ��ٚcNPD�,[Z#���Q�=��5umʝ6��[��A��h��.~;L7�G�%8}6v7����*�ǁpv����_��=�{���X3&�La�=!�]�JY���/Q�~���J���H��o��ʓ
��KyN���a{ ��<����*be2qI�͹
�}_ǆ;#��B薳��D<��(�#;��Z<~�E�H������taӔ��'�vP?�gq���a<�Z�h�0���~j�DS������l?%�nB=�8r]S��]��0S�0L#�h�,C��>��}�sbE%��F6�v�S&�2�v��W.b��޺"fշ)x
�MS��V�@�g��)Ū{ß�۠���u�ܝ3��M���me��:|
��ט^��˧#K*���w4us͈�^�[�)Lфq�ƌ�>���[|m�F�g�"]���9��|�L����*O"o^��	8. A��[���̎���&�pI=7c��]��� 	���Ϟ��]�է���(q�o=>ۑ� |�T��p�Fn�����.|�gٶ�4g�.��H�א�2{�E�5���j	ҹ7H� ��:�K��6�ĭ,�H�):�2W��q��Dp���ǣ!�=�kN����eE��b�?K�]Ӭc��?ڱ܊�I�zX^7�9C_��5���E&�AT%���%��O��r�z�l��?�Bi!e�2�#Ҧ,��±ݐ��XŊ��t3k=ĵ~��Uﾍ���%aՅ��H/2S��$0P����#��B��>-��W ��uIɎ4�8���m1�tθ��yhR0IP�f�1"�����,u�K4�s j=�}�8���ȫ6�RT�Dr[X��ȴظ�����E��G�Ó�vR����(pӵ g$9־�:����Ōy܉�p��[O�8�E�7U�!�T�7��``��G�w��w7n~��?��c���(S|l���"k6H��(Wy�D�h��_�z��Q�Vxr� }3}�Mo�U0V��omS����-����/[!��!o�C�O4���ű�
`C�Y���m��Ƴ�U�g<���|��dK Uj�L��14����8JI���։A��4�A����}F�F�=]�s�+�;1�ʔ�-�V"���40�����h'2��_%���d��1])zU�8k�㟡=�@�-�����w��:z�>���'I�q�šv�Ґz 'c��'MQ4�� ���D�)�N@��W��s�������x����xhAe�N����=�m0y��n��c��.VBU\0�*]�G����*2�ṙ��ZW9{����1�������N��'��_�[N�i%�o��D�-N���2 fw�R������[_���F�(��&[�\^���	��E��)k]>�S�{H�?w�+�0X;�V�s3'^lu-OX׻w������F��rr�zu�\���u�H�+��Z� ����c:TG_>Xƃ�#>CP��Sd�j�3(BU���rp�U��6�r�h�'C�����Н��_5[<}vs���.��P"<����xct�h2B��R��B�&�5��79������|����x�)�p�]}`%N����&�(|�4|��/.�C��(���7X��
y�"i-(���w�L�/���GdC�+�+u�J��ZIğ�G��)A�ǒ��m�Ҙ�l�����B��O^�~hShOŠ������J�#�Ww������V������t���w��P�]O ���B�ы���%���U}�����՚���Zar@�0u,�E�Z��v��RT�FU���E���~u�uRN���'���b%QO�rw#��ɱ>i*��i����j�E}G���o�P����R@�_8*���su��;���IU�蜰yl��$����a"̈3��p�A<�7���:��՞��>�]g���������l~��I����;��,�FGu3)������dmh$��g�~�[�a��菂�&��bI�ZM:|�S3��8��H����q����!h��hS2�x���e�c�]x�����4t_b&O��yLdf�}�}?�n�2�5��1�	U�:w���	��|<z�w�6���>�ej1��������b�mڿ����j�Wb�3��W
�c�����RPf��J��PY�L�I��I��]H����c���/��{%�3B���W��p{#A�l�ָ/wY�:HB���<h����L�5��osZX�q��z�H%�8���i/����:|�q~Ep��M��i&/9Q�:�k�J�|�WD��&-��������
�d|n�����SP���q�F�PH�����_1��e�J��������v.��h���t�P-�T<�P��(2V%Dy�*�)�u����
������o�⒘�̏B�&R�>�U�� ���7��	n��b�_��3Λ��3��8��G≾;߾���ȳ;�폕M��V��&D�F�w�m��LMT�c
�����i��أ�Hu�^ى��}J�B=��k� ���/�$�b���J������C��&��l1�D�,m[�ss���q�zJ��堀X�${T�ь��N��{��싴?읐�s�
�A7n�]�j.h�ąy�=�P�8���j����|?PPI��gs�����"�~[��#^��C=��˽FKp+@��$ĂA?\F��2�MĔ ]�hȧnc\]������n����3��`�B���/G�fT22~*'/X��bJGCL�qbVp'H�x~|u���Y�A���0h� ��`	=�>ZʶP��V����{��n�����HI��Cţ�~ea�;9Rv�^Hn�����n��"�.��������|H�?ɬ��\���L�'8q�ɽ�Κ�0��A����z�J"�lfF�����2Ts�M�M��wĚ��n/���	v�h�k��S�x�HV���$��2�᤬s�v� ax�E�ɮ��V |��*yn�J��/d�j_�>q�\J�g8T~�9��[C�d���7�+�rd��p!���Q�� �jOw���c������I�����\<�Y��3����Ŧ;����� ���H���6kYh�����p�&P�"�EI�`E���}���������y�EL�n�'e�:�D=2
	��U��3���| 唐��!vb,������1Yҍ0�yRj�gO ���π�GBT�h�e��oL���V��}�Ik Wa��"S2��_�p��s��ޗ腍a�eƫ1s�R����0���#����Z6�W�1�y_(�>��I������]���w�+hoN��O@��Y�s�D�%s��>B	�X;�"x��L����=������0$��H��s�piǻ5g�I$�h����(1	V]/67��~��ڡ�U���*�����;����ӬߑU�E�i;�v�fGz d��5n8�Q���݉�-�ɨ������ڀ�Y���4��;����#� M��c��(�z���l����
�h�Dp)L�%#�Y�l;��6���A&Gt�&����JTũ;��
�����Lq`��$�a�_� �-�9 [<=�� ��9�2=�>@�v�*�R�/�pP��PY��r��`��n�RQ� ��� �6s���+
%}f�cf���vb�eH�{��S,�wZSs9U�sP���A��u��|��R��z�h���JQer�kW}&�+ݛ�K�s���FvJ��B�8�w��g�ˏ\�gӭy�T��c�~9���{�b)��:_{(Pa�[��H&赌�N����B��9_M'�����~n�طߴ`V�kRa��9 H�&Hhq0fT�|1�����T1i�/�(y�'��^�e��M�Hf�;���3����Z(#��fP��l-Oa�70��=���'�˗�W���E,L�S��f%npK�̶�\L̗�v��dJ��r=w[G��KT7�w����[c�)��K�]�,Ò��|%0��k�Sl��Wq��&¶u�;��H��"�@]>����H0~�l������h��|<姽w���
=B��p%����P[��wΒ��4�T�E/D��?@����5AΝ��@����#8��K����SD*�k��T��:�F�!_����Y>�H�eK�H�9*�������.��4;�L{�-g��ͅ$�u|#��ڎFOo��O�ӧ��<<a�=�ژs@%�la���J�g���V��1"��5����m���=��������o ^�r��$xG��'@{Sֆ�*��ܰm�c�b�0�X���������R�>Ӊþ��#�|�k���q#���XJ�v��B[�v5�q[���I��^�з<���D��Gw�����қK�'u�}T������`A�}�J��{��¿��6�bA#r�}�]R���VD
���y��j��Q��N�"�?�@�a�	�\�n�����Ӝ6�5ӓ=��g3�,�����Փ�_��R�3���E�9B����$��%�^�P�\7Ϭt�x�x*?VU�����O�rgRM�X���s�O�(���9����@_�+*��ӧ!`B	L��	O�@P���wܞ@���R읩��)��}�4Y D�/a���;���cJ\�� Lf�o�%�����ZIv���f��s���I��Jm{�c�W݁�0��s&��a��	�w��e�(��TDK+�X��p����$Lg]fl	��;o�t�GP�*B�os����żp�-����f]��Y=o��t+G�ǹ�9`�-��f�$PU�܏=�9�
�ݷY����}��΃j�� j��a���߭�a8��!�y�~,_���w`W����7���T��T�N�`h�2n��TMxF���-��R��:Fx<f̔��7�?���3��$�_�����2��U�" :�����iO��I�ݗb�u��������?[�s�H�"%2#�f�b�y2��^�H��DHxj)�8�su7�����9�Vゆ�q��8�j�,����l'Š��
�Mt�~oK.�`8�A2���\�{`Ix�H��4){��H(�r\�^��_�$�b�L� ��~�W"
�L�W4�퀔�I�W
�(UI1���x�;���6]�]��}n2�&ME���W[������#���7�WyY�T,��qY>����%��)a��4��d7�ˊ�#���'�Pd�����xSt9M�V�0�h՝ڨӅN-TR̓��c �As�����^�ᅶ*2u_�n�%��	9哇�w1K������i�vq&RG����Y�h#�Ŋx���J�ם��.�f�jI�i+�K`e�JEbbv�:�o�f��<���!���������6nA�:�|����g}�1�G��݊�[��}�%
EF��K0Ljd���[�͡[�>X���M����2����Z�n�����tkb? �E�t���1*��w��4x��%bP�~
��lW.��R�-gJa�v��}��� ���	{	�HYݡ���1��l4)b����q���5�RJ�w���'ă���9�xsƇD��~5��3�n�����*�;��� u��9��(T��+�Y[I��'� �Ԫ��N1W�� �R_�����j�)d��8���+���^�h�+���϶`��ĉB�a�X0p����-9j���t�T^��q�v[6\7�{����RO��&,^��,�����@]6�b��}Q�#�>o�v��?I�P3����[3����?8�,O ݘ���4��g ��[Z�1̑��ߎ��-���(MOꡁ����]��j�ѵ��q٣/��XҬ᎘$9]�A�������M	H�'�oWB~�e}
�;�X���㻬V��e(E\	Q���Pq��/��W3pY�����m��A��T�Ck5�i�ң�N��k0��!�2O�YX
�1�*�����l?�lQ-�nߞ��
�����C���>�\��E����x��y�1Ydqo�s������\�p�ȕkL�L8̬�ZRu�K˨�Q;T�܂C���u�ƭ���dI,�	��$�W���Qp_.�;`��n�h��;n�d����}̊/��<}q"��B���p�����*����,1X{x�gB2-f����y�˰��Wj�[͍�l�<��u�,]^[|��� �!$����ͱ2A�K�C8)7B$'t�(z�!#2�'>q5��~�7����nq�5��Ѓ ��d��K^v����<N���8QP��@'T�-���wEr��� [���Ҏ�N��kw�?��$��kjZ��N��ݯKh󗙿L��ֵmx���$�������`�zȩ+�v�8�A��W��=��c� mD�R�l��D���T��y�:����m6��/���P�nl/�z��W��߱Qܫ��X�|��,ץ��̭�J�� �|�$���Gے�+SWj���6��`��p����8���k��@TD*6c������.f_�L��R���Z��8D�d����%���ݠ��K�J�MR:Ȱ+�R3�|xs���s�����-�:��Q���"�ic���B�@���7�;�p�ɂ�j;�pa��>�J������9�7�jꓖ�O��}ԧ"�([�BՅ7�fh�1��F>���s��/�mT9xlє��u��ly��RAW3�d �uq�@�Nw�[Sw�ӫд���G��B(����M��\�`#�΂�\a������h���dy ���蠩�*�pl�?�;��@"�3c;���ӯ$��M�b�wGp��t$>0��_�+�g/(���3�����#Ŷ���Cy��|EG=���O3�@q��?�_g��)��w�-�W�@Rx�AW�IϪ�6�|����z�S�&J��AYhDy�oD��<�G��Y¾�)�)!�?�3מ�3�3Mg�\��ۉ�0��6�Ё�z윱�m�\y��e�Q˴�︳�>�W�9S���9�,U2�k7��1t��	5Ԍi�Q#�\�c]njF=��Tӳ��5,t��_�8�_�*s$M���۫ Ƭp�v����Ef�.	Ĵ��椐J2,�g��+�ƥ�����+k� JZ��-X�ɧ�^^2�(p���(��A�
M�S��I��������$���
A���/�yW��кҫLx�ɼ��LQ:��9�a;i���T�/)_�2�7���)޵��ub�g�C�; /��M��yXx�+ևF��$�@W��F�јP�1�������&�r"%����L�|��(ea���᳓6��GN��9J]�
� 'i5�-߫��2e����tX��5E��������e
Zq��6R>���!~�ϧ"	ɚk�����`E,��7e��Ү)�wĐ�>Ru�*$E��E�	:Q6�h�a�Gmӥt�Y��|t�O��\L7�#�@�ů�x��������u��)J�E�q�{۽���Fg��b�֣����'��1Ng���� E����� #��n ����O^b�V?KI�6p[c0��տ�W�&
��E{Z�����F�Oz��p~�s�����
vp��W�ڇ�:�ۺ����T\�����ڗѪ�:fT�7,wčQ"?Vq0���Rxގ��WN��������v��P��X��p:�i���q���{���(�:X	K9L3sQ	Z��#��o�RlZ[nZ��� 56w�&C��H�^C�ՕtO��=�UZ�9�B��(�N�������5��T-`՗>�DM�+�B��R�L��֬����ؤL�e�1u�r����z�����B�p�y9�����X���kB��2 ��e���S���&(_L���`�5(��Ν�o�%�	�rS��7�A����T�_
���b��4�_]� z��ټ���nYt��H����R=��7�#�)���Lm��П���~S�����䯳���z1����NR�C�7�^�dp�tY�5� ��O��m��~�Y�LU^8���C��|'�3�)H�N������qa�K0�O��̣wGxS݇;�̴bL�k �
,,
�5�ʩ�G�2�H��ņ���e �i�.��C�j�z���0O3�&=PJ�S%Us�S�K�mM�}�����t=R�~� M9]D���!��
4)� q}�͆��H���U��Wm�
�+����O+ �q�oc�W�� �(,&�+	��;�A�}����%\E�9|���G���yHm]n�<	�l<_V�n�=|���P���`�R���,�%&u�m&� 1
���T�G9ܗ	�ؽ��o>�Rn$y���=@D�Aq�v�U�E8ٙădp�)�_���`46���sK1�<�r/�!��v`���h]�.�Ւn�("����cs?+��{�૾.�ܦt�@;L��Z/�.[T7�r�pF������p���Z��-�˚�ეΎ�1+E�7��z����Y/of8��&O�M��_�FŒ����z��T�x�ߡ`����D>�^sm"�gJ�?�$�+�΁�_�oS�7�ǡ`���F�c�xǇ;O�W�o���$h�-�O�T�	r���6	���� &F*Ul�^� ��8���ޖ"r���}˓
������0��6�D��v�?�6��� �:��mo;/:�⸵�G
�K�N8eW�C�����ޣ����:�÷a�������[ ��4r)��ɺ��M�L��!5"ܻ��IY-&V���J����N�T, �dgհ��F��=�r'�EM�]�R)��P�N�����*���+[I{T<u�}����'TS�[WA��(�ve�hOy�篩�b忭�R���m7�*1��m���kQ���K�s�?�{6�'F�^�\�
��o�Flr%�S]����w�&�I�_� .N]���~;��pjͶ9��ײ�Ԥ�V f�ٚJ-A�Z(�_��m�@��^*a���ַ!�	��Q�ah��Q�t�1�|O� ����(/�%?�qN�
����-G1q��F�^���*ggD��.��ԁ4G�6}�AmkkO�a��^V���g�i���TA��|���)��C&_#4����~4{�����-7US��[�M�"��T(䝾D^�]b%�،�r�����=L;�O*3v"^�dPj�<b@�scm���c�|�EOk�ؓf�����_(q��dP\5���B1���^Z|X�|\k�m�<>`Oq����0��0>ުU����O{��O-���f� BdF^�<���fQU׋��1�%{�y����J7�J�^�1kOA�jh��˜�����j��~vr*��Q����/h>�x<��#q���m4�2d�O�I��e�?��E�g@�Sc�P��$�b&4X�V�A<�`��Qm��A}`��b��bY�M~JT� ;� |�/�z��2W��T4�8�7J2j��h�lE�Y��6���KL7(��@����~/���Aoi�v�r����&��a�K���E��1�i�Ҳ�s#���br�hګ�Q�M���kN���)2&(�'4�4$ia@���`\w�hP}��W\ ]���اmg�*���˵��?Ub �i���baD�i����c��[n�����C7��k�78 �?���˟@{�Ge���(�,��/3�G BvR!�Ac�	u�Z3��7yk?4bI@���g��zV���}AŪ�=C����H9��4L#q�*�7�;$���d��K�섞��"+c����Ąٺ�۸�i^�)�w���-K�6�xȮ�h�zxy�-�k���u�k7�Fd�S�63`�����}���5kH���η�44c"#B��X�@�>����`��fB-����D�:*�8{r]�y� �BI����*MW��A���d��#W&���
v`P��~�e@NA��J$x��}�⼦���|j�N ɲ�B��au� /���:.�(G��G-��P��,Z�3�/��G�����"~�>�����)~Eg_�m� eCh���a���8뵽������^�_��BB&�[��L߸
�� )��
ώ�_%�-�������_%&h5����~CRG���>J��<�a��NG��5�aib2'���R�%%0|7��%jy!���$��F�%�7og;�s<�XtVΏ6��Wţ��3�
k����@c���FVp���Ի�:�f(����buAm�1�u�xD���u�)�D���� DK�'3.���U���i��(M�WA�%����Um����7c�_��F#�Kўp�u��\���7y�s����O������,J��=�!`89��-��z���0��KFK�R�v��w�c�L~�M-.H��^��m�ITw����_?3~%b�U�fs_�U�Tj���׬'���ZZ��]���s�Y	��dP�|�|,�� A}�J.}�s��|Yn_R���J�	��`M�cf$fv8B?i�[�:�:U7zȋY��ݾ�+D�q튏�����i\O̓��s�H1���
5Ǩv(o���b-ܜ���� ?��B�b(�7�� �
;֥�Ŝ����c���8�('<���͇3&��?
$������=?@�Ū.�W
�L�T�=����`�pw���:��c����M(�Pp;4j������g&��j.�ːyoEg(5�X�T�~s�6F���l����/a��͑S�Q�����B��y�}#z�f07�K�,�A�?bv�ҍ�?�Pӏ��k�r3���{A�����/���?��$����HO�*���gB�+�_�����{ƨg0�3P�
Yh6-���R�\)%�/��t#�C�c����j�S��U#9��c�P0�)ؐ�!�\X�}9.f��ԡ�o�~P���m��*����u�rD^8`l�r1.��P��d3җ"��V����:��ό�����S�͆_���D���,��>�yM���L���S%����{-��Y���v�3/;��BrJ]栎}�c1ܪIPݪTW����離Uj	����mXGq|����6k�ȧ܅6ߵ��>}���P=@�籜U*l�b,A��zc`��4���{�:���m�ST\���]�^�e�ل������MQܧ��S����J$L�Ǵ��,1���Yt.�*k���j�C�en2ĥ��4�5wJpqۛVv��3f㓥���r)hlE��������.��c�7+���k�o�
�ԩ,�K"[�늶�T(1!E^l��1�iT�c���o�ж�$����<�rwE3U��Ð^>	�ܭ�y�@)�4�RT=���� $�`����*���HB��h�Xs���PFl�=�W;����� Y�y�R?x��$���H��@��ۦ��e04��t�����(E|�Ӂw��.U��F���n�"A�`V����`��	�Ğp,�i��k�Ck�I�^���7����z|��aLyGy�z��^,��l�#����!F,���g-B]��I��i+��	Z�	���:)TOl�,m�2H�A^�TT�@�����Um͔�6͙�ZK��h�e[� �N��{��lQ��B;L[:t���pAC��;s)*���+2�~?��h�8喚t���i�}V9Gx3��g����gI�$��Y�ڠHB7k>�9E՘�娙3���> Y>��V�Im��o�Ɏ��)�~�Z%M$B-`:O[�E%U
���=w��zI�	��H�+�e�(����
�s+�f�S�1^�s]_���T���w4�&_����EM�3�Z�>iҗf,�i��E�����+�<c����CJ��ѳ��
���r¯�z��X�bt������鷕�;�o1��XV�L��������i�m�PӑH��3��"#2�(�ߋ�	O��D���&+�܅p�+!i�?��M:r���u7�T�b]Z�Tن�4�E���8k��}ݶ'͟�ƚlHt�1��Ť�b��M� �0�s�Y����v��5��\ScZ��K����F�#��6�m��K/��$�8��EO��!��G+Y��<ZyMz#8�;��	��.�<~�	����Q�	�'��4wp�5t�GC%��[�u�C�,�qs��j��C ʦl�l�?2@${� 4?%�8<�5X�UhMH^{w-���B��X�\�I������C� H ��(�ɌL=j5u�P�Ѯ�ݾ�_d5�,�܋S%E�'��� �T�|n?�7Ɏ���£�lhNL���*��������NzD��Ű���g���<%KN
Lܕ]|�Zޑ�n��yW�H3��J�R/�O�Q,j�W�?�g�sNΎ�GT\^@Vj4`��XQLl�o�q�����f�3�ĉ�N���q���W�iĴѵJu�
��e�r�Mz0;�oԲ�16�|X�A����(��4�bgj�)O��*��������D6��3��B�ƔN�������m�H���,�;��f8�-5�x���ap����
T��DUk�ǒZ���<!^r�0�.ώ _�|��%Jp���ͤľu�wX�$��/@>O"�,�n���J��!Gْ���r*�c���c���e�4:f�FX�/٠�P&(ʶ�]SH��@�g1w/��-Yh뽛�X��:�Q�Cd��x��T�1vM�7�oK�l��׾Y�fQ���l�۷󂆷��3M��0����+�g��������Yb\���R��!S偍����Ys;���Tl�aj�7�$ 1��b�]h�A�.���-�)���:�#vƵ�."��gE�Y�.Jx��)�f�a�r}�᡻k��th�`C	.IlOU��jD���|�U�)}5�1L���?̦��P�eE3��j�	Y��з_lè����̶7��~n�	y1<�ɬN�t�h^ �@�o
{�x�������fC�P閸)K�bTɮ�\@6Y�}u5��Vٍ�Y����Ñ��C��heX/�����:���x���EG���Q�g�q��sή�ѯ�n%��/Y������g��|_���!����c
�QZ��A��!Գ�q~���k�w�N��
���_��P��~d�;hS���b-y�n���A�( n�0&;�(p�SI�Ƀ*hV�7Mډٻ��1Th1�����Q�C	0%Yб��.�͖��-�M�}_���V�d�pϣQIz��2!��/��8�'��t4��CūO:�*`�Z%*f�߬��"����t�<���������"N2-�6)w)�2����u[7��M��1�m2첢�O�1��@�6�*���_z)����(�i�R	eW��BR��b'�!b+�� ����9�;x�o���G)O�����| ��5#kD�p�Z�|ɜx�ټʊE���Әu\[� �'���L������4�\�W�#�վ�$�������֍��IM�l��]%^�~�:Q�������Ӝ߂�Vq���Gw@��E���Ip��]U�5�����p�����AAZ!|���zg適�X��%����;�Z B��	��������������Q��Sm���X�%�G��|�Ǣ��5�v�8�z\q���ob��� �r
f������͍E,���lğ��C+E��:V�Нq"�YF�CaQ$�NIT���vW�;���Y��|���Mt��Y�{_`	�;��Զ5�ʼ+>����bT@&Gl!/A�̱ye$�b�Y��p'���%w=c�yG�W�Uz��"Λ�K��N���&5#]�m����$.�ڡ����/��AR���j키��i�yD��@�V�_�_���P����7H���hÌ�ڟ�~�л'}�^E�Ao�Ԕs���IB��i�Sb��VA�V�Km��R���fK�v�B�����Kx�zywN�C6̀^�u8�!�4�=��m�$��y�T�hG<���otZY������n�!��#�M�L�y�HypI��$!�R&��aU+���〱��2WAG���{(W��S5�K� ����	�s�^b�ڣ}�^<����ԍ�:b��h�F��4
r��Э�<��
�)�E}�ޔ5���r�d����f���~�����(����2]窔E���J�]�in�+bߢ!�p��:"��56D~��[�9]O��Ʈ�K+��=����0��D �o����R�`�ۏ�HǙ������g"�v�$L�7�\u������x������K�F,NW|I8��p����XV�ĊoA�Na$b�5�����=���+w�)�;�R\�J����._E-�ϲ
q�DmI^�t(�����`�NECH��$$�6�r����$5Z��_x�c_�i�;��*�D0��/�w��	X?[�6�q|�P��gn��g���������N�I��ꏝ<��y�����3B�,�Ȏn �R#0��_�-��R���@�d�����f�[�����a(�Ĝ/)=���g��}���	���1�m:n��yCg048��ltd�=7?�,
mYX���A�WyQke�P�f���XE��~���5E��@#f�-oQ؎r���rP�ֽJ�`��D�.�!�
iKZ]Ҳb��t	˒o1�.uD��H�BF���PK�]�Z�03g*��N�T�h�x\N7�^��H?il
7e�o`B���h��Ħ�{�h���.㢗�<S�q%=����oy�Bx�|�mX��d�J�%�zv��v���롂iE0~�w�J��I�3ԛ/=�<�q߳W����?�p;K��ˉ���B�܎Ƨ����s�k�ʯ�O�k���9TH�� ��WȰ����S���,��%5>��� r��QC�2����k��ݲ6>����H� ��t�}˒�}^a���P�
&�"'�v\���ڒ�\�^T���r�q�WB�#|��+.�o��k�<�&�
G-�3��\���֗�`��"�~��ԭ�b�������"Z��l�&U���`  �\a=Jv���)�˞V٬�����#�;goi9�﨟��?V ������G�v��'��U�����t]e� �3O_J<S�9.�>����p��+v�{�P��~�W!D������l�	*?l��n�u\D���2)rL���ł�Ri�d�5�9@�ϼ]��Ҋ��.����
�����^�qT)���SQ�3~�	,�����}�����6�x�f��Cl�WG�('��m���XIs]sDW̷�8������_E�ȏ�b����(;@D�x����w(Z��sA�
I!���!�"H��~�6؏�t�_��p$��A�C(b�O�A��D(�q\���P!�q
潗���,�N��𻴴<⣯w��;F�28e�N�����3�#�(�l�z����x�q�B�,�Fb\�b(�/����^��O=�G�L��dꃯc�R䐅�ݓyW7i�Hw0����'yC�F f|ȴ ��J���a��uӭ̱�k̸HP�I���W��i��
�Vf̠w�1�`�w:�w�,a���M�1�TY.�*Һ��?��L�T��E�״��ל-��.=͟-���J/��K�"`�3���O��)��蝯��$�Z���y�%�C�]��j
��A��gH]6�I;�P��b�e��[X*�*�/�I���G�
��_P��GB U]k���3��ܖ��1��<W4Ggʑ��Wk���(�iO�K|Ə��<B�b�����0�F��DK] ���:�f�<�i����_��� ��������`i�'��x���c���^�BƆ�Q��K�(z�V�M&۱���
���(0!�� $�я��,G�vuPʑ��u���Ûo1?un3	�|��tɖ�2���i����V�������1lkPN䉐� ��4�M��)0��4]78jj��6ō��VWN�e�7s�S^X�l��)��.<��bA[���~*���$�~��9mț�
]�p?v-{M��<��q��ZR3b
]���JC�> �FJ4�eMA�� ��1-���t���_�7��A��[�/�(U�lR����}0~�N���O�[Ԡ/�몄����H��cz܁3��'�?'��=+_$��W��or���7A��W��E5=؊���Rt�>0��@I?u�FWO~����{g\����Ɗú����dh�K����1{>9����䡨c�?pJ�I<�����k�h�������P���2<��l�nR������:���I��2h��Z`..
��X��.0�& Yp���"+�����PܥZ�:���4?��)�i�Q58=��l�ި�<w�����5#5��R=p�I�C��4�O���Ȟ,�əj���!Q�5.��G��5
h�^��(!t��˵|;+K��b����W�6C#���1SK�%E�ˮ�xi���!N��zw��������
E�!�em��OM�#��*��?++׈�D.߻�O����z�:�7���142���>��2�}K�T�x�%�=M��˺�B�sɖ�5�jF������� ~��ҽæm��C�qF��][�+F����U�_��T�u/���ɩĒe�`�3CeSi��qG�]���|x��w8	��@���8��p�����[�m��7�P�S9�v�Y��ʁA�f����J�����y5mc���i����v��K3�ҧ<M�m����G*��!�S�]%��t��ۨ���㩆F�?x:]e��sI?~�3I�lMp���ݣ��?��A��J�I(���ɝ������� �`w�N���ʯIJD��V��}�V_�2
�[�A��i띇�bF9�܈���|V	�1�h�}'*�-̼֡��f�^���02;K�����*zǶ�^���&<��1��o{�;�w�m:��������0�c-��_�y.����� 쳍��Wa�,�$H��}}�c$SϏ��)��iyt?���~5Q����o�}���y��a��'/�w�T�=VZQ��Y�t��5�����y���Hi����ԋf�0E�al_�[u����S:e�"�&�A,+���/��v����>����W���s(Yh�FT�s~~��)�*L�������gc�z
ΜV���RVng���k�*$�a�Йٵ��?4%����&�:Q�G�Ǖ~ag��z��|���Aڰ���A04l��T��	� ����Isӌא��+��Y�^ډ�T��̼)X�Os���'|s���+�S�fn���x�b�	|��=�$c%	����o
�X�tR�N����ge�4�I=���!�ƈ��v��%���.>���h�^�10��ݸn5�[d�YW���6y&��-�gL�3
�R" ��o�5��y_���o&>�=��9ڰ|�ߝ��F��4_�P�0Z�z�� g�
�z�q���葙$A�M����u��B	;8+cd��~/�4�x�9g��8�C�2E>�����hJ#U�.P^�D&C�d'�]��Xeq��>��p���ӄPQ��mG]�}�9F�PxX�i��%��P��: ����K~��'����`����]8*"�����Tw�]��[�[ï�'�5:��vc`�n|>������4��1�<�3��9�:����ȇ�FT�� S�>���
�2���S�g��N�	��.�-7��f�'��+�x7b���-�v[Ξ7�/�2��PR��P�@
x����^��v7&YC�!�6ky|q=ə���yt�/#K���t���~�G ʠ;[�r�#(]D�Q���E.��v Vk�)ld~�y���m�z��Wy�F���8�./���c�¯��b�	Mс=%:�/�A�U!�y.7�tI�d\� �ҚG��O$7���r���~���_��j��<��w��"y�B�0Sݜǝ�JŒ፥�X�j�F���A��4�1��d�t<��;��q�X�~N�&XT�Wt1�'��6's�LefQ�U(r��������v"��GD `V���T���f�s��}w�D=U>H��m�	)V~֥>���23�WG�P5(�2�)�[g����l}RwU<���9��=�������0Z�����*�K� 6}Y�V�	�}��DPj�[p�����aԔ�8�����@]4��k�v�aW�' ��F�z�wx"=y�s���Q>��V��[ܬ�}�S�\q���_4��B&��rzF�����bT&[xM�G>iy�r ���N�͖�j��Vd��@^��<�s:|�*X/߷蹚����M��=�4k(��'�����ũ�($C�`���旔Ḟ(h����񄢴o�����W������6����d����@S��9�6S���s��oNe�0�F�;�Z�nKV�CQsq�Ǩ7E�{�"k1���G�O$����1���3�_H'옒2����[�����{+�X������aIL���W�עє���,V�2�6��VDU�zd]?���>8�_R�A= y�D	NY���&����K����Kn>���k1�yr]��3�ro�/�?���F��-k���J�CI�c��%`Jӂ�3cV�Wo?��n��8(2�՘k��4�͠�Ɍdd�sLu�������{�
�!o�\sa�F5T����u��P%8D�| ���#~���ɫO$�� yqk�����~��@-m�v�n��:��?���y�F�k�IZ�<5��:#`:��ś���ٜ������2���"��K9`ƈA�Z\Vn�#g��O���YP<��3���KW�[r-_<N:	�O��X���T�ԁ���Ѿ�&���n���l:)@ �A3rL3XG�6�ښ`�8mF˟��~QB� ,:g�̦x�9'm&.Gd�����ď���� S0uhQ5����)o��P��$#�� �a�� v�|�M�����s֟�hpTvp���[I��+/B���@�ĚΛ�o���=\�o��)5_~�r�X�:�Y;��.pp���4wd9߇��>��lOT�\�]EM��U�,f\�H���Tw��V^UB����BO,�&M:����
�y.g/�j��M8�� xW�IF��qz4[[>g��#�����ۑ���t�ث��T��^ �$�뮴�JM����kL���;H}!r{������57�I���6�'=(����e,b�.n�+W�n׷��g�����܉ʷ/�,;`G��!��{��Q�(�!U�MS�!���"Q�<8�F���>m0�)(�Ԋ�$�ɽ50v�F9u�\y/��Noz��@u�x$Y'���'a��u����3be���ҏ���Sߠ���8�􊦤R��
�q�:��އ*R��SB�V�Zi��]�{�n��ܪ�Ơ��!�jMƈ�-ҵ{��>����u�9����Ȭ�B?��ec`�2��p ������HO�w�~�x>����N(��A�1ֱI(�Yx�[.��Hl��|���pL �LYT����	�;�,U�(h>��(cVN}r�?� ��jN��ܬ^wc\*�2.�tJ�R��ly)ڔ\��}#�BvO\�2c��m��J6�_ϯ��\�r�����|=�rCj|�B�a�A�PJe��� �+lF��,+mGV�����Vj���(r�'�u��>���:U7/Z&�üS�JRa�Wa�[WgEw\5^�P#��{�öm����o��y"� �"E�:,�>�>tTw�q����k�K�4[����F�H�X�e����a˿��m��4��d��+��p�����-��(�v�8��h 	7��2=9��~mf�0Y�����#�A����l~�\
`N!3��[��3Kil�*�	=����u�)�%1�󔅶sm׬B��g��!{̱D�r�&c�q#��:�t�l^
�DY��p��ofx�6q�*x�)��L���/%*�E*�-���|�0�>�z��S@I� ��݂�
�R��ټ����j!��@�����3u�ǼBT5�(�b��o��JH�n2��[4�v'7e�?���� �҄��E��f<�:סd9x#+ �#���T��b�N���C0�ɉSD�?
��d�@��<)�ǁA@��5���1�>'jfJJ�a�ez* }j��w<�t�N�0Ƶ�����n6��/]N�@�~��$t90u�`�T���:y�H��H!s���K��?|$���?Yѻ����+A�.�X��Kz����L��fœ�MLm���!P�8�C��̈�h6;��в����&��Tj�z��`_�6*�s�}�aQ��v]�@Y��|b��@<���x����,��}Tv��i��V��瀾%`��H���`�?;�_Vb`ޝk�Xn���Y�8v�K�����5�Z����*, �laeƤ�s��|n,j�\��X�k�����9����P���8H�DJ.���f��BkqTgAQ�{@�H���$�/�����x4�W*�Ћ��I���C��Iw�i�jz�^A��Y�s��Dַs]�X$|��g�l�t�]1�*��+�<e�ͫAw%��1
�>3�f�g�X�q���P#ifw�^�К�KO�y��
,���tG	DZ��uw�H
���ڮQ�,Ǚ�	��/�1�����]��ۡ�a�[�>D> �+_-л!2�QCOgv�ŕ�c3HO�u�?�i�e��	��(�%�4&k\q�*l%��W��R��
0G��ўڑ츌W���(�ۋ��0�-#G�6{ݞ�2\�PHNV�Io !�������c ���ҋ��*����m��s�_k�]-��@ ��l�I}/�G��ك��mR� 횴�Z}��XB�	J�v����~e��|��:�3����G�7"g���o�f��Ï��Тu�й�IRJ�	���RY�T�K�é-Ô�ֳ�%��Z�7��YߤŒ�����0�)�b�H��C+��4`�z�LֻU_�Ƀ�Ĺ�Pٮ�V$[s�Ʃ`��*w��kM�9(J7��H��.����F((!�x�g[�_���߭��<��hbƈk�i��rra�Ϣ`����C�^��Sq�)��&ʩU�#��1� �t�ʇ���%�{���b1�ơ��Sc��d��W��WC1��/�^ � ������/�����vpc�qAԑ�i�ݓ�����@����Nt��O�>�*�Ղ���\-�Nea�eI�e��THLU]�6[�o0�f� ɾ�����Fc�;P�k�a�q�G�>�p�BӇ���9W��(Ѯ�zJ�y���Xsl��Y*��,��d�l��a���t�b�o�o�Z���@OA��jiA�[��f�ab����x4B�Y���}�r6	
�dއ���P>��حsA���[Ʌ�_�Y4$�zvn� �4W>���j�@�E9s�I�q���X��J��>��
3X�ڻ���T�ڣj�"�����W?ہ ��)�s�Ï\-��0���3�A�P��qe��������HmJF8�#�&Z���=�'O[��V0Z��fE�\�ޣj�`6'�G�N�-��uƌ�D���+��\�bl_��h�`��^�=e)�����I����z��'�V�\o��l֋qU����Z��HAꎫ.��OK��.P����/@D�*.�{j�Z&K�R"ȌW<z$Uw��W�|2��Q���%��,�_�{0�>�V����.����K$�/�8����5uL�mb����G]�ѽ����3H&��r���=O#��ū����h�7�C���%�A��1��C[��Z]+��I����̩�D��"��US<XZ�
㦩ѻo'\��ی��4�9�|�1O<�a)I�[��O�aimO��R{;l#���L����.��&�2��nR��}��а7I3umv|i������mZ���0v�̖�(#JQ�w �ID��� ӑ�k4�_�`�#���8s��|݅�<d�p���{�|��S�'o����8�s��GHU)�Ve��H�u���%��i��k?[�Z��B�����?M,�yR$oH~�5%�fB^����@6�r�B�ݲ:�WZk%�ē�Ki����{�
�ȡ�S	���	��rY@�j� �Ewt�2[ȣ��'Z<�{�8�|�Z�T7*��I�����Ӡ��9uOm����D�U������_�`�L��x��&�+ ݷ�4{�Ӭ�ö�i�Z���,�^���Z��	��DL� �1H*�͝��W�^/<"68�L;ڢ�S�5�|�\��V+���0��d��H��$��st{�?���ӄL4//:U�̩Vu�a�z���O� a6��3�`~���,��S�F�Ln��'>W�$F|b�,���h�34���J�F�ˬգ��p����{`��Om�&��l�'^�)ERv�fޢ*����n�?zL̆C�]��/4"z�l�g����H�;��S|�Pj�V�k���������N	�U*����pab-�Em7�;;7�'/I
4� N-���5'��D�)�d��U��pI?��<��"+��{�)*����f�@��7��bN[-8�["$�.��K�o��8fZ'��	�'�2
�u�%*����jـ5��8�,�sJ#!w�30���#�����R�� GB9�;�f�Sgf~g�)Q�wN�ڼ~	h���x*Ɛ���΍U&Պg����5�	�u��p[��21�mp'յ����J�L�xYI�G�/�xӼc֔ͧrƓ1�dݯ��Cue�s��>F��Iq��C��g��Ƃ'�0���^�d� ��-�bT�"]�B�)4u�}&��� �'�*.��<�iR��Gꃐ���f��]�v���9��k�"0�׌D)���y�+Ϫ�;}[�s
Q����R�oZ��H���mN�K�Ha�]O�-鐃����6���w����-O ����!�3��W���a����E�B�f`�-�����G�\)x�1f�J����σ����4�ҭ����b|Fd��Q���Y�Kӂ��b&@?񃾍��M�����ͱ�P"�6@;Wk�R�n �+-���zE�ۮ�RD�l_)~�Фw}>��Q��t��h��.�gG�H�W�AK㉇�ug&�f������Y����N����2c��Z��K��������k�g�+�w0���rv�
�w�p|��A��N��ڄ�m$>G���:���^a�ai�C�u�g�����#g[
��\�w�a'ُ2�o�Nu�L�=+�A�Z�E��m]Jۍ�0��N�<�v��7Я�D@��\�~�S1�y��N#�e��e�+GFƑ5c�I9O�Q�f|�Av������#����d��y��Ww\�����P[���q��	*h�F��c�-�SyQ�r�Vd{^DE[�	IH���	I7��3̡��#�VTԉ��P�TSuo;�p�~�*E5�g�λ��J����sOϕ�b^zJ��
G]׫���֯	ki��u杊�s�Z�
�) *}JO�]�=`�q--\���,���B���<�!}�wf�9^F�aK��%��a8�g�Y�]��cf)�1s���J�^�Ϡ�#\�+n�l	`X��r�&�Q坪G%I��k-ʄq��J���鑛��&ˏX��X�V���]y@�G���g�#��&�o=�'jBk�g��YC���o��d�bZv�F6�/v��w�������ף�R��O�]�j%�r��Үd��@�\�/�䟗��M�;`_��o~��W���B�}���6�D [f#f�9j^8���������ye���j9R}s�s���I��3�#ǀ���ˋ��5����=��C�!^D���t�S����jyZf�҃�:��#�Yf�bTw��G�S28�5���ϭ�0����v>�9�f������#
�P�%krρ�ЈfPKv�$��i�m#n_u1K2y��L���)cg޿��&�C2�PIT����惝���������Äk���ln�Z�r�@�+<g=�y39��������!鑝��aq�ڄ�k��n�1g���WI;�Rg�>�w:xk��?7{��>I{P`�T}�{t��J�:}z�̐F�^���<��%0���>�J��ԍ��h�eJ9}p��#,/��s�fMp� hd�?DT<]�'�p���:qbq[F���K�U0-�]y
�
��ai�[Q\�ڑ�A���S�]{z�3�p�uRM��? n���@��fSr�`�1����j���̳W��0�E` �L�SO��n*Vh�f��Cc*)?�OgSi͒����Y��y^��>���$=<�!�^)���ጠUm�?p|a��7\f/7�ߔ�H��J��Vc��T�փ��)*��<�7���b��B`G�ۋ�h�-0�M��Y3�("���}po��'�l��8�iﷱ�W<���i���p�����fS��/�Ջ�����L��6��ؾ��iwA���Mٔ`�b+��h�	^��
į�f��:���P� h|�h�}Ar������`٘��NKs�FǢw��$�&���� xB�7�0;-V�O�@��Ln`�̖>��N?�()�2�"~�w����	Q�<8���Gh���,����Qs�!x.�q�̬2��0_:����𥛒#L��6�������3��P��\���w��դ5�q�g��3���ơ���)x�Bg46�W�l{��~a��&���Cc����~^WveDf���C�@�mrrV�4;�j�T$�a�Z�!���UnB
)뺄cÍd�+��\%��JMdi�0V	ݔ��M�^Ǧ��f����ٹ���]�������}�V�b 7-�6��@��*0Zщ� �Ǎ뽱���z�kA�n�i*��V�č���&��H�|�;��cb���Ĉ��>��N߫�eZ+�;ɑx�Q�̸��^1��5���p��de�R<�����h�#���\ ��X%��@z���i�T�g�b��K.�*vZq��Kp��*,Z%R����Z'�])���Cv�ru9:h��Q����X�ws���P�*��t�/�sA;�',�t��H6�3�(6���h�����/q�x�*7�`�� ����Ò8oUM�%�=T�õ��r��0Ĩ�D����\,�EJN:l�n�����qQ�!��x_{D�ԷȆ`��<��X���������l�X�Q�"wv:�aT�Q
�8Cߩb���f���'d��Nff�=�6Zʏ�@&�K�8��+(�$�1l�����{��@�񣿭,���@D6��<c�����~�������Uު����m��7��)x��H5ޝ�a{sX��`�� r�aR"�����$�)L\�"Q�O��i� u�M�
����s�I61"���,�O ���ݱ���}�:~K�v!덹��������l���ٮ� ខip�J���pP︯hlm8��MuP<�s#��ݎ}s&��� ��R�/��knY�< ��l) �͹\5�N<�#n����[��R*Cw�z*�(��D��C>�f�k{1s�3w�*��߮��S�-�4n�7�S�
�n{w�Ϟm�6�n����9D"Я���R���ȝ�BK>!ff�ۻ�А u٨W�v������ <����#n��yE���n��`�~dW{���S�k��C��zAt�Pq���"�����>]F�o��;N�+d��nx�-����/�ه��-�<�m��U�@����K�w^cK���,Z2O�ͯ�S��f\WvEE[,I���|�zJy�	�;n�}Df�L�.)(ڈ|�(W��.� �$��mc�M�sኹ�V�GcxvLf0gFX��E��V�0�g�aL}S)�luր�]��1�)�<�Mݹ�����'��pM���X�"^�!G9�t�[���f��u�*M�3A������z���� �3�����߀ЛT��ooK�ٙP�e��yM��_!%#7.��U������I�����nJ��#������B���N��i��o��DI��V(�.��d��D�S(�o�E�W�?v�i�U� ������#�g�f|�����T��y�9Mϝ{��W������GikH�/�$��DCn�S;{�T��N��^9YZ/+�O��N�Z����:�fs�GOmh7��F�D�/�R���b�
�CP������v\F�K6M��	ni�|��2���ʴ�Ԩ���ED�vQ쓋G�y���.�=ҽlLb���g����Ƅ������<�����`�~��ֺDD%QrD�*�����NVw�b,u.P�}�	�~�>�ح�mZ����^Ow=�ѷ7�C�B��<:~�u�ֱ��i���i�&�%<��}�ܔ����m�skW��?KJ20IY+����,9yq3��ZyU1	fXˏ��c`جc�������-l�ϵٖ�>� 8�u���]�� pRղ���Q,^W����ԯZ]��
����Li�|G�_�z_�x%�}����m�|�G���w�_�����l�e�z4)��Ub��Tc�0�or��9-R�{M�|Q~���֣�n� �<E�v�	Wf��U���+��$t��2;→�pm	����Jk�@lYǐ������a�^�JF}�Y������2y��jr"A�Jiܣ�F�Ux,\{ϪO��@�0r������b��{R]_�ڏr_�l]＋=pS�C2�v�������F��`�.:��`�}���(L��U�Y;�m��}8�	����	)�S(�o7�f=��}�l&y8�И�&�JJHX1�2}jJ���+�a۶E�n���� ��?�G1��/y(ֆ���P�R�Ք#Hz����F����&�C�A����F*Lˇ��?f�Rf��6� �oI�_�����i4(�$�e܀"ooC���<��(��P 9j�7�?<��MH�+�~Z��a�d���H�*X�M��g_�I��=(�AR���(X�ۏ{����Uw;��Mn�[�?j/��x��=)�o�/tޜIW 8�-�T��dx�v@�U�P�����@�з�LF�G}{��j�TY��s&�zd��?������qV"�`��Ù}搽��y�Q�ӡ�K�Xd�ƅ�g�(X�MK}_�5n><Eq3��Z�H��y]SE>�Ŵ�wK�ݠn�q�ǀ
�>q-�x���G�M��D�D\���0�πp>�`�k
x��땆U°��7�p�s-�@��_�%/4�WbT�mڂ���#c����>o]�5z���?�T��R7��E�r�W�%��k����M����o�2Q�,M3Ք��i�z:��*4@��y�<�����l����B܍�%,L^�g����O�^^������T��;��U��,i�!+��"�ĸ�rU��x��L�l��s��QOa6-��z��/�� �.�;&�j���U�¬�z!B ��M:�2��3K��@�ܦ?�(.X�����I�����+m8��jM��%c��걣� ��2� (+Q�Y"_!��ݳ�Ӭ�9"�̟�o��1�ͪ�f���*P�!Ml��u�r�q�$��a�`hc3�����-��>h���r%�Q�R�w��d���T��fTŧ��D.WI��|Kx��罛K�$΃���
�w�=f��k���`��	&T���o�齎LB��={����.b�:b�MID�5���/&gh��ZC���OhǵH�:���!rp��GG"��O�x&���e3�p��$d��WaK+ЖL��'���i�`&!��c:?�mF�����i�H0{tyReQ�'��Cu�h������cuf(�ӎ<ʺd,�(ڔ:7J⋚�B+�Z�rB�SƸ?0���M�ϱ2�J�5B�/0�ïi��l(d��xl�������nu�(�o�}Y�X��AW�Ồ��1��)�-ϖ����Lr�Er�ږ��:��{M��aR%�x�w��*q�7�.�C�#��d����!���3e��Se���bj��Á->+��R]9�%OA�B�����tƩ��o� �=�ѱ?���x�/�)u�#ᯛ�w-��l���٠�H;r�ˌ��)�� 
��@��1Gc_C�Ӹo��g��x�f��믲�������W�w�-cv}8��>e��Ŭt@��6ٗLt1�8|ۚ�3?�61�����Bİ~ೝ1�T���Ϋ�u�i������a�vs��^.g8�"F��2�i`"���X�v� ЁsUrI$���#��_��%�0b���lx��=7��1���� �"L1�ֳ@��`E�6� ��`ޔ,�GJ��1�}s"E����F)� �ZaB�S�w�Pӥw��ɷ�r��[H��qS��\ Tr�9t7�;�@�6�R+X�u�����ۆ���/âSlB�[{t��#|��Wۦ��P��'���W�Y�e2f����TKP~G�r��9v��v�Ku����lH���ӈ��C�d^�L	"�p�=I"o�-󓌦G����`%#�Y� 	��W|�"�A���k���?$�U~� 4s��d�|
r._C�2I��'�Ȝ�lV�56��ug����q?)+ze��GO��չ D��0���V�ω$LH��\�ra�;�~	�}�"OOv����g��Ng x��*�\{.0ٟ]7;���@�\)���s|bWfå!"��Zd�w���aE=;�pd���@M�������1�K�z�s6ǯ(����^?�7��RCRz�ܿ�m�k�5�?� E&���(#�L@-��|$�h���S�N��@��78�Ԏz����~7S�������S.L���)P����>�շ��Fh� h7I�O��P3���t��{��&�M����VEMjT�uQ9��.����}	��J���;?y�[(�ޗ�C8�0E$tSr��MSC�x`5��a�9 ^��*��@ ����%堳Ƽh��O%�F̠�J�;e,](hF�^>υ��y3>{�ˆ< ?�/�xuȺ�����1G�[/��ҟ%���$!aFk�v&jX3de��=t�*.ը`��svu���"���_�����Ҡlߕ ��A- y.�z{h�B6Ƭ[��E����ƞ\��Y2��M�5���k  �ǣk�y������HFY.y�`�٠i�LoMto+���H FQ�4sG;wE JxGǻ�j��SlƲ�	�b�$);���q�,ʛL��-���j�t_�t/��(�ҿ`~���\���7&�#P�����%7�@���g�b���� ��I�/'q�	�V&���?�>k��z�� ����Z��R�ޤ��'����[M�t��/�G�h���9n~��]�MW����ՠ��I�\��Æ���@����t����r#��-�l�r���Ǣ����%��=Z�vi~"���*��R�뜪��N>.f֣k���!���gd������~�7�9�P%�1:�3'��7�ħ�����N?u��BL��6h�>�\�,�!����g� �dL�/|�4e.�v�����6~|lcc�ՠ���1���i���'��ײaj�Hh�Gz���:�u���T$5yX�v�7�}���1m�� Zȱ	I��'��6��+W��̜󃽚z���? �~S`M�&J� ��C�q�=�7�.������ŵo��ň���%-���HH'J#ţ����-Rf�G�����(�`>o4a�\9�,t�ϔ�y�
�|�*�,�.x�Ъ�KY�����;��`ZA�2ܐF���UG$?�q��ӏQƌ|���A#���jEǜ(���n��|��?�H�چ:q�+/Aߙ����j7�d�����P��UC?AN�%�{��8d4�x�S'��F{��<�R����w:���6f�� �b��+���&h��5W�ڤm�×�FV@�-avC��|ŷH;�j]K#�9I2�~/���c�s�O8�X6��]�� �oI�u^n4nH�+��٥,�]�X0��'���o�y��Z"�[mV�&�J0����q��TI�;�\_�?ٯ>H������d��al��~p|~�_|9C' �/����&̽^o��;$�
.ƍ}7P�]ېqx36�a|��M�������xq��Zm��#�Y|A����&� ��֟�&�ѬA4�e`ye���ߔ��g^�{�f�$��-�7������^'���Ӧ�5'�Q@#2��_S(M�`tg��ԈTX%�����4$i xI�㑷��^R^���J	��X}����IR`1����-Cje�Byu�Q�=��$d'�ۺ�9�Sɑ�h!��0�}ߟZI�'�ΧwbfW*�È�0�m�n�u��y�Do����]h�+�ڋ�s_�ǳ�{P�ċA���ߙ���-17학[�)_^��<�#U��cG���5��6&M�e��Ic�0�q�	��&��l*^��A�{�~'�qy����!�8)h�vW��Qw�:�����={�>Ժ�4���W��8�+mV �#L�i�I � ;x����F�iζ4�ՅE%���|�s��(̝��7�,��`�T�.��8��B��ĩ�����9�;�0�-�ML6z��u����[��|'*g����1����`Y��I>�X�g�Wm�܈\��VT"P�!Q6����Հ�&vP;?�*�&�#U�k3���@�Uq������&"�^l��o��k��>d�Cn��"�]���_�C�������I�0� ��=qC�H:Rl�J�fO�������$������')�m�m��F�9j\^�*��SR:0|o��9�3�%f���Q
H��J��S:B�����9�-b��wH��gt�A�$��6��x��7���_�է��m
�5�e(d^�um3�߭� �O��\̚�i'=�(�q� .��ϧX&�@���V�u�{��Pw�;5u�Cg�m�	c�f�_���3�  f|��8�M�t�G�����U��ђ��&R�$�����YK�~8�T8�����%�����2�V��l뗾z���ZH�&(�	�8���Q�z��Pr͕l_ڄk�3m�����ñ���~(��c7<��'d��r;����	����Wa�F�r��;��h�ds���&�<�)�w���PL���S�p��Q��+���&Ң�d��ֳ�p!KHa��:���I��/��7%IC> G������P���e�e�v���
}���5�+� l�mgÆ
G2��N`���ٱL֗����iւP܆�C�ZN�]y��)����	�Ӷg�bs�%oqն�Xd籚+>����s����w�ڻ.D>R��f�N��"��'+AR9!���rb�o�5�Z�� ����~'�����L��8��!L��h�j�5�5F����8��Y�4VLk�����cI�fd�t�L��^�T�X�#���a. �0�BJ+��������u�&�Z����]��-9���=��9ĄH)��а���	d��m,�̆F�:�w+T9w�L9�p$m�3��v��5�78ٙ����fE7%�sop������	X���}��3�=���E������j@����n�PZ}�w
����OU.���"�L|��D�UB~��Q����ܽ擹L&(&� Vї����{,yy�:����#)o3��2[�$\ag���N��H�XU�i�=h��c�^Wp��a��ġ��/�7���1�fзK�O��E!��G��ן��z�)e�<��!�{́�{`�f���E�p;��^*�p�7�W��o�Tq��-	U���NP�B�͑[��.mg �Bak�u#Lq��-]8S�S^���X�3��a����PkPx%,o^֯��ߥ�v�}�{�Q$:a�\7���H�'�F�oN�ά��)<5�����/�0K�=�޻�94�C�ԺF������/�����z���hQW|[}w2j�JWj�;x�d���&H$$�6,�%Yp���q����S��%o<�.���&���;�R������hl�iz;����0o���Sw
���l����"�!����`��~Z̻��\�,� ��y�����ӗ$��������'�ȣB��fAg!o?��|�H�B/c鸹�6}%!�c�u�j�2l\���)'��c�V�	U�������|:JN)/.;_�f���:��^ٹ�B��_��rm��"~
��$ �dl3�1 �gE� 8�D��`��z�E1�#�2IHqX�=8��o�
>����ς�4�¡nۙW�<�R9���i��Nr�Eݴ���s���	ki�ͮ1�0������BZX�e�T����L��kA���5��|N���z�>�P,�O�l�/[,���RSm��LD�Z��Q��ר�"�RTqE��X�Ik��:ז���P�W�ݒ�(U��3e��t�1W�T�T͈;�cAu�I�~�|��o/�+h��
�N�J�J���zn���k2�}p!�}��7`�f��dd�'q�Ä`ݜ���SQ9�C�ģ�@�j�rL�É"+^�Q��#@Z��E����j��"��I��u�⺕�X|���񏔭-O<Z��[��V�6�1_�$o�O�9��<�'�T.�ˎ�/A���{AW?K<1~��*"�u�>��w��}z\'��d��Ĉ��}5Z����L۬�	9'�k~�~Hu��K7/���E�?��yMȚQI�>�c�5у�q��vv��)��;��#����3r���*JdP�q$R��K�a�V��}�@��6��4���1��s�W#XZU��{I���m�Wg`$�qH'�u���$�~`��} ��^���Q��b�'o��N�([�ĝs�#��^	KU
��tv	����xT��u��/5��N3(#Њ�0���x��^N�@�N1�Ǳ�x�\ķ�i=a�$�s
�ת\�atS4	u��ed)Hv�y�z�s�G���|%~(�*�T-��<�Ӯ�������d�9��7������mN��ڲxhq�r�G�����OSGL}6n��>N����+���Gϧ�.�����������'�����]0�˳W�!F�5A��&{���U7)�ˊb�FλO�4*]I��Y�I�Y��U�8�f.�b�Wg
��q̰"�SV]'	���]_��猽+~��*�I�%���s7JV;c}���zd�X�?�h��-�1oKd4�^UIXŞ��e�q��,/�29�] ��]�Y۠�`���� i�!Ir,�y6�d4?Nz�\o6 M"�[Sj�p3���rR?,�E�������_�^���<�B-O$g�p9��H��&A�ma���27���y�1�������<�99-$ �u�଄ۈ�נEc1҉�SB0�R0� ��"�C[�pxb�lX-��۷U��<4-��D,)	���{ m�@:Xr�|`�{Y��Q�$��$r�$P�H������k^�2�<�R����,�9��GDw�F����A�۶�d	����ȽZ��?��z�OvC�7���wV�s���� m����a����ėn�����J$,A�����Kƽ/%E�U��d�d�	z�h)qJ��̮�t�cU��x� ֣�7�,D�w�T�ox�/�;>b�^7��v�5�A	�(��{1"UM�Ҳ0h���T���`U'�F���^n+*n�,�2)`�}\PkЭ,��h�g�� *�j5��ZMe�k`lg�q�:��R����b�Z���G����S�C�z~;;�rJu[�^���Ѹ�2,R&E@l�В珰�M���*��M̍3��A�\�x��v�_
�.ȱ�sK���w�7�yE�D��WY�������_$,�1[	��}�å�%��F�	�?�u��=Jh�	W���#7Ԉ4�W��mQ�(�A��sc@�������8V���I߮�������3C�ݑFz�}�$��Ke�@���A���o��2����Mz\��EѮ���������A��(m^@IP&��x�ϴ1�W*\$���R}�?!���i�	h[�^��V�~��U�y�~�X��8h�H'+)�����Z�A
m+�irX�s7;V#hu�0mY��*f(�����.���"����M���X9��Wnu~�R3JV4��i�:~IId���t�e��שQ��Of'��.�&+W�jO�w]��� ��r����r�M2��kv�t���V�٨� �(�dy���k��}K�(��Q��eW#j`�F���;����+�����ʺ�K�PHw6u�8�n2Cᵕწ}g�_*H,b�[���Xh p�c$C���{>��;��m��y�Т@�-��!_ʭ��2�ɷ����cg;��\���)Lm:��do���rl߈�:NCV��Q,��ckCE	��D��&�5G��
�"8_��)�1�CJ�yOYe�Nh�Z�6m�7���O_A~��_��:���u}lX�����h��=���S+o!WV ��#��g��O+����3`�7�Z���G��P,X:���U��:xu�B�G�ڢ��'�-�����a�6Cv'k�A��ٶ�s����i	A�Z��y���(����͏-�$E�.$%�;�Sa�o��� �4 �IF�^�_������Y*�I�:s>62�s��,�~5N5����؟��B�?�����U������~'��fA(0u��)b�����Њ�6�`"��qV
$��9���u"%��Ш?�����D4���{u5�K7�#���)�t�[�z4@܂����7��,	�A�:�q�!WOn������Q�\�t��/]G�*Q[l�7E��5�1�Diȣ�V�l��\dgN�~��5� �92�x;�cD�Ҷ֊�$����:�c��3,~�o�qτ\
���iZ�lU����oe�Lͽѵ"�f�X{'\R��C���Ե�$���fGh��1~`�t�{����/�)�Eo�q�]>o�4�� (���1b
����Kp.kVA�]�H��p�� ��9�j���uն��F�wg���)�v�����R�h�\)���L2t{�S=Y�`���5��1�)δ͓�KƠ���O*���r/����}{��jY?.����_����r��h���O�e�=�����8�9�b�o��䔱�4��ob�5H���e��R��"Q�ղC"V��b,�����}0X@�c&��r�����ҷ�;pC���!�co�ww���Sx���)5��n�c	Ru����r\h/N_50��+,��6�����]r���Ȉ�8�_�j�w�D�R�ۺ ZRIB�v����@���.y�c=�t$�+��4�q�nbR�,��-J@˘;�yT,���ɲ�Щ+�Q�YDp��^�
��_1�o�����&@�����~B��; �o�%�HO�f�7H�z=������g���;X�y�/,猛�,$�����q�#�)���v	�	jSe�^E��� ����m7�<�6�~ޚY��g�4���5F��[�|Ok��W�ȪgO�e� ��vNp����$�\�6�C�с���9難b�����e� �0��uc<{��a��e��[�W<<��tNg@�n���`�ƟA"��Q1����B�~��;�΀
�?�%�,��J;`�F3a��""( �2>����4g
����T1�x}�ܐ<���ޡ�R� �NI$�1/��� 	5��L�g�����)ԩ��J�P��R�G�)��t��*K�hYv�0>��M���E~�1�D��������Y��"�F)�M���D��t��`�E�	^;l�V�(������2f�Q��q��(^������')������g�����!*>i$�l�$�~ ���r+��yM:��Mu�
��@~��2��0�fXD�AC1*Y��@��T�C�
�"���F��F��!�{��S� Y�N	b��9HM�s1�2�ݨ"�9���ޮN�'���j�����"]�29JM���s�L`wT��VT7�����h�7{���g�� ���]�Jʏ���%y���0*�[��/�?���3c �@]�F��4�&	ٱ��G���k)ers�T��5y��/��f�=$�K�T9^n�>��н��M��~<U�G��:��v��ѧ.׵�����}����|g�K|*��NTǧ`�i��I�� �r�p�_��a���7D��y6�׿^��%4�����Y����K���_|T��7�t>m\���.P�jJd
�|xH�g�ޱ�Wv2Lz��x����q��8�&M�\5>������3�.��$�ɷ�^c��%��;���H;.���MguB*l+��vPq�'��=�����!��^@ څ.���UOm��ܚ��[Z�h5#�a�Q'x��#D� ���l3^U�����u�G]��SHݩ��+ �):�zd�J��m#��(2�A��B��_�m⥘��ym�{�q�i�����v�$��#Y�0��a7��K�ㆪF2>p~rV��;z�B4l��Q���G�$�]FA'%���3����W'�0b�	�d��F������@c���]0,e����XҖR Bi۸`J�]]p׫��1�~��y2�*E#�-�%>�����4�-]=�E[*d��~�1(�SK���ya�͂�C`T7_L�[=���g�'���(S0P��Ο ��l�V΃~��Z^�*g�3Xʬ|Y�k��G�2Ұ��0Eyg�U��z��L��|I�����i^9d.���ǽ��3��_�W-��֙�ul�q���O�+<�-? ���̕�_���Z�8� 4/xB|����O�v��#�#��w�� �j�t=�	���4�f|�?X.ȇ�:^�6ė���2z7�j�ʀ��.�-��SC�\9p�aQ R~�sU�7��p�?��7g���Ms�8	c�����k=�[�*�4�)�_��0,9݇�����6����c����Sl�0R�L�e�K��ߦ��ǥ�<��4��=���vu���o�1����q�s�|��t�!0�"��X_U��*��v��V�^���x�O�(~�j�[��u��o�J����.#m!��`��v$�I�ή��9���v?~�;��tP���F�g9� �d)�\��h�J�{L 7�k_��\��Ȭ�y�f�\5�魯)sf}8|J���Φ1VS����;d��(���㹯�6��;�`(��ư���{�P�����c���l[&@e�G�$u�,O���U�O���Nz(L-g�M�a�V�hH�4&�徚$eYா�?s��0�(m���� n��뫧,\{R���e�`D���Ϝ?����#յE��9QD`�|_j����k]!�\����6�
��@=Ã�s2�riGʲXVl�c�Lǿ�l�N��*�M'VJ����:��-vΰ�D�v�T���!���Ho��x�� �;1_�4�t!{~'���y)QF�[��TY�B%�y����N���!�rx-��������M����Atۇ����l����V�^BL��Rn2���v#Ұ�*������#O�Rsuu#D'ʌ��u3H���;��W=H��isGԫm򲥅RO�:t逷��'+�}A���Q��0��7�
\07g�n�0�A,V����ݖ�WX�r�u�و(�-@(�ˎ;R�����X���ʻ�E._���%2�X|�������p�hZ�n|�5������Y�5�%F�/W:�i���Z�&���e��:c���!%�8���\ab��j%���z"��o:u�㤓����N'w���_[(�����X�k�\���P�o~��i�������jm���0�ea(M+��*�[*�Th>�{��h5G��u�U4% k7��;k���k���q�$�`K̟��ݪJS��*�g�	$��.�!9���=G��Y�ZtI�{+�ٹ��O�������ViH5�0n�t'��C�]ޓ��̥��
P�� �z�s��e��0�AiO��_�3��cUgJ=uD�k-a!���w�S�����>ٲ?*���V�Vڡ'��WQ���-ܩ� �x�����#>�67~�!�HS_~}�@�al��М��{-�j	�������z�G�Y�H�n9��K����7���o�͓}ȡ�\����)�Nw���GO�T��\x�3��[	?�b
&z�Z�a�_�1f�Q�]���/�� �L*���דu�l�4�l���{�%��˭X�pԢ�a�ZR�;j;�hQ�"bl������u7�p�� <jω��5�Y31C0���U��HjC��^�.���ݩ	oƀW*���� �C�ۤ���ㆂF}~J7W:�F�^ޟ�t=*����Kb��|���Wl;�Chh�9=,ͭ�5~A����{Ȗt�� NTWȻtᓟ�d��q�$��M��6�A��
�k&�����W�%Hwz a���p���:(�@=�gi�
r�$]1���F�Þ*obd�͇��9M�����-����'��������+鮃R6J��慥)3�LC����q���#�
 ���X�5�WH[�w^�̂�+�I&ږ��\�o�>>X�ψJV��(�l}i @�n���b�K���뮔iXKyްΞ��p���A��~8���x$ܡoa�z��K">c\����ưΨ�A���x���1K�!��%2&� �4'q�$���\+�Xڐ�MX.^�QMj$@!Jn�SQ��Ճ�<m���:�#�u��OK`f_�;`<�[D�p��sե�M��&�!�N�ڃ����\]ErM�N�#��~B�T;��M�;>�j�;Y��T9ϹF���e#d��Q�0F,s{�;�V}1�1�$�=}pu�ö��; i+��I��n�J����g�[��T�|þH><lW;ws��)��<&'���H���K{�O�����Ҭ�4�@:s9i�z�'�Z{>��O� �?".��Z�KfC��?�=���̹�����LP]���hū$Cͥ<o��j0��ޱ��kb�ys\���s�g�2a������-j���x��WM�������|*�%���E��+kD(��>y��g��	U��X�EM\�"��ś��LZ�sb�W�ޝ
����u��Pk>0L��qæSr�H=����<k�e�S1v�Z�"CnO2ބE�pӯh�����<1[��&�Q5c�左\>rħ�J|�l<:�汯yy�R4kQK��;ߋ��m%nEI؆��Aև�|5�خx&Q����J�d�2��".]�-ɾ	w���,����+ݤˊ�|��cf�rv���t�
��W�.kh04�*oX�i��?)����b\��N�))K<��t�����DG	xm�9y�[��{�6~�qJ���
�EL
��g� �̂�����%�VR����/�\����rV�~�O�ϻ+xe�
���]sJ"`��R�������	���H�ԋ�
d�K`J�x�LB{w撆g�j�r�m�>!��CN��-��_�t���k��+崕��ȥR�8�T��ch�'�L=�Q�U�A?��;�������B����D���@�x��ډ����o���}uFRvci��0#EA��2�Z�_Ex`���E�g��H�7%T��yL:���л�jǯ%��Ġ9V��7ZP^h��3�a6�Mg��jXA[w��e1��ՆC�KJ^N.���B���S�!�%�4V��A&"η?)�Yq�G�+t�:���la�X�5�b+5�C���pb����	O�"��-H�9�䑩,1�3dJ#��E$���~�xt���J��!Q��Ճ�3
�!�(-@ik������y+���w�|�$��pU"�d�<�]�t$NFdx���aJ�p�t�'>�g��l���Vl׬`RE���ƀ/�M�D���)pJ��	j�r�T���o�t��yh���E��*k�P=CZ�>�4T){64���0 B�6#�-~�E�DKaɃw��s۷�� H]�|z���o�婸D�g(�ÁaL_�`=Ƣebg��P?r�I^9��hh\"�A:@��gѮ��!���"�](DM��H.���>��d��J��h�0��8���g��Xi-4i���X�o�9G��֮�p�o#�h.f2.�A��)�{��i.�PBz���7��?���$��H
0�MOP�0�U�|0\���%d�].�~IaU^+;��t�!"�0w;�+�j40��Q0|Ofb�S
;i�C�E^�hӽN��A���QZf��\9<ƙ&"�¦Q���z%?��u$�F2W�_\t�LYy[�rMa��h�R����Q��m��)1j63��FɄ����0����3ZÈ��A�>��Q�Z~������k5*��������')1��e'nQ�Q������q�-��X5IQb�7w�QA�D
�m�ތt�*<�xB=X,�*�3�U 49�׻�E�V�B�+ƉhV���wqp�f6�y��$�ǗL��L���,j�i��J���,�	�V�*�JnQ�	�>_cJS�BIo����ۺmn�z�Dp�����hm	��,#W�����/��5�j��O�B-<zu1�i�B�{-'2X&����<��i#�|@T�'�F'�`���r�%ډW����੺i鳷��=����2��x���Hht��'��w�8�E��8e�BzQ晇����V|��(מ@s���Ӽ���{���1oy���sA�p-j�#�I�]Y�����_4�����OY�X�4ߒ��sa�_lAU�tqr�r{�Q%���!���6 B�����ڻ~���J[-��?�B��\O��W�%(��RiJ^�`�1�`<� ���d#?B�90}s�<��Қ��g�����w�om��c��`�#՗?
�1�,�2�H2���WN��)�,ic*��坷�#A�s�B*�je
�<��g�)Ǡ��:�r����%�0����X�ۓf)NY��+i��EL�cy)����mˎ�Y����U�AiS4ìIk�O�$�ͷ/	� .O�v ��e8$�\����#��R���	Â�W��!�x���:���1
�1�mO&�B0� <*���W����Z�9LC�͓��6G��o��	��3
�ēq��v�a����n�y�����B.
�(���7�b��T��.�n�Ġ�#�O�cJ��/<w���m��i�ȏ�����˿��k aNs��F�o��͏�Ɋ
 ;�8��$ckղ��#�c��i��t�i�"�]��$��Zpɯ{�|���aa���.?D0"�z̓�@U?6��Wؼ�j�u)_܍���+�5�}��q�1)4�}�ڧ�nq� Y�k��FP�hV��ǘ���!��UU��ҋ�z?H��j7�i��}����%WYzZ�߇*�m�YnFH�&�Ewz��@��}��rf�5�2>Ƥ��=y�=&4�`�;�2�i�Lh���Tz��TnU9�1/����E�MK��k���)N�p��K����PB��CzXI!=��!#�4��&jf�ei��-��9����I��X�K	L����R�M������2�*���;f�~�,$�vl������o�Ӗ�I%t3����_&C���T�p2�mѪ�ʟ̗�ϱ>�SV�6i�B'/��D�Z��cf/L��o���ִU<])��D���[S%�	�������#�����x@T!��<e*m]LϺ�TN��L���=���8���Y�m�K�1�Xѓg!Oyϓ�!����aU��ٜ��YN`.o4`&�Q`�1��c��y�睍�	�_<V�n��^*l�R�v�k��!��[�3=Q�y�fLa�Us��ǈ-�.��mr�x�K����/]��,0Î�U28%�ʹ��=�M��
9��.lU��>(�.W˓3����v�{]�;����c��e/i�^��2�a�oC��)/n����bc�s����5Rn����U��rAy�(�bk� :�O1��w�4�B<����^�<����ے����p�/g*�[7��')/Yp��r���M�f�&��4�|�A�hGy�����&�#W�� ��P�)^ ��5U�
��p&�&N �8�0�>eeG�4	� 7���Q���:��&9Vq��U8���
��nʡ�l�b�AR�Ј��GJ4�@�4�WT�&�t*K�n��qU`c�1z��7���7J�xC��R��)%�s�=kF�f: Q�C�����>�E�O����6`��v-��������ԩ	�a��À����S��cg(� S�Urw25�~�Y�r2�'*�(�"�\�A��n,��*_<�j@���i��
��d�������$t�������ʈ��(�;ןtN_�	>�0.��	��;:�e���!��s
Ex�R�g!��R��o����QB]Zb�ن��x�L��BTy�/.Ő��[�E�A�[.S�i��'�}6���`)�;���"�=.�~ۈn��ob���SƯ��N�� 1e�a�q���ܺ��� �:ԭt��v�;	�dSvP�wk����E~�z�GJF%6Lt2DT[lSe%�������yͮ ��"n�^[�5)0��^i�	{��f�S�98�F?�i��N%�Y ^,\��J�Ȱ:�s�`�a-6%�IA��iIɫ�� iY۶F���EZ�v/ ���ԥ�ďR9��>��v��활�'t"�(����&���F�Ң�*�ث+����&�K��z�AVAL�=����W�0A;i�0o�JG����F(Jj7�鑮�!Ț�xt/hn�B�P��nT�l��z];��}��Z��&����\�9��T��b�`K���Iu�h��Xl�o?:��\��/}�Z)����"��M2��"�����x���,�#�2ˡE�_�ژ�XL��&*e
��bR�0M����Z�Lm{+n�C#��<v�
rn3�-b@}�!h�~�u��r(&C�+q����I댯�)�T���ٮ��}~���ഇ���FYrL�� [��7�L��9��'��R���*.t�푥ż��P#�i�X���s���n��|����,��<�,ʾ�c��Dn�`�Tb�����.��W���5�@�2� ��;����Jl�F՜����}��f^(��.����t틫��:v�t��U1��.�S� ���L��r2��2i_�PH���?1x`F�����E�{"3��11�tʳ�'�5׎d3��a.�9X�l�gn�)y[Jr�����C�}��K��L~�	�ҿD�nK� \�nW�HO;n�� ����
?՛ڬSń�3���T�#�h~�����L�=1��N> pw�˹%�S��by�2��1��9y��V�V�>��M��K���X�MI�oc�2��RqJK�u����_ݸ�'��4��N��h	��N���z#_ž@Wl�^h��������>�u��P����Z��Χ՝���<��B�SP�7��:�7"f��#e��]Ms���;�L��ab�0�cѠ��ǅ�P�0���9l{����#@祜���~��އ���&|��_����if-�����߮r��y.��+�X4
���8��H�LXu�롕�w�+�:�����n�ԅ
P����,��+��*���A���>�ÿZ��A=xI�H�m�w;^(��H�I��/Vh&Sb쐆/~RH�O:��:�u��h��~S%���Y�q��s}�rp�|����q%Kl����䂹	�ޕ-�Xўn}_۲;^
7�}��ʚ��n��'����gnjet�"��؝Fwy��� z����?�3]4�K&Tm�I��/3�#8 �R�����P�*���dc�V�?D �pȩ�^��:,Z^}�o_	�b{� p����û<��TQ'�$Ӕ�儀��O�bp~�B��s�w�s�kA��E{�-�wqd���K��.+{Y�Z���q��bbo7�u�ͣ��蚻�	��2JE�c���"��ё��C�N ����zKPd����e��,?^ˢ��1����R<j�3�6�1��i���"���8��z+o���F����U��9�@̸x�N�qr�l�`�!/_�L���:]��K�Mid6c�2J}���#��e�NPa��c`dv<o�i(hX_���(���3����ӏGF�@�X=�\~��͈ai6�+$�Є�����H�)В�]�[�'��W� �����+�A�E&�7G�T�۫�j���p�v�R��j�Ʊ��:gc+��_���Z�̐���O�2wǁ���Ƀt)�GG�j�.1C-�3��3��R��Z��'�a{�w��u���/���K�W�v�ց	_����� @X�wd*���߹��I���M8�шsI�y�����nƱ;���zq~��d%�]�����B�Ćl�]�u��ꪞZ!a1�z�烫�����ZX��Wҁ���r�n�� a�h�I��}���r�I�\4Ł��a,�~����Ӽ���a��B�
	6X@�.���$��Q#$ɵq�!BL	�g��M�b��W�ER#�y ���	 9���p�0(����e�&^��a.�Y_>#|�a��D�g�?}"���y{%}��<G���u�wo?��%V>'i�杖+�J�B��<; �p�5Ԉc�����9�Df�!%Z���=~�y6�
:7�IZ�}l�Moia��2�(4�b�G9X,ex6Ӵlg-sݔ�d�~J��o"�z{�b����KB�h������hm+R0!���0�E=/s�!�?�prK䀲���ad�Fh�g~�pw��4�X�I^�E�@�ڻ�5�Aj�!��E�wd�q/�F{��m��b:�����"�2ʖ젧t�ʁp�������HN�<Gk����3��[��_�3q��C�
�A�"������Q�Bd�&�����=i��0���;��!�˓�u`&Ӂ.��|����c�U;lY��{R�Swt6@�WsU 77���]ս�Q����fڕ�/�;��ӄ �>Tsy�@?L?��Wv�Ki{����ᗍS����w�ې���A�-�-�����B�r��#���p�'���iu�΁��Ö�GJ=�B�Wo�/qV?�P��:$�������X4*�Rt}t�)n�X���^5��bÐL����<�kK׃?��
��7$G��$~��z�م�_)�?�1u³3���GR:I󋦪嚿:~8s��\f��ֿhd�ƣ��+q�xKm�+8��˴������6��	ME�i9��#�V���I�������@�K?_��E�� !+����c�Fz�v�^3�t�X��>��4�����aV%��[�Ⳉs>2C�l 18 ��j���x_���+P�����Ur����}��	ѡ���
��ѫ2�G�y�D������W��h�xWIJuC
7�׾�I������?aHRU�^6q^<�~�,WKR�+�#��`��0��k(Z�&���Gf�'� Cz۝��|�&�^a�l�Y��<fFq���*�Hi
���Bt.4|Ik������+����^򋍰C�_[T��I���V��b!՗�]M�q��gF�4�4�Ov8d���О��G�VŚ+��f�BO��
H�l�!�W��9��Wvp� 1�����)��ז�y�-�Z���A��r^*��䳐��F(�!}П�Dg�G&U�iZ_Fj|r����I?\˸m��g#S:�c-�U��8�_
��A{`������O��"��ޡ��{�h#,e�F�Ӽ���J.f-���VҶ�W��K괿�E
!�NE�IT� NQSa���FH�up���� ,�+���\7��5��f�*���s�ku���>� $pDoS��_��Q�*q ���HI/��*8�*��պ�]�Nn���}���A��̟`-���C�TK^� ݡ@��*����Y�r�/oR�K\�|�0R���q��9n����y#��	����9�T25�d��QL�m߅�i��]��m]��,���obɒ�JHQc�P�*t�[��
8���d�N�頡3ޯC&� ���PhX})zi_��.Hv��x�%�&�b�׶�i��] G�A�g:)���+�Y�K�.~@�}S�4*J	�h��}�B3��s��(Nk�^��.tTl@�U����g���txKB�˕$��t��>6��Xp�XJѯ#)�� �<Q��C�- *rQM|=����Q�5�PC׹֏~�_�bמ�G#��tVb>�9���1�^�������p����_v�(2��~�TS����˓�
募qz&�6��ei�o	ƶ�o�h��u`��v�zK,*7d=+����H>��[l��OZ��v��=���%ѻ$�7���x� ��VY�����(�/f�j���;7��Gh�P�O�7_��-�H��
��fld�\3�F��������M(זoP=�5yiA�:l- �(�)µ�Ζm�l�1���,�X㩹b���*�x�����Dw9�fc�~_;��;1q ���7Z
��g_��k)؎��^�:�1h��5,9�pC�'��lr�@�T��-o���"��zY��p[ɈjKܶ#B0�l;�D��\�O�G����պ��vmD�e�'cU��T�Q5����(��5��O	��Dy]�F�` 렒Bb��^���8�V�������`�~�� �lw���B��;��&��6���B����W�vo��ȅXO���9A�aX!4T蘕/]�0~�.t;it*.��򇨔[��0�n!��B^(���쥨�G+��G��_T����m��c�&UB��Fc��/�x��N˞��/O�HL����ը����1���j4�d���,���w+ ������<���f�d�;OD�A�)3p�^&�X��2���یf
����{�<�;p�ԲE-�{QJ)�D�<�Q5�>��:���o~��K4G
���┓�=�5��C�f81z�(�*:5SZb0�	'����G�]
��/���UT?�Q�����92��^�MJ%_� ��l�5��*-|@�����k�'�)�ݸ�[S<mG����X�7>(貛%ݎ�k'<�m�:��r�g8�hA���@�Be�U��GL�Y դaR�Б�*|j�T���H�Z�SfNd���1�;�$�LM���o3aվ�V��
��(��R/����9��q��d�ٛL��������[�B����_Hiq���2+�"e&�*���m"_�$3DL:������;�1}��|��js�ѝ=Hǲ��?A� 
��$Y��������kʹ�45((�֟o-�c}�܁ʢB�bls"��gv�>o�W$\b��3��0Vt�bp�Ľ�|��|��<�,>( *P��`�k
Í�^=��.��e�`ye�I-i �d+&B��
�	d,�_|:�$��S��MS5��O�r������N�(�qtK�oo9���b�; e^w�%��-Y�E����((�~��8~�k�X+Ê��L�����Ԇf*[i4�W��Y�-wv0�~P}�j�x�.U?�j;��R>KI��Y������69�ϴaB���L�]T�4Q3U_5�����+]����{�^ʗxPql�hK�ލF�\��R<���2J�-P�̒�#�.Ev�.��)�}\u8>�����b�� Z�YLy��ѫ�!�f�m2�������wGc?�QV[i�	N6�ٗ�������絔O�ޓ4��Z���X��Ac[�l�XZ���)Wng�l��
��am�m�_�rQ���y�[�pI;0t��R?a��//�j@�B��i�W�GN8H�����1�m/_��u���>@4YF����4�ć�\��A`��A[�� E�˻��b�<���JB.�k�<.D�N���˹�|�6�;�9������?�ІZ�sb��v���kq#�bܪ�e��@,��n�J�(Y��v�������,����(Ș�^��0`$i�5���"�	W>�̺��}�9����QO�߂-�^����9F�7n{@7ng*a��(�r9]"a�v���m�8�9ڰ�^!Z\FU=S|'���8T�E^5�Rm�-;ls�ѫ5ǋ0}�-��$�nF�g�Ϋ)9�p��H��AXg���8V�`�H�)yN3��IՆ@d⯪�_:�N��J�Z�c�E��t�ʚA���`�kx�	�}dA$�;H$�l�FRGb,H�E�h0�E,��^�� I��v8����~���+�	iD��ѣ��	��:��`7��w����/f2�i;��[X�Yv�xf#b�'�E;�>�`r�\����ՈÖ���Ƃ�M�,^�#�$������Р�N[���;\5�"�wF#�/p���#��Vh�#�&%j��MG!��s̥c[?l���?I�%G�a�X�.Ů�(��Qlc%ٜ(yFB��]S�4��#��ˑ�l/��������+��hqu�u�\g'}yk�Ǒ��R�p�T`��� 6�8��I�e��.�M��m5+�#�,t����/?���0�3��v���1�B5� sl���z����F��(��@C�ed�]Ւ�$E`P�C����v�V�~Ŋ:;��E9Ե�v��	s�]�J}2�M��R�Gaݿ$}�Oxm����<4ݠ�0�2K¸S�t�ڊ>?:�m�븇�)� d��2vp�ԏp�Ij���ල`Q&�k�~�0nǅ�ie�9�u�'�t��e��n:��D�$��b�(��wn���K��<W*�+���z�R��̎<�
�jj˽ZRE3�6�p�0��K��Wؙ�	�?��a$��x�
[�e$�8���L�c��F���r)Y�)'2g6���M������D��~񌎶�.A�Xh����lCXۏ
.|¨Mkj��s\TIS����~9=[�L�x�W�T93���n��{��%T�WNx��ikA�5;���i/<��1�/=������
��=��'��������p�C�.��l�i��|��2����gm ����UE��Dj�w�#=$l���� R��x�范�-Y��Ĉ����P�B
�O�,�r��,��o���o���v1�䗠�K���8.�9��zuh:衪T�����Os�J}])M0^�H�R$o�-[?ji$�:0�=[��&6]#���"ZF�U���L���(�$���1�q�sG::<�THl����=}LeF�s\��q)��[F��&�L�\�b�6�����6-br�R�/��b���9�(m�U�"���B�8��@GG�5���E����g�i5��N��r6����+ڼ��НHK+`2��9�Tf���Vc��2�l�]���A�ѱ�e���˞ ���ȱ���@Ѯ,�Q�1���M=��`3b/���<����L��@�y�n������hk�s�b*�����f�\�5��c-�U��z�g-O�(��A\�^2�֯�I"�PT�s��28��ѝFU��|��v��������5k[ a�/Ⱥ���(���v�\pM
�}SՐ����fm�skJ�g�Mi�&t{�F�D��_4�xr��-2vOᏠz3�)��K(>��3N�^��ڦ�j]4��B��"k��;��[�Ǧ��!�:u����A铕.�;�U��]Lu_�v�mMH̹"Z���]�FX��!����WA�<�#*%%(&�>�٥?c�(��9�Z��N��\w�7��C�aA��0e���"�j��nU2d�̀�:EJ ϋ$�%��fNADm I��	����X��?q;7�kzs��������x��xZ�Ռ�a8lq����U��ŬN�7 s�@C��k�ӡ5qD�A� -lN��'<n��0[͸�%(����Wd��X��2�����;�_4%�9�8=_�^�Ibv���+���|0�3D�����|4!K�7�V��:vb��7x�'˾����8��^��`	�z��,�n���
*-�ϴBi[X�y��Cc�H�'�_U�x=�z��Y�".a��<����6A����@��	��"��_���c�y�m���X�9̑��;�wA6c7�I����i~�A�����=��v����m�re�y�*���pa����T�y�������P��%\!ft�q2<L]������L!�������F�
϶��	U��q�����_�{B0h�K@��r	c�h4�-T�|iw�8g_��2����=z���J�'�n)�T(�t�dj�O��Ta�~_�}+z�)"��O�B��������1-�H�H�M�o=	����t-܌d��V��h�n�"
�&�����F�ui�,&l�7��8�@���K��O�4M6�P#�������h״��ʰ11 ���/��f�jK��I����{T�kC�g;��&woSР�y����m2��\fj�F-���*��ǹ*U�nh@}�$d����?��
+4I�� {���N`��d���s�t��S>��(�?q˄�n�Iʘۨа�^�4���Њ֨���Z`M��*M^y��~b`���̎e���}���B�m~$�����"�j�r���?��;.Y�H1����VW����1�Y	�	�h���K� ��R�O��1�K�c����g$V��	����e�m�V��BJf�J���.�ֹ�87�}� �5���il;V���W�]����7���-0q) ��+m��zpVz
�!e�7��{J��=�[(�~��ʘ�}�\�W[�A�f�G|��A�8��bȰ���� �X@�����J��5#GH�x���	�h��0�=��؊�l��s�H)�u���5��x������,�S�� ��� ��R}�_�C��n�{cP)�����@�����R���!Sa*6�����Ԛ�_b��k�B�'����Z�b���G�G�'U��D��d�	CWo��)qv�\��1�X���}/y��-�,��~��!���Ҩ�"�G�dm��v{�O*�F�9H�#D�	=M��Mr�܃����U��rd
����|&=�|�5�P��VRְ_�	��6�6��k���2���y@���A�1rq>��}��l����u�B.�m�!�2���X���S����_�V�u���AW\�R/��5H�����| T|p���C�zQ5+ ��ў�I��L�T�z�;ovդ���#.N�EW^�צ���8_$�]}w];��K���^>~�]��Z��,�W��砝a��(ŘvJ%�Q��|n��"2�x�Un��Sͳ�iK�H�P�����(�lӚ���Q�V��MK,t6��7�<Y`�}g��R
 �ڠ�>�%������.��\�د��F����P!)v�AҼ'�ӐM��.�/x����h6�"��
��Q�DD��$���1�?H�)@��R�jq�3V2����(8�Hp��/�J�EN�2�`rvz�5��W-ӴR���)-�����]��}�s�б ���+�'���	��o�X��?F�w[��qB�#��]i���[��Ò<fkD��e.G_����Z�!t�L�����c�S�ol��N���p�(���=�]�<�w���j�����n���M(ʒqMg�w�]Ȏ�D��t�14.�6|S��R������yª�I�X��`���"���_�Xd�M,�r�{�E:?���
ר�n�/Ο���p��@�����E���6'L��T��M�Ki���Azu��&88#s����6r3Ԩ"�e�5��904�tN3H�\��0u܎ T��
�`���H����S�r�8_)z�WP�.Qb-M�P�%�:�Y[O/Z�Yb1������`L��<��XP�,�e~(��~$E��NB�(H�`^{*����Ek�T�Qk�6��e�C���6	 ����-�"x���0h�� �V��T��L/�᳈�A	b-yYR�U���}�ô����/d�ƃ��5����B��Qv��}	� N�jÐ�S��]RQ��b(��إ�.�<T�~�p�,������	�٤ۿ�NK�l-뛖�_rYZ^D���%��<���螚�(�#�+y��Z[�w��L;y�|:^��B��@�/Lr���滞^dǧɿ�|W/1���Pu�Q���d��k��_�����[��$W�l��������NH��'�N(v�"��f��d�
k�¤�1��v/ �[���:�x�����|��ϟs����Eݽ�)\�{é�T�Afm9sp��\��}w^*v��j��l�4,��q����)߉t�������aB�П��>o��m��-�5�ΐ2]R����s�P�%��>Ph���=���K4��^B�w�t7�tԞ�B�ڮ��#�r�7�]#-�F�&5D���*��Ѭ�dr|F8�:r!D��yj~��}���!�OJ�ȼ/Wz�T�=#���'�q@��sl/���
y?���A�偷��B���R�K��*4q7�����:��1v���ƕ��T�X$�_��f��A�W�W�8nW���y�*�f9i{P�Nx���1����������'J���؂����p6�sܠ|o���`��F�q9~u)�RC  �֑���sQjrT�!a�i�Q1�c?�=ʁ]�Zff&��r��n,�`��p�B%��%�O����BE�\���2Y�w��05�J�񶜝�������=���}app��C]����D�D)�J'i(�����.���`~��7�1<��Sɤ�E(��4��L�kA�d�em�rLR�i /���kZ�G?�׿j�&��f���Ğ���ݝ�]��heO�^��{��o� ��؂v
}w���*�5� _�m��H�-��)���(@�%zN�|�j[���׀n�cp�x3�f�1v�b���GxG�IKK_]O���M�ӱ��	�i2~�=F �8]������?�S7��������v���\�W���U���vzP��
�����RV]jq��������KX"U���a��+�V\��r`�t�k��E�P�ADH�^!X�����a��Et��X���� ٣���I��LW�	��t��95��V�q0�b� 6��T^q����p�/���.��)�����������ͧ��R�f�@ٸ��U��0�{"�W������ۦ~�@�<�='�&�rwp��B�>Y�<�������L���uu4�%�	�$K�6��Q���ePc61��'�H$� m�TY6�+�3��X��Ri�o��}�����ǉy+ ˿5f��#�1
2� ��X��|3?[_��?N��lnS�b���2�\���������v���.8��݈�B�3����hb��Q��G�;��w����v-����x���ۖ�O ��f��{�c�K��V���T�k`�'h���zwrB�[����,��4�m�-�տ�� d4�4�<�]I0W�@�.4���{���%�љ`(pH��C�z���Ⱦ�ݺ�������W4���c����{���%#Be�[�q^��3�y�!i����V�UA�o�I���!3㙯8u��;��ؐ��ft
zMH�k]��5!T�#����>����k��F����nP)�N�y��ң��҄��h -j�	Ï�3�._%�7���<�S/��*l��?���٧2O��fs�6�ő��!� 4���w��/���@�%�k?Hu�Ob��j���U����Os�_6�׹���M���@v.D��!i7Ͷ����y6�)�����az�:�ms#���<?M�B����*���<�����,]޿.����@!� �2
��4Y�!����ͣ�d��N� l�_�/Y��)�)��-sd��-Ī�Ę��q)��Ħ8I���*�5���0͗[[�p+�o���ehs,�w� �^��-)�����z�m����nj�~Y'��PD(Qw�"Oz��aꨌ=(�]��9z�VR������Z��7�9J�3<R΅�>)�J�zBǓ��W��m�Х�U�>)�������)�Ȏ�	3�[g�.��.Q�7�{6:��g��1�'�Ye�,��A�M���r-c/�L�a0y�߂�>�F��G���ġ_n��Qt~�6mAQ����D?�|��������*	�b�Z�ǭl��ꢉ���
�^��c��o�#*�A���RL:s��8�S�@u���-�|��E�ڞS��p
/���3��Aq�E��q]7[��A�M�v�)��kt�Ca���^Z��?�b�We���G���RD�W�(G`@:Z4�6�a��t�w�l�1��g�g��edf�4�ձ�s��~���kKě^�"������ǈs����X���#�G�͆���de50�Y1F�m�*B��T!�����%���0��8mJ����d��υ�UL�_`��㬎a��EI���FMN�`��(9w?'�sj
L�:d�؂��b@R��7���_�7����g���ҝhy���;�:��ܓ&[m.���S��k�n�_5�R4 �F`?Y9�7�i�b�-R47���\>�Yf2���ħ;u5u�?��@k�+���&� Z�r |��&͵0EH;PuA�����Z�0��T���ۋ��.H	}�֤�z2B�Eӏe�E��{�'���k[���x���Qx!��0�Շ��Q�/L(JM�	_�QՏ���r[����u�c�S��|���!W�R�Fh[]�m�#�Ҙ��l�wI���_�%���t�ʤ1h�� ?�del�]�}j�@�OP��$�H�h�,e��Jt�d]k���]�;�k7��8���kZ%��x���~G~���*�Y<�?��k��k��6���D�J.'6j���٦��g~y�y� 1b��� h7��Z�H�P�
���l�w�]9�l�����p1�"�E
Y5�ڹ[�t���6�ق�Fʄ�[��4B�` �C�:f����,8��3N�D�h��{(7���O��#P�vi��n�Zf�r[���J�H�e/B׎�0d'��3&���H��tR�B�G ����d0���.��t�5�.�״�T�X�8E�i5�6�r��~b�����!�zX}��}�qqXt�d��K�W�A���-����i~�*�wY�<D��NzFܬ��C�P��9jǄ�'He@����2jzL����w8@a`��9䌒��C;�tk���9u0̭I3Q��9w�x�� �,'��^~��k<P��U*T���X�Y��d8q2K(5m�����j�s��[�#B�:�h�H�"����X��T�7,1S�T�����\�\������f�CA��H`��
�&cY�:Bx��\��)ae��'N4%�6<��FMO�N�`�Uu#8i.�g��2WƓ=Ƶ�J�O�2�H��>�9Uaw�˛tR)�o��$��Q�W��4r:,2+�Y���4[�_���y!�S�ǃ! c��:�]�Ǭ��%T4tɷ�FQ'���A����I�cK>��K��@��x(�h��v�	��73���&2�?T&���%6rj�I��n�?[Jծ�|{�>����ngy�1���Do�l���D�h��u��OΖ,K���~��Q��O�!Ӆ��Jm����SG�M/-��؁�:%@yL@����nLIu��4쬻�~ �&���op�e����~��|+�fV��4��{�Na�M�S��К�ȃ�����EO�_�ny���}���.U��weM�>eG�"z�@�>Q����{��SX�����yc2��%u�Xtܱŝ3'��n���Զ!y^$�hȈ��݃�lo���S�R��]rkS�u�L�����9��8� ��D���X�^���@�h��Y5�o�:I��<aYW �= !M`�|�D�(�T=�˨�*JC_0
f>%Kj.H��x�P��@��z��,���.�X�wRua��L�rG}�����lM�"�՘�=a�n��M����d6'nuSl������
h���rEmC/��$@<[�e�����h��w���B���0���7t�ӷ�s�C�N �؄7u�}�� v���>߹��µ[���p�D�a?f����u&H�T��и�Ë=R,cW���C��PΎ��Vfe�+aOpe�s7�SB�ZH6rn����'��	`U��
 )(���(���>��]4�Dp��]�c��VYX�F}b�������ڡY
*�Ky���
�9�R��,�B�QEU0
[��˂��������������Q[����K�&����h8r1�X6A��B1�WཹNBB����71i�e�9��l�ǥ[e�-�3�K�K��3M$�� ��ȯ%�����Q��wF�E�SVI��Ѭ=!��EN�7}u�w�M���״p`�?�N֥2�ꆕ�a$�S�<a�"P��ќ��X0�1���F%���]�0�ޝ��o���L���P�\އ��vl��D��y��W��-���ݲ?�Ǡ*&��Ҍ�0n�Zg��6>_멝��K����fRI��2��/XҠļ�=��'���W�������g{��m������~ �ďT��LO���X�h�)��(�k����O	�0���؂�vq����ШV����b���*��j&��8k3z��D�������F�WK��D3��%E*>�,����-6��������P���}��5�>\�&���BA�!�@�:��l�zg'jX�	�qiq����?�n�uM8ת�T��K�����Ǵ}3ǥ@!{��e0T)]pU�@.����{V�\|���26ă��4i/��e�]񝒠uJD�,Y�U��˦��t�B�
X�:ָ�q��c���T�aZ8����"u�c]^˘\�3�\{��;�H!��m�W�(=j����\�e�(�;�\�D���&%�^@��^��P'��W��[[�G���C��r��c{k�52�gVd���ߩ��Q+e�I��m�	 U��`8F��0��rU�r�tQ�=``3�~�����qupZ{��3gWs��B�n�#';T�⩞=�!�I��,A�ӈ����5�� ��_4� ���-�_����E��9M�Qy�x��VG~��� V%6�����i�BH>݋����]J8<��h�tSg��4�������Z�p� f����v{c�p�& �EƱ���f���P�2z[ 4܇�t�?��x�-l8a2eP�����y�:�b��q�AS�<Н��/o�(��|c��j��i%x]��N�3�0�.1;��
��x�Q7}t�-;�p-5����&��݌�Z�z�}d;�{���k��&Ҵ<��ȰRl��h�c푻���~�s�0]-m��8��A_g=���y��ސX�_g�@�}�z� ��\�@�so26Jz���u�LD(�\�rL��d�OB9�"����inT�&�.�f�������v�f+�cK�j�	�r�n���6���4�=I#%�wVj*�;�4�
¡4�y�1nX��J5�蓒�0��Bl<tv�v�S�5?A�R++E
kY;� �!}�>��dt̤Ri�������b�����l�a*ĕ?M�E�^Xu��U(o�TB�y-�������op2Hi�g�T=��)���r����r�u�˔�A,W��9�c����{�ș�����E��)���?��Y����)�2��޽
��ӫ(�b�hr~zBRO�W� Z��>�&�:�y�;�������#$��ں��O"� O����W��"�7�.t��A�(H&NꇡY��~�nah1�~����c-k������ǔ�ꏿ��(�G�h��v�Ńj���1��4�2��:�U;�2x���FTN��z��k|�^���w�U�,)X���7<����y'`���k��$;��M���Gߴ�A^�!t��6Mp����ܱ�l���eI�8"��/Q@t���L�E�rOPG�=�;� ���,�]����BRl�ױ�:���A�`#�gH��N� "�Ε\���H�!]q~?Ȓ�.̭nN���N�;WÌܭm��h��x}i��؛�PKN�G<r��-�����#r�@�&I��g�wHk��E)8��Ķ���V���D��˶\Z1Y�qx3EH��1�;i�������� !vTM�m���:�l�@�=�V��'(�Ք:���r���Z��o���T����c��&�o��P���@�q�Uꇙ��F筄��+���A
�8��zL��M�s��f��B	*���1(G"*�螥�g�@)!���ªc�m �҉Y��kay�p� A��UΗ�ҌL���ڸ�ej��:M�B�{(�v�U�D���*Qt#ߨ=]��'{������p�OX4b���c�&J�밖0V���� �bTF�wn��f�9����-W�%�Xh�>Pa�F���Ie�^7��6#�k_p�)/H��`L[�3@�#�P���Ez:Wj�~�ֿ����e�!��0w���8���������yE�/d4��rWM	�<�Q/���9:��-7��mC�e��Y����/t��NHEC��A�;l�j�{@���6V�'�6Kί�3��$��l�zuYb+D|c�g楬��:8~�	>��f^<<u�&���X�͝���>�Bh�X�S�b�v�}Iw�j.�qQ�/&�����ܣ2��8&�k󽊕����d|Y�l8D��%�{�ŐrLT�,h��!������^��W��cz��G�?���)×n�^ƠU�ٮUH��R���p�������y�c6�6,pٹ�%��CWcӒ+�_ t�[Le��&�5T��I�|[o��t�U	�!<���(�o���������G�*hz���ye>�N����@�4C�5+��N�j�]G��5�/�H�V��P�����,�ez[}	k���C��W��x+�����/Od���Tf�ңR{8o����-@b'O}{�BV��,S�	�{˙�+�ҫV�n�n_aO|��P���J��;{�Myb��f�Z������-q�c���ێfSZyY[��/��.���Ebˋ� \�JW#I*�3]vD�/�����o=�I/�cP������1,~�&e��!?3 ��J��ׄ� ��1� ���3D��o~-n["Ā�gS6����_楯F�_bp�D�H�w\��q;�Va����~~EW-EkV,]���G�G}v�-�w�1�� a {�� o�E�+`D1������]7%x$Mll����{���{> �����Ϡ�E���&ں��Q�������e�zv��/��O��X����I�1J�J(�K�eLۿA����]�~�*�&��T[�J����x������Qj~��5BZk�'캜O�����L�� �r>�=�(E���P����eE� �J� �R�>=���=	�݋���5�4bݫ5D�.iU� ˟|󜛶�4k����bt"���ګd���r�xM�+�z����O�%�-5i��ҏm��]w��}��r�$c7����i��i�Q
-��U#3��1�:�Vk<�։��f�#a����d�=��g��p${Y�Y(R���|���1WMΗK�M�O����ۙ=,#v�j#�qnvõo�R�*�NR-z��_�	@�����ç��*�Pe��&��!=���d�_�Ehm��w��7�ASvJi���fvY< L5�pw%X"�蚡�|,�:uwL�!;���k~��UHChߦ�Zk򡖽�PxKBh��JP dʾ�d<-����^P��/�����A��ژ-��n�I���8��G�A�{"e$g�Wb����x`���d���xkpW#�;o��.�hM52W����QT��Ycc���-��\h�6�!�N�l����}R:�?|��la�R�����(���9�7�]m�Q�9﷝�S��_�*(����.����짫OC�p���H��`	qtۇ0k�{�d���� �0S:/a£(WթD�1Mǐj-�|�UlD�Yh1L��4zvYT�!�<K�o՟�L�`� j��:Ǿ�[J�F�ӗ��<���rGe?_O|�����A�zo���z��>E6H�g��ܾ����`���q����<���[Y	���e��`u��Ү���{o� �5������ٵt�,#���:-7��v��q�rP�~�m�Q�.��I������N+�1�/�6�2��m�b�M�&JI S]n1�P�{�D�����Z/q�쌄U{���UE��rf3�2B��qЩ�@n���~'��ĂA1��W|W�I_fn�$�u�>x/��>�(�w���K�U��&>5`�q'�;���/?ߓ�rV^������;�R���W�{����h s��7P�ݥ����嬗��)��z��YF83y�֨���ff������JG�R�g�B�G�FX
�jV�ή���=�ϝp�����$�Ǔ�d�u��p��I�3�z�N#Яc$�/�ì���L��+����k�
nlADQ�Z���Ӳ7�Y�GZ}J�v���v�&�$�O|[h�'gܓᘻz@� �	�_��QK��*M��om�w�@n �r�4�!��\[��Zp�O���`�(�1}:�V��,�W�`䇴K!�7F=�k�����La���`L=�̯e	�>0�\}7]�u��u�簮�[c�D���l���^�T�|�--��U~�3�y���(���9�v��!�EˑԎ&�J���]��+���5XM%N.��68�`�f&�
�%�[��3� ɋ�}�״��D�����Iy*�h2��jՉ��L����9����Z��[&6��I�~�u�3l�ZC'Xج����8��?��GI���5I�W̟�Eύ��HG�����&k��t{�*����� �u�-{c��ѩ�1���+Tr8;��&|��*'Orz�3�o�,��������DGq��?����{?(��G!>��+��_A���M)یt��d��Ej�L{�&����h:[A{��;X[R��,-���Ϻӄu�{�7��/�{%����v��x��v�;��g��>H!�*���]GX���������QvP-�%Sp���CC�g0�m��F~M����a�:�a���d���8��o�al DoF���#����kw&^m1�e3���v�U��	Wln�^�IM�0<�����]�j.�M|[&ea)I�ʄ�����m�ԇD	c=�<��+���J߸O�M�F�����a ��Z�v(K�qRT�C2�?Yt\w;������S�g�G|S�n��Ox�y��m��˘�r�<�.��p�S!3��P�QϤ��v1[����dˀ�'AU���3���!c�$����^Α70�T�>�V��R�㉶)N���g��#�o��kZ��6��yc!�P}J�0���0j��U)6��%l��D2����S/��wX@e��/~�`�×P�T���3]3>=�����b�N�N� ��^K B����U#��/:d�I[�ޭ���
@� 5��"7��,��[�xg�=����O��w3�`�R��I#硈�1��R�7�Y�ɘ��
��ω:|-~�,�h8Z�;�=v���qV5��U�e�,Tb���$�-��3W�w�U�Qہ���e24�q%&��s�TU1��ư�Տ�yZ�6�N�d4���&�g��u=�-s�7���� �(XG>׹�7���h�;���\�D�,=9�" ��1��,�"�956��e��H��b��Crf-�jAl&^��Q�";6��m�e��fBT
_x#2�� }h�̣{f|�ڌF��p��E��F��7&�4�6K�?��*Q�.���A�
��,�2�/�{QT�,��G�Ħԭce����"H���*	�����eC}d���S�x�v��#Y��V��n�]�/]�^���O���[+MH��-�(�Q|�ԁ�6��:��ڔ��6��=�m���L�ظKk0��ڎ�r����6<WU�ps�v��w���A��[B��'�N4���f&D�,H�P���7�s�^�1V\$��lyxп�3��iy����>�Q�y�: ��v��YUp���
�$�#؞���]w���%$�4�;�$����D�D������dmY�~!�\�u��C\�vٵ�䃴�G�{�-J2��d��T]J�o���2�l^I�k�&҄e,eө�}X�2X�a9"��k�B�d��+9�U6�o?�z��r�c����^��,�(��E�����^�\Л3c�)���  d��ɨnw��n⬾*�Ew,��V������l��Ih�99Ͽx;����C�_�5<��Z�3W�boK�O�4g!Et����L��;�p/��*y����Ә3�� z�:pS����t��h��;�6�أ��
J#!P��H��'V���T�Ǟ(ʛY#�Ǣ	yp펶�AY�b�5��}����d���xJD i]7��?&>)U��,�/%��
E=IN�O
E���l~�=�������hR�c����Q�!��w ��GM�����:z�STח���#Pěȩ����K\=U��(�b��8Gį��'��F�
�C�C@���)6���s�){U���p�e'�Q�5��F�u���p|�{!��ֻ&9_j8˓w�L[*���m�s�.��"�Q�&
���eaޥ�ʃ�qߠ���[%��]D'��̆؀7�HWb1���erUkX���E�"}8�J��*jŝ���K��sa���쟨_-XI�Cx��!�zsw�Y���@��z�
z��.��
�����+>�WN��70{��H�����������j<���Qԩ�U�!��Y�`9Ck�����)���?�����c�^�\��)[�RN��݌��RGz~�ҒQQ���°�q�r�=���;��j-�<��	���XlV&j���U3x�w�2|�힯�_�.y৷��Ga8����Fn�t$�b���af�/"��>Ef��B0S��6FM��_b�����C�p����y��p�r�q*�3�	B�Z��������dE�o%�x� ��g�A����^3W+bti��:��8U�$;��z ,�������,ے���oH�;�XN�r����ӯ#�L�r6�1a�f�W�tj�E��I���ҖD��W#�C.tB#k��Hzg��;����EK�bDX,���~k�FɈOW:�Ø���F�}�-*�@a��v�́��4o#S�����3�u�8pa�c�$ٹ]\3ݛ��[ZA@���+`۩�1R��N �qG7�*�|���Q:�3*7����-wQq:n��I���j�b�UЀ��F6��;H�y���������O/�Zތ���'�?!n���Y�������i��p u��嗠��kSٙHP_Q�z�fp���/��A�#�[Orb��꒯���į|#jӕ���x�={���c��iKL�]1[ \�8��,�:�I�E,	^�H�<�}Π�y���Ś5`,���PlF~ew�h^��.����.M5]GAn��ud�V�(e�J�*��Ő�7���i��r��vA3�]&�3���Gk�SQ��x�4�F���F
�Pk�R�&A��̊�U\M֋8�݊��m�3b�|P�0� g%xK�hXP;\0=�Qҙ�5����-tBD�ixMMuwG��U˾zȘ�֏�}�d��l?���i4�l�k�9��d4��5v��+�hu�m-Q]/w�Nq}Ö���R�)N�A����S�m=�)tNA�W������
��c�B��_� s+*�8Gq�u��t'�%���9�=˽<�!hw]Sޤ��K?J���߭�q~�|�
�#�ղ�7�>�(���d ����T����ax�r���!���2)K'6���	����Z���N:�4�<V�a~�ߣ_�S���>j+���ӓbJ͊)9��=m ߞ �(x���N#Dp�z[M
v� �s����X=��Ɨ[4As���r@f0b�|��al�	1޵�b��87�z]3?c��|�(�2ƍ�99�ͺV='a�ƻS$�PVȺ�a��+ޜ؉&�ò�=K��:"��&[�В���
z .ov�$�̷{���P�Ɂ�E1��҆�7ߍ@`}�2s��l��s�H��L�D�4f�����/p� �Cog��ӕ���GHl�	�N�s� �@���K���#�:�D7LW`�q(��c3��;h�7�D�����3�f�.�^N'x�I\Ôv�/�G�4/䒍\��Bӷ�B.�u����d߆t��;ހk�,�i��R�kp�1�FX�]��	�B��`j���V��5��4�C��c�Cq�}�=F\9TOu�P-��W)���`�j����3��A��ѝ`�%Q�I�Ot�Z/��Z��oW�dC4J�=�ב�T�չ�Y����?���J��R��.}&d��&Ś����j�S�hg�~��$F���������jAj�ZSE8�_�v�;p�=p��ϝi�7�\.�Z_w��@�#�x1���N��J�e� ������鈊�T�gŷ&�]�w��6��z{a��ǀC�`�&9��t��8	�u�Ua%�H�)T�w�,j�Ned�E4�@���/V[�'1�����#�6�A�����WTU�!YT����J�)��܏�,VK$V��<Ț!�=K�� �=c+���@#1!2I;�h�/���#]����Ű{��5�/���<uh���J�H)0Q7|r��w�3�G����@/���	_�Uv�o��Eb��J�>�t�z�˛�{{������c;H'�I�A�$iY,�uy�q��h56qEո��8�3A>�wr���8>���_<�撛k-^�`M]f����ctO{��P�4����nW7c�bx��8V}�R퀒O�۴=�l�N���O�(M�&��92�y�9fL�ٞRz9�?�X9]Omt���F_��|�O5���pU�AѤO���Fʼ����SE��9�5m��*��U'�Z���:d6���3�O�Đ��T�jǳ��D�N뇲n���ȭh1=V(�S��ե�t4i�EO��e]��/�S(��[�r}8�ES"9_�9��\�m�S������@A�a�!����,V+�0,w��X�D��D��`Hh�tc�YOFdnǍ���W�
5�����������PZD�'�Y*N�-�7ŋ7�^6k̖Z�>+��{��lK�)7�.\�~ۜ�=��39|y��%f:�a�޿�l/$���$h��ۯ�0	�wF����r���J�5���ݧG;o����)>�^u�V}؍u�%����g���F�'.~�$"� �����>k��V���Υ�F���0�F>� V�k��*�0���ek=��l��R�W�*�N���#T*{���6���[�8h��	��dv�8[0��/�r�a�/F~�N��c,?�Nݵt�d�'� �k����G��f?Á��Z��O�)����	\�����T�Q����t���0#!��N킇1O�.@$߀m'�_�2�=(!��hے�Z���N]d��xz��^��F�������^�W���+�"U���(!�{af-���B�]'�I`_�id��c�k���_ܻ&%�2�:@���L�	�4`�����u�u��w�X�<��<�`,NZ��\q��ˌ3��Re��t��/>!P�`䞥KX��4"��8���g�f�0� : ��v@ao!+�O/5	��{Kcb�B�_;��/� �J=����|_���Q8u��.%���F���1q�_�:k��M��°�)☍�0)�HU ��مE�S?^�:�NM��t����֠t%���Tw��R޽,���Te�*� ��h�������V� Q�I�<<,�ڲ�F:Io� (�Ks�d���O�	\�A���Q�oݻ; ،�+�����jj�?��g��ٽ��LD銂5��h7�����.���7�՞���̴��lG��1<��)�;+F������g<��'�&�,s��&W=��� | ם�:�3�/�o���0��4����Ӕ/�@N�)s:Y��胪�����X.W-�p�5����a� ]�#��zT�gEu��; ����F�3<�|C�_5)�u�/U��^` �R\c�l����\��:���o��5��>�K��%��o�d�A+K�
����I\�iˠ?p��0Rk��k�
��
_������4��Fv�,(�o�7��j����A-Mp^��\b�$��i��¬e��iB��T��Ae@�X�~�E�?w��-�4�����"�]�Ót��	��؞_.W���ۀ0�[,�|�&�K��Y!���C�@V��ܓw�,��F��V�s�7�[X���З*g!i��5�*�e��R������6����k�3IU8L�qKR�/!�oA�#��U��0�C��tQ~�Ԛ�eFm���u�O�����VŪ��2C5��ݏC���. �zhe5(�Y�/�����s�B�vu�j���tMT����e�'���^����W50^1����{�q^UMQ��k�^aˢE�|�.꾝�;�4y�����p{~�΍|�{鄭���:����=fc<u9����J0�i~�x�FDJlו�_�����Q#ل��-^�u4����CMY�p��r�S�����]4^'�F��s�BNEq�?i�Na�#f��ԟ��ڃ��ԫ@�7�h���>o��(�����a�[	P+�LL�W��p�K��A��a�ͪ�@��?~�ђ��f�%�{����1LV;���z������	�C��Th|��%7��1���m�Y�**c��|o�u- ���yI��y�4;����.	x~�!���$��{V\t��plo�jki�+]R�<~�>��J,-��7�0�k)@v~�!�0h#L�X%��h��C�*�;s��B�����{c��$��8����ZVy$#��M��E�l�t����=�zK����Vl�X@B�s	�:}lx�sc�nI�+C��{��9��"��w���B:��7�ث�1GTbq���������N9�͐<�J�:��T�Vc����t�ǽ 4��01�}�_�Ŭ}�Qb�-&�zR��S�5��Y��!£Hؽ@�Na���v�Ի�	�=�&�Sj6�7���IiK�=N��
�@+�S�Q2U�J�b�y�MEܣ�����U<S)5�0S?x��/K�<�g��s�\�Kv�u���h�l���.�9�q��aH��-��9�6�W
R/6���s�(E�FT~��zs���e��J�y^ՄK���Mʂ��-����H=%�bC��6��#�6B���rI�
����j���k34E���F���?AR�Zx�2)Տǜ�<��-M��s�3G^��Yz�������V�9�mJ�IQw�H�鑚�}��f�n����S����������U}_K���x,��/ɽ���[�;Ac�������u{��w#+��_�l�����!�� )����h��S`Gٛc�1����á���k3���U���,V=��G��&�}��F������[�J#χ6��v�r�R���ח.�*}>��>emP��`��`�PI]M�*�!�'�[$笢aW'��w "Ƌ[˾ĸ�뷧�L���cɇ7~fv��J��+&���l�	{�H ;�n�߫�^�tԭ��B)Wd��x'��_���4D�Gq%k�G�l^��
�+�P�⢝]f0�<]��ĵ���~I��<C�K=�?�g^ib��\�����D{˗ >�v��(��������j5��>ͼ�:y{cD9�B�ʎ5��.V2��#UA=VlH���i2ʉQ�t��f��6�&e@[x���;V��}ҙ=��
�y��9x�R��|ӯg ��v�>�kp�"4���̨���1;��%��cK���ٮ�$}����8��̭������Q�ҁ��@�Z���ڶLX�F�35J*?���[#X��*Y�fꬣ����4ȹZ�2�`���.N����FjAľ��[Z�Q���
�פ��Ni7P�A`F���F����J�����H%��ߞ�(��Åus�/媱����������t�dI�
��]��>JD	i�ݐ��\`��c:�0�"5���,�<�7F A0~jŪ9��&}CQz��2�C���v�^ЛCV�x�o�}�>�5���f�߫~	Z$��1�*������U����K K�z3����F>�	��[U�}(��l��Q*C�$^��������&�˽��h;�V��t)� nl��)5l�0͍� �c'q#�F<�3�1���3�>�Z���q�&? ~M���l׫�%p+�~
q%������$�lVU
������c׷�x���T����v�:�a���	��s?<GE�$��s˓<�0��B���s����V��B��ʧ�32E��uЮ��z�d I-ԭi�[1� ��J��Y�,w���#5�h�{p��&&oIJ�F�@�B��3��N`OKM��A[/J����	3�?�n%�Q�:��oYl�oż�	x�byB|Љ��!�r�aU	�������E�(>��d0�4*#S2s�{����X��78}�-Z���,�3���{5��f��}�?����$�R��|��Cs'X�kqI�υ�����j5���I8Ѱ�U��E�z\�k\�˘���)�����q�㫯���e  ��-ۢ�O6&�a���tb��2�%¯�3�����7UR���Y�T�y������V����`v	��w�ʞ$�I�m�f�p�G�q\�b�C�' ��gq��7��g������qד@����?�r��<eN�}.�~x#	��O�cA
s+�K��Y~�]�mx�K��v��n[s�"�^�V�_o7������|��}�)0�I"���iX<�w����a���m:/\t��1��(�"Atm��2���J�I����Sta�LSM�f�ˣ�Tq,�$-;�[RP�b��):�!������pr�>���:%�(� z��n���sb�-<�ʂ��=���:�Q	�`�����~PDJã�9m���y������\�\Z��P��	��"Iݘ)W�o�u�&q'V C���[>��IX�]O:Ks�w����$�I�c��Zo�N��T8z�\�YҦ{N�̉*@p|X�n������c��ay�|]C�a
�xN�u��Q���1�����k�q�_7*T�Ox0N\M���Y��K���" �Av�E�9O����fe��u�0�$�����j:��P/�b��pc��8���2�Cf_�Kѓ�R���0�J��f8�,^&}ٗf����M,| h�C$_C .�ˀ��X�����W�;��6Z�(\
=�3�\�E�-Zs7��Ryq	`����z������`t^�iL�V���4g:����0:"�M��댾E'�$V�ZƑ�s.[��{V��"�d�P�����_z�i�tg�:��C!�e�,��"Rp&E��0)P��kl��t�]Ua��	��]����A��F��Z�����7�j���-�P�z8��$������bבĬ�G�
!��S���|����dEP�w��ČG�\yUm�N�M�y\t,��Fq3x�f�k켬w<����n?q����K��Y�a�j-��;ԉpן�^�!��Q��GS�]hH�'����*Zo:����G�`��ǂu�}(�=�B��������8X�)-��� ���ks�_��[�T����`O(���:�$6�FBh��R��l�ҌIIi����H�R�Ȳ,1"�vh�;��gC# q�z��W���:	Kqv���=nH�^�q? 뜐�)�|�(��h*nr�A���g�XLo�Ӵ�ئa���!f�i���يs�m�6��գ�6�I�����A����ֿ��'N�\"#}��i��/���bm`��֥v�߼�i��R�w^�F�f�Ŧ�F��������Kz9G)p����O*L/�����%C�lNR��� 2�����L�|�~��(Gٽ!V����;{���-�J��.<����ѽ R�2�3:�7�ˀ����v�\z�*�t%��ŦA��mϷ���,�w����n$��刱�0|�V�_L�/����ukV�*Z�b�LԀ�ޏ{�Ǵ<��]rp���@�q�Z���Z�C���f��	�<����g���k�;��1N�,����]J4���`�Hy��ۣ��ul'�G�>�I�ih�����B]�wh�n����2�׶�tj�u������)݅ ����n� �����[=�94��0����k�	�Y�q�����9\JC��j��ܴ��M�+gdx�=D[C�m��\��l��v��C����|����(��1�s{����O��E��6y�G �����F��˱ۆ겿;oApv���}��L�V3#���|L2F�W�z��ש���\[��
�ޒ���b�`��V�Z�P��d?n���5����~~�lL$Nr�95����(�2 ��E��$�g�p4|ߵ��	a־��h�7R.�Ti�+]��V�2L���"0�&�����
��I߻��m.Z�=~�.�V�����Y���I	sI�V�9��RTZ;1Jϓ�7T�xa��x<�a
�tѵDh�W�׋�S����']���%ۖޙ<�2e"���;���).�e��I[�_;{wz'۬���_�+<¼xͨ�,f�-گ������#�wV��t��}���=-�ty �H�ƞz$�U�6��Q�����L�C�6P�S����F^�<��T�ĦHg�7﬛��%��`a�ia�:�e��X��6vI<���>�8���`<Z�+qی��N���)�j���Ԗ�c��k�C��I��xn�@޴���Jx�5%�Y�['(�$�'�'�ԉ�ރu����u��8�̋���٬�`JM�2Z#�_4W��6%�L��g2Z�Нy'�=����w�lyAzz���s:��L����F��*���z��� ����i3߀�}���/
b�NfQ� [e,U���eP��z��cOJ���Vu.}�r%d�^�^�h�Ê�)���2��Q��ߐgB�u�Sɏ�|8K(��p�;[���$�ܘ���ˑ�8�Ƅ}q�ПS���%�F
3�A��rxߒ\�6�N���h-@:����Iu�E>ob����ҠgM�z��-��ciC�}]�N��8ı;ڿ"]���g]����DG��7���Ol2��x�e�K�4-"HZ���d�!v���e����OE|��PTt��1��q`�ඨZ�,*�\֓X����KEР�Nָ�x7�[/&�[��l��x��trJ������8<��y�$y��3�jQ�T���b �$SJ����������x|��}k�τ�!3+���:��t�#U{����3ge�t?/�pa�nd,2��4A9;ߥ�9NW��d*g��'��\��k��� �Qupq'
��h}1ĕ�{���/�gk���\)�^�iB����ޟ2�MԿMh���"�>0Yg.�[�DHY�Y�B�T������̎a��[_�^�`�7�^���y�Ѹa>�d��/�����k��|凯�E�h�񉨞�*Ծi���/#}й��w]����a�����{�ޑ�n�ǋ��d,�ݑa�Rv�A��d[�a0T�#B�Y��+G��xu����<��j�Oߵ�mu�w����)�cj51�63A��]�m1��
�ٰ�^���(R�׉��o@dE��rb}o����a�����MS�X`ށ�J���k���̸u���&F��(w�iֶ�-#�	�M��ij:�a!'<~4�Xus���+�e��ً��%XN��+��y}H5�3>=��)l).��}�C�����	ߕP�n(��N|��9P�3!��
�� ��d੤v@W�+��m)�YO����ޖ��d�hoZ0�+�c����8�u�ӱ&F�֟����y���X�fӱh��m��\���������\�-�Q�ޠz�H�b�s熢0��V>�(5�m��O =.�vgHHI�����${A�)4��3���G߸���_�/8N�B�c��~ֲ-�0�H�G��9�5��g*<o=��q�x��������:�e����IF��Q��\D��C4�[v���?ÖBJ.=�����\�nE>�#�Y����B,?ȯtiV�!X�Ѵ��Q'�ǪWu6��<^��ZB�y���3�C�2��D���=Კq����e�ڣ*L�0
�:~]��xH�E�����j�a�(��}�����u�?Y\�|�W���x���A�@�;�g�s�2�/J<�	�?�
�0�W��{}������f뚟��^��]��������{4t͔����Ƃ3�ի̕WYGl�r�#�F�7�
���� �CvO�l���3ĝ�R�;CG��|�Ò%!��W=mi�v6I;'��d8><���\��3F�Q��ի��VRݾ[�Dos8|�:M獻��o�#�O�bw�0({���%e��]뉄�J�tONΘ>�#*kM3�G��v�.����B�Q�\H����T��EΗ�o�Ed��c7��:!�!�A�O1d�8��O��3-Ƃ3p�aΊ�^����b���q�d�HȰ��4��y���
��u�����5�s�zB�4j�N��ĵw��&-��.�q6�9�{|~l�k=Y�w��%���.��E^}���l����H��Cp�9���$�'�-Zcv�� �H`�i�\lx�vz1�&,
|��U� �:�tt�-B�KDҨ�.��T�j�OlV�rd�1� Of��[P���!O�&�Y�)��Fbn�H\1O}��l����I���ÐF�DY7.��Թ�Μ�pn�P���E� W��?]ϸ9J�6�,��Ci�.Q=T��P�a�E8L�6��V\H���>	S=����m��}=/��]�wR?k�Y[l��Tk>�����5��aN&Ь�c���bY񧜷
���s��&ΐ,��0R9�
�����s��Կ�(�eŝ���	���A���U+;b����q�VG�����s7�.\�d n�?����?D+T���w��*��R��νc��(�'��6p�f�f�-}�3�b9%�:'G+:�H)8i��Kk�ʹ���������Q��'��V*�C�+PN%����"K��|VfVI	�LL���q��pd�%�䭂a������d�B}�4��o�z7��ɿn��ZIF�����>�;4�!��U�Kn����j@�n7��*��l(���=��!��6��m9�P� R"�J�hO=��m�nuK����[)k�|�u?؜��!�]9�.To�W<%~׾a�� S�_��b��$.�<�ҁ� ��h	z\B�Vb
��?�]�Ld���k��Hl�� ���(��N%�FF/��ȏ$���|��܊X�r;��{����L�Mp��bo��Q��9ћ>Q�%3��Y�$d�%KD��� �Y�6AI�㛿�S�������_5i���`�s�BSCz^�|R$�+م��n��x�=�!�'`�!�py�Y�YS��o]L��3ڱq�G�3
2BU��8?��T�c�$\(ȡ��ट���㜎�[żL�5,LБE��7?؆���s������TQ�o��z���=u;���X?�O�i�y�G�l ?1���7��ӠZ1\�:�Oe"�	��ݑ;�����u��릂s� ��๳�Z'��%�%V}[o��.2��{ʥy!�T�s4���L�hm�6T*�l�A�2tkq�W 2?�ڈ=�cR�m�ɺ%�x�*��Rj	�]�]��˭���\T�V�3���o�BT?��G�z�(l�d�6��_��{h�A�yuUW��,��c�Qݸ0�������F ���;���
��R�'"B}�!�����FI	����DT�K��Y=��rr^�!il�U;7D�pݘ�y���CG�h�C���x�7�3���7��a�?K`����q��JxK�K�j\�_ñZ(��E�7e�D}3�t�Fh%T0u̕k��v�t��!��J�U�|�ߑ0��z�����5��X�2 ��:�;�7r�ۑ/��䁄�"�����#:��a �킀�H�T�|Gu�\��Y,���d!�H��C��P��z(��jJ�g��S�U��<^�,�:��Wl�Rj\�ë[U��
`���iU�Xɜ�p4j����a*�V���6���O%>�ܐ�%���ս^B��v��n	�EBC;jB�>�Jr~��Wʌ*�U�0]�T�R�Qvvu[*X3rX�N�S��$1�Fe,+Y٣[�Y��c�c�ۓ��xJ�)��Z'�|~�[�{�P�t3�d2��2%r>�s��E&�*����D��U*)t�p	��Lj�%
kȀb��a9��v�/d��`!�߆�!g@*����H�tgk�L�����1�:��ؗs4�����D$�\��2� ��}s1,NQ��)��Is؞�8e��뎧�|�X��'�3.��n�wT��?��k��,���4�v3�X��{�^>��������$�V������C�����.Wov�f]~Y��T��]��K_���\�s�0��D�)�7�I4�Ox&S������G?��j�a23fwq��`xd�q�]w53���2ЀT[G�xk�+�ִ������1�]�.�R��F����i�R�2[�HU%w }r^Nx���
 �������R��"nu��3<�e�>��'xC�Ĝ��(u�Y���p$2�"�c����W��o�{!�[z�B�^�_`�I ��?B[�f���z�v���Є-ﳏ��V\&éu�֦��Aݨ�><��M�ư�`�`_��׃{��� w"^T����,k��X�F����^��bS(m�-�:. �b����/L�WB�ޜ�j�K�U�#ت�����F����s�Qx|7[ӜI��+ʺ�֐�s��I��5�<�����)O>LI0W��S��}�gE�|(�b������zān���橦)d��2�/��IRs�����F��d%��G��E��M��Tɑ���܊�A�}k>��3���+G@ rT�H�$�>a��Ѯ��z;Yoo=�ƣ�8ǽZߺ��1�d����?��GZ�����t5���@��}+��'�;9�?ق�t߳�Z�Z��ﳗ>������,��V��o��^���-H�G�Ȥ��O-���Zg�W���._��"����RTj{����%��gӣKy�T�27p�M�j�)`�A�	OhX����U�5���t���B�����@�SىH�S�D*�m�7׀7��5e�5oia&U���Bw�5��\��jh?�c�h:E�N���׌��W˪l�uT�.]�D���>�˼���`�V�կʂ�!v��PC�s"�QlC�=F۠6[��)�(zW��oa�h�=�Y��;[0/�N���K�߷g��������r�7��4����:6 ���
�C7�am��,�0�z�-��Ze�#�����S�l�IW׷T�Lݟ���U@�C���U�&"���{R��ﶢ����_���9�i�+�0��z�xL�;�ź$0˟T�:WD�:�R���f��H���o���XF �n�a�@N����CL3�δ�3#B�2�!U������G敀eH��������"�t���4�v�U0��㽏�l��F����b���i�X�3f{`u��Īۂ���K5�PW}P�r�|3w���XQ"���A�?^��IR]�A�v	�yI_š�%�?���s3�ꉽ��Nj)f�
[	��\�B<ȟI�
Yok�#����D�"�l��ᗬā�J��Fs?�ʯ��@�s�����1_�ٙ����� `=$���%r	����]m[t	]>��]_sC�Ox��p�^����P-`$��?���+�-���<�u�ޙ3p�+E�*/��� �`�7w�c�Z�8!�/�Ϗ��r�j��Q��qsRe�Ȅ�����<������R�)�ڤW�_���`��Ւ�v�-�\;�fN�6�"��B�P5tB/��dscDMEQo�D�u���X6���x�4�>[���x��ka�E�y���������� #|W�r�+�d>R=�4�x8_��*�@�њ@Ȑ�pS��!-5�1�(x`_�(e~�u�Io���xEq����B�:�Z"U�n�� nT�i��k�s��+Z�R�F�Ǳ�{h�S����f�з>�ֆ��n��r���sF������6Ә�ێRjH��Ĕ��n/	�wr�z��j��8��A؊� ��>�B	��Y(E�1�����{�u��Z�. �^�0ł���I�"�k���"V�Vv.���}���*����jz�'�oo��{n	t�zh��v}��m�H�����:�	�E��kks�F�~54�)��^��U@h�-��$S$�O"�lo���9ۛ#�CX:�o��Oz�@��(����9�G4����n�I�;����r"TŠ�H7KSGcP��yi��M��Jc������%+��i��'z�c�	��Μ:#R1�B5ًyS�'��M���qA��̌�m������ 4V%���{�y8*�/'W������n"[���*��mBҢ��Ҽ�G�����5���8�?�f`�V_��5�I���H���=%`��t�������·������~t@]旚�E�>�>-�#U(o;.=m���[1.S9�.�VL;y%_n.���a�.�v7��W�߸�u�kd��1U/�A'�������Tx#,l��X*����JJpM5�u������v�g��S���m��s�G�r(̦[A�- �sCo9@%Q}V�H3�h#б]/_�O1A\3����5rC��i�F��7�2>�߇�{�I�.�:^k�w3���z��Դl�UD��"�6���$���cD3M��Ś�CXZ�	-#ee���n�ꑓ��k���x�B�?�d�=ҮkZb���=�\��������ɼ�����p�
�+1����FJB��C-8yjx�J��d:zN��)T��V�~��D��-{G"���N+C����G�Y����`�*��9Q����)XZ��xq1� �3e�/*����s�$��%ܞ���/XI��.�l� eЯȬh��+��s��L������@�&�����Ƥ��U�B��|�r`X�ԑ�����_\T����|,��j���PW�Jc&6�yٱQ(1AԚ��$�#��	:�:��)�6��ќ�,�i��%��.��5�S��&ѽ�_.�<�73��M����+l��O̳ X�T�+�[���͌F�!�d�	�HH�-�!��GL�g��K�b4(��
�W��9�w5�/h���;�`�u<l��zY�c:[�����^�A�-�K`1RA��mJ�ǑZ��~����E�Ӗ���@w��I�/;���)�ږ\�C�z��Vf��"����^��mc;J�DS��A��-�=��˰I~B�{|tЎ8���e1*ۛA��VZ��10������F�*����`�/P'�!�Z=��8g�� �Õ#�!�N�h�٠=�xO�,�����x=� ;�^^DZ�l��|��ͯ*�7�4�E�2d�Jcso䤝5�f����#,�ӗ	�h��� ��W�|��#�����x�qI5��aq��{���� �Ő�(Cb�B�L�v��Ē�qq5ϟ�����O��f�#9���r͈�8�̯��FI?g3���9��x�7�팕�����5�(-s��]}�V��I�'��w�0|�C��"7zW�o32!u��Zlq�C�ՙ�����J�>����
q�	�#�m��?������.��v��,P�"u�E��F���w�v����N>��H��NY�mH��Q7��
���Ϊ�X���rW튟6����ɠȯ^��ģ��!9==�\����V�px���Љχ�u��Z�\�HX;ڐ��W��.�v�N�{1e�RD��眓Կ���Oo{��������u���}����b�8�L�g�;��j;�V�-a�6��W����/J.-���SF��z�nt�e�(YP������5q��/h�Xk��Q�������v�Ɖ��7�T��JקTzu��)�]���А�쿚^Vs5G"��3�&Y���KaW
�S�+��4�O�z��<������S�KL.FPJȮN����-��&6��d���4v8��1]7�¨�U�N����>ئ.�K���y�!�>��_\dGH~�5JU�_�Q����q�=PDU� ��LV��2�VI9���x;G��� ©��.¥�!:iF2;h��Cbu��Ǻ=!�q��0���Wt�uwJh`f�[�_S�1ڑ�����tq����3w���*'\7ݑ���J���WY%OD�J����	�>.A�������͊��ѝ��-JE���� B��v��?���T��Y q�j8����w���C�ܗ�[���:a�8��?E�줡�c�'p�:4�X|*��u�c$cH1�EWx�$��_Yv��dL��&<{�\�U`\���I�:�-�֚��w Ca�l��]��Ρ\W���8
�`C�:��)���b6��9�$��A���6L��BXh��.
�Di��" �%���<U�dFM�X}�v71"N9xɑ�*L."�r�Բ�Tm��D����!(�#R�ߦ00rw�m @d���Hz�%]`���S����dw7��t"��~��_��{��N��R�т2�ZF%>��~��F>�.w|i����%j�BP��r�:jCїxe�"��b @h�a�Y6kT#ց�!�x_��Nɣ*�wٿ� ������e
�'�׀��R-3�����ӵy�(��F��m�����"`���{�P��P���PG�Vw��|�>y�
a _Y�Z���l&��q^�\�O��b�#�&���CѓW���Ƛ�H�Hb��\�X�.~�짅z���Z�t�]����a��l��n�ܹnh����j�{k�� �?���!���aAkeeq���+�/i;Fq��͞$���NLj ��l�e0��p�	ck�}�P��r�ör���%K��3#�M��p�*�c��l�&�~Y�571 ep�����������q���OG� ����'��'��V6���II�n�W���u�j����P����D���^Mo�*�4u�����QA����L��3�f5�L�p4��(�l=��ٸX�\r0X�BO\4h;']�O�-�����eu�MI���p�Z�2��>�D����~�v"x�S�	�G�p�.�o鸞ԯ�=�-�?�rl�K�Zt̊;��0I�I��������'~�@�+=�_}� 
t��)o���Qa�""�m���Od�}�¥�}n*T��x�)=ku;�&m_I�+���݈+�	�Ԝ��s��G�z���M�=_��Q�����oi��M鞪y�:��/�<�!M�������$�DS�|C�(�$I] 3t�9�0q���7���)'�:�����Įn��n�3���#R�����5��G�8&9j}���XU�h"���I/]F���HG�6�@M��O�y��mx~(�~�q�0`��P5V��R��2\�:�p��#�G� z���/ק�Y�HC%<��U!�V c*hs���"���yb�Z=͝��&��!cLQ��'���쮹�����F��hk#�m�R�H�������=�祏S��˚���)�Tp�%���)�X�%E��XB�5i�d�6������y�h+&3!	XX�b�qu?p�9{���oJ��R����x���XX���F���)�ldX_�b�4A�%�"� #�I�U�TJ�_����mp��i����&H|�5q�z �s�t�`_��s]<�r���"�Ԝ}�0V1ӒKڥ#��8�.�:�X�p�^��<��kaf�P+�Z5�#� ̎G~�AqźL���Ӟ�袐i:R��=o����g����=�NO����%�D3�
|.�� �V+���Y�O�<ڈ�~��3��h]�Uz	��fCN�������]Ez�}�Pe�Jx|}`d�dAz��=?�f���T���:�Ǌ��4>�`���y2�&FY����f[������yN~KOO�3�ڄ_$�C,�J(Y�l��vi�&9B�iY��B�MKg�6)QV����pU�K����g����{���;�q�[�6}�J��1����^Ö��B�h��oc9�,`C\��U�꿜)Դ��-ۭCŮ�L�vض�EH���L��H!3+�=��iv��s{#h�ʌM���a�	]����J���<��a��9n��ȡ@�D]~e��ݫS���O��m8��&��a����2���g8`pmW�[��_�K�(z>	E���\L�5�G!ٹ��s��L��~�Jj`��~�7s�l^
�a�uh�E��B4�R��3�D�l�F�аѭ"T�:���|��t��$f�<���;���՚���&��@���޽+�B}f�B霡��
1;W{��y�Q��"�7u��I3�6feo��E��8.˧� �m���c�'.���<�UC�k��n�$T�����������>�;��6�¨�y���g���}��ht�.@�"4�8�K
p���K���h�&��/4o�Z,���� 6O&�<t��I�*�&;�p��8�/#�������D藯��o���ď�c����f�\[	����=��U=��]��Q��p�[��	n�ěV��j�3�{2���}�kD��D�����b����rf���l����p�V$h;3�?5����Q���88���J���:�R�#$����0�.�8w�&r$�� ��$����\q��AA�(G������V�⏽�h٥l���Y�2�FZm3vϭ��UBHQ|nD�^�\Y�
�Q����c��>yI�*����zS����a	�;��S|���`N*7��;.�%���75���	ֹ L���;��`�L0'�E��w��v��	"�䮔�`{ש�)�!���?s�6ck���6�ظYz�\�$#Ú�VV���$�;��޷����h��L�":�=S�uYs�p?�\���*����r��t��}�J����.����d5���U�	D�SO���/U:�"nr�
�f����o���bk�^h��AeW��<[4���	�J0m��M��LI�︥�Nfv���à����"d/��k 8���<̅�5�7������#���W��n�1�k$[vV��/@��w�#�a��AA�k#�Y�B%*%�Fb�N�w
={ΛS�a�Vwm���nu�t��7�]��^Q�~g��&aLן;�,~�w���od�o�ҁ�" ɍ��M��*�w(�˼��:峧�;��mV�#��h΢uAm����׭����]쏰����/s\��(#�=��NkG�/��L�(���a�H �8Cb��e�|�O����.gM�  �"��"�����Ix���|�k'<`� C Cu��!��g���ۻ~u��鰃S�\��n�2�XM��.�x�;�|3A^�m���D��b��n���%��{�Ź��Ԇ�J�ǣ��ȯ\��7�0�<�aSᴮ6���?�:}��y`��DDb��NE���ē��-�z�6l�>���f_XSa,�z��sl#ٔǛ�rm�$=TyH2�]$�/�<!�y\{��6��c�ʒռ���I }٣P9���%�����~�@�h.jȸ�eT.��f�	�qUL�1��G�U�/�������E�UZ�������&�~�U������ʣz�2�4�r���?�ĵ`cG}�Yt�Z�ix��Ҽ�C듷�~;+/f�.Pa�ry���Y��)�h[ء^d�� <�t�($V2��������C��e�$X�̎ݕ�/��LA/�U�FJ�g�c���C��/���জc99��vx&��)z��K���m�D�ws�_9= j�G!��~�Wxm���AdW���#��l����ϭG�����5�:����wZ�8�⊲�,*�5���%oS��-��;({	��9���Ib�%���j*~!���>ŚZJ���ɨ��ӣ�����;�"ne'�d��ro7�AV�G@?���e��Z�&JtL�w�}x��3IAچ�O��Al�!I�9�T|���f�|v����ƌ��WDu "��@}e�>��<t�R2�{�橰���uY��g:��_\���Y�u�d�C��I��/ד��A�+k�Qz������	ؿ�� �����y��&��{N��(if������hro�Q���\�^�K<%����n:q�B��UR����|�%�����ԯ�+�F����ͧ��������ȗ|��w�F��v�|��Ӥ�[�l:6�7p%M�H�HX�M��$@xaE��E�n�
Ez�P��c�v�bsP��9E�&����Z��bx*��^Ӈ��4^Gc�r����կ7�%��� �]k�i��3�I����i�?����T�NaR>|P��.��	Qx����[Hzp$�~�J�G(H�FܶG��*�(��4}���o�:��K�(Y� p��nBC��3��Òs�	՛��4��.�
^�i�]�p�3�C��H�����Ņ~W�)at^��B-��8�l�P��rB!M�̘�	S��+]��=�UOb�:E�.�ׇ�gK���6�F�]��>���a\�@[����|��P���o�k��&�XP�J1�G0P%(^Ec9�uG����� 7����O^�H;_��9��H���8QX����M��O-
�aI�b��?{>�͆X���RJ����'F��F`W�G躄h����J�bNՖϏ�}�:Ǥ�@U�¡\�`�Z���M=���4<j`_�OjQ���cH��!�AT"�~^\P�!��VX�H��.[Z�էꔺ�K�����W�]뢡��!	t�ܞ�k����o�+�B2��2�BS�'���p�s���i�tum/��"T�,�zM*��'_�	Q�/}3�0[g�~��r?�����w:������U�^z��b3=A�/��N�%&_\-�S�q#Mv-����@�Zun/�8g�#.Z�9V� _�Q���q�yޝͣdu��Ȕ;��=�Ӥ�¼[��`�^Jm,�*4���G�k��d*c`��!��Ht<٘��U%xΌ�[a3܆
��q��]?;�����(ƨF[�O���Z�%��tH��A#�g�N���*�d���a|��z��D4k���v�����R�����~��?�{<����=�=���N�z�"������*�ѳ��ReްЧW�S8wY%j��J3m@�^/��I��o�~�1�8�����3��x#�N���\_=��;� )�_���dS����.\*�n*f�B{�>�h%�����'��\�
�l�=���4k��w@f
^��_d��z���ϔF��:��nkP��L4�Q��)}�_x�Gؾ�]��)0�?kFi4�N�]��������ʿ:����$L�08�T�jg
L�Rp�����r0D:�`�X��c64�;>��p�*e���2i�����}�c��S\UeQ�Sg�v�1|��^sOY�EM=��t�`������ߥa�΄QLDq%�Fkk�ub|G!��Xf����2��XE�5t�a��m�u�W�_|y��WW�.Q����c��m�������.D��j`��✧�õ
����݄�J�p��6������Kv�O�I����$�C���JqUU�3��x&���;�rϢ&�Ě�!���(.��Ԫ�T=r-f��f1��<��O��q�h�g��T�%gMS�ۻ�:���J����31ҥ}|�u��ڸ/�s��񦬴ʘL�|#�O���t;d�IS�7�,:��O�G��H֝'H	�Vj�
`�e����V�]QFbS��b�O�*ÇYcn�3'�J!��f�[Xl�5��}�[3��c�[�w}�8P�f�n7�j�'z)�-o�4\���VMy^s� 2<�A��U^Q���� �|jq�;@��ɭ�5�7����YZ5֒T��,ܵ����R�¬ 0����[�*߅�V��u1��W��'�|�
Il�E�BKx�&k���������`[�a��J��yHG�;�*��n2U�+�o�j�ļ����m��zči�,!0Q{}&��3��^ob�m5/I ^��p�M��^�Te���t\��8�H h�ꕦ+��mR��y�ub�P=$?�3��������㴟�|>��*��-	G�j]Z�,�i����8��l'/�Z���h&ITJ_@����(��ryOሙ�8t2w՗� Zy��1�����4�T�m�ag���2;�P�:�ӠYw&��ϴ�I�+��I;'��
z♕'dN�`?�5�uZ�6����1��h�ȈPwL������E3R�ۆY��������&�Ý�B��'��o`:�si�H�>��o����pE�$�tS� ��h�n±&Z=Zm�^F����&�4��ʵ>�G�Ҩj(�ŜM�J}U�bɼ�$��'�ڋ5��o�g�ƞ��]�I�]7��	� l ��N����o�o�<��m�Ǫ�
�{#���宕)i0y7�#��5����4�q��*�hg�M��}��.���'@��Ɍ�Xk�5~��5�л��g�Ԧ�M����Tg��MQ5�c�jI��DR��鈠Յ����bO�~��t�*�����q"��3� Rz.ϳ�.`פa�G�",cI�h�  �)3%�H�A#_�E-��g�"h����z�]�'�MZ&�d'XH�=yw��g��(��I�������]�0��]o���:��+�] ���a��2��ok�<��K������F�K4�aҟհk�ؑ�9
����E���%�6���P����:
���73�u�~r�0�:"�rn!x����Q�?Im:�O�>g��]'�sN05����g���`�K:Y��w:��M�5��T�H��B=N�4S�����l_MP����rc��!�My}�f��kw���|��Y����5�9IS�n?�BY�A��H��SD�	�u����8��0F
1�iTsl�v�{s��[զGvs�ɐU���p%2@�+��we��:���#�C���� �� ���Z����w�r�w�M�sk�^�(�j�����".e���7T8/u��G�3"=�.��ys�"�}�v�PꆽW-2u������R:�5"��y�%�S-�5u;��G}G=�/A���t,�4�'�;x����I�ø�u$
��/]I*hd�� ����J��Ǐ�@%�I��_�'��j���T�!��5��R��u��X��3
7L��`���$�`L�Å��kV4�G�&����X�M?�M]x�8x�C;�mY!1��]<�oj�=~��H�:\x0l䩡Ԭ��*Ďpn��Q}�����gT�����K1ڧ^[��{�Byi.�c�
���SS~}�8F�OeZ'��rD���#r��*m���*�-�J�����=l��R�N��[��bY�D�g˲�3��a��W*󢋙̠���S�q7�,���B��&��+�����6���U�d���,�X���̄�w^+~㯯�W�(9�\��|��&�����)����������o`UyA� ������	t������Y:�~��Q�5޾�����'_�[�)�_�l�����u޺?p���TUв����xx*zq��x}����-�_+|�G�s�����c���~1�+^��n�ɤwsˑ��X
{�~[�����'���Od;���]Iqf�+�����h��'��'��x �{�	D����Uޘo��s��`_���eú���w(��g�q���w}�:�m��C�Ո#�T�� 3��ǺI%�XL YXտNU<'�3��Kj��bX ���]̃��S�)` ��ޟ_Z�!��h���j�̭;dJX��b��\��&��Dv	�2	�-9��%��I`�LEM�y�N���w$��́Q�x�Τ�Ƅ�fd������ΙT]��I�J���t�֔����8e$w_�!W����O��I��1V���%��@(?�5����u��7��ޣ��I�"�hh3�G8�b�(�|K1q�.kl������%�-�Ϳ��ݵ_9
'c{��˕�L�;��y�#͎��B��ʰO���$��M ����ĩ��i�� ��"8�y�'G:��F0q��Ϗ��/yXz%!֮~Pέr��S��@wƻ�o�g9|���SV�T,�����!Q����,�����].�p�RK��p�2"s2s-RW��Yh�eAOd��{%X�M%Y���(OC��<��l�\�Ù�T�~ާC'�QC�HN��uwN�V���ɞ~f��p�ԟ�����Q ʛr���n��xX���b�[�i5��a��Mhr����ۤ�I;��5��,��\���f�3�Lu�ǲN���p�>8��{J�1���A3��n�����{�<�w�퉩=�8̼�0_�z���5�5�/�������@�8e4Չ7=,YRG��Y⿉���ɼ�c��O��Y��Rrv�j����A3��ϗG��q���ʖE8���"�G�-%��M��Ț�� ��#����N�8��2�Q�^d�-���Lp�������J�a�9�U4�ٯ�v�?�̝8�~�]���'��P-�zm�w���X��	I7P�md͆�i[��''_�2�a�N�U2+�����_�.�~3��[a�<���Y�ͤ�1K����n�"`X-t��XL�m���(7Ж���$�	�g<H�A�`��=�������[�4�yUM��I��\]��<8䶭���(�5|�3��)w������o�����-���Ĭ�ZdQJŉ�Cj��i�Z�o0�1�䀐��d��s��w�nT�[��1���-f�F��O�{	��Q��N���Y��Q�rb�r)5�Rn��Z����Ɗ2N��E���a?�P��ߑ���{q��^d���hpʯ?@������ȦA�4���lo����X�j�J[��UǬ���6E�<��������\VC���!��e�e\}�]�Fec�q]b�h6�Mָ8��%�gEE� ?�Z���g�!�2x��$�*������˼p^�M�H�۞��Ķ>x[*U̢~�`p��:��R��.e�!��������m�}t�^3��Ы����� �̲ui�s��1����/O-c"�ߺAQ��L1����l��:��Y��&�:�g��B+"�9%H�p�N:����s��k���	~tr�M�L!w��d�fkU��X�a^�YK4�*o�p�(��2�M�����v3�.�+�n�R�h���,����/c�xH@%�5A� 3�:p��^`+��"<�4e�o$,.�P�hZK���ѧ$x�[������Ug�F�
~�N��M��C:�|(̌4��BT��b"rE�{�W+&���]7u5/32K9�&y��/��&R��@��@Q][G|�"�W�gR4��[�]�X�e�Is�_Uu�j�����TRؠ ���J�\�ޜ�V`�	��`�����fz���2rW�ߵ�3)>9_�Rx�O��$zU�q���w��~��ץ�R����qшj4����� j��b��c���s�P��^��P�J�����i~}9~$������H�B�(�v5�&q> ���jl�Vf��K��	}Z'(��Z�цɇ)pǞ��(�)H�v,�N���-1��d�F^)�}+�e���s��x���a��w��he=,M��8���.�(�J��V��S��l�K�5W��ч��n>�6M�DkC^�[fe���P�+aE�Uة��]�e��W���1�[�D1e
�W!�Mf��k��f�Vp3�Y����������z@H���/���I��TR��)8�g�2��Z�A�Q@Z�aq�Ut��UQ�RK���k!�t
�7򆹛�!����@Bi���קH�u�Hj��x���e������6Aҗ�kIJ���������N���C_���׆ʤǮ��0C���.e�i����x!���=�^� ��T��]�m�$��͗`P��?S�����n'd�+eN>ܟJ�;Y�B���4P�;Pe/WHa��-f�w�l��!���}
E��@G���Z@�}�0ip\4����12<V�t!M����6Svt`����Gj ��Wӆ3��-;�{�Sw��#@j�?�e�׃�*q��ɝ6��yS#�"$�~9��5�ǥ�>�GYcd{��cK5���О�V��تl�Nq9�0��&p,(i��̬;g.>�
�q9P4����� R攸����qOtf�H�����;kBZ�j�T�(pݍ���W'�����i
h,�	d�#�NcPC���WL��xjV��Q�ⱹ�L\��&���X���t���d���~�47u��I���Z��? ��m�?����
>LX��~��D|� �w)SgU�0�HfٝZ�t{0|�:iݩ-�7��i���Y,U�g�E����akcL-��v�|{��t�Ƌ� ��}�`�ڋ���W׆�����cL�?q������R���0�'���	�0��n12%,��w�|7֦
��1�n�<�8S�F�vOr܎��}����6y��JB��r�����D �j� L���b��<S>N���BjE!�ve��6��Z�Og��,���"t'��R���#��?��|8-C�2�Z���e�;�y����@�Q�-�v�M����l�܇�+VR��"�������ߣ�WB̵[����F�%��9���B�oZ�O(��<�%�V�qkS~U���T+�H��� �-����J��^�2H?k�]��9ڒ]�_i�c�p�8�DEV��¤��@b���'iI�2��������l�ǥ��@;���ȑ�@�Z,���Dp?P�ښfu��a1{�����k�ҹW��wϥg�YS��`L�BWc��*��|B���>~'T9�;���7D��lm�Q�v�����E�쉱�Tܔ,�9��t��
��)9�7>h��(���x�l��xƷ��Wը�/wCܝ�E�;���R�\V�S�7��gN�������L�x��ui���"�
���5�2z#`K����>M���Z�rH�oX��&��� �����9�`��bY7^�8����������pF�ӱ�3�� +�ᒒa�#?�+�yI�H���];L8Co���0�2bȿ��ll����t��y�T�c\�U]�ƣ%�H*��@�P�6�Z��t��H�
}P؃z3;c?�r�Wʒ�A�t?�h�V����Jnwb��<�V�7��6O��z�kIP@I�G�8��St3-�2,�J�l% H����.0*W!���{�ak��)�<I�J�}Ӏt�<��K�ׅ��4�3?a���U<#�p�(
`�1�Cn��E��2%���t��e�8���՝֨�;�)�&�+H|���Nd���F*���.�(�<D�Xw4X�0V2V<X����~ĺ ���ִ��Zy~mH���d~Y��.��o�d��g��p��y����ȸgQ�R[?f!��c����_���m�6z��(���
�;xLJY���E 9�I�hp����#�\fv>�h�~�M��q`���!=�n�@���ؾ�ʫ�[��6kX+�i����\Jw�]�SxS����ٺ|��J���}�Wn��~K�3������kEb�ah������J>�,��O�]y�U��U��?��sъD�N�@���-fM�aa��DM�!Z�02�襆�O(��;b�Du�Ӎ�%�:0�k��A�����n��D��Zt�t��2��Q��X��QTP��㤙�*��h"d!����,G�aʹ��KL��Ut���J�l�(ئ�7|C;ɥ�Bã�ǈU��'�����u�B�ȷ�X$˹J��`�WK�������R
�Jޥܔ�{�aW��0�%<~
�ʺ�ԝ�Z�'���3�sG|[wųe<�L�T��ǞfA�����>z(Rmꢠ;���@�|y!�U�t4L�$����X��	L	-��i�}�r"�F���C�#|���n�d�KH���bk+���:�C����hm��6�\P< ��a�h6ݤ�g�E%}��*TE6pÁ0X�J���7��3�0U������hsq5es�ļ�_����� ���Nh����
�6��ug!߷2謰�$P��+љ�ý�"�+�Q^R��h���Fv��L� �_�.?�O�� �������[��l�\h�F#��|�yΪ�A�"��^��A���q{{���fo��T\��pw�;}�8�U�Ϙ4ؖa)�O�@�8:�i�&��c��0�3�"���zB邽�bǤ��R�#b�@�2g&�'��{����p
+ȿ�;辁}��ګ��Ǽ��%����e<F_/�#`��U�IɮauG���;B%�냗�`���K+x���/O�;��{BHk���.
0���LC�u
!��zN:� ���`��Zd��	2}�vFҬ��;�X	��$G{�.��"�6<�鍤6�����
��vK[����^�9-���&�+��֦�D��|Ro��WR1�x1���V%���
�(�r�\��5��� �����=�� zhƟ�4,i8L@  ��\�����3��|�� N�X��;�T4,�T�1�p x�Dr*�U��_�γ6@;]`�M�j'�|I�ޟ0t=aQ�W��*��z��}�t<̂�6-�!"'�I������|M�?S�K}!���^@����ۇGF$��=JƘ��mP�z${Pς��g���n�}��Ƹ�·����\ߒ�����Nt[��]T�IJ�m)[D$�uO�-n$Ը���#e�~����&�u�t��g���ĩAe�2�L.�`
D�SqgQ��9�Kŕn���t٥�	�|�c�]�����VM2c�!Iq�(R��J�u���=��I�]���.+q-h��rlwO��)/Q�X����7w"��"��#����9�x�3P�����7����l�����$�za����j���9J%*�Rc�U\~ ��j���B�@���W�"&H�dK\ќ�|���Bj�"%O�9z航+�o��a1(,Q	��er�D�H�-�_��uH�[�f5Z��Y�pÃ$ؠ��%NO ��t����<��`��oi�^m�vF8&�(�؏?�l� �B@2ٗ1�����؋�[l.��V1΀��w�W�2D���Zʄ��C�s�c,Z�XEo����SW&�!$C&��V/H	�� ]�xED֙U�5��X�R�v)�¼ b��������'8��Dʮo�Gm]�qi��3��
�	��!�A���5����UF�FH���a7��z�����#G�I�u4�-��T�T��\=Jw;_ơ��;K�3��ְm&���+	�Z�7�L:��L9� ��N�ځ�oq�
�c��R%E����%���0ՋR�	O�^.饓 ���hFZl.h\z�c�Y���4T��� eh(�j	p��
��<u��qȇ����
�"csRW��.�L�c�:���7P�yap{��𷺤%���L��4�_�%��0�wL�P��v�[��ںhH�tJ�͢Edh����6�C�5Z��x���7��	���R��e\s�Ըm��b5�n<������U:����f�)�o����'��R�Kz���j��Ϫg��H:^�S�U�y7���1ko����Aj�DQ��U��?x�-� 5�q�x �b�3Nk�tE�B5Q���]�.�v6�N��>��� �K�q��� '�����|�H�Ϯ
�*׭�����ٰh���{����GԐ�+E�2$��!Ao3�@�Sޢ���Q五�o����~�l�$�=@�����i�XV@�E���C��7�f:��1"B�u�a�69�[&:
=X{��u�af�"0O4DÒ i����;�ܾ�-W+3�A�����_qS$�<G\8��}��]��	�����"�1�t��E�����`?A��{�(m�s i����N�;��o�6!�����X]��-��k~KzpQ�c���� o;�Ԫ@��j�X�8�l�r����֢�-��o�{�*8=���8�zyOD�VO��j���O�+� ���Qΐ?��۩���1_�x	5څE��g���s�Uڀ���0r*��_���h
���"�}�� QyG���i���4�>x�jKߣ��\�lz����4@1]����Hl��O�����k���^S*�_�w+�\Q�˿�!-K���+N�
v&�+�0:S>!�DѼ1d��	?�5�c+=�����Ƭ���H��&��|����P<�cä����@��^�����)�͂~����T��|Y�����P$��9�s�ؙ~��퉾 @"L3~&y�9hLs��I�4��w�e�*�`�\��?!�����)�r�7��+�J�kE�#4��tΑ��Y���Z�^�I� �ȏ<��,��I*T%ٟ�R���x��oSR�4sZ˱N�JD�ӁNJ�X��t�P~f�/��G�����~�m��@�@��ִE�z30b���z�傈8�K7,9ip��;Y`�-_*O����ä�dl%k�]�3���8��Ɛ=Cv��(�@3���Ckl���G�y-�.r�\(+�Tڀ��p(��N:?�yׄ���F�'��6�_�D�$)��n%8 A20ؠH/�0��n�l2���6�
�2���v�8�}gs�<hdq"���7BA��L����嘰gRv`�C̚/^aP�\?"����rrЭ��\��2�Q�:mH��k�����r�HZ���!�ὺ�V�"H����x}�c��.yE�X�c}��
$�ڸ�G�!�sf�����<��]azkҵ7�/)�ZSZE�]�M=I��� q�1�@�T�Ԍ���/��fm~�=.t�v�~��Y��d=n���nFq��s�`�&�Cr��E74�V�w5U*��dm�j�g�E_�.�������19�U�3dfY[��xl�� $��n��b�����eᩒ�.X���v̄�Ƞ��Y��f��o�М�1��sX�O�T@�#4:�'W��,���z�@��n�	n6H�a+�f4�U���1��ɔ?3��wxK�W�ߊ����),�
�	�_F�>W13\�yj���9��ݽ��}���?t���ɨiE|���Q�:������f�������Bp�)���h;d�tW�%�T���[3�Dq��3��ZT�Zt%(�P���h��?t"��3�'ӱw�j>h��ͧx�
��hp�3�~��t���5���:HZ�Wq|���I+��~�Q(���&��]�,���o!+uy{��L�w�&��tA��]Y�7�M�b���1r,�P:
�}�Dj��l:�'�7.�q5�2�%���ڂ�� �Y��r��7P4�y�;\��"�e^��4ۨ g���>J��F�yͭm|���|�!|k R�����P��a1�+XI@2��f�N�yi�1g,�̪�7q�	�|.M��%-�7���.j�!���8��a�~Tk3Z�e/(�D)��*���3v	�"ϳ�;,!��ڲ��_���cA�g{t��ځ�w����rYw��f�������I�-��J^�H�鱥��9����\�~ѿ�+n��wޡ���Fv�fW��I�e�ᴱ[*s$sy��&&���$[���aϪ�C��~v>�Bg��!�
����'���t!]��:WfG@W�_r��,���נ�z���j���v��yX�k��Y��+cL���8�w�ٻ��;As`�9Yr�AS`�������߿�ΰ�6�xa��f�X���j�Dē�Mq
��}㗈��,������Ё&4Cmh�1��Qݔ�l�p{%��xՁ�(Pw�O��/2D�]i�籺dI�ϊ��)����5�i*.�.`���6�]RX}�K�[�u�渠��\�p)#��EuU!���f�T�4�TӮ�����"�M�����^զ��r.�߇�⊭�,g?b���y����|
������B�J5�i��+�����H�^*kp����c:�����=Zp��(Epk��U?��,���DZb6q�.�y�d�=Ǆ�im-���B(03n��tz�U�rUN`��S��?�KMxiRC�� �\Ō>#�q_����ߙ�#¡�:�܈�ز>wVnɹt���y[��yV��\�T ���>��vyH��hd�~�0�y�����Q��B�)NIL��8��օX��c�У�v�������F�Д:��T��-��{L(�~9���Krj��_8�L���.Hi����֓�mj�:btZ����N�u�˶?agӢ������^��VN�ȹ��� ��[���?	k�n-�J��2���(ѕYz�>��
F�KՂ��o%��;r��(�����~c=/�]h�`014\k��ge�� ;�+t��<��	�*=����o�x��Ԇ����a�Z�	�Q�$W��r�}����]�L�m4���B,��v�洬�Լ\%A�h�o������c��чe�ȷ��>�_�A��W�a�8�: h�r� �U��/6t��(ϡ�9\�m7w�4,�?Tn�[�aӮ4k���/�LN�)�Y��"#u(������#���J#�X�}���V��=4?��b��1~m|(�.����D52whA_�u����;x���srV���x\@�
Clz�mX�0�Nb]�"Vy�f��D���2�#����M.�uuE��4���I~n��mR�ȃ���jP���S��t��4''>,8Z�u���]YWw:�"�
����V�C/�c���/|�n�e�fQ�F�v��^�!vFq9��r{���YJo[�7s����2�i���<�(> �� @i �����*߹e�"(j1s�؁�w�vp�9�7��SL��Q�u�˃W��G��igIF��{W�h1������^���-f��Ce#bR���7k��NM}���	����>J�j	��X%c��Iqt���b"�b[���u�N�������X,�s�;,D0�z`�t�\�D�/dj���i��>]�hל0�W{��k:H#|��'�` �^��Ͻ��xnR!��c�Nܯ�O%�"��n���{ɴSVZ��o�n�!�N]J�W�O��"N�@�g Hp<� �5V�g8N�ć�m���A��6�6�}o�� D9��!В.�0�w2�u���K�l��||"��{��Y �Ǚ�1+Q��<kus]i�.��-H���A��5��/�`�	VI��
�cmo�Ƃ�A�۳sˉ]���l"F��t�ꮋV���7��uQ��q2_m�mnv�ec�#:�Yp]۱���m�\���/"�#,���Fh��3��V�ŻA6�C4[�3@��P��^f� ��ԁ��\?��tZԿ�o�P��LLnd:��UA3��Ch:�
�a�3��'�ޒ>/�|�� ��
��B� �Y�4PE.�tCV��6�_��b&vp�6���G/ĩ1"���X:�d���*c]D����|z�;L�+�^��@��
��*?��+#�[Z+�Xxt�/��L573�Ф˦Uȏ�M��e<�"w�c3ٝ��TQ�����	�����S�z���nmQR� ol��$�{_�X��L�d���r@��bl�dk������H��>%�?QgS��d���	g ���ѱ3EGzȭ�G���'�9��]��Z���Jp�����y��B��Q�	E�v��HƏ5-��Q�J��~��'���7�؈��f>}	�0�>�TD�����i�TK����5/�`f����Q��Ia8�>c�U��"؁��n[��Mi�`M��Z��}d;����R���;+���Τe8�iῑ<������|9�t��1$�� L;��M����^�xw��_��pc%͸��@oEY�Y�'v�q���@Y./�U�i�F�j*���Fso�Z���ǐGT���������!�r5T��.-�0�'~��5�f̿@�w�Z��ilx_��.i�v���3�|;�e�����~���C�s�o"6�z��
��i���1��\��&���i+�&(�80c�]���~ִ�s�ٴn�,v��m���̈���C���7{#�d�v��;��R�J��[H$q��QF�,vw����{�7�a�S�y������jݕ�ʶ��� I����t�C/12Д�Dz���|f�A��SV�/V'�T���d{Rc4
�}�����k�=#)�y�m� ɦ��PC�F�w�w�F��=�vzzbb���պp�:
���A��$��řC"a4SeN��d�{�z�pEbWc!�C�2�(�`��ɮ2���(fG����'�q����k��>l��'��4�0I�pWY$���IE܌�(|��&f۳p5 �ͺ&�y-�[E��W|�
�,��'�!uhj"��� ���9�@���6A���\�< }�eb4|9Q�?�0zji0����|x��>�3@5I��m�c�hW��=#��bS@bW;�O��x4<���o��P!�d"}/:W �;�.��h�*낇�<Wr��X�X�.),E����m6��5�s��zN4V���W(j䔁�0��A�R	�<��k[ԪoJ�Õ4����v~�Q��t���H�M���6�
6-�����;;���i��r�<���*0�nƮ.�O��E;Z�t�Wv�@(�+ڪf�d��n��,�I�!�0P�Pmd�"^�	�{ݣ�CJ�"y���4�\ �7�����ړ�]{�sM��!�D6P��S^Cs��3�3��7FK�����hkǲ�5���m���:���_�y�X��lGi�f]Ա�!>�R���KM�[�'[���x�T�U`��y��eF��B*)j�]���deMv�T"����Ԫ�D89)�N�Z����#�J�e����d.���,a�ɩ̝W��t[x����A��w��r� �o�^
�݊��l���8^���.@��j3���-�|��怊G[������2M�a����A�Rl�,چ��B��8Q($� σw>\���y�4�t��6��vGMT÷Ȋ?h�aA��WQt�-����P�[�>	V�Wko��eW;��<��=��54�+j�7(�6��%���-�[a��g^���\)�P|�}�Z��	������@�}=���֮QH�����urû�<}�MD�b��/ز�ʺE��F�ں��V!aNO��@�^F�^�M{�]L���'/r�ܾ�c��|my	��&�;��$z�:N۷-�=D���v�%�a
�)ڑ=3O��1";�w�^�E[^Q�o�����*� R��}9#�T8�~�Dq�f��r�ݫDqS��wu��#�!/���rE�����H�Q�0�V��Ɔ�YR���(�F�/�s�"
�w�r�&�4��sci�{�Sl�	��=�	cn����8c���a�mQ�f��`��s,���S|���H}"Ch��g���c���)|�|܋�����K�0�i�)?�~0��PPU"���a��FU�?Ȑ�(2�t`����Ys3Ϊ����8�f�Nk�nE�N��g�,�o�2�t���K�m�"VIf.^"��	3۰��q2�H�������]se�S���T �qR�_qɢ2P�%�����+��xUS%�d�����i�pWq���kA��.<ɵ���c��2zV�a2�p�=�Uv&��'�ٗ�"�`2 �1C�����=;��0���>ġ�k��\��v	��5�"9��X��C�EȈ,���|�0�Nc�%�yw*�uB�Zb�Z����/ ?�s}�EN��zCI���~�y�ߣp��� �ǜ.���d����"2���$>�Bux?�����h�Vcr-��Hl��x�h����&Q���k��g�*d�0�P��s��:ͬ`.�<$O\jr�
-6܋���xh��nFq�?���\������g�jk9���t���A�8ݡ��nٓ��3j ߶�G+��`�1Lض�����/$���U���~��������ZVp%�����ìt�CJا9�S��尜بco��������/d,�X%cZsΎ�>c�9������x��}�'����CEy�8�2v��bAK�~
K��t�,�=�*mk'd��z�꯾���9x�k�CR[� (�J����J��H �B���Kg7�����N7c�y0���q�M�����d�ȯ���p'�4�oU��!ʟ��?�3s�<
s�ʦ����ϣ��
��),��|%{N�,�Y�c��"0�� f�v5�}؈����A�5&�T7i!���o�Ķ�ܦ��E�����$kceN�|�F��#
U�tj��*9����?����'���(8�g�_7��#,o�2��u_�X�`���{���U���h���r���"�3��nm1��5�D)6�˾�jej4�Dg���"oJ>,�=#���f�*
z1U�X�u[��{ �ן�:u c����[��~�>��k�ţ|���^'���m��E�2//��a?����"f!����HGMs��u���0����<�w��CURFt�C�1ѫ:,r2W��x9��ޢ�[��vV���I�Ϛԭ��>\����|��TՆ�vmI,�ƞ�F��)���ӫ��qi"_;5"��Z���dQ)c}"w/�Nf�i�,dl��Y@��أSШ�B�=K-���#����Q�����rhC�����d�Y�fk"y5O�d�2� @B7\Hnyq���o�0.>\��<��Y�^;e��1A:�cQ�� G��4�rѝ��ۂ��p?�OMLl/�y%��ԕ��k�NՀ �̹l\����%ͺAL�i[�X��x�3���D�Y
�u��I����	��	 6�p�f�I-e��K��([��4�:ZF�Ą���ǚӤZxK�.�@�p���E� �_p�5ĬkI�ɲЇj;�{b+��F=rm�L�q+(_��"�����-hƂCJ|+�Aiױ]?݉;���F��/��ܤ���F�˘P�ł�Χ\��Gp:�P���5F��8
=t�+��)�$���)JD��b���Id�����T+(��ݲ�`�HW��P����%�Z�.��d����.e��|h�u��uJ��u
��eY��/3��q
������<���
�dꄃ��rB����1�"1�)ΖE�S��
�����l�0��)~�Ylۤx�*�Y�iŨ�H�!T��|~�_~��xR�b�B�[h׈�?C	2�|�������%,�������_�ў�Av�At�q�^Bu�L�qɡ�)�d�V���c[`�zլ��rm7��$�a:�� -)&�T3و�Mo=�P���.,fV�Y�Ɠ
���%�rK��L���v�?��)��(vh�$
����k_1�؊_I��k)�S\�5T�Z�;��ǆ�;XT�b���䂳�x_d�W��̾�7�O�#*��� �wyt�*�g/����I���SRB����& ��ҡ�4t�%o
!ԝ���E�����#~�KC
�o�)�zI�:���JV"��n5��~�p4����y�@Y�ɍ�j���L����;.y6��	��X(�(j��ڞ�����N����/����{l�|p�����PU��k�;�h%�e4P�L�V�d����`F(j��i�b���^]�*���c<��f��� +�T�������]-�s&�D]��/���l�Szz�>�������s%A��m(�A};�W��0�Y���
蘝-0A�@��s5Vȼ�i6�����_%-';x��v}y���=�1��_�p���T;��+���>�.��/��ōbQ%H.����Ƚ��σ�J�[!�̩�	I�c��zTa龳���Ճ�����Q����cQ�^�-���b�'b�2�e�1�5.����u֟��kt4U_��	0p)7q݌p>Z���R��X�=-#�f%Ô��x� C��r��M���@�p�����=Rx�Ԩz�y'��2;Uj>��UՕƁ:�zo�&��RT��ϫ&��_�?���>�`r`���t��/�����^��k��{��F)],�	4�_d~���S���Z
��/����ۛ�����I�O@H��@���bG�����߷�8�'�=��zU��Ԭ]��f���8a�����$���c��K�W<�Y�2��F�?v��F�z=Y�@�!7�Kg
�?��@&`���/SR�t�G_)S���e+�f�)E�g��ģ�·}�����b�4OT����a���jB�������[v���dm�E�>R��R�p�%p��&��}�J���l��}�8)j�[�N'�*;�䓏ß@��]8�s�0�--�e��G[	���� U��i�HшѢ3��gm�p򙦟Z��YO�%�K���K���)�d�z?2��N�ؒ+�kq�u�b���31�K��.�-�_��DT2��<����h�=�[��S3nt��j����C�S��~{���Hiv�D����>i��͆C0�
Ԧcq���21��#56xԣæ�:$h���4G�{f_��ȉ��'��Z'���H�j΄$�b	k!�k҇u@sr���B�[L��iA�G��e��0"]R��T��(o�yj`}�������{�#h�#�y��H�W	Z����w���v��4��V�e[�=j��'$�@����Ag�enT�sX,ɡ?�j����VaД�r�ڹ~�����K�~��S�������o �j�xC�Gύ��.؁��/�5;��@�� ��G��I�I��HA!&�=7����}��vi{w�t�vso�^�H�'&��.�!�U)�J�]
= ����q�4�uS�ɇ�M忓���}��h|�Lw34����4�i5�˹�#�_�`[9��.��(�g��2�C�/1�#�!�IE����|���2��e�3��` �ξ��]��A��w !�hBͽ��<��"�#�l픦�V�Y��ߊ�ִ���@��&'�x8nk�K"e��p�ٖ��;NGE�1���|�u�v�'
U�4�t_�C��ώ�'�N�c ���(��W@��՜��g;a��Tf�tD���"��d��9R�,,����ɣ�M��T4)���rr�� ���A�R!r	e���V�H_h0Ċ�	Ѣ�a 6���]p�1��\cc�#�٪�`4.��p�� .����1EF��O)��ۙ Y���ۜ��\���Шx�H�����]�c�=:>�_{k�<y�G�[���%�����6U�� R �'Q!���������}��Q(��_��U�S����h�ŏ�V�#��RS��h��3�Q7�D�&�Z����JN���y]�����vg�Ee�gQ4�������ܖ�P$!=[�Q6d��G�}�f�9����� ��&�`u�ՠ��H�]��~K"� $.����ٟi�Z�i��7�cVP.��6���wxĬG'�վ��6f�/]�8��P�7�w���b���N��E���!�;��t���x/)K��
����P������1����F�!�S
�s�F�������+��uEh ��(L]n$��dr����|���\����sz�tT�7*Jm�+⺣!�T�c9_�&�^ȁ����
�Z��0��v^r����]O����c��6!+M��+I��c>fK�!b'p�7ʔ��rЂw�Ҙa<0�/�;��H19��2^
���W�x��6<N�Q�n-�bR���/�D�������)"h��}�Ȣ����k��3��|3l�����(5�W��a�g��Nj���D��z�\w~���44��!"���,��A�a�htjw�a6��9�3����<��A���9�S@'������1�)~I�|<�&Bo��$�84Z�c��ZYr5~E��A� n̓<x(n&fe���;jyǗ���S*��>p H��S�Q�5�j*���M�?w���t�J��}����*���tcW�]�R��=]ɫ)�7�v�P��E	(��������n.J-#��֍�oR���x� W�,6�������x��eH/�d����V�S��ml�o�h5�3Q�q��襦�ܲ�ޏ>>��r��j�N���Ƌ�u2�]q$���4]E�qOH_�����jv)N���ú�u��*�G�[�n�߼����(����7�PN館���t�2H��&X�D����#r��=���j� ��M���%$�Z��������7�<���Vn�"���O��>"B�),TQK`�Y����ư��.��j�./݌'����:�q|3���q������8��)���`�OJ��"M�{�ɧ6�RM����ءi?���r �<��_�(K>�ғ�G��O�Qʞ��+E@���Bw�o�l��J&%����z_��L	���ݺh�)�M,2Z0�1��~��#0��t�[�X�x���54X���q��y�:^��eS��P��(q��+��1"E�Ph������P���h���$�!�@�a(%,#S�m�}�/&�����7����j��;�z6u�XT�������^��O�E�A��B�O۫�3�C�#i+(U4�K{ɔ����z0l2+��Z�j��;�H�s6�y�}PE�1�&j3����%0�;�1��u����S#�����Z��pt �f'�#ըB���A�}DX�]~��Z#���!���o�ٿ�]��	�t�o���<|���
���g�����[%��!T�Bsg�N+wtr�dҕjl��^\R#.�R���+��7��6VU1�ō��D|ؤ�'�����m�Z<��)6ڙOU�$�UWںF/x���e!T�@�ip,NH����yZ+Z,	Mj������eŚ� v��#Y�qjp��g�V�b�`��l[���܈��{}k#�� �f�.�ն���b0�{g��9[Ω�mM�7Hs�1�k�'���C���w!/Mv���7y~Ѵ���ULkL�lR�E*��\��H��E��|�b�����%�ϻhtE�\3���Y�K�-*���a�����*��[���)Z\B��2&�O�K��������X�S����k��G"�.�"�7�+�͚�\L��P�i�<,���s�j�D@!J�M��׽d�KLG�ʈl����vђLa{�2�}�	k5#����"������5M5���E\�=L9F���	�De��ܿ_e+7�SA�hQfپ
cL��o$�O��^��m���x�M�;�����(�(��f��Δ�]����u>��]l���o��H��$O���G;(t�G�LO�0�@
��쮡6'ƻO���6��ۇ�q�2�� {�[<�_�@ўI���>��ѫ;Cu�{0�����ד���5�k�=V�	/P�p䳟�VzQ�t�Pàe$�������$:�o���h��?�����kk`!^���1���פ��L��r��:fn�qZW>Ⱥ� [�  @C6�%�0�f�WS�Cf�¡.i(�����Qu��7�v�G��K�e�ٿDT�X��߭�FNm�>*�e�A��@�a�!��JB��'hO�uӉ�sx�0�U��4%J�$��N�f�aDM]1��+�V���,�DGC\Y�Z�ub�_4]�N���8�,��Ƞ�Მǒ�Š�����?��?�ƓOݱ���[m�d%���t�	�`fS	�㒀&%*a�e�
gW�Mx�(���&��1�oZ����}�x]��jn0LѲ��E���	3�	?j����[�%ݝ��$� ���:���썒� �*i	�Y��9f8�د`��}> T�c���7=��ٸlva��c5|۫�/������΅�=�̈́W�3ş�����I�����	�;9����� �c���]��1�5���X�\�;�����F��g3�!��~M��=��D��LK���QZG(��gk�Q�Z�:���{{��_��!̆m(�k�|�$�q�J1�t���*3�ʠ����??����VZ��lЄ������ wO�`xB���-�#��tk��v4ߓ�C)�(��*�o�����x���=`k�#��"��t㑾0|������[��d�Aj<�uk{�`�-�*<,�恥��'O�*�\M�}qm�h[�G���mg��}g��-h�%��5\́Z�+a
�>GY���Js�oL�,�$��M;Ȑ��Ox�����l9����|��.x� ����OE���萛7Y��$AQ4e�A��a1bag�#VXI���,����p�P��,A i �m7�~����/]k�5�͓X�CU����H���y��q�la�\�q��8�,�l���|+aH��@`�J�����s���hXc������O ��`�� �['d�#F�3@\VB#��r㿞����?\R�/?K�ګ��`V{:϶�`Fa��ʺ���΢A�&��ތ��
�lxG+�����sL�d2�����햽�0�[�4����NߏA�QY�).g	��x v5�د��3�OlP��D����c+�W]B�jr�X�����{��Xp���{a��y�
b}�ײ BU+M����()Hiz0?m��d&��y�u)P��A -��������'�X��"i��\�y-����q���E=M�hu�<�I�>Y.�
~�`���6��b� ��ZT���e�^t�'h�p�ϻ�٘9V�A��7� �:�3�hG�
G������Dk���x���߀G1����R�7�/�(��F��%`Ɍ���g�P�[ڦL������q��
��^Bd����<��3��M�6#f|Ǻu9<0����t8�u����ꢼ��w�N y�w�~B|1��Y,�7�+g=)����	q���dv��J�/��(#��|3������j$l3�8w8]G�_�����(�M�1��!���t F��N��3s9B���_%!A騢�7 ˮ�4�뮟n�k1n	pϝ��őe�aA�Aq;vg�O�3<�Cn�Tn{��}��Qi50���}��t(+�Vqo�2�7|�r�Y*\��J��0F3p��#�����`��:��K�Ь�� �b���& 
Uz���Cf����D��F���T��Vl�������ùJ�G�fH���F�~:H�>ۨ��l�jl���Ë�������d0~�8k��'�S��QA()���$��l�_<k�b�/k8s�}�M|_뒋���(���/�t�/G5a<fP{"�i���ʺ8�B�7+!8���tJ�3F��K�qǅ��r�*��w�L��-KVNz���Q���b�e��ۥ���5K���{������.R�0n<v�%p'�z|�8��M�� �*��V������a� �%�:�:a��/��]��Y�Oc5��L3��,�j�U*�|���M�J��n�866��76;l�q�ѝ�>q^�a�p�W'z�9W�;��/��(h�"D���N��d��L��l%�H@v�����f�G���fΝ2�e��݈����<�ͭ��!������La+T�}|�Y��;�"�ث*-����8��>m'���h,���H��K�_BQ����S�\qr����҉'%�o6�}��N�Z�qް+��C�8��$-��hbe.r�U!� 5��j�\����p8I����
�V�V�$�����Eܗ6�1���F
Ev_j�����z��Xq��'��L�	3@Wp4%���w,��Ĵ��^�Br_x|b2� �7km�]I�D)Oe��O!�M�Y�E!+����?��W-/���||��RԒ��غL�8���$o�ʨߧ��ݺ�C��e���暭�m��,��b��#�fO�-��>j(}�y���\��L�(a�F�E��C��S���(4"W����b �����B�
q=�W��d�����/�Z�'��ʂi��ց�:�ِf�����T}�ʠ�0b<�Th]�A
C�����Fb�$�'V��N4�(��8���,|C���~�n�>��m#tۂ�ǈN������<�\�id�Αm�f[�Ц$�O��������S��P�u�kY	�I꛰۱�i���/%ɴz21Vg�G_R��C��r&�P�`�����f��A���⤗|KVЈ|�-��H}�(�D��d4o�=�M� uvx�s�����ܨ�E�F�IP��$����Fo��a��4�7�Ǐ���L|�. W��e"���VZ���.~Q�l��9�st>��b�l��_d��.�g��Rl���4�ŢT�{`+�l�Nx���@�(,��w;�`q0�@t�i�1��p���[j���[�Y�H�g���2���ÿ$72�L⛫��j�2����dD��ߧI�^�!yc�)��g���'XZ�
;p�$[���-av�e/8ePR0�y��:�r>� �%�\��.f��'�� �exb{ə�ՒiIl��M��v(S��#V�)f����rMLK�J�Y1���*�����׆ݾcCR+�@��*�ߵ�796�X��<|���2�K'楏�F�m��%��GA��$k��`��k�t8:Tœ^�a��u�ߏCJ^��*�����]��/��v��#^�:�x@'��F���Da�X��(��xv�K��Ȏ�����3����kD8|Y�m4����������	�"�{6�Zćzx�����������"{k�#l�X�L��7��H�C��k��3�7�cc��2���Ǥx{�;��d�\/�/4WV<T������y`��TCW����&��Rzl�9���lw?�Y��y�t?�rO��?!���9���IN ك��s)R<w�
��{���Q�M6�Q����L��2��6J�=�̍V+#Y���p�>��s���oAD�6�h߲6�Wk��؆����w?���k��q�`�w;��7�ös��T�mtW����Y)�l�R������o�j)~��d��l�*ep��%?s��H��7�$Mb%�tX8�J3�.>�����;�����s��_J9ھ�Y�S���(� G{Ď�i��c!�"'�uFJo8�O�����%��ޡ��y�2P̱6�53��ぅ~��2߻��SE�)��j���׻���
V�z���N���A� ��BH����<ؠL#�X)�ݨ��[m]ϕ �M�2ڌ�I��zd�(��%X����/CI���}�K--���.�qb[��`nj6u���g�b�p�����.�}/��$�ĸ��q��,R��\aHԜ�D�'+�`������`"Qn���`�B�:��.r��}!�f}Qt�q����.aHF�!t]�Za�i&Ա�خ�L>����lp'`�y&S`J��8ChA�n ����ꁿ<�)$�R�p���7$�.��~x�a�f�3ʵ�_=jx�T�T�oٖk^���^�`X�F�� �]Jwo�� ���/���V�v�2U���2��=�u�&���TwD���K6�B ��� }�lZ:	%�RΜ\���-L���Y4���~`-�dRv��Q�[�+-����D�;�rm��`q���[e��k�񋯐����
�����ys�Cc��:�i>H%_c+PX�F�8��u#K&��3�ԃ��E^�ݵ�I�X;�ğL�����i��#�$l�1�)���E��sc�f:�&1	��9�&���ǌh4��W�\7�����m$dԥ��"g�:�(R�HV���4�B�젆��/\>��$##�m�LgtÆ.�𒄅AɈ�}���L}�1ߢ����k}�(�t�Ss���-�U�F�g��j~�#Ζ�Ȩ;���w�9�N��Cr_F�<�����)��G��r�UjT�V�8����,�L�<��v��'MP��<�
_��ӺXv8o"?�S���1?)�S����(ե�zg���>����V{A5�pb�p�h�@�A��R��-��R��U����ri�t�E����9�9���,�,�V��1��m&��C�u�J�8)�.򻡀 )Z�֌����dv
!���gz$�Q�&�⽰ßє=�'�͐�띢�t"�� �6C�e[�(��&��q�w`yekZ�h��u� �� �E����r�J���L1�ƹ0�]
�Q7�|��g'�~�\w��T�u��	_ X��P��ޑ�:C�9�8C��Ba<��@ 1z�0���֕{'��?�d��4�Y�/2QV�NI���*����o�[���� ��ɿ�t��!7���FX8 �X��(X��YE���#��C�9i�p��vy<���@Q۫�ѭB�Ki��
H������q�ۤ"��NKr.����m�ch�"ή����_j/g��*Ҕ1a:���_5��cF�'@��i�j�����T,67�;��)���%�y7�:
4��Mb����ZϚF<l���'ǈ᭼����>�����Kv��ry��jT$�yF�&(�5���{~L�@�����uzT��-��y�9�l��/7���]�)Ӗ�l��%m�:i�t8'��m�C�ǐJ��L��KpȄ��f.���C<�6����w�D����U��E�5=��I�ѹnSEh�u��K�l� ��3=��LP]���U�A+＾�RA�5.��x�Pk��(�r��;��E�@M��.�6S �d����S �"��z�� �$�k��}��<I�����"�'�M%�������p�D��k�|�p�ދ��� �#%�'d���r��ڲ��~���f���U��8�j�ߪ�Ii��;��=��#kcN�ML��FU=֡Z<qiء۪�kB^�g�^�C�P�T�}��	/Tl'H�(�ASV�Q�p�4�  �g?���:a���vG3�)GsIɝ��xm
{d%]w�T؟�+��[�G5(X*�n�]�SŪ,?��5��1pVS�24���%�m�^/�	[#���Ӷ�prj�Y�Jㇱ>j@Sm�S4�XnѸ/XNӥd5L�����jG3$B�؏�Fh35-�������JP8�Boj�IM��V�r*�I`gF����9�S���X�d��PO�����3�x_%�ȹ��y�[����!V��k�fXv��� '	��  
��\c$�v�)ũU%}	�8�:�,�_��$�x6ɰFwє28Gs�1��pz���u:s�@�����Al�������k��%�:��J�D�fEo�d.x�"M�7�@-�pA����`�K��\=�s����Q�"���`�$�*��5,"���.mD�lkNt�#i�V�jpYN��9��rÛx^O;��A���E}J<!��v�1�T�
�<&VS�KѣI(-ƿ���>\]4�_���.����^������a��fK�ْ�AՋc? �6�`hh�(��8�(Vⶕ����1�(ȴ؁\ঝ64����O��/L+m`2$��R��̅5.I	�\��~��5,�5՞�BN7"�e*������*��/�_:���-��t���TIp�0��q3Oz�G�N5F+غ�<�x"�����D� ���H�F����x5]�j�$��t˿�Q���u?��}�v�|c�%�	�C	�ۼ69���97˟F��
k�^�5V������@"����K{���~y��c���Ê&��Ŷ&��4�^*1�ss"i\:�g���=.���i^�}�fc���6��N��B��o&�_A��%E#J���	����w3O{蟄]����IS0��6���q�j������w���8Ž�b�P}６f�B�`���<B��g��Q©��-:L�1w��c��k��Ċ���*�ٮ�[5�}Gqd�Td���+D��Km����	V���[ԅz�m�K%��uX�|�A��%rId���7Ȱ��:]��W�e�H̎@횄��@@	?vI�(���E��C0�'�i�<{�I0�R_���7NY��0�G������߉��ǒjN*��dg�W�p@]ښ�MR�V�,�a���=�P*�!�_�H%��\��*K2±S�l�)6�o�8l�o}��N��zyIdl�dB�R����%��Vl
�����+?���D�r��J��A�b�ΡT�~K�p�/7��s����QF�6#'M�X�RE�K�2��GCq�gq�$�'J
���J��6�o����	��"
�X�{�J�	ɴ�j�Q���T��]����#�W�����Mu���	�1����_z��c�La�G֢?@_��S��<�j�I���w]� }_e�5%�&�e`�X@M`�k�/<�q��Ѓ���[��Y�$������(x~��$��K��bF�q�����\��C*t���)�<2�"4S[3���fMI4���04jM��<8����\}I���7d�˔R�S��_&��\���=��2��X����j��Uf�p�F��!@��$wzSA���qTw��&��%m�̍H�����3�r���ߐ�I#k���3QW+0U}�ȓ=t�����6,�ό�1�W\!�ӯ��?�5���)	X����c'�Qkgk.�����NKk:�`u�/B�f��4H��y�
C�j�d�W#�M�?�&��!��9F�0�1����Y��U�5�l*㷥Dç3�K`@2��f3\��x:=\��v��?jH-6�U�w���3֡�)A��	�����%���^<q fp8EJ.�?��Hbu�}�|��j�_!���
�@� ^���:QC���Z�2(�<"t�-�T
	Ϥ�Ր�����ȩ+�?[w%�g�]�E��%D�}�TJ@j�A{��c[IX\c?���rsB��g��p>�D���$�ഔy0[1�cO��m�G0�]��ӱ�
Y�P�܀h��]�ւ�-|��4�P4@v���4�H�q�23�C������2�hs�mb�?ms��s�����L�\P���(����D0�����d�9��]|�+���(a��:a*p�0�ze|�`+Pi
�VK�d���ɲ�B�� �6~�� i���C�"d�k1�B�/V��߽a�IYL�3���A�:WFw�8!k��FUBDe��S#V��������6�0�{"��D�Nׅs�6
��32v���G���T�괵Z�|:W���D*��6�������p3c��<-��P������G&�"ֺ�s.�k6������vKeD���:���1^R*��ۧOmug(�*�e���$'w�:�|i��׼���Q��*���*�:�p��:oɦ�����x���s��G&���/"���So�cYp�}V��(������"T9�2	](����W���9���H�����>(���VD�G	��|w[��B��Yٛ�,���E�]�ă�B&Fv'NP�S��x�WQNɐ�Ǵ�H�잯������&�r���<��J�A����W�dѥqr�[��Y2�j:�I��D���4BG����S����>��8�`QR����#LIM/�Wϋ_�V��Kc�R?s�X�ł.&H��_�1F��WҵTZ1U+�G��z�h��f2�H\�*Ϧꮓ�W)d��^R',,i�e�5��,���V���l�j^������8!���+�G���X"xeߔXn+X(��,�ͬf���M�8�#�BEC?����p%�zlܲ�`�;�N�T̩��7 ��PJ�yCI�pGz�]ڐ5�;*��$�R;�3��]��xy_�SG;�W�`F,��E�h�6��O�[��M�a�i_(��	���6���R��'�]/.��t���}	3��r�<����~ hpu2���RW$f"L5����U��*q1���;��J-����1��3'��"6؏�U�7F�#�t3�L��v��(�'Z�M�}"�ɱ�-�Xؕ"��D�U1�C�\�l|)�0��heiL�������%�u�-�=�J{��b�_Z��d�"qFk�����We�5P��z�̋���f� �^�<�\k� P[S� �׺��|_�.��]��^�7t��yD>�#[?bP�o��]`�C*ި�YOB���P�1���R�\a���"��7x5��$�|ӳ��N���4�(a{!�v��C�98��(��b�O�>��R��э˙C��꜖�*p�@N[9߭U*W��~�f%{�|yc��~�0J$�h+;��W�=a6�vZ��qt�e�[S������~OE�Y��gQ���ɗs驊Ȫ���*W�0�0���D~���e���ˀ[�1쎨t����T�_"p��V������2i��J��,���	$�����]S�������̼pՠ�f�e�e	@\�We[#�F�lвc8U���j�3�':�,���I|ʀ�j�eX�W]�f]��k��bj��+�g��?���!�6��WZ�Sۀ%�@�j��S_Y���3�fv���j��uU��ￂ�mW�w�r�E�@|�����S��[��
L�!ߑ��T�y���9��'DO�@1�>��qho%�Bً::����n/�̓���b>SFX@(F�Z�GR߻��2t�;R#�sV�����,M�h�8�JjȪQ��0vxXdhIL�:TB�@��H�h�?��%�q�|�QW����Y��mʪ��ju�ف��p�J�ћ��V���o��>�$'���*�Z��$@��Dl	-#�
��B^@U�6o��b���ѝUC:�c���f��[E�\�&�NH�����(��_���ʈ}s�"�e�GV�Hh:� Iϔ$/�o
J߲�ߵP�ZmV������EUĴY��qѢ�����8�i΄�a==��4�!Ï��V�j>�`M�kB	!"�4��<49���:����(Βl�n�C�Y��Q�4i��;]�/2�;�K����s� �0!?$�X
i���Q�2K[ʴ�k��q^���l������j6�LƱ�k�ǵ@↘JB|{�T:�3U�䛘G����݂		rP��U�V��mٸg�����m[�F��ږؼ���jJ��c�����!Ы)��]CZ��ΈH͏"���h�.���8>6���=S�2�!�d.W���m����I4T�@���y\��4H���Da6�<�ka�>�!A��q_i�7f���#���e�Wm�QL���� [(<ijB.��+@��u�U��ۡhExF`����y������t�)��\�l ��+ 1��e�6c �S茦�Iͩ��7g%J�C�脹�n@!�<|���ӷh��\9� ������[ڢ(q���`'��*�N�J\�U�)�Κyz���eQ�kr"����;oJ�]V�-@��+�@_�^�0��׃��ޜ醭��哢1�q'MJ+��:�=��I��s58>1%�V;��a�2�م�5��XK����>��w�8֊"D�Sikk�xKg�ПE���ů
����Iv�^�i���{Mǫ9��M_�_҈�4�j	�I|��Тb�F��n�>t�s�㎩LLR�Y�Bv� �E:=#�!���+rv]l����zp����V�O��8��$��)	v�B��36��$tVZb�駘e�nЪ����@o�X�k���Zw�gP�� [GT��!ɳ@j�d@s���{�6����]$`Y6j�WF5=��@����\�[d�hC�Y�"%��@������%�i�g
׹�Ei�����U~r="���:@���Os�;S�t���S�h��ڙ&�W��<V7�AfY���8Ɣ���w;o*� D=M�4L;)$��Y�M8�E��d[��CM#�9�<���x�tД{L����@�/f�~&��/�V��[���g��{u���2��4�N�� \?�f�Ϥ�J����K��n_2��)~��`:u�?2�SLAdӳ �!o� a򛠛���k���rs������#ja������ܪ
d�@��/׃;�:E�`#�D&R�C�bF��,��ԃ��>M7�|-*�~�Q|q�-���ؼ�C�~�5�ND�:����,�jJ��D�)��(?r��4J)������\q�"���Wvr���$���ds��Ԑg�?!J��3�]��8�[��:3�ۯ0��R���K=(9Pi@�O�$lY�J�m)8��ȅ��"%Q�]`�۽d�^(�;�`��17j��� I8V���P7����PfG˹�+nI���#�����6F$��P�x��3�:����u�`���/��I���5c=��_��FZ@����2�a�i�|�|���H9��73/M<��#��9nۥ�D"=$���H�|<��N��~���xy�E.���������珹$�Ի���{�x��Y�UcM��%뭲�{���Ͽ��x����dt-�v����Q}L��Ц��Qʨ�x>��HT.HK�̧�NJ���[��Z]������U� ���T_��)����3����8K3E%Rx~�^��.p-�%����[���Fy��6&�+P;"����p ��މ�c�	�HXVlu|��#T�{x�^/Y����68Y�[��nDg\���ЖH����#�34!�$ ����u����{������S�c>J��y +'V*T����7�Fy�� ��NՌ�*K���i#��p�ӈ�c'MAT�"��	S+�tZ��-���;w���:� ��+-��q��=����L�!c�7��Y��-"%�ݡ7m��4y�hw�qnP��J�!�2M�F㹘�aI�c܅5ϋ�б�Wͻ�V��|f��pP7���P�z�/����]'Tb��HF�ͯT����N�b�z`����� �I?�	N�`����u$f���J���o�����S퍶9��ap�&���+����6X���0C9(C9k� �qr�Z�5v�r�|d�]�/�QJ�x�a�����Ut? A����в�G��;c�7pĻ��p���T\%��Z�*�
���ꎎ+��1��,�F����Zd���)2UԴ�Y���Ebj'�i{q"�J90cǿ?��L��M;�)a��: �^j��n�5�ۓ4V[��_@�0?�� ���𚣠+kZW�-coi������]rT7�Ն����~����lA|k��;�W|ԭ=�Ꙧo�}�&O9�I�t�Kd���r֘7��;��c�e~#?2���`y�e����C����M�A�.AH�X�;���J�����H8�0 #��d͊R�Y�	����,I�O��=&Yr\;�p8�ϝ��-o=�Ƨ��ae9�O�a
8�;?Zb�w�p/m��U�ȳ�>X�Ss5�"�} �2�?�\�6��_����H��F}%] ���:�+2��`��ƕ�OU1��<h���p&���bl
�^10��;�k�C�� �1w�pf����E����nTP�i2d��>	��{���آ~YV���J3^h-������m[��g��a�U�r�����	'��bj�Ӑ��ZEK˼�=���8,���u�J�P.K/���mMq�hy�IR����'���w>��p�������oq���4^-�Z���uӈs��hy��TS���p��c:$���l�hXK�.���>���z}�fg��0N K�]�(�\}bQ�Yc`��b)�����a��q����!2Mm����	y&��FPPп=�8뱅�Tb̀�>t�`F��W@�mK�$������Yn����֏v9p��J�P� 2�k9��0���޶���t\]az/<.foS<ξ�TL��Gc�@�r]����ְKzo��\ߞMn��ف#u�r��E7l������Nل�lעߖ�*4O~>V0 `~!y���k)VS;�߷%nvA��я�U�W톍ށ(��W|�@��ߪ���q���c��=�ZӔ��<�b���P�Ya�+�_�d<�M(�ư[Z�U�*.�h+x� ���/4~�b5a�͔pl�@�˵ɽEh�'5�s$UĔY���/*�Ƹ%gn�w�&e@˙!�L2q���k	ݪ���S��~R3���lW.��𧮼b+'�c�.��/���^?��`*�����.�)'?m�rU�9�ٖ1[G�bĬ�?����}�(�#$/U��<�u���ʔ�tD��
m���u���L-� �v��{/B�1��^3$Qk�/���2D"p\V</-/�u=����O�y�A�ihz���rk��H�v�U�X8�8�.Pr�P�x�_k�)��Y@��b����=Z�Ĉ}�G
�KB�t�&��ч��7��Դ�ie�
�0�d?�����D����,
��5^��nw�~��EF�(*9d{i<\�P��v)�v+��Z��1�p6�w2�����D���wڋ.9�"��	��d���?V�ʒ�Í�͡H�X�"Ξt����ri��X��k�Q!��;��cG�Լ[_��5�f�a��4{6��*�����Id���/>�6�y��74	�������bi��h����O�`=m6���´�P�Ρ�����ݔ�_�~�2�F��F�E�um�	�mP~u��~y��-������ �?��^�1׵���b�������P[�J�gC�~�I%�7(^��������h꯸C��->�������m%Z�pu��o�*��<U۵�Uu.��'+XL�H'3Yk�_,f6�P��P]�L����W�^;Ծ7�[�L�$[���S��ȇA�B~L�㯋ɒ��yF���'�K�"<�;"ڕ����]p���V�ׯS�g�_;q��sa��H��l (2A7���T�i��.���4<3o�A�������W�t<Рcɏ�=�P���x��;�^�/�aZ%�X�7�S�S��q�BU�롇�X�Z���k����9��o�� E$���jW���h�#�k���uWK�_����*��:��6�wJ�")�9{5m��^[�)R���L�rgH�o��H;���b� ��5��h���eh��C�S����H H��!$1�]u�D�b8���дW�.�����G'a����I��Pzz~���Tޙ�)�?�,w2ڏ��k�-�je_/B��	QՅǇw�U���i��q!O��H%�[k�p��/ݐ���v��l��e`��߲*PH]�H[�Ӹ��:���3E�.��f�Y��� �^l���J��yS���Ѱ-��c�-��� ���ZN�U����Ԛ��n��������V���E�â!e�޳X�q ����g�����~D�~!� ���)<���L���)���×�,zq&op�	��1m��5�go�28K}�&�`Ʌ����$V��D/��%] ��'��a�3)*�uV�rt��/W����t֮~���г��%a.�o>g���]���r��.O�ƭ�a���'^�@�Iy��C�Ҷ�"m�i[FJS��)���Շ�t.�#߮f%�dNek���L��J�}%�c��<6�@~4�H/\�8����`C{�X�AK
U�z���2.��GQQ2�^�Ǜ�tq�>	pKC�zG& ��Y��a^I�3v�`:�d�爫��B��b���E'J�� ��q(��L������Vn+�8�۷,Y�Jk9c�����WFh7���y�D*�-��]?2�r���Rn��;��9!T�<s����EG�P5@D�ݸ�	�r?A����z��[��wo�<0�B���ډy�OXݢ8�2�	���8���Ø��������� ��Eo��k���<�]ں���M5�qz�JlRN�Oa>)�����˃"<Z�.H2�I�,��>΂�]�F�J�L��^��l�������xh%�i���T|�Κ��9�>N�ON"�D��͑;��eyDŁ���%|�zs�ċs9 &ä_�T�U��k����c�a�R�|�kڦwMU�u��̹��z�
��b-O�!X_a���R�uw2�նx��6�tnj¸7ۑa�v�j�h���D�{.�\�0�¨;5G�8���	T��>+~}�I~�F�/�Y���OHxw����ߴ�żbI�i���]�������7d��5��`;��KSr6�\t�F�@:�4�p�m]���@N;��v:,tiQ���"�eJ�;׿����̙�r,�]`�*$'�C�����|ܨ��]P9��w1����|G�GigY��9A
!�:fI��b&���難�\}� S#�bG�b�«�|"�_H���]��#}�82��>�A�O���bs2�� �Ue�PʿΘ��0!ILѭͩQ��o��G����X!��ڈ�OUB��%��LՂ��L��"B���*|iT͕��@�aW��"߯2B�?�t�%͗��zO|��";�*Ӷc�d�{M��՚c)��6����!g���#�-5��Z�%�4�'�:�L=����,�+oIj�l,�1 s�Y��d�@(��h��#ޜ0$�����kó��-�YM�j�ad>'����@pA����Oh[�J�{��|�E @1�H�עc�7áJ��AK�i�y�Jb���oh0�Ζ-�i���/K��]Lp&m�A��^�u�.Q�Q�k�4̜C�����7��x���m^PG� ~��
����c��� ��u�i����վv%_�[qL�
�̙z������$U��`>Y�.�Y��4El������% ��*��$�w^�;Nu�x��}��7����,sܛn[��C	��ef$��)ԘT���O+U\w4��3<�f���ʽ��X3�L���iJ�_#��+D��ђ��|#@�x%FH�g��P2[�(��N$H��֮?>�P��4
��Hq9��?:�oB�df8"oL�^�~�4J:�[7햢Z��N�F�, �a�t2[�z�i�Y�h�Vw�R�[@�*!�kC7~7>��W��FtG�m�7�f1��E[�y��#E�A��:�.�`����9�����{���p�H&w0� ?1n6���YN"�4�8;��9F�/�O1Q��e��u�bf�=����H.�Z�e�:�<u'�sH�͇C���k�.(<9�i�@-ƞjy�]aY�
��J�
�o����̮���oM�a��Q�`moH�<�K�A�fO�CݩE�M�E�����3@��q���$�&�1ʛc�?����h�9Y�J̨b��(���o��߇�'�2�D���5l���\�$~�ʊ���I|w�w��0M�1��hn��@_~A���A�A���k�w� �mHQ�A�0��\��FC���F�E��8����(}��Ө��ұ-:â��OX��n�_�E��&��������xUQ�F���=����¶��$ڄ1��;E}��*�OV�ȁ�x;��V͏x��׈��ӽk_<$�>�g�R����P��:����%A�~*����<	زu<TW��2;;��%P���D�wK�NOGw��ENƘg@�E'��:��1+�
Y)!��xi:P�	 ��&KY4>tA�#���ߛ��uJ�/�������3E%�ik��Hz-��FɎ	��U�pB�k��8;g��.��I�6pu#�������E2�t"� �n�u�V]��dƵ�?Ӂ�U�����Zw�:������\?�GՖQ;��A��a��M��A�Ne����V�]�n�7�>f@�Z��t=5�ጛjF���p� ����fv|^ˆ��������b>҆���?T��'U!@� 	{Yh�*��r��5�����56|E4ұ����m��;�8��h���)*��������y%�p��iS~)�bS	-W{��;ƿ���0Cȡ*T��n�Y)����ᕟK	[iz�����!U�~≭�J�z��֐j��P�gY�ů�d\['+���2��F���X1��;���f�}�tT��T�Ǝ�\���cv6�J��s�<]��v���J���x��L�*�M���7vN4�<��g��	<텛L$;�q����:*�q�C���c} �B�럡r�6"�H��A0`cM��ˏl�ޑ�����煒��OV�63��m�8y'��1C��)y�G
&պ��&_րx�J�"��^�Xhꯃ�5�T�"�����&�����$�ɲ��{�޼.���4)��;�*���E߿U�ì(z�r��-�|������uM���JD���e��b|��4	�~��IAL�N
ܕ���sb��P7�i�����㦣�J+�'�l�V���{��˺6^�m�r]��h�9;�&i�/�f����J~¸l��B���}o�Ӟ%'�?o��-Q�����B{�VFs��!s0��f$.5��7�y�N��sZ�0����f��8b�i��_��apH_�c��ک:sXE��1�tn?1̢7�4I�0_U��G�Lcx~���L������v��cc�+jrl��b�&������e�͘W߻Wx�?;��iȭCz�D�V���{N�(SQ�Z@k����.��&�ss�)���9��`�8�H���^1-� ��39h�.�{��q'(f���B�M3�ٮ�Y��~΢�t����0�Ǣ�_Z)����ڀ�Go6u��n#��H�����
��}�T�@��.@ղ��r�*�6�B�ĩ���E�V��߯��X"��L7��$b
��+��8qŶe�M��J�%�r(���W`�r�e}
E�J��e�l7�����.��s1jfuF̜>�@���������~�P&m����lb��2�	�kǪ��%�_�W����D��� \W�+�׈ug�Y�:�U��q̡b��ⶡi��L ��u����I�]�]{��A�����_`Ef!�Erd����g�we�8��l0�,�\F�.gʾ�E����q��,�M��?!����[���1~�Y4�c~Z��J�3z�f�����G����$������RcE�dO�7�2��W��&t��<�(�q���邴��{xe����� 1I�+@#�du�E�3�H��E�֯����k	jP���|��q��a~8B��`%{b�1�I���Y�-�v2$������ȚE�1��n�-����r��v	����h ��f��4^g}�L�r����wY��F�vO�X�+�w�f@�
��T&�⁳3.��c��S:�����D�-��Y9�.\�%%K��5'��}&�G�2
o���wK�r.c��Q`��U�{v��bk#A�=�uRL�������jf�q7=�0�������S��f+B�;.�������+�ws u�>)���H��)M<���8�}{u���jo$�A(���$�r�����A?xgZ����Ղ��(�5��6��@�7�~QF1X�0,�;v1��"�h�Y�����@��3�������ﮇ�ЏzH3O�����Ĝ��E�TTǙcΪ������m�n�2J�!�3	�73x�5\4o�K���/,de��X���0ox_�?�hdXӭq;;���o��%����'��	:u��QO�c��#�[�Ě���O1�ߊO�D�{b?.��K���4� ��N0��	���l.Y�����w�(���z<�;�P�{c���*�԰��T�|d켇 A���E��Z~�X��&��0*!j�%�x,*,U���k�:�e�Q�SUڒ�M۴�]�(�{v2nY�d0��s��qm6@�*��&��ʬ�F�;�~Ap�
�g�w�2��Qko�?䙠��NXXU��!�R�
��������ȼ�jC&���#F��F�4��V�i,L�9=q%���ق] n����W��l���3sa7!khd�=���svFe�L�m~�2aaJ���x˛�R=��蛽�#Yi\ۀ�4����X�p�����V�#�����A��aL ��}d[{���LO#t^]Q�A��|xV?��LZ$���ΤS]����]�ի�'m�w/�k6�?.�g xq�$�#� <�~������c�Ǒ������l�>�l�G)Q�7Ӱ���]�TI��SK��u5{˧"nL����{/d�҉�#��2v���j��Ę������
�q��/�d�1�<�����A<ʖ�#rFO�?���x�Z��zh��g�UC�S�Ng$�����.m z�gd��s���h����=��[A�[ӂ�T��h$�����M�4�W7x��\��J_�´���͂Q�����lD��u�nk���h��=����Ԕkg����������t���+�9��	�l�xJן�U>|�L}���>o�e� �p����C��$$�W���j&�����͸{��Ɂ��*��u��2ps;ybW[��NT�7z���}���	��kbo���[�%[�|�Zz� _Gr��}-:�&�����E����A	%���:h'� ��[|Ρ3� ���*)U/h�����.�Ö&���6��56�8F��4bzA�Y
�:b&PY�[ź�_�gS/�c�q߻=�To'U1r���.~�+N�Q�L	-T�(YnP2�&�y]��kg��i
Z�2~���7M	�H�Jg?�%n�f�u�e@� ����:���4�;�wW�fLA�ηO��n��n�=�� ��qq�����ױSr�۰K����g;�\#���<(\Kl&�C���_�����F���L��^�}r�@{���g�VbS�*R�r��:��r�.=��|��=��gX�q�keM�����2`?{�
r��kz=��*���X���K���Ҏ���2<�Τ��d��UG�]1K�sJ�{w�����%=�5��҉j��:�c�pX�z<�����q��2U(�����W�
)�֣�a�L�q:p�b��m�J5<�?�ֵ�O�'�P��J<�Yh���GA�-L��z�\��
c
T��+�)ŀ�Bo,�d��(V��;�]���8-C�B̦��������y�p�ʳ�N���9�N�E��6N�n�ef�|�}n�V������sX���Z���$�nd�Ԓtlr�]n�{��)�7���#��+�����@�x! \���Rn%�[L���Ϟ%,?ZR���ӻww	,��J��OEzT4q-g�(q��1�uT�7 2X��I�!��3s���U�(���F��9�h���}��S�rެ} <��`��Ǉe��lit6;�S�'��V{Nビ��FQ6�G�����o����c�>�N*����o:�x����`AB<�Cojq�#��W���sA�V�
�j��h�$����w֞3n�k��<�Q�RC��f�(`�
}R�5X*#:B��ś�d���f�B:!��i������1�k<��L�qaZ�v�d}0L�$���Jœ���:����W@Q r^�O���}j=�d@Z.J�,�c��De$M������Z&IR^ ���
��������6 �1wS�t��:6o�5�%	���������=ȿ�Ohg7u��Ȼ#���x��ޙ�7m ��Qa����_l��\�2���$+';�T����ԫ�s��8���5�F��n��%S��������{{� �_���}�Qf},�5T����0�q�'[#�SuE�ø����%Q-k�Y���v%��N���;����&�褔���C{��49C=��׏���1@E1�ŧbj+�x�?��I���1�L�4���c�Djc� h=T��$P���ئ^��ϛ�7���5X�x!�T�w���j����� ci��ci$�؁)�&�=��f���xf��g�����^�70R�J@Kp�����JJ�R��N��6�Ske/���)��̠P�fK4�,�/����gw�o�F�*�צ�c�#�A�!�K� S�r�A"��I��4���u�;�V�!��m�v��]n����|��x|IV�^B!�C�(�%�%ݚY2�U�0F=��$b�3�\�* �A�ށv��.h��cB�o=��8�j�={�~�������u$!��0��j>�ۮ�T��N�8������,@i��3����95�G���}���}���I����m���#[����e[�$g�x�T$nuL�8Z{�������%,jl9��;�:�vڄ�D�s\����kL�[�1���-��� 5�O߽�>Xr���w``�r`ʰ��X��8څh@7�rRA�~[�H�&�y+��oS��{��!L5��|Q�Щg��l�C�O���������JǦ*YRڋ�atDɣ�nz���xR�ƕ�d]^<��cJn@��|��y�Q��ί��毞����=��O�ـ��y0���\����� �dQ�r}��GN#���2"eN�PAt�K}W�Ѫ�j�o��fNH};�p�h�
{L>}I;ѩ�.��T���k)�b�'�vD�,2�����Qc+���4:B�>�����ͱaf*e�v�.������@��E�z�]n� w0�Y����<��4���s:��Hϻ��e��n��9*1�?�.X��ſ�x�`�zAެ/"�j����8���h@+y�҅�{��9�X���mDT��f+v�W����1��
N`��J��K��r��z��F�wl��������d=Uu���q�S��a�A[�㞦�g�tgT�6e@S���Az�1���-L��͂j�e��ި�K�
�G�pu�`t��٫q�P�$�s�.��"�Ȣ�~
xl)�	W��7��@ʚ!<�I�����结nMQ�0�VN�\���e��X.#����P#2Bn���3����T�~��a�#s��0��	�i�Gg;h@�ˠ���I<}]8c1d��Dj����\�yb�AE���p��ϊC�w�n�y':uѼ�H�d��g���\*� =�8�`T1`���~Q$>�,"�l{���{l�[�T����>1J�LB�Kr�����bF�4�f�)=�z,ӆ\u�14^{\����Q�&^Pt"؟6���㟾{"\I��U�YII���=�����$��Tf�3�+	�tnTZ�_p���r<�"Vh`�?Nk�����z2:6JP���݆PO^Y.��c^�#�wJ����n�3��Ĵ����t�`� z��Eu�ۍ�0�S��ݱ
����;L����}NݰȮ�>y����-7����!֎�����gN�]'�u�',K�Zd����)��\��F�O��ݣ�N�������ۨSΩw�����=���RlY�%�aLѕI4��Ua����8��D�F�)"��9��ş��w�q�FLo���Mrqb�����\T�����
��ؐ$�@�cv���{�6VsT�XB�<��<7��R ���쎇��e�Y*�SZ�J���H��:��5�xq޲C8�3�˶��̺R]d��A�ì?���dIR[�!w2r�Ֆ:*�hp����� �Hht�����_;/�'0�l^�������@������UUe�����v�+="�f�}���Y�JLAQc�˨���v�ӊ?�� ��v���~wLi}Ӓ U���0u6B�����Ӡy��XGΒs;}8��8)4%-��D&�*�i�U^6�Su1�᳢Z�lF�E^����h$FD}�K�6e���\����P��/�]�v�"3jGn��D�O6��}Ύ��n�(�Y{:���=]�0o����/�e4�kO�fM�	�<��iĠ����N{8�6���A�_��`L�C0���D�"��zB�5���3)����6�J�c��h^H�r�J��W�P�\�>�;������b�XW�a�!]���'yp���818����D��`�nm*AԈ�H%B[���*zC ł�"g<+k�qA*�����C�����؋��PPD>����ac��5���:(��qn���o �QF.�Z&�j�:.8���T�p���KEݲP�T���9�Q��J�%�0����]���ꁯ�e���'�<1=��o��
�<h��ވ���\�P[;��ra��J�7�w���7�������T� �dj0�b_Dlt+.KK�Rjٮ�#��m@�T��?�]-12�`�w&]8<F����'=$�<�_D��Tнt�b�Њ��T���/�C��ݱ��X_���3"��5hø�jT�)�)�qv��zW�o�]yJ�d��L�E����	3�u�XiG�������o������`$E�G0���\BW�C��E�mN#��]��{o;K�B���ݭ�Rɛ�dH8<�1�(�ݬ���+��q�Ee`1���
B�� ��ߍf�i%^� E43����z[%�
4+����\U�&*P�6Z�R6�r�X#oBe��_@*CsL��f/�.�LAS��E��i�u�$$�gYMt~�|$O�@��h��=�
�7�TS7��b��{������ݚ"��)��Il�( HЅ��a�Y��P,D��<f�$b��kx�]�ا�>i7������0�p�6l�&��m��d5ũ�[�pG�|�ٹg�\��m��FE12DُQ�8��De��z[�/Yo�Zfe�ͤTxf�f*U�I��3�a�_޷�̫K�"�yV��?��jQ��8ڈ��[Wʷ��B�)�e�k<,������K�W)�l�;y2� ��l��W��!�4%�9~믲m����'Ǘ{/Y���H�gT��.��o�c�h�-(���O)Z�G���[�_��d��w�>�1�<�vf� V	��+p�2�'_��#�Q����Mg4ţ���<s%��Y��3����E��~�ǐ����s�J��������㳤����RR~�%�Ht3�ҡ���!�O�("����tDx #&sz�h�|��<3B�3�`���hF�Ě~�jln�V�t_���}�$�Ĝ����ʂ,;ڻ|��!6�܇���MX-��?]�f+�$G��n=���SZ^l��D����z�YS��@P ~L�@[-�)������r��@D���J3�^{���J1��!k�w;ٰ?G�`��Ҁ�K�e�z ��1[�lP߾*f�U�H�c��(йؽ/�V�Vd�33�\*�m^�0�)����� Ww�i~.�����V��ܱu~�pA�)�\� M����PU)M�X/��Sq�Σ '�@���j�s���lu&i�~Q�A7O�[U���Ӈn�Н��L�S��J�!_�՝�˚?�Q�0�,`�����Fq��a?���`��'�H�v[Ռ,�����.����O�`JN˽~;֛����E>&$�H:�L!/Ղ�!���*m~vU��x(0F%"�+��ょ ����YVd�@����&�����p��4�R+�}�YU?e:����ixX�q����p�X^f��Y�A��m�'^��+N�p�K�@<����S����3[_ۗf(<�lo�I���F�P�gF�����	��я����+\S�U��EǾ�{É*�՘[��Ds,���8|[w���s��Lva�}����%1��3���a�I3��ﶼ��L�/�N�7���"�P��5������Q��|��I�w�:B��y��Q~q�1��m)�Y'�D�浠t�T�Ε��@�T!y��4>[b��r�r�0��X�;*CI���x
�L�����J�>b'44UW$�f�+i\)���	4��8Ǳ�E�+I�z���6���j��ϸ�#��G~%Zјʌ|�����`mn������)���W���!ц�Y�zC��V\?r4�y!+o����QF��X֮5F-�Iз�]ɓ���ʇD���P��;%�2�V,���ñ��0�w�SY;z�l�r�"h����d���05sc�{0�A�� -�i�Q�s����i�;�qȾ{i��14�-��G�X󚀠�J�Y�v�N<�E��D�9�Xy^��y�F�́�R-eC$Fk=��0�E����U����� 1K�DcM'$:��uk��i� �)+���|9��k^�(�U���!P¯�	�Y�8Hd�f:�O��� �J�E9S�f���?�Rfy�+6�wH���5�w,��S�g�ιѝG�!kv*�q����!��	��J����Y�,��L�`1%�#7�-��_���p�����+�a	��TP�r�v���H��0�.߆v� �H1����|�z&F��3�����8���x��ʶ%0�`b��.
qn��g;0����53����f��U�ܺMh~�E����^	Y�QC��!h��U�>��q�z-��	uA�%NI�t�v���	1�=4:�����*{�T�����)�T8]�%��(�rR&�@Z����h��-:}�BVq%��믯s�5�dg�F�'��Hk�o-���55G�s��Oy������_�p��e�l�L[(�E�[�F�h;T�B�c���+�i�c�w��2�K��9/k����օKVӪ�=1Zv,lʆf���W�5�vF�@��S��(s�4d���66�ob��	@~Ľ�t i@����i0�|rM4�T��Sr�	��T��9���M=�g���,�QmӾ�V����>��+ܿ(kl�L���{V�68��Wv%4�IJ@��^��-	��?*-����ty`� �q�`�Y��o��W��̲�|��+M"7B /;�mt�r|t�0�+�Ec�Y�Ҽ�?����[<�~�!�r�M���w��bhnn*��_&My����N*E���n�_�w@-u
\�4J(��d���(�������=�e>�}�,K&�,/�R�.��_ H������C&��Q���Y�87q+#Mυ#�.�m��K�6�����A"�i�u�Z�ͲUG��ȧ&@��D1�n�e���hѱjl�x��En����T�����^����]���b�ap?7�KQ�7Y�ro�͏hVoKK^o����{���<��4Ä^�|g���y�������hU���4�BOba�H�آc�$�@,�p�� �<�78G�)�����E�M9e���R85�!D�4"���J�j������;�{��i�^�$a����y$�5T�kZQ\o*����$V�3di��q��Yh��]`vaZnZ!  �n��z�z�(��̓H��;c LU9�n�,��6gĨ=�ñΖ�\i���/�M�t�J��X�Os(�u�b�5��aZ%E�8Ѳ�|�.��8�x2_��h(���Xݡ�q�!�R�BT�Z�R��t̺X~{l1$�����,I�-HB"D�$��uK�Zۋ�w��{/�K]���?���qp2��ڨ�ξ��C����ЏN!�o`��Ww�67Ha�r������[���oh�� x0���5VK�/��,�*2�l�7L��Ww�-.��Y���JH�;\��zo0T�'��\4����ݚ�=D��*��>�di�G��0�s(��?� � �Z八T!	^�`�JoP�	�N۠ \��TJ�-S�`�am0��B�$īƝɨ��y�>��n���qG�VP����9��'�#Ǐ5�O;�5��v���W�*=�%�a#��D��OV'$9��7<=�šT;T�At8�Ō�bX̀�]`U8�d�g7�m���fc�QM����.J�R�&f�8���y�n��Q�H��e�(k��'�[�H8;�y?L�N��d��1� -��k�ԑ7�F��V�(�h�9/S/�芚rgԷB�%"Ed �r���u�Y���LBz���1(�P�k~�)3�a<)�P��Yң8�e\C��(�T^�o1R��!�!�X)tt��pP�IX#�$��_��ё@��U���\��F�bD��;$�k���`*��#ۅ_̒���9�p4�T@ͬ�Q#06SC��m���Eo�F��K7Nۀ��M��VRi��d� �R�p�@�BE��хp�?�[;~�&܂kd�pX"�7`*����ikEzh�G͎���D��P��,vR�o��A�F=��n�Ր�b#詄�4��E	�t�6{Z�9���n�RT��c����Ё9�o�NC��S���W���* 7~�x��px��ŗwۃST�|`����rqs�W7Q�'��t@$΂����~@is���\����L��%8&Ơ�]b�ǅ��LB`d뀩Ns��+�~���Ҵ[e���l�[O�uciÄ�]��ĳ+G�����5�>i|$�ȉ��79��B!�&-n׮�K��!��,��f�����P(1��@�nb��L��:?��m�/��� Nwz	���|���<1�r��$��o��A㕕d}g����_����A���ɠp��@�A���błΠs�+웁a0��0�CK�����&1s�̹gϓ1��N��šAo0O��MZ�!̈������ ���bv����an�g��W|�}�w�J�������-G���7����Ȝ�Ѹ ':;�/_��̝S=HG��ֻ��W�i;@�='��L����3�wķU��I�2�\O�j�rV4佗���Bc�G��bl,z�1��Ǡđ��^\���#�^�Z����Jz����Z9Ĉ&� kd�4D6�돠�N��#L$Z���jLZ��&Ì��+oQ JG��"�	q��^i>#%S`La�f9�ǟ&��蠔Jd�B��h���3"�*:/��j��,�!�֙��f����Z�_uB��E��lo' ����70Hg;�yb��,sX
#��,�)�3��הG�w���v�z�6���	����1d}��=�������YY�["���Ū?�u�n3�Q&�� �nh=1^���c�޵\⃉+��JX\��Q�_�X�U���@	�k��V�t���y�_j7�Y��9��lWn���ql;E�0w�88�o�b�U�\]�k��v�;2�TeA+~��Њ�?	��n�p*��ގ��)�
�Y;I�L���ٞ�
.�8��8�j�I���r ��������%��H��S���n�����ݬ��Dz���8(@��qcp/MM�u�� ]��D�䞼�lb�r|�k!������,����lzwn�'q'�Ɗ��5���7��1�n�z�P���v2U�@��I����m�6���e��u��M��$=� 5Jl{Wz�PZ#���}� �ǃ�a��=hy<�� :��`��~��^�Ѕد��l�M�2��|�'պϖ�xT�f���+W���* ���DY >s�4����b~�'��f�Qb=�Uv��J����	}{&h*)ќi9��kI���ڥ���-Ŕ9�sֈ�LI�M�i�C���m!K@&iB�5� #k���\��{����/�NIY�=����G13u
�Rǀ��\�ࠍ���P4's�]�jv'�A��LB��(�PD�*�'��-V�!!�S��;��B��F@B}��.�}EJV���By|����9��p`�=���ݤŁ���̾�k��\UM��Lbv��񄜣�X�)���u1=���ªZ���y7Re�͓�86�Sbx�J\/�U�Ҋ���X�d���s��D���%�z���JtD��DR�W��w�p��O��]��m�a���i~�, ��f!{ϫ5p���&���8��09j��!N٧��e�o�6�z|�xכUg鑮����1a��3a��|kQ����9@�?�� �z`{�8w�e�Mv���}��}��miQE�y�ѿ�*	���i��� ��2ӅM����2��{%Ea m��4�,݆��^g���K��$�T�&����U��^�Piz�즩\�y:���^ZM"�M~���$}�l��\���\ձ�Z���K��L"���%� �g�,;�w����WO�s��$�<��X��s�E��ԖG,����u���_��b�����L��jhگ(Q��oʈ#�G�o9|vf�O���!�l��>xM52 w�ᛒ�;̭L��]��AJ�th���� B�7��h��J_�;�#�>e��H��[g��斳�[2[�C�y�My�"d���PT��X#�v�c�}��y���lFV���_tm�St;O��W�����w\��
�) �b���k���ⵈ���+��(uc5�Vrf�6�4mü�v!$�
�r |���JKM�*���q��Q�f!<�,�Ϊ����'WΎP�}'����	H��&�p����Ζ��E �E�0��r�?FUF�f��f�6җѦ;#A�N�|N����i�m�fwpR�0#JL��'�!��N{�	�(�.i��'R�7�O\��Uo��o���{ o� ��9��oəm�P[�S@�I&o� �aH�l�����[ܽ56�9АO�^�ځ����/A�������~����(��x?���_e��ӥ�)I�>^Ѓ� � ڥ(��<L���J�v�cn��D�2�p�I�Fa�lٻۄ�Y��7��|���y�$�-���Zv&�F�9+%���O'�9}M|-�x	,��[x�K���2H��꿋n��5�c���T�M��Ǭ�P�dZ�G��#�j�ta ���2��|�R��
뮔8���ⶄ3ʔ�0t��۽��=�>b�}No"��o0	�9O�ş�87����܋9��e@������;���]���;v��MG2���/��q8�u}��+��qC�ru�J<
�ă�t�ƺ�=�I�۸\�QP�L��8>�Hk�T>��1�uF�|�S~�څ�8��m֣X-�v����
C#�n�z�ag:�ƖZk�+ߵ!e)S����6ɛ�n�I{x���q��n�%4㗸q]"��TR��\I���xF��w���3h���JhN��<N~,B�4��%�����$5�g�)��VY��Q�ڲq�4|����YYv�TUS\˶+]p�He��[��s����)8��:�VS���!#U�P}Dw5=s��H�xC�,�\��;�oq����!!l�gm)�Y ����}+~��{������u�~��N�Y�c���Mfܱٽ����#8�w��TH��o�C�'-�x�wD�xj4�<�՛by�F3��+���.���|�O����!ǐ}#9}TQ[�-����Ҹ��}� �q��h�44���Vxʸ�#��![�j��m@��I3�;6�dk�("/m���̕a~�,����pU7���V7���eT��	��=�MB�����Wl�FY�1=񞒞�SQQ��6ѣ��X��}�tT��}��䬌��q�T
`����A�:�&ȩg��H�X�k
q�=��g��f��eNFk$�9H��n1)��G	V6p����G4��|��wю��Y��@2���l���o	XB�˙m�߮�ȴ�OY!��K(zl����G�H� 	��MuI7D�ɱ^Y4$�od.�L�,Q���?w�0��ID\�Z��	��9�Z��!�/Y�΅Ƈ��m^a�S.�}I��©�X�Z�����H߁*f<���l%����8?.o�x)��4��������w��?�D7�9�w���.�"uȦI{���Df�ib��J�$������{-�����3~��+�^� f���>V��x�rQ����U'�D���Q��r~8=�BdB����a��V�\��5�_��u���(���S���d���b���.�0O3VU�����|N���{��ug똩f�t���k�Z�͉�C3?��wQ
�-�<���1D�D�0J-��H�RG?�uH�\<OmWf��+����ݓ>�Sui�bn�`���tu+Z����+Ќ ���0�HH�	6��Q�pD�r��I9���ٰ���*�
����� ��?��N� �&��LZ>MV�ӽ:-F�޺��.��@w�5nJR!�rJ��S�-�ME�Gc��+_�j{ALB_����d����/���U{�2��&"�̹����&���j,v�~=�cd`�������0lC�ѽ	W�i'KG��ozP})�`Y�D�̕�{&�O��mD�w�)�}����s���[F��ECas��o�]��ᶳr �'� ٙ�\�eӼB;��n7O;�h��E�̲�Gq[�4�9�ߨK]��#��_��\�v�ʴ�gy�	�tʮ��8>���8Uw��T൫�{��I)fkǌ�M۟��*�{�h�%�����gN4�o���R�Qg�F|��KJ��yÐ�`�*�M�� �̿��
)�2N���;��J}�Xu��(En�U���V �+Q�L�iygٓf�7�79�"�m��׾T���M9��gxK�d.=��!1ޓ�*IkBl@�%;={�[���Mܼg�����k����s�e%vQ}(��=���4�& ��۸A�Q��cϺ!_��K����l�	�NVK�]Ρ�ѕ���A��'��1�'�Q^�uF1��#T�}%�;�^c�2O����9���hg!2|���>�I����#�w	��������D�o�P�,��xL�9������V���x�Ϝ.?���a&�o�g��0�����M	�ɇPw51 ��;t�����r�e�2����;6�`U[�O���g<���-u2��U�MjH�x�z�]��������EL���_5����y�+�5�hK������Q����wI༩u�=QT�雧��!� �z����m��i�}��Y,�I��nc�yW��m���G;a�@�v[�V��b�G�U�l�㩁�Խ����I���z�Xto��*M9��b1��b=�-�p�J�t�d���3ԑ���!��Z
�!�h�G`���҆���Ph� ��H�jrmْ���<��/7�ȄO��HX,܂Ԗ��
�-A&8�#<[,�L��1 �I,�~%���|�D�d�r���Y�Q�9����0�/��/�e�'n/3�u�ODR�3|��ݯ5��"X�1�#��W������t`&��{SF�t��J���^���+������Jd��'��o��`�{r�e�=bW�Z5�D�(-�#�/��_�ϭ��T�����g��WQ�>�P�H�%��%���z�0{I�5�P6��a[��S�
M�~	��w[�6	�.��[[��,?��;
7D���;~���BvC� �hq�Ι��I.�P�;��P�7�U�w�>�kR��5�$Si���V�;��$�J�lQL�ǤF�SE��i�)��=�֏k��`�;8�;qt�-r٥�s�v�S-���YS4u8M�Ѕ�4�"��A��@,Ɠm/ ��az¬M�̰���K1	ZA)���p������MnV@�v��`��ƑJ�I����) D��w���	wd2���*&=ݧ���P0t *��`��1���xT"���Q�q�E �Ѹ�/����:h�������Q��q�A������A��B�?���)��\���Pʲ&�i0���D���5I	�?��s��"�A�O����u��J�T�HP	V����8//V��ߺs��N��}��a;���|���`���i6�^J&q-�eC�I;	TT7I&)۫$� 
=B�L�u���/p��!)�ɕK_��6�;�������5O���K�A�I�1�&�1,8ß�=�m�{!����Je�у��j��8��r��m|�΂��Z��	�>�:���/e��Z`�+�Ʃ�ɚsC�)�`/@����M��~�l�w��+�+[N�47�;q���ҷǢ4x.��H=ґ�
8�2���dc�`s'U5j$����m�<s����0�Id8yl���KLF��A��g�ނ���������~�3�oy��
԰�/I��R��B��L?.k*���9��k#L��_^�p�A�Z�'�(�����b����#@����R4��`�p�\]��򎿟�
�"%��@$En�^ �!y�8_t�W��?9�"�/��ݛ����%%�����pUƑ5�4ۘ{\J�I� �Ⱦ�ۏW�v vQS�"�U����������������oz�cEjB=�b~�=cDoVI�fT�NH�������k:]N��^E2�c4б7ұ5�Ӹ0��%��4�r�kr;p�밧�Òwxw[2E�ߚ~������3��< @�
X���	�pDV��U�ר��[���B�q4,�KUm*�̥f!)/�ՠr��E*�%�Wg��pCg���yd>r�Ȑ�}���;:�DIMp�9n��x�$�&��(�/J#K��4��E d�ߍڿ�ԓP;Q�ԤXQ��L��u�]��T9ʾ��k�"En=�O0y������gӲ�m�c+�Ɋz	�$[j�K���޿���ˌ���D���AK����,�G���WY�f8a�J".$o;�i�k�rL��n\H61i��Zq-�|a���a��u�c�^�pd�
��t��/����SIn�N�v=��dw��&5kD$���OI�Z�О��<��c2����_z���Fi �&�Y[/"j�Uu�h�17�כ��̪z#�.����.v���É�kd�n���C��v�m�[=�+�l�����u%�`���d[�Q#��.4�r�� I��	$Y�Zdr�T�0;�<|�o�S��D �s���z^fA]������X��=n�㫗({����W�:�~V�UӶ�N\���T��>A0�Ec�c#�����]��)����k���h"�ϲ���bu}r#&���-	-�����h���w�5	���$��G��l�dN�����t�O/1��#5~Uz9����َ4�T��<���kЗ��Uh"�\6X��~���!<[o��{f=F^�����)0U��QJs��"������dx+.��l�3FIs�-�F?r����ǊU�s�GxZ倽W9�ص{U���b�Zɲ60��tѹc�	?�x��W�f5ٝ3Ӎ����-��C�)qO���qd�� �x#d��s>��h���[��"t(��VQ�c�F奟�$���%0�T��X�/�ƺ��Ro~�j�@&V���(��,`�pf��%B%9�K.3��/ ��`t�&Ti��sR�p��)[�&M�.C����۠$z	���֎c;��穗�|���_c�=V�W��'��r%������3��8�:U��?j���+��,=����Pe����d�ˊ_��H6S�{�RB���G��m��y���ZR�}-Y�Ep��{Gc�����3���Ӄ�C��t�=�������(Xd�l��L5ɈBaʥ�3=ӐY�K9a�c�[H�����k�mBԆ�X���0�4ލ����qL˜AN�����R�gV���wL%�Z�l�ކ�3��9��0�����@�/~4m�L�h�ʕ��u `qL�����{�6�����O��C�b�B�<؊!��2;�$�C*T>)
$(�'�����D�ʕ	�{a�ॱe�V���W]<�:�Θͼ]�h�@&7����C��Yje,���Pi�e��`��7�]eU�A��K�,m���0����+�r#g��ۈ��Rk ��:��o՜�-֧����5���Q��b\	Cr4a��Ξ}��&P1�9B�� ��?c-M�75p
��b��6q�m���,���;���+�}��˞��7��+@�r9 �+&�1LzK<�(��!���*2o�p�!m8��)�O�4�^\���'jQN��$�G|?�ío6���ՈX�@�Ϻ��m���j)�����o7%.��j�bP�[���FO�"y���W~&z(�:��S|h�O�*X�"H�pm���L��@�r���#��*��gx�5o�������Q��� �D�>�����n �}�?P��������=3x�2,[si5{ �ʟ����8���G�"ⵇ�q����-xeZ����f�1NM�Li��A������r��7�at�e�Y��7�>�$�j��`d�Y���$B�Uz� `~G�r���(�
�~�n�uT��Ee���Tf/�=�{)�f��(A޲J���U���y��37P��B�1���� ���D;��iEN9P%K�H����I)vk�+0�˃�W��t��u�-c�6&d,�4��.��S}�bᩒ?$��+'ً���Za舥����3��G��gZ�Z��q��m��������5c�s�s�O;��Y��9�O��:v����$$�|v�	��^G���^H����Tf���ַy������iA16�JV�L�G��>7����"�#����Cm��4�� R5�e.�!��	������� *p4���(F�����^�p1�5�ur�h�L��C�@�Ij���cdV�sv۔�F�;�re[[Q@Z;e+�l�'K��l�lF������_s�y�ۢ��ϱ��Z�B���>���A�6�����@����qN�i�h������QWO�:��3�U�M�X[�̡ve����>�������ѫl�
�m�����Ÿ�6"��-�F�b��SEʌ���}L�'r�`L��F��H�r��]d����E��R��[ώ��H;�{��'S�'�H�W��W�����~܄���f�=���an�$<�����J8�~³��]6��6~i��|�?��F��,hH��P�V$�'��A{]�����y��l���9G�i���r�Л�L��ωEQ�X~��w8{S��0Y���(���,��~|��Ӈ8n�P8�(�S�������1�~�$�8��t�&]�y�'�x����O_�O�CD{<�_��:�0M%EG�Z50�~#�9wm7��&=�>�YYk� ˬ=-_9�%��x!u���Ͻj�v��6gJ�#ӗ��<w�p�����A1�r z����3��f�֙��w⬢���>�,��]l��x��.Œ�k9y <������^.8����JY��'��-U>��F�A���
���_����v64�zj���l)'�B�f�=#�y�]62MȞ���-ˇ-@��ol�L8��Ds�mJ��7������$���pMBb������I���ɤy$9���yz�ަEj%w��y�1�c|���AU��6]�]������k`�F0#I/\I_�E��=��͏yrd k�����d.��R��-��Z�;I��~q��2ǝ?�
r՜�#�E���}7�
���M��c���)6`]�_�O���U�u9��|��KP`����ԛXXa_�<�����uy�Jz�w��XT�똒���+���mݠ��Io�����;���4 L����v��j4��E��	!�ӯy��{/~�s�L5�q��'�q�Ė,S'�"U]���CRp�4��e���nz������Q��^��갆t��|�-{jT���W���@�{��<q��=p�w���!n����8!�d	���r_DB�����訛	�O�kmz���u�G����s�}���u:|�-E��OJ�
c}3K`X;���GE�mv�2�F[��r��B�B�[��&�$��ّ��<u��Xw5G����|$�#a��c��Nt�Ņ2E�p���R��"��YS�f��BEO CZ�q���£��e� ��0�#�����2���y�뎨#�R�&J��͐��몳��IGx#�p�<�L�4K��y����H�6�2�h�H�{��3r�@6W���;�����d�2�/]���!�W�Q�z!��`���k��3�o����P��p�\�{F5�Qeu��W�/7d}|�$��`�~*wk��fTKN�:)Sj[�؇�	"#ѿ���6���ޏ� 3��"*zf�h:ʢ�DZ)N�sA�Yi�ȼ��4��j0��������A�FX>5�b�����.d ��Ӳo"�O����������3��=FX$ ��#����@���o�����wv#Ҳ�s:�&e�1��07�R� �
aj�y��Lȗ,+z����n�A-���ߔ�Q
z�-����i�i\b���k�����Ͽ;I�s��uRz�EP�I��yTI�;k�{�㐈
`Ȳ~R�YnP[|�����U��~�7�Ć���"6�̀�h�n�í��b���˿�)�z���z=�p�J�f%�p�����5����=��3�y�OO!��:��HyI2� m�'�G�r$3!&�7K��`�_����{5܅�q�)�9�n�Ta*U�򬭒Tf�t���ط�(���!ƀ�B���@��cBT���9Y_^u��q�R����4���d�*2�och�^��2��A	���w��쨑��b�^]��ﴏ}]�f�,��:�M�*�7g?��>�DF`���Ӥ� u���U������OP�[��տ������Yŀ���=�3Jf��8�:n+�<��K�g:!c���z7�����-��0L�.�h�4�"c���k{�S̥?�rD�R��\�'K�����O�xS��-T�A����P�Nk �q�Im�D�1]�~�'���jf<���|���9o��h����7��{�cX:=I�b�-C��7�7���^dK:�0�7
����֯�o �^C��`n̛2 w�h�A�I(Yۖ{&�U���C݁������al1�$,�Ua��kM/�cu���g�z���	<���ӑPL����
:I��:OcY�?�
�S�-{z
|渱E�"�d
&d��q)�Q���6�~��ne�����{q���k��q��Ԧ�f��m2�u⎳v�_�lr��*$u,��s)Y3o�������QK8��k�Y�t�F�;X����O	L��v@�s$h���wR+���9���b�4ec������ z�	~��M��͋Ϧ���z�X��-�����L��nk-1*`�_�%�c4�%)�`�;��s������dY��p��=�~X��ˎ
��-�a�m�ƽ-u,5<���y�{�$;���~�Wq�8�H����ǃ��)�LQ��_����-��@�o�
��N|�@��?�E��(ߎ��d
Q`��CH�b����\�z���s8�����>�D�V�ϗ�fTL��M�OITr�vG��*h���6K���>IV�y�]^4NX��z�Ė���Di� -Yd��D����PDzu���u��<����7WH�+R�ş� ��	Q�%�9�|�Č!��+{N1M�L�fM�!u/^���Y�cU���do�f`cKaM�(�u�T-��g/!�L`�`9�Î ,�,S�W3�[�"Ƞ�uV<�!�Xz2�?���<n+�E,��-���v��# �N�V��%1�\�4����ֳ�W�|k��E{��v��+(��$�b�5M�3��jm�l�R=�-��xh�W��g��f�!�ym�E�{PHTE�B�C�����~�WITI#$�o`�A�\��i����~����v�
�Xf�;�5} n&S͊T6;>���T��\��k`x(Յ�	�,y��Ƃj�ǯ��(~y���)�X�=}��+/�u��y�xw#��vw��y`X\#<�/m��95�9��IJ0(�����G;̢�ܾ��i�eC�7�9H�($��oFa����˰`���F��"�c9�<�)��;kvv�'V�]��8'��r����Ů���;�#8�Vs�ݡg�kߎȉ�Y�<h�%ː�z-�@s���J.�6����S�H|�ƾ��Vӣq1�)e-y֌⩴�l��y�.�h��m�����Z`�V��c��jk��V*�6�[�����8�j�D����L^4���_˺����������o���� d*��`A��2+���-4Ή���\x��p���g�ډ�
���>y0O5�[���/��#O�Nm���8h"t�4��09y�/m��Ɛ�0� ?q�LM/��kfC�Y/����N�C��D��:	��(P������m�"H��Um���/;�\_j�"Mm#$	}s�v��{�Z��r�;��f�ϰ ׅW��黀�u���۞,��� JS��;K?��S�}��> ����u��i5V!��-��T�Σ�6:��E����`1�3��b��KsK���s՜�㞈���$�u��J.�D����#Ӎm�0k������94bu2Zk\%����ȼD��Ʉ�R(�����1Ũ;l��8�+�E���ʕ.N~��:�X4'��$�#�.���?z�(X�כ�b�@m��/�f��hS(�� N�T"e@a���Y�p�Q\�8D0J����8���*}�Ә�<��D����!��rw@���,��B]�N�
���st<Gk��T�	����\a2������kY���0�_���}i!G�m��<�R�~!�[A���d�&oIĺy�
���;L��yܵ4Eu�8��i��Y��u�I�6���Q]����"Ei�c�Y ��3��`�φDM� �Ym11�
�7{_@�������
�,4\�<T<�姶l�ͷe��e�a����iL��0�~q4)WG��g52�H,Z�D�`�G�ԥ:9��{d[7��n���L�^?�Nb=4���t[VG��B�E��KT�(<c�s�Q�>����
�r�"ft������>��Ȇ�tH�J�I�M��Ny��@X�n�"���U�il"K�#�N��-(+.���'����g��D뿶��M`��@��LĸHĬ�`��(�����T�͊خZ���\H��Sֿ��D���;�"��\���Y*��6�vBq%b5���I�s*&�� �@�zG5�X�bĀ��䓎�6���q���K����(L�%�p���ӧK�h�ܡ��e�Sn�]^m�݄��hs���
�1g�}�mMtqS��.(X�B�-����F�ݸ	z���I�H!P�!~�gﰾ�&u��Cc�Cg�b�/�ߓn/�>ۖ9��~�3L09Ͼ7��rN[��m��H��t��?��������T<�!4Y�D�vV2\�@�>+{#"�tz�7��ɮ��y鎚�����?L�2N<ªq�ʥ�!�� s�ƻQ�=��YD��}SOTX}��6~��T��L�J���7�;�4F��A�!ڢ�U��M��wU� B�$��:��)[{(���g|Tbm!)�6Gz3`ϒ�����4���X���b�K��DW����k����8)W��ayd�ʒ�_ zћୋ�6�����+|����Tm{E������ӻ㾦GQBL\��'CH�	�::�ExAw$E�����Ɗ�� 5q/�����i)o	Gd���u�;�6��-�����g�ݹ�h��k��%��g�4�o͔V�T$h��5P+{2��
�q�w�TCL�^��DDz�$&l�uLn��##��M�ǳW���'!��2�SI
����́�4v�XnW#�_-�)ۇ�MCdZ]�{bP(/j!$ĈYh�洞�ϡ�<��Q���}��	� ^@���#�f{$I����}GLuL�*Z��l'i~��,�6J��`����L�����UU�������9��z�ʬ�Ԟ�O��_Z�WJ"C23.�D�� �V�G�`!�VB
�D��1�[gE�vH�!�B�1sꉙ�qK����6��	 ��;�O����z_Q�����7z��N;��o�����\d�����@Q��4}��������P@�*�����elő��Wyh=���h������X�kؐ)��Cl@s̽�:�XH�y��o�S��#�2Ŗ�E��_p��:Ӿ�Ҙ�I�2��;��_F�G�K!�*	?]��J���C��A����j��T���꨽���b�':���=wQT�U�����ס��
N�g��J]�L����Dw���NK\Cjお�oW�����s}H:��q�NC��Y�<���Ф��W�:��ۺ�!iӖ���M�g�I�Tӌ��������8�BFRn���Z�
�
�,Rc�߶ Z���^2�k�.��HA���\��=��	�T�z� &��`�:�#,%&�=c��<��Y&����l�=����Ǖ�;w��fj��7�Mؿ�kT��;�GL�ʗ�jJ?Q�j��Ҽt���Pw)��o�
O�R�=h�K?������;3˛r�JKUN�����#���:��ܗD�����BƧa	�d�'�ʲ��T�t�~��MX> 9s�\s��-/��ɸ������2�|� χ_�0-�4�����+m��a'/,����@��.`�Z��Ch;{	�5R��_�+A�%�Lh5��+�����uf��^�����{���%�4 _�I�e&L�rj�����l������ �or�Uzd��QIV��LTȣ~~��G���u��B�{YM19�[T�XI�������"p�e�*\C�1�WvF��p��<(J���-_��I��(E���=�{��-�qk �D5�Bz��?ۚF�K���g���n
/��-�ȰU�=���OjiQ��~�I�i��۟�\�D=�g�	�1��B�;��Y�3l����ڰ�~l�p��qW]���K���xg��"�j5��b� U�ڿ8��gӢt/�N�V����>��p;q��v�����a�*�.4�Zq�K�J�e��U�Nd�8�g���Ȗ���0+���"�<u[z>�N�|�?��e%�=Pw�Vj}�����l�&#]8r��W���Sm�{^��N�mz��H�*c~�uƬE�B�*�r��¬A 2m���0�b�����Yqp��~���`X8��	HL��'H�����2*��"��W�=�c)��O����JX�x�`��nj�td2��|
�N�/��p�0e|m�)����VRu�u*���V/1-�\�xQ��Э)33J����U��DU+��`������]��������:si��ꩢqƘR�nU?�u$آ�נ9�E fk��Z5���/����Θ�, ���L#%�1����;��uΐ��MH�ƠV��� �A3u�s�=mu?`^�ܼ&�ʻ��%%��u�=.|��7)�D#Ms`'%h(��~v��J����q��vV�ŕ�*&����#��PS��,��ȡ#�&�,���})��g$�?�γs����pO������:X��L�K�x��S8�J|8@�������v��U]�kmz@�QU)���:.�i�������$a��F���Z���> ѵt�e����/�m�o*d�}n��k��ƶ���1��#����n������c���N�-���W`ʆ��y~���q����E˲�rBld�mfL�+���.l�Y�48�$��愸�ޘ�S%cL���1��0m���U�d\4�� YN����������'�A����p�}u�J&?-����9�t��^��킗���ӂ>J[m�����|�i��Sd,m����[����.֊ݙ�2����ܟ-ٻ��{O���W�}`�:��ž�33��]�7�2�E`"�S����M��}�*i����X�\�VO����h�i�ޭ�o'>x��jL�V������.L��ڭa���D���F���yf|c��"j���/��
v��R�'(w��Т�ӧF�Xڦ�)�Ե�6Rtu�)P�x
$��� n�7-����#������y���=�OP[����9]��t�����,Y�b1{i���H+�p��h�IT����>�"�����Q��62�W�Z�Ia2���F��7�/6�y˘/�l|E`Wwe:�t}�~��*���tN� Ax;f#JIھ���<7#mwY�,�>�@�)���Gٜ��-+����Y#0�>�wɠ���WE�,�E��_2��K�xKO� ��""�Jo|t�l����T����Փ%�} �!b�q�~1����f���\���6C�ǁ:������R:��R:f��*΁_���?��j{�+�F~y*�vy�J���{�*�z�a�N^х���>&
D��L��`�K�BY4"0�tTF��T>PaR����#Sfj�1�<���(����2,.�q�㦪	���|�^RM<%�,��� (y3��9��7�6�[���,���Y��O?�-�L]~�ؑX^��4�71�����r48�S��2�t�E��G p���_
�ģ�ፂ���9���vAt1�A
�S�xj�"+���$eC���q�����T�X0��|��"�J<���������#��-�"k��bzt?�HK�d X���{~�0q���r�� �ɐ�\�W>6:ytl+j>7��tc���nA�Bwط-_�>�Fo�L'ē�sA4��#���!5ɳk����X�<��˕��Q���b����hJ!��%�I�3�ƶ���}����P��%�/�7V�ڕxMh�K�9l������U������\�蜴�D)��(HYk��o�"����si	���=�3G4�.A�� s����͇��\�"�ӏ��,������^>�&R��d�����!�BM�lK�f_-'g(���e;!��7��5.6�N?Ƥ$,3wj1�cR����;��9��#���� ��	�֌��O"��p	j�P��)I��#?i�P�5��NU�T1�0S���e+x�t1��(�א���_e ����Ծ����s60ư�p����R�؃��4�_O^~O駽7#�4�a�j��3w���c"��܎��Ey�R>��&��9 �9�Z^FIY	I8 �wh��H(qŷ0�2,�~^X~��G蔘���Zس<eo�{����m�9�p?ث���X�"A_j��������~F0q:��h��q�d��Z������H�軞�rI߆{t���M֨;xN#mA.��	�(�˵s�(��Z��w�Ҫ�{�PQ�1f��jEr�����Db)���F=�1B%��i_mDh@�[�Q'����#��&��ͭ���u�K	R5���������l�������gb�{�0V`�C�?ۚ!�!Aٝ�@�Mj� Ϩ	�_!-�SO6-H:'I���l��bճv(z1᱀J7����R��e�ި����S��O$X��0iΉ����{�Qb   �hN0�3pū�L�H4�~�[3qZ�OXR�*��q}�:V�О�cC-�g�%��ǌ���&��T�����l��^Y��"�+�I�f�3�b��-7���'?]`6Qg�n�dNyEɥ�$�+��\����2�+�'49�j�����7�RB��X=G&�y�˽)D��E>O�����}o^�kT��^+���;��/;�cmm�m=~�6�^��!�@�rO�=7~��Zi��q�ZE��k�'=���K^+�곉����-��R1f+/PX[���]��ѣ�`�W�b<t�n���L�Oc��	!^�F��5���K-��qӃQ
)�a��4$�)lD���;!�p�U�ШEy_�Y���.X�rd�����^.^e��ӱ��q�&.�-3���^�~�!��/�̛tPyRݭ��S��h����{&��v�[�H����0Z����0~fPcY2�Hɉ�c˴c5W��F�kdIT&� -����|-�K����IH^ �d|	ff)>me&�4��%�TB&��)��I��;@ƈT�A��Qӈr+hzk��+jc��
+ہ!�W"�@rA��t �F�f��"��/�@��+������jA�)g�;���Yn�R]N5��CK�!�nJ��s4{8���gp?�!�BWU�D�EX����w�{�}���Hg����tg�#T��
^n���T;���rHU�����ހ��;�\l��r[-�a����!!@�zF�qE���`���O��F�>�����A=�k����|��>-┱��9ف��l�WLVzB�6M�!���<��eiCwy����!K�f��f�ȼx�7X�Z0����e�E�;4�W�|�@	,�wX"1$�G�D�����x��ۣ��2Ҹ�M\��Y0-|�dDֹ�O=�z�9>c���;�L�
aԜ�V�x��S(�3Hj�1BR��$U�2xߺ,{����csV�~�z8�9.���f�#q��\���/׿!�щ��ޝ��`7��5Q���n��j'���x�gmWNI� �1n [|��z��� {h�},��O�	�Q��	W�)2�ٚT�~2�*����^Xg JN�@�pڰHe7{Z�^|��$-K�N�$����mՌ��K��/Yu(b>�`�NBi�=3�i1�9�:)".!�Vdv(�����O�C� ,�M(�|�1�:�S��䥒���|�k�0�7�Zj�o��Ef��Vw����X���ZM��~�w�=|�_���L!^p�rb�9���t�F�`&�{���<���si�.
�����l
�7�#� �1���rbU���M���XS�+H
�L�,���	���C�޵�Q���(�������T}�Θr�+�*�ݛ�#�һ�����-7￸�)�[�y��	^�;�D�}�=�@���׭����N����c���ǽ/G�����,��R�3	:�иl���Qm5X�*�&��@��E�F��G*� �%��s�=sӚ�c��|�A���g���G'�� +�=��v�YĤ�'�<�>b�B��ֲ�F�.�'��[YC�}�x��N�~l*;2D	��������}^b=�?�-�Ț�*X0���ȷY`]@v��m7-h�ýҚ3
}$;#u�ߵ|��8Y�2��e����P�3��c��}����g~ � �7�ۅ��4��=� nwڥ:�0�BÓl��a|��4�Eu�i �+tӵ���4��&yL����Q@�Ʌ����fQ#�g[٬>Q��Lz�R�ު�逶Qw����4�p]6�	�q3;dy�!x-��s�� �����|�� ��-*�wD���n<)�蒧0�2�Ow�i0��G��Y9��J�!B.�@kr�U�J�Ꮓw��]����wpM�-vB�az3�$ԓ�hif�S��c��X�9Gw2:����a
��C�,����m�k�\����ПC qu,-M�X�)A�s %&T��u�\��R��26m�p��H[[��_���km�ր��\FW@��[��L:�Q�'ȝN&-���Vj����Ŋ�F�;s��zw��y�/Aњ=����)q����f���������Pl�<�A|�!F�ӲKO7���5?�s��E%aq�D2ל$5�^fl�.QpW��J�[E1�4�^F�cU|=����=���L��M��pf�3��#&!��v'�xs)��	�Q��'�W�<a�$�X��?���� ��D齦5
��p�\LJ����$���@lƯ�"�n�Ȳo ��ed[fg�G$�/^��s �&�ӣ��>A����WK�1u�hd�QM,����s2�M
���]U��'%�BP��b�~b������K�-=/�\p��E������8L%.A��D�����7הa�r���FLn�ݨ�`_�}Jd��{ױ�Zf[kյb����z�0���h��bE��r�H���h���]'[IG~�B8	�.��L1Vh>(����b�ΜڳG�?p�3=7e`uw~���I5*����Kߢ\���ĒFR���ba�"�D�B,�Y��#ύ�B�x1׵{r�uα�pޝ��p�aL�A޳��4��)�e����k�L�}<�ʌ--�.x�|��N�#�JAo��T��e�|��Y��a�<�Jy�W+�
����N�J���d�g��/_��b�WG�d��A?��3c�J����׭�?|'��mF�,W���wi7ק|�~t|�n�o�L2I�]ܢk,�w#c�$B	
������+
�L[�y��8GY���eo=�m�٤��Ɔ4��3��G߫�f[�I�W�^ψk�	������L�!܅�Q���:=Ǻ��h��2��Dl�����m�H�����pk��y��������?�<����zZ�Z���O28�7�IS��K��M=�]Q����y_ʰq�`~�w��ȸ� ��{ �f|�Rf�Lj/��Δ#�3����񭲜������e{�5�-hՅn� 39TAv���������w���	.#��,|e}��>�5P�C�ʇ૷�>�h��y�u���,����"[��2���JGC+Y/���^b���)�J�Q�yP�Bo.6H	�8�l��1-��P>ԅ����Tg��4*}�H?��~�	 ���Ӈ���|fL���쳿�]p�������]F{:�a#@OW��a��ݘG\g��¥9Ml�<���Ӊ�D�I����>���VwY-�U��>*+KF-Q9�Qq�F5֡��V��l�?�4�I�t����F��aӀ2�*�a���%8���`���m�?-��*�� �K��ݐ*v��/Oa&4��`=��LVs��z��]3;y(a���R�\*���Pz��3��O�Od_�,J;�J�u'�����K��*����b��.��W��>����1�K[�:�3,����QE��Tj0�f�,	qL̑b�h�e��0F{h�i���-\;=�(�5N�I�D��c��\�O����!F��\��2�{6���R/e��e���5]�Xz�����ʖ�҆��ᭂ��c{�Gx��������p��[J,��rBQڕ�ɋ���_4m���,gO}�<u%��6ˌqc���\�]�"j�O��H��2���G�V-(��QA����|=~}�~?�(C�[�d�t��������vC\wVGN|�Ŝ�4Mh(��f ��,!�Vڹ�7Ӏe��]�q�ً��Ʉ�H\���9�֧e��A�_�6�cB�Z���`�l���T���Kw��qO���%Q.]�E��1��H��/7O�cƴ1o4���`�n��x��^���D�J!Û9#�0�).#��k�������_؎A�`V��_������xN;�TQ�36��E'��NO��k�%O~6�s�!���L�3ǧ��qte�/Ŀ���I;�|�;:�`�!I���yNC�^��{�v�	��}Cv��1��I�3��]�vQ��r�R'w/R�G=<��M���>����ʒc��%�',1�P� H��u��λ�3�H��#�qWF��E��_��hgu��4�^�H�S���f���`��a4��}z�q�O�mہ�~ޞ��g{�~>Sl�����3,DSw(֛�3CKM�>�< �]̲��f��坟�d�h�0S/%�\�:"X&��ɚ�z���t*!.��J{D�mmB��7̍��mJ�/��Z���i�K����7\�G�F�`�QS��i1򯺑x��j�d׶��f�ɢ�+)s��d�;��*�4+�����7m��q�)ohf��.{����J?�݊�[MS�s(����<z�����.
h�"��<��{��T�[uHs��4��������s�M�����C�[iȣ�kjS?9���Ł����v�� �H:�G�|�+mz� ��o��l��W��4�8B}��|9K�<IZ�������r�����Jp7∏2�ly@�|�,ňm4�����g��mQ��z��i��ԅ��~��Dr�����`�(1ݲ�[Eip{W�-��Ǭ����I��	M��%�x��^�e���{��C���l� �** M�|�8��3O5���Vx�0�F�a(�m���4�I��Њ:v��C<)?��>u֑�����&�֔.����``=�=�=Vm�ѽ`�݁�T{~祠��.C���`����0����z-��	n�Qtm��8�Q�����fg���Y��y�X�aϛU΅Lg��-�*��Ws�L!z�����TJ�*��4��f5����#]��U�i+B�u=�bĶ��Y�:�`�%)|�R���V��o�g��j��/d���>��_���0ůT�%�˩dD�z�rP����9%3mfY�K�AqJ[�&P�~��N^(�qw��8� �ǟg���A�w[���N�$
5�m��jL$I1����u�	<[�n�4������#�N�	&좭˟�v�U�6L�>�ٙ'Nfs4R	��g�S/��U�2�^,���el�*	�W�˳�M�VQ���2��%'{'�JtB��!hx�$�]��M�Q!�j;�ӟ��,c��ն4R�*�wǘro�@e�:��YX��ZØ����Ǘ���HuK����Q�p*��B���_��Z�;�^λ��pzt8��5��[�u�v�k��]?Ǹ�!8���7�d��%87�o� ����'ہR?z?F6���SU�t��9�1���/T
�n�`�L+~���6^�+�V�Ħ[0	ƍL���pX���s9��d�a@�\�V�0��C�g�;w� uD��Em�W6��U��>?<�4`^_p>!몏s�V)a�{`��4+xB�s��()��w�q�T`���e�w��H�2ݑ{�����,�%{'���97Gm�'(�
F��Hq �H�yW仨�׺�n�W`ן��έ���@��%���������z"ږ�\�Rb[�� Gk;�M���a���X��Ljj&�=��s�f��D����B��i/rPy�i����1��}���w��R�3P�~l�J��)L��t����^�𶬽���]-��W8�˙����cO��[8�Y]�%��L���-}�&�v����+�=0�){�TLX4j��Mv�����3[s�5E�jYX&���8}"��>�ڔ��g%������ujP�jI�Px@�-9%�\v�HIb���F*9V�ܿ"��;�`�0�����=#�z�G����L"G������c�Ih�P�PSG>y�ϵPP��{��wY<]�
�E������o���K�1�'��뭕U(�nd��u�B��A�R�|�������D�y�W!�.�)zξU���H��9f*`�Q>���8z�"��i���6�_��W��(����9b�(������k8۠t���{E�,"��9��+א��䗹a�A����ރ��X�I�(Ԏ�Փ��c�X
�O"�q�0oɧڥ
��4'|Կ�c��m'�l��E��/�~H�d�|��aL�<h��hn�܁y���sm��S$��7��a�-��@��@a���(��#4R
J��E٪kyQ�"�3��+C��N����K�M`+��h�<g���o`ڠt�^,���L�Đ��Pd��bC�g S¯ݬ�'�O�?.أ8�߇�h�6�>Z֛����'�;e6Q��'�ʔc��#xi�j��4��Ѷ�IC�&�M(��h�t��]�)���.k ` �=bY�,4���=Z�weW��&�(:��#3�8NT�!�3�$�Q�hR���Md>n�E�/֪��{����o{0�+$=DR�G��b��g��`x#�������e�]�՗E��>�8�z.v>���J��-%���(��������gŻ$�-�M�D�^e������M��2���B@�z�
gjO?AZ2���@ 阔����R'0XQ)re���.:�w��!Т��w.h6`~oV���_ˇ/�4L�ɥ��:<��4��p���c�N�G��n��j��M�H��!�=�rU���9c͛���S݇���DT���ᔺ�ςjW��>_�nEp���#E�ؚ�X�zػ/Ё�{�RU�4 �����1�ىCr�����ӻ���Sw1�s�: �vw5���C:�P_�,�8(�o�5$c0��L�y���ـ˔��İ����fz����yg�����%��'����l�T��~��aX��,��t�e+���@ �Ͽ�ʶ�:f�Z`ܾ�c�r���ݥǲ���E��A����ECc�*�_]K3�ӽ��ȣ.g�l��joS�u��U S���2��" ���U3��Ռ��,5��zúݧ	i�Լ!g~���l�*L|�wX/k�����N���x�q?��nKz�\^@���Er���BѠ��WXX�OK�6��%%�ɣ��^D����3v*��H;c�E���s��H1�W�6U8��pN�]9e�n@��kGݠ'y�1�쵅G����6j�,ȇP��EAi�W��Q;3�5H����՗� �_<�JK�4`�~�V��QjH��A�� �3�>�:��AV��wf8�&k�;m6��t��y���h�mo\�v�����3�D��������f�x�4S!�n-O=�X�!�zj%�I�iЫ���&����i�/��e��gԽev�t����8�1^`�fV	tQ��Ш�38��a#X4;n�ڦ��]�b��&g���& q<����^@�1�.'����㙒M�2��iP�r���gt�H��>~7A �o�S��~����e��-F�;��7,tJ6d�>Cr׮z|L����+����`A	p�y��侀z�>b�-�$�j̨�,�ا��kё
5U�f���~u�&���� �)ج���(F B���{�m�u����#6��
����z�n�p��\mx҈��k��\g�}�W��M�p.�$�@�oL8��G&�Ǽ;��p��NG���s��aa�#����ީ�>t�;�����x&�k]�� �<�2Z�����C8#=&�be!�a4R�y��@��`�.J�|�lي��4�?��Z��u�D�	��x����T�?1ڿ��r��U�;��Á+~��r��ӳC�g�n�^ƒ�8ࠛ��%������p�@1����\�.��I�A1eiH�<����0N�È��DѩAWV�ט5�}���O�5h=�f3����\a��-��Q��~�u�o��uNm2�;��`/��Gg'L$�G��5�$�{_ ��%��ӻ�����G�(Q�"���3��nZ~�\��[i�.������<?���!�,f�Z	��>YƲ��	0W�R�����C�q"��՞��-f�I�ãˏ�A˽����o� �|w!̤��v�B��uX~�W��G.��}��6��_���C4�:.(�Z�̯!�s���O����p��,�|�m�ܨ�q��kq�F@i�M�5��1���6�jnˡ�f�s�����0F�ZN����4��R��4����nq����tv�8mB��B߭�[1�R5�gchv!`���c��YG��x�|�H��%8\���a���
P��vE���۞�a"P��B�Y:z��OOtⷦH��v��X]�g���O�.���r��~�Th�����*�`z�߫��4 q�ӵ;���Xs�:�Xek�Ө��f��:�U�NM����t�O0�2>ʇ)P?�z��[I@���0\D��#�}3�'����g5�\����8ʕ�i�s��a -^��z\���T�WFz��6��?1<�vRDU�$� 1~�y�턫>P�5m�=3�J�3+˄�n���'۝�J�ԛ�qJ��:�rNA�q� <[!i!����U.8���FME��ڭ���"Jka8�?���l��фH������U�[G.��6�0�C�L(�����P�=:��wb���}% ���45#[5�^{�fTJ�{�Yͣ�錫�Es���P��4�h���[Udy���Ce{D9
�Iv矼[�A��T��}١�~��$�����	($z�ܨ�+�����2/=mѢ|~�A�/�&x-�5�p�9��-�PJpt��]�`�g��l��MГ�5mFs	$���sk�Z���L=D`��.��٢�!"���H��]��>���޷��F�:���p*��N�+o	5�ب5ˑ��G'{H�u��E�~���Ҩ��VN��µQ�$_A���ۈ�=�}�����f�ev�"è�G(˾|(��峥G9W�1D0'?�Y'���ˈ)�w]�{��_b�E�Ζ��N
Y�d��ß%�hE�P�4�G�Z9�_���A��ilR��^0ׯ�1P����V��p�g�(8�4.�lV[#+��;�)���H&k.mj	�
TrL��[,n�������Yy�=�+�I�ዻQ5z,a��	1= P��NQ�ç�A�~_��Y�y^��a،$w�Zo�Ÿ�V�����7֣��L�Ώv����M�$=�����_���c�tWW�6��[�P;KK��-g�O�ͻ�X����C/��4����d*Gf�P1��{��)�����|D�>��K�U
�YG�=�ח��l0�H#(�i�R�\�c�,(�>_��JF�]O�?^����<JD���Ma��3�Ar^b���z������h1��1�n�����	�������w�ov�r�&��N��(|��c�4�j��+5t�.kPj�����@��JsP���B�T�5���o���N|��;��S��;��5v}�����^5��o���vW��GK��a��ّ���/����D�f�����r�#��=
�y���9'�:-�\f��V�W�AM������_HJ@k�>��j-�1��x��`�>@kDY�0�2OB��=|��;*�8io�����ʁۡy6r��z�a�E�ӡLxDr���J���C<�&t��sa͗I֢���#��C�(�-9�D9�i�w���"�fi�|���v��J���F1d���ٸ��eccxCH�ﰣ���~�W�Ӱ��\�e��e��Q}WEq��o�����u�<>��n�q=G :�2�l^ap"Lh�^Fu!���/pI��v
��bUE��/�
����d�/�-"��$S���Z��O�����l�Yz`ɟY��Y�P�R:uPz��LVMn�s�+�g1�W������`.n_����BS|>Md0m����l�m�"[/JwT!c�f��m0��|�U�}B��( ��ib%�D^�9g��� ����(.O?�:�g���2o,��i��J��4�А�ԑ3������j��pE>���{�*+xe�"���Nv�[U.�qu�|]�kQP�F�Y� ��v4�)��n|M�ܔIs3�W�2�c|��)6g�9�7P˶�W�(lY,_����@���"��cfVϵ]��-��f�j�n|���/n��<��:6�^���eIc�]Pp0t�%D2*(\w/g[�h6f��";͗9ojdXz���¦�/���"�g/���D> L[�W���=bM����rL0?�I߅���v=��
����P��F)�q�>��},[g�c*� -3��E-S^��gō+�a)�1����� ��T�p�)Z֮�V������pcP�icL8�OBg1 \��1��O! Z���^zA�j�^�D��u�gp�T�D�<MgOd��"g7u�cv��ΰ�ڱ�D�*��ƾ��TLy;���~�F��������{���^IӪfY�AH,&���Ծ���n���� �U�i>�ƾ���p�bJ��X���������w� א@N��+yr�/Ǧ|�Y,�F܌�a�w&kH�Y(�egSՊ��ͪp8[n�/G��$-�����U�yp���$!��3�N�iC��5zt5 S����[Ք�/�7�K�Fhb���Hk�&�b'�؉g=%�Ṙ�F
:��"ISs���:�]�ǆSjV3�BX���VuL����� ��38FLVw5$��g����
`�������e�~���Պ5!&�R�=؎*��E<�5�U[�5���9x+hHռ]�Ә6�(V����+�*�c����5P$�]-c�q!P
J��+'��{���Ý�~Y���*Qq&�ό@�I6��Z����/*Q�٢5����Qee�y)Z����(\E���$7�+~���o��	�}����Y"i��?�y�m����h�����l&�+���ٓق�S"��
�Hگ,X�	�UWe���e	���E{w��'����S��j��)96}�>"&p+���q/�!���g����t�w�Υ�~��a_��urr���a��Ѵ�2Sy����j��N�_�v�J攫&vϭ,�p��^��(<�x.sT�R��KR'zb?[̶S�3�{!�Że%��$�&
��:��������(�5�sڿ����o�6 ��p~m�J8*��17���� H4ƈ4��r�����b��WZ�s�4'�:c�N�!��6#��FH,�h�P�8����%I
��	'.��3 ��Dd�MV���^)�I�������ݼ���ǯŞ�D6��Ud\�t����	K7��0��s�1U�o�uk�Z��}����F��Af��`��Ao�p�^���_�8�S������M��)C���.��rCD�1���.�jz���U�H�%ѣ�k����k�0=�\;�Y�L;���@�?0.3�	�!H��~��O]8��63���?�a?�^�z,3��ת.��)Z�/�-�	FG.䶆׀-� הJ����1���B$k'Ԉ���j��s&�Ë�z\������]e7�|N�AW�+��|��	��+\��NT�j��j�J,�|��5�X�ҽ@h0I0��VA�pJ�"�,�^����|�@:�h��c���.>+����< \j^���-E�����u�mrR��O��)!Nd��ܝ��S�w�R�4����U�.ӉH'��F����%�*&$�A4!����\��Ү�n�P�ٌEfZiLf����^� ��Hmj�CUPEA\��^��e�ZW���U0_~AKm~�Q�<��Ł��(<oi� ���il�Ä뼟t��@��	n���,�z5���غ�N�k�T��-���z��|}��?�UE?x��J�����h�)�#�'_;j/Zؖ+K4y|D��&��!QO�ʂv(�f6�m��I�]��'��=��(�Ƃ|�S;~���+=n��u�z�$�7�H�N���|��٣��Ii�u�i����iB<�ֶlǎ����c��X���#�7'}�����E��:���*�l���[ҳI�*=u������J��2o�6������:�X�a�iǌ�.�e�w�{L.��O\�h_ʶ!�"��uz�,d�a�\�Ȟ��M���6е�����;Dmw���_�tD�|4�i`��I��^�/8�{4�=�e���*ij9��)���K��� Ҷ*7��1�ĊT�b\h������;֥!(C	\�q�?�q���Vd�g	�U�LYz�Ɍ����{=�;M&K8 sR���6�>Tl���B�$�"�O�a��F��ǻ�h�"ct��#t�������P�06�!"��:�^d�B(?��ii6�I���>���e�
�֪h�T�1ϋ �(U�o��'�rEn���D:�E:���L&�
)[ב۲9�����;�߮?�&��c�e�G{��� ;�d��υos �\q�L�D9���</�BM�+?�)c�/Db�bMf�����J�% ڢ��a-TQ�Ux��c�0-n�.���?'�B�>+�rq@��^�߀{��&����v����x�.��j�^�L+㕢�-}JaS��G:8�^?��×�L�,|!#���0�ʺo�m"�l���H^��-�
,����8e�p�%&��Cq�RS�*�#�5���C�P�d��!FJk�E�̞v.�Ts�Ԗ#�抑a�i�_���`�:�c����Gi�LŨ���E&;��W�r�ԥSx�G���:pefB���Q�M3�����������iF_��o�n�L'����epxI&�&�;℮������x��z��ՙ���$��Y"	C�o���ᕥƀ����x!���~8��P�jAPs��Kb^�w=px>CZ����Ŵ栌��`-�}49U����!/g��a L����7W�_<��呪0�b ����<u��3Ah��&s���r�Ǆ�${O"q��QS.�a���к˞��<L#��WZ��ԥw�I��LQ�q�%�c�w��y���)�r�����C�f��.�uD��{5k�GDRGs���� ��g��Ϗ�}ɵ#	d�ǽ:'"%�3S���j���#��⇶uwUf�*Ź��l�M<�sB�<���I�Z���s��.�7$�=�IH�����N�䣊#�d�6�ٮ�c��j���H^eU"$��F�Z@��Πa)�y��0TpI(��ԏ	@w����ݰ�d+8�T�[R�vW�%U�����l��E��aF�}oOU	�2���g�R�����>�ad�b�OFr�>�'.%�4�_T����Z_��0�x*LF���#	�X��/�~(���'c&�~�qr.��lȨ��
tھ|HE�Y�="�:� ���4z6�~*���{���^��6z�@���m�3�e��Tk�0uCI��	������F3J�w���X�B��{{0��;�6�с����+3��͵fe���#�`K9F����p�\opO�T�/.����Z�}r:�_S��I~V�L��O��Ωס�	�n�|�h���<�;x��w 0s�N GO�ė`����sb�L��j��c}Ig�N�և�lf�������i�y���H���]�Iԁ���)#�j^X���'Y�ٙ��w�x��Y��+��R`i&��da���C�
�cGO��[���_R��Rϡ����3؏���,V�u��K��zS(���Ֆ�[3Xț�ܦOɡMY`@������+I�n�
�"Ȕk9_7r�֚���(6����؃�ܥ8MZ�5c�BN^�*o�P�_)ed3cS����JŌ����/����<��{G3R��su�ڸ��̬$����� j!����ߨeȾ�0�����}2��m4pP1�,T�DySb�+�L���aJ�D.fyֻv�}����e�V�O��*1���/�+đ�Һ���9��@���`?u`ĸS��ͼ^�M��8Ƽ������P#L�II�ٱ*E\�`����UFT�c��|��]��[z�~D���O�eŜ3jMߊU,k�2��qg�X�Z7�R}�����x�0��A����F��Aw<�_w��/>-�ړk(:^<0���@�k�Fx �!�����j�v����:�N��5W^0���$|��2ƚ�G�I�̛��$�I��2��y�.�} �g&- ���S3q
���G�*dڥ\d�nTHP�[�\�'�T�67I���(�x�k�̀Τ�lj����n�����Yio4�N�?�h�c��ZU��Ρ�����h��=��S0g3�n�9I��x9�LZ�vp���%�\� �G�M]�>�� 6E��^��Ue�R���+���D�4
�U���j/���%3tI ��s���֙��8r����y�*j�yh�����H�O��~%�9E�W�w�fu/=.����~�?��ДLh��;Z2�=2�V�1��D&#��*�o�G�W��R*p}�غ��!�;^�9Oe�񣥡� ��<5T�t�������K�1J07%�q~�埶������E?��+#��=,`z�FY�5���j$���+F��}ke��U�TUᡌ5(�7�)HM���p�[���Q&�+W��t.�����p�pu����*�ax�)��/���K�̸���Ʋ����v�@iT��Bq1w(�e�����⻊u����i˔~�n	bm���n^��"U���,.���ܓ}]�D��~[���+�_�Z�3�-�,�/�˥f�T)w���!�M��{�S�z~!�">��9Fx:�\�-��������"ES@�eAjXQ����J�N���}Փ�'s���;ʃ�D�o�?�'ݛ����%�U�����G��q`+Z9}uD�I�9$JЍ~�X�l�S˭�R��4� �D'�Hm{��A���^�/5�ۀ����!޼�����J�N愽�1A����pa
�j�g5������Ci��>[��kWa���[��c�o��{�r-!���<�TU��d��=:_B]��Hd 0� ��5�S����x��FY�{��S����@��9��G���� ,:jշ���%Bh��O�a����Wv���G4��X\����Pi�����O[�P�`" ��J�����(��⟆7l��~�_� 	�,U��s8R=�.�L��v �x�]�Ä$(���d�f� ��f���]mURa�U��+�S�[6��{&���N�dG�R;�Z�R��jէ��Z�z0y4�?u�ɨ�5�#����b=��E�.ʐ�c��/�|@~i��ڸo�c���w��A+���	��V�.�t��t0��� ���n�>J�~�P�}4" ��D��� ��k�����-3����ì��2a篗]���M����Ԅ���lvÃn-���,���\r�\��ޙ[m���?�mcРn(�:�p���*-��ظ@O�*��z0}��U�C�,c�=�a�v|c.��yú���L;cEՖ���́sH�<��$�E�r��`�U�l1�)��,��O
P�1�y���8��[�j�SsX	M�n~����īi3�4�dp�)悥*#te�T>�P����֝R��KB{S����%�w.Y�C�m�e>E�z�B��]R����`9��ռ5��-�h�[�����{>|��7hq�-���_9Cg�4P�M�u$���PH��
�%�����D�U�7±��?Wf����сH55A���{gJ�D�-azc��bi�K�cJ�q�Ab�GTd$��^�y��P��Y�H��S*�H,���z��PTF6p5zq*B|̄���&@a5,}LގU�����X��
�s~������ʋ����03�5C2�J���;�T�;Fڨ�����!hWv���P��*8u�@	e�Mi%��J�+4b���q�L��O�kdh������>�b��
���Y{x�����Bc{�3��6{SR6T�ي�4@(���������'��K8)�3q���S�ɻ+�����O�<����0���\I�5l�h�^�[8��{<㩡�|�N�6g�-�Rb,�^��%W��I����QpĆ�=SEsx��E��}���C/	��k�bVP��ս�ǿ�Z��9�o�{o3��NX�:(��	Ƿ�4��a�bڈ�?��d8���V�oyr�������	4cM3$Cc|���og�+�^���p�P��֢����fX'#ga ��_��vz�J�l��lB��9����]�,׶!ŉ3�K�<�0W�d;�F}��ln�1��5�h5�� ��ۓ݁D�����c�PҩP3��?x�����X�y�?˥N��)�߼���Jg���0��d����o^��z�c��h ��v���q	��Z��""�^I�R��Ϭ1�H��/�{ԉ1�#ǐh�A�'���u��r�����<5f/�I����тu �:$"�}Y����3� ('w�0��JO��K�8��+S�ц��u�}R�A�S��`��t���F֦Y!����lhȫ��f�۩p�a���S��E�S���eJ)�Zb���n�7T��g��/
_�f��^Ι�*Mvh��:��؊��h��j�<��]����]V�#t��B�G�=d%O�y��9�P(��NK�"SJ�l�G�q��Z���ʇ��.�ڭ{Y��:sC��~h~��3�<k���kψ�!:�3k:��ՔC����@[dm�pgbs����M~�U���
i.�ǲԮ���5D���Ο�Q��\�j�0����V�_О�u#
�LD��|�0��N�1w4܄�!Y��*�/Q����L��:Y����R��WY}j%��	e�|�O�iXkר9��QB�8l'�-k�����X��uM)	�^�/j���5~\7з��<����ymi�T�o��a�Ö���1��W�=Q�P��"i.T��j��o�QϫVJ���|� �@�F/#y�I�r�H��i?�Z�2�
����������%���E�n��J��]��p}4}��e�B��M��J �B{ɉ�%ںf|fz��/`�r���4�C0�⭍��:�RS|��E#N^�	��>k� �5px�*��8�+�0�j��إ�8���E;>ru�j�S�	;�idW�m�k���D0W���nƬeB
6W-"����=
��8ڦ<��qg��.��ǿ7XFO�1�Ё���ޣ&٤1�nd�**��xʣGs���y�	7y�J�Ń^�k��Ӄw��41SV0@v[��|��!`������ ��s�V�����]@t�����*���2������B��b� �{ r�q�*�Qa6�Mp?���	l�]nW�� ��J�8r=`$P*-Qܕ����%b��� ���/]������ ��t�Q�K*�����b�$?h�]\��W�CqA䷏��\A��#����B>�5��w�d���Z�d#w��˶wu��t�P�;�Ok'њ���_��ަ�D�2��s�+�1���܈�ʌ)��X�YS|Js9U�mj�jF��j(~s�����yZm���Ϣ�y�B�����J�*�YQQ��+��Z����J���}XZ�ӥEfTl�j�]��+��Q��@���ۄ��Q���}v|�7�)�;�h�b�)���|5�Q�s<g5��P�k�>�@#87I7S��L�l��=)��U=N��>B��T �	5������Q_Ml���QF�4<m!6<ML��\#��S����*v�@ ��n	Jvغ>�&B��3�B��w2�v���!&}��:)�V����t�2��V��OǊ&5�p�V�'�F�zc,�Ɵ�N+�b��~2J�Dz���W���+�"�z��=$pN��~I�ҔBd�v�O��t ,	S�Vu�4�ޒ��		�Η:���F{���)�.9�9��v�HU��_/3������L����lj̇y�£���c�D q_��[e���O1M����~��G��	�2���Y��������0��ԍ[��,��C�*�y�L�L��H��q}`z�R�k�qQ�
>��@u\�k�@�1S�վ��Wp3�TnFӦq�+��?���?U�����"�K_�C�Kl��²�}Ί��](*/ga(}l9�w���@���f�x�UҪ�@jz�Nc���J�D:p�D�-LѺS���T�Iq���!Z�i<����I�Y�b��[�;��&»c}H �}��Cx����"6L�_L����Du����J�P�<��FK����S?��5����t���a��-r|���_���Y�f�*��K�n*��	��LG�,�K��ǁx�?Vz���Z���;0`}nN���o	�Y1��mE~�ay��:ЩyƢ�U�!��?Y82��J�p��)b�S1��s��s��nj)�3�h��d�,���[������t��;nj����$9�:���A��q�2�}��$�F(ٝt��.�b�1��f=�uC}w(~Н�ʘH	�wp��j�n��դ��?�4���v��M�YW`}b��?��F�[ԗp��(P^�i���,�v�#07����#��l� }��0��~2�x�ٚR{��#%���Q��������n������Ӈn^�d(�/�J�8R�?H�`I���I��y�f��CP�+�O�p�������-T֪�ϔ%��j @7?��L�a}ک+'-�B�6,�F��i5�Nr�7J����E�%;pvE��&��)q_�	`aQE�Om������ZM�%i7X����֜LpJ����CCA�q��dWW�`oNb��Yu���I� �^�f8i;���#�<�X�k2�{����QS��.@P�<��?4��s�(ܕhK��t�5�9���p."���J��kzT3�<�����Y�Jx�H�mL<��'�8&l}@T��.sAN&�s���MI7 ��#��5��-��K�F,��b:[��#K���[9t�pλ�w�odra��=���0.;;�W� ʪHSN�E��;��p+��/ ��/D���}C�t�����g��+��X�.B��#n�w�jW�Úk�өPy�C��~����[f	�d3�̮mD�ݿ*->��T�+U���Ǧ�cwͅ�!��)����I�H��~��Ĝx<��53p��
�ùb�z�,c@�j�Y������]�*�����\E�i/	Z��.��k9y��:����)R%���w��|�w9�J�1�ݢA��3dV�#�V�)�p�	cv���:�a�!�Ҥ�d��0��`�=Uv����~�n$�±�`�!Sa�ua��L�j2>{�/͌���v%E-A��b�5Z�����72i�g��X+�T5���$�a�/<Y�0���!��%}h $?ڰ�,İ��S���?��j;�SFN-�P�P��4����(��}
xbS����IL�y_�{�{��E�� ��-���N�Ջ�I��@x����M�w��e�w<��QzDc��58{ ��&�Bi�|��|C����tb��C(%�c.��L�� ��^����N��HcW)���n:.���J)j?O�~�=�b����#�$b֥'�����)zI��8�����F���I�����kU��)'�z�fJk�������?Cn��G����/7�e$�G&��u]�%�O�'GW��� ��1~+��U����$pq��M`��\�v7(!�[A}ɰP�cg<m���ğ�r��Z�p����v&��Y�D�?���5敷{h7�ǔ\?�0E��8���f:�J�`��ٯ�켺��4oA�\�;]�qBu@x���s�(u��x��$z�i�D��33J� +�X�'v@���/X��Q�]P�F/l_�8�}_B=YABi�L|�6lВ�-2I���#SCuC������}��Gn.n���������{�3`�L���m����Y��Ey��8a�����yE������E�$j\T��r�U�<�~��P�"��x5mk(p?K���,��`�҄����ۄ��=��$��45�:z;Q�8����;�*<�#��V�N[_ӡO��e!%cmD|u����Xq���1�S����p&�B#�w����ӽ�,�.�'��!�4_��Ž�l��.��֯ �KǤE������\�&��g�e�6���v��z���[ۋ�e=�@QL�J�YO*�ד˙^e�����p/ ��gw;����H��~Tҿ��F�E%f�=��g�A��`+�y����N?�mMvV 3��h��un���6���U�(�6�\@c��A�2 Y��{|}i_�.���!�s5&�����H�*�i���zO�" �5t�@�����.dW��T��̐����c�A��q8kߣ�v4�F�5#ܼ R嘒X965���,�j���JL�ہ��1,eD��l)K��̙,�J6O@�GP=�j�"�nA
 �w"` C��.��MO�TB�9)}�1���$ ��h�4sf�(p�^�O�����"��P������˘Z^8;H�sb謱x�}̿�;�p�I,�K�]���S� �Ch˧Ռ���/j���.�sF��9`0.�TH�����~�K�ɇq������x)�nEB��M�(݆����G;|(�z�e��q gj���/,OÞ�E����/i�H�A!ɳ�*Zjn��n.M�'����մ�C�)ퟑ!{y����K��h�9
�q������N����O�%���S-ׄ�>����k���}7��B1ڰ���}��:����,(.o/�:���H�Q��!������q�S�
��a�����e�c�Xo~�a:��+��̓��x�R���:Ǖ3�q/�f���nQC+1ƺ��+�O<�`u��Zn�Z��<`���Y���D�z�'>؏���P���հ(�Z�֊Ak>6��,y�J��b+n�K�0�'���7|7@�w<}H0��d���O
�/_[T�N��O��m>�1XImp� �MX�c���ڑZ@&#3��9�ҽ_R�Q�W�u,���F��Ъ�3�~�
o֚� ��8p��}�n��>ꤱ�#_���7���!�썀Ee�C���O� ��ad�1]�%[dA<��.��1ɑ��]�wȎN���U�~��^�O�eU��x���W����g�>3?�:]=���IK��Dzo�Z��Oߪ?(���(2��&��+�sKC(��ٚZ2�!�z��ҭ#$�ܿ��LpKI�:���iz����X������;��%R�Kf�{���E�e�{Gs�X��z�J9�ݠ;�,�v#��`��2I��ޫeb�����D�x���n~P�^��-������>.U���+�������!��Z��ThG_ϛ��W���}�m��fǗ�"��"��$��5�+�|]�?#� ��A�4���HT�]����yF>r�g�9Fk~�*#G�ۿ���kI����i_eeX�xQ\=��X	F�T��d7@���t�����z���pC�R붞����.��ת;�l�["� ��l�BZ�)0���Mh�J��9$@w�N� n�iމ�_�3A��/�}�g�)FY�ej�zJyM�]}0�k{��B��!?ꬩص��Bx�\�Uod��qV� {�1���<1�eE�B�=�cl6V5��6��)6ۻ�)(������lK��p�89z"�Z�OU�󪵨���"X�nnte�ᦟ�<�2�|��K�54Z�~�k?{���w\ +��OZA�sΈ�k����3awPRL����|�Dh_Ϗ>V+'V��Ѻf����6q�
n0}�vAB{,����R1�'�v��n��O���u���6��b��!�Ir1$��� �j�P`#�F�1����&��H~�:F9L଍�B@���|7塥�����1���Y�$����m���#fƼkM���:T+�/۵��U>S�%s��z�C6f��ȋ}�w��,H�{hcE9�U���q1x��~�3��`���t�l�z \I���6AH��:�R8�#���ʪ��O��k0�m�7�玲��d&^A~I��w Ҕ��~��,B�T�H�p	�O��{WE���r����Ҁ'YUk����W
*<�9&u�ʆk퉏0�9S1�lK5��3��G��9�i^�0b�f�[%��R����+\�Io��l_DAE�z���O��TnA"ք�ߋPi���D]�+UɊ}�|-���W":���gn|��&m��#$�I?�Cb!�b�NN=NI�7�b�]�d�"H�$� ���ٮ)jL>��HY���T����V*�<�s
 �D�=8c����v��G6;ډm��P���i| C*ץ̖J�Q�1)�\r,i�{]>�{��"%�����h�'d����8���D?�����vD-��9~/���p�W���Z^m�=��;�k��lɹ��+4w$k�ZE �5xiy��RyZ���׳�2���G�Ry��h8�g�CD�]�����kCZ���,gJ��y~��+�+�	<�rJ�̝���O�
��cܷ��S��#�WDݺ�[lv��+�u����u0�Ɔ��y�`���J���m�)[.��BXY]y-���tƋ-�[�3�ķ������\��o�������M�}�`J�ڥ-��kb��LC�(���$���l��	\z�R��BP��ȃBvzE��5X�}I.u�*�cv�M��В@B�ǒ����'��/�����L�h�7j|�����A��#� W�>���p�����ӗH�һ6�դ�h ���)�
v6��ٝ�-�����
��<*��q���y­f���E,��^������e�6�� 	s�ܙ&J<^0�w03,
�B���s�VxHx����6�S�|e� G��:�VI��"6]ڕ[��1�|ͥ�ݚ�:%nf���up�lf��ܯ�:���w��#��䆁�F�x�l=�wp��%�`����(� �u�)���>  ,�������bR���l6�s}����{s�)]�|��[{寗%T�h9�vd�|�uY2,/pm��C`�
F��W�����sr�"u����t�/W@�t7Vo|E�t�hPP�~���T^.u�F_97�  ���X�%�d4: ��gM��q�5y��?eW���jJx�Q���ڋt�� ��=�l6oN�ipѶ��=\�g��X |JX@[d���j5�:��@�����5D��ƽK����*��JBQ�ҎW��]k��4P(Qbס+K �v�w� Д�q
C�_G�����"��p"�s��Z��(�a���^4�Q�n8!f�3`�c�<)\�T��ur��ր!�-@X��~�Z~S��S���[�_���\:$�R�IW�^���o:r	dD��|d=@���L�s����,#V`%��>ۄ���Ibrm6>��\�~�U����?����if��C����ݑݟ�g=�ԡ?l*A������6ӑ�'1���CX���>�c�*?#�P��'�'��)�4l�wEFZʃ��J�Y[�5~ޕS�Ęc�$�TS�*�@u�뻱��݇�Fk�=�C��6� �d�ǀ<�t&dZTjt�(�����Zl(�r�8't��
�J�������0�8t�5�������N��M�9�qY�s
餓18���x��m�;w�)&Z���8�v���_� ?����d3��^֪5����3޳&5ڟng5�� �ao�?p} �T��f-S~IlR��#��!���>�=EW�uTb(�Ú\Y�q�PS_�=�Dla�S��U��LZB��)��M���!��B��cu{��p�"��%������d�g� ��ֿ�o0f/�E뀔m�����z������h�o+�\:�,���C ��P��s��a�7V$�,��2Z�~�E/\aG�
��:Vmܳ� �z��Ŕ�CJ ���U�Z_����j�C�w�{qfY��`*l�QϮ`ؾ�R��z�z�E�7�*�Xw�h��Pĉ�c��1�����i�x
^�[���*�`>����J����C�S��f�����<����M��ه9���}�ui݈q%Gɿ�X7�ǅ���b�O{���f0��s���j>�^V��}i�ḿN�"䰝u5���}YX3��g��U�D�(��Z%�S�̹t!Z�����v9-���	��s"s�FuH��uL�#M0*ڨ�6�����͹\����x���s!�L�� 0��D'��Jc��j0�������ο��M��w���7����m�.����	�a:�Y;a�O"1�]�tMԦ��}�~�.��̅
�h��h��Q�G��H%ߊ53!#��§H��h���E��Rb�ʔ�71�����~��۰�,~��QN��S8C���V�#r)_�`6)���S��b9NO5X�D5E:��8��#�:�	���rA��6k�g��G�q)���1<�x�()4Î+�c���'���|�_�}��6Y�Ўl��,���c*���sv�r6,)��˓[���|���4����ޭrxw��/8�@)l{�Kt��l�S]�
e�����.6C�o�����y��~�j�y��f��Fѭ-�8��(���S���N��ڸr���Xؑ<,�DzeBY�������E���ˤ������HK�e�e~�
�Q����_�"�:&K����q19t�ztI���3♍5}"�������z\�'M��JhC�����k�R=��u(��t�`i���39p�ڳr����8*�״��g�E�L�̹����&7ʘ�ѭe#����1���2�y�ym�]"����i�Sk�(��=�(FqX�E��(�[,��R.Ӂ�QoM.�����hyo�	/v�����*'L��Y�@��͸)0�ԭ�=�DR�t�xt3[�"M�^�t�-cu
��bsV'�Є����T�э�N�9�L�8|�h��q�>�-��W<ky�{ɨ�3��(��UO���y�������yX�^�����A1~D׍l�b�9�z�������]���c�.E�E2��ɂ��/Ϡa�bZ�6/�bQ�*ڃ¿�At�Ex��YL堨��;#���H�W���t�m��:O.� �1�)�����=�IaL�E���&���.WR�X��}�:4<9��t�ŉR7m�=*1TC�\Z�ߝe�5�o�:���lM}L�z��U�$Bct>�H�Dj�����⃒�j_�#Nn���"ad$#����AIs6S����G�{}�c��$޳���~ԋc��g�T?�u-)h��F����ӖH\�E��Xk}����R�N%����K/3�~Y+_U�Fv�a�O�@�m\�L����ۧh���n��������*�m�gTv�?ʪg�C�����b	C����H������N1m��a>$o�u<���״V�P�ܳ f�
|�ԽU]�)��.�s���������zH�$��O��C�A[j[��"_�x+tp����j���~��̞BHS�̦o���.�%�dK�	�]��U�C'g-�����z����͆XI5���!���k�H��4(��&4�`o�eq��\�������ꚸ ���� A/�E�h���h?n�p�[P�>CD���D�́�J`�� �IQ�tW{���?�ݤ,���N�	㞂�]��lY�/Q��
Ht�+�CտWʄ�y��)dg4mk1��%��Sq�����?���\��������R��.ms�g�n>}��^ r<��l�����.o��������H#SD�IM�2����]mmhz>u5�_)�c}�n��>���#9�<k�鸝%�6��/��H�c��f�@cvV��]ن~=2L�e	L+ob�ٮॹ=��2Z���*x7�}��kv�_3!`2u/+~<|2L5b\�5����.E��㳲��G��+�J/�\�m��:iӨs2��hh�DɈ��y�g*Jr~��jpL�eg��Θ��|ۂ5���H3�*c4����c�9pn=�
�P�r��<�W/��W��Ć���ro]m�)�v�}�87�ŦQ���&|�$���**SNp�C%٩�<sk.,���!�^��H������V�̲`G��W
0c��]G�	�5I��;)̍�YEY���<�l�t����$��u��9�$ �5���+ý�w��P	6��pw7�	}Y��AOnAf��B���ꧭț�x��h�/C����xL�WKv{�:]t���Ф��eTC�FP�]ke�d!�x8����42�Ym��H� [�=��n�j}�u0�p���qu
�:���G���u��-L�
b�:Ͱ�!�	�ᾹAE+�У���z{ܩ�?N�#b�� sB^��}~������b�����}kJ]�(���GT��>%,����%��~ӣ�FK��N[�gu^��/O�Qݜ<Tơ%O�l�N0ˑ�z� �B�C��-�՗�~�� �ᅇr��c72?՞� R^��M�B�f��jq*��N���$;��%���q)/�A��+�G%NỰ�(�*���4�c���9�Ǭ@1��wn�O1����K� Y�wZ_N=��d��C��bv�����z��r�g�����U�jZ��5��~���[y֢l�&�01u�2�ek�`��.���=���Te��Ms��}B��˅��ˇXT�,i,ˎ��)�0"@�1�JH�QJ��
��®ݸ��,q�I��<C>���Q���i��1��{]�rJ�����z��N�%7m�%� ��I�9�شd�`�:�aL�s��ӂv�Y���\����D��|ɣ�]G[f��`,AB~i[�=�*�Ű��kx+?4Ũ��g����}��AD��c.��}�_K<���}w=�7g����T�i;/=@]Y��U;�\�'��>t��B�(?⯨H����ɩM��6��ү�f�N�jk��Euu0���Y��-�7���uUl�Z���H�١W��،M��o�T�˴#�b��������U��� �wtv˓H��@��Ӥ��Q1�hz$1��G/���X�ʚ����X��,U�{q�RA�*���5+|_1�U�y�P_��TɊ?�����h�B�u�A1��KR-4����/�B��4�]�띋1���������k�G)��8��/��}���&0>�f������K�P�η�D!����o�&���Z�s>&��N���E(�CDa���u�3�@^�O��i��2Zuj��m����!���p]%��1���t{!oˉ�#Q��иY��`(�7���=Os'���ۼ&�	�O(��٥�ixMI�8x�4��P*�Tߤ�6�˕^��S�d�m|�{�(�Ӌ�٥@ӵ����_�����`HO9�]��ß�n9_�X͈�u�ծY�e^M�?'Nl6�#��Qі���ZäZ��f\��E6��8]qvu�:����K*��m�j�i�\�Q�7ћ>9�; �|J��/���y�ԅ������U���nٖ]�x��M�H�����p+v���ƫ�<	'����u���)/b�&0�;X�>O���=�nit5p	�Zj����̇��Y7��	��6�ܩ�_O6,����ʓ��RE����G/|��U�,s��0Z=R�:��=ڢ�ş�I�m)�K�y�C	ڎ��5Z$֬�ꤨԁ0����8���I�`w�d��Y�
}�!D�����@̘->���X}���4Zޘ/9��G��^��������]:hM��������̽�7���t���yY"B�c���/ O$[��)�n���1��P˅�#��js�~sՠ�p�|_�3��s�;���U����C� s����LHi���hjӍ$��l������]�?S�q�o�@�A5;�۰ch�<�D���|��_�q�G��zPGr���탊��97��I���h�1p�3D�39g,������~��*ة�"����=�m_ƚ/����%�>��/����La��7�W�I�q�i��򉣆%�t����f�X�'8[�}�4������Rt��8��]�{uX��Z�h� Ra�c��c��@
�_�G��Ĥʈ�b�o�h��8.�"��*��oV/�B�yvf��]��qʕ�d�O#��ؘ�	���'�_�:���=.�N���\��D����b;kF:��۟6|<��3P����+���m6���m��H�����Rf2_�җ&k�>@�a	�v��_�i���Q��w}~����w�a�ӝ[� ~v�����F��B�I�C�W.�H��w���a�h����"��	 E��/��C�k�����o����9�����Vձa��DKh������ѓG�愯��m�l�l��� M*��x�خ�:\x�/X��:o��m#��P-0��-�J���_ḫ^�E�������F��۟t���^�~��2�y��V��^�йD�&�*�'-���'8/�}�Յ!A��Y�V�'x�HZB`�;�b%�_�8��������A�.�c�:s���♗X͘���
�3�z�����l���{���?��|6���2�,,��e�|.]��l�O�>X�/b�U����UƓC��J�t� %�M���d��wY_��b�%�۬�Id��>�r J9J]`�4`]+����g�p�4ew�ϑx-����J��"e��qU�<WY�ߟ�ǳ>�!���a��F��i�s���U��ų��=�ش=1n=���|���OE�#���h��Ya��!ҙ!���Ǯ�WGd�l����㪦cn���q�1��W/K�8�&q"i�_��!w��7��%����b�W�I��S�9M�|�돵��r�e��ԱX��*+�w��i���Q�#��9�����}�A���"�<�|#�gkw��y �Xg�FB(<8���Mt�i#����S���g	kK�C) �u:ȳ������/�͆�d�F6��QA�K�:���(l��$dm��\!�G���+@�˺ʞ�<Q���}����u�(������5�U�(dXP�!{�B]�W��mԙQ|س�6�\�:~ݝ<�n��"j�^c����>*�O:���\�ъ���VR%h�������|&�v�?q�T@�c_�f��&�TD�|i�Š[�xX���-��Y�d%���<�6Dݡ��+��?ND(�.��8%g)E	b�������ڗ�(�w�&�'v:�6�ǂ��%�J};w��.}������`bmZ�����Z(���=X�7��mFm'�[��Xlv�M�{�HGIuͬ�]**��᜵���@��^3܀��D�]���+��x�_:�syÃY4��Ta�<E�G[�J�"�>��dR�L��]�]m��\�ؔkNA��������nX�%���#}�V
o2p���b�~b�����)�U�Q$yQ'ȩ���Z�ϋ���d��u�׿�T�c}�;n�m�x64�� �&�?pO�O(�A�!��_)�v�ٲ*�W��n�+�`?UW��y1#�5>ի8�%-o�f
� ��QB(R��C�#9,���Q�F1���>U"�@��?cuy@��ۄ.&��V+x��H���$1���N�R1.".��5���V��s����L��A
����g/wp1���^�Gp���QpQ��fK������~A��6�;��n��xq� �c�PыǢI��	H<i���֬L�Q�0\XѮ�s��pR+o��rw�V.QGٙr�������e6�M�
%k�9��f�4h]0D�h9�=so���.���'�'y�:Ғ���sɡ�?�d'�]��ѻ�h�\�+�y]����;����¯�/hlL�����d�1�ߩv	+��@�������>*bUq/wQ���Ơ3��.�T������>ދ�F��E挺���g�!�k���H|K�F����l~u�����Ϡù�i�uil#�b���b@�;��ȍY�c��涎�?��mm�.�t+��C͑�Sy�mPN��h�K	%�I�-S�O���W�50�y��)������V�ʨY]��^"s��:��no���K�.��zD�K!#�{��ꄅ���6̵KD�,sa�48\�DY��_�*э;9�jUc�u�,�z�7���q�ztj~����M�R��3�L�#W�'����}kh(�&��:����X�ݾL�3���_��d�|Pv����	��aY6c0F��Â��� �,��'�]65�jN�k���^;T���/"���P|+3�rM����)���e��εۂ��X���q���9u����n�V@�sQ(���#���^ZzV��LR��f������/�JFGJ߂��R��>�d`�P�;F`7�*��.�!���j�ɹ3G�$Pj�yԵ����Z&�x>t ��8T�>1&f����q���>_\�Œ��ni��5a��ڍ�)l��
j!N�{�=�g�nT��}k]��ñ[d��b��8em�Ƹ���Xx��uX�xb�-�@���$e[T!�D�U�Me��jK��D�>���$��+��a�ǛN��wj����0��
ډ���o�SP���ŷ�'��߆�b�ܢ8H�B���p|p;AU��jcIu�T���Yr��D?�Z�v)�C�oK_�B`%8\$D�9�Jp�dd?$�ɘ�:��xK���ٺ�]'AYISRQr��{�y�h27��/�p�!�B=�ZM�k}�k������Qu鋴�����\v���M�|U�Ĳ�1Җ�)�$H�Jk:[���{����D�Q�^�g����w����RV�ۜ�Lw.�oi�������n�sZ��#��e�l��}
��g�	�����������G����-�n��<l����^����j'�!5���;9ؒ��LZL�{KV���0e�%�ix-�{�S�'�����I1�+��$w`�k,���c v:F�,B=ɞ�D��/�D�G9J=�(����C�n�M�6�d݋)8z{�Fi�)m�=�{���V}ۏ��Bw�i ��
/���r�Ǯ����Hk�8���kh�<��O�5%��1���h��m&�R�(@�)T�"�_^oF�}NwP}��%f��b�����r<]}w�M&S��V�o���Bl�l�ʄ
��3g=��A����k����`~WE�&
O���[H���@0`f*hE��e�ᄏ�>�4�s4^�-v�����EO��`8.����ųa/?!�5��i�"[�n5 ����r���|�f ��X��q0H7q 8S;l�����Oy���}�����xGs���m���[�dH�A��L&ٞd���Q(��3�܅X�:�,t�Xz*>�L�:����[���a�'��{�Wr�$!�irC4�X����,���΢����~��8�5��W��ű~�G��.�AQ�����������V'�^ZDy4�F9���H��MF�`a��n���?���'\H�_��.��O:g�Q0�-wj"FE�2
�b�~<��]TZ+�ۀ,�	ؐd���5+*JepY���]/���x�W���Kc�(���ހּ��/:;���H�U�Qn�O<`�0[ e��1f9S�y=���B]k�!�[Es�N�A�Ot��޳��TNǀ1Ǔ����;�@/0�w�I���͹j>��O*��|;q�H2�̛X�- ۊ;���H���<#je,[7(��	���j���W�&J�&k��|�-��,6:��_��]�Z?���J,��LKs
���Cp�1��Q��m�}T���ŉQ�lM�6�����f�q����bm�/Ҵ��B�T'���z<׵��d�h޳J2_�0Ԉ�� �tNj�L�ȣ�{P���)���f*�X�A�����N�6[�l�&33{C�[+A\i�#����<R��b>����ca
�t3TIM�X�V�_Uy˷�(w&�īu.F���	j	��&C�"��] ����3*�BI�l#(��.��5&�Bk�W����{��2h�a=C
2��c5Hg���U�e���u?ޛ{	B�b��	דn�(���q��KQD��,��qK\a��[+��W�R���nŁ�H�z��c��k�ٝۖy2;@�L�ne�l^�2+�s
��=P�Uxa�A���&I��Lܔ��ȧ�u�[V'o�"Hѧ���q<���]�9y�|2��Ӆ�f�� �w��DS�s������p@�({̈́�Z�J�6&~Ko��/,��J��>:�	5l�1���3E%Ȉ�`�P�/��0U�L�'�H��0�i��<�4�Pf�af�H�bI���Uj��U�>�ɤ��_s�ۦp����'pc�:�:C�!{bwH�܉C�Q�	��DH�z-��'EK�__} �Y!�ކ�H�F��:�;�U�y�)x�ݬ���6��G��yWGx� -Fձ6���J� d_+�~\�"�8S(r_b��p#�=َ��v����Uڸ�v��"բ���?��2|M}Ｔ!����것�|o��E'б���h_�c5��4�<���Ï�s���9��l�}3�<xL�#�4�(�IӴ"�A�q�Q��:dE�D�v3��A`\F�[�j�U���)=�!��"I�0zw<�m��!$��E�)�m� ���J���؍�TP�9,k�,D1�M_a����2T�*��{��p��4�(�Bփ�^l���c�hTU�I��7�Mf�{  ���s��|?D&��a��q|Fブm�?̭�B����h�<2�� :CQt�_�laľЬ
���&�e�CQ"R�����I�� R�A�7l��9�����\a �����>='�Pdr�Y� 7J-b	�UL�ʒ����;{+�n	o�|9��Z@��]r<0�� H��<�=Z�j]	yƪ�:���y�+	��Z��m��wށp2�vn:����#�C��T����b��{�x����{�,K@����'ٍ_��@�"�0���cL�8f	�h�i��o���Ty&��(��OuFr���pzw
�<�K�W�Me�M�Ȝ����,��a�ތY��}�IQ�:��筼n���z�0ǆ-�tzc2��v��p[�o�9ͼN�ŏ�ݛ��2�k�U����|��`O��6�~X��2��?�T��> ����,6����7;��y�3����p�5���Ppu��-_R*�ꢓ�Ϳ�WWnA%��� 㦻ړsl�~�XD� Ò����dcОn&
�Z��\%$�F�����\�j���$H�t`������C5����/���LC��7x,SZ]�a�v��\�gorF+�����p�-�fDZfԄ��慟u{p5�"i��%nc�K�U����6�gH[d;zݖH(�+�������B�(K�W�`�N�0�)JYƿ�~��@�W�ϥX�~m��M�HJ�io8�>;���MT���U��x��ʇ�έ���:���r"_�u���T4��eD�5�#��;R,�9H1MKJ�p�D�����+W��`71W���qQ�!���n��8���1֠H>�_�]��]�ڙ�n��8�=/���������_o���9;K�.���}N�P���UN|Oe�҇ݬTM�4H�i���7�I�5y�_X�;j�jo1Ud�ޥ���w��������w�4<I`O<eG��.�Y�*��B���#�j���N��غ�,�H��m�] ���(@���B���#�J�x��&&��.2����^�E)��U�4��Y����zf�V�4�/�e�h��5�ٯqԮ��X�+Af���Gٛ B�E�Hg,�Fa�5��}���,q���HÒ�5�&-�RB�I��A 3̏�e�� X������aҊ�]8g�a=Qդ��c'�%�l�͏��^�狙'�
�(c"���V��{�V��d�������m7�iuXcّ�Z
⒐q�n=W���!-�9uߡ� ��,|�>v
�>�BS	�~�i�BT^��n���?*~g�`�@h����x���MZ����2J��}�+C�������rh��)����-�N��4o:@)v��I~xm�.�iDU�"J7��_�d-�3���	΋5��T�eԮP-���(1.	�-O�:�U_β(�hn_�E�[9�/�ܹI��ܱ$���W�аh�Cu��=A��������~M0�K����>-�����8ԱM����zQ&@g
_�q�A�8E'���J��]�ݢ��@��\̦��+~��G���ZU��HA�sg� �c���O����{_I�5o{K���J�$��45�ڞ�����(����eUEZ��V;�BB�d��ǖױc3�bc��^�~��>�a9�R�d���Y]���Z�9݅�YF\�j�Ǜ�Š��ͤ�PCO�2�$L���;��y�������dQ�\�G�g�@��A���;��Yɨ[6v|EP���?1έ:�����5:K3S ������ƕ��IRyu�z���kuo�Oز.����EOk���q`C)j�l[ĳ�,�����UX�z'�p-�iB�1CB�v��}B�+un�+K���Q@��ߴ�#���\�v���`
�d}�6� ���4���l��j)�/������g��X��e���S��y�ޠ�:��ui�������d�i	�<q���O����[ϗ��)C�[�$�H���.�nW�`���`H�if=$a��L�Wzh�ѹ�
����S8�S����l^6�cQ��O�F���}��}�'[�Tn��06W��$��A���ZG��/���(�����=��ZH@!7����^��f�v~Fi'K�T�����1�:o�~Ԅ+!����@ln�8�|4���ņ�BqO�7~um^��6'^�1�}^��XX���=�챇����,��+���(&��l�d/nJp	B���;��&L����0$oaSZ�����B*��\ts��'l�2iX̳���ח���LF�GP�D�T���)RaƄ�q���Ф����,��0/5���yp�
�0�n��`a���$��j�J�Z��7��/`��cb��g~B!��y�����y��[-�5 ��	}�?h��x�j����5�	j~�e;j�!:�K���p�R?�����m�ZM�z����Z$z۝��R�z��5����gl�]��y��3#9���[�D_��暩����YE��|���K�s������f��� ![���Uݬn����s��	$��J6��C��.���8*ҕ�,���������g�W�"ko�2�Y3���V#�ճ>g� ��j��z��ʟ6t�`u��{L�-�$�ؒ
!	����h;��ZA�+��-�cl�E�gA��b��Y�\A�����Pg�J1K�c�[#6�~�C���"[�pc��K���� �6fA��K9��%�=O���. �{ ���vV�;lc�?ڍDX�9�k��*��ҳL*�5=�%�^�$Mȭ�LX���b��6쀻���+��#�z+ی-�\�>��!Խ7
��XU�,�)>����1ݽf5�숼�Ry/�g��M�"P��]K�&��ڭ)��oU��g>Wm�O�7d��%�[K#3xK����An�#��2Z߾�bv�͕�X;�F�T0rF�jDQ��!#����O=~��q�̃����	ȳ���ֈ��.L����ܐP��"in���Hb�Q�9����d�賂�o�}(�2ݨ\�y�@�'�:a�6��3��׮4���1�(<2tݹv:I��	�w(�0�����T0�".�����Ci����x�h�|5�88G3z���e��)Pu��K��xz�X5�4DT�J�A��� �E8�������S�M0�j�ͩ���q�MX��1M2Vܔ0��6����9��C�{�}�Қ���|������Q��I��l+��G4R×�z�������U��q(�^���\���y�K	�M�"�9�������Q����&3�^�qZm9�Gu%��'�������v؍~��<M�Ϟ��+ x���$�s��R^��ؠ��E�[׀�Aʥ�6��r�j����'�������?��}�
�r\�����[D��Nu����Շ-5�Т��y)jv�3�<�5su��"zUp�9��7W�P�Ą�������y�7��!v�Ԑy�Sx_t$�L��u1�>���]~�ˋ��������S�!�Bm⯍r�G�6���F��ϼxPsz8�@�Ug|z��4`aJՕ���~�<�dEb> �����r���~#"ǡ�>P'����h
�ܴ���,9J�
a�/J���ؠ�ނQ� Ѱ���8W��5'��dx�6��y3�w�Ш���Tf�e��C��Go�h����w��3�Q΅È�G����=������iP��x�9�[�NP"��B�mB��R�m�����D�s�hN7S�0����WJ��&���6���\� 6�5/� �Y ��o���o�+�T�;|�!O�o��#2$���=#v��tF�����?X��e�\�coHo�ey a�u�Ǉ�,�]��ƻ3�	/�v�8�	O��6K�_*z+��H΂C�TDV�Ovk.F�s
���|������ʈ�����U��(Th�s�a(�J�d��yY��0�[���Ph���Jx���6`VVA��F����p���&���ѯ�]ND%�Mʠ�ȣ|�G��x�;*{5x#>�yr����h�W�T��,b9�K�o����_�S"��ŀ�!��v��,h��Ї3pZV��!!PkԬk�4X�αd�ǝ}Ǡ'�v+?�D����L����R?J2J*�
�ل����}�Kh� ���Ǫ�-B���T#�\^��=�:f��JST*<�p�ձ�vG%�%�ͮ>B8D»���1I��)�T���Ǡmӭ��F��Z3�w�P��{=�����v�����xKW9@t�R,�.)�OC���b���5? �D*!�#������\�#�m��}T���H^d��Jb]���(p��E�5�	���R������hTh̀|��z�����:ՎB�v�m�ŧ��`�9G�b��4�0׺G^����(��_��;?/���$,�4�X&\a�N��m���.~��1O�=���뿺�W͑������6!CY��<q��`ӫ3~��x�C>��ʌ|���$������F9|`�v�� �z|�'�E�Ƣ4�=
,'��$;3��y'��?�u��D�u !�R���v�ʷH:K�4,����j���T�u���]��9GfkA�ض�B��h�Q��0�)K��2��y,~=��z�������n�o*Wq��S��Q688���0 ��k�e�
`Ą��h����3������y2ꆽsh���ʤ"�>4���<6�fE�PQ��f`���&� ��X��nf���a$�$���W�9<�M������q��>�`T^B�ޏO�bOݚ�g{9�G���hI�6�5g��+-���isX���s���H�������U\�"<�����:����vag[�|����e���󾏅z%����n���D���`�5��F9Bb�)��\J�1?Qnn��w����"�u� b�0���z��]i��,�w�;��_��a�& 0���b����	�o§����4!h%�7宔����o��0���[s� ��"]��'���tt��D5�Up���t��s��e�wH2r��8��NW�O��Z�x�ɾ��/�󳅊�&Ç�j�ę:_��G��Z�)Szh����3G�����7�;��ѼP��"�gGUے�D�ħ뮤S��8^K �q\��x[�I�_7��̑����4�S5fa�jn��a:��>�)h�QfA!O���p[�:U��.'B���J���P���1+r��g�H�2H���y�S�w�l}j����SQ��U�(r����3�{��HK�8�,�����7[o�m��o"ŵ�%Ŋ�t~���R���0�p�<�l�>ٮ�TA�5O>��r�^Ȟ�����EG%����E����G�v�i�Q��'Z�y���Ŗ���F,s����Lr���7��k�KS�w�c&���l�P�5�wȢ	��%�߀~�?���l����<��8������vhutb��X���d�O�M�!�!3���@�^���i��C��\(K��F�NF;`�ԓOQ�f
T_%e�ܴ���������F��%Υ_-2��� �T��M���Z°Q/-Z�#V^P�Ki��"�l}��3��I�t4M�~�ѕ��W��C"��Ɂ`��Ϗ<���/u��N.s858�Y`S���E������ �1Z㪦�h�K�l�Z��٩�1���3�I=6�����|2��=�D�b�?��K����N���g���0������O�f���V���a0��x5�ᣪg�K����������X�&�8u�h*b/b�<�X��҆%��^��)<���Ta�#�̍*��*�S!�|i��Ђ�K�kB�1_�Nr�uLI��6��;$'X�(� ���kB�˜���Ha�}�&#g�yc��7�H��(Ƣ�;�my�e1֍}�C`!��=,�t�qS��M--- �'���Y��ru
��65�(gt�v!vw��{�|�Dl�Pd���D�=��Ʋ���ol[+�[*�n8�k�f��@�Rbw7���j��/����fP�Gݎ�^-^q[
��O����T�}+��&_��7pn�����6�C���x�=�{�{���jF�M�8R5_N�>�ҙ��f\@@�����eLs��'Na&N7��3�ٽ���w�̏���R�$w��@n�=i���a�i4&��f���v�y��#݋���@Tc���z��0}+g�� �o�P��`���r,�/	�ۢ33��C�ɪ ���<]�<6UZ�~¡O6}�o��>�)l1kE/�ڴ};U�qü�]~��?�dJ�R��֭|�r-��R`||��a�ZS�a���,���拭$Aݿ� $��Ɵ��y�H�N,�؝-��ҡdp�Q#���e�#_�m#=�D�U�������m!X,|Rd��Zى�p�LLCHc�Ӓ��f$��%������%��tOw�<m�_(��#���}L�v�xn����4�S��۔|�7��(��~���_w_��_��씟�0�)�87~>�A��^�`4�����N0��^R��J��K��%�[�T%%_6ԫNZ]/��LZ�I���G8y�+`hy"hGH��=w����B^ڟ<L�u��"3����B��Lf�'�o8P�I���sib�����H�6|�R�ϸ5����b��ZBe�Lm~B�D��ΊU�/�y}���k�=�t��tUX(��c�3���E������m�K+�4��va]&*�`
�aQ�Ec�c�`�m�ߟr������k��A`o^���r�!�����N�&s�`��;=��y�s�B��������7@_K��Wu������ ��q�C���Z�b�tٓ��j�}�d��3.�e��$�cE����;eK�t�ꦏ���y�T�\:��ۖ���A���K֔�z��k�4R8M2z�X���;���Hl2v�:����G\B2����t��?h���K�+���R�{K�̓�̳_��B�3��PbfV;�w	+��F���D9+��X�*@����!YW����M�g�+�$?��mmZ7Շ,��t3:�!x�/�|q�4�)��H���S����<�q󌘗�����F�D�F����E纤g	L63;6
����X��%ă*�Kd�"{L�Q���F��pc"a�|_ʳ�{9�$��7/	,���D_'�z`��Ǿ����I|:��/�����s~�v�V3.
��0)��=˶������:���ݯ?%Ҵe?�M��*� <f��hf�א�A����z@�fn��)΢�6��Z��#ɌD�����nr���ѐ�e�m���)nфA����9����A1�5��������U�}��?/����GV��z���v��<	��f������T7���̑� 
|�~o�l�]r�^j��؏!�� �E?2��	"�q;��R0����>�C�	$�c���KQ�g��
��3���A�Q�p}�Q>\D���6�M�T�0�K7��wb�5�q����a)�$���Y��)� Hօ�(��X֌��e�?�|K�����y^�8��*�}C��A(���,e��ۄ
�5��U�_�4.D�d���B=����v1i��{�];g���u�W)�]>�yɫ������Z��t�EĘ��iW��U@��u�΋i�E�_�
�͜���	6p��\ꇈP�Ԋa����B&��,�(��d�G�)��֭�㝍i�뚷�<8�{{�K�P�-�).|�v���y�;�'���FTV�9�/���bƲq��t�e��6�U[X��?��P���\p�0tTv�O~S��2��Cs�dnv�F�.�GS���k0�*����U��̻yZ5�~������sp��=N��I��t�Q�a	�&�í	$�j����:��;�sP��"~�|J�Y���'���dź����P��IL���ԏf ',o�\0�I��k�Lq^nڠp@)o=sط�?��!H�!����gM��o�U�W�0��%��RPm�)�j�
����$߃!����A=XY�S�*}�_7�TR��d6��b��]&��Ӣͽ�]���Ȑrs�w�K̙����b��i֟\Ǐ%��[�V`d��/�Cن��J��W{1X�:)���Q��_4���{ln�\i���L�o����i��Sa3�)ٻ�jv˰�_iq͊9�r���/�j���C�ԠZ�X*�PĉF-�|�����^�=uu.���$�q�;��9���3X�����$4i��]kJ���E�Y_/S1��2�~% ����hK�_�)�'J�i=���V�2�~��U�ZB8'x�����%B�T�?zz�X���ةg�ej��|�~ o����X����5���upx�z��O�B�������!6��e�����6�u�{�5��J���2�w��;�?�o�2�n����xŞ�)�����#�0)K�Hg5S3��'T¸-��kԕ0�7��Bx��f��� >'���
�86E~Լ�xZ�n5�yؙ=%z|�p�����j������
�0[���a|3����������Ç�A�j�M�1����>�=1��啼z��!��;�a�*$�Bf�WS�BM���_�Ng
�˷�2�h�Aˆ��J���kǄ$6���^���?40a�5����8V9�.$��6�^�o'b�e���=}<]�G�ې�d��(����F
���+;��'Ef+�;�;u�����
�@$�)r�ق�����Q��	Q4��a|Vc�)�03M�c�v�AYǁ�c���Hj�T�q����U����C�;*��9�w&�1�W�9W�J���ig���aH�`[<���G�ٖ�cm���!��M5j���$/��sx���
���yD_�I�{k��e��S���,� ����Ʊ�/s_�,<c��C�tm�$'��^]��j=���K���u��n_����oŠV�:���:�Џ�݋�z���5��z=����8�%&\�g���O&UH���S-�d�����=�V5�µ��<�Hs���`���ׇ���<ۇe�v����9ɳʗmc����m��v��H�h��j�����g��^
�I�E��DT	��"�(�3�lsV,\.�Q,��mʑO�P���V3��4ÎB��Z��<��_5Y���y�g�9T�u/��~���Z���aR*Hz��&<�0��~�NX�q�;��Qz�#1���4}'��𵝖�o��+���IJ�	�Z�3p��o�@Y��Iz0M^g;	e� ����z@G�J0#BBf�'!�1+����6du��/��:d�lf�g&,����I劦%q�XMa	�e��@����ꪺB| ��d;Ƕ�6������ ��5��{(p��� <a�2Qp�Yv�X���J�iPt��[�8�e��A+.E����
q����<i;����G5�}cn���t	�e��>ᜣ���c\<0��Ӽ��q������@������ѰۋaEc��X�%}�Fg�(���UWZ�H�����64�Qhc�V��~�oˤ�}1�6���$�/�4��@e�h�j��gc�9�BK��w�G����[#��q �?����VS΍���WH��߭08(b�.�|�r6x��(�%�(����a�#K�w;�W���<��Et�|gWkX��+ �E�Ұ�o~����{�똶v����X���rg{�RKqW�.�[�5����1&�)���#;��詘c�>ˣ�F[m�]��`�~�
DO&�*u�5;;�bsX̂�B]��Kh��# �h��@���^p�2鹚�t�=v3p|�D�y��~bpf�3|&�*[�SFh�ʱk�ɼm�`:s���ͅ��aM׮�����/�w���]u�S��r`�Z��"ѹ�Ɖ�:��$���	�qQ(�`y�z������Mqz�4�=�@�}�p\��o���H��I����cF�̋��]c�@Oix������:4+�!�cz'�+�c�Ht��}�uE��j�q6GΒ(m�Jy`��D��>@UB�<�����%
풹��R�ɥӠ1�|Og�_��eqk9>��K�?��|+��_�L[!{��	�92������[W��z�b�l]�ލ~�%�v�H�klZ��K2Dܛ�뀒�JRLF�B��e���-���{�g�jee�O�#�MQ��(o�X��p;x�I��d�qpQ�F��z��{I�n�|�"�+�����2�[��Q���!..�N�����k���`�/��V]�c��������*��瞊?A}?t��л7e�G~F7��>X�t��*X�>
�* �9I,�7ӱ���M��׵G�ՇSE�&��%&=\�BC�߬�Me7zFP
fy{��}�xzWaX�uR�p��� �ޝ��V��K<���K;% ���q$z���<��h�J�� ���#��0q�1B���}�w�t��w3��c�@�r���Z����G^T��y�Xj�̈́۝���d�B��L��� W�������CN�~'\E��8Ȱ��*h�:F,/�m��0�ފ2��� T��Ue^��2�q�>L��	l?Y��E�N6�Uu6/��4�(]�
3�ͱ�pW���6�6T����f��%��Ɩ�_��|����V(��h�F�E E��Z�0��y�v���fE�-:ʴ��c�<B2ł��_��
���>�}btZ�!ɖ�\p�|P�wo��W��ɴ1��Q7��)�r��>~
2��wLj�������|o'����s��fd��z�K�r���b��#�5t��Lf�g��8=B�cf��Sj[<��穚��7i�/�/k�m��,����l�yl��6~����M�eqk�W���"��ݭD�#�rH���A��9C�}�����S�s��rQ���[մh�G�����[�;���R�_�����>�)� ��k�1�,�d}J�W7����r<�G��K�X��%$N:2���'����K�B��R����ŀ7�� �t���߬9�>7ԧV�i:�I���n��溓����Tgst�*(7U&_5O���D��w��weE�N@���%���U�L��(��j�-̊�*�Az���lnq�C๓���D������)�m`��Ҭ�W�QS�Qe�����i�����^�TON^1.@��C��������6�����VlD��T���/�XQH����mj"�+�a�Ӈm(�9����T�KE���
`���H�}㱓H�`i�L])o��z�E���f�K�?�6�̪�����o|r�S��&����Tm��}]@��wy9+4''�O�[I��WG�=t�0C��`ƅ�H���R��]�t�W�@� �Z�����U�?4���1:�*?$�1��Ԡ^����i��9P�?��k�R#�����M��A��\���,�q��ׂS
$��T��C)*����N{z�t���S�iBX�A�t$�*1��Bu�����dA]���d�5Coݓ��W�X~>����j�_#�"�_���%��C�-O��S��v�ծh%K�F��L������f+�>:�p ����4j�T�垏.b��E�NbwQK[�\�J#��c�䬊�lTOU��X0�}B�M&67�D+H��D�+�|~4�!땇��e�UǱ�e]�ز-=Ҽ*�z�rnz�>�����Ω �.Q�Q�K�Ƴ�)vJK��\: �%��O;��o��opL��ߕ���b��؜Z��l���p�Oƪi�ʽ��"��� ���	��̜����w�Ύ�a�63@D-�v>D@�R��2L�{P��Tbs̮p�A���S�&ہ7��)x�N+:��/��!�L�o��?�;b4�ߑ��^W'����� �l�/���̫��\����l.m�U D#^���g:#��F.�L�5Vd!�缘Ȏ�|�1�4� ^D~1?�f<�H�Z��Gz����F0ᱢ-����G�/�^��9¼_F��Bэ:N�;��F&l���֟|���A�xM��x�=��N�X������@S���0w�PKǼ�)�Ǿ��FP��2޾\�[nxP#}2�RW��K��f�l���qcK*����4T��t�?����'�Lb�x�/�Dgje39�[�՟#Z�~S)�Lx�dgɺ4���榶ܤ�O����L����k:��`}1=�J*C�F�j@R]�j���Ϥu<k�Ÿ��M��U����^�fo6�}�+��*�iѝ�rɁ۫Sn�[HM�3�뀦�-\l�&������Ep����H��lT�[�X�߷��UdʙO5J��d��e��yS]�^[hzZ�(F	 ��k�g�X�"�d��E�F�����+���������-ņ�:�ahϊ���5kxq�O������A�o���Kh-+#���a�>�w���B�\���6�h�m��Ȱ�Rl��@��#~�v+�T����>��n��T�K��^[������y�F=��~@�� 3.m�g�������./��$�|��BU86)�9�0�U;�!�{�Q�!7�Ya%m�qJ��� �Ŭd2� 2i�q�E���g�S�b��Ej�3U�I"��}���V$����j���2Gzf�����y*�fQ)�lhʻ0��rEK1�'�W���eh⺄���H��������p��%�9ϯ䧗�BO����G��:�H����-�Xl�eGpq��:]j���@莉���&�Ɯ)�+���	���\��mXd��)��Dz�8{,m	���\0!��F��8���M@U�G�.C6ʻ�4�������"���)RNb�]�x���	e�d����
v��Pz�X� ^�]đ#��l	�T��Wx	6;٭O�� �Mg�\iNh��������r�	���_J��-[��O4�fJ;���^T��0�{�L;�z0�ڂ�G�Z`����e�+Z)-Yî����
��O���LӅ��X�ވ� TI�HU�o�����Ro�c��h�0���Vai���\uCWL����N�ޚ�05�ؖ��ꉿ���bĎN(13a�������O�?�
�D���(�O�"��뒈�t�� H�� ��"Kr}T�'�#nX;��K�,+>�빩Le�c�����}!�/���P��
�������VZ�@��J�;�U���R �n�R�FK肳)��I�D���'&��z� �J�*���@i�Y�:�?=kȭC��YĈ��2ᐰ���PD$8Z�-e�N@~�LAX�9�-��B��p�!�-��cP���6@�������{Z�N$�G�;��A`+��2k��$@�&�?�8Z$�����CϦQϗlv�u�H"��XSk)��i�Zh�y�%�8���I�$,�&�$��6�'*�1�n���J������SZ�1ؾA��r�N�Ā��It�,3D�O��iW�P0�f7�ь�)a3�^� �����l'�)K�Ǽsf�Q�t�B��{�F���A�F�GJ��w���W&�����vZv�Yu�wQ��(��)�o����a_���.���#��)0H�ݡ-~��SS�3	Z��_+��� ����߫#ޗu����j1,;�~��>���'��'G�I�bhzY4_�D�������"���,�jh�e2��'	�qm���X]���������IZ��A�݋�B�#��\;`�У,�A��$�R�f��NB����+ufZ<�K��o<݃Hm2��3��qM���[��񑜍�O���H�?�pp�!�2�#�>�N�]!"*2��*�]�*����`���d�!�Ȏ俀&��㭧�d�i��w�(��0'%�цzf�q&;)�*zg��e�>�`��G����z�E���o-���v������"�"0��{��5�@N��~�8n�n�d�;I��H��S�3Mt0c=��� ������)��|���Zf���!�ø5a+���`U�n��м*��0�gRg�Y���w��W���ӟ�W�kA�9ҘR��� 	~�Uͧ$�b(�Q�N픨9^�$O&	
���q$UT�1�'{�lR�ѿ��\�N���})�����x��F�B��6��7P,� ��4�u���R��CE�h m��"
2J� \�rE�os�\��n���H��P��-���Ou;��)�M��2^�V<�|��IL�(�浂�h0��/_��s�´劢�ƍ Ƙ�\��D��)_A34�$���MQN��G\�N@/��̽�ӽ*�J�9r��îƤjZW�jAv�ī��a�\yT��u{ae���n�����˼r�;a��Y�c��.ckz"'.� �H�p�p`�gMGSG��:��p�I���~�xA�w�{wR����V�T"s(&������~KS���
�_~�r�5���s���-\Ư�p`���<$�U���$M���������(�;Rʌ%y�!�hU��w��w�m�<j�<f�P�5�Tz������KN�[QҁqJ_z;q��nAUI�����᧠nl���͡b���S̔Gl)�����8zf�����ķ<9H�K��e�v":�G�$@��Eɡ�\�B�8_sg��~���)Fq��/�kH3]B��#ZAv_�i��f`���@x�H��E�����8���O�����?�`-%q��S��`,~áX����q�z_W5��v��qj3@�.��89�W�r�I}gw4�C��/�X��#���!5yA�?43�HG�u���1��	��h�ƃ���6���
4���
���q��AӺ7Ŏ<Y�]��;�Gw[DS�\��Z��Y�ϣf�K���pڐ�s�"�q�N_���*��ǡO66�˜���K��<~7�@HJa��o��~Iá�IS���y��h��5�I1��ި�c�4c)�T��G���ot�E�DωU�*pBU7iP 
	�)!�|CU�;�E\�A��h�Q�#ޯ���R�0�z���[p�=H�ˢ(����&(�7��b��<�'�؊���˽���ұ� ��N1�z��h�����]S��m��ժӉghsd��=3�,74�+g=+��	�����u�yl��5N���� ���;�T%�5/����1w+��a����3�M漫u�Q�ށ�F���uz�'O��A&V6��D^I%��E�I�����a1��K�
���m��z$,�ȿ0���˄�i-���u�Ox2Fۃ!��Lk5;s�����b^<l�"̩Š��C-c�٫�^D���^\'�m3��*��f�1� �@'"I����J-܀}*L*H�U:�|���(�,��Q.�H��$t��ҡ���5��y\�VRc.�(����NT�8dr�Q.>��	�"���k�������"G,G_�?C�'|�	��[cR�5|���wӟU�8�+ڧE	�\��.ٸ��2�r��-���_ɱZ�dd��V��t��L+{��u���FMR���~�0C��g�D8i뮲�o�O"�1׏��~��I)k}�� O^��}�@�n)>��1y�qk��>�r�|zIj�Jm�V�Q��ξ�J��N��0����-�ת���������n��~���i���}f���㈅��yi]o7F��#�_M��R:��ڋ����mA��ؒ��o������h�%4mN��䳏�ْO�\f�Ne0k�,���Xda��+s17-� e���8�M��l�34[�'=�툅 ������d�a��r�sl%ԗ]��P&��k�9�����W��C�U���h����w:;�q"���V��I�4bFo�|�L�I�n����P����MA�b�e����<���s������؆�v�K:��S��*� �-A#a������Q�Iv;����EHn!J�/���SX���b�HG/�.-=J���K�V�>�:vg6 �fv�����C�+J'�ύ"�+��p���ݬ�]��l��~_����%� F�����a��?��fS�Bl�B���q�a�qR�,K�����o�#׈�^�.&��o��N�
W�"��K���P�K�g���#��٫];�u��3ؼ$�5�3mr���������|��'�Vb�&�PS�A������� ?���������w��t��8��<%E�ly���'eD�b:���O�9�Ѫy.���h������SI�a.5*6���H<:=��	��v�՞�9}A�e1��r��D0�*ytk���t�`�3I�Q4�7�g��F�r$6��<CI �l�u2�s�0Qj~X�Ԡ�^*�������֩����EV��X�c�,
�
h�EA�<�,��k��{�H���D��r+{��,#�K��Z��B���8	�.����^:����mp�o«N�̡%!�ҿ��S�H�/q��*��`�-�ˈxÜ��O�ܤ�0A�����}��{��U9"[�����8("p�n#+Tnxe�[D5&c��瑮����I?&�5	$[���wX�%����Yu��\��������߂'0S��{����iߡ�tI$�(�H8��>;�lr�3]�$�Ua���%Q���ӅLv�����OV9EFj,���m�N�;�0��<���R��0r|sJ��z��#�}i������.;1��M፲�E�;�ZK�&W9S~$�=��<�7�ϋG@��i1��*V���SBnR���<t�J\��"L:CL��Js�ʏ� %������5�	����5;7A�:-�[��h+��oy �yje�Z� �}��rv�N3!=��l��ض���*@��W�4�jǸ�k�QW> ���g�{x	<��G"���c	��ԡ��}��gi�-u�2yM
|J�J䵤�q���u���|��8��'A�h�VC�+4�����n ��]�t��؛��.����������鲪P�~CϮH�b�X�3����=�ٖ��~��V���@]Y*�6��\�P^y�)�����4����MF�%M�?�C�u�䕭�YTn�u��$�`���~�5Y0�x|_Ŏ�O�dJ�U!u��<MTo���}qƋ�.��]ۜ5��͢.;~�SO�~��Z�\	�9��ƍ|B�,G�#�b�^K�պU_ ������KS�&	  ��XzU�)|��쐾q#E19��h:�u��n�E��@�B�CC˒�h�D�G����GOC��^q�+�D:��x겲�E�y���c	ta���)g��+[�M��ɓ��?��|������ua��λ�r_`�ͬ]�>��i#��������e����)��Mu,m���k��"�
��(I������S%M��r�)���訑��{>�w3s/h܈(-K��w�3'pfM��֒�/P���C9� 2wq�ޠr!�m����Ӏ������*w��xH��ו��dA�!�h��K��@o�����Fg�m.<qk�o�\ۂd����:���c��O��:�O/x.:��?C��M*�Bs���m��r�L���Tb�fD2�~u��w��O���TD'�b[j�O�@`�۳)#�&��C���v␂�Ϣ1)p�������yX'�ạ�����u�'�No��5���3�t.�3k&y��낆Ta�B>f_�D�p~�0�	5j�Y��G����ڊ��i��L��u��N~�����1q]%В�G�3��1�<,mP��)�rg1+8��Se$�(Xܱ����+%�[|f�l2�jy9��.�~(Ⱦ�L�,c�څ��ĕ�!ݷhf
T��ibc��7�i������:�is;u:k�]aH�'�"���\�GV�=>I���>�����֨!
@�]k�{	�}4��!D�g"����1x-�]=�iʅCP��)!N�3Y׷�]����s�-�<��LB>h�kL�5�����"#�+^��Mn�.�&����O�}`��D /�;�ɏf(ݿȶї!�.إQҌ^G2"��m�ī+��]{����Ś���^3��[?擹k8ā<�^�;����ܧxc6�'UF�������H|*�M�*92?Wp§/�"��X;@�Aa�mp����b��H��A ��%��\���;���錡l�Hz�Ya��Q�s(�;t@I�-��k :l�3F!2�<���|�0�}6-{������;Ӽ᫹l9����O��5��IS�	f��*�k�'e��l�>��bx�T#gO�&�ށA 6n�G���mN�_���d�Å/q^F�R{8;�iׄZ
G�<��#��
�W� ?�����逆ϋ���;�Ɇh�i�e�ǬJ�Hg�r"�L������ª�c(I]! u%�����P��}���kԈ��I��Z �DUͬ.w~<�W�7M���?�Q	`��!}��=�/����g�b��VpBdEE�T��t)ؤS�/ї���Ң�Ьت��? ���̢����˵��Y���"�ˌCЧ�����޿�/����(��G�1�W'(m��3��K����|�#,W�^�TYh�K�j��	Q��!��F���0N��Y�s:��͘�ͫ�u]:�&��=�3g��������o�� r�Ω�<|:���8����F�/ڣ؁o�k�������y��=�����k�UE����O\a����#|�+ߗ�r�Q����1���s)���˝{���-{��жMF� ����w���Q87�
4���!�y6_�wd��~<��Q��h�т�)l�\s���L��n��p��p�w�O~=�Um�#��B��3	���v�ͮ<�"�P۵���f��M��.�0(X��6�z�e�^��W+^tN�oxu*�2�4{���M�`��8��}���Q���IjRa4��ЬK�N��:>�eH爑�����&IG�1W(�!21	�BӁh�ѐ�̌�۸٣�� ���FB7���P�W�����-���uEf����=�n���z*:i�~F�`�v#	t8���Yr�/��8O�k`��f%xΡE�u�f���&\���}�6�Yd8�$����޺��p�h_6+xX� �[���2߁�,U�V=�h��3��x�Ÿf�OR��nCK�ޖ�rk�Yk���s�/�|��,;ԥ����9~h�>$�.e7���\��3�X&���
�Aw��)�j��4y������-���"�r��QXQT7�r3.�Dǃ�>���VJ<��9I��'7-��D��ۃJ�E�s�M��P�f# ��+3)��S����n��##i���������u�:�G#��, ��T����B��K|PU��O#��I ��k��,��z�Z���n��DC����Mw�]��U�Ym�5`�+j��M��J��5��+���L[�4n���#�
}��3�_o舱m,)��Z��Οx]s?
��Ʃ��J�5�U^��Ő#rd��\�tAu�N45d;��o��j� b���Ca�S�L�x����[慰���7��J��on%W��Ξ���IB_�,dJ�M{�W�����vu���'���-���A�=����-�se�H�W?�"n�^;��z��]��e�&���-SՁ-,�$�ƚX2jD[�TwH�i|+R �ǞFΏ؂�#��b���4I`������{g����̌Z��]�dX7��B�Hp�)�F��9��;I�o��K��ˉԮx�" �g�{/�M��`W���Ҥ��/(aέ��m(�k�7���ȅ���\DQ�3���)p�Y䑇�J0\��S0:5 +�īT�䶡����T*9���ߌ��A�,���,.'��:�P�b��5��/`��%�6���%F�UC�ϥ��ydF��R�T�kP��U������<R��DF���o{���<��n(�.H�K}�����6��d�d��Õ�(��� ��:*`��q��q�M1�����M57=!g�;������ozp��r6*�<��k(�J|�������,
b&ݛ
����˳,L<���4�ȧ��tqs?���l!��ۃ��Y-�H�2#f8��wΟCne���~��l�����T�lq=���Z6Q��H�+<�;X�^��S�:Ix�uh`P,	���	'Q���D��=f���(Bz-L)9�";6,ϺW{E;��h�4��\���)�w�YH�S��q�+�i|m3[���"5"�P	��4�;��,�W�a� �ᵒqh���"	K���͹��[��|����o\O���U̬g���4�˧ղ�������-��M0��mj�����8X�~ނ��'��A�v���b������O1	ST��,E�>|��qFM��x�<c���Z�
�W��G�q�yₜG�R��x�0��"�yH��?�<�\��Z4Z�(��^�4�tZ��.�g��p�)HQ=���B�!�U�n1T���f@'���;,�y�-^�dS/��I�G��]�F e������^�����d'È�%���w�|	xG����
H��������� ��:W�mͱ~�a�~�N~�j���txv��$����<��ʧכ�w�X��>�!º������T-/�Jr�� I*�Q�o�cǍ�5��b�ٙK�i�s�����&a*��棏c?*���M�NHٷ�ث���^y0wc½a����|��u��΅b)��o�9Ŗ���e��'�d��
(X޻:ۛ��XMê�*�?��S>*��P�k]�G=x6[`s3ӸZ[��G��9�@���ߡ�u��[���i	�?�r�wK�Z����:�=_kr��{�C� ����/)<�i�)_��g��;��`a�W���ZUAR�ȏ<�iKn����C��ê/@T��vjoj~�f�8��@�U�3c#N�����6A-�ZH٣G���m@����%@�xW�L��h"���#�B��lP�=>�-��Ǻr%a��
Ne�~l�s5��]�!���E�RxgK.}鿭.����{�Kcv�=
<�}��������4���sI��Gc��%(����Ƕ}7��Y��n��1�O=�؍}n?�՚�_ŹK籊�-ʄ[��K�U���5*pNݰ��7-նHI�c?���f���x��ƹ��p�	���b3�8I�Í��qMAˑ��!]�yֵ1{ 	R@�RD���`� R�K?�T�;G^��#�m��Prՙ���Nd@3���&���խ*�f�5��=&mi��]��t䬼ж��	
�	��V����Xx�'ՙ,�I]d��팤�M~�7k�B}E�y����E_�ֱ�nX��߀��j��]��O<,2fS�*�Y�`a.s�J�G '����F���襍'��pȥ�$=� �����W�'���bya�T7Is�<���`pD�C�e��V-����;B��n����Z4�	E���"'���1B��P�Քf�+�Gd�u%����<[��<E�X#��� �ʿ\?d]�Ð�)���o-r{�{ٰ&�d�_������o|��7ɪr}l�7������b�[�l��,���UkwK�,9]Ù?URu�Ol�"��4^�2`���m��2���XU��w@�۱7� |oSYi��2�Ro��@�eKṕ�w�&�29�_0PX�HX^�Xx@��Y�4�P�F|&M�?B�}�-_41If!�:�j]n�1���0�D��I��@�����F}�ݛ�}�h�9�e9����<�f������
ʖ/8�*�J�Z���	'���(��T �kO�,���A�'�Is���+�#y�dH�Bg��+������|,��^-K^�+2IÍ��o~a��Y��C2�����W:/)!���s<�s�t̥e�����<�M����������J�����/�Ԫ���a��r0���>�����Y��U����9����\����H`��2ͤ��YWx\�nY�e*�F�N��)k]Y�zpL��2zU�{Q/�z��^r<�F.e�i��L�U���PR�c�F�3�0��;��,�� �qg�H�*@����T�v�mL�1s�g��-3t����c��x���mȡ]���p����G���H�5|�.Z�y��SI�R��a��~&��W��-ߠ��Lč'��\+zq9qG��Ym���HFO���Y!X�klDnR��nQ�5��t��z�d[�.��;�.�x�3�u�Ͳ�HȴL���V�mC�W��V��rAȭ2��DF��'��ձ��p��W� ��f ��S�\!��l-��h^�U?�؏�¼�#�Lh�' �mVb��;�+mF�Y�
��=�W>�=��u��L���G聃�z��
]�� �E��W�|P��;�%<�(��W3�D��8Pp�y�ym5R��uZ�?A�?�xp��!DJ���Q�u�3�T<�PaI����u����h*��;�"1�:�s��_�f���� ���$?ΟvLMBkm�WȄb����T�G�|W������	]���< u�3��4j��>2z���:�Cg�K�Ef"�L��Ң�9��\U�9�~�1�f���p��Q7of9�:��0��Ϩ��n������K�4O��)(�+��!8�Z��&B�� J��^;��lrAը����dJkv5d{M3��͟bٔX-������N�ʇhn�,+�ZP�?�m3�M~�7L����]S-x!�b����rH��m(�[_4�ԩ@�6��9���b�-[+�$�T�������Q�=aRrj�Hy�T����1�Ÿy�o��RybN����k����;� t��[�wZ�w��^J�9�Y�]%�*���-u�h�k,��=sr.��RpجM�
�{�R@&��k�����y�N�3�~p���U_���������}�w�V�Pח���b��ʃڔ_�qi�#�^��>Xw�"�Uհv�^l�\+�^Qö&H�,���KrL��s0��ɀ�B>��Z�;ɟi%rD�����|hZ3@�$��:V@n'����@c�G�]�틢��Z�,w`.dT�]�6���M�T�xXg� ���5�G��zM��O�A$���I?�c�RU�{�^�p����?A���J�T�5�Bɰ����[a�^����]���b�xޝ��n�/{�y݊7�h����13���Zl�&�]�Ύ\�z^k�K��^q�q��|��r�}�eq̷O»�}�E0k$�0V���|'���qG��qd��l�E�D���xE,~��o�Hꇹ��ŒR籶5�1%ўi��&���|ӳ�R��9n��(�3n{�s���.�E/�O�#�7��ɞ7E����ഊu.=�n�s��APZ�^4��-#h`�Ik`�M�"R���]�q��ۀA��s�z;�m3s)Q4�",Bl޾1p<5�Lf��[T>��Ftx�ρ!�f����tz���4d��vU�� ���%¼6;�������=4{<��)$�ٮ��X5�b$}&�M����9�k~+��e�Q��%B�	5�ty�͕�c�2]���1��宷K�� w���䌟7�-4��h{4�� oЗS(-Dłw��7t��M�I���A�9p�t�;3 D�wx�͇������������f�Q&�-�_��]]}����&�)'�+���t�Q�4V;j��#��;��Tc��S�,~|U��b����Z��)°��U'oEغ�C"r���l����ל
���8��UN�~ߍ���TD�����qP�:	���J-��xP�I��^"����L;�T�>�7��E��Wj���Ѽ�F��Y#�a��T8 O,���EO������{��P�����͟S���K��pDDb()�5��"�B��6& K��K�Jh�h6����O�(0����x��.)6iQ�������[�٘��C&_���� �P�0E���/��x\I�b�C{�Zxx�e5���a1_\*e��>���f�T�����ņ87����/���<�I�lex[���Tp��h����|i����H��sL�gu�s����]!� �O������>���$����2�M������.bK=2Ld�&/$�Ͷ�+��q�	���B�N��L��(��o��v�R��.l��! F�~F��,��1��h�g R	?����V%�����uN&�q�'a_l�3��$��k�gCR�%�L�����1�Ϙ`L.�L�Cc�
ź
U+�<2o�C,��vʛ�s���A�b>��@/b��"ɖ�T�^W������*}ȩ�v�	�IT��r�o�
���
�W��m��Wp�2{E��k��c7c
��� �J����3Z�x6������G��������C����m�%˫��!�@�Y���\��<��{)L��ˉ�cv�|��x�l��>��t���"��w�T��a���P����ŗ�����\�ؽ��4���A��d�z�9dt�P����1-d�g(ML�}R��ؐ@$�K�#��s��EpEn��.�����]��Xߓh�Ed�d
o�B�BK���׶�T�� Y;��
v�v�0{!ؾ1TE��|X2R䮾=���$Q"Zb*�O�*.�\(c������y����@_� �v���X:r��$_҄��|M�Քc��+�n��b��E:	6K���%i,����rΔ_��(0a���%�D1l��	���9Y�%SO3���-��Q߅]���%��KYSr6l����L�<�O
=���E"�xrSLq�%A�U�Cr�-Y��íUEv$<�r�範"q��K� ��ݮQzF~�Ɖ�Й~�G!�wuQ��u9#�i<뷦���������D?D�������%Qd�������-���O���/��*{�cC�s�O5*�]��>8#ػ0얨%*��?�X*D�b�C��7�1Uj�(�S�JTn�����t���-�&ߐ^ݪN9g�
Y�TCV�b��{���Q%X"% =^9��^0�ޞ���3�h]������̴ߕ܉�&D��9�G�ݰ�?�r�6,��f��b8����d9���^Ɓ8X���Fz�)H��sǖ.�'��mo/ɪ���n�܁d'ǀH*�)���U>L�E�Ր��R]��[���R�}w�rn��`kE��!�Hm���m:���uݪ�`q����\/��0\� {��)��m'4D�}6q��EHFӭڔb�?达�5-ybp���T{��VdK��>?gߴ�8�K������/�����q�P�],à�rg�gk���-�`UB�z��j��>|σ�������^
��M�{cu��\���f���ה����:��u���>	شZ^��c��o�������c�g��m��x��K��vw+�'=r��~��]:�W� ��d�
d��,�)x1�vYJctZB9�:}˝��kךXyW~���K��~ �Az�PI���6�u�v�>���d ��U���+R��Ṷ��i�����-Rܛ/+T^�ӵ��;�������	��pM.j2�DlN��aI�&��%�K��׾���5a��9I�[	���{�l񏚛�I�=ᵡ��G�Gd�1�R�l������GZ���ͪN��.� �z������zi���傼PU]���k��{Z��_�>fw�TQ��M$;� 8���*3mOo�� T��aO��Q�� ئt�|_�x�� .�w��o�#��4�E�,��J����a�C{Wc�lȀhw��2�~r�Z��M�S�r�Y��XR�)���^�g".#��=Ww�YUMsR�1L6u3_#�h��W��`놫u8�� _^v�nM����)�/oka?��/(&�y�Z�=��W�V.����+�(®f�����a_Tc�C(���Q�q.�Z��U�:*�?���������̒�lh4Y�=r=I�Ph'x�=��G��Z����-0���'AL1��нu��(h���x&�]�����!�<��\$F�e�+3����[��I�γ���r&��KYD�w��?א�p� �)���td��(��޳r�_WIFf��3Ih�>�����1�(#/r���+��ǴF�^�>PU0�����o�A^~�}�/6f�.4���F�4�3�ҽ�A��*b����0������Gn	4�&a=ڢ���6��L�,�k(u#<�rb��*����������Y�A(���F�n�؋�õ��ob�4�>�t�*�"�<mP_
��g*ކI�3��Z@��s���В�Sf�-!ܥ�VB�#����7�t��D.�5����Y�ϖZ�B/�fiw�<���ꯗ�	�e'jwMV��5�P����ī�����q��_�r�!�j1����U��1뉵_x���$���$�c�F�͇�A�2�j3����.�FL��U/��"tu5�8�i�+rz��m��G���-d �
T���,t���nR��%�[^�����S��+G�����0m]�=מ��19<�~|�hf�,N�r@?W*	넠�2NY���fS�<�ގ�`-V�@�͸;_U`B�<�ޕցZ��yT�����%ŏZ��֕�q��Q���M��ݝ�#L�.+�1�w�����������y��i!���������_$��5d�}*
�[A��#�E_��M^�Q�N��m��{�?��t���Q�qx1哺v�D8�=�7�{f��.=��V��4�,;`k�S��>�5��Ԙf�.<�� �`�#m�AHF�7�9³7ҿ����{%'�N��:Ǥ8ٞ,+K$��,c��}Y����H�#��^|,��I�DC@h ��rx��\IU���]2jQ<~�,G\/8
+|vD�:Dk�F3�9��	K�J�(�e!�|dl�b����84��X�].��m_�F���	z߂v#�^�ͷ��6!�ݮ(�tG�����vh���R,Q�������r}�n�3�_A�/ò��`�qS�b�F���I��7��S��g��uU�-���4C[�������2͙���&PSԄ���\Ȯ3=Yn��'=^�j�3n��}>���Zȿԣ��b����EӁ����ȣ vD;�0�
T������¾d���#r����A��ɋ��\���h�&ո�?�U*g���i�1��%�����_h�����zfF�ΞS������Y�F�Jݥ(��*)[�2���u4��ؗl�S�ί������!`��c�������7�2L�
�vwC6���@vD!A��J]�a��E1�e%K�B}4z����i�6�ս������]�����i���=@(� ��J ]j	������A�V�b���Ǩ�S,i����8�L�YIdWo+Ors��Fs����H�����r!1�W��mr!$]�KE@X�Z�B]u��_�O8k�`S2*���5��CA t���S08�OgxP�(k�e��B�2�A�9�䔍'�oۖv�=��@�e/Py���Sno3u��X���� ����i��I�\,(�c q�mj�A7��7�l�m �����¶�9Yg��|�E�$YV�=��V�g.��o�^�a�ϊ"����ȇ�l�������#Bd'l��0Κ�D��v�����E��i�d�w�w��hC7��V&/,���#�I���Q��o�.����<�+���>�O����-���٬E�ϒ0�f�շ��|q� [�OJV�������Ϸ�E3"�v�z������:a���H;.�QA�I���nu�����̃���<璵�Q���]qs�¤:�A��l���p����?T�s��-jX����4��c-�ѳ� v�z+�*�3�n��^1B��ݸ�O}d�EޔTd2=�M�q|�K�!�S��7�,��Y��u䎝�i�� �zxc7��4�M�I���
+1� �ҚnY�O��S�� !+?�$7�S7���
9��G7?C�>�ƙ�Ս��:&�o�� F����˜��]�4�X<d���l���}	�� �(�e?r�͍�"�d��uۮ�r$�'o�Fq��7ؕ��
��1�s�y ⹌k:���B#�|ڢ�'KN}BTb��u�'�d���ٱ`��H�>p]�k�/�=.=��ul�&�]�Oĭŉ
��2n���	�c�suE8��/��n�2�:ݓN�O�d�?3~�2٬G��o[���OE}��im�W���{g!lKP��$�v2�jx{!��KXW��~��Q���'E�D*��Y���$�_징R� 撉i��1�pO��!�\�H��D���a
 �μ̒��a<��Sx��o���3�0�^�J�o�B6��&�}nA�>�\�}2�RS��Rl(<�*F�t �u�YoD��d?���T�vd����gSa��@�2r���
N�������"���������{b��C>��C��]��r�Fj��;�����_֬�:���I�y���������`��@u��}�JH�ZlN�e�Sx�"���+���X�PM$_`+ �o?0r� �r�rI��"��EdQ��"�hS�e�\ɉy�F��_�@};P��V�On�P�����R�gP]1@�t�4�v�Y��+��%��27� t���T�$b8�k��IE�E��@	�u�T� |��?�g� ��9vK5��ԣ }h�.>�B�i��
1n��a�X���j)�@����B����߈5����T���oa�]Ę		�b%K�� ��8�dp2���{0���3 -�����>c�N�MÿI�M�����8(eE+2e�D��5�\\^ T���*��M0?�D�gۣj�~c(�6C	���2	ؘ�c� Cpջ��L.��L�{r�%���0�uNd�R�Cˇ.�F���	�-�ʲ<�\���(4��{���ݛW��y���V�wJ{��'DC�FB��mU�X�<Q��I��mKZ]��3A��U>�Z�h~��%A���f��VH�![?f=$��*4�<�(̓������|��H�T�w�B7�}Y�N�����J����m9��|��!�ZU����X�2E�pqG�f@�?@ȺË�u��{��n���L�ʺj�I%�p�Uy[ :�v���߾�������(Y*��-��Gj���i':���]�|�8O�$S�7�����u��%d�&�]W�,����k����TW�>rS�n�b�Q�?���[�|$��g҅�fRYЗ��M�D�A����1�I����逸6ưb�#���$D'wFpf�iTـۘ`724,vW^�CSP���Ez^_�����l%����~�.P�K�![�Qd��EQw�}@�d{*+��k1˿L]Lc,��| @)�����3|28�:�7$>^!8'����=ےz!�>
���,�1��1�)��$��c6U$O\�*&��D�1�v�O�)~��^�w�!��Q����� ��ľ�����b�y�iE�Б�$i��}@��Um��;;��K��x�^`�ŗ�%�:���=0��a�(X�c�\���%���]��?�
�z��`.�bfg�%Pz��-��a�v�9}.;ï2h�<Yn�L������Y3��v�=G���6��SY���Ee��P�r��p��&� �{�?[����s��9s���?9%�K��7x-��)`���Kl��ҁ(
��K�A�<��ޜ.I�y�}�9�ɣ�6q�{������L=�q��_IǶ�H�9���R�ɒ�Qjz~qg ��D�"�qc⎋M˚�̰�@�D�g����A놚�����4�'Ե���),o+��i��W��G�EN_���'�oa=&V?���v0pX���$ۍ���L��@*q�܍��T��a��Ɛ�Ղ�]%�1wIaZ�s��?��x���m<���.�Y���M�<'�h*�15N�C�M�TXB��rpTm�P?<-��7g���NڑK��H��ҥ�Y��|C̆CQ9�Yk�s"���&AD�Kǟ֌��I�KO FZq�R�s���]�3�=��jpN`K��E��% ��N:�r��h����o}���@����P}���f,��� MEG'�$ ��+$�H�<8#���Mbm]���*��t;�� ���1�{!��˥!NI/cl�δ�Ѽ%��P�֡�!qR\I�
�us�����D.7/2FX�WNq���`��'��i���]7��2�l�n�����-�@@�����v�lox�cL�jl�XҤ{Ű�����4���[���M��@+�$����g�#q�n��y�Wo��Z�?G�)Hb�������7	��-�˦����i�i&P��<V�+u����"��-�Ј��e�����|Bf��j����������E���o1�H]�M#r�A��#=t�֍�O�ag2t��/%�\��h�*E© ĸ�oѩ�t�T�ja(�+�RZ�ǫy�Sah�!^yd�M��5-���z��˥B!��4LUN�r���̡k����Q�YB;��ŅQ\Yr�*jϹ�����.��zg����4������R�����)��aɤ9��G��+������� 4�eN(w��/����:�(�= 8���-��jh������������od^|'����_���!���E�:>A�A�a�B�ջ�JΥ����Z�(f ����A4�_!�g���.���8�hd�0��w�ʏ���Y�X��+_�)�v��4>J���V�VT����}��� �'򸱙k�4��3��X���
6Ԯ-W��`_mw��ٸU9�w���R�7G���m�Cۻ�����`��PH~F�����Y3l<�-d$1F-V*�B�!��r�2��S g����֋�a�D0i�2�$ O7讻e��L���֧�ٲ�P�ޟu��!W���?F3�� l�Zhg�"�wi��?��h�;�^[P�p"yxaҀiH�p��V��@ۋ�| ��un����xP[['�\HV�a�ˆ�OC�}1�uw��u�V��A�`��Ebx޷�&@�OJ�Լ�/#rZ�yB����Y���Tc}�^�eNwj,ϵ%�@��lS����˅�^���΂V�����#˗B�f�G4
�|� ��kB�A),X�P�`�lga�`,��m�ę�A��׊�(��̩)#���G��v�K�f{�;�o�n�D�n�^��ZD�;��F��{�K��MWN�S�w�i��0,��!�xM/0{"Y�{�(Ц/K�j-0lX�?�UN�E�h:������}��ɡ���Ş3U`�tsA�<�]�yaW��Y?x6Fz(On��S0t�Iqʲ'�؆����o��c����̟q�VuI�v���m�KJ��ynjW�s��[�Q�Ǖ���_D<6�0�(�߆Vp"w�-td�&�R~a�b�C��,:�s,V�ؾ�D(T����m$J���2nG����e��0@��P�nk��e�jM�t�+1|� 3�X_���	�_)��
�>�@,������6�e	_dT$�\�5K�e��A�3�y��{����dHr�à���5�]����b�f��4~;���s�����C���v[�s@�5ν�ū8g+����KU�T��=p�\0�]Q�L>�ԞAb��[�?�3m��2V�D�u���#���Vxw2�E�ڬ&btIܯ(䇫]/q_��K��q��l��%�@��Ih��z�B��M(t�S��(����ڕo���<�9����~�O��1ɢV�q�Ep9�<|@Ί�1������5 cӤf���2Ѣ�H��p�_.�Q�#�!H_�l�ͼ���C/'�J����򗻷pD�� M�b`�)��Ђ,�&*ō�� y'ݐ'�� �0�a���yP:A���e�*v
��z���(��w��h}����.�>�\:�Uφjn��v�Y�"��ё�/���:Ϩ��u`�N����	�c���_��T�-
��� m<����z��d;���!�=�G-����3�M�_�~�X�x�S�a�2::�a܍�)G�e�� ��5�#�9�t���r���_��!�$7|��uWí��K�0&<O�y�`7O	u9�+l��5�n ȳJ��H�X�r+b�P*�oɮ���*�]:}�fj�����IB�	���vB;9�\���T�+�y�a.�8�_)�i��/u�2���y���O��H���_:������ծ\-�$5g��Dg<�d�+{�w�j�*��M�i�h��l;���J`��r-��x/�.���p�[�0��(6���^�'`��(�rZw�N�h�i�~f���s7D��6���Y�y����t�1�ԍw[P|� �Q��,ЕsL"CA�N�`A}��[C�wd�ϻ�K75�eֳ~ܑ,�b|��p���w�1��_�6�������+�����h]�ü�a����(�Kd�q!�^dd[�U3�� P�7��{U�l�y$�\�uQm1!���CA#��z}�G��0�؅��2>��� �DR+Ȣ�:���ؓ�V`�|��\fH�j�֐�1)jf�����6���ƝZ�Fۣ�ZO����/G�� k,�Z���u�/�T,�HbZ���$��Q�c�k���U� �s�b�(��&�@G�y;yD�0�0���%�:p�S��3��,���Ĉ�?SJc���HǪ��!�>b��nyW��1;�f,���V�h��2>%&T���b���D�B4d�����f���Fpڢp­f�N�&��I��nW�*��Z�%&�uDA� ��%`9��V�u�0�*؂3l�$�pt���W,�ڴ��yB�cgW峰+��z���Qvx�\c�p	���sbk�^�F4��86���������+y�[�W�@��%0u�{p �eٷ5��IN:�k��Q/���?�^����y�x�x��D� �4?]ة
�{�t�Y�J$ǋ��:���\�#�gR��pd&{� ��ꅽF�u���c�o�-}�vʴD�L�|6�0���zg��R�F�iӴLĀu��K��YǅI��l���U��{ޛU	�٫��3��+�U!�đ�0qR��@?��ds�8Qi��'��D�)Hٱ�H��X��}�].�!!�96�A�K���(K1N\f9O"�S�S�BE��3�����yѶl��Ad������S�nҦ���9F��ұ�8��T'��L4���5�BZ�m�C��֝"u7˺�Z�)L�F�
��
�-�&����[���`��%�!i�q3ʦo��"K]�o��C`�{����R#7�4r�5ALj����l�j�Cn�@ߍ���y=�m��{�P�d6�,��j"-R���������T��l����s���9�	�F�C�>N�P�«vץ ��ǯ�q��#`��l`���!f�p���Q���_��C�q1�(Unf��Й��	3X����Y�])��aZ##��PIfk4��	VߟD	_���k�z���ݿ2i�U�J�޻�+��Y���қ�\3mR�C̬���T�5T��oO�M�Xxƕ�ǚK7����4��$�S�:��$ �	����|'Ev��D��1���}��ˇ����e���U�':#�R'��0H����7(��ad��Ϻ �� t~	��P^$:�.F�P�j�\��4Ӗu���Pʒ��N�w0"i��1�B��T�j�@���Y"QF�O-4�۰�|`�����e�#�!$	fu�2��O������;Yֿ��3~ϭ��
߀?PX�[m����]�=��j�0|�xD�S͋d�~����0��e�*�o2�;�ɜ�����\p�@��j�Y�N`��O↌����Y'q��3aT �Pj�r�:!X)���-�1<�֐����&���O6�|���R5 :!Q���@1z���k�5��Ŧ���i����G&�{ ��?C�T������U��ϳ���O5�,�i?�~4\������ÝN��:����'Z+����J�-{*r1��й�[N��6,�R^�����7�˛�� Aqл����{�ii�蛯�)��J�Sgq�`�U��{��s��0+S[|a�wfr� ����}T�Za��0�j�]|!+}��F,�)�����{��\H\�&#x���䁒���~Xڮ�����mp�`Kw��<K{����5��C�K��qC����N�]�*jP�=���&���Sظ���"����2�9�Au��;�\9 bP��iaO��	�E��VJ�^'i<ས�M�{ṧaC=,2§)u�!A䏜X���Ӛ��X٬y�[�6��l%s�e��i�~�����S��K}Tz�v!V(4�cz��D�}FJ#L|��S'���h�S�]#\�)�c�p¥�?�^ӛSVA�p����y����#����aE����l
��>O��^JZ3t�,� 2�6��.��jts?���=���P/;6c��5����*�/"h�D���;�J�j�r��(H�Y��꯮k�5vN��[*-�4�n��Q`	���]w��z� ����׃X�߁7��䘑���شJ ­?�?�7 -�����b:���~dO��Qk[�@@�u	�0�t����k��8r�6��S��U-X��0���rF+~8XQ����d'do��󂽠H851M �Pkϳ7	�D{�����������R�a��<�����X��L|��I�@5�]ʔ�Â�ҥ�^4�sF�~B=�V�`Sp��v������p����碩��[\A�E9�/� ���v۲g�m6t8a��n�L���K+���C��冞�5gu���9��Q'��ޭ����I�]�q��}F�_�}��j�QxY�־�Fc�����Ԡ$ � J\����p�
�a�'���ۃ�;e
��E&T��{:�A^e0�?Ằ;<R���`����h�H�* S�!�B�o���i�?^�m���@����o�	ke�)���.n��:�z��ћ��=��s�̦��c?�{�L��oؙ�8�bg�x}�Mlm�갊x+G��vC7�ax�P��R�1��%<�aq�K������%�T����a��] )!����k��A��Ķ;��N����ZF(��'a��˧�(/������|�Z���M.��7jp �BI@�a+�ThU��������B�#i��$���������#�4^�G�v�����2����ڭ	�N۠��4>�-am����UU������z�I�U������.��;7bP����	���=j��DdK�n��7"�U�(&�^��o�S¢W�<A��:�ZV���kWT�^O$lj�4�1_��B�J��U������/�O�!�E.�uޱ�{p��3Ê������	�	����䶈,$�S�ѠA5*{�Sr~0DZ��~�ug���
3�ImP�!G��#W�� |�?��|wd���5H��O�h���md��F��1�©�B�����S��)�(��.�[+��@"�G�a�sحe��R��(#C�(�r.J���\v�ɼ�~H��(cQsܓ�0"6e�O���}��V�1���̒x;vI��O�@����JCY1���ܷ
��uk���ܻ�AE�媒M��tY+��ϴNδ#^�������!F�A΁�ŏ���<(�<��^d���@��.���iqL7����u9�c�xۅ�Dg"�ȉ�}<����X�	wz�۩�WdIfv�Etɱ�]��0��GmY�f�Oo#Ĉ��҇�1x�;�s�2�B�h�oO@���e�#�U<��9�2�Ȋ���O-�7O��(G�)�;������R1�-`U�����_�Z�F��������d(��"��v"�m�1��x���7T���6x�ɀ���uO�b���g��#ʴ�d_�4{L��C��~up16T���2�n�(a 6},H<�Bub-�_M�c?o-_�`G�Ҭ�\�G��N�m�E�T�����2HdX��B��u������N��3RH#�^a:�\5�^w˽��}��^����CH�-@L��?�𝒨*�J��M �}4�����x����T *�Bzl!I����)�1�L�^�L��ȿ��]�H=��H�#/��m@�@����F�H��b�ӈN*Ggf!i������ɵ�%K1�w�Y�E�	�wkW��8��A�P��A@�j�V�1Qj�Ž@?��Ժ�R*�O��3\�=�^��1G�G�ю��������p{�p|�I8��I}��UL�������kz��T���7/ʀ���4Q8v�i��V��ֶ�� ��:�B�'��A�����k>�m*z�&@4r� ��n26Q��s:�3�J:(W|����6_�1�e��F��]Ua��� �H�9�Ƹk@Z��r-n�o��-�oG���QN�}��=�4Pan���v��qy�|�635E��tzn��&����A)����ۃ$��7���#�e��G8wI�W!rsZ�`Hj��~�w��C�9�ӛ��V��N�(��_�E�.XM��}�MI&�QkC:3��9e&�yD�SKj���{}E������RP\�ܤ�o�m}���c!�Aͬo�p�L�@��?�\� R�]����{�-w��<�`2�4�{9j��z�7�1"�x+���;�~�o�>;M\�纞�\2�knP�x!\տ������z���Ȃϊ������5`�o5%����UفZZ�Vt�� >���~�*x���[��ē,��	R��Q���o���l|f�b���9�� ��^�Q��������W���4&�.�I�n6r'!�&��[�2oL��]��A�>���ZJ�)� J��vHΉ�8�5Pΐ��J�n��� ����������:E�(�&���۴��R�JQ�'��!aʄ�L��m��P��4
��B� I�RV8iR���W�y��h��ELY�fڍ/W�/���I�w���קV�Գ3�J�V�O�.~I�&r��:�k�i����Z(�]_����m����^���w�]��DhQz����5%:� �Vײ�gL�)KOY��g���"h����	�;W�k�!��o�v�8��f�N�J�3.kJV�;��HG�c�f+$1� v|��{,`?s�Q���Q�Im����fͫ�+�����w�1[i�k�\:,�����UX����k�K<�����ig��YJ��/�c�::.�u;O�2�cǳm�q~�Ox`�
���m�xqWn�N}��	Y��+��	Dv�����Z���8f+h�qn�LƬΚU�����H�l�������I�8�;B�>�ϜAdnt�G,���x�cQC��2E ��m�Y��v���Q���,����g?��w̿\�| F��Rms�i��7�<U���W��Sc��w�z��mE�Y6��?�Rnq����L\䭹��8,��?�?�C�L�H��$W!�8�cB��
��?�s�S\�8X$��f�E2�r����kW7���(s͕��-��2Rs�#j��rE��E��UO�PI3Ƀ�~(^k�v~=+�;m��2vW��6m�I��!-D���?�)M*]�)q����IR �МΕk ������)4c���N$�:�"�&�yX8����-*�Ip�1vB�����u�tT���M}L�� '�>�>Q(H��P�,��u��~�^����r��@���m*rME�����'�V�>"�.m9�IY@�3�$�e�I`�W0�Mt���񮙶u(���R4@S���X�:[�
6�l�pR�Հ+�^\�3�h��,��2`4;-G�����M���`$��U��2l[����l��m'E��(����c���]�������go4�0�F6')�G�DQ[Q���MjT�n��M�g/A�^�� ���ަ�@�M�������)D�@�*eC����LG	o�H���Vٖ5���f6<Y=��
(�O�ó'��!�"C� H@Z���O���PЛ<uLK0m�Ĩ��[�h���x��f@�j��Psl2���4�}C��Y���k�����vW�qk���"���3�Ľvk=	���O�Y�-1�ǽ�}<`�1aE���8�����3� $	(�q44hh������%}#�j�	����kK�1��I|��U�2����(��r`bl�i�6��	τ 0�� ����A�:�X�?��3n @��$����@���A�9��|��^�������{�����c_����r�"�92vn))Ȝs�7l�ҭL��9�q�_�~���RXZ����k)ظL��{ڒt�KDf)�z]ۍ�TC>���}��c衝�Rk%��N�\-d�U����sCᢌ��K�J���uL��O�v�X�mZ@D�Mhb������L����8�imD1��"����	[�XG�����1ք�c%�!������LF�Q���n�8,�"Z��#�.އ�\�
pd���^�sfR��*[ό�t�S�0��r|�!���3�2�LdJߤ�	���Աi��n1n��	Wy �/�@�?bv����u��Ol��P�3t�g��I>�t�	������9�~��6�V;���v|�$�}���<�~�m�{��n���c�?��hy���a��p��v{ա�7Ϳۅ��P�_�?9���Q&���Z��z`��İ���l�3	pk� �E5iji���<������~�Bԟ�f\;G�Oćo��22q�:��i�pHm�a���J;S��Wy��^nR�ο��
���=B��۲�k�3:&'����WSL]S�;����߾e�	��,]d�Q��`ܿ�n���1L�t+DC��I4�җ�>�+��p��S��S��}�V�䣻�o�,,L��,���U�!3�pD}�2P��O6��Y8W��Da�SO��Θ<-��l��'bKUͽb��ep�ʟZ�������O��kYT�lX�<���
s�h_9�8�V���c���V4���& ��c�͓��X�\��[ޜ{���=50���Ў�>�BZ6�-�o�[$�>%��F��[+W8��������h�c��:5�-����h�!�9�ă�<1��X�1ޤ���n9��'6�:E$��}�Q⣎@��F�$A�'���������.~g1�x0y����wP>�:(���+^6.���0�J3[�_�;U���}���L��ZE5�q�{�x�X�U>r���.9p
� -'M�)���g��/�3��62^�>�=<���R�Th�|,��w[ݳGZ=�G�jc���0�СSZ,|,�g�hn�z��d�߰�1�=汎_���(�A�-YI(k��峨�y(��,iX�B��H<{�F'��5��-��aW�3r���.�K��VH�d���mp�={F��J�7��]�^������j�E�P���oz�\����!�"���K��X��:̧��y�d|���C>�W�d�LV�nm�=����at��E3��GV�������ԣ�L��D��v��z����gJ��W��ײ��߃�vX�B�D��%
W��9φ�/᭓C��z'�\ab����z(�	�	X�2;�%�r�9]��͈����WDZ���ܸ���~@h�;�X%z���C���,!�R���ŭN8� x�݌'���q���f�\ݘ�L[��.)欵�cK�t=�oD�L�\&x�2X�D�led�Ν.�Ig��Yj�XѪ�"$P�.�]6-m�4�Sv���EP)���A�(��v�46����i ?5�l�2�He�3q�`&���"�Mr�r&a�)籅�8K��G)��^�@�?�WA��gԢ}���8�e6VLSE�& �@
M`���)"��@�f�&�b/�w6��P�S!/`r�z����&����S��G7��!���ၩ�����TS`P��.�5�O�~~�Wc�ހi��8��Þ(��j�4.���A��kz�(���PMD|��_&��̳���
v�A�,���R����uu�u{�� ��g|�:?������ ���6�h��Z�aٜ���^)6%J�QH������+0���{8�bo�P�Z⓲��,49/Б�X���8fD��
��e�-�>�U�vR=�����ύ�/���7��qA��m�hH��#-ʉC�,D{:f��0�+-��3��mXҭ�91�C)t#���c���䘙��b9���+��0iaS>��9�#`��Ɣ���M���4 (�6�l쯸>M��Iњ�P��N�7� Q����/a\�B�f�w�7�gj`@�H�(H�x7�� 1*պsǶ���~m#HL�C��ZE.���g��2��x��S�4�{�Ҭ�P@.��Q�yo�C�8@e�Y[޷~uv��x�t,X91J��2�Ơ�/h��v�Ǚ!��P�Zcy�`wT�V�S���꤇p��#mKp�\A"���_�� ���z^�`.c�M�j�l�$��f<�9�����h���k�����+�����s�=2d�{kw�ώ�p�F:�rΕ��4��8r��5�To��A�_,y�u�;7���8�`\[8��w�d�:����F �V�]9ѓ��W��X��Bi�[&���TU+��.k�&�3�R�cUI$����ҳ��&'�1t�?s���f]dkx
Iv>�
���L=��lY5]���_g����/�O�v��>��7F��5��R��|m��r쁌t�,�+�Rk���k��@�.;Fj���5v��~�ڐ��#� S����@7q�D:�\�k"$愜|��;�:��s�#O�A9E��gNr���Y�I�|gŝ�� ��{-?<G�������?041�K+6�y��r��������	h�l�7�~�:��c�_v\�|�s�ܴl�7��������(����`�ͦ�?�C\��f��"�W�3ub��4�<�ɓ�Q����B8�H��cF+X@`<�ܫ��o	u)���_}K�B��ay2��b���pT�� f�*�;l�#!sMJ�+Mm;�E��n�5���^�S�	����a���[�4��6Y�_ޗ�^�\'���G����;3DCV-u�3�f�N�!ݶ8�� ��d�,���PS�q��Zd���*�Pw>�������ن𼽨���+��������s�30zcf)��^��_��G�������H���Ӌ#�%��Ѝ�ܖr��%9n!�-+��-�o�M���!eJ��T3� -,:�Riw��c��յ��LЅ��� ���ֻL�OzƦp�����]�J��Yf.�!�Ve@+Q��G�z���C|<�8 h:]@4,-��E��/�u�aU���bڿ� �e f�|�^.��)�\����-ѨU�}�c�pe�\7����1��Yi�>�B�^M_G&�*��l��LͯC葒j��4ci�J��<��:�6��ݬ���{ޅ���	���;���A�}-ӣ�z�L��dw�p��J��v�`��K1���#�"�[D�g��!�K#R�Q�v�MX}�YR~�Uk	x�&��"D�.4��{�����S�i?��Y�F*W8�d&�c��'�*���=M�P��-�&��k�����j��N,č����aafŤ��؛ ��Յs���u��u�7ў��Pkk�� %���O<A��-6�Q���"���W�˒�*��;�z��&�����F����ϼDF�b:�/�C�s��#���b1�b'Y��+~�,�����P~�x�X��,�)�{l��~ .Vk��~?������v��H⵾�m�% v62z�QIn7ׇ�Ů�����*A`��]f������Y)d}IY���"x�<��`���vx���N�y���4B,$5��KHi�9�Mk�g���A�9���;��C��),Q��
z���Qa3ƈ��#�������v뤯(&l��^��*Y�l�d4Fy�ݡ<rs����d��%��\#b�(���Y�!鼌�A�6j�뉫vȘDq���%��exܠ�To��N�Io����خ�Y�-GT�3�kj�A%��I��_�g�q�M<g2�d�t�9
e*�d�z�bWT��$�m�:[����p���K�p�.��`'Q���ny�S���>��'���T-��nQ;��`%�)9��bR�a�,0b�ٸ}�r��H;-��Jj��6P�!aU*>���0[.��k�R�.�wq�����O3���-�	b�NTG�(şs��������˨H�D����so�JÎ���J��a����1�UBI�`�ǋQ���/�2q]��a�,�l�[�@G k?��h��5�뵽${�2�i�������`{�;���A;��3���&![���_g�R���ϖ�2vs@ ^�?�y1%�*c.ǘwL��_��D�[�M��Ӥ�ߙ���F�>�A��I�r�Z��(��%>��ۅ5��_I^�J��^s$}��$Ƞ���Ae_+BaR�����e��`�lNO<�R�_�d yY,��}�o"�����#<�����̀��v	v̰�ÜIƽ��cpQ4
2t58�zk�,hFЂy<	��G��	\�4���d�QP�������:�ݵρ����k�h���g�& �7+������,?'8��ؒ$�M�bY�E��;�3r��b� B�:�3?��y������J�od^�İQ?"�n�3M%˳���lA�)������@�/�RWK
Abyf�����&��$ ܐ��\�2�_��̻f��;�e�BR_N����T������)��ўY��ޙ��nbt�+�>!�Y�{}&�R&@�3r.�Z�0�����a3M{�@Y�obO�@ǉΊ�E�RE�����}�TF���r�p�����*��&�4�N�|��ݒ��*�1\��`&m�"�m<�������>��`��@����P� ����,H"_�7+d�%�vxD�8�ğ��ǋqv��� V��MI=`��='�D��iK ��Jn8V?��
�Y���N���Ƌ	����)~��HYK�����̬�"�����/Q��ղ ��O\T��S�s��r������&/�Q���۪)[�NBxW>��j_�m^.ϗ^��`�*3�4 	���� ]�苹+\��ʽ)?�1�Zy�����{܄�!��36�
d���N|��f�(C�"^��/M���NÅ�f�H��9��7���_�Ȫ����M���m�e*��[c�T���Xa� ���>UDC[_]��F|�
&��N���+N�Hh�
�ڋt�
L��:�9���hQ�H����F��^�ĝx"��n�i6X�^�a��#�хe�z���+[�r�U!��6��o�^�c1�gV�Z��[���2_�v�Ec�&�E��YM�F�"���FeN �n�Ow{x73��E��\=s4�h{Y\:9P�3��~9���B�PW-h���gi\�Z
�<�ҝ��R�����`�G�d�0Is�/���/�N�b�|�>�_%em`"�
Mρ���eԟT���fU\� *y
�Ȏpݙ P��Rԁ(�Y��k��OP���2���`\�U���#�6��Ǯ��Y�(T�<?Q�4��vD_"M^�lX���95�#m!����B�Y��k>t0f���j�h�W_�8!�=��Oٔ�t����S�{�`�Y��|o��u��-�EO`cM�'R��Z���a4�B�謆G�4�In�g�;�s��q� �SmJ�g5�y�E�}S�n�D�U�����&�]�^+V��tu������<�$�{��7"<S6yU�G�蟢m���B�����ۧ�F'an��tޥ��8�j��)�ѻ���&��P�w3��͞�u{�C7�X���``����)ݟT�^f`�s��מ7��Œ���������o�SH�ؘ�J�͊iDJ�D.�[d��Nj�:��f�0�3eX��,��F�W�����8)T��M����6��Q�	�JpO��]�kq?.�q��`h%�U�v:14������>�����`�������žj�G�� �LP��u(���j��6�"�G��S>C77��yB��ME�	
3��'�����(B<8���~7�A��Q�����YE��8*2Τ(��L�f����=.��6�Ҽxk��0[��:"�Ř��gd���l���jN��o$���V��C譺{��0��#�7�?�Hy�zs���n���4�������;*�r8`�旼�RsP���ңް4MQ�0�{?�#�;
� �b<����w��(b�ߜ�\���b�@��\�X1ľ~�d�b�N�l�ޑ�DL �3��������PpT��	�1���cӒ�����e8lsB��T��&�4�y�U'��������x1%�^�^�p��AQ4��z7�����D�)��@�/Z��/�� �d�uz�jcx�0��|}�`X�ݼ	��א�N��"� qM7�9l7�w_~�H�Y�@�s�rעL�����j�un9@���HVx��O7�cdeΘ���ܡF7�J�m�]�u�Ю�p��֠���h�n<�e�X���[Nc7� m��0��R�V��P	Ftu�1�{1��ι��:�Rx&u8��59Yn�������j��*'?��μ��%�����w#��G�-��6|�5w���j՟Y�l+��$�t��X�V�տ�P��h�î���g�n�bi�k� �S)��ݯ�_ q�|�r (��)��| �#2q��(�c��R
�r�Hx"<��@]l��������\�A-�"�)<Nmsu	�
DÒ+�tI/bZ[������c��_?,l(���S��:��A��|�M_K�j|d��"�ֹN%��L��!��C�E�< `����'��5F��� e�N�.S�:&
��$ ة5=e��F�d���}Sg03~�⟛�0�v��dWd���`�4�.�f�rq�mt�u��<��p���.���^��u59��ƪ��#��/:�1:���IY��j���n���WT���d^��#Ʀ�!2�ig��5�{laX��m��ZFO��~v,�܇#Xt����������P2u]�����L���Z��[2P��;�5�w*�������]#\�g�I6z�"�՟b�5"�J�e���;���IHP���}g!k�df�(I�J�R�J�q{�e�aӠ:�N��v��zQ��[ˀ|(%��啰�>>Z�/�*\`/K>('��^ �ﱭ�f���Mx�IC���]Zx�.7p�"潕<����f�`0�YK�^%cc��6w+JbM�sD�^�_$#&���g�:�86�5@"�!��`�2�)� ��"wM�T�t"�,\&��#� ˘���s4�J��@����ϫ���]~3�g����KG
uE�F�e	�3������)C!���� �L���S|�W~(�(�~���o�BK�p�2]�\N|CTd�v�"N�O�V�vKQ �%L3�o$Sb^nX�1��F���x�\�~��)�O7Z�E�MAp؛��eG�$��1h\T��ٿ'���{B���TMg�J���և�V�>�[��K�i��V�����,{�Y�+��IB陜�5r�=DO�>L�)h��Û�D���N˶2�G:��%r�9.r�a�[�f��_Py�?ا��+���BSO�L��]dG�J��ϸ��$ �<��FB�M�EB��G\U�H40~��Qg�c��J�1�v�h���"�a��E�U�����
���|�Щ[}ՠ7��I2j��w_�f�?�7v�v9/�����@B��ٶs�����Hp�1
h�C:R��?⚱�Y�����0�n�y	�mI�T�����ۮ�D/^�?pnf��㹔��.�^�r�C[>X��2��ږ�l�Pn�7&���x��@������\��FK�����2Vd�._J1���Y��Ԗ��'��Eܟ�T���q3��cr}]��s��m��+��9fH�@o��P�zcsZ���|�J�=��Ϛ����[_`�R+�a�&�f�T�-�n4V�km�z��HM�pk��!����4���m#W�y�����#��aكXV���u��#$���jg��C#���Nf������$2�X,tpKI�:�Q�s<W|��҈hr"��|���-�DG3�p:O���W���`NvxY����U�T:��t���䉓�q�w�>�I-� �!�x�����^�>_�?���+��h''��B��ˆ���'.W�(�6D�I���E>$D�-�< ڌk�l�����Z�����Yzf�)�2nՎ�$ݮy�o�1��7�l�>��������x7.��w��d���:R|�Uh��eG���,i� I`H�g2��&�"��փ�2*���2��շ�sf����
�	����͌ld��M\�~~����c"�S�!�����%<��ʨ�!wX���	&��;�2
��H�i�Z��xp#����ĵ�lQ�*��o�>"G攊�y-�����I�s��`U-��l\�p��%0���'��-�2c �ک}�%�d�!��*���QY��%T�Žr�2i��m:M{@<��4/u�ms�����l��!�/���]jڝFTk��Ҽ*�q�����3����+v)�������z�oK}��d�r�vO�W3���9b�iL%������6ht�4*VBN���v�%[L��#gYV�4YAf�-w����ޝ���`����vo�aZEF���,��2L�)!B�~��/J?������UI�6�8�5������fy0�mz
 DJ���߾�����^�P��u�+�"]�B�ǎ���d�4���@M(u���f.�*��\�#���	�<���Tb2iѱ�<�?3���L�0��m9%�#���&S���ydM'1ڈ�kc�S�f��TgS��}ʉ��y��4U��X�\��d�a?˸�G�b��Fa�T]��{��]�؊i�@�����k����к��S�a��O��pjصֆ#��}�����*�S7��c!i���k��7�Bx�Y���mTuހC������dS9��Y��d؃��b�P2+XR�L"hQ,2Z̆/��j�z�֌78�NV$��s�S��ŗ��Hn:�C�'��|`ۯ{�=������~4~�l
��ٚ��i����t�\�R�LU�'cm�l���2��RZ�~��
��^L�f��(�)��B\���]=�ΰsV��ɍ�:�c�X�P���.�[�l���fa�n������T�T$��HoL��c��se�����ͷbH�U��N��Y��,��Y"��A���$3��ē�UO�Z#��Y��,�J���#eu@��?|u��hRpA�L_��s��E!J���G��͸"#'�_�����e)C����b7+3���:���˾����u-���"6��g5��4V��7}�cᮟ#U��j�-�|�"�{E`�79��	��V���jٿ�I���1F��� Ѳ����K�\�'m��Pp���G����?������u�M(=�s߯���M���U��B�&GS�Ft��"�)�[S�3	�����R���x5��-5Rs1G��0ە��:�����rt��)�&��Z�5� rE��a�q�hY��SHhؒB�H|,W\>��<���OA���~5Z0F�DԿ5#���k�M>eۀ���k��٦\?ܬo�lMF��|�	&�SS�H�~���%�8���1~5�v=+f�/V��~��0u�T,b����;���Y���,�eZu�L��+>7�n���Q��C�3�m �\x������^�Ș������C�v�#�)9���9,òe�4Xsұc�ä# �̷%3"��'�1E���v�Jep^��U}q˙�ej�AB� ��^�#���'L~Ai�����N�'(��"fi�c,�t�ο��㛃0�ǸN0�Pe�W�7��r�
w�k.ֆ�8u$`�ȩ�����B�Ԙtx�Zڵ�H%�H&؄�Ѧ_��t��fA����������w-Ṉ���T�Yp�^u&?����>�K�����87?�q!��E�b�˓��|C7��1ֳ�	a���qiR
�8i��2m�C��SJ�֧�#��)��	�¯�X�?���������u#�6	��V���6Q�|����V��;��w,S�H��$�+����8�!��+ y�6U�� yy��D{{��O��ќ�.�1 ���kp<�=�$�Ŷ��Z��]�0~C�tg]�b{���E���#�.�jkbZl�e�F*��d����9,1ײ�+�#/WC�`�B��	ɱf��l͑vs�@eA5=�S�P��
�� �W#�1y&��ΨsU?`Jb�C:7���p�x���j���?e&�<��d���D,7�2��b�����\܂�jXzR���k^ߛ8F��92�̒����Y�F��I��m�dWmҺ�_+o3Y�v�q��G+m��H$�����3|/�
�d���Q��N�Ƒ⤠}Uۻ��숨&�,5�k�OЅ�m����7&e-������r�~dA�GS�?2
��D������w��m�6=�v��+G9�7>�?�BD��+��tJ�2Q57��D�RCR��;8�/�9���
��6�?�̘�9;�d�ia�.��K�H� Ie�O����0@��X��-aAr��A��]7�iM�LF[��Wܑ�,nO��*� �y�P[���$qM0���{ɲeҺ"%pĴ����ya��wmL(�_1�/�~pH(���Y$'g�{.��>�]��װ�Y+����������,~����"�E@�r�Y�h(8��|�O�S����o�b��'`��x>ި`������2�w|��)@^����.k�m:k)K�� �L,�lvIj�Q����W�A̎�3[Q)��TqY%���;�
�!��nHy���8�dbb5��\.��T\l��bx�{���i�,�vj�9XYmd4�v(4�7HC�R��k��qQ(�an�\�ֈv��/��.��+3�&�fR����}����g�7�Q�j��`��WW.f�q�J���P���亨��.[KX���[��%	�HG�.�#�Z��1�Ål.Xu��t�*��a钌�KA �l)��:�}1L9J&y��c�\6~*�G�i>�GE�~:�̢��Â;k$ca�r��!9�0�YW���G�bdN<G��i�ws��!:!��%2�n,�op�D̿�q���믈�-:;K���̰�.n7���
�W�dy�TV?�2���D���a��ytG��/C<-����S�|u>b'����MЙE�3���t��_NCݼd���Ю��Q�Z��ץ�p�ӛ�z��z���M��.	/��|RaÓϋ����
7:����:����`cmn4�[
�8�u ��	�x|�*x�@�m��.�E*C���M-R�g�;�Xk֍}ǓS�Y��:�^p�tp2E?z�o7�%$N �˻�L'U6����ߵ2���%��8�9֋�A?��&�Ȳۗ6㌉'(z����֯� �
M�ŗ��_����h�7W�B��Ĩ�N	�͐1:�7R{�F���0K�0k|���[�����"��uB����~��٠�svT��R`M:�؞�'���?�Oq\�%�´�PH��IX'����C&4�qT�HƩ��wl$��P�ly�q�G�P1Ffs D|+�K�`x̎���t墋�N]�_����F{�I���o��_�v�ʒ��{���������E� ��D��?{	w��q�Q�ގj�e(Ӝ�,u���4$]�|�&�0�Ϊr"����$�Yܕ1Jd^�ű;>�XU��U,#�`��]���E,��at`_��Hmz{�A�M���돽Y�\�'�T<W >� A�=��B�t.[�[�e-�ٶ��o�$�����3�SkF�z�w$a�<�B����RRJ�WM�V��q��/.���.�$�:2�l���5��26X��li9�P9��������#K��-�$�MBC�������?E�k��J'+�e�EX�7����m%��K��GTje��'�<���͢���r���D��n��Pq���5����v�����{�x������4\$�vU�D0xQ���$��EB�D��'�����	i��*�T犁�/B�U9B�"#��6������i�̕ޱ� �> ��zS;Ir �X��,Mb�^�����'ؾ��H�K(tF�� h��X�d2YKFɘb.l���4M����)���pJ<N��������d��ƻ��(��C4�r����|{�Ō��5�qȻ���P</�DU�8��e�CmJ0����UGkg('�U���&�f{����DҨΌs�s��
4���ƀ<��A��%����]xPd���db��#��lɚ�h��P*&�[�|��0��U����b#����e�r�{8lA�O�>��"{�<J+���Y�!8f���q�z���k��v��:Peϔ���(V���T�8t������c��N��I�&�]�ɫ�t�"'
6U�C��Y�4T�k@?�� �B�!4����Pj��~56͔c��\e�P�[���q.~�q�����0&�m�0�:dOx�/e��?#pA7ǈ��/"�@���>1%h��>Me8�ܰ���#��i�����:-���IC�£�$C��;3zE�E��B��p��)!]h�Ȕ�Z&ھ��7Õ�x����-�sajjg�ņ����j����0v3��8w��Ѻy��,�����N1�����F0k�S�.`��A�'v���y���MGr6}�\�4"A�b�y��f��S|Ƽ�LWc��[�^ _T��1>�8�ɮ<�������#�����o����1����C%�z-#��6ߍ���%|Z��Sb"�j5|N�W7i%�1ڎ@���,���5�y��Xފ�Fo#Tub|��|7K��zM��_�6$���㑭�$/���������c����z �z��"��TԶ�ۜ�H	d�d��?�=!$�_�U��q�B!��
�,u�6��Q��U��'���{�Ǫ\��b�G�E�Gn�9}HD�׵`ș�X�N��2��o>�ɢ�ƐR@��,�
c�:�j8���a���(�����YHU�����02���cS�2�����<a`��K>��n��J7cf^2~E[/)����w!a��ߗ]�8�Dƞi��@-�(O��z���&9B��
�qj�|�A*�▁MIҟg-sА2�����	�[h�W#@9���g�(�D��P�:2�WV��?�:߀�܈a�a���/0i��'���|��O�#QF� ��"���U�]P`/	Q�5��y��Ӳ�*�k���X�3pw����9��l� ����G)�ű����̓�jy� ]���.�H5��o��1�>1�����҇a�� �2��k��� ���6|iO�82@��S� U]�4<Y��*Dzw�Ҵ�G/I~�H�o"?��,t�h� B��-rnq��-%KT�UT[��c�X7
�����>�]�C<�'C�s�(0^��%B�B^e��)ȱfCn�g�����y
vNۚ�W#$O�ٿ��s�KI^��f�4l��zz=� ��������iB�"a)�8\�+�������<a4���Ո�����Y�SQF�.��n5�| WA�@�)q[�s$�����4��;�2}� 
dvV8'p�G_���'t�&s���6
��yI�bta97D�f�/��j
<������F�ҹ#z�m�O+o�zE�
�&�O��v���(zعr[�`��+B���l39*�H���r�ߟ��(4����K)�I��q�Dj��r������$&�-�6�)�S�U�z"�k���U;d���B�,����^E�j�(����9g�'���C�f��`����� �&b�'_��Aɬ�Pu�^8���+��Y��X,�]���+"j�����sT;Tu{���q�a�|�U�Ŏ@({U'�%��\�c3W��@�汀)��%�φ�Ҩ��PY#�7���ܷEW�7DC_͌�~j}���a���^L����8ǩNɴ�)%�r��58���t����MhU	��{�U�`�^��b�V�TrWA�>��f�у���/4��z/�dDg��PR1���U}e�h���κ��i5��v���pr����A���.�u��!N��,B�ba�� �
�A8Tn�/]�V�o��բ箲��]�o��6�:x�4s��%��6�#�F��i�~L�x��^�~$�n��Fs���݈sN�;Fɨ0`�M	ڠ8%�ތ��(H��U��%�
�,7�Hl��T	�C�Qd��V4c��6�뉨�%(�uns1�I��ԥ�l/P���sk���n��6��8�R�T~P}����#�s2�u�|�5n�<HEԈ��&�	@�h�	��݋A����B�5�8�Х,�R')������.DU��Nղi���lB�9�`_7\���2����+�8'��ܬүl�T�dD�%����-c��Kw�$r���x��z�y:p|�W�\�eW)ތT�A�3�f]v���S�)�2#���#�����Z�)� %��(�[�C��-��� 7��x�.��zX�G�����>tS�߀T\�,���}S/��n���>�x�.)�2�ԡ�M��t`�Z%|�9�o��(�-]�~���œ�]��o~[H1��RH����x�N,�=�强MG����dd�0q����|����0�u۱/�s�	���[4՜Āg��.cll=*Z��ym�-�ؙ\��_ν�nͲ�bh����Xm�?�f�ʌ�.��z	z�ot����W����@��.^�3@��L�X8!�v�H��Q��<ʤ��h�J�C��H Q`X�E��QgI�\�aMX��A�������a9&[:�l�j\(YGB�׶D����v�%�YJP�6�%A��(���5�N&�J�h�`8�ȣ���ڳ*���'�ŽH}� ,�!PRli[
�Ʃ�쟇 ܨ��#�ڬT���� ��'�41w��L��<�iUP�=Ǹ�Dg�VEU<x�4V4�7;H���Ł��	�cl�Y�I^'�+7U��
�C^�Q��As��]�����}�I&'(6:֪YF�r���$��鉔4���Yr8�΂}��LS����v��HE����j�0�Ly�A��:W�>�F-$t���s݂Z��c@~Y�sd�{��^/�lf]�MAZT�ijB f�)�z�hNHƜe�<�T�?Ѿ�;[�-��Ubh�X,���cH<!w�<�٧�z~������0T����Y�U
g��U��{"zf}M�ʽ_�dH�dH��w���F��Lḷ<�
����d�3�ƂnB��m��`���[m���Bd��ۍ\���*#<恚���/E��CG~	]����oكk�_��W�Ĺ����jW�df�SQ�B�0�x�[
W�W0S}پ�j�����V�l$<&Y����k�e��P�����9�e���c��˥z�G�z�.
�c{�k.��lzX6���� G�</G�F|�j�+�1�<N���?w0'JS$W�d8��ퟧ�0�d�e�.��˧�#.��b㴓�E���4��\��c���ٸsg� �k��6������2_ R��$���ù����{q�ε\�XĘ.I,�,Z�ed�f���4i��!M�T�f2S��k(����N�=��M$��h)s_�����"GAjnf�]�� PF�"G��!DdT�Z�I.4E,�U�=��#7+7�6�t��]/9�..�1��Oձ��*�@H��_�v��{�wM��N�xd���ߏl@d�.��S��)�J�cY\iN����Caa�km�gjprɣ�*`F�6�-Vx�/;*�u�ћcb4����͢�ͳ��lY���ai�=��&����!���k�������I+��|�u��"Lcho>�뛐��էK��<W$
� �x'����'i��F\!5EH���k�P˞���\ݤ36B���B�`YiH�8�U�����P�T��Bj��ae'����%:����
Be*���Cç��i��d	}Y����Y�`�7]vs���'���g?Bf!B��ŏn��~oƐޯ���]���zv�B��'<>��L�F���#a�7,��~ �2^�L�gl�ʴ�{Le�K�{ȹ���#q=%��^T�����\���X�n�5��^�a9�
�c���6?�'�j�G��qb�r��|����칲ðya�� į�.z8��S~�� �Ԛ/�a�����[�e�KǤJKV^�!�?~���)�2�b~����ѽ���y�p�,�ݹ�.₇P�"J*�1��x�ю�ڻ,�N�Av3(DY\
T��W�&3YK�z'����"g}~gXe�1�s���̐s�բ�(L��	LH}\�[�EN��t/E��2� >��F�ð�g�!���L�DE�E�uf�W�cn5J-���Ϯ|����d��� �O�WL++��$�z�M�B����7���F�|���<���s�.����s���.R�9"5�����-\�p2�:���b�=�䭘�x����ߞ%���f�eZn�l��x����?���뀅�ͺ��\=#���x��b��m|����޽�&]�ȼ�]�t�s.�9���rm��hȷ�T�=˟	���e]ep.�t��g�[�0�� ����?��%9������<��f��JTH������z�]��)E@����[�,|PO�c.]}+&Iˮ��FVd�p��W�=�n`V�V�Vr���>�ϐQ�dV��B�W�J���OE���5��{����t_��VU�IY|���G]a!�k�Ǟ��`�o���,�Q��>��uL�l��L__Aj10π�ꍌ���׈,�Hw:��N23A+v?5a�g���s�6O�\4���6��Q����pP��U��k1��	��VO�v��D�B�F�=!���ׯ TK�bt/2* ���w��X<#��qg�К�,C�	}̗j��]:s6'���udF4kE�����n���&��?ΝY�K`w��Eӄ�2����dh�/ܬS1УC%Bj���".=�^���H�r��Es��� � �Yݼ�jc��X3\(&1��;W���u�Wͩ8_(��1r�j�b��i, �𷵜Ü��6�/�������vl���s"'���:�8y2$'�Y#�yO�~���9��c���5imt�^�@mQCEi��w?+�c��P�{E��m��I�v�(���KB�W����7��Id�J��Ͱ�1�ȇ�x�pX�FQ=�$���Qq���G¢� �6�����|��P�� X�H��Ҍ~)�[!�}MB�<�,g:|��V1�qV~��,�9����~*6݄�ٹ +3a��c�iu㦺-{�,�A�=�zL��"�u�(��r�������ʺ�9@(B�=��'���Ďl�R�F��!y1�e�9�ss�!�(����C��B�F�xim�)�\�Yr�z?�ń��Y*����YX�˞q�D�a���������� \���j���7h;y߬:㹅�@q#6WUx�J=�6�͑k9j7E�]}I�v����n��S��e>[y���&6ȳr|\Y��p�K����0_�24��Z��Z�TՉw�̈́�����GZ5�dQT�V 3Kspj��d���:�hl�?7��y彶���;��N���v��ꩅ
;X!���� �Z�-�tVR ��S��ו�C���P�8�vJ�K�p1ɳ��м���e����b���V�;��W�l��Y�V,��F��t
��F6�=�\d�ٛcK�䥍�Q�=|�N��_�8��y�.�ns=_Pgw� �;��۸�����k҇�̯�k��Ah�|vH?+�e�x�؝�ϳ#��� MxQl���j����e�h7c�I&a����}��S>�T�ä0O���C�(����G�1O�E
f�M]T���ҋ=Oq���W���g������#�b���7F$#I��$���<5�<����;9�
yF�>a�[\��qײ���t�}��х�/ڇ��ޣ��?�Ο��fe�f����, �i,����9G�1bP���Ȥ R@*T�@��V���U)��3�����g�Ь����Q���*���5M
���4�M�mQԘڵ���gQ��5!?n�����wp�<�K����NpȖ�v-i�ΠN>iS��Yv*h�xM�F@����w>�z���z��c�"��Q״��AMs3f,=}�f�����&"dY� ��1 ���C!�/�5(��n�b��=*� �C1�}�;�	Haq�� ӵj�Z�f��x\��F�-�E�1P-�x*�����^0��>��˿I��g
��|�E#�9�&�-�u�_���(5z'Q����H�A:��BgZ>
qc����H6 g�)��\��2r�L�h�e��Zw���J��|�HD��E(|��<��e�8]���$!ksW���̄�a��y���Ǔ�&7HѪjj���Q��9����!א��a��,*�~�n��1�C{&��r+$Ɇ�NW�c8��)`J����8~&5���D�6��r��T*ⲭ/��x炖oH��l�!;)�o�3mj�7}ߚ���SN�_6�r�{:�`oru����ay&܁��>���|%(�<C��a{�Ȇn���w K�����?\��k����cS�	��T��.���J�����D�[l	ަ���*���uۆ���T���K9 ΃aμ�?QD�]��]��0�G��|Nq���r(���I���if'�=W�����t�!+r��k�|M���`]��k����*�ج��8����elZv
�ӟ�"Te�N�?p�j�~��,�C8F�U�Uy��B��U�骮F!\/?�M�mԾs��b�t�t^����4yL����٣�wb�V >�����S�Rls;�<6��A�Ed����^9Λ���r�gn܏Y
��@���/D!^���߲��#BxY��[��\���4�2R>�{��m�k�W^��jJ3���8�oc���wi�u�� �Š�J��V�F|�m�]\�V0r2��=�PP�X�@5Ψ#gU߉3���()��BD�7�R���vu��<���H�N���/ �L�-��]5(7�R Lw#���zs�T<��Pј��>)>tx�������!������Sh	اZ�u��n����d7Hds�Z����4 cs��$�Y�&�7JH����/�Q�(R�t���7�Bs�|����k���"�!�s���0��j����aJ)��1����*u�U�����W�q��Wy��cs���<f�	���~j����Z-q�B��ulDK�^�s���'DDg ��'��oD�%��*�"��ߌyi͂ĥ733.!��ܢ�@���x���@V������n�������$	�T���h�n�Tq̶�
<�|iw���=oj�l���a"�Bڔ<��H��4<t6�
�VQ�=#�U�q�Zu��̨ȣ�u�G����I�o�5TI��!K>�T���ʶ��.]�ځ��eG�`��~q�_UH�-�����\�0��#��n�t%���"
?O��Xu�ҽ"6&��"x	Y��ȿ��g��P\��$��[k�h�c������ӡ�ګ���5T�)_�1_d"uB�a�@m��!�_�B⠪��ɴ%��Sⲅ�I�*�Գ���]����8z-����ݝ�����f�KQ0Ydh��w�*p��̬s4�ȋH��؝�a�#�#
�'���a?r��R�cx�����Ԭ�AG�����9̵�}uq��\��6�7n�6G�T��m'�l2⽩��S�����F��q�"D@�

�"b���ܫ�-���V�z=+D
����a�瘟ؓ�#Mw� B,;ֹ��Qv�DT姛�_p 49�b�ON�T]�v��q���8P�X��K�͢��%s�h�%��@�]@)25���E��ό��!�uԮ��"���9����Ǒ�VaC�&ܢ8�V����y��	�!ͳ�+�Q���� �H��:��.`��ZV.vdm������Ԭ�Y���aGZ�!�d��*��i���$�ٲ3�_^;-���M�^8��?%�k�r�#B��ĕ�ڵ�K�GU�\����~���m~6�ٙ� Լ�j_Lh�~����Љhi`a/c�+5Dh	D?����{�(����FRϲW�������,�x�K�Q�]m5I����si=瘿�FdEC����S꫈=�5�:�tH3/�݀�L]5�ޱԩ��m�b`��E=���]�����إ͒RA���ũ�?ݣ��^��PC�1���yB!�J�.��Nuh�o�%H,�[8��m���M������]�'����'��� !��J���X܉�jT��뙓MF��]aDt0����z^��9��è� 9��y1X���Y
nr&i��e����� VpJ��k�1���7��w^��*�ہ󿍬��4�����6r�1Rz�	ktЇ�&A�?�H��v ��Y��O+,���C2J�q�y^����ѦNq����.�2�B��=� �W�w�%n�������\��TנFN���(�5�\r�[�$����q��A�1��6��+*��k�0���f}��Ro������d�� ^�*F��4�l9�0~��2{�MVnsT�[+�d��?�B����x�.���5�%>��d�2� �T����:NͲ��ا�yDF�s�m�m����Q��+N�ㄱ��Wۄ�D��D���U���C�힇�f����)M�����w�h�IOƥ��T���آ���
A1�Y�����L�Y��jp�J�V�k�*�c {|
?}�}zƥ�y�1���	f�w����Ɖ��Ae��y� }]��%��;fGޣ(��_��|������r�U�gϏ{���>88�դJ���������j�M[��1a�uRr4ȡ�v|c+�>��48��/��,M=e+3V@D&\ae��ZM�J4�� M�R���"Rl��"iNٳ�+��fML�+�,�/	���bv������^ٞ�$Q�li:�g� �-�	zJժ�$���3�����lcT�Ń���!
�����;�Z����Lk3} !��D�B{�����kg�{�;�5W ���}/O����I�B�rt�w[g;_#*��zY��M�g!u��y���õ�Tj�0ϩ�!�)�F�)���<DI"<H$9\[:��/��y?DR
\�S<M�xd
F���]�"��Y��$���=�8`�nϩ��_uF�>�9�sߏ�����nn�~��� P��T��j�z��D5=k&�J�Q.�YP����J|̡����t�,J�yW��Xb�Q.�!
�&�3�Gi�_x�	�D������s�����4j���.G���E��j��"$]���O�&^N'y��*�v2�K$�5��������u+Œ�k�r�l^�f(����E�^p�=�쭯�V�S�N#�\��D,��i�~����T�-_�LM�O?�/��8�Dcv\�������ҧ�*!�KN�^�QO���Tnd�f?o�8��=�|w5�r���2}�?Ѫ��A��<�R�%��gpW%�O��c}�Q.!��(L���?����R-?�(<u\E~>׼wN���۩�%C�U�=ͳB�"�ZzJ!#n�(�z�0�ܟ
�dZA��dB?s��[�/�Q,&���E*W˗bw5{�|�9/W�����Os�m�N�4ʵ�x�k�_��)ݠ�-6��uS�mAKV1���n���}�R?�0�����M1�E��>�Hډϳ<U�:�=q�y����0x	�!�ШR�	D���|;�4¨��#L=h�:�]�k��l���r�;_�@�}n�M�*�Z�1=�)��2���]��	��sb�0���tT�1T��rd�l'�L�D�� t�?-�+{�8������|���/ �cȂl�n?9�V�(��Th	�
��sφH�GT���bu�������u��a��3�H�x�vI͸"��]U�UM6tF����0 �9��hX)��vId�V��7$����?Db>y+�3y#��[���9���އJ�ьǬ ?;#��!�'�������K��?��i��O��.z*,B]�_H�R��8ŋ�.��Uiμ����rԒ�K��fKOO�{��S���%���m�����5�F�TH��S� �%䚙�3�x9}��&����a������X���R�`��1|������^�{�4=-��?E��;�J	�,��o248闎�0�|��q�z��[���WA��q�����	�9 �X�loC����_��NI]�й�c�͎SG�i��!�$}��E2?��h��O8ҥ��K�Ḁ��>:|�(`�-�T���ZU�]���]�y�������b��O�X��P*{\c'��}��3�@��Z^."8���?:zӵ�3�#Z��o?~�>�~'!EUzL 4���p~�s�i����\x�����p��'i M�)}uj1d�a���3G��̫T�: c)r����
e7�^b��GJL� :�S�$�&�+N��,Z�z�b�iqS�٨�Q��m��C��?�u(�tG�8��#^#�
�UE8�`p�vy�-�Ev���U��e��2VU�ٿ����$��CTH%J���k�s�q���x�z�B� % }^Ǹ�{���T��)��b�W�"�<`������0X@��@��T�bU�s^TC��c�'�l� �9��	�m���oBDYgk�q�����s�*��	�1$ub�@/�N�R+I����ziRϬ]͗� �
=9�0�dI����b��,U��mʶ�3�QY����2̩?1�,~e��~~����f�_��io�ЂI`�'2̾�F��1\�ʞ����mC�ՠ��h�O�ϔJ�.� U�=j�����on2�B�t�e��m�[u�����̙Ef�XB?�~�4�r��߷G3���[N�g�E�0j����hQA5�av�?�*�������e#t���������6��ʕ$2�&E:0�9R%�5u�{2S,���q��K����l1Gt
ղ=+zD�t��p<����5���ӯH<��{C���5��e6�Yn�`�藛YA���ܡ�����v�j�|-���@HW�T���y�Ǿ�'���AC��/=�
���Z��(�,n���̓0�kp�!�1��Y͘t���~{���3ơ��1ڐ�7����"V׿+'�!2��	 f�*ϔ����a���X������ٚ������������ʿ=_���O,��V	��~į����q�!l���bH68p�7��6�J"�;�N��]ݷ��IK)�]��{-���C=r��eI�h�ʼJ�u���ި��C��/}�A�X7ɞ>�6)�-q��B��s||����ѧ�<tB/M���ze��T8����?I�T�J{�ؕw���`�"�2+㝉n��Y7\�>7��x6gc@Y%�5d�Ŷ��du)���N� i��R6P�6��'`��r��~A��O�x��~�fT�
_[�ܨD{g�NvB�6�ւ��m]oK�6�|w���¿��CQs�j(ğ�뫢b������ �+��T�:m�S�*Y_&rL0���ѝy=��$��*�!H��x��G���O�r�ɕ�s�)5#����T�b�^UW���������I�z1�xTZ�]��z�怂IJ������g	x�j�S�-~R �Xn&�u�Zw��t�F��t4���.&9*�5m9�dX�n���hCX>�垁\�	R֥ ��a)Џ�R�:�t%Z R��d�2wC;��ʽM�Lt8)���R��
�.������~�,��Y�� +�H�T�n���b�JA���Zâ�L�U�&��Z}y Z���/���h�(��;���=�7�zF�u�$�L\3��/ǅ-��j���3���ڛm}�y{@�4{�.D�B�l��N�(� ����jr`�����8.�:�hp�7
9�<��[�_~�x���Q������Xĭ���_\���QP$�H�}̀}K���NE�<���ӳ8n�ެ<�5�ʿVw�R�㥢v ��9�G���.��h�
�)��:�1j�@N3���!y��3��<�v��Wy�;��r���֒�#�q��$�\R��7I.����Ws�G~k�5>&�㷈���������sʬW�XW]Ux���� ;2#�J'�bXڼ�t@��k��\n�-Y����D��G�kd�}v�4�=�;�n��z�l>ꯅo��x{9����lłir�LL`w�H3Y���cD��SV���Az��*GGO��1��U<;B� <����C�*BE�4��F����(����*~����|����D�@�s	~����.�\���g��V���?x�ĩ!#��D���U�?�6>U�մ+w
���eժ��������c�|l�S��,�f(�{ܮ�C��Q`��p(�ɝӯ�H
�]
j�9Dny
�<9*Xl8��l�ƺR�&$_'�WJk3\V R|�������x:=��蝱3HֲX���:� �R%Q��f��P�f����rS�#l�҂��Ҭ�ܣ�\tw��Ĝ*�@8M]z'=�R��o]�<ܠ��m|vۑ��HX%:1 �����������rx�}F�"�U�IC�4��
`�j�����I	8���Fk�}�:������/ͽ%��Ƀĉ�%��\WV�a�[�(��x���[�	��07�O�C�݂1R��M�i!�
���1�� 7�o"Ϣ%0�����Ϯ�hT�$���G�5X`E�,P�r�d��2w'���,�t:�c>�u�^�Ǐ��R���V`��U����>j�����m?�a���pl��B�Q�O�oy~���>>�}~��ښ���~��;����ځ�2����[3Z��R��(��7}y��>ߞ�P� �GP&Y!m
��n��3H����c*� ���(@�i���{.6~����Ŷ���Yo�����.d(|m/h9��6O�c�=]� �ZӋ�T�F���I�ϲo�
6��R��!i���=�2�%�n��9��:Ωz�6�8��m�sֽ�p��7sijO����cU��/?�}dX��"��p�sF�Q�wB�T��Z�f���x���Sk�^�s�|yD��j�*5`}կ�BG˓j��!:�ա�7�4PHB��`�]I#(b�BS�q�}��f�V�ܝ��K�Y)�Ǯ���El;��\mU�6d�,v����ej������ ������)�R�����@��<�yc�p���s�;�^�J�O�Al�er����[���*+�Y��'ַ"0?���Y9e8��[�t0�#�`*)=���7Az�HM~�k�)��U,�vXи�Xc K�Z���}$�^�z�TM�R�^7�'�-1�F�P��팟�Տ�
�b��3���.��6�Q�� �ȫs��Z��b�������0�����Iy���s�f~�^f��������0j�[�O�� �����8.��*�]�dp�[/��/��Fx������"��EpD�EA�ɚ�o�{4���W���Jb[~M��` F�ssk���^��CA)	ڦ�\yh��̟IV���܀�z�Kf!�h�44���b��-a�T�5�����'�k!F��vr��	L}�I�-�͑�8�|'H,����>쇡-ٵ`�YX��������#w*�w�yФ$�}�͘�j�ޯ�����>-�@#7ޯM��B�����͢�E��D�`kԪzI���/���T��h8�U�E��,��ӝ���Z��jߺ��X���/S��υq�L�ē��v]k�g�_�ށ�R��Vùܗ�ݺ�Ss��*���ròxUM�\ˑ�}��	;)>�B՟���n�D	/�[݇B�M==/�ʆuz-����D�0�X��98�=S�Y4�"Pb`��7+�v�|2�y����C����}���Wg�uAb��ں��R�̭4B�7;�@C����qO}{	���Z�M��}Z2X�v�s��(��:��Ne�f�$ry1�%��o�E����2꓌{6��.L��t����/*��(�<�lh��$$���� ;�MVQ�^� yd�h���"my�<{<1��<�� zn��0x�|����p� b0�C{%��f�z���P_CMX(xC>;�۹9|K�
F-�H���{�����k�����]AO��!�yҫ��47dnSh'�������l7��5��.�5���ܽ��g������s���vV�����y���$����?s7aS�����TZ�\$>�&ԧXC�CL��;J�B�ϸ0wK������+� q�t.C0$���z����aW+�s78g1����?�����q �}$�S.N�W���y��K͜��_�LA�}-��í�Ȋ��t|�uN����
����aNG��t��M�i��t9����:��@�b�x���6�gOߠ��F��0y�?��NS6�H& #�������ˑQ?#Lp���P�:� ��Ś��=�O��ɳ46H�H��bQU��Z)*r�uZ��V�q[+0���g�1���X�ˉ�-Ćdk/ht����l{~�}�cܧHmg���7B3F˸�ё,tX�<DCFЋ%��XF
?p}���]z."[@G��R%B����q>����W ��ӔXFKݩ��i	L6�7^뼃��􊄫�NHqq��e�~�s�	���DMܷ���ʖ�� (J���I�2�}i�Q�aIt�T��P�u���� S%Z�YN�q��{dn�A�;ಛ��}�UD�tW3�1(>�T#�1ۓ�U[���>8-r�L5��^^�ݑ���c�N��o��~p!xz��Q�fMvkht�T<r�ȵY[^UM��ʴ���~��^���	58�'����~:f��K�d˼0c�g7n��r�.`�����\��ʦFbo�+a<4˖ڸf��s��4���1#.%����m�m�c�QPra߳UU8�����G}J�|H��U՚��˺*��`D��ך�O�߃w���a����_}nѸ)��w2��W�������:�	$�\CwK=��[�t}��U����cy�fA����ym����>[~8z{k8�ם�{��W����{�S�VA ��#zw��9;#���;��F��hC��k=\��[�n,�EB�C{-@���R��\C�G�����Qǻ;��RN۶�L�u�q����ЬL<����Y`ɳv�_r��@
�)��H�8�Ⱥ��
����(�,ш��dD�<,wi�^R���Cl����+��s�ξuT��Ǣ�Ml����4N��EԴ�$�,h�W�KS��1�!ѝ�	C��.Dg��]Q~��{~I�1���E�`��i�^�Ks�6-y�g��m�?-�S)Ǌ��	˻��\_����}��y�ۗ�5fS�s=�<U�����m夎�
�m�0�Y��=U��*$y\B'p�J�@�\�N^i�E����&��O�4Pє��RX^s�~��q��,'��|��� �U<7�-T��K���4)�a
�7֭{[��o��f�E�7�c�!@�G����Џ��\$�l�N-� ���9pb��]��Z�v����F���<H\/x�1
i0C�'G?�P|X�͠�A,���F���-4(��90g�~���}vm7�*A4H8R\&\�3��.asMd�fT ����n�J�1���J�u~���o��2jD�{둾)�F���I7
�C�J���GUU8":��Xk�4T�-扌�k�FSȽC���I>��d2��{��/���Bw�U�P�Q�A?�zE����<%�Hn� 6��e�c�̔����1�L���ߐ@�mj��e��t��D���N�ξ	�tAfc��2�s�g�5�D���yL.����L�J���f^>z�l��hTIF�������'��7��Zͨ��fB��=1rn?k=�d����v���q�4���}Z1�[RZ��ơ�,q�#,6C��N]Ml��}e����K#a�ާ��;5DV:��@�,�o$��2�� N�o�+�9l���9���}�+}I��,�+�\�/a0?f��k���t,>�Kp�Ly�E�n�S�fH�)a���-���Z�h�i(��w��aS�K,_�`8�)�O��G%|ҳ���ǉˤ�Ś2���x�Y��ϛ�D7b[Zói~����`�0|�@����q)��n+ffpp$��P�ן�F�sNP���o������i(�H�O�]�>�K`�j�;si������ל�f5��{5ę	��_��P��v���m�%�,i+�a�1/Щh�6#<�]���b}�Ɯ3&x�Wi�X�Ȇ{�O�3�N�j�U�qo�X(�aɝs�E}D�R��#�{�M*vR2̢T�V4.��0�ݩ9�fS�2��
�E�6d��#��������5��9�*�D%����2�e�R�!�|��E@�;�l���֓�A�~��WUhY���w�ײjA��6X<N�����9+�N��UU��x��Y'�}�a�ϼ�:��Ƙ@���s4��C�1 ��kk����`9Ƿ?�:t3p��X�;�+�ͅ�'�����T6�3�~�))��E��A�"g_�qz���r �C��_c�)ˋ����=K�f�kD����Rp`o_X� �w�Z]�di[Q�_.��R]���&Kh�Ǹ46��s	��%8��<e��_�8�%Y|�M)o@��w7f������C��p��dK�����B��uǦ���Ǹ�.R
^�~l=s]8��U�J;����/a�*곪�NJ�]^���U����ho�n%�YGwWq*�pu&�0yN�l�S�C�$��j{���SG��>7���z���׌zH��-�]Q�PP�X�S��Kc�V�J	�x(E"و	�H�O���/7�"<O�sm�u����[/`DNs2�Q�F
 ?VU�[��7�
 ��({aR�P�^��6�&|���*�v(
)���"��6[��Vǐ�+�� 	��{4k����k"xvݬ`a^٘�ሖx�[�k��m}g�J�s�Y�F����6q����H ����RM�8S����`�Υ�mi�5�3af�Aܫ��|ɔb��S`W	��"���+;/�_���QZ��������aٙ10%'��"�T�m�m���$Έ~�����??�j-�d��\v^m*��E��}LK7�n?R�=�j�%��k��(A�c�c�k	`�ӟ��3��������������?η�r�dX�t�r{����Q��u�c{l�1�"����aw�~��Iw��XB���.s���CV�0=n�o�_Q��쯹Ax�'��*|���~����A�p��(�����/;|�@�F���>g+�k���?��V���`ےԢ��b�'��K�qj�r��p!��F�ԙ%T�'��E�\��*Wh@���$�3���s.�JB�{b*7iy�������]@v�I�I*�K�C�����r���F��Gr1�����a@G�W��] �[I5����8��K,i�V?�J��,��Ωh�Cdo��HI�}���0_�pq?ܵ�*�:�ۇ�i,9����o��v��|ﲮ��������O6(*����/�X>E���Y@�V��u� �cS.�:Ke>��蜃O��,��T���G�K��<��[�X8$ƞ�-�2���.�T�5�ĚW��=�SyO�\�������_����L$�^�Z���Ӊ泋�0�+�*?���p�Ҧg���=?
����+�K 6	0���J�(y��X<��튿�޿{#�G�i1b�²��\�n��/�!`Â�]�_��DRA��u&5.4���E)+R���ҷ�EN�X�����B��v
�pG4�S3�n�m8���������U���i)���P:H/h�w�'J �"�/X)�F�~#w��~��J�%�#:�$>V�Af��]C��>3^��ֿ��P4�q�F�\ɫm��@��U$�Ӹ��B<]Jq�9ĩb�#C���5ݢ��FU�Q�(�)7Uk��&��D��:;'Ȧ)Qtc^O�رNBdC�����x��3�����p$�Z����MKoń��%���P�����oz)��������c��F��·� %�x|�m��R��J���а�)���΁;4�u�+H��[�F�<!��֒(�-w�S�Á�Nɾ�g���~�-���#yT;��P�rP����o������ o��s���BM���ح��A[} P�GD�#�/��p� |W�S��8T�.�Un���{?���1P�5y��?{U�%-�Īt>��N$�1yˤ�ӎjeg�S�l�v�����%0q��h�fT��<'M� ��]9x��3��o��� 3y��4o;B#�7'�S�bW�,!Y-+�/�>)�;u{��\���Mظ�4'ø���:P����fYv;f5#*�t~�nz���������B�L��~?aX�Q��&Z@@�$��ձ�b�[W8q�{�x���,�S!�t�@h��ɾ��!C: �R�X�VNe\�Ɉ���?�5��,��!�e!-:�x���3�GPy5I,1S�N]d�p�r����8N�;e�,U<7�X���6��P�������`=8��#1@Rc��մ��`��?����"h�KSF_M5h�y�$g��=Jz���HmI��ЕE벑W�/]K����#�iJLyQ9�2Y���.�����-�i�g�۪����!*�G����Ȼ:>�D��
y����-|�#�Μ��f ��(D<����������-���dj8�l��-�4��3X�Y�+s�@�@X�r�7�nCI��Z����v7���\q�ds�]��?��R�F�����F>U�@����kӂJ�_-ϕg��$�.���6�	�����sP׽������|#�6c �q�ˌҍ��+i+'gd5�>��i+�t�JFn@��X��ҕ8�)ĺO��V�LOj?��(͸���>l�g�*�.QX��Yu��ԧX�����/0�3��N��]�2Տd�&k�-��s/��膞d%�����Ĝ�"��'��8޵���	�>�#za�V.�+ފ�&B�� �#�0"��B��IVP��
2Ӱ�
,��.�Ŏte��~>�z_�˙4u��$�:�\l�5vy������.���u(
1Lx���m���XU�B�o�Ě�H�R�	��.�&��)�9��K���}zA�w�6VAm�1)�*������Nh�M�������nѴ{*b�8u�s�W����T��)�D�J�mƆ��-�͇TQP}U�u�6�x^�̎9�����6�M���Ev�f�@k�/�ȿ���{N�4�|���鍰v`�Ţ�
¾�;;�aCl�K�p���}G��G�CI�-�	�;mSW���Lu\LA�!H"1��:@�l&2f�t�t��H�Zq��2=�l�c��XF��'Z�
�*��(|����C�U�d	�"��~�\��Pk�����1�lJ� L2 AR,�ڱ򝃤��rj� �:>)e��&��L�و;��7�N%L�:�����q���(5�K�(�fv� 3Lyv�D��&�W^.�?�Ұ�N��qj1�R���<S�"��TZF@(�\�H��h���:q�R/���������"�n�Rަ���b!����|l��9��!e<9'e���.�Cg�}q6�i���ܐٙA�^�4Y�V�[5V����WՐ>_�+{mt�� }��8(��u�:1����p�v���G�K>��Iy(����`8*�ح2B��eg��!�l������#LJ�
G�b��תS��<�H?ᆤ������P��hE�3g�ut�s�KI'ڋk�X!癧`��7xb���n����Ai���D��~��tw��V��j�ַ3Bcm�8G���B�Qbw7�U��IUXQ#|�
����7�!a��۠%�z�1��c���ҷ�{���!�D��	��/��j�p�&n����C3���}���y�a�x��5���< 賏{���t_��G"���y�D��[��s��Y*'E�q��nn�Q��1�o���&�7ʡ{����1��b\ҿ_�f�e����K�����[H�r 9z%��5r�$�M��
	�j�1��7���Kfxc��/�$ݒ�d�����$6|ɚ�|&w�F��^�f�F��q�n��2�/C^�����������/fܣ 'Od���ݣ����#Z���_�j�)h8��g�Wx��Rk֞k�ף�J��s�U�.�x��u���\��Q�x S��4�%� l+]�Ijv1`M�_V��'P{Z%*��8��ي�C��J���z{��Yn`�E�g@�d���
�=H�9��=��%��
�����1d�i[���?�	� ��qn/�-a��Bn��QO�����8��66DY�i�F��{b�q0��:u�_j�[��E��&�nd���:n��R[�p}PS���v,�?�X=���Mm8�١e�c�[��\�b�(���|��<YX=��8ڝ��Ռ�C�i�6"��%��3Or��$�s�c��s�N��`D�jj\�Fp&F�%�ʄ�wPk)��0���1���Aʹ[�aW;>������"�L�uM N�F�Y�L�z��F�aX&���}^���5� ������	U�+��sB.��U����ڸ�����8s\�6���ċDNZ�ص�MO��ܴ��hK��h���U��Ϥ󔈽Ɔ鐎���A�F��_��&yG�6[k��_,T4u��g #4F#ʛ�>�����O�2���):�~5� �pP�"��%��㽯oUW��I�s���� h��
���+.h��Ц+a8>���ҿi�"�-F̗�2���.g�U�>��+�~��Z.	���H���K���dǲ���O�Q�C��.0ɰmSV:B�d�q���	=i�����׿��̔1\/�2���vU����dzug	n�������0Ya���#��f/?R5�K�W��(�����c��b�<bɓ���0�E|]�Z�콼f�k$�!bMr�]����3'`c����*�%��	m�~�:��������7�x;���{�i]	�i�;̆e|7M�dttM���~HQz������~w�����o�KY����P�t�g=\Ю���S��s�-��ݐK~o��3i��985= Rl*s<�څ�s9���2i����vF��ff3�$���Yj;�̓*�x���ޑP�I����F I�#��d'�-���C�s���\o�̙.f�����x�_�$G�d��)�̣���9d���;hFZy��N����M������
c��F{\�����C��=5Z2Q�n����l/�ەtkS��� �JK�[��f��l�>�10��J�2�y��Z���rTSk�+�²�����j���Ao�<���O�f+4s�	#�a��}ql �2N+�1�N��7lb�o������3�&J֋DPʮ�t�J����y�W%;"-^��ۼ%n49��V��ϊ,e^��gR��a׮��H֠��7����S��%	6��nF����u#��o��G3�}<|�y�������3I��Y<��-�-V���_9M�����tK�+�g�����Iw�AU��>��qәY�݌����5ll&��=4��o�ʃ��*�C�'u�>f�s�z"l�L[��=`�§�x�̝�o=E����A��_�E��B_%I
,�[�� �#<�u�����E��k�SS�'K�����~����'��?<9'eG�l����l��嘞6��
x^��@���}�����0����^PQ����R�ڐw*U���/4����(/Q��(����
҆i�ݹ�S���I�)R�z�x۱>X=�f8m�����})�1Ǡ�$�����܌���"dx����I�2�NfX
4*����)��h �v�9�*�6z���;q���!�Y�z�/O�PыC�W��Yo���w�tUI� ��;�#^	�Y�*촇�e��	�����ړ�f����%��_r�/a�ګ�98eD�X)'�ȡ����j`7��/N�+jUA�@��\e<�H?�kP|<֡V�^UL�r??�Օ�Z�����qG��{��~�l��6���i�GS���8Q�s6eU���i��x����]LV��\@	�(-�Nl�D-��NEIo0e+h<��t	� Wl��A�J2?Dl������9m��>6��_�hX�Q�,�ȍt_p��`yVG��Й�*���X�N׷\��>�Z���&�Մ0&�\xTk��9e��*-D�Q��U	���j�z����E�o��D�Q{Q��3��Ggم�M���))���؝tv��I�X��9�o
�[�Í�#³�^[N�CM��~5I��M&W�M;>V�?�S����D��=E�*gZ5j�o�e�k���G��+:��:f��0�u/'�ø�bڳ�����ȍ�
� ��>!���k��.�²R[��~\��B\�>y�C�'��b�7X���z�{Nl�*��T����7`~�u��������~B�|�Xl�T	�KY{@��q�`�bNbo�!`Z����gY�8�j��u<�?E3.�3V�����̼u������m.Sw��;��L\6Z6����2��H���l)R�����[|p��y(��ߺ�B�(AI,D�n�o)����lLk�۰Tv��$�֞)헑c�9�[׳@��O��CT�� ��yk��w�s�_�n��|�<���9<c�%1�؏I�,0d�$����c��<X�`��_�d�����'/M�XKA��)��CЄ����\�y�D_`���_]iF*�@��c��ǰc�����R��lz|g��E����ɹo�W�m���f�\N�6�6	�$^+M#��(�J1j��}xo�!����),q��Gg�]l�QL��3U������%�k�~��eZry`1�t6�^a�r#��������_��$0Z�z)~��1�H{R5ȟ��[nkf����\?5R�#58Ee���LM�U3D��]���	*W���r�Rڊ��D��E�OB�ޯ������)��#c��9�}�Xg�ʉ�2U�E�%�%��%Deq*�>�����M���������8�[#��#bd����M-�&��p�a^�!��A�ՆZ��~�J�4�{j�� <��"c�eH�J�?�Cdg�ˊLv,����o~!�6v��ɀ���5��]^�
�N���5s�>>���i��cG6������B���`Kd_�^�B
�Y��s��fQ�!�?H�-��PĊ���	��k^���?sh�'�͗�x�*٤�C[r��0�4�z5�"�i�]��9��.�z��slAiB�f6�|7���JV���N�냄 ���&�Rj]�� E����֟l��GJj�q��ާ�dU�%�z��qv�&��ꄿ�\_�U*Wp�x�` �Aa��dZ��zD�{��m��[��c�8��״p'�ݲ��;��b2)Y3F�j�5L�R1�n\��!@:C� ��u-Cw�f����{�����@??��qW�,�� �i|�	6t��J�CC��ÙDc`ڄ	*��2D�^�Q)p;Er���4������?���N%\�)�*t�x�k�G\~Jm"�h��eP��P��ߞj5��MA�H���6;9�=���HvXQ+;�FP�7P"#׻u�$�2�ɡ@���g�
�?�.�b��l�Q?��Pz;���t��9�B-�kuc;�^�����	aI}��?�R늄�Q�����C|:z%��F�lpci�ANĈ�~}��\t#������Gk�%�S 4�C0g�;�N��b6���]$�!X�;�6��7|$nՎ�<�l���OS�<O�ឝu��Xk�k:��2|��:�.��mK.��B�r�ը]A����l���B ����&K5I�Gb��)��X=	/m�H��bp������Ɏ2��Q��ǨlZͿ�@+hJum���N�m{�