////////////////////////////////////////////////////////////////////////
////
//// This file has been generated the 2020/07/30 - 18:15:51.
//// This file can be used with intel tools.
//// This file is intended to target intel FPGAs.
//// DRM HDK VERSION 4.2.1.0.
//// DRM VERSION 4.2.1.
////
////////////////////////////////////////////////////////////////////////

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Intel Corporation", key_keyname="Intel-FPGA-Quartus-RSA-1", key_method="rsa"
`pragma protect key_block
HJPAKd9x1fIRFcYv9A5u7az01GcFAMc7HFumMasEx1k9G1hhQNg3RusEhHqpnjcObShGEzLEJ+3W
OIDdL7fLbb1IFn/iKVeP3vRimfTuiZJsiZ88tLVnCCqCMU9J8wW0SwBda5JWCO008m9cbMNru+L3
VTdz3g3MzqwMo2cVYhSBmOttxfG7S8kEOt9pEy+6c806KxZu5jrQGBzDNvYjZVgxOjDpp99zRayV
chmu7ZSIpDH1cDQU/XliN+cx5IuEYJEK/YCf2ToMEb5EX//PmyVuRFg93Gv0nK0eajub4rGJBmsN
ux7lEFvNZUyyU2FQCItQjdWcQ7X2f9i+7YsvJw==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=20096)
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
VRTud+86yc2VArmTzB2voaXGVnzXCWSz6b5KcxNRjtWVSMuXh58fNAI37DEQVGCpsZ8aR3OotyuE
1Ju+Af0NUl1FWGdr3g8oH9PGaASj0EFcqmYMR0rD6Oj6YXGtDGHgpl+RdBf97v6dALRc8tzzHRPG
PFiA6bnh8GdmqQmrLGKOhfg+GBAjsyDkARDkNHR9IWRW/6AJz6JQQO3CarZldy0TkMl3u6fzRcF9
AhOQ9dN2fvvf+B7TJExf8opMD+eB1OwtXLa8qvq3zQVzHbIHmvjw+3tP58HR4YiXSnXFzaIfEjhZ
IA42pHvQnO+w3TExkdr3hITmWdgGPvmcR8HF1obUYkMpiKOzQ7ztV3LkOeXirwe70XHNcgGb0ree
CC3b+lLfYajnXqoVCFj6xzcnMh2gA+Yh7cAH/wsziaISZPxbSIYjeaoMhMsVT0qe5j/jY+8Gu0y2
EyGfh5lK20B6kvNKVa8jD2qv+Z+98BzaP5KrEit/RXRl73PiP1bXlkSQkNhH1iKWl08ZMdH140ah
l7W3j53ugc0pcnRWtaJ57cw+OOCsvc5X6AsiGqoGbVzBdRW1+MSyYep5Kj8kBp1JlRnjkGenSc1x
Rn2aGl9S5ctYYbCbNeEVK4E2gSGneVLvaIZxN7nQ+mAQ2+AJFIQ3EPwlRlaR6hjJhHm97ULYT547
b4ZiM3916AUT8aSBbYHqMl+P/vG/74DFZ6rthvoHj2sa6MSV8vVyOhu8HOWD9jews3egCU4aKWFo
E/UgHINgy2Vl0kX5KULft7Yy855DnfyLHfvS7CYwnzDTK8RPyUdU4sF2n4EYKA2lF/T1qgu12Ggu
bPr8QryBMFVu4ZbPx+e5N1Q2S8HRP11ckhFc1+q6I9yqQSl6LVfCL+AOr4CpRhMgCsZs8nKwSYgX
EtOjBGMb3PiwNsKYcZyDUPfGbG8+U9hoU62kqCy7rtaZbu+9up9Slg9wGV2v5J3wyIko0bdP05O8
5E0+1UeDa/5LRZprAgmvMCnuvw57UBzcj2/YVa6uuKqFuPE5T67/X5rl3ekdP0T28y5G0yS5N3xc
gHpmKrNKGet5TVfcOYN6rK+47ZAtBBr24/F31zxq2iQ1Oo9L62MQfhHXIoIFogVkhodV/MsXBXmJ
CLCljwWhSAtLPz0cud4HWJAQcOFngJSuyHCrQsAF3No0NPizmcznaP8mRYeDQGD3isUvX4PNTBLS
xW2brZRiShBQwgzWf5wIJjQP+3N0Jl1wl/phzMNEXxbxl9tOWLlguR/whRrucP01HN2BCuXBo913
jcb5L1N7cbaUF1+2fS3/10Sr3O/ueCXJgBSVvH+Y7y4Q8UzUX86we+A0ts183Z10UblT9g8hBGpG
BqwN0FbDnZuiDccwXZEMGm4JB2Cr2x6HHBz26nMfeiwPd8yiGR/gEk/4l5cc9JVGPSgdyj/s/U7/
35Nvcu+clETcMepVkEUMD9SPJrZJ4mKsUK/p19h59esCgLPn2vvjStSW2yLmZUhI6hHlPpu+rKBW
KOaZi8cAthtZr/BC1nIsUG93PYGrRLF2hmuBqxIFHtSVMGLXb92w/xhHEswsQzl3MiqeVEtNMaZ5
0g/ynjxAk6Cs5AY5QVCQp06x1Ewy1tb3cCEEEBPzWTcbTBaoU0u3VZCPk1Mqwrh/kX1HNFyGqzQ4
iRE3pG7/gieQUGB7c8GaSpOKQtcNYUS2KwLZ4JUuL0PtrYi33xExvopL/Z0rldVovaAjOvDhz3tL
KUKOc3BUg4Y170C9VHc7zV+Kmxcsln2sYAkpBOfofgXWuUvpohiBJOCbjYlf41fwGezQmrGFiy/b
bny905MyUgVI2YoJwQBP3Ls3oXKSrSwhVIiaiAG254kgmqVimKwNvO088a7qSn/K7p9LWZQMEmcM
0m2ltFnJDRKzt25lh8eIh97EvZHzQhAlc8N+C9n2gEfB+zYfzXv3XAynwq56tg32mJe/t21xRQO7
9PEOZC4b81w2z4Ny8aV9Qjw4e7dPByOtbcDcIXXr8IAxk5g/Bq3CoXSa4TxQAnjmeRhiiNxFZUqb
BHaMXmEeJDRuDfcHoYzmaXOyLm8i1lZivHspeHOXMb4lRfsFOXNdtERKVTlSANS5HUVS5SEJGC0s
UvuxOWMWWkHpO+PvVXQ2CbbsDFUw934Rtv7cyKWdBIRSHUaGk4BxnnLbzfi4S+3rnlTMc97nOF/B
YMDN/MXmKc973q55lbI1ql7y2hFr+T/hZNiT1/eDTZPyQY4PbB3Topzv+i/G9K7UWq2tOqorCE02
fV80oiXcrgUxPhiKH71QY4uy0dy2aByGElllF/uj0LkyqWU4EdgqcPO9uhG81HDxA0EMxhfSjELm
lY0T4CM734Jvi7Lfi2SLSwndNTUX4VzZTAhuBnUbQV/d/fjr3as6ePj6wLi/IpetVk49zl4HgKrI
YQWjw/Q+st9J9h200LobSsGxLxKGSdqOajsXFgys3QfztyUaUfz2I04ReWK11m9F1m6vKOAN4Do+
UeFQPc7QI5by2ANAmCqig1UYlKNzm+E2whh/A+PQ9/y0Ob493gwHt3q4zPL4CTfPF47iE+mSTngj
8YYIvqzQZvCiiohxIfucQT3xCNtg126FXLcNG/t1RFtiC/VuIA+sdr1nIWcEJS76x6IEMdz/oa7Z
V7TkldfyxqgpOq/ZsJOr8RpFVLi/G05kqexZQr63k54N8MMSmrsy0BavEYLkN2nexnZ4wof5kg5Z
CPcsSNU+XV/h88twgxvW/oAsL/Zn/34PDHgmEuYFxQMofKZ3vns5TO3G0Vsp9FEZoBCeBTip+YOs
4Z9lqDXNg0k2u61z7u1Ga4asS5ysxJIiaLOJq0aXviUCqzQuOPaKewJ5iBwJ2NeLogao19MDMGnb
hHCKYBtMz32TevWNz4e4wZEBYXTNPE/Km5fmTqzCRSOryDzH44/dOwvRPCY3WzCOMDO+6gQAQhja
Wx6NbA1QCy96e8MY+bhiOdyT40UzgFpXRKycLdOOBo3dKXE+KkDLiZT0NkP6TOPHa91ar9cnCAX0
Fqi3I1hkugqxYymY/KWbZsLg2krdfFFuHYqZIJqwBD69cdHRmPDHU1b2A1XUQN9Q0720kQuoHWVm
npZXMvEKwtOlG9k6DaBv6ARGl7V5E9sv8NsoR3eU1bnBMjQw4DgN2MVTIKqA0PVSVgD2m8ofo+mn
BYtkgcYiR9T6HsLjS0KH1AQDPmW9kcW9hgJvSKUGEB7YfAbblvOQf68P3KuIBwLLJLMfHbuSOWY1
bR2/H3AZB/PwVlzmKsGY1vzeQtGBWO5WbdSWtvrsydqn1hxHQkn5hHia8nF7quf88HlkMNDa7k6h
WxkPOLZzCNX0yuSU2ULKyM746QnHYnEo0LCQFZvo4xYqnpSAY3Xe1+ms3e1TFDvfTkkThibas/nM
9VkAGPwpHlzoOcF1xpMDoG0s9OVvUhcwvci4Y/6nDhxNHpQyjdzclgukZim4dmxpUApjommtx+2q
N/WdbdfDwu2guh6IXkY4jFE7eDnllE55mEKW5rzu2+BKll6vVSh2oaAsxUVy8nvBBE9KXAEtHNpF
XGuTB3pdbGtdox8nzHQifQI5JM7BDdLOGVTn/aBmASm7AbNCWTPkch/W4ym9M8P7MWjftIydwMve
PL/0DHH4EHICrFBXxWoDspBEkvQaPwnl5MxE0WN6D7ypIzTtFRObALWr3uZE2hEIEOWkNdFwh5r9
iIcqTbmrYc0KWeH34nqxF0AOYXZuLw+HKV9DuI3sHRkSlNvtUW90XqwZfd6MyeUjNyIRw0dXiP7M
dhBG4/FUEeig1x0ECY+nM2InkUbLWjrNkQoy5pBfVftVW/1FPk5pYHHrPFy3nvAVYoUkaTcdajVm
HB1c9Wm/E4Dgzd8fzNAAmzaPGvNk3Fls7ju/yApssEwc71a7jZWprkhsp5ubZXxFlOguVNcEQUXx
gGfJx8VzaQJcFPFPiwnMrxIMM6VWB0YltxpnipxInSNAssb529xF1jr99JF2RF3ugTeAN968Dt0n
rRx8+78YtHbwKeWgUVTa+xbdgHec0tBX+rkoPhxXbf8yaY5Qp7k/B/HdoCsPZeUoc8tDqXYzBYNW
6b2nfw46r76ctqnC8pxxFtXtL4RicN0mn4cYk4/8As5Snl1w+G9/VTg5ujv3zWQ78EQ24y5BSfWr
txVcRE8cK7Hd9q+I6bsWFbH6jn/ffxGk+BwHvz4pXgxw9ySO1gpICEtgP0MtaaJ92bnB+jggYPwD
NYSjAy5enQ4ywrnsev4klN4dySldKTefLGH8+x6eVaC1vG/KNhJUlRfP51GeXdw/bKNmYPD4Xs8m
bT8KmVIHVwZ6UGOQ+g+Y8YA72P7Uiyje0q0OpQKde5oXnv4e8rRkJRCbyRHG5RnUqf54tNcTYQst
7We/xCUaiCBHLhC+sMZ54IcBfgoBbldVqKKipc7nT5lnTzhp320gujHyjXQWnEQagM4l65aEWh7X
OY8olRppZoj60eFqYe+7o/v0/jXdhj7WiVIdQGSkh2TML4Z91Bzyw31UlcLYd40wm2PBZdCDYbOX
+BsLI5HtKM+7V9M6rsiZ5kJtiKSXb72EQaqpPMlFuAQDQS7iVnWX5miLbovEpZxrVQQUhVKDR49b
1TYn4DBwF9/s6FPW036cI6BOoNhAlnybPyMpmzBa4wKdW+X2p1qA2sE3BKW+5x7LgumplGgRGv1d
tSjm9sL3GCnVvuloQJmFzdoiKtttXc/OZJL8nZGbnMPMtLphl/5EvFaOH4/tkdYGYhJ7Lh2bD002
02pLTzKJFZul90fbbqVKKYHC1PA3tkn2hvMiTl4VljO+Rs6T3JZXg5Cf3uflDh337yzKjc/6KbcE
QDQibHn9VxZPrME3N613/bYGzH4HOJlAjkqOEszdIefLGXlThzwAn3Wec5e7tbUc/566xRKlYnfX
dqwU4NOUk/yuphiUGsDp+DZg1RFXvJSZijnf9tqxq8lAX0YqVrHlfPrKJ+Co7UVqyoiiT8ZKG8Pf
Lz2SM/bDOGZeM/sLWuWG2LLqAw6afRkmHwGt20iNE/ItifJFoibDApMTcVJ8m8vOM8BexivRB/EP
ufjsDww1iQsjn10Hy6viJFlCAZeG0OZUJKSnwuxSOe2qzfOkj97xjcT/oQ4UouqNUg9aUe/Mcvkh
sfV9BAeUIkBoqhiFN/iSRuB7wsHV7uGY40A2WAWn0qybaBZj+7A1W0cU/G7XzkFSv8DmitIJ5oHy
2k4EL8AccbtJfeXFICBCLV7ZiEthEAlGhcaJX0OcCCe0r/xtserEU+wmoTiRGpgzC3hQVPsDCk+V
Rew1hhqg6djfkXno0wsaF8BbEmR+36sEZv8nrRRK8mRdtREJOHdbojkQ3ay1IkBDKCTYD+nvpGxQ
bzrESh3UXGly+RouaHo0aFpObAquTg4p/+mwg/gGZCuQrC7Cd8MUbaY/HicHoE+7/b6hM3FyEku6
1hp0Br0p105bulon0L94sAZ9dc7Js4TNExmUtlxMhaELQbyz5ezvpz5JvCdSCcHF1Xgv7v/BCqLh
6gBS1OTBp7zeuLfI9KS/9GwG0GZ29OyDYvX6M++R08X+oiU7cito4DpSqP1j7gsZwEttF5RzSwnJ
mZKdEoD/sU98JScsWM3sf+e2qA3rFmfDdIBn4zhd6/HuHPK66W1GZZIaXkyZ8V6oN0j9MAaE1V09
NHWyIDcKTnN6F4uVJpYUoCcEZOybHX1eOnatCvU/C4FGzAtd+B1N42tCCRd1LNNZn29AoQvyh9SL
tlhmxDrkGnckSqSGzARfNwllXqx0Vn5Kqj8R6FhHUAdk7pNpw7ATeG6UfaoK3Z4cwDnwp8uvJyDx
w3NNb2WQqRTF3WAISfr1j7aq1WtykvFHenEAWvqXXv/SEoei9r1ZSaay1Tw2P3NHxqGpq/v9PHeC
0nQKgsBO1HZxk4pf1488D8Kg1mozowLk7hZMunofKspq3UIOYSHccq6zitEOjRcf2zrHEbDKcSM1
RN4C+s3KTw4+xBo3oBIGp4K3VBXYiUOyCpRfq23JIfnFmW9K+qqzb/SqQj6hat3cGReRly85gkYn
qWhZJpd9YheD5H+max8BibCK8Ii9nHFVZXnTSp5JZyLDRQrNhOPbVTmKOfImiKdADMoGMevSm3dc
Xp6MmJPVbM+UrliyouTFAQWMOUyvQ7Zs2gDkCDUx+x0HXMBFG398PNDefPrNWYdR63rQYnSCLq/g
/a+8/iIa220z6MX70T84GQ2CWNUL/rxqKoSl7a1S4FgGdpK+GFPJDjR8AFXqQGhxP61mMPtX7ge8
AuqIBkWCVP497H0jtSTFRsOOsuHfPHM5h1wBBIMzDD3YiufFJ2pvcqu6rQFvmtU2yPZ49qrIj/OV
J5lj3BjcEpyJuImF1BRDLlzIGGlyjs5EIDSm99QGMlhJAD3PLmz10u9G5CtL7wLOp2x8RokicDqq
Hy2ltWVzmKx8DfG18wkeFMdeOUMqod7rnNvXQIcXkTyzkjADW5mGSQ7BFQv/bGBXYxUKaUROeFnM
YcsX6XuCb8chLP5U8Kx9w2m3OeKEPKqztBHQqb1lmeXTP+Iv3D5XJRcRZYGREkmafj2keV5EnDf4
p0HkDVUGWPbn420iTOiZWdJN0V1aRj8hOvuhDUBhBtXEF0uNiFOelfNNnb+N3Z2z9FElTlYPXcz6
ZYNcPV2f9l0x2jKkwdrlbG1xtfMFQvitp5mlQfZvQv0XJ4/ddMzB7+4IT2HSFkcOKeSe1DGr7wp1
EsXC0VQA8/8WoVzp1w8N0qdgrCt63q2pJ1AfCp4Osd99cPJZuDqSZP9+3NbI0hmj4edyJS2Df+Dq
NxX7bMOJxGBqO7a4QstEk5uvriK3ummK7Uun8qMLd8pMvkdy4yX/jHW5vYJBoHHRkTUkEXmu/uXg
yMKZiGDN0r4dzKBn8TlAdkgNzLm1X8IFdoocaum+sWR4M0crVvxMcriInPfj9PD+9xMgKyG/QZhu
Pfa91jg2b40uMyQQSl0GRj2wN2mOjGZ6QHb4l9jVMf/zj4RxIrFX0gw+eIjOlguMIvvwumjS56sM
xaR4Fcc4RpAJDf/3x8JKYMltAFLypVjxf18sM5ayITV0n3512ignpwtf7WMxfUoiELjaLGo+Y93J
X97+Ml3EOm8ews9/MwU7oQ6vwSC1Zgk0fDdl+Gkf3JMTQm3jaGabvA6M22CCGbq12Q6F/hO+V3Vg
66dNBxDDPB7Id0XwgK+08NE9Z0I65M3hZvp0rwb66g0qf0pG0ZmmGWLJBiLy0vWYc2Pap//vcgRp
lS0FvqAvYce/Z76IGoTcMitiyVux9N88IRMBxwwdpaSziYkhFOFiQo7TWcwXJPJ5J4aQ+g5VOxAR
ddaHYHPx+5obFF/ZpTpahgmNr9EfDeZBheCUrjAtTJC/WYj2wVyAt8OsZ3vlgeqgburH6oE3pa1U
lENGXdHzE6rAhOzXQKUYRU9c/+90LttEA3zbmL1s5rJz4mfkMSc/ny++vyspmPTehQZoZK/Fv8dQ
+krTeP7spW4OpzvrAEeZu5Dfi+CLOkEUa0J6vmCrmPS70Bdgz5t02tPQM6EmxBeXGtl4ZJbxdefG
d2La7OUN4chblDn+lDth+e1JMJRScTgiu8u56RFtv+FriTwupWGVchqUs8kHOiTTLnv+hJLqMyRl
6jVvXbR79TYVx3vqPrRHXeyHCC+xv3G75dBz4m1Ps65A9E8xdgQ4K2gvPhvf7EO5wqjM7KNHtZ3B
95ZGZYceX+cDYUWlw62Fomuo0yFE2MTFtwgmFUkEzdHCNwoOgFbV5AHZJY1nwGBPUmqCR6oxbUQD
ociDtsBqyJpFzAzeq1vHl1FeABSu0YJnsLiLfthNF0AMrjgxTKzCghUXf527Ws2ynmcP1UorwE9+
D0ePsOJ6vobf/D3L5g+DFGhHueMyvUoRcKIWCDZ403QH1NKv2rjltFkUfbef4zyOKXf8LUO1W8hA
laYBcTH3EczYmjbaJP/HHQQsMhvDUh9n0X1ZyzJTMfInNx7mW3rt3PO4FGrGY+VtoOdszBZ8a/6y
t1L69PF3Qy+UOWm3vfN7LnXHiOEq3ZH09AjHRmKsLFHTVt7pGcbdfU+hhrF0U1zqDKpYRms22914
mX0LzTuTCth9IYQvCZsAXrO/gjC0BF5nU6FKwMwEtn89kFv8p5gfxwyuhCB3aP+RMzdIhHMqfxzz
VFAaoQo1k6jVsWDq3KIHBpW6ET+KQGlOcs6G/ql+hRl33Nwos/V7HpWPh7Ypd16hGdrH6lufMz5C
1ScSt3xDLVxQXdI/NECZ+NAFAKkLHIWnXoB8qYCMz03ciWlv/34OiY6Aq1bwQQ9/A34p9lq3XerO
cRkw0JMiPhKK/G3gtTGFC7LbfhV540kFi5JuBfQQx54Ws35CjwkFoPhxHq1vo/z0MX1+Gftt0I+q
gatAEmxnm7DdOK2dA6mlQeNfWAu+7w7CUGRfhzDq5SaPRlYK+cq+/bLatZEk1ZhxqTt40ax69m7b
1LWtPcj7WB7aGvdMLiwn/rXtT5FOZ1NS99NH6sKQZwpB60QI2guTJJxXKHui289EkUmtmuitY6Rw
H6m9hAjtieag4huN2i7UwXrza0/dg+JlbInYOw3vZ3i7mUvr3UeRv9lTB4AdInhzBfWxDK19LPrn
MtlPwD/7g9KMQGGn+gd12HunlXkSkUn/qxkdXKbowGPFo0MKLJQKlliEL9S42MBABAieewrWQQJQ
WSX5wqq4zcIb2Fk79C/4JRtfTy5cYMHYCQzXL+9UfWmxJvLPW9RTGT1V4Cvo131GFK1Z7h21leca
EywJ14eJqafW6cayjWqSfBEtKTwqUCIJvMQcaHng05XxyZwBXkvsCguD0kuqRVsG4ea4aiNhLqCe
LBLjMGgCmxZXCTfkA8ab0XM20FV/BcuYX6Oc6CVdWNqQsS2wnFfWHBJKHfY9kqokb10y95RttlYn
PX2dtgsQmqtp4sx3ZYTKakXYvwUJSbEK+x3RtUQpZ3n6nMjsdUCu+AwhRuOL/s56i0ybuqx93XFT
E9rbgN6jlmCWPVaSr5Q1yrbg3j4lptSkoSyLeuv3PhI7AewNcAPMYlkO9gSHvv+U8QvI84KmqVgA
lKV25jFmiighen8VQZ0WE4bYcnz5yQbo9YOMvNJadYiJ0r2aU6jt2/vyGrujyNrubFDjjlnfngbp
SU7bo4DlFm1xsk4yiiORPjV7SfOCkSR7MO5KDKXqRuaennbx4Hify0Kfq7INF+GwkZS4VR2eAIFt
CG+aN2NPyQ5DtYKWn1dFI5itXsVBRXM92xLV//KMun7YBMcMKp34z+9/H4SFyQ0+iBP4JGEkTtda
FjOUEIiPUccJusk8UlXw6492uNhNdvaLE/xrZ4IfNX5PfTiz4OVpp/OQLlQaIDhcUDxBElRFcLZX
PN9hwbtoQzd5iD0oZqFDVC2R9zObLfek7O0rBbmoogXtLpOqpcZOSmzbv4YXEqpYVLN/AVcoPFg8
f/bK2d67YEoSfHycNUW9yz27yB27CmN4olLnoLHAoEaVP0FYxpMzH6Ik0atOlP7N41+kCJvVGW74
wohqnLYy/k48Oj9/ZfRZcNyT4q1rsku4z3r6cOBOqnUCx9jZTVxVf2xE3vBudgUkyv/aUPKGPNVQ
kZF1XYrTkHEkW/b7qjShtS53Z/xXpJu8c1WKN0HMCtB/9K/fu5i01z59x4R9yHBEWZY745wtuW4A
B2HnvziYlCxQdQ01YCNQqYlh+vSXKmouZQTwj6yHmcF3QNLuCvdUFoDyaUC9q5Gvex19kLwBCOlJ
qakSNT8uAcakxF0Bw0gE+dMWFY9HgO4mOjl5mfDUXq/afbA5tXzc+T0xjNW7suVdvs7dGG73/TWP
4uj9nPtY7ji1dzLNhbydZd7ZCMWpIB2X69rVvXd1I2TZrisTYwGi5GnMrSEjfYl0gUFuEMI+G1jB
nBPuURbk1tR7zox3UmAg+7DJNt12o1Ige8zhzAIYW3by2Gz0Q80HjBduEdufjYuRIleKnNX6XQXm
33BAKYaVtVxuqncEP30xTtQrTzY9WpORUx6h6dUXCaWocW25z8xLU5DxfRSBrTUl3Si6dKFlLvnq
KEMvdtHPw2nsxNVNn4h9iHILl/Rz7rnV2gRCT5pWPlQuoKz38cj7oXxHhjeffBjBrFuZSRdIHHd8
VmJo1JW72lOy8uefwJfPpPlNAw8qDNFFgVp3rLQoumct4omZ1ZAB9YMjU6KCPUW6skjJ1d7cQqHy
Nejqo2Sbol6chUgPsRLSg74f5EpulVte0mntjFve/eWFhYBi71+m0d4GMw4U/flR2389pLMt/Ew1
Z8IOeYaAoZiVO7J7R7veXpVEJoXQ2Xja8mcrXUtw8GRQAASXL02UjSlMIXkxPUELCh5XQ2thge2/
H9rEPQSDvvzW+tK4HzNOnRBqWb7PfFbzGNec0jf2uD06tMRPAwFJ3AA1IjmKrqlLh2GKDbYWOIfu
4HxXMJVO8cGI17NAXFLrWOOXM1vm2pUA9PNZPpFxL1+mm6IM/hnpLHOcXNCTkWo57HR+z70C3HXX
IxPsK270jl5dRFV/SPNilh1gwueyIrNwsOXG1EE6IQy+qj+9yeUxjUuB/0PBVEAuyer0b/Jiv362
zhGifKq125ww3xK3Mu0ZcSYPHCHp9VQacsw5XrhaDoXn4QUB6VQw2ZaeX6gGIzndYuES0CBk5CeP
NPjNmIg+83BTZvuqXwKvA8BT7ewammt8cy7P96Prj0v47LOvoY5dR4k2YfUBiYPYQs3H2ni31bSi
LZdzMxibpr7CJY8yWiKv5dsjcaEdZEmeXCIjWfKJLIIPBrS2FU0S0mEla9xTlKk1TZQv9RkfbTBT
gPKMvfvhzVuQyTNMAx4eL0u5FZOXqjwUIG5T5FEiQ9QxJBbUYby2T6HcbqsUa0MTTQJ05/28Oq1M
NIExn46UgxtcfVIl7kwNosq9VHwRUAvRUQ45cxMaa4piYbpg5emMtde0wI4JLWQR78sIZeb6NtBJ
UaGavorjlRvFCFQlqwD8MEshSs5DXAJgeRJ0TPeaPymKUWyiAFL1dt8Or7q/colmNFUZh+qCNDcH
h1KoLWHVxuizoHDD9t/PpOxMuCOGMowbc7T9bazyJ8RdNszKTjmtNdqFO4aQlsl0g0axz7kVMmJb
jljF2ttij3yNTl/QHnwFkHbekhyQI+kyTL5O6O9qY4mTYo0qUwDAvewdKzC8QyYYvW9/f0j3KwJi
/OVy05qiZGGesU/CWgMrqVqePm87oIVYanBRHKT9srUkWJXBn7nhMAMNZuEMQGhmuKk++l1S6u3E
tUnEkJoFWU1c+6qcpwaNALPUfDISJWIi0Dg5F2K5tLDpvQ6ClYL4HDhcKC3KoTyrsmslwnJzJR36
Vt9Nde1rRXp/Ue2cBpYPcKQw+DPaI0SE1ME4G6p7+/sArBupFuP/HVLIS6QjtzyIpWQT4acMPY5w
uTEM4detxfXCUvoS3XCQ5Ggs2w0oA/5oYIz95Oj4brSOuufWEei63U+NKkgtn/l11ZJE+C+jaQWR
qvwoexHGrCVIwJBrbW5JGglOszUTxcs2HNKoKmYy6FUuPZh5fAGrnktHkGPZ1sHd+H2MyYfwB+R1
5wunjJkSYez0wBPs8m+cr1rgZS+X69WNlRpjHJh9V87LXWe2AosQAhsWICLXnHpANvfN0IGV2/Eh
GP0VmPLUhCdqCHe7WiB025udPBtyXIgPoO8pF/1rwcUtnrU6XQdRdjm5LebFMZLoCftKanQV7SiR
r+DdE753WGCthMipNsHFPP1NYUwBHAs3MoTxzqMYnyizbdRmC9+ptSd5WzZ6uK1InOjbvW8RpcEX
yfsENd0Sagleh/xjWgAuQoJ9oERMIxPWEQ6lB74t6NuPT3VcYsaJfYZdOu6af2iNSsHxqV0N9ZUE
6bXLmQNNdGNK0v934AyktjJrtmHDlu2zgcDCyqLMiGQnJkpr/KDo0Zq5tl18SbfdIMOp755dptPe
yKF4gOOfdoDNy+lYJGm8JoPmVNx1ITYaeAKaq807yIfT4JYlJPhCupBkiVkcSxuW4/DdRw0X0x7x
EoG1YyzXbyR709pUITqRurkMce4VtpxYfiINwIs8TfeVlDR4ixmu+ubqXfnPJoRHuSBI9WFDqit/
HaYUeEa799Zdhmlde/j4b8nqCJhuDYjAL6EnHPUGiRp8ErApYGIchk6Bk/91CN7eOi0E0L3U60J0
YnXV6cLtolnbXTmSpW6s7ZL0U6e7gSIk8AxO2TVLBAbEiZFVXW7vnlzpUlGshjoe25g61rywUctD
qD5KAQTupWCT+MvigKWeLFO938+QlYS8skiByOSzZn33n4a+ycf1dQ+t3U8Fb5rVdT9fYUhZhtxG
c2eHzXJHh42t7pYRJrcYL9TW6u1XUzLFxwcGWc9G3kHpJAsxhj5vjJpLsf/XReh4Gi546bCGWyv4
MEMmo0R7VbnbOze/TmYhjN6mR8a8Ow6ce8G/uQ8fpTlX/Gcj9R2RbZJ1Nz5C39P9nUzf+aewnJg8
ZPNKYPQiDreuLQW5D+VFv2E4TAbq1nXBzGBcxf6rYnJQPOY9Yaw5X6tQfbOzn2rMbqdKDSrwTZ+K
epeTX5YFr9qiR0AUKzSHmvMCrELNs7M/XZXnLYa8moMV/onzNVZKL5LkjGCTTg2NZKyM2WmW76G8
P5NWnE2RGL8vSoYUCh+f7rikXBP/zODRqOoGQewX9fE4ycCVzzMYER4LDV+agL/4MeFceBXPlt/O
kRUi9Q7/uTAo33QM5lDBeZ5Tc7+bkOZXVJba5AIqenmiqAFf92hkXTqHiG5nJEeSF5iVYjY2rXRD
9/BbsEP6lhUf1baubn9FbhHqxnmDuZrQwiAmVPaLNh3SeUqU90g+RpD25/F5BLTZrL7uzlqt46CW
8CPOK2Wkxuj2cSkOrjet7SxOqxTpZQ/ejvqzDyOaiU2/QQqHl9BXgWEOFUMaV2yE39jfOYabpUjr
CkhbgbsGwXSn8JxUfY1QAcU3JIf2JGuEpRwV+Gnn4tICOjdrBSImoVZ5RBMaWEXAZ04sPByv7keW
z57qJpGEwACw03hASw9WTdn0ah3S8UrHV86eJyDMCs3D7AxVmmBzkiamHheoMRapn6uLSpVQr0TS
A6mw5jLm+brpVjbTtFUgpmoVwxuM7GgeWhAsUQOticVqbScPdVA/caJD+gdT+7gAsd3MDIYFZHY4
m7bqpdPdnMzx6TW92QFuPmL0k947669boCRI+tW/P07JX1H4kbFd+US0GY28r5pMdWsHJgubq63E
rIsT19o1nXU0q99id8DV1Dv5S44krgrK4gM//PBHdrh+0+Ds4tM/QQC0eETU8EYoFp8WJWVHt8oR
EpjPraFaWTpDMf1y7klllLnjX6ZQCB/HME+UmrGcs7l7Q5Ry5rdCzBJEhO6njtVQTuXZ+rzldZQs
jxU+gceMZFzMiBqFvZOQxs4ffQvaESTgtEhrvDE+7kz6yYuaTduhnDfxW3qjAFp3aN2qQWtiCQPH
sPWC6A1Ne/8PddDwbYw1Mh8Z3Bi/HCQkTS2zMyaYgQXYhX+qSOYqSxzAzDqfb5timlquHFcnPiyk
FgnDsqDgwWMtP7Yn8G4ASSSP2qtrUchgKB/uA20kMAzjsOI9/4r4DbaE8++gysLFn5o9LD0vC8Uc
FEqUmoi6mzN6kQ1rfQqhXdZjA5At7/+/Dwgz6o97W8rzNkz8gC5K+TrtGxkNmpAsAmM17me44iSr
tgprpnfJuJnfnhUioJrUHC01vW+PLvXkgqZizPRusVOllHoUqWFka8NzHStGMqhdRF3w+Rpm2WhZ
5hlcsfcBLuHq/13zlXC2L05ZVvlW8OdIpO6ROnUlw7GxI3isWNcX1Xr+8nMmbvZJ2zRL7qWZ/du1
rQKAV3EzGsTbOfW+fzt5rShc9frslE/Ic8/Rg+qsDXqLmhGG8Zq/PCBkdXhQ0XUWVSGHJLm+3qST
L1OtxMUiTXWnScIkbLaC/0B85TKWHcFPQ6Ic3WTblrBqmu7MY9k53cT3W4dbxPGig3Z6vxFMDLSu
WOdQo6S39RXIYnTpOsVj8MnB7S5bfvJV5ebyRJekuPqc5CahHU23yQ5SDmodI4mnV5wT5fHxWurL
8+z2BzQIQhFLZx3wS78shrbdk1uK5e3hBYjBO7S9LeXfZN7WErsJ1wn7EfHKnNXJjlOqUfATXMz8
3T9H1fjIGYM8nY7J4YVbw8DcLFAz5fv5n94dGqQ7hURUG9elSekmCY2nJI+tDYyBh0ftVUdqvKHy
1tf/r0RKEzjdjhF045xcbXaw7ZR/fYVqWQ7bpQau728QOXs3Usk85yQFBVzfbuzdpuMLmPLzm3PJ
yaB1cosEKZxGdwB6Ks00/Y2W6qxDiGnMTYl0cIvQ21M01NUeTCJSpAPFX4Qu7yD0Mvivw30B2ZYl
fMQbSlB83OpcoEMcmaFnYkoG8S2U3zIIYjmAPQKa+odHKgPYQglhQ+Bxj73KgKv1hI3fgXDDUrgN
n9Q9J+kStIIE6Lgy6WGc9KtYRAmnFoLAsm7jc+U5H5VsOHNG4P0c/Rr4+jewwv7CZ8VnXrYXN+BO
9vgLgLD+6U+Olcl/rovzzEEhRa+2UGElt5srfe1xQ+2x2X5HQgqgcO91r7z2FdvjRJ1fRDvWk21e
dJn96SIhMdqoTj46jHfX1igibMnk02l3G7JWC0f3Om1G7JCgKL+cnjIdFzoZ9CKaBDbPotRdqTSD
TN/4PkhIBBTYcDzgXr3hWBw4MZf6lG7t6ci9qizmFlvY3qTx7Qc2hbekxEMvJKPmI3oTsxue654e
wOvBxkUnJTE/hUB4qWQE7daVKP83Yad2TBlDaFgakHCv61bmCZj4yqSaUsaMZF/wv2gGCzzdamPE
WjG4pYIKheRzb2t/wJzPB3Ppd5c/Ou2CsruueWW2P0NNiU8TsDUjzJTk4Yxb8RKgRCvwdezaCeEP
+WDznannBtYcJlw3B/2tDM6EN9yAPvKfczz4Xcd3zuHYE0ML+94PZbTEFsX5cc4ULt0rPDJVtjhE
LChCJQ5HC/4X1x9CYGbQyQVNigYz7y86r+ChJMEpkE6dSE7E4PNJ7Mnfi/aDLK77kFKAnhctzU3X
9qU4ayl3FH8rjzWQu5xpO8TPOFNtzw05kX8SxyUaj955jOoo28FZhvhN5f5veOUU7aL2tGeaz+bh
JXjcXV5H2SKatYftiaivCnyJlnv0idDBSx5qZtQ0/BBwfPazAMtRB9U+PWhIIjjK2erLhGQojZMX
6DFULYv0WXUu9Ft1l+MggHZFpESio2OzHVODotCcdGeNBtkDcY0tW5eiMFAZ2pIdVvhLIF6/heae
1Ezj3RORzrVeaKh7HY3cy/sRuXpLAhbcLRAsBcrQmCTfJ9Sco8zsgcnvnIqvgtxMu4/2k0x+DZt7
KSuAyZXTBNU7GwHGBfeSyvOI+C6eZQ8ezssvnYr5XLlYkBeKrwXaQW6XHbXIJCzzsdZ67FU0mayM
+OstsIodqwSQact5Sr6ER0NAdxbGS4toEuvJ5i7kx5yY26/tjir7lXVwNAvtNc3AvfYmEfYEChFS
CDOXBzZ9kJgiG68qHIWlMrOOHvKBkmrqP9F/+47NQw/T06fEcR3ABtnWBU68Xs0qkRtVYzwMatKf
scafbMVdd2k/7o746kbnXtmoDGdESXzpzUHu1Y/dXKtnxZz1xR59vlA+UzUHilFr6/vw6FrgD18d
lPDRjIlnKHKiLfywXS4lD5PhApx/BDds2UaM3eQ36mPIjCMMh02Nxn2M3+mZyhQScCX6FN0dgx5W
NPg0rcJTtpFDO2N65YFXTq96BgMTcxmCxoHwWMFDqP4gfZzCluCt7b6MB833c+4T6+T40X/r1pNz
jGdjIrJYzsoqS4ML8NlCge6EWlplRrujrWh8wOCkwV0hNUOKP+9RqRmKahGq3tydfc8l9Iqc6sW3
hylnLi2q0gSSBHjz7iYWd4sLuNbqh0AFghAUthbJJ8Ii1RSDGn+eIULuJJx/RWvzb9vD2SmLiHj0
DBtQ/7McULA2bhlXWkqDMa9uW0ByE4Q2NwaajQp19yU70q+XvgsidOwNoUOp/9GoNApcN69T2Fwt
ljqquWkRilrIo5lxvWqnjfgUYUY4WWSCCCZLE8Sh3LZzgWWEM6Igw5aVVaBcmrrIEafin9VWp0er
hPoNLHT6nFgSo/AvuHXDFU6NN8xyntmTuX42nlDGUeWUbAjZ0ipR10EWZMFHH8/ycy+I4hhUsmA2
fP2evX0rdLYgbCtUYxinJmG87NtUNPNh89ktHirUEhbJ+X4IG0x/7v51/ubIm7XIUvUkWqomebUm
sd6KRuRAQi0j79u3JpHohK3NYvyLVRF0lPQg0HTqULZZEMroLlo9bzCqlCu9K2P33L1OgL0w7p+V
Hs6F1mGxVcgoVGf4Mea+cOjg5tHOpxcV4zsxg1M2w+xP5caSrI2/b4U0Unh2TVPaHWMsXrkWNBgT
dxeE7oLkhpl4X/0LQ6O0pd4V1QjmgBBDfgCRw3+oWDOMOb/iV2HcWfzilRqFicWyowSPOd6gp33+
qMB4n66SeqILffIsEwYQg2V6V5DJrmMk5pJB/B5UmXVIOkCph2+5+1wLXw45NJN244VEdypC4Ow1
AmGO/ylFedaqPuFTpLkbwlzlc7CkPHvmvKDoMpB0hPUqWS1/AHlpgWKw1/WT0aWKzfOazyBF4t+Y
K7ATXhnitzAYdoB5QJzfIOumXGnazXew76DzgEQYybcIPhv4RGeqZkOb/cWN+NT+Q3h8VaH1rZ42
qf5TfLBP/u0Y0GAopasOg7QskGQGb2Hre86KpSTPnyfzkxMQuMkWWNibcbd8+Md5M3WWXc9WClq8
n5rS0BAmUFXrp37OsIuDh2hi6mdYuJOcFcbaDnwz5YV7wSYO7h39R+TZIKUdaOZOqUa9x94+KQiN
JISDFTeAggETIvgcpGltenAY8pIoJICXp5iEmw4Wspc6Zv52a2GSGbk5P16eN3PekePHdyF7dIMn
4ipwg9KxKTmqXHRQHcnPdwN0ofCUsSnuKYqgBGfdtAOxGBBRAaQZ2HFJmsya3ii57rjw1kn/xGAq
DemObZumvuzUYnHrGMPbNidS+IKs1Y04Km7Rr+hpnah3qMobhozNr891PouY2yA4VW+B54/4jDA9
81h8NzIDRlz3YrBdvpRQfpHYbQPZMnDONLWpEWOpi+hvaDH3xj590v6lGy5UT9Wt5rJPLE/rn5a1
6KrNzw6d0nERz67nuEbYztUJ5p4kInNcytWe1ksHohyCWDlttyWJwH/mf0VBIPiIDgG+NVA9U99r
4J6cDg3ZaW+M4SfTXiPhknLrSI4oKudecT06BKfVehg9T2efPKOEvDsIrCMEtHdmGwH7ap2lMLXG
/V896uGnwSJpvCYWhlZEb8MUtEPuzIAdhUFlaFiKw7whx1jG1MAbPWUvgHmEoLf2huRM8zeBGA+T
IPjNSWWS3PBlzFwidnBVxm5+YN9d9a7lAh7OzeMmJPYtdgGmGdT+HvX8XIB4avVw2WfmHM7qTT00
Fh0XT48z85/GLFhsrM0sbaFl17X12KR/NDrJz4kDmBlx6ZtHwd0+gma15OUJZooFJBkAToyehIIH
fVTv/DbGP/pZMvVIUl2CKVS6y8DVts0VyjDyl34TBGHmgp8M2+vg72xW4nSqKt5hkdMk2jdD/EJy
jv65QrQCzvvConcrF4lvjar8UHn5WJVW5SmxJmnHxbH7I5M3WAda8gh4OYlDRqumLbhZFqupTCT7
NRUUCvLTdmqlcFjatuj2pueBZMrHcuWa05mWVoUKgdPb7HnL8ZyQsma8qUmshBlt+w2SbLEPAAJi
Z8tU+8daRYMEbKF2vyU0iIr5f/5LK2qIcVPXGZd5dnJCH+whbe5rWi0ZX4wSZXvSDk6HAqRg3ksi
9MqofjXBRb7VJhTYc7lJu+jfHxxnqrRnr7VUrs2rwF0C7nbcKvBRM0RLTKNOxD444oa/p2H4FMcX
nvUT2H6Yfhugf2zEhlMJoAxJM+Z37QmA+Sua1JpKsSQSR4xtDp/Fe9YimwZwmqtZZVImX2XlsXzw
jTVux5DOgvfLnK1r7bqsJ7zirrdWzhLG7h1acMZ+J4KLy25t0snB7wMH3kVZE5uAbi5ogCKjtsa9
RY4uI5WU6TnyuwI3vCAbizYEc19lfdtPWlz4TCFS/KNjpTR77ha8EWUhiQlfj+lPTr1VCNy8J2WL
XUeodmp9OyJo71y/k9PsjbMXBgIK+akSIyhsVahQgchi8mfoxH73p3qYIbOxe9Pz8m7zTLpe98Dw
SflxavpNINDfoPRRJouuNQU2F2XnZk5RNiCRd/1SAZjsA/jeFKgyU+wSG0ra6ZpFVW89sH+rr82e
rOKFc2duiu53tSSdVIQCHdwlrAd7tGvPfMKujIR5kHbhIisMs7ApA5yQqSdeafJL25qOf6oxAr0Y
dcJ5BOVQfXNwsU+NiOP+QQ05KEkVLgRhgxgeEbQ98KGHy1mGLU8C3rWL3lIJRbUK7caI8k3rqq0T
9fH6iP+VTiwTlA2WySFrPElYsh57tUAa0tVhKDIHZDxVnSMLPFKxpe4RMq+Hgx0RY7k1ZMvYmm6r
7ktyGs2UVPejpTZ0zUILnxExX2ZLV2XCRlWj6K45uzf11SzhbbUl2z4cd5jQTbisaxrnyHtO3PFm
1K4jVER27KKhDZO4FoVzqza4ZSlXizlyDaHfsYVVJ8vARdA0qzck8MhOP8Y8kmJoRcdg+nwVFNt1
yh5LkMvmiXZbC5JXZE4JTJwJmI1Wd0Z91ydmU6tEwio0dXwx2pLt0JPqDSNNNQWAB4pMfIWYornZ
YvoUZTx+uRDY3ZCt7qSIQmSQmeTqCATfFjthLldbJsgkI4gY+QNYcOwWhTUP69kkVk3dzTJQ4zbL
w2EzjXtoAklNAmqnS/fX0fnbYRKvZpG2R71GSkL6/9x9EXPnGS3nlElz+C0+RVi+FDeEYZjwuKO8
fgNQ4wRxP3zL3zL2ql7mqbE+LfcR3dctHgxFQifhNlb0AFqcl+ujImSsI0EyZGfFe84ZATep2uUZ
f24+euD4bf7y/8cq7wxZunC50Lf/KXMtnVVpSUhIrXG7kIB1MKjNToQ4bX1atW0m0jCg18YVFlXT
4jfc4IHcKpriwhdfxb2pI45B2EIbmQeOL2XcqlaR2tZxh9wxLuhXnzcExFjl3LeSgKYf5KxnY0UZ
xsbQrKVHSb+QPqD7XoconXHOX8aevdiMFMDFw9OCh/S8vrIMyVsWnw+qhvBrkVTag93hLKZlSyo2
5g71FqFtbuEG4KPhAVKmRI/h9Qiw0AhUidlExNzeGYYcQ1geMCniktVU/hgJ4rrHijZr3a6xP/d6
n5vfy/sp7I67wGCwZwWrgBulITY7ywKavI18L8mWx6uumHcUODv+HJ9ArthWh8IQq1e6E7ftWX93
2Cas5/8fbvd9vF8vlI/2SC1uX5tkNuRccZao1ki21QwQRHDrjByQeavAgmOuCB7jygnT12+WCj3S
jC8utOzeMSGisMdnJAsTUsoK2RzvCpg7h1FYD545wt+4ReueNCBADPIksJCSMMoUxvkJE6bhVm0n
eRQVt6EgFJSy3gQjTz+xPq7gAbRKMxtGoEwuU2ABM4U12NDLk15AYJEv50jJ7Ct81pMgdrbLkj6P
YnOOfVxIrJ01EXFcBGeQDCFskL8VXsxgGxA8TfvD3YXqmwJbab1Ts3m76Npy28yREyaQY/BLLGjA
7BvNfJGDpk3vQhcgydTDO6vvRf6w4MNRzWHgdwYunJv7OIi9SH1HtiqmaIEH9kZnAJ3jQH1JlvHo
4pLxjYbaRcd33OAltoJvtsEZBzxcY0K165hIGxnVklQAmcjFssQAPzLxrK49WtrijX5JWTJa7nRz
urgVWkcSGeIMmI4yaubaBrqbCCgDB6aLkJoFZ2IEUDbshZglBSSjqCRxTtyS8SrIlUH7Mr/QGzJi
6fZzuFkVWimsLdfNRNQ50PLImwF6PTAFFvMZDqzTiQmMwEQFlxlHXxBGtYfz9Bv9ub9oCBPxONKs
dY5NDG0dmzh4wNPccTXQyePBGkBnjEwP6ytFqYHOOD/WfXGCMPVlelm9WGty7lgQgQVjBkMpuGXz
V3zx0tYyJhgz3wlHrrpjWSfv5Whf4VqblV4Gh15CK06zbPCR8jNVAvVTxeFukQSgcNPV4R+a5JIz
iXfCg3Nd+kXvIU3q3B05Z2ZeWR5kL8L9EUcDBiEC2HV1lEhV+RDB4ojk2rD7/f6zBTM6BWk8AJSC
JfLhAzFQ+3Gp8109sfxpQXmDf4b+PyVPi23WNo9LO7LAgYCvha2s5e5giQbPeDEI54v06ci3lhxf
/OlcPHOHhPF2EKEEFdcVobUzCID/1F2MBEa9k8iMlgIOhyRkNSq8VbNnSlc+4K7Qtw2sXlL200MW
J8rV5KbIlmFTkv0cgv/g6rzff32nIW655HFySnowDTD9t8QnOMe3+O7/1XgNYlcEH7IGoXhZCns6
Pb/bmpR3Mau2FWBuIn5W1y+UBG8f5EiS7e7w8bV3OfNS/d6vIpc1XLGTiij0T3t6E9/8QzKgM2cm
wWfeUOC7OhrAOJgHknRCaAUlk+O6ZdCD6FBhfof6qOLF424fFAVVAH2JLeRgQc9kmMwqVw+TwtMX
oy0dl6hUpr++qBe72ocMvqg3cyT1QHr25ZRemaQP6LrZtL3bXR7oMI6RxBnpkDU7j8xhiSiV79Dy
YPW8zhGRvzlXoAj/bZtyyV+Zn5N9U6pA3NcurbOZvBCI+NM3y4U63lS8jOXuPQ1OK+8kn0NbYQWS
mDaW2i/zLbUcUH8nzoxzOk7Mu/nwrO13eTKgx4oxAhx32bKfZBOcGi7UwoRQRP+/TBTJeAAimL0c
LLvtBi3JThhSD/bcXvWI2hSP0RQ58oBix3UxARtfMruqINjU+Nl9aZCswar+A+cMPDfLX+oYowx8
WcQ6Ee96NSkpixsaVtQSmw+Jh5c+2yo/c8nwiO3xsmInQ8dIs0n0a91eIGAvLmvkmaJSmSN227Rf
fpDiSNdY2ZnSCUgoBDmDmzlwLNaaWepntbBeQykrO9KCg7rP92x3eAVwnfvx7mS+UpBE+vGmmgZY
CQNKEEeqL240g5VkNfqhWWKEoKwENqnVWStJnMV+QNSRBhjTRwgAB+DXJqKLIBlFSBCFAsOL4BVn
/YtSFudevwXp5KRWLEmyIwRuShRwea5lfP/cOv49nfcYWq/ix0qBH5coxMJzGRmd4YYGY5yD+GVH
TzJam+/S//6BLUovOvrWTopqsWYu1fGSFA4GYYh1sSaaQLp9aQXVweIKL1/XKkPAFT+hSLRkc4CI
a7BNJb8B5U+wZel50GBSyDgE3wVW6XPTF2hq6wVgXIKL9iB0brixp0IvXZt6ITg2BS1TM2bEkfbC
Qt0ClD4hNYRa3/41pBD2xmIM2UTRLvvlXwFam1FM81E/+hw4mYMkAQr4i3ch1wSLGWTO47FA4NoJ
8idCoH06bSD9ZTIhZtuhykgKLoICn9ADw5etjPFCAsiD0o8ZgY99ARlDDhmkbL6oSq4Sw3YwHAiZ
AK1fPSpTanXFfY21Pz8ejIp01MrzJHIgcaJwisfis/HF3ucYdFPopHp45c/1FxZlYNqc+zpD+PT7
k/9vrFQsua8PJ8faqJwcZoEBHhv4bUoSTJSfy/diekgqw0SCfAnPTSKBZzhIlgh9PiX315AaJG4s
lTHOrWbLYuAvuCNcgZBgKAHBUlrnzZ2UniuBZe+6LJRK4tO/3GScF+Vv4kmdzO0Ulf6CaW4GRbg6
tn3M6KqJIvfx+a68Npjkp33pshSU2v+W1AKiGqtdMNOhP8CC+r9fNTjkLRU811gp27vKRckreS8V
3dq/gAuqHpsUcrdpIwvK7hfsjxs10SZI9C7C7dMO3+onE2LAEyk365Eu6fOshzjwwY2b6pw9tIJE
Bh3Y68swZ61FlnVJ8ejXsnroiqH6CFYPxVxUhweiQUt418cuLkvsaot4Lv+n2QM/Vk8eow+Zkpad
ubAhY0Nm2eEKwf9nm+Xu6FOhbieqjG21mGvYL5nTptQMoFvAoj1SnJGzOU0YZY9tSlh4wQzOckXh
cm+xWLRFZoH3ssVTDKojsU6ydo+uXLp5WpUzHMmvank5SDpQa0SaZzww7WFfRwcnAq406MmDMsFz
arWgraplWXd0r7an5TLwoX8B+vdG5J/XQuXsdZg44RuSx9r4boMfYuItpnk7WbHy/SUnhgyYswoL
G7yNODWhf961YC+NJufsZT5Kn3IstZ/c9sQSJgiKG8Y6VQ47BgI2duSilpHsoSz+apxGdA4vPFeq
Ko4F30VGiaP06TUS0BgRbx2rsc6OYhQksBH/hNC9T3lOvN+NoCJb3TH4+vK+YWotuuQnrPGMWQ2x
FD159pcbaL26ooxG+VgwbTYdc6UaoYvtpgWnW1WHWT8D/S9gLhrZLlfOLvvkUyDglKT8ak52IwxZ
NVD5VME2lROCU434NZUUX7hJhb60cPpkGRHe3EDRD58E+fNlPRD26D6QBsutLz9pxjZe5SOGiQJv
ewsuhbiGZR8jmV78xkGqP8y1YhBHXrzW3ADRS/ORZmDIBQi+EuVAQPso9V7ZZrppCiHU4dkpOE4P
KIyzLW2mBZVCTLnl7cAMCW+M3jUPB/CEUBNnUTq/1asV1O4EHd9Pbo9wHzmZupntqYj/A9AlhN3K
wiqG0nXqoErWDWgwWxDVA4BDRYThuzXdOvKcmh0ORFLmBMcrpRrX2dkUV/bc1/DFo/HGiIJAJ7lc
rgVmdMWp3NnLQR6nwY0nCMMDuciPid/h9s7ZFu6NXjWmB1Xi9KNJlnd1bKSOxyaXhNB3pwzFxDZL
Pg/IIp82cyeW2HiIu8IkPHST4fBG67tUIY+yL+J1unnk8we/U2mBWCJP+fZrMQLUtKtT5obO6Evf
GgphEA89kQSJCFX56f7s85KbXQ3cPhMM4NgcaeC9IksBbKX/E8VQxQOkVYrbenSiwGvZttTUBbnS
p/d/u2Nz+YNxIU+w80No3ike870K3dAQdlZaDD7AKSM8S6vAaz5yCxNXhbOIwQV238mU8TDTzVKd
VnZBBxuvLuR5dpPeMsN34owQ2+9G/jPElp7CQ2pf4kTpWjQpBFMQehE5UCYAvq59PjvONRuJQnBX
4GY0y0Qmkjcyv+t47GyRSSmpTclrXpely1vIcImETgwzt7yA6h23GCy+hDp0hWNrp40GstjOH7HS
wx0Fu4htOPBM8Eq0BQ8YVHSTz0aV2AC1JKRklZiRK3USUE6oyI1t0hHw6u46Buuj3aFhamPgbbUP
TmvL2TcjN4sB1ngP8fZgfwvPzSBg7937DzsEAHQTpyOUwciu/ipnpWhId+V2XZtRhELzimUOQrxe
uHZeldyY7OsrPuRI4q3eqZhR2SaZ/8ralwJ+/1MIRCkDldxzptGGFjTyKk3T3yZ2ZZtLy1EVGyOc
DgqM57JI7m4ZZuOTlATMctQ0xz77yq65VMOrSkolThSrDY6ajSVPvrNGSGk0hNPh0pBwqh2/KPtr
T/wKEELSO192bCydjZ8W6D3PgiglaIhHTLvHI7Neda12Gkw3XuwD611q6ALGw8WAOe1sO5Weux8X
pK+f0OP6RyCWlOTtdI0ybyMPABRuTM0bYpxL5D/SC1d6Dkx1/ENDsM7m4Ncy05rU2pfuMjq7tREA
Io8UvABx3GtZF4S5Wp6SRyTYFfC3NYRGEBjkJ6mGcfs5t/ymJRw4ILjScRJpYlgRbQ4kYNWF6C1j
2pOqnym1Vz2B3PhhR70EyvEU68Q0SDuTyjlRWzktBEwDv2ogK5RZnDd9IQl7S1nco73MLliKOraU
okiN+2bmfaFVdMi7UExU3GrZ+CFx9jf4PPZZyqKI7IQQjyqVuT5k0+H3yZ/E1ZiSsvqtBI8btvkC
IeR+URnGSPSKRMecNigNxIPIOrvXiNMIi7PUkaGBgitdjFG8jMFibU7hXRwObh1D3te47CPjIKbn
EgG1tyzkePiWrgqXF5Fa2qMiX3Q5UciE7scS0C7f7bsF2IJXlNt+UTCN4OqXqSpx1sdQ39H0qiye
8CqXlTLqeSq7GSOr+yOK998V7IlSdHKsVt6moALgbycEqRJEN0xmhxbp+QkjCfJfxcuMfTrWF2PA
vVEW22qLWZ4+8Qa9FjqJWWg8l74Unk5bVseho/ip2n5gGcBGjlSDCadHk0JY3OhkLd69v6+pjKzh
S0PysIMLzEv4ayGtDSKma1AOZNGlOXetsVAsraWj1QOBpgVHzlzSepwxNo56zRvl+jkv34tBWjlg
1or+xcTNBREXFsMGBBVIlvOPlbvBejqJDY7AJy/19z3m47l0wCmHfAOrKktU7wR1zDi/iUbq5ElH
ST3LlFkaIqSptLVDea9cPhU5m8+HJLLwYf09ZpTKZpt4AmJuSZqeqhTLJzV4iE1bIVufcmmiJOuL
JF06xAgQYZEGAvue/sQEgNQglOYjvMgs7YZdh+36KOVpMe+sy97xqU42mA/P6+m/xAVqy7fNSXM4
EAcoHF7zWJDtq/N+Rqm3WwvexIK8YH+0lJuQqL7uObJGZMqv0C3aDXBoO5OVmZQ5S0HwowTS5fgp
vU3ZZ51CwflqQt22fDoP6W3svGRrprHfdPLF+Mnd66J56CR3Bd2Gg0L9k+h3oMyw9y9TxZMcKNEw
LPuknCLC8Ou8YIY+wS9fHi/avG9Ls9U2s0fhCrxjq9EGFQkKK8WCbneLaLVaKuQbodpWO9qN+15Y
HI4TpJC+qU7xZlZ9Fl8FmnMMfjlEdWJIKErqgdxk9DX9VgHEN0g5oYOCunz4WhUb3hGT5V7S9UeA
drzqTiqmiwiaeZPX7R05GOL6BRKRkfTRumCF2VKbGikY7FZclM/hi8fp8g40BE1q4L60ER+8Y2Cd
fblviENxhauCccypA2tycxE3dVPZfOLuVQreAeCWHOsgjwxxrJFXHOu13GXlVl2AdiZwaHvW4p5B
hbjDhcDQPBR4I0JrxpIXuCOVGdV6Z5wMuGrAMi8r5CWF2kc0nbDL5lAhvhD3fp/DldWkBqai1cRx
x37BypjacIA/pwsHWpE5Tiyzjfrajakcq1xDIPVseRP/tApHrtkXl/vpO2bGFPqQ+YpvRUWm6XSl
ptaCgT5z/2mpkVQ9drdrem7buT6N/uyXAzlRhLQUfMdjH679XJzG6gT6ZG0zOoI5YAHpLBx6XwZx
Vr+edzQ+LYWS0OZ4VKVQDFPMeC6+45dYLoa4gzLtfI3NWNEudTeR3hUa6g3TO8tAfAMM84kBN40z
J6i5ZNhTUj/DJ2hW22TuwEsyBaI2qVoLGt0MwgfWZc27JKePdeWPW8Ruz306z0aeNZ6qZ14oD1Ht
VztCmNE2BLjLMCs0cnJSTXPv8gbd8RPaZrmyBui2siUG5Ud3O5TZuXuOQ39u8HHBnVDf8SOmxG8t
oAmwBc9FBL8itJFP6UQ1pNuHkQR0Pqa/48W5ejrU53oSkpKWIxMYdBe3kMyE/C4WPdmXhiX77CoA
+MrAv01sRvoh8hcnUO4uZ1gM5mMndrOuYJ19EXbHGrJUjj8EXOjQUc2enXMw9CpqHR3U1kTHpmib
LdvjJ2rxSpcPj2m7jAM0J/gxXLz5FRUqP6+2aOLb1u00kh/dWCoJoNX9FsM7L/R19zQYpx2lVCiR
sBKN+vM/KSQatUpzqElgzfiBvsaf98RzczEh9kXhzSBV9AHWdxgb0d0BJnZ3EnWB416FxteVSjE+
J3Vvi8Ux4IIPhwJwbUrXXZvYV8sIVq5nAlG6WDRDwBarFVCbg7UKv8IAr21HViOiJJfmXWzz4RU0
uRSO1rO+hmuBL2HSia9gczYF8Ya1jiXX8VeIN/K/AqttIaXA/tIxCN6WOBrc+cO+wOymm1xfHB4W
N2z1QcuQUNAJgLWwHeKM5tNXAfeK5fnnhijV0briISi9A0NTyvNnhvrSnsX7UmLxeGJFcFDH6R9c
mNBvk9rA7/dB9DCmCdqut545r7bHaP1FQPY5HOYJK1pljUQ4z9GxoET59c75ksij1HqEDjyHp1ad
Nj1QWBzW6zL/16UoyxvQOZ+RABGV+5o8ZPCauUbH/Fz8CUjMsV4NDzfdVo+7H3X5cdVCTHFfqDkQ
cK21zilSFrHvVselRfPdSbSZ8J1RTJAlNQlMaf3a4Z0G9HAoq87+ZZN3G2HmwJCRDp6EC6w/VdnC
bF2axR1gDwTqpvnp8xRB30LxnvXIQN2cQuzmSv/mEGeb6S6RihSeWQSnChl9u4wrcHRvXwWm1EgO
FaWDsLS6eY7BPqOeI/DTZsmWLxiD/bSv7eXijrlarEUu/lgPPV2wjpmx2f3cKOPAgEid7tuV23y0
u8B9axsOX6JbBS1VeLLidIl5xo0E6xbUDbNLDxVQzFW1Y5HrggUYUovH6a0uxIfidtOJ5X6tuqsc
PzYo4VTO8IM/rNvM52boo9L5zZc3klyJ8+aNT8lP24OJEWEBpiJwF8bsEryHUVhEnVhxeNOlRRlr
7A6jzB/yUpjEW/M/5heGhsZ1ZMo9f5lwNyoIFJj7eWRFtsuJFf/lvu+Xw7w9T25a9WFWpmI9PZwV
rQU4Bytgzxbgr+tsD5EvWkdK8+TJDyQjKCHrvG5Wud0+yzsd/MfdqCoFx9XYcSzrS3f5KJr7tY9e
L4RnIF/fl9r0ZhlIPzTv+T6TXPO3X2b1YakKCNLP2xGX31TPISsSpqE2T3s8o+ti4aJ+x32/C+XN
pt9c98s7IE+JVXweoFpnstQedzlTZucCRuiHfkHc/uk=

`pragma protect end_protected

