��/  ��Q(���]G%�B�C��G�1�*�$�^�Z��%�������[�Wq�~`�	v�.@s�Yꥱ��+[q�~�����h\x�W�f��O�盁G{b�]���i {����~.q}<�	���`�� �)���(�c�,��e�ط�>�KE��u�ɕR\Q�YL���PB����m�8� ��_�LJ���6R�vݼ�����b<�"�i��7k��n�.[����i�P.Ǚ������-:O?}��԰}DHK8�19v\P�X���xy�g�g
��s��5\Pa3Q��D��ʽ���+l�BJ�u�Ƹ�2~J��YJi�Pي��]�8U�~��6+Vo[L����P͸�F�2Mvș� �pX��"�����]u$���iJ�Z�oֵL,4S,�����] iR�����GJ���5�1>9
!\.��pU:#q�&���n|d� pnW6{Z��U�3u�}���eR=u�f��ǹ���P�>@g����#fm�k&����Q�xI`+��8���j�Q��e	B��y�!)e]K0*�s���c���u���d���f�ꦾ/��iݍSg)-��DM���Tt�Đ�JO��K�ؗ� Vq�F�@�:�n���A��H�A�ܜ�G\�}�����S���R�%+�4��p;��+S/S3�GA������2
f�ܵqf%� =h�s���,\a���R�������`�s)˺��j����˅���o�?���1�{�Av��vTZ�O�����������s�ȾF����tڗ�Jꮣ{����cu]G��F�x��,�$�D��*��x�4�m��V�W{��vB�a(��<�nw{�������k�Z����R��������ʛ��Dv�x)�vIM���,V�=�_��+�ߨ�}.w��ʶ3'��pe��5�e�k��$�5!��X��eK |v�l�c���4�g�L��X�Xm	�_ #,�$��v���A�g������+���FfvP5���!��Z<�� �g����~�J�;w0R�) ^� o_@���b��W{����\��)~��?Q��N���iɬ���e�|-�!���gG]��.#~�I��
z-;bs秧@�C�h�.�n�_�]���v�qGC������'�\�X�޶1�<�U�m��6>�|�՛Bwa{�wK����Or��^�Lȭ�,����T�Os�c0�[���x���lĚ*�E����)��W�a�t�M�����輥�O��n���m�К���Y,_P�횲����s����jYz�>�y�s�XD��?����>�asdAh�ߩ��S��M�G����t�����F�(tbz��@1����V\m�2Bm5��6�#nq��}5�Աv�Tp��Jƀ���"-����_�˴�#щU�����69}ُ|�	h��tE�Pf���2s塿�����k-|��q}Ӆ,Xgö�p��3��<Ǔ��ݹ��A�[d�,f�-f�yJ�у.�.�I_���5�n��*�>��uN&����%��c�M�h����R�Btcj� ��Ś���쩐�m��hH���Z�����J,*��Y�;�ωx!xC� ݒ8p��̯�Q�� /�N��t�8-`��*~;�\K���Lf����v��b��������xՔ��1)����E[=�]6LKN�O��!r8;y�K���o:��'�:���W�44�Ҽ���Ɛo�"�)��{��E%��j�E~b?���:(�iQ%z8]��kl��>a�W$j��Q� '��g�w�NB�K`Lv�}3ݑ�i=�&�"ȇcP��uG�&�T2"�����NNr͚��ˀ���mU$�
�����mԫ5 ~ф����u���&خ�
�X�/�����
fyQ����M0���Jr�+��<���|Lw��*���f*$��4�a�[�!���/��|��2��I�sɏU��P�Sک��-gB4~e
#-�s������j/�d�"Q:<��:�xR���P_|8�����ކS|�p���@������<�v4;�}�� ��Q4B'�/r�p�7�8O��|�Lm�'�J��>icN>��y�ͭ�A���Ĥ��B`��
�¾ќ��W����pV%�!M9�J�3ݹ����*�wY�"�g�PR�X��25��ݞC졀���9�BuI��}j�2��]�߻������u-q��ڟ�$����gZ����`g�t"�Ju	X������7��}Vx�����z�����,s��x���'�m��-;�O���eH�aP�6�1&�Z�;;�º�;��W�B2��9��~E���K�x���@jڜ�=��5��[Ŭ��5�X~��)�-����E�I)�Y��='8�->�q賺,~k"�����0���, ul���*t-eUa�O$R�bm��?�°3X�S���|�<p>wQ~�i�>~o�����5���.t��	U�������}��Q�K���c�v�٦����|��yb϶Ӓ��x��L#��/^P���8�]���FF?��go� >�Kk�`�e�'Ȳ(��*a���˿�lE�~o�.t|���+��{���z� bh���}�P���H�*CtlU������ 깍Sv�3=��ė�v���M؟��|<��p`q��0	u6CU�2��Dz �&Z��ZF曅)(����A	w����\���#z�V�&J*����A,�I(?e<�+_�_�!N���Ea 6@��mz	�╺�G�WŠEzt������)X������ގ�4�'�$��WCk���I�΋e� ��/�2��`��o)Ω�s���wB�֊-��I�3HE�Js���D�*�(璅�J��U+�z�Am6|�"YȺ��C��/rz�cO�:��f*� ��֣�=��� cS��&��d�m=��w��>"o����ڢ]���6� nV�2Yw؊��;�F�f��`�'�A-
0��-x�IYp;���M�zai�S+�t�L��nA��x0�T�;&�Hͼ1�33.�9���Қ�������و�����O�O`���B�L���4'�t��{� O����Uؔ;�:�� 4"��z�y�U�>�|�z�Ԓ�*�;�.ݨ�i��g�����f��y|��z�Z?Y���2#���ƹ��&��_e+�H���Y9nY��{��
�:Z�4l�̓{�|��@�F
��-�X/�����j)��� �j��B%��C@JoUWkּT�^j؛(Q�膩%N��^E�e�'E�v��@%T�`a��������qM
玵����DPZ��2D������+�b#�G���! �O(��&1�D*������{5Y�6{g��ߧ{��Q�bT5�-T�ѕǜ��t��0N�8�u5��]���)j�����:�Bv��]�؄ڢh���τ���[���eq�(��AJ�s�^c�\�Ծܟ��(&�F� <s�'�ɺtn�
�i%ż�f|(|Y�*Z�h��|���1�mv�}=wQ�g��z��>�ˁ�r=��ҿ��7Ҝ�����:'4��_����a��up��k��4qW�!�Ӛ0|f*J�����ySrc�c'��C{'e��aF��n�=����pv��E��r4�V�෾ٛ���Fݡ�Mz)3�����Y @ ,{��������L`<�b��z�}�b]@ExF�tm�B�W ���gGϘqv������i�2�"gv�UĄ�{��>�8�TM샳�e�k0�c3�Iv��S(�|���R6�P9c�a�����`�;��e�=fv�˂�����8��i��밈����@q;��/l6/{(���V�"��|1��t�Q�{���&!-��YU�����po��X�#f����l����z�ȁ?2f�ۚ��~dXf�����g��_g+��HZ0��쇣�#.=E�"�t���!�_߬^־�����u�3�G`w%_@V@���^86ap�ei���6 @�n��� d'�Ա%�ѮqM��*a��r�Fx>�^[�?fɕ�@u�����A�z�?$��'���%0+�J
�l�������1�Uw�y�@I�6����*�������4�	q�oWn����T���^�%���%�/E�Jbh�e�n��<�/S#�V����~[�]BX����yD�%K
�GXq��-KU��Z^n������GV�2��o���@�N�qs:��1��eܢ�||�NG���	�ن"W�\��X�ɯ��[Q.������Ah�K�����U ��Cg,.�L�0�� �F���-M�� Id-���e�`��$b@ZǵvZ�2��JJ&�{ EH�,�8��h" mS�83�"n%U�s�&���iT]g�nO�`��/A�=ʉ����1�4-I�U L�N�!XS��c��������ܯQ1$&x��9��>��Ԁx�6�-�$z7�
�gsa��6]�mR��̽ʍ��z/�C(�,�Bn�$u�Ϭ�~~���(e�f���B~>�`M��wq�`G���ϖ��JT��Rqb!c.��� �e��N���۝!���H�Mf6��VS����yڱ|�x�H ؓ�����+#���9<|v�1�`b�>�DQ�"Rh��y�A���Ͱ�ů�um�5h�]|�9z��B�`_G�n����%����e�'�Q�$7�m���$��Qna)~.����0���PT/�$R���8*w+]c)|�u.ύ�Z%�v�5�g�	<���j��.�>�b97$K%�*�W�a���'�3i�W��g���>�i��N�ܔN`f�3A��2�����6���P�miM(J]׆͓�n!��u��.��^t*��?��uq��.
2��wJ<ɪ2��0K�j�Ǩ�Hm�b7?�/�B�0�1�L�������V5�'n~]@���g���!�|�����L !(�S��Ω��aX�@����LJ����!}gt�ӛ��f�Z�jD�(a����4��J;�MI"�cO0�Q�e��"�/����Y4>������#���n������AF���h��Ҕ�ͼ�:��.��[�-
�s����~������[YT��kW}l�!+��.��Elya>�S�^�Ny������w3w��:�}d�~���0J��LF/�v�$�ϓ���S�}�e���hM��Ԅ�w:�5	5=l�������������k*&("�HÜ�>�Y!_w�M��gh���S{�.e��=/u&/�pce��r��CiϏ��5з_�&������+��̼�%���� r�C %�O[��3bY�*�%a�6y�������&x^�R��2I�:��=��TD�3A��]*pCR�]#z��O�ݭ��k|D_0��@_Eɻo�jm��M�o��M	c:���w��" g����F,!2.����~�hLU>�}��<�l���΄;�ޙ�%�����5��UfN����%Mi�����ټ`TUe�v�4���D�u�I�7���IQH���cp*��j���dBԅjH�(	��u�*�KO*Sa�p�n
�/�`�/h�/���;�T@МA��gm�{4��/�HR.%�c-�?�b}Rё�1e*����8��قt�"���Z� v���� �Cm�_���[;�&�,�#4��G�����^���V&��ߖ�@��*��n��~�8X�,
��$��u/<7%W��R����}Ȍ��F�:g������!2֌0'�&Qh���T'[�#~a�vٴf�~�Pt����z]uo��N_�smV߬��&v0�qv���d�by�ei7�٢7�풄=}z֡���*�B�Ma=�h)��{ a���-���b<���/q��ft�1L�S�0�2E��엧�\�%��¦���Y�&we�y���D�ٻ�hLo<$�Kʘ�'�Ǟ��#�"p��ay�$͒���ȭ��0����!�9�e�L�'��r�w/%�O	CFQ��/ɩ$I!�Yk��%R}y�c�RIL*�Tɴz	�MB��q4����Iy(�7=��j0�/��O#���f!�)/t�8N�B��A�-zc��-p
��g3�7IZ��RB��	f�+�xo��
�OI���t�����C�D�Սwj�NUtӏй/P�q4��γ����D�7y|� ]�����q�O=P���1��i��
�Xm=��34��u��$)r�S!�UY�K�&@�m�*n��U���������$/eL��{���C!��Bb9m��Oi+��[��-��v���m��U<3������_��Kĩ��4��a$��'�j��"�ଯ2�XX/�)��`��D�$������t,�8�Yȸi�Vș�!v(������t"&L�O@����M*��-�k��ʔ���E�i) (��%�v���78v�欬��pЃ�s��cƣ�q: ��þ�-��[F���tP��᧻Q��@>���Q)Z�E��Nw�K�6�n��*���VJ��ۊ�Y���kx����}z��O����`�֞(�D�:��f��J\��N��u�a��ؚZ��N-�1���^I:���&��'��C<�M�E�7=��/� �
Ø%Oe�`�������ǈ��p,�)�����`��u�G;�$���e���̿������n)��G{Q���$�K���ϔ���B����$���/���#Y<�25�����ˣf%s�(�S�[�<�[�P	�³B�j���9�Ց=vm���c�n�A
��3$"�V�K��&�Pש�*\{�z!��K�!KI���E4ƾ��јq{~Ü���&�F�"B��-���BOeA��+��Ȫ����&�d�`JF�s.���")"���`��_�lM8Zy���3�
8w��*u��ol	V@�J^:Ɛ2:	1
1�EPg�>-��#r����%�<V2�C$�E�%�cInj�ߘ�����a��229W�!�{��a��y����|]�;Q�ØI*Sj�r��̭#�5���`Ӱ�,���N~��Q��Ӆ�<G��-�`ޔ�S'����@�$%�w�1�)Gg��W�t��w�
W���L	d�ߠf�[m�m���{���s��x����jE�g��$���r�<�}U�a�R1�Z[�Ң���:���6@MX�`�8
��/¤����t�A�h������~w�q%n�m#��� u�n(�:ǁcQq����M�Y�R��3,u�w�q��'�ȴ�(��}M�<��F�])�2��TU���@��R�������X��`�^���=]�@�/ys��{� ����+��~ �Ey讓)Ht���]�N��U�r�P�h�1�`l|���)Ui� 8�O�!�Bs4VN�f�􀧔��,���oG��M�&��K8�ӳ�}坠Wg�Q�^�c�fIY���qHݭ1�M�G"1��y����^�yu��%�ܘ�A�Am�l�6u���j��w��aB����� <����B�$+�ê��,�fBV�)	-xDd!+t)���%,�K/}ۙ�;�L��hz1��Z�d;]ʒN�8��q�'�2����zoG��Wz`C5�q�V���?;��0����\���YH���X��(r�Opu�ܐ�7�#q�/ڑ��o����M�CB�M�#{�&�=��E�Vk'N�_��/��Ԯ�OM6��������S��;@������w�ZX� GB�trTT���0�����U��%���O��2z7�Z|�6��H@b\�����铷�:6+f�%h��g�B��7 �a���X^XL
ޛ#����Ao�בc����C��ӹ�o�� ��L�1�pE����T�L�FY�C׹�iItuQT�0!$���e���jhY�B���E7{5��9�m���ԀHez��bqjY�C:E u!\78�xʞ%�m��� |o:X2`�a��� �G!l_BߜEcZB���n��F��n�5�1�����z�5'b�/�g��7Zq��G���2ƾG}r���f��nQf� -�ɦ���B�6s�n���'EN� 6�z^i۞� >]�D�}������Xz�g�F��rgD�7p8K������9��{��[��2�(�!��\� �ip8<�I
u/yN=Ë^�z���`͈�J�1�yJ���G�DӐꍓ��:���іr�ݥeBC9p�^��ˁ��t��ȏ��ܢڬX#�8�Em�3�^�@R��3��SYS��S��|'���C����}j���KnL+��1�>
�������`7YG�i3r+�x�6��L�瀵��	7)E�}V�X�4������^ Q O��<_G���������ߓ��o逻��b�ux y�<S(�]�����(횋7���»�&��d��6��I>xٹd�\~�~��>Lډ�/L�W]B(����˘%�]u]�2�t�l*�N�>`R�e �}j�nr�0q���=�o��ھIU��ݖ�`'�����<����Ɣ�'[1첽5����������<�S��G>
�k�l����<AR�?�%�I�`)�kZ9GDK�LߺT���H���I"T;�)�1Ţ�? ��]^�u���'�A�>&����Ot�� ����m�?���Y@�$��c�;�[Q�o3hG�ǋ�3d`�iδR	瓫��~)�9�Q��_i�d��JE�<�*�leM֡˴��>���j g.�$NRC�Io�������;����>�� D�\�C)p7���7�8����Z�i ,O�Fa��7K"�i*h��8ﺏ�_m�l<�bܑ��S���]��os|(A�����}���6	�$w���O�"�.uǃ��r�{S�jї{���B����P/�N�l����r�9XA��j}���X�#�ܝ�#WZ9~�`O&���$�nV�� �z�M�E���7����)57��q�lه��(oWw�c �r뗁�\Ԩ����������|Q��O�=����[�8�Nm���X�%.�'�="��.��������H��{�B�oFT�H��ǆ���fb�2�c/�l�ɖ���AL���4[�X'/�H\�6� r��)�����	�4�:���n�T^��Qs�ѩ%���0u��|�U-�^�� �qО��)Ӛ��'�9߁pB�~�~8�)����vqsT����o��Q[��,F��pi�Y�9���m��Q�w2|�d�
 Ù7�(8v����X��T>Ɔ(y[�#�\���oR�mL�)[�G�.u�A�x�=��:�JL��͢P�Q���ڵX�[�[+s-�N�*H����Qb���M�a�d���R�*?ݩ"I|�h�y�տQgY.�O�-u2)9D?���hp����ivvKk��8n�1F����w$�J��m6ՠ��U���ȳ�1J�U`�y؋V�C�>#u���;����JLز��=x1q����Jk=*t�T�C���8��3��jw,C��vJ-ڀ{@U28ߎ[���[�=a��tv��`;�芖�"�`:�]XNP,��	{�<pF9�T�b�'�𸝦sdHc4��(`j~Z�����Y���T��M��)��SE!������Mn��T��2�fD,�MZ����~N:�y�[yu�Z��Vjm�<�s��}�U�N�C�l�#���J�L��O}-z�c���ՙ��.�etL��j����@׈��|)�u�zgO��D����3jb3��)Y&�2��8���o[|�pb5fVA�����"����'�C�wэKo\�6�AF���y�h@�]U�(i����,ÿ�����4�����t� ����]�D��2�6����#��-6zX%Ɂfy����c��V��e���K���W�z�47S�� l����V6gT��g���+`Y��iɝS�(�~�K�>\���W�{;6v
���慂Dݩ�N�S����aw%��~��Y_�!��\m5�r�׈Ý!��N3��xC(V��L����TY�Vk�������F�G�I.���֭������Y�\D�# �DR�:���6���!J�/za``J�:Ub*>�-�(��N�n���G����}��z�(!�J�>������!��
ƭJ��!q�j2Y���<ڙ�C��d1�����0f��`�9	X�����E��5�aJ�3���Py�
KTSYSsT�jd��#��\���J��} M/@�t.=\Y3�ȥpWU~��M�\���V�q���t�=50 �׵�!��~n-����Ѯ\�w�LS�[	�]�<����H1v���f�>��Nu��c/�i��ZL���ժ�R�6��E�씒k�6��!q_:��,�|�Eoq�Z��� �6� dċ�m�6l�M��{�\����B���d�NGH�Pe��N�&ub>�\I�
�S��,[/BƐT	"�KD�R~�{(�+y�6L�Q�&3��zh͝���Ck\l�NM�@scM�)��Ҡ���9J�)����e%0պ18a���r[�\'�st�Oe��q?f��L�rI49�G���4$Z�YM<�G��']z��K�0��[>Ӄ��?G34��'�$+n��?����@�V�{n4����cïm��g��?[��1m��z1	�ц�����tb��E7`*�}�
�޾nǏ����K6�o��o�m��#�S���D�� �����UY?N	ODbL�}��9�e��T(�ӕ(��d>k~ ��ܑ�X��KUt��DRRm�>%~ʁ���E��q����[o8����j)�-]��VLQ֎ZT%��y�lu�d����Vd�n��Pf�oV#g�X5�r*��y��b@�hօv�C�9�_sQ����.����Iv�w��������er������u�&��h�,��ły/T���\�]�6`��ߋ[$fi��z�z,��J���,Y����������q�gi@�"�QRw������Zو��c���hKtO�p�FHFѻ��I����K+�r�$s.x��/w ��a���E�ucgE5�2�"�j4���K��Y:����n�Sl9�l97�X2�G^t&�O}����y:$ ��<�7��4��ȋ�\TE�e�r(�}���]�'9l��~�h]iT�Sa��c>u��M`[?|0q����;M�4�E��ԍ���ϑ]_��B�d���b)��}�����L͠�.����K�G�>�TSg�$�	��I��%��a9�?ҙv
�4x�����R��¸��^��܊���pKa�r2��1���,>!��b4�@g'+��p��q��GS���mC􃑋��'x��r)���4���q
���.�K4��4X�.�`�g�0�M]�_L�
yS���w�/��=8��u;p�`���^"������,��g���	���&4w� ]�׊��H��IN�!��w�sXR����lkw�FErr·mz)��^)PI9�ɛ� �7wӉ��TO���}sق�E���-�� �ŔV�,p�o���gD쑖T@���2)i[N�C��<R+�;rZ�RC�jK�q~#��y�Z;�>��S!>v�f_~��tA�}z;�er��dl��siҨǞ�=�fY�CyR�SU��"y#��j�����l��}n���%�N�3Z���^���8Q����vӊ�*;�rl;&��x������?ذ;�E��-�c~�;|�i��c���୎c[�}�,�P��9� �m���s�lu��Gyg�+?�u�<�'P��]��JVP '��� EG���~[gwq_��"]���9��W����u���E~4��`�G�rpkLO���|^z}%k�ś���&�{H��j�����R��`�x��("��F�[���8ف���o'V)�~�!��B+k��|�ٟ��.�[�_�T�9`8�ɲ*K��{��9m.R������u֌��mo,�U+�^N�p�|��ӿ�ןAc�k���m)b���X������Oj�H�_P��}Ċ��N��0�l���o�0�j]���5���?Fd>�]��}�T��#9�ݖ�.)�b	���(��-s�=��{c3�@��>�tjIGFV2Fϕ �y�%�M�)��_��biUN��T��-�7�=����Tq���Wn�]Ml��͖ �x~ͭ3��~ �1P�uCB%c��}w��>$�1�}�̮<��g�=��o�ߢ������Hہ�Mj"1$���=�c|��+�J��ۑĳ��)0gWv�qϭ`�\ 2��K/�M���,��g|�ߗL�<�_îF�*B�Q6ZC('!B^�y,�v����{��F��@ym���4�Y��GT/�W�B�ĚPA���D�Ě�i�P9���7&3o<�>4ʠ���~��s�D�%��r��:,����D���#���W�z�����W��S��=(s(�δԢK�U-�ϸϚc���u1Tz���R�K�U�9�P�,�baW���b��x��hW���J?��������ο*�F>#iT��=OOHV7��"ع�q]�c��D�3�K����_Oôϧw����Yp���p��"��9>o�	jF���*N�����7�/�h�N\�Z \�F!�b�:�9`p9���؄鋫�+����i��b�M1x]	�9���[6m�Ɠ��*W}���_:�h��wQ�E$s^4��~��H���N��#�_Ƕ���"��
ާ	�Ѥ3�&���/�:�e���%*��E���%��{L�&�I͐���z�J�@p��F6��آ 7�K\�U�|��CV(V�:���i��I:��0dCվPA�*v/�\"�|��P�R*��~�o��cδQZK&�4�{:�ϋ�Gf���J[�Bfݴ蟱�B��C`C/�'�X��ZZ�_�ܦn�@�r��Z��W�ޯ:h�p�'n�Q���u=
������q�$�Q��.#�s��X�Ӡ^�Y*'�H�Jw�9j�&��|�5kz�jr�hd]k*��*7%�5���H(�j'���ʵ$�1�:��[�$m0;��"�d��rX�~���Mj�u�~4
jF^������-_d&�-o�:u�&�����1�"PuJ��K�,��fMU�|��J�Y�	-�0�!���G�o+m㶅{�r��sc�Kj�;�.����]}��3��אz��c���oօH�UkF^�v��|����ҧ8�3�&O_��H����%F��ͨ,�UHC{eNʶ|�"���T/�D;���{��ѻ���Q�3��hH��^�I�PPېn_H��a���x�,��QG��%����P�*�
ٍW��N����>;i5���i}hsc��X��B� F&���qb���$+^X�B�i�h�z���Q�w�B���=s�!��s��[,Pw������
�iv��;�Ji;�9�'=T*���Zna����̓A������	v4�����Ϻ���[O*wB����U�x�S|:
�+�
Oy�qY;�"�j�v�NZ�#α*��ձ?��ֻ����3G��D	\z=!�(U�f9e_C�v0����Ky��<���v��
�����~Csg����H����=��?Ψ>�Zȸ��:Y�C	?�M��#_����9��ݡd��uYt]S�M1��I�͈��f�3X-$K�\u��F���}��/���R\���#�n�>l������[�~���|Լ:`��3���`*<rV�Ų�&4�v�q$+.�S]����S�1C�GQRsnӒ�v�����i�����~ ;q�*�2NPA�����G~$,�y(���vh:!w�1���)�sB��}6���0(-%�B7�I�E;tJ���<O�F�������ܒ7�n��m�M�>�w0M�V[3������>-l���i��JE��V�K��e}d���q_%AmFD~UR�$tc�(��������{��ßRӪ��Mҋ�����)雡6�;i�X')dtj��<6�lO���| 9 �Xѩ�S��wl�p2�MC�:�q�K�,�f����¼�
���GJ��&�q3�S�;ߩ[����%;H߆:�9ĉV�y�)V2!���`\$2ˋ��Ьx���D�j��*үϣ%����Eۅ��ײ-$?9���#ө�ȣ�-)���O}�M��T v�T!��(��
�v*��״E�)# �M��Ȏn!v��y���6}�^��/��f��;j���RS�W�X6�Q Z��,7�@EW��6@�_ns������qʴ��������*�x�^IV�Lw�j�(�Sʓ�m�B�4��?-�ő�=���N�nƞt�f�D���Ϧ�l��I��Xwԧ�P�
1�F���^k��Q���k�L�[��5�Kx�I#����οk,���#|�<�0�;�;��,C�p�'5����[�*��Ӳ1}�t(s����T>>S?S/�|[Ot�;oM����$V��%+s^�LRv�\x��/�&u�h����P��tI5�U�ܺ���epW���.A�s�v� T�{��yy�w����k�COƭ��]��/��g��jJe���Q�Rv���+2*�VKXfAU �#�h&��ٰQ�BlnBD!��;��}>4L�M�%z
m��I�ȣUq�ٻU�k�WU(�v���8nz��=A�9��>�з�t&���HN}_���2���4�v-��y�u¦>ƣbݵ���W��X�;bO�T��|�崱jiKsۍUJ�;�zH����7y�%��T���ZոTt��N_����*��~]h�;)BX����Ň��d�9y���&�n5��ݠ"��<?]��x��5������7����֐+SMb��7<5H�I��-���7� �ҳNm���Bx�r�Kܠ�~b�q,�V�Y`д��1Z:	\!�����B�E1T����y��4�$�s�E�O���Gr�b@ͣ��-������T�g�_hK7����hiUTy��E���c��P���0�ja����NFF����ч��䨾)%r��\ԏN~<��N`'i%�=ت;Nog�M�ԭ�`}6�DI��\	�vO�A�� �sF��x7�#/�����E���]�8�@���j��D���Y������idi=v����5���������Q�y�l/���ߜ8ؠYP�;�剤�����V#�T�>�a[�:
�9��\Fb�u>_i���i������e�tr��ELS�o�	�ik��W��6��7���*�u�/�[$�h��'�g��%2�Մ_� iΊ&7�<�D<�?�}*���U�R���(��Ώ�IT��+�ˬr�.$?u��x�UI��Ӌ��^�y���+�pg�1<([��K�"<ٽ,�����a��X�ֵ�j����I����D�q�����5T������x8�X�BȨP�&\M�� ����Q��m߸�^/w��J!�# �������س�`����M��Xt�KФ�~�ꌙ�o^��)dYᷗ8,+9���ڌ�F�*����esJ\��d
�O�3!�DT�ُs���+2��;�J2u7�6%�ۊ�c	x�(w�I���^��pЏڞD
���&4g��R��R�r�v Ի�h=!h��;��K*���駫s���,Y���G��:u�H�[9g���ەe��Ӹ,h9����T��2.m)���3>���O�E6D�Ii�an�� 걵ŭ'պg�YB�a�z�_��{��'�u�c����歒%�R��� V0����2�`E_<ȃ˘B�1~�7��j�M�xb��!o9kK���B�^��{㨡�i����3���4h�*KLr7-����a��`ƛ����o%�IA��B����}T����<u��i=O^�'�h����ԍT0+]���%���9�I�����W�W����]��$�6�>�j���ڤŏ�����<�\��[x�.'"�ؑ�^p�e���B5���K.�W�rx��y~@��@ß���}>�C�7J�cC�l�!��mUe^�t[g��z�f�T.A�ty��=���v��;���SnV� ���	�D��z?*İ��PN�����/���~�u(g��	�Nk����SϿ���_v%.�e����(:8{�$G;;���j1��W����:���L�:3���}�zD�v��ݲ��oܜ�Nr�t@ eX�=���E�2�1��(@@0o�P��e�a�(��. U����b^P�fy����� �t��*����orY��Ԣ�&�^qJm��T0���s�I-�8��J���	�E},�g8H�Y�h0�d�*Ɉ������Տ�X e��y��@5���{L�]0=�U�u5d��F�~�����߀���o�&�����L̡!+z�(Q1}$��I�^�Cr����s(X9���"^�����-����E�<?���7(��zD���fJ{�}�4�� 3g`����P)�4�J'�h)�#~҉U�=�%bi�qP�k]
�T�5�T ���Zq T�ӑ�N�u�gc���������;�af��� ���� ��'̣�e��!}�/6�ʆ
N���U��|g�YUg�rh�M��z��_��/+����+�����嬥?�^���L4W���P}���>[��o� ;�@~��,�7%L&�۱��M;���-�b0��a�4bd��0ī2�]�Ӷ���[LHnd�,�]a6�C�����k(���
��&��R���(A%wK�ٶk�C�f�D=���|j|b^e��ut?�Ί�5'��Q��,o�:٣I	��ݴv_h��u�p\����
"�h�c�:#�쌟\���ܣ��Ë`�i� ����ymG�wT�Юy �k4a	yt�N@X.2���Vf�9�ٮ#U��k i8�P�m���J�S��v$q����O��O�*���?r������Sn|��� ���m	��v��+7��̘����IG���b��4׫㐫[-��Y�ø��.�����0-�.�>ʆ��Q	kU	��h�k��)I�7Ej��>�y���Lݫi��k�;��R<��&��z �>�zc����^1v��ȷ�E"|�5��������=5mɐu^,�00@L5�"�Lo�!��[��ٓ'����M<)oXn#�X��ˆ��xM��2#v���\�:%&���#H�H���<��͝G��?5�O��ǎ��:G�m��`�u��a$e�����5�ϒh���¼D���~%�a��<P�[���t �('�m��Ct�.��<	�S�>�W:h�����[߫n@�Ϙ�2w�H�o��p��/��d��2�!Kw^���m:�J����+Z��w�Z��������*Uc}0(��"��%��x>U\��"�R�ܻ��Bl\�5�=�85yR˽ɖ��3^)�3�ߤH9*�/��!űJo�+�R�q?͚�{Q�� �M�<L<T�^5+�h3Н��'���YsT��V�Jw�g+(�����듥#,.����O�`�2�Y���w!�;A���N��¸�O�i�l{��<�s6'G��]C4��o��a��/2ƴ������� 7PMj���Fq/��f	����m,�1I�'�g7�� ��/k�~J�Ү�wL�(野�5�E��P���K�ß ��y�g��"��)y"L��Ǫfm�x9�N�0���=/%'f䤙d��RsK��F[^�X�пz�SyИSλ�o������d-�s����s��þ�K�R�.P���ݐ&�j{���Aڒ=�R�yڹ��@�����f?C�}
N���~0��-��&t���h�2قV��X��t�xA��O��:<�O�a���4������J�n�e|��{��Ϩ�B�~��6�A��"��w����"^
��C�5��K�|.=�͕���4��xفlu���A7rv���8:ft�P�P\|�o�'�&$���1Ff��*�� �~��C��(B����{���`B�=��c5WGa"��x��s��T��o�+`��Y�_��H�=��������^��"���/��c����-�.�� S����{�>ž���{��-��#%3��Z�Շ.��*s��r���t��[e���๵$^�f_�;d���jG6�B6�/m+o����x@.R�Y �N���1��!6���w�4�5@�����&���Sy��(�]�A�ۦ�2VQ%���jIJN)����Y�ku�c=��S4��b3j����4Pd�ᯗS��ةY?�\
Ud���)�~��sD� 7�C����"��/q�c����f�J*"������r���#/HDav
�%'���I�|��@�Xޒ��Z�È��Z{h��������������A��~x�N���s]U�BK�4�:���]���&z7�������>�"�n2趂3��Q���h'!Fb�5��zK3�h�_��n�|���~��2� m�a>���U{�"��Hq�E�� ���u�,�ӌ�g�`B��9��(���]�c ��I}��&�jH\cG�M�|ʵZ1�"7X�Ef��2��Z��߭gW2��c��'æ�@�`p�A�>�=4g�~snsT�{��oB�U�
61o�:l��G���˅h:R�_�<��gcs��w+v�	��U��>����~��wX��<�4R�墻T*�0a��G!��9�J���,Jb�'����ȿK��UyO8p�j��G����Z�kF����������^��HԆ�� �,��i }��q��p���'�ѠS��&sC��1 348RxWY:�����d ���o/�w�'+x����]p;Q���2���/���E���c���(OQAq�c$C^|Ç��x�
rd�2�Gy)�ϓ����ԋv'�B�س+C��3���u��S��b�6�ALN6>�n���g�/���#�$uLd�c����Ɉ����*Mb�H�
@�,�_X.��z�f`]C��#��a56r��h���:���v�h�9l���m����A\�JTLo�����y��!��˴t���;wH�8{���_�D�1�>�G
�?�>W�����E�M�)�N��;s�:�\�R-V�_�%ٓ��^k��I���A/q��=�8���2/�_�������-1���#/�� ��;~�{�v���G�9�s����E���:̎Y�	�l�,�0�+`��@ �T��9�nƞ�����!�3äY�
I���67��;����E�.e$m�Z^#�{�gh����gSz��.#�]�+>I��(��GNS�b�{%��>߅��C��������z�0�f����L�h����>����.\Q�����ϱ Q�m���.��=����ð�G�����䯌	N��3�1Ҋ���YL�>.�����|��4w�J�T�պ:S��%�1�Ë+���H7?�������v��dp���t�U�չ�U)Oñ�*ھ��m������D�j��'�d}�gF�"� 6+�h���a�[Vw�k�	]3e칟}�mG����ば�뜭^����ޱ×��Δ�u��5�^E1h'��Pd���`��~	:�2Ra��;�����Co^C}�QJ�?��Gu|���[�9�q�w��v�)i����+Z���O�F*Q��h[n
Ӄ����h�Q �A��^��QvH!�oFQ8���|��%��D�q�������V���h�*P�<v�o���s�tД��18����:�D�$���$R��m����Jܭ.9�/�7���N�3�h6�֨&a	�R�7���P�N$	��Y�13l7�֢\��G���U����fb��Y���2�o�oҍR�w �(5�k�0>�,;h2�U�ͨK�kH�}��`�}�G�?w���*)�a\��{�����{	�yvN ۊ��~�$�;R|�D&Л��
�&͌�υN�����E��ؼ��������D�K��o�Q������p�0