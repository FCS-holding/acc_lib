////////////////////////////////////////////////////////////////////////
////
//// This file has been generated the 2020/03/16 - 11:19:27.
//// This file can be used with intel tools.
//// This file is intended to target intel FPGAs.
//// DRM HDK VERSION 4.1.0.0.
//// DRM VERSION 4.1.0.
////
////////////////////////////////////////////////////////////////////////

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Intel Corporation", key_keyname="Intel-FPGA-Quartus-RSA-1", key_method="rsa"
`pragma protect key_block
p6WixIvdweGqxn3DusGaAJNq765wrL9AwTeyUeNFydeciIFl4JvYwz5oU0/libRvK0IuRxmbKEQ7
+4grSDAbvB67J2w1GD3KCZ+bi8PLJYOzrjq0U6ehFnR/mIf1u0mbviPe5GxVma/vox+nLfEzylDd
a6dKqbB8VnfDs9XY/4EI72vgwloe+Auw9vvLl114EVw/i+NEWEjyPf8yBbmU67Oeuodh0XXtxpAT
2dwOvvIY2pcsgojzxDt147lAmlFtgUS/66Cs7We1BdMeJucfCsVYVIsXfDrBn4hI6dP+30JpY6QW
9Mt2dAoDsCUugjINdVyBU3H1sIG52EOsLmnT8Q==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=20096)
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
4AQ3WifCp9k2q4hM3mMXdI9PCZ30cOLhBgF+dCV2sRmAIWc5XMGiGD4vbLLOs47Qhh65aQOI1qiE
iEiivR355KWJoI4/+2WTCOuG44vs6dEjet05sW7EmrXB5nt1NBjWYVEOyuLJbu+P4Lnvz4tURmYG
/SH9CgvI08Lh7oPjdjWcdabfapRzlIPBoCCo4lMTUoT0Ve6qUB/gyMJAu3iI/ywA8zfI5mj+uWH8
lz9WT1ffgPZw19yVYpFGzjAqBOBL/0LBxZh7o1N70MXvsDk/H9KCeTZ++TFH06hNFRndltmHm+C+
0UfJpX1tXhuP9eKYQuhhSzQ5xgnEY9TyqduYL82/T15O5EjBgl+Tcp8y2MFiYVjplH7xTXqEqt3/
VlCYC5d6Io1cSf2Pvl8xVeyO+o4siO7VrnCSD8H/6AWxbhRRR5B/Qv/shQnC7ps95iLtvPdMuuwN
TC3aiiq85btBIyCJ3wHxjlxXr6YIlh/Y89X6Qq75XjyQzGwFIa7PsWtABb/+L+SWAkjPTtF7azYe
lWuiceWmj/JpHKVmVyyxekQLeLbdd617PujADqjiflWMBUxHK1YfWXi8dLLyJIjsq+NRdJCuthsf
FLQmIRElnbG5PZQJ3s6EDU49ZtR8jF4ehaG60i8VpcnvWeDOaT90d7zFFO0bkF5XmxW8BBQJaVQh
sIdN54s+waWXZb4jOB8lccvS2FYppzzCX5Yx8+2DD2jO6qj3RDDkpkglYUM4K/zSBdSriOAVYR95
fRjFyziF4uopiQScHHgzRPLhvQzgPCfHSkF8BlLgzcGQzkDoNPUm52pRJEbh8Q8nmJbQq/kAmxKp
0+Ngt0cmeZo3r6vkDNbfpUCTt/ja2z2vfkUEFdbswf4XI5gzBMbSbUFBO1005HTkb9TOOwHQ4cQP
VSS/YoXy6oM6yINYRe4slpSnwJKQ0C8a8jZmP4j11bWrji3hyFZl6ubckOsDiCHYGTbl/NailTYT
ADSeJpiXSpeOOzldDENPku2QNYeRNvG/YPNIh1BQG5oAgzoRZVUsRF1Eg04jgUvZjuO4sOqJYmq1
YoXizqQRyZ1ZX5MF7m2ykJ5vixEbyV3qGkcB+55DJZDobc+zJqmdSl4n3X8WN0mh9lI0fRQFZl3d
M7s8h8qFFbslzm9wzhKUFE4Uo6GEiJx4mSq8S6HOpcMjG3e39ChX5u8wVwOsNDz5Fx+Tl99wPCEv
ja1CZ1ep6pj66Fbgx/r55KQa6X4h3GjfCB5hSEXFmI0IaTalhdYEOJiFPSZwLKt0k884jBxtkIcf
fZtasgB37/Zs8imlfEWRf2q4Ns63psDrqH/TBSY5dJMNBkRsCECC+s2WMNbJx26G0bpn65NU2BAV
SXzVjkW32AB+5n/dLuNNf+pD0/QnkCgBE74yzEGXzAEfuyl3G8BGI68hDHhIhLG8H+oGsPNvZ14+
fZyrrGY5ipxOkWicp7gpXe8wmn5HWksMnEmhge9/XKbuCLuatF0VN05XnfYiTMhbmXsVdniUJF7Y
GQiyzhEewd61cR7bsFLf5Q5T1NWqVS8tof51qIA4SyBbcBnn8OmHP0dOVDWwzRs3VcqokVL5oQ8e
cNNIQ/sNFr4mfFUr0y5gaOXSH66jlbFHodz7o4QDiiF+6tIkrYNSmq9NGrMQLOe1iZZDsCm1DU9e
X7EvE2bgqH2imgrW4vwHq18aIhVYxoTefhZ3irXnT11hLILeuwabVqYI1+I4/nIEeLUM34FrDwSt
KgteApDzJp6qiJQ6rnDqckwgHZ4YnaK99f3/caqSFlx/rXi/IIqUspxUG/dPRG7C/GHItylqqx33
pJMzKY4NNNV4vgj/kd2vd3McgZEo7CtS2UDp6eMrPHkvC9FxLDCbzHHYUMuA1VOfjOOBA1IF2JNd
nk7CwWJYM71qheLwlUj/pJVgagArm1D4ViBn88X7/IQuxQOq+Bt3ACfL+P+/XL49pVERbbiiqLtu
9ScQcsCq8ZHnETNKKIiqrnB5msxvBQi+gbt0cedl/H6Q9Lrzvec7ycCYh/+Fuz5/KXdAutJmgvRG
Uc6axpNL+/1CLWE02ftPjlKlNHKAq3Dsab5TE1IS67v8fta2bmQ6RyZEme2s7PewUvkYQBEd6Ty3
Mz3+B/ZyFF7et8ravGTBmB2OppGVs5/Kt3I2/x7G+E8KSsERaNEPLtOVR4QldMVBP/BluJ+awale
9QKfWufOmUcl7iVV2YHbjH67or7UEFKqwDvKj/ZKBrHeau2RwpGIPt8oIsf+UIzx2RhHBDbRgAeF
ynN0WCHae7NxRZdL2GDhbH2M9lHNSycnAAw2DKY+cIhc49s9gjOsTcTVKwvA83ZAChc+BAQSwcj+
zJLHNFbDo1LLnnS7Yh1+NLBAqDJ0laYVk5xiMbNQTuYPLBhGn7fBm2z9z15Zp0DiS52nihZ0pb1q
eNCPku6OQiX+LwaPcc2gk5dFray/sGCh35nNEoJd8fR7vefTWbLK4wT+w1WzDAkXlmQXptoN0fVB
kasoLsv1bku+wqky5jLmT13ruaaiwbijwpgMnTZr2ViTMg2uowQaxj7zQEwYaiZ9A3U6/CLMbzd9
u1NwGIRIe3Soe9ADCdUAtSrCuVCPFg4E7mk3by9ziVDGuAqPlCRxXznjcQUAPVfZycaq4x2fihRV
mQUtY1OCMwDQGOh1st75YW2He3XLkTqMlVFF9xXSMFVDhiiTUJyKhE3wFtTz9FiR13vmyMD33bxG
FWjfW4cj5uMIowL9pklk1q/00AJI0Rc71T+KzKrYuw0B14hYnkM/Jne1AoZbADC49d1GupqqHtgk
o702lCXtFGF+Xtg+r3Yy4jtgiPU9z4iOp/JeaIkzB8dLUPS31w7tEOkFIR0OubaPT6yJ0BP4PAjh
R7/e2c2guC+ZbPCMRjTR7IVFC1Tog/xJMgLsMli5jtpER3yQumUOc08fV/EvApk0yiw5YhOPoggc
di7E4lBM5yelkk0Ls8R1By0Ctyaskuxu04JzH6RpyoTRjXG6WgE9fB5TxEwV6df0zWNxBKnb3MW4
2nn3vI42JhIBKR7Jj3LgKemo3D5UCTZlH6IX1JAXv1lCdAnoXAQTUgscAe/j2xrFzPHWL0ZqPteA
1wJ9tsAQIgwFBvR7XhUfY00ej5MsRoU4h85g2aJSZHaiNsiGSwqw9q76eZLh9D/EYq1ZSCxenIdg
Jg9PiRzSOubTdQ5xcnNTndxlM4kt1DuWiU7c354Qc+GJhiA1xeQkMeQ+j/9TMVLEmvuPqg+Aq+US
SxQZKxiwF+i9thKAvh6ER5UqJl1oy5Gf4jVbla/UJOMshD7fviUsTjoT/GUZ/3grm0PIxn529FaH
CMLcglI8Jj837exHD+MDToQYhe6V6JmXe7EojN7lbb8JwHEYE52Frzo+Q6XjKAA5q5qC6oMbbVnE
1dIkt9Sr+v/OyiBk2rNyTt4Di28F3ySprxx8rQnNCtxNKs9koMLpn3uuD+lcHPMnv8ZWJIYP+2Qj
UzrzQRynHuJoOTQ1/j6KCymhmuqE+ZvFUCJ9vjIaSY7rWtFonCtHvlXSXr6ybEj125v2t7ezpioq
jXi5/VJ1h96spsLfyU0+x8bpUR7QZMpdW2Ap2hrF0HFuHm5jUlb+DCyJ6SMRvQVl/qO9aFHF8Bcb
KNgdbUGf/gsQC3h9yfmipVDH+Ax+JfbmKmZTpvG4j9CfXq+0iqEjzLgG/7DIfpB5aUJOnGDNm5mE
3vboSzISTncaOFBeweSi8xHgLU53FDrou2FRx8miyTS62n0gp3/VbnlVQYhfh0idg+rLPv9eHNj3
EDMJXAwT1KyGs4T0YFkZqbVrXb/+lMLItwMWCHM87uSDjMnQ1CozqZh9f/qB1CtgtEyS8UsNExLS
bkxN6RE+pAbCPuHEPtsiaIN9BwYXdGVZhwshGZan9aFDBRxE77rJpPx4IF036x3PRlseSPkDhwnx
LR2NYKOAvEwhXFfcy2AcuiVD4EU+Yr71ipjghibP77eruY/D40IZLmcKbEDT7/5AJ9gI5KVcKCVe
FncWiMBM7Mm6SNZ2eMzSY//Igajwca8rQy3e6Ebw851lHtJgKseZDWc3pT63g4aatqdsE3ir8UY4
gNw3zxOGE6GrozrZc88hPhSMIw9q941id7Um1ZwR+Jdy2rQxPJWVY4803eG/aEDeqes0bxdeAQ9X
/oaOjEVBsMdUrSX2LhQrWPvgfmGwfEHimqDrqKFHpCCDeEIDqsXIYPRpZFZoc4I/lUyFaq2S+1ND
+sqqwNmytcbSOh5oDPr4Y99uohClVLwg1TZuc3HEzU7stAG6rOj8eRjyoW+YxbcFZ/OHlcva55e6
Nv4aMZPtwIjH5kEHETFvfu9R+BH0wPDP7jeIowUVaRveQngTo2wpGiVnLtAuoAYvoMD5WJQ3eTgc
ewVx1MK240OGYnAwj3C3R9By1Bc460hDEOwz6ebH76/6Ys7QDFYyXF4ak5UYr5/Qcfa9BDwyK1No
iMfVuM6QQgUvt8PTj8Sn2gqIyVTR0sNLc+Nn3Wtbg/8mwmBv7uuXtMWKbTQn6tDCiwOcOilh854k
FV+1Gqw4pP+jyRcJxJt87UJ2VN4p8HCvwZV/mhQ4NKFSaROW3wIwkn+Mm2YXUq6eb1y+T0xgyPnQ
dPLEd0IPsJ4iRhy2V+R1fB7kWITvpleWSKFA11qnbL2jthi/dGbxip021DQTMDHVmukx2kgMUc54
K9iaOOWraxnYC77/3U+bwrR4cvc6xlTZF8Z/ClkUMpByeMzMWLYgOfq4eZ54ZDKyfSvaMflw4g57
GCJrgoLApdKLAXMaxuBTl/nsB0IEaeoj+SiiOSQVs+Bj7ZDoU1bls+9l2qiOntp2mrV0Ow/4zlqZ
3pi+vvCg48v3KZLMgIW7MRdBC+V7DsOsh/dbeukr9yLYYhogVft5XH959XJosiQ0+C+TA//4sV1v
uh9NP+IvOjHjQEuqokayiEAxQ7cL8y0EryPth1nonryfL8B+qFjCsfWULnvaZpTGq8h4JRJC75q4
1Vl7WmQWnNyUsSoUF2+GHN4SpoFWKwTc/fyZB52ctZqiO0urvlwX4RbAMRgcYAWf6s7dTV/aITAD
i/j0qKFux+YRp1MPyup10S0mTB9HYGc1fhQF8xQKfJFNmfRs7bejF0amfPqA6pKRbA6dNgZrJ2U2
+HmpITNv1COY31ymQNKM+QICyAraHz0efXe6pXHagBUII5dxJ7AkhgkmlnTiJSZJcplH6kH/jZpi
4pxxLrtCtuuK8DS8yn1x0MOOlWQ6x+ygsa7sX9AFCm+qMlDX3IJn6Mc8+InuDN16xisec9GTVrcA
q/Qi0DQhsmvklmER/JSlPfp9pQWdsSavy4T1tUr7Wy4fVNbqrTNeihCLhKXC8M8RcxllxCPVU4O2
saF9CWcBaOYrdzBoslzJ6Znzc6i6fJtcedFSGhoTaubpaXU5xU3q7b8Ut56FJjNl1ndbfSO6rcb/
5O4l+wLRsH665xWYhb3p7LVr84xsjhQ8jZH1dD4uauyn7wiFBNz2cwXaHqEVi55Z56vj/ZsO16hZ
VHR+YnmTB+6dcOrw54/Cyl0pYpiFw/VPpdzWgO7C1F3/T6LISD0rm/EQhqDG/AXobTI4p1H6eURc
4dF7GqtZ6fUrCSdbBDo3gHALKJy8UIKHCP5LXyzfWFOIOBVN86dumRVbJKuPkObaMpJqMao+Gqy/
Lvij1zobTw0APxmBuqBPJd68xw1J3CyPEzZJuf2ni3riS9ScJnlEpWkLd9PU6ludE3AWLPCWw2A1
wH9r13D1JGbAF5UREkL14qDEbBhBNYjo/NggGlpF3tJaCl9RwoF1Of/k4w0vAc6niU1TyPHMkEU3
SdNKh6Dm1DwZD2LKKyGpXk+C5Wj/x13VeB218S49//nGRNGttNfINNHza4fdgp+7bfsI+nTX4aii
dyUa9yX7+rd+yoOAVKzmI0646uZjzqgaQdztu267XKqmw+XavYB5biofn/dNg+wT9sjP6ovf/osq
pcY9B1aeHbmWYkxj4JR3/Zno5hxtc1y+JX2WNhToFs00+GpF5QdB0VhmctPtmqtKRQKBBxZBfafF
CcIRF8ViBFQvEC2IaiNSAJCGXkmUx2KPWC8Kf211MYR+uFdj+jJGBkrjqp5oQosNk0PZ3hKfv/oP
sT+dqQoXI1EkFrO8Ly4Yz7XXnAGbhAoyFOklqaGOlDzue3mVYwauVcRtQWeULL8cbz1RGjCr4XeY
ouy4aG5DMq9jogBHnBAdY+ch7N0vFBZgTbikQP9X1NKpjCoWPzPv59+2gty5k8rEjkmLTFmH5PAQ
wrdtOZvyvMzoX4q3gPBYeQ51oFtayx3wJ2ep9Mnj/NYSSW498MDwy/xhBmLJxRcr4tLdm1YHNsXV
Z0ERWoRdVBytkUcbjxtVMxwGxnZpszf3KNjknbfnOVhgRRGls9RFwTK5Y51EDZqJNkUi1c2IxoH8
nN4Almb20Kfp0Seu7r7AoeUpv0ps3/foEJnYm2hVeh+wXWCoAtN5NH0G0r9nel4uHwJHkVJ0hhWL
4qQ2h38lKUP/krx4kxOwsWHh262JSyQbeqDQxFuLhVW24G/nrpKG8p+F6iAhbDLAifmnchdlYJ8+
/o7ykwW1Kge70o73+HHhlVlA0zeCOpkr8yBIq3k8UW/LE9CdTuFqlCyFvtdE3KK3JoDVLeDwfoUW
zkh5MlEUC0zr/D19Vo9v9nszp8Ct1/8b2IptINLSpWaZ24Ex1t5i59ZfCA+oNdLkRlM+4X+GhLq+
KNGZ/eL9zsFSo9h5ISPnwPTaCEoNxcBuI7m70a0uoCRsP/ZzAIJzAABwuyMv57o6DmKJ+ZGwsVaF
Y4mLnHw1Ej4KQDnAkPO2nG1WEzU9eLfLfaTtwuYvNDDwiqe/ePwgj7M1b0h1OTX2d+oWf3gXZ+at
I5Fk/IeOgnETWsoHngzsdkpq2xR9JQ4le3HvcF0bspM1J2IJlx60xuqrQmMXWTbz0n6/Ynepk/UV
H+fmJDEDpTThCPHxDygB1mKecCuC6S4tEOcCsqqRnkEJvIwFDPuxfKTEvwFRFXXAzMsiuDVEviR/
4c9UAmkVvvkEdhrUCwrLDNG9w+YhYKWrz+VHaItiZVq9aobmdnpj6kf3JnqomWd68plWi9kbk5qO
eJ0q6uvG33lOq07zb1fGoQeBt3YD7elisSYPMENdZyDFWhl569NNScFy19MbpUEammGAKgNfljNS
3U+hrcGHnEKWRUdsFdM+cUDqHaKCGo6Y6A7x7ZIfo5/Me2brWZ9C/DtpnAeLGRc1YmKEXVOXz8T5
MgIlkYzAxwCYp7T0hP3gB1JSQus1qQhoJh41VewsRvCmVR97bP1xRbK1J6KuJX3z9ORujCidye8T
se8Zyvmd7IQ+I88EDpYXeBax7FgOB1rQYM0g/UsQU0T4V3l/nbBMuvj7vgo06Gr8MpZMS5Nl7iB2
/3L8epxy4ThlyWv17wHCmGafsNoT6T2aQjRJQj0O5WAGYMlYrygEL+E23t7ciFQZoXH9qi0IOZu5
KGbl7bJiHyfIgA23wNvkfMBbmVxYNVvGcF2tI/1BDFtkgraILjbiv41VfIWWlRunDslM3Fvgq3Fa
rcHWRhJ4C9enniEH5cu1YQLp2TLtPOdUKHZgj6bqBP7NYjHAFb43pXCQW77FpWZLj/zXH7R3gG43
2zcSD8dVXZ2fa1SmdC5W0TY1YfHdeadPsoKYn4qf4zZD/+S9VHOTpk34564xdaryqT7nZ5vr+EZ2
f+Uc7Hv1rir91MIzIAzcOLrfcXKDfrdOxB7+zV7GgbYcWZph4F+tWtTEkEF0opx9AibWMNuse62j
4J4SZg0yI23NOUvzwrbgWYyHEdTcrTCqAFWn4zcxYNIEQEyDqUgcv2OLG8EtfX0DX6nTG4yNeQ5g
AyJ1DUmfYQ3wCu5bmn2jtdbiac943BV7jvt/tYM8bCTUD5C6P7WxBMqZQGxvCjhZKhwdNfuB6whg
BeH50TxjZGnDEYXYqxUkHlZYituhK+UZPDuunScqf/hFQqVs62d57N+SLAckWipckzPkM49by9ZE
zD+A0rrCVx+q5xd3NZtl4CrahqVmrl8+3KhVIuSQkxM5pMxMIvw7hjZHS/k5j2TAeApaGNX+LS13
+FNnIaE/sZrsjDZRq5b6pofS5gqdzbKuj9YbCo8bYyRbzYkgWxlekoJ74LZiXLGTIBbhcMqB9jNQ
FBSIM+IlbHB5UlR0ff473gg1qINPhktFOq0u3kjEgzMisOM9mdf+0FYWpyG9MKQdbO4LY5eHYSnP
rk1lc0AbOiKmZzkqIA6GVyRMRE06dsLzla0utq2VKGSmgR4GNjiVCHD85cVexY/k6L+oYHfNHjdN
eUAKyakGzjONRJp43w/cSD8GZWLbTTmgoMs4l6KSd9XPX4rRhr3h1Yzrqtqo1koQdQT9v/x9IE9L
iPDUiDSjwoGel+0ze+24SpdPobDd9i3iV9QOLosA3rPnF0/yT4rFqhhqoF9ylP6Sjk9yEOUbNPFh
5+G5cMhPFQ+1+3tZkzPwarLaoAY6Cu7ORAU7Tm7lCO059SmA+55KBhpXsAf2mBlTukxjbWYuioGj
rM3DEkP+6MX5Il5PhwVeCF1Rb++8DX2sRdQeSE1GeAn1cinQ6al25Co8bDpYhhoZiL3DEzgszkbr
eaf1HUVGUXlfbjP4S2uD1Bb6tevqtijwiQ0tiBxehBBswRdms7qBMH9yHsKod1n7QV3WdrK+Tg3e
AY9h84NItGh5ECtvusPdaZCEZTIoO1nuHWDlFNKnUwuoy9Crj2LujEaQlVRIntnRyIwtnQX72uF/
gdXruBA7hoiPoMAfkhm4Nf/5nNFj8zvtuYTuPvI15gjDjtwBqC3VzxhHuPRry77uTj1X6nd052YL
FRUCnEuPLxfs/1i4J7WpUGFmXNNPzfA4UpojV10YL3F5OqSW3Fq3KR3S97QBmk0pt64IsOhyXVtg
qOZ3HqdAfSmcPup46Xk1noHHXY5YoCnoTKgJ7Coyhul+b8sUM3yBdoFPg67fzu2QT9osF4ep34fr
GIsCowwAEgIVAgDFrX5CUEGLehcHMwMW7TxX5wgbKOjAGRSpo0WPv/S3yhj2uP66zIOUjuJSmSK8
VLzqL2WtsYMdtZGAcaLw+fvrEfZuHtiQdi5eO/ZvZQ8hedyJTWMvLYP6HPGLFd6zxKs7q6DaxUqt
zzPWHAGp6q4oUhfXbT17fFdmNh4Fhjf5FqQo+nCg/9CnYK84IlzhkWSXsFr4h3FhemksVKs3UrWn
bSIOQSpQ06/yFWghjDoH/O7oh0nKnjKCGbafZ9ZW4kKYhYjNRHtnxJOsIaM3j0k52bYCHUaY6iK0
CoCpbZGJMz5vCHmZBDhatlmxzv7Ksr503QYHg5AtjXseIjeZvds4y4uky/nElltmRl/mt8tuI3sC
VRgNf2DBAtD9RMGQ7KdCQ1gFM1AlSDi1V4Zzn3rXmdjCmPp9mIY2oXqniik3IauxTBVVdlne7nzv
0C+EZZpHUFKcGt8b4WeGoI3ghTgA48rLnzQrMGeZutv34OKB2OR/sGPuasRsL5cKeNVW66/u3OO0
z+DdtLvre+RbqBnhBWVUZd27/NU2ep1/zaQ1XhOPQqVDuDRLKLFrnD2QrENyKmYQVmu6DIb2+4sd
KGLs6+nTlgYI/L2GHF1QcJ4wZh5bfDhUrS2fv++7lRgKLFc9tMV7qOFAQeHgfHkAmzOsOZWWlRgp
lQXXRWoMgJIJ5ahtyon4i2f0wgKRjGTCsWIEMICewHRm5CAlb3e0xwEhZCcj5M/ehgO0QGocnSzv
+uKufubLTmI8VIGkm9fSPExQ6sC/r1Yi4hC+U0kaMhQlDo1ryKDS23pL1whZhdGbsryPeePKXkIl
r8iv4s+Sge2qd02U80xA8WYWXoi8hffTOcNozYuPDWzXmE0TfMEcRtP6J1vw2HTZMv2QJreijAA7
ev+JzUhcJk2ALNX7GfGLU6gp4K5b6Us/UTll+k/fYfyHrGIz9VzYbKr/nwoRgwTlJqG37d0Xi499
HOdV3pqEfPkGn+Eslfnp1sKI80LoZAYyohIG9X0+Vw48euN2UlhWTym5LUQKpF86wx++y14PLtvw
h/hVDaQy6SD332nFVWCQTNyw3gObUlx5w9KpX7MMPfCSvaUHz2mRizsa9cJzANYpZSg6juLfz2sY
V2HyJmMX82dYEeuXSqkjMA5+mGchdhOxRwhaenoJzeppcmgao/q572wvwbakzB5TZTRvUiz3OaBM
tB0zu0wWlSNl8FStASnkVYiDs3oPNTIqr4vFbprsmp37OX4HofubuYncR1UWI/a5GsH5N4Ub808s
e+jf84Icbcv6AYBhFPKg3xXcun4FGkDN67JS6W/ZxBQuQzpRzRvK+4yZVeMJ3fWRYVMv1tyJssaZ
SsyPHVs4/Zi1jgNNdmHHpmLQ7KzdNirtbj1AggIK5D9cViIOa4BNvmVbefUiRpkTkQdaTPaXYA1g
iqIEqtmOt2IgsljFcj6njn02vHhD7xb6FZ+YGcP5vWzv+v467/YgfGsamobYJJaEfZfASqGK04N7
u4EvLpXG/Yg91a4sOiIMnWs4QWPUnNh/rGzuXxpa6BXVfbBSIzpcH2z8OTEmOzNODK+PPUvaIGzs
LSCin9iUdL91OyWx3Rajn6VYuXpzABixBw5v7H6K2L7dK8hwVQ6Ow7vOQpvAfFq8O9v/Ujgc3Baa
huVaHy/og8aZG3YxBJxalm3tgx8OTWjE1nADJ7lIwn0/8Ld56MvGOLOmNJciJzBn+iak7O5dlzEB
EazULzJe8lv3DQDy7vgFOzvM6M7UV6wgHfScu4RC2Tnl9j6mbdEvPnMFln/y2KFWsVdxfgrrU390
uDngduAm9j/KMKHEB/A9+ar+Om7v6Hxh6LdxSXu9wE3mgCLzjTVDa8qa7wSL7XHm5WqWQ7FMrBJs
X0XhHbV0c6jpq6HP0VfRes4oYvHHm0LaV9vp0GXCq/dhJkjbTwoHjd7MfBfvzFqZkhnl4nHbIxps
Aq0nkeCnfj41l6GsDAfMNZN4pY3xfCcFLmaikmtfs4IVJfOah9YEsb+M5pPL4bEAzZr/NBy8LBAp
r59KgSpHhMgGZ+dUigH/mHGNKvjHW+hTlPFAWgO1oskq4RiJR+Z96BnU4nQpqqK39PBMLLjNQgec
1ayqKxJz3BwYGNDRP+mzFw4awfWMvKHZZRyHfgtEB+N+Uxvb2SOMwgkijhQgyY1PRiCiODIt1Oui
K3+SYdUj6gXvsVclmDg8SeYM6e76Uo94VxHJUBbozrIEH/px1XlPu8I95jziUW7Q7SHWIKiUbiwy
kCODE61j45S1ErQQxOfSpxwR3BA81MBAKFSUpTzCAv3n3z6Vmutcb0QvEpKYeq5RwAdXG2SpP8E9
O28Un98TM8/OyvZf5XicOOnn8YTPT3aXueXSXDmfTllt2GFZzhGwhAmDgvL4jkVhYOAb8xjnLjMt
2mU2P2YUVclBuX2erzWesD5QjVvy1Wn3C7aRuSBvB0rys5swE0p0bgEJt766MeYUajbUSIvMEJwL
6lfSUbnqd9u1HwHrYJaTWlk5fkbcPTPRbGAmk2aX4pWWqTZhlYyfZUQZidmdVZm5mlFi4hQ2MtST
nfdiScrA7Q//i9mNdp6m8S4hrMimtRWxD2d0DxMrWOZ9Oh6nusNZZuSrT5vtyPN3Q94kqaqLJDDI
x8w3fT/w9A8lHR94UNZtyrhDeS1JA/xnXh5/vAYFL3RCktrI1KsN3Hj9vP+PTO6ETRj0+xWn5RMv
SkGb0tbRZ9FCw9vMnbY3ZRIAdVbpAJehFTNT2eyWItt4cdwgATlc/KfZ7TAJvcdSEnJ3WVLts5lM
eAskdbHIq2Dr2lW14TbMXyhpFNtgg7BiS9Bf/aPibmTBTrkjCv+g2ivWLoeoRiaclzcIwaJZG22j
K1VtssEvRVUe0w/jBX/dPkdshfPQiEFQl0vpRVZVPdFYIYzT6+1bVpVeCp+P4QiwYhhvyiV95YHn
hlfZ2a8cHYSKiXYmlOLmQhPKjfzc9SIJq3NNVDIQU/81oD6Q1c82eY0O6rrkXoDxoXRIMtzUpiFi
7089sNadkCpl6LZgnAy3ftHal1M5W3ZiEzYTIqLFeMNsmCL3AkVdFQUeuaX6Fz6l9cToPCszCuCy
HjzxAmY42qC2FxjeFZceN0ZvcAH7vk6ErSnM/R8vWNmWfVAG/96U8XH5kLGHvIoxasjGEXQyE86y
aeALxe/yTyhO9mAwDikxEbTHDjI6MhA3j9gJUeTHJcgdYv2fsmfRGsUOO+vJMSBze/o53oet2+yn
DAwZAZQPYOWjDTJMwr4Rta0WZBDSp2Kl2/qLMdwoDAhEr231lPLWeqlbIRLuXWkzmvFu/Eq/SzJt
jmQO8Fi4dXjSbrmxcH/glP57EG54r32KKUiCwdphIJGkkNO2iS0maHhqgCryYlSU7LJxGcPRoZPi
YpaTF3ajVRJn7kn/p95QkTDF30KYmcyDKhk+mbknvpfpewJoppSrExr06YFxuaS2xr7NVZ7iVF1j
lGn4GJX1428JNsqR1NELO+4MFu0ey6LGysRNoh+8T3spE9/MnTZoH8VAClMIZ5CZerRJDz995yOH
vy9I1mc07UuZmAzJdT8qxfgUDB8RG8nLVsnykD2iSX9v5uf7el9x7JEZHLENFt2ZMdU/XEB/a8Ia
15emjK6oI4qWY6Z7O2P+lD9AR1aM7UsO00z8mp88S2T/qDo9r/L8La4e8j/PtJRMwdqzzvLRiqBG
ebrxOxgTct+NSKh8MjOMz0XoPheyaK5vsDV8gH7l+VvrQZJAV8PESUXT52zw3Xmv+4R6IUDGh2RP
XuNZEVIOdJpBo38usv/+YyMgn3IQdJ7aiMhzheWeuphwh/NbXkNWrTjyCVDakVpofLm3FcAxYzOb
a55Z6ZAj6XQlon5y2IcL6vWqgxoI6ADbCfrYjJEpIaCnWy+KzN0BsqA3HPaandDxML0XA1ppd8/B
1z3D5LJe+vP6E3/X6mfgVDDBUtbK6rNBR0xb++nWd8RZWofbO7cyApaTMrFvFhXPEdQZPdQto32+
YSFpIWrZdI5XkerNPNz2EMwb8+9yog98K1CF2IY5X1+463euejFqR/Q5S6K7n89drl1ZFYimypdD
myV/r/xe0iwka3WfhULJ7Pjlcidkr9Idh7+Dx8RJHFPQgGUoBZonNlY4DJB/Ww9LsrCxpRwpqNbu
6lGKgLw9HpZysPcxRPl4DK9Wj4iK/q6fNnJR8Wh8d6lGJuZzuCcqXRSfaDc0Q3fRI6HoBI2kuCb+
1KhswxdGxZmYU3wcl7coLl2HYR194I1OxR3ry0k3C//DXcjPjsfQAcAh+3WU9cCkGUsadZ2N27ci
VPsy/yPKstRYhYDkID954nUPDbQjmn4HVTKrRVzX6ZRnR2zZrgOsLPBdXtOniPYc2W+HWwpx4fNl
RJX9brjG00BdzEEaCXklWYuxoEIh6uNwKSJwx5TxhMVKh4vuN9iXENc2hdePYGAuFKmgUdXiEmSI
2LZlEGrMkqRR9VT/Pfqw8oD64brUQ0KCvvPauCv9xnh6kZlGysBqqj0FunpkoIDe3LWiByp1GaS8
VB4F4PZGJQuFQXdoldYSxg9oYL3fZdZsIBRxOPEk5sSTIchXz1lMhGdMrjxujQx9qXR3mOYb3fec
WVQKi7x3bYk2s2t4ambk+WyiZO0SeaNBesTdzTFKdI0gKMOt4E1ccBHvfzidGCoNcdWFBysICwFw
mV0FsJiLbTcpO6U8ZrnKaElvSxt5tw/wYzi6ITIC0SVrBATdFJ/kk+cSjOOV/xMPRBy2eSLmAloS
QUaIn726y4Ok8WTmRzTVwh8mm6F2asaYQeqs9ygFCSwUGDUw4RJAm/DdUL6k6MZkB32jEofVqZmQ
gtnyWBzf0/GGRc8p3WGObg9l//OAPEQMfGXVKa1j8mNq0cBohKVGeReyb2jarl34X+sQnDb5e9NG
dLQT4h+zmi94n9bAErimjl6LNcjhv9Y4KDyTKL1Ue/glcs0EIETlANwORytNk+j6hRLMBrkBf9rQ
lNq7IRAm63jzsZgtYxO+wOunTXaptJDfrt2du2FFX+7/6/4SX7OYdwXku8ioLXtQ0F+IFlkDLnE/
81YUkW9/zKWzN1LymU0etvoEZ/uaz2SBj4cUDHfMVaXjPw3s7JdUDeB4VelkQvNMweHEyBTRM85T
764/GIPqTB4QSvTaLlGFjwVYWBHUNdRKowuwx6aY7x+/R80EwisBvM0kvyFXPO3wIOKV+lLB0qHs
bZBKJYPk6OaQXU5KyS1h9qPh/a89UoAApevpAaKhxGPSKI7vk1F5fHTWl4rGVVB75jjJh+rd4KsW
+qRN1Tr8W0o5yVraH+ZwUeYc8oltvqtSMsh+2vPJzHPueHYGsivMdM/mgxoXfIoc1SaoukmNnhIE
areoXR/SYdvN/6B3CT7sVlIZVQi2t1FCrzMUCoNpnzQTIp9IPiKBVYARNJdAChVpJ1MAtin6UX5c
FdSAhTqj0sBHHp+w68nXaA4+qOQwFmkjjNSOWw0qYabZPvQVH5JVJa1QTUYNsaMZ1Xnw1bv7ng/o
tb+iYADKSOnABgIo2rpZPPfXnokS26LosPs+TnPLxz5YnLDyp7v5IAdNUPEMEmf5VIMIdFR/U0lp
+hzh6ApUGL2StqJkLaGTiNtofwFppPTQcWyvZf4zXbMgqZz40MA7ushTK7wAGAJAjcWyo1ZmQ6uX
9n0xIN++y4XshDfjdyxdYBcXWs9rn8Hi9y8xI+oP3nddjVD4Qd67kLnw3jPCV+f5UENWG2OycnlJ
x70ORKyyvGQ6kVJRf3QKIBgSI8yQahzPEPn1CNW+8kDJd+wQ2GhQYYmcwPpPapC02yBmOT1BZkKs
ErDrwunyp0r/0vvbsga2YaQ2HBLU22M1OQhLdpoAcLVZ9Ijt5IcL7PNgzZHk4z3/+hyPnmUM1FMN
LvM3OMAEAhmpcmARdRYHcF29Mf+cnj3+i8KZEADCCM50pCIgWVPQ8tf2MDiPXOhFedHsg7rGliVE
cuL19j9Baqjx/+j6v7r79KYekY3zXyKYjuj+OXm2GqJhr7bCTNibYps3o247fYvipwq10bq133t6
GIvN/rtj39xGwuiD9P6X016RwOAngURZNubGZFLH3b6+HOKUg9nCi7c2y8IZDjeoiH1o5R2WkfWN
NTyADYFtISoVxp1ANECqiqsat1UoUrPuF77dHDpst4fGdyNW/G9L9cjQHd6JVeaKqMp2dgpa2VKn
/qDrSnhPzribYBI9uoml+xEiyJZk0SQyUAnUI5ETvW//MssdF5L4cDsKqFgzg8rYPNXW5bJucxEs
KxTT2LkGcJAPGZdCyEObgTxr8nK83PXNRGRllF3J8ohrcNGbByZlTfDD7Y8g7XzgSCdJ9ao14a2g
lBx/EiCwqMx8IasuZs8X8rGx+rLXub33rL328k/NQ+nmRmffO5Iqf+UDxAQ1OFMzQi5O10YrgXdG
gZLOITSb5hYLCivza/yAyvCuN77SbdhMmo9QXk/3uFZk4eZGlHYUqBUw3ta27iBDkM1UGbPeYYXJ
954m1iLrloh1eCPm0hxlU/47Bw+I/JAK0oHb6N9KDlLCj7uSO+5Kg9DGRs6iCztbvkz1FhNS/fUg
FH1oH5hGjrJhkUkR7eIv5bwogjcPp1BKGRfn2GZyPIWmIxU+WMZcpKB7NO09tJij3ATq7uX8VfPl
YCjYTcsEfLVRaE71NWpDN+pB2VkzlkNWuuAtqOBx9rBmt1Rv6rVZ5sRsM0kw5tL79VtD/VZ3Kt9z
keSQR34m0bYOBB48J47VzKmAiDS+Syk99BNhZyjYzKQ3fI4LO0QDEVMHIsdofwVGaJ9HHzYmZ0Q7
Qn8Ua5iBfbLCdadq/srot33NTkjFTmAbCeEAr7WMukGs9M302BjyWQ3hMBfR8fxm8BifdPvUPSVQ
6iCJ9pj+QaovioqW4JvZD5wIIep092yPw5Gz1CjeJBlElJV0pMkFSJEYaBvor0FlwpbnCJJjrtYi
VJNh2s8LwNWjQ9XnRsxJx4FfPs+jCFGpMMqdmk3yRQZkrxekE2zNPEoP2kgl+I1c9/ixhe2hxNQI
T/io4UG+iQglWllpaa/uDjF7LDYbAXs6sOnhuFZHuCV4S36OGeWRYwfBdIfV1MLnZ40yUe77V37g
OgCKczQGHs8Ygwi9umnFqwB1I3xkCe34d7k5lFJbP0lmcMVJXnd1/wLidnHN8rAK9DR+skJe8Rdm
UdpwoRO2kzLspp+rYAsvJnmSWalZX5taaDCMhcrsUbCJeGRMhAA+ySBtzT9wVkVv9MPc13EXjdtA
9rwqD/eFGn2+niCry/OvKvXpcxbAV+9XFi18JUlFsoojQG+ZPp9k1XfaQUr9UyXyd0Q2mZS/xMy4
MkU+My4uOiai1C4FgYTb3LxBfNcqrAHWH7bwqzyXOtwd0MXTa1I9UEW7JlyeYXHPFQF9JWzu91Y+
xFJoJgyBU6SwrJNVYBdeF5obzZtlNfFns0FBq1MxCl/8ppmsfPLUfbyYPO+B66zwID6+um3Ah/Mb
+1SoyH3MJr8cNLKLRw+kD7mqGdUf6dyuGqD0N5XFRpxV3eimiYwYFsHIApQCEyKlWvZLPAJPT8gE
8z9bKLIxc2ioK1Pk4zTiT5+BxS5DorBJ1OvBmkYYvC/CdM2pXC0qkdeF2nTk4dFs96xNkuV8OUQc
4uwSNKc7LmDMzVCp4AdHlrZ8Uwv8Xx2q1Iee61GLqswoxhhRzSUN2XmPXnVscFSmqCY/JbDwMIuj
PkqR28JDD0ONbecjHj+bl9wnjA3YYK6ZPaXD1cD3Yeg3BSaVVnP7sukR4wDcXOqIa3BrypFwJoiU
wdieAEOVgZr+5LEc4AoDtwyEaxgCn6ABqgz6ONxo5QNQpfUgPYR8KpsqMQydr9v7AuK0nxksXOTO
jIHz96W3MeloBqkKPuJdfu95zGJRI4d4BzueYYPkfrhQQ968elHrGVdF1JcLVhO/OxDY0UX+E/Pv
9KdN7NdVLMnAH4+eRnfR6Yxu0xByW4AbblNbIZAj7jmTTy5z9KmY7KzYSSrXjMK0nfAdiBWBwciL
5nMKe08a/KoYmInk6J6OVlcQNRfCvQ/VMXONQyu722BLLQ0HhSoUeZ4NDDtOA+XSiXBpLXD5LQyW
eGo5I3HqKTGmz57Tprvc1+ofci8EB93O++qojENy1WZ3KJuZVC5cBqEbo5TG9NbJXYYL96f8LUs2
Bq0v5+4Xj6fPrk6h09j3nNZ5Jsu422mP0ArJdXCJpZwvIJ4x/LhsMK1nxvCYZsxqB9XKzZKCajWw
9kIu93d17Aq8QMYqCI418lN7Zx2gPLGAf+6C/N3y/rPoez3d65LZ6Jbpref24toWQWaCESMDtiwx
2dGcT3KT9pYcvmUtehIZhmdN/DAyN3MhgM4h7urgGwaZa9MCiaVn+KW072vYLSyX4Ffi6t2pRF64
pon3y4YEq3gL4zbJNtyY2ICN+oryv44tchV7082gg03Ipgs/yymYR0sWZ1VezFn05xyIklAkQyKk
CtF29ngtFyulr4Xwkoy8hb1wz7Xoj3+USOnIGiaXCLFh6qX4elapMsLk7YOZEpxh06EdnovhHPd3
GyQmfvdcQT9uOBgqP5zfLh1ZEzLueKy9xzV/crYqXmtSVqBlFbbL0+Lx2MtvgzIlsMf+Z/X/+zgA
aPDMQuEppvKvd5f5Hp8ycUXfO3D2fhDKxupYC5Arm5kqZde3YQyCaswpqpLJejlN31x/f1XCViJD
iV6Gbrcd9ESWSXCSHo/i7RBpv7qGFsQP/ZS7QzELwmEU0lUQKXienJEx1gC8A5lhJaUoE4/1P/s4
n4DOBadSfYd1iDbpSyvwsTmXGMBzTlDSH45u/yOt8m/RD4Ww9iECDDFR68LBtBFB1Uov4h9XLPKW
vYUyL6jnPLYHQnu8WFCGQRvK95zKVeQLa7H9hylG9V6IJzOce+TOUGQ33uSNVOl6sPxpqJlZ7QIv
U8hRdLvf4UaTReR46w5k5ggr7DmRYJI7IOI4BUsheb7vgVMBtIj9iu+3FZTIWN2VDNqS0rFd+GXY
OYkzVDa52OkUKoe6e8i+ZawgGQPEAdZMmIjJhaX/6LrGJ7c6jDihjoBvXQrDZsYK54IoW0udPseZ
plI5ZtxZqwL6qCBa0+3Affahv9bMBbD3M2DqtxPiE/izXTx8SZPWY4cNYs9xnRMJAXqNs25Lgqu6
yxcC0htg7EDUgtZ0JfltE659OL2Fr+NVMnq42tMpHTmDFjJlHD/9qsluJkLohtlfS/Pjb0Zx9Bm7
aCvYxHg2J0cnvCa8GzDIAvSUge+X0cPl3FHyrEsPYsw7+1ogXEkNIUPwr6pTDBAhQWr6VJ9VB6Wq
8ec23164CuM0EZ2Mln0/0zE+wZZnzRLL5va0HwW7xOI8nkOI7W01Vd01INzPQbcVKJ2BmATQ5z1m
9qUT/4Vglm2MroEf2kPW+UffJaG00jMDkpOxIQT4p+Xr+FOyC1+/FtoCBxUTNLlWAd37TZ3776Yi
avV5hmsYXQfvOVAwD+Tx3VcOH5EN3nSbEQMEx9e6rN64wIZNtHupC271yUSOF7PpIIko9wgJvEQZ
E8xvM1Sme9fPdaS7l9+UEKBIMRaTsi+Qzxdo3yo6b7BHSCE1k2fzNxh3O9GM8btV9KX/qguE7/lP
BYRj50wfeTw2RUWx1nQ5xJL4hXTR9PbHD0OUeNk59ZvPoav+gtquh5RiwtSSNCaaBXT3taaGIHZA
bqIjXfo2Bjx9bLwG/u5kGu+3k9WRbhayVWd8c2HqsfsDVLll/4DDf2BGRR5/0JFWaa8ZRxcLw0mk
VJ8D2xfw77FurHYcGc0aGMdP0VugiocpEv+QNuyZdzm8EDnI3y6bUz0klEOwGJkbA84/im0GHqrr
p2PymXYPduChfmpgOhm5MNeOWqFFdjVzVLXTOBRhmfj11FGND0Mj8DqhyyN/mWWrhYgZe71KOG/X
h/zcyZrotBU6P3keslanJgWnCqwePJI0N7LJaK2HRrnRqoK54np2Pomq+wJE+l7qa/4xzyOspfQt
Bi1ErtOp0Y4K+RIxesOjhB6q8YN4SGwTJupQKf7EWJL3mKwkNMYaEFFA1IjeNTII1xjJs4BActZt
PAYdjJe0g3Wjfarx9g1bTjEYaWPQfbCeXGAUY0dyB65gtazNlYHPOYLDAa3o97vLjoSuQAEc4BxE
aMwx1Vt4xqcfcLcl2L1MFRO1cfxN6sNPh6lRH7Zv/hszzgWrgRC9EvOpldUcv2B3hkT5gqwxU2Ms
WtxWOo/JktGLFpeIIMwU8P8MxwyhXF2z5NQGx4ZLn9JueUjW8zARUCWlhxu/GXEtE9s3PT9L1quD
9uAWZuEIV+ZWcQg0o3Qj9ZsJVXRIENOZxw/LDNWeCJHRWjdgy1S2qjCbO7ch/rdKj8AnWkfRITEf
5WJ0iFJqPkTrYT68Ceh+btV8AgNRvZNRn40AnrSIAM4AZJCl0VZZA8PuhwQ63qiS2pKjMYDK0dBJ
tnGJO/eC4brnJlNxpnMWNdU4Acbpl+8O6e+PFdUH7Ws0fbjaGlcb5g6MdzvRRDbofqyHv/1z+kpk
OEl5Le/FNfL+Hi+Xtu0C2tWhPH3AHB5cQHleCtixXND9CnyER6LIHzGxDtz6Zf7lh8W4xogansUC
yJqDbGiBbFkNNNPkcdI62q96uJtI0jSXF/Tu4oRvv1D5SrAoOYP3Dg00mhEXx+rkZlZj1mwu4shp
tk5qqkl87vYmwEeJWONZ61HwLvGmYJ7tgGAmgBYLLrucQvrbhNVefyLu3boKsbSiEF07CcsD5EuB
yfPP61X/J5KDkt0Ckk2HG/ZncMlpFEn4LkCIkv3BAR0aSDaRqfuhl3TLhfniuXOktakWNcEvhpPZ
HKJV8BVSun3e8xfkm2q9Qa9AOmlthI1dykPr1LLMtFMdZsKW0HMPLslT2IPpkOn8b2dZH7Q4rcZL
vZk/BYqltdmRGWc12jb+MCrh6AOIy8+OKu6VbX3aGrCfKhCkX3W/zuwZhzk0SaQCC2bpGdmiz4lR
UT+3ScDRjeGZXGYEmSnVe1UcIBfYtlpv7RYVRZrF/cYlzQt675dtFqURUnQZHRurStKxzl9ilVe9
YX94tkuvcbxJvL8amc5ZPDf+Rqf3tx+QlbqG0pUZdOr7kmSBWY3ceme3TStqOKAd6nRJTRgPNz2Q
5e6Cuaz9J/qWCAGN8WTq6uDNeEaqmu0RqoTDWJRBddIgy+CLR0H3fGaDeKlKKvOAGRLPMe1oRNOS
y5f+cznFnHd6mI++/Gj6vXuNwibdSuLDDubSAkQtJNP6Wc6OhCu01TUvhGm3jwajtLoDG8zmL/ZJ
gc6tdFPQS3EzVrFrut0MZ/W2PwGzaSrkhpsZMn8fLEGxVJ0UB3s+kB9gY0Z2mxoxr1GbnX9a0naK
d7LtN2ot+COPaL7/u7nYdm5/Cd/MBkUwWD2rzJqFShMN/xkMQFzP/e7qoiaZ5GOsmmk7iehGpxkp
5Nyi2+UfTZtE2The8iyObsK/sIt6AQNIUQjitFH91DtKfX3oQ6sDzOQq2YKXgV3p7vbz3WkKVMU1
5wXdqhP4PUmz8iQckfQWg3MaNHaOZXR4Vkyj8GErsL/BdpNvwxSWpTlfFUZSJ8Jl0kUxV1zcG71a
0m1RhCCEdmLtRwuk2bAWNG2xgBWsoy9AFyKSeZk1OBoYBIpfhC0HGj/07rAVhgb9RgZokZW1oEig
yijhL/Ma6j8lAwoQe6LCoEtYQfiZF+KZqYk4TmpbNCkli95zRnY3+hqHfoyaF+OsJuTTsIQynhmE
eQSBHiIlvxyIBPP3dejBlubF5tpM/ri7SESdFedcTELG7ZxiMBlIuecRPfNJqanxjjdV6XgWfYto
+jebzWpa9ZimwN2G5b09NdzT7eJmy7OeDY0xT9Ts7XYcftzCbI9DWB8HosOAnfaSe4Ps9vlzBGBy
pI9GOPTiE+P/OYH++PZ5X2oPhd9nCPAnGBlaxS4tryyKvxnIV6ls9iAF2ZN7JrqktUJYaKeuBY8X
i3nGHF59oJsA4jQxltlUTaCxuY2qBMeBUgk8Nc+JWHxapbXvMGcXo6E4YxW+macJvSxjrBkKFmuO
LVj6Rq/tA/oDT81sTe2fh501S8qbshc4pOT/fygcqZFqzhzwL1hIqPxiUAWT9OzWti4fjqeWfurY
FSA0g0yMsT8/R0Mu6G6Ya34XPDPedCTXJ4BK5qvLiqKyrwCWgVz63nrTS98QsD7i0rFm6n21FtQl
ebytNt4Z5YGKvcjZsazlLB4491jlLMjb4ZiEJHz9lZ40zMUUpmgTEk/5IAxzEDNC6PeF4hOXPNLE
bvLu9azOBGERSTvS9+kkLyLAB1EX+Esjc1vtiA6tfLFwOw5DSsnvK+YCUmcf2pHHBJrxSEQ2Ipsj
99ENeG37QRi576dA2rKn5YWGnVrprz9B/DjEZV95reJuyL3DrFTX5wYG+s2LPei8I4vAFsqkdIWX
GSM1vHZ/gfsm4hFAohzI/6LyIL7japuHtKvhknKt0oI3QPlS7FkVfg8W1GAP8PfuOC+NeCiBaLaz
rLXEycBT/Hn6blIwprEThGRWcmK/s4XGxzJuY9RIaKkM3umQKiABu0UPPFz7fSN+387U7f19ag+x
ZSjnHwBSbEunKezfQe/4QFfTR4U4jcFs96ZOw/GpwCSy2RryadAl06TM72fkg/2wwn5x0CdORcW5
CQNb4MReEDbZwt4ULaxC6ejKvBpo72hovqamNwbRBYzWIXAphP29MQ92118zSxaOFr/RgkInutvZ
JIeiTCLl8WXVE6mKc/OYp3OpNmbWuHM0/Q6GG6q80RfOx6gj/9gvNFlX1a+81+F31EV090iybRIU
0eIqLfsFXef66x81ksGPy/gjPWwTSWj2WNQ+4n6iWewxK3y0UTRH06ouo+yyjLH+gUV521mQkwTh
xCQ12WG8hGFsLUOPL5DPvNhLANPthy9KposScpezx0IWC4oyiY110P1GTJk2Mt0IYXJauKkHS3vp
1o3Du2wdfYDHYzFLbwMcnDzwPsKFj4Dne1l1I62He/qiPpSd43PnZA+qAKVnfq92ibd3WnM/miK0
RTx38TcbbEvxqui92tnUHE78w45j4BFOOzaTgeIwK5PLBvl8SB467UtzCxULMydsEUayFmwewbdO
5NkLl8yCpHXGO+iUi2lyAaMMrL++4CkYqhZZgSNUVZQUVXocuQgd2pWqivqMhJqtaLg2YlXf3yZ/
YGgtjvilZ/zpWoGdYlpPShrjf2oCUZQTaItfJbIQHsx5TjQeDO9ZOYsdyvKciO6Rpw98LwUZML4j
FgJshevpF6plvDuDcEKsZ192+pguT0om3/MPbrT1raUaV8OyLFB89WQw1Pm5DyoScSzo1yZx8pQ6
+0qV91qLLxkbVjFu9bjvTEeMHVAkPx+JgxmSmfDDnNYMOZpNQtEYCfBUNcd6NbAvb5PISp37MagH
1PJIvhl88bsuc86ZveURLYGHjVKRHnypfRL3Zake6UFhAS7VnB/icp3S84JTGsyilVozcWCSDzBK
QstdVzuYI3Co3kalVTSDAQWsh4Vcq5y79/mxCvFAKJpGyNuWjf2d+Jlyt5Y6BRuXUA3tngTIPtiP
UX5Ww5Iz9Wk/kZgYESzLphfYPtKWYQA+K1+ApWS1vkBbz3dMpSTzYzW0EkUpJHS5QGr625CfEGyt
1CgdfWLlRF/eRpaqyM1Nz7A9HacOnMbdb1XHANmuLTspC4ST5HEZsAvNwGiEyWl2zYq4HV3FisFP
B0GlwocSN4lCGMADpHHKoW4WWazDKq17nPZJH/oVpU/LRfRXV1zkoldbZh5ozZtUIZGSuBevL3p7
dTOo94P1Kzwk6wYJEAorMHzIQ5J5w4QzekAE6FZAXzPKFLuSPV82eVDy1BQgb3ahTKVn/FerprRw
gDvJfRGYAnfXbzxh+waWLtjtpmuElX00iu5pRaoC6D5bUFi2P0CeieeviBpOO+Q3Sz7rXQk9QsKA
4GtB8fgHmdg54J4gDuUeHlqMYNwO+lmb0smPCJsidgYb/mTDrVqEV/Zl1UEs+2lmUhuG+YOD6Mrh
erBsVMZMhCHMWOEJrejjt6l/6biYevBis2BV8EXV/zrKyVgEDr0Sv7UEGGwzk5cVYetCSjnEaymw
FVZCc/ZaqITWoUmyEcGVNNqKiAUt4Iu9gYxM2rrk2rEurLvfJn9NU6ru130Wji2Z8fadOzIOyZu3
cUpCaq6TZdtOU08rIpn1kbAtMlDG7MWVIR1v1I9haBzKpK76/CFYB8Z0Pm+wtHp0mrWNiB6hke3m
Anf+e+MimvNtV9yr62KQxxcndxN5Md4thFSJE8+TOEp098LQAUfLAvgYZdHKdN0rhyja8CsGDn82
JZTH/pYaWDzn6RE/UUvcBCE5oyoy1zB8lRHTI8SOeN4rZdttfeT2ddVLPIHrknmRHnbKCaep56SY
EUPmjPbYyZMKnjC5Hjlo+SVt0Shdw1yI8FWx8TompWvaa02DYtRw65YI31/rQPYzJ8kSwUHeMODV
bDCQLo1wImTbYm2PkJPt6y7eqhM6P//p0Y0hBmOfpb1hMxK3U3wRdchwu19qGek76hAqV3Nd1P4J
+uF8nqYeXNNNDVyak/asePUNu9tGA0+SHHUavqCe3OcHilk3/24lW1Sogk66Q0WuerVqpagJT3pz
iQgIgqX7nXYBt3gyVbiOF5nwkxoSBqsQ3uS9dFw3+uoWzNPn7ejYZunqihRHvSQsGln9/NubD8eT
P6oeVX9zoaX3nR8SKQqVYWfMOD3Dp6y442chYxvOAjkv2VRVjQRG9WuWlUMQz4uRs67ImX0HNbqi
9/Eg3AeObJ8QLlUOzC6kTA3wi7KFEPsgW/EGxewmwBFx39T0AFEkZsjDbTeS+Zab4yUT8W+QetiG
hbOiWzjOnrFM5hr1/7F/5URZUHlfDp+BKTCQ3emyvwEkKpAO/hVZiRV4nmFG2VP/t334JSGowg1e
YsI5OUNKygbXYfNQUG1Jz4huHXdyyWGrIWGI6j2gvgHKGkdR33M3yRqIyXKdWd7HUaJ/6lKZkC6K
gjiaALaGX3XIbWw55fuOXXgDq4GQH7OuJyCmoG8NV/IHrszgUH87sKZ84Qb2P7b9I9XV05iwD6Vg
v71jvuf5BdxCSAalCF6lDB6VZhl92l20vIYVlmVdGSoXQzS7t95FipKci1XaZ7XxQX/JGwe7pYMc
rrm0ypSkdLqs2brF6Q02dImYUg8xr5X4q6JVpubgsdbezfUVDeftb61CZa4jd9LVU8YvYXSJLb3t
Et0MUuhJ+X5O+JD3ZM2hgnCDDj/2FPdpVqyRWssKcLTQzndw7X/8g+FkRPRKro+dgdlo7RwACgfr
TPDIoO0WdtRyuavSg6mnave/mnOwzq7sbagAyzBm7shBXagouwBtK+Rxlje+iNyzVccIMrxl+W31
Hj78ezFxIwsTP468U8E9uwjWIm6/SmM3mU/aDOKnLUU7OtIfUJU66nluEujFVkTroq5RSr4DNoMZ
MaWX1Ns61xPMA8HltaHcMlG+S1x512pzPB3HFSyq0+eju3OUheknZpjYVoXXiof+lzPJWxh93o/+
q1rcFbHi44mAaY7mxSpywi8cz8Jpve7AoIDswnGrBit3YNvzLxdKEgc+0+IawJyV1+sjg1HiGFQW
eTGr/qhfm6rgV0/CIQxgGYQKs4ITQjFnD6OxQDhaXt0zDKrG9V6DriKVF3x7dYIZIxR8ZTnVus2q
pptQdEO9hxhN2hgplCQkq3cc/YNn/upGzQhSn9kFGXW4wgcExvTgCaK8SccpVtvv70uVfnDykebB
eToyfZINqpHtFx99jsF38ptci+a5TesexrjVvCeP+HwPA4wvVTbG2A6sJsg99teK75TwdAGQQf+q
2VJ1d44ma5+G6cFlQAzwv5P3WQC1THWsbxiFT8ZpJeo+zCGD9mEwU0FgzVrvcR+LPLJKXq2etBY+
M4DSrlCBl8sa3kXwlRjm3lmUiEeiCyLLUNv27ePnKdXpyHzzQp5IgRGeFfJEYB/xatNZn//S1p9l
gkm0XmNN+H8YG+464NrmZYQHj4Pr34CGPzSIlHsFUGs3rUaKV0trALRqW5kEjCcANi9YeIZQaEeT
JOBZnrrgF2qSkcbpKlg7DWXByNtXz+WUXerh1iuLMhkB0eUtf00LEMEDkhKA5OIzeB0uiDmsx7zN
yLKSjXeo4f8qVp47jV6kJNk7RP2T/BpLyYGZE/NTFLa2P+aUgcQFPCIcBuNvwdWbjAduGgYO/i+h
xi3qRtnPN7Do/FFgmeCB/JMq7872piSj5lCg1KLIcu3K82jwkljX4YaN9qOrrixwrHKrxR9ZYnXu
0vP4bYugYGHOs0+HFNYlb9E+Cu17uABnrMg7x5yaQMIykWn3cFu3hEdycsosr37rlmc81IGX8Moy
87vP8eowKCqrGNchRugRuwc4hv/UwaFkaafWtuNjbT0FxZv0isFKNhvt2JRPIyahr3Zt1Q83KunX
0D0M31ZCAn9p7JJ2cTg0Wz79JeaKlBlA09KjlPIgeSAy4zcKKhVOwyrluWmr5MHAhzfGYaDjvK3S
YNulU8/rKjIyB8RMv7oiNFaeUeR4gbHBtMLDc0xzbjtK1A0/cDyELKrEhb6uavyNeZz54Uusupez
s83fD299FXsE81KT7HuiAa9/SyZwGbCxSRxOMiM68Cn2Y5wnRGQAMHPM6ZHud4Pp48Z1voJ7TqXJ
YwzBVGce80y36i/J/xxNCb0fX4G3Uh3bec5EMWfdxlQ7bwwgtv/TLoUyA2OQa2owi1KhECjn6r6t
CC+Z423HbUZB/WiFWzlyK1rwn+ZZVVAf89Ja8ELvXrn/2otQGOBpDyHeSoVEBxTZrRUJE/ZFL+9s
Gzq5XI3saqjOFYaSyZBnMx/hZc0xRUF3wAT0PvrH214wVFVQYW7DPAW44RgHVmmX+qp96nRYvItJ
0HUDG5Tdo28GIF1CznUGqp/nkIcTOFJ6YDg4jU6vZP+zuwux2OPJ3pdQUYI4rGqmTsuDv0PV9R+3
LM3+2LSGttKCzzy+jjovQ0IbMCpbrSDiaIIIE7ato2AOjSTuZfv4fdJJoSR1O6GChOCn6i73Ifjx
8ErolxUm77eNXtRbpGWpMrwg47GBAjmC+3f8rbuJIvkdY5pAWo/xbzsP4Og3mu9zCevATBvug8Su
BaI7xScPViG/ubj68ljN7ObmFUuICH2+vWiBlop2qC+Pmknmm/lTF5UdrE3mqZAkBPiYKigCuYVL
cjG4bZymNN/2W8iYP8I/Oy0NyL54hIY7im/o2+l9RMY0I2JucLxb+K+RayGAmDuT+lVkPZTmqxKA
KhfNiPfm4zw/QlYokkNMF4YnxN2YUFCgnh6Hwp0GsPdjUGN8UvbwkIOa8xRyXnxGtkWkLwD2UtV2
CFR3ZRX1oNuuqG00Q9annnxpDM6lqDnM4z7p0RAAqQsHU3KxrJzwtVWPzIpSmrTfOCbzX5Qq38m5
gKqiNDKeQnuUzJGKk/7zZnfIysgBoLk09N+auq3RaIsyJkDivm11bugG1SOlnHMe56WJzi7KPPUe
evnePKAl4acT4TyTwJsQYLiukedN79oT9H9w4kTAHTl+ZilnqGZY9ZcIuoAKaq44Ps4rIeu2sQJg
Tsr3lccuIFu+pHeIbdclMAvnkYkxQMYEj3KMtmTuNfQMUMxA0Zmpu7c3thwxKlOEZVmyt8favIpW
AbfSTbSLzsxRvKmKDeAYSCboaCnw1FN6e9vdpRj22o0=

`pragma protect end_protected

