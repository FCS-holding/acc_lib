��/  ��Q(���]G%�B�C��G�1�*�$�^�Z��%�������[�Wq�~`�	v�.@s�Yꥱ��+[q�~�����h\x�W�f��O�盁G{b�]���i {����~.q}<�	���`�� �)���(�c�,��e�ط�5��]5q=ee4�͛�I�*��-�ѷ���z"cu�{D��x&г���?� 7E�R�]��B�K�CJ[�4?H]�̈́9�ۋ_Ͳ*ž7�iڹ�����%>H�
�燔�rH7�u@y��;
�oj��$ѷn�� Y0%�E��0>	�u=\uh9h�2�M�$/�8�\j&��R$�O0�|��3����I+�Qp�O�W�;im\��^��dքq��lI(^���a#O@��
]���#����c�y2������m�?�����;,o��B����P|�)Q��+H{�j��ǭ��0��1��'���8�Xu'E'̻������!X�M��(��3z��Ac�`/4('z��I�A�G@��q�-��K���_Gh�}}�T�F����4E+�9�iPd�u�;��6����Cgq��>`�r��A�t�|YJ����A8�71	�46[�N���3���D���f]}6�� $���㚙|m�� �#*D��`�1�6���W~���c�A_�ƨ�p�]��m(�l� �b��w�စ)�E7	ߑ���Թ��l���!�XL����|�N�Jg�;/�G5���؄�k�F3�):��ר��7ҡ�m������
��<�8�s7��Q��:+�y���~�� �jG�8㘮a��'�q�GQ\lȥE��m��KW&�R$~��R����$3�@cfL%��'򗽺�u�G�Um�t#����`�۵���]-��N�>\�3F��ǧ��K��	���&��/I���ՇT7����Y��U	���sr�'J��hW9��y�TX륂`@
Y]iT�R��ϴo��I��XmM�p^���Y�Mݳ.�0�Է;��"m��*;��l�|I� �˼g��ͿI
U���1��M�?vq�w�4Q2���ǲ��1���4o҄DW��[����=�g ����N�%���H�&�(j�%��^陀�IRj���	���M�*���+��������𗌸�V1u�G _�Ĕ�i�x��-��}`~@����\`Ӊ�3�����Lx�&�{����/��
y> �� �<f86�#*�c��բI
�ZU�_?hrfs�8����q	t�r@���%#3�bذ��崸��5D�̡�0y�l[��+���#;iG��_�t
̎Z�c�	��t�z�	���d�SE�1�s���l��v�i�<V0s��9$^ƴ��m��-o� �9&N�  Ή���crOJ�N���p<�W~���X@9�KB4ǹ)>Yi�T�]�B��}:�tb���b�Q#5��W���� �Ry���gK�$ �3쏲� 9"��|��	��Z�o�Q�x�����/8ts)kJ5��>��U�<Ή.P(���&A����&�M�1��)����%#�"ct��[R�����\��Eн�D�#%��<W���05���,��