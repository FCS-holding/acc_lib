------------------------------------------------------------------------
----
---- This file has been generated the 2020/03/16 - 11:19:27.
---- This file can be used with xilinx tools.
---- This file is intended to target xilinx FPGAs.
---- DRM HDK VERSION 4.1.0.0.
---- DRM VERSION 4.1.0.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinx_2016_05", key_method="rsa"
`protect key_block
CZooit/JMbwjeAcsO93z0bIRcr24D1fUn6/8hCyIijFRYc2bYgdf5bk43HvJVFCQ9f7PE1N4Snzz
e4KvlHA4VDVFxrsDm8pNeX1eVZ6mfPgbz8pv3Sr+7//oTYBg5VUylAm9j6DnXn/be/QEEEJV25pE
JQdQYhhPCoNgcJHlRylhVIzLLXx5G81DOl3N8AGeYzDFX2HLb/qOCbh2rVclfWF2BceWD3e2QRpz
KI357bqs8Uk2FZKX3LLENgMpb2grJKU22TNpT7HMl9HScdnnUps2l2cZDQuTxzzaKb8KYrDShjQA
ez2tUL3XtJiUaMLgLF+g/2KFWiYpvtgqEqqHeQ==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
ImmRyy+o/AQ8dWvdAgbC3cYogRL08EEgNDYXVPoBiFj2NLHy5oUTr10Ph1NgMeyJGyL/aA24ewOA
rxR8awghd9BiyeNEEFfKl79shEcFPBTdJBsuEBjxI9RwodP4OPdc9hIu73RKcY/UVpKRVbjRAbLh
NA26U7En/3k1JtB2Myh2BjaJYpHJqUiC6Cbfmo1XKerjRMl0cx21nHvh1Ja8sa8gV+h9hiFeC1MR
U9p547+wErindjxTvTRJHioBaVX7Je1dBmwA4ip4utSjDdY5GmYRzFVdBS5weA9yt2vM4owgfbjr
GKfsMlRwjgEPn8l67JPGyhIxP3Y68gjf57D+NQ==

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2019_02", key_method="rsa"
`protect key_block
l7wdPjKyXY88S1SHQQfbncFmBMcUZ0zZWjJivgBZSbAxND5U8CM5xsHJOKkU1Bgr3phCPtTDPle9
1UZWqdv67wFICKvnIPP1lE5JFiy4KzFCSp8RjcX9QudW8MGMMbXe+uhnsCuhytErrcCAs92mOtv2
Xiu+yPxnY95eu6Qn5hohzUJYTJi3rRCwfFgIBE9dXDOOyQLBWsMcN6PecrnD2A3GWR0EL2De03v1
RlEHOJgV2onUJh04p2nJhxbflsnJparQnKjfo+XZNzJs5QgBq3GzhCCs0HPOr5DMAWwaiwPhibnM
n2VZYoRT5Fbxq8arrUQDxOH7z/jmx+ciwHEGHQ==

`protect encoding=(enctype="base64", line_length=76, bytes=835872)
`protect data_method="aes128-cbc"
`protect data_block
KV9Kl20INYNPrE/NJCox1DajRwydpIgEUcZqEXHGE5bncwrucNiGfskuqys/6kBIWSapw6nSToV0
ZtXC+9dka/+788b4VqaddSMW7uCnbgYAQbtQM450igNwZ6jAtx5yOJKGp0bACzYn226wRM8vsobw
ZTOMjFOMsRvQzCMA7Z0uwdrbY9gSETzGihEdvQvrC9uED6V/a189bAs8MLQ98XJtKW5vTuhFsGGY
aiywSa/f+I7k6TpIgCv6oWLAkA/ev7hxlFmag59LGiPnx+Mh7FWIhLUxwfLOH5lL2XSBTE6vfvuh
/ovYS9owR7Thw4UthnkBoCd2ZAX/1IRIA5Uzmb98JRiZxskHMCekTcueGBFwJYKStBw7GPkxnolp
GtqYerZEQb8cj1PQ0j0PhuPxXecxZk2B7+xEO9RVgyeZgV/tKlbC5sWU4WoMa7Qzx1PyFMaFq4zi
jI+toQ6ZWTGF37/Wjk2Uvi4RMvIuwPsMb0evlq7FbaCYUeTWyKoaiV+Ae6Wua8na9OqeoRQl+eeL
g4zPuGJT8ZBuIQevpUDN+mSxXON2O0ZT98+wJAlJoEZi6goArU5n+h7qptQ+JJZHQW7g2O9xTVd0
nVLG8JAghH6u6KWqd7fNzSxY8QOTMO+/levxD9y2zrjcSwJLtZ902c0ya7voWUliA+nIkd82SedU
YKaoHRR4WiZ841fFDWNW/QYbI41IcO4P9Gy280rJnm/1aSm3JDDPecJfqHmzx1Bke0KYwnO0kiFv
sEFYPRSysacKD5jp4LFRdTiMXB7YOug5hW6PfwuQgLMizgg0Ez21S+JHBb50fOdY6LkVw2jw5dlI
2TtLkXxxPXcX+PDNiVOevkH0Ub/mPp/xWovnPJ7JdRN49uDPg3bGL8BeiASHS1S0KUOWzCOMzxfZ
yMDFFDt+8nJvN1OOy3xqSRWbiTSEOXbT6uwkKbxgvN3fMvvZkVg7h9S/OE8l6Ak+HdDN1xjfxODr
6SZyUY99x/0LSUpeCmS+h12PEzs4WDBWyv2KgaeIf52AmSy5UUhz/47BIHYQdQSeSQOOVG4ypOat
3GS7v3ljcPt1DKU27n5kXlZM79IpoLPYuVaSq9ZBFskC6Wwx+m+9oUJ/R45AhTWexQyCJ4V2LFeN
+mvBbuqMrKHwC+o7r1p87r1i6BOvYNZsyhMSPwno2oN6lKtwtOxCMcl4MXxlMYPFEAAHw9ZgI1KS
+0DFNI5HnUS0W/rNleApnoayto3fQu1ji7ssYdkqRIl/3vqj20gmtcVFLzt1tHk8teh6i7muKOm+
N9RtkEIYdSYq5EXzDqjydLWf0GSS1BNoWmXPDLBsYUnZ+uoRA30tOJhFHPkgCn/8/mHLFnw2jE2f
6vhPXPbYBnx2R6J2wX9kjW1QQxmpBOeSZDhv8K4XAQsX7VhUVR1eJsZn25yLYC0ll9TYTD19FGyK
L1bQZFhO5jt1h0ziboUTysEZa4chKOkYsuMAKiL/NrFZOJ2BOTn5DbdvlIPJUN3som9qwqFOnmtl
qeHtlZ0eADk4j1zLTXqoQjnLscKxvXHc3968mfBnRzRlHmcvse/3Je7U4p9j3JjfzKrpDwozp7Du
alKSrJMapxmNL8KtmdkuYPGvJeHKwxFpxbA6eW131o24hDTPekLOlnAgUW4Yu12HLaJJTpqsntA7
Gs33Vw4Y+H8ySLKY523d8CPalJtzzn7v72GkEB9hLYeGNBnlziw/RlJFABsR9xNMADryKu9ATzm3
1ibpvPdq3vggAZzppRc/Am7ZO6poB7IpPaiPtlJRyzWhUwHxLBD4ZctVuvuQZI8nJZhv8Vr3dOta
9Jxu7hPatel7LW8Y5zokiK1Nf36NUFV5XvL8nK7fLLjMA2mUTOBMwiSWjRyQzHa/yrgmwE0CSkCT
yry/3X1rx2LxhIS4mDfEhySTbQwRHksdU15HZe4IUWXPHDAILRHU8oXQTcd3HO8UAXukaDvwk26c
N+zoIn7wsLGpsouAJq4TI7oxaJ3HicSYC1uhZEognyBRxS8V5Qo49KHI3LN8Qgk1kZUDPsyUS965
RLmuetFu5did53Weun9qQbbFSKUf6XXDigWbj4O/e7730Tw4leWsfxF5E/eXwxbeHRFfJuG4ORjt
KOkGoijMDM8VQvPHl9aH/3gFkxibS42xwplKLVBMBQGgMOfGaxkFbP7ALFaQvNK0Hy5J799nopTq
SNJpUCbxuJrEk5VaBqjgipa9uXv1XGsaBbgcoZn7yLXmlrqEf7+KzgGUrvTtCNRrbQHFkHsJnP6/
jiTcA3aF7iNwI+/t7K8833/Mv3ythcJDjF8rjL5z2DYl00GkTUEN6l3W6A4ElVw+/LgXs7DR121q
3RBp9FyONywDntiuNddkS+haE0Bu0smAzPCkmD5iJvUhIsrgt6FX20Koby5c2gBgK0ehkd66QdQT
TQJA3F5NKo7Y5DgGHTGa2mHSIsHVgDTzsptrzy9vOrYRKjv4kQMl+yUuP7g9cJJSf4wjhSn9CsNJ
tAOftGtD0ASjzJP9B1PQf3FGTZhn0FBseDLnrXUlMLgrbCx2q7aT8IKKRuSjufSHTdlaUR/g0HlN
oV0vbdUzourJGuJTSzgIXZ5tkYR3iQmpWp8B9JF5lBdz07SEpy/AXz+NTw31teoq2UEkedKcpLzb
17n67yImZsM0flEvrtF/7ebznX1N7dr140fN/1OKA5wnlIL6E8KdnmcCv3R8+wn05SS9h/PsfORK
hB+Dk83mFl5J4GYHiVG7Z2MILUlXpSmzZ4fHONOevtnEiQh1mhXy7wZOCg9+VaxfDdcOh2V9uwIh
ebDDIuDbQSxJncAXi0jKMfByzzUVE2MLOCrby6PNAm58fJ7It4747xiqnx3A7bfGX5s99CWjMC/p
jDeRcMSHwxlI7dX5aHC+QuWFBSCqVjCAjSOFkeiXMJiGwbjFOTLWQVC5DsWl0s/ZIOLJv3t7pcJN
B82utfYk4mNZY1WkUPCP1cO3onHYQRX1KHd2pqgZntZM8HYhik3RooMg0l8NPBGTIbxoZRlAAPbV
IQhsbq6iJ7qg40wltWakb52fGijPBDuHfJtvcJEe7+OcJ4tDE8AzlkVLnkUbW8pHecY3crqHJXIL
Nk9LRE5Crc/lvKLaKDa7HIJHWe/MBHnPmO4p/CyteAFs5DXgO8xBYY6PObfj4wDCmI33ZXZOplNz
DwFCFtkTDqODLX0YKYDK3wXb1FwZ41Fi+M9UX7U5I77FpucyTHFQORh1wND2Nfw8Tk/T5D9Bfk3W
U6eARwIYYNiL9B8j1FMzBZoHxWjZ2zfD23+JNn5Sl5ykHZaiDKMWHtT31WeYJqIljIAVwnWLp5Bf
GaGc+nGFTXbKCflMStQVZRCGAsCsAm0e53qfg8iUgo6+0sSxIWAEyMDtAw8ZTO+Rxnsvyz4qptKr
9gS0yg+n9PPR403yK91gqQxMOvmDrzRJzNBK85Kq2i1Zvd0VQCLpDU6JRqOAluMNjk188QjXx6h9
7Gv4Xin+W2sYgtDMtg0TLkc0oPlBpZjvNSl1Q0UHUWGquLed4Wgu8UnLw4aHv38wAv2Wh5YcGk+z
zZkiF2gCKX5kDGPyyt+3I0zuUU4k5EnjRZ1kJDI09575RW+5tTL3fTtdBY2UQFBx82wYy0CVwnR2
CdDWu0pBqh92eHErW9+bIrW4r8gtTpwa1pI3id6rxU05xUElfBq1bYtGqw+O8r1BIFuXbB9LI84K
V6NhaOu3zIHV6612L/iny04aVej0N9/XHBG8cPIW0OkxHZ3jjALCrQAIEgG3RtkIzAej0tll8vY3
B4GfvXEjcT9K8yDTNIVnbSqiSmnINnkk10WAIUZkNZSTDooMq9vd0qQchK32eP0ckn1UaHX2K1f9
WapH+DC5YuokJFbZhCs3AGCjgE0hMbepie/vfLgrpSgvZMOJiaAbRXYgjCrT2k12SAP42iUWXUxO
BJjkM0mHR7G7IgbNjIcePVsRR0KAw32uQq2F4+lYHXoC25AVzyJJDqsCZEXKHe7poNBQeu7Af+lO
c6hB0rCL2Llra8K0XjbCGt1x+uUiUt+suLBSot5W8LVCZwe2vQcIjnyyOvxwNnzQcOfSLqzf8Mhc
Eww07qtH/1yEtB5J5wDYEqwKbTU5zq2r6ZTs5pN4RiQztDCkcjBroY/3Eaa2t2JPKFzvuhaagJxA
UckDbMyuitI6wq2XsyU9Euqc0493GT7z3V5EVUNnWjgVL5ZcHfWTXVI1AAFEiTT91CWnX99PLKL3
Bwv2QqtnxDsK4F83omuF/1IRJ1h9Y1bhrkSyX67OzZcrB9OxWi6rXxSQgQZBJ0GbFHabs0S7oO5m
GyNctcwd5MDVJjwoXTjamRAVEVQFjh8JE1KHpHPqEYb+fvYSm3pcEJCuvWIDhIs71pm5NkEzcyMf
jZG65M0uswsUTpjV4CiiXQz4pdpMRL5F6rcllrF08SEWgjeQg+Dy/ovuPY4qQlBsnlS34nMkZbK8
1FPZYWsOCEjgVti6xpjzcDcJS/1PGzHMLPwy3FvjJwUSX6z4NX1G2K1Avza+c1AU8NSO2LNsHItG
LcS1w1OU2saYFG3aUW4+ojKJ1reUaT80TF2DLFo6KCnv0Z5GUEgYxvGnhyFaqgcN8W82M7JJPnCP
XuGylILzrZHgnlCGpBYIATJrBlEXUKRiK15JygVC+Kza5S1w1AKVv96rU54njha3muksWMtkoPtY
+QCO8zTBIijjK+ibyv9yFUl3k27ZLUceb6XPfvqNsW7GHeCAV1eJut9H+MwgkJmN9ku4hbEs8wfZ
QpDG57vbv9W45w2HVJdcurtBaNl2vVlKlJ9hAMaeDPk0R3x8H4cOtvjp4u36v/IHtTBVozqfRUtg
Csu3jv/HsgrTunJb++oOfefNWJESD/3tJiWpiFADNATgr2bcYXYg+YQsc8g/xKo3+6w4D+DoMJ0Z
oxPZeRfP6UyX9N7vRxZNZblUYDH/7C9peQM8AAV6gcN4LMs7zPUWTl+MZCgNzNPML06QyovMTzQd
kb60Js8hLFO5Z0eWHZz+BSuNfIWSX9lLixBeGfAeSg9fKMmt3Uc1bcNY5/RomeyreavnmxdsgWV5
eRj/33skTi9sjK46npZEfTEI/pDbUwZdX/cJGasAPt4M102JZhVpL3DG6CFoMeR3xhEbhkdXXtgI
PGKoWKO7sqt7gDmiVZ5PKgLrV7ocGhiNsiaKa5CzYip2EcfdCA1enZCG8EV8edeGy7WSr91udiMi
7vfO5nV0Mo2vMiymW8xUBYsrDSc14UZzTjb+3VKyGMNKIfF4If4bCQOo2unWXyx/jKFHQdUJDQ/X
sXd+434H3/yz7cVdywJQuPZFPE0KNS3f3kPu5LOiwvbdrla7JguqQL7qpI9E/g5hCsqOxUSdqarI
f2bOC0hnclXrbnd5vJqCaqrlKvtGrZ7m3EEuaMM86WYxvlcAVOmcWKkde3Uh4ZQ0xw2SwKeYHAdh
HkrEhWfaxAu/OptTxRA5riLDp794Ih7D396amxHCvcAhb9BJXpEMhd7d28zIRExgn+9Ir/RGyFnf
mfr+/EnTFfdbZkM2dT/i7FHZBL4hmlSorZ7JmJ04+b/7J3D28ot4GBKYWiP8qLIez0Aw8rJgakFG
f/n28uRpcmbgAVWKEoryy3w5pR4Pdaq86Ein6SH4AA2TgLJcNa77p2euVlgDxfesOcXJ9arW4ttx
TaX7+1iI069PYgfua+OVlJavYOzziT4EHqD9fjNRuoIQ74220jTmhl6SEkAoAy7oMYMCE7fF+qI5
bKt2wHS6L94tT67/rxvsh5PE8CYda8rQX9bYW4QN2u3vOA1cR6L65gxC/w1nLnGo9AOa40y6P4QC
YIDUTStpfK0rX55DEJLq4kIKwy+JhuaK/818r4TAJpsPFhaLgmcG5O9XaRXrjMpxplpl83D8v98Q
oAJqLtZXuKs7yo3zvdMNk7LQhURVrmKjf3fJLzVrRVLWlgPcJzWCLgRaagUc5k6b0yjuX8nEUzCk
7vRr1daIKtjJOVQd1p2ZJ2VvdmdnwLGF7RVbuTojZ8/T8Y0sVBbeUKxddpuKgr9jl2d9B2eMHOPN
j3dLqg9eBuoRaxT2HC0Pbe9eLzdZE57kg4WRVFN6DZcQN65n67Fi8yva3F9fzQtSWXiBhG4Smf3D
K2OtGFc90ZBmhWocyyZt+kyHAKokArYSSvtN7HfodA6HkBG9Yp6srZCp04nwzXm6h+BcMzL6Alo0
tKZuBJWN5yr2hZtJpwO9FdPRgTAWzdkIUE8XTKj9aYq1FanYRf7Nr+OYgYXaV8gW4af26dcrDcSL
1CW1ouIpGEtI+6nrqd9ag6VZ7IVqIrMC+Fc0hHG99vLGNNJDDj3fZLcM2s5lLN1cVvXM0iy/5Qqd
ynnWnAwsF/UoG61xl7H6bSX2o4gGJqhIHeze8IVm0r5cGXSGGL0MubsDBw4a3IPr+a3tDJCVumSH
vVm25PMF/ywm4+DxJKRePSO/m6vFlluABwVEffzOR4PosskeyUhyTeUmBe4NXb0Uui2zcl8UZDRe
2RWUgzQxNwWrQ/zBx21UCL1PYQydkTf1F74DkP6QlYNT680gte/VvaJiF5ADeG0i6kldSGI1Ucz7
KkuVFjixQbS+OriglIAS+ERCGTECYvaDPwRpR3oLEWTsqAtVu3pKsvHPuUBvjX4Cw0bLK8d67SnZ
xD4wMVN5vL2vSt4wt6gd0/P6PbATcYdkJuog/0wnRPvswH8AJnVuWu/Nqn/jNMbvDG9fuA/2kXGI
oQRUvTrf4H8is9YAbXlgqCgApgEbOxP0qxjCmEURvzwS0b8Yd8LIsAn77j+4O6TpLycdQ8YQth9Q
iXrQDu8crHYyoXlZs+Onfijq5yDIvjMNS055jZinPXmFAKq94pLCi5J097qp5MbGQTBNdQjbhTfp
BKMYK0/JIqxGnTcC0/jXzBvtEu3GxkaK/77O7dwyjU6wEw5a+rxQFbiMhiOPZ4CmB5BGDf5C5mEL
fgaaqqfDz4VsvD7VtJpzCbQdJVeqBJuDmhdMq6yEN6re4f/moM+514BzIhafEg2Q2dF9nW2YO0WA
pbdTNfNZoWPQ9DHNWmeKG1aOJ6Vd9GCdmNvlyqKn9BnkhYGF0rkYQS1/EieDrUUqd+TqtguXelBn
lNu7N4hfoojicaIJ2SLr/zCMi1+qmCYra5Lx8ydt5pMAh3+hwUNEEmqnjutmzAEGFSWBwH40r3U4
k1iiFIn4+QAQe+6M0yRAAOEVWV870QClMlIYw00vb5KmIV2GP1li4E+U/zckOYcxFV/ScK4g1VF2
0yVk4JsAnbXbBMBqiDuCERMbrrczTpeUKJwPZBkgMJ1NNqjr9yhTP1dUZjqYmDB/KsbE0sJCEGhS
YSgDjYMuMI20D8YnmaKF8nhwe5Y0YQhH6s/kYjHSgJZy+Yd53kChFfLXckwm2r94r+WEvqEiTkUh
Vgzd8IUVvGyLR/A+MC7Vdi988fGVwPtNDb1RdQAlDOvuGY7xrxuwJXOplFeSFcaO7g1sMb8b54bv
yYTMsF1slLPeDPFbP9ANnV6T47ltYsH8onjrvze6ZaMde20PEJQWbOkXsmuFtChb19mQDQOGyncI
iy9fUE9ToDWtwCeCfOLG+b9fTTbHkDYfjXXHq/SttArA1dx9kwLeOUwg2R70GuIwlL6Uspvkqc6H
6ezIMuHghvweLXrSqUbfmHUX6k/w8y7Xo1dfOA5WnA0k0fn/4/rJR8D30Q5QmXFcAmBPAVkII8zn
aNXLZ92235h4j6gWCHzN5I2pIqxNcse6ipbcUV02Vl3IDziJbOzY7TKHMB/GPFaDHMADH6bC/W7I
6OO/3hm6NIQ5pPVsFENQEM9U9L2QnMDKw05DDThE9mFRWrGWYm48hvWmGBlRCpHVmReSbDIcouSM
H/Sd8bsIqTsOyazbgeLG9C/V+TcHVHoa+KraDmAUi3nQeQEOGDpCZuyNQV7x9Cb5CA012M/eNvZF
sUa9zPwtiyeaEA5NGh5rpiYDdsZyD+dxcZ4LsTGVSTWc4Hx/kOsKy1jUpwYSwbCgK54x3y31dytr
/mepaClnNMoNVpJ2Thr2g8jrS0y/z+cr/zwB1PZn7KiWsBKT71/mirNbcHN6EqXWGjvJxfzKqsDA
XF/bj5XtPjW1IMkbZjVNzx9E37YkExIwJclR3c1Ojp9/PIusHf5OpqxlvxLHSdpVWLl5a/XVaee7
0tdJNkoEnQGsAd30wpGIBVy7mI+N2ly2JekiHYgmuPK2J8U2rptwk14bJMk3zf3sm5tPj6TjTQ+r
aZV81pqX4olZIho5ASKFKx2Ph2kqidCP+Hduftu3WGRXSzd8KceYhlwIgDkddDX9IPP2LQYT2qQe
d9gEplFFkZWBQfO8dcIgTlgFkiZsNuF75rPKDYgTJWuwesXChEhsabDl2FDUSTjAvFJi1GGbCDBT
9EYnX0zSbLj/LMt28epqWEcuKRqzFLy9w6JNNVsWcw7z6RF73VAArW2/MPAccPtRgq8WwHCgtg3f
/StBinpaS836QRkncuoyeC0M9ulkAwpFBvBt+7rTgTRU3XCIvdecHtZhEq+zcXpum9mOgDLIqsVa
EtB9Isp48NJEQmbKfW0Yq4HDo7VhNHzFoq3jYTpAyfZM7t5xFlM+cAJvwnUFrd36Jj8J3Zv8O+Fr
SeFV/B+RNoGa1Dh5PEFixZD6GML3zn9JzxUyWV+dGQV6p4uqcQpD7BBgsZZdS7NjmpnzVNS552U+
BwyrG7cAGU4Ghb4jiZTEwco/e+qMwm6pXVCdzbdALCslWEn1apLCSk24PF3TapdJqjQkmnf5ozUX
GYnHNRk8BTk4CkMhQFMCjKVYKzE7P6kbhFOEI6HfIzyTWlCbs5xz3JWpGqDUMr989v5yLxrQFJOr
UnLrp/B+dYaMV2jK6urDMx1e+1FPudyzF2A/ld50aYr0ecEejIBi/gVf/Rx4cYLYlis+0kgeMpJ+
bA2Gw/XXV13ftR6Nx5arKe77nQMwIHBS6ZzcSAG4xb2RlNY8LWtFhPQMw7HRxQ/zxw172UPYegOt
QpUwDOkx1wEeI6BFKud46THQr4muFfBpTaRywP4LV1t6ir9qlilGp8gcTHhub/QR/ugkYs0tbJYX
DAA6EkOkC5sjyMIrgZT0uivJwUg158WSn4gOXfqIbe0eeK0qeMyCBdZzSohXue2sry35GMr1N6zi
TXP1jaauQdy3ZPKDZw6hre7HqSP6eA4aIInS7KvV3kV8ep45zDZcerNDozxtkvaFQ7rO3/sf3OlE
MEBHjDSRkyI/y8szGHOmXeXbfx+12GQofauQXqba5uuN27+S/W/LXSxfM0dOuv20XfeaNuon+slY
TZyk5MfF81cScEZbQwXGqrjeUIYGLcsgL6ohaOilI+x/I1G3vXa/IuDHOjbsV3kAPbmcxbDCgte2
MY0hRKEq6dVKfaG/650FXs/1iCzQjj/4Mdv2ism850bAfg+UsjoLK+Dua91uKk8eINSlNjaXj84k
lwCf8aokuDlLsUxkuWhuWudRqpUyCsfYsN+TWwXW6yOPYKzbER6csfpsoU/HuB/d6PhlKXWG50EE
mPvGC7Ih5i+u1xBGJxeQ//ZdMTnIDTiy0VnV2yg0unA98FpxTqqREDA1ilgLLz7KpnsTaGtxbYmB
LgKhmFwo5xxxal8iIG8LKP6iMKp1nV0GqCY2BZEHMeduEBcz2b97bAePLUZ+16hrzwJA6Ie5o8qQ
+kxhfVXFl8Zp9ftkRgxYcx/qSztZoE4o4S3Y3c5JuCzkDTAS5ShPp8XS4naGJWNNKQwQsPIsEipC
rRTJziJ2FflSbsSTewBot/uktkBm8+9pfv1F7DEKxm7Sxy2MB4T9QTVSorwNTqv4eRALfHGXo9q+
3fMegsxemEftyc7x1i8sVLJkOdFskwQgKRWmgOjm0MfEOulPAvvXW48gKeuewYH2q+6KeA7XujBu
1gOojqCAuKyTmmbQeVsPoHoeFuvwGVJ/4RAKhqdjApsq+kVp6b+9HM92ZWKlYg14vU0pFwHSDZ5v
O0XUR33tPVExhMtG+1h9ICCIVnsAffKfrMEah0SFtalVvowumBWYuVhQPy/152j1mJ3fNcrMITRD
7GKvA4os7iOeDWHyli9iQ9CU9y67DLfvViV5o28J9tOhzCaPCbWgXfmByCy2jed3s6tyOr+EDBQi
NdjR9QpoYWn8fZEjhkX7KaCkYuReuVy6yeMzyJQajEL/wwKRDvqc/vkePqcaOQAD23DNQQqr9LW1
A1xg4l1I08JtOxy93jeVK6M0JEPEe/iGUZ4sUwZKjUZZepkU5L9IpNBudriF+MSiWrz6CSVpjpq9
09VsT4jVoSveakER/lVU2hEeaMmWveVdSsF8Czci+tlJfyA6DdDYHOJC7qUDYKh4LgnCpBzZJtFV
jqoTQmJpH8Is9EuhMxvQxzO0mAh4lf9wdVucwa0pKh2q9HafLOB30lAO+eslDGXBxfGt2NRXSmlb
Gaaqpdh60BZ6LcbAGQ5R2+Hak3vkfx5zhjw2+PZLG76WDgRRM7F7TCD4JM4klnQvO71zC0AsTNbi
qasYp6AETkwj4ZFCHOnPfPeQFK/gkP4zirjkd5VNIPFLqL+dr/Pf9X9WEc+o+4kPLcNUiTXddlae
BkxIgMVbkCDWA/Y40qT/3GhGTvcVcCwDlft1eUZvi7Ff/tUyFv5w3zyUU7HT9Q38UHbj55i90xGD
FR+xc/jZuGwhW/9rXoDq1yuJSsjERRyI8dQQGz5ZpUHJlLbuz5wYr/MZ5w/mpiZv28brXKCW97cn
b7/63KAnRHg6c1xTIRfw4ipiMEfk7yY1+Ur0g1njNLqyWosrvUSNUnHU0mHqLqO386xvJiWd5mGW
Xhc2nFN2U/JlaN7kFstqdpyMkNJG1DDOLYWyD+hJ8fJ/wRLTWaRH8v6wEnfz/ALaK+OMSMsPraLB
AxgJwN5tJfjy95HiZ5cDKoSL6kT35PC7rbP8e+jEmD0eust3bVfzAG51dK17ilK2COYVlIWg2ZBM
JLzD7zftg16D69EQkhXGlS404Pkvp4M6UuTPFaV0HUMnyaGgDmaI8Zupj1jOSGbGh4QAKrLtt2kJ
TYiPrej7gyirbseyTLNZhvNK6egw4hIq3WPTh/8dafjoTqDZXy+oIQcERL0i47tQs1SMcowHKrPU
hVV0ulj8kV42oEE3EyeqhLpEA6NoIIDwspfDlpRNeMU9WTq1iXyFLEE9ON7bTVXqVxk6pR5KjXe1
TQPOHpXeCOv5EQX2naU04uMaiPWPLpgbyRmbjO8576ljRTAvkY6c3P/YktRFyap+lPuoJyYJaolH
rl5ReUK0OlwwdjbmR3LjkRktN/ah4FgCZIzppzPgahgdCMQfq9s5KziVIT2RP9oKuQz/E9qlyhL/
Q2bTYxJNFJ7pMd1H7lT4P8WeFmbzbdJmroFRzuylxFpIW9hzC5VYVd2/r8HbO0ZLhdmv6fhJF8eI
lbTY4LMtvGwkTUOuiYAhTaIkkQLLaUkTs4gSQw7RsPX9IopHcHRu3oC616etbqorX0LLBYcb3rp9
xFvhr9YgNZ+RRBQQdxUKEwnaUR4hq5FCDov7/xZNeXeYDrAYYwWLHKzdg7I4+nrG5EM7/ntX7wCq
fVhCAzae9Mbnt3CjFeSnHlOU2GQRvnMPpqmAvY1vqpxVoG7CGJno6t8qKkekfe+7RFuo/49mZkWi
4f5JsPXNfuqpoe8T3I8YrTObQ09aPp92R5wpPo5cA6JrzN3LoHK6aBb7q93Kv8imjiU7pgiph+t7
5vMAn8qo2iJpx9Qfn/Q7KYbxtvTqO6bN7x6entRpfa8Y5+RUkzbtq7O2LgpL4xIufMKfefQgkCOz
uKNgxw7DGAR97hTYwsKbGcE21Cm6E9whcVTry7mVm53rnmiXH6DLElsTi0HQ1eXGql4wFWokxknt
A7JLEtrMsoQWqWBiA8LyU2NAn/jomMggQxfYEwqDiPVDpy6wyP6PDMfzy+MsEKHfYa9UNrqQYwoR
0zbDZWgIyHKOiu3+R/J2zC9k9KtIg0R4zaGSOMo7EYknUnEclO2A9cP9+GyZA0Wqjo6PvY4TBFQ9
g/CHWvgbz7x7uRqFpYR6+kdwbiph22/I4J5Xpmf6dEB6YEgrglS5+6pL5gF7oXsVcI7waF77sH++
mNUrYG0ZvRRyFo9qrmAVmTDEibb3m6XJSC+l1+PTAD2XB8aAUmlS2j4P3Vw3+KZYY+cTDiYpkWIN
moQeZhBLESLAUvtyoMS6TVeTZcJwL2+bcHTbD3Oh26mieTsjzvrtVSqzTVerd0hWSxyjNVDLA15i
M3LAa7cagaB8KBmMpOD6H9UVUAlk0ytGRjTZLBE3zfoVLc1z8OVLEF1lJ1IJ/rIlvsEFXoG8M8jD
y6xpzivW37ae2lbw0oSy5n4oOfT1ixGh87zDI2wmXS6flGr6jcHg74IftR0WMIcZTWUQohb6gI3Y
dWqKevWr8siIZizArfTPrPoi7BAS5Rqg62+fmUe3AbYG0ynobXS6VeYFCw2CrZLX2YOmWYenpuv2
GcRpOo2O2ZkiwPiuus74XbbL90ISAcBw4Mp2VzlCNQqmCwmRvpk9au9/974dUD3mSQlKkymGKv1/
YPdo+AF+WgfyN+M01WKSWDNHgGTs3Hz9IsJHUJGYKY07kLRjqKEGxAO5+9E3gQ5Ryby8CrcHYcCl
LG2+CAELiIq5tRYzNEms7CF/2SkeKMgE6xMY675TI8FPCjQtX7RupbzLaXhHLL5s2u+xogazbdW5
UgYnCSMO8LJYz9ncAGU6a2la5OKc5MbedtIMQPEVQ86CQekj/0cOnRPS3KkI9Qm4co38G4kuHnx1
0RecitqN+3vQIt+iIJHJ/dQYqir58UrNOwMfo1ufv1HFczfomIFbE4fes+6SjPomKjZQHkdsugCV
pqof8Jr4noexsq5ipIJHU2gsoDCPHrgznu9/k3dnh1qTK4g+Xk/u8vTTtrWtADevnBRxf+dq9etk
ZDxxCqD1CPripUT5IvJi0diQ39BjpoSc6A8T4F6ux5KCQ1XHmtDeaqcDbeB9yi0Ta++R8/RBQSED
6Kq7KD/Sh6e2kplGTDEwBJvRkGcZVXwOJnf8gsRzelAZtkIdnD73K1WQSIQZYFRbUzSW2hScMrqH
wjar1MtjYylhJOwV4huRb2ZUu/cxKhYF0XMlWPsT4bL1y20ODwN6y0SdzR5+kdGh93Y2WXYsy95s
z5/INN+03+oio8yE0CVtJ/G/d3DLuizWd4+Q1+RRlp4SQWV5n8CkUS2Wb+/JsNmuocoSgnLC3OU7
wqcEFWkkn58Q8z2LTvV9FPN7DVHmnZhYfUSWH+IuaspakOk42yssy6CVaXImjT40i1q+1tmlGlhv
J+tabCMjj1XM3DENeLJQ0qilLFC+aewWAbT9LP73dPysqYD1n2SUhxNeYjVV5gzCYoGJvE162XBn
8i5vEVm1FMM79gExJ8IB0d1vr6UtXJ4hr/LMvf1UCUnEeChaC8+6zqgHb0zeACKePMFn0HiNqzw5
ZdGq0V2IpeQ4SQ99TOAKtxhfEDZXeX8e6qv1k1Jqk4zV4do5WRZU4rBOtVcI8Y+C7gP5Nn1fQq+A
l82mF/eK0E+q3aALY7RdJFMTNwsqLvbk2iUZ2dOiEDqhwrYNxfqQD3u6hKWPEZTPR5JMzMK/VEpO
QeNkp6IGVX1GJZExBvGrhC6/PH5vN3f57lF2kz/H3p+2duKGLBDxaYbTGg5oiAZ/ftFmJk7T+3C3
pM+SwpPUAuyABLggGjpGal0ollzdqmDaT04NeUqMBbhun8AcMsElRof3Xgk+tK98iTNWAw0aUo8U
hrvEH+5ngAlGBnuhtCwCNg3NSwgc38QG9DPqGjWARewip/d7uH1+n7c/opVPAxpOxEJU2JSUQBTf
S8aEqQ8OY9wNMHEK1n51PbAUJKuoq9zODXeGgKFVzvRbflT+mgySiflMBFZ3Xhtfy623zTHqEcKb
jx29uFlqQ/SgUVoJLpZjeePMqx0XJpjud0dZLdJuCOoDrVGZXp1zW1J458r4McSryHwJLvHq2XNj
YwlIHCPQ3lJDunhZT23+nTivjIqfM351NiF4DKmEKbpjknTV/Sya0sqUrc1L2bcOpyZIkMR32c/o
+Dj3+W8am2lfTjZX0Bpv6gqq/pqyko6TR+uU4uFb17k2J3Z15iG9hxpg3HWFezCoUA/PNmK9HokH
QZXWcDawuiHpOvI2paD4k7QIytEyUuVhIOk56cqrH/loa6xDcSxAEOHUL3ZwMiSRJMIrxCCEgW/r
+HvG9mIB1kJWnbENH1SpO+90R+bgBy5in1KFu4JCSwUwU/rQpWgg6KiYZ1ClmtbLXxzboF+H/cLx
g/IQGug86pp/raQkNXYXDe5RfpeDcHGVs6ZCJIA1Jl7jU7CAuzU4/F1sdgGFLOkJjXtWeyC9xl8T
qCisqUUWqxc353kxjYugJ4ak9hAPrYeBpGUYUv0fbmTzJ7kom1nyEnYnMqEkVN4B2OrQj7UituNT
xO2SqaoI6aC3zeH8qoo0igmN9JyKVi1AqzNW3FRQKzdaHq9YwN50KFnGnMEJ+inE78G9/VJ7gM7J
WX/cjrXWL98iBRx5Ai6K0Z+I8CQqF8EvvHDM1UXyQGntVvQ6PVLPit06hsu4Oe92/mi8752TWkE3
1z2fjSy6UE0AgSbmf2EqgtNb/ncjAoYoAZmvYEBAgMOnky21Qm3gZ0zp5EI4oqCNdBhKAR58nGPY
pvnicjkkIrn9Ku+hH3tb5Ny3EC0HJ1hEGtFEWNp3NhDo3E1m18rA0VbhzQX/vx64aCc/aOkklIjl
wHaXovc0v5mc3qKiYI0/zOOFhozjT6gyA9sQVl/iKJY0QF0DIDjPVpmVbUhw26O4fN3Jr6WpMGhv
uuUbL7943Kdo903tZPwZWsVPR20v7DavbnsDyR1PtyL8qgaR8wsiAEN5G4XhqJayYfsaFcCWymjg
1/c2tvmKkEjx1qunffM4ChJF9/7Jd1Oxs0QCLJGx0HQh3b/Fo0PuwKtZHOm/XXe6D/mhzdnr2KyO
GJo/UPnqGk8qyPbbl96AVAmp5IYXUdyX6hPsFi4F6JQsK9dHN/B3kcFckcezDGndU07MieRW5CKI
5+bLkcTlAjN4WBmCt15zmgj6nMQOCFlHjGnY495SRwYHv/XLsBYLn8DdEUFLN5i8WU+R7DmUdNQ9
zOuar2wj9XJ+fTwkrheSmER484ItGXguEPY+3a6ZnhVrb3ZvcClPSwvZdsevmUcEWlOtwqtIMBfA
eNTIfK9f2uEmEoduMZ4lD/yXgo2hryPZvi89yQZ/okTq+0HIMLX/iuI1cCLyjONGIpaU1MXPCdSI
VeY25d/R6VXFe+WZxPvb0vAg9MjIKU49WYRXhofRy9c9DIpSeit5b4L/1dM8RJJD+piZQrcoA8BF
2ue6UVwl/83+HC5+x4jZPBa7Vy8kG1r4Pn9OSfgvvZlb1wQ5mceTrcTghyLhb/1rDBJ5gdP2FtgR
rR8m7WI6QLlhD/Frp3hT14Iw67PA6mwt9J0hdl8voShqAP8D4nOX+tiqPD/tyZv/tJckZ5p4yqX/
yPIRzXOE0LnlDSv+19qcN6U5LUs8OcPQ/dxZJnMl0Z3/vpRUMA2YhWQouZFo+bYmpRjxMU6ZGaXI
iu5E0XiajWLVWRlpD8F2L34fALB/Zkc5dovC9/TaBvQsuFnicelBYAE9xHRD3/F3Z8xb0MnOhIHr
4nx3upuowFqpdh4pNdzkESHiKoluGVpOl5QsrgNIDsyChLtl7IZgYHF5Cz9BSYvFZzUvGHM/lv/d
SEic7sf9V+fMCdKp96HlODOahEtnxFvaqbexEyLAATKZxmuu1YROvnIezmcmqiNx7iFw/aJapj5B
MaDcmO/hmkE0IF+qYLNpz67SsxbITQpKX2U1zc/IRYppEBltyOORsSu5gka5n1L7Qe+uABHtGF4B
DqUvKyv+AAoRbjZlpbx6vrVKTgPJUBdo1Ae6G1Mb/wa571Mtnu2jgAEmoV9L78XhPV2baCkUTMoX
rGQ4aBiS0AiJt/WM4tYLJgyqURSlVh6AnNG0YVn3qAMe0oI/NVqfsHQzmerBfF2N7QON2hxy/hOu
RXvO6+gxoMozQTj/xDgv/YZPKjNatPhvaUZ8xX7ca55FyqbidlVVBt+9Zgj88fyORzCJeiDpwSTx
uaJtKC+Cm7PPCwGZX/dPrNJURaiyES5oY0X1ObuStvgZ7dTujzcjGGkK+o5QZGgicNUJi/27CQ27
S08hCXD40DqaWgfAkzcYA7SIGdG1AKTOYDnnqHfOcoKuz8ilSWtvE/iVYKlgraGDu55uJgeEOZDG
ezB+ZsVBLofeyZ6bWiNf9GZEt/1sSdvJjRxcao/0gmKB9shjYvFOviMSqpih+wD4lz1z0faZbDUc
m+sa1Fd/ilpT0dq5tLsAKeBoZvMkQRgdwLn7jT9tlJTWj/miQ9O6up6FRKUxSvMS8sV0CMyUTTcA
LgvNXXg2+bezCQOCHJaQiZZ+aZJyRwkV3yEaAvQRW5uSu9Onq+LWNYaBLu5Q5EnpFmOZbYJzC9H1
tQTMdrG26bg7oVggkuMHXVy7XU1025HtLUWlo04KqSNrkWE8Xh5r/gYajZPMjvjJusDBAiShj2y+
MNBtJIcyLGrIgaE7fcC4z1NoSAbiZZ1QqqQx+/7pmOnJyXxrVKaD+Er/4L61r8LziEcrHGX9dyMh
6KMz1xRmwV5+ZqCCWqK/j0Zcout2TIVz7GWeDfO7iHYtuYcgDdl5igKB9pw9RJxQ+fxZ0hzeGfX2
Vq9A9wgj9mX1GrLx2NRUBTk5v//jFvv0VXiSGcbmM2aiQwOe1BJKCpAijxNhljp5n19KTxQqn5yi
nrS88h7v0UFAn9lbrOCrRKPiGdzIucRpln0AWO7twmHhmreZOwyxxef8enzTwXZieIV3N6P7TH+9
fXew2P8CeA9sOezpp+UdGu6hkHg9Mw1CvZU/0GHrDuALc/plPkLpGEC2XEBbTof0OuckKPPPKTSD
uQunuuJ29I0R3zJ33mhcGyBVxSP9jSRh6j339AJW2cVpbubJo9Uq7V1jcvwGKV5xvR2qfRB/tGh5
3nWkhrgkiScpdaqmZqdPr59eKiDNUO3BjGWUb1bHksPZuxJjkVBnt8P8P2gozsqhxUV7yQ/iu96H
V53phv4ST/c1myWv4JpbJxGVaTI++tnAwh9D/lM5bblVqtA5s02xlAAwwmYqbgTImosoWgEaJLFK
dgmmw31cjvlZ+qvEffpf0JWaLxP8ul+5LUtzJOrE/7Dq0vokoqtCUITM5pVHCtBMz+u24c9jRuaZ
ED49UZCkGjeykVYl6n6SBnbkg2emdRZ5KWxf2YfzFTa2bogGRZ0KhUiDgwfumi/1bZ3XBb5iQ5co
UagOidYEcwKz+nUX1ulq/Ciri752gX5mKL2+G7todBW9CFydfc9r1paI5OOfF19wqX6U7CwpPgRx
KupyJ4o/C67vqRF+V1bWr0t+LO0SvxfK2O7/gEsggshPjN4OHuT3kgA9NJqD/nZyAeZjfZoepy0J
qpDEP0FPb7WK3aKsbd8Q8g2bbdZP7TkWotayev+smq7t6p/P9HiB6cy/C5+zvxtR+YMd61ee7bdn
xU9P40mFE5Dtnhd8aAizqzbbYfGPt6j2P+PhGqqKtR6sylEOo9m9xteF25M+oYUmRriSYGoqbZxY
Kuuu/YnojfOgtO3h5HPObGJTvZq9UbLaKwXk4CpwIiaaAqDcZI2iJkEmIN1nPGgVUKu6oXSQjJc+
WirP1YXV7WLAirNRE0fhpnqXdELWXKGtiXb3lT1g5rVxDt6sAlfOS5G2Xywg2Z1kwQQMp8k8ApV0
Ujs1EM+e76NQPttNKNpvyosaogkkaU1syjGRnmmJ0D3yoh+uIEL2SpguCB0W7dux6/XJkamF5ZoM
9j069C3hKNDqNCNscgQkhjrI8U0KsIiPG8fA9xvB38Y/fhHOdNuUH1loxciDXrYbAB8JE8ZvFn51
Ki2/NbTNlM/Y0gtVA15F6HaDMwdDlMgrd4QdDeDn92K5MaE/V+0SZDVC24i5RPT/7BCysOmhIpLS
Q9YzoYIGu4b7fWyZh34nOJ4OyAtglYTxL576XxHbLj29Fd/0ZKwjTMoKoXoIgehsGUciqvQyc4WV
xJlXLPGmlqtVqnmwZvlRY9zBFHhRKy34xaw0x6vuaEKM2PJafb0UFCKhKO/Vnmoe921+7vtFNv9x
/meUk414ET4e+wGbs3Uh2Rz73eoznMyOxGYhEBg1VfvGFvxXs1/qh2/4zbBdrumJ1KmOeXGxUo7P
hwVVgmkukBk7jSID+eBZtMeVUbckVQfdeSXozACpWgJRGinKQqeOYfJQbFsleYpOpKHdbJ8w95Fd
9BBg2zueM1JqNZUDGMz5RuOI6YpF928BsGlJ0tvI5p1QwVnOTowIdHO0kLb0lL+fSiTBQRVOrK+o
DnkyXkHf/eBmaDlyKQdPWn4UW5/UsuV+3Zjvf/D6VpjwgE0zihfJSpiUxVDc+N8mDlLmuJjiLhj9
C3olMUBSlzIZ1mu4s0JqQOCUGHWDirkNEo9SvNrw5BaG8IPVe0Jx447rMuxXeLI4W/tJnt2Bq9l5
6ROOVNBuOL86iHRvzBgJgBCzdg4Hn3x7XLIU6Dm7zF3Kxk5TsSwvrVUb/LL1s3dnvN7oSggTRqGm
Ozp6lIBr9CzdLqC0+jsCE/cDyNJ6glchfZzzsacMzYnF/VpYqsUwW3ES66Y8IB5ESnlUWGr2v7Og
8FZyVWNK3lO8YQBjpVDoasHcY+Mvok6H1kX8zXJaeSsrQ9acqcwObBWOXk//nvsfU9Yozf8fWHbw
VaePB9sDMyghNeA1nHkBplb0A1/nfDQ1FNtj0VTHsYOMoUsSd69L/8PXu/ogJJ80UZCmOUPDNng8
u0934wOM7KB282czDjvTVILGdoP2QUYmcJReOa1Td32FeGkv3xQLXDV9JbTw9Pywh4lGuktC0nN5
8m7V6SqxQEKFwe/I5Ins43eYqumIXxVfm/1lHaIdoRhaopiKmgdeILIViQ9mUmme4LjjfjSUVMzZ
87336moEdVxdknKLj1JO5kkqZA28DPimHFYfDchDPdTJinV5PfB1Wo4MNpmVyy/d69oGKKcEwK5W
pXncX1tXkY1eD/rkgVvrxznio5Nlnrey+LSSU+kKCG7HNjVl5mS4YXXtGaZJ844CS3RalYfKjh5x
5bs2XIVNNjhSZw0vS/jjEM+J7c4GuT1AQ2+afIPUI1R3TTMQA/XThd18fmZvCt7XVDeiBkP8i59L
UJoLxYFmnK/IWrlIaHic6GIc/qUPQ80R1H3clwW3aTVFM/314wqPxrZPSCp5hIHgb8VpJ9EwAbep
Ss3B0V7zQvprTtWepJHcpmr0QQhp4WmNTh+lPkuJF1Ee3jpE06VH53VE82s7gmldMqVawVrYX04M
WSycDv6FGVFXnddKsLjU0xHB3NLWLY4K1aEgTeFTgsQViTSaJQ+CMEDItsuVfe6A4zN3YGmkLdE/
TiI6DTFNd1Sv/835eQkkChXdxLDazu2/w18ODNAdiTa3P3uQf1FcPHA9pcEGiJXbKUmfo/PnNsod
FJ+PeN8JXivXhUh2sG5JBz8lR4oA7T2K+ZZlu2TatxDQ3dy2TlUhFDtsLtcY2uNEziNF0RZunvT4
BVsON9o5KCVlF17GmNIRzpatT9arSsmaf8WwbS/vnx7jfJl3P0OOGj2wbVu1STdUhfFWMPde1Tok
uMetYPEzb4md+EJsWIBRtdYQRINfWP0kZenR3e6y5vF4j9CLUGiTIwfb4ME8bgE7e1mBPYDWl9pl
HOgEEmCQ6He55FsL5DyoNgEhvmcZCYdUS13zaVoMN1d58uOzystVdGOegsYIpf1CtAcsNjhTD5tC
cZ4phEdExjCUj/WxUT8VTzFzd2vVnhOXpVqtt8dtUAxgU5zI5PIWYW8p5/J4xb3sAyTZFNxHFbL4
aQaYwKMhorXTzRM/nlBUk2fQGYmnABI3fd+aNc48A/tybHHpmZEc+4/IVi2syf0HoE661M7mfrQF
TLyB5CPIAUFWjf039gWHDyRaR+mqbudwZR3Ft71OVMctZS8fLPLS8qj52UFelVwr7GuvFtl29th8
rpbPUs9silTD+dCskECg+BhDkxwwg3S//00axiqOe+7hLgk8OVsvh8HrPFt6it3Wtkkzi+ZTWm7K
XgTEe4v1+Xjs3VHrpPauebrIGUH6oUZgwX80XqHXuaV2+zbdxLTqiDb1nk8+ay2rglrALp8YtCAv
2hs241P/xKIJ/HxRaI0qhTFOgA7HxTBhmY337f3Iv6AOEcFQT7ycp1u1+5MCvBU/33qUDVSaXSbW
ylchsxyMsZGymIWgsginfol0G0U+ihK0iak3xN6V0S6VJ1YyAHlCCvSClF5Aa+GvwEQA37eDwq42
INGvBudpjwVbMIU1EmAtQJrqKrEVKc0wBXIoggHRDeWjiLyhDpMADB1A99T+zyaFedtq9ivwfwiS
tNH2jz/S5iXVA1q5vJIDMThRmFNS+Wu5FKrCiQzMn+zo2S0Bg2O+GGqDDsc2bHyIFxXUlHJcXIUW
jA7DAY7eptgvIduD15YCaqm9C2F6PWLGMKPuVN1UkyLbAlc4+cozIU4mQ67zSlSF0LdXEm1Ysfkf
I8yg1Y+Opwprc4KEoAvrlOwKaaPJ9S98c0UBYIGYNpoWREdUfMsWww4Otz7jS3N6LEdYySelYJJD
gaAP4tgsAnYL9HZJhrFq36vIe8aRZfCV0hBne2YIdlUidf57PsFgmBPkG9BsCx+5P/Jh0l2gDVoR
m7xNwx6JNlt2jqpXDDF7H8KHvehUzYiLSlMoxprpM1fSeRKC9JOzMlpeB/buL3eXM+oRaaJ1yHsT
zSLunZ8c+h203RpejpWi41Dc/G1gdGMI1J2fgQUha+zA1OnYz05KpaLIu+aXM4u6BYLah391wpU+
0vqTgoFgMIqciJyVcRD6hittHUFNYf+bNiSlS1XiNhGgWXbY8CYOPsKKxiSKZCk0aqzSkv7FLW/Q
UmpTmnb+Bp/8gF9rZ158Io1UwIs61V1QyRmZTNhIxDky59AOrNPwEa6yuinV3Oc+QmSfV5waNtnK
H2OpTJ+dEaiwd0QOg760N9oZtS+cwtnLpYeljGR6w2En+WGq/5FlZsREkUXjWlR1sL5bYZbFkoNx
MZY+yAovKzxJCBuqm39a0UIULnC5LyvDM1g2a600pceYoqLHXCKWLv00UNwFLT/iCpINC8DlB6FC
Y85En/OcIILeJM1hTIVyzjnWP1IqNqcugO4dwMxTrIUvcsFVAbq0yr3PgwO3SluGxSTVzqdv56as
EmuYmiggCrNxr/AttEOA5RfPgD0sq3qbvi7bmRu/+l5MQreH+pKNb6K7mVmpxK1CBHQx8K/CyKVC
FaSk72zd/JGvjwdLGUQuGPsKfWtJE7lqj8gOukMo16muLBMBSzt4O7pp/AlYp1jG7NeVscnJgOS6
89pd8UcbwZ7jRc2rojyCqNbsyBxFE3zMkSLUaQ3YTvNmYTINAjc5c1dFYA/PwC/qhcIAePIXmw51
vQyMjTggDjLTXwfu1L9Ozh7aBETKb5ThNANInNfNlM9uWVScQHAlKgNj1igOaJglvqv1RKu/zw7h
0Ufy9RPzHOoVz0UBzm7FAXDsgAOH07GzAwa7DlLBM/Fv8OL+HWMYH2xvOfEkd0CbUj5b7VL93XTL
agILF3ajgTxfqAHF/c6ba+bqWWwlzArxPbsCpP8KeE56TY5oLl94ST1y8bBFHkl90eIl4RQBeBy/
yDgM3JD21dr05uaJmyuNIPFdXD2OQ4ieu4DwCm9bI0xcYnVbX3+2BWNk639t53XNySUk46JbRV4Z
NxNHbxgrNRicVGx13V4fGAldQQ4eO3sE+7gZAIE6TS4T07nJw/IsmRoFuqapRKxjSfGwWveRm+KK
PSAeHvsGocgL5ykrJWa6j3b/b+w9YJpVnyGXtmIZy8NyV8HX5YkzzZoW+RdW6TrD7GpXFaSyacuh
F4IG+H+/QxH8m6HxzWyUcvFs+eX4zYmN7dn6uFw31ilLgJMf+S8Ot9TPDPCOGbeL9gbOeVb3eGg4
15XugSM0WVMsOfBcTSuMoF5Wty47uTq07pT79ApeKeJOB6ePOMaAlNks5KlkOAeZSupLUzs60560
So/a3GvxXu+gajIRctDIt8Oa+JnrBono64EHY278a5mCrR8WltxJ9wwo5W2bDOr1Vx638RdjboPm
i33VkR1UzSp8bEgDNCdm2ZSRuDJD+j+D/RdPxYYgQSGXqtT5a/deUqhG0DEpNqcWGnPIbY2G04Sg
WJD+xIby2GFghmwbqQ3J8NmTUehxV6ZUbxpZY3nJ32FNuJmlocTolakpUCzvI3UV9099DRyteNGn
L9jZUNSzhHYSGgvHB97CTEpqwkIAtrdVglGLNNhtN4C1jJGDSziEg4cDZgQdDqZxj+qmPApexG6j
iAsOrqqICV0RCokPVsGnT4o1bfRalWZdXStk+mxKcuFwVy/VP2wUX6tAOlowxEdMm9YmTC419mU7
A9/vK/v9Edbcw7wyorpF4m4d260GVTZbqhxzcY5NkGdi6jXRjgCYwJnqKtJsnc66HwE99CErG61m
d93Ipbk8xDCGUdgoethxtRAZUf3OU9xbIZKLcDED/jW3vzRcdQi94OsMb9R3fV2ClbCbNYxPPNVP
cjTUg50RdSoY8J/2wEiz6dFOfOrGyRsQPnz2ZdiylAYvMGrx4wJQZPYh2gRuf+vpUcVpZPX6Vxk3
IdpR+S4aehupenD3XzCv2/RU0ycryiX7/2jisgXhcoaXRvU8j1STaLKyY1c7x1zOPEVfjvKe7wmq
zhk+G+pKnUbs4fo8OYryuzQkKj+Ee9vEVgbQA15q67f7veIhwW8i2jdCAFVtiLFnJrzea3Cn+2e4
u5DxYhgXfcTv5+T6jMXAxUDbk78IKJCQpUIen5NbSDuUnL3uDCAdUrvzlUCWYkd18+0An4rdUlAe
I53EgqML4o264m0fXdJONppve4lBdN2FvQrB4kESmHRINM2MnOk368n6z+lGgKeTXodLTb/h2LIy
ubfaUUWlzRANzrp3/Bek0bm+em4yroYDPQ5nmv49dkMbPH+bd4TxtBoioJTBj2GE2g+YVu3XH8bQ
6fYvV6sD9M2gG9xNPgK7FGJqEPdFj2DjntrlMqwSXVOQ4OI4oH7B+Kzj1fC6HjVne4Qn/5hPbCbh
VhjfVVD6sWz8ChgUAyZLnKafrlybBiCLhkJexQMHanWOm9PTFPlh4D7hf6faOlNxRbAowDwZjyJ/
HGt5qUezkx2ycaOblKn2WFkpCg/ikmMmEGI7dhfjFCKYo/ux+n/If5ibTxTEPBW5d3eEzW1rk9UT
wQkHTUh7ygtaAOqIUnHLuCEkklafVbFOvFi+TBSlFPsjGNqe5FQ+DHV0NIcsMeN5FhX1de0hBqGH
XQ/Pi9Tu2BWBCltA+2RFejHb8/WZmG0YEpgJyax1N/8kiy4nZXWYZSm2Ca2KIYIYmxsmGHIZubwt
pIhYD3WOUVxLKMtl9QsDSSX+dgBDbU3hSvWMYtM3vVEIeH0vMg/l4nci056n+q36Or7QoX1Wf8b8
gYql3MPDItvCobWngD8ISp39336egPajfI/F2hLKCoU9Pmq3SMiWc8wiejI/VsTDJOhX3e/vmkJ/
Hbmt1Lq1azhzLi9LScp9H5ypnc9SdHnF21emjE2NudfdKUmtNzQK5F+Wf3UJAy8ICZFXLSUW1Xft
+V7jHMiEbEj6a7goHUigx+VtQ181THG0Ehzi4p+5yR25mfzXb0a0FIhJx7AKcdeQvHRWnQSuVX2R
oSaeiTpV/0G+g9ajA+c1GaoHMu0GNFUz2ZL0Q1wYlnDhq5vhizUK6KONgG2Lpc6q6OkPAIqX063k
fJgESkvY5ogEB8NbBsc7uGQHQBP8YokItCIfhxArsQEgG4pICUuHTGp7i4e0El3bcalmbvqddIWh
pRR1T3tGSW88MLEAaGV7oprfSbS7eth0HB8mzt0+awDhVAG8mP0AaMnmNX02iH0BM3OMtgsqj3nW
KNic/desZ7NPGXH4zgaBhGck07GFTfSM7m1zlszEj6PEPBm0afoQJ89oiegOMhWfq2xvQwxpEROq
7KSN9dDLAcoMSZU+rzZDah+G1XJ38OtRI5Ei6ObK4QMzWo5oyoD608OgTUO9vuinZeVtesej2g66
D4q2rHsf41GlTrsi1M8xSwDZmAGHceHbi+B28etHj7KM8P4qN4BhvcmG4CERWcj0MDl++GqYp9Sw
nPR8zGUmhQOGaTxWGmujPWOvXnGn7KneiyHcfFN+8TiEx15ahmz5se3qVtXv/hOigo5vHPTM0F75
KcEHCapZ5nYaV2KIjFl51teHK9aKlC6hHlLAW3PYJxFGiU9NTjUr+C2k+p34c0MB/hOiADwwtYx9
8rYapo6xPu0RD5WWkz78S/MOtgasaR/dLndWDmdNg9TcnGQParXRryplQL+Ylv4sDGlPJ2LLniWY
p0GftnKvkI2AiXOzk9c4XFKZBelI0IxGjv7uwX1DVnZiwJp/D1lRfFpfkt/Xadqn1LGeaMW/5InE
1dYMDnqALqxN6YJYJCuT9I2GQzQrBZReOivVhAth3WHewYwOgPjk7mab8dCrbZLGg80MCM8vZY2Z
SMjiELIxSKBWPIWjT5iPbQTLmfSNZBtmtxZvBW8cYHbrA6N5EGOY/TxtFOCgVviKgv/qFy1tdvJn
MPNHTtyQEYDw6M8Pg2KHZK9XICreKAb36o3r7Pd8w12DG0yXE0iA22aQrB0eGy4vX/8CSc3h3boL
g2yOR/sTqnj9whLFWii3iDv0WdeqpHDFpcwWIi9RzvsUuRkl69V4Y4i2rwQ/NnfddzLkQ9AY0O7j
sW544tv9a0PmtTkxNQXJXVRgLxcCAQtPKAX6b0F+eBtHTu7b1xoOXZnj+gRvri17r57kc+ZVjTsG
wzASjW4z16FGkuIfbQkXfdxTCUttboq01HbbyJnpZ1KOVfmk4dJxKM8tfjvto2IK0HyPCY7kVSGI
GUwLyulWcNuxhGANk/JTqszuN5/Py5cuoiBfAZrBthJAMCRAjZQ+vcvXvA+DEV9/XideQfhyON3P
HGr/832PfsHXbHu2vqG4rih5YHUg8NKU+YNWAjFw1T3I3LzMKCgRKIXVuIctAXhOvSc99UkVvgJ6
EhRHjE896c9fs8ZyyQWhQPauyySiXXXz6fyKbPbpSmRPgchNh+pH1H+K9CQ1zW5y45YCfIqwUgwU
5erX+Gqs33z1Y4IG4UDuEQZqKqK0wXACTWjRBNXQNSNh0jPL8gSXiOnf+LgXaobMmHgmcwyDOjqV
HSrtmmzz+ToDS8vHqNPU4fuIS5Yb8q4v78UH3W0JTWV+ZGsz80hCYj28yuKExaspcSTUrNFpz+HI
QhsSqZeAgnLTiRRDqlxqkNq7n1V+XLs8V25ptcQytbsAwN6Ms//wj7EDxz/mHo39XAX0QUOHyn64
WqXlOZ4Q9cm4DBbK5S+yXLi7kgHKFxbVY+gEb5FPBuxawkZIMwDMVmOalENv9psqVverMRWsM0cK
Ai6Pvt7ztrmSBFeNM+a2i+ZnlZPyn5rwtPL2mAhVmruk4yfvCzfV1J0pXG/STzUmNgaAXafPjx7e
gD8rvdCcpWWmhBv5qBNnlPBqr0sDOERfFhFswaSlHJkjwYrSIu2MuJAW5Qv++IJIhFwJ0piWfpoj
2ch2Cwahl+GiYvV6IUcqVnfhoDQnrfkmiRtgDkE4jnt/Vp3jdNCW4Rm14LbI7ZvC8obFMPnNo1rG
rCzRX2zcaWqUxY4QlhcLcHo69hKM43rbKQVjYB+ng/K92ZVjNz93/Ay05IsjYsEJRd9b0lClojCB
FAsU7+hyOwZawR7TmwKpgCrGJ8cKE9hneR/7V/HBoCcQjq2sPrp7UeneUZ7BVFg5FJYFCFbM/19y
uyLFBKyAhh+M4wR634CKbA/R0ft1/qCrJr6RmywJLjs4HfGo3AxcNDe/onu/JieKuu7T0vFI+Oru
iudKeuBCJxoX/+47u4YRk3aQoeYZmIZeEPYyI7Xkoqqkq0ZAa7y59mg5MxP7j3fXTPZIB1Vf45r4
CV0hBsXND92msT3irnrap5m4d36ykE/Ud3obWx851KDji9GMdHqvXk5/rco5mWS55WQbknYV9u8z
qXyPTLGgEh6cNGGMLLedg579vnUcxzQjeVxjT1muIT0Ty0Ksa37KjzNzCOw2XPrQ3XspAFRC2sDO
c0LEVgVobbOXVrt3wGiho1ay2wKZ0jMS/X4hLmpKiskrCfR/mp3pd3oZM64ybgOzIGN/iWV4venU
K/mQBqIObXpBVBidWwpGnq25n6gKFpouFucEoLS+xHXwXjFxW61owH1V6VDd7XdzV18JfVgW+Jhq
rcWHR9HAdGckGtnrkNP6mkdanIRF6YwG+4dkov+kICdgpcleXH5Al9tqhG3/eQqWkY2SB8JuqhSg
pMhd3hpO+qor33chcNxsx761QqcaciyPqsA3f1yVkJKfdEAnHxcEpUBCY6fCUG9+038VeCB+zSdM
WiM8wUqL0fn2K/sp3nR16IccSsf3uYT+fz7HZDWjFog2/wzH/44Vofxsq3Y2Z/sun5NWEKKpBN4g
jtaOK5URyI8TPdxVRIn0sIMsNiwlq2oJzGlBTQCbPePrmIj19C/oI5SOhOcddSaqdJ+w8XH5Ykh6
bG7I9wWNgdIpqsiJiRlYiOPzLAFk+bgTLD2j+ps0vXU+tZsl9xTKhD6RUwMKQ6ckbfI/5JZUzGoA
G3oeZALL5027R5aiSd8TPA/VDh0m3RCdNTIF23sJ/evGNK0ePJrx8rV2zvzP3568rP/zPWzu66Z+
VWHPd48kvcYyndLZCnQrcf4ri7CRwlDlkXj26qNupV8Sy6dS7zWEhkXcI8/59ko73r8fybAPdv23
BIfakqiME+eLFI6o3lW9/yLgeb2WA06nhGPF7SUZyV5MahyL3eXHUfmHRWVfJmMw/3vhMDb8HxW1
XrBl1QPhSV+ej4bc6cE0jc94M8EY4kD8UnlyR84IbPFBWULJ6O+yQ3DFECUm1/Q2ejg/KzlX+Y2m
V1o5HPK6ufsdZw5M2gVNwTVPeosh9mr39YiqQPgoktpxs6jO3lAALG77dUQAwZBh0i6+gfdKQbqh
F+aBQLm9jREpbutRiNMlThY1aXR1jXOkfwV3Oj97Y7uZ2N/Vbs9tlJrZIGkRGYBTy+BsS8L7VZkL
/hFAJB8wDSq2meQuvovYG/+YfR3QOjDSBiU2//8enEEQDcZ6nJFTzHFOg2LJtd23Sg69o4lTWaFj
1lPW9VeKrkr3lDIhMOgb4iDcYUS8qzV0MZtqIDxDiYTC93X6xQcuqB2im1hg3+qbrgLn9q2iP7Qw
0ui94zh5DDATAeCfNdYtjRaikv8aIR3Cpc+TfH13PQguTUmJZSLPx56Nvkpz26LSvUNoiQYNUf64
Qlj2sEOTqAmDSdzlv7INlRmFZNKL9ofLifgzjTrj7K69bHxion9+FWwIrs5mA7i32sRkpUzt4GDG
tRbGyJSISVKtQ4zgug/F8VHqcm8NH6T6ZLPhdivKmezZq7QWT9JaKnNUIZNlWelT8TQzcNF+4MEn
ZxryMNkElcqzMb5ycRYB93ixfSw703yawzAKzbLSeCOoyQ+pH7Zhh7T+Co9OMWsg1LSUkNdxgedc
HpLByhHHIeS1sq1jOcZmq+w9YKI5whNogGEpmEga75gvWQUgcm3+XUeNB60Bf3mcqeAdBkWxMrtA
gEHGdlq6nd+nckmwNH4p1AahDwbf+k+ZC2cLS2rJ0Jn/0X9fWbiik6XFozkEpuYsla/3OaGZEJl0
9EcqDrBSThMQDSZl38q7ESgDfrvEzN5WBPdRfN/4ktWW6hZQtAnogmiJOCyBvsZ307lAHre1eEDK
xuRNs+JZUu6o42dLfCcqheTm7aloRYVmLbJJJ/ebhV9VIGn72JzIYmsSQMeCOtBM7TV2KacccgpW
qVh+/+qxgd1KrNlI9YNAzZb+3rBtLakRYDIYGyrydGEa6zDPp7vYW8LUcjx4hKaKJr9hoUd+8PPG
V6TUTh2QGH98fPCvSTbhwu6P69p+7z+RpO5zQoZX3/Abb6U9OCNdJNeOIjQeP8MWn/j0fe4PdNau
Zl8VwoAeExzI2j+8fuGfsZL0/YnCKROKGtjJGHZvIyF+5YWuZi/mikow8sSMnxu5Ox5eGyOrgNl/
83pUV3yk9rxZrQmS9LQkQvig6D1K/fAhPJdsGKIOOn1KMDLiN6fIR7gh5+YNFFhHsYxRDN0kPi3J
w0BXTHzui4GsU5/S3mVKBbgd+DR3cqFdEmHdxqetyGnpXVkgZ8vJbIPehRqrskdxfoEoRgtSSgN4
m/aH/c73SGMIG6mkfATTOJUwK4DYbjDYhNuGkSoeAARS3zremJitf8E478UadRQBTEb/deogiUp5
yN7fJjCPpoeg45qP6RPACI2rV8xy/hmt/4NXaAngGiAsPmN5uGoTOOF1eFnETn8VpeeeyOnelt5B
hikteCcyj+0p08aeXwQQidqhPPPbbRrtKZtrky5mfoZ2QUReo0TCaw6sYN45NHC4tmx7AHbfrhdQ
+ChR7CG7L0CVnwmOaLfs0/wMLhBpK1IH22p95OJimPz8Zs+oP1TzDboVzQnQZnrdc6yhgfh4qk+a
el5O+TplyE4q6lUg+SEYeJVcSopSTOGMuJh2GIrhNNo1E3HDT/JSe8FIt6bXzphIRQNbWLSf5Jn/
E7VJ4dIhaTA0eVRNuWGaDOYMVQZbtkPPi6DJEV45BukixgQv8spmSDSqRjGy3bGZaFRE50HF+lQQ
IUrGIVK3KV1ZPgg+xS8xThtIKAMN4cXJgnpgtV+WKS1dhavpZjKTAqAZOfGF9zj/PrOQN/ZlR6L1
aFD3QW4Re5Ik/xBrcGFPh2H3illcqZV+QSlujuBnlJF62cIqZpda6K+aUdSDoAcwvUa/2uQEraWC
FBpDg3Ngi9DOvFpRVw3mOrVBfOw9+aJw6/rUEmrrVmDg+B2ZULB9MmqYw1P9M35AtfcfPdnscI4E
r2vAAqmdM69ioxkdsYKsqjiUqEcC7oPdXKg+WHIdDQlGvSLvyaldXKl7IeTx9tQ/wCQZOnFgfGq7
9Bl9GEVFCwgpUsoTogqqiPcQROHF1pln/x8piOrOEqjCPaU877sn1jkuUNil1Dis2k67E0KvWVEn
78G85Uql3KFtIyopeFTDZ8Zli2UpA5EBCBHSdqS4LIMzr0pdCCIcIozxzGtEpc/geh4C79kbGl0b
uBAAajOFyFPaKIh2lHWNelplT36Im8abNsZRk6jfdyMxt7V9KWG8Wvx91PHp3omDs49d8SH0nFOC
72MdWYYJVH88ayoTtma0vdnHuipC15dSGby/4vNYtwnqUCS7g9nRt9sx7YFsd5X3I6v3nfKH7vMm
12IOhF6YVwLtObCOnQO4JsNBeRQeex+kxyrGfFvTRvCPxa1mpo6Ht4H1rRFwStlC6KC7JSP0z7M7
k1Dnj3Me2tlQfeQ1NNUKq/4w5vkXLCz9TnL0STiuRqz+TzaodXVSG9ODm/4+gLU0l/NASdqoF0YG
hwGKzyf0GZ6+Ya8CAKKuNwndy9nQntGNVqaQ8Y0bGD8BE/3+SKXkoYB3c/fDXQbuT+n0MliIH9x7
s6jicOxVWSqgs+dEixNgftc5qEd791SP2UQGV0CNs2yv5JoatgRHo3A3SZ5foZdjXXX2hodW2tQW
kmW2uk6/CzZfWrwyHsYsa0EifjBL6erfV59WfrA8b96Y0KB9tCmMDieBmO1HNPqBhELyFuCvOKWo
EMqtSdG6+VT/ADpG2gsTC1FEC3W0KZI16735ldKYlwZNhHnHDwkfVt62Mi3spUA2a7HefGDHrzwO
Qh9kOxuWCvmtHWb3TcOVHWHjMC27+IJmuOYmQ79tmm9Uh2R/qhJKXoM7iHuhDEOt9NfNOPWBhDkF
GmXmSEvOjMR9ekilc0lDMJRdDSP8XibWVAHRZhGlvuwh85qqyOv79+Ha/qWO6f4GNU7PYUatGpTt
RTk36nAN7bsWNK3hM1QVgbee75i8RtxHsvZapk2KdK8xysypDKW+e9LNOvESEGHG0fVryEUNR1gm
zZ3VYJl3rwQwntU1U3uEOiTVrJ1xhbFPCGMLNN0zz0UbXDn+VZ7vTmcfoqhegCAOQo1k2HJIGA+M
z/qsXDad4RVTiEp5Sa1Qzc5KkAOx04NbVa4sgMx+xAsdO3UhbqHODKKrGivxKKmTlKnFlECg+itu
Moix9Z1vwbzAipQSTuU3huWiP8wORFPrgerJH8DXf/XWQDz6pA5oZUfQ9phFJEBPkg0zGQNi4TOk
yUGznyEOR/GXCEkWaZjfSRwK9+osV0qcEPOV3h962jK851lpnadMb9geOZpfZVHO0+A1d/t4xqiE
sPKCElCaejeAVCs02cD4wl1lZI3aW3hS0xd5GkLwLd3kxZE0ZiWqZ5ymr6nNhiikFUxfBLzS92JK
pOEEFY4xqx25t1IUpyx+t/9rIAvpMPrO4e9fM03FJa/63rhUm9Fpqh5Qg/gitYoI4TiBFls8ImDh
ulH76gClwZnPdAljVeEqSPRF00HMgmI6Pg3xkwz/TIf83dyK4ZR69Rh/O84kD+35PWKZ1jEtGJTC
wKKBB/0VcXIOaDjlrx/NhYdHghjGkS7fkHrr1zfqZ1XqOWz3TXNkU3/4LmMpX2RXmKXtZAduZbHE
uWj8+LY9i4FOogdn0zd4ov2UHIDHB+vyozwdFCdaXiC1rhOgTXh4RhFK7V48mNo0Gil3vTAawsQE
OQALLMaPlHu3YtYUiy9MsnoKKZ2gB0v4dIW2YecYrfgSJjws0jbh/PGIwzLgmgpkRnpP5vV1HZPc
Bd9DjyTdZTb7GS/mYSSXPO3vk4/HQC14gQWJT5SiiZPowSt8nIqpSuUEP4HlnHk59MQGZqKz16fp
ThrOk6laivAjAaaOufvcj3HmtWR/9o20qxr80g8bmSEs0OeO6brBBcHfpSBGGkJwQxUUdcFwk+Cs
91pdRimDPiziRB4wM7IYejsjF3FkHFn/QfE5dC4tpffSiN0oIoq3kMv01DhQRQP/6AobHm5qw/Fu
v19oIYybvLlVxOXviFVOIVILlJGQsW6XGgDah4ScJFv1ooMgCV9EEt1cxoK9JCSZLUQKpKbNOqwj
aQ9bLUvGYQA7GI2DkyXELJlkM0G41oQ1VlMyBDr8bC0KjkroI3T0Fg0twMPrbsb/bkck0XHAuIj2
Z12gqefrDcHXTyp7uwtA2dmXaE+l1Y2v4KRhYdMBb/uT0jfQnso+/jqh+uanlkSVBCiXSfeBDUTU
HaKze7qfeTALbdehTCCdM8JpCBnROYQ/c7YXR/VUts3HSTEw3+pRxgQLrmvEwKZhDVmbRGB1O7ZX
asYzV6ODG5E9Bqte3RmdtDUPPGaWKYAzA2YL+RvtCk51aaEtao9gUxl/YHaKz4dWeDGuzrKUPmYZ
KeFMWqTP0D/GU0wJMaqp4XLaFeG/r1uMC9EUHd2Y8LCuGvOMmPphJRA/q0MxD++OU+q0AADoLxbO
EMdoHHoeo1x4wnpKJcX3JRO6PI99pyXK96fOtR4RfZmzpwbf8PbQT9sgrxH2kqEUvuNdurSLyEbC
CtQWPrKrwCyB+q+VkWcgSnprgVAzPufnQIP8RFMNrn8VtnrUwsFOVZYmpNDE0/eZ+XCMwQVM9iZo
JqWzj/faegVn4wmXqK47vR5uxFyUHO1yL9UyyRItK00KAn3Fg5ZMrjRoJQcblTam5R8N4by7adv+
JKUuMh6LGDDicy8F24YkFBzNHDpMImsQ76v+jBIk6zBNzd8vsAGxdsHhWMd7+Wb0q8zTmRd8y2PJ
lHQdw8indOSrrIVdNvU9QzgvQDvTjxvygz5tPvxkXtAImPhdb9vXlOlOM0uij3RYcvOYrfxUBDOk
q1AMC3hA+Vv6UgcZ9QgS5svE/mufXZXDsFmFBuG+bFqBrVoboYl48HBipqoEHzVIioMHwWH/xw8+
Vosea1Jz8c6o6AN4x0ngNE6kd9tz41+LxFrK9UfBKJt3y6ofRsmuyATjUaLPNI+ETg2fINtyxBkZ
4YszUbuC1I6OGcPgVGWHDe8dL/DwdjGJ2p62Sh9EmHfT3kei5zMhxIHyEErSV6lpWj3yiU39Iv2M
kpGOZTpKuB1hHYGPZb88F6posi59Lgz2yXJLsRi3WWExjkfMDtB+EOx87Dx3yFn6JUDTk8SIT/OM
DGwifk3P8pc2rTU22LwbZi2tsBZARbBHCSbIbMsXRsMWlki9USpWl3DQXvzOzlwuT+/AxrSc1IiK
anq4WrNlhkI5T0V8WTjOavWbmsLGO7Jw4ygMeXr9OBISR92SS0MASFRFMKjRMPyOyTGIJqUGncx6
cSBFzdMDvW8KNoHsyZT1btfsw7/7ZfQCDu9WI+0QMcDY8ysQ4H91t109aUg1pTd1fyb1DpvJZzcU
xt5uSDAG6GoJOB0NSzTOuwU9QETVeA/WiWvFHiM9SgxkXL4P/Th7ziTDD1PAye1JiowNFYJ8w3lm
SeNvCH6LkMJIAUVmlYslChM4aOk2YzUywRBNNhIDq5s+e/pYwRBj5MFnxsjxTntgVzqTK7QB2A7L
wFPHqp14Fb+VS4WV1QwhKVek8vTEYuvAUcqGqP8o3i3dgTKZPGL0TvClHDoa1BdQU/dOb60EX/A6
oUhhICr/NQ8bkpTiAJToTi17zqlAD+KMg5utpXhePXbXD3Pov1npKRVHTFaIFZdYB6f4U6Xwcomi
SYdR6xy/WuU49vKMbbqc2nnFNKsXxL7HXDf8k3bwuWXAM4W/D4e/qUqmjvDSRbMdYItGg+N5L5aO
3vgMvJMeMjWduVbedHY3t9Ev7rqeGzyky10EdhgNHV8UZZsSmENh3HAbiaLxvB1KSYfz3JbqDq/b
hTkVaUvxWLU4lzor6EY7AbhVmPq1kHgI0r7khNV6K1jP6QT7EMFQpbaNIPV0eKXp/ljPyXplY8Ui
5m5KQ1MD+zB2jXppGCNVM7DDNJ623orpDILF+X+V1YEupzRzJLlvkecW7ThGyJGuDQi296v6x4c3
8GLVbU8wj8uVJwxMXDwVBPNeTUgrFZA7qk3b0fjILK8hPHaytZGPUu3bJxZLoRoS2Vd0+3mqWUUp
Mq00zFpDhO0PP14X8WSDCbCVR064jycpn0wGBKkOCWwm+LggLmXREqt0BWRJOKjizRCWZrtwz8sM
tUOjCLVtqn2pOMvXOQw9OHjnWsM6vDS39pA1AUJl1NoRdt/0ojgVyXAdCR1jpqxj7uFXsVrw0TOF
xFprmj9YApF92xfPfYpnwuyToJdV6yk8eBFJZKa9OK62I9IJ5X8PYNVDsUrWT9nUrcbY8ELKWzHM
Rw+NW2tPyM5twUF1j4LZP2IdxVrwL1G99ul2BDrPaD1UDLo2Y2PvVyEdbN+0Vj5yzJ43l31NKUPC
R5vqmr64IRSCfiQJrhV4FabqcpsXVD8/SIzJyw2BnQwUIeEJrT4U/ZSK5mT5akgnI9p3NdfW98H7
66A8SHze6jLU8Gg5TQ+0IfpONdG5yV1UxlvQFRUcSsmhzeHcpRDe97mLHolrXR9V5HSmtyyz8Z9G
+10xTXFBPGdwoQA9wkl1L7NpoemnS2iGPJgPMyaFEeFwlKE0ziY6MHkX5ap4zUL3q4wiYQoh98uB
G+v7LK6RY6I9kpQ7/q8VxryBB3SBI59MVjJixd0MO+Cg3R27N9p3E+o3niKj7zxI956ALoPBzVms
N2AOYX2BwTZg8PgMr40p6xUiDt4ugz2pJkHNg6q3r4I1Zv1YwQ86xIFA9fjbd0s2e+8ZhZPV5qTb
4+abO/WpsltvIbQ7+zalyosEkLY5Q9dduJKi4J1cVavHCipgU27yqpag4isk+Gpvh9zrgoQ5+B4K
F3o4YN1WSqrz454RN6f0Cdg/U9oZ3Sbv7MdOahPpSMuT3v23dMwfYNkp/5NH77c/eLv2fUPJv/+3
PJmfdO1OfuFo1rGvO26FeVnL+DgNkppeZECekl3HL7UyYjqmhA6Ve2PjNxPK261rK+k7ZuA58Tua
tq9gMxP8M6uZtHEM3gcEmzNkFnwv9Ljx8yf9tq3qNo0VGo8/7MGy2RgH7IPvdsaM93roZWW7/Kt1
uP7LG4DkrakzR5Lc9zAcPq/uK6n4HFeH/hLm7PeeOLAirW7dYAI2DBk5nKukq3Xy1Goj6E4aNjj9
qXD9wZyGXJXTDLbq8EtfP5aTh6yay1gewTVBzfxzCtensW9JG/xbh77qEN5Qk50ARRzktZ7D5inR
BOlvzk786X/ziaC5FthUXL4cweQuIHJr6zlxKLJJOdqCbX6hXEjhnlkdTXWPbWGVG8XxSjtyLsox
UtlZVB9LhkX5CYIl8cKQdBMCC61K0x2szlKJZSmMlVwgJ1MdzMhsqVrS6A4V7yBUEJjzAtV7qr1D
tbWVTja4MWF7giVou4meVHpFhOdNayG1uIWRFtCKCGvC7Zi5WtvYH/ValuB+QUWB19PdeVBF2sHA
xvIjHnk/760ipJJ4vEmBViAhcN4K9V2kT82LWS9E8X+nnMZUvwJyc8l/Oo1q+AO7LY6WcO6dMpfq
KSwakz1J2ccg4UQWml38j8b6wKR+MUH+8a1uW1vIM2m7VbLRa58+3gESXRA8Yul/+etIIim0bDk9
XFJzgNQT/McYIeukU2xcFei6KBXn9y97hLSalMTrpdv6VJYVod0ITZ00eO7ZzIVYVuCTUFzNYLbc
YdPRiMEtHcqqM+gKpt9Un/hj0yC8KuMA9U5GdZUNlV6dfQdXpNbc0HWV99NxDfFHq5VMhdF0PsDS
u9E5Qq6LKBWmVHl0VkoWKbTfnCwqNfbFl05yIGlzXQseLgpB9oLzONiymQceae3Bu9YAY77JwcBM
1UzLoan8ZJt8dcXS12rv33noF6KmcMaUzF1rnLzUi9/UhwNR0l5jqlYwtIlbREIXHu7lzzh/CIpM
qrAMEEqu9qxDPWmyS1XE/SZWBJT8hryhS7VwM/GldeihaEwor1GTzpxewVNU0VPgaWy2gCtNUo7Z
uzqmBqNE6u4Js+vPdtFrZUJ+tJIM0CEV4IfsjP6hhpmlVhDYeffs8WHfx0OhbUtgC9EZGBELde9C
Iw2SSBQ/RL5ZF+1KomaIes8XsrsjAQZYqb5c+WKDDsZnsSFjCoo/E6UvyJBecVHnyIlPu/j4AgOF
HO1z60rLjPywNRah2bxsfg9LH23PNgfLqfvDAgBiOdyJz2n9q1+ZOzzjG7bKubKEDHtVH6Y9gU7P
VvtG/pGFUbBH4fuEX7DPAr9yk5K+YNLA9ZMVnEaZg0kEoQimM6hMR/1QqsjdnLhm8IPApge1yam3
9PCHYGnRNNJRuVHGj1oZeO80O66BsFGOf6jgbCmxI+Jh38EXoOQSwmz+bSuHuuoN4jhK3K9eFKEf
+QwgoKzxVPNiXO2fQM4VLgeV74GMGXYJiGnk0ThAsGpW+7PjR5kUIounw4cDmpz3bsk6YtutqhCD
8fqy3iTma7xCVLBE68KiuKQTTPrKkpdlpzXHhIt0R7TFzoQcuzlcUaQuTKj6C4O0Hhfhv/d8900b
78ZHGzGYUIbIng0vqAFv1Emop7a6xT3Iosr0xGoQPQ0wn48LszotFRWbOs1+SbPVP6NeHba/lJ8w
7CGpkdBS2iMGZZyWYwof2ev4eOn9My+nm1n6Ji26+5x47rWbEJs6bsm+nvF/oSsCbmGBYzkGFuSy
WUz54JHKEyz6dr29zugbkiFLpElMmc8JU00bBIS0I45bcigiNNzgJKJ9V5T9T/fxQSHTCD4jqCUr
2jEa27JRgp9nXraUmI8tMMzMg+t0cefdqlJ48jnmxEoZBqNbNXb+d9U8QYdpWtOSduSXm1nefmpE
DwAWjUMlAwOAKodRh+Ivw6UR8pYwEwYEGECABRtyp/tPUDJ4x94QoLJli8rgYaXXgl+0wwpfkNpk
YvowL11149mTEAW6dhE7vCQNQj1/jcYmrHH69V4c3OYo5MLSkSixbBC8Q3pNh8XTxvL50XAqwoIY
Jl83ZdhjQ4ghpfH9KQOQbF5COVNx9a6fGa4BcK0Jtaz3fWC8/hXwHxY8ulcHZNMTWEpNgmW5dQYQ
KGanxigCNVVBHmsOLKjeVtApYCv4Ll7YVM618Frw7QiHm+tWpjtGCfZO0crnc+RRWlGIEd/jIbn+
LoK8iifFQ/DXdPC3Ax32k7lc+2KgklzZkJCOjSHguu0rJO/rCYRnEQ1YmxOhWAOyI+bgroX0nmdr
/ihqkyT1e4XBlDs7YE7I/AcpSMqrcyWrAZpVsK1ekDOKmObeHVgz6RuSypNiwvCjn8KQ1nix6pYA
c8eM99Jg+f3WTV8pTBVHHNHbe0H8sLBX7hG9CmIVjcQymBePCofhleUKPddjBeudPa42bqXlGCSb
K9lv/rh6LULzUocYcxutKYPnhY3wJ51QxgP9NXDxSBQDdurEG5Qc0KVuEmZfmK70JxFQfUMZ8ksQ
AcxR672MDBKtMXt5dV1l+gQxJO3l6qLlYtetX80/MuZWwhNqglsllCpuRAqBpD4+B078cfIJbNPd
HabiRMj/XkZoGrZOs3Mfmme9zAYsKOcXWjIlF4ac1tjHXPDifplNpeB6wo1QpKfDdFsZfPb0zCQS
5VujopxEZ1GYUfm5+UA9OEdYUECdz0RV+r2XlJMlStNstcrv/nDbudxn7uz8psaiA32cl7CHLo1H
7bZC+3FYyQsyZ3iQOwJ9T6ZXOe/rhqsQYa2X5O/pojOIXYzxEZ/YcXq3BYLcDrQ4qmQpdQ5+Fgf3
X7qB6LhNhmIdGKKmi69J+Hhqf6nfJ/BvjvUqFN9fj9xODV3Ytj2B76hC3bKy30IQwE6D/7SG77/Z
KxJLvioO/GLrJFgOzgv4xUY6Xa0SGCmafWn8NnOPZpTUjBdfu/Bf+/i6cvvMqKVgOqZryvGwayyL
dC1jmoL5G56FR5/vidBM9WQnQtfm/I82lbnggpQvFu83Z90Or07VunWVfaFQBhYJvIk1+7B98FPf
8FUUcT8Hk9Rhy/HnS75CTYZi558ju5UxdlTXeuxfodWg27mJzxjOtwlM6/hQDZ9se4Y/UI4tHJF9
U22cZlHjrswK1EplP1aO+Cakkq7Gd4yqR152Yg8C9TYEJy9WYafVHWu9ikRbkllA1JhyFMmFlVYu
YlStns5/MOVGPrtfvbxUf3AP45IrG14ecXz/IN+kdYY+kLubHgd7tJzUC+8/Kme6Y/KLB5B4+20c
nwjaVEzgAxt2GE6R4HyzpVAvIluOkOdo+GHUxnbvtfbTCxKIvRGRYEssQqP+mAOUQjxYq0htTol3
cEmvyjRUKfhzUdd5y6nW+rdZSwUnlUlVZRKW7hAh1Qf3aJaehS6F9cDKmDnyJOhR0SuWVw0ytyfk
7kLoNpWL4OxbGnzeEKhYV9sZVBA/kcjDJh3muxDv4EaQn+nwP7S5lPyUZbEmYa2VdMaK+iDkY0ty
e2IrbzX8qGMiivkfuFxe71dSFjRLYDAIdMpGT2ZeQ+H7BJYSjMAtOd92Zj/jKqT+KNPvr9rL9N6u
/Alf6p49LgEPHBiEITxqPyjei5CtyeFvLZ6n8JyLW/+cd5msgcpoDXh5UTjzwRbIOTrBrvfsm+HA
hbqO6xWS7gRgTx6NmETBRdzsDBC0VWwsxecRg6ay4bM7pjvl4emMHsqAepAO/SoAuNFU5aYsMLpj
b+80JA/Xw1Q/vUPwQjz1089EVFDhlTlswB0Yotvwq4FAEZwkVnM9AYD2SgfqA/baTeCsw/fjZnDP
eOsCb6cDE5lhp9TEo56/+0Q7SbT7L3WxeXjv/TzHWt2rGs3iYb9q07XBxMdrMUMIYUyrujixElPu
EdfzSaUa4l0GYIUH3r1JksgFNWlf1mj6dS9SB7Rbzka/JFKARQuOsOpHBNPTI1l+kgymoXJY3quK
aH29QGBqsaTcodZ9sd0llMnCyRXWHgExPmxjlvBzNnJU4d+crfLNn8m8zXEzMju/9RiconmJRKsy
poQhNI9pZGFDgQ/rkjWU79MLDWObXQQQArTAo5pQ5sOw2g7VTALe0ERFxdKmyCAq9YO4RnTHSqlL
Z+sw7/aeZHAi1eoGrSUW06uv42rqBs5IAOpEDyOn8qe7UOkvLyyfubp8+F3PdaQxUdtuFlPnT7Q4
NgJMvfyg3bfm3vOf5lLMou1isk/NjlHYWJmNa5LX/w6JuQIVzHx3Cvz+7vYaPyM+SifGJN9HynYl
/4G4lWHAw+81MuxYlMvqRif26icQlnVBTDqA5Re7GiBKirBOLQfBxUa9oyJMKSIUcCl9EM5Uq07f
ciPK+Y2jNnFw/gDHGpuR6kw1MsDAa36tolgp6viBgX7llU+pR2DmKDkZQUjIiku7ButQi4Ty31jo
NlWxadn59PekjyGIHla6d39MvBTHQM/hAg4SdvvjImZtXe8cUIO2ug3T3iaMGmbjxmWbYZ5gxj0O
Z6SCKYnsuzoXXOOETyMco1yZp/OJM6PjgRkVKW4VZfTzAr1MJVtA3MbkNP/01sYLzul+1k2HXgdF
r0iktG7rWQ/TRgTkPN1dD2dUYacQ1Z0d8/hVo7I9S+V9s/deRWa32uDwIGQ2PLNx/0zXoLHHfbh1
57z0LMhq09FjuvUkZs2Ke87zPn9l4l3RiZAT8lcQ86TX5JvKSRU36qBgDkoiptbNsnR9zpOs42PR
iJaZyzagF2MMHybDMd6BeIm0k21x9T2zKQ3IgIfHyjN1IzckinJ7yazTyQur9V5qUVojhnmGqK0W
ANm2Nh4gHdjRbEOwbfQTTMBzwfelVlHFzL2Nx659ZkvuiBeXsPhAoJDT1qiPBf4DIfmN/8ohYxlu
UYt9MTJ7c6EoyvqQc55vTfEdF4CMBMERnAuzQp/k/zRxe0x3uho9mjftU9l5y4ee9vw8yGg1mb8b
x/EFiMCBg0INSo+VnRVxyK7GLTKTGm6SdQaxj4uR8M9Bde83w16g74J58RVLUPIBxXQ8jLXSB+cZ
7U4flRrB98GYGBaBBNW1h6B13xBFWNjwgVmFeISpGPTCuJnnYmg8RDEw4cC2n3A6meTYaYCxtJw3
ddO2khKdt4kwj9LeHIr7yb029V5Z9pkj2IHdHm3jIbt0O1dAjucPzOlebBD7HDk72W1oztKdHkjy
7EYft5msrPadAwlc9f3AMzyz/6KZmybx3H41hbSUAw39hJejuWDLJo1m1wklUxui8sMIvkM8sW7/
tMX1FQtaHApHgtX1xQSRS8qO731OJdZN5XuXWD4hH/GckLQ4z6AKt1gAa2ZJ5RO8N/P4vV24qVeU
IZT7W/PvlDBZO1jf0emC98xVrzFujWyRSuZcHFJYFC6PuOCL6nyzUu9oJ2GO09ic3N+pAzeiXZVT
nPXFWvKy6z1Hleo0GE+27Moqb4TtEYgEOeQg/XoEUhfsP5vzDXoCW0Fl+FELFq7TOPtNu4ePwofe
XWjZj9lRKVze8+bj9j61rkiUv50lhIHNFWoQJfR4Fk23gMehfZZnk2clPggNKc/R9qFh/ChxjKwg
3UY84eT37mJmIWRmtx2wyY0uFEeMTj/qC7/OAt/M9Vg1mr11h7SoIVmeHCREoOwHMBPyL/1Yfec2
F07+xsHsgvdqDSVvdBuHwokxL88FViT6eFGLL1BApFvKOjrvGB1fvxY95PBP00irrJQCdM4081n0
sppPWhyVb9I95gQ7MUJ+2pZMHhv6NihyvTIqaOKWLr40SdJyv29ZDqD6WbxL/PGNtszziehBB1Mg
Jvg+Rh6PNT6yclgr2xBPzm/EFJ5nkMelXyrURbL9pFS8FGUbLkWevDZMdkxEr6P0zoiuj4u28wK2
40kVHWWQVjvH7E31VCpQsO9UH1tT/ezaWmT7S+WzPN4OVp3taE7ed4azLTpuNTJkz9tjDPiKnpVV
698jiVQU/FjcWXch9YWwFquwfSjuUzmMz3bCS14T7NF4Dn1A3bCB52SM7G4DEWUaEutdYM832v3u
AnfnzM7/utZAyIR4NpiBOV3qfyIle8jUe2V7l2zcykaEw8YdtE3MMrDFEegc3lIjS3t9oxb/OFBx
bA5dXfLbzo697HOjGIFhsNLu/X0lVaYI1w7F7CXKK7azLtoCcM9f+7StU+4ftRjrreJJu6rsCApR
jzOQWsFYgXi7QmJE5JppQQ3gXBalx88uqFpDPxdFcysBpjcJ4IIEZxlOLeQYKIbJ+3XKMw2j1zgr
/pdwZXsux0D+nGf1WKvlBiEwPLvsqQnjVh/LLejaCShzyXyqIQ8ecpQk6E6h+50JYogTg8dxRpH4
1/4iyC9ax84944oC3HakOrkeEOUt0HUd0F+GjiQ9IhAnbnFjM6YXxg4SbyP7VwdQic9m8oFAoGvZ
p2PAeLPZa2qviscr3AlcldjoTb2lvyCR/HMCJHxuKz3JaU7FtMEPxdwRrweOYWo6cwJo/nf/o2LI
52l94Q090X/IDNUC3cFs8X+HKK8m2rIY3GnDKXJpkcITshnOjDrknwb9z7Gr6eGUsG5lbK/ngEld
IdiqDgGR9cFinLIrT/xhx8cAP3iBlDrBJf+K78X5NYQ7acsnlThwOziY1hkFAlewQG5FP9uHwXd6
C4Q48BLlY67gLEg1efYlo2uWmmKCL0Y0+AzZ8GYUSVxulV/NpqeiWg1ATFMvoFZ+az7yHOG/CT+3
z5yG9mY7h9GtqXQrJwhMPc2DZ4ZVeDsqY5MyxSlmKtsAi6UfK2Qx2KlhiK0IsLIz6WuqFmX92alE
qjPrmVxa/zoAyHakAQSE+s3zsA4vwYag/MTxkD+pjxg/djHVj+f/oeizUpruPxn1vsx2kzViS1eG
KJVYBQFHE6ddlNEzwYBrgh4cZAc86ZrGdQdKB9drL1xokx5CNSuwdZF25QxOjCYV+iZRy4rdL1MP
NH07kklgMRVNUBDGUqssTpTpvurizz5u5X9tYjArtmcgt8r26jtlK4MG/re6UZQhQW24mRRlE/OY
u2tly8DrWY4EZL/BH6gb2vsCJ3w7agD/zmgwEhUV7UeNjKI807uKFXBsz+62gh3jopbqjkepvItZ
c3eQqwSzfL2hXSqOiYdNoIFvaN7dM1kOiDIN8Xw7+Xo37pmzxkppdAP4DJt2JOpI9ooXdi8DqtVQ
NrssaSviO7489TCx7HLzdebUE6bNqAnp9UBEYijAUrKndHSwcENSzyqqfz75+uE8cRJNNXj53I/T
2r3BnYPla32Ft84T/Tjl44FjhLaPS3FHLy9V64ciLAwboVf1BwC6IKjoxaQgbd6LvA3eivfM7OM+
lXD7gI8JGrjJhm6kYQNjfYp1rsB2eljSQqRMjXr90+d92X7JkSpeiW/7o5rdekbNdRW6lxxCm31F
ix6DUmz7YFAXZfCMffdMzfX5LJ/8AIBacgnf4bkAYbwxGlt6obTjS/cDaA2r3qi+/vgynzRbzT76
e0Hjn8JSWef7BK9HFrvhX4EsAsp3mzEunVpbEQ9IwzmNQzVljQGGHbm06qK4z5sVzYWykWqmOWhE
6d+f7sWYxF0/qTxJw8C2TE4IDYwLxydySV9AdBJoYC/uvvjbOhchDpA/MjgZ/0oEASBML5F7PwCV
JB4uPb6yrsP+wDSPj8VyIgIO3JM7l6ztSpSi4mzlyUuxN12V95AD2LQYSsFui7fywy+1hGViwLL5
XYfJ+/6dOdeFL3Dpe+pUeYaDPEqLdz9elaE7qsegqRbvmxetxWwOJIkzlJenVV3ds6gAB/V5ojt4
BtQYucr7VVNIyrWg20lJXFQre3utqSqTs/DMoak0EKhyrmoQ5V2MnJ5paXbyBlsqpNYpV2n4BmHP
py9S47TW9yEnI5I5GH2yy6Spr0BLxiDjP5wSHvYlzOWwapuHlQyHnxfeyQhiWUcBl1uYOnqZPQGv
jJN3jBOF5ckNQybJC1H6MyBqBBeAC+k8JQ2CeCW8YCGQ8aWPSYEr1+0Fnb4FUeKhICBazjo6QF3l
GkeM/8kOH7YKDlb1cGYcLtVCWIdg20tixWpHn4RhthKZwTuVaDfYSQUtiKLuzEzuGysefsp5s8wc
UqalPI4PkPk0LM6KPuz7WPdNNKq6zYy0Pr7MjF8IjeaaC5O8Y+OhNYqOp13/bEbP7/dDpsHgSgsl
CoSo54GN1lqOLrnR7DTjNnLjf1V7PsKr+A+v76jm2LzMlW0Opi+yFFfUGJ7MjY4kiU12jDazXa+j
L+vLw6oV9Ewu5y+rvugbOkz+mEqKw+F2OpO3TOrEX9Ciplq05ThZZ/pXC19lIokuzvQYrMBwdUup
9akYZNfsJFh3k8SYsNYjN3kZAeqc7mJO6i2m2oCHxpQUix649zkJN9w21amEtd/Dg7DDa3GhdoVe
m/Qinl7vAdsqkJ36ANZYVoq+ckQqlcn4hSYzqEM860DQIQxUtZtO03nsH6L5yNPxXLiagsmjXUGi
LznsmR+DDOFSTPCJzdChrTmywEBfZAlBLp1FCW3FhfDhZPLSiwou+lE7M5tlRot0srhpqY0j1v90
cl0ag79gzCXveEk4m3aGIhHjzk+OXASW1fG534tatXUhRyEPlyLFZ+3WBCFizOJ7t8n2GnqWk360
8RHjPOyxtZc2gJZaM4J/I5SBxku8medWLZ/s6cELSS+QfGvXV8e0/khUXe6gtlBM9pHuyod59UkV
UQFzIn/t8LbNLVWIbZomUhggUE3hMMrL01HtEUWblHV/5WJwgwvDwK4Xrrm5CTLwtQz7W6dsf4tv
16wGvla5lukJJ+nF1B9hSWs7IvePvXZ+sPMnnzw90HSiBfsuxFTFeQyHJ45ct9Ns3rGI+LvKIwsg
g9lR6hdNuL+UIbIQx0+uH7oAL1Gvy7bRixZELKV0M5toVip82Eplnk/LQpU6kTWqAu5brQFInmWm
oTFfEGUCDDkOrL2uOzLfBq+YnTqXodR0cTgq1NCXjMdiLjO2T0UnVosfZacTil419S0mUr+3orQx
0pcvzVt85EQBydEjfOECKNTfCFdblDhByljqfPWPaFUB0qO3HiqmHfVAHpNSDWlET9+nYwUdq0yB
a8RWTCNx+xwnO2tYTyrI+BJGlJRdbRZccyv2o3vNJTTFCzjdAu2O0B8dyAEtaN8FA/feXYuR2tFa
E2SLRta4JEoNXHmSi4FlMkC1huwaw19LBXkpAH93RYHXJFpZVGHrcxY4kZPxpLB19EOQSo82KSI8
G/5Up3EnE5Gw6ypZLCvNIRAsQrtKBT3rjCdjR3qm2CnY+eva2KpNLNGsOLDds/KCfmssCWnUg6Cx
mDY9U6LOzDdyYQZgWDZxjLjwxpfmZjjjLxaJ9hX1gKAygis499NCzJFZMJCMv6ghowSHC+7GeQsi
EApDnNsHnIU1NMhpiU7ZXnIKq7IrLDXM5OwPdfv/NjtbYgOBwRfW0xIP+H5GhWYqO1dYk+9O5L8i
wm8nSBTvO80lnuMF2/LgfplxjuT6b9CHk0MrH8Oeskm15lW6EmQloHW/qW58C6caDOGQe26MEbTk
tFfbiq21rh3aKBXrXmHCKDTpNAWiQMF4KRgOXC2/a376sMWXW4WPj/dknB1U0JOV8btPF6mpk7k0
A7yzja3M0u9SlRRTB2ujaXVhDTWDkyAI41lD1ourvs6/xh+dHGzY7F1uhDR/XXZkKQOhOFAXcm2Y
54XHqqHYbQqpgevHTMh7dv/xLtnaW9/SDCG8OfmoupdMZhQdy0YLzLue/VbQFENmPcaBMJISpW6O
ZSO0FbCeEfslUBwbl1DgRpf0dDfcJe8snw0fw9qe4hb4Zqbxd3OFIzwITGzv48atsuYp/6jqIHA4
nX5fMriwxlOQ4GbsEeoXZEkndJoltXnJO8VsKJQWYaEgEBlzboMAhzeFmhiFBqSXkyHhzHve0Wsv
snsKeEIS9UcH2ZNgsP4b8zEOEj/t3mRE3y9TA2BT2JeKvYOybyk40gyY7/NLqBdjoZQeIbxPvQrB
vfDQIkmzcvnGwYnSqnfs7cd6Wa9BrceiNZOAsvi2N6XQX0/KVAf27ffswV61Q/VTXvKF5qev5YlM
W4o7vdNzr+wGfmhMOsYsF2e8QJABFWZ15S5pcQXg1KPUH/haamXbsYO9Lb1KidoTuu3ef64QbxX3
fKUP7vC48uoIB2HBSW3OE3Bcf2frl0MiJS0ggAft6U40oX+0WOtta1YiqQVtsd7TWPdT8s7F2UyW
Idb1mQLY8nMkixDKbgq07mZ9bdOGJzTv0XvJtoxbZTSCXwO0i5ITaMY/MZM/c6dU5cD2Fwq+ODaj
RebnURy9Lr1OAJv7PhXUjVDi0PKnGRsAos7IQp4/TA0zMllBoTYO76wBtsLhVNM3GWFHeTbpqkda
2vYLzWJee8liEwFXv9He/68TahwQasxOC9VV9NzKalL5iEpH9qRcla6T5+/81RVeeGi8vbGHPQig
LXBG6qPT1yKQF9Dh6sxp41hA79XeWzcq9GGtoVmRcG6xIaDzQLf06sCWUces/D17ySYjF4/Kw8HF
1nSHYv9hBz+2wtMEbaI15fVeYm+jGatlJGqR8umPas8X8Sp0TSmz7rp0N9hOGOGxI6aNJLRx8fIi
sCAQ83H0PbgjR+KPIcBky9ZzDwGM8dRk03AwMtHuF1a3IxWUx2X+edS/dcPQL9vrz27L/kO/TwTQ
PGjog5dX1wcnS83KusyLPe3f01G+O1TJq0dPvqRUFCxUu7YtD6S179RUcg2QUIXO3XvB1ejSgsQe
lQvdSOIxi1iAESNfRTeu5cdvI9W7NrFq6kqKo7+HVngcTIGizIq1XNczVQEx4/E3ty1mQhIy8vDr
hak2hAzxlpKBtMZJGoQQnVlJLv6PuH6HHY8OOckKhmq73iIvVfp4DzXTXLzKW8/dy18F1ZvetOBQ
0fSsJjxCO9+K4vYVfSjTBfI/O2opRsLV4CnBn8DkqEJlbc9HkFvNpSQvx+hYj1m39RLv9DdPXplV
U2cMvc6jsdKeJNNrVO7dnd6YwyGWZr3yjHcoduxVtObLzGuvZ0yYRd3w63NXAp5O5ENu70kCc0fO
KQda+v89wijxu0dqw5EKLH+LxWTCIxD78Ueoehv1CK4EKkLB9IjLZfyXE0I30iOvcdPWRug0ajlf
GIa2W3UNVjWDzJDaBZYjgDXVpSumuePg61KH2N6fMnXl5lSkIoUOCcEwCmbab4kH3Nj1Tf1J3uBh
MM11tP6tg8UHg19+Stq/LyBe6014gKJyRRHC5lzU90bMqPez5w2WoGif2z7wW+c2zOddsmes2K2T
HeAFl0NIwYXbw2mSvhcqUiHkW3DIPIzMnlSxqZGZZyCR4nn3tHzcihchRxlLx90+5cstH4zYOWRi
lEu1eRLp6XsjhuZGCW+rvUOe5NCYhNei+ttIaK0v6lHpGAdtyv8aKk1AkkycZdArEfYIX6N+Vf1K
aMsFdwZ6CP3Nsaf/m7b8kNhlYYd6XxzQO8REageQeiAc4kPi+BsgDbnJBzEor7XV7r8xogDEcjIl
V3nkbyTzcU4q3cn5Er1dwXoMO5a2mNzJ4LNM9Yq84bduTpbrHgnA9/Z/Gu9xqjFtd+sAwxZX72za
EAQMlYi+/Z+nn6N0EkjFhFKhT64OpFuLs+QiGv0by8Gu0oN7H7uIhfGS2938w1g0fX0WvYPqFT2I
ah2FLENDE0xJlhc/Epsu+3Wdq4jokfco2WFJyYGHPpPHL3dupVCmO/u1prJf8g0QajHTxCusJgAa
jQKw47AguNGHCFjpVhqbQk1co3DCH4/zEh3hchM9aX7spzMi7NFFBOFEwJVwiAsXWoP0LhT8iUO4
5Jej0eLVRMIo2OAUivfJ9cUGpocZ8TZF4u9yXXXzA/LylOLcT76NFIwILmYWrtL8fUsqgfhy62bA
0rt0INe1l2RrKtQnC3FVgEgwlQ3n5XiQOrg1NqPVPpeSqkIPhbHP6c3Su0fABcHgkkXBiOAlXPpx
rWFLFeBHrpCEiijOtEoQCNs+3TdolmWZGXHZGGcPCxHLcpuaaQsr2Sd4asG7SOnDVSVXobq4m17d
WfSmeCA5b4C40wDV02lWjYMSaj335+FvA7FiZmqBjPJ++q7Zgc0u6pWJNGVC9oXmI5LctYnwPm46
c5n+PKhF8nOO0X24aAM+jLWbHO+lQNwo7F+5pIlqy5ZQ6weNTQ32emdWaaKwGTKUVLM1DHEVN1A4
f48AKVbqPAu4hdeEDXmYRvOqWoGeEBRl4ExbvG/P9eHPpQBs7cH/5Ooek/ncWcrW7ucu84LF/rRP
GUCKgozzAI4onoK7Qw2K6o3VvW/fufsFdnDT53b05KvuTW2brdheozQRchTY8oaLIRYs6jmOgJNO
3vGgUIiVNocaw4T4csBXYAMFcenPxm5EdDmQEu7Dva58TIS9KiRKIsIItFvvUA+qPiofl+isriaL
YuIIMuZDX8Pg9wTfMM0AztdTMWubQu7Zi/xrcj2vQbGSuxvzBU0xjliSbOLMsvKvGU7Wk0/JKXlA
4yO3vz3nT7l/35IlBPoEcDlHLEANE542GtYbvu4k5h35zHOsnTaSoKW52l+iSaplJxj1uYwOaIOD
+WYG+inhKPjQUUAeD7HBE/OePYhUGOQ1AhssGA/ee0kBpMFp6Su+H2IYNQOtm9damALBuxt7xBEW
0RmzDbiv+vVvtqmMaKJ0oIYQhc1oTkD0GzeJYwZrXEnZg2a+bGkjDWbxczgUfgP1RN+/CvGeDmUQ
8tFRUkLxBYgL2UQn10ikfV+R0vi2oHKgjKmwPgDraiEB/AU0sF10CWFK/kLwUCAznKQCRuglnpj5
G9TDIB1ElBb1wTL+hOaGXONAKzu2IK2iFHi0zVlpm1GPJ+lk4rFv0NhFx5nXHHskZttYeq0z38wq
u2Ru1WMMHF02+CLNUIyc0tpIjGosPMfgSMukl8sjSvAwsH2x24kDsfYCrBX3uv8kdUZ4lpIa7Brx
DuS9hBrw8h3BPlgwAF8KvlBbwcIaUj2JSipiPXFx0irv35QJ91zF1uscpS+m6q+M44DE537cNwwk
/URmQTVogwxWQVUfjoov47ixCGob+PoBGbYC6PJHiSN2ox7NHiiiNl+m5CCVE4z9PhGES/kWbAkL
54MhyU117qARojwax1RW4r6qel/k5Y2zYbKU8NfawiFsoFsirTaa8AlVv2S/Am3tm5tdL+k4jOWG
nRkrSzNDVXBFu40dfUUugPEBSOJ7LaGIlFgziONFiE/kfxkLHVXMMtoN0HULy1WsvPnpQ9gqh5Tb
cGFMKhu9ZkphWaTonYuXDY9DA+TqGnkGxn7v4U8OxBQeExtHfy/m6xYZ6FljNTctc3I3xtvM6RGr
qYBl3qaIRjYv86nPQcZtWnRhThVVqs2LzACmSf5yUuewQfN1R6rcQo98kfI8GjeXeT0YahLvWbhf
5v+IlFoDo8CTlEaGZA4NmoMKPK+BXwXsOYqWFtKz3bZKoj4vYv+Yh0VOw9WPzmMHiPn4IGNpMbb2
FLNiGRL6f+NHbdRurxDrZJGKCMt4OnoMM3eaZoCX3ph1RfI/ie0xMX4ar38AYiScYL7CyWAiA7QU
sIR/bhpK+YbveEOd3aw3dgDKWs+plJKi9OpgHF2ZcQtlHKaLVHksbgQ7Fjni41SyEa45QtxuRV+E
9l0Wwp83/kXrafrlloy3EtHF0ChXzqMny02itM9iWcu6swA+Q45evZGGCh1FxDquIcscnNL30VH8
EW3eVpPKwq8Ou4f5fFD1eHvXTPIxyKJ763aR/r9vR3aKNTgk3qggODHheBf12mBKVO/N9cWHjBUs
LCWQx+uxhgGPwW0+cewp2fkHpUkz4YeL5EX2YBo9b4ZDkupd0763j+yKpOnIxpP7h+/wC2xmO1/W
zf82CZLz1ddrUb0gPWRSWp9d3gH0JohcXOin3aDh/0EizmDdnihY8tI9T7tOq0QD8rRbPO1bZfK8
uSQKoDbWYCJHaPLTZZOeccCHAzdkjBpueSJst1LpIk2Y7fuQc/SAPHMQUyF+LA1g9DHuq8reRwcR
5DTYIN2lJhP7lSqfO93p8Q+ISnpgwO0v+9mG0Wsbcl8bKXL0KubZmU4z+c4R3lcOn5Q5nPru8PgW
TxmG8muKrif+T0b9Za8f/XAJNT3DI0ESQKreOrh3fIgeta6JSHhSIYd2Z99CBH10NSvFBxbWbJ7n
6TAN1HZS5LWrHmQKEWCjp11Qf/X9SY7g/o4iTVS2ZBR/eA1JQcaKc35mBk+2IKxMFHMVu6CZld23
XWK7A0SvNqjlY3xxRIzWMZcJH+SYSn0C6VaRABDYDO3BgaQ0VnA8yI0ouEEkADnJ+iOGxWBpeKX3
9KM2aAXLAvj60vR++JP1QkwychRwBVeHgeNxbhbmN7RlC1awMK21sK5iNxe+YUyd3Q0B/AGgU/fM
LklJOqPrVbNVtVuksIDTQK0rL4OnpxNjnZqc44PkP81APaJbWx9kBo67PeHibC7vgBb684uG0i35
BV+hANbEaYVSFeVBHL4I4XXvlRG6DBtZiVGPdWSlQ84ZPLAeFIZswCLMKw0Dg4BZpKVU2BQn49gj
3EqIpTp1K+Ilrnw6HsXiF3e18rXveVZU+gefJtIXn4czPbieCgnN6rlSPmjU850JL7xrIoctq0X3
TaTalEGQz8URkNnY/Rt3vsOEtKTv2VcH9tT+85kfZUndYGSb7T7v8j0njia+8+ifaMn91ygm/i7L
txxDqagoPPZbBFhr3dT6Wlz7vPfKyTUWsv91dGVkonpXSXGMNjUAbYcAeh1e7Ywt69hz042cF1dt
mouwnMc4IAHZUbAQpFzzW5jg9SXWsaCxORjfGrlVmsFoIjKJuKYCY3qRSIs2SqfevblsPCAGQz6l
IVCx0ZszPocqArNx7PbFLT1FjhsweSqYCyXB4SENRqRAp1Noik1STeqn2WekDIvRwCKsLA80+WHn
4dntt9Ir0ZGLV2Wvtw/E9Md4mx7VdTBfZdvevEpuQNrq/C2YO6THtaR9DBVtdVEQOs6/xk0UC2bv
Q7foFsCGixRxtBFw0XTMLCi2n0/0eOjey5XTDovh+f3CX2lXPHhSgv7muE7y7T8euM4AKGSLXHrd
MMevGd7GsX01MpInvA02Oog1z0lxkls6vM0u/VPjxeUiDfnItN7/YNpd/2RpzSoa9+6gxbF8w5hW
hZifu2BUxe6c0KugAsQ8ihw2JhgQmjfMt5ndqulYeC9ZDTdfM/Z8UwpH/nr8R9VpXG/qLAQE7Ln/
2rzLizkRa7EgqOw8hKDTaJaaTXQEJWIkIYU5UFiO0oZef+Zm2aho7uKU0odOmRf11y15aJ08gjK8
2dLUK6BhLeOgVrhZiEHA0HubbTg5AXYr7Pi0AZWXeBt6fqBMGk1OhUH+lp2EY1qVWWTgNhOQpBPR
Cz0wD2ZncffDZ0zcaQY2P9zrJBVg4/d5SqBIu+ZzOJtIobWsZLkCGcexBI3Kq7sSfwVV/oWTHRYw
vXBSqcq2ozcd8/BtkgawgHiMDm4+vAgCJxNYCzP9g0maPdMzWLiAERI+g1R6mjR2qFeU7w1oelux
8jEHGrS/q96uQULUA9B9Z5JrLR0+cB74OOyaiqoZQjTRCBUrCXN5HIbLHujsAPyp25Oe/ufX5idA
2g+h7/PZBXBnB4O8+nenW4lKnk8y10HrQbt9utzRkFblSt+g462rk5Qof8mAMToW6kqISrOOBQSY
RI/hCdTsieGBLEeUVGU6dik9zmbRG/Ujpfx0UzVmlC+eVCnFMuXX9qRP8i7itLoKPAMwzH8emwYc
sNLwHmsdy6GF6PV7MwyUEPr+NE8RazgLfSlz9KH92qQKlj/kXq9hKTl+PLSrYoe2QxhBjx7Tro27
KDikv2M6Hw38LoKv9GJQDoCQeWOyORxzzdDaXFHSwBzxysSv5MGvi7CNTyyRfaAYzElAV8SSQkUp
qGy58tT9sCHD+sQZNWI4X/HheVN4NR/xvtt29O6ACKKT7TrgzWhpQmUWWCwOmT/oXuC/lefTvZ8k
bChxS9+xLGadkiOsW5XwU2AVy0Kqz0IAqED+p91fPa9OwUBIXACDVQ9a1x2iOGgFjJCLVWUQLK09
CQHCT2Bl1gpxcaa1nLaxe7ahd43z29OFvDegRIV+/3SqO4jFc4yV/IazTbmt37q+k6Dts9R4yQgD
QTrC/niO/lDuA5dD/mIqBb1KVkvecX018kUDt5h3k9DlCcvGMsrfYimeKBvgmCpRMSdx3rDxvitQ
UE6KtEgrOcXeZtjskV5bsUdWjpPBd14Qe0FBq8o8yHFcv7xVWTeDwScJaahjGdJKOvfdcQNP0Aou
JSXWxYrImV7M3fjDNf9lfNw+5FWpG/754uBOXaqtw6tOLFXwrT+jgRIbbR8paDD/OOBuvcVrv7oW
XtMdviMMNOlSSdhf/WXTQ4RdAz2xHHnKTezC4aNN5bT+C2fDSJL36qsOWqwIRHwNm2ZZvroyNG3s
MULJ/YOspdXs3eEPjmc9J8zamIVUn3I2+4U1p4PFd0crgaycW9PKIsaFC15K0Vb3H07+h5F77HyQ
NCH56E/nzEF534oZSWX1oWdq1ICvhW+M6B4HMCkoo4vkrjYQYiVXWro8JzLGp2t1b85IhijTpXeh
Wjw2douhzmjbkyVLNPYoDoE8sUXZrFrVBGMrGn2MKcpZCbhVURt6Yp2vndRMfd+F9DKu2x2a5AY+
m1i5hPowEJak2Yd00vJ4SnjYtI3pQgWC6vujLMkf1HjuuRjgscBmsjfaldkerOT4TDJq6Sex/A92
5No/MTeHwOzU6cneaSuU5XOTDK043H01dOlS/ITNOlKwlbQqUp32OYa64mUP+Un1S8Xfg/UzjNh0
iJBgZqtpN/VUFZLgPLpGTCHsucaIbAamzrE4Ic2BXibU3yMPq0kYEA4IQaDRW0JQ94aAwze3pPyW
klAJLq9AnkS/ky+TWVm4dP/IVciu80pl+WIbAaV4daEdYf7XizZ3DnKqjWG+HQtm6akNMzM05qGP
fvIhSGa0a8gY2SPIZv52dgK/MvnC1BGwUKYlpkgmpvK5893n7WrT23tTuW29VNyI0gOzax7RcW8O
M7XmgJWcqigSDQqyV0wkmx4rqMv5TQjr3qTi6aODckHqb5yIL/iEh1Y5KnFYOaGF96VT64Hermvc
nveUOcTTFE4ztVCB0ej+bFppfX1WAyNYEazFkC0eNjw0bqMK18qQ7xuahI4GdNjSmupdZYzy6ai/
w6/y0LXWcBLHe6HPfdvTKB/ZrD8KCddtMq7lpTe1k5rhVkoDM/d1RVyaLT05vN/buNXUuNIIlwrQ
iAgaPp6EjKlUKIbuaNik5PYOTiz6C6X34DYJPNUD1YgaO5Qpuqa6sgWIB2dwPteQsDhq0ibo8uvB
+RP/bD8N3ZzNH5qPF83sW321ibH/04e+uo42XV7cuW3s0Rzp7mEtJ5a7sSUG7JscnhHDCzVgOHUz
OcufMmV4FaDNc2a2eqVgPcB7W+WRWayimPK9Gc1igeTQkaK3DcSqjmmGN8AwWW8spvY4LSjRcsq3
v4X+qNjIqLYAIAe/v6+TcrYBn4zSVK+coXctdERjO9RWKR5mZa7GdMSNMB+PvLU/YNLxQAZt3VJ8
eIVhOUznr4bqHgcsDroTZtCG30W6FajoRFWGmCDvwS/nFP2wo5RRbsg6mQ5OaFAmR7E/EsilqMG9
B7wBmjUreO/AKvvGjItwez6eTg86L0zEIaFZGXsWy1f1f8aa3NH5+uelSo6qBhukzV9cUsRlDKHw
44ozYZhfqXyXJ3NSUWQUXsyYvtG5QuyTeGIe1Vx40OnxjJvHNAuS4pc8zZLkwYBECz2jO9VaUGXx
bkDI8zM31tul40rt41cpXJ4GLwOqb48BM1dQz61OjFXU0KobumBLubqnBOG7J9vBR7yiDuU3YGZu
2D38zJFlilYG48pyExLlJ/DlLDuBPp4Gu4czgyY6SLWXKyAH/ysQintt6w44CDKRRLCPRq77hXz0
pIFN0OR2pd4j9y5PHp3E7BFJQ42jfPHdPbH5/6kbmlnBb/x25Y108Vrd4/IwpTptDjtZ0g7mJFHL
q2x2hZFwWq6q4KvO13rRjnYrJdxwUmxV7LZE+dy1hfIjqzJyULhPJRooVnaW16DhvidbOLsIaEfP
bSZT4IARQvB9NI5VpsaNM0zPA3oFE8R6jlTIICHEGnRFm2/TkWIO0HEuiXuQE8NhQdnZPNrqir1d
Gm1lNc/r1b3ce+4xvEc8MmZ3smhMv7mu9r5o0HCWoCO//1HMMaVdb1SVxA/R/stIOSluIe+UAKDL
ZeCcACYjh2wFivMOkv8v3E+VhRNuOvKFbm2bgzVXHIsGMWVwzRXe+JxYJlECb6B7dchqwTFpoWus
AkhRskh9TP609R8VF9N1YUOyWP1WUNPOmeCNnQrSKrLsANY4sQbdQSOmJTB7TbGmJFqpC/tSMFqG
hSS2Z3CygPfGKQYrRZwZYUiQPqW8rPXcfFfYjd24plcMfWCCeJLhqvwmakeMSf9w6dNcpSmwyxq4
mQLo0pSOAEdNx8RJ7t0QqrPf4+hpEsT1w2tRqSRhbfPjxLDRn0MKrHKih4hHIzFzsw2XrfZV0hSa
WcI/FhJJDxxAbY92QE5DL9XZSwQg+ZaZ9QyZL2Z2X85VMbytwS1zbnxCdv3HRfxXgi+uE3eAk4Qv
UEhBc0KHQ0WBayCYwGP6WS/U04ZFICmZfiOwfpPbGtJfZ1gy++s/9G1nitpGFQQSHVBTnPSmOwNn
ZE3i2YALJMDiZBGHMu0uL3s0+h2BR94hwS4SHYvQLPYcpnotY1QKhFskDC34a502eTEtoH1VB+mt
l5pSXXn/z6ksVN5/z5ISYvjIk6EP0GvdgcXS7wu5Dkr51PdrKOj2Tmd8tNZ0sBr2AHe1MJmSV1Y6
fJ8iGZCec/RWBYEghtFAu9910sKhIAnoB29DV1foVDqCAGTa0iRom2P1GumkZeHPlz7P1cAvkO1H
XHJfyVK6dwxOG6IdRQvTcOJKf09YRx+zuOR+Hcdipqt33DYYAfTZoD9CzIbiyKkZRBSrQ+Uy1gvS
z7DlbxbVX09/qGc3Zjt5/2eglvvXLFTv9ruAMGdpyp7LAp16HW9T1GOw1j791Dj5Zfy+u7giOuKK
KEqPQ9i5oYKvX+LrIfLCsXXyNeF3iXidnff6GM3oO6CnaZEGiHT/S+Tz81//aK8XEOgQnYPaW8yO
Y0vy7ehFi377R97AtIFRX5Fu2IJnp05EszUiracsQNL9lklQ6V+h3DGvXxdE5Np78di6Ioh1BKG1
oBNW9kAec4nFhUt0Uwod8iAUJx6jRNTtMPDBpzNPULtZpn4kse5k/0PwVEG8bqekC8l9WJWyLhmn
V/dRZfwk9BQZ10gu34A9Yp71bvcIgaKmtmC1BkzkPxQI7NEmOPL3xr0jkog6Tv2l4Xm7bSlyWF0e
G+cHu9LoP8sAcVDAN1Nnf9FSvjiuC3S9VUbb333NjAiXjQcIhVuWlm6BnaJLfQ6bZ3mlX27DwYGW
J1xJjP+uYblcF+3RoNoADtShEPh1V1G65scYp4wJXHMu25LTxukKUj/CixOPQsxF9tV5pddIM6zs
Ytw2pSCvwLq6Qut7wi97NybgJHXT//Izs+DiOg9q82Ri0Jb0aU22Tz9DXL6G5xcC9la4k+LbC9Fw
nJMF208kOzbkHfRBbPOm3PPelxhn5wZyl8kn/iGh3vlNCDDo43hioeWD/gFiTecRpQiHDaWLJoPC
fS0Gf4DY0R/REUedULrPo/Nhx5bHmZEggwqvxqyDuKr01pTrGXH+SA5ip/hXmtQntXyA5c0vhL+b
ra6n3Ez45Eq9RKfLCEiDUhy/TblE8M16iaGFxA5odHQnwnCKXwUbD1QgA/wiTcbfF7xp2IlNLT/o
O+TZyEcja7mEgmTw7bAWkLcWUlb8ptX2JIxMF5Un0pyOm/S/C2VGi9mO6aYmMvbQW0JJsIo55j3M
iE0gJ21uN5Hln08DQ30K3u3M5z3LT0itnuNRPMpUlcImkNL7g4Xks2eDVwxITf6KHuJDfEQIaqFj
uDSkouvQnjTSPFwMP6EiKeNHedT5eTnzEfTJRTqCyVjSCSNLGxkue2NwC+zmP4PXHrCARywyLG1N
sSiSOqhpPVBwi/TjQJcO2JIG4GX3eVVH+6D8iOX07XeRoGPoOrzbEE0ptfsBdEMFoXGq9PRBonwr
syPhZzubeJbt9Gfqhp2Qm2a40qytbSYL2kvJwLK8sAhKnlfoxwNgVnqOFeU9PXnxTHYN7URTGeYA
hWOUpLeT5Ml+zeI2AIylhNrBe3HjkvK3hcF2PnsjFB3pe0ljKs8VDwcP0G3IFOlfHHfZRoH1sePA
8L1188khp0h3Sjkffp7cmsLEwojCWc37YVqbMeRvC+ZJLWhjnIn00umczghlGqLO/EDe2AczJP2i
f1GEv3LN0PDKr7XI+XF3ejgUOT7c771zcQaHwxZwJkbNkIMHm573rcIIu2fiymWZ/QsLSaE9D3Gv
W5m0bW27I+sOVksSRUPiqjwlIO1+7HjHBbBlYPEdn+PXpkBE9ZNQgDiukgna0/LdfmssDOTrOAQB
9shcDI/nyuxp330C/Ea+Imb7y9yTHETJTurEFEuwDKuBRFpoROOfYJv6nt43C1zwQX1rvn5Aj+O1
dC1QVHOuE5ymjqDd/OthxaEjHeo3y3+Ma1NGfwY2xlxVBOdryY3Fi0xHj2je/1kqCBHpVrBisewr
EV9b9hjjMRwzy11hboxRsvw1y9Bjq0h+1HvQNRV3Hw9JLjvVtowyCxFoy4SYUWOLNdSt8U1G9LWC
Pe6EnmUxcSN5xwjvK26UvQNSLegHaq0PlubitcSQ8tYjUZGosYwDyVHOJv4WChzVSFn2yfS6axJU
HSZ9iKHmh533WxJgQlUhIGSBfRPDaKbzjvwo1Pni+VtA+3GSJR356ZFD/NSkzSVtbDyPu5pXaQs4
nzs+07B5KgjktlRg5zjVGZt+8RnlYhKfu4LcYHI8WeLJEKBZw8FkZoG6aEjliB4PLvOrxkRJcf1P
qlihLASZQlvYJRasj/uwTL1gEyOMmvaOl6SHAZ51uedlsxEtnEQaraMY28/Lrb+8hSLErBmqJELX
r5vgDnqvcpd9+IkN23AjUCES94VuOC224B7HgwhCifiRp8sGf7MfytiVzHYV9bJGc8UXvRN0DlGv
ZtkpZBV5TqwexNPRvuozhz2y6ddNWCoUBNQhb65Bs7yndFGOM7VOfauZYElkm0FURitpLkrhYL6t
H24Z5+4y3GYA+JbFifU0aYbr3LKSEYr/nFoGDvXueh57cNW5CsH7oO4YA5Yrep2+kei9kTnTNeBJ
/O9bgU26QVz6r9gIdUt0LFaR1ao3FTdh8IEi2H0BdEASJ5GV8HMZ6Rn89PKgvmIUbn5XGyLUXqXh
DCt3CEYgVGJ0gFomgr15QxBSkPxZX2+tzHiQnSDhSxef0bUmFTL6psjsUkTOJIb5ho674jD+C+xB
dtW12Ob2wFwBdJOwBwAhta/6ELN8TZeCrWvfs96g3N3roeh8akHhEzns2fSq36LmavCb+2r6FcPM
iIe4U1RQDMXyFkAYlp5CVt6ABt3vxd/bDWzQNKOfHYA4nQ4KLjsMD9y7VMhMQUxx5qf6PT92X1Yg
jYmWPUlCj1IfPBK9sk9qS7Ek92vEBtQIANu+xQEhP/zc2wcIz808l5N84gglUiLFZLK9CIORUz7U
bkbhugubUYtFzFIKx/wJxsxhn2ofJoNdZ+c/CASshoW4Az5HNCQaN6bVnyVP5QpqbMb9V0LVhcdF
dT5Fg7JW/O0+t+IW/WODOHrcSxjfiaF1Km+rBf2SrKtHnCx8Z4wcwLvl4PSvf4Fak8T24F4ptlKI
o/V0cYeT6nTRo6E67NBB/qYhUfj1xWr/fcaje5vpiro6xiBZuEZMvCAjG/pdtC2zk3MY5i1ekaYt
AeK38jPQoP9yAkqHbcR3vGXIiWumO8I9LhBqxXTvC4LO1KzIVhz755KmM1+tIhFnEH9Jrsx3QUpt
b6AuXbVP+EPTrBsDTrJJiODfUg64gQpLiMpw0ov7R0UL87JrY6qbnODsRslKbObHd19YVxR4++j7
hxOstbqVCV4eEDRhvdLeefHulLlR4NE8hB/XGLEz420MGkbkockwDklcjluocHxWPXibIjLkvCOm
XddpsH/m40c0PVlA1HVAQfLplh4Tr+MDms86EohSafd2/uB9UXtoPfeDAWgSwAhPGyvUt0ANKlcd
U93cHDWAAw4sHAopCItjxsPvEneqGDowViQWOElu8uagYm3nZgXsj2Pw9rvpU2XWOvFX1YqlIpvA
pJUGq5mXol02MGY9GlEii93mqMHIlN7UwwmWpN76m1hOBew1V7XGqdHbuSqsnDNIkCPa0/xatGH3
HXp1EPVebkzJZIOEiEtK6510HDiKZv1Aq5j77u7YtLhytgYdWeblZRZLj8L4PaTudurW/gxLNFCl
aLZoCi0ey+Dx0ralYmwdOuJEdcJpcg62ecUMpZbcFwDc5EXZDlkbjf3rJpd44CVfO+ZNMxnBMDKz
rxF3cuXhNnOf8vED1zE+2useDxbdXZNkH9CZYSAOZmnLMUqqgw5OI2+ffbN6834Y7Qg4Zu9wVMJ1
VOZoqDH/wzypPLqdVGj7oW1eFLhX6bVE22WypRMcUaeknrhU5sYU66xqIFzVfAq4rWgASE0OCsek
Dav0ksXtwn4vyimKlbhxADo+uU5H0NKLcz04Y3Iz8wimTQbMFjcC4iwozZpHmE+EwQXzfUBW6fLf
bra/V7cp4gHdvpqnVY2gJJo+JGBSgJMK5QTpUlURRmeePKg5gonDI47+khRGBdLXVz1S07l0Y9lY
GAVf1MlG3MLpq9ZtDtSGh9J4dG4EeuHwsOPTobkuYoc63ROtE43FitJ7+OTvOQJ7xM2mmum+2+Yv
6630GzDxo4ZjPfRz5udRKoHn8wg9czWiJbrwgieqAqwBZxTKmIl6ew7IvEtxLoiHGE+Wh9Jj0Xqo
N1ft9rOeUeaeajOY9BEJqul4GpU0wFK0URnOeSDPB8skgczAOtD2em/gb6W3Daf1A2JS0AnjMJip
gE2zfjOWpOU+loiR50pbUxv6OyeFslBFvfxYOU4dCRm0RGF75M8g+e3dzYciMSK3Y3zRSa3an2iC
U1Eg5PG1rXA1uXYryqw1P09bVXubcOJd4hJMIMUmOxtNIhmixKRVYZaUkUCupT28yqjoW1RWznRa
jbtz0dkvhkrwPgH+1IxRtv+7E5QB9172p4S8eyUCMolsePWwCTCWBBuviIJU5NYkTHt0KCzYXVMM
apNroOS7JYQXZhl0wgVLHo/87bpngd5PbDa/qd/mstHp+ZxmlKO8RVG6B+2Il+EwbAqW/9r9SVoF
94NSM+d5xWbPPwpiLKruj0NXxrvpeXIxlwT009f2ICb54JCxJdL+1rJqQ7KQ7aAAgC6sZItBPUmv
xPr13B32+HtTPwCJKsIi1hHiTNRu8fmpyYyjSMOqHyJD0X55+RpV4/pOXFQCWA+hAUcAYUVEBpp/
JxnVV2KbgA7bzHC3Iitgr4JBgKfcBsyeO116D8JimTrgYT8GSXGE+XnJJz9TZGBHwQYpg2I+5B4k
KQVSYXHlFe2edP2wPbB0DBnRzimB0Cyooik6qMrZZa8ydGG+co93HO2vBUZhzQGd/RiEH7HS8uFd
hLCojlzSqY0zgDMHAMNNcxPxdNGCkDSra83OBf750QAyaFU9ILtnQWjASLNUI2nnd2LVmJlEO/21
BHLNgw89gVMp3t9UhWLgRF6FlHGjoQGs6hlHfDac0zKrg2rrwsF2zA/d5/2KBg4PQz/MtTJWYw7h
6DiwBL09pPExJiYc0T8I9Ya9H1YHQUwpRTfjA+XB/00KzYU/S8Nmmr56agRklmqPoPIV/GVfJs+P
MRXJ6sXJqNG4B5DCbUeeKPcTNGbWGDpt3N7lxdWBRifoH8Vrk3wHmi/2TDnkSiE8p6OgWYEZ4/t8
Biz+HjJn66s09vn/Cdwl+vwS3rggwQ7v06D8sKh39DOyi9fkuOt77o25Jh335z0Up8O4rXeoSozB
hpZSLAY3zI78Dumb1gsBPgIUmYY6+1TtVOq2f3J44oi+jrehxMMgtfONYjxkk1jA449UO0wyTAuH
5qN+UCPhzrmgS1gM0CAJUMKELNDqeGUq1S8WXim1uPQd70DsD8HObPx/BHiRIVZKrKR+85QXJ8MI
zn4lZ7o2fHVK6bH/WG6TpEJE0ZDmrFdiNJ2SqriGF8xANLorZFgnqljd6YEIyXe6n1dZsR5JS/YH
OnGj6hkAee+XfZL+aTm/ONQo6LmOE+BnunRJyPW4/eB62kWVaI9+s28wkGlaerdAm9xCihCLrFc3
LJHMyQPA8pM8lmkWQwYyEYC79OUEsZ3MwcGRmlp/kIKmWedOymXTTf1HRa2fDjNyswxwVokc1hnC
5A38CnKmj2Fw/OQoJm+hSVsRAp/m3tNd/dDLFGQFkoBYRRgGkfw0eQpvGAjYh9bHtDqUgn4iwPUA
y72WIGTU1Ndx3r3p/6l7+AxlYHSCwZsUpU4+LOAC7YSRnhzh3fqL8hIMkcXfHSTmlE4FAvhiCQOP
dc7B9z1lIh0fFTJTTvrMNRxhJel3Vx8OarrFuStenpoi2UYtRQeUZnq4k1tBRAhQu02+BhaLZQrH
M/hScNnuQDh0qUcas5bP1Dk66fyRj3vxs2eVaX1PnZVhPYEKzca4i1Ni1Tz1IzzUgMVc3fJe+9NN
Cj3tiS3twcDHBUpyCEvT0NkaUG89LRTz85ZAkIMgjW5TqQsmTHdmjsXH7/l+oU0PwQEXCuzrBm8I
R7eG1HYuEzUld+UbQx+69A2n0sOKpzpYWqbNA3/arBw/VNk6YOccG8h2R4lJ6zmrfmVLBcLQQENE
fHE6ZfOP7AfPlEogDyWpmFDN8Q118qo+E/j4uobfj3RuqN6/iBdIqV0GH4flKj9yJgK6AJsuCXr+
K09kAaot0HPYTMqwiCttjpQQfdKog4KAxyAt9FcQLGpFavMjBUmTAKRI3xH/ZW50Ofbert6nBzGg
jAmOJJsKSOOQxDCKph9hob5IP98DE2+VzT+FezgRmgUz8Zg72ooz7rBWNyyUdePhW8MD8dUwP0G5
UzyJcKQRqBtYKPeCO5s9XvLAVBHcT4yxclPC3k2EfGmLNxSoEtD++o2qR6YbwsRjgsQKCtpYy0Gi
XjG5pFSFB6FjQ7buCw+b5zDD8h8hMtmiApM97dPxS/f9mhBTv/ZuV5gHUY6BUrdiHJ6dfmsbOiF0
F2wsmRXMowJW7ZR1bABWH2d3y1ca5XlzO8E3yNH1tv/WBx7PsNBzdXz7sSGaNrd+elYjmdFkh7QH
J8NqbDqmKTh8ZLnmp2YmfBMK4Ac7IQKkGkxKiam7TXcD3vixO9uwqjJvqgz7cJTEadIDyr3hP/J2
PyhE36q4y/dbaDbelQ7ocOS1eSQqg602cjuzyW6B1Isz7H/JBYnCX7YvMnIo7A0WT0nArrEuX2nf
s1F/Zm7lwErzYRKaKvXGsRk1pcJ2qtnwZvky1VJADpHhvRHaO/4FM0B3x58FOAJtG6nhvXpXpFer
wWAPhyacZUk3UGK7cipq2SQIjWu48gXY5T1GsD2Bc7V7dwgSMRRHBbUbMWg3RTVQne536QlA1Bj/
IISEnCbu7CuPxPFX99fXAEMJCgMoyJqve2NYMPlw8d0S0+0nLBNqWnkH3I8bPxNhwRtK1r/aHtcS
5NOpVEp5l/5Kc1iXjFHCL/HHta1+yyPwQ1mOtrJ62dp15U/Yj4uF+hZoDZ5yaKAgLBPqE/monEcy
usoE4d78xvaY5Qfbzj5BJ/1YkinAIFhbt32QgOnYXErRatNQzTi4bCquPsR7jDTxOyjakjO81YrY
kORP+77uL5Zh+Yfy4QzcIQVsZuwWCTxYiD0al+UhIyXaTkNP902IRsoerXrUV9MNmI/N+LpL8L8P
gHWZSauT9v6hk0XfYvcDO16fAQPzKqROVNE+Ijd+ZyGZ4Jw7nsJHpBS6IYlBgGr51O3ScZIG85ao
b9m0NrWEzMEhnZgRSLVvBTXnGoH9KmUlyUrVqW3CaHwgDRkQxBA9gunwP0z5eMVP72qNdZIxg5TE
p+JF1puTMBKbXPAPaX5i3utsSL9/e18jWCCw8fWi2DqOr/v96DOOZCjSD0kkLJ+j7oHkszG3lpAE
g2xsX9EwuSUs3pQxZFQATD8IHUnepIMZy2uGNLxLVGUFWXpXX5pQD/+N9W/PPIVNXC6HmLzy+ihL
se4hWNDh6fCahe+fZdnMIV6nHmb+CUOmSBaHkcu7V3xeYjDwtKhygz7YKRJrRo5TZIBkIN4ppy2i
9njhq7HVOEK47wtTMsx9T6yZ2rq8w788Fi03GsQeuh83xUjt/s9MNxa6wCrMpSpXtzLUg5GtrRSh
MvdO2Tf4zc2lTvoaV4jIAuY0ZSUvKQRdpAmqrGu3WFycfr3lKyl3kL8CC0tgBEnjpvlOcu3ZTZU5
VJO4D3PtEstczfnGkGz28WZ84evCOSJJOKvsDsEyatufXHnCKV8rXIGcYxmnyxPGnrnhxofBXTa/
jVdH3Ru7m0oCKuZoZXbhv4Lb3C3TF8AN1EcDS8nJ48KOUgRqwYY9diPPrOeljiR7I6cBs9d+sSFi
l4ngsyE9OsyklkUaagOTNgtyQYbHfcQzq7txAJWn3ojXS0y8A0Sq3EcupTFrINBtHduA4W2P86FQ
loYkXCs9SIPApHm0ppywuTmkp3fJQnWEJezybj7FNfMlOJWIu93/jdIp3gTdmN2r8M4+W8S8l9Ox
7767LNNGSScB9YlVwG1aSS8gn+xNlk4WY9mM6mZ/atEiNwnpuVjXn5DocWohAMVveLlozYOeuSLS
9AEO6BHJQiRzaCt56NZXHf4w0eMWpsPwWKM5bkJf1ON5ES5QN4QDgYjnizgUw4yjiJZMAc0d3AbO
4Fzu2Gv3lrDOVFBMWqLFT1th5gfsrfFV11wxWekPmUenvJKNq5azOHEbdq/+wCq5FB/kiprsrRfL
e0CdZgckDOhxHBsJaDYCnl+krq1RUrhGzKe4JlOamwt70y8VYv2/3c07FsAgMG4+1z8kEkFRgljJ
Zg4eMvvioYVJ83/uc8TYjwF59gzHLl6Xe11t3TpGcU8f+dFvIwUdNQ9JpnFCf9jXNFbnXC5Em6wz
zpALuBQCKmy8o5FymatWFBU+i+RlBiY2aW8EODEGC1h2CuxpRJfg4aVxf13O6qCTpW2us38GBcG3
QYB5u0h5TuBbKUoCEVObdLXlFZ5wAMFyb60bN5qfgsDTgTC6cqE0ISBh5ToGZcBAkFh8Rb+qznNU
xGjBsXPLGusdJ8Zy2UfWvWurSHI7EtpJ/uHPDvE23YqbJrCDYSbnGA3sGrVT4x0O2asP4IM4oqLN
7XH4yDW2IGf2E3KM3XMKT4lDz53CAhAkkbgGQrdnvE414ufoOWuBdclfFBTrP9vQrZCPV7gvGSVu
b6nd1jbbaDEFUca2to+kNPz3qePEPFbFXhEZFLtWBg9p7pzDsgLbhoj+LcooqnGv/+HhAyh73Bwc
r+NjVLqOMKRYO5kbMZQ7CfcCHxPcZXG/Il8M2FtOVY4CGcDv5JTuEEm5P7uTlOhpZzYcTC3gRAgn
1D9TX3CPkEE+hM4/Rc5Sf/29UKq+gh3xZvVfhlOhyu4v7aTj0QxolqB6bo31ArjK5tnaJ+i2a07u
tlw5tI7nkoPcMcxLZGDxuFKBmloF58NWXGYILU7YeWFC8chq1bGbGSrFkiprn9xENVOtCDxY/IfR
7+VxHmz5a8uJiuhXYroxuSmndUGRN60btvPxaRtjOaC8ZOsHzPGGCY8MkCZ86S+xSzjDz5qOnufo
X7bec+cFlu19YyOu5JEiglGE6TWCg89ZK2wLU90tXnGcVKR+jEPSXM4vu1gjiNXVCgcVSQMl5rm0
WUfXFCO6vJkpvn2BsYxD0uVCvPL/akWSNPM70ZBkOjCEEm5adlJgAmtdA5Tail0Xlf6zQJWf4zXc
KivvDGg6989LgWmuLHzOjCqo4gqjIOiA0NW/SGrLrXvZ8ng3MJ6IHYSmcgSBSe4gXDnV46R902Lg
Yn1rLa+OYGWo/ADLJ1cm99pUergviXZmEJA3Qa0yzda4093Z8f5NwYUdCBg1IcpPQor/TzqobN+d
dhrJJ9ISOwNv6O8cpbFCrzS4mBOIPW1lmBRT7XEKaunW1oFinpQUWCNPKuo4rn0lj15/IhSa0qY0
FkgXZvNshBidSO7oXha0TO38c7PoQCoeTQqpCRYXCu1MTgVUut38f2dNt1eu7v0CPsAldFp/FEcA
50kgNOzxj5gINz1RtjE2Cqz+TrVBO2yXDBNPtzdWzsahz0QNDBwVPgbiVob0LTniqj9Q7WiBvsY6
8vuJZq7rbOg4J9NcTu1SxIOIYog891+dtb5x2MG3WsxnuLXcRVeJV+SV+verIkhnU0IbR4z1cBUg
NecKO0fvM5O1D30iqiQn7z2E+GM6hj2prfwUTkvnzICquF3v2g3Wuq2iACYoaSu0FaLvX2IYFcu5
aB7g9+P+L4qmy3fBB0aWL4bOJLTxlieyi/WMXKvNBcGOOXLhH19TMSlS+4do4qaa0Zuf0nQX5n0c
9Ca4CRVn4kWOBT/zLUloOTKwGeGf33I+ZGKD2n+52I+qGmAsnERJ0EDKu0EgxzWC2P1PZ12WCUO3
qKe7p09RKZBpcksq4xTmbsruphvxKWqyOVExtUboDuhM+86fC8154UJvKQS0ObPnh0owiJf/glfZ
QWtiq70MSQUE9L7p22h8+kfxg5ip1hFGXF3eIDAwENkBrTj14um2maErIj9goXZrDVsjAELL8L2k
NINigRB9ZHK2HjKz5ygqfiB7I6OogCDwVlbk9bhvevq2rKGUefPXnxiFDm3s/uD2aKdgzWefaE4k
HBMA/uzlzzMPD6dc0KfimjOcVcn33a06CH5NDhGy0CNNpI0lIByM9HDOMO0jePb99MnU6M5P4Sen
j+w2B+Vpw4aLWzkQdIK/X8IXEsTfSH3l3jRxQ0AIZ66IwRVa34Fn/pXaBzoU+NWrLfSOhhLjkL4F
msR3d8/MWBcmjitCxi0mJFdt9XpdyBpf7YGNrdyyEntBWoTvTvNfqFNIZU5GftrrkPXeSnTgQtUb
V8hsh6i9U7vgKGgKsmZtHSg2p8h0H98ccfzoem0shOlU4XncfGkO1AckzHofjjICzsDuO7n1rVNa
ENPtLWx/s+0mxegYtDH9bV5YyAqXXerr6Ov3xyzIS3m3KJioKdDPQnGw8VeRlhqUhqZ5rXept71b
UuwlCVajcZqcOuA4R0ysvYTaBmSgAdaaRhRE1/nu4RmxNTWs3Dv+vHE0W5p3oZQpx09XNGhxTvEk
0OJcFzcfyUaVajObmq9nuDTKszp9XVsANwjg45zqnN40tV76OSZwvCuyO1gmNcolh382DdFpBc/P
1U49NXvpn63QI3aQvXYMzMyqkmZHig0+/eAHumpuu1+O0trNogNmzNHUyTghmDd8IOJJVYb3rtda
ePCr0ye1o4yUZp29QQoxkgBsbYfDQucy5XJJJhkk+tHpJbMtlOAJ1AoH8opmnpaKYx6Es49bhBhf
47ycgGXp+XmzX4sPWed6hF9qqKdGcbHJACY2D8QBPehmOoG4mwkgZQTmq+sK+TS44agiS++Phe/1
U0K98faGhr1HfATMPgEOPj4v1OcINMBUJzNXmKZHBaiQo/yGXy77Bwmz5w13sJEx3ggt+noHFpFb
AJDBQ64ls1XjFTO2Q/q5xJmJhjmMK1hdzYAmlvJ4GHjocGaj8ipgRfj0Db4ByEvRDxIvgWyFg38K
vrO9TZcX3wdb+ENLJiTBl6w28uAf93D/74VnSBG9tl+9YB140HUB8K3jqZrJxC3kVU41T4mQTRQT
EDFtatp5ajsx1oFC/9y8Fz1uxw8kadIUvprENVZ2qOVabyoU4H5bnLDvuKr292rllOsWHgbEsTAr
+cJgjAIv5G6vwkeriAYaiwRQESIgtx1C9qSXl898cC6w/p5ax2O5JM4vDZR8ukIZG8pxBzTAAiQL
OGRtXVkqn5sh5bxazOiTh2w8cOqey9dYCC75qyaE2pJGSOhWSPzkr6xmtLak3xs4lm+ipypDgbpe
mgxwotZhtdMzVMRbqHPSOUCxTtzUHi19EfQH4BqPP5Zu7ajJStUvslKwLM0xLmvBiGJOaPCcw9yp
N3ArjX70d4PFb64tXRLPk9B0POZ+M4TW7QZ8WChyMJyBB4MGDSIGPNyI+s5/W0EYoZmb+USsWXXf
RD29xedW6Egv7VbhGXWOKOTJATaaplwNVstzmbAI3Vo9PCIFsniPrWTELA6TEg9vGB2899CzbVp0
rOaHmVhwf1x9UWIlB2N2mGxqMYl6Kt5/ImAH7ovIJpEvSU3DJHX436qO2bdZwKoXWwoEbPjhxu5C
cLX29GLe79+3fs9+1B5ugtBf9+j05ZDWKqqXU1AVjmocGhNMj2FZBNMs+FyAuwgx1xQD6eE8KSpG
5i/pACk8Pm0gzlFMEH57czHk4Whm2gOO5gjv8nYb4zvy9yQa+7HDoqSlFT+fWC2XR2xi1pafWTq8
H2azP5ienMg59dOjngxe46za9TAeGuqmtEQW4I3KdMv7VbBGd9IrfiIA708JFVHjISdHbHYp2AGm
rTJ3Aey9mQpBBkYeehialgCm/NO/fAkXrJDhteBnuaNS/g56zkj1QzZijCrEz+3WsxLjk0tpITyL
uOgiwDhPEXjockOEIpl6uLs/iO3KzHlJWt6EYKxOyy4AY7vJFX9Gk5DXOWNj6umiVyDD1GeC0BpG
e29cjHnEiFcVQC1yEv/TmqcttRzKTGJxphqb1XCMiR5TzyfQy8Cf7mEETANdZ6DQuzGTH13/4i5i
96vryLg0VRwT1aSM2hCIM6GOQKS2ITOZtaqEfJy1fSxnpJhNNEcyDVup5sksgUb73R9H9Jbpl2Lb
zTUbZBRV6pH8T9t2iVh/wBblARqBtslVpNGi1S9IYwlm2+oh589r5uhrzswlTweGYf++aqHUE9uS
P+chlXyZDxd7LU2YhGxeBlcSlubxWj/nLzmB1E9Nz2X9xdsURy5cbU3Mxeb0jOJeUKDVk0NMrBTY
BMmF/xRG+Qr6uRDADVtUIX1xWacSBN1kGGHgSPdTtHXoUsLpGGKC+N6fbWCk3UfOjdoKYt5q8QAQ
UDIoCl0p3iCbMRv0HtsjhbdFFRaVtgf2U9fs1hfTGsNes/m5QCAMZbvS/Z8LGsa/0oJsHS+DfvmH
z2Ne7wGsnVeIXtsjls/soVVO63ZRbXq2S6xXFw0Wh03plDBIBOuhVA8G+YgXMvD8nU0LdO8CedQF
dV9XtBfIf/DzAS/OMLdA7BVDTSnMYu/x5oE9KYNexgYetH/jSI4pmYgvFuKzOj6tT4H342j1swg6
HMyIu2kIdmIzQ6Qg03w1wuttW1Ur/esnpfYk1Z5bY0h9IISXG5OliL9kfBTYVxeuljCQspCRN5Lk
nbOAiWcA4uhwvfDTkOvYE0kdznIkPrDwphBRdk7E7QMkNPXZqbihSA5jMDMW01xNR/VkvIhj/t4N
g+vJJ5zZo15L1N1W0HNf8regEQUuvfUisc4wW/tJSjbFE2jP85Wo3OC9uGqo1W637EQQBfRxIzEH
fDV8TBvLK+6xM84BwRayfzcn02fD/Lax2BsiHaaLbq779WEK/xrNKNixjC7Edquzq0C1WeQX20l8
1bMV6RnRAz9P6MWnva93/ME47VTfYOi/uS17AtsTJl98mJ4hKyMC8K1wPi0ghwz8QR0SPYxsUgNV
A/HnxGqzPDEDIvp6drDczF3ryooZ5RqeyEJ585scibDO604tf8htxsR42Lh5FMfoHSflIJ9bKDvI
mO9JXLiQ8YzYYMrrJlMqyjnr0hTeAjJK4AKjt5subI38JxIKHVHfIip2mPtnf4E/kusk56hpNUNr
fA8TJV6TbzCEUE5KVu/2IHWiLZ3oEywHoV8M7vNrP55w7GzD4nA1GMbgTHTxe5Mxg7N/VETI/h+b
u5yqcwqrWTqBKQVGY9M2Uyz7sGRge0sV7SjqBquR6o2AgiilI091wTwc5uD2eyLl5CH7X0Wv7zxj
WIKL3seJn6M6kjZjSgkszH6w77915L4a71gEfp3U2dMVS1yzMuKDG3b5NZNByYL94gs7NW3anSxt
cGND9jN2/5jZ1UWdJxFKbB7+8cZ0Ev4LyLm3O2UJr1RvEZnX+LtN9W/sn89gK8sCBfZd796Ulnd6
Iqm8VZV7uxdOwUyd2Gcrp8VRzzcNnMf4q7u9QtnpAfjLNnE2UVozPOa+JWAlsuM703AJjz0dWu3E
14IM0Qs3Wj9iD96gNAgCTI8ZvW1T0bDIIr3FeOmtVz5zojPl3Gpg4F05zzdNAjhiWKb40XKx8/YG
Oalbsj3eCWxYYmUOQBK9O0Zy4SiJoci7YpZcSo3iwzN+7Y8ONhzW85s1ka/Dgkw4P5sQ5fpoeWoH
NDAGdY9Iq8z5/Rez+vcUixebFQTBfk2AarTwQPQ91Z2lwp88hm8UCwgoE0ylZM6O/xRWRwky4n6i
jIfT6SaTNmNLwUaTGQjlFv3yn62nZde3R1JKmoxJ4vqtBzuHXrVeAgjQbwd9cPteOajkAvyeX1OW
gohGaq9Ax94RVIKuQoluqRzkv5USGuBDJD97/2PkQIv317NwZqZTPFlQSvhcmCc/7r2l/Sh5o9X1
qekFP/3sLpkm7XrSagXq8izINt8peQboj5xCx53w8V/RH8YSZENYUM09qp0fOawRChCvBbTPhe8O
gS1Up6t1oiGOrDYYvtMGWOMTrVG0cq0HwzyQp2BtpTXwHHcIu9o+GcsGGOETd088+0ZA+uEfgsIl
oTBJtVvnfYjrQnwAAkwprOmX9QOpUbQWQEt/rthtn0Thwrlwy7hDgI3Ns1RcmnadCU2m395EUGBH
sB/7TL0zZ0VINssaQVJUmoTBo8PANOkBLwLKFHtzoOs1wIXLsMPvDwNs3xYvcArAf64RHvGbiAJ0
3I7k4sgasFXzHOr45HLAGQnDwMq5me55rYrMUCgeq+wWBI3sehyIAhwRAGDRNyjsxYL4GfJK68Ff
fj3WGp5Mx3hY84snPJ4QkrJ6ORFNiYaxkf767AK7EsBSuv+Mz05XTu5cRwCYCZUOEr/6/bZkfGu/
idpXbpRAwcZeuTRyJ0abE5lHgfg2wl7rmWgioGpf+smdiiaHY+6uMdURxJsmla6grYhrQnqHX3PR
Tnr6E+WMvir8LCwfFlJN1IXaJqLGGqPiOpTR15RU0EXKOG9AzpmmvKcqDml1oRNxPk0S4TX8UiQu
jOedJxUrO9t+jM9T4b3gVBWDB76CZOUHXFh+TPqxQLJmsL+tKhu4Z0cnf/sd0mD7oJCzxdBYzqIt
GDeTn4Qg361+jd0QCjpVT0vo55k63YiqOIqwSQyW2mKjLsQJnGHyRdhuzcCBBr0pfAGoIcFar9M/
0jSqAa8wfDUEibcaDV6BtqntzoqHX1k8v/3cSpIA28/2wW9bnjkol2gGw2tR4bvdNkW1kXSSozZf
/kkjw2jMmzWo/WcAmmr1kF4r6KVaSqvrj008vbRt4AYmwcK8mjnjJi7THejHz3xuLjMBchSNjSo3
mVlhTGkZRU/hgMhEJBr7Kp6RVTHZaniF+FWr8hDmqidkwuBlzj1yc+yk7yz3uHHvQvUb7lmArKvi
oLbhwHEjEAqqA/l3EwalIVYjJ2s9iPr3cExJ1u7X1bpw8Rvgxvu6GUXxBYaFFszAaWa/M+k1TUYq
JJ71YfFXGwDGwRcpq2l+xHsIxVnRWBiqyd+IfpYov2R9ctBVoCJjvu321UdewzGHgrWkfrzaNB2P
dYJ3mfHdLtiLMrzxWqF4a2v9P8NeOM8Ayb7tEz6o5t26OBXqcQp8X2+v40Y8MjCoPQ63GGnkL8fX
66eaJX35XVFXnjrxRwBkcHKo4x8+lV63ceRrGmg+5Q+zI0FbaP0KZRyQCk+0I9fS8DNxqrbduJAq
gcEdNiTO1HAbgBlnSHknvLzXNMXOTtyQwEIxr5YcLxCaRDsxhsgjEGVZAxG8uEAncOS/Z5BGOGqT
FHjrKpnTDgrmPA2u2tAZkvj/CQDXXPyU7CvqobfcKNotFMIfuV9eVbqOPbhUTLLCX/Z+Z5XXcDCS
WcezPsMweJo44m8m7DSDiaMBzi0AnxYUzRn+YkrG9Zjor0sh5D92A7uEIb7BHwesoeZuxdy7Nhbj
iMfgADvSiR63FHVsgN+9mG35KT3OJWlVZBoR9c3F4O6WU4035/kzbiZtg1Oqt+0Ty/83+CoxgU2v
pcuBeBXgtcRBaAlflJl0qba8XuKOsMs+JN/PQ4iePCcfXuDQeUwh2QgEEFkMfoe8qYiseofnFfq4
tuuzRZdEZOnFwYBoQwkdNC8ke9s1EuTA/6VPTGoPgAtjs/zaPvMQNFByLrFHRwoVVJeDCtBabpnZ
G+dwDf/3p67wJ8l9LNYEj3lFxAIltnJvDwQhNUGmVfgFRq6t6W3NRmH6je8ohHJ/QGChcwrAZBJV
A1UV4YZC1ecfkh7JoUywdNFGb2FSN40je6Sqy3RnXXFO5uBaLRye2UInXf+Tu1ZGsA9brzkwITrG
Sx/BKJXakXMJ8kUBvKTSzDkL/qqkf2Nd8t14lwnbxGmVYChI+1uGafK7Drrw77/IimRNH0dDWvyD
jZOFWF27cBAJD6THQ9zC6uR8a6P77acwz/hbLbmZUAIno4d2o7Oa2awdRy8FDZ7dIGycQtR3iQdy
55FRN4+3kaHVDEaQ84dgxXdjBEw4z/TD+FYqu4z8M7VjPTxhIroZd2eQm/q2Zu0Xo2uFTNUxRnj3
bBp+Kb+512E0y7JuaSvfHvjMRMY3PPTm2tO4VWgmZ0/woEsJmnDitqg9N94OuBUB5a+3C1nYHlDt
jINeQNewA1HJb3KMiws7P1Ks/LQQ+bOEOWIZBvuZg7TWEwCUVxI8JkLl8hsnJOkIwXExaghCMdQF
Y6Sx+pTv8pfnhb6iARQKVpXgaT0e+YSxXGoy7YUeCl0aUzd2eKP0UH4RYx5XuTqklLzhifIAnRuo
stbwV5cgOtk92JCYYyVWdlxbfRN7jidACLiYYIr9tKnAIDVZiAInNVoC2EqUR+DLt3O5ge4E18/f
jIvSxqqJIJMagt93mQ48nfuw0nQekgrSCbjCubHYSnAhwm7lnGhoQXc4ou1CVTqqMvJfxIixBeTY
gN/lqhJYupnM6z+oHQLLG/y59Ce0b2XrsLYKT29lZPWwKBkVQqmUSCeElbqDYlVvxPASrLyk7c6r
m36xdXDHLaW10inYngOExiwjnoyWJlkr0KQmmYBRJGWulFvkA0ayedXnk7ja39PtQZjbE19zm8yk
vx8XKfPpeASbH/VATEUisOOPcqdJgAEtstJMeDk0lPtClg377AP4tfpXk1ASAveCi90dsZ5VQyOu
mHgc6PGiNIgYMMAyyzYNpOe9rxJkDy1h4uToJp8WQJL1AEnHc+jEPHI8kc/dLyrMvH6GbZ7I7o99
zBxjda6k6xGKPuTxCKVjEi1CE4zqCNDTWbI7lAxYQsURH4jpPtElv+9gXNJRwzFXBAYsrgqlwtyf
MErU+3rr7bc23lpImiS3rXucha8P548/ovgCU3ypBOAmkBu1cLXV0zP+aT14qaIz9BjC5SqHGDQp
bUAf9E/OfOd5cMYQzP/vVh7a162qSdwXXyYFjYKwKQihGsmmyFyWEHfmRVtZ28fw9RJWicKT1mCC
NtV6XA5QyZSPds3Hq83Ts4P1xGGcGwriJPWSLICGRYouv579NcRyUviItTeX41+3FQgnoO0kc0fr
z1t0EjQWHON2HnSwFF+NsKxEMez7v1QPOTzCY7CsYK0/IcIgdJGdTuK1HCI3YvXeMyLsVTrL703p
zMpratluneb9gY/C5S2BQpngZ03Nh5Fnc/WaKeOyjadlqADihlLycJJ4EM3QZA52rTP7J52V7npv
J7LDZoigJzdqm6W/KSm/pBtgHMPZXz6z9nNvN1hjjSjGQB3s1vjzFAAD6lUxPEB9UOQlu77jhFYk
oREjQaHpAg8a1D//qhnuhAL+vGmo0WTGPXnnp/huCVpob+tiCv2OF5QpVUPd7ltdprQsRbSL0g9Q
3CsWf6apla57lwRIrnJU1oPwFKsC9ag4T9bLVjFY0XJuqIv9pc+JQiE35i8Kv6qnCJQtVtEqeDzz
MHDBqfB6eq9EY0ggyr7fPH/fYGmOozqLmSpac3Q+O7qch9wSx8c0FyGYnnbIVO+U44I9v/7FmEIo
2QyvwWF6Tn8+U2/DP/pRYpeWvNav+1ZXxF+CdzMp6RzKtP9jFjjAy3V06GbEOmHdq3L0yak9gU2n
j/9l4SiPE/W+8aVKgTTXNQl+/lJaqs/xf5gt54FbpYfMgWpy/+feXkPJlAImp7qbf+HizR6FHg5a
ECtoCBb/ujPEklM7seznAgcT9PZamgCH6vH0+SVCZ2BEJ3MpU9iTYt9dRXe1K1g9svtYn3i1hfg0
aEJrVgPCwlJuaO/AaaN8TsX9mDMHe0JVWdxGDmUgOUU0PeSHj9cQrlw+AFmWYqCaQIyJiJDWPalg
MEdWgxFLx2hb2Y1XA29TVXqa1fYM2hFfHK7k7rSd/nGVzNoI5XT9LbLccHAfj85wKkWj6ZjtBKs3
F4pH7fjW6mlJ5/UB+fVlxf/ZNhNe43EryOYGQXdeI262OT3CRab1N5el6G7dahRbnjzyBPQFBT/F
Lq4aQ6l0bR9bzBaHwJgdvsrccAlsAsku0NstKKcNPCheo2TvcSmmxip7CcNsRyn5XIGWwY64oGi2
nnYvD30Qr/dngxuoc11phNM1pAE344LlLUbEWF3zhiAqFjBBpUDMe/wMJ+O8BO1QXfLX6pBr4TX+
H4o161pAFSMVI+H7BW6ymrg+sOzN1gYRr1izGD0TDmKUdv9xR1guupESt5dEhVxzkEVZ1NCt4mHD
iKuivQ/Z5yllD2Gy84Q4yM+DoyolAFfbfjyMn6gK39QQddaHhiCdO7dfRJ89r0Y5TQLOzhKPQn3J
OSdIHOdKMdjCTqGhBzjeNnWIkPoaFbF+Z3JaB9XLKGyN/xq7dZjHK0oaS1RAZXLXbHnQY/nQbJMr
AGuqYRATCeH62tlJ9Lscuuq3aODOEmfyWbyI7YiejFfOcyV+Sjqh841nmsiYKsUE+ScYGuGpJZiV
lc0t6+brkrr8dfKBWytEVt2lQud+nV2FJkLDe9IICc/e3Xf13yJCcgxDga25pva6tNL259tz+Cd5
ccDZBKZxNgLIXDSjOjRKOE2N92obUP7/uD61eUrQC8rNKpBYAI1ZR57pvwvGF/0988oNlRz6rc7m
VtVykrEd/tGEmrL0JP2Wwk7kQcoYU4sal1mOs6nd5JRkRy0HzLYHIZrwnPkYU+ku1D6r4xfvv6kT
vMll6zVSltrTFgQOYQQJccld/PoNLCO1RKn+MbbonABcpxstIA/CfneY4oqSZz+c81h3NWth6lQm
COo1SKzXqqEZMvizVJjryidosHETHx1Nvr4GmbB7C8rCecHjnkNLd7Oq4YeoSbkGtVmdUuYHtQYh
CliPCpwEdLrEeYBWtVwYjq4QnRdeyjqaMK2ciDjk6P9iCGAbz+7YDBXgtG8Q1GlegiISpULgT17Z
OwVHrJuX87jzy0T7uAjSbYkhuY1Y3RgP9j49NU+hvaSSFZxKj5NuXFsaV9Ls8is3p0QHzzIMG4Tc
d/mKh7qX6s4IbL3YPQ7tag66jwvSLqpAWlDR8bGuVv5YEIdqoRQ0QwHLo+0oFQIbzgtusAacARbl
maeXuyrrM9TsM5H9QZbjcd3pQl/bRydqoAtBH66117K+PsBkfQPgvXdSalTHFiVTnJQJFN/HQb8q
6gorYzqm9mKEZ2lyQqkw34tMJ/zAKMZ9eogioDHP1BTCw2B9RpCh2r0KoNLI2VYaR+g3SWLdEqrj
ZwkgTeZ/PJnmvE/EyjWzA4jyOSf8MEOUtNjv6lF7VOw3OsUbpgGwVP/aTYOawody8fhCVA7FJ5We
vecHEjgC0gle/g9g+NiMk5O3rumbjzRTOmGF7HMp1yCYIidYGqbHnQ3RE9lq9zQrok2834X/iQyg
aMBkZx/FzXCdOwHSE7bH3KP3g8oz0b8lLupmcYRnm/rAC5I+6E6LMR8cWLGqQ7AXleSQNGlxKnzY
280XbLCk4VFXeV8b6Z3kXq8YhBWeyKGzGVSQI/QchzLM8w/S5u13LipApUPqaJK2AgXge2TCNJ6b
sz+AU56Lssyq52seYxM988jNn9VTQ5Vdjl32Dsj7K3ju/aABGGZrOuKQdwnNWZR7YOEEaLEb3xlx
Z1GCMvdJ+ZfRAhSB66G7RKCkkC5+Lmme4VpPj6CpRcWh8N75dYN7FQDKtvCIx7BcVvodmmLbpkTs
kbs4Uqw3KKFxAxIhSPEFHRPml4X5wpiAQK9YHS1Cs8GE3Nx7Sf2on5y4McY98s1ZqJxm0KZQZvIz
elgPtka6PWIlCcCGsAHbJePq2NGEc0CMzN5gCnhTMJAcZBSZYUOs0LxQM2Xmv8A44phT2kD4MjnZ
5cjeBIz+CjY8RCQLIILCUXpwfyUQ0G/tWQjzG96rc387BPh1eJtDwllpIJncthfckgd7naODZ/ji
ICzGs0u/jCfv8MppapC+uo69dcovDGQsF2UVFd9TdHdIFhelwYRrWxcIRoWGOdEO2p1Z9PJijunx
I85EIxBx31ZX0IkZZ4FuYr5JWD1IekG3GahdT6juTMj1kk6yik2uH7mPPXMc0iFvPDQMyOMvpy7B
HWFQPN3+7uQa1KYeswuVRy2xdwx4gXkazoWAYH1jZvstGyEAgLuvicHyQ6v0W2mML8h9Vm6iRqrH
jd+IBU79dfK3bciWmPunI4A1XT2zMaHIrpaot/sFIoRErG6Vjtn8js20VyAPTLBqgsPRTFfMUNHv
w6+4e4paajnBES0ondpzuFzE/VSSV11afzeH95Wgt63bYIAgT83f2EZ3c143hmWTL+Ls0Pj4tMys
2KYOxd86p8Ofd7c9n7NUoM9oAxzfhS5SFw1Fr4OJ9ktOuEvejO7RU7PijOY8QRo7ZP2gwaCY/1Jy
v6azXxfcJWbxZfEzHKwJiXdravG7A3tziyoIDHYgNAp/eWQPDF8xCqiHEt3vqzwFvblZPkI63Gpp
V/uUlZpGXmDlLpkXzS26kYEnR5JpqjUwBPGDSwlVXgOPDo9Jt0BUTf4GVFfHoOwTFmBHnPHSV3TY
tFDs5o7nPoWk78LPUgnUYvSEi8WSHE//dZklwqgCptTCe5l/s1OUCX941hnMbCcBLekqHLyaYQ8K
f9Y6L0lm+oitRBIxJ7P8nFQ4kxXu954mGMGQRxXnyuRrlTf7kQeF42teoTePPKUSpozsdwl4xbKk
85uvIRHP9b6d1la4HH3A1k6j08FdhI3RBtylA/jHDG32nH2XgPZ4XPbN0MgtYxq+KyEgNQkQMZ9k
A7t+a24oF0obE2Kr8Zw2XxPHOX36ALo4s59aFYVEFM7M7XhCewFMKPzcUUlScTnacrz9keF3dJJM
vV9vTtzaArSdRfGsZ4kocXdG3O2akp825Lyws2y0l0T27IstNocUtgpnuQ+HCJI5RDHxQVT2QL0V
Nu5/JZjXjLPtSI+vLe25VvpPkHHdlEyXSpuhIbqXHlOPhpeexJfOcvY5M+voLQPAxX9jxKWT1YO0
o0bUIIaSCs+eAeZiw1mgw6ohnxsAKHZWRP+26nCCgFT+02ocQEetMkdZ+5JBaFXC2c33BDu6Zn+6
GDN4H82zWiGkbgvO9FvfFvrdL28+/XVN2HiaZBNYjcXK+Sj3/BERAGzrMYK7U4gI47GEn7svZJvJ
y/IV7HL+bf9OyQRFkWa4nI4pliWXJZ1ILLzTzTuUy2OWyVeBYEjsuLSlYUs4R0Q7x6MI9quGOv4N
WjvZHCoz/Ttrt+Mw9m3HSt/6EP/74BEMgAL/0VCJKBWCPzwoQ9f9zFRX85cv9IUCJBFqLXBFElFn
xrR3bNcTmAyx1LEj2em51OvJwTr803HDhc/y5Y4gavPKANo57BL3gMknHiCUl3eICSmQtlZRXOU+
//PtULUvSJm+GUqt+RCDPStHP2yoGTsnJprrpuXUl3crjLIL8QwzPyEy8H0KeqOR2wl9I3gro4oV
w1PeN/QzmSEv0NVm7pu8SuxB0xqiPJ86LwTuSfuzQvwxHu8pTLeC1u/SWAJz4Tn3aiMLNqUD/s2x
KRs1WhWfxfAsnyjh0mHFk+gYqz2w1z1qWS2runr3wISXy/nnQ1VFe+EjcSHvNKM1MXyGmmzp2bxr
fMZh8Y5p2eyFL/Df6Mn5WHx4X+Rgl3XCoZtDlKK9yAveKbqUi0nb7gaMxzBao5cqxvz9PegV9Dxs
8XYsVnd3PK326L8lZnJHPWeBool7PI7EKKMPAW7ccKRB1a0d4P2pjIIiccTitqNL+Jj2WLLW6SLC
VGax2CjWRoGojPyElBpVPQGfrYPDISLQaM3u02XpkbhuxZp7nGy3FBG5Qx3d/VHy/AsWsaLsg8KN
RrEXmt7mTVvvf4gIMSvtdR5zdAevzEHg5kyVCdolcDKiZ2mD7w66Mw0p50bCEpVTJIlKa8vGynm2
su+pxhdIubW9w8Kah7x6nE8VvOfYpw0B9CtIDovnnevjdvxwehiYZhHvag/QkRmtPD9+iP5RTvw4
fWI8+cT7PLZMvBL3wiG1s0kpY1DY+1ECd+3OQLedy7HIF2Z3NVkMRPsu18lIbCVqOar7XattuFqM
gersevk+WZmnj4sflFLp+mKc44YHdEi6NKwTCNR9q9HxooMRVyKJxn2yRTDwQVX3xeIb3N2InZia
nOlH6TwnfSJxTZqTaje+rt5FQA1TVf7VBN1DZZJmV4/TAUJuybpb+I1IHsw4O8x/HeQLuiEy80RI
SqAPXe3+wLT6weMFQH6dnMx2Wk6WxcyokbxxNQY/oz2pirl2MFnWIqJDiqs5GKm9VpsAczW/PPn6
wiLAkyLorLS1H8WAOyoau/HENbk0+XkLFuM7qVn/V9iVYoBVuuhhVM041RFHwRzgjmUrtttRNlFU
UCtVpIV2rEIMQepfULHcyeSvToCOfxeVB+mdJ8UQRnGJJlf1p0NGN0kBWw/w74F7fQXMg9HZlHaC
Mif76L1V0te/5qvy3bAsq359xb4VyKsqiEDI6XWC5zolh4mBaFaKyLrbN0CL28bIJx4kR48dkT63
ImAxKRgjgfVDQ7EDJY+pBRWJQkfnSc0PsorvVtZqjlb5TyI7ZUQNQkCcWymGiZFMIhC9VZy+YIzK
u4w04Dq7ZSTiUcbK0f3mTpyLu8Kfw1+1AGFNRuZHDfbHaVX/3XUorSN/fWT7ePvVFMgOqMS8y476
jk+Fn9MQ6QMRGbPv1EoFrXj9T/N09yzXjFZhqCSCrbMFoFUaVA2zZBMj3Ms5lUSiPKzx4912wKM7
fKC2fjwDdp4vpF/d+qIGD/PWn5v2spWakwklkP+sq/ble+lsdhHQHj+UdHpRIuEFDIiwQDOIrfYb
pp+h+c9D3WcIRFT4/6NV9mZV0niqlau8aCXO4mTap/I7So8O7DZoQxvQqTeekXj/QfnQagT4WrKo
ZLpRY4FzDK+85khk/+UZtpUoH+0q1vKVyUUkFtpG9jn2fd1rryHtutUTv2e6/cIdNeRy6DcAMe7G
dNImil8/OZZateckjkfChqF9vA/C0e8PSJQSOvCb1mNxhBwmpnD5szUefY24UR1kzINo0stMXu8r
AbKygmHLBLSedDQenBmSHoqejUVJismdazVxOgYdeWVSR0b3nenoCWONyVCYHAOTkpX616dDg03t
m3337sX05wcnoIZyVgLSKpwO+b3h/JC7MlxJdd5Oz3eL/RkRrboe5vAvugRmZjFBoAmwalxhj1sk
pCxo5CRVy3GQRmR5Zv6jvPW3P6pdeRRSbFC7nqk6jgygrK7pxHAcpEXQlk8izcmzVijD9y3Ok+fq
TSpZ1QDSv9FlVrCZnBvORpedBHg7Ufi8hJmH+ADs2jf8oH2vp1JFOhwyYN13KKsPuhABiXaa1nyt
caq/8ZPMxt0k82qKNKCoU4yVlugGMjhGAv25uypHFThyurtElJuVSy9Goz8Y3jlnKGvuHnvBcIib
KhanBKZsbLiBkdz8H57Yzp3vjZpSOPaLgF4fv53fx6GqFXxGJW4fIZSIn3iV/596sYcJ2MmZU2Yb
AlKE3qDUZyYWE3ttUsIV1YqSo0O1uHXMk2Q0kF+bfOqxZyi3bHP5OnJxsnGOvM2VZ6hGR1atWZTq
wrTO5z36M5M/IbxZfVNpbFQWjJNzkNy/hPfJbqcH8xeiD1P2aeCHRl+Dsh73KGaPcwm1e4uQqRq9
ZfK6ugY+VYa/RECIolPHBhDs+tBxym8749XGBqew7DBYSOHlK52t89gJ3sFxw4/JjY1gt1Z6IAAn
vUzRa0geZqVdYez0R+gVL/w1XXC0oJeXgOAM4miDBL50mZUBW7cOaBy4Zgmmj/0JVfBLWwnR7X+O
25XsR4MoW+3f9HE4ARIB6v+Kor7zn5tpA9OKwHFEh1r9tuNzNolS7+tHxdOvgXGWjVgPpyX/9AZ0
9Gig+sGoQttMICegCFxtrrMee1paDA7UEScERu+1ZKnGbCJ/K6UfyJCGlsBLG2I7LSw188Zew734
CLWNWU6XTiUQQNTGQqJRCj2xejxEZCqAXlS0CVcu+evg3HDnSJegKCccQKpwHqW0EW6RHqfnYxc1
jbGeTaNQNAvzpd8pslMowadvr+CnoZadQZxVXL6RRmXKoVSxgutNcAvwxSeM05HNm1pViCDpVOds
M0RoIP2z7MSJRU8pKSbk/UpI9aVZNfs5RFUFZtDadSbLzoGh062qVUv9BsChrnsPUdHYfQDCtOyC
k9rEOyQ92IUq/2NAc4ISKMpRqo6BXSK+y5j8KLCDeo2enoaNn7LDyifWyyGBJJ+4iNV+selELeT4
d0J8Q/km7AIs8tjnEpTgQq4bFYteOyt8VHsFLtwC8ha5k7x+sKheP3P1qO4JC/3VNT8uXAkkFhyf
u+pkx6mLwV08QR3uNzH+R0zfnWTkvHHjLqJho/DQDyUw6onvUwQJ2y7T8HtFlVgWpIfxpxOKzbtl
7/WPcjbRdXeeFPhxhn4YijoY1q1dFQjTsFwZ+ElksSXscTsfsXKcWDYbO0uwRoBPIdh8TzMQO4lA
XoxLRTFbqivHFDRfihBYNFcNOWH0lyltxxw4eTWcZOKaM5oUzKAXabchS0WIWKk51PReLi76JAD4
rdRoP5bqLfX2JOtTIobbRJsdG7mY7QRzxetTLUSKAl0gxHI8Z77s/k6pLX4NHN8DfWAXIruGxPgT
d1ByeudCgZrcH8Ru6XdsGpwGicC6wr58avmI6Ny/kQh9y++VOVVnZc5Gr0NrY5FnLPRq1eJhzFvz
GxC89ATmrPOtqIDeJ04c99ybTKZTe/bwl8wpIRmCGIkctcpUVJR2JZia1322/83g0KiJKFL4ZTpa
43mUt1wHpK9fpu4ukUat5KT0HZoEwwY1DT0M9r6pH26kTegOqCk1MYCQQSq3bdM9b7YfTEeh1fZa
aTFj8ipC0xrmemfLJ9XvXXbMJZbRRHXx8MbCJHD5pwf0BZA2yBIVanLBKsPWZBhuOwGQoqL1zNwV
rtEbA3YbuLNrooU55pRh24mETWes1r3IKKkaLh4K8zGro8/yQSTBQiv7Ios40ZqlGTMliNWsCAbw
IKMi+LARYlmkb47Orq4yioqKX7X2XBg9HRg34pxAX8ILFAie1qdfNQmcml5nGxtqwFOMFcExNtEN
I5za/L+xG5e3uH2tc+JUPEwt9/qsOCq2gk0amBi5CFZMPC984r6C8xdMS+/rasKBVtI35/zaFGV+
XlxDIQzt7NK0fj961JXtvqxj0vlTLoEhT+tonbaljNkqfPUqozCp8oegduFfyMvBlbfk6PppYnxm
+LFSlbBK+Uhd+3C1RuMd4U0BHQJY/XrHDSBriDQfdkA/871AQ3l62d0wLIPBCX6hnCavAtTEk0WI
wb24Bx+wvFWGXsfrDGnZrFfD/m0AcdlpYEbmQ1IV6fM6JlFeCJ17jojpLL4dcQdvhoovCN+9c4k9
afh8Gvu9XUaqG3kSdS+wNThUfv/pS1BA0Z6LeW2tFQ9/ZVEjIFh5jRF7G+CFlbK330ZB6ZqbG4BW
pAfFIEjpiUUQRRd3PFpXTObdzuOZZcndl0zMTH5GOQKLnQdEG/DXvn3CMAu0P0jLErz5o8q5ttVs
hD+TfSWUGBKL6BPbenoWl0di3UhQWGS2IRtMTM04LyMIr4OWo325hsXnyI2ZzkphKXh2kRfxGPii
BmDroBCBwfj1xGprsm2w9dxM7muQQ00D2+7pk3190Al79ivB2OoFpbxlDNIQD16GrhKkp/b/o5kO
NTIVScWTqxxcW5F4FdHsP9u2K68pt5rvzrMSJjzvudvbFY94lyVaZovdk01iYTNxPkCuwMTSIDLY
3S2OG4VMKka5VGmCn+WKee/1pnjvK+6UPEGv1qIvSzSRQAgmvHMff4DGhQwONgQ/1zUZ4kJLt62Q
ndyKHb61boUlHSr7cWAOuDRSFXSKr/gGEGBndn5hKcjqVI9icWOrWhyxPO4Krll/e5wR8PB9Ucgw
nx65rQplwmxBligFBxum2BQePOIBf2MCTDPtaXQjiL44A3bgxQcjnnlUtuxul6abhIm2OpF+g1jh
ywTH7eusiUfOMlNyG9C2+WIZklfB8TzR8oL/7FpDyDbo1YdKzspgIvy+r9/nLpySXNd+WkOWafGS
OAG6KG63Yvf+8dHBRM3SQom7htG1CYslRcA1lHUcdHkKwWhMQyZHZp282vbn3pZrtMFBwyFd2XT/
d02SpYhV8zHXYNiXQXHEI1M9M4awuCIL2VFMmbQ3m52DKiwEDIMCen0UfllizA9UAFBBG1+phKO4
caXqihns/xvAUwbb5Sfss3DNW0FjZykvDXRFDbHbVdcVm37qpWb0VA5cDcMPlvJk2TOkfetK4QnR
CjQKwGSx1yCNv6qoZxyRZVh4XtYPODuqTg7QPzhwjCLKyfBoWhX34sf420JBb4YjDOS5ZUkYikDN
YJlcgohHzFxUomR/LbPA3xcvD7ZZ6dfIe/8ztrlGA0S6pIIp+J9vd09FXCw9s03nMNLVTT4PrXCs
3kQOFR3x9jCHLSXzHzVOnKU+DWoXJKaM2Lzhs1T69ORn1HehjSJ920MzzlhjwCNy170vV5iQrJOK
N4gS6vdw4jz2kufPlbDp2pgeVWu9Zd9VC0B0gQdDuqBP9I14ioSj7uPlr9ACtYNbvk5A8EAMu/vn
/an3ZgNZNade0HUQHGJMDycx7jfgVv9jehz1MwjXdGKci3ig31VG7mKsSQNmaVp3iIv8zC1sSC56
fhhU+0Anekbl7kYWFaN+Al/e1h32deta9gWyVvXRFY9+7hiNu2t36KheE6k6bHyNaAFE3YL42VVv
8fop09OjkuFmYVJ9gTyteovp1W/uUXeeOGvbliBeQ9vOrOOKMxUv7Wr6Svz4KK8T6dMN0zUeGw8W
P5h51D0ZMacwd24XmTBsb4GCv1amy0ynbClSdX0KzQuWxACtvB26mOgPBQ5tGvt6uypHrlBLIN/x
C7BE3JinSeyi+32lfDqoESw80Mn7mxgTftvR2UOKb8TQ5FEtsTtzQkQGFtI8F5nwhh4ySQm4+yIy
aEOafpR3inQqF8hf4n+pTUPruswlOVkjRSJ3t7vL6ckYVHljNuhEAG/4l8ek1UdGDSb9udFXyXzK
mfPRPwbJ+bIntzUtSZXeA0Pm/SX0co12LvfvT2YDaibcTFT20aLA6B372F44mn/qafNxxHrphRCN
woRa0yV4k5t1yjGvWwn+G7WSs4GThe7ol7lT5Ck3IbDs/lYe5N1Os9hUA8so92yHg02GWw/7FCGQ
2ZN3PZ0NH1tQv+wyxLTfYCKs9kl40D51vzw0qSkFhKBZGSMKP8ljHCcPxk9M1PtHkhNUxJpZqDlV
VWpfZ9X5U4V2dcDtVRudcQ+eKm7B3nWMOzKer290AYh1dEhcua75G63UtzEoy/p3tAF0GKGwCBR0
0dxyy4Vn3OcqDMXPq8+ik/lGUYL0urr0yLjm06eCg1UaLy6TcmDM12XPxMugtxPuqW4UCDevn12I
zTgfpS5le4gId4G1AizhSM/3NDtiu9H7NKad8M3NYYYUsDtoI+7YfzYQGGJs9PqQNHvskeKiitFp
6JHTU+Aj+FMYtqoxgMi3oxoBAiDe5GSm2/bOuaPe2ph0Cx3+W72Y+0VGhDl7s6gseJGBO70RCdxl
eUA7L3fkzNeFsM0jpKcLrll9Cy75ugipo3Lzg2bL+VTk+xWB0SWKbJe1e6Vz8Ys90xvCiud+/vuM
wYX+SnWxXC25iLOWScEcRpWSurnvAQ7dK2DfG92PZhCyr90uFbAIEiyAuc9X9sWjLxORFn1PI6Cu
vfFoRyT2BAIupf7Zz8kBMqd0QvvSD83RYuWnJlSZdjkUvsLjWRzJnXW+TLzUo462ZX0SOlhbIg4K
i/EuNItMDkSpMdCLtTVFgPtmBhEVWhAYHBlYLD9zvinW0c/a8aWwFoGdeyvTBRIRWIn69yiEU9QK
4R5cJAYXQhm5dhAR2skQKWod4g/v+RwrCCNZeVUpkWKCTGQZxVUzme/N/vSq+wC9LtB7iP1iTZkp
vNFoQ+OIS88LLOLb8hLMF/P7vhqhk44UN46rh/NiW0oGqCgp1bF6M/RtSqGw/4ICc4TAh22mJIjF
mNaBRvL7rYCcEJn4N7zO9LRiq5/1o8Z2vuCDC8nzg+Uyi9I4Gct9+6267acWVXAPN7hHlhvV50od
FwHaAhZYYMF41xXsisfvM3VJbl4XbK4m5FhhJCfrNM+sRhCoulTN7TTVeSjuycRPT3nczyf8HPVE
cxdDMYB415KCW+xx5+sIE87xFIxue4wLcS+fm+6gW0upgmCA3gl1A+sVlChtVz+kO+9GFpz8Fl6B
rGahGseqIYcI0V8A33+/RVjxcmONEC7ZRLgBZF0AGPIcadWBLNTgkyFHIOyDM4UlCmTaDyapsQRQ
V0+iAsTshTW94BA+SGHZXITPLKsJ1kO+huDMkB1Vln8UrnCdFn6VK1zKsVwXiYaeQrYBhE6zB8Fd
6RrQujtj0PcL4lhb+8dK10/WJ/0cSwNZUQrP/6jvgQqZg+xWcFAHmV5GyXvQKKz8wohgkTLL3Fdo
CeVXNyrjpx6lqj+W5s2T6v4XSrm7EssgTLfOIEdeINGt0Cm616A/y9YfRs1tUZth/jzfLH1AJu85
AzGANnqyRLyYuSIgdj5GA68TwEnKdyFYl5MCEgMi3v0+piiVwQt7y8IDOcTPcHxwEdHqzHxnaXXa
b1IH6u09Y858Hdjs+4DnG4rm5kw6UMzWeD59M0MFISlqguTFvn02hg5ePPU8ngVukn2Z9pAlpItP
UQRpKoPlCGo/9sR4oTtSUcSC+A8KpPqRRpov4fYsGERV62qVLiDcBYwTzAiNWgprbjXjcv3DILsf
wua7i4iRrcJHzZDsXevFYORA2cjklITsd6Y3pVNceGzvod/aq7EMg7uoDRxhxVhgCrPBxYZAa4Z2
NC89U0PJcPDrcqSDFsLj5tAjff8TsJjro+PIfSsZYc3baH7tGhzFkq89MD6RUIP3EnNVJrV5JOGY
XXcYJwRQjZy2JCCIZ0rYJ+1sr9GJqMGJ8v2dyME6HXJJlkh0GSJPJBxgMwPpMl8ydutxXJxWGRG/
YtCsQGJNnbwcuzQXhMe2ixm8uM9GfQta0rE4q0qHj7BN928KKfeXQl2KJsl2yHuS9kUTLzQz9L5J
wE5O1z9zLLg3hYldPvb/OFGFJ+gXqiZ0uOtjTeJQDYzL1oU5O4kv7zSCA+l2Pd5SKoFN6WglWK2q
t5EVmQSL47xoau17GEDmlkF/et9+BPx7YQfU9pG/y1fUGfv1D9wzD7SLZ1rLMcEkQOMUzM70p3yY
V5bg3GLVLQx5lUbNGFxNkRd5Ua/ej+28WuGlHpYFwbr3g+NuX9fm9q1rpqMoNHYSMbG0QsIeTute
FkPmm4gfhq6CttwNfOL2Qv5GHKptpAr1pVuKwsLyk8m2rXspvUtt1oBTLhS3Zj0oIqqYuxY5Lipn
N9zd6nESoE2la40oyKV6VSQgysdSpgNMKm7UHLJNWkb4jGwmFfJvX7Hs0P6yOJ/uS2Xt0fChsye7
S9wm1VCJprHistMcCIV/PFKjFBhbSo/CFGf8qH3/dnKAgI5B0m4NZe7Yyav9L5Q6oeNHLNKLasGj
AR3n/NtomxTHBEs9jsrbhtXRSPrwDklwYEUWzJHeFCheQZrmxDFkze620r7Jf/gbSQyhm3sCvuoW
LI2yjgt0wmqU42LkkJEvJI9sU9L/mv+/3r5OTlQuf8oJASQ0Y/5MjkTnZ0Y+HyipynUPj2Ig2U8H
ZwrtVQG1gEVtHaIRE/yNVUVgUYhUDrnmwZBXtJwYTrlufLKr0BQ5ZXLJ6Jb5szYfcGhCvlZthrI5
euPdh6xRssM4Lo7pe7Aanc1MA0aQlMSiWUdlHYzIxk8WgqQdaSpgf+f6E48kp8NNqKcqjvkb7OcF
WlRFFdW0lkcJ9xHxmOpP9Cp2tWMSf1GxsbYgvmXWSUzAFACltKev2so8oRnE61PtrV2FV/S67t0a
2O2cZglRsf6/8G/yLYIwfmEnAkWaYHwc+WSd0cs4QbIXsDYkOXLsKUyjwNe+Xk9tP5CJf1mq0bgB
uDBuLxnwJ/f/WmxuN0T/YwOavhogvyK62s0PKxksvPmytGk1jJ4yVzOi5W/kgr6wLvzF8oazUS/F
jkwIu6ySjFHkiox+XcOA7/N6L182pStmhV7i1sTqFe1M70teRrqsLeMYKzW1m1qsqK0NCnKdiESX
HuOC+rdpQFcthJ9u//+MoiS/93niN92FH3y6n7VMStwjxnb7HOaH+gmkPsChmGnDZJcJZ2gMz8vH
TKlqGn7bz1koZFbDIb3XA+xBmjF2NtlSbPGO9AOeBIIE0qXJ5Ic2WUkyiGTYxzOkNvlY7Z8wis/R
a+ap0uX9s7aejwcFcM7+qz/gnMHvMVATiIIJwSNPWyA4WACkbbspMpRqoKatsk2i9tOhG4CQ2tQA
un3VRNA9DJU2ev8elTCsXQ8PVHCEYqcr3HQBW/+IaL7e+O6U4bLCBrLIkUxYP6hmjXxdhgZ74RTH
pXmqD7BiiQkXYAcmFOGF/4Hgl1lJpchQ/2iBhE1BCgBGM2Co6nxVsGO/zfCuUL3T9GgIARPoCCDo
GfFzHAPaRHQjwX8y0IKLSrtm6Ondnxd61gftd1uJnDr0fPLYEzghPvlc4vwWVgNhFZ2VtLJkuOYh
O0rwfBo9i2WqxpVKv+ryDyhlKgkdbIkOfKzBhtmdH+l1h19XCLOh2ATlauapZeMu8XDWYlg7ZZm4
iZ9Lbm4cB2ouozu2BLfzQ7UATSBnzx/l/iput+jdLk1OJ2ggxOHLoHOhS4KsZAlicZS9icpgjjdS
eenZxFrO69RDwBOPZ9QLIu8OdcHtE+ZHIgaRqtTurod38mwRt3szfFYJMegiVXUoVEnOsDMFk5Vm
RWOWYr8Xa2S8oeYXrRkAAmTPeM7J8xNfa9+72r6qTTtY/v+A3e67Co7bWcj1nksgTJONXJ15dmCo
CGyw6GRJf9HZWZBOHlcrefCFcKNYZGdhModZAxki30I4G4xiC2lRhpskxQVTbWSKUj8tHj8rVYS0
sZIZjPkIcgMjbFsRWSJGPKcdezysNgCojDlcF5VG2Vwdm9e7eD+Isa6sTO/uafMasqSZBWHDZDpW
n1OEBGTLTaEh6rI3ufb44IaVjH0ECD/suxp+KQbYJ93JQK09bypz79TIP+dW/Abio7Kx1n1XL/df
8ucfKda//Pk3QeqR2mTx1XVtp1sAwgW3lQEF4My9V1ZRf453D90gQ9WbxbPNz2IPisJ7z1jC1idD
NSKktHdQH/hDmN3DAsUSSq0hwJkXLkzgqt6n1IJXjbP89Loh+bnLG7kOvR4rv1KT61Qkik7sVKtv
gWyYeAUUloDiul2j3GQmoMPNbrz5RORr4EnuSi3WPLlPekyQ9IOFJRqZmI16Pzq2xYu0bIlgSKd0
RW2ovlpEBnn95mVj1yAliUXTT/SskOITuA5GBNO5w8Nv9IauPs3UevzuxEeIH5gUI+g7NM9nwFdo
B+bus8OtwfvNGQcYHIaXl7joHvYE9TSZd16PJellPsF+odhOcmAHYAQpLLTILtBc7xnAiaXgUoY1
9MHViHGOgZ5I18yXXf2Wr7zr4hyjOURZXwvcqNxqBC89gpeLQ+lFR4lGfhbMEC5Hq9A3drBJ6YRV
mKB51prElT56Sxkq0Uza9gZMTUrCPd70PWqR9/Sctnb0DbA/QWnuX+YsX3r2JIvTbf7GoQwheZvy
52d2MnMKD4CCHL5BQVtCIElWlz3xr7VFG5y/xojeqvoO/pDznxLcO3OQUQX1D/yTr+5UGb9Jvi/b
l+eF97GKG2XxsyIfuO/cpOrJgItTNoxcqy5+u8K5PfrzbT8DKhFyZAHJ6X9MKn8Pue6d2TDIyOtv
TQkC32n9Go8TsRAqV00OZBPWiwVjeBsY9cgUybjjoHcKVHjym5EAz9qvK+fHOS7L/F6tmKEWLZmF
TyquiF2LHSxugdICs9JZimPCNqkHH59nUhj5umw0GEZESkylFajaIyDn0Ynp6agbxdFxa++gTu0h
C6d6JyZFWnuYKM0VkI1iZ47StIoGXUOHOmdCbz1Jcu4OvNTywi/lIcEYSUPoZ5SJPmpi07ZGn1KE
XNC7qSeG38KmUv0hNLPRy/xCxvXMoRZbJzlFnKxfhq1Cwkuh9+zKwUlAb7nojbqBX8daFMHn0+5h
VcLgSTByTjODWKq7BBR6ovGgdku+b15XI1S+PBQSu6ggb8toec3QxLLZRJiNbMC7HE4tmI/fWQGF
4vikoxBUUC3mWbOp5eTY88Ct3qpMNuQkVh8a0jQKujxx+SFw+QKdnKIZMiLEYILNs0vuUFZytpIn
LaMJ3jBmfvuzS03NCZUrpebyQIn7lrxstXSxzx0xt6fTcReFqlI/AFz79fbr1YrHd2yhtvXqqsnH
mjjbwxlO3+JYKsFPtEU637gvmHJ91mTdQNyDRQrkchDSIoTZBp0Q8X/1Ssz2JhuZPz/t8MiBpygD
fQl/3B/BBENCRBUrWVptlnWi/JWGV5jeOaog1uUjVCQtzX29as/w1Jq3cxX7cYP0rNIwgNuwxR0I
HNtzugSIb+fKc0WVOF6qPOEI5pn01hs7k2SoCZMiaspAdsWK5Co8UThg5BZ6JZ9WoIlp7iYDdcSi
6ldOfcgagA6WFBjmsu0FoP7EnDZQZ17B2iAQPJgm3GthXB7yTNysSFRMIKm/4+Vj18TJ20INSenZ
ycpvJbKi663cN44hsEbvaI2dxWU6wOHcRCue+VDa8Z7ALZ2Tqj4nr1xYkB2HxlLBkjzLh1vT7Z4n
MPEXDh7YkBHnBk9WWsr/uWblew3rHejomRLLimlTExBIY9KpBJngL7sejQi7X3Eo0iYHRCv23fx+
OeW2ulj/pm5CQ6wEm4v1nYXNKLgQgwAfJdd1f9zV1gRXDHDJn6MhgPRQJqGH2qb8Tx0Avev5IQeC
+KqUZ9TDN0U6Nimsn0WLOqjJujuV5TlI7rzQZCBBfYNu3rMYPiZkxvAnCWlrfN5h3dKZcZGXWddv
QYMaLY3FdPWSCN4DSLqrtoedLi5P74UgP9K3PziHUG1L9EtD+GilUdObLmlJUe5RMe6KXyf1JcZP
bROxTXYVBKer0nghfQAA52z2Ml28R7Cs3dsXk3DpscfbAklINJNPbDDWrjFpbP8jCn8WbKou/att
mCCXgItiwZS77lmjWRWzN4fH43gbFmfoC0UsfAk9YPYOuzFIYqbY+rGzfTT/Sezy+gw7p5K+aFOb
UqLc/k9s4Y0wclArqaFfZN/0zYzCAeKzQeSMH610e83k14WWaBRcWZ3suEK+gnIzJgcd358VByNg
4YzqfwcWyRip6eGQ2+j+JJjsxMJp1nalGpvl06wlmQdrqkB6zUlPsdh2P8nvqsZyDB8yyYFpoP1V
nTqfrRTG5drne3ERMzHcrxHMB9KkItx5wb3Swx20d2VyPQrbqQV7d3x51jRQgmtbcq5/Zv2CbijT
jttDD+N9eBMts6awXQJCXkiSpKGnGPsC2kujBpTz4Dqhf2gry/sAq70OYE7f8qvq+WcKqmkztOg3
r078tzzGFjSQQ8POC6w6NgKmGCuxhvVh3BaRmsqQRcr6Am/LAbr6o6FexktYjhkMVqmcht1c5kDn
4nWGAz5YsmFVX91GBN0OmyHbbil/jSC+fpQ9G1d97GMOzFno4+GLetjbbdaeGwsVlcsPk0RMcvGE
E9Y/PcxbhEgQYkCKj+/jryT8bGxsbs+/kK9FDyNSEQtsuU+2o4CCXFaFZpx4IYEKKinFjPB4CjW8
+HpR9yi3Lq0oUmyg7gPGsA4kMfIb3WnHiXdzVYenGDcV2CcN8TrIfSY5VQ8jnWo6riNmiYS1mwN2
AbjL1TmK1ySbwhQlOT3u+L6wShL8M7clurrJ3hwg89dlUe4evA1AHbwapvRmpYlgLlnQpxGGAvfW
CTUzD2B2UAzFEnlN/gKLxGcvPZtrBf2Nee3F+xlS9Kswjj5PS3ol/sjxxlJvRjmN8DXGHdfVjfeu
pxasamEiIFECI72ZtBOlKF9ecAbgHwXDA2on9g5rHx0jbq7Ha8jJkJb/6nBONMcRgqVhR/874WAh
RUDzOMKqO8r3gik2T3zBSSEXtkBGpowFp4wAXT7Ob4imgjlx39I4I0gUBefaC602nZXIWlEWcpMe
IOfNtc9yXe2wVvUtCjWDnwEPHcIzN7fCBfov06yFssIFNfWPZUZyT6gM7GOI83qy3GaHD0+Z4Hzv
uJ0SvMM1L7jz+ywiX4mg5AYdk2PY84RifxjLHXlGgUjEeCcmwwTr0sb3orVovYqCg2p1yldKGs0i
GPVPYWifvSFJyIrlbHoDMwWH7dfnoSLu2a488YYY6fZobOEYPjFzRakc4TciRuIdhkYT6e5Ne59T
STN0xlnVjs02Z7iq1Bv9ZluHyKbc/bxH73AGNNMYyCmHzr6+2jFjFimG8iFsNOEPyEo8QuZpymyX
3REGJVu36WzLB1AiBi409NB7q1kbAIa9UKZwn3zfwWIweDlAVZgtriLdKIMF3Uv8ufOmQqlEkoEJ
EqUm/JmTqWlI8k8BhZ9Xads4r4dNsvPH3QapKEjdqjEPLxfs3ugSYvZkQ/Oe/WMtoA9BIb4SQu6N
su5pIFH9Scfh5tGatrfuCW+w6FbXwUhe3uBPGksFvYI917K9zRiuk3KUO+Y9rkvLZYehVKD4b3Ym
Rjg2XwfBegiKSQqvJdvd+9lX5Spa9OxWfYxGV08huKe7J2OQ2KH/+SgLudCKZTpdUUhHoaPv6KpM
sKpjC+8wR9KoOCVQCUl/5ad5PaGi0FD+cpoCWAt9i4fJa9xF10HIDl6A/FlHaNhizn4dlfzkpOrf
Fp5ghc4whHv9XBvSzbDhbcjPlk5NzMi7YIiuy/wdlc0ycRX7mQ5Z56FD7pCe0AK3w74ZHnUOztCX
snzJxQUurE4xxhyM30iCLX8uC1MRx94rfe/qvui/tJZft9mCMRU9Z+iCxKbpvKNbDsrC5q4xIn0W
MtgLl+dbKmaRpKU4csnwcOIOzraknUl5hwnSX5crshhTjbD0Lm5ZUTxicVHvZJZjL3lSCrkF8pXi
01QlnY3Fk/h4emg+MNh1TDbm6bEYSrx6ty4SxKEuR2/0KdepStLxI8SgChVRWVFKrTW1JKOPLmzp
Yj+n4b1jGo+QBBKySR9/5vrJazAEXtZHg9yIsarQrbMRTuSC1QsH2CUEXNpNrxeYsvVKY+f0PHdr
vtlVCNNmiQxYWjWIGNbzXowBIJekGfeAyV/eyMNarf609t0gAzu7VTc+/Ny39E2u00D3mc8Dn7Nz
WdCU7ckoq9CQWB7EZ7w8euJKyqTbKk57zx8JeHTbIYaAzWlAvEYYQvJ6yhQCGEy82YYvcx+KeL43
uqD1ihaZ7iso/i6YRvfy6lzNQ+OfL6t7aGsxyctHEm0w1T0N56Q32Gf4wMpgoeGRwK2TB4endMlq
VA3coNm/s9R0fG8xX6rTVADlp3FVh3dlzamS3dA6Xq140Xip40Bw8NwjuMEghOzqe4EcOSCqj78d
gx2EKfBk/n3ZjzKoyoeqckkL8b9CqJWw8tbZA89b2rR4nA+ANvMOznHcwtWaI7Bdg/M13/vFQxXl
jeAwIHZEUaiAint+aQoapOEiKFNYsgMN0Vg6JoySv19J5A/t31GTsO2V6OEtzfER8P0mwP5Z0ehr
TK5eCLcxNYscbJSTQ3S8vi0FNDnqM75XK4tPTsaz9VXHTIN9jHkPc1T577+ib/jb/pLRVKkp8bAx
MgnZvMcpoPUf43nfZ9ej7i0aWUTofq7QRdM6M9eeErYK5/eHZ+++okmP8/c16pGxJq8UDUfVmxRF
ytIXkXRWNl4+0Pd311/Bn8KnPBj59JROjR7R4XI1ou2FRc3wjdvWG9eGMAPOAFadDe1gEV1eSJuR
ecmob/VQVZIpGBrceaqnTV5rfL7jQLPQ/mFwhV/vOfO2Q0SBr5mIIVi+ZhqSj8G6cngYBEtSZOZG
yF1+83vCVv4XUYYUdift9USFHjEqyZUFLz5X9TABwWBzA5MMtZNZ2V0YViW9I3e/RVbDF7ORxyb5
FT/XuPceFj8FEcajOaLRVA8bwaJmOgY6wutTBQKm03u8MM6v7uCaMg0+qZOB0wwljgPyXdwd/JfC
60SpMPZPLgQ0+yqY6HJPwHqHSj938XWEKd00+2mWGIisCLaovb/8ClZRu6M2sh18G9oOkMsouSuy
qBiex1RNJwoKYBc4rVfV6UzLnyyY0bZsx/fcf6N933QvldnA71epb0ir2j04XB4ff+CjMrcNZI3V
CNLvTq1YB2WHy0M1JoBctQpslbxjVBr7ds/4ko0mTSkNegeCYrEix75PIth5rTedrhLYLbVSl41m
Jy/uEdbM+HFgkPhiz3xVq5qiWJTr6hG8vglttoIQpaF8kt161OLcyEUZNlL9Pbb6abX7V5Eycc/V
2fawgx+15XeWbaW0MaVaIdEqEwD3GdkkiXpVA2pa5undpGaj6+FpEX/ouRIrn7ZXAttMfQiNaVfp
Q5XXKx0CB+J7YUMmK5c5Dvr6YGslLFRCZ5A5yPN0ncNeOLzxhMbEFal4/+Z6hLsoZQ4YbByWuUpl
udItBaIl0Ff4tfBPBxoMnSmoUU2f5SYQCYyrzyzPru8JhGTcXnkPmrAYb7kHEYKP0qt+Msl2gjyu
mn86rrIopttIwZsJFWmnGOikKKM/hdiX937PrGehGT/SQ8SRvdyZ7MigMtqo8xruOzbxhnb4T3mn
k1Gk3tfUAbUUwf2pao6CBr4slOHm8tPHFt3GxdetLbyn+1SWHO1PLbl1xQlO1xN7aMmu5/arWbYc
Y9COX2efqoNLFt0pKtdaxwYgtD3UdC++NhZhylYIRz544GHPyKG7GCNrClN+RtuFGXFQcSjZvkNf
Vf43I5QmDnC+lzywyPiwdMgeZ69Ywtas0m5kItjVtbRv/ercdHxFa/imjsP3gZPPBHv9rwYoCBe1
nvOe8yWAW8kLOWH1NytV6vjtvbnuoI1Xdt4MDOIczAr2RBYuwVNHlGhKNud8xI3sYtK+iYeAc3nc
FPkg5w0hU/bPOytJ3uCC/hUizW9zCHpdteG4CyPCsPFeyTlyHRl1p7QOClCC3D3QPawbNBINw7Oy
PIj6IkbdicdjCN3XHKf/ntkNu9pxihN3QsNzpQncFmTvmB6xSbole0FXqYSLlfs5eUus5TBaScE3
ACABtmy4IAjd+UOtMO1yd1y5IGU0cLhtJyl2rzI9mFWRMI/zDN/SQ4Pn/OA/Qk8tGOjvIZH07psr
eqxD2CAihl5Z1a5adm7L/ksh1LSD9gWvwbQQJSIDTB0G23B5QzCHxCxIIiNbJKnhPCSj33WdnmL6
cvvBLKHp3EmrxIxtjG7JRuaJ1M/odgsOjjhSYIWOQ88yfzcZ5tM+/ArcO5L4K7M8jlwIZZCVpmJ5
p/B//C8Zoxyj4hjWwKxtLEV30e92mHv9piw/NEB1biClMAoUp1wPk2snsqsrxPOJg7UHZUlKpiU+
Wkjhe2sakZIIX+sOsrcJkw4ViYWf96OUKCdBdGLzVGRKzMquzOcix9W/4HchnIuCCTPqh2HyIHFT
hz9/5fv3xkM7a4qQ5MGmKmaMU75FNVG99UTkrfCmJZ7RhHcv14ZIZYFLE9a1IUGAMzUY0CCJn/BL
1Shg3ZU2Vcm/QgFUv90Bgjk+DByZsEVt6p7HoDwjJtrncuOEqUdU/tCcjYUpFNIfIUFepzfmjwQn
1SA7z1wVvtsmxvcBhmJ0dT9RsZrh95XRwREunmfsH6avY95iOLvmEEr1szNTS0XMazGJag1O4RlD
5hdP6sjeYMsJ2uwtgpJH4zR3U/XX3Q8KNuSlPi2jmTNIAuYsOMVYn+9EGr8krkUcQ1a9q6+LeiCm
ZNii7irhpU5jlK9WE1bhPtJrPBoArUMeGhdurG+f9vuG6ZAyJ7JU+DRDo6hS60K+ttCJi/9OWtGB
EFW1X/nxU/3vhd8FJEHV32OwpErnsjZ0qHh5a/1DW7UZ5vMEfKx40RI3Agqe8zdG7kGZyS5D/axB
juwnyUaDrt2vJXfvga7Uge6pi5sZbc/oOV7/5qTWsQdJZvlevAzT8XoXZwdl+xhr3wnyiCHFC3Eo
PLv5xOMwz31sfdtncnfk0zWx3smvidUbNbnlKilQSJvueZcr4PjQ2obpqfkhSuJEmNkLBsx9Nzg2
0zfuHD/cJ0Q7+rdnXLHreHQR/kIqXGy8eEMcnsxoRMcu0lyzGY9P0+U50Bk3zGKp1in2OHyo2Uix
FY1OD/Jk0vxgvY5kDizkLKpihJPQ3Foms1cgwJTCR6DJ/EjE/jJpjBmBBl+ujahT30S7fsiW2oUT
t/9++0YoVfLQMaiTA3uapbmn3HHCCfncS+A4BnYMAszVz93VDnTMvrJov8re8qsO7GFwUBkSPTy7
vpr3EGhVwT3d1UyYYtQgmVoEzvI/b3v6IFHClZtUsxe4op0rkU/c+dW6D+Lby1iFU0tIN4H0cgoZ
3wNgvy7UwhQjzxyH+++bo8RgUNG7fyT33vMOxp7ToEQQypKBMAU48fQP7MBAx1368Eeaio7XFQAy
OQKnO/KdVpwkJSlcMiW3JLLU0mjESF6r6fM0j73xg/Mk2iOOHR9wRqjbd9cEjk3nGKlhe2uKNAo1
ADTkrvNqYc/B4FoXyKeiHFo9LRd4DIaE4SpEOFaC5xjmKbWC+0CgCvhMJwdhbid81fvZnrX3nMXK
sB9IfCmP0ewuEP5jLOSVOBXRUeIxZJI3pNseKVwUFHpZXpbs2keOOE2jp9wNJfPI6Bhfn0MCJUxr
w4p1LTuWRCk9IDR3ZsVYi2Ts9UNtCkGIiB+zE7lDHcQeSlvVJcpmmm8CiXrC1NsGfcw4Jxmskv/A
iT1O7I+ulHimudODkopJVB2KtqqVzrB2H9JGfogD0HjWDhLYOCgoqaXMcFy7r91nC5EMjxwmV67h
IPYq9J72EwZgT/mxbq6zYsDv7DCwHn2bFeURFWY1wsoHFa4r7MMt0J7fXHK32U0N97NkMcCEYrfZ
YjsWtQGpK6zrIzS2emdJXP3fJEYR7vybtOPDX4wcXwL1WALdhdSr6z7Ly+ICj6kI01zgiPp7gFHH
j986YaOXZv5cTdshy2fxunAY2laMuJkxHSpKjg/OcE4ipMXDGZsKZIPcbVg0qibT1iWr8oWKAC4n
lDIdM+yPiQrOwkUTNgTKvFn+9diXZs6CyqkQPJviPnMvjg2r1aexUfruTrfDykJLpKpL/52EwsDS
pKqepjakDvi0KDgNxH5EsnZmC9iYD/XXt57mgSmBiyCfkj5wUZt+sw4i/me3sVf+h4mCqBBxyqwV
1gd/syrV3HUwyoub0nCeVp6KkvfFSYdZN353NlYdzBbPpBV4YUg6VOcO3EbRa0idA9Q6Z95fhTDP
0FJ8cLFRnXdNvss7HVN+Y7FUCZHPJOYtVEacx9an4ExHvwR6UnaI/8W6Wu+BctzcxmQoBuNrRpYl
851OgRILjEOEqmzsv94hP77ME8k80DUnoqPBJo/+kIKndWdvs474Bz2BAm2iYzkgvWq725yLLuAV
rk8yNnoJnLQPITwRNrrSrL4RPJr1f641ooxTtZA0guAo/Y0w69iMU+5HGBhFzHLeLsrngCq4nZRV
RFjO84WIbc/+uiUz40xxsmJcg/fYFRz+EwM9twy/tlEBghx8TgvKpig0YwAFIaQ6QLpXG6YaFxAu
TX3pmP/MClPUqDiWX2bquIAvSyv4qu8G03UxGTQEO8W/ZSGww7Nx2bQWX7J/x1SMOencrHoimoJS
PYZqRnr80osA+Mh4VZAJHNA5hWytn7+VzECV4A4tc1X6l4lhfTbQ+5a8+8Hch58PMPi8DDQ/XOFu
HkzD5372djIdMflMWjrGtzR7zVMX7yuuD+zjag3SwnScubqb2Qxh4Pp3RL7QMjG6QEbsXPohIiwl
iqG6HwDlNlzQ/9Y42DoUK96S67bIhPNYH8w9meaa99N6aRxGWJ6xnSpYRVXTyumc8Fd326Q25+G2
b6lIHCQeGWOyPatqz7ORRdQhl0SzV01YDGP+0Cxe/g2t6TkJap0EFmf4eW/UwGlxd/MTzZ+KqZN1
DR9rM6Rj+rsPDXsUKwOXN4gJ2TT1gXGDPiT+YRxuJPXL62BD+TbtK83k56zNk/z4rf114xRaj8Ie
I3LWpMRsrae4Ekw3Baf2aRsIn7iwL/l6pa8pK7lqyvUr5xZ+5qPj8n4Nxc/AXzJnnDPxprViuRFV
IeXA411BHFqis1sC6BpsbE9BuvxxkCiQ8ApCO+2G2jOlISDPXeMlkq2Wr5SQ/flpt4Ize+505cjV
KpwA+0CUt3GG4tdjH+8z7BBs+Qxr6lmHV6hgsWnLn3M6kNfljFtu1VW7NY8S4WHobyQM7Xmv6n5n
vzXq6WfgryJXQ7IT5+0MOAo//DnzX9tofJylObRTud5rM6wv3T3nyIcdtaTWx0roMP+TwqkPENWI
X+19/o/6kHrGS8JMem3DHrd9f4haCcKH5z7yeLhD54AFCgSMqDLrry7Q9jq4iSVnxBIHMWN3iF9T
aknkL+Zms35da/w7e/0An3M4znbz+dmDYOQsVioLujQCkrK4QtJKIg6IRxGU61bGCB6smN2UIxdj
DQyeyInp4I90ZkS4AZPBXzIT7EFQhdMjMhGm1vW1WvUUtg5HZ4e3fKdQuI7c5xmgwundTTD61jVU
9DrRIJ9YPyQpXXdDEZfWjwz1+a4QnnfKuUg/CetIyEkv2SofEs43k1VCpQC9MULyTr3GJ7uT99QR
aj2+6NYi9Hq7lalC9TVWc2rrf1Jk1Efp2Ba13dhtr+kaO0lRiqq20s4DFuIYRt5RoRi5PKizWCMe
kOIu/Ba+i9iZW2iojt4U/pM25LR0OlWSgU1PBc1bPk5/w0zSchZySJROUS7ojwZcnQxjaPp0/fcM
BAwxO84UCDy1YjX1BRA6bh1JNQs+pFHUR6UhWJ3LtyJHtrjWQDU6peqWNsaBN66eXnBKpQ612I4A
c8cW8S/C/+/TmuTVsdjsBZWPrRLbKyHJygykzG+g45Fd5mb1RSWQ6wD3lejYbcb4rKvrngY75OjE
Au8fb+p705G9P0eSe8WUBdXFbN35bNpdXYRBpO5qqntZ1zvfh3GXWLhtmtSv/LSGPGhIrVhSgmmt
xjlSpaEfHvHzBlRVBT/Cbsi7V/d9AgiEXEfxEzebCPwUVWjqck7nIC+1G2ZKX2UpJGgSBq1xxNFn
jbF2YHb7M+TpJuC49qsyUfvPgLDK9RvpG0HTBQvB4caNkb6nygKl4EvgYGnFJoF4aUvOSyobgbGn
4xxDBZz19qm1mM9L345SMP4e39pGS+qwC+tSq9alZTij/GeRBqY8ZFxtlb9EK2EaIoekI+De0Po+
L0S7M/pGa45Jvyg8LsfJmcs3G3wbdoknR+N3oKT6HAMKhmyYOuHshQEO+MhtMB+HPSkfCV1gSGKg
FMLZDit+ejBOVHnEvpe6h7Bgr6TzYWD3PdJ1UWkcWA0OFTj27NxepCRIG/jDhAqHBZGGJsrdByf6
D3LYL8p9vzCBlYA4cOLKYO5eiIP2cJvHMJoXHx5rXcPNbmQ8i04wSD9OepQYO6fTv2vwxQHin2pM
6YwDOfuAtVgQFyNj8SdaUKgtgE+abbJgnL7I4Lo03L8ETjg66Br9odYZKJ1mBLJH9HqvmpHU39dR
0FscrgF1lMbhChPYv9cwlXf7OcUA2E/VVT2zjD8X1WEGSwApfH9bd8jmK6H4pfP1xNe19tM3/LjV
u92NUYnIreI/bY64HxrEETAEipeUJ9vMkqB3HznPyUevRaKX9vsXqSXpTrhAZQaTIcnG0W9pXYlZ
kNGuIFYXpLUbi+GM2dyecDgpevtyH3xFTSiwAGUm2IcJwKrFXQ8+iomCany2dxrAz6NSIMoHfpFz
smEqKlB9R5ZpoRdWdHfFgTJ9Bgnd2ALI3eZqE5pAwpHGUZ1nqFDKfZtZV+Hlg0g5qjP9p/if+r2L
Er9dbUgC9Tl4Hxn+NJT3fH9ndsoC55j1UpVbO52p8AmGwJTSQGpG5ccCkCikwEpN8/5Y+Fu4a/Di
HbWqSy24yLmdmP3t/b+oR9t5ZoqRzMCjRgwBd9i+wt+kEKBVfkX2hJVcspT3yh+J4oxMob4gXABE
IqhXC9UGS1ycfNPtLOdTJeIMQspue0vUAZpuN6I3Aq+/iJZxYq5Ddt42+ilsQ2wOs9rCmNt9fL5h
Y6Kk38FYR9kDvXoSlH/lIQWEgeMt4iLOcRPhjI62xRoMRHaD/zEIZ26ZzyXJETp4X8xrkyMQCcfd
RF/ZS7Lt7xrnz3uAY0SZoV5ayWbUSLLGwHNKC29vM0ZXYLaCa1hEyXEjegxZNNwO4qhndG93Um5B
xM6jbSkc+xS8jMBZYgXWt/pSNIJyuLobe+tLREmKZGVGm4QGfW+ji1fOKzyQ6avjHVBq8izPfe1N
+q/6NcRme0e0/GhocrdhNDHvD7RAna3M8jd68NCoVVrZ6ZMS2yjJ2mBbCG/EsLrq7dtX+TgORGvY
8csXTzHL58iew5ZLHoSk4bqsHEr2yLRN47SblsYNuhFGsgDnITQMswYRgE/LIDMwSrWqaUYXulZ9
792Z1ebHW/W97cOr8J/nttw58r38x3oIkUN9ZN21P1gXLgFD5CYCNyRp3zMPPRAtppRPdWY+UhKS
a8+XUt5AKjAELfgfGlkVfVJFCzdBrahhJG6GQzRfc7JXezQcRjT5FEF+qGy4uqm2uHqzT9ew1r90
3F1aArwhn6P06r7T//fDI7zeL8c9/HLpjZvoPaxDxc03NQSz1YU4x1nGWv1XdBtdGQ15cwhalcsA
X4GhzLJpoJaf5UZPwn0V6v+k4DNaAPS0x3HyfP/w3qzus7ayfrYz+kZ+WflZTpwdkP+ZYcZjalia
XKg1fM6iecHXMsQf7bdo3WSrpdd5AcmAHkFdGf53i+MHadwjQGnMp2ogeyQ4IIOHuUiuog9ERK/2
L/jh4FaaGfkAQUVXcjg6OL4DqX/H6nO7Rotp7+3zTG70DPYmOLg7UPnmeUYvSRkvwGxZ+1bLLXHN
5IpYKyk3p6SKJ/nmPaZeOa1q2j7O4eDwHqhHQQMx9uhsaYqnJzAazFD4WFothUCiixpQahk9/Dh4
NTLVnfjUsDljnVRvaNQ9y6q9CFc3+zIYq734jNZNVbjHIo7ByumqQtsv3ISM4t5fbmf2uxXN+ukL
XEkDqg9PllhkjkwHcjEMoOpQDhfTiYTjDV6pGhKCrXW7yyGXhzOB7WVRIk/P/iCAwOW09hC0SZl5
VFnHsGzm4EIqNvzECNq2/hlK6CfeaIH2fcrS4FfjvHZfc42zfldsmupOTCdU9aj4qXS7n/KJi/1l
viOyWjLtftwBSd3KG4OvDCMQqdF0RymkF6SixgdKIq3cixUKq7pAptkJR+iX/UEPwfOibK1XPh2n
GW0an1GWvo7fm2UkkgorZqoOUsksunAlLAsQ5fTGRX6IvFjvYPrl0Cpj8ZkBo4oQ8cLlGayhZHTQ
UIwlyUWjJCGLysmADqLf6vwLUwUgnKW9NDY7oHAuu76JQ+J3ME+vm7mywRFQieKUSqroSrulnwVA
l886dQIqx6/Q1YT3wK09Irvg4IW0WW0KcqpwErfIdXgxphgdmiuzEjjJ447inpFlQ56XZ0CyChJT
tnn0rFpxNpGHZzHvp5DmXt0/NHDAEgtJpm9eAmBTNert2zVCsVwCnp3dE8DEfGB0d7jlDijwxgfy
NDZ0pEawtK3bRTOQ5sJEWdiTM9jn96iMRQXQRE9/BTP/8SG19phRruSqQ9Q3FIJt+kE25xrTIp66
8D5G8uQIoRosnbjBXs0JuCrt3ZXu6yr2Lz6eANtISqUetd8uf7K9pPYegAJ89Ph5yQ1cyiXR0+t6
pbffl73tRRXVKAtf+e5w91LGBRYtD6guk3UxITM6xsFm9znU+608wdKLt9MpUxgayAMruFczV08F
2aKrGSEvFBdfRcC6AsMKdA8KbnjIKltoUN3heaORmd4x+892zDG4RQ7YJ9djonEUCnW1YeaO858r
NGnG594p4mTbABfLg7K2oedMrOZakM52pF0WH86Zf7zO+m+l6+bfYJrsS1xUjZ5RiIeH9xwRNQOa
vE0Of6No7V5RbMT4aPyAIrrzcHBtKK3KMpLCaitrsJbln+DeG6fiNtvUBd5gF6UW77UQ5ZuvKgrC
YjOfqbFM791ulYPQjU1EcCnqY2eoYZLt3xT3IcaZXeh8eU5h30/w7Cbp0ofLGNfGD/LGxZay+oNc
JhNmHROzq2FUN2cFcg6Teg316c/VuxSxobJRa0q98l7qdA3x249KnMM+xr4m6v0KZhqXHLSSZ/Dy
+2ynKxBNARSrfbuAbfYWXpcgWDKWTJ+zB+TF27asRFpNqRO7aPiAqR7qDm+sUW6eI/gnuwZbz8ks
n81jH6Jb2WisetOiecAohZS1tq7si4lCK24FifpkmdGyiOgstdV32/CEGMvWrmMKhazz6cZGfP+U
UdCogI8r3ovLaBItVoTv8kwD0J2P9jX2nERJc9mRwk+qrT+LaVqUPOadOJtuvrztrZP7Thz1qVkk
UjtItkfHeqh8QPd1VPhUxJh+S7qIIislFeGVQWd48aIUvanV8p3azPBWMFTe5Om7epH2M/TEh2ZV
7uHHX6y9CvrfHga26uahD6o/sEzqZ4non3Dxa8M3Ekqmhv/iAhMuuS8jEGXbzpQggISTY/krYYaK
8DyRJU9ZjyRlI2vB5IEmMALN0m9IUrmR3xy7Rin3RtK9HVb5+z7RzvZLaadnKla+Lr5IUbdJhUKZ
g0C3Ukf4nDixquqDTx+xNW+myrJ4U1l9WPQikqrHQTTZO/QxkC3fcRwaZFT0TScThgT3aF8UmOn8
FUC+7CRNzrQkWIkovamrKMeESTWkDXK1tp+0Z3AYT+j6O5mI/Do8yg0MV1L0XVIYtG4Ul7kCzhMS
CCWojwBTI7j72ngfocEokYm0vWf/BMCIDA9KzQyFl7IzlXbh6awVCoHEskQrEMx/JPgmwLjxBVEN
t81LBHF4uTMVNxxTOznYfHre6AfLJmfGwLZg73ddbMszG77qhP22pQi9k03aRJnMUD2hPU1jQ/zR
q+FVwgDXIXiX8Hs7/lwcj6/IDeIzrTqguDN43WVBdIBW8yesl8V42oSQPLeSPFrTUFM5wFKdqwg3
phB7FtkHE+DiRP3wdxPmIl7fvh0g1QbZ58w1l3Q+recPO4JW9cAH24JSm/4yzOrZpt5HOrpnfedb
dej6bDAEMk7X5YYo2DRDpxpjjX1e5NIMKLjt0l5Gq64uqNHNE78e71O4AfbCWx9Cd5mSohq2rgoD
RMdeCHk/uY/TN72IYq/zllcLX10F5t4+OxD+hI2vLitw/se63OX/AtLhmo0aasft8b1vYLVg74MR
EGaOeV0ZrDcNK/PwwYNV7Liys+SzEbu7PFgapikdsMQtGFpXTcR+s7nzvkR1FlyMPeTNljwa8A+V
S5SqtTbt3abgtww44MrLVbwNcQe5BiQ42ak9326erWuX2ZUUVJ6tSa/HtsR0ZM0ZN3k/aF1GjOZy
dzk74Ymhmo2jEaRmjQmZ2m5ZrqZxfeksFxsDSNXpkSvwG+9dwGgqcBorV7GSzEzBnwhL3ej74OF1
1u3kQEhWeP+pdbGj7l039aABpKzdqBa0lPwP2cPkO3b5TjmaY6jroEieguqjyHKWu7uoQCjF7/eG
uY/Seby1I+4uqKGsSSdjC3nMk1BmBBVlG0dknSOtYEntlS7h+Tq7ZjeeUZERGFzqYH4AGL2MuoOu
fcViQxTxW8BkShr7Lj+2afjyQhzD9GwjYUijECnAsc3F7c+R4m39tFIdv2MQrbfDgNbMUOX0F9p5
SApe4IA2JXxydLF+c6B34upPI4ICo9peuOmzZfYDRLfDnd9RiQ+3vd47aODQvaPjt9CS3Dd1vrPd
mxlgkGvD4saINmPY++rTmhVxn9Mf37sX+doyTDJWvhHOzyCyWbFGK/kYw6/eSbhgdFvUR8DMITJ6
KP0tzrxruLlduIGlwMhfWKvtDmoN687OditZ3nt0rZEomwfZwxtomprFWJG2GsqKxaceKhfIT1Zy
5ssPHilVbmz35n68X2GWU4/igicg1IY79wy1WxEsmtMtWufP14tdEKITZfAcxU0MkpPhz6GrXRIj
yHCy/LnkK7cclMayBRxurN+H9x+6rKNN/3u3B2te94AU2c1zOUodP9x97Xd6d2XvTj8fy8XafKcU
gFQ5aq9lrgD+AbU2xPcen37DBPfi0HirQcBcU6JlmbW5/rY2TA1PCJfEyJlxUv1oADbvjqfLpqTz
vJKItU5lQ2sxV3tP3CVIOnm62krgGP1ViLFM8BNkLKky2Fc2lt+k9i5FDGPkP7Q2ryETsVcb7scA
zyuBQf3pYaVMS64pwDcS8y56BoR8AI39KHjpGLpV64tsKl49jHXpcGcs2FahKofcXgKmEMgychkO
r4R3yCRY6eDX6FhVmP1dtVxGpEcwhG2ZGt7iJMHi8KhNi9A69Vbork3qJb9he+MDsBN2cjgr+MyQ
U4TeReo5Kpf1yJ6rkXAbqbjxuDvvnpd7WgFfRZa1UVRGlFRT+5GkosYZOVZcpaEkRGRbOP1NQ5tV
gM4+4Hiv2Nz3DbYpERmLqwEy2TX/7VIB2NyDboter95PgevQLdtRkyQV4KVIPzpth2VZtzV3JRv9
NQYILCD021G0W91Wv/zSOn4Slr7cZnWjxk5L0dP1d+eIhzN4SZw5/Av6bhRpN3nv4N0sJUIvASi0
OEbAlkFoXp7faarYjl9Jb0/Ob5jlA7cDZgUknZFY99Dts1n2TvNDae8Nz+4UfOfNttw4xgepboaa
+kzh4PTZG40B2z83109P73IMTOy3qtEpDG42FhqdShxbC7oMvkbqvpXCOLLyKE3mBo3V39X959jM
IcwV5UnhCxy5a6Dsj+Cg+syBRZ5HbbxJpg5LJ3/W9B5PL6UjRsqqQyKEBA07GKJYRLRnM2TwXVzT
X0JjQyGnfSYgaCt5Fh2uXaVsjGK62u5294RgNpI5tHKvBH5r8c675tuNyq7UWGW8sxyHLt8EKzqR
Gl7NMAeMzh3Z6kTH1PUjko6EDpvgWu675cNbiMAvJ4VaU0Nz15E0rSxEp0/vPHWWS7RhtZBwcLvd
d4hnKfHFGtfLIPTMTNaEtYl/cLHNWulAsHAmCHxnY58kv6fUnEdbqbShWBP6ACziMOLwKIfNHMwz
LmV3HRhSeY3Y7N17UoLaalqRg6JFjTKti76VZqXCa36E1A4pGtGimMWEWeWpFBJl5jNZYrJdMMIz
yzPDthe+uWmVjQQlMw/MiaQ1BDJmtlf8hlOHIP6/e5wGBcTUngeR63xf5nw8cyQGMQBRlDEPyhw6
v64qcYJW0welt+U8uq80/761mvqORtM6iMsvSuBOHFDMCtMxjdIAIb3nFKCQIJQr7rm9DeNY3IKx
xJ/N2m/Rk26+vn6MPKttV9SFuru+kTrg3xga461xBHvy5XeDgmye0y3+2PheRUzu3pnHIhBiGYoD
5+D2NijiFz5xG7LKriPqcVX8nMEr6xVI1AwwJcpIQlKFlyQRr93Azgz6tjcDoirLHuJn0+aSAuTV
uDkzEVvCe2+JTSQUyJckbFmyQeeFWTHDVeV5z13pf1lpGeQ2bxlEfbp8kPWVVeJ40g7nHdan3wQx
gUijXm5CKJ+0tZH6xBuUwp5DC9w4nTFv31b15+Fl7GXaKMW4XIJx4sGs3/BcJYhkWXq3GBNvDQkm
qPbXFNdq3yCek4mlR3htEtktyfQ2ydaREbINe8IDYZV67W/fF8j1lqIwXRWiE5C82K+WHc03EWR8
hlYLB0/rzX2hm3FEqvnGN2zhwuoJhV8c8pR71m5DhrECcGkLdMMEYwF5z9qG20iO2gc4r9UG3bEx
PFWMf9LAQ/roGVn7JyigZvX/LFT11MHe5xfpdgavY6UDh0B0Djzo5Qk2L28yTDYqtQWB/23BZBOA
0YYfQQln/DNJbsL+7bup/0MU4bD9wfrlnVC5VVfQxZNfJLVSESqbv024x6Wkh7/uhpnpdWwE/a2z
6++xwRiZKbdvQid98CXxdJd7pmidPyakSV8eDhuyBEH+/4/mAqYi8u1AXoo0zJaAKORMwLyKUVmG
U8Uuhh0sOiCRdKgjp+RqwwN4gj8qod3k88nwPzAXFUGfU+rM3whL5XFniMdxieqpyrnVuydysrHk
LUFJ9e1z78WO74Eh358puU3MQVuo/oPRS0OVs0APjKasdF1YzZ1xppvjFniEIHfv1lhKBnT6fQIa
u2gt2xE+sU9ESWtVjgv4dqCe1WnFrZkF4w/FpTcgtvQMeDHr7uvE7RwlDZoJw9PYWge0sAaMrH+o
WeqGf+Ki7I2NZcl5Cvngj4So2LYsD7sNcGAtCdbVETT+ICax8ftNyg0VIQ71U42jqrmp2fJD8bKh
G1M48ORZegsL6+j4jvwCK6V+LJ3Vh6ZTohpCoeaMgXIg2wBpJn+rRS0OHV3D68kAo5phU2wP5JNq
0Bcnj2THmGyjCJa8EKg//QJ2t5+TzY53XIPlfDdWQ+LSz9vSeW3VXjpI0AMMsFMafQcjjttbjw6C
RDIxcU/FsldCqByycpskbGGmusMQwWa0HBsUz91kNq3cQCiyVZy6DRfTx8bVlMHlKa+0K+qFm+PP
k7ubV+ToYTpWdhkYACwDhAerPsiEVRo5KkVPqs00rfDS8sUfcp2XUc8/smgHUGp+Eek89gbBxxB7
JjQvLmAUoMvAKBl/sQD98NPfJrKasUuSyH2YnkvGVtvuKv7XC9+THrUUDyUra/QsXdhKAli5h4lu
9QwndSaiXHXHn56GqGBRri2SOnEYpoZReDEJrxAFNX/i2mBJMJjzSfxNJf6eMNA2yvoeDXza8yd4
q9LdrD32GcaApOvo+o/IYg+BUxHekPScwiTmrrFj7XCFSHpKBPmcbCWVobc2tSaf5VxoM9k23KNe
SjYWa1GroGcW5Wkf2tAJn+JaK4d/LE1sm9/JjZjGqErsarosCHxHN9zFBZhVPoXFjiRK8F65U7HO
Dn9uIDNvIT1Tr9d+S92qHzvGCSef1xX0Lkel1wjNIRSZ9gJDL3pt0hB4Xg3lrFmFAfehcUqUUjyA
DlyHIPxKvqzPJbUtDRA5dvKtdxmmmuWFP81Mkf8/4Kal6MgX9h6aDI2FNd3KRjB5q9uUEI50SAUO
34ZxtI9l6YOqq90zMjicy+6yKk5lVeWmQvZERFpchXbjT9znzhHTbVRx/kz4U0+Asji9nD0NVzYM
yJSKeD8E6dlV6ibRK6rs6qSRhcyXcLt3N2FDUPtyauWaD4jP5vay/ATskcOzcEM51kBsRGcselAr
NqqYddGZgG+9nHc6E5vf3Rd0rSX0GueYGyIjpd2O9SCKZEdOmTgg/kIIT/m2AsqJ3nMg7x7Y24kS
vlZ/6FPCW6yauHQoDqxhnt10nLpCxj6x+3aazTbQ1IpTD4mcAqAip/EdkeSuF7dEqa/1rgyZflO3
n2Ldw/mRAPOMLj5gMoT6Ib0ZPrPMQtXMGPBArYQE5hkJkaIvldHRNZGjQ8U+aZYhHKELpS73r7Jn
IcNW9FgmvShvEkuYo6Lp+k6wNnts0H9Th8Ga7E0WdCzUo6Z06MzbpGt8hjhuqYjmlbuawGmoVQ+o
VQwY67IuplgRZoX06RnFEUP18KJ8OExkxUcmbV+N9lzJ1gM1FUoGB0L9AF6CLBfcPKz+EAa9lIdZ
+I7N7vbF1xR8j+LYAYAZf29dg9dG7918EmpL7vUSgh4x6+733trECtsyqzW4TcYrb5Tp0pQ65AH0
/49fe7taEWgTvxnoEKqHttjzKY1ak/zihlQYcqiqc713/QtfLns7fuHS5PO90sy3bAAjiBd5m+J6
lLkHnsRPtdLI9HkwHHgYVw0ZwnjROlr3jN7FI6tPakA7x4u2wRxXg/I25b12gOxMHXh6c1ODQmqJ
/hDH+pRSjTPAXKSGTvXe5ulHbJGXdCffwPEWmRmBLT0c7h29AOIYXxqe/ySmgwo6G/2Tv+cpVF7Y
quklmtn8K0cFARPuBfd0mWVcjy7EGhO5hVam5sn2f74Rs6+9NbFQ+I6ZfYtt8FVh1oP5nzAkNqDO
/KVMCer7/FFSK/jODpFoFAZ4sL7FDYrstTiFaXcffhXxp7cep989BPmcWz8zmy8XAFm0e3QWgXHW
gMt0J4fAd6459Dqd9dEMTIyKteM7TrdQPjqCXD3yh/b6mzJ7Vo494S0NkPuOpkxCvuku6OORs/B1
/+uhNtdVFkMxSOWAIt77iYdF0bAOaed4+tLcNKqO2WPwLTnXDTtS1OZMONB3ROaG4B103Vns3thQ
LzWxuKzAH/7UabhhJ50h1vuJqdj9Ok6lAopbqWPMsh7tFyUpC+aj88WsjCSgQOpEOQnRVtrkRI/8
vflo7cEp5E5tok8JCWFjGe/r8nYoDxKN3HRl6RGA8UP34aVz4WzVYObs7UgRR9YWpvKkYvr9bXQw
ypPPJWqCc2nV/RoroWkLXRLSjBPGCXQ0PZt2EWPf7zWGyMOYJJtvjrDu++GGws2eYjR77OQ687US
k2us9hyUHop4JRO4Luo9Kk0zqztaINKBmoNIumMHTT9x2BASkJRa5WjCnh2oD/NBTVJ5Hs52K3Mu
u/0pzeZyke0zuH0Do+YQHCx8wQxlROOg/1gyRaSgk+q1C0NLd92XVRchOF2ZB7C2seog7d5Kgznw
v2QT28E53uNCD4bfp9sMXKHESUsqIwTHbEXTMVy4a8h18JziKlFFwsmB76/ZnpCDfoxFb9qeDFIZ
+Ht/k8cCs+eG1VbJb/YcdLK6IyhOwl8dX6TwBgMagrEko8SAcESc7BYy0qa9tPCDzkhzd83xQ08b
NvUCUfr9BC3Do+Dtza1DYX36q1us0btSS97mV8WZjFv1DSevduOGbklU/jnAPXw64w8GDgmiNGB3
iFGSMFDkfp7lfAo5vXIMgUPqnYQORaRHfxK9MpgT+cVNeDswrLsGKVk0ABGCAzRUD5B7UEfDUIUH
44FgahVI+Pw7X9Uh/heeUqmuu2CMoW9KxWDera8yoBUEyahqaHUZfqX0NYF6JR4LZQUuSZcbI7bu
WAIgPVft/r8yd5qTxwPCyIDx5yMna2xC90feMl0UVTckPlaW+bb1NUNWEICbgm0Zo7710JvRf+b0
wOe7aHgqpd2R61fY8xV5tnW44fGqiPQ+tN16+J8oiyBDskEWwI4UgE9f5k4woXRRmK/0CbJHN9Jt
9wSztAimJ940qhBV5ZkUCeR8rS/WLDAyA6ucQXhIa2Gy4Jpjv3YyofUUl0S+b/eFG6hupEgEDQOX
sTRcTOY0jwQuwqDDLzQUcZq6I0ZjZBFqPyEdWUarlCqS2BHfLPTQQhnQeKMSHBYwCLOH2Fbi+v6h
I+fEcklWPNZA23RsB4y0H67rMWNETbU51Q5BpuzazBNNPf9xoZab+E0oVVRGRNrVtXsRQh6MRolR
UbLejWkCh31gikS+DMd6TDzHWS4I2Hp4LuMmh48o15OPKP/6WK7r8Sg4sTOg1ISssmW3769uavdP
1uYXpjyrf94YQDrpvkRYFas1AFlVYYndWGLNmBjZYYLB7eeVTu3mJmogFiInjbmRyRcIHZGRh41O
FX6TgF1T/qKPFTh4+9fyvEEoeVTTW72owybhEyTx5oCncdtSm3uwkVmY/V2sr13RsZDzzDFewafo
yL4Vlw23/d84YatPbDCJoKnmeExabloJtGDqucpgRlMvsnUYUS+YPJSKmOx3EL4h9l6UI4OFMYHS
fgeM/WBQv3AGLbbrkADlcmSu0SJ2OmtrWB0KyXYxCPX+b/f+nOGc8pIFRW4XQtuAxMx7ZsnsDNXM
6uJhOSjX+8wMQ6b7Rla4xZI60RG7sJZx5hOIdTHg8eR6DVTmrEcyKG/MmzzaO+NZx3tvn7zSNTwX
H/tNWseA4ougcaBQQfW/iZwahMAiP5fjrjivETc2Gc7UuPLUrJEmAcd9STpOZ4UYS+dtbX//JRwc
JSbYkqiIDe2VTjmoWwxbtZfS7ujNYsHT/ru6juiZzANSIompjoacPG3GMLxlkPR78N5kJEhaiD+R
EmtPI0PUsc51cRxzGIq9qcED6IDIUF9TlHUHGzkPp4o4K7TUiEHUzqt0EZFkl7CNmjYlnMUpWHQ+
WSlvs8OzPO7At7/0o2pFbIBkKpBR77ohXJ7IUdPl/YM3mgeBRW69EsTU9WiVqqYkeTYgK9Jifkks
s0lRj/VGa+f2zV2+8R4brPdnZ50bHBZ9nOpAB3+ED2bDUb4Td3lMoc8xgruf49A7LHKFKojTHGeJ
1NAfZtYekvLu5j5CUPSohjC80GsOBaeHecN8G0HJwzw/wNyKnVoXSRbtbnP9Xx6j8DfJedhUYVIQ
e7NcC126yQCHQr3zWF537QSyOyjXSC4anGWMLBQ81lweHmGZxFKbPLYAQ8vI4nutKK5CeCMQLRj+
ggCQcoZ3RPEOvM0mFU3/T4X+P/YO+BezIF8ytqaFGuxjMN3t106gsePfwfl8NtdzF68K6RJ3ccrQ
2cnzzwiuytEHpU7G76IwVipKSriujpPybOlcqaLN97/6Ba0p6CEZOZdVNE7/v7kLXwkWpAsk3UqO
UIEIpgjbxblB2bu3sH8bbabESXgqLsgLjnin4o7Ah8waEkpFDxK720OL0gjJwnqj8/L5h2NebEdn
+yi8HhTW2yVqa3HFsbfesfrTVtjNgn/hOqlAyINYa5cAMkPOqHDTkPZRDCUn6h8SFlGUaVlmljiQ
um5DAUKF7hbFGyNd9BPfQbsVFA6RcNn0DSZmiLIEb+XUMX6u05DEqqztaR8/bldQ8Gje6nVIQCKp
UVmj87bL3Qa2RKQu4Q+P3qa3XExpp1AGnrBh8rMCO92EIhJ7KiQwne+7qOwVWmZYBmXhPmAYzp0Z
PUx95jAAy+eA50CH1mzzQhMy7wQv5KKFJkV2ehFor/HTSydWGCDdVYazgzuKTOQjFaEhI8y5cO5J
vY3fIrSnz6KSDWpEqBdeHyjKvDkvhV5kWBvRUpmQBtH+SNURwd9YL002Qflsautg4o1/e+yyxfVo
ey9z6g7lAyT52K9oB92n7VpP0t4h6YAVUAlD0ytuBmNfX2v1YPvDWtflR5WOSyV05ynUJDo7PTO/
QTdaVrXyIMy0CzLTqmgdLij1d6u3rIwi53z/P8R7L1NlyakorjmMqPcsJ9U6HuTuTVKY9811K7y+
rwmrNx+p698/7ys8Q9T4499ASM17FMcdeGtvv6FOkWZllRPnVHnb8npVvM2Wsb3g7ap+o2zWg4Fg
1n3OW0dt/Wsa9Iwstq3fmJGYXidh0L/2BneJtQ/q6DtMORb1MLm9feX1t/ttP8h+qELhyncoBq+n
juv8j6l8hR0QImXhJiYrvSI/PpMC1m8o3YDKGMhDKNOWje8gROYHifbbGZCz/and4F/2dzHsZmvW
drMV0jXeWVy6PziuKgcrOy9M2NjVAHW96rB8rCsyQ4jKdxazqWW4Oewi4pJquN3Y0GgxSbDJhUBt
bem6UmpySgOUVg4idNagoK+szE0cWjv4QhI3ariczgTabUfmWcZxyXLINrgJj6zYcwUJas29rsxy
HKQMKSz0G4732cETyUFeit9UUSgUj2jretm/ZyHacpRZck4JDnimQkfc9m7qmPWz/d5doGQ4VxoS
PdK2mQSjpw6tDFyxtRv76FRijeIgzhpaQ9LXWYFq5746lNg7HEwVhx6yM4Aw7ytbNAeeK4Tzww7E
GmsJea+Xsl7fDG5YqL+/mAvSbJhiDdOgLaogTfdEIdCvtoLG3ATHyjeZLWgvkO5Uy3m98mFPsEeZ
FQBAOIw9/sxdB1BEFsCLD8WPxQpGzPPZ6pi6nv3bL9UK05kMULAceAfyYGmdcnC3D0TFlstF+fvW
9gixqPsscXDAovoJgNZ0w73qk1BxGGhhhzlA+3mi1sBVp9YTwuJ3WcYTnYGkpF1qz6xN4Iz3IolH
IiuP9ZsJpDE+MMBvyIumxmYsz5vzAgBPK7qELWz2SYMViZYooESb6cHmQ+SvottbZvyr5V0X5FkI
3w1fP4UVaUy3V/unrR4venk2c7vT+yPWhUOc61x+JmRdfhPrugweE39htkCJvv1uBQrQ2QKlshdp
72sOtqeFfyE9qWUkeyyW0EU4Sm6W7ZToRFkZNswz5wm0DETKIdBTSzyN9xSPjEvXC/bxhdUVQEd4
+e8PlYqzgZ0+1gyELV6ejK0L2D1wX9WFHCob/yPqFwP+xlXtRS63b11k2tTzvlhJBHfB8D1HYGjd
960aQJt9iCITKdYyLM2C5Nz9cQfo7IWCU+xtii/t+odrwJOjrJEsSGzOpYHe7v1axazpBqSOViG7
3K+l+SKlefVCH8Ti+lHmZVMefxw8SNbXey/NrZ+nCvwmynEfscFirdlPSzCVfEl2Tf3RbuYC5yBA
eLsaja099aErNHQ1P3BolkRYV7XnZBISyVt3iTYakAAyVS4pYGBFBN9vaEuWcE598p/3nRaAFesp
m9iWaEDlD7oP/AD+n//bT74SEhtoziOjPaG8Z3s/fm3OhUXbMhWcXL7gsrX6hkdMJVhgf6SLH6O8
EWRqox6dF2o6Eb/ZMEdVY6gDkf7aSyy9oXCUFsSmKSPKAlCnjwjjRz+AnaziUR6GYif5z3tVzxio
lKkBEK74H4eQ/pGtCPBJsI7VouBTlyMxDiprSqSoyqkBg5w+jmNbNSbagweCkhEpevnkGMehhqn6
uyaSgsr3kBr7s5LU6GTMZxoie3SCW10v3eAkGzK9Gf2VJDvL6JBpeEdvnRiU32uzNyrEXVH1vlfF
MXNl5+/bjqmSMMr/kJLoMSyKEFT54d+qRSJIrOGUB96ZvJLrkkERhFKt5AO7N3vN9E2HtolFArkJ
X16JdtGAYYRLt54nE6N+gZh0RFNeSmwnFl1oI5xcGIoUIbBSOBRNcW76J2x10JMNeJWClp9ZzMux
okxo63KFf2P3lcdr96LYvIoHlnYJUx9qPWcD3bCE5G5jtuRNH62tyEkZt9aLScx4u19WLWPsAQ4z
Kk499152KV7cFFnXgX2NkofZEuBFt3FywvVBY6HiiulWa7xCvQAP/y4TP8WQPMhimeH4hGxr+9FM
HUy7cz/7wSiAWYLmNfsvCee8xoSxRbK0VoKq4YTp7zImlrlbDT7g6bSvNtDQAIB9RalK+Z+6iQNB
AXVoST66OdL+illzi3hr8RdS75o/apkPWMkSEpDXuU4rgJKYqF1tkndVFDDPuKjzDxbShdhXdI5t
SscNLbfvFIrCdtyj7M0GOGshUrwIz26nLvEtBPx0fvFKmZIO6jt//zvhtllkD0UjgUsWcEsvGeuj
Bjjt/Yw+Rxi6CP5E7U1BEfJl72OUXk3XHUhL4VoKsbuwEJ3XHhj9fFL0cGzLYoWWl2fKGk+DAtc1
y62B+Le3qP/kdfsD1s96mZKPNn+pwz73ga6OoTyRHN0150mCnG1pzrV4D5rthx2UlOY/BRTa1XIM
+iefYT8zddSYrozYGx9GaAK6oPcIzJM2JiVUG+unn2AU8JmgQUXeaed8skKRv8tAUcZTNgrZ3FxW
j4SNUVvgZ/iTmCLBiKW2Ya0CuQ/z4hdrekXet87ZVIcAIazZIYyZUnShBmpLiUY06Uy7YB1rPVsQ
ALS9ZsApmg/GFN5W6mS4jkXoZuWNlIRMpU2U0kkRpLf7PO2GHRaMbKwG3+ziVWOmvhorfha2Qe4B
p+L3jg+LLlqVPJo2pYZgRpIWzhhF6m9MCldCb1yzxBkUFMn35JAyOT8EmQq546u1BTSuS0y8O69e
SpTq9/r7t3s7qouEwq3CSAI3tnkoTXscMOwwebAJPR3AELwe9r+CqioIGFpmdrlUL3Q4uulweJEN
a7842GvGqtBq9gjVQDeGUYWFU2HOFjn+wLucePxxKYOcL8L2FoH4u7ohI6Guwb/AwRZuPCFQ9CkF
pQ2pXWYMESuQrqL7TXdNYuj09W0F6n5ZkCV1PcLDzaLlGX1u5R82CTq9tk/5B55uoZRERX9ExkvD
Iz/l6PItGFBAPzRZAnbpHSVQbOLkPyY3TKmTN82HqyyPJANrq6wNJs9ZRxNdHwnrJA9xl0vp5n0K
GecijQ9B/Q5ZSIRxzwL2gN2R0IDryOZ8wp574evl7QumnZ2Eq3xSvVXzGrJ6cDisrIc9nD5tHMit
/8ljw60T7PLqarDrR9jig5GM6yvva0UWeLGs6/Q3io/jZyfaHZY5Gia+hty0Kww8Z9w9we4d02wh
KCBKmGJQ4lyhNXQnspew+fPMhyVC/M8Z1pzKWQx00U9VylaX2z+xgVfrBqgPCAk/iWomeSVbRJB0
pRn/UmjzRw07twOfaEHVEf9z+kSWEchFxbHIY9jujUM8wddYwkkpZD4N1dgE/yUkfY5pW/J8Abmr
wMhNtLG1+MYF7Zwn1UKiSdKJddu4QRq+haVhvgUhSMelYeK7+7k9N6d4071pa3bSXeU5vxi6DOFv
KMCQ8Y09kp4/qHZ8tuol8PIYuK/ABqn2D+kmhNiMmiFuDjGysyL+sl31n+CyomSnCwI6SXDtHanv
6Uo1r3RvtCYerBdA0aGRv9jyR9CuHjclQFAc8J0nodjGQ45p22SoH4/oCIo0/Aq6o3C0l8dIli3/
Pok5h99lu90VcQmCgvIsWeJbZV33Xa1Tpj6tm6quewQpUgRfck1gQAvZUcKPQsN9u56AgwIX+HQA
Xd0riSrwRSNKh+19suUUopV2tMuF7NTh2NyAUdnk5nchk6upqPOrt5cAR+ym4bbfLRCy2SZ8KEZC
oU8TVpaFOnpdWGFG0Ejide8l20bg/yNe3w+/qXbGzDE3CEpUiiiO7DSw5WZT9vldgubgs/9w4inJ
gNOiXA2Oe7HXw0boLygVTbBjwsye1XqvWgOx0h1QaMsh8CcvsdRweJ++rGZgkj98P4qF/OyaE3ti
Tk+SL4nRimOojdXEUBvW+Rk/3O+s9WRx6DIEShy3Gs/PRQ4kLbwDU+rtWbN59+WnNZX4ZThvpi3k
UcBNvEXnLny8R6ScxPj2A7F+hQCjzQFj79f/STgFU8krR2DYO7L3bBcV+fw3A4+3Q7ULMIykd8R6
T2/Y4rknHwOeGk8310wEVpVCHRZsSoghPQpoljlJHpHgMlHQDdGX+oP36EsDua2gniHADejkOnU+
mrevQB0pNf+4sSjGilo75hwhLTS1+6XQZkKkCD3RMc1UId7Yn8FUGzrzDPoTSjHKf9HL/fk3ggrx
c1Gdn0jSSKBljeTZ0iCzfMut2LgP2010nSMZhturLStq4HHuTQWBgs4Ac2V7fyuYKz+2KcOgysRU
NlY7ZA+UWSj8DEYxOrITaNdHywAyPwwi5pYxhZl27bfVJKry/MC72BgRLF3ufzE4aJz1xmMlRFFp
90NuqZULkGNeSO+92tolRRncRpMkZRDBoInMWedix/58b+zWD54IVb9q5VjgLDBK/Ks24ns72cjc
TqXvJEYPGxo+0BS6rDxRVriTTxMLz+LM82T5wH3Do7u9BFcbFKDgg2FI/4ESxGRd0MeWoqPT+3Li
ASAgeCvEv9cLru8xu5KabUVkCT6exHTy5I/Tp1q+/IPJxUrImupKbRhzeQk9QhSV4YfVqg3EuP+c
mw7JVK8jDXOpyHPlgdrC0nPPpOUHYrBE0nuz5bdQufV41r6oUvUCg0N+Z7QM/xd05lit3dRyyIjM
cHrXDZye5pv6dm6z4ZT12joMMUGc2gXS79bTmW4sIEmQP4kJEQOrfrUeVGvjnsDE+85bTvjRkfE2
s2RpejCGA5+6pOncrUg3vzMIRHZID2wLnCrjz1f2aVH88Kn5PEjzV7+TtWXC760a5iI78oDe4kKD
a198OmElF2/qfcv1m6316X3l1uMce5ahLsKBzMBBrKO/LdLwrpR24nhMpzsSWiD+z5PLEkbISHJB
GVYeGlimc+FDoqmQxE2wDnQLFmUWVzEWgRrbYEvEjhYM9Q/o6AYeUkT0eAyl73vUHyo2ZRHO0lhR
5EwnYqez9153iC1Z2TBtkDCvAulrcfWgsvYraZqPzbbOXkNaYOY74/cX/p8bi2q0GALvnHrX7uo6
xQvrN/ORZMvcPtbrMhBO0bDEiyrjR5ICiB9dIF4KsMptDlxKahXjjpmXPFIqOKqhCc7LzacNsbzz
Mr8j++Dg2c/XPVads7PwhaXf2yrmV1gJTz9SfDIU5q9s4MBL2yPGCk80buEhcUI4bZVfmTUAr3CM
LiQDy8dq/dr7wMOShYdcnOtu5fPg1TvkKDkQCikUEaukQ9/STPi+eSzUJJLy4eysowgz1/xY4EsU
x6rg7rYycwmuPobrRfGoOiTXYKWQlctvfa8eFs22YvHAoG14ldwStbi0zPKwwZHdTBEroNmksc5h
e+J2v7aPDjc7pXhYxp5IhtjWgxaeIbRV9dgz6A0u68iBttH9FguEd03OHFnBv4dnxcuRFC6XwF1d
Frup4BWVFI7cyXiqUFtrrHUaOUhxNC1VRErSQYdURw/Tv15vhd7m+HspaGmRxHMbmjHQjwdnd94n
PwwlDnYv9giv4LlEPuj6GlLjj7pvBaoNQ/QocA8+P5xznPLayTIiCmoZscRhl32++EwP8FN0mZu6
zI78yfaGufmmnNnTfKTRzcPGomvoYN0zNcrvOyovf8gb5AXDQtJovKOiXRFsw5hCC3ZbEnIqufdr
qoUvHV8VFXtMyvgkNDfpd/rtSoQJC720Wvn+qlc1mGbw/01iGwykhd+FeI+Sipbmf5YeO8Z3IKjf
H+XqKybakSqRr/rV9fpgqieoouZtt+QII85xtjI5/uUBZPS5MN3hSq/12KTX2WlFM+U7bwjYVeeD
FW7dwYesJ7CFfsXAMtsV1k4Ij7p8uNmdUmwTAd55VXTWO8TFgChncJLsaKNt1qS8M2iV2idIdjMB
fsoGQ9ZSVIf/Vwxlfq4jsi4sZL/xemDIMrLoEGiGKgycswlM64LwKXWMHJiVmjJ4eoY28gtLtrpB
WsMhWiqg5UbntObeLepurCkyLqfOChRfR5eMUFWrlZq4VIx2Fjmhtu93VYvf/xY2ZAXwpxOtGuTJ
U9RJj5l9anCtvRNue+NxRhcxzhAuVl7C5b4imS6uDZ9mnJQH1zyJ/gu76+GVYK0YpievZ/8W1nBH
8L70ku7EQJYjorIi1nq3NTr5+3fe35oyY+HVTnDD8IhCkTHfop1VGIr839wcLMuDzdacu8sP5kXM
ETrlikRU57qltkJsUpID0QgmASf5qaGecVjSwswo917DdY1NubOVfLwfIOzI8gal5NOSSsDN3iDL
c2RNe9a23HMgHXOedm+RnvIB3f36Cl78HTqAxKxypzn9ACWCG0ADoEc9lEdPw4Z85oMv7HuvdJJi
vg4Xyu4kGVPCjICFmMmi5LTPhH9fgjx8fnsdWnY33aEGBpQP5oCYRLnkvjOIOmMOhu2LyawAedEK
gF/uNgATUkM9fRkv/ijTL6iYo6A5iSUA6Dzb+AHr2yEo9/ubTilHqvoVTRvMP1d8S7WUWQIrLWj2
r7eJYuahLVhiJoBrfNyYovagZJouPMxl4NPlvgOS3P5IdamJYVbfC+hppu/VEJe6z2M9qNg9PfTs
yCHKYttRqdurmf3+1JFQeQEtktCJEmHUpqSKTWvDG0bcyGjbPOaPU7joGhlzDHIHx0L2BJaYYRdU
AYLR45xVMy9IF7D7xToZszsidv5AiEpfgWIzBxi1+JJBwopMDQ6b43wNX/d6jeq6n9N1vaNyL++5
k4jrZHWOJ1MFQRIp5YnzkXaHYjC6sxuXQiU+VrvGLYulXzO4TnqsEQQ0noJrBoRhiWrdkS5xl5O5
MGPaxA1COryUYaxL6fSnNaA6fkFkHfUf3on3zDPYk9eRkfuqg+QOg6yVpNOhUizua9KPoGZSaeLw
k2MceICQidjhvhH+avap032Cx31MVZANQXxJXimcTbb4XHSeVOSmTKQzcT5QLoyUnD7iIxvg507R
AgtajPkrITM6jsE6KY+sEpitw88lEpaoDv9e5mPyyu4Ny+kVBdoQjapjOVeJaf/bjx8aEB8G1jvP
L7mCJzvTh0kNNPrmPoo380bg8R6CCYFBISTXN59xThkLAihLWhqZf3Kqga+zs2O4gjwk/y9Ru8Lr
KMKPxp4jf6xmy+oujM3/38eKR3kK+BZfh/0nn7KMXSbL6qIJmst0vv5vKtvMiCX8v2AgEXmf9SDS
ZsUUjn3fg2lZ8YX3hcTrI8njBHX61opHd8ZtNQMy/oII7FdstXzrVtIeyjgS2DPpbFEtG5+EXCAB
sME0rbimQvn6wtaMjlTcx9r88Pbgx1AlpjYIiX5SY2X21th82CKkpr7z/AZfXwOg2MQjKH5RyXXR
VWSnTCFNBelkp0JPruzpM7LfVcQ2eB7/l+IVBf56wDGaa8TyXG/PUIJP8SEQtKVjgD7ZzsLc8mos
/T0Q0K+SWaWQXDmGuPUKxzFdlb6BoZ3IPEwcZ7mJIalS/U5sGoXdIm+xjvKm4uTAdWZS4mYdeUWX
i1b1sgfOhVO/pBg4UQGsA+n8Uu4doJowbBEcH4H7nEl1wJvKPiYHivXC21SAHsbLUnWAFsGWNm7i
GNN0D8BSgyxbazSGy4fuDd36MyTsUJDM13uiapRW6zltsj+6FKckNkReYE+2JBMv24suwp49tNQE
N5LhdMOUbs7AZyE8uUwpdLBpkoHsZnklEd3Sw1wdttFkV0jfaxSU1MK0S9y7RhoaRqK2qY+ah/6G
V6o6BaNB5EwqHf04sVV/7jmz1Vv2IFhL56lIqyybXUmn8PffFOjtn4gL3Fkjp9QJzKNpt3+74rwz
0zCRQyEIipzWQ3u5sOsNLXO94m7dt7Z902rrQEfR0hOLbaPbQWtXgRuBOZurB7nIqJDp3El5EeFA
UWpcRFgYUBghPOLGgCuWJZSMA4mkOeB7YefiXbdZ84HRqKWjN3jhrEl57AOAbeYp033rsUZYx5K9
LBSTZdECu/LH1MGQqKlVtegcP8XzUGdXwsXpWcV/M7MQisFO9e3GlVqlNUW32vVw5fruJ8PC1oHF
0ZatCnVagupjWjeM2QxGtzgbxhHQwd6yJ/B9UNqZvOXDtIVC8FAFYiFFUXnd5s5YRf2XSvOUu3Fv
juGbbup30eMoZy90cCiboBUQWjZBhFd/tq3pQQD/slbJos8Czw5ngBTO+di7QRCdvWAj6fCPWSfk
KbeuSajOGYkFoEjZfLoQLfBGrxDcmulLh0vCNGgkxLwZ4+glwhccdhyl/++6RGPlJDjehlcZYxCN
esdthylFNvwrQrhkjlShlOEqYzOfwXQW4JD1yslOCghbpHc+0AP8+OFU+0PRoEw2n7ZaSGwTdLty
Jdmfm5peZCBeREhoLJAHc8HDj1l0TppUZcKISWbNO/STPpAR+sZUJfqi+EK98Bf4G7lrr153sR86
y6HYEjtaqp0jSWLY29cVQbtiibUgb9MRb3qWMmy4AbPYmnBSAcHnLXzIVG5J/T4fQuQ0+VLbSTc8
3obL/jIEnRFVpEegmk8Hw/U0gWVOEU5kbq4tbbD7rDQi57vS8Hvvy1tpWUeFOgRt3SAB36wgf0Cr
PL487rFdabLz+XiYUy2lycfFLlm7GE441eH+kLvKsVggBke6KchdEbPscxB7qQ+uI2RnWtZkXlkc
iRDLLYnOLBccdEZn4wp+FtPQpEoEnsqEgU1V55XlGzc8BRmET8KGffNPpP0gD1bs23wDbg8pYOhJ
ixnkbfY1Qa18pPNoE+9KkpyNVOXM956n76oIclqJ+K8dIAKRKRZY3YaQBDsCn8BkRTX8WdhwOAaK
+zAopTrB6HXv7wjDMqBLerZyd6OscK3PoF3iu3p6xDL3KcUeoSZH28egPVbc7GVDUACAlCYQNSDq
+NomF3MQoXPrA2wjXLIN/lonLJpMdOzCLPjG9Fp/p9V1eru2IV2+jOfQRAdj26mM0KJJ56Dsr4zq
OAPWsVMKddLoIXzhWrwGfoNNDty+4L3t4iw/BELAdrn/pfBd8+kTt/how0Ihx+Bvgi7OQAPUUPZE
bg3JrAVTAqsLYZHy/LWU+FdMoq+upescaIjRXlAFwuSx0FQbDSEfswu2oEtsLaM/gzFbqVnytVLW
3OoMa1hdI7JWIrT2aNyNCXsndSx2oQRo1oksWagCSPwy+8PcNeDHzpoIdj19HfiVHEk44DbyPUjA
3HemNeMopNFDP7Qm3U3pjSz7Jq6LgUQ21Kopo2qnpo9kW/hpWr+QwHPTvJeoQ3hkYbVOgJHyVHZX
q+sQEtiWw4vODHVn/ZZq76pXFbdIzq8fkClrzmKRsurwzVLksdX2bQjb7gO8t+wL+TZGTsI2QAsQ
lM3ErDx7X3u1iGCrAnaoiZ8LTBQe1Do7NKYNSyNPbOzpdw4upRnQVUJB5mud84WC5hrZlWA4rP7P
JZUOthSMghCX7eJbjSvotgaD+VHqji1djf2chiK69GnmV5HNNc4h+wrGCF4Dnj2us/IWymBvyaTi
GILcwPbmPO5992/7xFqmrBDFE3bHZbuObgWSldDhOjfz17Ua7tyzexhZ4auwRbFnhD15lTHyUr2B
xGqi8+gqfeOLCwco1XgvzzM0Cjgptixd7b1FSx48G+CEUDig0VdOCOGYOvDiBt+DmJ+wEB7Ie4L4
EsgMwBlAThOa0rkurXWNB0lIqq9wms7v5ff4swvkADZ1+hxoloSDBCLtQG/xnzBkZLHrmwakDsSV
5AZ1LcA6Kp3vm+FoioEvTYh54mCYUmI2VLqqXqj9xy8DVvLf0rOQRd+OEk3Q953wr+YLNF16z77W
EyMIlvpDaBAvR+760ZqOkdsBoCu0F4F7mkX3SOl85Z/dKOIs2XUwVWT8HGXEfmNthIIcX9FlNC1H
OTEl7Wc0y+UgKnrrajdMgOvzSCWeM9sipXj15mAiN0ERX/3U4F158jHitGg+GJQvrE0NKl7TT/pb
86MihGpuajF2/zCsUnkEeSrSXcvVrAEXILoUl7FPHynjFZ7qh3ja2U/HYG6ImUaOPJep2WS9xfpe
IU6eoranPNvRJiWHwUlF5k/SJag5csiCJmuVvkPR5NJWLlMp1eU0vReBsc26CKoPlE0y3xmLAbsi
//Mmzw9nnX9xoa76Td0rz4sx7CDNrQfyToeoZV/fANwu25OXtVWo+KbelXYxXJlAe05/DumEfnsc
jWjTbRvbfPXffm385s0DbfTKOZVuXSC3EtztjzA8RTGpRE+0V5evejtWbvOEc0B7PwGB6FQaLyye
ZkJKpWdgzrTu99m7tvFN7nuqFan+FGfXA/It76moOZaeGE6IVR0Gv4s/YGoVS3REWQ/dQk1Ogie5
qgRrF2h4azwkY6nk7MWUZ0gB/weJqgeU6Z0a5RmbjFXR6QvxYJwFOxmju3/xjEM1wVoiUAMX1F/U
wnMiyqFtitG+OnmGaXeCg+YXFjM7gGPoR44oqsiL6kZKuR6lc/+LcMCoJ4gx922ibym7ww2RabuY
AJ+hT/oObAGHMrBBGQZV1l+KO7anbc/UosXF/VYhB83XUaOkXu5yRj9wUmkLsO9GZV31U6XbmSED
PdvDzYEqBz0y/fGCn4OPr1Un5URZYZkn5z838Glpytr14lywizp3qS7TwvQ1VTlTsQ9p4xW567PQ
JDEpbqX6E5UPOoTzo0fXc/iA3WfeuVGRAcXdpqEGt5v7Ciur4K7PdU7BI3gVkNP9ZFcM2nib+fp7
eUKREBwHkdW14AW1BhOvVNMLHUDl9QmswlcsbG/FXR9LlB6AtRTFcw1rwBpZeSjd58yUcmNsqYkK
m6jaBjgB54yBJ5AcWtgO+DZbfE/w9kxQPWSnm9mfeOYk0Bue2qeNP7CGOsK41QlbuXAK+Uj4oM+3
mDBdjaLsLoQJnnfXSUCgemh0nNgm/gyP+Kt5zsdC11hsAf21i7FytykK+D5PGZBSfrCU/KXr0lL5
SgppPw2tYOfP6E97EZNW17DzFO3ka3IUU/Wf8gwqy9LWUQ3Q5QDLN0bs0w8okdsdRYWrZQ/wu0pG
JcxeQoWMU6YIFM8ad5fbnTwjdKtdYTgv4+gdr8TmgZFnW9430esG66zadFZScTFwoAflq23V7xV3
DnqAukR2mCFmMuUZdMiopXU6gmdTY5Ro6scifmOSRnBp6XQxIEpfVkiLnHeltIuD+MMO/D8xnWQJ
DVH1GMXWvWNiqD1/nfp5fdxtyJfaKzUMURVgYxGilzMOujXCjKopgCrVIv+Pd4JmT0Ii4P2XNkA7
pmHpgfPMllFhF9/Qd+DzoXaqBZemBGyszaC0Pi1MxAYBCmvN2VlzI8JVasGKY1mtnH8HVZRq4rkw
2Ry7UTi7H3REXnZWq0tE7RfUYSDks4lU487sup00SzDO0As1DDBotdj5VJokUP0jFUz2gfllfVWH
N+aXaR34xS9MXneodH8n6kW7mUQKtot7exiqG5qiNPQ+f50g0Ccz2PlZCbMs+r0ML5F/hkZ1Wohx
GZjVJ0r3APzjFmNUHKlkjWZ4fneXLUcMBSwGwi8GgcPGTaXdr2j4N7X0brJmC/we2Rrnh61svZ7u
xfoh+bJFB8CAIPqEL+sW+mkX6y4F5iVhFMzsA/FevUej98SomxXOFJeYLaeLa/IGA3yaHEK6ujxW
/UP8hth8ldlMcUW/xeeDHhRZgfA0x5m9NBYOpQ7PDZ/pilnSfwlq4i6tiE8o0QrVd/DPgFA1LCKH
0iSBmKIO/wQIhrYiGTy/v25wwwGbiMGF1cWIanXaKY3sGKBF6sbzfGgSo7++y7AdbNSnXcVizYLB
TZO2IwTfHXjhD8HGvAkxurUki5jQrjwnOjix7KK31BKGLLCje3WZc3cpdBQBYH0owdefWWxkIcw1
+POmTNYIydb4bL1aRh7iwQiO3Ze5EeC4HKpL+KDGVXzuMyNTID2vZKtnFIvX+C4TW/CtQ+sRMNOx
SvDqB9r5OxGKlXNJi/As4cyi8pAgEBXX/rOkZO9peEMZqjqG6ATwqhyD2WFShg5B0/6puxDHPtTk
K7jK+9BwyGPD29a0L+0DtsLKru/lwBOvze19AbR1s4mImrMwOio7j5CN9xXXOY8WAdOWnuELIzAd
vqyJbX9+x0dJZHj1HBsP7On0vteKN/O/bxUFrnvU415Hc+jW2c6P2zQf/hrMNFpm1bSdMBboL9DW
QVyKgzHfnRi3oxsvVQ+nHkdMs5sYtEu5WO7V+rSbAY2yP5agLfHLFou4DVSpEDzq6XhVTkMDkb2o
2Tp/rIqYySzPegOiUNth427lvpkPZ0zSo1x1CdVP7yg3oSTYevWDD03lR9HwdCK8BQJT9RPFS1ap
Nnndut1AtEDW1ggbR1g8RqfHKU2aMqeHnJp/m0jr3G5c9BniAY2cuPtzCENXnBrEGvoRnRpXCMsI
FKFsQ8wFJ7lm7gk/gPwYdPJyBulxj4BWCJRtLZnooiJmEqQNtvBilWL1es1SIA2iuUg77dvt2WVc
j/0Xjj5Dy1PzRaG3TyEcqVHephtw4HkIOs35Ev9lKtFtoTLReVEAnzVzEzlCrDBFhXdelEDp+JGx
/wzfJSveG/Tpj3x2trE7AoIrHhUEtcH7so5C23f/lWjIWshi7lDnhQeh/xl385nbiIRLyiUMyrQz
fVLRImBeYJmu8Q8XrlXY/nuGLjvPq1vAaLlYT8uHEuyDgWndBFkosapZjr+sJUJ5x/Fj6ku+iPq9
/ekiZ5idCtidwd3gqzVrEhB9jbKsBMR1v61+xEUc9Bk5D4YEOKhqeHNPk0hJQO8aG60vcY2Nw6Pg
V9Ueu8fvvUlFpqDs6ZrY+OkGcD3OcXv2yeTzPUWGurBJEo2mTE7xHq2ZkwjKXOjtojt+0i5TdERC
clk5vA00w9EKOvnIE2V1YXmGlFp0mSwQb3r8hqFxxPuV7Jemnmo2dychj938wGebitjtoKRCRKeh
NdPDIvDg9t8k251R9Bb6QO1xZhYdECUvNlz21OT6uFd5epSRxMnrW6156Ghk799j1TCi0g7kpmnI
kvnu4ThdjiP6yitMC7r3F75nTUlUMokO1K4xmB1QJCJjCYhhsIjTildYRDqSfknbER7xrLYGYBZj
07Hlp2cpqofLIfObFWszpQjpZLMvyou4+IRskgkY7uTKzZJ2Bw4EHNoyTHL5mS6AOi6lmVXMcu09
i5jcXLob5gsEZT6eH77QkwvRwLyC33IqUPmuzQygCAD8421wmuCPYmbe9ztxnbR00hriqt13uj2l
YHJglDK8VrxzLe7pXxQY/vW8NMLfCLaGuzgPEji5Xcw23K6uRMsOtUMp7PXIIiupviiGlLXmVB/e
7Wo6NaaaJqVyCVJV2qjEx23HcdxnE0LZjXmSNAMOJkm0Pw2vnEComjhaO+hHRw5zPGnQf2wc3/7Y
AJwW0rR12AGq8d7K4eWz+RdQDZhGbE9mtaM7imLG5wb5kD96qoKG0P7KWjeaVF0OmlmxTQ2C/Q+y
WL0LWyaJ6X7rV47n7vwZqsYrODUnRp9Z/sSWYjXLfis1ywZ1ryh8uKaBj/EnCMDxL4UcbXKvjCeD
uaQR7DER1KPQCLZVdLZYaJkdiw1yWwygiNtn0+RaNAX8wO+siXVBvKltLnMCje9qU/TgktpgrDD+
12pTufnPJ4lKik+JhTu0GcSaXgUziUcgnq+kFUdaN9i91/kOTWVjQnjTjvUIS9crUmac4g7BlMiM
/S4sEo73lB1z8QnW6EDziSh0fXQmLuGTX4JbEwSzw2IyxcnAQi5pim8+BnAkyNOCoN8BXgynOgII
XRnHBQEDSrlXHhCa52nmg8YKm0zD92C1eR/QyCjp+vwP5zF10B+IpQWHxWHU1JBT32yDwez1sge1
2qaprtZBY2Sr6BhSsud4xYMVnowsDGBBn/oE+EK6X+vet/H86nOJAw25bmnULgXKm67OSE5vUKdr
resXdSI3GPzvJOFOw5t0rgRGE6+S3QcrltykIUxz1F9OjsZ+ck77D+It7nITDoAkwJmacZqexYvP
tTHD+YKAFQZ8qK2+ocD00g58iMpnWD8qJ/e3yyALt6EyVb2OGNQ0tYwGp8oN2bsRT6Cv3igCj1QV
1DwiKQPxcQ3vOyVhIY7fvoH7zNJTeu1R44KDvaC5qdFVp4bNxSW2UHjbYowYtrkv96fKAeHoWjxl
e8ucKWy3JMwOTP9b5Syya7rbQhN4FnYJ3trLKmiGkk0hKPWV/ZHBASxlfizTyyVMXXgCFrfqyg1e
IKqSD3sgUqICH1O/YmOk6n+r/hlpaIhOnBtSROTit5A744qQOzCuzDohZKUMZiPj5ZTjuVNT3uWz
PRcX9eM0VIlsA4FZNiu78u1OEh8kDs2trHLtSOz/K2BaJ2tIw8AoFHgtA1z3h5g5Wi+znFyKS+vo
AkEzwvOnIYamEAdAhtYI3s1JYcgVMnZau4GeoDsI9Z+RuwAxi5M+mFJ2dzj9v4GQHTZko7m27Nvk
GHqLWi3QmkbXHM/D+Uv5uHvg4hr36HBUMTLcshjHSOjSK0fVIpBJz0sUAlqRuF1pU1EAk9rJlSGc
P6ovbIJX35eL5qyZac+Kt+G1kTbpHTNKWCCbDfWOCS7km9qMaJGEEMuzeGUnHF+mpt447COIwoBe
FV20kpBLxWyjnJHoxT4D8THaNcBLCAAlha4GamfzVksxeK2GP8A55nIn4Ws4f2CE78laoOou3R9O
bIuuvIvRKPn4/qZybX09BjtrjpNeLGCA44rgvmpbqNaz2heszEW0ytQFULSurlJNiQ+x7iZX+7OF
mpzcuyo4g5ejPD3miwFP2hg61rSgWgKOFIC6ISnGgjLST/5WWEI31Juy+FwLZ45quijp/1IojZB+
+rfFu4LmSAvGLZlLh2gRTbvfE/LUX9S/PPR+b00M/vzIixnCy/y/p9ri57qAMoqz3+dlXqH3Nc1A
jdPNP6lObxKD7xd9g/eie/ThgDyuB8wuvixOyqrwaaJI9vKNAoIa7N6BTOIWn4SlnykLnF81VopP
tj5mlH6ALp4h7Fi6e5nXOP73In1cRwY50LVa8TEmucZgnQkLNIi9QMsIe4bfbSuSSnEmz7cqxN7p
keb62iyTudO0rZBRcJjlRrhWQeFXYehcJeG7OcZz9cdfVFbz9BhJ3ypThA+eOGgiecKQcndhwl4R
xlAxug7Qe3LD0YDGrzufMfnkiLZz/yCzy5rx3nqeiGziU8vicfZ6WJc25fUZiAYQu1gmCZqGQxL1
27x09/5vhrIp1QPyzC5Ot5TU+OJpxCQfsjXCliR+6IzyLmmAWJ/KDx4mbS3L0xSNjb+oytt0OGcq
lQRoD97zUkmCGon+x9hS3UZlZ7ln7SaS7WcWIqyugB9193/J7GpDWaM0f64EbbCzkUbV8oTuURXs
w8ve2dNCx9ZLEOvAsC1EdF/v89wG0h/oZsr4FXCNR9oZGIKwq7LHUgRmKS/CXXIj+sVoFbkMVfrA
UudJluf7f7ohXsluW0NK3vwkmFFi6JjLOjgpQRv7oTPzKhd/pRUzuy33zRlNIzy2hGuRik9s/ee6
yfRwN8P1C9yb5QVKOnmF0bU8kAJDQuCy0hMOA//RM8oeDVYZxUhb10jlUd7kYkhqYk/QVjzp6eu1
nxRHXqWNtTpFWpz6AgMpzrmtwPvKGKKEbvAb044FLxUibWFIK/ikGBGiJANB0D74iHLGO33hVKHi
6ZKZ5nzvyFh00sihS33ARlZYc5o35/cg4nQh7gwnKywNtWMDuOsXrk7HKNjrW9bKJ58I7jeA/AaI
hqHqzuPF3WU6E8FZbd+u18dkSoq2Xeh8y56czYe+hwBNY/MXA27Lpy61mDoUCirIPmIVG/BxOSdD
QPz8jyEBq0L7xKaxofV74ywyncwXl6roEHbtvqmywUdSwq3MgF8+HD27YQBnivumYEJal8GZROTn
GrqWlOGnTlyJYAw73+KwiVW5Jf4QMGuNT/8T5otiGGr0TLb85uEGv1yqAUBYjzuPcBVoooIU/mFu
vrak3LblCNjCRcW0ET7o6kCD4Sc1yrgvrqhwxCzp2q06E+0Y6ith/pai3VGF60lyIdf717/cKk4N
mG5RN4ciCn/JDYEcIrDtg1DMuAF8odxkC76X3AEsPxQ4aYunue5kxjc9aszkLwvvNKG/yfoPdCtF
HVKMvrlQR2gwhmjwWf4yL82MaqWOn1Vic0J5WHwGemWxDZx9Yfp2s7RK0X6zdRZQgwDBvYBWRnXV
A4GSjbdMpRfxSZ2btxFQZQne7Z+/tBCTdhlqcQFUIpeQZ8DAkzPZwKChMzKsfyBZKLCy2+JArTZm
gyo5nUwLi4aEcfsRwpIvGMkDyRRG0v0ZGUq7lCtf3pLg1qBWV/TPQ6ACgqCJ531Vmij3/VB7fJ5g
xgZ07OOBYowuwI5TeqPX80RQNSYLs4bVhwAFbOtVz+OhPoHglF6XDh28QDZHGnxa/7h6KP3wpCbs
uNIVwIo2WuCNdJFOAyfrVxunQMDx7zyU53mSE9aYs7Nt2k2Dl/EJJrzu8ym/pEKG8me72pnx2z17
/T5M0GpwxVHo3FgwX4ta1nWE3RSJBXpL0xxC5HP7Ob5umrjMbthaV2jY8+Kc4t8yrK3dQ1Q6NAMV
JR85ySlHSZ8JY+g4Mzxt17n4L3fU7xvnsJvHaUcDMO7/iRFnineuApwwNEMomWPbINa+641EQLry
tU6WKrjedqHym8uC9sI1VqduoLQ80wZkJaePeiDkV+vY4yPjzr3HXwv5aLZ2avvQ7PMvA+56CPj3
CPxG1aqYSJ9t3WNpgTceDL/xC37Pw87RAHfBxa+t78NmtOPp2OPgsxUcAFyAeQTkPF9yXSEY6au5
ppjX+8KQgsjfv0wgyODjSJtXGp9sUDmpuRtymU5wBvOhwcDzSmwjgRrAiurKFabrg7FouxITGZZR
ldOPA1QSHexQ3F5WZpERykBtqJmusC0ejk8j2T0qVf4mPjNM8qMF7WlFhzz8pADvdIok69xRGKG0
noS/wjru3Q0UHzFNqPeC4GT1thsIuqwH1OeNm83JVU2Ax6qrhYfhLU/us8PmXHI2+N8F+9S9/wKx
E43mrMF8+uSknBKrcvXv54Mz4PblAApNEViK+/SRRq6QTn2BZ9tgZAmKCMrQoL5seTuUYEEeYcXL
N8hTDlgJt4MFKcSy3Mq7yeG/mIXwXl+HxQnEEumtJuvOXonWGDGaUP4mpc36kDfvv3xMEsZ/p/cN
3O+i7fBiSOio3rArozgbZbLucYmiqpA5vKyN8C/rpz03Ytl0aNTsIGgHPiX7OcClnMXL2YK0QLDn
FDrqBqqwjvPOSuy/GYVXtqsHhBWew8ja7O4qvyZSuKGS6V1UD0np5dl7uStjDpm57/G9K9mdwfiM
EnTxWR/er5vP2F4DHDX2LZhevpk4br3RG5kbXzgFa9sO5lHSDfULjqZeq++CC5UOchxUFFmf2QTz
aRImRRSisPpIc+abTIXXkj2PJqfWTlOsFYZbRFbg/tHUMDdvXMDWP2R0wsSDM4OXIKwhuaDKS9Eh
gXbTILVStlAK3NCt2UjWeHE3cEz7hj2XjhAUAdbdBGqfg27DIKdryIDH2oHcXwt1vzHZG4RZ2nli
wofI+Oq34hsT1w9KXxAhoIteqjVEdup1mVM0xbpxP51NW5zouzrcQNTVqy5hDog7U8vbuk8Yoc5R
lxUIMccmHGZZ7fI3nzNyQkgYQv7tyUyICvCP/EFFXchnTEjs3hAUlmWuapS3lk9H5KdDAn5x3QEr
71JlwliaS1HAEO7PeNeaBdv3CdJU/ZeEzYf+swMFCb3tPlJNH+au0nKKSh4HH6EGKA5yZQH6YZmq
avKyTZgMwUsOkvhWlAKJ8NVpod6b8q0Yv+VHkHHHKDztv7ApX2JyhC/0CJYGag+21NuoFsfeC6GW
xjJS6Z76bf5ULEXm84OEHArMt6O2deidy7BhHrtmAaEd8VLey2Ll2VCrw4+ayXY4jyuxofLIdxCu
nWLLDme+0mL/clnZUaVi18erVzXuPBrGFuABQbKmY8IYgcdLSSm8OLMck8n7yLu0GVp0Izvkh2lc
3XcpMPUWluZRDk7eMxwsVcaQWwIKh/nQk8O+CEGH0NlL9oehjeKeHUQ4XoS5q2xispKhGilGoOnb
80vryr0evvOOTZQk6awzqjhqbgwgzpH6PoSbJuy+mydj1enS28dbtTrhuO8YlV5czfDLdm6CVmIT
5Mn5dvkkPZ4SAmEhVWWQZI7zT/boproO3YUL53Md/CMJZrb16TFx0piJyE01uiwoz6aAOD/4Y+1f
lb/ehcHg17JHAouDJbirFWoHBuMsHX9TgYatBqVwxAKU2Uem+AxbJUDhl9tE0smwsNj9PbKX9/Di
iUBUGXJBJ75vOyHLjPhRmQBXqzZxLTa5a633IHJxUvJuwjC9ghdp2cDZK+Z+xtszWFT9ZZjF0avO
U7uXjZ+7vvSMKus1As2kWHLvPFizn6YvGCxj4coqA2H8ateFZRt0+OAjMBih5Q5p6tlHmjxEA/Ko
IwKDKHDvAtNsGUeA+/EjLiOqcsl2i3WUC4RpEEzdeK83lqOVE0jDq1VM7ZTubPFKabbm2GC/s+nf
hbptEq1b+wBjfqxtctBwmWrr7R0+cJOxYTX/PJKS2JIa31hlf0DO9sd9ebUiHM9m8XXBepFAiVgy
MBDqEwvai/GzTcBZ/na13tYTPqcV499/K7nOctlmVNuV/qet2NOv/AlKCMytGJYmInHoxa2Rkol5
gWXs0gil+0jppCisfDC3hsqc3MTYrScV6ZjGlZfiNj/GIupsL3tiX7GSDmVdlwvXHz+dgpIPdptJ
Xs8QCgjxeKqoW45snQ04ia+irnlsIzJiy/cYpXIR55bbIOnWcFh3CcpgZZMtGDj4uyZWptr7KKly
jaQQrAyiYWxzterMbM4EPHCVD0bSYF3hvEYxUhy6cH7WBRNF0j0ocWxst++UD1OCpzligkYUt+8v
ZNlF0DI/3NZUyLOCEC/OdFCkaicb2xsJ37IIdpAHJ7qkd1ooHFIs9m/OuMqYQpuNugXqnj9PVSYY
x4ivhCyH0cHqBBTjuGIovEhAp3SVCmr1UHzFXeb8A3csutawh5CBhrW3pF+3v4pVTdQ9jiXjFvGM
JBwNDmIuCRvJVZCC8iZgTh33HWDTpv+li3teVGU8Z1jZ7ZwKzFdxProhzmqzlzb8wS0oy+5R6wKU
wT2WpEZgUN6TW3NDnE3htGv2YiEp3wjQLSUeznC37yZbBaIzor+S4ial05m0sTBrKRomOgh+wMYl
SV9b3CPSADLBJMYSrmo9vnnUAAqOgAaGKOoY67fABkK9R81D709ltTHOeHoNdG/XJD2/8WTMk8zK
w4fHko2IEyzA2B6Um3dhsRWFKJToREpFUiELszKkpCpabJoZ2PHZ0P8mUt/5F9BJ/o5mYo+u7cRo
TnlPRaxvmLblYapkVlUN0f3amPyNTHY0krXbCh1bBhoN/91/N0teOX761ZeGkMw2Sus/AIHk79Pt
8WYiQrDNrzBA/4UiYKZlh0sx6RFP1AEkYPZRX92lZFwus3DJY4kaZpdoxYwWeRgIDYYgPwR7oC28
She+WYXH3BHLeR73+8bvTGX71qefMdGCU1lcM8nguKnbiYkislySg/ntO8QVY/1Z5+13OhqkIRlQ
Dyzgr6U6lV2udDcoBS4lwi3+6+lRoW/r4b+wGDkpdQy21tDoHz2VDPQpuB59dDzNWsqBbsrLFM31
2aAtC5osqh/Z+VbjFXla+aGaDOCwdIG+gVMlMIc2oWjMc1gb2sjqAqtL37SaR2w2UZOmhV4XJGR8
e/S7TS+MXJvt21Y0j7NrxnILzWOmJhd1oZqJoZ7MYTmL6mJhjB+YCa3tIdz8IPMjVGG7/PAn1LR+
uKJUYBRHaqml4rXi93iPpmsTeFdakwPW2UV5IlwTBMnudE2tNnP3ClKyfWW/mWm8VSrCX58RE/dB
B/VRyt5ZlfU6J1NC64rzABkuJlsNfqm5JHVtZ31Kb1kPbJQQNtzRQgJkdi3dRXjpsvkdFOesnf2j
Y4CA+zd5yAXMXKbASo8DzG2A1dOAU84gwdfnBOPJVGEXYQQV5/3lIi7/6ybAmLcAs/8v400kog0D
bY6uiEmUi8bQnnH+vQ541yS0xN3N/+dqnfWu1CTjWwm3zirCr5yx/f/gLev3YR+na6qQhIVU4lCS
C5NmQH1K1tMNZrAHyjdZQpctdvhG3GPKeJR2+A5ijW7ao8NYv8geb4mB96Dyn06eGByBpIgu/JA4
qPrWHnujdjULCmZ8oZ9Vt+sZ5bP3hHZGv7bkEd+CJMDt3HgGAIExmWU3j27hDySE+sUo4IDyTxhG
VMN09owWP9SZVR3oEDxOI6NZZ1DLiiYphAdaV/FmxHlGiftI7Ddb+Cmhp+P8eU7JGQfPJYTaq7Qx
183w7tcnVnuR20DaIkM+RsGCA9toXCs5VTJYloygz8cSLv3kkMTJtygVvZ3d6XKyzTyd/N7tO0N8
KjRgBW/n/cilBuQXWODVmey0kwH5m7ppFBFSSviImtcFy0tAW7hT40x+e5dEF5QwXHepBEttWFmk
MDqK+vtrUlm8RFe041uI3Wc0S8IItYJyqQ5AFE5xFENtU9ZEnwpy+NFgBbSCEBPWruMoeAHq94qy
Ck1IZ+ynqLPR2fAsr/OfhLqGGNDtXw8m4UvyhBMYCRIk8UPIq6l5vKMzPPfq8GwOGjXzK6UBNhF8
heOdD/M2WJ21EpAYcxEf28nn9lVVlVEWStFa7KpdfhIh2rTmD9P2oULjkPAxPVQ5avWlojy715fi
jxyBm4SoCI9rFNqO8YuAyrGDDxqertwHIiBSRrs1FgxNFLDWkAPR5/ZQDL8T7eOjTPvjs3dA9O/8
kSxVF3o6Yb35tBVmip5iZVdYzKvMuCRYgB+Zdsvko1NwbSZk3+1SyHJJK95Fcy//ThJRHx2khSGU
FitltrtPQie7UwOlfupfM+C1TMquC59VISH1mZ8spIXr/fAIIjXsdcvQpKkNoLNew1sUgnXYaObK
rnyX54+AS3Fo49z3JCLaDvcyctUk+DTNhFAiFZlsLcJ3Tn4phpQaqrIO6QjF6KTDFIto2xiJPTu1
KCNgVrVQHAvJYoIkIjSj02CBcxF43YOLDlnX6PveqA2KpQQxQHTLcIDVnnh9vpSATE6hc4EhRPcR
fIXw3hEo2ypMign7IEoZvsJGbPgWW0ZUPjsQanohjbVQK6hzVu6CwJQu7gQyotV/7JftIqUwIT9v
TNCsdNZ+/OFTodrGyzeSReLc5B4nNZY+ivxwOedlGxDCNLnD0lagOCQZBZ3DkvFEEHdygdQ+lvM5
uRSfb8xaYPg+YwxRLyWN7wqFL7Yz6ulcR9rVCGE2Nwtu0XTGLvkMNLC2W33YzulPJYUHHa0SuabQ
GCAfh6/rXiPpBO2GkUmXWkCfVms8yDtzCIfct2tmUnL3bN/5L0B/QVAUUjzXnjPiIH+4RLV9VVk8
BQdAJxSisiU10z7fVFEfSL+t+iWa9lWwPTKipm8aoTANgPSngVX5pXeAb4oDO4giUhiYF7RJTwN6
ANEfxfc7/y09uGz6LIJN9GvjoTKLwLEaObKCZBG9NF1hRyVb6uAYTQZ90M2N+c8qZnfj8T1csaDm
2NjlgbRO9n23ENyjLflinU38LTrMycm1jkibjqDwf6ya+eRhPnFakRIWEvqv1sIZqRl+yPZxzP/g
D1K3Q90uGFSG5Q1TaOKvshbAmeOIGTBJLLmxF0lNN1EKSIIYHdxGO9P3loYmQ0dvAp8KfsaypBcd
qWguOZod6cJs/jHd9/huPPFyyEZfkmCyN4AhDOclW4+jjQ5gnDyOiUH66/XrEP7gzwy4zTnuljm5
S7LiokVmhNrb2HYjrun/x0RpE0Zs1DUhdAzhCVSpqogEuk+BvZw7+mn/O0Zrji1FQSyQK/SSJfot
nPPJWFvI8NpHWQm7r5TomSBpZ+fQkoZkNIcu/iKG9zQWU9vF23ZVRBnAQwMCsMwhskUznpyrQ2ae
T8Xr+NmGP4/Y7sh38DHnvMR1BQhGHiRIEVRKS+v75OI96chIjMCeio4vW5vFDqIp4NWIPuzi637k
7BjDitrX2/8mBrpGYBm7yqDM9Nx/AP8kA1HyaKwWAYVzPBpVKwHh0F1HSkBWGicJ5ASZ6HCrz29S
tvrifPmuq5cd/QSwv+boOBEByX4nXTc3elpgS71e6u/cgwNjoBiexs3Z72Om60lDSlYnzDtdhsja
VRFrHwN0Aex1soiKwlFG5LoiK9Z55DikMERy+fXMpOBBLKcBFth/Qxj6hk21FBWvsHzapYfmB35b
+uqzx9CHLWmnMMxcMiTDaWl20b1SWM9hZG5RFxiYy1OzLRiSoiqFUi80mqJObLt8u0/ETgJyuHjO
WLWAUfghvqafR5LW9J3mz1M8SHdSisD8lBN/zDv+cOkXMxBQN78f4U3hD0b15OpGa7hS2C5NRqpH
7CpLv/gQmmfP1JpG07G/ysh5bLqpNbm8HBA2UgfraDngzZ4aBe8k7SHuSyn1ce5f4CIg2SKUdqb6
jyMb9WEyXpW60SJVIsFUWpYq5SCl5M/Q9LzT8f7GFneNqxgSRpTqGH0Fj4ed4aikMkk1uZUgedqD
wg9zB8u9njY6umjC4eleSvNU4xJQfj9E80ZxS+dnJsDfW2q07fZbUw8e91PpGeClueO2PCcVabgI
W5WOWwUFsZaHq6ysINPOzG53ZZgxB6fQR4XbZhXsGy+eE/zAqfJM1XlO7mIrEWov9MJhdzHUoxGa
Zi7e824IAaSJDCWsVtk1+mQaKnSpYUyFHKk98ZCS5kc4hILqZAQF0RJaL0zKGpL4/SVv4OhZGX8X
+ZXHfd96iGL4mOyIWZFWglkOMbfSMe2wGYX1SCeegyI/aKzptav8qorx2eIM3h7mu0F5O56hZOWQ
OrADfrTvJyJARQ80MzHQCD0EozAzJXG7myszqamCutQ8uHbpYiRa+fmHfYoNj28rswz0MlP+Wqx0
n5XW92Vw2pEtAe1nx8uo39a+dmAWlQOhN8ssk3NMsX89qL8g5zq956ydTXzrl4PyO2AeAfjor5yg
mJCt0OvIHXSViBdI3FLWhpthBjm2yjWnrTEtz8w8IM4y9VEMVlALMIc/VB08jG5i+xPFxQfgli2i
TfMYIdsWCQORJfOtBJZ/WzLYmhFh0X2jdoMno5hbOQ1rXc3MCE3KOL2cAZGzDuvpvnxxakVKd1dt
SpZYaeEpZSaCipM+Mk8YS+O9Q598vPk1FRrX6nUIR1CCCIDijj6EHOhButFXF3HPalN/TAg5Kvr/
g3yk/PvtwfSqdWDx75asTez7lIZqtmMYEaAlI4CtIeeT6DrsW2XuQgYtDBKF9ctjx1hnL5OcjDng
FBtxg6ItORvf5v47+lbc+xS4Pg26ntC+cF7Te8n3ROglHhvXZiGG0PhhCCAtnbiJAWzdC8LJTcO3
mroMTrJxkTlnX+RCKuEHukt0OXcgZWmjk3wN4TrLajFLQSOhdVKHl0Lx/9aIjvL8FWmsgVV6LkEx
TZQdSUzaqMuFUOshMUl/bRDvubAJzBarTvTVFJa0cS59/kwtZPPkR1VaNXgsOr/tsfRDFGf2Ti1O
mPUBvD8V7+N2BERaC/kTHAfEXQsLa6cEa+WHwQnKdVaS0bdCDMxrw7fvD0N8f1PbnX2hmSWqskFm
s17CSFI/xcCr+NSWmZYqeOgQHCUd4sQCkw/l/i9pOpGFr6ha7SLM/eESgY7fKiaiauz8+bJXng2S
u6hNvxSsLBhIkA4K4DuNPK0G75HH4MP7xk6mR3HK4hVNvF7irS5W3o7eVAmDg1rSpGNbpFAolrFw
I7Tsbc5eegQ45zII1uBYzlHU+MoxKokzr1ZKyPFSkDIRe21RgvNildG7gwOzI+Lp7m6bhtXf0wMj
MvPefTNtK8replBldG2laJupKUH4LmZDn9IWm3gSV4y/QpNL/NPU+RNgsFNHgV1vwKV2xn04eiyN
e/Up0RU1PceB97ObTPyIopuOc/gOjcCkjSnR0GLtz1ontRVk2/5Ttf3wTn2Y/4cC3m81a8y3+Od8
J0FFYRuZbrDPUCpQY/IFrj/8FvA1DPdxwbyXagaRww/VSZR5so67TY836JV+RXMg8917AAHaoxsH
5QHH1KjaLpptYi/3+yj07u2zU5on+FB2XXbYjIbv1uN9dD8NhBLA/LU3E7IZQKaHeftkWxxlDPW7
fKbdw8sBk/c/n1WB1j0fjm1w6wQAiwOygkR3MqHfIlr+ElG9uil2BSek3lxpVto99OwRI+wdEIbQ
Bhl/Qqsgsc0QqsFMnGxcQn1JtkWtfeSyIWWhFMWPJY0TWJ5wCWfbj1LtPhQpJkW1RIGzpKZAZQbJ
z/DjjjvjZW7c3QbPm33OFAwzw5EnzsFl/AIkvhgcwc/YYFrgCYRUYwjD5Q6xemnqtmngY4k1o4O3
+iKy2RigSqRekBckLCBVQLoJrNvBbGHhg2maucNis5S7DxkVkTXTq6eRnB4LaiW9TRf+guL0W3mv
J4EOJ81IfcZzzFDQJBqdOvzLbG7sT7IjlJqVxW4Ltp0GhewKCJUN3JtS9ac14m5nat84VGyDyjWw
eLqW0PSpMoIaGCa9nVfJ6lq12bWnOybKruRGO6mANXElrCz0zZo97OzR7JUp3wHvIeV1rTdsFoa6
DIpYyKaxg+raZmb7tEle91aAPkUdazMSm7rznyE0KVdpfmpg/uQdHhDjS6RBNeyzo9eW8SI14P5a
U4N0Ix3PkH99+b1YFT9WOMcDQQpmp+hLc7CbucmkpW6kmXWAdQTHkhxCw09IBEWNnSp33HAstXna
+GKI1NqEP+n6CfZ2juc67Bngz33e432zr3J4UN2P0QyEXI4VDTF4HsoFAXLPzGmWNqmCXWGzdfuP
TdpOnfUTxl8/iUfJSefL15oytCRPXkiVMeYKJZ50xU/D6lHBXSVjon58rqbxObXeVAlFyzbxr0C1
ZrG1UfxOTjfxVQLcaHXTQ72IVIp+59daeCFlLVGUdCRGlQkX5ArtDZyCcLpjh+UUtAP4DJeDr/HK
fXwt1Umh/OdhVO44tcxmbwv+yoxfEVdyK1jEACsA9chOgWVVBiB0OXv1rNgiEJORLLKVA/LBsAB1
GbCunqaN1OrYzBm/lCuTnpAlhMaYdKtqARRiNvskeMnz+YIuUbKaHGmOja9Yt3XeAN6pzMUW2ATm
fCSdq5cjzzJ+HrWXmN/xdaHbUfaUjrjq2lNHiOOnAOI+g76bfl7YLcmhEEJZgLKPvgZlUdsFxpWB
EW0qEAes3rZnclBlh1NFQHYyM8oVO4jjBbYrb1J/yAo/BffS02QbeM4NELZlASFwrdGE29AmMtG2
siiCDTJtkkoR903ufGjZYZ96c7Lrw0uFAw+UfKhCVfaAqUPTFjbyjt9X+Iq4glmqxI3Syn+kO+Ro
aSMps0FrISrV/3KHpGpycCIPsjB5y+RjDI8bHHhG/uRdKKfSbKqCZScFbYVZ7pKfXSalwyH/Zzi1
8KEmMMAWxHsxhIWClvgqyRh3C/NDIwgKUBObAmtyzQPSasONn0E52vXKwzMqlwZecUrBDZ77lo6s
7/oO0VY20K0lxs6WB3bPXvlK/IcXVgHi1bK1htatXwE24Vo55Yz8JHpbA/CwC26maUDHC9ymxStK
CnzQO9zaUNNfSoBbBpD+K4Ji+7YPdrlV+ZuYbgEj9O4kqbE0xJVAg2u//YiNqk4pKfGsieK72zR5
zt06YRCAJYSdUkCMm94GI5cW2GyigF2uWoabukOD07i3oQAr3VfQlMfu/Ow3KUM3VHQ1mlaT7b43
3JHyoExe+zF08EtEK8B9QEsi15VVX7AxYU9fwYg0Xo6CWhC7cHBgyCz0hdTVTP/2ZfI3IXAMiVji
7EEwXBO/HZbcXneR6j221hKEcC0I3Nc4cNzcBPsaMwEAKCku4kwDxrb+Uv8rGOiHLUJMRdul0u9D
ObEgK8HKPtqIdArt1L2Zdz8L6H2uaYXr6zKhLFmJdKA+TCn4bTTV2qT6ngYSO59Nx2jgh22Jv5UX
zI5HJVwsm4pK5dpcQHnmMrakqlYXLTFl70cuijYR48vg9nBOiUyH/dsXXa9ESO5upZbSByFlyLDq
UppjQYDGvpsSnMnXaZIyTWZEKyrt4UDPmqNbHxD1iCVZ/CsCAuXvivTJ89WGIQOR9c3l87kOl7Mo
YfGbzw70mScval8MRJeTtDKG1sE/qQpK4mQ+/RxZbN+FCmuBoxDPMYk9DdiEmYbNFhS+rlH2GG00
fg5+HeMqnMOYzDPbl7pFVNCy7I4RfRNAoNM41igXne5iHWXUw1x+pevOiT0iyAGtjTCyfXIP6Ax9
NfYYPNr4zD/FX+cGaXC68kGLh6N3Yq89nxW455oGuQGAVmvhIPyJFD/krnjOznnYOMhvy5Ns5Y40
CaaC10+3zazs5xTUfVwJm+zxY/u62h4XCPa+T41lMGb410ISM8JgKTqHtyP0HTkT38J+bZ/GCjpX
xWSw/FCk2RI3PSNhcV1nXbtXN5Mk1dIGbeL7evr/DftpB6/FcGo2VyhSoJbzZwj4zCLWL9VdLHfg
SDTFGS1GVS3RTnhTGV/CdH8Eufru6aRmKg7TQgBRXLEKJ4gEcp9T1Dg36jDAyYYUykgGQ05y8vd+
96f+t/PjDyMHPBYEHndGtqEevsfx0272j/QKtjXCJF8Zpfv9Co+1Vht/rpe5dHwk/vnztUciU8+O
ZCOyoTrE5dFlNJijb2epe1xYKv4V0EKDDcoQAObhdM/+V9YkrCNlcD3MZHu85Ib/RyB5mffvs2+b
1fFW/XAxrZdv+6E9yWH8z6NZqV+2PFSZsFcN7bFxcDKDr/1D2YDthwREXJ44MqF9SfoAl1dos1Wu
U7SiJBf/UjI6tkVE9dL0prEorws7Wz5b3hykSN5FCuL0rC5F8tcATuCBNBF7kmtagOgdZSXf9BB7
TQbNnJpJ2NrF/FlbD6F1xkp2K+wytJcn7cgEXlePI1Qey4w/fgCu1doWlTsmh8aiibKvrnnVTgmU
BrhHKysLh4AMTHzVuH0+zGDvBRdumTQ4WeJ1cKJC/Al1byasX5bVuvVv9WzehyS8xDhqIuGL3FPk
3z3CtLTwRhXT3d3FhU/57XTuk17WCh7EFR0ORtG0lH3xwvxSJrPOY286B2miZT4WG5DWRGG+GPEu
tthHe5SyHgJPsbHGdZYUPnnEPztDgGvH5jTJgV0+oxtbb5zra2K7eK+kZy8Ia7WxxQfjPtGcRwBd
RWBzS4ZOvpmcmLHqWxwKLiCMeh8XR+iO7S7qLMnZwbA8If1Rx6nPpkEmZ4U2gowltyTgfbXUCKeA
7RZUPtPgiiKOMnR9ATyNOJg95AsUh7Ek/J+PRxh7u7v3ow0dmB4zNRdP2E2MWQOk1/8hAHy4r+v0
KC6GkOT9OrqpyqJqXUlcro/QwvV8jtTMlbB0dLqsIRwORorRRrkp4K+Ws2nj2mf/5UDVxgOQfYKJ
SbIJSahNE4CGSWiOgK+PARQH14SyVzKGP34J10VH99t8GQm3y8PApV1i+7hxsiv5Mi/IpGHYtKJp
Hm4lgI+LGbp4aQj7TL2QdJ2NJZBkMzJW2OWz3Ptqc6+JWe15cgctV/FjSlcW/aFkusT5EuCVzTUS
sHU/0Q+FhnIu2VakN87XKc9zPDHUYPOW1tdmKXFFPz8XOhy2C7DfD9vL9oAr3dsn032KsiJ/KsoI
2WVe0EUJKDWNZzdgr04jocCI2fwYC/B+cDQeM6pDvm1iBB+vOiUD/LMUn1XYMmvlPpYy0ODMK0tW
njyMgdOznIYYd8+OB2dnNS8t6ooHPwRK9ACg4IRQWr2EsvR8ckvYbxAGIe04zxyKR9BXdALmTd/F
OC/AChMoL5aOzHARUYwGCnPkaokuCZ6PLumHOoHeIhY4MQA+ypNsVfMdwRrWv7BBf1mzhFczyvCP
QwK7mqw+ei93aB5mBT2AtoW+FPDn673P6eFlRpqYYyCzvexEZAwf4K0G4JCwtmjLE3GbhphLjuQM
r0fMwMP06FqzKYFDUPjoXHPvqcm0vE2/PJerARGWkDLCJml4gFsWsIlUdOyqLr/pqGrfK/Sc7NOx
P7CTHNl3bcp8gJagbTYKvcEjxzW/MQQKWX9L+zhVXn+AHQd2stx5uDF7J2eG6X+63fiqyorTiiJo
F6Lsx43PEfspWPsIC+xTc/gEp8GiOi/fZ2YMbqPy2PAixOxtYrWqwdR3+zbY6Mp+lHoce0WYmcNo
8zNvbXNB2119pp7JXCdMqjjWEW0t8agHmrlFWPjr8XKVNTP2vaMBlYgO3CfFbyCVQG9lPffn41zQ
PJyzr0Tiqz+Gx7CWY8zsGmgzHetg/AvKNEuatq+3RuGgz8Xu5eXqYQA+2vaXjA4L1MEBfMjPGett
0HEL1n5waTg6yGXbhknWT52Jk8vcFKZYrzFFUbwWNwUABr8tdBrTsfqfX2bR/AW+YpG7bs6QN3b/
9t2+Sx0rVNGqI5H4+fUX6iPltcV/jGmVQHDN4kDpW89K0qi74ATSSKpeSjBXPmQl5w3lgflrXgRt
VquJmb39sY7gDAXBHq0yvKjHvF9/KFgMjvXkJbvsd7g4g2y2IuA5MT96nkWAOJ1LgxJQHsk8XIZh
E1ooMAt8Mg18dIly5npSFgYrTTlzKUjYILUNyvhr0/0TJUtBAGOP+w/e2Ny0pvoBUmlslQqh/fWC
AyzU82uW7K88EvP8cbEjSTzQIS3Kprt5tlwaplIiRKOiStcpwgPA8isPCNhL75OWq5j6gWZYC1pw
hkNuPWsHSNUExsDNeU9AUSxpirttvNAgAdxJjjPlrRgM1PrykKjcr38zfr4oYyeHJidNqfbxdVX5
vQnJZAfF49S3DLaQwqtXxIZTSObvOsNhGHKEr5Aly2Ad1MOdvHiAEyoSooZArgbRN1Hi/GaMAk97
e2O8xEfkVqRR5J3ZcVF1NJA4xjT/vQmaWz3ry9jKXklNnRma2g1jfDyzbYdFShPUSwzpsGbIW+IE
XfD0cJc2SzB/9IT1xMTmydZC7SOK5kbhJKpM/f97TkKtrmz8aIDjQff4NahdknCyFJoraqwpKTqz
yxYyxpfiH3Gby7iUYt6/BwWQsGO2CqzXOWKJJVA34WLqMeFRE4MVpwxHZpAHdDewfJfhgyafAqnb
7Q+R9Rwkn8FkWr+bWxD5WNofSppltcaGKHzvyMSgaGWfvRK1vFNluxgc4vEsAgeM5t6iuqvRGkW8
jqhSBeE0H+dqVhduCw0aPo4/Ez4OuaAqjwGho60gCykOJrVzMFzOdXTHDeLcti7oEOZhgNEG2GG2
e9ZafBrl9ja+LH+Z0cGbsJ1v283fnXUeQfmL54NlR6R1QyTNIJjL+duYdg3GKS28+e848PUDrUkR
ZPTMynGvbqWvnFU8I5gsE2XZgMFtn+HGZgF4NFbUvQiMco9bhrlbLaJDekKrF95z5GOgoN75cJ7/
/pjvbif98BRjmdIsZcPnSgKJzlKRqxq6OlXJYRWdo55r4JuPjS1vAMuZzKpobkuIi11cGhsY0kUQ
TD3MLXBuyKMvJooIevDgPhlhVTbDnBdEoMajAnCkrgkKudF7g/lCFszyGegRriYmSN/axmPWpmvs
CgR/WpTmI60X+BgLFmKIW5Q/gOptxgYprSPbrKuUH4XHFUE7yTbYtui/UjW24Te1wgL3n+XtVDv4
QvSBG9OCCkOfvyf3ohjOjTwRyWV4JSqiEFHj7obGWPrPH8b/kC/xlQvNgV+4wlxbq9uqzGQIXcVc
rI1n1Tcq0eN2/MdA49463pI90fa0g1MUH1yqgf7CCqff7n+o/IRrUMEEDj/e1ivAI3yvCw+q7QIG
pykGaUbFf5UDESPXVNUU8md8gJOuhe2A9G4T3cqRncPlKxyGAugcvyKP7i/9M/WYdLxymI1S4Mqu
2GUVE+Mj6F4bx2iErtq4+faT14gihwgBGzGprA5VI0wiaLKCV2w7ilOSkm0J6Ej2n7bjVv6fO3wD
DxhGJCbRPSH8nx89nwWv/49fap4p1ymR3TPEKrXS2rmPa60Szsa8ed/WAqA1gK3OXe2dprPLSz9k
4CFik97UT/HTGJAC4CDlLgI/Id7QlojgoMrSCiRA6vblaioE9oxijurLKcYygi1y2gPw2VSSoi73
R+zUszaw/HPDc9BX5qz6gozC3uE/twQXRWgglOusp7g1hpRMT5yfUsmIHLab4ecWQENuR9AdDNAs
02dv64A2HVG9bp8ac44eVJgHnCspgQfUHR1YZtT00VAF4DJjCKNbKnSrY989QK0sS18tJ/wafsHz
Ou0I+It91ufhqKkrSVTgFYi0Ad03Im+Gpp7xkPI+Vkk+i+B8fvpca445QbHANPN5dIYythPlpXUM
hO41lNaP1f/iSdkODbWERvLYs8RJ5CWApT5uSn9XgZlv8DJtCWev4w1ZpCLQ6Ou8GZa6DKfjA8SV
548nBmK1C1z7dKkMEBdSNI9xSU0Cnl6EmXWDNI+7MmusmziLGfFuhdSMPuRjCpOVn0NsoCTh3pL7
begfq15VwvdM149zlePd0SVFLU+drGjfB5OXg1WNGBefNfRrr7cQBP913LGVX3qwoDLX3JpDJ+KC
TmIjFKCtSHll0a7cLo56ZBZKrpa0nEpg8BiwIbOexfuxqEHL1KlxFtyO2ljXmvfQsGxuPtkw9qZd
XzjGK5ns0DHTH+2GFDDuihr9zPvP626AXYJgb+gLRgI5kpP2pLnKsXvHkoB8f1XX6jYpX+nvnyQI
2siJj5S11pif+l/HgSrnX+YnbrmhFhT0EUUYR0VGU1X1Ae6dzORgi2UtGwBq6TzTpOItjVTeCsr4
Em6yfvQBjErSdAx0RDGmkroi2hNAcl9lD8CAJKYN792522tdfFA0wPdLOHvd/U+dkLk18wFwscra
jj+W4Be7YMFLJ4ADx9+Ctajih0dXX1DJCgTGve5e5n4NGEfU7xaByFOOU7O8I8r744FFJ3/aQ2OE
NV/L2lhhiBY6L3SaxqKQ5/dbh5qzDKO15KFdGww27xkx1k4m3VRjtPxdXRWRoUezADWzAjDKR+s3
wTdU5DeVeQ2VGZdrXhBhjXc4Y7mjdY9ljr9nzvdwwdttdI57aueUxUljpXI500WessAZONgEP4YR
0vIphRnbL7eUCj+wcgwLtFKE9Crls0HmQ+00t7bDmKnLph7+1fFSEGnDVX964Vq+G3c5iGzO8Mdx
6mYqwHXU1jAbCRIMTpmKneeCvbOifQtUdq3ZJqoTctBazbmgEh+nliBIcQF0INYI20NJvaj8Wh7s
h9zzMyKRmF4+9VBs2U3ske1hmpKmdlnbdn4wB6RV3nhEXEgfP5IynZ//lcDJgWPz6FKgrph2qElI
DP7zORIYKEVLleNeuZG2ZQp1ZrkPrVh1/sYStdm4YyBUj1gYbn21Ct2k0cryqF0s+TQ2ATMpoF2r
q0rurMPwINEsNcGShNBAThPO8rrZkJci2GYTb+g1dPaShknRT7Db5oWGjAwiDpmFxd8SbZtX5cnP
ga4V8YxI+pzTHm0TyZr/eabDE909IOWuylHhh2nXpt+XmypdffaEWhUnHBL0lFvn7UDX6Nm5322l
BT+xF7WKszx3vLOZhgfAXrXyYM1qZEscvyvE8Pzh78J3q49+0P21hdi+aNhq382g+pyY3dwUK3sl
ziaURkNgkPoiYxdyr8XXMKwHf6FarCkUZ0sCm221FdZvBVujD0JOT7zkcFx4k8TWBImnVLS4gvBP
2yClm+jntmrqUUU5rzJrA87q85cP6twljMOlmJ00M2Mq3Etj4Gd0m68IJhi79DQuirS5YvVubRos
vrbcaCGWf2Te4L/qqNIGLflTdwtDH8iwfKZ4jWOpWvTFXHxJLf0a2TwGET94T1/r+f7ZnEiJICWW
UKokc3CJQitokzFNpAtkd14VhKuLV2AQExZfr9uMCXZ1SrDIhcrhaLbRbYuOjVCYeyk/yI/+1BNy
GqzJxx4NIuFBorEw51lkr7G44ugNRl7zoIFoPwWHAdxxYbxa80gMnQXktnvKBQCRqxx+FcY/K3ES
P+UZvcQWgUHZxvoPD5EqLpQZRsGgvYPljenLkcKhMQRubcrUOS/Mhtt0KW2BRl+nkFR9LZe2xLJO
061aVD5JiCKurv68t1SgprigUHCFsI8GTXfHXXqN6/fmz6PAA8l3IXkepmCspx1n0Z8kGaaNPks/
Q/PVe9V7NPmqWxo6QgQ1HygwwfY0WbFk2V5RvNARFHRigPY7uAvwMYc9eTtryBIwf5IgWtXeQ0gY
Mv45uqQRqtxR0xDoikAH3y9hhVMVRHfd0dYNXQjsAv4XRIz9eWZayGNDM4k88sAdfn4USkfferYE
IXRSnI2DHRT4MLVuAZi01/CV3KTUVlOWoXthB0ISZNcybjGYElp0+tPLK2OrwiVqBfPij1Nc25qh
6cWn4fAHNyal0HvNxqeIWqdYX2QrKBfXtf0p0wG3iFwDPMarMRjvfPVFDZ0VK2Vogtg3/6nTRSpf
8igbJfZhaTFLnDbfXTfP99Fy08cpqZVHnBOz/fYYxBwo7DXEoMfa0BZTAyqg25Jty85/kvG7pb25
PxTrUb0sSJifhb/ktbEQdMi3pPUh/cP2WH69rwxN5SnwzJbbZIDIVzj4BTrMjhzIdy1JNsbWwb/s
cohAGx68C57uGxPdr8/9FMOk6ioZuTzrHdks3KNRkdRuEPCdNem8HVvDBwbvOe1zm611mI6pZ4Tz
MROyJQvH+YjN9A8oFZ6QypI1hSENNsOpSIBaYY3r05QfT4opwcspHbMAAM6Ur4RprAPX8O8Q8Skf
Gw0HLrXAerapb4xt/yowtyhzypqqyQNWZrMz6d34me2t++avJ6ex228aYZLgE271OpQVDuKPwMvz
u1qDIKoHKUgbj92t8OBnV2I3+jaTibQXKO2EkJw37bMFE252kQKi5uKTQYtb6AbzaWUKIgbzIkgV
vRPBXCDBYuR2lBNw0G/f0nyNb+wNDRm1fvgbdMEWyx0/fycuFVlK9ngPet/UeTpGu4a5rWjxc1uq
p4kC6gOcbi948pMk4zFx1uFRYp6PUZkcSWCOpyO8Or6zMLYCVrs5a7Lh+w2C9aB+2jjzoBa2oMWP
as+ghkxe5kTNqIeNackz0qU2fd+WTH97cVTfiyQnuqsAMF3ngPj9NVvaI3HDpgKlPulqYhmLfTOs
x/RaxKn9IYuRmiv6Nct3iabQD02WgjxGVTwWp2Jl8Uy5fK30S8Q+VNTQfVMvffe/P/oxfqXWzE/S
5T6POFVZFj4WVj6IRVbqqM9aYW9iSdklFEj8hTpiAYk2yK5vcAmDpN++tGVWL+ye41eGmfOMV427
mPEX05M6eCy2JtjfSBG5oVzONoz2p1YUgmc80xwzvvWLFDKBZFf6Y3m2bFxAcJ+aQYtwZDBoeX4/
+VnN3y08F/Quqk46Vw8hj823hu+Bcbewivk9hP59RSDFZ8Ryv/evto5kaJwpeIhDSPPX8TW0iq+/
1hZs30uPbTQsmNKnN6Z87k8PbGxTjB/F+EYazfXmqZJ6P4LaaVsui92FldCgK6FSuxZieP932xRJ
4P5orm8DSETRA8aSLZZh0WlTFneLuGYganWsXYhKjf/5qJ+NWdPKIVAJnCShkxXOVk7KLG3IVXD9
PLMs5DttNmWmJt4kR13tyBNzd10X7QQw3kiVJTxv50xZhGaaqh+1WWXrKiTt4jpvKzNHLBRRsN7P
+LDEJZpkR0Ly573YpvTDrn0GdAGU3TJdoYU18jBWm7J/Tguq/WeNJEq54Q6rHXtUzNCM2f+aLen6
3HYUbsFGjSC6y3Yb51h3hWjIIugLAI+spNImhzKslDxsfUtxYS9bmZt74YFd7gAwQhvE2osclQB6
0VMtETqqEB8ynE0wQi60jZaKRieiPWOK/5MwypqCHsy6TIKIqVBxkl76VeRvQ6tyjqHmcuaEaowf
lXfxU59ScGlFwQx0+s7WKevDmBri2Z56/GN2Iprf/Mk9yVAD9OzY3h0GmQJ5Qyr0YoasmdreeE96
w/93Mb4aFxitmE7Y8//bznhQBhpwxftaV+55idYpS7EKPmS/YKhINqU5+F4wAvEV5jwctsn8key2
a+HqhGpVx/WuKOFccvMArNjSUiiWygR7M/MJfCQWhInEWLOqNZ5M7ZQRrFZtzwJ8D+Bm3AI9Kmes
sjUJamS/aTajaqiQZ2XKYbvaLmRQYVOtt+CkA6Wri/meeu5LhjQ63ZHaYv6i/ru8BhtZ0Ho2dLtq
H68otpTmEhuqqFn7txumkMRcmSTHV1HgD9GXhBNIjhmMiFsZ17bgESEwM+2n1LutEuefk33ReN3r
NKhMkoRny43Z4HSDedyWAOSBV2fbPRUa43z/2p9rDzqS88IdJQorSw4rYUsLZzqxKeVf/AYPyObd
mMgO9NrdsaPLEEBkr75RNBReSjdiKWZrvBiTzcMVoKYpX7PklcENzdw2SJbEryqE3nVO1yFzaf68
CLhadeM2pTC7+I/6WTQu4zNGUCC/C3um+l8FyaMr82qVCtQoR5hfJh6WROdHinKIZDMpJlB1YHWu
7CGjjvk4vt8kwrQjVgOAFf3IXyExGB0c369AjtQYlJczFcXxKtdqJK+PkZwSa90CGXu44tf0uzAK
ugIrw8dIERrZ7PEv/XKeb3WLwLtchVMStTKqE/PxIS5NKuv22WEqZBtpljXCOjG26K3dd2xV9ZTY
kBruR07bv5eRScEn4Ixm8nZOaKDcgM9flQOmefGcSprjWDCU53M58xoG0373IdILyhko2dzQ5f41
83bwLkWWZ/CqkUxJvxQYx0woHwGO07fhcwUALIBD1l2F3YjPoQP9aPeFo7ctNvAL3MOCKsC7EX+8
dua4v9avDYsGCR4U4ILSzewJlwtQjMKEN3annmnNSFdMKYc7AOBV+gHgWei5Dge1RwgOyTta0z/T
KAlvRDQFWPw3Ha2RXNRLollHPf7G3iMPfyMjCVVYvICuT6fpnrf+gZDvDVaWfMSiSVMmvddbhmju
yGAglS9WNf7kcRl8ILx+zgLzUXROk/mEJiw8/30UOJhiyRBE3AZe/LkzD0DcjlT24InGbXESVVb5
/jMAGsyhrTLfFgMuH6g6sNXeDjufVBIwO59jgidwLju1HiSsgXMaJAIROLxnjvXeoTljL4aDTdZj
k4U8uaoTsGtwpVCVv+PhzU6G3lT0irDsZCUnMG4fJ4k9IqGdY+pK+eRMc5JQzsbkTL8k6mWfOMd+
48aoiG99Y9gDhLGVItFnk4+RZU8Vx/zYztnnpUXiiz7ZiigoH8No3jTuG4RPf+WqUglugaZJwp+2
ZXwjOjN62E6BrmpIw8Nk9C2P239gK5rN7waLqdUZkUtW1UepPL862FIgEPM8baLsKAxy3TxQVThi
GJ+duRwHIjAlL/wUhPoVBTbHVOdHttWb2OiQUkWV6gR2bFSpaA8da0ij8g5QW1996H8Zhml9l5Vk
ztKv7JToKkmgMbzTWQsfLuqNyVjJ56QGeHonwTS6CwSarLWJ40JjJrE+Z3c+gW1w27gCJGaKWg/J
SyV9nxM73ITlrnXnyvDO6Exm+2OkwGWB9nnXKvaquWtkNCS0cbzuUbBOjeCRPK/I/40l5q7rDMZ/
vRnFOfpkcHFy1Yd1Ob3sRDKyw8KpbsViL/Yj/vdKz6SS6IjILAjVPr4w1G1T6YcYogwUwSdZ4p4b
gKjbhjt/EhOTshjrhQ9TWMGBnzsu+AKyUMb0bk8AKqi5PibZhWbq7jotrN/u5u6L8JxBpZ++M1OE
KeKPWl3sauzborTHn9KU/AK4gWXswhVeZ5jM6aLGZnEC4ZjlA0P1+KeD5M47NLuXOK6ONl5UezAa
WSFiNhSrBRkonieRwRSvygDq6lkOFNF1bXyq/skAoGcLx41CreJZ6V42ZZEvjs+yt37bK7j6x/V2
YIoI4oZAz0QNpXfJoeuaXlVmouoHXM1VjRyzJXaMkU0Ny+Kka9J2JY5BGXGf384bIP2R21YaRtCa
NPpYFI55I+23UcltNssY5w4O54XXd1PbI3+Q5TBHNPplomwdw0C2ITyrIYyCOBH/InLjsu+GKhNC
c+YcYCAgZN6EnmESk6vNUUnw5tG4doVcxvLCS4tUmUXD1mx2zdPPKhTgLODKrceFnMkozybiVpBX
5uTGIr1e2Lan3kWPHJjoM9df6Vlf9KD0OFVk01h0OZFuTiI+E/Gf1VAiRAUleLAa/6duxpog9w8f
bsQVqGurmRV+jsRyolChT04M9T4VPQ0OuiezIDGTntbl5Q+7XFbrDRba7v4xq1sLmK7eolpMcOEB
/CJsxbWe+bIT++gpDVLOroZBSbNLMFkoXyr7RVDOVS4K/uXLmHOw+frtStHmtmui9Gzo6aC5jG3J
oK+LckcjyYh661hKBIhoqgRVCjcPdvYRwYvYjvf+TzkiZJiEkD/yE96WpgyiR7aML1in9joIiyYO
+WwA6U9M2BRsxjJRYXU8r9eHmQ49OgCWZZEK5MPRQ7vBjvz3d2hnJWjnP92eUauLcOBFvD6CZLLB
FiSQ4b3GOMlcgrBkWVCXwufV85Ukdv2HvujLm2QdcC1NS9VyDQ3a7YHBSOO6ioKzrUsgDNhmBarf
/q47hyTtEcwt7CCsDcuVfuhNuTZsovZ4VP7b4/vxPTppPfV77HUN2l+B6i3S5Wa5Cda+KLEAp19p
LozIp/yek5PCLcGfkOQlYuFIfaMKTgRXSpUJOqNbygecMX+iFvDbvMwd4VxPMucrcH51Y6OJNKvA
m6NgKYZZ869Xh3FcYjlMNm+OXjIr/l+It6hfCUjZfa5+ROUHNFUE7mfW+Limixt3mIZgeG/gTos8
ceXekST7uYOWDY6/Uhff2H7fjIR4eDipw7CbKPEH6bHwXcfiFAMpfY/t8tKbOqrALtw4KTorb7rH
XMf53D+yVFVqut46cyGlchR6fZUgOjqX/dua6q8mhojp/7WMKzSP+589d3SQFn9Ns9T/9rubm7kh
lnEgIXNpHD0bmy4TdeiwOFdYRffARo2kjfCFg7K/DEwJ+rKwaS4+lmUSRX2pkZnYyu5FtEJ1UmTc
ENepRqLY7ManHYSMLF0u8/nXpgAsiWFo0vY+KtiDG/befwUsVonxQ4HpU5PV8Pc7M8C28ooACwK4
agx72amRnxuK+6UquUiZLyCkcOb4WPysJyca+7TpkR2LtsmoHbRcIAg0+lyeYb1MFlD3HRpsEDCs
HVC2Y7ygHDPbcc3jYNXISpd5107J9yRkbHbM6LR46U2HxtJcjpmlztEHkBTx7elqXw9IdlD0pIHR
uB1B9ILwCbbyMZJKGRkZsRz7aQn+vUeqeQhci6AXsG7R1EEy5FpVep+v1mWfooMNoJvzXY8ZQp8q
b0hicVwoPHB4AQvXSevyOQ323lS3A6MWrgKyFmkAS+nPDX5j+qnWfMqbneWpGYsGC5/iOz+A8IeF
15LyHG8dbEq6/QEfuQRa7Mzd4gY/xCuHqIclI3rWhjNTPtedGBe0yWECIZdZBqHZZQdzeOd8i2qi
t0mbGVsjlU3XTHa2nJkMOtdDmay46JqEzfbpbMaCjRLFXjBYt4G3M5RWLy+Kr9ymU/X0LDj2ZNyp
ICv/Wyte7R3IvjxbK/bB+lYEmmhhTxYJ3uHudf8bxZT1LKxFsg5/JyDj+k08Z9aGFWkcKSrnSrcf
DwbaKbzpD5rrP0dsejsH4hCsPuSR3kF6pameE+X9DT2+TCcApV+sXr5qn9nMoF4EIeQ4vbxZuB/6
jgYRHYh/CEdk7pHXIM2GO3AmmhMWkunPIGc1LU1MP09+VvziIYGg4NZE+cEJtraQHseZVpnlc8xc
UkNgCwZvMqp8a6ukUVBnr/JiwowiFVlze9a62U+iTAzMQQg2CU/bNnS/FjL1cT1MRtc38oqUuFD4
K8RTSHT8e4KxysmElhtng4/XvfAEypQp5CYX07HOJwgsT3WmkkbqrhR5l3r+7x6I45QOtV53wQWe
2vWMhvBSVmzFSZ41OdpjVqFwjaXBh7d+0KjimpWA2qeBwKolMrIvzJqJDsluPxswyIPcqUxJyXjs
fTjO49vf6EnwaSz+YZS4ob2HFKo5s3nrECS+0u5/zEYX9I8vh9wdTyAYUiUkUi5WRctk+bAro614
8B+0jQ3cjhqYF0vydOtHhCnFkv5H9oYxw7ChxHpf0yJdJVAI8yQhqSYZ0RvflNOlD6GMNIYG+Q9Q
kA5nVXs8Gw9d4YI+EifM3CwEopzIHQ177GWXAZ06b7eJFcPQOY+cmFgivYV1514eN76o8IOd/Qex
07R3p7UN5xPmIsPa/PvgIwUUiT4tDquqmmff/R/G76/wGLSd8oJ2dogTIfXLoHWvg0ASsbs8wxm1
JLb1dGM8yMCrz6V18jdDty1aKBtsMaGxivQ5xWf1bFlFLIS9uZK6OFhXes0ksdD5TjuPzuL2PG2H
fI5iXmUtq6ZV3228EM67DHi43fLkWI81UDQ7JzCNWnEhJSlx/W3AuauYGOGZQLCC3NcNnXgD3bPW
+XMmsqk8O8s/ifGWxP8NlIxBiRHUYMNa0/No/HfBd01Shja+ko2CAxWtUu6cCMF66bj19rpwSXy0
pUVPQjDYEi9GmETlm+w91RGDJnx0xgFO/BQOEzVrB0MXnfEw1wd3PzU/02FdkP20k7ZI8FeOIn39
4qTWSvSNRsiMrWsxDiK7U6yStqohU4hk905VzcNHCOMfdIekIJzFZ6myg91EiJ3gmxprixBkx07L
wIt/2aBD/BveSZWgt7KKx2pg7jcSmS8GUPShKeu9VYgrdXsxu15MUUbdtES0nvekZaqQxsqbVnp6
VvX5MU2EAjXPB0XkF1LG/QFcdryPwAxTyqRgaLCTgMB7PfJbyjaaSR6MH3vDrCbm0IB/PTLMdGV4
GmHy1eiviVm7yi7EQom/08wRfgN++LYhiqRE65FZC3b9psDBneGIyubczjitVWkQ/d2QqrOjuqNx
n2j6dLTwRyOXxM6j7EI1fsqpWI6cNm46Cw2m1sxt716N2rx8TWJJqy03/5UOhbIEN0dvzfCNvGYB
SRM6c9HeAFLaok8OXem2CcjQq/lCjIBNHADi+EpyjAuTJs+jOGO2xNNW+Pj0JhKXBdQy9LXBn42V
qAcLeZe9nT3EpAzVdfD59X9CMQkvVFt3fXx8CCZpfPlF+bgWcWXsoBNcytM8zHgRgGw4pELcw4QE
AiCl/jKHKzXZX0rE9UG72gf3UAio6MA6N25+Vu9dB60nBjGddOE15atDwSTC+cfOEL5FJbr80zrl
A80SB5fGaQ84KT5GL9UiUvjVVIyUkpTDf1KCGhJc1rJz4zCyRtEel1sBfWddCST347J6iN4kO7J0
ZcYILXbV4uvc2kBNKe5AQbpRQZ0uNM3FDAZtyj7//IFV1pZO9VY9Na2ilJfE6xv/skOslG3Aw5Cw
sx/1JFgJPbCW6tIE2MEvyX3W30c9gK4GLP7MGcG60RWlJ/fKDUpBtwTUVtpn1mzFXZruBLm1maOV
jLMJOXxgvedFYoc7U0orlq4D+6Hmh1GaziU18BMzBXJr3V4/Bvb3rElB8Pkvv+sfIGmXogdTd8d6
wyr3BMRvilqH9ZnZjGpmWgIF+u3MDy5Ue6/IH3MF/YP5/DJ18Uc5+cVWjebApfUp85aICtYiY/M1
Y4IXw3zzIsncqOH6JIRM+cuD/+JRnkfL+f+HXWR2LsdWWtrjgpqeyHCKJkgyb/PKY9oRJ2HExJrV
oOYtOGiNTgtYKblcIpTynzFCaKXqSLDStEIWvovjr4IM/ihHMSqPLIxHO30ornNI7XHqF1u1/pOk
zxMaR2mYuAq3Oc4fHwL49iqXJq2GPAIkPFMDarTMAmvcGs31hjslaz2MyYUIWkLhM1wbnSHj6esg
i5KLVy+BmGaNsR1P6q95q8TTvIsJV6D6JFnrLcET/NoXSDQ68fuWp0eOwjRSD7xJ1qElvylUeXzW
2bXnguh+4IHMePGwQBBq3976FbgACBuTzf9N0+XWmM5NCvm76K3omYcIlyVCNI6ePrqD38FJEghK
V0wJRgGfkRIiztmcS+ogZw/pTuMZ4gwdwR3GN92PvgZxaJktYulPrvsu6uDFLP8i5g/ovJ+sCpWg
8NgYrOiTBOsSqZ2E19rFl1v2oOPWOKGPkk9scqCfAv0QzvuI58ohH4Z/azNhNbbYsl1qTPqqRKHf
ReMXhl9o82MxHO8Ov+qUjXNWh/Vf56wqPFJhfS0yCwSY1i2GNC5REw0u0wPHA5y2roVCbP1+btF1
FHgkyr/8LJQ+0RydiJx7oS0EBZaL3hTvWiaDHUMhRtU34UQI5IpFRi8QGNFxyo0NzmY6qk0h9yqr
VMs3rhGDvY1rdBxDVEeNhqjPuA5kigJ2CR0K0cOHQet5MQlLbWNbtbtnNHq3GI9Z4hg0BKssXKXE
CvupcA0LlyDO3Kz8FKi7A1nT46Aw9eZi9sD/2QymCijW30y/Y6wFKBYMnY3dy5Z+CE5rK87Er6Yt
nnRCsW5WstJ5a94n8G41uTDrJbDreRUNk/Udc/Y6zHZ+JeLWGQFCbIOnOh2zzq9WUERJW6jb7Mps
kY5LqHYpefhan128JrPdDPqNEFGixg9BjVNv2/dCVENMuu2MzQ0+WSVIwhgykZRo7/7RzhmUFVJX
Rw3rNd6cWPo8/EH7GQfSFjiU+aga5MsWKoCVeoMaHIxP7xAkWasn5pkGqetx2IO65H4wkHwOncxC
N2FJWXcWoW0FohnzVWZSTW8NL/q+YYCTHZjt14WDmAv011kBMaI3D0aGYNfIGisPpECwdtOp6LUN
GOhi3VX8kD8JIZY7n7SlZTj7hfFCWI9Rr0am632tEdA1qX6idx8T0EdEAkaW9VvDbKmfoTem73da
+2soO6PDbR6nAGB6+jaXv7RdpATha4wlYFqhvJV8Kcu83DJeZVNOVgy0pPC2+umWISx20AiQPPlc
XRrlCLatCN61O6faqjDqdgFrGHxko4v+hJCa+ITTRUOAgNRZ2GDAteQSFVgTxThbwOP3DElAkUI0
0FG/Ixawsz9i8nkDMFAJhkbTO2okT/1Y5PlAjtTuczF+uog/6QguczvRHGJ7kVznJBwsJ5QWwmpv
pgoxAZbUWWqCBqKAZ5LMtRAgSDBls/hgQZtNVn2JxBi7pPnelV7gkbesqPqok+fy8pGyk/hrlBDc
eN6z1xwJTPTpvHFXY+CHzYjGPcXAoPZH866Re9N9a1IAYWcq6V+6A8SbEN9M8u9fpTbugPDxvTru
TIoULxfr7HnGZNC6iOysuX44grIsmPks/F2esGZa6aVlZVI3Mf29PX30/osuBcto9tZsF1mf9ZMO
/At2NKEP8zW7LsayCF/eiwZTkMCTCabS/52e3RQL/EEHX8J87tEVg/gcdFparoD03YWjStuvQMcZ
jUUEX5/Ci86mcpHRq3Vu+QZZDdMpND5gpFFmcFtm4w7raUoz594PEqAGabHL5wlhfbIHStyNJE84
OjQwr1jxvIoRtRxmNH7z4/v1Ks9OM6m+p7zSOVDHJpYtJZBNn/WEx6QPsx6yLAgxkeBve6NpKUYI
x6ugAOulXixejjuljbRbUE2Z/LTC36LqfvaxBiYVQ0H0roO07VkpmcpjWta43y1P+5/kqY7e8z1F
h78pgMDlBpCA46fVvpj/4NclF0lcHTaQtidtrDfu27YXgC+y/Ci1JRl5TbPeAsn+pd5ZKphFwmTf
VRp8wkxbU0LAAOJsQyoEqHx/pIc2MPuT5LF7pYmaLLOBOlOMIgogn7B4sZVI6P3SveoNH3NAHNmW
3XRT39TdI3FqjqVYznVDh1hf95d3BIXubrAPu9LazCJg8IsQhb9jSPojY0AcQq+UCxft6qQhsFjc
6P3PuEc/W+yM0QvWELRnMWRxYG80uR2dzALpHcpWPXWfXsitDyqA9FKX9LPSo+a1smY7s/5L8+yj
OIIx/a+zGU5Q13l7CeFtMmSVPg856BCeTzpZF5YPIfBgXJ7+8p31MOn4tBZBq1BFiJ9gWWqqSXkR
YpcnfBpx0ZE8xSa5rQi2PEz95w4RZPI8a6UG9TIvtF8kfp7HSZZSEn9x7FnWamhseWTOJzRwJVZV
8STyxN+3Yeu/X3pQ9BMhbGaAhmnc8/uBvstcq3Tdy5ptlBRzhFdgKBIdAjDTRxNBh0+d2UpOrfp2
dD8TJ01Wh+tLTK3Yzuj/bFKcAGRFtkYQ97wPPEZbRQqOhRE5ww2Sl8mj7jK8LqHCe/Vdf8KlJ28c
Hcd1KBfIoow/tY5O7dwz83AbqYD4Jj69VBTo7eprskT7WNrxQ1KWAl8gf+aCqgNgwFGUoPesWUZp
g4hxN7Sk0B/85cWDDU7uiK/mCa+vzVQczMLt8zrYB2zXZ58dWwJAUpfTNL4t98H4+G4hMHs+Y6o+
vME9ll3tb/Klq3RA0R2bVLrsytubQOfb+b05ICRyfpT5bHXz6OIgE1uW32dV1hRH7sYL5o9ePtVs
7xhKc2TpxnmXIwsiJphuaWTKP/ZOhklO0AzeZuT/5T7bH//DTgrBC4GcLrtDyO6iQytC6vb85xlJ
9Ty/TpzrzBgk6fVkyqadBFjWvn3aBbWVyFW5ETiOf45+C3DSdJIujykyLCx+9rX1rSwNhkZIi3bN
YrbjEKCpsYQO6kUAMONs6tzuZLY1DUSfBl3kKPZsLYhCTu2cAnXzr/pk5HfEIir6/5C4ulwq0JJJ
3Gt2ZSbSKC+bbvGzUaDhLrMH1k0SfK2sLVaxyU1lcMztv7WtwwxaTZwZt6V1oXXMIvTxm+o5dwQ1
eJvqHwP64uzG+hAamXFfzKXeU63gHv9r3LlldoqS8nneiyO63aDebhUiuiUpoR2n0lwBWWQNyU4A
E8j0joJpDIAo6fQS814zgBMFfs8UL+xMrn3VierB5DPjMv02Y/mv19MISnIXGpq5E93l9h9l+mxC
VzwgYLJyKZN7T7RI1oWA/J7EYGH9SOKNTquup96gYP+9L+lUz18XtgSXIjhIzWedvN+69tnuBP7+
j/b03g7tvdjYfXiZEaYTU+9GYOVVHP/R9Gl+mfTO0Ou1wrylJsGk2P6umPUVjpEG908AAsJgAL5d
qJVxN6DjosiC+MGyW52edXDHWSZw5JIJU96I7pTAYJgkK11gKvKmwvtDLgbHZv+zYQVR4jQOwM15
5qhemQFBj2s6JbxFr1GyiD4pHXYOP1dYK2jPDDV3XMoY7AfXl3ALrMMYIO/Q0pIYliGECCNRkw1b
DOv/SM3SR8RdsTLXiNLdzMsIo3G1Iw5XfXugOby7JQwsfufl0NTpMRlRyoFuB7rkrpJ4BeUO5ZeS
jyVTs0nr8PKhjbDwmMl8YC7n5jidj2OyBvLJ1wIb5vc6Au3k0dmTyE2xgtu1+vAGbfWfGCQn1oGy
4t4uVSa2PjGMZ9a4YTVEnjbRBbFLH0+WceWkjktw6euetolMiom5Km7MzioCXJLkgkZGWODQZBEN
t4kFqHCv3EutEY5Doy0MkYC5FLlwdAMviMhomzex77f1WvgB6GZT88wrkXIm7UGKnb2YNLwSa81I
nZ3V+lDrQv9GWec6AsGQU8+5EBUtssMh7ej4ZQnUsyBmIPafWlb1q/doSmpgX4TD1mwRRb6KtgWJ
TP9/gAQ2dL3KsAUL1XFvtYBsyBKuoJYuTjNpGDiLg2R4p3hAAV0CEdxZJcmTqZxOekmV5Y2Yp6in
jD+KXVa2wOVxs3LVbnqACZAmW1DJtJd4ZPpFyviX+MI1uV0DBzloTWJ6iF7IbHWqdbl6PdMUTFuJ
5z1hTLxu4L7qtcbnpc/WHci6UdhWq3Ht2oK/KIwqAhekThlqUvhK/lT4JgXvkEXz3k1hipBeOlJ4
yRV2AGs57hYgDtppzB7SgNt6Gk2sRBmZuk6Acg5HnuCL/nITcwjBvTsW454eTPePEaCK/2qfO7Sd
d2D3dhv8D3DDQ0Qb2bhLEtP1RPhrD5+NF4GLOe+ud6tsVkMA8gAqUNdP8CuboHvvGEJ9kKu6EQGF
BXaUM/xLRWam/NqguDN8840Pvhv/8WhN77GBqCfZR5V3rFPyyUI+fqVbgdN9t/SS9GUGgYeCOQQl
mvjULLK0w72Bc8gYJtB+J98amRwTaKsENI1ghGFXv61RmCJ2vZtxhXyayKZrjw/Uy2drCyeU/AyM
I6S2tacvKVgoDbA1Zeh2EBCca9LJ2zI1+mpsiHwI0Ssz15v29vXeNDt1ZQJlG8Ac4rCN44NwohsI
GshzlFkLWKa0UaCrFUe9fThALU3Oxh6Ip0zGwy+rqzpAvolSQK0ZOAo/ed3dZCsQcGMZDWiwvO/T
gdSBbZC6qOwKfN/ymyp6j1bCGxax4XBNDxNJ9egOin8eLbjinslbnPGiy5qk455zR2GltRg2LJ8M
5LmjLD7b1zrBeQenMfb1R09rXvctsLjSKhN1E4/jFdGaqDgTAe4kZUYkdux661TmJ5wWdvtefMMm
MpO74sCzUqb/wnuCS3YGPFeveNnsDqTMnMCkRqA1CgEeeD1n6c8Raqv7fuFB/viWVyvsT47JrewU
3J1UdqEMreIS7+BY1/4kAI1sgSKdGwseVQoPH16OaNiDz6h6F8SAuDRrRG0UISVdmOqq/BQrlsuI
HxFDEFHFjcj6kWXtG73Vf5QXzawFv7tUODDPEmLwjN2OvFyr9WhbX6UGv8XghR/8jw30JYJzkWuh
JziEFmrcKCbLK85sx81Pq1Ih/iVHcubn+zjBSjQncquBSc2oTCuplCy1sSGan5DcZoEcbKZv9qNQ
b1wxHOvPGCDsCMh06JzIVyRZ/LyAdITTvMQQCC9cJVLV2w48/Uql4l+A4F+aRva2AdQW0bBO2Cwb
atLLLf/xw727rpf52+VwnNEdl69Dhp0jdvIxHJY8p5cz0/GKk95MA8q0/NkWExOLtCclRj19g7qR
6xna2DmrL3VDmCj2vSM8WNFHfC13Z0MzTWbuzB2f1D6Ny+rsiBC5wmAy8yZhL9hitnkJDyxy1p/k
Ualjb+wIlGxZkfFahfp5KzoAEN1dUQQigoI9sAzNrPuZhe0Eod/NRfexo++IBLVSGetUN05jLQiZ
XLfnmwibVvYl0CVwAy4HXg6CW0Xi6PLKyxeZGVhUgKz8N0by6kPhJY8HSRlxDaKieSmUbR2vhS2N
tu2Z4AY14/9LZWFAgAwCcPEdhoTo+Dftm3zKh3VCl3EufgSoeonEdW9yefVm4NnEA07WDO6Qtkl9
GB4TGJ1dWA5JQxO2XJZOh9OtJbFlTBCwdbSpiqYl3YKu5S8Qr7w559N3LWfQkDQP5ff+BTzMzabB
bbcVO51kAA+hs3NnREUQBrLiZUjWEK6GxKL5H1yVeQRMtsNL0lSqTIcRsrQaADE8wZf9QFYTfbQV
9q/JUqu9CjcIe0jr/AnVZhFqpAYhusIUd3PJF5siduxCeRREnFzn4F2hxAIb1iF7pcMSV3VSKS0k
dDZQqdx1Ub4gm4nMa28Hqi9dDGALCPfvXy+t8n70AdyJWtH1+IROphKOJy4R5e6vm39ano+drvuH
v+M+sI9y5Movk3za3/Wx6Ljzn5hVizB8NQw4uqHSWlUP+mPjKhBt1vj5ooFeGIqqv9b9WjH0rbMf
DtAI+LNyVKJu/kyKW0Br6GKTIybg7TrM9Sfuvnf/+DZNei6kq1vW9U7w+iuQMwus0wBpXBvIi8RU
7wXtjUQtN/x9jAgi7PaNcKrdxaivrQQs1LBxgQAi/1128sowf2XVfD2sB1TtugCKsyu98wL4l1K6
K9yccsvWOGfgWC41KdBlW4MIfcxha1suW7kPhVJb3Nuov0cy29M3QBggFcCvcbq8f5PYBCq/3p/V
qUAxIOxl3mEpa1eD8xXEulnp9WNfvUtBMuNvt8LxFi43R6fnRcWedcxcJOWcQNSKL8lYaLFZ1e7Z
9iFI2hz/adCtougkrSqZoL6FJmtvPzSK6IZZMBGhbbY2QOZgFq6jtvuddpJ46yTNSQ5EV8Yvv9ba
4BE0azkvVBt6dsaf7C3ttKPnBwFN5LjLzSpA8swNFgJTSkuw73FAelXYFrrMUHNJ5J3NmK/VL7Wj
duJjz8wJ232DMnMZ/zdoQFtCKDtT6Ndqql0JMVJgtPbFP/hTIfVWSgJf1OQCTzS83p6yeGelqx7R
IYT3hx8kXPYF5GJs16LWEoKmzOg1UsMrCVYUno4IAqxfgjrF4O168MjKIKa+giZzM/uoboTDjQX4
fAZAqWnUcS3UduhdKt1ZjHXo6zr6578vVe5MrpqBPgdqSApbV94IIpKPoye7FOGu6z3yXkesUER9
xCEM1hp9EXa/1a/8NCDol6bRdtKVI1U+DnU0IQ3wmq/wt9UN/JJyIRHGObUbASam2KQC3dHn+/r2
oSRl0NbJy9/NdfUsa6ZfGMoeebkUndMdpvfRgtrPmSUB9ovVzulOGBWQWx6NZsuSVWkWJvIXFlHz
3LqN0Ktq+PNwuaGxCPsatylAdCiiLJdTUO4JZU3a9/z/cyrRhxRyDzHr/D96fkxr0Pfhroo+gonS
/qw1bt9FzhSp+VLMJhOuRslmW4V4oWW/yY379WzPt0aA6Qr/6AgtLToccy0EV2Al8gLjvnLxHhmQ
RI6h4HJffJDrQAH7TEevRGUIddAtbb39vRFLRaTm1TdzOxWMpmJPPpiBoOWnXzSGRI3cL5eQRz3Z
8ueIfWrv7IRkvRqpxMAIToWNZX5jo1oz3MG+JEZ7KOdJ6JIlmRJwKfMVZQfZP/6z33tHWZD91ZgG
0UDuBg9ImeQk7+LQHi2p3HMTR3TsniBQt2fes9f+QlIjE1Tq9y4QJsigxPRqSHA+G7z0Y5uoYn19
gneOqGwQw6kjzZwyi/LIJD4uYv7g3ReeNZpt5k/h2a+WTkiLtPj1w3CdgK1gbR65GRGUxRN+N1vM
TqkhLPbb1tZkbHuLTnClSgLZ0Rl+NEl0/A0Y2ZipvSVgT48Sn9dGZU4OYCE6ZKtVa5WzRLDuy/FH
/YkW8lTcvk1Vugsb/7XS8R2LWwchKZNoD/1i9L2xMtz4Y8GeZHbNU84GdjJG3iVm/nZ75K0FDzob
0kF1By/c1y/MujaFjJBaxxjLl0mgt1ulfKYc7Qfrj6B70/UjQ7lsyvPLXz3Jq5FkkF6aQYMiAkh4
APZiJ78oM8lmZZEampKZ1oo8O4RsVAPpoanj2jyLgYvGpL6CNsj04XbphBRyn8XavXHKSWRmMTqZ
UtAv7R8WfcB97cjoKMU2Z2aS9X36jL7JlGOoRS0xr7RtYEX/H+pHuAaUJCXL6P/b8iEjvDzysA/2
FwlIkxr5cuyCld4aYIGyTaHged0b5Dtf/eKRdGKvcbeAqHA/OsKLmkzpEqi8LOyKWCaQ5JOxOUJC
Yf9D/Vj8b8DokO2U+5c+fvpEMBxRLmeAdRLLTIAcjRjAf0RDMxeqrayAHI45rRmnvSw3TClpMmrG
lJCGlOiMS7QkvCnfSUhtWTh+hktU7yMOK9UxDWUhjcBytr5MbNVBQfF+1cnNnqpe03P8d6IJw1Gq
dgsGDbxj6UpGqPbNyJo8b1wsqLtSwE/9Fe2eHMz6QPBK1uoC3GUISdshC2mEGso1EAjj582b4Lxg
SDt6wU5vx05AoaPaBHOB0hbZ1Kv32tQY6grCRznCwaorsnc0s8zdL9yKP7mS3FbGpMZrcy7kho+Q
L3sF1/I+9g8trL5Vy4q+efhEuozmfuKQzgpr+oqRVI4D3sN0oNWdv/bLHncdtCF6dfPyFQ53g3tL
hRAMcgR+BjIk9KOR9jzv6uI1AzZO8eFPIxn3pUzhptMuhyHvP60YDHB91toxIMBATYl4ik2nGqtU
tRnSEB9aFWfqp9J5aDn1qYZOsjsXFLcSt/MxcVeo6xdvUUBR0WkpG3l3EjereEqTi1NZWo+wTTE8
5qPHQR7jkgvvO7IKOaLFa0aiojCQ597c/trVSVC06JA7KPyk4Rbw1Pa6/+3mch2J5iiyrpAVBA4b
ZU3qORm7x+6GzsIIsJEUBUmAdcgpbSTjmw2dXWdhyIThhjhOCRkvbYKp6ox1va2B40Uaw2EFAgUL
+r62Q+Pf59XZIS3ETo+3wLBPdVzJN/zFfoUsiBxKc0ObCRTrV10tf7N/AjUmh6Oi/9yugiBqjxvF
oZP0EgoT6GkTj9TM8+TSoBLsLgu57h7l3ORfC44nFCC3xqsC5cPEKWFyiVHoNTT9VtrCdd+Qzqmq
hD/4TnIAICD73dcB04EiIax9EIbK43XkCaVZ7vAGHhNdepnGRMWavGJ1ZwY1o3jmuUQ+HqOGsMS4
wjYkZfVsaOshXAerghBWizx1S9VBDc6FU5d94LJebdVAqQfMBMfoFpakkS2tM/YnW+qFHR7W/D90
ppYQrHgw6wowRSWf7j+hoY8rKlZDtNXqu9H06iIrBsBQJzP9ZpGb9tzvrPHGA8W/Nc8utz6LKr4+
RKBZjrXe8MRhjMuSRcZRIthF/rINFCdWpq9qZ3Dim+ZrGDLmcj3YDhf2qFS74hbmf7fV3Lf8rgev
fqvWjllccKDFLAZG+eIE8uyhUfPKW+xY/Y00hhzrQ7EtMMUOj2YKl9g9NJdAa8rYnKWXEzLHPfHQ
rwupv0fUx/CoIpifPECKvKJVWjaguyWWXayIg8SlBUUMgz2sCO3dKajqfI8VJYcjvPGX9zaHUOGm
WnlJdTlt2UymlovwK53p1TIcOReDEYySFDbldkgWwK+mqJh+vSH0z9+sFzVM/mOCpXG2u3++8eIQ
Qpy2qELhxxsP8nlqy5mUcAC7gNfOfxqFv0GyIiWpKPcOhW3N6DTe9QmV+HPVdn/Z3hMhyXaT0V0M
Cck/47vdcM59eiG5kQukVCApoXsOV80dTdfwqpqejVWa87kHDrHt2G2dPrRy8xa+55/qdMEYRTbg
ouGBcBSKzYHtDiQHEsfERD2ljDnryS526FdWvzWEDy5cGDh3Qhu+jwDZqZpOGK57ZBqvEWsPm+Sf
W5PZtDJpXaBmncfXi7cbLScWt/EpuI0POZhngm5tD0xe+F81JNI09n86u5v2BObPUr0n5MjPEbKh
EQGjySn2A5X3ojnx8k3SiBwUt7ctGJS/CM8/M2FlldTHAUeYZLGvHC+l+m//CeL2zus/maOjBPqs
Orv5rcFqlAyL600TqJau0VpmJFTQW9OTch6Ge+Fg3gMsuuXc4UTmMJ0XQEc66w09Pn4iVPyM7MCQ
WimfIlDzBtjxQ04Ql/Henrz7Z1Aioa3ufIAbTuxpL9PdJ61ar1FBHQkSgljusJJgulkJUNnPdTQe
qBwPXa6LvSII5RGwoX9L7mvmHTKB7K8xF1si6RzexOAncVS+R3ru23NrYUd1JsL27an6k0/f75V+
/XgPTQGtanICm5yRP2wzQGIEZFfZBEZmenj6cVDMVw2J6x/GYvSpelQGAN9SwMeomSufw6/qwcNF
dHQ62QzuZ/q+VSKLkfYb8aIr50MeH/CefAuXBgRngwBtpS3qlFJzkVp59g1FjKI2FQJ2Xg1Z6AI8
qectNeI4zQaOiMuVBVbDo/3Oic4OZCTpBsGC8qojn19XFzLFMMgMRx3V5t9w1Vzf0y6Z7eO4VB3o
ug1Y1qxoK39u0WD0EPJNDvM1RHtLFBnWJf9sZU4lei3NgcTRy0eRCEDN8jPu/1f7C0RqaLdyG02E
9zJ1rLzCjB7vq9vBkQhfgAj19eIQoO9UmeKwKwk0c1p3NnfrjXmGAJWTicVLDCwJcEapz+vjdWir
2Kfg4ZSybPfg3mpflfESHzBJwyuh6h1X1WCs60w5qsH3f7WM+/TfLOFi893kNQXvLNNiRccWTad4
UrjAWx7nM+TV/6IzPB3qzkMC/h4jTT2SkaoZsl1UcOQ3khJ5jPKKVNyMU2iR+dL76RuS4CdSATpP
XgdGvM8Ktt2eduYLQoGUY3Z1IOWXbCkHaH1fOnIkVlnrCYs6Z1pPciAapoW7ob6JebKyoVvVefgp
9b3+a+UVVKPeo7qzW6Myd9VbU2FfjtTmi23V8/30eckV3jMYwxyinEJCEOP5XzEtyTJkCMij90tZ
nsgiB5QvMZ5/Z6/C/hv0Ormb93LXhdD69E0MaUVd2Y1ZJNjuEgrt5p58rY5/JNkg2/9Penmgrw+Z
szVl7ddGCdnheVHgqvqjCGETTodNieB+6fJSpS/GgxVDphkJm/lsgSuzbL8SS1Ikwwnwj7Efk6g/
KTASQnZhUvCYVYMn9KIY7shnqtOYFFBAlrKyMYh4uMHc2atw8SvnFP9n1qhPbpCQwSg/eD/VJWaL
KirM593DOoplvS8laEsRlFDWqTBLrW+AVY+IzwoNOEzp9IG6aLu3Ci//HZkdiyc4EUeM4W7FTqEV
jvOpwVYXuKPYIEf/5KS6yfx8Xw75hGB6CQxvuXYrweVYiBSHfhhuxTKVEJLwcd1q3Gf++kD4PUz1
nBmGc5F6gRwdolXWMZwFnAEfYZtY7TQD3D0SGX+x0I6zpETMz1wbOy0y7kWGL5XWXBWxud8y9WsA
f6JZeIUgJ2+mJSG7KcPGdvntycrzThR5EgkahUmt3YO+AUVnONpUU4TTOEhHP4RMI2RgHRVgxIHc
1cW32JYMfv26Gq0w8yVZ16EVTeVQOdSsn/qKKxLPgYIPH0Kk8J44DsI8QsCZQukoTXLG5se11sts
A/KQeqKRF+3+Z6NF9kvSHe6WtKZsn5m37JiZUBbWM4XXiR7xXNeDtnz24JIlMzOaZ3JvVTCWewSo
LtWNadQRnQOx7pWh7hin2LSIjhHsNrlVigHLiqdtDe9R8PFcRJQZM3yNSu6vuhoIcz9+DoHC8R8x
2UomK9eg6UAXrfbwCG/Ubj6WRc4SJcsemUkscIPRU/2XAJEBPNglK53ikrWixNd6+UUz8AukvuLQ
2bJ+HiaPgxwnJghyRq12Xy9fjRGN+SVXw42jwWdbBHZDdurKByLetT1FSvETBnyWWYl85cPYza6I
eDqUZloAa3BS6NqEPrXU3MlSmkzZUAczd5NR926debDH7zURBe/L69xK5vLBgaFi7utQcRCxFfgl
BJ0QQNXPB6QxIWmYCCSqe3VqCLV/jUldeaIGixLCVp5b9r6yAPiUfUIPoDEjgcpBlHH9juRRhQRy
xe5Yjg22X9Nz36EqHb2tDwzw3omON+x7Y856Qx51V2CZ0tis+Li62PV1k3mdqjmAcgW5iU+3EdtK
tuoPROfhb9Gne+/8NeXNndslxBhpOcYZgiNKXODEHcu0VvgrlkjurG04+RJWVFImKq4rUeYT+NrD
RUi9IyE+hu//zaQ+Bz9Vyk1LNY4tCkINOD3G0aT7j6PZHHL/DX+erb2JpiSYbPY7GCj9zgjgMTuk
LejrUs5rW3XChRuXhWCiwLtjklzHTSYuo0LRTIur0kBzdTwL3Ufs4Wfxi+TGZLy1i8855xACwHI7
hhA9q/WDu0iwwxU3jQuJx0rkGG/UMHov7URDD8Sc4axOujGoRCsmw4VwahkhPy7cbVrP18iGAVsT
rhiO8HYPKBb08xTI8Kg+epwdpOkv8mKBkBayjUlLNwb7gDVSeXgzPWcxcrVws+dcEcZKLNosmIhD
v3y1S9YzNcsab7Mw1klPcBiGcaQzhJzDvMvcjqPTnFIveJ2tvOV95ux8TjhqMcm8mvGN6Q4g7f6/
HtPsvAQ2jY4Zi4dx2bF4R2qqMN8tinzI+RDqMSPf3N2IYV+cO68y9w+0/2pFp1O8LlH+WZ/q7kdi
ZnAbRRN2sILs8xzVVit4LBwPj5yzNrxlCC9V63cFlqOBJfWA/RV5rarIJrbzVphdHbgX+j1Duf8A
AiU3u6xyEfPOjF00s/QyInHd8VT2RP8SY2rVcKMd/Aw6tWGBF/5BFq/9c7zhhQIYgk2BC9OaT8/G
+xEuMi/q3PqnYfRsShpdVhkpnpfVbe2hwnw2YZVcdFi0eDYzf9c26mBvgURpmnAP9oM8ElED+cOL
ZxnEtKdKIBC+RvWTFMnKVPx5bessreUxJHqiz0c+ojjRr/nhg3mzQ0j0zV8W24SM7LDG+CejH488
O1Pq/DNmHvJNkbSoetk5KvQi0LMCp9yCpa3u5CGZtVKxICaQroiHgAfUcYNY+Gv2ILFEgQ28uwOn
Opjy057Nbv6xdw8RKmgE23fhS2OrBqMmCa8UKT10YWfSIlaW7xbdkjKMfMhgG0NgbHr21US84haH
jdIR7FCEYTOsdKrgwA4AJ935xy2ujy1gWbciMJQvF1sYBtnl7VWh+WWZqzAGqqliVr0gzL/3za0q
2DEnCCr0+8NPgJpvjXkoYP/InhW2zmU1GdhlB4DRPZNslAcbdiPLrDzW7cDPZucNoaCVUNsUHQo7
Yp1lMHHWT3zmrBzQEok5TCkuGWtfvOOxN18Uzcz1t8Mx7OHZgUCpMnG8HzinF33YEYWvtrh273e2
c/kFtw+IHs157wxBdfFcv1zKcc8xVzSjKm0fWIQy7Qvbo2bgLFq5BIUTAFAZDg89lr20zBHpahJq
mNBT543z1MZpEygcJpCM9bA6gd1j7H5JM87nn8CpAac4UX2j5EvLNXX8kFgK+zjxQi8FnaPl2qEu
vzzGI26Y/OTncs/fZloJfj2oB9DmHiPI8yJyrivEeC3U1dhFZBuVTAXX0gjrrDGpAOXE85lvZsdF
E3BLu9qz0A0Tim2sh5n4jGKXfSv/hRT5nPPVSPRqqYujhAmnWyXwuSsv4gTT6dNPKtNb1fem7z0n
AmCom9Bei4BMmOsnnbK2cx4FM+aRSKaz1WM2QCoG6h0tHW/pxOA6SvpNXBXZV1WCYIUycTHHxej7
s77fCj3b1wR/S49bFOYRjX5w1IBAl4WPHI0DVx7nry78ZNWy7/hp8OsUAuklJoXt/W7kYJNMLmpH
yxrmdLQ3ExPctf7b9ncXM2iZsVcojsPAvsjyNmm/XeXKEku5q3TXi8Fdpr8xKNzM6SgTI0ZIij2R
m5LbwgFxzvSuX8LtcrROdy4sfSMvN5PktDtGrooshH9R3s/+jmGxYxH+45r/T2315CN+ecnz5Bfv
1HBz5MBWmaMHXkEzvexPZNk/Jj9xZP4JP9hbu8AoBtpN15NBXe4IUxk9EmGH0wiVfYiZVLu0e7wD
0hHyX65bKCqeKvYtQlEwcx6CqWD8GkQvB3I2OmzATRcgm85gf+U2IhdZMZbqdnkmqk1eoUn+W367
eHvfX8vtTFVQTVGohTTqg1nO84SWI+PMa/3T/okxVIfwqSANo4/mBdWCjIHplZfuvywrtnNfilJt
8EAzVVwJY2rwdyE+S8B3R+MrU6C5gNDWEtOoAwCM8+0gZNAv4V2PTC/LYR3q8v98TNWUVWqIP04o
sz7kw6OnoN3HpyyF648nfT1m96basiVilyI/K+Qv0Gv9GbDRuDB0OapFhfGY7pPQGN4Oc8DCwDvp
ABowFyrCbN92zzcNS0clmDxLUKFvP6s6OEiPVkVM9Ca1GScqjw4zHSZXxQ2E66IWknkPDKpDkwfU
JAqPyQBKoSaCYPO6c6VNM+kVAqHtM1tvGbgvRCD5cVrVK0J5Wf4OAvY7oCsy+nzYpIeAuSItIxE2
827BtEt7kr3osiDb5q8Vb2oFJhpw6U+AyrmMYwDXUDX6kbT2TAsLyR1LUuOCzWUPz2ATr4t/1kuc
iCWhHbOTkL1vueJR4+aMPIA5Cfj8uKY2ChUp7ra9l8ujJ/Ym9j+hW57vceya9U75ljj+Pd/pVyvJ
+TjOC3aq9nc2WeAjeUDOyz3QFSJCnUqs7mI7XSBz2a+IcRksAcSg5htzlNdIwBU9M9RszdguRLBy
1tZT7pJTfQj/YX0bSA81NbEiZO1ZkGb0xgkIh3pTa1hNCev3gk+PYarJin6Hg7yhumJCf+w1M9h0
XHvuH2zh4HB7o1IumgJze8rz1F9rTbPF7oN365jIeNpom2EDfUzAe7G9Kos4bUIipE4l65sUNv9D
X9ZUVhwoITF1J+gD5i+qWMHFqk2q49ylbHgR76koVLnKstE1WQJXqDnwdkmcihxazqrA1PRbzoWq
0TOjL6gK4L5LQi636kUZNq9BoZnucPllG9GSh9yqu+uUFE+xUg80zFLarP/088ITo4mSTH09Whfr
lWVnL/279xxMresKQ9NSItpI7w2tO+nDUmB4VXo5tEeErXcyFDGZvMT482iYaMfpAOKGdYKeq2uL
c6V1aYvyj84gamiCLj0K4mB56lq1/j5wNJgTa1s4blPoi1V3h3e3JGqz+AH9Iintb3m0EqmB9h+V
dvZQQLWLmzsMEKl0fdCej2tRfMvOQ+wdtZ6qF6RiUJewVoBrLClf/szKYtSdOMDddZfJTVIulgTY
dGdBv9zOhj7ciCsNkiQIg2WVYm1uq79nlNI8na08n1crkS0PQv3iFa57Bl8os4p1mJpQHjrkW8gI
aKL/amoxq4UV6JDxztJellzFZ3d3snJ1DfX0Vp5fkZZVRNfcVF/Kkve94IOPDgjb5bu7qVyAZPJ7
hgm4auCCdgHSAsJIqfi3dbsXTj4Ipn4wVdhzZKXwKmActBWhJ/rVbo2X+zf375SWp7iQRuuYP25w
ZTG4WGphFpYK/r186vy7l1xBCRCKaXm4Jmg1zJs4NDbCJubFdIa5o1HDhAQIE+Qo3PUgg4VJFYj1
WOLbxnWrJ8jWVYm3ARyj6WfTdlpWvqqX8nv8oMae7mt8L6ROnTsEobRCOcCykipmHsELQY9i9SXs
atWu4oGTq9XjrCU+LrM2eY/cIwFzGIBGciAfECRmYBdwB6ARJYRORt7iZbMNXBRfwjv/mQBhApvH
kLN+Hb0d4s9sQFc9v7ToUdFJJM2fpvwb9katrTnjd2AB0cvySkZ1Zjhih/bc1MjH6ZS1MKtzQhWZ
onqoHK0IuMKeiwXgqt3AuLWsJuCgIYeW38eqYfQK6Jp7wp2i2NH8//EWus7aC7S1nfiHPOTk+dcc
T7lZXN/AY/zRzw57zwj1xblgr2Lya63ClKp14TAPPJcLWMlGJe7PIKdnZ7b0S1cy0QFZJ5KbgkO9
DxnLCLzDK0OzIjnnVjaPY3BJmqVzKpUyHxYZVKgEaOgIZSV6xWgsbzGAHlLlz9N8pgt1wqN2+0ou
iUkwnLWbHGb6ZWnQ0yB8t3DOIiLxvuqTU54tCU8SUQT377uwoekeqFVCGNxxiRtvAnUVJwKeUHuD
gYBUnn1oPvKDVGCyRQjBbY/WaY4S92/9vwWw+JgJTW1IjoUnhA3D7y5BYgm1CTBOSsmAmLHZCxgW
OasW6Z0Q6Y1nWpOoxe3WOw6QExSyu2VaI9v5X5IJx7jMXAQYZ2hNj7FdiiAPjvYzQCrK5EWkZhdA
OBg/eJmWubYgFjrf2gAsR2LuB1VkNo0jNBtfCUkRqogb3Ncgk6CqXDVTUPD+ssWx9fcDb2y9T2zI
6qM1vd5wcpBoYpuyJv2qpuz8NK6HSL9+sAXRkTCeQWdQkqtdoiXMJ8FYYZ2aUQ3dYCz0kcNdcyZe
azrq4BhavHicNzNby/YrZVuJnYVi8T34TaCHTXst+CyFuuy0q8w5u7FDpZsBIejCnswYOSI1gV7F
7weA/CJtvn7zX5kh43txdc8g/G+Uv2WPWCktvbZK9qfdtyX+8Dj41wN4z40wUBx7BA9t+feUy9n6
l6zSb1W9fZuILozfcllO4ypx14VpM8uNKL+1nA93iTEUJxONfkXAPqmKb+4DsDU2Ufgyu9N+hGvi
ibjwCJopyTRSdh1HyL5pJ3V7U+PqvMU9yDM4TFFAvhOlgLabHrL+k+g2zBfcCN95h8KlyZcMdWWG
n1zMLpUu4+JnJETFTiSsFxoueRN0ZjRTzKyKZMEVrAuIZr+9JkqDyd8nfdUKwEGghC2058UyT8ay
7REykO0D+vpagyrTIcpDDS6HTzYS3GWMG9YeV/g4AzSkcuhHjsJ5XgIL5VohZJOm4622JzQUj90F
nLSGloq2iJMWSD+/0myeKyBoXkCU1O/O9lStSnoTtwQumKYqFe8JSmTETPqbHCPiQh2f6maDN9oX
xVJ9Bqr2WxPwes1eAa46CJ/YGMRuocRco5bqeesfhy4yhlQ/o91jY8mZqm1GrnOEudF0QpajX8Cz
QHyaYJsopbAI44gHX6sfs4CnkE/8yoLiHC5tPMbcgQJe/jDRlRY7ehlavCERyuEIYKjYtUzOkaZB
CQbJLr40J0/99WBaAWnarQ5IH4igF1lCHMzUJO/ck4XIzdgqh0i1x6eM2h2j1Luo9g/15rXUZWDw
gwe0p4tBh6focQesZv/mIrhTAIIo1XaBLkMC91PBpsk1281GLp1obP7QuvnhwVB2tMgQbaTySp89
eD/CYvzKoBvdmu9nzpFQgjNlwJ4ANIHYIhbDd7i+V4CAXOlBk8TT7ufOo9IQZotX/PZvnernQvuN
wRKcOBwqmrlgS6dwJ6vtIUhroagJkcmtoh+2V4Db4fsZEkTLSdszo1WPI8xlsmA7KbWeLXLrTz6V
SqdhXCwHOo7m8sGfxxDtZI6fn3a2WNmhti6iAQT5J7T5LBihQv36CqT1M1keb59gIXa1bHeOMIq8
vMheferq42E1PdmF+KWn6mPlAnd9ml0VHAOv2TGu+YrJkNJejupiE8uk716+veKa4vYEUVc8FU3v
/s9HZlDUkoJUhyA14SBORmuoePRr3W28FUSH/uhcw31Ea7nisYCABG2JW1hsTAanZzddP94oReli
C8UogNPcTR+5NSEhuwM/j+zUb+Aa6j4/eLb0+o60Vrvbg1Ap3AQFMsGrvktTpIrOZNcCydlbrxQf
VKfNAYrPWfhGVEt9j24Q/nNoOfmALMIBMO79RUcS99U8ZbIyp46S+NKiTqFka5RNWK9SS1q9t/UU
1Tr0ZSav9JUpXuXcmI1GsWG4J7IMyRNLlbZZRTGQPVezBXO2QeSbIXAQpEXrxiplh2wvu9ja/EeY
hOIik8uAMiV8v/KEo1IqtkIK/4eXCG7vs+X6S40T9cg+YwaB3maDE6VdBT2xT669p3U5K+jZMRrz
ps4avuHO9Fd9DGWvWiwQy/MLuwCeYVEOyVE/ylJEvO/K1G316FUJFbXwNXkG2WZsJ4dlEFh2FbiD
B64i095PfBVYuu7z+mTpMNwy8ETT9YnXRF8X4nKAYLb+ER0BHMKBAulXEB0lnxiKAuj/LXSZ/CDn
BRzWdwtaBkhWSji3USTGS2LkGF5Huuub0tkTWd5bp6NV6HPmBTozCI/QvTjTuPixqhpMCn82Gwlj
XuTi0BuhaAUhvYj+ntURKW87d2UL7SZ/ZC4yVea9e8HlpPVgmfoINndZgCquWnsTrCh9opsBWRGO
/LTbV8aDOlEZpop56ILAkQahVh5q1cjEo3i3dgjTwJ9aRT4lBVnw2StiiHiQI63P3iXlypkg6jVJ
XxESSoa8/QMg1Hf37qyU2RAdPSKXee46h4HJpaatKgBuLUn/prxwbpDeua7AJzc9IXwBXuy3TfX1
y4ZVCRlSCNqtqzdn135PptCDah7UF9WmBSEwN5KdnFL5NsmFihtfKaolQoZdBj2ZGkJyLOegvNqy
QsRhoUcQz34AMnl7gEzMHzKcccUe5c6uD6g6kfJJq94qPh1I89JxuaW3Rlg4G42aU0TJLrFyfD90
WmVWFlp5qr25U1kAsda/1r9+s5NcCbHSXDH299/9LScbx17QHp+Jru9B2RXXui67PeXuWaluBl4k
6n7Qo/xbbTWK7wFKcC07SwTmcY0eUIRG9Fs6TV1tfmEzC9NbxddnVS8c2T7q6175v6AlKX/LJZk5
Qr6c4BKzV8nMYkG+wWtrbf60bmS1RpRvcIIl8jmcphtQgTfehK3ce8oe5/cUjeigCVq0OVePw92I
xTUHNLJaZHGrfsAOyktfL+0mC6PkYxMhNWpGOceRnM8mFxSx1edx0BATLZH1snvpz1INwbQHbjwA
Q1+YCj67qxBxq/wqlvlHNTp2021cZbBivA/MivkYP+n/VB5Ifosmcv0Xtt1gQLM2lyGoVximjdPl
cJ5P5Zm2EXF3qJU04AOeCTpbPXtu0LsCUVwZ/uLeD5InCqlbdhs7YxwGzWsUYNyu3+pMXuzFNKku
mIJ17jGzEOWPiUjNeVEUbKz684jMfQrL2m+D0xcwVrlhpMkDcwTXTRoZNtIZLLh6t3L7xKWxSB56
D+RhVUu7lBgcT1Q+L1WC8tlCdOJFay7Ky2duMiLL3GrOcqKdxynUydkVcNosfhioR3UgtZR5KMA9
7tNf+e18LIxgrqfviVngSLEZkmtiH2oryweJW98M3u/+2lfGFbqrkzDRUJqVH1C7pi1Uf4vhVFRk
gwHEwlFIMmClsAS65n9roxSM2WKAqqADudy99vgkV3yfJaKRpGaVtEk1NGjAQPH/D5iLtKcZNlej
3nUmybAM1+Jp8gLSIxL2B0UP/Q0ICDsF7wEL2tsH52FVuIK8dKU98Y+KM8B3MumIi9oYRx1OP+Fr
7kE93Fm0BGt8AWHWkHaZmitnsSV9Z21EeyPRw2ggfx5UDocDV8d6wpkLBnXevRDvDutX976lwowz
xRRfoTRQSpw+73dm+HyZC81jjy012cvv20GmeaNqqPhX1Q2nT1RU+btb3XiWwHlR8oLELZd0JfrG
nujYwuXmHinvO27xoEHYhY6yh31XnxGkKJLi5IxufBNIBjH/Ud1CgpSo9PJCljIABGKRCBVcBFbn
ef2cjW39GUN8QoMEGI77W3eIG7iB2PKrRkMg4I+jdMDL0LprpXq3lSUYuJ2irvYjhcQ67Y2QTWr1
LV5AdJMbRta6lwU/zeLfsQSokhn8JaDJ9CF3sPl/Gs1rItuSQhbmmHUN9CbBL86OPKvBjBnGqfCx
caZoW1D4LfGLmJpI8gwq0artK/+e0lbGZ64X6FUnHKgtnw0EQu2r3cbhAzwcplshurDnWCTob3up
ZV3DSbWkDrdGOfXxi3byWdZINQ+hS8Cn+PG2M2fQPd1n3j8phD5lWmr4EoLjqKwIte+5w1ANdlOi
RKIHV0wIB5RXtC72Jg6CLZMxZVBBPRRx1MKcYQPJMlnwxSR6OGZjtZ/1nuhvTr3Lu0twmwIOnXP7
ZyMhM5/zUlQ3OxvsM8zBuT2R0m0GYDLciAaZYbfn03XfE14+iIFhlpwNh/Oq+XDFdApqhTuWvLck
m9qvG3d5qbVtwzJq0q+L5eGG+2ii7OpNht9aRHMvZgnchI090ErVQIBNKwZzaE3YgLPA6zBd6nHy
o8ZBmjkg+OaDeDBZN/pBqjQKpW6U5vn2CHcsYSGYweeXeTu2sxOP+lPcZHHU/woHvXhPiU9axNuf
TFfGFcYRPyW9WA0foXbWOJenUUb/Sr2cTwiZVRzBsam2WWOAu37lkZPz32jjzFXTuVssGm3GlChs
pXG9EhfQDS4+DZD1WjYK8efiQVeA6T9Dj9wRMy/okphi6QWawWsxs5cv3nm2lhIspzyKX+xqozST
BLY8erqrpaTc7K0eUGIcbfCL6y+/g24iHqf1RWW0wXyMNADwUHJAX+mBTNG4IzJ2TbsU+DPsT/Jh
XGgnDX5yilwKulhgZC+iV+4CwXqTHq6mdcY/sUAcktSe85+EaYV52w9wQHU9zaMAaIiGO8FpDwCU
GMaCJqwT+Uqf2ZsXh1GdG8LUxztCMWWCTS1BkfcenBKG8x8TsduWmQpEQIAGBUZ+ygfFNtkR991g
VNniRlhC8khUTu23n8xyINtAbkOUUOz2L2lIBiPlwJKVL8h1LA4ehO8PpeJ5edIIgle9uoF+dfgk
RhwBNTBlXregq3Myx5yWibJ2GnqMD216BNGei8LDHg3xBqticEocPndDlECZil/dET/oFaFeFIq3
YcpiKINtRNEaFIEcNNuFcqTmp/HbKtQWkEIyxFGPqO0VxREEaOFbz4bw/m0f1dcgIRktj1ZPHoct
/Qp+/SC+PJNG6xamQsf0/pNZMupVsWgHYidRHGnLouD5UpCQZD1cdyYCSv2cMQgiOvpmjudMwSRb
nZoFNhQU8LfLMW5EUfr143YnMvwFGHjCgMkzt/a/qTBC86cZesgrH0CGAArKxO62GtucHtp3vn+Y
eigsPu6M5w8XQy0ESEP+LSPQ8udqmxkfcZ9PEreNzDpKowOdplQkOh0Fpj62ehSofUYyR90SiIQZ
QRY3qbGjh6JWHv84MKVkx7GeWuDat2nqmzcyTiiIFFloEXumoZ1YuIfXOGdzgFlg0Hn02xZHCIaD
WILmco3m0xHarlII+1TD+z1e/UE8GqaIQuBT0tTERpjkRGyd8DucnKwsHCu+z01DXONBU/EyGBDf
KdLA6emvYT+ZlCFw2c9D7uiLeLcquJoLkZ8EpkyC8ltUJL1M2YxlEajEdqQNEmXCjRYp6istsiT+
D1RimoVNUMOmfvfbMJJb6sZQLduGNTAW7tuWI9IOMI96suFpkxySRJnDE3Oy9tdIcRFETehe5W9w
L2mouM0MvHJ8s/vVEB37X6Y8R+b4SGadQqBZhXbS8Uk6VxUokaAJLjOcf6JaFm8rJU583ZjQZ+0Q
baa9iWwuESzCVLFo0mng23/reDg4akeuIarap+VhwzQDrDth72Pka6y+jo/pSi4qUkX4XC/tfbhj
I0R0vMjsGv4AUtLz+CNBu3sq0DcMCaR4d3ZHvMioVBT9akyW3N4+Ll8QKRayMZjA7aezyIsDO531
w1hogkpiG6GE/qRW3r4Tlqcb9VcTd8MMNP9ddisagFbwkLIhG3a2hQ5oB9Pts7pFYTt9tF4HWcXb
wzkFo9EmECq5j+Wrl3CQ7pgWp/VYmtsdeVvv4tpWOyVuKCSbj18nDFfIRqqZSD9nLCPTbZgfy+Tn
kxYa9vYLMPXlpujFrGpcBvSV/bBCqOzat+F7eyGNFLyeJDysdijkhgDxU5LfhAfBMxuD1HXnmdfG
/+TwrZXz9VmaVtzfzD/rAx/3L2mHn37BMQ6ThOUoFfiXzOIkfsuA0E7n6ILRwmxiqh1V7q9vtOyS
e+lSmSiRwaPtgVWm6k3/jc/jfMkXVF1itCm+KM2g0b1uePGHIzDJTIc7xVV1nW5ids+mIWHuKLcB
lSaUmjQ0Lt4vzm8YEOWOWQPnEahrhtzPMHEw3UDOMTgas5FcRGdoexu/kKGRrYPYpRIihqHz9qpk
w1YOkRQrzS39OTxR6+Z+fdpa9Q9YQFqwWENDx2NEe618zOpzXpJ5gyJ7/lzrKMW7QXEG277STqvd
pd8g3OYQpokk/4az3ciEHhnOdRrXPHRm5DVcW9XX/szdZUMrmJ5rd61eHOuTs+GYBxZciVZ6MsUc
cJuIXoX+h/Rr9b2J/UuTEDcdGVO6+YgBYYdzl4b+HT/iwvP+trSSqG/wGtOvpCyAG1aCjla26B6t
7VmqaneWlfaXstpD0mLvGditbtvr9L2c+hYjYlf6WbAKmU3DIw3YZdR+dkLcKSoFPmOFE+s2BD8p
QhHVpm3P9QdhGwAEJEC5i3wa4So2V3BMZZajW/ULye3PMOMgBmYjhcOG6dLizOdUO7kMHsc6+uc/
LUtzNh7AlNPCkl+OelzJbakHTfY3s6PmA8T9CKSBnn5AY1LoYyDmIZDd8Jxh5XZXO6I80UuucKZZ
dhlgIeRF5vBgXnxy206gtH6A/vu01HCVqGybV8rOpaBIkGTaL9RZUrOx1Y4yOw3ZZKuCm3l+XDOy
YHWw3PUFO0k1deo3Zq5h7D/axIf0Lae45J9P6nWJyBvex7J39SqDVeTXB0VwJK2a2+1pQXvXw3Je
1MqKEuJdBRBOsop2tZG2hqwjPrlyuf1tAje9+07NHevUxnTZQYoJ0HRCzqFQp/s2PKuc93+Lu3Et
XR+yZBt3TP3QXvm7SxZ1pwiHHVZT6zTyoEYXt3K5U3Kz0lUdrKqIMmS1d8FJ5QHonYU1Ku/NO1q7
WXd4kC6GiJVOLG197iHimvOpBthk2tLhJcInwoe22SqfvW7TcQ/fS/Yms+QSLcjWfDhF3/3UI8jo
8nUfAYmZByNvb4nlCw7A4Fo2R48ez+Wqxxsr/hD94X52d18o0J7bscYnxihuNEKwLGorIgVgLsvW
9P+7DS0zO4wAaXNKxwzEdJ0Ehlhz7O5WwKDtBpcdR+vZXr5O7ykcWO07WDgAw7Ii5kqQapNYTIld
6dTIH20Mvl6LTuhju1KGyj845HNrFJI14BaKWLaHZJ4ayPXAhJYaUDtE+kHDekHM3aT7AIz/B+FM
4Fe5BFVdjFzBy4NcTFe8FnbFJoRhfra3rub7+njdq+32KOWKaGLE5oKsq0AoySjXpHjseXcokqIe
wHTCaPEf9izEH0oPV7lm2GjNhgTDcD3eyzN4VoH9ebAZf/hCsnPUqeTB/k5cv7oZModttmMvOvAK
ftSiN76+QkukjHUEZBSgwcE7/UUmmh/GqXfgqxlBJoo2NOifdAHesWZRvkD8rySLXmRV+DdJ09T5
H7icyJSX2YrkqY6tzMFkfcS0l/TC98pFAwLuxYkK0fw3viJOMWjuyrL77o/cakL+x+kYlHu7AwAH
FGzkteVp0eZTzXd+K751LprBK6udNoHmpAJ99pwR/O2cngPn/1w5VXyby8GP3WUVSb4nGfCGcyQR
OFFV7Bh8RLzNCP0O+EuKNwoULvXRI7Hxbc5SXF9ua8Yafz3DfghWK+0yAs5t6c27Z8EmKKrOwI2u
QE875PHvsaq6JxHG75LZVAX0KdpWCjTkmDb/ndg3kOlZYDREiqU5WeyfV+VeCVM+7iUdIrz/kGll
fRhuGMz8X7ZtlhOENSH9Z524blpiHbf83QtH4+pOBENoPsSARomqk9qMKdG5+arPGLzd700X+ULc
zBkHe4Dvn4qMip64PrZACgC2kIOHHhTsBf/4HD37vQxeRIYwUaxh3ENgjgcQLELYUKDjRwkaqxo/
4HQktWB8qSJQNEit6StNVuDBy3ffzCb4UqA6QLmjbRJ+pXMZf5yseniZylU+5Yil+YvkElAadjPb
3Oct/tUtWU98nrlWAKocKQnVPJFQRx0J+SIrMMYsigHgCL+F2A/kIffUvAmGDU55PZ9BOOgpm2aD
RtGBgl8wC520qdFtsikXxQasJzLArOzE+Zv7Cl3+VuUD+yrq1h6KJst9UfRSa52e/tps47PNa8z3
HJNbFIRNTDwBZj3x9dQ/UsmrErUI9B4O2/Dk+g255kTfShPQrNpYS9IHljh0X1u10F8dfODLLgQJ
kWOL2qP7BclkT0LU0YNF1KtMgNvmM7y/RPVDC1ABnohajmGAptsTpBrFUTuoCMkQUoZilz0e7Pb/
HVVz2tOileBvPLFdXVfdUWWYCCjtTdkAtg+m0lkhEUQSgn1k0uHVMQ7t3k5qDPceufy+3IMSKuUO
q8yYzg6zg44wUabGR1ygTYsYFT3/+EnZ2m7X+xFTo8LHKGydIp4FoZAV16beDgiInFRJsNcolQ0/
qBvAuf4sTlMvNCrheQxGgC/uJfH68F7hAMbZgY7UkRcyKhX2m3nfZB/2nEg9bRI/lA46H1WvX2Ce
TkQ2NyF1ehUXAZRvpNbL1gj49wjhxK4YfTWFqBer/7MtSk/YUK3UR8kD3w6+PoOB+vLSkjHJDt5L
IlL/fJAuhb+EPaP2J4mC8v+gbWg3xUAtb0rk3Wt53Jj9yy2ciCKlXuUSTgpbAz6JdaVfyTfeLFZa
x4Nns+1TD/OxYV3/MJl9PqCIq3HP0gVsKyvCHuSBmdqLS73RfaMLPxhyFyCNgdJ0wTtb7wxokUpg
9WGlgw85S0GiuQiSGp7MhjL8gtyvYXsCuKMzY2NKkuyIcGCT7n9Upt69Yqgfiw6miqNE+JQOrixb
uDnuS2g2VUVjDq/lnKKG3josTCYF7QC+iP73ddZ2rrQCnrGFWkE2dwTruhy/HsiN45pQ+321uBoQ
XKcHXH6UyXGHH0p+7JRzYyK3b8/jZDWI7lz+5P5JbCZ1xxAtqv1O2uhDXJ+FhqkixkUVyEMkJKIK
8Mu3HRYlBchRfwXGq5OEmtBSJA/oyw7KpeFUKzOWFiAWttx/XnAnX6ke7AmZUBfFlbl+T1+dIj8j
dYKOc/8CTdWOsfQX2yhVSmW6lmmtdwpKEXVH361oM8NR4TiAvTY+urF9f/j4Gm0ncJj1DdvY83Q2
xUSsFCqG4xIwbS5zHKQP1ss/ffrm2rlZ5nn+xkNqzDmFiVIaZNMEkTWrcphBmgHrMD9jWNOio7fB
srV9+6eAgckD3EM5xbMgX8KkqUi5xFghM2eJLqDTrGhwTlw67RaKnhz+2cRvjS4hVhYFDrAyuZ63
GFph9EFiCOZZoZ3j61fiTR3FKBc2HdAu1GVuuiu+mpRvBiEGaahzFO8RQtYetYqltb6hCorTfzNP
2hLrg1M8L17ovPER1IUyUvC7d4WGCLUgWIvb8i7YvLwLko5cQsYqaQ7v+Y4gA3hHLOjlDSW8Lrvj
PA+zv8cqOlibqpaHj3oRmb1GIRqs4Q5rdMkBLpvugurAut89Ip2zcY3gsQwdXeI8Y2MWkbRv21CE
Xt/yrPHqQZ8zGzhOwoOkqt4tiGjsRicF6VQm7SbzkdI4KZQriLr1T8/vbOvZX8yUTn+DQ+2ZEfRV
TVv1hwMwSW3HnBkyWDdiOUi3qQYOtBVMjq8Yt90O1UlQxIoxf4rbTjFy0TPbQ8v3hWgad2kBHKzp
rzPHf8TJEDR7/bPh0V6TFB5ocr5565gxXHuhdEk87hlePHiDZC+TOpVMqswjaMj/jwLpoEJFUeC+
ldmaOhRN5DFs7WlAjdha2wQx1n5xQD6LLQ55+L0ssIfJtn9pnbdHgCQ39sC6G0PAXmnR11IfYAHw
GI8sS0H5U1J8UHrPjLjnHS8Bi6ngzoDLfLfcw/AVXATOSM8/cuDcsv0WZR/Au+jRsbeN4owT8hlm
oKkmzpvpnvj2slsFP5nremWLXR50X+mumO+kqxhHsEf8XKbQGrd8aTcSiyN+rbaLR6YFQQC6lzUo
NZJovK+wIjhzrMl+hvj0cuIO5YGqOC1KJytzk6s7U56sH/r9wf/FuALk6xk6hijl6tits0cdpGw8
EZYrGaDZ58uotQhctRdav1KLg1PkbgB0Ps26OvUB0DbZQFtKU/qoo7rAkpxIpTzjWllhH6hEcafl
Z8jlyvFAY9MaXhnD4vlxdT8p0g/zcIe42aYJSozKxbyNwLXrJQMdc92IvxlFsUCBwOZHWljpFE60
jCbiPoy7wO2o1qSoSiL/7RE6cKHbej1VhcCkm1T364xndK5DVrt8LLMJmyWbAh1SUCiSH7V6sgEg
iGotxwU/heWX6R+iV1/KZ5nAV3KuczS9xkFC6y2I/1d52UYgTGEkHOCOTa0cIB8QxXwlAkUKENoG
DKLJuzsUHDEZtUYUy1NLW/cqtMf8Zn4ZxzB1tWSnb+tCXWT4Do9LCjREevT1cV64JrFBsABs2SNf
Vihr8xD37eUI8AWuQxkSGfWcjCY+p5ZHhXebvsg3BtYlCDrS7AUyO0HCKNPqCSfhvs+JE8t2kDe6
ozFHBCC8PchMtCa8tvALt7YJTFlDRLO92FcnyVaYgNCHBxCe4jun6CGcTFHiueNAsYUQe2ra6crB
5ql695ZNWow1e/r4Mr9qQKz505ocO/tvqNJ5LUOd6DWTmTETfuwpyCZsy7Z5I7SWMqDfMkjGbc7z
sCHr6++EoJj1KTz0UAguRQ3PlQONcFKcBSxvUBK7MKS5XKX2pZp3GV3v/FgW0rUHt9y88ytymkLi
O1ofYRazeMInOQTRJaGNLfIrJVtTCAMPQCZ0enWOeuf5U3A8QER1qmDuVlgJam8v/LqGHtxip9lN
rD+G1ImOW7g6WQ5s/g3MXOsMYrnuMju5cjSNnrVBL5FI/h3LGLR03E+/CVg5ke4eIaVCWNOFA4dN
Jp+WT/Cpj5exxs6jQeUT+/QOilqpDs84glTVfxIKd1cSHNKmIUvd8vRFwisK9GMx28+miGEj4YY9
a557z6dOB1F3d9XfY2IDhw9Hl9OIwi+IPVjqllAAj1BH1lDfJ+/RtM1sCC7dj9idDq5tarPXThf2
dU6muzEJ/lKqpY/REpn4HDd7Jl6fjlrB6f1JV3fokXHJ9i+lJshGttpmAbE/+UuwJ4AuTQNTTwB1
E8dYyTSKfQiSivi1Q5HMk4s+kiGAXsEIW/bd4jx89DzKbfTQpa3R78tBTvxaOMTsk81sk+QAFqIQ
frK3LWbbS/j15XM/LT+/Kr+gDe1s6OzgjFR61PeOgjj6m8SC5rgnULxRPdgmwAbSL1n6kC4YreO6
+0u9bij6zSnulFcPSkckWxSjCJAr8t8QTMFhThUTPLS2sny0X8PmQLITlOl0KkI5AWkw16DJP8RP
kKr4HTGQLumdh1fkJuIvU0/YVsHMk0HmqKgRfbGGyDFD6Et5HgMaTWfBPLBEkOtt9zdIOvI0Mnh3
4iQE/xCh5ie1Ze1g5ksJbZ+skJ3/oFEyz2VVAv3vrHGYb5qt7jMBbBxf71OGeG7f3OZEAEO1UGiY
5qbZRexpDh4aCwOYw5cV8pDPYazQ7rn2GR4NQY1ldgA8yPcTwRGFpu9y5ZsbVH7NZWcfF9KgpatB
Bt0VKtXTF3kJSbkQn5mowjMfTUGRPtywe0zCWZerGbuPd+AlOeXb8JlmerCc4n/rzsokJVoMTmXt
1MAHy1sTY4nRiC9P3+Bo/+CPGiD06XhTamAsXhrSGA0BDUFN97WhXkQqcbtbrDrQSqs2SBMMZQNN
zzGSo8QGq9DsY+YkfQ+VLqfmoxdilcxnTsjaXnMndctpTxEnS6Pn7kmBQGTkDSESLsGybT/7aCs9
7L6FPWzXX6MPDdgnl68W772bUvOIpv4C5luC3FyUmkQRPjVJ8fux9OZsOZmQk8VtAUofNFvNTHnk
jDmNwrmXWyX3pL2QULlP2F+Jtdm4TwTxwntwMGNqO0GztU3gBdt+iQrItPimaKSvQwFVrSt3qZ/Z
1aGkLqJEUWVgEkl3gtk2z3k8AFBBpqnJlU5PCl5T/BIdu63mdZyr6lXDtut1/3EjKildBI3qHARX
HkZ5hKWilFb7yOFfwCZlJoNhGiImXVfodk7U8mVhQ7/ERcQ2FGYikEwaWh4jnoko3fx7t6O/OmlO
1prTGw0wVhJwbIV7D6MsfvZD96ibS9sfx+RMLWb9iaJ0wPZc8yftYjC5HmgX2BEbEFjyThz2KK0a
rpMA+nYWc7IGo2cJsWSQoXhZAPNaHrlGuPo1O8Qz3FmNf/UFyuaT9HBppE/iwDSuM401PtQmMfwe
J909B23mW5QkJmn0Sd+dbn6p0J5+ZxYeD1ijpSBxRlpcWyfN8fG29IY52E8mKryE37fk7jP1PR0X
kAyWnN4T7oO9ZeDz5tCo/tkruz0ZKbiF9nMbyvlCA399AIPGsQ4PO7h9odLl96ivZg224oxW2wQM
nZIwVdbBY7VSQ14r+AKaqYPHzI5zgO5C2hSmsfngOs0+C7TBw9uQkgaJLcvZ/sLYi2+MxCbCr4KO
YFOzUEgGHGdPRLqWcDAtslJ1d98Zb3gPb85CflfU+ra+mqgMIwixhjcH9sIuQWMcNygJst317X4n
3LVwKwJ+zqkVPHCA5m4/OmYkqO0HJkNnH16tcrsAcOmFpC2tUB2AxEooQ5qCH3RlLTf3/7NdjjTE
Yt6Gte8MrR3wI2R8oNyrqiJiA7evZ+wsYQprvOSqpoXk7Rr8aAXTMf16a1t3HE+gI/JGc973YpAD
YI/n16PPmAdXws8vN3F2hk/uHzNc4TWhxFQl/zVOUV2SeSk/RILKvKSN8KUkSKSbZQ0ehnkV5V8a
4LH4o7Ep9qURKHF6qrluzccXjDQ/mNm+TAmlLSfCVcVAzXyuV/hiB8ChR6Uf0dObHw6psR2xaFeI
IWC0G7XczVhOgAQpNKySUrTJLnza7Mqixc7MASrCHKJ77rH01+Pui1d+VKz96ezgQA3fp0groGXj
6oj4kf3aUOHWoourOMZ/T9/ZI2jU+I+P/ojgA1SE/AyhbnGQ0wAmj8V5oKm5JonbMOrEjB5OODu7
e9oCswY+atK4ZSWeQ8z6WuyzFGaPMOT+mQhok/45YBp3cRur5HfSnvJVLEUHJRp1mA6XfVK754rz
/walaPu1vCFN+b8Gn4ZqKmTZcWXEldE56iss3xa3ooMlQz+hUn9DGozTzkjKYSuer+VQqngzpanj
lEE5Fy7sDFPAca3wXFWEF08XHyqfuXdkwUFVNmNMT8EIrwooqRLmlvr1RsvQhLSlJz2R18L1OvTY
MfhDQpAGyzRhb+2Im+xstBuGDRcgAExvvOK9aaVd/stv3AaEr3ANNGl1W93nwizvdYhvKD9sFOaI
zC8utNwXHEijNpsJOKDbUYLif3oq5FCaAdr6BeunQLvl47t+GlApZMQkGuVC2L9/PoXZwaoH+VK7
aPS/3MApCyav1su5HmqalLMN0c9ItV0nq7fa0sYF5Xr+QkV9VNE9Mgwfw9gsRiOyYFlTeMSGL9Ou
7SLj8/z7x71bRu8DHThQcQf/3ABJEjc3M834HebNdPTQOrvzipBdJHtuCO57G9BbFvDmb5gn/y2t
1cof7ZyMdnOSIvq/8yVN+hgHNU/CkAgkoiWLwSEgKr5a/KW//awL/JadwHYl4/9g8lo/uqA+EJnS
pjP7w9/KettGldnFqsjp4G/ejGLjUvpNnhSv5FvoVP/lK8NFLl5ewZ69VKAaL2UwqFZ4EQUl8mLQ
pHliyVgH53DDu2FnrxUprFGSgiS53WYOYCOqkGUe1uEOpYxyR5g0uTpK+9mXVAC1WBWskCDkcLHM
pw0y7YyvKXL4uFeEhNItIiVVVoHavJ1OIHwMTGMxMVYUkhtjIF2hGKWXNRwhxKc7SBg/G3Izk6Uu
VWoRlhpG3yjq3bXJks/lE8VbLiaaJ42K4v7D/YF//mnk3v5SoZXkG1idHEnih16Bn717CY39BSDO
uMtjVFI18EnLj9xdkIrto6twwPeWsPamDbu+U2LbQyLPv4cCg+dO35Cq/okyRg2ZbgOqmY8DSNrR
PXpdhLXz06vNkMMhN5+Eh0QAAq4ff0ccLDm79m+IORKH67NtQfdp4Lt3xY3d0W6A4lPlulRTFowf
9h3TYgmLTBZ9QpxarEslXTy/I8LSIMTJKyj8DH1zBNCURqhbQXi0R2Di5QnEIpLBIL0n4BQj7lJ+
AnJ9uR6Bk1/vnNJn571zSFYu7oSMQ6ZfY0oeecS1G0mqA5gIqBh/FUNs7AkLOh70etzW1MAkGF0+
/ur7NWKr32xJGWJLHJMqJTFQsv0TPyhduifff2J02TeVHiMyToZlvqX/TKu5x/m+mXUBOMzdL/LL
CJ1HNWCOwWmLleRefhWkfbvm89W1FNwwpadRupZIOD3COESoDLorZbrS1atbUGc5mBL8VJopBAIE
tX0ucBVfXIalU1JLFY4DhS7mogLg0i5jn3ZoaqTHyyRnQje7o1OxaYfQ76DEXhCV4hQ0WynlWqLu
ujV8BNYBLzM7uZhedBMg6FfWiGogLtpwTWRhCWjZGdKLPMciTnoil6dXKBV5wab/44D1MXIZE9c9
O/JUVEclZsQMyj3I0/qvS27zOys0e6fTdmTPCYixe9CF//WNUDzFgiBu2rNGyKMH38wX9GviMXFR
mVLJSToDGAg/UvJWwa+CtEPSP69vCbd2oXpYpCwrvNHxzNWcx7oY+V4jcaJL8nHsIHPdk0u3HkYB
1AfdUqC+uyeeCU1L5/4+9Z41NHMhSLi7RM3YVMUJOeqJTpksx15LDfWfkezhsk+OvXx0C3xxw1TZ
qa6BaSJ4zd2pTLOp1QwNYGtlcmMwKTW2kXqeQaatd067dsNZYBsOjvTcM58pCm+4j8YPkGKsjKZc
TUF53xn8ggw+EEMuwEYMFiztskN06fBk0d6jNsy1DAOb4EbkkXdEV01t1ysVc9f9wqp1jOVMoAmy
w5+Hphzn/3SI8mQyT6GBccdneDP7qkQDW+f81PiJhBl6UbYqz5KsSW2m+GSGRTEdKdKv2uVPzPb4
cguXEWzpqlyIcIM0IZgjvRXpiGGf6ddOkcwcU7LNs3ieMip8qk4GeBr5NXlf+NVFV04mlNxuEsI7
LONXDShtU9q2FJnTefRwip65/ADRFg5lLCUgQr+OnBw9G2Ye2sjLw4B2aHXyqUtCdoMAnccG6LX9
kXrfwclREDGDKm5FYlkiVPoCciE47o76MnVI1QKkHaaJ+YzTDwIzTzkEVbOsrrge0BTfktlwBklS
yeGP5eEzvdgIlVa3F9VNe+xJwgTViWlpZDlgRZ1vswgpJFsVCoY6RNGHRUCTR3uAT7RJH5bXRk28
aDYG+zn4AwhOuvM0FxDcsmOX3+Jn4cpRL6UJR2QDyvmgzlInUrR5nGiKbImih0Z9BIF+kg6BYm7w
gZ3zyXv1xY6XmCgPx93yf0OU0ld+dfOMxUb+GFlHUnvVwiomOy44lTNy2OX4SLDLN3scBl0lv/Nr
fkgQOjqsJYoXlqUJ4pYxKBsOVsHQsqd7jepDkiNUMlASLyoXc9a8odY4g1+BKUZtMhYfyEbJf37H
rH+TCpH4ioqQKTZIib1P2cXFxLw+sNGmC3XbW2UycCXkGXx9jGOXktdw3j7pZUUK0NDhXc2366of
+B4Hky8m8wYEgCVA1tkI3T4WXOPZRN4FcbAcHg4g2IjpwhSr7smGL+9yxKe0I5E7GbLwEF0U9FqL
9/jeHU7r53eqPjZrABBQ2ft5OR/17RQwC+tnClTArruUbRqJtrcQYWlpD/kviOCXBGSFE+FztiNb
+fvwKdlwB/lHB3Gd4AlsYPBp0Xdr3XwbTWTmn62nFRCZi8x1pxGv+a62pMPR+mW3UHIm3E/Zj9bc
R+0aWBccLFascNeUKawd15N+z1FemnLft3+k9gMDIMy/DiXe+sESc1uKT+HXqgolVNXNrEnoweIX
AOpBQDIGFrWULH5BV2s95mbqGQcsnWFo/t4gyToAc+iwlXlh/UKm2bcz8sVdEoJk3zESnJSSHJmM
9C4RGOeVPY85GLXDIXQD2cqlHp2toa7ISTA+xYeIw5wlOUs0/2JQOHZQj6LDJCzx8cHt+aBdmtW8
MKDKqDRp/uJmC8I/IxfT56DXyApYAYy85xkXi/6rw3ZcYFUVLz/VbpDIiOAod2klAZi2TuvADL8F
P3cKcEhRaguJ534SY/maFRR8PPNOwBhk4GwkkNU3vxbDzHIL1jtQbqyW67/GUf21thsimaEMPo+y
r0HZER03Sc2GzlWqFYtxj0MTinN6Rw5IKcPH7LfyZtFJZDEOP0fUE8PzZZRWssMaQQ5bUoIy1OCO
/156tqKU6ANxjLXUkwmzb72Op9OjQuN//WG7WQuvqCeRtLZ3sOcsge0+1C/1I9Mfk+S48PFH/Csk
uP4RfemJ6fsmMZ+Ji7cc0XohB/UDAoYLdCODbHtkeA+kP/kPmSPj3tHNO/M8mN1S1aWg/mVgwUcF
WKQUVjCdHW5zqEbmZIIVMWyYZ6CknEwU4CU7CvbahubcXyWgjEfEZCbc5A4JviowtVyiXImwZ7FG
JB55g1qJ+HACt6UT/B6DXGE/S3zGTZKIlJn37f51MCsXxwkZyDISCMZLduphSeOPGhCDIinUMgPL
0AZgBB7YU5uLAQSUhJAm58rFDibVgT8uXNqSj0pjHPZM7z37/1kVF2WjWjx9am28lxiaWpwc0F6R
+ZkcNMTkkIACevLrGW6MWuCPmxvY7DKe+msw3Ud7hFFbe3dmONXg3GCQl9vwPf2e+ZERYAhN9L3o
uzhliQFjyB+MPQCDuaMZ9uSsqAwKsE0fw7gOmNqhQ6Antjww3gefiYBjIIpA8CW4LWXhRakxiRAt
5e7ruDsT47mSGd00+or/dlZagoxxLZE2KfhCQGXSpytHW1pgbqUIem3Mwn3s2EgekUVWlb1vxR3Q
nqtmhGto1pEnYrfnFGuL2qONGCwmAfQpMmR/Ri0PhDgWeh6QFCExBVFDGCBkKbBJd7l9//YFgisz
5isMxfq3IZuOpMo9oUUse15cP5ff0Jb9L1y43tN3Z8Au0wkvxUaau1db1LfZGGIyKucniuXQL7Mp
jS85XUhwb2aLO8TPIVjl/o1I04of1j5FdofQqGVW6rfWqqV4lgg9AGA6AY4FU3TmTgMqlgAkUaZo
A/7eMRY/A+r0523DwqUHEwULA7YVR/yAPwiTrI6Jc6EMQU+lp/CcjNNKgXzvzuthMUywmFoNdlo0
gAPuzNB+o4/yfhl3b8PGKKmQJVjc8/Mo7qH/n13PN37E3x6QS5+kJFB9+Ewo9avkF8E/ufRDVnrF
xJ1nNz5QoMfgAp8BYB0AdxAh3CKFWW1icwd1onmtouq2BK9NoREAFK1Gx/qGeId0Mu9kUQdFe8sQ
qO6zZJ24cNGQZYv2mGcrVqTv3gGCDdTjFfL7wlad1/TkRZAk7Yh5p0Mgmb76KQm2Sa6EpB6z/Row
w1egHOLLB34jy9l3mqS3FNd/TjSFU8Ma7wReHmuzvjo7xMTK74k9pJiQzmU4xXe/K0TdkCA1bPZf
uVN3smx7NMp3Hyv7bMELG5r0byGh1BvVsOPaTuRJZxSU/PO5Be4/IzIGal7ybYgY19umhnZE5ZZp
SKOyVmDnu1KnkhlTF4ZvMWCIUJhkiF/K0JUeKPjYVmvZ2c4DzQHnwqCKvSxOwx8U9fb7SZyRr5TC
1FnHJVhlrtFvJkT4GZv/vjwNtCRLFMtA412f9ABnYaflWGGYFBpfjq0VZz2VamPcDTLt7zDpSrht
UYKyIPWyOMi328GhZdr8CEd3PLJei6nv3SjdguWnVwXIilwQVFLXq5SnaqHuJfbhAPfvi2TZoTYu
rJxONCQT6nqDlVWsBVQLGXrdPAZXs5fkbFe+ot3TiVEA2zpVX4JtGfq/YFo8yIcXRHBncj7QLMk7
lOzOVoF2Hl4/j6FD3Yz9V+zUtcga+ezd7S7ecmegNDK/TpGMvWDBwODtB/cdUAJZts1HskbLGUaL
Pw7Hr/zAed5Wxwz9jyXekmX7rKreqxvksEBUg0u7/z+/5eLutBMpFoXMgHLJ7jtdyEW5TZyA94H1
w0fxDHiNeVGwJ4/TPxT0uLUbR5aDZqNCvjtPR52uU5QZo87WZG922Qzi2y81t40irs4yHHxMo2X8
pADCkr3jTTlpFwuac6353zq2Kog7YjUvuSmHxJIaLwpkFlo4Eh3xuwjhFkNNRqw7GSABAO1mD5lU
9LSfomgYq+0y67aa/05PIOJl2n7VnO+qT9ikGLs0070tKq03FNpelDuP0KO8LeEAryW+IeRAcY7i
Jj4W0Pgj8uA2v6xCOIIs4h3/tV0a2C/zcQoEszUvwxLMsWtzZmv6dPpgsecxNthLWZ/0db1RqPGC
DIanEMyCTMoAeX6qxw7gJaruOOjO6udtP7zpgcbZoVOAVvnLQZdN8mmc6M+EXMoW5gsZrSZS03Oy
jq8iGSIca9OijGR8/H2+qQq0Wv8uL7dycxn+3xnWO5bVXVBPlKhlm6rm4oiQoqUXoqPA6Rp/CDU4
pUCTZUhc494/181FUXQU+6lDFWepi2QJpu40UouZNv07Ij0D221pCgIGygEWAiokVTkvOj7a1sT4
bK8HhyXtv/LJU5+EEu9fnSxznTb4xcNonUVVLGMXBUoAguWZyGTDyv7xj4hA4AHakRXM9CUHA6x6
WZMCTNGHtD5FcrTwFlK3BpoXzxiucwkhZ+YmqkFyLab+qumnFMn16LMLRZ6dBNGHeJOvpFeTOYlE
U2m9dwwZxCKUkbfbcyhHUssnnH1zzsWs6+QzNYWD9QOTmK9QEF4jM5UOAIBQet1v3lmkH/+tnuk0
n1DTZ5M4f6vQuTYlLrTZgIexuRMK05QAswudUR6/ODv1tNdnLMtzGXBDwQYM8GlOhETO4Abd9HXv
dRQDIj2g9m/miVrzJ9SB+Uomxby2cpA5qLSJXrlzL/11blBc1JWfo8+VJnbbRyC9rW+f4fHkhOVK
nQwe+0ufMf+NCETROgUBS5oVYmee2hjkNVkIfVe3ojEywkKB+oIdUTZWaaBPcLPhRf8ocAExU2qm
AUSMBnCePtScALt98nOT8DExs1XxS0HizCsC9WDGPW+8+npy1zeiNsc7o8gc8d9gfzTOuM7OucIF
16vI7deZYnntosnaUTuOrryJnmkqa67YgicTQhGCQqma27yFUCHXklDEDbzsPtT9hg3OhkNowbRZ
sS8xvdOki4/zsOg7MXRM9jFU4wZZSFe+bpLgOWPrMogaeFaEi+HRDLkGnygjx6807qr/xX521rgj
W7ggsOvLJW+HyHmDreXx7eTL6BtuuiV+3vIjrAuErMbcSXESbyXg00ITaz9vtgMDSTUZ27/QrZHd
dDC38mOkgPGPi6Eg5zgHXK5zBeV+Q8PuACMPWubGl3Zm9NDLrJKyO+jKzg5f79EA2MUMDxHEH20E
UQ32fdG7zVPuxoHx/D1nICIsKcBAeryWnsKYvv9Jkd4QJduISHjP+TIjNEl3iip8+e0GM9APz1ws
F8o+84EOW4QfrKdGdySAxHzPgYtKai3k1pBzu4+XvJdi2o8+NuwiaSoKS6wfjsg23REqvvmonxGX
NyHdOc+yMTYi24mQUyud51Qm/ldSgYOjxkCd4YZruST09/by618sUQz5xtdFawsO/OsMqaJilkxa
JTA+MWZ4iYoSl0OAhus56WvcVSuXliwwEv+kMX9nWpOsTzJ9gckTDrCR3/yl9P9Ja9RndsRTEOrv
E/xVb5yD6BUyM4+cFLOb8FxMsRWaoPs3ywpDRh1hmjuXKkD8VwxxOxdS1o4G0ZZ2+GQXc5Sxj9xc
7p+Ci28qn6gUGrH2PmGTKcgW4Z4cXIkZDLibSDUjmPojfrmadgwgzKcHrTiQWtGQIyW67tS2jAX1
sItilVk2D/KbLcolwd8PILE3uGsdin+0eBaG3yIqxiIJ/pDYPMGQSjqeDwqBz1kaQv7Jl17GRb3G
ftCAquHvH2FZhI2SBcNBD0S46iiD+6+DtqFlHGspkiyrZbSeX8RAx+BGOYCYRQideTl+RSfL3HNP
j4sX5/54zPQWJS23wrnSphWAaWKLWTLNgjFCkoBw+V13IRfdpNKbX3uKFfxJHdd4vEippOaiG0YU
oL3GtL7h3w/6M/smphxk9t3gTUEB6WjHHWsfRsTORjeDLSvPMUprgqxjP0281zWhVfTI8rJsfHvu
q+apojI7r8CCJDxY/fW+17GTg023QouvARXClYziFKn9ZFvovpnw8V7O2M+szlQo9xDasttaTZxq
IIbCTNlzJWA/zV8HnMxE4/+x76u/ksr/BAEN0YootxtbFM1rJpR7jI/ybBjqagxxSZlh722x8uHy
+sNKtjS02nEMVFd4oFVtumqqOfNn6A89NwVUjZGcLNPTx+9h3gHKfSgFF0RebWMBYEurqdZ/Tp9H
Qptv6+YF863Z4qkfp48Rac4kgbdCrUawlW0EAJ1Fe2P+bTWjKP303CrcJV+lzbdL4V7MFmwAjU8w
7XvyWzdaZ26G/8mfq2wI/cJKW1lc3p+pS3ipdWx6MaoQEe+lk3hlZtU7UM/fvMA0hBj8ZHEgNyKK
xOPcGqm/ZRIB2X22rjpVAFfHv7gDXrpcfTtMl2sS1nE7UMFJxtCNyYip/hwLiJVKL75MgaqwYABX
GU/ARnXmvWUvXjtp6Ce3LCRXJrG58mKWQa2yNKP1hYq9sJkM90MVUg1EScukIUa5bsBChql52Z5X
o+JLCIosYifqiuJpUPleqONIYH3uLyBjiJtHHNCXHI4iw4cXtj6i5cNrsm2jVFTpfWDMjVFjG74p
qF/jiytdoAh9cejvryMSHK9Si8RXLBED+Ax9y8CiHuD5qoYnLJHk/RPbqpcxahmn2uAeINZsLHzI
Q9uK6562HFdMB26o/6h/NP0lSAGe/w+cRAOTe4HU4DkHbgLUFUoKN+AnR5hoWZr5bMjoDld2z655
7u6GLPaz2rO8BTNJtVRykBayCMnqCxwNopQqqdVfBa9SEiL2Rnx8ifUoQbQTcImEl7AvpgJJIEo6
hBKcaXHNxUd19IeO1e9I/aKiE2gH5ZjDg6yfTS5JvcJ3oq5L21kE8xuhEVVolN41niosNev/Vdoh
jXDL7p4fNX5zuYO8VH0gQxDRmVNdZHlYozwtPaYRi14XcrJl2X/Wdmj60Sbu2trjlSGEYSv284t8
5QYqGFzNAQkF5GjTVpcMyGSe/J8JqvGxz4nM/yXCSdKb4QuT20mj4JOv+GwXMeGcxWBvR7fCu2mn
edXD9pSnjT7uoP7dTz6IJ5rHVtHURzFeoBUsIWU+QT8APQk0DUrxqLRwCyq/ZuX0gTqx1obsmVn+
GLhh19m21no8abYxm92xJjIu1R4OP5oIfWsFywklyWXO6RBO7+6im+b3HHxQd9fkMGHVdwPEg52K
HegjDuvsLepNMxeA2oDDhVx9F7KXLrlW+dRD7yCrpwR/42VPseZCuAKYTdsjihKphEObWasZ6lGJ
Zt2y0XsAHIOKRhR35juZV1lF3PxqXOf2xvdXi7fU6CpnEhCaUrImcRXwATNVGCefVtlX+RTb3Lol
yu8zIlS070G/uATm4ebgxg0Sjvl9hkOFIup4bmDal4/bZ4AVuYwbGiY3p4jMQvTRxmNxu0+heNsl
QJyOZT/q/T4bMu71cmFGedFeM4HUQypO4vt6P3oP/UC7IiQhPvV9B7lCMIoF1eInIFcQVYmaUjXl
i3OWIDMwA3bbWfryYKNBVPwNith+7xRSgHDNO5zM6+Hu+oOFJoih6KAjusbm6dlAIJ6rR9CKIa5e
4Y/D6x4HzHgErk3o523Rho9GmXXxSfqDBJnyYu+XDdSMruDu75zF/7RdVSlUwAj/QaBpR+7Hu4dN
oxqU7vAq8N35ns6SQgsGlfgp0mACCwty9NNM1fHP5cLVVjsGBt2N+NRe7V7OA8Btfgey07NNbJ5c
sm7XSQcbx+TEOTyY9KrYLnhw0bmTPNK0GtnEWme1o5xEr4Uofk8OAjS35R0/2no6891QG9YAnqCe
M5t551TUxE7A1qVeFsdY8Hm1qEdZqD5YiKApc4deKfuMtmpKWMhhmQLdRdFA0cYBhv/It/AYmGo9
rc4Vip22DidmOytyigu7YhRMfwowXA9rjnlgPr5/ofrcKsGsWMxLcdGtp213AT5UdMIdnqYvo15u
lv5NtiMxkYDbYUZ2ZYQ5LWk4MCneAqMw2sQ27VuNX2VQpiWuzpMgEWfH783f679ELCmieQ5CI1AM
mf/rpIfTFRHlmDgbhnOaYhYM5a2xrEv3ZZGwoQ7gVBlLYEHuukKMXhXCBwk9tT/wYFAx+FexmehT
aDuVHb1kbgROFJnbBsROrnMaQCS1qQvNNU0xDhuFI+y407pv+L3F9tsy9oFzgIAJGVM+vbVlYlw/
aiWar3bI+7V/81F1j2d8jhRU4fBnstGr2xvOm/T01QsF56PwfGtoHAfUGv6gQQlVjiK7bVgf1BZ6
gshfajlJwVnwcLbENXCeAJ7O5l1zmRI8TkEV12lyXVH7iZvc+TLU2AaGilqn7ngLwnGsA96PgeNz
5YS7OCLx9GBXonw1F2D/SQYuVascN/2+kvijHFxfrsPaPN1873wM3yT9uMSRmEHwhuXLidLA25wV
IAIwCyBYtW+TSDtILea7VxAN27zbYrPSsEm7bUviYaupLt2N8OH6hnRZpmge0N0W7K/0uM2JK0RA
uoryiL3dcJcjqRqyS8x3OsOivvYE05VrpKxtEYizkt1slfaTGY1piXBg/Xk9ypNPoPuAxoXchNz1
8hIPuvlgolhuUXpmtgn2ttbZKwrZess4Pnq0q8v0/HV8FMOdiGshQI2SnaXJ7kQ63ykQwqZDImcp
6QY/8sov7MlHLwG5zJKiuWgLwxgNc0bSdJ+ERrvB0NGmBnRbYoby5dxGg2v40eMgccQW4F28joV6
iTOgVjnNbjp6oXIbqq2dAQjyy9JyxE434OUZIzBELhcidnZE8wV0u4Rw44/kBvTSDxX8qUIwNbnZ
crw8KggKOjW65rYDFxdMMz7ST1rnsQCC65JWdBvAomnKcBQ2pF87dXbbBi88hZx7uQDd75yhI0O8
VhdlXq53INGOGAQgoKyxpoEPnYuJou7RrGEOYv+4RHUVpds2oMrrKeIxyiC1vQQ9+6bQ+pdSpqH9
18mVEUH3CSbvUcLGSS1ZGn3bXDO5HCxsk/z3o9sWZNFHroRAnfr91/jgQd6A7IoWk8qJfnAo4+Cq
FHs3U0zIarOhKNalJ2ME1WccQ6+K2+tuGeOhsrB8dSaTqdGejO112q4qBi0ewrMde/UcxFNHkQa7
DSr/9G5Wp5SfV0YU3BHEwogPqjnL8pqrz0+QbEpu0MNyv2VySzzNjFelESCccXz+u6ye8EUxsBse
/fwke5VZfWLHGSbuZ+NWVk91FYAsEmV6SZ4GWLuZ8YUVQ1JxfWbiol3qoXiMHj6DP6s/xPKRP/hM
nkEMHYAWf0B1DNlR6byoI3AJBEifbZ565u3LOOgVoIiAiKHF8pbVnbRrvjhTAa8dqmctCAph/PeE
+QtR3ijbNbzf9yMg8ldTR4oCb/fosDnTOCiA7O+e/A6Efg/S7s3JtaOiOLXO/oOMwwP7BDwn3XNh
GuQN/yb9KxgzalSq8GlmN/k8cuRflIbfN2svaA/cNtDCuAhSyc9oiLPbClGPcSdmf7tXbeNXpzUn
dee4i36Ykxk/zu0sLj5Zgu+odWOct2qp9hXMD6fD4OFpIau09xC8DVOaL2qBeo53qLexa3C6qWkZ
++8OBU4TEYgwryOcf9zzL8nyZWnMKpXBCSsxpzLYQENUYzAscdFVMKTw12ze9kIr+cwnxdJVanfq
Mbjrpy4Hf2pGaCMx1BzSWaNTo/uQFoISjPNQO0+fbpgGZ6Lvvj7LLjuLYr6hgq7uvEp+JSnIXO31
7Zg+B1jaDjr6I4bjiOTi/L+BmlS6yg4K84LCeB5NCLe8Nw0xMTz2vVRJOHhzu7dC3j4Fmtin2RsA
tOHJPPIbCdMXVazpr8tXIIVTEeK5A9aR6bvFeMYdTCFB5qi6Vfn/CQb4ECVOBVX5M3rCSyzbCOTh
+iSceEFobvF3oQqRMWoAfV4zaKKcG0qL3RqwYphsIu7y41RjruBD492vILqaHtmAdPA3NnyTTC8q
0WjcUtmIv+J3CcEUSghtGwVbTOQnhe1g4+ISShijJmKpHJ7mhD7VriMAhIwNe4FfTIG1Je9zqn+P
9qGQxthf0Fqwx2NL9cqZr3kvV+UG1WkTS7a6dRGqy2+YYd2G2BHBTjG8tBlyHLNlxDfqACDPjmFi
rz6YkCITzYjuJonc9o1DZvWqFO8N9XZ45Rqw6VkZidHxFBgoHt8WGoXWmRiRVN0jCofLB3WoNuQG
182ZtqNm01s6B92q4paD3+bgViURpiTcL37ZIGDe6rE5xpdjCI3XKgLB1s40rVK8hqEC43UHpKyd
zrr59KGs90ftYbnQOsU9e8NWLlSv63WNQGIWdYMUGZrUuNqvti5EjhOVnyKcs9L01ip4s2lbxawe
mSdKq23p71hfBmUAJQuOvjF3kfXv5GZGCKHDzCKPWWgVExnFZeJnfoCv8sjEc+5gGpssTTM88+5h
M/jQs3FBp1+i77GaJewqoS2SO4H6+gTL0pSP8tOu4iNez0fGiuk/5xC0LEyybHJRInlprMPp6jFl
VznG4Zg7XYn1DFyRDC2QtW9pjY+Gizl5//ZMGwT6Ji/+auqM6MFgYZnUNwocIvVV5Rb/UZmbHjSu
1EUs6+zjh0JdBFj4+Lw6xccyfSMNO4Sxee+dKxq+vJQa1wmr3n5YSiIBZVzU+VD6KSug8DP78boy
K2ytQapfdx3Al29vtYqesQVbLiXP8pWz9hu0JIMkWwRcHX7AWFXDLdXLv6fFxoiH0jcxacNFKZv0
9Vpcc/FYK48kWcy+j7qJnSlI7d/c0hE55DLb9DRs/Nhjaef6bcNidXqPI/xGs0FtCYmO2lJXTdUw
UjgM5OBgKbNNKwVVgMi2Fkh8lI9S5MsfsyMq27gg90zro+Q2dQTr5dvCFCS/PY45j7j2hF9Y8Pat
OtXQKXormxsLcZcP44gR6oAr4YtYL+6lCSbLdQ3q1QCaje966YaG4qvXUVR6XBO8Hze0y7bUOQlp
WtghcoRmY4Amzh/q7dGu3AB1fZ7z43/36KdbPWPjEGXaltTDeOUKkHibyyy3MDQdnvaWE8ZIQCPb
Cly7vap0bn9r+uclFqPE+N1nrfxyN36uriCsspe65m028R81dVlcwrk7DBXG3AeF1SzuGhb8PCsr
OJxjaf3Ioldkr6d4FkBQzlyIiAE4lhCkV4kheIa/EKOeMpzm70jWCCdEiDhImVF/v64310XTfucb
vmGSpWl6HzRl2D434DcyIfx4EArO23+MQqaMDQeBP0AzFQcoF7UFqSbExxckuU05nMaUYGspq0zO
zsvKJG7esQSpO4wvrhrtnynorm/OGmCpm+GOLTKJHiSCGZV+Pq832e5mjTq3ghSqTL1ucjPu5Y6f
nlqizRhF2LSxb9hSGe8UlFij0BVTPJFAfBMEeJVIvnjC1JG82NffeDukn5vhXLtiMrbzD/2LQWyj
l6eIiC2Frb5UtF7cuDafXcss8Ts8f1vhkLur0kNAunxkpj/dd4SyEm8Nd+hl8kHBOqatVCXeMbxF
ivb5WspOyBSkUXLnPqbAe5Hh/zyLNU7pZfIJ1JJkfGDF1mRp1RdrM4eVDfoc9BnKA/v8eXzsCWvn
FibFJFsy4QPCxWyFetxKVgIJS+r0K+tl/b5Lkor+uw8KxfHmZnDdlymzyQGyClf9KqXYyTi+sFwd
lhKIeuxiym7ccIKQluwxFQjyghc7A07HEd7FcFF7EQLTxGLQHAyouo4XfUdap3rAxyt0VWcSrhFR
MG5wydlTm4L9W2EG7LbQ4RGiEBZKBuEWp1stA454ReH+E8pSSe08vx7eo3poDY2yBO0tBJQ+5KIb
fsPkL3DcKzCYQHacAI6tO0wtkyPchCC1pPwkaS0ePe+q+6FXD/s+GevOGwWqqfuu3sic6LZE5VfL
o+s/Y84fjo6dgncS+OTCScB0wO2srQwUyoZa8fTnxk4DTZkpmMUhL3Ib4yWw4SqGnN7ASNbXqz0T
kmK73+ZgOcosAg4Dg0KaKWrnoRyuD9V/VbTtJK3K/4PoZ0qgQ6l9p76SKwP6EuPvCJDTRKROGhQa
6BfaPu1E2ZT/1Rowj/zlJJ0M9eal55D7kIY/Zyu73ck4OG5wFQTgXYZjF1RnSHNBBd0DokX8VvEU
cj3cRXtCGANYyHI4fv2QU9d4tr/gHV5EyWdfE1ddnTLeWXQ4uKwaNUNmfqC4E8ZrbSV5p0VJqZTM
y51G6yFWtBg8BntlHgw0HkWDKNcOv81Gr6AfnU7mFAQIdYclHuwGy9fjOFdXR7k46aLwuYw7rr+s
ZniFVk62KR73g7W66dtPqmHcr1yfKCTfmJuMRAi1srEV/MH3slBqZj8h4AW+DODw4pu9152ZOFjW
mAib1OmKalZE650muC/08rZdfGd8w4A0rU2Le/VsutDiAQPtuqjo+2+UH69L2nSy8uv+nObZzJu7
0aaJQx/qo/kwHOZbiVQPYCcrfQiNy3wx1k34jFqXg12XJAJ+8DPvnChgTN/gooLDPZN5QKQqpal4
3mzvBk9hwupFyVu5w/Hs/qc3LcCIS/Zi3MzuBA7qmXabd1I+AflhksgMG4gpivg4YX0NgKqDLPHJ
qgM3L7uMr+e+W4z32A8h6mBFJAdHnFMRB8OVgi+2/kGrEMHgmpTl7yvXMHysU2aep8iniyme+OUF
dELJUvRRzYxxqKeSlrKQHRHjJPtc1XJrmQ/5deLPSTYsFhJmaixanLSCCu5zPZNktfpdCI5BoW/Z
upjBpqq1JBHzsAKAmWspeJHGBeMygseXWv3rUIqfdyGk6DPt8NB2SehlrDh3kO/nsDxVJd2yWPs0
Qp3Kfh/GXcr6jnF9wR/9Y/vVVM59wD4ArrM6vkWMvcrBhkSWK+VNANDUj1ZZ8KtQ81Ig1vAqiXBD
y8BaojMufp6IBNU+aoSWzi/QCeIK4dbNHrsLuDe0b5spIAwKH36QPBSDs635HJ/oK9ffPQ6ZZpdS
KmBDXJ/hYREDtqQEkvvRaSsP62pvEwjzoEYTTIWbTgsXh72JZugKGYpBX7PYGRAV++nBwgV30FCs
kXCPGxG4Yf4b3ypguFEPQrR5voqwXn+n0pZt6AN8QYLaH/p4jsCaef3JaWRFiW3/c08vwKRXgc0A
3un2jbYpD115oN3iL+3jTAuO1SotuvgNLbHQkX7ZbrX/cGPUXUplNR8pM2qDtEFX2nSGzCo8L7Pz
3jqZnHTngywWHaY5YGdaIxJBl7BqSqwAWsWONV4FCR4/c2uYZOUdVc0TuRZwkpbheprpwuQzjHuR
bqjGhdZiq9me7kVjP70jDi+oqHYvfnnvKFdKgU94UDbPn6cpoKSeX1AlYpbLikKckP0B6sVXUf+r
r8uu0JacdAMEEPqH6RbYdUrpgGyBzUoNiQC1AJa8dWCgHM3vMOArL6MsC2ox6nGH3injjz2U79mN
SIwBdetLk3qU1cHI5qvlR5vJZoI72j7eeubOHwGd5pW2iBmtR4ncePBJZt8mDjEplEXtRgS540RV
rmPs00GGFD6agKrMU4CTkwlksZ6bqBC0Wu+poBuCgFHSrSgOXpud9SC29ZOjZ/9CCdgkNLiQRu+n
jPgLzWIEKLw414Qzn6fl/YTvJ7yXzON6NYixI8qpnxWvllDh1Ja51SpA4YQl7LtBE5HpKNR4t2Vp
ORwOMbl5g75xBIlEkmc5etp6ZAw6iA+cQUg3F8L7I5bRKTizkCmFn1tCEU4cvkRMhs4RfLzZyzAb
qOJ855wnPdVTDamFgKgElwBuWVCNonOnmqy5UbL0MXckUbVLB8yGNhHaK9kiLp7rIQIUxGzW3DgL
bfIMU2AU9Uy9XvvDR08IAkclsxVJm3xk8GKa2aMuIkA5x0cZWjqEWZc97GV1Kco8VBu2NgDRwITf
gTb5KUifVFWW8S0ttpi6ppukaAuDSOLLCd8qV8GJ8J2L0z5Ch1J1A3zWe4kzTn6Ee7fVPaZ6whBc
xs4JYllWxnfo/wElImIJKkltdx6cy05UCfjLqQAiXukWoxiYx7vHDn0qSLDlZ0rQ6I7ZFSy4MfFw
QUXiVaPWd72c/J+n8XIWMbP1GMDMCkigMpGUGqLYqnLB8UWouIMEC9WyT+cML2wGlImLOpu7VYRy
O36wApBGTM5B7xMXe0IEIpKeC4Mlk+3+OCYeZXLKMGFbhL/PKym2H09JDowVOXdyLaYJpfEEYRnG
/Dxvkl4tbc4F3txoWWcfotjy7JBGLlkj3QZ6+YU+YTcOC/FzL6DUHzGrC02Nk79pRmp8/lgYcZxS
gw/q6ZcSaurVfDreSfuReqnsIq/UwCA59hvLXbl5jGaCLR2kXgIgTYErX13QzQ+5GPOmHhh2RHYJ
6FO/UHfnZxM52KR1hsHK/fr1qIhRooAjs3XK/UT7EJn1KcqRrUVQOIn4G98yIJAAnVtS3cjVEVHN
iG4tDifyATZ+grIseez4Xu0O+Gz0GSpafXzdX86buasuXvrm1HtlR63V49EjMyFsRbhV6GAsBZQW
K3j4JbFRDTErvIXAjs/AFZMrOwd7FmTsnrtlhB2FsWBV7gVfHV9OSDVjXrH220JCNmjaq2AxDiy5
li7S0HRA03rQLfuDgzvEC02E/af4upUG4GQ0d5QwbTGZ6kp9n5RT61wlmHYT+vWhg4O+aLUJWBcR
D3dM5Mo6T91TpxzPKOYNkM5KLhg96AypC1WZIcTQMrc/UHi95TqynZsK0r5fjnKq48owV9I61Juy
MwhCajTAr9V7jIq+IKWkrT8223m6KBy1uUv11TVr7wIUdUlm7GO/H76UXW+vWvmbBqs1H2s0N4D2
7Ab10C1fteFKotWioYy2liMHyadG8Jj1MSNv5zZq07WPo0Az+CMzg5LhQftpxk6plw4uKQE/5ymZ
Ier76tKK78+jLO2kN+1Kretvvc7C0tEdYDoJMpYaLGAMpnHd5o07KO17pY9lN0nSRWbMofOMEK8c
zbaT9I6cRi1romKeiYW8P2ArZD4rgYTpeJWVLN0h09Bc5n9osbMbkwQnVarF8t9KXpKif/t4PPTk
pHab6rUWp3jkJr7XP9BQ70W0p5fvvAaN0UNHKIFo0f3QNqoH6gMiUiKupGEj4kbE/dppNBSOSdic
M6CP6yiYl9HDVY95BVKmOjXqx0187g+GnssNRPKHfpfo190ikd23nbPjJghBo2/68hIZqWaD6nAW
X5oYnU/R7kA7n/X6LG70jvDfOL/dswAtd68X1bxrv0TvkjQMVaC2wy1KHQCqnkizfU5/3rYDVGTZ
cvgqcgxGvZoRG6/O1TOYW2NxQLNFdUGAbSMBrdst1XMsPdRJ2c6yzQ4B2BlAARVOv1ZTOL2FTga+
bHS5c9ECbuHRee6y+Ki9rG3VzCwbSfLpA5g+OlXR8fLRLWSiUmPeavQDve3DbwwTx56fm8fm00Zv
UX89rpsPPWLzdQwszwMF1pmjhWBX0416XsyspALKvWSUUW0GTm8pSHPDirLAC0hiYFKYfXirIYzZ
HjSu2R5IK98P0yolMuzTo3s7vcWzSQJoH5yeWGIAObyjBh7fTwAG3fDlSb4RMPZllHKgUmoy6hvW
mCcA2MU3Ov4PCKjcC/+y2JuEJykyle9uO+PdzTE5TilXGXvwDOmyycUACphu56XE8+LlBAnRSNVJ
ghmbED1psSOoQuIF8fXxBIDmFdfDXZYdJ6+SH5c3Se/omT9uwGfdZkTh24UCNfSI4vz+B32ZKkHr
Vyapiuk3OyKyeeqxVkY9zj1HcUfBvnnVs905catYi1YTVAX6/WUlFYkdYbx6jZuoLNaU8iOm+IXF
F/eMsLwljS+x45GtnIzj3VhaM9B4Woy0daCPaJd+swsaiWnO4qw734nkRuFM+di9V2WoYCCvhxPM
Iv6MK4zLKLyNuoZmZqaYmW3uZWBwakdYc024sNuXG5QBb5cRxgU/imjgERyea506y9/sF9v57vac
v0F1UuvL4rfy5JA38oiTGX0vPfoO+m95NQqGYZlDJTCKFmloYPhwxDk0ncOgyhYVwWZaVYrZV80G
F2g0HwrJSZk4pwWDhuubhGXAlgVkVNiMXXwrFzjR5BInw0pNMUSJk4N0ahmtgs+790EtOM0ozTyv
wzcT7nN+AwAxhFZsToiyT3oGKsq79UsBmOOtN136YneC+8KqzKB8fJ9L6EnqqD8DHyWa2Q6OfYgY
dd5pMt5XGAA77j6MsgWNDUOMM9AC7IM+J+A6cP7Nv5UOJGJ0ZbhQNkiiNT10eAQg3rjzye18VPza
SShCuZSHBnfD6v7oAGFuOmz8KKYYv3dZbSuGXbmbEI4v0BoAbqDjFHLhFRhSXGppqU+A32Udfakm
z2kosD+jGZEW4hP0SFAyA/98XMCAyRGxraCIAfyR3n03JdHVZmIaFEDj8iV/VVIf1NWu1H0ML2Ej
njAXnR6TEC32KW59O6EsNd+U8OGS/nniLIzMFpdFTIixqnioDQs3ce3Uz8bVMdJOdYnJ6IgpVTSv
o1qkLb9tp48Zmw1Tsopljy16iWRudRHMvDN60tDSbncPuxElQjyjvfPp98/M6AWYcPRhCK/14anf
NU2khZZV3/xbD828HCwZeLD2NqarWxdB23UXdvt/YZtrDiPsbztaDhGv8OJaTXvzZ5He/t4kXals
BT/d54QXkjzHhpq9MktiGP3zmvMOeH5SSVFz48+2kk0yXwnpu0yGCNU3aPWpudQVXSiXOPvjzcFh
Kv4AtMbpNQt+r1+HXOvIqTWxAU06U9g3Rw+OfjsvIa0SLYuSGxpa8482S1ml4/nkAR9C+KNHqlrY
Wl1yGa8w3OP3dVSLvLHOPQBvPIehpwuze2MjJw2y7iQp66+k8g+Ep9v6JB/C9L2sTMOpV4BC1D8U
BPq4wLi4Wjm/S7cp2mSlwv5wn6Bf45iO3aO4G9qp3VWLYXzWCzPQ8n1lJW1CmmFUlzWT2OTC5G4q
DrawFWjCXkw5nw0anS95bNSKgWyotDDEoB8Pn3kXBANPbq3AhezgSoTw8RVY3q0mIiRUruMs04wT
wmYuVpOSjE+a3005u68uREq3khvca/O4xKqrMOkYbVBhlA4U5Va2L7FerMO2VyiisCMO8/VC4rLM
v99ZvXKZIdvrpp4T9DrJLB36JrqXNbYdldxjn9fM9wLVdVKGnYCBPo2a7rIoWyo69GiSz8B57x3D
Oqv20O4WdTIYNuorfNJ5mHJK+V6/ClWPA7jrihhfIbNYtUefMn7Iyk5UIVoI1M1Nunu9Dqf498SC
Tei8caGraXm7jN0nb/FXpzaVdMbuANvBu/Bg6T4cFYl0GrMBvvVyjMmTCJbIc8iyfr7TkhVcUOy6
qAiT2wZZd0lSuys2CWVepF1qqVhmv4v6J0/j6SMPYSgWEIbshHwRjkJ1WvKMOGXH/3u/lEYQhqvN
lREf8YBJ5tkuDpLtr768VOQmPWOv6MOzP8GRRgA/5rRrtoLXkvSe1oryKp98QEBg5cpkQHwlmAFd
Ca6n7fJ8tdqzR0jTfPY+jA33VvYLjIV40uWdMolFxQUhkDlAPVV6OeyPc4vB72sm4pFsGKtCQ7BL
ullRVo1Xa9jyWv6LbAjnXxsTUQ+sKdgKe5aaJ8Sc05duw/I0i9rxwIZ6HQ336NGuqugr7OyYIQeK
zhknJKU5LerATzxqS5CmZQE02SXc/1ESdEnuIFXLHeRz2L15EZnxuR0QZVbjip0iojf08jBCasNM
Pk+957nBsT6IJQpHDwVoYOskqa3Gt7px+IEn0tmspaz9j14Ia2cwGIyNCupoO9ZCmkk9CE4t6GYr
LTiBcd7OJ+GLtB9Y11N0Ho1mKRHd+3QMN5BoMaDZZg7/PwVR+b0N/+JfxhgteKXeyXYwCLOF2+a8
c8g6nex/9TM8zCbdf3kZTRWv2RaGNMaIx+kGgDLEVwu+DcwsIJrd3Ts2jJFROfVXCgAH//gFzMON
IyDop4Olpje9KDvfnwEXNMpd/xWax1cXGfHv7otSwi+oLcOMEsJUzQK/+A1RqYcal1WJV3qzayAk
rQHRgbm1Sh1PuT6ia11B7pynhA5Eh+/wWQTBX70xkLP6hZ3y9PT2sU0R9AwpAnWv48e71EvKUDJH
ib5MfqWqOzFh55ViVrI+izliYIgd000KD+16fNMO/pmqJs6QKrhU/rUpmmubMhgPj4K3z42UwvKh
Yvh3kjscqggkbooZL1ziahh6+9nM8pQ8EscqLNuOUsUnBFdibb6l7SS8CQRUaXby8qCX3Xdb8Egg
qcQJ+iWRMC/lCcoZ7pSN6DLhBxYEJpCW/akB4RpeE2bs9sRw1FjarbSSX6WlMSeAFFLYjsm9hd5F
JBeDl1CA/93w6YT1Jzfjh1PgR9JR6xYTh71Fl8al5bNlJ0KX6I1R5uFFXKsxhI/V7mZci6iUP3Ze
HbDjegxzrKeGpHlIENClzvBhrpahWVLjeY42q1pcO8CZIEKkdKXEEprfn66aVq3J1ldPCS91UyQ6
0NRxWzMoyoM4QBrltnhlNI9Ehu3TKxfmV7NnYWn2y+N9+ANY2dXnJtBo7eTXL4tghU2/NzMA0xXF
m40iL6WwFJnhdVlJwrEXgCa2xFCdirW0a7fJnMVeV2m74qQLzjzjWTm8RdIz/qY3lg6rUSOmLKw4
BB/vNMKzkNWguVnfIfHFZvnTZCkQOXjt0Q8V447cHd4mRVfwc+F6Im+6fLl8q96aKiN/zD+gGWEH
YYygapd05BJ7SnKEaR/jMiFfiVpffxRp3smPlCN6wbKCZ41GRi3ma/gVhWiggVADb5lONMvLBW76
dX3Tpf9F+gOdijBAL89vjO8ePMrE8izzU+0d2d/42kSxzuAb1GV+YGJ1yM+wkVhnn8nqrBRPPWzy
VvnYnSEGUrk/MzjpiDANV/pnd8Q8ZNBDhzMrbVzgvi0un85/wLYMGk23sMa0ZBJu2KidWOT21bs8
Fhrp9bWkKLiKtlVJEyFexr9+QiCEignJkIXiwu/YjqZ19FzSE1Wbeuf/Sk6fipXBPvyug1mxRgI7
U4AHM+ET81pxNjzzJ7rXx8PJuyd6eOdIn+YFo8qsP5EudWfUePAH/YCryQKQFShgh7F1xPJUcj3X
CwYGvMWrXhXtia7xZ2Pt8xa7g6I+LAEmv9+DRpUiCQ7Mvpumam3zAJ8v1WeqR38FqK4w1TBADmU7
xB3Mb4XSZVOQUtn2Bl7Qc+siTSOSmeTEGXqKEUbjNfFbngerFAg5MiyN/usmj+4L05rKbzpLnFgB
gnHf+isllS3CpBiELeBaBrXnxrc42TQTeMTtSw9NDaUm9mWhtGBqn5JaKX1TZTpJlRcO8MfJikrZ
RH5Y/KiFfKMODiHOb7q4MLYxoBaw3YrV9YtAby3hq1nVaJ+thuwMcmloteEMPsqczOyPavcoxxDM
j0X6xDyIj/Rqn1dyUILzoJ41dpdnGZe6t9Rfzpum3NcXsheakSgUlqfukTEw9pzxFA2kquQnO6im
hNQ7tmhCMU7/SNrpl+nzfG3/kWj22litDnoXg/C/GTb182m3bGpOOHn9T9+51/PvfszIi1uhlX+K
LQYfgS461HzXkbxf+J6Sq+uPuZj4DPJni+fieMKur0MmXKvB6su7X8IcMoNl2gZchVQfsMnwX5Gv
vAdlO5+XBLolRheQ2MYFIavRg7+iZ11gIy5uYdVp5tzBEDzaUomFVtexK+to+TX+t1+hvsLl0E1z
9Qm0vZ9+4WFC27c8XQZYZwUIY0yF+bjLOvU8EuEqRszpRaI7fRsA3q2IYL42X9epZ2DIgYcdeT3O
91aao9QKtxK99QsYwJ0L9eChwV2MqGQVscCSSlgl3zVc5gG1vSqPi8GHZNWSYF2uqxuReRCrlzHz
IgIFf62V7+1ZpoMQpspo9rLpyuQB4kG3NcjN7KXJcUBARWnQe+kEdzjRM+nXrpKBLYA5xQa36VIW
wHwVViZVPXO03k5T0dY2Xve8ze2mONycBPwmVVIKRyJVpwZborCVWsJM+9L0PIaws05NOJ/I8Rih
kpeh2cAjQ5LB9hbnM28WfiZkq5JCOV4XLeD60qFMv1xVIQjs3cVj4H9iQCQ4PRSVk6T5dRUAsyx7
NWS/npm7p4VCDJk+C/yCMwBSFC+EkscodZxt3z0gQfanKYsI3ktT9VyaSFLvHBePpCNhGE9TYr/q
mZZzzkneXN3Ewe5TdQ12uyStq1viA1ifM3s8j2RgczPxktB7PzrnTxpx31xjT5W15Lu2HxcVNMyt
Qy2/pasaYOZQEnGXLPnM1yplwWMD7HtrrcNDboHFt9xAA8GBi4bnNF2CZ25BbmKDX8gzDCNS+vMU
5M0mW46WFRWM1R7WQdLCbJ3sxX4YUG2hfCRKteVRo3CgHv2KktujdssfkRJTGs2//KPBZWahXreL
xE+z9atBJoxWybgeGzDPKbMcI2jcFOV77sxu+aKizzAd+vRPjA7H/Y5Okls3YWzdt1xnkIXbeSvQ
ILVcB41TR3AdaoccvfBnIXOMXaBnm9JeTuzE0Ay91cRtg7f2QxpjvnPwolEY8p3vMJLrFlNoRmzM
1G7822Unklt+oFEa4nnObn+R7sUI0ZL8DguGHBKmcv5SHh9HG5DKNVBeLfTuEClaNpH2FETQZCVQ
PADQ+ybLdAgPdUOq4brspEkK8yzTYMNzVwaOohYJ7VrQQ8cMIbYWhroFE0qOAYPjbBew6M/hlLBG
XJOSaZ+cqoi6VInh6558Odhu28R38a6ToV3W/RwNLu/gFTStwf0BBM0+oQ2DdxhIuTQJvpQSJIuK
y/l4+kDIVQvmoJDbwsRZYKk3mFw/ikyxmKQF1BjEpM3fWH8Or9ySzXOl4xuq7QEA7IsP2dz6uj8S
pH+KK4R9Ws8X1yDwzZMKfxZBng1QvCGRj1LHS4jeQ0yImKrFIRpsE7s4sbl7OhSd0AMNJSB6ehE9
gbLR62IdGu8iAYhn1Pq45xOp9L1/JVzd2ZQlSc9hlK7hes2gvpDrh3WqEiQ22CicJel+m+0yzi6J
/ur9o4ngCb5PPL+mj1vx2gAD29V48PiUIFiQjYglDlstNnEDAJBWusWHkIg8fNERbOitk4UjRScb
beQzdWYt5nmWR0vICmqaj6AXpEmE6rQi39+emwkncef3fzQJcbbWlM7MbgfDj5/f5PIXXKs6gPpQ
qAne1wrB1qy2ubdtsy5HC7lGDnW6/XAHogj5Zlc+EP4p/U/vDgvb5Z5ODOmwRSMX8SXOkqdvTHzq
oyilc1rt2TS0cdDEa0Xje0Bb6tWJnwayTPmfT4gOVNKFXaXrs4cAZ6b7QEzBBrcDvNOzyoRx7L7Y
lEt9ZIJTmm2dRnNPFvhzPWyEOKbvxToGdZIJiFQfE72+133/SpiAR4O9PkRsma3mBPLDMIkFW1AB
5O6kx/CKKOMTJF5gcGl4MGP5qXFtkTHEp++GwrhhgNPQaFvZSUK0ZesgN9LQxQU1avvBGzDtVRxP
P/W4QMXZ7lEqkTv4axQanBfqsvztJmy+zakRPuw6ncYHE/dF/xtqqpFEdbOVYaEPiTXK/38joJCk
879VsKRNO2tX6FaQH4VnvrNuY/9i5sYv/ElgCkCYjq+G0w6Wyz5bTtQ9jXI+yiNImkLxH4GufLFV
CCRpaWqfN9YipfRpEcmYi/ikFCx/nbjWDRXcFdx/F/ebE9G3lj6uJsj8l9o5lznRZIK0vFn6RoT5
T2rYkxCVPoQeospwNgTgz3206+6iQSQXn52Wh1yv9KDb/MZfBKmpVXmRYivB/oCYtPT90qUXKgtg
1RfTuJBDcULJZ5fnvWE3CWw4xXbIjcFe/GblHqcUTFL2fykq81QVN1zcUmC9tNoMnERlMiKlMZSV
vEE/oLAFJQNJdWgpB59ocCzFrnXJelLJCgi6GcE76e2S3oYuz489rZ5LD6TJRX+OhYkPBsv6B6VA
ExSh8kUWFew2opntYPtST8qICuMNOVM6ZgkdVwZw6lAvdfihpyjzO7O6Lx1S2AhPJg4clN/DP0Pi
F407JFtCr4VX47JzT5GkXxXpRane5TvfBTeEt5Bs1oeYVnhVezBRLnkRBLDXsm5wW82KqBKTxVB+
ktpY0OSNfR1iBWVJP1sEXUP2PldCcONb4Lk1163z16ITTf1f12XPRX0kSwoWFH/w5Mt37ZaJUEsk
St3z7iBRUt/DiqOUoFqKJuHNguhOqBa2CByYZUZeXpfepePsNVHGHNE5QHiIpY1YfVxe/aurYnwf
HzhQD8DIEbmnzTge4tE98o6YtZ1ZyVfPtAMiYDcE8MEVmEgGO1xNX+WwLTvGuLxcW3hf//arkdXA
m9MmCkxmPTDAG3cOseToBv55VcvvuC87omTOU6hpZjY/vA4uC0EYaKmvMFePXfPDB0VYiWloli9S
M3F5CWL8X5Rb27MFkcvWwwWxybCREyZbcIQCw8YL/B/8/hXZlMFClF2j7qRvtxTeliy1gwtyMMqP
0jQ/8adZ++4so8kkoJt0u72qQakyDVTpbY3Au5ZVDarYxBZvb9dGCvkTxGwaykmLHIOofGF1e7M0
pM0qQN25egCPOFnsx2tFssUWVECAiknQzBsXf+LqEzZIeDx96md41GhqLaf8ETwZlSA8E4lMYBlZ
MLAaRcg8IQvJZmBDS4rgwxOZ3ksnRuL6HO8MFLV73c6/DktTeC23YOT4Z2BBBp+kn8PNt/1xyYrn
3m3nFVgsAq4BxmZRO8eKTvKaED7XDGpCwxEBGOc+Uj5sO/CpnUSwl8SepshyKplLHvPO7XEhPjZG
v/NyisFfkUOYqzXn33dm46LOTlTnBK0LtDByTY/KJ/IoFpkSWmuB7bSAVY2RfCHa03wW4DeRMFWY
wMZpXzJA7Z6qcp525EnlPN37Uh+wkaVzftfJDvZP2Wc234MuZBKRyGVwcDjD0+Vo4H2PuY4xqQRR
XQMME/dTtn95BmFqvM9PoUnCWNasCeCWVg1s45y/VtGgddyAV67lcLga4r4Am6u99EU1ZOVYiWbo
lvkJIRzvjypWUYh3lgAZDiIDMF2TUMGrBXE/5hB7wlvKXd3subTehSZYZ2rlPYxupu8pfMz8ug7E
EU2B/ehcPIq3CyOrecKdmDdrzsQhz2s792jCOc7uEFrOGJQA3ggBpxtuu71vKRUK0nNLPdH3xUdW
ugsFkhx9qKROKM2MzXk9AtXZVmeiAn8Fz29JEMa4aXIED/5nvjGK2rJifxths+EVwLN5GhKxiWHb
KAcjKCm2/GqD0N42hkqWpcUN4HKZFH24kVF5CIMsY3Z9BlMjGzQmKgoDVwt0NnFTRCZ5qfEHgpiu
Ne1AV0KbGypeKPonJMBg2/jizdVBScDQbhkjmEllcUnns/TUlET+9mi0rF4youOuIYAOUX1aWziP
87fZLOBiydu7Gd7+e6xUcvZGMBs98oleKHfWEBV6k5xess6ROMTpEk4HNvz4wWDhaeNUchTYt38i
kXFqxjV4NXoix1cp+dxmk9DEpfSKs+XRaUI94gX0RD4MpvkoVHVN1VvpUdRhL52OmIMrxyYbYxK1
LdN3YYMmBerC0get4DQdtBidOzYzwrkzhaGzdTRcsDQ60tdWBN2Rp8uTbmFCjiYUyhCj/fXLCSZT
/06K0jdpHk2eDE12xw/C4ks2RipNcPmEeKf9LAFXAV7u80x4lDcZ3QCkt2LZzLuO6kpthtiM4EU0
uEUu4Q0b5K1yb3hq8cWi2Rs7UbV8hCAMDULHFeIUlMofnsamfThx0HcNKAthIIKLQConZ50PGGUp
PowYRwd0JjbgN/bA7SGeslaAfHfOqsXvjd49mUEhF09tHQPxPs7l2pGdfUAQeKYlbfyADGxn5EB1
hH59hQzVm+iN1pnYORdKLmF/L6Ijd/gJc95WN4PlsYBneSe/LjRK/GeHPj7mqwNwq18Lg7qQ5FEP
IPMHp4FmVZ77MJXmbYk21u3nXb9moIqXHh6zY0oHCMj50P10cU6iebDCMiyg1SQdiIMwOEmMSR9M
wswUbDVF7b5pYlhExNjYeZ7QLCmYX/uAcO8WN18ZlcOrkbd2UgzJzdZvM9d5BCyJfh2bNtNkAEbH
ZfvhQgYz94+oIwNgv5+jSNWm64/Z/dIAifIfjtR/ByIZNNkUnfFXGCisCp5AdwZj4Ywjyrk+mtgk
zJFu8mvSz7UOCnGFJD9/VM1yaXT6ezKT95u6nbAQTbT5syNQzq9JVY8y3ROtN7JsUoA2Xw4DfrU+
wnZuuiir9Zefccwir87hV+IWB1SloOCEeRPZKa94Y2ce3G3S/a11O1tdjt7JDqId4Sz0i8yXLiJ9
uG+zzm+jE8Vpie9s79vYoA9wPpEQOpmfSb4kCSEVH9NXpKCNe3yHUaNFvy7aiLPEsuocZLDhUlE2
2C2pfU4s3fGDbElwLyRK6t3OpG/kdVFFH+HyRBJauGu7lucFlc77vTaVNWs8M+BgmEg/MnT3Dh3t
MqtnGGBKyBadoYR25ykLDa2yRnqaNqhUtZh0NYYhmjvb6//fZbkEVNBkgrqDxgvircOnn8JlJPkp
9xUAun9Yy9gKjzajbSek8nDQvl12yvjfaMYRa2i/euJfVpV8S92I9uS/FayU2BCoCCAOoOATcI9+
i3vMNereeUH1CnO1X3GnzTyf93lasrN2IAImwuMSA2P/dMXuttp8/rwbgk8ZSORXY9Abxw1s7U0Y
/zTiXLPjzviWlB/UO5WVS5pJXXDaAkQjCKu5WElEpIafOrK/+NPp8KxJq/EsP9mDLKgnFzGilOf1
S9Ez3dvHtRQbr+cj04X73YAYi7d2fPt71tMJsDrBhOn1uDDweZwCT5UdvXjz2KAGxIly7E8O3s4N
gNb6x0Pmh0J/1VrxDuuTnj9sqOjZ3ncNlA1A/uKRoMMkRO7xqgGOUaABo0m3fZdDI17rBQ0LRMUY
fG3LNAGbG48BGXposxNKr+6RH39RqDljiVHOl2mfgXpLTnsyzh4UKHq28akkNpxQhyMbKR+i1Pbx
l91FdnWCGhZF6DHo+9y3WixB6v549x49N/vWSfes3q0Mcx8FicN95hnXFqilkWUvcQw0gBRzGTeA
dQgqCWG8pPGOgfVFo5zaHiXeFHdxsxNBIxj9EivfM9ugL2MIAq12SWHshQNVthCI9rWCBdmBm+FZ
5+h2+Ree4+vXjxT3XufzC7utInmCDlK9gRretbxn7WUFN7lKSZhpxZ2s+k6hookoFPP1lyp0z4/n
3amNY0TB8RRURD9y1c1MINt1iWBIZEKgeZghAnoQsO/PHS57ednJg960YjezArVS5E6XTc90jS4U
3KLIdrGOvgP2tt6fFBkjdBvBJnrp8IH+dyxu6roMWViGraAMPA8TrdTFHqJH1tCja61y3z+U3BuF
J+vEeT6umQU7ZCVYn1DBc0bCD4Gmre6YKrQJmVulpd6qDdi0neAYkcLVln/1XCbQMrR3JYoR/QWp
iHHFkXqGSyBQnzUqmR99qfZrD6Y2DnMFgvaSyDQfuuajCX1r6qdKy5T9MDktx0h+auYawefj9QId
JBOOFw14rJSixcpr9W8tubgrh+ZaACIbHyOv+hR93ycv5n1HXafuCfU9Y+A0GRqopFRFlpatc7Rh
iBUK37NsAvx6yHh4IvjwEG78X/b/diKkmFRg70GO4cR9k6oIycOaLjet/apqQUsGQswgDnRLJxua
UwfTT1NoeSRANafPixiPydvrxRGjcsNI3oalgaRTzWFZtJFyX9KnweEfa4iRHMZsMZJWB6X0VhEM
Rzvk0nzIMi0tkwbMokhiBr1qq3AuF7TAd2QvaU33T9EV9/hqQQbcYm+9XcalehnYpUP8Ptusak87
zyl0Plsxztc1CoHLCpe/nwPXVi08lTXv0sHKRX6f2HkS9lzCWcxQE7LBzFZbVMdG+t1haoSFx5oj
zEXrCeFXAhJaNai8STOtvJaILb8pIYp1MNjENmqJ0F1HkM0j+NgHkzwlg3mJ9iwGqU1KKnTVZngp
2HYmuQkT/7io7N1LxeM0X09wh36w2Ib3apyAPMvdBS4tojemFIKAldSP+IeB2ltW6YImODBuxtdZ
m1ucrMhbi/kxeDqz477r0MOQoX4giW525CkPyxl3NnbR53mHowB3fLTwn6ofAH2PvmL27sRsVwvU
hszQQut01GgOmwV4VFQb2bvLU1mCJ8cNQKd5UnQL3V7bCq3d4mE8GUWyrFTnV414UAVzf7DcdVlL
RriMZHI3PmytORp1C0K4XhBg3E8fdhgI0pqepwzhD+Ib7GQQkmIzDUo1v1/KoeoQRjhHvo/ArE/B
A8JkyglpOkuTNcMTjlgwYyHPyV3tZm4yyaxgdZhSTJ+l9JYqVi8rrAMxNfva+4VRyfa0VP0P1tMC
SXSkrFj50AAEBaFH2M3FeX6ZPMYRrPzOxL+KqzuQc9B18SCCxj20K8Mqz2YG7a062KvOlDjnFzrp
OZJNruuf3iBTUycWYzDi5HTckmHSKMJmFiyl2/cC0W1jbRv1IS2yVxS+0zXV4Dk+8ZDZ+550Cmf4
MsYGXVEbliTyRL57w7Vra4sQ4/fqcsjMY7HLW3wKl6lSmdzfOHSW6XFVEAXbab7cKZYImJh2RqTm
r89TksveE5z1IkXF2JSkhumjh0YzXw+25okmAPWCiyuGVs11HIJ9HUU9HasnqhotsI6C/cN5IbqT
T61gblWYUZJsZFG1ZuDb+Lri7372fNIvmp39JTzIYpO9G3KhntA00W1+M7cp2ezBt4m/M4XEOhe3
siApEotCIH31O0dNVeLlvmuSg29vpp7aD+Ucz8rHucBsjZgx5t3Iu9CNR36I1RHZGvEkSTHEcCPl
QKb9hj/ITlHzrF31RfBlBfAIfu/xxsdPpkCSvGK+qzlmMCGdAqz9K+BE767nHOrSVtlvKm7wvLZF
J03FtsTJTvwSeNWrU5RiZAvTkU6ZTyAkOFuOuUPIGtM+aax9p5tFVN3RQRoT018zZo07ikg/gRJ0
udNnfXU/Nq9iGJLtnP0Bcw2Q37rtTIXIuVuo6D6ptvMznFGJKUKh5L+6R1aNZwJo8U7k1TKlK8bL
YHBdzhfmBZ6X9VsyJbx+QB9lVyhr67xE4S6zSQhQ0zaZLQYIrXdRCfEJmPIvEE76EXvvuq0ui75r
jJeEP1D4sIHq2tVh739TJXaTqJD9npLnmWTUf9fj8B4uNqvMf76t220re1Syfebd7ypOHdo9+T06
kHVVshKm9oOUwjaas9GjxDTSSujHZp3oQiLTm6POmDx3WT+HhkBJiOMsqtdqMEecrwIRJt8/YVc0
COoU8JQdGugCNaXswjaM2HbXN9X6qRens/46k342VJT4KUPwDwlglBmMnL0i9+4Cy/hrp1qoXNYf
7TdgKkPPR9k0e+TmNF5NiIFRjevfaAcS/ID/7esSWI88eBCEV7lTiSE+hM/uFIn5V/irHDgE5WNz
KgyJ8NdvCgDrRmMo6LNwodFY944828mO6jreSwf3pDrHfThnqjLDA0L/pxNOl7lEpakA0b14eATE
v2S9vAIg0GuW85FT8dKcL69CJrGsapOkhc4FzAs4lZhpEXTrNO7k7KvoTGyBFhGD74QkxGrJo8lF
XOS6B7c+LHGcKenhUK+oJ4Ww7d272+KEBWWFxDDf61e+tRIVCpK9Lq5M4qhy9Yz1kA4gQTPajKNT
yAoQtGgOuWUz1FlOiXzquOqCQeF8Cg8utEs+ZE2sfcdqvJU7N3+E6SqLXUhv8+8D8xhXDiO1G90s
UnhybiJXVKC8LMpRl01YG6tFQRJ5B4NANUITZrPy3S9V2Zh11KZ2qyX1Y+OByNZLVY52h35P/84w
LouVpmkpviC4ulj/LyNCG2KXFbIT3s+INp7+Cq0eK1ZNA4070InYs/PvDzmnsqm16BCjLUyIH7bm
zCJ3oyN28Hht739TgEwQV2c9J4/i15EicDQ7FigDoS308uTp61umgMV4zK+hAn5dpOd8++0/O5UL
cHb0rc5NBtFmak14oVOtCiHCxwd56gnObuuMXZKh9R+iQStE+1RRxk2ItQ0o6MeK4OOCC7yvCkR5
6pGe6NPLTdyCnc6ICwBVRR83TfLcU0sacOyolAhLdVsfwH0eV9R6slZI1Kcwah2Kv9aQb8szeBnX
TZicFl6iNMoCB0b01ItfQp3HoQd/wm+nZeefIYWki5xJyoor9wA9u043gb0WpiAcdzAiCBPgt7vZ
0T9m2qBhWVC5xKkPoOn4z9DI3TGkn9WRCBhg9vQa0O7py6tPtMQayNEchXihdEvGJbCokQKa7RBs
I5FuJmaAI7VMD8SguO32svo7mlzNMhr1LcgTLx5RpmnhtWDoMZWSIF6AOsy1TdcD+C0Fm1uehSEc
SX4PM6kK5ntUo+5bXS2m2k524eUUz8Va8TFn1dTG5zfXfeDlMJwDCObgoVr9tBNeV6kHJPDqnPvX
/sVuyWYIXVeLky17UAzWJQjtfa5JUb726j6GUjSUi+EBsMdbzE1WobyzpjuSXGKKFpEJpaBN17eZ
tjFaDbkKLEhS7Nwv4cRqQmkKzZxNOsGAVkWjjBfLFXSP70PujWp+xp3Gh7lwO0XpHbRG/LPzLX6b
TeTMOU35NMJiRX/Ybdb0DjNmgWk8YXO7qed6F9+u458OC25fbfBe8VlXlWkHGxZWcui6U4AuBVeg
frGQbyxg9KonX58aBUzYV4XbWVaJHozykIXsI9LwtrhdKFH5wWnrRJwytLNmvQxSJpzhThVMNSeZ
SpmpAnrlB9AeRjjXyMHPi4O7tefxfYgaFss5sAr+T7j88Ed99Ovf2b3ihe3Y7TTeF/BV8VSGOCP7
s/oUWsEBy2xJmWIl5hzMPsXc6nqvm7THe8pqMfSv6zCgYKIrHhxaDVzqarSVhBPeHqLWUJA82JCZ
k+RGz4cEbBoeJmmuEjlCwLovlYGQGXavbKnPZHeFWxz52J6ruOy8fxDmCZ6hamhlnOl+VDS8X9m4
fl/8+wthWoHfF4ely7ppltn4lM+ZqQYx3ZMRyHmOtOkwmFyrkDziSZpC2sg+AonhsZxSmfx9M9D2
lEXtWF56bdMPJmlvu0HNrSQb3SJazXAkJRiTK583j4HguxNY2IEF9r5QmvwbgHrTQYRAFpaLhoa9
f/2Ps51WLEbkB5BC6HyVAP6SnYD8NkiVA5Th+KGsjni6P7AygspzUxukVeaRNXCtgovlcR6U4qPj
wjb1LhSGPbHFue+IejGXoUgAbur1yFdsJZUSI4qOHbV7RjGAtdUHp7LFIw+rpzeizJMJJpiGCYgp
1HDxVLo69nQU6k2GudMN8kPoCkTmXimrSGDdUBZygJVf7ZS8fDtN/05XSHrR6DVaSkqmtSNIbiNC
N+nrN+9yw3gXMrpPuaLsDGRq2p3zL4hK6rMjLBTat0yJHGTGgtuBO1vYMUNEl9U9e4JpUncM/U8L
Qxgvq7GUc2eIawAdV5Us0rntGfhiepxns+M3LDNWn+A8hnbqAVky454EZAVQteGVHb4rvmibd1dh
qvxvjuRJlJyDN+NOX2cXamD/Z/LEqcjxPuogI9Iqz1L0MY0FCVcr4Mz602tO4xD1pzG6uoqK/xEO
3CGk04cR7nUOX6IXRHVYsB8Y6P3ZG8czk9gGf3rep7bi4/V/qcaZCkt6nD++aWOhBot6Q64YzndK
zSnKf4wr7Ony/R9jWQl8annU1y5v9x64nW7uz6H7cuprunrKNdT/lHX8Jqbcv+XOYczizYH+mOBx
a/XaCqbIn0LA4I3Ym1y230mACgIwOlWPSh8ftzpa9zmxCKKQo4e7UCSasgwjBvyYRzsHAX0iMVHu
iM9NfMEaFL34Vh0NjDH9ERZjnj12taL1VGQ1WIhPaa1sbZMhkGzGpPNsx530g5oRZ2AiC/K1dT58
Ee7aVWgacpVj0sgOgzGDZwbpp4+gbm+hdKZhD0O4+RwqdnOboi2PnYQjdrVDoOm3eriazMJYTYy3
LBEaViRH+gYHyLWqJPxH6A23fvzz0n1O6LcTD6WqZZM14od3aiZLyCHnhfjJu9gPM7PgErUY8IWZ
i7RhJB0pDKZo7teT1nV0dbZft7gevxpavhfyFhVDmwEdW6eO5n0biL5kMI4DI0GEDmen2cy3aZxn
9hveUxkqwhx8fz/ML8uYkSjq9WBmUK49J8RMNbfX0RBoX2jWuug6CXX5/P13siyiE04AHqiPUL+f
jjHgFgpHlx4JJ120JZ0IZsfi9xBqtCdovWX6tyB4ztBnFxNXQSUlDfUiMsFrulvoGESQECWZ06jl
QrYeFR3TY0gB5RgOMEeDW5mahWfgjhNUAS/Ryhd0zFXDq8JxdIlkUS/lXVWHCw/u+KdNElwHJTjt
wYVkZhguYBWUP4Q0/7SxlKA4VsS9zCc07d+k5AS8+p6yaYBBqXb5gWQQj367NotZNyJZPxbJEgJ6
aVgbybvtll5mtaxM5b+zmHCQdBZDgji9Ltl47ySuY5TKUAYiWwSmeQaHdtMashM+njr17hU5dlw6
nuskKY/eIVoRaFLhbAEIy7mz3ltgkDhlsp14A9gfSfAvMDGpezgp2HYZShSgsEkBUW2giVZRSNVp
Nggww+Iu+HQNHyzB79pTuJ3rC379F5neIo+gmWQPUnUUtuKFk6EdxhWWfViktV94T6tVe88kPF3d
UkzPITUrNnAMv2p16bDIyy0zgIXA6TC/pGt2gcaYBISLsBG1N+MVrlS1oQUNh/ddhcLW90ghz72r
Df/Q5sn7nW9Tr8NRlhgvxX/bzPAKVRXdPPNbVafQ79KWd/0AyuNlCViTUnHqMkkAC4tVSFHOJBG7
WvphySldrF+G01pmF1FAhfqRP+FnLhNBQZQXFCC1MjGv3G3gQ72q+debTkr6Hs8qOISwChICg2+S
Ins8DfBk1FN1KX+MuukcplJ+vCn1dfXrrjHRfwojNdn3tXg++KcddhedzMCoQfpc1KyY57dCEI7K
i4Lyla1eOC7mtc4KQ7/6pmZg1srmbpXbyZlZuio+a4PpvF3e3CM6ADmdmvoPxGizLJXnQTxsFrQ8
zL+nu27CzaXVSVmTeogZJliM2BBXpqZhz4/TEP8w16J82ksJMgRPMvvYGGAFzMBGqrTouyYKXD5x
o8F8o6C69JaSggO5JQ5O4CpwujEHFlNhpQ0PhOyUKToflqeSTiOrAiDk0E268NVQ1vtHCcTtEduE
5sizaYaL134QXDNf1HlDg0fWw8z0m4exRWdk7/B7Rw4ZLN2rBv9ymVlBfz+IDHiQYnXLwPNbWBcA
YChI+CXVVTMDwv2UXrJPmk5Y87j1NlBxoytVCBsjQjT8IXiY31foTmwv1m+uzFRvfhFrAzxetuv4
0aqNDkEdJCEDa0kIVVkXAMYp3djAfHzVTKxvdf5dkJplfGc8nwsxV2Zu9TgPTe29bWyC+hPExdfG
jU5xv7Yqdk/0v1D1uw6q7oe6Ei9YgczG0MK0hKmYnQlxLfC1PAhmEpQcF48dPlwalawu18DwcM4P
sR7alVwEyQx8eGNdMJE/10WhjXRH70q6k+h5IguGhy4ypU5JgptQm1ngRqNFbJ2OpMuMfg6XQpIG
yLZ6to0x30SNExuvbPqwA7ycBjd5rR+4y843Y5L9GOkJqm6/l6HpBB8pGzk5XMwLjsDV3yeHJ4Ur
H4bf+v5BzwqJF2B8dbZf55XXJ+MRa1Vcki6rDFOxhV4oZ6kDkiIeaYqx0babE3C60HDTggaerCmg
LeKTffdTy3MDoSMacLSvZVYVoZ2iToTL2yHqIDkC+6C9HEfm5LbJUcm83aNU8BC9zj6FHyRI3kJL
xjnx2LnDajIL6godPQ+Xy2KOh2mNagZ9HT7lzWGsUV/arqKHePdt1PJCBLviCpSPboH0ehkoHTpm
DdAQdlGkzc/GeAM+NzScQ/1ari0xxye0eWpQG8KIIDvlzSAJ4WZGrF9wzCQiWVVLN4DtbfZv4H4a
cwUqgokOSaos77h4otAL+iHCU1YuV7p1qOcwnKob3P2spzgRbs3SCzuY7KrHSZPhx5iVcKp8XZIW
t5rOAuX9JoSHerIQP05NsUQbmIv3VPbujgoxLv7beGSpzxAY/TdFjAaBSTqGDWHczhMJISSvFCqi
KlDaejKK0Waw1FRhxKLtiedSaGymmLsl36/mD7z46Z/aAHnPYCsnvozaZ4bgLN4pda09Y5k0qgAZ
SCnK/Th/qSR0RenP88/l9KzEBowzvU6c6mTXb51bHRvjaQJnQO+SXUPysANMb8YIy9BaEMJ4ZjD9
tcFrWJBhUEqeyIrKcU1Pxr+lBPtAgXMNvWvjnKSpDBm8674DTF5otrqBdeHw6aRUU7JFtd5VaDff
A0CFvJsHG0A0OzJeMvMHv9dU4xmRnJFrk2usqKJVP/H2oAMAR+vERj6gMXD06ZijEx5++a4PDoZT
7eMtUmAZU08TGMC8WONmyQqrB0bkUU5UV6kar+9i/66/yc7X15duYNGzHqmAbzlZ7bfFVwM62e6U
UrtqCfQ2YNc/g1lLQ8S7w9XMRaJ+iuVIlle+NvYT6P71IEaleWOfEkZ6qEn1Uik2Ch6Ygh3kX/Gb
zZUuu9LwIjFbybd12oFZT/IsFdkLeHgNsZxgaoKu9lKbNF5Jt9M2ImKk9OA6iEsHfCH/1yLB47KG
f9da9nMuZfb9kLNnXx0enc2XhYC2RtlOSQtY8eM6/b4FMF3u07b+7t+yriXmYMS/xxgLGsqlikq+
OvftpksHagOhFG7VU5o4HiVnFrdQMyqS+SaPdFhci+BTwBvOzdkdmuz0PTPYEo2316J+hUqX2oDG
/7LTw3GcUPAsB0gOsfY52O4VfMQts6MmyY494qQtmW+z4ZYHo8ioeQbYjxvGquFfzmXzFynOrKX5
YGiJD1wkU+9DANjh1TerkfmHHbF7+JaGBJIaFYymgnO6fGsixAvY8PrQfT4UYN1SSulfoer96+R6
swwF2eUwmAjNSSb1vlOtHup4kpG970nIOHlDX6In7L4bJkZQWpedy3D4AfNiWqB3IHdPafICtPAx
hPnsDzpPnaRJ7rmI+Pdltya92j8t3oonVAjJfZ7SDBD1Puvkr0MgviSLMZTUl2xD4b3q+2tcad+a
kymxTteNx5267ZKSCJxTQ56qS18rOY84KUlN/8mp7Fux7qLziYKAMsRdolG2t/4bAePaijwxHAHT
k+7B2pKyR4zewSjvgMyvmtkSC6hWprpAlqk+unuHMZnNgfhI6h3rozkNZodf9cpVsgRhGaX+X8VW
HOTtqcuwbQ6QqdNL/p4OQgkdfSIEUS77G4uyPIlz3LIsw/GjHDwZUSk/UGcvKvMWuEOGONJX0q6b
HTF7qQF0982weVOQmDFebS5KPY7qpl2if0+pnyGNgQypGa2hCRWGdsE9sOw0UOLebtpudkk7MnmY
/T1fAsl//NU4ROoJ4FmpbNfbV0psyVZTNySrS1SIYkeLc4W360rfmJx7XCS5pXMmqrfNLmmMYHc3
aVQOgDT7qQl/uieexQg8AbBuQtK0WSjjlhwie6M2uFR3K+NVvZVnYnnHN7R1A2LXv1KV073/mr/Q
LRFMwCUAmCfT9lSaaLI9IBhsbGzXD6TpZeKVusYSPlfyWkLynzi19G8sH0cUVmr8+5IDJkooKSRX
Dsc9bH75ZyvHa4nANIMpWIRG3+Vm5qNFK3yd8AHQbjHKXtuVfTRoOUwkjF2xFXce/1N+SOKnPnmF
o9CSjwGdyTfymdb2dl/6MawJnZzx9gVb9rSTyZz7tqUjIfg+pdMHWPhmanmxeHSVcrbUlXYo/WJE
ACUiYHonIeKx6TlgQZeisvLKm/LWPuJMRYKuY2kwjnNsOwojC+kK8wNSUpswonP/N/6f6JOHZi0/
gBBEkxVLQsuwm1WqKscvtCG3sxD8y1Pz78yHTLcEbvt8ncUqoAHtXwwBVGzAvhCAVSuP3AliLT/y
ueV4BMyL5VOHrdzi8FLp3iYMHk0yS9Ppmx8WkMhGpILwOhEWCuYkumBHnmzIzZA+QsjH2v3bE7fy
qCeZ7uTnaU6Uc0SJGWye/Nj8C2B6QixjH99BYQqE/FMtr7Z2+0LypGjKGvarcivjitZ552mCajO5
+0fO7Jziz+dwoflav+dtni6Ah8azW1ltm7ocVApsNx7dxKvO/ewltS55uWZz7ZuPukYe4X6ZWoa+
CLth1DqamBgY+s/1RL+WkaSS7TTdUQDg0f/E+2YzduOtnNaB8Ow3GtU31fbqGlL1ACG6g+Jl/ges
bHKiLT2KHRqelLeBbly9xoMmfZGg9UpFcXYLQcvEqciCc5e6cP5V5OinVrLuBlnChjRD0PiKaPdh
KQHqyMgqh3A6e6wHctoCfgqJach+d+dxWcfwQhan9tQHozEMWqAakJOABc8FZ14mD1k/XXdplqtc
lmLuk2vElAPTKVbeimXZ2mbrm8Lm6BR5q6fi5ShmYYGoFwDC1FlrpHR0JNgb2d0SSZ2tDV1wUxZO
TFReYy8p+SgfLujMqQC+9G2069P3oFNpEtSYpujMQ5UMs5IuZSu66ZjJQek2iIKVTHzJozMXlZlx
9uTJWVeJFqi2A2YX67D3SeJfcy4JJEXO0hTYyxJGTw4q9zwVP4/NTt2tG08Tw5GDOo2rW4jIn+9P
eyxuB2gjgDJJ2MCmGYspe6Xw/W+nf08gT8vEx8kucULzT+HAlfqwg4pJaVHX8CPQOba+P4N5c1/5
8vqwHPYPatqfjori0Huv44Q02W7eigu9df2D6ryXzA4LCdAWQFH+uMPwufW/e3LqfYa0L1EAcSpG
l+MPC+aLsLKqwA0hjmmepLHK3uhXR2gYZqlybuAXojlRf59tJ/qZ6ST1gAJwtoQv5geHvHtd5sIh
xLusIDbOKqxXX/czyaWaQwfSfDxCtGUYYn5H+azsMDUNe6t3qirqLI0ei8bC/xD8NDzphnslOaVU
BoJmYQ8oi3jOTGjPKxtf6AHsKiM41Qmyd2P/U+bgA21/f2cqxG/jLhJt+JuxTpeLM4VDj1z3wjAe
L7PSywRM4flL8c8Sv9pxxxdUKRClG2tIWu6B1Y4QXUQ5Op7V37kLrmmTOQDG0MavBIWaUJEyfE++
cuGkZM9r3uyRK/p/1k45/lNiLjSUX0ogEfuw4IGnY8RKRbDzMcdavdEecMxkF2hXCS3BZSMJWIgv
i8nt3Sps/wJr4rlFYjfZ3vpdzNr256kxSz+Z700BPzmKylmVmRG8iB0yRhtVWp14dmq2+miAjdvc
KXil0s5znu/PrLDcR27K8KVWgmlq0y161HtYfhKLiYDLXx3eXK8HMd7EUbaC9HJFv0s4HApczIqH
BKgMpqOnpPNOTQ40TsB9vwLGlrGukyrXWqSdLZFlYNZhHNKqTTEdLo0scirDNAMCgpUhPQigC7iP
1j8+mL9/nGGOpFDubbi2lz2Z//tcfrpyyxovsWoD/XWZokS+B6pq1BKIzWVKXYlSDGRkwhI24JzT
+Lg4rdLMQ5epFL8sAAV5fXXV4dx6peEDhCVOz5bsnDlvgt5joKpPFu2WlWsnw+Wpm5RHoqK4wvtN
MiDduilU4BbQhL1SbdwQTvY5xRSXOB77eFRDeA+yHaYr93T0uDvpJyf0j66wjXqZm/INsPJ1T+m1
WyRNywc7lZpcGWrXwD6gUcBfBlLC8KWg9mdygOVAKotzWW1SOuJiBoGrhFzBl6TQewV/SVrij51n
n+BYjz/T1zHJw/nFvSXsMduNwh0xXTIoOgij3tFqjU8frLix+2o8Gd4uvG1UMs+vu0s3kjgzGvYu
n2z/j0rrnBEJ/ofuEHjS2f9B7qGGMpFsMf2pesyRk0pGiwAhBBVDrJ4QzcuM01elY87ngkah5rJ1
wJYB+LIMyGGYPRdIznWoTrhaAD7h0mXTXcxG4dasNrlrYIXPBboT/BVtYRQbv53YZuTDagXRU/Hc
OWU2kOiQHgVdMxgxvthjZ4nh03XJiydcTL6CX6Pj5zwfepFI+TPklrpj5ECutu+B+/cSVNmF0yv+
gBGZ5oyCfSXzBhfEAWMHgiiZn8dLoORIqneq2RcvjntyfF3yVCsB/bD2hmsMbDxUTsp+SZcmWEEG
IBZmk23cNxdf14ddzrIKldbnGfhIoxUookYlFc7eC/XdKEZkpfi8/zEdnHnCgUqINqn1/DKHe6Kc
ugtrZlGG7gCrfaCh8BqvoIWKLvrCLnuMzt9tkVXN7QsZKUgq/QG+ide8cXzB9gfRfHCFAtaFOxmv
oBTLj7YE8KIW4jYQXQ9VTXmEnONNYf/lozGfRt/qDdAt4193yUImR5LltuiMn9h1lIDdAMUbhYpK
dqhTv9/pjFfNS3qUg1pQaPqz7EbVbcYB8SsyRJNdfYVAOta9390G4Uxe4h1vTrl9MkX4EOnF4b5U
SV9YN8BafEEahulWArCSFf0VAKOuD1Kw6QldaKVtSKbF40DR3OKfFLjbGd1jyAYkXWhj2NqM19af
MMRdtngvsNqyrY8H1xVDfcMM9rs06ImusOehJzeE+gq62bcPtPug2mnMo1GGWUGZaD/O4N9Xhu6g
JqI/xzR9EIonp3xeBdwoRBMBfMmjTW3CZPhqhVlpFLutGq30WV8rHpTRsbSiw1QpaBOzxoqXR7oI
E3AimkPCKgRWZYhvK1FCG6U0hWdsqHRRWhSRUTHP4Gkf9uVG9CX8gPOv1DEynMZlCiAwwvCxegC8
9jwCTvHdsEagIA4Pxj5OeoYqtDVlvKMEfMiStfHwIaxYaJQlhRuWNcJBhVlhPkPyr1JgKTDUpLcK
7JO/m9J4w3DJJhCHScSpkL3bELSkbaFP4cjPOrNH25YVKfSX01bwK9a/cF02qJAgo4VbS+kHC8SP
+yWal4Apl/J8/WzTyzbo/ac84nZxMBrkeZRM5tkjZ+/MRVV/xBE42Cjks1MFXNIOarvq9FIvbF7L
fuAB/vxezgZ0hlOUD/X+nUL+KdLJU7Il+41aEYQCW/mRQUl9quorGFfqhwM9rsm23uuDiujpFfdy
K6IBTVAfJcVuOWGDxMJ9aOF4gvJijWy+bioD84T4jHXOEbDOe00kDI/LtGZe2D5/pCWkdxY5LX1L
0G7313fUvxxWZOxyxKZRu8jzIcIwLvcQoDl3+kIwk9O10O8dm+ePMCunmA1Wuu1nFLrulFI4ez8R
5ksY/loBDH/03g1ecP9i/AXpTZmF1FuuijAGIkuhdIzxEmOxmkHDjvzV8iwLOvh+5eSr19BrbwrZ
GEBN+0q4R3cqLQnR8yEC/S+YQZT8h+CnkvZkKCm2/rUb8rQrL4U8DzqjhKd+rpXp1NnqzTIvy46B
0rOCAhFoouTx0tswfgKp9uiB9t7/fLTFk2vGyyv7awLJZPDOplxJ++c2AV4GizTS+abTR6EAaw1w
m2hXyGJrml97IxAGOFHdCSCDWLsRSkyzPUxjhCnDkWbdfyPzM2SmHWEi8Q2oXetPY25DnBXzWWCD
q+4ahTpLUytLoAX0v45IAX1O+3h0SLIVzM3JigmXEPqlsJgWjGro6WF+nAhK1yMijo0KUE19N4iI
Uvf7JQ7x0As8GpFhq7YDjtwMoGss6R1IP3t6YB11CrRP0pzymEJhpcEqRqqLo+E4pmTg1ZO8yjGV
12kFFwD3DzjZtMfFDBb+oSmc+Ob7U7crTxpMigFtUIu9f0sKrpgNlHw/QlMe8xNqdY3He2L8qcl+
whhR+vOKuAhk0/VZEzloDyD2z0612WlU559aL4KGhIb8radaGeU1FpYTFQObdFCRdZR2MKyc2byd
Q6JrmpFMZRETdYgQZ9Ij6vdrXOZ7R7RbReIxpNBBHQaEeqSZngrkMlNPsvP0UMn640je72EWHuPZ
NhRVEhzCGEs8tvwRHjbcot1SgmERwYWRQvWq78g6JtCFZdY/ZM6+a9l8q7v0UQObGfNP7AbofmVU
JLA+4L9HnOngBb4mdDsGGKiT87tzzKpsEPyScNGjj8A0l1kpY0vhgDX/Fuh6eAGQO0CLusw7CEHB
zk3+swnJIXJfq53CkkS0nnKeThO2MX41b2VKSlkXXPZe8QIF6h2Dr+rPk0jCg8wzzHOMwBNu8ijH
gfe2ByH6Hn7R3UuyaAz4VYDVJuL24/pOzvF4EZgST+vGYX9d/Iq1XDEuXt9BB9LzSNuhmYdmN2uS
gFXoxZTXIX2sqvTHI1FBjXzZ2r4rtyy7DP/pa3OzZviyIxkTTTcRX/MzdAO9PM7z1GxyPaX/Z5dB
aEUhsJOjfe1rFCJlfRftJQ0MAt5j6PQVJWBTRIQV50DxEmIcyNvgMIZgARpuClpnAW32HWe9yLMK
CCOwXMVEQNKzZ7ggcB5BTfcrXqiPv+BGayUDpB20lwiMG7zkPa5xAEHvDURm5y2mIlm8VKsgkJVo
pL/b7P4SuSdvFvvbcDm8gvrv+Gzs63YbBhn1HoIEDS+bVOCpkZwlPIqMZ+3k67WAsgwTJx4g4sVn
Rh7Gb2jNONLXDhBGoZKkr3tvTQulzvjJKZLycVcPmkh4Dl1cEGbXuIi8nXV7AuoyQExJuAXfXK7C
xNDFXEHaIyOQmeJgEseXAjY1zB3DhOD1bdFOZiaCbqv4nNeVCXJvNhsR7xgbfzg7ucZdDbGp3e/U
YX6qaw3Ibu+h58irUO6cBP7tCfXttoIQFRWUTehVzAteHUOJKF0M+Tc2vUTkF1kImE12VfuCAZkX
wTzI8nRpNsXi4wqxdNncIrlxUx6dXQ5gYED+lsPSiFNzFLB3ve+1qQZ3JPwIZw50tLN2YViJcBFZ
rvdFrOOA8/wWVpUHoMs3FwS7vCVeZ7ouy8NaZHwwBxFP0TbQAMyJLxoLb8XpxyeBGBTZ76J1LWT9
dri1ecxWqW5rQNWzETAO7T6BDgcD4gP2y4d0Sv3TPDsuEZ+Rrvi46h/+okoaLxa68DWG+5KJDzIz
wjnHXX5ukOptR1IE3X+alLPsfG+ADEooCgOBw4bo7jOxlDyI+gCjDabIPFY25rzsd5Xh6DyfajX0
bBDqJeD+2kMGqMzJ3uNp2LTXpxtSD2nhljN/FXQki2gYgjvi4fg5vp3mwvMCRKQGd95LBdVLFJkn
U7T/J1I1owkK7yL1nyh5BEBjIcPvyk8wbGu+4hRsznTE6RlDm2rV8cJz27mqAriUZhF7MJxMulTJ
x1W8g+t8HeLmAJ7GHGRsiqvQSX9xzrhTej6B/O43d2KwSgqITkWXWpHdqFk4SkHnFuGsID2npsCt
ISENsbo4k2FnIFSglEOD4dLJ5Bj/ORJi07V8iffRPJNNZ2XnRlJaVGXCbLLpGMGtyndVCZtLInl3
PQOpNZ2nmGZkcnFWyfl13rpaGgWHub7+MJ1JX7pgrUC5L99Gk8ApGNdWiMf2Wpx5Ot0qMHmwvodN
G59Z2A290IMHdoKJ/SjUZPTyqmFbAXEDfJyRKqoozIbMXqaWDiLTY5sQXc3yZ4W9iPawPFKn95nK
oNrlh3N7PUwQNAhx3bgALWHvAs+bwEOoMB0FX222Fad9PAVL78JJTAz9UNk5ZRqA7yM+Gyg40UIa
IpH7PraV7WMYkWhEZq0lpnBBBvtf7aJYCVH9P52uv/ZqyHiC2RxvNDlpKXKAR1ASkc+YBwXWg2PM
QZptM31EwP95/a/EJ/az0ERQs/lTV3kT1bAAg7QnFSiZ5RR2HGFNStFypyFDsnPmQXSUpYqF+VyI
Doal+E9ljOPXvS6hmm+jaLRIGBR/2nsUerBUsAaNdMH0LhhPrV54Hpf2WeizCh161RYJKtzqrdeE
A2WaCeJv/o7C/Aai8t1g5YkiJKJfmjZp6e/oZSBCyzHNwDgUmZNuKj/PBmCq3f3Do8khYtyEx6Pq
+uHK9auV5F3EDOfNMcmHz4khHIGsqX9f90U+McXeNWy7hZcy+bfmzS1SbVsTBzPUrHibArQJMqOW
6zBhxoY4W/bHg518iRlA7+QmL+DIjDY5kXAg7IF5Mv5CEx1oATl4tgvCAz85VVqQXeuIAPGGouhp
3d+5AQ1mCIlR+AB5p7cign+g2cvqzYNgmjf1dplqbKAHjjB3Y1hNv0yVwB1IulJvTN738w04qyTF
w6cjx3ICUCmI5qnf22HkdiKgAadw+7r2apPOJ9wyF2fPAQ0gRvY68aVoUNqOD7zztw34BKvHqXkA
D82OJMpP6MOdcB56mqFtFGtbBdvYtmoYXUxCT5tbJnJd9yCEdjfctYBj0MLb49pw0miZXqxlOYaw
LnVvSpg5tioMs/fXsNzz/58tAU4N7E/HtTWNyb8/1MkxyKKkBz550IOguRm2Hpmg85DGk5rsPMOH
H5cdhR6uTyKHV3JQpWzq6mFCc/4ycox01gmKzX+fffUeFMxI57B/BFLurloGweSEgqzuswOKwDsK
7fNgPD+hGPxNuEFD7gqP9Dw4s0UaoL+a0JhQ2H/qr6+f7SCgjy433Ei7DjcUy/6CwRYLXEUnumto
1grWHVD+PFDnxNDNiLTXLgwsGj7KzOVwTRtS1mugNPCYNgVMEyLuOQm1dTI9a2S0Wmpm0MUz1skX
EowcZfVmbB3MZotH3J6FarbxH423tXxxC26mNfAthNTSUhrhJsDS/Qq0s4+zAsekwFocevVndxmh
V1q2q1x25JBYo38JeWpArtyVFIUZkIM3rJTKfmPLc+F26kEsz9E878QEBuKD9pWIEeie/kD0mL84
uWNgw8gJ6qPxNyBRqao/BzTxGHsF82nJv5pokLqFIP47lXvJ1GxRvywJ1aFqe4rzzjH1wyP0c4px
HyV1cjm0fGiSPB83W0YLYHbrTxceTSMqQS67aoqLnMQ6HOSMwSfT5evas+oiQeY9gdGl50rBS/9M
9ZwXQclbHLqc6wevRJSK+5kamiGBFmW8LKvXUkfAJLVKnRSkaixwqACC9rkJoyzxTa/rx38ud7ys
94cXVrA/rCsObsxm3aU3H9nlUnH4n+LP9NU4bnDvNE49gfmhwXdjZ0aSF/W3CL5GIqcmbZ9DhcGq
5vLR6O/zUUjV06urXwc0G12yQB/TpItigFmnV+25uldEMfn1U/G3d6smOi2oSEF0PxQNXCZSYxEJ
eMZEs/FzeXf46dKNwfnxzmOVRxzcdjv6rR1wueOJTOK1Rxhh6EzYICwuFBlZ6gpGHafqE9bRQ8aZ
Emz1ahByPlnFCiUdTvoR+fulwI4QXxdWIMg1TNmsZAcvjYrukfMPq7ye/MWfhSu3pckRMqvfJ4qY
0AycKSnkoQGMt3yX4W1AfzRPHAuTHDZaCM0uZc1MpSsPXgwyy45sL282Kg0sSV+kd1jPkbVNFAV4
Hyb8VadADYSlXK6SN1jpIOPYusMJ+nn/W8f5tWA3wDgV/kXv1lxhEFOpUwx79Rvjgry+L+qIixrI
dxVW151yFxmtErsrzTSdpsgwrtig3vs8azkoWeGRyCy0POc6d0SQxwBeqR0lf12BUsb8b8ENivHn
jUww4okRB/S5/L4PP9CV3RJaPXb6E3d5wwDmh1SMzxaTHw993Usr3tujdPNT85bCPaVcvSWLyvq+
D20Inavu6VjImwOh4/Z+Vwt4DZ0WyjBSLDVNmnIr88ZR6WqK4eC+v5rI0O76O1eohjtIlQRvOkn6
pLBHisvgSNicpMpolw9blThW9m5CU+SQ8RfW8SyK9T3ZTmiByki7yWRpOA2Fogtvc065zq1cHDjx
OEhB1e3zaUnw6drAIPFlcaCotjCBzeIjwimoqlAJG0lYQvVHgBRl04ovv/07fJra/ZqpLTCiIxTF
APHttv36wfcqUcAk8lCIYSpwVMmUJklQv2SC4MAVz31TZCPHmpNSenljYGSTOuM+jVDbSzgDylk4
iYY239ULFnMpcsBBJvFVndBSL2Zc3w+0Yx1T08II8FNLEwYw6I7c/igmqV0+r0qR+uvDEjCiknge
3+hgNgWtykK8PnGrHx9LmmHaHNC++uhNs0cStxQpWy7q1zw76ZH4qyOmSVmlQvLH4bY117tVnYt2
ELeL03f+4bBBEXFZfILE/WDkdJRGRngzntuivVSrvdVs5KgY8UM1XfjkT6eD0654QOf7RSKo2e2t
a19Uh8m2whghakIMX4nt5jUZAl/x7K2/99XRGhbZk9bA5BAhcLX1M5urDh1KV5iCqapgn6xkB1bd
bs7+LUd8rVUHJXeL80+G3nCJdmCqfDI5fOF3WJ18CIyHZn+UJtgjcqegDbTh6AXzHYn6FTfkf9jT
vibpzO6taaDD+UBP/tDe713pSw4fdIg2ORo03RSr8qmAyChuVc8D0GPD67R5GSBOb175qPs5reUj
Q0FdGHePJaroGE5OwoXzgScwZQBrm8kXZx7/bWwnx4GFluIxlWVFdU4hzugLNwVHzde6cdzlXute
i+E5xKDvxxUmY/gBCtcxxyj/SjfqMbLD0zryvsZxIQDfsqqwReqw6L7ABqsNQzhqSayzjbHxpdFo
LnKUPNCa26+ROLxOn0Es2U7mTaC76AJ9ItcKxQm7ki9rMzeZaVw+JmQI5dM7z9UwgQgC0juO28fA
kjKGOSa+y9Y7XmXlmqA1/yBI9RuuqgL6YXBquhce1QYKryNqIGJGx/htKTMVyyfg5hU8/0B3Y58r
WIQZFaaq4ezEN2g9uHMqkibWhO3hpoZ9mh9gugww8wBaaUdTcchwCTSwBiLgRO0IOj9bgIFv6xPG
5CtvwdZQwYYXU0qMtzI/oePt8MngtcIM6S4cx9Fc5eZIxe+3qBNE04VCnoX/Wk7JHRkRwRnA32Ee
UemlZm1AG7ZPGSaO8sYSFsSlyNjypSgdmghid/RAyOQkpX8aSin++OBg1A7pDXYGnzFFYhdRJhmP
5p3HMMsEqIL7mHPOJT1QFIHgPs/lPBOP2PC+5/zchK0ST6HkbmuxOMbfaKCMcJSBOyXUGXOp+P15
8zJwDR00pwkbqrJg6XxLo9tWk73XzlVk6gAe4rJ1DyC4O90hnme/ypAIV9QYVTg9naDtRpS2omOW
NelhOLcKf54WihJUT1CxbmYrjX1LrByw/QD/Zu7yesHN4t8qhqWMIt57g1upnnOoPdIU+YftJ86F
sis23QB9IGQe0n2Z90ryTT0JOmf7bmJfrqcakI8GrDVGfTA/MXU6ikxOqDZTPCwQ0y9DXvlvnhN0
IQZNYDNAkqSMpmMIXajSgGbLM/s6YHBghObHv3LFqL0E7fN76a7T9aciFpMs13vEbOQoKlp/3fXg
WsJI09WhgbB6Gz2MJYSVO+DULJ57X3D+0OTHHX9xJEgf4ROPP+Gxr7i8hu+S7f2pYlp7A2ECbBmk
bLFdL/3PqlSj7Sx7NeuY1eqf/3hbzOayCbxPmuahLf/l47CrlllTgXmOJjz21xAtQjvGMeiM0mmb
3A+/az//qVuTWzdubZJ3wKMDEZPHyItnKqN33A0cicdwxr1dOg3mALjQNHHW9Zpf3nINx8VDcGPM
+9DYIU8XLrPT81lgoShlOc+NymOWWFmGBe1u9kLobg6LeruKncTFczAAxUntLrmmlnFy3Xf+hJhE
L+d44vocF4vySr2XHNJvizZ5vDoYRnm8ugP4eO7kPRel/6jsO2zpRy6Jokd0QYORWjD8b7wMTqjy
e8aHBvnlmH+hReGCu2UXr5Pcuy0ERgC9tZsRl54m0gooD5A8QhkwyVSVacu7uOYDiEn+/BMyMHCO
NLvscmn+kRsIx2PgGp2ne5R9g4XHE171UEU5OUU7ATvrAk01RqCEGOxoxqFCbFM6eDExhLnAlkh6
zHSd7B38CN5iP+czmbVTARKcOczBBfVvNtc2EE7f9aI+RJA/9PJv1KUOdDzDlGGCKK/MC/Pekm2K
OjFoYGFBApIGo92cX1TO5XnSENdBV6B1HwmkN70/vWQsnMd3e15y0irwC9pFioXGJ0CyY5bArNTq
xR1lUabaD1DwJvcOw0W5OxijXB7r3nKQWCG9GbflIkPkl4rzrZuxgxxIzO8T/7pb8zDei0emuSR/
KWAQ+n/BI1Z2hkm46amhqlEvaBC8N+RB4swaaOvR0rBSZ/Dtq7ZEEdiZPehdLaOM037a4nhX6iJQ
AvtK2MngWiDEKFepkNGIOUt2joYq0d/8YCTOjhJzdsSa7Xxye1i31dSbR9I01bYT5LiKoHk4Wrj+
uBwqVNQ9wu/+gJzjsvisdYD8mB5Kgq8m8fPiEQicgpubM1CoEm8aMuq49Hj3j6Dwgu+hYjTSDdH2
tm47x8xnVtrNLn6Big75+ewRm1HoZX2ibJKmEzii4fQNyB2xMrO6OLNw0p3WZvPxRMPzOiSE3rWC
Sw2WkMgD3OEcvYmLbkYYncZYVGKchP6cHnetqWeCQXPd5z+4RhWjQA3xqe15zQcJtzBln6NIPD6W
cIiOJlSClnR7J1NA4BOIaX01NClUGarIXWpyyinN2mrpkfW+4cuoZ5aABKiJuW0tcESkWI5E4diy
wem+SrbQiBmmZTnsZ8YNr67VkWi0cE1RnPnufKh3ym4Jg2gdyTrfunKruVRuzVTNjYIKFO9207kS
YmSMauDkJIlaOf3wJrcAfqpHCV/POQlxPazxBf+Cl7n6W0lKDTfeBKz9KZxJYjNteMq78plnnWnl
XYrXRCa20DLeU/CsaASKbaNLYKSsE3E1m/55oW1NMNVBN18liNVtaEQVWSF79W5JTJPZGYI7gKrH
cLd0zUepwyUbvxlP+XUJR6MFBpCubDEZMZl7kz0zMAfJcFsiYZKa2kQTnz4uDAJFE3GXRRQMg01S
qalBOhNQPDj0tiAMt7hDecFcOGGm7JBEiWoLg0/P36LbjBK4JfCmQm2out0E4NWGV+WajPUBoVo/
6xIuZxVvA9SKt9XUrDLFu+SMn3+3ROBPusLsYnDOywex7/e1Pa1FEgS2kZdzhS7CtSeE9E/dGsM1
nu/xhz0Lma0V0laA7Zj5Y86VRWSN7ZNA7780R2+BvcTGvdoKg1BlmOz/My+EKnnD6SsIOQZvIGpC
7Q7EsB6G+vfSAdJkswyz2w2QqHpFML9SadmEDfbOSbagJwgZrjaOP3eatx1DJsEZZkkVpCW1EuCB
MUMhcYXCQ3J14lM+RgXDdNpN/PblPMGNUB1MnlX5cm1Lblw4xeEsYhdwUnXfUxh6c/a436NMgEqt
TO/7Zy9n1CLBmC+3W8+dc547IMjd566E0+FP2KUwa0TYAq66+mFDqU/Nk1uhtp7joXBAnu4zaHd+
F4j5AkRXpWG8ddZNd3RqkzgFtushogvWI2oxqgtb9IlR9x9MnEfhbIPn94gtWlc4WTFzUIQlffZi
dClmSoJqQRvLFjJg0BtQC7WopEf3BJTqmBQvy/uxkNVQ0SVDt8jDRE6tdbcAQSOlT0M80bGVWIhD
mz8oVOEkk9nlfWKyoggERrgiZcUT7zXbD2xt9v58NJ/tgda/9xUyeRlqm3pqvC2B3VMYQtMf+sac
SAsAW4ZseoX1cUpOeGaw4/uOVMq8T6U61aBQBXOGyxjb5IuHftF3teX5jvS5OdXxoOD1JqTRbwF5
1bM2VWzcEjBUbnWjIf/KH0wT2CAcapA3nD8TxP8Xg50LG+uhmruBa2NDoVG7Rp2CAzMcD/iaoyIl
h1pJejj3y0uJOFZJYpo3k7oH3A1VILZgcpaSk2+GL0VUfjOEOiYSz7+zbjKyFVBb2m4xb8tnvw9A
D4KgZr04s5nUGMlhuiUkm2DuycdMqOW6gT1djv9NcujEgjOeNs0/+fCiSZFVCdqbhb5byZ9RB8W3
lfI4UOucJA5BHKnBAAq++nScy1YfEMaayTgY1oRFsg3LsziVkIDz/bWwIsyZtN4+3t/pr2YxTgYT
h9RREwbwgRaHUeiTlpXXXlElYAGHqpjgnDOD0nukNkMwdEpmJ4ridmQPCu9JWf18UPkY1TColmPF
4mzv7VExVsV9l3Sb4IHX65Vn/wKcnDOKta/dOlLFaVFak05YjnwurhZVx4QXUMC4Satjkru55WdK
MxOz61gPH+LgokguPI8JMpIM9BoZPNLiAPWcCLmFv4xR0XNKwMeMGD/p5soz/rWOM4a8rRVn+1wF
ZvqdNnyCm0pLrptWf2Tn8upguXs5N8W/uav3lvyi+yQ1/r3wEBUpV94J/yqsQFmfQWxzyERPsGQE
V/mf9mDwjs98OXIbHOQk7t72D4pqD5CpQ6wAzS9NUO/fTjjp/m5KA5tyrYpVXs1UEcpYMwL4g7t2
GZlRem6AcPIhy4j2ZMfPhBRg2Ms8snUx0fXdofjm75CQMqsIe+L09XOdn6U8qGUv1r2SNWCLhIKS
9nHdKjtmj4UvxeoU+e1ya+Hh5g1RSgkwp3UOLvZIyZe8Jlu3g2cfK+HnT51uIpLjB6VdDX4aWkld
JzkRjHD2WXVcTX/sbWUN5kAWFZlk8OmCMsyVl2diRdJEJrvohFoelyUNvRVH5Vjx7s5ErpmhGhDJ
Kt2WXpAI+7bRkKNSOPgAGxToF6eafIlirl0eqzO5/o+3TkG8ShzBSCzICFoCJ6CGrVRycYBIfN6k
ezAAYRJuG4kK7RQtNfBdIX4leAUMvhZXEpnfIQx7kJQDhrcjtzookfe5t6XJLoVb6Rpa1CPOTbtm
CETTD9xtf6oMYI91m1ssJfrBVbSIwIxG+LrMb/L9P9A+mEyyvuV3yfyIGoR44sktPxYzcGmYUUnN
+ueq7Hc+7BRXCxNL4dnu7O93qH1tHmDkUtZq5arQ4oZIigc9lgIpcFeBmOZxCa12kataqUbuIoqz
zm164ch7x1o/Vj32XNs4sg3l4FNYxe+0CI8oBE0H1VnYBN72WaXKJk9by2vHER6cOPTTvDh/2+Zx
CbkHeprf6nHfLPjWcjSYzbvAnJDUPIIAyABVXbFwFpw65jCX32v4Jn7A6VqNX7GuWuqIFB6YtpuU
fHL7llhKaQv4nYgSs0F9aGfO6tlsjk0a0zWGkYUqFi9Pp3bbqydGhb5+ZzB/YFgGvSk7yPoF5boN
+P3geV7LCZuXmoo8yulDrGxjmEGPBVGfitntntDRehT6OX42/8BWg7DJzo/RBrqpU9GoQ9DezrK5
DzqMDHtr3IR3IbNNWEqoPCivgzdOZSzV7Jhkl/RAGafF2jg73ol1MZmcBdyW85TE/j/nHHU/Gmp7
+fivbMNNBrYk1z4LjafBm2cbCn6marQRHBWPQZTFxUlb6gr30frsrQdJbfJZlQsLcogJU4OCqWaN
9duD6bB8WP9gmMrF9IfhB9yulb26/hkPb8TocirVd7wGnpQjkEg48y77NRRokdMIfJwe+AyFQtWG
ETR+KHrNgQyLrKIhZZhBj49oKLpM24mBPz+ggjSbtgEdOFglvUI1qlrobLqJWT/XyY1pkUi8mGo2
ycKGIZnSyG4kZ3me3eddk9S8OIyUaYf1gzJEUqkywdF/RhWipAkZ9yxKZAAd7H3XQOU4H5M2bAxA
4Dd8cHtfL/s8eck9l69YFl105XM/+EVK4JAm2I+1epZwzzGRRFNY8pvws/RbjPXJeqFgiG2X6adl
bPEE2ItgPz1kbSJku0SiuN+rhUl/1S2mCKYyCSdibhb4wvIZyoLPjJy8mwt18WrLtyHvKsJWecju
xMzuLfyidcZD/keyC/buiVw0GymV+IcPNmNAI44Z7i2PtKzt96tD5LsqtaD4Gb+KgFXNvzM53sJq
ZJFzGlmpq7ycg223JSQQ7eIq07K9ZvPUxsLhnl/QjZqdYecoGYJANtKSUpofB3/inDmQlCi3KTMX
fulGZmyBKKYn4JMqbJXOCHLGW+PlSrwPol5mBZx9OT2xaVQUaSWewDFlsryYgzttaj/daWu5Bus0
WEbr17+O6Jv+CCYwDZe7lxV6jROxHKwGfxGGcFApqK3G30G857PtBCPiNpb7JONm5P95BtDHUDW4
G3fiTYLQiNUQ4XACA9jNRVpSI9/Pub5+g8XApilyWNfqKDDTvumnMoR62KVDWUvO2R/gpCCaSkd2
YMtNl93RmG4KbuVcmU59OoYoqpgnkBIIX3sgI7cpOhgUb8z9tfb5NavweE0cm1N826TzI4yxljOB
85oicMShQ/EEyX2kcElGIh5cZoGQhC6rwnpND66jkS2M0xa3ZR6soF4MA79CncLTF+XjNF3FixPo
5lwTEPq6IqXyr3juriy0Ck8xyRxx3NowKIa4LXu09fhclOoLYA9bMm/5QFTBcGjSo8HRqO2/J1oE
RVve7n9GjpU/hOcU9xH9/NkRwApZwG/+XbPowPD4HZ8e06yxNYKDnX3shmM+jIByIzPTua7wwMPh
6GhhVXeTdspIMJ9z+bRcffZYg5UIZXYYE6QHvYkuBuQneTfbj4JQI6zUW13SkFipAC+ZuJ93cNqG
86MoqvwAzEWYqjTmWiWU9nItbaxNsa4Dx9vHled6ZIRdjR7Lj/dy/ATbUydOBmm2sQdWewbZqhWt
ie71d1deTD5EruujyLfm43Kg6UGE8tGMRyT3zVIU95H4spxrJB36vhuLlk7oWwluq87gAcV0HE3+
VYc748o4s5QNKL5uF9+RgS6YilcsFMLXF/5AnImQP/GFyHkq3yq1Zdka6JDKOH9CM4jV3UOXdfnc
YFHH0Jc76AKg2BCeqOzWZtDDkGmDvkynvFigQ8gN/8uHJFqpHhwXJQqc52dUZchl9N0aKy80DD1Q
6LvU6kPG3tFBDs+vLoczoAsVcSZq8t9i1qWKiuz1cTWI8+O545LxPKV3UO8wnd3wfKRPloJ+YEwe
ZuxF5gyWE2VNqo7LcsOISNeN+qt4fAtSMXQ5DZiveU0d6wiOEMbstzKAj2dgKzArM7KF+pViQoEt
MztujByhwoBGII3OaFWllxgIDJzISvmaDnL8vh1L1Z7scMFCNSqljHFtZ7kiCpeRRfqHmzxu1biv
xvUXMYp2iuiQt8ebx3D+1HbMGbWGJTDhHymayHKJ4QIDSqJOYyUUdc8VRoVTIoe3qmLq66HLKn33
VoV2Nu/HqcSj8ztlkqjysfvq5XS0FRnZnkGgUAZO41PK3rRFI13ExzkNqglmEF6YrkAAYnuuS/H1
aoYPK4+rvpwWRgjFAq3MH6vUzs5+eaAEr+rNnegE/NKeXBx7c9BCCwAEh9Q4gKPkWV5zuF7N+z8L
uSdjy8K510+gVOKtQ+na+0JX8GmXJLoDFQ8dg6YuxGgkrAgeWVpDrraYQBoZr+qf1G5tKoFr8P5F
gBnWcaFPf/6Oa8toKWbjzataM6I7ryuWHN4MCgUOnN3U5laY+he2VgCFk5RszFO9VK+cRPkG8zI4
NDHHf+d/n7RE4tuHa2d8sC42iFYlVRQqG++wiEjb4CyKNHF9YqAGlz08laC66cK2WklGQPsZ54Kf
7eV95WaplwO+9dUf/6T8ns1fHbg4S6WEZte4i5WYZYt/xia0F8HrqsUkoJD8RJIjeh89Ogxv13JF
HyEUzXAX2Nw/2PkMnhnBwtDS4eaHZeXyl8wikmKykJ/V5PGMMHjOnOILTzlwPTh/2i5x0Uk7118F
9prMzH1cD4hf55idUovJ2Sx5PJEmkUfHQqHEBY/WASsrJGdTiQDr9cydj2PyVPoFj2y3kQaMGtC6
Ds6DDO+ZnesOiTxdzUdTXAnqlOYASUuyd2KKfNBVbcA6l/js4AnUCVKvfJID11M8vpigtiVRFZg3
qz+9RlHUWxfTudOnwOb9jJr+AxVsCvnWqIdDNZzcDm7E9142gT6bVwOgTs7aNKNx+kNuJZEubwPK
MVOnOsNXbIAj72Yk/EclzOb7U3Yr02vtaISRZDDBgi3KsMo/vVbznmMutR12JSfrsa7mjPZr0nrw
m4Y9hcEgdnARQU1dqjtROHtMOoOeAPIgiqDIxavq2CVwdhpdqL0Plzvihw5XJfA9cnNnkJAFvegL
pNC7jiYOD7l05N2+eVOhpwlVYXs6kyzSScVIWrj839u/srpilQ/3YT2Xz52UKUiQZbjPSadbzZrd
LVL9hcIgVj1vsOyxCKXW1FM8TB3zSJTDgJiZe/q9CZS33aijopeXtBUu+WBerK2tQNJByM5PooXK
OmhhKISBi/dxX8yCHSNgqbAg5er85mIa7Au5r6BlrdR1iiWY1wjbJ3p3hddrfWHZK6F48Ej205hM
rFzko/wpg4qlh2WJg67siu4jzfQqMqAT2bz6SLZ2X1B27A8dl3zCWkg/Gg5pGaxo3GOKH2ydSOeL
jnLulfE8Ao9Ovu33Ps5yi53p+Bu9R/RGPCm93c9P/lIvGXF/hQg6rRtwLB5EyQAX5oqtGInRXCjr
0sZhf+lvQy2K211VRaqtRn17o8RMfRgGOiNvOUjDuzwtl5BKeC9ak8BUKzBl07I1rd6DDJARuo+g
qIZkA2EEPtkrnc53GdO8aDCkAUMrfpA1inrVeSHA/jiC4L2HCrxack/70xrZMZ53zRI2cytJV8KE
Run7aER8CcgBH5jSvmekWuI2Jt2D0ngPzXXiJnTze57DdlygZm2sfSqyzEGtMjhTjv8BlgS1I4Td
oM4kdecfj0zDfRZK06pLQ7BlHI7cDhcbQYO0Vv6xhBqJAnM/UzVfSOyksrj8TMkx0FOKzYwO9mL6
0UjDKSv9Wua7s1H60Le7/k7uJvH8EVK/rCvavMTr/LXuR0IB09gJ0Tk5LvPz7XSqAnfVois/o2dM
rDs/4BJwzBXsz+OHzHJTUhD5LcSk4YxqWxgnKxfzHqubwjz+uCCGNCTtC7PEH7iZmNxG5QVWx2Pd
bX68sx7Q8iVXHipLKFi3CTiI3lvPbUjXImlcyFpYX572dT0EMWYTz5m/SAEToJBZVfsvQc0JFntV
7lb4zruKhbJootLUHdcVx1ikVuTr7izXbtxgLng+ZoH3Qu31IH4HGxsp1veOxO2y4SlfQrl3+Un/
Ld64mrdr7sTEaZQtOK1lfyhvQt6NFBDxYYcENwRNncuSuBfLbqqXqH86IQ4H2jU/A7hd0HAPpVzK
E7tyfn/tunyAyv6Z15MvSO7xuJ+qszLm+BituaebGobrgJPF8/PtvAeNJMwYmjP+REwfnGBQLEwb
W+8FslTYJKmP6aodRwGZabMqW0mzkjdwnKxKLH1KRai/1D30o05RY1lns4bXjgPLxlZMyBL88raV
8xN0tRk3/f/jtg80umpsLBz43Hi4v81DLSlH60mDRjJpKf7O2gbkbNnHYDG7VZ+FXGDPOaK5jTRo
iktY3W+hgw4WR4fVHeZRjd6A+GvkNmY9ckyh96hf6YuuoZy5PX/MCtoPRv78xZZu4vz5paf281HU
+086KbeL11MATJ+PPpJWOiXAlA437VaRgmnyKCjOGXfcndiM3x1UHk2GS9aA2jJ+Tdkxyb7uFwF4
NgueYpPeS2ZCP1B8HXfWnhePm/8r0Xmbz3Y9IifryuoTxmJpLljEXaaDEGBQmTYu/vRiPoEf4c6+
bmq7kbr7K2DOC3kQPkh/0e1fWT5+CnqpSPTuMyAm5jppDID/V/b3CsrU6htfRHT3QbvnS2vqmzPi
1rMPYKATZkdezBrSYmyau1I4QPBlHbGKdrIBlqlKgQYLl/er6lu+QJ+eob5jxqLjQydYkE8HC6UY
AjQBwiBtQ5rQC6Fl+ziid0kKG0bzJM33RbkVmYiA1+Bl5y1aEvRLLaixeJif1LAa1vN0l3AeNLBc
2HuW2lxMhGlqKti7hBK4w0pHY3YrQUbFrUdwoRns8uCgXhvXqezmjUXIpapypO523NSdqiMa1+Nb
I+BG81RxGQuhMpBAgfx6E462cDX/6g0mhgtPEmX/QerfnjRtITMo+pd5lqir/pQkLdVsuS0LN9Bg
Fqz8kMZEjXEPfegQYsnMvOk4c/T5XBEFV0+GCmUc9rdkwKKQChsTAdYwstQBVWpKV8Gn22ibKTl0
jUPHQXKSx3JQgUziuwjpk+qTF1Aa02ggoZVE9gYW5GVJ/BKQ7C18Ng6PeZwIvR+GGQQcyHh7MqBa
WdWJfgzju8hue8py1mVHfx6c9gQqvpr2L6hbdGGp6gZadld5JbU4r1EHYdqpNEko7UmU5VFApys2
WBYdCZtGjzNIX4GPRPpL9oVUtV4P49yhO29HX5fdX+7J+iFQpDmsScomC6K+MBDzATr7IISHdl4q
3OKyoHsQVAWCEDvUGhQkm0KPGuGoiCzTGTpye0itvcE1l0oYD82ANC706B0dKGG3mfQQpi3yvA0Z
ZXQGi7JXULrpZpJfHoeBSVk0Swn4eM9xCvPneXRuslnOO8KeTW9QH4DRUhJxzppykf1PgjL5B70U
xpauuUtyaQ4CcNxvfEnDNs3DM5xtogQP4g05S3DAKVjktDQNLLmtVJV3SIF9sc5IjQ623PcLuKVb
6R2YdoQOJiBtsP6YLtKZuVaSvFaczI6A/bAquXm10gmAG2yFdmvI0rDc+mPtM3tniJOfKfB/l3vN
ynR9kQIrx3ZXJqJANHbkJhhMluIR/w33LufLn1yeGQA5kAsU6fbV6aIJsikNGG0/vIp8haIYO+lW
s/a46yhLWWMWtKvHLjn+RNP9LU1MG6qmRhw71GdGWmn9j/zuHDCi+VfMEIfXdOh50uZKDrvTP/FJ
rFIyETy5C1zo2rMhJdyB3My6RctaCYYoAPmBqz99/AECJcg6fWQRy4OyaElYvs1sFV+kGqB1Vp8p
yHi82iaLPZoEUwsKrDU5pQcAEdcXVukKPX32p/Kr9zJF4fUIXmKwBs7S8gyM/+mqnExnOyFwixl0
rLX00n/uSRtpbBQaMdQDbokWiqTtSrDcG1oOwvpd4OzB6vhUBt0gdS/YOjVIJ3LIX1EAOikdwPGo
BBaFPWYjo6MaGjkereDO1D103Pa0RE1EjNjxvpWqHRscZWn8d3aF71Lk4JC3Q/bdP7xmn4iqVED6
FdWh4tMLmMWsanIss9PP8IsI335klYjfWEm9+SwoqeBrKTFOPf/HyC798l6iyH2zdzk7T3XWqUe5
B2S3nuxoStAMK3NAwQEqUkv+lt7zIatXV/IMfWhEur4gLTVRx1P+GbleYiqncwdMQt6t/2SeJVj/
9xDU6iyIswXBrHqVPmYr3sHyW6Q7SwvCuxLFSIDTTcK4DxYN+7W9DOTWTIBbACjNRyIgrB/hwWKe
A1Mtv7lSOhMkrIz6lVyp+HLixJE1rT+bTzQBJuv1icu+wumEohgEb8dXyaUvluhS2SFjY1NLk6qp
H68IAcC2I07v1BEv9w3voQ/ZRCWCQG/dVPMbutNekwHZt3h8ZyZriQWoM4ElbVlBswatKaWJqyoI
K8CqAzBJvWHgPXzQgYw8dJ/n6oqbPLgo6fiHKJu1mUr6vzowXZVx2lbd4Jo33db5AIA7V6kHjR6O
YQurjvrgRRJk6zgcOWDeKomNFuCRKXmJUO9Hm9iwP2akHTynu25ho9z2iFVQxh8dncFW+nlEAoan
zux4V9Qed1xOELyR7mV9O6WTs/wZWal5v5UcCOdXUbN2nIpk3PmNQpa7j6UalC+IUVr+OFLOhteI
LCl2J7K4MlbHNzqtwXytczNFTQ0KixHf5pNnN+L9wlT1AWLsVWS4D8XeV7Q90i6dA/G8tqzoub3k
XU6G3o1+C9Esc1BLqmUrQQnNSrrD/SIks4DnxcqXD5Nk2UuXcANm4un01xoxeAAbFcoxyuHtsbT7
Qhk6ahQsmm1pbPNkV9YTOEFdfyHtw8AAP4xD/7zrQtDpZp73xmnnXCVSnjVE52I3LMpdep//806x
IZE1bE5x1w7u9udp73pHG3hcNNjWX4bhBdiFQj0b74X3raF7sFesI1M6EiOjgTlHREsmL5kKJDgC
A8KuYm79OEUG+Lbnx+iTeriTdVjPIXjYhIYgyR2hwQK7o6LfqJLYKzT0qfOiZQxXwSMMMqRfEeJE
lNe7lbgpoxDqNDMB0I7CvGmBkX2UFNWuRaUEYam7nGLbQMTEZ1uR5BQobglUahNzYoOoq+pQj+w2
jtuzxWsaDF/0DurjkyoOeHY81a7QBjw20jEZcvlm1CwOcWK5fwBfYMlTq3+K7j/dNhZQ0nWEDtdS
Iw5hHwyNO1FCJodtJgNc4NFhIJQBIEfMd//rAx3HkQ6DUOFgF5SmMoLQ6pu+QmfOL899zVayDWuR
0ogdtwJXGCyLFH1V7SgBJVPHEdIgw6I94q2IPRw/M6/hjP6HV7966acY8jGbLjYnwNuLFpDxR8oR
RjxM1zdTrQz8BO8ovTNTCWkBOa67zqypxTL31ydFv9LNT0rGY86uQ2hk9fy8/I4ILhiThJC7iS9K
aW4tLBjN2d9IaIsSZ+w4HcLsQUzK0fDKSWAOWFuulHWkknz9XpJzcBh7YlhYHqsvjXdQpq2Vwo/R
uZSBYt6K+zXtGZMOFautVh+R0HCj3UDOhOnegG0fX10D3XE8hcN5vu3s6ldPfv1KDl9kRxsdiIz2
xSu99xbeYFzmz6WAjdRi1XMxFAzP+MnQ172dcFtzTu+RNLtOJBUFGF26dd60OKZ7QP4dOAteTQ8W
QNACP6qnQy3PvWgGKxIFr+wZam/BeiZIRB9vgLpSmhlk66rmQNeTy3QvNH1NNX0kQ8zjFneRZYiE
vy9UsnitKFp0aGldj06pM1sd+OXvFkqOixCb9PiL9HLrWnXj2b4SA9MniT1udHySTCYqXkBnt/zG
k3mRqtFU/9sXWQpYM9GCyaVKtggyHyf1sc6AHUFvwTQd2PaWqJliyFIWlvBjptF9R7U00OAsZ7GG
htV90P5bAHp2Y+sVxg1xhGy4aebfvOZaOOhYnBMbO0HG+0Am5l+50MkAggLrc5mlZh52a8qKbxAM
UrW6lGqgkTsVkXu/8SnP8odGfwMzfKDhy542TvNWyR/wZzi3vGj7/asrz6NCqu8L4x8OTVCKm5KQ
1dxYRDzExbrA1khjC2iTJ18cvNU6ghvbBkJqL6cI1GJNvf3v+gTRhSJmTIKryVCE8XTJeKIkNhlW
acylTAblRBtdNdvSnUm1ByTEVZ6zVy8FPlNivJOPl6258dz75u8F55Wgjp64JKN6VZq8v1yU1r8L
HRifTtA+yM25vmI4Xx7j8q0LDyCRoVIcaEkEcEl0FjFze0iF/d/iHieAW2k0QYW9bVZDOzX4oUwL
032xrrUmH4XcdOX6y5vBnFFhmJNpOfyAMeNnuqpB40kth1eKfb7efe84xMkFFSOW7gkx86VLNU7e
wd7NkxiJsIvzD65OXDCkPDbwZFaMu6Dwq+o4nNwwVsIjMB+TYdG8cyUJ+elfVBbmN/o5wvr/uUft
r7FDC7r0z6LVeclo99PbA33aOiPfktz3L+G7HdMNzOoXHMFFkJf3zbAz3WWseiBaXW2zqORi6ppQ
y7Sh+V6MPzkT080QBmjyDFNNCe2Thg8Tmss3ZovUywTumhgRQqfX9+u36YPxjW6izL6ccUOlBsEe
f81ceYO337rrcV8h/Y+B4sAp2HZJLsU8iF3CqCY6k78tCw7VhLzYCvXOT4rDJ+h8Ra3wgNMkwfkX
U2ICQM9UmsonyxC94oFsSOWpvh/Mw4rtK2zuHAW7xQx+8dEpRIYPOFcyZtTCDIRFx9Fq7Pvelk7s
QIriN8wEgjX0NiWd1z9yvktNzicrKMr8ZnP2M7QmRPmJTEL/0cbEY2HV3FggQltOLnoaUoUco9S1
hDKIAE9esxaOD5lpNIIAdtIfTRRbUfsrZzBnm9DvwXKRTNDiIVbNJh4oKEfrJVNG1nEYj3ASI1fC
j9j3DycwEJXgFP8cVRUnaRYcOMxdagkPuqj5o4vlf6lYSVVTO5nmghgxm+T4CWD/7OXV/ZSHneea
PM0vL3TaYSpo10FFO9misaBJ2r0kpjcj+avrnPYNxTl+rg8cv7Ps9KzHlmm3b2zUNOesGqqh0iE6
lhg/TdDqb1l2cN3HB43hgLuNKTcl9/nMsUlVWbIOGZ3wG0W27dbZmrnNKtpkcEUpPBh+k5uXppR/
DU2kUojPveqmhuM6XjMWzIwU2N+nqTfaFb9yzVI3D7NtXluN9hSSDf3BXRFVsKiLDsXheWFwGqiU
qY8HLgzj6DGxvpeiUWVr0148ZYdB7uBAAFgyxifMIxLtQwKCj4CIxuKQLqXCPqE777WbOvpTGEe2
IWf2T+46tXM094HXolz5ACBLrq5XZmMgxLY0R1G726p3kTJJ+139fiw0Q4NE+v7v3GPsg85KbN6V
wfks+f+UgBrvR/NyGEoifmddk8N/Lpt9Ab7GhNIoNpXZ78MvI1lccGzBYsA97o43YpdMw8SeYCA8
d+v6TXEGpVCe9ZdK9iBrVLKMtuctmAHehYFQVEEsl++v+n7usaOPDF6s/YUJsDZ7QYOvcDPdIxlO
XLvm8B68iukOeWUl3agjTFdBFmcfQ766x6vuIAEZkiY3pue+UCmrEicTjQ/BqUssdWQuunNTDlQg
r3uMfUsUHuOCA5V/y4U+QhK2WHBpigXAh1oYnrnoNMbs1uhEVtvTKB/aNUo5YCOwvkM3g08fKwmM
hpkmpxeOnfktuhRdI1csBp4inZS0q3mdLH8+QDX5i4GA36AVFCwy16GHJGFQ9qJUJd/uilwcjdkv
U0bidEjqcvAhP0r4Lx6qRZWUKs6m2ozUge8hrgyznwgtpvR5LrhmXiLu3ZYdkvN/zRkTMUinb12D
6Inv7K4Bjeitm5EG1Vr/LmUGUrl1EJsB+SbV+VObinHBuMNrfPUfuZhn3eg4f8ZB1172TjrhIxMx
oiqNQK+MQUZ8qXgiBW7tguMjWRUVfePyzzOthJK20B4yrrgpjW7FbUfIpKjKJnjV85tSd6o+hD2f
vqfvQbsc6z3ptCfAiT2oaiMeaqonxZ5rchqGV5lI0BVhjEgQIIWYLVY0/1wqScgWkWazRb+CiZ1F
FcLZWqdfKSfCNUeVTC2CSYKAwhMYBkbc4L7GVT40tJrsjdPwGBAtMwQ8Jl5+p5fsneUQrzggstMJ
402P/iauHUtSEqxjlV0HPq4iVxeCWfpcoc4G14VOHta77bjRsvzfnSxhGQ7ReBjukqoRAbur07qb
Bs12KxtTLbuZ0Pqyi6pGb7k5Ev5nct+ueuQSV/ZmePCqYgPFu4oARGm9PaRzy5KxuKANSj+zA/Z7
A902MFAUHs8KlgTOXmwbuGjp+EWI5LYr7emz6YvqLq6rk0qUmQy9LIQBJEWvAOCTqAqAH+BZBkoa
oy388b/QW3xmZzGKdhqNP1f5PPvAgKiru9MH4Qa+rZ4BGOXr1TiBnD+ZKOXxWnEpHtP0JIuJZvmz
wWXcnKFr3mHXIm4I9b2GapQ2VVKBpROmULz/RqW5iRzWtwxAJq82wHNIw3LBJKlJmUGL0Picc2hH
J9OE/dKaOU3zwFsVp8ip1FRyDmTKpvy0OJrKcC6xMY/Y77wok6LoT7H4ILa2liq0OVX4Pzfajkx2
bnOZVdO3YnYzh1KVLcaYK5mxI1ZRaYEEX7Z46LDgnA0YUORzer24aVzlHm1k61gMOG7wQVW2AO1n
kdhg04YPiDJ+a7zAEtn4UQD8jNDchI4FrsSm3daPWViAYeyYABxkhPiW1I+sH7YPYK8TXSccAtCY
m1r4lIQQ3aEPxLlqvgDYBDKO4n1QREPCj0bezkfqbJhWb6aBzgCbtFTEo34AycMzgMQHaLHxVI2W
IIdH2D92LmLDkfY5zzmIZQkRPYKElSOEZLZyvGjGDMV17M+5sZwS0ZFU2rpQ8mrRug7PqqbcdV4Y
Bv0FQCLNCbHmhJzbJiQa58ILzwjtkMnJNvRgKcLm8URnB21KJDeE8eMnsGaBr+S3kDEpMJTvQSbx
MiB40T3xZefabPdkiI4mXH+Qtu2Q4hnm+aRYJdbhEQX69zXeVfzJBwFLrpDhM+xqaddNgTi0j494
RVRQC2vexjHZvwU0KiC18bjHVd0yWuSWuxfw6VUFGuxNkOCrprj/N60OD5fQVv0SJ+FRQI+Ismcq
mnUkwxpQaqcv47dcPeA3bgSGmPd8R+XmtKHVyN6prTYWeU6Or+4LqRfXlRpRebgroUsnHno2bQNq
fSOTz1hcTCMrup90xf4B9kzP17ST7co93jQUT8vs3iYSJaCjMKvn0u3Kr6I7ahUYDBj17wbdAvFL
f6NBLGCxUPxWs9jnSqqDy0bGqGXkfD1ECNFfamoXOD4BVALvMjKQCK455EUAvEda+cKujNxVItFj
8wVpr8GFa6JoffX3QlCda48BwgmPoEU1jPTP/yIUgZdeVESgzeXnatAoJbW45qSGRrYAS8K+3b0Z
9kmGxD+mwMh/PIC6uMabcVTNMKaiKg/v3IS5phlwBnLTNWWaBpr4kzqowLru+TLyF12kWjQTm6nB
ozBJT9872SnZ/2bLbOVSDK/FOMaTUkpS7S/qG6AfpE/K2Oe74XoTXvMXbdjVHzDSZSiOWExLViUe
O2QaxjBIk+U+sIPnJSUqBcQI3G6tRtwxVraYbfX/JV0KLK6zQAPH7vAGZaf+TmKQQD5kHSdbui4z
Ql/mnDd1HWe91qZwPgxFeldodZXY+AzqyGeG9LNDdkvg4oEkPtvPcaIgp3Iz3uHfTdD3LB2qXI6M
mVKmwYHoHgJlR0CjrhS5HDn1hs7xZCjLwzqosjG12rzcq7CKvzvuw3TD0JEtMqD+MJiWRwTtlC7B
scadaDdkJD7oZD0RnGOx5LinCNIaUaD85NDafF7AK/Uq6gDQVC+HZKN36IYVp5guSBu3UMwvfisg
0HlqboLA4TyMO2W8OlJQdbF8ASy+CqxHA4vzxDeLaowP70Kv4apY8WKELzY0LaEVU03wRcH85kgj
HzHzTWsZq4HHyIUl8l1DlGR+BcInwfO9Hcq3ML+Y9DnRkXXVpTVHH9kc17G3egpr10D2hbn4pJDy
IfSyhIz2kkzZZ2UL15/qQvQJQYfZ3/enTPaIG8Wxu6Hqp7NMH0c3kRxZMSlWtEX6uZio4en4Vs8N
idhuItiFMqTHxqzCL+qCGbbOWoZtwhg14FryI6ec634fJ6S8ZqvIYoy9SZm1fzQ9T+2SB4kUOGKP
Kch/8xYZM0+ROFP/xw+xG4rZIip6VYvWD/mlt3v48lWWwfDiC4EMWNbxQeTub0bE8ms56ZwyS/74
d08Hi1q+MXmuPOMyBqfF5gz8FMtbH3MgGXNUzi7WO+3xvFW3sVciAd5SzNx27By09ylGsiEPp4PW
ISBc+JWi+g1hNjMGL4pKFR2PfZvCX/PZyoJ3D4Zd01G/vi41av2+4jQSlNG0ZWv6d6ssyQBLJ+29
qS2tAxC1EP5wlbG3iUr2STb/8ZTDvfza9UBcdviVtX0MfW+RX4J0HKX7s+yIwT+XIYUyPDGTkFU4
WtX4eZPbS1zgcL0DMulBIbQOtXjQ2G/R4cRtUDx0b7yyWGJZVOyuV5m1D8pXnptg8aE4x2lzciqi
9FsO+HIfHciENe30hlw0f5+v3cQ6IvmiDMUFAhdG7pe6EOBNARAaP74vVd1efZHgEIgJm4SujVuW
KmX9tzsBDgZoH4bJjy6+vI0xVoPc4k9VgiUvYj5Jlpc6YeQMcPJIbGfkymiBYTxn9NkLRAvNtT1Z
JGGCqnlsmtBgr5fEEsEuq76oqvHcYPBM9BH+HSmPEzFNHBO6bBsKbM6wZGOdG2u4mAbBc7bI2x7V
m0WMKCzuSvDqWg3ljmwfyX+sVs6crS0izY76migbxmjs9ivMUwn1EW1WORQ5PI3OX55vwZP3trLA
72x0aWrxqSKfj6ghcnAdx5+EKvwNU8eBONkh1tLb1VQr26AaQOj43mPCCdUSD1oNT8+gvDIg7tBe
W7h401VB63eY8GPVT9HlN5dLR9OfNyP/9XkX2Yj9HGa9ojKpXEcVQ2qpyadhHwjE7dYgas0V6it0
rIaptOB2Cgo4z2N38E4YsZeKyjsK/bDpoQhNL2eielD/9WFuV8awJwIul/awqhMct2+SJYp3KGgr
kAL/pzHigRJXw4+da+S5uRRvj1aVcu16y9Wy1L+12Gm5ZlxCkq+qj7gXXguWaJC2UzA2RSIgGQ4M
I15pi3sMuoGwukHsNGAq96Sj8emN9aS6b6IEZh+vkeXabOjXxMmHOjg1mqp8hSrr30sek1+n3hxy
GUzumeC43QeanNVbzuMWcvvONr7u/sz3hX+EGMCUcgmfTRM4xuJCe3vJQVToLVfelayVj7LHZ5B8
nVKTMsfGHO3uP9b/+xr4MGbbWpDwFSxmLVvk9VTgp8Snl3178yCWz3j5Zd23joh2+KrbaRrqE0u3
l/HUm0yEGuHqdQNOXY80QW7UoyS7DUAzMHULyuHMZdjCPLznXXoJnCZLAYtDGo5QGFhih4rDpCWn
X55y47nWdVjBZfla1i8j45weYGtOM/FR418mBG6x2zsbyz6qdaLxFVszor8h0iKXzryO9k9B0nLy
t1dd/6ycQb3M65tyB6UfAv/FFMJrubzM2nwcGWti+xZanYb+1kOiu+QbbApUUtUPBZiIKZ/8bNch
o2Qu8xhlJ6v2aNBqst2sEQ6aqgDHz/aoIEqYxCM5fFz6xzQdZJpOahw3xb4kIUXTo39EsSWu+ZuJ
NObbl3DsmxDylx+sEkuDtWU6QFT+Jga4hoE09+H7qfzeHrMFaRiPhW34eus/1Nfjn49oxHmBwMc4
ajcoJ3qr+MAbZDxY3ODQ+3H7OcpyLI3qn+/CVsS1+erYSW+a6QRSodqpzwxmpmop+45gLADA+Cwd
+ZMLHGd+PR4DQPiZRAfOTfT0y+c0Tu210bTPrHalcwPkzE40UmimnTQ8bymUhHxf7IIzcdzPA7Mb
ME6QZuIP+gVPptW82A3aEb5WJVcyzrLUAB4zDjIs4w+XAWgOKFIf01pCcA5ho6aCwpXFTqNQUxKH
dWzlRBIoNzGU/yBffhSXxsPdqFTXE3/6kThsjnqzvSvoSONPNDZg2lrlcFbZIlwc2SdeU7j5s5N4
b4Zu+kYg1DhK8aFDFhMLQ0FJKdUHYKbnhEXY2LkF7Npp6tNxmaAynYZq4VaBcjSnOXBecW0a5C0t
9qm95HFZMzfKDkxI6KLUb4yjtTQDjONQCM5z8zed8pNkMfdxFiYIL2j1qhpSCPuHht4iJ9VKaaEN
WcMCodMiCHSdztS1h4yHegp7apowtYq6Gh3sFV3MhND4TkkH1Nn7c+vAg3PKX+Oi1+xvHRZ37BaX
zalq/zI9hsesllH3O/mJlxcsGF8STe4foXlKVT6zAVqUF3wqbK0J/3z07vSQ0V0vUP80yVElAnwn
mGJtQyQbP3xpR4G4xCm8tSK/1Go/uc/EK0p8847zPblvbfo0Pgn6ua9f+juMggglqsI9cEDeIeFM
zAzCr3whnLUAhbR25it8d5g9DmOYYcOhYQMLsZFK453fq2zLBoehmOMvnOsugyenScEKWEAOFXtJ
5rThkZBx5T9irViSLtEd39cAOV0NGVHTZdp8mRm1w4VnDtofI2EVjxyDFr7G5J6WhegPGA7zBUwR
eI8zg2ho8KUXy1uAVVQTzxiMtXTWpSBXP6NrXoK8oPfglPJBSqUcEyz9bUfPrsjk+QsaYIsfVwpo
TunKPUpPCgdk3s1vBXZoTSop1j+0g7QenP0bYYjrfQTf6kso0mDOywkbc684O04lFs5mJeiUAYD0
+ztMhM0+seekaZCmn/rWpkl188KoE62CFB5E8pelKNycYNKzkNbv11SerdIoSuKu9r1HuqRgouHJ
o6fzgUU7iR6XaZPvWzKtqjswHWPQYzOSDTUqcvwt1SLgeq8E3rpah8+JNPdZ45yLehQRoQW/HpI+
whRjXnkDi9ogHdQqoNdQqwdjjnv8OE+EPYgPuYuHz8fxW/xoVn/fOeP6D+uvnVJkgJOdzPTQQcLY
A2d5OeBnpDX6/n48nM4eHlrXjgLUiTd56D8RTRahT/K04YjwCE/oGc+Yp9b2wCBLOmZ/6X760/wC
zh7MY3iSKq+V5Shl90tlMdBBSxwaU4nbxsNnU2CncG7j750FWhpWGiM8tVZJKZLm4ITk5wwqO8dP
gdBECYRP5SPq+EYXQFQ+XGphPQicdgOgYzSYIYs8Asc1Hpfjqx4s0GQOnoZ5nqX9wVccZi1Q69fr
np+R9wPpVWmdBiIQOOaHjN8MW43qb99Rxu8L9D+3oS4Hpcs03JgkNI0cqdVajqOXu+mdV8Xt2S5+
Y9hf0cD7mtVuZWU0DeyUcvnKqJijt84lzYBV7Tws5roHFXZL3prb3LYnzat+/xiLIFYU/A9Ziskw
rkUDi6DWxQdDxByJd8Srr26GvmJmLK7GecdKvz0RdJRJ9F6MtCBcMG16syKhpd9ny9aknQspXq3Y
Qbfnt6YyCX9dwYcSj+67+csTLzcuuuMjFU5X4pzbduO/DOjsyFnJG2ILc3bDJ4iuvIdZAmkkDLFA
4qoMEINs9dOIpFOlFr5QWmEOEVpNC91V3sX0ehvaSF9uY/uwFSH45F+kK9G8LieXz9Ct+Zpt0i+1
/PjNVSXRQWA+YJNPtWSBSUJTlk7SHDrXHcDYdfNL6pMsirOOuuW+DKcyDWNMDszlS2WDFV4WNxJx
fC8Cn9Vzd6khAeV3GSDtsWFtaxGSlM90yifyQ+hT78mJZOz6zffwMDDRBNLqIXtTOtZ9azh1JNu+
SuOubJng4wOkzE+ICmarO2DK5js9DAcNeUSVuI9cXNjIikFi6DybZt31yuSQI0nV3eUw0U+LUhVg
pcV7GSFUy4vlhWGQdc6WrrdZuK+OIHfwyMKnO7jIQgXp+KJ2eMiy8Np//jju93b39x+FnKKPaJjC
zy6nweorr8pqKSWhq59L1aQ7vGFOj2Po6e2bf8x6gmg5se/jzklbMAdiSKs85zbovNfSswqpzpAM
bXsGdndsvGQw9EzRsbSDBo48OcE4fkWOwqrI0fDLoJrZ6Yk0EkcnebU07HYiHs49zKf//Q7/JU7p
aGFjtpAl6LPJgA+UkBYNgaZEitDA3cTKbXVVC3cFX5r+W3FIySYkzaLuVQ7pe3IKGU9rmWAfuCSp
Sfq+cW8wb0VHRfVDGY3JBR+XNKIqKmIq4vGR1jnmjbjBijGRtw7tWhDsSgd0Xl9LWAyyH/DQpiMM
p7gb+ii/kBnKdQfLv7cuXr6KL9Kk2ltE6GHna+eRTURsg0MUBU3JBdE32y7naeTJfQQdMOpi2cFA
rFruQN93xoSa5Smgf5/IYnpMOQyQXLjwr506viUUgqteN7ffhBVEYMXL3IiKL+NcLfACJIvJnbjX
nXLsi8ZiG3PiO5UoiT2ehdfrYQSju+QrvairbsLXD96Hb1FhIxpAvGioXp2XWTdTgDcfNwB1khhH
6JZ90omdFuKoDIM6olh83VA5QKS05+pe9CNmjCw9PSqy56HT4GRk/WQlZBDQTeyI+H8k+wBoBMqD
wKRtu9LYiFiO1A31jxlHAjHntjDQiRvljsPH9cEU1AqXy1hl4AVbdQDEg+9AO6vKP2iiSCMA2g40
u4T2c3X7c176xgWc4uA0I8NXisthZTRvqLJwCGEGJutwP9Y8DNrikZmgsVq7EU3Mze67xUqndpk1
nYjzL00k25/PoyxN62qsmCBmR8eMZz4FM5jNbsTMRx72YpKd6mc+cxc1eiObarJuUHVhA/nnLn/z
xhoOJPI3RkNurBtkgWcjnFa9a/gkDrg4mp8N2rBseUENt4UoNNrS91JfHHsKcOBI4+52FQk9zGa4
Um5NQl/YfjFhGdOxvG8g+oMzXlpwO4tuysdCc+xTuqkVi9MSB22e9wQOzdgd5WsslpH+dPpWaJN+
65k4yybx7dEFRDgl5QRldxRcL+HqZXnzO+DYjNdhfZWToQXI0CfbwzfiFyTvkUJ3Eu2g8UyP/GO6
8EszYaHQFe0klI0cu9fQATrbZwwQpEP4WlAFKMZmRQqsBo11S0aQ9q1F8+4tyD/DaK+QS+3i8Pce
992dv7PYrqw9mbEvS2/9MXIloQmfSrPxG6FnoUchUroplOVbVWHU6RQG+X3Z+gGWK4Q89MX0+mKT
WJ0sTUdGTr+6y13BsjPbPlEB50SYdOfMl6TINTJayB7ddwp7JYcQwrVYloC2zI6Ok3kCC4uRdAZA
MjJr3DlSyKGDnKApmzxhWWgo9C5uM0KDGpSjcGgLHqXKGmvwuKJ5cStlgPl0LX9G5Og4bR+vmcCL
iPN9iRJHAZJmZEoCNIbuWkRChW/vvLVDSOk7DInE0j98xw1ru+aD+/TqMWPDGHr9MBnr5bGk3f2z
TrG1wMbuQyJhUgl0859G8xXSx6bsV3Kv+bwTch59s3Vr82dsQPa9Nhoh35iYiyuCkmH2VTwKNVY5
AM3oohnmZSabjH8xCSQG/gsHUrJIdsGxdKiiFV88aJaBHy4oeFZ2siYIi4iQGjreUVFV3mSt8r+r
suJ7EmsO4+eeMjXjuACjFyrEIunK3DwLm7DIglFA9U59fll8aqiXRijlAMy29GLmYL2FICVoiivl
M++4JJ/0uEsRIe1XMR8uByXjyZHOPfEk7NrDJ/AhpbAdK+Cu7m9Lynctdn9zkrAvYTFD+yvF93T5
OJF1jwxZcIcmglQDx2GevtVev52TS9e5PXdnbmDg3A6gsesBhUIl6ZYP6OGx7NbgVhw7KO7+dVXu
vmnUHAPdkbFIK9jXihoyqOQQm6y9EJadv1N5TKDv9hwQo4tjkfmDyCVV1w2I/a93tq/mZlEkEFsf
XSd+wEyE9dAJSUTZQvg0eIoqAXt6N4Le+OFP60+7qOjdnJEkNyRkwMlRCUZZEoYCe9hIcD9JBnPy
C5oDqUVO/0LzPbR9ddOv/biliLG5bVn/snlfxdt9t1vD8EDiOQno7bkGsJQL7SbyEKKBDRPoK8dz
BArbmv9kQbL/X6piIN8vgqkkpdwiQeZmfpV56wl8qqTaP6wyDH3aAw9NSjQ0Bk6t/Ia6/viSnwh3
EfS1YAghIk9lI7tCvGnLCLXA+TpvhCrXhFNESE+7H8rYjEYQ/IALrX4Mt3gkXs/5CvSYuAmzHGl2
eovnM1En1SmywTN8Ntq7uCB48me0YnyjQ0NiDFF4VhLE+4vvGzBqvRjYKRvX0NTUE1+VnTmXzzF8
JzY55oiAHUBh3KAp/uImHGo9YJNtVgc3tZOg5AeOGVuZ0nfENTKaTUjlUqskhvhpRYE0b8RvFH5N
hq99BLcwzq2VPwrlPlFKIwhKKIv80bb0WypxI5WWuwe3/m45d7Yn1aAuuel6jH7oWXW3+wSjKoCs
HBlUU+bU1qTWRyLH5TmF4s4oT5OqT1Kkq4xNo3I0oEi2jVIpI1NL4kKMeKIlzNgpOkR/7Qo9evAr
W9mvbbd7k0PdKBTJaJ2iSu4n1P21H+nGR6q0RaqHx0CBksWnA7+Py/w3yGR5vIOgx9DoGfnIhygw
w2fCJvrrdXGgiHY8bTvWZxq9cD/7KElCckNomSp0Ck77lbsvBTa/HjCOq+pE9mMlFT27A/FoObpu
SkC+5qLTz5D7uIyJLmaGssJ7H6lb/QYh90xQiaHhApE96VwQVDiONEPwGhbXUH2BXsq+9081H+MN
T/N9Jy6iMGEbJYCs5rwoFDYcoQUENv0f6y5RTlQKJDVs9LOHkwIQ3BBRBe70sDqRdh0QIMIbCyFb
OMXIeOntXC8QdTjokIeIUtY6NgEBZThrP/Q9kiK0SeyNS9UfIiYxh0za+8E7uCoBDF39ItH1CiUZ
mu03IJ7o8PYgDvpQPP5cWrjvhpY1PONvQePdjpak1ynCtT/pZqxKUy9SrUvNqfrU1aXnwNwIJq9g
0WKuPsMt+/jwGPArgpujB6BfIyLt77Mlw4nNnFZcfbUvpKbg9wuvQf/yp2JHgNJ6hVrnHzyJXCdU
IKqvQ9cqC6KMyaEgzV+Y61ZsxMn9lAfE1CoXPzFpMhKc5l0QLUyByEZNv9bIm28v0H36t8FS7NTT
F0++e3PJRWSKoYZIx8rScslO+4BtRcFZrbVmBCkTizm3oe8F0jdYReEC+iuULAWEZOHt1xnpvOBU
NOo9MpXg1V6Cm4F4ZdxzO3xeBW+zqwl8FFx8cSZJHYg1pOERPGImrYIOc0uQsvPi66LC8MqRUymj
klMU8sqTdXHkgggQi0MDLx4/6ow0RX0PGuxaI+bKxfOlrhhhFuOGrUT9eqaUVLKCuQtPZgMT4LFu
Ty6/3Su57DG1X1zQk44cRYWwpK9TdP5QM6ZznK6ct3oi2zxSjY9+6wr2BEjCExPeQ8ICAqe5fogp
cFNDFbQ4Em0W7COQk7W3UZhOoGptzti0a9jk5EbQQK7kI06BxAgKI+Xh6949ilYV0fqRGyRO+yZ0
vCSq1fRAt+H1+PqDVXOVsjJWVFi5f5NxnvPnK8rgudQjac1n2hkJSq61OF824y8Hyo43kMI2+FKE
uL/MuTx3c7wrCOh1QBzQNJy2ZhQbqIII5StV83dAYCDF/exQbIYKpqY8rucq/ZU4u/fOhm1F9FMk
4iE5N3xeHLTA5HQHH6k+Y+6NiYyZn59sQIsBWeRZ9HWnl6hCImSw6gVGe8t+FGy/0uzsHr0Gj2ra
yx12S52bO7xwcs6sUH291qg4im4uT6NP/YMX76txbr6W9w0hujOOKEnelC5uL4Zf0pbORPyUgLaW
TtmiJbYxat8xIyoTXgEFdMcNeKgvkxctCrj2VVlZ2sOQnDfj2gbxHS88ftBrkNIcyE2swEpkqxQ6
ZX19Qd01E+FGtB8pyLJGbx7/Fcc7RlSgGvmo/xRWqSBC/2v+O3l6zYrECbCd6wmDZHBtNkf4KNlx
JBCw/0lvYBYX7GYp/qX++ZlMOMRk/LKdswzgX6Mg36vp8g8BFglP/o0w1StDhOdd85NQbYRZ87OY
LLdMLvvgpTsl+MJvelaHrS5cZrAiNr34qT9wtmohoTZPVX93iNYVGtXB5DL6y/BtSdG1PU6QERss
LBjkn8JZtje19qRLPLR01rQsMS69TDNpCsTO7vC3TiN6aNSXP+b9cGJ5xPtEfA3P5UImPPttI+8C
buRNdvwpugkoCLGSWAlL09jZP8LpUTh8oCkQmGuUqaw5e7LkJ2MEtvM2M8FqWvCiz5C1erScZQGY
v198r/lvG+u69HGVNitPVDxqvPkPIrUTjgGnWF+/4Y0fAerdfkbcb78wryht0Kn30RoxSFCTkAv6
4naP2w1KwZesSBLQ1E9SvXHdLKIVd5bu6hXuHfXUie4QVqAGl4fQJ0HYvWK0Nb7+KFBsHYW7Rr8T
UIoFaOna2CA6W2ySxzkhb5D1swRvyv41NfY6SbJu43wR+wF4A+WhV6Mn3Bk/VxsK4RXP2+v++dNU
bFs6Pu119yNhXNuM6wB3SeyMLgKVT8Ts8xSQIQD2CA74yNKKwXN0tgLuXVJ1oJpSZ8EJW4svVFDi
t2cVl66+lNh67ZBgjrGt0MFYIJlUyYGAy9Wy36MqhfU2HF9RpEc8+wn7gNyrQ7cze4tIvV3nVs4Q
UN80EpE4L05mFZFhji7FOOpSLK9yWUaKVf3TBAQsH31Jdcr4F3GUmDzxYDDT+tbkgOAyn3IHWl/I
vzt12hnMtD9dL8TAylkqW53VhgbRTH+gEeaSeGLi9RefEe9pbDZd3YzxVNfw3fdNm55O6CHPz31u
1UJP68RQwD1GxHakGUPD935PAu7DkSb5D1ZHG5g5w99rn+EaiHsiiPmX+xUGIrOYWwEA5PHTP5Wo
LCggv2SdbU/2d+MBiBSPykRViz7c7FI/tgknjW8/XYIlsfplcmkzyEJ2o5gxzVGA+7GLGpiszINX
8la4b1RAwvhntV6ibsvDp70ba9GN213m/EwvvZawJNOlG1BjhUORwyasnEJBPlot/C3QR5NNZN4p
n8uSPxHd4PsCg4WRRYAiZTK/o65WsPrLFlmUFRBBM0r4a6ntwMaXTYPAI6w/16vwlx8yBmfmdDbi
64YI0xob/N3/6X7ZPh0HJVXabrb35JpjDAzJY0zmFpv+LzfbT4J4uKwK1dCW1hLRQLmGXemLmRI1
svhwQx/IZc90gW6CEC+yzz5gNY0O2zaPeDZv7rhEG/w83r6XigwpbwvM2AzoEfOlhGzkiQOWbkMi
w1MwgQqOU4ohblzt6k0PcdSepgDdufnZ8hipmiF2FBlE9LJQQfvO+nMO4VRVebjRkRpG+PxjGOhO
2yMcWzaRF+fslpiYRrGYcEnRSq9Alk4o2nOLpJuPtPfbbUTKYEz6WeLVslrHpCojS6XHR3kDsO8P
PZ7U6JbEbbdn9Ww97eDpRRR0b635S9X6lZfe5yiKWgArr1N2lhW8ysyGssvjcU5AFDiuO+kPTvGO
voP+jGeFC596SCbEIpG+j7/DiwWcvmG8UsxWtNCJGuB9OdspsF4UI0+RAkIBhfxXfjMZwS1KDA77
Xv0XWYn+hSdGZr1WN0xSYVmyx7OlswmRGJ6wxWsambUxRzo9qRvf7u6D+FSy9a3FzBUGox5eoBbE
QpKuDz7rca+44WgFlcFOCJH9g6mDXacSv6joim/OIqz7hgyYqc07JwgmMoaHcUR4FwTwaegBmLXI
MdOxFmp2GkcEH7TBfw0E3QH/MLJtpFKnjnjNxThPLixYl1uOneDHPlgoGi72kpdBX9RPB7Yz6Rjr
Uq7Hol+1937qfZOzpCqYMo593CChzID6//qQQwiodzMyNsQrRe7AeEjtjS6EoXPvalPLyfceuDuf
iWtIW8tWw8Ll+TQznP0brjXI3WTsLoWh5vpL+WgwRhqGKcs0gHGEcKaeCpP52DCS6+q/uHNRe5ep
QrI+NXyi3Uwi1PWxol0FECc9NGH3ANhzOJm5K/HaEw0Hz408U6euU3AOwwgjolTD715JQmaC20Cs
LTxlNNZvjQ8CXgj27vcilpdudNDvvpPctpJhjjGVHIyuwZbT7CXyCXU+iRrfiwpXzUs37EO0cB23
Qqz1xfGhFhrfNps3eSREbIVlyLVMMvO3hafwYfC3iHKEmbt3duhR3Qy/nAXA9WTwM5rQGFfcvgtD
pj6od0EMFU9hsXSy19x7YgQEeJfxClYGttJbY0hpzNCGLXY/uZf/XQaCoe755jnnp+xD+h7IRasi
YdEZP0+q+nFEPnwFKabFPPCoL6p0jAQIEQ4Xvdf5QA3GxD6Hb9mXE/4LqxicKTNLS5pEawYt2xcr
dPFTwm/FphklOC7zhfiTNllTIrGyWQk3LNpSBQvhTuFR3QzozSwQnWbjW0WWNXDyRNRco9Ibi4wV
lZBOkd6x7jvIy8dR0XSDx37vNMdiC0c7j2iTSHVagXlxhwI7gqry8YyFI6EEU7jmi9+7xnUM+Qlc
whetYKfA7N8FwVPHDhrih1scqQ7KB3z4U12s9ZMTZQhT+W1bIkY8AyEKN8EdzPMxHAtD3PCK3lom
9oMB6lguE9nSjkAxi3MZnZreZZBUjJgSMZgThkyOy4CfAekDc4mhgZxABtw/szf967nJtnCl7cW8
spjW9GJXUqDPolteumQtCXVo7Z90Qj2iz0VrZpXwmAEQy2AwNEdus3A7laMJncWjuQgAAL6kuaLj
xvM1z4A1L8FtszeZaMfVG2tZJ79gPbQ4SOhQwDh16ucIDuRoCkjGKxT1LvCayFzahLUMEO/nWghx
HOeTzsSMdHlDLI5X1DG4ME8RaXgmJUo7toYOmMu0P0+QUbBxSLR14O1+KXVueyk41f4svPDaOC/E
StlfNtr2CdcX03kQOM5pWoH5opOehdgRbCtdWd831sD8vno7XpEwS3WRnir4bqz3cpTnE9uvk7Aw
gMasYwKuC0C6kqOkC69I4cDsMdjda/tsKG4gLKrxQp4pFgXkfNCaGghOYFTob24xy9f6uZns24G4
ZZ6wKf+6a1/7fVY5oAah/YKZ9jT0BddyAvVTpHBGrW6j8UAxtchuzpMASnYMZ+2c858ATKbyt9Cm
jmUrLxAMUmkxmZ2nfAvc8xsVQNzojaFadsHeXHAVVidJz0alFFZ2johLb+hLQFj36nQPCcNBEMsZ
isjPaIanqWPUPRzlbnbuYlifFVskTJuuZTVYz1e4k13u19YcA4+EApIuXscq0Az/qjPFeeMwSw93
lB4HCOhNMZQ2NkN3CqDBDA0SHPBAalXZ2ni4vLEzYoUmFt74GCknkXywnczF94fmThBaJKKfPzu9
yGBAuJeKVsXooqgyFMQtz1Jivggu79OpCFenFnD4m4EVQjJZmsdANd6R4Doc2792rYw0fGOgP4FP
ncMufdF0FmchGEKRCKN5cRkgStZ59wG4IwhRk4QluIau5STMfGJUBRpKXs59SApT5+J9nubhnSfE
PLP9uxSUzeFU43qtyxAbvzhCGW86gAR0j38Gu3NF/fSx6GsJT6GN04//TUrRKzHLmdpmExgqkTz/
bx2DxtR/K0S3by88rIsuoQmZV0i2amxm4pU4OXNb3zG3Xs51oxEk01mOQTsUvJh656KsJDWJcmed
iv7A/tKFEt7mqRiZzXSNjpN8Pvb9LpO2Ze8MWr+qS0j6LzivBnoWkiY/3F35lJJq4jTm1rIsNw7O
wkZUBlnDszjOdUgrwVfYJSN5aoA8OxfZqUAXIKI6tC6BQaVsFTVGEZLXfQcLiT2h+H/1jOj1cJb4
AGcR0kHs3jkKbLwXSgHkoyBz2HtS7NuG6fLd0qU3TXCOW+LJtvHc2fUCfdtq+iMVRWoaeGKomovc
eWgHgmyNqa9MPardT9M44ulXWMUFezZPHEPyeqoujmZF/Ts9Ux85Hrc6JF6eOCWoDfpZUxpZFIsh
L43GbYpuZkIQNkgbPKbpgQYsAO6cl4QHIS7/YUG2L0zmhBTH+9Ck43nLBfKM7I0DG8tiddlYw/Tc
nxRP/9NSxNyZcaNpT8QgD45Z9CRo03MmmFPqYATqejSnRjXebTKpMbqWsp972YeZkVqI/iM4kpc7
rbIfoRmP0HOZxx3KQ1VS+y8nLp8BcjsgWIuwOoUqgjsfUCvibFdrl/cauOrG8f9L2EMiJFPo4NmU
J/cHf9qKwQzudh+kV0FS/mb5wusLwzIJQjE/YrFauxFIMqA0j71/uUEK8MqWhS/yJklqbePF4U6A
NR2KNK49UmcWvDgb/hBKZYuUpYQ0gIJ8M1w2/miRxgtJ/kSGJ7gac9h5GslsKlEqfzzdK/6Y3uN6
8um7+Lyw4UIYII2oGR7o0L8s/eGpYLam+CCqCklw0MaMh21V4WSmb4a20eotcjYHgCPt6BTBx9Mv
RoeBXWsb1RZbxpf5g3ALNnnyyNxNoITdqCXKC5hplE+sq6ky51lAzjOBKRSp+3bWAF6SkjgayLYb
LZ3gSBCMouJipXdplzI++FmHZeTAjwczEt36igncrcu8zfrsElv0sp6sm0kGD8CClJjL0YeafOHP
wZdk6WY6MnH9Fw/XUdeRv+tPw28MaM4gmuU16UzyUJJHbInafmCUdrUzPylx6DFeUDn2Ip9SiwtF
wJy+5vHI8L+JdhmbzUdHXzchjCkDdzEySfOEuGlzMksmoCyoIHiXCxfArtPq0ZWUYbG+G/9j3BZ+
1RupxP+KfrCKEqT8aA9wSbPOUplN7K5htXssP3wNNGxr8H4+xuA5XxElRxWxkljE7WdGK593a/E3
qUBR41ph8HidCqP+KoTF+4RMvXnhm7Ht5RJiHug3KyYkqbFMTUjzv4gnxJoiiiJ77RjILtrtvgd2
X0gPnnk5g6v2dVN2r0l7f+oLJsW7oHbRr3ctQT+V+TBMO1p9j9qgAP6495JynnTOlsQTjsVFef8I
8nInUuYnf0VAPVUVfkOH27x6lAcB6Wy4ejcBhJV7KXodokysTVy4Hm/pVDRaG6CyfLNlRlasPpf9
39vRzy8ZzHwwKZWy3G/hnCssZt/ribuEQkK45u0KlbLyQBx4np5hZR/5RuVn79psB7Omuw5OA+SC
dKaNr8zkShL07cDop2UODi4Tdgv9+t/tARot/eMIomPRi6UYm+3lUGNnNuE+WaDtBjwrSIV2NIxt
6gJPagi34TiAoUj3X3y1o0T+ubJ3ZIj3Hp8RqKv+KSW5LsJ8/7HLW0xI4QKQ4XBj4L+pInr5dJkh
Ye8boNnoft9GdVEh1psaPtd+Fjtplm8USVoVMlKRKF3Ged7TafWw67Dy+/A+KVfHVv1vwkrqwDP3
E/TFRXZtUB2XDH7mtRQJS+X9jlVLXWYN3HkaFepME9EOGJUlkIy5DZAaq3BeICLmGhRP9KaOu676
J/EL3P+gXBIMVheL42AoNFFKDzm8A26n86rVvrNNrU6GUnK8DITPFC0OjzDSbLvM8jlX36oScLur
TMcqy05zRhfdgGtbNBa40qYhq7BWY8els0mp0aQAW1tpCOTHkWSwR2fHhgvFL+0hqjvbbYPL5fQB
gSgwMxOXzt7Jl4adf0Oz9pB7mSMLe/YrE8ohNPHxg+SNhFoPJnV+GXKPkAMG0Zwx8M6TtxeYhXYT
7P/UVWkhIEDP6EDqZlYO2+uCQdk7Tuq6BhF8xUlctp53LkjsLg/9UhYwJAVIfcZl1Gtqy6Lr0GGQ
3da1aIQtJz4TYBZaBNean94tuCYViOQC+x8qsntQ0DMlyfE0p55jyyCXoCSvHSPHmY3L4RNV0Lc2
/Cza+vGdi0YUJfMHCUh9GdJva2Utke1d5kFcUR6q+O4zBzsTWgpt37wSbcf83ddkj5RQR9xsok43
TWRzpF2RrheAY6KLAgeAoZMpZr9wIghUi0Hw/n+wS4aRe9ByHVu/IyTFlcReLxorVgvWRGpVLMAg
bwJLZzmTPlYspNA992ze8/z54gXXK4OWTexzd9ozo8MJOlo4N6sHv4DA6PG/gJe/DtQaNDMMdVi4
qBjh1pFzKENydRJmVFIRNgnD0gZJ1U4ViMMbN31NEGrBX3bgUh6kIeUdy6VbpS6kis+tLjK3lCSs
bTdsAFpLl8xZ7PwPVvpl1YFiDYo8SyOWUFqV71NzNZsmw5etN2y79wNhm0yttYfzke7yMGvOvr7m
nz4Iir5nXFpUnQQsP9FCgBqnDec/u6VQchuTBzFnR70D7yWnbEAXJR+IWOOqyddDkJScCHcHutXR
MXguOA3wpnsHqhTKzJnt7rR8P3b64MmP+BPmWH8oy+8SoDzZRoGxqfH7Ux8Wm741OrQjrN6RZ1mK
qYevpcYuiEM5H+oP89SIV85Vqj71hW21pG8e1UrTMIU+o2ESeF+iHdVTkX15eEBs12Ow6JDU5KWu
DOehtY6TMuaxhAu7I1aGap30ZwOx9yfmqhemgwCIzEJgKm6hQx5EC2Dd0Dqo2Huasi7z/7D8VWsc
Z8AQifscnu44+rbakPl0cSXfx7U4SM21N5IpTUS3jtO+w6ZNg1ExC7KO7HW+0q9pT3rRJy5152Cp
s0sQiyGjicHz5KPVrmteHO0puFMTlwEza6V+6xEs8OQpv4Z9W9/A2S2/fIsOCN2IrFfbe7jKbwFS
GoTKCV/aZQYR34OUOkJ+b1diN9db9jVdxRTBRACJAE9KHYZnQ6BaE+kQMNxUdSezsow4Yn54i7jI
wTOvAB8dacdwZGScsENnhmf6JcooQn30rl3Teu20gt3D+hKUnsbF3fO6MIUNGsOX53VtyDbe2T4C
QWXIc1xT0tIlS7MEaYpBEVBqM9Gzyt9u2TOVOBpJnChPO9TRiRCAg5r2M9yMd7r38rEACzgaRdsE
nJZg4Nfyh4UT3ns7ZlwPF5//OtVNU33IKaOxC6Qoiz1qceb6d1xTcJyndEZYvpiw3deAgf7V+Cv7
ISJrQG24hfLWS87t8GqjpmIl4tDkM2Zy7wL8IbpfhBbSIt46G+xFhSPRYpFS51DioOmXALKkXC5U
JXCet3iNy6CCJx6NA29zCoDptQUgkS6WfUqyTo+Xhhvls+ksEHgYetWmdDLF8ZhlvJeEhwknD3E5
HhPoe7PLjuk1Nq6iBq20ny+Cz5hiMq2ffuGnxtaC3AE3yo8SqBl9/Fo57cV7Ac3TlytwxrC16Q1Y
imUtLKIJ4UsSZaiNc0zE4S0U2m/SthGmO5UPmr+QDSXfrgnJ+8+IHh6hs4laee/hcxo6aq+owmME
QHD8TUqK0ELCgCy4+H37D4Z+GwNKujiN35V9zKuDCbah/Bo9H2jU+3drnt4h7kkB9KrlHuvM4h7/
qVEbUOKbIJIN/1vs9x3qRDvoygB9btkiClvTsoQEWWAO6DrcvcGnlKydnju6y4HztjPSaNGfbKPh
5EgW8fIc1jatFLcebUrU6YgLwmIaQMIk4TPjcCiy2pvmo6C3IdJybtTQTCKlcjnmRiwxPEUyvDKF
m0TE8oUe/WuQwKQBdWnhSBtE8dqj/NR3C4tcKbjWL3XXE2iw9JcpH5kZCmafSGLVNMfw35xxodT6
/RqsI3qsPEga/c6hvfmB+ctMTSsG+2jPvePChIX7GNdyeZ0eksalEX0BVyleax7oY3433R6QuRls
i4VhxZq6OUHaZIqOvH68QTpD1ipK+jJbSd1rzPwfIvr6MJ9vuURthpdGTCx0yc9jOl2FC7Z4foou
sNITV/DOIukfqbaJxp7zjLFea4u1RhFUcMZtqKCa/k3osAYVC/Z+c3RBXrc7Xr+NQdNeypRRuqwG
u9VS09A+UkcA8lZICUZFsIlvmg3p7DfxHnKNUhH9SxQb6hkNAf6cOedDx5z7f490har27lprCzN1
SSew/cDgKZlgrNBfNmjkOefeHukUJp1PrZGN5JvbAcExUGzBt6JpUhmMsUyDL5kFG+6yKmfZoOGW
+Otq3BJWpsrfGrDm4uCZvstOLTYG6xF6f9+D1v9SQe7XvXGC5YVegMN9S3Q/JWmFhRZkSGrcGavu
+4PsuLiKJ2jqbOns6SPeWwBZCVyQfUKOBp0rcBrkOuF3xZN/sMDw5xr6XzmTLGZz4DkjjP7TcC5R
90r3duX6hN6+3ewsn5dc+/0qGoLhTko1Dm31+XkZ+EvXMbIBQj+xOuls84Wjz7ZNXQ0n3SdZkZlj
1KUmmyQf/Iuvxbu8KSDGbK5bWip0lnqvP7PtHahpzykhzcNtfTcMtafwv36YN2EdkpyajV5DkDYl
1F+ztrkOFB68MSG6nC/6hhjAwyXMflvSkMwYS1CksKATdCwdXCR4tRFjH59WhkfFsDQbMnnsRm0L
6ZoyED/z/QlGl+OFt1Vu+wa2j1zw/24kmXpby0dCXTv6Z3KTddcOwcAd9B0ju7LT++cXquvgIiAa
YqnAFPbJIStiNSovzbCPVzq2wok9KTmgSmS0T1gZIMM7+EK50LJ4W3jKnhyZ0zan8d9MIEIyQv/R
oV5tP6FBfy6D8av+idH+K4V3NlU2GjRXA3oWYGIr/MH9Ln6+cuMNI5148pzwooqKpZudpOjFYHUm
dTch2njEUXKRpLYLk5VzBoANijcO8acMq1fRiFYErG2/COSW8tdvfXU0ARt+HlIPv9N0zxT+9mcr
oMKx6SOhGRmVlUYXY+SSjigpPlVl/te+vj04EjhL5+o6K7LQcsaLov8xmbbLuebxQ/fqWDudtLm4
bCBxtiyscqncu3rlK3fkhfO6DlOBBWoHaRAuREhy563gRSRifLxe9d9rNIE4l2x+5Q3WFCZR5RML
w3CLHVs8L3azxPmiuRbl7+sL6UfOVXnJAqZugHKgQHKN3sclQBr8T13qf9YAQpcrPpVGKK0c79Wt
p6OXmqOIOZdkE7xi6pUXR7OVxfG/BjFqjlgEQ/z/cw08fiVDB2ju5l7MV0HRNPofOxRnLn/U0H0M
Bmc/M29Vgm1YSftWVTlDyGkoffxHWoabNNrc7SqA5ZBBQjMoKJsxNMm+sS1ByhuDmIvpnMVYV4WV
hU+euR1yYNM7TnEqrpk05xFm8q6duOH+OEllMIh2YIsiHo9kW+SB5izrM2Xpu+YBBHRCJfuK+3dj
Y7m0QHxYh5cY8l0U89tUONpitc9hVVfe184nk0cDd0BUz68m8xwdienXencJHl6yJSJtF6pnPiPa
n8RHYQSgY+wSlx0ePTTgr3n2RL8zv/FiKRqRNIHSpcv4hDlw6MSIHkZ5yJ5UdSO3/EOkdi+Y+bUB
waPsypbJtcu1qgg76sbau0WHfTGQOQ/QDMKr81DXRpZPpfYNitHJZBTundJae6duFJMvqFOXSfrQ
TNkKDT5oKzptiQyRxuAuXM9WnB9kjrr55BY4ybQX4c3A2nQi2nBW94LWgNW5jj+rxVoo06fyuwe+
vLWqohRt+LC4JY6E1ENLNdE1N7YuopBm7VO1jlaV39GgYG2MPFPRiDMH9ZNaMcqd9A2491DkU0AR
NhRAiFH6FkZlCDJpXKVUBg+KMIpOcU0PCLjx91faVmSbLs9NTn2RS3Y5T/0LnigqSg1RMJWVQpJ7
7czpy7zOd5h9suqQWQEZCNm8oynuRL4iVLL3U4/q0caHifb4ZH9nvEi6yZ7h8EbEzqb1s0KpSzzQ
Q/uc77zvsdMtzmVYLbjGbiV6EiM1cJV3hAcRM6snSfJLHVMW6CulqHHgF2IDyDWEgnypsX9Cg1yK
rnIC6x8sMXwBp+dVOwz8JOhKSTWlmpay3o9lp342aGRhCTlImq2K0bojGr/rdwa0GLZB68fafFxf
OTYWtRiOfMd5862f/KLwYBi3uXq+l5nA9EQn5GpQcmL/B+G3BwTU/3sJ8L3tqgMUqYf/ktssPSpZ
lj3hhJEgEXCPz40qkUSXVs4c+Y9w5dYsDK9tV0+KHI6CY7kJc3qVp4oR+ONJbTvSGdtj/KqQhr8v
XzmNCu4Ff2i+C+1CWarlB5CoB/Kr+g69tYN2PXfCK5bfGngOEyZtsJJMUSchCfdpfRFu8rdFlUE/
zcrdxbtEaF/AgWYk+hE7Nx++4fGu+A1m+HkEiMkhg2khFTNeE90IvIjHt3iaglRbMznGpzjr+yqG
LYmpxgeIue9QSJfD0T7vIp2eUenghst86111wIiW6Aohanu0nAZbCmkKu+hzFTA66xbhT1wxp8Su
TDR3nk3fzR1PT3Xi4dUCZj0i5vE8QktSZgib/5dEybTBRP1UNUEBI72G002XwHHrL+JNKinMKOgc
/dwdCr0bcfhBzfz+t3osJio70Fq3cVY5tIHJL0bcClr8930mAS7vU0Z61qWgf8Ju/zNLmw7K8GaG
NtLz7bLzERxAIy8gWI9uRfOPniXims/K5NjGpxuppOWRC7Y5/LV+fLTsMsTjeK/9MAvhwjBDP0l6
o+btXlPclB0vM+PTEMDuR/13AClvTFYsNOqQHVgTvzgNusNdIrNJUfDHGX7sdk8t6EH/r/7o6kgJ
4XJ4CQoyGprJ6tFUR20Y8PzUMPUw9fXA2zWUFjAbxZFKcy5DtQCmwpmJrkZbOVJLWNJ95Q8s9L2x
qqXhXcJlAax4cWV7fA/SzMicss/atg5+JSb4IHNBgZRBO53IXOubB7eDLKeaiPqrtaDgLhsA42Z6
eni0dS9tdyYe9soDIlRy7o3k+4zAberXiCtVT43YxZVnds+aCa7NurkZbVfoJ9gXW/2LDhPLw7Z/
L4t5kWI2iERvuMkHLz3VaNtRUC57V64Meg773yuG9L28jTXLbUXxplkZ2TlVGajh5VX1WP7M/KCv
7aSk1VlEuBgAMPPCyh0oIVgw6rGAo6+vXskFXJiS2ZdTgf7k3DtPnPlhNa6wqa1CuCJf+iON3jtw
7zzwx3oD+qDWYfkv6/NIcsM5eTa8sPt610OpyxhsqOAENOF7VtxK7FAov3aM3pMrs4lJAP1x6Cz0
c8S0sZeQ7xWAdNUIEIv9HtOLI+/i3slLl9p7sKjrBfKs/fCqSB/3tqF4YQ8lBvNg0ojEEwv1Q+tm
/T5R2NWO9HIxgnfohcr68DbJZ3z67/ZBuDFN4zqbjCLnLkMeHsuDLXC2neGoxQGyXnP0S6e1qwPr
6fTNJv84FIU4XI799ZKTuBY/L55znxhFcnNd+Q4FHEVwgW5amGbTgLaxOq/0PfIne3TihkCkwx67
hCfBkRFVW7kVlmI1Ka3t0IX1kpKiu9DOuoLTe+LAoX82kEjsq7iuoHUcqc3OlrpE3aIvqDKE2cR8
qaroXS6DnWHXKnj0y8cwwgPkLVjKEfqN42/xGJdePF7pB1hlLRko5UdNeiL9R6ycXrLv5lOtNkfN
vRcL2pvKVDNurc/HEmT2MyAHJ6jgSN/lLGK9l2EsxVFzvjffW4//leQB5bCqnde19LeLby4IAMPZ
TM3zLBSllmmNWb95Ne6YupTHY275ETbXY0ZMI9VeqNswnhIZ2Nx7QD8Jq0UbkzKKuC4Wmx7N5TzV
8BquATV9d9NxmD/6nf/7nixu1XaNLfA1Lr16MEFSuP7xOb5Be2tcCxkyYi4mEbUYDJToGPLizkj2
0FPhie1px6BJdgRrIHYa2FaRdaYb/h+gP1RICeqY6TTrJwkmlZMGjRiypdhEY0xjD7pVMniybYnt
+1NCXrim0XsHFQMM/cxOfuwmNmMbnKJq/oYyhu+synJC6KGc6D6ai2uhdRNVeQvI02Hh0Frz2ofD
NwoNrNkUD5AYY3N5spzQUFIIlNarpgTImemnegCjTxSlCyAlk5Pjc0VQorYxCXUIldjsbbVPOod4
F0sGpiFz6SM3u7IOfhaYqVdYSmvStaOQSz/EjFUXUawLg78MH72HGUn/Gn/Pzrq7x4nKOwCRhm7M
nUdeZBzgswAqxCTZmWoZaK0FJGtWmo9JqoebJTwFgW2jdprW3vTruJv2ZSH2mmWDAR83vJ3SRKOu
iNVNWl1xFQLZg40Raou0YMiwZJBKcfDoWchdC/Tla829ccX5jq0Gdh/4XRHOiFwtmRCmlIe8KTwe
yxH2aGkAYg2RD6axGL8F0MAF2XAWX+9jngH7wyyBn6/fg/JaLDZBUDxT752qnQBBnsdolzgsFfQw
c9DGZ9J1qLetWO+797qf5W+VVxybZi1O+OGpq1qKn1ZbF1MwBKn/POEzSi80nF6Jyxf9LVop7+V3
zni4Xd1faH5JJQLh0dCByHuwQdYOAYserYPtw5OIHw1YIhsDMxGVyagQX/7OyE40+qJrYhsBOYoN
CB/pEWPPH+J1T9NCWhFsUaEP0FEwC31Jhr8hufKTFcaqiPB5PkaKBbXowFJ/cIFLL9S1ZxAjOgQm
ji4eDLUERwSCgkk9mE+8lGut4S4K2u3s4lj3PCBDErf+8hZOrv/CfdFpPBInbQYIhRCI0RZZWSOR
jcSxqJYTsnAqSMVHrGCFbKT4n8hhhdqdrQwyafpcGsYw4p5AIjGCpAuR0If6fKZREYiFRMolyy4B
puxC0VrOQbwJne8F7AodDAjgGHGSeSfzKCoGsIyETf9u5eVztgBW4G3eypwvQ0yfm1iPzVHuZUvN
WAhuXPhjwV0IrLlJtD6R2BvU2ut1NUHiY2uutNbNH/i8niVGkNOdTYYsw4uhgkHW8SLrULkemKIr
orHPKa4uHcfQPAEtZMAh47B/o6KYhJh43blLMzrvmR4MXbTLucyA0WcEo8dCws5MiBne01gO/tzK
ZnOdNYOkKicBA2XO0FoU+0anxyZ6F0cY5LlyddJdhjnFXKXJ3TIASzh+lLudCiZ3GrbVgDdYB/vc
w59VQgCJ5FPSmncECoBlionK2nu5QsZqgHsffrPnHYmDGWc5FrEVGX7v1lNgwOsuP/Joic0o6TXR
Df33E0FInd6WBK0I5xcS9tTdaxjdb/zLJLPEMBqPE2ocfHv1IPT4v23l33iUcn6mKD99/9QF/Zew
oLQnziuRbeIO2vpMC+LQVW3iMLkyJeM1vRaJBpHe1YJhOe0JZhL4+p0scr8thPYLw2oOjGX0uuF4
N9S5QtVwiOpPflR1c41/RXO1xcIs1DMNWCt2QurGrJceDoVAKxuYaJ2VhNuKDBx59O9UyuKDPnOr
HMCQ0vr3VRYp1lnDPJ9Q3fLStsa6gS1QFQwIG09TwitzyNeyfWI+ThnxtAd8sWOmEViVzz8rtWw0
zQyazxEFaCbL1TzRREHlaWVUOerqfVu5Coj5nkwws4kBlouEd9e+tXxB5pXzNH3NRAI4ttI5cqDN
e8rKoHx4y00AHHLSiPio+3gmipssEm9oU8C3NXSuh5CQGWyaIUDKNbP86yA7ylsYfxPswymmyRmA
Acu687lpY4SgWAxDm6SuL97jtXvxBs9KAQf3hP+/eOb8QIs9xr04qTCMMtOIFM8/+mu9yq1/De7Q
4FrEqAgi55lUqejrN2ycPFQmv7gFOiM8zjKlYKGGc/Y00MfFkpSD5W8IWLWYMEVqucYlZacTWZVx
wHta+T/n++V/6rmvBWCcz12kOErh9tSvgdUvgqymGZhyhibtx2GpNLC2bsJfy3Wu5YcXMSopCGyv
ODZM/U7dlSD9Bl21fS6ikinUdba8XY/gNt4nCYj2qYI1oMSPpmETQJAjQKzUxMwqHAm0oMk/5yOf
XLdw92rgB1pJ4mJVtUC8OIoKDGZwNb1iD6m8tW8VBE7foVHxW2osGWZI33UzNAyCTG+Ae7tOX1Rl
usraqkwOi/v25SEKZVc4IPu42ma7KS8a3pigT3lSLIUjKznjas6FQn/eAxtbBkX8NpsD5fUpfVdQ
cgN3v1dbVQM4f2vYCk7winmrg4kfDGz61kVnGg0phzLIx7/NyAA82ikRB6Of/0sK5ByL1mHbg39z
Qi8Hqyvfd74/PLTzUBLLkYnWO7sp/FE/v8qk1qF1cEBAtcrfA47wnl5bU4imRrC80I/F0UeHpJYX
2cJWUqfFBglR+4tYjucRWYxT2YVfA5W/S4k6pso+ipJYBy8bPJu3Y4v5+Wk6hJZiitpfgSLn001A
EQ2Ntta+xe+synex9dyfe7IsjN0ny5BYLABuZca9ARRXPUllzbQ3luL+OwlraeCdzLHzjUT99Bwd
XKVfAAdFFNtxFo6ICj6iKZqogpTxK7mUX/pakHhcBsVlGRcx3uSZna9JZhhEgNxBAKMEZRXJInTC
cb5GUsiRN3b8RAlzbSI2f/EI03vBkaUVR2lt4WE09EcFxM4bRJIdp8GUPzto/KI0tTHvutV1yvNJ
IG33VUvdyHYUKhlH3TQSGA5YBEg2mGwkbOdf+C2f2M6veBmnqqi1158bNisUt4dfCwALHY7qfizi
kzyMUvZVLEbLqIKjRTLAGj5r1ZIlSFCcOm3SKbFqy3clG4mBIU2tnNJ8A9cwVDs28nlGn9m8+2z1
Fcbn3IbVLc5wx/pJyGvfKc0mtloZSIRB2qqeNxQiWdJIdyHmLXT5opyLjOtzJGvI9XoxS3xG4a57
y7CryT4fRWUJFjBdMXta/R27S82fD9TRBijuxAmik6kNznSiFfiJ+Cp5udLxMGrHOViGO3e1K8VQ
pTCTftg6uESCBatbrYIAOLOAN01zW7UEa/RnwYIcorcxN0CXTRL4Hdg6aHKP0wYun2n08pKzUpqp
P8XQ3+AUhCPP2kAfA8OLSAVyGrI+hJILHlVaZ3F8Tq3tBbGKJMLtMuWgesqpatfTKnvBt1xZEJW2
c/XCXFvJhxxK86BqP6lvYaSEytWTNY8ZLhBFUu7Mj7OcjnTLFEyqVT7AEkqLy9jTMVW3jXxaCKdU
wWafqG8NTHN/0HH0k7pYYx+E8XGDcfYbnq69ORsLlUf3sVtE3CIaW/uDyTPHzKWJQMLlVbijes+L
XwYUbhdZdzGrM0tTeYYfuYMMrEQSKQEeXu8xj+6UZ8x2Jli4THzIewXWpj8L2Isvir6XTeDXx9tV
wzjNnteCtxTXxIbjVGcjPXMSxI3deJqyKNR0EuZRbGFhwykSMHA9n7FpnQyIOwxNWl7IHlzgllci
ldrorlLJMA6AUFAEwF23D4OGcYkvckrlEtYhehGoxdeSPAX2UwH151estkTIcwZKeroHYoZNSQTB
IepBQn8tNPp9BwwJQnUKvHHpYb6lgPnE6VWCdpxVq1UsrhinvDY/6tdYlc8hsVv0qNP4Otz9ePEh
Fb3OPI2XZwT1uGRp53pfKmhXAWTnQtvHEuKABn0ZZa4PUzAt9x3+AMjvBWbJnHle/ppFEiMxQLmF
335oXtKfvyGjtuP3p5jwyDlr/rYtpWoqJML+ftL997/5Vz7m1FEXghIV9SaV7VvAixd4qp+v0W1o
26SQERKlR0yd+gEmUOtQjTBrRfJbA/7sG0YKmu7W8LKwcg14pJD/tErXHsu5kVEZO5t4P+XCXuFA
u7xI/BQY1eIhGdbRGH3VE9CjpHtdYoRIF9iZAenBpQ9Gm/9lrXTcfPsL2I7hXd/yNGDp9nfsES/i
dgJLJhOCYOQc4GrCtuLLkRPAr1vQDU6bS6F2r/3eN0mlYIc9Rk1GxqCK1FaO8xtM17D8naci8Zuf
ZRh2u6kWLChHY0qqnwrph+gFVEZfv6VKSGl3OUOkCSZWkWzCxDeAdBqQar6PuaOAb12yvkSSnsSk
t0YLp3lj+32jmYcq2sdHs1ppbmr1Ktj8m2CPh1y5FHxxLsLajL33p9XrCF7f0T1OtNptSsk9MkTV
xkJUbwqXbNpnByOmgfzufZRZyjAtbYL8JXQ938H+Dq1NT5gTvgYY8HdX/4TJ7Gzf+E+VBmXyTxiw
XaCsvtncL9PY3hk2dEpyLXBH74nqqM6TCsEQilhfYRZfuX5NL6O6zPfy5pelxX8rxizIqhUA2UNH
/mRGCT+esVwiyxNbZRrMtWMoUTSN0j7QcYV/fkpSz/VXax7YywT9KDoV+9iBRRTNZGOL1YeyLnBE
RyRugmptfDugsFlLJXpbEEJ2EQhXzowTSsEh3ffUoLsE/ZwClK/4jEozxSoiGbtDv7fZ7SQ7nQH2
MJT+9ZKaQ3m94v6NUrl884hEF/5YnbbTkPD5Rmm4c32tHExglRIPozpx6fxM1ocltx1Tkm45nR+/
MmyIvqU1GxNc9HNJq/c7udRUmbVYe5RkkeTHTpTqM3IW4nQQ7WAXvT1aPHuJHzUtpN4Zh7ru1X/v
XprVS2UO4gj21Zv/fAJ6Xv3+m3NlOLZ+bvJcIxxNPThf7zokTfPvaXyvelD99PX+vW3Gp+e1wdUA
9D/tsJHu9RGxTkWLeM9fuTpw/VFxI0nd8CkvIuUfTNXB79VsqPPexBa+Z+fOldSRi0SrO7k06j7M
P+NRBkkzpqtm2wtwuW3wpe80HvxSc4Uxgg/Fqd6J36CTynxageqmxELaE93OPnROMMbdBmK3EuKP
I6wRWHxBDcnIV4wX1DXazUu8AwgsJbcTWXkzR654XUl7ewZRHLk2ntaq+ZfiKc2CdpG5SkQ8wjM0
/hr3pQcV8rqbv4lUF//9OCHBTNboS95jUv7Opx1mesh9FEyqs0U50DqXdo+9let8F3XFWUhvfMdz
ULHIch3xbbfYGp1g4vDn0K3ORG0GWH2T2ZXjgjE4zYwq79DxjizsUU+Dp9v9V2plJ4vcfn8meXQG
VnVafOHAi5jaCuu6dQ5XRzkf5vvOlmd1jz1BqrRCpd9FoSjDVls5T1e/1egYDenJ8gwPoOHbzjlQ
O9+shoq+YYgJuY0RkSb14FZlu+M7OmmNWsXvzPVbEN5q5Q9rqetpe6X20eVdEf3x+uBSMvntmDa1
kWpv5wm1esGen5LGFKfMzKs7JaFR4vwfnC2m38cg7Y7N9ZRZeJachY+e+2+8ZHwQShq4pYI0TcvG
2qXXRuuY/97jT/sZ7WnxIW9ZaxJ4/NSud4ZpQMvzeaBsss4mRHAZV6yVJl+xcc7ojbNKkTDDwdef
yHQJfQugAlHaKBgM6x+AvgRSAEme8NCA3on0zutD/je6J0rT2MQVVcZ9bqH+H6AEKKGBLan10L9D
8eKZ33CrUdGKNux8QXCL6JLonCgp5RktmRVXpDIf787Kp0jvSYKUzfkbu2f2Woea7g+8B4hJDNlg
pvTXKkgE4v4lEO0igl5EOytV8AWgYWDgN3ADZDdECcwMM1hb9qXg4EFe2bcSoYpeXfJugvo8bUbq
ytbjzWVL733Kr9MWvlf0sHeCygWE3kC0Jry0BvT9H29c5a0nW90qR23jvBQAtPI5C3ly7ivFYQoN
N42+KP+OxrFnnMlJwGTA+6HAsPY207I7r/Au68kpNSginer0zlq9IRIPk64P2u2u1GrKQ0mHGZma
LVoeKNZ07TYEbNrUuK88AM2KeqKn7l3/rNsDgFm91AT2bm007qyg991YtONnKAIYacexbDXOdh8V
423t4K7L+8OYlE1sRmhxSUPW+FGr+vqUEjmhf/gFmwecnY7Ca6G3tMn5qzQzhDODBWbPM1iIGGlB
odqET5MJkew1v2J8KfA+OXt1C3lBuE+Iyu8Z9EWe/NcBsefKCwAGP5ycVdZqqQMisZiYYlDQa44E
nCMWjAbj4+1p6G5ajd2Ozq0eUoF6wZQEAfzhggalCCCIChECdLrlkr8xUHK2wdweU0c1SCkKAn4t
1zf7Tg++3jZ8O9m7blYpvBFAIVsoAYcz8d9xTqEOs0cXRGTeTAl8/UNuzO8dcBzRkRn1hhjuAyjH
ew+f3eK154je2Z7A2Lsa+ghMD3HpBZUvD2j9TXycdR1RN2ClyOuYGlGRpwmGQCusJeeWzIq+O4nI
5cXk7aV5nCoDD1/mYMKmbJxx6K+cTQ5jTxNPMbExG6J/+PPoKMvKsglFkFouGA143QVmWAeylGbp
bim0CZ0S0dThFt3XwLDqD79k7cBNbvw1+PEGVCwLqrajnv1uHaN/fqdB+v1qnKlhYW2ocmbAwvpR
t/0gAAK8ygi7SRoJO+UR2zD4fioozj/nzRafJymHATjxwwx/6CMwoIy+jfuBOuYnErEiGWv7qlrz
lsAupCtL6EEDf+x0MRxcdVolJ5aojqntv90M3vhvf+PrEWCC5oC2uWp1NGbb9asYzVkIwFxkstAd
DESnhdbVH6SR45+/VSASwGkVfA31KvLbHbkbkGJvELDv0PV4aK3Rc15dkmEGsOXHYTOGBVzpuT+q
Vz/aRL6CTUpR/zSlT4DCPXOanCkOqyIIaBKOnV7CBB2/8N2SQ9MIur0CEZgvwPttOSsXUJEUXp6o
RXoiTOja+Mzh4RtMW3uSrwNZDOMC9yzl9gHNuSt6Y29lVGm1aNa2FlBQNUQRD2u0amRqMTNGPeY3
tYDQ+52amoGu5KGPrKL18AVxBEGmUEZe66KNmFNuioAC7VoYoMlGunW8MGcWwfAKd7fCRicOTN5W
shDiaHaCpzJR0u0+dOaC+U85pyl3+VC2RbhhQwdvAWtdHcAxeSoXckW0GmKI2aBF040nc0u6A59T
apKepUWFdQKb1Xo7Q3oojVVa/7kF7kwt6md2HvlmiAthcN2Df2diCRGAilhQ7ybrWDnmhZA6+4Ly
2wiO9LmioY4NihTyyzVZQguFhXyxv/zdolGgOe0m6Khmot2Brh81iik31M/NX5ddJPfYfO19p+Qp
NELIHjPg3k4iOs/um1X7fkqsYI7iSVxxzXlTCGOLyEHFw1O/aIdyvzBO12Vhf28xop4hO/XE9XqB
hPZouhPh6TrBehjky1YA4S1LIU7Xs20ItvMXgpDtbkP6ycnwjFvhQ/qd5+cp/rNofbyuY1+FtWQa
gA2adM0ZRbjS2nPFuiDXDIx4b2MP9FQZXz3q53fWqwBY+lHvkhlye1rqkiAnFs5q/OjiG5+8xbCl
IWau/zMeVi1cFdgotx+1S43mG/D3daavqVlMwCvuTMb11ZSMbFoCjT6RnJUDXLzyHADD0rN0nGW4
z/q9T0ohR/DUdS1BPNvpYCITv+7X3dY0iUFVRBXKgVg4anSPqyf2Er16+B/6fh3ho3dhYPHs9rUM
FVI0NoIbnKXxkTlpJj2m3TAadFTg2B75SSYH9x+Mpyi+qSZtId4pqVltmkhVaIr7PP0/pih9sXF+
n9TsD78rx6LfDe/TIClQ0T9pHitsD0IJUQJu2w+7xSP2kKmvOoBoXRErX/3yl6pSeYSBn3Vfj1Xa
bhpGPORPIxDAMo4Uha14fW7ZNOoGrBjXNoa/lHuypf+hlc2Qf8Qv2aCtdOoICemelNo5T6O906o9
WXBRnbEEkMXOBGlt0HR1Ck5PQyNc1j4QAEAfGOnJmdTe/kTx6vaGjL/FfEcApJjs6gNLVqvo4dN2
j0QzApAKU3BY7kOKkgLVaWoyeBXJWg0f0MJ2/SQoM46+7XT07ARr7mhE9ruyzbP8hV8fMH5c/qyG
xmarNLFh10jSX2KfcinK841+4mGElowM63KwZaLT4SmmwxP3eGY87wpVaQO1XcpU6y6hCbJfHags
j4Q55bgSxWcH+DOjuR824P+AGtlEMvqde7FcI1VXQ93SWOZyzmMuBwxtCXZGdnPq4j+WiJCpX8eO
C80GdTDHKK2nag+7FRnfkN64GuB2fSo3K8b2MP2vbVWVMPXmoF3UCYq/nevFY+81So7WXQ6aZQmo
wsJ2NePVrVlJgEAmmisxLPu7tetF3ivkLf3u+PZGtqt/oqPpE1B5dnfl2K6UHp23WeO2+fJXNa/o
qInGa2bvc8L+Aq630NGMGs8fexHJvKMUoMixURrLBmXrRDLQDshx37Kr3P0bu3xC4uIv1nLVHZFb
igt+UrF35zGRkBEoUjXSz4Iper27dw65i4KKWuCtS/l3I23w1tMIo7xQFAOseUMRX3dqOVLv8Ogv
hdym0tg8YgMP7xImb+XJWJ2bm/QBH5VQey9hP19FBSSEQh5Eve/THUFbDKoTHQ7/h/shbt/K9+7J
9TRldu4MKoF190W7i2t7atLsDnafKAS/f9sqGEfw8Vk0S0CvYbz04MFrzlnbi1YcJfWLChfgsyaM
BViaTBJTonZihq89FJ7XQLCu0zGZwle4FxgtSp0sF94/VdSkk6FsIb9a3go6JpEk6YS97bDF51oM
g39+S8eyrL8GoQSpEOQgDaJjnE4uHit2CPFQpvds8nvxnmr/EK+eIMKFVamp4FHRvmXuoic0HDRe
9Ub5ma+WyXXSwDe42B/GJc6J2MFh+jzyBxU4wGq++Tuaj2f4tPf/jYX5irUPB51d/kam2i8fZwJV
Oruo0NYYllDQGhvJF7qCIKyg/5Y/pvQHIRB3GdqZirf91dMPKjEwOkBQN98hXc9xP2eDhQ/P1/81
3HGWIBCp3ge3neit1+qj6+I3jkfPJSy+t+vJdzO3zV/leB6Kuc2aVEBVpTAXXWMRhRWc1/ltJCRI
j6IiR1yFL9Mmerv7O98pyKtf4FXSXCeYQkgcCx4a8s0TdJbiWYsNBf/NE+h0SzlavH2uGE4mMwLB
vzizqnHi6fW4CGn2Vt1ZfpEB7sVgJxab5yjvjf4gXxj8ULUNwrbNovPCUwHRgqsF0HC4G++xrFV/
Qv/jqJ/CI6oXBdCGr8JxMdsO3zaJUHf6mlYqrbSI3vn+BHPl7P6qJXFePvh6o79/0Y+Y2ieGcXnP
x5MU2wTXmFE+jCGJC0prpV7mQOHPIRmmkS8XLiHQ6gnGgDwmFNIUds+IV2attoiurOsxRzJglZt8
2r29Xn5pYIkRlHcqQZklfhd275xITeBi9711eXyxv0nulshmZCZniGY0d1Ny1YopqmedIgZnV8Q1
MtsSFhQFJDnm6goyQjvkuhU+VYpDswZeJM5Etj8bcUVNokminltoE+28sZBxtyyt9R1yEUXEeZ/P
AY/k78rk1pTe2ecv7RwwL+uwaHHUnh/Q3TU/7WLXji7nNb7adZ++HO5qVkcqNXa9n3hP0Jsup1kN
qhaZluMN34SNdftFoBzKQmNnsisVFOJxuWC0yFGTPYuGSy6iTvQH+Y26+/3h2NIE9f+306pFzQ+C
QAdo4dhNP1rH0csHkVXl6mdp78WzrqKGz1PhnwZvVhAirTWOBY+vf9xs/iWOnAICe8mckqDNDGG3
1VeoZDCPHwSt3Xy5V7rme0qokvv73fPxhKCFvpKKz7JQs1jsA5ycEaPPV1hOIgUGwkAYLXDyLUNk
SP6tcsdcC/A57SPJjLM8IC/DaukGF+T0WJmebB8t6WXflT8wLHLiYMxYVcf85m57s4BXy0/j+nbF
82JZZ+wkTZCvg4UjYkCwBALowmIq0Io5ffs66Ezg2ypaAzqlHOWWBUbLvw9+BSXSiAxVflZzJhu0
D0uqJPGytBchXP9TIhqJNAbN9lE3J2ZuV34XmiwLSlFdZZCF5yeAZUqL7uQimjMCoE38caKbi4bJ
+OAkVgGHEfFLv2iZp09i9t5ZPI9gOTNAxgrRLieQrCQRKrlvVJFVS1PZa72QfdxnGnTDTrjvJA41
uqIX7D0fiK3YW5AgjeMeAIjRogcQP1K3zjmvtEWKYqP7Y4DOmilM2WyRfyQsKpc20kkkweQVFzLY
95nlEjjis+z+ihXn9NEfZjGB3FctIDn/jOY4HDCQIRRlq1lHpH7g7yjVGRh6tIU0zw2ASrnwHyad
3PgkiItT5nNX+Wwy/6uqWl5cFTC0glMN2s1fvFmPwJLBCBTSIfmL0SJRBTqPytXDkiFsf5G45ger
1s6J//1cpibgRIg0dHkoy+Du0YyG5+65E9uQ26TM6GCHQrdTvwNahXGuzmS9sId8cioba4bv3IrO
9B8DOVQ87LclmgxYLlH41x/c5WmiM9VUTAhyEiYmziq9HhujjhGCYG04IFPmGTwrAkatmLhnBkB5
B84xq/XVhYnh8Yhf5CfUOYdDkPVWtsUnypVAsFsHHEGaqV/cwvyZvr5trB4nZ6bFa2ay1Kigj5/3
41P6rNVcOMmv45rVBurkxGP+plRGGa3Ge7hmsYp7vqaZYQvQaZF3u1F1z/gOTZWdfdYbOdrnev7T
jxJTncHQZGqfZ0v+799pJe2mSpn3yR273lQfgm0LKLITkZemModGdF3626ZJawmZ89ocYzGs2z4o
u97LwvPEKs5zIySfrgxI4sKyV24ezg/51sK5H2eTsKguGlVQnfTx7LGXC3Evo50aYmj2zzmF1DpP
jv7X23RZ4vxBTH9HHdofmgVraHCCqazIcIKUK/JSAn+LRHcmjJUpUjfboEFRTNAcnpbRBf+dyECz
/WpGNpXlyfP6rdD3aMwc+dRkuHtJC4zd4LdqIviStpr7rltqeQWFiFmygG/fggzDp6brnwaqdA2f
CbbZkIOsBpQCrGP7NcRZnkf4O7nXMKW6tEBokzCEHOQifRMggDYZsWEpRCsUCAXCCAPV1ewmVdMg
54FBA5unhZbeAwaoKriftrGuFLZs68vZpAHNElnD7FMizVsAUZpbPKINadqRUF0oYnui4jGxBhkG
89z+KpSGDiLx28wexdmjmb4Oub4YhsjYgObws/hdpxyPJ5VgaaZBxtvqh6brKKf/6yLvWXYkukgf
btEZ3J5QJbnwpTYKqO2rlFBRHHqnyX4yJSfTM5ceEng5lin3llAB9/LgjrIRDh/3fh66/05EIAPR
8ilOP5hlphOGEhKrYQaz8Dxj0arV8Kc86HwxPlvStgExx18IybwtvWqerSwuVX5ok9KHwIoxFpxH
67NMclQXNSYljfHm7wyXKNToOQRzjcKpEZYzPZ2JyFg574iWg76boxeFv6lUq9N0F5iJcJwa1kg5
zvUyOpbeSfdY3O5AQcV7D6KW5F6OZ/9WSUl1BLmJ0ezvxT4Xt6yOy/ZNsoR+HjZ4gZ20Ul8cdt5D
DFqCX0GZz8rj+99WcrchoYDQvwArg/ZtYg0SSfJGc9Byebn+yIxnWDG/8dWxVe4W+k/Et5d5S79u
KS79/+YwA7dyARMUJ6CLfRLGDQJMrhscCakCCItguKaudJqHAoFTGVRFIKD4KqdidL412ZJu3DxJ
CNpiz3WYoNm5uDwSPfK5NV9W/KlLAXG8235YvgDjMpFS6KRqR/L2Ez1sF2/6XXztqq2Ao38brgrl
BjtCuj7TiplVak9p4+ZyitDcdKAgJYc3JTMTfR4o+HcTlSSf7m+gj7f3LEsOTAvUQhQ3xuCV6+yj
Atj46/inpuD5V6XjlYd/RtmjnzeTCFRfuohqtPKRGVN+aVHQrINRKg9wfDFgqtaR1EKYrigO2X+P
7l1QgXQbfxtS9PX2+UfcuC4tYuHFf2bZQMxfM4RgrEPQPpFjHbJzrWjnbVYafaojBtVOTc27gup2
k7OMdj/IGHS1PAoFS4WfbJ5X+YcxwADGwDN8StI78OniyQDv+VA6VUQd/hx5J+v2oVATj6YpxQn7
sZFUNSU+5xFrgfsI30saWYFn3YfpMSBqP6asiAwvu9mNtk7RJufmltySwNJgOIUCrQHhfGY7dvIr
h7yb0XwqMrmXPe7Mu4NwEMkaOHl+pWK5OUROZeN6/Iumayv/0axNOTB+Xslw12TlqTdD653t3Rw7
AekfwUTPSxH9SDv+u/xd4ptA6MVt40zy8BTBSMPQYjfMDo6T51OHyOBZOe3Xec8agnj+AbkjZCEi
ypEreyN993p/X41+PAM5COb7wqufUziPtJpOITmKqD64eaUC7zjqDOUZH9+uVhyaMSGjRiIBNQ0W
mJDjtbvxkSrum3CX3SHdn/7GRXHR1as2legoJg+U1BCWvnTYGyIgryII40tBs1gec78WtvvX/ReR
YLYhjlRnZ/qAv3TxiUfATUGhc3/rBsfgFiyJ6mSImG0tg8rZ30Z807/56HRBo6OYvbZlTFVsdLFr
ZsAgMUW0KqyfDedIaJh5SyARXkbS34xWakIJS7Cc9vr2RCwXne6jvDVk/wnXWGALqEDN5qBgKCrA
RueuArI9FXq9Px2XD9bzwLSxQXo+Uf3iiN35q/lPCPTxE+E9CXYOBdu2ZNbmQB9C/Ae8eQWGQjrD
my61Vlag+QjI5IETDcS9Vnx73/H+omRvNoT2/szedpUCWOjEIp0gqlJBjbMbV2g9GRX9FkaOnFtr
1w3jF2/6LbzIi8Nc/gO+DTZOVv5M1VeCHRRy0FPWQTFkxIKbbDeSJnaHh/jp10O52IK9fNpJlaKc
4TzWxphScYwKma29PvhCaEZcgI2TBkuJFFwXw0uIj9+hKOZjm7yZyJ+UaxD9CTLsMNKxS19YPxwb
OJM2MXRt2c2RAzl3MGeY7eb+Y8lE9/Q1+MQhFvlAPBI0XQH9Lswpqo7Jr+dpZM3NRYkj9O+H1zbP
iMxvEOidXPamsESED3Mtyy/nLVNLOwQPMtgf7LT8sQrhyEK+UNRDeHscAThKi2XASYFOjsBIFxsY
pwozXE51j5rXdvxyxe2K3bhOF3DaQmxb3BryOIO7HILF4a3nGGsHb8eukqVC+VvfFMJFXNkiqge0
S54kI64BH7FT5Asv78NmEttjlk+n+cxyvbGnrTFFAFBjnR4RJWJRBBJyR/09vL21q09TNLK/0I6L
VRTqE/Nmx8XdIpyboRXAafxE/GLudKwxDhtCITwcCCPLZwQ/RRIk9ra63TM7peCdLSRdFQ9fVzZu
w5Wih41I61K0h7d8OhzQ62u8MEAnLum0zcCjokTc6PrU4H2yEkmiiTNFi6aw0mRDpesg6tZD8W9T
AHuBY5tumRexMwYyhQEB7kF3RgmIvuNSiMw6fjIi/aJuE+cROxTXf22mjugA2glbuDYB8CaIlvOS
YyNEfnk1PYWLhtcs5tUQefQpzRF0fS70uW+AaEdl/cq0h/Zuh2r2zsC02KxPiPJtFVKpkdt3yjVv
zzCMg/e0oF2aB24m/IpOmRMmXqdQ90I8cCDjNoD7MIEbbatLFt3fN+TlD4VACbEeEt+AMESMTY1Y
GZRw1DMTjg/gkxb8l/hAIQTFl3hCUlFcTQYF/r02gnXJpB172VOBFp9E2mlVyolaIlAlT6lBkNya
AJgO8ch3xLU1HfQms5m0d9d+ZN68nUM8lxWMLEy5TsLR2wYZp4tISTbi4+9tps3NXDeGj3fMGB9i
phe0/1ROCE5xZNcBQmOUQ/fjOt0rbqudftapHugnPJviBC4+VrweHzDZlC+a3KO+FuTZBX/oUdM6
5nir+Xs2OfN2Bm4dzzBqL4zpuhKtIWWA+rRlxAF7p3xsB94nlDyklC9X1QmBBdgLtBPTq9r7uvu1
CgAxUTjq+EM1BdPd+A2VhtePEK2igXWYAifFfD5tqn5YkuU4nCctYrR3DffuyIYb65+6pHbSDk4Q
HTFZiSFYjdLgQfkPp3xrggX3QDg0vtNCf9Yu92r25jVFpWjCVTu+5EVg4voeK4TLo+jRvJWa1H50
EOZbACLStKH6T7HX6pGJPnHNDzrrYeSLOpIl1GEUkkTDuFqqjDtZqrRAL7tURLOpeVRg5uyI30vo
KmJRSe2aXjNREMsJao7RxJaxluXi2kALYWAKX/ussBpfA3n8pwoXCzrjBqdhfOtFECLryNpvCbat
YAkB1iUA4Syo5gfYv7XyTG4YZpT6F+LcDayJkBKF50Bl8PbdaZ4+vxcbVB7tN4mtZ/SY9PwpfJ7V
CNygu7BqPldFjvey2IKW+JnHLTIoeFPAG09k/TShgpN+UCUyYoH/MhB4qvBjNEAhfvJXKtFvyfDu
vHWA+vJfTVtQ8ULzQAh9iDZzrpieQgvdrZm/h1hcXWgnCXzXCs17Cdjpybj8fG+HW24yHxaPGlxk
SryOIPqKeqC59q3+WzmsOuPo1QB+MKN+QF0qa1ieINe8/leybseQo1Us9GY9hkuUZDTMYm/4MUGz
M8JxH+CybmjZSNzMCh0IVaQ/1ZQYDwVNqkPTP/Pq1w5uzAe3Olsuk9h6zOKVvosYp/lJ1Qhjqnn+
LCjzQj/VloKx9poxxWP49b6WeCeGSexkj4UWBdnzOSO7nIj1moiTKUtW1DKH0CJRS9MT7moEBqva
q0/smfgS2XZjnjiYtDb829BmoTdMxvwvQ7bhWN1eQNXaMWyLigbfKjUS+nl4U8z/NfPFNHa9aFp1
UKIxNipZRhVdy9VsotYpnhcZpw9XMs25g8XyQy6zSLX50V6IJwnmIjzQY9JbnbK0Y5fRXeJfcWi/
4+Mr0mlVsG3NG1eNNTQvSpL4kpwnDLawuAGqn/PGO/bb0Y65EZW6Ya6/DWK8VbM02ROCTD1UFjZI
fp54Lh0PPe2yyPW1fN65zsQg8m7raeKwPmGTs4c9jQ+2CsOnGe4VoqpSf15xYXQkd1DFJelhd7YX
d76Ic9wrRsON/Vya1jduk9nPxWCJqRL7Ozfc9dtwqIvpm5+VhMnapFLdCBj6LBNBQCKcFDaYd7o5
DD60L0+YeW9O+WvCr5hJFW5JN7kXT54MdUzf2hrYQtMpc2i9fEXfglMqq9HsHI/aNpuDY3kxKWNl
tWae/VM5/rIHqE7x9cZJ62Ix3ZboolDAJ3nqUTGGMCT2QoRywdh+hiVg0wNWTFAJxLzyH6H+iCjf
eBhC+q4qn2JoH7vRBgsQBVR6Z8hZBqYsEaC7Xi9wBdeyYsJD36pO3kpS15j7kIZOfbpLfw9wNkDm
Ylz+yrgh3e+Sa/G4xknlyS7WDVM6U8VqPfPfRDdtWI5xovEs9sQ+xFPiE7m0pT9WSGrhYH4gSHUJ
lMwYdefeDEIEu/DQuFN1itgz1wGmWWbKPp09dkYjZw1KnkFU3FELuhLGzgy2Uc817kz0DLI1J/KF
BM6Ns916PBly2JAdeE+skIajGCYVAqACRxhUqEkRoOpo/YFqK6UEY+T0ARk1DNkxavXAOLHCFeRN
DGDTwr9z/PJ0/eg1DH6EynxbjdVqy2JyKnIvboyHxqWx0bH/aKZEwZLO6VP/GMISjAQaw1y8nD9q
gy5V4bjHBz63H0hjE8IghOzFAoldrKMkSMTpngasOffloc6m7G8kRYUalFST9ZJrOxBdJoRAXdb8
VUS2IoledEjl1F2QRpxU07mBAOTD/mnB3rTchlNPKRl4YclkX6Wtntrtpb+NqECrUuenkKRg1lir
+wySUqRBBRsLkgy6LYkrIq23vtsMdHY4aFoZ4llUND5g+WV9mOPYoN0Zn7fPNN8ahh/SjhE7WQRi
bfpv/i+deQKNoA3+b5i6teBTlw5Q0Uw4LXeOqLH0TinkxEIX/XcR6PtHyiB8ygVMzbYBjVjIR77S
S8JjzfXxGMXTO90qoYsod20bSmgXkW1jEYzug/4D/3fWVEaBvnQT+ZCu5kGkO+ndDsrejwRu0O+f
LIir5R1QrHy2IVbI4kOBYrVZg4wg8Z3+ySlJ2drkKUFeY2BaAr9BqZ72BtgNQPYlewHmKqjSFtEK
jre/AQtjmDN29A2tH9B/j2shIE4C3ufm7xVgvkcU6M4jnTZrZmUhKFu0+5NfIm6Jebxg7YM93Tv0
qDz4qBQFbSnKSrQg9k+Vxzq6Jhg2VEMFQqo84xJ49GJgec1jZn7xNJn+XUqdb1ibDcpVTNorTkeP
VtE3cnmH7CUAWW3A4mowdUFQuFmANTcVxPflz02F8eseWiaO6unh72fDujxC1gUzvqAdhK2izab9
v/rsoWoandshUG7Cu+3/gPCdvmqGeJxO78MxY2oO3SWD93Ym8BRAVAQ6kd4ye3mZlPIq23oE//C2
5W5iZlcGjl+vtwfuU4MgBdWkkd3HorpzQQTECqVfTM8IXGF2A2p3OY/mQpcYZCMl0eyeNQvmgRxd
eQiTV19AmiX7fTr2KYIoDBwVkKe1tF4gbv7AD3iYLeX0D8/0bIYN3ghE50a7RfTwxKZ4bYn3fZsD
afe39In1QbC49cGlJbazdG3IEki9cHF1dizDPAYAv3I5AUt1dQ5NA//N7LV+OvRrcu8WgEq41IKU
9n/eUakR9q/8M6S6W1lXYQooue2P4s5op23mxWW57AWfe61mW3blolNXZ0WFHW1Z5Y+Ogq8aUg5L
QfTpK5zFApL13pyc/BDyU7JSE/2yam66oyQR3LCkyg5g5G3tDCN3Jqja5F0OFGQGS2rAnSjoe6Wm
zmTsaLEh0396CYwx4l2ekNUgZ6yHnyjk9ElT3Dh6rqaES1PcpFHeplKNLm0VkGSV2ZguohjhpODy
t/Bgx8GZtCwx2s7QOr+dt+LgDe4R84bwLpjWxNvG0ur6ShQWpAsZioft36RmrqKpdxYPxJ+3cks3
bf2dWF6ke9VKwgUfTX+R48BVf0ro8FI6+h1s0+kl+v51OqhsZz1dskhtfYnbS0vwF/petVxY+p23
aSs2pY1+28JDcRY3Ab77GtxjrmFovqezTz0ZDH0wyxigVGmOk1Rrvwbh5qzLQUQbXU3mOamxFvoC
ITIyt9loBuKD3vH74AzGAvvVsL8cdNjg9/MV1rz2oAxotUQWgjIb60V5FQ20I1gHee6uOdAoa7Q4
NK8ZuZ6gw3071HeaFkSCY3oaaLwz1/wU3FJmg4oHUQlbfHwHFPFYdwtwmz/Ss20etayBHoG9r8gh
IHkPkHBMD3Nkh/yWjHCOyM2tayglp1F8IR8XtbUW6fCkQH6kW5unzTUnwMicif6ZCjwl/Ous5+uq
JSAEl1d6Fp5Cb3lOv7t2V90oa4N2cFXP59cJQ1MPwSirp9zfjapmw5ogldIFzKwoqWCbwqxLjTQ3
gWmP6mlq/8cCekEvE0Mr1bNPe5ZU8mMQWYxGuO+0lI5ZPpks1PJlvOyhdgP4qzEWD5vrpLd4DFiT
6a6LoUat+4dLL74hji5/SGwamHzivqympMolNIfx2UDCVcTObpAwBRvnGbu8/P+ZBUMt+ooobxxy
gP8S4D7tHPUMP7Vrv91Z91KKHUbsSmnjIsF26mAHAAKx6TpZbvpXDKIYVEigUEY99kyBbTBKIytu
4WvmMDuNv9Xy6gscCvlJxE4mDft+XEuWiUIDq17FC9uqYghSqgmnla6M3e3Fr9LxBSLBPXFl4ccs
6ITK2rG5B2DFGb7r9oz/iMtWCUV2SR/1f4cmGLYj+Iceu+8LmfbJfG2Tl6mO50AW+TJlNbM0//C0
HwfGhvw92be/OSx1czbkdal6orCf5Wya7Io7gamHouunbEcas4NsGa6Ks9UCqh5mTNHcWnpWb1Jx
NLq6EpYC91i5oPcvbCEcFve/GzpvXEbAvuHV4F/zpS4/VfxAwyp8jHamQ1pCMqepVNaoCn2eG/9+
sRhjbMH1b75B7CExlB3QpJniCpM/w46YYXUaYCfzKU0odIAe5EM8KS8Zx0SUjD3EYeRup/FEnYgm
kym9ehucn6yRtg+A6oUmv9lExsgB2mlNS3Wo1TF+Zdr8s+LcLxem6HTTgCsaz/DENgaodX/+a4tR
wHzoZd5Z8EpqBu3TchE3gZcVUIHIniZ3mfdhO+o+IOzQPbxzu+7cryDGKADSJ2hvq/w7B2jaq/J7
fVLyO2XbLtT7/s6sDgn58cIOvy05NxcRcGpIZcfMoXJw9CsYYb/AQcsZVGHVnqebFzeUx5lAX4v7
SVW4KSY2c2C9qJ84ec3tk0EihbBd/JnDNtQd8Jp8CUnFT46YIENNL4KXST9fZQGbHkS0s0C7NHhb
0efXhZOOqMhQcv55ygf2iD34OdAtiqrFI6+0n6dhtAFXHkLJw2ohXdei3xrUEoknW0YXExHw5W91
c533tzzKNO5D6EPvDFsNRZ04fw/y8e6vu64PzWX7nLE6ZmM0Qvf0WBAJAzIPjpKDuamH6UVv8XAZ
OM2BDOZ8ArgPvR1j7XSpqluCGyw6p8k5C74cKw/ppQcdmtXP0ukrJ9wr8tBLYRm/S4Vew6WGgib2
8Cdr1zIH0+cMG/Hr8fN6pWDlnzndcA/Lu/cqHZrkLnB3VFp0KfCN9h25rKBMd2CQtub47uRmDNh/
o5xQSpAm/UGScaa6/m1QI4huz69heAlgzdgynzvsE3mssNxXDBeUoia2RUwUNAM0YUo3J7oWiyy3
LeMo6+YV7IneNkDU5Bwn/8cizZujbnrmS1b7ySi+pSkHFn0grTpGwUqWc5SdgYR+MEp1SRHoy6mT
gsEIICzCJKhg5JjwWr9c6GyqxBAZZEoABkovUFEUJYXuaJ2UdtKvjL5xc1vFCbNoxDvMFqlqPPHe
SXbe9LKDg8Lzrp8swFqaNtiv45ChSzIVP9cQ8bjhcoZADpINATgerhbE+LnNITrD3M6AQcB6uqcC
/1euizp5aW846raOYiE9Sxny+hVeKJXxrc+EUnHoklo5NerBxK4ZZGrFWLzIzOkRgTrqFMJ+lK+h
0NZYIk/wKLRtQcgyMCLZFz0Xh0ylUbGC9UJTqEimjxHGEAixoGWZ1zyKeEj0G2ewlkf2/n5uZy7B
azhpU4MAUnlkMT+Sm5qteHMrV50HWbNRkyCkYDIFNV0oh/GziAD1vH+M5HzTnByBsdmof/kOyxcB
pVS2Jaljr8jGhZ33LYNWvMbcQ1byHw1sTtSIsZZJ1gQOemen7aLV32NuEAMJc3TUll6q2xoTyaj4
J96tQjxxIHtcZlPIdB928W53CNT6A7FxXYG3KAzQoE6owqVdk649xjl1P1nVs+GYkRVArNitQ+lW
VWh2QsOfo3KRk6rVh5jY+EUE4Dl8BQHwCPlHXT1+mJlXsTanokKAvnmg9Y1JHmGkoCjNMUqfW4Dv
MoudbITyVpTSNjutOukb75sUeUCuWHkVed4ihLvxG8oyI1y6mujc0JNd0i04nrx35pQ3UTBTFomY
ESruc4WxNbCP1kimzlfHGl1pxJHnBLSDVzCGaPp0mmGC/ig49t3qo6kWyjuVH7AJ9F+1E8ObCh2i
2RNA+HXHmVUZTuxXtfp08VBWDIl3OlUdHre8w+Z1rtC5Y3J+Vz89AHpFDwBwKs50+aF5DlFCnI/g
VLLLKGltcEgTpSnR4gvOn6R+3zzLhoa3nYiiJifWE8/0VbUzlHYauy3V1rb6NX96Wy8a7hZELHLM
Upit2fC/RLVdELNTwdaxDU3tBEkSqSLG08652aoJrkbyF+bSn3jacMeOG9K0Pj9KFgOaRahVXV3d
Z6BtIGyrKsqg/Tiv42ioaXfaAnM9Wg/UJU5whMXUXN0bAkjOAc0C2Wi9CNF524ppEdBY2OyOnupS
Rr1SpNJ32g7rqxhwetYNtRuOBm6IM7HIoxjzdthNnJ9USNQjy83lHNVVCEXxEZW137DMjmeIWXMf
UBNy9Y39dcvxa8bBI7TozLgZ0qbjW7MW0T2O7AL997aLFQ3+io4KHDxkr+TEw0PReaG3KOCixk4s
6PuvQqEoEJs2LzUc3pYxuopQBCiBn0gXeyM7Rl+Bq8P+OSQLuHiTMQV6jWdxAiA/3Ulf+5Zybvw1
jt7JOiYHBtPjzZ2Jao5INqIGjbVPyoh5jRtMWR+P7E6ooQkqKOctkV8ROTajdaQKcZ9N+DHsHcTW
j0FGw1NZ+T8x/3kpTlMGTwwY4Evu+uUMlkSz8naIBzjYMyniPuaSchBMwPziJo3Sh8B03x71rPDo
MEvxoOcwV+ZSMuKUPvPcEny9S4/lI7BUpvgk6X2uYnVUeqLbOhgmkJi32wFsPQ5Li7muU7ZRv6K+
D+FIaXgKfXlqN3PXTNURXyomfQ2WKPNISLQnsbLIu6TwsmWKCuOEBdgPR8fzHlGmiLsUQLM04iyi
Sl0xW3hJZDXRfDKKJYVb2owV6dSFV1EaAq6TcdZLXcazh9VykB+VwdrEEm5U7OHuss3yl74tz+V3
0TEM4yZvq29R+0A6kzbsBWy6ZOjDngG7ZoFUN5jgOfrKzwasuoeWkR+UoX7VhDQM5rWj2heNayZc
k11Du6JIxMDJNzFvI/8nVYY3aGoW9Dix+Hf9bmvut5+vdM80TKrlrcXpAKQcL5TqdIx40RyiUw4x
d5PprcLDIy96Xt/2YpYEpkRauY4p9C+sK6ok/P8YkhwUD5SGw4CPm/2Wn1yASzKrHzBeSZ7hcCcK
cyB1zGybrfzopkUJB8jveb0SgvvHWrrv+A3Y77BRIbqypQGLw4/scdV7Zb18nPHOpT6+4HcO5TNH
iuc4nLL0dx8F6/iKdh68mAXsEZqJKqxetr3VY8ws6CD0a9eQj5qYO1rXQZmbNgJgP168dtsRNklX
96EnMEAzbn/H6rpSQKfvqDK8AS/6hPH9zM3cWG+tL2LfCVInTdhoBr/w5m4t+LYq/k9leqLa78gF
ZH0si23T5tH89/XC95CwUOkLjYC5U09KTG7FwdawTdmBpW13GfhvLCOZy7PmDPiwn9vurmb9Smcm
gBM1qtKc7Pbe4OByu/FAb/ANych8xwrIQVU83zHxNRJJt4/7HzBllz0+RzR/etM8/7B8mpBRpd1l
IkE623rlBOmlW5qyBGm2WmFCs5naMdPklt+JuioE3ldVjw9DFn/OaSzuqwpjkbNGvnGDRZO3TczF
xhTp5BDEacezJxq5Xto+cTaxzdPxXE7ibgUeWr/rI6O3KgiNHFrzF60ubzbmfzzrANmgbUBOtWok
h7+j11DFF04WsN5fs1P0R0/Zbz1mtoDlj+O2rbyoftJaC3jtnXgKsTxRWu+x6Pq37a2xkJff3LIh
at0FBdxtpOTecZerdfC/Bj08qAmJiMKDPSonteK7p6jqb/XkAorH3Sg/6ipDaS8wBYq7IZtdoihx
XFVeOpttZ7yiRMNwXcmQD9dua/m3ELqk0M8uhEQuwG2dueXdjVDv+a4SlJIhGWm5ZvwKgFw8xplv
Fk1jbbN+0yRlvPDysmr7sH3yJXGvQPtAUbJleF8m9yRLdrh8TqPVGZ4RX4xmaIQgDSyYfhjgTvkn
jTUaMvgm7OF20VlTAFzhErySoowS8BFLCb634NMh2+FMSOdHgdurlGz7H15Vrz+tYtT183zgxW3w
pN6J4XDdFR69CNXdTVDfG+w8qBT04bzowBRiMdwvOncXFcmv8zsymqk7oT47BdHyBm/qqOok5d3K
KlPd3FsWqZ8qO133kFxmJYJW8rwstpKRoSbugatNRCnBDyj1NtbhIEMCJNpmjHccNTHJzy0jUSeR
KtlIgKNIvfGsDluDNJc7VipWXl29LG0diuR7kMK8mtjkEkeG20mMYZBk6tKRChx8rKg0YCCMcuwr
7DGFKaBHm4fjGw6DVsnEv+0P5SHPGdwPktNOoL39fHXeVuIIzAEsrI+QZGPc7pkUkDdDqSiQU+VO
OHMI4PSsGMrYacojFaGOhxClBkC/IW/ttrMl2MsI5jopDZGNeXQWHUOEjPef3ah6AdCKTx7ZShvq
FNw3GGrL+Zi4zQZZ1/Ju3B/N6gXCAvYmgDnrEiIHaCpNxS+EyslNtkNobvF8+sDMC515z1DkwbSc
LohDUKasyl0gvUytHfrZzuYx58XcsH2YVo2I5ZyDbOwbJ7lQ547Ro18zIXGuz0EIdFWiIkI+3Kzx
GuDuGpxoi1X4ejT6eJ37G4h0JIU4u8LQV33TZ3ali2SPeuDPDgVQgPcoC6wHKmL+gnZ8UbXDxVcw
Zli0n8L22TPYEmKyehPXaix89XP9y16BmpY2ItxQo96IyQZUWdkV6zP3p6VrQLEeLJd/jEhW7ssl
LScH1s9/QGA5AccYHx2FU996eYk0ckvVPdaLv4ke8RFMQDFl6mtfxeZMYkwE/2J2wdbztEIaWkAX
mFajtnJS3imZIQqZox+Hi978BNUCRczCdHHA2qfDpoWLoHxmI42LlhFaV0r9HS07CpMZcGLPluf1
8px9huaeawyaxNG6+6Wg0kEnN7RRA/D8Jdqq9MJ/0jGSbMGUPJt91osh10ECOJeb66uHtbQzFfyS
ew4fHQ6Gys6GZWsBLFY7lrozOQO9IlOb8Wuf11Q+x2cK3o8SE5Vvdjn+cwCuKj/8ZHMusDmhWEwF
/NbbUR8XMI/mROra0EJimLFdtNx3rI70L3q/sjq7wB+zbAtDEoDFp7pgHLSPSF6C2GZpH8UAwZLP
kdROeloCKXnMWUp4/a+1JH23M3ZNwXAaPTVbJUpfKpI7or711jxEfiR9uYZpA5CBmfMDKw+DRUCm
KWii0qWL3V5GXmQTuNU06uovVZTfhPe122RetSnczDxJ8kdbq5JqTwV6+QnRY2K7wSG1uBocc+3I
pWZrjEBxFZYiJt9WyRUKHnABRDKHT9g34DpcXZt02TnL+a83Vi310yjjyh9zzIRzBKEcXmlltWg2
iFrCG4rXxVoiuJoFlo/LjqlZzewmb4xL+2qxG5ylXlMS9hQFShN+71BqM696ucrsduNUmAncVG9n
/KUei6Oy21HdK1NUwxDbGWkvXktSR7d4Vs234yAiRoD2J8t9Bg4sFHlHRdfb3p6WLfb7KpTKHEBm
LGTMq58HlOCxaay4XFxRLe/ueWMpSG3vbmMyTUVld8LLKR1A0Kt7e988gD88lB8TjOiMLPYlkqh6
9cBJkMEoIU5cJIJ0EhJXz9GstvyYHoYlmKO7uQ2TOSG74gfu6D0FbNUdrh1g9tbexf4f0X8qs3WN
EE4PMQj5zbYQIpcyJlEeYzBty9KRpdVu+nQBywnhMW3FdzB+6orAKohDejKNbzu9/UZLGjFfG0FK
Fa2H8lj+jHDWuusKCuq7VUO03qQvX6AO1mRw5LFBHXXxwdk5d7qWRj5VowNsZHDUe2wi613pcvbS
Yxdo4HrDXj1WMoYEqj7r1swMMH/RlmpJaVfeyv6u4MK4Otrydgnha/7XIpZaIJp7QXLheIh01lNW
Orm4bZ7pejoFOpZ/tnzp2eY5qfffLOq4zdcyozC8p186p2ri9sZHtJnHJ/hVlA3f27PSPN8cmtSi
rkj/0Hq93PZc2ZkoYP0n8HUK4H8m67JKif9METzeS5T2ScO7RJkSwWQrP9cs/5ZgtNwDq3B2fq/7
SBy5DNl+YEJjyDFDbHWCz4AAuVMlLgGldbCeZE0dzEpJ+W+w9PRtG/9hzJ9Pgk+Lvuu/75OpVR/4
9TnP3rqKaxLWXIcgWGEepB/0uCRALQLo8Rn4YoHVWA1pJIBxCY9sDJ2kHMvZH0kjnc86UYQP5CoU
2NTv9cXtFYuMU/gAUMxdLWXODG/p7EubD5Im+t2tQ8ZSuLa+twtJLw9XnBKZ6EeZ0Fc6+9qRR1Ka
SLMYq/+z+Bxfu9Tyh/NCgwv3GLTrHv9fGZA5bBVPNxW6DGTfYVTyjyU4jUmUvlUFb6x7seqjI4Vg
Vre5A6GXM872jsJ0bYMVd2GAGqtDCwBQfDhglUUoVHxbfdE2BV+bcBD68hBmmAIlq0bHqrQJTl11
hbW9Rco4Mtz9guUcb7oUhRZ4+gT4uVfTG2r8Eo63tm+XzHQ46jZwILavHlu1o2ZU1z23r3yQLqy5
Q1qK4H7cC48OIHHahv0TZzhI8voKmdMBR4t+fz0O8hp5LMcRvu+ggmBxjVybQ1UGbY9VTfW/lgf8
mpz2LEsy8PEgbn2Q0DMikW9sNgqQQPGHXj89r4omYEERliOGfw4CdhqW0nXzK0BDDkv/NNd95U0N
HARF4gzhGP9dq37bQPKTI2yS8kNivWwvyn6Dvy1OT7CXnC8lAjDb4ipaDG7qtA+i7SUsq1EGFIwS
hEgnc8yNrzvMRSnAetu5JinE2NHcpWwYMnaJ2F8BbzfJ1SEVs2BoccQBpdVOBW8KV5yxxF3o8Nmi
RFf1vNSS0so+kaP6MlXgXBB7syGAIK2suFTrVww3ZKxj/2NUs14p2uMa2NJw/+/bc0QvY7wl0zxA
PMcXN8CphNNt46lyYa2iSva33+w4WdXn7h736alkBiy3/3iseDAZqsZNEFvJgAdNGXxcw0xElx6q
nChYtKPjkNLVTUGIP1iy+RreB7eF5dvzU2UV27KVoWSwRDXW8/ANKHkBQClwVJ93MdM3GjOEz3Xu
j1rEQ2VkUpwFKwuVMBWLGvm+iLtjwlI7XE0vKGAXWOrLK+CNNZ1fJ6GEe+Mp3LY5dm5RM6o66ow3
zMp1QGJ36eihjIxUqTULeZ3RnPBWgUTyIGP+5xJozeKuhtx7kB5cOmMQHG+x3kMwXL6c6bUBmkjO
UxbgN0SCNwFqt+j6vGX7XEuXNtCPoLkIFp34nBx9eL6CAXioYy1GvU2k53q/7I2Ajh6Yz1nVkmEh
kmBzTtn3G0J0LZH81Vpc/VyNt/b+DBdG/AwAFKmEuVx7rcGd7/j37zaM72eqW6zeZUwxO6D6eUzQ
h+MFaZ2esaNpQtl408/pieMvjw6s4kAufkozU2qEykJIvLREIG/se9y5KFN5f9ad8xEMZ1MY9KEK
Ki+XJUNx6SJZfsHGQHIHfoNLJBc4ZSfwjMKwyfSEZtlllE8bOqh0gLBoG5BwDrD5wTleX0o/kQyR
bfvY0UwLqZTaBgvs/SWmBDQYMVx7P+w00TEpuSTa3X9onrn20u3tNNsgUdAtT8Hxo/Nlk4GZE//9
2+sfrJao46FPpRO9Tj2Vslf9m3aHjPJMtAfS7jX9AlwlxepDvNFHF6Bst1zUdhOsWDAwZj3HYso+
kcSNJhK8j6NwlzDszDATnzHVCJUspkk4GvperYy65SMzc6DkTVEpPdUlHEk1TPvXkJjL31HMqHZU
gI8KusFyAhhrNj14ZaTMGSkeNuu1+jqUZnur5SaHe/oW/9c3H+INPbncm2fj2Mp7XscJDJcjZOA4
WhMXPqQPbadrebvJzY8jn8fMFmEgoVcq6fywW65UPOK3ElFkDw3ASCvba+h2Ul+od83Gv8klSIMb
tPkjoqRpdJQoFlYxXHz2lOylr8ZKAB1rOGDoxm3Y5opVYZImKtEhQjt363efDrpxJpzmq7hXpwLj
oqvVmr2jSBjNGDJAOmJ4voVsWaz/i61rdIXSIVyR7h7IhxVvTowd/guuh5a4DaaR1jrZQjrRI21f
mOkl8YBRxdQoatsQs9yTciBqlkjaLV2yn8DLNLgN4OdyZKp/Ss5GselUoC8tEewytR7y4TDTFicx
46gQup2FHWoPRMNIExx+wrV+VN9WNVvlv+bBiJFkOKRgb9o1ebNEkaG988jj08PsWyuAoQYwe4Wo
bXEaejyL2r1WKJC15rSE2srwbNFrXvINRjwsS0m74nl7che2saG+LBpr0ynEIvPgXtRFM079PHLP
JdzxpMeWGllYvJoR4m/DE3R+oHro4Hs/wZ/Lgaa5B8aS6i7Y0j375rYgLv2+Z6r2qIcqPXmDPBGu
d5hNYl8HSj/9IePGouEoksQcB2d29QzhCfgyX462Y1ie3xgFGymQ0k9VQc5kL8cXJhbjbtNQuUir
KtOiTkYt6uXdx3TglBfr24DIP+vQLCpk8w1rwneCeJDJmxgocKFRMNB2wHHCP5ExgYw+DFgSn6cF
9iZsfp24g/1bj9PWjPBcxFr7byuPZsqNY9wtKdLAJ4+vp/vzKqtzhtZuCFaq6c7seOruzZoPrNIU
mcDitXUzSqtpbJo2KttODUph+c3F4xsINFQNW/9P4Sq3ZmDQH4JJgWbp9VIdkqxBHy+5o/557mgF
wm6uqznKya+PPRKEoiQawz0p1oR3rTHKBWuZGyUoTZXwl9KD1Ryx7DipKnlOEBMSy8qnSUK6Dkp1
bsmZZ7NcO7q9/PxlRK2RtItwNEgfhZIlmDRQo+GglWwFkb7nBaiXh6LpY5a2F+QIiMinfJqV+e3B
LehJ6RzuBtB2n6C70MADsSLce1XduOBXpeJD29B3a0DbXFKhXgoixobBD5cFJ1j+eVzL3Y3Nmnl7
AqLFXlFEgjnyddJP75n3+6rxcQASK3qlrUWcNSrnmqxH3dris2l3eU2VPKDD5E+ZIh4tyD38dEhD
P7Fkdvbh1nSm9Sp5aRnktDw8D+L0FMfH6PmyuSyhADsCrRRbVVlNDkjAskQJ+zWhLQevNjqLCbY4
ZnoxmJ6u7wrN90QEONiPrHcHzNtX+87FMYRpz035uiUvI1ue7PTT2C4z4GL3HTuaSNDcpbdWpd3A
7U8U0gQydEqDVss182gQw73hW8u/Qj66I22UomZh0iEm0pxxR4z9uRy1KR6+1+T6PaNIG0V1cmxQ
yTSG8p9BNGHAzxv03/jy988exrl2FTeHHBtWpFrTUcmziqYdCSIg0KG4rOxZd0nlH6Cid+Z0sZ5N
aeeMXkLv2fkRStumyiPjkbfthIVNAp2ZmXr1rvpDeL8SOZb3TpGfO4imzo1f1D6f0EISXdfqCBaR
M7UVNI1naFeMWng4ULgoYikFOHmhP/XhCccy9ZetBbMz5vGpCH2QFqliCk+8NKfXZBQ8QeLJaR3z
i17wuQsf/j6ddNErwFvI0yhAecLha3xoi0DOMTKi07bQxzcnkp73+nq1DdE3te5x4CUogHH6UlFE
RKubttAgiYFK/hZ3k840zC0O3SJeG9L0oDLxJjbW2Y9x06ymX1eXAmllrzycJE0L/Q9aUjCJYp8h
8WW6s7sm3mdwzLSUjZjm+D/PT4r7x1NnzT4sB0Qci4NPRybmOFXSalihQJF2fJTZ0+NdwWRq0zsX
MAX65nMNyh/+YTRjoHawWZNsofqEhFk1JXYAgDaCp75/dht1PClx1Ggdy2EwKoJWrgEAdZwfad7c
PCR7kmj7VS2q75MQNIHdqZ0Is/kcEXHXUTnJCu3+9n/u3z2Vux1gq8AZv+QEp8T72YMQiUUtqw0J
Tq5pIZrK2DdgA7uKrvqiUqGOooSLEUZ1jm+51fcq19TqJ7XRx5vSxJhn8nI09AboJUWS9ovgQT8H
PJEj87TsWx070STOpvkIr/VkAIlWZ7J7egtJTiRb95Iqg5qMBzawLSSQ6JQ5VOlPPLmcDp89mICv
qK4RcU7qIGiaMoAO0jq3pdd4o69gLB22fRa4y+8Z6EfHfXETtK3WDEpnX6Kb7q4ihbmSrnhPix9y
ykuljrOWKBgj89f4zWVwNdk54UlKmG2kd7MVddMKUGzgr0QeGBx6stIbS9RQGoAK6/UdiR4zB8GX
Fimy88TRKHCwqIg9w2bZI8+m8EyCq3IQXzQrTyGgaOMtHAEqztiN+o0LF/m0PKcNCXZx1bTHVdj9
IA+2mqMSyKOpoSKPCP8VBMjv8U5J0v3SXis3blUzVO/XrG1ccZex7/TRjDSPhETjupp8sy2omyD7
m7IQPlXeTCe9dTj3DQYu1YTn0Y/E89tDonjzdxAmp4cj4I+Z8lJSwZ7ahKIRL319sgJQ9dctUuoP
evGwVkQf11IIwG32iy2gXJgxSdJQECORMgu34p9pAW4NRU9fwyDoxjZbTtuH9Domz0mTwQe2IQQD
B9gsDNvMjCH7OY/dh56CilwgN8E6bzqPoll1l1on9WgF4v+9n0p2jZF8UVzeJbEz7OoAsOBFlVYg
2lHF3qDSxxc0MoMPS8wAp0o/LsW22h9RQf+u+Cm7rBMJ1F6OQjCNahRGYDwHeI4GZ5+p3OzXwlbO
lStQBEzsLlTczq+V1jY1rgrWCjDqX/YN22dny4pjcffJzIWukzCt+DTsiQr3Va5XZMby0C/xddwn
6De/AvdmPFJEuJT0RP119PRd8yed6E2A9EgW9dNtEWT9sbj1vqW5mMDAK8vrQVTBSdnik50BqmHd
pPmEFnRyTIMzJc0jLGMbKzmVipt4Ao0wIfvOPM7YpJelJpEERw9fOKcDJyTMaQ014CPBGoOhZFLw
+VB1dDSDcy/xuEXva1Xpk2s9eLSN0swkqaBgU5SAoOyrGXiMRxWjKrw38pITBUNEh85clkPUmTPS
WVhJrLDCBj3NzPg94OKsyxh/Sxj+KtvqZEQDhKlVFwY3hFJnCv58QmzbDI+3K7n9bMW90MiZf9dR
o/ar36TbmcEbnkMBatUYELEgn1F/73Y5umRWa2RTykSLs+PWqcnioci/XJMFi5SmIf/iW6bRE8ne
8amJT81QAQM12hIab5R66rBzRB96HLEAuUkS+6YbZ+wtwYHiWOaeYeejzSiulP7Kfy3k4tAoQG4g
muN8xYkMsdUdzluVIy3AVgHYnnZ3JZnsTQdWCHliBB7IiKMW8MzNVBGae5WOoF5pLOzNSStS3c3B
gVeaStAfTHbZ6lUwtaRJlKVVrT9/bEyz3fkduRfRup8vzq4M6qXnBlqfaE7vji41af0glHeqto4d
dQIhyX5U0ujC0VIb0sAtIq/v9IxBToz2T8CFmKgX04eS4/UVNeuBT/236FlP03nigqM5NdaPey5C
VUb1hPlRw6+wWXemAENaHmTfqrWQ4BOkcaloXd/lfHieaD/12Ox7CHs/oWJo+YBLCco0YnqjoEJ1
ymKanSgbgPdlLQ+KJ5i4HZVpbKcp2SIz4rGDPLX7MgoKkC39VsKlhnfyFP24w8FstY8L+MmwC7jD
BDsnrsFHg/Yc8naNxioiUJ8FJ9QURCDou1BSbp0E2kWCPI0Y4/Kektp9GzltSeVJUaf+kXhL2+uS
n2wQLNGQDmLkIQFFHpq/cvn2CtCRAFvgKXW98Uu2wlVXDQ1XRYAXizeAdxNiTvVNXTvOSeTWiWlw
RyS8FvhOyu5VH1lwPQNbfyWXPXdiV+jnk+Qrv9U+vNh3pFUzqNL43fBpHIkS2Sdf8TVuVBc8VDU8
2GStsnz5JG4RtufXlH5Zl09FRvUAAG2wGx3PC+2uUvm/jNctPJcotDR5oXT4AYNfVssuQ7zvaeQn
pKn+3bUMf4+b2W/znQ3lX3WZsFi/c8Tw28iDGkxraHL7D5aMYrGLlQysfnOMqjLMHGAaoogGH90n
QXLOLcv08smyPQEeMTclz9BdnL1xL3rCQgv0uNbjO7Wa0yJhXi1IYe+Fj2HOvyWTulHN5qEZa4IG
9ZOG1S14ia1TtL4NTfmUgp6lMvE/a+jcVn/MX3ydO0ovv8EoFX+1+FNrSAy5DCuKFYADRr/go/Op
7TEZDnH/2bIe4P9x4Ik7jcOVvkC9O0NguDVIj43kAxm6kUEUwGdkJxog4B4aFUCmcad8L84wj7iY
259nkCI62k9bHmyYr/1c/u1jCUveKdwGjJ+54hAgNCrLJoK+VvF6yYjJJTbKC/HnRryUmYVM6v5u
DKx9OuqFfa5s9kiBGr7o4ZOO32xY8W/2VbMuYoYyKG7JmTrtj7gT1RElN/dMwuiZLGv2oPoqQ7Ae
d18Oo1r5yigHFZC+wjKecBm7TYt+1R2IV0pzY8tHRu9iGC4FI3ZCGAH+Bm/iFZ9BB+6G/H5o9y9O
expH1wS15NGC56bwbwmQt3Pph851qAvtUCPG620axDdfb8u6jLICN9NxnHMVO6BG3oU+LEVH8hTg
kcG/UwgdhheQqV5/7PQjmIWO9mXYMzCNfHzdn2A8mLNa4VKnisR5uWFjxovuCi1RZyCRA284dpdq
SXHLefozdL+SoYfhs3VS0MrPzhLQSvP47H0/IaQmsBwFRm5yRRohf53nXFKv1aKzU//o2RfhDeYr
i2DCxpoC+5Hh3c+HHEyZWx41VEsIQApUXqOdspNeHDGsG30ESBUm2Ka+5zFen9F3TDSc8Wf3izPP
ClJO8cuLuxROZ5r4RwJi5xbwCOa3MS4xabWufNgEC3NdpMvubiKwt7RNAshX2RKsEj99mhR3q7Ei
krZcJ1+O2xmwjBuvuINDpgmE37tb9OrbA+ixIkbEzgtOCxCErV3MYsYmhBsm4/k7aYDPh7VJLBqI
zOsI90YH/u4f+y82Rv0gMo44ancx3gQDfVEGpz+sxszuQoR9fNn4krgCenaCCgrHSb++BP2Bt0An
6j4HxGF6f2ndQqN8B3qElhy4rBI/5vT5Wuxc3Z4PXZySUzEjYj9N/eTMbk+j6AVNepUcomQsNE/T
vMuiSU1vXhidrhzkMgxUpZDh47HYTlHkWbEVgoHgfm3P+QJJ/6sAiTzUbfelRsr8+8CpkOjmda3s
NCsxGwsfJg+ZiX7ZOANOs+FOkr4IEEbwcu5gfG1Y6MpepcIHLJM9xnZYvILPUjgmifgPiZib7kUv
NK6v3id/IF9ky0LvJ1b9L1vUvhyW8uQZr7ZKda9AVQH81blCiKg4m35qJfIKadM2PVUlYKW3y80b
hKp+TnvuTX9YZd1PlKvAexTWLfTJMoUDX4wYiCEw52YlUNv06l9m1pg7tU78AnJwd6ZOrt5G1oyM
r0Fp46+ap+onMRrw8I5iJRsJOrsNK1vTsG6D1ipCdIq2m6GVS+/UZPqeKmRzdXH5aWmI3BBUL+lg
9gcrwxHhg3y1g4dDdp0wuBDDgIDpTxJ/8Vw0KIKm5aPJFfk3t4pHeX4iWuBMU/I9nqWiVg6oJr5Z
RWWp03M6li1pywNaD8NzG+3c/Q4Hr1u6UvPmzD/YuYvYxJf/yI3/A3VG5sc32AGx/tJvcxMIubKW
l7acO0oqbTbpw5yHVda5JiIX2f3ZXGYb6UZZ8lphm9tKpNZlNGRkMJms52yFMsr2ueZGrgHmnryu
cWSrb6689tQLcApQ3zV5Vpq1BWbWsmWp/xKnOUav4zPD2Js7HaGzPKWRCdAvb5HO+dk+QATnSZv7
fxmJwUTVTcvIDHCo50sQ++lJOZs3cHDIQHVKj0XH7s45cD7yLcexRXGF19z3ti5TBBvg2a1aEGyY
UiYvTjnG1uT2M2sg2AgqTYQeUPpaCpwH/PCXg21zUDFPdDTsov1X0EZ3+hKJ4hurLsaU1wrTeK9t
SmFfcvaTDC0+YqAcs/6Nfddr8vgChdSF64TjOmlIoOXbbqtWL65QdHuh7GB/vpW4ZdeEshfxfEE3
Df9zAgOaqpXAf0BJAy2EQBihQB8U+LQpU8N/3jk5Fyk5LmVfiWCAiJ8F7tc2v1oSTLlNO10ymU5D
YyJuwb5X7n1bcnEljeqb69BUYIW8Nhxvfeye+q6EJSiYwCVBRTTHuFKX9ZvyM213+ef0cuMeapWg
zqoKlHI4kc1yMlfWFIRGPOYZALzMly999zQT+pQkCX34Spf8Bv9mobXab4sPzbTlarIdMAjejFkc
ySeHuuGmKTc/a4PrvF5ULUT0QYt/YEsNZ4ijug2veIPfsiCz0CkzJtifdQOU6kXSpq9iD1eIYSO7
lM/JKFZljEp1Ct0D2z14kF2lrVvLjE4AFS8G/mDTHRsALue4ffSwMjVTDbKuew7Qgk4T+/M8dYJj
oKGm2Rr3OeyWPwVBk1C62EMv8Q6tot+CvMQh6WWQF2+CYejQFtOCBm3OMeYKi0aK2Y530AhtaqeN
J200gZinwYHOpOT3BQ2hIc3i9CENABARw9cCwjGxnVzr0HeVzFoCZGDWFkfymtPOHOQ0zTpbXR5E
lVCrIJC7Ng5c6wWu8qv5zc01UDJq4j76x5aphQDNyJr36N+XJPdbwyXmcuOXaQWOOcz484XdsqCf
U5kGSvydYAevlj9/4hSgBRjwzhWYpliRf1ZI2fzUO9dIZHn9+ktcvX1BzZGzihGDK3b5uUieQZFg
Taw6HQT+wN9E1g8IfezkYUCq5DJedk2IySfvCYy2rV/fHWUPTmxHF+dgk2Y2sdHkWGPXYk+XSNuW
G6WVu1Qw5CeMkLur6H+FyiYLLcw0QwiBoyrhr64JdKfgTYMGx/jZVMnfrTYWenW4YQvsT2tw4fNX
Nefj5slYx/LbaOv6ex1volAVdQkLNZYoyWvYzvRZ2up2WURj97Ysv8giUEACIheHLhtN+t6mNkrD
y5DD+msAs3XaSxFTETWowscfc8SFjdTKkt/K6q7oINh2SGMeQTNUXy5+2cTO9NYKoZubnBapah6N
aUtUDzvOCKu2VOwUsjQWOIc147qjHS1d95naF2iTlXkisT/NYS/kvDocQ38HT4FUy0s6oxhqeen3
aguUQEjsxO9NE6qLyVohDkalK2YzBbKbjSZbr6w7M6N1zYvuN2Uvv7hIHFHgyggukssbTClihMkG
tqpHYhMUzzUwTS5TsN9NQ4Dq76VOeIM9l4cYcV5ohrxK7DWhmg0i91/BRdJBADxOQtxkRSOUIdtH
F53V/mCaNEq8lWZ1ZJhelj2UkSuLSY3RWOUjvJweR7yWy9BmLWAgbIW8/g4CTvpFASb3C0mEGd0Y
22QGQg4NnppcdvVG8rtToqpmb8Y5A8+NVRgAzOOxi5Y9hljNQoQZQwKEJIIHv4d9h+GZhSwIrjNJ
HEquW/FFAQSnl0fzfk4z6SULIu5AFfTDRWoXgkxxZr4+Y3Mr4yeUbGYQOo/25T+zcCf9luztNDDe
2haKJRdqBpcsXHw+SVmcC7xXiNCV+sVXRMBvZlv7RSqm5QzJm7YX18kXcVh+2m9/6K6OZT0FwiXq
ifqy7XFj+CEQpqhOxz4DB0BsKdT3meOGqM6UpWZPlr5re7JYfCnQdA7hQXZ85VdlELMg6A3mEhqH
3qAj1DFrYdxTloN+MHjxkOUFgfl3Fs6D4DClpV0Ay2gimmLG10MH1uKR8UndABmGYi1bm5UvPs/E
jH3VUtO1GulGF0vZLPwdU2eMEKEii33Y72mT2hsiizFoyjacLWPi5Yqb52t6rZB2XxDUzTXarxXF
5JU5hpIpdEa2Mv3YiFdfsZsfGjDLrlzqKIHkwzT7SbXXRANNoKL7R6aSU5qK4CTZPE6bitGk8kDB
LICMZsQpams/tqnxjRfrP3x03OeRYqGVSMU+Qw1c8BLU5JYK4M2DWSs3uC0Fw3wn3MvGYeqS3yQ7
NGLFqhm8JrewcYRlgH5r6AO2vMvFvdsWwcKcEwr/HKfA3kwyhZSHl1be+kmjmtpjAzNYhAAgmSb0
35mV7HFavREgY67f1xJBdPXvRrEJmDX4+Jo1IgHf8B01b1QAJ40nhq+gegdquQAG6qlfwQEYZvoS
CO46r7LL/cLu3PewRCeg6/2Q+ktGaTdnAsXPM7DQ4R6PD1+Ouz4f75hjxbMjsSdVqy11/VwWnqHs
9IroPA40qdqLEzy3+obYgb4lxhkcMu0K+fZId6mWym7xNuMny2rYBhYjDvY1FB7S+XqqZV6IvijH
F/mdqehFnN+HaKQMcCm8qSHJ5HUjQNsH98VFT56aAH/uBpSTmJbHMf7r2uX2FZpkSY2ipE6MaPx9
pMONBdOjLTv2bQE1yqG+jVA6I0TMiDG8KRhI/u5dSgQo28vTf41X686qrVaQ17fKKZrfvSB7EW5g
oRjyBEiDnvM8lCCYRM7tcuPtuJ39HySOOEsc9gZqHve7oT+pyft0ieeonMHJsse9vhcNKACbcZjB
anz9XgditzR12QIFL+85tVusmU7RiR10kXukmqTOWZ4CWUQ3GonhZWguOslM9Bg176Fh53To+fvO
bt0pqW/LILtIqE8z8teqaxLErjVHvD7tBpI2q3OkuHSDFQGeRf259gBGJbFtmpTOz4TEZ/YYMuZf
MoUa/efoyrUoM/1svrMICLgjNzCmNs9m3SWY7+OzPPqDHMrsB3N79y2iNSnSXWiFAx4rf79GM21M
J/EjwuLC53bLrFIxhu3LG2BNPQvGA7q/XtDdN/1Zhrfht5AtmvYrgAKoTjGd1ZOzODCclnMptMdn
vuFbbf8vHGzdef4TPj74JgKByRdb4XOOImSl/l0fOqrig5liqCWXF/o1N7xFYm062ULjvSYfEY2n
ND9uDMICjo8IuX1Zo08AQZdgOgVRd855JDxEqrNWqGq9HrSChZe0cdLsRhbSUAmhBM7Av1XDEHaG
35oq4mz/QYg/6mo/K73af6jzBFgWaaVonsWc2QmQU8Tf3ebXnF7f9lNWriowPJx5/Q9fZJyTj2Ok
ysvn+2TmHK5jj7PM7p8fWiXo627i1RylHCbIxEPBOMqffXqKggyYf3ZRnUaybyxNSUGltFWrtQ+Z
ABMlnltRk1UxDT/xPZBaVmD9O0cV5X7SgOqcvbSTP+dFsNex9H8Smfzns/Q3sgZQRIwPa3FVfbe0
J2h4G8jlVWpRwhn+nxIlwW5NL4E5tDsx71Q0w3yLXhw6opARl7k6MgfdTChMh51Exxg7gwB2AYEn
3eSf8LfGNUZcdSi2/LMbKckdvaq2YvQa34Qyb15gTshLEDSZS1N3DX/fA/yKglPZPMoWzSy6IQ8D
jaBYce1WBiMUDHDGiOigXQx2l/zPajUqx2YMj+6gGBDSj/0/yEYZyP/rOEDLkw+xZ8JSbTX7qTHR
IJjJ8p0sKnRoOBmPpzPaj0xgK16kogfKR/WFdnG5EXNUiSig6NGCM2S0yTyhFtcHxYoltOTczZzM
M9Aaj/Y3J6a7LoP8WA+LJiPYV+J4yRS1cowSNikfcWR3G+9ejfChrORQxGgT9YmUKORTzbDUptPI
3t6XoSs01dWHBUVHkwH62T6r2D12bQdFE0WiXFGry//zGj9EBuTVGSBRTByWwW3iMuE3ofK1ltGU
0AOT4sXdKv4RPl1u/HAjP5brBF1V9V+O+ZxR3AwMnuipWOCD25Q0rEmorwNoLCN8dKm2+Mc5yOfO
1eMpVbBjfLjHeAc76KHPo4z0OCsLOnCCprRIPBZlngc5mG+pJ04uzwBax2vFgj7FPUxCU6V436AQ
EoU7vB8e3fHCnd1Y/FO0bwSHzx4kfX4F27ZgjCn3cppV44qobW18nnD3rDmJiHsdOA4MVEFVmG52
GrlspFzgbEvk6HAFmFWHOlbtgpfx6Io2FrGErTM30eo/yf34KPhlJHryDKbbNrzsZUVgRq/0Wwh5
fER+zS5YYnglTsXM4Kc94j2YESIa9ZniA6CNSlcJEhfzcECybCpw8xY16fzWuRH7LsbGwI0hj88y
wfQlZX4RyAC5aZVq/ijOG4DkTIXHJGVwxmslamG84rNixHAVDDkuJOVGXqbf2A1m4DJ4irpmzZDK
bXqKrf14nRrCkt7ewUpowRCl2elfEW7wSzR/WM+l+SzjGP25cZaGDqTZ7Xz2Da5U8tvL57PTzE4T
AcsIrV+KiJiu8jq8NjaL5NJaXNRBdBPpzjcbysNF+bZznmZXLSfZLPum4ceWXzhzpgvY2ewZ+rkF
6seIHnDZTppt00kv6Pn704t2/HvHdSO7iu2pN8eQ7w4GFjAHm/FCAS/ZjyPzZ2EyHwaeQsaw3gv2
mySNWz4aYO7ec/bjTL4eJBvoHNPucJX4rAGBTfonIaRiyNqBF+B1xDFdfHd7xFeY2koWilRhXdJO
QKBBB7zCT1kB8LBVmpA8bBPUWjHiqJTAdAK1/zcLaCzH7XpD4v/AETzSjFfbjv3v3n8QPTiR0CmF
hPekWk5KB4XNNMKoYjcpkzHuf9A06ywUOXxD3HVmZ8bAu/XaMXyU3KGB/HwNk98tonYnb6ZcX7Au
GWqZTKWsjdA+Ukcmm/Pn00IZgd3E3ltpL1D2pBKXuENxEmEpd3NlZrZZwuZvlrp0PKpb6Ye6gYEq
4fvoGNu89W6NzKgTDvZBBmIzjWk/MX0d65sOnKLhuEIPfnbVytlCgSR9deHMGm7SgzLmbNlB8C0w
ivrkJECvSr4ztg9OBEPjpghHpHsU9gdxahakmPAE4xfDpk/tyNn0Vlenx2vzXQ2oC3976mBdJKhl
s32A/qMIK+47V+0yMwi4mayEcKG1R5p19ZgfIA66h9eOlnsvn9xwuti5gJl2X7pkQdX1v4SeEOci
9WQtuWzxkrkv/0Fprp4Zpo+zbHCudqIItghAZE7+KnXOu7M1KZXHizG8JZpXh7Rlj2x7g5PwzQCl
AoCqCSVtH5TeHHjeh1yEt9pOwpCQ0bzbQ3w0UoN5a+8wrS3FgC9B810ZxmDlHag82W0UwAJh9PAv
fim8KBUdTDz5LxV5KWC37CHUVZkZTrdXZDYxxr7qgLgqkhF+zujx4A+rmbBuvFaOKiu5rp7NvACM
U4edGThPXkuds1v4Zg79zx8CaY/eaomsSiRDvR27PYfDuo4MroM0uPhqnAUA+P6l2nPEXOZkHf5l
rgBURazAwoHVgs3IYebpz+kphAQUy+RON33yELHwFsCuVsXmP1UwWkFkX0Q6IWZDixkrkECl93Gt
jbY4GLbQDx4GrqETT8EbcqF/3T6EYtt8f8512WmNcbx//z5HPnuj/owJByqINGc+oFmBgHB5ObHz
rkVn8Og7v+AdtUZfNzu9QnJRFOCj2oecVy8MPoq8hBvlq/0mY81/rrghAOdE2517Sh1bfj/o4RT+
hS/npFxI0B/ziuppnExx7ja8Rku1qJPMGUhXJy+mDOVB0ze1TpNgU8hmjBxSwfSRYQo27qg4QZie
AuGxnFJIcwDR1pBov4fqPwEXk9p3gZ19xFlKnvjHLhrLPEg/XV+vGVhUFKoCl4rXg/GmHwPM1s7G
zzhWbn5EsqqcdzaYgn5z5NNy3Ni1Shr9V6XrFX+FFOqVpULpNyv12AGufBhdRH1zf2jbPmwKMjIF
BjpBR0ETC3Z109cPKn+C0cj84cV/G4vRSPs25AcQpS8Uj6vYhSmFl23XT9weiC4i5W5M53aVh4K5
2QJQAmzZqi/LK1HW1IaR3zQiU3vt5sG6a4iuOWPG8NlX4LdG+xqZ8EIsybe8BgpHxvSNNl3LoEc+
MZnKQQX9ThdcuopBVJ5o/zqq+rFp8Podk749G5uKeGqPlGqM0dpru8YQiB85fVbJhihbqX4YwSMt
NnY09hHhxubOu08fZjvJjDNTDvkdGcrp2sYppOCjj2rWQZCwYGY3VNvj3UDc1KupQz3TIc6g1/To
cKmfurQYB/hHkmwC/6YSSNR2TSRqs1JdP8/LUaYEGCGy/pgWKtRPdrlNh6cwOpZV8/NJ//oRpUIm
704i/MedL8hb2cHRxMHp1ntFXsBGJao3b4D2s5pi5VhYJb667kmy/wYGcdzhn6Bi0/ddWiGAPuGt
IbEPY45KKxA+HK8PpBYL4h14ePsYmB9704TM0bFDFMFMJBzgiw92UQwQFXgWutc1Z6EFFOEXN0zc
Y6vM4VhV2bsE+qs6vXMJTJ4cHjVYXVO9ODQKVHum2UCMse63L/1oH76EVYSSGlpL4GcmH7JMnmhn
tq/fLBiUkWVSv+r7IYHPuKOFBKLkBK7Eq/D2kJQjPy6LsAiqZE3yF+kDh7zFv+isEaaex3Bd73YD
HuK8QoHx5fQ9g01MzvVP6hPhZ3pU6E79nkjFbh7bx2k0gfuy8xA7wFxphTSlveYBzFszg6eXxLHj
s16G99gQSxYnoUbJcS/dMO8osgrFkD5HfA3EyofYct0+IN/lNPXvFjxJSdYOw9dli705y0gULhsr
TDnKf2HEGku4pJHc7mNUT2Ftbm8Xd88xSiNYJs3Xzzbw7ssjXn1ATeUhUy2dXiy03yjG999EfirS
lr7uz00ImVo42VsHWvI8l0M/vmctKrYGDaB1Gf5zFc1X/6ykD10BXU8YPOLnIeJ5/daPXqlwt6HU
kSW18CZGdd+bBaH31f+4kxevWTVUAS9bzLo74skQ2nBP0fF2nDMVGIz3hKLqoeRtIJtght0AFxya
0Wo8CeCen4MTwSsYJsAQZ+PpbAuRTJeE8eW1Xe2ZxPKspdEhi0IvdZ96uo/XeNTtZn7KtVE+EDSX
HPyoqhMZlKIUQPVE+uxFuKZgY2CmgC0YUghsXvJrqW/AWJLlC0EIPqoEkz1C8wKJDpl0Lc0Aj0Ct
UcLFT2HntQTStf9yvJLKZDeTxQVKhxNYS2gb3ujg6soRv410tDdshU/3U7cUPbZSKbyUgIuL3LL6
tl06nLcble7AyIksfyRTeCvn+GhbAxckzsHYA9SHjiPYhO3F/ouYn/uFHOAreo6Ded6dhT+3bcp+
YcAR7Jd9SGIONeaOTSvEPXbs+0hc+X1DM/11ZiLRl3aMQ4IoKI2oGj19SSi0DWxLExQtUFMQHM//
aB90nSjoQ1ECsYWOZQthT2jkF8YciQSS3vj6LGiqxWuXvM5An/bO0GnVC62+AZGA+opa1ft4v5j1
WAh7hEiTnMFDG991EDfzArBkcbEX2Zczlg/wM3esJ0LMCnOUmnm7E4+tsnqVcvqJn4i1fY9tmoeI
DadK9B9gCyLLkMYoVL53/fBeIv5DgFowlB3B4t9+NHI3k0PyOjzuFVf6/ninlVImzt0Xf6sMZmD3
u5/WvYSAHWxYEVuHu0uFHtG0rUYSQLK/Vtf3hPfdV7dPuFs64/R83Fv/C9VHo56d0hkGAhMgYBs6
GNThWHWi+nu80fA5b/6roHp68yraprdBJ2tJPOe+GjodfcWuuukZsqZVTPR+Qg5cj5fPU5v19S72
6N+kraajP65NL77V5cQIJsMeT6K/MKXRBQy4/SEMREEE4QrPS8tR5Sn4mAls9laoPDVFVrK5FzlI
c2v87SD8oCqX4tP3iZP8XZ2/Phyf5OOB2KCRp7OtXJiktruWy4+VUmnIIFD6BrUiPaONOqMWGPMR
uNSJXvm9ppCrkBRZP0BDqRh79ObV3CzS3UUh6Kgbe+EfivQhCVqXbCv316UoU4yKfUp9Fc12732X
PqwUBsBs9RgaMbX70Iw/Mj2dpUJpk0LP40MILZWN9WzBShQRqzQz69n2UsnpH4o468vAKR5bWDOz
H/jW8TkKtBcEql8c7+t0l7L6d9mITdxXa40lMv1WCO8oPevhwBiC7Gnxo0UaSSa7oG39QJW/4pBD
NhNiSaRUKvJqNjWBq8e/hnayiPEqoqLhLunJRjHjz7wSd1fOgDehwf98fuq9vFJzed5zqBnoKBRn
G0bZbGL+7rSmoMftOC97Xj1PTRPUF986wPXxQv5Q+J/a2o1OeRL7mh88DVY1JGY7z1OzKdSu0E+0
v2nMhVpAJasMxgFN/VSKK2VWEQmP9hu1SXutKFDf1R3w/B/sbzC2ur0MuyU/u4CD1bqblYj0t+IT
vOA8MFGLS6D1U6lNtGe2hKvPlg5yP9i0ieVd2bSVT4zEzb5wTBE3tdqIVHyhM3/57uHasuLVFZ6J
7/VvU5L6k0dR4EP3Sr7PjzEqVJfEvOHsI3cqJaEmxFnwh+HaLJHhPf40+ZlP94C9nDciRmSFVAF1
syQyt/mE+sCL8gS3ERqcEvf2VsUtmW0CJ6zwLfI8YcFJWzsZMZvtVBYweSw6FdsNvUMXfjledqzj
Yh7sDBlBxxQDzi15avtVsuqg4/ftbcinZzyPkxIKUm69pstEF45UTEQ5bPbvQQF6dUt8hfTzjaj2
D1U6ybmUN0nCAjE7CNdwpflYnZzge0/2wCPydp91CO2MZZxcqEvs0X0Uc0tvaKHGCxWkfoX4dDcE
KrR5eQg6H0EmEH2oCGmhxe0a/JWNa61pMtXkpoApZh87CyWgSYoD1WgWP8OwM0i3bwNAcAJDONkz
YYtIDPIdqV+Rv5J0pFO/Niwn19jGijMKfJmwwQ7DyybBYZ/4iC2spOvWYC4azrAAyH9Td8Ack0qm
kzqY7ufB2h/I+7maYJL7Wt291iQlWiGm8EV6ru6kcS5Hs/zmn7mHZoZN4BVBaao2J/Fd6TWuowD7
CDwAF+ulGmRgjeX5jaJ5bEPUuT6kjU2o/2jX4mbEstdtDO48jZoYfAimeaqjmNp44QleJAcop4Dy
54qTi58R80z26xuJqAOkQPFbsn/WiGEiu1zmwCp4QLLOFBRyqqImCoScziBoHjvSsSY4AM34njk6
kvMTivlNpDZkJtJeGK4ZDSnb/6pwl8v8nVuDLgn4CzG/Dh66j9zTf6H01JA2g/MKgX4wTkLhzu5v
iNiXfzbnZpQ7lUVxY1WZhX0Pg+GchuFLWE4KImWhfY+DNainy1wNoXa8Vjqis3gIEU1IywnDZUjs
eGMuyC/sWGqC2Uw3LrfhB/jVsm1kQngNbzZewnGPfOtmAuJw4gXoxlE3quKvz/aN1jMDI5y+kRu9
IB9FSLueUT86FOU/Hk3KTkNXELlVGKhfvaacfXpVBAo30jwkhb1tczxIvZAkqvYw3uGl9TOG7dla
J5LNUWh3b78wL671V2Q9fCHefQPTJZQ0OuT5M9flC3AQg/sUwr7hBWoHMHV8i/ER7atvYrNO9LrW
rhv+27q1F52eQ2gbzio7y9x1fQXvkBnW3jqHSrH1aDGejwFTRg4pmaSxMbmi2hPF2SjRzKkTD0/Z
96IZ2pUFxTf165UQejuOfUIh2N1C5WtKsYCQjHtpdBEjQeqP1/jZbK6LIAtTq1rPnTX72STR7pkN
jfS3VqLRDp8uPpG0eEfe+WIsQDew8rB4moG+bCSA3LpOvM89ok/GLM66VSDv6iURV5x66TrZesFg
tGPIyAwZSyB7JXEQXlkclI/Fr27ryNpmSThB/WkT9Dcm6Qn8TE+BTOWN6H/8ZviY8cJbnOSCLA7A
qBN8kmI5omYD5ZjCFC2M0AiIxwPhWtBCnMwvpDkVskSoW+Zk9p2qRHjoDTqoos9RfmdSypXK+Twv
tjnM0LpPehrOKtEak2yB+5Ff2aPCTmDTKsNfk576RVCVu/B6nrH2rRIpOI02KVy2phcfCO1D2yGl
9Yz6qP9zXNYLplc3cMGI3BGVAHMRO7vnRnlG0S6uNYxkNzW9BM6QfayQ3M9BnNoKaeuMT7NJ+ZEc
QWIk19MGmOPMe0uuFWDngN3rLRv1p5KeyJGgM8tG37BZZwFQhAw4yI6ABq6+AWbNKVGxPKOtln5h
xS+u77uSs/vGxFYwZa9la1Zw3VS0/2ZlATuOYMOsbqCfiGKii6jh20jMejwQcD4Zj38UeBJ3dS7a
6uv6vWcPJmw4rt3Uf0bjwjWx1hMO/RDllihek2J88LC1+iT2JeVgLQtNwAMms4WRTLGl+bh+Pdu2
UqG6LRsh6IEF3rOMRgn6EwsayAfI4mPDvEWRmTWJTsGbXcz3aylPR3Bk3leprayuhrFIzUkIhEU4
1n4MUeToERIYTqStFuNC+TD7Arlm72vguZvt/SZWZTeSk9VIGvyWdgkW5tVwIZzP62Q7pfDs5WpP
13OlcQP3GtBFcBZ+Grz1YR0rUlGtvk2JvZXqCmQyyBjIS6yyz8TkYWEwz2LGsmfTGXoou5o/ISYr
fKmjKr7htLs5NBLGBIdyuB0bjvBfGirY7rPynEsaZHa1GMVR3N9CCLQIwK6+3jx3nel2O7sVZCCS
zX2faaSbWx9QkWUngHBDJYLZqr3xftiL1hxj0gGrOvNJswVTOYclJNxmn/iqBfl3rcuSk3bMJ4JI
AF7sjyO9eRYdPJlbOdePWHuXZPCfwmhLfMre3rcr/BGBK3PPKG37RmN0dSRdrRJ2A62gxvZgm5dF
2VGzD6ZH6tAtbW+fMOQy4JK+6+FNdyEf27zwzM4PyBub51XUv6YON9Lphhu7BdpCQtZCZqHoG/NZ
jJWNSrhHlwcWZIpfQS/3vqnlNKtcoSmaE6chDTyJ19/kJd9e1BUnPnC8FUprmSsvOuh8BqhpiOqj
ZJaStgC1Ble9KaEQsjKecwwKtHvzCwk+C51tVH/jUWYVIh2TTYB9VMRq/2kHwNwo6E4hgmE9PWE4
IUdQ4QwDpYO3kx8NQzpeL5oqfcSIP420LWZXnBhWvUpgx5GbBmScPUrcz0L3S7rP6Q1zZNXZGfHK
dgilpsjPjyDraCr9SBi93p1Nkq26h0AmiPcUm2rBmHelT2cb5KX0y77u+qXI4MamdbOULfmWzFdL
Bo7XmTeXX21Mn6Wr1VG7W4AKFNm/QPIWVugMIavZ4MaQt7fT7df8Qj10tr3CDENuzRAXUSHsUY7f
i1yxSzo/dEHgA2BkRASDuyvBORqVuDQ3WV4+UJJMaHtuImp9sBVC+W+/u5YMnewnuMz88ZDcgQNo
rLkE0Or8FTLg9Ln8UA4Pi5zxqJ6orTfCPHJHP4Dk/5y3EACh8N4EmCUkLbeTpJOvVz9/JlnFPWDF
3fQNAb+K2pg1ZAx9j84MoZICjZDGbJOj3xJMb5KCtPgnR1jrdFhUD+j/qaLPMu2tKNNAy2020pbb
B1mRi1ESieUi+j7DPLsxC9F/fOTmRxRbHctjLLJFCg4npTEw1vKJ5RJey+4QNKkMqhyFcRfeWAsI
GOlbdZgYhyf3QiyKcX7JvC6wcYHmcxym9ZzOokNkZrunAtyOY/FjrD8og6evjpGzvmEarDDN66QX
GQ44CdpeCiFvw/4KTj3RlO6nDh+s8vMv88oY2H/eS79LtHSvnBFXkyfuU11NWKvss9VaSy6TIGDQ
/MDpcQMcTUjQ6B+0fzkjtrcdHWjdiAR/vRsvbsnNmnCzxvyqb+sdXKb2IxaEahytQn0CiwrIUZy3
nDZbRplTafGwcC/IxDy/QXctu+Dfzbu7eY5IuHhPREjxmSeqEYj7SlURnPOK88vAjnwU53kH8ZWf
NBWBA4rmTl5QzUFo/M/LSfbfRXLf2bRXIw08Ld1XhREBKraeKOTCBvK5I0a1ENJvIN1IbwYX3Mlj
uyePlZrSr5rcXTieLNstzFZ6kaJEJjg5N7+ggrbNHCtDQ2cGwIGnOj8V5BS9rtPE3MEVo8HgEhLg
aWAw4ej01TP/5TUa0n7QLfbKHB6oy5qYQBPJ81Pc0LyTyWYTsEnImlODLgKBq/PQjrTm9tASMqlq
MZFberkxoLBYFHmoaQ/SE+OpHLBWggU3vWwmfKmlveVkBbxsGxLo9goeh6F3VvFf8TUf+B8EdAF0
GtDy1kFNqfU+9UrTjeQurny+k+TfDIjuCtfuwfuWHZ4wN3i8vakX4hcFTcfHzFh3C4wczZabpApf
t8QZ3HCfAr41UW1sTrPwSWK2paK7WprqZSJGynixHqBjIlchyjWDlAvbGNlgLVMV7BXjHQ0kj1it
SMU5324eXGSA+XSnj3SOhZyh4O2AgQvv0tWiu0LNmarL0Odpjxe4oV8FySBVVn0kIoEX031L94KT
2fGJ5HK/8BUzbNc7u36GPQbW7OqLCMW5+zp6JlWVIPPtiDNrU6NDyjAUHionyd2YcEf5q6YU8bRV
42kPvX59tWSHCbtU2fmo58upM2Oerg2PriWjS9A03W01yc3E9D7fPB82xtneE5zB1YUdMXUV4cP2
Hi1MhxIViPQwDl1SpL7dhMwAM0+S3IH62VB1Ea44eJYwRa0y5DDRJ320ly1eIpbW/GSKSchHWAZF
6rwl6O7Qtj2t6SdNmBO8mxOkV9gw7BakQWfvu2MPF/aot/g/ydfLaZK5YvoNTia8Dv3Xf23nk7wL
4sjDYHk8p7JXNHqctHrJJZUVemWuieVRZX2voMGGOOvCrPfdLXw5lMYJ7MafzmVdVGT+756PwacU
Dx4IJuxTEwXOb6WeeKBmKeqRBxNVtAjVBqIXVoIUkhyaCjHkq6XyRkXsn83AUyC24sBgjrAf1p25
/2b96gOh67/vfNs4+rZ6GXXTW5mb5ZjSaRfsFTxJaID2YoNx4rQA1iSYQc4pXFmGgIWFMmVVlLyD
qTzUpr62+0Ip/ej+Ft/1GB7oWF8gdZ5TmfceF+kiZAjVNA14JxoT5Jq7cQqf0QM4SZ8JzYDyX9PZ
hwO584D8My3BTOdal6938BTvHWHEqiVYTyPeXr8KE1vRje7EeQsxFDXh5zrhnxuq+LH8F01tn5mr
eRwDzP+XLN5Z80/IRLN0Ffl6yUrbfardQFs9gbac6ve6ejZXspjsYUlGpkXC3am0f8zAahQSrHf0
LX9vXivZarJtLrF4hbteycHRFEAegYzXrkPzFPpFH0eDNKUFiPJVESysmNMODpPi8UKMGn2w0axm
dhDTXXS2QNQu4+7bNb5DoPghFPauXLN6TTcsDWLU3AHqWrnNmq2q5iTGS6m5I3JCrsUiXp559Fg3
cRkO0U10FCvl7Dvn+W8qU018j84pBXn5+NF7hdDGbGQzGnYt2otL7vWPl7t5bavQ62EwN5tK4OWE
CFzdxUhLvi36EjT4QFAcAmK9r6mWXwxK7tLSq5+mYOUMR37OYT13CkjAfCbFLi9aVrbFbfpBzluc
9JOriEq9w3FPrd4aCQf20tdrdW44a4DNf0kq/MiFY2AJnqlN4DCX38XUmQyPtklZzKSwAL5K8SpQ
rQ9B8YukMccbcnp5RtMeZUkFUngaFmMLeb9qSvziy38uzNRD1CkD+jE49av73pxEdb3AJ+V6O7P9
33t7k5x36YzXTffu60xOg5aCtFZmjC5GuIfPpRYQg5OIVR9CB58300OLOVJzCQZgLxRX924nj8U1
u83MeC09k3mJLhM8qXf5+0xFBaWB04Gddn8ecYjm4/R8hPkagYuys74/KTxXwML+NzQcum5UkkVD
n/ixY/7+2urneAS1jSiCgYEZdbVRSfCvmqLkAdMpajFHXpli1MgATAYJm7seCtZ69W+ARD5dKmMM
uFrxoSB+vi9Y9Gn1+4xsDZFcuDMSql4PKqEWfHZ65BxpXUA+o9sv8KlQ+yxOGoFLP/F/7l2JyMHc
b5PyC1gl+Lq23BtERKr2IUEb4yMuq5ycKY9RT69GCWF9BfamKYfP+Ll61b03+CfXSOcNS2lfYrYI
sARRCcHtMaixmfL4Cq/DSbX9cLWbZBZ6g7+OV+J8NapsBdEPHbocTNtP+TSqhBSMZTIBcDuj8Mx4
cp1N/TlOsIz/0VOje7RRycoZv03wflH5N1Zv8H6fRWHrHBLIzrN3BqyNgECO0+PO7hVeAKDWGo1l
fJCgCHnzlxGUXue2wtSw9WSsGKreOHFxItizaLJkp7B4+xn2hZzuJpTVNggeL7ciHC9wPjrRR9XD
VUmSJXq7D2rare4g/8xjGefCbzRBayxjFn1q86kIvTzccA3je2dvcMSz6tJvTTPsthODFAPhZ7tx
nEz7mN7k6Nf1xdexzOY4/TFd0pg0Z1Y17RsnNRfzlMq6dpGB6E2LF2VdpyS0z+tR1gayHbjHsaNQ
wBh3Cc9jKesNQI0wU8ZatARTJ/6JMGVKJ28/oaia4YE07JMAc9dXINpySKFWrceg0qgX0WeZ73oP
7IBTNq9e9sNQE2gBIa64QPP0fotPXK+EVvvfgPhDx0BtUigEBtWNiA19ELxreRB3PBFUnbTUL27F
oAsXTxpvvye7k9kiAjXExlNe+PYu9u6rjWJkGAF4413YzW3dmlIYYTgo+Dwtj4zIDF9+1wFQBC2K
93ovnRzmaY+Y2zAsDljnHna0C3iHRuSf7hPMWtYQE5paJohXO8+67clmxNHjUK+Nq2j7Muolwz/L
+CJUNn5RasRuR8dLPUQjoExq7gBkK9UTR0RfhqqWRw6orsuS3kwyWVgCmPua0ouUq3VLBHxrRa3Z
/xHdhnY60xciOc77bnsL5TNvWzbY1I4mPrhBsWQP4OT6qDa8nWqU6qV3CEiBQYsX42VVGtLxkVNt
P4DGtKhs1+VlBXy3ciAXxt9Uxq7opZKBxatJ1ppHSj2Dcuh9+6Pho/44z2lZIZ3dH6SLEU4BNve6
2VdO+peF8T7uBcKIsX4RX0II6u9K9/23T0AHqMviXgku6cw2lPrKWa41aDCljYTiE4nWIKB5Uam9
+MjlPdjBoXm28PRhp7PVjEnByfvbUyRe7jtxc2xtjLCCrQb2FwWJC4vZla4dyBqPfyoAxhgh4h7f
d6SWBkppq4FL3bfGlNtgtsZKmbPw3QDxXcTtHKFIMrC6GKqSo58l6Dkzk7eztJ6Aht8KSssNyQ3F
galWeKZk+xmiDdgXXB3VJBGmEZwFy8zXt1cQe3tAKLaphVBV9jd+EXcUUDuuFuiFo4Svi41eyNHx
7NXLmgymY0B/I4jPj0QC8wpD3WG7FL6Fbi6y562SVxVBflN2J/xDIvRfHn7/71klmTOm0VeIkvYv
2SZduY3vCtxXJXwy3c8EA7sB7EJ+UYKr1X4M2slYCiMVsr2R+7x13HDeCZXvoVbI3v0FVWIUvPc8
XhFDUlCmdtR3Ads+YWyJUZsxPhaSFboIXXAOx/t7vstamqWXivOjHMadeh1xU+Za/iylq1EuDVZu
q8isy3lADFN6gxOUvU+ZCdGVsmfiuS+gdz+C0zHWKS3ujFYnz2mWWZf9hOo/jlPgW4VPdJSXfSMY
uKdORYbS+DbRlx86VgrlSzFndLaDCuy1ZTNykyRyQNW8rRGWqU5804Naif+2IG5xjT2lVkWd3JjV
oXUC668MTppaEsG/78ZiZdSyuho0IaMowe2+SmFDSlLGzBxR2khFpAlI2y39fB9mKKxg3SaFGf/p
TOnm1aKIkXECac+uqUGqe8vwNOS8Ld/bE9Eh8GOzpbdfNcgfPFcKk2np4SUBSIpJ3BM7wdWTY2a+
JFtN50GbU7gPS0wxo7g4vJruBdLhp08oYdAFtVGfjiUCZdyPpObP04+a3gwyFOCSB3fGHwPk6Sb6
CP6NYMRQ3WYH4JhbJF2U24Dns4iRlt01yR4LJVenSp4twnNu1JCXpAA80ECRaRWGGQNyxHUNmCkj
v/vjs9aQhaFghQP5WAnJuxflF877gUiJou2VwtJjVFKgxSVQTQDxFF5n9TmWUO/0j43ZodODKqOI
/VZrXXlE1KHLluB4vchRHR8Ysfn454YMkFugsiRIwgIqvSqKZZDE7B84om4LhTbBJFUmyHFvlwkQ
O9eD32a+f9yR03ST6a+PojEibzEXodXBRLl3pGAIAlGq3JKKgEjBSMBFvExkSGwG4EmEsIPZvrE+
tqfwd8tI1B36x5PE77cK0Zg1qB0lpFjjsvwKNZgTXvEeFvEyS7aajmY4w8aaVsPV1Metw1zo5Tie
Xi8sydkXRwzP7hr4/HIsyq+PlUOQvGTAmM29Ta5BEoxIYA+feHsraDGT0AlyhIYMRu1CjYOqNX6Y
DleiNV+F3qLDagXL3lrtNGO5Kb55MMhxSZvrHN69PdMCfXFCwMsyAlfSTIjrtr/bGI/twpQL1l7N
8D8GmhF9zEGZwON7veIRLq9w7uTyw51fbkNto+OmumISogqEgv3HFTD65GpJffQruEyhIATgmdJx
Ozt/W6yql4gyVQLMRL8oVCE5OGOnWhnvCjADD7p8YIRa4kDU3DK2fhL4UIhdDR9oZD4E0ohjOKY4
REGC4EZDYmTsh8kZIKc9WwOvspXCBcJpzlwkle9SiQyfNzHM7aF76LmIZpbrYH95Kab42kuS+Fra
SVzK592ubmt8CAojG6UBpWqhjrTw8VpZ7uat16X6SA57mdApm90bPc2UeT9kTOQ9lwI+epEVj4wk
NweRIUjqlO0VdZqlKmWbk5yG07KGg5ZokaKAZeWasW711aA+Gwx9tQDBH4aZCzQUykzsYrKke3GQ
OH/poa6H7Ikui9+2TxRnNwGxlhq5rOFBEWFiULfPVh8yqAhtRv8kO0ZorXXu2Ek4vdrxFpxxFuxX
zZos41BF2qxHH8z0qPcDh+dqJMvylvBZySS5bHb9linFZN0gRw8TrI1GGjRhb2A2zYmjcvqYPfF0
v2e/OfUynbNoVKFOECPNF3YHt/M4kUXgZ5/N53f77DY4RwMwrbztAqZ84xG9aosPt8qzfyVIxw/0
8MJsWCZhvPvKufmj2GAMmw6JFMomooi7LKPuceKxS+yJgq0B+SDzwf63XL6BYNXU/LG3KsP/aOt9
EPi7yeFFm7Y8dmCx5VPpPTIPv6nidEtayCnVqWDwp4y6penIAbkPwDgbbr3LtXfRW67XXz6srNwT
DkiknRTAzbB+KnAsJMlTj0FJEhVrf6XejlPS/U08mnlIsTWQphjrN14eTSpovmj/G7IuDj0pqJ/f
A7j1AvnH+6je9pARozZHd8zK97xKnOsl0xW3Dj4uXM3lHKiVXxyIuklJWcMfxwbjY/RmnHQAsyEQ
lOvhAtfM2bzfmxgb+cBa0mtphLK4tvj5OYla0JftETmjORelsfUqlSznTh4izb30gMVokR28Gb+7
Lt8BPDY1k1KjJGIPEwI/CQ8AtPTl1YfLFsQIDlB+TsltuqxDSAoyDylNsd5oR0y/zCQS80jBpWsK
f+NWz9P2EMdFwc5DaLjYwxt3OdM0v+yDxjwfParRdWfh6ffYuGLyw61lIRjPXs5Kjn7Z2zFyRdol
0smT2XU7c+P+QelZV9UXSjyorIYazYQUwcU3cnuZ72Nz9v/Ex6BAMFiy+xFR6bXyXBiv5805O16q
QOSE8BsIIw8DjhqFXMzYGrBapOHE156ux8vM7PscNZxXCE3t0gfDJcm8d9rrzJH59VmJyWYhKu23
7QRcASGeFzpiVzpHNmuf/SjTLiBSn4g/Z7AEUh7q1PStaOOKL8sUk3eZdDeKmCWT4eYSG5r5ZQZO
AVdIL4k964T1llG5yjtNoyjUiLrbX9WqfRPzva/GzeQjZOMJ/4s7NUlEYvry9lDIDBeuv8qA9AeZ
BAKVm2KoFw/9jnhpArLnjOHJC7sEwufYP8qHTpXVTbxciRn/Sr32P+5MmovO2njj1Eso5PXaCczm
0gGm4U4MSgLya6frU9YyUer0CtFCseji5djxNkokkABFSFNUL1T5bWnEA1U/F0tjPYAk9AFIjb/C
SnekDFJikvFpSitB3ANgTZZVa8p4ZFqxqRf2hGUmfbSnN/aNuaoC7k/CwYjqRU0OH4gxp6jlmovB
cX5JsGvbYTly7L80mcBrUaSj+bZAO3Jl2MX29Igvye2xs2WOE0MaDdQQ8Q/MQE7woTVRgaxfnSrx
kNC2ArkEo70la8V/qZZvoNcmjuRtbvE3nZd1YCye7f9w1o/NH9tld53Zu8t4pwuYGY3Tlkd2wC2r
hGU7Y1fi3POQwgn9GBtQxg1EcJPMRok7fCkJVovdIHDMstPcprkFhuzSDirSfYhuLA+hxzlFbVEq
12GEjBJ58eSiqMWQIXMYxW4B+hbhJawvmxUaY9mOaqQFdvcrzMReg+V2uwAnuIdUAlQYlZ4KWnME
Ezmyn64xAn+A5RDP9I3ste0ZTvTpKigBAKSccQ6iQ4IbCbjC01Sj+NLaxYRICiUQTT3PoOUDRshQ
BP8jZUFhJ4yozBAMp/nKbTQv6bLvYyIUzIvJno1G32P7GHTyuvOfd5OP727mKZq+fuZVX46sG27Z
MGazXcDJkNznrOUBnsJi0lt8+RitPJswEUhwXW1K4PhgzmN6NsTl4w+1kDe+kS5Uj5cfJfxFfvM3
gyGyepgLGS8Y2wSD7eS325GdNMSSIwVLqZdjy/XxoF3YsOqdAlFLNwayq18HjaPcrBXAXXpgusTA
6/VbAXxcrdbRPQ/O6kkoc75k6NpNEJFTi1avBm3tX8YGXBUL6QPgRdUCaAbxMUjc6fLVwrqlvAIt
qMH4ePSqGBH0+hUaLqTiPtKEv1taV9FCkiUZqURW+DdYHNQfYP8DKvYZ1wuQBwhuyL4IIIrjKpvs
zuymIpQz5os4sLsmT2pLZ7Dqv7IQUhy6MOklyCDyDcDf7lSBUiNYNCJG+VwTghgb41FwxuVRgWNw
NgF7McShID0y425rwk6oBFCYii7ftFjiqnYJQwJIc2VB/32U7FlsSvu3lnQRFAfZPWqLAKUMoqv1
8iICuxpvyPJJzw2/DLXlDae36WJR1FV3f5OectrgWzppotBWL/Q+ha3XbxAhnl5UKzsVQSGuQb8n
8LS3Ov7zkQWVp8NdLHUFHJNN+oAEBS//okAUiNIZNxYnM1sMieBjsE/hGEvum4/Nf7ixMOEZWFPs
9rBw5DhP6nWieT38BuS3WR7Od+TrU93gS0VQNaevikVSCxJeRWJh16d2AnwmjfraAY66KJrCqjOs
I+yvp+ZUgPMfhpF8ITQLQJaqEkn65XuBGkgwADFF6Cxd4Y3CpakBpudTpDjo2qMwgx2Dx2uxGP1b
YJGOWVoiCFQuurWZRQiIiyLBFuWkoCTCKObQHFq5lZ7tKpRT2zh6gTcxq9JqqQt1kXCLiu1pkkFK
rIwr9oRzF0FU9Xpzkv05jWGl5BV9h9gnDjzUHPV5b5LDRx5e3oz2EiLFAyvhJNOTU8Yc6PU8V1mT
+XAVPyx9DX0AujN6UgreQz5c/DSRDbXPlGU2Cz7r5GNANlekvHGJ5lZJv3IHbLz5NUtj8HMeKYmN
fMuwifc4s8s57wXg57lP2ZKL0foD4f6Hs/r62Tt7UqfcUMIEz5SEAcW8U2UHIST2Qp0zpkfdvmuv
dy/wv9m08Ji1K6KtdSbeDthaAikz+LuuG2zoGkLN0xlkXM89wQ92jQC5YdrYe50Sguw+M2gA8UKH
RqFW29Kfl7C+D5ZrYH2gsfP/wwtLQqTOGNWrqul9CnF+hsuY/XptqVlOWIso957OwooRlRz0FV/E
P4ETx3Vt7O1pciTXAAK1UeD2N0DxUPVnkyHGo8GJTU4aPveZJ1boWXsvqI44TnHnxDLbt38bf+qV
B4BUCXPKOzT27gFOQ19WOgSsy/F3fBBrHMXvhbC+OefTQgbcbUL2QGis4Y2vtQdUgNrK27nNROry
Gtc+rgmR+9Klz8Z/qJUMbp0c1jXZWPHnqu9qybOT/8TIclmCxM4gPzuTgMleXoj7IF8EYyreC3HL
QJnCcpiQlDVSk+cIDakdWs+672K6YBJadnHVbo/jog1fzCoUiHIawsbHNF9LC8FhcbJWHUdiTUHi
u6ktivHLB2j52dQ38tSduVuzXVHko62WxZvhWPJAp29M7dml9TapOSa/LD3pIjup5Sbtic8fokdi
bUp7M2CspsBy1u2k8d/krcjxWb3ghy/EAMhmvxddh9rYGqgCJ4hMfivjHV8IWqfLlDkme2kYPxVc
cYonp3FDe54ytj/9fJcBbspB4hMpY50zaWNoGjxI5Vzz4Zw5ttSSu8mx+OEwiMS9eeBN2sGAGxAO
/9TEKJ+YvaS0xF4G/Su0rcJrA2LWWk87yBd6U+71nN2j7Gh8v5xhDVzomnBnbfPO1Ic3pKvjsa3P
z7SkzgdWnjjTbIBg+/uiknc0h9SSEz4HE66/FBTOeCT6p274k85K+DWA9ZMilr71n+bn1O0f3ed5
8Pzb7MgcFQKzPqNxAwvi5672Q8O2zuggYaWw/QvNRhV59J4riRl1Njb7wXd+g5IWnl4FxUij94ws
qDnNk2rtxWETGw4KHpQJE1qp6bFF4qmQJF6pudbObVC/6CXy7EWd1XTPebhc/fIRAz0yt0YD9gPh
KQDDqW67SHeWU3KbzuqAjbNK3qqp2vGRcPgUPcoyQyquYt+y95smrsdtvKcXABp17vj1ctIrNvGw
tbieuzolQ4SbH0aSyZ2pD8ZumbeRrFqtB54Mg4BcUjyuiMJGwy+1Ey368WEVeYXWbd7Q2YsZ3LBA
pb1G2m6QNIoXExDuzBAEMae74fxFbFXD11IjMiiZZjvPr7+t93OqED4UFX+dte7qgwUURtUvATAC
vm7Uo3qcTH5AwXmNVPbRVtjSdHs9b9eWxzbf8Ue+OiyFqPQHnqrdUrFNnVJcrEdb5jH/W/z7Pfke
JsQU+BaubpgsFDNmAeEOAOsEkrz8LDTmcdDWhpAv5H0PdDApvy5ecZhqCiJ3D1FkarbLqZWo9KVi
XbH1aTTCJ2IPMojDskLcECsdc7NnvvYjHXp/wM/rAnU61I7tuXh8XuQJCLjLdUqSFVbiSPBx+drE
IaKMesfYwarIeFV1ENT14UCqglcwH2uXhwE6OY4ATQMHTYbN1qwMzDvo8uu9Pii5de+R99DGfy0v
xPGLWwgE8eSk7vkqmFm3tiAdziOzanCnvXAm5P33LjR/qz/bph28r2LvWScwqB4/WvZ4vPs5ctHd
R9NKswnIMyNZfpsbWEsoGgg9LZuzYp4xGoQ78uScpLd+KXbjM5akj4N0QlDlqWSkxz+qEpBPcIOY
tcFKmk+I4RkzOUswrADC96rCdI4gCj0yzY832J05LrEXAnYvjsy/7ul+tURWhkhCTk9dBqjkTp96
BHAdCE3ukAzlPZ8+XBna12kJVjAWg7w98N72wip/OJjP84zSyZ3zNDDBxBJXLM6IokyiRF6KkL5F
sUJyGVOvgxwXkURfHWvQe/Dz+p9iiRu82UA02OAtNrnN1Wz33l8bdaIU1boP4cS4n6OY4zLLaqKm
lSAYYGMuwRNFaJ7Vl4ExP5HRL5ialIHpOVKPLmppU+538VOk5SQOK2998IpSe7Jk2gF1cVh82L4o
EAJvO8j3AGigFNzcitABEry/jzPrZfGJJ9BO27e7ifY5v5PONjDaiHfXWpQ//JxZYWip7op6/ZNc
x8AUoA/3h/MZ91u2OMgN3Zt0AjLZJbodugCWsSTJfgJWbw9Xr5f8B1JaBMdqPSby4GyJwTnHQPQV
NNKhde+DoRs2CV8D2EZ+teVD65+P3UkCg9ENtyQQpxk5OpV1zq8CgdKy1IvWjYlVOf49pJW7gWMJ
wZW8O3OIyEEIyIV73wUN/jGbHPmDGFAVAzy0IBb3GjuksmQ/olWx8Ytbh8+l4f7eRAcORXtV1cJ7
sfOGZ5jqJ4o3STlyjlKM6UiYo7OODrphi5AxNcYQiykcQEGRBELPINsy2j0tDyyqisPA8o7P8jhS
VRz1lUzABVXDuaunx6GYV1VQ+JnkvNUIF9DjqB126yg6Mo7N+ctFPsAdmwMg2f1+ahYBYreYUzIp
C7SqQbY3vQSy0dDQhMZIVME5r1A7fnxVfherD9pVGxfA631Y4KIO1Rg1kmw/CODVx/557greJ0xI
ANzDSpeY5Zzk49tztOyMDSRO8TXZXMyNnBsUBZGr95iedacDU7IL+E3Il/1BiJCs5Y7Muo4LqFnG
z4tVKJtdbwc6HUAPu8CGpluxcJHUv/b2GbDUGcQKM+P2a0gR0YWQ+XAOsi/X7xCyI2qwqg+VxoNT
0HhsMHsz/K98PARRqt3RI9CxwdKm5GpPRKKc1s+4Uizo0CqTQuJ9iiILucQX35UDH002m3P3HnkC
xn6C9Ftcj2mIMiaU9c/WnFbzZgCGhq1I3phg18SPFn8KMGrzPyAGqjxzkClYXm7VsmarfKtU/W68
6wwIiKMvLjNDMgD3k3n4v+EUtKFZH3wSHxCqNUo5byz8EguU2QFN++tbH9IPNDfuhlh9OpkpmePP
TvOJcAjO4gLEmzwZXJWHTvMosAd/LxhjiymKFkA8lRv6k+EN26Y/dAQHhw5l8MwokJrGz71TDalN
v9mY+FZQkXIJ5LC2P4Vun9W5roGRw9OghcJIa8cyDOHHIHvGCuPVG6kbgtbZa3Z6nPq/jnslcZr4
DM0KgfzFiTSXWn2rT1XH+HvpSxzKZYbrPnh2xjhjn6vRc61qZK97fkZivLUAzbMomIJGs8a460wx
0shRqGX3hcWpZbjesKSMlN/6VuVoaVHt4An9Gslg2/Uj+pFUWUNxGnEz7i7jvFPMeNIFBfF5iZgQ
EVJnRzLZvtfqSLbncC8X3v3tSfMk3YapwWBQkCjRiHCEi6l4fmkqE32hwbcXxHydosTg8n7Hlr3u
a/ZWDNCqSkxcn9g9Ml84lNM0O6wuyB9x7inVGjrHZ27QPTTRT7u2uO1mJ4SBeXBhWyZoeW+fxxDU
GwPigQUOOJZKhST5wrwq5NG8SyfCGzxSq1KXJnbWzWNmJw8zXCHvemATP53kDjFFbaOnRY+mZzKH
cF3YlXvpEOlYqUUT2yBuo2EzI//FhVuoZFRivFKUpRpEjUpcJO1pvYNolNLPnMrK4EBMzhn0fJUy
+N/Dr9025heuhdAEyF2MzqrM27re1QxEA58NfVrF6Fq6kjnKWfKyOs9oz0kgReBWI+6IPtE24hKL
H5d+sOn3e8WuA1Bh6JqHtfAbaW5Z3nqChkE//u9gmIEbxXZvj8CV6evbP+/JyvFvWX1sXuNLl2x4
BFA/TudU71zXibWHUjH+p2Zn4OKJOnzv/ZQvuLDpxvw6lEAg+OxrlFeihIBN0q9gHSVnKiBvlxOT
weiTcOikI1i5HH3i9AlmUGr6KmO8oShFFi3e9vB8omWltFxrTGksHfFaKWn2ZoLb40AVQ4eDWCi6
JXfigZ/hKi/1nyZTWCIYrckvPMSBo5dztGxcBOccS1F50ur8swMitRyDSC1wYP6qy39v0XAd5WK6
31A2A0ia0YvfsHVOiUzTUlWebg12stOy74rdAEQrhf8VenApGWkSZyrivmW/BUfW0/9vIquTE1AY
eDutclTB/re8FkHSc1aJI8eMUdre88rVkROEb4Snt+CX9bybWRAUxigWjbfg+XYXhD7EwkHytV3+
suNumQAQoGRQU8VvJqW0XBWpVlptF4cR9ksWaH1vj8Ct8Op4j92QI1Xwax5CcfLk7gnaiiWzZ2VP
KV1GYiwNbmegIvhqRvv0XYppuu5S2UmSrNmzuCZ9SDufPzmPGrmFkf5czuaMQvQMZ9q/ekaP2X/4
72RvTR3Hh10i/0+1yvIB9lViZFgseUDeDXlwUVYE6NBqQKLbIK1h7OKiBF87xovSA4ZjXrOOetFy
7h3hRzoWXTL6dhVAg6fQsw21iaqlofN5zYcT0RfeRR+ucQL1/8oRpHkXi43N/xwohsAwlF6uaxJL
OQNjvSC8ONhWntIn/lEqsCR9P94hOp5Qd2eWmPoh90JgEazqrz/+K9EGm+qeNgtM5hZeTsyKXuRL
UkaAdhiKNi/Vi0T1vpPVUQ8FQTbbLjFDbkWUMjB6f5l47JbNdD5zHoll7No1wX1nph6fvThU3Ef6
EimjUnr1OeYBqjZd+GnTKEBU3rAKQb8zqd1cBzDlR8dyrwCDF4s6Nzd503xXETGEm1k/JEe3BP49
pXrA0Ef8g5ec8Fw6/3LRACoQwrch+KiNzXPKPLBZ/6ZOKqToBkHR4KIgS5FXU57eYM28MlsWCmKn
45MVJL+Q3+ShxgX0MYNpR+WofLfI6bUhR51HKo6lAaAta0Dh5nAvicqar0hagXv/rqsLTm3giCx1
w3XoJvOqeoq5doJzJm44clwqV0EcjFy7ao8PCz4ycpa2pMZnwa2VsHsWMivAVkB7h6Ba0Ki0qqUa
2FtduxPQUz2Yv0z8053aVmkcomYsfMWIy65Z5jU8uJhb5P+K1nCc0KlylXQFPxq382+z6zqNaEvR
YK111esc45bmmIqSM986i/tip1N/zX0AZYMaOJ2xdlaJcZnoUgGRpzxWwMZhxwoX9mOmmaEQKWlP
xgwtNSqwPHInjBQ5Vbd2evQZ8DJQj/0//rLbphb7+k/L5xvA1T/pESOIfIHPlwDtHb+pFASGSlCe
BT+P4R5QVSgEzg94lQq/wCMHNvYIUsImctPvXiKNQ7PYkk1qBpgjWOOLhqfbNc0SiAehIvxTZXZq
4SgihyPLXkVFFyD3tVEQ5aoxJUMsyQN1uS5va192+1I8fberl69jbiD7IzPzKyKgUU+MGLAzPz0U
4v46tAOF2oPcnTTZWihaJkv9zrx64hTNtUq0esnripggepxH4MEDJA6LehUcbsHQcRdywLZGW9mH
xhVwsqeP179c/B2YTsMYZgYdfaoON8bNGOZhCv1UVxu4FK+AkfxaAWUfoJYQgzjcZtqd3ZcBdIoB
q5NObkj85yeOS1KcKGBdr5b2qCBHQSlGBfBDvt/9X2+Zep+wZ1mwlfMJQydR2E6itfNz9jBKoDHD
ZtpxyuIiNPzS5Lcw0+VGRL1t+uFbsTH0V8azCUaW/p29sNgI4n42jOIRqG8icqTWacR9n/zF5RFY
68W+dxoKOnylWp6yMsRKfl85CYXMAwZUymwnm9Hk/Hctqx3Jpi4R0yYkCACXs7J1WHvCrsG0R6QT
zZrTPmAFG8VSjtFj0crXfSQ3b0QsypI/TrHiIiWVAEcdU8YlhXo8qAu5DZ/tTd+QWo1tggUAL6kH
HItjWoGga59Bw5W8LfyczCBGG6G4GaF04OALNZwdVO5H9zvRLBGcDQoytiXA/Nl3EHVcugzA5t1L
YHp2q2GSd0URvfav1GdftYiIaopADXDosaB5Nk55YZvnJQqZRlPaagRZJq+Bv8Wfm9+D+dxp/uu8
3XGVB2uwUkNgGHmuK8rGVevogrLoSMEYHihwbTVFfE243wTprAUeeJtg7csjtBhYGc+xxwzwt1Ss
Zs/e1Lj5czVHqJ8wccJMY1Kl84CMWVr3oFK4b+k+0C3vp8kzUOGF9q/6AWVwQM6MePI0eNVRf2aR
NP4GJK1zKvTEQT9HxzcgETEOgbmBKBB/NqIKItU8lUpJgpyba+brnyliHIZhucNjSO9r1w/0YD7o
MAr/B/FrOrzLNxeelvoFqOHKnxoKY7ciVitHy2W4ICXbPuWk9VADZl9yj3ORpGdSzwQNXVZCVX6d
U/jc2M90My8pHTDjZU5sTwDBzrZE26AjEea7KHH8vm9Pqza3XB8Zy9SADl4HNanmvCw904+ypH/R
MJJrQaJLK4WISolkRBmgi75m98+HUksq/JLoR9IbMBY/B1y9xqKBM2vpbWUrYFXCks0WjwRt6649
KTEB1EwaEMquNLl6UKoQWr5C9EjHtNeu7kAGJMhXB1xHvCED9h+EzzMZ8G+XTFsf/BX/bC1+ZIQS
/OyMThoT4+iFBdmv9AeREh0vmh5EieAD13ZMwsBOTmwTIcm3GUpeQbl8UJOLb4FG+KkdvlC3cdKR
5dgk7ZZ+hZSABaRd7b18GIr1TLIc6eSVhNpMfRxJmAVKK+XzyJTJZb2vp+Cwz8pyv+CtGFJSA0kl
BGDUwa3JnxnvkuHNAys3gbWblvS8WKLWIu6etktpxczaJ7Zf9VHUOD+M/wigEzbjgE90tNRae9Cn
WouWxAqM7gybRfY/AJ3fLCR3kLB7b036ODIfMP//j4XfpRoIzVzQBbOexoqXa4CZngbJQzJerzdz
zW4yN4lnqrUabtDq2+mzbuGaEdhXAyQcwbh5mBRHnb4CFyyaFgipdj9FOIc4NKpvfIEKRYdfAfvw
BegkZHzlrN0RlwIVYWrhRznCYyUSfJfKGJOjOy5tY8Da/aKaeAkJjhZm3Ge3mewU0OZauHrXdG5f
3A1oRtj2ZPufd/D+tzXLiabQ46U3tIa0/BYXF5Cw9tPU+Fbdm3AYz5DeokemUP6fqjXIVhHFkBnq
CqBN/I8fUl4IhTIyVtiJSjfn7MiHDvu2qq+pzkOqyzwBN39yFstn/C7dDCub9N+iLokBqyHGyDsx
4jvC4aiPd4JPCDb3AEsRBWHzeUCflVLOaH+OTGvYc9ZpUsdK/QDS/HtCnJFRbLdZX+r/TWMmFad9
tykjGgYjLdeZ0pD2ItcTQasiGTGxYcYTfxVBdktzppWvZKU800f5hkdFkD5wMTdu0v66wzC7+iZh
c39K4eiR0zTg8XjhADkHwVjIzt656YLlALAP8JVXQNxkqkK6mTvx9V0En5MqPHEZd/SyXtXvxu2D
7weShY7XgrET1vXSoKEGHUW1JlpkXDLSKx1EHqeM4Ouywrb0iHCpezSHp7BMBR9QGjMxgxan3Kpm
/gucG1dUkCPkdoyK3SbpnGxfiAM7AB6kOsxl7uEvuhkRKc1l+qBAA2SxG3D3VKs0eenBbGPXh8AW
gIt/LNTkbMMOs6wbOcSxOisH9vBRpNux/wmQNMwk60aWVAzKBmKSSs0ardRPVj32gsDCAd/g43V+
+0tGwzZwj+JHm2Oxqg7ie9RxkbhXppA5HuEKW6STNA5WHktzmEfo+uQxjmOsHZD5qt+I+E3BSeDe
L5gtF954uGMQp2JLuYHuRhVWCCA7RJSsotvXWCIVW157oHASG9DgrBLdK6oCfR3AoAzfGKBaj/72
V2LBVUk1LH8YijGQhcYH1kUsFsIIcM9egnP/XGOXn/fa90pwcD1w6dtfv9plG4iVCwBkaGZfxkPH
LoaGE4rseK3v25BFVDDQEFSixzvZzsSSoFiXuCIKoJGrrZxfaQnoCWZzgsqK/qzXyqgA5IKAvyYe
zoFmLrKVOKZUEgltAJ4UIu+V9k0VCsvWabY156NgfWxvqYR5kSmMR0ratHIdueWr4hQRjmYEoja4
N5LGXDoyOkcjKr6kK2tMKf2F+RInWX173r1jVlN44Qn1zqmqDGv3KFDUBIsJQ4jtMHdIpJWZxA2p
YlLyhEGSXbInUhp7KZCt7mkY8RBG328ZPYrsXd0x+6t9/+ntjPCBZjNDOcPwxb6H/LkO4AcIyTQO
vUs/GG91Ci1bMRGfXuGGPeZsG0mVFyiAi4khOhUeDz+PkuI75qDNDUd85F/BN8pboQnVqKf+MiN6
QBlD56EyWa69RIN5ktw06Bmo6ISR5R9KDLNAzDL5WbbeVf0+CQOKt4Zph7KqZY8XZtVZIZmsPPZK
zrCXsQdXOsc7/w1Mifbey+XILbtA/KjIe0aTb+RnBbtjawamu2w66I6/7MH3VdQdM401vTtvFTkj
hndHHUAqKj3nMBtmBfXcoJcP+t+p9b2SpjzEUujsJrBRjKKdRA3A9tnNiV1RlwykEHqiJ2nv4MMI
aJlUb3x6dG+jfUYN/6xSoGgjQOUFUvI4/MmPyqYUYgFBbbF1NPfbkStKi0TtI2ZoovvW3pPc7fyC
mxPbrHZNLR5BCPk5WrMIMj3v1Oqz0QGlTZ22UOxijMfTTcsUm9Qv1TwA6NRDisTBpkFXbRhVZW/s
13DIOs64CvAgxZf0fp5rxQL7Q63b0mFXo4ljJav9EpbuwtcYHSnq7nlMXFCvDjqnl1gFvRobmsFx
kva4WD4Ls2SLz5/8acRBSnFQkMG8CXf7WSBpPldAoerIbdzRws21HaReyqzarqsAzMpyYNipLqsa
nDHUF++3rmPcCUXQognlWmFHY7yKTyRA2Qk72PpeAPX2r9Y4oJy5uEKmRTrDe1BMR9nkmTeYRAgV
47KOH5AHIJ6nhutfVSF9pAc2ZGcQbq/408kxmFL46zliCgNYIWl4u/CJZoBv/cZnyqnMhooRslUM
+etDTu1olhkBNjLJnjpcw+7jTkiCqDlzxBfTgfnadaMWJcwlZPYeivBKSmJwkr9ldN+txNnqazlw
jHTsn1yT/rtmS749KwuTEabjtDV8OoSys33TL1EjOtqNaVsyd/C2QniCMh/yT0Dpy14F7zY3COrS
1+9AnIbSsXEwkC0egsHGuFQHy5QTiAwRBwv24qs0q5CRAVDXfBniL/5H2C5Dsf3Drlt/ylE6zM4m
PE2bxyARvRNvJ/zubGIM/FRtR1et1oKkML0+YzGaBL4tGHCWzV2AxxG8Jgyp+OFnpjv8It+7z1ys
W2db+4bpWTBfl+UVU1+Ya47LaSHYy1hVTSsjQEUhVL01A7gAXHONKFu5zob4wGUSBksKNnhBBVT+
MOCWGHBnh0KHtXrWqiu4VNHyRwN9XviJmQUs2AjR4I164VxDoQF3+seGCtRNtJDOGFmWxsMgsiy0
3fJqOJW9TmQ6tW+NvjUAQ39ValngghnfC2HA/oXr8/E/zq+ms3lW5TdSSPRMLtY7vHgIrPwKlwUo
wyits7tfyc4VFxH5sqIgCcZJOxuJo6AWW0LuTnIvvPIgI/v58pRNNWudVjGLZIbkUTIvcT7nrVHU
vr47/TSi0UdvM+n8+mnPHhpsaZisTiZISBKoQKH3/hRH5yJB+a3VE6f0AUxCglqiugF1eZrZaAPo
uZkrVJg+mmpdn8UE8F1p6V8+g/N4qeDb8jz4UQse1EcawVQFFzWs0nQt+4IVLsMMC7RIJq/pkM+8
2DdBkinIrww9rR9tc1DOhcI0WNPIFboKNduDvT4bSJDSyqLFKwWcqM/oNjs54dYEyqPno05v9beI
n/5hb3T/Uhep0Cx86eW5aTgH6b1bajy/I3fn64R8a8VL+9MMcuwilBav7rfj1Fm2WtBSDy2FOxgc
xPhwMr3BCT+qRX1tV0Bte81uaJDweaxZm8JFHgi92lAhr7nLodWGm3qz4HNTZTnOGIn5dpNOJZxp
PGkL2n5SRI3UXsmLy7Nn5/imViuTwKB/i7dXf/xoxiomoHayg+jCsStWtfnQNxofg1dEpD2kbH0Y
gdRJ94Qz9rA/ZXvGkZPPzVEsllcKrL81JqLMXKwq2tb0iXQ9RwRYiK7LO2D69xUBxjBFazIwyf8h
A9yOYvXK7zf2giXp1Ra4dGYCPH+dA8iMv5ANJmFZ81NSsoVSBr8//K8dKEy140llR3zZAUtKQjbB
L8cHbXhu1xz9oFXgNaqdGI3Cf2pdXsB46hK/UVotnj62zrQ0aB8LMrUJ3Ilgcpm9gShvCyusHMcp
gUG6BdmJ3UGnOTaxv1cfAnecrS1fGQmrDgL+ETNSkf4NhAx7TG2rd8Yp1V302im/Z07PYVwML5+M
nC1CGwN2bZ3WdFKoV2ROLgFEfeJE4MRKxyfbVag5X26emARPnAK70o2SstN+AjkY0Crw1Q9aefxo
UVsFkJt0aj5OVThwz2pRhl/2eyoElZNazv9VXIhuc2PnrSS+dCeMwIvkBsqDP4Kj0kqa7basMVkD
JYG5gyA8E1Gt2BoGoyRloDskJw4EMCBRnemgu92ic3u0fWMRY0PIRBM4nKlVuClZJTIb1LyVW6Uv
hNfm6J/vO6eU6bxN8w+itnBgcoMC2ugoCWtZVlY1R/DLZLZVfnQvGm1S8n/sWj+TblF8GXRKEJER
A5YQ7HLdJorGrrUxi4wCDF/v0D6TUXr9IDoZyKAgbsVk8tv9SOwppiSp2W96DwXoM8EZLM4Wo+hO
q/Qo8AYzt9lcg4VPgpV8kf64GFwb2wFdiHRDG1jsYDiUowz3tgG/DWzSI8E5zBPo2taVvVHSEETp
pKAL/UYETS3+zy6ZJ32Xz/5eCql3W5a+ZmDj6Kv62427iPwvjgGcha+llBTLAWJMjjdfvLUKw2W/
SIA7cq5J93Huvdet4+f8cGg7YTrmZbL7v3yrZSh/8eV9ybJWotCJnU+ak35tPC9NYiGtuOg7BLlL
PW73rpvldwnh2QBQg4UoTDPpkQGBxG/cNilHGGE3/vCe41wnXnQXmrY+vzBNyIMNM9HWq3GWvV1p
YX0COb7Cko+zra2Tde6gqP7wr84qXoMiKc9WcmbNgah11WasaOi8P5abZJ2HFajxDNhVVh/YXjY3
UDuDWT0sKhBzcMTnR1lRzmEyNFSF0xI0Wx1Bwtnterl51fhe8WJgB3DeeOI3FIbBIsVoo9u+/I4K
O/DzxCNN1IAxX5ECACPGVAT1yNDja5muD818R6LhZQeVSpOsn6X3Nzn2qInN0TgfzUO7jz7E5B5O
CWQG9kEzbnovO+KFgRpz9EM3ns90fhlgB699GW5KJBzLmvwXf0Rs0HvL/lhfuZFZbt7xXiXNfeqO
X+OgOylnADVuouTDUNVv0fy36sae3U8BIi6iMk0DnESYxMwqYUM2+5Lq01eBZWofp8Fz9KHDIYlj
Cv3Cd1iHEvSKEdLOyuA+NKKxNrLfuY07wvlT0wn2uBvwYktMG82YDBb0WPCCfrSVz40Fxp7NR4rv
pxgpY6WX8WQH6Qu0Nn9GOw5zqSH4IX18iPHzdbqh7WYbslwseFXY5RUm38wCVh+fMjnkxHHld7TD
ZRKL6JkFiC7J499OO+aWAALNQWbOhW0TCCv6gMjNRs4g1fxbalyno/z+F0dSDSevovh6uPLm8jjK
CRMFBVT7I7qjAlffgnv9YK/4LUlzgIFaw/H+768ilo2A5I5QC20+tPPkO0ZcuhYvPmBUqw0NHoGx
AWO6l2NnKslgh5HeNYkCb4WDwzPuxkc0BwkZUPOGInhl/zvYG/fg2hIZqQz1QGEa0KOTR+Bnj9WK
1IwQ7sdhqluCbGmYpcC7v4izKNhQnbv9GF1ZRlTl0TMLOoDszY40AuilQZRIffndQ221j2luuZAh
k/+1EEAK6w4a9zTPeewkRdxac1G1bNjdCNa7NRhBcAhHsYx5sQdLsFWZBdUJn7CipNTFhQGNyUlJ
KbzlUNtx2WtEn83Hqest2WRAkE383JCCX5irvwpH7473nRTK5USGKE1E/JoP+C9AUPdpx5oR3SKr
OV7Dc85bXWq0AM03e3+8l1c0BpuUsydnkFK/8Bq/29bE2vVWDrSO6dlmSzWwFHYy524n1HjLKdYg
kVBL+PZIEs9H8JyqVm1gLbBBkWnKLyPU83RbRb4fQosNT0qku/4/DbLB8oUvCWkryPxfQpFN2VP2
151R8jpwl07Kr6E5QSCcLaHoaSN8DChx/Ep9JbHf5Bbc3jR9NGnhDYwGzVxNyJMSaN2ib/GpSJxo
VE2/9DmFGX4hl0m03alQRL+O6PI0F5pfuhRX3r3IzRxaR0retgeMBBd0/ftVewZhmPzQ79CKej5H
hyFi9DytSpJSj6BQOVKT9RCDcQjVHtA6672lyx+OLDVctEbdkfFc8zXkh0mVyC8rEYCuNpCgOjFa
SvoykDTU/Y5Ne0QRo41ZYX9Bw65/8jx0bcbt3brSbEotUBWLiJjJyi6nr5adqILxvOyPPoVO+Wf1
hqYes2UcxWlVxMbNU5hAfbIZpK9qw81BUnHfhcmAHFcyHzDtgC97bTrAC64Q/LLhrJbwhQ4ff2tT
yLH952p2HDDWXnMoRvCldSSLzkqgw6VWpKwzyXqAzh+POcgtnMYCsMZuWWV5h4Qfu0JlUdfcCr7G
MdUFh8hyH3Zf1ENrGiSBw4l0zMR8BJWAByys3YCohW6XCaJxCArern/C6iTkF6ryZyjCQvrFF6IB
v/RLQ18Fx/x/g9B3NxNR7qixKs4ZfhFY55y2/ReJ5OIvAd3lIUWqdDdZwK/u5g0a/le07PzjbvIl
mt1/qx/nmh/s5Cg8cdOCWJfWKuZUrMHR3v67UCMw1YCH7vCC9bxV6vDLAd5t+1hn8Ul2JUVZANAl
SmopFn4oQN/0EctmiWXQ+YF+1TxmJfiEZrDnZvG6FKjphEDrT61VfE2usjQT/MMMH4u+4Nftz2ux
0ofVC5K79djCQ4GcEQ3IjpzMk5s2wBBHzYDalNk+ubW/Uqu5otXTja/Dl/jPVMIRGlvfkmprnA34
HkNCFLTJwAplC0DvM92w2xMr4uJX4q6fYOniLTB6086IXfwYw0ARFsJCeW+eEELPDPlrfQ5w/YNf
CriI4ja4smUDJZENzkm6o3px4OLdsWLYLkhuC8tYONO/du+2VJ9zV1tWuDMhUFeCWJnaW+ezt01H
KRP+/2+eHqhmZXv5D/i9stlRfCz9Corf9cT+L1N9Pxdwm1/RA8nz29QUGiFUizfkh0GqdwV7P7pl
Qtib8fDGLiE5FBBylS8GKUoJWfFCadAD1yqwq4Q7hQXttO0hN9WaKG4cZO1UHqz/X9JysqCYisAr
Htkp9kgftw+u9V1laKWkRCTpPycqIv9gqQE7D173Wwt4c0sLLXdBS40yf4+NgM386Npad7l/g9fi
TxHhcmZkE40iQNakzWOYcn6VXDhT3w5NKj/bEb6gGparoQanbFuAqqmHiUzHXUTWijC09lNnCmbi
B6GfrnByhRTbco8sK3AOyAjtjYqiMvVhMMg90Qckf0RRkzkz0SsMFSCqJwEvQKw/mt4sapQ4T81h
AgtKnkAaBx6RDzeCfd2HVo9WDvo4VNvAKAQpR7zlMMvZy56MPFhqj7zZfNWxKzpC1Y/Z42J+VZDN
faQjTyjZZBbpqXGTfzlGRaQsSsl2xBswuktg9CEq/t+PsD/6LW1BHg7QI3rrcEwxzY7nFSkbMuw8
1wGD+xvHy4GKq35bvo3mWbpLwcfxag4HA5ZXp+8W0Q/thLn5g6/oFRXuuLr7zkGLpwupDnfJTi5E
Bsbxzpu3tsUAtFIUY82c1nrFRpgHXxcKAsXl9PgG1tNGS8/eu+H6xvY2Z/h7WQDDcvNfUUjSyGX8
PItMn4E14OKpGqCAd4hQuGQfErrSDjJW96Y2dr7jDwRPR7KPPCfJwyYof9VZLzK1Q9cYMzbXywUm
WyGx3Jnp1g1uAvQTZJzfvAY7RIbhhUo9bJtny+vSkf9QsLsm2y7mWmgbefmOraOyWlmrjI+Mxp6R
ZwjzTIqEyzFH8FVOMAAEqYFxpdz6DcakkCqhJZbKakKCgW5wsQTQ9J/PuMzqdX7Lp2SlOZ3iN4Mi
mIDj6urzFEST5/yDTETJy9FltRzrZyuFKzzoKt82ri9JsAB3PN6WrRtDj1gO8Ss7zDQ1TJKGZRAP
lw1w0ZK5ldv/RERxH3Nu6hhJRURP6tjzwj0rmu597gIXs1oxHZlLEOZM/9wlDqLqGDtJBi9+Ibj6
KLPI8074Yvb1ULwOQ7LV/YToh1NGUqbzcbNTafaCM3h3R600iu361S23zEn0SP5D9fgPqj+3xIMt
X6nIfBxRee+CffBBjWUIEZHbUfUWRb+H1R/ICWERsD7HN2zSIY7hJ3oF0j2t3uduoRKY06+TsLPi
eo02iUmbqf3mXJ1kmbz9ijRphMQPRbXIoy/sAZEAG1srlxt2c31KfXX4pvdHThFsLzsZ6eG64J7/
pXudC6NqzJDMMzSNK0wi3OVOLv5YM9CJGEqDAEYWGe7SbIlJw5FiQXK24nk2pV4SnAeFcALQC2Kz
VGfIsfGerbfayFtcHBPKkBMPIujbOCflL3NmrMWudCuIJf2nFIcepu7IuskLyXsTLV5UnM9ShRe5
rzsdLy9ex0t7d5SJoaUO9TS7QbiBwgG2s+kR996ZeqQpbteGQ9v+qNb9fcGHIKm/1ONW3klSDvc9
Z98R2ApOX6/kq/iVVqSVI7BbmhoCY1FBO0B3uBUYmGobXNwEimUKi7+ut2TuT8xzQkvYrMoRd+nO
+v+ERfpG7YgB6HSVMiq55CAppDhVG9w8yyj7IIV2WjoMMDEsTGDwfGWFVIogOiHzlS4a6BYHYlne
ehmWY7hBH0BD8Yt3HLJroEFVQ9D4soPtWZQRWECTdN8OjYFsS1NgGLwwPGKH10ZiQrXRXxaiL4fl
rghsRx2CN6xspMeQEy/2cdyJIeQ6JKOOa1nOtVNcKH7dUtingqbIFhzRNdtGo8WYXAd2KmfMVyRQ
xma6nqYl6kOITlqAkJrl/GTEOHGsKFgfhMXNZc6FTfVQnbjNDiPPJBap5H2cKJg4LHEWlvRLpPPG
rff7jbvvDM5RUyubg4BxxC/ts4bpq9MVu1kiygIccveC5uzXyDVeDXzWkXKPEyAGDYH4VqvUof2K
VQM4SRAgQvL/U1Hrf3ILRS5+X5oBZnhdnfjHaQSCHk5ImXKmXue9afsBbwwtgFTezmVAgUsWD3TE
tjA9WWDz1mr9MjKqOhKGbbv/HR5utIe9BEl+sNcU/unHpb418AGAOSgPBiPsMF3GfYIpsL2KvPJs
k1REjNuJN0G6spseG7fIwuk/aFkJS/r/pPQgY7/YY4rX/HSQBwf3f8lrpU07v4LjyPiz/5l9jjXP
C03mmHBOqTVo70avv/O5wDfDQ/6fbTaMVqEmMb7Gjy9EcZP/d63maVwhvuP5lqrF2gX9SI3szsJu
YN1HaW0ftDHHtPatgrbImUHktbw6KcZzalufpK69hD3mfnfdH7nKLsSFjRgYJVlxHC0MX3l2W2Nw
58Cu6m1I1I5r9Wu0Df8Wn2klAKHt1vJhOASa5N1EAerEaz6R3D/E/lg/nL+rHGpxGrVTSMeMd4HS
GiTlqcMkr8zVLsyWVFS7mp6fV3VFUaDahbly8Z9+3Hzx3I85b6JCoPMwCGgZYv7j2gdQcPYn5Ole
RGVDPAKmr6WiMfKSxki0BkMtvoRJe/P4ZCEWPJ0eDXFsd9pQKvfsL1jOpVuFgjNWFYqUWkPxbFcq
t+NnmBjn5ywGkpdH7HiOWAeVq4RD/YhVaAtb217xI2FmUwWGZFFaVKPOaW4RdjG2Ugian2/4X9XX
OOCbUHiqZ83rRKtJpYGlxORKlbEY+RmhSERfUHQrIN2BjOnDMuHT/DRkOMmO/UbkJ5EUu90Hx5Xh
ZMJTvHbXvplTMvieckC3gc3LCb/rxzXTvs45lOf72MHSrcR++0C7XJdkKWiGhT1U2y77hn/jw4GW
ToOlHqdmxrteBiA75eoBgseGJHbIG1EjJf8/WPd1JIY3/6SDwVorGRuIj4MW171hDAOAOfQCnOSo
CYT7OimxpXxHt2Y7USyN/31fiHyyYvZQDssUwl3VWztTJVyo4FqxcUqR2vQlFaTsIqIvfCh9Y3fg
gfEMFPC4F84zU0xEap6Zj6MjmegRLRqbjkq4h2wkyRyO3nBnsdvst/gZ1amyYZR5NhEEPqHOPt5i
IHew/ezWQZwhoRMzdV9JDc0iG0+yefVTN6IQ0UNVtg5Him9qCkUkqmZbI874WIXpU65671YqJYwS
PMu4GfVAtsa0p0vj6MhG6qJkDao5tJTsRPRW3BETCDPpdhR68EH/qbIng9rScUdCF9hYyozZuDKD
s5hnKhGWmeAG/FJwnBHbAskhv8nZhAEfxENItk071rUlMljAWqUpseONUkEozgv8+A/XPuJ+MqpE
ShesGvUxMU5b4FH02mo6bHK7tY0IltS65i+OysQGswSfCT/p3K3pyUqYcog3gxGibZXgYiTZzEr+
Oy/XRQPEup7FGM1FUscw192OQ1nBt5gpXfosuNP48ia1DnuxH2PMsKTLzdylG5BgTsASLMAzGvkX
kvsfwt7i78jrkBTUz3xTUzxwLrw9pI3vQX5Nfz7lF+VmTMkO+L/OyaocMPRSvqWEB2KK8RNty4Eo
552ju3YL0vp1y4S8oVXqz59Zo7NVMd0y7JhEzqhXEg/IwtxlCj0Vi26h0iOFm0jRCAPzo9qHlF2V
PLhmdzFje2JRiUH4JUFhsoSAqnMF/P4FkFYv9OrNSsmTAk8Xuizj0MJZwR/+AMXg1WLvb3N0NsXv
AoEhwLglZHkOdNE/ZBC7rbBteNn08q7PEclNOMqNQFNuOKbefVfUu36EPkl7iiIf5kK1Ea29imTa
SVMw6iUP2I/eg0HXc94wqPXc803G+2vcadbnOtib3mIbOlKY8pxIvtC9preGiraqVO+7fzYQ/+3L
yLZ6LJIl8J6sz27TBlSz6Qu3eKug2BXOKqFEFu/p75ZsMJbL+ebDpDi77YXHXaB3KLDRoII6zTuj
aA7neH9iSazWu164LZO0LlAYlYKo9GiZ34LrOufMntM/rQFnisW0oZ1hgpT1mbBwD5qQ/2IHLy0t
WfnOeTe6EgpZ7vBeR/hOe/TYNtwNOThbv5LPumzDmRwOqzDBfRAAbYrrSt2LJWHffh2j4XdUFvhQ
a1Jfl3e1NP2HZzywKgM8iEjVJPQ8gHSXTSzNXUe7E1L04cmiLeblf6kp96rRGNK+Z0qx1xhYW5gi
CK6mIMOOnELQDQTnD1hiOhDuXrlKOmdYbm9p7hvxITF6gyXPUQ/ox95pLg6O95ABtS3h5UmAX9af
9gb8H6Cs++T+WKkXXYaxjAYgUM+aqVAzAYNGh3upUyicmxP7gTghxwGX7KNRU5IpaZUKvykJAjIH
7ekWMCQPy4MA2/2usqZGosJJhiQq27VTilkPY6lm8Nh21dJob4wS1uVTLCQ5fv4x8+DqNdWovsDi
P0GnY9/l+oMzLmeiojJHNnPVLNYQhFGbkakZJPWWHt40NMyf0TJ/Ox6q3hvCIdpUGki+Als0DILA
oT/ua+q8NU2SHii5UeHcM4rs3w9V2kCiWt0nAh6SxSKiTQADy2Hv6orUjkITID5tyWfcVJFGUrin
zHO63denxe4Tkddm3tNYDZlbN4jgHaukndjT0hGRfe3yLLWawiW2EfmfSa/R32Mw0v2BQubcCWUl
oCzwwnL5W1AuRMILO7r7AD8Ws662ZxVeHlBAf1RKeQaRQXG7ozl7hUMxKwNTvJOboQz6uk2ku/Sw
i1RPHpBFol8nXaoGtKK21U0XCNUVeY5opqYIxHhKunB/h53aj2yq1aMyGL08t7eLAytnH8838IGd
LLtVUuBDUovpBee1XZyIPbYmefKub3jDEeN2TI5qUhrci0CDftzNm2Sv4k8dXzBWDMuvtkGSpI0V
/pfGyrhFe7LmD728e1TZ0usX08822UGLShVKa1IUjfkuhzh083ZnhQKBgW7gloTtzpPBu9qXVBxe
WlWBY+KzILzv87t9DaIli9Zj7p0cnxBJ2LW93f6Ka/B8oDqdT0KrdV4RTKigPpjWu0Vm5BWKBfXV
JP0rwyfg5gJiLojsB1ZRd7BjX4/a0m5q+2SykeIgE8Z17ImzyLU/jK0m5CE6TErpZ92Q+GvSRZ69
gA9KIyim9UxsmueQUvuh8v/PtmMrxahmJNLyHLdHvSBjS0yoCrkFUVoPq+jfBOjyRKscArpM3pAc
8NJ43hnDnrMh5m9/h8//BSN8MJ2w2IYI2Fe8y1QF4bMRygXbnt4MvqVlQdvGH/hp/I4xXFiwOybV
cS9G5PRR/PTcl1zT68PeDnZfFk0uBwkBMlM0t93JgpOugtuUWlkeoZNrtf/17f+nExB2mdTZ3Ynu
qgIasf0N7darixiRkoky2OTLXMwKem3ypJgY3457cgWzWZsmXNfzfa7YO8jtyNZqICcTmcmnp2Ie
W50EINweEeKdvVIair1YjZYZCWLwr1zin2lR99wfAvv3w+NJy9cM+gxF9DL+cueVb2bfh7vMXIVW
ulwkuaSm4Fjy/kZLJRIwIeTwYO6SFqeu0kYUqEPhQ+VxXxW6kqid04+2eBaay0NUrMOqyyB/YcSJ
+Q3MjIGwOXzaWO6y6IgfFGV5DDqlzLezTenTVvLiN6bJmbIs9joJikzWdkTeJ7LMMI+MfzMRqiyU
16oncE6FrMdNCIl3f5o+W5hjk65cj+tUjrA3RR/Qsk4RSPhFWWehb1jwUzHqgpjZUADCF0D/qX0m
CLcbPsVhbrhJ5MtCNKJLw5gsl7dAXHjrtZMlXkDBr7H5Qw7+MFWP3s7cOo2BZP26NPkHmt5LdMaE
Ah3m/TkDsghm0RiwJ1z67GC4DEx87F7rSfoZurCBTGfHuaXzXwjPwvN37ReDzQcHO2FPaL0wmYce
0q9s+3QRMidMb3m17tUdUIxa92w5Dw4MRuLrtrCCqvHEmg6HCiMDH1eTPAfoqrBnTeUToazv023Q
DbPeevr/TcK5KpJrRNsKJb42hblLmzuuSe3Ul4vti9QXnVBUnPcQnCSfqsXvqB2sdL1MOEit6rmY
+8jHiwE+y+ivAMyVM5gFAtAGvmknZUiAWSFmWeCoDHPpzr1aCY0kMl2SPSexH6Bg6HbkRVsDq4RN
lq3OptcrUQZuJ9PyoO/KseULG1rq8BEWoxiCP06QmCSNund2NQaE9blaqDewPIKbytaajBkbRJhr
T/8Mic86cxffG1QnV+CZotpaXplTeCbjexTuZYBUHmYpUJFET9q1jOypEqI8hSxTtbTs9StrWvYn
vKD0p5LkSVbuB5/Xib63dTibsTSS8jd/UszEl6P6TyDgupwfk7vU3y/cJBvYHQzlR1CxNL3v8LWA
+Eamau3kY1PZ/pYpLfY0bvOyhuoVTnywz0TqDvB5tREFc0djbIj7FPaOWjLveHY5aElaBQTECYcC
rcyqwCOnXgj/ntBB9fS/v///WlhYhBEb/Xr2tWzsd9+gtJKI9kr9wQ2WcqpAhkyHzJU7B+PDk2kY
WRyl8MWGJ932bAxQbWch4w9dPyoGGWWGVvvh5wXPicl3ggO8+EiQG8kH8jnmqtsLF+fB7XKzj7Zg
Kf2nrlQYeBCI1fFiviirG1FEnzaiaOgwwGXiU2PLb+dHLPFqU3ideseQoXiBTacy0omOceVoZRZ2
hnw7tOGf4AyQPNtuVQDMSD0qTLeu3UJEn2Dcflkzrfon9OwNIATBo4qJsX+ks1u3Q2wf1tKwLD3P
/rczc8qF5DBqyNITbgvk6k7J89HJ3vi/G0kiYHpLkX+qC4tRvGT63FaE0g4ZVadzOv8amJ0R7GV6
pBkrFAw6cQbcNN4Y81DPl4xkSBk4+tGhl+DM+FIhjEp/DHIGJ3y4Igk0aXbypvPn88497PGJQFnW
zShvpRkbNB2fcM9TWigBDBylMWur+JuYm4tRIiF3WSz3QOr8nJUDhppPw0wNB9rLTlBZb6JtpP6b
dYMSfO/VWxcdYsUHai1pqDLiJkLnjFBC6qo61QXG7NWV7gYh/OS9gk9uTXmF12ZUUYLxcYfugKdx
xB690vS26k+Ez+reWJL9eTV89VjZlr1jE5HJc4p8s8Mwpt+/HzISXgnZnYJRXbnBiQX/ON8nyB4i
K6OHeo7ua2l+nRqSnG0sCe44UyeIP9QII/0wUoP8owYurGNB2nDkGMaYYt1xquS3aZUstiymYMNi
n/ZgnI45hVlBwtH1RHfn82CkaUFeS0sPTYXJGK/smqVk7WKoc2cVBZCTBfi3gFEECXT3COK9dAq+
aPgeYCSca9AZQknCH+lLTKp0Xh+uBUj09x/U+net2FOoT/zpZu1Jb3yV/2goBQz6qABTiNw0LFbe
EKCoKc/onqJ+bGxn2VDPbDOsFbOkBJsMKWmgeiRTr0kSKeqr0lpN5ysvz3uwFTgs9IKEVg4z2CFy
kX7YvsHFsIgzw/+qWXEpJdCADVl/tmk2YVNAGI7bhxw6fHqk88Q9CqGHCUyimYfviGhtlvvElzr1
JJ767L/l01j9u6eZhKafqV2ntYWF0y4dtO2etPNPI6QBS6Fxftt+oTPZQ8V6Y98c9NU7erL9qSvu
qYgrp1PM6w+XD/ui8WneQl7uJNzwQLi5crokBhMG984fFxcL6fnmOsd+7G/v50jENzPefRL2PymL
xlSobWHWUAF9U9hJvLq+ZJQlDRUtZqNvnYO8DneWfo5fVBMUmydsCbUySEKEvxdEvybEmmx1CW8f
YDQowlBjUrZZS9fV69wTTrhI47OKDoa2q75gfHUSSgIxOFYrJolZTJlN6xp6uEBk2iuGNf7BYGt8
yhTfNLU6mAoXf9H9njxCr2m9aY/j0e9gwdyAcGywsT0QL9baZjE9KDPw9niw4rDa4ntvfFYoOM2x
Lpu5EDLEP7UlcmZ3xQRVPOUQ48dNVM5jLfwkdQRbStClboqtG8BpFVbVWGdhLoBvy7ywE0a+/feW
KEf5r6Wgh9o3yWtSzRps2E2LjaCiFsEgS4M9m+x8r4bnJWFbIoMRaIEPpq2uLxlY2pzdx5w2U4vm
s4pXpKeTK9J2l9Zb/TZ3Qf6ZEuulHcAWLRUtrfS+BztbqQ7TWcEuqTqLjnzc85B1iWCdZTAt1PAt
qtILTCT8jQ/jH4t26kxXSYOZiqbt2zBsSowolSSvV2DNM3FDOd6e6anxAL5GsV3GUOmx7TAp8aQ5
hYU+3dRHAsn5nrVGyJk+sQpQABfpP+2X4Kua4mdFAJ7bMCD7ObwU37kYqCuMoNwpDRKMg1GyaE1h
IrsxzieEXPeHqVpmq99RSm/2+neh6I1jfGY4KueqZV/8bD3tidxmRmAEYZU4sLSETYRT27bHTH/D
jtnS03XXdJW39DkVrzKCawIkKtCg0v0XSWQAa0jl1YRTShJljDvBULYqTOquhz/KVY9/enVL7W3M
KurPtCviNYa2vpnO6A6c6tjhuciN+3/H4tCfH3Hn8OOYn677Ih2G+zHGHmo2UMZ+6bV1OrhsVI02
PmJsTm/cm+MlvIxiPdXCv4WPQdJTXEY/I8WSREsmJMghCoUWnqcIfzip6YJcH875DuDu/su7KAp3
7iairLMe1wdtuKRCWyRIpfEcV9rmiO0ooFeB4/BorWehHjn6sftpIB+xARTFMhlal1bwX9BO/PI7
pJ8efaStsfrhYirf+IycoQY6fnqAy9MyB4n4Z3GJylpnGM2K9CzjXC1I9dDC44/V5cyRpnL4+Ad7
KBLl+x4izvyhDXPWHqm71n7YlRjnT5sRTxerTxWWZfPFN8F+NSUON/LnQygi1Md3+xPq+woZJfCs
hiAZwCtwfa3qBwEmH+fGJrAmdkzx2RLb16YvsM5rtNKPQVcZtQfRW/JnBrcNYip/pc7rirDTdIQr
ECVhZk/lWlA5E8+0VRmuwn133oNjyW3qbAA/5yXBS/yjTEdNY0WN/y+dpIhgFipEleb5l92Roen9
/HDYSSrFKcos5DklUe6zg/PrFtszwVXzJjgmTtaVxaBpEqldOnv+sM9KfLwcG3m8E4RIt+caH2fp
TnE6LkAMkQOrgfhMdwqgYd/NkN1SH17p0Ax9ta5q9h57x0xjC5uOo5ZvLpKHpKCJ4yOgf2PCpNGO
IkSJ1K7yMueBhZiAfyx9CeGVcYU6I04+ZUWcVW/lpNfG/6YwGh9yuKDY0upoVvWGd0SAkwwWJ0Iy
wdxXj+Xx1wPVRoP0PLo4jKCYsY+wtK92aqQSofKiK8wa1FwpDTcf7P3GzZD+CKQ6u8lTfcn4ramV
Z50KBkov+HEGiyRcxpBEJpVFySvVNNuPhIXcwv67EkB/kttBe7MZihez0NbJ3Y5J3qqxvNVHrwnR
M42gxZ2HlUnnmfuYopO8+PkyIhHrE7nlsBZrfDRHYaaec0Xczj2lf6V07SrjcRyr7G8dj6baSRIW
/EhPgl0CVP7Y5KJRNB5yORBdolZDKxhceec7kgg/UgHVFiKCS/ooFcD7pRY7ra2aM5CPogYXCIsF
tzare8ae8z7pEPy+aIBu4Uji0HJ1E8J2C1qZd79qs17+Y3SRTNtV8nW+okbbpcLBxnHTPlPixDm0
oKP5Qw4xQQBLa4O6uuSVlopTdhGjGucXBpgkL1eYzCRlK+LPvrA0cDd6E7YTK4Z4eabXCvM5JWgi
Or35vwAaj/+fez8edDwj0qzRNjOui+V90n0XXkWnEeLIcLpzqkQrmgOERmJQBuX/SD8cWeMyP8QE
mCzRmqvueBdpfw9ga+ryz/VEDFZT9VoBkM+VN4OO10NLKswJcKBY94SFVfDkUJtXUnWyC0JwMKEq
KnGXGHg/RklwZKt5okRycYgy+e2H78n2devGq4Tl9UWOf0Uh3tN8MBnThfsatr6cJ+tjoe5zx0So
1nXmvPAHYzR04tFWSmvd40ITP0QjaL9hlrswSFht7v8VrzNpgT+EOJ9266U02uI/GjpFQhdmJGGg
/e3driSmiL7Mt9J5Tu4wJBSveEieIFlKmmm7QNA4Z86e2V9Nvzbp5Y5yX0aEGI/X/pviXJ98vsP6
y+sAYj+MpAtdK1/mrH1xDVxuYZADxDKTMWZfEUQZtuZGnDpt7n75qz6tsmXF4mVeOLffaMVQDvHW
CSrxSJNF8iKVMjCHF/fX6RU4nzl1Xl0K8zGio1pIb35McOyuaZBoMm9JTguBdAxUF/qJ7uZH2B+A
rYMqzyKjTvsrZZPw7aQacggXCqwLyE9+4iem4orlmB3LJPZBZLnzYcYATNqgiO1zzyArbm/X1nWL
qGZGJycEFssEdPh58doTmrV++ZYHjXmF12anVI9TFgkU7sRnNfATzWXKMrr7vrBHu5OIC8sbKf1M
Yp3uj395qNFEx/uf8M7ks/cAscASR6XwXnUBiFamoa5OKuuEFhfSlpVNiHH7SG3t50HdSpv/Runj
RiknDYrMTUuzoSlfahtfORyDQ9EhIXGqGLX3EQh30WRHG/Km/ham1dsCcsxchwcLtMy+yc0ENHzh
hSnIWUj20zpbHnRIstJOahbw8/vL9fbDHShE7PnZRBTZZyssLrxBjHxwkgJXSFIHpodGtdq+yOBk
PVzOyOIJD9jap94a/GnFiHs7ppJTqU0WTnj5v0m3ihVWyFYLcUsRnHcc5YxgUFCs44E1ozXZEsvo
L+jNj7xOsKfflmfkTqQVN5EkC6nnVREqjGsufPHhOeI6X6R1GHK6GsMVhUg/U3erC2w2/b/7BEqp
WdJHuNjJ5yKEp1u38AZWkBNV06UKbqWqwL85DJqqx8mKa/HZMV1Ka5Mm6441fb/AmmgJUM7sqKe2
Os/E/TGzCXvoPhQlVpnrqgOfKezaKbcI9gBxs0OQQaIGiUkfOFnIIKu/fm7lsK943HPpENl8RAMp
v0AipbT5sQgPCSn2yJPJNANa4vEZN1/3MjdUWgToMBQ5SmC6mcEbH8XQZLusRWycZi33uK4D8P2i
0w5fzCEfwdDshx6/JbN5FRZkCgv4rZ9boS8tkNk60ch3OcdZhcGyiT1m49COrOhnIEazYV3Qn+P/
yiQ5Ed1PpRJ2Ovigs4KSzPhp0dEhk+zTCfpRDaYnHORCxXshYr1fy6ZRxG9Fby/YEPnfV8n216/O
bSEY2vs98WXD6cvDs+UVcdbfgPiNmcNGvdeEsqhNEAQqo/Xw6bU7iS5sVsLGOEsggV3HvPlXi4OQ
/TTXjo04bxCmEme9Ou442bvZN9Y0EFNVlaDGnLG7Kc18KMtT6CtfV+kABKqoUyV6A/0jjBjsjRkk
BgdmX/F5WnwvPLf8w6v/BYUZOlXgt98BsyL+T9sLFYP/33ZK2yeZtCcUOaXynx3FXuF84dNJCCeY
wjutDh+OnvWbbWEodAaewOpbvgBRbwxZEAOwXFslg1Wa/IK8gkXL3mhWnuQbqu5MrYEbmiMFmtQh
g32W1KoI4jJmsUDdbxwaMTevkiQpoYphEAJMMRtNGeuPBM/ovYsBf7eRJvadCI7F73dDtKUjnkY5
7Xvst2Cc5ZdSY4u/XDZ2iWh4DRDHgettZNlL3m+quQ7+XLSoHyQnrCiCPIAWhDY+Rbdzif9TMtiM
T4OQUWU3YUYRtOlTDWFW+MwWgDq4ruKx+JJF2mdlThWPHI0KvGuS8o4s8JCaoOLCXur95tDs7Tv/
BhmHWIwJoCXBIqGZcqR1YbPQ6zs03HfEGelYw8OiFx6+K5SUN/tQE/smE1sHVWm688s3Q0df5YSU
jn5SdhiF6CpbZAiIH27MjrIdJfuAn9pL3cvwfs5zr8qOBhwqdMvqeUbGNmPN0Lwp51gRYWmMhthn
UE6KU0TWKckkTq6B55WT8iS2LBSVJzdr+6a8oI+VD/WiEVhhnBjevbWn8l6tf0grO87NIDdlpsjt
6iqejgb+8UW2hW9m9x/vJDpjeocv0Xeu14WeCNke/aRkWkdmdB4fg1nq2/YTR2/H/+P34yOVfwkX
S4odPt7Dbcj/5H4FfSHhHnkA4s9mRZZrMShhEsdh5I/BU06kR4HnWgcxf9Pvn2guqOeC8DLxVwFY
VPepkpIMIHap1VgCMLWxvEyuhVY8Z+ldexbrMEz7atRH+upHCxTeBfDDooMBmA2TiCuE33nnLooT
ptt7sFK9EMuhm3aqkwSig8UXHrSJX1x9d/wELWDuMt3tJ0vFXWVEI4DoEd89EwfFaiuVPkkyL1ER
PJspadAi8zOag2ozvwdV+G0RPIKo1MaqxePJd7R2LbAfu0tKz5pOW5YJNjJWtzmMVycBVJdf77xs
Qp3fYe41AhQhMHGgxVAh+RcpgvHCSM4Ebpf/1GU38+s6k0Yo82y6K1Tl0840KMfksmK70zMeWdo1
S642VUkptIIyF1HcPdSmeX85xJuhdqhpi8e9uWlBkCj4wC7KljyPuhwlGrAzfaF8QGHGSUAOJxgz
aqpPTxZo5XfZPemS5aLUBO3R/j/RY/CEx4F670J/nEAMmtHmbGsxpsGNAnMrGRpvjYdsgkLWnJsW
a7KHXo7lawnv/zE24pt+LLEG+JZFCYOfYnVP4wc4Rg6GJzNgd5v9w/9eypEqq7HhSsYsAhkVJPwN
YkgfFWa5QePAM87bY3dvFpfEHeW+JJ3Uf73IdxNd2pLxD1B6CU7UxgFwL6KPkWDuN4zAeu9LTaR2
Nw0l8RALblRHyYH9F/XEBEoHjlLpFavXC9MCtRo504FI9EiC8S2A5ohmjVffxvTMprSlmJd8OD18
EHUJH4et1L6t8RiuonH6QsxpBLIvDQOtw1zzkWQNqH7VSqmSUgmPt0/F6BqcWuug6mRj7qOJW467
tKPDnTwpyP3VsevrzL6zyEjUiFDYihRuVIYlYiN3z/LN316bUaJrAUI2slUz05zHhumlhE66TyPI
6Y9j4+ywN4xxgzBprtB7oKqBdQicb90P4ENhRqPpj2YVgDg5MoMQDHl4KIcSVrrKYcKdsrSAZd0u
8NUPE04rqOwgtW17ST6S7y2uJsPYi/gDf99NYY5PBfnQdhdzOOark7B7pEAX/iLhXmpf5MreVs2t
d0WjEQmHCRKXp0i9ohEDJUkFYR+sXsUmpoLObDglncsIeFd9hUOXgx242D6/OLDZ33ydJ8RA8Pfy
zKVaVpVX9TNA0DRuB2ROQVB9Z8VsCaVcjvDwlvfEIvFfwLnj+xxNosuJFVABsVtGIDwxws7qZNmt
ymYj6ovZ3reRhpWig47wixDiaYHYlvvZlDhWH07BiZfhHfRz+OSbymikHL2CeD71A2fe4ICF5Fe7
G+NvReOySbJtb0vBpo4NoRZNdTrC5VDyxgjuPGvhOY4rvi4vUzcA8omGuuuQDFc2JFre4QDYMywZ
F7LI250ODQ7+sw1DTSlTcg+raeT2+q+770UwKOgszmh7/bNj16mrOALlvQZsCV9AiWZlnVz2wm9o
olbK/4kKKmVwZgJgDN7qyo8HKmmVtFOvSxFcyyfwJ5ieenddGOOMOjpgHVp9d9lLdXr43MCxwnUS
O+91VWnJt16azqxeINeSa6FXeJi3t5+onTlzyqhKVEFazAfLQl+OJBWHCWRGXPjByTrK1H2fGn7Z
vDPAKJjOOytQz2psIC+3mLLKHKwR6AEut4gklwRgZSnVp/YXXzlnBCOdmesLV7g/q6FHi2OXbaKF
qqgFGGVBumdHAC4r9vlW1J+lb/CGZSwGDwTSPNmfKw9b+dqokG9YuemkKZg9pVD1+yY2m4+jADTB
BEGuTIOS/mdTzeM67Bxq16VW8v5lyx2H9vHTfaC4C9h6QnT5fa8SoUN7oKxvf5Cm7KqrFpruU9EL
OHE0evGT7dcHhtuH8kqbhQvQ7NcV7FBcD7OvUR6A3EOKxdKA5uV7HxhGHKgcyH9NP6tmBGxZih+S
RE59ELJ1ac6uOAAd7ilsOLnXpcncZFDzIKJ+VOEQtA/5SaHref404sRtISV9fMG18OWpVwvJEn6H
9Qpb9PNwbhSW1WYn9zfWyL6RiKIr0ooTAo6T17v99+DQLJC60o41FE6hTb/2fpKjQUV2QkK0oCQ6
hEodHWTSLzlyA/jkrNCV4E0wrPs6sBpdk+8IML+LmaQAdcdVUCnPsW4MIcymvKELY4JEN2vj19Q8
6yJezKdLpYOJLtqtqExjZPs91W2OHB61/S+OMPMe+Zr50Wd4qPQR9HfvttluWFLXYQCwTGmcpE+d
5VRtHE45sh4oH18OeU17C5TGY5TURFKKrWhmqKvxBX2tJgklB9YdwGzJPwmtm0/sPBpBj/uGYRoD
I5KIrRBZh6uof61/OmhC9pU/StDqNWNQnVxT4KVA03Ec0YTy6PBD3oxbVio0dT4QhhznYcI6r3LQ
Rgzf2j8XGCmDWSoaqtQSqFFieaPXEn8Q5zzlj3LC/qE3E5VlRh6WX1ZTIkPwlVz3KVH9EwfMF6tq
W1XH7PJ2frBsh6sASdaoZdLzTX1VtiRhhATzIraLh3LkoZRN7OzjIidm0R/wdw1bYssMyJ0fswrV
3AAtUU/slDnmMWufFjmQHHVfE/iWG1zxPzX4vfBVtz1h6Ny04f2qFqQbBN3ar8AxbWOCBL85aYaf
kTLOph7i3yWY1S5oumKEklbebQsrMv1ykRrJZH6of0X8Kw0ngBHJDLISK5hjrXcPv0tkbWCZsCAD
IzydbsrmcjiWEmwoNDJL4xqGY1jVMBufbQt4v+XNkNIhEg41flDQEOvZMLGbYcfcLMPvMyIofJJc
Iea1ny/M/DM09jQZ33GWIt/eOt1aJhqZaG0h7ABc06g7DsnwTKfIQaI5d1dQrCHFRANxZy42qekr
PoXc5JQDAHj/Fb1BSpDZP1oYWGig+XkK1mB5+OoGJ1Mm2Dx+D1F4cmSSQQXWdwsAPDXEDRkH3sK4
1loMrGhql0WDMvt2YAFcPS6YdhWPmD/ZyXp871WDPpFBP59U4sD3oLm0QIE+p+0qmz6BSOrBR0Gr
H3Aur0b8UKbNud3dkJxkThqlJ7jBbOX5bY4VvcRzFOg8wphRF/1VR5PisMcQGlz18IOzi7o1s3wt
l7ZCeUBkWsvUG4a48+vIX//kTl7pEAHVXRU0BuvNC/sVS93v+kBzO0pjCBFUlNEoWoFlP2qdmQLD
a9GOUk9R1tNdqIPyBQgGq9WNb8KpO66LE4xTQZB0JkE9Lol0PmNu8MLjzkp4x+4sXub11tHQfVB/
sw5nzlpav+2a2AMDTpzkv7DCiCimtw4EKA+83+j24e0pyEw9H4nUHhMFVTdzTui/ABpJYq1wcraU
UqLYf3b/qgUGt+2hlEN9ZDH0rQvm6R2UCoMdwtHOZ3BkfgN5GQipgzBYnq+bBWWRxN5OFRWYPQKG
2MstVjIXkeIF5+m4Em58spLiTe1RfCuSE5OyjbQb69+/nuDZr/zJrRenh2xMwykUkZ3QmzXFPT1Y
qTfDWuB6QYYsnP0b5JiOUzMI+ZsP1fvz+/3S8LotRhC3CSu8uzCswKKeD+id5DZRiuLGMK9+fDcK
1gRIharEE/4j9NJex49D2nG/d6sxWk0ZMKngjJwZ5X8Fu6660ffCZ+TqOJXVfrsbo9+0TOKElnWk
co3baWXpgkM0i4xBiiA2TDA5I9pqCfP/KoRkTKQ/4mPl4oYk9+nmycHxzrsDSqvRWKVw4PTlEC5Q
4nCPYpNXwz60CAz3Ni4Ig/2dsl3hGzd+5CEUS2LohDLvcJAfuYvernUaWgx5KiVQMz2LfhwA5FkG
9c7OQR/Ejzmdx+ue9T7HcNsnEpRKUbW0atz3psF8t2SyxOOABgu9+sreIb4U2oKPZB3HHYiGiwRb
A/Ep1ocyqXms0NPtf3TIMwsGrqyc5YD+gCdrgNElQ53KwZ2eiqTDKk+XzSK6yJOCjzzmbfRN8FxX
tiIwknh528N/stZlIVPvK9SnWDBsS3Q+ghJetaiC5qpP2jKvKBV5nYrycaZh07wMr55TeT3IXg/N
hPz2hHN0lHE2USCj8jEGLfopX54D6aGjtQ/YICHGhu2wjtfM2pkxpJCeL+ZjycRb6iVjQh4izbAj
fZbDlLnETFiMzw1Mb8H9ujb3pV4WO8w1Zyoroac8P74uu4tyvwbHkQ9ZeN8wbGB4feQCKcCdjAKA
TlQlkHZgksB2iAdEXfzRVxDJI37GMQcj3B6SdglpIEKIe5TW9877DYDB55yLJbC7vsBsqWKjMDA8
fsvIr2PfedRXCeyK8QXzkQ/1g4/ciD1AU+6DAHESKWbkRgXLCbTLnCTqKsZcwwXEUY2pqHvJ6Dx+
EFY835xJIMrX78pzPvRxFF4rgyJo3lkiMVlnnRC0WbeeuZkiMZ3W/ph0D3HhTIOinq1PV8/AqAS8
6gRm0l5+zv5KjzcLSaigdhEFH5QB+PmDSlgGsGa+YlBIDMaZbV6L6iFmIbD/aLOREY5t9J0+e/Dr
v3P4B6REmQNqGBYbRuBzPrXgKcLpckRIwQeDQ6aXj6+f+kNLKVLDdBi7NpSAAL81M1GP99UaSy7I
SK8GXdGpJmX+s+r51fA0tbQXdY0dMcG9zhTni3WeWMNbc+oSCf+Vr6iJEZGGdHi3HHybHI9Fb5ol
Y2JrpeuAV4Xc9MH7Ows9zIoLvCEvcmwaYy25hTYvxwc2+soHlptBtJhPNnpZHRbhARtitWTuEFTB
dG4SxcLBGYLs48PrZboYQWopIfrhSH25Nx1DtTvASiHIWsb53VJuYvZW3IXBFrdMt1bMaz/CmEUD
+toLZ16XF0TpSgSrCwOYO99JKlqU5gz64+Y37cb8buIyjdIx88RW+RxRNQgEL/j3xID9faGKRgXl
U8js53RPS+gWhi3sFQrkuR8ZUek5P0781Bvr67yfIMHK9wnppu7EHHmiGmtpC5WmTLLIXMW3w8ch
CbgZXSL4mLuD2Imm2K3dDofPf0cJftR722M2bHSkl3Kix5zwzTOLgj87J3CctTf9ZYqEY0W5Any5
rXj5qm0UNNG8n8i6uhXeSkaw7YUm8MedQzfKlAggloo0LQkIGFgMh/l2vSZQOHINRSU6GZffks9v
sqAGroV56fd3yIoJDoKu6fUVbP92jrcLTyGmgvOFTLO36c2if406P8eIKJbuIfE7Jgq93piBXSHS
9cS293iPShL3Ad4VRKVgbewF10JRa2wtPZiLOASFiKBx9G8Jn/NOqSmfOV3IJe8ZVFNEAsGvtlHG
VP5A3AqmIeBBBMljSTs6d0ui3voqvDF3euKilEt+Ouy80lD5UjQnZpL3S0OWVtvXY3byMhLRv1Fg
CDlzjZXhkEY5fq+IHm49DUPyEheD3A6E6kXEehNSJ8YNg3wALK/6lyFrdTJau9aflzUoAMscH3Tx
nPfAwR2nbmZefOZrJsAdneeGm1jL+4Byz5JFUPSYHL86yszAdn50YY4VbxsdopUXLv5FAWLvXHUd
WAgCyXfsWzliDftAcMtdv1iUTlTgWJgfubZQMuDPKG62v66twGhV8uVzM1q4nNzrWpIhWruMgC8x
a7Ei4DDti06YT4ZAuD8n3tqAWkUfnogP9Nh9ckYLlndjuryAyau96N7Z47KKdEYKZheIF5z9G8mh
6V8VMMMk2y7BwYDEahPJoFDAL9OnNSLcVAe6hNe8tJqmiB1mwfrS1q7WCiGDpkDNxxm3SdsqnnK8
HOyQ3o/uh3g4YHakofS6RSQAUDFAVF31NyXT2zM53HpPmhmdp7bUme87hf41M0TYbSV+Q8kS08sJ
3VRbT8rblCEN3AIEdbOlDH0cjwCL6wIpKykm9ZCg0hRCKDVzkVyYSOOzA9iG4GOoyBpJg3kBwXQ3
oxD0tUGicREv6uhbKlJmPjpdUSktNCMc2CmQbIlAunfdPTRzUWGceIJ0ZaHuOIhXy37XOZfCkJqr
xHhvitvbN6QTMqxVPBrVCbfjJw5aPZNPufKFqLIUKRkoCI+y+7oEYwmaNwIB7f4O4540zQ361GAM
8yEOcJRnp21YaeL+RLutYr2/0eUMs+dvkGKEVE+SoPJhADTq4JE+7HSPcY+VL08zXvTZNVpdwrGp
j/AVtGiy4koBExRAFJa4XpPIGLQVc/g334lNlZlu3U2WvI2Cvk9gouT54CJ581RDbPcW8H5mn+Qz
RKFWcD7t8skzp2u7V+EEcNBtvK6BQ/ObwEZFBCdodkzYBHYOJ6ki6hDGRjudlFDP9CZUO5fchpby
1u+AIw5lBS0D67HoDKWTrM4hG2LPEo+i72wedjBwvAYLA38s2ApHb60U97rZ5TdbuJTPL2cuDWdx
xeklfGiRVGqKx68oG09BP74LrxJiOBQxzpq/YZvitT1zuZFgeX+YAzhjSsBLw89SA+85QOTJPJYo
0Q8+tFnC0O5VuShWU1448KlNz6jeu1MQU6BDJMIGdKDUKO6JvBOnqDLLts94itDQx/PtcqneQaRb
CcnuKt7x60GOtLSXhrSwPcUf8SbBBr1fAo9k/KZBrmaKNriDw/5FcJFWMy6pYVHvqb681XJzgz4h
iazgrvCJb6EbZOLsTTaq+lBsV/RWqdZkJqzY6puOW/0uieG4WAoeyjhRpNddQ/z5FuZNPztMS2CP
vW3O2N0a0SZyAFHhm3JyIxSyAntEF8jCcH63tm7B6p+6FeQYB75e0Zy02Xl30DeMdYUUuOxeh6CV
2wPfjTPlRK74ADrks14F7YNsadWcC7rClkKN8RocrKzid3pO1Hl+qteRa1/o7ukb4LX9iuTNLUO7
vZ95vDXsiOdGmAeYkrqiuTLjRobzDe9xJIbmsgp7QXdeFExNARK98JoFwn2SWdAJyV0Hk8rbr+fN
+y8B8uGfpGoDWSDyNmv3t9ZxDhJR8wQ/0dMBzOg2UjcvWKXsrWsVkz/bgqpEpqoQDLtUXxvsWABo
aHKfYeAJSV6hpuMI9W+CV9W2zHk7NniZy9fIAJIvyTy8YksOCH3xV9WWTbjxP2CcDnUPtUPFuP8P
ighrEhmBaswbINdD1CKkRusIvL+UNV5rgcUlYoJr/yrdYdrNp9kGMSlaVQggxBXIz26Y88Jb1mrs
o5cbxYokQB66S46bEUx06UKfu+ezUootwDuY+vb17wVTBKM+c2DvKboYtFNUCFWKwlZeQoC85SSQ
WUgazqJ+0nXs4BalU5/Fsb/TRqd4NFg1DeHYqsz3NtpZsnGbScVl4b9NXBL6Ur6bB9riFqTyafd+
qIqsa8U3YETiprx1b6JiA9Bs6aO+ZEMHM4okCqK11740Y5FAY+WJs4o8VyJTfMGczHHRa2GTcxjL
K3qrvtO6T6nXqxgXx2BOz7HQUWUqNGVGhDfZdHw6KDNc/nAGrNW+nFNNDZVZ7BsOwm/UvnUGrOUJ
ClAHZayOBRvqFMqxsQQL89rFtOTxiTmuMvph+nydqJg4cgoJfDHVgjd2e/geklhhekBJwKSKawp2
uhNoKttbeBI0DKePYzUTGIWHCrdSAi4e3knH84qI+VGgEQ4n/jRKGG8ItWt9MnOAt4CrCJ3y/OV+
7xPqDGrpMtbZAswcviubzv5AFxwwNl0A8BSPcMHQDGoyRbtOFbMChvfRRkkmUOuXQsoUq/CGIgmR
4uySPAnHZWYdZ3lSDUDk94LhPZAoHWj687+7P+aq8IGTtfOtBY9Mr1eHczOP9eofzHoMuRX0mM/3
zslTcOd0Xj9sATKO8MTOu9SzcQvdC73YsrVNdp7yLaa1mj/jIFMBzBhfwAgiz7E9KmB5eCJUiPuS
5Zc9smJtv9UfwibeMNJ0rBdSbiJjiQ6FQMqL2XgA9wea97MoahPQ8bdRGKHQCuxP9CgK7dvurC9g
8AtfG9SLjN+PVWXPwz2T2NbXaIuHuWfHkYNIqPZuZ0ZeCOjD6Hn8HP6homY+qQ/R6luDEPNlEIKh
2rZP7Ijj2SoorQXJvkOAjvrfW/X14owlwjndQZWSSnJ8z38vYwQNUANfxWHnz3b3fBRB8hFgl8aj
xHCSLrDxKflh3xYgK6YnFtTvdxriGSu63nOWAl8t4PXSfcRbhe7j3MJVagHwjbhzvg/+yHGVeB3q
ALmERXuhkk1OjTWUjh/BiMXCIb8fQoJrMvjUTDHVvYCZBcVxAVXWrqYlqfIh36xIqVPCf6sVnPSR
AJnoOJ9GL+3+bVy8pnHOocgusRi+Yx0lKr77az07q4y+9B448+Oa9E/x1TpfxYrR+nOpGabFC43d
0i0fJkjTXLwQ9HLzmqsdqLFWBxCyVlkiLFns2BQWlCSaFmjmOzOkcw5xYChZo6bJpwOsN5JLG++w
rtTRCbJR98ta6BwAfNXH9YOdp8QucbBuFVZNtZ0XaQSycB5SCNjn69a6rl384juTJ9p+4hsKv3uR
zeIFCYcgkeS2Rfkn0KJGvdt3UfKv1+zV+w/kKfp59Zdko3W3LN0NPC18uP+Xk8LAbgn1n8uY1L9q
Jo0j5sBv3ODhIi9o742Pavr6LiS7Zn+wDG+HrIQ4/mmCcoUASK5UQPm/Y3dlCRikf/xeHTVqeDww
xOdP54k4WWh5DJpIG5HwaTlCpgUuCfp01YvGPca+IKtm9F70AKDCINwOaxX7O4/G4VY7sw8nleeY
wRXwfihsWsyQ1J8AN1JWTZQTH5iBKHPk70UUbBJFo7zfeqsM0cQVIIdj+a39gCwQ7ItEtMHTjiLT
W/8H2Pe4vBc8ea68l5Lxsaz4tCVQh331UH+1YcmCW2uIfY8aGqkRGnwJ3n8pa/Hongk/8Ce2P5bl
Lm/g5rGMQrWat7vTcyGEp8WeRRG5y0F7pUA/iNuiyI6wZJvC1yms04rKVscdtSO7Ud9eyMwKNphM
dAdHeSOGEsrvufN9PWFrdlhSu+Ao5cm9xia79EUFyyOUbXIy9Dd0IpUrnVkr1JDKina48fKuiHMO
eEBCf3YWQgk51y6X37Eh4KB1IsEfQH5NFuEZLE31QlExexRXp0y6Zvvl26Nt1CulDzV5ZD3l0cfe
3IgamjDPLH9mfZN9WPTi8/AwK9k6uP9JK/Kq3Ze4BzESjzl/Ufyh3YDFlBa/Dt2X6kiY2ID7OB1N
pHdFdXLbI9x64DszLBCqignBLzVvTC3lR0vf5P6o+N/wNlcU9+JlenSXboeqA+FPRTocknOIblGR
91+0wmtMF8I5EgLEC8uSDP92HmwEuXEYMEfA8SBHNvBo5KQWKSjZhvxuG/w+LuEEapKXYhfSmUNE
nYjauwkl3C0JlRFPvz6qd72VSLpSCtZxQVAl6ICQXD/WTSFbl/MAt9Zi2ssDOGsgWJP5BF9zV7rh
A4cSituIC3bFQFPp6ORCn5/c4pp0/S6ykSi0M+6xoX/yHaJ6M4JNMXoE6E8f6U+lrpjuyQpoUWEp
53UPj24eOprb+KbLq6rwDZnfrh2jPDuefbPx1lVyVe9jyj37LYAFnp0MB3/ptToMEb3JgHKFWZYI
Vo6Kims1aGgHOP42SfOOHYTBGXy971xRfoYFw0/njJ4b+lHbXbaY4rZt0xV4LgSvsASOG0yWLGZv
SnLXrL2SojPy1WNt2lqb0i4v+vaN7tUO+IlQJ8aTvwD/TpQBgMCdkO0zcRkwTa5xSmZVI8qGcy/r
3S8aU8Kg5pc8rLTr7xX/91R1EuOXMqZGzZwcCf3KS91hrhksr6tSl8w5KpA88s3B6t4FdGNnyQuH
5vEMJXuu8GeV3aWwXk+UwafLB5uD02SMec5EJgYyyUWEX9C+2x5gFTOyLBvmpw61YFnweRdZk6LG
XNv7Xrr5ps9IRK6QRNfB4x7HwHgzh/2p8wDVsbxlYOf+RipBGNbOUEpvPrLo8EsNm2gYMP/9Ruf+
gz1voMSxyRy9qyTSmUx6NKZJQeBv1ZfeiW8rtl3JlUfwhR7SQWdVa+nc4thyMTcCXl0a5p2jnJ9l
/zhQ9OObmpzmLjKqEYA/buiheoOXHPRTatyuxy/VW8obuEcxj11A6Jciad/imDA6aqWLqwIOxbbS
ztqiGZpu3uSm9G4UapbFV0wo32pzwh7fnh/ZpmUj1doE/bzRFporLSbETx9f/aQDCbidCGZT5ZNP
SceNz9Kf9sY2gPXnsmJRXW60yd2lr2QsQO/G9ZtGg0Y44RY7SI+J4e24XllCW96/sKiXYNe1LsUf
8Pv/QOEAtZC9+DYNSPxhpqo5IyImg7jOCS5zOKxcYrkWLal+O2C2tI3NLkkV7hUsRqfREa4un6XY
n4MNyrdYSgmx5uLi8Bv2GLNoVgTiURQ4k+af34phHA7eXc1yn/pUjAGwfCJR5D3CvJfe7JfGfChY
vzboMd/Bxjd/6+fpO3T6nzLlip+q9p9Ale8+ZcFM/p6B2KojpV4W8fu67JtUIH9dO9UW2pMNTcEK
e8jixcuoJofUAUEcVcdz6mWIvZ8LmZ8qTPG+Nzvi/v9f5xEngog+z7/87gBRgBMwMY7jQAt+Zgtl
RTrAJ5xw7kBQmu41VUFxcapn1v8C9hhd6dGvE63IHvTkoXgkQAHeio9E7O2VjdUzCeywVbMLtJlV
XmO4AKkmEhTVDDaACx6pw83sh5PeGCY9ynUVWH3pnU8Ny2cCioeV+2qsJrQhrMwnl/Ivpcv7kasn
a4YEOWKGQmLpb+c5+j1cYPbM/rIbF6J0unoDKPEtzb6SdJi/HVvBCbQ2mSKirK1J5nlknXCbZuwA
2JH9Hv66YMTGf1agzW70GJZh7kPc0mokDpyzLejWTMKFhUmZOw+t9NvEyFPugrrwDhppLghyqsPo
pVYdfMmQtddeLMcuQQBHQfA7XXZjch8MWGAnGvMZ0A6n+tFzKkapAxTwrQHM7angBuPkzBti1dGL
+vYciOu8c+ltw1LGz2BK6Ahm243CtPTdYduMPdqJIB0dPbV1SYU7RtdzlxaJDwfdSjPBxq+mvMzD
o76bEbEA0v9vHklfhV3nyQDiXotGlrJ8umcOwt5EM/5Utagw5jKY0wzXGG8CIJAB34GaDsOrhuGo
tSQ/JTpQTTb4ecfAHducv45LI+LQ2TzbBWL1UmudDRSFuemeCByOtSE+SjdOM65JzaxqzQ20UH6L
dU6MeGE5c5gFZ0yUnS44CWvBo3+bQpPB9YdH0NwucuYebBrQkXXU5OjcayCQTzExU8SswwBc216+
lWXjgrQ1bfAIOtfnVhko9gqsRcp2YSVSszLcAvzSOlyK8hYJWkC834KWCoOdA1tvG2iML7eUKbHU
Uz0hGxcaRawHOjamt2PEvqKWvuGNhNOFPNymQwUt9l5MvAQc/VegHUIyRYalVEXo2++Y4VLSt1qD
zTRnFGqsSqAsWx1cLg8+kuzdi7pthKFHheQTj5NRCCeVztAFHf4b4Q/E5EAdK/gSjKfTiaRUoDKH
pUTrfgeUcfoiNLxH1kvpGSFsvHUa6SxpAFIwiNObvwtfoUdmPYOEZML4IyJLxP+Srp+++wgyWnIa
G8hIrlTEMRJ+QcMX7dNsQ9cCgzBH4/cZNLO4Ei5IW1262TGkGSf+tn26+sQ8wDPtNdKXsQVL7mMU
xg9DcoxI77vKtg5eEc1Hw2zmR25uiOgkmyk3J2koddvt66cyAIWO1z38BRzW/gtOk4+GKn5nbFTd
LU5sTKH1g9ah4Y4scWhZFOhCQOhXGSfuCTw0mXfupsv1/YhqoBOd5EiV3QY3QCRpSkvWPE/pk2j5
/PSo2oueMVDFj0ovVqwxutC9cETT6bBUbvEaW6aHmo+QVDDr1kFtH6iKiIWcFxBz7Pd77hJL577u
go197RPrMpDmrWHJ/V5qmjJLgGpWGe93xRbgK8CxG+f2ta4VQONI/DzyQ994z487ZIQvj9rNZC6w
lxf8H2CWvgOy+1bmT8LP52zTuqdjnBxog2RDQ5DNJ8u3fvffh8ICHZGNBzVA5b7cmlzRVSyl9bxL
Sutzr43rOJE6JNIOGiYdZI1IHHB5Lzd8wFkriScdUo1NN6xeqSqxc1Fu6T9upVejYV7T/zyUyJH9
a0e9kDUP+GEXWFWsPSpi+uF9WlfTSBM0WNtYen76ImWPhaYpd4JW0pFYOq3upkeHCXWd16DtbS0w
hkCZ/gUFc/Zoyin/dOizEpkPH4kwHdnPICV/Ch2jAhSPfuuP4+3oXqJ5pC48eJ4iWDkQxFK42Sbb
afuXHkemY7Jh0OyOc2bHTUpqrwHv/ANhZu4V6zgXQDyj9lpsew0EN6uhtbwDvsEGBAdRgdcKSIyj
EvpWnI1zUHB9b9wa9E7cLokXxIJxrOOqDhUV49hrgHpIG1eVL57e3DO+32X6dvuzqp4tgsG1fBMC
5D3w6PsESD8VlEvt+cgBeQVvuqblkWYmiNWIUhl2JX+u8ue+53ET2GS2JJ7vEWzcBuI5ItItsxoZ
u9NvbFXLg2405SkeQpiD3wrUYN1S/2A1bdvU5U5fja0kUZrbtVPEdD92yjyGcya3MxRX8pytIemw
RYP7xt9FdbpbQuEMjKfSzhqM+7EDtmGj1G5WLJ2zi9FC81WCJ4wNzM0Iwamq3g7KGGFkK7ozdy+F
ecnq8YU8tcxgbBpj/gVGLppc3Sd7fGMSmNN1o3a0vVfXcl6eTrCHNYUw91qV6YSDRRdKbH3nr2JE
b9f/htpbTQ/lRFsWGSuOgDyEWvvUwlrcqRPofpvJoXN9C8LSYHpQlvasRrkELxcurHr8tQohJ19U
6ZiWfsmGLDgUp57/aOMNPuNOwuPR4UP+jQcJJx/+1CO+eZSYI1KfPunmGrKpAsnI78lWoMrVqtzI
OqDu906TvMU6SopUfDas2OJW9lLL/EpHxJJDVxFDAts5IU6Ktuyo/++1BdxXZu0OrpMfPdnFx847
uL4xo6YBoOF6A60sW63pJ0K16vg82BEMWHa9UghIxNqOpKWwx+q8LaTd9AzQ1isEB0iWcytFD9pv
vsVR8kdbUsyZJxKBsfrJrw9Ls5YzjPes9rCHYySTR2V+6iTsGGZAnRxOzhqio8zqYsDfrk10q4F0
wOCtxubkKGUVt/onqyo/UPekqEHBIkK47tKNS2w/Xda5bBrCMf+0naNmjQR2iKQcZLo3eckjvvAW
jDfZPnrTrNh5pcIMAxiq7bPVnq5Q3gleKN+UX+zRgF3XuhFcSfWNOG/UrSoAsdaYVF61b95krFQR
vHujfKU5yVDavmckNAGTqoxtARr4dBWhu8L+dbM0G4qiAEucvfGN2iMQ88l/A75EC3XJGckxEQdK
0PVldDUYYejL/ibsdTjEQohTDN+ikh2TQtM7SpxrIiOEHnX9Ry9HVFAYnyFutw3ywKHtFppyCGey
LzBHSxR3VWpL4TL7qKrzziiIkp8cU92ZsaiL3UfNqdH6F44+NitjuYfac5aKFw18+mO/UvqUbdbl
Ou+Uu94I7LurTpvyIY2V/+QN0IIpgpptd39JTo5uIe3p9jvb6XLYNVCGXwyNtilfRl7GukMMWeWd
aqrLIyQjDrTGj92jMDAjxOFWL3Io5OC/j3/B8NQdQfRVaGM9sYM8NQZj4Fz+bf33J/1hBKJsUVYW
5ajEV04+7FlhpE+nGVhy0Mk1329rgKx5TmrF5PbaMmx6jhwRp1plqQFU4j6rQsZ2Xs0yluf3zp7G
nSOjezoFGH/z8m8PnVKEkhayiRDNDgwkjQSmwS+yWf3IMQhnI/0K4QcLWwI6hRlh0+qo3GkyGRwR
+Tq1flQDjv7E98/3N4IS4P6DMy1L0ukyGU/bRkM3RAgAO9JDa6G9NcK3RI8QnZatGXj9zeYv5JwT
/hljH/PF6+lbjTSqWi9CzKwk1wvJ+rixj6MCgCgpdpnMAs6Kj3LtKfv2h4qIZCJ+hRUDXpAWfRVJ
Jentqeat/pgg5dbgOiUV4S7rebRPLacL2CYTkWlUF8NNktgdJOBE++yi6opiZaZL8jZrvp3FqKid
7chZmTGBvuH5/XDgCrUJip4/wVW008OZnVZJGtvTwG18CyhxLgrV4HiIUe2n2APb/R1uGZGi/8Bq
MT1UXwYqe//kTaexuRHWrhCR1y+GrN8QxtO3d/q76J7rt0irqvrBT1s8uJdloQNyXAVMngyg72WQ
buuci/vw86EmvRyGS2BYWXN7oyWIO5aQiVB/O3BfinaeCtn+SnsVeemzydNsEnJfyhqV5mxBWVx7
HxiwnSsDC//TiB4mH49rsihb6R/qjMq3ZZnc02UYQKiCZww2hwHwjia30RzPMkfzy8xamKCHkQWA
RU/sPRQuwWdfrX9cP3J6Yep1Mb5C2mjpuJDr2ELanA3e/nJ4mFBD64WC3x4dMkvHSnl/yoyRgJpo
2CR9L0thNTrit7i/zgA66tYavBVp8znq0ciPCOIPdqGbBzf85nXzrO5yN0BiJswRx8nG3h4/jX5g
1jXzdkR03MO5HfAD01cPn2awcrkiWn5jaNeFxzfzfEUFa+pu5P1xdjaeaNK0V27GmybW3YNGrH5p
Z9sq6mcoS/+wHfbrRIk2xkC0l6vkR3ugSFAtaqegWLL0KmToF2P4hLl/6m2zvtZNscntWZlg+0WD
RVOaGUvzKWiQ3lb4+cjEhDwCzASoWxnqCc+u6yy580w+Hilj25uS8iN5oYBREI28twFsJM1bHaYt
wCaovkbhUnaGoHJ4UZcHVhXFztYNJ0iPrgZ388P8TyEiO0eGnHnVFNM4Q8PUBoqfYnNIlWF4tk55
LUms5QcFB5TXjh7uZZAh0sgBJTEVujAzC8yC4m4T6Pb2lTVpkF7rfnsq/4DShwtA4985zZphpa97
ZWWdfcau3KIC1yKIuRZAQa2Jfs66oYHywMN8B8TguV3Dxc6IRqeVqW8w1n+m1hYk1nyx/z3iliGa
hp+D3ZGe4Xt15a5zUYoL3JaFTcI1OWSltj0a/I7f45hHVF1qe3ok9bN1aiaT27bZxK9s9X0thvmk
FLXLx3UKu/oL9H4SmhTTIny3s7OCPpXqFKIsnOn6exA46qOuSKmcnv4qBWze1IoXXP//bG94PT3+
Xw0sEQRzsmweaFbVHd3k4pUlSg1yRnAHoWsdrrGK8v8tM4Y+41xxS9WoWU88eHrVQ9tI4aa7FUwu
93y+6v68HRvxfblpmqoKTuGvxbTY/4d5U0hUjllb4BIeEZT5VKiRESZ3yai7lKiV/UJM7Re9AjaE
cy7XhfVfULQs/MjwrdXX/measfEQGt5jvr0d4enrhXH9im+Y89KqOP5IkgMw1/ihpGtbleUiFkvt
bcsO98OkLY0VmuuEY9ect5ssk8rWe/c6KbzDNpAGwpw20FzNaeQSVs2FhKY3OpC5FqUuQiD6yIqO
4SUIN7SwqPALsAFpgBWk/qC5JKfCW9gmrizdqqBwSbyLhU7LM1JPAMowYYzGexG3P5DalUlj8KwA
Myg5ObI/CGIFqtZsHTd0DPimdcDkSjI864eAVuVZg3+MlPaKtLwv6vNL1SvFu9MvJ2hxPsO7ckYx
J1S/n9BDwEbUzkmN455BWF82AgybefJiIcWu+cWzUqS0Jbzvw7wuOApGWG6GjebILHcS15mhGgTk
KrgfFBYKizC7O+NUMmEZOuFKo7TIXMVRFdQkZHzWyPXMzK1r2WleEr5poCFuvG9VE/VeMsu5PSQZ
+iuq9KOXsohA9KRKqE9XjYE4eMOjEwmbgURQMFBTKdo5px0G+/ElbXf3aylK8t90iN/eVaKwzJez
qdleJsVMjKEw2HbGoKw6IWozm6WErrSG62H5FxN/yuEOyghPl71nTE2EyXGqr1qO5YS2Q4zFdqVB
LrCdCnzxzwC9yYpP0x2PXbNK1uHZJbBLwG1lVubEnX22Up25E+OuBdeW8TLIz9FQOFCJN4LLHFJ9
r/W/psWdF65PshJGDGC8CtdkWs4nKeTYntdZhA8cMKuZy4nUwLd7JSE7jRRHwK4Aez2TfojHdIPQ
NAU0IsnnWg3cP9tn8bxtUdX+RTbTwpeRyxHIKvqOiAZF8solmdbHfpBo/nRVW44Eub9lbt/WGMiF
cY2a8pqgkDbJO4N3duhdBnETK4YA9p+24POVcN2EiA5E5UDN8XkzyWLnERp7+6XxyrEfxd97y6Dw
Uky4Cx716FoBe3YzNA3TYgUNHIKnxq+bWV8mbq1RnN4u7NUwAZURx7sIq8Y8Emd/FudW7FREzFWp
pvVsmJVZslVy7tWAz78OO0wtqIIwd09ojvbaeGv4p0srazvyk0oS36WpHvZsXNi6v1sHboYkw6x9
hWnTsOrj1tirbGZAdTDP6sx5sEiyHE1g+DwxTCAc0SKtPw4gVkpWCFoR+jxFhU3AjbTaRkZN/AHV
hR2ZbZZsYeCSXft9WS+GEraXmRwTidk/J9vZrtnYTzTYY3v+kSg5+PWf2IJNpCcTNQRn0/GF34MM
EDcuZPwr9p+Hke0wK0zlGvX7TkousjPjKUTP9BSzV/BOi0qiAWz0JIjz/1WJ85sFz++Miee2IAQ4
GQtMfXvEMqI+3JN98/MmX+U6/CNCiVKk672ICPfGiJr9UanPW9tTN5ZczFd66juCFXdKl025wyXo
GepHYNsfwZm7OEMD9jZOR5E/wpmw7joblpkryJ1AKDfKccS/XRdCIErBfu9jv4aaEPFhKH6WBzhz
kRWGE+JkPU+g2k0+eQKqSuRnnvCqQzwDGHMH8wWqitKxOsmapEfebAGBFA4ykUtz+0HYQTiu3zv8
buU9w2194I17FY7ko0BVRoE8vc9F0eRBYeV5VQr78fba+0zhU9lJJ57v497OrAXClTjKq8glh0RL
0aBsz0u8AYQF0EdHsupoctIiD/eNxiag5HwX4B4MH99raKLN1s2aAuqn+clYBS1XBkJ4HuCCtgQs
UgGkvKCzKS2ZiJTqlXf4szWwATyZgB9m80DAzAENszd/Lv1unSqv0zTTJzsww5jNQsAzdPFwbiW3
vUGt0QlDqDphgSs3e+6slx43RTKHPkUOLK+3SsEqatoNVhCkVyfUDY/LJm89K+FS/AMLSJ9SZ7XQ
cV+2goYHm74CNAfQvYfREimaU04MxwxecZqbmf2VuxWB5Iz8HXMYVvNPZhSg3c902NaTXhu8i/rl
SkC0tdZTq+1GUzHXgh1PL9X+MXOw6JI50pW3wkXqByZpxOcAyn4Q3epKKZnWcZsz+QBdKb8Xu3lS
55fZa6TLsRYJ37Z2+Lt1GYFRGPqeJVdkCI/XgdjKLIUZjj8Vk0ezVsjHqhFaMJcO2Dh4SCkFqOHI
WwrJYhQxGl5gY0BIgcPtzNrIQEGCjs5SyTK1f6mwW3mpFuwJL2QeS/KzBjqWaDR7gVMxT/Tj3Uj3
4CV522rYmwro990esjDyADBylm3CYfDcHNbI0qnwF56gfqhZL7UFH3g2yditbA0bRjB3DzIQU6X7
OntN949wCW+tTqljkpMJU1KzpCRh6aAjt8zwWk3Qrd8qKVJZukW8nMXLZhDHRqi9OpVj9AktPyJp
6knaGSYUg9NqBxbBbqkPiw5JKesBpGM2JfzFvFQ8PqD5yy6E1v3EbCWGF55kV9n0JLg4GKTzuMIu
GQe0Gjvg6CUKguMZezkd9dq8jTZ1ftpyEgriDleyeokI350UbG9DAPX1QPWVM6vumW7Z1d7dEV/D
tpMqFV+mq2hYI6xJVvFYdIakUasfOY8KUDFejudn+cIf7wckrEuJZ1rkBDgZaiYekeTWPxKOTMOD
XT9Yac42s4JyJZDFmeg3dXtYamb2iCAbPKAJ1LAVYLOEmEIfWaNI5EjN49nK2bwev03EXYo0VFL/
yI8gc5IWOxwfipHacqscK45hyKpqsR/ymIzY6I7JaVnwpAVpKNYDiPSz31XpdXp70KA6krv6H1aM
cQUyV3YHVSHo8Il3D3am1MHHp/hJTWaceXcUvsDeyVVLiD75eFPzflnj3haop2hqYAxu8oDQdTwz
N+f69fyP5t8/MRUwp8MBYGXkw2UXBNUsELmeDlTFGIUItjbikiZif+cBELulx+YVZb0BnRU9Schf
EFN7AdMyW8G54YL3yhqhTJa0+nzuRAZOitWtOcQ3NwWQfKcD0tkZ3dIJk9zs4O27XFSU6wPaHXXm
GW7YEqqP/11J2gi/tDHGsyYnsCa3jQ1xeXlCcKutligdg0fVGNVvTru2Ye0eOlXw/+SFq+I2WPAx
YGnS4yHKEyk/Vlp4Yg7Y8H2pAJMQqNAP7hycjz2aT/r12omVsqyanTgr/fji5FYmBZG6RiVPi4oj
nJpcksx8NZrXKHayNTjcs7YTdaBZN1yK0ru46GDaKOgXWA2YUQYoVAc/4Ph6Jdon/4NMQ9pd5LPl
+Rqd0Phss5wO4moLvsVovlgqVItccsljJrnjpjjmD0kW++pFC6OF4Urk2ccltIwgmnp+ODjS0a2f
XCh+lNlqgPdlrXCTLe5vZRY4qGUf/PgYhlJT2RNH/kaU81Qw9q589fkDpSTcJyn8fGJqYdEpKPQS
77Bqu4oUQZGgzpJ/0JLs7f8Jtqm50RuCNtsvKaveHVMgJGao7T/a+0l3LlttKzE1IxvDq+GF4JTA
L6IV9aPxLuEYYFK8cqwpvd64Ch1YL0di2kFqvvh4F4NJhuqiulfFHJOiHYyrVVa/gFDzGsJPDSMe
UdOd+EAgzWg5NYRcYa+jrRi6DWC7ReFmjrvhHYecRBDpj1F57utJ4zNzSuMueETC++4Fo7/D2KJW
/T+Meu6t1LaH/HpPQHcFjv5k+RLZ1L+W9mnmIS8hrJjAiuH6nM7BvOzWpEHenSXwc2+/BWBu0ZAx
GpNzzTh8TlQXdfBjbWvKxxrCQqdwAbhEh9kbZdBf9ZB3WfS3jaA7o13M5ojpJsVvWaLFFY+iEYXY
Vg3AqDd/SEEk216nKPmjbwbETJ+8/xTA8IC5OSiSP5pOiYN2LipgyO0lfrNEjWReLn/bpd76AoCF
Gs1KLw82THLQGJzyVPhsDj59kr9JTyxTYHAouVTZlGne1OxyopAknyyTv1e/sfnj8qN9EpJw+YtT
J4HbBKSJEn8ZSC6x7rPxKqV2i53LLF19kSdR+6xm9UYjc11wfDU8xVyTXGbGaLgPgf9FoiojitIF
5PLZDB8mhtn3+FY1XC5AnRGOKxu+H3eftRVNo8mUOAsKQCs5l2PeHJ/uMZxm7sncw21l3Z6AyAl1
BrPDHijwdsQkbNAml7HSKZEg35LmcrfgV96X8XaZHcEm9ACmXZMh3nJBNd5Hdhbs3rKbNJPy4py8
41DNlFVCjBwbbcMrGmJHqBYISYDLG7NfXOkKV4VxRPfeQahaNIgM5ExwpGxJH67qjvW71FSFC9BH
NHdJO9lCgua78gBMJQrgdNkOhf9OjTCZxnmek9y32ASXyzyuSPyOjqwNN/uGoPfqzbJpsRkHWsz9
qqin1PPS91UxNDZBfLUmtRNhJ/wQy/furephfnTDSrAYMmtnDj8jrTMcxTJBVFBv08HRQiBXkgPe
1tEaMpm2uF7ApCgwdShCZJ4YMUT7scl6MZLfu3GIcUeFQxR3DXLB7AsY7FJzY5TGcdhDc0oPgX/L
4p40EDbqiam1hvzAJHZ1U63JgtbzgqlgyI5geF3sBraSLA/OUDUabOMFu8hiJh3N5bNvvr8B7kh4
5IHEeEPlOhgGZcHQLC930Js+uRDJ3hDWLnuB1hcaHdEpdIOj3+f4oGUDRgNzxn9ALajEOj7d7puj
X+t22bVKhsvpDXKAS5bPTWiIab7ZlhZjC853bHKcEkKYeVKsBwzgc5mHpfH4hwUl0sxpz5UWa1dG
9Drj5o4d93T5EgYJKZJIXbKs2HnGIockFi7ea2h9SeywJ8UZJtnU9g3VlK/zosxx3bOr0lvl8dcK
pKpSjhT3GdUlyKvZtMuP9tJ3V1c+JJPsKf7QdHRaCR+NPjBjh2fEVQlh/rHkeEhR1KZCTHCTraiB
pl8lxraVIFbQYvv5AK0DiBwQ4QD5IFl6PRvMmwXde0H5fckeW6xppWBsFrCyis6WboeDi7uhIc0J
d5ee3hPYxfBUhavbCoglfwN/x36xY2nQjKcFYnEbgCUMy22e29TRsozU1pm+MElGBXKtjffqcMPI
VkHcYFXaZ1Il/CgpPCDZr1ju1qYmKaOjPASeGMGokCPtLtB8TaJs1tudCIZM+tvaMj1vyfyacsSY
yck/F0QVE/oC5WZJVm1k4kk6qA1FnMU3yHVpfaPxN6GXOIaf4KsVu0LYrPYIfHTSLsV0tID8VOEW
JR8ozopas0ylCAPbj+Ey0iYGjv+rQGtQH+PEcFRSgM+HVthmzUTWBuVsHJ5PtHprm4JmXLOswNB3
DVBJ22DkhRoonB+fkysTkPZx+llN65/gSXHxq9qwt3PypLD/5NpkEeK08oHH+uU5lBri8bKqwT3p
h+Zsr4MyhOmTRLjDQM9VJKZrN2xWAQvgFJ3IRohEMPafKUeom47tu2dVTUn8DhLf5slwAhUgeGEQ
e5uUppXTO+LG4QVK0N9lioj62xplc3doHcyjNtHI4KN8Zq50VbRV+252zdq3pCGPQWWjdnFLVmKa
zym+zsjsjbijsrfmTdTdM2OYcOnlnmpdE15u0oe2ifziaSigblWqyIrfdH73e2mg0yBFjSvYCFcG
W++xo0mhHIR1qDK3vzif4xpdPBcULGv+C3AIcBWBM1UyHy/fRYtLYXqv5T/YscHDqeOjocbhFuVD
aWf1za5lu+96KTNFXZIn3/5FPCtM81N42RiTFVyTIhT2CCsW6eA5uw6BuaEQPuODTvtqCy5NZoY8
ram3fnwYx+deCnpHKeF+mC6X4y7Z7DBg2OE24s2kSXzfSToOyjAVfGbPmOeIGiWExSwBEQd04cyF
pGDRE6af/nvAZ+M2vYqSq5pURxuCI3myX3QkVzByWwXvwUhNUcRKAA9cEw8PgGBz1WTIghE/fQ7M
vtd+sdqg3vKCYih7d/2gYqC8sLjNzVqamIRrUZ/kS5AycjzBEFiDNc/rL3PvEvHNBHjTRYY4PDZO
PkH23M/nfSI0adJWxQ/0SaPw4PDgJscLfsMOoyMUgE0jngzRwI4sW9oe5Kb8yk01fQ4+RGj/dmWH
STI8NAnfNxUDt6Z5PwA8utg+OiJNNepkS/uH4+zzz11qIPi/NrrwR/wSqMfh0ITwCBq2XFon7SQ6
89VR8fIv1Ypjb3fkHw5fYa6iycnqF1lqo6agmBmPL0Nmx+/mei79f/r7xeX4+UuJjDAeqZjC2pLl
zztR1QkiwAU1ov1hYeglEitd3ri5fgl4Z7c42+Dfb8OBQQmRXhYo7NIVMN58lB8SDyFkSdZPhAqk
GfEcym/CuecqpQtlEbYbMKi8gBEYqBU79QSI52xBsNn4Rui6MyTFXEDwjrgCVKFPGkP0e6lzTLmD
tjucfwucTFaL1G0Ptb2Q/Zd+IXj1D3d74+yRcuzsoA7YOf1RPPkfqUw29JNHhaPPO7BQfxXP9c3G
mB1sw1wqAHO84wSY5rgdyQ/a4mlneNlhsY2hmVJRkW4jl+nH16DEOGz9Kp+nr348k7jWEp64Wv8e
taMPZdduL8yGnHintS5pPpmErIMIt1vliIJpWNCZqDlC9WVvF42QN1UEXEkvnohmAtqIq9/c/8bU
zfIgHRAjregzGg8wUrBarB6kRGwU8e3U8paaWVy75/gZw7T6ymrTXT7IeRY2g+eYwiZTKO2y2nMJ
SfkAJN1TspeQWgdX+v6MEzQZSKJsbOsGdsBEqJcOSytilo0HJYko0v6wDzO4cQsuDPe9ZvSxbG3e
mn9FU6jmi1iNwHeFXz8E5yygwBWLyy30YQuR8mZvqAfvk5csJx5IMQXH4N2ZK+ycmiQTpI438nxt
FI9+Jp/rs8pQnoOPzWG4FLxqeIsL2S1C9up7X7lkyiFAZKiq6MheTk2OX2QDZUXjsESETInu0xVS
iqrexzl+BDBvXQ1+rLMBBmZasI89hy6y5ifMekxvP5EexPkXLq8JGq6njE1IhcjrCLij3FTzXiAI
waeJnTWAYDD9Oss2KVLGq/RrGdlL7Z3LkQxSJiJ+0PCJJXooAqjlfVTNQFpeunCcimgAhElhe7Kk
EwTTwy2aC+Gbv79mPB1vZZHcYhZAzCECX6mGxv2UNVn9vjgGdFkdRWsjJAQvsmQGTDevTlb2GyRp
Y1XGJbSgfNkWlhzGa+DOvg/eLSH4Xaiq5fJ/EFB9gZFTE4HV+g62+G3nuPQKfcBOGU+to7pt+arF
jYVLC/7q0BanSDXLvvao9UvvIso0UMGdvXfJ9QulbuD3XGssl5BogaqmOReCRQ3zhLW+Mm5W9Og2
/uND1FR3WHj7X69O0DRsB0YmkDrazOBRkjaRWKl30heGFMweLpioQCuSoTiTBehiYb87zXjjuzp8
ysPsNVzbfJupOtMIABVKnh9IHIkN0YaLtx9VR3pTG9CgKu1xlSehNXHvppPXo83iS8q4TJ0Pa/W8
lPzdSbrMJeqJyAPFk2aNYFt9F5133SMQRHYoRR3XInvVOtegIWK+f8wvio6a0hlAFTL6vNqiwI9+
X7BxBnVvN1z2xrp7yO2N0I77O7Uih0+TRkiN46gE+J15ywoAx0RgTFApi6xGdHzEEHZFnneGuOIW
NQMpsDGp4/HzxX7vP2em/xD16mAMqAeUa1fn+/1CVrjY5VXiY7zU6PyHIS3ObRMYytqHTd8kvRTP
ahBQyyfbK3N8OHXvUTij0PTWz5BvS+dMAyEWug+Xi6eSRsWXOShzoDZS9WB28HOgRWARO/8qXJ2i
y1/fXKkfpSZfB4aB2EnbUJkXpsNb05bb5Ysu2WUSKyEP4LkCe4gF39xI85xZu/FOzJoyNJosH9WA
HG2F02vDSKhxOqao7/ed0a+8/JS9IY0zcKBoPmuNxIE5/+gSlglYT/3HRUozAYOq/NboKZK4LWxE
/ER/Km+sXEIY4IjCbivJksNsqZ92P2KlTn0oKGNBKFnkEXYTVFBHU0+OsQ5QaoGs1P/xQU8vXN3k
JgiNSM1jMjUyIGBLBDLaAsekqCj1akXZdCl5zk8f4Jj5yzhGd5GdOhIxjqswp+VxIVCbYw07A8Nq
laHrzdXJUFOij7Two8K0IAvnqzpSt6uU0/dMRA4VJJWzR4B6o+Y1ngQNXtaHWjm8jgDp0rIISQbq
iw2rxSd+0DTSO1MVk+tPkgk9jiM52pdhqc6pwkMik8yZVB5YPnkKMFuMA9p4HHdsiQMnhuaiy4Js
YboNmpF8/mD65ay+OWZo8nNf738fk6hUyAjCSlcGYFu0K6zW69wjDm367kNLva4ZeVr7PZCg4uDR
wVQh5RfThpsZayh/9HDjBfUIyYRZ/YpH691RgixCy+J+tgPT4PEjNfYf7JqqH9mmRZqD0AtQTKt/
tNx6BgjHtjpH4fhj/UAtU8Qe+bG9tvkrifJPNI9slvPmYt4TDHG9VximuJ6R13rnexQkVQcCJpik
+oXreRnLjK56EMPW1wzcz9vzUUI0L56ET9LrCLF0NQOCae6/h8RizJWR7L6gULPpQFoez6Bss72M
WzARbxqGwJs7F/tgXwiKC3I8AoADstM2868+3MF68iIuI0AwOZjRAtVeB8Vs8pk3kFLTCJAZ5Jzr
rsEQy3d+m2TPDir0u3OqfFg7uQNn5JuE4d3iJECFXs8b7ab4k5ui6DLjvKgAgBuB+brLzh23TYFb
HDqcH376Qh+MGtWVUqT+WArirSovnUkb6NB8jDLeTc9Gl13qvD2yDlTBuhuaBDUcawQ9Uf9flZD3
l7rP4HbSoLbhXiwBWxzt9HCRJeA2vh7XCPghq2Q6Yr1POxd2za6OrTrpH0KI6uItAGQpZC1Oejj1
ZM/ldqoy24Hzbe1EDiwZQXQLDHREoQNTVtnl2lxoSFjj7h7e0QkfQU4YSmv67rRKjj+FmRSAcdOz
f7shzM0B01EzYnV6s5mhcKpVi06VwgAMKJqRopUBlnbA4XyFSvC//ujuOgQjLGkw+P/lBUr+0sNq
x/IrbLmh0SWHfZSp/9GvyBNF1QLwNDcGHcLI3MZ862LqTR3+lxcSBWbMB1uiR+FNCxLgi/v1JjDU
KVxlehqUW/5kzkTmBWzMVvJmeDzedaGdJGz/v6S/4ZjavYspi8pJs0t/vaLgC2Jwn3uPqxvRloS4
+ITAXkjZwR5x8KmCWRu5f1b8uMHETflxt5lvnN3MqkRzSG18f4MZpS1uRKRfGfqA3xiprqwBGWVF
Oo6MkVUzsWxQeZC3lJfGS+KDzXBRI+/vgwwRgAltrMk84Bli/1Tr9ZkzMgEQ05H+xhu2s8nluCgx
TexFvQrPbHc4sAou754dDJGbkbN9pGKQLbls1mVZlaPyUo75sqJGLZoFxakB6W/ldfrpKenVKQN6
fo/pbqImsam5WW0CO5YqgU7fzLCA7XmLNysd6iK/l/PcpzfiYPehuqsUc+rUi9Ezl/08OEREWd7l
FQcTINOCsca2iahbp71IH2Zpa+8KIgFeBfSK4TmjBv4sJ0tAoqHilTjZlYTXhdNePPsrDQTuKpDn
4eBWdTcsUYDjB4A5TfGQbdR4dPvaS3CgQeYJjVPM3fWeAiTlqk8xaiF+nDkodAgQMGJQFvHJzYup
HllQ4NYAtF3KvjuvSK38kVt/nfhMMXif0ZY2gXxf7e2Mi/CDy5Ah7e9d0fhxk5JU4ZF8nz7BjxQP
Q+yt5n0Nf6GaV0TL05qm8vcOy07FUrewB7KwGpY3wwcuHEnvj02znHachPBcqRxFBdI9Ujvq2mu8
sW5EwtC6ffhiVf4pcOfZCkSqdx8cj8+s/Rew7ozuoxJt9zoeVLHvInZZxuLzcdMhaIyn+2Sarr2a
nJfSTmR24AEDr2Wjc8bw8rikg8m5ihczjLL5a98hdOWCA8rO2JdwQbIq67RQ5ROMdZ4au1vQPrWY
sU32RQb8B76uS44dya+f6l6xhEbB4xYiB54AMZVvvhEXs2dhAsIGY1QWnSM4FHFDq/9NVzO8T5kC
HASXeoyNhKykTFsBvJbt06q1MzIFK6CxMwyzJ8+VAhrtDeRTI+xTmzhalkuORQSZOGYnJJMQKSvP
XtI0aZezCvrkD7JO069ANoWU9U/kRu6efAl1LySxso8m2eDc4ad2z/tsjbOEkLnoNLNXyMIQmIDX
MeOrasV01SnEQ5NPXAOMQfLKkwIIS8JJwpVnVMJrQEc/8H6XbsuPv8mS4Y09C1jYDnX9F23kSmXg
rCd1R9rzpqroTOa64XTgxFXnv9glX8LGuafK+ZEHeQmhqABN6t3Gye0+52EN3Vtb5WGF0e2m2eXT
Y80QKJ9iRuvRe0y23ivPX1SNqaRTnL2m0n6jizB1dAIsDdxM1JjujRu1Yf5U4n2p6rGSmxGFCxYx
XTt6TXIdnSXPMCmaCoWyvyufTN29NVuaVe1LC7f6wySyZ30lI2tmKnHS3A1D2jqmHHIboXBLabw2
LoU4lImPhoh2iIJ9uaR7huVafsJCGDtWPO3sM3/9HmXX/bPmYNppyyRsIe0WxQVldf2yhIUtssQE
Jl1oCW5hnFTEBeq/KFgJikwmgrgR+qzEa6XourWkayYwp5cDGsNQ2XPk+DcFrYgmIgNW49Ulk3io
GQvCNXg+V95eLAyeBZ0Pxs+q4iwsguzMGgzmC3LEMnrsDzrPxjhAXFTW3x93b4iRY0ksCaF0bq/2
4Ei5JfoYKb2Dszl8gwoXguq+rAtiW7WDdoxM7rcRB5QwO+kJ0kZ8jfUni3tvR9l22IYTzeSOZ0z0
kA3ZXxvAksEt3pC7WoB5D9HFzz16DhCC7NKA0b+mdwetx0cI/d+uboh9Aixn2RSpbx/ViYXXljyb
x3pNzhypyXmiFU3BWm4S+YTKWHMk90QDNNbgjvHp0QFc21rQdEgX7rKIrxkrzS6oeXWHz2o3nWNY
38O7MxKYnw5hMnDPM2VCYNMCmjWNQsABANuIOaEu1+WUMegLY7ObkrLeU43gH+qIqZk8KWPeSHmE
wdniy4Qpt/gwH+KCc87lIMwiLqJlw5QQq2ZoC/VRI1+a9Fwx45hO4bZLrFHeu8yDSVcOIHJSlBo8
Zagd9e2LrB71hi3ZSm4sB9J69knECtunqd7C3kKlWKvw6uAsFBK9CgTv/8kZtN9HgjkAxyzgIJmw
wskD8xmpOSLSevGaC3/sSuWqkqcACI3MQzY1YH+0RRkrUM4RzqbfCC1C5UvtcIiwXZwc8BlppASk
GhKExg0K3y1UIAIhIzOUW/khMrRHcxGgHmkkTHMhbxpu25DfmNpnyu8Isj2mgnAjv0pfJZCp2gTh
DQznbaPP/+OBRt8UBb/QoSHVXtDL3HWWetwWNt8vDBc+9hyXqGj+RvztWY4FtCmcOEfM+E9CvLvY
Mn/vn+ibhXw/8tt8A7pMFJ5LLAelI/quVHuCpu2bfkvZ9naGKA3cLh2FRZsTdwoeF8om/6Z2FUIR
KjcrnY+M+PSCMtq1gYTe7925H4rgSEkgv9tva6sdl4r9j/TysKeVmrt0PXbAU2bDNQ9hjjKa+EBU
KYtgS4osGlYsp7byyDJd6JjQYw58jCsBJMBgfCrevQnE00ieyw0Ac6+ayjgfF2nsFKwaJT+lhL9V
CtGv7UzmtRDF0EklK7eT7lRQ5YbDxzZqAJ9R/dz/BNgiN56nYAkxIo2eJQd1RSeOX7yin/3sUuHq
065eA63hUsCRK0zoj26UGyTsstXNDq7AOoqegH9A2s8CUuvarEjqCFms4B+KzSU4e/GXzIaeRDf6
c0+lWAOLW5P0ZHT9nlQEbVPtxPBMEa5+F0TITI+UcY4WdhN+nU7vE9qUWCh2RYxjDOueqV6lEMbw
eqr5oJ8px7Fyb0wUPFk5YEKWlcKmS6cW6cvIs4E6B9xsAEQ+5Wz/Q1Jg2mMjRv9Rm4Nz3+ybsd9c
8wFqgsHept40x2g46TlsQXxjIPvZxGdnVe4n2SJaMp4/rZvFA2P9MjfTQ+bjWbD66BE/J9XRmhVP
dvO6F5w9nD1lvaXipYjy1AU2W0Mj6Gj0s8+QQ+psAQdVtUMg65vg5IInRjvPZjShLMy5nwU/jLgT
Isvq9qwTOokt96ZeXYWSjC0UiUVo3roEX8qvxfovBBo+lcJ3016woZFBlHTj4acEhOc1ZCz7syqX
f3DPrWfRV88V/IJLgkgQZdUNCmjPFmvko9Mnon42xUgW8ZO2yDDzAkPjFlvGSw6+1YAnZiSM7Vtj
A6PmgkysbtFH263x8u7kqj/aAmiRq0gtnJu1ZV/YXTtGSJ88NAy1aGwXHp6WIBpDvU29OlYyyG9I
mE6NGwC+so8ZCqV3ZEYQ4flzZYdKS9gcx0Uz3m29FGY8d+PUis7PWS/u5Ut7vmuqTxLFXJDVP7Iw
Yw1QfzjsmvmvSf5NpW7hL7uo23Pf6fG32Of5y7CYQ/xvLJ2OzEbQ+bq/heACq5xAoXcd1Cl/fweS
S19Ax7jAHOUAwDy5l+ImrxbTOmtipfby0RW97KRkb9hD1sS1g6SKdK1vq8KxKou1k/8rFn50sVJI
TYsR4xsxPuqBS4GIKhzqcdRH1EPe7Z4BZdClO26b29ieuj64Bm+PvLWSi+U46IpxwL6w+Xwe7D6g
Mpu8GKpPPHZzPcrvalpLpijs6OYjFn8HIROTXV3KUwY23CJBnhDmgeRqDkE6JklSN2cZyDSRVf6t
P1eRV1rb5FkXerWUfT0lfo7N2JwR+Pkrs+24eL9By90PKhXulT40UaY9vHVo0th+AZ69k1vqdX9o
aFtxUsYlRoIW+34+0A+AvfpbgzUkVLiaZILfUQdYG1G+cDhidJpS4+1B8QhpGwFe2WCuBY7zGgUe
xB5tLxQid/qL7C1DgjMnGxRpeWRmcPR3ZI9+jMBqm0Om8vIxhVLB3QRMnQ8jqiA+5UHZ6I/v/KoU
u+nLz+/11PT3NPXtR3k8GJvu9A3/bvEW+YmsiNrID8FQkLhJAv2Ilx9w3sQf45GvxsTQPTmCkqug
mxmYDct7jBTlakroLsx7MwjIjlKUemmsnvjVR5nJOXu1rZVaWe//vS1aJu2Lu5gLDvDAf4XVWkmf
eX59SOSO6H2jbNRcA8+JnjS2Y1URbKNRuiVdBVPi05z2tpLrw6FuTFKaw+JD5YYYZ5erbJdPivgW
OHjGtkESU6GVA5hBdxxrL9J5hYmznBp3lN73EbuK4V2Y4M4Xwto9C8kGQokZu3bjnCR4IkUHNQWF
KZvWcY8mqkL9hejUoEAqyd7748XTlR4Y1LvS1bYs0BL7vtTq5JmxdcZmUxIRMp8PCveSlSiwkHZg
HD1XeNJ2jSvACqf86+zCQ+pfoa3F3s38ROZ6pPiPLDUXM/7Hi2mUwre7eXF8oYYr43kwhereVdrF
L4rueFeDglKa9b27kpoFXhxxAm7iDZxZPDp8qKZB/XzMJjN9MO+n3inntDqAMZBeHEGP+REKPtDf
dwhSzfUmaYGiuOFg8GINcXpyf2P+TKxvnnmLH2tmSr8V0KxGAtNQV7K3lmIP/DmVfbvXfRhdNISU
5BOJ0EA7ELG/d4WJ2hhCDKNcYtslpISnzGXE85Nm8j1QlDUTTDWV07RcdrR5nXOVEQAteItPYLil
gZ7cdqRewS35m5XEhcJOOKutKnWecS/YXcHhpzG1+Mrju6IlYeUOjJGku0LV0+qc/j+vUNrcUa7w
SgJ5in0Ss+guGmbCmSq9sHW9BeQMIqoEDw5X02WqUpx8yHDBlATYiFwUZ8iSyZFradCsRpJnqfJg
NppLkUssp11Gha5kZ8taGUNTA9KZMNu7h7KFup772EOZMvRpDh088yWKa978hB+juAKtpRTq7oGg
doDesGVgXxkrGZIYDaj6/A+KN0nlfCyTBGsPIiZWNPeIpCXYnaJNbuztt3mxGFQvpCQOYygB3Gij
1N1c7tYSKAyUYy9wbkLvSW2CifCBrzYeHMzWhbdOCdUKV7erso+TL2QaVM5Xs9qwiShCrWKd5CSu
n8+OFIlbL0A/XDzpYDRfkxKciOqbkaFvu0v7TrTMddlxcLj+eOBB918xjem+SzCQEdYwjzf9eikW
QXHjxeuzDJSfYgE2oIekK/rsFzWYBnQdW51TA51iewByLyioIcdADp/oPIHgUKV4QopTzH+7PvEc
T/fCsi18LVJJp2JjJkqbMUFrH/IIe8YUZeOe62ng078XJFVdPT7UCVuRkTAY3rHNz8xxQODd39yD
xPXQwDZe4NgNpJtfV+BcIgk3vUp4zyoD5j5RRar6Z4vvr3wk3GqaXI165zqMnwKhiNT3XDyW503s
gUpbmVgNls7ZJGvU1ool6eo4hh2f+DMEQkK0grMm4V3Uf3gx2c5ucn+4kkQKC5zeSM+nYn2H5Qt4
peSFNvAMz/LwxQfVr8W8E4EWXhSnBbfCba371ByGmy0taIC2pYxtqzR7YsjpC1axKxKKKRMbWlzb
eF4ErofFyRxehfei257faSn+8mHZrfGi95GDHJHQBspT+gm21DjqsMX3aZbqTw/nDremmWpwxuZo
vTSVcVlBrr280Wf1NTNqPpWdTvUkQSTIFc/r/+jUwHWLo69E9LbmlL2A0F3HzNQvqyY4B1rnMTwq
ZsoqnVQwsFvnCUnvQ4iBYoSJyeoKkr3sUtGN3hcaCusUr3HUNXoPnB1h655bg9CJ/A+pZiJtnyEb
3Dc/JhRUZOKcpds+MBlZPmdvYOj8tEjTMkogjiJ6rOTk2ExbCogadcddto7UFsYcJIDuUPmZ34nE
+98bvKUJinHFyzEDZA1aKKAGsNFEnDXHstlzBgCj++NYuRx7BdRefR8zB4O9/6Fr3RVIke0x3ayZ
vBpvomVLzGqg3MaB0DVkTiq9KQ7upPX+qxURnbIgjNNEVzWYUwFF09dW+6Qxjk7QPyrGPw0hLm6p
padW1ZucsHA3K0ZC0bUd5bTe6cPGPBum1jxwRi+hNmF5YkVg0KJBOjqnxu7Vau5tZFXY4VJ5d9yB
RqY2Gww8syPvDigv+E7MJBeI9/dCADfoIqFBt2v2nWJgtEAePURuPTJzmk0fC5CcLMw/WJOFT8yV
aOJqoL7U7qxVGKTiiIFfwSM7phSSy+rM6syfZjbtmLcA98/M6uh1Qk/wes4dNJ5MXmC/wDYugJoe
kKRp3VPyZwf13kV+xyUkAHRARGN0+jecZQd5QUIshDOcq7mH5bUeAkReiZUyra3zESAY+xluJ3DS
3JH1ZeMLTVa3ctyWVOJUo5PnONU/fpEoodWdJslccEVv0UMWxZUrCKNf0XuDy1U6XXe1+yd9Vro3
L5mFMLSbvs6WQkOnsznioBdLVhT1syghAWIPoK30V+ZSWmGWGZiCJFUXRqqfVzhyzpkvx1ujciwz
cbWIa58QP7zN3D61peRIS2LSDULLIoIf9aOmD0cnHUiPOy9a+Nd9L/8ywSOCGnyRAfqC4+CDcTJj
5gUwqKkP/grbfPEKp/vdftoyA7yZkO+T+i8d0ae+dxJBo39BZxLzWA3Zhamn5fCBvDKCoSjz2rT5
cUSDDeHdx9/0vPHkdiTMaweEUVCVxr18vEfI1U1Gc1t5gDJCDvC9FmVy0/+fMqVEK5j8LXOBmwy3
f6GqqBuS/hznXtSvLE7VxsKtBXkIMJrRKSsdumXcBwQcE0YGfcofEsl3RPJY6oLeJFKXJ3FB2j2R
4JsjWinpsudf64BBBKLeUYeJndpjeB2N3DGYDVC0THFNzu7L2a1vS4pRkVqdEjKEDsknNU/KUOe4
BNE6bsBQptLOwGtsBuppI9ftBeqi/sK8gIyvbUjtEIVHJ9IUwt6RAl2rQuNxILYdG5M/rL17wyEp
0XKPFr+cPpYqckkUZpoLmHMqibvSvH/YijAGpQ9vy6lALIzFOVzX7GCFJVSfMzPOmG/dGKiZPTeh
boWkSAgV69EUCykC6DCMaYO529/cjWp4xlanKQCNH8u+1Nfhcmn5CDKTAa8p9Uk7pwoC07jkh/zg
zSln/lOgGhD5s50GitI2+/8Ojm4kuu84KeE/Pqr3wX+kFh+GV/VQn5GE5+tTPn0xwbQzgUd3o1Qc
YRovkEkqAqZSw8914eeB5UvrNtr7pIHFu7hFk7tQvXoFCAj3GWjCIRqAe3TvkkP8ZqYPCPSKOxda
rXVI7Z/hmHVp2sjRF+OweesBz2pAjL/nmE0DbXS04WazSzJTJEzOBS1Of4YGK6//m2L1/3mF0rTm
cFV74mvLs2lBEnIixrB3H8eW0IqxuQVJMazQhTUxBCDYbjhA2DoMKGQvhk2H4AeH4mwyFYKwKYOR
dMnG55UtK6mHRAoD+XjxTTU8KCQrfjzd4LrsEeFqueZFvwlyYrE/JivPl1ZfGrNk/laf65kC1npv
Y5203I7iB1C85KTQPvmlulW0optxc3nYM8mka831/7hAUTj46OOcYf0FnmH4113B2EgrSROK74VK
lm4F3gwFYtOwU8uzQkPYLK+0VttZyIZu6Is6RaUDo83t65XgNhn18a0DIdAMj4l9xtk+FAoeRpwi
qQq0lrCCfY7CiLzvMG9ds7uUmfpjFMXhzOC/YvxBLN17Rc9C+E0MPO9rRMvNRaSdlsT1dLGHxZdU
z81l5i/Bv0j2Jzsd7qSCAEwAKhS1VlI5/poW8yr5wfT6QmLsOYuDypiBJiRFzLlXC+wF9QIkjkGp
gmFoM0WU3KZ94mC1WYGMNjfZE/Dai90B3Zu2bYGin3ZVgvUGwBexwq+DPS+OTRKzkyADS3ZxmKVZ
+5wh2tS8+aE1B4gEkwyYioG+YyN0p1bm5OcILqHmlYaIMWaD6mRQnGVy96vrj42U0KlszgBsLeUp
ZD4ecKUH4L973/2ZaPvRkA3Cr8LxEs3AZ+6XpQAANWpcWml0+F4G8Vdac2q+oDt/PG1xCHqi4q50
i+HxL2Bl7i3MPeshhiKCVxmaus180PSrEHaF79T8jYtl9WVxie7vjRxqWhA9GtevoERQz5chOJO9
g2ZA5/PIjM3ANiAaYFu+bUzT6tMpfpP+Pp60bq1RpoLkJAXrBOyWXGoK+VnzFiHrroCTa1TDxSpa
ImZVv0QuF99/gq7QeJ93GJoUdsPb+OwL4DM33j0FG1cuZDIU/2jsMC0t0052LYqtVvKeR1KfrOg8
OrpyQwrVOxwuPI1ACpJrjXMqwtM3HFpB/TZFrVyleOXJj0Ez1OOX/V6qLPVJKBb4VhrfoxP0kGiC
szDgkHk26arc3wsorPAlrTHMDE7VKClsInPGRyWL9BUO6RG7cRiSjEemMi9jACkobVGuhPm2kg83
CpZV2QU4XEknocbDsvTCGWVOnSjrT7KBpjS1NzPEdgMHvECLdb3LmxXKBdUcqSgS6F/Q/GlRJ8mI
RfomAgltw8gp7oqZAKkISv97ZXMIc2qPUUNE1p8T36Bd0V4BgdE4vW9W54+EQ8rb6ToHYr/LghRH
S30qvIwulEJPFwywX3k/Tq70WcA4QpZTbYwu4NgM6YreQeEOqRc0bafELZoz5NEWFhE+hpA9Q+WE
nyk77wx6YrQe25Ld0BJtyWAnnywJyS25ypHjQBs/KsbdpBNOulcKi70TfgZQFIbABwWz95vnGSxr
SFOSaCQ6CenXc0zHUCb0y3G0jz/8r6VT+4X/WaAAK4z47V58I19dZkIULUP0vT8KNsKq7/RR8wTG
CxCag1jEh7LkYQvGeVMi5NMMAws7jDd9L7Bkgv1tdLHybO+e78y2xsjudNNXsPy9p+ENA8OU/BZ0
CrrljtZe2KNnFrzXmu1oLKEltcIYpYjYbTArvM8QoGI5DY+BkOMtPnlbmz9LTF42eauqiAkze2yH
D7XvOgTfOiNQz81zyP90KpwkAmuFVRBJALT5fhkCmboL/UCKUJvt6Hq1gwWgBmTR5hEfKJKBg5Z2
rmJ6jfqE9Zz/X6hKFA5nDa5EpUSwFNpyvxgwRBU3JwUQBOCi9Epf0mopMaXqI1tVrsmhq1VCKPmS
lchJMSsd3pu22k1xWXMSGj34aNW6c8iKIn5B8WZAl+5j27NA6m0zdnVCS4Z//K/2YUF2s5cBp/dy
HtaBMbBszi5kwKdzAwsi0pPBgcyfCiowktrOZgwSCS6ij854eFJs4+MQMXH9dwkq4UaiO8/M+3w3
CZBiJRP1zQvP02jC8uI8ditFuqfTq+SDFM7KZm0U4O8EUqiUVSHENQN0PAEPl3vyA3AdZ86ciwPy
PCe0+BSEzLZ6bMmmCnQSTWCrIX7YwZWSKeB7WaFaDCT1Of7JxVyZ0uAm5ouszQEgjHt/rAq4g+gM
h4Nq2PFbCV/3k1vWlWaQWcgzD7T2B5l8u//cZae53uscJ7W05ROSV82xJHJZL53sxLQvWNaFBIJV
UIjcvqGwx4Eacw4T9XEfAwZLuZfTDin8dhP5IrRgyGBvX0PmM4X2OBw2qlUmYk85EAXJGR2Ujzd2
QWJDUXqGa/lMnjuo/nginFoi8va50vv0CO6BdoiEeRsygCyk6RDPDDJML6Xdr6EsQ1N2JVgwfQD7
qY2G6uWuYCoWfNz9YxdCZq0Dcgt4NaChXlkKNUF3WhUxfGb650xxdbtJ3DQSlCNwLyGavvX4Jh/5
MnSAmhnwnNtEzD0h0JhISNg00g4uI0CLJ0lQmmWguSXIYcBYxIqbNpbCfmJx4V2zxich5PFUxzxS
ZCAQS3KQmb9JsyHr+XXMgHjgxtML8UtROIP71R2+1yHrrGyHoc1dGV4ImcJo+10SRLkHoNssRN/D
7jGuN26JcWiBUubfUvIDozBa98BKjnwXH8HpDy66CkXhPZF+T3M2HFaV3EVRkEoXkBbOhtZyQnw+
5iZuNYcA33ScEaMC+uvS8pjjWmhObXfMMsp2HIhpdlhIPi3aKDcI0kzS627zKPED+5dtvBCsLkl6
ligLmv8xDiuB/i1r6vTkpiPEiR8rWeHR2Y6emHjGtwEomdpNDZjGsgyNC2C4kbLuyVDWErUu48b5
ZPUPLBEJjPfuyicqg/W5fgPimBx1hN9Jr9oLihp4rQY4G3FyUU0zmX82xPSh70YgVE+hXFuVwBP5
0kQOeNvtybiv4EtSLKN+8+lxnPsrSmrzlu/9Bxyzs+3QkN1/97wliQ5lUYp5KgOUsKQWuvYkWWwa
Knop11U+eVbpFEPmPt7RSqGHyOa5svf6SG1gnQ6x8ORGa9HVM871anRHDth8/YTDTbl96OfllENL
bfJhUhyQoEOpmVAVgccNmQVTDhxkINufCqeZRA1YHbDMJfhpZS5UtPqm/5Up3uknn778d2m2Bl1R
koA6KMtE/b9jxXR6sFmW3b8IIvGzq+zWPsMsomPVBwsGdlHgifVU0IJ8CsBoWr61ESeCL6DZdFgw
p8oNON7jgdUh6YQ+NLieD39kqExG19Cry3z7N7j11UrSetN6RAS4D5dErg9RbVJtq88qdk2tklj1
5z1PFjx5UNKEorF2Pwvwed8aYPo/Kg93gBMb6TD3N9xWOJ6v0qir4/BIyFOrbW91uyOvwKqHu73i
O8lLrAqdudbWnZ3k4hPfvIrZebMSoJxw9ymsL3mUZ9Ndg6C0R9mqUNAzEvFMEZ9iFNep7MSzOguF
6g/qwvKLjJRLbCe85BhM1JvVarC/NCbwgqqBgTKxnQelkZMPeY+swrY1EGBtk+dUn50UK/5J9giP
Yte51vscib/bWqn+iA6nratSedxbIQwSDnzoNX5v5TqI2HKZxTTebov8qG8KxLn9I/frF0RB1pwu
uQ6BEotam6LeQElSxJZJ+WJYFXwgQGCgDNuhx53cCMQltzZOeIyOHXTczo154eGuenJyrM4hrliW
gNaWMr30m4y8Fr3foM74GDykZvLHYCGWnZjsitHlTYjuK/idF5mPg67fpKzM68kCubRl/Sk3n9z3
SAd8Insh0xSc0rsF7sW2fbah3vvTE9sneM7BhhW8w7SXU0Fgl3SzWjhubpsWFdMg7yQvneWag++0
3kXSYREe4TCeiNny7MOPZkX6x2ByhQWRsaj2oWftvRaXecG4K+htYXpNxDbclVa+l1UzSk7ULmaD
KGDDnMtCoA8LzdCDiQ0UafW3Xkfmrno5mri0SBEEqvSmuR1r6kg4blfPD8l6eE1e5s44Atf61Kbl
uVF+Jh5P9YzfiOC5kXiUNWj4mdaD++6I8QJrJAaG9yE8mXoqEM6YBtd++NHpX1jCPXrX8Sl4ZENm
Brrao8JGaBFyaZ+AdekA8SA6s414pORcvKGgTKOClAX5p6NYlPDdp1SpMViaO0M+rjcnsEGx27iz
cH4AQ6qqysxs1bPc4xQ9kZ0H7OE7lkhR7/AdeIogBC5sxRGpioaJ6lEgtXrcQVyNBOlO67GvPBTa
1jFw361iA/TPGcEveAgf0wTcsTZanC4NksIhUFZLsgEw0EH5E2zIcrhPSQ94fHlkuJPJ0BBMP7mt
zgAmBPXm9cteMEYqDSzqXHVb+hRKgQDIcrEoCNWI3btJB2Zx+rsJDCVT1FwtV3byFbQn6pXQm+cT
0741HX++7TNgYaBqya8lVRxO2m/hYn8QCl72ICrAHHdNrjUIZmfskE735Qz2pSnCaDkuO5Ejdqgo
OPKMHIZ32Q1WK1lrnQDPQed10eGJurw65BIS0ozWv3j4Fe/cUANgDnS2Zd4thd6UC6wrvJ5Mlq2a
Lpx+4p4lZbOp+igH5EoXmmednDGXnC0jSla4+7BD68uLRGp/HOi1kRGw/E815xUaRXdpbzbvABA2
QBOOrPpWMCVRezWg0V5JcJNdjOes/xu/V0Z3/1cH8YoefJfkdR4uRSKusCRYyOiZv8XqGGh2aiPa
PSqKhh0oFA6Tze4BFZHkHt/AOFre2HmJk/4d7kk6qsnh8U2eANAgk+mrAU5k0mOXd8RAcjTX5/XA
sG9SqOsHSf3ngC5F6MwZvgMNSeTSj1P85+8wyIXf62OSlg0VimJpxv/Ygd8ACC2IpQN4Bf/9Pemu
/NNiojbtSUYLlFiGyYwNp2dg8JzSzhKTLL5ccFAANL/2ykADZxnbWPM2i9nTXE4qFthOmo++rchi
W8V81ojB+3jXJk5kCITcqBBgq7/VLMLXGrun3QbA9X14gMseCcyLuDStGwH0Q2J9NCGsD++2/Q0e
tv4vLpYMwirG/ho86bUtb9qtutGqUeZQw9CJFlrmXlCqBPU/3OJNF40+8+caswsYrr1unypTVECe
AWK7SbpYUaK+zQPR7xHFYmgx92jaXXQbhYChLq+OsPRe2XzLwvpg/byR638Wh3VJPr5R71EvhHpF
MX2mHFiivLibUAmEUMpXCWt69bH/tLRKACCilcXNIAhHcoQEtzOWXZoCfL6LePW8tHqOFhM3Z6xb
M6ARWI+41r8hgFlel2vHoUxwnsKSJve57tNoh/R03ppFaULx9QJ09bVplyySz98zeV8IN6NOT1Ad
bwO7kf8IaPVOT30o2RpuD2kvkXtrMnZ6Mf+VnliLROWRaTFsjtfUB4gkTcB+1E25q10PN5hiwQlG
WPwIX2g87HvsB83fqF0YQ1J8q0VVmIjy3ZwQrJ29Lg4w4rVWtMK4H8I5hGSDDD3nN/GNcCVXmWWw
uhCfhzF5i3QjBy9prF9jGY1sRNSRayWjMg4PQQqyLvMJZ5efPEnSQMRjm8MZMo0hKe7/wTZiRxBP
v4ySrMWzDgMAqgInHw1EbbSieqwTBzgkoQQJAFsqDsp5NufGxMzNGRHo6qMQpqB1CI9P3IVnYGnk
VK6ILJSpECeAKVwTTpbo971BKvZiNoGC6zofrfBTNyHGKBKAkC/eq+D1molLPN5vXlDI/KRoOq3w
4ZvO06PjSOrt2E0MsufDlKTjJ9rAGP4WCaeBYSE6Aqw6aukeuyVqQe/uy7BlSqMTMwI3Dd1uRUh4
ZUKVICs7srH76M+aX3UMe5LPz+OxH5z7+8DweGqGDgxuNfYjF8arQukBnvPuVMQHTT/7Po2uGNET
Jw4ny5w43t4T3rNqjKFJ0+qnFhNZE0s9vb/rJ8CdgukNjLsCvWzWYaiseUTaygYdi766CrHKq9sW
pqVqOsxEHKDBceKiOUFo/vjHgnb/tY/3TNyUfGr2gpWIpCHsi2NDsHEDOZkEKNvZ3MGyEOLBqM6K
7JLgN7fT6PAj+9qBNEaN/IQuJ4FedKDplcOBaBgMzozi+u8wP8ZhsTsnTOm9VVRQ6ZL+A2FkljxB
xQf0Rl18i41kJU1cOrgmwZjOl650iIXMf1JYEEZsh48TUiLOcmFbZY3cJF4DiK0ztH3xv+hG2Gba
qnKkZ4RObMqFUwiiNS2A7YeIcctQyTKt1g285iZKXBkTUgTw8rMx1T2pZU2CYwtgFuKhP8eGQYVl
NmJh9BXeEmq/UssuhnD37JILO4ciZIjJzG6JPv2GfQwDdYcUfNJhzyOdWf2fKEsgU2lTxYRxk8Do
arb/3X0wCUFm9nqJf3M7vjtbOn6SrrWeS89lxCXSPp2uozh/mm37wP3JEFF+kOn0MGOXqa6pcSJu
LQqhG97QkYAIRuqbVYn9bMSq/JjWqwyO3LzB+v7AFF37NWdiDnpDXs3VdL3mriDMuXzRwMTIYaGo
2wizqAbz1gDjrRfEJ3Y1QN2hs6XGw8DwNDkUZlmp0touiNay9Ye6UKuMcPrhSt7DNzk+3V7aj6Yp
VFrEgdEQoGzZRII9vC5nfcDRNbJ9bUIIjrYyO/ywBPlWIMPOrPlgMFOCH3wfPRxUskWLgOYJDxuO
8PJV/2+BzGDy251hBrdbOl8O6TU8qOZIrponWdIDdm9UR67tyhHZh6Fa2z1ftLP0JtZteVthCF3y
9E/ZcgOOdkpc9V4uiJq356eVCzcv6zH3+NDzRSDhQ8aiTWFRcyWuXACo/YosIiRmmziUxQivgcJl
xUSgMkRpxqFnK07RkDKwgtqcA89D7EbjdgZJUTDpI9Zfv0V3S+L6GuaoSzkUw+BSXHmJT240u9HI
Cv2sbIZ/vBT7eG944JDvJfnGTeF6WQgMQqeO1asW9xq9YgXd8YHvU8/+sAJaijFpClIbiLmmV0pF
1UmLZh6VK1jL5zA6K7WTdwlzHUtl3tZ0j+8KckJF34RLTrj1irpUCv5eIpkKUvvv0bR+6QZCvykz
pKabWKm93+DceRRZIFq7JWI+LaKZjc9xU5ip7PS9iWkuBkHyJt60PwE+koDKwO363nI09r0D9Jea
ZdHO7ClX+XuOGlScYn9ZZUFjG9sNj643nI50uUHalQEWaer5rDq1bNbHhuqEsL+adG1LURPtuf0V
EqpUS4upGo3KV6dWPxD+XqxMk8FarzHkMfI1PKF7ZIPFaLZ9usendKhcWRfvk8rSe09fFAYtyZM0
XNYopBiWE5ovOLn8WqpW//6SnK1Pyp7OT5+dsk/kTYL+99jnXqxv2Kw45Av23cImcnUwiXPoqgC6
PqC/mmCaIJuP4v+KxLsgrit0ogamvtvKYnz5j1Pkz7KZCpbcWWgKMd+dqSF4jLGdruPBL+/Z2PdY
MhJO8OKNgJQKo6r7gag3yphju0MZdfDXsr07TMoS+0EDMdcJBUhw08BiloZgqYB7pcevWB96OaiQ
goPvZc2O1NSjTGAL3mm6yMX6uQ5+1iuYkyRZd1EkkH1oB+S1q4WczO0aAoQks951DfWQy3uo4tjX
m96VrV/opH7LzQaQuwNs7r+zP3oWQwblTcVHPj37vXXfTh3Q/1TvD5cykKtkzsbHVi36emoyvyxj
7pV4rr+d52LR+bSxXT1yxspn2OqJMSIKooKnMPcq+C6rtMU/4qTAI9WIP161T8b0JfD/f8M1R5XV
eswqXbzc29whOF/1i4QbnKB4EwjDg3oXFWbmjpRPyvTUM6nS77vwiKMsrnQDG154NoTclL+vVG5b
2mDIjNKAmxeNG5zRmbKnDLKZTc30LW5TV8K1v2Fb+Fp12XpF98l/Pl0fi8yUAYwEtLhPOnuvi/f6
jEuO6G7W8+QGKJczWKuQEFD9k4u2Tid2T1FZN3YWodAUKF+nqVWAl9m7A7nH3REAQ7dJ/8dByA7w
vYD8ZvUnZtu9sZXWaP9npbuXu2VyAgtEoGakYr/A/feLfN+70OKVnbwZ09hm8LggzjF5A0GDN8xx
E6MPi9MUmG98DEOmvJgL4LWo1fgNMW1YBFivFex/7Arch0K2ciaXp327TQmEUqB1MkVENaKiqXUG
TDsD51D7sSTaiL+clr3Q8rgEvuFx2DRUB8g3FA5B9N1awPRxt5ZELoRdCDYBAD7Q6+YGzR5VhUZj
7TxoreIk6wfyIhsByfSyvUv/y6GECx6wPhw875LPJiOTTLeXmyvZolZIueCI2nlkn0+eTSAw/A/w
tbwfKIBv8xiGhpRhapHySgRRY8m1EbFizC3kP0oY82LR/76qyvrp5QLuXJP+yWt8dfOP5hT1FuuQ
eC+MxlhfCoDHgEKYdPfiHIJPr3nc2VBooCvnqgjcn+hKdxq0Ho9JxqR4+IPvdIkEdoVFEysvZ3Y7
V8NkIQDjvkYqoTNMBGe1pQ2jf5xTDnZaMnWiCLPBKvdzIFyRPTc/+9FKmV9mINvMlxXK5qYCuDp+
L5h8jYzelRjdhg4PPVZXkd5xCJbiZ4sBdomwiMK6bdf+P4hl48HA5rfHNp1m4qWuFV1mytLm8lSN
IuBnlZNNsR7rtkDQfnJUyMD2TP0SuYzUykqRaqq/zhM98Sux81UIx3FvKqjuva3pN0pwcCyW8k0T
jgi8hfNJ6zrzgibd4lEH+D6kg/09KX5vSgjXpbNNh/MPp/R0Vg/gWTOCyiP/Qk8lGmO4jZKTXaLd
a1r7wJ+J1yt2VfTJh6gsS0oUemE7yB/q4cNke8pdC5Zw8CZa8X5VUpdXNxG7l2lEndb5SlQHR+xJ
5s4ppP+L8s2mZOYD5h4yCWG9m+UQJDJtXsbe21x9rjmnGzvc1c2EzxUmZ3N2/ImBQ9R5ye8FG9sn
eAGukALH9a6XH1xZsnYAjodKPvMCejGafCnNJm9x1gmP1q7BgqSyNY7IWchfsEB78jw+N8wgPARO
jbvZ2EXA0xOnU+FL+740WufH4mRchnx1S76i07SOSbcZ1NZ140WXW/H68b9iy4EVH7o5dSjRV+RA
dUdnrdEhBGJ+RWa6pSd8raMmORQmB76HC5iFtpDSapMeGVSSdWiK1jeQ0t05fXrBEymktaaCY7bM
dkoKAH463wAD5Y1y0t6BbAn/PpLpVSppgZ/+HdjeYSTVHtURjHg0uuxd4d76MqEQbmR1lRY6q0/r
gpoWa/wO83NrfamCOXU6YSVa5aFTWOW1PC5ZkIF1IcRNNGlCSnU0nS95ejLaaow1eO/Oao6gz7CS
aUmACEVaRltFbuF5X/hIfiZRIvZOscg3uCXSc7MhY/BNHfNru0JfQzxPow+/7faJcrDMZSmYhQMA
egG3AkE6lQmv+LDv3EY/Iy44AFmUUKa8/QKBEuQhJOfNpo4WPZeJGLsYt6H7QffnEexe6KyHfV+e
Sg2kaNQ4dyJyMZ9yNDVojV7nSHG5t/XOn2t71NNk20NAkjvAlRuwda4cBQaRiZ4tlr5TUWSwNdUO
tF68p2XhvYhfwidt99tiO6OuYQ8JvN+75vGWwC+Yk6EqgRneJXlXm0r+Mc6cbAkMaq8N0tyMFXnk
Arz+vN2xJnaNlS2eJFd+cuiZFZjSUbCqH65rpJ4b/oCu+Mo7LnXQm3uTtgQPI0TYkg4a6cB5IB+T
RGP+Z/jWQv+Fdv+no0vUlRsFVbE7cZJCq1BpY/Y13kpgJ0WjU4m12arJa6ec5ACA4YAtgXdtoO98
YaLsUtHuGjFLABd8d4BymNbCiVpBh777UnPMAq1KZGpozjC9MAkZe33lLV8QCdvYVXYtbmxkw11s
r75ZLSYT3ZIwRJ+AcmGq8Bbi87gvrP5Nfh6kLpiCOlAl0rKAdf+RX2HEEqlvfOO4Aub5zIYATrBL
4DtYZeWLbebn+fK/nTPbdLgBQR2rMyfmCAPPFx0V+eR+mTTeuqNcAZDLlgPtYgK1liDFuibbHCV0
7g5E6kIECo7yG8qxmgGSssSKPXRr3l8ZncfpxqiKuzpo0xumWZcBAXX/qzfwUu5Mxke762epSXYm
jhkL3etBfoPVloFqssMsZl2qkrnom58VQwntnBVjJrAVLyiJV6uhLBX7liuGZEaEiNyXZlbDRaPz
CYLtz3qlA8Ks0CVHxDi6DG03iKHAXReXdqkD8JfDwImBIfn1KGM3v+EMYrCzbPSHtb8kygjf1UzG
oeuPqz3p7sbGvcRFKIBle/S2/ByWQIUraC61K46pZlpp5ovz7nCXgfCi7wNg+Gf4+Y6Lv97iiY5G
JDqa2dytzlED8+G6En7+QkvxjI1fGlVfT6lnq/qPYoCa++/PHULf4gU6EKlsEEuj0bkjnHvwfj9a
e1G5VmC8jCVopx0IG09kbJYlCF5wy0FeHTbpGwPA3yGIHu/PZGKXPwN6RFCv8pvO34zVaush3vi6
gnb98y4fRTrhCUGjhwjKuxc0Q0G2chANIqg8W++lDA4VqGu+gvxYzr0MmHGqp70K1HXUm7IXuI0Y
5KwBKiRYEsJZrHL2blM5+/5AsqVOGuWt9UdEycYQtErCfoVIrenTmSIOVbmst/yLSEy4U8x7F0IC
o2aW9sFsWvkHxVj0y01PSdbGr8/W3A690J9WDwGqpELZR9ZD4akV2QZo+E+VG9Mxj78tPgcPTvbB
5BjxhqfPCsExHfvE2hI71FIHUz9LAGCnf/uM7rXkUkypYEpcUqVtjBhzox9hzmR3gQVzqwiJ5rWI
aXHohDshGufzRlRQhACfCAt95+LYi56fL9k4fbsyock0/+YRoYbNXXl8A8w3JKmRaYWOOnw90Ft/
V8XisBchtpGlU5pWi4SKihIT32WCqVw134F2VN7uIzFA2gtl3IOWum9MxNFFed4bamfVkR/zs+iU
KIYJY/iJ8kQg9UmosdQrDJP1ZubZ6ZELHVbC35KesR2RP/HQIeRFGj9n0GEcFdUBd3pzLt9B2DQT
RzbXxyb+dB3GhWw9LVmQhl9t8LihymFcfUUk+MXtKq5nkj1kNqabCUbdZjjzzT4Dp7PmCELFr+/H
l9SPwfLVA6L8SOD1UiWq0fumjNqYbWZJzTfel0FOQ+eTYNLqrBWybj3VeZe4KZCoOg/MR8CHa2fv
3Ex1AqreLrTr2QYI3BTMFZrq2zfo/Fr9d1H6O/bV447ueYaB+jSfsAzbmgk3ExwNkC/eNhS1mTbY
0VcmNmSfX25ApeycSmIoD/NIomAF1FPRAmf1jYPw+7gbJNnXlN7fU2PPcr6iEptX60Nzt6MhnKTa
YNAhuLeg9qHREzqJRBZi1G+HSr1eQLjNc2IdbtEj34KMrwl1hGXZ/W9ibv1wMbUjBZmEKzYi62k3
elbLMVNkW9WZIa8VPOtbafGkWgQF7/24SKQeQagu5Zl4gZo6ciTdv8+uvyWP5MD3rz6IHQDLXj07
a0W6RkQs5IJWbGQk7V9X9lJCk8J3aVC/elbywJHTMJd2B/CQVyMKGw2jsVVtAmqyqkapehJ4c5yB
KXQMQtn2yeEqwKN/U2THxf+YBXERsGmetSQaTEzfG4ZR0XQXAtClTU3kLB5AhKbbZto++mcNkhNF
XxqwIXjQi6S/G1ct3XPj8MGCeW3g41fl6MiqqhKIYjs+Wo6oFr3PGmVd/a09dpESFoAlhcwo2xJl
nznW0vKts8Z5Plwz9U9raDb2GACG8me5zgY7BhnUfurN7bAjAq2eju6wD525PVoeHUYtkZ8MyyQu
ltPLajXmCb6UWOl/uYOlzKSsnNIIShFVVnDI5RARG41UkMQAzQR4M6sqIlTnI6hNOIW2ozCPzuae
1lEl3chsqcWrVkb/hxeK8qeFH+gIpZqAXNi1JleSA2NY0Nl5Sq4cycWiKYu7bn4/z1F2oBr4dc/T
cK/RN8iCwCQcP+s6TiiLcY4HXj3vKxq3OrDtqmXYniIMj5Ipb799CdDE0O8O/wSoOlYg39QjC9hT
4YiFtxszSEOwQLnqIT18AWvw+sRjsWN76p/V1BAaOr/XK0oxAPZ6LFAVTXaaV6zWaNcX7G/9ira8
9TU7Pli12U3yAt8QkAyqODKlKt9d7k8lAmLvdG3Z21lQRMZnFa0ZZbX4oDNtUr9ackED75Ow+ZQJ
8HsQlXTySpDAvmQzWO6aYA2qjmyNDRFP8uiANjwZTAPWwzS/IbbU0IcspWcZlUq2RoAbcqzQEgIq
+Ojvf8P28vy0ou11v3JqtmtP38jmVqFkmhToK91Vc7VlENg3n0SeeJcgYDk5gkNT5KddGQmnWHNt
9hl//xGgB9TnPMVGpQ0AK5mFPPPc7HMxLWzJMm7/OsewqpiNz/7MYF2Allrp8q6Nu6k3Wg2lvVco
jkXeAcdjQ154iE6ZP5KU0bUmZF2QNSm2LqbyOPeTi2oXbMApch508TwLuU2meiqWk95N5Sk8Sdt0
PmPvZpy9PMiyljUhbYtL8hpx+dNo97RW1oifGCXSORYRrqqlUXYFvLIUJF5vDCo8n8y5j4oGhD/b
eOswQj25ckLzrpu7xjOIMNceFhrRDgTrgZHWMWktyMLrxze8k7NC2mOk5fE+3enhpomSIrF2UflR
vVlvY0PWxG51fR4zZQ91bKsCoouym3r5yCJibIuvI/777FJtew9anfNc/78zuazSC4QZBb8R192L
CIhvWzXejedM+LirjpQWI6Th/zbcWOJNLDvtJIW2/UF9j7elLNtdZ4t9XDiQjWeTvgbq/L59BjSL
KS9dDsj0ElK7b3XocmX1CdnxCzkzASB2OZPDB8/lEesb7n45/sYWmBmLTz3QD8ZgJ1RLxRNMBXV1
NSt9Z+h1Bn9CneuZi+z7kf3CY9+tHTihWGWt5eUAIPiMCRz32RSXaqxQJ3ANF2dF3jEuvet8xN4g
VBaxfKdp1vF3JC8vIliU9Xb2Sl/Xuiu0aeAWQfnxtAmU6Qq14SedhgqSBDnMppV9b0EATAgBKv8J
BCgAeKOA1S6ucuOx+RPGXvm8S1SQXspMv2VdNTgOI/rgOnoCiuQuxq/sTK3RZs3Z4TkQGMRrE+9i
dk2e1u6D4JTu4t+4ABQv2qacbsfa9lrPnUtWEWNJDBXLfW6/fBcZuqTnErvxYk+ZGGUgf/UcwZ+A
zXZehfv6G5LprIzu+RrxFZi1frys/abWPSjRK/GTICp1w3ZdVQLvM1mb7bJ1qFEwRBaiRzP0pObQ
kI1tTqDkVc5YJE9QehbiPKUW36Wk3YlRmUNeWLDqNYlHDU6pjFsbrrM9bJ0nbFmsoE8dC7cs1bjH
eKF+j7auQf0PPnD17bjtQ1SrhBL8/+zvwF4225ZoB8bfg8ArVTY8fm6yhWGGQKEHwb5gbZ7Z4N98
ihzlSF1bIA4x8E62tHCBa3kaLqlF/4hxaS4EM0lMHFS8ktPZXYIZQbYxftmGjTB1QsIUUKigVRj+
HGADDhpy4iWE37zmwZczwd5OSjX2ET24V5cu6xnZBC8CUNi3/VghW2MvtC6Dx45fFWrspsqKHOQP
1oLH22J6O4BScoGvQ3Bn8ghNLtO/CGux4wEpFKAy9UdFL6SedjzaKF4PAzUYDwARr4FhZwEUThw0
ZQuB26s44CVXxTiMnvtAwacxjZereeIlJcTD/ieDO2PfyNDjquQ/z5btZeIgp3/nDiGvgMSiNuXF
pzW+ZuaUb4xv6eM83xr/FH1ssnOnLxR8h1mJhmky0M/itJCWOwEpLCEKZADUFDDmwlm3rm0EtG5D
Etj84cQwfRrkw5I/Enjli/W2wxw44HRK391Avazdvw73cie8gBmUsdWn9A0XOJGKWSi5ZzKRRrHv
hRvq4VbzUzTIbRGD0/iG0lPFHCTHMybMGDMyyGNcip/TZApHd8SswdGdfVR4/3/cgQf/KuL4DwOa
TetKsx+dyj7CrIzkPnXua/5Pz09uzX+lF0G8SYtA5UxNlEZNBsFUTcCH30zWllP69mIkUs+lkigU
PQBc6dFZ1LjiJ59UGm/t/B/1ahCuFtsmyWUEuMJQJH+4mHEcPLvtMjX3qXprD+1DNWmM3TIx6Xsk
hXhtmWGDdnDyd/b/qD5pNMYxcz7xijNLlVnK6BRHl+nonWd+CPSojtbdknPIm247ch1g8Iupf6Bm
uaqSCKTsJA/m+4sHWVNq3Dem0il/kyEp/5wsDkAa8Es6LDYRhRNJniH4ECjcLBtVGeQKh5TUAZ3P
LDrn7jBOsHYPX7J2ywgym5ZZCk6hue3u64SxeebdWdXEikYrZ4XV0NOAM5sXtY2zMrbIoYLgE0+9
aC8ba4VJJ5tIuSgwvKy4ys25KR96JA6OPG6eqI0E6D55RwboTIrYLutK5Bx80nP+aL1t+sb0TGRa
prHQrw30gERlAhcCfu2boPqHUqt65K66DlGk1anIRwuMmzF/2o0bpdlqruA4es/V8bkBg59sAyR6
FLaKShcvJPacd0oFDrbJCVuV0ng+wf6Ts/COZZGFuNOytWoS2LDwfOMkXMaLeIBnAYrfDEO7uS2j
Bhesed01VPEuzI8I8ZYk1sA80JK4aEf4d5En43RP2mNS1/ldJuH0z1aiyj0u9w/hgfxz5MNw0spa
+VL9caY9+Jcn9OmIqmexXUOchYE15NWtPc9D+PWLnbiTNEXwlKoIC8b3jYz8O5YYji0/1xjRdzrU
+0YaDsA5ubO79EJPfbzyzVHJLBREmk3Mz9rb8txccAhIDnGReR4LB9p6J8zhuvK0p4a3B1W15Ypd
UWGIFtPCH4D4h1UxEw7nhYK0W2Kvhkb/Ug+5sqaS7ckDyV70XSlL2BKtQ041HhnpepB7YLguLNmd
pSRCpS4qPtOmXqIxa4Qc5LWKn39TtRHLJT6irs5IrLvf7X5RTV6ow6zb2dIHD1lWidFW9bkVdUA5
/4/nOw24NEOM9L4xwyH65rHF+ylVUwn6XCZP4EjagZogxNS29O/gpOteZz1jljCHZTZRt5POGZMJ
gUAvLRRUdMg1wZwYXxeCfTp/y3/t9Yuf8SZwrzv6pHdO4BmVBKsYiMHzsH/QC7Dgc6HIFcECPZrK
VrlzslMY4UbUaqMm69ESEgfF6UB8ZIw1O3OzyXrl4C5hESjJG5OyeaHK3myksaaHL7Im6KFTzsCp
AWWyWMufk1aXshYrB2ZXa0YOFNcWpYmokF86GxFahz48kYAEZV5++wQfIH2nx1pYHnFdrJenTcjD
LZ7szCG4YN5OclCzE9XJRHGiEvBDBgnkNUEJNxYGNwDIX354ep2ww+L1g3M9/yS1GTS8sIdMC24b
nlpeuBltZbLwdCHO/mRebGRGMrnEPg0T60Wo6UtdiVX91SgPEvB7u0LC4iPJSF1RzVkitjZgX6OO
ZM7cEzIWH//Lq7rgsVb+BnqgyuFNpYMWKl5Gw+W33eLPEsPshBfHq/uEh1vqWGzQHjU8csxNplR5
AfNSDQMRWYk2SeNHNLiljIPiApUFbQgm5UoI451cpDycBBPtBowsYnYgV0t6CD277SVMLIge3CZL
Q8ITtKQHICty/csePHN0pYoX7NRGGaDhpYuCuFGn8FSM6oC6lslLZ3KOhCqfueAx+USjVo9yRjz8
M55d114AuSYgqDGKoHcwl0NFIVPo7Os+SCyt0t2U6W9d5htlawDS/1z3C0ywpgSVNgaOMPxgbTAJ
80ecbLRIUkaIfUxY7Z7/z051UUmQravsXUYgiGGQeSySY6g6uqs9JN0Xx9YzhJxJnL6OZv6qnyCN
tvXs5JvvXJdX5RENrJs2EADVfWVw+ISW3QU8QbKfTJdzRBCvInx3keBFeAye+L2VkmGYGvwhDJG4
ftYcZW9VrYJE19TUi9Bh6XZSXt529+NhaDyFsa9yD2y+UVo6O9NnLLGDWOo7QZEw6KXlCQD2KAdq
rpClZ1id8X4SidFVVzi424rq8+9SEsQbmGBhJkcarHk1J4LsTEigyEhh8eLO2ymG7U3nOYrI+P0w
n0gvvKizU5msfEoLbaXgoGoLy+d/LELtlYZmn/l3pJ8vBhpVCTbAw4wM6hdmFQY0LeVJkHJmFxRX
dmKBclw4mleJtb7GM3qDzzVk95dCDP6M7y0fO0p0z3EijOK9pDNOcD/k6gsfrC+fZ5AMJVgk12Ri
teISEYmXgQ/J/q0rUCQlnf/TI4CtEoF/taAiNDOPiXNkT06tsWqDUm2NdVb7fHSAmmx2lXKIFkFA
jiuwHx2TBrO+kWpBq1KCB+0CMJzb6sOU6VEKvo0y7ZeJMuGYmxugNuMbYI71thgZulpUusvOgAdr
+JvClVK86ggC4c2qnvib3D3VQUCRAnj5iljGXbDZ6n9CxYxcygFGi4/aBIEEWH4xpMI7sFZ/xhEn
OCK7BKHDwca4gWYMvDvv7KBp36+ilGe4b70RiL2uaH4UyPTxSk+af8qYexKyJbu7R1Uiguuq8SXk
WFuLhWEWFQxEeEQIh2/9JWxPz3XQ8KF92JnoeZI3gL61fr74+sFarlNPETOvbU45XsEp60C1Tx2v
zsSQRyqrQCzQHicQ2bpmHfwOPkZ2UI2s/L4UiHyGgJPMWU1ECYmTNU/VxQ0FAzrIdRTGtCPUUE56
dHOEKxAVhnqnmBvSC3KqJ6ELDHP1oaiZUadlam+mxCwPOtyYxrO+uo7QyffHxJGSYNnum0ogEs9X
Xso67qjDL019C31E6mvMCeT0aVqfvuO6yc5DseUGA+mdYMw9khhyvzMGxddHNWniU61flnP+elLK
6ouE3PHTU9avx6FdNFDNHCqaPrlKlxsZbkKtBMOKyQ28HCL2VZX9vGO/ayv4aozf5QQzz47CJNZ4
sqEAxLTFTe2o3mFPkK1scRMJpBBMSP8+PgmzWI927J3pk/tiU6V2TXmWfmGosrSRUSNsop5pvDKr
86bVZdAk+1E+E1GjdAjqgA+A+ZmdAfGKAvyg+IX31HGlfwYEPx5Dsd4SPokAl3pTyT7CvammXrfU
kioQcwLrwIYW7fNzag67bfw0okRSJC427GvLYmW8fhTPxaAHxVPGPg3rJZ5gESHFseRK0RwbD0w5
UXYaX5KFsZl+jRn//9JdzDABcOmoSzww/yH6Dy0/Y6UDQrsjo1feYcsSqAijgEYGdlJ+PZz9Ji6l
6thukqQJh/JHXN+RHWhzb1QySkCOBoyhCBwvADJKjJo8HKVXQYrNf5aXy1RTWgjz2CTpOwGAQq4b
Hz+MezGvjyLfpMQ4oqDksjksu0Wlvd3LfnhgC2LnQWM1i/mLmu1XtQdM2P1zKJhfKh/e16xx87nj
FP2+xAdUEIArEMyPL1dEiJ+KtwivWyHhqIBzRojZxfESwGaZ6qfPpFdRg/vXf93+eqQEqrf7FjfH
aQVc+sIyYVUhR4gYiTg82/I7CPFAWQwPkDTZxzm1i7gG/7WftmglPz6S9YESny407KtAW1XjIBSq
opztvLfC/QjcWClqMG4tMIR4120SsMfCt1Wv1maw+rVY4h3BRU/Az/KsC5dRKQBI+o0wThl/vhGi
ehPlgVcbA964d5ZS77m7FIVT993qGEkSulINIU9oZo583jhE6AfIs+kxGibkPNTNGapHCQ/NpnJQ
Vec963mjiuHlp1VE7yisQnXOpERzHL/7VMBC/LMvW9KLXMqicsXzw9Yx1O6QZ/+RN4Qm21bBD3ct
UPfsZyqAGBZCNDic0eillxnuI0RcAWLS/nOvMHVS3/QiRGxXLdgKGSHG41HiZU9wbWg8Ww+iVI64
dfxvWdmzLiZkMCAUDhbVcxVxDKKVRDuO6t0cZjx9NZm+cd4eIKr8zPW/3igOK0Nbk/C5ACu8qln6
KHFEhqxRF4AXb/Ka+T2SN+o0k8s/F2HjtFXoGu2+gwZmlEeR8AtsfjL1A6QCc3ELl/VV6CJMAr0t
lDbYbdZxt2OSliNBoc/mQTTVEed+uZ6ZX2AkxK9TRM3fDQzR8BDfZMAAbeWNKFBlhl7aPNdi5+eE
SGCGYaGVTfLtYIyhm81v5BwQkdqU4YbneKfsVA/HbuAmiSjD4JnFQJe9jOEL5C+DaOdMLL6xwlwT
NUf1zllDRkLscKFTNHiIclM68DpTxs4aASmXzeM6wSr2xLDOA2marQRpQW1tHf1doJOPEKNwLgC4
cRTi/xAYaC/sR0Ft/1U9E3XHeFkO8bhsnpxYYBHZ5F58bynGexiBjyIp/SeQ66nqMhNv2REcIWQc
hgYWFWCZuxVQ00VEU763eskeDpcyprWtJBIxj68imm+0O4KAqknnlZP6pGBSWk9wnwDSdpHMSp6u
QGFj1SOjVfiOETdkZR8k7Y4rFl8JpVoVaPZ0qLBya/s7O79a9yt54rtxvEe51/NwEijXAf6YcReU
RGJCb2d/KEFE96Qj8NMrBnusnZwOOIOK+JxryDgAIwfglBDWoURJlL07bQsKCOojc0udDZahHLKk
QjOjs8ikCpKSBnFcjrlhzw/TTicI6ru5l538UKdVSGQatvTI2jo1HHw1Cj1ORli2y/2OXdfO5bkj
9ezsd98ajWqZRn9TISZy0ZQOb/yV3p3gxPxH1NV4yhEx+hy5bQMbCiGG80wNLH+52umGiSNqAI50
vPbtXRxZGYcFw9F25OYpeE2RoH4aQ0efLaRXriGYn1EdEzi260eXY7qYA8/XDZJh5uzyKEBQdUoN
lGfvKWy6IyEgYmDddT36rCkw6zTcJEdvdsaDY59Ehc/bTBimyC5h3QjdRuHnlKrahaM+oc1wJnMw
3o/R2HrzCHLZir0Hv10cz7MmMh2Cz8kQXY/IdznXY5Mcde4nTgDzEmH05K+BMbTzMHmohZtDoHPM
5Bo3SomTAsn+QX4U/Co0Tmd0nMQpkQ8zYPQHBLdU0AXRkqCHqbnhMieroiX4hnPvI0IeqKIpPvJp
/HRMm4EvEGPEHmHxYzirIBrqrCHsSd//pDT89EL4v/t+DkoG02MmW1Lqd6mZoyuKd6r8r0VnKjFn
1jIADYINSQDlz6F0nr+vGubL+ktP0vnIamd7O84ziFevlfhsVh5u/FEhweqf+C5MjzhbS7Yzp24u
3kNkFrj58cdMlEqYgYR/jSME1uXYAoD6Dtu49fXh63IcA2ipMiH17m5RjWRUokBTXYUPhkLH5AxJ
Icstyjyf4KiO1TXQVPlTtdg0W0QBdv2+AxWHmR2i+2NtYSnc+PTm0Gq2eQxDU+BJKGjQHXoC9wQk
v+6aor2BBpgP2VRAyYSQo4qmZXVhq66w3UqvrPAGd23St6AbWtMgy3ov6W86xe8UedrPnv/feuZ6
IOiFHEb2BKOkL5DXyrCBxPh8Bvf3cBF2Vd9NEXuepyB9OazU0SfQIwEhc9vbeu3KwUsMXcAl0Yxx
KD9NR8xOmvMj0uEZ5Yj2UWsGnn3KuE9s+tNnG2ZmuGggoKBlvuhMa0wnWe3uSwlUxToF+dwv9JSl
Y8QKf18WvgiU+oO1FKtHC0UloOKqpFTBDKoQYSTvISKTz4UT6N27LdTvKNdNnq/MWKknVH6qpBzs
8hskUTw0qZg+y+OnoptaxiKnWe7C69HzJZR/yL/bYjUzT9ylJlmCFOVHx6S78xzzuxz2nT9No5rc
dZHGworW48cYjc5Y8a/nwVjKIlz1yF7mPWrsPZdUtB1tqZtu0akZaVLXYoMaHZlaq4pzjj4/MSSX
mJiSlt8KZ5AyQb6H9fU7mwg0aZog1djgCiFTNjzixpZ8Gil4hVbpwvkO43JSWW+9C4I+fU+aBBiM
I9FU59CZAO+dadNh5G0KpPo5zjiW+gFXRXe5dbr0AV53H/E9RiC9YhEhSN8++qTI055ckYgekqEG
VYugpQlWavr3a3GfWlhXryLiVRBLAHBP8Kd5LkJIAH7tQ8vhPM9svzOQSviYDN9Voi/NYbaNygUB
yfA/wYsRUNOPYBaY/0pVxax2j1NfozZPpjwDIcaPbc87on2TlFhsn+ReAKRrMs99QAKXs8slZE9z
n35NJwY7FYbQSQR2rVPRT/dsIvrpBWoakaCJS7Og3xdCBk57vtbJIALJGHHVyaFuYSOHhcu5yKsr
bH2g0OpS+PKNPlMBd2hrpIapDcID/ld4rUytjxz5Yx3Kf6On7ERRw8ki4/BUKwi6Hmme/9Qj4IbR
mZo1qfP5pMk7X/dxDz/ST/hYmdwXTVYg2ko/8itxz2qb43NJ3grUtngolHWYpxnVqYOFCug41GgY
aeDBxJc/7XVxEOe4f2aaKfwADxIF89fT/MxFP7u0QasetXlZpQ866d61dKhp7/+HDzWl1Av6tL7l
/qag7uprgyWE8mPmuETUMFj/5zCGHF5TRkcU6687zhg+K/SOPfAEdwSc2uHKvuEJNs1pQSLEyzFx
CgevT383uiIOuWNWDsVSZgApe5b/x364Eboqy01ypm4W2E4OqD5/cVSpdb9xaFkV+31ztXFEdvYx
MVLyuRc3p1PeaZN3sV9TuWDn2FFMicFRMQ4W3a9sBsqZSkmaHW8enkDQU6RO2chA4ptwQw9I4MHm
Ml+aiqNdlxt3ifn7gy8D+Tqicu2Ilhqd7Uk6CFB0SCDv1JflHPAmXyGXg17Hw/Py6QOxp+6/u1yd
8QQYKcpYCsXXQ+cQKWy634oHdHaDlbCrtViPSBTy/+7j+y9ELPawhHd/nSQ/WdcRVT5VuOb7IXuQ
3ey+caYJJiJQyS3QMK1Aif9l2ofUJLlkjknHY/CZvnz8IyGMPxQgcIdBu+2oEiWr+877VnXLoM6P
0UBwO1RUQMlg/9Kwr/dHk8/14XMUQyCRnTGY0xDqogjvOAUdhq/SxHTvPncjJMp6JO0zND7ccpfd
U6j162NweYWIGDpSbQozYHqGPKDvLwrYIP8lOyBdOe8u+jZuuZnkqd9edZAgmVk1BngsL5Mq/LSU
vDCe6M+Dlvlekl/f5+eBkJ6q8Rs8L07BWz26VXPJhnPyHuUf9jSHUfCw2NAHczcvUcr1DsXRv3ka
USsS7pzFjwKSiGo0T2BCKehuqQoQgu7OqysBaJ6tEeiatrhquzYVXBCbyx/9xJuNp+tYW1auhTsN
eF3HelERK6lAnh/WXJl/SEnfI9iRY1/XBPOJgARTYLbbq+MsBbJzBah0akh94zl8vNXCw2gDfUWy
QHTv/Xfqms6AgIB0uwGdMP1X+LMKZV0MLkjCH1Y0v9xr02xB7de6Lm18MHR1ZJZNgQZz4RN55S4e
Jl1nPwmSuIsIWDpVCwPWIQnTG+xpJWDOZC5M56HRdfd3yn/uCNrFcWzjTgPVFp9goELE/4bpfo44
BfsDJ4klVCa3MGOZeXoyRbcO5VQ6PThxdLaI6Ifh7Z1wQCGIQ7srWBkUw2XLuvGibhGBPfOxfZ3T
2hPTym/ns4behBjvliM40CPL+RkEYI4cOOuOGWNOcaIiPNBlDD0ofd/+zVaOUstEMa3CIaZSjpCd
n6+tHluvd8muPck2BT8gHV5J79lmAwowLwwTlcoqnVBlmGl9Z5owiINZSMih3jUg6hTIH2Gbx92u
5kpaeichxm9mdYEKGreVGZd0nSKFRfmetUZ1I/aepqUdVa5VQOGwatvTJtA6A6KbeRJGNN5Rye68
CrKGa0qY8RR/sMx2zQtX3EKdhxxN+hGF5t+LP+Pg0a2eIHJrAescgjwFIVU9mBoJA1LzdqFWiiC8
UfN0wfD/obmfbDy+LSjPlkMt5uRkJWCWEmmxeljX18fXFIFq+O5PYp7zmrr6cMIp4zsGNHtl+JBU
z32iaEzPl5rnJwY8EAC9isiqMASRo2mo8I9zwpR52tK3k3E+3TysnpOvFT5JfQXfQu4fX1Sv+zPe
p8ygLGhBRNIg9z4RvohFK4m1UdN31kNTF4JQr7gbYbKrlOOD0FCRFcMVuxORqFf9MMRrFQ5Ztovh
J3DzZx1/2FsQJlViD2YIIEjShYdgOkPRFOB2RwRAPqHWYDT6bIU64XeqTPNKe3SQhy9wTD1uRzYD
hcmjt4wLwVzGW9AXqlI4sq6sQ8+5GaYaBOVhkQu+DDq5CVU8BoZ8EtrvmgSXS0Hi96cGEjHfN57X
ooaegnbB76VCTT9cnv0kkRHGMeAIpUFDH2Lb1Fionhu0Ie8JYOXwKi32YpT1HT2RvMAkOFURZufp
3ym/DWAfZiILy123yLHcnCpgototJhHUViwUTeJes3/kN6EL8o+7njFtpdcmTkQ4OfKrNkM4pnAf
WaHTXvk0BJxaEWmvJ0TSYE9lIp002MpIQT9Xjm7L2iFGWWxBrMNGOVMGbvMCn2i/5RXes1W80wBa
5sHPGjnA2EHxeKKU4vt5YWkpCx9L/Z4jRtG7hkHhkXEAhoOu6mxB1fvNeJLusucDTyQmqmBRmrWm
wrNn0d4GH+7RwIAqJM0IGZDp4EG3YZJVUBffgnLkbIKAC4wIwn99lniJPMsOHo5zcY/oGC06/PCI
aBl0WJggJVMb6rgPcdu0DeGI44ZUTryvTGvXlxy45R/K3QX9Bqm3Jd/dFqhSFi0KGU7FAoXigN8g
XSvdZ+i26PY0bvkYUy1VlsnT9SkoHBj3e9NekQK3nItNTbBBZSAjIoCVswoCo6Kbu5zY+Ox/zGq9
606tpmvWnGJOcBw58JTLXz3R9fzTLrctDyFqFwvNb7o06QtBWr8zChYLx8wyJsPL8NTjS29c7tB9
A4YQAQeQvFbTNpneJqW0YUNz4F0utK0Hp0p/kCUUMZeU0S0yqu0NjtedI85AsSqiRS6yzPoN8r5v
20MjGJOS+cbhp2DY3TMjl8EdIduz5CJr62fQv6XCodFtuJux8UmCCEqL/Xncw6x3y1Sow7mTZzZ2
Lecw8LcxB3OJ+az/kUG/TxFBT2kuEN3Vgp5UQzsklORxqNCOCv4RvEWGApzvjqYljVwZbRtJa97B
BwsbbJ4l7L6es8aKTBK6KHuUEKCtcPLTTy22D00B1PLopUqbIxpgBSS/HRoD8Ur0qGiJGNFrzLlg
g4NmkfH0stqlxxL4erIfqkXuKwRTSivMBHG4li6ikV+liIudpz2eKP8iHQNZunb2+ekFLKkFHCwO
dYf2iYwdUSHMmY3DKKD+zjsjrObRWUDnTMUPHv1xuJz1JhLBZlpxQtd5dgEiFKRglwvL96EocK+e
cYek7vRZdl8AgQSDzA2O3AuRWym7UL7wfp5YemVdEWkMX8HKxFxCXC9r9qK7dpI5cJpMIfIME4hX
VOcmK1cWCBeV/BB19doJteKNinMU5MdNT1xN0ifkLlA11HTTGgccEx2xgA91cdmuG16qIQBrRuXC
gnFbdpYJ8DksuoBExwFrlPFummphIt0TzanOvD1BMa1/rkOWaryWt3xf6g9eQBfbd/DeYCkI75L7
9AlUMCrhdvFFyF/6GAxCD/n9AuV+/JkvMlpe0rFTTYjolEkKuoB7bPaLbUSovMVIxchKKsYc8bZh
OcX5SfxCWqRtGwdPLs8FrjlP4IlSsTbiFoiQ3T8nkMgBY/9UxTmsRjoWapERzDe0oOexOOI7tz9w
nrPEzSWooF0TZbBkBSBpkC3KVHe5ggvHDLImmiViVTVxWQFBU54Wg4lnMRv495trstaw82SMfgv8
/MdH2yfvb8uIvAkp/+k4kQ9wk4izmhbWjwgRYfefaxmitT8IOZO3L2pQbvgyFjwaJt7IfWl1qRGT
zF0WgB4+8B6rqfAuTtNEGhcOm7x0/pMogJc5uhxqaQ5NbrOCMPLogoWsgLrZm7qGkoEWAOxj6e9h
9OkNeEv/K0nl8vbt1PkLwxt36YIr9QYpRywwu/bA1b5EmRHgpOetteA1nJQNaoNk6p+GNTGe3xOH
3CA956xt81oB9F74tbnbl8TUdTsWjsN63ZVgmA1E7imTkTndj931acDdUM5HiKiZHY0ZLv4GrAXL
IReiAZ4o8O0AsixAJtYb1zmT8HHl8rsN0NrjCqOi+YxI70PMRJS/30w4tIvXAXC4haJHEoj+jtyq
rlnIgVsaFbsvz8Ml4V0UOuz1J9k+AvYmoSrKuEUFcDfgmurfCHCDIfWvn37Io9rb04Oyzh+tZE8Z
STseoMs7/20xmP357mfrFQJDIaalAcXc1kwDNynBHV+W09FsSby7v8uWSJeGDy/ry2Q8YzeG2BNi
JKRWlWsd+p8J6k8Re00Y4XGdHhTFPO7DtcydYT3LgOUXho3ydMniQq+pZ+lOY/tbP2yqKIovLxWs
qhqvuqNt+Mi2/xgBYKYNRsv1OIwsbfqcD5n9DmtvMSFQ43rPGRDxM9ly3lvL5DVqpUhMMFf36Cr0
yHEoHLjGCRdiaKx9y1lcpwp9xhHWvQ5zd0OfPX6hYogSSwLDjk3sXVk9XHRRGVcsKBTGryNkVPKn
fl/o7qsJXxZM2MIAYjQQCGxPlwBDNL1UW2wl9n7ieTOWBWOtzJOmZ0rd7MgSQ+jdDjKbXGcHEu4r
07TUyTh88FlfYxGP+FRlco5mg5ETY1AkIgPJDBqcZSBe7al1AeD3yHKbPt2ZMsubF5VOGLfdjA3c
d8m/P+4gtTmXQfUZclBIb2x02b1y7LkdI2QlZwegxiJzLE7dSa/0ZtC2YPKz/iyWjJTp6H9VuChP
Iek9ZNpdBzP76i4wtpTbWeaRmqNkkB9gmJstwVNxAljFgNqA1HgQTl6uP/s52JGpKhBgdQTmVIpN
O2SsZacURG0xp7DiZcFUs7WnwrQYRqfS1arOV1pOkxuR+XDj4A/fSmDf00+UsBrfOauqZrTKsAt1
24CX6N5QWiCUF8xUIhPMGHwDMniVMNYIlf5F/iGSpgsncz+n0Aqr5aktcLlXtwEMel3JYlX0kpzW
f0BF2WJn2V9wvdrR2xJjc5yYdkpcl4RGdpkO0pn2kSFHT8euMgVmiqmDck40hjusVnpfWU8eLXLZ
b+4ptW0SrYr1rlkJ3DI09lLh0q2L90UZdcEU0D/QQpeNlFnElW65jbLl+KCguEZGNO6LsyW0AKBV
Yf2Rf3E/84/RFEmUV8xFz50ZpEKeiyw8UuKq4bqTO5n3Q23Z+lubU0T2I0w4nJzhSs6Rkv7G987c
2JQaH3NanO/qaQukiHoQjFfAQb7S50fM7ZvXXnrZkobfbqZx34j0KP1cYDoV3RcV/tCLY3vxqgWP
hIiC9IiYAYaHI/0w4NJ/fKZ2t+sbSl9D8cc1ZNOPmpQREkJ3oGc0ZLpFsUpntJbBo143e1cJOyDd
JMKvsjQ3uRuECKOcxsFeyDV1hmK0NsqEhlLE5KVw/gPIhApejq/q43arR8r2YvaYYtScVUml8mtx
rzflkxLhFV2SANt66gSo/2iNbx2zWt8pQ396pWI2FC3956KvIZsANXDDRi0H67wd/oqXu6aG4ppZ
NyHOCUcwu+XkCrITRIBWZhAgq5QTyfYyld4UTRweu11heR47X41CJlfn5mlzeLfzSPT/P9/+cXw8
mMTD75XIb9KdfswTwTgWnVOuQrKg/eK6u49Xdxgk3ZpDAyOMffie+a0h1P2NygPwFu0/BLB4baBV
2Xg0E4tXsvBenVA2OdPJz6h0aoj3AukaRPFkm7t2D19oyvdYdxKmwet7is1d4jJtxMxElV1wVtj7
i9G30fIbmjFNP17pV45/k9yGqsDvOQQuBWxs/WnIVLI2zS2vbl9amrxUXXpDkTj7PncnMo332NLC
98DBRad91sT3mM+6m37GFM5L19nXfmVHYTeADITr8JlTFt8hDeHIVHh+7IKHw6iaaHnvLnYi7AJy
dMVzKp/P12DUKSXva4N3BYkLDOWBzmIMwg+QAmAv51LlOcNUtyCBiVIFRuxNSNSi5hFppuONqA4i
CWn9WhbfkeiImO3iRtyv74eGfbOBJJ5Il0k67naaoKeKIoFTG+xAE16wtGZFUZTkAHfOxrQCtPTM
PgSWTgoij0MWd7PkYJGBest4vdBJid5xdSYPo6PiS/+1RAka6Q3JhKDJJy+trS2gg9zEb5Cjl8XW
T1uT4wx6CKmDgJ4V06Jpiayw5MJjxeCUOUdeKHJHF3idvMaWyOK4Xy53DQbmTHHBLpjxM12SdR3v
FaToojQD6GRNgHTNqfvolbYzQz3ahU4CZKxCgzcWPJntCdWjJmTsOEK+1QVAyOSXzPtcb14KvlkN
ZiZ/5UISNJm5ZaOfW5KsauFo7eyArHPxQLmD3TxT8P3S4YBoxRFndHKz8Ihgcm/JvAvlicM1G5a8
H9AF10NaOF68m4nTW4eM/DI1VVvmaFYNIlIFxm+SeBHD+9hVW4wXEfBFStFVAGvi9z+w03YX09i1
Deqnq+kv6KRZtktKWWTOtafrtyXsJBu2hRe7LTrNnaUKybwOuo6OBGOtimH4gLKAFCq/a7rgKAuX
LozCnv/+MO7YOwpl9JdCxhlfMaMLd/QAGe8385V4hzcb1lVlwNuWhbJnVh1ItlJG7dHzoNp9Og08
qV9HtgcKFc4RWI6utEEwXdzrwLFBmAg0B3wMjKC8J8S7oMTA+nr5w2QZvOU2xmAZVjz9x1jFp2UT
LU++BRJCSWIclCFo8cDGrsR8RrcCYWyV3WHlSUAi19aqlkkDiAhb/Xl5go4OMp2eTPlB8vWUkLps
3a0iv1ON/+P3ILkWwzf8eJi4jBQ4cBTCMulf8Wcg8RUci6VZRspU/D94EVeMW7qKYDpDaC8GEzee
ycOyV4uwXF3aIfPMfEYfbrm8PYt6LRKwsZELh5FDQdM/d2vS/kqnv0XtjgwAs3VOfVi9OMKv7MRo
RpyTjH+NxmRSSkJGtuvKEW8ugY6UISQSgbuyUNYSE5gcCw0AkP0nToo5nND7Vh0KBH3+toQBzgp5
l+/g4HiCLrA9KMMCpryyeMm70ApEQKTZzH+FGrgZIszuhhe6v/KSUby5dAtmBd6TotP9O+CvJzph
PGG+5NsreC69mg4vXPfjp9FCKYYdk2eUgDYJXE/NoB6cXJtKG7n1jZx0uXP5xz1m1A0zZvIc5R4j
hIdZSboW+yc2Rm30uhCy9gWQ1e+VPoHo3uBRe71VvJN/LJutx26xs54Gxa8Lq4zsuYs8VHt0SC4a
WXREGiGuqtY42z7NTo6AVlWtJ5eQQoM1yHE2nIRlTp094EtFdDc+JAs1QAcUddIvXDN7WQ5dMJaD
8+ssj1fYJ3ZN3hsbQFJ+IX8BcvMm1YY74ZFQWtd0a+AZ/joY6H7Of7Q1BMl59pXi0OyTLE1QTaZ+
PUgbsMBfWghoOTZ8XhYrrDcMVlKqiZyAfuCcYYS2vegib48EkurCdfjqOR8Zq4wakRNMTyzkOFYB
m11oWrAuFQkpk2MOLGJypzY5QIr35g8g9+vRzgLS3WftRpy9lwQPZEigBwSVa7KbKOFFEhwdPZ4e
XFGw98hnBVzzRh0yuag+nQ3YGSKezcIlwhH6NG05Vz7U0HBnLOEhdqpXqWWc8RN7MJxYrewhckDy
5NPKSz/5OGNf5XwBSSTlkrhqf/AXvR1sBiHc2O7dAMtRzY40DmmS/r46P32N+eM4KRbaSu8X5dt7
f3joxNFtww+tSc+VuFOXfFI9ktRR+rQUP/0SGnyVX5jJuh28I6wJTG/t+DTXqYq2NkWMVi4Nqnv3
K6JTTACMAtR4ODBLHkFFvFMnFsvHvhiEfOp0nupgsjglDrtkD3jNEYIpzOcjvshW3GrY6w8kX1b7
4AOBdKYQpGlV4lAaaNBMNP4XmWN2WQZ/nQPLA2VcmeW0hheguel1xHfUcnZg9CI68cisikHPEp+H
A6n76RD81ZZi1WhsA9xc4Y9PzsYbYmwAf9/wLtPCv1IYXsTWSJLcXLIgCYEsOY/YNUNu2BeTznV9
4tw+O6dWyVdH8PiuWaYd5NtV+xWnGgAlebrqDVWBZBTGb4VfSs+ln8eO1DQHwGGH3NGmzqP+nOhm
i8zYt5QlDjK815DvQVGsn0eifXV9jlHz+2iZ5XqSP0mTz2KtSb2LGSeCmnGII/94YRL3DR3CpIph
ZYDrU8madnxEtT4gbV8zVseJxV7O0TzvY6SKMsbQoFZpPMbtkYOW8tEidM2MWUBAjRubbZVQWsFx
henr0vYDCVc+RHTFAuyjBay5lQ9V9rnXS8TPiuZ6c8KxJL3wlNhEvH+an7OkxP+0UFRkxaJgHFzf
VmqSYA6nFLtKd+D5u6YNViFLXpsdKy7WHQOgxGa+LG6ZkJ7VgkCuYayd5ryEQkxddzzwqHvRp1Ws
BUTSG5o69vSHUloy0MKg2jblIhjcBIupCc0DkRClkHaKm0i9VGyJuXxKc2ctCwbKvI5u+IaKWsPK
khdJQLND5KYNdx7jvWrrIYxzBVHpWuPX8RawrD1yZGCfpm130rEXca4Od7zIOGqJnqOqDhGxyc3e
HIako8yC7kB2KzmR83FGH0iBZKvCe8OSVoIVh7O5gTYBgfCYNuhzA1WSQueyMJg9U6/aLiVEBJoa
3nbl4xa/hsRxJfL8o/ieZznVZrtp2PReyfQ0x6tfHo3AND/AdLGmlUekz+9PFfdmt9xLxB0WjhTS
j4iOVskOcjRPeaX4llouk7W37lIaA3GrlmGZRlN87VogF7DEaqV0B1FNfi58laHaUheo9k0gayrh
7cqJKSLO4c4pOGLBajjfVPTYl3crPSGM/Xm1TAmdYCn/K8Qj0nQGzGpqei9psLXrBZBrrB8ikdeY
lL6+EjVBZXZv2jihosd2eov0T/jV1RrqsxiZydEwJaIuj+Bx3jwSrD2AulL1C/vOAq7hvea7Kosl
w4szi+45hoZZ7la28kyPW/8xr32QcSuroFbd5bbxGsrbB4MZd84mpQ31qFqTGNyZmgsiunkhBCDX
vSaPAvgE/xnGIF9deX5QEQG3Q0x/Wl0YNqduk3C/MzRc36/KgG5R4yVG/Voyx5VNNuB/ntWe4zg2
f7KjRlzJeQE94mO8+RqxCZM63vHJyznMdTRrbcRFxzEKjYoy2Ek1E+TG26iptkHTg9FrWfdDyTxx
t02AVTFRoKiZD4gbs5O6f6bMf+dV2qlH1wcSi/WMaemxVYl+IUXa2LSf7Tq3PMA6RPs4qDn47Ylv
7XJXT3jR5dD8IJNBI54PlxhW+a6TEF272eVfTs9fzdMXFbAl/nHv9zdWFmCtlPW+XoFWvBgEhdjk
RqA1ecDJjqlhad+OD5g1hT3IY+JJzaVQ+XeVuavU4Z4xb6JWgaBcCSKPkimkIwIg2/ht+izhm89s
DsBjWWvoowOJelq4A/93R51R7OciM7uKdvh4T04XhDQ2llRbwnc3k10K70zoBuZOXa4SRfEIGyZ1
CLyWP1NGZSaExQUsVIxEAw3f15WxMaiGNQ4STozyldcjmnnmbYDKN7/Dxjb/ztk5CVqGywGRJaJL
sDnYiLc7gLCPhUeKdcspb1fCt2JM9rxg+9uo6hmg1BJL7nkwbeIv+zlIe5/C4j4QSkmrt0HGvqZm
gjVTE+fS0EVtix6GJM1W4QwNaYxes7eSb/q9ORn1a+JQm/3sRvihGJuKs8+7fR56rinxtFajFWP3
Rr0Vm3YawLz9SQZekE96qIGRd180lT5sKuiR6PfBsRt0KmqpGdvBLIaAj9NJgWvowd25gTS4j40g
DUY436sNIhNDRXNQmY6ZAmzT8v3z9z+xNlzKy2daeEfqe7d/KU50+bZ5eCW3aB/Gih+DL1GPikfa
CozBa4RKawUDdAEXUZ7IHGi6Z1DMRTsy5S28M4axblZx3LvDMvGswEeoTpGjXyBf4vdkESzQ/JXe
uBkMI6Bt//23g0NbWMa/OFLU+5ocG4gmxLzPTSDqCVE7ThZKzXSzaTnzJXe8ZUVbbAdaLU4/qpQL
PIAuUUK/97zC7KK7JAuR59rmfV1uQcC8xOc4l6dcoObS9b07Z05vyMz8T+1szEKNjZhbBSXm+9Vr
QJHzy3v1QXVUuOhHP/fUOb33yx3WjkXcr5jWW009BSEGWbUw/6oKcGq21frB8rQOedrFe9RQjD7P
MGX++9DC5ix/lwO+iNSjrUwTbN5XpzrRVxn8lq6PbB2qMHmSLltl1RglOc4Oc8eXuIZnmqmcv32R
a7aYzI5B3iCONfBAN70sI2BiLyN0DRtXxTzJblUhvTnNbPSHYe0+ZOzDEhH/yE5uY0dAs+e/l3el
0zCOCt88LfRE0hwCStQ0Yh2jezkCaq5L5utTdti0775kLakwiI7zSSma6U7/qoeRwf4lkjSwXIgB
0wReyYCs3XteS6XbkNyQw4J6R1aLU6kWoEoLaEBzNFHxY/oNLYqzhynjTEJqbSmk5bK9Mir3Q1MF
4l8EJ9K6OAvEzqsmsLAXvMNdH9jk7G6sG69AB/TpTo9zM1dTikrhPd9cLcxX4p/aZFYEL5gwWjOZ
lsq7JClQGP9nbwTz8Wg4+7XuUccsqL/7RNHCm7JejdW2+VYU6P+07+ngEVVELec02t+1sgtqBMi3
++HtkWu+UOMN+QszAibKAQEluUVv3zOeKwYYhYXaTn/UykzmLXCvPfmxTTFmbrxi+/ctOAeusaOq
l4ybq4PRYaErk0rDhMfZ9LuUA0iHGEe/Upr9Sg7Oq68mH/OvyiOA8NKcQCrReo7MqI58Yg0Lo+/x
skistDvGg8fjUfwaT3Lzf6NoyAeQItQSvDgkYTxyQrpFWNs9s2C2wq/t5tt9pE71+GITwYpBxkuA
OcYAXi5+V+zDiaorsNyPBfwKarW/fpOBut4zLSsSK8XldXFWajyuKz0pqsAhuCQ+Jccs4xWGEnMW
rAOsKqUWTKX9ZMml6D6/wGPPPDc84EpNvvcRKj68VhHY314ORGRW0FsNKEiC9nHU4uWkmxBzhU4N
rUFuy4eNIPqMg3A5zPKunLuU9y+UW9dom77QoCh+TfpFYibrd82Su2qYWSGI8cCIQI+oBispQvc9
0muedBMbHlnmdGJBiMMQ7c8z+gKGC/WHuSC5PZQC06WiAhtdHR7wG0oqnPDXhMAFtTgKJkni7NQr
pIbOtnlGySzMlcMKaAmmgj/xPmoYOgjCqVtWvXslflymRNsLdFNfVJ20eflaqyLGX+jrzZXK+6BS
hu7uO0TYBKrQh2XH35hz7RroOrBm7qkMEzPAQBghGODm5II0E/g1aZ99oagJ/li0kaKTtJnz2XpP
3MYb/4Sbpu/aHO2zHcn0dVQS7+B9/83rh3BCWE+Ew4XKdnsk7HDVUSIqW/TfnKC2pZZGh3xcJ9N4
pwHK7mJJHB+BuRMxID9HZ77LhHRw9IZFGjMMpqmTZ4WRqg1D4BIgx/Bbtl7sTHhLUljXASJjvsk2
ciEcrI//jYrsMGA7utjbAGM/HE2hMlgLzJ/A1d38VQwWD2vfRyx943X5U2EEHmfb6YFshu1dSWnU
zaf+ZFgijREbsU9ANlGMYW0WACgXf3KmPl0Dp9R6eLzIXFMq9Z6ODEdH/Q7NmfHnULh+n+pUe/7g
9wBMd6U8L2hPnpdlIyyrw+DYJFI9DO6ddnKOhajj1uQTgAEdRR49vrU5AM+iUL6Ebt9TYR+5cH1+
NaXQIkJqKlr7kvHMqUDHmm/GSPFP84CO7LWucTbTig4WYxtlhBfXLmx6C+iU/hq0x3nSyT5zOxEC
2otLs+Leiqgp/OWMWAh+SyxE/CwPnidD2aGfEjNQApnunzAX6VxWQM4zTZWIc9jxVQi7DJjEDFHt
skFZGRD3HgBvLD9nDKBbKMhC5C2s2F2Jv5ToYZnVL8c2CGkluU+9FYKtrcVfW180owNqS63LvMN7
Ffe94EFwU+jHHBGmAaSoixcOLQkZHDrBcb+b8vd5Ii629kGy804pPKqDlYsuJi8QjqjXDiGNiOEX
d4do5OOLMMPiW7vgBpP5tmbwHOzowjmcodM9fjCvZ+KmdPp0DXlLBhcP878UkLf5LmERDL83OnYF
XW9Tn/YvEHt2L75jb/fz+eYJniScWT8tk6KemIzbqDHnSoqEXAK3zwtFxFWd7hN3BDZvX3m1RA5h
GzY7kxIrGxZhvteAJmUp9o9Wqle2xQDnsML2+Hb4QVQ/y16LCYb76vO7DYii9NOF3mHzHa8WUc/t
vweXCdZA3AUyTz9715eKU+62LLoPOD2wFlWJ+7RQq4mXiNMMMK8uCMicdZRW3h8kMWh7GJ3vN/CU
ym4y33iCiUESg/iTnjv8z48r9Gu7xWk7n6TRXIm6A2dUFDR5p/Ce4FdPUvfPzTEREYVyV7IYnAVV
k4Ln6qRwytruvVu+JMkTuGCLSkWwnxD/ftH+vLYnv4Rs45OAGpavCdOkVDlV8rHghsqDp98rCU9Y
SZUjkGrClQVZNnVEC+StUNjCi2NLSjgKNEcZk5a6FHG9sk16VZ7C/PYxh31WB5H8hNSPnuo72iG9
c8pN0wEyPfoOuK1VyVTaI39O4bEuUWuxY1UcaHVlIJpy5TYMCg7QB5FomsuFi9tZkPGVDtavJS5d
EcrA23sIe6/mpdpyo0QL+gZ6IjFPlHt3maLH8vKt+jrxhauWTwHAJTQP4rvsrat3OKlVmwVmz8MC
xp5nRZy5eaidUmEI0PG1YVe06cRxa0rePT+aSDS/cN4llOkCKi1hsUbxF7Y2gWFX/CsNm5ourcfm
0uc8+dw0FvVV6FgJjR8qINmWSqufQ+qVN4FrNv28j4wLUVBcuDsiN69cpnz7RX1qy4qREM/a0xnc
IFpEoTrBT8zzqWqzJyUe8GJA6Z8PZJ4xKevuf8815xFYKGeuA6NMjh9+eb18x5OMn5VHVLQRTZnB
XoB0Mh9wCdCaWN257hshoqY5Tj3Zqftj3Iuv8aOft+xjW0tOr39DFn5CDDvjCaMPT6iB0kA8uqNK
gNuKPAjHkvGijc6G1FnoBixgAPjyvTxDG5DQPO55NH0PNEortAouZFOoBQn70O7F3TQVySeL/0F5
QGbEe5MuyVW6AN55nhKTdRTDw0dF8EgGKkophfvcwdCVEzXk66tFttRDaR/WlBqjx+kufRtLxUP0
CjUGpnyH5kBxpy0o6ua3gxX0RKCnUSm+JBTy9ygYnUrUaY74BVRui769jNocCZ+YrMZJIaXfzPdZ
upGkQZofVkTRHDrCBLHY+QKVKMquwnn8dzjXQhhi6om2QJSYCIfSDH5/3YdCxjM9q7SY+uxnoCnc
p8HXqoBYQdB0b5he9c9MmFCS2+8gGCVs4pe0vNgcKtDcayCt4rpuI/lLR8GRVNwMnb9MLT+sHJIe
8y3Hqpavy4Q0X2kFWRrtXnNI0Lz7YnOfEermeGkSZbZg32l1V91y2csnH1qD3kcEjUtObi/FBEP1
mnd2z4lA5rstbCpOw7U2SWqTKBxcnF7wpmMxePTsvCvdMTtEDwxEl/uVeLzfIXvRNWF0Fl3qMRVQ
74me0pQi1nHQiTx9/pYEqBVu8DJeLzdJ3RVl9bw1NTh+5eZeHkKmA60eFGn6V3Wo+3FZ5ZEDTJoy
g2A0NuigblQwS8cuQ/KRCb2D28eaNohscjUkooakoJfXLA52GZ0gSP2XK2V0/BlZZxIDzyjRA/30
Y+UsceRO5ptJxld8srJ9Ioao0RiP7o+p745t254pDhg0gWIQEqwwbKCLc+0vkc36jdp9/lBAHXaz
uHz0uKCxRF7Km81gYG62fsFjwJYs+r/BUC5i4yGVN7HmDu1vLyd0CzDuK5gDNY6+Ivji//w2IRFR
g7Q61uhl/1b92LybYZ/eOw3NFXEJry1HyK/9RlfhRAvXsgQRE/Pu0vYHPwUIbOGB8VvDv9clIJ13
ZvctCRiZlC8GC+MCoBxoxq5TbwIpRqS7ZVgvk+WYQ6U9//9Cusa9Zu8+YT81DweyyyEZNwtcLgVw
1FWmrxvDA/UteksLZ5RerPGRilIGBjPeq3mbg9HBlgr9isWdtnTQA0LLNM2xQP+UlfpTr6uuk2fB
soAAU9Oq9ZLV9slTI9SMhzVgHCDWfnj11gnYuou4T+gOWS7c4zrsocxM5C2AoZMGjJGIZL0p7DFz
GTP2BnTYvj4YReJG5OfBRZD1xxQezwxJ12wEL/3+W3LKBQkKoDQ/TVUcRhhbTfJOOH2KUgT7SQfe
pUeTQ5MkCUvimiKb9oL+OhCa3cwIb0ebeaeV0SK717A5Vj09O80H0Pgr4wAE6hzvhHQgxcbOysMm
mR2QTtfg086aK3jOb02luLhzyuUPOttMfex2PqFZYrJflvNnJnjZloAhLBxfGkfE9r8G0S0/gAyB
NlEzXfzdUSp0htFX8H+y/2uvfcAYe8UQcQONIeSUkyNbweLcwYoej7b+1MxyLVL0/7nOhtrXlgIc
tANkTGCVuopLkjvDBzv7g2ThSDARo1RSu6X4g7W7+UOtNin0y4pOYMgjheB7yQkhJbFbphJBZvz1
k149WV5L+tdWlw8ClOKRmwGew65UrxupSDX0OjkiWiYsPReCIrztxF24bRaATOK/ion91m67WoFb
1CtrAwH5ND59qasTe+BGVxMqE83hdPqar4DPbrwIhHd4wtGRRV9PWAD1lFiuAm/V5ikTIO+s0X0z
8IiCD9mg1Eqsiyx9qLjD/WLMsWNE441nnVQT3okVtYUyHzaK/DPciTqBbyj3b7oPRGaa8U48zTiA
YVozjRPL5KR4PAr/3AooV0R9ed3J6i1ISePvYyWklfpYrAHJEkIYlT88+fUSpOwcD8KhsXquNvPH
jfGCTJS2gaJJNpVUY3OhXeIUrjJoF0YY/XeZl94Nebu4SmTRQ03oAE8FIWf/+effEZmghMgpF3Tr
Z9fy7o5biwQjII1k5pN8u5BG1J9XdCisrpXPTkEn7piqr3J69pV8BGZXBjiRrDYXj2ZSr/Tig9Tk
vp8bMl2KyoaEXKAeApJyenK7Oz4RzTSx/zhR8QOVMHPpB615iG5GL0Ulys5h4Hc7kTuCPqol4kWt
Dk3NFDdbtBqvgFM1O8WDbX2FAcc82pmlKd7FqM7oCxRNgh9MiQMHyfqgRttamoAhjZB3dqjg2mpB
7kQII9MH7YGtxDZhK9/xmw6VzuTFScFi6iusEzOwbXAvfgMKpnL4gqIl2GafYYohELuhZep1AxZz
a7J3doOWc/m5LU+JnLvvxpHMaBYkTa+/4Hr7QNbp+SSLjkBUMAAtvY5tgt4Hab5GoDZ2tld6rm9y
4C3EQBhoTaIeQXWMQRXHjgEQiK9pKZFgJL7Dr1s9KYBVpzV5ZHRHugQfLqKxCKThP64GYtm1S1HB
stvCz26+8yFIaDGavRAFMojBGWP2EDAMy92BwBGimPo/FPnRdMz1J8/Fl7ZWonmjsE2DTj+5Ux3G
XXskyEbOC4ILxzXxe+i+WbPCZVpXyFHz+SD9PFPunIcq1onwD2YEjP54l3kFAXnZx0MYnEsPaAHc
VfARqdd6/FEQB1s4zYGw6CKktwqjD6mhKNDehQ3P06E5w+qvOTgVG3cePUmfDivLzMJq4ZYcMmzo
hAeL1EqxU46m80B234Dp22U8XKi3+KDU33/XO8G/HWfirEvKwRe9QnK4xjEgf/ZAS7pIFQ4z7Msd
DU6nZEwRY9afukohPW8ud1rx3U6bly1+7nK43SFJlOo0Gb8l66ttzyqfn1p375xmfOf1DS5kd7V9
BBCLVUhL0jK5XnZ/NVIuIfsxQ09EJBhCfl9r9ItCPruKH514bqlX1ybfrXfIbhUpVwNw35afrc0k
0ayQKARKgPytZ8hkBccpeV88h6S+EbB3me5scSyh/dmjpfDIAZpcBlHcEuX5xMh0O0lM9CF8YzZw
pTLAUuuTzACF/HQL1Xm2RgtsPwWaTYjyJwHYisx+YWnRJrbWRP+apmhZpcAaw+lH8dMwNHsMUB3F
9gazEaEThTWAcCd2UT+mtnG4BdElLcTlwG61V4IJiiAlbkmxnDaX2ba/LK4mjHBZIG+pkqaMoXWh
kxc1qWYOTkNW5FiqbbUR2dqQseETP+UJGmtUYEmuhPr0rqkCqd6mAiAJd0WQsuFC+zBUhEcyNUVP
myckU95vRsdncjcxFQXgh10zSVZOgYlFIL2cebfqOdmBiA36oP4eLlxTtjHgxTL0TOgvp9eUgxS6
M/2sAsSRB0Egfl9lqCc1OarwOYRMXwXrwoHKDo6V1H5thkL5DEQ0y3wjRjWLisQ8QYN6TfBG6XkM
1qAhk6dUCf9UbIejIpTyw06zOS77NAX82S/B1OVrJYpEunlwaMpMLV8VLZa8s8mq9wyaMvoHXgzW
nrIK4cdgfYSLjzxqV46VqGQgBX9VdBFIpIXNXfSRMT2VedEPNszuljvBkk7uv1/wHGl7hd9ty3XX
rZg8hvo31WGu41rG86UYthJw8ACOKaxKSHsIAA6c+1Str7B6XToA9Lf4CSUKI8CexaMwJbsv7P29
y3EBZuQysm9CF30Z8nS4LZZbyVbj4Q37xJghBHAM+b2lBvs3L8Ts9qzzlyR/oGFMnZ1K8cfiItCI
8nF0Iz+pLVqtKiyvPhCA58xa0foVtHY/W9n2VROSsmI+aQDC5MaLIotIlOGT/zAGw54k3DDdvD12
2VbyKkSnx1GqjW2sgt5yWFLuRaT3oyaAoP9ioDCcqa1So9ScQOgRBV7S5SjWWrDrkUvoevV3k7nA
uQ+5GMpjeAW2muvfAEK1vfXUwXJ2babEW7LszZrjeVZAMLSL2A9hB6CdyZwzXYUz1pBhjJkUljpq
PyHqLOvqCiyUrL2jWHBJXow4KuaTdO962OHl+9vm1B68El7/xL1GYmWFYg9bsD3b3owFFIXHkr5u
ujcXpASYSkOkojcaMCS1xC3zOQJz0ItGlYmswZLM952nyoTlKayaa/9+A2QqVZ0XjpO2Mnfs3dpY
Kg96mAstYE2IWFheqGBfu2v3ZKo84yWWHFYpklHQphxO6v0JCDCn1Z5479rgOTjt7gnmCIQ096KM
pJCzguGUOs7CkIPu9jgcw9ETZgz2v2o7Pn31oz4XIWa126J/tht7ZV2+v6QRH1U9Cx2z39DULMcD
6EL034HGzKVRICELRBOHa0CrTyo0jbjd2zWRhf+kPMuJ5pAXNV8/WB9qXVqFTWEHK7kLgF78Dk4i
KdYWJcsiaAts8mEjva4Ev+eLQzw9sGu0WdZenB2bJl6Bi62qj9f2sbQoXPWsVlLP+RE4n3htyYkt
TFgSwVQhITu3QntafuXy0jbz8tMGUpDOOLsKYUlKBSwm+fQ/pyiPZL/BzsmYAYOqo+16eduST4q1
yB3RX14rfve5qW3iWXFShq5c7GKVcPYIeaQ0CumWlYHr2Sll2vER5CluKWs9qc/ZrNnW5d8deZFE
zHsooLFRfWH/B6bDPazb0C+aHIW3QCfXRRpYPr5PO63wku709QROhITlFION30oe3jEliouAxW4v
42AwCyMYbffKICoQMrwvn339VlK2ZYdOtO6LsisSRGFo7LlKuRO7ByV8fv+WYP0WJcEkYAmV1MCi
spSMJt5nb6igjyxcsNomDZQvVZdt5x+lG0zHUWgyY1P+P+URi2Gk8pwy6dfMqLBa/wImQeFzjJMt
qH4P8KQMfyp2OOUhE2eknCZ35K+EqdEvIvVF8jod5ExJVachZiTuFnXFnAq/iW0hkbLvEdtcEmxy
Mst07DJBJBjB1ZSV3fjsLuYba6KYGhwDXEXEeoqRXEiirftneDzGlNq+8rgKteZ7CxLDw2SH/SVb
k4kM0cntcQ/gxlxOSddkFY+Ck7PPxwD5M63LubkWh/JoHj5kvJlzgzS0cB8/eLRtwL9TT3Y6KodC
O6W6QUjpSVwywaUHGsRgjciJPcdfhq0PjLvXwihzfIsdkgqZhKjzOC2j6FNfy/erRQwttry0KnGm
sJUd4P3zKFfzg6C/cmCumpYih3vec73uEqpsKSfMWrP5zG3uL8YeRMVm9EFxGoUDTNgHZGqYaWFh
w8Vq2baK8RMSgW1HqYb10hl3gl3tYmz21amBp4FcJVyTrmq2UOglg9VWO7TCU8lV/JAiuGbONhI/
uvPzCiNoET+yat61Lf5zYd6eFBOVsGF46NQnLmDO1mbv11+MU+uPt8jjfZbN1apIbQ/Dzh83juwM
Q6lVTxgjaX08WoZ6oFezQAgw7k2ICybpAjK+e7YBLZjsn4jIATL/2eDZRF3n9t/FBBRadrdjGtke
+aFouOLi5m86vN7Sd31tQlk54tVM9pgGRlrk/hlyxYi+fstSXKsA873s4WqIUeN94AOWHXW0pDj+
7wLVUWTGxNzmtSLFUU/26eSzREl92a5Zprom+K+8GFn/Tin0xXnnO4VkQbXSie6nytc+DUU6mCyd
kaVNZkKhlPoojH7ksT72OUMNfOE93Azo9IYdaEAlUfSAYNclnWENwGlfPkf1I6jwuZJEcZ7GJ9BA
4cfj8hCvIok68R5DVeDKGRP+dLP965dSMBqT+QH0CHGEP7z3sSnf3hzW1LoLKDeijujtucGaj8Vr
o7zw0HEYRhpSkGCiNO8bgAGDdAvbQ/Q4tSUl/ZgVmjFRNSxdqQ06IooBaGr3GH/XxbVInogVV3Sp
z+V08bVKPcYef1Zf+YDDnPyGprMnoRQGo30fHy6InkHeP8IfsDEehasW7gIjPU5aVBiwBeEhusB1
JvQrVD/qWHzhjjHisCC5DuQpxniOL1vUdZa/CF1zJkgShahqBhTo75O7Toml+Q/zH5pUdKO7MJ43
jo+FiVZb7qKBO30ofUQvRB6x+hhsOjNGbOtUXJcaOCT9zQfx9ik0cHB+59ZuyshiOV9gFn4oTQas
HPtVySj/UpJ7I8elnXqUdtMkyEjXM0W2d93IA896OLvdqW538mIyYxasO94h3RhO6+o/sZViLaXJ
KvlFA5ovrDZoSh8wR3+I78vPbiPY28yqQURNJfSt6EE9lIkpjO4JQrFIOFvx5UAJUY/UQV9iMKKd
7g2VifyXuPsdR/jzFMwH8k4KyMjIHb4rKRioPEbj7VKSR5ttCKx7AqU3+umFHYkM4QBiDZ3X7moI
o8VPGvWMIWM4f2yNJ0UvWUjHCop6bF2ojWck6HTlesIT77xSsLB2rOnFknWceIM4tzhrQlRTC2gn
bxXM6Gx2so0DMTz/5x4RgGYQh4AuYkGZ0/UcBHRyDIjapW9MuG6iaTBFZvZreB62H/UGDhOCpc5x
7YL1iSXzP/UFgMA4TaBna5V/FutjgN4+erhTgvIHIoghmNloTI91Ios2PD1Bu2SkdnPUeVls4o6S
gkS5HtqD3N0UVMGiinaMyBd/zY6dV8EVgcxTiguXPZJ81HiwcKfnuH7djG0fIpa5apvtgtKqvUVk
IIph1mBj0SPa2tSSKtRrGyvEo/cgZLKUbXiMK8kcimcYLooGB5zc1jLNJYYBJwTgkI4M+lgW9SL/
R9vXJ1qGi3eAtTiOVnHuOycOFn/i8Dmc6AgAX5Gp3Ge/r4qTw6z9CHYQ5zYzh9W9XTCU3nZDPN0J
pRNDffyR7QvHa0X+yjp8tJ46XKjsAwjF5c+qXV8VvRllxL6seD56/T4M+5AHHLPflhYX/2Oqz5Ra
mOR1lZV9p3fAZNzK0UWL8IREmGNaeK/jO9SFwmIZ8YxzA2JdtURQoVCpFli7pzYCAHcdU27HNXFy
A7FiDSNBNIwMXW+oEVwVUEByIy+EJPOXVTT6ywlVCp4flc1AqvLkcew6B38DT5RNxKecJK4DGBxz
SSOPeNjpX+QR+yAMqyGMSFqMS+qTqeBJUJtQbKL5+OZRk8fk6BQPFQFWmzWNJAy6EMYIFKxikziC
sZ4qni3PrgS2zsMnLZywOcqubxRyqweMyN6tPPtMF/bCYn4IMuxG19zREI+kpUmEHw/5HtDOyiH6
a3burFAkLZcjgbRxV8dO7bjefCr11P/nqaldUdD+TneYHQNhoRkbhqPIrKGY7uhlvvljmO1+SFwH
tiUyUY9PGQOgPcU/LF0nyNDopsGp4dXxeyT2gkf9cU8jXOZp6tSBA+L/3ztRXwUMkOEshK6HHMpf
0yqK0PWEZjiPaUT5Cw4nCl2qZKFQOIV6VWXdQjfoPFQz83IZzUtT6JHCJ8q+RMLGtYvsxNCHXiqs
zK99v2Xm0+dvNeUqx+yOJYIW9oWOb1zfH/zb9LLExVZZZsEkF3QRMfLzn1UVjOeGXUIdhUCq6aS7
ZjJ4apknu/j/4pHuem7W1o4+XNhwQ3Gv6PvbCloxkp4rISo9TokIGtHiMeVXKYvxxMcYrBQnHeqa
R0GafVTleYsjkJ79qgbnhTr1F7jeiQD8FmRXKD6r1OTw/QGZiLI6TGgYLp4OJ9x0yOO68B+qiDk+
nYNeSJDihXMwD99JU4W40WhhpK4wTu5DOOg5KH9m7tcwsbxsSzUBAgn3P3PPjwpebOXMr258uw9B
3wgZmxbygSzCjbO69F5NR0+BxKn0094FQTyWFyoPq6S+Kn5YXNMarBfG7i8vagrJkTOR3vUpz5Ht
TNK8jV636n1Tm2jJdqrqMJOtnxqaiCXadWW7yAqyry3awT4jgkjUppOdY9ocqFVECefpy3rs1ik5
P/4RMuGrFY5zo+jYHbS906fycanMknorMDEVfqFj6OAZ4uIsjzgNPWuf9RXwGvBK68tXgoxVb9Vg
Ptxat8pvEO9+STauPSiaRYYciQcTzAqHy8iayPlGJLdyvYT7q7x1C0zbdsoR6iObb3IYXnvvc1sg
kN8fIa9+QCcW6NEugMJfQvt/j2ea/9YpwmYjHwHem97Em9isOffR1RwBX/LSujrIlCBzG4F3Bred
icxsss7nBaX2sbgrsFfx9wRMaKmDSEqHEUxENHz5rLazmVlLW7CvqTF4AhAgC6NTUVOgyeegWMnr
5rbnDb9NYLW8fOP6KS9NMszjwdtjvcALbwqG/k/nWWjjH7mKz+d5mAZ210QoB6JwdEp4zW7KFJeB
T28F76NTZNJNd6jk1+A7BUXf+790+Drpa1qnzBwMbowfu0pvDEuUGdXNd3ozzplcCj0owUqKSYlQ
be2bOmOGeyx7/FUekcAxAUez0k7mpntoVkTVUrwMpUfkIBx2ex3w1kJduI3uW7QZno8A53g4fP/7
fEFLYIqAxh7lL7bmIxnCWZ+VVYlLgHHM3QyUErnDAtOAgyodUcRkKk29pdADXGnse4aqhyjhNyjv
XcrZKFtnimOA41OOkKp3dqm80u32z+IjvGJaoOh26hpp55N8uQ20zfCkOjuhz4OrO07VxWb1K0Uq
9vXBUJbNIavEvJR1kf3JQ4FvruMvaf7tPvzXBsw1PQaVWNu+pEUQiF5GuAjfgbsxNe5d17RwLV5O
J8pJSOJrPdnjz5L0/bm197gp0il6u9YMNakJVWi8LUK5r7p1fKPxVnD35XUQFVQlV7vFStV2g1xg
UPSOohdyM00QGeF+TvPMN9k9SmAAtzYeoETZ5V3C/NBLMtj6cnoro28eqKKGD/e/fnrEHnbHcJuq
IYYFGoRYzmhHWydgnrbhiACe7CjrTQiFfLL7m5ctjxuJAS9uCZYo/+D4KW9TinyUChm1a8c8JgjD
THKyy5otj07WNALgBL00tIQw2rSQzTaAJ6uc3i8Tz5steYwq4YJUKKTYGjGD06DDNV8VGl/5LEwf
geej9kwZC1P7t8APBZLV4WQZ5GxDs7nqhXIG5aNeUeMTG/mX4Ds9izsUuF9lXtqrS9LAbWm1pprU
xZoi9Ao4eVEi3mMzeCa75x4NUBfn4rwDXdgthuR3WLqf3P0qN9edgywtwyxoiVtx2aA21YJFYs1U
PQnV5CgMxBWYimyGsMOgZ8f3BrOTR7e+sQOsfmvHJ6ngCAFS2V/WTtVJnHA681AkmYKPdm3cVV0p
zZOQR/cWcj41Ivfx9/i2IXq/lStq2EEfJ4OIbdiirTu3F8v9X5Tbui1S+NV5E+qkt7XIebrKQCp7
JM0nt/M6P16YSRsUrPmS8AALlFv3znS071pTyaqOC6lqpjUWWjgxZnec8ehvooW55XP0+F5G6UCy
Dw8ZPVoeL/bm/IboW4cHTwu0uurutWrYjJdJwF8wKNxYf3MZIX94WZ3c7ARJtkpLzM8Hv2aDp7W/
GvYTh29EAUsOwdIa6Yy3BIDmNnQ5VwLFJHmg4A3IzcvK9QqLPc5Pt+BfOijp8hdyoyuHjfmcn6Lt
Gclqd9SJpCr2f2RP/wFlgLqJAsbbQfMvQ3gBbWsPaHzUt8c7sgH07dS5fm1zyyQukiFAh8FE2MmT
s5clCV5G1zy4SKWS7knc7hi9Nr4eMcBLIRTSI65plAZcx5S4xzFYmXwCUlUm3hENbkPBkhYSRRMJ
qlZCFsXhfwkzqSXf9qukZnzIcMoO15V9xLux0ZGzQFL8fsIcgkPaJNAeOKZL3dEao+aGx/2JOmGP
qYohLaWN0P4Maew1drED7ZbE0bACFRyPltIihr8KFO00X6PDctH/ykDwVhDE2S80InM3hdbrdNi4
XfTJkusVdOjiAqvV5ioZLBRRhYA8WWVA3xq2BGXHBdrH4ZYs6LDt2tUdm0mi4LDewVQjuPxgOjkY
Ifn2nrFxfIu56zyy/e7nrsaDpMasyKAy9Zp/nYsnx4aG/5FZ+7tHFL/ltOsmve0g0WijlcW6uwwt
/uVbP14KB1Odr0JzwsQ9FoZYOmH/H+q8qXdUKgYM0wTcJDsWyfBeVTjFYIpSZ3hkknWoM4UdUofS
zEDzZY7OoeSnWt2v3QFXFYd+S1AP6NCYt0fVk4jv/K7HuTNw6VK0ubFcFjpqD1sTng84S7UKT0TA
ll9+FlpkWeKjG29pO/d7LTZxdHClcPJUIu7n/hwsLoibilyR2tO5ln0ZWyTjJaCeGHdRpxTnP/4z
y266Hpyh4hcry1jOuhyuc1xD0kzzokjGqMBh3oSLKEpFCMHuXopPwwvkqMsRh0Jy8ZP0/1XJYqqn
cxUooOCaRMRyCVsQEl0CvmsgEJ1Snh58pc0cXXObtfl+l82150WxHm+Ekn8jBIK3I30TTiB5ul2S
QMojyO3JiNvcIvS01Ap+plaRpS9WAsWZQWLSR/FC+iI5K/nJIEcbBevUG/mvFQrCQgCVDBU+DZhm
gR/M9HpU1IMqVXSwcS/nmXmSZ2pqIZOtpgUsMd9cvrj6af+hm2N2pwI5e7CAmU/AhhmJVY6FFk02
DxEEEhHeOeYfkJfBjDOhLew1E9lIaHJyyO+Ko4d4sZZ1KFYjai2C0tkyCVICSxLPXCi/p5okpxdo
9EmuLpl0Km/C10WZsAV1aCAWaVkhKETYkSo1c1ZJxcKbxWVyVgBl4P2ApX2tM7oH0I+IDAWAerzZ
RsEzPvq7QXMa9K2SMXGIyx/qTDcavh4xxCMD8TxzvKFxbnw9dJR2UxCj5rZLXZiwCpTBpOQhUjWH
Y0obZ3l79Kq0QfE0nJqDvihhev0WFR2MAOEOlzrDdzHuWRpGVg0OLzdxsf15/s6QBRoi6BebDnzX
lJRkIReZMhVUuyyL9DBFeYBcpaMC8B2l7WaYRGIxxpoNJQ7Wha9YosSmFwYYlZp9Yh1mKCtWgZyo
Q3HkQPHVpUXtCZcE5+FxXBaDrLtZIpVy3dBEHAA9Hq6dAXWCp8sVhYZuvpOyp0yrjuaW9ww9VbBo
/r71RkBbrwhMl6ANikvJJ39wezbhUiCoJLNPLB+xaA5E1fpd9cCblI15IsL272tzY5C6QBMcs+5t
X2tEDP51/0JNoBuqo86rqTRpDVFhATkV2fqt6YVnyYcGh1tluLAM7WVjIS5kp33GUjRaupoif3cb
WwLNoWssMyzrZO5y7DGaIE6vxKYXMnfQoq0jmG0XFh0IT4QPz9I8Go+Cd6Cm4IhOSH/VyhAj77N/
BuYPDC6RfKG4NmSJXiMVYHBWsOHTGNlO61M0I7XkYL5cTaxV9QqVY21C7FNq/QWfIUlwjqL9Frsc
n7QxyHiCrgq0/l0P1QoHsfmISK3F4BqjllYaALoLxZ0cWGsvRsn/PFMX+qRwOh33yIRS4zaivtvT
tex/w9W34RNM13LjtSZSrRaIItNFY+KosUdFenIzRkDJoQb8r38BbjUfF6wppu3kl8/K/gkPiukF
ECe5jpYwUAgxKrefLqhkL+bAAdxPefSfMrzmo+uK7kn9ZF6SAyagMV6Gyc946ruV2nSmcyE6hSxB
XE6iYuiM6G5f76QsZytg2HgneQwIH23Jph1UonyFbXbsy0NSm0sUPW2jQxzJzACn0JLYMCfiJJ7s
7tvf5ESpvRl9iqcdoqlh4P8kYXxjvAa/cXocCf0A0nz6T7wecM/oXrHZeH4l/cOl1FhNgQxO2Cw1
dTL3F+g4oKFrvD5gyOU3qeQ+APKwF++tfW9yfx0H22JLqI2j7Dz4LR9/L9apj8R2E5ImXB04XfeP
Md9c4UTvBhibCYKOdSeR0AxxikXzgFI2dy5pfy7w1ByjoqvPNFr3vFcg3DF93FrpdeJxV5JYPypG
rsfu91Z/l9cdPJ8OC+6Fou2BS7AqCxvxaxQ84lWEd6SxsYMgXCj46OMlhoXuM4jmqUwZ3J+zjpNL
D1B8cFaKMMFr8lIDW9KQpfvM9tDmU9wZK8h0ea1RC4nxkViMars8qMxQX6O+zoJlacF/oDzaqr+r
LkO/hydoflIdZwnphNGEeNC3GzVlcU7ipAw3EaLVwLff83xtrogsAJX/CisZBDrFKXs90jjiJ4kV
OHjgJ7uWi99zp8dDv/j5MnR7T6LbQsybhe7nBywDQ1l75RWKQIFjNdWQkTFmmax/4p+BM4gvMmOz
zff96aOoWmPT4mz/XfUK0NvdEGkUT08pM+RQBq9ERGYlEuZw1X/qfhjI4UoaBh8nEV4mSJLzGa7b
sHaOTdd1EkfVXNlfwGfScosk7R9qLZS1YVaEdfb4yJbtrRJUpOD3wPytHA9TJRQ8PH9SrPBfYdCb
Ip5dcBmvAEC6LcdJu4Ag4C9Ri18SkSK4GHHOmRTJLShsKtaARi2ryUUc8KL5fbZmIWZ4L7bH4ojQ
Xgjke9qH5ILArrQHtGoW7b116w891FXBKYjqPRyRuL06+IvNdzhuXdjKComcjPBCVbs97H0lqhXp
spVRC8rX76zwQrwy3/DcAAvdSG8cTbbQHKwRWQw975LamfFf/iRLA1krjsZ75qE/F+kFAlicssya
yGU90AYwjh7LSXIHF+xcKoXfN7NonYSX54qGYU/XU+gbLREmHXnKpOf/mYhetlNicUyTa2crNbIp
5/tT0KnZWFw9mc5mjK+4ipkD2hRV7AX3XXc8Iw15X567eOacHvbQjYY9gGIaSdw+p6bgQSqXfjZt
7In1/Np+wtlfWm+gWiuNEseIKL0apjMktnu2PFcNGUmI573WFWpPBSx4OfEbffW8QXWxxarHxFdF
Bs4tkFs50Q0D/g4reymT8J7tKE+6v65nZa53bWtdMbguaN9Zkw6jf19flaPaUNqt5FySG/aw+GnU
+H3sH4njDq30cVc5ChNdn4doBsYRACETAVGgjHKhdrTSYm90Gu0KecOuwSvgHIIXvwjIukQnLiS/
szBoQgdQSm5bygTPlBcDO1Ml5qcbu66RAcWYj9TNNp/0lBQCmTQ+/CwdSYMlrKTc6zhqXWPChYEt
8Y6KxL3y9ueORJGz77LkdpO5mSv25cBy63CEVSM5WoyzSEUdt4FxQBHVU6NJ60UEceaywhrxi9jn
0RHv4xbpY5SBlTCIGUhxvJa9borUPzCV8LE1FcclaJWHw+heXQRkgoEBFRc17hsY7Bvw2AWdVCdT
yCxBfy7B8zfJfcj2ujNV0jcVeg7xYzYpo00gGuKWcrcoC0aeSeRu8Q2sAe+VYOeWUVmAPRR8vyci
qNL61F67wFbTHMR0axXCYY5pVgg3lUOU5eW6e1zenDPRXoR0nBWI6+3Wa9Y/vEr+N6Se6jwJuZvH
vvKVI15OVoQ7fKgBT4uamDoIDxkTvkR9Ako1tomIKjRafW46aEUrpqTDpRlzwsviAoXiT4SDUR8D
+O7locNqkZFrZEiflivT3SZjkncOMcEIDpJ3jRRBtM0uVMgXnUBPoUckX2pf3gQyYXCgvw7cYEJh
9pme+lYsyQV1ZK/Bxql1zmw1sdOor/L0KyKPAUHu7LZJWfEchuMeFqfXoYioVVkv8BGp/y4GiYrI
36mDhmquNePVuOGfeRCHI9qJL1QFIT2EPfMC1GEKOX9SPwFfTo7494gUrOwbvtdQQ5vI6G/6xfSF
e9bnPteQUztb5gygugpFAbwKSzZR6+1JW81JQQWgSHCqiq8vddcHAI4voVqna6tMODV8GiuUqxID
VGMtscfjzHlhQCdtnv7VzHf/9L1ABWobq5VIzpbHi8wi8EXBePBEKh7k5lkbAM2uj7MiGkLwGNSj
1o1VjGqlG0wEKODtyLn1KczSljlYpxbkH6GPva+Yti/3Q1yEmVkDKUc1ZHFJrLxQObGO0+DGSO5T
RTy4sY/GDA6qOfi6CiF33M0ey/rZ+ZqQyIGRszy6tBvkg/7Uy0zYPQISnG0krTj/636mAV+zC9uH
o9ZnV3rUd7PTiqT8mB0IPdHgeHL4NMJWU9VJuPZ8JolfpYStt2duTcY++uyESQyk8/493Q8VOP4Z
cqhXh/SIjG8ixiGjfOl6L11pXVMkWhrfECB6VYx2gfxL4KC4maJ5HX+WdXTEyIYvQUgajYf9Aax1
uDNN3YNtGebSV/MPaBTsOzXa43w94dY3qBJUdpwtMPvGWmcMg2BLmpDQjhiBh1qEoHlCf/cpHGVu
CxB2Tr5AfKJowX8iUTW21C9fn6o6Oyw3XxAQJuuH6wtYDK+9igX5fA2Ao2Hz0kiTsGlo8eq/Tzun
b376ktHSP3EtL/sqnl35vubXIBuPIk8RuXJvJqtD/KMoEELYa/YVMXZ5s5igJJX+LZi7OgTqSdP8
/DYn9G4WCSdz/gyq1me0xTJFUXICmOL+02mkNPoapriTscwUZowRcvVAlaZDU8ZhRb5+F5y8RYPw
E+U9dBeOwVjuXu0LU4I4GZU9Q33LPRogKnwEfhTd91DriCg2j9flyuKy0N/7CFYvVGdF419FvDto
SxbWepSOGaPrp8W6EMXI1InAGMiyRYUr3+aHkifheBWl4jb5rPU/GQXoe1LXIBC/OUBHSTsITGD5
6UlFy8k7+JrGuyNUiWbDmypa1sz7IfjqZaZfF09OsIXjuHaZ7i8vZzbmDt5/9BbJ2DcsSU/zZ0bG
vZDry0cN8iiXKCUbMaJgrpTtD0TS2MiP6bL76/HAUL7srDbFOPC8C7T8dJ64dRSzE65/4QfliYQO
3W6b3tUW6Hwr0zf51zyZkuu92AR3iUMWzSv0J9wme63Wtf1YTMZj8nd++fk1k/REiHvfrkRJuxhT
KnEfF2hyZ7XE4kc9wdt/8iHJ8Fa9XPEJsUn9pXwsmSfoJRhRQoqPyo9K8KNsMXD5SYFRK3d66o5d
6b22heSUhbC/Hf8zErSqPAxPz6+u/Iz8fSNZ4cqzQK2DUK56T9j+UvPMmu8JHZPmhBBXowYWZc4n
V4GArB+YwI6js9ZXZ11fX6Srng2B1mR83wU62xXhY4WRXTubHILyAe39GxPHaY3b1nEBFMdqjnCX
E0m9TTEiHrHgwyDCPpta3kngkKguvGKyeGejgIXieRZdXH+VaoCSl6QCx6BeMa9WgYQKsrESUB1E
BjLYT5ZmE8B/c9i+GZhD7ZGl5rS2C4/+zCa9rQLa8jSDeFuQfFyAtkPOYxlE4qU0yoDvLhwTEkfC
BtJa6dcjA7SmxaPBGNtotMRty9/vHxZiR/qpfP8Yi0paMY1YOWZHsZNiyPDe+cO29I2eZGZ7y2/P
Zp/SjtoeSBtIlwUHJSU6Nk7btkPoBaj8lx1WrPZI4N3gdf+ZY1gKjmDgLl54fGaF/JfmsgbMHiE6
SJEeUaga+k/HzzGzQ2a0pNVNhZiVRAIM9C4vV1BLCOW4LVyK5x2u1/aikLPWIAOn2feeaZTbwS20
Rnbc4VYlpg9AsN1CGlWMGjaDx04IytJXy3m9MN2a72CG87M56Rc/2NRqDUZOXLylGOwHXWccl6/c
VsH/h9GWRvZ98yOCOy2Mrb3my6wrH87dovbOLtR07OwUhDgfKT19fcksTejelntmL5xaGcxT7OE8
yCaCM5fTLEKz52HXsNmCpkFE3BRCQZR4Ec1yqpSQfHzxWTx6PvGXZvc3UmrQ0XtmEPrWzub6NvFq
2srBhku1PDQJB1fDEPW2lrXWFu+E6bBXWxvg0lIizUsrDTSMAaiq98MR3xNsHnHeSlk7ImtzDDLW
Z5O8EhNiwV9EXvnyeUFhMBBvpqGagGfh+fPjE/tDrH1kIHqDlFBj+Wo1Li15WhH1eMnEvM6FGyYf
x8zwxFz5G42KjRxG8qpt57ugeA9pUXUjxlEkyzuJ66as7c/rqiTHt9iwXBh8jC3SIJIOSnVvqf9a
nBxoicqIm/aAaQBj94TT3saymjIiW3IAJsAq52xyym7VCrmqsiZPftnxktO/OK/1SO3IbUolCf8C
BZgJsTqIAEamvbwHcAIXsqYhLhBWtXcRPWmHAxztvrq4kkDedb/Fa6L4HYQWgnmsZLOsdjjBCpdc
uQsQ2x/P0IUmt3sXbtHHYGmy6HMMdf5knQ+5tTC0JPtvUSgArIX0rhRUcremFymXgNM0wWS9g5vY
cM2F8WJ849r+mVZ5200GFyUN4rHOqYhvRylEB9KWw377JMJusp005v1Gh48TbrJSJo0MdtDA526q
/7ZrofH/61GKJ2KLE72XrHnrPOCIUSeVimuzo/BG+S3T9uwh0SYVhQ7B+isdNwaynMo8pKWo2hp1
XQKbRV6MPwx1OXveh+XKD1ncygxVyIX1Sa0nmyin2KaozJvunf+KeIDIDcy3hG1nNLniK5ty9ehi
8vXJdTR/AWqbyoBeKPtJ70K9Aphz//YFvk75KeKRYQ0EbvRWUFUsDf+/hcsbx3CU9edApr8fH1e9
cSR0NfX5DcrGrqIYp7yxLF3GmaC1URK3WaKtCRkmVo14Ix2yiDFOxeCfFRWi2bfYZX8yF00b7RAn
7utTfSM/7W9ySzY8Lzvf693lK19UOsuRt55vQLPUrDCueK9U7cCxV/g8YqRgkH4sSzIKEWTHr4fQ
G7hSFA7Pf0Hu8aqQi4U4d5b1omET9CJ7Tyal9HZNqQaFRtjEXa4D5C3Uj4rZNUC9OwDKfWzZcB4w
QyXWRCzg3XGCf3WVRRGxr2O2ix/uTofkmwk52ZRa8Q57ONcnwSfVf2qxka/PIG24FUl+NeqmBZaH
fRsNRGbZH1S+MTiSn4JSjCf/SfkIGYzMA7afr98WNoH7OMWS6GyUjuufyqPpOde8QBM+CigiRzS8
aO0Lsu+BFulB4Ot+6THiSfVAQXLK1JiH/VnvZ08mNjjvMUPBuVFx5HcmbMo97liJGrc2FHLggbNr
DgmhMWroDbgscxHiTUxNZIIUyyZziu9Vw0gYelsfDtFT5/gVah9gqZi+wEObxd7/Rjb1QRvId/EF
bVBZoT5hnjsbOfJZnjnf4Iv7ryJ0oAp9h6rrMcHqEfvwqgkerYCJgGpAd8JJbwl3eTZuwOQym6bm
ezUeZIHWAY2GrbDz39AOpgnTHskcwxojEd3K/vWw7mri5MaLjLMvn09IJRP+ukdwQ4PUHyF3JJgN
F3qF7QXp7V7gsEI4ZlQRHfoLSuh+oTWj/3bINXUH87hL9NeMO4ZXTGkxMhbk9Z4rJUaphwPMyO5a
JUFeWcbRrqb8X12/24L2JHzJtIBg0Ue7mE9tiunNzZyLUEaWtJLXjWZo4GtefGYyTIlgMDvScIgh
mpUZoEo9b+BmRxT23fT7WD65WzD+qw5Iu6ofk09rV8PjLIk5B4Dt6WnGqaO9mx7s19c1Kk5Vy3XG
9BcRsTuz7xPmbgh8HcHgUs+t6+nBTfWeW+8+nKzJBpu7gd0gv2JyykRTQyXiFRLE+1qAcJFalAyT
CVswBifguKN/OkapBwowR4ZHofeaCN/OxY8v0zW8X71gUUwkOIpS8m0O0LE3eqB3ZgG2bfupdf00
lrOTqTwVD7V5ei/V3Be4s9+3lRnhe749U5RUOnvUcCgv9YPDeN56MsztnjrjI/k+ioLQJupvsYAg
Rzs7MrRHZsxdXS99HfCNiz/iTgvhyWOQWynE59odH6pFa1+PFZNcdtLYcAVjNd7PHy3yppNlDX9u
YvOfDzTpYTNzgdU2vDCbeTrREZLBUKDAAdNWFoLKXbKFh1r0CJs82GdzkcBvmCkqJbW1qizXQl4i
6zzmZ8XK4i9EYNESIbc+v37gLCCbgzfu9HYEqE0iRfwf1dNdkwHG6cIVSFBthiWdx58LzUpic07b
PshQQdQHCruheosc7PKBkgxVM8BgEIBQWx98GSU/L8js9h77LFq8qrHByKrzU3u+tfZebRkWz+1S
1z1KFSd2X7zgADXtkGodJL0Mt32kOmT4ieckubweXWJhjUl7HEMhf23wUtF3WVoCSIgGURZO4p0r
S58E7L1mOeJKwyq7+v6S1aC3wIxjFah7GZ/ABk8oXy4H5HyzydZCe1kcw4N9siiPuCWYsJt6eACF
SBRk2hUDkC6NyJnwjR73/MjstmVmhfktbieu4z6wUMxn5mGxOOgjMO49yQjvWT0HalcD89uPnbqg
HFXqUcAPDUUmMlwaHvRecex1uZplDkQ6QQgVW8s301wbZ6Kws3V0asha3ccoU9O5S+sz+hx0w9Ha
qx53kAUJOathKK9hZsxgdEW00PdHdvcKSHxuppxmQHk854f6OU1K8pLEMjNvL4m+5QSA/QQxwglp
42JBHonor8Y+Mqo6GmnzYXvKy/b/p6u2SCNenGPGG44deFRi6UUVwB0lPAbwx4/LI+5qBsnVfuAF
HHQKanAUdD11LIvZv1aRExMw3QNM+GNvt00S6kHaUaUSAGwCKyyCvsOG8UIczQadx3ZLep4jY2DA
YuaxMqpCX+VyCJ7OvO4Y1AU97q5VSDU2vwto3nUfCcZJBQV9nmC9T2H7o0ug+9F8ExQbKnVmZlKm
1Pw2BIjf7mIJaX/BQHjn3eeiQ3A9RNPbUHUJRF5gLBY77mKJdJKyZPLcXyc3ZGWu9gUynUNviyWZ
X83qtnfNUFQ2RsNTFG/HHjG5o1ZHZGUIShBSPznWf6rnB7DW5Ex1MZxi0KX+pqpcPz2qusIe9Mhv
tnTc8TOzZug+l4ofeK4zMinT3xy8lq5CbtqoGsLb3t0dC7zLdHETIT+pV7jXQ+bwAWkRs6fx5Hnp
pN44bVlKEkhRpCicz3ymrXlITkt81fs0+06WH5Ztv1UhIF4uUKp8YxljvAv75WV5XBu9VosUH68x
k8D4QvyD2iwJ0lONW5sLR6pxmeWjK/NNVPmsBCURwuqRTFj/y9cPW4f+BdZrnQVw5TJSyzjlM/Xx
qBVMlBEYanTIPSvflUXHr3CS9kMjZc2KBKWFJMCFqhwXNLU96l/9QbHvfvhBNf2PtBGMivhBhT7i
KZvRnRIi2OlJtqbV+gicWVDyNLDvL60mxoh5LRpRWWFsT+P4YyZHpqG2vEo9qk7oMR3zsGpuvyof
8Vk4xlCdo4dh56Nu7lQtAZaeTg21FI6H37oaNxhQyipoRId4lttTa66L7S1lu+6Hi/4nqEuIMujH
wXlrxthpD35MJ6oz91uwmEdFb2RorZ3G6hVVVdXEK1nNikug9e77UOOLNBNY00eRxj/T2YqBNblY
xfqyPCddZ2zHZOUAv/C7WIdQE6c6/ug5FHQvzLw11ry5Op58LNlxgqD5m5i2yhlWyZnL20TiCJs9
Qrd0s8rAvMrQkGR8sunWfQkHQDdFVxhELdmfkkBjiTsZggwbKyp3W+dENg645pIAueW9DTEHOKVL
NljB8vL5bScoc77NCV7RnO3eO1JtiQBxWzbcpk7trt2HT9b0PKQjyEp3T4/43Zfz6Z2BR6IV7IMz
zU+Ctj5lGhy8HPbHgFj8TR1ibGk0/T+ZBZ8DOhGV1TSivjHp4lCsRssXji4q/XeFtTMHiJjvm8iO
g0Qxrf/p/Szm2jMkNQbfPqYwNom9242hlmYi5PqpEk+e203mVxKXdokQxG60bdMxXI0TP1xqfT6a
iIBgoLSFIzb/GdeKXJTFf2LOW7Rs57msGYln6YgKQDRH6t9qWmld/8kQTbP9/495rXSp+ZhJkkKV
40OljoFazVuhQqFvIzJle+z2fEFVcRrwa478/WYpFZCxetr/RkHJxJIHd1mQV6wAFtYZWc+fHUB3
Jbnrb9UHcNtZZyzIbaIte8nzloUT3uIkasKs71ryZxO9TUGUV7dQ/6Z8aUt9aOPsIYPENMuxlyAZ
d1JnvOJYIEwmgtssZKlXMfe5o0op+z6skvN3nK6wny/sGHi9wpLdUeERzDmGNly5mQFTzp5mr+Fv
W8iGEAkPuwelV8+BLsF4XdHKASTk8bhT+LmE9EpB3uo9NBlh+3N9ESKQ1JLGnVjvIYldT24GTAIa
R2eYgNWu38kKhkicalAcaj29IxDFGsY4SgR4x0DWt0SgZ5YjLNimOR+6MZ6muwcnaHmPrdxAsHwD
9gaws3i0ET6Cs2NHvMV92mnNNjOxkToEVQaq/5vc9hOib/L9I0NUw6BlHV6mSIjQevAK5X3ZgANo
ckdn46/3yvf5nJdAU3zFqjiCHWLIcG9v9Q2eUSDS9HgChwCLJmPpgkZ2O8vPYT66Uu3wHFDaAQpt
dI1k3GLfYywFm7Ofc8Y1IBTwKDRav/sxFCdWsAunx5rk+2rtWk1NiU6QZEwixl6312NuMbB9pa9v
DO+OjzfI327VHTenE3RAYah4JYeD4ItnVxrjThusFI0/hGGWfArON37rSzAsHI/OK8dn9kE7gpQ2
QoaRGa5pQFBfskSt81ph6VVuWmBOM0ETrR9cGTlieCTCWAoMWVxNap5gpMdszQUdSjRl49N3gUpi
SI7D7jhiHAqCxEf5yaROzlMBRghsgXOTDdWyLG8hgAt08hTHCwB4Spgocizo0jOzuwTzohk2ghG0
4L6tfM0gb0zHEuhtU/a5ojmv8tabzA7FWs674wodiqOBIXVV4xSmeAfZUXj4XLKD6rIceqopReDa
7AubeZ830Cn0qMo3aZcHRi2TtnMr54N1OKOUzVpUaWRT2QrJjyQiimmhqsuHs+NEHiRY84YFiXPv
HnePff17MY6a0QnCoghWLBnSX2zckVwo2m24WHKHKVKDhi4+jfzTVtLOQAQt63GzY95ewuv8Y9DD
yBieygLwDeVLMS/lO7dDoANdnOJ2lUXU/h7BvRndLHytMO0CpvJVnsFsSPO+JR91sE1iQaIUaJ/H
ajnqMpnQar3rTNk+Jt1JTzaP07SNzi/nt6w03hRrn8Pa9WwYokmlzeVdxoq1Cq+tFjEAjpvvJ5VX
l3vyQGvRdRxgySdBwexs02eK98spYN9XfBzKizttd2m04U08FkmFsz7gHB9rUKXompu/aicrH3Hk
d9AUpdZtEi3r90R9m1TBYiiVI8Q7au/tnjROlKXjbkx1MFcWWboq+4Bm1V24S63inabo2b3KgKQ5
n82KIzAaaeJdoe/xBqnYFL4Gq2pnI/yer/iXplW81TFpqQCTMh9uQhVhzSFLmlgClO5YKkIYiW6P
o/7mfLz6xWmrOG4XyHCiucflXDup3Cwdwx/jh2UPpz9OEAXz938S+5glzVeHlg79RfbeyF9PPwzO
teqWAYNB44gwwQdYc9VN61lmBVLZ4v6d3DoJ2X4ulWqZKN4ZpDF/yMLRGunMfVtX0tn0AK2Cihoy
WALM6be1ABwCcuW6ZAULhXxE74EuthB3DJjeCzM010GOC9Tcd8w65DUc1O2ttgQbVlMeOWQETUt1
cfTi6cQrvbTxnbeV5+9SffYyUSk2OwHLbY0PWWGwPbAp3lz0AugfYeVn12snlBBLUFLY1OmWE/JE
kmeuglhPGZk2Kq9Zi7QuY3b2nbdcUd5r4zjak9zmrQmjOahoNzjLCPM0kchbTUEqlOnnW+ENouXr
ZG6NfNqmhhXiEUtLq69O/ExQ73amDHMZrWBCbQAiq+zEkHqLdCoeZcQimU9R15O31w0JFjkcKCwd
3m07YVMrem/sVBDWJ7LMSEG9NIRG19ucM8rC6H+R98jeYWuAYYILXERIM9RSiEfcmpzSHplwRcFx
OVRGRlY7ZjR8sGbWsN5NIBKm0YBdrFbY/tbDiPvUPIKszuYMcJRCnfdzxL1ylYpClTFGUk0ihoH0
/EfA8GEArh/6qH1yQi8QWc/9BC8JBEipmEXgl+UbiBpPD95IMwIgsdG4+ku4/uyrY0D9Jhy5WVYr
GuhnTXrLNl+FhJJHI+vr0EsdvWU8URRg0bunMX3L9SrMvV8OfLTj+eIKyxb4ez17X0DENAqIIgf9
RciiubZm32inNNlJ1geivR7Zblp66wLaaPUYFIKvx4Q6PDqGHsuzkoNSdtzvx77S75mGm54CFp0P
AMTLW7e4p0OAmBKp4XklATHPAcIoNpAAYUBithnLWxxus3WJuyNmQHsuoIBLM230B5SN0M0fGlsm
5RlsHuXBdvvBq4/I22A58eL7vvB8t4RLs6ITVEKEoYse6FtI78qTYQGfn7kKKNk4GD8Zi+wCcvMW
EJYDjti6VpipUYHWPbpfMWr0mt/spI/QxI7nOyTGN7MYhV1p3Lb2nWEt3ZglMisrh47ScKavB72h
txrXGsLHi/KkNkuXpiSRk8GHQ1buP+uoPUlSoHYf7PTGz2EBAI/guZD0l4ZtQFntz2owJn3II2p0
rbILF36kOUF9eQWw/C5E3xYvOu/KuuCFHJvuEjP+GdAg48HzvVTTGmKUYMRMlZs2jVIG1rh8jopS
XMn8zIK+dK3Rd7FKp8E5iWDvTzW/1RWxWjzo93J61iWDwY8GLsebQR/zkaoir1RFAYmDcMJqwhE9
CJnrwaWzu0qY6QJ77pafLfy3tYCNmPZ2WpfCV7dSO62EfjV672x240BzzEm/PnYuF3jhJFM1f+Ub
51p33iUR7Pxu6GokVTcUMnCXQ3/21bFLt2v9k/LmoeyHUQ6Xj+2uS8wRAsV/1uv4hVjp3Mz8UQ3R
CR5ZsB5a4QpueizmxPlmUHPfbcjUYlr+DELik1iNzoeIRX2dAcjfLhucRybLBg0qtepcN8tYaE+t
NhxgUY0zBv+NoGres8fzaydpuAMeFe1nbYZu82CholAEUDxmfkdYoZI1xj2zKxyOfGwsnU9r7FvG
3oHNzFZNbXK8QmDET9rIi41von75rWO/rKFA8VGv0UDYoiszUv1HaBC8KM8V/1+OU5LyuUtYNCBT
O/R8A+FsK80cKF1Q9vj9ZsYGPqFIgCFCVI7NrckkbqeNf1ihShbF7g/mB4i5Ai68hYfp3lKYtMfi
2Eg0+/SK1oEL+BC5ozp1JpHxsl7BJUnwU8kX8ym2gtW4AJP1v1qo9e07QPOEEN3R1nyjWVdZwHuS
12TEdqhzFcZHAOc7pATmf5aEKROQFGwQ4ZdTPOepKSiZXVm0SviRF28OOx1rBcP78d0JVAZ1ZZcM
J6LEEr5+clKdKoVfdP0g2DK0u6N8ZgMtcFgS/AtoHp018I720VaVrRrByqUBWANjiKGA2Z7u6Ltu
vmFJUQbmAjdspwpgQjMSMgyar5krBwQR/BIkg9p6e4dUbSM/uIIvSmmWUL2TZu2DsVv12gotq+AQ
U3aCUyM2jrlbEeyqR4A11JE4HTUOyTPHVXpRz0WG9dy+9Ghf54Jwq0WnfY6uT6RIfTBvOxYbhwaN
Z0g817Xa2Ulx6vdljbBPymriq3QJV1S2KJY5in67BybtLmY/8ion5xeC7BjbnEPssS3a2o/D6ZSo
GxkRUYKbe+SfRHH8Ub+ZBROxmpR6CCESAC+K8F9dxpGXA8hMXaGdCl+DWs/cKucrPmaz4y6evvpK
Kcg07/+qeq3fceIltQMSvm+hTvJUa9mX+9/reEVzr0cXPZLhLXNiVwz28KWl9R7AyVbtlvOR/lt0
kUJCJ4hNxNkNfr8JgygNH2c9VSv1XVCn/E54yYDsp2e9/T+oknb+XNKGXQa/pZQ2B+/ymLS4FLeQ
GXZFj2p/rnTcJwUniDI1NBAfRgUw+kZWU1WgkwB1W63OaZ+/ASHgxiBbQgaNX5/r9zHlrzC2TKcq
18wHXDyUnwfbvO23BVTl+PWrIxRf2KxcvrYhEI3hfA3BEkZ8Ax6g5MweFGin9k54qCFtNKRa55IO
RReMCalQc0LhD3G43TTnPfhYN0x/hkL4BHuvmt3ktz30gX3PZi6Rq3Bn6Svd/uQOB5lGFbXYfs8Y
RrqYgtFF5RqZVKox+38j122KjEsDZ9qrRKzHTaD+1GynuT8PMuOuRQmMD8b6d8vVsop4csB9d/jq
jxZ5rBeESqrWKgS6ilz6AczHj110qy21TYoWPGPt9di4sSqbMp1SLGFf8bLHH6rehD3WeahyIoSh
XyXoNelcgtp6l7/VhUEpIrkFp9doPkV/tdCfukQcRjYZxXr0K1SkaDaSImDsU11YGezy7tXYIt3L
kIo7TRMHKImuYi+PmdLHVPLn82i+TYAHnewGlesRMpTvCr5sV/82ZtoMfVBqfZGAr25EdWpFOEHo
8wey228wQ89vB1PnKkD6ieW8X3w+BPjSi5X0t4XH7h65aJnWqzbDO88ZMh1CqJQrDEeRAx6pNmZA
+OhVdPOr4g1dF7rspEAZQJKbPt5Jy4Wad0IjFutw+2/clQ1pdVKEiFJXZJsT/m5R22AnU1th0oRk
C7nSJPV1f4EBM2dL0P9C5aBMNV8bRexVW68y5yHq0lAy9wJj5mPxBXmVg1MIsoQuC7bKhC4Y6USN
30L2DmmClc/pCIyMpZ6UrWhZqhznS2AsPWc7RHn85mSUC1O+D+pvU5owKeyN/pF7p3c0Uq+vAPSi
XEw6xW469TkRgTFNPG0WYRrYhjNTD3vMI7mFkDzXXnfVdoEc/qF50L6tWEPymNl9q4b4AmJaFbzU
WoG/cafZsheTPp+V80n7MDVAUQkaxefVVawNSTawxavaCmaPYe0YtoxEwbTBhwo5qLSPD65rqwZv
t41yCI2qUDum7Xdq5N858eVIXoNc969ihTlrprqp9zqj/NyJRLJWrM86AOPMGYHL7J067xQztmTR
ybyN/mY6NoqbE+oBMgVBo1w8J3JwCQ28M/XiJdK5r8cRRPL06MODH1RAZ+c/bCArqQxeZyTbkxyl
7CMbTUHyx05NxixKOTGCoSJ6EbmThdoN/+oRFBhHu5yLyq14RIavyHEFN8hc8uyinU5krLajiU/5
dLo5hUqi0Is3J58PjlsS/YdNE0drUvQyUqA8C79uf1HIvE8HpDV7lwtFGAtQsVlF2/OWyKFCBjDI
GwW8ulRvTXaBx37VeU5+ygU5KNTtlbkCq1HDnOCU2zNojYvFyIQh+0332Jq9KM+PStEFZLmYZbZ5
0l130YrrXD3LKMhCoBTUWwZwY/lwSIzVSz0xPi3IOnb22kWBYNwV2GPyEUMPHPCyql/qpyuF+cgs
BC86DBOqAAnhE3yGoPAeKkZucJRrEeLmtE8irigh55S4nm3nlwHE0tNsi2/HthLDWWmUNQ43Vbzk
oeYEFHEui93pa1iFRPN47Q+dnWM7SYV5PuBLtBdPYxjzbIDUImRoZKC2wbxxFpLxkD5m5G9Yyemh
G/JuLjGX2WzZOp4YtlPFSvxNb8nN8ZQmSgb9llraJNpxeiXn6OemKPeQsurgqbNHFtmyYlOueflJ
w0Qqw5emTlh6+4LqWQtAFkEzamaFH26dxWPYbjEup7HDspMDh3Y5yg9p2FhoXCMzyTyxCjjNJaId
j54mmL1oSRgYOt26173FZmTV0u5CHj+5rS38oHG3sqQHIFbosyyeo+0hUN5/Dp+t4JAOovCFFYTm
tO1RngkehAQr9KTFIMHlI/tQXry5dNTvbVZX46mOQxSu2Gfcj3VJOAUmyrwjbThOgIZvDQ/e++S+
2wREAGniEg+ciaf1nU/0sVdOvwCZCj8AL6jEzN5B0rBkf60uZs5RjMl2PAzLhnSkPWGHIMAocIU/
l8UqTrLzYO24CYXb4u1SYTRMAKqK7GbSTsycyhjc7g009FC4r5Uz89vij7zplhJbLQQPn+Y8zB96
vypVshKQeyx71To6HZ9zIe1n3cipJH2+zhqJE+iiqyprC8lI8gC5nbli3xYwJG1oq4YiN1y4UctC
XydUuihnqGZA5wFsdamAlx2GMbWTSKgqhwvvtnq5t927f31EsKtxGi3jwRz0wdw3BFVYHXreRPee
z69XUNuaXnt0l91i3P31e6gzY8BPI2C2ZJoJwslgivlcgA3jJ8m+Y6LA+AumtmZBcwxDDF/2DzVL
oucKpeEK8z+nbGB0FePKkeFnAkRHH4sZdYkh7J8NugYShaROJ/JgEl4T5P5gJRrttZdtrE8oxv/1
JsxlYlKK0IypSiOgOKJiG8DmDJ7yiHOz2Y65erUzpZN7ZeuxZoUxFRxqzgMI6397BqOk186MFYbX
hguj+Pmlqfx/57sNgM6YoHN7YgxaoMVo4JS/HAiuko8XewwsmTtmV2G5aP8oJdMEWRUIDksRwzLE
05zYgQo5oTUZ4lnvdYrAJWav48N7bfavsPi7wseaUQEIvnInc4g7jXXiWM8dBEMbeTUxrPc6ykVX
iwrtU3xrZ6pgZ1tIuYAWf/tSj5zC9En/xJzbup4YAh0iuToe52OB74ImytTpD1hM0O1aR/mma9ul
XRF7XUuzGb/9zeLzQ8q72l12jrOcQnBJ7E3LW1aZRZn617BuD/XgRdvgiilRfYgqzAZSqzm9K4Ei
vMu1qFIdZ7GFPpqpJxWeMoPDpijh+mTPrIEgZc7HlEeop3keAw12dp+aNZ+8eUlGUMUmtpwFDmjR
dX2iJGekx7DSfeg7ylmXjimI6T+B1KDNRjSOdhOjlgdf+kPld9z/D7zP6uXdk7MhRz4D4kPSUU/A
7TjgP6SxQYDOeKbmvtrg4JEAT6gmHP+Awg0wjhKhza78bjbvGhTuwmNv0/qU8fldwNbUL1W3Rm/M
ZtJFezB2BSsPPBfv0xFrlF+dO5HuQ3kwvRqRBEdo5Lb3Ly9ufjPlD1DAzBxUIh8joFTq6c4htBU4
qSOub9R+laB+CZdvKiB6KcveF6E0A6BW/2RkrQ3EjuRI6bXxBF0kCdklzQUsQYfbT1xwu3oH5JKU
LBr3SriwrKpVePDHNxmUqzIJ7zlmoBre58ki7IrINukKeH52wg+BewS5LrH5KGtgSI1oX4JlTIfm
Fbkpe3lEXA+5IUOpjM41WMmt8bx8PPJ3Q4CXg1/M8DI3pplY1x/LZ4igea6xV7ArO2Q1c+5B7ZKT
hSM4EcTrH6G4eCwvwiHV/3dQ+O/b8PGu3rf/JO4yyE67Yn8YbX6hKAiYG9wsQx3gnUhWhKP6Hy00
Zcn8JVT7JFBn5LJNzZarbH59nhAQZdvg8W/4gxIGfrG6EEFr2CCrmAI9kBxaBU3X+S05f2i8539H
Mu2VpQtukmQkOEwLJbtN/tGdFZYgrGFXAy0COcpmwHo1Oh5Pw+TXHVNO/v34WMLlGR7e+I3vPaai
vZbWM2vzZX8+JOdSp9yzrKD0rHSLPtdHBeH+gLlnnu++hCEvqA97esMfH6HAAzJ4I+M1zz1GLvoZ
7FD7ztedCEPFU/6G2evG64Lam7DSNIrGaA7iqUEiq2CsEYhnP8Atm/BbQCQCQzrJEi4285dzXaz4
0uwOKwhiyKzjUAXMZZduvdrLwQokJ3LW+8kvRj+lk2qq+y0uFGujli4CbXE3cfB/L0H5JiAgPAL+
q4s5fGGAcRVyNNltEpy2nrqYk6vWqK8ieC2E0+fZekSZ78T8vSge5JbBF8W8xZqD8r/MJnMwjPML
4WqRAyOCmQKFqH5tPy10DT916cnv1iAYZaAHiCs54bQDSY/pTaH4fmj993s2Fkzsyc2tEc7fac+c
hC6MWkgtllHxuL9Fsx2sU5hz/x3Pce6Wt9Z+iSVWTUFkx7WTQptki7/gl90Xa5C6cyjji6WBqw8C
DvsTYSZ66Pn6BWH/G2UmS0tXpSk4jLRN5oPcFozR1oZAWOuhCBvuVXI5OIr3RHjILmkzqRX6MNjk
Wu9SQx4LnVmLu+RapFVM3HfAaaY2vq+H7EULY50myPFwCEvE40Ofhtyp+8o2nOcBdLi57BAKqV9y
AKO58N7jMYDWFkm/AQFRFulsp1JwM5MkSZ0UAGFCmOvSyI/N9x6YEGHXDN9K1g0bYgs1uekNXaUP
UWXcEF0c23yN0z9KhALiF5mi3ndYfUvrQfpxMq67oOSogjVUdq2bbCMDEjT3PxJfGA3fE/GOtzOY
pq7pC5TQSSecpk01nXegUsCNIgW6G2NS59i0gAjgXM+5lUiJIcpXZnhMnPE9tUNiLMyhnfgGMaYK
ch164u0ZmRQ4nRiZtbWtCioDFl5N/VDyky4YDXD+KabOET0cxVWyTl8hMg9x5LKK5Wn8IusrRIVH
iuFgFHn6HUzI0ZwJSNmzoGN/M0apt+VIHeWwluFVFVZIBCNVybL0gyX6ewemRg05SNU0IHmezDfD
STCXpv3Q7HOEQ/QGFAQbpLeAb1C9AD8Pln7OXCITSrNy9YJFOmTD+yR7FlvWpV4fa5+MzG/Lh67I
xtyqTo9PCOXHVo7bcO06KCDUppQMgg7ho/hetWx9pvGSuZEd6oZk+0gv0Tp/MSkSOC3p8pbXYxBC
fF/DeRsW/gFndFXbSy+AUx3kUzcZywVFVYjfGQHY9qQmvJeMcf8dFIzL8fPTvnhUUm7lTgMt5ThF
DKSDMxjkPKT/VmCvid0RhoEx1EEIZafdJehalLovJbbJ5LsnsigiCfZ/gonp8PouekHEhy4Rzssl
CLu42Nlk5Qfw3KHv2QZr04YBVIX0DhlQ5Ix0x7feNN359GfAlItIRt/6U+eku6368zpDdOJV1+TX
5OVMcW2B6noK8yQ+nb4MtdVE4GlSCRQNZpzVdqAGzmgMEGdoqrPyZLd0HDg1yb0tJixLOxYTvdl7
okf/8QfwmBlOHR4hVlUdnyKKXsinGMUALDgWAPQ9haz0L9TtMd90G0FVHrhgL9CHdNbUNCAtGM5u
ie11TKBHNqiJvoUbJue1/VpekoLUj3xfVaE/A3JVetl3gCau157e3/g+cIRaUVDhzn/RwmZmbkQE
9oEdklrEh61dotYwnEZeBiLcL3DJILV8/vhf1qxEi9qmHJO2FPjtHnbkksO72qaJUaUvP1lu1KCv
vQu8I5v+CGPlZMOCRo+C0qRG+BkOqXZ21sT1nGTvGl5HOvCHpf+JE3fnR80my64ofoa0d7qk1BI9
ShJGLKZmjopgO60di+SyOIna0D4Dfpegn2xL/vK6Yv/fHIfbcGDVV+T2Hs/EkFuSAA5/MWREOmeO
HvVQt90x+E4axoE/89BrF4yRDvkc0PShXU4L5VqHlY/BgDDHW16gRZ0k7t403DSS/J4TZHrK4VoQ
7UpEDmZsgfmEwRXtP6YpxQGx0n+oMX4CoGmThXbrqReqglQrKIpgt09FIXilBBMfAxtMDwjv7hn3
A97VUAxrlCqgdqgpIXtxqGKZx8SCozwpLldeZmlnFZdfNf09qFOvZoD1xfBP5kENEQ6Msjmo7CO+
KvIJ4nPJEqhUO9smbe629pOv+Li+uPC28+u7pSppyWBcIvvp8xYn9C6qE9bNP2IpoE5ygzI11XRB
mWIE0Rv1k0XEwVKZmeI1qEQpx90K5bTM79VsYtBvw6ysd/lk6GrfLmfR74iya9W40l+AsaoOX3wo
fowezhwdWO0OrFGjf/lugCvY5iUvJk6NMBxZIbyXWqmQLQtvgh41g6rIsPwyIerT5vneWncBDDq5
mIeE81E8n0c6LtCHFv7azwKxTdeBbFT56f79v8zQica4I73d64E7E/0Vg2kH9tSzldvww/pnHQBs
qZrOXnR2vEmysa0JK98EApwe5lTZf3yLe1HEjDvi2j6S8RdOtExEK75orp/xNkk7gTimKZl8WD99
b4HcytiPeMF7yunV8Y5+sOg8jOFIySQRB6bb+PtkMoEpIs4vvm8ORExr/DHYIKLrmJfgyB1abWeA
cgOHDzQcCSlkHm5svgGJb4Mib8UdVAqFG49DxB+bQ3gtR2Vm5Y86sc5xcIASQNbdmoFiT+3Gdw1s
U6M+tYnDSptMnVGYAmhhW0YfPuf08/7zRlMTxMAyreiOqFLtFSeFMzcnShxEP24XBuqkI7YcRde3
vjXaSloSt1sW/20PtEvwnFmLyBkAp/v1C+r2N5gTWfvZTWKjpitvMialVRslnMBM+40ZYGrq74aT
ZUdcsO8oFsgVz6gYsPV2hmeogpareeoMxcMhUlpddSZK2j8kEwm1z+pvKhRfX7Yk6cjfk+0zqeBD
6CMwnt9tICQP2VbB5Jn4Zzk0Nt6LPrsEuypV2zgudfGeTpL2IXugCNEGYeqWyUin/KUtcYzurGEU
OOPhaxO2yof2+ygD0LvxCCrvJZOT4yjTDbqQqpgW4nK2Z9OlJ+YJaFEUjimix2Ccy3B3G3wIhwR6
hYnUoTmF2m0CjOsta/aeNT6lcfxLVYBjcxrtpnwFp1shO4wHrhVnYQquKsiiUz1LGkW03fUVciov
X0vz36/aOyzajnY7bUdXJDOhv+rLaQ8GG2AghHw9ejwK+pzppWA/JRtpJV/L5H9/+uFpFkvECJAs
1rWlvCFp/X5EVY3QUyP8rQ+MXpNMhm+AjqelcGOrKjxf1kid/JVDoJXvFI0gMu5UGjJZFquacqzN
2kWL5Uo9KvGRdr7muU6VMoFL+DAIeMZpy8PIYTR6aujn3SeuQS2cJUqpGOTXHxBxzgmM9ACCUW/O
XvMnQ4Ef6jW7s+T0HH/GuuBa3WId7ooiNflC/gMOkfgUUOdQxQ3PVFO5qDl+31rXS5K5xwm2gM+0
90qsveZsAyfweVw+n7ohynWiV0CspGtx0dBYRSN26FqSXjVlPnEHiCil4CDnhC5cxhyN7nHlJNOA
ij6rlfbFqV8MOlRqE5r9BHLxhDQboF3iTNuPm2BLl3tMNp/0gcvYj5A8UdE24od8WoiTV5Y6iEsO
9YniPM69uzIrOTR75h8bzZp+43WdjvDa1JhlkKJpy0WMhPp7ghBozwKhJZZ7ioWkPb1CKcHjES1O
Tq966Q8bh9tEemXH2nk5Op0VDwTOFAZeuwez/JD9RM9TSsVxSeITEJ1gnR2KJ11wuEd6crmMflpg
x9qFvjuspemlt96trmd7VOSYhWDtwxSl7+l2rRfM8CYmto5tZVWkd/xNBd1UvniUHTjQxhOq1v45
HrbK38bszVlDVb8tpLWpFjg/lZJlG+fTTol/Mpu8kKcxYhuoBMo9+2UoogHC4/w6M1Yt4CVT08Em
r5UOB7o34Bwi1sEP2LJ3whinL0TlX2uRlhsE2yCGgRfZ9+I1OgIps1m99fXyYb9NzsozrlFGeUhV
pcGSITbaZPVoPNmwS/qxfyfbzn6+Gd5v/lrU3KkeW/6z2HSup4RHs68DdRUTWBSxjAhb1fJcbNTx
CCnb9gXLdv4RjQyBAa1nNDNkWT91ybwPhhsMyllks89y6HjoioWHZJ7CJJsaAl3n1QFR7INGFh3f
/CDqFOouSM5AQAxA/4ZhpXf7S8MAIreGAvlDevJYEfm8AzEMyUHjn5bOBE5iWaMDo9ZaHi7npvqQ
czljG8NoLc0PfKZzxoAqdMhFGIPWxk2DhekUt/MAW/KFpKVN4Xj+Rlw6xCCUzh44WGNcWRNH0Y7Q
Trb2rzB1D4jZQtnH2quicl7rxy9NfPkv9lRpZELXoYMCvETqnD9rj+GwY0Sj8u0L9GV8RWigMsmR
tARdaKqzDEIMrT2P9OOpbb3V+nCaf6ko0oWwdvOwdj/9ggq1EC4y5H+1ghctkDNLpyRNvFktmLgL
J5CrgGHcDm86vx8c0l4uv92yXgq6aGQfyzfRBcjFkgAY7B3QAOb3dlCND6ZcDXN2mDdbQVmnEUlK
pMmqJa2D28cm1s8wUQkHrHXLzeECR6ZfgXsNmnZwAx/iD92y8xHkMuGxHQ2QaeZojkSheVSTUdhJ
egJQtlJXTtONmMA/kTWwdN6fB3MCXajMlxmADKW0HY006WLSb0ORaL+GzqQ8FPf4X9KgKTDXKQkJ
v3gqLm5c91/bFFZ1Tke8fL7l0iC8tU/PeyVg0I2jUNUib8wJjB+tCr5BPDuT1iYCd5F8eWjPUhUt
mzAF3alsJRRCMYDkm2nvnxt/GOHc4pCF8jzVJX3TE9OYM80udKiOWPRLEIpL5J2PtaRoimgY9497
jqMnSffWbGXREKWnpR641+YLXUIFyeV8xqZ3LRClOLgPZ057rVYpCmFXtOH+ypAVD1nRGCHpp38H
S9lRMIiCtIcmkuQEve84dj1vLOQ2lFdzVuO7m5fM5ZIDg7XU83f7F+Th68LHX7pQDaA28njLFYvE
jfZBkigNxAhWT+zgo90+WLijRctD24CQLaLOuAiUKU8dQYzwgIicerDNPk3NNZzTxoniaaHKOL5X
NSeg0EUWYGW/Tm2wn5Z+uJ7fGxS6TdLaE0aiHEpZmzBaviiIoe15NcZ7Kb96dOszEDV5ZWIp3WK/
RF01KKXuphrEvvrSF5D+I3Dz6NovJ5lvaUPSKVDRKNgcuTQdEJhTZiqmb/3/q+s9no+BE041iLGf
IWsfU7dfVg5wKaFuqzjD+dg03b7ZQVbVyj0PsoeQEUiITtbdw/SlMigN7547r37OjHJO1g96IcvM
gAKAJs16f0RVgIvDgQVfW+Texd7wSfd1PPVEbktZ5SydKqMjmbFKT8fafsxkH4ymE//nOGlf0hcX
tMtOMS+dHzzMSyFk8nYE69XWScKeM2IsFfjPcl0G++RyntDRs/YkQ5Q2xRiUrrr6RlTvL4PZ4Wz5
hqq5CZlpRYPdi+aZIUOh/zD4MbIAd3YgSR19WOaQ1yBQpUSb8hIIkWFLTbiLcgAvqwtu8uHh2jF6
0rbM2UW37u1K8Lf27lPc3pcvGSEf+yJL8lWfC+ypjcW47z4lryIo8Yo+H0NpmJ1LKFl1RSeMaDMj
qLBiDv0jcGZaiY5/0SKhJUDOOPOfF7oQUXQCoYdUJhsTdC5nfmGWEDXITgqWUZQLjortuJUo/D9P
VTesrf7KagRLu0PRL8ZZy+HuVxGiYiE2ToLXU/+IHhtoAwzi3KnmEJKeiYYY9Cn4ypwPiOVYzpkC
/j9yJvveLmA2ablAeA7vKwrpvkXRdsq4GgSUUuLraCqgJ6EfRZcrVw5X1YEPw7X7vJvxwwRacE+E
euppqjk9MhPb2K2Ch+8+Z+9ct4swjakWa4q4AqTE+ydu3um2NykmnenyZudA+hpeV0I4HVXpmrcs
v8m/HV27UIQbo3tul8OuqcZVi73LJO0zdPvXu1BfJVN0TPoz/sY6ZMNqm/Gr9eiIk/ZDA09JfR7Q
KUXRdH607ZSR4wAbvL1QA6gc7sRj3rTQZgoWILFN9AvlUFscOBrqCzqTfSA2g6Ud40u8ON3Eao6j
tGUHTFchZUFsqgJrYjfqyL0o0robwTEie/LufCMCizT7Z0rl81xLQtW1l3VUjgawynu6Uj+MupGz
8ey/ulJU4Kl3psjxp6VJcAnr3KtD9dLbIocGNvdfZFxZwnL647IZQiuXeWyUaeLcA6qhIbf5ncpT
GLOHMSuOc/x/L/unu3Te9O1BFFS8PPJWXOe68ER7hO0MVHu5i8H3fyBnGqydGO2Z6fz/e7P3NNRt
CbPi7vM4I8B0+UzcIAX45B1DtZ0grFXojaIX8pdG1By/i4V6ipJgndewqV4O1hZg9fENaTayqxf2
Uu4S5FF/wSogfjsKPl8/XQd9xCkmTtVwqiOy45j3eX9UoPG2M1QIWtmnm/dfh2EKYdup4h/IIMs0
zIEGcmfJTNEQZS4hd78hIqPLanFl1BqKRjke1W8g8sVSdTK/jT67wnddz08LFmPoieyD2fsnt8nr
XtNMC3ZWL6zWV8/OdncnobXzdwCZzHIkRrPM410AtX9NEIFG04owiuZCDeRlbSCZ1iuGEg0d6Poq
r4Yy7ihb3ZLZaKpfUCime6odOTLxpvI/9kQgMIneb70YRdsxeLk8FE4CVj45f48L2BoGxNicmmP0
dNPNOWcsJ/2qVPWGaoG+ssOK7aoJoGRulG+RkXVS7mNDjBnq22QRz+fcpls8R+eH20asnOHbhlpg
JIOpNyJOiJQptSVfaSFtf6l+rYboF1FjaNPzeW3PkuQlq54+2QDB2U4V1fPLcT5b+PKpuXg148XB
6ijf3eJ37zkoX45cfbztWgbN5e1kC4Q2NyyEeLERc/5QiJZi+sMUlwTyTNCGB+5jDWd5fuSlIdJH
+SnxFuiBC9MA/Kazo6np8Hm8Be82eu/XKoZUwZg9HyqxvQRarPtXgACnGlYL1zxjE3K644+mVgGd
xXRDAWKYo9B//qHJcfHVflqpO6ifnMO+tyM6hHy13+WA1rR9nqa0muq5jFVg7IFyH2QBixyP4WK/
lFQy6kJm3HRscC+I0WgvLTJzJiEYgYbDJQt1U6WFHz187nVZRJN4fcQkUuY8Led3Ud2G0kqVo+1d
npBNRy3NfbOpSs0v7uA+RCZkXCpHMyFCuEtZbNi07b+BUyNEz9v3kqoJ+AKDyNkUZivdcrifYvk4
X8J90Yqa5i2X8iViUDNMfqGUez8gYGzMuNCI7yNl+w95R/duEO+8K/Ldqil2teoT42myaCqSkkZU
UpBZAfgJOc8v4mlYmuUypc+3VJLFiD3PpaVzVs43UyD7zH1CsJH61dqHh59wWtDgbkv++1LtBfuB
ZmqgOo6wKwAi/cR/qsq6Erivh8LuS/Z7YceZVT+gCOQLhKA4VPWniFfDRNLPVdeT7XgXv+DF7mU5
x87XiAIVGjN2+WkcUtXoKIzGAPiNp602EmKMcJbwbBw65tEDic6tYQkjzHPFH2zU+VhbC3/aOuG4
Ot0zy1dNH0DODB3+LI1PvLENE4SSmcL+S3HoKuNX/KlAC5uk+5Ql3Kt0wNVsmRlJyb6w7p0Qkp8m
wF2PPfLjL7I2GrCizJttGqfCsTp4sgtTLYVmfdVaGpWbR3oxwngIpOhiSu+1z33QKi1gYYk1TisY
A913Rusg49HPo+zw0j5mvFgLXo2OZIxSpdwvXcbXDf6KMLTnWPhAlN1RbTcORPkfx/2c9EzL3qAg
aPw6vCw2xjcezyt2+HuKZOLi7X+XvdRJl0Vij1x1rDxkWlml4udEKXlmFxF9ZWqd1yaBd2g9jnd9
O9lza2TKGybYEBhWFh/CtHDS+8thMQrll/Tl+NSMeA7sbDPLZo50qsk73IAqAPvRw+kO29UcMe+4
Ga9Jka34NzUlj25zYLdjqAJ6yt+jaeOKoP4SGe+uzMMgzg4yciTynsj7/FGBqgBW/zsSH+Tkl07f
sGJ2AVr6SVWsSschbFamRDHhkTuoprP/FiUw14GuPajo7eHxENQHU6ib6XyW8KMulT3ULtw+OcIz
GnUzE9Uh2eq79Rsg79Wi3zU7iTuvgN5nlXqqkSjvUgWas/+7r/t+HHlIteTfL8IO4skW0jueFpxO
lx+wYUnngBY1/h4b0l7yJC6x/AX5f8uMqrQoNEa6GpRWSD9EVQKNuTAh2lQUE5Yw26gE6vvJvBIi
JVeBuru5ua/lW61A5A8V06+ZEmk9/5VSKgS2Y9hHK1gjp+0j2ePV+pxfuNutRXM5ZUXAnnWcMfMh
aLUuVeuPG3R196SM/yTLJWsF+WqpLKvWLRGvlLK+ll2Sqt8Efp5sKGNqRUgENvSTB0/uk/kQsLf0
tBKVJV62vfKpJrdvKIzHBVkES/XxcZ2rb38ptR5rI1VcukN2JGLllHUgjQQGBo1tVwHFgdkij1AG
BRt/vi+QV+iyAUOUTpmqmpwU9HefaCTyB0b6S86tetDZIE4yyaA5CCRkpOOR4zwBRB7dlB1WjyC0
V3AJJuGfOxGneTHSN14KrG35PCBDrYmDLkVXxruzMs+Ovj9judvPWqzZX44qfjn61jIJrK275cq9
stNlgUHryFR71Xka72JU3x0vjNPJOrKJI8Ds3IA0fVF3oec0rSW4w7EtUomNJaDfE8wt4Xmq/nxA
V2GXfx4BFu7KYSQnZeCAHtFmjmq3nICdXpqDsMb2SN03+uWKYFwLiMBW0J0KbaK6LKg4GpEG9+tk
gGBYDk03ai/03C3NsprqQfoxKOmd2wIYCkCOdDSo1BrCAKN7ZO/eT/vzS54RQQwRagSB6wSCr92M
tBGefl7MUf8R7H+8LA6QesecnId3TQmzle0g6ITIP4VJCGOxFpRmmZu9Xthb4jiPFZh3mk6hqjbT
v3EF4klUEgjq6o2IfRmiy2Ld3ZMUuRnVZsHvupuA2VWl1E3SMXGsW+p6kj8/afWmmHpvtT9aQu+k
vMFQlwkMIpzmLRBhVaapxvmFEcfsJ8XRLnjSpVkOhX9FpRATNs4/DucmNScHrgWUQgXA/iWu3xDC
F5gm1Sn/LIi6Hbo1AhH44kLtE2qnkGgL5+jB0S3Ag1NwtuCjOxl5788OhlTiQtK2cef3SZM6tnxT
vvVZp4pgSPiuM5608+O0anY5AQWS4e2LboJCJzOpWQbmC5LJj3h7X0++XnG4EcDzf1TAO74eM/+W
FjZBqNdKGFpwuOtooBBohRKvzFynr6tEJ/yG2IIkp38yUC8aq+lyKmNLr3tToYe1eoOcJs9obIk0
QjCTkAnPq6VfOexVMUiexp0KPYPBP4jjnR54vSCUQi4oLVt/VyMQ93fowQgIj2vLXjA05lJ24Ph0
cQNajpmSnbqPjuBAAUi85E4xRYPihyms5EKScjqMyxkD4ttfSndCUPUVPBjQt1v9dbGDIDLLRYKK
AhWATnw7TL4XR4IB0dtFTqjW1W5YVJvooY0+WcbqTqeg3DGA2sSHwy9hn+aHIfhw05YXtEsuTtkK
bWIYUc415pzuRUfBCN9xlyADT9ZdsXca3rlIFOAteEyJ0wd+CP6H2I2L/PqQ9aN4QYxvRA79aol/
rRbAbRtjcOsinCElk9M6ZaE/8pSqJvDRnH4ZpD4Yvuw6/DzcwZZz7kNgwJBF99pJYuY3WmucHusD
9NftrHo2+LMGVueyMTaGBB3D1wmVeOEUyi+B9w7ajs3JD4qJW+exeoAjFVLFeXLPqCnOUNs4tZ4l
EnlYtlBnuyw4Bnk9nYhO3vXFeoLMr65ShcaIIL3ZtLyMexgEB8K3M6CioE6Yot3QcvHTcIIixP+H
BIP/gEpJxm/Nm4SZW4Z5874BT9WBPW3ZWhvTn0qaH519rAF93eR3FIFTcGo9/vzMybjWK40H0Sxd
Ovy8blzUP0raXEO642v+L0cmI8mffjIERIDIX2/NpHZJlaLwa9NbMDoIrbr3KUUrMLggUc1uFQjd
M+j40SUEJWgR9IB5QBJIBUp7j+UHnIiMZjjpomItRHbTfDRWf/YhhucYwJqPZP9Jkp0q6JIoZCt9
qve4af/8tfZfl3odffZUcqlcBSMucJn8fhCwhEIUmK8EkbPr1hOHQj4JyDccQNQC83B3KrerW8V1
1ktC4HT00Cn0QlZ2W2UTNjrAX4NeyYlPNE1beZ5TBrpE8EjDiOfYzzXEtg3U01qog2fFDEaDp+Qf
eoOwVy4+Zt8mr7mRpm5B5TGtZzEYkHGRcM4ddgdLJ/ZhyiY3ZC4tBK3Lyb/qDHjJYn44gq47w56f
vLOqzad4lp/dLZJZqykaHjSki71ao+SPX0Ksv7oyb3+0aLkFYCvipccHOULc8tbf3d3XX2Otc25U
3yi6ilL1QNjGPRiTZVyTzsg08ntbbIlBTLHZnTmw49u60andGC/h5/vB/UrCzS//mjiyhrDz+dE7
JPMXnUOl3WtpENlrgY6ET0ueMrqce6+y+9rcOk3B47ssNtoE/MggkLfDetsQvrsJd3KZGs77pus7
d+HhmgZSXycky7dUwvutFN72d52jpvWoN/fbBadK4sEJIWLrGVdy0Wln4t+LqsrZ4+8g59RgkaC6
snRdNo6xAOFqSIGZ/5OwIaeBqINVfTqB+gljZOTnTlsqUgys1BO422cqldW3g7baduCBndfjnCof
6XEk4eRZvHtoXVF38Ponh6owLaWPtOJtY7z/Kmc5/iaD5iYTxHBCf/4XllGPv9wRMGox2QJhXFMs
lPQyNdxLbUyzxIFdABnKF+7xWWtn7UnYyaK2KQQfHCtCdPxI2lOygbaPKGAFNNL3OmvjHmOMTL7D
bfqJGo4T5ASdrIhTU2W/RbOU03xBz4A3qOkNdryfPxcGWXjaRE2X7nVQxp3m4HOP5QZ/LEsarfLa
Lliym49NSQAsxmSc/0AyOFEj1ueOPWyQlPNPFv5etV3V/W6ZnmwfkLk0hWv85vYyGDN1GTGvYsLV
Gqkzh660/jLon2zUqzQjbvktyD51v1dCkqNzFZC29q8hJyT0qT4NdZmW1/Wdb9+rR9/nmOX2o0w0
5i5ifehWer+1/V3naFACTanBDqZhdXGIPoWleeikc6s+WIObbbZE6yt+8Ine2Wf+03ipYVmW0DnA
mysQRwZ1N2gjX1e9cq1bSMk8uOtKUvsdrbTscHYVuLyMXKrDK++SFzmyuJIU6129LglbLb/5dq54
tneVxj9Yt1qh6m8X5/aSg/+yd7VHJmH4sFCjWOdcsjOA6+d+z8eMuDtcYJqybHx+EDUA9ZJpVseM
XArx8bg8LnneO9tKZuu5b7WkTNn4vrw05L7E0tDh/EQmZi1f/H8vQwiLtYk3kPXdFsYNxrj7U5Zo
cr8r3etsnnlEhO188o4jX1j9ZMx699ljwka9Fo4vppj3OdDRQijJSawOEDVGFZ6fC8oOLmD8YE+/
JuQ80RWWqs3fA+wLJvR3Ecw3JZoKzRX4oSeDg9JenJwcfDXsZz9FO+gl+LQXQlwUebcArOaxr7XR
Y84V122JpqIw3nQcIE/5jcWtrkPV/4g0lSjnGdCEv0myYIRROb1UqGYmHwqrptobZO5ranez3OZZ
9+QjBTJEr3Kz8dBn79jpZQspYxUaLWeeNRHNGDmQvd54a0x7l6LPPBu7FKh9Z2Hz7M900BHJ6C5t
1SgNCx5vjH9Ir8dQP8Bvsgb51vTCrnGV3rfU4RFs8veV8GSuWl/jPMWWItaHV6hBNfk6RQMPVAQo
XAAUSSl/DreMkVInCNyBPPPA9xtN6U89ArSgckIZ244YEUIZQaK+37nOyNWlnzqPnl535PoV//l8
WATr+4XeWZECRQAcJFl4RFyLcg05BELjrvCVCUs2T3AzD+8UcG+GxXnMxbYL9JZ+gtnP3065uKhy
w/sFMTG7wKWkqEAg1/MrPKHrhXijKQYLFGt7aeFlaHH1jwdWpJp+3oeTBeJCdTFK8MbrEwRUhW8F
xRp+lxPezQzs+MOEfsoF/POTp9Ssz/EqF7uynUpmBpfNVfjARsNvtJHr2Yl0I/sIk6oFOBPh0O9y
SMJM8EEUbKkJI5s94eJLxv/m4kFMr7UQ6HgkpMTjwyz1trrzeiOcvKgzXGasu8O7BngGhF4sOBoY
f7aq31tR4oUAXWTx6GAldqtoTLAWDia/Ob9fn1TXJZ9oteRzVokPjFl0TaB2d6Xt3POuqpb0uljc
v/kqwpy/8qDFtxDh+PN9l5dQRKHAKH2IVfWIyAUDHUDTvOxG0JSMGUc8qKRhZsfH1X0i9IDZuqjt
ix/H6sBhiw3nXpkGYe6Fzk4r9F5F+Bs/i8D1mPwrsb5vPBOierDiNfRIsHH7UBwO9WQMkGwnL09M
LiAakGMwv53mSyxyv/mwdVGHEddsJOoo31blub6tfaHc/+URabrtBm8bfBzrH8wGLWBy2CnEmO9J
SJQ+30VOq67/gl9RnpjFlMOjb7bAAdCFboTCFE6oxRSrwUq5RHtWjtM0KXqDfMW2fY9lPc797k1i
W7dwc1S6g4KgOxhhL91vObEFXmhGeKFvSm9ouAHSlJhmIhtD1yQZ4XTqOTw3MjJrw/hUTTmNQ5+T
ja2s6d1v7cUI6kTb4KIyHwuwjIw6bRa/GZcDDx7g1o6mHXHuRV8ulvGxhTAPoaUZK/WEqiJO0u6h
0yZSmFL0zyvNlxSviu8r/pIOIpR4Z651JZt4iNQhmuTNjj7akkPaftl1A23aDl8QX17s4+VwBPe3
UqfkS41ZPmQwt3MV2NtpYOnVuAHIRRzkUgYiPNfkw8bsYWX8u1VrkK2W0HfJwQAMeL0342bdmkEF
+BsFb8WFvUpJyRynT3FJHdFSUO55W31U1vUAGwcv4dfsva3+EGrMB/BwiFD9N1Pyg7cpXqo0j5vF
5VASV160g9ZTaWfLc40v7I2NUFHzE1MLMK130T7ZPaqi3y01eZ1IG2Ft6gBnppwBk++VOA9xp1FI
FaSVtOgsw+QgUxMPZuCz0u6tDZB0eJk3veywJ+GzCVn195XD+VbI/5oKVxKxZFtO43RLGXRiNxvp
bJocUk4odjH3GoKofVdIfhm/lgmr2slizNXYtBKz6Trdoa+Ca0jds1cOn6M8X0S1LDWQ9TZctLO9
qchKfzwu90JaFif4Ms9cxcMkvsNl9VLVqFtp6feN/x81nJikXwf2sa8VE/mC8EGRh/VBWyDPSrXg
xzzkAMNq4KzqESmoC8UpXFV0KBGLFPi8blqGp6rXHHVMKHhljegr1519IXuMA4S9Vr3gWpKHngZr
cAQ0lVao41x81nZoSLOb45KhaghKe/D4MmPyx4sxqzi6VlKcQJOSGfmMsErW8gRNFC2WSQDUx8go
Vb+MCaCI0UmwcOfaYW1aGCnvosmCvLwiz1a49c1yI+mLdO3QHVIXtNYa1cjpn+r5A/srUUEi93f+
v4drk7Xr4gOxJcts9Im4h0pf1oljX7Q7ueIsJi/p59sHV0uFVOjDHN8aHPX7qMK61A6WJwPccfTV
y3+SgXC9TmdKuPNhbCWppyMTmp1L+mN8wNNn0BGd8YgbdhgCwK4rb7QNgAUCGK1PQZY+vdxypbxo
0AGUNWpCn/9v/OSAueurnLN6BelDs7N/VqUaQVikWB1bUvWeV+KmprKg5jWcGc9Xu6byVpMTBhNt
5Q9S3HWAHfEEZ8JUqBCXW4URpdtMOgcQVM6plIUu26VxVG88Gh/fvWqxOH9hxzxVlfTRJaljlJSV
V1cJZNE4n3vtI6RpGbbvihUb4oYquVJGBsxzOhB377MyTX3+EImKdYMv0ZjK/pjnavhSqpMllDv2
RduCikCxoQEaxbCR4Y5WS7LsZCyVVBOz1/uY/dML8NB5yTA/dbjWGIW5yRNcNk7vy8q974eDXI9O
2h+1nstoX0aApnj5Dsa2A4D5cmI5XGEUGwmyZ1SCcEOagJiIEkK6EE/LwTKPuQ3CgQwyaQxeW0OU
iKJE+WEOq5LUjUUKwrjJnDLgeLsyeolA2pU7jMhLMjU1M3uzHRsvOMsj3tX3wIDQtUTDtalDDs41
oDcFAALSXP/H1pu7mwbe7/PLtuQlgM44UIkohx1X8nViURYQtPvlBgS2tWOalARnp0w14eCzPjI9
ta3vcCXpwdZnIy2TZiMrwLi/MG35NUL4UawWPy8jqEEr3jDL7T+9kAn+Nx066tIDRiqhPGssbpOv
Hrsc1QjTey19bwoFziqGFwE/guIOyL2AR8gJqS5un3oCf4QKGu7ejLLrOVSlVRzdIneG4PdA1rXJ
cVSiiGoCZp1rfZlbEAu37w+L2P34GUTptxD5xzGA2AhbOHD7LJ+CFzRVq3ogDi1us7nTiE2k8g74
h+BhFWYV8d+DpsEV8ZakOV0c9arerOIx0WjWvIGgT+EE+fwrHkOzI4qK4s5y5z0sj5ksI40Fjejx
jXLSWpzqaSku/MUrJmzeEaItS9IsbNvcij54s3qTIvuyppZooFQYbiNW+twCsN+CAOfwPfU3nbOM
8Ne5TZYSA2uE8OegyKdjKPxKq4o44PdC68lSwsC447dq9+jpHR0626pKViixO6Sm/vYL09EIEK/1
Q1z1LQ0hxI5LnjIXVqCegVzhIvwll81SGVKdrjLurozXERE47CMuSZ8749KEOsf08trJiIRvg0gI
CqYEfH/7S9yHNxKg4dFcMqEumy8qBjURd6k37wnj/ZPcdG4Za4SnTImX0fBYR0ZgezpcbiwDseX/
N+EqMdJ0KhZlebltg3VxgUXxYNP2aSIoBuckixLfm897Oy0h0O8qGYRbW1U0A90rlzYDev8gRrHL
SQuHPX8oIR6Bufcjmoxcb5Wjjr9AR1mo1w2j7Duo0hUaUVmXo5TnsCrkjTfgeJzqSuIO7gI2RfZF
S4v6gfPZuZe2jhkqLdn9aY41qr9OyqR3uvMgjx9HRhlifGcge6PmNlBWrGs/PJXi5GBIT1LOaYCB
OZ/kuNQ4Ia1+ir5EAcSk+lYAXTkMFyYsZ2ZNOOWvd5b6G1gVrGf1F2wkN7CUGsOOn6JUEEhoFknH
YEAXg0mnAeN9BtcM/LrqAwE+XkzFhdhbeEVR7DxS7E0sZhNwMItn4JcahrKI7JjKdCrLDJ2DF0+4
/DLll2hhhf1KpZGg/GYxBNAQyeVXO5MwH3dUFNO0v9ONKcyDxlsnSvNwuCHbb7BKG7sJGMcZxXv5
RzFPOj1oHWjvnzpcRK9TTwwNfJuzU/V5/eS7GSl4pEPk+tc8fPIi1ufPk4ZGichQSNxAQIW0HJ8A
+KQFpYJO1nqbuMrZrAHd5H2hqSvgCbv8nMk1lt4sjeTXDE2KDXv8IZD1k5FoxbcRbruPdtAjvIED
qnSI/+wzlJ4yJPt5Q/zjQ8VIp0Jfd89P7t1A8cOGlx2CDHZpyCnTyGTOHlEcsCCpeWYAgMcDTaxX
+lSaLCUHONA8HHnM7OVlreZBP5TG+tsuS5Yq4LqfL6NUJtckUSI61FxEiyZS5vFMaIE5xvQ8MFJX
6m+uezAtesw7bDEakRq/q9gjsUVUR1zMq0mUbMHyS3MqxizISt0x4glKGjLpD2ZqkLgGzD1Vqifa
E3iC61OgProbUgbIKX880UZP/SUpPJ9lS3nOknDIfIsJK3w3Voz4YwSW7N+rMowLnfBG9yAmjIBN
h8sdKV6MRttFv5gLLHPK0CJqMazKvfywOmoqEvaLcR1TYZzk9z5LrHbhuux9XPiAgrBCs7srJE1Z
4E3qOU8N5wIK2eMY/klhrgGpZJuFe3QnUPKmxJ8lTVDsBM9If//zCGU44ZAStqja5xq0mxUfAEC2
ms8kxdT4tR0jIFsM1F1/vkx24xEylXYX0H58gxsdwLJE24q9Q7L4pj9xTVJGz/LAgNvpwXlLK9Li
cxk65l5IZdAe8fgZHIQ7X203Yfjq5o+2qil4r4kVgc+N2v4RVlj25Ehy5U+BPXFSkpZzKPT4zIN/
8GEKu2kleMKGgXMPqPjoNqOPRFo2KTDfqR1VQh2gwx1U0TRLomCsYC1zWnERqC4srtUAMnsyHKDJ
5+Cou1TupydYiq3VRozTZJ6/zwiqolQ39NIEtc1uFoSC1K9nUb72mX+x9/jAn7sAyJdviI3rjMBz
a9yCh4aSH2JYrR8wztcHhCFwZzyrH6CvDAcQqB1Cv6o6xFg1T/tfNYG1qpHsvzTtfy0xJiWp5Mn6
YYDBRRmiOmnolTqn24DBRjpKTEh5aEqCMWMZBnBbffTSm9OUnWRNuorve43ykf6/yT4yzbsQbTHm
P3zBAUzBbweALLMBXAlQiccyGMawZGK0kt5RBAP0q0ZpA7TKtzFwpu+O5E8/PRhT6+G4d6XQngO/
N+/XFKB0gRVuLY62b4Q6wn6LHuafv07+QPyDaY35v3VcnJguhHyItId2U4JV6lx07VcbLpV0ts3P
lmvp+xeVf10yabrm1jP0bB27Fqtjzwe4vQXsePbLpydA52EZszvqDVaYhjcIJVJdAUIU/EO2mqSg
ZgkFwflC7blsMV2YnKubNayCEG06JxkvGn+qbZJ7CPawzIDZa6G8oS+UbgzGx77Pl98GuNeK4+pW
LFuXgcAql2wcFyOfm3C5IKNYATgoQSHpBqLWgbJWRUiZx4p1IuWJ28eYanxkp9t2oULsA7DWtgEl
ai350qZz+BNLFWjB3ZNilGc0OC2lw0YsixUfVJXLN426Hux4tgSam2fmv/09Mrp0TOw6+AO9rOEK
IqOYH3kstwsUtLlXK6Mem2X/pHcVxnOi6420P34ZBnPb4TTW4QnYId8ET1Pte3k2OYd8HKPyrYxO
TQTZsF3W/cq8wW9N0e6AjWpPfljmnzhlmZdlTfJV+kzl9TTVWfO4f0plf+TiZM49uuJaFH+b24tX
BcKEdAwGDyQEoSHPhcwazNy4ktjb09Ncdejp3CDoBxivHrGrXn1gzlazJqYQyzChNf3KJHEPHQ7C
tgUrrZ+PT89dnDjyxZ5zQyIVU6X8bo57d10q18fZh/aveHEvTx4avr+tClCqUjBJ0O5wsXl76SJN
wmLF+W+6oH+5PGP+oUhtw6TSZBIBaK7L+YjzpX61b3sTMFJBp8Q1PlD0XzQmWeoGjaseTSdU+ifd
mb3xKnx6gGAxuB0kY2ao+MLkZmqPjg1c9kbg5Ms/lGo+uGSlbE/ASX2TiubdJE+nw0OyWu2Jl76w
NeYNLfroK6/czHZOCQCWqKww+pX0ap9bVyNaVKxkqAn9P6Luh5OM55uoCc0GgIWC7JLwUEgE+gWF
8Py1d3gzTeISyC9CSb0mOo12yCC1US0sRnlxgl9IgSUi5asd8B8iiuGLUt+05qBWo2nd8z54Kxjl
W80bFtJ1GAvuoc1gSPchQyY4xWB38movCp7nmyFTC8xUsZCFWRYL3DNgvjwVQEp6ECR9dokD72lJ
f8UbRWHC7D7d9yAv/aJ9ncjKr5+Us4R2TYPPA45NciHtcIH5UA8ei+SHJI9VITRmz7Q+6tGvydg5
Mgo8bZoIOWaJRHm/IRM9Z5N5+DbAF5MZc9C+TW9zVz40Z0KoVUWdnoSgAVzi9X5BQqOOpgNXu/l+
KpEJSlu26Przdc/KpM8CbKkvzVq1ZY6aOo3bzsGmm4sjYtOLFjp/Fxb2lcD68wz9CubG9mm8ZsLs
ILzs5u9gj7wEiDZzphCDz552fy9ljRZr6dhjmIZNSYk75uSvrk3ZCh2v7N/zJnb2lC4+WLeJMPGg
e/7OzdIhzgZoou49Rrk0aQAcX/DnbGjgKNe0W0lYlgxkDxNioLM9r7anNgjCJGe1rqUiHTQOyWWZ
SwtaHXRdL2gQCGSz4w62EmiC3akqegq3f9BA7JYmY2UOaIQvlWQwV0uJ7VW4OCCL8TvxicW/zGm3
CIUPtNffoOfBjGSQABH1uEJo67GDxwDM0+RTsKAaF53NY0SCjELbw53I/fdA1Wrp3uK4I6R+gcEM
bBCHWTg4MawhCBNdYXC8Evs7d07fJoXf0UBmQWd+dZBkARze8sf8q3m/i7+scSIhFITj2xh6edXk
FGZdxoyzg8unfw9MkP5BHZe/10Dlky2iNh+iTXK2LVxOzAsV2d+taYfX+PvXSPv6sYccs8qXrdXh
0UJMc+mlHXFfDHo5Z+ujv6XAVj23Os+2h95KNUKOhcB0lLFmYVbv+4ecxD/409TXu65YDLdD+7iv
ZT9QpRvM8NY4O14C+vHOf7+w1I8YiEQBp+UbSusXlmsuyDCJbtEDchZXe1Mhx+zP5W/TzuG4SbC5
hXOUwxGNd7kECFG65jUkToPRf2Qbn59/hceKap5Y9k0hIpNg23wYrLUc2GkDs/Ssmb77J2WIYIeG
5AVchQ+gAevwpVf8Be5wenvyFqcYx9dxMI0eKiq6U6ebKLonM26JoXwdneAUjJme79SAybGAQOWe
/vTwUaiefCrIjlljL0cQoMpbNCDJ23q2DvB9FXInG3QxE4p6/0a8SufNVv/PgyrpXwPv9O2M9QBD
CgHfqVXs/ohosi8s1UKAyG85YB5MIogLLr4Qk2kByqYB2hPEo9KlqwvS7yjErsQK3pFYnxZVyDHe
tEAQD4VZBuc/3vhVXa6Oy96GGBorJ26wrAUhnpCpDC1JxfOYPHiIkfNxwS6lNrm2Z1iiGo7lCbr+
QAjtEyBGQqqhIrzhw2uutDZDnohV0pnjVPudLC//Km83/EQ+S+/4kP17eJjuic052Lz2o2Y64i1l
bFy9iJCKdjOuHYEyHKamMjNoT2AiY2lPA3qIvTMB9106XmZ0qXQ/9cWLh+OVYQIYqb0i53990usE
BgkH2HQDpiwCptAWZ4f+GmE2dgo+5rsX0BMXtmHR1Y+1cbOzyJa89rVvaZVJQiZXMJl2GDz0iP9F
iT1XIluEwU4FBKt/xgO9l62SBjnA8FBg6bycN42fTVQ9WcVkgtpDa2HBkalOLnosGXBHtAUiQG81
pUJnM8vZ/YgTT9b8gTv/43OcMyNzylP7FJ6cDn+/+j3WOL+JGb9m0QcOa87+WSVsSa+GHDD2LTou
g113ojFSvwyS7PazTP0kpg/tPnbiEqKykU5VyVXqxwZU47ccR58SJHmsUi95BHuKQ+S5WL1uc+jO
S/9QdVONTVNT5Chuad++KXAAejyawpzm3C7hlm5Dyhtriw1drkv+EN5aClUyGF3KlCt/tr3WKJXe
JxLTpAy3jBVsnWG7RhkVBhkdApohB75FSbAih6yfCIRlDETBf+iuaqlsvjBV2Em3qGn08Y0jUKi1
lgwWHowUfGLKO6OwYn6/kyRQ7p2NWvToOGeUu7JSVMVBcXurFIck8gTbKNTLzRXmhRN05GKuf5DO
SK3rcaQnI+XiulCxMnlvvZB8q/xmoecskxwYu+kReBOCx9RCjK40cwHJtuSG73izgC9/pAgKSfxX
nzc5AfobhrH0keYekQ8CtNHn6MtzckuciJJz+gTuldwOG4Wkjyjn3QrrwvEf6GJMeWcphdMDQeOc
t3iwLiEOHZ4DbXVSCrNg2ry+B7jbXPhm6nsjfgp2/NIAQvaL0ri/TuLFxRd0zXmqI1b31PIX87vq
rEpmM9H9kgAYiNpDgtqFhGE98KitQpnP7QLCw96pY5rXJqBt+wbIp0qp0L8A6oa4RL9q3U+ptebw
N8hWfsvdexuXGd2vAVfV8qBnP5WbEZSgw8UijpQjvoCaPyzMya+2qGm9J/kiFUsT+T2MV4ve6U2B
vmN6T9Ir+c8cInNylv5lQ2SjtuJ6iR9DKNeCbZv1oSIiBMJ/EKtIR9AVOZpf83CgmdoJx8YpYpMl
RIquBF+YwkrTn/dM3s37MDyK98CxZwxeeGG/SggKcR3toMfQtU+JbJ5vo1aVki+LPZ1TW9NQYZeJ
HnEJ2t3Zv59TMSh+KuuYLffFO5INH8goMIaBGpOhAEKFapjlxV9MOhzHJAyeral2U1lYdL6Dj+F+
xkajFnONJytHPv6sMBrodvepT4L+PLs5echDxoTOlBEJE2QEZokY4WH8strk2r5t8qQxNc+NTp3q
QG9O3FOOg4D3S5beZOFvhRBwUW1f3yp2Yej39VFAeCE3NyB2usQCvKW+0x4TRZBM2bVmj/G0ccop
p3cabFGy1RkzUPeeHDpsF1hSGhdvZ2MFI1gjleGzG3gcgRhI196GcXFbGS5wWhfQskToiN2fFZvs
9++7nBHbETFf9P1IOq8IGC8qSmCPJ0MIlCZsO2Nz6EQvy0ki0Nsi7cx1kTMvr0sQWOof22/3vKTk
5F2U9ed8GZ1ZYmCFx90E1E4ZVZKWDDuxSmCcPZt+7JjpWQ9loSmNfIxXw8M1XXr8umGt+iUBWA/P
9+UHZUAILhncczK1GV322//z+FRtvmiof5r60M6xaeOWnZ8PfYmR2hGzlKjS3uF9SZmjA5q4SZkL
7rY1WHsfW3GmSULRUVbupRjLPGMP0BherHSi/ojGN7IcGpg0o/Jc1DOs4AsC0lAjEnEYaAiB22gL
yY8mCoXlXsO/Tdl3qMsMWIhANHo2PjIk9pE3OvoQByktEEL4+GOXr+pF9Yae08/X92xEFbBwkZYT
eVv2YXnxArdPIuCN8MtBL+ZT6PGnkcCd6a/WdtLftvkthoCSvSmyHoDW991TNjYOPXW3f4M8lemd
78bSeebtdj7c3SrGiCZPsAXb2+XKzZSw4PK/bK7D7s0dzYuMa4f4h5D+7MglP3Ips4ciR1fL+EIm
oEaQThb41i/NVR9j4FmbyV24LJGsWzLA/dZ7ElUj2UWHn3fXUX/omYv99lDhxKxe9AjKCvJtQRpr
Eb82dsKTIqyjQlp0N4PYgyVIrxIToFkYNXT5igGKUSjiRBihyO1q+xsNentKtJhQrwBcZae3EPm9
4aHXchCZvhgHggSOTS1j0bUY4ohNqm+zZyr2TW2dFd14d8f/se3nZzdkqGhFovEnh84OyhCm4Kee
Yl9yAZPO+M6roIB/AXVzBRG5fDqw37heyoEPJwi3auypLZSVHUVRQxPPfpzi9nmxHmspD4YQL9Q3
f5sAiSugouobXKaS6OsB0kFfS5Qc7joEn/M/43Mhx5K7Bkjm+eKyzbEIXrLkldldWbo7uEFhNdE+
RZVgWWxPZku0y6d1U4NVNKzqOHDJTpyRXFZ6k43GyFrjkb8U4hIXLQsHt9AYYu/ZtWAIZw6DtlW1
ExbCz/POGClOl6p8wVjHEsrXDfKdRnmpUtmFK1Fdr0Ez672nfRS2BpXvAatxn9spsu3svGdvIAox
vytJeS0AZde+BkcynOQCBGVTs5u5RiH+D3spSEUvkWlOnXP59YEKKStYDGJsGAMiF9vbVzAh7fUi
fvnhQ1OKXiLYBpX683Y8+iQ4BD01rJlhSyDa45fHihQuucUey1mT5tDvWa5LvHRekikshhM1blQt
5Df8Kq/Vx1KE0Fmnn9HsHH0mFrdhNs/rRcutNws9ApJzftqA6c89N5cBC8OU7JYO+RlWsNvKD5/p
5RQ4p8d4v2BdMe5kHKjCCNaaJOYB3CtL29cwF4/QI/Yf97z99/jzwy3kid/m8VeNgojPfCGW/5+y
2GoARJWAZ3jRhkiAgmpBhNI4n33m6CKcDT8jjNQObgyh578x3VGdWYmS4FTNcJ3UkEVQ+IGj1/YZ
QuC8IW5dZc+zMCneQU97TI9CbEoDiHS+5tMzbosIW1TfXCHvwvdbJeZLAoiKstceEA5G8FEs3TXl
8pwLi77I7bIsFXH21sDATLNnxtPwNs31YkpFNgkfQ1CdpYy+77iWYKuXAGHvBnGYXuA422tqfKse
GlO9nYdxZMaKjo73I3B464TUu5ryNlSPHgqJCchTeCxMIG/BOftL+4ingKBdcuwrLJSp4vRie+tC
WfCGcoyfGLkE9PeAf71ST/Q4fIIo7Ab8yFYDzu5UqO4KCpYfmR+krJd1/pJ3q0iVd8ZU+ENe5iMD
5fkZY6W6dHlm7panWIgrJfEInyDL4rBVrWAmyiICEEDGnPbxbE0xQ9fYBFFJzGjBtjjttqVLTyCf
GXz8tusSKEF20ddC3kiQjku0AjNCyDfd8FkdjX/bkCnYvCFNDg+u4uZKIhBJ8uKycl0q7UivVyil
IHec7szIj4UCtNTztJNyUriyoLJTYAl4FTfegkIiSwob70HLC3lWK9ywAUolUvdzLrBsI8PTD0/S
bUOved2kUZ3CHINwFRXbkRC6Sp03JnmKO3D9hNieWEx82LmvZJ+SkAA4GD4cjA2XpDGA5gxPtL1C
DgE8yHA5LH4Bq3xIiK6n/RLp9cMcFKJaPIEUbyAImyuy+Bap/OBT0We7/6g5ZWSNXhR3ceLAKoWe
1jxBk6RO2m2owBsHEG+ih6mOEDgW8a8ChIZS6Ubj3g3xL+TvpKX9s7XipnV3dBEoVfYi5potYRdk
yst4F8gfV0HEVGb5Qo0jkoezfufseclFiTs4ZA9D5axwGzAdgjO4fwhNHPmUGb0LpXbEiMQzRMYJ
T3bXqfacKiXRrBpRRlGb5WFZcifLxH550IMnzPboRycBfVdIc4yEyMjD3wWJy1qci8IhGB8IWOee
Lluf6jrpf5QsZwWWOzOuEEI0N7RZilulb7INJiK/SyaAzP6xDj9RVD8v+fapuhBL9YJPBYoxodnn
qL5zClmj70bjDoiN+CollprNdioJDxDZkW/4eSES1hT0rAWVSkG12Fap3jNR4z/NXW31qujIz6e2
33TBK6YJkXIl3h44vyidTBX5P1H6ANyVn12+bZqkhACIiIjNFRE/eW1p9VyQ8DxO6zJsfOCzJ2Z0
3NTeaAFdH/YigS+erSFIPbsqzVhJh9/m0yDi20YV2iVPtIszJEKuiAa6e1UISTeQIizw1iR2K7lx
wYCgtTq8AMxQy/nVMK/62ItJyzdnZrQoN449TjXONnXuygy6b8qivL19TQzVqbNAcyXxeW7vdZsA
4GRwy54pxCySUpKxxS1Apf+lQc33b1h4fzxnEVR5AQ/5aIONYGh6HVuDvfJgcjHHLFmUb/NoJ0PB
FmnPrey7j8koj2ZQwaSU3ipo+y9yaeqcl7DiI/1BVxKvFkLE8S0jseccGdIcB1j4TnV7B8F2Z9mB
nxVx6xI4+tsdWhLE7c/yT6Rhb/ND4wMM+LkF9KHtBNe109Libn12uBLltopj0Y2AdfOHFh/oNg1Q
sGEayXFFO8RuEGQ/7YRHFrNSdz2JYwXK9wJf6Q46q+HDxi2k1HV7qjEXPRC7XtJctK2svqCkV+ZJ
IsdcmPgX4JO7ek5f9AmMhSM+sYLd8qrRrJyHFjGwoQPK9O4PYxMxaupVp8msO+6VdSXUgEKLRxjQ
1/2ElghY++SUOuw248ZJUSck/nZycaodPGiNAab6K5644BEocDYy2vgOrMHXan/pSUFLm3ZCUC5R
IIGIfvMKLpXoqhk/E2aKxq0210O/YNUZF1wmTbUyJQY0b066VQt8rAx89B5stUHS12pxMbQCI1kb
Ipn9V9HLN+gpix0h947cqvzyEM3Ijd5Io9Pl9K5qcNMMivHEffcXT/fT70Yr7gdbxr22Ws4DcLzU
ck3VnjZGOP2oUSfEqJ7Y3zQgCukvnqKdDfpMlCBbnQHiN3NUxihO3fXuBKbScNAW6kqObVMFbLy3
+5gQDmwYg+NN/T9ASFQ+a5lso99c0jjEKPdQq3ETidh8MBY2DS0D8eYbMULd91w5PIDJpEdw+PCL
RohT7qhfaDPhLUL6uys6AVni0fAHR/2g+r9ULMSPK0rRip18JiybKsDfvVLHNvrns/Dw5Hweu7U9
jBJCrZHrACOphSNk+Tp6P4h1tMTgJ++XOYou7STQN/9CbwKOfWmgSzvWM7rnStcIQD6yxpdq12nQ
tvnIn+IsU0fTHOVI/b90341HuyMY6MOr2gfq9HBBCdBIwqZ1yWr3VSkenZU4OtuY5nPCXnWz8VZm
304gGJETkh05TME2/3T97cbbkIbXSNeR4i77KV8Peg+9ErFJyU3wQmoC8ip2cJzzstTqBxoZWp7I
laKSXrUfXZQBE9MUSJgG4TqwtZqMCbnoL3GucXnKvclRkxFyIXHXRIzFxhrZbuKLnOpgzb05LP36
nmycTK44VpMrryqeplT1IBlj01m3Ay9EG7/Q64VmCtG8t5mztonZvlWHdJTZ57U84D1KyySYgJf5
+ftv4F6QunMWiL8pXhkjRXOR5Du3KhU59OHdy5VF4i9JHkN9KX5XKiSwfHDZMUGfdRqAiTve1e0D
BDOQ4LcE+vWlIIJTn6V32KgGkjRGUZfmEfSy88Y/vFDpJDtAGCXOWhkEa2C94YSKxLj0K2n9eFcS
7jEZBz3mbXV+I4bhUna+xrqEqy+yxgFsLJZbJiK1sehNVZ7eNX8aVsLCmb78Y5H2JlifDm8vvIKi
d/jNu0YFfK29fPyzqXCV/kKVh/WPUX1MZiQO4OqOLjBv5lKaon6jTtzpJJ3TbnboVmCaLgvKRjah
X/y9KNx5QaEwuNnH2AmrxfjjPY0zgWnZFJ+cJqIMst+GJCXnJtKYPvBU7pjbqDNhswta3jEf6tgb
Wd5ojcO3skR2LrxsLltBQtYO1pTe8dWID/e4Mfq+agqZ97tVmIjdnAQs1xtLcSdOxjdXzc14E7++
v/5BDPgaeAN+lABSwZZs9BlG02LZdbVbQrxy/s0PoKUWz0fuY6B5N3Ua8SS6UmX0aufS62s9wajt
is0tWNyvSHCUJUS2dbZj9BTLkGqwPmK1LiQ7nq6Lbeg7SzPGg5fN0B6TOj94+zdmwbqw2ptiksUZ
EvMKi9S/l0knbQc6wQDdd3hrLOnqIRA8Q4w9QosQ/p58c0PloBU/URdAQWND+uCFCFpuBRUv33DS
Y+v+Fx4lUANSE0G/P4s+V8qtMQm+c8zPSQZbMz9P5cUTaL+H5qTgg+GN57oxguxjUoKKJJGfolON
62bty46LPKZIPdLGjbo/uWXMpTR78tmg1U6dOmF0s0Z0qD4NO26A0xYprL01P7Zjx8M4zNb6My9v
Dfde+uJrlkEsANcRgSyWoE+qMmIEplwZi3GsNoPtt4ZICdATme2KZU94Ki7kqY7QQwyDEB6LGW7f
HtX/f5n/VUrw6eE38fsEUxUfrKS7mvIWbtxIfTOq2jXUxWfwn8zfEOkbiWvJKmPSrQnZQFuo/oFH
IBPzPfD+qfWOP33YK4BUk4TEjHmKBmUo/9nOX4ZjpU3KdG634QCdbuRS7byVrDwTqvlMRRVlndAT
rc4YIMxHmj/u1TrljpZQFuSdnBqW1RwZy6aMW8/4KLB83MKhWvKGtG7kCi5ve42uEBUMzjFfDVX9
9ztLPJY4cfWCod0ZE7zVrTMUtLljvYYNUqGzDcINPj7tTbAglLTtTk2xh5ynEPR+DVZRDluZdfEK
9aB5PIf8STnZoW61FjMtMCxQtX1kDQr/cd/5akJ2oUzGS3P1Bm1LxDQYaGgeEgVaTx08k783ki0C
w02T9SsmGCjnJhvpuiUkYobdG0dcF/Fqw5UdUuFwEhnZvjdOEktWrAA+rJnN4KAaVUwJ0eq6S7am
R3exOJLIRragO1/cIDNOhkQ7VGZ/jv22CC2y4uaDt+Kcdd9+RsUu7N4NyPBai5sr2vzgKXutRv1z
4qJs2jfvhowvK75HasvKHC49mjECPVR/5dYyzRqzvuIlap/bgM2u9Og0jMMrch7MvH83bjQVlPjn
IQ5xiE79AtzZUHs3CUXnHtTLp/BKjw3P70YGdlprKznRRmSD3vxgzHjHDW6vYsnNy5JAbLTq3wyG
nEaGQcD/0O64Fuf/NpgQNaCfnUs5C+G8hURc3QLUhxxlzDgfdV5sRXahkFHuJxWXriD1HRXcb3As
mhfmSiXyuDFHgf4403iJhK7r+2SHttq9XV6xrNe+zJ/1/hbcHzCdBmIZQ4FYhRa9XFvKzdq10sl8
13J6aUf5nmG6cCvigKGIoNegCLQ44SIqfUF/yQFaevAF03beSA11PJaQiILq2LC521RNAJ2hlfOG
E0OXMFPjF6uILIskbwi0kcSam39eUBQ+TWj+dIP8s5q+Rwj0YUENY9Kuco7JeBrvI+NJ6b4OKpca
FawRBEaLmUKFGaYIfK08pKan7fe03b7BzLDi+l9q5B/0GLDBG1LAa8ItdWa2zamXIV7MOChCng7g
tJpUd/mLVrbqBai5vNFwCkiSh6r5Nxa7+8wXeaHVfyr9IoK4tFMnCCxyp2y/Mki8cU85/rpSFPq+
uKotqUjkBy8SQLkkSUt+fZ1Ujoyy+MRInZm8hkpTygOvq/y+cu21/9kFgJm9xf6PaEvYFLeLjs9y
D2xKMd3cZnZpm5oCuHoP6bnob3ExhPYIwNQiJx5g8Ox7FVjzOQIeb1j4rXHrG/nimojBFRUFxFf1
NK4vZDhtzvTPRuhwek4fbcob2gKLYzO4TbxIBW6G7vKiDe+GO0cf+o4aLYWNskZAiLzEZ3zoNqxs
By2u+URI/Bzwvbdb/jlq5WbDq7XRcUJAUsznW6hiOHNFcRCQpDF58BEKRZOSU1wOislVU5sGjqTP
cerx3lJmEcJCaz+jxQlx5J2QGMnKKzGzdqhNxGFBMh/NMx2B45qg7lNOJm7k+IottRZwMYFF9GXI
vuxkQMBpKWylgek8p2ezA4vvgdtXIwe60uYlYXPs7BkBV+Ocs5E8o3yt8gFizaQx4+5tTs5CW6i/
zIxiMqxO6fgLJGlwpsm9FFMYNPdCqRkza9jm5RrXXmCK7GaDo2DtRrHsH5QgP5HOJWGrG232PcpS
z2neoOWectekasJvNplbFZI/7R9XyCbr7M0wRP/XSRfwz41soxTzEHbazILnTjZDs1PoFi+Ym8He
3NBNHq5xmZvQnUSEd0509p01LWw8qvwafJTT2InKsNWApfBkQpErXlX0/R4v1lNQ9vbLg5Z0G8GT
iQ/wfuZfsmS1NufmXiRh4GBZBEHSgP+8a7DPJRYwR18upNh4mcu/Rz1C7OcSDglswG+E2MYnKyxf
pUVvxYyrfTouzmlpRwEqTjB8vOcSrzyshARNrxTZ5kvajsd3Q0L+VgHXdGr5BUyZWpMQtH2yJi0Z
lxaqDQQvd6OI6wO3zQWEjYHihfcNCBy12FHvf4DumvqD5OXAkdqDU6G4Qn6d53Is10VvxVRsEixX
vnvUw1Px2M7U/lYp0tEweNmr3fcq36KxDbVa9coAyaUYrqQlmVGWEd+riZMfwRlEs1Y73UGayP6D
6r/4/NVIPJfQaQeqLfX60nSEU/qjaMcPQKIA/aqh3lfpIclWwtmF11IGYrLKj0Oho1ZfOWZ4gpN0
1wPAmEfsgedc01WkgYmpQEf6+2ItlZRc672/8F4iV3+wArBDPSIEEPgCFrGC8y5fjAV/BW2ICi1B
BHX2b0Bddgr+3vLzSnr2B4U4ikd3SksxS9If/kXyBsVBl4avln2iJQvis1gzPw5BmImQgD4tMpSX
tlB+PvdjTq0cnJthBZam/Ttd3/1xucc3kTqPiKHw41iHtVGxq8y3JkPebQTQuQsZ8ikBzK78HxAN
FaNG0kjERAD0drHoxH2aa/l/KPyRInItE7/q1/SLwqDuzvbwne/g/6RM5EiYdNTtiSsm3FQYqcqr
zE5xM5nfQafuqYweWvjqYSFqqinmwldGle5dejUTsklu88f8VKQrWpFZm4RJ0B4+0WgfvLgrW+w+
mv0P0meQLvpIrA50Y6cdJ3xy+KgHKX+jUSG2ew650lTl4iP0grVFcLM/uKE7soNmulCOETb2VoXR
Qt22xayV0ySWHAtQzZk0RqoxdiYXhpAyjzrPQsYPPISkulwbLPQipa4u3Yx5fIz8UiCLUBg4eqf/
g6EE0ev8orpyL0QhxjBAd6Q0pQYmc5TDvfKgCZYCa+woM6joSrFC8/MrvLVvTxdN2bWBn1e33VZ9
wI/i6mVHtRsuijOFws3Ynk6fW/BvNG68DWoOhy3UskGf7AahneygJNp92Du8p9tNeHNYKEuu0Ubq
XrbiCxTx6w26BW8igKZZHmcAoFXuCYEEy4LSFTD9XsACeDIzuT64+9W2gIincXLBNhVhPRlcq2hM
hYKW1u5LqC18mmUx8FbLEktiudTnHEPE7QvfkrWq8NmRpelG4xiydzaXNBLhPOj0n3jNXvq3UaTz
g2UWcJJGP9+E13OmY9YNl6WXYiuPDj/hBaPYtXG9ePIWlbFyoDGIRbZhQvX59LUaQUkXJUFMWJvo
JjCPgLvgNzm8EkUsMyJ4vYoBSBJHQqqVQW097cj76hu2UP2H4968QNk6ydpoJv8rNgXxLM3to0o9
AfbjoTAhoYpwa7lOx3DQmL1T6wflA6KcTmKaDM2+e3qKxgACFvfdn8mnvEGADP9MS4RL0Dtxj/gj
MurwrsW+3N/gU5qGGfbMmnMkG9OAtjdVbD9FbIqbiWs4TrBskLCL2euzA6IRsEyBqsXRoUbBQjtM
vMzy/+s7PGpWEiqNNzL9DKwR6kfZreMrT4/dcBmNjwkb0HUaz8TwKwL1zfcZ/co+usak5F7+M+cB
yPbwsfLA2FZe822uQEbLet9gHBr33jgHsh/VvTzRYbqdDbFteCTV0F0d15DPB7dNIJrdA7f3Buav
BU8bBG4aHd4YISSmDmFnb2ocP2JmDQudANhpgoU+ol4KX7+fnuZGG6y3oEBNuz49CZiwZovGO3Hw
BnjLJR5KH54ETOon4cYYDeUix2Lusif+OOIQ+UIsoPeOYwZ6uyq0XbVwdonGDKEzlyW07+sBxxX2
ird5gLviOmjSWy76AVIZyoQae42cTo+mU/3R4vPrlnx22DNxafa/PD3pS+jdFDHmxy5lH5CIsOyK
T/lS3ermai0WNbH5uxpyH32cLhy4paXt5yf7HZBK+T7UZG/YKFFSUaB0Wxot427UnMjcWCfGyVc5
ubEWlq43XS60UhuSpZVg5VaLm+yoCXkbmo7YDqDsZEjaQHz3JHsIfTBumuRInLr3dPfvdzzqTVsV
0PV+aAB2F9hiOg3NbviDEZ/e0sI/3JnwRLutV9G07sXqGw6oLvbKtmFekZgtyFsxELofj4BMluyg
EmCEz8GJSBvEORfaiZAJh7Msa+J0trRoVOObpZpQP0PrH+1YGrDep3W7lQQJ5C65zNSsZtv2p+Hh
dTlMQdPXmtkcCA8a+77D56SjEv3pLAd4yhXTiO8Wj1VTRTPGLdvxxJWpQlFN5c74mlFsYuUxvF0F
N9nLEYDk8n+tK8SKTU9lSz4koiSM0HRIVlpVOAWb4XaG7OJYPNRViWiX7+/Mn6cls+pjTUHPZDMp
H3Mk+L2345eF55F1YGoShZ4FaAytPqmXE3mkUWTAMxi1yZGhirne3LTguzXWQz0APslBge0IGfg6
meytlfG2wKIpu+8KVUYHvZxZJdmZ15smaqq0LI9PDinLYbZfSRMpeWIjEeMoQJ5s0OJDndJdiTMt
kK7p3YgZIwz9hxZhNYw3PGWA3dvKHUfmKjwTStWqAA5ADp8GDq/m5OAEnxqqaqcCCBMpU9ZAjr8s
ZjZs8JC61SSZM3l3iALtGILjtVLc8ULyLWht8AH4S2jPIQxPO5PcoDIwbHXSqltZZvMjPe/Qoz+O
SxEnLTDsySkAhN9bf/GbHnO2jhG9IYZXpYoxVwQHcjnhDaoSTUQL5yYKWWfhBGI2Hx4YrkSSanfu
ut7WHdmPC1u5tYSjCiYha+RbZWWaChlc8/dw+Za0DTx4VkUk+WMRovBehvzwa1yOpgIUIGWZPT04
Ssk3sEAB4pderhDSdhj58Rz9XBC3aouD2YOKS98JD/t6xfFbhUy9VanMwa6oaVVzk7up+gc2b4HJ
UNxI56cyZTIusXhZF/z3HbP6Ax90S9/FFtcIbGsdzn35eIyizG+SqENdm6gronA2oWZ3VDAjmmfu
TfaxzNGC9kt20MAlyMn2BJeL7/SFLQf0aSTk4A0fL2knHscuokLFQkX6nCZB9ngte5Dd690dt1de
VAH9l/n9KYZqJMnacKiyUhbH4/Qk9i8F95VBwT2x3hOJz7Tn/jcMgo8306seIU/752xJMFP6oXXn
pcQZqRJFqdr452p5GTNxcD4VzLkWw5MmjhF8WZC+VltporNy9unwNRqJ/35BcOOzeGfUXmJx5/yf
YbJE+fnKExVsr9wdFbgY9y6dsq62+WHxKa/j86wtRlHT5fv/prvmy+gc/xzezf346foDUuhjUNqr
bvPLCNPKiHVaBXIbMD9EhjUmtPCZl1DmUiK1eL+BQU+Nt6u7ScPwZwuG2uiBkurOnL+IPAKi9ADw
8LW9loa5ZHoC6fzsQTaxg+m5u+xfASCk5PUwqBAoCNWyLMEK3E6D2YJEF3x9Xa+ziDr9ia4wUfHe
vXBP/BtfbsQqjEJ3/BXDcB5Xx0RvpQCdAmWOPRUXea/GnwZ4ppRUw48UgYLUwC2HJXD6mLQkK2O9
o8RUFnAJgWoNO0cDs35gS8tYXbFcuVXxX1Trez1yw5NYtVhnm7t0pT+UTH2zyhD2HJoH0XuMa+I6
i/4OEo0wuMIEEX2WjPws7Ui20la5L8CyuO0cOsqK0Wh7tWl6Uc9JFG6SQNdlSK0l8hu3v8TQkenq
urMulYrGnlWEhMxnKHfTJeMVLP26A93Cf7NJ1zuVUhme2jqYYHj00SFFjVprwHULLXTx6hEDpf7B
hznlwits6WASOfoejs2Kmw9O2S2281p2j3bXeHMbDaKX8Q/O54Lzovz+I0y0VIfx2ee8FCtLBm35
ED36rx/iF1ooqM6yoRvxbzx1Z+k7PH/OwMOCp0z02R5C9nPHaDjC4b5ay1OdwdYviaH1BbD5/Fik
UYRgHHQ1yW9HQhsILQkxFClHAB6sikok4LW1mkcwN4v9jGR/KPpabRPR3HCt9z5hDtRnQ+xkZykV
apRq2Xfa5eh6nXOaBlWfj0RteG00aHD9nVpKOlKXasKhO4Z9Is0biPmXi1OSRJOSFDjDa6WUZMs9
jsrvfHwPCKZNCpKglY31/THWDSF/MFxeg032rC8fKJVHLaYPJL/bCLJmixftCzwLb8CMQJ4wDfml
c2yAJUq+Rb1aiTSnzYkJ1F0i+ZnPsCux9OY6EesQvN04+pBXxwn+aQ1Hl/nk1S/JXjgE2axMzWDk
sMLcmw3TfZ68uKs7VQPtMSCuzmrwsPB2kB5J8BWYmwfWFADPLUZB5iLaMUFoc4SzzbDWE06sbAly
4yPmvlsocgyzqYpxQwYY+D64hMWoIdleRwq1dnvQpWmjRHw/vfgNOLuKmmAPJOrMV6WHu3iGnsXe
iYvEIQ18DwgpMX+cWwVraYZPkC+EOxq+7MuCQM9xMFzGqmCQSakPl/xweIKv/qJdaRDABz4W+2YP
DU34rOyIOU2oib6cJjVnfj6dxvrufSQVHPtyLhaMx3jjgYtw6hq4HUMqMf9OzUOkAJHbk9WKa31Y
t9zB0HgXY2V8JJgbafMxge/03dqSIEgmKx/9LohvdYYZpLlnxqUmCpiAKvMIhDq3KwqyA1uMDkqu
UWRnTrxkoLJItJjVB8BvoJwj583MfTl9kfr6nQrr3GOiYReif6pMAMTaWAHqrgJP92UtoTb4FGy5
enZXKgTApoA3HyJfynOsB0yTFyimLPx7b8s5JqMlKV4TBNSX8r3J3yUNPVsrRzKE9/I8EPRJoZ2j
2XMeV6PyFxYKz8xYiewty1XwOeC21oyrqn1oTvd5b2KzGVYyafaVfXy2wP/VtMYwTIaJ7rAGa2Cz
OUwWfBFmBsOYZgjxH2d4kObCae/QjfAYoHUYAIRTfGzjsbR1ftZuG8/zZQgMikHRx7upZtTNVeuR
/BA6AYfpyrvGkMX/iPn5mmi8KxUibtN+Nu+Cwxc9fTMpywmUKnEWvv1cGp6K4r0qowoXFLvGC3Br
Dl5Qho2LZVvRSYO4lY6sFvh8lPqN/OhkkgjhbIW4PjNI53sqPJdD0ulcnTBJEk/uIiTCPoP8H+HC
xQjKoCwTgOKW0A/obcTn12h6XjRCt25mzH05Y9ukRe4BEdZveX/zkYVP8O3WIBMvdE0EPkl49i0L
vPYsms0OwwcBIxRx+r1vaT6bM6Tf29+Cy94IRNimwOu2DjPeKfTyjvzMdJA2xVCtUOPt9Dh+Kqsa
JSz0UMB6iiQmtgYgkEEtoJVgrGPxmvp+9y2lxVcMxZaRxAM9uZ3YPCiwF63LIk2vAA1CsdKaZ7u3
viypBm3GM4rqFlyoTerBAiURt+oMmT6LxzB9WKeoCIuqvBI8jBBQjkCphKbOtcbnuVS6dkotyvi1
yOqGVxZu3+HX0ujQ6b/0E+59hfY+gp/VjlSjWYAWxmE5aEaKX0eXOI9u1yrOdqJC1xI6kbB8pzSw
+OYBzh+rcJDwQHgZeW74k9u4mC7u0lFpdMIj6bFrMpkYhYERipE1sIaOWeALNW03+pVeD5dvGA2f
VTDxZhZ6EMcux7V/hE9rNBvSIrJkq4+GUuu3IVi50u9DrP7l5BQicL+u6N4dTGu97gJXXZVu09t9
X5O3p9DI8JJPXm2lUkjV6e6mAt4Grssgb5Z/Hqg+XMga6QMDk3/jPP+YJkozLJ5ni2T2P+2uidIr
RcviQ7pFyTsoHGddWhJkWjiak8aHpPkNWyOGoxrynIuYC3ln5hMDXHwfzgA+Z14daj1vgYuKKqUZ
JBYl6zY52qfLabFd3NR0rn6izrb4bw1+z+7JqtUTXzMdG+shAfrm9VgI3h1W0wvHVcEOhZldvk8t
BwgLJJMzqG/KJfs+yICyPpzYX/LV8Q69PZlNmcqG4cpZg/uNbG55mcW4bHkJbObzydaLkifnt6wq
MM0ZxMnAFDCrswIlhZc0Rs7stWCn269nXOkZ4y6Lw4SrN67RN6++t367xYE0g1G+aUo56NiwSuFW
Dyu8A3DCzeCc1ZNLKpdquf8A8mGXeaMOm6r1f0A2ky++bbt+c18RcYFOZZWw49seUotg2usoUm4e
y/3IPAIZBjPpPtH07XUqP8NKalhUrxs2OPXeJaHYRoiiBlZT0r+TvPnLVODeVSh4NbNzOFtgrCfd
6NTZVvlNtEPZgqPVZ0LYRqUI64RuthdRrzkzs1up8ho//OLWymv02sU2T6bUYbDnWHCzjS5mLxw3
Mz+eBLxgNI+0kN4T0VHk92x+fBQgUm3hsQ3fseth0Oi7WXs+RrgUhwfJP+b7ujmjJFCjx9oufBNv
IF2BYl3MqWM4+qPbPXv03oMSQoFnoV/Rbvn7vo+N8qlDJZrZA3R9yOR6bU5n+82yyAldM53fE7c7
WPx4iNG6mXSH8+gRC8W5CKfS0ZZ/2sxlh/RIbIgk4halm8z6Z3NrBrPFtBOv0NACZKt6XruAAyE3
Gbqp2/xu9l9N2qL/i5GYG2z6Aj7VLN6h9UZVdQGLCacZMBNy9i1/QCdMtBvJunDblMr6KBxcx0YE
DveG6XdpHJvT0x3m+W/H6BVIQs0h2C5GlkoDfVfsqTriqunGwfhViQnB2AfhwZWA4K+fSkP1z+PB
hvHHU+6x8+pwEZFe93pSv3cnkcDTDpoNmiHOxPZKxJFmPqG7WdpTOGQ9GEsu9Gjj2k5YTrefRfvb
OKaPlxmQOW0REls9pmAzd2HrOE88WCPqCb16hFp2nloKUl0jilUW4gDWBC9TBHd5Sl6DpwBMPKEf
q3GJvWTnPfS9x1iEzwWqlyBiIGJ0i57VNPIRH/iM4Yxyd4OTthE3YA6JRIxhW0IkNB1FI+w1auKV
0Cv/JGwsiDuW9CY+LMRr6F3WrgBfWFULpg3WzsgyPCVlrk10Oo45p5jWzDdXU8zlIdV8DWF/xdHM
q42y6v9/iUfq0LTcbY/h2ESHEw7ek+0WXiaqOcuLfKWcNUdQ/8Kq2W1iwDtF3egQFAib3DH0XfIt
2EuKp1YvtpsZXpW3VPmC+d15deoVoSejvVuI8wiTuoNkrjVsip4EfTIV8a6L2sRz/T5Ekf2hZklB
QRxNyzZ8mZNCRHM783nsXMU987WLtGdyQv5Jrxu9UjdOrfEzPWQL0puhVgH+nH7dE9rGVVqY3Ul9
rKcrcyneIknrlOLDoE5pKX4GHA8WDJLP4eJqq0jcprAbT3ROgbM2GT0g24rwpvLgPTfz0G5RPEFs
HRPvD4cAH7Dmk+UFM8N5T2tEgtn1m+GEEnJ0xFIEhN8/NrBRmI0U6jXF7MDlwMR2sc2UvQIGXqFu
LnneC2yMNwMWK7CyOrbdjPGS4qoAwLd7+Tkjds88E7r7rQH1JEGc9lP5+Tvwl/o5hUiOv26vcZJ5
+bgxRPyrGZtWRsUYDZg1wxAR3zlc1Z7xoKDR5SPDbfVagPM5Kt5VMa7sOf1C4MA6ips1a+8yCMbv
D8B4ZIjYH4FGLfw6miwS3etWDGEPDhyABFY1lGrxtLLa2ZaP8hZ6avs0Eytq/Z3NUXd0Eetef8S8
W3y1vvcPXK6JKfKLG1hmZ6Ptr1YMGV0Jrl+dBrVEddP7bgkV1lY4buuVhYRbmwsDNPWk1AjyeHHx
bazw5b93HT9WkKybSlaK6Pf5cqSxWk4V0DD0MmtFZkuemws8PxVPE6k7W6Cx7HqEMt1TdaJLJlc/
n2nXrsdQ7mBmE1eSMJLX7l1wzYWc0vQavG4ux3yCEfNH3KQLHnwYnRCnvHmAKfhfXnvj5xgl63Xy
0smRIUJgQwioAfHcNu+Ryke2F7BwO4frTKEZXoYEl7Ypjowxmb75+0wdHQoJEx94igPwYGSkbaRM
Kyu2Zc7MC2R6pmQQDrOoqqHo0huDwYblxQkfHbSGcPUXxvWZK7V2P08Bcm/Ug4k5sn5qx1k1GRu5
0iq1RZOGvrQx85uQco3VAbAQrQVg3jePnYsA5Jx+a/RdvkJHvohXCN1I8V3S+mScN7iE9SOMDl57
6m8N7E5KEdvhz8GFLHNbLhtpRxB23Qq9ldwyGQaJ6oUg2vxPMIes0csi8wJCH0S1hdbu9fuAVt6Y
0Z4mhXIFeN6HI5cxPKRXHWel0GRrcAfUDBHzIyKyc/hPj+RdLnTJL61FlVjFVGOTMuouqgsCs537
qDU5DW/o0y18JsOe1fVbxwngaJ+x/xdTphgJ2gjT4RXxXjDxnVCPW7xPPdmRb+KXxabPvTT1dhTI
LwLeCI1XHBllxnO5O+aLdWumnZiPnTKh0J6vRR5UvngLxzm+RaFgIMc7DLUEqeO4VM63S92XIodq
oaSGyjc38xnfboNoPXpnVvnI+i9iCgjaJhLnjskr8wryYBNg6TiR+gnZDNN/YE4FlDuqzutvX+12
DvGe7OFcu/TVaeADeSkjCG8wwvbBs0VU6yer4Zqf+3ZuPlu3A81Mxo9LlgUhpay4312ga+ptCQZl
3qURes2VoZ8eCYEIWrWQUCZ/PsxVRqSn5Ckdz28RNyfSWHP6pstUC1a1Gla/Gf1g0q2j5WOsjFkb
8HsdbXclFD/OPj4ubYx3JyOwxeKddqFTG7IIvkg2/mxGIzaEDZ7PKgDHS4x+68IiW0txip+p8Nyp
nbiNtgHrBNrHrWDGwygxLwBeBEyjeJsYJIHSns/jytAMUmC4OiKo4nXCIf+tmKiC2q7uYaxSr65a
J1AGIe6XVdmsdA11AP0D1J6Lq40z+6Fs5qLJitRhcagvVHuoj3HCmf6T3xZQoe2NSA4hEg2cHFxK
70Tdea/SL/qn25xovC7E4I4D8QoDLbVHusd+fsS6APhObcAUzky1oXTg2BUPPSvd8/CuhIgIEDDp
cf1YjLlHxqWlN8zvOHeBLRXb51REtDT5FTUzIUXEFvKJV9pdWI48DH8IIGmP32mWLlxZGfbxsYHO
hPxRcvOITcI2kVv+rmF/+bXZwPM2cCAvNEDRXfcWOPC83ci28XsDuNfZNh1t+Hb0aLGQC5F0OUDA
X9j51Gv+J1LjzyzarL4aa8U8d1dxZUVnxObkmAzHOt0zb7/hrCu2Ca5YF7kfwZ6Ioc9E8s6z0Dlq
g7/rcAbzIachNWfgTESJtBKRbU7kskRs2FyloB3sxu96PAaCtibHnRlS4+l2rZI4mb+2oA3ot8Uf
zuQXBB0ABq3+TJsWDYIRCYwfRPMCS21tcBJ1T36EHscyVKna0eL/EgmMhyAYOQOqTiz//ih2H+4Z
YSwnW5zrqDKQhmhn9uhw0pH/5o/bIKyhAQ3b2VRGppRNv59sWTo/Pgq2PkHyfzRpu6Eky2ACj8MJ
tCFisUt5rNmoJ7tH55BwAceo+dIsRNhj+5Zz2sEn6e7MbbiQvE0RALrzobyB7O2Dob2oAbTfIIVZ
AgjSWtcYTOdml75P9m5UenuB4m+xnBNqjd3H53nYOzXanDpGEQTE+feodYgR32qiafLDZw6zlMci
+jHx8LlntRur2lyeZ5yP4lyHDQ/Ipz0A7dMCxUhVk6htuCIs4GbXQNSa68QeKpggmoR5ER3w4a/1
+Nea8GfB7UyZlQRCcVk7zeFekqR7nZ7ASQ92RXtAsK5k10PiLfpWzmg4HzUiYMC0VVEaXppjLLXH
aV5kelh8h/5y4tEUAV6IVs6OBv02821WlC2IXU6GuqQcDLYtl+LVgv2D/nt1xWaTimjd+IWcFbRg
YGWT6juPsLDP/lhK7lypvCovnL9P+9L1rjojbKS3ksDrWmK5CS6ukkG/MG+h1ONnAv5OkGBWMvtp
yljKrt+mqtfb93Efk+0tIxq/XD7hn/TduOIf95wqx37xcs8X9HRI6zo5Mnsp+3cY+lLB9Ub0CcxM
xvcZ8jNa1sJR8Psx3Or5SZql/+9+8tQmU28hEPzBh+wggmoDRyVGd0L+TqTlmr2/NBTccrsjmaJq
rfLu+pF+Bh5giyAVfYTCayTKrqIHeblStr8qxuJJId2aDTr6/mlx6j1iX5CtqzdmpQjZO+kXhbJE
2Ec6jUJmLjLxlX8+S8Wrqsf3eUs5jBmS5D3VnVsp3g6bMtA5NR3dYB4RVAu/52aP/UN8CBEkGOD+
xt4TO4dUddYDQXCnHJnggYmPJnMJ9byoUSdcKQwOhnUnHB8oeyWK0SM0OkQQ6WzTZeP/B9lAeOaV
T1vEFlLYHJnOafAvCx8uIltemJ2b6goHd4nKQp7DKmEl8DHp77cP8q4ch/vs9X2yIedigAuYTVjQ
493qpWQASHWvvX4RL3aDIRqq1d2Q+TiMgB7QPyxBWJsn+Tx+/zEZyo+HD+9pFiQEgk8n9dnwngFy
joYekwDE5d0wvqP12gXf5STxMPwc/KY6H0X04n34HFhPtlVvZze6Bp7p5cBGBLqifDkcr82fb6Uk
IZQtH2vaDCY9ht2jIQaRfvkW+MFu9eOEiVAQkNE38LE3wfn/ZoYLBhIGmoFxgij+jdTYLoaDqxjM
+9b7adIyOwM7vFQ/DQwkj7HqHLjisGmvItyFn3McMNc6SKej7IhgEHk4KWK6eD1YEqOjPzny9fDj
VN8J2f6CoVgkAnR5A71k17l1g7Cp0bVxDzjFEqN+H0Z6a/S4vALgFKz5CtitS0VEd6XQUspruDO0
vt1Y5jf3etyvXyCYNDjDimONR6feC0hP3E8+KqvigeGteKqFrc02L/HQRqe2Z7vqcCENUssYBviX
Ptn4g8iscZgo4LRJ5fAYkew/LeKsnwkOycGLuchPvEsrRyBVMMZBHicDi4gqJ6tPtehX6Y/P0HLm
fkbtIGmofZT/iLVpM8EYi7FKRMK+Uh4bQwkD+gAyQo5+yy10ybZ7oOXRqZRRhkCQfBzXTGXPIFZm
W2hGxh86GANob4EGVZmJk6lyPX2a5fwAvyFjcs6n7dizcid9JG1k3a66IyPImO8fZIH+GVzMr2DX
XvntxKBIXZftI/+nSdj68gE4E83Fc/By+2nKcDro8RuhMhzDGzp7Xta8sb+P2NqUVaiqV/ZPanJz
R77LKC4uJEmnnr+oOkILPZ/PvNvCrcaBy3HOeLT239CAIQP/mq4aJzsR2+S6xZ9SHhZyNnrDuiDA
bvBmcgggpcIO0DeBTVkteLZ7OCTlw4QlcD7AJdH7pecncA4KbQ6YPmbQI2QnP8PupbFO56tNoNKu
B6eZylVdfQjH2IHUZS6Tip9hI+/hVGdOG/8EJHsscw5se/oMv0brIhHNlI1Q+CI9JEsRuzenG6iK
hMSH47u5NjcvbcvHSGJ1YG5GksmtILFmKYT29HpubBe3ryWa7jF74zDXJjE6He4UxpmKjyMgFW+8
SXKwlkiKQdWRRk0BIqSwD7Z6iALEKSiI2gvZnZbpM89d67oEkcJ3RTu7CLaoXDybf44RN6sv3hXG
eqM6Ks+8OlrGlca8GQxXsc1gnzCwRoO05EMuqHfpEfkljxtcvndrlw2AqkhifWPfbTYHhRfebPy4
5TNdIOF1XNB8JC4A/LVzCgr1LlRRKrsNPVg78l8XB7/HQgV0i5ZLg5butPjY4kpQJSOpsu/0+BlB
QMSA1OCEgW3SdegjfCr3SYm0pTFz5HQzPLaFTQGo3abc4nPSWCUggfgagumDx6ysfYJsVTD1E9W7
zQsPfLliTMK4wob45RHZTkhHOW1kCoZ/rpOgR2JNhXPdANl2YPrw4tKTJKHdToqyHs+c3OsMV1eE
5sz04Wt4GFQZyUXSQg8WMouVR0CgPCeXNqho2SgFbGLixnDZcarhGWgxoSqwTVHfn3kJ84+X2X0W
pwZe5c0s8d2WgvuZpMDNu2SUKCDJhlyC/g/uE3Tw+YCRDcqzeSWd6rNFkOpQDzN5jsg3g0mK0eaM
CFEEU+KvyZ/es+GSkAoz35aTV4FZ0NHq9hevBdvvpmmiI41cmK3DbHWaN9H+R7J5e8POAYVsrZKp
OfLZAjUIpMXltWb+eF3r1zAiUCSYdv2ufZtUPs7xU+9pbZ36CnsDh8eNDN/twSDKcegd8BPdeIig
jxN93j0vZ05CoYd2/G2o28zSVavzFTB9NLuffRyb/bW4QGh2gIoNNRpHYe5R68dzb7XNGhPzKNL3
06bLppYElSdRwiWWRed2NDMEZCryERXl9TGDK8GeslQIC1loDnGN2RUweXf2VrgEpw3shLMM2RPe
drjxC/jgXwyBI1Q1rLpLtow/ulQPMm+lN5yfQ6fK/RThpcGMzCUqTKBbI4LBOSI8sIuYIqKEQ+An
RNl7gLrC/u0KVv2DNBqbjz6HYjHJPlbxTuuMNH669RjbBJhRegbkzKjBFruJmZI+auOJnUFhYK7S
6ffTg4RQyC3lfp7lTKW1j/kvlKdqNzmfJOt1WWQOBwi7SfJy8GoeAJ3jUqUEJgp7IR5vDPQeWyYi
gPTTnCinJqBQitjvK1bVITo4IyGNIhp8Woiw+5S3rzwKMrtlxd08eiCScnvAU8S8hjB3b/8UGDX0
qIBVW098k/yXdEIErKyTLJmpAdTxfXaspoxGpV42GDFJaVK/CBwB0R3iSurGNwsbAMwT+tlaN9uC
e+zf4SHrJo3x3MMI17ffohlowKaS014L7jkqVPpfXX2xmHqgmZhgT5Bhldlss8Y0+UsyWki/bBwy
vwBdV02n8FsWZcrJWuslW/HBPhTifZy3kzPsQh3rGFjxlUd6wlxX6gmG4g+v6Nyyn5SexkETHHnq
Ye61dUuXD358qzrrYZKqsAIXTmxrteLYGgSDqkaXS5pSnsrsJGVPAV2CCqLgG9hzc/HHpywmiSlq
LnIIaY1vb1VwSOEeIgg9EH2+bVwOYhIJJWuEHjVYKC3EarfhKOJK0OvvEYz9/1D6BQhUVkm9fA7n
pj/sq76ceyR4kXCIPeg1+MEPvXB2NrqDWXL0SfNyuW1UhgE8/SKULdyLRaaYPe57M9zQ//tSv5M5
HjCYn6oNtd4gyB7Tw7VNC1sDPivKp7uY162vdYHlkEyBnjsdjFY3S1djVcm5MJy3wVeOvbr6++Ge
kdsew6q5r/KEMt/vlUrN+XfGG9NJyUJzYSlUTdnb5LkHYC9bGKBjD5k52IB7sOncdgZlRICEMbDh
2mQ+5LcJsdqNDbvXNe8Tprf6t84QgPyMwKxXsLCXXihxWXxllhfVAUcYc1mIo/7bAFLw4o9L3NxC
SjGuNjm7Eok1psJXy9tyL8uif+Ri1TcS14lEfQLD99CZlmHPW3iqcJLCEJ9enffbsqL5GImoSmCt
AduxINsNFqv+qcHAK723aKZb+AZd7vMsKyztmAvqEtkffaE8UXLa8ELm+MWpeErovEiUagwR0sop
NLzqI4QCE8kAj2zbT7pnRFj7kfjyC0qG0mr3CDiW2tkp/FGgKDeRWq4/KwDgfhVJQGpepmsbygux
pvZeR0o1oebnqSybnL9UMDiRLL/lgRl1FewQPfRwA5pzeV38AzPQVh3jFCF2wEDXb948xi2yEJEI
l8Ywylg0Yjmo8bEc+pcXKfXCt4662I8rVX2FD8ZtTA+4qCs4jYd9sUaxOzbo+6+fNrTJATS2bjVc
9bB1iKQA3YYvE8Dx4BdTrT2oEh5XnTEdOmm1SEiZSur2krMACaWZxG/5Z+ixoM+8lvi44Zyc/KND
Y+amqE/pWwGHXn9S7Km5e0QVJ/nkGZH2JZe+ydol86L/ewDHfiIfwDLav3yKCe7/X+g+MDVbmu5d
C99FR0Qu6W3W+d03xcdpKqRZS8rX6PpqMWDyYLa3puDdUSVPfCG0rrNAC/nWUG/JiWZHsYdB2sqt
3GjWGFXXl+9PhEllQRg9OLQgDYrSxmhAkzjgTapQGC/fueU4aPh6+RHsr0H2vpZgsC36wE7D2kT5
wmlOHKsuWI9bcAAkqtp2lxNWWcVpSeKVehevIQqzT/C+/HrsneUh6XS6J+NF7m6eT+oK0ChuQ+BH
Ri08d+kwZ/4bzvPkyUfTu8RoVgtvFhJSETuemhdJMAKWqDPmHsZWxwowQtPWfuGHuGt6anbxHus/
3HFyrZqvnI0Sh1GinuJJY2OzFMgfi9H1/4Q8+X6cU/rwETlWf2+n2piJaPSulvC9XRtB8nmD2Ee/
2aGwhK1TsZRBCxar7G9UEo23QJ1V2u5kast6R0CmJTx1IVw40PzURK1RB2bxdsUAxpHBHYaP6xdY
fTSAXNXvlr1hZ13OQtzwf/zqj+WGoLIRRG7mL0l5HtlYF54e83yB6nYtFc1lTlVAa34MLuzaj73G
TJ3kW6Odv3mGsAPYP8ZoQHJOmkbBH0jMfbFY2G+9PwBVtavA/1wDlnSWOJOFV2SJzCeoVcB0tVHr
aQhcFpgRg3tsL+xc7wZQETZKQC48nMY38Zh7lP5dn8I/n/ZUa9MLbB49i+oTwXtBMW6/WysF5Ope
h+Z+X3pxkV68W0PzwZvn2A+RKNJ5rbImkNQA9NFDfqnxvgC4jSyz77TyZXnwGO/f8BZK8GjWt4cK
1QOJArEDW/h6enbPLiT4WrPvSaMX4qEc9/6Yu+/P9hTeUlVlkGpzndJnLlxPNSHEkWdAy+McInnk
KJhTWnpUH5J+6IsDlJvMu9kEzyW0PhH/2vHM3cIWbBDTrhLhlWEDrrkyOt3ZWm7FNIaLWhgN7k6w
J3tewKjIHpNvgoTyqSS6ZjijHZiMpPxRhm0WgWuxMOrUTxOlnI/Aiw5dCyWA0wH+l0Zi68adoVir
ZQqce2eOEPgm3ibHmU4F/B61F7v+RnMQu5hJ68JGlYgCMtewg4wZQVafOjoYljnFexINnrw+/R0w
W0XqqUiD51qrJnOO+KmEX3nLCVVZ2WQJCzB8ZuDnHxuwIZdujfY8RbuPqHKRzN2N+lDGcVAQDQNh
5HIi9+mQb0jFiiWMl3vogDUkRQ473g10rLnP2BdjteG/jBf47c+YN0N6Am5N3H9wvVuiRBdEhe0e
6CqZwFYqDh1Xx46o+OzRIlpT6kPh0vhO60T7+Nif4OHCleGz1i6mWruvwVkLEBU/r40ovRgp0Spv
zCJnJSE2BLAVMZAwI5fqtL8pwHol4yxIcxfGqj5+2l/TGQj4pXU9GQEMseaTIf/Yw4qH31gpaOEW
/cBC8m/lLVlydrUMTrEYJB7iLhwTmb4OmsKlqxSAuc1uUea30YiMEogCZ+F9BXiP1J1JJVQZ2rij
LpRkBBwCTyVA8EVowEJLKXlKhPQpYJZHAUO+QvaSvU9hUOd24G+Iv0a6Xs439NgeXDLNnqTBipAW
O5hQq3l10GcmiTL9YRGgDEDHfj8x2JCgr04XBXL75u3Wf4cfpvA6TaHCyouF0A0GBN2LuPtQ6GCr
cU6wEeDDLUYvDLsSecWnj9rhusnibBZEtf92kR+RUtqgfxLolYJGrUrEieka+YBUeXQF6qNRrUWI
fxzZ/+hZkc0CdG4I7t9UfWB0ov7B4mSeCbwcP5t4WIlSxdHChdv3ch/LricWSzoR5P4OfezGluLH
r99TzB6BL9ivnTH3VAd1Lh9vok3y/LRoJkHfyPnY9jiKbtKt0Ubn1YXUf6KYtlHUhFH9dIodLH++
EAsvlNcLY/F2uzhwCvK6p/iqZkpzcYkpdXSROvFyH3LKimnPEWM/3CdxArldf5a1t0bj+GHXVAdO
rVTmrT9FWviTxjGwz2PjoxFEXqmy8sbp4hSsO5pQj9NJF82jLRvlB3rB2Sbgpe9vH12RXwJCOg/j
shRa3ihxp/ywn+5jo1pS8GYu0GkaKFPC3XzoxA4qaCYO4goSRsgLU/9LD4KV35M3TcJyS4llPTqw
93J8q0GGovPCv7F3mqAHKVGELota4AO/AcvfAyQPmfUSNkyAYWEFnIrBOkN2XrnQvcwVb5Zs2VsJ
fGNuVJVpwZdcfrwq652LjcS97uftFVxxAVtV3YQb31SFfMhRTHcii0NI0rDDzbUi93NQBz02BHJg
w8zfUlRv76zsP+r0PInrFShk2Z4b1PdAuVVDUkW3TQOieJgGQ5+QBQ2yhHW4+f6KIZ+uTv3maSYq
d1WY9BFs64ZfGtmmAUTrrkIFVTSPfo0FjuPpzT6JhhB3cBfDvUp0UIUW3xFgzwgfERyM0QLrJ7GG
3oP7wi4FENTXqNXgnN3C0cNNCQ+r1XmeoVGodN7TyTshnlSrNuVnpeZQ3qVH0sB/oNAN4X3j+enC
/7GbDVpWKC4/btizMEbAFEwXqLl16ac61yoNYHJEBQROLvPHhmqKHNaD1cQW/IjzPUNiWek/mNBr
gWWbPzmoesDYebIU2NLR4OTSI+xgHrRQUN0UGVpSP26586CpVBua+l26BjZVnFRoLP6YYFqEC55E
gtHE7sDdK6Xve3p9DpkkAiQirUuzib0LtnDRUiTJ0I2qs2jQYKKixgY9W4etbQbi+ee7rwAyDqHD
l61RPKPlOIWHPjxUJJBryJoHhmqqbHJiKb8BCqQk52+dyPdNoLqcJMpqsaEqEWsRUAgNRMw9Go3z
mS7jf8GcPEH09iXFbBrU2uNvXFDVSh5EV7M0/7QHLcXHKopvp68MXcKt7icf0qPjXECfX4m51goN
f2rUNahe976c5UtOaorVffQ/QqHonGBNRLaSXETIHnYh2fe32dktTui1yAj6R2br3g+AGS41FmiK
Vmgc1WafV8sZoSFfnZeCiEZmEDuj5Zd+t00t1KMXGD7IsGkiKRoeJ6xYoAM8gVK1Fz7VPSg3J0W2
Pg5z+RBCVTsnHiEwmOkzPH8118g4WKLpZqpD5qZBL6sj8ouV+ASWGQHDgV9r1WBeYU9zAd8O1ga3
6a70CEtcO0RGiVj4/JTku6Rd6DURrOQkO2yoHmESRecOS/slMwNID7KcSYGYsgMNAWhd1k3UZjlv
a4GHIBeKplK6nO8haV8fX0enzIHParLq+kNXivxUZj5Fdy/qvKvq3BwN4R7G3xZ3f41f41o90OdO
czc1FuioLRREWW1CDRPAbmDSaxR1ivlS5xPSYxlpWJN7l0qzkdPHgk6Mz0FoVni5TU7BrWbnDq6M
neSolYuMULjLQkyqhJvu9iwUzL+e6ZZ9JXpgY5CSIpVvftFv22sbj+Rsdq0QwjTExhrduT2vAL02
BXskvFzpiOUxHEQ2OkUAVMAvEtjWMbUbb/0nmkuqQQyWuh8dzrw2TWr6GArwoqeNqxSrtglbEA6v
2wAQjhta+kBR0fw51Ow6e5DPmeofnGAhCIxXak5k8YE3X7Grw291AuRotcvmd0U5QAz39kr+Iepu
EPCMspJN5rgRmh0jLIizerMXNq7qZl09fD0SUtHnw4GDXcANAK9hs/kRCs+/RcWT3X5q0B7vXn2i
oC9wRpuL497t8WMgfWV3ClESOTBEuYUmlphEGMcQ14mPrUaREezWCYa/CAvoGU6jdFEBVe9XcDi6
VAFSGHx/P13E9mJIcrfTb1/gTnkGt/pDyN2hJbsA3uomXrFNrWTrvEMFsGAlSexxAhUhPaJf98j9
ocCrUwoDVFKiPSyB6i1D36CbMnFsU6EU3EodAhUXRhO1gNcAp7iMl74T3UCienj2jvWb85yzfStx
N5XoQWTQQaGo0E3+iL1pRSi9dKtrwEYJJlx4t4BV0qT9450RQaSgJccn1wwgN1UIA7+pFzG5ruPh
NYZ8hMpKm/qmQoOteoamumnMnAuxEs8tOCAIMxp1WHxmX9L/0KLqId+8X5zQC5tW118GFysahb4B
4JS5oEMsK//U0FQqZlczyszecp7evb0Cotu95J2iwndTe77cK9Dha9yLnOFMdjZsttz4vENjLHUp
BMvazfo8IOcPt40kVvq5KoPjXc8Zg1Y8taCWWLMmvyDPfJECb8z9F7FsHIzimh3k6y5JI+HqytZp
tx1tqwjA7CJl07plAzU6h6WKGFkPdHYkxI9Pmfg8HZqVeimTs1bPlT6YPJijPq+81+SnfurgVTME
Mnve1GUt+uF1KK6FnmeH6NGGGRhFy/raonUJtj6owokBKp/u2wkKtoW/0egeQtQbVkn0SJnDhTkG
r8/1b2MoWFVGPdQatysQ9tU8rbutpaVsuqsufcWuzLf92Eq7hR2WiN6/592OWmvZ7wKDy2h0B35t
8NAg8kGekWAPl8JcCrJJ74W7cugRkrqC0otqKDpV7mrZlVcg+JlJx963niUKx2M2IujGMAv4Yzeu
AsLu1rpwL87wf8N1wKd/Fe569BAK1UzqNU7+4hmUWHXxXpMSZCTXSyfFj/zQjHkdXMUaO3v3xZIA
41gEG2oRFHtBSp3J5Ee4XwcBQ9iqCgTOur9GGZ5+dBY1x24xnZGMi4WvY38P6shxFACUPMEVLMVc
Bk5EgCC3f4oIwUMcbzcsTqNzsI+56BxPc8U7K9kboUBOIMWvRN5/v+BbCIWDwN894I/NlPP6ojSF
KaD7w2dKPogKpqTW0aveU0a6C/3naRcRP1JH6kT5Se7n8RQBLHFhLEFE7ilFntecnmm1Wgv7BHAP
5T1kOtz1b9SH0bWGsivkhjn0q4cgiHDb1yJoLyObka4j463VK0/KTKa4wMogMATm8+gyY6xkHZyh
eW8nL5Zs/5XX7ITsUiuump4d9jdJA4nhCzuo9SAR9ga4MSW7Lj3o/ihH4ecOqEZnlpulV/M/rbTh
JTA2i9MB2C7f5JxqKxvrGcTGPMawC6u35b9jKT3zpDR9AW6e41JMM2xSDh3ucsVYlAbQTXropEcr
EourDVBv6f+5Onb9okT8agzkTEN1A1VlKkCcTgLGOuQphra2rxmA5QlNs86CQ5sjMJJl5pb3horz
LbM8szXaHe+ySroCNdbA0kvylye9YkYnhQdqI11NMGjo1CR71aDK3SOTZm9CzXz+JRZ37x4ONURr
aMhXQ3UdQAq+tnfOrFT1mEkQdocqjxgMDDbjGOGNUacMqLjRzS76Gkf8cohKkwCYk7zz09PECtOM
aQ1dvYPjZWpebgktgRu0CmxfODq/T/efi8L27HmjKt5o0BC76mwNht/ak58z9O5aMgRgjjscStkh
WG5fe7cFaCzh3/+t26ZFRz8JNa8C1HsdqqKQosIWaX8SXWlO8JMp/C+3Tz6c3t39T/zxwU1zH7Mp
I3tTxZlGGPJCvvWY6CxIhkaI/qxG288jNjYiBeK0wZ0a3ij+OebIfjsbJakh70bkDhOczUlVBxOO
EeooxNZDlDqB8mKBhpuuL+3VokaaCnrJnB4Ew3PAgKSd9htv90ISIAHjs05iSRSdsjSK4W2zrX+i
tzxa0Ca1fPSgXFXEXJ1qL5TXsfmaM93Zvds4Rht4dEvNpEHxHwrWJT9HHq/Xphe4WU1oFsg2jTtf
wXMP8DXSHG7OOfQlvKpNvAsu3iKcT33w95iDS8qbta4nYuYp2tBpxfkK05xcuWT/FfHWIbtQHGqQ
rgwQGzVwRybmh8kCscb46Wt6EYcALH2hkvjNwjdkXmH++gzdJRWF2W6dy5/QaUd7AFcAdJQl/GVK
ZdaWCndvkqEkE2qI8sJa2NDNQkAfhMhaLaqi3BrpzI3fE3y6lgpGNHpFP3omENW6yZAcOvOIyOS1
7oYw6tgQ11GHcrktGviD5wDI9EbeaMpfj+cz2OzVyVjX0z/kRTudH7LgYH8WvkQHPUTYuhpGRNWz
+g9vPjMDJy9YjWVa/0Yu2BzqE4Bv0Hn3i8g/JvwKtvD8MnRt+RQT59j/Px8quA2wCP8u5icGzoPh
aHr9rSsoSoCAdWWGFUIbYbknsMUbRZi9SdjgfwNDWawIh93tLJpDftXOBA72bn3LXTpnoLsoU3t1
zFjGEbbFILDzNe6CmmVqMuOXr76lD34xiP5lDzfjoIiSxnh44Yf8GpIpSbpbhz12boiM+b3Qy+1I
hAqwSDRc0PFk93lk3F2FwzDB7Qw/Q56TkQZgGcnobWi1WfoG5RmyKGZDNgB6SzrUvGdxgtp32DqO
U+ev4JAeHlDLLrtAD1Pp1lrXDxlKwdCT2gqztOfNWR8mFmbv4HQjoV0Vl6PNTdQ5gZ8Rsl6ghA8l
yfiVvCmlXyFFEQlYcv9fs0V/qrwU8iF+WbuXJcK3DWbq8zCFV21VzDpJ8ZH9j1xQxxmGmNYOMkul
5Jk3Nw4UaAJxO4zmiGpozcWXL7vpAPyPznuBND7zuw0fnu0A1WcE1Cfpv5VqGoXMfIdCMjT3mcvk
MwJ44YKFJk8y1MFiUBz/5cHfclj8FCLksO8v633Z4e8r/0kKy7OUQHf4FGJMjIAEpx+ia0F0srDS
3jYILY87rLBsEFgjKEKYcBUtONqAJa5QJ81eNUCiIrbzZCze1Xd5IvyKqrvdKlWMRJRtIfHhJfEC
AqS5qZO38SfnNckUwozEckcSt7HEsQkdPnSpjHqUQsta6iywrZTj1DcreNa6+uouZlUMfsWTXq6Y
UB77UJ+3pAJpSWXWYOG2QK0jZF1Lw0Hdo5so3UvafgK4csybLRNq9ft3wwPLZdzBqFWtZoeBRPom
Nw6pXSEqXJX3/ibZ9Pu6owVDc0hBiGmuOq1DkkXmUI+ktU2KZferaT0ywVPTms657YFe+fdrU41g
TTmNhhuYFFIK9EYGuZDefJBGFqkXQcd710LWdhYhwVU4cMHJe99EVzjv56VaWvISZ/UuK+sKvgZa
VhcS7grhFJ92MPbmNG5jIufSOKb23uZtPBpmSBl7MhozIGmG63fZT4S+m07ZVx57fXSTb56fDvRh
rj+8qfZgiRa0XV9Xeo74I2qaJQS7sNnRHKGtwDPiumrbqUloT3PxAgxh83Ig2H0PieEo1te/V3JP
G5C3B31kgWVHNeDLsjCzr4OY9gRPZ18yd/i/2AXUY0L3hM0ZSjrAT3tkMN9/94yLRsdXCXYK53BD
f/It6JbIoUN/0GR3c84a6FkEX5sEPxYGXs8AIvOHONDJm5XYyjlozQVpJi1oNktmWiQcuFulUp81
qg3PjBBUG6PHG2F2Zz0yAVe0L4UtxFliefVKe8mGRmzxQbmXtMCx8wgwblM1GSsQ1RpnvxmHOw+r
wao2ivDmoXcBxVvho8Z3i1LWEiNFBxL14Y0QnievMpTxrZCJdBsw10sK64edlNIDwwtCHJidcjUh
zuTXNVs7/jzOK2ZuyNaxaVKeumnKkAqhPs0CHVRUdzN4FqkVtVVoT5sR56MhAIXd3bM2PdKtOJoz
cjvSjbgQhhNrFfhCOrBCKAaEs5VkR/FqvfZvL9Y2ZYoRUpwZ+WY2FPZ41qO2gM1HiAsDrby0rK55
l57xcLXLPwFHCd2IpJfM6JNknMxJ0vUJTAwFSDCIipookFdVGXHXOr7HPzkmnlz7fBsZnove5dWj
FtGN2++m34JNRwpBWSWR2FloMkuOCbCyvfPVFFk8yHQd4o2Ox7U1z2VAOCX5O2Ij7Veh1OF0vcY7
o9IsVHmIfXSIzNDYtJWtA4AlZ3wIRusGLz6beSQjfj4Qf4w44TKZD+EtyZSwsypdfJyiQW7Z5Q7w
4/svO067xwQHAuKe1hG5x9QTrR6elE7YZ0P8oNak2N9mD3sL4crIJakQ636x0A/73Nayhxnm7fZ/
QElsceynyAf9iCu50zuVCxWyhIK/bOJbasE0HlopbLxQckbm3l5YXty8p83xC/cQc3zJXBfUVpub
HoZcOhlP5W4JcWaaW8Ot5tpiS2Jk6gp3B+njQzRwD1akzFrvf408LcCKP3Ozie293aJSaM1T+she
zzkQulAnFF396iIOSdXHF1ZKI0yThs0dM89sXDfJXiAIj++/sFgcx1WNl1v+BllrWHH8g6EiAwir
pIwRJPor5gJgsGhc33HbBGcgRpMM73Inkfs3YpfE1hVUD4KSIiqrfZ4HhSgWYXLWYAGP3yf3FLnU
oY2esY6hrpHoyY9IaMGYjzuhnUIF90qKGeLqDVJYpAa/+oSSknitB2Fdx5j35qrLMbaaHW4E2cji
X4iPkPceqB0YE98RhGAk84nSajgyMO0n879Ly3ORrBauENmDDdZsITdvW9ukzFfdqs+f9XZyI5IG
vkgGixWeLQMPbWw5Lr5cclHl3cZzYCskbJkl3oUShTa7jWzuw8NYmZCxyn7LQIVNO9C5LRIeBerW
k4ftZnOu7XoSPkpFuC0q1nX5wFChGExFY6XFy74Jb/wvq5GC/OENPZeqoBjWhku2mdTaM9DhPr/q
Q2Q1X8CWgudcMQ6qdt+rvHJ2ezMl2NPXph6MIRV9pdrlBSAU0F2qAQb1A633kOZNgyK4rXYvMec0
TWlNMb8b9/gEOL0/i1MV8zxi7aMsclQCccCHwae5Mbc9Q1pgYyWCbVDmfU4rL88DH4pi8sypnexx
uPunz7J4D3ARMgsbOsxLjMPkygfkb5oGUqBjBTjdBDmXvqu/pGmzkLR19buWcUIH5DsVePngPIDZ
PzS1lMLguZdz8ww6w3XCtFKl8OCjaSMSpezluL3Dd8F64RLUtp3ZbToZLPP71NKOb2UD9c3sscLq
SgY7TPhkgzFX4beN6HVhnqAymIsunaiq6uII8t3aBzXv6TKpZovFEQQDhJq7ERdutSBoAwQXbq+C
t3v5tqsARLwOfX5Q8EQG2r/qZkTH4CjzhJaz+t6YSC5hKBmQXpDl/em3d4E5oU2EqhWnRD2t3bLs
X8oNqU7cDlEYtkBJ21aa97CwQjnHd3k/StnLbQLkPtpIkbSnzBk1bZFqB6MWeHmbyg8dCPjNqmxc
0YJedAIV4NzAMwt5npZDRcmed9cDjpiigvkjzeOmK0Jtui/3u/z00ZbB3a16CJ1oQXGOqxrHsVIz
exMOZX+M6alus7IHFM98niEWRmtIm0yHU6+Ye6YHjBdcCCaWYaiHg9MwptF1/4FwRf9+Yn4RXcMT
x2mCWveFhwMwkb6zH6DKWB4FurIJlRWqMa6YwCIeds+u4StZGTrlyzmzE1mU0qHtxvwxKePHjx8C
Pfm9hqlDuY411p+DmDWNqKoVCeM+HKwM0DVZ0XsSKcofQKWJVcg+9l7zbaHBJYWadtWsArv4TRMr
u7zOyAthxdQ4i1V+pDOyqGFQsXitqao6ZmM829dHVF2M8Av5flP25VBqPEId3OoEy+TO8+bbMgOn
sDbeQI67r5W6fBH2t7V1q2qBGlmcNZ6OIYmJucW5xtV5U3udzgECPuqTcymbX1y12SSDGP1gKs3z
Y8gtFu1AibYdGdLjaNnG6ghCecB7zNT5laN5seKzCP1uxbqPnAiCbbUUvLTCvAg7L1crqIBjd3jB
oj6lM6es2LFRNwu42fQZAGKp1XaK4Yh/U+RnKXZgId45doD/mxXeNfS0/2twV3TEMPfkmsfCnek3
snF1FxxnTeh7tViMfvVYlKM7ZdHEZWsdwvP2chLxPc5i6tyMjYUFyT/IBcs+jmBqK8KxSiLnnIg4
xxI1RHQ3pQWCSEQHi9ssEDNk1gSHl5UHHsvwHW0dbSaZQ5S0UotBk+ggJg2RXiaY8tKJJOa5lbHV
oMlMbrpLqxNmhM5E9yYQvb9DHDr2mKai2s2GnuJPRNpzQh7/E2TAZkdK85NZqb4uW8lFCpZwAbRG
j+WV7p6AGQpMBp4r7SzGJOdzxCxZG13Vrr9TwdfwAoSHWFFugPbjYvtoEyFkdNfBj+XNRhGtuzx8
cDiODwbDzvKdAPil62j68A3/lBC7DIWjXhqtquoA5Rb4LU/+7Cs37yN4iLalTg871MAaVNvxty/w
3U5ERNeneYwsPZcTuoKXNh9LZGzhl2E5qy4bHTfTjfrH99Y932VPyHwS6CAFp/ATNvUksqyHS+Ea
6FLbWl34RWXFNxAxylp2Ls2UkiivyrOI+DQ6409OuI+AhdkpEoHGIvhLnkxlIrcR0m7czAPa1Maj
KpBYnRRUMM7eKjr+twEpFLr3UplAkLOzumQojWjQdRArIj0OUiwMTvCus3Ucsj8lmWifgHlOTzZF
ZrCkzJXyyIIRCVKdlAiBEG+vwBmsrlHhqbMGMrVR7cm+44E0N9sDAMHwVp/KJMJ+SclPqBGbH4Jb
rdG0EzwWQ4ps6XZ8dT7TcLPBMjcI8pB9ZPUIlLZWx2BAyvWiNaidfSjh/ufKLqsFlm85SrkOvCGW
8Yz8GsvfI7bzW+Pgh21R6RVp08Hs0d0J1TVgynUsyQlyfdt9uYIqlCN3x1Cv+PNEvxD5+LlLHKC9
7UGgs7xV5KLZlI5t7R6nZkiQQ5BDOM3S9PlDJNzJMauEYxZAa/fErnkmRQf3KQLxZrIVn0fwnlCq
Mpc2FSchX/7C6tTMAsm6uAfbstodXT7iiknBUH65p5d8NB6/lWpYOOT28o3aA+Y6GlnV+jegEcL6
A1pdHYEwc9ULHq8e/S7vvjjJoS2mb4ZvpJRziIfoppQkoMsPiqBbdmq8dAIqE+kHXkpl9QjtGgzC
LeJimMvXId5OlaJtv8tnZ8mSxJcbvZVvBjCaLU706qiHxDS8hi6JSqWbVrTM8Nl4AFDmhiWaRuUt
zErjUTQP1V7+hOH6ZMML6fTT7tenShJM3mw34u2eGzTTJtEZqVBq/Ra73014Lp5ihdDUrRTXC8+t
xm2EW1M6gFuhLhHha7wtT1MP0KD6g5nyiX6dMVK8hq06zPwkFl2+Sq/2ZGraU1pdNpquX0CeD//i
XrzxlG9mNUgELBskbMGEF2f8qyZp2U01kXy3xsQ51u41B45cQjy+kkKFkPjj/cAAWvu5xuAfi+pH
GfOivSaM81jZEz+rgvumUFe+ijRXttptzM0ehuQ9eljP/ZboyzyllQOWREx/YUiZhquFFGdAQbsl
uTZLbc8A9xZ3MDmGo+nGbn16j8F5PTbl8um/PisLx2I86C5N4u1JuzDGD6bsRuqc1tBCi9+vAUWF
fCPaVQfGfGpG8nowNvv26aYfYcPX93bMBp1umZ5oZjlp4ZOxzrIu0W6ObXftHA1ytvfANvVPRAyj
K2uEyI1R7gT3FXI+1BRGx8t5w1T6GERGmtQxd7gNcvvtasA0Ny/xgsDKqV180Wvd0RMcnilfQ//P
tIek/qTgseoJ8TobiIs8q+OAIvCPhXAq2AGWCubCVfStByLB7jznAlNGLlPMIl/FcncS+eN6xqAu
qMoYxRAzIO2pOQrbcXWx2YcPYXLKXwj9Ndip3kvtCF/3NcY3dsxTzSlVIGWByCWlNblUuNH/nBIt
egYOQbOHQrsvyaKuf+6HsGk4puyzBGYK7utBkNhcLp38yOFi+tGwYuMTcSEs9QURPdg48oi0ArJr
nCQO1ktqFqyd6iWKENG5LAAZ4sY95k/Uiak4YpEiXzMFk1hyKwJ2HJoOHiALVOTWi6D+11XKeOpm
8mVXGw5YT9LxMA+ZEdzL1j3DbmDHfIEyabExIuJONnjQaWuxOjAuak3byHQslkeF/KPlFc79MfbJ
YIpVB4pmsJWZVrF7yDNbr60JfsL+VwtBBvooEUBU+NpS5IF8fIWz69QT80EL9GfLsjXpBUs48YIT
2r3iOadL3nTHPKRHWM4gBvjJatglDfJ5GXWyQQEztlKeQVJFfGiHTEaYwhVu6rXKxlLMdGsc+/Hd
Wne0bfhwvXrei2/SMYxobns7E50DcnWucTgDjxEusO5Ak8fBhAY5UcIuKZ1CtiUBtcI04YTXhvuG
pkKv/12R8UnBEzpiA44NZm6GasufQv1ql8Aecqh/UdvcNrB9Tjx+OhfR/E3ni6D4NQ/UJz3npKfe
xws7Pp6BkbTKYuBt6EjRIgga4OiB2kdXiJJadJLQDcqY8PIFvJ4CRXsKKCy3W1a6WexjQgGvNaxG
FKn8BT+/kUDRre01bDjAxJb/BODJvfkfzAC+n5QET2Qew89h3zbUHUkOBqzbYUhJAVGwrzgwxCyV
04W167JgKaqX/26B2atFUClKSYAK+E7VtBBeskNqb2DrxZyTX8xfWMUZC+Zs5YWtEdnaQCSJkGZp
FwWi5boh4n0mkM/8OSVGNgj8X81kzrW8LaSAdgJW8uvE6wRkYejw/7bYO1xd3pv7/bqDkeDsHgGb
cei1DUK7ZV5in8VyVej4PAsph+kf2QmzhhePACRBAZ1kyWVZ9UIkAFfy2Ni1DRbr61+qTCLg59RD
gFPOszezZ7e94/U1KuKxvh4bdtvhuZbqOHvVywqxD0+SQeE6dZW/11z6YkgPJ8xTX7hGTnKNtiNu
E2LEOeG+mw+9mu3enjSLCVqhQm3JdsQtwJ0YK9MvaAyklD5LbXbLZx/mGV1/LEncDpFbsRNhJJe1
ik6lxTjvekas6HtCKXa/ob+Wun5LpiHwaPwgB+bJvhpF83B5Lo3xa4GGFcMaSpl8q2wSYWdaRxRo
Qjp1xnKyijjBBH6/K6Re8xgzOfFYQ8TOGKKdD4z3UtGF+dwF6n7IVJgTjRfrGXkn5CvSiMr8NaYM
vAQq2MBF3/QgR6DJdbDJeMx4xtWuUAhfogMvIl5SXdPCiWWzHt9aeOpi3m2bzxxPRg448aVY1fjn
ubwlKB+ngkF18OPjZ/UhOcijq5yzoOhlwm4GDneOh3oSQLyiesGly+LvgMCN49giZmA0m/8CaPPJ
a/v1UUEnNppbY5BMIf4Wjwi5M2gHGrgtHoeO569pXAG6hX28sKihIMZn6Jzu5h+LVUqy3qThJc5U
Nj8WBuogmkm2aAS2F9wvV/+abKduDvO0+rXTsfhZEhujRkmhhjQIGapoFwFNcxttgGtqQNltsvJ8
kPHsFbedTrAnMrOG9z8zM72mNqkzFK3iuiuHeKLH6kKtljd97onyyyDNletqqInZ3FMppxU6t2Ha
jt8r15xZwj2egtKvrI5P71mDga8n17/DcEIwvuoLGLPHigK7PyJsu+VThtNwJjx/A5wrj/aPRGYY
AiYwhLGadv7gHNJaSgUTZLhJBglHIfLgCgwgDoVifpt7YbRvHUNIQgg94zJzeA02wUkOoXRXCs0T
nn39ZQYMZ/nhdX6qbwylTAG8wfMrdkz5buzSYRjouNFXPLnX9LfAMXM6y99vTMjRN3aimpCkNQ/J
NeK7LIpmZToIQVJCa4O6r/QrVT1mnj7cJw0nvpB7/WX9dQMmsjcwhHr24PPqhnE7WPM9EwghBrzt
3ga8phw3vdqGk9PXqxzCc53zJVgC8dkPXJmhKlOPINaYuo75Iofku086827yr0BTGpBTK6X24tmp
LuSW9BYjBTMNv0n8laBO8HumDjFZ8lG//yrd3aA23CPWKao6ycPSxDKiPOfXonH6bO7cvF3DDvUj
KNvnfsdJ8ovdwzUIbplxvmF+g79cC0i+/0ksFI8IbPC2tnfJkJUKQMptg9eRexv2UstDf1KOQJq3
t6+BY6fTXSKC5AUlEuXLYjZgdDeLjNQfFLRpt1YpAZNfld/duz0meP9XyG18pM62Ia5qUkobPdX4
3gvDwvGdSXWk+qvk+pfTPBi795YuwEtMDc+/k7S9Wu2pGaVRiEPYh5szqDSlJNmCu5EZQYXz4h8b
bZTPRfPs7zwtHC7XZ0kIwjVCu0m+v2569ciSnp93TGCUjT5frKEVLmlJQuCc1lh0CAV/9wgswV8v
wVBlg5Gn/I7MuEI86wtbt9k6Bi3fxo9kDWF7Ev2pTDbfg0ykIJgsCkjSJgO+3vpcHTdcI/MpfHfA
mwgHpztve9v0cIxep1iGZhqtaXGd80edRYosFDWAyduG1VEIZ7rlx4wPCKhPLHAj0FQTXce4mtoN
hu9kzntBT065yTliGY4VB9J92ZBkBDrdKgRjMp7Vz0f9xGsiLmBjPryNh0T/fF5bbq695Hsdm59e
+Y0pMlK9Ngfdvi60cig2Yb/JmeFwl+pMaLC2/zOlbsp1ZnhGt+tg+P1aT9edzhpGkp35UcILqUDE
yG5X0Nfbim0mAKt+WNVnbWHGsNzioaVor/VrMW5JS0YVvJH2iarncua1uJIOQCb9XJK5NT7FwicX
GRMGGzv2FiJVRAO1fcmbetlqWgRlu3tDy0Kx8QSrelEBjrff8esMde542T/NZlc7oY/X/DGOwLFh
cDnAfCwj3MGdLuUxddkI/eLzm7Xa5nJUzXZN5dj70G4vlWGIvtqnjE+t5G1P4AF9d2HcDohBbyHu
209V7MirvcB18+U5BXGtFrL5BJUHWHStJpzQgsvIizewc+EpwJ4CyYeKnHZGZ4d5w7HJjoQ65V4B
15JFma1gbV/vG3PKuBleQY6Hy0fLrPn+N7DOUrj2y685WX5Cbqy+UWIK1YpkxyzmS2O0my4TqPT3
5gqbyHACy9jsXYt2O/6qKftt+WL83vpL+t5eStn0IIcGca8VuDH5W2yqBqhATGIoh6tA7to8yMB5
jlXm8juvcr4Ypd6LT6YZqy5Jf2BEGwIxbbLsvWDi3H9ZhwF+IT/xOrN4O2nV5BM8xVUC0IYYuGeB
xAuIgqxqv/2+VY3fn3gWOMv+dgGr7Ag8r23RIPYDZL26TfFkcvds4vJvzYFFbkC+w1NvaYd6XWH0
HbE2IcRlt4FzwUgdgpddJ/KGdPJWAjYzCfBMq2qvo8ZoPdRjkUGicLV1irdtBlJLHQ2qxFBweCsF
1Dw2Xk9s80w7i5x5uRyTwzlq9wM4cws34IX4pR8rK8+53mjMlPRzdl0cOyLWRH6H9tR3VE+Ptf24
wQX/AlFsWs1cXBwXRDgM3GQQPmrhjSD9gUt0HvIVr+Csb3SQ0Q1HuvPhHFBQcySozFmydIi2x7B6
pOH6JHue9br3GROxcf51ZabJfd/cUoqtqSSPV7WDUPnMwxZ+cP3NNtUSWxNgShuT/qXj5HC+6DbE
nkTrQC3NTg2l3WXFo0G8cZmT4d/esxLC83CTzIlyqyekN5siuZUZWeihHPFclM50WLH0fJ/cUVIh
eBKgRM1AKHKRyknebtoNLGkkjEF0coiRJE+TRHU1Nqod/ZxXvdnB9MuPW/FXMj1NML+m6Rx6xf9k
c8giHfgw9ptWeCoFEGMToHi/4eFkkkVfPrJhpVCTMfrmmDm51RuT2freIl/QlU5DuPA7M9A5UaSG
IVKsTDxEt0NpC7/npR2ome8XgBeTLIcfqZ/mGlneFx0euxhNQ7txEGPIfHPrJX9r/mgw9hPTUMkt
Zmbd099I5kAbvHE2/mUkoRx2OBy2/Tj4ycC4HZ6yc0IOrT5LQhWL1CSxZfP5TFe4btzHf8w5iQMQ
3eNeweLklOWRodTsh92X+NjLVOix8q+EAK8S4dPdDpl7DUcC7s9DEhbmFLR/HHuSAJvutq9EMIO7
01Ff3rnzsNOK1c6FoMTDjEQUWhswqJM+iX5vzyTXs+I7PotmT2fCSl8eJ1nf8w0IuUqFO5rqi8Z1
qFnrOA5knDJ7wFpsyv2YjN7jIuaIBwmsOrIZLAQ2t1mX4ix8DimvghHmSfwQNy0fjn+uhNI6ascE
6OEEcrQJMlZUi9kIGD7YLlEnIh+FfVVcouFTgAbzq6J65zPU8f9MxtoJZo7J3ZoMta+RE6omQQJm
TbEct0oGemdwkalKyj2CQVWP5iCVJQRuSyYtORzIopq8EtW2DY9wF69DHeOG1XkRY/IRf676CVIa
EMf6P1x5bgoMye+eOPh/ISaOoCXwLrkR2yaK/PNts8XGpOwKJUzURpzhwnfTL4i+VDiaDUWo3oRW
o/g1i7y7vA+qWdtfKlNP53GeEw8wcn+pv/lX7XAI5gTe42re4uHV9rLmI/OseFjiy8D6yrzFE1QA
IZPgNUet9drSxAhARbEBtTIgRgEtiqdeAC6bjzDyB5wd/cj2Owi4q8BO0++WyxzK+7B89ACeDKpA
HbG7ZMwAavqVZt2Yap1oAaK+IuZlPBjCvpJnW/k6LFwCII+iNynJ8y2Jhb3zXHpfXIQOC27nxlH8
2A/L9H2xAUdjBimMI0bGVvviScFb5lhG7JcY+3/FS5dUAhW/gq6CehRz/2B2ESRv0GyNkkfXDLO8
LXJyTdGQU3Gddz0pIl2295DRLrwnWVYacGcNRYe+0N4KXQ+JTFc4m0UFcg2QXEFJTK4yoXBmTDX8
aQaAzIA+4GgzOiSyoTeS8kbFzD3mDJtNB/jkcX7dM6GEbo7ESTgHanW2JvvfN2Av6w5dIRW5qvdM
J3eJ69KaWF/rN6p/ygHajXXLFh+ndjnjuTBkW74e1tHcI87VN2tZJY4hQIBtwb8fhz0MSXjF1QKj
TIsKTtNFNRS3TQR3Zw0wcnZ9W/YqE8tAHwha/4ahS5TCHJUjUj2Fnt72ERtO2arK856g4lkfpTWC
3CS+5tuB6g7wnhHTlb+nQeTx7VQK4kvW30NJvY2AXJAbfOWgvZMdeGhDGXVYgSI1lwxdPN/Qe3Jy
WwWVlU7+Wd9dnDZ2l+seACe97AdqCXNDrlIF7xp0BaRm3JuIu7GFvRiduFn6s5Hl3uxYiA4rM5nj
pyqpleSc6xuanjZqdSfkynAVqlLW7rGuMHj4DevOoJ3WZ8ojZHUDez3pbhQYt5gK1vy6hBYAi8oG
LaGNEANZ+j4/xTcu0sfx249Z+Pz0m695nQjEVLa1h+WyfHP2eWBj0WVuXg3jnbMviAUOSwwY0Ppq
JytXh8pBdW6q5LM04JnpvQ8nYa0CIiRB4WJ+5zxMY1NBkPU2XzLELh9c9QFKg0oHtZcFtrDka23z
PgUv53mT/VVHSOPZPYCoT5ycUZipxbAf4u+G7HfiLLr1FHt0hjDfAd+9UFmLElHGIRejEmxaDXec
lpP1dFDAA0O5eGt9Bzlg6fIpkAzACneGWoOBTM6ot/hoAAr6U6hzJ63Xat7Jn5HQoSRBVdbOn1Id
tFozjMl/9pczutmq8Ro/irhmQf/AFB/YlqlQCLAr8QaX97/krZGqM9FHfJacRUhEIE4K7eXx8LA1
PHCLpLNdT2+hqZrTN8/bOL2kSzKKxloGAvAfuGo06+NGQ4vxYZL3UvRpwA3AVDI/MelpU9ylIsus
+qQwDxbBvlljuPTfVaKKovLmtGMihCwsfm2PdAvpJ+qtfAdTUuSS0LIpIZ183AmIAtyh1PDQII9Y
REx0V6x4PrvkBHdtmYFI5jQK4Sk/cFAbGsBpZ3HrX3AGWMrLm9F5lHQUW7JnFIkeXk6CG7MMzKXl
5mudQU4qewUZj4Yhe6JEPAPoWaTND0ET7ZNA6eISJIiS5lQEsDXkflHiOCeiA18eER2hZrCZBDOW
h+Ky9RHLpW6L848cQHE+ql1M59Z+1io2jK8ehi4vqoq7VqUN0EHuFzglo9tGcRhXaW3uQJTip8E6
vLpnjjabkuHJfj8DLHzzfCkdXOqR1Oy+z7+rhquNNQdtu1m7lKVZ9RKlKWkWPXo1lXrWobaZfRis
TnZRzBelzIT/BXYcZcuQmE4+4pZBufUJtrjBZLZelFBAa+HGLXe8NhdeNQxhqPNfVZr1Qn4vwOho
STP8vzyiFr9cHotKegrpQ1uCHMF1LVKXLPwg18+cppmooCt0dki1aVBPQULT/ss1z5dUnWGop9kR
+Ke0khDCNBG1e5XcB04zy+NjWKT7myzP641yzwaAb1Nq2u4ADi1WsXJYeUlGtsaEd/cPsKuSb59l
pHE/jok2PEG42tM10LFYx1WC9F5xZEFTG5VBoIYLidcIZLgKWmqL7Rwya2P+siMtDgWNHD/IONNY
7D6wn5BMHqy3BFFW4TD9EI1DvsaEqHjtKroU+Qnbl9O3BZVpFAtqNWNKOyvd7ymODSBNiN3Y+Md3
ZNDlopZbxFuDWOQZ+7IcrPVL1uxyoNugw3c9YCZd2tYylqMMw717Rccz+TGFrF7S1VL2MFPnDRmh
xZtksLbp6HalScRpzvFkz0JQo1VGXTTKYX+KD03yyQfPTi2Dj4klla3hfxOTswIqlJJIHksfQJ5D
PlSzaeVL5OB33p/dYasYao9Na/WgFZHMOVpiVggteKJYX7fioKCZjFvx9HNagd6A0ejh54DkVfQ9
Mnp3IfgTsDfj1Fsq6p6wqZSmFaIyCoqGHh+/p5CDGQMPpSg3WyuqG+C3TY+bKICRObjzYykeeBuh
xX/dGve1NJqTN9g+ezYndKcZke++unMcJtErUNIxuoaRmBsKXCZn7xyNjvYz76YpgfBVLRabXKLf
dl2auyqy1MWkwrcjvK3wvvgAb62hGpJVjEgWPK4RQsUkXdoi0m1jCqBvs6ujZVZjSnp0xsY9gvgf
QTf01Nje4GQB127UVdwy+JpKtJwRkJS0M6cTAQ7L5otXuY/bhn5VeXgWvP75S++w0e2P4Gt0S/TF
bvuQvFs7v1ZrDDLVD5ZvP5QZyEW7zEWFB3hYd4TxQtRJ1gkFdCvfpeTT8Up+pRLHnuL7j9rmtuI6
leXNKMhFiW/q5nkTguk93IQAmEG8qMaJK3TT9x0rr4lY/p5S7BrOFFLFuP9zx1oTPBRfU5wjMLZt
XWz5HoJqXQiC6HW3mvVuS3CVzf0pww8cGWwc9G/KnaF7ShTY+7Uxj6iDRbTah5zkhCRCDecEwpTD
tVgGAH6hKtSvatCGxG6Y7jeeHRQvp3gtnXnacurjm636VjdY5CuqACdV3pBpiDsH7DgOZ9j+G33Q
1DlfF2PKLdaW96Cwuf0y5VBpzuBNpEkmVbkll/48yK1ydJyT7WkobDEiunELOJLuoGdBKhEwaJ3J
7B1XlpmxQSX9Sje7QJ4OVQZIVONK1V1g85BMORLFsOcZ3n4i95f8ChzJBqDSG0WYiuoTpg0PyHdw
Ii5U5qdK4CNVNHfAQh2P0Yr0AC6//PcutEHb+d0WKeM1nAGmbdSQ20Xdg1Eb1fbKWjjilBEl3OWz
1bHf1hAlmWnf4X33org4l6b0GK/G/GqztI+ma/fNfCXnlnCjwtP0qWVDFTafsm9QIEbquZi9begT
2/ZL5ydAFc4vLpDMWejErJn90/qgGf8YlR9a+/W0FuAmzDzHv3yo14//BmKdkAU7eP1ZuAYFVqh5
sjwMeT+Po5U27Eouh07ZA8dD4KTfst3mvtGAzC2sETfcQPH7H3jz4O/oCwvtbSFIUt1M70fYiChv
08wuprLRHyJ3hpWqFw5dE4USXGrtF58cuRtGrNhmamtbOFTmVqIqIqirYuJXf+mMQ2j0XNdqWTuW
jZueqQJbrDmRhRQT4pP/kA01PGMzrj7ny04uXeSK0avXIA31pNkiNICvTZLviuLrRlxt1CDGqrF3
PrzQDVZrYqZgWjrl4wpGmzZmnjDoxXlwSkD5rCoJBzTRr3QCW/Q5sa/DAwpAonfV0ei8UBjWNyRL
XhTRonUjXEjgiwxaJzk5LBF/kIenSBH673kBI90cDfoiOYwYduRqPpIymMUr2Q7gfbeRtXZWI7hH
ITPcX6BWYPEprZc1u/5MFfTSYQ8Z8dVaIHxsBRIkcnjy4JgHT1I5VgqpapPj9HUioq6oHpgZrMdl
SRtRBK6y+D+7vlZNXkbYKHoDCPi1LuO9PWzFCBArenVLTil+GyV4oZANlNsRYgg1wJ/smEuk7lId
kd+1kH3+BZJU8zxJuFAHzzHEYKh3W4pCi2NzOTByrBUeunlIY/OP8tJYOrFrOX3B8wvOka564N0c
6e/Tf+12Mlb1yeqg1t10I6JxDUurbyEaNJq24tFlLe8CVkBA8aueMSl8soVyXf+5KL+PYbffuBXw
cAOflY3ZNfGyd2/3SbWfkvzTy81vJj73iaEVsAJtbUdSApOLYhTHK3qD3QldNC1KLiudZNEGxVmv
3ZD6bZhNor0r/MdTz3Azk/mcyD/bylcqvDR5+xjeUhNmcQd1dwuscr9pKwfjwvyDQ5O/PZS/L+pX
LCbhudqrqBliQ1YGYW8z9oVCUsRFqXgKOwdsO+CezceT7zcnyjD84+nSdaGmiozwOqgvmtXPoo/M
nak8n51PLxmka0ViXl8qaZNk87QGJIDCoosmb8g/7RZk54CWT91Za1L15t8qnBW5sx2aLRilwzBK
N4gmKpNJ2LgMov1yui9mY8bIkp2cLJd4cjTfL3B6JoBWNv83S0futHxR7t/s1Ok/VrG1P/ofb3jD
RqulbKt9/b3gymvgBNhWB8DUq+4SnyXhcF3tGvzoAQGtKXiiAR11iekrzG3BqK6Y6kPvt8ad8Fyb
npMd9LcvPGo1aP5HH0sAvxjJMpoKt0yDrsBygpYQuyDQJ3/S+K/kWw8zlyaJramFV9kDjHyoy4bo
7bELW6VHJw/yx+x/QHCmXq79CbbnW+/gA3rjqXinhKPrZts+uwIuUjKtm5Nkl3GwcneG1ixvuO4w
XcOl7tAs63/cqnT5rVMxDoe75b954CGOD850QdWNbnLSnTwN2TSWy7x/HakA/1FVkcaGEAFIvl5S
PP264afCt4lve/0U9FB6r2VH+tZi8cW8qwR08P08h6cCGqGGQoulChTKqn97+GO5vTgUB9EMHSCW
EIiY5Ytpmcm3xYOqaJFa0ScSQIjGNFC6sV64qXJk2vbmZCGkzq2F4x6/m9ILhn7L67JUQCy7Yw8t
z9uSuLKGpbIa6G5u80vlZxdClwHQ7b3Bial0WuyVrXoW6V7AjIuw7zDSvcGU+tI2GMk6iPWUTAr1
ItRGjFnD47s8AzzBa4orSydtjNjHUkd9KFgV2000M6ptfH8TUeaegyZv3KeDy2IaCQ4RYff1q9qK
s7u0aNzbnPJr7zPOFEIjTXoyJUE1O6l/SlwxmLVP6aJdJ8E9mKZbtq0glsZuWfJKOsLTeUQIfH2N
ftn0wn15TK9uF1oFj4PfVEkxemre+fUdqfNSjKcZKi+XHo1/USI34yGiRuXZ4Zs22MngXYqjUrJ7
dSGiwk0A0K/IYUyFAmeE7LfqoGD0k/ki0jHN0doq86MUusMQYNiPnhwubjrpQrPoeFHkBunYxq4q
5dG1bOUaGSAixP2rY5hjRIYEGio4vTnxQkp6pSKNlmuSbP1YucKN7XA8DWiiBhEbybPgefvouu20
JG/T3YrigINiW0zJTh6XKVFTTnGf0rDgIQEVSdBEhGjFMlewQjeqVYOTaWwjLVHmhUeZi+rJdEiC
4ZfCvzERD3q9MPM0CRqNwDVydKFBwaJ70ACHP4IhbK0Y2u9jF5Nqd/ygi40DWVYbknldsegd/gZh
+Hr1F1esSL46YOZTSBT5UDX63CUO379z8vNqQcbERivexeedKsKE0AMOVDhWO8f/Uqchq48YJQEh
vkT+X0i/o2dKBGfwN9IX8xLVc7SbDk+VxMCV1hcjg+dgfjvbqBhGUr8JRi4hhGQjwgVpNwFA0bsc
4hi3K+FMTxzdYEFa6fUKYPhYerLnKusQRg4d8B2Adb4b0l4bnvv3sTKKCVIf8sgWtUiez/KFHHaR
dPVX/u6J87vwSBOk3Zwr3NbhMEXegSQI/ci7KwvEY5HzGyeM/UJVzU4Jq6DvwYtIrY3kai64T4E8
+0/lJWketjItBgKZiTNMaIvulY5rL55cM7ajW3qpvHKyNa3B5rmHK94L9pF1vQqdIspDuOio5NRC
bDKXHACuSlyphdeIch166JxaYh/z8z29k8AP9p7UL16jTbXaPhPMcEouZBtyRR+ySNXyIUrnYOVa
Q7P97xdwo3PGJ1MqvDOYu6YHPnfJdBml2Ce2LWx7U03uZdpj/Yi4d4VO2QI8aR73zWmRicvyZTGe
mcYMHJDQjPOq74IQealE8FOT3ymFRvcWc+5hBR4E3zaQ9FPB8SIAzNg+UxskhrN6/nIfD0Lfraas
rLly5J9yT7Bhhidk0hLwQLp1TKcj9Ao5zWygKEOwYmneYZDB3khe5pa9p3hSuRRNZtQTw2iZVCDT
A3ng3fEIVxaewHk5majJkj0yUcaS2c5yYls5gzjO1rXJ1900O4sUsciMGkmZv3QEQumHYF0B057y
7TqMRKNHxf9owC7XThCsgzAbvn9U368uGPjoLhIeIQgSAQlZ2bR1CaRfbRnLdsXqdKSjigARqQFt
rI2eQWIRgeAVFkkh8UzAwB2Cr9f7RrAU6ShgvR2RYoOebjdy2i3wIbDhYLK5/WqbWeqlBrvPyBJ+
pqk5OFUCaOOp9Lchw+x8NuuN56+uxOZ58JrSLRrV3gexWB7NVVUOPlsR3p5ZgrJqZ8BZIDEeu4+4
rxfNOGbzEb+7daQwQ6vxNRXsJ9TxLU9wkq1tbJw+//gFErOtJZu15xIF7KoWQ69idsr5Xe4gZ1H+
iQOOzyyzggcQliHsSnl9UIF2f7sVqS5HZZ71c7KL9rs6G7cJ/Gqnokis641uzGJQsfLonNtSJwx2
kwzori6nt/QzfVvKBtrFOIuenP4iVaLf1PJmfzObXx9NH0bOm/fVZiwYZwrfk3WYjnfZ4x949vZw
hBztsMK5uuBpQrit4hHC5/TN1qrLY8+kURwk0Q7OtAO+qxWJegZdeGwipl92W+yzhv0rr1SOaaqt
ZhAlI/7S4VV76LzmD9AgCSGTwcTDtgyOvZwAtvjtVxUFox5Jmhn4cm4lgoH14alcOJBQ8Lh3ypJy
IVBroUJOHW87vdfUlN1AX1DVcoc9sotDu8Wul/yppY4dAEEd8u2JMtnTW6BdnCwFSM8PNNiJ2MUH
kcfK7jejXPGSgZL5YVOj2LwC6Ng1TqESNH6xsdEi5omVUMlEUTxZixJHJEBYsnvgtdhBUC8+nSVH
o7CImg8XhWSo8Gp9NRPBQWuhfhyI/tcm6vaJIslYQuxsIGHscyCQx+xlc49HRy8eG8A4Q9cF2uUo
uvGYXxiYiC7AR0/CPEEiVAT+hRSGkmoMC1Y9HJ08oLQ+Cq5WJp9pW7Ae+LrFunYfX/h08G49Qm9U
VdJN0jnIi4b8qPt3WAnRIZRMivQx8dfMNtMDRX4q5Oa6JekjYgiixwRdHQDSFtfwS5cW+HOPnxdr
AWKGxI2BCXCBAYvZL9OndPmpGQuvJ84SDyxU1gZKygdX2oJ5L+B1DQ9AQ+aDxHsgxsEosA3z80c1
8xMcmtaMTRBxt9vlzYZZkTW3CgZ4t6a0ac8GZDtyATHSOlHfraMPFndtsKVINIvwMb/kjlPMFiM4
uG2kO2uRpHDZZp1j1F1rDcyOgmOZf6x8ElhcAsTJKOE5JvizacHTABJCnRY0TNWDQuvCiLvjqROg
oUQe/6WrrVoRTz30GI/qN3uKOw06VZQTvwSU5HUyNVCGr/Lz6uwyKHqo9hFdtIZJSBfK1cjxUZdP
wNexhFh2mCoLXbKuAzM1pvrInpHu0OD6VwFnevTW6KzO8l5Ekb2cPB9lMhBTRWZ5XC2AMGYwRP/Q
qCv7UeZ9JNxddu5J4YkSmZjOYz8S5COzUae+GjJaAWs1oVltskv3AHanBfswNuwFhAgrSYd5lIYO
XXN2YszXpEkje9f67ZBILV/jNBgCrS5SYjBLGRwE4fqs/Q3Zy7WYTvmeuI6f3shOsiF6giqj/Qvd
OxxzBKXCH0+hISXaS9HsB31/yoxmpNGgfVwhtzVIvs/vq0gpd5d+ZywFOtlotaQddMXOn1ORtQ+W
3rWmvcA8qDvffi8+ZsIjQRouSmucZSog0v2oECWBNOpJYxuKzjE5YIFvlpZMsAL3KPbJik/0DsIO
fe4D+QUu6zF2Dlo5dg4mRusIbnyGVliQYDmbhAunRa8n1iFTaVzDK+PTDybFFYv4BlX1L6rsHq0x
3ANIkcyopGvD56c7iWh8FlHE1+hCMoew5A24EiYMNn3W0nDCoBs6a9gaMkUcRl9JVsooP2HdtRi1
Rmy1fgozOs23MXsS0AIIKKMt0mEkfDjZfS3AA0JXJ4pcTKUphVrtS9XgGYbV9HxKHCtiv3+x1WIT
Itw6S1UsOK2SSHsBNhwNTMOWmCWPXu+Hm7k8iWrK/ej+RKZdNHWQUD/bnCJUvWQwS9ciHT21jv7P
y2lZ76+SOEFZHx/NRFPyL96qgul2t3QUkb+5Z8sfITGQyx4a1lJ/TUFtnrst2Gj4PY9+fRt3j+8U
k97HMLizOQ+IIJm5QCi+L98iWXyD4Ol88yLGCaATowWqvjzvBbWxHd5t2JSFg2OEz1efe8T7j3VG
MVXdEu3jdcRp09Zi2QmXUiOiNdNFld/n/GqkgQV27TbGBffA/beAjHhkwc6nZBAjGNWzzWcq6jb+
sdbpvivFbhJcm8RqRE0teLlDEoSW847l5RMQQYrZYqiooXrZt/YEppOJ0qHIrG8ugMXo3fN/lKl2
yxiGDLoY9/kSxptr71SVJtYfOmPlCotMKZ6kyKQLLpxg3jeDvSFjMUrFdrf8P1vAlbdlNxJ+wnaa
vPCqbGaeAdV93tfPgVEZCH/1CduSvAYhWR+/N1MX6UgTxP77omC2JgDyry3xqhZxGCZfzzNRn4sC
/d2HW4Iyqp3LynBt4H2uzdXGPRPLGuO9yKTeDI0InjSnxb2LTh6ZutobBwoy+lvDUeQXSk1VzFiv
IjmBDU8tOHU7tD/zQcpgaQ9ZxEV77ilzGMb+ZFvEJuvlbkojuGutkzuUuPTJH+D8W2+/eYbNSRax
xlmzo6SiupMFrWIq7ra3kQAPeheuNTRAkIusiHzVeEKFjYfP/KgN2qgDcGdvnVaS+9ZpooznTWoe
wvT5y92y8LB2AsVJWveYR08CC6AfKuli7eX154EjIlki74uV63HET8TsaH8OG/ZvpXl7pXloJqEH
8iZIZTp0WZEVhd41bmuCYSOvozxqV/zKs6DnTWYuK/WPwWZHJhNkbiodpLCw7hOX8zHciQFrJxnd
qgFqXhPbbuCgqNg4TyDylgXLBQt0OCEE3h/6r6KF4N7OxsR8ceZQFmT/IguTrGnCAuK2okNROlwn
qK8b7N0OMdF1Eqqrt8wj9bAk+6ZPsYsdGpc7Ypu0uGAnrtLDzFDUPVCJEtFxwiNY66v2pyhsehU8
1NRTArjyVgNI6Wl55SEhZiGFKiTcfkGOyQSjJcDSVBOhzd0r1ULWYDPB5ZgPsI8JcYtAtkIZHAVp
97R5wJbCXr0IUsa+pFBIiC0M0C+Osf5jGgVh8V2f0GmZZPU3bDe0CVRE/2FISDXScynDnyY1tuZj
jFYNVFl+RbnuzZFQrW8PpHk4u7zRJRc+SJzNIxFkX0K9zdJRV4k08oipQgA0rq5leAylAUXPUqs9
Ah0ELZ0V1jrBBHbPnFjkeUKCPVQpqn7pVF++12mPm/IxoileJLB/5H2HXMLceNGvHP57xZNwvRXk
ZqUIMlF/edaiwrc3icGFsqza6dTuuFuAMSTVm1yioHSw4wBkBCb5qySxB8QBijbbwRMTi82DP8GX
CayW+75jOqmwUr90FyfDjNtpAr3TFR9RtPtSLxJC6R7uQLUgWcTWp/SAkLn1In1decHy27Pq0sAM
rlO8H/XpTC49sHdOtE+tjDjHZNpeu9f0VltDsfMV9PxC+uA5E/X31ulLfl7kpdUCOWjlc+gDOo/N
pFDlkHf/Ziw5N2InUzC+YwYo2SVCHhEUg7xAk92cDCKMb9voIFPM/V6wQWAo+19kM80hX8DTlLhI
MWJoZBiYJBkDrc9cN/wGVafZf8Fnv1so1fLZm3lGbQ1FO4bp94YmEUuV/2EdohF42Ft0GIv9dExC
fdcNIVQVwFGRdqoaYtOybj6pd4DgaOwrbPJ3lMAYZn0xvmTqG79vzaH1wClaJVLOR/fwT7875+Ip
oLJ+YNHG6Gn7UHDe/9t4yW/WVj9u+5BhgZFsijA17/i1SY1bMvxViBLju09By2c/Q60qvwTTnMVv
KqVExFU14Ecb+Ybj72pgaNNkDIpl7w8MNSPdLcSuTL6XF69nft9tqA9MqDCicBWviuzHRa78hRwI
wpP0JbEbEjZrAzTns+HOejAtuSQ0XST5aeQUv8zsZQGUtv4b37dO0fabptssqoaJvhqzZTj2mHBV
zuvHyJrrkXgny0XWh09yZUg2XRer5uCzNUl/xZI6iKDeag2XwrQmIe9dP1cqGymUrpmgBov2dusv
Dmmo3Y6DIC/mzAf7MmWgwXgYv+D4UTnr7gBGYcQdifXmhLtsdrDFQl0xQ+1AQ/1DZXDu4ZQIVvX5
txQKfX+3veceuuleDhYY4D2Hp0Rknna3g5DxCxlRtIAXUMMedpR9czlntHpL1IOrIvvt850PHkP2
CkVc1TB9S+HZWxBSFH/utCfkPON3XzIGENcirLVAFRUHZzfSUnhax0r52tLjkwPYqGCsecC4UQ5Q
AaEc3cle12YfXy1+RhgoO9FlMsFCuu6etCJqKsaaj751flbc16easZbKFNsYU57TpUf33206j2GE
hitQrv6kUrchpntJJ7jHlLe7Txsj5MOIv14A2/u7iCr6R+0TQY5pMCIfGuAXt8Dfww+CFsJtM1FC
tM1LpaxXs+k+7etEEypCq+wPbtNto1o+2xw3ynS0cWs9mSmbEuIh8gHedmavDEG11Dk+l5P3WP5D
Am8RXDTXJk5IFDJq04JZEcESpBbKScF+HaCqfLK4fAhygi5wSCzfd1bl4ZBSDeRAwk/XRrNze0Jw
253v8kjIaURZS2g9uXVgMHiMUi2Wpth0iUPjbZE25ltXjblBIoBxwYkODjbgje9WUWaiHlyrDDY1
COv6y7+5oXHF3dIW4s5MBoLB5Os25nc227qMqteYSQKGhutsOWdGDKGxrPufJIiw2hpGFc7IOmwN
gLsZgmUJH4Fzj8lIDGg7aN4slz3kM1vTIUp6Iz+bDAcxdUbFdynjA2Q23/waALDUisdB+ioj2w28
rlz6AOu8FG+I4xwHcRc3Uavv59DNXXUOJg2ounmbs3H3pjgIa1m0IXI+uYvk+anO8lID48/GQnf4
E5mBwAldkFhjvv2q/Ruv0BhggnekezrtUNA07mZoE3Hed4Kw9srHpiTezK8LKov9NUYq59+kffNt
WwY5b4yuEd/opyDKI6tMSW4fU7XDfaVgOxWAfYhZlQU3jJgQvEsmULJvuuZQuEyrwxsQzzXJdWde
79wTMDhiygpCrptswh6wBH3n9OTTksvdt8Ttba47XBCnkhRt3nAoO46x+R+L1tXkXUv+r0eJeJnE
SNKcbEUnSGFc+BrhRQ/N1CEQuaPNyUhqOgmJEmrQUHWqMaRlHy0UIPhVR3VmEiC9RAOM7x7QelVJ
0v2MbnbH/9bVPCXCHx7OShEGHNHYOsBtTwG/fdq9X1O2eWUKEET13Z2Pl4FpkeYJZ01bfNa4Yirw
P3EYirR4G9Gx3aIru0ETjxaKZz1TavtiQ76+tC4m1Gbjrn04rbdUM0v98bJWoEq1tLbVgSrSxswS
x0wqgVbE0FmzyhsZODi263wQm0TT1E2yjsSpw//+PKblQcXDy/+YUspcVRV0t7nL41ocFSIdhXrK
3fPHE1pnTtts64V7Lj49RWcheLRX1gfOet/wWROL0V7RgBWbncZrI+xVoVogkdGb+4F0VIT/RG3W
YcfMcqpBZQnrOG5Re109DYxKs/QjGjAZt15ZE79uyP+1moODGLFx84OrHuidqf8uh8C6t94OZj89
hlYuxqUxcEc6ulb21RLYgQjIdr/90ipm2qrk0SjmiE3fHJqpmOk79CSBQVyMdJvCBMQYBMhGOOVI
en6pJlpyWx5Jak5OLeWpYjATsanDKj1QGbOYlhg54OapAfxbRd+trw0pfsckeXL/TYdcfmTJ7jj/
CBH3GXOfIFAbBGEulNR4kSBQfD+OnEE8yxl9+ZjwCtPdNjPDc6Kszl/G4ALLhoeVGTR8egmeOLF2
SnE/ZA4JFf2c2NfqewiFI44kUcefLp5SrROcUye+kjY0bdKBpcwXytjxbFPbKdxfq0tvbn/+WuR7
lppjDzHOjnjz0/g4j9eVWtB1SJ6+2JQO6AN8jhpeDluaMkLuWWl8HYYYHDBoPK66IdWS0LRx76N+
OFGK4yNt2iI/ClILYM0dMg85n933oO5r/59RMGTJBcpVSxLl7uMzPdtHgWG6PCriz8DQOWUGi4/z
cQ5aG1gPIP8yVC+Sgar0Huqmi9Z1CFWLwHMDEc4fDG7J6EjUoPgSXruSkN/RJ70EBlnlnkfVF5Lt
X+GtBEASpePrBuz9ZwhzfszqoPOZYI2bLcXPqt8gleyApn8fyXq11McE7RIfR7RN5lvzU53be0R8
7tkqIcz8AT1COykQEKCrjeoC8nsT9WSN+OaEw60AfEFry15dHbPyljopoq5K33XPNPXhSkwXMIH8
24neS3a3HxOUS2574N3uyW7IzRU9Yho1paOyZfRmYazPvMQFHqityJmUrjyA+BwdYPMgCZ9py/Aa
SFfeSPibmeq149WS365JjOXMWiOhm4gekcEdlKYS4cAoVVg8VdwG11ffYOzZuil9Dg+thmbvfVTr
adKEg3uJjYBC81k3yk4CZ9E/miOkorZnpiM1IFNmKXrgi9HX5mhSr8VgbseyQnBz0sirITP6Vv7E
eeas9tONChEQZBkHZtHoa7KzqgDECTos+5QrxP4aYh4FeJLrxqQhobSK3edq348B9mnYCsGlKUlP
euJGdqn9I2HoNOqHF0bcHirVTdYjHcQtvsQvo4F1t0er6M/3HFvvzAPtKiPUUzej4dJfuyzWQgQO
5knZ7x3IGwcAlYreg4Fkq2ev6fgkL+/aXWbEREjUSaddXvmQ8pK1X+kvHKBaURWbbY9hg9wPvLGD
/jq7mL4J1daU+3yffpyV9DG8yNyp+vzppMx33kZYvCoKn9xmUsu7Y6ckzRQbbhxrkpPKuyHFWNoU
W2fJX22YejTIwYAR77hvteLEWogsPYzRXE+Zzc09UWsTskb8jUBKMV615qlheNHHL5QLuXsq7KaW
pv2Q8ASWkFmJsRqZrAg5J0mcwqMONBHDJBooxY5ZvJcSZsq28QQJqrPGVUqTXg8VaTJAgqeMwreR
wayw4lIV3IGnfhXSMHyFy/bIwZXU6dofVhNX6asiGZ52NhmwyOQPIn3SQKaoZ8XlRyXTVE5fzJiK
/eSwPT6WwgICbQSFS1ZpWaIq6pOLcDCxhrOTQiM153LY3TksYmCmVMFae5PaM2BulEaqLxLOZWIM
sWGkQyxpZHR09SrgQ2yrnZ0ArBZZ52MSubF3EOlpzJOOEX3QJc/7xgr+nRTOjlBt6S7muXU6gjdt
IfvlwYrV2VxQGexaIU3fp+GRQ/RMjz/Y+vBfdadfkli7mGZ7QLkHMzkhZuS70BcE4ds16MzYz3kL
bMsb6qKMHb8ygKResW7JuabNKV+dChZ7QJHLA7yFsCseh0MNEN/o3kKBkWdYvkh1JerFmfRFrN+E
/jJ6g2U3uzmoFXLNB1f6t39RJ7slTM8hQmzjpvxP/yxD04bCq+twzVedeWc1Uu5l5mQ3wkd15xRw
aSPUnZoc2Vj+8dICmEr/jRTf0O9hSKUc2fUyNaP44BEPAh3Ydh93ZZl7p1m4eMsRZ6pZ91wvsDI3
pzlG2UaEjluVN9lw2S6rKScSoZjsXh5pXRso5Qy7FvUeq7dQqr47caFzUX8X5T/ao2iJZfPBGQvW
2Pc5s719PClAnYWJtLZGGlHQGYcaAiP3xwSOUkfK0HdSQfIHliZztWxR4IFZvORfA0DHoYvQocSU
VlY+i2YvP8a9szZWTjSZcJS13QBCNNSAy38YRYgLYAe4mt9pezKfQGEaLtUl35VhXgVAAet9WqhB
iNFBLsv597JkumLiQFF7PBtiWK0wkhfrFszAad7BJIIsiCIbX0zEkhIjTwhL0MfGJJiMMJNT3xCb
6TQsy7DrZh9BIUmIIVma9271UsjL3ew7A11gx45KRGYzq7NSjqzF5FYxyL4CmfRDPQlPHqLvbAG7
YICIYqAEHXl4BTo9RZUPTOxHKJvJLsNhGOMqk5RKyBM2t1rnb7hE/j9oTJi3t2jJoMqld9jLoGyT
yciSxqZ5A3RsnP6t1XIFkF0wdok0Ib6LbYZTjTwRzlfB5rc9ArUutbAGZbEPr01ajcIC3wdYi1va
3y/duJwiyLm81hcz3MNU9QIoWqvjxbPalpxS3Tt7116p94lQEM88isUAZ8ULdY15ikNy7GrloPxE
6mf6NOAL1TxfyAZVRWc1WfDKKyTLHH/H46Sy8P6iAO7P2O/QJQgL7JnTxV6pqatvP/aTnG2PIDgJ
0TXO0bhVEngA8XXFgsnpY0z1189WXa7dIZMoKV7GzqZQ2oXpm9qPA7JbfYL8ZLmsJr/zUwz7kTbt
1z9QZmfeT2HONh9x8YTScPGYjoGqIOZwhEqyJ5kVGWJvyuImA/HmCGwKVJ+dmCNU5lGqkn5E9XGM
iZxNLXmTihbHMAPIawS4yqBryJcDcZdWntc9FiVn+8ByrD5DbBQIk8TB+cO4EOfDwMVNrFoduDjE
m2WxspNwnVQ4Do0hTTRExiZ0MA2O1Hkj9GQQLRq6klsIVpj9QEIciwbBLnpgrZiV0x81H9KFRrH/
++NlcIxbl71kNP9g1NOl3ex9VkBbFd8qmMZI4tXD88ifptedbboCWVfurzDkCSsAw3UE9OcHEt/a
zaFC07dueuP39yjNWnQML31maZRoSvD84WsuzO/lxaaNJxLVnAzD9g/r+Z2TWPJumaQNLHA/kpkB
P3rPxHc8inaMb5QlvAZq8ygtsc1pFcU1qjAu0XMffKv6iIjL1WxYXlMbZXuLbhgs8ps524YWQraf
tjbnZQPza7vBRIr0s8llQ6bMiuW7ZVmiQo3c6mqIeSAJbh2ZN6VslUCIav2v4zmFDwniwLujc/nX
bJURC4Ktw3Vv8T3tsMzMXM/MDcwtRStp7fQB0nKh7p4oEthFT2VI+E6Rt8uDvm63pMhzEENTz3uB
ml248hE88X8Fsw1EIg65lS0GlIMoyY+e5dTf0pI6Bo3ERbbIvosh0/iJgn0B7Y4Feg7UdepgHe+4
QQKj0YMIo6dWT9Ckg6c/n92kWrFQKO7ab2Ha4UrCvanxhYPzqu+jzffhhU4P8xxV3htWgM6feTC1
PHoKo1p09aUa8qOcGlVEdkffrul0fHk3/SfTJkdHJGZG8v/3j6mKAglrdTEfAWDS/uILJZek7+0e
C2dmD0hJsz8hWO6iwYO1I0JEOtsZ2SbxyhhRVU11TALQrW+PghUkadHIPUXsOgI1/90berroeahS
eANVHiw6yS5VNFSM0EHoKYbZXk2sBQkFCcJDQG0h+cVqCXi+ApTRdIn0uKd8X36MJhz8/ooi1zvH
c/o1ALPqhP1otFVmzLzZgu+kh6+c5ndaWu9NB5aYQLLn37CvEGRc5V6ylb82IR2O7CeB5p/Q2FQ5
e/SjM0pI7gfAGiR7UR01U9qEoLTVVMRwu6zv2Y9um7ixSxvJb3wnTRu1Vu9gNLAQ9wfPnDJbBdod
DeHaS1QBHrQ1hYlyhc9mBAYS660+O7r5/mcQfBxr3m2dSzC56sA/bDhiQ4t4p48SWG6LmF6XOsGG
TrZte18Uay/xlLNQIRoz2+J5aVlkF30IgA40zLxBU0I6PC10sSjyeOJtBr3l2QG81ubpuXiJ7Fo9
rKaLiTuWz5M/lWSJouBYgOmDJtPTF66959VKxCJJtB3Kt5pSLdeAywsFeDHS59e3R4IxT1GG0ox6
uWdb5OI2MDP+ZB4WMwT4dicevdFxTZyQzyVSYpecU6ZCrwag+YCXQZEojbO+TRQDD4N6I3/sHzKF
S8k2ArWHLk8rZyNwWHIvHPjGqqUIdP/tAWE4RklpSpu399cjjS+B21lb04bDTYH9FV3wVQTYLpUx
ADzWK1qS7nme+4RQCeeACvuuL6D05ZXvppkTkK0uSPNTWTCGLPSZrE69K0/ZOja4AMS/q+ovk4tf
s3BFBAbdI6MwhUH5Mbc0gecsSxArMiSTTeS7sKhB+q34Iol+L0HbkJxOX+P2J1MhLNjxUtZ3rVIt
MvSDKXfv6wkDU7rIRB3OR3twRiUTejFarAUGh5KR+Jd/wRrV9HIMAlanENWmI8Ooq16rlKGBSN+3
pHg1pTVhHTQYvcbQtZHD2xLzRm2gwQLw5b8xYAimsQ9AAqGyT97VzZnnAo5aAoZUkL36HUa8JaYB
/N9f6062FHhTiydE/XJR8w+duUkvlWZASStqRbosZHvr+1bqBsFO4Lxpa9GSk3RyfPJr4axCE4n7
j9I+hz6DktNLQAEMrp4AM/x9u2O6sbMrRcP1pCnqq07w54enDzmejLqBTIUqYdrjfeBGCm99TeC5
eFULYJBtulPWSkhQKay2auzpzC8CyxUsaGkXAVDjFiAdn01Ovjw6En1CdBp1wHrA+iZ0EoLHeUuE
F/yznq7URQ0t6WNQUGizQA9M0stCsn36LMC5BbrH0jNQQV3L1pIQMJndF91HTmUL/Y59nfd5WL+J
Y8I+/WEk03yT1uRYSxXA0OuJGz5IHySA5215CmXGJN15lh92oMofB/gGKd1KEAAHCoG8PAix79yM
upHxhEbm8JwrV4ecsPH9rF38WlKL9vP+OPfl87k+qTviA6ulBBq0ti8P/rz9iiTYCJFz0h0U5rWA
R34cOItGzJA4d8i9CVNU6H/7W8tvUsKOLm8wt1zzIos2pSFG/lB9N3FA4L3TFx5a0UusxS1z6m+w
VeGSEBgix7CT7lwM/Y/PO+AqSDWht6kEDW3L7RuXqPddIb21QnSU2r89iJYcMfNYynNZ/SwDB54c
ossB18+bF+R1ZuPEkWt8Y28dmfF2a0t7MsxX4dFlemUqfVBU0MXXumoIZKF7QXlvMcWPxiN1+UcY
V8rCEzEpHid9m/C1UdESKRhfLHTx7HEayS1v0UUhmbqQ3KzFmNGY/JxPglwA98+6N6qzXlp5qaUV
mcbrS74hnHWKX3jmw1hjvongBKIcpoHShblZ1TyRIYZCmA2HjQIwm6DLvx1dHlQKZfNEwuNuTPHX
KdS2h7vcXocEYtdR8H4unOzxOb8RDTcbqrbHhY5USVJGB+xg5Mf+bQFXHbxljkHtzPeM5fRuJS9g
ITgrSCio7F5xa1gPBcVB6xNMylDAgjVmuVs9zPU/+gssPymO2yb9Su+r0GXZ+sDPk/pofOd55ZyO
FktOaAQLxfVCPiVUVXLfIxFfLi6y0fSG5yZ9GKuah7pFIFX6QLQ6+yGJULWrdYPl42VS8V4GeC8+
fTAz4yJSfyVm+NYPLhc61dkl+/j+IkSLnoXDlj36RwPmwl00/8mccgi7awmFGQAxgZYiUaWXjyhL
uhyaLMiJzGYwoc8T4/8c817qh9n2FucT+wdXQDrpZ1DbS9Dd2QT877vIR/S5yrfNqpbFhfkVrOxU
QYjBU7VyGaJNuvWJshHIYkIqL3egboZZOe+E589McuMwOiWFjxjdWfoX5iLOac9pos64TCP3/3MZ
PSrONrGwkI+QtVa9seA8gpLdEe74KDlJv6HMB3uh4P6Igkbdc583+Iq/c7GbqZy2yL13xtjgYhJp
oKh/Mq6y614D2DqhpyZR/Rlcuh2e6E+ghAnAQYMXLNCb1AA+t5QqhVP2J6f/Tar3I0LM9AU3PgTV
eX/YUfMh8cg9U479s7fEZ2E65SN+kREYIiP4GLZRWNr6Irca+gsvOi3u2fVmUpwtQqsmYYeUzMqY
q0ZGqf7vSjA09FYzqQCOEo95BPZ5GBQOMWUHw+YmIMVgFTtZJhFzY0gBWkThSJbtZI7ESNv/2Pb/
ygg646TyXKORScj1S4eBR4ojSr7Ec2MIl9vnfgoGBZdyUCe/GO0IObFNawSE/jF3uMtSGK3YSwFX
tRHQtBldBZ2ls/Ala8WvK+NfG4hfUTt77zeiFZpYEwZXvRz7wJygksaosDSf7gHcKYe36lVwKhqq
aYD98nW/GiCTzRu4AUNWWMX1tgNVv97Oml/e5WcnEltfT1j7SXoXhIEq6dLRewXGMtkyOLJOtKGG
xs6qTH8j6YkNeO3YYMBo7cMCqyv3aV5LPDDBjmH+FqYss149vERKKFrZkQdgWQVR6ndo7oJyZT4N
0fjkMZRPPpo3SZbfSHV7O0iAlot3lzHNs3PFqLQ75XRWu7JZa5xCDf2H0FgbM1AbCKnbSyfy3FBA
qnkSxoXJFJVNrI52I4tIGsJ2xXHRyBgXOmJ/U/fxuHnFEcvoPdqca5/r8yVd5lpn3H6uqJrCYr9r
nejqYd7vPCYzTANHLESmR3iUVG7bjq96GVYuSTNI+5rDy9+DJeiUJ81JN1GjqjClTK2JMYKK8y3s
AsdvJodg63dzx3El0Hu4WxME707Pa6KQpmHz5ny/6+tlaoiHQCnTnALEDDyPVNfWw1e6krBIX2XE
Ugq49JzaTLvrk1f3pDgHv6lN50nkz6r3PC/1Nkdb0f+t4gH/um5QKYDpg2TvLjgmc2I3Vnh8iP9d
/ba+5pTKLQHqSJcpLHIFbW9G9YeOof5sCQeS4iLhEQyShJCke0ucDq+jbsInw6rOlS23R/ghb68q
vCeFMDEeP9aqHjF9mppYUhEJZh+oMRFDQsSTpafHlu/nlFTmOltxnDRfOn4sVBLbKbq1GZZVJ0uY
TusjgNNO/31jXTrI27IZyAYjhqS1lCRewqd7s46r3SfS4R/J4RPhPFtfVTsSBtRDFGvBrOstVLIK
gt4+sqxewsZYdDBWvFLNvSGKXR4nQ1ZkPlutW+ch1hkThc2iJk8BUXTiMnis6a0cjpn0pMwqJJde
1zsibVFuuh6sgdvtBnkSoxN87BeBQI8wOMG+L3lWebjqXHoxIhExz7Ym1poDJ+RbvrbeTo88Ear3
lwIjpZvPVjsePMauTPRNsgXrGSI8KNEKKfASnWDsjnuqeRWBduuihBLcJJts5wVyWi5Nl/Ei66ku
eF8PvHk19+uqG0nZWXPunU/Qj7D9gmOsyFZAiBieujGDr2ibS5hnpT9p30Ap150iN2J7M9zaV85X
KqhgsLvs93ZXQ5/28lxHNfe4OshQD98ro44yWgaudOWX8CkZKHW9fBXLKCTPONvHNtkbv4iiHLH9
LlTKpQCHKqujPPjojsfTGwsC6V4Ad8AwCQhG4r+Nep0ehB7Mv4iTstSTReWwX32loh+bi7kwR0LO
Z/KcGschuZbKFmIHrclvTNbHV/E0i/bcyoGr5cRHrmYiA75we+rw2HuyAhhpOMwILQ0DfvBBpmq3
0UEjgwwZika3ClNUErrvAFF7dTw7zibAurDgTDFZdECdwWocqSfIlsPl5jfP+CL/nYr2cAk0SBxt
vvWYcxVsjRmvfhmJOhAhHhp/HYyZBu+JaxyrP02KO+yxnvU2FyYhszSWrG4fFSAFVADm+3WWEo4b
1cIIRQvbkDXIEh7UeKC5UHvqB1RSbKr1HTt6AvbrRQ3dnEziZa31Re50zHt1JFOxfVy/Xn6Kf5Oz
6n62x5LW7zn6jDdiOdKWafp6AtX654gKinOQqj3221XzGky5Vp02fQ+xeo0M7CNVoCLaV9Ba1IZa
oaEQuMIYI5TlO2GhAtKBWg17ArA6DwePB/nHHZpUJSuVtORp+4+kTUbumhyvnrNS6lONewCFZAvC
uB/Pplz9RWS68S8jMr8vFaMXHUUL060zXocsoUFkSq8us9aGKCa6YCI420h57k2i78nuoybCasXR
doAKQnqJScXUjhhJxb0xyQEMSDMLQfcBPn3hjF5yQ4QA+injm1MR9pB1hNR+Mo8SzNsl1u66qJ+T
Ud2roFDPIubnQVjBun/+jHTml7ClkKHISgETKSoDBi/S4pVd66Vz1Gz5BGSvm+5d4s+t8BEd/52k
uT/9drg2l2rHYX5hscApKeqMbR9tTLcOq+BRP1Y+IpD0sj2KA0FkGomq6d22puxCkvL3pWyOUzqg
71ynevUtYarP3UzygUVNFAeegP4o1aKQBIyClL9H0s5is1eNFMpZ31oQPXZiA96RtIRtpg1C9rNo
dZEwrVSlLSm+qKviO/RA+ZHpZQuPg9r37Ly6xKMdAXacFGb92RIlqAXYna1/GM6/iFYTxYxZS2YZ
Fn6LXrB8uolix6IfbnfOIZLWGNHuKSKQzO2cKwsa0Xyh4Zz/VO7O3xE1GGtmdrtjy6mhYFWjjhgn
CQYKTDZLvfcIapjExQS8/MzU7VpSKHfhviYI0CM9CZDsj+H8m6ImtzAcaUwg5L5csOr0ApMTs7UV
RB8HJnLrmzYe6dvuRjN7fgAnjgBoCblTk5XdQLbETKAuNhPMjZxngpeXq5E74yCQw133BFsBBy16
Lg1Y+QmuiNmMug2PfzQqu/d80VfwYoCPtwF6ScUd/p0LfTpInWIJlzKCIq8jpdDzUHebUccEKFTr
VKa84aC8oRfzcZUOHKEOmMs8Ef99Lr+JcJZf/p+ZKk5y5lADyZ+PSdcfCabl51we3VIhsf22p8tI
iWXdl2nE2X98RVHtnyCQtPiExazC5TGlshEGJlZwZNdGLh2kB5ceukfHDMPa7BvNer0GBQD27Agy
V1/SiPLWE0u0o35bIU1Vl/12jvgJlO7k0MyqEr3MbuZj46I7PAPqhysV3DyvQ+wgczuUIVg5BmfD
7efNXXEoqc29GdtcJfOwegZBBxsyvrkoYAVMu5RTCPmP+Nq5KFxdGbYSwZYixRljkMjIjh5a/1L5
Nrdk7ovM79VxUgJxdGm4faLja5jP/mVbYZv8nwlxIeDWPEdfE5uvmD47MfndQgc0wh1qBDF27Qqf
AUwhorgfjC2T0xsAFNQurFyojauPK2N2NxWSyUe0ZJ6D6mR/6wcAMwNSQXBfEWb1JB8MD1raIZB5
kpZ4+nUHfL9SLnxDxe1c+qMkOuChSbPvafiK6i4/ZC2mXitep2N2rBvm2XTkhDDRgcUJ8jssdmp2
XrMeFOAIye34EVenA6rldX3BJRH3F10FDih4sInl+rijZtgFEGt9n2P+a3lBGBP8ovMbkTeJ0yaH
LanEnzCXNa4HOeoOV7JgLQcGbQlGI/RV9W94U/KcFzJ38OMPqAulYDdWQSDlnZbtd7nHHM/y879P
vA7A3WJMVYp/5rieOQwy3KC8VhM1kbvEaHhrdkC1qYj/00KvTJoTsnoiXjy9IFFUCHbPi4bhcAu/
Nd4iAcoOL6irTl8b6Xvy+IYvTW2XSY/YogFCV7CFlgbFVL5kdfzyFDQQWq1+3xjhRAeyq/2O58A6
2IyroQXwIpxXJ/O9kmhP9rBwCefukQLE9WtGj6NrSMJx5TPuyu6E6zoo764oCUCcMMx1JTJ8myvF
I4H6vWY3tejEcVY5O2WOFqzV0XVb+Qabwb6qIttokirG4lzlk25wNI1947HVIn/KZjLIlz1R0vYd
NUuvqt2faLheb3edqYY00Hyg1HJGcCKpiH+6NwIrp3IUmosvXc5NPU23sj0tDecM4dNAwUhryF3l
B8TmUfEcHsZaPe5eiZjsGQLYfWJqXyGZ7T9zY0/tnJu6YlKZ6SLv1Vt0Kz4RIhqLScFblfdQvypV
ShR9hbv0GwpJc8VlwKJJ4wsO2THb7SMs+MS4zxuQOiuqicn8kw14mzNxe0SvlIYKeHBLdKN4Rlwn
y2G+G+fdstnCUR6+5xGG4Zf/rjCtKGe/K4vic1ko6716xkIKYxRlWbG0M1q4MbQpR7DIcVtCUVji
VYBZovhpnUWDG/6sG0qsZLB0VscPXDd1oJ1R91LeVaK0NjSkAZGtAIziodEq1qozMmmCfS2zN/6Z
RXsz712BwsbPYkTLK6hSmJYdFJhbPedd6qmFMMxgIKdF5Qzg6+klQwbWLkC3sOIIRVJ9vHwkAZQp
35V2Ql5Elv532YKWcnw+o1we7mtPpGM8QkUk7yvxVPhPDo22QXvacNFehFEyBTSt5fVujpUiWuVh
uhRItfHhnTdtmMLXV5qIblb75i1caLXQBSYk+Q2ufLHYFkIjSBmyUFYUngQvbwVYwk79UEQW8eBK
eddryvaauZK2CAPTl0x4pj1gDyDoS/Vg9GxD+P3w6QrOTEvEN4PK5af8tteypdHrEky3RXMZnsQ0
oLxvKMql7Wji1xESO3EUha1u4Hst8wBkLg/eq9QuWnxKmfgFzXBPdwG1p+Vz235WrubHUCXJhzhO
dA5Ohpv2Ff3oIDAKKAEFa9la73v48faq7nJgJlmgxHy0dIVC8DtC/4PUE+xvug+EfSYpQ2OhDPro
M6rUBvbeKV/KtO/OcZe7zPLM09FlLukO43L2tSiTDOJb9NkKpJTmTDPCdkDx+vk4zh3C92jzcRi+
CQcKXmiYEejaQi/a7U8YTCESITw6ngb3CVFgqgJoko9wa1Y22s5l5wq+5uVzoEpMQiQ8BdNC6zGb
80jrs4BpC4jh0QdXTu4HJT4XuZII2ReAmW5PYG4oATS/q2wc6WizvKvlp6XX82b9Vc3KJG3qX/ct
S0Akc9JkXCsEucZVbfIbILNrsHiErJZSs9GHGKJY7vMx0yeSh2JfjBwwo2j2kosqV6M0zGtBdl7l
2YYrgQ0nHz+ItCv9qsiua6gd2oPGxoQECbjtUHbMHcaNvwNPy8PbP54cD1KtyeBN5F5CsSz6RNZI
gcBUtbXM4NkEnreKCjEiaAy0RkA7zvSpe2lR1XX5L8amVnKX6w5OYupn7NOyi3lFvKpYT9fWKfOA
8AfLyBhPHr2ZM0svuBUXFpuMtsLf6QdGDkH7xE3+zkQ5RLMQ/uVAHKK+rLI5MlbBgJd+PpOEjG75
jYODG7oFTe6cGznbVupbi9H0mtWxDUO3WJkw/mUzNDNi21A9vMI1lEZksTRXcNkNfWl7FjKKrfFM
myauna7nEbbR/wGIEE20olnlKftWvOVme4CrtRtBHu+AvA64Z2ai9R8ERxpFxzz7b193BS5Owen4
kWyrGX/PE/G0UjYq7xHvzPjshrH8bn5i8DGpcVYDL6Fr0/MPVqL0cK0O4jeLfbXN/Gx7J8mwYfD0
4JZUDEsoG0S2Tzguq5w2jIJ6YVycsvbw7n5mWvApZieoW56WFf9wYdDkqjz2FUp9GcOkxRY7SsxY
eBnzAUKP88yBDbaCEvJItekHn+rxPxHWNCKBKv/B1YF/lCfQAZY5S/CyCuPkZILJqF77OVrULx0H
oUdZ9iKHaYPoUq2m9jEOReX11YlYsyN+3AnKyUAFBAXdYY2qkM9JKBXQJPfGcjGymTqIJWSoLz7m
Lt++4zVYSPeE+fkAVXdESP0ickvnCqH204s1voKfeSyOyz0KVWPqL+otMy+4mJGHh6kx4pyV0byf
bRmm9nsQBxMN2ebRQw8lXUiRV199e0xk5qkzKpNgkM19hFayl2b7b7MQppILF9ZMcZ9BFDGHYj1f
v/8j/yS9bc8OfVkW2LSzaYOFUdjbkD0KuSifX9cGiPrlfmyrKtHhzv6FTt8SrmYi2XnSGoPtdIA0
Iebh/I3w6CaqntYg8fn1+3ZPAQJvJTFOe8QMn4JPjqGwvlJTeMLOJ4iKH+U1xI7bugqSE2lTDW0y
f11Bv6Cfpy7hPL8/WFVr14nzSdkXAxQFmX7ZK/x07luZtUzlNbH/i9kbldg9TF+YPszcaxeXdmTB
qZKxpXrXOt+Je/VQngXgV6kqIAd9vHNkcFJzk+Gj8RMC7q3HY3LhrY+V7iVqbUmvoS+uBpV4mN88
aWX7Aj2f0sx+wz6mkvG7WdagRvTs1CtuZvgQxyLmUCHRtwV3GFx5e/x1+jyhmrceHnZtFugBF1LW
0fWEwzgCRaRayPUHXwUSnGc1M8a7tBFbCbe+hRWPsFYxT2F+trqtLAUos7WOkNkhMXjL8A0vtqLe
phxrL0HxHMd4Nz/QnjsQSlywNzQofQk98QnaGw4ZXOLg3ZcIoOqP4NXLKTQY9O7HoQI4m33Hp9Fh
gtxf3YbWoZjnjli4+xOInEXtxP0DF60x8YoR5qpmfXL3jFN/2xN+8WSKG2L2fMH0VPtKQuI0ZkXv
TLbui8j5V6r8k2VOmzIrc6oOUXI/7p5LtXSq+/FHwDbznKVGvpRBi3Ja5OGcLR0EFCRSpf0b9L+8
NqFyC/CkfIJ4hoSKgWDNcPYh3+c7KwfTdyRmdqM+zFlIBIg2ARlPrW7exq3QGjxGzo9UueDSdAuh
G/AlKOR7ymSnYjTVlJKvdUtcDOJx4ix6MSsS9Pkgns8JTuNoN2yGJzc6vqrkGBB0n7vGhOj5ITof
x2HkVCj4AYefcUR5JDOGOVx4Fr0c75WxQRdtoA/pDfODP6pja7f6FOoNZdmiLmofNo3pYDmW5AQp
LNh1mGS5Ob+VFjBteMXMzVf4yKhVpLfoe3aokg7vLcgvsaQpbiG134sW8vCMQxFpWXyVn2IsaM3W
dCwpYTTVi5FJS1NBx6mC3C59i3n3n59df+5o0MoZSPGnZkSKr529Lph7ugleZfV+edQYC2q2aFBO
+Sv9qfur3r0jbF4lQ45upJrJNDcLQtEnai6J8n5OLqg30PFYQXRGinpTdi3fkp8Z6/7C+ua35NQV
0CW0IUSYbpvGNd4hqcsn5lKX4q0MyoDdN8PKg8JuaJ5yKvIXsQy4vDgcgrjO1b9h5O4etVRT1io7
PLiqB0snsqSSsV0ZEr38HibscrpViYOzO8pmXKsdoNPCGlEQ6/56MXbLCoRog8iACq7MDWkLue/a
NNyotcB5xzcCOlwOI2ZiOIYCKLM0sk/fdCgCi3swTAl7LlAel6JFm4wg2EgHxUKaosfXqC45QS5n
RqAGbfEFLiPzVQYDnUEKH3ajBxfSsDoB+5Dkh4wAb5oqL3XOuRJ6ZPbQNUg1Sq2AThkMG4sFUOUl
dJTVm3NP11DY2twoFp21QBEQPoAWEurTPZSUIVz9e+/2GCRo66TLIuutAMEHEI7fm4bYrK5TJr0p
th3QQhZXyYZmpkbs/N+0h6e3QkSm1n6SKrqqFtd73hVvXwbz+xpC2GpfPkOXwtUAZP5+X19QHxi/
L2GobyN+xUQZFhDlLeaD6wLjHoZ5geB+zK+HvVYInGEa5EwK9WV97yIMhvbSjJYObYPApWpmHBus
GC+pApEu1I9Oodbv61pV47MC/Veu2Rp7UY0apQqTP8+zEZ5kvNRb2gwOgJP3r+UBHbURB6kyGo2r
Li/taAHQSotifNS4TvfPXdOpam1RbyvU7m/QGY2EkqfYvGjRksX+Yu4p+ITXNQNwpyz/ZFz2ZXj9
hukXKyhkfKA0p8syoPg7JwFn3uoWyPoXBPaw4x6o9Gyn5i8EoHZYB3BfFIvY6ERsjuyxF5qpVH5c
mGbKOzu/U6OIdfvpE61NRE3bqoqlpwJAFo0Vsqgw+LprXa6LmjOAacKBTaCeB4E/yFE26DZfmPEh
Ua6fpGotgjSQRXtEOTzeqRYe89RyD3sAVAf606owyNgnzSMI8gnvN0RUoJ5Hw39m1d74w2PH56AM
jkxiu1AsZNR09xvJ5yVsHbkbufzq8q6NaCxELxo1PFk3dotyTviu4Hmu5bksWbzCNePFA4mvs62n
7yhV6I4FEbiL0y50ASF9700/+uArSgE0sK7zgs4L1iY+ba0CjGKcpAMsFD5WPpmKYyTF5PHYKEQp
hPMVQEQEO8hbX5udgWunnHWMwjtETjYHz+9ug4r2xvNSt5L58FOAdT2IaRUIYSbmnZIJIpsge0b1
8hXklcCmFBD4ZZSQncqf1iKT+o6cb7Umgm6v/cdIHfgy8VnIkUUPzTBNG2akINKNE+zNmN0cVA1n
O27r36LAhKbI6i6m2r9W1mPQqvM+5l9/CFghbnzhZqMGlSLMT/56S4D9U7Wb2SEFJDb0BmUjSmMi
RzHOsYn/O31tiYpU+w0ye+KUWBwFJVmERTzNoW/fsVFuV66xLvC2afj0onp6a3Nyr8NLrg6ioDg1
HHCI4GhkBNEh4J1+LT2OrkdkPct0Dy0uwVBFlZvDBAm5NlSAHBLJH6OOQOJ7SRr20Urjl0f0evF8
5h14slHnJGO1jvbmANKQNeHcnpBrnUcd5ZLTnhkn+koDM5RaYoQ5N/C6EB0L+FRHnwu9VJuvdEtf
qLKBPNjDerwCWWRJo/FmEG5THAMV5kI5VyjV3zHatDYQswI+X7JfWURxLI5S03upHT7LDeQwL3b8
J0dSd1ohoyKJcLN89GOcU1HR/CihY8qyjRYiLBxj2WMum11PiEuQPkoNxqzK+8vvA+7mmNymNAPK
JhEQgULRWZIbkph3u27bmjrFAw1rAbP3uvfLvCvZO8WczlzqDIJix4N2lm4eUaQhFwH8lYtrdmMe
0OdWUiE8vJkeO+CftEVmWCIjeHcisWvzkL8x1vA9u4a1mjDHOfn/owkp96ZQ+T/kRJtzrLXyWSSt
D86DSGP31bRqhEQBaezOkr1F6GcSPlnN8XzDIKyGA4xLhZJ43FGvZjXfcMfHy7fnZbOyyu9322HH
fV6Mq/PhAbQHSq//K5b56S6RmejBmzsNE9Ig4uRJVPtSx72XprO//WE+/l4zWv8z5TwPxWePUfN7
cCiRE703/5g9Iwae9btuIYSfKdpLIDPJYPhNZWwvgWI3t/Q6T44scV9HDDsgSYOWWAU55pNx/Uni
WWluH08akYn9kbXfpwMPfCSHldDttXr88fQgPTZDhzNc3kD0yIcZ8+FQqCWSyClIfgnCNCzE3uF5
I5WHOfvvgC8ekKDCpd3vdETpNoNZtbaQHm0VXJch1mvMHVUDYrt81kXRMbJ+ynwVSVOBXlaaUlsZ
cNfIQrxcxDVyB/uNnMR/nnMVHBADR2uuTevEs3oFGYWwqUG9VQqSHQUK2y7k+bfl0unhhw011LyZ
XyR+d5vyxpTWWWN50tjTuR5Xxdnt46h3LrP1WOrag6iTBnkbcgBbKRo7uhcsQKdm3NiVt+3WbUkn
DUpg1Pu66ejaeLwQyzdK4sTxQCDvY9a4iUKlacxKn0THw+GCxsNWNqB2a1Pudq0HAXLQUpXQc6s8
cq4wuKoNxFxijp+1XcMDZ/NIKtdAHpOPTTcepCSbNuu2mjRQ38y/6QmUOgWTq75Jmg74KDIql0ze
B1uZ1rJCWOtjvoc3Yqz4ko7jLl0n5pHitG4n0tVNoYTlskUSWG/N78JfLhKQxTDiWY/D0xwVOUCi
0FvAGZ/bX97GnSdTyZ6nnhWUbrzsn53PIF8Zr1oBWcQm81V015YkKrczSVxiRI6NNU+c5oLyyptK
v8DhYzi6ro7XveL+9EmyyWCiHmhw+zEYLGlBt6VDpyQDFvLACO8CWAn4nMQqjZFbVCHMBegZGSaY
ppJfs4iUh6tWNnbhDOL+nK240jBkmukvvjPY/L0O+Xw53QSp7Vdk/a+9OsWN3XgSpYRLQbv4e5lx
t+63yhMcfuzqvpBOecPXwBrnMM6vmmGKOntAZ8nADqrUb8ZwoHta0eXNnkwNayQEzZQubwwG7460
tjJ4ixfQcDnI+Tk9fVvD9DFUlI3zeSCuHn3M8XkdNmOsig8GrOysSPubR0A0N3dGJKKFtSO5KJWD
ejdh/D5eErrfhXw3HxnOUFfqDWqtAB8tHvs0TzGvOS8a2ow5mR4oVzltkluLuzPJ268tPvXr5wY/
pqMePnvSJHYQtTvZiZOk7xOLkYdW53HASeQ1wmnEdVvV4zkISfyLN3Jow8FePjY5OkOFQK7pbsbL
xyIoPoVBp3bFmzD9LH6wuVOcBXOwFAbkZP6v4EWFi+o3xsosq+/1715V/2mhAwYchaQdPr+3z7CF
YqFn58puoqlQb7SXGNturFidDSxcOjbinMXoZleAtuB80zUrrMa4VwMHumwbuZ45os0V18a67kHT
V0FRk/n48m2dcfCG2KnAhjaqd2QABf7eaybuCMoJPnFZJ6UEQ7YmY1Konurmdrgt0NkLR2TXfVa4
KneBVmTTuQWBWiiescMy8vPhrMU190tqKKGBf/k2nJJRz1QPG9b2JqBH0GKwFCqeCN6kyT6qLQ2t
ebdu0XZz25p9DBCOnqMvkwjwfVqq9p6H7W+xXDcDuMfJvuX7dgqFKp6ZJzEYciV4aXZvanm41cjB
9lMaMZKMskuMZNvJjEN6xDVSxwob6AcoBEMTrSb2NuDAwkee+6nyy9hpq6CTNJkMgTo2XYzYN4ol
uS4q5ruuGg+4ECCZJnDFyvI5m/pieV0rCCEaAKzSbb23E7axgWSAjUJfdS+66uHyb8LQvVHPxli1
6UzT5xyWzMcqvXISxDeEKHc2HxjXOyhxbeAWnrqH6/TzBL/M8UKGQlNNrt1kE9mC8PBU6QtC8sC3
Dmt8pOYdjyp1AtA50W7UqefGVcfjkK2L8FM+3CsQeFBfwv+x1msNnm7nQ6LrpudsEMo0Ugxua0Mq
yvZWoFtsLF/6KGOb+eQKIgH32bDQB+MuWt7zUHWyDyP+Z06HpWToq5sYtHCB6Sv4V23sAZxnupZs
Jm3wzJgDX5zQFRkfALUpg9TGPG5dBeL997zuoNZCGUx87PWw44nO3znRSd6otSR7OCWStnp18i/h
5G/kl5SldQO599PmYSYqGF6RJ6U+uVvQUAo9CNLbJ1q+I2rE7jdqDE4BUI/U+THu2JoHEaITMYEi
qjUQfXMPSHdBASLsLg7VPJsvg92xCeTA59+Js7ku1aNBlf5j7NOGJRqXqgyUXbvs80ojFyABc8pH
C4fNX8bIPwg72y7GpgcOfax5HzIGCsI/zZSIq/CHi90rxVixsw+5RbgJtPRPGusUT4tLSxSHtDzT
eovbKbCzEMbsPPQ8x1wu0kT8H0cUX4UZF2fUqhnxoOA+CpGT0ZEEMuI7AlJ3AKUoghpyaZH5vFx5
sBKwMh1LVztjUOfiDyheCc6KOZWN4agTjNuJzv/ooS0Co0jvfQxQVY/ZqQfU670HdNd+AeOUh/6r
X+30hyBVJPteHLl6CgzetoM881bv08DbLWMi6FCozZ4gs7DheMSP+xXL3YRcZiCvEbakSLlGT9rU
EVrxlGJENP49wsGPOHId/acF/7qu+5RQlkcQ4IrmGglpRYx2PsnyzLNdmuWeyFWc6ei/XnWn0ZvI
orfY2awW1C32SdY8GSaeclAhLL+H7ts8ebo7iEmouwQClAvzTe0GCedEwu/v6WT/ts0eWiLFmbdJ
wx/8F0DS1dx5zuEJEzMDcxqxreUPRKhU0r5V02FWeGyNO7s36qyNFjcji5OgBZAAU2abM3eDkJYM
bYbsEmzWasgp73RPxRC2M+rIrwTLbMmbwN9in/Mq90xH2rbuMylTny7H24oX5PCG83YGnDuZ9EV+
tLElev0N17mEmREXFOfdz4Rq6Kl0Fg6BL9k9Me3rFvOHv2/JLxDzQJn08oioP/dsoJ9O7DOPM9vK
ftmjWz/ItrlJobz8FaGVeKv9lduCNMfunXZKV/EdCDiDmF1zkjNJYwP9qfZHCUOt5nqJ8O9btBfI
MVx4xejER2C2Eq1B/wRmG4YsW7lsaP1UvEb10N6Wr2Ioyv8u8VcBVtWABFruOnmiDtUeaTHzYiG/
A3ALxDr55nfxn0WYi5nSEHHonATL0+l4q1SGTp29IKsKEyH7LFpTl09tPzR1gGtJUNDcmTWfxqUG
39naWwGlHDy2bcZDvj/dmdsmi0Tphvn+LjQ+Uz3+pZ6HD81lhln6vgUzzVb0KGXKdXw2jmR7BYp/
eEouOlD4hlNbAHOapAjuYIcU7bvVRMjdaThwS3f/l2dEdJmX+dmVHTe91q9U9tR2DS+FigjlztVR
Rb2WZ2FUzZY8b9slBmp6KAB8WYDY8ORVKLsME2XrJJEiFFUiIuozXj4H82De2TgghsTCWCeDlAfk
mxXZvBJBtMaHkdB9GF25JBrXkCos+AoW7j0gYmCibKksnkjdMsVcy3FOvxUrHEp1sQWziwitlt2r
g/aEfUyd4lRY44vicL16Pj4jbLRLg2sBWbPXh8y2odsBrqlKOwhG96kFkoS4GHqY0DmzpQJYUivy
xKwpTc5z7KBK1c7nztvEh8obvi6rQgrO9MR44Ky2aBk3iEC8fmEjy967k35cwBDTUdokj0OFZxWr
hXS5DdL0BgRE2TTv0nLsPYhuE9mXvlGL1OBR+Y4rmNb7I0Q6HgqSgzSt2xPIn24zXqJ4KfFAb4ws
bzC3qdYRWldIKT5xDvlkpopHkiGaJmH25b0ZZbVyyH0FkvyNTYs/Bdqk3M8E63ocpU4R2zcienx/
BhtapYODr6HDmJd5gTJkawsqvIAEjJrbYM8OpC7XZxO4rktA5zwRf/Zv19AnEfkFU0PyHjwrvh9i
/r1ZA31IGXM3XqdwcGJMYl6D3Fdk83GYlhuX4KK5RlV/J860YhWTdhPtj2ywrLgBoPJEm8ls+MPA
FyqJtJElnl4+sfsNKfLcY22R6clHMOQwbDHmyc3wrz4xR42A62VNc8m2czLonPNi8IkLo9KvD8eo
1nzMSduKQMctpwwHMxTUfxPbPUIlzDOvZYfWhXmaMnaRN8uoHyGpPLirlqvoKEYQPzXapDu+930y
delyTGQemuAcXS0MtZWVAkfLoqi3Lql5VafPf3qhmiFsg0r9CCAkCKWlrNby3sbOMrggUcURGy/M
Y00bzIHQeRi220PXZOKmqjOUxtziQibrhOcGbn6TiRFJpNLgrm4eqhnurJ4CC6g7kTL5/I9UseTP
vubVh7c3rxMWXW+XmOCCFdDg4Q1Mr8gYYiOZqdvIajP2wPFZLO9m0WBjZiuG9KUyoalbU9oHr5lE
8VTLKGjDaxIMdsdrvcIEv7T3xqMtN3E4VjrdpC0ov52g2w1f/spacFJpEu/S5PLeG2dy4xmGnvmu
h5Y6B0mNtoReLkn/Q7KVATbSn7oMBGdWEE8JARtfhmQkArkH9dEupP8cg5dsKXfyR1I4LhK+xm3N
98CwN3rQvy33av/wzTKxbK6UQJrNfstMWHcjNSuTXLz65mAvXkbtyipoVJy4oxtcOqrOpZ1CUthc
mN2Boh5jNjE1BFoc2znux3AaF3kVe+rM8+WIzK32fBXbx+CKZaB9uEiXSnzd2Aio4DWxhVacUUMy
SsPwZmFMf1kO1JzZwpVkLJFnzfQJUJhZy9XKtTs90k5BNLZJGhAvCdt5p3RdloRx3cc78HAA4lbs
dZDp0dohquwsL8KwFlf9W3YgyWeT4M8B9sv6hUhtlD97XeoSpvG5qh9/3f4E2dUmpu4OvSUBJNgO
rgIZpqCvLKvHh7K6YE0fZUg3XjhZgYlQEXY6BQ7QXuWWvK2hiwrYkK1XuY8LOQYK+UKPp2PkqI4o
G1BL1dITjbUoRkHlJX2KnZmrvSqxuSo3aTVNlzCvkXQlT+7wudyW2d3p9Z9dv2+SYAKpS/x2eJI4
1v7xfaygpMNHkx/88UmDSngbOFiVU2ilGJHEco8nfeictIyWbg/0PC6gxjfB9I8yWnO4Wno+Oa1h
LNuDNY5pwVwFipbTG6miS/N7f2tG0U1EEroW6sBbKOf7WTbmBavZfDEQ+bB/uCMPWDqJAqLUSHqw
DdRl6eGCiH0LBc/Yia5ohkrLjTElAwAFDHLhELOfEifQvWqtIqV1VGH9hSfX6MOmNl/gHMxAkFef
0Lwf335fq1UoCay/VHegV+/fAYmuz2ZMiM0SZ477T5XkyrNhpTxWKtZKtNR0Uv26Zd5Vxgrw4YqT
p4e93LwysbL+BYIxBStHgpKgm195nVSQe6rHVl5ZLizaF48wJenBQ9bFyu3vh7afK1e11KB0Ny/m
qPIl9h1FpT0H4Pn2fctLJ7IrzAhK282tifLPaaPb07nI5QScm1pn0+se56GuOVK2q5kN4h6Bn8Y1
5PC4v1TcDUcpxPQVVLjfSV8uqEwwIwG348vAVsfQJT/k1P9dB8OxqGT1/TcMCGWYaFofAy0vwTY0
EDy8AWRHw2Cd80Eip6JL8X75kaFNQydYeoLCYMdekoHN5SJXPM3Z36XEEuWEuqjA9O0Sus4s5yhw
Asiba8eUmUZTGcVUfrj6INfssDnENkek6xRdEPuGzQY3ApY9jkh6vYPNljg+8iY0C3J9U13zzTby
fKwVBSxj1DQFzaPIPZvWqCegV/kLjaz8WeZrgg9PP37id2MyJb5sEhsVzI8SosGAFFw6AROM6/iK
XEfg8vcJ+Yh9JV8fUQFjNu3HD1N/d//bh4ikk6FJNdUr2nkmaeVvQyqCQoJLneUS0ANmAl4L10AF
+GLAplJoIrw+lHdgcHD20gzddJ6Lzyn4HtdnXyU3+THqnRkMAaYwiovV7JkAT/HlAo40TRcQreUN
KJuFYGhzOVJPtWN3gurYyyIHmg0xgJhgwPKK53KO6iDt5xWkpFXMeb5WJ8UQ9x8+pmvGyhpR6o0F
Zs5d+N63rUujBm31M5gTkeTqtIWOFiMR2e9UN9O86DRqisQ2mv3fqvPQo1v7YaNWOOCk5ErVm4qL
UXmGtol1qqsl9GKUtCLqxG/7mJIAJmzpbHA2Rsuq0MykUHC5i9i9eHR9v5qcBmWhB2IUFdJVderY
ECwGfU1e4lrU9yrIxntYR2NoRdBsSaBymytPAUz0pF6WUdz87wVHvUxu2YvvThkP1dTDo/88TPnK
51TeIbdKNCZPv2Mjzv5/mHf26hmYWQ25vZe3OkJGVDItuIh2sZh11Nm2UpgIP0Pje0IAf43duqBW
Utl4K/9ip5eDZuc+B7BV2CRxfN6ZBBj890W2oyvuhmjp+KX8oYNVNFmmyXCbstXL/0vo/C1knZnb
6XFmbH0iqAufqT038NNfVGX0kA78CV8b2tubREC02EnBEqBbfde5NEZSiZxOi0J4+T7iCCftjG6B
+G/KahqjPu1Y4TTn7S0aMeL4YTxIDCNkQox/vig94OJBBfulmadB1cDas/gDgGTZlVje+3+YY+nx
/48ZOyDewdbkoPNoMlwgxQONPbj2wsPAKgyGMd6WYiR/EdHNUaj+gtzsMsimPjv/njvMWarTvfHz
iJY1D52YXKihsn5prdljWYq2Z7k0jP6iLbabbzBQMK4TwpkRzCnZ9GOZTeKnvoZ/eWsuNKqFEJEq
YlUTd9YNZHfBGsqGMHG1vIUGD+bu9egKNlVnS9prnLUItL/vcOFHgOVBQLB171o4HKxKgmoTK2mV
Yio7GHS7hW5Qv/XbHZ67aaQehy9keoc0Rt4cEsvKABp3VKHuNtlBUgnJxBP39jm/PQbCumnmpYsi
0WFk9X+kcBTg60ofLkSrW+1w+MIiSLKUP4PE2ODsyAqfZbaNvhLtpNfsPWJhCmnwoTJNdi7lVREi
qAgoguA2Q/HE9sdQi9PWraqQiI0dmM7BrwAxMn2TcNQ8jwCe/S4punSxtMONneWoQKKOasdpZmUS
wtClI+Me131w+qRwgwVtgAnlo5mBXDvsto87Slh7YS/PdLsgBW8Nrp18AeR4OlnhnoFfqG/s0yXU
Gf0BGhJ5xXBQ9LkS1fh0bWAu9oPfMqHTkFuNO2NTu5tv5jIjdvX2ljCBZD3wbwOancFMupeOsWl/
aVa3IQWhB/N+J3nETFvcw5A5h9uzIfBOssO2Xxju9HuTLkvKvyt3B3vWQ/o6UBfMneiNLQhSWRsg
5NfhbOPgUg1bBGZHnhBfn6tZOlrHy4BXHB9czOqtlVcUUXzsbUXD6sUZaP7yhfgefkSbNK0Hp1UL
s1W7WM316raft7zxFPLn9+urwMybk7uKAk5hTXh/GN8FrHTg84o9geEbUlcpfMv8L9qdtIHPDpXw
9eR9ng+2Q8yUFYk3qqQqIZeVwYt6tIUQFfdWVwozrMcCO3paauNd7UyjkBew/Ui6mkEtJ6AD4TqR
NDUl6pwTXUrQwLmhehWKxt4xcHXgVx7KNYm9GpaH/CORVJVng0idbp3uJGVWEZcBv7LLNKWwlkah
vhts539VoyJt6eRKejMm91FtT3FMcIjAKwOY8wtPy+hgGMWN13Ft2RA84m9a/CkITBmzXwfJaS8G
j69hXI8zE/Swa40fqZjn2KAFnNFtBe5VaV1lWtDeSb4gErPO08IiZ4bUejeHMLcu/LZNa5SuxQDw
lG598ScywjHGIUnwMLoCoZqC0PDHBjI3ovm9EkP9TKqkE0ypqJrv2zCOjqUIJ+f5ao72T1CnryX2
zOsFT/oAQOfl5/rGTZzMf/RFnXcRdi7HSTI1npyBuIsgkvtRJgXKBeB/uFQYHnTRDzgZTLJah/Gs
AyCeJ3lVlFPrh0axlqCJdQ8OIEBy6CCeT4omlK+LNBwYNhssUqtrnavGGAqMK2BmebQJV5tp1L6b
VyAAOyiK0b2wqrqjpyn3vI/yMpfJY47EEE2lK6o0x2mkgmWXA/M0G+tf8pei1XDoPOGd6du/bfjm
iquHPFReilUlhcJB36YH0kp9/YJG7lUgqAAGEIPfMGsRIdRqSqUQ49e4O6kWkQcfuOf5pZhJogVF
0EoqvKxYjMNdmbg2lE/7ERI1Be6yDyt/sBOIiagMkHS9tRhe9a+CknuD57XyyER+hZt/kYmr3NoM
pxvqRuVgP1qL40n339Inu0Y5TxXHan/etKH5xZNn+P6SrtLajwAVt+B8Lu1QIFKOv67CsRS61SFR
8pob1a6OzIoN6/4pmSia3TgXhw4UtsykJzQUQUsirabnU22vNVo/Aq2xNxjUg4ad/VL2CPgy6cZz
IZXjgQyA6SVV8nyI7kM6nDgqNiyZNL7VvO9axH6DgtSEsX19h7cr58U/1NHG66gkGabwPN0e1uFR
PPZfrZFT/cmKcJUIf/jkYfzSFRIovR0clTES9VTElPl7UIgJfi/COBsaR6nrTQvAaPZdd0pDZaLX
mUTQZ1oTm139aDCCMWRjuT3jxXoDcoN/4dw3w98rD8FZwl+GaW7cyOMOMN2KGiFNcvajZXvhDXwh
m9yWCsUcFGPRY/TAyf7KtxT8zH7ePl71CAeJd/YPSO35S769zHhoARLZ3RmHeNCBu6XCiBFuJ2Mb
RMa4Eex3SAGwvuFOncVO+fy8L38JiSx4j3GLZmiwY8DaepLy7tJEFxzlGrihRuBXEancM0aNciB4
CFav6wFjd+l0y2PqT1DdAjbYs9VE3JOQzR1XOnTdHoxgRNBXpdnYxXjpnwiL2Mvq7Huhm/zzbp13
2kcEU7WTuQK6nSgLNCtKkz0TGNolEXs1dfq32IbDaJ5bV1wKYa41yzU+U0c2luOh39kAhzSI1Quq
oeFNSsPkH84mNOO5Q7tucvJ7cT0m9J/aOtJSy6QrV1BKEU+MOutsFQa9138zg/b4q1HKn64I8EF4
3iZcNH+z2YNymOz/u6L/kWM3Mw9zLYKsEE7iz87Lodwzbw5n0OISaexBSUrTWvRVkj5tEYmPXuec
GujQDxzvGffcUXP2QlurAdqMaaqMYSET5SQ3y5mgPU6Yc6Gfyn+epM7oWZukuT3zlvhYbvg18rAy
1/Rz9RCytTJFVR0CwQyhXI5ucpXjcZL4oPdI28CTAot+H0R7lSyg9UwxkMMy2/3lOf95lUzyWxdL
nOHRoE81fwDRT4KFv58PoJ221Cb0mFS80jgbkO+SbOLP0CoWCdm1ue/AK7Fm9Ce5Gn0x6lJsK8kN
jO+gOS7CuHLYJUNwaOuPFpFqIU20d15fqiOnrB5z6JVZ0inDFCpWTnpcxprEblAS2FZ0Rjy+590v
s5cpXRXsc2oaqE96AV+7P/3ZgiszwMBbLP7v3Q7kEUHrECB7rRubOr9OJETFc9rQYfPGnx4gHrAF
q4SWC7LoR7cv0aiJBLoM0S9mdd3DzDF07kEeRrOZqI3ClZn7a3zVuI7rnVnwNm2MUQbWaEWdzfHp
1J/pSLnSIhYHjcxcnE8ZyKpFJQo45oqSf5y3J9UZZakS7+OL4zHnrDvXEaHQ5MbzzHwCNGAs+LXS
EeGbrH2eSwuW+4tAEo519IUIocbi/TyeXko29h+1igX4Ru0jSrFisp05ucfgKZM8tUxpQsw9cjfq
LCpNKhcJTGfWUf5xEjQCggzJ4BxPQJ2zc5opMzg/yhlnaPAwf84qv5TYuz2Z0Y8tPchBY9ykvN90
B2IaJJ/W0PEI2VLogRKMJRBm4plR9IgxIlamlx8CoyBjPLrPm25wZPjQv3drMjyIly+i/U6ageRE
tagrp8knxyn2d6kj9U8SdtIdChjUrDccKO4CYWVLkp4dxwlVBiScP/EBgIsAN0Ls6G2LH0WZXG30
x3C5sehyeuTq4hiZCuHCqVaSXEPCVM/AF5bCZ3N2nsbJzWvpyKjSFSqATdf8MaPvU7VsUMGduaDX
e1bI+y/6VwOtp34WSppaMH4es13FgigB7MzRdo4rQg4S73eUVjL1Vzo5fN/+BDZRx7XeakPCFLSA
5VWfRUdWODGj3tHzm2ZGaR+ikkCWlUz31fRRv3pyT0rbW0ZkncZ2KAxafYAiTyseGzLRTN2++ZyA
Hwn4A8RytP5CHohtzSYTzYU9Nhy7T6oYPvF8VAyAvr54V+Af6CJaiXBN8jD5rXtqjrCZ0NT77QNi
fGAYCMTV76FBV33x6Vpo/322r2VKdRawtTbnKCyZreqVGjOZ32acHUrs24DGo9p3GTfLsnUVoDfs
WgHyeEZOPJ/4k3gMcEJdDSGqfLuLfMG5hXLpVpMsOT5fZWmSbGUgCjx+2mM5nM9alnEzldXxWbV5
iQ7FJVd7cH+Xxp205lfsQyCrki5GmRXbci4/xZPKjJAlUdoqsb8tXZ378n5alkCWFlcwEmkWrY4N
cTCHq7Dt8lOUBht0H5DDX2Oy4xgTW0JDnieubf4CiTs8dlOK49Kps0eMC8wPUn1ADSqDpHFD7wIq
AFloS3wBap/SWmeYmGOC3Ooh0KGDfPGAr+XrTc2NsjwyzIKRIw0woh4tt08jz03GqZH1WlcnGYHJ
PdBTMJjqnJbNtW0FqHA+74SkCbrUNMTvIKZQaHytyEukpnyYmPDxjzawNLx19dnet6yWR2BPpPHu
qi6hyD/b2/AgtYwGWSxJ0SilMyhd5puQYZXYUZY+ORnYLGZYSZJZIq/WMQ3CLlKPVVRnESE0HJX/
dhSVj75AScrtcl9hpxwH2gT2/xF5thmjLGwrZYlIlMIHM+/bb5+WHWwfxeQ0Ht1KxOwklZAUbOEi
u65vh6UGJRluGYGUxqcI1PfqtMw59fCJmLcISow6iTIT+pegoYEulk0zv4Wksx0/yMcxItl6afia
9xpXyh2m6BpMI++ALDDax1IquV7LR6BiAN0icgig+zEiIl0SlBJ3TRPIimmgnxKF+kbnaOyYNVrv
T5//whMyi4wtP86ebQGqK6EKKaDXE6NfAHTsObU/z1/WsdVzZjYIDasED0Gw6c0fvH3yKr3q5tMZ
bJCxLIazkq+rxceEkGmU3xSgRz6cPkq+4SJpODCqJYcFGN5AKQoxOJjXkJKD42hZsddw9LDI86lq
R4XxX8GjY1pr/em2hDssPk5KafLkyisLem/11lON91RvWBmtjA70jkyE0++5/wH+sIVRV5SZZgN8
mzSD2UbPEIe2pBbU4gChDz0NPxzrgJsEh+HYDm/6w/QEdexUBQp00ctEw7MgXa8XQvBLkPx40lAO
wfxtmBhobNWCC2irJEtSowY3KNK73ERlnBCxhSqeEXy+TSFAGHEJBq4iOLkps7GCad4EeQ76SmmE
gdHLyQLFL94QUR3UOz3YgeakSkTtNxKWt6w+QtHUEcrFjMxOICQBhldPSbAIKgLnC8VDgPfqYej+
SQ+RSYXVFOhd6n6u9Fpp+g08DzVXDteHW8wV/uAt/RlukpWG4GfHjr8sFJ26QoizTd7v/yfstanG
CFC3w7/gEB4Tv38U1+CABX7FoCnDTVpddXoCiID/5SqzD+uQemiQ1dpqyyHomw528UcfSj1aYgum
pSl1dU4Tc+UJjCPrp1M0rfMUC25AEb80Z6yLhNYi679zOP49MAoZE5lBS5ikEbMeFeYM0GtLtdA0
NN7ot2QCXKlHZWnOBZWdGI6LOFCNbj83ssGqC798bgoXmTucWfjaatwdi3t7VbQBd7vlUrT11aVB
7iAz+XIE1zRmVV8K9127jqUgj7Qw90oLD4A8TOkFAi9iFm5XhJAmUL5/XxuFA78R+FlgefoAkthJ
9hzoX4zOvfYZmVRp8L5WpRCE0hRTXipnjXnruZ3pDwByz4QTZ6akoH2mvXAONS1kdoiu3sYYnVzr
kljzl82Bxu2g/WFBolQ3YWKcK8rUcY2cJ5OtiGMbJuT7OpKKbFTtShMYoVDvKLDNM9cxaKzNDmM9
H2jy6OoS3RpsXhZVpn/nPeni67EBaGJzDLA+Z8yCOjigrazs3U1Hwb6xc2SwszwYDvshViygBzff
toiPZ/aeb00rDyQIDygGrrS6rOGwbbz6rP6jt9qQUWfHCADaZNpQ0eKoLpwJi1arjkRH0e+/Je3W
lNzryX32lwKMsOaJai16p6uuHSO4CVItox4tQq6TF8oMb9r141jwAoAQG9KNg4F2V1gelWhWFl20
D7Z1GTVQ95tLgYO3bn/q21TkPCE6gBwlu680RLYyACoelhWVIQfwdrVl6tyKTU0t+foRNVGcOYhn
/GqpIQOSi4DQsdravF+YfJFKQb7wgwhCQCcDfuNlyvSJLV6/YC9WFarmwNNUTA+Srsy7MbXSfRUc
s4JE7+JQrQ0QSrOio3PcZWlTfFkB2uEw40Xa7TuIlinYdp3epYoktqhTb7r9qsCTI/oVgU7co3b+
ujqbn15//EtbTXnW7efFPFn1jd1SMU4OaeMda+HRfCxZsLNlmGDV+INpjMjBwPLFIYBsyR9AuUjD
94HE9bbc/FFfKQzCFN/kGry1lNw8eRvX4UeHf+fyhVaUQ7S3FrW+0iY47PfsntqFJ/cZvjaS6NEf
jPoTjZqqRkVUI5BfyjyYMfc++fNbR5dVlUBaD/I6zmNVG3mBEY3534UySFAoEVuRxHHgAt7zL27w
p7vSd3XQcNlFPF5YqUi+RayHBv1RWf7UY+l053lep9YuPCL/r4QuGl8Q8uPvfQq6GMA8ogGYUot4
mRKAWkAWsL5L338rHCsHkWZPEvuIDh9tOzbxNRyTOtDy0VDrieA8txpzYboP6ZLP5XtgMmiT4/bv
9dIZ7oGqDwC6tqqm6BR98jQQTW47jGdsNdBG85cEsdStMcFPEDyfq4rwgw79DhQXLsZtbnbWx7ZL
7ypkAtw3g9UeSv78BI8O/5uSzo2FqFFtX4b2StBmtLerYFcf0uGEKzlPC7a29K7U2ni8uEmjAbEH
6Di4qTq8McLdiVmgBcOebGyQfCLA609Yypgsy1hX/cHv9V8/f9QhHS+6c6PCkF/F3Pi5baGKVm0h
z7MQqj31FwftJ/5eaSLqe3O1qOoRKH4u9o8PWd1N5aW0V1a/6eJ3ZlqnQ+xD1l/6lpyAmB4ngR37
2bFpa5z1UDOaxn56r1CvWvrPwvOkBcKdOY+qZdr5EIu0fl1z6oCz4pkmHfqV7kZppTPdyhlJwxOf
B4YO/sey3QNwrOksNVMtkDR0WOSO3QvqNgqIRyF2MNLNFL+hoT4PM4ovfT9agTGNuqSqAEKgRQRM
y5XmwUlXMfZOXht+g6dIQzaRwMfZDlMutHq0VwJcmnrD8s6zBTAf2rl+AqDh76XkxC2OcYL2qDPV
8W6GdlLpC32s/wDimXhDc+F0qv1wy5W0MxAXC7akxeSVayKdExEln8RttM2iCcojYSjYi1ZErw7q
o0wVIHKXCWNbi5BmrxMnijP5pcSn8EieRvP4q9zfwBESqzYnbu38G0OAYpLJd8ucy33LfuCDfTwC
Jagj0zZ0Yyxu13tFg5YTR1UAap5DQar5yzHYoGWV+atyEZwoLHO5PaFBjKanRPtFMOmPoJqRrcpa
ZdqCpwOb1oCGlF+0lNnmu5+xjsh+MB8D9hh9CgIFrIxOhWFwtMSkGoq72GghUb20MQyOmrP8jOGx
K2KCt/IADI2RwxK0HIPdRYobTC+eo7AsHW8tdyvlwQwczk16GBr3y9Y9UBcrVry2NgJ97b6Nlcga
Ju6wR2/efPJ0pjeoOF2s050fJmmCtMaM7S636P6hy6atFr1Q9/vnbFG/qX3qWqM9QdY7qD7lAHow
9zT+oDu68n3mdK/drPXAsOdjtxbx7awunT3FBVeOZMFdpdLjfN73RgjRW3+bnqUEmYTwaUqt+xvI
oTB1MgnRnJSZNSeM3F5E3WYkMfmpvsHa4uVR2wUmLyRrSdqVF/h0DwbzUYZ0+EC7c5ZJTGO87WCB
Xuj86rMPTfzLd2P5Xh+lF4uPYxsXueE70EaP4+hUDa4F98KgvqzE/AR0FAf12q7wXy/ArZmKccVq
nybRv4X4NaE4eBzgmDkFxFvF3aSR7nKvBLTS+9Q5immNF71AKvK6Yjp5uEs8WtpjFwPMwhNyz8ca
xl3qJuD3ByTImqIkl2n76FKLh/KsnMKOJc1u07O+QVp4wErCmAyYVJQSBQrPt1FH0v97WKrcr2x9
29+coALu6suXMGrBeN+FL4ZIf9PD3Sw+g43HaRwbE9RFkxwhy4sFCdqsVxLkb81sBzsj+WUL1FgB
EyEo8bfjxTMkuv3WOGQpitQFsGGjxlAxp1l1mqZ+F+WFVJ3bFW/nj5+mR9010pw4bbjpKvoLVzis
bkESktCLiK35+aVZNkwqkU0neBONo0LcnDqqEDOW7Z1Y9XR/cVTZUHzDWFAxm4ZhPXGgRopIHA6Y
Bvtuz62+MOb/85krOKRV6utO85gb8JqLFHM8yE0XjnpSdQWYrex5c5f0lvAghDCQHfKQzgFhqkst
cqMDO5D4RAg2tX5sn1FvnSIa1sGKJfFos6sz7O7hkSnxER0Ph2wFtXKrwdhWfK1Kn8iWUv5aad+c
RSURcdKEUB+5gLxRv8TcQEDkqVBScsIeby9uNR5lF7gWM14wltmH62OlC1X3zqSsXpcykcuz364W
8Fu1cTBzGf66N4Y7aFfswrKJ0+xnwe1XU/uyjafeBQPaIhkRSDrNOThQ5hlKaLST1MQZGXeEl5DQ
hV5Xx/eHxumxwVzvK9ikRcYRRFgYERyg6T2ptfUaA50srwF4uugSHwyYhSpZmsQL6ZWBl1k6b1lV
hhwd4dS7NeErNk1atKIJEN16BSIQhJSINGRD12mjtJ7Z5Tkek3rbKX54hFhuKV0tRP/ajBKNeNCD
dGGtD1z9xqtZjVNnTzJ2cO/sOrMre9MrIeMjNmFsPGJOqF9cCoNr7PGOldkqpKr6MCSN54LDvYKp
r1wqeP6VKuxJls7B7ucBPugbsZ551yJCysRpUwBE7fmU6ngYolYDUoWzEMicmbhcRjeXvFlNQ8LW
SOVxefc4oQfL8BzQG06gvATZIN+mqv+jQnM19HDmSyO7ZcM6S9cWsElw8tstr+cquNW0N2ZlF/Vw
bFECQLLTIZXHi5Nt3uQCA2zx9VEoa42HHm1+wvoPK5sDGxkiqviJLGttXowNbS1Nvixt4Vx0wIpO
lvjobkevCS6UgxsbV9/jcIlrd2td4hRZ4FwIvYvF23DPoDso5Gy9MnxandfRD1EXojLDiiaPa8Dt
mX+vAy+hQ3boldzHNEG0McSJo+9Xg9B9jN30eV8I7dX1X3tA0PJa0J2J3Mj0v1x1QOIdhjtF3u9h
K+Le0s2olLF5q1aVTtGeWBvNsAEdumiLDmcSvpxfLuAGTwAby4afjwe3tnYOD00dnwAIPMer168U
9jyM6m3ov3cFgB1tJ0+74EnGxLwrpcINQv2VgHwVc3p5DnCImif3VgZmM8V8BLKqupkhWLXIHDqk
4S9G3ICpV9kCxu0Hp/FUF2ThlQLw1/dM2Whi0N9s1k+Cn+Nlp1o+OLY1Fvldk9IgBBn+n0sFTpxA
sROy/8XEsofH1NdGnKnKQ/BuZFEPGXAQxLzqE3Dt7tjogU+UW6nGsSii1DIAV02i/Rvumu7cbjZF
k/rV3Ui0fFuG7VERXZtnATeJdpTV5yoRuqvPV6OHh5hSuj8gmsZG0Xn1XtHecKp+yIodbCPrNSYk
pQaxKbSNNnb8XTtvx6V3ShfrpifaAu/Z8BAmV9SrLAGPg/yoFbtkUCl7XRVsDzwqpbGgyw6Iyhqj
3WcTK+xSw7ha0FfHcdk4hjDMJB6z1vjlFojk7kCcUKQFzsaaHgQKNdTlXrOowZ1IPZWhuI8MjS/W
wPuYvHLj9a4ATUVi6m0DTltOAy033n+/ZcLU71zFo2KkrYtKKgfyyNezAh7SUD5IG5P40L7FmD+p
JfK7HiEMEmHUchhgfMKfQ6Ck+fipXMye0wVlHUH1xkG8pLJMNw1bVV6YOsFDfKpY/Qjb/tGBp6jj
OVpjdDlUIAn36z6v8pgaIHb1Hp4Vzv2ICUcLUTLXmVtWIa9cmJQW5CUwurKvhpOJCT2AWmwDSeoa
SDu8dQWhegtE76I06B8WJvfXNqYeYBGW7/GIIELhFTyPZbOCa+x83VcV9eHWJMMRIsC1ITOuuP/B
871d4VWB3BjGzksHE6N0iZXMZQXBidPJv3EnA+W56VfXuEDNVAWK3ce2KwNagHRbmSj1xdZuai3c
IlosuNhNs3MW77wVN6des+AzxbCv9qA8NUcQXPQCrJsNOjCic8AqalBfq0cLHwK55Dnx2rP6R21A
8cyYgNlo49QStp6Zvk5Ag/tGyPCyYSbu8twCe6AwYyVm2tv6XBsgv/BRmVhLG6DqV6/DD9VZEi1R
skhqI3Yi5/E036IRe5y1bUKG1drHG5ox1q045K8SuDhTKVkW5sAzZo23kbMAWny4QLbGlNPs9jG9
G0FhulHAqcttlzG10Coj+c5O8iLFPWaxU+2z/e54SU81ughLbj3o02G+5nBJN7Nq5odKqNuxnUpp
mwkmRKldUZNg+bAabTdSexRmu+ZZ8IKLSEanSz2cJi/aMuKOHD1TPALzLq/ErWEIk+wDMpgr4R10
md2x6SB7wEp+KTBU05u8Fh2pqWw025CEdhRfjyU8Griww58/rzRDm9+zWsRpHTH/kUf8FepXuKaj
IF8ZOSAQh5tldiSlDoKU/DqPndynhU42nNPm5MzMJju3j25O7MzPqOW6wfTtqyffhAcOWad5QdNt
d96ASyGK8f0YgeNSLeo0FuEtkPPS5ei6V2W+98+cEk6H5KbK2QHRwx89W+viWrhGwAx5cb9Ly0Q9
r3ImRByRd62Gg9HfIPbAbHCujKZpz+RXfBslkpI0R+mG+OYtg7lOez8TNLwW+3bfCag5XNNyn5xd
ehuiQE2VxSo15NqzlrfF5LaDvvu5F7SkxqkwcNRlaLOXx/UaG8Xbbf23LC3/9yMziKleSHXdvfp1
CTsNg2i1Dr0yNMhLGu7UPsfQTP5g3YFTwHPm2HXWW3OALorZ+LiP3WDlJWRSn8zCBWJ6FCEHthVZ
6GiTIqu6W0gO43SnSXO93n1UpJ9ZMSM26fldbQyTj/ZtQ/KDKbN6SnldnwNaSsTDiOl2ogChU08v
e7P24+5yj41xBkChN/43ALsGkXOVB33cOmke64rteZhclw4GlOm8dCt3tZBvjJgPA4eZf6Q59w5K
Xkp4pkzbwIN2M2bj1wnHIYwG78qMM2TeA7UTOC7FfCNQ4zhat7fl/r2OuStC3Ref2et5yKGty0Xr
5hiAAl0+SpBeUs0ByoaNQCJG/Azhan5xjdeEA7b8+Reu9jJHtQpRu4HXepJAy/w31ln0NMiX62lZ
xHVab/B0hadBcCo+kH702A2S7MuBgPMDnDWCfGXiThQksbKNrOsMXz8m5jHPfbLIreRSkuo4/CbP
ra+zDrz+YfncF5h06mXDUN7m39t0D9KQnYFxMrNR79TgFH6gE/LLcUWvo89r6FcXIpItV8Sl23QP
4854Ga7SG1sB/tGt3N3VuBznQhs1zcTUL0HOAe4tJAESxn11RU8DtwFtqo1Bq2k1Jd3Zs6GbDILD
6fB4KdoIDLTiag6+KGIwwsbgL6jOhWNwH2HhthfVufwvEPPXmfXpIwIOKGNmftMfuuisQbg/bT9L
h7rJt2WwFI2anjnhFWYFnq+DJM72LjkPCByT2z1lSO2FmNICevIZdKWejeAJeGJY+TTqcDwljl6M
sX47xTuPAnIFfWR83oDpqTKAOaZi4QyM2hSydxT3BRdaMulQsUct5G6TQWK328vWQFkmi/ZphzTm
qpLmyD/21h2bTGk0NzVRrzEA/Kjo15APgGl/MQLrxlX0/gnZ91NQ9TRFFzp8F+ijTx3pu61WMxx5
kh5QIoVXvrT+Va2nO4ZvR8u5Ay7u71K9OQN6IMZ8UU2ztEoIl+WTGejYd3snhelnop/jCdohhGDe
air/weTNHbNosYimmdvGXopOeqBl/Miujt5T0JltpGMZm19UdM2ckRGusYPUg1ruuZOhGRgpdMhl
Hu/yrCi3T8X0eZsI8PtyYAJji9OxOwC4StY2JJA1faO6oatuoHeWJO2pzROrSteNpgOUk2cQTvJt
dp4KYjoK2CM4fpuXIocAAX/noPrRJH7Wsyxl6LhXVEYClsgDU63e+2PD3YkvlTpefsU9QfB/zHeM
4EHT5gcOAquzkEBI1Va3tkMsmcw68FtKmpgWCJr5h0lM0cv16hOrNFUJi6Tg7d9961omoZv9Qn9T
cg9xnqv0kA/h0QMKrwfuDsmc7VwTXP2ldDmk5/1SZ8uWB42y3x1SV81iAFoRttykFU2D5tzLZPiW
l1cQ4H90WK/xz15AhPtbY9H7q3I6iF4S5E+8LBs/t1SxIlvbuBd6W011302NHFlxE7w+hDA0rZDK
4iVIyHYY3wmDsKZyJFschEn9CR5sGVKZrJBSaiHr3HuKsFAua0Xy9UqpQkSUILW5JT9aR3upKyku
n+e5xSchvXSoiPlF8rGVfOEE9LYkvohfQpkGWSCv23McKhitbIG/XoApYw1RuIX1dI5FUZefn26N
uHqOpeyyNamIsj16y+5mFzSCttyCRJRS/+1nMwuiGw791MQRmi19HBru6d6Ytryyy5jqVcA9E2bC
0yHe7Rh+BlNDs0JBhltrR94kjNCbrRhA1mIQClvwQa6B6g/Omu4a8EF3NdYjTnz7PyG8fP2QenUO
kqa2cyqzHXA0/JhA7nsrqs6cbHxDSRU96zGmgZYde+gk/hOKWKruh+lZMz1o3vLsgm+T++dmYLeU
7/RvKG6y5H/1sPM2WHIwauVBI6GXYAz+mIdMQ/L5H2ZluM6Rsk70xeXvFCcmBh1/SDSFN1begHC6
8aUJQm/EwHf3Pctnwyo5yCeE+JSNa9rzhs0vsEbexuuUWNb3IOdrcTlxHwGyj7zCKsvNY+izhJTS
bz8vTwB9zUC4bylNT/r9mHab9d8ot/Uhy0awpWHKRtXI+WaGsgdSk6De8T49s3oXq5LCEeB0/ZDp
SB1Jsc0Rm+lmWfSZZv8QDJN5JVJC4IvJj1KDHkitYZ6R//Sk3AkJx/f6V0tjJWaO4ZQcn19vPb5B
EkSwlM16Ir0ghp80TJNQLcBJRgIhI1OOFmJzZAdOZkJ5uYoFR8adOGUw/s0NGBZq+MGg35rgwPyH
HqAvqV/4B36oD0+6iDEUidl52pwJiWlKRoKIAWaudCBA/ChJX3ACL378cNz1HEdudGbbkV1u6XMM
OAqMzyCsuc0+cx4+vHubqw+CSLQBgnOJnYBt9hdaQ7fMaVuJqfViOdz9SFSZW/bvPYEbngNtON8X
CaozQsgcKuqiVtwazhNjm0GltHoNDqs4q2EeclK9oM4KiOWsBEPp9V8G+2qO3Cu0LgLYqQwMze9B
bl9MZ6FPBxRfKVuCKm7HNavXggBq/csG2/jeWuwLvR+IVzXNNMIsr4k5dnU6oNshHADB7hp01ufv
/fKHabHlMR20LnkLWdib2LzqlUModl6h0Sq6TAtpetBb/5NAOKY+NMs9WyoiowFGKZiGWU0y26Ry
0vOpVeHR06x+SW4EbgG3x1EatrqFfxi9+Ff6gU+JgFX+h35NGqUWVePLOQteZfoLx5mVQ6pZW7n0
gtZRrK410HF4waldx4wS08MvSSJ2NDX6iiMZ4R5/j5+Ofz1DBNgAxxEflBcU8ck5Iy4HtCj5uT0H
GNTJIxaJMJq+A/KZWEyTJuZ1SuDxvw4dFBvlGJrHwlwAQDT512vJLU7z+70pt+P1C42glusBrDX0
ZrxFbD9ixjbZUB7bXvW4Lszzl0glkJ5vkoa6p2szMa2q9zAVKybjS0GchFY/KBQWuDJvDQSVQ0Ey
2qBygAhKL0qHKc4f+uEMQiqNlvryQCnK/AVot7LDK/2p2boGVutoOc+HFHX4EJMePyHau+IFfw7o
zd1WlFVGjr5xgZ+m0X884OUdZIHr5PEyB80C9uXFc8Bv7x/VXCeg6FGbIikaezBD1OIPYtDqOQUK
6EmKJpPWUilpW2OHYE1ZrJ/FlbYHKMko5dR3NtF52YkZ9s42MRwQcAYRTLHk1nNDmZfq99eqq0Rq
IKk6UJAFcMNvzk27wzlbrCZ1J1zJqyKb9Ma9/xmq+KU6j+FDJkRl669C8ASnIAk/1pQzSv+5b8Y5
hS4jJN4pwzShuXX6GrNl8w9DnBQJuZIjKMok7AdphVY+BQVXqgqEY4z4/Ql1at3JzNB1RqjNlaCJ
RlQQZfiiEpWzCa74/qY/snsXf9eLozg9HdH8yJ8EwEdWO5RoKjsaBaD0TZiNiDVKmM3XfplvanjG
Oaqdt0JPFKomzSJ/EGGHVmEEcunlYLPlOyGTZNFKtlz8Y7tiCoi9Fg37HWMBelVXCTWirjC5EbPA
8+uczeAtPjYBPkIN+5MbVgdxHC7V9qMqDL3WolBMFlnCe3kKyXqSWnO3jXkdjGoE59gKxtAbBDby
Lxt8qyVDMgfvhzokzcfaO2cLkPbw8Slf8Tev3JjW2bW+MFBlaCkRK+jutQOowxRO502YTP+H7Kfh
Jj0jBUca+woJsx9TMkapVixDx1dHmKZqWWDtqeIioIWENVGTEEhIjAoSkV+dQPvya7E1NibwHo1J
llHJRQn+mVzPsDXKL6h2TZUwnx+78PdkWCpJ2DjNYfUc0Pc/ScGHFZS1YFKD8NKi1GNF4lOQC7R6
OvPHMo93YjQh/7tn/4+/QgUJcOqmpsxlU/cPYmFrO8RNRKF7qnrXyXycjQi8NuoP6SuM6ORfvgEY
S9wzDuXDV1qdfwSyN202IFuHQsuHCmWoEi5yV5WCgo8tcFHy1alD3nDyIeJSAIV2zJjNcymRqmn9
C1BIrfTdCfHduppugoqMy7noarZQ2DhHD1SsCSjkQ7SXBSg0vffuAWI8qrJC2zsi7U+BPiXfac6A
hAezDjn34TNiZ3+yCmkRnXMBxh90fBEKiKtKsZITg+F/cazb+OwLdf+sawBppAfdxCHkz6at2wOH
yGEKeHmsJFYhA1jNBWzP2bURhPBcy2E8K1x/UzqmAHwxiOK9Mh3qFTYU5B2Tm/563eowsWd0QU28
HSp+ZWvt2sbYf3JcvihOdVSyXHJEmygLOvg0ClK8YJcXb/Av9F1RjKjq18gso6XrdHHZo5q8RuMq
tfoh1qw4KnclniwVbzFTHh4DuwZHYsYcpBoAclOxO1am4hoYlpFb4Y+rmXx46aWu7BgsuCGgvXnD
3V2gAQVWBvMmFYQfwmF2fwCGxjzaB0x47zWrPe+JLzPPPl/h/kCj2x1/tSl1//tmnEJWAgE30fuj
BSqx34q54wvbMwNXWeJUOz1RXvhvc2Pt2LYrltml7J9avbqLyiieZgPT62TyVqM8flHijqOIGdh2
spbG5ZTHyNiFmkAjjaQNZYfwRoHn7WdQaO1jmGKx44nDnBHrXL3xyNP3FCPgr9k5KLjrKmVj50ij
5po23/pbvPIZH9AaHHq7hRorRPIyHP5iyynMT3o7/RAT4PqZdRoizj3BWUMcN4+TrlCId4l+UdE5
zpijul2YFMhgpIdGJIyb2xsEsiOfr48DWTTZHQxOlV4XxjK6kPkSRRUxQ9e/LV7o6rnI+Sdixczq
HGLWdojLOcmW+2UqZVlHoju7Nw8Y3c+i3ov4+xQ6QILPs4cdntPRI528IKalaK3AWUI5MD1Abj2B
YwtpNwSvt5tdNjmQSOhi17qD4Zx9c0ScHh/vFGoViaBQZE2DDrWDJP2ETWBBw6i1qEMkQGXZJiwg
6L12jP3B633NVDvkjbVdSZd+HGYUwt/+MWjv8ZmBg+8G7aJrttJLIfjo/FpxgM29QGt+1EkRpZwA
brBEEETLBes2H0jLKB+plVyCGRe1MDYrVlZtGCKOmf2DeJ8nKPKQcI/YsPr6ceiPe+NaQquqWbGv
kzAy2G8+Hnzj11+0O80o+8lXdJwZQCMoWX41epx/aABFWlAb8MX/yc5Mj2hfLFYRhdH+jJuga76K
16+Zh6/DK7cE41ILubRjIW7TcsUYlOozB86/uOfy56VUcFpuWgA5ACUrT8jaisNEi9NhTbi73c2Z
SyplQqUeJv+IfOUeMTxXWks89dVE2WAgp4nbyuneo/ppufWkwq9UnF6TQ6nc+XTLDWgFDC7DEnON
O1XlE9Yrwb5azsuBdUSX3y6iwTjy1KOGw6gWgyruYGqIHfOKuen8tMQeCzipgz3i00z2QSFnsRtx
agj3mijfUukif8j0286JLPd52qDdA2DDJaByMsioO/WaqGZeOaOjt7v90AF8/uwUvI1gMdTNyKhl
h8dGU9wWOLaEMoGC1jW4Fi0ljSRZ1KMX+J8QpPzxOPZ/B40eEgSOnAlnMvUP9ziRNA5ZDR+qgaIg
MWRPnnY2jbbbvcoApTP2gz7Y+TBhzlwNf8Wo34DkqaS0cPzk/XD4OmiSsOfpjhk/cz8DTIS4R6+R
Wfj4J/47oDpVSDuNZ7cJGJ3d65Vhq3tR3hEauRRVgj48stYqifgkBZYP5Ws2+kJXZVfkFZppwuGp
+YDeKW5nFCGsQgroBKQ1mcyYvMJs9SfynAs3kAxnEQiTKm4GvnpNLy1eLDxmgVxJqc8qXL/j+JQn
xyHo+5wFbL8hz5wVBFaLcfPJMsWXKS2PQGXe6XBUvn/Or6NY0OmUMYeRINIM+hN7TIsvaBQXCw9s
RGeS6gp+xiEIZWr5EJEI8vJDMh6KwF+UeVeFcCBls2BF9qXXQ/f7AdmBV4vsMVtUnaNXbImlWYXv
+PNIBdTR+RSgAwQZWDPGNnIULnZu855RJEbrG4AhVrvkFUtAaJslXDzEJBE7xHjzeOhgLl+zMxbd
MT6ebzsZHeu4fTjw06AODk5lq2zNP8tgdCegv8a9bN1aVIXwBLyCvNU3DaacKJDGk2WHuVUlUga0
Pb3JLhTVPiVQYvmBVv1ryb3sgQwcalZXklukWNlheba8e0+PQ4uB+u942RYD20KFTkwNSRDZGDzT
9piTdm10msR7vympzNGLCtR0+34iYcZ14TGe5IQ8Zq2CVFcTmu0nWXQtrCWBYF7LRB46D7u12m7p
bCzHi56nYk9bLSc1DB+YLlxhwRNAeF6MS/Iuu2Ll/nhR1iCLd776hP1u6hDUTJL9gPTql0tEnSWq
1+FqtZSmjIq+9XLC8gb20u3ECk2hPVkuZHjeTggkTHbUr3+Xex0B2loxTu2tkNMMmTdpv4Ud96Bd
2TeF5aIf2wiz7J9AeRAyVKZbyqGoD0JM7Y0TKSeqkuEj6Yki4oz6otoY/fhl7u6th64tBjrS0H9F
NeVX1T8yuCoW5Bxf+QbHahWwSrrV6PFyJmJKHBkGP3H3j5Oc4BwP9j5g/M2w8Gi9VPbsPVDB9nOz
fbBlukhVw/ub3zukvmBK8M/EQ75KsLcDRyD7wkQQy8Niyz+brEfECZxhgFanCAglbhXXTEvySQSo
T2W7SOIATM4sVazXkL+7a7orlQrBAIa1zt3QzlY+UgjIj0KWDP+1M7lRRm8B3dgG4CAWgBi5HmyP
FmaxcSt/f3qP9bf7x0CjdCO2tt24t7UVs9Zua5OrV/ppFapv7KnAiTwtkdSiFHFOGEYqpkebtf5E
4K1lTzUZTgd60WnvD4DWs8uvM4wOWoEaQb01+FMkf5ukIaHQIg88AlTW9EVeRgCrklS0uJtfixwe
YAjV1tJ+ZQDngRTZYIbtibVk48Iq+DPrDOxZ5GQnea/WCge5GcRi6jypz5maX45cmb0T2YJ2izBa
JVvmVwTvINIh4Z8M9g7fA/UGdEWHklM3TVyEgctSlUga1eGdGXPSa9Z2NbSL1qsQ6TvLrBUNhglb
tXDsrThZLFX/4Up14F0IQ9e9oGh4glx2SbXjiwbjrJnvd2LgJNh467gN5dKm6IzS1A6VFV39+tAG
JbmTDVOvkhh08h0hHcx0zGO/8kJemmgOSRo3Uxzi+t3HebyDBPgWqd+O4lMD48aYGJgmUGAg9goe
xeoc8AXpau/lulGmNVNK1eeezl7KaVQPwf9APUXpxiQ64odBeOyE6TySzvO11nBnhIXvWR2rnvHI
DPnZeDfiDo6Jcjx3iStyXQKyieaiXCCpKlhvxNXJqj/NKeKxmgFxhUlqPwE1+agzGjo/+/d++JKd
3/U67ZNKUX9BVgMOYoOC/FTRXxaonWaLl5hGIZDM8sUmO7Kq6MZjSVry+iysZ/u5m2/eBl5UndIS
87dAyoMdjwysn5rUz+EC2tPj/O28fpOm8jIyosFbBaqMhkEZ3+pLTMrEWYnk7Xr70Ke/kd5EhYC7
KKt3kTBsRXncFK0PmlOaPG17DQPlAfo74WWVuNITxRBCHJKSXx6/M7FB1VtImBgBwOwqwifWGiOJ
fKNVFftVFgnltSHS3YGBEkBT0Dc9yb6+k4YuVlIAIMOkLbNKpomDnsDwbkGU6/JiRTQw1NvlVZ5o
+mZvCww2+LUP8kWfL9YMjXPnVQeBoV209cDgmGkTWKvUvfuCOQBtzzfx/R9lWRYfQC9/ON5MV1HU
1qI/uNHlAfX3dWpg0f9k8bgui+IWab6+G6KojLUyQZ/Q4UUeKiYmZJpV8ePoLp7niK2YfzvMTR0b
rYnhqHIcuUWVUR7Q+jvUDLLFuCukh9epvnixD9maAweMBWXmD3TEJRd6uBgddeqkBUDsmykz5snf
7eK0JnPXJKoeLgn29B6za67AHEOH+glvuwAx+ooRCi+MAi2MzlPANyLzdi56m8dm/yo8h3tAPADa
SJoQNYEwEsOacqst1XNBf6m2QgmdPJ+cP6g0+F/aokz1TBPm7Ge52Z+774A6LVJhSFqycB6ahnkR
ixyJEJClyYVbSYZsgqZCZWLAW2dwuZUf40MRa80y0WDH1j3JOA5VWo+Nx23p/8FezyZ04zUbfRd4
n6YUCCEauHY3+c+inTKuOJ5nY4p94Md+FfMiH0l5seSIvyfZiq7KFMj+5z9FNNuZHSpqMgnZq93c
XFZ+qs6UE4IGPhMm0TULFtX6dlfZveL8EVR9oA4/KqUMxLB/x37M4HvQ++Ev7P+bo8fr2dEUzrs5
1/65eO6xGzZ3uBU6/IbekarLYrD4Us5vvxakTUFxtir1jGg9rrMXM8eBnBHXirvt/D5NlTr+cwbV
AL6QIBJnLDR2LSTFPzxw2ut5ZZN2C+LvgVL6zgQWE+YCCpPypknvlBNFaj2C8E9DoAL8XzXbsA7s
yRSBSFCASE+44v7o/C/2sX0CmJnExpy5xa6CKAfFKllC7+cIWRXaZM80xJ3RM/iYpu5xsyqQ9hMq
FKBdm0nLEaTEYr0fK1yICjew4FbGlyyRsV9QoL59uQ5fqbgFIAPwyFycuc6Jk92/iN86+KM6bfru
+HmHY6ftDmPvmcDLYujH/B+CWynJWHm7Ml9gXTLFeB3yqfmBFzyu9ZxDvUPGLW5R+kGC9PLWjpE8
fNvCIehiUgqcc94acgXkN2fi9g+gq4VgzgRpQnOLQRIXHLyJeApQWTxAn0oxTrfmhV0r0PUL5akn
rSnKTlyb1RzsE20r+UQ1IlbGdrV85A7JZ3d/GU3oYge0qsnl09cBkeCshnCXDARl/FLhzGPuxFku
Vs/InvjpcyKxv9DMYdX1N3Yb0CGylmri5tQ0aBOfSgC9KKUqv8JEu1xUe6so8JlPXFq9ZKvRduer
HAqBeRB45geT9AO4m2/SPnxwEQm2ne7+26VPzNTBTxN8A28gYTe8TIT90sjzgzJwyY14r3yP0pqz
6X8tgUvqxK8191pxgGCsMA4AsfhL9R2dVge3rh0DPezac7mRJ0WHlM9UBGlMheYfh0vFEgAiRapM
/WZFLFEK2wv88OJtkWio525+PR/KMxIm9FC1TKb3fhrxz3+SWIv8lHg1/0IOMJAA3Hv7o3mYtQ6l
hBOoMksl813pb8ARc1jRPDmXdcDi0g6L8w/M/aWf0VCbymzg8AdFh1mjh0CuBVShfGl/Zi0Ha1fP
56xHNYRWxHOcQo0Qhf82sZTi2nifR09y0h+qzMnmJthAJiQPThhFiiA4ge8Pzhg/dTHcyhkmwNRr
QIAkjgSC4QaEKLOUY78gbEWCG4+JDG8nvIkxy6nNnHvW7ZUE/wTNHnAIV8IQVDRpr2anZx1UoAum
9iZrpLVm0H89USgjY8JTKpoQfaUCQVAgndKlSybFEaHawkmBmGepzxNgRewES+5xecGX3mXO+swF
+IOTWiHu0xE/p1qTVN6G38oAaBilCkJuAEBJRpaxlSWC7e/NqUAKRHx3+ht4X/n960Axg0FK5nGj
7nE/v4+HMIWUFSFEm7xKbIKD2YIP2bWoDu08YcROvcmcYewqihityMvrfXLwn1eVh405xuqZKh/E
i2Ac2lrUW0URaCpRe8jMtjKlEzBUXNmnEqq2bC0Qh7fbSUmoMg2sC3bDT+Qe44Jzgqd6W5mk+O50
mouNjF3fAVCHKS+qX5HaJanWhLYrCUWs0FouBpqWIT4NYH+Q58F73eQWIOUsOAseiO+YN0QoFUWk
l5vriItTCpiHCraK3DJbrkd1xUaMbIH+U5muuc0qmUlCPOt6d3hCCKE2MTaE+BekrBzv7CHrOARE
BHCKnrmh9A6j/4PAsDmJVphkvgVuGPyxEGbr3FK/1Mxbocec65Xd12+Ybn0i2zHm0JtoNDxOx4z2
2FSk+YSP7Z6Vz+l6jPM88pgz0hKeUYcaUeAKuRAJCt7Fjcibb+ERDtNPR9n/lnlvSclpuu5COSXf
6maNYYrvkTwDy+cnXAg3FD66eFqyXGqwp7KRmi0ZQuOLJmLoBrF+uI4BLvRrV/no14eFBvls7BJQ
fKTevM7z1XzHD3p7fms3ZTyf1s+Rolas1l6mbp1JB5huHCiNOwfJ/VGa/pGd+9Bt8leYvo+6AElG
xyauiJFfYFCNJ17ZqgC3dJXbNRNLyPPyhvNnztsDZGe2cDrqdzbdCXPJIBuIJZPATx+wYwd9ZLYa
WZ7s3n+GNPZW4AmQRKNd9P0cAszOwyoHOt1Jq2WMYfhkYbUcWaqFp2ZiDtTZJ25qC4UqMC35c7XJ
lLJkpxroolhSorTwdyvcfbgJx+Huf75ByHFl7xeqTBq1L1D8cCHRquEUeCKzXj/3rYV49mqoovfX
EOowTEGgxxzQCbodR636kjd3LqFuiMIvPoxFPDuJjdNQQAhFzgRi/Pd9ptj2Sy3Q910IcvL3+DoP
yXm4bNGG0iprjTOR9NiD6gTwDim4akUDrzqJWzZVOl2EZB4Q00rAyPCCJ8+/6+lpkEmRPXubeAhD
WnxAqBuEhX5c4gPJV3KYBqKoJjSlhxh/xYQyYFeeaDqa+12AJyH2gDtAMw+lm1158W8b0FXUo7Xd
7z81vnbhOVd5CR7NOminViYLgLvJm6s1X1fpaooyZCxUCDqjtvDJ8lLL0aAy0iLeQ4+iZTgM8N5i
6y4jO4ZJRwwvDZ7V2PpmV9zB4Q5RQ8tEoV0fsbqEqpPa24x9Qn/Dk7d4bWZJ2Kr3wVO2mwC9X1ku
YPz8nLqeUNFCu+D96GTLqGaknxZbQfI/LRfeKzsKgk671jwkVRgTu1kA6HzmS9wD3PGvQKFATEcj
VNmX/f4G41DdZd9aLAs3B1Zncch+DJslySe/JmJDouViY4HhJKxccU7ozLlcyHxyV6Dx0/YtI0LU
LKLHj7xr6YHMq2t/SC6sqvH2EmsFl/L7LEX0yZgY6hGmFNHqrdec+qIwiLp6DHhjbN4+DUrjTwbB
c8mdujKLkeJk0FRVrXM4u2bxyY0lZf3D0qRDVTCUu5ZDM1eeTIezQOm2BGPIExVhgclymo9+1D4x
fuLUgKmjRTTet/Kp8BZtCk6KojsXJCnRJNUO9FH0JUQ8Lnw7pndt2aRiho98nbJhoO0QnKfmmTsy
NtX1Zb4HQ+3tvoSSAxOZeaRJ2WfwIisVm4Zds9up5biQeiLKI36Z57pceZkzzHxIncsAoYbZj6WA
nMhtb/e/B0K2peGGE13EBpe75FVpqzTzXOcrJ/NcUagqtAjvCijlToJBVsNWnowBlFzAp+FA9Rk3
E6Qtz/qSSVmWtQtms4P8lEYAy3edF5Livk9uTHyUEsD7L01pfcLB+8bTjQo/R+tzlwtSGynpbPFM
4p4my6Ljlske22y5ttAJYWiJntJvqAX5Fdh1BARDGtJcQ5mEGAIkbzCU6i7xURETtjgclN87uRCw
JZYoUZbhvfA27smInLDwl+057o2wpClUT3HSi2rLZDQMy8l3gHFaVO1NvaA1zyM5eTpGg9vSSBoW
JfMgY4kEopurhZT9HVorQsLPq4hfHC+WuFt3KJEesOQ8+SOHw8b4QR85CNGhdA8SgxG5GjcQzx82
2BFZFitGEX7nvVfFEWuDVyk8t9HlLrjK1ikFYVHCQiRA5S9aYZjwxG5xKvGCPgfZxJY6xFv0Jn2J
Ton24K3OWro2BwhtQB7ZPD6EtbZQ5B2rBFxZQaHnWW50A9SX6EkV8/YgiX1vOo3yOdmNVaSnRIy7
RI1GdnaVk1x6iVEXLkLFCwpvgr/Y4nQJwIYrG/ttRaMc6vDx7u+jQDFnMvsMcTisz50ox7imIcH2
CwuhuC/NqEN1kbMx4eWj4hzx+mhyZcxFm0870InnDpaN8oJHOFFeJHw3lK+NQnmvfMFLiu1MpJ8+
LEHm1IAo1IKOJp6uw0oH2G/q1wOMXn40tveleq70SPK5YDwgL+bKThlw5gb/gN0RX3NACy8fNjMl
4uiNzIPI1bLYjQ4gQ2eDpolTHNTIMFCQAu9b0wme/NkNUbb85sMUhLcBxGu5kgDyRuX+EN8b9aPq
PMdlEsHUlYAk8AupKvXi5bP2isJji2QWnLmmu7QAb8rIoM14Aa1eCvXXzZJ8H+2JmcZ+MMHiGMvc
KfMqr7lrVpuS6XxfYm6dmCtOlC2pF2uiDR/QfZJTxaIS9agLMbeCjz6MnJ3AOrlU58k3cb2PTHYr
TNDnhMM2yeQ8f7qSkbKAAR5MZiftN2FEkU2viL+itAVQhVvvd3C94R57LU5p10+xJQoY7Yn1BvIV
34GtlsUqUruX7WvJgZg2vpmZkYe8qTt4E/4EeyfM4MHvAHJw2P+TiwjvnlW935e6FA/tArIQWBvV
0Bi1KZ0KW0PbARGWMTpw+7syJ/wJSRppJX06W8EyhNnT8CaZt0Ve81vF8NQVE26If5KwlVSiRs6J
SfytsbEGRIi/1BLgpzIE+vhaLR4HArupQASiu64+c/BA3BrW7K7mgzuc/bi8UzMHyOpmsBlsrPEm
udbh62aXgErwH+NdL5KmsmZte7zOmrycxeS4QsNPMg6gjtdhBAnACmbyOWukSuliApUQhgH6bvxc
yD4BZc6BSX32Q8UwMedKMux3m7EGFNADCbRqk1ZaLGbDeOa1RhQ8ACw7yD5mx8sD+Si0EwYfh9aT
Sle+vlmTVcEvpaw+QLClE1KZwAKKIQ0jz3PXcfilrysVrLEH1Mxwv8hNR2eluJPIB5DUkIIMVf2u
lhS7DILK+n7+x2CzAZx2hPjO2RONonzKkgxW2DS8q8R0cyahpP8w/ZdAAKmTRjOV/2A0+hIcMXC2
MKLQjs1dPoCEKZXIjs8P+tV29hBAQkYRgYh5spnnZVohKLwT2h3NOPE+Y4AquyMv0PEFWSODQhtE
jphOTbb9uXUQuw9qMEnDmvXe9W8dxtPea9PfV1uB8sXoguJ0nAqK5WuRhp3Cdu7OCp9QQmxQtmcg
nMWGvMwbLTPvHrOIaEQBF1O80TGdrTEoW6A6XBfrc8GLNno941iLadRn89cXqnquJOG8vGX6pneT
cy8+wMN0Lk/kA+kUQLhGss5Ge4i0KI6uhcs/Tad0lkSJtW39D34m2HY0ryFyY2s5a1j5rgr19a7L
8q8hSsKXJKt7TGUC5wJ31Ll34icN2CMpA2JZb6G9+6ulmncl8KLhzZuM10g/m5FGN9zrJih7p4ks
xzEJui4A9aEOu3EDpEuKYpw2Z4b5xlq1QDGomnhskKgnTXwwGhrS0IBwp/bY79po/w4KS+GeF2FM
9Pr4bISNn/34ckhQZT6NM7VF27J8FcfrHF680HuI/EeyiVN/a5uT/eK/FbgKQE8P5xesGhh5dif/
4Ya5x/ZgJUhGwKHAKtfC5lK/eStzAqTD00Q05Ok/Ek3g8N1HcprxLpbnK0mETAImj2lfm/tiSm7j
CnJoW22qV3T5jRoEvGq+2qL5voTOBXZvT9MOQ7Ypy8h1zsBAfUu4IbvYoYr7BYH55CbPc1tQC2nu
5Y4HkV4vl2g8U9qj3rvnYw3L5/ZxRG82l7rVmNz74iI77Ui+02x0JJI1mT3D6aEKuGweOmTU49xq
Z/3DGIw6Bq4kp2KJ41A/KkPnw80eSPMQuqHTZJ9GUdQ2RD46ypP7XP5IEcuQSbiXnx6a3MbEg87a
nc3u+OiCZvceKzSkPj9GcYAWWOIddCTshfp8LvnWEPwknH+hk7r2TBgPqU9AiIrXUYpRuS3IvmYq
/AtdhLbk12WzM19WhprprVNcHEU6rJ3OWMpMIsj+O8rN44RTzaeXgdKaeUT9yf1bu5dZ87nwX4tJ
OrOVKJB6rK3g/7+mKdP6piacxocMFSlzYPNaZCeJsS/rEVoM/xRarrNJ2/K2kZyDGq8lKzn9fllB
JFqIGXLghnLXym0zDTeDAUwm4NAZT5TcN+Tm1xDcO00hww9+BLvT+DHlkqW/WL1CaeBNkJgFhNDI
XUDsgpBtj7uaX8BAzU/ZpiFz/x8b9gfxcR0t5bQ14wq0/itAxhqezr8Hezr0uquuJuK2jO1/AOaF
N2f2LOZclil8VEqyDucg2JIMyXFoZ3ExYNqjrFw9sXmEGmlwd/X2+bwY8GPnIqIOgTOTi+qNaG8i
sRoL+b9Jwi/xHwBrHCKH24e50PxLdUk3XDJbkZ9YLjpnbiYoRsPmq7BZZvtsTPWeeJuhcKmi2KvR
CiBfiQ58ollwtaDJA7YE5KcQgAwWaaAPz4uIgr5ki4GmTgIjeZNNiz2LHoFn+HG3DIvYY0BIiwjd
w4ml7AK08phjvWqoVUWHP/UzGtKGyUTn9YPo01L8bd5jGNwB7OBOrosPM4cvPdBlD0QBOrzyTVG6
79+999N+K5l6BN4yqOxou8XU2spy/Lcs8ocKoF6MWwpObei9C2S/wFhFkQiLGhIDhUVYSm+rcKIu
BkS0BC+oINfETOYevEcptPlOa2mT69go6b779w11E8Vg8vFjwwHYBKK+yHRvTXZuvSuPgqXwU2Wa
J9ECehc/CXC2wRsYk+koHY8onEww4OC4iGOiERuNjWfKNBQ7oeaTtUXX4oOeYQGhi3bz5+V74GdD
W3iH/zQmuGsXWjAcZVBUxePMKwBdwOxySmeLODeHbiwt6TAKmukE6XUgwG3hJrIxnHvGrbDgwZa2
fXOyMUfy38Wy8VU+CVUypzZA2yfwBS8eOLCoim9yqJ1gxzBFXN2SVUvgk91vtmPXiAP1FOWEC/2N
tWMSgWu6FlTAJ3WZLLb7rbrELrJumdCXlLua/Vr0eb6d32q9Dv8Ir21KRqWbn1DhXYCj3HUNwAhM
J5bsZZJ9eHBWjXgSyxeHR0yUqNkfpDj0zIjgtlTLoH62MxmP9fowYrJ+xtl5RPJ933L8QoFa0860
q/UiVBu6QBcQKalHABchR33E/JGGQCTzJriCM6m/P+a0+9BLjLINy4/MSY9ufvoEPLZypf00BLOr
heFfaV9S47/Kkp71DyY27tvCbQgGR8F22Zb3WVaPV4nfwGT+acSRkHzKg1ofQctgIrkWTGBTAG3b
eT0skxkFoOShN7B+6bmXFFs0bcDowJU36XWFcw0e9GVwdq6bWphPaJV8gGAPqh4t0T2AqNnT221f
J5t6wsWtzIDGgpgcX1pfQPha4MSrjmcuEYCcdq52ugl6JcALvQPtwl3x95wChQpBr7eIg+hzfROW
RUDd+XLpDu47UmsgYlCxdWJWpZ66LjblVDtCgGlX2tDi2Upj991f79KeU1RsJDTy9OIkysQboZyM
m/Mn0Ejlalv3FJ8DswvDUrfWD+lYip6/1huT8YsxLNI/JLwironHljvQImPbZea7BOuQKg05qrRn
0Y9J0KE8HX1lN+Z+NcaztzlJ/XdFL8yLvuyB3cO64l1+8zKiyx/7dhQSwqBzPKgAAApKTA3/Z2a6
RwGnNZkZ3tT19y3peERmCpp6MY44MZn1h/6Ut867s7eWAbUQOZCBRYgbu8Q/9KHAT/1fqupVT2dn
fLkF2EiDrfny7bEdV5AE4yAShCd+YXdRyswuukA+qjbyFCmmVho4rQskWZTJP2lUO4xKmdlo91qa
0ngITB3MinJRaYQc64JG1c4d+1iMtzysBhZ3ZIC0UNVQJcBsxWkkKUc93xYuCULs2+37xupJvuMX
mpg9n0LmbkxZ6DMvp8ehyEawfHdODxnCS9X9FUsD6jstUV00FzrIbJS7HUtu9aItHsWPaEUlm2MP
qmHcPTmBy3109Bn4qeSUoTtYY00D6b7owAFzKt/jvGJlzOVhTaHucgwEWxTbFyjV+AqDRecfcGgG
w4P/XH/p1s9NQl9MvAAWQUtKbqa07b4CfgSbMNF5SZrJAnG4zhXS/2fV+CsQU3LFxz7UNGpJBgo/
Hepf15nXtgQofIGAv7eSW1Q8z+0JhSmQfj3guxIMPPwiBsU+DVFhupGvuxy85s2K34lhvwmuI4fU
GHfOwpMxUdsSUkTmzVLDlcE0rWFzEOwXGz7vAVKQI1T3Kv5OeACmmY3lwnJugCk60gkQM1Xwi0md
uJWKq4UkJZFhweqjIWeyqfUisfSShdzGomIV0uVzw8OrX3AwiRpxaK12oViGAwE1NtbxOo1wtYpX
Vz/h2CImw4l7j2u7LwY+gpC9aL4/0rkKtSr5HPv6GJIjW4mk5Uq7lsoDC4XlNM8iAo6fLiMy+PPm
4pBkXK4Iz4HhTH/oCNyihyvHRZP6GoNR30IeKcbT2E+dh6lkBA0+zx51szjsudzvhIn/77TplSy+
1uvwN6M56oMr+u5NumVbgZUP9TQfx0wQxGXjcjTkV2r+B5kb/NMz9nNiTUlWjQ0lNvEMZXiyfOEO
gkDiPyYLQxkuWy0oJGEvx0Uxl50RTqPikcJ6b5sk//KRjDkmLMiwFfnvIBsKNxYnw1RFMfJVLFxi
m1e5xHA/K19bttZsdpST5aPRMeDbi80c8NBe9WR01b6ovmyCIomC1/u6/3WRXORcbCye0N8Mr0m8
S0yPexnaDOoBONvSYCtPH00aPy5ASm1xUGRBV9ZdyJ+EiKXJJ2gfFUloQsXbL/G0URGDZI7U5R22
xqEI5iHSMZ4sKPMFiwXQDvfY5HLCI0Gtsic39kk5TRPm8Cyk8EKL+T7H4QAhPvSJNRukKYe/ycTU
7f1LDFrmCEB9A4zllLRKuqkFxOwJ9mr9J6T6cgmfwAiUtjm6BfC4Yy8ffgUVN8UJGyfVkzTTqKvK
pDtVpAKkPEuKYihTCZAOnuVtSn48KtL1E5w97sQTg8lZPg7f45WWdvpPMDArGNRFtWNQ9yt9LhIF
C9a40YCuu0lONwKs8NUUwMCIxGU88J3CpCj4HqlIs+8jcLu8S9HsiT7OSCUODafYNMOhuHa6poHu
j0/cfQJMO8AUHRkHO+KoVmPVKuK3tsrhSK9V4bAHSZo47wdmtOf+EoAjKhqLKjd48fHjMU+EVyk9
QVSdaxINlZd933V6lZ+EiQ+wxurFAK9kGAIugKkrjADkLBe4bPYcOCoF70ceTSo3XaIQO+BcmlTN
5Ssflih6mscHxWA26ZwP/GZoAlsWLedsW1V6bzM3pTnIQBtq26/hoBlePt99AfVDmgmVVf/3jsM/
8PCGo1+1PAwoYi6QuNx+X5Hu0V5eM5jQY9c3aUWX9MO26Lc1d18dzBPdpMd4jp/2RRxh0XUN5t2e
ULR2eABKwAW6v4ZASTsZ3Ahcg628XRj8yLu9kQ51dnYo2+Dv9tKoF05MS8cZbckdKMANVkWNT83P
lZllUIpH3Vfaj98enL2EJ729EsxHhHP32lZ1P/dsmOcEKeXtRmxesQK4Hw4Uvi8DQd1XjDfy4S+8
08dmI6L1Kq648DYlePvsvlZ8+8wZkSfhCnehCDJ84LWJUiKOuHt9FizTfbZcIIY5D+mWm+t8W9tr
qLZOv0GBRibHeRZBcsZRSZfO+BlMYYlNkxI1+LLh06WyZLU6N1me6LUaMd2EamvICQxzg0Ci+awj
UN+MsCVV415FcBtd+mkIi1lDSbqRAv3y5NU/nzP2CCvrLms21IDpCExDs96uM8u/EuDa5vpZ+bIn
lD5a/Z4qzNYEGBZBLa9kJq3ZxsyI8QjRZz8ydRLutwdwiBjOCkIoqjav4J2Uh9b4AkvEe6nHgArR
BS3OQj8lMzPKXKn/OgUBrcKui91JtWWkz4GHTXxQZH+imPhg4kjzlAH8mjUe1UcIMuzHrG95CCpw
IInzAWy761QkHicbnpFVC0kip3FlQExWWS+Y2vSUjDHpsOUP8r1C8tGsFXIDFQPmNcgVpglHRtrj
/grCXom44kOIMGr03Xwasap3t1B6/SvowLXYwpL6WSgpPj6PchJzadrXVI8Y/2cT0TpAuXDNBuPz
fYdlD1sTeP1VsNvlEelrUgxvwiXYLxtPNlSTLy4fUSq+rdP3jj6xV+9efxAZIBm11NZVtfi/xh03
lF/CZYpnXGck/Ket7Axwl7/mDGSQTQU6WrOH4dxFBMdHDiu8kU1cpDx0xNor2T290LdJp2YL68Mf
AIldoOU91xo1m4MrwwPth9hAnysTBI9QC3wCNBJ/Czh67UXw2NF3CyEQN+1z9LDXtzt6pzewQgG0
E6/RjIPDWsCNVV1kd3EltosLdlNksNYDoIupQ9oXJMCnTo7rqvSvMHUOVAGCT2lU7swOno9/iMqR
CKmJ6ln0Bdxq138v6nDzHFj4F4AZjpiZv5Pq1VMVihnfKT5h8j3g959FFuNEptc54pOyduMYjZGx
I6wr9Hm/n+DX9ot5QoFVSRcO0YV9VY4izWuoAie4XHFcjFEe0KG73w5FY1HSwNT4YasoA7xZejyB
Z8INIQLzIbrZBbfhNEyG6bWkgpSO9HNphIkPTq1L3npncv700CAS1YW6fEhEAc+/wbiT2er5CrCQ
AG0MKa9Kr2Vp/i81nsEw2JCwVK3bBZK4Sg/C6HtCh/NUDdAIM2w9Sud4EkKc98V5LqNLH2fOAE8M
734247SxRI0grth6LdD3bsNt66KtxGzwS9Kr5vDJ/CaJwCGNgAJPF8owsU/7+/0+kgwV2obfxAxt
Ikc+ASjBFHXlbml1WJwzYIelxNq+exNr2ANcZV00JgwG67kMY4bwSKv2ot9QCXzKeWpLQFtoZg4N
yzpZvAq8QV/weIWAAr87KPEv+5xegsxzY6ZT9Pn9rMsqPBtLzTbmyZ7A0+tFAj6/VNr/OV5d28H5
2mQyQUbGd5KROLhIIKdy/R4kGLAb0CTutRjzzeglx933w4zkycEv0g58MT3O7oTDWJyI3DN0f8lx
4gGl8V+grJjR4VTFWPXWn82nBEin+bFLRhpyClU9gkr8aTYWmBUwW/lVoDopICk8RhL62GtkHQeA
wZSKQvpYRqTNDSU6cfNeT+BnI/ez+KlNID3yO+Iuk5LLcZR2HB0zDA42gDBKJuRbs8JUzCI2UfHJ
A74h/PIh8AZR2vTIKE9xnDnMVYeoXzWF7HkLxNMlQaa85LFUdnpjdPQriDQLUXonzmau0x29ADEg
1pZEJ+TC08fnghwgYPk7rZ0yzIo7PJNFcqu2R0ccRziFF1Ag2jNmwLl0EYxqPpIFxhtZEM53hXwW
CRpln9IX+OP3TH2mYbvkLD6pyDBZVqYQIcSgdJrNEQhD5Jb2tWQeh7aAp8guTWxwcZ4Sc7kCZ0Nm
mf1LXihm/icnX8/TWQLQ532LqPZYI+aWZtiz5S2K7Ujp/8EP3rf/yLcH6WRf9+MFeDOItZl8RVW1
fGqvNOJBJYt/VDZ9SOmM58obz1J8jsikjp5BzBuTPbxsstZjhXMfYjvp1awq6xw2splNFJ+J/HEd
f75LgmvXmTZwOLKCTuLzVxTVvGHgvZbhocpeWRDBqgjkxFNtj+9SpWbgprDUpSktybsXufjz3eCZ
+4p9Kf6cp0qtJCeE38P8iWReMZrh0f5HXtzz7xJj0UyjqPnIPLbqBejMxSE6m39CU0Ng+qUd0gvC
Afybe7B+35Du6K/mzUvD1UJ205QJXDggU+ErMPhczbfDp0ea9CVZ7p40C0ytg5oPg0IpQ/BS3dUE
sspu9n+UdBSEzEBuX3QxUjBsy8+RuX3CYsNoq7+WJrd/y3Kj/hHmIhK/MFPUy9DAV6DfEnz8nMVw
VZHVTgbDNI88hr8CrJ3BXySXuD2NS8NOk/VVKVr1XcjI4ofcAezLJZZP+hWqt4nx5zRwO0E6sUFA
V1HCErAbcS1U3IrsCN8PnOv4Kv70q7gMi/9SHmK6tTESON9I8lWWyjHBKHsH4QUjIvHQfTniiBY5
6ZzcYsAma2nocvMf4cun0KUod15YmMBhuDaGakJ1KaiUoBHtDbryrbZ+DmwPYSWBK6WHzbZH5biq
RofUuQdTTa8Z4jXRQMZtoshUgtX6cyPIHcAD31IVy9xKN4dUtIa39A5jIG/HO+noCUFeAHuqhfSp
I6ItiKA58ISIJ5zyKhhD1UPcoJ/jPJ0WZLyAAZK9VeztEnR7iXmtGe+GO4eeUQWPw7kS5o9UcNIk
nwHRhwg6UNV+MBG4MxxHUX6j6/l8N7cKXplZJByGJsQdRb6gbvS46/iCMaOL5elgA0rgwPpsiboc
rQwxrt263EKIowY/89Xl2KeujZ8qxBZX1xtL7tdTHouCLDwRJgHiAJ6C3l/tRUBh6iFTtKV5uO5J
1SSBCs5MEcrj1MR+piUVttoYO0RwJjC6qw7CW4Y++rtZLw2YAkgjZrWyYmoX88hAxvSAGguYvZZY
MLgxsUWqcYySi0/aIHa/+/E+97+OcwyKcNugrQRfxeFwAZ1NlrdbBR7OCzbASbhc7TupZBtQA5/z
BL3tC/c7So/0HB/IHidpanoyp6vE8aQwFFGTgOskn0vX3M11p825BGWgCHi7K4KnXIHw7f1xc8bG
bMyLWXlDDKlFwENED63uzdqMbOTmJO4LNGg+d4taN37M5KDDvOX2B6y5sKCkZTjW+DhmuxC7BcdH
riDquTT+KT6esVDpUGknp0zDDADR63SCjgrTnqbDQzda+ZumTwqUlin5Se9sQPO/LOlsuLywBPNv
d3qQYpRfW8hkrWzQtNAFk0Uh6DKmjz45uGvIIlxA9l50gJHG1CPvhmnsx8PVFMiu3stBrrgGCfsp
a0+68frB45Ye3zYY5TibmTgqTD+EG6XgcdHAzklPfxRKNlVOhRJdm8J29QDm9+TMMGnT/VVAQdm7
SG+FUiwbUd6KvMIbYu2eCHzD9s8YxgbTzbVEq0PCwWtsaX6ocEmHqiDSOBesLg9QNBDTReBNBwXd
okPz4x3eEncsH45mgt1xflA7POP+xWB7ShJhkjN1boyHn0I53i5GaUOL7uA9n7aA+koNW0nObSYO
+RkuIewPxYhFJEVPu4KP112SmC01Z3osDofaR7WEimy0RA47Xu3IejmOJZUKdZHLXSzp7RyR8waC
pbzr8GzQBq8IbovLK+gp9zCg2STPiCBstTHwq/dVQkKt1GZNQNXwIYUdv65kAKeLJjBomTAtu8Il
oGuhsBFWnTS1MXptJfh0LCqY9a50LTlHZtqxJkQFu0/KK+MdmZFZ1UsW/ELmKC4oXmqbwL6qHQO2
RFg8xiXmssWIbS9VPtafBzxbuaxVKUHaUGnIHBFMNsj/rC7sjsSsGUOcpDkIn8EeBvsxQsPS4Uly
Zt/D0JGf5l0XPRUkARRANpDYuO9fPvREaa7SuR2Bc9pAB2od+g1Hgv7I5hIv9qd4zEPG00wB3RRm
V/DVq4KcTpSw31Co+w3YJjwFHRqkbNDprMUwqyiaaWQVviJZN6GXu735rDqtywc74gREEDXUYUzB
wRI35W4xDFQ0KzbSkeREv/fzfLdtFkh53xL9Pm4/NdfFhTjyhXwqR4wd7Tz7wmx8E5+i8oxlJJVi
gPwmFYOOz+2wgNB/l0uZCFhvjaI3RvAghGihnh6m/HkMb1mH5TgPBTvnXG50yAYAjBPRNea+TbDb
XaCQ4r6y7kgagSjxapUuQAVJ3h1eXb2FmdOMny0XJPkVwGfIVUbtF5ZWXEjbVh9zOjSASMDIPUmL
rPjSdjtGQ6YqlQD7Eh/8jceQP7G/wjNR+Y5QUOngoM/9f9oVEHCLaYskwDWGx7TTErRSWEEwsiPr
bUUIF1o7FeRzpWVj5ZIhHlPv89Hpp1IRNQDXP5xhzE666qH8kU58Vddc6ufqrayVEHASWNLPMcI2
AYvUQYN5+nFQtmluHM1mGQMKghuRjfSr0gtKNAjlioM5cDK3L1svqv1fagxj94uysljcv+79RhwT
lcv089rYxM3cbMWm9NGNAeAxuoXFE7DP8FYC0ZUn4nuMWzOfNWug+5ySmecFl0vISdEziyvGZCQw
DpzI/GU3ADkeLArmNC2dHPBFltuoggbbrnMI6DGVoPTnCpBZvTikpqz0n32HC4O3hjYyhgPSXnSL
tS6Yqq1BhvwMn8DtSX5rFI1ngTNdyMbG6JrN9nQm3f/sCgyRTH5ID+JUDobul5sU+o9zk/BC3xit
QFOOlwIcYIJXYYBAKZdTZAh95PTgb5CiyH1CSbAxuObNOSRJrS+LFkQDZCZMvI7wBuHyX8DDXQwP
JrUS3SvlmkFcIhmRt/igFwD5CSIwpwrgIz2ouRUM2Kgr0pFBdqS18QTw0h534psSgri/VwtWyufw
t68CaKU1U+vVUGW7jZ6E7d38X44EnRJDfF8tAsGatSfNDzfnO/8fcRuVRkCaE8aFu3DpXQJZ0JrG
dgkKwiU71Rn0imvSCLHixvL6TYIC0Kec1N8amtj2cRB1SgEAb8G18XGuXXu4S91GxO+tMJHrQoXN
WK8k+RTTahzrekgO7B7YeVq5+hxIVG8moFSIi24YXXOBm0jeLw/428UKdt0AmM+uOt0IHga02thN
RHj57CwCccrWBLyMCyh6IYimtWvAXRkUD0x255n6em9JRewSxGHAFIfVBcWWsETAarbnPhF2DUiN
bfBgMye/hok66xWTgMFFKR+VM/jFS5TR+/xVznImUA5NjaN/N8C+iD8C/rdJN5e9ix8pnSdiiolO
RrqaJTJ4oyibP9Ywjcyae7/qwaEh29WrtgezgI78+J7PuOyi17izd+3j+K13De70eV7refzkQ77s
l79puwnTAbeDpU+ZfUXuNBJj9V82rSrLNxrYQKk/CDpfTgi8tJxwDGVGRFFYByJBJAHxpOOM3p3v
luTJvEEvzOwfVDN6ekii9zwzTWtwoZNCEw2b7DGVp8Nfqg8oR1UKN21MDZ+DboervBhrzNLpIyKV
1wmQY4k7NpHNC30jC+cOou4/mB9cnLMwACr1GpZlfuYxla42YXXg9jRp290AXwnzox2b7OiKYlGw
I8ORGeuyHzSrDwmjJSqaxBKGlvbpMTk2G1ZBQ2PAwrFBh74MNd0W5rZ6aupA3xMPUCLEZIUMA6L7
LOB7eorFalQ9Dq8frRH0rVeCBFLq/M3bMNZyyVtw5IV4T+jyKbr8puOOxMUyP2pjLMJ9NxF4FYp+
LEsam6qXVXZa9gie75UpMXwQBuNqGZCeThrBhUCFGwnb8BcxLo/TXFbhnkAVpI8NJy0VKKB/CbgN
jFPfRBLFrvt9trc3bZzqQTZhPW6ooD4g9dinPhfIk6MRuC57ChUAbAYPv03ZvrfZwdF5kA0OO5Zn
97tRn6k/cKOqn4VTOoNI0BCsgO0+cV3y/bkl5RlmarSHSCj94wnOhjs0yqRkLcUBZw6GvGQMFZHw
rZmiMDKigl27zqDbI8/BiwnmMctgccidDQMs0aXvjttugQGM4y/bc2wTZ/RXxCDHghbpMbWnlGQ7
hmw74HG8U/rPv/4qjvUt6p27JBZLcyUQ/+GFk0RHUqwFqEMUo5B04HIU4uJADoNd7LuoiXdXQly4
KCZUr8TQFULHYovvIcuqhqeGyThoYmvliGjO00yu/N/fVfEc8LEGCbF4xp9n/JX9AyvXyhv+Zz9S
Wt1ABfklv2eeXb4gd7TU2CdgAE8dWvgsJsQobjMkWuxKowLFK4Zg+L3lXiW4JXbLXxYr/8kUcVVY
aXlLJSwbTHqTXkd7mFFlHKUAb/plfOU4lWr0qfdvgqs5qfr/EgSTmfsEfj88+27ZNW2xF9B2fwpI
uQjSFUYJ0mFgh7T9MtLUmUJ8xU3033BJcW9zCcLUjQ2kbBed2s2pyhrkSt9Yczd7M01ZA5/g0TMt
oRmRgu6SyYyzC/U/xOm+hbGJ0y8B7zGOhGmTEryOI30Yc5vCK+DsNVkpEDlfGnwKvAlEHpDYvhp4
JQHO6w4axPJggnfjh3eUQruwsiQGwoUH/+tCSjwc1UYk6j5vski4/pXz+6uBflStddwqgKjgmIEs
CvfWjaP2brHDBJXR9NODr8z9bIO9SM1H12svHgjbTMTD0F4lDJ5i7Aw3fukRQPoNzoEmXn2sonc1
b+Sr+fxEN+jNth562QZAOxIfsTsORQdbiFUJvYcOsSIBn0WDVLSGWhNFBqFhym5CorT5W8RQ6p4M
Uk5wVYX3sIJu4x4aHGlPlq9v4fhJgqK2qUD3yh3CHNV1IRoCVtXhtIXfV/wMJNZxA23bKik3kgFy
IrY5kP9imRTlu2yiL8Dzxrao3c32+Gyujp/rLbHGMFO0E+ai1Bkc/I8iMW1uNFsitVBJyCPjTx6g
xQo8zMzQ+JeiKU6vr8q/aBK6JSqmCsEkDuFpuojiiPdG8hvN2lCuThVJpvRim/7v191ohnx0tQ1R
xvtOiGydYdRsf02L3GQjWOXtzpbTpnCHgHFMyeZnQX7zrJWPJ3WU2pkw0N135O5K2//MSmAglloL
MHIUK50FUDqDISqZX/TpuIQLTj6z8COsdXHipu6gX7Iu718gAe5UQjWi5IftR41Ez0yLWA8icady
dzzxm3fVLUrGzzFr97T/mJlMq/Zl1fUMRlzdilxGapHfZwaITFboEPC3tYS7es3iLT9vTA0lfRPr
cJXpXxmWmv3qAyWloGSx8fT7RP1OU73fzY7GSq3pmH+GLAw2QKHAmps1n1wcj0xvY+Myu+bpS8lJ
KWIN02Jv0Ecqg5a3ACuVPaOMT9qzszdhVU1hu5IJgZFyPE8fY/7N2aULMTlBdxC8bq2n/jz9JGry
WC4INlZFbI7DZspqKD48rhCTJlm0TbPRpzGrix6YkWk4F+y0n188VENV4iiZpHdnbg1/LMqAjdni
8+gTN/M4aPeAYripLBrHoBw9E1V2SEHDxfGJ/A87PEt4MNopyYS/sY9Q1a02QKjAU7SPUFbPlXJe
kXq3XtzMsNg1mViBrd0Y/U3pPxi5uABuUuUZsUoLVl9HSTiygKlUsEwAQ31QKDyQTImhOvvqlLvM
82DWTCBRcm37APl8g/L8ONw+pqyBVCQm9oM4gFQAMaLJK+cUcooU2Vl8oEk/qztJtYgQLGjsob7c
mapJMCl3UGJ3tQ5fDE7A1WePlSFi/tJGWkoyjNkWtK1bZitVO9n+l2dDhz7fNBe7MaPN4pT+hBid
xajugU0otH1mSXH0sRFwtXwklg55AnSaSaKSBfoXnxw98kUTJkzY1oOztLMxGR0jrnggmz+2lemi
YDF2qOYscpMIPq+TkVUapLPySJo2H7W3WW7BTwUu4wS3ektIcURlYCk0XRE0FiyUEeFDaTwML90M
RdFhQJ6vkZN3tkE6pw4Oz0pPMziicVr2vHlIneu7WcTGtXLyepjSD0ZtU64CGbRTLKvazRQ9twRq
v89YWSEvwL+O5XQN1Fpskdy82FC13An2zPSjXzYmyj3U8v52rXYyIwHlaVYSubE7dpn7qxYmOX0P
wVeW+xczghp7SpQ4+OpWJfo3QnCLyH/mESlB9q8iv7ZZhj+NqIMSQYEOaGZM1ru908j/Y5O0CQXg
FACDI2Pmlm3PoGxtMs3yZPAiUvgjrR9pgWoiUUp7QLJ7odjHQCc2eMEVOTMpgtXdGKx4EXBCo328
QqmfsoffczASdEcfrKfeOySPGp1NudBd5XAD9kgAOZFfOwQyOKXAXqmWmHNMcbfxXuErKev4C1r2
qBvNC26niPLSvHI40zoGDwW/HhxhgXasVCSwT4+Fxwu21bNDrsvd/EopvjGh7Krg1bjJrQLl1Fgl
p+sibTU3Km/qfg3Ddwb4/svrY9QlmCxx82d2ipA0n+J/aobzaPcoKHyXwxmpvM5QtRaWSafiovw3
1IAsiUEYc+zLt1IkPBXsSJAs5DlNQy5B2+sEP8wYF11MqSv/iFAHnN+YoQOX0QCEJ25pqfiJHwiz
0NCYGLNt9UCBqz54seY/6hOWxY+OPI6xGfEdghek79Vs4Mnttb4OXnDqyqJJ18Y35/qdjKQMGPwV
SZeIB+SX/CdkRsqqXgt+xL//HbgkHh+eKqyIp5D+nCF7k62qEcpcTSWI8U+rJdCPMw3cYjhbixxH
Sa/1i8vbX//3nWDYA7lJhVqC1FB9x9TfJ2Qkeg7kwjP9/dsG+frgGIkkHYUNGlXTxCBp3Uauw0nj
cR8Pl7q9GI9je7NsdghiysPljfD4xeuLyYV+g+nlyhpEjt+aW/0UQI1iQiOC0oahPxYvleLEz9ra
ciHu2j7oRgNHFtCxadJXv4nrVkgR67SRaoQQCjBCfTMQExrQ72322XIQohqJbhjxWgVp9okIJ6Fk
Ohv98w4hSct/kTutQY3cHQmQEQLepDvnkAHB+Mnf/tvgXwEQjH8XLzhxemysiJoKOfH/UGCqkUV7
nCZCfiMqFbmlRW0Udn3krXItz1Ke+a4E+2TTqSuRZa7/BMd0N7AZW9GAlwtYLaC6EEVjFFJWGzyz
pNsLPBNojbtU+1VakEwCD0VlzVEjUtiBwEFRynH91a6b5aU8OWSKUwTahXT/JeUxxdomMynHEcoM
iOSiWlXxNjpGwfDVRfe6mtrvWWYoFcuxez0AKSZDNaQ+J7pjqeuJdS4h9GXfDavP0l1Y5o1H8okS
OfYR7U7bKdVs8/WwyPMhkY7jUs42kRZbTYyF5RCBPR0I4TNeW/lEmycl+0S9Gyj2HXwYmxaSKRpq
XdSnE+JLRD/guosNSXuahknIENrTKQvr9Q4VZ6e56w5RyqV26N01OF39Ozwuy4C/0hMZarAl/ujs
0wN17WZnAX63t0l+x12kpW0nFw02ms1BXtbvAPCB75XYGiwDbYRK3rOyprzq40Xrq14DX9WL1wpY
IzRa0l13dhMECMP04l4nWNhSXMbhiEhxx9Q+4TKBtjdbR0fkjAojaxMwjOPWAM0fPhXlpHQ6ZpXP
8uu449Feb+clqWhoXARchf4/uRW+jbuact0nvbJTniy7IXkB4jakrM4uayBr6dCEJI0wE0NJQSf3
QJCRN9wGk2c9rkUf3GFTWL1ZwR0xtDtkFHWeAYdhZVKeWM4TV4+661AP8uaoLhRDvpQ+/pfIRHEs
ZKZz8Y6T/Lqj+aczFkF8JN5+2dJcltUgN+rLZGSu2YKS/r4h6mQNC7RZQNTYXXKWLLqlkBrhJSaR
vnriG2Utq6ity+LvFtFVCaagH9QrocPIaWwJqZLALNqWq4ckiZfQC+r2G14ZkzFXsZ7Wxm459xaV
0DTV5fGXO9WBinh8DWee+Ocodq6CQ17o/JfdioVH9TkRbTNuuVa2CuxW3zEESC+OIwLOfteqDeWD
IX2BoAROD2uRFrupO4hChMr4cy0DQL6C8sLlA5OE9AUJaaHWlh5vSo8vDEEaDX81Rj+cp930ijkI
1Qaudoi++uJov7PMOu9I/3aYGTADJMJbk6nXdDw7DjC6+eFqj0KVrgW+UQ+gWGZysF16lELSSLxk
IVNYP1sl8hlKpal23MWweiGgXK/J1GO7XrvN8G6nOAUkupq2wo6xXiWt8MjG22jMy3n5k+ojC7Yn
DDLjD3ZOMES/7SJjXOCfywKN5EEuD9AXmkC2Bb5zse9FCc7R23iTOGdS7gjB2Wi4QO7f390lDzcx
X3iWy83Oj34GuXO/oxh3X0k/NV+KxD/OEn30Uh7n/OUTRSNK6cjVWy4t7LgmjKidh4pmFcfV2Mi2
EuFV2Vx8cgsQdVnOYMo9+qqlAVtwyShkJmoWCvdKvEjK2epEWTw00xQ0F/e7iWDOKxthUC7aP0Xv
IhzJaxXqUC7x5LrHtKGXHpa0z9ggkjuoSUfXSbSvrdka9CutnHTUcEKs2HW1uXCIAagEU0Eq3v4N
1uMlDaGXuXHJSdr9z861mjVY7n76YYfEEjEmpwVHfNOClTRXGwz4E14G2343EVYavtYXorqpt7uq
OBpFCo9QfdtIvbBDd8MRlGVBj+XGm8mAYXW8U/AoJruKHhYwJlz2/c5N0xkqMic/kv3v2FnNdPKH
EG2isXiRvT2TUa2RlphWVMChEFf/pwpR8U/ELaNIaw3yXLYz9urUWeBJYmWOf1UenpBNabYrjYxx
BmpRqgJIPbn0JDRKQyvVjGuO/mxPoDqa+RG7XPhaXT1c922mGNgF+ozM7Njx9gCLI3IC2YabgWsg
SXDoRfq1fRtZu1PXx6YTpBcmdtmAnZVVaYAl1mpScEbuaiRvTJ8Uc+CozkZ0N196gnfOHnzzjrwz
/9wsmPfbpzmxT69eMpoCL9xUDMRwbbes3/FOyeLZX4tzQ2ofY5b8ocfxK08X+gus//By4m8n1wkq
BcgWDyecLMDX+ptQQnvvNmo0ne+gzCxHGzYAzTP+03UBB3I+A6tB9b7uY+KulznG9EbXrTiThOr3
sg3adx7wVflnwlUiatZ6DhkwhM9NwRq9UrsysrKVJuklazcIVLypaN6A/FQjicFYBeC+enYj+FzX
ezJvFSDI6CtmQd3yIyLxT532MFDGUcaNVy9ZEzuGUo6xT2Obq6h9t0uz/2S4tCOd3jPCdJSk1s47
h3cVquaIyOb13H/mgEEP2X7Ogx+ZKTpKp2yMD/+l2j0RV9YkitBp0yvAEstlKpSsmojHf6SdNGP1
DHKiA6Ey8iC8bCZLeP1VEdFyBwGrzlNSPvwt81O8R+whG0h/is1QSRSruVkGjhxfIAPRXSxC4eHd
MH25a1R8xRFO9s/EIBDA5nNsB5+Z4i1ZLLVAE5C1Jv0MVgGVQjXs6RiVbbFqCBSF5QrtM3FXkqMt
pG9nkStznUURbwrWT3Lxxzlts0iE/86ZfV/Xq1+yIiEusnq5x7JJMPOrMnmAxniNVlMrlpOKNbqj
M3tebOMvCrq6LwgX3ZnpbJdJHIyOosoFzzZqMPme+OPbmHnlaJKaUHTRTe24PkP/gllH4SJLCUI3
9VKLcgZdekdHE8DDaMenYaTZXOsXLu54Ub+v72pLPDndoajFcqL47yn9fyEsqHiV5zNRpEiwjmNw
4S2R7DdwKTqBTTSxpzv+aigIoY6NfdbFoZXi3vsCdqkVXRROeu0h3o8jGSG7p3VpL71U6esDvoOk
UTX41xPAnvvOf04p8X76+tv02uYlerhWiuKMMosWDvJkNl7rvgIb92efqxQENrCF+Jh4aZ2EZE1u
/xL38qsqAk8P8Dg6CyRi2Vs90iWMssoKUoYaXmJLZ5lfpqGw53+UqyM6VDooiz/V5naW/8zmtYaO
ob4iuqTFA3cJI6vErp64/nOQbmTTs9RQf8koNqADjD5Wv0wMzMDVTNjyinfOvMjjYM8gitPvp8og
kCJQk+4cwiC/0qL8Apf3Wms7MyKKO/LAVNa/fwfA7BjWabwm0zuGYfeX261If8gImId+LUpktkob
/jSMKdpay6CO/vVst9oYgk7+5Vn+19jcO91gvLXRqUmhJc7NDSMnNR05Ps0i7X7nFtwS41BbtIIU
WU5/DZ4Lcwtd/nb6zXkuoeg95tSz7VzWr45hlqztwD5MenXrOAJ6ZcNLFhd0MlOwVWB/9csJZsHS
lJYdxKpwBvTF2DOh+t9Bw9qOBhOL7QYsLBil5q0gKhd/Y5afq9lF5QGphkG/GXhqOaak7OZeF/WI
S9OWWrGXq7rLDdS76ohkDXEl5WpNsgSpD2hmv1Bc1AXrifw0nEC/lLb7N9tv3yhvPlt+vj7D1u7/
mjZiockhVQnkfJo1dycM9gWfy1UzAePyXSar0WyNb7SIEZWoLVHGvnjzm7OiZUyKMi8gUPCNDypS
NHXkzlRphQrsEoAJFWjuwBPZ5lERzkxL1BHqAU8gyRzmkpHa/+UFDhlRe3KDOuQCEh2pl7rMHukh
7GZH6Q4bEm9KHp5wk8LfR/xt73BnHwxV83AmKw1l0PHwhT7ZjTh68L9496mfVrp3FzZP3VHcpwgD
zD25BZeLr2lzVLJBPRUewBALk3OpRqvYf7rn1w0SlKLm/PwgQVsfh70YKMPaasHjti28X8/xcaqA
zKjlKa/cGO5nePw7fMONR1jMx+ITtRQa7gFt07qwV7N4K6P2SU8AZf4OQ1A9wFmg/g3XH6uzG480
j8ry1QTHl0bOhzI8mGFWf3QiJayN/VkzpbNTmH8/acT4C4EcsCdKCPV0aYNAMxSOq65YJzA5r9eC
x2+fBT8WA+p8D/62H/FK8uS2haRBZvlmzcEOBEkLJJZuA5rWW30oqbi+b6AlBM18eNUWxinX2gZ8
3/TkL5xJ9AA8Hv7EIv8DRshNQ+wIL6ERT7LrTTpgvIXacMv4oh9SRhkE5ZcpZ9iSK3mTipQMXuel
0VRUT8Bq1MbzARnwhxwP+AWs3iAl1ku4n5GxYdjGd/PiK9UYhuwbQKj9v7EG/hZE1sCrmy/8+MHW
WFBUr28VuoLul0Vv3RyELB3lRjYFWA3mB9F/WeHH/zMpLme1hVLcciO1hkX1F1oaSz9IsGSW6FkK
QEkuM0CcdzTpcEIicV6AfD4oent/MyDBWLvKmjHV12l6iJOUUGYBeJ/kqHROhPQZ0SHYGWQa2p4K
64AtZjfxb6mqQBV8E/QcJEk0GjDgEA+Ky4ixlQFIRhYLEEnbJHslTqowxPCKHPSjqsgpptKFgqlz
z2OjSqTBGM5DNuAmyx7yfK6QxqkGmEnI7OnjvOkT7DYb1B5kHYWWFBtQJE2Yhb84i78eFV4Dqg7Y
mQuugWGe7sysoRpE234gigsoSpPAYNLQxNBlArJHHssEHc4aByDmVuy+y6Znq5/Fb/EssvKuGjPC
zIoHqWV8h4BxLJ+ofp5ecJ0H0tMdqVpVMsdxYwDeJH0DOGFl3J2I18+rCFFc31k2NCssPp/mQsYF
EgYBTptYd51qv9YlhvynCNa/ibIFeru9U/H49T39PU6+Kap9bjL0YNP6xsvgxlSGdbj1Rsv2/apj
+eXlxe6uFzIrJGx78NLNWt45K8U2ErC8JwHFvsAn8zSLcAFvzmMV6tGDdh03WdD5ifwoT3hQpM3r
YacIHx2hGdt4kuh3a8YkNy4Y+BdLAwNSeY3+s2N1/Vc8YhoKJI4lCbBpi9kWcnR2hAlujgysWYRy
kRYu4BxJUd+CiT91NwnNAqRaLcrPPEt3quMsq9fziA7Zfovy2QcHlWHET1lHYO45AoEw/LFEzYBE
YCjDPmLwCvA0DRIkGlxGMEehM5RUMZUF9mg0Yt/jILylQYQciWq6Ephwn2iAC3M27U7Du9zipsRZ
Kbe3zkkWoNqu+415r/oNZk5nVe0nWRxp+Iifn/erJVcA3IHMBe9vkoZjXGQh+q5S3QUGc81dI1xP
nsXOu0p74+QbDG9wJwn7Xr7s5URoYGShqzfpBd/0bwA5L3AorS+S9vpY0qxThdvFrMU+jgK6z+p0
VADIvrRuQs137Zow3KYepzJYW7C5Q0bOVm4ImAeYidoyhSg0f7ToArDr6piKk7y0mlrVr/lIbr3Q
eRG4+aMxhC0ZuX2T+0YFWvHCL19c98Y6Nxi0P6pc/ym96FQNLoskmX8GjA3tqMFnAY+vO4REz4qW
GMOQPaozRdrJ+vY4x2rrZ3/lOGsvzLKNNs3/Q+MCQyq56Tl15Te/8EQOc1Op9HVLqq0FetgOlBU1
2ed7XRiGKgaChsm27UBmo/4ecu8ivw5QJe+4hXqwFWpg12ccpbEjIsaVYXDJUJEk3r+ttnCiou25
yiU4Fc1s8tSR9LQj4fanLQpEKaHmZYXdvezQhia2ivbA7YXyWsrxn4GNKXTn2XiSz6D5dAG3uQII
YdTWQlgoelMsARCMtpnlsbQWUQGUzJ23sc0YkOPHoBQDTDT5Hn8Mv5w45PipB6zi9DDO5ZMz6/7C
1FNU1mg0RrcgmAalo+C+LDSYr/Y4WlqRwZz/YnmNrTQk1ECzlbpeHjVciaN21oE2w6ojGNqNAYqf
CV5qT4wR6L1xojSiTCvopdwqv6j9vYe36j9bgQLir5NCXFQ9h5PVrFWfQX7zrRqJwQ/AbM7zcAh4
BAPPPO1RGYtjlkDqunLrMBvMEgNxZlL7G3V2sgzEG47gf6alpxJctJrLVXmH2eKJw20du+ykoU1r
Up7cTAgWYIGn1vSbhA0RNx1A8cyG2gATa53fWTPAsfDwsHgWd+h0VwGYW0ZR3wqAgvfzFddi6mSf
sX2uRU89iyPTQDKGjAmrWVUi7yOVUGZ6vEVF40PsLo/lEAcEd3ZVidC7ja3qwx0ptK8bIXn/LWBz
b5ITQ7K76Gd7o5PRD1bFKRzaNJB+0yqhziGM8ONTluouFkClRpJ0MBkVGCs4zBHt7UgJj8cm5/Tq
bWIM/Ff+EshEvtOgCm7qAq/8d8tMNH2eqIxqnhHNJY51eaJqb6Ss8dRmPdch/Yqhu6btcARO7aP1
HmMsY8tCiNr1w1/+nZej+cPptMkPDptn1nQ1V5x2ASrRy3nBk3lOFFQOAXTcDKsczEK+KEip9O2m
XsVkJ7dj0YNm8yf/gk9rK/4SnTwdN/VBxVqx7DmU+7DpmPHU9HIB5KLqp7KFfpHGkTnrQOm1WcFT
DWFahRhiv/rrGJbSXD/5sSBFwYsxjYzxAo55g0MGz9O71T5jTCygLdVFxyUcUAu66bWzFYn/f0fi
GIuU5BdHRdxX3uoxExmm6yDWut+D3zyssYRa8oOTOVFVvoxLKPTB4e0ZhT568AJbMOEmp64SBNGL
KyUSmWz7CRMZDjcwO4IBq6JfCTCJQZ5ccpQQ0bcKZDtSTk7gz57cAP+19O3uw0Kb4Se17nC4C3z9
///NuJQysZm5aGwItAvNQYNhowWJi2ixtOYbhuXhOqHdMtLSc9YDzk1aLat18GDSeJJhf2b9ZYFp
SrlQkio8QcrhHg61Z5PlybjkJwBvkwGSprdCgLAZs/6XL1nYwm1GTFXwPeSBAtaQVq6HOZjlJtea
QYOXlZa8BmojqEkVt529AMzkbrnw6hOaeDDogKyR3Z2xhMypS1Zuwre6CiAhgi6XZIlahz3Z9LM7
+ObZqJPWaMokELLiqqSeciLHr475bL4Rqv8sU5hlu+eVN4ZCceb+wzl7jut6Yhb+5wFoCKUmO+MK
VL+5XUbaQIEF8c46VOLJX5sCsjGT9I9HU9wxp/YFI9yr/YVXurGPvdXfxymutcqpETcxJZR/0XuK
Qg70AyZZtFZr6rcEJTuSPWXPpzYCHHMDApa7dsZVeVlrpMXTG6kZszWXroPR8zwCQAzPVtF/2hyo
u9/Vjd9f2Z9e7Vf/4BbMx/NWc3tCIyZZCGDOwS08OSNtEVQBq5WqjBwmqXDrMFMaWtwCEGDOz09f
jaBH/LeR4zbGp0G0C6dMwb3rs0PpT9Y/2B+XMbRqWoQ6EBD/l49a3BBMBZe9r4nIBwGemcyYFs4x
STFB7pKQLdF7cuQxG1LUSU6AN0HoyEeiKbzIcLKuASGquxnJ9tD2PlpDt8RGeS0VsQGaQjVJ7xoV
JAHdrKH4OM1m+jfOXydTSmXRkrGaqsNK4M/10Qrw2VYF8a426UB+kixKu3TA7kzRRcCKW31ZVcdp
6PEZXnKAaL/yIzEXhMQ+RlRGvduVokAKR5SHUGFOXQLlNKluMtA2YBKT6UT2EA6T57SEbO0JPm94
bl7fwgLe6F4ThUJLtbtqaebDBHtL7YOooBJyPaMiqUrkEtW9WhfuLQeehJ87YhUWyw4XkeUl8tDm
KTOslT96bAmvfSiLCZX6lD4uwa0Bz+iM0K8HpGIBro7D0XkoqqftdWmR4wwPYy28hPbKaE67JVNU
9OL5KAqBsBtp4EZaEvSiiIfXgMwfPQ5wfWklgKmkQ98KiVd+tbNkwb+A2JXXizGwu1n591BuSOY8
zYFvyQ63AqOSFtt2PCHG7zQurvF6766KZ/dDgbiWU8rMHbkaQJEH6tKZxaJaqWYMRNGSMMTooeoD
9Rl+VUwiHp4BOX77h35hrhN1lToJeSSBtaIaoNCKbi22Xf3jOVX5qdb2YTgLfDJpEhb075pzCBzp
KCXhczuxoQOoM7mowH14kc0sNbyRbcB7y/APqYusqDm7Sh6y/f/4+XQWLvjefRSNAUuioe2ZIMWm
YM6WlvBTYfhIpXH6J04OXnWwwGzFwZjjAwu/gg6VCrsZXmR4855eIdiptWeD7LXacw29QhuMBW4c
91oZYm0zx+Apen0LtNvFXI4QV1/n5T+RPHfjKT7CpZo+8/Q+gzMUNh7Yw/NxeZImbmpGk7jZfJjO
wACkeOsTDjqZOv1LV5QSI0i6XiB3PsuSMzvQNowiDqNS5Vh/B4nzvYmWdatdWeGzMR6q754zQ3C4
Xj/65ZkCcWwGllypr4KdBETcUATzRM/yzTg/eyL1kRDX34OQ9mQTnkv8jWdVwkmSVo7IsTGCdHnt
jikKBFZGlm9ZgaxQJssZItDWT0feRacYIQcPXwpBnq5kXC4JmWnfaiesmU0uOcmxKzinr5FPJoAV
tQwKLuKM1Usnw3ZX9Z6TgVegJzJ3/T6pvocuCEu+wgFy0DEZ1xXEe04uNBOV9CzkWFN5kY24lOa1
FKpLMOBPqmuJIqaocLyucUHyCvXXi21Ghf2SaeBGXbT61KCVgZhKoESPDCoJVgwUVX9MlA2HKszk
VDVlTSIV4aEmL9UKtTtbcHpQZkMcvRd9d6Jg1w36ZMHqwwge2hlW7J0uricFuvZg4RJ+a7U16Xzf
DTi+YMwSZamGJ+KOfNljFusE8otaa4h9FbXdYkxLS4FnQ3C3jSFGu4gwwK82FJ8pIQ8SuWXoQiP5
c4tO72Vdpbc8xzQRAvR+KV2qW2v5LFrDv+zaZ3pndJ/H/PbLindTLkWL02pN0/yj6c2pJk3DcI+1
ZHhF5mebw8wQGMLGoWz8ezHfrt7hFc97XnmUignYpDBcCmMcNjHSktfOFi9Sxv3joPYlKEdSB85P
mNmr+VGQeR3sSTYjyEmy6+7ANCajBQv8R3xOshxvZkBlETaWiCcEW1VUvl8OA+MJ3RTuBv04VBBs
AKRdPt33XHjN52rWNP8fZjEtGHt0NAIz5Z8UuqeYlr1LRBK1xAwWv473kELjjAARn49QDxeF7pJ9
p+B/e7VayXLfTWkRngB2OwQniFpSjDbcjeFBRBCoR2k/fAw2X2mTdFyNV8B/MGQ4N5gEyGwmVIFp
dlgyPc1r8XagnPtPsUDqHJGCiWGRa370ghRWcpSG7T5D8PDhAchiI8NmYsw/39lhqEai61BJCK+7
qXOmwj2KO55tPUMdHfiFVfcYefie56mRtqBYO548axf7HTPLobtmfnVDu7+aiQOlayozwDWwqLJ5
kOXZ+PRrzFgeJVDp42xkNcEMJjQNbqhSieppwKPTgMFc/WycQpJ/FjM/Rr7eJnNHyCYqkKKm4AiI
pyqfcQIC3lZ87D/yEAOByGyPaAJhh/FNnCQIMy1x08I4iblqe5ETmTA7xihVT6FyzkC8rO92uUXi
VLA7DZmyCEjozzbuvNP2BWLN8w/HbCUBpR9wVDFau7rVyG0nEW0QOQnXKP3YLqSs00X7UuWWlOaG
h/iffSkM9ub4/m/VM3UPhjWJk9CSsg03TDUFwgx27yfImAGfM4gU7eKlp+rbkefGZdyLKVJLhQTz
tx10d+lGGyjTPJ/ug6kzTFnMtotczbM9h96kkmGYYE5/ll5tEHzrKZgSD3PaSioDrcEMmBer0eQw
1H499wQjnq3bavAY3KRtR/Lq3ZJ56DYToa6Zu/eISAUq3bU6II+da2Utw1FUT/EzHlE+bGUCrPpn
prD9A6I4z3BUM4Or5gl9tyIuHFje70Ko7IPHTQ1JAsecLtHhi3/qRFGMExlAi8t8kGVHoObz6zVN
nZ3kR5I9yF2T4qolroTTbP2GbQuRfE06i+U5akY/Pij4eXjNamhvLikYuzLQoMIsItp5DOXRurNJ
LPIaNWrqHls/SAAhVnrVdch8Zq5bzziua+wzvNNdSRhU4sz8R3UysdUranszlsR3p6/cxtbUTPWQ
btf3acOw7hP9L9n/XrlYnAIrFbRCIvX0Buy4FqjcafK9+PyklaA2ifdm0Yt7FP+z4kOuG1x4c+4v
xEr9xzTpY5wQeJvcPbxseohsOwDad2qTQ/vyCqi3mnbzmqbrpNaTEgUazveWbzdUwmOJoBWH2DMi
NrcPxh7FE8Uqw3Zsp1iM9GHsla0PGKGtABsUreZoWOIxKdEPLOYY8aiIv19EA32ERWQcuvkkaBbQ
XX+I9QVQzcyw1HNW3LpT3V7Cx8GmPuZko/MXfowUhwZdsxmUXX13kESMxSGvrbmAOzFHomrEi8zs
cWC9u8ZW4fIIHXx842vL3K0xXGxX88Lr5B6RRrWty9Rj4dJ5Jt7rsaQ7KlfjMUuJred68DD1Uz+z
9/GVVpTZXDJyGiSsXy5fCVcafeStnblCVnT6KYRBLn7R78O22ydCKUtnobRTtmRv90mGMSzfhLS7
iBPlu4XzXHUDqJ6PhZIK+3fxztn9blpBzYH5+d68b0/5ZOnqeHt+i7pDToADd3DAuB/myIaC5hXI
0toXGLj97Wk/zsyQncvJ5P1wtNcUDc1vPhoUyPVNYV5qeHWW5KHwALu9T3oc+cd7wDKG908wzDQ9
yvVNQH62/Jtb12gqa5TRIlKNsZ0vGHtB9gcAaiTqzd70UR0XCXq7AkCyJDgQJWciRMNCaEHfTX8b
dbje3MB/7jaCksO2vetzgqkj4+KMkxGnSPSp78vQGLEPX45AMznwhByw/AIadQVxpk4kNVDYxXKS
wgwI9FuoCESzYpDbjU7c7EQ4zI5gYZzjV7aWvc3H71uqs/qm106q3eumVOV2V2o1GJlfiuzaQ3Cf
i3xLm9/mG5/OH0avAazwcCafh1tQlkAWYeXkvlyNx05CTO6IC8e3m1ntiqrkrwKHiLn2kssjayDJ
gV/JI6y3JaOVhl5Ea7vi9sfLOaU1EuUHss10xuscCkYnr5Q5pykASZi8hg4YMzAIKeezxEU1bFoi
Zea5mTKE8uDYPjt1y5J6EloZuo+F6fUWkDDtnB+hXvz4x1eHEeXwZgYdlmcmJ7GwB7CzvJqoy2tp
jPFWu7wNrZAR0i6fdJHpIi7p/DL3W5nLHySXSppX7OZnoh54/EdSlktJ2vqhrbM/J1EFaTbJbgEH
aV2AJSHCLgs0P1lHa2uDivH/1UToWvbOnJBiXhFVNzqtL5zuRDyt2KpLFQ8elh8l7rom2xk/oHbA
z9C7rOK5Sv3how7VDZ+l/UofKSKyjuUm4qLgP+Psa4PweUcEDSzBkMNt/Aftp3Vq35ooK5mR4/5K
dybP0oQu7DjBlsxTrZFLjEiUCRJwzKCu0Jb9TWagpVmZGcpO0h3sunPOazKL+HpMU0s1N/oaDjdT
YONsJoBXT8uajlb73SmTvsalPy5VISmM70HyA2yownmI56u4mwrVAHq+MfcpZlSLlLxUml7kNcIO
vwFvDlqtCWzGPmXogfpj01dLTzmATGvkFVjVYQoV1Ux5sAiLXCEDoPTO5FOulFyoPAMrTEEnQCTP
lnupp2uq6DDyNneQkDVMaBrnfgRcjpECT62mJ5kuGTj1H9JOIt/BvZR8kSlGjzoRa7WgHi+JgLqf
oHJCs0RWlNPOw7WNz/HZFmIL6+Q4wpA0HScrZmjRDuvLIhVI5ZUkmhcBszbMLTvGEX9BDfpUCDy4
enqSrK/E/xo33ZLxt/8Etw8Ajg8CskO+9Olxc/e8CPBE5pMQtNM9edLXJ5rYvKmrk2yCeYLW8INH
SE5pruZbJHJY8NZziR/yAshl4ugCx5dbcz+5H8M/7qehEF9qZts8sNvSwLkyTVxfuGRZKazDAPNw
aollmZCcyOPrHfGDsAmePNUXB0gLzxgA2fnvbEzV5XfVgMxf0aT+iu1f65AWrPBTlPljLR0v3AaE
zcgKYD2cPFjSyK/CuzjgsJrMf8+ZBRQ2BDOtWRtAHsH96Lc5RS0QZsNbOqjZmdIjUQ7bP7TZXz5X
qYEZCMHke+Rs+K/wZhNB8gqIO47GwIP2YlXBJQeWpQCnab116ImRGAfPM2Ii94zq+3HApR5gH5w5
3n80ao8GZy0751hQzXFy1ub8Ft+tiABxwuKJ5FbOi8OOwyjUc0L8qVxEDA31aZ8LOag/iUnxnA9D
/Kh/ifraeLZNzFkxR7Pnwr0eUD+/jViVadR4iYGN6YplZDo2iAnkayWxrz3MSi1lQIfTfaNzXwIJ
zz4xZEPNIMG3V28+WBz4NP9Iqb/RsqsnfrTjytnuTVRaHcWANDHA7wla32INPoCnvH4/286HVvYe
Se9p5ocR2qAG9kIkBC8eDHL7B4j1d6cWT6gJsoUaSlB4RXnmwCDUwvWNc05XkXIIgIUHz1a9Sn1i
GBCwkGLHywno6Mx4jD1s9YClMfaySidC7bP1Vlju3/hxOrzzdfogFvvNsxiA3mSoM4RHldBfOBen
a1f4KlcnxWbasTN1G9Tf+aXp0muiKVZZrpaITok0bFREfyRysfJW3ASs61Yye0t916jCjsIDMwlf
HqSRSpvD8H5TPOsEkrNhBBh2tSiHijojHi9WlUe3B9P6lzLsZFvbkg5ZXl/E0hIWnAjtcHcgruL1
hoNIs5IWnaiTw0MzP+Oq10ue1DEa7jQz+l4PXDPECptnaKb+G+Hgx6SYI8ZNqcRdxlNJ3mGYPRHL
ViA5QHims0ipDweqk2cUMTBSCemIGYwsmCOB2iPPaTPn6u0bYYERsqEk/DzWBTVOieQp6NfYfQYE
ali17v+2xCypX6JjdAQ/8TqGSVP+lUlDdreRRO0fYOK6iDdjAgOm3q2GRObhfbpEsin+354j9W40
mZVuWzP1d+47GM6f7WfJzgtEhZnMnzoCnbK7+cBuhlSQBJRXLQlqTZDfpnbqv1xTUWqJGg0UTndO
NuF7jwfzMA3t7LJwd0a3KmLMZRC55QktlcguqyRQxCIA7dxzkuklw3pHLqSOHZCgo2Y+yS7EoE0T
+GgRorQxUEnvZrv8LUODMuo944FIH+rZA7PQxrgIKXPAwkmcd6dRiU2VEMmV/iCOOxUjNVWl1cSd
eW9Pz6MDNdxlQ30KJiIsjRY6Op4b/RqyFFDBiObotvCrr1A081jGFE8/JQ0SOfUrbXzTkzNray7O
YAY8c/I07Jtsz3O/bbPkF3Px/Hj1FVyTn2jTHzaCVQTAS5Zbs5/yKNbsWfZwEYidZ+dRpgdWKwIe
n45VkAYCYzmrjb5sfLH3h+wi0JveHD67Qd5xIcHYLEQmGpszGd9cGVumi7hSkj16Vfh4AYpL7cKJ
YiY3Wb8UBGvlAYc6GxpDDOUKjZ8yUEjHRUjJlG2LGio4Ir7NfvYSJ84kum/g8fzhARerBzJgM02w
YpoYQe5asY0/NhbK+f2+OaXCfN79VnA4ZSHPLAxDDKjbPgpBK9tEaxpOAIy0bhlP4DfiJt90sSwf
XL8Aioqspzix/kTDZzy2CnpoXpQuvF6lzZhv/hGZbw18yke0bw2AEbRpVTMpWvLj/b6NT0I5nxI2
/g09vcpb9e8Ay7niRxOcWdngqpYud5bRGDNOITWz5ttJrtKOd1SMJ0+Ndekm8zEHeGUgVb1Q3dHT
iSEK3xJO/ul04D7L2Zupsr0nskiLc4GZ05jckub0/tljpwXYoGbwIH/h7HRq3cMVlD8TjqZnf59K
IdNfBZUyh1wjtUVpKGAmEK7GCSm7ZMxgejkbhc6yr4bGzZlK4785mkAsWc1QDBrVnc0kw/LFCx5s
/PE1bxrPwtz6QTL/FtFhPZoMso2V9AajRgLsO2QxpaJBAwf2k+OIPXi/BfjmUyPb/9rzWHMC843o
mz+5z6Ij7ZinoyJzUOkK3RMGNisvDsExqVqM/0oSUKk8I+N77CGVKZAODCbQVQklQd6hq0XJkSFh
ztSNe0DYKbaEpzxBfiqk9tcq9wOYcLSYCOIvSBWtzkiC00kotnfi0bcweDx8Udwo7QD1DA2AfD2t
eXz6GFsB0cmYkfnVvikxNGOpj6FLko90qc3DuCLtNdydXQi/GS1vJQ9VN2apf9bX1dkE8Ddersh6
JCEuFOZej6SynAnYMryu0HgyR3X8pB77OJBrTCGkZbzLaMq9vL2KRGQLQS33FliPJ8GrOka+hbFq
tC6FYfLAF7uKGM/S1CQQrR1+VSj6ZvtKfQ8RNOzGXzMwL0bPCcchS2IE2eShD082YtkgXKGEXS5w
zmwY/FW4RjUM0F1gYDPcP7cf2/oUwXyDi/cHguQPi1tyi+Ldpxj5uVvpaAn6UvqWOWOB8orQo0gp
c/SPILt/kh+W+S7hy+UIPRLVLhihtysINabFlDj32ThJFzP1LuDIrBSlhQ6t9+Sca79dj6wD/Lng
QFQfE842tuDbeZAKJ+sBQ+lYKPgPI3PBJy5e5JKMKJeCyHq+JJihu4u2lib9TbV0A2dOVQ8kEiLT
s72ptapn5gbDwQlK/7+EAkc4NMU8lg3R8KL4V8nGyDTXnvksL/44CEpz2K9TZua71VW4YZu8qB63
cIfNTinU5+/L2FN+27QmzKrHSGDVHb7DGnbt0s9LOa7le2/3n931EuTDPavWzktE0t6MNchkLogb
pyftb9x1J1zFijW+Opk6iiEUyMYCJfxbFdLkwpfbKuX3Tr+mlMZisspb9y2jlSN7GdReq0RBpX/M
T6U2s4mL/GBOf46nfJipMRsRYpl2VvekPwyIQhxuY2QVXTmaL5oYA7VTlLNfQ2LbAqLl54hOS552
wzvlC4hfYYMht26PPeI2o9r5j0kjHqIeYswvosUUANLmDszl4+GkC5ePArIvH/1GffMdxawREV01
Yt3R3jY8GE8eyp+xGkC9C55KWhn/gRJ0OJWfeG4MjyxbPKt8JzVwc8xeFlaXBTbSsUqas612f1VJ
CRFqYs4RpE4PubgNCEoh9W4NTwHEWpGf4x01x3LMKWdACOvmBNVyanzcAvpltktKoJT3do6HjZHq
+YgyYws1KPHY5mWQEjSWsxAScHa7foiSQUKpPgH/Tcy5Hgur4DWKlfzfYzc1YHK2zcpqlQsSPIph
IhC/QHPaazH2c2BHBnamUPxlOitYJ0Lh/zcVVr1JTMvxbFjzxrl4S5hA0YpyWJdzsrngFqaJPsGc
SNx3oUqSZvUjSTz6VCGXpkqT9dyWNSzC4L55RtvqHiZ5XSDOAZIgvehU1drmUuXgo0eADDMDNXEQ
f1WkIUyjCWEVWvykzoGoSfHURrBDPY9M8qFghG0RRxwk0AhcbmIhMo4b+Zy5qNmJ/w8sQBHJBC7I
I5x7WK4OssKsYseHQHq592+XOnDoirhdq7D/UfpsrCgokrwtDbe/lzNV6v51QhlLTM6HETblYiF+
RHGVULrlTXnCjSeG6DEwdTE+h5liXzE9KWcdxmUdbRSfJ7Q/ELUwkuFLIkLwLTnQ7CzGmaV8cnDC
eRFHBxYRnVBCaRf3MT+M5niFgSWa90463o56js+Fb1GyIADIoWRmP7qdlV0UzCpT4reG/Dzp9Qez
bGbwyHUvLtDQWMOVK5M5CgrljOBRI7EVLdoFtBiJY08a9QqlS5Z9yzgfoKUex6gLt20ryHboyRjw
obGsyCg4R3yeWxVnYOmSxpOgaXW9ehgsaZ9KjvdXHdfDrK7i9bO2aOFUT+I2z9FUl+7Hr8+Cwogn
g0Sbu8zIHAYGTIG8Leg3wjoWOwPG7suF1EXyaAEYRE44hOXh9iDapOSzMmpavfYGxN14SJ7WOFG3
zyvnPF0FgJYbLvn4vTb5B5Gi9BCmIfU1EgCWQwGUn6khsBoRrfj2Iplj2067EaGC8RC33NSaNzg1
mh14wBn3unmrvdMlACzvg/qzzTxbzWmqppqjLv7K6ScqipICD1IfBifUl7hg1/peLLnDrVU1NxOd
3flBGLi1dh6kdlUanI4cQt+5WR/UtqE00SMVcjSMyF6dMWPg2Oi3VtIdJmmdrmq5z6H6rIm9up5O
vp+Guqm0KKLRXniL7OMMgYscY7W8tXbVFNFYDhc6cgRjQyotZqZU849XeK4ZDaJlSPzIFBuvaJu9
a16FHM0UR1PMYriQP5KeD5CYvwo6117tnAYdvl/NkmZsN6Xo/RO6m3Lqi0o/YZLDbh1mmQO7ajTe
A35M6ZkWaYFKTKHIfsyGgnHWngYcyBcLpt1xvm4c0LDFQNnMVls1qgN5fsngDxKbGcLb6qrNJkyy
1ngYhrc5GHGp4Hd6KvBswcsesL11EWEehvIuKNzQgvK65u/Z9v9FkY5DGmqEByaOlMwJXHoozGVx
1QLNWf5WWTXD6ugb4uQ4UbF1acP2JefGm0RRWKMV04X6NEj1oPI5homGkxxQfA2fmX6CMEatu4hb
t+StSKBGZPSAiBdV5VT/g+5HLSdYHzSZKiLe2Ji2sIbS2MvICxM0ujyx297LKM1lWO2V39AE6rOw
c/BvRlS7cuMfxjfL0CZoXtQKR48hLx/vqFYyzqcYOUcWY+48EYs09d7D3CcgxW8TFou022SQQdEs
9aJYDzImVC4iaOGbU0xTDOhHOWZTncaPPuTdph6Y6+x6rOmvFzBifKyz/rg+qOgOecJm7WQzqrk/
nkIJH4TeXl6hnm1QLwsmuwWKZ1tKzJCob9eiOV/6I5RrfqMSf2gENPp5vwcYPt3c1/KUm5wWOrKL
1W9KD644SWOGOXhPUAQfMUQcJlXTG1CZg5jnNRev0ogQDw9AJUGljIXZZs7XjWyqrjsfePo2fv2c
IyxErWhhu/bf/LBmvg1L0vssmUHcPCsplC3vai5EqBiHyFjTv1HyipOORe5uqlFpvyIHpgHjy+fE
PL7C48NMmkQSNx3YihGZMemY9sFXiiM1WPgwlECjD1imVqW2sxa89iXzK9k7WqZVDHoMx1TCPiFr
QhFiW5t+QOA5eXFAIIGiOt/nZNQOV7aVT5YTnSMHU+l/XIk4ipMSk81f/YAIWVd0J2F+FvoSygSD
eBomZX4LeVmyBFjRlXYoHEEzBexMe/v+aa6uoPY3ot41hFwSL9wk7GujbDW9ThYJxFVp2jml+cJG
e6QaiCFSkqiEjh23acTZBPey1tvc/xEdnfA1aSJhzMPQZjbJeUWlxPNtD3L5ATbdRqdWgEVy/+7m
NERdQExljS3KIfXC4zZmJERiMWQO8znnBAkPopvtAYWatTnmujBY//kGHt8a72+qV4/q4Vr9PgwE
2CF+qcYYwXxpMvlHO/G9KdtZEBvIvNPd7ggr7Kq0Au/ieLplqMJ7+LSPYsRRaGX5uV62DvbGnm79
QfBpX5CGUh5/OBV0hrs/il0uY1X2ky8+ra5gbJ+DButrO9YjufxcpfqLp0x4UNXguhQXyFR+W4yI
l1Vrba8SGNBN3Uo9ndk62cGB3L2BAeBWYCGvgwp9tR3ZTP3WqG48i622d9SCWrk2jzFXXo4CCoeZ
TmP4gvVl0KBPCZmTgqFA+Z+jKjw/uHggcxFPw6txd4STMMf6smlL4WgExPsQ1859BhMhOG47hAQL
ts+mIZSLI8UARwPcM9eDgo+doydPrN1oL06Bzdcwj+vIFCpdNVGGZ8WMMEX1x4M6/l6KjCdv0Sgz
e7dyxPrOd8RTNvWasMW2tfQFLcecNvWHybLk0rCyaC1JlpxsApt09PZ8JubPEwxfl8xybVFo7fvU
LF8iX23zdAYF3cNOF3qr8UaupGsFGUjcIs1aDFwmjk+d1/KGp0u9Zug0QGF3p4zJOPUAPbcTeo+z
//eehhHNg3Q0Qbu99T07XsS21KqV3mrxEFI2jXPgLra9z0fNs3/vmyoQ8cxdilfyo48GMc3uS3WV
BeS/Lefk0krTgZs7JwH/TGXVu0SBYk9htb7xbUQ1zokFs7DFI/5oVChVNcS0C+SWG9S2/piMK0m6
/toGMM4ZTG0PPBPqslr00iodx8fD5eO4DM7an4au883luJi/VbGnpC/iehxSXTx5NdzFq0Rk/ezr
+WdaydS/w1tY9rHyXrJbBriB9mL43pV3Y37GfB4eNKwafqN8k29WWvQs8Vh2yZg26wkM1p5bum3P
xj7N6wPAp/cfhGFC8eo0bMvUmiU+hFxOTjU8qYqW97XD8WjWohWjaowfs436D/pjOcNlhkFAN0X3
8u4Cxl8mAtNnKmIjVoeMBDyyxil96O5CF2OvysMxTUFmMnJvK26/qmM0f7BOPgraohCpC3shFwIA
cS3mMj7vEJWC0mmZYf4KMnKRYbFtZxY8vYAQG2TrFoGYc/0vUtYuswIBrtVn5SHXmgZSZixM4yvJ
FZWrN1ZBxFL4OsA2WSI1K1UOdUAGNPB1zoJz9CBrwEAq2yFhqyTWKlPOleRA0KVNMUdxfwTB5M5T
1kDH6FTJfW7vySJxr5Ot6YA1w3eBX4NURuL9d14Q/WgZM1hmsdMJUvffOMLB6TCR1DOP9Bdjhbwu
EfGW9PQj8j0H+fJVzKp49YMarC/R2YqqoG8ZedS1chbvTXg5YmRsqv/srs967kv7CmZ+QUTcy/Ls
wyHumcUvDAZZ3c6Whh/7Fw1AbpiztmPSqthKaf2HifuyAd/Z23QK46NS23hMzZd5v6IOli/1mJsI
3Fq1+vA7sYoC185s+ncq6vk6QFwB5MYMc/x9ZDijbfnGXP0z/wxje5jYh09dmKQ/tmU2Br6G2aPy
VH16mRsagVQ0LqwRcfQV+gKjVW40wY1Usv/3jtLwwvAtYXM3VqJIgb+cZvO/Ypmu+qLJhpqco4qh
cmcQGgJLaQ/XCExE/s+ZS8aktpqB0rjHXEc0iFEFOSFwR6GE/gHH1ga0mKLWj9oSTuGO4gzaElXV
S6igE2eKiFSX9oiNuIuOUzBClOeV0Xg5nT9KlPYnejNF5n3c1yg3uLNBw6ZBjHugREKxDn9NBd/t
ne9jQKU67n9/RlAn+WcFKN4tdJE9lUPFoDaCvoW9EffbXaAHI9qKL5lkPNo3DN6ENrhyCWAgB475
gUKTCJezg7Lzi+24mSGiZAbkhyXdxZ6W5HfbpZ+KdxlxJxaaonMZ8hc9TqUtXlQFF1BEdzdTV3sd
TNxPiq1we60Iyob4XK/qK0SMqed2dtCfxfTQbirCysjM/NvgmcgkjZG59eEKUYz+kihJx9KkOlNR
X9Qp3eY2jo3r34noPxJmbeI1+gohKrznMepjt58zJkLkcXbrHQ0BjSKs8YKxhpBFSLy2wzpRPPsq
I3PM9DdHOLuA3g/XEaTJDuo4nqzTm2ijX5XY4e519TNroEUU4haX2BEtrJeLX5vwvUXoy/WXYVyJ
QJ5LVYiZLsHR1yMb/H/bp/0Wh3cy9/pwEOy959FnbYvkobgHvzMa20sJeHTrqd4tAuyyRMXUYI0R
EYDFbYnwnUy9/ARXFQpfK0fzYf0rDMfL0u9Pqrypy9otC/Q7zxYw68TQ3JqmMgQ6U5dn2F4mhkr5
H0jjQa8uS/N/SKeXKAbAxuRh7NyiP2sOkMnlBTYA+LIHdOG+6ifKX+hc5cEZlv7zzo4ta/POcfcG
DZFJEVeoJQ35ke/xmgR0zMAkoBAkbjDstMySBckoGA7wfNC+cAcg8+4bhCNFWIN2KCSiwI9hWljH
hc/sYkkq6/u6oT7KV0BMBD4QWWEORq/2Q7uDNFfNa257uXypu2kDi+BT0Y2Hn1W7mtyZXnwxKCtO
jOIUHm3T2lHr/kRYxoO8x116YerCjIVP5crmvUqj9svLSTDXV/KbIjyQ2EGmzbYT4aerq4xYm6bv
5cpBGDn256Ftf8WxxKUO2zjKB2wRzMQoZOMcG7Rb4itLKaBHWMmvcoFQIa7LXmtGV7AfOicKUxx/
tSCIEK5bQTkgS4Pfd/gdWA64EL9qbyHRnTY+8uwiEelBWEOKivNt/Fr6QzJtCpm+dAEBVzE+0IFQ
gXxpLsSblTC0s83LVbNnEbwM0X5I9JLLwPGtwVjXP9XSHZpwp23/MxT08Dgs9Y4ekQxBFoQRonC+
oxq/SvEYQiu8pU8g+vGPukzLWRAcHEJbE8+2Q97asoT1tc6ETqxzfGwLyC4TlCB17ZcGpr6glSzj
j5/DIjv4vzlTn2WrSQH7onoRKBoB4lMyHppD1NKO/VpLReFFZGFArHHtmyUFAIpC+6qoHq62y2Pa
tMbBFZ7RKZ3wNw+RdbLOX0BNwp9jT8v4Z3TdNpLWFBhJA/7q/ODZNJrfvjb35uSHWdg6YmaKWcZv
Y9AFSdwZe46Ic9u+MXXZNBK8UdmPmKizE0EvOoOQq0vctz+nKCxqi1vHKHatuCLsLQYiQjgBfu9s
vXVCcsFBXh0ZgJXFkrScRWBTe+tO2AZ8nO66Yvgt7dFEaf379EsRyvzmZGWr+Q+A19CcbnBN/ODn
tryakhYmGkCBJAoKQadCulO+NDTKD947pnRE9qZveFUpxvy/hNHS8w2YT0nXvEdF5OLG2VuPgGIK
vhIaPlG5bw/ZugmNZdt2aQZ07lV/lx5AZqZWz6r4JjbU8S2VL5Svyr6hW45S2G0uxijyliotMoA0
/9lHfvjYIRVqzkFTi692fUISJ8E1M/02mMfQ9n3rb55O1cuw5eLHa/xmc7q8s6u/SIMgPngooK7/
HbzWjxDE0ELB/A25goN27TJQCs2sXgbmjCTpvnOf0staxUP/Dx385cxTitTne54rxsUsxx66DGpN
n2vZRQjzBtLVOIDgJ0fhPMeRyDJCpC4wrE/Do7Bb5dmEqzGSFoOzzoP+4DHgu4ILWdmda2tPNy3L
n1nrUKDkmoW4h2jP1wgk2Nznavlgnu0e7BXbpsTqxtjII3Gyyif4XB76A4UXcJD6NC1HGtRDmfaT
vuXsFaUirbQKUvnXRb+UsWmCRbak3pBseBSmk/LxaWq7tBK5Hs+LnesIwXDTgPy/dh6bIE2A046I
7QWYPg3r8887ItdU5OPjyudELIArISsr+O/erLqK/0weL/F9TsTmLl0zLqf8LNSmJGVMnLd7Ahad
/PfnnXpuWW0Y2o3/r7WYHxHwAjVU2G+yRLSyyabzmaFT4hHtn8XEbOcBzC1ulSX4jszgG4DGmaAT
qE1G4hQVVQ5I6yRTNEyzdjZu4uF7hlxsj5weKdx3hAetJW+3EiniZlaLflJngexOT4LdUwzTVbco
ZIxPHV5M53M7Pm8VnReejyhzDvOTD01YyUYLWzXqeS/ASFIYuy8eP+wBciWWcaxaNW2qXoxVfw3r
FCDbkbZpx9LGT8zF2TWmUS2GE/Sk1aQPoFc7DGqtKqMlN6h9VMFrzvoHiqMghKr+nffNcFL6kUaM
kC4qFjSNc+N0b+73h1ArQytfhtT4mtLQH01+AokFHN2MssuZyZc4Xunoi59ltmctaubKwrbAk/t9
tebfumXD2YBSOXOH4e4dZem9+sv7TGGNuH/qvrorOTbSbdQcaJCJrtR/6wkyDJUo7K0k2SgjRc4s
u/Bqq8Pe6AvYySBTGsqA4snv9HZThpisL7xR2PMYbbqaJeaO0IwbWHoJX6/oVr3XrW6HNIcglkov
8iYxfAsiT5T4Xx/LLI1p6XhtEUUC5vQcKjsbSuzmmRHEQ3sCFixvHXtsZfbN/EZbkjbRQLGo4Fyt
LfvnJ7JKn8j3UGpJQRVMPc5GughhhzmzbNR/NERP4pdPrRSvdfQvyIhunEwK8fbLNsO8sz+C1SG6
dPlT3f3vxbUrU76wxsUizPsFu+CE5ZUArN3EkMxKwpn4Wi+VnlcUBH3AjedWsqlwzu3HV3y/05Hm
r//6oV2hHwQQrtgNvVukezqo8EiHxj8W74BpWPemsbJltoLQIu01TO1VceOv7KIx8bz0kYlZgBui
KB/rOt6QZGqyu9Gu/Iw3ToqFrU5oOnpL1ljbpcv79w+r6qZXYQOpOd0aWckoxBceYsXD0mGMhTSB
dYC9WsnFEugtHZtaxUWG7NYA4ylZq/uU4vR3nR8tvfC5zktXvLAg4GQqswdtx6qtYr3E5yEYD0LK
0mgmssDAU7DtbAm74Y5tmQhck7gYzXZmQamYANz+/cu2RW3hVx+KTkbg/J0+4LFxGNGTjG/lo8Yq
b3zZtoNdsVTQ2YhnH8Zygs2qY68njNrIld6kCktQkYw+dnt1FwZvdUjCmojND/s5gQ2Hg0v3GWDD
cFseZssZTbiI9xKoupEHQ0GGeLCyEYyD25x70DKWq8nMrhpC5enDmQ+m8sjzMHEpibySfLN2WhDv
1vvBLrAYdPqXxcC/Vv+lqpyzp4AFya51uPXJwOGBuM3OCRZ82OQvIHIEtiPeFEgXEe2WeicqVawm
KG60AZNPHl+oqH+oip5ScFp8s+5+8a0MdCwnwwCO47EziQn2243BMuafwajS+ZIuUcT7sqtfWi+E
PxADCjMFBVS+KMyT8jSj2XClTocEHnHR2NA4tP6S/eQvoRW+E6i9WS/MRJ+0t8udRdi302dah6Xw
2hpHpktj5nMe9KMO3zd7NJLMUSxRq5wZyNVD4DymMvlp+LCmXoawRDh3xR2VBX75RN5peuJgK7vo
VcaJ1v+3B7LmB7DwSP+LhnnvaXHEgy8AEZMSfB/k17UOP7Y45wsXX4AA36PQTIB3glRZRCu3Mmr3
fomFobAdMJ/Nooe5L6rsYJDQYh7P+uSqGaSG6IYAdLSnTjHRMf2IkAMb2GB5o+f/EkIWpAg3xAe0
HVNtLUMg+umpKn+p/kzHMSaSl2HbvV3kYJgMEwbRTfMubLp33ce2ZZzu7pdKqv6pZ0mvyr14/yAr
wrihUF2Nf/9o8dQ0NInmkhrUPWKr6yz5JcI3HteakybHQizcXbqbNiBCWC0SE0Tk6bkdTOE6RGfR
SM/OAu3SvizOrbB5/w7mWAtc+XBTQ0aRvemEYYE5WrOp9M0YMKqjXy1OKRH1h7ncxXU+SZ3KR3Vi
T91j8EdW+Z5v3yLzrRyBlBZ5lxcrn73C2tq0a0y6+z2C4g+mBUIDUQ20eu9q7B9UL7+Zns1rfgP0
HEPTGSaHPOIz1iwbnm8P88rjaShAMaDD0RM9Mytn+SSKHFVt5sn5a9XWPgRWKDtDljbUqgQ7X3JX
UySBk/PBfIzODjEdXirDOnT5LJsXmwThHVBWhetskIgh2cNW1UtRD0igunDbfOTyh822AvQwp26p
eRhLB3lrQvtDJhE0dSH4xDSWs0Pg0/DpHL1RMFN8R0BUWEnJ2TqhyR3pTH4UlpetHD3vhfd0yuFc
i3BI3ULd+4F+A236+1XSLLolLqeHV1QGYdevJNEqFc1o3LtiItGcRMAI8ZT0r05rDGsAMKV2hX6Y
KwzqZI5qjpIBcoP5hBQZf/BLgpUiUW7eTQkVcImfRc9x0z0siEJ/UibrqSz3YfZCDz3LWAZtP95/
r5vHCHeLwTG34oqFzz6ByNYc3+GYouZiJnqhw656s7AcMizY0w9S7fJvjsdvRa1sS/IjDFDnO5l3
eBqjPW/OEYGtBNvERsCEgDPBUkA+SsTungzizuE1znkByVsWAIg8o28z37K/yC17ShGD7r4yk/yo
e+wHMZ2i+Ln8R7uQrU990ZWsDo8yebNRHBQCLQJYE1PCISzXvdW9F1bAGLhNIuJ60rbKDCiBf7VB
muGLSd0PvCPEoAN3XPlo5d+JG8BZpiXA20HTexnqTZhGQzs3B70QBwhZTJQ/sBFfaWnlud5w4okA
MaYxCnNV+ywNmmbKUrC5p+OuOuV/QHYkjuVC7EDWDyhZTmmm08W5xnJluh5Bic/SoHETucbwBBKG
lm2+PiA56G3UKinVBaxE44A7kjZ4PM3ZotlOhuEvrzO0ayaWy/SRGwdmJZpmuHLZk5c3nL37NqWp
ospyT2z8jJVBFqoIaMGWCHG8NAqkxDC5NrPmb7vHqtG60u4xshhpsHxnKF7GCNaIXJWYH4gWZG+J
oylXV7EhoLq6+gl1nL3PEPEZHE0UEXNRoJbrDMuLCz9yCzggTQrEjimnB+VoEQ0fnDfMEHeS/eMF
rlaOvO3qu5X3kQNET1olWnvpxpg8TvetCeh0tylQdaiCaPXe3SC6xTjICo8WMLW5hzztDNZtpDkC
EBucjOlCwhz81HUBNY38s2JTV66XFhVM1AfPG0X6Z3qHXeMUygaby3r85dXBvkkYHhcD32zuKc1w
mnvodHLSSglWb2VOXf/trQXUI5IF+zSlyHlucPTB17cu4Tll93kmOZ4KGhI3woRAlHNL6kxUukxv
sjwRBpg3bZw9JRfJVPv1r/bUy99v8sx5HgMQYKsIBbj5JPV0vKKimtFAiQmWbr4odu0I5+hOl25D
lChFQowyLnhVmR3sKsJl1fdrs+S08lgw4VHKTZHB/3u7pcJ06WAKf+R5YtavdNlWO8Sg/27fFCwp
xc3nkbm2Kl71bXAXHUkobLWVsAMDtS00SSoF44OzBO1c9s78uglZ8mSmjjIhmcihq8F4zwrHFjMq
wXZTpOkQWg6cv6d+jy29jWvAP2cbhLcPTFlT8mGDsgc4RzWEewygoVIozL2k7/t5fq6va+E7y8+B
IBtSByh0xqn2K04wWF461YhVIrFcqHvrDBDU+lTarqb1s1un3uCzjW07Q7Dp+0DHGtXYPBEAVIIg
LFK9RvbxFt/XxtstDVnZYBdOU5OwEI9LSdYTYALltfCgSejCQtDEhJNPrJj0A9Bz3UWwIoW6O5vP
KGYF5ksllKLrT0WbWO+uY7+U0sJhWrbYguQEhj0m49dnkiWw1IWHE5IOcsqDB7RkLegegPSuUZ8D
G8mvsPdHawzJy8O9zacimabuQFedLLMVSJiIo74f9zJ1ih66KGFh8sEw1h9mWh50RQEI2YWUtdU5
Fs+qGtSIcdpuFOQE9RQjMVjFPyLzJdwS4TVfbVGEoDU3rnuWRdSpFyHVdp0L0jDUJpSYLCoYpPml
JFt/mzdQH4xQu4ZxPeUuIsB+PijbfHfxGXUsWEgdQDTs9nuEscneMuS0XaZsu8zf3sA1RN8kYR29
dKT04v9scd9eZOA3enoKLk45jHosV4+rQ2f7j9Rgo/Cff3RsJGtrCdk0RFYkHiljs5UDVCpG5A06
SHYuR+iOgdmNbmHBofHzGR29lU6Shp+nZs17WDNNaAyEGtapRJTGatCCinK1u70T57/Ks/QhCF7b
IlXiVdM25a9gvUDyI4zgkpKrtho1fTOuwrQcnkDd6ZiFU1JNSyNkeK7taeiDyROH2FHX4YsBGtHo
teaJY0qVMYGnqBjrE63cNOClFmhuo9m7kIeJJkGh5IP5xMHBVgUkRNWchw8MCDZyEZDTjnfhdpgV
44ZOovQajsKkd1Sq9M0BEdk2CNt0GIPGk1ytbgqvVMo4vKBz3wGZCWJMhKVOvUoACEph1qxxjS1T
ED6k1F9kM7HeMBW6tt/677VB2IflB/T3aFJQKkKQpwR+gAWhrZDn2g+uryxS0Zmjy5C+Tmc2hgtX
Q1BEh38jCeieD5U6ibC/zAHH7C6xsnYy5LaZZbwzfO5wPiPKXlwQC6e7iENWgLV1t141txsevThQ
XtSItRbkI8J3mx81ap5pol5pMotz3epML/dDwQiKddAOkhBKVT1s9hX64IJ1KSbGtPkdt2RFMsNZ
OB7wAv79dIlWva7FW7tAkli+FKNq9XPqZtFKyRyapKa0EivO3xRlm8CNOQz3OXov6mUu1i/DVo1Y
b55MT/89/4dobA5Iee+Mfo9PgcLsSxaGd3ymOHmCUM3a0NRXPk/CxpJw98eIE5xjUeBJ+wthESzD
PWL+AWw5WD8z1/wvpBdobQWSigeegNiV9Sg2JbdmIMW8xHvdWOz9AiDr6zejgOK4kW4FGg/VIHB6
Dt9AHISY8rY6quc9TMmhfEkVGQDTNncEKvizZ5nQCjE+NaelZnt6c2NkFsa6RJquOGnLx++QQp0S
KhGug7rit3DbePBhEy67afJHgC8Sl7ElhPCYmaGXJUWLX+pg8wXtFgbmlXvZ3+s37oUyp2wgOSXO
hVxCXLyvOYrgfH3uqKvH4cgLlQNg9aryecdPnpMY8BDxRFqmsrWDmcRlTj0vedU5SIpIgbOWA790
Q0fGXEsgd3YLhiD3KKnJ7a9OCUijx24WMhk8PG3CMsEOhPNaN9sJSu2oGv3PMxm8+mkAJl9V1dfX
rSzhCqg9x8JGkzuLsZ0KzKQYMJpgTDL/hjVcQ3N3YFfmEfLX2NJWIxnxENJwYuY6TyqMqJwHDnrJ
FNTs2eKpQVfyRGupWu7/bD2QbdWSLfbXIDynGdufimkFV8cLdYISA8Kssa7ccFaCH96NR6RB0ZHj
y9Ai4AR0Pqg7MDSTe0CrN/3Kk6doVAz1xLQ74icYC2KjItT3ICOvJI5PkrfX6XgayFjSPvuyJ3gQ
5ka0PqoY38TCY9GP6ffUV044q4iJOkpRHxmFX4tL1emLg4hf7oIYaRA0ieIgn5kM5KqtgGRQLeST
E3uBQoec22EXfuNhVUBr+RgiRO2GT/fidI6V4I89H3lHDxgRCYS6uZ+8UPfJGjpS1wus/ADIXuQV
aUV1DGfS7SRe4w3crBwvnPgoRqjSxKkY9fI4nyZFLsCtNeFKifuY3EOkJRzWaPlEDixsIxHTHgwT
P39x6TpnsbmG2jcgjQhvPlW1BxEXkD9TG+4bG8zeB3PpXjBIOw3vrvecAl3ibeuJIQyDZfngh0vx
w+imGuynq7+ihDf9IDR/I0GrjggEuVivMf1KbDqmIoDspTWNxPBbns+tMGg29OZqn0ejUl/w5ymh
CmJP/jTdc9MRq/I9WWX7q7g90+/M2SWPQhrGd4DL7naBp/ZJCJsxoKga7nbT2bA5E5i6A+ZWe/u2
h54LfwqqxSOOBLULKBaJF0mYKEh2Wf0a5tvOQ5AGa6EfgtK9ilNJBWWUgNbGk5mybgky24UpK1IE
9QkFUOh/iX0Zzk694HFwGpqn+9kLcF9HVix30uQmbIHMQcwsKgEuw4hFvFg1vTttijwwkrhzDaZb
3AbGwGjdRFvU3X15Kpj/uteFrNvRVkjvI3jmVIvB6Ee9fQzLYjkmrdaxq4CujWKX85N0ROvxu4AB
s7cvAWaTQeBpqP0koOOG4j4YJf0O8v2PQ26gdzgp/l9vnxBYt0CfoXqz8rJ0w6RrdBKs7JVVnbIG
EjPxMkl7ME00HmF1mWqld9+RhYIjixb+JwF8ZsYgerGir723umSQSwrb2VyAhSTsrGof/hFRHEEA
noQWH84QEq2YPgtvIs9O6foXbiQd7nbiun+d3BVkaEelZrgK0JM75/DIs8nQSk5+7NnbnwTpKbb8
I688TgEq71uVPe2ZbWzrEZjIODHdIQmUCt9+DVlsk/t9HEP5vna9U7FrVIuaby/1aRJGy4liDx63
7rCliJh3YieZvxGwuNpz+BHVe1nmECk+mfGCGXmtct/+9ffeg/EYijinxs2xl9ZP0e8qanPh0Z3d
lCBTVmKeqm+r1ylceBJE28bcPCh9O5SO1NjgOrTvfot3N3V4SJfN0laCWTI/o0N4SG/NglcHFi4b
omj9J2Obhy037J9AsoSRdUt0bOLzuwASxWR7u3exSt9USzKpsiCThkfMiHrukpPj0R7vIgkg/7mC
0w3E9lz+Mdsp+NXfo0EA/9URdCjH3UjbmWaHCJI8Nis1xrm1J9IaGttFXtNya9QiRTedZmISR2MB
+2EAzwIL94MbBv76z7j5Tix/mD//Xd5uWQVPH52ZPltybO2wyGE1RyV42cwF6BMHj688GhmQz5RA
ksWgjs6aVva4muQT7Fdd28qgeI9ITk18bMBkBzmkGdzBRh9Z7ciPfLJpLRO4GZUYutjw/Ky1CEzt
hbAqLoaHmQxz/o1gbpJe+nkyLzwFinQvE0wqwBOK00nr4hNYRrQ6csVKk+TBL2ho9xPpVewtwsvj
NWCNbPgbmV6BdyAetXgGJ0B6Q91E/aARzNBWu/Z/hpS+ZNJAskc0LUOlf804cY9cFV6pSMte8vSr
ZQKNLS4Cxui1O2se/95+QfeR3p95AH5GdQWG5CITL/910JkupiCyNQS4jlzsiumuOHL0lgzAqwJz
0j1yHa8N6wJZ0JRAHTt1iiY52LqtxT7Jl3ZF6GhGJaA6GAXfssy4CaBRIiphVbjj3nDaqNhNW5Dy
UFzLBUu/uq43s94rU+GcDNgh1+YmZAMZmiaVxKmX4f59nfAL4WglvNwaxNNX7EXMXH3nvGBUX+Ul
xYZ2XBfTEVmusRXy+eTVbSgKPpZa24DHoW6syJJq/22kYGHxwtzQuU+t7rvNLLIw9zk9xscSbGUW
r/5CN2YF7pSQA1LFrvdEktzoEe4wPcls8eW8GyWpcxfiBJR/SIiJ3/gBGKGVOL5WvwlRXpD/BbgU
dvVrbbUKhdqNkCIK0p+Mh/gfgOMRhs1Y1cy8tpFqdnWV5pKJXAuZCGzEmvcY4My+a4Dysh+YuBbH
D2CvtkLdwuXFl+Ge6nxdbW7gE+whz4iftNaR1v56XtXD73TIg6FKOYrFhBMTx0cqU1v/3k3KDJYe
Xx+BaZIueeYAEzcag9x4QKwdj5eUv5JPqyPVVMYX1PsodGJY5H8TFrbjdsaY1Bx1L5BwwQ41zpu0
HHGPInUb+YrlDnkQR34KqvfEjq5r+rdzGqjMLxAdhe5UyxQ5/qnRtMZPAT3qWZSyjWx9oCirsgeA
SvwJRRFD2JdG0D6JofaCiFPPNw5ZQNOx3nt1c4ytRUgZmnR8415IC0sgyEN3Aa7yEelR/cK0Maam
87MXxkcrjSCjsvAStm58F2/Pb89buxIiFllitDbz6z5YgnHu3IbovGK6wxQ1sRTWWWD3sv33jmGb
89NKSBF7+527DY3JvS+2ov3PJxrtOJlLxr9ggOD7RUyFDOJQ+8PN0GeITyM0n1SK/cK0ol/SqcM5
4LBbhCxb1qe1VKeCyj/9dQn2pfO93sIObC90bmAdmsTdg3geODYmTybbL6v0LT75ibFS+RJMlT6+
waCM5h1zJxX5gql4ctAlrek8+hi+c/WMmmXNuUAOOkf89TkcI5A8wJa8mgZLetv3MeMb2mbgUnmN
IblHdbYUOINqtl62aiX1QFHM4ZelFxMVIBM77WsgwmVdR7DW2rABa3d414bZl3StROf2Etod3/po
U96GNeOvGsSV4drktNWexQod9uloyEUCa5pmhv8f9w6S4QytMd9T07dwCZsDJHiyIV2F3T0lhxYo
WjpsAJqodMXWMmTe86u0nXg9qw9ru6hrzh3WlHLmcblqkm+ONkEMub66vEw4vuuZJJXWp6pMDc93
byf8xCGkoNPFa22P1852mWeT7ghDhWCaxa5apiQ7j1/6bbeTmJKhE9TdjYaOay5LMdbVOMMO9hwr
SH2iB2Glv28NBOl2hO04LQzwXSfMW4QDoxcEwQmjjFik/LZTh8GBqYRavIkmNQkDJMf1OUHJF26f
6hBcbtVR37ml8ms9QHXMEWp9d1fQA6aI80MITtKDI1TiL4l2HaDjg6qGR0JHSCwQh79DTagcGS3S
/nBJYSULkp1qsoZDf8EdjE5z5Do90l4kYmd+wOmgkhW3xx3AmQMQnw7xAH197riLrgpNGiPhuOVJ
uowNr4CEP7+TK46dJJTOHQHJWyZaAHNg+uDdx/buU1Q5VH/ItAX36n+7mSFIGZNAa1a7NX0MK/9z
PIMvMwAzFm/EDWEAiC3CKcBLDHHMb65yebYa5HORY2eGd5m5EDeyki4t9wLf3jmUEm/jJGGwi53C
uUmTiMIgXte0dAEyeZl1WzKaELrcwgbf0P8npR9pFa2EwZrQ6aR2zCSaWb3is1tKbF6Zyi6nNsnG
TJ7fOF2F2sZ1KpWWDSyalfSCsuB+6mEAhwXGD2LoKBYclGEd0PoR1i4RxITXBizVIiAaU/NBHLdJ
qUIqllQjFFrdNKFKKGBmJXMv8oipJ81ehJzii0WNXTmtSAZTuV2kyTjTUYDO7Z5jowPwiK8CiEsf
lhrx7OPFEe+44xVDoY0m2jLiKrjBUy4ic7RL2wTq98ghjElujM6zZWd7JbOIhwXI4wbQ+x/9qso6
vyFuanbGWOzN+3f7IV4YqJy48wJfxQNYPLGR/TzKX3CAfmaOFeCMGzQkKkN/Kcex8W3P/8MjV8pk
z/K3HikGhwFbKlLEdOQpe0ASX0OJ7T4cBIpJK55S1tD188HvLsbb4z6H14LUrmS92OhxseUj+vG1
DRxnW1HskPwq8XzPehiIY68AIhyzW6oUxspEJU+y/XWhPgVA4mZhcWktEOUA1d9GY1eNP6F2mxkr
XuAsWHCUaq9pcnKXHhggH6W5/aEpAUPrraDqBGhT0DfPg8W1MjK3bQywkm/QHpHMjjmPtLu4h9dk
Da1rRLM7g2WU91i8QJBEtOOgjgBrDhPHFqyoZaD89k7A43UBofPtoo9TICMNtJPkcuCHVB7cTv9M
V24uWPmGpprk2syYMHH2+tOoE0Hsc/bI8hpUMbbdqdz407u+HfwqJziLmyzvvO/PuMRjePSONKhV
Xe38beF/SSA8XIM6kmeTYUv5FceRavyAXocB8aiOPo6Tf0Hk8JfgvfJiZUoM77ytWYr894TJsK14
92xmDdKXZB2VzMv53UPRfGmT5fFz+jmBHkcwZ/o2YrUrH20YeJuBDg4nIB1JH0tDd7IHGIZO+loL
B1kA7iuYu6Ku/xzwOXk12y1HxjUBJI1xiNwzDalv2k5MigFijESqJvV09X6rnw46zQbjqvKQYqER
1W6Hl4wieSS/UqfqOa4e+GD2MMqABA6zKZhOfZoRA9bj0YkPStOTbKUyjfzRyuECbG1X2he/vH6H
W5gxppRdGrUvEpCsxUMKtFoVCZnaBstvvOQYspQHvhBlReXct485IucxG33DiyBKEkwjonIwhk3r
C9Qx6pmAhXw8l6+ROKvXQ0XlZCoJ8Ws5iMKaoH+GYzFh/sJ4Pt3/1HKuKbmYoNHmVXSP47qeDJnP
9y+jS+4oL7XpXJMCoWfSbt6UbodZG654myZtyCjTxn6GopM7t+6FPnS2wcVdu2NBmhGz96Ye4L9C
COYp0uc4dyIbtbr3q+07nebWSBegVco3L6G+sKnzhZvp+7EAySdXpBphKHmCzowKuh0+q6cqTTS4
mTpS+dqgO2ZXe0ZEBa784r/SrrFGoBvhPet82OfiVx7El3r6/Leo7rkP19bHKeFk5aC3AZ1uKbke
KTGfaz8O08Kk+KitIJEF11h5ZIdgoVdkADm/u6OgaoM1NN2l6wvNH2MvXKRMYnJJhc6/yUeH4/Wx
fF/LFY3bMMGwv4Hwadmdq+l5bRU1w+n7qJmURLOfw3EpBNu9ttk4Z8ssfB3ESbDoI62mKN3B2xgt
g/Hxs0B5RMRIoDFu6JZ3DaIXkYWkejbbBc/LJnURbGMoA72D8hGaIT5UTUsyvJbtyDcHg1oQJffS
ZV2vlDqx3f5ZuPc1pBDd54QhpOI7mb34Dor5qGFjPutnxOx+JErG52El1r1nCeo/AGFUyK+jzlIf
56x17utYCFLF2ZG7SsW+IjRKpWJiDtB5yXpMRLg6jBv9AIG4ew044wzym56kBOo3tOuFol22jix6
lEMSUtmcVWPxvjIFLONZN9yJMsJMy5AiGkp1U/gvS2SAObyuQ9XFcjZCmmVPcv9Nz8vc50Ty9TWC
FJ7fovy+NWOZtwGA+soMCsBWWa48Hr+qMhf1yiQ7VGJMsx9JQXiZuS1YP5P+3JbNgWKXbFtlgorH
2GnKPso16b12VUsd7Z7SzSpSxOko+xYA7lehcyOKxmh4sIMHeQkJHi0p7T0oYS4UlQsz1FoCKA+2
WY6CMvo/WIudWw0eUITq/uMb8dm3BG/8HSHDq0lFs/Ef2fLG2KZIvGaCuGHfP0aFn+QtX/RSw39V
Vd2MTOpf7xcTdsSC3hvYmj7m5e23+YVYnwlMaY06M1sXIVci3W3n5Wr1IcE4sF2T+V22XJbrBQw9
SPl+caJTdH2gXC5D+X64K2ooUsq742fP2p6FOwpdFCrqwya0CDA+e4t+nOn2dGWQuE+qPAPQwep4
jQtTC+nDHJgbXTItRQzaKIIyHf1nKvyQJ6TtCMoMf99i2sR+Tqkdd+jpQtTDbpIm/hEjru6mJcb7
2bsmBoCQZxikgrvQTuBLJibMD4bXbSJR9EPh0C+9MUQ1vJTPUhPwLd0YtVir6+R5guF3rqoY4xb6
z/N2OuRP6EuhS3z51G4QKbgUo6t0Q/aSnLaSSOOE86RpXIHLr+yMxqY5WeMN0IUfk0EAj4e6VWMU
hoQHMtJpVaiIFWXbJ1evO35FdmCjWH3XKoiOp2ZDYv1lIPFgdn990YuhMZsAD0ovN/W/oIpEni8F
P3+CKur/X9cbFDS9pyDLbsyaQ3V4dyVNYWK/REN7ZQp0DGbI+HcL3AB8iW0brzaBwASbAj6J2XLE
HDzQQ+go7MMo6IuL/gALa+qapTwnZMg/dQJohA/+xojdqm+JPqRft76vP22hhTtyHtyiHGW3CGco
MMPlE2h6t58iM7HDF3Gr6JVf8Np3eHh4eqOGE/2q8wT80rhqtRIA+ZNAQ606VbWh1nXa7uVywwGw
56CAf10VGHu8x67ENXO4pEN/k1H9t6KmDPH9RxkJAkWXK4drOyh5n7AsfKXfcNvzDOHaxTCOwjyi
o/WfoZKYv8i8vjAWnsdrwwIrH32woWHk9RriBMA7dAzgCV16XDivmhrwwpxdwYdq8o//rHwLNkSd
Gx+5++GJR9fSC/U6BbhuFhAG+Ahy29DNkE8XEOqQXIzMpzSuIIlHOxM926Uate/V1hk12241giQJ
39gXYqhwLLGZvvjQktN9DTla+kmFItF5oFYRNeKb2vxBKvl16jaJYeZWfezsNRghTVmIrRIUVOLL
f9EdhSI2LJuhzf6qoQ0RS+uIUdUXX3KKfr8DGbuwJJgwj7TMHK93ItASXjGmrIUJM8b5wCwnx/VQ
fkLTBB5xt+j1D/7mI9df1lXQunPdbZcbkM49eCoaG/ak24uChCs/0r6NYnhPst1ZOCPgWePZ7h7O
NgeWxF3Z6aXqr4mz7TzJ3pxO7uxmLG+8ewZQ5G3iBXy8VQIxQiMLzqTtt4BkSQ7MLzVfOcltT92U
TwlPzC1eGDleCqWGz6150VdTbuIZTijXjtzJvXlfyLpPqDvb9QFhvIUS5apdk7DxPn5Hvlo1b+LC
uBZMTmCa6ITDx/yTTopIwH+x6qOoxT/G1548fnGA+PJoLwS8yoiymI7UZ8Pf7qsOxTPfSzSJ7g62
FOEqvAC4ykSAtur5OoHrjRBLPvxFb4rPXINB2myRO2Cf+o381Slfp6MdiQAtzsWgl0Xt5RE/+bms
TDmO+SpizmLShFAbpIdpD4G1QQqfWBrcBmUEs26Z/kzxvGV10W40xUp7f4vB/RAf90Erq/UNiG1d
bnEjFM475n284YmJPJC2LW6iTfQqTqcBj9tmMxw7cQPhG+OSSQ6D5GdFDGIbU+M8uxH2A5chT/MI
rcFqLrRKw4mEqbrd8ofcToglYzyADB5HHHvLBSoPNUceCu0ftbNwxGe4c/Ozq35m84f5ofvhh6KR
XmDFebkfA6pkmvOm7uOyRS5EIoe1wRN9OpgPlxTlk2OvJ+JqLmZlvWO0FbHjTjd2k/zY3o2nUB/o
bnCoUNUSoYZF2gGKI1rD2CoZh2fxtgP/iNnNmX+ZDf68Kq/xr5RQHDwKkBQ5ObxIZ47moYrqKCEC
95+mhSiCz/0IlXuFfN2QbmlaqdvbOQkrB3U2q5ncK3CqK0oXaFTYsDZAcH+GQ1kd8awQY0aeCqs4
jqyEDECOcHGnhTqRvv5GI6nOiINB9XvFJq0o8uybMUI/z8aSbLg9HXA3O9/g0bU/Jok2GwqZFe3X
hWDzQWuG/MZoasgFMGlGWnwcIyvJEAuNDPFn3Tl+0cS/nUU46Wknl0Kg1jAQMEjqadLp+eyzTtcz
JJS7NpKZ8RjX87jOf2Ip5UNPMIwQR4r3WyP/n75Z9WPiqUztflHbD0qA+LVtL2x7YN1Td1hMHWNv
2RQ7Pqs5nWyCMbz2Fnu7oQFj66GiqZXMjXfmA3md9XBDw40j7YvBC3q/M1B7qPt36s5qNOhKBkYm
T8sovRWH/cM4lIEHw9W85p6TKZerlEUhxlzNFe8vEKfwdb77rHF+nO/+3jdi4DckCiNoOpn6+th7
kicAiUPGDvs1zpYLt5ut8+y3VyLiTL5fcvUPXsgYxmv9dAaa+F6FJYgpmwUPHTcpL2WR5oGvMFPV
cX3HXT3JEK8ZpSFwglzxN7mjOj1/WoO2QI/AQAj1Hj3iFsCOoe1NWLVqXQthMpnT8mrsuEeZvciX
aR9VCXlQGTqL92E+QK8QwX57I4sPaINpa6CqPjOg4GQruMxtFVAhjlL66jd1EC8qGzq6eJiO6yHU
flbxtI9jbgD0gvBVep5BTdm4cmtAJdAoHTfsEiYQqo4n4NTeIHefQk/ifUHbNQIt8FWS4C7xK6FY
nRPlfOCUllnYTk+oK8jlwW1DYAe4KsB8fmuWrrylbQb6JImL874sBPLh4MuxksLBUhdTiUERu6V7
V2NV1PFhbxXWxfhOalXxCtELLiHDuEMI6ZfcceoLOI+s4S14Csy9oFSf70jIAZuNSA21/EINZkPk
D0aYg97QCGjf/Owbsrd+6qR6SH6+Zqk7lPTd/XU76z2VPCvAvqNa8GdsCeqFi4z6ZHqewng/L7bz
zi4VtzuQ6zhEw02WUF9q0pSu10K14RFvGL6LCG0Nlq5+Z9l9qDRDQsVuFCyZvbosBKFqNRXqVi8c
2FvAF67O0bLpX8BSDWz6GE33ng7YIrkKJDqXDukQax0TphJqQbCdWeVUzhoXk0nlCvLt1Av3gKhG
w9zdzswilYM6GNovYomTfm9AqTZV81UmhuWUSJTGX6fCAi+UbcEXK/bjvBzWnhj3OhJaS+oc4L3U
UDA9g9RhAp+K+mBmWGs4o6IxfTUSGV461UI2yKIorShoMHIPN1SrzeMTcIomUAoYR89ajJWpbXs/
szf/OiiP5WZmKwKRC2DgzpijeFQ+u/4Wg9KmXL3cWHp1W19fyprJoVBCu2k6/ZC6DmuZQTEUSOeX
oY4zw+uKnBEWeKSSORbvUmlqinfKZxliB5Wj03CjTXm8e20VLvtAp3IwbkxlWLYYmivGBbVGu+YS
+72ZCugpxlN2OXzZm3ZViwBI8vSWYiYoZrXGlY49zGncVEouBIyX1wnpIICy3fH4X5OvYu30/mvC
TEOnsgb58fA0Ays5ZEQobmT6v75M7WR517+fPE9+Uf/86NMLfID24f0tQUjLuABzgWoxU1Thc7Ak
XyBj3BskKdOx+Bz6iP0SwNtTPzclFi/Vdok4YyADZzeOunCZZY8tmUSkeZ+pTBGV43X2cuApuvER
CVw6gQacG8Qwdlu/+QV6FthSxlM1mg9YsjdsV0ObSUM2/Na1OjBLQqTunEQoNZvPEOx/eHEVVMIM
/B8r1lrHa99AHDAMPBd/MzLdhpGyOTNnvPhoexCKVnAj7Irag12Qcu0Q3VZ1jmilwNqmgBa6Wlyq
RsjWfo+oHyR3ErYp8zYMYtQJlyedrA/JHaFAxhMjbtz9BxVeMgo4GpAdL14Bp/NX/3pCR4f62sk1
ukT7ZSz58C4f7RG6bHyu8mTVNIu7HUXfsYSizOmQKLkEAGeni4lnBMqwFDon1semLfJdqK6cYBxu
0PZnM//7OSTXzvmDtP14cbsPIi7h2Y/+gBbGOWBz/ZacpqbjZtco43vHhAhnQRNEgf74bykEYOWF
T8qzxvjGQIOOjdCUzyE1F2k3LqyD8E39Mzzu/3j0p9xDWrHgiqRF+fzitG366xYeLWVYjV6dtnC2
20pC6pBv8tnwkILxABSJUqVirVsJs7+Y/7hYdf9oHTSfmFNxaZhv7f25Bw4cY6cIOK7aNxaEINdL
3eCProWoI3GJ/GpkQd6qr7d+s7qEyrLmDWkBqKNRSWST6FlIG4BC/V9rD9b5HG2vzDRHo31Yphwl
sQDa9ZbNUehRc/j+0DcJ+gqgOraZZRR58cFNwR4JVkGSLl1dY3aJUD7dAt2r1yfFUaXSylM9IWK4
73BOskrDZDmXqgrAlSrQdzsOaVap0YFojyT8CU7mClWjY4rTOcbvy0enNApr1q8fTKTZWtYRxoJL
Vh+gabK9QkOtC9KxAP0VVH8ItD5BhN35Ka43t0iSSh3lU2IiUMYdblJ6UT7+Fd/v4REn7FPG7ATC
PvrquW5ePzqHq/MdRiWQM+Y1Or0c24FJCmTfkqNOhgboV3AgUs4dyFgUYTMDRseFa70kf3HePVII
ncoLflHL2Xz4sVj3RZqiSho79oM5n18RNq8sx/gk6gRux5uVcyOJ7yy7WmsagX/+cleZBSOPZeHS
Ezca3bTiya7hyKfn3D8krbngdvB+ibz2qh/iOIA9vzzxFhqh8A/hSix2T2FKqfqlA76rrmTLDl55
SC5YtTesOMAhgqwtgS15GGL1QBrOSIQIbTlc2dB+qZ9ZBVVXNRDegeN9zE8vD5oibt1CDnlzk+VZ
ZNQTSNQVLLaq/3iTTHVzPUYKt+IC/p9n+BfxzRQo5K1n0kjmBiHPVlx24FlrcrLHq30iyP3EFdSI
AoJVGPUWmC/RS/OFLjqXeDbeJX28VKDuOWlNHoph2/BuGgrB+OATGg1ZhzYqX4ET2s4KajUeZ1U7
U3sxylhDAzMEfpwOPIL5h0tj6m6dAFGMa+xYHojb6ldFEFT8lUbIgWzR0mCtP2shIgOusZaBYFg2
Au1dbpRBupmnE+AkCnj7lVC6l0q7I1o70YO1ktmhs2vTyxKNB4JAu9vcsCLv/SbspZLIpa95twtZ
id8SWYhvGjK/HOuAD4qNfPyx2RSOBmQM9NIL8WEQkT4k9d3uwreTlk7peCT4Qu+GGkJ19oZNQ0PK
kpXpi83u0uHn8ys/hiRlFh0582XAgndmwPbiuKITR+uj665JJDmnalD1LVkQiceZj9jY08e0kyui
bXTBa1QBzKgE0jjGr6htd4pw7qwAv+BMZnSJUDmgz8vUaUfLk5JyUNPj84PJtvUpciJyOfP1iFTW
0mSyVyM+lTo8zKMqci+IK4fdjfhS2FxgDlCgQhMe+SS+OaeRcnq1bpPwLXQuaJmRhBRko/TBDjyc
THiDOQq8RuFT09A3QbLfq/a8LZDiBJ4w3P0R2mxuHF0XPCnj1EaACwmobiAhwH3VmAQ5ijM8pk07
0xSBgR1E3N5JGCxVcmWe0z6L0KVXFKdkHya6AZdfxKDSh9FwgnF5Sdh38LyO+TDO3P5AV/wTK6yC
qSJPh9sHPxRHamx6caFvxOJqWCme3mnBjqh5VdHLcojGXrAEdKjfLj7o//Ocpf4VRRnDEIHVjwC2
Hz/mVBsBP86b5G/DRChqjWvatQUXiUjiy1EFk7iqaHciuHTMHOCbOx6wrAjQMVX76355OEOui3Jz
73KifFJcPoiLDJQr6Lb63bSDMiO2jXxQ3F53Nqrmamz9gGcM3KIzG83TcTG4DkathiitcBZ50c+u
AQmoEjQVfTXMjzzdYc8bB9phE29LdbN3oDaDhvULBm64petaznSCJ/i2jWtxVIrGhvwnv5O8UwOf
mpAZqJ3OjvLZGl0VxIsdNEtV/DNrisNJAOj4M/zAuJ8GgOTQqJve138aehiaryxOy/hGIoh6Fu6W
n7ogzfq8GsgU2pcFcCty2vu4Wf1uJ3Nua3i4zq5qjKNksE02+fPh6rFY9RbYGFaNTdtFXbUDhyQe
VIcT+EIfovAcexok6FSTYcMBkU+7f+MNNJm+4bINfMWGi3A6S1DgG3SQz2O1r/maSFEK10RUPK8t
a9KC6scdpLdM0KzRPaV4Cee0rUzyBdKtmJ52UdSYNjmYmXoKlxIRY0nLazqmdFDMxPWMY7LjG5qd
/77qWOa+H7L8IA1wIh+EXsCt34WNb+saW+ub//yoHcjEPAwyo/yr8pdSlW9CD8pMqyClqmEqnrZY
PF60CicsxxpUF/f9H0Co3ytwHAKnYjOAm1DCr7wkpgxdRFWXbU45lJn2V5MciVU/hwnHotm9XVHI
PQ8+XSt8Denx/F6zGzyTZrEf0stfazdnoh2iSe8/lj7l8+Gqz+MQ7IyATTgupZoTANHWcDXUO48R
c/YJWKvrS0pKAZQbpPQsfV1BdtuErzT6XgRIuiSjG9RG4rVa+mWuVtlhkZyPrq5yKx+a4ydb4FhX
7fhO+UGI7BIxYz27jdw0JoLcv3cF7lF/quWbvDaDgfpl1jqHjwFEmv41Cl9ljxER8s3yTwJ6mM+5
gzdP1iIGnSOiQsqIrnaOtc7AeAj6jtjPLMezRsMUhiSzv8YnxO73q/2QIWCqRRNeu6lh95K3Hegh
heddAYdRLUJSqRwpNjmMWmFXrk2UCD0QEJjmrAfketx988LBy1YyfNdXx5xd9DJQYxNDmzPOg7V1
Sp1FEyEs5BqBfzkLqXu2EcrRrFb0oGSO6Xf9CVIGB5TT+xTicf2DwFZfG03smgVfoldAwFVhny3Z
4QFD/ILfrwIzP/M7fQQ6AdYHKUxxFdROoXZpaKEPVT2Qsqt2mx1hgs4kxbNKwCpwbPObo6rxFC7w
cV0B7x4qdEee1KGGROL1awTHja3lSqlXq5E6P2uHqVJYay4tTx5lJTyaq8S2J3SLNh/KX0vZt31P
PZkep61zA3Vm9Eng18ltyKqJbu8oGCh0S4sL5ZXXDE4a0QOUzv2u2b/zCl1f6GO8wLl7BU9KH5my
FWAn6WqJOruMSGFvMjHNec8EjkTjcUSNJEOiKIvf5N7A1VCf2Ua7nKDWRi22vh2fajodvqOIbUV1
LJBDEMYK/uNWWiCYwyW++Vq9PX9MsrmwyU5UIVa1PtYXgJXJMw03+sJmp7DJub9Zz3E5qFcGn4cF
AY0B0CkNok5kPGbrOMTEiDRfAplsefCDmdV5UInCJNzXAatFbc/U0GWT53aO4feDEwys/F6k1tZe
Q0Zq/duGLzQftqJxAMMp6+CgbcOmd1WlXNpuiKpHx2DJiUu0bh0ceYNt6N9a0rdCGMpYh+l5PytH
6fD24bL3cDi9WwyrpNtcHqsiQOc+kk2cY7n5agwWPbjp5GkTWs1O7AwMjzpNqFkfCoVdguQ8cAqd
tn1+0/ohfZH1vn5vK72SPgtt4+eTO/5lGJ6D/S360KUDOk0PjcYVE0TaKgfIb57nyOHyZayGH3A0
qdOOki/kQjOqX9Kwin7i6bWyxOgyhCjKmdrY/l8Swiv7PEToYvJbZF8BQmKnAG6bNMHNUG+mjR4t
GG6J0YaF4IyXCD6cKR65XFk0N4ry+yyMzoZLg8mMDspNhogvk7Pm/h2BW5kmFkWx4Yd5uW4dfQ1f
NlWq3GJTFIYMaol6l9IA/2u4FW/s+KiYeF+z4x1nUSrjoqr0MMmNa4R2OpTsZIdcpoSgy3A4wCu5
w/lsRmqM9kmZQ8z1gPNAQKP26f4M95djZs5U/AEi+IrzgnGTkCNlwmf8kNaR2W1tFmc2XpRMb8kg
6/jZ2zIZp38zO/Ui9WO49a4/1gu3BVeKLyoc4k61G0rb4G0DPmo/K1eZMKnC1bYTg7Ljfs1qAw0g
sCg90qqP86Gm/qdoypdfPaACQignrI187pCqRxpV+mwoJ/4FSiThUCa58qzZ5ls/+soMZgqwPxWL
zFEulcEPsVHG9xU9sNaIPnADHeNqci4k8sEIw2clujffjhHYN/6P/FbIx00rZcbaR+2rG7tgBHPV
YTpWoLqytrYj98QFqzJMafL81sWsVWmxBtObLBx1ehIYwNFOnU0NzOBuL6vcEO0zFLNB5PsUUmTT
AWyAhPA9isvqARcJXH1kCmR+e14BWKCRaF6uhqVYW7fTsotdDPRz/ChC7edcoNDyGp9NAAnLJxDu
baokHw5gpwh/o2yNF26u97mcAxj/eZ/n/jaiXcaNbW7yPVEwCKjcRSb8W4Nb1O5AnJ4y47RuCGdQ
6ZTcfUo3NBYZPgNP6un6N5jYaLCuN4tnqHIqphUp6VsKk0UuyOkaESKlXUF+SlwbwBN7MaiWg0mD
eKnd0FnVNLnhsdApM8u87Okm7M7FNYwMFduT9zajwuhj+ZFolD/2uWWSdK7fNp5MasS2CxBGTTbi
7XVzmda/P/jNYFhl9K9MVXM8DtnOXOZNYL9GNwdsVJXCMtTIcD32DROnWOxyMGeoKjoHQRpCxK5E
SH1TXm/+tlRTk/XGD+TToK8i5K6Y15ysdBOerqSpufGhUUOVjpEHoFea/mQQNjvwmveh/Z2pwMsm
lZ1Kl2TeSzOgLlmYLR5b6EtwH0wLOM6/aEjT/lgTkfft9xc2oBxX8q7rp+DPZD6R++ecbLsO3ciy
alTJlvFZ0gFUpgacl0nHqiM3R7muS1sWAR549fx/CGSelebC8OdOAM9RaJ8la3w0oLVT5dgIaaGC
zN82D1TCK8hkSws3ZJBsHiyx2pmvUoZGGQmnJ7RWp8/JIZEIbAbBNiOMRR4+NUWrghjlTyHpWT3r
rrrOv31qL87qYf8tB/lztBBIgKCqKqGHV2KwCxMgZEq6LT34rhDuRz1AfN4FE8qEBNM5FeU86dNg
k1AMHnxcshIkLh4lX494+yGHneAl/1XRthawLyyaxjcpg8yMI96pr6rHsAt2siDvSG0SodB9uXHd
etgCdRmBpvxc6UqP2nqQo6vvk2Lyam+HacB69YCVAucwxDiDTbhiA2lKib7Io7jbZsOd35alzUi/
QbRPfAgmwgV4EVg+rnovF03QvZWguKBwsV5jGSReXoYgyVZrr6bo+E+frBsowgg8LypHVt9+Fsaw
WU6g9Zm7Sy8hUzq1kPrQ3QBxGuW4sBZutKsNuD86qR4qM9ndo84aZxSkN6gr4956NIHgw9HeyqAt
e4NPGCLuOgF8yTYGci3Cm13mHCAnh3tDweYNsmUV5t3PUWtZUhCk5+SdevEm25IEXy027n8oXeiQ
Tf4Yl+HxilsF7c3kRaj4rhtLPMVWrQ61IWdlfwOWOFDh/N4FE3Ths+hQjSvUMo7Km3FlaJZlyMgH
ecm4qzpzzJBBU38ZXIQMjeNICrG4LyHVEFjKCPpMkwXEyy0fz8WwYl3Y3wAES7Ef6jN1c9pu8xjm
Bl5IY4g7IgYR6KFjxYDDKgs4kxXeSqdQa18Zu0joFsXrc0xYUzCSlkKk9sWjx6RfoQ1xxCqQ4rs0
2+iwlfIt4rxUJ/QeQ9f9Y9lPc1apkNj6mdPDZKpW4w148IDoitPtvpHRq2b+JESc5YSO9mOlQlRm
ttHC9V46cY23bUGBgCdBDr37MhwuOJ7o2wGlX+MXUJ1h3yIeDGTfurkV3ePNGqS3aHcLi3rHFRjy
wcybm+REHyJ0HvzwzSHHDYoUk47VTyHbp+TQuoCPJirQYs+qaWRilAzhDF15QxCS0pZ3IqZIIX1a
qIoGAJA13DCZeIqjrqZC6NXiq/pluPGli6OfeIU9KOjgc/vQ2hrCnIe/OieXXzr34wPbJpc62rxA
P962bCzUWoJCHIu4fSVzBb6kvRagE/p3/W4ByzwFx1Cm14yEC81g4EIQIud9/TI9eNhfdxUOJX1o
cA+UoFRJ7VDzPZOt+UZ/r07rrERmJu2GBp/DKRx/Q7hJwdz7U4Plk+pAgfagERImxz27Gw034D5+
HYuCPbtTSGFrvjqYc2IJZpJaf/8aajTHS2mNgaYTWV7aWFoEXv2HjHCkSo1wfZUoLao7tVYDqG0w
JmczgmTQ0uDKRsRgBU3gInWkGcs3Koa1oT29GaJgH24mzPd3+Bo7WdvwtChCaJ7ASre+bq2/SYmc
jVDs4B8zwPt6FA9thHp2UnHc5nr0o3C+wgxqRoTHdvnTnBrgee27VXoQufSvOeifwYQqS7N8S47X
DjUgzwJWMc4Wo7J4lEajsz6q3xqjQXwKr+ck0Yw2qnAOkxUlnBjw/EllbavgtCD0SCn5Zy6QI1Aw
okSXpHOAAk4aeILBUrhO7FtklKlXhQJGPiE/u3D6IbwZkpVvQrgSSM/FtHUGZGIKbr+/B8jrCaQE
gRsUelNRHQu5p4I3KeC+BWbktQJs140EITgWOc1KhmErkzPZzRRofRPIBaJgv64vwQs5gHzA16X4
BhojtcRB++E+S4xoQhhAukCLdLJqZBKyQ7vs4R1w0/uVQEQ3B+sdXMlGnk/ogk+CaKNTDqb/gPoi
BGfYZfCnQOZH+5ekBAaSUJ+arQjmsTcfY2sSycebTcbL4SpCk8/JNv2Wk6KUzqA7/arqQpzPEWCr
esj+kWm1N4a79HtASi6nREWg1rteuvHDfoxT9mQitOxmAjXd6xr6Dxtt00McUxCGw5XgP11hjlcD
elDRKOG/En7G7/C7fFWCaGsdRPOgrjpZlNrL0eku/dN3o8sMqKtoQvTE9aJPi/hFP1Z8STqanquT
L9yUrlRu/0jh7O0olbH6Q6aKUG5P0jRRlT98xdOWcbjCbAOuSs/eqXEMujjEMnyD1IZiDoxYgPeC
X0Ii+i3zX2jNiTGWgzjO1ACF0F/9/Gdh5AxJ6IOTKDTs+s3LgjstRbEI40qfd7Bcx4mYObNBTlRO
vj77s+NzLt3JIzljqBFaH+lXuZzjBaJAPSAW9UPxZfaK1STk0f/xfnhemUtBNNmYDJE1f4Z5QZ6A
nP2G/qslKw0jB6qJCY9GoePqLB/gLM93XFOTitK3i+2JxiMoQgddeJ5aZomAdhoz1rSRxWoG2DS7
HnM+4evlbqf15LYwn1N0BvAhQXq+C+CgVSPi7bgu8Yz/rFRSYC9tW1xctkbsO9XNtzM1Yw80Q/Mh
xJ7jJPf8g18cqPRudCgv9FxRBH3r7nvFrmuib1m0TU87tqVdrt1KcEyRjlGtUUfzLFturriAVvii
0Nx/D9uwAc9cDUacTcpKl41oQ6XtaCjuO0AhFUXvpkVyMF433NK62l/uisP6tO/pKgvLv6zfVhDk
iNjFFs4gHhozAxCgKV0lKaWCjDPuZMbTnfjpbt1q46F01UcVk2mSnDzVQqptmenFKfJ+wfHqk9vT
MKEiu9KSzwnmBvE21C5J+Gw5k/f3C3ja8KSfsFPzE2YKb0Wu405k8nuvVk1w4K6DIdm93rfZH8j/
WwpExQqOTfcMVKTQcDDnunt8qKAAv79GG4QUCc9t89NeLC0vngNe2KBNadSz2L78xD7aPmLryrhO
SDuyIhjP//mEX2Jh4acvLEOjMETKjoANr0zHh9aey8OkbU5IVnzzkX1ufSq2ZiWlVwuOX9jCNAyP
JyZbXgJzZdFcRFm97sALeVfO7UEGn6WLIhR6kDnSChYSi/d2QGlzZN/oU9BvtPCY3E7nCPmAeV4f
rWuFF8670r12gQP8R0JizYSGzofJu/p6sFLz9fdc4rDa7XYvj+F8nWOC28mkFWg3m4D6jgNQKS+d
hh/xt6czo6ZRwthmD/VjOnim0E8xqNZaVVKvAllbQQyQoJfcufHy2qIZzyiQLo8WD++Bpi5HPZki
nX0jhawSu2gNSGtmeE8Txz/DSK1QoTC/acjWuKxofwmRYMqOsimttWX+PjG2FINu37c+NkpOk2wZ
x733UWHUiniTSvWjy7WAOnZoriWmePCbjbpTWxcKv4efpt7WdBHVsc/E9m4bL3/YjY5lFRY+0fEq
X+I9YouPwb02WcDTtsw8fb0NDF/Phy/AJ86UVmeMhqIRyk+EB7nTMaSKlKElt+B7VVTv8IUBQBOq
37lk8SRbTmfit8YrXsdkqkUhPWJGNgDpvr18h38FCAt07rGcWya499JjO7W9kZU8fFwWeDmF1HUf
+m6brd79PwNteDWqHAcJ1og+E4pi5FrOoJgQaWZn3fWqPySYQxTWfx+trtPADonBsFbQdtCP2gfD
goUljNZuTEjFYzNCLlF6Tcu+UkRtNJbKFDjs7ywrdUdqPRbVb4VkyyNciBMq21K0BxF5oPjroSTR
/IKfwFmKTEgmtmeNszRZR/vsWFuSrBMQQCcengsR7t9Mjacdz9Ete4h/llvl5VwoapqXIOF1/mr7
bE8IdN6NVqLStjxyZ6rRgNEx8uzFZ43KJ6VpfaPl6kDVevpDvldKiYDrjE6jq6Vu3TgXYLjF7WRp
BMjZ+S6KsSAMxU4LjP1TOXp6gvaWQ04S4r9Dp5gFleBOzcnJAHz1zcjs43//2MhDkQ+bc4AijfJk
9YRdbY3nf+SNEeJgXZff5awW7D0dPhCkf72PjTO8Onb8NOsTAREHMscJ+Rr/ffc5Ke0faNe5nFe+
phSqCibkssJenIWsCdg/KdssjmZGZ+gr9XyykLMzD3HtULk5PwdeMjaLd254Ed16ClzY0IahqTHQ
/biVCTSw0HDmlRbSoMUrqTr7QlncJ+GEyFv98XABKVND2tZh5nk7PuCXreEsbCb6oOI63DRrbY5P
MJX8NgpPHfE59947NAC+sHMAddOYdIxHXz4huWLeDzbSTFW3YvCTPUWoPkT1r17spyefp7UiXFTV
+rOzefrYRR2kqxLegKgpthinhLvta4/XdsS4J9vqWSmdrx6xb70lwfNrUEcGyw+5A2xQiMuJdYlI
4IeuUtFnimfzAt10MiQSPC6Ue1Nf7QkDkGgat79IQPzVGshc/F//N1a2osKhmC+zo7hRJJmk9xmF
o27yO3j5J67QDWk3tAOrXglMmlYdgb+j60DIymEO+whblxc71NZxq3JOeerJ2T4Xg/wkraM3X67k
AhdbNuk6Y1cqXW5ymJMkLdSXZCixzVW5nll3EpMseZzaoTLsJu7tRB3/OID7i96unqbDtvqw5Rvn
CRWa9H2Ji1n/Kj3s/TWppPzEuKfW1aqVbC0IZXUnd78MbCDewGLYe0bknsiOPBNWnm/QN4bQpSNJ
0UYywwQ+31eY1Ju3B6D2q9371MqPv+FqFMfuVyMhQ3lHmdsNPH5JC8aSMbQ4EvfOLluM5UBMCRCZ
QktYwF1cS7OFfBrKNRmTmujvpqArSRNTrP3iPfe68sbdxV9s2z4Sa0GXopcU3KoULnxjwZJjCiG0
BTkIvIHcxoEC9KVt3RxjBVgecb8bBB8oCcqZweT1FKRSVQSaR1FdZVFIRGPH51g9+o5umV1BxgpG
kXDMl/kU3tTyiGEhSOz346DZPC9wknvHAqByIFF+hP1/NXGBPlfPvYk9ScLRprqbQ70nuOZ6r8El
hlZxYMVwTSFFXopQa9CecCacVo0x9736VtKnfoedYNqYJQbTTU5yzOEqh7J0Gu732iO8483ixX6z
HXZzgokWgZZMGNkepIZR9RR8aFWb9d0Ig94LX51COg2CUFoZLDeAo1dCk802rWAL3FCz9Flc2Yt1
RxAlOpqmb6a8NJnKPnEUNvHF1RZ0DCOgKmAOlnmZDPlTs+Qaw/cQM4ZjyIPOSvsdYqIcNxaIEKF/
vTQTXfhikuijMJFyKIJAFPYu+uQrlDS+RRLOe6QCV7wXUY13roLggM8jj3J5Sh/56f9iU9SlQNDm
5u8ZZb2hejNlSzVXqc5mZaFDnfb1ing2KolgftD6qrzDq1+2tpwelOe8ys4W6WU9uLbI4uVOrfE4
8gyyViVOTvUEgHabqdgS02VwkbHIiG995Bwg/YIqWhhjXjXk9ZCUMPnii+b7JoOBDlSWRrsAqzJe
7Nh4mY5+Z8kXPhzTF7BzG3Z5oXmZ9DIx6EwLl0MjjgkZQtpcVnDLJ0nymqStiZNoLe+V2mlPDlDS
S+DgDpmfG0V472+e6s/qw6cpALk/VC9ieMsNRUfbHuWUoOnpQQmsASbzEi9lj1B6R3pmi+0JIK0u
6O3/4P14xq67pvfSqK1pDu1PRJOMG6J9gmA0tqqWQIB69xxIVoIdYetZmyhhJ7dwHYJktWeCrdCv
gIpty3JiDQmTyHzi0iQRT0vrupWp2AX3T8eHdVLJbIVglKAu01/eytGelEfUY+Edr0n3mhljyYwy
kcO2T3uf0fKcxRCHhauLXoR1DtvwoGM3kbD+BGfkUR2EMuZF9p01pPf03kg8SxuSAIk1CO2v8pSI
B3z/T7en1IwbsWsiOTF7DbO7tRvk6t1Owy4Vj0EmqkuzwxGsc5h+abtyjY4BjbIkbRvz5OmPX35y
la6l8ktCZsC52CkQ2FkrC8vPOdqvGRlmh4PrbmheWIL4te5b0p14o2VfQOlcNYxIITehc/LHTJx4
7EgwONMdZtkKPSorbQD4PZbbHx488B6sAOomJP+/AWhKfYJ/c7/v7oEGdg3w9MBcjn6mkTKdo7AM
Gm/sBJl46feylEWyFqdfcKkVgTKOEY6cQGSolNYS+/aeeG6o9YInxuruyHgZsQ14VauBVkzSV9Wr
4d41LEVYej3aQb28vf9PZOQFHYZ4QQZWrPDPquU3PJFIWnssHj9beVFY+iN/T1ht0WVcKoBMcrgp
vDPsRWbaUkqmasvvOHmAPpcEfZTvTi8li6awp7gf+WH2WCgZNIcRRPv6PFm/hZcOB7u6Xt9fOcjF
Q97Q7iNsvUWRCrlTAjlE4hcVKKNgsAsI7KiCgZHSW8BCIYnnmK9TSthpoyA4iBAPSij4Qd3jPPqi
IQmscjcqJORQhjy7S04NGJ/y8qDpPfIp2OHBBJtL60+/WRa2XU60lXZFfMLTqczRGVlHd8wb2vvI
TwZH/c/u4MMegHG8lISYYXUec0qVei7FDof98+cPZlizenM04gweDOEKfsFSwA1JvZGRnyp4MFYA
E8bYmaqG/GGCnYR0P+/3w4PQkqhovVcfvxI3MzWuGAIJIqwfxUloBZoL9xWqobw+x7Bq+cjuqBiF
9uHwRVF1zEN+OLN9lwn8HiQYPA8I8/k9nVyQfvbSendQQF7qNMMlp/hdqZ9pV5O70CkpF4P7XqcU
t8gOGKzvJxj58MhmnwocUkXMyJaTgug6BnkPPAvl8dNkP/6Bx0mw6eBQuFtBP4+bUS+Lqy8cyFgz
Mr0yut7jvmzQWXxD/KrC388yyq3a/89fX7KXJttP/b1B4ybj4PqTaLY4e1CyZGmmQvOQI7Q3QzYa
2bR/1XfKcSxLG+enJGfeW4G7rqYmPGjbbKlQwxHntowCpmv1bKGjtb0EuhnrbpAdaTwy5K7VFFfB
jJwfdH9Pvd49fnz/vdD5PcPRNufYAsfjXG/R28TzV3lo4vF5rsaH6Q76/7q8ngyb07qSivCLa3Vi
QlEIUBuwDK01zNhVHZXcRIyMT1/baXQGQzPUaFtGuqiTN6hwHAXmfCwPhERRnO4nxCuw9JjgZTdJ
6th8SnJsW50ajq6NO2UZ7FOjV40cop20QFox0JeHTdWD5L+PWIXhB2wb0y5RDmFAlvek9821OCJz
+i4e4aiNJcKuZ6x5I69KFEUqsmXVzRNJFLQpjOdl44K6xUAvZFMiiJApraUNrofmfCx6kqNFt5zN
s1eHOnzH775qHt364lVShRI2C6KaljTpoqDjDgUoV2HOTS1JXI2m13ZIhbU1eM/5z+RaRX+klSTF
cQVSfiwVmc/EVtFM8gLkGUW8cM+kBsYViz2Zlv/+5+cYyiOB/T5VMWLSI+w8K5osZZK2+3ZfZ/HZ
bv4UuM4Kaif5ogjoQ+xImtpM2BkaujkAIiLlF2DOHHYQZp/kwK6b2pjfYMpvcqdPkVmwcvo/t9Fg
x6poI4yo5y007Gg8eKlzDg87U9MZxQCFFF7opomE57lThBbnm4hkKDoVS39fjVulZp9joTAC98t/
2sLfJP/X7T6HvadnIuJjKChR6+TIBr0647sbaeQc1mBEy6AicbkAo7oEvodRWd14jOdJ2zgpmvt4
czyDH4Q4D0scBYrZvlDcP8oiaTdkeqYUxlk7nyu5SvxgRQYY7JQQtAJ/8Q4WfAh5fqY7aK4RfQlc
x0drSHIcP5PkK2wVLupUfB9bngjAXfwXU0kg5Z5RQdMJkYKN8vZ7WPLjjHTPQ33e5sDiQss2P4wP
R75qMc8WZiV+3mPN1Uwht5vC6ovPwZ3P0AnDP7p04VJ3K9DrrS5Z2cJ5aYBQuvjvYRMdYzs3N/eR
id9MiNIk9ACyO627FH3F5vz75/DYz/nlm7jRVsYEhuV4s9mCIZMEt2WTafJEnKPouMAuBKounJa6
c8bDLkR4a+e+3v1OW8b2mC7gINfy6UcuBg0Kkn0pa76ewESRKxjCQbpxD3+S7YZAmfzkhoz2Z1zF
3S+WDJTBbWdiMFupsKFhCFI7sXQN2Ngvlw4+hpgE0XDWw2xfvTaDbN19nqYaTh6DQkzGNZQY1h08
nAWkn5qJzFQS9GjFjJ+dt68/VX8ph294OZniIVmOMPu7ahcwdb/f2wzql8NEBKiVvrfN60s9Ps+J
nB3tMmw1EZDMne8WB/ksVmu5Ymscpv19fDY2+/20C2eR4wuwUvYJS1j1bIB0jHhF2nT+vOSJtUyU
EpZELNyqq7SPfkVV1BzYSiwA3M9Shgho/v/bxUDXFF7hBK36zHYDUvUqu2FfUnzW9HNKimJyRK3X
7Itv6HKCcdN4YqDcIhV6vYF7iwCFktjE9CzllkpaMTXWArwOfkF1UNr1wpNeqDZuuRFP7g9Eg1xP
/TOMRlo8icbDHLlUBM8qWUCbtSeb/p8cMcwsbhTW3sJMb2wiyuj/V6DAs3WuEIab93kxVdapl3xF
hNZDZG5pcmOOmM3hhi6uIAZGDaoMv8fHvzi76fbS43fcBOvY/JggOs+8t1yo9PUE7QWJG5lTdGey
dhTPdNFY9qAjcFwcoEzYSCAfDd3e0RRLI+NN8Pz8VyJvJvKKrQqEJPEao1pYbC4JF9bxs5Ic5+pa
VgW3jE0d2LRRQrb3b1sd2Ku2UohNOU+INIe5FeYI1EwZZu9b73yXTwHD4D3MxD541G5Am1djU3Nh
GaZ8gjbimUBbGKg6zUBqT7BYi1fTo3M2DxAoSH5+4DER1mUUIT7Ca32uJsozLeuf6PQimTmcqql/
3LC2VPg+4xX1j2hd2UooWrX5tDnWH5PCrCiaepJ8pDM714jvDBhdMLnkl17+fDMw/g0lCwHp9cHO
v7kHgOeG1Hs66sCEFXz1bqn/JUfLMGnpOdfZh0vESI70Fy/X/prsWVv/9mNhADBcaiFAc0KRxPTF
7o2+kV1JCHv1qwsPILDEEjDm0T4SDKP86fiSWtuGF8+14f7R1a/d62Ol4qS+on0aD1ZhM45QeL/K
tSkTKPx2xLQJ2Ptx8TImngzz8QMZXTtO4PLILPQoUURBrVVHaJPl4ccOozjsLK7+DzoNd+iTz29q
8Ov2B8HbZoiYLGNjTzKZd4eiCKDdm4Ml0AOY0yrTYHVjaBcMQplBL2m2B59i23QBAG5ZXkMy96Ed
xr0fx+K5XNjWPz/KMepQ0sVFSx3bhYMfk0J7hLuhuJj4zOe6O/xqQHIuD9oJUT8nQncywDPimNb3
ulEblT7fOAy8Bppvl7NHKZpY5dwAQjYVVZha5zbHHGZvuNaawrg+yWWKVVaAAOlzYJhl7zod2EU5
jATU4h9Y9jrhMx910UKiZAMlaMqj/3X2D+dqriKu7jIw3dRb7ujjk1XSi2pZNX3zIM8kXVKdRq//
2ZSqoSrePIENIghnj4tGcjPF0Nh57NvtV9pC6kulVjjXbVFWKyFssXoiW3BIbBdqeBnVq7aM+Wp9
jXjz/89hlX+r3HKhlsJjPPczE6vU4Pj7Nig70HfsazFItcCZyN572mMASicn4QFnTBft+oJle1CW
791OztNIJU/AvmjRrs3DX8oQhk9MsiPmWVlGD9LfSVCQgvcsFMLshJkbTS2Ou9Pg3ypt4XtRVwXF
F7gHTqGhWwNbV7vuSnNNbAehVwa+tqxaDgSmwS9qiRN7D886ThoWtbN7PQZVljFYbas4NXeGe/A7
NVHVvQn4FRPCJCOd6MO95dJrSbN3fmLfLJfcEglAWVgUd7BWrX7LqZeaFAfH+4FGmuc1960tmmw8
T/dPWNBocUN3v+GTcqcZqNb4nsmTbzexLK/QMP1yamolV543VQJepZzA1JflVGfBNF6PRHjNzuP0
yGzulDPwli2pubsz1B5SrqLMb02etRkQgIJwtrAoa6aBwaRFlOdnrXa8ZKGAXaFM96VylWxoDcUk
j2cmJRR74WDiR0toti9KhE/XqbzZgBDdzy1jyNVD3rmLNVzFIpuyW8XaoQNDYAbpLlBrE9m3yR+d
Z7x4cyEZn7avXQ+Z+pXHDr6gJANnS/B3U9c2dMX+w2T+Ahw4udrypE/FMY87LtFfQrsj+TsTU8Pp
rCBKWdHTcWK8wmz/izfJMDZk7qjnZN07YlnDFzbsGKkDrEWXFyXRJkgWYA/yHanCkz6ZftslvYi5
CxdoXXw6BY8MC428CNKt14UQW3Dk/hBtKY+IV/MFmDn+Z30uH47mMaRxKGmdbBs+HLw3L3ACfrzv
BH+kcMRgFDQP//rbuirrpipifvL1L+ILf1BmBPKeL6VcOTxE6tk0cpzHYOMUzrBN3/lt5yQyJySG
ES0A6eY3EVprEA52dwoghpxezRj0R4xImuH7lqekLRoRGHUVcdgixZI+wXqTSUGYHMAMnkmbbYs1
PvVIUc0sn83Bwf9OVoGlkK65lDIrswvco3bq1kNedYymdwAv6Gk6IPeDUWbm9IlOKOZxB+FNEfo5
R4nDKiVWV8ZlEUaJb4QnA/yFaIktSbjOfbl0pHlQxi0Fsr0QiUa+fA69ovvryTdl5qZdFQSn0O2R
ffy3D7HIRQ3/FFyiGmmHb3cLcEI4fOzA0cGd1EQN4/Kdgq+bPinfV8u3IR4C3lxB9nl8HIsn1F1a
E4YWl2bO2xpaxjJ6QtDswv5g8DfS68wdXHW3RP2PorOXwUSRMZ1kbVRUy1mtiBo5k3lYeFvLvALu
g5ucEYFUjQ4y5SIKRgq/1NURChRmhupN6UlbW9OkIv2FKbZVaz/EhulG+GRMTKOnVWQBsk8Vk98Z
8EkrMkI2KCMnxpVR5Fcs+cJKVCokOj6nSyo+zxqBMM1orYe7WAy5CBA5TnGz5kpQNSRS3hBYnWf7
qj+tBfxnjaZ4jslfF+deNlCRaMPan12WaYd5usniZhJpf78ydPAdeMpL2luUwA8et6Ywlf1QgzZ/
MBQ+WmAJ+HjFfZMj1igTxcMoK3PoQ56mbqsmd8WCrFFNoGh+rF10mWSJ2JBLLinbe1tu90cefu5S
2gDkoIuZpvWhIOY5wXzPaUK+wVU0wlkPiJikCXTR3W/VlgnJJrpJzFq/OPfHWoonztq5mjn+I6ge
uP/UnFzgLCRd7rWi3DNtVNjZY9NQHcVV+apAmCjOMSO8Cz+BskaklGbXcHTIBy1ndW59vRdQ4msa
Jftd56OJCkepTHSy2woD4CfexytSilHp31X+rGqVIHLkSkpaPjh/9v0zJ6vPct5Y2CnYjSzsOAky
9QE16xPkqJ5G2nQBJckjNCeegyZWHD5Nu+ELD8h7AvfBflKm2i6SdglkEl7K8jJnkHysl3vh6vg3
g3+SIyHnOPA4/cGiDCC/okxWnuV+q2/dFLYy/t0S0O5B4DvlkiSENVwWPLf57dspinW+Y8MqUOEx
vTx+dgMUS1v2xt9NbAqvgnWB73xUH8eNtZX/TAeyN9vFBbykJ3Lv6163IzyHcE/8T1jTruIPo0q5
VcFdyqfjji0clrjD1e6p0sqnLsUcJV+XLBYVrqs78bSzgpZPsanD61WQhbzPRoHkWlnWh+RDBxnh
D/MyL9+j1ArtV/iMJXtn7I+eRl1GLvwtmGH/xsyUyVlWsRghgOk62LPGIszKY/ApT3E5A9z8eOk2
Roc8H+z85fQOTSz1YjWnQVsJFYQ0X9jYfgCPIqAcowrvAKeVmYDRPRJDnsPBdHbShPZ5vjt0jwrj
f9w7i6v2hT4xxRo40Mzp75lxHfSwodv/5yQbEhc2a5SW2SDFErTcNc6PVFG5tyWcGiwbyBpJkV2o
P6ig+OgmLTZ89pu9GQZBTyEmnyHjBvTeb/WCL8cwuU99z4Hd6KzOypHzvaHL37/AgJkP/t5O5Kia
eGYZ+j+Rp/08grYZ1u9W7xoLnIbOdc3ITLWXfdnarpMnEMqDu0ut7XYslmjqy3+cuXflx71G9lNt
JgrSKp7wap26o+CoAuG9fon4Odvjvz+jKxVYgWvKvWTDluKm4vDxXphFlfYdw/zui2Vy7NUA1ixi
BlkDn9AGdkK89XyZI4eK2aOMr9QLNiKsckzuIHwPmqnD2ahaBrOLiJCNlzH0x3oARor+gPGn7csR
ECXRGy79afO6Rx0s7LNLy9rdPP4IR2bzIsv/g8HjhhSXmqoJPYEptlW7U80IvHQBW9pho9wIqUxx
E/jn3SX9i2zc1kCj7d5SZ55b7XwGqQiiQoLyJln3qS02+k6ZQ1L2hZ7jgrIajwmQZdPI0elSx/Ql
wt1LF0fghhXmlzoCIVFjNG9g093rLEQ0L0ZFA6ZdYAp6Zah4W0i/hfQdKCmnd0lprmlaLaynLhKh
I3R8Rh0pWP7BNziiVzOOMYr424m4Jl5wYB3cT+hYB1VjtpOgh0CWKJkp8HOxc8sSG9+Xx/kb9YrS
mBDdDPAB7vjCvY65gZGVFX7IdghUQWsTsRO1JOUfDBEeI8eyIKIlmQFBlbEN36Ly3njYrwsbo42g
82hyR9g0s03oC+MqmelqwqVcestUANdDnfKxcIZ+84D0D8+yrE7z7h/2N8ANg0sm7kStp4vmxyZE
ryjXvelOx4bj6QX8HtUfyVS4ulNlpB1NXWGUfGDpz5w/WhaF3CSMJucMzy1Wy/4ZthFeSyYLRZtT
hKrn1pOGcfIjj1NUD7wIACxIHH/6/P7J0zuEczUHaXSRRVoaLaMos1ZfSRgCU2M0TWJrzPRJaQo1
TEgZPbuqgmNZRof+4VtCS6/qjPiLK+Q1CfetnNpx4qFzyvQ7j2iMnB26S0vvnVVNxH+dXIb24L4r
fzpMa3J4e+PySjqWOtHmJ9Tgo5DLrBjiiIWCBLVf/qxxqs6ZWzBswxIP8rXH57bNeVo65cK955q5
gV4S0BlYWcPBopdTezAMqQ4pVuZ2gLAnd7jNYIKO6+ttqa9wi9q1CqH17W3tYsCcaZdTWYJIoeXN
mU4gF+6CqZzEiGH+zgbQ8uexxWS74TTIFuSeBkihmOaH/3Eae/zWNW01IZzxEDbtjS3mSkbwkx8j
jHjUC4hcCfLrkVq/fEkQgYGRw0Q0V7f8i7PBJPoVZZ+xwyVeKg9hQpDTKBPmmjNEZjYsEk7IKcIq
e8FvB1kuIEztgqXfSlR8hZ1ETGOYSaFB802oLdpVOJiSdxWr1zNENeUv4KCdBq6iEoagMyIHLOau
JIpuS2LGgK1MZ+eb6TQ2toBYS/w/n94V7vrpWb9yfxRExmRu57ty90Ry+4X9tKA9uuynVxUKTeq+
Ipt+yIG6uDjUqGX2rMwbcDschGjhwSZu23/MEGFcpvyJbwqcSIfVQowp9VK3HVxnVLXP9CuUM/BT
Ldpuq34EaZ92qfV0zt3DwuJUeCmN/e1MzQEwE6DdLD0ii4f8OZlER/rvaiwT+DYWlJOffHO2OTd0
0oIYOqrj14mDXFFOIkQJLN6eQS8Y6XOyh3ODP6/LTudU+iKDiu/VgbzLU2EE7WDNI0DSKAqitel/
Qhpq1EPvK87cHRpEQ4TLmbxWxGt2eQrDaGXkGXgCQ1IKbAnDGk6X5mpx4hL19jtITnXCFEo1LQA9
RnSSIpwYpPzKWE6n6Y01FfmT/cCoxjsxelbWbsesypspzhlS83IUaGk/UaYvWlygrchqkapGEL14
cp+wbFdn9/lAEQI82rqqM0c29PO9JLHg2G9WgjLI80W8FdIUc4HrMVP2r9NJK/fpKC3/pqaYIpiq
KwQ4NnwEO3v//HnNfas4TfEKERnpksskKLTVSxtEEqZodrLFMzsF7YivKeA/tlCygf7DA9TtmiGl
qbD2gZobWltpnLb1G9WE4jXJ7IDRcN/IcUcMntgtQgqKF/v9n8/w6gV2cEd255xjP8r4a/uIrcZH
7KWqDi9WGLKG5Yo3pYgksjtG0sjXQFPQaNClG2j9iTB7UqOoRVB/koqTTsyGoFz31YASLoq9Gvra
AXuP0xcq0AMB6RdivsFzTLrlPSjvY0WI7juN8J0Tngbe0nZHQdolP/xnszWGD7uDwdeeN+p9U6o4
XGVaRp6Ohml0ghF5WgTlcOMUhJoqAmy7bMn9xaAMnCQ829/rTEYtQIMdEgzifOF7GHdl/nyZYsQg
pTv+87ZjXNxQXzjP6oE6EiBmX41TZ3B/xaBDSVqen+DYrWJeKrSnhm8TpW13bQCIhWtcujWCQIkC
gRZ+6CgqaYUyj5ylG4Q1N9+App/jkQnJ5bEge6xkgY1y2OPzTqFPT+PP1EG1AWuJhKecRyoKsv/x
EYhMqpkwgFAIML1zLpLVi2BcvjSGAg05g4dbWyjkVPqJ2WayNjEPFEGWqLOnpbrNFlHV7i1lz1G4
DitvwZaLtpeIM2kyKCciomdfmJ4HvPusuv21m39QzLtOgTY4YN/ZhQzFNnRydOV1TTazIK8vGpfJ
OEDOWbbZK0wSQYtyJn3l+yqxX49axJEabouMPL/VZ/GALZw6AQLxgZ9zorBPfeaMH0Bff94t6Ep2
Ow4QwOEz7uwF7W/sOdmV45zABA7SOIznxoqCxLYVstuDUR2Wk3Yat62F+DBAdrUkpyB/RxdfHQ4e
+a9PHRbbkW9kdDr+5p5pjhbesNUvWWiVpOl6J0YzmsQQejse4Z7lgQZ1YBzANqaVfx5AmQgXY9C0
4usxJUu36c/XMrYlo2rXmsdhoir1oi2ojVWDl97imbxo1ki2uwLbOplAD8QotLYwfw/WGPFvtwYW
JOB3an0HQg7fvL38rHs6vKsRVi2bW51bdbhXqYHuNJsZgTKuSsCZhmavIYhiO+0qe8g0fFC+1vVS
dedG9zf/8rVfZAUpIUn8XIXmz61U+FmU9PiVr4bUmi2vHPIJFHiY1UyPoOwxBMhQ5xNkWV1Z+zPy
gLlXxpO0Y9pTtA4cmFnrqV1TtxRYnqRoKQGIURpODEVf357NatmMFeqRghANA7gAZ2czInkbRymM
EnN8E3tnOU4zzDj1N6VQsHOlXMQ0jaSP5m23X//DErF26rUeX/5kRnXySYdJAKp5itg8O+TwflSe
cGBEg3zfZ2RZhj9I96knJjS4/4u+yOur779YHZHQltkGFN/LaOif687fppCFbGRBTQubcv47DEk6
uKvjjlXxuN5nnK+W4QaXF3VR65yM94nJxv8rt7Bl29hYh9lfEvxCEZEahYKd1AC45MGBRcoC7znu
0oHuzJt7c1w9FxO65uhZ0MSEd/lxUuO76+KGCYgc6gMtp+YYHQRGGvAT0Aa6HCdm7MTC26OSQkRU
4c0LGQPUZcTcm2UK6+LLOc9TfyhWdzmcZlqHEyC+9TvwnJjDzp87IJxiGm5yrqh/LIQSgz4PRaiY
WlIozEeP/2YlOn6QJXhzqkbEmy6+lDCzl+Fc9dOAmKvquUk5nPa2UeSpJpHBOzaUcobDlCOXiRBr
ybVptVWC8v2b1F5vyDzNvDxQLBs0o0gvSo4zN7PkRgt+CJ7yPsgcN08ssmpllo+m5xqm7ZjkS3EM
l+GTWo5beVkB/LnS60IMxM4HKtWHGX+SFJHHLrW9sQYE5GJdpwLBr2+aCH2kt9zslK61noEMO7UK
u78YboroYjNrVWOderWBE5P4mG53JstL6qYe/PZmocr0jHsEjkdthGiMYOCF+1ox5kcmiedcmJsL
8/+2fu5DVl+gkVcDXtD5Di2Oi3LNPO5zmhK+cWEOaY54UkdZ3WSyTcZU0BCheyeX0/kSuVc2Iiei
tOYmdhmnNqrx24XW6My3GIAsnzNKK2q6di0gjJajodz7n0oP550/H93ctfJw4+GUk1LEigoPrebE
8NPcsE19hqGtZ0ZS7QhGAtTX+ImPYqudEo/HMthfDgUoQ57fmBmUyy847imgCSTYluMC+G/9EB9V
i7h4p4bQwki3ziTjb2/P5ZrpnCMArsk7+4FgplMbi2mP2ajC5H1+qb+vi61gCse3WMoqukvfh7UC
hmCHHUnDj98jKSCyhNHnaz7DPvv806eQzjL1BxJxOdZ3SzsDmlhtk9WFRIsvPp/1BMYIch4C8bMS
DXwToNZJkiNyp6vQIRY8TH7rX6+smDiPpUy0GsKUjTiOo43/KpNLWxrt6voIETMpo1JZxhlHDIiL
28zqFIM+u0q/Kn2ftwCjcgftMJzXEJJY7XR70FUdQi+tCz3Q38V3ad6Rj3SrXatd09i7FOWBmVIj
21jQP8HYN4z2Y7PumaXKyjv/qtjRUp15b9nafczNegUd3kKiW4fvvvULrT9E+rELjCzPeTTN4P+p
/Gk8yGxhjomL+Ft2E2ezksRHC68ugae4LRY9R0bUUo46dRt7QQLilkLTFrSAkSVunJRsO/8asKyl
ATbVMiDQH7GW7JFOKY7URke/LsZts6L+4yp/0SGFakurCr88A7twaeYA53wMapadJ8vT/J6yjVbA
tgcPjakNlCWorLiElSz9SL81FSxnMxkCP550UA/ssRadb28CpHrmSZ+4OafTW4FZZN9xcZ19bifS
RE1tTx1xXy/fys++BfwPE0c271VfwQTbulQna/uVBklKbkSWsmUldOcOZWqvmcQSy/NYlYPnD0Ps
7rS9pajtY0EywfQ07Vmj9h+FFANScOFrmINeRtjCECrfPahg6ABKW1/BHs/JdBSIMtULMq6rpcE+
ESNvfVTuTqZIJdu4qX/lXotXd8EJsoyKqCBQddIpsHJ4OmS9+PoQeaD2cgzH6oxVel17rmBFdKjq
ICyqY3mLB/B0uFs/53kXSLmp5YaE1kh0p2gF0rw1Ko4krRcZQEL7pC7jWv0X2Di1nAyh/06ladYb
EHf2inLfuAF8U09DuJc5ZMjM5z02PGI2QYOslCmQYdaAUNzq4V4oukxSsBPBaaVk31I3A6Co/nSH
brUjyAmjLidGYLReBtun3BlUaqZnWFuxgh4qDit0UqPGyYhPdcy+J0yw7g8aHS5SP0OI84sppSbk
LraiKJPgI5bORGsk0Bc9a6OG/mpwCBp67j/rHqy6vMWkcXY/Kha0He2xTcXCQPfaT6pBS7JQBK+M
hQvfcU0F3Iavb3CHE2KZmq2za3oCHPh/QmsevKo43ZDAbPuq3L9gd3WlmrErDOaL0hm4QYxj/eXg
w+yBaWDhyfAIkOApQwnKnCd401bJWgZbCn9oSzHCxUUKthMC23b9L72FoVXla4VS6tSzYwbhajug
djGcKxeO20lZshC1cRtXR2qd2XqW5OBQbIzAEuqVuu2xl/WyCKPEdDfncURBLL9XfHM5Q9pbFmjp
dZKSTauMFb0Y+gGAM5TzHZErZPo2MmYmorROxw9shjn8A1AyA66GbWrCwDTvMUdsmOS0gwtn1qcw
eGM2aY6f9JCn6cc/RSk+63cgYF05zkmID1TySD2FmRVUCzcmh8+3Zwt3EkSbi0L+NL5TNIm7gBLu
2wV5i0dl0aRNksU4kFtUiaqzI2zhQ9BhyuqTuFFCd4xCMPS2K3OYZcBPsuwDskSey2yfvMB2B0ps
LIfMh3jpGsTdabC4D7q1n5gEIk20jV540ipMRwN/1MfeL96LdWw0HoDSkWJLcF/r0gG+jKIXnBOM
MgD+ULjDtGZErUCMIWP6Q0W/7TFnpI1QTSo9WlqTwDOnWxZrMvv2UuGLczR7eNpMQPb0UZmz6gxR
n4isUkyIuYPdbqNx1xGg0SxG9rQTol8WwQo46+3ygSKWjiZkl/qz/b5ZNS24ruYiipz/nk0RcXjG
C+xkOp9BNX64EJe4XyafHtItTwfBqy27fTBGIH2X634NJODxmduA9bNJu1M+anHz7N641VS/sUuh
DEfhdIuXjl/lAQNtcgDo7iIUzTtZxZCAlfNxLfREba/Hngy++xHe98yRqT96lPzhZ2odJDLXzXzt
+j+QiXPv4EwzdLcNtQ1hSj9L/qS/A+Uk5fxkcI7XtmN+C0IlLH7N4j9e60Ts7mAf/xvQsdUEblCd
123Lgp3l0dLLzSSiGTbwyrTFqvLWO5vxbsw7zq+XTcDGIe7g2upBFtqIJ1DJil21+KklqShcDtk9
aPZnStwaMcWvHJTuRwGe6wuLXmzb4dnqffvd68MrG1HQMZC51S4BrMaEELBz+5F+f/u/v+pVm2i1
HD7X/+SBz2qJ0FzIHecuNHKlJu17ddWzgqRDS69OWfwWSmwArYoGGYGGv2E1TkGDVQnIu6zaaieg
2mmFldML3J1KKiDDB+ulpy3c1iMU8CgWsXqFhTpJiDDCIpwvF/D7GQBIbWv5YC8pTKUruwVxsoBz
UxF/r9Lubp/+3dCU8CGp7Q6ENQbaSBs9i1lBKIgfr82yCs2o49XudTh3s5m7epIX3UiLueIcPzp5
0A57vTkkqDprJoFHZqCYazyu8DoOZGYeGgBype/6yh+R11GtO21uJhwTkabQbq4i86xrJVGaVTPT
HMXYwTeel/2j/RlZddHFzVKtKaAQsUMfOrdLdYsHD/9jb99UAbAp2XyXCzGogDWHirg4WHZ2dZDk
oWXQ1hNoZytt72nnZnD47WQC0n+O3YxDTE9X7CB/xluYPBvuNlq7ahn//BYQ0RqpVXd0j1o8jzQT
G5E673vEkq9pZrkXPVpNw8TCmf8x2bgQ5n+yiQRoIt5GTgfNyGNeZLg0E1ycL+tFy3NNF8bIVH1u
SV5gC0c9O57K2dPU7sA6UMiKDLiwN+VtfBK7aeW4s53Z9IIXQJdxMeVatkn06RDet1imaRIK0Ytt
jH81SvUCyXheEtSOkOzGUyXsqMmbqBYJVoGTHP5E01vKirA3KbRYo/19qp8qMyVbTwBnIB/tUa5i
4q0X1vUcIiQpyBb0kv3JBfsMY7LGjDfHn3Um5w63uGl997pnXYhcG63zveLWW9Ns2bcUNvHB9npk
FuolE6e4d409KErnMZOOKnpxX0pvfVEddZ86pbvuQaJ0mBmOahiREV5bC9mXbDLcNdcQgtCsNIag
VpvZgWpACCjPqk/p4qQOEny9gZgOfn0JNAOnGtBxt8e6HgCiVn4FEYOb/s3q1HxRRXfOUVrVeog0
YEdMbnCg23xoPF0kYKxfFnDtQlalRlRuOUBzw2vFTVBhB/c4UcGmFb4niulegbh9x54Gog6VOb8y
NImLbuGQNeS3HfMN+IzQbwtj6uOZ3meimLfi4O1I1YfcQOxRDTr0rpKz6dJCt+rcLwQzXzNpQiF6
nQ4cT/9Noalh9SSSVLukKShmJDuFwD2JGcabDEizzGDk28gywIWbSMD0P8vxHp1UeVW7Qyn3w/Q7
jb9icj+Fcj4XuWSi2B9Yvy7HuZs0+iyRf4d/RnpHRNSs+mmm6CZXo67+mJYfNBm2e4GhfITahnZt
GRxy/aGtPsAO6YXPB4vwJ4u4sDHQnBZZIl/FLsHoiME6N+bPS6doRZbNgs4rtJS+EGY2Fla9ulir
WJDdODUcsl4/gFErotWMmmC7Il+aCYu1uhZYI6wjjxTbPP8eLumgKzW2JTxuU7JVyE8v/vNprJog
H5QpI3UkyXsjFseq6+fk9b1QXPPXXOcuflN7x70DaNQYf5H2gPWaqfF5LCQBPusdgXWfLeIFGEm6
djBbL9GAHAO8+xlKqwtI+txi1zB57NNwZcg0czeyuMU4lrPd95RZbMcwBJkqwcV/D5i+x8Jcriq0
kA30+4pabmvvWxATa44Se2Uc5qSRlijEOsBdPaSzVU2AUbSS62NmcQhTn7MPNg1BzelN3i/IgCPV
sBKy7M3Dn5Z4/OnJkKImOaeObMq32wYOhrNrDJAJHPREFUA4lO0yQn+sAGjfqQbgdHGgYND5EeCR
0rKwYsrsbr95kP/2pjhSOBXIwFMv8OpGeuUFGLKnbTky/56HFSTaOQdJ1jbS3EA1YIH1/eaJRBIl
Q2yH/jrhtg2aTk72ORYCUR4vgA+u2deQ5TxTqM5tGy9afi2GO6fy41DaMrEVV/YcslshVq2LN4IW
dh7RP9opPs7ecaKQpxmcfdClje4AMD1uYGGxQL9IH8rZOxk7mkCHQaF1CWMPFNyoL3s2Os754JFS
t+pS36mzkEHgXI7k7S69YW2pU5hsyJ0S4+sh1jXMsWjeyTHSAjZ2s1zPh4ar1wxZ2MxM3iIkIvms
Umj/rm4603yHKO3DDxafDNoKwIySd6fRHTYn117zs9U/cjo+Z9K4ua77Tm1BA4eesONhNawYOHiT
A16Y1SA6SXB0BFLQToQyfhJZst2ms2dtqjgTnXuOqqc1vs5iUNLKpDc0ExYRJiuvT9eXO1dU8OZr
rgEdNtOeX7kUZDd5YVp+w3Ifea5Zacue+fLOln2bAmWB1idVUFsKu5n8+K4iGTefO2Bs/GouEayT
+Qash2K30k1Bwo7EDLai1QIsm2TzaQj1lm6AZrqWgOCs3s3r2Nzs3oEucEeVzHHzCZQ9zERT76Aq
Ll5yRxThIb78WUNQgBGAbASrHGGS5iLwxYMn1HQ/sjMgByQ7tCAAg3QRvmMC3ovJSeJ2Yjc01oXR
Jd9Rf3Y+sKkNXhJ4f53wNwG7/OlTmXN6+6u1+WR4z5d60jtlp7Oe4+RbHR2Aa9ySsKxqx16RtrDs
XQNiViCtqTtP62c8qPyhvzTjRDnM0lsA5rGCKpZUAw0wzVzLCzqFHu6y8aVhFMwxQ734SP8AVMr2
Z+Hd2hWX88CNmhTdmfw+ZUJd6IZUbQFKCSfcvx1wMjF2I6l8qhPUBRZwAZS9wj6la7JuTZaNAB/Z
ZP4BqnicK8cCZTmKqe9iSFbko9SCrd0kKca0P/sSgyteF35bQ4QdXB/zP23/jggPDI+DJi1ZMkY2
zO4x5ZPgsC6OgSn/FWZ8iJXM5v8wbjVX338MhJ8ImFFL74N7QnB0jLyb8R87cDvy1WPAnflLh16b
WP0PRrlaPI9NCpv6N4Jdd/PdwtFqqHjeq/jItZJ47RI403ldjr1GJCfEbehckYuDNuD/uWgRv+ZE
t1Pwr5oJAu/FTT9WpJy2sN9BRX+4KrLEu4HwZx9og9l6Tlxlt3HK6N6JchW0qIsryvpIDF3NoSBQ
CmFEmQSahdACmP584iL0L54cy48vTzh9txTHjwNmanXYD82gmMPdDa4oxjHCW516u1IXH8fvlBjM
0VNUrNyLjvhu4sYZsg4pe3JgVzwUG/B4jM1L3NKy6pBbMl1T0CUPpQ79FBfr6rArrNfqwLIwX/qQ
A0SHcP2VjQYb6+jelRr9cuEqbUbWkwuL2u+fv43wH1FQUsOrl8hAgOCXhPtgNH06W2gOyM6wruiv
89khcZpdgNtHaKWccfN72nQr6c1K1ZyEsxNnDBcaPCJQ7fkl94KlmUGjv9Ag4bj5wKYoIqrCbA9U
VmJCsZVJM1RJwIszA2bWM8NAeBlzeY+AoLxj/fSCZw0J7eIU3ntvx/OpyaMqIdua3jo39ibITevY
g1taJw1l9eRO0vvRz2ANd0tnLvhqWg3Wu4gsUnENaE0jD8GJjeRX4fPXqxrNSh/QBFz3v8OA71EH
pE9jx9rDar7ChAZkrT8I+vur+lxbvqgzuV5HCqHLKJ1RJJyo5vbvTYKrW99HLK+yJzEqfUsBAc7R
LBUHRpO4KKHaAjb1qr2p3sM70932LCMEPgmZvrqS2qGVwcMJZo1ecGqW8xTGEbAjT3MrhrgndMai
sygA66PErz7WL/x3ysZO/43VnO7oXnt1RLmntNWXtZEFpi6beS8TlBiLG6LwppdSEtmfeEOAo1h1
LgXqJFExC9nA2MVFPg9f3MfvusK0zxsA4eKvlcPgXMV9zTPveBJRlQt7Q7eM5W5dlVajeRJXU7hC
uPogs+xsC0NqpM/xauOEOXmjqDsdRM8GW4ofR/UkW/hsJq1yz1wsw9UMfcbgKkIXjcqNamEJIHMV
vOnGC3Cwav4/PTaSHnC1KUJvxSnRbOyUpGHv+iyIBJrdWut++YFS2Yqmkl4sLHdI6bsOq+8IyeV/
ZH232VvOUKY8Tt+23fm0BQ4Eaa6Om8fVqAT9Y6Z+uw0g7Cas1oOUchlNbKAoMQdw8vJZN2N/jojJ
Xho2LwXrDviIalT918CD8KbfWDoFbuIU3j2sJJueg5jCA2OqLt7ceWfM/kdWQvx5EmKpliCzMVQU
HY760boiowQGTCnKYVDu21VKD5thcNG/vKYLOXhJ0sszsDzhMl6NFKFjkkfvYHppZjZxmQeP3B2u
4pEOo+jDYisnBqajZeK6S35Cmwk8dIv09AFFIs5MMm39PahIXco45s+4EzAP053eoRTzPUHmdwDH
045zi+SPhaTtaraHGij8cID5kv9PlFnMVDn8eog2mTHrCqJgL3sZAPlwhQUSb5jb5SbK3rsmXkC5
iHU4AXNhO4ZUFGvBnDqNtakJORbP4vQzdWF0g+D5uYOTncoeg8Fx5LzbwQbudhW1Nnk+S0O/UkeO
ge+2nI1iHlGRPjVgBs6EIU5bvJVMmFqulenIa7P3URQYXdCdWluSJJLU3YLuNCYtyseBr7ufJl/G
grjQf5HC4ePClIwz5avQs3kdcErD8MT0hW1BjLL0ZO6is0ShxbTIIzKZJ+dRvCIj/GnfTGEQlxKf
lDjrFBS9EzLkx4oGB6rS0pbepn0gf0Q5ZUj46/JEqj7eGZa4yMqWzxMSTKiFZ2ETZqqJeHKRE5y6
vA8v87tHzbik7EX7rrWnizgjtTsQnOFDVbMNrQJXmtEd63dGjj0pp4xEZgQKCdZlOSvONGUzH3La
AuIUfe/98/c+xCpbjqTok4Pp5a4ouV7GKdV4xLHcukTMksgoCQJWJUQ5u+UCqYnwYPaU+pXACDhd
46bqf6jJslWc6rheEDe8I3arChgisQh8RtA6Twelwoxgnic6gWW/RxuQ/5sUKuwj1RC88HuM8fQJ
qTWVUSnkmf0u35Em6cGX2PKAq/z1dp++QYm02C/oGrxCR0SI14Eec5nUzcR34oNRUD+kKThlFoN9
lNmntVt3p9oZLJG+oh4VAPfle26l/4+WjAGbyZvvo+IRnHoY/lcgCPGdGkHO7sc4D0VsJTLVJlAB
Ov2bHm8Qrhf8lJeD4vmMQR3+NXwwlkpy4t+dD99tSSpaY089tvxyv8ehgau1aMLo6QeX6H8hs5nX
9MVkQeKJw/PnyEl6vptCpJ3/GT21ujjXPbDh8LPrPVaJgCldQOstcVpq+Gy0Rb65JMyN25qjILA9
yxXasE6x2JHRZsyqPcIAUGGCE66zVRtPjR5K6IyNb7CAfQh1QdIkQZRDB5bzAJG09nEkUOk4rWMS
7Z7MK3ufRf4lDjh1abE2l5iXGM/OB9xPUXf+j+uL1YdmQqnusLAkCnvgwdLQqI01MtKL65b4YQlR
ir1YsYzFGdWHuTH51RTe2QD9QT5GFmZeU/nXUEnl8QqNK8TMY+LvvVjbL5WRY0cDg51T8etVufdt
VieRGGkEG2TKNQCBSqgxZ5UBMgQ1tJ8ZBRr9HrcORArJ0Pq+Bj1AYPR/n3EE6Zm9/3N005BvvKIN
mAEdCO8oxJIvUjl+iBQa/Z58AoRe1HfsO0pQTp8QDVxXAQjJrU+qREwh83tfrC1CRnA1bNEABY0A
0kYYfgXdI0wRT04kc3Y4cU63qNBiwcKH4VpY0Ftd335W5ErTBMKW0z3ugVVkF13Ys1D9HzQRptjp
f5388TK4VR7LzQyiPF7Mmk2zBXpSjROzK7v3lLts+8bT0DLtWtTjiuCEBo80RpxDYOjt6lBfExbx
uh/jH7KxkRIehRdqVscx8jEqBy+QNxZ8EBJBuqpiOrYGrpW/ykx4s1Fs67bvL0n+8GofLBBgLEYd
ZmbAm537SJ0aqs38YgA8co13MaAGPnwSiEU7wd513w1slCIccIhh4Nua16WOfPHb0c2YaRQPtCtO
2tqrWFYEn727qcsiYtXfInhOfD56EhXqzstFELhXyBIU8fISWTksQjrwFt/Fh+xy1STbzocBL7bT
X79syf80ZAI/VQt2v2Uw49tJKCEfRrUp/YVV1nRfebHCbUB9RIOr6131YhF99UTE9bIb2jjp0VRG
4oUd49ZQES23eseLAOuTlyr6alThxwfe02v3ufw6C1Qkf27UCsYPeMwTPEhBo9qNzwBlWgO83ksD
SRgc4TMRfrp1Denc2Mvk55Ru05wRXpGxsPWjBR4YtoBX/XXsUBiL1VUDW4JL0aEANUd74/mvAXPH
Wh4QxKroYnJvomFZW7XM9P65VsK3JJmI3Bekdp73y8KzRekJqARJ99Oa9T6X8Zadi6DxgQrZvYJW
RP1tj3ijXNtnOJDR/nQyY/yTMppyrLGeHkO6aPOJLd+8G0F4f4WO+FeAOMdZZm68c0/DKBgNOKbz
4CMwLB1k9vaaLBdEr9dBwmX4a90kDNczW3w7yUZ88JEpvhx8ksRtg/wG7jFc241P/Qii58wpZxo9
2n2qdbHb1G8Mo4sVZBXwZ2YB6rLIwhnHwajSeRCK++qggKnAOlqilFkmxryiItCPZ70pP/yDlrtG
Vho5zt3BWd9GC50lv1mmnEjiGPc+n/MymtFEsTaDHo7kecQT+Az/sOrj9D7AIcG/vWuTvSy+wTEs
iynsmLZypDeBK5sWInw4Bm/E50dmjTxr9osoIKt8v1vefRumbChEbF8EPH8mBBWoXq5qkHhU124q
dCRKr4yZeT3XwKoHnQ+3kS7VtdeWTAkCVL2F9WwwvCFTrlh9kHg0kdMG9J3F4HPMYa1ClOK/FPHp
iPTv5S8lprUAi3gNs/ZWwI2Hd3pyAmSIyVcxEevNDzheJVxjzhwuGirKliDXinSVfzAIrmEzV0tN
Ao/cjfQa9seRd9f6C4hpe+tixBIJVXlkqq+06HZv8A5v4XaWJnx34OM64Pgha5qy14H+1hbNw1I5
yI28or38QQjwwwxYB8zX0b5oe8BNoe+ZaknXVaLHkQ6RyJEyoU7NgkmcszeslyjcytejXNeiNZvK
9C/F6ERfEahwQrNop87Fy6u7BdQ89vffltVP8pCQSko9Icc8JqJPl6kYORdj7/oOqdtKs2dsalx/
kohxtVHJV5GSGfw1EdaU10QtSyITJwvyjxKaQrHcytkuor9zUchR4MnBHdxGeuMd7Bs1hN9K0w+M
q0NHvX1ot0pUwiJD9Gxd2pmslWefioxyIuUjVdTGGL+746rt6U0SrxFR4EcG/F25sb3g+XHspjWz
c5PYWXTi71u35uvMof6TW8P7SQvsQbcazNUt1m8imEM55iC0TF835F6EIt92GjSZ01WVla2jDu6k
a6j4fLe5t28tYEBc/siZIj/52bzU68VvnLw2F8QM9vk/5hHlKdI9MAEuuafTRUPq1NVs625uDKa7
sZG5nIb3Cm8x3o0OWeeX/DRYHvNla5iUl0WnNYXly+M48rro301xaMTMzeXq3bRfWeFSTjp6RWKt
w009uK0otaJ2CSb/XqoYYk4xCkHkC7b1+sNc8Ct3Z5qhmWQy4bKVPSpOXM4FmuYceyObjl1iqvYc
xrRdDBNMEkZb2iYSMHjSPAgwS0HLppAg9l3TfEQTuxvUMAeIobMsqwQ0OZmE1Tqyja4QzOabFOwb
wkhLwziEP5ZP6WlucJFFkBmtUwNzhtoIB3LNi28vp5t32YY3r2VyPsycF6kPxcFR5J8bNyBHtsD9
+H+/PGVtrxjmrY+rEzUSKDUsC2UbR+diPOH5rMSvzoGz3JurE+bV+SIfqUIW297I15sduoHtwMtq
0fGZFnJC/u54CpiwpSbRY6HNcCLbu5+pSMCQsIuMr0YaI1FLbzr+kwW88szeM29q2lWt6rcVa57N
OPRFudlUBbaSMljYcw5O1gCR6Evx76jx7n5BYzF8OK1TXJmndwhf4Y5JVFIqygHgVTdwQ5sOF4Rx
tr5mG0wQRnLbcYalmI2vQ4b1syreZ3HmeHohQ4oSJJsbdY6fNrxqOrLcTMOLEj3Osv2cDSNVKJ+m
c40WPs1xdJbWFGefcTIHUzvw4w9oIQ5gWoHIQTRdzMVBOYd0eno+eBeC3jZE+FN8sncDe6NopTIJ
YA5omD/JGqexxcsKqNwr3tmnuN4tZRTqk/dv0WBMPK2KPQI8O+aVxmFmWVXBbXW5tPvz5kw5QNVF
FHGA4W632MmgzkK6HCenWEIuvFKUUw5mc5rsdgvejIW2M9nxz8nrg6LLEwDjRHeq6sKbVwVIvLzB
Qmitwq5fP07nkqtc1D0RVW55Gmhjq2J7JfYtjiePBp8T5UyMK1eWEuPOrom0ndkc32diNo5hOouT
rOMF0xYBhqNjrVVVqwXJ6Q/aKIg/FMX0+R+j/ZT251968TkHu/tDa/7P/cpGrBCxr/lBOCrr9OAl
XHDDTuj1ax4mIX3YN6uLU+th8Gpkn1YT0NeZGTAOP3CbKxr7OOnf5b1LQ88eJIRhyJW0HcZt9DrO
nx4HREl28zySVs8yVyDbawN6fT9WbjGGfi6h4MBsuohjv0ZLIM13yaaaxOy+io7oj3btUxDbT64L
Pkphs3BYVxN5Qw60C0FiaEHen4eLKcdCSaA51wHLsfx1yBsbYTAQomJUYTJHsbpZfX31U9gFn/78
OcshR6hAzdXM+rIt3Z5X+qcJsLHb09asF78WnxnBawH82GW7AX+DqVzeAmDvV5jIpIG3X6BxfDDQ
WPYXlPupIi/TIzrRcAX+CUbXDHSdtuJkG+LuTPux9EkuZZ3pbOjQ2h2ci2KM/MesK0Ekv8fBzFDN
+nxagyPsruSLVxEfV57XydYU0ZTnbVJKeXemaZfxeE2ke8eveXStGLS7tVKb3XqmNJyuS/Fsw0Nj
9YvK/fPxLU+A+nnrISeFyKcxKZ5fY/+MImtPqlKZ1yfSIicBn6yxxMByhAe0rED3EEuxQ98pSCpM
vAwD9Tlgdk53N04vxBC5r7xfHC5R3F1LHbup9PIPXWQzl3ExRSje7/7DnunRHyhV7qq5mNgdJ5bF
2Wa7nJJnYtCqOgVaFEqIUgr4cECk/otV7e84DQtJHWFJesJnqF/i6R9dqaBgStniAhJf7lf1gOGO
ZgLUYwuPUhshYcEAi3viDYUXECUA9TkRQyrpV7LwErh9F6Pp0ul1xBA2kttzxmelV4t2orD4h7oW
ugovGjtV2Ri/9a+VuYpYe/MqHCOJXcl0ZbCo0eCvT4N83E1NpfeC3uCrYmBiQkjMftOe6aAy1lXQ
P0Oc8SPrLQsxGdLFsBj9xpGlM1R8Kdh12RbGmbTXvoAfv4o3v5fTDalDFFHe0n6JBR/Cy0RpOM+c
MZU4/ssol52Kfxrs4MXnN7VjYgaYBZm4+drQH2XfaMhU2aEJ+rFSc3TM4ja9JqHVk7Hphi+lwQ0b
yEHqVTBDGtarbpctteGWq4ma/dsxvleG16j/N6yav+COkz7RNvM1ABo81iVzIHnv2ER8I1gBAgb6
vFN5+4DbcvCo+Xv4T4xYV9z1RjNL3Ba8TfgVDt2gcbkiGHv/UdWlghROsCMsrzDUY8gWI6lu4sLL
ltLU3Q9kxZwHsHXrarAkZfEk7nmnosY6JG8x++e69R4eWD2gvIxW5vYr0JypMc/Qujf4oRoyBKur
bpwqRFG4iQJBGdbqIHX6zRmL++GnWjXlrvB0IyzRmuivRniAF6L8ZctzIR9RjGGmostTC+kYgLrF
fltiRAAKUyzlFKOnHKlspCYfHhRJ9MLS+Nw6VDEhS4Y0KsW/vnlxcd+4JbYdZ0PMkZAciXualEK4
tLkjbxWodp1ZW1Xc1Jv78rUlXJpgBzvk8QqZHq9T3QN3SfKhu0qIluegYXYtSisrjkbvI9miGF3o
8iByJ9Dp9VF4zMpqibUBsliwcxTk2pmNLB+YVZvYz4P+I3ixU19MxTRdRvrXEsBmX/7+aPBsNRbP
QnNIh/oFTZXk5WdyADGZ4ZN4rWnBNQ3aS8tTRzR6rENiE1dOEYpRYXk02/rpSfT+bU/QcX0cij/Z
FAFnJUkKGcgHVrnUo/RlibM2gRVnSEaV1dZGmf7dbckWwJXqnjmNcoQokPlOnevk4kbzVWHy98w7
HvzgxwzzxgqQVP4r1B45FwqkUeun1/jCrmfCglTSqFMIkZTjTs83eCI0pm/5Wr55uoMi49HZPyQm
+rJyW9nWJQgQEjR1Venq27WubQQ0Xggyz5llFQquDhJCXe+goHOo8QFhec6aN2H8k1hJVJqimOPl
pwHbHwTsogppB9lNjLeMEdDEqeT+f0BOuJskwb5ReFPL6QItjHH2h0pJ8UICRtLKY6A43K+AOgO2
T+kI6HZYUMce4tJsDeRwTM82HhV8s+b38nxjQQXs6t12Y9BmIts63pCQ+R2RKYlhEG/1AHjcwiOv
DIWDcIzoFxk+Tpu1KeZTXjijsa5FwbltX1RVo0YLNX3DmUDSDpbOobxCOSKWJMy+jdtTeUz3FaJH
iKSAVli6Hdg81YaKhZ2FL+m9dLMGgkAbzKq5eog1kHqFpdIxM7OVXqff/A5kbt1IaYSr8IcCmlbi
heopEN/ly8piknShjBIu2YmztlhLWGtFLBMC947tbokb8ILS2oUnTl7u/SN4QDlvxWerSzvfIHi8
NIG9AztBm9rVKufZyGQPHEk3bJEJkYaXUIzZChdkzX7kFmKqo6EPrUp7uDf8eqFXVUAYkrdGTsmu
B8OAAbJ9a+U2pEoRQrOBJQP46eaY2LRwc9vY6M0JxjEkhNAsZl3s7tMl+HEYD2ctORzsqVIeuVYT
UmaABGkrhnlRY+iLlWgzTYpUtnkr6V4UKLT4Nevw22CENBd298Sh7ssPgy5/cN1mCoTB3k8ffYJP
gSaPhBBKfwvLYrxXvxYpU9Nh+adwDshgNVb/1DS9t1MXA17yKLkjZOYV9Sm5tT5/MacYlfmDtXOg
sFfdlUzcFwApqGNHSiScTfPZxHEFWA5GnyZ/kf36kyZeKuiTGtJgDUAXk1ClYjllZhiU/VLJSP1k
qJ1zVTN8kdEZGbqQ0PNKOuiBr/cB8k0ZvizWjJ3yT/PyU7cw3+Af3OEwE2AEKlMELGxU9oZ/Zcri
beiwWcGc0INbX5HVpNPiJMCnHHILvLNERK9z8/Csmjj6FGqleBEF9D3IUMTcX0Fg8cACwYb7liHg
ALkjOhpsmrkBei8UhmTQTAATanolg0cTucIjjst80H5nuj/sBw5SFxevY6+R11UZEmHV19LkSDYy
lnl5sVBVhASpUq1bQiQcbJ/ZKEam78VdSG2+HfZzj0b9lwuGlbXcttamIA5BwINmzV24FPm5GbOT
PfBvpe0hR44JNWOi2CL4J1xUO7RvubFM9OlXIFxyJmh/55jCEoTxu+xe/goxkbP1yXv13sA7GKnt
Mk4etTOi+lPHNAa6myiRw8KzwlYliWHG6MMvREY7gRG9MEwMljlyR9Dt2/LdfxQmWJCZIqu/Gt9l
Xr7+gOm3R3ia00UuX0Jmk0+OOO1WMwXMZ7Kdg5fLQgd03c2dOZkK74lQiNO3I2l4v67ipO6pNIsn
o38tdpBzjtD9cdKDjf/c7TvLNWPGGZMuwrB7z0TU0f0xOYHcoIAWKwx2BZfPHiQ5Oq79cgRXle0v
BYHZvXQtQ0w6HSgVke+iY4YdEiFM2rF0cPVn5q3zepce+FFnoO/yFjfiJY6cTR2LtmQe2EkSE8mA
MBRSnJD+u2rvSBEWkVn+P5JUcvyugnjlk7aM+Rw2VjXMHIUf8ovDaWEoneAXGk5bJmCuDND17s+s
phjO1LmQzP39nSW2aie9Xc6UMciEF/rwJRJLdFpgJuP+hCQCsC5XnTE2psnZgoe2u2mhPQ75TpBV
Ut994Ei5gAgToFYjuJR+4Uw9NYWnOhJt+/VQceagMWVaDE7ymfwEAHIheMbDN3gZXBtOx4/AFBU2
TAU6+yLrAFIH+6HmpiRYR9xanRhdeN60V/UrTaaaH/vdLPdWh641LotHd7YHNtWcfP75LSnkZ1y9
38gxaT3T9MrO8N8KxxJ7iTV8IS91fIQXf5a7TygBdF/5lKqP/1/vK8bJQIQN5uD7kc8HTKAMjRQc
v/3S+nfsPw2gID6gHwHaTSvb6eRaiODHrU9EW8MCfp9KGLqqMqI+JYz0b0zLo5VwkQEJnQPaSMOv
g9h3wAK40zt28KrPECtflxok2lrzjvpPCPZSDXu01FGvkxX1o/VD/A2GODSFS7U+RLxnXcXdfjiF
+P78BhUCsRWeayxdVllwYU+8DvNOecSBv6nWWOpdISwmAvm8vUTdCDXKxBJgBSauC+4LtUre6oMz
BRUeDugCUfsaBeH5FZ1xMnP3cOoXTHqQ4wXYaFE9gtXAoNLEYplNI9dKV4lZGYWo3nSVlBFWjDFf
iPxf0oa5QPbEsNo7P5ldbZ8HuZPYmYWsQhsw+bfr57pxgH4mjowF/BM9pfUgmp4/u6acKCDniTaN
Dj+d8ZT8RXs4yXqNcGOKwBUiDS923JwD7NJpSWwVjqyOQcR+8X1zYFmBMkufIlZR1u4AhHRccl3d
Sp0qu9MxT2RA8ZyUVO9bW/CjY28v7VSBnl+rJkuRomIIedSxaORufHj3/2wupYlGKXrxflUrKfIt
T3yhhfZkzObYxhsAf+OSsrLk6ShiIVE7KRZuun2x6EwsOfRMs1kDhsvfqQ1tB23zfuMwKkU5nDbD
rZjCDYgqV+2e7QU5LNx1CpTYkqqwx3G1wKRZp3/aLmRcFznEhxpU0jejsliLlTF4eYdHX8mRX/tm
8ff3zgShr9XLSxccvsIisXvdyjXqIYbcHzJDymmQLQOXWULoT4BsJyVQJiwWNsP6t5dPQwnHAO1h
E0sGa/xdrQodTrhXPOF2xoG29xYi8BdO3e2qLXMsWgdcjhYuWWVo0OaMn/ri1yA8N7RIWhQFHUZn
GrJyJx6kRLgRHZU3/fbsu4DTLzAtFseHASAMswtYcHocYA+tzBssCiwBbWUD7nENPB9n3gJO8DAL
PXvrRSK9tEFJC6GP5GbNVWFdfFNqjN21+27BSjadcm7y2GXrP660aZiBnD/EmBFQ5Au4mVSBwaVc
izMioAYqd+ZUAGh4AtGuMJfXx4/2xmO0t3J80ixuxQAHZ2lgHJkAI8cc27NWHBXRaVQqilu0+jma
i1FMzCWb0iW3l8pGOSSTRap310pnbExbNtbXkfqmdY3MufD3h28eKqLG8YdQBdFi6zXG0XStH7ey
m38q2P6bxxsuNR1kwks8qVKUdFf0sOCadKZhpMu0Hhg/c0D9AGafqLFRLAVPQAqqcYsRL/N6I4HY
oZ5olrdZz8zWK88bb6YFjxmaBUczRbWKlSi8QaqnG71kXpPZN6+GWoPMlUWqb7ph2f9JNJ6WH0us
pVF83vvyVlkz5QU9ypaBwuyOR2lx+2Tg9g6hoCdmuiDMGZuO4qeVRZ+Cj7BGffUDa1EMPsVpVbgB
hMAmCNjEQwBEXmqnnruo3/VrGiHW56Hs3+KxAxuRkKUj+ttsXAB45UnaocoWe0zrs5Zhb/gfnbG7
9CH+ZTZHqFpdxBk+kp2O5NHs/PQcqR7IrfW3VCqwMb+JIX5VOvGpFZc2VZrFJosKYOCww7ZUQYQw
MW3SvHhv8VMAV/pfyK8QiKZsKbhG+bpgoq2u2wxJi2aA+CW8z7iIL5PkHNMinSesN5JlTgJ5iYqF
ou5q5OGCMJL8shwDaT6C7Il815e+TXxoUyBJYt5MAvWI4ljqi0An/Fku4tEcTC+IC5g/jZii1cuf
JSMJ5eYYVzRmBlfGZ1aOiyr0LRM3tBuRcyk7hySUWxZ/5x64Z8huTo70qx8psPAIm1EOvkMMMeWO
h0NmaihNfwGZXKPX3s8NROFL15FhvczsMn7YwCxaYMd5sNYNBBi2+/5oc1AEGIE+iW/g2L68/agN
mEyCDIrhigrbUMMM7IahAH2+p8PzkH75Ke+B1/fD7SEZFwZhO8OQtkA20vNjwhwhLhh0S0LR9mst
YanKmsV4fMdVpBErvGrCskPhvEaiT/knRtOt9ua3uunzotHkcrTsipc5iOuiQ5/c4HVQCZ0CxMyQ
bgvQ55ar8kERYXUZf4XNxSHdWoJGJvckIHGoGhxaS9UTxsT5OSYNtyXBPkj3dHJ4/FKn6wexmAh7
zXMwppNSOSU5rulWwX3ucaa+OXSLTZ7rwX9W39Tv4aNZZz9ACjHKd8W8NNqc1auBHiaA8L9Fmbam
pypOwHOfDHgtWkoEqDaex7yTwwr4EiJDai4aalEBjr1hi4/NegjLIPHGtC8SIBIaqhEd5+/Jv6rp
6O7Rkbk8teY7BGIjQsFXKCcPEEkLLzepO8xcC2LguoWrsxXMIt8a/Vb7Cg7j5v4FinxsOphXg/13
5mTXnlTH9j/JjDeBNJSAgO/UTHO/6jZ9OqLTfHcqvukLsQWm4ATDA9wgFSEyzZeugiUy0raNz+ch
WrBUiZd1iWIYlPjpRicDrAQtzGSYnrP73dho/MrChQnq57SA4tdxOCPgWVJQshDNRZxxRp/45H9B
+M7YbKd1W5u6Nc35WZXP2MuxmCWJ95xe/pWPs6jXYn3P52a5yrUKpnuGSuonzUdJOBO2tjjkUNj5
8LBWUDU7GUDAPTBfFFOoGE18gVruWGhFv8DOln9R0fHyFaGYcMFWcBomTZinnmITkGyncHEeEFBt
CN+nW8MFtG7YTFphBP544jxc47RyDRmXaB3re0CquYReRTPoakkRFqyhJNH8DtZzExYQVHwC+zwn
a9qBG4hOouWs6eZG+OWGobVU/C1QmTVDVI8CIMr1fHEtyHHfP0eFiiYFvowW1NmCG3xtKXTr3dGq
X6kXr+t8lSyurCC7ovJk49V9wOC0pC5ynJdzk4aUxLGgdIt9mc2Co7M/h32CYT2YmZghcZJby7w8
2PX04byBBMVG68i/mgU2VVReq4wevWTYFHKFwxs35Oi0DUyMRwctPGoWy6vixs4Mpp4r21ENmmDV
JyJt7YO9W0Zlh5G4xQIijsuqBrTZXe4WAKWTpYCQCar6DLhHD613MFmbluTDwjTq09zZxpMU7aH9
plSjeNFrbIzg9r5iudJO78/2esph3vZgCQJHzj6E0pG6/OhoYez0nQahyP0HCYxHXIxbrWwAXRRC
KR89SwvB37er/kfc0mnbV/bEQIyP2oXLaXZ2iI3SQmxjhHmWUgUCDibkmFGdvstQ10Pa2YbQ2qXo
9rr+JcZiiocS3Ts4hRChHLBHzkhDxi7wP0oDUoO1JyN9dW5+MhdGzUMMtuFKb3demUPw6mzMWxz4
Jw0SLv6QkIckI10w25t/omVyQonSCWGe7zyp8NEpN8LlTRCheydZI43DC+n5gUsGGV4iaF5nIHb7
SLV3HhZfg1tixqWm0kiiW3IppENPmnj2UewukHJ6Y9JaBU3nNe4eLQa7nvVohhCTCWPaJ1jvXZtw
R/o8izfhyjSAoWzq4FPZfF+zN95sLUchhK7nQ1aObwfVrgwHiNfGlsLZLUU5EubtGq6dXgNM8rec
fPop9RM9ulwJ/8NBE/OaUiiMAics+eERI7KXCazY0BWjgR4peu6I/tasgsfwpuBblZag/Wem4Tzb
dfNgAFSu7D9Gwa42f2Xc/9y+BQuBdclV6bGY3X7wyJ1BlHycJB6MDkZbXc/s8a6xRJ7KQW3wEi0/
zofVhYMxmLS8y2OWcjj54tZCERmAkSTUUzPs5dOe0gGxjDDZKbzKBucxabtHYz2LfLpm2kNVIxCM
8AiizB371gKGAxXNBLq/6rHUx8ufhKv5tW3KzCdsN0WaS3bhR2wCJWxtOdSajwieGaR8GmeXxhku
JjXPHEAQJDfgRUMv6MDx7ilkHCn9BfkxgDnW55r07P2z4HWxAv/KXpCBHmT4XqsacD7Rx+AOyeg1
fU/QZ442LqhjlxP1d0oFL6Y5vI4gqfGSaCliiRay1ROfTny0lAI3cIhWAJ4C85cVeeQ3LRKNw5lA
Kz2e1LQR6/lniDvthospCzCJLo7uA9qEev5kUOHUywYnSPfsNGc2qRCdSXv0iV0LmZLLaK6Wy7D8
zXa8nh0e02j+Pmc2WKpQJ9u6qwcUcxonwxumkNYoZhtZt596JuS0OuRGWVKhIwuCm9k0CHUsLYRh
Jjyp3aN7aRitEjdl1JGSHXSbVZHyOcEEjbYWJ5ZHGm67uzUQUB2kVQC8KD2fA9YlFiWT6Wr6R9Mq
rTlT4KXZT70OJSvuitst1itWjH0Lm01OGzronWlDFuhA9HUg1Y9Vb1hoNYKZhTL6dSXTv8pYVvbz
CUz5rgCXwLa3TQO6UWyHx/wW3vf1dYU82/HjpVfDvbDsnvHhdkGY3M1Zy33q0iT3jOfKnLVWWKyo
KducT1KFDLtm8mu/shJQNx8np3jKjAhlV6IRT0PTt9OGfjDudZ597saxPjohoiuw5ol4qdeUv9yJ
jFXj7+WEvMk4tK/ZffI7VuDyIB6GR1JFP1CUrCbCMEcuesirSrdpB6aoOVLwQdFhRYuFoC/QnTa2
XdDTblr358ktpY2tooITIWXPKkid10UMk+alyo+bhzDN+Uh49fdDjZ++AcZeUXg+NAvLkb0U0Cri
tyHPgHP7Fbs7kT7GQTTFrxeK5gW8OPyFP+OinucWWeouZLo6vdyksjHbISY8MK7I6pzFgnz8LKKd
bjxo1CkIl/T8Mu7vTO5f1i3S4Hn7l73VJgVbgsY74mpq4hBulY7EP+Whi8hikEfbC/4Psv7KAaC6
BxWZeXatfzKGCtub0O3G8XZia1wuRzziMo4Y2fO7P6QmT6UvqUer2q4YRlTdZu5tVnY22gNJU6/d
jzEJoQNq4so4eqmUmTTBcgRaNlUkDQjFX7+BhblVBvBcRBk7lQgwYdP6M67YLEKjYBXA1yuhw2Fn
l72RxgYJbiInzIm6m0n6AJHqWrXmdaqNaxkWnjS7HtgiIppW9FWHlxN6fIwInfrrgQ5uOZIg3QQz
FEmKxJBazjKv2KiTUi9JALm66aA93spBFBMcJG0Y1+usPVMekbC5llvbmAzbBaign6hsPxSHq0f2
kdMp0qCe2eF/HSquSjYmnZWXvBx0LUBILMwlhIBOQcs0GwC8V6FQI64t1uogxIy9KnkwcEmDaS2s
yotHwkFkeJfTyf970zHlx9XVj9bi8bjXqxt8J8RYW8F8wv/KfWVp9bnuXX5LMa2IofuIgYNfJdXj
LI1Yy0SZUl6yuZetz0/nAz+Zv2yuMQHVcD+OGuKx/HMJVRgwJKKXorHs3BxdinN2ktCdAvPo12A6
HtoVSLTjHTdPYMxcKSANvzasIsjcX74t09tt38/7hClZnOxl1Z3EQKi2KO7omC8K1AIR8wy1HIao
+/Wx38oGNhlHvewXJS5loqku6Q879IDnYjPlRLqe2mk0KCO2JLgH2CPS1+pUdyQrvBjTIgBkc9AF
9nhBCGPgD7YLAx1FJTWs0qMbqIa5sLrwiyXutiwr0FOsg/pLsHfUKTBGvv8igIT7U+dkWVw+i3IP
8r+tr9G7PZulypVleKg5PXG9zBqf5GGQatdJAJ2Po3TKzPMwVcGrp48Gfw9lSzD7EGpqsIwQTba1
i/q6BVIzPTdc4DnpGROEANSML0q/RnWpRcsQiDFXdhq9bJwo4s5MC/JWxwQbjaASdplCVWbwELBe
zfOlobC7iQ2zGGevJezbpWZ1E5zg9x2Ek/7dN3XWbXSM9UDyxFXE2/zK9kGNDh+Oz7qaOcV16nKZ
HfQnx1Cdk4QcSO21jg6c5sujXGrhVzlqfbMIOQd7riKrMcT14caI+9AtuGW93z0CWNtKyQ+StFZu
tNoUtpewunWFi2YQLqQkANXmysAmI2qVZF3vsun7ByZM1TOUkzR0u6mQAU/A6ptC/iZ/tUjYUAan
S87DholotAD0/97FmnNv1YGqu8vUic5Ebpq9FzYLNp5RT/PgNMWhchWTynq02qzEyeHpO/gi5Zxe
WGNzHVdIB+yuJgl2uyOtWxEXCVT90T5Lm78REDLOAQDDTzVXe5Mn3eRO+UODe8sBnJrFOLhwcfF/
meyLQ5x62fZR4QwC9a63kcfsBA+sF6f7JHz6vQReo1rnPYcKIWCtDOS4+AaEZLqLtwfcRFvAkG21
e8dclqBimnyhVPPkHOWmTqhYpOUfPDNk69s3FqxFHbBbFJObc0WAW/I9LSsZ5NixPqH8Uwpf1UCJ
55HeGXY5dUiN+GeJXqFxGBO0fznLZEk0GBrY4Q+xq2cijZ1SHUlNOvYkE3XtDgnYmJCr+g/qvca8
7wZPMvWvKTzQMS9j/eoV3qy+5nrx+BbD1UWrZI/dnrX4nP2sJ5T1Lw+BGyT8hzbsV4DK8WI5gtHB
SXsjpKQH97Nx8PyF1PFJn7dOfHQNTsMXlorHdl/JOnpb4oB87/rK54x2Qp3eqgtPUhNvmTlC5fEk
Ok0UqR7CcyDRs2xXq7awvHu05HwZFXUU1LxMTp4OY5Q2jPPwBKZ5YDHOBBuXMj2y8DcBObhAPVHQ
GxG5/sQoX6s3WziTEuF2Jj3HXOPAw2sEdsG0A4otbxO9DX4CbKpmq2F/ybqfvo5SGuRIUNjo/uMO
bptYOg2OAhG13VbFQvB7e20LV1WuOSZUFp/jwWB+Sz7nMuP3u1M8kl9O/CXQPczBNSrwkfPj0Keo
rE2QlUWZEl39oaRBdjWl+8AOXuewcUBSXXagLsiw+hqpKDEArPmhqliRl5Qfm7wCAMgtOUth+3QA
vjNjtkxK9LKf53+9kg7mAHUevDCVfUlhLGZ88zluC6VPiUwhnWNKrMUwRlcjkVMwHk9d/4VvofzN
bRL2m3G5slRhaUK8ykj5D9zzOfPGS7sd9ya13B7ZUMc96YK+fsQEmrVDlBboKSUO/lzK3vVHDSqR
JuhIzlznNWWrYTAod4Pdjj3tA+7CGU52lLlk5sam62veCNlG8Z1TK2htjjodTbw9E49XA+1/yyb9
2hTRUAj0tCjnfg0k2CMa1ZuFWPqET6DGWDtU4BLLvdoo2EHhJhvnJSXNPOsCYhJlpfuyvBqttxDr
XS0HuS2jFd6gZfIPsUosWAWCK0UnyM2Fbqz3OFVpLAYnWXEdjnAxH21OihHqWBDievKXJTXQLNwF
waKiKHe2fbe2vuTGVE3qz+wtghV5rQ1DZKc0fkHjTKR1LiA6ibP6eZpWSBdIkJNm+CuhwNTXNEzh
LkJXIpQ+jLIm0mt4KYfXNfVv8EdSnFiA4GmRTxWIOx6tp4dCGqKxhxyeyy3Lvs9/zA7M6cZz/rT4
0VlzV7YDyREA/dA/1zSyVM1re3bCLiGH9KxA553zmehBe4aKrNGXhstPbS8Z8kxIofUt8VEAtCnu
w/vBYl+RddszPQNVb2o4HmBsgzG8cLVqVbHn00x3ZYw0MWgQhm2TvDuPJGL6vHAd9z+4FYdpMvPW
dk9rgbKNH/HGd7s5PEqyxx3srTD4j+cQH4KmzjfgCZA1/VQJoK6yMtSfsq+2DhzF6rIl0lfOv0H5
QivcIG+Ggue3chHtbTSSE9d/wMj4qm6swKUlDDTws+iSevphU8YBQLsFejV0QjFpe9VKl8YaELi6
IKrWSjVShJa3/Xnm59UfO+SWJAGwajlAxU1gYDS5UkCk9cmh+w8fWyrVUbq04wne103xDKIvCzvZ
bR113lDdI8YY+WVbPjJouI8zuewc1ef2z9QzaVeOwYYFPnyTpvfca44oVzMGKkrtuviUHyHIDUSK
dySSmXpZqGG4OJroVeeZKjlGr4oz1M8PqesWuM1+NtnBzSqPF/YL/LINJDfvXc1RVM/yP1pnk7IE
yp/tTJyoVAFd0gRk8WQVUKUl3A61I1JABvvC3tjkz31LfyE6qmpo3Eyme0qiBmdsN1DdkgExzR35
1veGB+MSigvUSGq+HIrivTB4Nk7EytaqerZMXxp41+ns6mjwAjf97EypPLNQqgn7YlA5VtIU5lL0
1LX395vH1Vh0O89gitGHFmagMy/f3N3EhdFHRUVPZz9Axbbw4LD9qkKDP2RFMc9KjmIhpby9O1Jn
/KAcI+f1yNw0Bx/VQMCcpM8vpUbh+U06mkmDE/pKJnY7h6gljbuvjUUswf7HRRAH9aTv/fvXU3uF
2pAeJZwHVG8pUc5oJAdsVTxHZhatJajmUvj7W5dAOUnAVgFHg/Gd/nRjSxSsQeeEoA6FIRV9LUPN
II4zUAKDZ4RGvXdyPkS7eRoMHkmTUaMpf0RW3tj5NREd6NC31zuB3WlqORVy8ggZgd0J5GBjD0cF
uXTi1z0tOWF8DRCp47BvIAHYwO1J3Y9rrurVhvyeP+/BPmo8wkLoPezDeUsqIGmphg5oqtSNcFud
kq/xnb5/3khPkmnhDiyUrSzj5o7EyS8MANvdnu42K/OZslI4BrvnLeR3gMIwyII615LpeBNi/WxG
lKrWU57ooBqluOuNuDqothTUe7mJGU0A6TJpeN82A8FwdNTl15EtJKGP5GU4uiEoncFaPIu3/074
BXJnN1CDlKB6llvKbHZxtwL2t5DsCe1kcrjV8vuwSIPlVt4Q0kEWU5rAhfEYxpFG5Qhqwo9+FpAs
kiI/Oo02mFTWXbuZaLFELe4c4YQ1OmwG+9BSeYzKdOQLB0XVEm+dhJVi9nL4gskpsmhu2ua4I0/v
ePpFABpsi5703WI2zvMN5ciWwOnh+e9ibHcTQpmcVrBF9EBE3LJ6DPICKfgNrHwh52saEN9zkISX
Ad9ZeowkWSSZeE4EhorREL84AUk8861xShm4+wVf7UIY3euRtbbbSDy3YHDG14qnXB4y3u6yudax
01/CMJCiM8jIybzJWv8urPQSWB+rGPmLj0KFqvxX4G2hO3hzt+eZ4KAvsS75d8i2JRiwBTz7Dz3N
rGKosZr0l6W2jKXJ2l6CNbNWb36xaBfPMYaTc5m7C0QHGJJ5/rAL2Q6U8g9J+P9dpZBEQpxiMSfw
iyix5L3TQZ+3WFq8djmgrAct2GjCJdDFaqaVtBOKFzQFk2Gz99gK0sNwLHsQ9nlKrzgp8TusqPEs
qExzlcXx2pn6grmq5cq8+Xvl50jF73wen4jUUfNW4Q31cgA3QMJ+lZQfbfI+0EEZmJXmloelU+mu
SCZ2OSptPRKoQFYIep6IZ4lFKM7JkdEJYQI+0bvuEXk+Z2zOrYNQgujG5WH4CkvmlGBHfYB7TpRR
hbBIvdvzpFu+zqwoG8eTZrveQmESqaFo4APedF9W7TAASDYaGTAiaSJ9bcK1PJfrPWWVMBj4ZPX1
i3/yVHCmpga+x5HnIYVKtWEbKRhzPu+SOaCoS31Ao6s1FxeTWL+e9Trdqfu5hEJIi4dIxSZp8MQ0
a/vSF6pwfXgUDxcCYDTGGVbJv1FNkHKeQA+I5VQYBxSNMuF6u/aX5+c514KvSdUtiLRmfMLohvli
b8uPKWdM6lTZZZGaN5NtYxdCO+67MdrQ8nZU/21E44WGh72/9SyDPFtrbJJH3lEgN0bFRczIXSCu
BAi5can45ulIrRTQTqrZAN6aE7o3nb7EDl7bIIsOmNJvSru5IWyFFsVRasTu9JqAuI2awgZmToPT
xKl3z+cYlYaAj2/Vqh1as7vI4bJs+q7wSGgHRLtOAXeZoVGyFnYEc5fBEAtWm8vcXsvEW99QBvd2
CcPNuH/Q8HU24KkxsZrWgFmAlqWnPx6wtagSfPdFURZAZTCHOHzyjpiAiQ4PXL/BTUgFwN/Z+mad
sLSg+zD+o1L/g2cNrT0UmYux8My9pR+3vk5clfqruWM8+M5+9GrouwY9203CQ5RA2/3zx70PV4yR
pndLuLUUr2DYFL6POGkLtlcGoq0ndYyt1MoNXBc7R3UHp9j+ysN4bBJeH2I9Nn0Jyw825WWm+aiM
mypH7SnRSWBzfe4IfcX/DpWZi22TZck4gB+uhCwc2qL0FWEUCsv4RG5Q90m1UmObeV73RSIdV5z2
15mX+BWAm1Ytwmi/RnRzwufeWkSlW7Dhe273xot1afL1gu3Vlh9Tw6XEAdKwC1hz7LOdJHRTRHDr
Vz64t9WDdqWJm3FE6IAL3WXV9CjlfQrfOfHyhJnspLtpfyYgJddvbuoeM5KxXDgkUhu6NwtYWW9c
EqGnDLVM2OCDa573b/1utYW2eLuV+PW4iTI02LdKJuFBejbcTZzWBuTSIyxpHuOCXAPdI7bzRHmZ
dSllDzEFlh3Jqq1v3moY0ZBnAYHAZgPyeneMzc/HMYkBU3bQ+m/0hlkTEm80nK8jISmawoddyZTe
7/gFYxZtsmFjoA7T1jv2M8f3WQxHBS141sBwEUDdnH8pMi5zE1acAs17GKbB/DYLfI8KHm2Vw+Ba
LKlnw8hPHKXsRnFAwvIEKgZJlACxQR44hMtmOVa4WGSvlYWsWRujT/t2iV1k8uVkS8fEzX/lkIiC
OuzAmewcmjnxUhsOkKSmnnb8IH2cLdfZZjcUWVROrQ++EZlsX+TD2ZvU3y8UGTTTEpqTZaXizXId
QaNzE1vboPilox/a/jrCyiAtmCuS/DZo9xK6TpVhzYR/NeUrGLDSgVBKQ8CB69WG8jyUqaK0RnM6
Td94KvjDo0OeE5xcdaSwYrgUiwybrp4UFpbNo6S2J29ZQNlgAWjcEnpBoT6d6Y7gSVgJHLHLNhiB
gEWfMC8UCkiIXmKJ/3wvPxVBYl7xmh09YyoRxCLk2nOYShI27mUmOQtV+/lqNHxj4RQ+s+jXM+xo
l1HTrjoWecTInf0AIniJPK/+uxOiCVVav+dZHM1OGXi7jvvztdQkBc2dXnGsma7pdolD4rO5b8EJ
9vJVFnwq2F52A+3IXUr+xcGi5f5XtNHLNjho/XVOFmaq4a3e+gcsFidthLJadQPXbagJGbAsvTQ4
Iwhs/oBYhc5Zob+44WwpZ0YJCwkjQPXjbMmfTk0zSWEWp7Kgj7sgjfwxWfIwA34gJS+yJnn2Dn86
GU2zJfVyVZfweE8wrhoQyQ0i53yKve+QlCCP4c0aVxE7JJNt4QhVKH50Abm8ql3lgywiqCXUvbCX
J5wUUjdrExgjlgtRI+0qxowJr6ymuK+MUhViyLpnola1E9RS4EzSQQb+Puxcu7P7OlJK3DgZJmye
xM/qWsylfd4IvfaTKcfoeGf1kzpYJ2OEMijBWMxmlmtXWUVBH5NhzyUT70+mT92tgDG3w+hVLzhz
I9pEmkj0Je6W9u76CrdnN+rhkJ/29urLqyS99jATTm/6+3zGMUluSoWYxirSu2tWSEteHN7r85QU
Vody/ceX7Z2fLkManRf3Hy4ac1Sl0k4hmcC1bcu5XGr/nT0J/w09S/3NQ5z1exXDc9f9T0vbBrpm
RxP1w3gWLfs0mSAPS+ochCQ1h1NWSXza+MTMK0IF1Cg1T8sxp4J55cL7mFKHcYz4pzGdPP7ncBmJ
0XNOQzq1YaerXNgQBVw+AWfMuHgFP4Zx+1Yk+00bkxpfScJO66lmX9uW6vpFLgtX/8tWpRnNejsj
hEkVyyE/efrJNfgvKvchCXBIJMhC6xAfDQbARJBGFF5fWl/i5fWnzgyDJ9RuQlFH3qExYyVs3AnM
9dzz+mnRcNu7FITuGFfcybjW1Y7V9pjT/IvVS7MFGAdOSJv0cj4s4pZXfysZM1BF4FeP8GDyCFcy
sd2WgWZHhixyxE1bhUuMHd97s80Y77aYCAYNif+O82vaLLFvePV2mumdFBPBDG5933F7G0JrOfww
nYa/TcZUemYymJfMq1J2y3U2rodIluxfKaBStW1WXzoJv6MOyHwf04PiMF0fugQDpJcE4Z0Yvcuy
73qThPT7SjYTEWkbmr7TM55hdftofoVyi5QSPPH0yKe0UIWkFpUxZQ2rXhXJxRiVsiK3b3UIC7qp
dRpIlNjH12PufxYkwhFRkjUtScDnTr6aFbVFW5fR8ff7a+U0FC/1xcWXySTHimNIPwImcKO/W4Pj
l9jWKdo0pycpnr1DpOQVjbI59Y4tkQFtca+UFX3m/F0rtVVUTn7zz6qhpSjfc/u6knqrv3pL1jAZ
9eEPSUGgjKdVXQ4gvyOzMRlOjw8Obf5CS2i4OS8ASHF+bsuJ/xOm/zbFKLygrBj3hw5NlkScNtXz
4UJnTieA6MopkQFlY8ivfZI58IqskTLuBD9o7LdJTiUJu7aWpWovszO0gEep/s9Bd2tWsVBT2yIs
aBJjbyDmbANIh1SzgbHmYo+GW46tgWTYrrb3nxifCIYu6l8yF88C3WyDf8fEUkh6aX8M59U8v9/O
pNAqXYIq++LFdGTQqbCYAW3iCduyBTHM2cXt0fl+QJB/AeZ69J7hO4fBb+bQFnU8c4tSw9dbdK/R
Pmu3cM2vXoFn1lN7JJYzmAekrxdBR2aV3wLnJTIneqt+w6Y4IRO31/ePx/AvbGEy5MR4fRQ2KEsb
LN6XA7gbFhHZyMu73egfLx4F2mz7XmnsrEatBRwIoAeCRtiQpOp1oAS7HV/+1gmZFFWWybLYbquQ
K2ThFIvTO6I/06U5h5lD3XkST9fh+NBcfoWrGDRFrNF7a+cfgXXMMvK20c4Oh5hecBJSyvq78nEB
HPJOJkiCfGqLs2C9Rxq0jS2nCNWJlIxPuYuEkbMexdb2RURIQgOqzCA9tbUDou8u7tIUY515tpxf
QqtwJptfY0uB9NuxdRQgRr44TAu3mzajlEk95IkywW+6Miq4RI3eEQrr+naMkOlJyBRneP7ju8T1
S1qvK2SC2+YVJEaJjEyaHy7vO9q4sZfMJZ1JQAXBSS/16n08QCdpZ735GQeEuws0z3FSqWaz3VPZ
hbIdClRHFk3rG8lvD+zsSaUhTkdwXi3Bl+r9tDSTjtz1tq1X6SZ4hQ317zuhq25JAgAKHVIe4T4y
ZzpNWBcuUHMCFEfZCr+9UfLoZnd2FA+I54DvpUdtqGVFRVhu9RLNKhQaScMy8pzM8vpajiRBLuPT
xQrVESXP84tnScUpec85DZqvyRtgxGveGWhMRe9mIcCtWTtuDDJGo8A/Uz4jQ2oUKPapzxCcjs24
Z/4H+a1bFwsxgeraciUqXZDQVNVG8OUhly/NKSUQo+wfutnE1yoDtqkSLe4pK+wweX56OWJ0/5jh
3Fp5EJf0j4pSlSEw4wjdgWkFtqU0ilR84Qaa1ugZtpWlv3vbXBVRkjrOkyLMpEFPvgw86vJtJwGa
5O06AqOC0kYJ5m2k5MW3jifL3296FF0pEgqYm6FUF9gUqLuSk7gwzyD18kqFVxGObj5yO6BMIeC0
9lhTqF8fDz84e1Y9FI94VX2JRpUsU+s093F4d02s7r4ntX+jWJQ+MlWH2B+G6l4I+OrVt0DogtEb
T4XvCb8VEt5X7FJHpgYQX2eCpQX2ode17s+n9IIo7YB1VM3N03oWX1rNpsrP1dzbeGjk46vg9oJc
bkkv9hIDJ9AznFbkGYmog421OR41IiiUtm1hECoTxFIA6rjDhkLSzbwqgGJ9J085TdHWqQByQBQj
MoVtGzfkLiur1qq3rwTFlpjT6sP5c49irXZnu6Hil5ZCf5f7oyad6Xo9jPyBtF99EJ0nYsNCth08
JyfAc8Td0BGKxzl61aTVfl1TTWk3Da4URCHEbYHWWKn9/K9Gn2cKNfsVaeW+aNPGyEqygFVgN7Gl
FJ9YziK8vwMqOnH9x0G7wkOIxr6jogd91ecx3NBjz7N0n7hwLG7oVjmnSybqzu/IUYpXIXMf7UD4
xWZSatZyBLF58p4aNc3SyYc1SxW6qjBBz4A87R4Kixvkno5zwL9EVwxJ4p3NfSWHKzEwRN7gq5lP
3Rhgsdhz666V0HViQyngIIaUuhmWODPECwrAff7LxtLFAuQBSJCPblRJZOSOoTptamMnUJjyo3XD
i5La3w06i6uswAxrAQHn9zQVSmvL3fzAD6sM1AFzJVgicNT0CdQpolT6S4rPpjcLrAZahlYUpN6n
IUprzh7f2Jms4SCfMAP9ChFZx6SVF9rU4rkkmArq9jiKTWgm/VP2czmJa5wMu9NjUe+j9SZGFJEt
NCuNrjqLEcdA2fWN91MtBP4Zlj+lb8b40iw+a0NNHhg4ZLy9z4eNo4+ik+IjhqhvW8cWoBcZnC0T
lse/6PWZH98GZYUpZCUkSA6gB4JZ25cJ3BYFlh/7hRAz4oQelrw6uJ2PYix6W/jo0oreAGBRK6Fh
Y1wH4NrXO9HWY71v71YTMG+FuLuaQuIo52u1i/3UU1u4QO6UvkHZmL1frEu67NH+9ibKheFrS7Iv
BiXlR9J6pJy/WgbWKgnQs/TvKS9sReyp3auvFQOO8Y3lqIoxHQsUUnx+vb2ux4K+GA/jqT7c66AE
Rd8iaMatizNEVhDu86svuga7lEb/QJFMTZqIQOjzgoyiV7tD0op1O3cGHSVgS75q6ptvA4jvTwdk
hZ8M+ukXZ5rKEcMY7vmrdDQM8lPHY2YzT0PmqJBOvR5vdfuf0Yr/cwzgPrEEFsYI8UwTrAve983d
uJ1KUc6lgHi8jnc76WWDpv0G22ypCYqmMyC/2H8toEVE+SNxsIhkmlFzPj8l8BXyDz5OrNgJIAne
0+nAxXvmlN9wZZZRnmFi3KADqOnLrMKIfVuBS4w72cLJho/a3o4LO5ia1R6Eg8cZFNd0MdLyILfK
CmkvVKPmvSzN4MoRugcqYZuMF6rRpa4ceL7INBnGbF740TAG/nIqjRgz/ptpqFcwkZ2YjtXolSWw
dfNoSi5xFFy+Q2jFiMLB3beHA/rprekJGJkesWfX/KMNpf/N0vRkcngCaYehvGOF+cTtUVV8CB4X
z5qIZcH3WA33eYo1oVmA8d8NcCxwcBQceG1SZuScY7ZDIwnT8zGADE4QuN2dQ4B4kE3YYIBEzXlK
UjZZt5tIcXluCfjnwfzCf7O+sOYC3X/Zt9CTWKreSedkD8iaDCk0eiSbVOlcLbM3k9LSzI3LoTLV
jdM32KCJhlPloR89mjSNrfHuVOJMr9r9qVykr74REKhIfqwPPODEhQ08MtfeP+3MXezAggSmf7Aj
NDZ4Ti4uNqeMZnfO2FzdKDqWj8Hv9tSk60OrbnxrdR0GKEzIodSJ5EeRvDguRi4SfTDQedOvYI6E
FfBylJAnF19KizKxEHCf+qaxaq1GkxZ3nzJAZmUOLxep60iidNkBy6Bwfv/K2sMJql5YenyLsnPg
PCg/CYNoQQJgUQo0Q6KxSx9t9oKLGoGlmLYCVs/m25QWoGv+2UeEpycnC+TBqoqNofzW6R3bsOVO
DI6eP4p/cC5FmnO9R5ZahTd8r07n4twrvlaG4kjScwXVInkJcjMhDlqmykOWAlTPkcpOyAr9nqPv
tUqiZ5M9qBk8ovm97eR3gFdAZPY6pecOAVymkqltByE7vjsVzWkv2AVyoBs8r/LiD+8PVXrBzRtZ
hJFhrobCWxu4PV45soH6g/DMo6EC7ezgak7fmpvDzJuyDCdbejZ2juy27YAxGv6yL8U5KJ1IEQLD
HOtsBUUwWYHE1zSF/QhVguJimqZcq6h0NHiZJdjmnAQAPaRaTxhUr2RxsUqwBGA3eKkAO0naj4Zk
P7yhz9VAeoOZv44d6VJZrB5CKhjnnDSVQ6sL2T7xOvaj2DDEf6IiD95geApJXiMfSpF2znLOB33F
EdOREsR+Vs23itHf0O0h4uB6Zf8kjWawrWOA7jW1XUa7WMrUIkFBZ391iEhT9TEOinm2kgiKy6S7
ywRcqmBR9ONUA7wCbtvnlvAb0WKG2XzENNSt8ftcFQQOcO1BWQlR9rdbiUo3ZsRV1waCXyu7nWSV
Bs9qWxI0VHHtCZVhFapG4F3K1Ez9/BJG1NCsClzxZEzbEeYbwIuU2ez28huSwXoqCTfYeMdA4rEC
M4F099b440woW3T85hmu1GRBEdDgNOnqah30FA/8zudyzL/l4pztzKZUalwgve9iLX4yCrgWjzUR
E6B/XKF9YPbirOPoFKD/45TE9sDuZTXwbfCst3RDoRC+mbPBr4M4hBwk+OpepBVbwXmsgbSyjNjW
nneC+YL9VghE1DwlUX89vky0L25c2p0J13lrKmTzT9PMEQfY/EhT5pw0JLoVJk9oWdcHgD4TBZkZ
towasKvvmMeGqmkOEOsu3MiQ4SiQVzJcTwuRSCns41HuqDpFDrXBs9JePzwzwfMSB6EVC2OaEXcD
jSrIkAn1Q8Kd2ji2TReZpxoeuqEMvaXUf+/wzB26Du++ufqMFZ5Tm+ixIZj9PEO0e0vTwCsQB4Ui
SDuY5qvbbFW1tvUvX5XxqMQs3tlwgKhhPTdoQyCYRM2c26EHP8glApu9tQ8CfJdovQPCUWMP1UgD
l1/4XnlOsXYTIDm0iN8R+Oizwz2RZX0Vo7noITwis1k3UV1Trzm+yYdHdxAWPZnStG/cBYHXt3ER
yb0AIOHQ/8ZYZTKotmW+y3xrUFuAtG5I5+/0ck8LcpTXgorenN0M62S7bma9L4BD771xWYW4aG53
Co2BYdn1RcG4GopIp66faIQEaiaYKixpPNfXHTsAFa8OYBx7iW743C587panGDysIbMt+OAGYqod
OLAlmnlmylG2HuZIu+gr15GitotoM7DH37rP8jiE4W31kmpcTUXvyZv5ERDdcgAfuCcEAEXeZeAe
wxA1dV97vjBiOQEh7W5guAh+auhUmUOZI+1+TbBm8EqbUXXOJ5QXAw+s6LeZy7l7oQIjXNQmyTtK
Bkbnwner0reHZvaoBw68w0M3NGZhQQnutXwDZi3ISSaylM0WGxJgCBBL0rFf6vjMemwQE0uEdz+x
1NT918Ory/LDt8H9lHn3ZRaN1Wx47xzkC+YYlkvfU+eW8ln3s2s2ethwHpwOazS2K5Ut/L+GCjTX
aSrVv5SxwzDXCsVHB9iQ98acUTUDGY7QwgSmRAIOrLhBBsIa4ZKlitmE6JJO/MRvGjsB6Dyl1/Fa
3hZRDxHoXmECHYgPlQTqHjOx8WW/ZGQFYU07cRa2llQbJYNz0xvdrAnHPV4V7nQhoyoXI4nDT3RN
3B3j4eUDNx8c/oEeBKllB7mrKc28KNsaVxc+VoYjdISd2kK/qps6Vu0VyrZURewgeoYATrZvdWrw
FMbw08MRv/zCawXgYVhl3ItwZfC4evNSxoeHKK2+u6D3t8xUhcBkiJ0fIv25kQCVk3UHKCGAruv3
hWFxjIh2XcsnDmnpjzjxVsK56ybMz4bLuUnH2pW9DHC09xRzRVOVqZdP0O2hupgKiXnoOBthMtew
7HcG4rJc9HxrGZs6Iex15owtkbUGBq301rcjMCDjBKHX/imUYtWrJq5KSLSg0XG/3ZkxY1Qx8raU
O+Gf5YlzVXMKl83on0I5+qV9Rz9getjrZSL3+RS6J2u4+ffG26F7nnPfA7+oA6u0h1Mf48lqTyyd
xcE8+2/1c1BAqbxlU30qWqoegUMIQpU0TfVDv0Uqfq9vJMo498kBthgnNUmZ+5pgK82POm3pK249
zACRPc1TuzV/6iifz3JDslyBudg4K8xkZY0zWeu77owSsD+2efBvObdInQEVXOVqqbg3gMBfwgj7
ZwBqJbSLxNAW7Nt4bdEkTzw8IU/F9omlc8u3P4VZYJu7Y2Bzdy8dch5obqgepupSk43XiQBkkJsn
nvlzFzG8ORMmEWymqu1zpRaI6YSeF7kbyHK5gxD0Zry22sB+rr6+5Qhf73+F9ABh1N/Q13g948JU
YD7R4UiwEgRfrDlyRUMKiAssmDeg1uHOTp1saHNLRuXCb0BO20q/3Ubldu9BLhKlv+Nt8hz2Mdtu
uUaZXMfn+iU9XK1PMKrpZ9bBwc/rWS3mHEEvGnpPQGjqeVbbFHTk/2AFofr5u8lOqAg7kuHSC9i9
5o7pWOS3HPVJ2PwB/hj+8HaKcnyUdictX1PnUF8CaI5ngSTw7VQPuWP3aVEHJczz3J6IZB2ohWq2
/DeiCIGkh09gEIuQge0YcuZ98Pu5wlw2wem2KdRb+gvIMGtlkAU7E7y5y07WiI7wKVLtahpMb1vc
46PjbwJzxGAVwbu/UdfTtl41m+fD1+8BYfOTTnt25W3c3aWTqnZaNJwzUO2Foe/VdVlPKDYNvaSq
rXi8N1ay/9yf7pBZfGeytEJXIFD05JmrdyodgQbp2Mnx7qid8pfAWtY94a/1eEUEgo4wh5fB8u3g
5qfvyPP50fX/ROMbt2Na2xepXB9lYvOpc/lyimIQ85esBOjY/zUZm5aEBebZctCLODiEL0n8ZdUg
Zus9iAjDeGnTfJnnl9l03t/ovmNIWHpjEFM0SXhHbJgmqJgVrfO+O3jGOt3I6scPkf0EWjU/qxAB
8mh9CcYmHDtMqNCZXoGTCN77eGpSGRyOK9EqcadYcxC6B+jBJh6mEhiVoQDAjrOiEgG4mzDSbqUs
vYE8yKnaTtzwy1d6DlZrhyd2Hks047ClvW6IevuUoT58eGtL7CqRzM54vTGqpZ9lPgIINSSKTRMg
YXc4SP6SzufTs4x4W846ValZCn9Fa5B2duwpnDv6/0B53eJG+x0rACawkMohaNbVrEFuixXZu8eU
khJRgmU1cjNx+eeBgDqozQls9nfNrXWmtBGLIEz/bOdDAZhd75CQO2bN0Zv9YcdpoqWj8+U33hZr
L5uEx1hD7syeNmiBi8gcs3HRLe7i5OY/Z30iYyiXBuuT2c9YHlVf2Penk3HvOuJTtzP8FwLMyi6w
/obfimgjdRLFjdUVRsHigNUwzRSvwTCopRXtSrbn0h3Aj2ssY8yWv+KyK+d4TUIJnEG/pi9MphMR
cmmnv70053z6+uXFuSo6e/DwETga7WyFEQugBkba819BgBbYzY4GBCMWsdHFFAvOl3y70KtpQBYj
BsQZ2VDkX51VMgMZZS9h1i8ek48/iu8DEhkX5x/luj0KTdIci1G8ozBDv6w43tO3ae61odFZgHO4
HC7spC0YKghBMg9wi00KgRAPd0HiRtrjlJYOQRoRgViGaAOySFwyTAxw5OcknHtwG+Vild37qWVk
eJyNXa3RoCHXZqnNCVE32ioqLMZAe3v55ThiQVpoZuAIehxm6thU9/28oyY5dzAzYEfvd8LQfjtH
cn4u9fCnkahJs3mHOel9gjhxpxM+lsU4JkpPfnjOYO4oihzXd+zANfg4ULuHQc5htMIivrotcPyK
vo3rS4G7b5hu3EqkLLGGd6hT3hXtKtWG8wMV+TmlBORiPJ5IldbQKxUeXmB4PVK17Uajzlo15sO9
+4fVipjbV/4P0gJfMWJ5jBsqjl83GtrfRhm6B/yHE5OJo1u9oLCx6+3ZEUDNPZiW8Ki3yVrlnxpj
/Bcu9pDG5vZB7MEsAvkq4ixs+Fnl/lKwK7sHysfG7mfhPFerh5mqRKWFMczS9uDhEV5qAEKrWcyK
3hrpSF/QcxmWkWOMOMFBBrk/++Hi43teb5pU6w38PLSYRpiiGwtJwOfwunZLviqo310QjN1sq/ve
5ojovo2fYM4goRH/GQppqNaeUu/MAEnyNjM3WU0GsI4b5ty6+We+tIgD/AxULB0D7mh+fK037GuF
0HfP7DWskVS4H0LWaei3QchXtFGcewKuwYv9/oVjd9oLDOsu6D36VN3Cf2PR67UrNbhliO0mJGh+
rx6XWghHmJSuRcmpFcaMYOtmM6gYzWrLVzExL5imtPYOb/nAvJFEQCsJnahKPL9PsB5XW5BNdNJM
qZJ7aFkXlZFMKIa54cts5KobxsQqzKDHUOW5a3JLAYX+qBsLlCCdn2dBSd7Q7mHvdBLaWPRFWjJa
FCm278whqjI7UTUIsGBGO6VV21+qBa4HdueglY9e007cXLZ3wKU2eKZ0yfb3P0puY3YflXk75oNe
OeyJigp0TojNddp2UCOg9+ThdbDNkgwnUk2U72pa1m06mWoN1p+oLK7JyAL6RXu8tk8pHjjio72i
TMcmwKzbltah/TsJMF9NJGgUKHVfl4p09gbyX5fmTDoedY0Scvvx/jwlXO7U1KLqmwdh5b5kJCYT
LA80/z7vFRBqb+qx7WCKiH//kgKO7QNUhVgLQ4sM3jA0sxRx48+jB9wKC3H+az1B1w4b5FqjupTd
PouvgVxT5joghxWQAMZEqgqGxA4Z+vry6RJKKb8PDe3Lz42HGeVE6di06bCqvz8vLG3V0veTYgpD
+PbOc9RWol9Q8zCnSp+Pn1WIoqEoKyZsKI0xIamU3HZkCTA9biWlbDFSwJf+gGm9kWc+ekHkvnxR
0B7YO991d5zgu91gGO2K03F8K4C/bYSmj5uTSghY1UgD4gZz5hFRLNHYo2T+zw+YzFhyGWWo3di7
nkiRK8Z8CrATUCx1yETtM9RwByzd6fELU4k326PKknDVAZOhjyNcQGDhvuZ6ZsCQtgE0mdSbtPrO
fV7IyN4D6OSLRkuzIr3mXjs8h+LX/mFWDjWCgJQ9jZPj+Kg9Jm7EbUHNDscw6lRthOw8ozYBYKQa
91DWrhm2I/UPiZ/O4eeIdUdFsx4eWemSNVJTY9vM6ow0ar6SbQfu1HHiK8fXPh9vhWryYfAPxIH1
wVx0YQKuYUpLxJupnCF2ikiYGuaVmzDaBJc9k4LXmxectajm3QWoJ+sBkXwEn26obUeKpSm+xVJH
Qs3HorJwkTfxgtIHk9nn0afiRYxvFkYQGINYRM8CG94iEFsDpFjXydCAi61JJ1uBbsxMQHrq8aWs
9pMzcpst5cdshd8GYkn+S1S7iYr2glS/lJaXsWE8ljSFpfvAo7sM2a826YpOM9MiAzaJs3h6jCnw
oBwhgW8w1nfriwTHoJC7WQvI2YbZ2bvyuVJBJ9vNpmZZfcxr/PZAWDi75ScoDCbBQk8dTeHuv7kT
GiLsJO5o4OTkJ3RzBC61GTtfxXjq9/MuaGtijlFlRdGQcNCyLZLJRkZ8kNpJUG3syPt2j1iMvwa/
cKzDeaFkrWZp50s/CBRP0haZkIAezAW3zVT+h9W77RC8UMZHM2MEBpXSGLAi2R76CXTnl31ZqnU5
epKULBC3Mf0pc1NB/v4unujJcH2RlGuk4cjoIbWuaXPDFqwv2E5rfrgqb9K5u7Hzfvq6OxjonRWc
DVkAcxtBy00RtnkwCThHKdYaOTPoEBY2VO/SsJ5TTCNUNI1NOk/4ceG52G7XWMc6Z0dHH0TKjJ5n
3wHgWPrY2IwCWp4se3X3uwB83X3M9du7WcCZ68QujMzP27l2iz9mtYhFn4gd/oXn8xkdkLjVZtKU
iKznbn3G5YS6Bsayc0jCZMOGI/u8PXLyFOg2u1EMn3hdosSBNGTQDtB5CvsR7L0QynkiYqWX3E73
aRzjcAhWC9Cf4eaTvmssgIf2Tcnm4WZHhFBS0u4dm8CebR/OcgVkhqTC+jFZaA1rjKVk45WQ7Nxy
g4UcqSfXGFNe2mxt83Ta/S+Qtl6+6wetJi9bx04BSQ6RlrDcAH6CQInb7qnLx+IZnJX47qFn5sUR
uFp1zZ0lDpsZsPF9C1rFkzdlC48LxIx1b2oSAG8kEPXskrSq8b2Ve7ta6vqkFPleVUIJRBNM8wCm
dAaVXg1WPMYQLveAmIUQkavrUjxt5+G/XBpdTzfK+lWrrHq7n/UOMZOq5bOvgK+WG28b40I0O34L
+ogI/MxspfdPRHcggRrCY8AmTApztaq+8k8NdmsIAXKEFsnTHIVT8GJoGFIi+bniLMj6hNCkMiZM
k0DthtuR6uE/ywe7cuBJcwsft1PwMXiPTud6k6GN024gZ3PPFcPvwSx79Ul889R8+jMUT60b2GRI
Mac6Jd42UzWnIPj1WvEWc2fwpyCcsvB/WvzWhbiFtJeo+H6qzIUG7X8MFJEVnCKfhbsQZQ0dV1I3
zpIwaVvYEWaAhHRmvgVojetZFVI4XwwC5i4wyRoNXOG1VSWHWnnTVBT1Yy8zyzKcQumAYIAvzFE/
mvJIA68mNpz+rn6QYRoObymZZy6IVTinE5lSWgj6n0o8x1+iYoKAdCl4vdsWsgj0IaVlw3tUPyqV
jassxsbDwH1VI5gs8tF/q3s/VwE66Zpel2KIg7j8sUmKLYDvJeL3hYcsaR5zg6RArtZNzFqOrc9G
teQ79bADXl+IA8a1thT6WjPV9mV3sY9SJT85r9DE+mKyoY8bPPwhWR41mbBxNpiZCk+1ph4nJf6r
izMWjVIIFBNmh+ih5Gojvo6nBHQJIYmGLXtAHGp3mK3S3dvw/hyqWanzauMt2o4QQXBUDTtj4b5e
hgio6dxbp8AqF7COSrPo8ivPMLJL7XHEzxywMaNFPBCxm9e6jjbAcB3mIb325J8nJ1uwX8qxhJiq
Wl/lL6/vfcaJZJ83layIJ3R3DowQB0gVC17txE9WotYiB+2deBqnh/3gII7CI7nuePuniDO+YqNT
RIxHWY5YaVDU82CbUowHcI17NewbSw9cto0/8hZtDxSemBuNXsdJNB9k7saf/YlH+MkAsmzSLaPQ
t02eY4ousVwLriAExrQOQ8Nj+01KfAHb/X6QOMpC6iY1Iq/XXBNindx33Sna91/fvW7OYfXk4ZWh
n2JPPnYVjR1F0rCQmzp2eA7d+CgHQm/eEuYWN2z19LH6KT3lKmUg0jcDUDgBVcGnygefIUnQ6k3R
nY2uf70VjC4HXlVtCn7JDbGUZm8+27x9MsKlSS/tkFi6I8F5e5uya386NrUFhgUGJp8e2D+CXm4J
7oCIm1cT9MldFpSVLPvDZLcb5T+11ZwqfF7pzfaroM1ENbuVTpnb2AQh09T/OSCnQLuPz+ueIYM9
+FCPoEUkkHZMPF/cUjsCchEeUzslKIDy9WVmZx9Q/cHT3j2gyjWBJKye9Y+3nLCML1PlBGFuaU57
lfPVofTsNnPLSOFf/oy52fRAbvVWwkeZJ83zT51LN8NM/x7LyxNyh0bSG/q/t8EtyBO4xyvhXA8g
StZJQEPoZK1v/jJrfsNB1jWNc0+4Lh4t9iPfcRRmUfQGTGIa0t6BNv8uzx+VTKL+QragCBJhHObK
qtzWIGgL2X5Bm6NvEdjYzlqSNoB+hYUfqpgeL2zId5lD5h4ZqBiQNB3C80vgIrZp1XYucmT9Javv
wQ64Lpb/Mf4gENfLGmETIxBgGWGaw0Z/radyEnqutrWgpKuwOn1AhbmbTtz1xDYHsyw/V7hnauA2
KwoH8B5jszL90P58PUN1k/rrDqdl7jcFO4rOeKTxcvMTeSLEoII8G9qfiZlE2oJm4UgfdReyFCen
jxjtg0IPByQkmdQr3emHaXXGvCYdPS7nUeIrJjEt3eUXwnqvJS60EMykjq4lltQxG6Sp3/vgFOH3
+UgoHVBj5/ipw0fNF2gfq+ikDhG/PPbA1aLbAthNc2wWvkiNLiOOlv8MJzEPvl1e7+MPHXX8F1sH
AZGhZ43fkl2y3CugdDuyTFWsIo9vJp3SkpUN8G0+WYawor7K3EQQ8sQy0FoCHQQHmIrlgkhOu+Ih
wN2CSIaKjjMkz/uYdud9Jl8SrSnBn3WOZCj+zbOJnGM0gqaESjhhAddFkB7zBkluF6aOGrVlUqhe
FnUwlYRpO6ARDao3ZS2a0ZgsZq/EalB71YFvH1RnspPVtlsUfBLDCKBazz7+8qJxSCRvIvfNDTBL
wyz25Oh4gt3GNfSjWum0mSxFOyrCz75jxkfYjnLrcuBjVbnmHixOYYvaOluJDr/bbDwCGfRvjwRe
lgYF1OqiB6XizXSoKF/Ti2RHd7fDeVKadIQ/NAn+KBnV7raN46WH6Yb75OU+H/Cf4GPCZWbh4uwD
44ncht5W2c9QPcuMnsfVWQLzR990A8MbN3GadPF2vZ7XyMAuV0K2+Ka18IWhauK1aYPdjDQ7PxGM
ueWQO7fVvqgWPbCkqqjX0XjazjE2/ri50LVWZblL9xrBFLbXoP3gZMMkKDQ92WuuKuOpuDAuQlmu
fgigZ55LQsJ2XuxF5POzAozoxSawlemH/EolACTnDDgG9lKeAl+DEErKunspZATe4bkItvCNTG0z
KhAr79zaaa00KqoCjJJBGBYL5Lnx5l7YIpN/C+YEV4RAgscsBf5MgFVYu92krm4+VGyMoBZPTlin
+f75p6haRie4jXldSgc6BJk6CbUw8VSxy+mPeK9cvYhOhbu6aPSKC/+0pEjR8iGhNz/J347CvBL+
iqn25sv+UF5Scs5AxEIVfgTRAAIDjrxPyyKG7+ExWEm4a2p/KLHo7uMso+wMc6tibZ8fR91ap46U
Mdl5Qph8toWn747V6HxpPAT4oaLD8/5GXHjVlXP7E9nU+A3x94SgHAPGxR7OynRaeJ6GkkmFaDHE
cJTxC0P2GyeO/wPTeb93ojhYDmILD4TKJG14GsRBejOxs3IrhGwWOEFJh52qJ5kcsKUk/lNcEA+A
qJZ252a27Z08WfFWZgul+1Apg4nSXPI65P3fglWWCN0VCxI0/UpmgQ2IHCNtrIfQ3XVr9JIETA7x
U/YTsglQleD0hmu5LkrBaPJU0+IUo2aXG/mTzElxAiWysyley8PmLtwab/h7ZGHSg+G2ydl78c9I
Tu/IH35NHpe5AqSud6W0LFFhL/JbIoOAB+RaD39ON/1qE00VZwIyjSKs1qJNvpV56KcQoy+bj9Pn
4k1DZI8DUaZc8Ua/vc1TsXuOfgmzN7UV35xK5+cQJ5g6BXkwQ1Nl6uWggoYgQUjQANowVegtLfid
AsmaSEdCsJhZsqQ0qL5TV2k2LbSZK0OhZ2sDu7bRNKn7PdiL8qAqGOEhLrvicOIk7MycCSKwFWoZ
wardczfbYIR/17HzEXdjTJZ3F44/AQ8okGLdqeOb26R/LothHkPtRugEy4RJbr35BvXN7Z3QlI6r
m546l69KrqdJLlDzqIZWfj4EN/FfPaJvijk/QXylK2OLe8GNrBPt1fHj//wh8GJvsILlpEyPa9F+
b8rFSONB8NYtlUDQ5DbOUiNFz+mDOsyX/R8eyZ4K8S1RWoXlwRha4/5VVaMcf5k+3I1kNt1A6zbW
pOWyDgv3RFshGPVAU+yUkqyB5gBPTKNAtG6GoPrBlYoUAQ3eQVt4+ipdUg1/jVXfMTemVt1jrCqa
ja+FBbr2TtpTw+fgz03+xXIFX0wrUNqgGw6LJSqzyUc8dVot/YnQvwYmETfhsB52egI6DNN4wPeK
3SG/t1rv89EdKUa9YcxwRqo1twBgf2auAom3Xc4Vd8vhsJjIy0EHzWR+PIlKXTkkCa84cmLy3NZ3
2Y+31vzBbUA/WGJoBGFV+UoAQb/rxa2tFKra6sCyPjFdJJbzRWQzRnc/KMAeD+BCSzIuxOUCm9Rq
ajIjPTUu6Nhll96IR9Agkm9cbXk4bViieCqeXNseFIUOTC6HX1WKiWRUQELsJONzRqcUEKY6fBoW
kR5V4dNDp1m9TeEygDHU6mnXeVGTqtwBUTeW2V1nuJNoJ82MEQ5pQSndWJHn2tpfJGkwhrht6nbB
y5C8F65Th4gamMhOGewap37cG3Qkyj5+gMSwKj54gG240ARcAmJv9Y/ib+L7GYbtCYGt53UkMix2
Mg23eIwFYzMptf4C/2+6HlkqYfFAkb+Ks0NfAXTTYvYKT1sqh+MgDF9Fpi/p8CYcq78AMKDGnBsQ
K66uiRkPh2KBJ0AkrQNoaKVccA4pxxq+mwp8tVcTEVajDMOBicWwJaaihrUf9f1VTCD+KzwjpHNt
hCne7ZKPf0ZwdBb7ZiDCwSUMBfIL6HvB2BF0ZZpE2Wo2p3hAtWP2iE5dPbpjir1OJvPy97ikRBd/
i/nTriY1XHQ1bxXDo3DAavOWbHncPS13XKtS0GKaq2erktFEpjE8JEC3+4LgrpqO3ETO/JOqXsf4
dq+wMPvRrJLR2mhsw9Z5qXFA/zcyxrH6ImzkyKZBgDxCKnKYr6WDPKj2p6wsu5ekLYnbiKr3NNFF
0bnrM9u8jwMWPTer1sU3iPxgUkU4uE+aAWf4LB2X+/FdGC38JODwcVsZOvZ6xkAb3V0V8l5G3JcP
DaouJ8mVLBJ1Sn00Qs4DDBWFHF2hsPK8Q1radUZNOYC4NRqRu15gDqqyOGzSI4tUpATswM4jIaTm
DTM7I2GPpvYq15MIeQQpKsIRhay8FIPkRD0OSe/B1wBZ/y5q+KbG7etYZ1bgRIWWmVwcg+XW6hHU
cve7Lvi73u0Kd4EN5uYgytV0D8s/sx4xS6STDcVb3GLLAk/FXMwPpE1DNSM+eV9ZlSzrGcgfXZlB
Uo/r7e4xWE5qopwrV/pL67QfzEhI2WgnknKezMTmEspRsZBhGGrY4ZJGbjcamEKqyq7k/kXCyBmv
bOsq42TI6nMBqj2GZXRtu2x3PTkp9mcKE7Yu1z89mLSC2z9xkC3PT4Sc4jnNffSUIPxa+VEtDlTp
gCHpaje3XPJErpk/VMfZo0XPfV+8p+u/wV9rwVqmtVR3jtmQYmnDPKeM9igZeyOmOZDCi821NO16
ukvFLWtw0GQNEeqNcSIl8C3mRuZOwsypAeG7NK2LGB49+0Nn7jKHVA93sUTDHNNGOuI2US/rqHCG
5F2VxvqIclKooIHUbZ2y4EF3mp1NO1vpqZOhxVkqlzhtPGHLCQShti4lDhsiRLLdMcBs9zRkbr14
aeGirQisSXWQhvulJ46vv4Mp32eaOYoeLP34Ko42i/JWjUJHjA/V91c2DuOQNE7DTVFVdcpM+/4f
2yZFPJ9sCTl5O1jpPuSOVvfFAMFSiaMKfAkfKWqVQf5XR5f7iffJSydRpS2LLP2zshHlTLTvxT2X
hPklqH4i84vaY10vxclzhPusaHpT9I3OHOHM0YNpAZfa02PILCLHxfB5Kjcdrye6STb4LUc83uZp
5U0vApaoH00kjrTRphACAy24X4hG28XtiscFi7lezdfjppkzlwe/UZ2v/232vfAyTbsQSOU0NaaL
L/MockVpG7YLcZDdTlR24Wgnn8rN920z0TZdbFT/QMtpd05eqhFmu6syVaWG7NAWJr9YaZlht5Ri
uTnEzLp1QZ9QQqt1xstcqwtmHoKpwuK+q5aqVQq/WtRxnVAtCTI21a1j77aYDsCsyz/6RNoWUPyv
vNt9Ldy974VXBJ0ozKWREZX99ZhiCZV0MSIfg5w37vorN38fa7iDDDkPRm/r9iDO2+FGfmXOPFOU
B55drdpnRDAFeploufJHz+RSrELsJcC9PSqY7+hFP7be2w0xbBReal+Ro3i0xYVW/NTdiZxFBtpN
fs8gcHWD6Jrglz+hr/+6+9Pj6mAXQucdxtJT9vHeJgJhoLpQQ1sWPjo+G3SPbqF5kbXfISLyUfTS
RteMC5PS2GHWdx/GrRGZ76hgRB/2bSN+Q2FGlXqeqzvoEygJ+IDJzf2H7d39LqvACfL8r3WbvcpI
K6MIBF9FCPRrNrVTQqkkJQdxs9ngKeffET3p14CsSZ8YpFonwLbtj5KPYgqQckDhuZdAIKuz+cZ6
muCycRcnm0+GZCGg8ooPviu7aQtSeCHghYrv6B/I3Zuv3dG2nNaeteRl66nNxZ7lD/4gXEp4w0QD
T531HwjS9FH8QlMzTcnCjyxQ1tAvV621k6/m9ebPUZY0EL344ciqmhVjSoW+MI7bDUADdet+TRkj
pMgR+Me6ivtAYiZ0YXGLUfxoMzWSBvk62Mxy3sKul0NHPvyXNqKq7nrIvNnuh/KrvpoGyZ2RQFYk
uOU51+tbUf9o3Bcr07N+19VjzI9+01YXsF+Zc2AZQlCIlDAQimw7eNMWBygTnpb/sCMPd83eCGJ+
PsPA6Tj8ED7FfIL0Qnlir8pfzLbu9X6ByufRysQ+qQv+L8tHA6zbD3gVmgPTIV4kUbgmeoPFkk42
KLrnSyjaXMwmAC6Sp+4erUvAJeYxQln1pNEfEbWTwJXI6Nffk/wWaN83jy3xqPhREryxxlQkHMPN
aAYxBsNsc/20prjlHNCnHgg4m2i3HyK1TXV/7V7xed/Iz+XL60eNIU16A7NPrmcNXH5Vx0X4JIKf
k8d5tZ0qBfpxoffWWO7ckFND4AOCz7zJO1Kks7Pip5PMIuDh8gLvAwNqr3PZA9FqppYR7iM0g+Da
gmCWh/L/POPd81SWAAU0+iQncTi+vr2pYidBKI3Z7iOgaRnPC+KRT08PaS8E0rLYb9niYfXMIZ2F
gFfGgKfb2jEi3Cy+IqkqMW56WhakfNcvriuo5EJHJJz1LRIOANQOCabbkUZDBfzmVE1KH4EYm57z
KKQRW5qAsGVJ/+16fNEEsnU3DTqPlv3sPO7eOZMYxLsv2d4GeHdWSS++a5lW22Hti68sIRZircVz
oBNCFWRh+kUVjc/dNilSVFZx21qZ7uu0Q8ZqfIRRtQWFZ/pOadps798f1JoJ9oK3whqNeDJQZqPm
/rQrG9ikNp0KHpHDNDm/oUd+Sfhbsj2W6mrwa3taax4UxfvuINSLhj4Ra4fdx8AECDA351vPSmvz
Kx6vRNaGk4EthBZbaqt/6xsPiGlBve88kpzxHNVjoxj6oAa9/lIFcNn9BoaX3s56KrCKoNRwN62A
eghSQJK2VMrssOSjEHAQ53YmB+Eag88dEeOb2pYzCbF8fFdb0SlH3Ln+NyHvYvPDd5pvzbIfqYk5
BqOpYbaYxN+1Ff9wdUmiBZ/HPbFKTJr5AyzPPXJ+6WipJh3nUWg4besQByMLaFQiVl3zhNA0+qt3
qnw5MFGfVP8XRXgVIWl4Kwur2PiNfqbqDnPptaSm2IbYcuOwQjthrsCryU4QvIZaoeBXlMnbZfnZ
0AO269vI+UQnc9nuuwGc2FBkXR8nU+qf8bB2v6KemrmOtf7J/RVPxxT3CY0EIsHuzDmOIIsw0uGH
rBbA4RdXKx/XKv35lEj+McDQHgKiDEMtS0u1C1DlTx8JT0tp0e/yV7hQ+b9xFLI5w5W56hdFVBoZ
5N6ZDdhPTlo4fSPI4XAyJZ2VmgW7lFtdW9/tDupwAjggg4uxufT0yZC8f+j4vxXGY5bIQ/tQ+e//
W0cfH5EXibiBZv9HQ1vDEv4iauTnYMuaNpEAO6kEp2Z3WOYl7tQl5QEDYhdvfK3gwszZviWeH/X6
LMsoWLKxdCQ7/pxmme0yWXsACtU+yPbKeUF3RYFPejJ3o4km+N5Lp/s56bmjOPsE6xPdUGaclTdL
N03aslbeftBrJHbiRdN5SsshpXuOx5i+obCG84BFqfAeXN6ikcgds3HL/3x6xQklWfTZeI9svBd5
3uOjenwBVqyi+q7qqZem9yro1lB4U1dYaAdtA9pAQk7guIVbx8qzqCe5K6fjTb5NaDOZ9rJ1G4Ze
IMRDfhebuE0FiGwvjPxc3vjzmTZqJ3O+35TRup+WvvFU8aa0erTb+G6GVOpxbCK/OZSwgduEjad8
tIRGuJP6qhqDRWA3CnVxr6AwvmMzuWKbf5tcGGJ+yxC68EqSP46WZ21psk/FvNEcx1NORmx3Xlv4
v6GvNpokUDeKP/Uz3G789oI1yq1IZC28L/LRxDXQAP4X/0U72eznNxUammQq2u7HRV1Aor/msng4
FbDvirW/LKAqAP56FLExrGPxwbphyrHX3IAIDHYsNlu0eXnr7xsz7vwhuF1tb/YS9UuLJltJuH2x
mhxCd4u6/NCGIBr6xwtps01AodSduRQy77v+xurMuFFcqg2WLL7y7qc9X1UyH/mhGuemcOA/hzlr
tilmvhIu9O5gl7+V5EGrI06pSTq1unomDcM6NvTOeMYnqbXTv3xncv4HBl93L0pDLp6009tjOfdb
kj+uQHS41veT0ffiXA9ajS+Gz2W+YcxxmWbPibedt941dDWtCOa7ev3HbizhfPBhl5F5prOz3XbP
cYCBrFhaL5ZlAm+op5XqFeg0ikHMrSTskKGFMoKmjRXFIMEBKgd+bp7u9SWacZEe7do7XkCmmDWt
IcmwML57XFJdfvmD+E7wBNOUT7ZnZ0ik8nuUlsBYcu2hQxMvl3KXCUsJ3wYwwP0zv0pk1roReoOr
NV9co5U+dJJ/3RYhN9Qoh8AcyHQSaZ4lkJttGHpbSIdV01BbazmwKg/R+LIaEQiizDKO9A5mYuF6
UVb7JgD1z4jgL8P7OZT9T/1k+F4gEiCva9TQHH3TR0S/SviIvkqIsIuPkR+dHo9X4az+tnr4hkMG
owUWmcJilLuNOhEUzn5fVjear54AAaf6ym6JQq5dnBCrYANxCfxBErdBFDAWE2yW0IKuzo2qDT02
e0u92J8BgtIRJKUbjlm8jS9tLrzVpo06gaZXYtM5TeB93xUNfcgIIR89kMPu3LClSFaRd+7m6rqs
ywvP533DBnfVZdYeSufneuofiAPVlgJoMCurg5qVXLIPBbl2h8/eMGS4Ot+OioldPh330ofcrbBU
rBxbfVpDTAeMkz53EBiKsdpABNMc+BcGt/+MKYt30L/+DOMWu0SdZ+8xF+zNE/jK3sCfxtS9FW8O
rXHSjXHW0iZ0hiTzN6dua6Qp3rP43dkh769R6WbiY3TH/8O+Sz3JURo9WXqSZ/LeUI6XlqwDioVf
rWw/oJwylxme/4FGJJzebnRiViwHpsZtW+txKfsSj2KjIGMkLgsMuVWRNOT+kgEATUlB4mZf1VUS
MAsVrCe7WSb0Q2LrNzKnQRwsBmNv8+cV1gpNUNgEKmRv/Wm6kQfiegVWazYoDqT693b0ZTIXqjdN
2QhsPVZ2nOMfE5Fwt7jhBN3ugNbYChACkv7a/l8GzmxcZ/RJjdXtcdiGYaX+GlWbz8yzvYN71QIs
9gaoZZJ+eYiIDw7WP13xscl39NglDP1WXhsHnX0I+C2P7kkR0AB1tTZS93H2DPnsbCvLPZK7GHMa
zLyWA423qGkhEbjmbRBrVQjumwwXeMAFYdC6XZGi8XJv1stdURQzqFRQyaV/5A08sNQ8xwhqSCpJ
IphEDBPG8gBnoWcIqJ6yWaC/sTEOP4ozuNrBgt54wER1YW1E8yr/jxm8U2bL9tybkdLTrh87p6qm
iecHtY0ZXzr3fOIaFTXSzWITaNStrC62xSmQS/p+4IdZk7x2I0W8aOmQ/+Au0dqxvJe4LNszqKV/
05S8CZoJMuVn4jkCZVgPgpVPZErEBE7eAVMIX8OMGh86tgy8CP9zkZhzKA5le1diByOmzSLpHrGY
h085xBPO8mlhSIPD7z+GNkt6Gs98sdatLQmOZvwFWh27W2t2ZVGzCbwmTAf5SGW5aFOB5VIN6Img
CKn9fUMSmRZVMGAjN8NO4Yi+5Uf+z9TOtZa4C27X6DjBl4ao75XhNRv4kNrhQU7iJGgZcy53a/og
Gke/p8V8JrHx8UeCwRJrJROdCHCmV1Xax2NbxJZkMzXFrtPyGhmHiDHt8PrVkPLWK3nfL+NNNK/k
rud1Kw1skBtIhJQDpNz7EW7SF7zvW9l0VK5WfR7LhlcflJkst5kGaMBk55l+zYnqWvHsQ2xKrHhC
MA5BzTK6A/o5ZUua5s7SdI+0RhfTDKmq/RigCD86e3ZnhwkatPxZT7Rbf1RRVKNk+762AdaFm2eU
32XGEI9n/muhDQa9sG1QED9s4EvVoXbCu/+AAUupzOOtRq3PM+tPsqG40o4ToYw0Z8due+oDXfrp
VP5fJB1laFSXf4KL9aP1BZAH8vsMEJUgOv4zTjWjAI98VxFFJgm7RSmo9Jck4sj/0b27buQjmmWo
qBkr4CgjqVoY1xhQiC00dTcWjKIUCXFxmae/S61FMwnmLtE9WNJUoRMC4m4Zrny0RX29siJ6BN7E
06Srxh8ITkuxlv07zSHN+pKFY2DzuFL3hN5vtwQLJ2o2ZvvMxtffGee1wRCoiTcJJwdEVG3JLBic
LfimciAMUuhnEcymirrRmV64kpsaICgozqo9MieTioqSBZExMU2ZosMvZMEOUiQ4+nD4yGrkWyQq
PD0f9K+ksabsIH6KTpdq6UX458PXpUNwyx/vPdGqlVyjdCfGBH4PrY+VbwgOhwVkfwccXkfR60Pw
V6iW6CjGSOdNvPawh1VMk6LlVGMyfUwFeS1PkCISHsc6n/b0XHouV1F68QBPkNQ3p87A93zm2LSm
Tc3f9DWTzrLJ3dBaV3sUxHwydOX3J/uZoNviHzpL+GhZYet7+ELBc4wScrcXNweSR27BXMSuQc3K
n9vL9PCzIgahXQ0W62LUuLGprfCllYEH4XuOXhfyu5iaxu3czUtbR/rjV5gWd2SPgnd/wXDJ51im
tqBOFyNIPTRkQAtd18EgXmGlKjv4pFs8CG7kzpJ+HriWs58W+/bvc0Hw8n5W21D2/lfan9rzfZdc
scIxhk+PBg1jspHgtptxn0it35Th/UZ4J+gnj+c61qnQqSEObFURoGI3E7WXIDN9t9d7EcqSuNeP
zUGnGlDVe31l0P8dAOAC7j7veLYb5+rZzv+suIeJxgmwXphxM0lq3NsC6Mc9SWgGqKGMW6MQ0jsw
9UC8tnfRw6p4+p2YXjmXCWdrM8VtVKALOFMYfNnOmVfivNqCUS0dPGxFmGWFhoz3q+mEKDUoQK9i
MmFJ4PtS3+WYAannePPatgl+aZM8JOu4+Fe3yOXE2y3sdKwS+z3sm6DxhZpaDvRZWD2EjPrEoCDu
o5EOMBb+ejcMffEnMcc3ZbJ5h1bmHu2aLCLPli4ChLrS+O5gsKZ8eDp6YXqHUrdfaRkqDBli18Bx
yQWgRtUGcXXhW9ggyIHcGZ0JKsT6SslWEoniY47LeaJwVxQn7BXqVXANFqlVUQU/yu1NVioJpcDz
rOCgverw3CU3tbnmRIk+ZXlX/6Y/eiqngf5s5kKyrIk0pfaDMn9HcKLXeiSeauBf/WGuqqvVnPoS
gim7LBdN5hTlt9GAX0K64wZE3V4FM7qAWT3H0oNfxkVhRLY1V1P8M6Q5YYjU3JkJdW/xtojN4Uza
D2o57SZ2ippc9n8Ms3rIVn93b2xEBTe/HBGd62ugfvfYF0961Wt5ZNvd3js1wC6ll0wuMqpN3E11
wNvexqb5OXL3Tm0p4NuhMUeKJxYALVzwnW7v+/i9UsQU/QwQY47KKqIg7+nSoW/fnfWI31xpyaJX
4UKM7z9FK570MTpmL1MN+bhkIU4l9Pa8oVBko5mibqiWf6Qn14lW4i0QSifAR+lps77TyqEdDU2w
4mH6aZML/v1gXMdRO1QDWhrHvmW2632Uzc/Fd/l+OiHZfBR0H96cjpZfy21JAAUQ02xT9P6oMLdC
48cusP0q02Ywq/KC+ayWaIwTJ+N7GthmzbI2FHixmNbI0xoVyHl0HOlx7c6o5KsjWVJeaihER4Ot
tCbtc7Izd+JZ4k2y4t70sia0stDEFzRw69V60giyJKSdr0nbmKL1X67IrDl+lTd+LNlSj+qFyR2X
OOUrKeMw1OMJEHsTWU9k+fBo36NXjFrODIH4OjXwjzDJ2wzbLXWQ+2lL5VUPueW/CJAAwYILJQuR
AuGioM9gKTNO/OxTuVVyK3X4e0njxDvc6vC1I9ZpSsnpMVBoKWFjluWsZh0z9f0+clWsaHhr7qyT
Wx1D9p8rCUwFsKTe8JjV16CzQ983eYkt2K6ETCY89ezTcw4YnEh4wf7gR+G/jfYR7TG4otuAIAP/
me8Oc2/iSJrvQl277tYZRxqXHhBGRm3Jjw8Q8wdoiHrRZMEdenyseLRt8KGaMrkm02ovCj8cOiLs
xybOWCvt8sOt0BczLTOwl4t7zqG56zJUE/lTTHn/fa5JopKb4+TCDDSQKqd3D5m3GzxXSds9uZ57
/jtbG81kKsS60KfPcElpC0QYo9mHxv1cfSWN6Zcklgr1VRRJomu+YUONADmrcJLOCS45FswcD+jV
rOij7xIF3wDoX0mJQzbmJ6cI4Jwarto5VzoGTsJnlzjTVOI/aV1HxJ30uL5CqGlPqRKkYOiqSlH2
SJwx6PPbSR25wcCoqPoT8iNYIcEPxrakJiqMe9qc+8t0hjtuN4E8wUC7XUzhyyBInAfHRUgLTgXl
ZVi8aiEgT8ZoOA2LCn264qWxnPU5Sx9Yst9n720QRM1VjDgQ7UfWA2u4aRpckaCFQ9sRqT9eyL8i
rFx/JDAfpLFmyxASs91AptS9uOaJhouabU9s5J0T53i329E+zjAzWtiEqLyMBgKKNY09mGK4iz/5
B+5N4mxFlizWUPpScwWlSaqNwJcZMiqsqVr5nwkdt32+WQBlPgxHTOPOj1/sRpw+XKynIR0J5hO5
9V58eybf25ik76g+AhhqbILpx1Akc2eWhPsx02y9pMrfXKBAUBxyM5J5d0aAwn/ZQT2eTZa6Uquf
ueknG8ZEOisvm+j+oOxTuXkDbgOaU8UylBUEwj61g2YuganECzusxJXpIqOho88AaHLagF42tqU6
Zp0NVdmWbUO7XKClefjtgjPoL/YTnnGtjatJife+EVWGYRHrIx+NYo0l0Z2weaLJzgJ7oh6X//A5
36fmRgZTi78Y4PmeDltIIn+CausjFvEUsexk54BxExr71Ygca0xU7kfr4cuzO6U9X1WB/3hIe4i7
x2X9eh4ZeKJEsSD1U3aEusdocdnGRLjMYqeH8UNBCEXFlf8d6v6K0DVzrbyOE3rTJ9tPG1MQJAK8
bzC8Bl+Y/uJst/y6ABW8FNikeF3f0SVBP0/Q3cOEbXFMe/7prUChq5Bw+db++jVajfAWt6fduFfz
oCCW1lf7FNl+nBlZsg/j/KKiGdz8rx58RoV+ICl+YKyCewdP1U8+hw21k7rS4/W9JfDqLk7M6lqI
dyX5TQaE+SIFqptLJ/vPBY1MI3XEk4xXTw9Cf0lGEVGwg2GHkAIXwob3lFYhXyfElOJyJqbQq4x6
lTr4MWC4kNiE3suSh+2R9jSyIBXMvf3mTfg0jIbhbuQYSXij2mbiFZZxAsAzjW9F8eCe9GIqwZIx
8jfa5CvYoYvWwUPY8/N6wv1xHR4DvCYOFsQKSQv0drslIgXO+VuUira3m4nfAxk6BBRaRwwys1s4
wPSaP0/WxIBsJVQgODn6JkggnmjV0yCkhFLwBb2aw39sTU2lsNnEdDcLLOz994V3szbo0HWhXH4A
irLu/rE3BF3c3nttzljmT4G+p9VRZpls1Y5QgKsnyl9AY5OC1U+hh32p1xPqJiRSLfVrOuHiVOdk
tOVDjf1omZrfMdfXQ12XkIs6BT+u5PiXH78V5zXWlGxE5AGfHdz794yVFotX+rCRT287N8/lBvtk
T29gKqLHW20Kw2CBQDNUASQDTXjGhVmC/boCIOuzuwyeYsrg1t6F98P9e4gm29pYzIhbGr5XrSl8
WkFX5JM0z+pTbR5RYjCFLwU1AY853QxcgsP0YCsc9a7TVoNT/M3Av8CDz9MbHEGK/+kxYz83BT0U
HP5xN1vpBbEKYJ8VXGCJ11Phd8QCUMnAS/bcsT3ZhFIt/f8klhiBMmwaWS2Pb8yblBopEPWIf8cI
ivWagUD0UPOc0LUk08uVaXmjMHw6zqhfkdP4ke4rYVlCKNqwJsRkf/5G4r/WB44Uy/tk4glvyuVf
qby9pD7iliUm1mgXme3LhkB8dafYR6pY9JAh7BXGOlUgJHXgqP+UZjxXvVlaIBhFS9VvYMIU6vS4
oHZQuAP5VNvrCnUxTrQLcTFyXxBCOl0SYFjmWErKgOtCbdYInDXfb2wUN4NPUVFY+xyytaKBveaz
ACdjQFJmujBBBenv5Krh2wFTraNM9Rdu0vs7lJNPQYK8Wx7lCoNVJ1yC/KJfKegh21FTOciilsxA
sasqvvVnrW2xvGXC2b2wKrje43bJdJH9YVCTyAVVfMVun7iiIcOD5iNpjBPhO4UWQXWL3mPVtb4v
VjVMQaek2pLwyfEJP8gLPTCc2ExZdRkV6YWHKQNj0nauknSCWhBcZ3caS4QqviiazhqL3sZoi5Nb
ZguTcNJ6PA4NoyOhTe/Iy9eUJQrrwb/2S8SYPmJ0PKASB+zJtv7qIDNGuVIV/oqeKN7ptdOx/9G+
35ofoDX+vw+QgvpCAlddhWobuQ3O/j/emCOoZ9j0Dqi+3SuAO/QaFiUy+YCuAT6TFMCCMOE1XvFv
4WjbMP2n5tr48t5WZNq4RF+nmHlEIXV1O+IRzKIqKDAhYP+WzwAMVohK6IRJXIzLkfOhyjDJWafB
p79lmR8PuHNROKWWnDyhpr3mlS0pogq89OfVBsM1IelVD6Bf65XV0jdcVQegKDL1mzmOdJWxywSA
Enya8WkK5dzyE9RHL6wi0Bd9Q7QR7cp5PMB+LeNW4DpIiETtIuzvVcx5gNRia1zw/fHn7epi0m9f
MP7l9Yd8sRCwxqlydZWF1o0XIJpzdxCMtB/lFSQ9wPlR+3793llTn1GLSWcOL/qw242SW5t462gJ
AqEso+Fri5WLSaTw+3V+Ps7qIW3udI9HNoeeTk/f3S3Fstxc2/5Og3li2OZDcuat9iYE+Y9iMDSO
JVTmOoGKnJzN5Gct4hXpMWhKCgIQ9YnPRmWhua4HGs3TSpNNAFuWsUgNIA566RThObsBuemJ585U
wqDKjnjOmzH5R/T8kiu4VnCOxJQ6en+gd240gq7p76i1b67RVZpBkYPc5EJG47tMlqu99jnsPlJD
v9Sm4yxMBxZpzSM7nKT+MbdbbHt3VGQnAMmL5D/bbmYkfCsCjYOA3UceI/Ud+oRSDXWaRR6+0h0y
WXrrSySJrQV5+EXDHYQrJGeCeEuu+VDtS2vAwY6KeHI01uHjybI/4EykueoVxuDgUeUs8VQikmvY
CwZsmrVKqpX4vK5YUof+QSgErGKHfEtl2hiIJcKlWGQ/TcubItcEtR15MTe1+aWY6jHv13PKJaQ+
k1DtsMvFHyXUiBl1Z+UPHCs+sTmqydXqd1megI7FmQ6LOnUxjmpi9UPzAJATWOlJLU7XPrsPrhp8
vsDnBRU49m0ZoQQpSbanbWfcudiiyb7j8JtKNxSX7VfrkgMRP9lrMvHRBG0DCSRHV032wK0YDV9O
PA92NiQlqrXSSKRWq4pEbGsMuuxX0v6CB4tWlw3beOSeWVpc6OUT3Hh6+AT8vNMrhWJRL0t9whWD
hoQBaVPNbBzWxbhZuIug8z9aiP+Hi6ZNf7RUufD/2qqI8sNXaCJZr68XCZTuMXsJb3ZTWDTefsy4
Kn8V7QFX/v6Mh5e2z4YZgneAjpseK4p+1ccQkcVbBysu9UvklBOZF2qBjcUFBFjePfcs92mlr3Rc
PNrUDrrEvkPY/0Foiq6Sq0f0/D6/AGYICm8hLK2z77vHUwIG7TSBcajOnMjFCQf7ivJUc8jo/rpg
osVAUq0I9akGSL0COo6if1oasyR+r+Q5yecuu/S8HYdzw07nwJBJLfCawWXO4dIVQfoH9reRy5As
9WMC6FZJOcyZ+kG98WGZavVGLt2JD7bFc98w2o0kZyyM6wyIx2bkbBwdB5Sycoxmj1O7ryeuNGNt
eL4Acc+6tBapQzUqDDGr04t/3R9qfSOy1RUEgiVwZj4elvysJ07AsulJALXnFdNxXngwCkcSlZcC
qFuBc25RV3PyPiCRl4I7NCrdfYLXdcw7rzDAgNPdsqmyExRBCDOOLARz27t4AuXh8AgKocE3P5TQ
IgVx45Gt6Y62vpRuMKvXDgQviUo71UCku5HsD8QPa9ysF1JRwE53pfPzp/9p9PXCLQQmryRRKc1r
r8/cA463qeGGAExoWNsKor6Gh0ueAXLSvZcHiebYtZfn4N+VECSTTIZOlzzlv5UDR3eGqxDWmcRN
scl78z+GgPVi1xKRoKkPfNtWTGSX0BlJ2gcmCMGV7UdN2NLU68pEFeGpwW0A3r6dywhxZBA1yAxs
6bYwIOGevy3zmWsEYFGAOsg0vExvvQdHgCVtSpbzBjOfEsBpcLU5XBJyhU6I8ghLsrBBOYrJdkHL
mzAdJ+dPqizmWW5FztgPqLyIPzYvmU7Qc6ZieVBAGiULw8OIsdisFqriCWvCvaEdK7WW8vfWMito
PJlnA9qyir6tngszjzZVPn1OIaG/bX8DtfIWbTPuSoe5nhzHeHDoed8uCp38vPPQCoFDffX3EHk9
oFW4jlFJXREr3vNHYLuvLuWx3UHvCJepAQ2gGGyHC9847CxOKQZu770rNc834YkJXW5bnmTvDntm
sO1w0r0B7qak9ETGVD0CZx8K04v1XxNKkAmZsw/1FuvkTFOuQWYl0lbW+6UOB646Gt91Z6g/r0b/
RSlCrcsLp5Bke2pIYfiivEqLBH31P6PUFSPkunEOj5n4pgSITLoiXgDV5Nyb/kUtrohwiEHsP5U8
696XwscJsRhSje2owf5sCZJYtd/ENUwVIJmy7+dIvy7OyhTGDjOdHC+q6+okhzitvR62p9N8jyuc
u/NTZ6WPq0Fkzi7BFC+b+rs+Y99dqEFyW7n1tdtLluzeoxH3uW0ZoHPb3AQIxpAu+1hH0paEI2SJ
ioBzOIoqDyUXUA8N65vQJg266qFnQOK/y7uMzSoQJ6/uMWq2qHpTg7mHxHzY7s1MSmzmkgVp4dPQ
TsmXu2ogzu3YA8r7/XoSS00/viSoag9xiHyNMnsl9Dj+T0VSsyNqHrNhB4AFeTYbMT6YaaN7Fs3K
UesnnwyXb96OJmXUNTO6Bfy558kVgNEzTWHGlYv/cmni2/T3X8GfhY7RWKLv/FiRSwWc2uYF9Pod
zqd/FTPVmlNb1ByDbSNJ6p6cGPp8bbW0RglpmLw7UXV8ZbNtueEPklYFySpaoqjN8RoyM08geRPG
ry7GRFJBZ47zPjdgyrf5Rmq81xPjTWw2syQ5wFboUYHi4731wPoNENXmrnVjjan6ZqQSyiBI5wRs
avni3j0oJ0XZyzch8cNyF5te32EHdcwIcrbU7V127WbWHkoy0rgyPJLI47LlZzvsRBrsl7yWibjL
0Gis1Cl/iw2ALtsQAnQL73DHUkoYz3wYsHUVlbGgsm1CB21LYW5JalgLxOibfyWOW/FwMxk9ztij
beASmbDOtU2dJKEjddxKtdKNOwlAhifTVJoSZ4rkRboo4pPrhIgljB7527m2gPctKftts/QwJl05
n0Y6aO08vOh+EyzH2NhClz6errvylqYdoqZbt7s9h2zPIHALZw/hjwqkJH53ngI1qYSYZTxCF0D7
B2lHUpRZW3jNsYmetWdSR9W+LR62N3OtpCw4FFZPVNYcXHMtJInwj3xMBKUiHN701WDBYQcmSHtz
wcX4FNIqO4FEr0gHp8/KX2MAW5W5/3EnPVDEQeKpodQzu/MfuYh9WfmUgWinV9TFKEDRufOIOZHB
gpHqAmU+iTCTiUcBcTRrPBynPkPyGZB3/6GrYksG/dTaYIyJ5hRJcGXcepWsLk+RWMpaeFkxVGp2
572FbcgVmAFWWtnD16hopPSBAvUAsfoEXewoZfUL+uXLmhLTXujCd2Ea7t5pYqBNK2aqHl3Mhk7v
Y6gjMavnhngbpjuoqAfZ1ORUWXCQf6eZWyUTV/tx92ildAdV+50t9e1H1LMq0v9cdZnHMzGaNgjK
+ATqHz6uIS1seycquWaxu3vXGpVJm5gM1u7IhSZuBUzVQhFalvC3grj8Vj9f/oQsbU23ki1xgg/K
I6pszqb4AOj2LdGcHN0dysrbroP0Xs6KPR37PrPK8e/G2GeerdhEU7f3SvdV5sqyAse6fDLr90Yg
/YR6+e9D6IXaUDaMN7Cz6/YB2PqBd2uPpNDqDTn/RG4iFdkv66jTC+iCVzimK8Fe35/hkeBMdka7
FbQZwCv39EEwx7nSvOvI+JhE0jEBUrQWPlmmWUclxODejgrOanxJ7a1GsjIsvXIl7tFdHhGExWax
p/Ch80FP27/cdpBwDiFdGnYKiUcfMQ8opKZ6ejtZ1/rc3UmLvyVUgPIzaMIzkjfrRts2yv8HMPVU
G/MnQk64TP6HQkRrx3U69Uql1363SKBKqt9LQBhdphDzKcn9XAF37xANA6b41g3Lobp3+DyZ6L6w
68qbwASDqLXAjdIyXhMiP9vzb8t9YS4lDEpg0NuvbmVlFD3eaF8E795FiAKtwKR/sEsENKZQRueU
GKkQyPA47s+aAI+9stmvpPca4XMVlhEo3rtP2fRMYBHrppicgBVCBAwZH/brdMk9aNObqkF09ueA
/lH3NETm0sXEL8ToCR97jbaWZnI5KWc5MW9C0O6C4mb4ZiAXA0EGSbYzc4HmxWRlWXwi3GCCBM5g
WCQK4+UJ+XLC+ekzzEwEj9UJO3jMr/7FajwPr7aG7JhSW4x5nx0/in8DjJ+eJY/rOutuLpfUmKpF
18y4EvpvjuiptH4V3eiho8XpA3i45BOCGZhNSFbTPMx5fFkE7XAGDKA/ndmJtGRnol1jdgOY4XCq
TIeR9/eA8hruu3Ex5J04abUoJSyoTw8hUawDQaFghH+ER9yQtW9Y6/oOZ1cnnCIckl6srPTIkMvy
Xj/tJ+udEPssdFJb1LxXF/vGBDY6MGgLSjIeVlDcEMDi016dlTA8c+3s2eIjqU0PYFmcdcZ/47jm
PbceML4n39KyqhV43ANCxggrfogkWzRR33f9ewqjtVy65JGlTGevqMxbeHds6CED9YNR5PCw6V5n
3y50frnbl3FG31RcA0rpjduBjScx/vOZn01642XOjKoQO9c/Mpj+4fCKbYWtnDTQFZXAdZL5BP0U
7icPN71ICFO6VDaUfsrKp7VYYwiYy9jrE2HPBLkXExP6PiUv+NQ4/yAgxC/Jo5hsdO92gY7f+uEg
YmDu8uUvAtF19+hPB1fRl6Z2rs9Gc2PharGQSf6uWtvCAEqeJPUR+zkPeLkHL0Ef6w2MwGPXZqOU
xNzI500Wom2d5xt99ddeRbTwbEZNPaz7zhD4Yd+sWoOgRvw0NnBbxqVGdeP4S/LkWTMu+jUJmD7B
wdzG8IDsi6VfFnW4Sx5Q9BST4Zfih0Je0FTUdS6TbcqB0N5R5IzFQ0Vxy7RQfhnfUOCE9olHfkIm
PTHCNgnByDf8zVoNfp6LdnA73Rnnz+znLxGqE4UPk4RHm379mOWRAF8wso16Ve8GVy2/uktCYt+Y
Tu1mokEPvdfNXJwl+/0mx1SXzN8eInjQRLDu4cDwTdw9oU1TZXcqQmlj4wdhaevi5fcv7hBKI7kL
Ko5WSMi/bucxbKbYdZKfs6qSgwPJWkMuA5HLo92DwDpGLFueLjbaELhbFzJwUfZljYXGQrp6BCVN
prj+4j65Pl6P05J6PhoBIP42pUSIJaKFllx6pHkOegUMBbIIcpQ3AZdyvCchdZHXc+5TazcqfzsX
9U7lSgzcgiXga2pWQmFkVBUifIhe2qdnCMwsrQVIR47ZFtnDPYXqA7IQSnzG7W8Ty4blXBooflOs
THT55dtYAi52lHTuKVa1GGIgtfRaQBfh7/TM9Am6L578ECKvBAsmTrE5wBPxQOplRcqUcSEetWBN
ooclIKiZq+XtLAUvTf+seG+v24Xaghtq1c+HhVrQRmoL/ShPunVT3MPkjLfgPjSyI8ZawK9MKU0Z
8hwwP06XClsynSM7uqvzNgy0QjlJNCOAmEehaYdhoZwWqt/YtNWNVffb3WgmNabS7/kDahzP6u5G
0WivFXWodlBpEBacbmm3Si3ZHngbavLDg3/5Rj1EtSPJNx3hmRZpQkGKWx60UETvqrkbeerDFgMt
/E3ZIhLhBmwebQwU26FZxLMWPbinWBxtBhzV4DscuSiHLQgf5IO+CkCJoJspA2JU/2n9/2F1wrf7
Vvw2Xp/WGJXlc4Ew20ojPkya5TY91XeDJosj/QszvCT9l4x0bsz8IMKSVQQxTf1gGNz6U3Eo3dqx
Itft22/J3Z1pCgfUMeNTghPSr9lkp9Ec8jxrvF49fToKYIoukhPbRsnezi0zHQJ8y7TSqt5GepJ9
LNRFZkohK6t+gZ8IVKQgfCTTgQChJ4M4F0eLJ64NDhnXhAwEh4JV28/ygr1Y9IKpCZ7Cqi54d6MI
XdE5Oznl/K0f2Gbl8QItHGXr2nvEWdLc2IPp38ul8pKe04jC2bfqbpRKGD+h4OrUOlXqPRmLR+OT
1sVFd35e5XMjKh5KuFBeOW4NO4NtYH2oAwqALl9zINMuvWXEIPMl3zPX63BMcLXA4RLf4nxoB1+9
XXDdEbkcxylpawhUkXIoH/4GvcdKfamX2dhtY2EVhJ8ypJ5vcOT7IXRMuxV7zIYSO6BLUtKLJJ9s
K8pTgMrcr/R+8WDmgJsR/radlzSucrK9ZRGnKDYC1cNtVM+V42m2f9GjbSttKzTEODBNEOKIDHRq
BuS2LeyXUAWc6TRBGd/hHFVMcpxXi37K9/RaeupS6gSlESZKAEvXDvsy9d2aeIrkU+34dUnHvkeB
cKzBrth6Ot+FyFvE5aV3iKa7mkw52nO5f24JpOJejZMVgczqWlIxu+D6P1CRwOKP0DDKz7yFokd0
b5/ghGNdo+YK4f1feT/KGkRI3h8kVg5/0tszm205yJjBOUrKntSkzdX4wQ6u6NasZ6vNMkg2tEGs
fE7CBjmlplxUrkiVIO5oi7Or8UxbXhL+BUU+2w90/nVbabV3qyWKShIpo6alyCrtOimO15MheWjl
U5qj3gN/HWrwIS5Z3hQaM/TsrM9MtKrKXzxlr15I+0ghi9sPVRi+eA8E5zfrAUmgUlPXs6SdJzSi
v11o+DjcTNcZjH9cDTZ55/ylfTE9xaVAuLFCBomLIzCOqTjsQUeJ4LVng/Lh58IDMua4cfKyY/Ry
5vY0cJ9P0gtSKWEx+2qHU7XrYsSFJl12XzKRhUYrGcchv0JhFDYUwFOVuvvCiU5o0ePjRpaM0bRQ
VgyLKEYuGGwUpU/zwngXiMH9Xi53zCyz2C5nRl61RkNaWj777o6gFgaOw3sU9/hx8TVNioSWKfEC
mm5/KoRfCBq3oC9ZepZjDucUp7kHku1QIQS79W4rOS4rLeGnnTrevpm0XsXuma/4fS/d0FBSLpdZ
0a4CghX/V3Rcpt8f5LZWf7hi8Aob5MNgbR06FFxZZFi53F74PmwSBG2bKh6E6jE+72VkRUu5tKbb
ZOJD5Ynpnm7HSYExQ6jatG/amRqpXovPQESWg5sUEtam0LLPdBeNrGyhe9J0KJcsfut+2SLHJAwL
sQ/9epCW8/nvkoLeZ+JyPay3sabsXlNi1j9F+/GxxcL1w+sp8nmNsqoEAFlu/T4yGoUivCe7Qxys
lWh4lKCDD8H2RoHrU6UQLcy9urAO+atKczj+NbL5YJ2VQLoiTteB6X+vAwAjz0glpKZupLrb0xwe
j56otdvY3yd3UP4e0+TVWTjg2sz2FqCwEOTzvtOjEJ9Cem3EZhJOnRvFLfNNqZwrVSNbespbqFa6
py88C6lSWejTNeS/VrBKRKbBdyLmH516/tszCKDCLbh7pn93HTECNaY2LV/YoLrQMn/FOEIrW25W
6pL3efNGCCVZoPHtFFe3qliueEZbMYbqz01JbtfhB/AjWcoWztavLW8rWLM8+P+j+ZU/qfb2Q6Ty
UeZoZ284axPXfp30VRTmvufI0tJ0H9lUKfqUv8DO6ffvVxGMJ/VJvNhFfqzMgVmzWyWLgXEmTb28
0Tj8pj/WTXIM0izsRn37WNUGXSIacWsOyO52VcwG/QUpxYXrIfXdKb+0YdPVJnlLtwbpTts1xA8n
MZKccc+h2KKofU0TnQY5gSZCtqfWVZZA3sS9a3h0ztBem7hq3g4uj3gkGb0uIL6EpfuwNrygT5St
TV2Xom1USjNujyLn+jne15yR+OXenMxDEZuBrv4Ugv1uU6zSyr8LztBa0/MFzU9Uddcqr2D66hHL
yM744eDmWKKHNom7Q/IlgKkenNkZc7cx7Jy8w6Jq0xWFGanZhp/B+APJPfDemJ5HFCIqSMFNADQm
dDk2Y4P1Euy0PNelc83mB6Um/Jxx7rEXVIj+MEGFUsVM11H8KTD6Kqo5MQxKe+chJfJGLy16JHPT
9FH4/+f22ccc/m3dyB3ULkx4+WQO3Lye/ENKSkwSWXHbFOYKQPybTbLSrh0u0Be/coTvTApvcthu
rAQ9YS62jjHdF8uU4pKcSvxMVgyH89mNRjjzRFhJYSQOPQPnVqFthMEQ4dGNduVFUIZEPlyVyNcz
9WwtTlBlMpP15Koc+sJQMHLD1O/2SXa9md7WlHK9MFij9JzLLRwBBPJcS21aS6sqFC9tVsS00XeO
Y3RHS4sbmd0erOkQTN8ens9FvGqSTBwljC7FOT2DDHaRKh30c1HubCotcdcWa5EU+Iwa63x5MzLZ
Nmq7YWPuNTqyAxINGH2yvsXXWXb1dpHZZx99VK1I1Em54W6yW4+i+6vmKI70CQz592hY7+/M9S4u
PkeMPbyxg74imzH/YTSPVAk+SPhEQmObh3i50fqSCEeac0gexm+eZwOdlmQBc1QH8RdPeHjH9zoc
c2RrF+exGtrYEtnG9TqsvD7VYETNXixoTzuyvkFpXh+GsjegSany4PulVn1gU+xmcvdebviGTtq0
MopMw8oUfMcKu//3SxXSUUVWHp54A50jZSee3MJ4BvVSfDU3FeV5hebT8Uo5jI3fnWEeZgtm23wS
bjvjOpvmBjq9THiJkpV9BM7FS/2SjUzZmCDLpUZjibaME02WgHIH+TZXX27LjQprx4m4CfwKMijr
oC5oRAjbQxH7KIYzS7JqUc+TZd8Rk8K8LQD9OCLrO9EMcny3LG8cph9HSjNyEUH2f0eY+Y8nk+9h
HPpj1QQ3XsYOQ4Z9h7nJOX9awLrGW67SHYZTag5qDIFPjJmllkA6Dj+VRrHiu3UEJpRZFloqBcXv
09IL08BXcy/528RcDySNvvhMzlQnnE0s0EXoIXSnXHvB23gNf4vNGs3opY/MfU2de8SNH6LaE3SQ
hdKIlZRgmIwQqDHWQP8av6IE8ZZf+1BovVKh5hqV4Xsld+dcBjX2V0N+3U1MsVB1RcVuzVl/+35Y
l3CEkHIS72PPjC8JsR8uCWzEjTaV3hI1vp14yka0IU17TAZYke2Q61FJoHe4B9+PnvtIku/lwkM5
gGyy9KQ0YZsSnJ0PXTfxtJE17a80VzQRjhBhQCl48me/zlfI+qVvgImN3/bU0Ph0PpZXN9HLXL8J
U3f3J8axd8O8CEH+QDbNu2UF1WMic/+ESb1hjykURFXXygoMfsAnuTthHso4rnWXR+IcMyzPcA2U
3MCbAVcCQp54ARh3yiBkt44r2HOBS7TwG/iKZHbYgW9mK/5FgI+7aIb5nwwkivCn4TGbXHbh+ZSb
qlSHu23726fzIJ3e8eCojFKMgbpGlGe95eNtrKh6AF4xk00JjmtQhkkO1Vo6BqvIwF623cXW0wU+
p2qD1I8bRgGFWj0xQeKgq9aHCvBab1Sh8KZ5SGlZ6hCrw+MXMDs/YOfzVpWZfhS4nmgr+TdK3KDK
E1N4bXQMfMdk4FK5lo2yQJH2boO0TdVSjTBVIAwNckqgKm+QuldjWT7KkAJt2mfnq5tWv2/vxcVU
EJO9JxH/nGtWvEa7sp/IBovKhvTt/ElbA5LZsdKkWwlUoHlDkFvBiz6RkMV6RPzFb4ML6ndmnE3Y
JWwxGjClAIk5J5+xyVYxiVXpuPSX+jDWMqhEceCie40xiDgtXTSvi7GIY1C7hcLkls28hEdtDhT7
RtWD+kj3iOAnx/1PuWcMDpVeainKdQeOVmlY8cLZ6sljAa0IOPIE+IaJ1WZOq3T6qxfxsFXt8th0
YnVTBbknMkxMOkJmvKrQgaPL2+QjBjqVW0t8QP5NgA8Cz4ZUpa6P9YbVfA1j4Ai9m5Zc0k/l3LN3
Zurc/A0ude5JLQ4WnrIpGslFwj1405AgB6lRUh9D2R4dlRkcDQd+DUVMLrmUZ0XkQKCJOJOfCx8M
xA2aSgTkUcCJ9pFD8bzhOmBi2FLFAfvYi8262p2uCyAdqLpZwe6qQzLpSRAtpJInuYTU0zHw7+1u
EFd1SL6NRvNN11xzhDf8FAI93MaFu+G4ndA7EHKAvpVPR862GvvcxljgCmSj16T4PoVXzYds5aiF
w1RneHdBxtPVV340ORUoQcNx0uFguiFrU59aQCoxy5Zycq+jqFfY+BO8q0u4Qf8sDlTP5jgqkNJ5
b1ypKcUmTFN1zGcE3U6DBX+NW2e0SIPdyTvU2Y/ZzdMc29wnNOcaOTUshIiYb+hXcaQo8Hh0ZwWs
Ux2kbY+ZACZOrmvomS2aCxsIPGIxfhvc8FZN0za8ZwMiy74EXtDn4X51FEwW4k1/f3OtKUI00yv0
SV6XVN+Q/lIB7WGXBIO1vTiu7Jhngwtic0iNVm13aqr1Yn1Lw57HzGLm7eahYySBR2QFKDN1W8bo
OOhB/hDmmTIQCRs27h+sKEIxeJIQzE+c+/mSXA8ya+eiid9yZ4zMiK7dNFZPj4MzRLmWDS4oQcek
hVUoUhmZ8U94naYSoBQq0GyL7ArPUe3AaSBR2LraZhFojOYx/sx4vfhsGpCKERVTLkrC/k0jmglL
Eoe9abdhPx0gHvX1jw4mN16559xWSa/tG2stPEEk/t5eNLxrWWE+iHGlbGAUbYFjMG7z4dF1ucHf
GyTvoiiPq/N/+12R2XRHXo5UsAGWVONh0mDddpFiVhOzAl1baRx5YPNm+utjTBPoYpQZPSqHUIBn
YovZFdHpzJWDVddy4DsHz2vs2K9BWZ5n3shk6thDfDdb11opalRwfX4P8vn3prcGBu1iQMQAEgN/
tKqh4nvDEa3/l+EDTFqp8r3XV8AfBSQC5FkV+NacxGj6EIm28tf51PfgpQMusOvnfftS927f9mV5
1j3b3wthwx7XsMPb4S2tzpm6+dINhlLSN8CSxkiMYD18Es2au7r0umnQgY8rj9AYL2i7ST2fheRV
QAFF7rMaT60bcjo9HDUr0Sfsenf96a1GBb7s0aq1j3UtlstrBp1j5FzYpFrsZOpIiWmUk5V7EhwR
vFOwSY2OTllUj7yNUwHb1QXzv7ObooNHgGX6zxGMdz/vlMp8r9KcDnxmcYOUBb5jNozaaBJew6kk
ZyvjbbMt/Zs5DwQ5MpgPSOCh7pjXvcFJT6Gtd+z54BSkcget0cASpw+07w4piO4Xp3ALwazTGoBT
Fobt64VGudnv1fhZj2d2h+HFT/HluqNthLJNQGxaV7jBgqgkiAs/LBAwSDm/uzooqd9+gVVW1MtB
elyAWWuq/dYYsxF8EypP5ZBrZFELtPAHdhwtAJ82y37IhsQl7fCm9ZMGm0d74HbgWAGQ4n4or34J
CgbNybyGljQv9WLpn0eEmHtARX3NR3ab4D5/2Io6s+oPKMpPHi/K9QrkS4hJIaMZYhbVjwRmBCX6
9BP6HLUFacQAVyJwDblNTmYkBoyQrLoFvNDuxlmsZ5dhddePFGZEh1Qi1uEtfZO4eKm7SbjhHwV3
HN6sxpN3gnLS2Vp2zMsolwqQ9K8c2b18ARJ3/MjkLCxeJvgkKod9fuRqREB39wZgVRUuZKYJvYX2
EHJmpe/HU2FVtXDfYwuB/J8K1CMQUBwAsfNgRSodM5SUxLZx95TGjA0j/G4RuFZajRsFfZffhDl9
hz4GEvp+kRONql98UIVK2ZqpkeguJNyAOiTS6MimR8s2uWFnlktZuCiVX42SWcNTnqUaY28Kywl4
PAo6khTUuvzYb00wU6cguNk6+MPyYNYszXDV9bt7JeiyHI28S31i7hxn/5FUXduI2OdeZ+c0veol
eyL4KPjPWAyBXwBZZ2cBMKGfFCsy7LWvDQei6vlufPIi+5B3KLyxuKVWcZKPxAoDAe9LeN9EnZKI
yOGJDlG7/mZhu9UYaYhb0Z+5JHXuDsykH3f/orfRLtbguMQrakUWxMYbzAbVnt686yj8PLkW2iwg
GuhdJhJp+mjxg4wzMYT1jnKwOhAVq78PREZXID7a99guJuC9h7koCD/qehas9cmAs2m82PurG+w/
g0qM73GNq+MuzbDUD3pZAsnnAsm2TXxfGLDbY7dW/OuBapWX9JOI6D2Nc0EqmQVmtIJjGp0XCEj0
LOURe/8bOm1iPsvL9j3nz7AbcsCEAdSZrUAGIesimcg9hmzxQgTI6lXLPmfm5K3Sox9NKR9bFHJU
mJKhrxLgR5e26UU0SLShf910KCo0pa5/TIYwXXNLVSUMuNno5DvVY0zT1XYXv2IFIQRbBdMXiZb6
ur/OJxz6Vvm5/Z5cwa8yrfwoZza8pG4JqwE4csvwAJ8uR1yoWaa11GubazOne+NYjHqJ9WQkDYdy
USaQmtDdCw+BzTHcAlU46IluwFVgq0ICRj1R1FXexcvdQbNBIdnLXxRn7Y8Co1DBm5sT8E22ZeSW
XQDl2XEwO3CCRVFSKvurSnPaSNQi3oeboBFet6JvKBY2U8iQuZBFsMaImaQdOepgKIWho4rnnXWc
OPt5QD3Mk8abL4Hu+tXMl9Jqfpv359bRMHH6Fk0HK+TwbjRczhBNz+EkZ6SNNtcvjuPckVPozBnZ
QV60bO633qV8uhY5pWntWPp+q1VSX7vPSoJQCHFvkrjVrX/y5YGCP7WpB8QqdiLUB21dD5V+c1+r
+se6eaYpyUjZI+BmBb0556m3iQKt/9IYAbLguTcLd8V+7Z9B/lwV5GaPW/5RPmx+2TFk5kq8c+mg
0aMPCtXv94+R/RQsSIInaKqwerse8gp1wcUaqglZo6wbqnD7zNRH8dXY3fGe3cp+gRC2ykUzzdsr
5jXHZekcPXDQfhH2wmaj3PDh4zDpqPLD4G09pnrxGO6kn+l6w303rcwVhoVgodNWQsFlHEg3I8oj
AlGXX1F45cVXFYmwOHVWvq6BA1gCbzxvX1gXJcypFQwswIpevOUt4gVEWWgDdpsO89Qi8PzOmb0D
x5/0PSDrQX1iphRL0iFxCgkmbTL6ohxURh49kCdQny4thj2c3iQvHX0UFG17Ael5VcfD6Q0/TMBw
DDeFKtAhlkKM4wYmbEq2kqjdsEqCv/sHZ8LADpS2A5CLcjcy9F9hnCjiVQFixXpm2ot+DynXZrx9
Gj4jd6kh7HOg0zAWdNtYjc8yJaTD7eYQGThQs+Yp6pQkJafdurFc5gA+0YQnJeP41J/C/dOwewfg
k0k8QGt2xZscr1ow61VmcuPSL+73UpV7yhRDgEF9OvSaBRF1KAB+KDFxSgT+J9CipJoUnuUGfOvH
pxJmfkxZPbcKSRMqgiQt+VIfFNylClhMxjACpJRYhv6K85dZvlpCkNJQHkAa/ooUT1RTwTm9pqA8
/c+nzR46l2uf07TB2yBlCo1MOKw8St9FSHXKMykqrDFw9G8yHy+v+JhFemADxx1Gsf2wErjel2lb
UaK1LxnPePhEP4D4+daJOGj1tWTWJyuPVWJzx/vfJb0F50ITx55ysXroNUNFQaIk3bQV95lohXtM
N2QWDqSeJjJxT0u169BbOwDuggNGxOUZmDPyN9398sy0CnA59wDecbYnwjxlxDAzA+ulRtua/eNv
pl6Hc82lVULFWKVOJltiO9D6X8m+VPd3di3FkevFP85kSHo3BhpGWZuMxxAhubgPChmFlE/yiKNv
P/sG7WaQyEGLz3K/si/CmLyEn67st45pkqBKSa6D0rsxwznMDnDDjosgIzrzNc1GOjgIpMAtrk8e
bRVU/z+/A5Ugx2oYOjJkk8sBCVbhXtKDTQmedq3IP6u5vXxd+We0UNVIqkvr2/c/5pGPwW8GK5pF
Jv8OjbOrek9o3XBj+u2TE01L3+tP0coWyZSx6ypNjSiVJc54A7WdgXCiFmkNP99mMM26IcwExwNc
viD8yO6VONCqLn/gR+LRnhh9FXhfz4SXDVlmk3wJaaJoNvM8Cs7CF9vEnAN+El0xkx+Qa5lgHa4Q
zg7jLUMR0LwTiak0Co2o8i8PxfgcNF9Rfh8HPXyb3AqANXGhBbJnZbZm9QKUedLOIao9H0mhYA9G
whZ+edGKcbJDQ3bzbgfiiAk68xIHC6SYpv/vRlxzCAu6cDcKAhB6GOIH9i3RJPXykT5ldRszz3Zy
Poez8RD1tIyKu3ByzTceK8hanxP65V0HRGjTAOZXITTAY/pxeL/hcf+RxRWYnX1XWsS0qqHmcIMk
NCMSysO93oeH592abzIxwwhaD1X8b4eZSrul/WXqH6uel/Sk2qOeISItnfm41JAdeYMxqhxj2D0k
T4WKEXAAeNpKsD0EhY/aIqaXkab7xTfKaoJxy+Wu3hZx3TMrgHD6UMxGa68OR1sAaveTbSD2XEJ5
DpZndtpQ8nFsXgcx26dEXEswuNb8l8qNOFfh7VIqhbFYxVedL183dQtcVz5O8mF18mioFQf42uXY
0GTM8gjD1A2lGnFFvCZQ8mrfmybBgHPozIxsbu99Y+OBQuxgBW3iIzDy56HuxCwKhlEvoutFRMfR
u1zgc+XUsVEi9QO+8E0TJ+aDfuHRFOQyvmSwOAHjEvpzBVwQLCjMD+JYa370/mS50x6l4/38y9Of
K/K/7HQSiX+wALZmRzZXZ28ZBiYTzBvMSUcZtRnJc0c7SCa0HVJVtAV8b1t7yiLBGyna8V23OHup
io4S5UcQo8+T+vQF/Mx1Lu/yjgWYGw2VlXmCZVgZ9rm1NaHKfFDXWOGyExl3qvglS2+jYuLhg67O
mSFWP1rE1ATB1lTP5nolh5sz6g7nGI9UgWAwzMxbdVSLZ43XJG8/kMgvnLDetqNzuiGhwEcxTxsV
h09VREGFrk5VGyXdMIQpEgez8/kS/S/DDIH63kQA6muw5VkU7aEa1/A712Q8yUJxpwuOJ+Wl/zcB
q3v96wWlrt4XvH8hXhqjjTIlCul0h0alcFX5joSgYrmUSVf4WxrBBUeKQXXxSdsr81FZk/kEdyz3
0F9J6zZkaGTFZ/u8n6LDQvaNLlyYD56GnKkRjmSbYuPKKoacjL92oYLPKXAxNXeZ+zgp0A8MSEc+
f3KgpL/D2rUA339zkuyHz7n44oAYekP1B7QN8uAYkg2aJa1+maChWWPmMW4T+mF/UDWfW6V60g3E
Yq2oApBKrpIAuj/tPGHQFqu/Ujn54fwFgoLMmhNDs0UAIEq0qVayQqZn6Vv1UvHLfNK0eXhmB4pv
Ey+JWqXj3qqT0ji2zJZOFudhegheRJnGpj7nmG5nXdIMQhJj4TaW4a7QCgbtqBD7tYthG+oEct6i
Ba/x1y1rJIkabA7o2DWjRaLetDhfotTkVeflHx6A8FTskqHyxyaRZ3HV0HccGFbtkm+E9u9ULGL0
KZnHz9j2DLIASPsCNOtXdFLqL//D1seZwDaszwc5XWaq6tLtSGEytIumn+GijAAlqcpOBHBs4Phy
jIyAe4q8tPG3I7rLanu1wm496ycAGIXk2AhTh9g6cdwltw4TOXRGFHMa2W+A+4exCRM41Q/wZgRC
8Vhyj6cG/Zllzno9NhTEa6QIlKJtGkbexthgKe5nJWZJX7gLKuv+xURzqXJScit8wTtNsr0EZFCD
tH6/q757D6/0kuCTd5+1cB6DKBVRL/WQlH2pNRQbLl6rWK3Ug8qBjVTvLWsy55fx7CEx9ERzZoX5
d9ZlGtmkdQA5fepP71Xnj8npRz9NR29WzJsGjzUQ/44DGDJRxKjWlPtHWD8EklgBdeOcabpmJZIW
9idRCN+hNpxjJDdSypH/38T9P/VUrXkzxQjrAuaU7wvC/e68NTOQMx4kUilYlTHW2B3yVO1duLt4
cOEfyarTgFI0Rsw5jvzrxIeZoJDeKkA4DfaR0JTYZTzZCZSEKA88ZlY8hs+8/3K0HAAMb0nFHmmR
+GEIHJoHxBz9drVWAi/OH3ICLh0K5UJ14NeAkZJKE2+XmLyp+biNEdPeIJz7NfTVCpMFC9CtccKE
6m9ff6UyW5DzLJt7gkN7cPDJ7EAgbF2wlS/UPhL1dXPJyuv+OkUSGGRQ+040YMOqFpr6G+3wW431
eYPLmziktd22Yr01ZMmOSkX5Bkv2qIv8sTN6WdfjN1EFDCiXgOV0Qxsnny8BRg7YgSMU85G4TmDA
NcfSzADoe75BXuszQD+rnggLsxf4cVg5dtHIo8XYABwYg1AA9AtKZx1HfuETrIO3PSvoQtipMJ6T
3EdzK2VrsPSXlA44QHPuhRxOn+iAJqPN8op+OZq45u8m5BcUWDVGssooxIhUJeNYgbaqOTXsEAbG
vACjUqDWOJKyEXxDJy7YCZ+VcAPBmF27eY6+YpLh+Vif/07wrQtEYqLwAB3zLMBmOMQAJGDy/MAc
SJULIGnmrikCavlH5x/ci9gur3Xzk3BAMqEypMWfcO5Y8kdsxmRZGsUn5nR94QpzsHUafVZpG+/z
IUuB219zXP1rijRpqOVwK54p1cz77ISy+6GBW/QT3xPTo7OwPYDh/RKTVssuah6ooHyjrJi+aMIa
CZQkPpOYEP4TigIFx4pRFFvMhM5Ayvml22aMRQp1iTJZDABqJRo1uXKEOACVRVHX6Jsy0eJCTTNZ
UlDk0AgHodADtmrRJi70rCWp35nfLhjffJv995kmmEz+gXEzo2lY/xVc+PwVY2E5QpTV4/iU6YPb
M3FJliPcwz9UdF2b9YLUMKGfzP1u55tZqKGrxggkYeV5dI01QbhdRfbrwmpkfBfA5yZh0eKgMAfk
SkD7nUfbrOiMTqforx+FXUgZe3eRtdf+SsHgpIGZPxSp27lWtV7gb6ZMq3rN4iDeRKPSg0I39i1C
9PKBpqZIVXPXP46EYITGoKGwvX27jB19kzqpobkvAVQRUhz9U1Ww3Zn+QjzUp0Qzi56BQQPtMkDX
AcCCa36uDpd/Jm5zjP9sbqnX7dczPbYjNWBZZz48sJ2sV8UvDx0fx6HGqqHUzyU6daIBHjeYQWkP
cVBL2cUUi5fcvxTHb3aOy0MwVFZviur6avr3HI+L/R/SckxL4jXwqtCrZT+k89jlshhNJKA8prYF
o6udWj8lObKCI5y2PHX9IrTsOEcQVQ26YGdDeWdTN4JB0IrYCmy8HmOap6aEqgqLPUR6ihQYscV+
jRE/XL/wP6wlDSHwinDG3s+uVO+JZKTjZfZ3vQVggC/E42bGqFOh/mCVCwjPeGPvTvAED2c+DkiT
IhWWXlAN/4yHY1uGn3CG2TEusP7uRKK+FK6SxsYD5IKqanm84Jri7etFsNjQCa9nOScavnIo16lU
kTLPumN+EO1vkaIxKUliYXUxlSRRjI5SC4+8qUUYvMmHk92uPiNe3Pu6t07G4K7mXq6a6tBWSBzt
hwSMRLWN0rNKwqBKWpFV7VRO0KDRFFcM2A29NwdjfuuR78VZPr9F4Ti9i3pQOH1CbKjuzyLhxPbw
sIyRtFJTOhR0IehCEmU+pDJIslNtXFPhVBapoLgb7EgGGmAB1+KX+53JPSnEfYFjyUseRZz/CK5G
lW4nC90wGXSq+W7extwb3LM5fEOtdjNzrrPKyP0UFtTsgt/3ZTX23lwOL++0KHVWWXiEoDe6U90Y
eD8kUiVdDS9uDobtPGRtvvy2vaJa6TIpAmtB/khbrrnlHFQroBrw9VJKo619r/lNY+Ccg75QQAcc
Iyq74OVZmRxpMQSAqtHYHkTDIQa4TPbaemFhqafG7cLrKxbLvxL5l6TKsr3YXIiIjXJQ8yDpVD1A
ug2rIeN/+ri3zkNzmU5x6zqZSms5xwzTH25T+b1PyoE2p4jPZ4WCSaRzx1WLMJ6NeGP/KE6Nec6n
XiJZYkHiaDh7g2PyVcbAe8S5KNUUuCKPR8aJXBlgYIPKLEdpyyBhTpHV3wmS5yFlVlNrvda3lmWx
UgxjXsH4LxgoWfTIMTt2VFZyy0l1EL/1b9aH0DHyJtv7Tcj4/D0LWuytfEjRqfc4l5KFb31eT2jG
A0IaykdVrkbZo0t77L3Z37nWcEXc+/pQiZ1FsWg4KXBvuC/6o+EN8ONEfyOx80Iv4NekTwbVCnsg
31u2ZZDziDnl+usPLsDCwkRHE1s2PMIOSHB0laNRRzl2Ntrt/oSS5BbtB6pxFPTBOsEBqNJi0ccT
zCIsxmXRThAs56JPe3rHvlqcIKuNkVp4oRF8WcrvG7D8pMtG8zgUo00kkU6K+uaI7z6K70V8GRRJ
RChabUSoLQlEKolIMKZDdvYMbay6DGirW848UBzdoy45cqgTyWzl5MH+WMF5PsicKlMJPhIUo02X
9hS4Dxr4N7hsPLxFMFdmQZY8zZ7WsVZ4a6Tbho6+sPbob8NEatmgFNdW8ziXwieHUhWp91CAB6QD
IkkhGesM/7jsEI5R+e4ZkNUWEeCyrt+WzFBhrkAz79CLbQIg+L7w5x/KIM38ie/RCQQGqnKwPQbQ
fGnaJVllQc2ZgZezrIoJD+yHb1zEL3LBhZ2Y5A6XN3TFfPeNVOPfYWxC9rCeeZ8ife+s7xT5YphU
ZyngnmmeIcH2f8D8LLWZqqZRhcxGZfDjz3uvD52O5xCUPH0JbsR68bGEKuMhgBD93GpG1OD6h2wg
ylbWLUSRPNxvu4GvB/ynmTdhc+OeXtAs0YaoKVHG3C0gQwmVHG0sABc3ETz2VMSNrZ38AJ6l7QXN
zIToZNBOsQvln1vTvETDkRNnNx7W8R4vFs0FENksUGVKBmuyfi0YC8BbJi1CgiyHm1J43jFif23y
ma9Ark4R2XIDIMigOoKnCx98M0ZsWtmt7pqnbT9EDfiXEdtmhDUcPebH5hqH99Fw78HYdspaAsAs
fIr1ZFGcPB/RfdAm1yqWUiaxVax/Liy7Mb5vP47+LOblmqvi8YKe1USXlrOC3tC/B5+RjBzv2At2
omuAMC0WNuNPb3ab0lRaFuSC2sJr13AqHJbhz+mI+9SGULbNhjfAG6oD6KrAhPmLYs8gCirxG5RY
qacvB/yf/J9I5/cBu3RUzZHXsds+7CUauEt4i3OQoznr/UQyw5Tn0duYRzYVG2n9JFk5vrBxG0q1
8iiiFZlPceulrKoPuhXEJ/7heluN2duCXcrLvLi2t83lpkWiM6QQb0qh0mBtVZiXwsQ8GcPdpbEU
6C9czw9NgM6QkYPw4Vs+kPgKsZ+NIbE90hqCxugSWyVGJjAAUZDMJpTLZcwxOAZ1WqauMw3Bkz97
b/rt4DAWah26/iNK+Rt2zims2F/E7xbBEP+NVj9rcFTsuxc90KBDtlxRoe7+ITuNjbRZXMkThjR3
ThWh3QjdqloUjWMmcDcg83zt1ebFdFC9cMZADs+KLB6leZaY+fptwpcP9xUcJBTBQ66cCo0oetdd
FT4bBbuuoGCIfR+7d7R2Ifqgs+1Jf2gQli4Q1mEBQVC7uGqrqG5taAG9Y8uQgKsafjiuRiXMlhOa
b4GBlun9K2UVOfXRizpYYfZZJbuP8xGJB2lqoIN3IeB4FjwTnuSk+u6V9Gl4Cg/k6LhlO67tLUCe
ZRt+xBEU8f/3XNSJbaEwWXjvBtF6PEY628FAwG+hWuQjY8vU+T4KCocSbOpEVaap4mcaZJrviRB6
yJelgCcdajCIPhtTXXbvZSSHpI8pDl8N1cje4kVqD/OBg5X1i2qi9WvspqpDOqfbIFHaY/dm+zv1
93GJZaWQ4WM7hU9tta7PLf3rnwH9yNYNDJzDx+EQmq+HtZGjwmE7MhTeeeK+2psXeMQkbh6szXor
cEYQdFHLvX59H6xMXe31WPMnqH2X6oN+Rc8aVdrlY18fVhDP57Bs7R96QJlaWrhLUTXgJ9P+hF1G
tP0X0aWEqcutGJqK38sn8N0tA2cKGJXODKJmv5V8jA7gKIz1DUdxRq/clsv+u6E6lf/7zsw+lUO1
3mxlnlDTkjFGvHz84qTKMGooCIQAO2tV8UHcVt/L8Q4NDBr02T8EnVQ6nVyqQ+cZsAT2Yj346Pmx
OUg/Ozr+0uoxdJ3RI93t/YbO95o8G7VXaoDA3EFnYzzVINKrIpvj4lM0qVkRoqgRPD+9TYSqN43U
2oszaHhECfWu9bvFwFwIGPQTCGU3mPqC77K83kT7EOODNiQW+qnEy5rcQwmDfZ5KNGv1LejCuzoA
h8k3r8RRqBPtGZdolSIfy7UpqLyLjEIbtbKikuMM3zdGPr1gZU2ka6pgkqQ/lEwItTKmq59WhAtz
zV0l/uqPFDlxNy9KYNeDW5WFpNaiw80FzWDOwMtbTk8ILXEDR9bwClP2lJdf90bDMg2k/SDGC0ht
bne37pPvNzr6vTIzTyEym1ad6LQskTS/m1cnzVPaAV7IzdCHO/huiSkVBXF3GcSROYnvoSUzjCfT
opiZ7YyZv/Yhc8YsZ2XWcY8FgIxPNrY106h1GX6Ocv4ijQK5M/0LzSd//w42D8lsWNjkwOUq+Qhj
dsU/YjpRmehC8+WApPwkW7z0LFzacCmDylopcm2Rlvg4L7rNLuK7QscIJYI0pIBuXYqqLypXMWmT
YzoNBTK35ocBD+vyoWRunl6Pd70PvvlDTzq9AEdS41MbB7huVSMmh/cqLUJj5THsdYKYQYD9rNyX
5duXWHAkTa/cxJG4+7XmQ8xcAl76mhlNT6IseLzHy0JjeKzTI6bseC/gHEnQEOcqRva3YczVuGYJ
SYBpHrEqN+lV8ezxTCoF11IQpMwc8y4BK8r1k7xaYr9EB+OxEBAnpq6IIZ4vAX6AU9v+7+KaFLWo
fbwef0M2sXlAyT0JS21HbPVtp0ZsrMPyhpyM/Wneco+K81s7ohiCRsuX4LUn/LINsxLV2kWO6/Kl
alOyL3YjS7UHBEgRz01+e6MZxg69mLLgfvDMdIpkBmTybOJT5KfC03Aacxty5ucQugRmwGRT+6Oi
UNTHFTa3449tY5U3dd8yZ3rDEbgjTi8ClYMjV2zawY+u5wV016XKi8UR6YoGUFutlV9atM73dV3o
ZPHyAyXu/2AYMPg9meM1avxF5HJfsFYXta4EMej86izTV29T5Ne+KoUDGQE8Gikb/ChT2RbEw4Lc
vine08IqoDYYbVILwO8yORN6ufYKt7QBnSa2k5kyBgQsk4xsyT70rq510SBOOFRc+G5YvexEd9lj
6buqAGmeheDFmtIyCyDnlUEMn56JSxS/xXtZzpD0nsQJErbyM+UdygBqpUxjve9gGJjxzgg4maK2
/eZKclGtMjpe5SJmbuvSUXfFiWvhZRLQDbRb2phZig7FSk70RWhB1CGkHpqVgDTzmA1WFS/tQdaz
Q0yxZF4tknJdn70bHIBoBKEOLnXRbCMwVjcqlfz3L/qnnR/fVdo71qQID9RLHCZ/B9091xP59Bf4
KCeePi6XjUA4Yk7U3jAJ/Dl8P/17YzP1zNzvAcz4tO+Al7d94JQNVdCIo0nm5jRBXxKrC3Dj5azK
a6NA6XdD0V8TwrxPXA1zr/92sa3DEzdEWbemPeZxLcHpdASIietWit9jUdMxKs6AShXexHhgEs4F
nN4uhbVjbFIndWhhZK3kF9sjjMlgkYyhc7qwtXUduw/VjaXL8JyyxvdNAFAkhDohlge2rhN2jG41
NFDQm+MvfE9FipzpZbxNR6s0lzcoV+jbqvHFVa8UhrjCk4ZMHUBO2MSFV4mNrcNabVjhl6EjV941
MPAQt0DxygPSN8Z4qlHlw7zHTtiSJEUEiFW98TcuKqGx9ECPu0d8AoE9JK722dp9CravM0dKWVUS
su9KLOoEogXGot+WvQI6NMuNRGuGkH7B8as8iIYjESpHMS2oaYSf0UQ4KexVzDEtSsNxRg/9G8Op
mQlAT57woZx3bupfohz82VARj/HKyLUNYyiS/lJFBVw2s9rxEwb8luDXAahVRiUc4FpTSSpA0+lg
rWf0kukHP67v+XHGtcA56S4GAU7wn98gXqOLRPfSavqENggwH2AvsaS3pIQl0CTs3y1yeApFGk0U
1I1vRujUrl2virPFx+zU5SCYoQ27GreJoK28/08NXtZtxGA3hsNisLnn5bDMc5BhDmK250U6CE5J
PPpw8jYhfVpyIImmCO4vm8iDFsAEf6x9IuluqKb81eX5he9PQGwiEtRpMFKP0D8SRYXRdSa8WE7I
Fw11SqAHL5nTjXMLBDIJAYAthJZwL+ZqI2J8CG/ueHulFT7GNSYdbJf6DqlgFqHfKd8fQEHa6rE9
sOXPjR9nD+oaHUXOE8YJnnswxsMT4pAirngUgkmzR6jzQrQDzP1Z2YjJjeCgi99JxtgzQmnpohPa
Hv6ZiCzgX/yHiVpuTZJNBGIS2rhr8mNPMbHE3G7Aw1hL9BxPm0zzOEN/3BF8UCwOVn7nUW+Zx7Zg
eEHeL6YJKPpBfaSf22UxNdXJxC7cTg6JvaYFeU5MlO/kROJyM39l8Q9Kwd5+J9qe1KQ+kfRBmQra
K3zINi8KJNqcdoVQAjBkzkXTFyLdjoy7zlPiYsRoRjx77G5B8uqCnhX9ir7v3+gBb+oqwEBGn9kH
PgzO5UgA+aFYB77LRIX9dwGelGlsCsrYs8qY126nscMHPLvTIjPKbre3iCClcZi2zCd07P1qK7+I
KV5E5l7VzrroAWjYb6W/Hh6JlsVLL46rp4ijProYFL9jWrf/0elzIWup4kCwdgKCpqH6B7J10p39
vnDFBRqnkeJ1DQ8W+trDCVuuZ0yoj/U3UGMW5lAOvVSHxguabIXPcCSnR6prxOoKI0OOmublcMwk
OcD2TrUdpsdNJ5La/l+dGA5dcK6we64c45yb3ZpZQd0utu9HrXGw27//KIKsvSaXnQIDCkYNwO4s
sjkONynMd0K2gNcjiQx3gX8qZgI5RY6Xw6Ji4oZqjkuTJHH99zR+I7Dl+CeszdRKZdNgWQNWHukY
qSexYE833lu9wJ3BDBKlGbnyifv6XEJUVKlBWE7gDV7UlbX3MCJ9pvA5C+XygN+BR4hLYaav2yZp
6htz1tTka59OlJCsG4jdRSfzm4s9OS3fvAEJuGqlG+FKB9kASX3Vf3QKHMNkNAnNdFSXC4mVwR0f
QWGy7WtGvowFF6qJwRqRUYVzFl0xgOYtihcWGaqcNR3Ypqpa+SdjUxndBBxPyslHUivE0WvW2Lhl
CORkB7UxsXvwPTRePq4Bkh2LG7ib98rUXCQzzaEy3jkNxTauJvdde98zHajQHEXdK53y82/vJfos
t3DwhE9+jhYehG5CFG9Hc7/2AvacULjj1WyL8/FeUAI0K5RpMwDEslwtRoXzjUxX8k4VnycETlAm
TgUn88WGrmtdOFfgto8HyUB/UkWJVRAYXaNaoG7T15d4q0I9DXRyqgE5xgK7LY5Ctbrtrfu8pUa1
sWuU6j0TAql/xNFXNiBmsNumE8OSHCQG00s7mWa4gTg8HaAiL2IXJ0UVZuXsv3OB8mgcbZCykkXj
LiegF1e2jwTCZ9BDytVzmJ2jyEFiROO69vOWy/r+yOodvnVH8Q6PMctSHqVW96HjljkEKgbQTzny
WWYY74yDycG+P59aBXeH1BqK4EaNA0chYyOrvsSn397/paQ9Q1mi91GW8h1lKFIFBdYjVsYli0RB
PWXHzP2fhrhKj7AKuQ1DtRKPRuJuYoUKFS0BXxRduRHRg4c6vpWy1tUA1vVmkfKlghkygvuzSnWY
kC5PENBC+Ikz8Tuw5soTw8DBz2BSOywZwDbDBmycRKJH/y2qE/NaqHljDsHiqzp5d6N3Fl1nbtzw
tPJattameMvqcelarbuhqu6yaUCGZHZ3iID7CTU1D+69f5jGYpz/SwtyFAVGEjgg/w7oyNvFB5DR
EHqR7ZTXXJzTa5mIt1vt6bSs1l37DrFkEBS1XOsR4Iztj/ndTR2pp3NreqAA7LO/O+DS8vBlCaNf
KEuDxRhKyspuE/sp0lq5paooS4ulh2CdouSIL3JgpbQEXsK5XPayd0fcNW7Ug7whyqKrG8i+zAuD
n/DpwGoTggte29JZ4Om6GLiboYhtqElpy+cCowZt77JPJtkXFXgicfDVl+nfsnYvCOnApWB1mz8d
YkFRc+Bur8qRQCZyNQDnVYm2xBrFr1R9+E4YQfTaziYdJMh7/bQ1gS0aMU26haH9URikDJpRd8w2
cAq1Fne+BERmzEXIrMW6SgizxYQHN9kS2hqp9dNfsQXZAKSy2psVOCJS2+bQOvOZbcAjfFsNh2O4
gA0EmwgRV5Kffwgc5zTAWSk1YTMO1BIwpofUT0blsTMnBZmTfjyKx27FsXahWMH0anvI94Lcryiz
CYpov0oP1AAgIM/xfnrM41PTvHuKvwfICXMHXRaAp3Rd0qYrqHWlV6BEntj/s1X1sVmZZwVxEIRb
4+T4zK8H2/5+lSm2gJouQUJl69WKgctR+SAPM8ZR/jRZXcLQajkzs97/3qc3Yl6knRinogkc+sSt
xJUDAShwKlca2HJadhNMsX4MX/5oo+WSxtCYNG7YC5GCIAMXKspxZV6xttyVIad/igW7j8o9vIA4
EfORJKtwI9IbYDLEiHmJEO6Z3DgA/YpPs6whZLecgupSHeAG++1w+3WI0mEKJTfKCUF32lAZmjCk
O67ahKcmAAKNZBUpEDs5yHR/rv5JElWm1pxLXMWUs2MDEasUCeBHV7HmdSBrtUDmSgnCTAGnLmNX
R0zV77ucNOO+EGIiDtXLIdodlCkUfsCLoUNVw7/l342yo2KhcWjYcjwIoVWp8J9QLG1rLnfnkMip
6JN5TOpFBFod0JHwwwXdl19p6NA58GBBzty3dhK4njVOUKnLLv6wIRmnuh4a5WohSVXayGcGeOW7
MnI3wPVlLhX895dsaGSotKkwHF6pCmI0yEpAS+w/RFzlOx87ZrH/9UrLb/wwJnPiaVosjkNzbvKU
KR9iokBn4GweojfFeeM34I87x19t5/tsk7zOKYdfkigxhiV+DTi6VRIKy8M2s72Zv/cwrsQDtvdf
MAa7quzuviQBH0iMbt3/azAxrwHeYZEfzS9byAxwcQ0OP3+SJMbgtyQF3e9Y7qUjWRH64Hm94mbB
co4TWi1igLYkYWw2rhBfK0HhRQ+5g0XBezBjvOkTiNDCuXHCvOfudBmgtTGMDlvrWMAPUMQfwyR9
tQLvWNP/If0Xhr7Y6ZQiebBgipkL/QJR9DtZeEksRF0Tpffn/2LuTaxUuUi9oUivGlkrnOmGzgvA
JQ8EQOqzm9Q7l6OxKc538SvxMusWzOb5w0LSThRR0fbkQOmT4qd6XgPUguf+h7Za63yhHRT8YwAm
pU1lcqkpa8Du6+Og87UXR8OQCOSSOAp/58gntkStH79UfWkK7tHjMM4+WNL49dMYJCpZxEOMeIo4
a5KpAfIvgHja+oTEMNQgH998rCQMtsrxqLJwkTFxzWBR5ZOwwvrSawtAN7OxAL0CCsZPIvR5gEqj
pfSU7N8G4/dI0Mhhf5AYbF+GZdLWeGq5w4BdydT6MBFK314WZl5BzQvInBdst7WqqaTydzYwYsZT
hKVzGGZevr2118EvQ7TR91U+lZ2wTdcQ2NRbMtxIcXYoq9P6rSUPe824X4M7AxkNYRM/uUc5GS7D
ElaSCelGHv+FNPZ9wLhoeA1y8mvCh5P4rOIZaC3PPf5f9CNEMc9cY/JFb20lTDqweqHK283ay+mM
2n11ibvUeNRy915vQiGsAe0bcQJVn8d7K2+9o+MfSBV8gWLqhTXvI0HzTfprbfd33MhXaAmsNpGp
P16ZEeIxMWIwseXXEW/UoBAP50F45npHRGTL+ZcPwkbGbBSDhbT5eKqu3P0aSoqRTDlz2VLHFw57
D2yoFGLKsv1MwDtxFKX1+RNRNAlrft9yUYJFl8IFTcSJRrgGD8YO9BsTa339qiZP3oPSy22cE5IG
5lrJ6RYpDyWIkABcgpfBa4GHxRP2l8HxmJhpZOL/GY/KZ3t26a78Alc4k7eWXxYvBgupHgu4ZmBL
dFtTYIQMfK6i5Ag6FhKv60f9wt4NmJxgYSbGsWb98+QqQ4KxBg6LdvUcZClICzxbRCpplnNwhpg9
wMeWM3qK5ZAXmSBx7FYitOe3RRqxWhX6n9g0096+sdBsUIB3uDiWXoTQ+LcVnIM1aeA4Tz/1wSGM
yi0u6lSgnSfueOWaF/E2zSnrM7Jyh1X+WRFkh9XOkZOIHYBivVUnNKqDZq18aRJJrmg+ScV4rz0H
+LYGYM/+g62kVTIMihGizFAM+BR8/X1roCysuui5yfHRvhVQRwaHiHnMqkjrHG/jACsS10upDklh
hF1ugTeObNipcGYlgXPaSxZ9ggTVEiBWhKVpPklqUzm/+mSgH0OJIE9ceriQCZftf0fxu+cjQYQp
HP7Z0+L8lIKn7tYWKHlvQZLM766fWN4Z7sphYZuckGkuVtxUICD72c+X08h69qN+o8Y2gInZwZGE
s0hP+biwVP6Y+knfinoWY7ZfQI0ThhAo7PC/OVrPCYh6MiuvV3G9ECCG6S1Xl4/q3yvYReWAolVc
weiUEOQ9RExD1EuLEWx46ZSAvFWyY4yEHQiwlnEXPN/VHZ+2KewThAObS/myNVstEyCQAhxQJkQU
eEgp7GyDa5VSmliCUgsAxRd62/NQ3s45xHlggYAgVuDm8+PN8uLm4DyZ4tcteXMQZ4yk8bBECe6e
oHN+3EUbFrhpH4Rf+CqY5p1VdUthcf32rTw+JDLEqatZlGeuKr+3kTt21VCNZqS08AhKAHethnXS
2Ak66e4ElnZaYu+8YZ8oZFj/icfRiiBM+HeH9GxZkKlgr2cJnWxjzhbAu+63bNJLEebEpdoL+Fud
YHhgsq3ECozqQOARlFxoD97qRchGNH0iySTeOKT+5ZkbJunlBitRHD5oins7rBSsTMXzfC3THqXa
Qz1YZGYi3hq+cQzTICYzMxLS8XdCLHUW3IGYdlSbPFlVNdeX1RDGL/LLCyqaZgVpkFUC3DEOhZnh
+P4qpZr+cy6w2G7P+XmQLGAOSv6StFAHGH2DsFZumH2+/ZnvNDYxtRdgNtsuex4Rz1D45+T2YXAj
Jn6MzJlavoV3JNLTg1nimkSm4PpPyGfiZoplw9S6yPdytjvjL0QOHguwaYSvT3xxBcHWRTMX90i+
sqzVmFizW97yNJnmGOMuTuXoUAwVWqxROLnYs3aVGBoeZX3MhdzMsGfJgcr7NzZENlwN4NGJtMlV
wlWOA7umoQD6ipdatYpcnBbOeMoPjSvIt6b2APFss9Bgy0XGYWH0t9tyRJCTAUbDZFmc2r4aMEsD
ufaWp4Bk6OIBOZpadXOMFfbWts3dQSKHx8C1qzlv32V3LM1HaL3mxd3Wu2A722RK6JUTDegzg7Uu
BOrh0QdjGFFc+XL7p9Hu8BMcUvL85zCQl4QCCzSc+fBq9AN0BhFST/gQnbilFBgHt8QBPEoUAGEz
Bpr48p5ltaLCC/MV+jUtzA1XUqJRnjVKDDeuabTmXn/lRM2walKCpJvS0a1f9aqNnFCR9Bh2vKk0
I9jCFBsFoPnMQfTK/XHKsYp6S/GU+3bqUJWkZmoiA2qAQwqXNI9YaZ67VsbghAjrtsBCXsBVdbtA
VAJvH3ksSiKdU8vPp9GwTl0VK9raJJRSVkCnqq39g9oESbrRauBLQv4N5PveUF9bGuv7WKac7Tzw
FksxOqJlh9LtMueAI0f38C+05Bgo0PfcqXEol9ekwdMHZTXtbYfrcik3QLXISmcHU/VpUh1DoC/O
4sOx1AU6/GYY+2ghNpHSO1glZsitwwSxnuzNqsONJwGhQQgJApScQYEKFfZjFD5HneMVZLp+4oKK
Mp1g8KhPezuX06o8cWIClqZsJCw96l/8MNF3Xrbj6EDORl5yleIPUnbSTer+oRdAL3CWvLZZb7IV
CumVVa/POSDuYe1nJHIlQt85edFEHw8OlBIXF6vQ4QniHS68oGMb4s4aTC+fK0Ys2yegfN+OcEi3
8lDb4/+S9XTMV0kCR10EYXdNVxdPlveElIYbP84r+AhAMZBpBAuEoTsKxVMLjdKsNbpIXH8fDe+0
EzVOA6no+2cQdSgOtV3FCKpgNVtQlCJS/BuD4efus8GgojmFmo+D6Re37OVNAUc4Pku8MXXtb/kJ
K4bGSnjt507YhRHDzYwX6dKxElw3uKGja7ULnuINCXpEN9jFW0/2GruNkuakHLi0RPSoAXQ9j8+e
+ZHjErOzRgk2alA5y8u9CTM26xd8rPE4FDdvr/Pv57ZN/rXGEcCB9Qqk14jGwgD51pAs0Cf2zNDt
84pCPPYW/cW1kvSSCkzTNAq37KjWYADe2s8X8FN/NEeZltvp7bjEePDeneyxjti123fyb9+doyeM
Iklw7meT1TI3ma3nX40lbjbvhGMjRuskY7AAR6hzOR9zAdHZhLRJIGNoAnFZJP60oCFMVu/Mos8i
J3C2QjB5H8Z4IegPWiuQnlz0xLnOl7YBoz7Ylzm3RHg6ThUHvwInJzs8OnnnivmbdnbsXBee6KR4
bsmLDbH8s2xqS8Qjpfvw5dj3qvXpw5yTbhTm6oqXyJMHDd6jyy7D9kjDvQADaULaHmn26tHqH4kC
3Pqw1+i7+iCsW8Qy3wa+yJTkGYCVB2KhS+FngBw5zTu96xXIeh+mEXGeVsaMPO1WFJ6WvkAaMBdm
zqx1Hf101O8uG5ED0mrFdfgVPKoO62OnUeJ1a+MfnaHBCpe/vKhZ0FANR7JMLWGnghg0DLwH9uRN
tF3tNZp1fktv6hcxKBKyFl0fEuvS8Bd8x8vSEM8ja9jvr+WEuY3ZCUsb6z+6mf4GQxRhhqKFOp/p
XfnHgfBeIdTvZjPQjpIvj2Q39ONlgdCSPmewx47Yzk4atS/hO08YumLzaCKLnF2ZbC7HXjndoX3B
DUtUm0hQwv51JiP1HNFdA0EjsfUJIKxy40xSpDuToRN2qXiKR8HX1/OVSe88SrN0aCwoourBRG5t
e6/cswF8tFdkfZA5PeAZpcfl3yDZ2yrL7g2wIzJtCQL/RXol//VTrFAHiNmEPHlZ64jPLGLot4/+
xAY80OE+IMHHRwQHv67Y/qS19YX41ZVtX4jjlsCtAv8K1Gn1nvuQVz7ygZe6Lj8ElhKfVWjAd97/
pjuwgE6bXXRKyAEb9P1lWy21T2kH2DTF+2pSBB+ddLbCtb9dC0QKk0D6r5idCEzJY1IpSceWeyIe
NYK3dIHNzWx6+ZiueO49wnhENHAGouEhyeGKTRb+ndQSfUkayGoNlABa9ZCAGFMu7DbrgfoGxdpC
LjTuJ04iDKHxAQ5Np8nBBI+R5BuaPwJseGGB0oybweiPGzaZtyhppg1XxIi6ZAAceifXlbHbBP0m
tG3C7kmIXjhNqPTFOMY81t9hRt9I5CMHb2mhd9nf2+rcnqXVwoFYWe+PY/Po4LrRf0zmUBcZe2MA
gjb5aXmaIvqFFue838Y5V2etPQSB5kWzYIEwAuJ7D98E4Lj+LxURS6ZDLVSr3KGqjA9M387W8IqJ
UQS+XA8sfUaJBlCuFIbFfGqrZKkJpNWpxKx3Y9fSZOXU98kb1675kI3QfNn6LhKYcI0KVpPzmfH9
cIe78GW7zHXvT8MBamLXAfx5hYss0MF+3M4OLphFYYtMaN33eJ7sNHU7msSOHRpKaW58xXFnEwBv
XqwlGujjqyN4cNKWalVYH/00CuuQYp0da6teqfaLxqMwV5bMHgFp/PxM/LbF3AH2Myh7BsvtKimt
fiKb5kDkIdx5GUjUn3RcwzSRs/tLCJa3E62x/ah2EsRPonGox1w6mBpcPIv7XF8ipGLsRhhdGJsW
pRUvl7c9kXr+Ce5IlvDLYF6mAwClDEq4n1m504zXuJjRq9284n7mr3yKL8v4b3dR+PziCV0VdhU1
cUh5bYotEbY4AOQMcRsgglIIQb39mbso1ee/D44Ov6KoqMBi/jmwu/9jP/o8X4ATkVseFMiCl0T0
+eS4XzXBtCHvdpoeZKdeU8sKzMMfbLdaOzjjXsnkBwuJO/axqaB2daGw/CkJJpH6igBSRbAsjK3g
Izpg/syUiphxJth9tdS6x8DGX9FhXdD5B0qijNIRAnWLNJjnFhPHx3tb8L2m/mTrRBvl6Rxe7x3b
QbdOgk5fSUuLFPkFcEE2SEpoc2dU6gEaHxKpZXM6nD0HT5TgrYB4BY5GO98GvCJBv0zH6hsgqfNk
6aXitP24NebZlJqKXpCkhKEN7EBSN9b7bJ0ZHmfIs9wZcvUbiNTT4deNklZfHG8QAWbmr/QQ+Ysg
A0epV55oBr6eiqZmKmCh9eh3jmzZ6YIplXGfghQX+g2k/kukIGKRW7OmtIHjnePlfucc6t0MR0+i
weKbo0i9hU/r9XULiIpJfZ+ZrgsO7XalQ2CsVvZPTZ7l6Q8g4xULgDUM7CimOd7CBmjHMj9I2eps
cDA2OSH5ShZY+PFD5TmXFlIJcKfgq/KfiZA+aIda4uIxbMpq8Qk8/RohZWKnBpswV3ZIJIv63Bo+
KTipA9bNn/594bpibod+N3vQ56uplFrlgEhVwKCHKqcj3ngK/bT2rVGAAzYN1q8oPHZii12+LiFg
iuYWVW1BJraX9rhjMU8j00BAO9ioKQomSUwTllkrOHqNo0WfvRifvcmSuEZjQbc5EMGwAx2ZvEO1
WFwDaKBk2SCULYR61nSlXNsjge29F+zdG1h0Dri4JNfT9v6Qd7BTU9YQ9WL+C91QblAWwnxsO0YH
gqZG+jU8/t4En846vyc7qmrDEylmRlmUuL/kjQcfwiZVjTicXTgPez19QEVBeCx1uM7QnUg/Sbf2
Ei6/fk5T/6VqrQx78Qh6o8u32KoUtpoEODjMFsrJbgzZe6sL4YsEDi1ofzC+WjAhILJZ4nZGn/zL
0oza4vrCP0tCFJoCCtt8sPJwMK1V5zxJ7D3hThCXgRf+BJWlYIAxMOfLm9V0T/6cdOctop/LtDZP
bT6BXmEIvAulO5ny6XGH+mJDXtzGLxBe9FfCmLT0gDLn9DrmhEg/p9lZmfre+3FOQ2vdbJk3QZJA
LKeT6qSvzA3GjprFoCeme0B5x+oGrIbfN5+EQdDhU0uv0u4+XrGTbL9qfY+z0JjARnPMaqMwUvmt
0wZn7dV6N/fWmJg1i/dbIAmCetjv85MXWS6zGG6f9HTeVPqJtz4esGl+o/XV4P8PVEzx6D+mb0SH
j6BNFHtWC3HElDQwDyCxSindCjS7Xk1orBhRiN7p6YmTdv9E4B6+3zVkSaCVq5BfkEXORL5A4U2H
5lr9VqDJzpiYyeKTczwvEdvkJFkWwHezrDBNJeeBqE+ZNfhfpvdIr/qLn88HRkVnQBNFN0K5Fx+j
kl5B+xz5UJe8nXuQCaLeUfnvmCda2iE8/I0KK1aS56X+nx9wrbKJ1QHyG7+TtRa5L/zYop+6u5th
j2uuE6uBiSIFFOxNm2vAN/Kb6CG3Ti86DJvUF8QFRVZgDVzMWGVXhGDV+cdvGLgzeMtRCw1L+k4L
UoRRRw6lZWNalmMZgPyCTO+jVLFYa2w/k46/0AfKnbP2BvykmyPqmgmbDOiskqYK6yEz31x2pyzR
10EOO15pYP54ALqt7CQ6vdaQVlTo7XSYwv/9T7CgIiv9U7vpGt5BSh7OeGUWs51QJ36ffb6h9+70
rbWOtvSwTN/4L5JrR4CtzGSKZCFmajSmWjhpBpXTh/VFpjQzAa+l2uXDDBtPhEHElqNTG0TalrHg
du4L33ypEHh1hrQIhst7iJ1IYnI6+mSJ3/GM5G7kHT4U1sNF7LVn/72y300BlLnjA27UUWU6DZz0
FbSPuH9lBvubpdSul7YUwWEWGifVXimUin9mSDVoJ4oXAG3z4Z3IhtDdK/4zk+/BCPWu5PsE7vtv
BeQu9rhtxLnxQ5dwtzq4Dtl11UEJoLtHuHpGsPlL3W86730Xr9LFnlYTv1pRBRmgOL0JH7mg7/9Z
XlsPZzyfsf+tmyKMgtAsaI3/TtBF+4hFJQP3mfkCGeRgrrcqX0BTcRtvihJMlZddr+7/MECjlGMK
4Ld26QeolUhwE9JlIz1ovEDYCRh2wd0h2uhraTHl+CzKvVV12JD8y9QFNG5ev5SUFlMZ6vtG46zJ
0R9aQ7SLimJC9bp7WdWTIcG3W8yksb4/lNfJ7qNMEyGAkLqFgq5dwVVQyK6mvbMR+yvauGjHSL7u
UnSm4VSdOn6e7MqHJxKdV0WF8PaqaaWWFjwQbQvN5JV+YTdZbjff9HgFJV1ijC3XUR82rwui2grk
gibNAydN1mmzeIStjCPvgxvwdosFrUgI2f4Hgn9jRnnozBp/yEuZLu+vYVTP+WDaRRBqykF38Fpk
ihBS45DF2gE+pwXYynMJxgxzIcdCKetq/Ovonxy0J/TO14uLSRJi1pSgNT2UINbhqu40XFO4r1OO
xiy+fqKwcbtSG+Pim7Fsw7lDtB8pvyJ83OYlvkxQKGp4AX1tTShtBQPaoRcl3iOvfLGSg5zZO7qu
1sgUJPNIh4o5DtmL5Pf/1Xl+eHmzTAZKXgIm0mQeAVW00LIPXf8sNWTRTIESbdAusntPIcjdlVDA
BJngh73G3EIUBPUmnstxHTTEpO+GTK6Csh+/PgKcbi8IrCle+Aa4S0XQWYvezXwS8tayx/YvUkeY
yGeMbE2k/gS6mLTyXT/8w9h7mtQE4zZhiHGcVinocLEHwbqEesAoZasO3Ngth7v6CyhrXgsazlDP
qeBBqvmpOfJgGTylt+wXpmk0T2VJcOTqCCYsTDiWjXcCVErDgLTkuhNGJYkotV1QApx52kzXZX+b
Ue8YIw8UgNJprZxh6e3F4qN4ODjNOh7b7/7CwlV0jyJzs0ScmmeCsGJAbdyt2CeR63pb+KOY5GaG
UgSs1/f05/rf8lX7n/zpF3N2OhdwNRHcgsE22Dc1HM7sknyOkN/0jE8axQro+oCpbPIzUIZITFYX
u1ZO4h96O4C974vsXa1Nypx5YExt2SIDMN5W2QrMadW6cDXC5KdSl9FL88nyE5e6z/lSGoP0Av7n
r6FJaApmXanzfENqzE95iUEEIgYGqlmy1uTPQIn8zx1px9JBVBHAUWLE9HIfXBhn6cHNCo+s2g3m
/duivwTrLoIdtwVSRwJx9MUmF+WcPKzSyxBAty/AITuC7Sqj4EQ+nWY+vYqI05VvefixB5f0gVur
uCs5emJEugYbae433f/6w/4+Ub7XRdqy4jRVs5nYegDX38yB5XGSx4lyTpcbqEDrnNHWYYAiUuqt
eUepaa/8xf12dVfUBzzUbhJeaGgscAo2n7e6TbqSapY3FFb0YuG1+WyaAfWvxYrn0nCbmV6PJaAe
yhlv0cvSTJAwilpQhPZBVGJxDoxNhOtYXtJV2Z/iZjsjq8yXdHsbyt2JgGi4p0A0PmPsJ6GtIjSb
68tJZ3pCqHAgFVjrvVjvxFY7Z8NpXcCgShuy4bHw1rczGECgh/bFWU7rVOU+tktjXBkbL3vceEVm
cH82OvbDN4MS0RvFhWtFPyIVI+vjef7RPTe98Tq+TcgS5GPgBzQ26YYS2RHv/D37pbgBFbBb+ZaU
mB+BjXCSGaFEyg/Py/Sy9MSiERRYSb9JWelY4PEl6tqI12QH4d1iDjXwAVIV79UdRvI6HGY1zWud
d1yjzwtzvHh6Q3tUTSe5Vv2pSLY/7ixfbIiaup4xtO/0mKToCK6xGpx+ZHVP0fzIFrCQDUV6xmi5
tY6B6ua+lPcFl0MVBIVASDN+8deuOeVvAnyqftyaQFVhpj6kilMaUG2Em5yThUsvJG/VqETrIsjE
Ke0vJuo9TA5fANscrHEVvnzszxLJl+26GUI4qwWj1OHJLA8uzZu6UL7AmBMMZ4/kxXjhRkm/pXB6
AB7rQvDnVLsFghxV88C7Il8dqx0wY21DVn8iandejrNFtWzlBZAp6JeWn0+Oar5h7ORIJ+6O8/Pb
l/SjkIOh97kd28aFOYPlIh5okrVHO4BJ38xbAcdKQRYhKndizxRupunVMoPHgXh2Yz0azEWg/+Fx
8rygXuTKFRAqqDT7Egl+j+4R+GVyMsdlwUz/M65D/0wKhLGLx/4OXyU4FJief+UNgBvyrsjGRjmg
162ZtYLBVuwAiBqiRClyl0wNz9IT3AGknAmPvGnu2Ae2sH4UQJXoU3IcQqflP+81FBP1wEbA9NMp
fnpTvQUTanWwGUaEAL7ZFpj6o8X6iSia+xEFCTbYl/U1riC1KVLqBaBa93Lwl+n4sxF557nFf64S
e1+ct4bbcSXOZccWe6N3uMGNtArMe21cd+rC09SrVwyx66vPJU8zxeTgnI2jBw0dsXmwm2FrB1iC
Mjg/SHp84F1VWNVqJGNyWwkZwBygk0V+s3eNXfwwxb2um9Qh47VDVCzNjgLbyaLzDYuyJQHBs3O8
TZSVvRM1fSaNkLHvU13rKSgzFGqrNSVcolkJmjiL3SbWMJEgF/jNdXV2iDqBTOoBMm1niFc+2LLI
IWoNYtuW6OTZcDQ/wVdvevZFFpEiWBuS4kL09dmNj/wZd+tl+rrRppEQ3bHDZCe22OM6aEnSgq/E
Hlr6WxwvsAtGAOfeOU6bW5BqrjdKpchqBYhEVz8cu70yg8KS2razxMRDZ8s/ge1orGuDu+hpElge
+abGToq/ta5rPOOwHJrG3L49bRB3tYXUC5ujslAUfK7mdtaFMExY1+ctepnwVYIr/F/+5xROrtpU
khhQHyU6gg8nAmyCiQ+JgfP2dNF0FbQT1YqcQp6vgsGo6feFBqC8UghB2dh+0MteJcbPicSUonfU
Qo763oikQSn3EkzLdWBLWdobxkDXSiLQLrkCLeJN7yTHU2xcsSmdDf6lLq4vqZU6TOToe37aQvVC
5TIXdizgHp/rAt143EYLNT9elOAdAxBCCImIy7g6a+X5UT60rmQi3IFGjNZgSUJYvf8ZYushx53M
J//IbTsOfyZGWQlGdd5vm5Tf+YW/R16/TekxtE+PwVXYgeeQbEr93M0IgBQNCTmUZIP5rjMgZMsg
PdgrYTOhdRAtORFN4FFgF3W7xH/qNWLSkIyTApbkta9qwfdlgYRXmEXnnC+iI/eiLD6UgvOu2JXY
S2yk0JeJmrEOJjrHBEXYBMWqWSwuJ4pmpD+QJfVfdJMyYZ9Iy09ySMtN/msypXjLfoGdFHTjZOXW
SCcOXgQcOTEiJnpMqu4yxObYtMuQbs8R/GaCKclEh7RmOGc7iMK1vyNmACTw4hhH2R5Ld3bjb9cE
Auxj1cdlEmz3AuvNk7Fzcs9Uw6hAmpWeRiTMRDgdRxCEGO2+rfAhoL+3Ztt2DhSgqdg/5ad2gCsG
gPaKMzsc9SpiT23nYzycZ+iJg5n3rYtC0Xfv834j/RpsU9QqpRpvGNdfJPp6MgVMDdlpyOopp7Dr
vA7aOx3FaQ1tJw8cGJocaIQOYKq2tsyw4fKtjJKa9tRHo9QDf0Mm699FCiimUTULG6PcIJZtEIN2
hNwOxiGhhCUoLU8UWP5HO8ozN9G40lgKwwWyZD4nrJggZdd1ODIEDZIjB4OYlwpmd/sxeMhAlxBT
bRyTpdNrJlQpd4BTdjKbUAt3kXbpT+RSVtUTtSZ4x8bfGo1+3RSm73cYXf15JaBUlL1q2VWlV6K7
2qJDdmtNaHvXFdl98YYoui3W9QKNRu/YGual2BGLXtnZbJe57ua8ew3WG7zEyY0j04otbPNAcV1b
RBZ/UTxrOwi//Q9/UgdrLK6cNQxM60Jec5yhWjSh+dvp+FqCA1jkxLvuLVOT1JNE71CSLa97aIPV
7MPUEWCs7GheJ9b7NYqHUN1KOQbm+NLiMbcOE34rPlrzOxId+0ww0L6AfI63AgEr40fK7T/ei4FP
SQznlM6BytVzp996KVGdxN1FtCZ3hnsbda62nzbRVaaIKuJkpFn8NFCi/Xv0eU46R3TV93PsYBmX
0Cfum36vmfG8zqHXWr4dTul1TsxI8nGEVW1XKVB1HM0yTbURy72HbfBBTzmxMTRsSUzfmtD2LT1h
szqxeScdXS6cKmJoJtT9SgWQqHT3AjBymTzEdRaLH9Vc1RO7Pf4j0CGUVqsXVGem2xma1+GI+/tC
mqkBy0I5FfPRDhBjAICIDZmcTfEh4lk52Qm/wdSZ/amzlyam2WvUs29SETXtF/uh0K+rP4NVXh8E
ufBKJqmLpHmfti/MvRsOHB2vOaJLNF0rJbTj9w8C4wKbnX1/ihS2gK8x7a5XEW6bniMzOue1hwX5
5uwqXLGFuvfLCs5+Fk902Bfrw4IdWk/jbHNvgs65ifG535aEN8fco0rLdo0pqYiyT1b+wiDjUn+N
4lrJQ6NOXXcWPR36EzouPKQpODNFF523/nhLXjKm7nAS9REC/z9K+StifKVVDlrb6jZsTOOCo/Pm
Ic/QgRgx853uCtIlqUmj65tIB9M2afmmoxbFU7byZVD6nR4XRgNXM+9JAmED4N7Kr8xsWnw641VJ
b4L0PA/2FOjzAuXUDRvoDM9mrVxWn16mIrTXQH8dnm3vULHJTwFnstphW7BUlO3AP7spmi1jrKa7
LkJC2hImpM6AxnqUJLY5/O3JTKvGG+cZBT8/QTzIrwY0EFLS8CTy6zORYJhwzhofYf8YSVrH6JtD
SG3awXxqpkhVeGe9fFpGDSnWGlbNYKS8r06qCBNHEbzSgrX8FOgCv/CZkauELzO/2PfDhBKlmjlR
ZZstdHGl+IQuLefT/V6u9z6uI35S00rMLYR+YAmh2v193nXgYx3MjT14gMwE0B6I0ln1S2VQ42ZW
wyrYBkqRrG8DXu55M0RRKN6He8LJ3D58oHvatvnHqxE71qidTTkNT8qqzFm8cGXhT4QWPHrbgJKF
sOHNWge79kaxhlbKZOoMLCIVtr97CjNuhVjk25qIFRMtdvTopQsfZzBvwCdQ5tqEkZNcWl9QTXUf
1d5lYtVSxNuDHOYHZJAU2/xWghLGYWUuBUaEKbFToMP4ruLNuDweyy7wrWtEdWXeCOde4acIt0xU
RbpZWk0YpVKUCi4kEUrhoZnkiyPrYqGPU85g79wZnrRv4T4K8dSKVBlzUcfVIz7I596JHMpyTNUo
fLSzOREGAJQ9E487KsNHmvceZClmUJF5vYRk87KUqt7+uVSxbtEnapis6ruqTKpR0jsbkx1WX/cG
f/VOi4hmm4Y2g1IWHfGMYyYV83vE/nNDs90vbjbDuGc3y///e4utsTEg0LFAIzFohVS6e5uqexX2
OJrX+Rgs7R44HH4g1y4Y1kD8p1+/58q77EvMmkYSJ0g95PLvKju9L5gKvnJA/Eai1alxjI0Gbw2S
9NV5AvYNq2ZixQCRCaScb4s7pa03smQ15+T6e4Riyj+vAqo9nDt+thHoMpGgYdclZjuBZ47k+Zzm
Dju5OPFwjEBdD4KbPt4M3VpUbgKzTWi6TxLuNXOJh83JwlDBeG7pGmKGGKr4iWVuAVJnXgV87CHV
ipU8S3qNuTURHgN0KDgYvo1ZseYx1pQ0CWSTVybU61SNHgPj67BrySUn6Qw0rfgnZj+ZHs+0X/uU
SEvXMy7aD+s2Tcnlj63RswyxhtOBXnYKjLZCO9AQQrRs37eyDbDzVobaVi0Vos4Pqc2jdRg85NKB
MMFtztizxwaEJcgLzpfFTZMUpYX2enrjyL4kbkcSHDf9h5e32uJxgCqRIBRcW/iz76SOcNM9gvZ5
QYp+QjQuFiCEa/P2rI3q4bTqSdU2H42KPD6FUJAAvgx6idJYzOAdt/IQRYPfww8QmlfU5wi1y05C
YcpSX/iGgmjcLqW3Q9ZMJAzfXGkIDJ1tTxAIvSX9Y0xjG9HjaDNJRIg9v0CxsHMzQA4iB3Z0VONU
mG3UlSM9MZ1mZOmqNHagsxuNHiJBp5bAZMQXqxHAyoMEv6kHhj9MxATXlL5yAczQ3YRscP8WqJ2S
9fJ5C4/Hum2/C8vAOVV/RgdMv4FbPnKuyv4GVk6xDqyoKok+j8XBoQobgnSE4Uay/oIPE9NjVp2f
cM2x3c5lvz2bdBmqJjcFK2wml3i394QvEPnvGjtEb08PLlG1cZDQPSANUkLYdxcH+GlVJbbV5Fxt
EopDfjyelRVs8tG5ivKZJrin9Y8OKalCSXiK5rFcR5GKaqn87Jsjw8DZWXkiLQuBCllUooVmyef1
12CyF7bUgI3mFg7VVTZhFsa1QL5takq3IZXxRqTryqm00Mkc+cNf4B4smZF47XU+OyvzuiIwuww8
RsmLgLM8QMYT39cUYiSnzLQCxXsq/EFAqi8gdP9ZOF/8XAly/n4/V3VlPoQpY8nzIy6jbhFwM1Nv
GzEFnE0mARw4KGXRSomtg646BwOjMz3c771VMGKf+vhyRcgbTT8OKCH4M580AeXSTzbEBVyII1Gf
wGt+bO7PIRYdX3ZVRgO1pR7vdlBsLVjSnpSROLymhOSapCsmiLq8aX/nxF+PQsBLyy6DigmR/i0J
llMBkHXdtu7QsUCG3HLBrtJLZZXJ+0RAquWUJ7UVfRPkikqMM/LoHzAgztSYcbrkBvaPwQHqBYpm
NS/nsMids7R3ud+vd1j1uzJtfObP4zExlRYpWogy4FbI6ttoNdWFOMuvhapTxQA7a+JAvvJ/esSX
TQla565oEbj5L82Qpo3YBgJJ6oqf6AXbswb3vIH45VdU1MLmgU90czAU0QTthPUjHxTsLcW6LDD/
qoB1dWNNIK/OcDGhGsyBHUGBpD2Od3F5nPXYr1gHBJcsHxERAulwfueZshIQfwvkten05psbZ6FV
3UDfk2+wyZ/rOpy4gaq3V0kqOLWJfJdEnjzVMC2RmJmJxOEssV75cCZAkhzWwlJ5JBeahhK3pPr3
V9bMGJ3c0ztZ3FwxJxodJ2/bCDFg66/RXSmqqqJFPuIBTAzP99iAEsrbsO4oK70BNP3Lf/KWa7ej
JgaFemrl5a9TGk6iTNWrE42eN5fEx+bbH7jo60fyKgNh6tat210UM1rEYbzL3qTee1Kmo5c0cOM/
cA9EPPCF5uEmTOXj8N+nX8gehBuMdOTjS6lNhRYklm5BD3NSoiA7IIwLETdRQsBYbXlqX5lCLXDQ
Pn6k5GuJew07oVbHZFyRJin/fQy8ZZuW6RmILmJOXsdkhRNXRJFid673tYuxTxFwzhlmxslV5RQe
zAG+yZPjxMTeB84Wi1ehvri4Md/NHkCnVhLBFKyt73AU2TJnpHQ0SFPbAuWBK5YPPwyhfZuf7FCW
eUb42gW/U+HR3T72KZ48esw52j/ZntFQCSSaPserSBxTU2GmSG+qJXcdxPISKqLS0dUNrfO3VrYz
HUMs+jdqNjnUrwlMV5XN3x3U/0Sjz5IlnvfCm3cjDS7ebQZgmqaOv/6bn1GBXvjyT3lzCIcKfARf
vE0jb8lXUZdaX9qY9YZwFWFAtnprW5lDXNaaRIemU/6S+mO4m/qBDhjD4Dweu8uwPjT+xgnCwZkv
4YnBTUrsvnDGu126er+u0DzMJDohwBQsqrQXCTnSUCNLzWsehFP7iGYQubIopvfBNo46ZVhzqTNf
UxNA9tZ9b/O0SCrjnUriI1iEuSH1NuV+XpGkpcoXc9uMWVil9RiuOnv174SzW3aVY2I6m0m7d4J2
vphowweV0j8dBtUQK+mU5nWc+Qs/h9RWB4OE+AMrpfYUkVCkuP5mXaZSMOdLu6bWeCmgaPeWSrCe
2wqWrVS/g43AT+Rq41xm98xmJlcFUD0YZnGrt+fEYh7svf7DO0zrEBn7hmjqFCJBYMQuIkGz6RZr
Tgm2q8Ws/X5x1y/yhQcMCz2M8OWpF+mL8hCCSTpMs662jGsXc+nfc4U8JYWnyQLVho1PI7ABUXNg
/6F5NteSqkXyX5HAnkHMK7051hGP+iMoTw04OimmuP1TY0J0p6ilujDBpsMNjv2GZOivyOs0Lfhi
SicEzrBxsbimu1WCkXHKVPDLW8Rw9sOGGjRcNS1KsJgkZVvpdTtZBCEMcEkVDRSVAeQvAHqLmdqO
F9jNvUKmr+ocX/3sRu57vLcz6ix33GpTIBtLftuQ0TICxtIU19+tkwFBh3/4K3d0nGZefOtnhxRU
PWCdBQSlq3a/kmQNYoO95ybs/oot/aIXTdJoRzi55/Nj4Dr8cCQLi4AUz7R2r5NeuQ1TG5RzXU3M
vQOcQvH/ck9NJ+7aQz8sF1VZCU8XILufjvNp9GvS8jghG3RfxhXk9rkQ0xTphHS+Yj05LFz0Uthn
It+sgbmXDn18pvwPfqvJeo80dUv8Tp+P/lxlbsH1/1+c7MuOCvbFlQL2/ANJ0NN0Zbkk/xLWwc7p
SdKPzecXi/9uGNjDG1oSb/Zrj89W9sItFUkh4h6i2HH1IqzUpOVszuGnRFCx5fJzykxEUj1YCVSo
wqzvxVgsHxbg0MO6REIspJJUsDT0LQtOWUJztPnl4SEy8RoUkbTkojcyLIecz4YBe+8gv3qj1LG6
NDPpTZt3zyKVm3MHVOFAwJ4AMASbGNOtptOMoBKVvVC5kl3n2bkzZC9CUFx5agO2saLC0p5lLVo5
UuVWeLeUhV7k9WrjTMj14zDNsGfr485S5Q8up799tsO5OEQImuEDl3h4LqrsCfOCzniX4JOBrPwb
VDshjTibyOyvqT6XvrbWjMSBjPq+UakBU2VlckMQFQMRg3WcMEvp31pewG3WW4PQU9aLqBe+YO7y
M5us7dL+ka9PDSCuWiDiEqqx/vSMVjjfaPhj+AG88GOo3PliiV9KmqlPtE3GxRGcbFBaLQYeUbr0
QNEPoaCCXWqwGHM/50svb9cZ5QDiljSNYhXP2QSBUaqH55imzYjrtNTzy6hbkE6L+qegKaIewXWJ
kx+4ftzTKdfFHJ+Wb6rbvxsTf9NHiy7YxTDfdGGDpKi6oIwhkPLYabzNy9ttjBP3MeaJ7fe4i7vE
EuitcPjX2+s+MdLpEk6TbYlpShj+U3dBA1ChFfwtsurHejZpbTKxD+zXFpd2ztVokBLhkNE5Cb9+
FzE2trB8m18/kWG09reqia3+shtEdg5WaigPkd7jjWv/VYNKS1p/ias6LMVGyIxUP6ay92qR2KXK
QydT6v++iKEofoDXKWFDSxaqFDmhB3IYfDa79hKaqQaFS8Wa1DyjZTung/vPXOxJD5S5DOsBN5x1
a75IQ78+ttQkzmWQI6YFd2QvCaFIKqZ88d4Tjsh+MjmymVinqJcR0EpxQzxrBuw2ISQ9vvTtGcD1
3stopjmVPWSA83JPMsGJ3nBA8bGDlEGXBYldZ9yRJi4bNpzJMZWTFhWLwYYERXsowYVQ9RQD0cFr
Hwynns2fhh2XQ7v1tUUukyRp0yFNmulJ20VEdTlyuT2uJzbtF0MGGl8GXV9WViDKrzAoFuBH/wAK
MLFKFB0IqEVIGw/SQGfqDdr9YxamNqn9AJvDlEk55IHMSy6JVrL0E3vwmD92vmpPqgizPrdSXQRC
SeLa3W9+cqvEEevcaQVgc4fdFewf7OIKRKR5F/MDVLt3B8KlHRnMfA2uxay7peah4DzudUZTAwS7
YbzWzOU7//7laZPaHlt9UmXnnyEZ8hp2y58OkLFVU0AgFgLwjguTPn7waF2DyLY8NJ/mbprD3f7v
GJDac9cQo8P29T09J//MDwe6e92x5eoh1QYlWHdJWepCzp5bCUWkfGlK2N6w83IiovQW/hPu09hQ
GhKoVLiyJ+/aamMStkZO0WGIJBvUAaw6M+NPczQk9Ph3ZvCocQh9ZV7n6SVwSmu7Z+dIF3UcgYBN
f8l7znnWiD1iiYGtdMu1ZMZM2Q3LuWDEaIE8XNlqeNSlmvRWEllJbbxPRrBt/wYtXQUWQ+Fy35Rz
boDF2whjCH6KDMH3szeLLjeg6039VizzpFDSSxzJGehUNdtqRxGqbGFummEOduk7QKFmCZTDHCRv
XslRi9aw+v23nP3C4p8wtLgM7//mCXxfhHmWusHbj1qnnkM1wlO4VlrpNUC+gVKvucLmpQ7BWNqn
IHadwJayS5IzAyHqRZBgKKMIuZuktab/2cLsBd/Mr2m4dSNArpjqzIur5qSzU4MjLVe6HvC9xZ2S
5YbmzLwZlOuFAP4Dh42bXKUL7hqzFGOkZ5DY6E7mM5ivUT9lxCN7RupBFIN31aXGlFKp8MUA3gCf
JZzIrivvWZPsxCPvkk47k9kZZJAesXaWXge4dkh+rWTzQ5ywKTrcbnj5XsTiFaf8cNQUhdvGcplZ
HvaJquOVDgVGj0D4sd2odJ07EFw9CKz31oZTzzglPRChOBZHGBM5cPDIyb0IhY/msAuCvKwU0mvk
dtW6QJrOz61klJwy3UrUyMafMAHYELymFog+ODZMhBpZNwGzNnK/w7rvLbUf3rILx6OzSikTZWvQ
7qlHJY18CIXft0mSGxgB5T3PUMsCJW+GfHjBtkQQDexMplLBvD2axOYmQdrQKtoj8xjXpzIFCPYj
auZzh06lpxPM1zp49pPuHhZVaowiBA+WJYIl9WazPVZCyrvYP+VPL1AZKiK0pYJ3AcpqMcg4nC5S
AR7bctjk91GqJxOa9eUsBVZGRxGFrXRKK/l71f9ZTChagff8G7yuE5iloKUHcMkI5q5CazwaIvJl
8m7VSh4EFc95//wqWkFZFr8xtEFd4ehN2tvJphyy1Q0h0u42tde9FDWWrDf6O5aaBvguzRiItvnO
73Q2rVgRxu06P48JV/Iurmr2IhNtlbIoxk/hj9BjmyINCKBrWjikigUj/MnaJARcZnOyWii3Ymfj
mLeG0JU9AutTeOvFjHVh2Soj19ydjfILXaLWsxzbEQHjQC3PGyg3EwsvSV1EG9oVVlaD3OVKXmfA
AIMOeHzRtUzS9cU3pcM58BT851mazy7TljdBfZkERZaE68e39xwkMI5YR8bjLyxkoHUXhUxhWkMz
pbWhy7/jWOtyxW5nxlThBd/nrUI9mpDmvOaEG2MU9YwFHvxNwGkT3OTUeR67IEQRT2Rj3IHzEL+c
HXBYz9VTOzvBvQyKYOPAbbg2XJnxluwDuZPV6x6yJT8EPBpU3LOn6v/sjIQfogBKre8w20qUv8Ro
2Xa4/IV3lPfO2C3qzCs3hfBtzihBxOj63ptAm1xQc9sglO/sbXeXikjsxYExTtf+D71+hFZ7swf9
Y++acWnObOk85TLH4HBPCjZCWgIx3wfZY7SVtJkMD/KHuz/s9I8atoFwI1PZiDGgKipGG28fm7MU
xo6umfMPOg/iF74wKeashsjpO5psoR0TRuluE526CsT5GhiqcupdH/y4raGEhoCWl87INA6dIbtP
JwZrywW5VJi47DfWYzFKwn7oO9w8/HXzg96NRBmT/hTVpukq821dbpwnfDbK0pqEfvmexcQQpQVI
xSCvOxLicHePQXI5D4Nj8VuNSW9hWOMuXmtRYnpvlHnPDHIzs9eYpRp3tegO1xhVXhEsxcfZk/Lf
mwbyHR0AsSsNTHoClpf0rhhBX0ISNeFnUTCi+0VGnrKUC1N60R8aIoaYFzYPbdf+ifdaq0jPmuIb
nm4RnCScTJY4EdIPXaZV0I8ulLhLRsIAwEVL2rXR2bnzu84eWcH7tZ/70RVJK8ws5sRIl0j4YCIa
t5ZHsXQVH3FqSjpE0gcdJpXOcKmNE6iWjD9JSwUo2LY31o8SDTEzKR+PaN0yt2w80jr2rwIpkbwf
ZLGNgrBcfPyuncpGcR9nEkZsx8+xSY/QvTTuCmDoPLaiTC99b+gi/I45GSmhsPzUiaWQAWarWWWg
BVCsZykl+n7V5/ohg6HJxFmWwNiKamgBvb5dZKDKjup2DuwuHhpXb+eOmrg9U8hZWDWsIeeSwsCV
PxQC24CDXVgZwHYYytUbrfRx8CA3gtdr3fRMwRCe0rIqRNqaCpIj5dS7+yeps9ebMg763aZ1bQTH
RiJIBoXeOWUEL9AWpW3RatEmYZkXFZaGjOoKfjv0ptIafOCOaGd9SyhYrXv2um1MVspedW6lTaHD
vBfQlwY0yMi38Ki/fdtk82EZNn4CNDtwoyDnkELSvqNRhrAxXiWLeCqpqyXa7kHx40WsrH8wpkqp
3ZpgnUebUyAYe7u31wY4ej3bvBqHNFWuRq18lHttE16uQW4R2a+/4Btx+5x/wNndeUUV3A14X3c8
uTLv2RCsIJBl4VmYKMmoKH5DVU6DhwSj+fwXhEz/eJE7B9Ms/mi4EO4VW0AKBezbh2ktL7c9RtsN
r8cuOboINdia0hvUa6kmikVfppqA8R7inNWIF8/0ITgSa761DGlMnZWaP/TBBwyFbQQ9FcH8H/yw
b9cKIaTy+oUbiEYQQHBNG2cPawhUea1kUSJLBCTcDSynJn/qIE9XpGgzNmXU9ZCR+BHAd2JZebq1
BH3pEt024V5MgTQ548rXwp5oyF7aP1OPjWAolW3O8Il+2CUtIadGD3mLjitlozyfpya+DQaEkRKt
O/ZlaoY3W1aCc0Thh9tne/EzkPqUeggoCwHDUlsW0Xg7JPwsaEzMjOO8h+vuuyxjacjSslZMYhrL
UV0YnMqSIp9yGeTVyTCqWjYQmtUlyQCB6g6V8w4uoKVfZjcQvtFc3rOHDklHl2EozkX6UPYZp8KT
ydPwerKT+HtNG9pyYzSxINYMnXyrmAEA4J/g911Bcg8yQidm1i9FzaLILGc/0gWiG1XDkube1XeN
/TA8S1xrNC2p/JkA0ZhntZcp6kh4SaYl9cc5iRkDsTB87hVXWunHqrbVunnqPixcHJ+86bFg5q/r
eC4jK/pEis14T3/lfrHQ2rzXN7hv8+qqtbJQxooRq2W9r4vPdfdjQQkS5VhoLq60gWVHC/9383gM
0wmg8GAvlMR/e5kWikuP6ykwP2Hdtva/DgiDnE7N1g+9/Hr/fnIc25NXaz9UaV732n1bQhvmfNE7
OipiG/hJQQmQW1866/YXLlz71rhaVlF23VbQ+/t//uP1CJWd7L1YNCLZXH9OvPdQdEei8EUVT+D/
csiTwlgleKNdp7Iq14Cf06i1pyN7DFOkkub4RyBLDqV/pDGsyTCBsg8MiP6R5kMlScX6BtqroYb+
wwfg+vVMDc7Ypaax5fhES8u+d6apKncziwmSh8P1xcQkGsAdR5YtwRqiKSzId7FITvYvXfTSYzw4
qNyZVkytXUIa1HVTtVgu2OiykFuHGDI9U0SO7kpqkHTq4eLoAU0At4C4adpHqX++nu2DlYqPy2hv
oJkw4iUvOQ/HbRymAyJq/ChrwJyIemTPnto8kDdqFjqj2uD1Lj7GOuvKbjbRZYplNB1uEHAshjcH
iz4TaWh1KEoAsPcqiwHENMaTeejszFNYG5wCD82+ZGxMq+zSe8FZfZ/SbME1x/nCHZ0RlwEiLLUi
z/47voXWd5sM7d4xt2uIy0A063TAX+MacZPEpQBi7Khn6spmvUNrPv9tnafhGP82UckBt4fH/atq
ya22qM0I/+6n6/psj+tiHG5fLEO/qgBSWiCNR6IS+bTfAvPAGo8GDWIrsq1TVSyuXu1oDRkHui/L
53YAkPXzaDIeynKFPUfPyw5or/Q+92nVnLNwCdVH5UGhT4TTUrdrI3a1+iHdnfr6S8nhPBbY0bKd
/iIKgUbu5fLE3wTfMCxt6kL6enLhCeeopfVauvb+pxxFOlRiZoLcRwoHzQgq0CSHmHPBwzriG4O9
PZuhiIwhKBS9TXk4oAqmZepNJ4uVa3R5LzNsenbcXYlSTFjP/nHN/Fk/09Jm7NpryWiObUECjSz0
AMOGLaZvunykxYf/Ot2tUpB53v4hFT71C5nLMOJNcOX+g2OamJCfIpceJQ1zaDctoYOtPxGU8lZX
Ox51meTTscQB9cs1v3v6MpJKlTSjzCt3q6vJDv3O81Rz8hgpVStVpxMU3oJ6GbsFySJjWWJFFp+s
M+7H3etV4SI+0glJbuYJfl8kClR9CwvlqekHcMrLadEfiy6YjzUNDeUu96oPVg0i/mEZ4Z7CozIF
vG/rUiAh/1GHshSuYoWJsr8h5xsDst5awrXjO6G7X1RvohKBFL2LtX8UIYe2xbAxQwVUCbsZwLsO
aUiECaiUdBn75Mxcm3rXC7BdFNSmllcyODO0DIbDckc6oLY+EOGBJ8y1vEIi9OjbOdnOIereZUQX
K0Tb5XNyMdxElgEnHFcgfcXSs+yj0Ho6gSR/X0D85ymeMJ7NAR+KJw09IUe4dEF7Lqq+0FYHEKNm
FmSxd73wK12BaQV/ULyKZpXuI3+NwTpnpBXx++RkuAdY9C/GjEgTjf7IJx33lWY7CL+fygOXX/WG
EN096cbcC2erZtL/3NkcE3lzPtd3m6hSrsHi0ESy39FUHZCjX3Z6KfiRUA6K9715J9AVzk9qFkbZ
fXgAA6HjXXNZweLCG8DhMc5wNOHURjLhMWSkB0KhX+ZrH495InlbfVOWmLBYuplDLM5M7nG7Xpvu
dYcpQ0B8DDJzf4PYX4g90SprjXz2r2yEotgacSChscYD8/22frOfxwFhMzjKUG10CHMVIZt4w7Em
LMlai8JW5rGWobYNMiXKznFWs+fcROggZiGjlG9eFEp4Zz+iyoC9QQXVkDo5nNDGJtffWfwOb93N
VsWVanFBRoZLhS5Vy3W67BUh7+u7lif0dWlwFPsVBPbUVACJef7lPHtI6+57xE9E/p7phJzzCo2q
VW1VcC/unK+h9GA7abXNIEG1i6VOxJrfsl1+RLSLPCwY4J2VHnyZYomd7wcPaxwanVPNusSjdEzS
FvQ2xkZDVrzpKD70vqf7AC8PHrWF+Z2kOkXn3YQh2RmGytqfvtiJv9qvW0xsmAsUBqiLAi1Ww0AZ
Ufdbf2UPAGS6yYHJfBlzKj4akLV9H8XTy3FXQ1SYgyotEr6DgjM9OHdw4RI3w+RMYAZTyWGhqTZC
a8EC6GBX2xJC9Z1glCIqInztO3EVJhJZEaKFJFlX60xP8nsSLs3LpLhTwGyAyt1pGNXofZGcuxen
fasuzcQPp8Pj3WcNM7qt+v7fHJ3H+iVAN5+TqTg2t2ge/oYVZeHD3WXytD+/Xt2nmDUR5JPZD5S+
rAQyk4LcJSVhfzAacSzGnLdCDghdlJT0b/QpH3fBp/tQ1D2+ikGcAkiuqvDOdVeo2ugE2HmVyfNg
GOn8XjdLe9fLM3w9GR30ddh7b8Y3aBGmELv0FOV/7FK87TECfIUmaSyXzA1d1P7qcIx4F2vP5Gmo
uyDzgbURyEiPS9xAaiD+WZDa1heD7lHqhF3+mXN4WGqxj3ExXOfT2AntpoDmSdbPMT5qngQzQ46C
HagjoCcpxJWyP6y4HbfRF9JuTsUCbL7mTVQExuRofwW+cGzzK2zWSrGZVTsDJWAzpH8zMNMXW7g7
czokhzAaUqgPHJTMso5hydGu3ky5fOfKTHLtexDxqnIbwcLFnQnT0j42p34BUzhF7RoLiPbxj39f
i+iizmL9YB/QLh95h50wDOTA+4J/8fBk+nKsy318Vq0mIUh4ri8K8wvESS9d/y14/aRBjp2urJ6V
62+gzP4vkho8LVpVdiDYVznJofMxuo30LREAimKigF+EhXLwmRjEDsIWKj7Y5AzJPJ6TkNw5rDhJ
Tgu7vB+i+nwhl5sAaPblrCYIPv6xRDVdQsnBAPvppe4LysyfnEe3TWtYD5KlTMIYWz1SSxEwDOWW
vQEFEa/9pqkO0eNBmbf3VOIdQFnCJXHrwmLp4Wg0A96dqUEJt3cZpcPVf5tR1Bin3pAaVopeTWpv
/1jtgr3MG5UrmFF1STEOsoVnNN74tavtb5BPOzjOg7Ie+NGcLWVund8ythAkBnxB2OOirdXHVhuq
yBH6Z5ivWYe46H4UK8HPvTIiM+mOwv1PkdIi8oKHQEOkP8H5nVZj+atJuns53EU46HMXuLtUJ5TA
eL75k9KSsl5djs2Jsrsg55IKgahd27OnGT85m9kkvPG/qnQlmH3DmLO7OOv4JgbgyqJ44Br39vqN
0Yr08NLk+4Rnhrs3gqEvGpaGOJ7VQIxS6qAJhn/spikYfVtUcCczL8m+ZRBUP7+tsssXXfLqxJUQ
KMmN5jo+fkMCCOoC01Af60+pHFG0vh+BdRJrXhfJYB/T6gT9vQkbQTB3ziyYFbh+dxNpLmoyeBWx
l77rZeqe/63GMJA2vsHRy/mErX0VDlicr+C07Vx4KKM+Y+I5dI7lALGVO84kJvrlj3nsqFomt3NH
xSU1k4qdWZ1CHbXQAa1Ye1mnsm0cDYkkwUjvbIrMH7bXz4mYDK2w6LIPH0e9wdaxaiQZHjvo9uRP
pulXXffa0yuCuo0AOl4w9jkbr76lcKNWVkz/ycStiqhHAIwm4PjasP6EwAy9vUD2BHLHUhh+hy7j
RZ4fppYx9pbzBEMt673yTAypRoynwfsDtc4BgtC8aS7tqylapHiaQVDQRl87IaKbSFFrdpzcUW2f
dsAPJX4lNMXB6BU0yXDiM0ujzyQYIj4+vOilwqq9k0r0iUDbTn7oMk4qjIO2xUwHp7qqu5ivHJcj
nPEGdTSqVM48pDWOSV5PvsUJyB/8z7xgCuRNB8GIj3Ry40yP0EhIgpMYFme2UPvTw26eNiG6xTBw
8WVzrrCpgv/NVf91C/hFDEX0Xb6eQmt+52eenYkk6CcoD9FhPsKEmnOy5oX0FHYbD4gd6OnGBGGo
2a7Y+5uX/E6yvebh3m9je8XfYyeslzqW8PcmgGml7HBn358PovzdCqxfNXd3HVf/vvVTvwBvLBqN
GXS9xgQzfdMt2Qv8EQCflAUzXwVT0d3QOAz0uQfIeip5glKtbWRUveTdJFFYBK4k3fWO20Tjqelh
o5Muva6y9k8y19xuKNBFU2UPGsj1W8j/hpRX1yYZQuHXz26hR+Z6Oso9CND78pUKhgkzliusvzbN
uMgrcZh7EOs7JA2tWASpZDW1qjJHK09kdXIZYzxpGBPe8Izi9q0GzEVwioMMJpDVfIi1s/HPTj5u
icPxL6bQYkLON9VlGOB0Abw41ff6/XALtDTkGJPgQh/xL9g2MuHzYnp4suUbWacbfU6BdRaGjROq
zbRFMikCDtFzAUsX7DGpyV9Zq2HulNztuk7AIHqFmVAZ9eSKyIrM9a/8RF5DWNBYTVO1aluPBhmj
jzG0BlMtyIxzHvj793Oo/fbdxkLNSNtVeQUh96tJUGCJXUw+KPaM9qhaqGUfHNfIwPry3J9Zv5jc
v3K0kyFtH7AinkNdJ1An6ROlsvGzFIBw/qZHFq4ht95NT+cOumaPziFBGPlqzHiH73hvcXHRtOOA
g3P7qs/NDCa/zVmH3m6K83KgMw8xiZ869ADSOUA9tjgPmCt8F/ngq/eSe4V3WaWUmu21IRPT/6hf
ZWExecqwWLKU2Bwwdn0RvJhREXbeZnejZUD+6NqlKMFUwvnTiGehGfyj1o9QzLrXSn/UIGtcF4Ch
gFKOjFz53Vpx1QQ2Cueyfwnyo3/rCI1+4rItXaccFVLwRQrrYvbs9QGIYNbToCCwenRa4Nj2ZEWT
39Cci3EKQOfYNQyUYIEltV2qoNILZNs8jsokc/5T+hDft10QqDJfBeC8622ZJh6VRzIGo4b2F3al
zUjSlPLZMAOhRrLzdSMIBW20dGcjCxVK5UFCBnguvaeLLTHf4KzCBIe55Si3ZisouMbCHViHywa0
Cr/PTakLNYfv6XDE64fdaTiXdibeNh3ZO9PJMM26SkCu6x1ZMHqkmMyFNpFMrT2oiCqMMUINJNE8
UF4RuAgKGlJJdUfI36tcn/UuOPkrKWemirywpCkIIB+mlRUCboM4uK1b7xFk2NZXT5hVnyjtoRAa
t+5COad8ztDFYqi4NI2k3GT1Ejihxoc0qqNfwAsovlnv1W6WGvOiDK9zE3e8r3Fu//aOuYsR+yUf
Fuy7cdQanLGfY4CDqJwtB6XPfnOaOoz5j3xvb5b4i8o/SWjhW23E3UmglBW5II4KZxd+P7gccMbh
TmxRTIcl4iHyAUUq5eDlpSX2apb0nYv8+kpgHIv2FuaBFv/7ntxkQ9AIvDYpku9e/xoMaoVj7VZD
ixeUixa1ZKuC5J8yyEZo1tORhMvJw+kj7kSFZi33t87d59rtM7YPBxhPDWKCMCbmmj1+vFZDb7S/
b8kDu04SReHzopl1jihM9IDtfgVIgFRWHCQRc4kl6jQMZ3rENZRt58I44ckd98e3K7qRsc5EPDcc
eYscLISvYQRnUc2Vtwz6xtgffPIwf/ubfSgpd83+NhpX2UYBekTXsLaJtPxm0XPiu5RxWBHNeeIr
8DskRGnOu5u2P/nxf5G/OTROu+im5JdCjJ+H3CAf2AzvJneZT/A43w42/Tr8LQvVOqeCrZ/C0pTv
M894AHo1KM1XBVdHi8EwL1VKjtCmV/ba+W4d+VnQRA4c7kOzaGRPRuHuva6VUM/pDjlbFHtRW7Dy
RsH6Q6YnqhifhaMrpACXQmGuo1JoXrmMV0bk2VFhXIedS+2/S6tx7rSvMlg1hgoSIzMS9l6ScJ+S
peWwAyukB2DzvZ6ejltWXMQdvyCMbFlkVxCdzbDiQlBweuVApMMqEOXeX3nkO1BEoElz98lh1+3a
zqejCzqD5ob8wiPFCXzYieuiPnajinvrcaQ2pOktpLKLbvhDc7M4Y3UcXqKNG96i9tjTpkSaIAUu
cmOo+IYWhsqYy7wPFEeYDrWPhHEjhQDRuTqQZcpbbwBThJkYk+oRm7v7xkIlgu/gQbPhomEA8gGg
pZVRUuAceg1DZRpJiWDDcyCHheosZzh00QcGmY2wkyihXliWmAy/YfY3JWeasBTMHCCYlfTS2kC0
fbBXLgQqQel9m2AkDJ4ts0priPMaugifAPVEB/YSphuGX2hygwCZjgcOpeCoSE+yVrv6Rd1ACSwq
FPrejGWtDamIwJ5fzvbD1dji/Sg5jKOsDWk/p6LdZwLJig01Ch3goWdEava1wQ4qixnABV7swy4v
/bF5eWJZLEK+Bd8a9npAHujkI8KwIiOLDZK5/JqgR3ZlyPMP0Fp4ZEixzIanWqgNb1OIEJf1I71o
GXF1NBsSwaSgthvQYyGNKDVxmsL2sq5JN05eLnBefEAaCEW5kgNk1Yk95y65Mhs1B4u8VadBUP99
Am9kVv06JV2p1N55qNtyWxdTrc6sSJ9z1IUH6YRcTQB52SOgxhHvE8Rzbh+5/QwDo/SU/WsycGpp
iI1wQji78voJ+gmTJyK2hH6Dw8ISnarGlRQsYEwenC8V2zPaN/ENuDn3YujNylrWwSiAE8XzyE2J
yB+MMNtdTIm8QWomIUG+Ew01oLRtOeFxd0RxER5Ng2cQNOJJ0kCvWUI0owqWhWWmNNqfwa+LsICd
CzipUjW2Pz8eWFhZ48uR6+kZdUE0gNKf1Ibckya+uuoY/nc/zdrwrcNEt+ft2J98wi0bU+N0e+t4
tiRF+NwhVBOctmR3g3DEqBhhDeIFvS7EycHTRqgjfr9RVnzswK+ZyABcu0LEfymAWhtfZxRGMJqu
9j/T+P+Slotil3VeEywm3063qyh20x7R1C0bJS1fwxhDFYw8qO0DoGAp8Qo+DYCWOY5/6xG5Bt/D
WZ5G1p68bAMQVL7Ow7eNE4e+e+KRIN1FalLY4zXgxbnI4SJYedPCJhPw7CKQz9PR+LYKTm4is4pc
+HPNB356QctPiUjrWk7IZzBl0R1UCa/Wz9l63jdTxuJBRN2GHXPYWG4/tKhtDre2thjVQeu9pk0W
6lOx+pki8T+Kbm3b6wwASyphILBDCmJi6jQiinaxU3KcNFp8Dt0XxozcDdjGrKW1kJdKo/ahoN/U
VGgeCXIv9CgPqu0K5qqMmU7TTr0lWvcvg6FUgvnE+q6GQwkA9Z/zt/tTyAdvMgEno0XwWnmx54xq
4MmRHr8xWBen5T6CYcWSqJSmu3Hf5b5n9CmvLiRyH51sr+WGqEaIIWKMTtbFs2IYPHJwrqocFhyA
noKlFda8tfY6nQr9S8oxgwgnr/I1HcFmmh8DMr8WgGnsb0EpUDzbI7uQ6fqXLN1H2kx8OmO9d5Si
bXFvQCOhT4Q2d5g0ohE+J9I0avqvogy0n8EEKR5AySNGXkc47irWTdxHWBuIStjFRQISYtnHqBTJ
bEBw3P28cczjX1ZaFoHdbmPiQWhrwLHrj5drdbaS4k63LtH7k9k02pz07uJtdjQE/XCsO589lCzB
HFrV+LI9Y+JKY07gePjpNaSrBfnsbdkLbAPeymhKRWVVQ+SgrDkRoGcb46dxpeazK2zfit9U6bTo
wFjihxYhfup3l6S94ZGL4WgxA0Yi91ug5Lqu4ixw45zSIN0I3IdQ/rqtz6a9kixEl8HNlSW5Kfxs
3HXqK2rB+qqJwqx/VT+mXFbJCXAiVQOP3AGKqOSjwSSFnZ4dt9i8BzkxnTxXzf6g08i3jrKIAOVJ
0d6cZln2vOVfX1EYmk0YktsqxSCh2rnh5Ie0DTKSKhfwenfXLtsTeARe+NvRDwjbsdoPnzNJr1Sb
w+YPYCyg+mdhz344n/6rXj+abo9Xz69UrgNK70eKK9m45SIzgzRanh57WBDZvQsJ+0SRAHdTfV6E
momiCX/pvKp76C4t4qiJn783m6jqGa2jIN2IK5/iFbznCAGcFI0m88iWXZhc1YnI9GVKOk8xfrQa
8yBpXu9infrKdYOOCMpu0x+e6Si9DMmbTL5ZpBOpotht/OcLVduB60QPWM9wNjvmHoGJzBgwYuB8
wvyHRL9mzG9BLXsidJXYnQQH47yjAYDzX4D9SsaG+ArltM5IirIs/PhDSR++HEP5/pyA16l4m4OM
0wUTdzdnY1qlaHySju7Je2lNFgbB1ewdXYI6N+Kj4+tRnmXb2/DMSs46TpA1RfaBFwCXOSZm9CWT
iTFkwhD5rJXJSUePI8tyWKmle5hKSXnBleW0n58Fktrfvqo+A9X090EjfgNCqwPV6M6ZlxermAJW
dYrj+3wfo0x1U/gkFpoq7lTKMsMWc638w9AE//Wtl7/5+Zg+WtCOps4YVMrNTx8JCojQXUcdgz1v
AFM5Ie1bcByt3oqZjykYZy6wghV+vYEZuDhDtt83g6BK+HlK1IGP/oB1hO5ETuuHAfGe9wDqSIF3
CQ1IGhYU/GNsEJRISoaa6LW4APcgOx5DvzMqqlQf6bOdgWznQzRcrNS4gheUPG9/gkgwIEfI7atF
IazXnxhdliuQI6yg1e2uQORnxr9w5rqm5h36QKCEd4fNbR8ysM3JG+m0rhD4EFPTAiwrSnBLUfpW
bIWZtyFZwpYGLB3nv8cnZAYDUPi9OPGC+ev2WpaNZdKQDPovaJsCKTzWHcEK7K6tBd1Yqj6q1fC/
fBJdF6F/elSitDtLxZ9h/SxBosm3hRRZAUdJwpgIqyCLHGj5W9ssqzVkMkXgbcTPxk6rc2GqNCeJ
XatZo12y8/IHPQGV3+xVMHN1/wxhE347+GseCksiNoOJsJipDbtF6t2YMGJKA+O+WTVb4Fv1BOAe
2jVUl6IBVHPU5HpY41PO6MCvQFkL5by5P+xC8wmHhGIJmrcJl0r8IeoknXrstSGo+QzykqLSzxph
CfpgzlXrEkPWgZD1kp0PuXsEjQYFGgazocHgxhutUksUFRKXHzpDL/ZFo4JWQ9pP5vQPla1UbVn+
uwQvpZp4MFStwfsr9JnlKGGsnH3Txemsbd8IZBnzRAAX6endc+qYJ6P0vGJYDUK5XpGo9bYgiomB
CEHyEASrnob1Rj0m49onC79nKj/8LUg/EjpfmUKAKbK3YfF6nhtsRg/8NbSiDv+jzdmRiPPoCwht
S9KSfM80bXWPKXoTx50ySLjuJH1F/qOND3IjgzS3he1S26mfbN3XcymU7LRunpTtYkYQZP+21Cyz
4xJJJMYwkUPQXE+X7SVPt4s+qMh58mWYr8CluPukOSy0qkvDDUtOMgrZgxWmW2YplOmQJUXPnu4U
AxBgh+bFmHa24IplLCUsiSrqNq6Gzyg++Vd09h4+phI6Z+o8y9MesylI7PuAaW2FZxaDnGVkHBbL
N+xw2yL/jgbqru9TLYlzVSTPVXHEbyBvjqy6yNgkEY50lhb4zA981E1selZ4nB5+jsKKfz3iMC3B
crFHyg2zsexhpsEA7iIhwPnwZsokYLZFA4QI97xunj0LSPYbtKvyLSC98uDd/eyJchL0/nUI3ojC
eIQV4dqy4cu3vJQTFKvikdo/tIvgZH+h9gXDRCS2AGLXHn54u5EPJkN3yNjU/rAFoZzBtj0xbqqc
+l7ZIm+4EzBGnWCLXrQclX2Gzg1l8HlSw6VIOADO732BxO1Lzq8qDWVGW4b6ExLEkGci76ouHJoZ
synAdSrQuTuhJdtU+3j/opFNkWr6QqEzxtfWcCJAbILsR9vI+6NlEMAy2Y6xWrtptOBPchPrtdc0
oIfn9vmBDmW21evuKc0OOWy3VJ1tLqBnaLArEjFgA6kBZyWgb3Qk8OV/VyTjyxqKTMycC1QY7xZH
uKjmKsRbUHDcaSvtfl9E/rsBlXyGdQUR6NOf1u57go6hMNEoRe+2ckOPEVsGDeRKaykCXqbAysuB
9IBykFdUuTMIgs166p3sDsKA00yHxWBhZUtYVPQC3ZBM2E9zzofBAiRWRmNreBr2b9V+Tn9f8N3E
B14l9QbrcMjTbJIQVVGsmX0XOCFSmRBUNxC0VWfVl+jsuC0A9+bPhwPRVFDZBp0xgnIagGwm3/GG
YMkUVVbqm9BnwgLyQqhvDVice89DcRdubKYcrC6SNACVjTTFjwbne9V+rP28A904Buo2+zqfU1XF
qv0Kw6TdUMob9IL9GY8zN6TIp0UEcto+faZzlovdEoK0Iw4odR4owiBlP79dAIzIrRky9vcVktcb
A2/sM2Jj1n5YGEh0xfORcZ18ZNoJTzvMEsxYSqgkZaLzCdOYxXhgSosmIdPGbkspTuLduQ0uiyDN
ZKR08ixRM+JhaBFC/uq8Rz/2A7TkBzLDm1f/jL43yqYabhRy2jd8ONmS8Rm/3qKeUE6w2r3IYaBC
sexZ8694UCBQrgC+UPDC4OszvKp9czNZdvwAAFqBtIcEwjfB9lcWPtmUpwhmBwv3kSw4pQKKnHGU
i7EtwqtHAl+xrGEMGI2EnR5Pwy8Reok6ZBZtAKUqNQ7WUhhcKpUwbsW/cyZ5jXS8oTTT65UWev1F
kbjEzQxHSsMppxGhFTVZrY4QsJs/htRfgWCakp0QVN4VuGfIgN4ExU3tK8wGMzt3ydA/W1b1curR
f6SX8g62ttDvqirdENTRYgeYzPMBEeLmDV527b7ouwZu8rOhteItcdJuXae1xIK8rQeedBuX8cJe
dgJqODkyHgSt9QTor9/GRm+pBSajcOFRPkDymNGCPwZKHcXVAZhdORPXrKT2aYF4gt6Ml4NytX9d
I85Kmn2v9WLhUBfW0LJ370WBrFRzrskYWdYMOs7lMiqznIF/Q8PWYZB2OOLL8qW8xDmm9tRDwZ5M
Z8J+1vs2uyuVeuDMJtznrIXxmXeXvZ51KrE0VJOluMamy292Mb16KYjNOmTWhpX8Up+feRBt9HVH
eUHTdHUJVown4KP8MhyRWKx82q43Vqy87GkD/NMTdKdRsjvfOh8l/dgpZEeGiRO6S3vTBAxEjzQA
zxFgYw1wzaucMeMI3EArxiYnEIUdUA34JQaEigWfo6AM/AX6GqBaTbUbcl4JhiL6LUCZjp6oqGva
f/2ru32QmAAm6RlBD9G5nJjPcmmic/sGNebaKqe6o9pRmcESiI5dkjgKKZ4pf+R/5WsNttVGqTgR
ticiLfevKU9HwfkQoJljbZeVw0j+vN/h7cVXbdwxe4vZZA1YRSN2HIkZXtl+lKuZeLqUa0uiq7tP
plbpLtK9zBdQA2b9r++AmZGeHN4+RyPtD/juDCTXrTZsvt1LrwCUMTVsWmqTCVnMy08yzTR2nrtF
s6/iSgsVmA96xwXfURU3Q1eRj6JD1SSTNwla/vWVpYN/984UgDaABWhgMrFQQmC7NLyIy4GQaxh6
l2S08oqCBnYeZxWLnhCsvXnYx+2PXLgQdkh3yay9i07e/phCMZ3dNowW3GxZPLRCl0L5j20UGHH1
QNv7noo/ySKfVujjKFwDPWRSKjFEyHdr8qE25JYJJzUjrrRFI41HdnwRoubn/wUMgyVqUTNEwQdg
Nhea1aKesr+yY56jcU9ZJpEtH5aUkUOAnlLY5O1P8E1LD+dtXM/0wi/aPmUS/aW3NGN9wlf0kS5y
jEMKv0WT/L2gcETLtqcyqidRVBrTB2LIhMtPMkSYgY8PPnLU/edfjX2fh12RyYsCbMoz3rFzQHlK
GZ3ZPLI/iCp5eGElyB/IXg5GRFHu32Hm9tHZeONqV8CkjHkVW+59I6MS7thVcrsyZVL72VR3SwC+
9QEqV82YkIHhecafYl/Iq3LAKWBKWnaVzmGIjxCOB/WLwsK9uF/pkCbP+m15LZlhhQ4GMBnGCT/R
l7y8e50xWiNdcAByToC5/2ImV0RI+squuv1hP8pN3fVEhMG66V5E5V39V2DY0CMqYX9k11P6mlYJ
PLae8mEerEeEV5zh35imje81PlrSKOr4Ve4XlQt13aK9YVXxA0SIluKuqkTk0KxmuKopMTChaXOV
gjtJN4CS2MnsOW5So194sVTX0WGHi8/4K5WQEXpktxAm5swsE5Un/dIZ3LY7ERAuu2kfNhkZ5Ylh
ep+shJtJQRhknPmJF18YnrUbYjndt77SCTuMUOsZ+Sa8jLT8GM/BFkxZfjkwfWZCfgkRDYAy2e0w
Gbi+kfEI6Ijtza+cSsgz7JZevfmtlKxmCvltV4q6YAD/yT/0J01VUMpbO3ZGv4cS0RIgKMJmNh0W
n9kmTJDUW7Qm/1VZ4j8ro441ceaOOzW494ca4MEzy/Yyb5E5K0UMyUO8WS2qJM2Hu7KYVOzASrN4
9q/gBc2LsC1MmMalP3wJ2GV9b57rGP0aJodk7h/n6ebThpsovSSZd8AYaOEN9u5xyNpqYlDYINeh
vz+QJ+ikm3BzMJJbz1itlxkBpbauds9P2c+kg/xHJYY+tCDCniQGQdiFmPVp/MRtchjaUogx71H9
OkN1VfmbTjqvXvjsIc1RJY32yueop/65hwhAk3sFqjxB1R7H7XcuTLBHcSjE8iiUUPKpzTSAzoJe
eL5IwBDsqkIisEe6MIH3h127G0ZatJysBPJ4kZZxroQCTnH9jkFAK0aqaD7LmaEvP6prmtxj5YRS
eCaUoccJVt8fMPccKODqKrYu9Zaoh9Lu0eLG7S5H6uaOAduxdD8Ym4LzhEOcp+9TldYCfRUPN0i2
1zW9W2iDN4O2aOJjqJ4K10BghkLVAKsvuNTBRMltAw8V8B5Y9MjR+2ZdX+MdHqiOZ5zWqW9SClny
Qudj6PTFmoZK1CPBHzgopLC9DF6ku0asoIlx/63hHgLLjlAf1JCTVOz1xzmpVKqW7cy3zXFHVSFB
t1aisgVXIofuX20UC8XHM7/nQipkIPfftZ8dRq4jbH5FLQWvbIBiEWox2MVMWyoUrdrX2VeP7KMX
qjt7qE6FFcrsp6sMZxLHwRYNPMJr8GqeM/F1uxA1y6nn4+L9sCJR+QkHLePcOFZYSyrNfGJ/08Pq
pWWJ4oqeWgCx/OLnW/Fc2UTYBSr0EbEDwOEcGXgcMdfvRgp8Kbt1gmzOj5XnDfP8alrL8r/9Urrc
Ffu0craleLIuc+FqXDWd5HGWyEQOXS1LoQRtGfiPHJVO6JphmvwHeOqIi6aFscfPFojaYWFQ6HcO
9kiaEcJ4i8VmVtzsZGwSVKCbYMxZH1g+GDeOnEmY2XIAUhfLPr4f5ldnNhgWmjPB9nsGbeOLH36s
60MfdQY/rlKrPuznRBj8+em7dZlWPx6oDMGpaxGrpvfbPSJmf0caaAYe+DqZH1uTEe3h85APPcFE
vnaexoqqto12qP+/Ovck8tzRQtGD2wXZN9jL8X81haeSdcsgxdt9o7GIPouXXdEYTA6xoAhT8OU3
DYNEtnqN4ksODuzPj5TbCF/0HpKVItInDMe0SmYzpQYUpi2eKr/9Bb6i7D3BKWrNaODAj51E8cwh
23weLY3uBs91HRWgtqtwUeIoTB2iqiL60WZLTn0K223zQG7nAuRiy25LDzFqvfRe1SRxkEQFGlBS
3ewCgPXUXV9qdsPuQOytpgVPYgH4qkj5VY9RGxj61IU2xG3gi26jV88RBj9GLIRIAP/9Rq2fgKto
nixSdTAizomH+zsya1SPvsFj11geVrU7qYFqlFE6aJCJlfPxkJMPosSFoYQNH2n4nt5dHCJsheOi
YTYce6W7JSt4bnm0n/WyioBQKUtMJd7rfoVZrweXAyzdp8xCd5wqEKHwjmB0UnsYiQNBiXDzRLzN
XwX4XFlyemivpHazRpugvSVy7U8wUO9ZVRZTJ4ZXVV1QiPR+3YoTKbUgp9RqUAEKnZPT5+vF8Aqd
2y9oDeegixQz/hrohWKSDDi2IrHtKlNHowzQYerOP6fjRzivaXdm2o67QMUYKSP65ZGP7aEB5Vzw
4NE1wkLXbD/1TqZLAuaqx+qIcnG/YIBbX6FpvZ6gf8W4kc6ceOJPXgdFQE4kiUaI143A5zfsRI4+
COJ1UxYHzfoc70FNAnffq7VgzwT91bwhYiudX/S+7pcKDsqWXZguxlskKDlAVPi1QR+prPGCP6B6
A0mS131hU5z3rbcKWT7xN/Snb6AOhbBhUAds4xSYUrwUd4+xgGxZBjkFthp3TkW9WsxnFEMN5Twe
E8SpZ8yVe3MBGIzySduQqvaI+HPVCzAUwEcklXpxp53PBCuWi+VtpqnJdsKANOQ/DP3mRn9o19GZ
fNrfLX1xx53xcO1mHa++x0HbbXf3DVso34ONV7DPEJE7+VNpOFk1BOZWXY6SS8ewLXh++FdIPkMS
hiN0SWBwkeWiyLol+Tz3o0W2GuUVEy4dDKAf8p1YC1lkNfY2QkKdo8/ChGYy4e1YYQVQq51hg9iL
Sz59YN1TZGBxddvXIyLjsGrE4YWrnWSQv5vu8Rky1wlQa6vGGFxwvuWpjgTKdIoGiu4VLHvo4rKW
aM7LFArAJTtQRbtcsrN2OPTaVmr9oFcqWvv1nEoS47KdV7FyE/3ir9SxEScrcg2amsA53zR+/1A7
Jhga/oA7Wq3CwC21BGreJTwIEoAecjF5R2Jx05g97MJpJJ4zcKCrbjvBbxOUIGvd4sezW3zjhM2X
j6ARe1DPbf1+vWWPt3xJRsk5W4LqDsNFeErSs6aSu44enEi1V4rxTbm5lmMzoCCQUpbcWBo7BunR
wzr5djsTMNwMInlStJZOTwxJiswVmXQFQndw/afdmXlV+sRe0kiHs7n60GRhXrLEKNVufporrcxL
IMSPLSyQYlLWOrELICNWnsSCQRNP5Vgyy6+3YkwO9BlnHmyHPQt7T4gRkEUMHu83dxM0n6I+I4FQ
/JxZAknbUykMhK4VUq5NXl1nwKVLbganNjrjVVfyk01265DekfpAupaNgEGEcL+g2niooud/8u1k
///VwWN678iYO7ONA0oCtn4cfQvK8R0FjZnWW4Tie3PWbf642bmXqa5zrQOd1HzEjzgTyPW0EYyD
XWl61uOLnO/Rj6sKE6j9JJizETkvKGA58ylSBeiuusJhquwsEHXvaKinFeTsZRRH0aZN1Fwh82zD
y+O/XLuFEz/FzNdcVmss6xB91JUvlny/0zFkLrO7bjgQlxEB1ruMM7jKOKs+i2CjgSpJA52jArgh
YFLyBxGAVx1UWO6GnPVNvjQZV2mpugJrZg4DkjfmNhroAfkXGfldoks/+ufMPXCunz544lHmTLvR
ynDw8P0hQmzyxQX1yfin3oNChVOZhRK4f51Q+wxIwuFhPE9ouexpvewmCDdGQtPFofAWoj1H/ZET
m0UnFFt7U4SmmwUKyo6WwmX5DigXcLjogY2vukVdaS7pvOMZ7XHewF0Jdlt4E8H0WWxQciKfMzvD
6hCOgWUz+hWjSo5yYcXk4YKy7a5Ln2U2qJ2TBjSMOGicykutHTcbs0BvkiMgL8cgvblpJYsLL8m7
gSClvDZIT/YYvi2k7ldWq0ockK2pz38oXcqZL4DFpJEukbKYzAm3OoWUT1VcCQ+QBA1Q7vYMiksy
t/JqXID7cCUR05b/vnguM+tntrRoWw9aOJ4eHWYLTHlEK1SbFRTmmhEhI43bWjkWgZlEspR88zSO
/GWolBFCmW7GSbZ1w7s5bJlg8X6wc0Fp2u45mdkgaSaV97KjHWTqgVlLLlrwNa+eHgE+B0MQUSfC
7eozSgBmUWCWbGyzpMQnZhiSMuAy+fjtADpC72oq7zldYr8jFpn3vY/K2J8wG7cxQDlkLnQH5v/K
Dfp1pyyY/oo8bpi5kuZo/0Ln/2Zaifc6Nvh9VhcRiJujjUhMU0x7mkkKx4LuOnGhU3uMBpwokXoN
tfhRG5MkDkt9bUCWbSrqcOxifWYSaP9YY3rxapRJj1Z6Il5WNd+c9S6rzG+d9r/FCgyfj+VhkqmK
lkBiBbbNEcQw3SzVYYfjkwHFJ0f1nMzyvMHALzzsO0yGCHmPWBzgQcMbEq+tf2FvNm8tw/OkoI/a
0pGjKrb5ECHguNvMjUi2OQXtb5vDH1W1siSxJVtX1ymbbCLIlYUb3AqMdUAUznuR6kNb1dfXlgnr
N9p1YwghwlRyXfsDypA5JhT+Kiw7WVyDmNvxUwanQWkbItcljj6GDzjVvYqgjxGg44/auajXxf+m
bQYyD1nzMnq/hse8gzPlHKyf6M3uVDLkDnfpJlsGsRnrn8UKSCjMG7QdzSqu5GpPGE+t3YXsF9eB
fNkvsFV2+C7G5//tmfDIYVp36CzGZm3afJRTrXuFqbju1KuxNhLvq+0zCI9AU7nlnn39RFzL7Ekm
lM/5gfVFiQlT1ZC+IrVHZFinqVH35RUCIKwZFKpltMgVjl9Gb7l9U1re9c1lAhP7J26xSIwMvrhv
IoTNSbyjnTUyObcdatqfePDbmi9an2uAb7fEQuW1cmeGwW2XG4exTIJsGgTeuFASeunHXQbd1iw+
HPLtz6Alw35S8NRYqCIM+KOQvkTFCzKzdZ6QClX86ZQbMRrR9bCtk/y3ra5S5EWfTQhKK3hZtDcc
Oq26OVihDjalekRhC49bFdauDLfTHaB59Bxp+4bd8qarX9XXTVl1hRTqw17IfnCFxUCfUfPK/NQs
XlwZCFk+aBmmsZQXzX6ahzvD0GtStaXdSGOsjdMeRlAYhJNVagXrHRb8ZwFeytwgk3hrtO2bh36C
faJkRDlQJ2nJJnHMZO1QnWylCyjDL5arWJD3UnCnp3p8q8J7q/PatOihqy63glZqNUyDAg6hGZ4m
7to2vgPXbakSznKute/SnyzGZfQ3O2dN/NTpNDfqeBoUI6t0C65pSgQSeWyYRv5Zw77KvkhLx+Qh
DKpcFYyehTZ8dQV5q1OzsHG//b0i6UiUevDun4SO0dA5AVEn+qc3UCISXUPrv08aR0sMZS3x1xZv
tFUlLutG6nuFugE389XQMwzRCfpLI+yEAQneXgRp4SrkBTStthmionjDz01jFbTfi2+VMuICpP/7
B00BZIDR7BWKevCh8pffykiikWfmGcsuzlthL/K/C5Tj14UN+ZTH6CKKeigx06ywvCvFWCi4hFoS
2nwjWGHQ+22Hg7bS77Bw7gb2M4S+tsZR/xAjkUIWlbtPS03/5mBa25Y1ASzLXN8a52yS8tEi5QC/
JhE5ayB2+zA6gZjCQwmrrYaV9+yBnEKF/+zzV6eDG1jnACyrLq5yTeu4RUjpaDfDPs0vniNMUlBm
/owBv3cELExq87ueb3BazZnlGY6CA0tBbpKlbUkw5664Fp3l15/EOZIoVTDj2IrhEypE7yS27iql
GDChXz3WTcb4bA/iLTkhZE/iNpMIx7QJSltmdjQXie8KskFvTUZRv7KgKRwVi1u+rxnCSLM71q79
BP0YS5KEUQGgzNpakzFTkqmskEnfjFBll+Zj1OGmEPPdkDvqZ+sjIeD8lg74nJxuTDjEDSf0ObC7
N2AWtR5m6yN1uU7w4f5UYF1QZwT/vHYg8UZOJC6b5yh5/hKX7VV3pkGagrsDL/rur2NppnaW5JGx
Ml9OOrcZ1du5qWdvUumajufHUf4reao5VA0XoLv816Emmt9i11sHmTkRg0BsAd56gCOprWogkBMx
MOFpUdR112QkfNzsqOuRJE6YeZQV4Ze9fY+ItbCJwdKMrTJWEByhlHAclGeRTD9WtpBjqH01jH4A
k5a2GC2WY7sgEPAWYlv2vwfodkHoj/702cL7e4L5thmVVnk/SRc/jX47BKypfeWChiwLvi6dCnZ5
7rpKC75fQEQ/g+LS7P6lAL9SjvxSikbOYxwcqWwV/UXjcz4tSzVETEMiVSLO/2y9GjFEL3e02/Q0
+eDXfczYOB1vBt4GX727Q8rLFllMAKi98ocbFQaOY3pdADMVvfVtlp5B5xJnvzSiMDoDRGR9EwmI
JbESAQjiUDQ7Lcdig4jphxsV5vaToQru1PwiMv2tlGuL0K0QZYO3/wkzJsjD6y95mkJIcaxOraTh
KRLYjfbfTaiYkPWINQLgZVgaWwhLliu3vhJPI7b/GU34Jl4oXlkySytNiOo3ac33Vef6yGh6HWjb
EmTHsmTn6VqWZXU+iboBr4m4FKkLKgkHBxQuu0YfL0eJlww4EHcvEwRQjv1avV46UdEPID5qC97f
ChMTROqrfaXRD/iZOM1z40qq8j84AKQHnTZbTIAqxFJAbPgqTtgAR+WxN9EMNHm4VILVBbte3kK5
2jsuR5TEz8j1QeXpBYYbiatgJnBJX45JIg11DY5ba6hQ10ut5L5fnFJ+tRSeNt4NnFHR63RwUDUw
xEgL9rw/e2hDHkpx4WvTvUGc8qpUjJj6ez2W+dOeeQq08XnML7+KKWF5Y3tNZwKuH4GgNTMz05ql
KiV+Jb2bihQO5x/gY2KZcOfOqyegQpJsmh5dBiDQ7zYTG+8clBi+lUPqyzxd+7BQ3jMhx0H14l//
VtTiKM6BbwcO1oEOYCcakCdhN89Eu7w4kHeVb3UE5zXrMgee16TVqNcctuQWoLen5pvFKa6YcXP4
VLNZyW8ODwuGn/r0u7sdtdJua6Lf/tQ2ZV3KZahvN8OxnXkJmxq4UWlqGv5wuvI5fUhM1ckzRQjN
Ft07jbOnDvFIbqhFoNaKc2xPgqaOpYecQEVw+cxdDKh9qSG7O8mMcM9koX51V6azr/4eZd1dEkLG
ZwEJTj5Rv8U+s/re8SX5O71ehgFZKH5S9vJgsOdEFkjmXMlH7yUyqSLn3u3yaVTDo0rlmTMKjoO/
i3c+G8zeGSglgUD/xQZc/OBC8ukhESCD0QrsfId1ZRHOlBNNIOp4/4wA3310heHs4ha4bCWLw6Pf
aowBmgIDQscMMXRFEE2NSLVWwW3BdY1hcIB0EhYfeMySLlNlU1YFM7yMln6n1ZjacvdLgdRvQ7Yr
27odrgEeeLvjO73PEkF4LW3KRvat2iNhM3t75sQMMHZJXRaytjBRREZPzqcRRldzfKw863SbkgqS
zpV6ptpzBxYjO9DdvaLUEU+SOPpQjkISsVTrJlff48frpZ2PdEGW1EToMi4TxQVHqA6fdjzfCbE+
XmZyY8A/LlwZqrSmiYIsFiGV2IaRREvzZxjiy1svRxo7RM7XkGoMAMjqYH3IqfYDsSEULlZjY3cl
JIsjk+NNlXlUHDjfIXKhLOzPxg1ssBbPUjtHyxQRWdQu4HilsMA41puB09DbSFfcR9qnM7W1lN+/
txJCwzERoRUYSIRXyMG7iW/D1G+4UyIYIgyuTujL+yrcmct/QYaru5TNuGM6R7NwLDhHuZadWc4a
7PBJE9y5CCXOKAmBNUKbPJNaTQpXrELbTqx+ggy64pv9+ljku0XmYyshIuwwtMYSa73WimcEFd2U
G8AeSEx4o8bUR61ZeWU36v7WSts/vygWmCTfbNzHaKer2PZI5g5+0/L2pWbqPjelqDnjWGFW7byG
9BuOphlLuYecrzQk9L2pqiJS0MJQvSMnnP5VO0fsjGi3Afq1b6Gi/ez2uZyouEC4A+rmAPBxHcKV
kCQGYsB281pHXqu/7ncfAdGyHQ3uVeTlJODPPiynFXBFWfelyzIr4jXBUq6W4rsDQTusO4meQZdE
CY8U9JlBXw/3TxRboySHfhcJfxFI1m/cJl47dqq7WidludStPMfZ8xNfNnQv3dd1rTmuvCYljVCq
j8OKUWFEGZQpTvGibSjpWP5FSYZKrtB4gDTZDRNpqYGIcj4rLbcZJYnKL9yjE8vuZsoDOT3DR1Qn
qnCr9RqiP/qPGXyuGuImRzAzAUqjsy9L1rMBE7GpkYv0NQWVp92rH+QkFZeLSjiKm7KImRPEirGn
Ehy74ko8XwE0vbRXH9UguebYZsO+WCZM4UgvW4NSlAZp8iJOv0KrfbQt38MPTJ1zT+ELFKZV2Tkj
GdAw5T6EtSFqHgyN+GRcKj1lBW6A/u+GXu5gNVmz4Z6MUzspjolETZLByEP3Pfja5IWZ/wcmTtJ8
LBKa1mgDZuEd01HIrFUTHFh3czar5e8hq49FXAb3DpdiRSZQyoht1CszW0RNfpkboZ114tLkwYS+
yG64mq6Nly9cwucKrgdY2JYOYrcxgY8DfMJbmodmwZ4W+YaL6atETlTgzu2rwnGaEXKR0a6ydqOZ
Nmp1IQTfqBOEuWggf85eUC0TEkO63GH/4uLeTF4seQqNUeLP8djDkbYFDMMwv+4mNkMHxD40OCk8
fc/gVWuNQuMhzx01ay5M4bQjUPBsUUBV/A/mgH/puZ8qqRp+QAZCi+Nrn67uz4sOiVpcIjHooJHU
kYL+vH2V6YNf5BKdwKxmj6J8TM3v2uKAy+npx4Iitw/NpsP00YKIZeKBbQ94Dt6M+6yuZkHBwGqL
W3cERnavtrUPmtb2RS81d1oPI+vALaSnscX65w5zOR4udLw9LAtmBg5ij0JfKN43tPemTa0LH/8C
Ih14fkburXGaE6pXNDlHl3Q3WIGy3eVduWbh8r4idcC3kFGlJlJa/2vl7twvtcJHB1Xt1tFUZ/LP
cZ0Tx1ucU1ixGLVp9cQxF7jBUPYsb+4TDP1hVDk4VJPwZ5Hces/pK/8tgwzaI/xsQC1oeXinb/o6
3a/kA2os4dK1L8EPd4LbINF6SY7Xrs1VdnQIPQ+VqVsPh2WZAStB+p6hPvTiMCInre4hXNVFdu/M
rZ4upVixrsQKkyFVt/3V6MuWP/ykATryX7DCuFtqUQtP6AFrJZ5sAYkNwMTE0Bf4v4j1KI4JM4Mj
RDZAPsdmljb+QZG089BcgimALuxPV2OK7UgYsp2+QLA9JX17IlWItnlz3xy27xPHcbMSfOQlR+e4
LZeFLWPfQjXMPLG2MFZ69WF5xPhlU8BOQsjrKoYmhQxJd6E8BJZTK3leRlEyEEY0aPfEBv9Npp6e
xaxTMXB7ATqOqLIb29+iJL6Jl7nWrtoxVe3hmTK+kmfjxSWWra2V8jwSg2nB3O8pfIZeDaCWXt8f
Q8bhmB1mJ8iyC0QeAH3i3ErIsJ4qJQL/wNSD6OUMsnz3UFLmBywyMjJCsWQ0QCCfAEHe2aGzDCkl
rjW3Os75io//62pwDPNHNdTcduq8qvMJjHhAMOu0KwuadZ5pYC0QR6vM50s/fl1xSZlTPq2kcEeR
Fn8a2tU2h0OvHnxQc7v70dKtMAzWeFEzjyk9TALJFbBqmsO/5s2INZN52vKx1YVlfpmr1ZxhsgyL
NcG1fMsHVNcHMqNoLSdJ48ndrH0aGF2hWhBht2B+ElNpBQK8CgqnDolPr1oOB3BBsr/JuW6vnQut
ERyE+GcSXlx20vMDu2ZUPj7wXUPPi6AA+4P9J/RMrn71S5XrF9mroChUK//Y8UF/4H0FUB1sZ7pL
y3f2nTmoiwYGb5r7Cv02SoN4ysA8V/he8/7y033TRYL2fj0hPBWEvQArv1ajp5icT9igZeK2+TgD
z7QMhjl1ObX7lHpJJNguOsphonoW0q1e6bOfFZdZDDKJi83sbG72l9S+SppG45BCfomyGK5rE2KP
kj6zU3w/l2jhb8IqJIweje9cWKkJJ52pMqC0Vgg/TZYp/k9RH0RujNCfR8TOA2Db5HvxP+7zyhXu
PSCRWPYw9lUscIRpHuion/eLp+HJ8PxCttLGOdJAPT8u+srnJ5XuUoHzJ3QhpSgeJVSOwxy46fOr
1cfR67DwQwI7wvntbX7JW726SugmqhEBYtMLZPcKcra3Mtsk95fxIITo7DQsS1Ei/vBVyFThzJW8
F0P4esplyLAOMmJ4tuLROonszE13HveUjpj8MwuCpgbJdamqN36jtJgLTkqLfektMmBNfVjcJhto
8/larmtVHTjLgetVe9i95I+oF8B/UTYQZ9AYn57hs4TO8CdGb17Kgo+Lpvzc7WU/Hq/54aM8Mb2M
HMUIRgvwKYq+VFe9bYPN0B2ZCfDXjmxqm6oidhjnYYGfn2Lkyom0H4QccZ2uaz6oSZChySZrOmj2
BHkUiPJGK0drakniFgKhr82XMuceyRsXB9KGp+r6CdKiJrb9kYJwpwji/y5gM5M2Xpl/Fvucptwl
YIkdJ4GyXq4UGMSQmO2rKipmcQdkJfjdfrKRV4MqRg0eF6wyy9nJ+f27zMOHwJcnQuTwn9osEtsN
hDw4rwcynHf885inrMQ0M4cj3lgQMSEV/e/9pkRNtI1usnpvoUjjUw5iFpZ/75P5P48gZJQ+eGn0
oKmnQx9svrgaxWPe1YcAyeNlX7TYNFq0bD1OAM0ERXCAH3mJ146AilU0GI8c0M72y0GcXmEBpxAl
hNfgX/TYGqhYbQq8X7pM1IEAbtFxBzPjFzCCLlk7yN2qOA962uMol2xJw8XqJZJUYUq0rR9Ki3SV
tbLHPuiU7OtZGe1p3hZJAgb7UXCABcg0nnM7o15Q6M+X2Eoj3IxUy582/KOPesQAPWEooStCFxf9
nIWoYfj1JJkrdYgDYeszAqH1QsaCEvNNR8JS9epnf/1D7pBEXewlbFgxPnDbhHI8lLva/FyPRumF
rL6N9Yf3/QdhaJ5WwzDzx3LNsM3vVErf08S9phMvkfKaJpVhff8PZiQR66q65nvcMoYOuO1F1CSG
nqoa4wzG5La0gBTvJLdZ261nU4fwj/dGL2RGEvqlbNbomB/x0u4ZB6oyPG3CmhFUqHc/R8EgZlup
gspmg5EXUD0kSHQKL5it3j0DLhUyKloZQ3urc55u4KYNZ21QORugZ50ixkun0KTauvWzgp0/QoM5
tJGpQXIdVPywHzqlKY9dn6vcsCoVNntc4QH0HwpijBXDkPKqoo6WCkoWJZZFQ659Oy0a2GSQYn0A
ouNN+ajNWl2qvfFOlpEC6a71Mi5ujX/vOgUMSpgPUsF0YdauryDnXn2giqNnkOvM51lApSPxO2b3
bNbVK+MjTUDP2I62jcygYEAiH2vk+/YRsgYSklWbtcXajxLKmv+tPa/ngISAJTT7P0qDqhGlyEfG
PrBITAIZfpldPdDtVzmeO5vQJ2A/uD/JSDPBkMaCmju4JCN3Zq/UXjZhsuBC9NkIEJ7feNRgEZEu
zwOVLwAwCRhPRiX/0q887sNJHhYSwvdC9LhybxmlnrHLmCiPaB4olAON5B4APZIj2lgymukJ+FFs
POUIo1+R/kQxTPfmAoEiEXQ9qapuY1Cz85p/RrdXtVJkk7SLNCfhKHPGfvMwdNqxbIU+i6qWYIXP
/UcXTacaWOyy/69XGw2cuqLdn9Oz/pNfJHeHfaJcfYfz+vBN0oCay1PrTg+P+VbmDyPJrwZbpkl1
gQdpMpfBFRUmtKtRsnuby8xuK15DzA5RE3344IWB94aqwR9P06r+rUIOttpBBiBQUvtHGyZK1g3Q
rNkjgAd3N1evwge6locN9l0rfIXMw7OrFYTnLX+RIfMRqzKifCLQhZ/PbU0JrYsKlql2MiQfw+3H
uhDfwxBLZVecEVQsf9tL+87SoGU61XDXrYQn/CHoJw03Y7UnSJfI4lS2rwWDL3bz5jVmjkgggFJB
y5WAy/soPRWJjQOpT2oyf0OJmpNi7geuVa9YtorfUTkYZveeolRCKwSOARwPBYAxsV5cSrRbGQJ4
AyeYd2pl2cJJjwrZvff72KWMFL6v3hpoYFx6YW4Nf2l08mTKP9KQ0dA3gwbMWBPW2onB+OhXL4+S
Mr4ABQnt14tMqv62IACDDfKIgP7VjgVyHlxISAeXoPL68ad8K8AyvGsseqvcNuLm+A7YmuX+vX5B
OARJHBmdoAdOu0JoqgSQws13T2+tbuYHFu1KDQeCC//0IR5zJjel4JhfLJ1u3Cre/P3zLEdc+y5D
GKR9Q5K8OoPCA75tGNss6pf6NbdYN8iNTYDMi+7VJrOiwWG5Zu6y9a3sADifP75owkibSWA3HlsF
El2pIqibquO2NAzUcKEzIhZ3nMRBdGdtO4V8DwgS4tbuwsxdIho8L88TnzFnkMoZNzYBYZ21hwHG
br15O1q98Jq+oWZWjm/Bh7A1DF+/0eA/oZ5wBlJ01iuaVpOiNekPQJehv7RvvUqiwIrpsbPAvbK6
FmUnNOg+UDYEmNoIm5Y9zAvSQBqRhQDynb7nTSAW0gZjP26HxTuQ6bqjngGa3HPGBvVrkzRypm4o
NIKJX1iEjUSNhMpy79OACW1FWZejVUTGJPSvbAI5zjfUHOWZn76tUpE4pCJQupUFcpyubPn74gaM
q+B/hrRrJ3oq331rGaIPiFtyLQwL5d8lvqY0hYb9U+ghCL/yBCewjxpxa80RJD1gp75zc2GiS6pE
/m5QhcEjUakBZ/LgOYZkPYKJT4tTvkWzm3/OI8eODTcj4XA0uc+0gjT+3yTqlemX56dVxC907D00
Q5f8sI5ABFVomovwOsOl+aDt+HLYTJT81WtsGW9cJBZZtyLHybFJkRZ2EobDbb/GP1e1e40GTUno
eUXMar94DGAMGoikVVRnjDaEKDFDAvdD2nTgWUfQyPau71ZyNRersdWMX1fWjLgRt3QWt4tIbG2a
H+2S4gui6xKtbU98RzWhQwE5P2W7Ef3/HBV61kRC+TnxkQaTHjEm6LEuxObufhjjNeMl7AprALS1
ya2DmdmaOXJsTXVUmK9KciSx++garUHepdrxw4rT4i82L2d/gFu1b0q+LmjnECxJMm59cK+sX9po
axzyF0Wy/7iQdXWpz9ykNILG56ekhrNvZNUH8FvqDu4JVvbI322zac0dlvUGXgwOSX4u1hRV5AJ3
Mjfx+oIUhk6dOS36thIH64YsbQT6xRWMPwl2GMXkGAyD8Yb0wwQKcS7D35Xe0Jd3l/ehsIxlhvij
/moS5GrajgwNP8yFBLt3IhRJ07XjsbzE0Q2YcWBWDKFRcoGPfrNVabKbIS1Xs+nKCSnduBgv3Q7o
9XfH12dPTfAwWr5A/f6TE21Rug0yTdY3BXm+irbDriGN61oGJOPGCwM4mA61mnoDL79m9Nwyv7QG
DGp5ZtXsqaSQdHmh8BGh38ZsHo030EIXX3JQWmfYW7nvSe3I02WD5c3JzyOBuDldyGzkZng1SYj3
ODrjB/oQxilsbx1d2OztywzmNqytiASOwvzhX76KwqVajK/PN0Fve2Q+6EPelBb9Zn+toHut576e
Tj7vYvbIaRPLWMLfq0cYzJHT09NilRtYa8Is9exTGlWcVySMqs7JGLGizP4vKxldzjYrUnHwerue
0bpsfMSJ63h29uuGM4wKebha0gLsDN8U/9lLeR9vx9GYBaF1xG83izk9laOOz2FL1zTqD6XfpbJk
jxf7z4V7BgzNy54IJk/6Bg4RhN4xVULSL0SksRrkSBTn/4aosiOPOeGbNUfV2Qelr8bEzTS7qJd0
JkFjkPQ0t99E36ri0mlNn1/K7/CWzhOocxynEluc/NZXItjKoDbv1nyJf/yofNfTIrDcLX4lb5qF
yEVmeHvK9GBRk0RqUPvXuMBiPrWaIQ9jXXKSURWZP1Fpn7pcE6Lk8tkqiVQ/EcPiieHkVZ+PNwA2
nnWBUQLXvpq6Lh07w6qL3kKxS83foc4IhWw79cTS+qlcPFpniPSnI7bwCveFA9txTOc5hoP+aA5u
cdzfYi82Qwy1N145swPI7VcuqWcANxikxDdSGAADR3y1VhaTkZah6liB8CsCN1UbRXhKuEkYDnqH
yxJhZyijxch8mGhI87yJv135IqEuq7+YFoQd77ZYZT95A5wWtNN2AtgMwv7AKQgiUn2P7lER/FXr
evVPdxy6MzQIaVyxEUSRL3CTr80Z3c9tiIEVBRXMPCprewviPA3bGgW2xQWrPJpuSugNZ+QqXbq9
2JoIakqvOFWJOzd0S3wy3OuI2ewSDi1Hqr1bSZisw+vVKBrP9LGsBUc+FPCHI6pNw4SCCBr6j97Q
EaMgR+20gM4He+OHB2HAvWgXo7VFuc0fPO2KYymNKPbdXRi52typvB2t9Vh2f+t7UbKxmLIZ3+2M
eke0+qsktogsAIyE3JuadORs3FT69SNRALeBH54GnQY9Qg8/EhZTlg/L0TwmOEUGrhE5PZ7RWKT4
0ULLGMmxXiYpiX72t/rjt01nHHCeIkDNwtgg7e8Sn3c3MOHM9i3qs8jhle30Cg6sVNg1VzDB64Q0
6mGgjLoKbSwyNmlpD2WzWLGF2uYwXnBodu15QTWak7hWyWlzjRDl5AK2cMnGdCccSXBCrYIpbXaT
UYlOl1ZYl64r0VJcscm4I3zkZ0h6Arz0WoBShzEb8K/71RZKad+EdtQa4Dwd7ceTTesk9FHz7yPf
+rTxxa+IpSR6nnb8r5WJYCremd/03Dp3kPFAdcILXSF3nwJT0A/EfjMcPs//zgOwEpluxvwbJbdM
egTRL8vRHmJi4NqPsDhTUQxWUwjE2ADjOS1FHHHvfanCPeVHQaQKnqsHn/at6YNjQJb/x5g5xul7
2pBxpHrcT2Pgz8F6hyen16RjSI5AIpLgrLcD6O4iSZ/Y2hgUS0jAGooSrumqROoTyZOP25FJvgHZ
tlw5ghAHsWqH9DhjH10dPi/RRK70mZTbrwWr0b2XlpQvm/VmB8njFBRxx7APX3LJLw1T7Od7Uy4C
SBGFVDoBtbrJ862CtxOD4+AIA8fQmy6OYBdnsp4iEbyLSvJN4laSvbKvhPBg93pXP6cSdmTfV1ws
AofJFuD9cBJqpGj2+o/0HJPPw34CBe7CJORn93yBhly5CWcKH8QAF1p6idxzjaP01Ije2AZk6XYP
g0mtQAHzJrB1zUfwa5NLXBEh44LJcJLqmlpMj+eyUI+E/kMfgiE6TqkfigGsVfueEI61u9gjbkcf
aOyyQhpIvt065Coh/hxrlEaiofHHxoiadu6AZK+qPI+oyXom5adbCdaepe4zf5G9OS3mvCzpLs1y
j7Xx4lbAgimOoR2ha6hLMFYlWOvjoGjhpRZ+4aITiR4Fe6RXASj+BTmsMLvBqXY44Eq+IhL45FP8
1pzB78GFHoqBZ2wvxjqvIurtArR1qY+wdGBGNg9oGh3ynYQLH12ZSPk/dg0XttduhYYr5JkwY2ac
i51S6ceq98CItfNLQkd3Z82GaJaY0FbW7c1+PZ1Yq5evZX7sFFxhlrfqt2xgdlGY3QodB9stcrXF
tFEw/5TkLWhgjVhrjxLIh2DrX0xeVgZrG4LiITK1ysWRbpfdk6qSZFNoJ8mR1QjRLeuMEMbO81WD
YcCCSWdixUmg1mtsKR+15UXZEB7yV8o0Hnl1b4f1OX1hyVxp7wvrOwtKdPw9cfhn//e/cHO+YHp1
KD3m43CMmfJNxZjd5jJGxpddN7RSo93Gz9pskQlGaYkPRrHlWCWp+4efhMRX7OBjh29sEf/2r6Kc
TrIMhdrBApOFMA+BlBJBJK8RuoDgnJw58RqHCWNVrmxoAkGpohW3XhAjTMsK9o4hG4RHDuzlQ+wN
zjuBuGuZO464oWuo6dWfSVgoKhieB44TEOSEtkZrwcpDpNzGeLNGjAP30vs0PfDsmLk6ClTGS6jq
2uA6oWce9aAx9bdjbjjVBWfb5jW+NqSw2GqU9P39tvT/z5HMkVy56yqoMd4Pg43jNI9tXdNH4wqb
D93rJ+N6GHjUbvUsx8+6JHqTvGRNWVoNyX6HxClZ/RybGx7Ah+mDi0D49eyXAmm7w2w075glAgqz
7SHx3T23H51djlC2sg7K1LCis5EHPHPGNewtsSiQ3foKjR2B4NRwRzmJTk7y8kdRW7VtGbNTsZD4
p46MOugXHPlNJAeMH9FP11nqrAFsqB6sIw12ypswbdulEFiDuKX4zC9JG5TaQUt4GSKyWhb8DBBX
ruW2lVgGr5VQh/zf5pEofwZTDA6p/4YAyjbLuLoH1d7R0uRm6gWANqG/EPyWhEvjKnt7zCcmWtqW
L1YWzgg6IYKKCjuZHei/sIepT5r/RDPgMGf0bdyFtxUvGN3RejjmljXEWAiyRpGboeZdQlyEn7rj
4EBYT4wPHOmrxU+vTykdRY0+BnRzWvK74Ug/39WdMOXUlk5HrzF7Eba3q3tDP2f81LsskA8Bk9vi
QmezdAXgwTU1uSGVkv7Yog5RAE+2UbGgGLD/VxjcUZ5rdfoFaN1YFYJ8577mG/p3kN0a9azSTF1X
EUFb7xSAskC2uzZ/VUq3+y05a57cjSGkCDZ0Tir30hhk5DnchO1NgQ0I2DZBH8xqiekoHFi09Y/6
KESO8mHr4fIhNSDKIOKNoxkaWUG6xH4NSFOkw53z+NSh8wJDlL/X+/6IfN1GmNCBdhApyM1w9Qhu
RCNbncL0oPFkIS91Sh+5Hfx63ObK0DCPiAckfWPr0xYcIgg7tHtveYFVPNq/vw0rorUejdf6R+/6
p2/nO1FlNPOiMjvXbLg98k/d8k+ARsVO4gD5Ybv7a/06wUuGwraczV4KocpoVetQQINnsiqLe8yo
yifXhTLL5fyII0s53GXAuaJCYNial8ImU0vpJYmA3mDo7zLLYcVmQSRrMxNZrShyF222hBTv5jj1
bC0Hu56110OTF58gVrkqxMBn7i7vw/5ld7yzjwHUhypCi3afNh4bzZOdH6JFh1u+lU3DJ/MAppqB
SJg0zdeSu1v1GQ3urEf5yj2QQmgPP2DmT7nW6V8eLoJ6qgQNTs/GXX+CU4RBV98yMVEAdP6+ibW4
SuUGW1RQWJdEasJQjTwjzEPku57/vTHo7ecbeYYuuoz7VZVQs5tj3oonz4aWde0sZyBnzHDJ20Zl
qHc21nAl6uxbheklPb5LVv1qaQYDzjOr/lqCAWyiMlj4ImLDFyF9lOLrI55CRSQ93IHzKo9T/JdH
HVXX7KfRBMBNcg/BZdA/fBD5CTxw5Rfj56YHriQjkNDhVg6lYNkTZI8OcH7uASpw/HtUuN6KnwRO
KtMe3AXd1G7erIrH2q2z0GOlTgkMAVYlOm6E1dPoxCbaKmjZV80+IYwMOUHjP6ANTqGSD6GIe3iz
bStkRiolaV9Xw2YI9aMIAs1vGphRfRe/PPFa/pNrYKe09icRDCqXXAiOzsUHLTWfYkaF0c5WY1y7
sTvS2MbSeaxdP52LpnkllLFUJBXLXeF1ZKrd+hvZBLVER4eaHrAsXJLxi6Xv9cIgpm8d3ZbM0EAn
FMInGooMO+wCP28CQQQstILzDrN6XG1aUaK8qXuqkC55TS7mMOqutbmFdLSCqNhJbRNdvpBExjoR
HiQia3+0NvnSkyg529Hl+0nbRLDuYVImPMgeaEIejLeG4SWSYMOLCjMHoEbQitnPdJ0/h69PtxNU
Pfj2vhakg9I7Khx/IFFHjyy6UMe8ROK7eXJtgLun15OJN1IErVnoIY5B6fO+y7TUnyN4nfjLjhRg
rBnrayrdRt20fbR/tQGpS5xNTyJIi+U6vHYckOwZRDcc0Cctarg1IwIELA1Jkxkb6qUHCHHVd3sE
ysqH1fSpfDQRHQtuYsXekwIbIkBJ0++t/PODRboe/24QcTRmOqeIc2c0eqVmaKJg+Od8DNXs7IlY
NTk5aG0r4t20lJijxccPclb2FA3Kdrd+HM61Wpxr6gbvhWfmiBDAnJwNvo9KlxzUOko7+sL76UJ3
nii9anF8AsvQH1WTmVdQBtie1kBWMYJHjBZUkX6mdc37IvphwPhfxv3VZkxdBSlpnse/zdvyKClQ
Hq4opx7j3tF15fkeRDYhHpg9NYlv/hqQ/lBvaixLIKT4ktoxeOqxI9UI0csxlDm4y+59uIbXmQed
GKwRvUw5syWTdnEYeADZIUyK4Y13JMjrp2VE+Jq8Rr/oBoo3Ymb8bAW2ut4UcbbmYEEqlafEeJ8t
vBCU4iV0lrQjLf7GduwxEXojJGwjEBPkfpW7XNC/f8A/jMqe5tgQ1UXmh4Lv49jvzd89iDXrNk32
CAU+PcLtcO6ysxyWPTzcqWI5j8ytL6Xc9bjHiM4i334FmenUJSEO8FP4mF2zaub0WbRmI/0HCkJZ
zwx5CaJTu4NQKkq9S5SLHoPMnyQC/mtfkB4qKlQq7hFyT5PrHULtc/VmO9Kh3hH2a6l003S3foAf
Ct6OtcRzVdj1Bwn+CmbByDN2b6d1T3Jg2ddHbUzrBUPSqElfVMOw0kxphlw+sn+tBmotiUGKUUvD
dUPAOuoetN249hfQOHuJutkVfICS5ldadBHv67+BqTUU0mr+q76KXtN6lde3iR6Nu+NX1X32Ky6s
vrH21eXw/hbt4ixeUR4K0OC/pdWgpf+0nv22ru0wJLAcCGoFF9FVHDrBVmFUWSxBkwLULWLVYfGY
UsiVF2MwdrffunQyCgOuRmPJeGjH7DNVnnEHcsZTMxMeONWC+SC60WHeThyR7MHDqXepDDX23/dD
KOAj8W0mQeb6fOzQR8s10yS21ETjO8izXpKQkRb4hnXDbVWvlYgzce0r3mfYBgGmCsyM6BMKKSM6
BZ7nGPDNATTLDnJiuvzQ5CI+avW2mvtvWkeqHsv70Q6z5fn6WwFC76maKJvl3t6Tqe574tiGfYXH
3gDTNPbkc0P9T7mBf4StxK0QuUViUc1U6alsabiWqs6wWGIQmyo0n7qFOTPn/N8JqCMBRmIwmB46
1Zngtk08659gd8InakMl1Y2oxnZUgs5D0Pj2gPOGl5hhCO1vgOo5xaYyJxbOoRc/DaBLuNgjR/W0
bC36Ru52DOGnmVjo/J4+njU5/QxTzBr7IzyTwuvLeko/Exp4b9zCyiTpRWc3+Z5rDsnQKpK4Ceoz
JsItjPSp+kT3/Th8OQmHjiNML2+7+sBkwzX28fO6TwEULGcdd4Sb/ncKgmhDm4oXLowg3lxkel6o
fn9ywt1Y+DhuR37Ohrxd9ZIhDbtr0LPh6pTI+AprFIHfNKsRhxdVjzKNx7tll/uuB7ypVenutEgA
xylnJJHa2RoX93SAyZ08IqfecP0wrloj3GrI2c7aMShLqCGUTjeNqpzPlsVeO66Hp2bDE+1lrDU3
btA1arKqPWoQ7CYaTBCmFQ3F+PDSwu6MdDrXZpbOof9VK/OavP8lrzssYcjjqdXcGe0neh04UnJh
oLa6s8CPxlaK7Z7/S2banbDO1i+kDJ9pcnPP+jkOOwBMfIA0LbnZ91KoK4nnonFYquxFgnTDbW3l
xmFpGYySGs+R984CSFX5qy98szUcjUISgYHZwEJIwv5mMHzHHgOFuQiPby6dnvOEQsVZV/NX8j/x
MPDJjEp0Twe5R4sKRRTTs4QiED/nOSsf9cj7GuQtLfMRWI6lIaghdGiJdV684s7cN9tAzoQdcnM1
ZmtSbQItRfS7mkhdbPB6/IH/78c9eCZuY/vVbBYS9XiSUe8BLG22WBNM42SRFFK97QnnDjL16Kr3
tVshZlQWAn2HnrEgSiltWlXE+ZLXWX1OPO2mlDuu9XP3PwqjBWPD0LKO3fsGHZyAKybmIXdv88xh
F01Th6Gf1RuQzX9O1a1HVH8SFCu2cltfjBRbZ97unR8ljKiljf6EsijfeDhuqv62IsLFGDxLbcdJ
e+GgNhULUkWPHT8lN2pf4FqYfHGfgeMQnATXtLVSH7auUl2BIW2aaeLH8MSnblQrQ8d7yIHhDvfA
ywZXY9EvVpQgiPbUi02Vng7vns1JwD1f+6YiBmEDbMU14/7pgHQqQr98LSAkdLeWgm2AUhGTxP7o
z9o8s0ssIkHZ9Z0c79iEn3aQuEn2SHK3lg1H6n7n/YVvwHXe4HyWdEcvmC9X2r4fw6mncnoatcwU
ly40/hTtTeVn63yHzV6TLa8SWF2KMeJ60kwqheDtQWEFfZcUNsoixpNWMczudjBRnELAhDcuwO90
JyCWNSxisE/zurG5yT1GVH3QUcz8c9C8EO87LaSNwzFa4cfFnPo9HmaYyQkJDyT3TBlgVLrGBD1Q
gSYkHKFVanf3MOJ7xZ7YAuQ6mCjXlTswpLrcHDkEsoPjtlaMZ0iUqCFjC1YrpYEkESP+ZSxgvS4E
vk6mN0YZUOvvOaswNvMcku6e3cm5PtxHfWSGxgCT0DGUykQuQmkKmC2oQlrBcgD/JIAoZ3MWHkKK
YYEOEuV2baCfir7PoidGMvJ526qYADU6n+/yuFz00B0lbsCy1fQU6W3zy5fqy1Ca/QMV7+WDHa63
FOK3KLlFsrgyt2U8hU0kyKMVLtCnPnr1zgQAwhmWVVVe+4Lc1lulNteYVoeN57fnXTcDAPyo0rlh
AA5otESbLr9U34Um9EfxcABCzFKLacGl6OEfxTnADkfUG7n0iIeFUO+YMoagnKINXwHhL7IBsthw
g6YxrjeUU7V+pwRh7RqDbVRH4JsLWTbB91grNfZI7HjwpfcQuRYp8+CHI/KMPk5VCyRcpYaqwQ2I
oq3cp+OG3unsaz3JErjkFdR5LhX+Vq31gIVA115N0F0r0FCTbPuffYB+/LlWbKg6jGVi2dvNlqJE
q8as4gZ3twalxckpsVwIFD2jVhp6M8KIe5//jhrt89PH5kb+x/+qhJMyYBKeOFlfeMxs+4xuwRlg
64cxrr+cGLd4Nd/vmOzGHKTgNGQ2SgFcttAt80xcri9xF/xXyWJoXWsc38LrDa/6YXttrp+b7oh0
fiodX/p6Y5qoMUcPu4jBSTwgwejaWronajudp2xXXu8d2qYYv6T3ytqmJUmdBmWHF5NJwE2IZoaF
+2Owq3TooOblc35CcYmJbREMjHH14zIAj8u8dyYnIoaeOUHCn1lVY9Hva7mRbyGyoDPf9Jatw69D
iZdWY6OX1bv3oU7oJNKJOnZnnAQ6G3YoGndOMB9/ljPSQT6PYgDK/dxJEV3l5UbFu5AJGy1qnDE4
2RHBegiXyMu8c0piRyc4yfOERmEEhC6YpUlsptxPCKm7hNxtNp5vDl1ioQVjJVNkw8EY3rSwKVPN
Vj3pQhMhKWabJuVxqeDQ014nfrX/mV0qGoGW6vg0YJleN8J9Bn9d9YsLR+AfJrxPfeYrZmzLC29O
i7aNYnJV4RMOO45f97DaD2nzNdMl6AI6kwXbD+DQF5O0jhZsUeEjLgbkSllWNuvIvSA+2fcrx8xp
YYry00Mhxy/xfxX/OcsQRIHv1z8jgLC69ifi8U+SvDE4HMTzLafAW56tzINYfcb9yt6GxI7fhqU6
XVVI3yQTVQgjGTo+vWWdGOYll85eEMlY6bwC8vNid2nwXu1ChPZHpjpHIy+SnkmoW8qqbz+0NGQu
YcGcYbBtGNXOLsnqkoeJ+zhzdMlcP52ylX0LjCm/qNaYHHcrAhlUOtOWjXEMf+DBgsvA+dMl4mc3
BFFhwzEvb0sueg1yD/1fCjtPz61tweV/uLIcSHBXeOPaA37Y3/+Brxavjnlyeyjqko+8fLCqhFRX
Z2oANe4zBAT1TRdQfVT6wGndA6UdiiX5sdS0xKItTnhfWhI9/AnSuBHu/iyIcD2/FHqc8yySoHAt
ksCwYEMJ7EJrLIg+62cDeIZ3FfoLNwi9d6RdIiXJBzDnF/cQSyJiyM6EwSdNHz9MMwrMOhy24Rel
sLVc2DSh3EZs4DCNlasKaBKTLBM5udb68AHaHpcO8SKM02TRxz+qzRHU34sobk3YA3uzczecV0VX
/ahKHxojjzENJXmsq8qNWzGQlzmZ1bcADfBU+dwnpZABswOJj0HlPSnz430VI2cijrA7bqNegzuU
c1UFlvmx6Tu7BdHKH14RGMF8Vb+BkdG+AZyGm4O9cJc1ADTqpw+vilGSj5RncwlKoD6EdYrmi608
63qd/52mT0dPn/3ktlGOCFfZQZEVyCnXBuF6GCXk5zrL0LsRKZgwz+uawoy8L3/KnX6Esm8BihcY
tMLSH7D7dkSjL4esKhs8qdi0Pna6NHSg5K1XRoUWYyekWAiTF8BfVuqBvM92SZCnMEyG94hqt+aF
Y5mXlRznMpPZSiJGokgDAukF/m4eG2rXZRuEfpmc2rAMZUkZQfGGGn1+UqZ1TtVEfQGjW1hWA7xp
4IaN3OP5YmGnrb3UPSurn5xZ96DdSy2TC/4qwa4M/D6A6HKbJJzUSFSO6WkoH9sORoilbDZZ94+I
qhIzgxNxb0PC192dIDA5CTEXbAxD9ZhIaOPzbk+QttQVhLwc9bSTdX4L67UXGK2+umLMzCwnoW6D
8RFzV4sJHor42P+ug1q0z4SofI0Mu3rZ5e2ut2MJvmsvViyXVvTIu9DHP6nkNqnBakAYipCslyaV
8sEa1ib5/ThYS6vJkqy2kwpk/j1GZ+/D6bBt1HGWKXpRMvLu5/ltt+nfyzPSn9IAJQogL4/PS1a4
T1N++djBQneumZ1WePXBAWy8MZjDHDoZsKW5Q70Epv0PQ3gdEfmicAz8A9Y4Nxy4iGk+Ht31ZHmi
zq8PLHjihKG00KkLIFlhs4tPsErrx0js+npYzJqNb6jrZndaovN9taSUlaz6ep58SW8bT0o4Esgf
j/jEWdwdyVptLa4JV5myjjqE23MOxxijMF7SJu0C2g1EWWcwdOYe3cBB1g5J8s0rSW+kZoUFp+CF
HpmQHkIq3NxX3zyTf/eEvJKUj0ZLw7xei+RlYHmK9j3LYOlieNXfuxDTt+gSqGxj+B9F3LpmEwTr
b8S8ZjDZvxgn0ImHuyldUmFXjMIVOHy8h5KKwg3Sj0/OEg67NMgrgYvUdu3RoJufQNjoVVMXrWKh
bZinSbIr0ECIRgwDqMMaZm0K+X+nxiB05TfQZRynuaDItbKcXopK/ezMRqRtxAgFMIVM6Qei+sCO
4n3PO7FA1CyT/2ggzd+RS4ThjdB2KH5URO/0zyYX/yh/p7+uxwxEfPTcUTxNEFD3YBerp8YSxWtJ
XccjWH8IvLUQH5X3f8zXi/UDTwynJIi4jdSH60LXzmFigTgdtYF0SvrmHDdWfB5/WgZNWc1rozV4
n1lr0f1DmYReSD0iKA+TB+EfxejzCfPZTyNSYI1WVt2Rshp75j6SZpGBtb7O9HiRQH/vtSA9c0GY
jSGF2EZWZbdoIPW/dt2Fg4odvgBOmoZo94eoVIS/N+a1UdKF1hGT+Eh4OQa2x/o1Lnz85SviEs0U
d8uOl1xl8qpEjdPJhbuXvf4bh0i9mTEN0eTvO2pRRINyNYVcUME+f82BFplAXs36Ev6vYFQWKeSS
kPZ/8jQnPUk32NhH+C2nb3xvI5tOXKbwxouk5JPAh/ri2nLf84Jk6dVwMmGZ3TGdyYZ+V/t56Lhs
fouNdeucBcSs+gv4XeLGQZqFFItYJQMMixsJr2KvHnWbNVd+IOt099bSCmXLyvrpfx6qU7VWti2U
2u73OuO7yCJbGPqIRL7nY4HHAGS39zsFHzFy3WZGEVb2rZbAt8DgKKActYHC4mA8zL7XA5oTjKKl
MUpAG8oigerF/yU7v0DT72ZyWNHeLqKWs2+8wKVTJZ4iDs82i2Q+Ve8r7+n+yPyNxb/on7qzQfHJ
jkFJF70PJKC2KUGQyP2H2AVCyqlQ0eHEoZE/HksE4/+HzVJF/AWarZGkaBhWOl+WhOxxiPfrB5zT
2U1SANAEE9Ae6sPYg7M9VAmxqgWn8B25xIEoiGvaVQoi9htG/mVMEYEdjKnd8IAR7Rgt7a5BUGEF
avmOGVx7Krw7tLuvaAboqb/GwDUrIhW2CNV0PuyGwHSGUCy2D0jAKo7zYglJoHLbmw4uozSWEDuG
tRL4yZILn8Cn8cSUEcZAjXRlLa9Y5Gy6iXXi6LmNSnQVf02k+rvs7hYngUl3BbL14GtFbQe/2oa6
s/m5kswInBK3ods+7N+R/Bu42LAc29yCKWkNG2F1iOON0RTvWhA0YjRiO/GJFWIRtpYRk9n+/Xgl
aUiJbB/3tpMh+sbDOGXNkSCmn9FcEw4wR3alxe9lO3xQY4L800aAiWVTkIPlGieMhaDuOB0gpSzN
FZH+KntpUNP1sAp0cYHYxxsaz87CRDq8zw6twhiqbs86qkcS9+wd/M/QoFvJPM0rFn2em01lXCAT
4QCwgYuV54Rc01/OC71mdwNt+oFgE8fu6vigHQcd/o+XI+3LsNsOhp2Hn8bBDkWDwRpYsff6+gU5
JBh81OZxHOKNe3ROXXYo+1f1MpGIGRp1H8F3sa0F7kFa4+XIAP/XJQoIxJpAtDFMfgLVNYZOowr6
HUKbhZSLqNkCfWeWgLtDlXfVm3sM/szZJ4UJc2n7x+zs/9QFRwdeGrF0HjIjnFYq0bVEundFMykR
s6g1zN9DajomxGQ7DpOrrYfNgFiEQ5qGenH66JIOog4eMWjVy9CdiDG7ddFISGpI2gKckl9T4o4a
jND6LEX5Qdt484bBMm8ILbAJHZJKfh4VMQ0fo4nv0tI7z+R9U0/ECGd1t/Xh+iR/+bxfd8GIj6bj
hXB+tVvuCPEVr3kszg5vkQL3TMkLfRpPl3lfJS8KqpbI4zWhYiOxMzl88Xngek1W7KShcaVDK0MD
IwASqtcnvhBg9pPiXYHGBfdpZnMBFJScKNsIIYA8OGZjyEFhUqqXxtFJM8gMsRGj9xrRigJL0KAN
u+aVt47cnPW3P4DCqmtae8Nj+iuRPcQew+QQ7Te3jzFOVtcKJX8hn6NDyu1vlmYG58g/Op2JwJRp
oqAZoSw+TcuVDMTrJ1y4R602F36m41SwQvJL+h1+ZTcyVV9TRXRKnmj6m0ilzgKIz2qHVuK9ILeo
QjE77TrrRYmkoJ03AlEyMlgvUZ1fQHRNRhBKSNiHFNTbQbm5HoTsfEyfwzU3Nw1dQBxbhsE5k6B0
HTkvrEybrxgj6tt0+fnlhl0mM+mCknDJ+dIbTkdls/d/z8dGh9rqCpMRZeRDZxx4i3jTTCpr4ySM
+XbQuKi1iXg1F+yYW4ei6kfM4g9hOOELiX4lzm7UH444msTB5eAD+CqetVo2tHQ3PMVhDOwo4Ba7
q/CyBVxp7grHAJVe5n1AEiWiKqbD0arle8SqHSDzSuiTcQIzMCoEpJbgKLfnSCJjSX79uXs/Sn8y
fDY5WgYl+5aT0OYfHUmzr47sgBAE6+qDbYrrXagBPuDY1+4Vo6Bpb30c3fR9BOqlF8w483XejAEI
g8To0mCV5MlsWNML/GG8nGKLbohv9HkISZq+DzhKPpQMbtlJKk6JgQE6U4WLdasQjxn38ih4ONG0
7nkgZ2wd2roGHo8LJIWr22bQNvtRnuONOHSwds05rK+kjBgEsrfjXIRIxOFXSJAqkZwm7Ib3d/xa
peEs8hEpKyb6Id2inwHkAtkVAc7Xk7Q36335+Jh7KaE3Swg/dfdp7mirByZWFTRGaMudiq3lvXnq
/lOK9wTYxKsNSvC0JdzRyIc9f30dZbG/2cqnBbLj+58SU35t5IZEBGzwDOZO0Xc1hKrGpwn5T0kB
BSWpDhl561SB0v1ppSRw5fTP+Ju9BY6PP9qneY6awyePPTSS7F4Uyzvfa251drZDf3MUC2zD4xVU
nAn3ww9xq8Q3UJVHXcL9HRyRuXCXjYsmpFOgXQeg+ysczqILOa8PUQO2LMHkaey3PALdR6e/U536
DEdhNAG7Fuw80EWT1NeyHMx1x8RKRy1qroBx4600q/VQBaq8RWfpaSu2ghstKZhoKyZ/zT8fYQdl
5B4Zfj7HHrenuAwzTb5jqixpgOEVLWN4OsPVvmQ71p9X5xXEZik80Om98+WUX+B4OMr+F+N/jJjb
h2SvlRxQwdtxJE1s3fxwRlQzbqk3FE8QmxskqvBGgXFhFBb9O4W5QXr53uSOqLL4bETPHFSfNTlu
7K1Hti+wraQOIl8EXc+LHp0gzAxmG1AMXx/fL0yFhK+KIHvaKWhkTClbyz6YQnuoanDtCc0OSTzE
IGN7KaXDXb7qqZ/nst9Qjvdn7IYNhDIPICDbhx1dis1/gHoP7Q1DGAB0NNUoFHR+qOS3YZ9d6N5V
sncH+Vpq+apXwsx265Vn+ZVO9mH6cTauZdzMEi0bpmbX0UP9EIVMriZ2Z2k2/qNW7WaLoxUpLlWu
kXAnQpGM/XW2XJ1F3hOrSG9rHoI0pwYYXfVAJpTqVqtI8ixY3bFsvErIV3LhmF09E8YwGf6onA7i
X69tZJBoPUvJUBQ4qquOBXdaAuhc086MT876RBP4B6oSUMd91VBlMkJXGa4QBqWZF/jGLA5uykdd
s31tjaUO9g3L9NnVIydX8BoBkNBisU3fUqb0NCW0pDX4OgGbb3VWv4Ibv046D3PFja6zNbTn9Tuj
HzpQB8leswYvHstlSMSRAafZnHhvQHV3Me1baa+7UooBCB5hS6D699ilHiqzSuzKCQ+x4zAh/w9s
MrWkUKiQ2J0oA6SCGS7Lz83o5NCOVOBpA9Pz98GWV7WgErrh87VVR6ir0oQxT+omwmCoBcP8sLBs
n6JgidPKBv4c9rnKDwdLPZmjpe+nfFFBXuRiMiwV3Ir2JJKwo1YZSyrSmakMd3RlTkDZNFATQT3S
Z9/+ZAPFpJinMNKfuTEIvzhRGJMccYbZs9FlN8nqFBPZ5u2JsXJ0If/ilDmN5xyUoM3QxfG/EEtx
x91gfelLqTt02u1lZfkGZ94ejLcWy2SEhMaIqK5YkR1Oryk7e9KxC3VwQYZLyJmhFrn+WaIjveYU
jGUcmvHRvlidrOBAthvNJyxCJd666SAajJTSvRwLhKgi/PoTwSnzjhPH8v/uyRffRiB7t4RfdMEJ
P+4503EmSnr/Ww7hOtjmwDVTFJ7SjfkiqVTpX/IXi0AqTARylaK+WSXC+WEhRTRMGJ+BGciYJU5J
Sq/05kzYQZyLj0EQfK2jyFuQrxgKkTLjhiFq+euhXvyeCb0tWnE/bll5X9dPhWpdXhNNQV5wf6ms
1ifv2nJOafqaAVcaiBlB6oRKxv5JPOJj+XJmKy6HkAiSdVVFwa7Yk9MJ88enE77KRL4GraoYXzbV
yI3IVl6UhYralcVHnyKF2w4OG5G698U68CX1lNXlONRaNUWRNl2r0SA+krYc3iSexLaTNAKukR0y
Wd+6UVJWBfpgz1mZ35kAi/CppVhF9hFcVWDQsR/4Caofwgrm3/hSbaCG/Gi3StQvH2NOt2R4Y6Py
Fn7aLssUIH/3RR2mfptp+VSVh23sXZvPzPGBHBBySy/9TU1mVytHIIJfeTrldhFY7pStDgBUJcT3
Vr3pJkVGz5RvwBUAnul5mJIMBIOQ0aCn+3YproIrr06ULia6Xb7+JGSSCDzXrabEURW5EYEZORGF
UbXJlIvoLu5CSKj0wCLxlvmN92V1kFyWy4ZlGhX1UQqomIGlObVA0EvBmaQXhKBMxkAdF0WFczgj
UVl/xGbPFl428qqaWp0utkb1aSDmUZx/lntg7uY90BSEog8/LO4BWh6ib5Lufoao38Q03/gDQAz6
ruKzFNNkqvp9CCIduz1Capy4/fWteOHVAagCUrdpzI9xnWAGSLYVv0UUQdndb4eHS0dfmBFrNib4
foh7XBX9EU0GCouE7pRcaU/PEllmntGWj7J5U2/SecpXl2CmdFNfaP85fZaCBwpiW2rkcvfTwYEo
eX+1LVYiaql9v2k8T58UrflcEzw1ECMQgySApM+P1fwilyRc16c4mSCoQtU4HmA2kUQEDX0VPlQD
/UwL8bKMKgjVqvYKLvRb1RYBC1VpMnGMlFpIMsiBqrVDoORzhcu6pldpqjVJy78wSGf9blmaHbpb
O/d4tnqHN4/k2WVCemSjvh8ApDtNeEPkz8ITfGgi8jP+0umJPciO1OgvaNBvHEO5r3tNgS33tPEs
q+j+7nW9Jq01nk2bSpzV4in6j1Uz4ENRqixvUNBVq9AYGThuHSah0y4GFoWrXpVHSQlWwJB/xBq9
Rh94/3dWbKw760binIpNXmuiyqWG8rr/Vl3gtnxe7tSLpBxHlVYx20TMhNV/7FYesOnvCXOmeZNG
2SecJWsJ2Cuhh6A5Mdj+sNcpytrXKJDYgw2LNaYLgVWuDuPVWtT37rm44AkLmS7iRYoCSIPnz7NI
tidJaOQRRTHwu2cVNNUDrPWALIEccp4Gpe3zazCknp5lImt/KGwY6Vs4XCTVzKQWFppG6ZObr95z
vaKy+u4gSMlygzKJEpbIlR+souParjLOvE4P8VAEJBqOAL9HmA03dSsCXzptXf4ncL91WXBEFZos
l1+Rd79P+rlkLsFrH0eIGCtyNXmH/4U1Kex/cd2vdkCj2F8YY+izOgCo83+DuG5caYuxN4Tdg69n
02E6aj9fQD//ha9LOaX5Ug6zVEAZlzRE0fGL/jmc7QlVGNtv/WyiiGT4dg6qjIr6JC9iUBuBLwac
9bKH7fLCFqiLoaVTlhAhCpHQuNHRkW0yfLa/p6oxmcybdilSeYljewyMHgYNlMKVpOea/YsIkMHp
qlu8wT9GW4WB+nIV/4rwo1qyAkpCyfklFXN1tVAyj2AaAZ4a+oTUadqrB4C8B2efWpEGSL1S227u
eH1c/CJ8R9OZht9Nt24gkF0DTZBNNcRK+nEQLgAxsdwBS4aO7u5FSqKNOmFGjiYxaKiwqDlotyMD
nVeK4VRJaJp4zrUa64RtIQnYfoU01UkgC2peTO+AOuE8t1BT435LYSM3qfToIjs/pseorlvRajLw
NkvOSuGJNAv2ntXUvnAduO9hHXsHx6TfBbdGRCef8soSdPrlvjOjldKBUs2WyMIRBHRJWh0QTiDR
LZnl7wcoqYazVWSfp5qrOYDutrs1z2uFXW1LsuVj1gMSSZ8HNl5NkRx2+O5Pdmk0MiNOz2aTVFPo
qgi432fVs6m4NK/9wsvcsMUNeFEkKD+N5m4dtO2baV8ko+RGm8tLDB7t0ZfEjtI3c92pMJ2S+1+Y
bzRKAeM/fWIz9wcApyMsuKGe1Ih6UQTCJRJQEWOzGfURL2PKwgZ6tzRO3tnuDDa9qVzNTMAZYkTM
mwnZJ5zWcQq/dQ1GB3s4zLsTZFd/1FV8b7IMoUzhuCKRHRWrOMBow2UQdZ7xomc7azfNrGRhru4K
v+Tfpci/+Q+2aqmkdxeNCa5EwFgT95TjfdbaQ8LE5JGRS8YiHXaKCQLCt24fxtuY36axFFCkhr9T
vy0hbNeBYQafl8HZB2E2spNjmYGXiDXinav3Pvl6x51ZcXWK3G7uKr0ZxxU2z5CdRYYMQwZLogZN
KUnBHxidCOv/RsaV0gz1OLiihLvlEscTYO4M7HES/Dwt2k3IBNUxYW++8xkyxxRDMlg5TDXtpzLS
MQ12i/+prQKbIQJLp2SQdljUBDgnia/W06bKmSgXYHXhuUyuU8nU3ey5nRRAeXSPAq+WggKY9vd5
Wxace4hBGjSkZxT5NjV03zqLcTBNIAau1EcgNR6RxoBCz2OAudOD5ZLcy+QawcAUXJNLfL1TvYET
0Uxe6YO6CkcV32hoLfGQ9j6ou69JmIBCwtX74yVNNh5AnEnkWG1Yiyjx1/kfgfvqBY7U9d7slp7U
ibrwWYUCJ5n+KmIJwHEzJWM8ZqPXr3uw3KbiOBiGleOWMWHOGFM9zLIscxDuDT+NvqAYqteI/GGO
gZzAPuzx3PdlEWF7OAZWepAHvMQ6T1ssQG9/VounKFT65U8yGypX0Mvt18IpnEHwsDSmKnwlKcdG
RDvUmWxA7F4JzWYIFsYoW5TPMJ/mrtxCeYuNCGRUj08hmnIkdTGDzm0kPpIEsmT+mr3kgIcuKFns
S8bO4elBmQ0raG1pDGM2SRg4eTVrZagjgSXRBlxPi9QfcFWHfrxgWAFRaEj45lIg+yZpxavwqqJ6
tI5LzYj4z3ViciXSC4TnYp035cH9Pp/ifa/x1IqDY+vJHzpnRua4j8DHkjL0CeMUZ9l0iqHg+xzk
jh35abttofhMusNRuqhDLlH1QN2ymJbmtYCf+zk8YWv9lUGslsTIHwjP5bmf7kbvYy+wHGk4+XW3
NwLu6vXbEGvXF/PEo9cSRYIoqG/uDo20KR+D4AIf8doXX6LTuhQUwXFHN5Xiu0g2RQHnVe+b3KqZ
+OBvU9T7T0QnTwS4ZPh6AZ9XHch8mtK6cAAygO2BtLXYU7PAVECQiKeRvRmmW1gRY/zSMrzuLZjU
gVZnnwYbrZa9XZvSUy+GAY5q6eOyUu4YetL8z92xY3ZjcanOXX6Q9eXWJHYF+wAuIyUwGDlueqq5
eSupe3vE3BkTCmy9uykbQQhdManmW3FiJKixeV7RFvnAvIG1DjvWL/O5jJYbDk+TtFCqK6otkIEl
g51GvkCWyKZ7A0mr4Q53+M52/yCIbp0du0rhY2F0cllsAbUZyZWUYUw1Sx769j0WxefAg9WgwF/b
CR+DpOhVj0SVUA/k4Ci2siAA7wPPekcaBMNd+Wm0I9qcAf6XTm/efR9HF3Gr+j35OMM+8JmlkHKp
Pq2p9Tf1ve3a3LuX98JYgb6Xwu6zcvPqL25DgYnY8iBo2o6lLahcNiiH0Ub00i+J+n+1RSFlqnFI
LebBTDiCyiQy0VDSM9FLn0PHEl3zQ4HOHetBqNiqdWviN3zsOKXdRo2/nG3taEuoynBnhtTO5yYz
FTFRwld5sMCMF7IE1ROG02KLz/iTXDxZyAurYHcJAbbu2v/nnR4u17HwGyYYj+TnY2+uVo3nMrec
2SrQBzd/1MITNorEgCh7PwzMVxEjNa9AZ1ZTohsIPCcNS8Gh3T364MciunwdJcsmW/VBDDF5BKF3
lCS4TxTkgpbpEq959ViyeZkQIEPNSBEsmVOpymDEUnD8Y6xjVfgjoH/AxKxdkK/q47atvb+WY3UE
D27ABkBQFamGASH6d8h27HBDwHeqv/WpFDI5FKMRel8sOjjZg5pWTKLiIJ7ulzafdAiVL9fWScm4
YLB4EKFgSxZ6ylPIBy3h2Zfmg91UqJB/vJs+QO0eRgb3e5U6kRL8S83ylS69hLbAUPSSDJyJUCxL
lF2l98EGr7UnL1klBIvYXoVfw826q3736mXvKWC4JmPZw9SaaY+mequS4CdCmOwc/0ob4OWhY1Z6
EDgExd4wSwuNSR2ves6P9RhIrNCnYx42BZbhQnx2v6lNTPiOIxiH/8cCnBqf9uPFvAmkRipMDg9z
HZjyA8NA/3lqoqcDHdLcWRxZxYmTFrlkzt5Q/pN5lMuzJQoUCS52jYWWsOdyfQux7qAfh70FODPn
HUiTRaLd9UCYOi+v/2oB/GmsD8qSk/6bR6nyGMOFiNcjX3apz8Q3ZbfdjK007yvrVoU7ijIHwIYP
8DYwCinrioHEpqLLH3RL4nb4qSqbnyxHnIgpxy4ycsDMgsnuBjp5obb0isA6r1Ujm7LWZqOFEHw2
MTqXAUdOlS5xz1J48atZdAJD5Ks0WEarHBJAPZ+aZWYCDgKuB3SdydKKs3cAJnwfNENohn8ey8h/
s8C0U6W4xkM+hTYxGQezVZuNQUInGm5vytl3GVG9zrvP6H9zLgkZXGho5wplynAY6VQh5kbPdogn
9qUEnaoqOaMUcp9BC32BGJnNfCyn/lhaHynUGJIFQp3yH4wFjfjr462d3MhVLudVndTfjbAeBUWe
ql2e8PTM4WXFNJZgK4QKjdY87VKJZq+Yxxp9LslCGESC0MG6aInL8Z/LcIk7o5+raFzR9gThHjJp
vJiWXCvK1R/fg8VSD98Jo+/p1zoHzv47Ae3g6F8liOIW7OGIjJfcMi2YTiIrZdHH0TcLsaOfYrI+
cR9zioKhgM8ksNCr5EIqUfjD1O/HE2VMaphUAvI6261z17jTcjZODO9xBejme8FMnCHSeR3ZDKtu
zp8vOKQZWEW9NHPRiXjuGzpgvu6VMfhh40Nc2+K67cMzTlfAYkqc+g3PjrwWNDnvwa8/UBh9TWVp
wEYsfBCY7uotlueYLMJBYyTnbCgwO5dL4JlGBAKQZxfLJGwMiOtdSLt97SoVEhuxRTn5dCyXL+v2
mPMV1lh6n/Ugx2zXH9a+ibf9iLdukSS6JMNm82E2OKeG45f5MLqyVUDm822Sa+cHag41jUhZQgcQ
ahOXixQqtCw/BPMy4nVRzY4pAvbQHztQL5VAzz3q2G6/EvwRrEuViEz9KUgTBiGaDgU7TYys4mIa
omRTt14K7ogp3nNS6FIs7etWKwl6poR4TPTE6NgUaMqSEvuX6Zx4RmErggCUW1PP6G9M3RfZ/jV9
DeF2RTxIx47HYD9ZHifBrN6DwBiyzyHszP9sv9CSXc3IFFlf3TNQLY83yThMzJYVxVH8nh3nJfjs
8FQWpqcUo8Y0yPcSLcP3vOe0JGQB9ce6hpTn5AiZQ8We/slwzpdQCgY1pLuRYyUcyQkmL4FNTnIK
PqoJ4z7WRSW44ZTDK7OZ/JJxm/XEUsRWnZdTIUf3RE9Aaom1lc4TyXET9czWV/AFw/JjAbxJKrIX
MSq0cprjLi1eQER6ZfJXyCxeFuNMOslS89nBBHIE5UZrTHXn430zzTJfarTWk2R6ji2bNbuaHP9i
klvAypQZrCfPKXOcYzqPshdF3TLgej2PJvslvVC0eKp6FQr+EBToje+HhX3heIyZFsdywMSyXpYV
8+UQub8hBxJCUm1ymo3N/UQKCeBewg81XZglcykocPs/gHRdWlrArmKeOeZRQiJ0v/EpYI3zsxf9
RQAhE4dYV91N4EytgFj3+rQjtw6zhCQDXi17Ce3Axf+6aU5DzakMXSBUFmdac95DktND/7B7oPRf
w/nYsYXqLwGJ+xsD93ldVw2neSpOrGUkA6a1iiuQNXHSaKKLBlYNs0aohoHASgKwk7Mr6+Te6DSQ
RhibKd5trfgOtY2Ei0CBU4DPpNGRA5q/sXAZ1MfAkIg6Irx4SQH8sw0QiCNpGad3xp6OhWh0++Ol
3XnT2DZ1A0wlxUi2hrcDeuFczPaf/H7GjZ+Azo8K18+m9sLA4bD7TnQhfAcTkakRKfbssQnYtXbW
0AggEpsSHQybN68YDVP7Q8i2l7IVMKqTfzlHi0wokxknaLKpB8bOr+piKtdxoWIEVvU9m0D42C+W
gX5hjhsJsqbdjBY+pJOhcCp1ksjKrV0QGcRQ20uu7RwDgs4XTsoYmCTqNDVWx3dLoerSeo3xtyIa
uiNZxa0+FPXKjr50jImjpo+SmfnujuJddxkrC4NP3dsklDaRMhKOH2SbcbqL2Ppt3ioK87i0wr8c
Y2DqjPCgFYaXuelpQoPUpX9d8WKLn8UkLT4UD8Ha96JkaLiQCiPkXpstx5UoVSZ6OdORirc9+NKw
v+8KgrlCkn3j3n1WT/2hNLGON5prCp2baVMPBbYqb4aIlbB8o2N0OBbXZBfevZ2hsb6rwfDTvJoC
PppMlLY20mGXgXRHV64k0iIdYRAhYYxcpQjvCunBdsnGc1FNb+eNgKstkGf5P8w5avAqauvvtOKh
XCeXwplVcxVAGSQ2lRRklU1diMWkTHu/rRUYAbzePwbzXbNJSsBltsbJTTVze0gIc3PffkDjl9In
U4cXHQMmn8RvkkpF589itxwXRhquSvIGQ0o1U2l60zb5V9y1HFBPXIqzLlT/elIGSn+amgmBkwYn
iUPGgMwTNdqQr1YNVeL0hAMGcrhfTrtFqjsLk+IdIRiiLg4r23PJZ9dVTLceTYZwmpMrZCLLE5q4
lpVV91AfDSpEorbMkSzjk3GzjclG4CcDFkuVgP8AIpcgvt9fn1ZnTo5feMkFIw8nSf8tpM4fyiK5
BkLLvcVQ887C7i+zEFXHzC4fEb7fjYPbGuyXsx0l8Ibab7FRHdWgzPnSJ7aykd6hcAU6g1OaopwC
rgnD6stYKyQY+nUz156CjlUoRyWbpKEj2CMFRvZf3MDycr6AdP2sfJGEIdE8RF4Y3hVTGgYQ/jNV
jwqzK2/61CslN+EWpvTvWqj8pzxpvLYnWYPthtfDyYHMn0T5XSalCUjUCuhQ8fWMQi7BfFqZi+Pi
H5byUahO0lJsZoDAF/jGHLKmHHh1i8i3JHwpYjnlmc9SryQA/+U79CxLA0JGk/0IPVWYnmWXT6pg
Q+ym4HNDwp6WldSydHk0FI2N5Rn4nzbE+sFNV6fSBdKb1ZlsKjXSGVNfAbshZ8kAY8PYe0xz801n
a5WQ9ppDr+BODAEfjsNnDnqdMbs8Oibso1PGhvLOOpweCgo+NS3wRsurKbweS9JOst4bGw6PnphR
6lXIOE8QvINwEf3gS5O+triIQQouAE57ur6up4xe9KF9zTMcJT6iNS+0k0eNO2ZlVg4/dY+0MQ7I
ktxx8TOekTIysv1lrlebp5SCrtHhL7PZaFFCIeR592hsJaGMf1HF94D4El4po7KMG1Kep5g46Xko
YFF363+Js/uPBLJHVRMPInr7LW44PWxIw5qo88zJI0E2BHW99Uz6RNsFOP6n/HkuK7+4c/LFxCIe
MEakn/ZfaEggn2+v3Nzdo9qs3OZWkXQ2fqPqS6b7OHxatWsFGogaztmf5VohtljKDrW2HuPo8YQU
9qHDdQFsoJe9pDHqKbEXMTSIUFiw1gm/uiY4AGGpnCSEVsf6S/xWh+whI1hGgkDXLDLXZTTRjmcC
PxXWuYC3yQVazwkqYNxMEu/fsSdwYW7G4ketJg8AGv6yLK2SVaRo0wHQxdFNBs5Gm2TQkfD8693A
MCPSwE4t0rVaYH4RDvSSkRbXFXrkxGfYV6zfFQfmQ+VxOpV0Q3uC6LpB+wmUj5zD3WrY8D3QkYi8
ck3CzbTz+qFS5NUIPFopCUIqW9/83Ik/R6GJn277u1DvZZU8a7dS/fjmojVDjv+K1L3ol+RUF+sB
9V6oljFC7Zt23Jjn7KeH2G53SicRoOZ2UKLubnoABCMhTY8QsFEm7GyNmrOMI99W/zGytcqfkGBv
gbNl7uUBhFw/wZO6sTLQNxImIljec8ZXdUEUAUMWxkgKO7jwX9w7OyrR7piq3lTRIYQQY8l3n6rp
w2SRhGL5lO+8jAsNLyBbAGwF5ETOAEqPytAjQhRwpUZoMWhGTbJsCb0hDNm0FhC86g97NlFtTxyL
xXnTCps09KKbrT8WmomwuqCmA9UKX669p0SfgoQPm/2FnaFB3RKMXiSrNLqufaRotjy6H1tjK8FK
lebksj3LlZ2s77w2NQBpIrywvJ5UcIDDx3owhOE3vHTNpIUbPjf+tE+nJtX1QO0BiD6uDc9He4MP
VisEw9h3DATX1qLxFTZlp+U5OkqBDyMJMd/cg9PPWrVZreDF0vPtY1mMkcjnYC0bdYhnp72VJ+z+
C6V7r7Bkfu6+i0N4icCZOTt6CPeHtK0Fm3XxHfshAIRdi0+02wSG/U28bZ8B0ZfkuvLCb1b4uLUU
Apd0QzEv5/wXbLpB7ceM/OBCveiMyByQeJvQaG/w3A/ZEGm6x5HeyY0RwXtFN/nKNpOyIDJhiEgR
i++PXZxUX2yGinEaxOMYRUL+2OQHInhUrxFyKrAF8ZwE3UvmhAb3vig2Utvgbi7HwhCTNDNPJUAN
A/r2huHvsXf2UJ1uXywzOi3t0QSdAIi5TQbwRit2prwNakAT1Up2U/y/+cATywP23dJT2zAmfiVL
ZxXMsQe5/gz8rOnZ4tnLaaoBzUbQ+16rmEmtHYh/dx7vzUmlZgxXmZMHfrfZJ5en3kziBfXqfd8b
JsFzKcuVXxlULKyoXutBeJL92fpUSZWL5JVoX9oDZGYJ5/XrdVu96avlMJeFridYj7VhC5slmNQg
+QACL5ttWEP0gC0iWroerFjmhXU0QxYhJX9jkp70OEfRNq3ACPP/ezjfgFW/cAcVxXNnAP6tBv8F
b/Yo6eT65j7fjWY7kVtFS3UHBJBRvNi0VosDz5urvllHj6bCr5QiYwhvJnahQ0JrdaL8o64v+vlN
ZsAP7jeyMS9dLO5vVWpjkOeTqU2MqVQlMnFUWQ77ikigOVxhZbxhc2xIsrMDq1K1w/h/Z5lM6y/r
6BcgrfmwdO0PXx1Y9NuIpyXy8S1Xf+ncu/LMlOjtnm0vX13/aMJCAu/Nnw05E2TkhTdV+Uk1sqHC
fOK247A/KH97EwlxTFdoZUnodyv0Z1iIkKji8w//GxG3WKu/ixQF1h5oUjSqI6/SfqIhjxZW8Yab
VJyKzVjGh+/vbpAfoTdFdH8ZurBpcSwyfp0ImmM48xk4+mQtql7XTGmlPBQU7qxf/H1MAh5v6RXL
3EpcP7SrugLbzkSbs1U8LJfwww6K6nP1mCZi9gMXlg8BE3r8R+hlLp7SOH3TzztjrfGAVJu1XxCk
nUWpv54WELiimps6eweE5z6TU3YWNxlWg0ADXD9lGd7rWBFnEdilzOPNNlRvGtsMnU6FyuNvThAP
cGUrNRa9WHlRZCemlgMlq3KxaqISQa/XE0a8DlgflUugW2EAtMpvjrKLBL/KBX4A1+CQIX/9MNme
D0M2bIMx6N6RUUMJhOxsIJeFkgJBIaygiobI55nqp3t3yuWRB2IbLlXm7FWYHxD0+j7MqWo69h/5
6pDgRnKCd9aTkc1Jje+R3rMZoWoBiZnfnFbycYzbTfkwxqTSONuIVRUAINKmDbvOOv6lfKHAx4kT
ZY7CvzPPtGjKX71s/2qjQM/N7VmFAUAdI1Qe0uBf24F3yQGrZYZ4jw9hb0XKVPlmA3EKHV+6oZV4
nLZSF8wk8FD7oWwjI+iTBaZmap6hnoPqyFGGseEXCzgONwgoG26VLjJm2sFNU8/eLijYgt16JmEx
9YZdwYS8mJi5g+6wvDBAiLo3NjfoXFncsYF2lKeHRFU6qgbDu5URluWC32Abz3oYqOK8wC1LBiyh
vohy3VBfbhiMdsCp7N0cqnqnNBLsIlTJEmHyTQzvoAb5U4zW74tIeZpsYzh3aPGOepv+wJItmjpx
aJNrIpfzJG6YUw4wF8XeKw7ucz5tBMY/p9P6wt2qpKGtwlypHY2nzMbRBZoZmGJ9QYUUYTsbchwj
5xf64dyybVsueyszNPaHHpXJtdkaZyCu+u/rE2WHp4X8iTj6mwCq1nY9iGtoVmqqgGzMm180qi7G
Iha+AED9ynenNrBHl9bKAYfxeVE7zLZCnHKZaqaDt3tilfK94Lbpi2xo2hi/1gWbmO9LAFlP8vmw
0j2hKEiLlxgLRQVwHxMROslfv09Gt4uE4RdWmwYOfcHE2/X+zlke/xjLR2Z5q2xtgfjVoCS+zArk
+iVvbqZozA8vkdKUeyV5FP5JsKCxAT7sK1nzQmSnCL3XNQmB81Q20tEb8cztIS+EU3ekk3lBtWBQ
wRcycd2GCvRGAP2XrCRdbt1TyxZh54PCZFpWgin64+RjrF1xuz7s2QaXd4s5NPVqtT4lGHxUYq8/
jHlN8FYDJZ3gvMKbxR7MSHip1yYOMF9hRBT1xbNokktQDysCAQpZYvQzrOJt3sR9mrCqbLAMHeJ/
kEAnWMnFovzhMUn9OKz+Fx1ve/cGdzuhX7ZbeyjzFZ+LBTN5oaw4iiX0Mh91R/0pe7+gSdZWvUE0
l35bN/5js5E6vKG6JyB3MJhEc8ntqWGyCj1iPzF7pjsyUm2wiHWF1+6s+g7qUPQOfjwUtXILIpVz
8AH5El/4GYD6DU7YAyi9J16Vu7T6ot2J452jzDfFfAVKvtaPoXPXik8oBtqAd07bn3wxpuUR0zqs
XMvtovtG6UcyD+SwPnmGx8cFwMNTCIdSlzSm0DqocfE2CmLvf2G3mKOpZiLD+22Oik0nWGOfn4B2
eyhYumQVV7vnawZf2lnatwM4kSJEhNmpn8B3aOS5Ji7ruWRE3gJv0SGhXK3EVu49sozEg6xM1tLJ
2F8IAoOpbZokjjffGkmxmD5Bzd+xggPjljCyyq701/Ujc9JTNEezLpSnFAN8r+VlDvEaxGFyTMOf
7kfEdEUtdNeUYPPw0axJDVoWAQO5B6tZmpyyj7abqCkhQNzAf0vL5zNHFdHEkbFJAtJZO8Kckqed
vhirTUKsxOxd1iNWgQy3lXde6K+cGmfFuPVZZkdhF3HxWLtyxEUmA4Ue00ut5pR4fDfpr90MlozC
HlfckzOvklpvVqIhA6MEFS8nAyfswTe9ATjnJvNrgaqa9lAZAwAhEudU0i5BweJLcd9xYfxNSyqy
f0lQ9oI+bxehzfJgv6kCnJGQVS5zaa46sCHnw2TZNdx+K+wKOz0vHqVUWI09Bp489I4sRtfsOutQ
/ecK75WoADyv5J5ZOwhORvsM33Q7/4mHxov6DoM2eMPoaRMbYUoUBCT4iSXRMCPKVdGDflJ7lW2Y
Yt2TUOaXcjttGl5WP0nwO/qp0UDJNM8MCIP+42djSXnq2wjzp/abCQpBMxG+Q/6ujIp+KQJLZZIZ
Ty3O3lnkxvwWqd4MBR1vDw6X8XhdPVBSvksqZLShseMTQ7ZbPm2X8eYS/Yt8Yn2BE842b3ADymwT
CKzqpJqO1ZW/ZPmuznZZgW4tFZ3MqEAj0PYFuPFChEJPtWnEyZHdmsi5Uhh9Ak1xumWJroB8ymsz
+c5oTUYnf+Rdx5dPyEsPazx8lxGDZiCs7oJ+0s8ntneprd8oluKh9IOFCDhmrPugOM2+Yk0RrONC
rrQ9hYlXdW7QFk2iORjL7oWc5Fd+6nGiGLxWyRFJM635y11ekx1AkSouf0gsGbam+vcYtKpu1mPx
Q6P5LAaSK5DzhX7pd9p5jHE2T60ImTQpwWW7yZ3Ux6O/2Dj2wPIrDxelbSQ7P/52qrNKyBD0TuHP
MMhjtClG5xoGLwgQ1CFXFU4GNGkdN4uBMI77CB6+6HatF9wRLEwsP/Q8GCgpoFdGLgUxrZysDJcx
pDcsmPPsjQ97FnrUVS69oC5fycApQtpMhtpnpOI0TjtDD1hI1iZNL8G3nJ7jZDMSfvX3FKpePUBb
/tqXQLmFXOO5/rU0/PMYCQp47kpAJEANPMwHhbGLOdRu8qmP9QY/56/YGcmvQJB7QuEWspClXPsx
H51PFxr3Q7wYj8hHfrPSTOBcdl9cbNTPr2UvExiCWL16rNaOBhBZY4TJFlULY5tcrXO9d1+if2m/
zWoJZDtSHmOten/jJMj3skFcBIcc+Mc9BtKrrOXuZSgortwqDxIVTlanHzEXJSMTdUsHK8zAQkCL
aytrEucaqP0r6z3kT1SGp5BQ7+5hBWVgpQopUpRhx8eHdOmeeumJlop/PtTEtMMtCYlHs4vqlv2p
skB6mco50WppeCxPjgh8e6n4SND9lbLZxXQz6Cu8roTJ8+IsOFo+7zCvOG9TRVW9l61ORM6o52mH
18NCxppAu9LCAeG87LuZW10baA7WvvdddCaHsSfuba5xqT1BETdMwso30khWQVGg1y/YssvsHQza
VWllNJ1i1W2yV2Uep9b46qVYCK8WIejibAKuCNq+zESUbmz7AWhCHUbNDDQhXYqMw+VSvr7hPnfi
hRpFWKw5TTLektgXBeSiVLGxMmRb9w0ozmzSZtva686MImZ6kC0CFlkd20SB7NVZjKth41a4+td9
kOnQbwb4gGMLd3HRZ5syvm4mRUyA05mBIF1Vri+QgPgiB3VQWZHDehfLV31CG3w/DlHO857xFIs/
2cIgae8eYkyAD/+4fBSqgjwofNBZZXv5o4n9cXImqH6/8lfoU950SV7Nj5OvbgTr6GO3Iy4zuU3c
oMyJAyrcUCDtH8LMGyNbCPs2pyl7MALqBNjlZfqMr5EgrO8kceER5Fp8QY3Prj5mpNq4MHO4LSpG
y1T0vFGdArJP5rzUO85XfH7nrSFiVN0MGnp6uEgVk635aUIJT1CR3VamUAcKY0j15MhtbPxYfxav
9PYA8NdaaDD0AnsCfLyMSd336lWNRhceSUjSC0YfOhGLxEq3AcJHNEeJca5/1k/NVmGpUzG/nvHK
fgz/5OeRaHvJbmPRDEsjRuCK+40MjPPqCwQZG/jTkK3xAjO4U1gYm6A9Mx2qFftxPzed9uoLD3O3
8ZjjXZ5df20eOBHFcRCV/liDkmtzEsErqMfZZaxTtSyL6okkK6RwCkEVMXTMAbcSgAPrmfj8DtuU
yFjL4FuYBPmkwL4eUSl+yVomWwsRnCewB49Shi+j+HkOzdkN+E2qxQ6Qh14Xma3cVr/7aYi5P1DU
rq+uZ++s0YIogRvLS46b/EpPNZDxXwkV8oXIC5n1DfLfiGUXqBcW2wnkNNvkf9i5o4LXi/Y73lnd
HHNiTLkdmAXGoe7eBjdSwd2+pQ4C7T2zfXS6ZPgfd1JJO3I/9gof+jeQhRZHOIwhfCGY+urYjGMM
LrpfFysHqAQvsBr0nqMqjW2rjBu61i4+rt0OwlNRL+TpAI3r+P66G5APbp3Z/RNACILrSdBb9mdZ
9SICON5GqpP38gFU45BXC27tWiL9qBQeQAc/Ank4P50yZoqxHY+jrbjEIsBMWUd6RAhQOWxGc7/w
Yd4koBSC/e/b3II4xoJZnnPHFQwlTwIUON1PyMQgycCZ4SiM5cpEYmMKCKpw6Vj0Rdiycyb7r3rD
RGWaeBwe3Cxmfcu6sQG5kr+OB8IgT296M8KBjFyyakh2CFYseY0TRwKZIq3MNaUOyB4DLT3R+OjC
vbAhuPfjjX8RJXfQJF56/orUKO434cLvrtsIZDq60ji6zbdPBYMyL1K7NW6e/dziDMRG9lGY7U5P
X8wQClAEYn0jnc+X5js0aKVz8eezTOIL0bIpoRdtslBeW15phlV3xaUsFmZzrgc8Nk1XSlWHQvPA
bdpo9XYPMmBkkDbzkq94n1afQOwIAzsHx0W0KcG4sGXYZK4mZFC7HL4kXTM749ALXg1sQma7HEx0
IVc2SvzXnU6ukdlXQobJQlDN764+n0lzWM0MDeDjYXns41FRRblW0m6fo8XMXuBBh4Vs6Q3Mw6Tu
mhTzKLP4/IhA8wM1s/wVeyH5f6/BEGz50c9YtCBDWLCyE3HlSngmSCftXBhW6Gp9kmdY9x5md/6+
3Z6HbShiao1STvNFQPCdDrb3McEY2qcyhCnn3yKkAUYqFOdQeXDToIqnjVjCaZmCjDwgvNLpy4Bq
o3LhSkYo0OxjPr6X7a+QGHkKZNR+DqjNRI/3j+CVnTMu7qRGDtjMpz/8Zf0XIQh8Hcn4T3SB9ATG
kgrlWE9+OUK3eiwU6lQwIuXv56r3W0e4ywcssYbFg2anumnUV5ctj08aPDBvkqbCtPnfPrtavrgG
H3XZ5FlSQW2zWnvJB/JV3f9LzHlI7wtWWTuX2TXqRiDoShYgaD/GtAzuDKFIiDG8oavTP/oFcGeB
2dBzfwLueGduzOuPoWuQxW7AHU5Rv51Xu9MCHqRSvjaEDNfKrj4TNcFeenZqrzRWwuHqrPyYuiMK
/bQdP2+QbZ0kI+bcGJZx1SGIHTTpuRdcihIsaEUfCczQFQVhRk3o0OX1685xqf8GnsA3zRZri+Gy
er2359b4o1Dt4WaxDm2kHg/AFNT4GeCM2IeQWIxmtW0iq3B4ZKH0It4sF0ySo741BdoEb/3Sl9O4
MEtL1Ojbx3W4+D+EonDaJqddxq9FyOvxs2IWt0BOtp9V+fhSP8veIbz7/2VhtwnFTh2R/CpzRqvq
dt81GSIVjUd0QeMyTHjy4EnQ13ckhNQ9JLJMD0CHtJZ/oxspS4/jouOEchsspoiMf2ykBd2GMGnD
IHxu1mNqNVlTe9WImjFOzgSOqYazM3J7DZc3mzilfPuWlT5/pUx4UilcJSc2K7TQlzDv7cviZLMC
DRFHBoJ4EXjVGxpBHLEw35K0a3mu1KmcsxOc4whMSh7dmeQ6+Pw4PDFq0H2PJCG9f7ODxai8tyZL
jZGsfzGPpYt33JVnWEk9H/h78flZww2NYgBkVYqucU2xeGvanWKPHRLebKpe1Mhu+u8tzhBnhV+E
sR4LwWktjz7s3a9sVTaXJ+njq+bormhzmFmnBQnDVPFETKh/QLtt+HxJTNbxDjG1+qiz8ULdWX4o
jYuNrd2BnM8jJnXcPD0hs+rEq7Zs8RWAH60lCxV6P4Fz3O7Mw8Ds0O5TOLk7uUDJTR2tFqaXVqcH
wlw6d9kHfaWXZufzYFZ/p3giX6TEOKtLTufQEp/tHItStN3A44oahTShi6eLrUUG5Qpm41WrbTED
u2dvXTmOXPE6oIbgGy6D9yQQFAWPTlE5EXIgWkUsD6co1UElUIUYDSE4Bams4VX08SKlmwQOwIu7
w44+ZfLAAhaIbEpgvv7Vbt38Nv4dunTJR5WAoIVUBHnqmMlEJ3E25wNpTFQgB3uf/GL8PDn2BzfI
/pLdM27fu73tXR78RVZywWf/vBCxWwcYM3pWYXd3JtqctnUH/69LF7a4aAYoiFp/SohASveQsSJW
XgHg5O1UfGtgwfFGCWPNYcnUrHB6rm2za6l/Kwiimkz1UvM+51RuNQOS0YOPxe9mXVFvcCZmQM1P
MJo3+jd8kWrJ8n4dTGDjNE/wzGzKh+HBCVuwMlk8fIZafKW4ON4MX1SoE0FjwongDrNPA2AeaDWw
idAhMPI18ktm95m+hS6nscKIYA9hRYjcVv1nt0KKHcdsRN/0p1wzYjWlvvDK3AGOjQURElFE5YBe
2hxgccqdyRbzoQiPuyNIcQN3qVvW+cBzheACNJS4DfDO0K7h8xWKam8Rq39YXMtF8ZJFoVTd7hYx
4UeIWB4Tlp/tJkdJAIbQ27Pm1HHqbguj4mIid8KenTYZ0TBYg2EdsHDhzD0ZVl6/KnMd+W+siHfX
lwusDSrNrv5N7p3BtZIRX2xtcZWsGye7maMUmp0hbnQ9Wo9vNptiGPbLUwac7ROt8qqI6DVdQiNJ
wjhnMss9BxJd/IE33APhohnfrtQIF/yxxfJmCDYDhWlfvZAWZ3IokTYDEfA35HIDKxoEaUnUU8gN
tiZICCiNlQbb3m0N3AUh5b/H9QsbMROPgDXJUh0gseABpwrKgHIMwrboqzyVN0wS3ikV8c9MTL37
pt4eqVTmV9nMHOPgCQdqZPwgexDc7FNMeHrFOYf2KWDt7D24M+uObkw8vrypBC78k8f5k2QFkeea
fttJgFsdQYlCCinmF+N5SBUp/aMRL0nBNxaP7d32J2AvHCDafmyHtZzV/x8quN7S9c1L2rAYG2XI
mXYcsbAIKnfwSnqjYtQ1ydAqW7kX1UaImO+WCCzyHxrP6rbA6OeoXmqvdATQh2ctifUWzmXzolw3
DZfXPYxHWCkxYNxf4hAWOf06c0wa85qnZB4LlIg5+K/K9z++5Cgm9xLuTvWHjSbGh/Blxo6lHTJ0
CevlPJfYdIDz5ZDw3Y/Luy0/uUoiRj98STOl7qsiuedRNAj/j7xXvGbm222MT83N2jkwW1Rzeugp
/He8IqWnrQdIVOzjQhyL/qRqPsecL8LrVAGUFsUjU7Etk36vUQwjpOSB89Bof8esTgc56OIp+6c8
yihFnf7pfSoZts91YYOjo4TAWpdYerWYQ42n/hLvK6XOFkMKHhTTDvyL5QT2953bmoNZD6sS7FEe
fTc+UHN2ENPHf+G9FlC694oTANdZ9Ey3+/6WU5osTKWSz/TNaVuBR8piMqI3PHUbxj7e+qecGroM
3TVrwVpVrnGoMpoDkfk0kn9meHhi4D2yBPqTR54fkCZF7LSJcAprAMHvm35XVefurWzoOmBIrmjv
QkeNe8dLA/T6joPfcObpl916oO4Wgk3S0lL31SzA8vXNaYvrw3pjaWFllhdVyxlbXT+zhD1qAJms
S4jELJ7jLhH4zdhZHFSBThqH9lME2UEcbzJc2w0OIq+s4rfkJLkwHlAacIdUF3Afq9mN/Z1KXoD7
6oKTLVBRuCU0N4J9yQczLG5ogtbW43EwvEYhg1qXGrcpszxJrTyme1q+oy5kH85PkB/JYwBNqH57
aVe4OJDeo4oScsYimV/z85HpVvdR5JcLKWa+Tt9iSrWji3ScmbV8MoNPNKJLIRwk05rq7j2G1w6l
4YUc/4beozbkUEdtS1pDsipUaq0lAwFYi8fAQikSxyX6luxyVg+presPbC2UMEqxZTndcitvOcWD
zk7eL2y+Xhz3wOOVx6UP1uXZQ+nFuabknpDDh9CjEUaXLh5PTm658JdSz5vEELHudnHBx2AH4iw5
r4IfXvoSFNToNBm0tox91tYu80mimuujirm2LMGUya2tSd5ctgTshQIk2QNjNu6s3pohC+7YV06k
rAS28H8kbqbc3YXYewIP6cAVBV0kn4Zyo0eqcmQxkohGsb27Apu4pU7qWrg6HzPBXcrVWWUBvI/V
iWdXt81csnLZm6qGOg5ALKTGqUB8gBAaN193VEaLG3KM5ptsSFc16JBU0TfTkxmA2bLdcLfKHZHL
/4O8PF0NGPOJGq8esV9XI680P8K0IFjzxVnxNsF84MCTX3L3tgJYvDmzZuGKGtXmwm+CzcewcIQ9
W54vAPBlly2+Zq6CipGtYleW/ZDCIvy5a/ttENeQIf7/iv8b+O8kh2s+/wT19M+rMERqFXl54A5b
5JmPnPZFJ4Xw2JpL/yKE0zLmso0LB+cnaybD8ZtRNYXaVdFMGbiy64GgCzokfp3aWj86JMH3CtGF
JGRU7tzmMsaA8nzUg3Mi8AlyC1uXo8a0Ok0Wm5nU427larBc1PE5yPGTvB9KVJqCeRGqpBPUlCKi
e3/iKf3thBakixKjX+xSQfrHuilJpeeLyKhyGQL+OoeH48Hd0KKPlhbgRIAsTnGrZ/WYlvA8MF/S
Vvo9U/NSdg0SHEadgI7rZ4Kjoc6QbpWeKjPi19JQ5DSiITM+MHYo3aMiXpiG2PUs2GfLg0It1c+U
0OrVvJl7fxKVPFMCVH0YaqaVlQncuaje65V2fj10dxFIkf6F70mAGnMgt+Nz2kdzhLK0hqKAPYVL
QhKAe9f8LF7xIUx+l6Q6IYLSZHxBsu5+oOpbXUrc2tU1C+wdVYN0+dEyHu/+UZwj07j46LJVT5zL
9+KcIP7AH7zQqEgtMXvbab9qSSNl+e/rjBHrrgnmfWrGzrAUlaQJ+LI8QK/xyhamnEd4o4zwsQBF
Rr+KvayvQaDf1alAvBVEs64aDL2XD/v3jUFBDyBvk+A0N6cUbFBMvc8rOVKcVzMZ+Hgp4Eih8trg
6YPi36yjGWnnqsDUbUp12iiIOwdqg4Ok4d4Rz7KV/UE0YUCiTE+Jx5p1ESheDRj5HMr2gshCj/yz
Jnak4WgDu2h3JljiY3oGM633OZi83/OwfQqZrOSO9k8CJuPC6yIE9o0Li+3+DB1W7e2snY1rGXSU
Twk7az1/9kYo0ACzXaCBQt1bahgxsFRjBIuRmZOxDEeFxBstiiqZttRWVlFMI2xFxx5xNsvXLyM9
foQ1Kx8b2xcRlURttpKW1fBg4I7WQoK/TxhrzA0ruqzJG9MsChZqGzHvphCboKR65/1Bn4byLlEn
r6U9l6zSks1zWAeYr5Hr480sgd1ulbllDxTq6RdccYq8aykey8w/fDLy/tFXn5mguZEfuYd5v6sS
/nEUJKVhmWCN1uewCySJHrso3MUvbEoYfjOcA8B8rnWq5UCrlZM+7WoBz7Wa3U4gCKGkI0TB6WVp
dHU2MW1ao9mD0aDg7ePfBmSm+bt5h1FPcqLAlqJeGI3xz885ZYaiDzST0/hhNXYzbhABQ7KYLJ3q
IxcPbDobZd8A/jbH9OQZ7KHNYVE8/g+619UBZS/4ViKE68iXVAWxndz+t8oLK+tKo7Za1KtO5YW5
WTdYNdkPSyua7MRpdbTc7M8YJAUG6OTq3RcEPbSYustIJWOgTrBhlJQTEqpyvhYOXcJ4TUqatuZu
EcAeyehjESwE718Gv5R6RekAkrYve9btidROPb97mGDOtW3ePKsbDOxogU3EN/bbrByq73DBwejv
yXrFwr3FmCZghTpYRO4U2R6BxY3t4gjB5SUA54ZowyRvxauFWbapPdo/e/qtPniM2CzzlMgW844d
YpnbQ8KUosdLgpEEpxlhTGnply3HccBBuD2/NkOde4gVt3qrdtdbSYFkD94kb2e0yUT3XiG5/igf
EbdfN/HaTWXiOJKzoPOzGIkqLn5t2/XP1S5ywXnz7TgxnzV3JgzeeJzFR62sCdU7P4mH6z1C864q
tGapx2sscnp4/1jbX6JqS5K0thcbaTpw4D/VvvAz01Pg3LKnJkrNGyLml6pKtg84YVbr2MzYFYdY
dCCoOGiqMenIpVtHfgbyuxWxIlFNk7NxdChd3Ws5zTTcXtGdFM/hjgDaezhW6SkSGp4p7VXdAYSs
eTSoB/72//gqsSDXiziRpTg0by401ozFxwz/800+Or0ndfi1dXLLhuuXVKRvJ75UQCt1eyuYU8/P
eOfhdlWDO0BCC0/vh+q7vEp6lpBcZXZnAqGEGSAFLXyj1a0tijFw0k+MTL9n126wAwpDckmxRZ3S
sRt2IEZlDJlWwssvSbE7hHoWvvxC9j0f3Lh5f8Wr+Mqk8cjHXVVTcy2hNTQsVFppA0aDNSCMkGgP
CEO12fDpdZfRfq5BzsMEVV86m9YklshPtDzEq65luaNGDdv+1Fpkl6p2h4lupDjHcwqfcV2xeL+n
xxKCN32QDcGhGY8TPm4S59jrc7KCZ0KZ1vZkDBxRTfYVT2hYh3CiG9kt29DfDe+B5soqyl0WyLtI
uYTTYb7p2OjuG2z2T48SAEpRVAiElRJo5eYN7ckxiRLwBzbVnhQg2tRlSDm1Vy9kMXfCreX3oOTa
OFUIfXG6u2EZqXEuHO0gC83tj76qGhbyI2e4dFywkeYXvn21ZKNSswwwkobUHBpSYwOb4LFzFdvL
SNvKH3/oONCnkDgtgqiQ65gEOvkE60iDy5T1QQ6j4kL1AhERagJbfIgIfzFaq6YXDok/PJ/n8bb2
S6501OaKaDy7DG+CYHGhNIPUlNhL491ZVGSB8Mfyw/TjHYW5aghh8KDcO0+kC8POxdvLQUL444lE
4wO6zs0fzCDiPH8W8mff/yC+lRJ/rcYvqL6IifYyWD2BHwEcOIzDSvr76tAxo98u0ty5HY9821NQ
6at2JnOTUMTyX+Sze6KMylfLkhpBAdCZs9O2lhi1p76GWvtSVtZdeKOn/O5BdBgSFOzbdckIPbAw
WfnF6luXwrlUcElfzQlFbWsYjl4YxR3kfrrLop8bC+StNtn2MHWC6DcVEQFFzQA/ygs4YAni+6yI
+L38oe627UYmb9Y+4H1DIRYH8GDwfGa0+uduke6hIIs5Gv1rxLbosXBg8L8cLD3Z6wB1Tnf4XvoG
pWNG8lAh+TjO6FMwDOihx2xBvV8LhTAU3Uu9pWmsC+XDgWfbjGy70DZEqY8145gA18BL8sMe75RG
Wlj/pRz7gjl+yl7xz6+J4XBuGQ4AcZ6Dyx5nOEihO9d08g2hVN6YPR8JJ/UOExOj13vHB8iKWAMU
9pLGyvIb6L4Tr/ZPZddDhDgWs5Jq0K0aiZimgrKQBJdEsTZkXXt7I6iohEugVU08nj/h9ssoX6K1
G0r2Z2KQSamZ1AGdKxJz9xIfVF+GCw2O0oi9dSMywAlUHVjer0XsiOCeHJRoKFI+G1Tv2clvm/YK
jG49Ka72qNKDn6iLjg1UZz7KTg2uq7FvJ0gxBpa9U5/pec72UKHj+x2HH6vVk34L5Vt0npsRrVta
ltLneCQN23X9ndoHbrp/6QxJ9RHFNvZBGyk2dVuoqV6/L5C4YGszLpU2bQNndniG9WWbUWVw/eTB
Qxqkgts+JVmQ6hpafr+fbQitqkD06s+hEhaItWAgkRijEo8KhjcE2XL25tiWMj1psft5DzrY5o//
2ebzagpHkflzLpswhopPoOBXwo4QYhq3NbeQ+ZO3g0u+yPO1yrdPNgHRSljgqLSyIXR+rik3TwhW
uDyy0m0NvEN5O9vQV9v8jxdOaiJZsQXfpYco3n7+TRVfinX+1AqnQlB+7+Ef4J6qe3HOaACr4g95
oGljFk+1o1sHIP8YY/+fvJiHrNU0jk9K8hswVmBb8PofFSvQZlikc0m6DTNAP/VqFOphaNNBuvR6
mBIcsq4pBwf9jq1d+WN2XD8b3kadtyPfSQ0rbR42fnThudu6JoODU/uaDT0y4tpzZbu7YL/yAZux
8bTfE20UWoA/7eQvWPTkO/mOz9rBKc3NyQYbH7pgZwnHbS4/bB6GkPVIdKiE5SNAG/mdBKUHPSvT
rWrvQcw5s0Ssng6u866QoZc/nhN/eo+62a8BNINf8b5ooxnlzUOZLsuxD0RkZDzLVMdD9Qyrc8S5
D6Vphig+COD1+Yg1ZLwbK0Gk7v8td1CGbtmuyVn0+SAGgAAo5ns5OHXPf6WDPmPteuBWEMvBRXZq
pNJcixTCQeuzaPGA34Tw+ngJ9oeRuIpViV74qp5APj0wMerowzNvibUedrImxgsL1mZMRIO2+l3e
xuHZzwHP9cQIoVxG5evQlhtlbPap2WTSUcCbEPOLNEAEhoQlKmNEV6SHW6a2hkJMSDBZ2Cplscfm
PFHLvBaW6n3+PLk7tCnXL6ch05kwCHSu+JKJRsl64gAqQGrrT+c9WIvU+RRX6q4bfd0Z7j84ABaA
CXfH5W+TmD33OBaZku8P2c53fCLLcc057Ic/YqnEcsRWbpXUF3nMKUNunPAL8xIFoDD5YWiSfiHM
cfbygyVCywSUUVoDjTWSr37peHf0jSgkaiu3K8aKYJ/gksyF+DT1Fl1poEOAjr1I21HsV05H31Ym
G3jW1PPIqSdfoUz5VNZQgs2M93MQHvu8E7rgecsb6H+M4QiS3p37UDokzieOjAP/nGkwL9T7mXCn
/nGEntrmmstDZ7KHMTt9sYHTR3EcvGNZr37EQnB9kjvn405Su8MGunfFIX9GQE2KbdKFz2m9Dyxb
q2by5IM+tCdwx2EOqThM+4WF1P4hAYYtVdGJYR+4PCDCilKtuzCywFd2O4vq5rjCbFOaB/gKMR11
Or6BDo9pIR05Jt/BGiHqq8MVDEh5/DxXy6N5vZYl2pzZ8zGPvuxa3nDdOAgJIDNIQygzHYgKjUTF
R7JL02/A1zXvRFM+rq0bf8rZaDS7f6E84fJm6dHgwzP1Ag+7b9+zzsOEMT0GbXV/e5jWYA+RzXSJ
Bwo/65Cy+447o7ioUAyXwHIWQcrGzgWFvqyRQnOgmdlaE4YvMNf8sjYt1bxNrjALqjJz+SWHJv4i
SqvYDFofPCfbcMNBajkcpeMcNz/pUu8sK3EGFCpk3yK9wNkTx8HOTxWS4YFenKymrpSEtwE1MojJ
ygW1ZTyZw558WmMUeB2qPMhwhnGHTXTEdCe3BRgZe5FNXx2G8Y2TMCBVxOuzrON4/mCzMVQJFfHC
43w64137Rqtnuxdjuh6yQ+Go9aGsWiaLvjrzkeXlxPmRcr9SQLvzPvkTf4pVc/uMicOfW0839arW
JtAFP4wcMWxotRbNW/DOBzqDdIWsT8wJvEFsgAimqMLO4EWn9nbKMtGqjUpUool3UYSB+bcJvvVy
GLAhV6D+/BZALBy+BcbWha2GWZU0XblXXjfx6rpV1vNEwh35VXq1IzLWtum9qaroHY3Lxic3Uvgq
NqOeZtXNwSbm6JazsXkbBOCU8ZTNShcKcygYFyEEk+qV8El2Auokhii8a+Nt4obNFUlqrSkSAgVT
reDXf+UO3bLddXWTyVZnYSbUDaPcnNxQcbv72oh7RzbgTDSvW9MbYS4ogCK1i9QsYWihMGgJY/MD
6ad6Zr9rNLsSrOhbGVk/5mZUdG8CErfO6G46jqCzc5NNKpjpV4SCF52wiwZdd5tB3gdpX9Tt7Hld
MkgutIpo+qrLONleOTvTp+55CKXGaQ+nTzAfxb0ZwcDSfG7xHOCrNcuzEkfD+f6mz3ttdKYnUUrE
OCSdKuBVOmq2z5vYVjNS+TfV9ndQPZFqvhzsrIRnFEISZAkRXQQbBxcE9qCWihBT8aQ3OybxG3+M
mMTQ+H0TeYj1f3sLdkdwGABHArExMcIOYKV2/9wxxjyBYmq6lbIt5+Nyth00vJDcy8WqUUO1f3yp
FelC9Iq6pvO74ueGRDp54Ana9g2XknW6k7g92EVNXRiOurNVTx3nATg7X7Nz4mCnhgFHx7gAsJgW
If5lhS5Wjo+1z0po76R0ggvEJZgIqP95lBgjWmyuMWFqk7RZ6rGg8MYfEwOHKEtR82dif7F+JyTe
J3QXj++58YktvlWgqMoKAhOfm+YcNxpal+yvjEpYip1UpK7RNYcVBbeaQ3Ne4PtnJLhAWBbMQLpq
vUI7Djyyf/o9t67QnpKznQL9esUomCXaxSgG8gT9jpyIfE0vFEllsXZ8tdkk2RlPzOwc5P6g2N3U
O+StrDCsd43tI3jl7KA/r/AIJyU3c8xGxuJdloNOnn5XMZm9MBthIRbPqxPS6zzCL8F5Qw5X5mzQ
WsM5WWz27xapB4TvcvDaSQO+9i6TnpIvzIIoYvOWYYCEDo11E1UyRYgFtFja2BHfPxUsDTV+kjkM
YXGCKTwafIPvez5xrc6gHGrNd1Lo0ArvuqpRL1YNNLH8MHTG44QYfS+6wvydgruUgx+amxTfymvc
1t7ClxNh4tt7o8UqESEWQgpvLX+5N6F0EorQrB9iNeQrDAbAp+Lu6ga7dj96KDfeNXMPbS63qwXR
9F0fWYdXZolFU7irxjc2ajwUkLcT+7PCWF0xUkUnF0qHB9qLarINoIDkIB+JXHSzprQOCvgwFs1s
E6X0VXVxDp4EHhtItF9LWNgC2SefyND3psU77GgCuK310e3GhhJm23waCpiB0ym1XwTq6yAJxhX/
kJs7jrgcW/86+ZTZPDKQb+2TVyHuZDabZlQ/8WTUL6PKfrlww4a6HP7v4lloid/K9b7qwEenef0F
gP8gbknBJKq2r1BZ4zJ2oCAoy6HrTgKdEQfz9zDTuuNeet6u/jEX+z74N7kVu8tBKTdyV7lTP6j6
+l5RNYND/d/p5RlAQqthrtYilBgzzGHlaGViZErZrPCd0YEVw4DVUVrQVqrJmVnUC57iEXFSlg4I
TTufunYMOfsG1dDvuQyH8Nat8e65aXtRJBbD12DRTyS+sKR8hVKw9nOArfc8Fx3Sujyaz6CFpG9R
83g8HYiP6E4taKQBgg/qlN65+0ewfgAdIHSo3dYxIvkmR5EYo67M5/pysfnlsEwfvCGTx1aFigf0
CD7bmXB+ksFL7XaRfHdbD2aRb+j12luyQzkQwVFjbN8iHiT17p0XEnIeDEPMMmo3HqpCH9XkH6DL
olr/b/aEJ7Mbsl6rIDDG29U8xvOSkMvsHWpvTTGYNXmXIFOIv6k0prgLYXsSpyPWe76uAIpGtrVj
UqAfQayJXqA4cgxcMuK3gxkdGLK/JiIGVy3xkquygp6Cv+n5jKJSzm70+q0JKFxqab0b9DkpcyFL
JmEqZUHuatGkeetqMXfPLXF/yzfiq/pIqlfmt5kGPQuwrWrc+sCXnj46i4MFq2nuO0F9b1YpNhNj
5XTEn93H7HbHOcm+/CQCKQEoDdpGZ9xZNgdVxXffvpoSpse5hJb2BpU8bvvNjV76ls3NPlEhxh90
BUTZbCzul4J7Lh+AqcDWehDVdXeDUz2HYVuM6mT0xnlmhVr4jaby6uNzcCDhBGa4W7xQhpByyBfh
jKrEwWprhBmn2HS6LKK9GF13t11eFEchpwho7S1hExFnikP6i4QRtZxpCJssPtbNOqmJn47S1/Dv
RBqzy1dh8N3Mf1li09FUf/srUEMCqFhGMT0lKZqAiThUbml2GKOlffQlcSE/Ka0zZBtuDari+elM
wBG3T6tV4XEcYhNHUPa+xFxYeHmeLJW8JDCYny00+6yNYmBf0Acj5dhqFxPXCO4WNmmYyyio8PBE
woDYlk5CpdALNwjaYn9zzXkOEN98stNjAIF3xjAhlSNDMO0Vh5mDCCdkIo9lxwS95UACJUQQmQ91
WzhEObne9jRcdV//epXnmiikk30vb/EMOne2JKuDvXUxfIEAKJ2WRXLXKmxbiu3rBN1BEV8C2XEL
KipxDoR5Vj/IEZHvp07dLL1/HYuOmptv8TxnSjzoctAVH2VMhBrJnS99QL4Va3pt3Bb2aOxqmgEn
gfp03ti7Ap3ETMvK1l5y3UCBqpMPZICIJ6hbQugK1ANh9q1+R/wE7TsW5GN1wDP+0Ghqdj476Fac
DgfRFU3OXYPaPb0d63RWnoCyCiVB6TN2LHu565tfUnEAopz1A+phtrup7YnXscRskygCcQpMY+1C
5EBhVW2UyG2LGqb0kZvW5lh5G4/BTTmABXjTYsqEoqTOm2OVRVWpWpX+eRrIU2viudFm/UPyXi+q
JorOpefxhW1TZwEL0PeI66kV8RRk53wIvKoqG7r2Zc7Fboa9LYYubtIfbc2fbrP99aqYGY/fXhw5
mm0Ln8+n/BMHI/zNujlanGxyIUcG3l7xkPrwToMEm2uJYLQyZ2NMFcWtdfTX+Tl4+CaCOUiFJ7yz
+2/lUoisCx2X4GYiTJ9Jv9dqztv//9XQFki4N0NdAdKzS7FhjqJvl2G8ReJ6P67QiAy6swqGMwI4
rWgzo32HMSO7PAjC5870JjtEAJl6mjOTJ64fjwTZxu0f4sUXWDPRRbz54F2Jr08ZR04SYDVv40gw
Ldkf7LX7tdD/Tsfok7nfMOcojqjnYU9eoCKhkhLJ0ri/+rlhGHKifo8y79pQcW6+kd5/OqXmdMDE
ZUie7B7rMz3I2uc3diANPa1eogCQowLAO1isVZJDX/4yvv3zxnDRkYsr/WoTqeIL/3qveOgTazUp
4g/9YVxBzzO8T3q7GBTs6HLkQQNiw7jtgNOiK7oLldiJHdlWLoNxM7vR3r7IJyCd0CMpOLA6TjyP
KPBUP1i1jXaeb7PFyVOtvbdc0C8oH8xkwp2zSsISDnDG5Rp2+cG1LQVqZCyAcaANkoOYqHIcL6VN
B6E7kTUMo8SdKUyFGNqRoAvuIBVUjS4PZJfJsjcBq68EDLWrEtXPWXnH3aOo7HPWZMJuqtR0+RWc
mQqHjtXlhp2kCWTvMHd+OQzRGMwLIec4AgBtSvEODv9ZYYPq6pi6R1AuR8c0UtpfyxqCm+VPEFE3
EIQmnKpbS0ufPyHd1ejvpkJQiAB4GXAyGr7vPJij6DqWNwjNENTo3AwSvvyrvdlyR5LXgDiYfcu+
cHOFkBTKAIzF4q9N0qAOpwl9M2tlpTc4ZQ2rwsjtJ9fg2BGuURBUzSXwXGycOYEmV423yFjIuzCR
WQP2x66t03afsuLs3H4GY08IEMvJgSqn1B2haNRYSyzk1YL2pj3BJaMoou9BQ7Go5jWO24qmwBG1
9xnVaAWRDa6JECv59RPcHyHyggF6cLcOYoVepM4WC/1ejq9WYccQB1fWXYixOpbGbOhHmnRoJkdK
JD4EZHbBo2SY7NWwNVFEIKZyRM/xMqVUGYLlDlxGzjM5L/3gU8OWtZwNZdVA4RvCijoJNLvQ6C1s
lx6KT5z0a9//FCGzQ29W+SWIIdJ75exFoizwbBKpeXqInhIwbT9ewSH246CDgNvnvfDt9H/2hLey
wpSuNbgiUE/KdyBhWxDjLQGFuDceal2BgWCMhuRDvX33KVqZMU4L3YFIbxYVHmkeg81gro+FRiVk
4r2uh/FPj+Hs9KIykgF/1PAnHeA3lHPaO68bjknTXSGI4K5/P6aW9HOoupF/ofT02Eml/8tuMAPL
OTazHLPv24HIRqoZhzR0lodb9ONlBur+/Q9/VTMzOXV7o8425rDSLSJgqwYn5lA4TQFxcUddug7w
i5oA+H/5wi5O2VHkNedxk5jydZkbAQT2XZeT2Bg7r06pPqzRjriWS7oOXJCeHN9WyaiXsbPWkHKs
WR2pE9gdhjXtYszCOdVAH2Vf56K23AuhjoJ6GyEtwSvdlU4s19FHDHo4odsJ0kGSG7yfZMKWzyjs
vGA3ZgY7BVbq+2wV49XWxFhBh1KUtBAvuIISgJW+OuGUqnWtIMGFBlenuqPZssdtYMPUA9mhTNi3
y6pogYac6P9V8j/6bVZHN1VgC+WY0j9SzDOY64VI0r7fgbPfn2ENdEzz5vLE5KmSwDNgkIzw2W72
mZKH4LNXCsJ9LkgC9/LAp143AOQ8HVw0MYLwMhTCyfHTh7brkKXvmRh/xWKKFBHkBYmZtYZYATsY
n02ys94RuTSoZPcFcwVIWQtviutd9z8jOE/CzGG9QsFSce/vxdsjShTjVrL/M6zLO0yHebvNu58s
7sLznYu0/WD/+mgNo93+2F6uvCziNT75zcdWqwa8m9cIXzfJ6+V50O+6ZVCUjkBQu+GiTE2/iaXM
ALyowtGwsGFndcNJ03rShRf9NHoPVZ8rKoT+ibtATTC/jaR28KNXeTPH/SbzEMU7pOI8K6fnoJCG
AMJMK6aEsPMkK1fnFQF3vwEHU8YZySt3klNce14/ERMmhBRRxiJUlzj7+bba4iIL7tDWcY5mxrpN
MYdsfkcm5SiF5TenPMQBhXuvXmwPR68Ufu1tQ0uBjd2g64K1JBbS289G5e7hhsYQQgPQDPPh0/cH
YnKRez1Xq8FrzAELqNKZq7ccx2scwyHthnj+BnaUi0TUb5fz49MzkUo9WHRdotH7SOAIfvHiM2P/
7H1tGYiu1tvsf4+M7EGChet9HOfOiq4MAwAo227UYsJWZn6ZoCeT+5Q3w4jepBpiu7EXhkevFSd3
pzyxhWAVOP1lQZLSy8JJ7dKINnSulRJHx6SersPo5r73oyZ0gceiibe6RgvKyMVubnA/5WUUa6NZ
HkMaEA0sHXkUS4GrCLRYSYcSbfCcL30100UtBY1QNwFjLAPx0fbTu0wbnJjmNYzEi2Zsc6EkkqvS
y/wR6GQdZMEIhphps1OE7NeXTSGKaWKaKMtJv9eCKrzPS/1ioCQwvy6Ny6YxWtfWyHLtU0eTipE7
hdmmiBPwGCGnL77ZW6ZKun8gwkr/+vy4goX38YGQeDpMbMw5wIQgElKTkTE6zLe2rl3rRS5EkjPC
w1wRlIl3Cu/9umsuX/EMY5yQvtoKL29+66zrROGSKCHXAkxUUyA6wdsbU0ozBLSenBCE1VhEM59P
316wvxmtp2OJy02CoDtX+pcCm+JLouU4RXPECbbfbJozP7dAjgxbO5/LSDsvfaz6d+9PAJsNGZYM
jC7+CEZzfj8n+F5MpkqjpXCKAw1/6+QcGAbTZHo+GbBL05s32E79OxHtvDq8dQwzKpsgcFuRo0XJ
i47KswlaSFOddTRsnV3v9SKgPrCBSy9zt6mSeChA3Hy00VoBlOCRSIfOdsK1j87X0qUaM86QqRuh
ZNbz1sT6Zc9oKC3u2c6mMZyoFKb9XDeKz6kScUuchTtBuiGmpwo74gq9fOmDqQHv/k2CIloXHFSY
YAQhpIyp5kaQCp/xo8KeWWV/KANt5vhCjloYDc1SMFr75kRpWPX+IBI2JoaCMHPiezr9O2qpHBqs
eDHneRamP3jRi0LrjQsVSP9H9XVRO6w11pQch3RBurIUgFbZW5U3ZBMvsva9BEGJHRUkm1rNvp4o
UIGL3SfyGJd7bdpXazAHpdzk5fgVt/7l1Z99wfQoaNsfO+H+6pPHZWNFxLvMi5cAvkxCZSjROJB+
IdQpWH10NJ066dmYUwwU/VlTyf2FqqHvkgig0IqSbi9t8tNHasGqyBz8W0kIKAYWNNtaOX0mFIZd
RS6Gghjo7JoZF5/AF7CfEIhjqCoyny3x845uY1nEsLBGr0m5R3z6qDQqeYkR7mpKE7jOpwXghEOF
WtMsyqdyuZOxSqRvnH1X114VuwBUBQcAfzADyvNiMLpG2Jt9oqOV2vnEvi+dl5UrDoLgLzunfGEm
pyX/8a1VMShAQBxydqrjTbxYgzX4x02IMPQ6kh/Gm3icm4VLVx4lS9ToVhqAxDZ9HLVUDK/g4ZPZ
04dbqGReJ+Ql46bQqU4N1AWRcgeE6H9/QIHbjCW6LljHEWuZC6Jsg704acMdeWkKuI/mhN4Sf0ae
LK5FKXK36ESRyiQJKYGHSpONX3HgzTynghWIl/dLua/FPbhCJyRpO9yr/kFaN52T8EN5jfaFRBTv
VYarBcWgUhNDuN49wdMmMixOkEH2tk8EGySKPVaxE/UEkwtMSYxS+ye0ymGWpkxrxJnL5Zi6fPTy
WmB/d1mn44dHE04gUlq2b5kGxYeNHHF+JZfiYTkYfL5JcTdx8zzashGHiVwGi7ehMuXry504MOpj
vyaTbDcA9atANXm2nYZ/wXH0nX/ilLZ8ZeL/jZyaMcXCl3OLKhUgT8RxNdbwiOmEjr3ypbqYCbln
K16yaqY+p9raONu+hpwyonpImgFfIcasYtNxyRFpRX1/PUVzePr+8H6ERavP7oaP317lCJnvRXJt
D6jNb5XS17pm7tcz9QAui/HXREpusJ7OOqK7dJaGFnBOLrVTdPv/p52PdCvvy+6j8OldbIcbVdoq
FgtNKHe4QKBQ2AzWuOcCA9yQ+ZZJafiJSR1a/70B1toVIE3HWc14NObKOiR1Z+ShSxaHcvFD5PA9
UJ0RdfiXdsAf87qkEnagLPu6XIIMpcMQOFoXL8OrH3zaMr00PnjxWUa7miTNcKHAFXHSFusEvKri
P22Yz93Um1667mjWAXn1A3e96fyFL46KWGUdtxzdl5xmUBKpC7mE+TZuBt+6EwMqpPRXEv7zyswN
vwQA1M1Jy5+e9AGPgUYXBVBHp8gvsNsCHgnbKJkwBNa2eeVHSkkJDwbi0xUL44UY+zwo2I0JCd6n
PzzpdyauHlMk/2kZdmrADyibcKuepCqqhb0XVR1QH5et3KOr2kRHwDEE/8gYVu/bTfQTVZH+pfPP
Vv0Nztzz7GvlOWifuEvJ8SPQ6BAUEyal/1iZdMcT5Z4crZfdHDTTektqv5P5WGYEl4SWwx7rSaR0
TKdpFDyqt68ogH7CqPK6mwWypHXx3h6P0SFUaryHdpeLklBIO+4Y2jGPEUcamtrhIFMLw9vCKttY
Fj2S+/wzI3xvpNjNHwFyGo2eygeoUJxm5z+WZNBtocdDHE+H4RcRMMg1yfVmi0NJdu9BwvZleYcQ
Up1Bed5QJ9wNwH6xfV72xXdXHUJdSc6hLPFI7GvO0bTcoIOx2KCfcBROwaLIzdO1Ai4EM/Y+7b26
bevB+ssdmjs53ykIExorfjMv9Kk1M0pDGMxNUvPDewBef3ues0VD63HBgIHhc/Fv59LzYTUXwC7K
he9tQMNA2GFax4XEWaQ/vP2vkZr4AsMACnhbYsb8WpZ9oicF+r4TO2v4mv1iqKFC6eH+R63WKG42
hrUjIw8TczrEFHVAx+mbgj33cginVh+aDg7OOhrjxS1wcSrdoVhs5rVOEKj2D48mkTWanfHD7Swv
e1gjqvIRmizFNBXdvw1ZQVyDo3v2g7IfvWp6l//Fr4cZ+v7vQ3a8qpA7xS9VoasBllP9RIu0LxDp
qK/kGCbMmEnpnu0ru9Pn1lOSV/M22gWx6fR1V4aFLi0knMYvnsIKjS1fIhbPcYt8Gh+XU2MrFMVY
HCK3OR1dphMul2Sm6fXjx6RkQm82TEBsDnaG22SMmj9gU31trXGX0sGCNTBbFW5rYg7hpI/T0O+k
AmmwYzMW7nQot17Vk/sdVqf4PaIDgEUqG2LLfl4qAo71szy2UW5vJmYRvTxSN88Egu7h0dYNgn5x
BH9Xbdb2KPM9uSi9zUVAiv9DgZm7yjzrgrjegQL6uh2MpjGI2a0QtTSyMl5j/zUhLSmqU37KnH4d
2NHbmXxcnwCI66rGilPGnQizDvzLSmATuLRMKZLlZ4aevnUZvQl+hmI/hfQ73VmyIibI0LzxbHnK
S7nQQqHuTh7L90YPZ/e+KoMPNwTk9J+w2wdUqcg30RSa5VZgYADopZ8Pf4s4Zaa6MkyTL90fRgJR
ix/Kv3VuoU7QSHAIcC0SyMHzZp1FgJDJWBQn7Z7CHZ164HViy/Nd0l+rz2UNu0a3ZnWO8v24ZjRs
JGqABnYVLwhLkpmPt0KV2Hna6Yo8YuHlpo9J1ZnN5Y4rzAIokKAVxxUSuH21jWOBmExy+e6ATcwu
kZrmwAPYF6GY9Kd2452IAP3WgdKoJ6KVKrPWOYOudl3SiJANHhbty2DXb51y966q5fnm5TsbNcHE
cvjHXbo4l2+GwKUhwhCOkPG2QCMIS3flQz5SO3qmEFksHiy+CorgiaJ79cALmtzI7OtcijIWrtNl
EanpVfzIe+6V/z/rdDvpnbd/pbh8Kr5xboE5Jx4oFTZhcjb8wd3Bpo08a5PcoJd/nhwGZ6sUw6YH
dexEWWH/uBF5weWm1SjiCUt+9obijEhKoCQxpCmaTEXFwaU614QEk2DmEnTViMD1cN+XJyqB67Tn
rXwSTA93RalzEPeaBW8Y4asddcDPMSDtPi3kKp3ZkYdEuZhMWEiShF8qg56J2XgUPSsjtTAWEk3r
9Rj9PvZQc24KI91gt7FZ1VxWYmDExUOZW7jTjoPh7ihPnA1dCpe/pcT6LSpnZc6PGYPE0Fb7DR5i
Giv8cQhhev4bNXl+X32GeGPS3U0RPjr0I6LDLxvIHBHsgVce/zeExAnr8UXHJwqxp0tVvKI2NRN4
QzbLwObhiodrDNGkP736RIi8jgACO0K/xGeaiyt1AoWqNkKIUXobVN7vcJt2cRFQzBCva0kcUHkT
pgd4dt5QFZvfCVIgz6ZyodZUw1pj/hJIlPPtILukYJ9iIjOOG/s8sSVa0FTKPqPUJnw8BaHOgy+k
Vk1+qd+mYMPCw/o3HkJ/MxP4/rzJLEb3jJNsUbqooTm4msJDBxJEqiRaNtTia/nenFM5jY+2n0FF
ZyEm0H3zM9x0N+/1j//6K0MBOmZgdub6pyozqvbGmqPl/sXcjqubkzsH0YmRZ+Kb7jrxagGz/7dy
Qy+ly9DjyQVEUptxRy+eB1inY7I829HNQvq/Hh3NCwK7N8A2ZGj4y8uT3w1me/zYGjPzo+BrgvOq
uz5SwUcjb/Y+y8JxU+MAVP08e/YR5qZB6R1NrCWEpkrzvGUePtRVo0JE/qUzvbTirsb1Wfi4BmD/
t68PPzh3yMzmDjEM2yKw2lKWjMi09IPS1pqxCGz9ixBRAJSEsF/HlF38JwxOQ9VJN/8DdSAaWHJZ
NEz22M+ug9Uo6IC+iBX1taaI+SQbJQGWgFw9QOwPUk0qhJJNehY6oo7J6eP63D+eMP9PNnugW4hh
MIjZEIAh2WSKrRTyTKp+KUoMAFyjedMXcRjzqnd7B2J+OPSPpUrFAdQjIj0mr6G72ZJ9v4v6+FI7
kFXTedOdILb5lr6GO95HwtRLr+qAuHWd0KgkhRfXJld4Wu1dTLwUw3qYo86Zww6L+oyyO2IqZXXO
W+y6AVXx7W/7/U0RQPP7vKRSI9JcR/gQl/uBnnkDI8r2iEi0COwHEkWV4JxubVzHzAlu7Bu0ZI2a
73QNqZrbNggpellNTLxzrs54X9mK/gfDCcTpF+s6hWrKgpS3lBBtr2Dc6iOTI+fE6fZt/Zcz+vQK
+4Pecb/zDX8s6Lsz6JD/c/pvIaD0OdX++IVlGgLe7vEUn1V45+8mr3PbpVsAUh8TiB7ubra6nMQb
hFtTsd0rUZ1GM0UxgUw75zJJJXxesShtHXvEyUgDfahSOMwUPiJkowxIZ15JsobpVP1zozZ+xkP/
z95AGB/WCqyrnQe6V8joWnY7MlnFifDsm3/bEG+lfiW7Ig3eMsEV2mV/LqnWRz8NOlbDcvWBfFaR
nPkZIJhDzPz9wZnsj1+RmYBtB43YzpCdSN8i0OfbSZxIv0R8y06hlq5z/PtWRFQnYnlQHbzzuivi
molnX4a5W0xGDbEC581gCykpPoBKMkWWwlvj7gsW1u89/hlDoD83Xr2EXdOFMUVATP72pTywztQN
Ne8PdGSCkQNusEz0/ZT2Yf96ocIWcg+ZjU523oL1YL9dI3x4Puuv6U6X11CQJcPuJ8z36Q+DGV+I
KvYTrCS7ElaTNbv7yw7LgSd1uMC3SVkirdUUYoEmFWnGz911NOtbs3YOEUG34EFidA2ks0mYCf+x
om1amH1751gTJ1MPqQICaTFziK6Q+VRpvOPN9rBKr5Ix9vuKZ0ApEp3Rqx8Q3WjeD3So4pTlJEK9
cpfgpv5VvwTqwk8Z37v8OM+MOT6H31Fac9NhECjebnbpH4xxBSurP1IC2YFRKjd1U7Y/WNseOZbz
DUOS+Ky5NOIqOuJ6Pi74msuYDiwShuRP/B3yCeusS59Sge88O+QHGoiZ4UwRr7Dj3WV1Uh0cxXaK
4PDPsbvHW/I4nFGMqaF0GChnNpKAxUJIpNfDIduLzN84QmS4N4U3Zj9rCQa1av6WNYFFbu/3opoT
RO/EOQSP+KUuOClQoIiBz5lxAaFsyTIHwAZK4z826PWA6VPPGoXNh3R5Pf3PU2HyVNO8VTkY3yuH
qLdBk0AeVR8rYWXik3OWu4h8F6RySpY7fgYUp1bkHlXhs7TpwwcBSmcjXBlbXu1KIf6j38qbM7w0
JWOmDNb89449gDhlEdpHUIDlmhv7tQehY5vHIiGzO0fhsHinP+b+XSB2WqN9uGKwQS7uduzHj+1f
Qo6jExUBRvdGVDxtqyN/iK7mtEeAYKZQW071yL1uaERJWepZv5JRSB3Cx7tyWV/RDJUBvjycrlQL
AHYi3zwZki4gc5VB8sNgVoDokCpO2q6ZOfgECK2p8/T4EkQu+cC3NY/aNn7bslypLFPNBZ+SghWb
ckIS/39SCqw66kpGjlAo0qDDzRtMbkbUGjZfp//jfbk1YODaTNy89DbjIwsd6ImTP53EDonri79F
gX0Pg3LBraNhVyQSykgLNXpUjpU3Nnr8YIcAfvJpXBDZzTf28O47y0aBxo/G3Oif2KTe97VPz0KI
32pR1dMEDqtTM3T/wVJzH8RrNcSS2ORVvud1bOgCgVY7w0Q/J8rvwVfypA1g8VX88qzrXvGM/nE4
dt+pi0LalNBDb5Y5AQkMpXkewS2VNAmuAi5zqe0I5oTbELZwjSbN1kCn2zLkbNJrgmEWFtNIO667
pOd4er2iNdoWxGEahye3Qp+Cd/wurZ1hK+CEedEjs9ir7acsNvsqiUoW5Jfh5Sy2V2PzO6MHIb4P
4avVcC9J//uNQzce1nQDvzbUDzVXvRSUkHzflgnKRFYbY0HgK4cUTKzHOC+91rWxBUeIq5yQ4sz6
PLfEiKCl7eVw+k/eozlPPIaJQRWBulzc4SOECKsmRWoqZCvYFNui4YMYqpYzUNmGma2qEd7PqQRm
/7noyR2+5SyCXcNmDMth8kcEslj5FKpS2nag5gwqeT+eJS49kowI/VDl2AWmxdEnW/fI+X5bMEF/
enHd5t/9YaoNDeE87bt4HI3wUl8HtdaSbcDMyvKixg//iFUtFRHLxdSG/h/1gsMNIjrVKTOiR25H
q8CErxEUCdicsuhB3GAJOzwXAI3t4edVK7FfSYzOFZ7BVC5oN6q1BYQBuvSwpKYluQlFENr+nSG8
ftqc+3cqstIU4SVvXx+xV91XPoif2/h3gKnWSsynMuMj5xUtRKcV7Mmtj60FgF5kHuHUqsSq5Nlx
687B4QMW/X7J9kGxLWBBT0mLQnEBxK3IjHN64oJbfPsCTA+JTLLm23kki1PozlWGRqMRFAHk9D/g
4zSRFwW0p1VbziGW0TbWx6f9hb2BkBdb9UUE6hmPI8bnol5vNff99k5VxXMLLIEL3YCY1oCpfhTv
RItms8OVmqihA6CfnZ9PRpYmQhnTeq5Z/Q05GpZIyD4hl3n15VnAU09eXNDmkdcIfWJg9mITwuxV
hiGjF0GPe0yLWDdCe0IdZM+dhiDu7BJccvQ83hIrBo0jOdzjzEfaflZBLCzndtOTUlcK1n0rgHqT
/X9FtZCzZR0yoK/CWSwcGTlQL+GMOkSrM7t3Z7W6itAYSmr96qTtFnmaokQ+6JXfUeXrexZxiuXs
AML6k72qWcmYoJsMz1ihcha1e3E+H0JLDWsp6KRnlXIrxz4qe6dvTv8nJwJPmQAMFnqCj9/IJZUH
dB+I9hnXnOW8eKLta4sSi8MwDmXoc4vq2PZnrpi082vvhV2jY2FU2dU0IPPbsv2nXOftN9uBoGjY
o++gFjLfNBBb6qVCdtbB8xXJzZlIZhR4HU0CilwErVKkaimBZ2qNoUqvtMlEVLzEcpqDKA9vLd4m
qadNZjPTxYDGLy9bfhV30pwaUThb0E2RJMFRfjsiMNrIAHd6SocKIgHjuviyMun7qZ11w9poZyzy
A1JJj/TIzcH6aNkrQineW0XyEuHcO7m/zg2bByS1Q8bFcY9TbAAEPU1M0pKuO+oxikdQ+HbZT0mi
0ZgNHn2BFWi4juwE3MRZE9pho6rcTma2inYS7LXjLL9Jd8NY5EV/vsgR35hgDdekfVFZw0A1v+GC
ONccomMwO5vlVJFgJD74lLbO660O0cXNKxrR5/zoOzQB9DUyFpToHx+o0e6UY+ZE35qCtV4Djjdx
xn89C1Ca6D+sYYQtLfHekx3tceTfJzb2NilaqEIidPbji81J4m7y8gmNRUNgCE//0nWYGauaPLbo
aKOK5f8s/bMOH2NJ39Z605qX4qQxaj45SjSDS99AcBeiv2J7r36LvoH8RCu1NrKCidf1N76t6NPq
jfOl9sgxryybuFJFFrJC2v7qp1PMojTxnkuwByMc68qNyURPE/eKS7CSFy9QXeT5hMalw6bRPp0I
GMr1Zc4LAyx8erl72XV2d+2jxnZG6q8Qqo6i6z8mzrhzU044g0uV4S51r50NRkt8RWYmTpbszmcv
QDxmIzmODMUN+yXhsCMWtWCEgCJ5/SD1NB7VqBtUs+PrONMFMTBsVQQ40P0STZ/ccDA+oiJuX9w2
tI2U/4bBIbysVpsnTpKq0rvIOjQVPBsjXLyu46zFazG99Sk+EAMuDpP9DsejzQ+6v4dCjn36hD9t
/7FaLecD0BjaAGbGqULwjfDm1AO1EJy6LSnQd1TC88VGtDs0dJTpQHmZEqtEnGH91BMOcypLEW7E
IZ1HDInH2RB3yKblC4xyBcnS7CXxlPJF/Vs9MOFstRxjmDulI9OORKTu5rKpjol4t63RIx3sYlrV
h8WEPbyxB+ygHFQMD2OId0XzPCeRiLozLOX9BmHEK+SUzW5Si1QSXCvoA/dzQMWwxjGu5YeTuZtM
gH1HhK33/I6dPdAIbJUlEjZvvVJRoyI+OHDYINGA2LzKANv9wJPEHR+VOmjt9wK685PtX5PgCZFo
pcQasR4cXRoXWRbjA/JBIeclP9W6dsSbuhRijgMZAEtbAmYzBCdHkQNIB4A/8QPufsQEhDcz0+Wi
igfv0aOimJFfEjYKhCVoXc0aQ/+uN63ptBJraMrU9bpBxQf1PDq04r4JNARjy3WE1DWql2Nf0/ay
gU4+n3n5hAgW61TKW0Hj8x3/12fJcfDtHYCsx7ES3aqUnxYJNEMiAZ+8bH/seU8WXe+om4AnSZEc
/ezdMsKLO2zuHWTBpmyUhRSHc6wIcvk4E4HFjoHYicCRVpMPk5RgHvs9E7stXs//Z7PcCpozo6A0
m/JpnV+6i1sUMjhuMD1EPkrQ0WoiN/aILZulsrJUTub1OJ98FxXwymZpoj4NcfHcQm2YeN7A2xga
BRRHGLBFys+TvaPUFzuwZi7yP8y120zDkwSbEgXU0Dva5lmoV6bbAhvnC0x8P5iAw3uTpRL2V1cn
Emc+Ey5DBLWYFOODpDLLA253EAkuBH/yAzgxbYyWiir+nkzCxZRnRuQPgw7zxkVuRICx9K5PhFrd
5gt5/J/9vgoh3IEMJIB9D6RfLZeFFogFA5IgHMPJa+xCc5p6pVRSxES6omko00zwRLvjJTV/tPeN
zNfTVFv2dw66S7e/AccROIEobD92JPG4x6/V2kfoFzu0X87b5VmSyrXHl58qdTIe781/ihBTNjj1
S7hBHWs8jPzi+tYLMWIJZxekpsd5JxlctqWsqtQKWmPn5kNxIi8F+Ak9728QC9M4pSwPbnww4rp8
lNxCuqfucBduQWuY2uNMjwK8ZZFEA21tYHdsokhy8rm4+CRSkRH9lo74YjX4KoluPFuCiDp8Nby4
FctNC6PYEjRLFtKoFb614C/uOF0qtt1v1CTyhrwbPwjPZA/d2UoInYel951D24ii87eG25IPRDe7
nBu6fGvC1n1jGvc30dU7+/pVuBSkt3zMYxlNVygo3fPcr1X6e4+emcKRhbk5aLZ3BjqivMseF3vJ
yZfldu90tWAMHJNpX2l07NPafrAkjGTND+ORBP6KnEiYZVN7I+byB/bDKEaTvRdoQdNPDVtHQ00G
C5Mw5OX+zbBbSVGJdXB23NWM1qGeFs50LFS+HUnl0K5RstTucRse3EfLwPGeP48JhCgB7H6piWor
/rbKQW9WNe026fpWY+kfzASgy7Y9UVQFPZs2oo9F97xAx89dlmxRuwn5qqIu6PvMazYpxmlrtwSQ
VUC8Hhc8dCVm38QcGX18Q0DEvGpvrE6Lr9DA5zh8GHKS01Yk+F+l4vMY2rRlebBInSA9U9LquRwZ
E2Bg4JeysjphoAm9YVcrefZC6Rc6VIsgLxB8rdFPB8WUR87e/LDVQS+zZa6T7bUvRPWkq5D201Vg
LAxVZ60WNrF5SR3ObY+TldACPdyjBvbGYKib+RxSsPZMG8Wge9ys4oqNPO6tTQmOypUSV+PROXVG
PsoA4G+kaLiVRYQxkGXXcwLd2hRfofWYydB5z30pRGwhwQzgcNDokd1Fa97GG0E9oRNuq5ZUd36C
EWE+bizH4pwvTsL6rS39FFbijVc0onro3uUCuJYIYGFMAsESBzg3qLveOkYtL9rtcFnG+gLT4Lck
CQF2TA25AEUoDI+snZG/gPbCghDNbnQlL1mZ0E+JrscQHYgcWrsOZdl0YjjHsD55aWnDD5Mar3T/
EBOF2vEmB4fqY0iNsdG6pBscsPnWapGeMcnewGqnwrIOTqTzGDOtBZ/955B203WzlgFikbTge5MM
c+c3DoqBk4EAAy++mKZSdFCBGlOkj4cBF50HzjQUVC9SSFjx8qPK6lAk8J+wPZqOnPoYV/6ThCps
d/6u6Lcs1BjvZIHzACCwY1PwEgRBa4BXhR1FciKE+uSCkFo2B/xTBRjBFWML4dCNP0+j2w2PtvG7
JsXB5ThpXqVfaoQpbOcpVOnNygwtQQi07gWeWYBh+5kK9x27B3c1UEwcssE/9wXHTvs2VhygWiH9
S/iXNim0eLY1zShqWdk78Ra3rclaB32SDLU6XMZeN+t2bSur+ePWGPWEEVujAggiAuPWp1v9wglt
zoIM8wkJnIR6MqMuzsVLmriwNB3TOWghttplgxvztIxDroKR9fnYu85U0VNXZ5VE4ZpQDSXr5HMh
ABZfV3ZhwF4sayIwCGifNYAcGtAKBvBjIdpb9ik2sA1QIFTTQSpUPeVCX4Ah+9Ryqru3LG+lsGXe
I5Rb7BOCUsqs8ryQd1sarLcLLLFIVvcJRVlOFFR0+EQIxMhb00mM0n6Q9IxlsSjzxGoyD//VdUzT
egr3vNw3TDttwjG/2rbsBa/OWS6ZaWmb0UQ0Acs3TsxZJ4lvpWQ/OoO3A0DgmpruoghRzAFxwvH0
veMRWmEw+vRABwtOZK4Om3utDC4qqxRW9UubtfjtlSl5QnlGE7IJQQVaSUMQk7JGafWv9pn+82FR
DXzGg8a/XwkGnr2bLkvqBAIZYAF7dKz6ORbAmWRq2f/af91Xg8ivnskisIo4g41WdRLyskzVA79f
Xza87+vNYbWhH/Y7yrpThr13zUcphI+URM7WCwcSI0u1ebpniiKW7bHr2l/6fS+57uQCfP2dT3Os
f4lCWIcAHfiVD0XRkhOJ6dmeombcinUu//5avbIs1Rtkx+xShzPBXbZfNNeKpywk3cDLgK7nlTjF
WfFKiUJ8P3VP6KqeInsWbd4qyZ65kFCQRd44jIUqUcZF1aoSiEIKgQ2Q8YlxFC5HVvlurZQvSciv
l0ImAnxQe3Eol3dMbsY88rhh4QrssxA/sLBxTWrHAG2Di/6smRpNwQ+XjYsj4UIQaxdAQZaid5vm
rHYyDC1Jvey1NB6RnEmqU2qbazcSbWm8W+Zeb74XTd43cKsO9i6oxs9acZTaM+sxOhvc8u1KZTfO
Oj+Qpv4e8IVut4LVD5RMAXR0TzQiq/mFCdky1F1jMZKd9gPbCZuaht+/vthFOCrJpfec6CQ9JBCe
09rVA2djIO0WnGZeh3h6E4lUH7IUp0wePkyFWACqKuyWGt9QCUSdK2a1eLQDY/DyIjd0svI55QWg
zwZ58l4cETblBfxmKFplk2kAHE1FrYUW3bPSQ7yXrZO4JsYp26sEI9iERGfe82SyBqFF/BPynf4k
NPh1YSh3T37lPZSfp9Ae8NuzP0pD+MI06H4ZF4Q3+0VMu9tKK0R0sBV+5h70SitdMToQIEIhsWir
ZkLRFxL9ix5I+9JXSHjBVT4pwJrA0Ks8tR+/FEXVCJJplNkOYEwRpxzhIaQ1e1wC+9M6K6fTCHpV
xrh9MAYkJ05aO7HmLh8wjDap51DrWvDXGWabpRKvyz0BSZzaSLrpY9vPjU0xMTKiYLg88nW4PWRT
tg/fE8pMXiFENbMrtfLYbNkO6prFs45jKYK0iqRMj2tf0iCbTOHk3nqLV3HslrOJ1liu7QkrJRln
AOnTVSGbm7cZ3T2xq+4UUDRI2sPPSypWxZ1eunS+8eO+2IpFvjJw1vy92D8OVbLzLFxi8ncLrsz7
MAlNY6FFwm8C4lC6azkTl74vGlczDSgS0idpoMTbOtl9UN3sA6N3QGBXP0JLfRkKfG60TOSAUJJD
DIUGLJoibEd0rcSrCXQjE4Op7YSEduNaO2VK7IEa9xcxgHr+euUpIj80vdv01WdFKmPg8tUKIsjL
m93rbZ/fsd6JirKTIVi93qlwtgb7gUMeckqSw/2+CwG4nUjWwEjFONN2km6g9W2SJujmEMvyexnR
Gx3oFvmUcSCoju3ArNU0EqueIJl2eVFtYjtfmLRCoe7asAvxLztA7sDKeXiSVtgtYdfOdWml7V48
atx+9Ix/4b5SujfnGaKSgYR/QqSWZE2GNoWrjU9f+s+aFdxY6tpS8tXIuLp3jVRDd8UcTzSvNSRo
IJAICLdoTtnBfaGAj5TUZgouFM+GgL9GO6oeDoG6FMOlkBNezdQIeezsnpf5UmcxtrKoNdwahH4o
6RVmr748b0sSIJe7ZNxevROZJxixdJXKAjChqSvdDs6gx5QJv4Cg9fc180qeL8BHg3P5g7nZmo1Y
BTC4S1uxiq2psMvzdGF3NvF90i1/Lx45PNxOoP1I9+TgqTe1s9cLdFElAd9yxaYXhBLke+E4Xubd
IVCNDz3TeVsm6g05xg8gspGr6HdlDsv+hig2+tGlRsT31rwnTCeiBa2bl661ZZKP7c/FRdExMl14
ODLU/d8eWphtPMzeZHePZbe9oDRsdL1Wh+ORFldij03BKYFWafJZWYFvVnmvMTLnnZYxJQIuYsRF
zlP/ZYcuU5YQPVAttjDNJ7PZGPCozMEsFkuWTrexqFfRKREMx002TWJRzJe3NPMCfJrlF9dzc156
/Ne7kDTkR8EweSJYdGoMLGmuUO4/CZShFHc0IEUw0PP2cBT8tgeCYpNbx1YO1A5SsE9DWQhUOE0A
PumflawphDsX2AwLkr2Y0DrwnO5R8U6KmI+GKn/+69JgjEFxuJil3jVd0h8LavOJNl/dmMEiIoJD
MijeEJMjrTwjWW77sLw+6BOBlgBqQZeMWNEwNm8i9WQC3hEqd6pg/6ol1Nnh1R1NVdKqrbQxjDxo
cx5VPodoXha3ktof2zNnom8q2ERDwK73BFQhyaKX3aPK013+akvEjPlJonhu3IbytabBVEYJQuM5
30Kz9CXE43sknhysNOoC44xmtxL21e0c0S81WI6y5aXtHDytfq9bgq1uAtoez0ELFLI+nS9GSrhO
H1IxApiqkRN+GyrLuyakLj9OKt4Rg+ASe6u39dHi1fNj2E9kRhwYmdiB0B069zT7c59yFvsiWNTL
fP/EyOlLLWDeiuMD8rj1so7R0+GcXQTX+Mymzy/SuMSCHmL/bG5YKwoGBfkD12jeruIKW2BPcW0R
x9prurCRUUsLfh9mR2YHX56tlnrERT4RF6ihe+KrrlbQF9bR/Q+QTMNlNGAH0Psl3chGlbC4Wz5d
NYKX5DqecV3UvRh8YTXK1CEg6LXlro9ovskahOxtoDDwlZ1C18cT2KPgtA1PjXSQeVh9HGLTNvU3
4dgHAraXfys/EYaKA2Acu+U6rD3KBDYyW7VnoJMBdTKYlodkFJYkSnmB18CImBhB/H+5q1Yeo8h6
JhNLHPcYuojBKsMcjsfXKAxscXiG7PzX0r2mFzP07kJyiedrQ6xGanO8W07WvM+vf9FL+gAtCVM/
CV/a+mariqDBxUdI1vxoPPHm/SH+92/7OaCr/xjhM7dvIv/j+Sd4C+mNrEm7k45OPmPYgM9zF5AF
tFZ/9J/EXaDt7AFvow/e1kmiI1VXhR4vE7GZdLWIz3eZSYAdZDNvOPNvBexhzSRcSFs0pmDcMRO9
7PqXCALZXwcIXOyDuK7rUFQLz1yFcBwoJEXqweCDMA4TraxCAnXh1xZp2kcMeHGkv0uQ8Ou5HavO
KA2p2Bs8kHH7l2D5AwJb05qYE6miSDD4pV9MarAGLD3wJlhlA8quS1TFQG17Md6Xsj+h51xTasWL
dUIxdonWimanl2omuhA6GhNFvXde2Xh2IX5xHXKQLOe82kMBZ7Dfhxst2jArDc0xdW20iH06pEy2
MY6L8NH4RNWJ6NrtBZiI6qC5S9nLco/dRa55PnA7zBVjl4x1R9JrW8sFvxWvl196i5464H/xQaRB
3aW+9fiFwrXRrYQB789twqHYUzgE2SbxFfCvpS6sHyWhqE007QRtUE/hDGPzbQ08TANbftoV/cJ6
pUKIqx7j7ejgZHqNZVAKBcXlyXVZBlhQz9FgIZh9caitRWE3J6YOQCnm64zJtcpiX5hQMIxKsCU3
dAIrDBUq5rKuPmxwHBoLde2xFyV+SxGjRuisH1XIu3B1jF3xPRTrCvLha+Axwc1pvZc9YEfDCBCS
Ra9RM0+uEzujNI4qhWTrMkfSOAUA2su5lwmBNBrpWbmTOSrWOXw8gms0uY3w7bwysqkxCbPMj5qD
3CPrjjPORnbxVcFtr4PH/Yuu7QBSOsne3fmgRUs+l9s3Bq04t/m+x+evMo+chy3thd042n543ZWf
V4pROuKPewGwahimRHE16waUHqhoaB2YvpDVl1tCFtM1p9mmCyhWyIZfWCGZEqc/sWhgNOLkb39/
DnYYpGNka2fs+a2RMy38NoEXImLemjNOebcya1HpdUliSW62iEhL5wMMdjsdbxr8iw4F9PuO2GLD
o+20uyRvbeo+m4jkANd8zc2Zms6vqVcSX06r5RH8uVxqROuKREZPeH4NpZV/51YK81towBq1MMOj
VcrR+c7JnHW+VEohuHVfi28B0eN4riaiBi47vDTHp67MlktoRBjMCuQ+cTAFHRvbZaN6qvStlOpr
pXj25AGzduN8oWOQ/eHM99UCVdW+wP9c7sr2Y6hCmhKEPU489Z1C+jU+VQOtZDeEOQU84FxNbEVw
QxKF+4M5Q8XjahThMD2nMIHK9HDAkShSFDHY0fgROrVJ8ZfVRmjFRRX6eQbXGzHLkmJkztRk6Na/
ChLvOFSvnvCrwXXpxghp7VUDjY/bmmaTYFr1imiQqGvBVX5Am7Ko+lca+cuXz6n9Tpj3xYnUgk86
UMZCAri5iNqOKFOqfystE2MVB4bosiaFAFIXR8Rmnwnf9nYuzWIRDqDZ2YY8PaWRRvj+anaEU8CR
+QSvRfq/u2VZ+e//BwbY78S8rcWzKv37VydLxA/wwgQe8MRWIeYRSjA+qtonjoltgyIHfTpcd4+A
s3sFpq4ju4FFoY5qJpxP2lfODpHTNzRE+UakhVyeCIexZ034Ig6qAj5pNQOELQnYVJbXZwvBHbEb
IZrsy9GOIAk0PCAvMeKgdgrgrmj2O/qPoVdL30Yu18GrZwSovXJ8o5wutZMSHY1nNvk+KCfFPYht
9G+8njDxl2gqBRMFpasoC8WNNyn51z7mM4hGjzUAJh134HLUkKTRYLSlXmr02yZ9sqqPOgwqC5yQ
CEJLzXzKVwXoDevrRjA0C66ZxyWoRPIWzN0weNs0eoCmen6zQSk1WVpBu9aPdNyxVj0rKjNIks93
W/Zqr3tqO4360ujs3r7Xs4cQqYSyN3pnk/agM7xq/eIKJEX71d1QIVZm83EgVNkG+c5xHY4oE03I
MmpDDlrhTfwq/TDcgs2TfcSwDSup4s9nitKkJONtMJtv7malc2CAlZ6Iq3zJ0YgtautRsj5l2s5L
7XpKAqIyFmtM0JSrTK69ns5FxymK2nlOdAJAfTzCkX/DNYfkPt2LDlRhgXk0KeONFECSXi9NP6gB
ps5tvFAFkNbiXkIKS84dAPnFmcDEO06otw/wKiXNf1pLgp6DGvjjwlL3It9JglasosvAqDp2vMTR
NjEJ7cHba3mpY2hV2mBz8Mm6yT1vdDr7XE8MWh5HsGBdqKduO4BRJHaD57Yy9qMorPhnyqBIRreM
DZ4G5GAVkbJl7PfRFLiD7j/QdhKUFLn/0XTBdsCQvmbNZBh/9IuRYAAXQBdT7qCg0rTyGipoMjBp
abVeBLqQvLMuInTE+cm64bOBK1Uce92THWljuj8xz88Mk5aMkUCOOhe/gh6GPnP+txyUvAlywg+G
XERugnAxQsQVu3HsSR8lP2XlOEhfOGg9x3/brUxzjFzdJGwZyHXIPWUedADz7XE7/iKijxwJtBc/
unLtUft4B/pd03muyTvKeJ+Coics/ljl76dQQg4+Y4RTU75LxElvlJMk2TIJJy7914hwi5Bwljev
T2aeDrcvt0IqFfAuSWb34UsyxkY+qCCyI2OvSDZ73E/Xx2fN8Qfo05BoKowwRnj17KMw8i12We7J
0rrX/BfHyMwd2NbLFaBYBLFUAy0a73Mq2M/BIQaatxeoqxqL1RIBJvCgy5r+84zgbyjv84Dg+h2e
ztI4/ZiWFRE8xutqOYUuggbWqDffWn3+l6MEHSJvwy+nIs1EirN6tjo8AtTDP4gzMom25+g8N82z
zQOrIv2tpAD5X27FzAbx6BinfAP9rdl0fKi+VH4jc6f2roa2ORp/ujkIh5Lb+5HqLdxQwGBfgM3J
ts9ghrVUXonUnabBlu/QCdVpOtqzYazcM23oUSN4bNVcg6HOCDNUbcQhLl7ayn0IleJp/PeDp4fF
CnSgT3vfM34fXYUAO3npbZvRE0fAfyWHzzfv+Vy+RIi1de+qyVks5HDQRj77hIcdXyC8MWw3zxcu
VviovsZuntN79zCq9rW3I+/2BONCN6MpPARouTDD3pKGAoZw1KW7umTYFSUKdrHy1SG30GLhjUpr
ArSQHCNS0AZFYriSe2r77gvr1btG/zzvxBgbYClxTwpkUdOTQO4M05P7vhloZiUvbiI2nDi6httJ
W794ujivhyQMAS/o7dA/u53SN6T3dyh25fvnmzR/MyOZyMAwFYmEA9kchJQVCR87Yopv2WUYfFKM
4BhpaXdBCIlUTNxPofF2WobIoYVcXKHC42MF5NJy8JKzfHCLN15JfrCm8vQUAT7PHQw3XUZKZl/O
dkJQEkEKpffbBcahWHQbJsg7KkOuSE1wDjrtLP1ITfjDGQ0HX6h5ly8+IxPQrICTZzwJFX6cnE6v
jZqq8FG5bDk9XlZSdlsca3/QSjEn7D401pbuUYSv8GaYZ7hwu/ALF/5zS6yh2n+ftXQJD9k4mwgI
jC6sMypUP0vMjJVurfrEG8GHunE62HXOg3dBU1oEcUmaz4ZZleWfQFc1pVpjDgdwqTGhxlFtjeuI
ex84o0cusdkHfPpht/ncxF8gSjaZQHcWMXrZti4g4xXNQUxtEfbUQem4/Y7+4SDaJM4gHvqfIyhc
G7WqAeOkphhrehOMuAuv7d75sZxiP+vm2OA8wpzu2xG7iTO+yIEmWi4nh+9qDmsjPXscZ+1zr/xW
+5tG7lYRZ0u6N4mGuuZuT/H1kYGWuxVCsV6UnbUqXSty2NLmpoy7FPS42OYqaFrHiLjdFS3pliNw
NTS9g76PSfatatZPOf3VpBRj0nRoyZVJ4hzeTwBnRYmNwmKZdUesfDDtfW9ySC2TV/rPTA26WXRa
zn+bCShjF/7NUSLTxcY03/42fZsrbeIynUKszW2IIwo76coR6YOgJ7FBLlQoJMIMC/Jd3DDyWZK/
B9ejyLYL8XYiNksv75BqsKjJzc6qR/yfb43iwGKnpEz1h+rpyrmVzXzSk3y4+3/cwUG1OcI+dKtW
U8e0DZ/SjHHrWZZuZXakIaLpliwKjFsWCkzHixkQYXTr2ycHdxQEqYeWErD+95fjJZ636aRJ8dmJ
cY/VaGM1OFOkyUFFY60nbB7cJyshRfSCdKNvTk6F6k2CBEuOJxsL5Rjc1bt22JjyAptAUEXel694
gTxuhSf/ZY4S11zqCaMnRQwuj7V4zmHCE3dnefaLCQoGubD5SXy2krdlaAIeFC8C+sOkhav3mlo3
jV2IuyyBDqeKezbYcsd3qSfcXYsjsOAtqby+gXqBgYQDOn6jqHUdaFsy+XKagCzTvrhYFzA3dVrN
AMVh+4DYT8aJAJzTlfjYUNSo/4CzHA4V0V/TPZgQ7ew53zatkk0PfCwnQGEtay07Qa2XpodxDwn7
Q4NSRAcXB6i8UQuqEuQhpexIOBILhdqmHww58XA2XnsP0/xmfKbrTpPa8Y6IXIzcO1XBjUcqwnlp
OM46mT644hLBXlGgSWVco0/ZT4n/CxcMD2oLlUJg5Hrj3YBtPUgs915cuSdVs+Znms/pv9pWtwwc
jKHsZNlq2X9xmqwyJHgec+g7hlwJoFmREoMcPvoekKIUPBAIG1JZW1M4+Fq2rIJYruPrYviaJR71
QlTwxPDDFPZ77/aaLwYi8e381hX84UiVOe5qIQZqwCyNnnlWYI5famDrkmWtK9j1LfG2Ou9BEL1m
0I0dD/T4whlvGVBwx4wfsyEVCunRV0yUmzx3UK79vXUEl+cz9C7vXMB2kYg29TYY5Itj4YSqx7/8
nZ4Y4CpT587xWp2xx9IQbz+q90yNbfO5w5o4QC81sBkiwDldlik4yRFiaBkkx9L5qhBNTVMm5Qx2
ZfqBhLh3YL0mb9w6UrykBkyTfXRsVZbT2gSfL8P/MGoc77qLZxVgZriQOAffHC/OEERJf3AkfKcD
Sf7HXUnuKbwPSrrY6Qyk7gCHJI0Yf1Tc2Ekoi4otCKeDZWSCUyx4C7aZaEDHa8Xm1scTQ9C3pwxA
mGL94QHwBWEhwOJL2qkNa7tP7s9DBvTEE4iDoffV4DjkHQbOgl9Y0cK8ooScxt4E+ZyjCbliLakd
vSVebArS044xiIWu6rh+ObFWkFgu/IJzNIljbpmIzxhnyu07OIGKktLPrv/+aT9c5LMeRo3xndxc
NJStO9JvpYYTeIEpgbpMV4/BRHs1EfRbhgzqqf2EK0GIGktEHHaWYClkLu88MQqP77NdlEAMoeqN
qVdefxNu3x5UwlFSknuBytl7vomzRxidUjmlCueQANuvMxFDTy/a++LREIzYy4WX6DzBxiZRmLgP
5upnA532HX6eHRsaTOrDLAk6qAtI0ZS3wsQQ7P/sjlfgEu45BnrRvam8EDJoyOnXAqAMaqVzEcTO
fJcjk2C/xF58buia0CMVGREhcpbD1+QVGD6NLF9Fq3dPqmqeRDFRd4s6+wzPW3WQ3JcJ5VxYPxn8
/qKf+hp+CR/vkJY+sg0zr4rhoTTUx5TQ5mqDDByrFSD3g+u+rv3Okzv+gWGA7UE1vSsfQnYg3vwQ
VztcsxWa/JndnTqsSD/aJ1xlxjDNhu0buWW8b0qPfJcsVZDv/mjwAJ14fbdKxpS1l0lY5ZJvRaO6
4GGwUSmUD2dWsiWoE+H5v2mMzDCzBtkq2WeFCcnm5qjIUOdVyaS5KOi1V7rl5nB3DqfBj+JaATPz
B6ZFlpquFs/mmV+JoP5kKDmPoKffVKY8ocnBKiCO897F8x7Fum1GfXXsB0zeBUGnprrMWkk+SqiX
r80OTX0RBe4nr40twc26JzwF46lhPJmv3TZO9ZlQD6QYzzQY4UMTn8ukvduazwH50z184D57ziN6
R4lgApyr02I+fzKpajoST/tu2+3kfcYObElJJzuBAk+RQY/cEL5m3kQrDOxXPJKDeAIt+7Rrx9F3
DqlkYxo2idLjnwv8k8p1VL54gAQgC8pieXRJfNgD17qQOZFe+TcXNW6I//LjiY387uO70STFZRUA
3QIWQvAHqyyZfeOdtSr6zw2bu1QW+VTq/BN0EefMSpdl5QEp9gsHrid5A8X8AOKWN4QL8dhrwFRZ
zYjOAiCFCGIyC1K2qXdN2m7jUKA2XGk7ojnRK7ng6sAxX5Zusq4vN8Ye6ml9TmBF2mbFhITi86Dn
VnRWPjTjNFCiYLxw/Jy7IOWZ2iOm+BT5ItPxRaG4sMxFNHVpkmscxKuTiGeKlze+SfiMIutB/Bfb
fbM4W2nuNKDI5uqlsZ8lItisDvKhqX3umKtF5S9EkINr89uvsPGc9MsdJuh0Z7VrCKzhBZVSwf0J
v6FfblZH+FHUfA9stxy7KnK+UWEmK6ok/5rr0yWaYtdt1oAbkQL+2Pw3doGj7uFZJK0L2M/tgPuI
jIc/CORPa3FpMGKo3bnrFUQ08bVa9FmtUn4t2HhwaV1m3A3xxh/BpmSmSb806OI4Lyu3k54Ertpq
xFlb3KV5khHracJooDI61P32NsoSZrUmhLmT7R8kXgAMD3dYmkPQodZOEI1PaO1rLaw1IDQmr/7f
IOYazKtN4YBNutju1TSoOLRc2Carc85aHFhw4WF37x9phygxbgPLwB1xmDGI8454pF8H6o/HLN1Z
ke8XtFGYeDPnGNJChPerpSX2xXQnbRktaNe2iG2c//FKuWOsfghtbtoMu4IK3X76oDB65i0+rqFt
WlXZSy/DSbEaO9i+20iQOAquLzc41hK5jS41zUfO3qTgHrt0XQLln6rEzgYv0l3hNN736SKBUvgl
zqaUj6Sk5Ryjvehyx1hIsa68KUcIe1Bz54FXK+cquXAcDSHVp140lHUs3mlcR+WraTnadh5PhZMZ
K/u1ihvE3mRCGoFgc1YW5ldg+bb/yc5Byc+QVdo50B9vUzVS4uCA1gbOxtFhA91fPLDsTkssj99D
sitgCPxv8OfFdlPXGG4Ppss0bH1+fNZWYN4+Ljme+gINqHgrxxScCuPSfRALdTGaO0YGjy4WOY6+
dQHU7zJPFz6aDGRkkqJer1tw+CMN49IaKSTZbtza2k+nsdu+NRXPUsmGfA94EErD7lckWX5iMb+3
OP3+MsfUy0GgK+Qd1rQvHlEB7mpGxKV/HkqTkQTiWPcJdZH5ltMV03l+0yRbuzDhOKZy0gyVcDbB
ZYdPmKEueDwEKSZdXk9y+xIVPRy1k5E05HHlUcfryJCWhehZtaIPU0NgbUP+cFvAaj7sLk2SDBpj
ZicC/nmr2VexKjbV2MhiGu7IZ6w1FPS59pIcyixbg93euDCCU1IWWCNimiiikWeKJ6LVn8oJHPmV
oVTjN4Zv5oN3mK9mSynN0QFLbf77OgBxThcbHepW6p9D6GvuIJy1dkkz+TLiwrpMxCkQigMKiayi
YPm6oR1cYOPrHwNO9kKiOnxT4OlCPZwdNrLynZhlSscHduhPWHpa3UgaBa7meJneT8B1yyjWN3B7
kvpWd+EtpjTzEiB8ip/5+tqlKh2OMzqa6/CE0TMMPiCgDDcHOKHQwRattv7DWpZvLoCY2Q7femAw
7pWiaEH/BfYhRJWkWZl7jJmthiH3W2kO4O2dBRUWTmUVNF5ZTPw08Sl9wS/wCjX8tOXHLV3jIGVc
yy8wA/i/M/jNWFkwaQF+xrzf9ISyRdSbSCBN6OkjV1swByMJ1jkLmin5DjnH08TKmrlE64q4X0ti
ncRmps2PL2+umKCl3TNASpMTRslzyrNICW43+VHlxEwYZMESQMa+0vpQ3MFCz4gZF8fBx/YQQxka
ygbffcxvkUFG4BF3aJV3t5jFcOFaKejjwdaLro/k4Al4lSBeRbBcP4Qqt1eAxiJKE1Y7u4u5FP8q
JQC8Ck+qqv+6+OccB/uwcKbXg3xTvG3Noudv5gklKUnRVYBgR+x4PXHrKQ1/8+BzCYh75cDimQiu
IQudyVIotTHFmn50AFCmhTdcxFvV0VS8K5tQu5qIAemQaBVF73z5D31ZxdxDTsMXA1dmVfHiWoTq
FE1HrJB86em629TyC9WC0Xw8Z6AG7V5UktP2x9mh22O7vT1ujE4S+T8bYxZd8VHyLUvTKNHGgzpe
wP6SCVtekgv2k7dvwRFDiWF//WAuLT+Co0Fmh+b1BdXli/nJmVCUi+LY9NcSTdBIB0beGdMuJlC+
tK67PKd5QGPJmqBDmjSzKgXk/6bTH6PepNxUyWKQ4LayUujVI5jg8Qid6pxJoLZlXoIxpave8UBb
mqid7Xv1w4ZtUbGJdf5lo50P5vLXwi9Ngfor7AJpG3ty9fSeXbyNIYtfF0QrMUGXeoJD1bBCA5IU
OaRfPmJM/YBkmmZMoscrwyEhCFXOak1mav6tCJ773ogG8U68b9DAK8W8rLcRKAKkGV341g4/J/Kl
nZfjrV5OTSCaeey2LHed7bB7Iwsz5S8Qc9mt4Uw25OFme1fmHfyhBmJ70klvyA/WNIRZw31ygGWS
q9mfxC6oqaYwGsSOJIaJZXIeb3f4bFPwxjKuQluiz+9ORZSbsl+qn9k+GX1jUJQ36OiDRKwsAdX1
ZilFUL9sMfEIHZqIILCgNYx6JRd9WmneL61ZBSKp9W1yGqbShlIWFwQlrNKyXoy3lR8q9uQ//+nP
vkH0+1zomuwm2qgLy2IvSRGNjG8IVCu2WknLaR4W6f6Z5erG0vzFQr2/HKMh9awtF2uk2RVlYjDn
/kxUKcA0LUn/qVv0N1NxLt9g/6x8nLQG8h0Y50RNe3PJrJgk8/4QB13/mpghlHZpFnI7NwOCn/fV
Dh4xpybBAqDvMv8LYO4SPGlxmQd5cu2TiMJuxo2v6z6SNVuWXlDkcMGleDbRjXWN+WepfArnr0Im
zM4wYEZBlEm8gSiO4mMISOIkVtDdagt4hhiVTitTHyVTaAsCYGjvps+FkNdCc9tbx54hx3Asa9P4
ajaK8JQxPSCKgX9jqkyrgWpLJyei6TQKHarpmoWuA5Qjoo4B2fXOIyh0/g2eBCsyWeqr1+1SBAko
YxKV1lak1+GRluj42sN6Ro+dpLMnoxo8tHNkzhSaqL3j4Hm44IU5i8MyITVi8Gsj/b9lxrIMHTr2
/5HWqO2yvfSiINHE4Ugyia/hX+IoUqm+ewhzr7T9P8Km4GTqcF9PalxNG1MvqMgYmcHPtB1WIs4I
HbXepLqN4NyC7D7zVGGX1TkcdBSQeGno4MOJ7W7fJm94Ds6Xo6JW0G7UUL2+zbpTfc8XadhgnOZM
niAh+yUmeq/tIaxYPXV++RsWwqc+JsmPRiIgEVHydYjHI7KWmc3wpTKFRlck7aAjAnjfhqhW7JYg
JTxrymPjwKPIL3ub+pFC4O5ThaAulcZvpgwKHIZpTgpg+B2CbhrHIugpYI1sA64InswbP6ZMVZP+
pwHR+BkZrEbBxZ3AEhgQ7zdDE/RkB+9DcnOF2vCWhYfxhYpc0AZHGksZbOwfvDWW/gDHkXrvzXFT
vndyIyugRX+CbwmX7SOk/eOhl9ib5mvjj9ttzVeJFzWxUYQY3b1Oi5v5xnzM7gEGDK3EqmKOvI4n
0oV1dQXB4Y5DuQyEz1Zh8NT62qlGFDm0JAKWxtxpY77v3TKYvnuNs6gONWgLWW9LPT++ULko4k1T
E84swC2F2LKvSPMRY4JUmiu16w50VOyXVw+P0hfY947jpHLUmFEUZRe2j4+DoP5FbPXotss8vAjk
JMn73XM+ZaDQD/bPwD19mjhGAPlE3Lt6ySxKrrfepgHyinQgASZJxRepOOShgO6CZOY7qlrF0YMX
MyHMIVarVKBpv3L/Rd8uQePrGoC+LbPqsb2ea4zfE2To+s7fsUiqovg8IbeXJgZLkbF39lXre2+P
n1so0GlLTxz0GczvToNF52ae6ik1bktfdQfm3NWjSYw4OvRjIHyz9tTAL1t/agL8eoECwyk3ewcg
01THutARdNhJYmzUZ5beoiO9Q6oy3DOS8WiddpVybyNzPrxiax3MsjdwYracJmNeENwcBMz2r6qV
nWJHqy4W5BE0ku0uE+GKUTRvrx9oto8jaEqtAUc3BDV03IB2JuKq7Sw+VXoAamNt1PcKaLa6NbOP
aFDkomVWyf/FUn6O+CKETkdCEY7oGTiCbrP146Z9QVKTVhjhedR0//fxpfkxLChJtw23UyB4a+h2
C577QvKigC0eyrFPRQJUFGp0zWu8DXy4c4hchcxlKAqYmKtvDpppmA+mYfgBePEI29rpSbSQUFRj
U1VP4egbUa2C500v3CaWpSjuV48snBLybbLAYGjuIL7E6/RHyjfoMWYZQO4XLQY0Lb+KO0bVRGRx
KS9WG7aQRAew+Jt89j4yrElLghhk/hPbSOJb3C+EUS/jSUuqI3giPjBv8d/naba06Xgx1vpc5JCb
Z96fhzXAJ7neuNzzH3dRMhpqgd3tl0ZR4M8yaCNjWR4L/+OxobESCPmwBqdkX7WhSVahjZU57B48
iGpjcy22e6k5J4Ean76VExsF2IbB/F/YnjsnepEhnDcLtDCaRv5+mXDDS1zaWyxsEhaUiVst2Tp7
nU8R/8X0Rbwt3j9JNa1ATjBxUTgHzRXrCzw8jPER9LqMcJ6AujQU4M3GIOioIJgMRjdBsjPvxxGj
ESU5wx9KFe5eVp5owwBR9IvXNVxuOuYhL3pgzAdCbuKOST5RIHKvuHQ2b1U49tO9vzJPTwSYvsD0
ToAzKoubnwyV1BGHMNmgGHNDjAW3xDLJRJsbs5FZxxA23ChEs3D3Dt/hV/vrQt4ztH+UpFR5vnAJ
vQ6YYjCOmqd38eUgA1P9e3Z0oRmDSH612c9UPEDEkQd+Qn/dmScJbxJgHcjhgcLWkksp3jg82GJQ
IrR7gKDawBQDFs4XZQmPEbte5dsP8XQdwgQ8t0tlki+8v1ykIUYyWQlLVtFCDWh5HhWTHSTmGDaO
Q0Dw+ceuOk36I2ZyuIwXB1T3g6DZBxTpNFswmrF0swMAQj55gIyPE8ImaDifQSVLozRFbE6sw1va
LAaBh/iXg8lDotUpP4UqPmYFTcN2JpieDrGtbxNCBPfLq+agMDcmOmvwFkoHknRmSrkjcXCXQY37
Lg2GmjGzlZv5mrSLJfCPcN0eA9VJxbeNtUYA5TA3vBiWAOfZTqZJlpMYDK9G1HgO7rNjS1fnMHDj
agU4PBvqRls2XnbU6Tc4f6VdD1NzkL8vieRQKJOOobgEyoC2py4hADfW+EOcMBA5htOrrv/9B/Tq
ake3ZoLrsEwkyNd9wdkE86J5gh1rPGbC6HwRQ9Oq3r0YaYli/mP8ZgYch4YKBV6xD2wjx5QCdCAL
9M/812pPknIkAxPUoblIb9s4BTkXDIitTyiuQlEooP5tF5rjfx7TuQxaNZDhQzJOQdHp+y8AdS+H
4DcCe+8Gkd58DwD9HzKyd21vmXcPC+eOw/rXF31ZndldlwL9FcOhdwAlY/5GbGm44dMUOAGPkKrw
zN7de3dIUEEvmDJ64oEiSYkksNTR4/7rLEBo7q14OpKmp/2smlQjuSQ/xOkn5p2nltpg0lb5P935
DqG6nYNW/eOD6XoPaBr/PG9JxBLLynGrIXI908dXmMevszeM9z9rN/3F03/b4tiEFeselDEZ1gqD
Sf2bMJGCnzmhWA+1L4Qcmli+We3+C8MIvA/1jLkryJpLsARHevyOFV6Sr3XAZKRvh0RP6lH8Yrzg
x1hG+afp5Exlggp8TsTvbRe9B9NZdXrwtkQQhaTLcGbsQdAgM96XXGvpoh1YSQrgId775VSs8wPE
uSuXiOnIMuR1gU9nL68wK2SK57AtBlsOeUQALjfcSSbh8Sek3w24YftSUpFwSrUu81473JkF9kBT
OaHWTi/QXUdAL28uGBLNxo+6dmjRaYbDh5z3w3s8I4/5kjxLADE6y7y1IxctTREyP8+I0b8fZvq7
vVgvre/2vnrqvj6W47o02EXDqIKoX9mClcTON7H3NzCe0OZnSjG+V5gOqMfnwQGPZNp2fXHBA4m3
f6BFp92KGIicpoM0VcIYbiKCqqUVa2kHdiYqBgPHb083MRIIIyfXcoAbYcrh9uJC56bHnk7GKGuw
RUCcKxj+WpVPbjE3gCZTgsty70z6Thr7bLkbImJWU3plgpi8BgjOm0e+ql3105/Y8z63sJ8vN10/
9hPapgbIWGxjyRln3Y04ItegTK+JT23n5ArLjFYYNAsCA/Y3Bnae29LwZZ84zA9kXFgmlu3WzoU4
TXXw52sdmX8SwrcCjRux4ctinEqCblpFBeqCjosvT/rfotm49vgsJvBN1MXJoVpMRnlDolvpPfX/
viRl4dITcqb3pmaaCFYqHptqof5KcidvQVR8v0AEcFJZY4CRb7MqRSzsL/uXlG2rRMVy9PzaSQGD
J+YRT99+wxOWb2AmBQ3UN+r6c4W5+UYBL7M3xCnR0dzCQs1iVxnh3IFWaipfH90hNYQS34OkWASr
p+rYxVY3CNc+4Vg6tofpKmJTanF/CDXlJipweLeT3Z95eikckGTg8n2VOlUERwpC9Hp9lW8rvv1m
SMEwT2S7cfVCigWB3UoFJnY9wG9ikX8q3nzJzRcEHf1kJGspzvGUZ/jY/Uzz6vOkp42eg4jVzrUW
GEbQUUicCG1J0DELLpofczv9I6Uq6IzH2FE4qhpOnkzXlzNxvUAH/kHv6J2WEmXRObVFsO9QB/Mz
nzICaq90AiD7LH8yUz9UdQwDsS69Wdme+2+AMEneMyGDC0VHWsZmM6LglR5hZeoR9Jbr+5VLtbwb
CFzUVkQm20EEXmpJ0dedAL9Qkt1fehLRbL2rCXAybFgslk6VEsaDXHCGDTU0NCsbTlneosEkRTzA
YvbaI6WLtq4yMAIy5Toxvni6mU6OnCJ+4jSjdgVL4wYKuZv78EZBBj3Ylt/BdkkBQS2TPMHBQdTc
li6GRhl3mP6Qohtu3HSKileSjeafUb5tlbbZPIFyxsJ4nrDmtxRbd1joPb1WAN+wDcFgTRuRbujU
b7Padx9lJDW4lo0Cve+7tZrlbLVzdxRfFaUM1l7GQsNtq2FZIfxw9TDSvJJCwxqCLn1Sr6ToosG7
/f7cr/S8YFbjy3RhMfP3mLd6jvomrL71LgnZjJM8ww1gBMx6im8O6Pbea7Dv01HDfZnoTuiU3h4U
dsJvayTJZhXOBiKFPZo5bwAfMtb5mIlBerJAR5RCl8V1CYRh3sWz/oszfFtT39uvSxZ7Vbc8CI7p
PKXrPOQ18IoPqbPD7zkVQIS/IuZzqY8W+dKLB3Kdo3ix+uuCRDyHwp8sECWZQiXMLV3Y2W6X0kVE
GoQvksOWNL8I0TEuHAhQX6cyGVrGIcyd5g2t9WWwq8ygxuwL7cgPbGXir5gmcurXOZ8tdmmUEWKF
wQxCc1vt2G0WxTVQjBZfc+ktjAFy4mchJ1LyOUwSY9IVmvOublg8vu0jY6oAjBc9Ao7kZ3PhLub+
bwnCytYFJnUfAHZS6CSZiUicx16ivGQWGmxkNbReL+KliPTBx0LPtSyLyr9PEOpEmqZVee6g1pqK
bRbiUm4De9MW8/m58EcNFNIKORntF4rquDduxVEd8oMwIBhDMOp1qyY1uNpwNkOLNXjnHX0mFrLA
biY23WgffjAia8FSIXUj6J4OoShFdlXdOQhEU1O1KXstJsHAsXzIndo9Gc87I7TUG0VhITxdgFaE
/cq0Fw6uKxGOs4rP/ajNM0nJHnbiQI5C7JRB2GSmWhXtJCm6mSHjtr4qLHrdQUpqL54+/ZwK9zD4
or0mjUxtjt6PYMC00Wgw50+SZEITNYwUhZM3uXgzopZbpn8oMNWOSioNEIlVe+MkYOuv44e1ubz2
ft5NNg/aH8DaEnO0QeMOHn64aN8/CIUfvfB5pqE2orn1sFqsq3bh/+DOH9vsw5yUjpK5hQ/qJXie
ScMIVT9u6Si5g3cDbk/1xoWzbqSRoICyyayzln3nHx4UJfP0X7nhyx6RrQkIFWmzwVdhR0wIZwNK
rmnxrgCj1U+2hLKtqBm6nB879IK50Sa8tKBLsrNuu/qwfC0q2k/WnUBEIRFy19jq4DVjm2MfaZxG
rVHbflrYLz9sPo4MtrcXL7hQXu6KnTy09u+x3UNfiM8z6WmOBxWRcOHq5D06JXCvG3oVAraCYLh+
ZRTDNzSSU89w3gRlVDv721xpuF6/Za62ppf6hKpmGLBtykS2LfEfm0xCO6UOIVLxMXMU1ynjkjP0
+Tt02Mn2Pbum+85F527gzq06Ydsuvv/8jM3EO0vtbQIKpFKayNNoPaICsyhwD0xJu+fA50htzzqf
pBritppCd/imJc9CFzev/5dBEdXOX+fDhJJC7fuET6XHQLA+OenJ9YgjKN67PCg1Hd05oquidL4p
atY23t7v4BMW2yCWKiKqiuoY04Ul2O+zQH93/FNVhpgNAjkymBf2Nq73s9GdKXFX1F+vX5PF3nEN
7p/lwsDA5hdbp1fi5EYmC4gJn+jLn2sC6p162q9e8AJnOUWBp+dySU8dDgskqIOTvTkBoVrEqAk7
wCtgUjOL3U45mcFDA78EC7IvNUga/MeH5taQAbefje11iBRaiP+44OmnSBzDg4MdEmB57hsO4I2y
al3mkK2eGUoc+UXYzdCg+t6ERho6yrzccQQeeWp1aCuIJPv+aA2AjJEP8Ck4fbmRJFGC/2XLZ9le
6CwZn86x3Emon65eijV4DwPWti7Gn4ZXDdZwKYfPTuDHbvUEOrGlQu2ED7HVq59dBRuEVzqxfNoS
AoM+FH/LS/2T4V0AeZriwdtHXOkTxgQk/uxDGN5QpO4scjrjiEOmTxtbXsHSjhWanRGA52qLjtAy
qmTM6E/0fu6GXRHYtPHZWonZk4SdjEp4YDpmhXJwg6s7t4IgHe80RX/L2JTOwFfaPmwr30U+3G3j
dJz8rtlJLsY3CyrE8TxmxlLFhMRqiZzu4EasDZROUcAtgQpT87WSnH5OhXUFm7oHiQlJAGWeQt33
BqtRII9xZXTymBILqH0304jqLUYfpyDR61CXo0nkgHrI1gcYTyx2vuoxRlz2BUAfxLUGiJQXSyfJ
TKPkzzQ8osdee+a65x8AZmWz8h2VkLd2VWnZIIg4lCzcVvie/nRerhsDccJx5F7Qk6qc/4N3N8Yg
0eW3Aq72K+YlsluD7/Z2gOEJ3ezp/E7Gi/ZFnhGS9t2Gjvf67UGp8bhiR3vHSaZphAUZgGnH0/tH
lF765KmZnfXwIcXPEJBegK0yIvZavbS1LRI64IEFqfm1/IQSjzkL3l3oY5ZGaz6+LLxOeucQOj8U
Pe8zELrzA1XivSu4euQ793AmVTECiyRHdychC84APuQQCzvAOz2IyKlJJ2fu1gUt3/p/YKadrkBx
PPa7+sTPd4Xu7VS8SPGGjk2jCLVxpn/hXWDxRgk/KFCy763UNF3U/sVxbscZ6AVz6bBKFearH8Kn
t3nDd0R+ucQkX4dg/IICDgQMz/KBpYSO2Pv7PY1uoAPdgoW6akzWoFDIbZde54NvWceuHG0FTQa4
xFGVOGkHQE+z4wAhs1/1+0ggiJ8B+rIMcNON0gORyu2DZFa7xbdrk0V81Fuxgu9ay5uM2yCR2v2b
ssLStjy/5Zwgt3ZGtBX8AJnMdVlHlr/eiYVrKLigmbuNOsm45W778zsYBHwTVlb7juqYH6gx+PXJ
wupjxzn7jERiuPi9JJtN4F/4rsq3OBbRvwApYfrOU1aVi5mQhdlv5J8PwIZuFzYHFt1XrGRkMHrB
JOBCeXxWVy+igK3kDog2QqQRBEGnBWgQZCfG2jJBPjkXAUpi9krAhpP0gyoKaVvRLATWnfBrUVsD
uNshIcobjrqRI4QpmK9HGJN/Y1Yj0prrHHYoNHt41uu43mHUx+uROG79IiRPzpFsD2QWXn1PsLaL
iyMbNGAQxlx60TafpJdYMNygWuxxW7LGaTMBiO1qduhwVuMYw+lL+tLnA7cZidhOE91IzHxXZJ9H
xYrESG/XcNHNC5dD00ZFV82OmPIHG4hnNUtHr6eDHmmMGrSS+tZ0tAVS19++z5pzsKeBr2fFOXJn
D8R359ISNOWHqc4ZDhw3PRH755srpJqdPTjE8/+mKQ8kcUe4LzE371KY7PtzCsARhQ37j8UuIR2D
XVNBW2jSZTRUpzKAR6+iqJ3TXdiIND4guSqTa4VmO8z8WZTkO/wfq2OW2PvaQJja88+TStLzEPcY
a+tUS3cQhNqWcHnvNIEKhiaJdC7W87hQ1zXF/WuDROosErNzXZhUoYSrp65moTQntw+wGyz2iIYK
j+/hm2I4frV79MOVoyVBwYrLvuGHzTw3zLkMZOgDoaGzSMK31D5iyygdn9+xt0TuLqTPZCL6sGoZ
I3BPP17It/dHaJrpO6/XAqcim0jRhKB5yCf9VIYR969D2e6j8XNvPEnp/Ki0IN8Uv3JeaRUQJABR
TsqJ8VsDDSsRN+5kgAuGLZoktbKLxh3BYW5xq96uqilKAhDhdklqKg1dICA/3XSrG4eycNB4Np6u
j5OWCGpAOjlKF0axdhjOSrBo5/G4vYeBz0dcRHEBG1DmNbUxUfU562xuuBkVTCTkcAYYCJyJwvKQ
Pkl+2FRMjRaTInF7jrv8byTD4vKtSBF5Qb4NBhLN1AvlfT4UXBjcvYbuP6NqOBN2x5OpQEBGFGNm
XhpSyohzpImGN2tzEMvPnq3nCTGQWLUcXmIaT1cPQZMlD2nLFL5y9Cplw9eGGxiI+HAnO6kbBqvz
ntocgMfDmSn01htroVnaf5EzOlT1exB3ulhGWqW4NHKghYGKuxK05FflccndEwWZPMW7x0FhyPv8
5YOlM9jMMEnpuMsloqqxt05NftQO4zUt/9yBSYMM/0+OwfXv67QKX6EY2P6Hf98aBIUraCh8gaFt
ojGuVN7ylyIBxFx/ADXzHliWcmEgbaf2v4TrKoe9LHKT22CoRFZzIdutG3r3dDWrinS5h4ve0zCO
dsdsuWEpcwBN8JQNRqZrH9iqpsPZrRUD7LCftV9EyayW7Iw7a2ZLWEPBl2+k+DP7OoeJW6hbYtri
yRTjiSgvG8Mpw8U6/yPkI7FgRQvQ2s/atfmDJFrhemfXtHk/gxmoZCXt5sEK9OoYMS1EaM8BpveZ
R9/gIZ+ktoHJzYoszuEJgNPOEKobREMac6s+7d15r205sUyKwS1KSz69m0glXjXGnPuW0xmUWWLr
1fNo4qWxDVYFfzK8zOxD2AMG5+UA97PEtS/W8MeLASgVcu6suTD25UIgFlUlTzHZJWyLuBPcMbZ+
6RKcvK2UhkCGNnDa3TJMnkz/rMoWGzGQ+COPRw91bCv59qUyppVTtOvO8VKEJIGjIU6YwNFNhFS6
MYYbV6Gl2o453PptedlB1L/z+lIaoasFb5ZxhA2c532Va/3jQN/0GH9Zkll1r48tqaoIs3yf9tKG
TReL0V6etVB42S05UPPiNHP/8Fu36ssu7G8v3vE6DXHJ9TojTML3Zr1N7rVYjYtaWOZOxdKrtRw9
fD8rDmX92JHtlGI8Y8QobwgHRJ8Ej/ERVoUSopEVEGh5No3PoYyggHtoUDIsU+eKvfj8Ig1bCuJ4
AZnutSYVd2eyseG7pO35qWjIeWpEJGliUH/YR2BhuKHmg+6T4YWf/DUfRWIl5Vzx7/O9OsJ2LdtI
cebrNgWTWgEQq7NXLLhsWPdVHoWgYL8b7sHS+pqaoWPcneQ+6SlkRPRrnbpJ6voYELIwWDfn2q8v
unTnE0NQfjyGA5QJMTRJCY9IpI6Q+Yho4/L5oi/8cwvob6HTBunAj/MTY6BqjtV6BHO4zy5w3gRM
Tg1csDtTcg4KpudqtTKisxxwIRDcHQX6/xbvoVLkqjXrOD2tH32LZvkiOYBykAz7KJAoAdy4+iI4
cV5GtkHorigZAlxbYpQeoIWZOQc5X2JXmWukficRb1FpDuOGbXudazB24WLIXvKIMHyY152LnO8P
ZPOASeXybqDC15WB8Jc9B7zzMx7N314SgscUOwx5PzB57igxduuQmjJ4T3dDn1eGjwPQfoWugRmo
kTgz0Lgw7pVMgsSRNGvV61WNlMvWYyF9MllkOBySUp0eTMNkiO/DFVB6fB8bg/diwN99XgnqBsuN
LH7llSFFMhgRiWaSW/xPdWFdlJI1FaKIihKcJvGBljuKEkNMbViL8+6bYljdZBcZqeFhPPdPd45J
z+x6GV+iLyWxs/C77menVhZCY6TQ6TCDyMbIA2l+wxgxkPIkDx0wQYQP0GM1C60AGiZySaMAqNhq
gUEG0VA0hk9L655oI9iQmoM8RQi7yGnxfRQnj7UhOmRO1869PM32Yzp96j69jLdQiRq5c/FJs1cO
YynmjONBuWqbVWqoWa8gvp95rhU6Cqs90kBtx0VvK90SyK9iOt6QhLBotAZCSi4vIev+L0q6YXVq
986r2NXDaZaCZRxADnDuYzIkN751pA+u5T68/Wvxafrr7dXy5f3lyuJOQUDaqVKAwSEpQHW6D93T
15DPW67qmsYaO1UPsTEuEPYWx5wDsjJ1DlpV8UhSGUZ7++3hMK2T38rJu8orDWHhS8QqRZ/XbaDv
bDv39bv1w4YDKX2gAVl5DcO+QrFTnpE41cT/vEmrWRpzaAK7/WHEp4jrObsIiBzuNImEe3DJ5Q0f
lQh73PRtrlsXx32q2343Ud4RO9CS+Zak7uVrbCLFHpdRxOHhJuSS9SJvC8pbgzklXXIHHgM0LZYR
XGaEyX3X9Emq/AF8i1gnrchMETSAjQg4AblUgsep9ykN0FTIo8+blCbd0uF44iDILB0I4fdtRQox
uPk/fSS7NQrLb6iKJa40W9BrdEtHIclb2I9hhec5KmyHiqhTKK3LJqMm9Um8beFnbOMnF376+NhF
0PrfbZrn8BQ7ev1KWgK37IH6DPYRFkXg74mdMnnJhhbrunPvMAfT8svKFd0iOv++dpwzwxw+H9yW
b/e3y64zhLA5jTg5Yv8n9BFF5cEhYt8IONXLpXv2oTrv71dNhKWK7W6ianctZMxGPDTitngBV6NT
WjVh/lKeRUgpVJq9qb1kb9TLIgwY+zEWH9nogtN0Wt05pOqha5QvzKqtH8IseSYfqonBkH/BzsK7
H7b4wzs+lyONiIKd+XMvKbLa8hkp7XJ0B/sRhTXPu+yfM+mgDc6BeXxzfrVEore39y1y3WMizWqz
WYD0d2ZbhYcSJ3f7ASD9+0aaX/BtfugKhv9BaU+Z4yYpPcJ7vWDFCKnGaZlBhAJoeOaF3/GZ+uP9
kT+qyPWK0BJeB07gVBZewvDe2h8uXhtKUU4sjWn7o2TsqL2qZkJyE/ABMrOi94Qly6kdQrwRgq94
mo4WtXDHJ8qyBy48dZ4IbwUhE9M2ZoNkV7oigDvXRqFkWbl1PTKlt1MueSg4kfZW+E71/R8ICdPh
0gjGv0TBH1f81UHZ/jAUZHP/2GS9DlOhL9xjp9B2SONqbbNvkvrPIvX4rdQBjC1H0f1I0SJI6kVf
ZlYdCLDN/B/xvrmnogZWvLSXw9e2noDM+R2m+wytXjvwTTXjgqTxhUMTTz04XXGF8ISMaZHgttv/
C99spOSXlljbPCQnoRaXXhWOfkD8qoqEldghDGuYiWL6whgDSjdQtF7P6R4hqOru3uqAKtd8H2Sw
5mQA/R3zia9TVp1wIsMFH3QkosexihHnzsHtMhYL9bEvKSY/KmzSnb8w2N9jmQUSp55XMP3Xx4Rn
bgKLYRsItg6nJgzTM6D6C0E/lWJlpnh3GhF7ZEsBntBbn9uwerT/7QiQs2nIZKaCReHlQmOlSekU
c3eKdOejj3Qs5WJD12lPEv1nrMCea9loyRLlGjW7PDFEmdOnDcL49Gg1KhcUgi/80tHsZUhRixnp
pYRz+ZGHc0OG09dlP7Bcih4adpvvHIXac0aos8EkTquJXJX/joA5AScgyCs/6nUy5+IZDI9Yge0N
BYnT4ugmWMCbygTDzBP1xRddRpEgxNHE5tQkkuBjCYKg8W7BxrhuUFORAsuCR3p8/bf+b45xOj8E
0qYD1jvLysEFbiHFGsANuOlK9OQXocR7Pav4WSSZ5KhyW+13Tv9A4DlPWndRu8o4YZAT0OnTCmxT
f5cAGfmHIyVRFF9/8Wp/9UqGUkmYxGGWdwz4G6joNFnwg71m3BfaIkSU7uOfmv4NDXqcQ1NZEQia
hwRw19ZX0yXPRGagg13QE4Kb0wLuz23KRwBdG9yBoH5nvOwqxVzAKIWcKENiaNSVLEoyH8Hqzycf
FfhQZVw2VX9hOhkUi8q9HZINqhAhPW5b5BHQTGrgzIROcJJhfPp2bnb9Og5p8nDmAr+9XM159Aw9
leoF/xu28pwrEZy8FyYHi6yoeUEmW/yXk4AtLP1Ps++L5Ml14xxdRgEeSczMfTgdIhUrAvcBUS9X
raykJLS1RjFolRcBC9Wrl23Z0uoH1GzPuZQJ65P4P7sG/mnJNwsv//b5fHdaSCzJ2yCXufhTBVO6
RFQVpN2T5lFttm/5H4q7E7d7BFlwlVCsCkSDdC88bAfUlNp7yo8iZWAydCeb+7+14M4wPoLcGi5o
TOw/yYFECJ8u/KJOqOqPzqRK4qCJmZo0qytFd8wP6ocdMaJSlS9Jvkf2TOKvpgyja8DMpGZrj/al
KuW7zs+GmcB6dfszEqqC9+kiLX49WRCtPhe5EaSRTWosOxN5muvLU61Zo9I7evlOaoLWLKYiyr6F
1nT0nurd6SwOedPVw/98v6MLjzDJiQE2EujOo7e9n1a3JHQypDUcser15RbVffhb+WbEbbdrT8F+
TEheyxsEmwj3Nl3CQsg6ow21Exn4OsbFkNsaedt91d4ZEl/hWF8fRRsvDKllqMnsK5ODMYm5Sf7V
0HafbhjNX2VzfGxulXai3kr18vP+PbC4m/g/ZKPEYM9uSclTcg0g8sAzrkOWYQKECXNDMY/2RA8K
TH8cbd5io9PE257b5K6sCQX8TpVdxPLkEnv5zRanG05S3pNrKfDEBZFKLei2wyKljJikF+Dy5CsW
u/AZj2nj/2niWIiu8CPptw3D/OJqxltoO08LHTqptw71cMJxybu3eQJeHgLKEwjAVKsWK67ll4Xg
JX5mDJQ0dr4Rx6WSNCt9hxktEV8jzO2bjCi6VP5X1iH6orNknkuKLEglCEp4PfNizUdlmD1lKWo6
6HzT6sawserr67htDHnH7eYJyuJ7fwJVqeoXPrkX2AVc13vvLwPDu75DA8DQDetAUY2HOvHIOV4i
emmkWdDWpDUd2XbNDu661DoT8co2wGxTb2CegNX3GJesyBeZGXhyQZWIWkdBt9/wKuYu0JxYx0k8
L4BnwqTucEkVbZkwLMkRR5Ujrg9rSylub0UYdPXNb61P+jcm/50AOsAEBU4g0F1gc9zh/UCgVeR1
RPy3CHg0TA1AAXFun6+QeDHEQpBTE0o7QT3/U2w/ruWDdqWu0+VaLtgvzjoIpKIE/BQLGa3ek7IC
mx0iRHX0dCb3RTWSLDAP5ELy1tFHc6Rg5XcSXAUVsUDRC/ko5W5DUwfIGBhlvmUawYsCN4amBOWE
RiLr2XDxnGgSwvWAwAUFWMT3AYwApo5MkIwt6sIqIe1eBsCGRUdJqYENhvmmvTau4+VnG5UQl21I
w6gb5g/AoyROHJGhYGzJL7qk6IEjXToPHRw5mTTl87gUfVLbFO28Es4ISKjK3eoj9f0vmCV0LcCN
ViFE3WioQObP5Zt6HR/vHQhZs5AfExSzdyYI/D1OH4chDsb6YsA2579/L4lGXarzd5pggYIpX7b1
fiuj0JZhqT2K+P534NwOLXIggVfdINtmi23LX5WpWxJmBQ+kCplIW9xoI91xyWa99+WJR5Uzslk9
b7vh/3pJrqD9BPq2wcC0NsxSWiOGBDGhfRq3l7LOISmtmZ8d6HBFhPW0snxwGt6zqWsCHkDZ8QbZ
/nFsTTx0mf/JN8hAt2Ro/QNyAnJMMNC+1k/YuPuGwn5DQzJoqXG1ng8erseWaVNNd20RzKiYp4m2
r5ugdfGw9DGwXZ3bGmncqPaeacNzJbsGUqXhSu7E7tfHsyxA6vwVPAn36NKW2v2Fy1hg6jVif37p
DjyAWd9MMgVeta2Us8LOz6tZyxMhuN/Ui5CWNVF3FlcpaZFTccND8W3UrcZegUaJLO24HPOCfQUw
bQKesmbhLffOg1DCidXV1Sra2atAU0vGa3+AdU0wvUKwZrQpCw7UiEHinVcr0zfW8j33Ss1ri7NH
fpIZWu6rON8qvlqokhEdA+PW23HSnb2kE2AOgCtXEBhhogUUC3ahOuqCAWBMLx5o3kSxjNPwDkG5
1SqLZBFbWR+xSBil8jZQzTj2l/RPy2xagRoJG6jU6VfCWlnrShIfTh6+bYu8yXTnlwKNQGh4yNJ3
v/GH4MPvM0aXnbDObR9mzNBGtgLSq5YoYu53W/fczp7/NvvhyeF+dimSyZ/CMo6Uz/H2hxLytcLN
+jz8bH/qUSi4h7MD9QAZ4hQEh+hLRxcFzidq9hXgsEp7Qyb2XWcAk6lxhNuEtLA8wIbewKKQKdQP
8WStSZwHmgR5/a1TGN7CZ50mqjUvRso4b1vvgpYaYu4nFVkGZGFy7PoplcVsOfh6m6fTgqM6LkVC
ub6OvGtT8A1XHzNUdLISjMWhjuy4gIiTcsSjUxUFuI5hd2YmY1Vi9FBeztnIWYSjmMUKI1tjawBc
HrlOkZ0hLKlj2KY6n4VOQ3ooa6tvJWC8YHzeVa5khHAVj59pg8hdQBNfj5FqDeuyDbl8NWen5xQQ
9eJCDkEnWa+JJtFfcf9h6zIpkn6KlnfYJeOuL7GjE04ivrApuMW5/iO8TVLsZ5ypUwdJSq+5TicE
Go3trQ1IW4tFlXd+sEihaxet1AWJCFTlM7vLPaAgg58c5JPWy4Im/gDDFNWge0TUfhjKaKAXo15p
9K5ddMGgIX4/g8/hDcD1Dk8WLN/zdwyOTOPp3YPDSnV3hqCyl+oTzZYI5wjMhglf3+5w9uHyztSF
e1TAu1j4mASQrNxT0j00+OdizQu9xsPFHOoOIX1YzHbPIB4BWaafqC5K9KXRqlVXULayv8744i6Q
JrogvTTgdXskdp8jzrpc8DHZqgsUp3/bZOTiI2kRvBdmMFo4yOX4EcWd+vYMsY+PCASB+HaV/cZr
x5a8PVUirUeYkvAmhFd3IwV2lbQHHjdEo/an072UiToM7WyRJ4A2Uz94WWacfLmy8LGNFI7U6dVE
RAgEiKUvaHr+hpi9jeHm7ItOBtDz9+bT3o2AgYSbgw6ET3ma+aP2VmUPv4FFghx18XhsZIuhVBvH
5bpx8o/0Qu03Ojuc4lOoZSNKbZGfMqQeMDkyU/W7IAIgU/K2a0/55ogyZC8oFhDSZo34erg5CmC3
BXMWMBzlmwDmGYsx7Kgr527D0E2j/YWzLrVh0qR7nP22+HmOEnaBdmZrYArcj6mitcxnvUpwVgmV
m2Pjv3E4cg5K2NW35xhBZYxqsJoJKrP8lkmvY4MbZfeH4/O36HBi95cJwyi/kqYgwkYLjWNjISy/
+kvtDcJgtdz8zDq3H1Y7YnCSlLtKJ3lZXXbYBp73HvoFYIEwsd1Y5F76nqRZeTMnjqZ5rGui/3xR
W0yv1/2iHI8qQX4E0Ed9aihUKf/l1UHPL3Yxfg4bpuF97OPp9acJNq2CyMOxfX32lA2d6jm8sM5H
ZjXIQ3wq/r8BiKyLhw9CtQ/ECPpBSWU0NUwin8Q8+59yEeV1bdy+i0zRQDYOMKdY5q3xqKtLnta7
5KYiMN911jj2OIbd0lMhCCVhKlEGajjzVTOHEJk8oCAZqtp0j2GXPAW0idC2z3cUE+FbspcFDlFb
n5BHbXXsVIa9fXVPtE1wF7RzqfyORNGIhy3FzlOIbBeofaioSbB7Sob5b+Vams8nIOmNftwZZl33
jT8mpARZbk5EmIwYdm4lT9QFOEstHZN6BX2mwu6aNg/xafJsKrxlSlwFisxOFlbhXoXrJYJywR0z
k8dTWINtJZzoQSCya0lj4UIc4aLDVc96O06xIOfJhbm5qU0aSO2rd7M4li7TpFkxytkJi+UPGg87
ILpZrm/hC9qDafhnskQLMa06/vZNVucHG9PrdFMxqezR6Kj+RSl9Eg+9fQO0YEIkeAUliW0YMh++
47Dt69j2+EnOBOYkaBQLfzSzdXy65jmAuitJwa3LRBJEG7Knr01oZyM1Zlzh6ZwcnZU0OdKI1lux
1zzHTrZa6lb8mWJSToFWqXoDMzlvRAzPDeWxlMDHz1tUSxgyyLqE129iv7ZJiP7LVVexia7PK7wC
/q7kSOABgKGg8q6ywcyQycn8ZmZqXjmlM4mr2DH90ibEI8eV2o0chr07edFepDxGDrAXnl78LC3O
m43Z8Ge/EIGhMnYefpp6VGEzIzN6qEeFG8sJ9EubGJ0CMI0TxNvkBV31Ot6TriLFjoGjjqzLcbRi
qwbAiMggfYIvjHMGVzue5Sm3WS2hcrmhp9Xja7pEmdTitfhtLCcHJiMBj1FzANbchHI1OPuWsD/o
zxVSsDeBA3KqaEoej4eZ8ZJrxWdqN9UOK8l/BsJYkC6dfeV9u4psACcOMFBqqd0g00uTgVE+Rw75
es4FHrlH6zvpepM7NLj0sLHG0aCjMVSBOLUSYYHyuWIoyQukPigv/DX8zYh2LBZ5h/HSR8QjJTIS
3WR2ZZ4UB7gXeSNhkK8yP1XZbDSeNXpKU1/ZGimtIvaGk9RjTLOoNs1ICBwmV3bRWpc0p/+Cp9vS
8pcEtp1r3U7mwPD/ty3ym7C4El5tBLG55pTB4Wrv3yL+yC6J8ZYnBgLpwrLl5KW8yyjoT92x0hVS
dOydwRtpcqy7e/pShMQWeLwr8KuKXsqMxBaOYenUuwdQZPCUfCshWU9slrzf6Wv03dzm9t/N4lud
4KiBDhwBLjpch+H6ISURXB9uJ/qjKDmGyzRSnzLoC676ZsVaaYucEvobdDHf/IDuKUnnr4PAdKKz
bpQrcAXO6iqKYLFoKXf/Y+Hb7Am9X1C+9ZATmna09L60MYn2Wf3tYTuaWVOWMYxqsJKvjdMc6tYm
9dtXKrPPKd8ul4It6E+HbeKjmL7UpCd2Ksfyzr3JyJfDM6xnwwztpffASsDTt8p8JdpV+V2cHsqm
r1lMc7ysOpS+gaFy+mn3BCtJH6TuMRz614js2DN+l1Bdk2G3Qwf3fXGggMWGOTf99pSGeBeiij3g
bdTK1McM8GZKWJQBzEizk/H1ImcI4zdGWVZ48DmFWq1/4HmV7W+cmqzkL7gymhDHqlqpWjW1Lu80
710nwcCDo7L9+HMCbWUJsjyg6lEPP9AlT1OjgSXik+YiH4JevioGfJkl/3aUTtgS7cB4XtdDfdxk
K6M2qz9uZedzG+IoP6lXfGvdidCAGabieVujvqEnML8rPcZaUl4He4rAxuiYCMpAOraM1HDp9oTK
w2CMhWL2HSXtK1rRLV3Do92UJDoe3Dcb6RQPmX3w8KCWGmx4fjIIYhS3JgxvfKBtioMbEMZhL38K
CT9uArA8v/tJtiU2b9EYnnYQq966WwNqu+1g+kr+7tdQVqFq11JB3UmWhPw9jD6DBezzZTyebA8k
EL/gnJli5gqULRCZWjcQ50bIGtr1T8m1xnezPq7yNwSBilnnYHbfIyYiK3afBed8437ylHV6o6E+
db4kuCKtZj01SW9EToscw1tqS93vefnxF0s4hEqpXeX2c6Xua+EzVhjRVKvzvBPFgtsgpBSNjtys
okZD2kEpwZKvLomGKBlMD3orAXIg1KRVRxCOyxWCRaGmIO9UbblSLS/88anUCbUquxS7PEiipLdC
V0JmwweTunZpkVyAUC4vVkgknEDaxmghoM8F4lQaJKkhRIH+1Hx7lDyYHjoqC34Nsaa3wsAGmFJh
LNUPPOYdC3zryeqMhNCY0t1A6gKWiJpWlBaxLt3xQHtE+D9e7YuDVLxfBE+KwOhU2VQ9rJhZpEXd
8qxRs+IJYt/AtUSMvZhmEoOv0Vx+y0J57e4seA368Fw17xUPgyFl6g0QDX3G0QXELfIxQ1Lk9Lsp
9hMnZTXO8+AkjHUophIaQHmWQ6PIGmS3s7xDljwVBhgpd0hlwKMkvtJEuXz/FeDetTY3cOrRyaUv
wzeCEEU0zeujkg/6g9oVc+ajuQjjRgwUbpoegb5FIwbr0yY8b8BNGOhHRe3ydiHxVUaceUnKECPr
JaOTupEGHL42mb/kQqGlB+oKNzw5gEXdl+Oc4Qi27c+2/LuC9l2DK9UU+IsIK6HWWPp5gl2E9oQz
uY/FV//JlJ5ZQvNV35XVGfwYvec9QI9EJj0HORRpPxGSk1ebytwAjJ1dVFceDfpUFsQtVZpBt2o7
ZLV+8zoJW/FrFGnhl3wFU3gqXhLtpeazZo4CPWzt6k7OKal93nUD5buQACUKVBNf4c3cy+h8KVkJ
J/OT+o6h4VuwIfg3JdgEVwD2FTW6GYN4OkXBrL3j8S8jqroIAys+KlfC5yHmpE6zsJFpiriWGkp4
SMfrgxcpizWlCEdpDPaxR5IFZy53Jd+0FPg+Af8FYmcJ1wBww+RdPRlq+WSaKGV0XX1m4FNhJagc
v1xVWYHts1Au8u1NFpt4l2Ck5pnvSfgkpaEXNGa6GsKHaFpAT+9iOcw0ldeKIX+yVL9nLKa5y4Q1
rhLYiIaghCvFqtEiUMgYcpzYKBtv/NVFa0J5q1QI733bYwukPaHFYNMu1dDm/emMN7Y3AZXpCZ+K
vxRPv83mSmguZWPiHT7YN/hZP0SLQd73xBD8bzTj7wipj/gn7X3UBZAY7nSeGIYmQwyNzVa9kRko
Lc+t6aqRpCaOon4kx/o1FlB6sip0fn5n4HM884lDhnZskp4pXJNo+ECTSjtoiNaT0ZXcM2VGV0TL
M+pL55cqIGhSsR0p9fWwzZbmHE1vZA4SNNXqkxOpqiGZzYe7PUoH1h1FaYuZAr81YazViscGgD5e
PPnu86KM3UtZnSC5AEEL8Ik/1OPTchYAjCK4wC95jtGCfo7wJhya0P6xSNFkeq8wXdbPn8MXI6FE
sCsmc8+h/PguRMK/NB6UcddKZ5MhyOLOYBjRetwN6Zs7E4D2GTKsA+fRyRXx7Ln+rbWK68nmYh9S
UpM+UI6NDj2XahruX3hOlmzNosBJtStbb8uaxtek1hOPNi8iD5W4JPdsV8yp0b2BF24/Qh+S7kVV
StIVuu2uUaACiSchPg32U/RBjTu1SuYvMozGa19Yndrgi2KvPh5V8vyX4f+7zxZrRi/KkgWI4hPX
sFPvQwK5/D/aYKs04j2yMMAmSHRAZf9VIfTfaWyxEoSQwbLh5hFk6S4ZedTL7/mQQPQkcf0QRUPd
EsdF9/jSt+cXGtQa9POdial4R9rW4AN0cOX4AVo4gFc5wCTdNfe/zZ9bWuCxExYKR4oKSvQ8/I/m
GKUXQ85H5JveOshHjoVpeJoDzX4X+iYo4yy257t2n2XDfXQv96xBAYu1MgPUGg6xi1F/m4bVlzZG
2gJ12+OwGAOpv87FkGWA9eBEKAs7fv/wAjGQjtfGtNblxQMHse8aNQuPvlr6UD8uVapSVr8lWk68
HvovosA/h1MK3+ZpzdxMEw5jdpCD0bT/ewA3+3n3PdurA7+LX+4HeJ1igGNUPGG+8gpcc8IJBc63
DIRoIV8MVUE02e43P7FNvbq8vt/1A74M4gObXIdhKj+F9tYIBwRstk+0rb8HhKan/cFxiL3mXSrm
U8hRT4X8+XMX4fYT36riIvp6cKQMtJsDlwJOa0Z51aMmoBemKoBvPl440iYfzMLoVDUPWsAoWTpg
jVV10XL3FWok0d83tTP5cGBiznBc8n7l7Fx3kkp4WcSi+gFKT28CRu1sBRsQUdJL8VD2wGfuzTiX
HQ/hWnd/Q1u7iLlnRibElmViYe3Ji55m4S/LtmAc/Jqy3odY5B1qz37XwmV10off1/7qxRQDtBx2
G1XQ3hpzbHL+ASbxTrqg655h1Ya871+ulu324WZxgHWzPrDou9gYUEzG9AiXoMIGCaCQAcXH4O5A
napeRrbAeZkdx4TCtQfnnwFt4uryVV3RoQy+jz76sVWCWK5uYSx+xONRyTMyQC8m2RdtruESmuCj
w93ldNFIO+nHpVQBdaeaIZ/B4myPFRlcqZqtbxzIMhg2Xtn9aelughthS8XNn4C+J06hHOkJ7lLZ
4qPlbr7lhXCnDIoq0Ixop9JRhmrhtA2WW4wm+/wv1DyGW3wpV9c+HKjcEwavTdDQnsVeByaIpaKw
VkKlsRfPqubueSkHv+1/WZaVWkJXb9qq2FZx2qYsYfHSBsthBkxp4sydNknuN3aZ6ihRO3wzshpe
44XgQlCMlfrPL85pgJmqEC9fDvtzoG+IcnPZH13kXs87N/a0W9/HwI8pA1RpYWtvgpHg1fMyzekP
AbLSgmjlh8rSWVTdAfgVfuA7NNaCjUIxt0BShEoGS9hIznPh36q1urRjuc1xXhPY4ogvmR0T9DkQ
mu4xwRWHatjIqSLKDpKfqfpHO8dgYYY0jQqKhbKzjs0SElJwunYhK0QovVq5oJ7KsnqI2pMXd8dt
H9xRVpoL0MzddbGyo5cYgmGVIDmqOs9DUrdCUSJEHmDDIQJATOB7GpneXlcM21eJoj7XY2lD9MsP
OqxCj9kxqJ9gMhD92vefVrlOXMRD/VidVRnb6j8I01kx89ovK+klwGg1cfxhJRh7rh1tq3nVU7ZN
nF8Jgp5gzONpHXTHdJ97BGECPCetgBXRkbkEUx1efD8Lmo1gAfHs6/hhcN3y9gTIbDaD5xApWU1F
2stUIs/yIH6+5/9WHXfFLAfKBEKymFtDUhPh8uTeEG1Eb1xtBvJqFHzS9fxXMhPGpe1Gje2xU9Y5
RU9+EK3oFzuHpocTgKzz1+jIMDR87H/ifvp3uj7xFUpTGT0JvuYykygM6vsrLZ5mDYa1CPfFEvgL
D89vSuRwf7kwgE28qDvLV1CS+qkI+MwYHEt9TjCXVsJQRYJVs7A2x3IS32R0rZJBSFnR/lJv4VVR
v4DFzDKQH94GOyI+D7EsmIbB7M7C20sp1J0jxICYqIUFEhmVyF0F84EA5nfRiL5Ituupec3KhCPh
3ndZb0AMZQy24QmMRKxEW0YIlMqKJwqlf6l3L1GGcYoJnTOL3GY9cCBhlzJHECKbIIiLZC7pHI8b
rQ5Hmo/tluAsGdadrBUw6Du+BlShXlUVt2FT1qBSj3/V0ZZ5J45s5UyrH75vPDu7N1OXugIfCo8g
GKiJHK0mABnL9frD98qR+IQJ+fFTJJg6JOXIY/KN6wRzSmjXR4gXrjoih5t+iZ7Adt9IvvEbE5+E
0fP5RHDNLbF7xTrcY7muXpuM2+SxInZbJlayvpx5ZJE2AJ3ED9tIxU/5zKk7Lqh9B/ikvXrI8SFy
Hzor6KXZgm5xjf5a2KleUWuGg2Gp4Lo/YsEgoykPzPvhivstFer75nKFPRcmPlD1Kfe9iLn/g+Ao
dXtFO8TeOTU4N32eSRi9AdOkoaVvXGDl0E3C6ffRfVrfOLjyLbL6TEBJEfCpfGx044BNCyt0/NdR
2aUkuAb+fCaZ620b7a6kWkor5GjUpVByDcNun+jBG8/rCaooh2yu/kLSF0T3BUKvJKGnhLHGMwK5
ab2y5yV9J5uruHLy17/pJjr/ZIymT0nSEvsLF6/JZf6zL9B44FNkhIE8k06r9CMSWLLt8tFRk8KR
agWb+m960njkBX4z88a4WtdBu0WJ+l7CFpFGlefbZPBih9QM4auYm5nWHN+zNS6h82c/kQoK1Bl5
rP8XtP+QXACtR0SlgfVmzNeCmLuiJXtpzwbkcFXoxraGKlEXaLj2tz3tG9bxOHxl8nlsQ1nXUKUn
AXIamTF1l7KB3+Glqg8vW/84v7W4WhS+F5HPdO5jvy7NhpqRCA0lLbI5lD/HpVoL11lFI9aD1hJF
jJyuWHoVJw+TkB3QW2isC8r9v6pSTUu1YurUu9PwYaA8TEe6qRyVyCXJC1AWyWHkzekq2Ec/ZW4w
XhW0OVTH4Q3rxgX7mkc+v2pniAJ9gdl/950MOxMEBbrbnHIUVBos07bV0fp3450qvwPzgZiaXqov
aMmxK8G3/wfsjOSDyLVUhJK4HQ3VV7PB93Fd+FnzD2CVUCIaIgQHp+Ww5kJhwsv31VYlssU/i1j6
bdNt+6x22EZIdc3HXKNGMnq1si4kKgysABe9OK1GhJJ7Jr42gD8WVp5dFwIBBXaBX1nADNptTP78
+iL0zAWgvWb/bFOY/I6acM4lgoGZG6xarCPANxi1i6yC9clllLij1wlg0IBPEi7gV27ZQ0Hu6J+z
9qeZgQJrJlI/zcl1/w41V7CYr8VhlEPLQo71Zz4G/2uqGF0EBwFSmUxGkaJnl37S2O1+0GAN0+9K
8l5CTKHhMgFyGRlgy/otALfYFVX7PfYwOV+vLvFUhYiU0DiFTFq4wrOAPiocgAxxCVRGZL623nSh
oAJeTAB2DABjTmRPxZ7queQy4A8F/mDcEQDo0ZSkeEZAN03zjOM1v9nJNW8xBMjgCqpedYmQUlOc
LSSjXmgc3V3ykdsxjOQk/cfXnsNhg1tHrVcQdupkdhpsv6YayaluHDaZBcwTUJbzMDXdG8eruoZc
v4PlVp07/hJZSYr9hmHiMrqv/NryHkBz1zLyfnQKCfZ1tbBpGn1c54lcYDV7ZhgvA6FflcUrKUQ6
lOVdjOCnTy/z68A44GW3rNQoMlpBPrlRMDd2NtYbHterHlWO+CR7lgxh9/fbXf/HGUuFxeDDDXNW
oGBsgG7EetoBibb7+MCbylGdmwjJjubLWdM+EoTzriClWvbUpG949cQ0oKcJj8ezjQot3qhqvyhR
VZFbqILSZz8puqSYOe6mR2hTI+kU74xQol2p0ZfQHLbmaEhqnUrq11f6v9NkuxOBUdaFHYAPNywU
3hS4hELRfG1AIMKb3MjFZaSud6SPTM7xJ5XCpCZ1PUoHQGriUNM9xKTGUEo3QYKiOiKfB6NcomET
zK49CFjng3KaO6F+bf6tNQtsjO4+/FESbeB2jfzukFVzNOD41ekcoFO26m/YS+ZJI1ZtGTBRiH7s
v+Rf7x7Z/YJuFTkSzuF3+fd/91ToZlegk/8XpvVBcPh0FYtJvJRvc08tC248BKf9hosDoKYDPPRB
M2CLPRs1H3suYOrkePXKwlcBXw4Yok9MZO3CqRE+0dFTVc4OVLWhhDpVKLmXdGQNuFZAb3EgvP8o
XTeXd0Bd/jUsXUmhrTmdD2uzqVCxW+Z88prbEyqwGe4BOwqQI8aYiN2DO0ktosyynPH/hMjJdz7z
/NeWXF7q+4y3vtPPLp7Or9B/yTvaLdQFOUJXXOR3Z0oWNhQmUKu+3/1wdHgkbBC8sLWG3ekKhDO9
vi5ZntbCB4NAahH+naj8j3Rvu48DTTv5SHklo19BP1pZpwqxJc8ZiPit4bpdoPwS7lfXdfhe31Nf
k2LxHVfPbjg18WJsr7FGBibDscRj/36AF3jkElLjaRs7L/TtLMyupEaxP3ApiSSXindSc2Ai7IKI
RJQpoDFW72MRB4Fr85N3+cBOX96BnInO6I5kVSgUODZqchQn0PK8+JTiJSDbL1W2A++HyChapM3g
MQd8JYGFJ+4hZIAsc7jWeYj1UzczBipya2h6LKSZLlj4omT+EAtVAUdBPYAzZpYgkXbBygY/2wHu
tX7Zqx3/UXNt1VLocfcnvxBYc7XgQqf8/iCKicRj+InJUy4NpW853Ft/cX7suFpnbYivZ/+Y/dBX
L8EwRGTcUkPo8mQIWq0lNrWmHh6MzmTkYUQJs34Ol4wX1xzvgjxkcoC0QMBRk0Sp5eSnuYGSSMoT
Ux9ZZ9xtBbzQd/Yyka7eLepSVMg1yOC6Zd/hQv/oOfDu5qdIQaAe1A4XIDVXky6skTEVySHeig5d
QPStXMEvWadrhfyhyXAcHW9EQwu8clnbRT08g+3y3jMQRVunR7nM9f8ykptXmtEslrKM0MwiL/nS
wKRb4tBnA6Cw9qZJHB9BlAi2Uw1tG6lEDuJJWhPAH9UQxGxn0YyoU4mJ4Stp6bIBpXYUiOZE5ucw
VuZTAzoPA98s4J+XRPnFYjy9GmhGGsm//lj51yHkpd5roKYLx46jT7e1fmJuU16vdMxEPRRft00K
wund6ErhVR9WCiY1MbkEVyIH0bpEHOJJrn7EBHC1WYT/Cw1LoP0/5quT8bESxWi6sSEMBwvyRR8P
OL+wVQ58USENqteAIfhax+/XVuF9nHiUzRRfhHbi/2p1uNB9nGQ+vorjIFjugGLnVCBZUQBJ6c57
0s+ddqQcavIQkugfEugwsSe9+3MaKyOljQo00Pj3yYf58CHsOgqyvprd7ys5rBOL1UIcWwVqTTUK
z0rzXo3JTZmwwFXI+x3OWaUyzfUAu7aWjqnmQyOTXQaSbnFlxAVaMbrrt85+6i6n0mnUcbHtaR2F
6YdC+Foa26NHOpYy11cSzAAASzceb+HCdB9nS4t47CtusgBQh3SCxlrz5ALLB3BFW4sgPquG+t+O
um6FX8ksi3virK8i+6AMbc83N5sZ1wxlO4WVAQY08YcxTTSFfHuOh96TAMBnYSYCG3BIc6IUNBPF
nSvYQP3hF0wbM4Nq+dX1apomVcgswQeGlnxC61oJ3QoHUEnJ6IEV9OkS+RyJ71UKGE0KMCATi3uW
xor+PEK0KlBDKNjqnK/KJ06ZheVRI/7YlH4prDoM++iyP8iekslQW46dUVQkWMl2tr5VJRXEBKzE
nXtrIXB6fahQ6WReFObAUHl90X1RDBIwwuJqNu7SKiUi2SBecJNvJzti8zcjh9+HGl6FBTw7OxCF
g6msNxYJ7Fv5Nstpc3jLOgL+1ZWv/eBNpzWCiemFInfsjaFuEq1dwRe4P4elpjMSglIVaKobumhg
pa6jzloEa4SMrRtIckfYG/Js/TrjEMRAhadq9Qu7JL4jehpC+VHaTBOw8aI7hNc4oUrx4yUJCAif
47H6J4fCgerhi1XojDmQmg01BmXRCt9TUUswLrtJuCzNan0ebYo/Ays2HxFoi1FTT4w32mLm7MeR
tdK5tfXWEt6iLRV4pOBPD1qhLyxHNWrzbgK/DC+vvMiWtCMVgJZkREErxekbbGSjcSEtjHNHedYj
cIlcfnz7iMm3oWu6oUdUlvVBpPxLimP7HdyRiBQMJn/mQZexj8XCa3N6ztuKdYuXt/pEFgv5+Q6t
oJsvE2l2k302WB0t+6msrpeoRJsjpqy6NzLipAc4QOpFHV43s+Y5hlJlVD+W1Vt4+t8Zz2GompFR
ztj4082hZNJESKq3t2cTXjKBqopLmfSxj8G+RlFmTPiSAUjDNg/MqHJzUrVIYbzYQDzpTJcskYwK
1sVBzYFMRWEQdgwoxPvfCclX9nFv9zlwXJOKQ+oFS+i6aZz5HM/cHVgvi1HuGk7pj8ic79qLo3cc
NhFDsP+2Zi9zO91IJld9ooKkUhoYANc692p3bRXuR3dKSuYADS5FXfP1IC2WxV0w0tEnmbqQFhVg
SLdnOgwP8zLa6vVYrztXhcOxq8ozJ3MgeJvDgyEpYL2CRlZ3PzHEyGXAiFhfzWs91aZrrjZlIW7s
dZyyULgErJ13V/6YCh3Bar3b2W0h4TVi4K8rNph0yDhUkRMhtyY/TuFRzCA36H8uRGToeGD+HBLu
vhZ3dl8qKrtHcoGnPIH3hguhmQ90AOuN+Z/5To++9U4IodjRnpnvbiifl54rxpkDqxpmMAHgQHfO
NGInTC7AtDV9c9pj3GltvJ8ysNIled8WofRVJHxOTUhV7ljyq8+FFbuo5Z/kUi3ta2SBz11JtDGW
qh7E8HLASx0O0G0eRPHl/9TATARv2K1g3LNrQNKtiPOqGTEp1siwRTFJCLQ3um0ps3I0P9wNGOaB
x4jRWU6dpbgb8tVEogsbivjKw6vCcsKOwsMxX5a/bjHyJjV4s+NhNPcGVzXl8VUm3GwmSYoE/XMv
AloKfLdQ/Eq7/KhowNdWyqkJttzG03vwBzLKqXpFOQGu1wu5r4kc5qOMt9WDXUtiG83apEhFs09F
k06Gh7NkoPY3wHmvtsV5awpA/FojfF9Ws7vJva4JMrftTnQq3KVtJSQM0LMg4O0NpFKM11Jcggvg
ZZek5tC6QsVT+W3TYcbv9dL0olu43/ap3lW9phLq0PJSpk2R2SBvL1Re/KD9wYkw7oQQlJEBHMZh
PoeQpp6MnrOiE6FHeMT1CLAeVjt4OiGNxQ4r/YVFGj8ylB9vDS9w59eSLP81NPLPhP87nwKWrOcV
yyAotQOZAgG4Jh85QOjcuV9LX7BTaNaMG6sCy9KXO6v3cRLzhZ3lR8M5vIwSl2Q52idWkoRugOPV
I06kWuM743O8AZbquPOXhy6P/EUgxbLD0FZqgbYpXb4sHzbZl6Wo2l4YCnPs5tXhcTlBV37gpNBb
/0nLURFvnutku9PZXkkGLeyGTHAkyFC4fvlRcjkhNH5r2yNdwiC7jCboR0A+djdo/QNzjcV5vy47
7qkGxhIIzTxL8hGrJzbjRNEBbdNdkoBDN7P3eDpiGXNl9es1krzQmP17qKgpxKhfzBwZL9qPA4Dq
5olJlItUcun7A+6qrYS5dg+rNVcxbFNNfyrO6C80f1Qkf+wAxRCZxMzRDQFHKjvk5PDJc5PdHnKL
wV1Rkgfo/KrJ4OSa9Bt/T0a+Tf8AxI9KOqgXIQaGWZo6Kt9jTOUbByPzZJok1+STT59twt9lngB9
8ZbQvIXZkc64thA51YEh/Q+iHBBlNeFVlKNpw13eg1FyDNDLBYEOIkL1R3nEv0OIxx9fU9JC5ERd
AGnnN4PKp6i0f4IzxHZvxmEBEB1t2OvrG4/O6La2Mk3ECN8hsuUoXJczgK0P6d4ORRnsouaJeq49
da8a0w7B5JStIyKaodqWhi/4T2DxE+z6S0+wSkCfiK8+M+uPqTAD9zRfGkrYbRRIphU9zjorJEjK
96cHfZ5xDalxx2UuICoYNjGH9lipsNzaZVANdMBi318uxrAE7fyfYUNJ+m0P8XKRBcirgunP2+LX
O0HqGxELcde7fqpemR+41JZuwKccjtbKSPfzyQgwE1jlDWNXGDUssDlQ3XFTnt7PMCM6aM1e9UV5
WqI/fXEVRN5wqV/iHy36T4wPnDsc6c4hOl8NY7BS8mawc2LnRp6a3b9YazLLkJcnoAWUlFRyOXbL
zDUoe3Sdt6CHx6pc1pWBYeW19IKE2jwzivVZcKooDJ5i27SOA+mRpeoEWOigsq3Y70xnQgjp9cbl
iOUdXkgpenl/p2q/6Dhox+HF8nM5/Grw2liybdkpyeFCouKhWj7ilACIAFC7DinJhg6o1wvWXx+7
ss1zP/hZ7OdEy42dMz0FobgStxzdXjhdFEGg9W/fYxoOitylmXwjS9zViS1ehdej6tFJNI9e6csG
HEw92K/d3bPRB4+cGr2kOIek+DuQlur0VvscDc/33/gibgjEHp7aAjTc+D2TYOl2Q3qXHyAFgWyM
U0Z9O1RE9HrUJ842wGAwiIrJoJYjyPBA+6aqbII8VHlHNMFNwlcCkZT3J4qTDLdZWKLjKf8UQfkT
bhHs1c5JhG+5RopGa+PUqeRbFqNV47EMO0+4aThwKiV5rdWnRiOyT4j6fSSVGE43EQfMLbmrpry8
tkJQGAvx+ZdlJz7J06Rb1Zt/G2AoBW+eKXWUYBntcbOnOXKL2RkgNOc4WaYJZMTFYpRqO1yCAxR7
VFAvGsU0bE6ZhPBSEY7hePAiAE5mMgrGIlAwW5viPtKQmytYhVChqxoi58EuXb9KiEDCjkVah7Nq
XJTBVYFafV3pmcMPhQE6krWCbveXH49fShdCUure6PW+6lCPUDC3AG3/YTiaZU2DVvDRoFahRckW
mwXTN617QDJfsV4XHI8CKRh0wJH550NcQKoBTknZIBfYcEXeE5ScxK0rwQ4Ky1sSdW4AOsRWUfjT
QGlQXhXGoo69aacjk+ICO+aQsBaIke+a30qXHL78YoVucMAJJ0n/XvvaBdwjFxXsrbG3mGmg16MM
zDQ5X7n9tYywvQxQvBKNyhtZgyh/GaSB42bR45BPqpdMsA8SCOIapmrtqSZqgnUkfwEb7+yYHq41
Ghy9lGqvJwqnYR8gAZ8d5z+L6oypf/N+p73lSgXbgStH+u51OhcuQzMG5yUfLEKyWThNyEWfRzIa
58vFCCEPyE2Xy26+ElyopynHfkwHKDDq79srr1HtSEz6Z2V1AZNpWBw4y5rsqAQ5m53+lzGw+4r8
ZCMaYgp1Zzyk6/nU4xWb1wTVXO+f3rbem7aZ6eiTaHjAb04nLD2BaXI6iQaddOz4y39ycmkLvAz/
XKfmdcMZicVz9KK0ZMBjLcRKbLjgPoJXUj/3p9asblXlDKTsg8lGI5BpV7sN6EEbu8fCqaWvmI9V
0iGw4T5+BxBNRITGNGfUyu5IEZYR58cB6Ce0tyYuGHVij34OKh2Q/7cmV7oN8NFF+pEeH1s2Nu5+
8YXqWghjMLaxF2gS3zlAVqwn5keAVIyhrZvNnO6rDUaTiMw62HBeqq5e0vJhDvq8QH29aOGreKOr
+73g7TmP2LhxXeXe2Vl4Ob8kTagViJda03xKaSu60XdbumAlwaB04lXI2Iwa20HRpuwJ5JmuGqsy
/FpeBXu9GBqT6Y16U8IM3XDp1Xg50+OhkfazBXJS81RPmRPQVnIrpesbHUp6jBkVa1qk2s8LiZ3b
I14MKMHskmMmdxRVIlwT1Yr2V+krWgqotzy23LxqOXG81A+yrSwUyglq4V6a0qsgkxM+v7RNC2EY
J7Hw4vs1hPf8f8DpxGH30eoxh7OkA0FDfNshrkhNc92JGQO0oZJYmlLRZhXws+mPVj7ApMrp8OH/
s9N9DR/As46eERk+zTEMnYt/gnbhAScv4r6iiqHV1p3OuExL5vK+VZA5GVIYe6b9ZxbQxgYT3PxK
u+t3aDIO46HtckzTeV9bt/oPO+U4maoEZhZPTNkr3YZ1L46O42HW4FEe+kicb70bGLUKbGjjVW+U
LS41L4qGyGTvgPi8zRq8BRv5Qa6t+VfnS/hOExDXDe4j32NpRpbMAN3KGaMFMeSJBEziaMM92b20
Qz0lvmv0tXW3H/GCuCUWgoSzF61yJgq0BIFzhckFURy5HAOH1CDQemlFahgo2L3ZEfPS3qANGM/J
LOpuMT9D3WtxYsQjBIOzyGwwF4tatnso+wwcthEko3LRCyie0Mb48DgcG+aKqHoikeTpUQY27qho
gl0Fxw+NWBHSPtiehmrmzQmcmQjbl9faVV4irC9z/nvTV99JAr7GCvVG2qR546i/9G345mppKQmx
ui8nC1s/3dZzYgooE6Netr7PxYeR2+cyYqE2KRgnhxgONfDBt0/Eo1dh1RGMBvKNIU4EmAAW5/zG
dvjfYIeDG+TbWyzoQ3+FVCo5lktQeshz7OxD6IvfjjT1yH1qQXunuaJm9014SnFERDKHSwpJxQqX
UjjfngvuFH6bo/Z5GUbKuoAIWWtD0o9iy7g7YgjWi47P7WQcB3IYsNF+EeLZmFifehSCGy7P69bL
74BYRkxxNsoNZLSGTQDgAM/9wkfWgELiXSg4Zzi0vNlAqlWbmYBawuJqAuN4TfU2AysTzg1w4e61
ooM4+b8vsfndnYUVPCoZro2i4K21qoJjzjsGw20/xiVeeSG+DkmBCqo6S+9tA4ACN96euN8/JkDy
dad3e44c1/miv8rfvnZpZtU2/hCxXg6oYlKlrq2yZBibYgAflkl3h8noLKzGKyozhg0uZzMU6wuB
Lfp6J5vkjMQer6hqoFIfaduHd8dYe9fgfVCkaNDmdlkjNC2qT4gFrhkXwhkHuUqXtSUpP6fhIc/z
U97vEqJt9zR63ia70Admy+DFjvsdjUl8etEcINcKwAXRZBuJTkrq6n46a9AR6iDV5H8Nh+isP3P7
7Pz3PipBx/gwVQ2ZC4xIDQknCa8c0udIxRJgiWXAYAMyXa9S5dXwsEDeXZA341s3FgZIMt35hv37
hFiP4mu95YLoe8TZmclceUMObn6k1QCASouObJGVI3cLQmw6q6BZs0JJn1BnYR8u5oHg4ACMLEcX
5a3c+sEfq18dtrCeF420jsW4HzCuKA8zVleTAcg9+s7OdCif+M36EZiTk+H7EyLv05U7nCNGJ1tV
BaKPxa+zYfMLulBsADlfq/re6362LKcLn2NQxE10ofMVpveHmiHYuvpcrACOBYrvj7A0NTFz21AK
8++DVdjm9QjzwTuwfgmfPZtndmiuJnVHKEmCWeiN4Y8oaNtcq7bKceLecSPXkQa0a+JgbWWL6iYA
QDNc/5Uy3fMreYb+b5DYYjUo3tXr6nfy0/hPbTp2sLB4BZSuUi2UI7IHzrBVYlknaIBEpbBvtSVk
NuXPa1fs135LIWSV2lvu0UROkJp1PT1i7jvFFpuIot1lzyaHyJardtvz0GrqTR/xuURIjDi0f2Q/
jkMplCuYchoIFIMJkidt6nvrU1ebe6IaEKKXJMQO2ZYVxghyeTdGlo642o2d2GWQF8418p/fkZhR
9Wajd9+6t9bVJLSIrHSwpQVcoR0b016MUPx6nD1SYfHtB+y7HrM+4pXFl74ZgeoAGKuNo5wu5pe/
UXevnnj3fRPYZxawtyJ3O38hbyYPjlBk5TPNm+3Fzt4NzLmL51zP8rc8UE7QXf/tTweA/2iZzyEz
d99ZU5zmIF33KRB97FB0xTtPuGsiJ2S1SOF4VbDNP/9CrQsfsZAHt5k9caUpZKOwgfjQVAMNd5qR
it4kNM9OzXedp5LZWmcXXe2+Hp44xKMVpzhdbsYEePLg2iA1K+1H9gUjeYeNujdbwJFn6rftAwNR
IbRWxMbFmFVou9V698peLUlmckyQcajW82OLVhJc3/wz2T8CDo5+H0MFss92eL9VTPGPJaiNjkxt
tY0QwMPsPO/iBG7fTcsYjqbVpTaDKnluKJOKNtBij2jFtYkEqvDcUgzkn//mZLSarwqRy0QsQC+m
RPAgH/JN519s/4vnUldG6BaD/Q5wyVo0/SedAaKgN7np9RKJRQZSxI24//WkKbwR89F8NAUUNR6V
AHEkOkmOTTXIlKhKOXCiaEEsMaegKB+DLFd7V/NWmrq59aiYPQyT6h5GlzI/4J+wucFeaHvnRmFz
Azj7Ce//efEmzOIt60WbcyfRmx1opKUV05BXG7bZ5dvGz2/3FWsqaCsWOps/TjW8uSMpiC9CplsB
Di32RloorvgKTJs7aybgyo9b69eMo38XmYtGH414q2gJRdLjwFgvnqAOsBAKwkCi+ApoqQditY8a
wiCeDszQ4jlSrmQXu87yT4rgMhFsygGHEEcXh6XwgURo9yNkQUxrjnct/A1TBFqLpjzXvIIa5wtY
aMlt+utGUV/6ud1IxgSBXOsAM1s2tjJ5QaoPSABRM6SrHxK1H+VcrkF2k33ZltOxj1ZhvKVLAg+Q
0/arX2ccDwdn92tOIVv5y7pdTeyEW0lGYFxjm5fh5GNPAOrbVCXpgK7li9IGAr6ENY4XwNsq7+eQ
bCiXuckncR6yPfUyFd0IjLyOjYLZ1I3Sl6WcgAkAS1niaBc9Tg8ICyCFfmxPKdVcf7Rqbj6g/+Ff
c/GhxN5CRJcSTm7i8ppGukIFa//zeWBiIlfmUmz2Q1zEkQyJX9xoj9V8w/s+2rAVgcYsFtTG5S7g
kEMKQgZYTl2LgIz6mfYc+qtTzh6WiTUmQSpiu9h4ar/y7N3ubY9pJgo40mRXw9Zo/gSF04DbRuxR
77j3YoQogaqfouHr6Je/sEzQjAM+z6Kxfe6SHNkNp48zOZZ/31g19pOP0WumSy6gtj4zsI5vbiMr
XkUDs1ZqbZIyFOnLYSDrBjFf2oq6o6LB2oOuuZOYvgIpubToYVicvcqgdsdUeYGb5G8k8RArzZBq
QfjpgRoHK46mzO0Zi/VnNR3dGkyOguxwV37dfyoXbrSfvXWmixLAJn+Kvw6zlgGmLrSgxjJKLGrA
9QwyTK/t6M7g2L+x7sqKCie47xboDd/Zz6p5kYts5BB6xw+KGWxxQM7zUCWkEqRZj1bkk6oRv1ax
W7lcaaaEzM+AM/kNfoz9PtQ91yFvqrA/Kue6rRrBXu5OquDnyS/TKjZGYb1zyAc7esS32Ab1wtBD
f7qV2c4gTcwlFfkAVEwBPuovOlTxK1pp5hwyM1bfdkNC/LBwTjlu2FRnx6Ci3gCpxEQuPM4XJho9
ncRzOeEGCw9tbTs4WeL7bxDPw3JkBA6ogv8i2HZyewXKMkzXoAS8XqACdoxfIMHpmyN5gKcX9sV9
+24Dw/XhDzrolKW2b05icvjVy0O236q/B8vUQG3M8nwjECSi0DSv5biVohWlo1Wv9rPGgDhWQS6p
K/doNbgQQJ5IDEoCV060eAhAHC/41nqcdHSC5wvWX9/d1mK2sMtKOMaP5Hi+oQsEX0G2tCjyGI96
OF9WBm8IE908m6NCS+avmPNOWA0JX4FAZuJMSygKJ1FZIp2PLNWMuQO5XV51Up22EImaUWSBgbN+
LVJZa8+Q1cdsdT5FnwGHDBg5zU8y+DSoiw8DNVOf3J7FhTQElt6soCWT/md/QxPnilVEN5eVs02r
0/ozNo6rf5/gBh2JKT4gytlPdwF5Dw2XiqjDdVYF0Vh34xl1zrO2G/A9k64vRitxd/RVv6y3wlWl
MmIjNB3Nj/F2lgGB3yz72m0kTr0f+yPz6WqPjn2FVMV+nLe64KnEWwMN3u7d2Kwv6lzGpN91/DOt
4IOQKdoEnCp66tiLsJTrMXL4Ee5N14vARdKJr4M97ZDpLxwuOaRU8kd4kM84rqTb5UjZSWIDlKPx
0AwFSltXiSowIa0hpWKnscgcSBcK2keImMbi56jlvje95dbClf3bLxqQaQNByQx+LcuWTetnDg13
W76NZgZy1gfOS9TQZOQd1o2HapJJ46K46deFFtRq0XfkE1pGGCpsYRGHi0sk3eZRlHgP/4Y4wCbv
B3IRvuFcYkqL8YR89t2ps5gTTx8I6zOYtPxeSU1w33m1jAlpfg1F0ajWMvLhnUomh8a+Rq7N1VgD
gZVfzgGaj/dJcPoVWRqY2oCzXcVQIqIQ7X/bzKw5idohZtV7KvAQbBQlQZh8P2tMJx+jOOKWPre2
p5Py4WV0z8G+LE7FtWQNWL5gQ+A0Jf0/KXEwah9YqjrQF/vXtXT//BfTgyltdAAwzm/NwluI2+9t
zzM+6Qzzpqmyd/0c0CpKUOBZrz8wWzd/VUAXiHy6NEOAIE0Kyf5ICvpCzO7MXoNZ38rLRogEsOLQ
R/mJNCTXCCdE4PYYRb81/aqIyuJU6eUoYlQi36PcrFereDT6TV79VzyW4qaTf9GKI/J678fOnCgp
vUYS28T13vgXh6etFBM4YKriGojF/HzMwcosOPP2pYQiFZ29izMdX6Bc0b+sFEbK9p9YTKbX3fLV
o+DoJBXOtWgOffUtxrkXWj0FPF0VMGd4/bp2WEiaTKAFX2+0/mGxXT9WC21mMUojwxYdXlv+xpRo
eomtEx4zdMGWXcHSvyOavM683rG2Fo/SpBg5ESWT5KPAZanB3nBAUh4XyIT+n/fYp0N2f6to81cj
BiyrxR1F7/BoYPhV/cjR8ddhoI1T0ReAeUFWumiM8N72s1Tla6Z4IEgrzBLZfjRxoqsUdAJivsmw
DsiKjitC9ay0PCwwbujl3Lecdn0bSXGoMiW4C1VVRtc0vA6KzyYD1ic5JnoKIPmhSExoWc9LupX1
Wrxg36NHlFnMkimeEwq6I/3McSKwYnkwYqvN5X+pFXK4do5405bBlSiUtD9d5oN7uJnSbK7bmoa0
8VQ9aJb2/f50tChQTSzsUj50/wLVXTWVx1ZfGktDwUOWnR+8mgTlgWFIEfl+daE3hLn96N5IhuNl
jY5+rJFPrG94AOK3bWrA+ZpFoySVkJoRzgN+/HuvPo/aC42PjMFCBWqwNFPBK04madS2OFkojfXK
CkceIsko/TSRwrbk/K14jMlkg3h8NE5u3TE5lgS70VqoMtv9uKpzNnfqp5wkFkyUvlpma9xvyxYm
XLcRnUKs0Cr3CN+4njRviPnGfyDIvl1t1K16WUdIXHy1bHB/xn5OensKNoQ7YeAvnSjD7+2duLAL
6m1x214k8RUkK29GHAd2N0vCqa3PGdy0EaaXJFROY6Rel00kRpBQXHlJmw01YGnfKop5ldJ4Fi1X
q1Ddp6emAGRAQl34F2OjDUuDgRhnF9PnDyE+2kgDXMlnRuTb7d2X6/sdaHX5WagXJoW8IVDExTNn
mhDlt2T5lVOj9KqooMf4X5Hb0YSZ8rWnltdQB7QfgnL1tmBnGNEP602Iwe45H0e3zKC+NBDYT8kz
bZfBBtZk3Q/Cu/JJG0360REIs0ESiC/qB9+92oLBRLE6lBhnUQnVNPxiV530uJNzJTnZWZRirRtv
OUN+XnqvPauqKwbc9NL/2OzLySjweaXJW25GIb89B8zq+XV3Q7xWpemTtkFe/OmggnXdY1WoC3K+
Lk2T4djHpiWxfXcazr9GvQE11viTrItkF6dmalyDv+XRGIjKVGaBKRhnGETwTIAE5/t11iPASXKp
RekB8TJBd0UntuEGwasT/voXj3OdJoUFHQSAWShatdfNZIXObnhzW1sNWc0B/9cj06+14m6FiKSd
+uNT221f+vtuouZcekQH7m00TuNPNq7Pgi3pe4fXc5qxRq9pSIIOEMcg4Ig0yBODtU9+TejA13tn
1MkS93v2TFISUIrANfJiBEKuaac5MUgynBTvJtijdvoehEm/nzgSaCoIhiscDt/9Mpl36eD6geFz
6y3sj3o1VgcgodGPZpD6ITOs0dew1PUo14G/4hJe3RMKmAJhJJt77FMjnR9AQ79X7P6fRJqPNhuz
c9bvDydlm7RjyXIAmbr/I3ZZPtDcKUOjBrv7ielX3AExloIQu833IlHyWgA4NLaJlIUaftWrf8vf
h0ieGpxbl69PeUUjG6XKCiFpQ6cjVF3ySeftUtPEb6vVpesp0U4lty+GD0Taa3BuqNUkQJep/mRP
ggQyyEeKrnRtptDP9py9rqkqeVDbwwJ/aosenXhP+uMjpevv/cRtQBCKK4GBrvTy+zhPyIDxucY/
qJCPsBkLjC7wB44D5U/srurvyvVrZk2cYHcJi1nv1wLQYACSncIzfjYq7oELu3yTA51tlDnh9QxN
FEo5EO5ie3wmJE6PxZAILCZf33lGRLL8Ky55DzfHXcUSO9w3khnYMarQ1M3++MKfySRAtwSk1HKh
kFU4vKoj1Zq3qqrLgGX6LT59WOZMbG+dqHKOuWSIbMkVjhRE3Wfi+dBbrkfy8QrEJo9bXfwtCgmo
cTlkJT0lmQWUCZal2smNh0uZELg4YftpSeNOKp4Kbt0pp4K+ebGqce0z/L1mOVm+eHlB1lalGPGF
rKQf35SY2MnnvaS2f9Fga1eb9mL/Mgdo16hyqmjOcNl4T8e6N7s8X4NupKpr1hWNp+XcbSRzYY64
6qwHSfyrN2j9XvHTueH9Kp7ZwUxcvCUp11OaBWTsQ0+s5TovQx/1+xH5pQ8IAlq8hevUKoenmyEk
tqyY+EvR/THm/i2hh1UPQ1wMKwOkl8QqQiihsmfStqG/srVgB+yzF71pejaVZ9fbtNrx0kPsMVPl
DrvlKjlmJMHg1iqylE2xy/WvQdZA1wLaFllKPTGQ61rl72ERpJgz9H0bDsag5DVn4uj2NcJoUfIo
NnF84va2phBShM0QE0YQ2xNezr4/ABqjORoY1Jnz44iT0yeupHtMo82Fxi8/XHidgYVyTnu8KT6i
zkagITDAqORxWQHN/teLNhB6lrcfoPF8eSn9cymvbs/6PjAJ9tD/OzbCl2w8HjLKx+6aCx20WLtz
9bC8jkASO8DpVj85hTYUr7rPOnqSgSkCSKkHgbSILxk6nzkyiG5yu7BhWjcWdYHJP6GUlYvb8Hk9
y1hWT4GQ08Syau4nWh2nAGnokYWmjYZuKwX269aRIzr7dvBExCwzcphBxIEZSlhFEdEPduA6LXHE
6RIPwIr7JAGRQNXJ2tHDQ+SNnfKlKpWffQWx97gzi6zh+aXHVDZuvduUpGSXnzsnXlmeuIZJXGNq
FWiAQAMU1RoX9jB+Hs+fAfaQituUSVcGO1jy7HErvCAohTcakiZTZYwaX6wVfoeEQ8DIlTI5VAIX
6ETBm88OwreB3SKrAKA/YQUlAIoD1cXmO7YNhDwmZr0xOZ6kl11QvxasHy9w4ygBZTlhsX6gXTGB
/3qUyVPm2QJGQEI21kXSkC+LHBNu6K8WT089LK7ywWU9qK1hPKk80g7C3Ur/IwkNghoXzjnHU/sI
U9a4KTUtUAd1ivYYTiTXGTUetFgJ5Cq3E4+J3jlY5QTnYE6d32IdKaKQmuPPbxP51jCTiA7ksP94
UZW/YFJ794Y9yIaKA7O3V9TbRDvNUPggMAuV0m4Jq98yb7Oh/zw+E+eYh8by2c8bQkkV5oXofhyN
fLHHhGlNRGLaY5VIWgjdVaFZFkV5W6S9NQK5tKO99Ho3IPF2TOpBUGlBU5Zbsu8/voc6x2TCkqSG
NnhNhXTj326+gRYpY63qg/FOc1CuZmwNbPPG8jG6/wjW/HG3u62l327r+yXBU4IfQkHEfAvW+MLa
qU7ncQTvEh+f8fBr0nCDdXYTJe5tO/t+lcU0b9QlXXG0nbhZUhB6P8lUmBbCx17u90HshazNiTWX
+x9iy70Se3kZE9PaoAPhJqKd9egfr22WrH0/5Lm0TpNClCORAM2lslkAVe9wcP9UJTTL5g7Cl7XA
77B68eRpUs9FCL/M9ijJedzLp0NhJ/v+XC/rsfUxgX3HbZ0Tk+AJp90eWQxaTVBIk73gp1vF3SVb
4M5v8YEr/Cw/J4MHDJZBKVOuJsFTUrMq7/zjd5g2gH6gWYzvN3763O6NHSb5Eb4SZrvoabC5GMxS
WdTkARe3vBMYZxeWt5QZvCsBnLYqeAR33MY4euZ6cPIwKQvf0NLmdOVLxrBbcFcREoq6c6JFiwOJ
AoEpGOTLb9QgoJzCyKK29+VGhxae9ag2RS7j/Zvj329ejZROPjL5oGK3CwVgmFmo4VWKa+5kxew9
UZbODMzKR8pY0XYKLL167aP95cijzV3T08mIqb8MisdEl2/NwV6vAJoovrEL4Tq2ojBfS8fdj4nA
ASjQ6iznIxuJn3cGyuRYSVxyUt0ksChlwfEsGzT0npPiXxc9ct26u7B0lA8a2N5mj168VSIMWchv
X569m7HsThe7nmEStrIZWh1YaBhOqIryYnGrxAei/4U3bdQpweMNY4OObkIeOUZuHzWfcAVeR2Bw
eQ6gb+tzaWn9whoXETrjkgVnOuCuinUDjjJYqgjk5WntBcZV/oHQlm0G7fSsv/cpWiJTxlwZ8oS+
qnzSEE7Cnv6JA9IPaU0edZxo7DM1H6mP5Jarxu+hLCB6ZnRUW7yvCDLrcKAtUCn9a2/AwCI4g0bT
ZoB4hPQVvsbgAZo3g+Esrw0pMI3kIINLxbmf2v9ohCY/+5nz4Xab4yZqbiZjqY7wBzmmpGjsG+fJ
QqRly+4lqLXXqZEOciIqq5wt673em571RMqofokgpiMf2VM3qPAln72ONpvc3zS106kEDhn7B0le
jS41u/8EVJIBWow49lbQKLZVdVwm9e6R08SDbbHOguvvAtfrZjFvy/DysNj5fOgv3QuWCCBzhJVM
MrYkoJJfVrY5gA2yWo5t0sV+pbO6Bki8HcSiwaQa2XdHpmUEde4e+imqEz3yWz88tAURDgcFPD4a
wYCPoCFAgmXxvaORGw27S80hYYH82L6dtoANY6FvDV5K921J4OJl+4CtxtN1kvbf9enRYeSwSLkK
P89iGhOWIPiAOCaLmzon/j/1kdwi8/tLc0s6u3y6BupnJpV8p+rbFox95gLi2gidm7Tk3A29ES+O
rgMH8hHu9ty7wBhyxPyOTdnI5vcxRmdii+uoXSU+uzP50CmO6758SkP6bCzLlm3W/ZNv887QtJtP
PuWhBp1UnC4P7HtolA/wAyTOVRZ7R+oCVoY3E9dhpCfIKascdPtgqWfkqVNOMQrLwHGskI1oMNrn
ZoWxy/aI+HjixbiHWG6gPX/w0npiUCiudPsshlN/Lsc4WT5B+vbJ49v8oEq5hsNXHF7rL7GhslXP
tP/8gvP4TgLdmX8t23tshUo8SEq1GPeoc0F6V3TQ1ywn9+D9fuKgQvYT2NKmwVvlDmmOLoSHtNC8
Pd9+30mpRBckaT7c8Nbz3wmZ5t6VfDXDwzMWCXBAfYDi5Yd6+0BN3bzShKpvazpqH8tWz2+j/eiR
RPm1iEueti/c2LkcTvjQgft/yeGIskfPNIVzIWE2wNJ8guHguRAdrKW/O6vA5MXUsl6NItmBn19V
i6mot7DjJeclawI/KzW6p7+jafLSGwV/9WbpgnpA5VCVeAnZ+bekiCu7sqyqwPsoiX1xc+azQzQy
VqEAnkAYXvnzBMk69w3f2+K+z6poXk5DrxXxVQHpB24ptUIPikn4M/kbzsflSnTdSLHo4m81HglU
z3320B9K899LMovhIIXtBrnOLT1AE4b2pDdtKt/Qz3g6o2z9qoQK+1rZdBdZKFktFEluZ30KNGih
BBBN0edu7ynsVLcbrpO++xJiuG7xcdo8lkt7kCg/FAdjeuH4OD4PwpSj5t9VbKF7zGdzq0j87auw
fuXg8vB0AzhVDT5Gb4Uq44DEe5qW+9apHLZwgHh0GaDEp4sTnzuKC62mkQ1+V3EfuWtMG3ShSMna
k7zi18+6CBXOizAes6HPTjxzO/scH1GRkrSIGg0hdkDycKBlu4oADbcSv8ovFosnnnJNSpEGPcox
FdrmrIhnzjO53OblmW9BhWpoqiVQu08lZezKsZUwtYqQpYP+U5LslMoCuLoNAyGb7A/s5tkAEUtE
KMtCRnWn8Pv3zI8BbDbfSXlq4FNF/kffKxLR+uDnvhF0Ix610BlPjFY/KDpaW18mkBYDy2M6JQ4r
bD6bj8O0yng3xqhF98uJWFYMyjf74AFmaOjFaNRl4PbttSiMBKobKg5uuxlnMINLplX5c242Xntk
N5mXattEXPB7YiyyytoPKa1NiXP2kw0NbxRRy2EvYKttbhzy1cLN+B/DW9v7uvd8/Qmbp4Ae6I42
uSQ/OrJcF6juZPMUa1c68NegzFUTWLEkEcISSmGjFfvSy+/5tHL1C6kvKdcXfs4d8IVZSGXkZJHU
kkRMPumqBX8PbzOuPd6qVD59isGEmEINN0QCOePjtBmZ1NU/DmgD1JJuSPkOzk2KiHO6FkBvyw5h
C+7kvupZYx4rGCukKjDi4uctqOUGEOvrm5XUgrELR//VQ+7CQx6QVz/f9K/OOdCD8DGk+ZTWAjBX
wLzVPnK4FML1yQVtKTBf75fLRZOj/XQq+JbwJWIwLAV3aWeBOZ6bOw+gNpJN6H7KsADMb0mJ0zMz
vjVrs23h7gXpybUkQjprrXE9wSj3mNlj2Z44hLQLWiSTJvvGg3XD0/9U8aWKmdeIpfiKIVxHd9Q4
5VKChHPez8yCuWmKRhT9I9KXPA85Cpbiih0I6tz86u1B04A5pQ1f1sqkNGuPyTMjGvTmfO69+8u9
2JJUYioQxdnTkmtBrDURVRctsLeT2dhbHuUAmfE5oyKhgiALKGZx+ZbaKkm8xRmNBKw2i1pJvDpH
HD5+Re9CjOFH8xrsc/Ttp4yLMDTb+doVPRkmOLXZH4jdI/aGj/KrZ1ZZoesdUmQo8qQpQjLuw0Ki
A36PAzTtcThfg4WxifXaewUU4A3f8dzY3hG85XGb3fndws3M/H/cDcXyfUB5lC6/MjFoyzQAKyVn
t5hK+2NgLugHvIknS18OWirkrtO4Cu9Jyrkc/TNfZETF5DiKnMDZHkJabIST8YRiF3lqWsH1xrdG
Jxl1gRNhYy7ClRLrDYFMU0DaFnPe2McU/sReejERucmNrqzeSoysrGy67C0lwCQzY2F6Ffqo/hZc
yy9YZAqDdXXcH82douSF/2ziATBf/EcWOHQlSNbfhG/7gfrd0wgWEE3+7Y0XmOAV0aeZVU97Ji1n
NOdeNxnBRbbGoB4iFK1AOXdSCeowJrJOApklpui77F8jzPb8uGaarFkrPkh2LJ31WkIADHnKtdwF
xSMwAH+BtqGv7GQSYndTFVscBXWtWyOK47j/olA0/EugNChqYyD9b+iuklgS5nXb3n/sALunHMfb
W9I7P1d+NLQgMb6YuO7DW/+25VrClZPH/J1TAQoEQpHpfBIwJRKDsdPX64Ip+6N2Pfj/7Vu08gV/
nkwGzQcgqtN/n+tmqz56BCIBkvZeUrWEGh8aiWZ487UQ6ZvHrfx4fjlEUZsTEExAzvtgiLptoA15
FFSj/1RaEgWeUU9jtYWNsqOmZ5op3tUm9ip8vK+aCOAoMgyi3kU3ULcj0ptqnF8c+WPlTmnMryY4
3C0NM+tOGVU2W2TXcXlz4oP7g8+AWdWkj7QTixHU9lmdFclPMwjhVh1Uz7feL4ujCYOd6WuXNQ/0
GwN8E3+v2Z0UCXXRzFUSmiqBcd8D2FcxS2qhsU8fd7R6vh9S0zt13PT5TvsSeKmGmIBJJseSgJ3R
y4K6EauciNLeO5PvK5vBNldEaTBBEbhykhnmMMEuLeMI5rRNnDkSlXwbe3hgP0N9Q5FMIoTblKHV
+nV5aJWUr59P+cnrF4cNfx3CdbQQhJGNUt5hHQiZ221anKRDcOKhvP2jM0wQkb5XA//Y0wxMfM8I
6zR0xo4KfcCPxINghzffc/3v+TuIOe9X7ZegVaDgYi1J6uII5ELs2Aep6dNVahNsi1qEO/awgsVq
xz7jTI+CZoKS0zCudEi+7Kt2aWyskA2zyib+YQkTnzkR7GmoeeF1DEqEPX7zhCqihg1w8PDqeYKN
Bd+ZQaBpM8j58oE1TqZSty6C5olYpd2+pgyMJz95Hrtt+9B320KwsL+2N98l5NurlsEKCbJgRDvI
WHx7GyMaWa0VBbdhtQWGeCP2rtbxEuD7xONeXxPjB42j5ov8AoHxUotKRuG8UvQNw0dsMTLMd8Qs
MlcxZKUoSiXLd2JXvcONrP4hMu9Zoxi8j3VRRtpBCky7uBGH9R4VoXuJ58TXXgpo0DsWa3VuriHV
N9PnJNYDug5hrboTBzlvJAukvZ+lxCWugyOq9gDcUEyyr8i4db/7o6dfwpDsMGnrQoNpEUbu1ryP
4+Ral3vtiLbwWD2+zTpakQ+bGT49uULhYWrDbzLheBKf982ZKcdXQ7ZUFiimAttUp5GL3fhzb6Eg
Ae9eevpE9OgqEwkgvZJtsKEG/D9sefj/cZesPnLIG3okRqt1E5aSivqxz/Rzg1ss3cSTjdMDxKrK
eaveNjXauFQWC7QzUQ4JbzqJWd1sd5k5OsQEdjeGDv7MAQ8JaHKM3IGetwmJqT+LneKJD9qAaNDT
d5Pn6XmSX4QzqbJy+eTzhJHlHC0y1vOBm1OOI3NPgxknVqhZZBHzIRQtiuTuz57w+DRnOF9JnIjn
eiBZe6n6R5ZOQoOHnhtxgoP06WkaBjALReSYo8/C2x4q9ug/95aDuK1G8mVbc6pAsmxhRWG25g4K
wh/cMnY/f/N6/Uu0/PvixC516+Avztwfr43v9O4O3gIATdZyyCegK1sKBxxYpMuJ0Bjxy0BRnFUe
gqcFuOad8t6lynoFGSpnvyoHfDE4ISWUDZ0toK8oMclA7Df5djmJaHkNt5yw+/GitwgUS40KeBhx
GbBTHlVDujdkGSZ0nA2GHBTTFR5AHE9Vbmv1iN+OGaTpiyEPE4vB9Mpigu3p5m1fa9nepZSV5tmI
SR+luWLtgqqOlhfhxV/PF1Tyakq4imKMTKI/7Uul0k1/IlVOPevKKHlszvtYzbn+T9bEetoqCKlk
/aTki3YqddobZFqrh0heAhUiJ3SmKswLzhkt25MOnP9/M2Mw6udaF5lprK2f6uBi5SgkrZbRym+w
q4x3ziLJFVnDqqtOYJCVIC2PgCnSt+CunII3MNgMYDNX2S5gpIGy5MXNL1PF8gEFl10WpvMr0urt
NG7TSax5gKCasV9KNn/jxjtR34B8+PIE0z/jK/Lo0atHcZYyzPx1ogbUl0QaOxQTBfSDtgUMeEAb
NKkpskNUeZQ0VkbYnl6eUPJmW39t/HeLBeoypZNb4beF0JRap1rWjDTZmCkQsnIr9SeE/VLIF+Ki
Fu5mFUIOm0XCxDWAeOGyeoq6dqzEumLsphjek6LFcY+AjRKDPh7V4y2VgeP+qcR4LRSGIkb2A366
T8EFluRYjL+oEO9vz3e+Wi2prW7HviFJdqQl5f9EQzaEKZDoMpSu0Rm6EaWwonhC4J3D2QdhA7Aa
b9AJezarMZbHuuD2XEUXezgfMYHVriHtc3q4o4Tz1AbrHyHjrVyRgqa+IMnXTEWJRurYMWwG0S9X
+iivLJirg/OQOhtPbCL0gOlFL+E/kwvTFA6VHixN3KmxlodKllMc1duGEzXT1hmFCJLQ8Rz/nXMi
O1SOI9tLtcVPooUsqc2HoeDC4savWpoO280cbwg/6iALNc8Yr2ky9GLCwQVXoqYw6aip49KtNQRa
SvyxucApwXYiR0AA42dwWJVm90ZxmvW56RdtZEHEik4cjARRveDR1zwYOgvCtTnoTpgce2Gt6Ri+
VSXxsGgNitDYcnkWXfUOrXyzddMNblQa2gjItFkUII+6deT6wnxgyipOibDZesTMeJMwZN5F8DiP
lSVHfFdubjzjJD66qJNUC8d+wSWdvX+WNsATHMTQ+/SsNMC+U0PqXMAHsRQrVnD2HfW96BmqtDjH
Um9hIpg3fPlCCyEGtQHfdcXEK1ZTVtjp8UK3s7tzZFP+yyoF/J1r5OBcWqBOWrKrtpehD2oTgKiz
/GtoUmtIwZ4aQcNzw0V9LfajKtIDLBlpF2uv3sZRbLRUe0YV+RzM9vG34FOwH457ANputmzNKmJ3
1Yr/6ayltJrCswfbd4ZHBnjZfxFeKR1HeLvbL55VLC1hoMzwHD7TpARQyPoLlg9bWtGiSublZ0An
QElSlZPWeLVtPLb3NXtuaXPAUQRLIuCkNVhbD63TXomoAmzXSwnpXKLnND3sADGicND+yN1IPmvX
+/hMj18rhce1IAHqQcWTUf3k8G7Pvvx7tF1tmxbswD4/EYreGFDvxsmQFJt72tV8qzveAeH0jHWs
XTj9ZSLzJfLslyQdMkryzDUoKjyEvFJDeERuiozeJZvZqeh1Jfwm6QBiy56srYu+cbt6PeerXIsq
RyodDDWNMTTdBuzAAisndaObRlmYXrl8hfZQOLh9VHEjelLAGtE87KPAcGbI/fRnHeGky8EahYs2
W0zgikOS3lHxEYVLgbEMDcqzzcTvirrGsYsPq6sWxHplSQbwD//gd9Dk/inC0lMdajdOM2mAu+fp
ny93thosWSPsqB6stgycoZoNb/nUsPbw1gMxztt3n8pv5VEE9GK5Sqe4glE5DIzRuY7wJ0pN8eOG
LkT4qhQl/Zus5IRxlVtzMWMOITLraFcC1FLxkG4vje4Sz0Uiuog+FuLvJVwWey6X7jle4R4l+hCB
ft80UWqa/s+OE70wWC9DGeTO9QvAolQKjcy7ipgTm2EZJE+2t/yNrw4i639qGiY1MFDMT5SHKJCy
+mteupUnaoMevI7Do1vPaWeZEpWvaho8YgMNOOKPbHcp4TdGPQui/UF2tC7y+ixu9VqNcKHVBNBT
hzo4xtupDDM+eUjbjpND7r3Pi6GhhyvL+tAdHLy9RO+F0MEUzYTg4Bgxjs7fWCK7GPCGED4ijfGD
jNqYNwNmCs9qTgXhKvC1DleoapWDXsyQUvHFd7sBjgc9QyXURl3Ut/Yd3dk0zIb3rHwcGbQRomlw
4IJleuA5WXAQYHStZmAG7x2SfeR+qdsY7z2bDCWYNvj5uX+Lc5yg7DqHtiwTAFUQvTv2/zQw8SqK
Rz7xju02R8SxymCJp2ciyjYbgtSgmIicgfDiiMQH52AKYFYFimwb3xKaXigf2obrFS+JYWth+9sM
nEN6HT2bYjwMQHFcgssXIG4fn7l/dp2KzimrIa0A2RWM5YL31rayC7HGBc85LT7q8H4XsB1d9ADh
2nGcwKcdSFeTTLpW11kqvv1kAu7oW2XR664zH0GQ0G7p4mUTvfZ96rvTmnB7lmKeQqQk+XGwtqBx
8hqEpxvSmOumkept0ev9kECSMJie30/fnaH+n5R/TAxNhghy03R28kkohRZWCI5r7SFEAdccWJFI
ZA3awXNvZH6RT8doYGByFqsJzorVpW46WswA11r8zBTyrXNUM10Uukv5v6alRA0DGt5GHgrUVEWv
wJQ4YRJ/51K/E2YdHLJOM5Ym3UGqcPAvqc3Rk4YR0uoXoyDK++ZuJdhjVYTXXb4RS72A9F7yMrnj
U8RqSTSnhFiOYY8UNUhru5289Blk9R3V3M3h4+u7vBSRRB8wiezFa7zm/Nb+Xbb5TD2P7Y/Aqzcc
IhmU1mj42EuYYvuMgcL13uS4MoS735I/KMDDL3L1DH+SZO+sD1lTPkC+3vLTRhhNqX0eQJhjK0zG
wx7520uIOGySmWexHRjwq0HLjTjD8rJ+KaMxIz4N5HO6/CSPRE3KraomjWU86uoM3EzhyF6V7bER
IMxUh9JiXHKB8DlInzZ8Zj1AiSGWFZupo2Y75jqBbN72t5otNKO7Kj7Gt6hOtuVJTr2HJldTcUay
ElSLAB/vI+sNwMkFUZYzU9cyhSUXMu+VvO0fe+c/5YHQFjsWk3sj6v8XMNRILeOFYnq/om4TBVjq
9gBEM3TE8dapuV1xqcmTKcDN3Qo9vgugxwmyXIuMID1oJe+guJJ9oGkzU9NRtTC7pa7tm+HORo8S
VBAJBruFNZ6BxF/pcaozZkTqsAG49kZSxMmSLQgAnY8C4H5b1bj89dmNfzJ6WsHCidifTZRp12Mi
Ehpasxwq0WYkvH3/G5esiZsXqmoOWKaQGHc38hvkqqLraKO6fowIYT24hVWVAMYy7o9klKv/rXsm
yJw5eySKS2BNG+nj+vfDNqZ5sHtGIudY6vpTLeWZWXqDaD4dV+7fYzR+F0WfRlKLMdmngfxGOqFb
zpzCDLRPuuuhyTRZuXHp7AD6SjTXaUgUZpWhin0znx8UFsXesI49YWLyF6dPvTa5k8/cmwnP3uRH
zIoGcviNbSAluojX70q0VSZ/EUeLREz2qVLTix7kbLbz1sfBRl3LSot60l3kmRDCztz/1aUpiDxn
/1u/4npancLcO0t+bR2V1BVe5JHxdF5rj9eUQDhhk257xYM5jZOSAvHTYArMTiKK9hE2gth+zY4I
PVbWRnWy5UAJTK3hlXPwy/Z+uR5V1jhN98Edw5L9nCrNfqXZMaAqoSL9rMYuf7GXGx/PN6/aODaE
xEs/fUIBOzQQnWHYctSTMoGfTM1KVrR8wF8Tg1JoCaU8X9JKWFTiEl+P2HtArbV9x/CUfOnGt4Gh
1hsW7Obtq1hcFQyIlfVnev1g4ffsQ5/MzifDkSeeVf1zwI7nrJe9us4fmwLjXOTVFo0tRKJJWdNO
D8MBmvit8OmtCQmLBMhruXMJRY32sWZBt5t081lmjgSB4Wv1El4N+ScFXUTfnBS1N2P4e2hhUZlj
YQhiVnDibZhGOj8ycmhfS/lQ2vJ1kX9R8GhRHUNs7gkYeij2V/UZd9n0KUD70TmUtmWTuryKaiwg
zryJmconPl2aCoJtwhjjRuifphASJuB2aHazwBpy/wtsXKAN5LDkXV5I+4NmzmQSRAF9XIz2SmfL
UIBhDxQuO8pdlUPBfo8fv5PYkFv4d1qBYWDys422QtecK98ZacgHW2oAMgWnDMKHQX+N0GzI6Inc
XZnwgrhZYH7he1eDSw1VsKMdHzMlb88uHqsOEh5sIOk9nrd4HzSlhbMvOihUB2/ThFNPVTptp+lX
nXDljr25E+53+Hy0X7HN7DxYJXUyRhnGT2ln0c/foRN+ac0pAFiO0TnU6tyfkO8K289xffMpV+sT
vllDh/d+oUdkNOh4qzH8qIBvoVpatbe+RVWMl1nR0OkR3LJuiMaZmiGDz3RRLJc8oQI8Jik4jQ7m
UVnvfCLAQDwfkHqo51XcdyHEh/kNDzMQan4L08FrHmi4c1WwnJHxpv2BVZ1GcapgVrrx8a8nNs3w
1w0SqAqJc5J6eTUETt8aCBTs6iIr0Ei8mdc7GDuyfIqHEzUQW6wYpUzM9TklIJMNqaeRIBqG6vVl
K1hGjbGPdHogCOW9LctpOazaegUZVFf2qbZK/WfhZwWoU7AWr2IK8PtRIagZ3UFyHSynyOkPfJFj
mL+p2ixw+DQiKCaJ32GjmFYTf7u96/gaxq+l7KzPpGQUAE4zWBeZUm+hiwEbxL6XPjhaba8smCEW
ryBwgoem/orbrRmRYbd1efsPmAMK7D28dbSV1J6TwOf1iEOPQ+4K7nogC7gdA8mwpyTg9urAlR6M
AtBqbj31R2c84cwsb/OZq9PGJD3B1/n2jStY0OHEY23/bwIHN6+bE8nCP6iTZHTBygLMXeWDJ80o
+KW/8ZkgkhAEJy9x6ihC823SZ+oAVfC+uTmuu7OY+bfErzpKL6zUwzTqCxPZbYyqStXl1A/sl6Cx
1CkBSaSPNBkiXOO8k8/eCek20bIaazp2EmCFTBvp5ccge6bOfowydJLpz614f6g+mpQ+oawDvciM
qxRDs37wIu8w3E5QOtTQsUNaIK4jGXhYfJFPQnFK7zzAv2bUoD6ocS7LoDuZ1ZIfXQ4O7rgVt3pG
r/bCy/4aWbiYN/jzWfXJpVW7JfLjzFRZtdAoyu/l0wVY0sFzq6sj+gvobeT+WadW7D2WEuoftxcw
kjQ0JuFqpwCKPPAaEP9wzLVmXoEg6rtnKZsxL2GmFjjLv+esJoozOYzB0PFYv9ynjh4vEPfS4kC7
VfC7+qNxVJQIcv7++LB7QmROS54GQEHYTHLaRArBTU1Zvz4CyDpNbHhsLezOxCKek+/H90lnAWzE
lwptu0w2PyIuT6fpgr03S2l/mo+FrDdfhgpGL3cv+id3pZtD3g0U/s3wwO91wMh+jXT5u5Zpbn83
CuyOiSdVmI/YUJg7hoNkuwxUqmxwvfZ9Y32CJLIL58yH4rmBDafikkYFFkhQU8+xwFDUvYUKGC11
vWwlM/yd/IJTdCU2JvCo7j0S46ikm4iXFpWxyOUQSzAE9R8hGrnunPsDr1XKn4BH4eQy3EFwuUPS
qe4+a6QOMHeXErataY4EN+1HUnQ6HdLZdAU26n8Yhew4diZaO+jYbjcxyPju+DdQMIL9/BsAqXcY
SnX75J4rULMza++J66mOyZxAzxXp7+i7Pr7bj+C4p6RUYkVR0Mp5iNio6KpJwpTvCEGY4OAStepJ
Xfvks8Zv3qvIIwTj3xL5lWrJONnXA86kwtQgi0n/Xlshe9ZpUysBxBcmD00/MMIGZoEVTYAwH9U1
8kCgSXf6drpgfGLEXKrre76t9oOun7bAKXo6AyrU0CBMU92puDRv81wVmxahvP6qiK7Ursak1GaI
VbLjXJTpvZdAc8QDL1EkAtV13AvliuLXHniZYkIYYG77YWrETvcwuZYgIR2pKpr6esHvDqHCDhSl
eYicPZ+pV4VNlR1xbsHbksWtrjRQh6zNlq0ZfXMp0LAc4IhEMoZC6cPXd+xwNnoiIu6rc3sqdgW6
DnuSLsdCIVknNLEqAgZsTzr5FbJM1gQoKpBaYoPh4qlEVXuOaILk2kiLfUAK+bG+kZyk5vDZYdzy
OsOKANuireKkrlkr9BtX/zyVxUasoY2lmrwEUGbOkXF8RLv+64gwuQiDYM0il+lKceIasNALRwpJ
bxWkP+yNyzGzCc9NfXxoRX4pTx0MO7s2qCrepFXzbKw7db9uvTirK0VYnR5CFuFrFgD3UDSsPz2V
JUMyPLw39yi0wa0nU+EYTn+o1QeHOO1fDGalg2XA6ddSU8LxjGk5lmaIqyvMZVgoCu2eIDHFciXL
qyCdG2zZCYN9PlvMUPCMYpRvGxwqlw5IggAwDuU7y3WYNr9wwic4Jpbw+0k58+wT+idr+Vj2ECuv
KLhVVfyJObgMGPpkkojqHTWfv13+XCfXmj2cH0sMxQRym7PIkzqWzAE5G/xKygUbYhZVCBIHwlKC
+Wr04HtFOeYJSlnEHPeIgdUvrTr1yRWbGqmCmbI38jxrDRcL4byVlMZvn3IdpXyAku0RdU1vfSVR
jByF+J96D60Z/Sr6KPcWrWhZnbw5TE6c7sD2EynNe6MH7rmi1vRFIIad+ajDsoLcdv/y9MmowDNx
Z7NpsdB75egoA0YE8IbCRNnakKIS0tzgyWST0wBK27aTafQieCOFwjRCehm2mwLOznfuftk/yU9s
URPEbBKh6K6qcu1oF0HAT4gpDIZEvuL8L8lEdsr3lbHSxFeZVabspwTKgN3k1XfJxKLDqhY2VpQt
zFlgpzAF+oYUFBsB7vFxGHN6T49iD84sgfUOhCdKB5s+840hgaBuicB1j9Zz5513XFu8oSNUqAa5
b1JbP6WCvJAJW9wKtRhWGmHoONE9oySMH7lcvWyiWr9w82VFggURZSvBfn1N233engY0i09nwaHr
LxT1bHA/ElM2jE21j6VI6E8jrzCBaL+jh093vgmMIuFDhmjZgW9xU/pw4RXuFPvazMnvTCQZIlCm
ce+AGjZ3s7neJilxz4b9TFawQskLUNlOpKPQPS7nw1ntvU+T/mF5RNHdvkc09r82c7j6aJX77mCY
dsX96TbuaRPmnAtQH/0+JE577jpXvvnMZ8k+4c/5WdMMLyuPIhhBQxtYDbHDzn2UGjjTBW4YDVCg
ljR2VWwIy7jr1OTWlNTvdrEYzGGOD5FQiws/2hNU7XxcOcVrbNG9iR7tweT08vE7ieK1z2N+knUR
uyjX8U6OIYgu4td9NC059YuyaebYZFuSgdQkrnB4Bg8hTFYvPMa1LW1hnYhHGEK1KrvCmweSHR0g
69FvwqIpXD0+s4hJbhX4s1T7CIIbthZ60AVJYIRU0+iNc3hmwknZjuEcTYJrht+esNefruq0Q1bg
R6TsiNfnevAlEjzzGCwMSWc76Phah1xNyGkJcdo1UoaiP/rZCC0A6J/pWj4QOn/R09rH7oNlks7k
Rr9Uj8JG1d1dp3eiuIT8Y5+0rkJ+yaDxatZCcmbgVLLJCW7M4QXH6OXaGD8qDyjV4rUof1x97L2N
m6FDu0+V9+Ixf5y4Y7gqn1N1ZOL0U0JT5nnmQShIvbeeB4ENB/5owf+zc3rF3euyLMT+VfSscMD1
YvWuXBojvgJfSBpE2LNYvQaCB6Ok3Cedk2hsJJwKfIzxJPd+PSSNPSJNKXATk5SNuKngbARXJ2g9
BN57n13keIMOvRNzJebyAqX7EAh5UGizLLLsLzO5v+c7qB6DUvWetq81rz8nidjVlMPpFqJ8YRf7
f4zjBprW+4djA8/Iqr4S1/VK4NpAPzlk5QbCn/vtkSWoLDRwzkRUgk+EZKNJvTBFnUgHmgaJ+c50
BFBFwC7UTYHbFtsxdQilEZatiTPHofF+Aj1zjsBMiYof4jUseefxClfF3vvA8T7ihNeaZqBuI3VK
/vf1fzT0UydpIDGNHvrNTrK9vMU8Gdi0FkyMcmCQTwsTXvcgwrHD7Xwn7bkGY4PWLSZyHrDLUqkj
dku4WC/zWjTdOEvlBVc6dT88oUyQa9EyU1jWVe8E4ftgpERZbS900k8EFk7Fez/Ytq1Cf0eYffA7
LTZvUuCg64eHyMrIZtGlwEUYdrlfZ6fzMMgqemIamJPdQS/PX2xd7DfNUbMSNFDAd7gTmVTsdn1e
zU2jiK6SEif7qj+j8nfck8PwVrRYtTuTw6/x2PD6Cbk7Z5dtUoYWZcPPgZBhNFky32mGZuI6JGhn
D+cCA0LF7x7qjqXqpTSV/BOIP7HmWmK9tef4AmulAi4XxWFossk8Z8iugsjdhmUPzbLJlty8ziCl
Ym1v1Meds+sQrI8X5q/FqCzB2nH/DTYYc+0NRemuJnnNZawaFWxMPPM4VzWLPc0H5hHZiGSymF9a
AzXZtWNbzSvOwULeX7cZy3a84lNsWo175urMeZJM47++nq76UGMEZ47y8k6yWkz3kbAzovIbDwhM
jywppPq2p1O1F859geB/rBR2GPtNT6oszqZek/0fOlmIo9HFuj0xsSgW0V9oi0Hdg6zpCpQG/dmZ
Wg+h0x8z0kSOLti6uumVfxMEfwTVksp8R44A3p7GDbuW5KXEYJR64lzj8ZcF7e1Hg5DjYvgfS9iH
TAARxlV9TOdJTBrxchZOdLc3rsj6jBlG/EvVms2VOO6BEr+1AEJ3ydOSMgyMmXfh8DrAunPsrb0U
IcT5u4Q2iI108EKWbo73eYcwG9LBd3v5qxtDynRU4kFvWKyOeldCoaID99BItc/GjakHNHFEvPqs
MbagKar6bawcsc3s3X9svO8x5aCdpaGarC0j0b1jlLmcYY+NwkpXXT/Y0CfWt1MX3h/PBbFRnhhi
kk0FpNEk73FrzbEQuxjhK3/DrIMNz9s0PM3Ysl0Cq4iRo2EIRZ/ZviWUZxAqsgjGn39CfyB7mzR3
FXsOjVhnlGQN7jo3pNVU82P2VGk5Dd3RLq4H8rM5AIz7rOsvLmfMcX2yRjmAQ4KMzxvmNQgCUP7h
UowBeSb+ZeKTPUFjJLyErJ51rul3iPf0Vm/CYjxICUQSkIly6oBByzGIT3SevD5qrRLQQMifcNQi
osDsQjfRktgEmzLwSNaccNkKwSTRcq9rbZigFOTEaEp9mA0Sb7fwo4/vH4fXuOd6isT1yXBETuWi
hCFMfaNPnqE+pQFIxHcnMvhExcp7ULBK5QuN09cvx3CuPm078odab0GAVQa0c8tQSWkO3+X5fdyl
oLFGHZ+NxIFvTNLtE/1LjRvnBfpnWWo1Y2WtET4Tpc6UPUsFnI0fq/shQYwk/qc3Z74fuJSS66BY
e4ylj8l5XOa+5B18EAjl7TOcAsL9i7JWOKVZ3hdwt67YChYhnwwGfU/80FaAmRDhUPgS5GRW+Krg
wCXosY+dRO0b9N70tvu9+L0zehk/q3VaC1JS8Pobsxm5BDJZ9o21hcFaMn8e2E/BGt8NeiHGmqeY
nyyqMI9xudQYuYFivTwJy7GGwp3z8iZ/yhP97YjKvFW/Tba1mtumiBQt/yrN1NJnRieGQtjp78Qa
c2wWD5dCeT6FIXUBhDk7d9wGKKf6m5oFsgl21MEwb9XySQH7msC2wCSvvGvI2mofiRDCzROpkflV
AAMM++ViQ+f1pRezalo9Mp62RJCg+MHgV272/bgsL016ms/MOtYuXbDXdwaXwO4uZnWGai7MtoSB
Dlb3nFv5ryrTKZn9dT64wS+bxR4vax28Haw0qGkGSTumpqER9vCi1Xoq5DlSVw3xH/5VDOAQRo+7
H9+OnaIwo7TaKKUF52EkqWRSE2FqVC78XY45uPb14+sX5wggxO7cyeNvqQ5zce9tqPJZivqUJlcb
Wi9hzgxwGRhle5AL0xW1/HJNu9tvfLIFVEs8Wn3hcsYGjgCAJ12nOgUKq40EkWfWEfjSgiQ2F7SQ
0VRa3bbbbp82tQ2DMuK3JEXJ5bN0jR7YrqJCZLFTDk/XUBq8yBJD/Kw1vYrJayv+gRsP638yd2vw
QDnUNchBgBVA5oRVJV7OL8CQaRjxEusJ7pNSNC1YWGmiuyMka01LJJNd/YjpUpDqI17C2HjsIuyb
v6qK+D1GXYOrmsgOX3v9u4cm/GnfEIwTtA/IlluZ1MLbNyil14tkoPZBUgTG/sM+S5I78SV7oMq+
rJEHPIXCPdqOnAPf3nE7StJCRqAtxlu58vrEkmrThSpjYQtxWYSqj4n2d9J3N1JInnAjENcEIcnn
YTCGNPKvGvHD7aTJYzL2Nw8IDBemcMd/HF/1JOPfVJa+CTloqyvsMUR8fgXMBEOR1zEs+tBdv6hx
L0eMkS3srkn5NyWweKBFkjdcA3Vmsw8R5iRtEibXX8kECNwcJYiwYqT1JNCWHyxRyyEmDb+pBXbk
zK+BaFgANfWCHadAJ7sHlFhvyiMBA4br+z6Rh0XLjVRq6H1SmqXxOP+frSAk3ZE7tM0VC+rv6ONP
cnUApMJWFJtGQzNVMhjg0vZBnGSJ+9N60G7dTknXKvGNogNlApvMRhSwI5zH3D8uHOF1RirzTFzr
vOh8LdtTkPq36Sw413lC7lGC65xUa4F8XurKlFNKiIO+wjwJCpJ6rmZvBso6Nxy59lrYar9A22/k
Mf8kd1uF1LU7qrfQ3RTkK+p7FXPX/2uJb3HDvK+BM0Au8Qdl7S1hgbsKTT1T+BZW9x4Lj3XCgGBI
vbtCTjK2ydSiW7VCUYClATTvrbe5f++Hpsct8d771ofEaVjOeW/lBWsBSYQ9sCAHSLyfnSlXHm1S
BQl6KgVT/FLjSNZkSf5zNOv5I9Wr0JKRoUTHNVGv2rTlk9uZKfiVpj7y9qqbLP9tArXyPFa4cTea
KgBNXnmlgfh6ZykDn9c6HimomZuxVyqP6c8BhSOk9yLFmzQ8xDYktZ6Wx/z7qOhblwWVnF9cQ6uf
3J1Xan5nmaVKA79ICThyZ3NGP/2AEg8VPij+bq8n1X4IQLgl0iEiguv41NPfzY2D41aEiWgGxc4G
Ayug3NFm6eAEBCQeazqKI4PkOse9RKROF65myYn+cE3ztRIBGUh+4cLplGf0hK13v6Yjr290aqyz
bvMi3lQ/9a0x+gnFJakbC3WcLJWDe7wqo/oWJivaCElnfY6GYy4RO9G3GXjMvNswbpLRP97TFjbk
JHtL8ZAPHj3XrcY+MYTC+FnSFQJkkSpEmTZYlyRqTFd/5QwscaBE1+1egcxDkm/RUVveBEjRADhB
XMITVZlXqpJk99Ir25Gj3IxoWaRYce8UtJSb8D6zpHhjZD+Fqt1dD634niCoSP+rNgEmhHwIuJaO
JwalKci/j1crQpqht2USkRQNPukPYcxPBRYbF/sXaVCY3S+pm114PxYL/ytIzJs/p7oJvDvRfIXh
EVQfO8P7Mh0355QS/pr4OUIT4/i3TqRmaIO5HuJyts1PVBiwqs/pj3j095tAx/rGPJcWShaRaWsP
B2Wd0i97kO0v1Jp0Odh6spcTmL5WLTqz2u2mWI/EdnnHIjn+H5hXcAWihJys9xK5+PqQIFeN4ETN
BqKUoQYr+uvSsUMZ0l8Xl8T6jS+JGQXVfl8Ib3skxYCQbTR0tbNCbIOKj3LnkmH3asJEyuc1Xarj
f0GcwCKjgH8nP2pZMdkFyGqTKuie41cg+JXJXp1yJ5W3BTq1XQtLyDf/djeoAOCcRr0gpYQfad3Y
G+F6RwVMShPlItwhgtbRFCtaApzIQOUS4uFHV0ul5kUYsQNz3Xu3gaB+PAg3E998g4eH27EoSJno
Bkwh7dMrL5/4zKiHTENyTGQeLnMRS4YGeL5B/lFGabAlZWRNKr70HO+snqPqhI0fqexIkCxCRmfj
2Xph89VtXJ60TnqI7PKgIceaMvr/z0FTm4SWuWg9dVcX5pz8pKwoDAojTF4ULB5UmSLXPQFVVDLj
vI/yONCHRrKtAKa3JnKzbxfL9e3CuY/PQeoHitXpmOKrc/z529qoOHaHjtFaFKe/oZJ4LVN10kla
fggiDwLbpEqKinEyNejVQzLJtf2VPHXh8lVOcZa6Cpx/IZ/Y2Q9MZyhiK2CMsTujy2ZnJMOYk6HT
mpKMHM3UeP7aDspIJVeM7G+rvSQzwtXI6lZH/vaunN/hbpevlbqxVFYEaQKuMAw9mEfEgrsIyaRx
CaPy63YDKMjpK1rsc4mBLx53gnGfUQGZOIU6SMFpWDWDwO3WRIofd4eR6GtZgh04Jd456cM1wna+
i1gEvWPUqRvziAbtThcOgLSmHl3oxu6l4uUnzPQWUlZMoAUv7/g5R6JmhJevoVTwI2uzG1nBakee
Whva6UDh8drKCUEI9TmbJOG+RMSmyzIaSYt80eF+9ZnpAb0+npcfhGJvdyBgVhlxdqJGm8iEKEiI
U94qMortlquaIg4zEcFICC7EXxw8rOq+O9XF6LCSvdqXyrXSmN9bdmECVte24RoBNe0La4tQZkvE
kCK122HuXyRNMaZy4fiIK5uu/kPZk4Of72Y3ZeD5VuAMf61HJhlvA5jjF62stIMMXvdMLINf35/Z
P6bA6ftIgoJIlth5M74TgGZtHMsX9W9giO3kqcNbo4EyNbIYHLGGM5PBvHbq5Xe1T7vKXyvS2zMv
WxmCtA4C05xy7Xn5v3WozFJpovfWsvIptH8cbTAWRbAMAAoGvJPNYp19iOz/E39x8QmU94dyAWjC
mstsPGDuv7x3n4ItoFQfwQlLkGtjzBZnF2/xL4SsXMwhPxdStr9J9rWyecbh4cPhEYExMKv7jZ/t
olkD1YPUzlOtba2EwTb6f9Osnlr2ZJ5KSHCUkp4Ga60GAvTnDzN7m0Ljatk73F2HAz9ruOB+PnUq
UPCqrXryGFgJHF1gesHTdZRNs2evmJ+sIuuu539dRPimJYnsdrgs0j6ImpQUMJUVyW2IzwagNFJY
2i+Sh9YgjkH7YYyY4Ef/8C47/yZGeeBW396dZmT8zw2ulZXiDevAVqngqvlbd13/Q8MPgyFBKkPp
L21r2C/krm9zyGunJKpGvoIOvw4xqjpXdy2EYunmnaPHpaY6gUTaPKtnz1uj+h33vAhpwFSBP/tV
QfKK3/R2K2HBe6zBAmjO3xPgBIdiDnOlh9YQ0QLTpjKdjLp67Y9xHiAaDAHeDGN7XDHnR1VlYoOd
JN20yOISjOHetUuD8PSgDHu90FnA8rEkfQKJ6qEMLOegGOmXfZbuSZcbWt+EstRuZIoO1CEiVEUY
C251bYniJMASt0VuZbf/TnhC0/ev/dqytHI/gRpCKKdfFogxQW1QMzOigdljWjXobP1iOtbYVnNu
cKkoS7crZNWj2V2WcdBicEogKri2uWA0FzKd3ykbAZFCbA43Cb6ercvAFVxKPln+YycORpCIhUDG
S608Tl6o5rblgnCIBScRMbBSkHTSDK9woIx5Hw4f46GDbbQpbson87dHzW7ujNtetvAjDvWlRIwz
s0N4vzlN4hmpBmMb7JwVJkoJBNQvlu24ltKTCK98Mkrdk2e6R0Y3LlNSdXGo4UM6clGVUSlE9vLI
dpwtuuG7wRuL2iZvWM5GuNiPh0LX5nwMYbTKjkWV3S7QkLsWmm9sHuYAQSpbDX/hSfG9mvXbcxdx
uz37OiV25thiPThNIobCQcykAUAdSyOdZgt0GTNbkdBKhUH+N0SOp0QckdGu6V/rLiDUUcuns2WM
avrQsSi1QFTxX1wcFzvCnmq99q1pNpvyp+x+68COvgiOh3t+roRugqS/7lLlTj1TjRHGx5R8Oz5l
X1fR+6IY1J0S4GTRzP2sPQs7FnOGewEiTEE9AQj1WkHb6LKqh+k+LlDBIF66oZJedguVlLwZ7l4f
szfvKNzeeY6VJ8htO1fo2gCRHxWZ4wDupTa3K4rZejdzdFOXVpTEZyxUctGGLPfZqIlatVULiXZ5
u23SD/FzguuKhv21R7eW+WUXMZN+KFS4/8jkVxc7OUibOMlEztnhSAkPioH4xzQZk+r6l2hc2trL
L0TFbIkCMSHHn+XwWJe7jqIvvjqlP0gCb6EhrGsVfw06ovLRr+fG6p7NFh1UX4OR7EXQ7o9SG0TH
KUCRd9DuuF+gb7mVZyuhg4qBOsn2hczXUa5vBT+LQANO6xE8fwU1yvzdio4HsTg8cSS+47ekldn5
/XeY1zYAYAcBjJ9QHUiU5mXA6nGBr6+TTI+NKRd2+MnViTPZk7nTT0eW2zDL+BtTLZuwsmaJ4NEh
eHsClHh6xF30Tepd2ZGiH6fIxuzVG9toDce+8iVdgJgGM7b+GyNKaGhXkyMKzZNB0zFkzGzJV2mk
S+E8LCDOiX4BcZP+mqKgqvBkt05P/oHHBXAIr+0RzqTUB9UUDrW95br+DkElVKKtNiJCBGUW96SH
jvDqTgKM4V8vs4AKoA3zcJcRsHNT+lhjzb/WW5lLxotKblvBzzfmeesbRb/wLFHDO7tBRgkPtFKd
nHn5KmjjlJaSLo0lnewizc+L0RGpCKeoFdyovUPTltNEXBkh/9GrhVB4Jt9UjWqh66Cqz0cG4PJI
xuHzg60hEsRjV2vx8vEwShoeReFpc2Zqv+c5So2Kga2zhM7NvuGZT31h71vhp6eiRx97I8h3ywvN
tKkgBMOsrnWnzJFMX2Y4Npp3sFfqoV1sXdhAa47z0PgyNZElLK0V3Prex+MdrMEHCswtNTbhUe8e
zK3txgOKqLgGZTiCLJRAaPn2QTjOt75ZrjkeJN205cuFQXvTC1seLf8rmY0WjJPSWvooc1bax+aY
ZW0UjV3XeEnNfK3mAwc3fh3BRZc6mQlxxxymXyHmoFbwveCC4LI/3C/2C4dV2BfPs3fGUwZdOPv4
RvDGtH/0ipQKL7i9ODP8hbXq8/Ds1ubrcMkCHzExNdtCudfyBiOTPAzHB0eR2ooK9OJ8Qj2glIN/
owdj1xAAOnKt5oi5WjmN2XDwX1fl9pNCcbTuI0r8umDufGXXdUn9pSK3BY84+uXbGmGc/wf6miOq
W5XCULkA87/2dSOQ3dlLcH549OVR6xEtmovDTLeVgtou0RjZqX7vC4ceDZriApp5YhAz7clKOpUO
kWl8JVAgEbZCew9JhFEr4MoRudOSxXWPx5WSgtXNFpD1HIBb7Vlt07HRd/pUBclYkDY+qSVJBAf+
yW2MibTNrITrfTuQAuV1ScxpV/vLFN8SmFvDmMEN1rYunURPEu9GkxlOnBlkmi7pupLSzBwPKxF+
e0ix7Uln25JR9CJpt3x2XiMsBOG6rDmX8uMhxd9/SmNqklZD7ByaQn8jSyc4V2t+CVxf9DZHjTEh
pjjJZ/vuqLGAD3vFiRIAv7mvagUy5/cNe4W35i8jVZRu/TWyZ21W52SEHHkk1ZeaqfHr4kvzUbwt
tGv1cSKwPzKFtpCNykSDOd0J84d0K6exdavddMv2WEbeRL2CG8vt+gDYvRutiT5UAKOjSdO9VpVi
Y5x+3Ge04dLgHnyfIsUeQBXFgzLUnYaRZRniYVmsJY4EM1aPCwzcZ7UXdK6PKz4TV0E4Naj0WecC
k2nGe6Q1w27TQ4OI1EpwHKK6afUtWoF8lGHIKYqJNQG+BryCUYsD9bd8fqXL9jd/SsXMTNNruYqP
69DfwKgN5gu9gigJmWgmVn98WdUquxy7rrSqY4HG6//I9RGiHMOYllNv1/P6mBac9apvm28nanGp
IsX9jePB1ZfDaw/7NK95TpfoUn2x0PTtAtUYLM8ye15iCkQH0JNvFOdkzvpvPLrJgwrpqZ1wcF1h
nxG3QiwEy3MsdiGc8zmlFf46luyEvCFcnETBC7L843JS3LgoS7ekELe2iy/qNgoKPdSWSpZ7Q++x
EJI2DdyYVFnuYZ2oXVyO4ddOZKyEYq8IBvVneRrMk/C3/Yr/HylWbDWLVFDMrt/iADmbtmwrP+L0
JuniRNPP6VD0cDcWeCMyZSZ93pbdOLWjkm5+Y5CP600k3INtbjwAKwAUfRykmb/IMVOx9j9eZWF/
EPMBQdFmpCbs2VFTC4WewLES1ZZ0Jp7ryzSLOH3i+T9X366N2V0bH0Oa5CRE0uBxjG4Lggl1bTTw
faNObf8h2DXDFe6vREDQh+h9EIk9q14+Uy8zgNz+n+NBr3AVVptd8f4MhyHYYE0WGA8ZGnfVRe/W
AAXts/kPg03PDdq7TBQEeexnHCwtpnVIn8jtlHZ0Xr32gOo8X28DqtOxTqQs8GVHMQBoTkwqtGWN
7lYMINM5LwzNlTYpA42O0K6aCQs39TnV9si0akuTg+Nqq21kqSgpjkrp9W03FumqQ+6FkJOCNise
LK/ERUp7QOAV/HLlmb9d5k3j+yu+noLnwlKeAWuwd/Cw2NOcXHApCygBBmA2ZHfL6icJCW5RhZHU
1e2ypTJzm/Sigu/I9LJ5q5t8My45mpTzT/dmBSwgMoxXtuaVolMVHAUJkb+70FXYrP9GlPaEh2MR
1UvqIgKccO6ZEzI0iAApoq5QnpGNmmxZrLyVAj5zLki/HlYF+AL4maCKK3RIlmFB9YEMVQ1L2qI8
2AtjYQ2GN79exAyME97l+JN7Z97lKmJ/8ecfZ+ozzVL1Ge9q139eB4YE2JHdsADtIxCdJuvlNgR7
krMfFolZbjYLh1k8k5KBphJYXabcqEtQbNtjOMul+R0Kvjvg565E/kcIvCJviky/8MEWfbH1YRRg
ESwLRoI7StDfKsdoXHHFKsV5XRcQw889wPXdUJnO8PnMOvEINy9pYvg/uO5NPd4k4H6+DISsA/Nv
shhmaZHpZvk4qqemoF4Ra1UPAexFrdiH3TRbMlpICqOGbkY9mLTQf0xgUDVGvoNg1YpyVuv9XtAW
dT5sKCvFJrW3TeRI+tL0NFCWpL8p069IIBxtRVWWkeY/11B4NcyUJJZb5HdRg0NB5nCqS702uTdD
qUhZEE2Gah/eVC3EDB7GJKY3lXnwCIp8KsH74YdTqOGto4QTxLFcsgWvNRueNJ7ZBm9L5jCvAZTo
fzgaUEuhZpnY+TbMR1m3j1LnwwpaeCX2DaeMHn/HGTFZujQcU4u8C68H8WINPJ09LneUSftTTpLZ
C7afF3AHOwZ00hy8vZh0n53vOolNG/TrY5FQ0HCgUlwq6gXREQt3MtBDyZIHOCxAKrF9VZ3j2wX8
HPjJfD2u2v8Tnqs71VDQDt+b1p7Xo2kNDxIBXyDy304KYwBjUfH3e1w7x1+Jzuy3+AHNr/tyEm9o
7Zc2009W4kSa323m6rp+EHyl+WAjbmZi0inIt3Z24yw2Up9DXUcJEtDxztOKFp5PxyQ/5VFD2nHF
SpJzl7Qm6a8cWSbVULaTKu/1OBhWp2qufQ8QX2uQkg3D4hwfv9Hmt+hdz9weJ0KLyBfIQaEZOGBD
yRTas2fYxK0H/kSv16YQ7tlxB2OaZObfA7/2Oc1KUVUnwb5aQdZUl+wd3jxFKmA0FeuZplmDYMKV
JxJIg9RhrZTfhuZC+55UgKAcZCiqDCjzDelQUhNRbGhzCIOYGel+nz8njOJbGZHNIzoWfIdAxxQk
gAks0OSbYE8RoSgYgz2IpFvvM8oGn+CCJ0LHETXVbE8ehNB95QuyZnOyJzyP0Rx67aLQdFxfofm8
XTWB6/QoG1BvJ8enoGd8OrM3X4sVW+P1VavLDziO2FzWiXp6mxuQM2/A4mDY21MAcVwKEa57IlMH
sjnoGOY7k24gC9kq6lmgT0Drt9AF9SipyhWN4Z2YBMlss7MEvP5YklvqKkNQa7Dwaqv7Sglg8E5K
Dag4tr6yXA6f50LMsu2ksLHRzBBJACuKF18uVIHUqgDEGjvMuLkTpHlkJrg3tMXBFMeY3PBpOl//
Tp070jpEncPcXfLa3Xu+z8w9kZVW0E44JOBWOuG3G3P4sKq7qK21US0D2R1t4KdNwNmFBSkAdejm
8a8EOK1guw2PQBKHqDaMWgrb4lmgCtCit1tpbJwVS+E2iKW+DwinFWWFBKy23jF63x0NLpbrPO77
qADf0CrODD/we+ajDmgBJcuXlL5RQXSa93RKMzBeJfXR+2KGpVJEj76sUIBcBE/zygWLFw/BHkUt
XQ2jXAeryM/rKVOFp9BrySgv5y0Qodzjs/npxPIBNUmw7GMlnfOdGwSzedtu9Kijg1gZfRnoliFS
gxLRAyB98g2URVSNv9QyxDaQhYLWh48JHCsghqC2IP3SsvL3k5J6f3mjMIRMAhVdyx1FSmEpnAHT
8xSIe3GBLIkiHQqCa0KPgto20dc6GvDNR2alFKaTErAPXRtrsgeOE7twhSfjhrVpaCIyaQ8quMMZ
8Njc6OP70j9oqOfQQVdLeeD6y90ze1+hI3tB2mEllVGKRnZlspybZWkmm4kfiLIB5I8KKSkAKCdt
bsUr8vH/965HCOUA8HIv0Ajs/lBXlBxWTXk49MaE79TDRjLURzzElciJ/ZJNSnSsj8VPF3KGfZK6
knrzrsZG7/354RV653biFW/zvXma58unABgdZQ2JPKYPGQnDqUBi/iP3PWhy9WzPMyUmZBLjyIXu
GLEa7ac4iW4u/soTr3RuMncxXkcWcJ9dnPTe/vK+OzrQyk7bzrNJ8DS1rsjuTSByJFqrQc5sLGgd
kGTKhm/70BMBCl5f0kPvualrFNLIY+BgRV/wg90rRmQj3UkoaOiBaj6P3NbNkjiqMCw5P0nIv9DD
txvy16pQG5Vzz1FU1k7h45uG29G44pz+QDX1f2siQInV/0EIWjPGxRBrfnJLT7kYvXWhJO01QuCM
xkQSjWut955v1J23RIiJBYqvkLK3WHuvZKCO9t8meR7IE0JazSkK47FI0rW3BK9E5YGaQkjmtcb1
c2su8HGdxHkFXDXeJl4F6y9J8vSP6ioC85bEME+31qMvC0+YQtf1/mPyN5bJGkAF4x1Hhe+xQqv7
xiBQKTVlDog3ZkDWP+MSzT2N263D/xPiqN7cWyxLO2GEysOE/uYBq8DR0IEzySd+ky3Kzz2efo9t
9VNhXF0EedFbBDMEdhlqdJDxpGmVVgeV60JsJN+3mGxNz4++sliwkn+AQN7MvudtwY6ObLikCYTi
6RRWMbsQ0oiXsbX3rQGUrGMfbR4i6rYMGr5XmNKIidsO0O+3ErD0y3srPimV+w0wruE3R/TRKolB
4Uaov3WSgidJfn8naERR8hW8bhNDAiBeCPzAyLaSQ6NLaXp6vSFXFiMxBhLaxeF3vPA8FvSEIw4o
3StqTmucEYZBKqSM6gO24usQrZcg1tfKCsCJHnObQ7HCi3K8vCw8kFPGuvC390ljE6pgJZ/avM2h
dfrVn7TyJL65n9HdFhGQU84rpX8g4xqLzhuYIT9xt+Q7TOFF6h/ZuyS5iUDpAp3p9p7/Y421H1Vd
isLS/E4ROTlGiUMSBLhHXD43FsMvc6D3W96UyHxAXpthPKaB0EtvYYdpxqwrhW1qooe6pYpCrRpX
knI7NCrLBgxljhcqFZ+vxgcax7WVhsxN29YQvMRZHYR5P3gQha93gfGu9wMTypv5XzbWqiZ4rFCh
35qDwcRLaY8LkEkMl1WFHXwP3bCmy+jORdODPt+jXNBL7lNscAjJYvDknqiQaWIMDcvAQG/GI/cy
+YBCwEub2rkFrWsSev/8JXLH5MkI0n6YlRMaqcVSK4XrPYs7ZKQU+/k6UH27RdXIzgVYaXiQiovu
oawzpR7DZl8UjiY8ujpZ4F3Kgm2Yi4c6rCPNBvCCvlEJ+YlrxnAFLEeOeXg29Zm94MCxieHpWsTV
pD8/3Iq9a5/Zi4pm8oiO8bWQMYibj1ONaI5fgarWt914PQtWFuvSfZw77bXpu0bs1lnjaRpcXi/2
y+3MkIQbejDWbxGsmKJL7+FFD8O+vHV/n910qC8ewZBs2nNcWOzzNwV05xJv8sHITaBXiCt8/3iU
8pevZdldrJcX5ak8W9/17fFN2uf/4lLmUmEbCOz6h2CtygcU+4w1+TysA7K6Wu2yJQvu0eV6XIa3
sUIJerict58QkQKXZcu5WMPALl5eC0Wzy6RTxLGLAmN4Shmtr8U7/dM7tcyjiPixw5V2vi79GX9i
Uz+SE4/pIOKPHr5i5lBPlv+JOKNRzEjOEbzgqm1M59rDRcE0n1f9ix+ur7B/Me4Uqlxufjcp3KVU
LZDsruf0iVOsiGQF8FBKfdy0gDJUOGZAltCzTgAZiMRQRGIi7pLuMd0dI/zcgmt2Wxnoxnok55+M
6Ufo1N2iOeezPvocJCkItYPkgO6sSzdeuuVIctN7ZpJIc8mNolWcLEgmjlHQGtGbQGLvD3hGMBJu
mYROflxcriPB8jWLvYy3nFGh2ZUCNMPPrHkgnMwYlCs6MrdlKi6kCNMdTlPY8NgcHTdRd+fwwQQD
Uv5cZW45/QcW3iO6SZ09Lyuskwdkn7bEjlAmUm/5QD2uEEyDZ/337mVh+L4iJm2qKOsXDe5/T5DZ
kten3nJfLNeZdc7JOwSP8CI9cmbsd0w33EsiKbbYLb+YgOW5BFX5KmugyUv5q84I97s8nfepbUCU
kH9i7qipQm6D4UeiJ5bDJFLB07vE5arbQGdKT6TmPHloApbq6jyzM2CtbbqRTPV77BB+cNqrYOJv
ToeYqhIMK0SGJ09z0ywSDy67tPnJ0w+MxqyhLIVjrvA9DTGMDv+rceVw+DlcEZ+QQfOfyULIDFAE
8CC4ADNHR8tRwl4BGEJPY9hA4Q4qZnY3zrSBidBzagvcQrIOb3V/vaRy9N+KbicS20YuuyTy69Oi
xWKIhYwBSL5TiUXbbcDKvBqjWtJ1WYNJdM7flc/6KxlCxaoFN4HhJyCiczDWgaYPNzLP2/56k+Ph
106V14EKgAoNLkaW6bX750SmFwtpSmXd1vgm4xa7Lmvmjqa3HpcukJa9mcBsL49YKHCpex2iz9rU
Q3TNd4NAyPgmVKs/Bz2x5o6YpLFS87eb/j2lRs3P04vMabtiMU22owjw9W67w5IFEc8W3R0oOFEI
QFtKz3FKwu2N9yLOUfGPSMxJ0UNKJkwfqMedVv6WrHI4oMKEwsKvLeEL+2YNCkzt0+s+/8FtMFi3
M/RuavdrP2Uudk658z/QMUjcsyH6xvtLut92F5SbYQiL6i6NxddDJTViFB31aY5J9ie7SWcAa38o
H60Bz1mU8HQ9dYMKthAVfOA3XqLjQKqNU9zS1wKwJEAxKSCbsJZfXsWJ/oDnvMTs8cs8F0RrQQ/Z
+vZ2poieMRiWFyLtQCGY+meABM082amNAnm8Kq6Xzl7bCgAkkeELRHvaBO/ftIB0xn+kt3ou/kiU
4OIM3Yqdl69CvtjXVTUJyGr4Ruh+iF6kBNQgp9FRrrChnpXdB5gvtlfGyvVNgynxAp0nyNVD7UXc
RwLp6K6l8OjlfPnxBdzeulC2886fa+XyjeomSJmp6DEpVzwZ806t99e1GRs0eUx4kFMhoAF9YSx/
D9eZhEC41160pg+/KZBKv/qS+SHnbRWwtnraB47BE1YypWglLUDm+RQ6Dvt59XlNjtIVYQ7Ywnjr
HXyq4nAXBaIYGYOOOh6AkDJ0uesNbpEYSJCOtBVRmeSmMsNA+DJ2oa2N4m+bY61i0ohsgd4SFaXl
8ypCdxueTw0198S4AffHkNQuQRyLUXdtZNzrQadeWUVV1S8Q22kDWd02lDApkCNYi3pnWbYadObB
g3duICVU8iTHFTDeFy99nIXeLu3vnoORwtYf+ZlAwplMS0S126p1DUP4sZ9r99yMHw7EAGXPvB/W
0W9YoB40IHu2z7NZtSzgsl/Fu0ETCP16ZxGWm21mBgiIYbieAIhBDUPSZ3cie+2+oTHVhlkz9P/e
pYTE7L+B6rzbpZkWRgWZKz8TpmE7W6BJHrc60rRD8TMbyS2ighy1HhFYkOq7Py7/MMmSkWM2db1P
QPIgJd0+glBkGXDxFEnDvDts12AWtlmsiMGhzOC0K7Ro+2H+bfSFjPwFf/wlTezqggNow0Iylvp9
NO4P3K753BzRN+YMAyw9tNPkR2VJl44cMa8VhiYv2GpjvYd5TnowCilaHO9U/nNvxoSxm89IA3TT
LwVq7Rzx+Wx0KnlpYOsuPlY6q1pdcWru+UtRscR+V4jk/MjKbim71M3jQGC9kA3ecxHtVoKDkepS
J2fCZHiNsGVoeu9KeZFxVyu8hRThEHY4xz8ooXYNx+bhEHm2INRCR9VoaOLYmVJr3uyg66RxfMl5
09dUG0m0+kL6WhCs3z59kRU9OOH3ehQ155ffq9MJIAms8xPg3SHGoJNN0UT1g7mzhImU1OzXsUGk
X9OjtnNr5CBWlYOHCNz6TPF/cKzOgxFy7OCWIjVfrKc2micZ3b6m38rAsmP3vhdlgkerlL58FDHW
jbodEl6S3z1n5WBezINO3u8S6KeZvdPXGUE6MpXWn3qt8aNBTUL41cP/9Q2drgCW83qNZPTHAgHC
TA7u4kT0JupnYNY3rqlyXzwR+G3CtoaxM53NGq7epCDjjgVvhgJ9yMPoVZZ0iOm9BiQEVeG4/3p+
0ApEOnC9lIVCFxfZFf6jZfXLCyj7CcgJb0cbE70NOYSRgbr2bf1kGaduRT5ok2ef1Uy7NEp4Ca/L
5CK4p4JMQDYIcaXWjBUDfmdH5qs9yKbaSVfYhpb+A2YJamEw891lrX8nhv2cVRMDGU0IiRaxkUgy
JYehY9h4f0S3IhecDshRxJi8Z5N98qC7cc5IyUj/wGZhURcBzGmaOmOOk9i0e7EhTNmsOPhqyuAt
WqYmiKgchDahs3ex4QpDTkEC7367n+TFWZQQgqss6d2olLfAxepGPXRPkNDmASjEP9aOgrPhZI5n
32hVSga2/JcaB5e8+YJ12TQ188C6D2IMOIDR0Htq+HfBCz/R7xCWM8Cueqp8ixvw4Cz5PM8ALMKR
eUtPoX5z3mHXobxtisDgJ3i/e8HEoo/Cxcj9rQanhQ32/ZLUCziMfr6wPN6ZMp2pGtQ/RmytDkW1
2UDpGxnR17x0WssMnPiUzHisNU6yOFBrfpCRKHmojXjAX0G57lEVq8eOmT/c28QieXwRvHM79Ty2
0ACjSjfv6+aEVK22FVURbYlgDiuOvNkrlw7r9brWarCwL1Gd7xLxFok4Rq0iM2EvdRaHgVhY7zDk
uJ8nQYONAwWjHJuXs+It8vWX06iyR25sW78Iin2QREZuCvD6fOioEiNv2pAphAtnMnZ6OzaRdyNz
3JQkAIMtHef5CSoZ5riVA+CA+4Cs3Wt54N5iHybMm2SXS/YDZy8EGjDBXbXmjPqf2/gCuG8+anXj
Ub4Wbdu/uzpfU1sn7gzRm7Z4yWXzrti9ILpjZQA9D36n9giW2Q3dGChpV7bUkB3/mg+GY0xKdylB
OMSyMIELlzLnep1qfn28ZtzcyuYFSAJcy0o8hEV1FwNdOJ92TfO/0mDX8Kr7cJocNPidITtx69j7
UdarpQkBGm2TO7OsqwugGN/mSHjbJGR7rJmSHf+NM1aKtmIdvZTsRHXVZtHHrpk+172ClIqjDllG
oBuQQX6q5IHiNSzsl2WSOEXrkV+UXVXTT7CD96h61XrLX7hpcGK1L3grL8X//5hBExLH0yCr+1Wk
TANWUV4CkXqlc2UxJEH5ih677RrZBS5hh4YseZpSD4NYJvXuQF3Ad/oaiGh12QYADLujfNMbqKap
p9E8nuY5SZPPpAHa6qHjabb+AwyWoGq5+Yvdf9kQpYkziPjAsbx9G/K1uRfMEQCduD5jzpdTkTqz
vV60rqqAl5cv/vZ+yjdsVulopk/yHD95QYQ+pgYMhaKTKfSud7UEmL8txR0fQwJckEaiRh+ELvZZ
7TzPiGBTQ9wn8BKDo/+aPp5pBIdP3z9/tbxWiR6pUusdOypHzQ1MlNLbi1f7tGnwAQ+mAz3o2aoo
rNTzIMcl/tGyPPdrjb8AlleQntsqdB5/BtrAbXqQEweBKSWAjz6JpBB+sxKbC8x3OLYdKLbqFwYI
p+OR43IdfvfE0VfrrHVwS9Ya4WiFmY6ffEXgAjGgEI4U6k8MdMlIe4YgpAw47TG4/d4gzUN2kkoY
ALvWEG+m5IW4OUHoriH44aMWY+9M0BM1jtD4rZgshjKT31dqjEf8cs6I41GYng3hehWxkSeD8SPS
gU68zz1efKSzIfR2re11OCqJ+/eFHdL7y3Aob+eb2d57MoMzGE/2s5P08Jojx5Ppa3AttIDSz6do
1E2W2GyRazfbANFynFJyPuYfpBSucMGoq2V8hkF1EZBDuYC6uXXHdJ89tGKTcpIE5UohC2jIBBVe
dCc+QWaMgI5i31Bh4ippRqrXx4i3vqCmEO7/lMy48vjqNl70E/Hvr8KpvYADMj+XOP94hhPtdEQZ
ACyi0hBS6FYyhyCU7D9F7SoID5RAof3X/6sqRtcHG5oR7KHfxUAOvKJuVZqgkHubNQKSvFl+oT40
OnfAp/6TVdUFL4QZWlowmawXBWw/dU4oMOh+0geGgviEn7bNF6yjkXKVDFeIoLBvd8r2Vzz7fbeY
dtCMA1rcfuMuqIjPgDUWlYu554xDu7Ub9F2mQZfS7JJ/oZw/kSomdHYSzIuS/BU91kYEOrjqkjKg
ZtvNFmLXTj8K2afU2gkrZKbIV61rKEGWNrgltsF3lDGmn0i+Uh37SXADPgDQK7gJIQFbOWB9mFgT
FY74GEdRwuDbvFbY/+PSfDiUWT+nG1pqRD3o66WhNHkTRIrIt/M/gDpIXZmUbW7uOWuKbyrj2IOH
f2lD37R+26JAqiQ/L7BXyCgBz39k3n/G6fFYJ+r0Yb3nepOITpYZ1+hliWdfq2AmFfyzUvLbGhAQ
fTSUkYcXsdHZuGr6nOmTnN2LFqf6IRsf3Sp3qz7yJZdlLFBLdfUSnVhcRA/qEevqY64sAf1hPlJ9
YUp9fyOuqizPiy5uvQKdOoVJH5oNzCX2JyvLDD4D6WIbFY7miWQ1WiBUXOndLSRyi25h2f+rmSE6
oe742ydK4pUR6w0uswXrX5fBGQZ0kgXOZDOjn2FPZXyRVdyXVG7J68PctKIdq6wZM0T89jOLLzRc
Kp9KXuG4DmfG5KELFw8g0aiJNuTp/rD5ctWONzPnhvJA/AA33O7AlJoOh2kf4tEkNNF/+B8+WDV0
7Jf1eBNS+XMvwyhFMpfhzV8fptcnnAj2aFc80we0rlFdMHDAqr5OpiVN7G7V8DnN+RA5g0xyR1QU
l/7gdJFICSC4QSRy4pGpkPMgAfrAI3m8pnMGyjUtq+vNomD+1L3WjBgfnmRIpYKT+nsVW/fHEQ9F
sgDMdw1tQil0iEQLCp/jMoKxewpjz6nIsm/Vc9+aWFqCCdFdEOoFBXHZqAnTdEDT40sIOLzBiTUm
rjBDBOKjpeCYpKJSBgLpYNyRlCAK3GaH93LSLh1rmyRk9CRdk3dMoJj4AoWuFGbZHlb37kovIk4p
775KU0lHFuGYy+2F4ZXFgD6JQp8W5eEAmRZVWLyhpioXe3MuxJNAOW8enL5+XWpI2oZ1mG8HsU6+
1CVJDIis5fNXC84x8Jo4QcztD7paRrjS0h9o+huncgLEeGS0A3MB39SbmU+XmQlnKEhtL4bJWJVE
xoBd3r7y/Qnf61LKlxcPwkrKwSKEbEdeg9QhPzY40pgWpIs/jwUSIGF5fxYVxWM/4TeyyXk7C1b8
r3Oco75gGtDkfiAaqpl3khiyw3yfk90ZSwpTFP6OFKCv0FsYmCiod9L8JnJVkK4qIsN0LH3i33ny
MFX9pygzFt1IAaduarF+AM3yptEI6kNLcvSu5UHC5f2F31IyV/KTkrnd8h955zc5n6JW8p5h8ISU
d17zanGBAFrCYcJLUpNLUxSyd0Ah4MON390hKr6jwY7KMa2O2Hh3Fi6S94pDw9zvTSxXbypa08jK
JYUD0Y590dWHpb4PKhUFu3rgpbr8QHPsdo1J9vVnvbF3abwjN9jqcJ1qD2PRgz2uY31IIi+Jgk++
dYrsVgt/LxO4mwPVYD9GOM/1kn+wIyH1JjUSEy4U9LkCEoDLkSZlS1+yBleLwFgf2ULPXgYRKBsh
sDK+r1fw3rnpGRLJ+3gW/A7nQMy8kZuRogcQuOxcdIzMJRrzm1Y0cLhfA+HRYIN2x5wnRagdYKip
9xE3NAyKA8ubsIlqmUqLDZewZaLtnpFKHAlp87pkVttE22feLuGk+OdlGSxY5E8jh552Q0zpOMc8
Z4XkdzonnTA3HW3cNVGhryri9QK9tueDTsiRZ4myCDG879BB/7elE0KVCL9W7HgpnsNcKT9r4T8y
uDO7SMVhrkNYBTxy1Xa8OPE3TYEjhQOi6zGhbcgPQW3pTi127OPArYaMzgZvTBQMxvzePxMCywX2
WIGc9h/1DSa9tYw5+Exnn6PEo3SuLhq2IyuG21JdW6Ae174HHY8XO9tb9g8vb7lBgzmLZZoHN9r1
nkEvMyQu85HGGjpoSosl9vF171HysMaHCXY/BpFf7X0knJnykL+zE1+7TTUuyzWCQ4dn0fqX2AFR
ydFowBQdgGMKNfgR4l68C2VD8REqh+YuY/X1H6bdum6ovo2OW8TCi04cdTZZc9PKuAU7fyarwdff
Y0M0mQZMfI2VVw5fXBRWlSLUnMNEtewvChAYBCQiTBFxBHIUGLQthfDXjY8HpHC1ZzZz42ALTsMe
KV4lFVG/5FTffnkwJZM+9gQlaN+IYBgASezKTPs+QP6GAFZL4eI0+MqdAq8TigpE3GOY0DazqcL0
qISxZP57SGO008IfDmFKUwcMAyDDXAxtRbChFGazm+p9i/PjhqWO5piFnj/P6GFTKWInDx1y/vYZ
UDVulwUuA3MwtHsQcIKXUmDfbSx5aOFRWa3BPt21WnyFmApiAYWuC7kJN8O8qlfZRWI+ww88SCjE
E9nWCdcmJ0H1sL29cVQuDOaLhct7gIw0Ed3Ih6xsjIOv4CH8uU2OmT0589Uzqe9TQJ4b9twnftjQ
IJL84wgQ/GK26O7MP0k7aY0u2hOV+4UYNw0C98jaSA30NGhhZcoGW9ElPKj4Uo4aKg3iT8Fn8KBo
hmSjk/n75W2tD6Mt4/4WxUTUTp3Wm33PpU6b8NK1zeVeoCYRzDEuNkOpNOWnNnR2QIztNgcQbige
a729sFws1mFEOC+pSBCQA1SR0TrSZCCmrkBhAhmJ0wbLTawnVYGRmVfW0o59GMvG5WKN67uxwaXa
SsvOZ8Dy32tnd7kAE3hBQyDV/4ojBvboPa/3AghHWAnpuTfzYT/kqM30eQbvu61zYX826i36MDt0
uVYIAJ8Cjs+QFqqL5JTALhAgA3xdh4paCFdNClelvWnmgUS71WX4ug712HSd0s2aP6s7mayDVpOU
HV3d2LoiEqtzqdCLvPKcLw6YwryROi/PYQnQ+ljaiyPn5zZ3XCbfhzQg/JITxmUC0X9dn4UfM3R+
Iy02zSRhay6EPrCMS5RNmJBaoCnmIX58kbWBHJgvCGf6Gy8pk9RHcxglByDWf6Zlos4o8NPw33wj
LP/CadIdJazkPPj/a2rwKZHxzZvYUvYM5TMxZ+huIvjnpnGdgO0fl2Nu1mSDEhbR+CUTJCmmNHXI
HMOTLa6CrqSEGOxjjTso1550z1aSQtegj47SFj9dGnUIzmWvO4I4FTUnJOy5GrL+xDDBEYjk+MWT
hmZgkzAPV3QeFVEKzD1J/ysJ7M7mrLTPgFA3qKB61IcX2gd/LE/Kxv9RAfEu7IO8QZUspA5DwbyH
k09xhM1mYwdlfodMTWfwU8OJcD6+10KwOYBr11/KJMnOY/w8bAKfoZdeBHBsaWrvdF2Vd/9D6lWF
ugUFQ24qdvHriCY8DQWqvlWaUaXPW5x9SGS56TqfUJb8qWPOXvDLofHCIQEwR13I56RQMv3E++mr
7xXtbms1UFfVCzD5FdCgLLzP+URGPDILT1HdvywK8IWzJ5Wg5Sxk4/RF8g08oE6dlFGcMlteJP0W
sMXS/yu2gDdE8VVK9tW88/SDgjRyT6/V4n4rpxz50OnkWrV1oH9JK7IasZH5+B7Y7ZTeD4FxPfOx
0fuTcWt8sVBiphI5DcloefTDiFK4FuNDRRgo96QLb04eReH/lWjRcMi6hVYzJtb1pysNar/pmCKZ
lOvF0iLDso93HJX4TeL4TymsjsamklWOBY5Fd9FT45jjz1H+du/phJePSZdV6RDIgl6qtDcXR2Io
dGJ4YiAgPevcIqrdumua0W3eYKr94zJ8IQv/gl+M1J+MZbCMX9NTuNP2Y6XtjU/z/3e+7OjbFCgy
6jTzxbIPa6QJomL2g0d5rl3P+LCitqqb3kZI0mNrOa3KsEE5LEWAozzNvHYkIPPHC3sVs26oURfG
Cqaf3wcmtHzFEcSYlJwL7lWbu40CaeXHJiqlqNTGQ6tWv9E/IeVds60Ch7q63nftKnhIHO94qcHs
Hd/tu9GMDoqYHp7U7HjLvuaXyMvQQnwHefIxCpFvkLMuv5sp42fw/vi5OVluB5MxEJoJuI5ejtgK
mj1QHwvNXcTyVNhbJcp39vmjTIdur4xCCUXh6mC6nEryi9GEqIcXKDPWF3STrmX/Ru4Ar2VqszXb
gunElRh++9al2cmPW2POWHyXwsSn2eAWLzkoXHEQ14bvQXfIUpY8YpFBtphDOK6zEPxH874wl/eY
fvnik94IOZ4UreYIQEso5iQiurgo161thM8Nw9Me32CIRMhyNM7evmfcwg6zfkk/JL+9aweJHySZ
ZpVeLlz4oo15L66uE1l06+NSQPJJLlBoef8c4CVADwvQxvdAdtTWZU82kNI7ynOEMemBxwsk3dzQ
HILiWcAX3zOLKj4ZBjUORMEkL0NcaxuKHZ4GySOG13YfEjiEIYwYBF/Q+gpVuYFiaZPk1Mk4lVRX
00L5MM+CK8NWQJ8rfLHQ8iqNQr8699m1PW+snuXwCu02CoWjgvT16Vlj6c4C+j3gAM5JfAWvER5Y
MdYqxISDyAYHYaHPxeVGyK2usNIu7hZR6qsgyqW7R07mCXVyiYnnmfjY17IGc92hDfsUw3HDbyYL
QDRKIwzalSuZs92gZ/1gjTwMiKl68Xi3HCXfsa9OcIzoovAFiOfZee41d6Dzq4At2i+vvFRAQKN3
/jBAQoaj1dCIbZoM4z0zBQOMJn5DszyuVcu9Bp1PN6r/ncu4lZipjXQQPFD3mOZNGPiPtFJ+l/+9
QB1MdUGjZcKlhrFKPCXD3f9xKMIt0/Sa/1UvadmIh9brTKmuvtU4QO2v1m3f7IgIe4M80bjrwY0m
GUH5NYrjx0ZqdJVgxpND9x9CFN4He4blM7zrcW1SqmWJ3TK2NI6z7m5GOAssVKZqnqSCMFFy6IrA
X6bpJvgGy/aIAHe43xH5AcLJrAgmh0oBeJQphQwB3Ar6Hjq2kqACLOk5L6lYYFau8eoXpTGmBqlQ
9Qfngme4RmYq92nyCwKvdjy5fkorMUGqDytbTID5yGxuBRys3nXuaJ9AbnIrp0WV8ox9G3dK1B7L
rEIQjNGNf79AjgqrSd81HKner4Oqpr0zbgNAO2xqeF73MEVofyE7XAOwhkzicUX4MU3U7M3Y4MFT
KlkSArUiRrqUSafnqEEC+f0yD2USRp3ktQwulMZ/k7vUQC4rCyDN7ENIOnftZrDZvP0FKg0NzAv5
U5Btsj6h514Pq9v6MuLsgRljLMeF2SygUAQd+6L9j0w/jd40n+PrOEemUEFHuKIvMs0fd0H6MBGn
/qf2ZbKHnds742BSP6+hpjMIH5+kj7n61je62hrnQZJflLTr3IXbDXXDRGvcnoBOtr5yNeWc7kfW
bTYLOCTBPS//m1D3focMNPkT//bFvwE1ZsMkToTHHk8XraBb2wNUPep/qeWsFiakhWtZB1P5BuKr
u9WrzkxGncL8I/tHpFBVKLwe4zur8taOm7hP0hgfGyigW0tFocE3NP6asusviNwLFjbWFBNZQMwm
u5E0WrvGVEn1KWh7UetyhuQNzaxyy2zCBO5tZ7t+xIhdTfp5Ew8hAlegKQf/Gh5kRrfG6VKLTcuO
r1439xePUeIoHUsqIs6spBcEvMOLKOZYTPQMUd9y3y+rhrK9RZf+15uKFV6JilOSDxwCNoNxfkUg
dPTd/+g4DEJAf/NBkLLE2d0ez+ujTYv1+hK9QGLxFXaM49mpXk/nkFPkXAWPaNU+NtwzpClqx/Kj
ZmfsThmB0aEFzQiw2bAIl8zCwgqrFlN1JGsxoDIH9F8SJlBHe4sVsnhJRRrAX7Q5li8SCygEwY64
/f8mWQBCFzighAWIPLTbMu+04+uMLvGg6sy7+aT5saUSMyQWWgx0LKJaPWozASydCz8ZKyutavsG
8Crw1quzPK4hYQcqPU3lGr9RutjI81wIqVDH2MRP5490yT7X/6pm0rxz2VUT4AmNtY175a+9cIa0
ukXJjR6p90g/vErkZ01EjqhdrlYYLBc5LgqqjU4B1OgbUdMCr8SkLjM6iqN3BerA19g3s2ZicIpS
7bqa4mbykBP270x519OfITb82hzs2VfCMFMzofLroygd8YaTVLygOYA9ggx6qIao14mO0eO7Rt1S
AjMmb0dWQRLqO6YJvv9vHUJXq343eQkTPNnVh9u7J6RvtlGmM7xahyQW451a6kfQXXvS1Wt+ql+H
5MNd4yatHj1gflxvi3qLt7tGAShjtk02VMXWChv1xE32Tro6833imVvOsBTDxuCgxSkVl1aFL1va
4QVmUX/C5TZcsgOZ/sD5p8iwN/TQZ10Tq/wRQNSVHF9b2GwWllNgM0jHyWfk6x3kWviB4y8DD+II
fIgSwSmea1gKk1zGTdZZ/4FVO2zS+u3EpPRTeMiQB/PkBglYeMVEP2Kp7htKHMZ9a9N4bsacRWBU
1sqblqbPlQr4auRaskzzylw0zdniGEXBdZRgkUwLGCWRVrxY2eW+q53LDdwG1ODl+jGmmP3JRi9B
C/UxuKD0z5I0Sd+QsyH68Ca4Tig4jYbMaB3ew/oH59uGmxG040cad/qLlIueOYt65RUkHoE1ZsZ9
Z/5srpnhzND496onawR3mdK1mS1C6j+nWc9iVNG5SWe3dFWIzD4YDB4/TKKeCAdg1v9tlzvCHXeI
hsAy/5LMiEmqlDSDuJYcfJNTUZkSrV7kgWD46Jc3PaoW/HbnOgBpHXERADuBc9k7fu7J9X36ecKP
llKBxXGgbX/+/EwBc2Buoe2B9ZPAY8lB0nM0VENj7MREogHHSdjjIr4vaOqxW1HymtPY/n0BAavU
cwZZGyndbCCS8sJo6wc10QA9ok44p82AJ23hV6OavZWrvvsinw6X04QFaudvZ+pT3LJa6XflpMPQ
RaDuhe+1qB1ROMEkczEgh+tx0/AzXlHNhLc8M8gBZ9dXHqIpVSotpVWJdjW61ex3Aejvemq80Qcp
Gi8GSW60pCHTau35EuUK4nNAWQl0bKvLI6kzEM3sNO4ht8XXTCAvmFGn0lerftyj5tIVAXPZQ2h6
OXKO+pB658A9N/j+RDsWN0EUcU1Y3p1QxGO9xkawz8EsBmwCCrU45IrwcbUEWx3wZ/EGiZcTYEVQ
V+2uUy+81of4Ii0YoHH0R/XDyWXhDxM0hGJUwI7cag8MY9Lvy+n4iFV95Rt/dTcTj7s8i+cMP8pa
wMCFnSRmqw34kgEPS2l3HxLWQ3U7f95491WulRIY0OTT5vWcsOGopcJpDwH8eO2IKDg5etNKacYd
WUsgSd/PnNVsK8g+bMSmgpD8/6ySGNe5NicHUBtSyhhDg8QjVFYs/xmBxr05JJXTg8lZR6QFDY/j
Xc0edTURI5ITaqFc4kkyY1nMjWvNZLEGtxtH53c8nJnCpBwlw+E7iBtdHoQE1C9LREFjqj4Jwsv6
htE+EjNNDCfYjhS7iqKQ8LuP9ahjfpnU1Q4LziKZQvH1TQFrqy1VFRSV56MQs97VxB6teo013zkb
IIaDrSEZgwmEUq8SnWIFAIAFzh/3wQwr0PJzQNvot42NVrlFCpaWBcfYCuk9nMyznXDyBd4HNx16
ieHLfdVRdKWBCLzCxA3jY6+/m/yPclWTsi0W52WSVnmWICHvelFXdPsN8ktO1cEPo/yR0ZQhaw2B
wlzC2UERE80l+2gdqzDTZe2x9OXvdHS8ipKMVQTuXhr55RF9UabNG9OLDE/gNB7Indu9XWsNqstk
ZInSiFwaH7uKcvtRVMGzEZ6mV3bs4TtACVd4qfJl9JueIOwh3TfVQtxwhNycW0tjLnr+IH64DKP8
iqEF4lOHSQt/0K+vdsDfbFNhS7EJhXQoJOIO+bCr7v/5iU7PzzsG2HE+QSb9O1NWs/FvqwmMoGUd
qBre11J/mzS89ZYPu3JZj3gQPCtUJBUL7tEjZ3oTx4OH+7W34sI6AeMgTROHDe/UHOo0hYBHRaXD
hlGzCRhNab4HM3whJLu7Fv0cxGUO1O51wzaBMfz0wI7y/cU3KMHnb5Jd2l6kQw/CJ82TwcgjDrTu
dqvYQQYRhmLS5wZxuDpyFdlxEzlFgspH2v0eIrj8HdWN9Iibn1HI3oAFgpywZl8eRyG0otLUlU6c
+9fIkrfANpBAe1pwJwTTV45DOn5vO+t/F+ynB+oEgTIznuO8EVx9Tf8SvjCnwrqamy9EFvOwlmEK
jQ95MlKdShu10jfTlqCaAZldhnaRgz+iRrZs99OUhcWbQ/gxK/EtX8+HumMnuk6wEcg0+9U+gycj
ayYMLI4S9n03GSQ/0XFXx92FLX4CeQvG0T2FUw9u0l0ycL03Hk3ThcOIi6F0b+rYaF3D2tgDLp4d
fC1A/Ochb9kfVisgR9DeRyJGa7/kVPqziT41ZjIUwSM7nu3xr8M2vFFHpqDSzqcm3c+QyoWgU33g
dnMuAV9BXxVPc3bHwpfJRJinRt4HnxmahbbqHHkob/NwdC/xMbjZoLdo3K/wa0Y2qTdF0RGsHoUY
bJTpr81Ky9IFr6vwdtAZVtwz7rmFUuOd9RrXbC4/+7aKIqEQHzUjmk+K5EWoqTkqTbw66iqiRHs7
rfD8n36yRdl3Jt0UGRkorUnsbYuFK2HLP3oCusalJN2zjqF4WIK5iGEJZD9klnhORfpl9eY8gQdk
V4022Osx4ZRYiU2rAoMrDMZllktR2pUMoq/9lKdj9pM5JteE+8suwohMCfWtChHG3rMW1DgYnix1
GWZ/ojgRE3ceIcRv/gwLU6/BgZ+7uLV3d6Rg1xLdc9OMtvnJ5uemNCEldZPopRV3dOdhrOCH4NKI
sV99fjMxadxgl2QjzS/TAUWlYH8A3/+/wLGZUF+zmzjwf66bUQo7Vt1nSa9ggsXDUnxchIm/KYWf
1vv9LE909bLTHdUT0+iEQeeSXaOwn2gRaLy6qyy/GH4sxJVUAQNyi/nG51oti6HG3N+CPTPSX0sa
or0jlB0FRlhf7pBwNSGhZEJk62LGlhSvm4iJjyBPkoPaaGc2daMgxJ8TdCRdsSgzL369R+RoILZZ
nUeCSJOsdI3dYp3sR59t55zaTQkH0DlRzRdv/uinZr2DVTV1bpml93XSTXgAGhFqtWvNQ5LrpWJU
VX2gm58EWnnJceBY4oZXdr4aIHr880BNJ5FTlCrj1I5HWSvuxa+Az/R4iQVghh74yn+okIHZFgl8
PBqG5xeN9mMP4x0ZArLw0h/svoRLD2R9hC/EO99bpbyJ3g6ygJXFxFzATeJyfsLvg2pweG+wc0tu
iMaG8VqgVwznJqNMhe1MdYN5y7zr8S+TEbyh8jAbH2dUUBhUIOPCYWCN3NMHYPI9okKSAdSCzicb
u1sL4CwDUnnzrEfSHKN8dXizcsJ4w56l+EJiu4EbjiAWI4snX0ydj1NnOXp6pRfD/GSP0vrH2iv3
9MdT3l4rNd+9ITcxA7Mxf6DIyBQD9/oCAip/6Pzi5ktnSE5YTuOQkgD7Adqfs7DkSatJPlLhKM2Q
D9J1XkL93J9SYawlr4rcCrDKt/XjedqNOnfqFirxBnsdnC5BhAHYRmLNr04OS38krWbwiB9m/m9X
Km0vXqBBQWeNWOj9RfrBM9scfPeTRuCdd1WPO0PtTW2bUqJfXaaODfToOTr91KDNF9ZezMNDOHQk
tJNjE2Z9CR61ygomT4U1vhftjehsloPkXGcb7Mrw66k1/DrIUc/yPXKn3kXUArG8FPUwPMqJpve8
9blmgSQQmVyDpcGmClE/P5n0O0mFCaZF8SHtZvnO/RihJt6NqcgfNAus/Pn/y6EddE5o6ZRhccy/
OWHOWQt8wg+NW7PUY8gC5/u2szqJkbnnmFDGKAQD50Y8dDyhhf4NWEsM5X/y3qKjNdfYs/FzuvDD
IGId52hSLEBWsoA6A0xjdGlVqc/tIt4V6aCUQCFYDqWbF7Xo6zGZUtpXMS7bkFvRCJEqnQqK7Ksd
wv+ocIph5jMSDlsgJA8mICTG0IwnvYunW1A5l9QnKKtv8RnGixNLI4zP/1UmmF1DQSuRbNobOAmG
N3ck0OiumCSvIWSBsrRSBovJuiY8Xmdbpzci2G6iL2B8tUolRP8x4cpPDjns/WiDbL7Tl8GIbtga
iVkWYzYnUCd/gBiCiFqoY2gXjoeIG9SY/9XQGJ6YnPT0Y5kSgJfBudOZFZVweYDltpQAyIbhtWTK
wViBT+KWkq9wfdCvErd+PNClSSDOW1G+IMlva7shbUFmBinsEViDU3frT5rTlUq0vswypNViZlPr
qczswcZE8hrgimK+qVFsclp6rHa/MMv+brFaoBqu8QoFXuBEYlMcdbPByXRevinu7ZEfmucmRT01
+PRDSxmrL9Fw6GuHO4JznkF5xsBxN+HXzvP/UIgzCPltOWu1tC1lowvqevzkZwXlxwXZfcI/Xmik
2zePRNFqWBfrY8dP0pnt654vXb8cx8UNxj8aElZ39TyEZdxui7JcM/XRu/Zs9zuv9v+NwiYVZ/Z0
KZjrCkLTELKwG79TeDGnS7p4ViFXDf575wFCtcLjDDItvhLCsug08TdqGrW3Nrlq6Fm/TVkdCB/k
ngWN/v87z6gp7l2XzTtxOSzsbkBYi9vLQqfNsJKQtUlVAOQg1kbr6UWjWiBfh25X4+j0iGkwjCGg
kNSfG6qPg8onuXlxdEze6auVwYUrqbnm+8g4CT7amQ34bSkmpIwAVOR5ML4uGPCQQ5lS61c9CGvW
6nLcIIaxeDFvBQA9thi8eJqmPizrDD62l+jd+TA+gp/eG/dZdeKzTWLH9mbK1Rz57VDH/yqEVrx8
rj/cMNm0gMP/JP2mJCASKQWamfsovit1poHV45+RMX3pDQUHnnuJEy26fLIPGiJLosWQeGES35OR
W9jTp5T/ksz3sHMcz3TbxdRJEE5k5fcDg4y8GdflwSaL0o0qcubDohdNebIqPmGZsNYAnS4oFB4p
/MTlxQKtiDYb2ur6x9QWRmrEC2X8ESsQaTXWw7I/8LY8HeQFrtr/p9eJjpsdX4fqFHIjBVlZk2PS
LmTdIR+4armWRbF9Uqi8Givq7TTB4gA6Vnqo8l+RiZS2F7a0F173fWTXC510ghaCKQ+m3+cJQnRz
DvvYFcQfQC3bkcPyIjjvOIJIXuEYOBxdXVx5+Hdi9SdOFIb8zSA63xBFvTPrl16emCuqhr/BwNeQ
ckugSk6/I7OsbyHpwzcdYOnBG7QDzDnsuMh2kIjjsnp9Tv5ib9EEFzExGXrJ/6HfQEFB5x6BPx0k
o1bN8w59VnPdc21lCLwBL2KYs65nhZtkMMWNHGAqKZflpnr2gIYnKtWYEmnaU6AUftKIOgDa5A2d
K1OS09GN16wEfNjGcw0rBGy8k0VPd3rV8Wr9pYXI0uy34yVnDk8DuBjJj8SWBEPU99mARjLA7Cpe
AcPRWFTBjpfO55+y+yJeegv2zzWe4OSgB7wEC3RwZHei8pEztGsfn0olkHX6FjDiDljOByTjYRwK
idlWtqGasCQmABDr9/pVwy5m662upK7L88HlsTmn4YvjGOWMWelQwxS5r+ntqcKeV75isaNbvHk/
eMMxXkPY/R5N44jDTC35ZyqIEhEselRd3F6w/j8bHpxZsuWcT0D6La2QxuWeCKvbUP4EIdRigW/+
rHNb3gb0jzORjUJEPzql/L0q8JjS/EAVyVtFICBDa5k/QBtZbgBFVOYXAhPsXaInkBrjfUdfpFvU
TrRM6ZR/HSSIa+ekwjcTn1snDTZf1ehuVI9Wp5K42/r/6Q25gtriV5lL6VUaa68t9qFM8iN4tERC
aJ0z55X1ApxlY6EYGOzNU0eEnU3q3WYW3hwL/5HLroiiN4MfreA1BqYw3Muc8SuAB72e0TzTXcfq
Qw+nrZNiDiOKqjflOg2Ec4TF7qNsIC0f+7Ay75AGYwi7yQZTNXoBziDiWvSoKcyTM/4csu0Vt1g9
ZSnrEncFNhFFNowFtHSlQnCv8XuL70wBkNx8APx0nj2JCdDCa/DEjmuaDDfrcYKLIbWokuDLDq3p
OdLa/JuwEWDTlDH+74pqZWcZkl8oxZHzY0XkCl+B+TBtJCPIz4brN00Z1OA2zrFBG0PcnnFBIRHC
Ezq4lpjzE6wCePrYhkG4EX8a3tVQRqOFfFwFW37MlB26/9e3eKD0HXGoNsD33+Au/8DcTTBo2BJr
9/A7Yz4VlEKkdic5blSFQd84kKKvy0UGS4/bIzq8KHC4CIcwzffE8wiaJ43EwXSwO3Qb8sBKhyNl
zqS0HjkCgM0GsqkNO/FMj8f7lXFYqs7GBB/JtT4afp760qTB3Oal4vYV9tjEGd5Uf52JlIi5lOh/
25oTdTe66M7jbcSQsJL0Ccr6+0UHlYt6RcixKz8ikHtpUWAHeQdoGuXsmDozapD6oec2LHgY1w9b
mOnboGM9E+zTixkOE7WOVwNU+R+uMCriddekg9IH2Sqy3qEC+wPJjmFCg4dRXOSs5qO2zb/qeqjV
uIKrmfkJU2aWF8SZ/xHQpq42cO799evbdLi26huOof66bCBx3vnBQmdbBEQYHW/WeXPnp1gHeBQ/
BcvtcPKvO8QLSEqc7nI/ADtVU8nWTBC6KFs9eOQhLF5vpDg0AQIr1ixdrWNXtGG+/8W7vA+Iop+C
8EfRxTZZZIzuYlNzZaZs/4N8OZwjXdQjAWq+qbc3jyJHhcUxU/LIJ9PqFIB1971gpL3vgvclOsgS
p0O3FmixxBJQFzzpiu7qQIjJ15ue3k20C49x49KbU0DH0EiCz7eVQgPWhRJiNchlbGnDRNXmEhjD
DN045T6g9X7PM9w+qG0M8PK/Gde2Q4dYGgaimBDckKuyv1ZETCyVTEyOxJ7ho+5LnugcF73avtZO
ezidbMFZt+wtPoV859QZKbJlwSGvOF8LttQJTOdJdhoRiJuMfVrOhhZYI7johgVKAsahHr1ujsp9
y4XCFiXI6xesP8k6aLBs8YdJhUULkeNZ4AYoXAe/uu0RQuYZWS3TkLaOEYR0a19n0CnAZ1va57aI
3WwZ2kURW/NVfmvxnUFnWwa+Sw4z1Od21XlUXvjPvW7A0EEL4NrkNCIjugGKGSmiji3nHSsNGKm2
MoP+9oE6Fbj9QtpYV1UELhNjHJuuHMNP1s8/OpCKfTVJiL3yZDEdnABqp0zchzH6g/Z94YBlmTUY
Ao67DORgnygPJRYi35Lm7EgoOvJWH/UWYJ52DLkLITtp9sXPY+KIV+uxPsDA4iFWjDeXk+SFdb/r
nk/wKLnM5V8PoaGZLQ6FIvLLHBerv/FbHY2kTdmjDvT8fMomaryaBqjJRrF8BfzLwpdtfjTJ7lX8
t6gLDC2GAArC4+9oDMmnNjSoJUhb5GtMVwoLtZvAiLy7o7TUKRvC3AnKAogwxskkBqchXxnNEWhU
XCIBud1j/Ag8d2uI+lYv1hKvW95WgEgQomssBp0FIrgVveat9JEd8DgL5PDSm23gQJgC88xt7Wou
x3sK21fdghGd5ZT7zZRdvnF8KAMpETKR2UyOCq2oKEFQDxdlhqRePQ9VwEjNB8XxEz4chrYTzR7x
uGt/lf7+8PsbOinKYa+oxWBCrGQT5YLBYosB1wjGXXUZM0mIbaN7ThQBgdH532sEjbyaWv8DDrtP
y+1+ynhTsv1dduep9wAFuhSQZTnMlMcZS/5QHNASEVRLR1PdZkVhCNS5T8oPQdj+FUFt09BbXAT+
sKMrafaJDPkRnE6fXwpssDK2Yi3YR32q5tKe6vY8AbuKzxA93onk7gihIIlheDhchDJcl18VhvHr
/zqnmnsdV6kGNU6WxYyyGr4Jkl0kolxz17LEAKf+lSGRSIKpISnH6gXu+Iw4sD6idRRsFJsHIy+C
C7optb0cAbehWdjSG4u0xEFgkMF02o5+vY8Au+QOhJHbvF0WYRxqbFP2yCrJzkBcyLtCcQiJe7gE
P6tANstKe2p4JtjzH7z8Gek0qiCjQxCRIZB8R9rD8zvPuyHBaA/McuIo+j3+RDNImSO+79XGVD1p
sZWwfPJGp//NsoOVjTmsMTdnFg76ilQQAjKuNB9i/FezunbaUThJgRGSacnI1IeoXcoqiyW8VKYZ
g4b0duQiqMGhdnCOjPkcGSz2ujdC3845uPQtlwm4FpELCjx+U3hiIkqgLih1nay+x6oIawdRhjxW
XSIREHeKhBhK6Zt1Z3Pcj4u1R7Ojf210luW8hfD8T1DzNW+J2qNKKp2+KtHDJn7vPUegQl93OCmn
d+1xRRVflLaHIf/yAB5y53DNwjP4dae55b8mJxB8jJIo6/p4rc5kfT6o6Mv+2cmvpsr5dAfCRCLd
0sxb3Oloof2l32x89lRiMgjPsG4aNdsbSIdPLHAm2xgToWIDFkMB660BjVyyxN+myQEHh6n4xW9/
6665IEqSGTIbk2wDzuF12PkzeROEwCVUOIscmgsYmMX8G0yS7g7UIPdqkLwDmN54OCp209x/kzUE
2B1Q1Zk2ETAr0dCsqrK+4FeeLKofdnffTPAC5BZnpOxJr5NQ85CWAGypWGF4l1quByII8Y5XNtpC
T8TcBbdhVxXG7y/EnszuRFqtSLjlIeTuXEydVl+ogY80vQVSXpRXy99l/JLUTMeAlOHnBTAa8xUh
o1lgjd7UtsZtVk21kDTYEwjUR9Eo1f+oDTBsNmbrELZQXVSjzalXdbHenMotMWw8kCCUg/oTYTaM
KmUnlkl6GDceb/D4gvm46Xee8JAgd07fsovmyVS3Ie4tnTweJAnKJe4kU1YcvydtekVJmzhss/53
/jMDcw8zkuerKTQylwGdFRuxU8Ycm+yk8IKBYK8BtnP/21rw99BgTidoAmzjMfnXtqZgukmmLIj6
KBJEaeaMCPxwth4fqnbxX2byXp72IqbPZUeCzpaZrlUddK8IBeyS7UPkweELQFHtG8ijI81ZUOEA
yLKflP2PMVptg1MieNUcgxC0ZRODT+3CVvT1YINSonlHS24T1eTrA0WepRcTkiAcnCPDvR/H5rqH
NF60NzK4tr2I5Ajw8cYQ1Vldy2INQp0YR2VJaSTQMXSNV72KZxfH08qsoTdHgj6qu9Nl5xQxFMOl
cvut22C3qyyNiZPsjvwr2F3MnbKbqwmOd7Fr+hPwYvnv4RrXmU7SaLiR/W5g21GQ2p6tYhOOl76a
ytFNhRVk/PojK2z0t6gWaEYV/+NBbPxKmqvYDly87KnNuqU6cW+KFkA1gFcWNkN62TByDHmv5OCE
Rg6pNJ5lkPwQjm7hCedll+y5rvmkKMckDu5AlNQCIzbftIHwLV98vF2UWG9huhPmWZNOdAeelEQ2
MxO4k+AOX7fKBaU4LqvbS77/A+QTWD13xTwNxc7QzfDCAwggF34YemF5VVclg2D9gd6q77lJ6Blp
njGhZD75hdCp0jx3ILv9EJTCi6aSdxnEL13l6IjCJW+oZKGzgYvU60udWFRUn/MUTHMMhH+tFXUI
YnuVXbGBLx0gBev7uEswOBI99W8cJtwP7gMDwP8Bs0Ui2Fhpes21LdAaIqBdg1PgzU5+RFuLBm8o
bCviKKHYILeX3XiDm3MhkFjl6IvwE4zCTl+B+iLiuRY7+jxfXbtOEE9h/pAfXCSU3t5S5tXio+m9
8dxw6HD0Ge3hGp+pkjH+bkF108skdYtzsDaKzJcfAEF2BOKmndtMZLy5mCCeHCiMTDE85ZXKKsYp
5rrLtpVubrm9etFii78A1i2UxfzDvJIubm0a4wWyT6nEN2xNlk867dGr7aIf65xgvlQdkzYTmYV3
/2Q/AAtu72caONStPyUI5pNWIVb5zLiQNID/GuubM+xVfxZyyhY2ld2ZNzGUOeK4xnq9i+OYstJJ
giRuit9SxGnoJEYDzX36aEgaYMPvsk3sPzlPQ6/CPRK+OtnrxbuOifv51Q8CJ91J/R5J7+Vcqpkp
jzjQ8O7hMnRmxTZS3HRiBSnxCKnEVmgsfcszJ86bgwOy/prIOObPpWm/W5ivWZHD5xyeRMIALqEf
Byxlx/X4ATAE0Hag1MCv22Ccq6bmaWIL0BsfjoTJZmJFbaT3onOEMZcjsrgSyoHLDsKySogbDoMG
74pkdX1RsyWxelBWw0dR1SB5yLtxcZRzs98Mmx8uhyG0/UGy87ha8mBYRlpuFvrWkIxoLgvb3UL6
ZIdf9PGvlXJaBNblAEBLPaWUyaAhX4y0LaKRs2Lp32VoGh2RT8y+JuhW7UIQX1nOvKoejK6M/k/P
jBmMEiaSxZmJVZXF2wqUYfaBpZU2Fu54wT1OvtSYtEPDB2MxZ4OtsXUAjd/A99ZAzU8QB6dH2UY5
fDpDEUCr6Yr47yiDA4Jizhy96wFi7fWdxmRDBUWF2OIIEOHRvH2BILC64KYBlkewdtQlBsnq6qE3
EC7dC0c3Ncmw3O0JWRs10y1bjOQQ1ub8F192WmBnhrbXc0EkaRMuFUqLXxPULl/EVlCQ4XyQrmJK
KpdkQnpWSTZUDeM11Z6+nJRuLfPvWk9mfBuwwFbbe4nfNQCICqRqDZxjvl5dDmUo+J6P+7HGfOpy
jOpd2bOBIIP0IA/jqdbqG5Ze5xIFcB/D9j34ArWcU7wX9rv3jo6uFN1h6i9Y4qTXsZWHJGxZr+ER
REozW4UYHFTAxqFsSjx2ViD38Pd4BeLPhEWx2URN7vidObfDYi17YjGhQWjctbJSfHocEC/7qf65
axymPQn5uq83ECN08NR+vcMSuvnzEjxSdmhX3NEs3rZO2vCOpgX6zw3hacGLgy6foAVUrcqigbl1
mYWeokIjDoAfk832ExNfkIH9OM1UezZbKzV6UvYAbFLhKShCncVw2MXcuc62/+bmGOcvv9ijAYY0
VmDVoBVl3L+if3RqMsYHUMzCvPKvjRvjE5JrJ25jKV0gEqfXcmJxUPaCEfkRbu5utskt6dIWENP3
EDavfFwYmxJv33NjwxyDwR1EdCWamDJ63YKFcOnSsYGSbbHc5nW89dQds7C9TyUpJQTys8Oe7YUQ
KQnXdHF+HcgDIQ3ThYIP191nAa4CgiWiy5B+3owiigHh2FXEt4IFfN1eyFfvE+uO9STgK3n6oy7j
sVUJ6dRXECl+bkfpraj4dpMETod2PT02KHbHot4nQU0ioCMu/YO+C0C/5JB9i+YtX54E3yiMyGsp
Xb2Z+rQ63Xrk6Wwk0CUCyj92HCJf/cPJ81pjpAvPfiZjRFd80eYc7h+f0NMfNHZpc68RnE5/QLET
EG3e67b/Nv4yC9/5KqFlK2AS4cG11iKM3ucmJ0BFNlu981vShRwCn27ewIn2NPz4oCJ/OslNXLYM
w9jCb24A64HTkHJQgXKEGvCM2bbIxcueau3h0ul/D6dqwDpSIzh77iYS4hDlXyHJ6zXiEnLUTPAF
qyDjsB9DxGdXPudHxyn0Yqt6k9QErCUNECkS8POyS4HAVnIDK8haUBf+V1WV1ksGb2wuEbCV6CUn
/BuND4/cR9so/nWdChQUqGb35R6GYOwluo2WpGNZ78XwMMjBHiKbcMuSJWb2C4PbdoklFPd6Uea/
ywaAye9fILMStCzWChOqe7Jqeg0C5zl33kDGo9fOYD1OcL2DQkujzFqU+bbmr5J7sLcMlSLqFCOx
1fIbux8Vg+gUAVvM3+6QtGpdfu+hCK2zTmR40i751yKkPc3RUVv1ksgF9LsFc67MxdMvi5Zq+178
Wr49NqeMw78lRjjsLz15UQqMGZ+jLS6pAqQ0SD1omjucjpTsT+maXPAc+92sMIt8AnG9A2JM2rFX
oo6LY6FeuA4i3A0EujIfPBwNkeLWxx7z3XHDb99oE7I9h6Xio2Gg4zX9yS14OXgJYl/se4RmI9MG
VDJyecO0mJf758eKXZ4F710pcRMG2+Q1Z+k1RX6AY85KRBjxlCkiXIJhbH3Z8HYJaXEJaF7ATuZM
0a33hPBIe2U2bzncGWwazDma7a5Q6wYjcLAhNp+E5R9q0nkOdsD/q+KFSn3XyrtfpHX05Wp9r+Y0
PJjG/rVU+jgAXTaZ6En4cXICk44XM5gbZTsSo+8yYcciMgG0sLJQW7aefobzFBPajcIcSJ4v85Gp
yBa3COCarUL9v7gGPRbbbLAImZWManYoY4iiuIqriOeCnrh6GyoodFXevMS4zuLz2Vn26b7A4QtR
uBeH+hV+r+Fo7iXXJbqQyO0dh0fZ0LZW6gdM8wlXafJVD+XA1N71Z8JQcRzNHmGqOl+7J5H+qvZM
sRL9KeC6RzTIPI1icyWukRFVZDBGfODUBk5FjF0FBnCnurFXkaJq8NwWhUD+xNpTq9UAi/d3HlEc
aotcGIjav9jm+grJn5Mupnnhh4GuG67e91yEewy1kXIUPyiy41hLYDbtmAYyKIOyvmWL8b3sbtcz
AfBhynbSX5+kC+Y2Zncx5CgxgdUzSlzTHEo/ZY5XbzCYmCVGix3do+2mOTYY5Z2OjYLjZw7NA8La
N4AWwdpgB3IiJKSn9CDXjt9nCUGrrJEM97zeWo7QYNvMJPnxVct5ZD9Z8RCDUMAggfu+UCVe0kbG
e4jPbn2C3cRrk+Gtvy4Fs7yMhq22vxP+aQOwUDRT/661lCnymBzKHWvK0H6W4U1grZirxr8Q1hU+
c6q32nCLehbr2HF2+n0yNt0DRmgtrKe+1s6SrgQ8bipvTG2HSZJQggLyjBZ0xJyRpHeynPEPafBO
b4GFj5XLyEPG1aASwcjp/nx7aV/kjVEgQ/hSugYSAxj+eauVjdjXRrceLcgs3M0pfEp2elmTCrYF
f7f1pNQK9hbFZeicapjWemTIbzwjTrWWG6Z3QAQlb+yeOghLLqQFI97qRwB11ZNm4t4PdQk4qutt
QQEqNymysF/ao8SVwZ92Oyf706jPiz+7FSaeCAke2V6N//rnu7dBHLJ0cvdpVc7XJ/QO+JhWBCNP
gPTbRr6jnWVzZ/sxeM6v/mQ9wfmhEMYa4tRnfCme0GZ6py9xKiaMDje8d9PD4Dt5ebm9Sq+5Kcr0
Xuedq1EWf5VVDkk3+kPgAaKOLVFuxNLtt7DUdEZkHI3wP726L7ThQ1pY0jFHkIF4cCUepohk9Pmh
o4m5VOsI0QehYHBay7B/ZtWqUa3BYXWJTlrkEowCD7N4NQeoJ3iy6DfTVxIu4XRAAkFaflSegH0p
FxgZDWbicmESu9F3SJl8UnQfxqkQ5c0hObS52cCLBdyS0X/ra4v9rTnPpZyt7NNOyrN7rlqxA4/n
/7JEeiblJtyX+RYvrFDwQN42P+8UqDyrTx4JjIhE6JL9ziKJjNFqkjVgbsms4yRHPu75R9zen0wn
TEVdHHZ0L/wJR2oIg887CuNEnxOB5FjXuRv7AliB86MgGLrsvurmyhc3QymriEw3/5JruJNilUDY
Y6OiVabb9703LE9ojgZ+j9dO6u/HrGZyttTWHdgRgnIaJh2n6+zEAjB+I2P4RRxGvWpXNbrfnixW
6AzgALFphcKTnWyUdsQx2Pjz9bgP0+9XvS4X0H+yYJ3M4kUdcYTMWX+Bec1Y/XpovXLoinB8Jy35
vMrWqeXzCFgAciKFwAcYyXkgkmbjiImNIx1aBU2YyXoBOx+0O0YIcV3gBjVJVFbkVJBItLUNap8G
za9f6eeUKK95S8CDu3cf7BM17zqsyvgI6e/x5y7V7sK1p7rfWuU8ufqvF8Tjn+tXrqdLLa8R3r2n
MH2WAIpghSiT07iHxB+nxLRFcNVemM+6jmwmdlKiNWN229PeEzt+9ADCaQ1BzMyeHe3blW6TlDJ8
vG3rVeXieLgH8+1kuqkg+w+5klZkW75VU3y8ttucWH4RGBOiROVEyk+Ka1AZI1kHfN3h1omK2goc
UT6Q7tSHsMRTx9ubaZlIMrINV+qtRWyPCL3UNjGdWASJu3x6rP1r7Sl/5mLx6wgHn4nBccqvw4oF
cP9SCv8/gyFcKqNVLoXFv86P0KSaqXKhLlv/NND/fswdZHpN+scxPwsKB3FHBozkkOl+ZdY4J2jp
4l0AhKEgsHf0EjomOPNNMDcgdthEXU4ewuSIeiCk5zijyk71tfW2GuRBg23gEHDyquSYr83g2SGk
O7KqoOJukgeYSsAwo6Gbu5BTERzF3YWlrsKnKAkGKpJFK6kp/Y7A+wIbVF6SUqqlhoRwL8OItmUi
+eq+m7qvqzXceAVVs8qS7P2J6IrFmdEKgAoDo2frbNs54CAkMeznvQNwCfsNdL6WyVucOMQTVIbI
SNDR7FueSmJJH76qB0qz0hXIxvkgJs+Si1RpcKQ93aCrd/ZgFVqCb7x19vtiwxIKWqQxmnmzm395
cjvcPdxKfLsXeTsG00ta+A/h6LcODUNey4nt+mK3v0XrFmko11d3LIbS/7H4A4tTBh0HHkGsZs4g
S8fkaCRvelHloufwenTNGuR5ljidz0ZcKGP339HI4hx62IoGMbiUq0ObxBHOdClXpJkSPpKygzf7
ZUqrHLOvQLWfZ+mwi6XuaIxnPZa25zxJgOG+m1h6EEt+/ClgLaU19bYoLyZFew7HoTAXzdqKzxN2
tVEAMddi77IyuNOxB62218yTNuCHILfLP38lOSTceX2jJ55uVuUWkuHm+amN2fEiTJ/GWS5IpM4l
uqclwBnUln23IRECOUUjaCyl88sS/f6cGM7tMag76POz376el3CPZxvDJO8osILp5YueWYF7k4V2
YrhMlsNNhEM6PdHw+qLmOgnTccwbhcNeZ35y42NDGUI9xyHUgcMdP26tGD1ER53zwcjJWmPuvrk2
9fZk68DMEc4RNMY+vV6kv/X4wX8MzHK/cjMatSxE8kddzrppPH270fOFBwgMSlgOy+pDLCwoz/Hf
FAV34Lt1KJcXIziw128plDnNw7kl4ZjqL9DbWf5pj3Kck8bVyNVKUDPhfxQge666G001nxuf9+ZP
RtotxRcnCIFGIMt0LYZ12YNAfixsc2FNEobcF4YJYNSObWgn/uOiV3uyVVRKM6U94a8nwV99K28A
t5sB20bxlMFXX/79e1hOupOJCBAq31lfaF/Z6IU4vpaIsFqfO8oVsmOtUwZalW4Ja0BZp8INMn7X
XXzKkRlraEAHrU5M0PGOUKzxrm0fG5IFEZ5T/Eeen30sRr6WlOSts6QHK4IbmTdQ7BAFEyHRwelQ
iPNhUFop/yMpyuCx/ruHW2QSOMaKVGbofFL01GtHW5vSHRv67/lvvoVEVlUXADiOI/DjDwzoZ8S7
VWmpU3AwGO8LIWGB3zoGVL7OX2H3V5IhQWAZl6vz/sESAea6a5ncCP8Mni7LFpb+KeZ+fJQUgHgt
vxAkf6ldQeOof05AOX2CSUOxsy1OAsY0qF91Cwv8ejJP8Jj6C1Ihk4a5L7rJtGmazgvXEmJ7N2f8
4dOjFKHPj0jCJCwhV3b2XLIveN8cdb/SJWRid2Sys+TCK9JfjP0gyAmOSLIWoANJSobG6tJSo2Qd
sjkO+tL47ArWcqfkun9BzAxuQvj2gC1ZsDYbtsSD84TLS4Ew3pUJSBnRFeB1WsWrJAcIoQYraGf/
PFYKujWjxB9RNr/hORMAIjB2uAgupK+bhx2FtrD70fDFDx/zjSSLUxqc/ngeHS40QAWBdGM30Vtd
wl2+Hl85tyOST+79h9BFB3g92+w1Sj6g2Lf5bAp9aUDrm+CBRUXOL0vNgHKSnbmVW7mKM4CilRQ1
jg88wW4uzj2pGZCYA0XR//tg4EJGv9g4jsp3pZbi5MY2LSGzdWnIyGFPCFdMYybMTZjI48pS3Bbu
V6Yu0fyLBRsiQxc/yBRF8eyyXvDgZQq3CTU1jiqrVECK6PqN9gDo6KdwFhELxDdhHoLWG7E96Nvz
ItlH21+rZ0cdn+MsVIZ7VAhCyvQgShSH/naMVkWZVdIOtsxNovJrgDlAqpH31r7P7YQGNsN93/KV
O3BTunvKS3IzPNGw56cj1hj9Gg9pC4n/uqRupA/79FbWb4ZSP9/JGXAOOL6eFx1M3PBPSzWA5AkR
+xq/2llDkuloMyVh6QlIj4fMUzAgnsCTnGtwhcOkhqQSPM6ufpyU2dRu1UHtEdTEqVIWst99Jtai
LGduytvye+Z31LuzViJP4zDiNvd1/lat5vhKYZf0f+8LWmjX3fV6jKBwUwIYx9mLV7vwbVWuu1Bq
23CrfsbrhbkQL8iNUC8Lj6hT/9bkctVnaiBPDF7A0aI99g0fbrrvL7Eiy1mNo7Q0eOENl3K96NTX
C8AxmRHObPaUJPUVuCuQaRfR6QKv/0XkTAlAczOCi96A9QGoCH5Kco00tfnNNC+d1X/an3cPNyJl
8aJPIkCs3a0H9reTsFixYo7+OlFC/eVYQa6fOe76OHIZMMpujgub62QaFk5x0t6wqZHABxOy6cTO
w4IljKOhnF27lWcet8zRrkm2HMPNdfjHyigKZW9XL/6wb4cvLXDzyslKlBL64kI1ogUjyY61UauH
Nq/vkMvlZEfiLIz9Cy/me/kzjVT2fkMcc1HNENxgKEScXQZf2jNM/kM3czkWSuh6b2ZLvtAZNiLQ
e+IrkxbkdvZz8J0ex0RjvoV+xtYTyvvXn65LUZUOdWdiBed+d5bgB3UHFuLOSc4aH2qBRIn+b3vr
9HlFdrn8LV4vNtWvq6l/VDrahSwdXbKJKbBMZOWZIkQVaKi+zQoKgCYXUjJf/IdNpInmhZxAxVjG
OUz680ZoZKmCxYKMupBwaqv+b5pdTZXfHtAcpdR+bgVcczWJ5rjSmvVpYF5aj4Tnb4xga8sfyVdB
GdRCD9mKmyZxWp1YYnhG4bQ4c9dmMg0Ke/86E1M+qmZwCIiwqNI8N8rVmkt2NtkJEjWI7XWPSByf
qRoWzgTrIwt2l3QtFKMzJFkA9v0KFT0nsH6Gsonpl7/smFHOzjYjr5L2cnzRjhG5sJEM0rFEj+Gg
1K8rjfv84zqwCTM9/4jcUZsXlG3g/MP2GHK3VMIGnTOalOIA0t0c6ylTjJE5dMc2PutZRph7rpfS
uafYNlVqKyekDFJFRjNDT2omd8ziHkEg/rbG/Da59MgYZjl9/m/Nl5KqPSr8MLlvk3f03Fgyv4io
HSj3rkuCZITFUNfa/CPkMuyJVMYJ4ooHKh25mtOJS0Fcqu4Gt+Iy8atSrP/MsVfIHbuNcWQwGvcA
D3ZZFqpWH2x3sBt9q2E0/5sJm0KUif3H750XSDtm6kSRNhX0cSQAiQQ1a+BYIu4gn7zvN6Y8duJh
MraeGM/hsdE9+yPSmf4687+fh8qAR89XnagBDASA+xDaNVDAoRmtqyE046JAcywS4ONRNhf/n2j8
jlhP655lsHI+S1bQVFUgd5sL2XV3qaC5nIW0Fh3Rjulxn96QTEEMptR9ZDfz0ImdOfh5vbULzQJW
7Sattx+Hd7Azy2pW5IxKAO4xC8YO+f3TpL2OG1bl/ammmgH992Fix8e35sjNsB+RynQb/AM8X+Hi
TVUB4blhyKsjZx6mh0U2/pvJtN0kkSZQILAuMnGh8hHKbkjCUb4sEDee7i/vi962nrYbeXM8s7pR
7G/4UjjM4+3URdoqtlUrQCbN3njad3kdQLFAPPT/sPQjVHuNBnvh+EmRAyTiR4qDa+vHy9t8dvj1
IpAuXYUADZUir/hC4h7UoCmfKMwxFyL7PWg65qagxzPZlthcvpMLUXlXvSbAzF6lDomNOt3mUIz7
9CqNsIs2zwrSlTtJfI0TSKNB2ZnDpvtm2uwaMpEFabSgipsplB7Xf1ZCNCYjc6vtJiIPyfn25Dm6
J0rdcONuUx2LIh+ZDZGUIKI7aPDDXo5tbZ7MzrvkRdMRz4s25i/fTUf7ad8bie3QYYBBSXa1ptNV
PXPtqI8Alp08274jU4jDrD/L5fInYVNuckaNuPsIVn06iHuUw5N3EG8QCWnYD3kjUPuuYXxfr7y1
S5dQH9UPM/e9iOCXO4WMjIQdDMmbRpTmAJmRuUG05Te6C+3auvaKp4Mnu3j0kxxwG2OqLysLsgJg
jnoh3J3PoUxPuqq2aKK3+DLXnm2nbyRiQoChAkGm5d/R1MG196ALGYAIQjeU9dkyzmQ55JRsnDGQ
7LbF7i2mv1ZTKESZ5yMMMByqZ0bJmW+6dc6s+hCpSn+2wvz3QZQce3SpmQmwPA+Pl6axVEFFrUpW
jdJjnXwSOLH3ke/ngU9PgoIM3EHrYhfoTuDkOfyf3GzOfGHbic1JllnZAc+J7p4MyRUVznAoCqx/
2Ogxt361Xf+js1owPsWwGxhRvQWZHprcRaS7KFq/Wz/KacfdSD/Jj3VsBuiohEGa/dV5LDnLG5YU
bqYya4bXSRoL/+atq+PQrq+3NYFD9LSELUjgspjExY1HjBo1vQBPBybgp4UDXfdmSrZmSv6GK8Nk
ucns9Ig00uinfdIU4sQtHArJkkXqgl9XAKZHrIEdgYnN2+mpdJoEZ5KCWifo7T9VNdzmrxbhvAaV
VClphgrlZuLgB4byAqmF/hiUVQmd3wzkowG7KVvxD5XRQlhi+Co//3wS45RfyyWK0vuMeS37HPWN
XgQb3vb7aYJ96HTfpAjsqire0lzzxVFchRzyWtSBdBl13EvlaLk0OP/MiXjCN4u8koj4PiIORMxB
2MVRCbIAkgudwCmPGq9iLVjwOuSHAM8m/7vW2DKYjAAWUSdKqhmPXvqiCjRImxC2iHuKdXmlSBOt
/x7a6MtqPJ10OIJ8kZP1dUkveiVv/LK25J8MROL7fQmbymUDUL1z5wnNAD9jhOU8bGgO3izHeK30
LQdT7JS8hFBGxFrwkjSPE0iJik1y4TOKEwUscJf0TVg/hSO4osYcIdb898oXPlUmPCDq3D7IAqaQ
wahQ3POxUyAYOmpxwHydrkJtsrEzro8LMU3Wj0p1PCk6XM6QknwRjUl72jNSdvi/H8NJQfRD+cFD
0dEAhGt2HRFMfEUduGGkMgxaFO2sr4bKhzwiNEmcFpJScQ3t3emWQkP6rp47fBT/kaqwQpVoz8A+
Z3mDvH0b+/9aVSFAsP8XdqDCXwbubkY4C8ngrIZFnaUZrR1nZkCB0+I/0gsGfYPtnZmsyIkk6VJx
jewg+9AKM3eMJ3kUuJ/QpJDf6Vvnj3nF53zn+JtxYM8m57BTBneC7b9nViOBzskgPsL6ekdIQP5z
4gW+RLD4fsP/Xi/3QcT2xA2mZ/m64tMejvRLISVNDAzb2mzPcqbCYis9l41DTb6yvQ0QxLM1/yPk
bGN9Tu1c6UTYSD9I5aTzkkMpB/77Xpx3nrfJXv4497UptfFIfcP3+C3GSN+GVqxzkvREzJe8vMu4
PK8ukALSK/Gh15yji49SSVbSYMuhjT2S+yukyzjQ8IZRXsA4C9lOCKsZIlTD/BTjFWC0gZS43AjS
dStiqdhk2LvcZBoUSdLVskdU9FSrl2hW9zdLhBPgIbag+DWgd0pl59KDowPAx381iVIi1iRtjnKY
18T4jdxI1Rf8DH0aqApMy9t4rJsYmwFS5zMwTHFFtaCCl4UyERYMudc4tM88nhUMWi7DD9Y2tdak
YRioQ21qnfg/Wo+0F2+vhBrSVBzkpQ4bEMeT85u5dj5yoI/v7TEidemi3FVCm0dgv2cRoL47eDN8
hxFkAD4JCAFtZdw0Y+3l/ITdzp0Mq5GSHVxZCXqrhUbde07sKcSNpxha51M7BAiv2QVRuyL6V5R1
xREKK9OV6zI2pMZrk0ENnSDmqWN/NKy6qT/oVW1Ah6d0JandRgSBXo97HO7CdMlzSs+8Z5aYac6c
uZNsDQGdtK1sYKbAg8Trl3I+3hIGZXbI4HO2ZE9otiQnCx0ZKUv1kGDSPRo9cwoSEG/q1OIb3Bhe
3t/8fu5Saqs0O+A5OlncPN1KRq2b/cR0w7EFMKWAb1K6hiAIdjWhJ9bZ5BROa8D/4LWcifZWyddi
tOoNz80bA0hDG0eLsj9bvTzhHNiqlJIPrnRY9003RGyTAzk8VPWiuJlkH7jQYaT0hKBxVnNtkZD/
RKqBZ7Z/Da+9fQpqT6xQc9Htc2195bkfs6rUdzVpTr3wCCqSQDbDBiRx8kKryZhw/Rj4H6NNFUtC
NhhIy0Ik93A/KUHZRWI97M7dKgueqsDAP8dMJ9Cac1ETsEW929P6bJGRyF7HDiheN/4DpM94qQRK
g+pPbz/B1yqLR9Gx8F9fRi5tTzrV8dWdnIGJ77XQGFdt2mlUEVoMeL3uh1+hIAjOOt8pDXd+soKu
+zybMlXj+LyTIILNIhWHLUvJJAVe+aXNaBpDPnZO9uR1qtSr8cgdO+n9F/n/NPDqa+Pr8ekpwZPq
6YiuMWvtOPq9fjBvF0HQkgynDj9+jjI7YGMMTodFnEe8+xYpx6TeOPliMFWM8jBR9DfUx++N/ngy
IjlvSmrEP1+EKq+zCg7U/6mPWrKbLrpPYuD5DeZ8XJGodyBAMdC+7QVWgDC3MXEuGfEeZEk5O4WV
JV+GlUVUlms+Ht3B/WK4awoYeuY/G6vqKVDBOJC4XantNeASsrMDj/IFCzxokziOyqelXRU3Coyx
UiBctq7iVPBubPwhZ6S1kJARJS4E4XsvvkXzMZqv22qe5g+0g+WLGMVNDegdCC9xa9NNqBAQvwdJ
lvffVPbZpsP5ofXK2eJxs/0u+VU6/+HgfP/6KQ2QKA8n7fbQUJ9oaLO9LexNQia4qrdYnLvahozo
esy35eT/Xt78OIjV9cR9w+pTw//j+adWpLDvYOOhvBmPwTjMwgQAZagjbdKBYdbivocfwEkfVzP+
iUrA/abWwdjB82lOLy88ucG37vLgWRsSpjWqpxWn9b5RPGsqsiJ1C/Fu6cBuYvcoIXrgeLe8MgvQ
hKKTwx5QFGEHq2o+bmzT0Ltwemepi4wKQFqXMc5KGQ6qpdZVnuHSC6IsOns9U82dORmrgcRji5u5
XrG6qWcsx3vav7oakfc6zzidupMWSR89gwoDkVfkmL0zIRf4YOh9V86nzSD/SDIMbolK/dkfNpMF
fBnPAKlwl2PxNo1BCH4bXr9ABh5QsETeA3aew2xq6v/+p/tWHD7sGsVnF69SjnPvDegrbyumyAGd
mCJ7zh1SChpVGIz2qZRn7mG5t1e7hu4LtYlBDokfasykDR29Qfmk4i6nNQl3+BmK/0XcNbl1SbAx
GBMEnEpPzgJpiPoemTUwpT8yjWtNNkcgzrsxDHhdkn35Bbdu/VEXnbwBVK5wrnu8dEJqiEFjfWKU
H003lTJ991nGYOaMjYKGIsXkJ+SVoAEc2A714q2Pvh7i0aUrm5bvR//flNKwWA6t71aZFlX/PgTS
fls2On7MqzeIoUhT6Uhs3mYmo0wQmXQ/w10rRxfiYaxlwAknl1v+oSK4zsC3qJ5LkXoxiNBcHPLP
WFYuxl9jYlxNLsi54AiT/RFazTxJ46PdKbJzLfdzroQwsunIfNZFs0kNrjsCPonfAssbMjQva5oJ
ulsCDLROkdXnpaP1cOWNi06bohOSr1opB6NtPkDzcFOwzd7OSAg+xF4YfQC/J6JrUATgfij3IAV9
0z6InBajSMRlmRJSuLrOz8V7oKt83jgC0C5YdRNE5EK46hgWF41vuXrh30rB3pkANl63JOmwsirJ
63GWTzFoLpeSW8fvTpNI/ZqlxPmf7epInrdvUEsoZv2m0Zbd2hmv0smBktBNw0cYAKAHF/qzI/g5
6zhXcffaKPZNALiIlwMq3KSm6yp4oQXLQSagQ2PK10xgA12Qfnfz0MlBz53jL8TT6HSW7NtFbBU0
Je3Jm3vbPzToC19JZO7vOd2/vjKc+fvnyz5Uuq8J1bNtBHNZNAOsT08/tqVtsDrQAxM9MGqAXK5V
JWwSTk7NhYkGrnVsiIgYpcBCGvv0xSYCG04x/jDipWmUX2VlgG8I2Lb+o3nhYimhbo0yh9OOkJ0T
KlUDl5nZbqPRBLs1m/qo9h2AJ1Z3KpUPAOvRMWZfv1awQX6UCr+NoxmUnZbNueMlr3MaZPWjrIwf
empFrnBrZMLXl8b9v5yXN0Y60jy2cNTmm8/NRBN5nidXj1VbS0h5tycBnRyJ0a95W2IewkaG+oo3
nucM0Kvr9VoyxT6Nf5A10Cmd5OeDbxU6JL6aWfj/96E8vC99B+KtY7NKPY2/WppaVDeRqHR/cRC0
JmE6Ne7+gSFBAJrT+KQOEdtCbGfTUXqid9oo0VeQ+XcbaomDE6cKlNncRthLvkV7hjWF139Mrs+Q
pda1v6k2eQ/6wLYZfjnYl1rYTq6udcBd9vOfucnxZWRFnctpXDxVS3nTb4p+8pdusfeg7VkqWpYy
WXU6mJaxOPIpCbwLHYlQM/uJGOEHF4LhdgDg+6sAcl1Kig9OqdSE7lJNZ1fh3hZTOuV8zsGdRfvK
zEIhD/OaG/GtiPbFiC+4xhceKhuzb2PlAWuBqUr+DN+3E14capMusQv5Aw6oc+skFZpquknvD4lo
cBjkqzfjey6lpBJLLFksQiY52LGpcopQIkq5gavOKHyWtQXijFMKH5ABrxfIpZA+9lhF7Dv2rXvA
eyXBH1/oiKNN9ejKf/T0npGggbjoihsYnmjcz3MIgyQqqSWTlhyf4zpA44Zqobiwi+cJUp9rFmAC
W/oCOG5hg0KVVmwHGU0Jd06kXFMyNHGoVBp3V1Eo0rCN6wFUGIgDowFVCY0mkjN8dhrmJvdeflVr
boTrxK2QZxYdhhouRzfPUP3uIEt3fe4f+MEOcqtF+/zDdHqIVxzB/IRZMPz2hKdZdPafMTpVATNk
08g4+n7Tr/lFvsdruGxH6/jhIr60I2/FnULZR8v6DM+pZkvidZSYnl5D/je69rQFo7jhqd7ythZz
E7CEWCSeeVxdhQrHYQYpp2PT4soh7DgdDeGf/5Uy8OrMPaYgskp1uDJ7MbzXLz5fj0LTk1RQlKXm
244484k4arhMtr9x8ktuSAEiRkD4kt0Fs8G69Init+diS6OGESy6W/d4g+9B5y9tqhZUvaHwCRAD
ujXF1W/FuP38ds+MWXgcil4Sh1HqlFOyVh2wUCg2qvrSPznMRjzWbtXBY9PGWPlHV1GLiJBX9MNR
qWwaOH5Q91PIhmMzx4UIOvCTT5qFWVmCGbCIuGnfM7WOeAERVqiQLTJgt8uhRxbE0OogDmAu4Ky9
kz6/2wV+BUVobRE+UIOe5ZXAgENP7N4NrqMCJhXmkd2IRFn/lC6yb8YCc4HmAgfSwspCznMrA/rL
AHcQNk/XaQ+n+ab4tlDZDbLPbaY4HrFDB8ueJomKJV63qByWF0nYnnySP+fKRcYtqSdirIiDZ1IF
JTvUNX52HXNU+cKdTxTYbFqJvw/fKVBs2PjR8CeM8/LO+BMZBrbNjk98iWbTS+2NNhfxM1GVNT5I
rRH038ANtv9zxucjVKpEZIr4eWZANOKLv+J1+CmTRspM+GqENBXi5ljWmxh0k2D91QL0f+bFgA9C
KiaIN/Tbh2NxYITuCyNz7pnedONX7wUAeIjUS4J2ZkUkTF2XQlTb/UdMpt+V77kQg3YkEzGN5rE2
PoRMbEavMLCZIH7g47qjPnVMbJP32IbxlamcsYDTygdGbG9SwXWDuaDJslLslh2lE65oypcEDEzS
SIsWTu48JIxcMnzEceZ45BzTyqLiBTk/Vvcz5px9Ub0wSVHU5vCDaqhKqQFMmwxFQTyaEYblyBmu
Ze1UGRDHk2q0Lecv3mHEEoexXETUjKLIlsAjVaO+CPXKN91ytwsTKlm+k0j/0gTL17/dwTStZLDm
G6wX7RuLJxLqNb+1Hu0T0ymJ8z2enKhRr/YoAMvByVWd0iWEl0NFHZPYnJ9hVXCs7zs389akDKf3
Hc+cWicWI44lJAB7I/ovD6UuwJGmlQYXSlfPypHnxZky3tHrvOOcVSvqJNjB6+bLcfJDe9HNMl1W
Bk2E8HMPBwB4NPnOi82HVsbUmoHWXnqAeyl8ufgVyDC6IODUz6CEEUsP5fTaTZrHtlu1S5KZLK8/
U+FtV+yN5KHehHJOzzBxGqcuzhi2HQHDOQ2LuTPxAFSOHBtiC1hM2H6ax/y3nJOAIW1m+l02ta/U
FWrcXUUoKnzu+kkJ3KSytdnejS3nEQrP7p20CaaSbb0aucSHRy+aB/0kkr5pcR1CeRJjdQWd+r/C
3kfVogiBUSXWt31DmuQHXMKd/m/LWw2RDcEaWySDHEOqdzHNMNMpG9p4/hqi3cEhwhUVquvPi5Or
u9kke1GRwVbkZ1QDGjRX4EBfyIzBAyLj4Cq718VKlo+GldBiv4Mwxm8rO2zWBT0kECpujfgVzB9O
kAVuLPAe08SNpxPkxOhcUPC0mDi2VkgSoplQwUviT3tBHUcw9AuMEd2DzevX33YOETUSMz4yFiKI
+hZN3tdTrM40S80EXjshXN/5O2fWK8oe6/oqhMgSOuGnE3lMVVrkLbEdug1UkznqSAGDTix8XOia
DFEL7IKXD5vyorfH+OXrEgDKXWQbgQ6F9J1AWqS2H6izhfraHSnV0RHzQiTXG5M8TfDxtXlI4jqr
Ix7Es8YgDgsWZCJ3M485I+wzxD3wo9wlfyt6TwOqG4H3yLb3ly4RjBac72YZWLVQ6IGEoGU0QxN8
P73GwWGH7CMlgotKyECQI9fRhByWvX504ocxh1GcSGrpTpJLsr4+ljce7XkJjAURJ58EoW8hqgf1
1iggWlPD3p1Y9jesXVgEEl2+GZHL7pJAGzum46GvWd3rOglmFphqVrT2iam033SZx1+RzOInQYL4
c57f31D14iayTQAUEFIemf+LHlL1VO2LoOMk9J1yFw8WKJSMynZ9UjBBq1xex1TQ3YtkCEWMKR3R
Z6emVrrVhjOKlulRC8g1VuCxE7hQs3R8OMHPXa3TRIbzHBQsKa0kNUe/fApsxV07VnSqdrw8pzdo
KaAiYjqNSoiKHRKH56/xoGWbhFJuIUb4xFCyrIxvdxqnm3+TZBBrlyqS/O+0QLbIBDnO/lyVCVda
OxkRqK8fYTWbCDmuivbGBeVk+n+4Q/CVZBOnZ+uHADL2sAHE4BFJLP08zLSwwVEt/a2Ry4em+92h
I50g4+zaQ47QSi9lg7v3I1vj6Qi89zALPpWG4YKelesfi6tadLNuAiXJq5Mcv6xpibQKtPNw688w
dQfYUkyO/zVpgl7m9RGCK0UmbFXgyCQTONVlaG8FImidiODqET7gAN/s4UjzfzienzOP8Bgha1ys
e9OTvfJejgSyDaAfTApf51ibMiJ/+k7Kc1I2libmdHIOQ9h+eUpP99Di12iDybQGlbwH7knma2ZU
+gNWYfU1eL8EEtdpnwjfQ4/pQ4VJzPCzVbidpobXYHw07Ed+JU7tIMOu8iZd3YWGCgxSjIdPX0Jh
epOj33he7JdwQwHpiwzzwOgRX9fTHWyFgu9dLIXR3tHJe8UccqZUg7l11px1PDWUuUn4ZNhz7Eib
FCeD2bBHlDiiuPcHDRNfl4+jCZOrWKPePu0skOfj9xnYRfiA7cLDkLaBweJl8tVo0YAPxsmu29eS
DJh0jgpdU1xK3/5Xud3esbRt8J5oDu0gchfrzGz0kRf0U0YexyTBgaP2VPUUWxLlF8SdELep6XKT
75vkxiHOz5mZIAZSabsrZ9vRmhZog3wvc3ctbGbQG1zwQ7jNTwyoDyavBCkWzc1TT2dBFRi0WU8V
8jq7EwkdtF6ofpkcbYtym3wJ2KgWedO+aJq1LcpgbwT6O4xwt5kRWPxHIA3hNfu1Z+S13F1MgmAI
DO3BFfi3c6jrzbeWBc1vAZzuuY8xaR5cqDzYQMOyaOmw9+ce96e0pwY+RG5k72mCbulBu/zgxX34
ikO9+Pc8/p55MpVXsEJX4SzqZq2wb738xsZoJOW5TiYk1xFrXidMS3dVbOTFFpJ0gNM490a6/TKv
VsnikJ04bTNyvMm//qaOXp0E5DxEtSzz0eHP5YPiudBuxqokO1hh5yaavN/j+3R0pPX3gbvnlP97
Ja76tufMNc2zkDsH/S57pe6onXVYrTp4lhYfiesopFBg0iMBfyFWuL+0jSqBb9BGKLkMXxRdiiPh
tTDnBZdEaCmmbDVSPZresFewaUnaJyokV8BURRmXsOzH7CN+fqm4+1zHk78ub1RiHmNJJaAakzTC
xK1lKY+3doT/J/R3KqLaTQT8sAriEEFq7IbMXmGc0gUtr3xKLXOiSas05GFbOQ8lnOJLWa5IeIC+
HJVbMPrZGmaF7Fc7nhYxw+tiJWiOM1wyzc10eESYDhsvTGFGShXBNFP4jqcSTUXB0QGCFI+Ts9BR
sWmlWBuzHp1yJdEd/m6dc+6WrLVT9L+w1RLqX3PJJ8KjQLxmRXouY4DhI0q7FyRMNQfnUjGBRwG5
oRk9BaWkOBcyIRBJOeKdByJnXREPLglY+N23SZmYHRvj18nTW/H7jLKu2jiwzt4+ILBs2BS5E8hp
o/R336KJ2A8of7OSQwSB2rq5atRFmOLTqYD62smEI3UDl6doUgtYRUVNeqbOsUdHdz48CB7o2Acg
j/Yb9lZNCFURMo8QAS0yIa2y9PZUOEzw/nxLfkB+bQ04tZAw8G+JolKfNl4a3ooBkzaMOsQ5I0zU
ebd3SO5HMa9s1tbQ7uPI/v+OQDs1rTA0IIAbA/Z62/v+udOQKIVljqP4GkQWnp0ItK4LMn6Usq+6
Q34krzOS8FEnCugezxKO18i1pOZ1Yz2Xbz2OJrvNVbGNY9i4ynLpnokLB+ujf23tsJ7bUW2iz934
WqKdMf9nLBG9CcCaWrlC1Kopx2/AAr2axGeOe9ReZQbrN75Ph9prY9HdHXDis8Q7HGaRijhn1hUh
G4OIrE0opZx1q0tdlG57S93uXriZkNh7/kl4NVFIX4caYX3n7r54MATq1TwW2gIOKM5wp1q3wh+D
KkMNXO8gOehcjpYGO3fxt8nwCKqiItkORXtwJMu5DGj4md9PxgOueprbrXuO7HYZ2XMhT7KnEhry
LPZ95eh0KpIeMG6jEbPlu62GFQp1/9PbTyM45z9CRm7FYxOni84Lr5aDHPP1+HINr9ACIHO4DG6K
Qfib8jaVeFvBoV+0fzYUPHzWrGPBYioP0DJe8tty5AdJMjA41SB7S/W1/2kFASIauDOvellfNjde
5bgL232C6zz7EtMHFfDFMpw00CrSthN9fUuEiKkqI6E0h47ikNStJEA2VjvDddxjC1jkkSrKaYKO
9KOD0R+rx3CCXSwATynWTaTyE+AWRf0T/ib1H03sk4pqT7rJUDuEgC0Z3uKG3FxSSfov8bb9AHgY
UzJCatCIIyrPtGmCHISiVAMks3dbdZxbFYS8wEdgVDamXNC0t5MUWju8EhCQoXOq9CgjkgS7ktoR
nwf0T7hkPmf6gnKSCYlm3Cw3V3n4bHyNEjbkVQhmzKkHYYbDk0Nr4KgZxhfKJG7mkDLQydpbRFLm
5RxCvttLOI3lsVTMyFwX6YHOx70Z//SFSFUC+u4GfSmxxQ4bDasuJM3gLO4q+FIrQ4jufhZnUs20
v4I1ZCTyM88WtMW7O7h639K8cP7A1ygv/Q5P9+obeMxJBpqhRQMR/kNY/cHqqDnDE6omKpPebTO+
AJv+8cy6SKyGBlXoHOJtvB+5IRujmpwihgHbI10dK8QixJJaOXq7ng4Bl3hk0Oxf9Rl6Mm9/uSgN
Lf0Ick/YTw0rXHEE7gasFpM9U233zxIl9Kqv9X/ob76IVMLSGj/YpGz8A1v9fdPu0vlxOYbCiEV7
zI/HiFMqb/eHc2f3b98N0AAQ8MzccSncxswgsykkLQfKDEgxv4KqPoZe3W9+4JJXret3nrZ8Qm5Q
91NjMMCIRVfaLKtw9fz03MDNUNK5Z+whT8k3X2OgAlAbzOLsrxqxGxmiVu3Qo52iwcUKE5GpvfNN
EWxbHezqQxLdX78tdM85m/dYL4Dtn5VETC96fXZYiMMNoRX5Enw8IWHKfMCK/dFe2DKnDeem6sjZ
h1PKFgx5mEJ90y7IU50J14e3+SDpbNzF3kGD3RT5DUjmbcpYaQoPgPL81Pkrm7cDV3gIx0VTCWH3
obWZPCLxXhnY4EVEncFBHVUC+2hL+qgmVR2IcaZEseYEYvrv7gccXBPF8ED9+J99ljYZmog92kwe
lrCZix5P0udkR1atd9v355zVT+ryecoSu+JA/LLdhYq2CHg5wlGhkK4zac+yrXLHDGOUkHygopbv
nrWmiUYhOKnMPDQ6BsAjuCWKMyA37xdJ2IFVmYblWQ99jIsNKjfT5UkkkncUBHpVbiX0UHbLFpnP
yE+Rl4Ad4breKzX0WskryxRh2pFObKtXTD8iXOLpVfm8G+ZbeoIKTqeC9M+IEs9UYerW1epYqv6E
Jn1NWTrtMXPrqjnGmgFcDof5cltgB/ib1pgQ32DBIcRsOkNzLzvyGJyAQVef6skJ2s+8cBwen0lD
oxq3Ty9pHtrxX2gnX1hsq0ZMfLTxYGavwD1ltFHYcQz3SDEpzkByHvWtHxs0p7+1ZL1k+JsjjwHf
TwaNK1UAtNa+O6Pz/KHJR/a+yVKBsbLIjaR13Nwz4lt6S1ZC9dFtiai3y9ZUoYxsHEu1f46s0GXp
dXcwivuwXjA26feM4yJbRnRXQDdwcuVyxW8NbMYplhMhue7beyk2WHjO0xqAEpqlQ2mleyCZq9Hl
glyEdtDbS3GTkBql3OunD6MuNbnOsq5+lLAoJ9jighaxNZ0E/jrKLvBckUQ1lWqPj5SbZ7Y0MenC
LXlMZoGlX/371XgZ1YnFa4B2kmY30x3OIvx5YU2IHBrOYm4mBC5OlAmabXND6YrXxqbqXa0FOmgE
tLWHFyZAaZ26eqlTLhB6K/WCABrj4whjoQSgyp5FsGO6Qqu+7Xqt/G/puTGobegnKzssuaPmZoEc
jiRbo675k1IT6gPN8D3d6M08/8G03iAbA2L7C/pedX2MsdzfxQgSs5QgDqkK4jrU4Rn/uQN8M8QH
2Og9MMhc7B84CwWTfTH6e7i3YkGVLyqvJp1xPtFvOWLfj5pEJfDoD3rY/ATNSUEAIALm9tQbhQeO
tJee0n1sPWSFk8TpAsW7yKhKt4S+AYQDeZT1kc5OIYrMqSuWkl+uRDMNnlltctep4VW7S37J8XvB
6852q7Yj2+IOziB4ysH5PKfKSG7LwvKD2limaNSPoC7Vq2DQ6t15jtuBGNxRfk3/1/RVbctXivjh
IHvBqA9XNnJPa7fb3uyiR7hh99MppGixKFZBcs+l+tvABelvHY6l+IStLz92NrLFxnnOq+7t197m
lZdxuD/NKamn7YuQ5ZAFsjDtpCusDlX4QC5Vzuhh71PXLSEnkQSmjo1JXWKxvEzoLMvHMMtMeHxu
NGys6+6Ipd3RowEsa6I9ejg9Tqw2MV/bGvve18A2CS2vMYqCe5WzLkCO+xDin2ylaNYwxgmk0U6C
azq1BnZHD2SbZj/zqm3lazDuRRUDXzw9LJ1//tVbFVyY5kNRa0DDb2r7pEgrw3F7P5XsoeYX0AFP
ixLbhLYMd2BDmu1a+dyLe/n6Xp9nsfuUbYHh4WZnbgc8+0nIY7CN4UiKFNzEjQRltRfqhhabUgAp
kRemVebJ7IyaUl/Is10RLhSIkN0rqSiKqZB8mcVGTLD5S82Jl328XUgjjaH5AYPtJ+1IU3mI3o/g
Vql9srxBOYyr+zEh8L/+nK8dPbgDCd7iWgD0J3xYLMZ/h577d9ZhcGV7c/Uu35mikYBSD1YF2t2G
t1GFODft5vQ2gQSbWkpa9wgIySOlpqv4vToOlNPlmJI3jagNNzlo1g4RocJ4noZiOpnWRsNnDtwE
3xigBFeE3hfP33S9/DHXkx42eMv9loJ5QqZCwpPI98hvjjVgHSnDC9JeemR7gmJO85POQpb5FKii
1QrhZSkudw9BJZ0UHRC8CettdwHdCdvVKmywa6Fv7cnlgD0E57Fpo41zyuEqiF0Pt71s1JCYcqH3
waBnv1Yx4gMt52Z4iyQUpQbHMgKvdFJs9/iZjld7uk2x7Kf6NG5yBZssbhnC5LYd7k66BFEyW4rd
Qc3OBpKE6mgUYQWZXH6wdZ84c2vfadPdfeZDv26MLlwL6gOmjRVvcS4G9pXV+YEkRXveodkddxkC
x+6nGF4FnN641XFL5EhrFBJ7bk/C0lCXBM0/Q8RihSdPDJ5jXi2boBYRarDGQv68w3MAzQeqO93s
UyjiTmPu0V35Bl/cZervXg9dDZ0m+0A73YcX5yYeufmcFc8IYs+wDXvYVWKkohkbD2CbLY7zWWnr
bbI609uii5gQRb4t7CuaTb1cLOI3wblfh43BMWOrrHiyl2EPabr5UeoCTbbeyfQpVeILMLdfDvxG
dGYzmBQdSwlohhoVrMvEGtym/wB8ktuVWpLHjgOFgAm9np1mkaWe/dQU/3k5cLs0iSDk4P2tdUK5
eQaxoFXykFyKE2zD3fvWozjQsh/mSpkaNPJV7E3uo3uGSlRRjwf5rHza1Mn7yY9sc9Xl+ljp6ihV
CIOAI16SHsZWoqRJlUU9XzOvpe0MByWYn83xo8IVApxKvJ0BAYTJRmuy0pCWA7XuvSOlxifSvr2f
NGwkiWjFd1M8csF8wyv9ymWgwPyL2pGDJMqNE5Mn+KHn+cjU9djDP9CN1vRiuxuv9+biwF8sTyL4
DGXSsG8Z5L5OIX0BibdsGVhAPpAgonFHEqak3irXebpCxRh4sZAbcax1CvFPUH5UK0gaaD8AMJF1
I7NPBXkkK3fxGOK4pLcHkvyBt84iHUA4duF7WNeO0WAzsukF/z8wVpZniAWBHkEfS0bvgNwXTfcM
s21gD/r97zB86Pm79EnIV2pIe389bTEGS6W/rHtGIMCNmSz5HI198Qgaf9XRSddHt/9ShJaMjDKl
bK+mT2XFcpFxIiNJk5WujwSLiDJ55/5T1r7JgUR7aQVxuo0pdP3MORapPQi5LPSUuqUdGstrzr5j
zWd/UdVAWaoxlCD5+genJCIOyOKPyCJfQTM7bxenRGnNKhDaJmq0uneM5Shjpot1sfamdhdNjvc4
wsev8d1e53v8W6iDVGJA2QoN9ZchZrTDX8BdlGac6h+uU8oWuIiolQenMwfrjQYrLDxGSFXRiQtV
rotuL8NkqI/qVB3dF0Mg9/E5kNLO1z5x+I0KA7zLZgTJUfL2zNRX1btfRKXdsGKiEBu487wA6Ugk
c1lRqHuHXTsVto4Yp49dlKByQb8UcC1UTFLTt+b6VjZLe8Ovdgkxp9KB5eJE/SIIFdcd9tqEauSL
wDomuEuFMH2+ZAFoBK5IGKboHp1DXd7kbQrbTOOHHrLhlU9gdhAxM3WVFtwfzSBRFNjBijufJgQp
I8HYD8Rm5CFC5BP0QZeeOc/AZnHHkIQ3kRTfO1B+fDqHPsozq46SpcQKQS1xg4RkVGvJUq5qtvua
4FHlCGAGh2L9rFMmjgMlbXErj5B6Cw3vvdmoqcOdwkzDoyCeHI3JCrd9hWGckI6ogmCQT7lMDK5G
i0JktVm/w6fuzbrZI9olLWrsf0YONIowUN+5kyQg98ajzTitXcpAwkkjsi06hf4IPaeu/a/x1EZz
8zB6CtJV1KqA91JQx4pMuGIRMiKrUYDEDEOvR159LBFCiux6PisA7mJOgzaStaA1MM8cGqhBfDoV
ndKqU2a7a0SlamXLF0MrdnSXJahpTaxSUzAbbuYZevoJ+kJuIlF/LotzspKAPMY2xKc5sC8HT0QD
v3kvoYcjJTmKKSH4lrErXKme1CiYPW0vNJnioOSndU9Sq5YuOvL1sw0i1dDpVRhybRnQ/iE9Kd8x
w17NxweXRaXiMByPH8bTLEbu03bttx0D4V+dA/3W6FyskFUr4maN9Sxlx4eSpRX5otkdTuo5Ejiv
e+HbghQla7YUdpGeOlNsqwfkecgeggaXD2ZFC9lEPOAT0DeG6P7VBFtitmmzvEkwdVHEnQAZ8AMf
ZFVv9HVz4a78DkfWlQ11NgkSCZivbZF2s7961iYQ6fo5YqI0OOmfUqeHtxnWxKCxSGvfxU7VKMa8
mHifpYOJLT6c51LqX4BE8oxMiSLYog2xERhZP1pnjgDBjA22pgoz6T6zTZo90pPxM7IpnhQS5Ik6
8oNzfpZZM+RPfjMtNQIxlrunRpphj1+FhAXMFWN5wC+xtzshQ0LNx13LciLOpDjOJcqZ3D/kIgVs
Y0OWyvXSZti7CBiYDoekwYAaFqwo3qMBxdORDxuwhxBPh1FDp89fhTvcqzBh3yyUQEaviYsB9aOi
P6UEcqgxc1TcOpoz/0MgcPObb57RxX4enm7u1Pbe0ef3Y6ausoZYLR2T3X53ANZ199lTzqvgNLhv
eLcbpiwEzpJqk8p0rjsauX12947BNscCn8XEt7u76wgOsJfdWimR/+lIM4YiI8LNJETe16/LpuV2
+QXnhSFZr1VX2fCzNKphdyFMSo4nNlxvP5bP1paP/nmU8bmbvWIt7gFPk1jJCO1qtepc9GL0ILvS
rgX6WH7BcaRhiAgDmqggGjY9JBAPw1cYEtMQ7dwN6gapsT/gKe77HRvILKVupz4sNoUnTca+twla
uzwdG90hoKsNgNJ7WrA0zVIAAW4f9+kZP1vZ2tFnhak+55j0tgtKekj7Nz+dob48iQW92KyRMLIO
mhraM6k90R9EG7JlTXbD9DiHxdc05RmYzaSTN6gr0SUsViCLK6La6D0YgNYM0NzTen+M6oOxgROq
lxO3jeiCU9JDGblxMttAJcHvK9rWV/P6MMMhV/DOXES5Mw9dJKIHdtq19nIdck37WyrNP2ax6kUm
X2bDc7lCmMf6qeZZplFFvqaT2WJvYbF4U4OzwoUTmmdktKjiDRwnj5tYpZuSKHCeeOLBnBxCfBlx
XGOwF8xmcxCGD+QAiPNgCor/HD8XYeIcsVefBUlHaD8yjsQQbruN8mm4UxSzINUNWe4XvMPAcRXc
lCqtsVx6BI0F0XV8aGDepqxWTLr6DyzFla9hxJNCrgaRcXKdl1hn+LL7/BbXx8HuxKLnM0Pgu9DD
J9NkuL9OFcKEXLE0UFPZM6DPHc4dVis7WtTMNloSmeostbdUH9QaiqlA091U0QLCjTX9QRH/Jfwv
nnyouCmm2kuzTG6/LEjp1/7jMnMpGvuhXvJLdeQt5s1lW6Ox2Ugr+ICs53OEzb3AAzYQMUeF2l6l
9uTV84Mf+BAJ+pu8Shkk9u98Ku/vji9Zoc5daqwfHofwtFZNDkLaObxhoMlkJ4z2loOplvwcjIvp
ddfoNI37MDajsz5cH2DxiW/zZpez3RH1ljgrYCwkFgPBFZ4ycBTZ4bBbXgYhde9wX4T5Z4Lb/sl0
SMCk1hTaya515XYP32kUNYyoHljomYshTiqLqIvGsf8Vtbo720crsu1E203Xr0nw0HE/PtdJnH9I
S77XXjUx7S/dHJES2LpkG9X7fbSiWvX3n1QirsThYSLmdYB5l1r7a0qmuISgX9QuLAcmfvPTPot5
Tfhx47PRIKLorbwLlBJQxIolCjUeyMuSqZvqSx0jzL6wKtbfM4FemY7uvxft6MyB3kBXsgLIpSC4
IO3E+rjlTASvVTFqT7N8mXmveEsGgymgIpqOm6iL58Sb+WfbsAevGwOLcYoNluWcOeUerr7DjL0f
YwjeZweEIctRWN13kiH7J0HUbNdWdK+A4LlOHbo4mG6oztqhJPmIayTFFBYJXXuwntQchnpLvk3E
XyLWj/TvmRO95PAWDSrnTyPnGif7A7txEx3Owpe1ZCTazuVRg4Hx6mLYSWCYCBd8PPAFobfLmZTD
QADDSkcLwEvEOExHeNkgYsTLgbVFZHPyMHG1C7n7YWfTiQfnAurhPpmgkjFA2968LSSqyghbwvsY
fo8ekPfLJsmQEYRUSXCoEhQf2DXNTZcxLlGuaussUcDGTveOwGeqEJOmuYl4FD2OAUW3L/JstSYL
Jr1fPDyHWsamoZtalUBMZ9c/yXtvCxtdsCVKriayv/nT06OlSkn0nmfo8TO9ekvsIEoUs4KgA1q2
L3lpmjFvfhJTPnfiF6MEZyaY7gXEenFZJFqZpsk1rwf0t+eTVHriJlDG/SpCmGSZ4wOu0c2VzJq5
rNmpn49AMt0hOHhGAh6bZ337lU2x9cyMno3hfI4v6RGnKIuEmj7oIEXO9e9FqAckGfvlKfOULNUn
tEngL16Yfanfnhmjc1ksuw/uWE9PGYAdnQ0Yc5c8tySs7fkdLqbbGmLacGfB074qkeKNy+Mahd10
F4S7RwnVErnxv3ilpdcDfM6V0eRaqQWExDPfSnKDeFASa5o9bvcdr6P3M5oQhdIUnrZ7zKm9i/+v
G0SN+doAPKO2++UITGjO1zxW+vPKXmqhtBwrc/pwbdnOQpewIXztG7JknhKd/zbuDQqn+CYQYCs7
7Qarx3YeZatnPaYK7ckrIOTWvvRYYiRz3MdQ8w9ODP8iQZeiqfpMqRuvMu2ogLHfduxGqIANh92G
2PznXmGxfd+vky6LglIKZx+cXXFz3+e9BxG5RtURqK5pRxIt1YVHy/FX91Ocen0j/SLb9EOZEN6G
3uGgX3imWNoabpUUxf4RxviYjK3pwrhh9DRzjT/nwGXWE+bzGvGnXFAgf7SOrj7iTF5JWU+te/xY
Ityr9QCln820CAY6LCFuSyH5p4v5GatSWupY1jld/ipt5qcXxLWYQrhfgsuQ3pLYrS2RAuhWjTZL
pxSMc3QCqWoyw8s0xOucuxMa8s3skdFp0asA1wszwBew3EI638+guha+Wwy/61UuGdEFA7Z+m7t5
UuC/4xNISzA85AYaCcyiAdf2T4aENdSyXs50XnNV7eHTEi+G1ZSO9zz1bKS4U5micw0yI61iUkhK
8uAiCW4iXXscIjkvCzb0/2Ttb4rYm1UyTxgnjdUHkMD8PexYE8aBbyTC3/b27mNGZFW9e+Y/aD6K
atV+4VRmEpcFgStEH9v+gidluRCzM2xR1t+WnCh+HR+4EQD6fnmLIU61e3tXt6ssj4luKzO5htUF
tlOSM5WDwN1yexZnPEVD/Ae5u8dOb5mJ4u6/FyJDvI4ApYqM3kBgUngwl1qCk2nMYd+FsdonTb2j
S3gPcIGwvONnrzhHnYafhXe+3Ev1SP0gVWWVGYbTFELRBj3rY7lUNS1eVbjHMQiEKnb7ZJtTVEKQ
X2kRAsb+XmEpdtovSKvgfwjMwnXQB6h58TOHeu1KpB2SBCYcnVH0u482m4fv2MTiU6EOIOhpnh8p
/y7RreVMEPXrT+0dV+BNDr1zCHoLu99n+L/UEm1V7MptAZzQ1vLEJ8FDwgURKRGUWXZY7BXK0b65
6PpOVDDdZEeJmw6AMpfaEYJluEz1JNwT0xDZPTRxk9GOLzeikLMoi50q3tZKqdi6eh8LXkaDNH9/
K5qzjkdCSQM+y6D+vwGCpuhpsdQCb5NpyzjPOxIFhzUaxCfr0+Hw8xmsn8INofXcB+0/sqUNa1eR
HquCJ9ZUxBP6NtdAo1QKrx+g+ZNKuAXOxu1J0vDcU4e7udVgRY5k77fbfv7WaYlKKuhMNmGYDk0E
MiH42fgqKqanLeBENTvzM6n46Wymi1+7UntewaB5/0K9sJVec5QPVh7/Iaw3boY0KOOTyNinvvWD
XRoE8WBL1C/dn7W99sK+6VKuEMlWHbqBvckCmB+V/6YuPRGlAXVAeZvljLypbUDde4mvTKGdDOE9
tcJwv1wn+ajwcHqvwu4avselnVeX6PLXwtpZ3uI+TRuCA6Ei9EugnbCNEdRzoA+PwAkEsj6toayR
wBhcNJ7g3V1jGcN/q79km7sAUjvbTnV+j6Uff2wjrxsjdStFtYaFzKBBvwViaeeoVA2TTakuy3Oz
O6IGtUVKzXG5K8zfIUdoVwKvfrvBfgBac8qPwnEzi0VI6OU5oHC5NKs0Zhd2JoiJJY/0HYpNuVD8
7rSCJELtgEZFN5dm7NzPL0od5417cnW2O8kNj88PoTlj76SrlKzOjeri1Y9NL7u3YXmunFMuWRbG
Yw0lMSeXTtXQ/12pAQfHgdd+MsRLPYePiKV7+wOlxGf1L2ILYR+jk0iD9Tt4GmgirrMWDsguRzuC
3P+tdxls8Ed6cMh20SR/VBqNSY5uwE7QY3jRxuNtvuwNRdpz3Zgo7rtcVRpwpzwwPXfSEcmfisO5
+DoRA8rTdgsRRdBPUXTu5zL2V7yHgxPQ7rLQam7Zet7iyixUBpFaRCqmG+ds95Ghezc1OQTLSlgY
CHl0AaFRPFAs+Df56I7YrrEwaAkY7fRTcrLYWeytuAVdNJUfsY7fIy1arjbPXB9cA2HoUnDauYxd
McGQPF1y0OFvw0jgsS0GRtJrzovJSPHlUIiCj9+9NTss+dQHhd5Y3K+0DNPHcW/Ea0bepi4fXXX6
G5W+HLECCsI2qQk/UISN6dAIJWpgxWIZ2vFpSmngJliyf/PbGqZ+uMg3SaoisBmcpoBeufyeRmDo
WmnpqlbLujsVQa8hTZ6QbO1zEkRpnzc5gldWpy2r8eYFYKdTQMiNiQjERJuF1CbyLy8M3ouBBM8w
FrpRTzxOiFDp+6S4Rafwq12RVFaD1SXCU+IDPVx6la7E1vAZmBw8/Qbl8R1Fd+obO9fS1STUu5yA
vr8Xz5nbd2sRsfNWU1jilbKiL1vghYNxH048jnxM4dFuj2OXUAOw5N/6RvjCmh0s3XOwB00PmcPl
XL1i5gdoT28RbLDQwagpVEbM84jSFPyAjhHswHqpNK8W/mKWH/WeoHhCuVsCsy8RLEQNXo3g7LaR
56tpAKm5NTuN+GAFkRxuk4iio6QL9Ywg8f3G1bXeN6HQzKoxzL2veIi9aMsCoXHIjvVZ2lKlR8wE
E0zLJ47bjQ/HX/z8CG1u3koH6eBxlnNii78UZOkvuFIsXO94fo/xYCqd2bHha0i+XNx9i0zRgl/a
v45TUzcOlDFdAAyb2e3PJL41uNqnWMXJVUTfqjUA7HonWvET+1Bi7D9QncPZ0q/G9nF6l6U9eHkA
r0gJzibePhB3aVLstPTAnZc+RFcaHCSZLclnyW5SXV9RgodkMmk2yHPyr72MiKak19MwCuzYZEuR
PLAgvnDx+dZMURD8NEvD0oDcvTQRCwuk4tihdHB7iIaWUyvnNUbKaSJQ8qocy3RJefafk/s/WiZa
pmxrhGvh6EuBgD/hh5FO88MEXu2SLfTNUBMoZIhS/95mI6nHTqzPZzFKM09g6mFxl26eiYfGwuRF
5F1f/DrHiXSnmTtxLWesJrj0Y8yk9BptcQXEyXKh9AYgLADj0J+LW+g6aEUeiydcg8LnxZRQPrnJ
0jiY38Xj16uSWnDIVTXSM4FK7PMSNSSoIbeNoKSjx5q3YeiRPAONrUWaO9VcsWOWfumKZfSvvskd
/wF6pzLmr0VDP8s2nVoh6+MQTN8kJHBk3tqmyRflsg1nXu54SJjQGmUPPWQZ3xx4sMT0oWBydRVB
m7yy1yG0zy6v2LjFww7Xj7k143c0wv7a+7Fwtdv131fz17KhOoQr3uhHtnRDII5QvYpzSBzFtpdN
exRsZtUNnd9AGu6pC3X0vKGEd7Y4O5thP+cuM0a+gZbE42ewXJ+VuSacusPiTyhygdWvNH/M10N3
TTXZOMzFmH6swsc9TXnxi3ksDK7M46YygaLnhIzSVPqKDuPgFGe31ZFnX9Oy2xpQhNJZ1jy4atkq
4UPnERiOUMy9cbY7eb4wq9j2UU9UnkQ5EQcbmchYjd9bCw+J0s1EgYHlaRF3+nJkR703bMHGlmFE
ioWp+Ek0TvMP9LsCjgruyS46r7Ehynu6iHLxdOOgNvfIS6Qbi7oUEn1YW2B07lAKMc6CRjltt1Mr
cS+XHAotAMN7mHJGSpH7RN8SWWWP9pRI0sqRPhSTKdSuBB8FaQoGZiC/LSECaCx2wnGripHdW006
jY43xTDb0E9NaZpSsbTTOIxy327U5Emfi4EZ7l3RTQZOTnPbfsydkCd4L+dfLtTZHBUiz21y5uyB
J0C2XAQnZbQba6JD5sDMOHLqtNHiK15mkzmWYcmfR+ZFAvCG+ivFGZ00IKeG31puBLN5WQ5JEe9H
fSz6VuJx4+MpCicFXnnGFV4/MG0N8DzVMvVowMXc2gUxbwfNQ2k8vuJfvkJbMiDeNoIuFo3OEtFZ
Gk5i9KbZusuTW3GeIildY8niWglD3Mg3LZ8FzE9QdJ5HHoclPkRDhc5uwjii2HY4RiLOhjyQKpOt
cvN0wKzUirH9PlA92ps2ImYKc1sAbn514todN8tjZJKyIiFcB+70T90iY4fuDhbsNNM+yH3mOZL7
SyBO3hV1pnRONQEKpBiYB50Gh+3Hfd6Z26EfkCZjd6nghn5T0o5K7hsg5tZ9bzyLghDW32UPVbkQ
CGV+aHqdjEjcl5eBKvbBnR5NOOWF5rvS6mzn7XTU1MHcC3Lk1dAezNjdO8RD7dmcPmyDYTWi8UvK
lqdZpO63d5qBfjBGeL4ijo5+lVN87+qKubfP+GhH+Lh86Vxxe+4QvusOC+wXIbX/+IZW2eQJTKfj
zq2lfkQ7vWbSvFJBJinLEf8za/6WAD5f13/uf2LhOVmVZ8qKPBiBW67Ut14IhyxzaoYYXAaQ0Nss
z0PiNy8RnJ2KeuAbC96kF7Zk5bKifmqlZeJKwgLCRoGkw5IV9oJkWc2AtemBV0BbJNpx0M0fUJZk
MK/iCLVsFWTLmqFOdM4RguS6MRfVm3gTVdpj4NinLFKn8te/DltlIp2sceaQSWCc7c1kQdpmTa4s
AeqdcJEMVwRxpKCgPupCyoP22C5IK8PxrWJfB6eGFm6NqV6yHjWwSiJchVs12aKciNMbjrwr44VE
Vm6gS4QOoSXSv37I40BPejYG2BASlMDrunP4lJlzAqtWDhhyxjdvwuhDzOLDsvLjYG0nySLg3rT8
5OacHUn6iSA3X5WXL6TkZX2vMZmHj+8XvaU8KPmf/3toIMQTAlGcZbVXcuQa3ygYDkfog2msXgfG
El+xJ9qwF8/z3krB3KHzJfLJ7Ryw/qMuqIfaqVVGjMMnuvhnuhiBOOi9keaI5Kxuyv19CZFgIu0M
Ul6jErJ8rH2vN4Gf6z759NDgXEMyXdDwaoMZrzLuUjjRNaiF9xOWOLY0ND4ga3aGwBApNWlXbEc4
OUXgXXQbWK4QVBYkCivW3+vcbtiIodDN1wQZ1LMs2/b5VdFHGczuLRD0q/FZj7ilDJPlzziaYG/q
p1EwnvyHBTBeQBl3z042JwcNJ+uQH0AMr8h74u3F7LiYEP1GYjKiJ9RVOeO74KAI0JgjoPhB4ijY
0+LwfhemZYNru+yxE5CD7dH+WFYo+XnHmcHSitP6s8hJM3iPgkXqb9OfWNvfSy/PZ2wBVkbVEgQe
gWgBCvoYfx/bBIN75wrtklzIat8kwvyO8YoGORJxIWxNqaUDCe2sy2mnHTddDaiy1mMfW+I0Xr8A
h7J5Rua5mzw2nsRZRYiosiAo9XMlXxajPeYioYLYyw/zFGdHfhAfX6klFSHiEX4d66LAnITfF6EM
AhiVc52i1PIAFrDlGoEBjh982q6gejVs+yQaA6p+f9ZPs/6CBcAypmIHxou+V6tBrI+//Q0VKQiB
KI4EWlnmkkIuGwJ3BMFq8/4Oveo9CaUE5r5xIQ6np4/7kTxsg54YqUDSqpKD+Tsb64ObXlNqS9jk
uoApTmvzXCmwTKPXb+5xd5rtqWzGAFAETsRxsaeL8RLJ95nJHaIoDyiJ/ABATQt+uIjDFxgPZF4O
Vo7FoxkElYW+3P9gjsQYxqjC0Mmzi//aHIh57DGyWFgu3C7bA5QGphgXhx71WlTYWMV93UtG2jxY
PfMe7ae9mGmfMKpwunFVGMLDFfU7wBLiE1PwWARW0TNNQR+KlAbU4enAasMwrqowIsZMNYB6GEKx
8OhXV9vOv0N/cKzB0tVYgF6slVbXa7Uv9PGKbLZ/ua7Nj9dE9wuZyI8xHCn/Shjw8DUZTLoWJzCZ
KxLhwROiWBLE1ReXhZ3/J30w9HQ0Hs86U3d0tjeXNWPb6dkRe/iO5DJsZX+EIirmB7puCgrr6deB
xK5Pm02GPzn2LrYbOmqKzcpvJ9+W76lyOz1vylFPpxSMV3UmWoCmNqanafMIIqk3AVz6cIY6HtaH
rneyKW5MjVTcwMerqi8qBiaR/u2bI32m+EE3v+0ew70a0iiHGZSCnaRI/jrgje9NCmswZ38y4ruY
3vTnCkVsfLNt4sTn5G3Dtv3wiEc31o/Q6jo2f0IPIg8917MuN6Jk47PqzQW+W7nUyoCGbiHm7y85
nSO/GyyjcNFWp6cbLkUrb55F5wICtddC8SvqZNKYF/rFEMMenM0CvBQ7RrlAEktccpvuO77xqvO2
TDt0MQepll15fRcP0q6hypbXdTg3FJq++wRIZMznvhxqGQzoTPXb+dardHvQcf5Upt6G0iLNj2Hx
0sFNso6IGfDnAT/r5EJa0Xg/mQLKzQjGXhZ14dXT5dI89LeHnicTYVj0AH8qkR7zwVr59KhgW4wR
yiMSg21515M/YTFwBH3gUe3ER5ABnl5ROLjKhEtaBYFBu4S4zBDImBuW97w7HqMJKS3x2VARCfg3
4eGpXZfXHuW8PYY3Y62m+hdeCWrgP6uZtbBvakzStaQ7o7vLys1qZs410CC4xuSx3d+hIP44JGlJ
hgWprI2JZQ41MGSms+M3ZzjPeEtd6VRWTyLcAhgZyBW3fk3dB7zHTrAvGXzdo+nDtIxslc6/XIqa
De+HNWd5we5JCBA7sdYWeftJPu2Cm4VyZ5BgTQUOGGPCNPd70s1K4DxamOygmM9/6RhYXDu4QZso
OQUGgSZ/Y1cU5ySdG8GKKJED9iCTdaj6rry2I2Cbx54BQzyNwlBI1d79AuyJQufdx7KKc/u4vRi4
9OX/sf7ygR2VhxHCnH/Mkbx4dxjnHWjUoa93FR7mbPyeIF4jg2Z4hcmPmzzVewLoIqfWVbAFV0w+
QljCOZHWegwnpSLfXo+RclOCdrPscXMJtSl0LQTx4Ye9LQETqLJrm52DaDM9Jj1Zm/fOiG/cofj0
38dxLKiJ3hcDTwLh8uLUpcvOY5E3eZ6Do01nt0bml9lPGCLt68maLHKVvelmJ03aJHNGbcpNTfVp
Zi6fvN44FPRtaFcaDmDlMGx3Cc1TfZb7PT9i6Xl1EawBEqKm5sUXtYXPV4TwXqx8G7kej9ZN+h0C
r57BUeY7lrWmmajqtrYoX4i9SeAkIASkWqZ1VhB8U4Q6+duuLHIjfeBiKGI+TM32GowkWOkaiFq4
av0EndkLxMZn9S+VAtD6LqLyZXWsal+XRJCvKOF+IzoATXeMTZXIjMJKMFxPZCyQB29QXL+QcVn5
0nZlDYm1kM3rVGCA0Qou896QItVvMs2LcBiNq7VYthgMVrQc2JY3bGej6D+veIVfJE19RgbllBOo
Kx6g96bdrs2zRXH4ewde3P5bS5jetfEzN5sgqi4nWnRWzNcdlfuURnxngdD1WOtHbYOTJqeE4tMC
0azYvlueXkPE9JlIIVtiUQUvgliOaLfLsaVeOF1lhfA3t9M9C2mQdaTJZeFhsMnNm3XB4oJL+iob
teJwPJIUgnIVnt/N/KVShlV3Llh/ZMDIO1SZ4eJjK3FYjwas4ttYu6b2fF2m6vWer4YXoJb3EQHw
jUeW0S3UdlIvtRgai1lasJWR25GEVju0IL73iJPbsFv9fscpFdB+4ENhxN7AsS/yrxnyDQBj6Nkw
E4a3D7Wnft4qKlrXR4ICigCCvuCaJS9Q+59TYmngPm5gzfM+uJFKCE28w3NNCC7zRX/DapCNp821
/i3IkUPxbsJ+AaormXK++77rXyYOryhYT3hbQjUj13i9iNa1aiVYU6gtFRA142cwpNM9cxIHjr2B
sW2B5eGok9xK56Rj7Xe0yMUZSTnMjeKvSzJKSgxAhcbRD7YPb+AhAUanx8JZlu/kML6vqgLo2/wd
dA64bO47cKUpW6w6ZTtHV+M5Hh3uKzjIgpdtStQf3kaPnV9MZwAxydtH/akfc+9BrAqijEsHvFjM
Wy0hOfC6q1FGoVbnl7FkshKKx3c0gwhARXErUnNzAa6SpZkyssBOk36J8p3pfFyDvZL/Mgc3wi6r
3GV1YFxRzUn6I0wBGEh/1dPj44ji+trJ5WK/WQdPFwOw/fAcbBYVAPdp79mwj5+fUXYYRDZzjiHz
WkRBtkAA2bXipzzo0NVet+R24k6lLm6adZQbmkU4zhpyzL2SVr0LK6uSB5WJ1FOQlmnJJaozWqoZ
Kp//Jxi6JGwvmR+C+h657YfKz4FWbwxW6NrsTkHQynFhKsro4WGE7lrP0WLSbnXOEH/ec2GSpXbl
NjMIWpSI8QcUwDwkE0BN2nfCH0fBbus/lF41AhKln9hwL/VsytAAqdpNpM+ikaZotOYNUmVd5V1s
PbSJgnuTLoESUTCXkQYtZeoKoOtkZ6sxfG/pZBSptDsdDQNzEP2vf8zJJ2ULwJzGXGxfQcwisU15
p2mIGr2VEQe9VfKa5/6GqIRzuMw/lz4p6Bx7x2yrg6FwSHsqbzPrOTiPGm+4J0DlzH2oaiTilGlK
Gbb0oG3SlqhMTH0o5mqUpaodgBOV4F1iZgN6snx+Kv6LAskygF/pFQWJCav8QnxqZ5xBeGYsPu6d
NfuiphiZwLvjA4Xrl+Nm6VYc3n5HpMKvXiS+HAB+6A9yWiZzNCdi+nB9i5Gn+tjQ0p6Ht5j4u/jz
y1z8Z9APMqbZJqS7aTNHnkLoor2gl4W0cnuVWSTQnr1LZJ64uMfOg6fOJYB9zxFUHAmmaCXa2ZWN
/05k3vd7ydAWAV4HEY4M8dWUgiX+2/XojA78597RG94/Y4yokk9+v1FFwI0hW3/V4lB772+S68jp
Wsqs4CG8uJcQxhAMSFYj96ABUUay8xeUwq5OBexlvbLgqZRptjDxYgSJ/T/lxzZ50mtDSHTtbBvX
zL63cDhEvmjeNvBo3dMVwZR5EHWwTTcrU8/m4g6dvkpBjs43baNYmQBc0kph9zr+z/h3IkylT/md
IQwmex+7ENoKex42Ahvl0BGBGFDakoDlSWYLjg9UTN/S3c06U60d5PoTcBM7uRNXffQF4lWGOkVS
bP9GJkjRWPvFmwY2zhg0FgZ0OCBczvkyjxY7KvGWvvK6WU9GqI6LXtepujgyq9tAUQ0EcTcyfcyh
L8PiUtLfsRRCj5Fe6JgEry53pfx4MWnAoppC+dy1tnGspTiZtymbjFHT+RLUUifuJPh3k+Y5YHsi
64gI5JUBK8ty3JnJXrIBOtreO+tS7XdOk8pRdjsLos+dldhke5WrpE+8HjffRUQJmAskGSAsgete
i5g1vdevxyER1C4gpbupH6PU6UwfO2OCSsMGRtSrLjud4mzV0MsZFDfaOuRpTBztHNJfHEesH288
tPE6lZj2PwgaO9Pttq4jh71iN1UvsRnC18wrvQl2knhUTvovLkH6dRl7HWDfzFGBREaJ3WsIU+We
oAaKcj/bkWmk2h7Zt9BBbWO+dggIqLHqMu5LYCptaGdDfWuLn5oZOSu+c+hjZ225L+gVcQnquOkV
sLowZUTkWsWrC/qElogxAGBT6HBi6zzKJmsAjNQOwn6KZP4Tzx//BiN+r/hkUdiBITS0N3kkzD/s
HNSAnglgjgTHTERIKOdYpu7oduK4fh57p0PDdi+7JMgpz1Lp0N8cE2Gufadhc4vsuX2CqTdQA2zU
+FwhfQvFruw8gLlN0FL+GDKxeEU4kXEhl6yIy0vOli5n5aWQLi05VE3qrOVWic2XKVKXZpBfw156
4niAR44m8QdEYM1W851SKMsvdy+cKdDNwH5dTLs9Vu8YLUq7FTc/vTfvFun/m2gKSfeqAu/OTyLE
cldD1c9ZjaVg6wx2xLmhsL+G93xHZelFxVFI4MVgywZr4OxJd0iHxrCeNQ4AjNxHOjQNVKaei2Fn
5u7x/2SWy0nqGxJ7u1PhawD8rNCVnGmnoCpXTdOH/STyoXCjW5EMrRnXkORXaxmlrNglAEttFSdN
0wjAPRwszJ9EbS78AgUlIaZxOUdg/IiDiWkC1nQsoEjNNKmVBkXZ80HMZlc+mxe46tziiH6GxRoL
nVCwF55/vSQjttAhFR1JMP92Ar2Eu9yHs026VHht0uwH1QFP3SYE1YLdWsbinTu1WQjr33fbZZ2k
WV3YD+hxvOWVhAucBAoWE4wax3Z966O1dSqYNzHffQ57x3RyJhICrPbECQ3jENWvJKboHFA09JGT
3QDe6M5U2ENAKPYCnSim3o8fUHMQQHmRXvalxYsZCGri08D4achHRE+kRHlEqNJHRU0dQne8cV/k
biCHD+cvKJpXnM8y9qmJK7mhDcWZ+VzvsXnGWRr4umd45aOrh0khnNHKyqZSBCB6DXSCRmKnic35
AcEtDbsNSAgzifonelymj5DYZ4htLXw94edDlpJVfCFpUMWv5YlhLiljVu13bnW9SuUGkZ7H7y8o
8Gi0uanos6bXb+qkOO6CE0/tO4BuQQslXvAlbIv1mKaA76qYwC32KpBg2f1hZjpy/VYySHU1lKAb
LBbUqjvQZe6gZ1lslLzinxgjA5vw9bqdRe1Ou+d1FNdPS9rifHWdl7O2iKt6zy6CgT2BT4MoTYSg
dkbnZIB/6ZXfRwicC3+OV6/8khE7zQ5CYIBVHLLloEISU0BrNWH4g6QQ4URJwADm8b0381nnT5Q0
EvYwCVpxAwcMynQ+3ssHXnQ6h86ToJPE2V+sxt7YPnRhtkbZl7ZdXbD7YsxLUTO3d08/ZBo8gBF0
WoG2kIicLVWc/1PLsO8KihaRxoW4DCuGgeOKUsz7dxvdOJ/o8YEw/gA61yX0u1kObL0IhyZszLBk
Nm+ZaMNI7a11IUxW9Gu7mW6p8/7tcjZIE/2GvCgO3CGryIf8VKR4FWIwqlsQ29PCRSo4MWmMJxIn
XLAmlhBjez7+YgznfFO8ODTBrfg+uWlt4uXZPdGrY3Hq9vuvveHb9Xeyls2KRhdk1qGVMvhVKQp7
RGRFhuUg0gcdM10CPeoWufAw/4YsH3+myfH2ek8Rl8fA/xvTPeSTej1pB72i93A8qXiswb05qo7x
ryvthWrsXZTZZUthGR9hGR39ueeWQ6ZF47/HWeGQt1xMkY/W0XoRf7wFiXZk1NOCF8KcO1hZT1Ne
OYDqOBVTyVT1UQ2Lhoj8f242KkboA+aB1IT/iQKj+YzQazxhVtkdEPBXWo242SLAaBdjnxyNmPmk
VD0XIFcatBrHlVn8gHw1OnRCw3ZA/FfI4AG+a/Fal8OqOv1qL8dG4Mso8R4GGGXxS+0KaXbcMiop
XYMEG/JjMRtcTVEQ8ituYWkJbyAQny6gdyWhE4USw+7HJzppFLFZriZE3W/mlPPMSuf9VAkwrBiG
DB2A59L5/d6a0v2/dvsx3Gs1DC30rbZ0ovgfBIakWjBM0kh9alB8mmsMtbrvCiRRhIFwbmo5203A
//1SaWBpCjbefujBygvVBFSUHWmZNUX5caoMoESIUm2pSmXwyHD+HUkMF9bQSFU5CrwqNA1Eh0/N
L+mos10f8e5ps1lRKM30RE+8xpJqI+Terms6RBsRzq6V6xEae5dVnCtHH0uZEEatOK7iYdtQJ8cA
Hl2AqPpDGAr9/z86t1MbfvsAaE3Vla9+EVrlDROV7vTLqCayHey5IBhYcWSVC+ucSXg4YdS9x5P9
64zLqMgc6+sall1Ac9XIZQpxuguCdk0KdYBXTsuXwLxUEzXKXIi+CSqBxw5bbVbrBTn7XI9qmdXL
bbmlNVzyziZBdbNK4PAuRqoCEorNfuaXErgQqijE8BpcGpl7BdEUc13YZJG5rb00D7dJl4vLL1g5
TC45TUXm/MBBSxm2RKNCyUGfYV9eB/o214gEVZigKzsm6ryEz0vPZfx8teseuMEefnU9zlPcW4O9
DYz8uCEof5aYCwnaym7NCqsC+VzwdmRttmtN/HgMV5kB/Wkx2Sjy8Xbe2zN6GATyMekIkyyVgyAy
WLqmTzHZAYVQeR2+Hp82RKMNR+a0Ke7MrfbMI0f6sK3FP4Yfta93qQIYF2BkDEopjXryK9EEAnoE
aNI+35zbEzksz+44WRKAFWaKaX2Tyq+rx1Dj0bPvTijfhyBRsDJn53GT66o6l2tPKHxSADpt9uBi
UOQfBmZ0MFM350hyqAYrGA8fM23omeAEdV19MHDzXVAw5wNqFIj12SFwOZFS4cj+2nAIqFkYlGKZ
3LGV7lYU6F1VZwaKpR5l/GFIgk3jrAKyaok8hk8oxE3R9z9KvVPkTfgCJgN0q2bdv1nnuSLuWJHi
fvWtD/Z/qJIJQk2YKYg332M82VtB4bR0YUBTRVHBOHxf4VL+01XN3L3B7ObNQmKeuwkQ6VhomXih
xhwvsve1LbI2pqhMbdk/9PaQlDDZyGNo5r0mDwz+6Imzqe+AGoXWCg+Wn1wOq/hMOQhGH3CSpDrT
smsB3OmEVVlgBqTU7rBMx0y9zY+KiratTIexBnpYzitOp1NmmyuvCfLgtu8lwoJQXTgj0Gg48qva
t5nisJm76jl/+ldUOHTnDaXMJQOZ07QGDhcW9VP1EpffwOPsynZa6lSpERF/p3rff/RqzwMPwPrH
EXQyi6yzSteDxqyMNXBE6R2SPBmVyg9Pqp5a1mJV6czAen60aaS2AdX7lvKJmceA2l6ydh5QhWXX
d5T9EpqF5xQHOwkClLqO1G4kYU/nWrR097GAsd1DrvI5LuEGPoQG1pkjxJlv9zQJ3cRAOklT0gPt
sXLsyORdGzC8eyllKRBPU96wp2zxNCzeX3idbJarQtXz6CA+rSqrY/vwo8uvLPjlYDWNQ0K7RPiV
EG2mHcFuGZwHPdbTTuKRCyfbQRI0uWN+6CfSwMF43GogzkOufmCnOI2snRB+mhMXarF0YYFH2GJ1
bhW6hUoYWGTSwjsIHtAcKolKBhbZdmcxYs61nloKs7zCQczp+W0uk5uawO9nOaphAtIasBjAUE3z
QKQViwLNamxg74YjBO47cp80LUmHpOtxlhNAJahNBtplpBDC2Proz9Xtc29hYmG0b+d8eDtd/aw/
D/6wjPgP0/N8PWLZfB/hWlhGE6WmDvS3h5HTFHUceKKI5/XZNoKJ/Iw8SZ43xyl38PXafVHvZn8m
hZiZTXyQRydTo1cW+wS4yNW3mFm5JBuhojZKfMBdXmsCSaabHSoxVq60t4ZgIQ77SPVQCQ75QCW8
m/0kyC9NqljdCvqQUBOCRi8k8/uoLaSJlI6+5twXhGRCatrbof2nTdRT1+LecnJ0XDEYo41ZkLn9
swLu1y92YwQfI1RInzOYDuFyfGQNcrXNPREzUs+AZZSDNDdISzo0OX+EU9sZL96N0rOkil5lWRnr
+7zvg955tgEWoKZ81RJ1toQLWmhHFGI9aQmAP3jE1nE3oMb7f0bq0hv8SkZO/4qjV0XAXbiIqjy1
y61EwZOrefTUu277Cm3ltyjaRAd2hDCHAVojCpgLhXS95F54H3ADo0nZJZcmFA2NCBpuSe9EPfGp
O7yyEnMA5i4CoYGhx6W5rMf1Ipud0+5YtDjMTkuAABxj8jsFPTTeciPc/O/lELQzEQw67ncqS9tn
EfUdJnW45z3DylH1kfOo1UUjBt8/P4iMWlkihxqjyP79Nvsu9cpkfIj5gHugh/LlTXaKmSMXdFan
uAAkBDdPrOXd0VWDwBbWmLMw3UDp4nY8kRZtPrDlD0pphae8pJfkKXWAQ9/n2sKwAlxZmZ2sNCZ2
/pJfA7q2erglAKgZ/hiIjHelr97+dq2J+1yWmqVkqQbsR3+wmM7RKRAlEas9OdWv9fsFDnbfJL9H
4EUHvrVPz0FQ8Yu3ZTBFdRMagsyloJEdWSSIyOiz2cOYn1i+67htNYVk9sJmw5bM0k8kz48XKI9Z
wmQtJv9cqZQHxQQsx5UOHJxkYj38hCtbqYrC5QFL/rDdgxTVelB1zjXzqP/1Ro3+WC3wZ0nCFMdH
bLp6HlGrNcHXyldX6S9++dGnVdpZmfuHu9XfZVneLHMiksi4WFZ69rbBSuZvFYw5uCQI1FJ/bAxd
Pw2++yIaWdGyP2eXElNLVNRhn9vJ1Za9ePQdDWXPAxgOKHPHEfIrRY2z8O7pHQE6q3qlLfegJrJf
FEDnhYucQw6i3m4RMOzSpFYjFKE1Pbo9rLlKfJ14FN/lO7k/6RctUrulYrha5/poRlPNNPm1ivgq
WUKdIqjs6YZ/jG5izMkB1rSMo00jaVtJEMlCdjPphNKKvuZNGR/q4ySpOYv2pScThUHBTLdw9uKV
Tr4notlOxOgGoU8rb5KVvPgZgjIBIBwx585XYKF7kGr8+YvteZ5Q4ln2IyqSuXb89ddoC1zNllYf
3DpKUKaGzCXP14i8cWdpNvdcgaONhjOL+61apLXOvWih8RtmBXadhMnOdtnjAW7s1TEKda0vWt+1
/ZSvF3DuePm3AK8GpT0YnxEJx/e8qRiVcB9cI2A516ahF3ZG/6+JeP2fIdPsDgPxMIKMeE/eG2UT
DsgWuzRklRkZMQMvXWe8qxk7WibxbhPajUys4s4t10sOXIfbnRM+R9b78M8xeGbkZJcSFOz9TxT9
3zc3KYx6DZSwHQ3dU6ScCtSTpAbTByRqKtMhM5Xo+IpFiAIHQk6+VnobfzOlrukIP5TFLk4j/MVM
6rzgvikatYv9RTXDim7umxDy6fn1C/qbwuLEvQRFNxCYvWR26QoD+z6WYZkuSqyEDlDkJD0Z39Ix
46M143b/vR53qgsajq9VwM+VbgMkm3qJSn2VYuq02eEgOvIu9vmym51a4hQJTDJuP5kPuQLTc75k
Y5HOL8N01THOYxvVSPZpLeU1oFMKlr/bUzRp44IhJl57LU2ldVzOLihJpeCg4J7TxpvjdWK8Cqz3
2scog1+tljFi/PhVsm3ksLdH+OVb85Xmm9H7pVdCr2h2Tq57v9iMi+uj3Z/UCNuOg71vEFQroH5D
jJSMQz8sQf98j1/s8wC1qbteYA/b9Ow6hkrREotVhT5Ud5kQhHyXrHjackVyJGIWFnlSHozYhDww
u791mlS7U333ZCi7aOQvgZgRXjPS4It+IpIlHap02kOdOMLc3JiMUPkZKsFW74oVqfnyl4tl6vp4
kaLoriYIlzxMHgBSpLfTArXp9cSrRqfPXf7ge4J6MaIOFv5K41SSrKtEZT23KZjIDXA+tsLdfhr+
zT1lFxOzjB2vse7+8kfa5RohE83m9ABAn5HPOHe88MSrgUlH6GmVcNIZmW80vZMyuArtwei4FEzh
Ur2pfa1DIW3HsjvT85TtnzRIMyENjERF73Is3Yy17nPZkmZ0aOif816B+Xo3OKfs5x7Zwpmc0jiS
q3eMsN/OXPwyXdrMcoSgC7rVmlSYdyU73jltcpHDv4qAKQ6z73eXy9NvtcNFMEgzDEriowWQ2fXf
cbntxJdLNVrKJfhgzJkhsJZfFReXRghGgV0jEFB7ya6kPrBxsEAG95nIic8vKUxrKEwEHxbHLj15
92A6sb76se3VB800vxG39Tt2+JxkjX5lC/sJKN2z1Ixb0nFdnhNqshXmG0FbAk39MgNSatfXnl0z
GCSMrjPAqodQYzF8eFmCY6AU6X4DdZDdSQxTEjPNX+YDOMyuXr4R6aWfLvHZxdDl++jTs6i83bWw
e2XgxlrT0/Gr/jVZlZ/oBFLDjAB3F5WI1dcNB+IYLz3g3lNdPbPdbVcCKwof2hmsj914TXCDF66s
ZiOVqVIVmgcaG3V0xbU/oXu2xJGKmXuLv4d0TMADPGJ0laBYbDwInRBw5GhS0f6uwH/qHz9RSa+G
2L4orHZrVwIMKJStNKNjybdH/1e6KMtWFgZH/bYGJ1JNrTmSnEY2EfNjLeeE7PRY98Z3qEVjU0gV
TkTXfni93yTewEt17yG/qM2LnI6TXThRktmURMd9RwcvckbhGfixeFsJK5Yl1tuAcrrP55rJf52l
3sO3abZDc/CheaLgeh041uGOYnDkda3/At+r1j+LgFXrws3lFjQyK8KCIamB2SXgveuGo9b47N96
q8AxWNk5JyF22Mk2Du1wzH8u3j2C9l/Mt8HWNcoLHuGdg1/5KmL19OVYL0TztDgeXpu61gsxv9Ng
/1cZ02l6o6WPafM5oPX0KkJ49MjFvG0jaWFJ9UnyuRoDEebJFMfcjLmA43yDNJyXfp+uDdrtvFOP
TEpke7enx4HUIEnj7CNxDAQVTA4Q8nunJt/X7IgiqDWxMFj2qMw1f9hZQS52ffYf/BzxYbZLQmX5
Qpz+N9VOMeqovadqMXT7gI69OvpEbZPpXuDKzCtXvf/r4ENs3Ng88Z+lTpkLl1Uix0rXuGuwQP0R
1lLd+nyXBTobvzMlHSusZkUNjKvoAmKOnX3qd6GG7Nzwxo5KeqJUPThy+rxTwwqgb9EPnka1wLRO
afwVG6028kC9VqroppFJK0H5w8rDIeuRVHO2RhYg9Vcn0Cew0IhnJhp1FAiBTMJWsypwbEVF0gyd
VV7kR7RexATb9ajUsqwno/jZoZHV9OPoZySug0AeTFEiaWuqDtZY6sUh1lZljnPcTyKXS7W0ril1
8mufDeHxZEL8vsNsw89bOjnSDi5snEv6yTU2N1bUhlcD3WDJ3YtUMgnViOCkkrcRETUJ2bD5wawy
s4S6uQXTAp1Kbrp/667qex2S0ihqz6iFmeADeflF5uNoczCGt9p5RNWQnDJRDsTuqGjow6cwVvmX
Zyo7h/HtRn/0RUS5cnwo2N3+6GqwL/iBOP+rBfI+3WApJylA5/z+LJ/m5dUx6PijcNefQh6HdRRh
i76DfljzLuVXstMszbR6+E2b9HS+G54WCCYsPQjglTK52+uo/lRcMg7LYf684af+fy997LMw2Kio
JKxNGwGJzOiAz6YrAwloMtqGf1Z7xVd76sJVpAWu+XX3F8S6wVELalfZA9XEq51lFapLe3qSj+Zi
SBV9c+BKTTp+0gY6ylqnRD/FMBIr4uFCaxLRdgamRN50l+ErKStr+IAn5q+zqgpP5bwFG9rEOLwi
rWUJTp803EcI4IaABsuT8S/x2JortkF/7yQRggF2fg2BF8tDdmzCzdpxBK3qfnVJsx4C5jpL1bli
+hJSXr+Xu56iXolRnLGrnpmrlYqxWOTNrjaipihsMzZIQwZ0dizFZVtx3ivuX6ehKb8XR/2OIHgw
EaUbEMOWxKB1T8sBiU49sMbQS+K0Tkd7OtVN9qCwmwycafotI/kh0VsEZ7IHwsUB/W5iFJpyyRjF
bA6VdMJ+MWqOJxC0oFvcHrn3I2w6MkwtUuGgiihPHkIC/pi27co5/Zp4L1Yebnq8d45NnoXfEy2M
Xfa7BPGDirlplCnGB8ORn7cq+CVGheIYfA/LPD4wHWwjbRltJzaFCobzqTHSxsOME5JHac7xyLCK
NBcljsd1eP+aqWatiLWopY4LZnHkb4w1RZfCYB3Wj0JhXqxzjzVd25VdV0fsm2jK8aDqyoI7CP1o
b/ATPJyTYbCCJh5QuZMSGppb51bBSZsygz1mvL7G19bSFjIXlpAZME07KzRFPUqFdr/7Ca2LB9He
f/Kk9XPtP5i6C94Qv3ArJdxOjyWx3Q83h81E2xwFl+Io8u2ui+n607uHSWK3tQOZ+K8iGc6mUTXr
K3N084ukm/8lvc/wXWmbFpN1sFRI2+qeVBgrYCyJtBQzWdj3N3YT3P+NQLeCdKMHwvqJrAyfsyU4
Z9x80pCuk1TplHEUqjy9DeGhysJ/nCWYHCQGQ8yg2LQrXCDyz2erRC+qgmoD3dqFu3d3TN5/2J/X
3+KktXjp87+sx5b8caKFnNiO5H4tFm8C7nEuaCsMsb1YNfKiQGZiJwMRCJrTCD4wlKe/h+lc6o09
g8Z7v+eFfyGyetAc9ZpTplKcIdU4C60fm2KjU8/NTHNU0Basks+ve9mRpJMuOHbDCJnaD+jna534
9u5/xXGhM2IG9AOcBzoF6yHVlxqa6vRH/AG8i9IKqgvGCM141IQt7uGG+c3U5ZsIn9QG5o/9USWR
yuArrxjokMVRYWlh8qnRJIjb9beSNrmm6WXapN+qqRYOms8KPKGizC4iXlBnW3xWxWMZ7e4EKtft
K4kHwafRszcy0U3tDa2cmR6AoOMPBDtI0f59tlB/VZ97x+Fft1dnUZv95LVX4CtnEnnWoShppZIh
EWIH/xutslOdQuRLx/Qcl5v0dJYjR3Hv71AGILo6mQTsV8J+42EaL7Id4Z1dnvyQZ6/0Ep7PL55R
D48onhFjjq9WugPbbmFbBD49LMKvm4m54frvDz9HmhnhWGB1v+16efjYRBmJ5n8rtwJazLAa5YOR
CZiWPGR7u91y1ruMFXcZF3gKMl9615MiOl3OJ8XCs/MGzNbmDyOJcZTioqV7KRrd4jhoSEr/WijY
oaWPF/ubUCgiwWP4co/rubDswvPtpZ/wrc3/5ydYPJdP6rxmfn42dM3xIPMy1177eRUA9CnCHROF
1rcBjrzDjOMEVqvioawmgvIov5KJaafuHDxKUu7/E538LNxauAqvETr/tjwS4cJK2Z0EcqfEUUmY
nNNjm0dCFlq4/BL4eCXytprMS0Uv9PSBmb6Fyu7ISyUb9VFfww+vZrlz88DXuK1bbdq/F881HYkV
Q4CKb8noz17a/IZ0X/zRA6Bo5eqXD83B3H9MUEfT4dqL3/ycLlpGK/hwaBPWtRW/WXKp8peVk1MV
3cMPwWlvLZ/PfWbcGSIT9nNsfUAL4nG2rTH0ur1PvWJmb25LhCr+HfKsfXgDJDMNqmjVgHUleFP3
DigK4SVFxZinxtgrR9PDjB7Q63JRIQNXbSkxRL9u4AD8e3FG4lPRT1mi8d6j2oewISEGoD+ZgP6E
15eSlLdYXiUwFbd3ZKL3kHEd3HFkXjj0YJ1bXCBF27cwEa30tEkij1wk9+Mqtiv3ZOuwu6nBWEAg
EsPYtlJDZ9zXkCehYA/QSDVeaAXW5jOCrhGRdVYg8Oj9h2xmu6ftcy6NIkcdiKfijC6wSUD4u1Ey
0mQOVP+shLYVkurvk4eK8ksyjVtrCNwTxUKpgC+ZeqJ0zvz8z8iyrxlKW8EaBN16lpkYANZZxBrh
v9fFn6H2teumzkVFp3VYRmq+OtGt7eqYQWxib/ld/mwWIfHLThNoPTVQt8zyOP+FDozrDgk4AYkP
NfQGlusntaCMDhdOL4b+KcESQ9ix9luxpGIrbIWGat9otpzRFm7ENeD3fRQWyP5eZsBECKyzR/RK
90mpjOyjx7Bb3v+9iaISclrJtckEIzQ5M+S2D/Delwb+2bx1g7HTRUg7uy9G6L8U/MvyLXbYQ6cb
NHLBMIkJcZMz3J7uDA9Kz5Jd5nis2BvQFl4qotZmVUGUfORKAhcUlzrTmDLiJfJMQFR4efozOoHh
1XIlFiJMxoEdfAFxZX/ufiqctd2GKT5n38qHAFw/Mv18DMPydHczpoYFrmO/RjDJk1t0OmTEG1yN
FHtNqfAAyZ0JqXzKCP+uwMf3k7VgJlm1VaWSn+80wKeeDr2bDv+EGqxo7cX2uxMo1KawLOCFpArP
/ETGWrlSZWnSeiAziaxU3QKyM7CCByTx58v6OBtck02zqNejgA9w7jRR1c1vRZsrCY6UJOBaKLPS
FFLX0Aq3nCGy+l6KPZRJBiE8fDj9oCma06yrwtywpHku/PukWJU8lcwbVpO9NxyunHAC+6gEaFBI
OqlmLPVxjGQBn4L7PyqEI4jG8mCFGQF2PO7Ax8TNPmWOzTllaH3/f59+5y6N8sPUF/5kEVV8dUS5
8KQmpIO6TbyngIzVv/w5sT7lF+ZHL9JsxajA2K+Nbwki6ReVcM8BO8+Z9gLazP3xU8Kg2hjEAl+V
Mlc0Cx76VSlTCZ07No8701EStgrzTg9qNjfCU5fpZCiiNyqv95hIbrecGXvNjJ+5mHanVGklfk1R
EG+hJMj8p9WUcGVEYhU155UMdeQ+zKrk97b50qASuPXDoQJ9Zypmkn7r1skJS5kK0JB9ZTMn4jec
QWp9CSKFhdH2Pv6ZQipRXXXF2S1XcxnUfLV9Ut0iEzYO5GNzDi1mluKMMFcXIWpwI56stqaGhOaf
d6cNY8kNRiWGcY/K9hFUSrVlVKlL1kuEO5OmAVhUKxgqBPhMWoR76F4Lkd7jjAdWYB4Uw1X8JCAn
ujdQPTOOa7syJD4zzG4bkO/dbm52FqO3sHstd8kt7DyerPSgR1k3ESWR2q5IIApnwzJOHVszAV00
2JtPkKJS3TyeJrGi1gcmcn81ZDMXJDcZKyxRfUBvVylwRGg1WdzV/MjjpoXZX312BEQ8T9R5IqRv
sZWIU/nBi4cH+mWGoZrhU4K4Cei891YvSHFFxs/4tZjk+S1b5PPfyMhJOwupB692l/c2enRbSST5
03PmEaTBQYfrm6MDCpF3Cj/Y9l+SIJuCKn+JDWvG88fmUeUlOUeyznOry2APNyoS4psdAAaria7X
gO62gxQIJTvPqhQsjrdllkdKf9ni02e89tf2HrTDX3akP+SuAaYdJpvLc670vU99eEY4tR/C3mbQ
oDerLqidEwqFUT6uFfcsXyFVjnvQ/f9uvL1Ozf2T0d5egs1C+skqnovoznPI6Fci+PGh0XZRO1fK
d5Xe/oahtjlLcA/5hyVIAGHltwxqJOTcIJuhQekfpT3ignylAkTH95dOPC5dBReaIDKDorpuHmHk
VnYglO3SIbgnoyKkLejRo4OZziTeA9ApT1eRr7Hfuni06YH1w/bK+d8sQn46sgEdXHYVRrBY+XFl
UXiyIR3Z/SUAAJe1afLGUEee+td6MTkpIb/1X2qG1uT4fV+LkRtKmCFy4poS1T+1pAa5XDxFO4bL
W5zBxEkzUyc6J7Za6dZnn8wp49wlcuemX5tirCnJw9wsHiIyjQJRSRLt03fOeJMg8aN3T6W8/C2B
lAqzumnSuWS14V4S/ZGnuvEKniPeEyySB7HoyaIPiFMElkHZGUCoap748yefchQtTK5KdVSBkVPj
UvWMEVT6yPGPPJrZrxSBEww2+Dy+w9iD2qvolQL1Ju8LEnt9miQbYEjKXktcHnSRBmeqRc3YJzfy
yUCJSpb0bb1b0FlroHJq6bqnq9/j9lUQ6HecKfO8zMHqCzEaw0De5oW4Ubt3ceajPL4ttqA5K/jU
2FCJx1sunnD4cv9BvS0cVviHzgoC62wWcCH9fWXEqxJLFFSVKRwe5/I+MRzxLWHUATQ3gZYrVwJh
EVZk6ZpLO+t3bxpSsw+wV9kiuZkkNHBO+UwtbDJLdqme+9auzh8P2xDJ6xd8MdlcPhtVnv8xcMiE
wi4QUMahu7RH3qqcOEH0cVz6XqaH+iO6Iaf30ZpbrWiaoDfwr62KWFJRYf297eLe6kCnf9MOS2R3
jTFtx7jLzAchvo0g0fXThG25aHpiNfI6EFZO/39uPAtAUY5vOiAEQg8W6x/98SI7YYp32YZusPKx
0jqSVi+ciq0yRadLGULscj7Z3bpr48+Wc8Mv0HHPVe/A2XQE8Ux+h3kzl5e5zo8+5y1ylk5UQX3D
G8Y6vK2jjtuTrGwreAkqDgsqi94ReGYDvb4I1oU2bw1vqxGmEAkqFtgnTHg68K5AKbooZw+SlsDA
m565eSBEafl4XNwR5Lv30E8x0Gwak0nTkClyvAscYaonPw4qSfvcPv6002hnHWwrLtpk9eKwKNa9
oWYqwLS4tG6Mb/DfINXi+ZZ1HdpdvpsNiY3JV8ud6jjpWAPjHkezlbhaBiBBsj7P0ygeJem39fsn
I/JKiv3GtnULVciJMcYh1kk0YXJKnWj7JdwSI3td7ElQ00fPZhR+FYpV0SZbLkNXFkGw/9xjen3G
TVwVqxyDSobAy2uOWl/XWIenwCZRYl6nZo/VjT5ahQhr/UagumP1SHe5PUfVQplIq3LgTwKbIWdv
m5+qiX0oOB8vehQgOamqyToJrnfBbw9eV6ne6gBsYrsJ9MT/ckthnwGqzIF9CChwABFuB9XiZkRb
TmVTqn3oS9ZP597qU6a159ItWXa97eOhohwMh270L51dPwMzR8NVtcsDJ2nDj0jKUnvLrlteo5wq
83ryLDqcv8RMfnh+95DMau+x7BWMyDpU6OjxcSJyYK+/oZftCrukY5J2tTt+sKDFoD22M2IuI1Ac
oUCiIfrpFHYzF24erz79XwpDp8g9+9v9ianIVb3MSJ1qNM74nauDYnmOl6lZIJyV9KJZDS1PJV5/
JEwGsOmcaRVkVhV+b63ag6GOVznMdxyYVWHcDd35dUutumyrbKMvBK04NcOq/EvLUPGgD2X8yJKc
nBDlTHyQfv1QwZutDMK2BcZQwN+UQJKmTes4fZjj7yjHDSYF74v3ZdWUbGK6nHaOr+LGNT38/PBb
ZK1UHzsz8rMqWVL6vAhJI8lS/YeDhezZHvS0nxIjXGtK+b1XPgN7Vu77jpj9eTa+jn8LWiXSjlAX
ETTnYvSu12xqBDjBLFD7+ta3a1rxtXvOAsrfqu588CLGEvxeT+VK0QIB0ZtHhdZDwl2IPwBXrZyr
R3USUbBWksyil7NAwrfsjen7wCo5qR81UiWkIZnEwXOE4OLfSLXoINoAJw7q+n9dEnq0S7Aol0NG
w3XBMNT6C3aRwr68gQrirj5h1qKEzY+3xfbXhI5QrZCHSE/wm2a0IHYhgrpvhgiGDHTj6O1EkRjv
MuvwOw7MvW6N/vt5o/8hyEUVEKfKXKDDKEJNPcHBZhCTWlLNDRQ6ZYGIhYcrtVTN33N+YMChUscs
DJIRMf8EaJc6U+qLg4wt/JUVZnFbHv2qwiMek2CxYCD16v9autMnw0tbAucOwmo88flRikW7KtIZ
VotnhHZphgBZ+MG4VKNSB8PIcOA50VAwHA+VPEbsE+jvHpuES54GmXV5DfjODdYraNWVs0j/ya7E
4mjpBIFLMRMoCoW6SFYSNEOyKqXRYLDTRC5CVAxxI8tdAeQYn9KsnJnX4ecs1WKXS9M0KYJB1U1U
MOmi7/l8NkgPM4yRRUHWFyQzRPhy0gcPkuykI4vJogT49Rz4AYYj4COe6Xuq69rWItyO+fQG8abX
DXuCCo3icq0hIpjHSbBqjJmShetQROgeodiptrY6YK2oD4staGZh8eqqRrJjVbptPHLxJMOlulMA
DHvN3dCyje/zvvrB/tc+Lr9/n5hghk+AiN/d5DHuS/me9M+jtR9rwGMQI2aePfm1Ko1ml+EoZaIv
PYDY93DsmacKzYkqwyiVYKBWwcot6oPvsKmiKHBHIZL7gotJonwOWueyUUnu45Xg9dlKBSJDrQK2
7tLkmnm56z1cylEn+nrKX5RtWtmKOp+uNb8/p7sfpfgoZueBDJWCBZ1W1aal4bQtiHfmuvTbraTa
OPao2cHthCQ88JnUlIazws4nYkV0RnG/ICsznWm9S7YBmKv2sktOlH/Q6p9p3tXWy7LC5ztkdW7k
kE4VAABLleou5JYvJyDA01K2mobzKP/HadsDTZPIeC0hmjjf7xsrlfkzihx2V4bJ+8PRoemFn8HC
8MlGROo3wEBBDNJ4pXglYke51H1HteQ8YiI8/z4e4QYqGJyMEL4LrUeCQycvsBaKjNKSu46hsvBT
2wLhAHlQz4PAmzOL3y/V5r1gEA1XV7iyY4YbKQqbBxC158TpDroclSuuLVYECl4iVZnBYt9VYkOM
WaVmWnMaTbS89lIX02nBTqxvAZc1yThaosAbAWdsDgol26Ad6vfiE2T72qykWWe2CW6H2oiBjzKG
6wenxA68EpNwUrY2rwt0bnTGCJQphLJfiTth7/+sAont1wQKKeQfNjeH3hsGdhfE3gzhdIJzbA+z
VhXGx68ERoVnu9uSeOXH5NzT2xed+ScxUR2tJYYZAv2cTRSx6VRXsWZ+Kofa3t6w4sTZd5bBez8v
tnN065yiIfPZgrfVxw4D8y//Br0VaWyFATg/jeLkfr1KfUY+Qv1MdoUcPo2Z5weH1pCbSMoh1dVe
GLiPTFus70jfQSRH2tIrNA/JwtByDlIuRb8Yz8TmzHonhiTZ8ltt9doMOphFxMpPJmjYjMtOxURW
ZEBhOzEUHecQGJouhWYNWZD7CfdOVdQVk+sWqnWt7x6TAWVDVjZPjDCXHkcG8X15Mzrvdasa06w+
GQV/y8hdaIyy9oGdumgdRJSo/WqPKFL60iaPp1of0PR8GDb2aOWhtLAFZLdmpplEo310q0hLUYqh
HEBxAUC541dPulRAqj0/ibiGfmkVNIvNoIRjeiqynBk+NGLYwCOeK32809DC/bfh4nG85ZvyhhXt
vqFaWo7aXBwO7Kx23WsifDIWHyJaHNTV8cWgjdR2XZlSKvCrgc9uEYr3+zp9s8K6VgHi1LZOtp1a
GEUYS3xTtLtYp+DAKht10VuRcKbmW0dn3i3Wdrmu1EMPpk3+IhbllixH+uMk9nSXPKy2UvaCt+Ee
2799FZIHeL/iO57RLJdpn6UAjTvTkGCIIuYDrjqEtR76RUSFyq7CfpiVl12Zm419cx/Fa3NNlWte
eeDlh+nMOkggaVlBKgAvri6TcklZh0na1DskYmO1p4rJJJj8cszb+QszTJoM6IC1Irr/QJdz3wjW
WD/eQVHpsYHYtqHiFPokw4fW3c6UJb/CqEbn/4V5kwmWx8aktuFnQI9Uyj9Nim9jF7JbIbR6S/nh
CCUk9bL9zSPs2Z17rLPj2BcG3X1u/jADRotJ2q7pHFvic8MITGxJg9pqqmGOnWBnvUgXX57ILFfX
SaoXiFS/L8bs3ZKuDZYzaDlMIcvnt+lzc8m6nqDuqL8wig2U1sYEF3BJNsiRHffKO2LYImfkOucG
TFF7+esZiAaAx8XV8epoldxTkdhO8PUOjpIEgDth3H1KXCTG/SIuE4eE+cpjuUfl412JASYygBqg
aAE+v4qYB6lSGPLn3j+Wtdw5pNRVtgxalDitHCJlxzYQgEWK5dskNBeSujrw2XTLPdztHCGRUi1A
EiBT+qE+5A1jNOIYkysDHDlrbC3B8TYGvfKrY/njyenUXhiqF4KROaMmtDvO7cIjo44cf9JAJ1Xs
Pgx7xSlF5soO9mvXPk91U0jmXSO1LQroGwjg3iPVOtvWIgRsgbdLSKmZqOZhPGnBLfL77hfilmKs
pQtaPmlgeIALAoL9uDvTJliEpJDHT9avx7sfsm8wcWdEcAb3RhE1UbJR5JT6W/3a08OU9wgdyNA3
S62LEl6B5/YQhuZWdUJMcZ1o4aCJvrDE9BQnTKhF6sTdazMXmexseeZa8O3aR7t0JaGBFxzcocCg
sWZC/47E3Iyhj5p4EZOJDzJIfR5uZ1OezA3z1QT8/pndnqHh/o4oFD02QoNx3dOC/oWST5N/aVke
S3v8IxUcoD05lUe5aoh+ZJmsgGVKR+y2JiM8AUJgtRiWPmH/Bqq6wj7AKA3tN9OQeJuV0/berH03
SnLXeWfkCdX09y3sMe5/40UFCwnE4cpFE/ZJWZCtmDI0qX+AWuVSq3JrDiEg34jcVKf1MIYuqLXU
UIpvw2iiKOoKP9Ak13m1DSK1CQuTx94ccof+7Ve8Uim9pYefSLzd20NOWWsCNKOgsNdUlmikB3GW
boCGfxtOrDdwZVvA2D9/Y/SnSMNvR/ht7jR/UMRM+xB8NJrPOby6NuVsJNHWnH1xNXojMk4LYIuv
GXesRYwqPPDuENvDQsayG89Z75gMAS8r6EeXhKZTuWvh86XxJ4KIbU4FGqlC8T9gTSQaOoYA8Bt7
ML4Q0uC53lqXxMzwjJknE+gfBjL76xPziPmTwVxz7otWqdfE9O/FvCtESSeVBlBIZFzG6/326go/
HihXH4NReA7Ow1P8IGm7dH6zSimT/HcZGli/yUmKi6aMWnYI5jTYqTy7emhQIEf6Xv/4t2Txwkxv
6W6MpiXiZcHY5C3ee7abgKkkNaNrshsHKAExxLKhHsulisTYkLHRjPtN/byM4wlI+R/BALx+L12v
08tY15/Wj425jtKrmAgTSUvm0TXkpe+tXQkJ2ZRO3+kHp2MaBy0ywyO2Yhp0JFf0VABZ03Sb478L
GBwSvtb/XC6mrXyhBsXBljxdICQdIwtMY18t4ruyllacwmlvSZMFtODbSsTuCSe5dp/U+gq3tZot
mZ/aiAyOkoRw/gZPb6GcVqilVN9xnUEC9k+j3B8EZzCY2G9+pI4Vxy7nKSOnDY3UTDov3MI1sZMf
lmte/+0gC8bNVkomyAEAdbu5gWl4TfjEkHW2is3V7Nq/h0ryqBjCHbjvcSsXLqxfKSUu+I2rHd4W
z83TZfTRwcwKMrpzRhwN3MlO0pXgZdIfNsDlACp+jEQEobZOWOcK1Pevuusqch27dBLOmfevyrBw
vMVOnkxTXatlp41LOtSkF2j6TdlYW89EjdJtEdutYbzQ7ZOjVrPpNK2puIgA5PjZ0H35KtYmfe3r
xAo/lhB08HW/Jh2ayiMjXpm3IfyCjK+wirkZ6LgOJhbddWYVrJZoxPLzztJcU7EEvhzCXu1pR6vR
yP6ma9jCOxdnP3IK/n2y0plDIZ8WQM5qsfcB66kZUwP6i8Vmx6m27wTQBtmRvuldmDtngatlZUe5
x2usk8T2BPk4wquP+q3zYT5m6BajIZjYiWTe8lW8jjO2U/IV2s32sqEZfdVujBz7RAKrvH1erXXS
WiD5O5Ky2FQQ+kWQRcYYtydzbbsotw0sgyvehx1SGTp9067GXHUToXSakmqTSvfRlU+3G9fDf5zA
0GyMI0VbW03C5UIZLeq11pHhIrFDCtEECR7v+IaWngmoIjpvEttyi/mVEzF8V05+lRzjYM7lD7M0
zGB+802zHJEeZz5QnR+l5vQo+oOCgJoKIsbQ9E1giDo0Q7cFM/V0BjMn04VDjGytVNpg/SuNl21V
EoEH9D0LeUFXBKxqAiFFmWOLVWc6Nur6aMnA6e9Mgy9BdjE2xGHsHWZ9B0wM1iGmHm40HXg8H4JC
EACmLpQn9Ir8R5ZTQIXuwJevArhIoi1B1NYkt8AbUlQmEjziP0nQTy/P/Au1Fm04+ZStwjjSW+Bw
/kiXRyDSc8Lh/nKtnA5bzIyp4Qmg5DQevRQ5EAyUaMuT2PWODq35A7MxAvqhCfIWv0jY3pH38vox
AMX72UHnA3t9w7rPVr5PGaPBJYdE0Qi1MQBM7mfZDKvZqdVBmDshCq+hrCn28B/bxtBe4orJAkc7
ncfCnIqMpyiATyjwnd2jT8S4EdaaMu0NMJsla038xqsNr/DA4FRwwjDSwm3+pmDoH8Hv2KESbDae
dBRGaxMbgNM39/uVmg6jamei9kcJT+YmUo3oiGvybywD4CFjmSK3uDbQmIhVFmQ2uhD+ubUOhkH9
SAeD+M0SoiXuPHc3/iaWOfkQISycgLxIlAs8fH3fEGDr7VDSn8EHBCB4A2QHl1MnRHWoIB8fpArM
yYv6dTifNgfJi6STlMwJPp64j+RF5CMWkUasQz+Z03f2VwT9Rayu4hJhXe2XgOjxQ8SECiBQnRcp
sYDqTeOfKC+x2e78h6HJDWzMNONrjj0z/BV3AZXYkEj4bDM7VQPPwXP/XDhdcg8zaBxLjOJfYOak
tWvujIyyA3oey9p1xYMx3tZohxGAjPLtPQqEZEDxxwDESDdX9QKoLEB4gw02mkD4m5Tu9ncYCt5/
mCshTOuPIBL38oks2o0yxuUpwgsnjX9mtF8bcKPf+xXTu531D4tNS4oAQaBfR6MxOoN5ViugnJf6
CElWuwXbSVpWhVoKV6ZPJWmQhfRX3dbi02qeCNff/IDGzzkhxYcr4YhuF8TPUIS1zrs3wlQrFPws
GkNT8IyIfX6SAss/b9eYIAur7LWw5VxD9DhTWEWWS9vxRZcOhfak8K5t/TRpk1GQ7TcRaqlGmF1m
QGXvFebsEzo06VFqTIwFYKJUNu6AwTfZc6Kvf+E3LoIsc599W/zQY067bfgCMu2u2S8G0Ull51MG
21ZMOMlS2uxLkwcblUPvlifbYoB+r1coyS0LPuaHQylFcVP1WDabLT10ulZFQRg6EmpAp6gUHaNd
MalXnJGESd6zIIirs5a/8eWm8CLLAiXgyjtXZEy0ZcTZ3pz2//xGOElqmj+X1rRca6veStGU/Ho1
XUseUA1Gum1zlXWK/JvgF2hFnZ6lU+iLIzyEhyn8BcIFepiFG27Sht4Y7IAfOV720S1qy4Q8akwk
UlcjfNIqyn+qA05ve/brsruO7tbIa2JNa6etMbU+dOiLMYBN35s8IW7tVQlDnw0XmSFZztHyftdY
3tCppMEOprMIZMI4HreSjxLBjhtrwD2IrKawh868bCOxalHhcYEBZkKlKHwtd7lxxehCU70AATft
eTDU5ofIJx7EoS591R+6e68zbwtwuxbATHJGscmizLs4Qq8Z+RH8cyujkdhh/P2KYy+tu8JXeypl
EPSvc8YdgYqFntUlPtyFlOwVjTH6QQTX+bM8IspNn/RED4l6anyzGXu+Fe4Ykv2wn9Pkhif4yLHv
T1PwCiyqAZ8g9RNnIp+DDt5SKcbMIMMWeeC5lSJkRc9TxwwyzHq0ZLWobWvneQGfL76bAg1RUlRE
n6/hKPYneth7poulrcQrs8XR7gSGOWUK4ScGzL2XNqz8eHpfo+lbPIBlxaWDKnHNGl5MTZNXe8wC
ryvtfuLoVI5ceXQpexCtdwfDaU3kiwFwH/abn63GicUvtJzTPFR8XHbvXNr+TZ1+86g/veY20szM
qAU/l93v2dgCET0dXpDJZZqBrVmE2b+VJpJ39KGxS6RPb4qB4jWK8fHLzaEuzqwzxhrx4N89aUiE
Utq6sra1JEBZbiOMkUb0rjaHgKdimnd7HZKoyoiNO3UtfdaRlYREyjwe899Y1ukMQ8iqJMMLi0sH
8RPQ+Q2oYMy7EkW6hpHEbMMUFpFE8xgeJkc0qiz1kCijV3KqOzmj0cFi5F5NicytSjLyCX25DzdL
6IITIX46RVwLsX5nHfIdiL4E847zRuC9oVvDoLhAd+CPLEdiv2bd3OoMzbOYjqysy5V2YnQmChkC
7r/QjKZ6fMlAa7WpOHXHH+460oReb43ttPchD9lKkKuRgzS0osAJqnNbnDud0yxd8h2c8OOZDpEf
VUvNu4qXrFrG3x1ohPJh3gqJerMe+tBRda1kec5WNrRHDE+fvrzcSHy55KYR7d1MW9BuV2vZnJfc
Ova4VodSLGuIm5Tat2LOuvxUvGEMmvm63J8CSfgA/Nh9rnFSHvxoeYpf04gZrQ4HvdvusEzcHvnF
gYwvxYaAkk2g5MDlR0g5ktNNT/4gbh2GVrFYLTEeDMVUQcYrGqVOgLmu1ROhvTPhQPHgM7pT8wp1
YubudlL/STtb3SioM+tBbPUIDbDxw8P26cs0tBsVGF7T7rMIF1ePAFtLjfyJZeek51gFC1Ju3e9K
t8o62jX9VCz7B1p2nntOuK0rd0gUN9gzoGvX7NlziCZ410qptaUfLGec+f4HV1eq5wW31ZBTOeHk
clKrtY58oSfTcjaL4zCKQvl9feVrG0ZbFZrGIC6/bsuxuK7q7CG78MCeDXkIDPKnbXxknZ/sntCR
PWSGtgXrTVqsdK7gQmc/mfIpPaA3ZgwgBmuRPHmQp1SeGam9lLFBL6UXHpRGpbYacSPzSMhvtJ77
ZeWCnGJEi5hbAu5eA2HtkFLGHhGKBaq0dezF6+Etik0VLdnsGGwPJS2bjr9wnfwrv3owdJQE5lpo
KX6zLnf57L7tciS8O8lMTuGlHRAKmRUy+mphoJDfUJRCNTgciZ8w7SOeh6k4YAtsdBmPuiHX4S47
JhTfzQCh0pNGGT/MaTMBfvIyQfUaagl9nxvhFb6MNAm2mbCCFB8t2ukmRvobdqbvNC3DmmkHplBt
bQpj68f4Vnlr7RXQC/p0g98auaTwFpMABA01qwObaWew2xm/JTLe0mj+/Qs990gxTSFFuBGf945L
J5rNBtV6OQa76bfaPs+3eHjTaP55S7z0/L3rqI/ITjmgYvFsjtr06JhQ34DqhV0x4FQ+LcQ5gB7j
+OdpdMpmNpb7Pzd90uQjyBRNFzuYPrLkpWeSyBQr8Uvli//Px9oAuKOmHOIIUghLBn75MpOeXVYt
xtnzcyB83pn1Qc7uNrX6yCIE3JX7lggzTdvtOzdB4ZGNYx3h4yKSHQ7bVvhK16uU0DnBZGCRMZP/
l78IeZpe4JVpBfzUVsePGwokO3sWLIw35aXa8KyBWIwILI4xfUuI1AJr1x5ki2KfddgFpC1VmSkO
W95E5ahObIkpUiW9DFbhySViKpbnmRwccqxl2nM1kkViimcSU/LJ2zVQB+1nZAtHODMAWPdqhljV
HLNB8Rv4WT1mEZTWnTLYybyfBDqxVomYCmrwgBrWQ3JRV3WD2X/TN2WzXc31U2yxWAGFDZxy1R4P
AUm1pKiVGt5dp1dhlrpI9au6DDAnT8iY55DMTH4JOooqR9p2hF5mdTkJxKyS1yLXzTC9/C7HVgsF
2M08ZyCGPFX/AfxOktcH2GJ1et8z2a5ravG3inESIS2llwQZ28VfWAV2DY2XEfwvWrgyZQArQIWQ
AmDGfkjyB3zHJyw47CkfdcNUFUzE6LZI/nlMDaqyOe0QWEl/eGSVK4/GpqgFFbxzpqfYRCwZhjF1
z1yPHloTuO9uGnduRos2l2x/zDwm3fWd2EPT2thRkoykIIxag+c5gxYcorW+MSvosgQqwRn6VMIk
sBqkXeQk2QAruE4Qs+hvEa/UJjc2mxpBAtSngG4ptSYVcWl17VygcmobX3i36HyBQ3bn2/s7cxzQ
AB4Vk4FALjdJG3AqxJyZH4yj2sJOcWpy4Gvt2Ydra13hb+lm5/Pdm7ep78w/2VAqpzwVhBpX1/+f
iFPQWhDcr2MC1aSFCCs5Z8iQ/my3TS62kYDNDe1lcDcNIw1TWXDIV4Uywjd2QV6cCPFYHQxUPGdj
ha/C4+ikzbFuHsTqRqXIR7AliPg3DBCT4HQuUZxyMCTpiRV4lQn+tKhc1Z6PjA7P0TDeytZDBL6T
+zyJxLuGheUfDrgfHgb10HMcsBb5aiyyeD6yQTBvRLVw+GIaKYAXFdbpS/1CUE1dECrGfqEz5fnw
AuieEz1kk5hlxakgRlqTtPLEvrbNv9hk4oz/u/FqCKadECOU4IdjGciij9G0RHif+B7L5jL7vSpy
oLTJsbugjk1lpSL+MlK9QXJipKAlaJ+LOgIdSTIkyXB349yjAaOxpp9EFc3wdWNEd2UgBlL/uWIT
rTJtNqpPX3oog7anHBepg87uLd9TJAQTPkHqRrcW2klRM4V84G95cbGDkVFZyeBPVPcHxcMVHYMp
IM++3dyLkQGShZ7xC3OvoM/VEB2zSoIbHp/fbc+4fDp1fJAVuJxh5jnwodlcSLmGY3MLUkHUon+N
b7VKfMJPPORA4uhHnLdBqDvDp0pkJA+Ny5rzGatBzLTcEtg8V8VZKGR5CuPiS6+f1+Ke5NNeIuD5
rrck7HlFgffZfWIDz2d6kvyD/FPrFqcqM/6Cj0iWiIdc2ZR/hT48mHyXmERWG7T+dMwVdEJQQ6Yo
WhiB3P/JbWLvovO959GzrC7PgiNYnjcadylZjJT3e9rcmgj+onLyTWod+CqBNCvee8f+0dY+tsZT
bNiSwKbDKc/9hu8Bx9cWyvh7Trt0WIDi3JxKqtJHEIcjgRgksbAfsaVuUfj4fdZ/sHvg7LbXRsv6
BWZg9jz3HYWFqy06uiskvy7Zz7gvp0TVJHcyuZokLx5H9UaCDTvZgWmpByetijY4eTAEoGSgRDow
0UQsejOL1R8MfFRWN1FWWEIFQHuOVcBF5UZoJZ9u+kjmV+XFEoj5b7CmBTVmadKKrFsI4sNbofpg
ionCD1771uWKkjXcTCeXti2YJIo2NQncG08ePD+0Kcdhnq7z2Q8zlSbKZwzTJM/ocgdX1hSekB0z
LujHaOPkhXjujC5iNUJvLxL6p56NpMu9Z/yujX9ov+En9DxkCgT9QPqY4eIHzFn/TZkMdhkFRXrd
BiABoxrzpdsXFucKM9pjXWFOWYPNEZg58ErdDweQtJMyGCRkgoqAsIPBfl1/ZFandUByClSctcn8
ha7lvRfX6voisMYSPjH9+DpvZijT1/RPK19hDNa2X5B/9frH78evWqAx2a14RXiHAzeR+16nkQnC
RWf24wzCQWvjDoPGkFQRodtE5/2RLn/B1SOhfP2tk49LvLlnOBPQhc4pRlTVNh+QNSXLhiokCWhS
Mtxmf6LnXA5Gme45GMajXKVKcbv9aYL/TDKW5jhMX0b7of4eGKot7Zfb07c9wLfRL5oEQWJ1AMqx
CzyUZg/iQlFfaQSQ/BT9NunRYDL2xIbzECv1vtv2Jezsa3zbxZtVZTwV3n180EdDV/rGg4lP+cDg
Tx9smT8gPhYqmGtrGA76OBYEGIJieaUfCKHjrDCYU6zAjisixoqM/KSNtUxT3mGKc364Z0eqa/hJ
LDKDTVoDmrwwa+lwbiI4kBQOgfBVG0iHkrvt/2A77LlqqkOPDlhxR14oCBlXkiHs6T0mqsWqmJ5h
bf2mn08hTR8FFmLsqUykNScPeCn3Ti5cq9jeUfQVBH4qpPumBnuOuxZxGX8IMoPSrnaqDNKmNBll
Su+yUU1J+jxB9YiBeH4UBu6kxS2SmwWWW8ZvDPCLQwEJrfgnbPafFd/nMg1WYUA8Y8/e5Piy1pku
ccbeeRl/WPeXDj6GkIA2F1Vg3v98Qu5QN1Rxcm1C957o5SJJGhSBnXbH0ZvDkXDgpDyLjVf87wJX
hFPaWEKASrwYAw9GLfuhI4vlmhT74Gsbg0k3Uij5tmdR2lfNKwaDuiva5hbG4UxK+Tz/INiAYw/W
r4XI2RvcsRIAZVVLgRMVwhk2Lm3unvMfMP5sUhUac1COOA6gAMAPHzp4GYQ4ttgNDm46nhRPQvWy
5Fu+z2vlTX8rOPo1X3mCUd8aSZR1WPpie/YZzb5+yd+qyra2oZDpHdPtkJ/cR8ZmpHLBIW8S8Hlf
eIg35zfpth5URtlzMlNVj9oLEU2foYg/uY9CoocmR9iRqHB0LSKOPEXzSlLJ8l2GY4DfaP9jnKSy
4OgBG36qw1CpDotGvM5AvIXSby5kZncouZRCZThsgoH/lmcyQlCvQpdPclH9Lf8RCpL11W8mVM4S
2I2oFDd9SsupWiSCKcrUOKQpFdRy6HXM8sRKiKkw4BDRv4p/Q+Y/dteKv3gJ609WWgwIxvVk66+W
bvnb/kBV4T0W4LMP5uqJfI4qyJ5mjcbIYxeue6itC9kL1ZyKp/uA0DmmjDf61P7NDSzYO51ERE2G
3Ii8FjIj9AqO1GK9cTO24t/6GLZPiu2hBkiqExVkrbiWD0OMrUhb9ZsSDEb7vUMtzKxrdjXhIsYi
8r+TsH9RAALxSPCAYVL5fY63qPbleFB2aQn+or5gkSsEgWJeDGa4Z/6gL5kiaEj+9ypy9PrgyXwA
MN/48GEgPGr1kCO75U99fZgVe3gFsV/dbpe8Bq4emJlKZgWCj1110iuqNdyGl9KM+JR6iCUeb6Df
EPUd9z8pfbM57ckRs5BB/OCLhxSxkCGX18Yb5qnCpdkGRymTShhwqm0N15loJkbiCpKnJQsSYPh6
GqyCIduuCM1EgvD3aJ5wPvUzAyTgGIMpYIjcK+wyKvzFhGh9ZGgqMC1adetHaEIyyf/kleqaVhZS
2V5fQbAgWBFCHSOyn8kwv+DXBCzh9puUe3ui9j3XS3dG5DnUzPY8zkq7EDtdvNurFkq10VLEBFmH
vBSKHRABjexKRxW2lggHwpmj4mZqIc7PdrNuVg9sOZue6wvo9CXOw5j0D1Yu8Rk4m9d9q/byNJmT
XVOqbefBtndsoZuHRqDBnqncSK7VUJdR9IFOh4hvJSOYUDYGCPiMxVAx3R/8KUigToQa7ryuc0m3
vo1CSLlEXLaCMPIWUhk3eWwwYgP1OMeSnOfuXGFtlDO9aImG27M+8V0vqfoLfdgAJWWJVI9+QFK2
T+6gU9Emwm2DLqI7qyjPZMUfxOQz8tCEDTYs65JAx3IdcdANUkz/ESEKPMuw4ThjADm/27eCnQBd
tk/EW/WQmb7P8dcOe7V4lZrNTiNxAE6vkFbGZGtX4g+CXNNtDNjovtLjuMEFS/D+zFiuQPFy4on4
X7iSmpyG2ze9yvJ9hIsThg52oUenaHMac4QwC2bsp/54tivx03LkAjoDlLa8OwEMUoX3WyhjA8RQ
9f2aUbdtrmWZfcY+xdyD3v3kAZEUvcbIir/QvVgxH0Vz+IyHfSmeM0gmdK+13P9WC4KGR+KYXQpC
KKFVCmEDXNnDobodMuvxkTWajjLIXGTFnXlc/EvKlyDXZPIbkQYwJ8M45+O3itLjvKWHkdVb6toc
XOZBOnnYp2Ge78mHDUi13qSu8aIIxIvC491Ru89tfnL/OZBfRtltK//KGiAf3rAl6hF0NhOZdA9a
epwg9BQGP+Vt/m35ABjYFpszKsAAyjm5TMgtf6EAMPHYEQnsjaRbpLZzJ38L7woPUBhjQVQh7FrB
FiDwj7F1EjNsB2lkg6d988uU6LPwB1O1lW09ym5FNhzW7ScFFywxRGHd43Mw6XmTdRjpwFwuWcCr
/lnjMSR1YDhUy8MHablTKSnsHcmt8AOfnkZ4ogNnlN0fAKQHy8qApncmobD7bVYEaPO1+vXz+jIR
GPyNmTHIjtOaLvXLvoXpLbefnkefDVZOUG63hv3k3zc1/4VC5g4ZyO9GJMdXbcnCGwtcZdRv8+mZ
6YJ4Mviw7O/h75LDMDozk4P2JpKYpn0+EBv3CVaHlGQ1Uhai8hceqETfl5FvygtjthCaTyXjsepO
tWAoWP/di9Q0tazJTtohUAiqr0vtQmrPu9JuZGWdjp+Exo3Iz7U5NCJAAKs2WsiZUHS+st+0vYhq
XGmwTUMWTBtcrg1lF38lZ55CXTjsshjl5/UOYlkkdxio0d3ruU75QNYSa6qb1sadYGzeYLfS65o4
hJMeCYr2NUpTKwacTi0zD1eKWeRU8nXN/auFyOnKJfjJWbjfqjPagD0PdxesXPE5teYElqVvGZo8
wuLlDnJaUSmEpe8r7HsUrtkBEtpN4Q+oLplrURJelR7g8hTMgmkLIQzRTYInNMpW4SFqGSY9jSnj
/fxoORXRN+jorHvYXNIBK9x29w1fcM0XaduPF/Wiiqm4AXNcRV514a2zPs/fUCoL1Xw/DbtaDSFk
yFh4JX2X/z/RcE98tuUi/3uJ7OQicX2vYF6naRTKB8Jw9GkaG7yyZp5bwaidyYb4XeGLeyMamtJA
w1bZmpThiOaCsS3Rp5TYxC7lTMCvwjKXmlUVR+tQPBJu+TJnhVsDJT6++qJwxXbv+SsBptEQSVV7
VnVve1cck0oLfZCDZvvrUEE90SvdkUdA2vUYA0q/5mp+8/IKnR1NOw81HOdQhGUYm35+vDP2yQjR
EpLOcMynOxOMqYFtVK9WiGsrcM/2q6fA4kWTQmnyLpvOn4/L/vblWF2fKnm48VCoOs0GR6N15Ht1
yw2/RcXM3JwPQpVU06lW/9R7hpmM/WrM6Joey12ZEjIuNqxr0bTHR16ZnaLrZ7kxNBssH2yDIecL
mp6R6IrtGxw3TKM1Lii82bNg8DXlaBd3p4l1ZjvQVHbFBeC26tdEjWBax4wWElNYQ1yZcA8Gfr9e
buGNQnbHEno1v7JCy5nQPioHpgh7dhFSAukZVkVtoXhs//hUX0GkoZhoq40pGAvwpSO2B7Mb4tSD
oEn18VZqeSiYWJhR6jfP3aL2MVEhWYociatBlOeWkU3khxUv0TVX8K07odEai9cUGP6XC1MNNlC3
2XH880VRXL/Lj8sa5K48+8X6CJ9a7LbZQ+tlO/AkpH0VW6P1OiF/MykTPdjDAgvaLV6Y5WSkppaZ
YiKZbvoyJrehE6UQYbnp/nEPUyK5ftXEcvoXRSYVekKB+aGMOCeZbwli9P3D97TjFerWLGcyiwyk
iJBu6HlP1+xVv0odoSGTVr/+UxgiQhSta7cj4f0+S4lPxjN2mkuk91XFbNMY6SXI+Y8Is9+3TZSB
OA6dIaT3YHtfEP/Z7byuwAD5iPDRdEqXsBk47qZ4F161CvzRJMg6rRM4xMs38bIxStW8JysB5e7d
R7fWOwtmVTAfBqHGo9vefulOTC26dFX8xN/hmUy1fggssqYk8Mf1w9/fPzG2OFSnShLTUEssQtWx
I3MrSpQGHG8242Gh9WDl8sd1mgklqzVkKHRd+R0CwcMINVAhw8urIWoL22p9lj9pi0ZhMiPzQLjG
ihKDWxvMMZIItEiaSlrZ3QGAesEekGRQqW3eS1Pmtl3t98aqdn1qcB2l8eXZE9znsIgnJJUJbiaD
NP2i41JT413ME+Y1x80i3IXWVjC10zyU4z/P8pLP9rrb8WyaN3Y0bVjQkJac/rH6iZ41YeHfll7z
fwW7mYZ89/Lx77Xbl+Q098ZLwyi3PPi3qnSAMK6pRZt3vANIZDbofGamN2AU9lxg1g6VF4+Z6u9W
Iys0IcrhN69r7gRQ1w2LNQTtH1UImyP1RtyiKBYccnnxLPftFEQ4Sbvu+reJ0hhNBcXQIbeYtlXm
8N/L9vcVj4T3YLE6Ch/woinhUWEAP/MtS94JKKG/MLpOSRLQ3wOX6YEt/0RwXj+WvDCOHVCsP5GG
+hMuasgT9EjGDzUZd9U/CAM0/dSSrJyCtLscPOqKKuhOAXxYY/StlmVJMsrxOTy9UmPNcNtsSL2Q
INj3HbbsqFDrMjGpZbBOygwrZZc3TKiU7KVtCK6j0g7E8zPTk69ci0Le1+RbeDolDbdQ1uPWdp6a
M79APXCfWZVttxtyDmVq/3kKfh1f82d8jpoGcqptWJlKmAVqLmdfeH20CEiKeJHWDxGntqKxW3t3
wt4gmV4X9bEbl61B+rEkhnlq99WBb4lIAlz03agN+3fxUqatHkfYuWyJWE/MzBr1DVZh/w5e/6Qm
nAK7e9JCu/FODS19dGL42G9YAkC6TKQWsJdRD6jSIv+CvI4Q732Ft6j1CbqOq/LCyUTDYdKLnoGV
FwJcRIr+MhTzAIx6ku5jdcYCoD4YszNS36do3IiGFF/NiBb9QkjkeHdxXUpU2qU7ngXMP8HIOWY4
omiGEOFFn1eHo0y9rbx7X9AdlMsu7ott2JaMNAw6akkKVJrLkBNRhQcLT5JZji1FONaQOhKlTFdw
KN5GvA2+2363jTdZEpRqx/Vu8yHW99WPBXFNrjYQ5Bibfl6NGKUhB1PKE1q/ZVk8WIvjwNpPD971
OTYtxDB6dgdR44fNdiD57n9JytxEnLXNuP7pqv64vOagiWmazTs4T5IYxyk+FSCQNbB0Gah38vBk
gbmgyByDjtUqZ0RvZzZTwYf+jdox/IQJCB3Jya0KBcTXZaCi3YoqNGnShOGJ883ztVCV2jrJP3x6
qwCEkX7wK09g79RIIxfW5TgulYYAW/yPy8cWSLpWyMraYEItV3d7jpIduDsAkWx31kBI7kP6jP/A
RQpFL5lCjjk5zxh0lSHfC2gAguFm+KR0Uc6CjU+ph+UT4zXPszrpSY5ZqOLS8KTptcVbowN1dvCR
W0nW32CjJCAM28swd0KxwRpqJhJHdfrfxpV7+KO8wQs2XjPAm+EbvFC8ljRn3jcMz2cVO4gpHyN3
IzVZmIbOx+r0aN12od5FHNOCfd+tr07+TA9VkCBAW/Ic12Hm5P6iUzxKtlbl3fHweqghHv2Tn2as
0tmK0KUUV2uGNEFD5Wp66xPu1A/ml3BNkJdLugf7cNm0WgrxUiPqJ4SR8KNivtLRt+dzuVnCkFTg
Svbw09//CGXvZucbdUk+WyZHUVvHNE+naSbiPrC8GXbE1E5quhwMOj33SmzQQgPxY9N4jpqbOzsd
JZ10ZNtkrtacDME/Hos21+5Tv2p9OoaGgW1tnJH8zGeEk1lqyskZyCQqBbVCiiP/nWFhysOLRjUN
MtpKIQ/ej3zPRd+UeXRPJQQomyqwgVHTG4BckvXkXEbgFD3xKDTbPUuCzLL+Cs1h+rpqdK1gjTkb
VQ41zjJuRGZfP0VH3CYVXIRWXwTQU9RWX+12YJJYItIw0C4XfuNupzbxa100WjzAmLhWIKdJi4g5
gK/+cnMHHVgQw7XJQ1Y1C999GFEmUi7yvnqaRoXaRCZUFT/6bp//pA4qGAdYkSacT6Qpjv76sGGh
10ZoSkW5JEmnsVth+m43qgFvcg0TGXXkliE7APojsEgHFW2DU1QimZClVL6FRHBxzeNZv3JrQJrF
yDlqtSB7ENcZ3E6SusqGlGDpsAdwHelYSuHuls8509MYY6XJ0R+NQtxntbJSMd05v7h/T3wqwFG1
q7GidkzIeQS2a/E34zBZnrEZbemumdn9TK7sgRxFhxC+L4cZfWhrB5PERo6dOSimZeKVwzGkvd7k
nCx3JUf6HBj8ClpIH5QGG4yHCoAO3yfifXHEkIN1mXyBahCiPttAEuP3ifg2q8Uq7QtQa7XaMKdO
vntgQ7k4rqo6QmR0CpF3avYXSucS3Ni/qtHhKhe9fMR9tje79h7/M8P/4CDcFGyi7TdOMrJXKXk3
Zxox3N8FQnHmHlgGTbuHF7WnNWmlm9rIcrtK84Ywmcpg7NTI4uxTOV1My19T4Z7Myx4StKy3dNBM
U/SuziMb0d620w4WqobvhSmbNqy56meuIiivlTE4BdsQh7DASuoX9qkLtXPreVOwvx1T/1niL5OZ
r1b9gSei0gPue/gjvMvqisBwBUL5DX7qZDuBNeWHunFqLsDR0GqaYMvQTmGFxei0fCk2DPXdWAxL
brA6dlYVuGc0mkUX6/2cAENXpDV0ilppeKQ7W7/mqCMWJ7DhrBaoq7hUk14Z9N5C/taXXoCtT9Bt
ZZQy8swswmM4TUJ5MaK5cSRLAgD6taJ/V8nP4HS7EZ2JUAmMBaVKDiYw5EldjYf/VnuF/tlWCcog
xzFMYaXHPlrwF2H1Owdq8+V0nYg3iFv/jWV5xU1fz4lOnEXtgi6QPMBmncSOffcHEIBcjm5ld7fW
x8YWzsaOcic+L9+qW/xJB/5sZ+qDDY+d6HdGHiqer+fEBLyvbyeLFbLMrr2Ful2q2KTEPG7zbBFv
OH/Q6uVH4paK1eIIjMG2X5D8T5Z1tJEs3Ix89QD3hy7ALirX2+rACP18HICod4aurtfzNrYA1R50
UZlDB7oPFAXB6te+IyF+/beGRIuX0j/YEg/88KXygLgCVrLsmnRfQ+y+S2syD2uRvKtDXXQCU286
Yz9iByvQrvpwrT/n5nITGYRYFRkJh/WF1wfvgKMEnwMHo4JJxfoFneoH3gfhtyriZs7OLUBahjzv
1VHiLgwtKHsH5x9CkEidrci05IDrwrcKrr//US1fCAkidQbswVWM4eOYd5p2JgbcLzYk0zc/lVRz
qUOCi9T9zBtYtWqXnVToirIJN7RjevbrGwUMjF0tr2IgRVzzZ2sSeIca8xSKJdR3mSeef84U6SFo
w8uHr30oZkgwuNpCs8AhywlL+P4EfPK7blLprs8f9uuOzLxi3BP51Vl+sPOhZWXheSM3rswzaXOH
SzdOCfruX349bHvfEArnY/BBOnsoVlcrRqIjqcqXSc69zl6WRqiqXwTkbPXUimtnbarlXYbcXV8F
2adSpyw/cctmJPO58BuxZznX+iI3L3/2k+oDcqu8yKI+BkgWbULp6xfX+RHGZlKPPWGjpxaNj2Wb
6J8Ksygqiso2ksUjTjchEB6cPF2X9u7mo0/y1yI2xrGnNxTGRbsu+kAjuprAkC44YIbCfNqw7Ny+
mA2AyWC/8DrZLTGQKvlwOp9dS4g04o2gJCyIZ64yi8ARqNpfKEhSR8DNKUhNQNLAVawRmZIyJ2h0
xHqiw/i1T6jtsQDr5qZcsBoEbCImCCCn6RB675SqbGraA4/qEy+J+lRAwQssXji61+LS0B1pX/hd
7XGIkd0gEKpIm5TF5+462oD4ZotJuZ42/Cz1UKRSdn5DBbWu7JQ0USoqsamwzuYDVoq4E6B3Mg5p
4wtkA8zWFjatTF/PxzilRWp2gtznEL/xemT7N7+tXu7w4I0TbKHpQU+74KtODIOpAFSB4G++dtor
E6PTA2ZtX3FzQNYbnlMRII9IDI2/Iv0MtGjhjvwIPrXbJ5k0VKwhsnUsh6n9iC0muWbqA2bq3+8Z
N7jsj1Xw4KsPlGNCk+e6GyRH/kv2S1VpIGKNraHG3tyvjSL4OYkT/1QNm83PW7F2ZNHL51rUWyeg
GI5Vm66chwBkL7caFp92/ygIU2A6/NSvUklF6AA80AFK+rY1sLxBOo6V7qC/LuJzJR0F3WIDQ6JD
jwQu4CjDwEOJzgr5IyNMUWSAnjxe/gCr5zjBZxAZnYox2RivTEONBhV+Q+5iI6o+YcP83OvGFVG7
/ziCxk4M0xXFwHp7Dla3PO5GjcrkmGs7Z4rq6BNmamNPSu4DzaDD2+vB2xCP3PbJ40FG7pGan2b8
WtU+atcCoCSgLI1gi9KPRShC15MSUCDfvzpc0fQK0k38QOWWJ+Z1huQjb0YCJ4O+CSoIKVatIYGo
p1ose8moNKDTkcCu+4i5dJDGtFBqonuqFUSuZW8pMI8hoBpvHFEtN3WWqXTFRBtjCj62PsIMkQo7
4X9ikBVIMPex7KEGThIUJMt8VVcXnTazrI0klYdlst4GlYTCyQJGEvvZqIM26E1qaMGNbNyAWapC
1cNOsUbaH8RKrGlrZopidD56ghOzmsCAKZUd2QkICphDaLW0sHuwpfVmAZXZ4n7OlviUHGOft7YG
trKOtqgRuk4lTxc0XfqisMdRgLRFdt2z2SidIB6WY5tAe9URrWvI/MRev7dM8d1BBix7dok4hII0
yvfSc+RBeLbUuuTOafuKwCnKpmogP+pEcc2l3NfH5qrp6JPetqdRfqOZ+zb+XhXriEWHrHES33B3
ndpzjZ4ET6S0742kx8oQT9uOTSLCA1DqF8KrwkxCzuOYou8a/0CcMZszX7UN8XNMR6Vsc433YUEU
rxPLV+A4V+qenQZ1NHUPd7E+RPRP2/Sfi62Cx/FvUZw0jt77pQkPF6qmlxrY4CDTpqEVmgmneq4B
JlodSi9bDqGjT22PaAGfkp/Fm0SOVFjXRWP2skzsYPnZ5IiCjf7znT8Fuehn2lBMgjFSeLCowSvX
CE8icT66YKNkUMhy+MlAzvjXp4DAFNdHlYHgwhO8+NocHHS/T98zdIei0p9ynYfl7KpDhAT4s3s2
QLlqwdr+mZpXj74uzEqNwbi5g4DFgC7NlnzO1W3cxCGnXQJh8cSICK98l43vvJeZQzNiM5N9IkZc
xsaUtZwkfGMT7iAlUzikvyPuxHdau2cBhVypbAxvz9nyHS0x7xMs1bIwSRBwDgY3TFkG34YZZ8iI
pV594CnRovf8a6J1gZ/0T83y+2chjFl6FYDd24xAiDZY1K643Uu/WM8+B1NKjq9yNnK7IejZzqFx
VgL0Dr1D2I8kw+on41h4/V76Mn+ibP7ddzKLMuA6UgMfeckMzPzz7tAJ5KQQlk/eDOSCriD+arIS
WMTgsPsxAngyJNVQgBcZrXmp3vJ0X8Z+d2SYb9SCMjHDznXgGKQKu7jdX3rxMHBncKHcZTrniMzU
mwUDI7azfUuSBGnbtEhNe3fQFzeyUBr6LxwBdsLDdgbAitj8bx7g4/KavkiiFhNxL8jgO+r8XUnK
WpckVh7LUrx4uqF6KuU4MQGhJ0G2TYeO3gf3huo1t6r0VLFo4D6wJT8E8nx/nhQMtGFD4HnqRydl
f/MQ+/mSFeyKhheQUAEJaYhqHnPnmTBDg6u+TSp8XVlWjoZ9Gk/RI3dpkP6wXVrwq8te29M6fhWj
57zpPKj5jE/CG/chpgiiBmSdT44PdWjhaDdHVm/iMU5syVLn+gw3iknhAMRf72W5lV3kNjY2u2c2
VgAgkolXjnM3DOwRv6rXCQ/h6rxklWeH0w51/RenxDZu06VD7Jax3auB0HoSlP0FjDuiXbqcxpaM
QKkSWSvqWPexG44cOrLsMET6jHzg430otqLBgooXl/GNHBY5jgnAJlAqfSvfnDh+/mzN4O55Tf33
GxSbu7NYyUs1KkwSnWan+IqNI0zOBoE2AZ7Mlhc6bo0epAFr9gIhdhkimvR1rQ7ZMSxW4ruLjJo+
V37Mz5aLI+S1FD2BQyKOZQh1HvHWRTXeBAvCRRI0GGTv7SPe9Zkd80nVY6yASVneVjAereNSfKNN
GAjLzsWiw5pvn0u4TcIUcZC4xMTkbM4LF8DbQvefdGo8N2SEUMFnGyzVVl0lU83lx0mD+H3RYrEy
Fsv8rNuPxaxTk/ctW2uHJak0QgJY4Sdg64xVYO9uNBno4mqtJHi/ky/fCwHSNx9qP1ZVSMimVV69
My7y3Yl5W9uHMkyXLbo2R9A9W0czGTQGsmHb+K4jM0K0tZmbtYqLbewjnLgHbra85DZqbx7S/u4/
JpCXSUSYRxDHwkkJMhiquRhLMM1ua+Ozq50gUcl2NYs7G9R5sLmdAO2x2rQDHSSlLKhnsXj08aar
Du+riwSzXxusY9GcE79WqnorhWt7LH76wa8jfgepIXuVtrtEC7Fzyu9Du3AdkHLHH6XdGXNT8oys
1jml8O1ZSkgct+WQOALQc0ds6kHGwugqKkQKTJs6nvDxMhpuSbxOafGHGVIINDix/vt72kMNQVxp
VtsIl2sZf87NYsDiDZvO9VXK2dEN+3SdXGpJtztrAFXHcI/hSx7SVq5HD+Rs0SzCFKpNGuAESzX/
fRzjxE1yw/6dOc2qQJ1xb9aVcyHL2CvkgrKby0DQr/LgWS8/ESSG53iuZ2ecEL1Sfj4G/SAMbfR5
WjNYoEP161y6QEWfmM0L/H9inRkqDoharrDevHTGu5YXXms4pNzUEY45arBrKjgSVMYnabMaeSIX
vNCBLOlgYK/TUKfD5keqGBclGylVAKyQ/lQfYbcuFlPUdTnSn87jVzpqKhK0CQrBFMJlKJDG7e+Y
uKFCTFS062b18qxIjN0a0ObKieuTNUgCd9RWUIu0AgajfiWpIkiYwUBMdratXMUsjn+n1LgF047/
XFNFcVnvf/GEz+zZFG/gYFgAqLp9ynFTdT/48kk/BMr9HjJCcuvEPfVyeRrFp9xpvziDpbi/5Zkp
OzI1t0WYgyQDSsTVYGe2gVZKi5WJ/i+tY81LXL22eb64vGrXBfYtm4Jc9Igx+J0OXWs9PZ1F07ga
z5HvoGSO++j3AYNBv0PJ+zifROqRrZQPWi2vaq5g/+2n9Je9veh1+qe2HxWaF0GnGW6jpm3Mq1SL
59yB8dTtuy2N+MlPHx6eryHpRXwEs1SqJcEIg7vLcxTIAL7xGukB6TZiDCPxm2fkH62cg47RTVzC
8byOdLp04WFyi2kF9s4aftSpL/KZe+ePO1mbo8s31dvudMVa/PWaBhnFwZuLpVAWhjCkCMYGpHev
I5A4mT/glO081FKn/IMSdNXioruy88zUs4z5yG88sPj1WjQOvLqVLgb3/qbMHhIgkaFr9TZAfSRt
LdWtlPmkBCltvdVgmdx6GEY1fb+388jqPDxFqGBmoDbhNffmQxlBwJDilpBh7xr6Lo2YQOuhdn/1
H+G+Jy2W7r0zYgFpCH1+GPT9AJ3jU4jmJ/uMvXGisHSgOlOL6wOXSZiB6FwMTT/D8C02Tm+VTT7D
5TmFuT1AMU9MTVBIZcHFPImQEM7fCjQH2i6/+uw5eVj3+lECer/HTNK8E2qNYeOq1IvuJ/UHXAna
/77laR2oNSZqUCzNp1WZHxMm0GWUt/6x4Mkgk6PiKZAXzKTZONi4MRxFowe3LwLC5ZYK6Syl+pzW
TxSJOXghObSkKE5n2zrVvO5+nsBmu8RLOKcIYT/OqXUOnvTHoosy/A8Y2xyPu2YCoEzRuqM7uwgE
qcn8evvVujMeD2bAcBSM6c8ZiNA30awx11SaxUBS/n94SF38fQJpTDcuKFoGnmPDrtKeuvKgB7Dr
iOuWET9DYfCqsg8IKwmPAJ633PWQY0b7WdnP50zwpFQNk5e8Z/3gKR9t10Q6Td3kL1tlQu1BvgvY
c9Znd5TlhmrWr7V/Nqs2rwSuvxS7vVxB0Uyb1xvuGBo6pqoSad8iEYkouLkzzISr05K9QQBGXCBb
faYdf2VVyu6NNQma8dZgYsvmMoJTWJYU9DQlVR52tUoxbstWbgAUkceHDLcWaINXxaGudA1MRYYV
WiQJie5VXpc4kHnTSWul3d9KUpYqGN2vHZhbdfOfzQm5PBLred1rGHRtvRB5QKDQFb+esu/ou9PN
RmBg5dHN1EgS6Tu+kjlFgzX5A9wjL0jizjqybQaKpDV/KcgcAQTsQ9tYGkxkkM6+KjXKYcby/Gr5
E2KSR49AcPYUdAPmo//TtTy4DoZyX+OmYoSFj1n5KT3C6zMTomBM972iAOqnorrgoJR1hvYogeIw
NqJPsgHzgxqORRw+3YOhGr68xoFtk/oMaxBQbnFmOmWiWSknzkmesk5aKTA2DKM8VhXz4YVFo63C
fGdPHxzVhE84Lqkoz4TFTMmxv/LlDnaDgvMKZFCKdTUf/92x8ofag8P3FGmmbjEzZdpEcpuMby3N
ym47nFLM89ydAnHkl48nsyqjJtHe964qLGM7s9eZrNNphAt1/HPtcEorX346bohrcShv+V6059tH
GxuFBr7VECRnsPIA1Wtv9mTYP2AVXishCUEAu9tbG1tiwALR4A+bvNoJBrmf0jUMMu1RkDyC/i38
gXLLaZ7vJBRkQVnwr9AgK63mbg4tVTcVLM6WiTyH7jtGloeX23boHOgc9TZrUEAMVK2I2BGykTUb
1QgE/3Gk5DL7cN4CsNgyR5IEKKjlzsALY9ty/4e0WjCffdSLpwAtQIjQ0ep0frb3qN0z/5nTU3+9
I1YAgTUVV9bniR0FERLmz9m8HRA/sMYyoUmzfFq5UtBJSOs5cyrYmH1QwU94YFKe5CoSOKugtRej
jwUAU6hBzuoPWPSORSDHIAs8sBKmsUIET7pgZDQTYGF5csJuNBosBow0RZYr5XGggCgC39JW81zB
JwdwI9jvubEtRFISRcYGnBl6AfBz9oXQWN0OEAyva1LAjeQYzDyNJAYMKPgsgtnnjcW0YE6sLwjg
jo+QTHgwId8/jaf/tiTxDj4DDRuHWiWx3AN013f4qQnjY+h87HQNOWPcDKIdWvwel/Bq7BAUQWGU
f//mPENun31mMw4qFrKMq8y1tYY3ynjOBRe//ThmHUKsJMPx3iwlEisQiNZYip/KvL6iOQxxkjsy
TIbTyx0uO1NDE8YM/nLSz1B9XxZCM7sLOzpyqh3mCmCAb7jUXKVpISU9oBRRs4iZq/piovtyJ0k0
Y6SRrGY4I4GBhAcIlUoKYxKgEXNP28fLnMjUarrAgA1sBKKn1wOAKlzDVzmkaRE5y07hQBrs+4Md
1Nx5X7QEo/NEjFg9I0kJh/0wuR3WoNse/Z3pAiD4Oe5o1F/SjzF3k1cCjFQIcq5HH4/Kjqo/hrpD
wdK1dPVSKnkd7Spz7q23AyNNefk7AEqjlyvm1+AzcovF/OkQ5g18GCN1BrfETqSRgP59M41dcq/c
GrnLj4QgGrMK8A5YdJaThQnjVYBffbdJ41efE6WYRp8lU80BOB/wE2f/QO5xW7caiRRLMRQbrA0B
tGaPNbBtrQuWF697/RlPy7xauSFyS5wZjcwC6WRbxUCBWsPjAITcJILzewMFiq+dh8wSf5q58geL
mYBwA2d+pQUSeMb8l9TxmYLOoywNw/yHBZtZjG8/aQkzfmm1h7TBBKtxMOl5iAyGnECByky9UHGL
R7RORuwLva4njKhKfZtib1jMjWUmbjYCpGCHM2Nq9zdPU4o+91xtjaL1qvkSOcIpz/1WjAUkW+7q
VQOCvbGMN98p+B74kQOqVP5UzMKXIUcZWf+uRBN/9y4g3m8vnEA+pKV7mknljpw8CUFxaHJv+HuQ
0pvQY6WSezeDwVtHNGtwvqIVXf8DIBielQdFpF8fjqgiKfrG65ILU1UWCcMVqUnZApLZXvxPhNoX
C/k1e1vqIGA6Ds9kIfW0XA6BrKs3cyklBi0JuVW5IO4uQhNB/wPS3em6lwbMt7qFjjY/lYzr2gpN
k/2/LVsVq3caurCVwg+/FiEXhKc4IX4D8azLQMTAm64tz2KlKnzCW750a1tXS5FgPrqf8gtfQ/a1
PMqVKa5VRYVvRhiYjq0D1kfP6DEHIDIoQfid/Oz7kogdtzqvL/bbLY6rOdMhSSIh5LJCZ6AvrmOE
HNFYeVFruO4l3oZaGW3B3j3/kngUnF/B6+ctQ5VJu2bnPmm3pEVZwo1tMqu/Z4XtLEJgagCpz1DU
59InWomd84wP8phyMVNYJLObh9oF2hiVa2AprPm9APQ9YfPhKpMrDvOMkuOmsYQ3MOU11aYytN6k
fsJmsES2nCmfKnfJeA0CNH8kGVH5/zrwJwvCkUpdRLD2rD5VmzhFzPXmMsTByHAK/Z5hIuTuD1uK
rs2UcpxeCrcwXagvh7sa86VtolV/6NGOAbLBej9fCq758SkgzW7WVq/KdjrnDz1Mkuwey0ryWOdp
7AiMW/auxU/69PnGRef9/hocLEzRK3Zrqoj4DTnLp5uq500JMBKDn8Eq0hblDrbHHhob7yuY8z7Q
NWaxgFLJeQQVXxd3dfmHs2SifRI4H29ggVOtGTv/TZhJhM0YexAPUzWxVzrZIzgqIxouY83PIcYb
TveyfvVIXggRejHqzfnz6HHJI0iUlfyUYgb5PxfrGzeR5kPcXp3pYneMAxBipNA3syngLlmycB4p
ab2uH6ECaIu2n6i4aFv1SUduyYK2G+TYtTJwMpMw+8I3XwR4UhmmOOSiMemmBlsUXLzIapIqgvJP
RxaIk08s2/WHKkjqJSbfVP/44RFsqGq0maLJnY8l+EmkLtH9ON9DaD3DeXeQZ2+M+dPr+XedSpx2
y8nYFRIuil42IeJrngOE2zT8yaCNgNIJgK6+mN7aE0ySYWNwGoCUP36nnAf3ZpbjWAnP8WzXC1fu
4foreGNdioRtc9MRq2a2zKkXGR11n7Y4iEsELwKfZMN/wYEPbbc5/Ba7YOp4+tIpNrXZKJD2H1gi
XOkQY1Q1ivdo7yc6tze5IJKjzpwr243lS0lM/tva5LKP93BCmmZ7ySgLr+C6h2bTGPSXBnztbbmZ
joKla9wCgzQwjXWy1Jnijl2pyW6Dq/qmli4CHn+RDRCHFvKSEWez30MHttBvNmaxBbrYuC1QRj56
ck+P5eNHdlNkIl+ptbP45OEG3GF/Ml8yci/rC7jhUgTSlbAoj2JELaShOpl1fBW296dhcZ2FEz8a
SinVGZODw9f5WragzQ9gXuZos5r68/3XapUkL3pYq2Qf/ZETjowvykWK6hs9Zdqn/CLm0LV7/wd9
6N7AtYpyTdJWUTsAigEhpUPp7LAv7K41Z4cRy56/jm+ZTY9Na3RfWsZhgmRZIyuw6qVo8dykribF
1yR4gPPx6DtTch184vjbgpW3i6xgPE12lw4ZBxOJnOcGY4gvO2jzFLSRmSizFVITfkEFtJXcF2M+
TD7G3PGvXa9XwptzfCc4WEBjjou5lmy5iAXgYNPphslcPU0s49eeyQb42ecpY3UNpk2V4c2mwQdu
NXNgnDp1mYCfxoE0s/VayJALit7c+/mmSRXasIRY39mH959+ThCq/77AZ61WYwYc6Ut+rLTOTncA
sR5PLjWkPZD67UwonkZ5n5uuY924+rg8QMWHa5RlBJcx63KwlPs09MB29xXOpLJRlikBpiBKb60F
CACkcN0wq7KsB4tpnZQUKaW02Xfo/byjgHqBZlP4oSBTquXxpp4k6WYC7ap9iswbQAcdIjr/DYkT
A5WXOelJ5MS/OCx/iBUsDU0wpDZ0TXdYkQpRS2uXfCvcyPu4TtwYRSmW4mJo14H0DwpR9+ekbrnV
NTz0r2eH0L1PIzGi8n1ZoLEYzThwCaVUUvWZn9BWII/lcFmEcv5nENXNePqCzetkHVGfhgi00sk0
jmCMsTp4zOA5ANKA7afCBz8zmGVmayK5FvTJZtkM8DSfNAwxvY5PJ6YqhlNGpWZ9yUq1xVg9Aul1
YXpZgcaag1AMj1NvQM/LC6TjgHAQSDpsev3bWW9ry/U2ttBhdwS8r6k5drkElax9KIi2emdyf3Ua
jM63rHLQ6wff0PMe9sgp23RVdOqbrytNAZ4Y7dUpxAG2X1wGboxLVOXESyujyuqWgShOp/BrkM+3
zIAL/mgWMjD8rv2n5GdrdSOVocGe2yjxzo/0EGJ2rB8NQvT8/fXEGmQ+h5UB5ZQNQZF++tpz3Hq0
22NNXAL0ne4e+EkrjW7o9TpzVrmpNKk/pzqTEeq4gQDxIvN+GKBVBlrTCoU1Z5a5tZyiElf4ynaA
/2VRDyx55wWdH+hpOeDaK9M5Z0l6A2N6ps+vnizW595KGN2ns9hL/b3RU2mysGgLi11canhz+eoF
KkLZg4ExV5c5nNjoVSSdi3mQJfaoLrk9v3BRcbTXZp/PjRV0fdPv/QTL/7eL8HEmtXqqsDy55kzS
UROYc4FklDG13qIAgQfg/XftCmZLwHoL+y8XhSpZaELt1Y90FIPumR+TG2Og3p6mOn+iDOELyThh
SE7Unue6iV8tbKjfBYbFtgfvBeGZUbkv4dGvVt1erf2LZ2dwYjMI33V+W1M4nqqCvvjkQxifbpBM
Hvgtdv4FDlZ3VH6rdrFCazk1qIPTU6Hj6hU/EgCSY7Wub/sPrAKxrtUnqowJHwW16lWa9dP6Fm7r
Hs7B+losqv9uGu1fIr79pGseMIHbXN3p/NzRjDcg2x/OdFFI7sOPD9YmoPyHPl//aKjpLjZctAfg
S2QrDVkoNva+iIUvbZCkYyu0EXCNZ8+jOqvVEVDlzogfd+lE7qu+ashxRv87emSg6wZXM77bW+Cy
TDtZZWWya5EAlE5MEuAtbdBvhqJSe1x3rDqN9BJ0vex8KBT+psV6dr8mxaVIxynbS0vXPZ0kq2GP
xVcYx2uNRdT+Pzok++An0uWdkVknSamh/RLnFZQygx6mEmNwZFAOOkwirGDGB71NMGyAd3IJpt2u
89Yb2zA/iZdE1vJCU++olEi+0usNwaDqkdh01DaW52xtSIKaxAhpwIALNLbKpsZq34K8OSK6gssG
i5ca9se7LIUU8QXAyZ2Yxw8u8ZJQkpK7qIurT1Ru3Lzr8NIJgA/qxVIxtx6mWaO4BHrIzZIkrNy+
YKJBB59I4mcYFHSR28tOWtEjWj4tqiasUMYiUZADiDud/Lf8900MaaiYUFXjRCJgU7zD46LSTOMw
buRHH2n6sYTz6Tx70gFwXolt/iMbmtqS1vwf2jeCeG0LQy5qU68tLW+NX+uhLTkW3/0wIQs6fVtA
Q3+imAKVsNzU2m45waxDsE+ATCxNTyqhIIHXHlhy7mCHqPm5WnqcOdGq2IH03/SwzAsOF66XkUem
p/CHATTzYfPTGHo6NAruOqS2i6SXiw8bM55nN9ZwIOVeG96oBtp3EAu5rnaM7pqhRYiFQAxJxMSQ
2nFG30PENb+4JrVq16gs14HvBUyk2p+W46FlPjpBOEwLncSSjzzc6RjY54K3x+ANUBv6JFb0QBz7
DJHopQNCZ02hF7S6JBEv34HCOU7BR9vFc9Z4N76E5uFzTEBu+46xNEjM3BP+YvfUpUq/uFssV+mM
A+RBHv7sZk2v+zXLLEHKqp8Q9AIDdPug9Qp7f4Ze6LOBZqcLfhkA0YcvxwfGyQ9IT/R6zNn9IzHK
f9Rf6mTy0IOakhhPZCM6fES/cyXxLEbm71A0ggVCChSp9aVrYSZIIr3kdY/Lbs3FqsO949DJefnq
PD5eA+GnhaDGmlb2iKjrKqTZTKmRZ5vIKYyKqwVqvOthLmwSgi7bf0ZVCcbx/ibJVCsr/e8n+rDV
P2tzJTQQGpEQntRrKChX0TH+Yo0l3+6QXdUSJaomdjZnSdsH0fgKE+SyAKrZlF3a5V6smiOF4Qos
n74DyrWzQHEvjiIVbadgs/kJoGoFZxKdyMJY1cnYlfTHF1ljN6NlbzWw/jmEntvAk/Kig6OghfyM
83eekSv0vDARFrPeutwkMp152MSincyQ67COQx7hNZAnHJ9gC9VZtQrEQgDP8bVHDVFimDukJ/5p
zYv6DS5nKVCTtks0zBeeA9oONB9z0LNLkuB7xsz547rl9TSm6FZEhh43h2UveJ3VFHjAXem3ECGk
rt4QVkqQxXHZG7c8ldXaGJ/d2SmTcDkTea/VgQoSNpsInI9OyZsvYzQUXlJ0RLcVNzsO92LT/ZLz
xTcgAymzT4C+qXd9+b15zHPKEKNFQ8sVHvi3hMaxOQvkAzqYe9I9371a6GaSHP5CGeugrs484j56
lC/4l2RZ5AiLmzYEJX7kZaB71TM3+moQplqYNlnjbvBiWMt8Vt8E33gmOAXLL6yOtJR1c5zhsjOx
KDEVbck2j7cE2Rwp2fxmzwsaqnCXjUBlfD0yDOVLOOiBhNMPxlv78edXJt6HZ7cXLMv3sh3X0BBn
ptIcnTk5zmGoTO9we9VR3tXocidqiFXhhlrLKR69V0tpl/0ndtD9B/B9X8EcjhgTGItd0i4pAqpe
bRv2WubH1C7eRdgiDhE3ccMUyGTxVRiH7Vu67ibO/YOb1SogjtDOIP1tFNvL22x0dv8rQjEptK7S
x3AHtaOVGZRywG3sVZP8UgGOlsJW3XVKGw4D2vdnbydsG4hlvoiEvNNX1OO1v2XUAvqyD3uhMFo/
XppxkUQRjm+FYHERfRe9qNFpC5eVCl7IvH9WyosloCL+qzw1ekwa0xKCVMJi9+Tqapblm85Q3YC4
/296h4ME2M7O8JIsQogDt7OXdRuoGSbhDVd/K/jcCW6NyTnf05aY0zuQffhCs9VsYeg4xEz25GTm
eENhI7aCf3pjExgOqVtAOHGo3CnqDaPLLWamef31YswgrKi2dG0DLwtKFXKgFNaDA19spu0lHiK9
ClipIw3lPzw+xKx+mtZL46XlS/Mddgbt5VK4IRA61vW9HVpReMS3PjJl1nc0JGH6V36Qs4k1gOxS
FMx1tRfZgslOy52ac1N5UXlrfHcmZtJYyNPMmyc8Hz01T8qN1W94XqlZlHZz56pzO9bnLl9L7U0C
fbZ96QvedVttxo81qRNrd88B9Rw5y3nFEawknajzfSZaHdU2C91uZFJWJ9tq72bRkxWOHmbL6v/y
u0g+554OOI262WHsky2MJ5NL7/s7GE6I0at04hSWE3djZoVdGiWN9Gmwzjxu1/HEKJwI7BiaYIB5
BjP9BJZRgSoXgsQspu+OcNY9UKgY8YC2Ns37KjaO+76t78k9pb/xRTlgN07dPa0J7qfv3mMHK2Kr
fbDZXhYMPMb9z1T+ZMt+KHsKcyfrzGBmPCtGDg9JkpZp4tFQYLl9+t2Bl99OiXNJfFx1Ltrxuuhg
P4ekPVG5QLWBlumquLwizlrUMwdjlOng0zHypwxkQET6VbDK06/IbWd17wMN0UNZa8SE83IzG73M
jE6wwXHFUNcEOv2fAFNhe9hfVZ0EF+UUlkJZeWVUVStqlQhN0QxZ+7gDKxuK96R/t3tqJtz4pAxS
0mEPnfPYgx962L8stzoA8ktyRvfoEC/dCYCQn1Gz+0iEcaDm3ceNlWfOVP+wVs20OWDYmwO6gifx
dIbpMrN/TbBPuDXz55NLib9NODjk0zeOcNvRgQUnQUpuP3r09eOqZfx4TO1NlMUFGLGpjlNLYjgj
v15rpDmFLasKRIFdeboLg+RFOLK7fRb8QoBlO6/1u40kkOnmWl/YjUMcjXJbvKgeQwzry/PGG2p2
vrLrp853vg/jfsrBPYiFuJM77TNLWZvDdJjkGsnnwr2DhIUMXM01R49Q8Q5zw/0EmfNaMwqOrHro
iEojOb3dcHE7nyOXClaFKxMqoTCIT3aZbgf2W3P2ApAzVTDWf4RC+/4YBjYDf/SJr6TaCkmrpl8I
JY3OLGZp5vN00JwaUW3MU6D1Y4Fo9ceThG0iIlGJm6ASPZirCquXmRULFNeSTtaYCLb2pT/BOfW4
8OFSRaXtoqChXprcMiWz7xcLb5P+L84MDMYoVBTu9jc3wvZr2TGVAHrHg4uF9Pt317NPYB9QkxCP
i/p+IL4zqEm8pRU1iDWdU2Kz1552GyL9ueAEKmMyFE/lojK49mGr5/uQjc6g12zqC3zn5oeJ2uO8
irNZ6C2VNK7IjGmwBvB+7RS8T3Mbi4fmC34XjbC6JmGkak4P8m+rG7mf9/oEUGN7hgyoxTavA1aR
i8U8tDdxHZsrbDzY0WHhxH74IlDEdWvx1M0pSm+wCDw5raXRcOqj6HCxl8oB8eXk1NkbIX+9Ni/D
40piK6QCLHBTNpAYTLZ0AvFhO8Zx+qA9N16cpRp6PMDBVLl4Ix5Qfxfs7oWMrvdnQidhAMn8z6gj
Ypr5C5s11tWRT0SorskL5CG8atgeb4wmV/DtJyh6wgPFjENsK81zv7R3ClqyvEC+Z73DOCL3S1A9
OImlBaO3vcE9iCHybgd0N4bfhOo4dplQdb6P2q1yp3137HvScmYcERcGdIV2tmo9OKZcLVPXJPdx
q5djM3kjsJMVsKCY0CqgZg5kFhHaO/ug/RPUO/vEn4HDcx4mqsidAGt7S+8s3HQGer+F5yHN1AQc
WvfUjQT7aQxDK6GN1mW8A2eq3NT28uU/cBleNNrCB1MQbM4mWrR2/Pke6nAXeqmM88khzj4YTRHi
HOQBh/nHVZWPBK2euwioPbF+Dvsd0Xi+9+Kl5mLBiexbZS5AxuJvkck0sHYA49sp1eJBj7b7sgM8
gphPaQdq2ISLTbVM81EN8FpGRNwlMp5yuziET07VpM1i1LQw84omNaTfdmhwQa0/9SA7btERoBlZ
RS21PwHAE50w04iZbqtVJiTIImga9tVnIAojQQfwAUUvXqsFwr2zemoTCEmOgqDSIhY+cylPpMFG
Cigd6VINQMsCOi4ush1cUEuOCSCH9EiJKAc/tGD1XwItSxAUqHQYp00VPaoFb05qrCwNhdATstIr
lkSMvfJGCATPiNl/rlgfagMWmm/PW9V1uO1WGjyZamaqonoo8i8JEXvgpvQFg7MTb9+SF/s/UZKZ
EBf9/LVXmH5hMWWjeQVVTZRyBNqI5V0h+3f3Xejr9DLcyiRsNN96ZzjV38HXTVCfy7goNHGiQUCP
Jht6o4NVW6DTMG+JjnlPSgW2pxFvyavGWNk8GBzmTBsyP0/6zS8J4pEgOOO7tE33z+qmGdol70R/
zNq41HIZ/19AOckBL9t/68yUwU9sKdQy+ymox2HJpE/5Bdtf2xgAkVBKTGDcTLr8CULRsa5LfQ/S
lOapsLIC7HfLlxjSJvTwMv5MoAyPF95ixwwQXguGYF7uFEq49YkO/i5y7Tax6TanyyeyObk0MnTP
5EPfi6S97bceMFKq8gkZLHit9RUQHRaFpgHKzWUu3NYSpfmYLZG5H6ZVWHOAeG8Db7ECo+P+GpVD
VzYGxsxxVSctk/VUPY4Z2JuzE/1KoYHJoUy7XNiw4WYDsNGcY4sJxxEDEfCrwhpombD0yXKjfjUy
y9UvYehqdeGIi/xMKnFyibEvXt4nl3FpoDLzn8pIOD9NCeW/M69mT2JzoYAKKV7Jm5cSXehIFwet
gKfZBNLsIgRKLxyegWN0fhEBa5JhB8vU4M5AscV0wH+x/Azj1Eceglu+FhpWYNm8fHJMtbY/+Ewl
nPgkUDfbJ4mA0IaYfeN3kPNp8DdwVQaZWvhV0O/eFDSwL+GbQfx372mgM6LRWrBxRfWx7Ed0BW+U
IryI2wLx2abx0BEvXAqKt5EtDjJWnSiy5U+gZJ3DA4DR+sQJrYXPg10Ylv+GAAbbkLajP6xzQsNL
0MJYRDjFiMAx29q1Gtn3396ychxrmXR50MP6w96TZWplDpC9Qjb9yBRQwYS+4ZFokE991J3q8ayF
7Z9TJ9ZbYGP6MGSHY+uIdwBAfvth9ImFFRzrOVnZDFaFK+b0PzAp/2NsPqaLEIRAKuv5/jtxYEsf
8TXAxwR2XO7dS5JzKoOyGJQ8OF/t5dFuPPv7IDQ8PY+YGiCVslcA1Z+S4DJOQuFzEqiZrr+vJ8lp
8+bLmwpL3GR00v7uDM5lmOYdKh3m/uv9TsFL3UXxKiC7RWt0eh7F3bnKjQMR7Ag2k+x4LeUxfLII
rHVXDSyCwjUW7zpqQff4xHLywtzywqfj+81vGJvv52y2bEp+bMeR1NLHPFBc6eJIWuKeknTDIq0B
IdKatSyn2xeOfOHm17tvHTAq0Z3BN4qJYmqa/n6Fd2gXv0lWqN7dtgjv9VK/GQY16fJG2v85d8B0
UpF7SUmFJDiodPIxiLx2DzoAi3zuE/Y3WKCuGR+09dok9fGE7X+OWen+gb01P9yJf7kilKkmMLHY
CCSZ9KWmqwo3irJLGdrXICm3FxCY6JIdKNhfnLvfNhSYIYYqL+DlIiADM6Y9I9XgeyZxm3rfdSIc
hQYXb9yrb0gBMiprk5oUFHy400Lk+h+KNSeQT1+ocGF5iyD4cJkxD+2lceoBobJCe6DK3CLTgBYX
mQOvxSVQa+Z8l79O7MVKll0oZ1IQyx/Gdh95xPIMxW5zG20/mX2F1eGa1yHTM3GpP0knpB2R4eRE
qPD2naUlla4OshsfdoXszctbo+0L/uGv9wCwk7RvpqTez2/zM44n6ZYo8zpwFoEUtx1w9AjtGNu5
Pemn/bqJ0ylcG07qYHyJuXnMEzL6ttuWqZHsKcDlM26+TblqPMCu7CMg8164H4vO+XuJ8eyEXi8E
ci828oIG/RXj95qZ+0yM3ISsAVPV379VJIAHZS553dpt41GOlVq+F7C7Xw2dESrqfc6MgfK8czoa
OUhfSxwd4qT+skO8tR1Jiuv+Ik0snhniPvLh0dB58c5HeUX3eD8UREW/V+59tmX/3HRkCsJ57Dvd
vwuBbHKessZVC91XE3MJeaJr5KBzqfMD73FFrW7PqyvR4qppNd9tOzz7EdHeKmf0mb0cXQOT7SV5
Rlj2S4Q1p3+Vq3zq+uY8BsFWe8rDjRFuYRz5CZRDnOLpskl9qjBOV/ZtBSuCDirbROtgchZB++ZY
xp/3RyskBa01IRjJC62fAdIQvZLnXeKnjB2MF0zOQps9tnjF4j631LkVm947Hu+dxNMM+paDla/d
w6OP50+imeLZjfh1RnutcS0IncQTF5xcvo17MEXjPWQ/8WgM+IyP2Un3jqmudaRRh7Mv4TWsNINJ
iGfqrl+rQXoIFYdUJ+PpL6QKvRSpimaqUBXa+VQK5IkrW5jfeZRz4tYEmKezJFph7q922VfdIzsv
v8UQmPj9lL4RN+j2q3dpTBPzxiDetf88Y1huBKTD/WzYIQdhIJiLNzy/qpXJDDYTe5qQzyGyGbod
NOGDzooKLI+arYmnnmX8Y1qeJ66QYD+h4YTLKzogCyzJSt85/FokkP+zHFNU4lu7EAEKs+9r3w5Q
TJf4kjLjkWFwO/+RBqqgxKhoqflR+4MKwtdxaJZV8G7pZwyBqM61pHfa2F6sMonm23Rbsy3DkSfJ
Z3MDQhU1lHMZYBJmDABNbYezL3/yQUk9SmYwVNouKmaFSbveyWlVUU1gdE11iPvtmhuKpPLMqEV5
PPE2wRHtRyUz96SodwhweWvbf3oTUQ5rpnN1i1nk+jnsgQFsk7ImwRamkEolO/Zu9vjxkXqnzpjS
Xpl4g6uB3Xd7cZrPkFp5p7txv6IdSn2hzLIzMu5m/30mBGlE01glmhZLS8LJKwuVpnIVxHeFwc0P
VL5LNhfomX49k00s4+5m/ZoTYb+O0CgvQdVuOdqV2ao6qmjLIZrvPO0EDYmB3Pg9Dd4dtR5oQmWS
OYgdljO79oZiEikVLCw+Q9tOy3AAzgINpJrSDL2lX4TlfDa6iW8b9il5xNXk9+9o7osWSbCRhsGo
CxmtfgSFtEv2P8QrzoQqv5ILfcfEOHvC6HkdndJ/8Q+nEYiOraizev22jTgdGOWYJer++t32UOZk
5ffU1GVmsoxTZFOr7cCpH6c1B5r6mdfRZHE5Jmb2E6ADNWjewdPVQxUg5QOW2ERL6d7w5vQfMpQx
dx0I0f5eMyX7hEwzvd04u6HTXEBRq+rMhGdqp8dygqU2JuLOtBA/oB7HvRoVSdV8xRQrQyCVufSX
rua7OFG5dvLHqV+RzA8lGQ/oKWD6vuJo2+agfqR8kUm5ZTbHM2xdCxDhi//cTZlgnaZCzY3QHu1c
8Jh3+A3UpZK/KUR0FegzVXHw4UCf+W72pne/Jbwsil1lYab5N3I5XucQgRwjrWP1D34xJ1DGIFKx
UyWMjNV4ATK4WSA9TsdXVWliha4lAce7Sp4OkU3YTtankcjizaXs2AEOn18F4+uD20hhsHU4hgz8
Pk99Lu8HDSi7Z7/tbY9wyILmBl/+jdu5SaFEw7837NWnC8E3fJ2mk8cSY7xMGMyYuOj779BZ4h5h
9egXYgqAmrSOFKYbmkkR3utnECFAsEgot4/YL1X3OsC/vIabMsd0JL46AVPB6tDCAI32ztTaDWsq
4urfiL+eQYi1T7QFY+aPckPEhV8P/gTXPXEHH2vL7Z7SPlFFDCA2UVQ+tiFeezS16M9i2IsISxsB
mARl45I77kKXH8NycrANBdrdDNzvsJ02+ql2lGflwbCz2m70hy7svcJpaTvNqk5Aodt1qut+/zBr
wZE7HfPbGSZ+coffVcjjm4m44uEmbuhmE2PrsB+G6DEHK0C54KLmtFi4/3nOVaHbYyfeEF80Ooln
cXcHK8f36/IJ9NGqC/hvGfICnrZxY0kjq7TeKCPkBXL9+O8Izf5hutFM/cv+ck6C2dny4Z1SdEbp
6y0ndCDQBHNtngNEoD0JUmawAHeWOlaA7/sMiFx2nv7VWeQLW+y3xTHnIESD/jApvsY5H1VowACK
eZCpLXtSlKZKUham4Rz+P6sxvOUl1K4I7OjEwMBwlvH5QUzRGt8iUPShwEDNaHUUdEWqjuvAN8RH
9JqpfIKtOilX+Lw/On7lDDgpCic+r2Kg3197fmuZNMTDMQ+XqPour52tWOb5tW6CDZupvf0tFFEi
5JYJIXy7j0wGmon2MR/+gXPWCbVrvZHk7IrTXrR9HrzuIY82HU967mRux0NeHM6OOLyjDLMeoc+k
XZQF7mkKhMsLWA/XV6jajkGuVhrAQOy6HEmk4BnbTJcukZSy+dEIe2mb2WVN6l/YBU7hmefPr3/S
kct6nVEh1QSEwiAYW7GJDNsjtX8DalbClRtUfl0BHzMHBLOo7hXnpOFTNmuS54xYB96asPsvHCD0
kVqbWqROrtP6+2DjnjREJkm+8RDsX6TsYTHS1FJ31Bkgdxp0iPi9F67tIXrpQtCTdXuJomAPfhWo
uPdSgrN/FFhsH00Mbgp1JXdChEDW2JH+JH0fcX0BM/230YZY3Nt+4qL3wc/Emuph4tnRO1wqdXH4
WI2Hizpu21AFoGgkwMFwRO8uCskemymG1PwFgALCQLllp4UkMqrwxB6W7e2W2kjRQbUuEoW1vbWQ
9n9T/41wD5upe5xWmVo/jqXLk+9bvpXpe0VHtUza5pg9RIdveMDOdHEvnFCy64dexaD8yosAJ88x
mzJRvVgAshnMbDlGNbyvZJbSG6sqD5vnItlClFHTQjqJmgnFW/DBjqD+bMA5CKSbbBHw/S9rZZVg
8DHRmsQvzd3Qf05xxPmALFuNdeN7cfd3iS1/6vAijFTz0zcc/Aw88mmftDqZvZ7jAwhxRnvQD+/u
cGBhW7Qe5g9vcWC0+6ihqpbbdcrfm4aIretmEHEhNMN9CiCYFwwc/2fMXUP9gT6EedzGC3irrNz+
Tqq8nJxryFuzM5o+/ge8JlrA7VHwUWo2J6sFEjwZzutYx3OBRofVeosXkCf/SAAIVA/c2c5rckGy
4MS7BuNr9EIxLvV3YHAPoZfj7axMr2VEfH/p1WQJhb3Y8FVzn7E0kigz8McsptLul9yWEHUoY5dC
WLY0SVEMBDxMk0UXBkFMuhGGncVBAYDTWNlWgT4iaiAe43JjEf5xbzAQ6/lIRRjc+zeefBVs0e4v
BL3U8zK6J7YpTrVjZGBvGZPQwyPwYLpkHrT/GwfcFEx51sT9aOrCaaJeV5vP8qh7h3oBCwZK4mv4
69/CPXJwyFz6a8MeyS4VnLC2dkTF7qF4UCR+SnjYkVPSy3dkeqT9AkUHlwfrgOuJ4YTFlMiL2jOb
4oBHEpnmqiDLsJuujUWfxETf4HhXgtH/rrM/CkfLhBAUHNfLFtqpCBXBGwgjLIwhLnf9xyebPOfS
qup/IYMjy5bpD8OAMIIme/blRSMwbMw60OWITdYdjDVLhlSXFGWaKdi0QL04+QVK/k+nOWx8USty
TioiyKHUsA303Z3Il/RQ5k6lEmA7RNJV/iCC8rUMgGyAc1RMx22PejuqZa0URW7Mi93a55aDZuPv
qrdXgOtd2dYhBDqzJ2p6VfXNTikrbgIvnw7LWo5euv3FrPx0bKVxgwyQDs6TrfDjF+jGecvxoWsx
FtnTgmWzo9OqhR9h8fl12YdkpOU3/7f03/xDAeGk48gjCjCDlHF25ocavpRDYkJCNDZ6HL+HhqM7
dhv/YYGzZXgdSS6vtJ3T7TvcYWzd6MfHFIwkVsgbtth3VZ6ld3Ml0Ndtu4tgoSE3LHR8vGoox4Ke
vSLJjCKe1rJlqK53bxoSQBDtZ/Btp0Taf3G5n5DxfvSdQnOPXclArrjk2dYulUg/QokVoaeHi5QP
tpBGHvKkKu2ZguwKhyzIBD0pwpRTdD44xJ3xSKqtcENUYaKe7ewp3NuJJyTXhdS2Kx5LsgVesiHF
7XHIP5k1iDxS71gHPmEpKAT3Nbbxo4+L9LkPYA7sttrQJIeY+zSCSfxv6QEOwgoQtcOAEFBzmhhx
7v7Fd6n3NwJbh4p4ViEzmxhtcF1y3OMwr5pMJl+WrDKvrWPPouVisHTRkMnrhD9t1APu/SbQYSGm
sa4Lh8hqYqmLKSmSPkd70e8QajTeCfj40OIDHDKDPO0vLrspQpUgKbNZ/Btv/6osLHQ3p6zSpaQ1
nDRALCehVAgh4KroL9NLMannIPtYOrTayFd+Vx38ilnbqX27Fi1PSZin7nzGHTjCoO0Ntzrk8ukP
LjDC9HdadcQ4WC7w7KBpIyzDp/sJUIA7dMuZ2wECPflzqDw+a2EqhfwcB5ZJ6gyvn5ivhqXv9vJI
YogfAqK2iFT/Bbvf8nvrdQVwUM1/BZtpwYIuxvqLfgCRENBKNGZFETlBN+E45pqSgfFq9YB38ec0
dzdfKMenr36fY8PFeyEb/kMEegS+aDeRiTTn/Dj3+NR+hPgJvzplqo5jpyMWGSHoxDMEPHbtf2Hf
4xmElxseJRb/vzxQ9NCObySmntJDtSrCR91wNStINMexM4GyqoBTCfJZ1Tg3Asd5/mnLbo/UyOud
8iOcPNyTPa4awZ/vchgQkjOkGLxLVDleLHzWPZrejmhCeQZovpdiSgwKKhfLx0x2Vb8SsSduGQ0f
Qi1KAyYcKpy9AEy34YFJ4wBU/Bg+XtPP0aP5pPvPFGDi2ELCMB/n13mGjSj1ZXBIM9mGV4BJhyDU
cwTgiviuJLaNnT7/ADBedDS6lEBDMur7JDw1mMeUpZOe1QAqS2g8CQuD2QueVBzId32rAwRCita2
4D66epyLdv80VFXvcl1H1ZhGxGeWERAHz1FAPPdeNyTiGtwegv4/iFVrjsP4Bi78bfI+nV9+J3GY
dDn+Nf6QVpbClAWhno0YCKRSMsh4RmL5wheVDgTXu9sX6ty7+kz1A0KpsblvFWMVK4YSyL0YD6mE
2mZ3Xpcgr5/Ik87wWPIOP3uCyw3bayV6/j0hfwqFeBuCial+U6eqPtex/Fbcf61lLxSG5/WjZhhf
qnTLiVX6umdPgIDLfrWb0j8Y0UA5WHZcyRtQF97YAWtIddoExc6tJnlr3S4HfC0cK3oAAVVWfLqq
bK1OHAIyXlR64qvIHumDD/QSMTNHdiIhRgih1NO4uP1ieCd1JPOVxL/knCQDgzW5heporf9IWLHE
kHJosN/unNN/ttIAzAxvvtkXXMcL7whP+Hq4NJoujhxmMrGNtUCvUBs9sLir72OzIiORhW43XITV
thd9jZF8+BpqrVuPgs0eoMy5gTx51i4Y+jAq8Lct1XbYTbdtAZLR08ef3mL93kiBMvMZrxJ0hkx+
MreB1uRjNda/3gMJvbik1dt4efvXpGAgYi17NmMlcOGjB089X5721k86pYGBQzyHn+/oRCQ1OWPx
V0AKiiz/aSzODQe7boWK2oO6pgtIJUQcF1GKKxkv86rR7LNSzXUwNeLWsU8OGsccRdMibEeCOZe2
SAmXf7I68aFjQe7Zqy2xZCRlgdqtPQZa9VwAbc4NO1sOy9A6040GysomaiTA0FK7cQtzkQmJ5TEJ
egOxyPDJiu0/qXd1VqGQdFOZ5b/9LhN0zaGV2DTrgQM5cnVWspsHdu2AIglrpcju7p9linngerzG
ZgaxPV1qS+Ag1SngSh64oM1/LgybJpgzVqJN8eibMkw8L/VbrgaDIsGCb8ongUnoc5/sfy4YvEYO
dL21IbVy7heHwBfmIzo9ZNAq3/vGtIqSfVXYj2efLQzDIhjcr6F7olaGUtb5SDXwxokcQnGq2J7H
dWdTnu5RSZFCDhSTpCJUmAdMevUYLvLzTXJuAJRCWenL3nbwlZXHUabUP7P05jRog0Vyq2PwQiKa
fx8NApqAKIH008QrpBjxk2LG8X1OfN9l3hr05y+goN+O95OEh2Ttya65vZtvi5vvHyVwskR1TgNW
NEa+TJKRgcZcDOFKHQhEn71mDJYCThmQZ2vPT1NWOlCJ5uIbyswGiN3wtSMZRjrq7YW6wumnvJl4
54yuJpIQ1A/E5Pw67qYmFfb0jCtlE3J/W2/0jWBTKySO8uuc6jxm18HNSThWZnfFQrkbY9Meap41
R7kRV8TjOWJmxmNi8VGGhcHGcPdT1/16R1ZeFFW2hWe95g1SJZsWgfm4aaeXBui32Lfe2sViDBJe
RuFKhi04EPRe6x/OWnPVRO0PeVVNVxEcUHaSNJXF4BLtdYIkBOVwaJ4m5wiXGh+LhYWvS9F0u7gc
gnWS5TnkBjl+piHlJPYnY/ffMt4LnOXLYV0rCokE7dX4+8A4Rih6wyK8BKiwrr9kGkyW7njHgrlG
yc/SaW3YxJDem8Igc5oW/qjg9SVLcH2xdX9NBHxUiE1oVJBEGcZ7kcSYZ2ZRDgdyzUv5lbGNSwD7
N3StU/WGKN8DZo8AmydMpC8Uh09hZAqzq+5vazLxvAjh+lTXUMIFKQQPBUNthqSO0nC6pobecWbW
fLEUkn5cw4Ilra9EyXk2Ybln7jeDE1XjxYcOKcvpECcx/eyISitWBILgHdAa6H/U7BXqwpUs5WkJ
WzeZ73RKwV77G5lk6Un28dqkDPN3dhcRgMuxrJ8QTeZ0NnSVhRfjiO6ixHveeMyIcPr8OpyFlsY4
HVAiSjPtMKvz/E+chj9idX0qhJKTzNZLRYtFJV/2cdbjvqS5NMdEgV/OMnjgiLx+o7QELyA1h1wu
5t8M7VrMFCjnubw3W50LKeHF2Eqvd/bqk1katRkUBHTENqIi5maWvSRbutMnvFUFHDV/ENF8z71P
ZSINliIJlNMzTUd8tMnKkuQR64YyR/N3BGPDfK5pZc6b3fCUCGeZ1r7cSkYM3p64iQk/bZnvv3Rc
z8GtkJIInwxLx7ZkjumH+5B7yAUAP7c/xtGVsR1YhfU2TA5wP6Eph8W/JAwu70mddurWkmnq38mP
rOuv6oof6mr98KnKlKBDGUu7hsct7YTqnAXDeFzvu9DKSZ4rdTQENRpTqg5dNNKtdmGJyCAdTNkB
UA4t/qE125UkGO+C99deuFf3mUgHpcMVbaT4gqEA0uVfvHs3rg6OEDbQjWE2oh2tbbRaTh2Tl6P/
SorYUx/bukP2oTttA0tTxdxC57yrUCanh6XgetOCLYcaIOXJA1r6Khjs63fwGA6WwqY8D63dTM1T
WPQMvbFMxOjy3rqedOR+S0MSIhn7nbbnQTeGRLAvyIPvbiTw4lvZfBr8T0V4z5ITRd3qHDKA3JH4
BJ3C/9ZhrDUV9J98VkwrfGdRUqlboJVRQKhChLIxocwcY74vsXC0VBXeEZF6tjxvvZpsYv9uFcVD
yShZJ3fO87/8eyNM67+3hcsAl7gTdNJ9mZl+KsCE7Ow8f11hVjWPpUozi0MQzQkvniUy+JtHnNYx
18BtbiNUH3+YJTWIa6eOlXQjHcnZVGy1lNW1ePXxCMO8z8dLvIqw/Zy4EbwQianA476SerYlBGpG
5YSg1dGA23/6o7fS8nOUIZG1xQt5WbxfHdGIQoPJzNLEpB0JuiKfk+5T8TWAlRR7WYph+CduqkRr
6Yga4deIxMq5ki0iZ2MecKrM2BtYPytngesoeClBUoC8uKqOaDCEEmsiNARlGwUiP8a8Zf7adVSy
DBMd2zufjQQtJ4t/v7+wUm16DciQBbxsUv6bo6X54bzSqwNh2UKfvE7FuBZwmqrzpK7aG17dzsNs
qmAcC0hFkfIDv64+4eMjJRZmrnVRVoH/WzY/NNiKocxwR94KrNG74kP4JrRYtAw/7MmaP9oosYe2
nA1AlNoexDYal9dWxiIjJMIcpWZAVOdG+D1rXrEcTreLrli7Rp2Nau//SuVylTJ+I7vm0ezrli0q
/Lf0aEJULpGata1eywPa7enGOjDgSDDb15dRsvLMQuNqdUekMbkJA8dWU4QhQR+CUMQsMl30uKaM
ISOfufMG50XLui9FKRvfcIUTZIVOcg+aUC00c+7nRkFu1KK/FaS7J15pc1SjJHpZHma10zGjHZsT
uMR4pv2xIz85kJqCN4bhNJ/Pgca1eZfv85cr1UxFwhZyngCmO7wPPGJpXrlRlXewb4wrol8vw57z
iCIVljvBz6mwuw7Wf1viZas6trlQmzAK7/cKQzFOtvukJY7UpnS/rhq9Q+GVn5qdLuDrZTKPMs+a
S7CVlzh6HJHLfE1YMGK5cRP2Q8I1s/s9Qby9RHExmu9ZU16TkThY9N8wKPi7BV01NThLkVM3SFIX
B/khnJrL6sI99khEQrbBwU0Ks+NNLcypu7xQl+amSA2YSSbfm0WdavzwbeUrmSc+4YL3/6ou+xE2
JpjE2EuDOKCJ/4n3VwwTKlNFsQd+wPfN/gHN2Jp/x7X8P7jZRbBox/W2povwG+/YY/MxMR9dRkvg
1A4dUlN+h4KcTtYouNv4gBRHJArO4qzR+7gDMP9U9Mu8o91MeKRUqsj4P6ls4EAlD8dZCpZJ10Cf
eB5j4iHY/B4rXbSarkMt24aTvKNDxSi6bDtNLlCU+5kB6SOlDQG2ih2kHER8DSezErDmMmpsQIoS
QG1518rbml8wdMhVBEMjILxMJ5THAD41mcGEjPLr5KzFpnmxBN7Pp+9Ly+WacRkQnFDe7iTbXJy8
rT1xrdmHyNgi52nM6V3vlFlq7+oGvjP7OzGkIt6fZ8ABoLIIyb7Ve1as+wGbakfRfxjCqJQEuqE/
lWo0KWihvod1FEog/wRktpvU0G1toqqd/W0hybJ5MOAr/tN0nkEqarWX0/LaXmxYadxLupSWVHoO
l3Zy1BUa/eM61BT2ZmWRUP/GArw6maWEIa75arOb4+mTcl0SBK5DjP+eC11oBtKBayxfqoFzjyl6
mmQgTt5H293ZWQgQEgopkcNWiD1Ri1zMLRWWXLlBOhoTnXOmYYZVVhPhf5cMlFeVzVaRtj/OdG9f
dXtrl4J1yY6WSf+4viI5Ql94LrdzgC0R8C0nQccWNaYhRFoVB90tnBmKa2z+xzON5GVQ+kX/0Gqo
mofwUW8wEfuWEo1Fx5ekhSrR78Hr6Gz5rMoVnMaFOHREsQGDbkpezoB7WrUQFBrWDWWmwKw02Eve
pd4dbmkbr3hkCrb5qtnM52FZ+JoC0rSnpiMQRDtpIgzmN4MoIHNc1+n+Txol88XFPrSiZnlWi3Ie
lNvJA1YNCzVpJponOUvJZAG29C88Ugauhr1wMIJJCY5VD9JtnNSbas/OvQrAN9HjZLJa7ecR1zWC
9N9qZUhwvvKeT5oa8B/ZAGD+nuM8PSNGi9wVTwcnyhn/Np10ycgWEfQdFhtV0ErJNzeRt74FCkEQ
TWDQg5JtM0A8W+ckKqwuawxpw/8JQWX+LLWdthVi64ZqZXbW52Ocmakcpl625RNv+2NsBitoIGj4
/p426VWxv1smptQ4epW/uGrQeSTn6H2KGiSk5yJUtE9RzR8lpioUUT6GJ4IjFlEB8NirQO5Yk2Fn
wWguNCktVqY591GqTXEdOBFrDSF5NFT+JM2AyFlJV0Xdm4KRXul3TlkQKaDTuuzUkaARz3PoH/C6
vr+EnDog3E1KN45r0WfsbztRbgLLs+yGCtGF7Y/P855QwDDs+nFTXik9DdZN+pqz5jaoFBNyaTmV
fvYIY5NGYPG2O7UHFzbz3Uitvj5wu0xnpcXrJIVer7Zb6fwYBEKrS6csEO72k1OaSxdVkwLq1a/K
WFOwiEJhaNxDQnzX8mgv3/cEel7KmJhGp14zoAMkkrhAK4ubbA4btVLOwNVCseai7pCgyjmk8mbN
Vk+0ucDqEHIzUWAyz1at8AXRQjkFYtBAEKm1CDeza/lRG4wvPSDw6LL/Z7pOOYKGhJOVq62C4GsC
TIlCiOtLLOMbIfnDyEzpWuHDesmh9gZDjeRRVTHGTLkaJUlpDp1F9sxuPhSjF36ixUC3tAUbJPWD
0K1YeMQxUKhCmN6vrgLnnOhbtO/kQraQhUlhRU4v9uw8IN1EYUSc+FcpBZCk9q48TQoJv2pyD3gD
YkCMKFYltIa/ZixMp3msbRVh7+IgpWCU4MNuXQWTA82qZI5M6bH3cKvRSsqJFCw6lw7QqoVZ+SWW
T7iX5MrntqHnG3o5MRiQF/UiJM0zVl/UDcipbcRFae3y4Zc8x1+nncieVmndCTTpqNnYn/9I5OKP
MV/OB/P0EX+BpayQ7IsDP3V0enUjFaCWVa/UDfpMuOjamhiI8pV26/DAMahBMzhTf8vOSd5ydMiN
D1Mhvm54o4TtOzCkGxQWG2Vic53FQMlvY92CDZ4Phn8AW8mq0Llqy5kjO7nIdG6TaBe6otk8bJq3
LPyi/D7UJXB14VwFb3JVhvwGUUUckKd24aIOnokNmz8jcxIS8KEMCSjJyD+2GyS3Rocr567imM2X
ZxoV0D36lBZ5OEFkrorRc1k1NUYYrxJfyFXoaS9DJDY3cAsTrIzZwzUWoIxB3tK5tqc7qnUw8naj
kPzG5rWW9HnYHWAF5gLHH3Ru9vZTkh8t7gXi1PwMTCOW3JKgZoMA3PCAl6hxS8YpfvyrPZhYnmnZ
6XQp1VpJwLjjFRNyND1GoCKL+gGn00nv49N+Lc8pjoaaXrGeQuyjl9QZ3NeOBt8lj1TPsCgi94Sw
W3J2Sd5G2vtsA6ZZcxvC20PB8Yc/gM4cqydItMtYEQtUW74FIfSIbGN0RjomIk6TXELu1Qe8obpS
A8Q4gQ6AI+dGRcV3mus7V+aWxf2m0Tdg3NoF65UKJO4JBQlCGxbiuvVj/J0Ze8gFTXn9RLiMdabR
fyF9TDs17Cu2ks8wWMd4Bkzb/P2xi4ROYqyV5F0C7mOuee6H8xSJfYhpu3UwM6Un2bkvefwjZFKv
I186aTLSIL6QEGJcgXAeylH3h/9JIsJ8VIhdS5HHRk6X6iIeqCG5OeonPv/lzwIZbGWfm2kD6hpt
PQHGB6Fke0nGzh2mYQXgaQ+iATiAuxf9xkoK9sh/ikNjEPdGvReUyPt3pZj00+d9gu6kCqXPdvkm
4SWsieCuEvWZckVFlnsive11LchLW4/Sz5kLmFep8pDawhmOxXYjBxPktqGudFPtDbR6bD4Ld+wO
NYAzSqTLaFLU38Fxu46d3z2zunfkJFy2L7J55GH434eBBSlO9biMrRgPoV/z2b8z34/cCUYvkUW+
MrFZnFCIuDT/e43sK+hjCLCdmlcoCEpksRELMVQpjsX2FeW5Hp3BkCjMfthyka/SxvFGkPnw1YBz
GupFerHY0Xu/58G8lM0Ujr5AZRxOs359brN6qzBZkRoCvOI4siJLz/KyqzLIQeDMoTF8BEeShaKT
vAu+PuoktDEUTBQtJX0PsJPtfgGJrKqWzrtiYb2VVoUkBZx1hX17JBZRCo4pdhROWGZ3SxM6UxpO
TQwpF2v05P/tcwNI2KL7YVZlyEulKmjI2Y0WqfePFC12IYGHiLIfRLoS7ukmzO7RsV1n+zsG+rv5
jPZgRojzRcESo6Z75PhsNCsc0rEQ8BMrcQyD5rDuFZZZ9ihojFMhaxg8JzIoxg21ADiBizDa1tdJ
AIWwJDjqvqncCkw6e7ofJ+V+XGCzbpjomBzCMalEJIMsQ1IW9oNHpaun8FGhc5RlxBB/+TJQv0bp
sjuDVy7PAtMSiPQ0g9Roac1azRgs3snmupBOcp1uL/ZKSLaJeWRAGM0x+9/iS1y+iTjcxJgLCq85
mislnGlwRB337p9pJ3BjRYGA+d10+H75umfH8OAdi59xclHqlt2/oGO6ix2YKcpyL7sCX0raUxGr
PrF3Z3JORCzK++zFYt8nGwfFGU/LFUrpRfoF5BJVMfkOtZjyKioSLdG77W1haNjEC4m2L8CCX+vr
5UMw+ITIuOrsQDv1ngs3CzDCJWBxRtXHnT139P0d1/KzKU2UlmENUMbKrqxlV9LCFN0tdeDZjMkQ
NvlQfjNTTe5cMs/CdW68Er5Unf22G6EWN3fxq+14/iFsByJ9VWYdK/0Kj1b8GFKY7Qm3nbtjlY5m
o9nMjn02SUajViTw7YjUQys69ifrJWDaPfEEjv5d6jdaoJV8yBa5UjNmm9WmhjvayW8a8yQ4X0R+
WNNoU1hPpgOX/wJtj3/RbRJF/JyaBmirSfXQznJd6FdiCkFtA323gnN+ThMtjvbb4lGnMMLtUyeQ
CQoBPXFHJKGn+EKop15PhM2KXbLvEB4Uix68aA3eFAqd+h98krTx0sc7o3I9B3583ztTrpxG3t1b
Oz3zm5bE47EaXihp10rKfnDoowiMIfec6DDMNxIGz8XsBZFuEeo2Zz560wY9knvKgs7yeSaMZkpz
+dp7HS9D68B+hAXS0rM0d1ND0OJmavZ1IKRIUAaMwlGdeJKpxV9Fb0OnGG3UkxKXQkqG5CwfLpnG
+efj3/RvNq0Zk2MPnRGjYuLRcfOEruocuhQUlIoQRpAim6cZ3xY2Ckj8gI0cHsaLE0tcvuYDTGi0
GpZBi4y9gV/M18ePSqkiJNxEYCtqNZaSASUY0H6WIFCd6o1JgIqS2acgIYhWsTX3grrlYxA6XNQN
9ymj4T8O/Thzz5i3v9bK5gjIhEz8ZsgJ1f+aLU47fBq/wJ1ljB6KjtcieVzq8b5LiUe5AauDQ1mi
TenuNL7tu4Wb1FzQeM5SPVkXPWe80CJ9ufZkGIf1YDMV7LqXiXt+Kad/CNvCO1YqHckSHoTi5zg4
7tlMro6TZT+5+fJR6fI7/t0I2EjZ2UkVKt5GIDFbiu1PCdVUIYoLaNz8qhGDQj+wMWQG/c/SeOi2
1WHLtWgQ+XXBIAQim+AeGT8lPpDhYSizyEDxtdfnvAAEUX88yTzYP+pAC+xrnNcWb/50VRW6/Gsl
aWSJ2TcokDz1Vcvk0MM70MZPJ55BA4wpfuzFatVUmcpRvkv1lgk3Q/FQrEGHLXDhSNz+7fCYmSo+
snoTLB0N+mYw2mnEGSoBEgGqmGemJXd/xVfudKc+UrsrzKJi0D89Et6Z62L1RTThojJJhj7TzQPM
9rka5joJy6gNO2sKtQy89zZ90W9oARM8m316BI2w4FloKcwAtfPThp3mLMSogF0tr0Et5e8IHj+8
H36nfRXO3Z5iwO810xHIPcbd3yOTq3FHbav3eIz42nn6Fy95ak3HKVTCHh+wAE0wciCVY5o5bAYR
+ozvUUS/Ls2aKkFJau5iuR1AbsK28MyvLiDl2JUk9gXDNwHURzm+SZRsIq9u34RM2Tt70GpuJSIU
7KJoT891E8JPr7YjdLqjF6djwZhYyEVE+O4W4PU1V79TtsC/sC9UYEWWBYsXjGSzS5xed7fzPCLj
Qoz/e/ABN2+ZRtz5zMdNxUVoQP6j6P03eYu7Z/bOy+BLxqgyrGKMjouJl67C5EUms3HXVeTE74Mh
rCA3TCiYplP1IW8ht21Pr50FftV/M3e2FAM/JZlksWOaiM3NhccJf3VGMqEnVj8xLCG07fMH3s1J
VFIKiu5fNig+XScta4x4GwvhWzrB//0J1DzVSUdg0tLRzq3C0WjfXCWaevI5afqNTt0/8vo1m6yh
wnMCmCYT/RbFNeveRZ5H44lxQdvKibEBBns2GGJEv33Pp04yUYJlY7n8w6VOQR+5F8EqH3jW9IbA
Z7P/8nRPcsEIQMwc2Y3x/6DN6C75R9L39j5cwpvSV/64y/n79+oA0bT3i3S8xOpSDHGnkwOzr5SA
E3JbFFJDufpsHT22u6WVQQw3gelqLFagnYyAkeQEiF+lbJFXbfyzmj4wUkVUtAqP9MgAxO2Tfkmn
LdhWrcnPvY62oh5mGc3/8eOGImoVczS5Ci7EFkvfOGiim5W7nNp1rGzMLGgPGPuCGPYV2Mr69SPC
WlPxwxDdPvmy3uEbESHaa/FkAslaZIEG4w/UlXsXm63f7XsSUsoTY2Oof59+TtA2i272++tPLbV9
iEdDkpVcz+0FHPn4DgNkcp2wDULSwwqk+4ZQ1htNeOeOxSQY44hKkOk/MyQLqFCn39/uAvylya9B
laxr58spD/vd9x7wshqqgAUglLxfW61Lwfn9C0YVhLMxc16LRfQ4AjWY7vrYDm+OfHRCz3TXvxrO
InVFpBq7QP50Vl3inxOrBMqdJUAK78/ZMgAj+TJh4YmHZdFtOGtDwI24h47kF5bZDhDJyTFz3Elu
aU1/ArZSzvDiZRd/s8In3g/COEzPk3emUE9/1FrXP1wJIiexX62VltnC6YepQGzKZ68v0BB4CoMz
andSp9DekyW4aZVv5Yy+Vqnq9zSt5Fi/B/C3G8sFDYouqFCjYU03/5XA+CKSl9VQEpzjtoePzTtO
+nF03jFlzpeV9/p5sLejqOGMFALxpC7wysBaef47yqX1efA9ONUnvBzKp01vPFBX/EcFVKIN+uhp
QXuGzudHlggFtffLyARb+v31ron+a/i4nJ3vDWcriFK09Dmz3S+LHCFaxkLFnM5GgH9Zncf8ullC
xnobOd8mVj6LHW4iBOml78JTWV4LigSClDKBwj9ML3BK9g4acA59POTr8SvzGyOSu31DZ7zU5O9R
bdlHW9QC6mpqNvOEZK2wpPgnHSljV7gYGsPcZ6bqVBWxdGDpE0Hm6f1R/IG+y64+Fx1Ar5O/F8mC
FPsRqOcNfTTypwtCqStW8D0KwS1z9q9PxgikBAQuBobJ3ElzUJ1IFDtChj1t7YlpLyygPcx5i8up
JoFREcsVa0gdarC7wOPqVNIo1J+twlSt/gpH0IMPDQV3UpI63Kkk73KMVD7oK4199dfgyS3veEzJ
KSvFN8IRKW+oGG+wwA/IqVnmB3/9D3wjVPpRO1HbR/H0/mh8pRn8lAhBJhaSqrte/i+mYW5lIxGI
mYxenm3TtixNTw3PGo2xm1P+ioHalmiAkBixNTkmCn0Rrcb84uwZaCEp34QessdEwK3oK8TwbDJi
u0oFk09pCOFqfAcy5yeSNXBQD+mWDnUbvmbbRRpwqyGYT0C1KMSa5q7JHfHG/13nxyGJakx8Fqq7
wWlQ4brQAobo1QRgBsWlYKXMrHvr+daeoQZDXjHkeDAjy7w93pgh5Vncs630qcLWCYcG8KtMgJxZ
HU19Y9tgE4Usy/Z2idJt1M9UtZrlzL5P4LCmY+ls12z0Vojii6DOWXJQ5ZVVMQmax3+yn4Cbx2G/
YdwVlApJfY0gyAF59ENTxoDhDpIARVNg2kZ2l4jWiYnG0d6s333slMNJtxYCycvYyOEz5dVORtWY
8mjBKLmRldXBEKGrQ5Xs08G9D30jjfpE7u5bLUUYLsjjKppq/9GSqHZ5XnFbakuC5AVGG+szS/5y
4HHpulSqjX2kL65XXo+nY/K3r6iBjV0rTYp30VUYjVbko0WImo6PiN1nRKiAyzfJQTHrWt7xMSDZ
Ph8cIXpGUV5UbQtjc8r9bH8CLKY7t8X5PexvkXDHAIWJA7WPHsQvahyhw6eGT68fzRLDfuO+DzUO
2vNe9YfTbxz2a9jehMJ5cxt+vUnYYAvMm8USwTFNbAJ+6PctCaABUaQXq2ujW8fFTcqkQ5v/OelV
mQkoFuZsSkYzNB6mTwSNIWsaU4A5uxi/Oiqjwnh+F0PQC330stutkN/VxBjf6zQMaY2/Jf8CIWmU
gI/zuTLlxl7cWuoWr6MHRfqF+sbM3qH95MjbXYKIhWxj3f/k3Zvsz5ydykHPI8mtP3j/kNuZtfkG
a7hyBxY34BPyiABewl0/SiaFaZiy905JFS0TmFZze0NmhBJdw+bU0cj1bAGE8HtrDLnVnXo/Alg2
+dNMVwJvJA1WO3BEbiKFd4DRchma8qXzyX57uL2C10TIU4y67v4dW94kFKJDKliDa8+Fx5LvN0h9
fX+SEhakKacjd27kWq88iJd4DiUH+Pfz31R8NiQvV90dtHROCULJbx/0pBhA/hw9hHGZEoaRnyVo
v3w9Rky1PC/sPgoYGFFEUnEOmEnRnM/jC5GEoEmQZdqmTRvuN4lzGDgmo1V4mNG9MnNOOWnrRWGm
sHV/WS/xiVYPHbfuzm6D9UfMe1yj2FHeNXKvPFbLQX0wwAjA1VTsXsvDG7CDRrNQfm4+E1ZmtD3i
CROgVdWKqQX7MRFJTrc9JdBaxenwcV+TS3iQ10SrpWpmL7n8XO2Vm1IfsAK+deIdKg1gbA5GfAlv
PUrLngp5+z11WAu/ArfJX37H7WS5YyzMHmSuPnuvRqLxoV2otrSf8umO0Lygh7X6YHS5Xs8b5cah
9GRLzCIQNLQsvA9b8AwoXEpgPsJMKCX3Ds66k6bmmxD4uipNLwluj24QMUDOxxAWNU9sq1ZaI3ig
kZYxTCTH6qS1GCwaY4vWx9BB7RYvGMhptJcoGIRoYUeV1OacOv/e/DsYnRHnuUZLRAn5bZjRoE2q
EISLt6mclq0GB26vrCmkHz+MdbZ4SErSWPGqRlwaaruSlHQ50OrSru0kphBFgmjfMKzPlxTXlliX
0wqGTQPQmMGE9+Oi5f0Zfy/N6abjcfhEegxFR2qzGG+6We3p68FO3eB4dHvLiPnC00Y7qBBL5g+R
H/39ZvSa4J03ObfS8T5KBUmF9QFnsKeEeXhNIpECYcBszQMbSGKlSkXjCqRQEmFUeCXBMNJjMyg2
UtLs03z/3j7XfyDs5XqzO1j0RwNhonIW5sXHfPQHLmr2RhK5b/q+4c5pxMFneyv8/5ZTpkuP/zIX
EbyyssmdtATPv1he899MONC/EPVlHMuz1z30l/hM//GU5IfrQB68V06WJWByrNlXqndDMDrOqwJW
Bj844Yt/FOne/LjzVYlPVNT+G6IJP5AdvVx1hXT7T5kqc/ehZVKXTD4GNwQEOWgXYDp8rP3OKb6Y
JhlPy6qUBuLTA3QB0sxGmmuhiB4sugp0xRNZmcABJQf/cL9hCdj3g+J90fyrsYHR8+mjxFFsuou9
akOl5RX0soty1ki31PRtMeEDQdTPDVs3FPsR7BMP+NzydhzuIfHRup33UmsETJbB7HBtmlCDVRpM
bGk8UQFTwQsIVX0UXkLWDeXBjpj1MHSgH1AoQaAPadZ8Kwgm1ayQxPFcm+disjWdjnpCt37txMIV
jCO+pF/a3ePCYB3bsrQEyS0LukoLbs8Rwe54eb+SB5oufGwxlL1sSrYGvPfBKecyuivqtUETkUY1
RNXI9HIFPn4yrNXj0tlgYf5ahnx3+By5NhEtZhLk0FryQAe2UqLJOD3WoIMhaRsvAMm9oz2FNK7j
ekDs033Lk28vixQuQe+tUzurU7b9ayyAX7+imW5d/7hsX9Tf+RaJQXeatV4FUhrrGAxa4QLqvUbQ
qcjstbVOdM40bQS8FzdyWzIGXxUvCGJrDsk45cXRHucSk7gnlIPkhhLxTIqkGC0BUcDPVFX8/Pvk
dUo9bAZ1c8/7Feeo3Hfjh0BymrWotPBmJq36yGjdOv1MRlbx/U9XWgHg9pCH2jiep51goGnuhZwx
ITnCa1yU5zUEthfHcfYYkIozI8tNqgd27ql6fxArJk1ALWTjQvMgJCnqugmOfRAWVzVW1cP/djoj
zAVQpoF/H6hAGC8ypHRYu2KwygBURV5rWDfean0Drfoa0qDf+nncXeq2oky8fs0F65nxdNGdZkGV
Ryze7SDEikyI4aUkgU/x8FnYuZc/G7CN1msPk+y0z090LCfsz/4gkmoSOKkJLzYBf/WeTsS7O1O5
t7OPR7QltJDGipHY+PFRczGsq6GpE6erbSv21z8kaqZakbkVlukgoiSlBwJmvnlXP05kb9ZeC2Ek
Ui/VUbIOIXMdHP1szshaCHiOEy4DDqYTpk30LjPSq2RbMpwhtCOJZ+lMuqmhI5liE95GbRAhJZn+
tGCJ/Whn7OqrQ368hpKwdJ+oa50CjfoebAPvhmpDoNPxhXh08ubbhkxmKLedBL0vpmfUjPub9J/o
NjVN1tkkdXmPX9sTQu/Xv0pAaSDvY3tdEftm3JQFAA3u4CdvhSrYLIpepxyQu1PHZ1PAtb7RKP9j
kgPYtduFhv9nzEFUexmoR2nabOqW8W3gNrL+WcsmcGe/lf5296rQYIjUMXb73L6/XYV9cqKtumES
HnksR053Z6CD4Cf2wVBqNtX7CDhcTHyENL4wr7EAJMlTvwoUzYe6WZEvuzZ8dCYU09v88AyNwZHW
biPQw87bnUOr+yiJZ4gnmx1E5vDqg+PBqh992WoTvudgXA19cVSmNbGRZzZhd02I/NFBhMobxGhW
3Qcn3HXHwgkMuWiYZcdq8Ecgfpax535ohJf1NjkeThkX7W8P768rp6xDjA9R4pk+cs+/+dP+//Kt
2uDBKvnnMbGwYQSbPQahJ3OC+57xiWoYbWGoScxRTKs5A0M7c8W5lAD/0xDldMz4TVx0KYJhVORU
4yVdg/u9z8oyoInxY4OF9vdavEmvuAh95yKuwqBnrAm3xqZGxF1ukqhb3YL+rMFsZKaBmQe1254n
GzqP05L17Fk4SwNXpkrZ1ldbZaDYHMyQvkBcgJIzcacmgcpKQu1bhkT9NqSmJlg/rHieFC0bFmnT
fZnOH3Pl/6maIKJEU5OxM/ee5P50B+jQsCanxrQsk1wITnReHmO8rXpFuQd4msTV6Gy2QEG9nKJo
OA/HysEwqVunCXReH6XLUevSb0pXtCWacUj03uLa+Vn/8AHwZ1cOdStm4ZA12e6m54H+NDn9wGyg
1PLRCSS7XiUTn3Rrrpj95STqrZH6IOJug8C5y1Y+y9w22b/Ppek3/AZpLiW9bW9QBtqFjs9z6amf
S5Nf28rlZ14FD5l3tomEgeFrmoq5R+aaiFH+4N9lCMPkZE2PncwSQoJWAVKar0j7TAODOHMSF7yC
LHVEvABLf08g9twK0NiGK6rf2cCJdOLZuXgHxhHEYVNWDxilkq832AXgabUuv3Hw7jjTmygLtIvC
qgrjuOnw4zJhMU+jEvYG0A9aNNbhFKmjuj/GExWzqJi4BRDLMLHlAj/QKN6pcN3x+pYGpQXlNQmy
nKBxdnBD/W8Hht4Nxly5nQJ6lG1abvfU6v6MDks6P7xM7LDEQArEWttPpXhozJvNDw7p3FcJRdaH
uqe/z1d7w8vh4XiCCyigiPvdCKmbdksKh1Kc0X2QXBvuQKrkDAXQsuKjIvT9SdDu//Y1H2D7h6ve
mkW3yk3/8+lHayRvX/rxI4LqxFRYku3+cWt6GZSQjR6K7bFTgNqXnSsjzCa0A44z53gSeOu1xBed
zmhP83RYC9WPOYG2b0c30+IRb12d86HL937XkObunUZw6OQpQEP6vaa59tugDEXG3IqwNM2mqAAS
IKtPTfnmdvOj/k+kHvTaJU7Z9WMDaQ9DP8cNt0dwEA/zdeTqDC8whx1EE5VKLNCjysSxXJ1wJMnx
knsWiXDejP6Znl9biH194I5r05bAriBRwkHMi5rb/ccb3oxYJNpCv3R5rlAV3mFYXn2n6hif7esr
6L3CjqOCMBlzu90HZAV6rx5MIVKMN3Y99eveRgEnDPur2dDQt+ftyRmlDf3/vKMghlEuxi0DPOqc
xsZK13saR1ZP8HLTSVYOF3RmSi3kl/nreAmten7chS6DqfOzMi85wO03JPUD9TSYSMeL+aZ+bAI4
uU9uTW2jClMAWVW+chTWGXNBaVLCKiBAsHil63Xjl83es+0SzrOLk9lBHIObTce6Y5t5D7XyIN8V
P+7fWP4P3MqQlmaSSOUZ/kz5oFApy1acQQ7/NbUFH2Mjw9lBFLf2Lvj3gGqa0s124iSlMEJSkHwy
uO9HObqVK073Qz4I+mQnavEy/R//hiinl3d2V3loAvURpVPuq93y5hv/osatLFr1OEhsb/07isuN
3D50aoVJpUqKTJ/tdg2ff0Obuwzk91mgm+7n+TOwl/sfxescsCqLbteqR4YH12gvkWFEOA2fo49C
Ky9SvXq8O3J7A7YMr9XgnMaFmPYlYWVIuCrSoOGYNIz8bf1inj5EHw9Fyz3GI58OOYbO6PlWoON/
542sM8A5CJBDPQg7aXKNdhWrEK99kcp8LJC08MfiMcEouu43NXrdru5LTIB1WB1Fi7/ojfAG2jke
mroqCCkJxW5ojzyxnrixTotJKApMXLvAFDL82G7uk2SUV+t1DQsIflJKOP9CHXVZ0gLsSsvecfhr
jVlDHIl49jrzODQgCx1wUZ2gJMpQdwaDfnINb9zv6CfMWyGwuv1MPAZTLqMAvdgp65Z+3+eCVIqU
61Zl2j9AZBkTYqRrz9QwbAXirLF8TO7vCSW06HZPu3KNb9biLCxKPZJi5RQDRlrWoyLCl7PR3c2h
6oHRTi5AzWkxTNdBz9w+D1Jjb8artkZc5yclU4yEXODTvPy2capZ0GkkC/PGo25HjHPdAwGGEbv2
gPd5jk+8JZHs5ybI7lJbusmZzrL/4UhLdoT3eP4JMzW/+pE4jNjS2IYD07OS3qrS30ggUoQeHkhN
PhAmLgYfIOsD9IbB7+hpxHlwF/LUUs9u7rvxBLTR77lanubmDDCC9uws7B2T+jZiEW5TrEtE36JC
8l9JY/FJ//sc+ZLgEFlTIhsCVsjls5Rw/7RoVF0wXp+T9iye48Y4DseoQrMaaDk+9lphuXCteqfW
JLFMjAxQC3Gm0jRK7K1n76n2dYKp18PPM7On87iVhx9KGRPgphrxabeKhDBQNlVIqSV8AahLETIh
1voR6eIVYrCGIiPGKx5z4L4VisxoyhrGIGRy5zy5dumkbSslpbz46xXYIrTnBoIW25Jky3iJOCui
HDP0N7mvSHUJHHVgZd2uBsrxBiUP+69YsptNTPNJ8jD7a3prNV5KyBz6qJxAQgwFgciVl9YPQNeE
EjOmyLgnwZ9vW4isccgVOX1msb2pd2RYVR2Da2D0aPjpFkhYCz5BsOe0XXDDJiXlPnTM7qloWFzV
LpqQgtFq83nwPnJTs6gxJictw/0mhsPXbX3UjXcjLuazEQWK82npM3yXHNWR0fm5Mc4Kkw/IEYTy
qyj4b2UKOISHVx+XIzlwho3DJ0qXl0oB5i6x+5cPijo4PdG06HU3llD9AooZmTyi9di4aEqjxWJN
oTGWn4te1FYj1T8M4kRR+PL3np/GaxskvtQ7cXxhv41dAVPqVLHmmXyyh14Pdt5gdqtx0G0Nei4A
EP8RNt1jPT4psp2FSXC/14EgQnSkWs/cXfsB9aCSdFWLNZfXQVSX/7oFcHM+AKyvV1HOmo5XNRwx
4HHpZabIbv3OKwAJslryV3AUud2PuO222o06v+c6vfCjarTPyxfK1ZL70khygYNttD6wmcvih+mS
nTmit1jJ3bv/v77f8itIApyvkTlci2udnnLACW2hY9hav1a7F+xLzDx3t/95kRGxs4Cta/ZO6u6b
iMEkJPXVDZMW6caryvTphM/2BTTXGMyaIxemyzERqaizCE9biMjD0mRfCYQ2piwM+9vTAm5qGbCc
C/cwI7IQqK27UWFlS4ofMugHvd5noWAPt7Z6gF0QTXbsJBLqiFrTaiY/7Jomew4O7qUxYsZuO31+
07YIBAwyanQJrWnF7biT5CQOHurB9rWcG/ojsI7aqXVwonCJOlMZF8wlF2Cjs/gFsIlrw0XDefJx
mIuZ+sTkPFKtLqrEcbdL+iy0/TO/OYcQBoiEDG5WpUpAzaXQkjIPSZor10ODrasW4YYExR7UIQp2
f0gyejvd5bgpt27swGmeiiG/BTtRQoW28vTEDi0JksJXgo6PKHzZcUnNJ0grWF/7+MfRJ+niUlxB
ql8i6fjh/B9cIwXDMR2F2ObpWUOr8PN8L5AzJyele6DV/r9BLRrpfpzG4NRIpmcittzGj83ahOgF
8f0p59s/0k6oLcKf5DZ0cbMNJOPC4tNZjx/dSApsy+VonzDw/wy4zlNLK+oHuKJq+14R655Zi2C0
Hc5sqP4D02uBnUfFkhRhrGM5OW6gDkkOVPaU5W2By8rlHFqpvDGGYY+WPcRykfqvGcvXVypzGNLK
B3UhnE7d974dNuwZwa92Zw6saMYV1lkA3PeRym7jRLYXVlRqVONWKRl0u6LTUE8tYdd9Vefi4Rdf
0PAZFnpc8kw8dPQgxpu3aTU7srRi+eQ7tyoRgM9vqIRsm6MMgBJd3mMJs4z4fOLYjwsurdlUPXDd
2jwVIBADo50kEVG9NvkCr2CkiQCjGnKhtFK9c2AbFSoSONNXO0bJ5hxxqIg1ZpWTw7W/k+JoJYzq
M70wejetxCap44fv+UVNYiTJGJwFjTTmTWTtpJ2ihUhGVm37Ldrj56fa8UmP7KnXYpMmlf3HSS/B
uNSnRUYgB9/nvI55wmecGmaMCbHqamoCUgT1zjUT18k9+FsThpxcM2DL7pP5vxGmAnoPvmzakv99
7Y4LzmdKcWtz8uTtzmEZMsA0lRENdH94H+zl55WhIMkaxCPZg3uxzjB+bra+H8iJ2zkCsJI0Kwkn
MUpiwoZmlAR+ORKIu22023g6MZ4oqM2/O1MTv7Sb9CNq9MFIRf5b+ECIB5sDCBybTY1oi/26bv5y
NGTiBetW3KjC5T9MyZwehcrmSA39y/gctoTLsM3WQoZ7NPTr5X2LDAe3OB72sPBqUs0Af8jJKZ/i
wEC2G9OEIW38Go1dqw5W0T2IphBHxLSOtdC0gZ6jWrltdvaUlOGgy+ChB02aFI8x1eVBLLy5fKlh
awNjB1Aue4ROHjSqutu7NmQ1Bnxjw32vh4nYyYdHSh8hQu9awf0vNfKMAKLGPpQqsuB5MQlqntK7
D4z9vW5PAl1Y3lDdiVOjU0Zta7YeWjLtx28AWfBsnyjI83Tm20nXBgwTDyPdb+5YBcjFEB6ZHhtB
nNNpO73TK92ZSEpJu3P/mCkry/4jLwFYuT4dBauZ3KGwxFHiALHToH0xvAmW93fgCvz+vNXB7/EZ
2TUO7lw9syKMhZCBJtXDr1tLoJRZsc4OmiH22apv5DV9h10NXDxeI/9g+JysmWtreEPXfaik+qfL
db07IAiRm5QuHoyHZehumqCxOxIEmOVvxS8BdyIkp6al8ZSQMifFFkRvtIQWQvwpRJDCivsU4r4E
kXCvlznFik/vtvlCs1CLmTY53qEuvjNQ6TfvIcC+Y6SwahdvdrubqAEv2sUmS2csNp2GMUYzexFk
JOFv31DlNgHBE3R9+hcypHRmOH35kAMPf1/IARwG7gZSZSvfMh+UHSDDLuSGLcBYtpNh6wM4mNok
CvQFM8WE4EYY3Q7la5EoJ/pD6/RDrb7w6NbcS+cD11DBoaAJmRZaBfoiNerX3NKA9gLKujGTrR7A
INkshS52y6n1HEHCL+FIz1xWKVEHz3j7CGjpXhUWnSqoVSXa3xWdyTBB4i9jltBXUn6eXImA99KI
QVtwbgCpIYTFDTN2ckyT2oAWHYVyHkHP4m3u1W3BqfPUXxJjDhkXTe6cgVUNrwRKSSAhjyJ9yN9g
pKjD9nbV0J4g9AAGW/uAwZALgWwq/eNoYV3/+3Yz+RktFPPQVMNY0rKrTNtrhC+T4HH/gzzQ9QzY
OA1NIJU4+CJgt1DmH9oTeoqBytvSwux8OLwbF7WmyrIjgb0TfzZu01nLc82ASFo29TFLF0Kf8/Q6
RBckzuvTdIGd7fKkBxW5oTVJ9/WZCN6V5cN4Qmsarn/20gAw3995HSMzy+aBTV/jXUH4ZQhIwmLK
YrJ2VzbX9dafyGZO67B+9wcSv/8Lh7Wg//IkgwwauA7OTe2ETcSW6Y+qJSQromBTwMUmoiXVdTNl
vL1P38Xiw1Bm3MymI6SmIPNPPKCVQYT9AYns6wm/08Z6o+/sBVeNOHzaBfde6PfsAykbqTpZEOtr
cug55rKsMYbfEP+MN1qjD47XK01/BeevKHGz+fu94P1Ei34J/slSeeO/5mtBIJNGIfjdHEuMx60T
hZhMfWyyKlf6SyVBjoOQIwL0Uvk1tZVcsBwNISzR13s2gvIjGB48O+61VgAkDF8vxfd+1LLM3zyN
7i36ZEuWT5JNbEWcdzuNLJq+gYv7XgwzOTWP9TiSImUsdnDuVzlr+kVEXh2MiiJZyyAJBOzHNbhu
xZ+iLt5iHp0ErP+Y08BYkYBJnPI6xEFPy4EnJuZcY5+rWruc6sL7hv8nEhxMuD8hu12fEZI+m+Ou
aetuYrRjeLXygYe0mMSr0QlbjpvEu1cHA0DnP1RpT5YJ/AncU0WcibVM1eHrGyNS/SgnYyIGdoHN
4oB136Lnc8EgxuRcQAMwmnjBC71nFICYlxZS3dDCOPy/fwsEHBrvoxE9nC8hNKga0hQhq2EahS9L
DPLKTw5ykSbuVkkTGi1zdbi1yIQe6AmBorSQt+TMGTvgJPoKOpAkRNiyHoLwYhi9qKCCDcTIcJPm
5RyrwXho3aCUWwfejpvQSy7DUcc7oJ3dk/w41T4v5FOOsm/HkBpQ1FgapBONZbQdz8Cp8tKchec1
uo9i8Ztkrfp5cIjvjTAijUnyvzkrtDTgjvP+mR85UHYQxsZmtlrOyN5dauycBVLFCGlgUr0KIS91
UWo2gvh9fZGEKQlm4f+FPAdrFLXabgb8iMPMApmIjySz/oRzQ0k9Zr+1OEPnjrE3zmdy53xharcK
aoaVukGSX5BVqEMSaHiCiPSHOguotMh/j7uCcfw7W8h4TDCMllyl633WuDgnQF8Lg03Q08AE73q2
e9gXljMyymWmgzuvDsCiB0/6L06cN6JzZjnSf3VT2YnpMFLFR1hY0LddZnd8UT9UXBr+LV24gAe5
HRsEQFsZ7RPmocYic6d1B//3Aq2Inj10NOdsAly9QmoQAR+ZImaXaBdozx+Ongicw6uVyAhtSc6o
7UVn6Sd2DjCqHYVNtCrrpRgvjJXM1mlS7/zFUPY7XwfMXIFlGkKj/gfbR0NWO1FQlNl10cwzAhp+
oucVxwqVOO/or75YIN3bRPd6JgkjaSLrlMzRMRAf1QWWsfL94cKFP3CaiYDkEO6c6BdogKU6x6uD
IysOsf2RUdzItTLETNhAcQQIRvwwc7PQgxn2fAk6/KHAeJ6bJSebM1D5htJfaIsJ0fyIef7n+yyp
nVcGHFnApRfET9PhjQeN25oAVyZDXqbmkqY1E1MYizdnqzd0cbXI7tsy0mPjPDod5yL8J47FgVhU
fJ62gPX+hYAGYTfgVJi1CTVE38nMLANk3+ZSf4XxMk8tUGmhj2YQOKwCKyy8/ZsSuIF/4LgdqqN6
FOjkb4lh1ILXBNvk2MC4sfW3erYLAEtgsjDIhA3e5LzSQdUDZOdOKZAHxheJFRRZw42ey9IIxDt/
IWpPnzyIAk8dikKrl1SITp09vGrWl46DQnVdtkykBNgquqi23WAPb+DuJ2bxBPMIwVCdhqca+ujs
VgKzAO/iI05QO5JfjoBDOA+mZiz81mjo3fhTlnawOLPmNzDK2WCNkPkCPBcjARUyxoj/kt4LFA6e
MZtd4xDKiLDaAF8q8RX3eWJH12g19wHZEk9+5GeO4yuo1HEgjkemJv8jMGuFCWT6kL6AFJS+UXx6
cOF4N0Y70nQLQEB3NgSotZEWlvabTSJpMNeH+1+D3m4dMz7Hzp2E4YH18ARupXrUYqip/IHUwPsY
5flm3bEgVHY2qlk7JelzFGayyIE6bPSAselvL7zcdL5t5CsF7txGVE/Ze3Yhw/BXFN4ihwAGdZG/
xDoOIyz1o0MXZAYxPVg32R4hYA/aftNGeZTPEMEwau5Un6w07cZeWFs24zZDV4QMHIcKlqAzRFVK
eHzk5wUODTSwDxfOXL4i7iptKtkxQPhmz7jU1gP4RK0amqRbThB0t7OAqHjXE3kEZ/miVd7SHDAs
UiFrv2pjCeQLXbQiqcDhSY40tTjXbnWSYFgvsDRQ++wR9IIvLyzWSlH/j/xPKOUyt1G1e/At43F9
x+TeS1Tk19q8M8U/cw+ajywytMH4bCa9jqBy5WYCyovNoTKCM0QY9DvqnTuWq2XmZIoXwQ3945fZ
KkPHwzGbn2Om1/ipSoAA6S5NTHut2BzpPi35Uqkz4gPSnEZyBvSV+5LeKwDB4lChaIZWwQ0jvdZ0
fWJHtH52goxzfX2MPjM2LlGUSTLDYTZaifqhW4yT3FLI0SByUCKCsx9MMzkUWnaSN3xcM7V1u3Nb
YkY5CxZmZx7Tm4ZEF/onGNxzDbjS05j+OZ0awa1xtV+Nkzo+D28vAJKz1hg+TKR6WNqTxy1ElY2l
K/H2qmHYY3c3ltnf9gqV85TA/aX4jLdYfWG6Yi9hFsjfQ5v7LimSpJzYN8QfWNGeoi/JD3wIa3/Q
nHgwbI60Cr7sMfFqr4cBj0BaB3/T7mELbcAsUa5TC+i1gr2WVbFh9DMcPdP7yCXaU1kD0GELWxPg
jpZ8M3vbj3nXqZ5P9otoxaLRgBp86CituV9NksZIzKEhq+fyvb1CxBRdwmvFLT9aGmIz+c8UAqtH
ZAN2mMG1V4DhVibwjrW24gSwTxIRdt/Nzwh6bh3BS6A06TGdNpSt09b5qvgDhCDGN/dYmJfUOTFu
Znz7Vziw7vtQCqHe8xUewDFL9Tlbxr1rqtLrgWcNDRI/5txIBKvwjbhm3tsEaCGlntChqRm9U8wg
nRT6svpkQMIsHoosnRIeoB6Wq6e+CvUujgz8whY1Jn7mmLyyjlq8xavifn+0HZ2PSoA+cudVRNrM
m9AiEgiuLgw/ydBHF5P3jFnBZBWsEM8L3BNKV/OSLwMIz4ns+BGcYSrMGHy4Ph626jJQaf8kPWOG
kbXwgD/UvS8vxzMtgF89rq0R4oYzs6LzjMmqy2GmbFiRTdo5QSKGvmS0GFcEsWNiqphRihG1ePup
VdcoAdbOD9TQq6lY38qiQEs8dghbAobIxlVvRnQaSN5waP6kdsGK95uLtjO85ukzguDabxKSoSko
p97TC88rFPkfbejTItdC7ZskhgBphepLBOAFmj0QtUa+fdxXSoxFkn4wLFIi8KvN613iMEaQNVAi
b2IizKSJAa+W1FSRk7voM6YUC2tQ+C64b6aUrihLaU9yNYnJLRILoldDFt4nY02mMFwHFoSY3+iO
umJE67ZAAIZsa48gEOlEoTpiHdgJMOSlLGk8KaAY6XBDmyXqXDMS8eqJeJ45HuD+XJv+LKPtI/Vq
zOGleVXdptD/Qla+/D2dud9RXkzTomyOaUKCr3KyiUtDbwkplepeSVaVY83wQPysu40CPfGrrZwI
ECNHpiMfW9LojsDTL+faIrxsCoPtVqjkfNSN5iwBLNo+r8gsUsZV+4D9wEVdOcyAbaHXfGUMdv6j
osC5eRW6bMVgrbmMggu2A7vYDa/82vVA89unc1ariTZ9opWClEVp0rhPhfxDY2OY3Uxej2qau0Ga
hkZ0e4de4HN1LzQ7co2Fbc7uMqerKi4/Xg+R5eEUAptqOfdaQNkT7CZydKkarP1HP4jtlC5gdoFg
rmrOx4977TtvuF7rWrf7ZtBfvs4U0EB+qd+ZqT9RyxSAfJI2dXgb90o7w9097tCrE+HbUgwTfm6z
CebHnAGQRFdFpJnHe4o7ojLRtRL5L39Gii3rc1844W9OiIjGB40DrT6DklpyGAJ8uf+w+VEvhFq/
8PaIj4Nz/u0RFxNsFX4cEPa4KWri3ZDKJFP7wLlYxhnztWhGLMqjJsYl3Ls1ewNmdZNN69EnCvPT
WnMiTep3jfw4QQFj+q/nXTDT6RanTFGVMjKDjsDTv4C85JR4nEpwl3BpHzdSu4nklSrTPz3OG8Ni
I61xmolIphuwVNc6R1A3pSDIDMXD7ruKAPHxTNJEShAjalnENkVRmXGDZ7C/D9WFqkbEHnV7Yqs4
noN4s1/BAW9lCQWF8yCn1z5PLKwO+5GSpn8mMGxlcUuaM1hZjHe+d618821YVm/Ag1DA2BcKdama
21id9JDv0OWeAWQQ8UipauM8AsaT/R1dEozaNrKAGkbxP9L8V05roczb01MVPJ/F2E74mMwh12Hs
UPRUIfhedLNsyIixbSti/1JeFY4mm/ue1hh9XEk7+eTIZXG+m0OTWA3ZfFrGUem9GtlmFDu2SAFe
dn2QUGPZxHVKI5iw4wwJSl1LpVsEAdwdqLwh6GajYNQ+tw+96IW4xcnQrn+LD1P5IyTOWUbRK6I5
tcsKU/BB9jvfFOpkz3tomPQaHP4RUBvB6BJaqo51NmEPagnL9FkFz6/kEQZqm76cqHZ6Tyrb0Myw
iXvlvA0H5PxWOW1OcWGJ3KF2dUwdSReV/QAfwqHMhvHrBrSbkXnDIVadi6XmxJqmvri5vJ+zTrgd
dXj++x9I90yq9gn9CyCRsWSOHoKaV77D/hB+LMqdaklGzuHxse27l2DQIw9h75aIkrsckxYNR8ea
VPwRRHXr6ouv3zK7MlNx2deD1Dqt5eWQLSD1GVmuTTgNt47VL9f+VJEMjr5o3znFAGv46USNJE9y
qfN+6R5Cwjq1/kDzHSuZqP2+8vjPQcBGtuIQPk5CzmBjXRkdQfy4pkf+WeEIQwHCut9nKs3YIj1X
OLDOwlgILo+O1D7xSGkLfi7b6va+akRmXz4T7u7E6Y6RH8GR3DODjQl+i6POo/1m1pLHUWorunlf
hnOMi7nuetUhsYnZfysJDwTauLD5nsD9SekbtoGXEZ1j1ofG8yPX1EKK/9lzIQKtw2fQaXF/5G/U
xv2athilENQbCFXK3fNmDcz7uKbqDvBNrIvD3BVfEjbil6QJE7epv70obMAovKAjLaTETS7vnrl6
nuVXRIO3evW/tuqkXXzte04o/V/Ag6fVcb/vConOJzVwL5JodXj29c+hmf5/VJpkqia5z/nfPPcP
DBMFo2a4vecXij6PXGAkAcHnuvwLFQ5RbPKhzMgZ4cxzjMvzPN5oT3qHRhUhXUl3CVrO7nGuC++6
xWlVmlwp6Krv500aoKoqWXJGwN2HA58zEdsG7AXPmdz5psTVUi1zL+gZvK5dTRiG7HGh4VrHP9Lu
ZFtvtJ8ljQQlQtN7EG6SyBFV16v9/zFjPZ+0JHFrQ7LnUg43iwQxWrvaoTDxsROP0t7zSHBoE0qT
VAKP0WXdq05+pWU+l9/LgGzi5UnjK3AUrnrWuToXvvv6qgeCRE17vwWa/EiihL6l60mcNlEo3ZE8
+UtArpj4qBv03qULYvZVdO4gq9tscmxefIUPJEFzT1Y7P1dc+idXtBmCWC5IqXMKxx1cNtj/nlhV
0cEEhS10f28u0cwABWqFQ9SfSzLJRt/PKK4Fs8AwUmSzWUXD4tPLwy4TT6/kqb0fmDXwEJxE+yDy
4DUhSBdnd27ULu/Kslo2bujVIoCa0mYlJhALaNGJVejPm7Gk8NoMEVJ7G69nRbOmiBWe6YjYYU1p
L8h9zjgikaTY0blAC7Q3cyCjhiwzWQ6g9RwC5svRdEHNixr3zqxWQ0hcDSyXp0n8hSD/LhvxuBcQ
n78Gio+Fi4SIPY0cjXEcy1t4GV5/kz1p/XM7yRff0nWizYKO99BjwM67GPlDsrUcJeE8LU1lP/Sz
q5u7q3bRVZg8qjjJAZr9fmFgrSk82FjiGYYWHfHM1RgomeAnoz2lAzJFr8fLXEo8kdynbY+H13Kr
foaN1W6ULuQ7JLTyZSKyEPOCdJLKNoizflM+wVpaJx2B3TfqdeHLibxq66baM9HCrT986mN6c/oE
x+RzhpP8jQJ39bebnYkUErNqVxbypeQe2SeulKwDab2lGPZmO8/E9dmzH/S/uCT0MiW+KEFCaFKO
ce/wvVWvJrSvrfBJb3KqZzulAHSTUxEaKRRA3yuVKB82K+3GwvdrzCP78VAI3yuMQoSLg1sVAUDh
19ZZGiLgtraPNoFm4Af+rXrQlbCbC+RhI86E210FEu2HFYt6wpT6lecJIg8peqRWYQAoq03653PN
3g8SVRiYhXWeCmG2JuX8Q3YsO3kuxR3tTbVpb9wTY+TX7i+eV4TMtacjh+8Oh6RFBujotwpe/4l0
RG18siazUqkueS4J3ry7TXvVTMTPgnGSez0YHJz9HaZWpCgoAjL6+t+zGz69LokSWVKjHROXQeXp
QnXzz/Okt3dk7qwHykF3evS7QmpVtXhtiQ7MtfibR85HoqjSvflw+b/ndfGeyDA721qcRZRWfkOW
TyYG6gqm6XMgrMNRq53Kki1nSpc6LbDwvXed+ZZbK8fGLKUtrtOBcxb1M8fl9JW/KQmIHqYDzyJY
ozvGTb35+hmLN6UJhcGrO2YmuK5KZsR9bX2zd0AAo0ideKErm7QdqdsjyXEIrFM5XdoFJx9/BII3
iK+VG7OCwPj6RGmwIg4u6mFvMaolYjpqSi+/kW9lcIGQ66xwdtN/Z2XSKNBzWt1UqUOg+BlbnIhE
34Jy+XwVpJvHBJedTOk+m8Eygb/Y8GhpU9ZUu7cHkc3VcougsglS8nEtxTxiyyLM1sdW5JTxbEG0
3YInOLNkWdpW7m50UO62r42QZ0uO0TqxZp09k1aRqni7QMW2DGmL6yVTA12dKzv3VgF8LjThfc3/
GYl7BgnoJbr8u3MFAkc3pcri5FgVKpulcUXg91gXJ6l30O/9BCpjsmyxOPJcoJZJW/bhvnm+9Ii1
+T+UxYjoLk+VmhjggQoeMzR4sG9TpoAGegh85QVhqS03WCoN+O2JXKH1jmyW8PlnTCjJ5XqhYmYQ
MOclGVBr8EktDWRwYDEdZjEHgdt7u2ofDHZ7Gik8aXs018hIMgXBOn13uqL3/OlSNS/ZdqwbMtbf
UCYiJAKbdZTNv2LpIjpbfSBNlhMAC+qRl3ZhTifmScdCixf8l9vjHM5/I84FC0t/EUJpMWtnvKEx
fXixGGZYOskHpo9EZYQoH3Ngzm+hGdncP8v3QJnUbVKwIe6a8X64X3j54yAw+XpMpzYM6fl6mh6q
cPTpd+EbA3bCayWybKvIxfEYyk+0JPKUSdiOLDGJiW1ba+fljmxHNrn1abhiHQ5EzbXKr8swTVbS
UlkTFsJqA4wUCFeOhlY14T2KstKkDOuzAV0ATn+BaNKu+zk7oH1Jb5uAfOh/C2dSgM1JJqpprkCq
0F36zkNtNLNwe28iOWWp4T9NR/DSt1CnR1tfhmx9lGM0TicvixpDVMFvrVfmSk6HDqvr1in+ljkt
L5BnA7T9G/AZqDC8MiNOzIs9OctpjbW21/OiseLkNpLlGbVbOtVSUnl8Sx/84Rx4be5JVM9ZfsUg
zL+wwbXE+y9bXgfw3YMx+QJMzrSfZ26xZS1xDUPrw3GVlOYOOnOheQeUuzVSBSGzRMqr+liFEJh3
URYuKy/fSf3wMZrGBVF6J//mpGIO0ZhKonWUEoOTprCT3ybR3s1d9wfFiEYlxALiqxTmuZAh4j09
BT0mb6oForHv9WY0ih2xfcHQgV4P7k/GmgVYm9W87ZciGGqbCxs1vfBg3RFGqrjlWw5Ax4Iqo0QN
sJQMXabsA+IWUUDstAC+qRVMFw8uBKq849ILf7q2Z2Us6bQPrLAJnMY2ho8XM7A4xQHFy+0gwWzo
ZZksxoDAhzvBMRxdVF5EOFgh+/7vPdiGDlk6PEPYm+yMBgkB1wvq+UzNeKYKrDuhjjv9ahYetuE/
6K7IUaeB/j2pOgmqOOFpZyYuRxtGJLTLMBILRQzqj81RjRjlSqiTNbbi/lWCLRCkBzXCt96qK6rk
yPmNCYP6tMmoHEzGicMmy9qbtN5ns0H3Y5B39fNV0U0D2QwHTzMXDmCJGS/6QMY6BIhUn2uBquJG
zih3pW01ybuPtQptzqQ8Tg0ZkGaizRFRLd5cHvlEtpMze55iqPjyeeC6co/itix/CVV2YFlMEC7z
PkJkAdUkfnUgG1cG/IwgMQnQNLYXm1m9xdsQoFziJvYUz+lgNwjBhQfS/oVhjhlAvKmA+iy1UeHq
es/QsrGwYdHaqz3H5z7ePWsisuwzIT5/0fPs0VgYX3vZUMXxJRsDchAX6XOnlx2iWB5E5gG+ztZf
F/8CxvdG8wRkcjZDNGc7BGBeu6b/FhXq1nZNajwuaSPqri3kiRRMwC8Ik5DoFfLnRxL7uKErbgqy
bbemKbm2aBJSTfsHfSKcIa/nnU1+aow7u2v75Ir4gRSMZfahDI6x9yB7CglDC/M1isGl4pBARugN
zQyKAzGi177MDwwkqcmD5433RJK4mibMc4rGLfDD8M1683n0Lv2jzZXqihyP5C3F0daZWHw2wayD
PDhDD6zjiXIq5PjBJZoWw3kN9p79HDfVPwgaDfpdMZud3kI20K42mtX5pVxdbyTUZfIgJ2Tx9L0k
Rdn+x677a9yN9XBe9IRcNR1q2W3Lt2ku2+FFe7+gKZF6LRfTdYMW50JIN3yiwa9S2D0OrryAR0vc
3O7tPDjR1TRWwSAciPZFLibfZ5UywiB7kOL6U3JD/oD7o6GbIRj6gqwfzn8RMogP+CS0J5zbx2a8
xIQMu+Ym0iX8WyNCUlfCyCH0mUOyrGWS7d0j8m9Zm8+3e0o/YvKac9FV4N62uF7yxu0F+Sra//Nn
P7H7U/jepAdrKmZl7iIW5rjxLuubQS1kiW5jZ57bqKxKfxMti2INwKbNXZeP0J7Cau9ES+zXXhW3
nrXWogpSfTOC1hkgpk3utIoNRUWrRTTEx9CFO0u94SWrpTuMSkkxweQWIDDHF5llLD5vDBfn34YZ
s6YWDAdwmjHY66a1jXHjVHI+h/Ey4sevJJEDM8OQLoWqARKwwFhgpWMabD6di4iDs/ilU2D0TPoL
JD9l4xN9vXZTBQkxF7Ba+5kk8+TCN8O78l8u6RQawTdlTM8Ygu69b7aFebCVUEz6udKEf9WeYqo0
hV49PV5e1A6Kmrc7agtZYDnbMCBo7OYdDeWSGgwM+1W1nGp9WavHBmrl23/P8Vd365kSPKAuH91T
SYIuqevIjxBTuioqwH4P0UkQhvK3/Zlc2uwPIVGBF7BTGgVdM/IlFx+dkJ0jZyh08LBMww5aEkbE
D11eq3PF0NYdTMFCq6aEMrsJ6ZECf60LokJVm+K7OVTZzsijPwqkvMBEncv+DmgQzQIuSlkIwje4
I+8p0A9tivbRKEoCJ8x1cqzRtzyu/pEA2NItC+32JBKJUeGZnp7mhdI3VA0xa/1CWM/FAndKjaSs
cgVkkV+ObM/rgudoWWi64Z45oNmIEFn8gE/lL8WIy7+Sm/gWJoDacqE4l6ol2xnMD9LgCYFsSMtw
pvMEsD+Ni02FFjCyhyr4RNvHlRb6NvQCyvHPrh5gqpTFRRe9vTT8pD740T+jfPTLSRlBhzlZxyf1
4tdGvTBrR0oDhbm04ck/4ldsu1s3xCEWNEWOjAT+6lt0Al85JdEvniBqFCvUy9FEZ7jigZbweITV
XDFIPb0mImWqrkt/VAh6CfDua5JcjzCAaLS6Lcga+RQjxBIAjQqBUaLPlKUBdTlT/bbn38llY6/g
6rCMZSNedoNlsd5Rs+iubJCtm0OMux/SPryfPWuVZhHZW153n1O/jVXz+7u9qq5J36aLx1Rbl4uh
BfTBiNLtDJvnj2G4Q+DtNTp7c2XuzenXXSVOtAdIilR8UhubV7/x5mfTOpmiNQ94SS/BR6PWoMah
LmcNVuwL0EfNfz4jehtelE2h+4Y0sajzGMAfT7DTkKr5N+mUDC6pmmKweA0RNmBP5yozvwPCXlGG
4rC3ra0wvUXnhG6AeRGGNh2631z/mhm+fRlOdxsxalF8K32rwcFvgxt9FHiZz4gzttxRV5onCes2
VaZyA3F679HmvwCdqqqRm42bOSSCOu1IZDlvzKYMeHtrdGjXOlAZ/hD3xa1Y0516OuNOTXJXElsA
Bxm9eZY9ORuPetE6xfd9ihVCHKPiphKcKndUWY3ffDJjYVcGlV3vRdENXvwKEFnepuafaskLWxk3
gCkDqHF37ZMqp6wySaladJMjvjed5Eq0CAXu+AqCeAXetHsYIFBDVTODtNBPkAzXyFdhvzwpw8PD
ZON8ViMcr/z5hPT6sbe0iyhxPn1IzH7qdZG7rEHVf7mAm8yFm7e3oMlgZPBiiujLmz2kXiR0/Y20
wteAa7Qdn2wnYozs4aPUFPY3zsk7g4j0nHgTSLJ6eMhSe+f2p/Fsi1eeD6AzTAkEco0J6lfsG5iA
5L6L+7CZl24LGuBYEkMR4+hAWoEYQ9uK4TBBJCen/WKoNXlmIPwN4zikHpd4WRCliOkLKoC0+XZH
1AWUuP4LTxBisMmvcc/nNmVFo9gOAmpHbbVvYOos6JeoiQIk6WqaaXhjr3dPoFYd+2vdFTLQFrEN
WXUfuBPqRj88n/ubDZE8A1cm0yG7oeD7g8ofFpqRTmZWpYlw96wHSI0OLWmm9zhK4TyY/mn0RrxT
q+9xRMM1KORIIu6nQpj+xwKOnLWTd9RoaExikHuo9hkuq9685f52Hc1EpyDB1HK2I7gfCxui/spl
QEuWg4Ohn9x2jttk8EXHytCtK9EZEMqbXcABu3deqa7lyoD/FUnk3W2oyE/7lenSLVDOMaDtuyqD
eOzVnxVwa60o5M1iJzP6sClloetfsLqk71uCsYzBLCTdtxEiLFDk01zZ6jUfTpJGokyFmntswag0
HhIkuS4MRMeHYhZ3GVNxRVdlsIKs5d5p0Lv2A+hmkcliNTHGRM3VYBJ9aHBz+gMXO9xaiQTu0WpB
xGDn7C1krXXR/Xp8VE1aVxvgXBFdIrL26H3WwsD70FnHmxSsHRloafT4Cpex8c5O/DoZ6vO9CEFT
QRUJOh7x/FG596rk0eS+flsRtaOK5RMMW9MqT+mUey90w82YXOkBVsZrNxlzCNLfrlVnhZeqvm2I
5o8xSk6x99s2LOrlmERLzTdlgfLNrwNenuAFPl7NfCySG5pbe3C7q2h9Lrfr0YRmA4hLkUsllBUB
7yfhsaYYWcYlxb6T4tFgR3ogARmAZZtbA6P/IB/IjxMq3Ls1EwTB5CH0kCxifF8sFkDy6OtWL4v+
TPugRV33L4tojQFbIgjq01lTShOSrrIW/h0LExZca6PJQfEbb6g+wrdv3CYgm9djZMGREOTtRy3r
BjoCXvGgtBUMIu4yjoAIoBq8+ngr5bRiTBAOb6mh8Rw9mQkyAOFwTg4wP0Bsjw/kSiPhiTcnrMrJ
G9Qcy9nZhS9fDRJ0QSPE+l+hoP+FumqsuN1wT6wmgcZzVnHeDut85HCc+a/IUTq5c1609bTET7JD
eB5SO6iQ1YjapiJ3AFS6OFc7x/kEuIXPM5qnPmKuEnPgBNUj6duDZ8Hx34IFhv9ee7fJi35Jc+nq
GwPK0zSocnL2P+dvnfH30Pcjccwzva90nwSvi6SAas+0bxIxtvM2nWosNP4W5Runr33zWpV+sMk5
9Albx0udOGzHrPy8/W2eqGv2pGMGQR4BE3KRvfwZIWbmRdrZlKXrczIutbVs3AhHisdbHCoFVb1N
IyIzOevMjfCXg7H9MdakbpUio2NDuXGnh/wVF7cznKKYqXTKygjEYtu65fVgMzsozelm9R2GK/BN
yUwCsDYJQ0AP+vEqiX3zex1ueN56wsJDyhTuBAFeOir3yc7g4Z+SX6k/aavb+6d+zRff9DyjImJh
dOdozf6sWU1+gy7IdK1k6Lit/xCs2uDHFxd3YjR783CakpXYLImW+Tn/2I5cmDKr2+AAmsHnBfFV
DZqaoa77z3+j6LE0HLxrrO3qvSFY2A/LED5iBxmDw/epK1wa0/YJLh5sIuWJd8w7o/hcOtM1YZwT
XMkqd6yEoHSZzG4O6kEQT4YpS+UPW0pskipQKYYprCvSw1K9oMHMHhQ6LcprdUeABdZmEEZTgjeW
oaqmBL4nfeKVD3iM8xki/nQmmkil4jN/nkOz12BA7bgi2tIPP2MXJ4eG3LF7nh2PD2Hg+4PcPQwm
dDF/YxnspdW9R2v+QNm2zfp5h9ijS1fzpfwdlyqb4Q1r8iEcsgb2rNIvoWMkE3zngc8LgzxacNd1
izliC2x1uLn3NyH2L+gGq1g9tpM5A+YERPvWmy0ASANhO+JA9YyZfD7VcKQepBe9QQ43F4lNiK/M
Fmmf8P9h09mrQY464kNtSJ3EQvEymHAhdF+f84m+Eoh6tYyr/foDIuP5vwCJw51tkuXUQiroaEX5
MAB7lZj56y2YX0LyYamnjmv4nWFkMrNTV6CAyOygxQIKz7XO/+z7hxvMQOQ1Xc0nTTPLNOVmhAYc
bzlv8MO9Qqes5iYkr2AArqPMqBYm9cTQQ+G5UQEl/zsOQ/wI+GL6J760DqMTwaEW/XSBPrZ3tO09
Klch0eM9rdwANct8YorbKxgb8M4mnOgte9vZViUzVgbhPi19NUizuB8Qpg/Uadzx+sUNCJwG8C4n
Zdfpd85PoOXAG8YD3D/uVROsAYYsxrZg4RPXZOzbBLcaGbcH0xZcRRToxc1otmBzBm8jsgd3S1TO
y8wPJWyIKW4Qk+6rGplEgHqhSpsArzK5QLZ/VuuJ8x3jKzC4sPeQya/CZ1EMCHhEPat+ZX1ki9P7
kyBCytVNfPpC7CpDo0O8Z/2S8Tdt1rVppZjxqexfKNvVNq5lZhPw/jmkW23NxNII7ODiMdFGbpdh
zTOH6/oYDi29dWsnzz6D7lbKWlvrJVhGVqRpO+YLQKYtBwfYfQRJKPcr6qav8sPXEFv1vOyKWYmP
VtXxuhzqY0uwadz6wBA5by68dFc5pW3SpQoCsps1cWeMC32U4FsqCAJr4JU0z5QAv4XfP/qMF0WC
A2lSL+XgCUWOSE8mB1iTxUbpSLjIn4DLDIm74XAKUX7WD57MInxb+EgOUYo0NbtajUOiBP/dV+Fi
LGC0cj0QnX03zpRLX5zHIu4lLUgwDglrvwK91ONQMz+UcdW2dYMF+ZnOyyv9Wn+slOw3/fvv8JNC
HmdVBMsi3OFRoL4tcbMZt6zSjtOZjvdUVTZ/RDtGB8KjiIFdsXjDN1V85UE5P8rV2qO2a7Z70Kz9
f4ReviMkbGuI/Bw0PJH0CUL+lwW7GJf3EpILC316T9Lzu1m7t9BfKqTWUtz14ziqJva2mia0DDLi
7Tv1rP9+ESSryHuYp1cXD1Nhv9udj5IeehY11f3flC8V3sFC4IEUwilzPw34EmiDnXeaoWH1IO1W
VoN88Gy3Vc5T8mDRcJ6y09nXO3WbmvVNN59CMDDnlHwKh3jJ596GSZqaNGxoPbFq4JFwVtqVCRAu
Hio7KeSNYYAkUH9U/fRU5Pg9QrAEpOPA1+MtU6pLKqmhBPQQ8k7K7XjeomrhbtIgC+feVrUzWrI8
cnsj6DLuyTZDnt/iQU0J98OjskicRlx47icafQNke7+aITPHqNZf28rJp4QgjpB/7IjqcYNp/XZH
nW/F3hQe6A8rafT0IGjL/pvQUOP/hQ89b9OvVk7A86SvvI/OdmWj4F8qQEu99uM60yzomL/ntHCD
zBq8dx7gO60wuetcT1rhmhe9uqv9+amuJvzTQOvzayNhmmGVQSELySq7FbVzaCYnY21mzC9Z3efb
w8B+zNEieB8jHtAvu6Ze6GFxWhduNxZwVFL910AJnWacGx0erC4MDFbMLVmiaUgGz2GTtaSoeBu9
X4EyjHWu1ZiMF1ZkyNM6xJrx2Sb6KOrwGJfSDy0u3efRGrvnp7Wyvqmhv+nywEUJP0nbZx0cYo7O
8iVKqD0WdPAgLXJSX85YUodob8/GG/gCowgbcK82/2Bvnp3gq+awaSGBNXnMSgC8bvQCHiToedku
Rr66LbCl+pAJICuzORSRlzLBvf3ItKUaUqIp6YwG6LDbc5ghOACqYkY58OztNLw71oz2vfU23w2s
O0fjGlyQ5kTUif7NWazdrO+IOjveXKWXgtbOq5gV8hL8Ew76PXF8HGksVkUVt3H1QgdUOtqGaBht
V2Ng83OpJVUGtKPUQukFw9UWDM3+I0Ib8+1Io9wyq502rIRfr1DQ8OjNX1VxkVJJj9BAlw+Yb0jt
glWxiyfilCyiV6NZnMkflkDU9tB0EDDeeAIjqaOknv9/VuGAB30A74YEntKmrDQL/ISvyfTodjv9
KfZu3pTDMMCWU+58yMmcOKTbwM11BAeoCeKj3dUr671tPis/RnZqFEmytl79+m4T9PUcIa4IpGB1
um/j850EmdHDFKvHfi89rNr6ZMSE0/X5zlGm9ogmqWQmUsy4fyzmRYFCe2YJ1C8I0wxnD3xlrlZa
ZUyeg8TG3ZRvug+8jrO4womTBV7P9gyaQrLFRZjz3dQUdnolHZmtIE6/BnzVTwKxVTEU4iiGajEW
QLJwOhzoliVR89swWWTnPjRuO5tjJqaxC24syFhPlCgtPy8TqLDDkBMQQaT3rLa616MnsHgo2uiG
6xvc7nvTK6IT5PpRHBvtbpNi22hcBNnsYAF5jsULXU1BMCMeqRmkjflqpNEb45mpjGFF6/ZGN37M
WxJeXncIwDB11u3U66gc7TgYG32jXtg4Pk9GGAOdmIsxKeg5OgEHB4FGvhAJyzMhyfHY1qD5aDTq
hkK5SfDrFf9R+VaRhbcNCSnfaLN7zqfgxXco3iQDyxPLri/rAvEbjSwJat4hTtwYz5MDu1H7qTSD
HcFy94LzVm5haV36zc9mRNsaAUUcnNh2oZ7G15Vl1rzzkf3JYtxLKRa6LhfsaamXs8i/GhvVZrL0
UTY+7BEXA1VsTkaeDt3f5fP6N0sr5IY+Y/wXUDWBzHbGvawaohK9cfvNbZ11/vanOFbJuaBwRiSM
5Xrw9kz0x6cdkAScJDE9VvUaxlpRryYpIItEIHTjOWSZbq+w7mCo0OuK6yVrmWTlk20ztTh64P1s
bcsPiu1ak7oAfLBuQbbD7tnIrfyn68ne1Cd4/49JTwxlCrkUkMfEqkGo4NFOw+Izz4ja7ImrwFEp
It4VwuFbH/esIeVo1tEKrM8uzFmZO8jRUQyHH6Fq0hHVVKOFVNG9DmcRBZOJMsCvAQ76M8EI/E0Y
c3Amu1uR2RSt5NZdeZeSoSes49FEgY8drx4R5MAM6rEN3n3T9Y+PE6j1ME+463vAEHQyOuLbdhPy
vft5IzYbPhFMpdIqI5Yg7/LePwR+RJbY1MLDYaY0cEmmxBJVMKpxoWSYKwS+e9alM0Xe2zz+PCXt
NXJdRuC1EX9M6qFeuDo1EWsxlTkE/UzcXP4ZVg72SkA9VWr6FikEcxJWf0VzMfmTYLacAGODSplt
4jlWgngRoualjM95ubVfG8KVLJY2GhTNysMFihgmQq11iPaaxE2cuBdJiecLJ88ceaXYnw+RsMsl
ZsGu+N0BuO00FyosbtKJ5G1CkFHKvUeQ2qbkHTvpLYza6Pl7kjlGFZgkkkaQmUOA+aBAhLLYM07N
xlaDbiqhyQDwE7vDCETOabMvNHVcD2tGc4XwAg9mwxQUGHsErdYqoq7hY6JqyVisLBUwFLcWKGdY
tmnv5YdqqvZK9bt7Woyc3z7vRk8rzyBz6q/HC4xJ9QzBp7RtSfa45etdwYrbVD7ofS0aThW2/8lt
rBfnAby3t8HCWybSotZqwGzCk6KZ/yBk+AUqgifnRvE+uOTwkYds5vZ84UnloJG09qNhRDGqxuU+
UuwD6wVCcjn03CI0gKCUWyQ4mzn/5ZX+WAfc9iYeDIgdY4gp/O5z3hHu528hkP3s3B4NUpwfrdiA
UqB6ZljJaddd6cSx+vpmygbjPQBnPl+wukViWvMuC7ueDku+KC0iponARYqg3MlEGHvhCbBjC/xt
rkiRBkKXivyxO1bBZZt8pXbpww8cukSP7lBB4s8q/oRCIbXLjYrhj1w6Q6P5ii9LlZ+/icnCB9G4
pnmjqA993edz0WBGTF9r2axvRRbOzwAIcLGzSlvdr4ZnLDnHvyfgzV6DRgmG/Zj/qYVyzow3SXl9
GljaNkDtUIeDobjZDp053fhMY5C/6Wd7rnZwZlYaYB6AJjlmo6p0XsQFlRG/JyiLRPuleN/3lL0S
/0Hw/7Vc770z2/YuEeHduJ9VLUf4j4QM51mtZG4Yo2GtaMdyuUhBTFzd6+IsRLsuPj+M623gQEyC
VEq310rmn0ZmgPAN1UHRePtW0gtjLlJz6qORDtWse0rZZCKQ7ZJns/Xev2rS0m4G+Me5CmMjlyqe
Ih79MLGiI3KgT6ukOBdfpauVCtPAIMExqvnpjd8jCk2fHFNvuXt9ZFfdvv07Y4boLiw5RVtpU5cO
CGowPTW98w2z6sp7WlNkE1HyCzo8KKUwRugrfWCUTDOgVmCH9+KsFd4oYrOIg2wWzhNcxIJJoFRV
TzBzTSt2IYxopgFFtzc7xGExF0PrYPs6cHh+qlXBzQsHQt20wJ7aMVW5q8EG84hwNagfSJs8GsPU
kgu1U4pfBhcQuJJOhfPuRuXsMasxh5MdUmubCePc8Rn3Zu4wIWvkcx5sqUSInemrtPXzvF9I1+gE
PzQz7tuPjaRcGBp5j0WbXBRVfrYUw7qOo+dcNhnMWHjC3jZPprLQHCbRE0bPVRmgj+plvjtCLHX0
Ml8hxHlF/aKlCzTHbawqoZcbywOH0wfVkyLGecx5BHPyq3ffSaLIP7P73Pc7iY8CQfmae5c66G8I
/TM6JHtgjNIZUv0WKEwskgO3MM21fg+UyfnrGd0HCgt7eSolBYRp/5GPkyB9KATn/lWXj1V6/NJa
5TWkDJBG4Ek/LVGnhJc8d65WFJi9EhlkEyO3yp51eJs5AYQpXOpdj5u6V5IkQJrT+GMT+HA0p9ZT
wYYTA8AYP/WpxE6N4yLoVBGvShwk21AYiu7i/EMAVULvKHVa9RJBVg3tntIwLrEHOcF1GvSukTj7
Mz73SX+FDDO7oZKpghnRmHwK3qV2wWXfgAdFUf55eXOBapn0s6p065KhGg1HMqxRMWPTOYrj47FK
LiKE4Flw/+i1XtQ2sxRfPCEFHe1NPT7madnmqLI0p98v11GO/Us9FEGDIyS0OzuAG1QvHowjPuHf
b1Ea6jsFG2UU7m6Em+cdwIXMSHw3Ufe1viP0/aS1MZFAaF7wTzWRFapk9bQiQWuwnTYGwTuhOIh3
P04028A0ovmIgnGUq/aPiITe1rpEacmlfz6c+Dh9Jd+3HoUW/OVm4DQTE09oZy+8a9Ns7rkZ+uo5
DvDaFdbgwEFQ7xxxa0KrZhu8hFv9dol4DN49tYO15fvQpK0/142vyArKncfGn1mHhSEUivDZ4loF
I+N1AnpkOtwMurzONu5CiZoieGvbiOGhQKyEBlI3AoetGRMO1sRsa9B5VVOJEgqMwq7t/nVC8MQ5
i5ZCEB5iP163o/AOISeZ8ikN4T4wDt58jzoqKakLmg9cjtC7PQ6z6t/gU/AyLmDWJZiWhTkqWxmy
2nDJIjChOweQPg7knGaxtDea/cDghaNp7tHJbxKbGkepPSIXWBU7lGUehRUn15sFNWscok8bOkqr
w7A02YqGF9T3pL5xW33ZK4FwaYKDhN9ur9vGqqE7swIkg3NukWoreQjn+T8pMusuTUUEx/C/pwgT
WHJPKgGy/i2S9FKaXyCnIF1aNGeVSIXsW5G9TklyHJI2W7bkAmJnSl2n/1NU+ucMd6vfSKp3t68G
YQ+K7St6C4RglWVsGREhVVONU44+OlddoqwkCG2+PKa5eVI7B4Nf2IAMwWa17yzhHiCUQ4dVQTUo
bzBZamo3cVO8IcbGE3HrEqpeIupnsQ+ieVE1NDXZd15A/aEGOEVJFSGE2Q6yKFbZVihEh5FdYxqg
v4DKN2yg2MIXBLShUgDq9MWgxgAGtBQfvs1QP1GuyDQ8YvGwf9GFWtb6KlTK9m0kJFKz3ZeZKnk8
LEN9vlPgdzTe2Yg8brxixHpp4gzZeCrdzup/2tNDa5qStb+LqYA90q75WMswfPsjii+HJDwBfFE6
m36HVzXCMmwxeuvnw/IWqy96qSUioTE/SD8covwOPTuXiNXjWI8AiSkAibbwenjHRKWkVdsLBFeL
zlMY3TXeqyW4DyHD1GmeGX1IQLI9n43Uy0HYGmInrESrACh9OAO7rDMevhTWLNCuR965ymDyulVq
yAynjCPvROkxir0J6CklNf5NVtp9f21acgykYjNNNk11gtSeYp/XTfC7xUS147/DkzmkcnKEkvsc
WhrazWLExLMq1L6pWdn5FPVomhlg++RSjB7fRMgk/b/McyL+93sjsPztBqsNyLEXS7xDQ0v248uR
pOs7alQzmKRgyM6JET39yGDox7kQgSy1bSbDNV/8TbRQD2LdifubzBVb74tyRDTWAhmt1DRhIxqX
rD2nv6YXwpohFTpALVqYQzhaJW2bIg1zMkwSET5n1ic6jlML2JrTlV7XY+DcMhSrOWyBzyyKS7Xc
7o+lhK5ePjMI23xKlHv/YVwVdWBLnGizLRkUxXc//eazdbnFgN7YPrfYTtiBKjCqq9y/doMjVGGU
tp7QII5Y7luqLH5JUzvxaGPEPrYCtz/b5s6SLh45Pbk3UEA8L01DZwGQTzKxGHMXhnIoh98Qcg6p
Lh0rOqvWV26GpIm7W/5Sz+NisErMlIF3yQi+ookYx18WnXI2pURIwCkJEXu3e5gNkRCQHv/YQqco
ZAmSKSrx7X11JPx/RTqPAqu9S6DSTEnkcXYvD5nL+3uLoAu0nxGXfidmwLkwDXS6mhmrm9UBg3XF
1ZVuKltf4fj1dCbGN2hU+i6IyNj4vT5emBt2OGRV6fi99yQh9yX6nex5yT7wzC9dUxsWcd+hlBG1
usCsq9FQ6eJCiMpWT4p4UoXlbIdqkZNlS8fRik8ElpDhKYxP/3is0TedeJH9yKaJ8/SQqTawU+Hg
y4bauOtuqawnjHIKjCZ8ktc5uzIasqtmNwbWM5/MSGXofniiONloyW8pUjsX31WmB0cgtykqx1x9
XDScSZV/qPRDIQ8qbkvKO+uNKF5BfhOZXJIOM2sXKX+Rh9mBAcAZO7sf1fVYceQtV/gpWCGmQymi
SFV443XHDATyaUP3lXLXkbGfE0rkujDnKl945Q8p0EgwwvIWx5Tw/ZNsGJTWEmbL+/pfXu6tLk12
ZH8gvFqTE2pwetdoAcY2+Klg8jz6Z0kW5HlXNlWZDz8lIalAegiBwKRA+vIaI7okD9v+DbjCrPTx
7eP2wWBf2uN0CGLK7j7YbaI7KUy9weRx36/L88iLSsAncUGvU28T2hTcmyw5zWVVGGBDfnKmmwpO
KH3YZSSE1C+anOH/rauzL32DlXLdHhdqR2N8CLSeTivlQgrY9OmtHQifEfl9ndL4IHRhCgzMA8nT
Y6O2DlBzIiPV4ja4IxA3o3aHYgU1cY62quljctzC9v4QbOTy1ni95oxWMaQuZKXYfiSF8l4kNKhk
hI5onh/xGYJB/ufvYFkf59lTyMyFztMhuteI1RCxl1JSTVHaTcJtwaXslGB+FocDqJ1lMrU7hR7r
shERZRRh3vURIQ1eraIaYTqtqrL2pmPt4oboGx632OiR4YJgHx4wPK4D2cSss0TdVKVQXl+QUSxT
yXoGChUq5p0nWGCV41oHDM/ashWifjAgfmNsar8MI3Lk19YGJh7gast5ziNa74DNuY0CJAT7eRQB
JYwRhkTlIMt7kPeoCfxAPyFT0h3vYyLZKkQ7OcbOxuYe7rcygiJbYMnriu/8UYH/vvA5/8HhkD+s
lEsEftsW7qtijr6NxlNSlOCDp7l38NcOFLqVqjlBd/d1Mf+kHWbOKRV6SHNzvNh2JtHOECoW+Hn+
sKXors7RYp4uS8n/W6AW2DKOy86LyzruO8BRZRvT06Ioh1YH9C+xUaktIihtLDGzfcgcMERMSJ/J
jQCvZK9PfTM0GWhwWm5I9Jt6oKFC+dmKtwJD1pFrNETSYY7+ufZsa/0KSIi5AL4e3sbH3phNovjt
PYIpTv+naZB/D+zekEUKvrdQ8xdxhgnGhIDJPKzHExy+6fHIUXHCfipf09lwA2Duj0FRt/7iKJi+
E9CIpwAIY0U9RKtA5HLjTUzdnlU5Z8c/IeVyZTxk+hsxgMh4fu/D3H0jDMaS8abVKs19nLOrWsoH
cwMLeJK78q0XUEtmLS4iY/wyeQw3kg1g/7m+SHjXiN/uE9EB0r9iE+uVwoT6ilJ6cEklS/NZ/cfW
tnoqJNkFGfxdUolzhhjXdo7aYCVgio2ad9wlSSJfBX9/t3lR6jhxJT8sNgzxnNIg8ixKpZJVQ4yr
Q3775+VjjN4TlNK6s61rw08CPswnHpLJJYH0PFQJPob5smdPsV0zRHcyjip8rl1QXfjeD+WwCpjQ
/e8c/WnpDE884G7JLCmCgxQGLyZiLLmUsQRoxjAb5Q7I6jaEP1djgRzeoiPkiTEv+SNaAaUrFGWb
u/hFXtoxLOI4dsyc6Um/f4EhjUtCwthTBLhEWqqBj8ZXPNJ3JCBcMVEoCMMj+2RBp+nhdsEC8fXP
N3hIvxl33e1q0KXA54TZIy6ZPzHckbVR/jv/qTJUVgGFV1uEhbnGsoTyk3qqs9guXdh0f4T0yvpE
1E6hzDeG49k/mg2qw69c6kWRExor32dRxBPlVaFc2yciHs12DT/5rc2vkHbep+zpr2DbND2FDHEl
1wFtrzxsjBw9xLPBUvgUWKjLaX0Azf+lb9z3cQ+U0Qw7W35Bx+egyhfawUQQBg0g/eFpdija/Ggy
C0BYLKjOqCx5L2Scuj/CRsCN1qy5CZz+7JNg/a9+8k39DppRyXSoSk9VZeu07rCVvOvd1MyVJsbt
bbSONeBSq0IBbK7RcLYGYzFQPnlCWt/lm8ZSzDTzTtLHClFWVGoPJB+BIObLFNys25wLAa5bO6sg
XDpOllctKWg/LkdzkyfacF7ceJrnGtXnBczyrCaTG0DHYkdZuCIgjRDU8OhVpjQZY2eYGkXtuX9g
9s6BLSSZd8una7vNHSRyTjPaXuOgU5oZ+L10szTS+20Hn5ceEgmJyul23zSX4g7BsVlh3gAj3yRY
9f9EviBrbgyHPgQp/TaiFyDOboO9RIRzqvM2TL+BftF8DM5w4uL6EzmMoxTgq/TtWLHkCqaXY58C
dErpjWi5VHYh6oEhKq4axMDF3wNdJOcy5C4H3mXcMM4RMCUtlTSH6ZQqIqlAdRLZ0EoFADbZ8aCl
INHvz797Evrfx5bZQMnO+9c/o3z7aKoNTWwy9sfQpuiBUiefnHytuGhZGC8m52h9SAdCBEANYdQs
WH3Hijx0Hg5M+DaRpajCEKYI2KWs2X+W9A39fgvKuD/MCDNEnKKWjOw5vQmnZ9jkUEXWMKPTWamp
rKKGRqVH49AsWPCuDyITB4zSePxXhbFmRadV2fGiAPfEjJz4pl/EF6asjRGRyB3J4YO6bB3Wulrs
xH+LvvKlES3cxZA/1sUvsiQEdKd88QFrALw0v1AiWB+ZR47xvwcuTkh2MrVNmppAlUL5MzxDqlI2
imfgJWXRyqAlJu+0h0jzUiihDREeALfaPMM4fsAE+PhmEFc0QqVwKbLRRwb24XRkq64pWgx4gedS
MXViieaxA4rm3e5XEg3idqx6c+t+VnShjpV2gsKjaaftYbhwXjMc+2w3tZCGGif8Zn10iwbKTDkR
kaNPwPMEq0QEvVm2lRmvxmLQ1fqlviX5FLJDUw3K/VhQu9PPgQ3D4eG7jA9dlcDh7B8lhMaNjzWZ
7c7E4QMBlx2AMgnLCTYKdwZeY0tXLCa12CIy1rFXEgXCZhnzgF4SlQTo+lrtbEXxwG/yIEUP5j3u
gTEwXhvp9s2umKFV1oCrRs1GC9wYQL3e/L54QMcfn47IHt4XRIKPtIkby7HozAWP9Y3OUhv4OoSh
o8sg850XR9jLHN2AweWnZugEL1s1T1AstHsUKwegXhRZyORRb3FKKgtu2FzVIuz3d7J/eAXefbkn
RO+vIoLkFtjen7zBkmwa4Q6SbjZ+hbirBbyGPIVvbLoeX3z7r7ym/+zjUv4G+nibJWsQyxsLBfN3
rSol/Yd9YBqXZJoIm8q+OuvGVys99qR8yTqAdXnT77+Z4QqCqa/wIeni5ULKnVRP1N0gnfZ8TM/4
IdDY0BIx4ITVvwmmlHUxkAA/wUGkgLaVP8YhuqDaE9UuCVYa82f186rrv6IfKzPilkWPjDuf/MD0
Et5cV6OMoozDv0I9GsSA3IkyKwnVNtSY2LibJPUdnFg2Ii1HWZCaTMAU+Pq6qgZtBM0wc8aLdizG
813oix7q47O5WzATZQfgY1xqQE5rAY9u33edJD17PdM5/giVnH1x0S1EZJu/hNK22e7yfHYNzPMe
Dx9w98CUGv2YlbyBEiJFlJ2YW03sQ5/isoThTVquHdyNJHBtsUnwqJn5EFiEzAbEbM0XRfZZ8vBl
8RlqAaI+EwS8yMoRI9cnzgUHjXiHdvWFluhhJhnq1dX2pD9ENg0sJ3vI/Cy2yf8pTQBaebarSh3Y
QGDRZVW9LneHHwxN3NCZ/teJH2uKzd6cNoRXRfMPJtCZBxsweRMKSj2wZpkI5vTiSaB1lS5mqIeI
6vKYWVwdXSBHcezL1GoSeKbzhqZHEMAs+duD36TVB24TMKHjIBbLvwE45H/5Os3tBzCcOK2D0n+O
dlLkaYHPODiTJI0lHPpH8QcLM/R/yHqic5mV2EWNMDaD5+3jBRwsIT0SLOluk/gX47LN5fwOu4/P
rdWAqWLVYpZzZqFJQUw767IOyzfCOiZeU5D4/hnOyujcD1PewY/rF82BoNBUj3BGymR0ttS3b/nq
uGzg1GPJJziNc+EnCMToWjl/rVl/UnQraKGa0olCmwCF+0RYi+eF7W5DC/cWhg0ROQIH6RJftRSZ
tV8d708YXSOOnqQDSWvxI+OFQnGrU2aFpHb9jX+XxW3WHFWZgwqxzLzcCvSlr006NZI7hNA5Ozhq
37ZN5nEi5DgMvMKhTRh8/NKmAXrDw/gGpQzSXyd7rojUpjPRulr5mBK4zr/JDrUW903Ou3RGOvj8
fmWJrHL65xQuHj5Av78GVNmGYNK4Hvu74jGDsVzzC4Tnvh1A//utiPAP1boUSvOpjUkOA+g+2b+K
jPcuECIYQqVe/5bV7SD54iEKRO2vq/SsPTFC8xXJGLZvjkTdBX7ceM+hYvYMH0PYlITaGAc7Fryz
DZ+Dx4nuF5nAg86YnrJtcwYr2LH2Fm3mno+v5gm1GQTwS/EyuvSFvXtve/tXkXBqs6Eh8VtyocWE
wrMZzRU/AAdklZi4Fpve8/FR/EURBDUN1a+hDmSOzb9tpFWHgZyy6pVKdATC+cgqOkJKSBtofxv5
2l4WACN+cnrSPhqoPBdX0OMUVWEoYQaYXpF6XoWJ1cMXuI+54TkbFPs2kvWD9kJmRUkrP/dA45Ik
43yg2kmDznlz0M3/a1BSVyYRg2/0jGmfyczEf7IPy29mYh9v/lDaXgXWBUSV3tANASQry5OY8IWZ
27jIE3tW8y7cGjdu48TG7DJvpS/VaVYMGcES3+Gc2nqaP/7IwuMi+ucL3VRqdHX3s+DAJE9ksUr8
tBS80USF4G9gc/TefPHfwVLcPtM0D1g4cG/V3fOULDz8KqS96uM1CmAcvIpzk5j4Tdh0tJXOWdVP
hXatntZvGzD6PqAMhitPAGA9dzs1lGzeiy/y+CPtO/UOrMYl+uwoJGvJFP/7jpsIVDdX3mK+yVvU
EcYLHOfRrJWcAZ3yZwnIAug2kXiI6CygFIX8uxsY+8zbgnPQlQG58H2mEzn657Qq4i3W3jK8/AvT
F+Q3q1eFVMq0CkaWtsf1p9NAbGYRm+mZZsWcn93tFpahcn/l1UN0LuyOPYi8Y+JOwjjIIEDRRwRH
42gaW+lj2lLrx61zwcwvhqHwXKxs+tf/yTsTh/hMjTk+4UlHzUiOJSkQhK8HbEsisl9nFzptXaxt
q+Q9J0wHNiGUnripnz/O907fipsL2rvXQCfODF2ANM99qPCxE0NVUga9WTXsrKlF12BRaweYgkx5
KMetj38TwSZEVqT2hxcDXNc6/2ZeY/UepBrsVcRBrsL+DdQ7JrmWUNKifDN1P8H/5rqK/CFz4grc
qZbp9dLya1YcA8cGvfHb9vyy6xKGRe3ogaV+0Fxwcg4yqzDFyurA+OuUYIZbI2ugJq8kzKS2euyb
PcQLc7TWNTRgoBNawBG51aZnkorqE20iRgl7abj17HepGbQavfMtgiu/JJeit8T8NjxoTc4/V6tR
u2ibX5Ay7jxVrmyJelDYFK+8EviUaaQMkCnwVnfNkuGGDudb9HuwXn1IrhDBKRIWQ06LOIY20oBW
ycJ9PFk7iIJzqhwm7SgkLq/NstuTC6Se+x9ZTyZSeVg8cmJd92CWO8fuv0Em1+Vjufs+i+Var+ok
BA2pifxKkYWfwg+lytObrvWAuddeDXtqPfENbjQkgnzTMkAwndTiQIxY2EnEFcnPmQ/up35xU9Tx
PwsyS+9P+6CEKAjKrZfzURn6IgimWSEWqezuMtK/BJ+9b+ws5UtMRxCzuEjkjSAwHHEDfqh6mC90
Mmaj4g1Tpii8TkgkoZo1HDbQrN5bZ0nqt8f/tr63cg/D9KkzdiXwhR9vrZKEDuIpX5FChnwNUUYm
bcjtsZW2hkFs0Y6jx5xQYo+3v/vSh3Xq74oW8rRgUa+HoszqI/VMI2JPcUSE4u35hYMt5yfgo8eb
zEhz3F3fFnp8lXqF3iZDG3vyU/AkZJWl/0KbXG3M9aJJdXvQZEvs1D+/WQLnya4uP3JDm8rVOlg+
z/gwd0XxR6SlvubZOHgifeGEdqVJijCxUiPT/PuJEsfsJLAQf2PgPyHP818dTc2Po/QZ7W1gAPHq
CFq9E/G+0lRpB19fVKcqdWkof3AgCBy7INlVNw5aXn9gicHF565nuxVT4nQrjgLJEuocRHARX1dX
vYTsG1U9GY3v/oqd+HHREiHo4iJRVnz7sZ9ZRsJPr+iZ25MxvXmk9PxX2sqAzULx6hEhsjrk7bI7
+RMqdxzlnDLYOG5yiSpDFT+hsXAN1QFoaPBA4jVb1XQXIULkgAhd6GqtMnjXhYZYFhiVzhVavuWI
/joQnettyn8XNHiwHs1iPtxCcKNt2djTjCSS+Gm+I1JwCuXBP+vz9CoDxtqkJmIP8iLtEYiSQC/Q
1SG9907Hu2qYDiwqXwSZZrIS7wpuaA4IKY5sFvlGSJLTcBOwhPBQ+dXoZx6kZ7esEdbTxVh7DyFQ
G5aJMCNeDttNOcwUXvhPHy5CNaMRoTt2nFzG4Bt2OutkHr5CJpNSb7i5PEDC79eYjsIoQ72rKxau
eohqNhYbu9vK26jwNdW/E7MPjrd+7j3YBQmZr6laJXY1NlK9GMe/XdGcOfWjEM4bqcXdsw+wF65k
EeOz0KvAMQhiuwbF1EFVnjX22mjljlyXy4H0q3Of6yLuL3ihI9LiAlLSOXDrejIQUEEDcWzZupcv
DxJ3TE9UYm67GuTUkkM13F6T/8W+nG0QsOgJm82ZpBTR7CPzHOjqTYC4vmvrkl17xYmn8yn0Bw5w
u5jk0dKTfwVpNa52ndyyD5TZqXeEeqh3zrFX2mZn9YxZZn4sJBu5lEZ226Sk4uNRPOx6eZ576njF
DWKbvhhfHsKnjJ18yBKobIezF+ceJwXZNCEymPei/PR1ZYsJHmcY64OF61nzPyCFuxwy+8dfPGhd
fR95cvLjjMU283JRIQlrHayb2swdFiOs1HPyusgzZ6oOBvKvGlDNk4a7YPXvkwsw2CsB4IA+Ic6D
5fQL4nDZp0ve3MyzggNEJIvHTxS8ztpZ61Vp6cPdTkZ2vqtycrlFoUxJ2cPn80wr211LmIzZoSNa
ee3/4UFE2i08yE4Bh4U+E8KGdk4vOSJ0+lnrZSDnQtRFWZYgFJiETgvMJkd1G37p6gm/XgGA+p2a
/kWMOi8hPoCJXmlQBn875sgM6pHa+lPx6WC2oGbDD07sI42Zyq6NkCGWbHdBKkX8gZ826QGjOSE3
4XtOr2nvabtaJSdDjg9+O/9Z+FMrhr+DA5bWQZiZcG8QfDYNpBKC9y6aY9JW2qCXZoMrKBnC8Eqc
YXyiNaRSp8Xc4g5U9ntUUx5k4K0RywpW06RWVW7o5sln7/dN25/EjjVYG+3McZdIu/64yqHToXxE
OuyCNWHkDAOiHj0cj8dEnnyaZ3uMKHYAkrZolPCu29648TCxWxa1Ct6t6NC0gcmggLDtCtfk3Yyk
RGoTeNy8UKVpLNVWSLkPytf3Cvy6gAcBWe7SPYNnbHUwt83nassI7DvKmOsGN3u7R21qiMjlHmGe
gga+2Z6YuUVmV9H110Jf0pNB9q8W1/d9zNp4OMcFH53K4CCyYhwNv/gAOdiAJSQpMFGn03s8wVd2
Z6c+pl8tlV/o340zVZ3q9TtFti84rzHt1Buu7B4G3/B3mYUecVI7b274CVyYt9MkEOc3n1T13TDk
cX4OpCTcJ3z2cquwN0eIJGgP5woRfA3umlWNy92nlhvwd1Wb/IxZA6LBrPW2lBbzi3nfCVcfUM3/
MX5kymcVYOby2hWrVpcAmWXYWy7KMxReeILe/W+AEjWxUicRZdL3bB0uPA0fCXhaw1n0RvKgP/S4
qOZqINoj1dDuHM18IP0m28OQ8uU3hhfrf+AQnBDdS6sWuSF69AsolG+YUhIF2zCtwo1LmrRUg2cv
CqB2ZkZ58zRMZOur+IWIswHmk+mPMHhX7VYcCKK0NxrxvsCO8j3mA0Lc/z8qHvALuUCIJLFRUKsc
m5yjCZQnyMBZEwEp2Eyxd/DmR2/60SOc/14uQ9mqv+dLlXHtEq0iHRiTI3g5oXUU14BZgfCBMGbB
4FVYXmoi5yt7djHfZXz/8aosYXDlg7mReZvZaPbY5art9DaGp4EdlLSX4tKcw++T/vga44fiUUSt
QkRGHxW4k7pLySyR4wpc9WgiZx81JNJWXcYj1ZwiTrR0V+rodcGEz9d/j8fJhVR9L/GrNyPCzQg9
WHzZcnLQVae+kkdVwxOE85W3JyhLQZl/lvqUrnague7ykxByxO9zztDi6gGjfPGVeLr5Jv411G47
HqrtNyVdcGT6rBZUr70F89n+YyERbxl/r0lvcW28///dXBeHdHpceHYi6ouuCFuXgNsC+cB/Zxur
0PGAAlNL6y9gGGbHAjfA/x69SRcAFcVGDs3012+maEeLbnccKmkzzr9wKEwDnZyHK/JlzWxz5SsO
2EnsG9beCkSpw4TES70QNkj6pfyAU8Vh/iO6av1Mcdp02D7C01Da/JcFYCBSAbFNSRi7Ndi+Em3l
DSyAsfHIC/RhnEUeLCIPGez46HZjcXx45OoifJjpLq5RW7ZcnFhK+zst8CMHj3sP3zHnh5EncQ3k
ZxHXcEMTtqbYNUL7QhCPmvimXVrydXe3JL5/lLGhya1pIlP2snWLLV/CFbljeKTQcT9BuBcS/F8Y
gErJt6fu85OCYXOY1SvyB+TS0vt6KU6n2p7RtSVDUSMrQRxR2e++cx4iIAw9eiRYyCbjXXmi6i7W
/SaMzMmt/Y2Eamlr7Q5hQDoRUzBN6vMCYzGprSLhIJ3EeI7xKaD0mQzkfbHAi5Bc0jJNuCqAKJyM
XIgfH54EYqXM+lEhwrtm3ypRuHbW10Exeu0llLCzKGyVJg0hn3Blbne6I3VP7dkDk0pLBI+urrLW
sipzBavnvKF0eyfvlqo3lqvjI6/23X/UBnOqwR4TG0PdPBHvGbYLP8/16Lm0LBQuMEt6Eo5X6Ile
CbgWMpIQTdUKsjOe+Xn+c5oKXDgc0E2YoupIpCGXbGiqd21VcWRQNzpVTpcsEMMgPYOw7hluvmZG
C86P42Saxdzc6hEZre4e57RvGrw1qj02ijRQn363IOulpPkmRDrbbB463lmdbFwxF+J0ndSw2bcE
3/hW5Yn+Czq4nimR6Rg8fYsIagEy/PlcgeSCQKtYbe4RNIAR51fyAe2P7S+GpEV8imrkaN3z1Tdv
UTWkrNHR1Jv3dxXOkIcsE1YUnX4tZne4/1olxq3qu6mBmqdsFcq6E/9MZcjdcR8hU4PW/KoraI1s
f0H1N+VwUnhZSkMvRSjPYp0ALBqapMK7sxzeFdjXngtAFWjCV8VAuezngDdro/gNrd4Wjn1qrjE+
Kheg/FxtqvzslafAdBa3+3sfyQNxjVqNEG/Gl9TIAKkQxdOxootn+l0MKqTsA1gIJMXZZ+OGU1dI
F2EG6cV9bJIXREPefqR5pQTaTmweX6Gbllde56t5WxEOX3No+RcYmEt4HdYIXSs+IHHWyq3B7Kvu
jNYfhnOanJE6VmpSk+UgMOJZv24zc8eoTsDXq69Q/ZOW9uaCELiJj5mXES71vRZ7JCHd+y6qHzRn
Yzrp9gy99DZFuGUm6FhrRUIBM629Sr8xEaJBN5jEMDHOn5H/pIK4gQbBuVjHr/uexjbl1yKUdkKF
Tv955AqYb14Utf5+yRDzrOPRaMp08vny0TwpG5KMEoDxGOCE1D8w8yQLrkbDWBOPDxu0Tf1wRoWy
bo8u0EBRsL0Aa+jL0Hi+/uVcMAn3JdV6nGSnVIdUh33kfe/ItOagvkSYlCC1wjMnZ6orXzgtegKC
UiMZ3GBKMBkV38y5rgt226sEdMzJna2RH3Tu9SlXvTX2NMbAXR0gQ1XMh4QyAJ7H9Lg036HbzPRi
kN+RR1BSoeHbKkYDgVjsoZDFEXMKBh8/rOuGY2nvDpIRpzWhwTgA+vDMYNc+Hb42fAtOQrHPKpVq
uBvDlsASxBZ/fTiQRv5BDJsVordcjbAi2UD0evQp30gwaXqg2HECp4t89YJgfeBrAKbgqTBeUQnS
3BxCtUDGtO5FT451DX4YfiQqckjpAHmDATppwOJ+plK4w3h83mPeBmfKUrqg2rlKimb0wdSdfm7r
3ddnAJk1NsVjvx2cardrHrkqIKB2jiHvwyUCNM3PT8+vS21tRKnEB2RWJCOM77sz+I0JeYThGbzI
3Jyvw0TOPIQtANRV1On9f4q40G61wzgJTMhs7gp74lrsvII0DkoV9jXX8oSLSQN9I9u8TYZwprbv
R5u6De96smt1Toh43ZKCbyc+yU96cL2HbAyv81oKACMwMqwHBiMZ8FtcCteXsZwI8er3CNxut4vW
1zGvU+xgpi52KSv+I98uU093M1TOFrDjTV1qOfaaa4qFng42RlxJKTiQVvFitbzyJVOxngcwuf7R
6G1+Cq6pwnV8vUXxPW92ohaR7jzXInkc1XSBOZ2ZP3lGQ+dvP68Org6bk1o09X0YrTd8bdY9mmlh
E7tSvGkZYMVk3I/Vcl5pOAHZXyIrZgLPHsa4YW3sAHaVUrW66ehr9K4IMru5GaHvOOkDz0t1hv2V
CowvvoFC6wHzQWo4/srQWzBs0pib+AldVhJzJ6ARGYqjJuZLnT1tQvn53Q0FeINIi/JE8q6QpH0r
6Em+madfPyCAZxnPHDTNNr01jKDiFP7HcsC6HG0dmSxq6j0Bzx1ywdQ+QfVsfBxdhnwsAgyNJ/ht
Hxj4auSWZZPv9KDb8rjNtdH4L29TuYG/IuX6qehhJCfSM7PRR2eZs1BTkcObeHh7dX6PfqyrqJOM
V4qvUEioU0xMVaXqDOZMY8TwPWD1jLfwdZyRdgJBtvoAHIJ9XfTN2U1rlkQrIm7BzAgVgoKVwOY9
bW0/i5IV7PMWpGdJSiau2kaqX1uKhXpzMHiUvn6BpeTXJGCSi4t2PzfPRRBt9fzKj6rhd0i935R1
9S1tg3A1/BfRABIAymrmaWfM1JIzERK5glkHXdDQSe5gaHTTm9FLcivN/o/Yappft0C8tPoXgQPl
Q4FUdDOrcWRaiVCQm4sdh2xIpGU3epLAx5CNj+PvsRKGOTXOizfIHp2VwCMGCxxvdLpZrMjmIL1e
Rot3eV2bhV8OsYfsA0YdTJyZBOL+m2g5c11xD0mPWL7F/i2ts2HpA1VLIWUUYfwCRfBiODqQ4Inp
J7SGOorWDlcW3QltDTdedVEAu6nlx5vUJCry6iw0UILVD3ZxsGkHtN+KHsHoYZEvisQpl8GZKhRY
j/MK7X70nDWlZmbk5dA739j2qgo/kwB+zX3sFMc5N2Ei0aoVNOPrpqXopq01AsWJutcQFx9ZbcJF
3n0Svyi4xHXzJWSM6nipD3rSSU4VgPmtD6mVXG7e7zMij2rWtggjQFTvl+1moOB8FZKcx545dWn1
+JLlg59yN13kcAChE8+it/7mAIio8BOuCi0KyZTHp4TWtpfba98T7WF5R0Lk6X7w4yi9SEPckqLy
9hLfT5BGs6wL1w61+Y961hvIqz8xKJ3ajPmULa1wcz8REk50bzn9FLYJpIv2E6Qjf5pqr+iVebnM
mWLZ2ft4EX7S/Pni62Nvo62h4B/VEx/9NWan3dOW5Md6I8b/Lx6beABM9FneKyNcR38+wl6Q6YUV
wHkoiY3+Usju0xxQ13WSq55GIKT7OYwwpFqXhO7qT4vg7A35LU9oWGz2oGtKjJKyC+sm90KG6UHe
wmfXFdWMHIrzfaRzQTsh4rULxFVBY61rnVVq3kHHFDoE/dx7MMpgt3/k9fHspkBBajqEHHhtS1na
qduIfHaZc5W/8ahEhzklJyRQlCoYLUc9LsIqYT0xpSOnGz/2Bsm1UR7O1zQstFk3l8oTuQhDcv2V
JOBobCaGbHlp3ymhinabOQptyb40Rr/tx9xTDwrQnEgInfSdZ9pD8oj8gvYgkxmb9Rc7N3WZcMeo
BwWSBWBZHqxQzDCvOywmtQ/FgthMOHLXuA2EK42Yf8wFMUnrqNO6zSguPCEturUgHegucfokH34z
N3cGSXCMtKNDuzxVISMMDkTcq3NzsjaIXQwYyC72mxLSaB/yLJYU/PkfM7iITiC6NDcc8FV2vusm
HigDmjWVFw+nj4psh7241h1iEzXRa5RdpSy+vY/E1to9lN0EwYtpGZOZWLEHPah6XZuZiTOotkYU
GUxI7MDpT5e/X4HLpBh/UIrJ/23ywj60rOwz73SPPFq3LhIXlJmZ1VpwVdNjN5AtUuk53GYF7l8F
V6UPBUvlzODXvIqy6RiqS/MOa6Pkg2O/keXpvrhytHZnZfqHOikomirieJzoaX8BJ+DeqZscgxcO
OvGrLoehwheS5Ke8Kz3GQ/gJDABbFiGcRFE5f1WGMCzlH1QMtK41lOHUxSe8l/fHD7zYZUxBiE4m
8qbuMFimTrrpA0Fb3CfDbopHBUWfPe36st5Xt4v3nbv9rXmSjBwqgEIPpgSFkv+bQqiR3VMbVC+u
yTd+dKTD7zL7qIunWzqiHzLdl+LOI668QtZ6GPb4obn/digZe/fC0ncSqfyyQmCMAVwHD6xEHAMr
4LXaTNdWP5ioPAeWnTc/MZMQPRx/RTdam05BCLcVhHQYuBRCsptPn5uctMd9aWXsBBCxTVkD60Xu
vqkGnX/MxvjA9uGjmsLczcnRsf5Z0qvDn9BB64uAtaPH7q+1TmHXK5U8jA+C1shuitTA6YxsorOH
/HO8Af+ETBx4aNOdkV2o1Xj7LH6DfYVMZMA/sxXKfIqhj/J5R75NbP67/Fsk080dbZ6IuMguhZLT
eIRBBwCOUk/PtKV243HJzHqMqngylNrvvLvDBz5y5kqRlD8iIfH7d1xheqUKqmJzZnQUw8WE3mss
JvyEGEuF60J7Py4TaAgWFq9CEzmaWkSKSQmHovnCUm5uao0ib40gf6/M7K71NfvXyZ0Ruu4DHB1O
ovf/4gPPcRb9L1QbZ/Yah5vtxCvMjsvEtWiDDE2HtWL+66KhJfRgeUN4FkTZjlOy1y9yo1OKQeSq
o0veWDMVa7s6sX6awannwKtma9B1/EVzpMklXEFh1K95SB/ZpntI62FA6vib9pLihjNXMVo+DT/y
ljwxgFiV/RRsHrDvVuTm17wunMdHnngLqCDW5XLYH9End3WgL9C+wrzaan/gfmba+oGQ835tLOK4
rJG4NUj5KA2oFiDdV0az83ax9/v1EHrIFhW3myaT2BEfhWNDwCOnQKvb5EJ4j4esT12BykELW3as
K2tBtKPEF8EekbyekWFOSUXS5NTMBIOrsGm21JogWb826IzSiuLMjhOSQpUDy0dWBAahQYfy50mx
j7X+VW5mcog1Cd9R+FVykksAAfopo23Q4xXLefigZ5d0D0MkjUCjzgY73/0TJlDhPbkm3TzyFdoU
+FCYyan90PbOMJm74pla5+HgKVNbN4jh0sXJaQjJRKRlQbtt8gSMDME2dGHWfuQsHtdqrzYIRvpK
XlZx7rizh2Uj1+CKV5jAejK9NlXt9cTOpRRG3RPl/8S8yCPsMPPit2FC0b/eMUyqfdGtYnMY/OFS
th6tAUuFrPEfHexx1dkWJ3gbLFUGPcH/xe2R0Kf3WZR2Xmqb0Evff/M5O0abo+z/U67QRdBu3Neu
5svOXmOUzkXXdZmaJUD2lHBVuJGrlwF38BIzxo4iO3kX9PqIh6v7MuNspb6mCovNhbNDeZFYFm/4
4MAcrjCKN8OjGyrAHPp5rKD2o5x7lhy38IpjlbH0SBBl+WqIyPPEaKR2ZbRcOuacyQ6SyjB/2UhK
ikxnAEzgS4vrcfDtSS6D2lfn7TJlzN8p5Ubu8078vpZFNicDeq0pIxM/HEXscw7TmSn3h8qV9d9N
OY/mmbuENZm9VaLg9JpamIHo7JWg3ZOMo/h8RNgui0+C2xgPDSvg19hviT7Gn0RXSFqUbH8LDDpc
KqGUUvDijf4maxL8GNoA3xhjweJlwfncUnSx/ITkhhDiqteuq21NQUGbc95Eme2eUHtFScy4sGbK
4HJ4EIvfgq4eeDMxf4EssLWL0Kl6xtChWZV6nmIlCYZgW1IpXiS2LLPVAlcRHapE49f5iMy8H/Qb
vxvCuEo1CCSUhUMumqcZZJoIMTDvI5VNFim+4r7FTJ6xVR3SHHJp3/qbuwZJUA2ZycG6S/0n6Ucf
8QX3tyoX5eJvb5aHLsnCNMowrdGiKUwETuwCT+YA2fn6yEyKoKF+rf98V6qdY2QWd6G7BX0zwT09
EDcsTf6JG38MVflW/oTFyCKToYHWt1nBmCIeI7dmEY+b4Du5bARaLNsSfFx6OQgoqiZCUG3c42Hh
xeeKUS5fxVaOoVxmqsTCIwQdNSHtG11oXQ77/2sAGMnjFjcaOdcIY3D98PWsgMBgJT4mNDTroCR9
lZ0VRZmWOMqhACxOWUf0wzOg718v6YVu4sfDig6AQp9SZLCO64zu1Gc52YNMMktNozJHwJmtfp5S
rjkul/MEWisdIUUd10FHLiNbYCAI91fYC/+7OBAvRIWRzWY7B72pppp2SyvvreFNbPJdZZeCRSpd
aQb9MaX9J/2buxr3x2iewfuFGHiqD+gN1x5OhNYoZlhXe69alS+5O6gSj0LPGg1hb9CngJnr1Vtc
6k6JCM8/mWBGHsk3iST9a3OuBrUKdjXfR6EJjhzAeRDy2s9WUYmeOAWxAsmypK7qzn5qD0bKO2xs
kw6eoYiT/qiZmRwuTlgKnZLnSHn7fJQ5XjOYjLbZ7Y8ssKG7NZGBXjHtuBA4Vqi5Uj5KHUG4D5Sh
ai+6VPnH4InGkxLkPN87PaLdS2UfqGtuBLM6artuo4kRzkUEGiy5MhEYiUTf3oJYybd4Ln1tTcjB
fQscghIru/iAnlS2qlITsDABUW8OKpogUyYGe/OCT3iw1YKrwKi2Ykm/EpXaNabjjTujJdrf+6mA
tXD+eHt2ynniVC10OsFRPGI8SD/ag3uPVYEqeTLgL9H/oGhnfzDjpQtaEXFXHUhlzWcKTaSP4vfL
IFrZREHTxUUEeiaumbyNBEchmbGcLzN2hoWFNEDJcJDaXvLnvdKSDrjkoR8YjTwFJYNGiPraSZ32
TskIg6R5z7EfHw1ilwT+k/kkeOmpPnyacfq7OVFEl6WMxZLR/rhdiw0Dz4jiST2WriyAr6otczfM
ul1xGq+u3Q4dMzl6eUIxafVv0q4nnQ8aiBcTpIlQiqE15DZXoh+LFnH5H9kjDqn7o001hS+wjj14
2o2sOtEPGBVcPlWySdVOx0Pou+L2ouT37PceVI+Y7W7rKJbQmxaHvgGiDbam8L8NCJvBb9I461Gr
YW7OV53WVh+90K8Eu69ZHpMPTUEMX6lEv+xdEiLb+wVQ/bvs7pASNw1eFZ4MeGJaQyt2qD9sKotw
vHU5fAFy1KB6sexBvfyqDyUwpDAj65fUJ+mQZJTjYDs0mFp6/n/FsxdWkrYImhPCHvZGNMBwkEwp
1yWjkeG2RLWABj0siDuynrTXh51MwdQNIvnCzXi6ZHxoylm7Ldhd4ki9Gbp1YOtUpsjkwgS/e8sC
M0QfZ3hk3buQQ0OB+lZugDNu3LcdjVmbRN9gogTEtk9wSUORhVNoy0E5DrNkMRZgOcvSUb11oRP1
xcTMgW3+K3No2IcihEY0u3pEqyH3AouopcdfFULr4EUprmVthPQlP8NvIBQs0gdjowkn1WvBcThU
CUsD4+4tO3LOLJIDvABtia0fuIuP/58XTrpsihsUexPghmuda/aKrfuenadZ+zc31r0S7Ilr6uFh
808S2tEPyAvnxmd2Mw3Eo/Uol8YiiZGt69RBTE3q08WFyYvdcqOsLXvDft8K15vl1EgPIOqyG12m
qxgJNPjNyueHp31f1e0iaEsUgxgmsQbm/TV67BDzzJHzou7L5Q3uWpc11GAOSqXbFlnHF6MtnQSQ
J65vFB3KFpjjUFAaOJVO7eIrzUSG3S+Ys2dqyuw8Bxcd1QH/Y0QCEoVHCP63LcYylMJoCY9b+Rfv
mz6OQLzQm8Tw5DR8awd7vX0fCFRDMkf6QntKnZdJ6GFKSqI0gAvn9/ZB3rbH8+NhJQHANEeiYm8Z
ZQlNlQTsPEnI0t2hNBVjPK94R8Rqzx/s5egscinToqhukCU9V9Nfs1WAwSZx1croQaFyz890U/xm
XibnHx5w/ZIGSI98/m/VsREW2ksJvgNgRF7/UngasJshwJxMJxELsOzs98iE0Pde1G1Ld4Tv3dGI
kam+NC4Z9JoZbKAIJQZSpJhr3VhEgc3dxNmPUD0EdJsvHvPymsc89GabIzjUwPcR/qK3qnmZiGty
Ls1XZET66nzxTPyIHYPBnUscFbJ+ojl3bcP5hYi5X3nkJvcNGc+06/TiWews2T74bXeXL/tDozZS
1R0AJOQjU6mp6nbG4OIYYS2UGwgQgxf8y3BnKdkH5YjOGgN+4TA3QSUi+PIqDmTJCH8EcXdkns1L
aOqW5BsnFq+DTzwPbg91Kpo0wCwhdd0SnulpXpowVpdkuY7Ol2FKZGQ8+idKByZq3x6xy+1SNXKN
uEhagfpaFUZ9CdpKgPCjY9ANpDD755aj5F4QJePUFqgfEcSMLVDEUHFskQHBCceDjToWklKUW6r4
P0uct5ZOokQkbnHCAfJS0IuSuGQozLt6jvJlWNZDQK96yOwPJe61WMyJQRuqRLHHhdjtvloYul9G
uAeh0Ibt8gnQKn4VGPjTPDS7yzRycllAKwYOayYBGX56wBCfsmbUNsuxOvzjQg8S8YwbiioqO81D
zivi+7WiJ+Jz2s41Qt9ZtMyiopDYiGZ0ryWoWlzWLRDiPehaTl7aN0/4qEZwEQZ2JQcVaM1apkI8
R0f8sdId/191B2hfVlSM8mWV2709ij9w2t7U/nPU5EALcCffSMy5EqTjFLEve7fuWd6LntJ/SBnj
Yw3IkJe2fC05oT2yXG6REjrHE0GRkEaswylvO+6ajW+HpUTBo2lsbG21UuKq7Msm/l0aOPYf5g/L
Hz6J7wUmZG7RxD7DjvP/nKBDhpJSOtUaSobMYWkHYZx6mbworKFu/AqDsDp0pTm2c3B/YWYl0kLo
HdQA7d4JrwWwd3owHOjGfX2WlxAyheuPzM70VRYvlLu10W6evmmISwGp0ZPmGpkxE9nRkeEgUcNW
1c5mPzw3smnnWhM2Ce1AMdMlA68woMxXKYJuqx9yv4yktbTLlw9jcJ9NFndRFBcuTBtNbJdi6bfw
43eKj2HVRdhT1p7vpoMiE5lghMr22jU5H8QhMQP1RhAksvA6jWS3F6lMltQTjiOXZWUugSAN2pU4
Gh/0VVlS3Gr2x7louwgDttnn0PXXNMcF7YoHhqafZvtuzCjU9HfuiHAHxHN8UBLG20tx7qX18jiy
ymoho9fRyzt/je2Z9saKtpA8iBfIPuRqbQow+H0pZOB/5tArBQIaXHucwjr6P38MT6KmKv4mEwgl
4xrcGa9qEDOpWFAEVAKd3tIiqFUHAijVMWBrWzaZNQxaP+8AmizRnNekYLMuW46pFRYzz67IH/lN
n3stoCW1C1V+laOCQUyVDTPWrhkCs7XE5eGpL+eUbnCWzuhfZWPC7KMqb4E0jWCjtKDfNb8DIIjY
srREdLQMLMqTHdgkqSNQQstjy50vM24IfXqaUrkpvsQgZXr6n4BSr5WnSgA8oqUC+QvObtMXuFlk
5VPPNX5vjJT2biCp35aUlqDHjPX3EvdXTi4oQ3Ce6tSwHT2BulrrMqhx1uABT7fyhyeixCKuWtzm
+PVJdZZLUnzBiaTHcSUqWKAg779TngdCjX3MM+2SUtPzuuqOfiyNKqMHdsqX6M3uucPdd4uaVZ7m
sOHOFmWnucwExotYDWtiiJ3SJ8s85H6QGOrtsGGvAaB9qsUIgsIRoWOq/4AH8Nj8xwtVONTFuRSm
emmD7Cm4SkFuSHDHQgQAJ+6NteqQVGBF6d4MG88YFJmySBKYHDr5qBFmfHdItY7YyuY1y6obWFUy
IgsQm4NuyW7kSATJcTVjNVZOXBevcchY00ksxRIHwjdcRMivGHD4lriuL5UQgac0BborGXgUBCbC
N3hUkcVMbryCFs6HkfvmcunYu/TW1DOWpY2006rDrWzcy1sw5jnQVPLnyxdpOrweLxrE731rDlij
FK/x3pCeCl8G8WDIlbgi3L36eeHvyj9Sjkcmd9JhXNKjxZ3Iuu12UHqcjyjAnKPLFBkCDLskUtFI
DSHTVmyTg69wgz+aXu7+TbS/k1bcv+S2dsxoDLxdLN9M0+0Ky/nhG9o1Wi5Rtj3plVK8NuN06aQ7
yry+Rpj7tEGeRSUlOd9OSwi9fLrvSQIGmVVeWafWWooZEAAsPq6RJYcu8JseVxGyjzcyyInBOsqR
p/V4qRzR8t4U8l9w3XzJ2gFx4G5tlysuRATDvnMf1qAJtmBqDPqDozU9QY7IDausNDKE9qpvDy+v
9vnfzKAQHEq6JOhhfYP4TEsbOSAOhLUcbSmcv8LMKsruBXLjmH9qY7oJunGB9+FyXd43sAfNL0l2
A7GfMa1+E058cV2+ocgr4hUiCLCpvc6p9AHgQz3tn/xVSq/+Tx/QEyNZVEWvYBKo2HlaJg5WuS/6
TuEZue64o32LZ96atayahe079TBTXPzH9FvwQcK8aFztyvuNhXS6cb1lnNEdTnmMJhpf0qQ+nUIJ
frpikTMDInUL6yoYUF4S+zhRs5njN+CAwMafYRjmy7iDRPqN9HdUbMAmYpOvOs/5uyWcnG1pFwRi
6D0XXdvFKirmL253eVpiEKpbV7PXuZ81hyufNJfpghZN+Rnbe5NlW0H2Jv8WfzxRHnoG7KYk7qrQ
yPgG4Baa5nBkuYRF2qUNFlNoZUURLqDt5YzKl8XKMa4GItzWrR1Fj0uqxIM/of5T6Fi2RhZNja/x
aWr/GTmc0SBV0k3zKHvoo6K6NNyPD90JrS7gCVzaoCpU8eYs3B7bdz/X85ZEsevzldxpttNU5WLy
lbR4EvCrlfJ46d0tD3NHOY2skUbWFWqeFU5vC5kI4CoQxTcK/bz8crhSbRW2czYzpFkZKM2dTfCM
MvZ5TasKepw8fHoaKyf6TMJt0A7PP/sRTLX/ULzHKGUI0TyPIMO0cz4E9KRPGiTLQa/DVEX7kKqK
KWT+U1lYDf0wFyACYvK9BwScgqiqMybBCYwOmIa2vl+0o3cc0QGWoPcXzV3Xxw2aAya7eUntmEM/
Vzw/utPZMr5jwmxVPF02eJww1mET/TNOT9WY1yky7f46tcKw6JqJa7ObG/aS8B31wwJHATfeBPES
YLHFvTIchXf9ienNGGM2/41WIiwyd4ReGTM6fR4KCJyp350k056dy/3voKeHwvmcumudllTOwGKi
/A+QDBykjm+5qS+TAR8StDZE5Zd91bQKb6y0oEaRcVqyVZsRiD/J4LmXxLOIgOaTgeDbK3BQio5+
Pf/xLP3KMH7zvKxd2mV7BYGBLAaOeGysP0pMzwm62fDaQaI3ZLbPgZLpYY9UcJA76z1q9wYIs9Ze
RFuMlNApBa+z5VQtWP7zpjF7kCI6m4o3XC+WCfDi2r8M6vBm20vvYMqDDMO1heJzda4AqOroSX/R
Q7mFMIYOtRUZ52UwAxnDB0gkk5gZK/7n1S3jbVTs2vPAG1ZIP3kXVVKFQhtDzfBz4FhBFmRDwhse
HcNUkf1KBZB4OZQ3wElC9F5clLLg6AC8EBPKm2In7W7VDE+1olSVWar5vbHgRjLBS25YmGEmfNAY
6zvhbFa13pkStmkq0Jbgu/9kG+fUvY4FOVnS2voGbFHk62BwWnE4yJu1psVUoeW42DNmypP5KpJC
6jjIyOYp5jr2O83uuc+49oP54svgfWFmEmYFX6NzwTLOau+e4XgbHbbc57DUT/odTPljoYkBEDUi
4NvAy3yERq7Gdp7uWYpxokDYRJe+MlIATH3doQoEvy13g/2bUGd1EY3k0MS/9hd2GeIBqM3Ldtdb
akXLW636tusgYMZYc2+sTxo4jDXaW/cOQ1H6abAHWcszV2LJhGcCF2TkcfFBqWriGtTkiAqR0QMj
OHi86iJf9misDhMrWtfQrWFqRQys6dwhP66zrpqk3QcoaH9dGQXL41yZuozH7+pXAlLZx9iBn6I2
Fu9k5GRA7+mIKa5wuLYHOXsY7GRn3ofRf6CzA6Wd3B+1coh8COUwDwtm9qUP2HAcxa9T/6u52T8t
0GVP939aQ14WY0tjP6PWKOUWbfSXBDCzxctHS9uwrw+EkupYpDHLgelb5BOniY0NAQh3hQQIkLub
3qxAxmfLRHe1TQrOoM5XfXGflcXBOKyC45Wv5Gvq2xMS2PZ5RWhbr3gDT2Len1jqoPYOWgRnn7Tf
P4WIH7AflirHg1/NVBRIi85HgNAzhFexUODcfbfaXkCNEskIjAM3JeHc3+geEGfcvffmsZsCTmDM
L1qeRyXaTJnTeMlaEg/1a0ynj+tZKLOa4r9py0xRa5Hk+tHcfsmi0WHN3kVPM4WWokl5ZRdGGE++
mw6Q3miCIJlpIMhZCz2ZTtp6geTrHv5DjrnGlZZ2ZD0Vs5lObzpjlB9d/QkoMsuDoEHAT1zdwtTg
44YBiky7S4KNaRSc7wDlDYhfmOCzfJRXhcH8ShxuJxMgePBt5oEz9VclxM0OqDPOrspRh4whYhHF
IviqMJbiynVnEkkRa3CiBtU1qL8eymm+HzfqNvS1+q7O/4gq3jmqqbLyF6+EcmQJfZbMtynFKkaF
rahKTG+3vuqPI06aKK0L6AOK0MslB+am+N1TjdBJbDvcIVyim0OR109odhDPUoRbl3VhiVvGKqUG
Sdkx4hnKma1RZC2eR4E6rmWOAeMCBwHuTGBfp1uYUFK16V+qQGtMoqe9jqcSPb/Kveo3kqEC0Q2H
OphAY2Uo/cM377C6bwrOxxebpUcwPkgt1ODKlV8ETZKm+TQqeiWSVex3JBoC0XOX1f+vUgZQFFVa
OXnmMI+wF1O9F9EIanL7L4FnRkaDh7NKQPfMx294CwLVplHBGqcQuhShrg91bPf0MWFwcqckFkv6
hDFe/qtbnZzADl7yk8BO80Ti5ufveFXBrJekkKDao5T+e5a2NQy1tbexHZrrIFCScdvF1FtMLyS5
QNtmvDWpU5PB+7C1pUk5TfpuJMGtd3QdhdgDf4xDoc5TFuCQrRK1Nfr4ZGoR/NTb9jCYozQ4W58e
5GMxCSdU1efvjNJF4ZQvdZqCvlpo5/B9sQxqHUvTWUQ/wW0VNklhUSqbq/fjg3e0LT72xScC1er5
o0DSb3mmJEWk/NEKbeoJgFBTjrFFUuTq9CYfDqzyQzwioUbkSPesRP3r0uzzK6WWFt8y6qgUNN54
sMWz5LwrKYz8qX5DTucPSR++wp5xzlXp2yMoAWo/T60owljeqTnltoPYESs7RYWYRdkpGlZC3d0m
uAkR8xH8PvSxZICi5fmxHe7cCh99jRMf+Dq8Qun14QC2ZhjaJTtfnqnM53CZptYnZMDHaBQ9K4ME
J6Hvo5SBC0bMbP3ouAQsomxZ7TFeGFc00yAoOvG2z5h0wCKf30Ifwfk0wYcZiWP1yapCWTRaYFGx
pNMY0OSrITdEu+LHliXkYEV2bujBCwYUdoME/OhigyH/bgw6U+mhf62YRbitiQ88XcHCQq0p4U5n
Q4XRXu8CWinyJ3WAKaSLoQmmcWdQxbN3a1sJZfP+1bXvOlo+2F2M+a27zib7UQEZrkXi2kPXGIRt
t3Hx/ZTx5t0COVpqqOgg9Nz+SEXa/Aro+An/kizejTO1XOuWv9RQ8OnH/ynsksfCM2SSTJS6EDMA
Y9X2/FGy8XOpWygWKP2SNFKl0GXjwbnl1I9pONgrQwErRPGloLH3V7Yy5M6E+q6joo0cjkr2Ucjm
vgCw3wf4gA01kub04Rw5t/lUA6jCB7VXUnTAxd+krza0iVNzYHVOjH4+85U9d6LE0jgk4YGTTK7t
LCSFg/q2c+HReEVYljhf2yEbluxGLV091xqz5f21z/XMARJErezIDleldpI82fZfe1lXbwbAGs4f
40HxkyPWz/P2tl1ryEhG7wEKYJOoHR3r3QpjWnX4V4l3kBY56jqlWm/KeoqNuRiWEljKIscR7Ltf
DNxFE6a/y5RjAnV+HRF0ZjZYC+tlTfzaZ8eLi6sy3ksGYbNLh1z2qfGpM5KbaJ1M+T1BeTZ1mP3S
KUoo8g3JaHN/4VCnQbLukl+r/Iv3X2nqYhuWp4QE+n27B88ixzli4/6lNgOGf5JSbJC5JbpiQOBx
y/1qSjlF5g3salCbzi/N48YsGnp8xHqOPQevixm6rbLUudLNG6xaSkGsIRa1ABvwqvW7KlDvpSmK
lkFhsSM6S3mhSvAca3nYgM9IjzPH/EEfvqS+YUsUkdP5GgHUlKdt9Iw06eE9qr/Iyn5JZQ5I3rxt
PWB1rv2vq290RhqQ30SQFkK9e/GAfVwdKsYnxpN1iSA5BHLycrapntPsdoyT99CpQIjIfQ/QJUSZ
om0+hQVpwrCBdbinCyS/1+/I0acfrLn6KmXvG2X5Wq7n7wYdc6HpuqcWmjhj8E0WY/0a7lcY2PpZ
iDSnDKXD6168xnz5Cdce7ZyNPK+NTGH7VVfz3GA2BLTcD9K3+++oGHH6VI+a/vUw6v2L0Ei1FPqH
7hyg+z9vZq5ACUSp9oam3rLx4hGChOv68eTicxoFeeDSMygpe92rdwK8bDTW7Hrtpp93U/R9zCtZ
qBduh1Yu516IWN6rjyuFC3gbhdfQ6slEbmz0I70jz4dcTYactsY8y0I1S5ZcRW4ciVSNsqh2rwDh
JLcm6vyxZDBY+edwoP4OsZKVI5FhcWBeiooF1d6c3Ch1aE+xxOrDaUavbntWd6IhgUZacYNTMZzY
l9vQo/85HRfvPGuTjwZkpjOlO/Z1+ahzJn1kYoAaE+dA6KVGcdDb0X3NRja3iGmE2x7nRgBRKc7g
tAp/pcrN286VKQB1sc0Nd+mxkG4WJMr+Txw70TjNE1JpcTsJ9Io3uHFmuqp34TvJS1knaq64n4pX
sPzg3b+dJzQtMzgBWRW15AtDiXa02mkd0SKTHVcVdNDfeUjSlv6S35btAS8pcCNZiUyBQPz/xJDP
otiQ9noYDDtYIuW1FvnKlwD+3Byj3Xi4OsWYphEKi6eg3Crc/aqTrxnRNjF/INEGcmpG67Rtpoh+
J2DSCRlXCzLt4zuN8up/Hknu4ReN0MF2Rivmjz5xsz70Zc+uUIgM0s1UZjazmQ5aztlOBBDzF18A
9OBQrYgAsAXy7avAXf35IDgjYjPi0ewqLN8O6uY4cdckf2ZpCKv6qVj4XWmmIGEykPY6R1/deYhU
91w8zairzA/xVU+O2d+U2+lLFwmRSYtFUYk60AyKHU3jmjVtpobfcB+KwDp1XgDSYvDZnaQ2VgFb
EnBkAIwkkuhgrDg49LZGu8nPSkdrM9xmpbNoXcBYJXDrCYyB3X5fWh+2YeTXbGPDNfDUcGSVvi0l
5NqdpJpcc1y1q5keE7OTaT3KoCN4q4EKBZZdkrpQq9xYDMORqvA11WiT1nAOp+eaTLZ5+mwnfvDM
iMBcjTve+wEYxsCtVELW6VrE5KbBzTM9rD1aC0PqasevgBEI8mx+Sp7mHM3VuDc5ZFB+ejp226PY
HUT2oqxqePmCyE9BTVL+TyatG7KItcljUH6HT8MYSKolnxGhR4dwBnj6fofpo/O/LTR+Rgb8dkA6
Fn6Rpfvz3ISvbBj54r4QuKAWf5phBIh0jZJV1H00OtIoEDxTbvTFcZF/FsY8M1Bngz/r5SJgLBz2
0UO9eRwSqPTkdri+sYUsGijmIqxFIYpd+AGzC0xADhUr1Yn8DvsIk815ZYhMJPP/HyC1LcAPge7+
lOI4AOVygDfWxHhMifdV611hSY4hczE0KheYpz8R0h7VZh86dtWn08P3Wds+xllnrKuNdAlOVba0
xHxNOxWV9NgeEXXj1vGTfyo+vxr4DkuktHMZtxCWLViXXKHzYkUP57kodIV+khsat/7x9Yrs5ueT
Zyb7EkNjwpmFzkWJji1UYbwCmmjDQth5scbYO2NbtMq2X+LgPX6TiUzJ9KpJ3NHo2sLbW9oi7GaV
96DpfPW7bXgbdbqce+PfjZr+4d8fkdiMH1OV1P8h1yAHWRmAOlzf9Z10lommXl+LovEq39b8BlQ+
xdws/rNydlb8uHZpytELudinmpFvANP6butyvY+iSnULBdNAD83ucM3hWzzQ/cYqtFKZaXq88+el
QBJPX4gtWfHATUL1dsiJ1Fm+o0tUgVDqcRltTp01A+iswhPSqb6AXaW1PAoX+VpUWM1gQqVZ4yvJ
Olmm78Ll/L92j1OeTa+OC1g6vj/PMWkFtyvKbGKhj6iVS0Shbxnk4aHBSiK2t9B/ZqjXyCBEFhiO
QwnSbDxgaG3IGjT/Bx4+s8EthY5AWDTvFMziVNNhmJzzuZEFVmX36iOOWY43+nywGis+bpc2Q6bs
NDQu+VVdTEutXMkf+2+b7RnClCxbu57/w/l4VlNcE7P5+x1f66RhV3V1nMUBcVWF3Ve4MzvNuyy5
Nfe4dkZPcIDEYYvJt4CEe+BkgF7R4iWtpc1jCIHG7fan/+C7INd24qXeLY0EQuXE3F0TQq3Q/ppr
4diUoYdespdJ1YgWVWYCRXLBxsxUn9VQrzc/oC6n5mzB3tpiNxdHBQKhahNl8XJvsZDKO5FoT1dP
8ZM35xGlclV8gbUnIXVZ0li+EwYjg/QCq0D2uDre1m00mN8mdkJH+IB2OrGmoekY9zsJ6+VjjECe
89WEbfLBYliV6fXf/gQ/fs+Ars2OtCbrIQJpBP1L8Fgo5l9MUDuuDFj5BEhYZ9W3CvJskp/zkKvI
kYrNtuVlyu93Is9k3aO+3ioD9ODVQmD+sInHCiIlz2mm5UE/LOlLX7awVcoGBiVEO02F6Hy1qUJ3
ylDBmijFcMlQniCrtUyBI6lD5JfXH3sQQ7ie+yz+Q4LQyDrfQuwXsia4scuHytT4C2KUyMvShQ23
x9T2EkxkjYsTIOvPYaxTFuBEzJKzu3wh3I3N5BgIBuWDzC90FgMkuT7poR3j56y2fve+lKUsKPlU
EDzU61Emx8Gqdw2I0m0muqLNiS0a2Dqs8Iy9UdizUHalCw/4FaMBXTiSppxNJHkU7QhQ4rdbCt+s
wbeOU7wfOiaGgI6P70br65Jp5JsKNo5wDELUSMKK0OVlPKe5YLwTwIiKNnDLlm+FaCPGha7oIzRc
KPL/1czKaiIOzrncs3Ms2fVRpkQOArykbdXQiE8DRX9lAfr45pTrTJW8CaOjFkT+xaaxz+9zQzle
R21AvnoVAI7gZ6kVcJf5asrc74tOjUDUJB/lRzcopWqCFYRfq4q7AG48hmjqGbPxESis5vODpH5c
AuhXwCg8DLPXGHzr+F6OWX7P9n9L/5XJjPfGRYKawQIVPpt+jrow98+AwtchUbJIZP72KziEa8b1
tCHjMkGdQb9M933+owIxhSjBdxxgiDQuULuViLtWaIMiONO/UPJaMigjgA52ujTA9XFu6DaPOv9f
7DYCoyEIdN20zPTHrh13FuzA0N8On3epKazmuqxP3W0mEvanPwwcXZqevoLheC/A6SpOJY1LiTri
IF44Ssuj7fhAwaLabHw+rsbeHr8G2fqTLPn0uMPv3PHU3rUF6VU2mkCABzwENQINLNIRKZSpUWGf
kFCR6mZBf6K+dgH3G05PXL8VQdwH8JpppzX5wx1iUR0T82BYfkpP/j3maPR+NcPzJ4OSo2XOroGO
yuJIw74YWaH+W2XnLABdVf0oI2pmsGlj19R8NvwnnSOgSDmtUwkADvs9ztWS9NUfN3dM6v+AgvBD
KrJAZjxD9W/P2jdXEp9ASUXFobSHXHCf8VwpU+6CJH1NjAv8ups0ZR5B2AHot2sdEbRELHanI7qu
IWZPVRNukRWvSYgFJY7EZOUzOjLAYqG4Nt2jwgzzDV9rvGb7LlOOJlpXe0ScKNbthCJdomsKn7pP
W2u9A3al4oDR+LTl2wdZdG9a9mc252W+eB2fRQR9VZJXpXNlcy044eEFYY8K3BvK5cuFW+6diVxq
wNvDpz3cdRf/E5pIlmnsc/3xzLsSsmjIspfJCq7K/+YH8Hqeb658PfHZjaUeiiuqlQN4JqnvQzRg
Z2ZIii0t6b7rnqkNFu6trMe2an73f+OoIh9VQiLSHtTgg9N219flcP4KbOoustx/blMOM9sKD/yH
NEYHYojbQty2gs9ahBXGwady3nXkaseWtETvz/t+1OjW07XC51o7RHiAbRKUrEpeHL34ErE9UooE
+cmAUr8hWKYMoCYRm07IybBGRV+0VeegPk/neyhUgwGmqWJYVFM4Qamn06PkeisbV7O2mutQxYkJ
548U998EZXwe2A8lCrMw4xTW1vdDriFRkHnjy0YTl63Vdps/0dkRaAgnMxIfwa4hCIBLffd5TI7b
NgbVB3rvaxE7lYCWMX31MrxOxp46VjB8Tni6Qba7fj6PI5GKZV9ZPgZ01U/z6a+/rscv5cK+qpJk
a5z9hMhXsKNnsGYYyOs+MNzO3YVOuGFUrAM0AIGHNoXhQbrM+2sHwZ4s9huPMaJCMUEaJaVvVX6W
MxEKP9/EZ9fZtNVJ3raz7sYTs8taQ5GCG45WyJ2F+A7TeQM2ltmSq4VQvi77mtSJf9s5u4Iurlg7
OzH5dJqQyjvUwRdfSCA543KXqoWS39/Yk+rPQ8ptqcE0MR/g7/2z9D6Qk79Z95I+X4gF9suEsMw0
KBebOgV+fyO30fDyC47YXpQs28C9/XIZ1yMjWVqEidAA9PcCNLEMFCZzIg3zNAJu49o9gPl7JgFX
Lg1Hgu++4TIIWuG61oeVWNlQHo63q9ewXVqw6YnGuRlPMtPsJKqEdsQ71oYF8x/zaWBulFy2Zioc
d7SK/eZGXA/FEJvzqCmrw0nv4Kit1IqVYG76q9J1khyshO8hls+s0lW1C0/6QSywO1kGUEt47gZG
/N12GfJVW5w0HNqXHZylabGu9PxblP+xNBjTFWR30nAzPChrKWVs449Y9RBfGBCPXeCWpdMWt14E
eLgXEnZddWQxq/XCTOvGbiB1XaxtgrnSluT+uXZkFVrAhXixW3hstuyPqJ5YArtDvgRO35qI2kA8
zviCnQM1sNu9TGdjkqPmSTwOXtP9hyZurf/bPEsbyOwW/9fhpAruHoVIsEa50tPEYTuKBkWdxKx2
RAm0XZmZNzSsj+h4ydc10zPc5g6GohYaTdlpX0RxsbwVygi4NVOLgGqWpDpdA9El/mlbk6PsbKS0
B14M6qrOv+H74UH3Mz4RQEb9rDoo1rzSw1e4IB0lb1GyMVh36fVWsN6tCrgKgFlhCKesN35NIYb8
xV0sim1a9N+I/ReTd5XG7Cblviznv/6bzzGa4qOsYI16EDqyPU/h73gE773OTdB+QOC1afZm3JQ6
th2nNyzR8f74Te3yU3cRcqT8ULYNDI97kr3k5WLYB64z/YejAcfKukDdVhPUIqB1RL0QfQDdMt/y
FeM29F+B0WsajlMTshhCRl9nGTuu+c/C9q8SI2KZdzc0RKbkVHpYl+7Ol/RBP6SnnEFtNVxwA+7Q
rBOs8hHYQw1+miEZSCfdjFDrk4nop+UOCY4SJ9kvgBU5VG6j4B/uEBhUWfg0jVPPeB4HSWMr9JLc
HE6lP1M8KIl/8spaBgcqQ3bBew8DDJKgwDzLCg3Cl1cdRO+Xxyyu2wZaCSAWFaOrS6zZQJI5WCdH
ZA7sLx+wKuy/x7iM4Z+HM8VfrMo2DEGI0wy950NsKgUyP1zKJLVFzZv23Gcge1v0+JeFD5Vj19/p
q/5CxKR28BFd3sH9dmmotgiKfqLwGIraOsbl8dr3U32oSGHeMZDhgqcwA+kRWR24/aby1POoaLd4
NEwFv+LdBVOyRiTvbJci9Byjemy1gctcpNkMVRjGhYP71kIu/mDyXglLk9dlx3nAn3CioNJgTzkT
czZCLoiuaMA5R9sABQ7X4iU/zkO+vLBU/t/QtXvYJSpSx6AC+T59OUcuRWV3TDrGORLE/a4pbX7p
L4EZ/iidbDsUvIe6E9HRHzH06yRjv0OQo7pUChq84bZrNapzUcq6rocsxLw4j/8cBfzsb/lTg/iL
1zW/spGfdpARPe8Sb8Pv7o80FnVdu2CS4iHMqQOvckHcg4gmUR0eYWuNKiVOAepWW7xtuV1P1IAk
OnxiSaWUkYxmh2EIeCcEVSaQnDgu2U/9rz2LWQIRhlgWPLcHrpSU0gm9yiq0DkiUyISB+ehxbUXf
w88OJRhbidrmVi5bRiqyiaSCDQu5heioy8duzALzzCbH3umio+u9SKUYUMcZXqh8HA8ATdKupBNp
MGcvUt2figbge+MWoY/TY2ZAa9PuNoPb17LalEa0Wv2t65RHSv967ntMoKXxEXeJBiGe1TzU//Nw
lVbIBuAbCJprQi0r7LD0EV2lox0DGBzyauixB2zuo1V3RkOjxay46hfmIIOe+/5hI19WW4gI7bBQ
flV2bMIBWNUaz3oGGgLCA8TvTfcjqnOL1HB8yrIGrLxUNMkrFjw1EnUfvpGLFIxXsj3LrLUOH49U
hbWs/fzNaGf9MOJEq2jBFNbZwvmoSSibFr1zPco+9ISX7TAV09ZyBRhXx5+tXocyYrb+usx22wm6
bfeCTR4jrPa/in099lmO6nFXMtzgFYSb5U/flZZZO4028CGnGKCYIYlRkYJWU876TXFZdPS/veVn
0LIp0TcJFDGKokxzPPg/T3YUjvTf0ZEWI+sqUTjVybwcDmpl133L+5jncdlXvKoepQtAPEuRZyAC
yFLV+F0bhZ0btitT/nu0N89WP0aH6o/KLOPdPd84T8icrgwSafGxeUrVOEjbQ6c1QjPjCQ6EHN33
tOTeSz8fpacpEEM2F7clLJEfe8a0F/u9j+KixaaslCzj8i4DEPK3w/NjV3o41PwsmN70zJDaQ2Fj
zZZWZooysoo9RmLq0LLWPk88UM8Evna0aeONXylSIk0BTG+SKTUgyleqa3LWDZxg+RdPOJ/D7gsi
RWgqyJl+npJjtyQZ+dNxEJvcq86xJJbBkNMxmfxembq03LsFg7Ko4iNUkaYC5fNUSU5S4VaWQQJ5
WxXg+2nR4ntyWamTLX+Bd+tGDgcLUK7HicjVmSfm8oeFRxabcNPoqZx+JoJoH8ZGcc4QpGxbA8Xd
N8S6iGLhPK7kd8xAvirmorRiiDKf8qPTlCj/pxX2gkJZNJuxocW/NbsxAhXiw9KLBafMGfOh0kUP
YG9Qqt9gwgs1vk+G2poapytPA9oY3iRVFgxLO1wrvK+CYGj0nb5CKttOjj/gQ5U0lIQoDRkKy6Wx
E/x7wwMgZfmwtKiWxQzPERI8inZfJB0Q89AZAwDIhRsXE0WJfPxKSeGfArZhBuD7+6Iy99u1IvzN
mvrM+VKKpIa4VcyFs7GOJC1HxSkkKDb7PhBlsUNJIkFpJ5Ce1Jk++9Zy92zH04ht27CjoaPBZ4hY
gp68hamhXEIyn39EF4tSefv7cuRUWtsMEtWsjiWp5EdVPtUHflJx/YbpY5IzWlBW1IlVS+rIsEQR
nNmBSRbmU7AX6/gI0fVjjt/XiJF0qn7V/zeZ6nbbCWMSuG+0/n+9yfZ1mx4oEkQHcG7VRutExugT
FHaqFxFdqnZ1r5spLGC3vX84TyPj+xZ255X7JpBBJ5biL4vTm/cZNvTH5E83K+1ElFyPoVpWC2fe
uPahnyhWMV3pewLT6jhZHtXQN125dJ9upIxTg34j8Lfuj0tTTXDe+xNqofqs1lByMLLlyh5oDloc
JhwcDp+c6Wn7rAr5cWRxLxa4OqhAZfuqNhRjH/1Qxz7nXKZ96RLZBigwCWD7UREg3NrGIkuhQrQS
8Beh2Fb9t+OVyQuCOi2gbEYebYAaqWRDdTlzkEn2Aa0yOCvrs5IfFX/OB6rwKDW1b2eZ+siNVc+y
OCM/mlStJuyVWG7Y9K6zHzupiKqufyTVjXW49eo1QLDxeu2lQ4nS9vlDM1kiKGjRDChc7kffaDJs
gv49K8bEyMKFBgJx//bEfrozCVCPkFQ2jCGUOaNLa2TWskixxPfbNXNd65Add03yH2JHKXRFx01X
kBWoNMzifcs/nZYdnlhRCuTF+g9iMdjG45T6fi5igkAxPmgySOPjXT0RGi3XQJxP9PzKPRyYBkXh
wvVj+hGsMvD8EDaYzh4unpukVYCKIn+6k60zq56FERwScQWb2UvS7ooSEbtAO/E4DP9ffm4WzqId
/lCgmNtN6Rs5e2K05cMN1YIeoe5r8Pvhv8NROsGVfH+Cr+BjwAxxRRHI96vZ9tTl2hNbDCDUgS9W
KebwwxIeCIgtZUlQ7OlSJOGP24Z+qJB7bM+n3PsCBLWzbmPmYLsQT1VyKZxf7CTI8peTb9/b1kVb
eQiO5RmJ44CtUZjyfqSUBKEiUVT01a4Op38jODVuhlY4rQ9nzAX0VFsY2WBw2xzWQ3TrNzpQGRKV
QhRS2vNxPCXfnAUdM+M5AbNxPUXjWa6c8kurCbq/eAORATRSc60O+MFKmMC6JAVVtae6t9MOXofQ
qyZUWpkhwl2GhXNVz1QB0522Pp6R2B9TvT1tayNf39iMTTGYHOh/qs2DRnZs1fH2vLLArmIzlTnP
qg87cfbFoOV8Hzkddkupo3tJ7KgoFh2+W+caVgHd3E73xOuCDbtZAiJN+qoyend8SAmF0xwf4UuZ
jy94l2Vvsjli2kzZdGeaVPubbpqJleVC6IYoQcC1PhwnDxQvkl7GrAwRU086LRQ1+a99SnkYiCWq
2anykOvm3/U08QBu3IvhfmN1weV5MLvcN452ndurE8bmk48B5KficQdFwbg5J75M9/LFmrwk+BPI
qox+QZ8WzZgH4WNwHDbp+vNKoUknz4cQdyVScASXhOJyfKj6kOQhINb9vir6+0RUDIeNrDMFdwVP
vfyogWp6ULM9g7GzfQWTKEWmvO6h0yXTMCm5fZ6uFaJl2UXc/gjlWX/+CW3gkY91PnKis780ge9m
21nJC7ER8OYyHqh3fg83bfcKlRaL5AmkGylVRzTJKjhQYosSLTFSgMwCJUM6arH3VG8QTfiI+UBq
suAlJBZxbXliCdb7I38zdYjFxWZhkunT8gOv4oMPYb14y5TuPFsnlEtn7FSnZUzRO8nJTgP1jyAS
EMN/UXT0rQjzyt1N7dE2ihFNJ/CTtD7bNXzXJ/9i1tMpJalj3wTSKvx8Px4blBoTKIW7rYH5jadr
/fAji4AmqEWzCV/tnOFJd091FQbEL6YgSlkcY22mtKdKWaMgba/+ACCyAkrrUhul3Di2lhS1Rybt
zrMXzLIQ593VBJKKk9SUY8avJL7vV58GOsP3UPDMmaWh8XJIy3OY/kg3Wry2//OiNSf7znZ2WtFm
FuDTuV67QH6jHSHQ2vmGOC4pl2za+6DdO9fG51jIsKnsfXEne2CRv0RuRO1NXtAkSARPRO9hSBf/
PmZO1wvcC3AvCuz7N4ZYjeTajLGgALU+MGuyH/xbtsozmK8no2owB9t4hivALFWiCvue1QTGSilv
ao64jgrD6xLdYbGe/BrwwibRSWFLIaB12onWN8LHrcOlz9jZbVtqaPnOdzBIS7tGbE3P58NkOegG
MF39XUW8ZjhBUWAwD4tcdfTQZePx9nHZRYnDYI+SJjcpn5m2fyZbew4Z0FBXxwgDZ8iqXCLCvES2
bwQ081EYK8JSI7WxVzvyyuRx5Jr13OYeVyliwKZoW5oeTTOrLXF/rcA0/wLK7ykeWtl+WYqsFMUA
o3AcFwIPTO3tjM7f8Z6xzA/qq3vbd8zrV9ZofNOrK1xtBdfGdTCgMfePxVc2lI0HyLRyZMCqvWuS
vlwDR78o+Bn+O+7p072wjfcG49NDEFkvRcmHBbRNNmDnkZtl8ENzCMpHcwXG2HZGekMweiJFR5uO
nmNPAKzh7kifQOV+CFCJI1xbGGG3CLeBiBhaqhJd4PE6I14hXlOKgSq8q2UjOW/lBSNCS2VGpMPU
MUCu0ZGOxRfNHesBDLGhb5m8guE3TXplpq8yA4ZmQulvPm90KuDd71yMAezP9kdglqmBoXSC2DbB
22/gfuQmr7DTLeM2cyDJ3bOX6e4sS9Mb+WpZ9B83GV41zqiPGVDGhtueJvy1V+SsaqV2fsRSr511
czA4wX5oAANY7DHZEsNNEixt4hv9A9QmPZk8JyMZpdV/OlG3rAJQe00xV3cM7lU5fpTJ3eYJKG+M
WthCXCa8RvAREmiZ/fHKUNsKGzxf+gpN3HtWjuCrY2qn5T/+b/wv852IcevhGlY58Tq51AjG6yAU
Zi7VFa+ZbeOLjDa2sLtEwkjgfU0sGGgtVNGHoa6QNnyy3zk+NOijYSc9/kJdY/P9fBVjwSkI+H1G
bTO6qftTMy/j5zAzNiS8ACl3k7fnMslJaBpZlXzOSPmXyokgIOxb5EWcXBCistqLS5STPXhBlNYG
sqILb2raCGHYlzLevIJLFTLiqErwOKShjb81e9DJm8GdL69RuA8x+ddmT2J8r5oRGL0yL2eZTqkm
PZjME4/qFDqYaCdiKppE6Cyk1D7MTcLK0SP9f2cPEyvgXlZpPkqzWKFaDyM+bzrjo5rMz5uGJbSs
gvTVnDY1ZMT4KFw+dGjex1tNK5kzuOpnE1cO+QjIrlbaxkNOwYvdwXMdqwf9SPmpZQxLe3L1ARYL
xvpQhJaLqfmflGExqgQ9nUBd0zrLBcTyR244IYc1MVuBjyvH7kKzP1RLhFDEkMWKTgLJskqW2iSM
Nz6kCMelemxBhSR0FhQwUbP5QmB8TrNlQIIX9f7j9O61lkcI46WjgHcBrnhvlH+Zs3otwDIDj8qU
69DESRgzRkZ95D/8ix7siCsI8wI7qA9XI60pOtuSdhPkwpaM6OLL1E4xaor7GbsnSgk2Lj65NYRw
tdG8usjdsOgolDrehVaQXrIFV9CWkWMS+VsJUbimLosox2V3sdljrEGc+0qHxQhdalfDPKLMVbo8
qwAIJi8KGeT8XSBCorjRQH1n0tIXBkY2gtO1rw04ZudyEwfgCwr6R6bbmnfYOyL0cMbklAX2fYCd
CxMxPC55FdOSL32Iif9azA3YC1StyGTmZEIX+npq3YjHR+KOWKJeilwWx6U0XG6G0J7FUb7ZxDJO
oddBMHs/vVQIDfT2CAbgWbdpKyFoFLBBk26osz+kCHJEqFkcMSQQbjsMDEzD32A/lLauaCMiTP1/
IuOY4zkgZs7Ce9BTKNYoM4F6bweU57lPp6K/7ZUlFd+QJNxVEmnS+i509GXz/kYpcUOmOQGSjo5Q
wXkQKOe7ZALtM+DrWCWb7dFaLYIznmkFbSh+WUmP/Z8lKf2cxTSaLWV1qKqVOciTnja/NpAM+w9P
eP2QgxDzMBQ5v2/9/jvx44VEAk4RO1w2IcI/L89gWy8c+R6lbdKg7xegtUwu2SRN+qYw5j3yIfna
8eC4QmIlegpCbeiAqsNZGZoDP+cCMJDs/6AWeSX9OV8m7o7znfGYDK67MmLifLmfIquqrgman4fe
AdTRQ7FAzIL2QYN1GlSCnndC2RKmnMxdw3Rvx+tm1k92Kj7jXxlBtJsWzV5RXlj9AuD4mTAU5NP0
0dP3PL3ThhP8QchijrhW1f1EFzjKnJtDEyQL9Z2+o3hwqwYUBe2fI3OrfOEjkpmRn2/cqWQv1yXL
Y5DHw81s1KJQLR5z5hRlg3CYr9bg/NILp31LCjai9ZGdErifSm/57BqV01f8mlUwwWEu+r3Yc0aU
aCi156nxOVgTT5AyhBHfBRT4tMQor/pjpU78MQWabklsy3kDIsLeTl+xQAOhLhhjUFZSy8o66gRf
TBOP8w5ID2Is+RNZ9YW5qCWw8COYE8zrxCyd2hyIOvwgMJytQAe12YmSau+Gty88GEgzIhJMw/tR
ujVmfb+q3rGgAQa7vnZSeabJnVpvTgudvMfwwyvN8vfdAmvtURnd0SeCOmvNmLIyFZ957EfT7vKm
zi8YqRqMr/Lg7xfilAPFnEVBMfUWLuFRKdap28Y5/bihEE7sS4YLiAQ7jgCRrZKQL0vz+8eIGbou
nYX0iAFyqpR5beyR1t3T7nsYLN+qYHefq0Zk/ZU0HdAdhVR8QUY2tQaElZtXuGgUBnUvbrJUl9QC
IXJX2LC/LNydRNwbobF943burjc+7GeD9w4k+JBWpBTVMO4vVHitMXhjUYy0bpvf9UWccuyMjLaN
bRmG+3L+fhMzdysvm52F4aTv2HiIdfDBVHT93eJzDEkV0vuCJjK7dWFNSw1hB0Xy7z05Hg3Z4fcN
sQ97ISurZ90INF2CM2fl0sCFG/flB6VcS4EflM9G5gamcQ6JQv4kFNYbUYCDLOSX4jREWqoyvJBl
CY3gpiAvmafZ1QB+/xS+jXEwwST1PFdXHaw0vnZ+GCX/mpi3BzKm/dIU3iPcwLd4ATwclfx4ydE0
GFJ63AMUrUoqtR2c0YFHDGJFxO+ctgu21+cLH0pTpyT1dz5guJbpeRmvLoNTGqbY8tcKnPJypYe/
s7x9yl2l7+7ViQIU01YaAqnTanHVJdNUdK0ywWYNDlV89v3WgbTbCdYFnhHRBQCmwX2qyeT+c592
zjxkmMT6hdVWrUbxuXwCwQSL7Hh2QzmAubGFIK/PKzsfgFiAw2JP3K/xycpdXRZgo+fZT5uXxNwJ
aGXt4gUL5P0w9iVaSE2Htn7o8/XqjmD/he6vOC8r3/XG218E7/kmn3TzcnRcvaX8+7HbrqgBW+sl
zgE/Kk6nh1pXO+rZg7VzkohvzbUFTKdwgmXMoXTi4NgIfDWc3amAS7uyo4j6/VGWROBB6AgPmfbD
jwHRmv904nMJlfiz0BsUI+zeU20urxwp/5TR51xBIuzBtPVYbU3vAnD03nYzUfgCBl7tMc5wfcxn
QgQmdpYBT4WDvuh/5RxXYP4Xhg+B4iSmO2X9Ux3aI6jsoMt6A6sLkfBlIhwWy90x5K/nt+TE04qU
JIj8ph1HcSbhJ2h5bFWy0pjQXUS/amBpSAcx4LHDtblm+tYJR5Q1U1Qh0wMcVIBidvMycPk+Vzvt
ABxJ3rg4EUERG7Zos1L/FD+49gu7VlqIFwcojC4WI8/TTR7s75eJvCMBArlEkj4jaBzqAyM053TI
yXzmuTCrwn0ETseoE7VHwwxJvg5QX14cfoJK1Tc+7zp1PwaF7rc7vxOkSQsw2UQ6hpu+LfpKA5CL
F6DNNE6O/724qFJjuBQr9neyQBMK6GsOCxFV4IEJXrt4ObqUGq/S4gS2f9QHiybQLCimqfUjLRkG
gNruhXxt3oRAdft8nG84cWxMnyYKJ5UskuGTv7lQ/zC5cYTSq6xOZt+MlmAe39Yv9v9zQW9lplGZ
yNGtYXs+sOoVzdltp/l+6CpgZ9Ozq7f3kRnqxQZeMYZOEJB+3ZzXG4IyodfY6FpEzf0k9pIBZZWC
uieXh4dTiL8Horzsn0UYhh3AAAkspmAJkUH37j7VFZUJQ0o5vYXybKy6ZLYr6f6jK+NvB1Xig/TB
VAJ5Sxx8NZx+P1OqV4gzkOtm22C0JLPdRR2Sw1UbGUMRPpatpTVs3ZpVcIvWcuo7uiMwcpejyz7o
2equ8p01UV14eJ74C0iSgwVlWcMwnUvQStv9zf+6sMHQTfTpr8NTeAyogYx61dH+DePRGaDbMWTY
8lKjCVj/R2Cy7/Tv6llMepSHTqX/Ut8/fUYUG5x5AVXbmAjbW+qL6c+AzOIqCf+x3unx7eShbNef
I1EfsBeaazH8Ee7CQN8PbZbm++ZMk1eLc19JoRTlOER01eDWoZkCCdyzWlH4160bcz6O6AaTMgK+
/gX5PWWxwSHRWa/y26mUdvuPcXjsgimFexOi09bQzIaxuxcSR6nDozFgy0RSHk7x6rxNxulqC8XC
kHSNhOevkSEcJusfsUbKO4dUW8gsGf3gPK25kOkebltoMIyRHxau9Owmx9pZNwoHPTqHfQVbdwnJ
/NbMwUrqxHmzHN2O6Q6cqI1zTYR6l1aR7lc9GN4kQkj4TPuUeUVi0Tr2qPNJh9JzAL/2f5lRTIWS
1kOdsGSglubw7wjZ8ojAqpee0y72V+I30ivNBpPHppEx7QlBrOctl1QjPl5+T01yMev0NT3HvZ/0
cRAdyPXdnQkazCStchfNCxQRIIbjjT7gh7CiymI9Vt1eDfUtA/WxLh8XKkhqF+8GcxfACFOIZCn4
o4YSN+9xA2NGzATeb9UsmYCkAB39jpmGFGMcS9DuaW6PX818ZsBAQBg+btrXT4Fa0Y0JN/0hcVjY
vPZE+2MTERivQL5jSwTSx7xQi/+JFo7k9Nl8x7L6RddTLJdTBd8rqmDUjUqnwrn0LG5SpSTqYo/G
gDTeTgy+4edIbbQjOuCCOwiu8zdwtIMGAwmT9ku7kduA4FmLp1C+vkHxzVYEjhFI3Q2olTf3Hj7v
8jvwQp/CYREh/0lFD+h7sOhkm4qILS+cgYsNZXiaqorRxM2MBMJQiAMEt4n0kO4NsrdDZUpqjyZo
jZHzWnJsYkeBmzoT+ArVScPt25u4FHZbyji8VCK3b7lxgEsL0v/BadonPf+Zjky5BXfOzBCMUz7I
IjrV5iSqHoapKjM+EkepIlQp+AKvrR1H75YRRtKm+koKWEUowaLB5FEOZ4KAnBRKgguS6GMrbaN5
NERjwclmdA7cLaIuP1TAZqHIUSo5REg5JGC/MgoviZiAhDulzvty4+yuwZdjq/uxaZ+TaajOiVCb
hoBZDerx11qQR9wo28DMnkhhL2N/WFZgQ0+s2svnI0pkC7+qKrhvwNMqSTk+T5FCeZ1XUDYh8X9t
t72zs2bexZ5VBQ9KQyF2LWvVgHBthBXCMCf8yKweGKs3aIUY/G10GoaM8a3PUrwDHIsXIA+bBLAV
XJyibUpQY7VJYVvTzJKcDnrEe6GXXDMLlJZiozwRTke4NZG7Z79avEcLsigDLJME2wrZRMCbwmjf
1VTHUIojdHWm0VluNBcLSBxaCASW40GW2KKPConRp4iCBzJ4L/L9jW26Q0QC97dJHyvq0vx7b+Nx
mlmtfNa7rxxj3822kIHyetPq8wt83HChmRlXiMZSySCWQOdN+qpWiNZyGR90jGfUFCOou5iCFIXM
L6PsZGfh1UMDQpD3vgOgYw5l3Px/7hzEW3NBO/JF/fBz6Mp7f99klAh9wKh4HDLqW+IZY8TimX4w
2TydDkq/r6AWDyKD77K0MMAe6Bf9UbNdyTQmnncNvPWpLlsc49nKgBIUMJECcv5FdJSaczkRKt0n
d7uAUmEGrFSEgxJXeaFwjHpVyB7rM7yp3uV4jVxAg6c64ltja0763v3JfRGxHPqiWDnYJ1Wj7BBA
LCGD8lyeIw3ksiQ4TozMh4pxZLQAiGLUqiFv0XLfPIq80aYvKJRQAmcz7KN77q+Ihw7+vIXDVpcj
PoJ/LkezBuG3fw+8X7sSCwr1USlFL53a4sK2B0bLPAbaogKRUWExxf3FBuW9HhshE2UxTOYSNkhY
IK0+HQMEEKzEoln9wqgQdk4ZzWXL+bjfxbkVUXQodnKWIZ85R4IrQd0Mysr8t1jWT16Ag2Fjwj1n
jVfa8vfleAXtc1Sg6LQn4XzeS+ah//01SOZJ7nXNfsbPuy1H3GPc/bSy5L0I7WzMfPEipDXlfKSS
9fD+BPCLp2fuQsfqoMFR/u76m9iNVD2jhGg4TA6Szt93++Y17ZAG0zDt2IQNgdujpWHrbZZFm2o2
bN1V7epUezVWv9o62Oyp49C65VMfd3lhIz2oKotFVmZFe+zwxb4xFP830Tnj3heNnpRPElhE1t8F
dmqnVR/ojq/hy435PtTvzqzZevPYG4YGnaFG13RnNbPhkID9dUwtxRueGnoLoaHQRjV83W09o4rE
0PELUPsLZ1aZLZigoli9faGgulLIJ+NG7DjlBoaCwBlsm7OcWpLX1DftQ1sbq8SBiYmaLNyTvWGo
PXwp5Qfms/1CuAjMXOewPmLPWK4qKC7F+k7plk0v1P9xQv/2687ag3JkpnPkV/9TcUDuHkK0vaJs
gUj5qnwNNUqO54SxgGOZCzeCmk7tFq4vFDeCXui4zRiaFUCngRTygrv/ELZ63OB0HKDITOMAwdIJ
nq6RzzD6WtwUCo4/+0P+fCwJyVfdmbVZji/+9GRnW7e3F9N+Q+ZwoCP8J7zqvHKOjivWGfVqT3d8
RF0m39Bc/3mOaCZqBUEe/FQBzv5fvXuUt3BXpjoR2CytFBW2QyYEpFeCHsPwpfpVTyVXfaAtgonf
HI6hwgotyo6rFxdC2Y5o9HSqXnd/9LcK4gYDciZwl+KtL/9kn8JNmC7wfAhYipk/igz9qo0hztsw
yMTjcoFK2UPgsyX2Et4pbt8Z5d9imp5vckn1MZ5qmQN9gULrf/TFWX3mZeWHlWZjAKNDPFzu5Kku
9hnWbzx5AeZ1UUp8kWbzykkeXCVxbZLsdql/z1h9Hsk877lXpSepfmHXwbbDBrp7l0OZaMgyKDDX
i8il+VxvOuNU/yH9VpQTa6Ufa+EL/es3LI/yzhUBTFfaktzbZzZyqylGIZxn4Z6iCA+m40YWRE0w
hXfnSJBqlmmvL0aqtL3RQJElHhvP8lifENKHCxaZCSp+kGWkqVqtM9rk9vo7PXJKBO/55qoT46EN
JemSeJOTyD6tL5g3Wxa7m3TzOaeYRC16cnzvEiRW9muw8uVM6BEnW4ZujOncub5B6rBwSLBBBYTH
Yz7TpXBvOtLixh0cSQNikHBgE96ECPpRBkYL6xI7A73324dRunHTWxlvD1oMDiCaG2uNDSviooEA
mzv/EkIoGEFLu9uY7A5O+jLLJR3IAAkvhDZroAka4+dvwKuzLsT0x10TrHETJk8GCD9MtH0scsvJ
J9vyrDkPB6kHhZfAQuT7pnvAyMwFzpWeinBXlou4god3P3N3Pq7aN4v9gftt3m+h9sHlXuC4TB1Z
eEdYwmLAMuaGtL1hPLiuOhxXc/gGYvsdGJcSGj8+ypdetJ9gRsfyBm9o8Aalarwi3qOjgQ/ZMhNw
mJ80bbrbX9rZCMEsegIJ5fTC1kNvVyfhlt97P+7hKhiXFMxGuUP3toG1F49+ZHKEdrA/89+NVt+s
1xfLtyIi9MLiE1XS3GiHMJUT44Ka2+S8KuObu4PFC0xR+8o80rgj7DMEUld+xLXIkgJ9qwimIy8a
zXvKspKiSOuewXPOi+oWh+HqEYWoZx3ZJnOJwvHVnx0U4GxtEwW9elu+bTue9Yyxwj+7dxKsM1Ud
FokYVUffscxq7F01+yw0iVg+Gs6GYp9Vossw/clbt5YKdRyxjmwYwfxdoN8QP6h3t9wL3BcwFDyG
Z+GuBGtXJkEfk4sXhczjnDbf24PphjFepiWG+USdHNPnEZv4egKik/xGhfH+yvqw7cvuVp4ve5pG
+5XmdYiJG4RuMbKaxhDTopS7w2zz9k/7gucNMFDPqN5z3BiwiWLKEUR+qB9x45/py/MPLUaP2SyI
Bp8FSa13l6VMw1e8FtIDA0rv3UTDu2LTatQZUDnjVqB5JrGvm0ko4Rqkp2h6zEzlLhJXOUuDTNa+
Q8HnZTngda979juCGFnDXIlMGaN1Fo9Txi78WlqA0ZXfwyx4V+EF2n+m1fhetmJVHUHWFwj1Q/wg
Rtnk9YRQDIHm+Wx0yr2X9z6VxnfHDpdVBA/ozW1Nr0FrwJAahT3JsJCfUEfQY968gdiW6VDVjW8a
Y2xORVwDU/JON4BI3W0p1lq3ZgkO0ni4KNAYqZ9jqLE0CFttlHrdWj1LtMZT0IcRMrHxsX2XHTLj
3z8lCimxQUQgOcViue+SozS5ycqoCOiUg1pgmLF7uvAaTyV9NtnAnbJC/OX60M3Fx1C2wieNvlZ2
SE/UJXJB+U9Uc4BzvJp/TFbYeyBsuif2j8URQmDFjYfzwZPEJ2DFdsoIk8jTfyrNqVvNQ1IccxCf
RjtsI7MRg8+MLCCQWeH+xu6AYELngB2fu04VIFl0BZS3TCwfg5o21svHjnKXcD+KWuNWRlikCath
lXanSafGECAE8AxJbMYlk1tE7fgH3gAJB4SUbb0BmWf8+VWDAOlCVEd3Jd+d8pYu9YzukY4rxoDj
ynl+3A2EKOEA4Sq+PDPrOu96JVNTVC56svqsSz11jHgoVUdET0j1j8hVTDJXcgiJ31xs0Z+nJo3V
g89HOSIKrWQrB6Jzafn2VXnCLyXYUPPHFEyTLwH8j0G/Vk6QalHCtRuzw+qeCJzIwxD07D9Tk8/+
QAfUs5SjG4594CfoIhTBvnmsd7yob14jNK6+dA1bQCWfKhHFYIs3QrmFEDcoPkwubnaZUHEXeSab
+O/dNMi+vkoRH7GelXMBYyHje1dYgSCdE1/Cy+K8wBVjpRfoIXI1AVXABZiLAfuo3D7ZUbg0j52Y
jQSeNSyFutsZ6jw3nt6PPVX62/dnfUyUsrYDTspimxKw29bkGJojizeWmVFapJQvaAyCIXAKwmpx
PdVEwIPjw5wllCTLWAO2mzSA2CXZEUa+kikTD+ctqCgxJkVAymjuUtqkVM9zGMqZwvKueFW/YwFv
UICdcpGe4qW7daZ4MTS/l+QXKlUM/VPm62797RCKDs2jRU69v2e4P9ySGcq6zEhafCTVDLjhuFFK
PCPsJ3cnPqBJOvogmlZKDkZJBdBJg1W1+tULl544TlsvxBhQWhyuuKi2fygtBhC3ZPTRZvQes5U7
o8huCjbVLB3TLgfeiIzGqudnQ6Mcly6kDT7clxP19Vc8b04MU2zL2S/ZyVsMAR4VM8cnYhcYeINc
uekpckk4iUxV0XMQDQomRJi9jfL7s1xiHXS8NU+2LT5gK7agCJa7zRSGjY98H8k1zHu+UmG77k4X
VBmOVI2pF2Mgiz/d9205R4WN0dFz1iadN+Sw78UBdzbZ4zxcetNyUSOceqO/LkBWc43TNjC2I5Pf
ax8NH5IcoFgvFPTizU4sQqnZBe6yySCAAnHmHFgn5vNZvH/PXVCofyHmvI9YPgw0sdzC5wspe+oY
sN7turRGvHtwfKicm/kWXZJqz7AHIZH5Lm2ecAMx5FNLtgVqTzgdeqTnAOX5LRQsau/vUTjI4Jmd
octBo8UzU0IGClt6ON9BVfJeXtRmRVMTqLROiDf+w8bQtRpBByha81b8TAhZUgNBajFOVGYsA1tv
AqUaYGdwFVzIJXFlGTLNPUMil3hKRRCMvSp14XwbbBTgZyXmiy+rCR1Lyrbr01vntp3srfT/5BIQ
b+VkR1QWbuYftG/aqxaXv7cVhruXfctUE0yLjf1o0ZIcQENhsM/YI7vWO3J6KIzW4dmhi4Nbaa7v
pyVJU7OtkSmkHG/nIM1+IC1UopwXhpPUoL9VdDJtKjLY2VOhgRhKc/AX1bKEAiaig/8bhNGNYoU1
BuE4TM80jIazrzHHeo6B1HQj1GN9jnXETeJPzNuIZQ1VJn/uzZ3pSr90gywynqZMyfS93/cIgsQA
ECO/HSdYw9pe/iKhKEhvQgSIOXfsTiMbzOP991iCTVfxOYGIAR4I2zifbMHp8cekCa0oGjRzjCQu
FCacVGzuR6XKsHrF3ZIwLXjuzGBVbhJ040yVnyxlA+GFJzm18v7FDj9Isdo9RZxt+1sr6qSwJ6XB
DfwlCvt/iQKE+CBrA72ZnEQg47W9PUQ1YptIZZ+ZE46D+PoRvgybd0CwRaodWbOcw61vw/J2PR+6
O9iVbIzQsZLanpChi6cMC7TBygGZWM3jwoEmB+pPFzriBVH/E9HmpGSmKlfzlpppcuxeUKQLOJe9
X34343z47KTx+keHOf9HxG+G2UcM0/K6fMmNqo/KJAXUqs+zPuFVgaVxAH+BV0P1raoWu63hzq9K
HbCUN0Gd+HDpJOG0GPROMxeg5vor1Spf5q3L9MQkr8r9KryaaDuh8XbexzZr4urMBjGwnHwZSCcs
CMdlyS0kmuHnXhYRCI9HBXlOF9u83Wx+b61c2HVzPZt7D3wPt+BcCuDYuWmEYT/EnnQDzcX0295D
MVn7SgsFSvlkFdOtgt/2AhqXuW160GDsMtA2tOtRQDS5C3jE8wpDHo2I2uI9KXoVxjnZoOlQ+Oo2
ElzfqvOzlDvEd0hfJWzb18RGEx347uP/TRdJCv1NzLp/UgDZZw7xWK6S/pardjyum8PITlpornVk
qG1d6MkTeBiYfkFsdyz2Z/wKgg97UnyzVnjaSlVdpuKnQhG1YKWEieUfqHDRbAYmqtlPWgPhK/AV
tBuNcQSSYcoy9edu87mSl5TMfvqnc8BkqM2cYn1jbZgcr6S/uaGbXkbnSGQ4AtmZBdfsyeLQ6AGx
EdFu0io40Wxmbs/zXkqcapxVJgB06zgAmOZ4yF4uRXhGBUudueBVQBMs14kOPCtmax5WlWiHISbL
Yihfc7/pBB0GvZFyX6qL9bf+tzhmw1cm1TKCIgY/4+4JYJAddgrNPkZ3iF2AgLByOaoW1wumu0Ag
g8PrfzXZ12hGF8A6G6l8bcMUmhL6dOXhKDexdsZV+McKnLuAIyCa5+QuJgILEauJy7rQBeYXzn8f
+F47vEdAWjAoLHEPGWs5p8QziqDuB6ir1EI3DpurZ4DiStmPR/I9EJflWmg3a0iKpm1skIOYpKH/
BKF4DbdxBsL0zv2TQKzOzWsO+QPsD28J5D8DaycOw0UIrK+Z3G1x85PWLtGA4OulojPZsmb+4rrs
jKvEGx00tsDT4Oye4KsnPsbasTMNSg4lGWaMTVXg1f73/opa9IM9JrCEGiYvJ0O3fM46Yk5lpkTo
eV8r7eELoWnsCgSd/lrTIxHs+kfawbzgcUHWlbmODlpO5ZUv3dLsN6ceA0LmtI6ASZYP36/BFPnU
6Rc660bGAZsKIL1keqZJQv0TqVy8jvkzkT6xB67kJD0ldSQ6iBXHpRMEHLmdkjW2yF+LMcHjPaRp
vHzfxz0xHyLg3zVRyLlKHFU6vqxKhEGnF3cbtl4/kMh3rIJ3nKsCPvw9LKScSrIvm3oTNDX+2QV4
3naktnZqIjKufBwjfed5IMFA5SqwymcV7F8vDbV4aTJcWCTV7tBs9EObAALrxHiMGo5hAu0ilZZn
aJD9bzMMKxhkTZppDv29HWTMxziyeHTQ4hhIMKXMNmI9xCDSRymRwD4A9WrF32HCo7i1GtW2XtXP
3RBwCX95thLCb/lrpJ668gMzDJgnA/ygo93bvpr9qvuZwIt8dt47EMTrRoT+Mts7ApACNQKaRgrl
Zdosc4LEBI2SAm1g+R+Isn8wcmp5yIs5xUaxgwJKisP5mJUyNWpEkt07mRB0kZnLBVRokPcRgp6/
SXFrQqBP9jjoxp0tCd1RLZoArx+RkXBkEO4MDAEN0VAQEYzBYsoxCgQ/c9hmI9uyemNaPRtvr5fL
EWqC9/HK4hsTbI5LE3OEdPTHS22AgPVtaIc8LCOxI5EGIqtrBxsHjoCq6NAq1bN2FWyBTZ/VdqrP
+DHEJyyscqomlkDPY60LhCsavAXmdOV9GnT2uK8JSxwPvL2ZWAF1A9Qyi6f+neMK7SfO+rIrDdgD
BU9tWTsDLPrlUTnFVDYALAoE9dEtx+EqrRqPFrX2OZJvqp7bMGIMRoWwb4+fcogbT1yDRhQ0FY6s
iSrAGQZSzqxSX6iuva8XZk5I5JiaI2WBE3eueEfTVxTfRpO6v1LHEYogGcn+OggI9Yl+rwpTnj9D
N3MXxPG22CJyTmtrV+CRGX3DspdVQ1bIna6Dq396mDK2onbE3b7aOJD/51wbkF4D8uHxM5D6c4iW
t9e2QJtQMbfHxFRc4Zsb7q/3w0zuwZSz2Baa1p2uvr4QXIwWAOBG5dKLoa0oGM7MIxOi4bu1DxIO
JiUUW+LNkgJVWcGk34Z70beilAZUT7dp4S4sWNPC/WMEubFeBRwrsZCdAAtTKXf8q/2DbATp+P8o
BpqJZS/Vb0+uIk+G8unyWhvO52bwN3uS/c9mDQJgmH/0jbxsMY8cITtAa0n6Vvof1cQuzRKRcQjv
jvk12iWoEsrleRrdPSimSKKEwxsiV/VDjNInuHeW+X7hdFtG5TdzVH6zKn8czt98I7vz5zWpQOtl
lAreVA0KaqqbA/lgDn8NOALV3ocNxACodsVkz0p5WAhYraFEY8/qIA/gj1zfoiKbchG+fV9eUtlh
FR4QAcp+g0u4VgvNkFA7Yfko9A0g1tlmr9+QIy1cXbksExuwl0XomYJuINrgIYbWAF3kAx/a93NA
Ulf1d+4MMvwiGeUjHY/G4o0wUPJQe0j2nZAHr2bEhQWimhdqWkI12ghufmkfnP7p3Ri8ETiVesCd
GtrVMA3r+Qr1d3CQN9JGgWM2W6IkyTUD18Y+ex9S/OKomMRIaZaRwyfK2TMw5FmX9t7KyrRgxl6u
Zf6ghMQ03V68oFuSOdz0h2AbAzDJ6RdbslJjJC2ifdawYkqn8TCu8fLgGxOXvnw+XMstouhcE2xd
ovRsdBU7cVk5OOHP7fr4UHNzRvvedWOyxe5ND77bo0v0qD+zipk9qDkpquxh9FSZxZqS4YoxjFXu
/PVlFofS7qTa0eRcL1JHTetj3+Gu1cyJXzluCRZ+tCvZF3BtQiEzYi/Jya1GfUtq10hjnqXlFHKz
EllIv0SVLTErOOFK6V4Wd23LmvZEK5uOMkIbhRAkKGWeay2RvkbmaQ2mCoRT4XsgDD/mmWk1tRY7
f09s4y91yZZf+sQW0RqjHEIBhXM84CDZy5EpRVV1pZzUUHnM8kH1r3KQYTk7JOzOSqFyGkPQr6L+
mwPf9xuyfaBdF+ZzpOHIif96pqKic30y+JzBAID5tL1stkByLbcXbWMrD+d9QvePQCkjIf198t4Y
AjY/DPIcO8qgnoTQMv3PufG6ZjU2nMd3fhLEj0mfrc1cFnHmdggaU1Ax5l+EfFjGDBvxcoT74y5u
gAxhKIa/OZfvxrNqayIB+8v/czB8pC4Fq/U1NMPn02sesEMvh0zdl6eyWzyssDtqRAxDEHOrCLek
65GzkEeVbkRDSxBbJX75fu7N54l+BlAkBvPBubTv2OtSAmTQZrJDwu8MWno+p6ISIva8EwNo4R4g
6J12VqumXH1qpCkKju58CKPznz9rbLsYgetl+dnYOJFz/y+6isD7C3xKUGo6Lw+HLzTEv0Hl3FMv
6n/A+nin6Fq/M3h+lGzrWu988PWQfpSFHpfweaG6pHx300maUSkNspbGGmZr4YM0UKT0pSuYReH/
wOPz0db+gYGRq+ubbuPsBYQmcXACwk8TxYJ9GMIh36gG/wjM++oDAaBpSrJr5MJJxK9oZThQEROP
C/IIoo97d99pLXFzKTI2GZeDH6OcsR+rzIFYkfFLnistOtCZo5KfZpJR8P4fmCACsIHswgv7hdMS
i5xAZVKkEMtYfvFcdcC9jj4nxwB+zLJ1qQ+gze6rapk1TsWU1SWZ07HoDrzgEqsEAij36ImT//u6
hnnTDXy9iFNlN+5M3H/chRAgzVPBQdpLM0d3EZYC9IQx3DeRpbnmYRjRfuytTDmI3kYqTPQXK4VO
/t0jcOPLU2ZJAxsG0qTadRPoRDgnjV/aL9OWCa+J7jF5/BlmS3NzOgvBL8f2lQw6+l9zqbzkXboE
qkogAYZD5rnu7pxEy0vTR8vxG+g2si9US7HOOYvov8fPrvEC+uDChBRl8DSM2JBZajpUSCgv9mWf
2CgFXNXtm4O1jajqMQZ2lIlX4/8RaDfWWGWqbn4FJGsksInIAv8z9u33l/OYdw49ByEV7RYU/unG
rvx+XYytbnaZUpL0w63kKG+GP9FdPAameH2VgTev0Lu6nz9ZvIs09hQx6XLZnu/mkgu1fOVxNSFa
H4iiLY13+aRERjTZhtVxIcKso3tYVc7aVM4ntTzRYebdKZQytRMRc+tQtcTBz/6D5iOlBzTwh2i2
0TcKw94ODVJZ9L0kSEFRyBTTgVXZiMcklWNFT1t6XYLaN9G4o/krLGm3X/c2w4fOiubwCdw/fqnn
krRuyP2vsGl8XOkhNBCgE+P6VhCWKYtCrCWBZXddlnUcPU1rnzZl27tx0Q9UR7b2U191zi4kWz6v
ho3zsw2NBzyMIXnCUBL+IYGlUuZc42XrppqzcQCiHBrb4W1g5Ft4qGfd6WjeYImFLUR/IWJ24arR
CFjZ2EvDl8mt37xPd+T23PwvLyxwyHir9ZrAHXXslZ9oaWkFVJtFxhjQaUbaoCuIXsZdSpkGQFud
ckFFNleETKvqjdk0+XFNFkpAohZmIp1Qxr0IiLTvwI7cK4fjP4XyHux3V3im45xQPDUIu9GPIsvf
U8zbPMRqmG+RF5dGBtliw0dSC/UGeUl40dfpvp1VgxCGxFTCWCS0uLu90f8E3bJevkGlcYLN6HVk
R3t96TWwlFx/Q0qVE7rJvr6t4ccPM9tDTqLaQjhjsbpGhFxgkVgmVU1BZ5hXSXxrQwPGgVIdYUv5
gbkyRUH0DcD6FOvhHz1XhMxuqlKho4TvcxBxoBr7g/kYM7PJmnjpb3IM0ptbSQlq2YF7KX+mB7uT
NHd6TU0gT8EOyX6Mdlkm2125g0dmmGiLrVUZ6n75Nxp+eMUW3iMeJeYGXw7pmp8Wu6vq898SEXy0
ntwrxBooCYyOHhOw4uAsfO+ZJmvfnsTtkppKF09wr0NVApahjWPMzXxqNVO2M9Zl9gYyZv7+/g5L
QkWUQ0NGD1GUAwJaPYjncpMAZXvO7zRTFU0h+27w5QFxgWnEI/uV/FyhIMP145x9Ja22aaTtroZ6
EGpkJkJA+BRQnrdOAsGpkYKjM3UOlbV1YZUhfkcLlpa922CTEryZ+UWCarYxaTv6acavRvn/SQep
9IeeIW6oYXwI2ArdFIGTCJ89ityTGt2DMpbxtKFB5bpYztTkcrvBtGdPgwnYq1Cgi6/lF/16ZrKY
lQV70nW+W/xI56fzBn56FhGiCRqdaOejxPZB0aoYsQeuyyLNrdJ3gJOTFlAypo2+9joGs9J7QZrv
Z6hgVJ5R9NXrgHT9DUAwjXI/5PluWkzX52ujO3HJ9tFkdHSYmFxoFqtYuojmT6LFFC7+CJue9yXZ
kC+xIvetL4lYYydyPTQCPDRShFD35edUBhS8dFbmC8E4D6SRhOhsiMrpjNDdSHmlsyPrMujEmR3P
sSlT7oJXM1/0tZ3ki60O+XHN8Bk/Edpy8o612VpM8UqYPuK1g0szFyjlpi7LLlUo1UHLYHDs8zui
7Yl9rVbsY49lesfXJBX0LLaJRHaccIORTWApDGMdMJL5tSog8vZp9cfWBqpXnK5LII/vTATdd/wA
q0GzUi5Y2VEPOhohKVgPRRDV/di2VGHDnU+q1xS1KRc5oV25ifHcBqjMHNTT/dS9VmnoQynk4xLq
1/k4Yqos287RSPrl/w0m6/ryCm/UwMfYcIye85zIei27f0YpIgQFP+mQC8I68l3uQSpwhRIjfgtI
tJ4BfwYat62qbSjOE1cTedxNqmHOkVm2XKGJyOHVUxfmoaL3DNRKb6XfXDUanVCJEZ43/Je5WyK8
/Q6Kz73cN3kAC8C7SejydfnHOnw9BWIz5lPFYWcw6tMJkhZt8yjJf678FDwzwZbVYE7nsguca1dc
368lOat2MxIhvTkUDTjshyDd3BZqFNT/B/8eCV3/ZILO+1PQvpk9aV9hs++lzn98QTvi7yMhVBli
0LB5LwuchtTTy1G0a5tA0DhHaW3qCCUvm9XbWy99FhAqr4uvvhUwT0TY3FEkADDxLntXfe8Nvu4r
GVJA0u53z0+sNtKU3Me+5BGNT6v6/ifxvzqkpvrciOL771SNIZBwy6Ozgemr8XCIxr80Hcpr8K28
WZm1kAUwhdYZ+hRLjIVUzcyTZA+fi2EU6ZPdQqucsksrl6BC5O131bKUpq1w7AQgn/apNZnA1KdT
+aMqlzACye/w/1SbjfmTnMdb6BoRKQCaTE/ThcBbolcLZHHQ+CY2fJZ3sLKlPE+s9OXxkoRuEP0k
AlD8U8sYdBNzyQNLlYjoeYsiqf348J2nN7GzodAzJqiRAiGvjL8MXG/AHFWbmRzGPty/SMQSsgcU
OvxMxryvO+DR+znzQ+KpSfoRF8+EKwbesCHDng78tD4joQSEP6I3R5ZHsB1LUTcOgrtxYWyEpke7
/lWr67/Ov968j9LVAhOzhb8YmJqQEPZONZw92xphIzRqMzsIDIqMw/Ajr8KcfDTnYM1ojqEZfIT+
oRJULS2ip6T3zE72YTumbuW6iFLpXoB3fVAW/+X/rpZtHvDUnJbfqsO+yM1IfkdbHN934F3V07dK
2FxzNDJwmmXnDLR66jTsishh7ukUPvChwoNmLGa3/PM07n9wL0RUWmjZ6XLbV5pi8KAAGIKoN5tL
ddMa0F01bc9L2uoNiphK1IVJV5xz2k13CnrnK2Ycuv1uUEbVdWhOErsUmD0GsCq5IoLqNqqZtpdf
w9bKl26xhNBLQ/y8+yQjE1Z1dVlMoi3KI19wa6IqQDGGdw1oSzkiIZpe4L5GdCXPgT0F2oGeKYj9
PLF4En1SFEU/1apQ2HU3S4sDhQ4/9PcC9ZI1wj5lI+0Hk7vwimSNX606R+lNn71RQKjv/l+3pMN8
ZAh9HBHX0LkyOxqlk/l6zz/mrFSZlhve3ZZ5SXYEPqy/fsIqQ7lIEOxR5zOUfd1anStcn45763o5
LsXxa8CynvY6JmVb1ImUiqZ8uLILMSiqbyiEkNcGyvobNyEy91EN1ltyv39dxnmwsMfO+E6EPL27
1CIumvN59iLUANxXxrbEuTNgbFFG0v60wUlKsgM9hE3XWaOqtOQ2pxwBmTsNDznsftADFZDzdRH5
7Xx2/lCi9bINJMjKoijPw5vftyM9YqvuT+921vMSgLB2ioyKRPpnkDd780AN2+LIxP8Jkqh/eVS+
RdnSG+Ui4nWOQee+wttClJB435ktHfmQlpx0G+uWhVZqZjT2f8BM8vnWt7z/2joMyNVhjpA66V9o
prVA9tnRLbRcA2Yufq8dU0OWagOnTRIyVHlN4EnfHhuUE+sIMr/MOCw65cOc/t3D49YwRQ+p5UuS
airgv+MUB1a4qygYthKY1rKpDffMG5bwBj0ah+jF4EgwlGNYPjliNH+ACesekPXYG4uQNP2z6nTw
PAY42vP324b/MLNlF8sr7g/WkTasl1mcgpDgNDouCE1Gzt3N4/Doxc5KynZ6aF6FGPkBMD+f+cfb
PM7FrJ76pZ3OtQMv4KHjL2S9c/pgYR9WJ2joVvQspwsHH3DcPnc2qD9YESAc6IiMWjqS3E+Dd8GI
Jb9m/2wTWii+QScVNjvIMGvzOqwogCzmlJaRfwUvEx/1ZEb/eWCzGTLvckNjOswAoAk1vzZE/4IM
PGP4GbHK9VSW5RNFLXPR1rwOWWeas2sUVInp544ODUspUxA9L0RLIvsQlYjYn1O6LtbflNYXCw4i
FM0eGfyA06sic5eRmtJ7fbmjeTu+3eEyUqIsHJmqVDcD/GJtuLRACIcFWJOab6W56H9wtLBH8zYS
7EeqYTmz2e4DopxcZdcvIJT9GKuLOqftmwW+Oq0lNlSCcpNH/qeXX/SeVNuWFG0G7JGUd8QlbjE+
FFbdp5JUrtJipUliuBQjyM+z4r/rnJ0IjFP16I/HVXQb+oZaWD6iJsOEwu+MWkpadfATdBAYAzAS
n0EgMwgUkhu8M9I6sYdwNx+SnocZ0j/CnqlAA01QH+ZgRBfuiSQ5kUdQTsh6ykWpa5Bsfe1u8Zlm
SFoZqEg3TdZNuSH4Jw3pT9o62/fcRdIHOfrLe0exelCtGwLHWTktx14syhBAhorFftPM82bL1Zk9
dizd0upkiI3lFVbi+7KwAUYX4htJup3R6vXItQS2v15DhqMrYGqgSf0cMj9y474PMLmx1KO/sElL
98X0ANs/qjiGNX4dHMcd42XDqsdQZRR4NSDNXRPAKFdjcipNGsUW22uud8ebY6shBCv/jqjxhUzy
2XHRW8t/nw9MM2mcgm/bRDjI1imI68AxfZCrWOwMMYkOFj+cLtd7epMPdWfaDodyJgamSSK8qp3c
ojF/0Q/XajWS9fGuAiIrL1uXhCjDjbUHV9NaWRwFDI9BykttkIoOZlQH/jfq/jHMF0c27AUWkt+K
+feQUIKji0uYlSq4z+fpLIaJa5brIrvOl2vE8G8TIyMtRm12ma73J8PhjvfqCy5iHxldO4cbevDn
rlQMlA2oG4dfmIDf+CyPbz8FQKvBMfuLl7JxUeJYGqucZ2oTLovwuAwS5rB2SgYfBe8Q+C8iE6sy
WGJU3SN/SvbsSv4f1icGCIvUHO9e4XwTmZrWR59QFCxkgPjoYGtPj8MobagwYZwvhqabsc6j/G/V
KVxTTV/K1MA3hijZcYGjgG4AT/UXYDDt1+U9givUiWqn6I/zF5dI4jN3cqPYVOw1hbCwuOt05xOP
phkJydjC/2ziYy8o5qPNxSDK3Yzb/XXFtZfBuhGTV8lsUs8R9N97HFCSAYOcNdskIfNkmEf+KTvQ
zUd5KtHwXQR/zVfSBDI1BySYsK4kBGp30KkpbS+/qSbdPeFc+y4LvhViC6E6azDyVZYxUCzKhyp1
wHUxXLvEmLDCMTDkP7XWAil0trHAEIgY9MNKCiM+op8VrKOlR+Moos4GCmuElcSvz6caW4nyeLlz
r+g1XHSovxHxmO3MJNY/5/OxttDspgESqw/S7ccPH4TBh8QLkSAKEMfHLIzDlmzzoomY7E96Qkkp
fzz6RNZXG+/e0oIP2mm9FbWdqIbPRFTV/n7eiplypL+D3VL/C6D7FuFxE0lfZ6INAbaIWQjHuCNg
PfscgFhA+pSr/JNY5wGPahVM3aknjhWYW4aN+Ex/EX4zQ0I99o1YXUesOPeXyTYzbCe7aQ3tHi3L
+S1nLQiljoEt5I1S7FWdhxkuTikV23Ovq8ZiHxexBUt0iEUSaRBEbqG8rAXbG/Jn3apTnzrED0ir
J4b1c+sH2HnXkk9HUTBBS0L5f+HqWlHTMG4hqOYMzbEK+zmMWB+ii9a2pymxHbbLcXHyW3+p3LV0
2/ku/bBOwr3wgPmKwgpT8r6ov9hv7sk/JKajB0Khx/ySemW/xq5yvYMaLu/9sel1AFIguwVFpY2C
OJMlwrh7uN1eHAknrWWtFCGprA1TPTaDpm+3QmnsqfhL2rdWYnCq7E7QVoke423T4IHfhuSanrqL
cFgqyT6vobR4jhWvdP+75Wenmm9GK3CigMsSVdx6Pn7SxJ6f8GF+dLgKq0Nc2AGqgpbuWzyBKWGa
FWrglDyer6BGTL2QP9jw0Urhv/lsvLH/itamrmD/8SV2Vz4I59iaf14m+Wxx7nLVQINrirUwO/Pe
jrrluENelo2ncCueXH4Ni80XvcoFpAKi2xT9698Nwi5rDIeADDVg7qpMufcB102bQORP2c049b1u
3vWFuCqiFXzOwSD+tlU9jN2wiHgbGA4+8V6zWU7lpDSJk9UkJH61CPZs4DK/YqgADP04GPBwnCAo
dW9+n/tqrOn28n2wV4VQk/pIwqjkLgJtG8GuY55hP+bqNhlhOc14LAecYZDgr0GDf5tscggs5oU4
lp4EJk1gADUgCuhGsLBN4+Zvozo4HwlUgjP4dOAVZpB0nubvXer8cChu2Mmr8/nIIOtBl3oZ5PHB
rtQ4/HxSnu6yztKuMQD5jXwKsRkaD/Xq9JvjN5RxBMouoArCaB8b4Mk4ON4b6eba9RrBv15RX10C
c1AWfQgOnK2hvZu3e99Xfie0sLKwHTCJUgeSoqDrI5EnRaF4KkVpJIi8EvEI75Meu42cTn295fSS
uO6Ss3KslvcqiQD9GttPJJj0wJKGvQ/DU7GZ82FpwbNevN4CSxx66KWn229+oyAujB5wgLPOiGsU
w0gHXS6rVS//5XYwmlC4BJXLiAfBQ3ZQlh6U9bDrutfNee5psp3Job/VcRb2Ff5UUiKHbHU4C3jX
e/MKVxx+LuNC908K09MpiETwirTPZB315aquYdmIcMJQOdKyfhMa8Nm1HgezHpyLpz/M7SCFN6kp
ZqZiVvdCyVLz8iHmHXEAErgifkQ6/JkKOVdatX8xhdJLHPwdmVG6wvugx1v3tJFemQv2J3SVoXjZ
Lk2aFP+MzS37Aw6tdd0KpGHQHRYY0qUf5DAbXeXzKc0qZkQJ6SZ08V9LG0R8/a8V/VPf/4bsdNB/
EdQRkO8hVIQvoEknEpBOqsET4L354bMKkXvqbE5fc/BWj74h3uVr6rjylvQKh3oAA4X0P7omZSXD
meUT0gpV67i7aIoDQKZxTlr9C1/kF0OhlqKNZd3bupZyH17sxxWPeEwQNIvEKc2lmfFzAR9wxpo7
HREL/dw8I+O+Wy7WrEVwUfmsB60oihEgUmdpPfkGxVFzC3JxdJTyY3Q1UoFXM4/DlWvsU4gd5Rid
8CCBTanJtRgCpa0vciLviiDoACE7ZjiFhN8jBY97xwWoyTbBLp6di/FqnlDT1o7uCUnV77U2CqxR
/5OGldKjidX/07djHkST2QqnahfSI3wiq3DBTJsRKgFbYyHFV/IVfND+y/rFs62dQJhoC4kJhy+C
tAlTdjRsaurxDBL6GOrM1nHG47qOuY0ZLFh9COulqlRezDL/fMkFpG1biOxgCrwPzEJtIoU4dZ+v
E3IOQXuLmWSLp8SLNyvl1z8AXdVIAZY0D5yYrMD2hnvJbZNicaW4BR9CMzsDaSxgcS9XvUlKLzwk
J3kkTQk7+KO/IAUYxubU0kuLEtLwsKZrGCE34KMN4zif0IM7fHe0VlCxTVNXdhCXRGLolJuEb5W4
//JliTNMdDajEAqrTMJvLjNfcXHdUznCqA85rk3OQuA6wgfX6Mq7gkk48AKt0v/mR5HAst71558d
d/j5XxM9NOoKFA78OyZvPJ5apsxbxM9FkQhBYcXlaQ3V0cOgOxzlTTMRBw9A9vzzBKYUD8ss422O
F1yXxe7ZNeIXpWojbGQ56cL7F6fd9AzLvHeSIQIphJs4z8dLTsQ5TdTXLrL/jlSuHYQddSWY++Hg
ToiQvnLoTbxEBgeiNNpixR+e3gIWNL/3MnmSsVuPNImfIXBhfHFIc65dpRvUqxrr1bpcJXUfugks
L+2jMg5LMPRbDAqIhCX6XIPGlx+y6MGzqwAMiauQRI4LW8GcPHHT+DbZmNhoWCIDT3/hX9+Pchd2
xZQrl80bHFvvhP8rWD/Izz3OwE55qCl8/EGFehf5w7nNwHWfOTS9Up13QeIBeUjwYY11tA5aa7xE
C5wIdPXAUyAhIOfcsfPhiwSbngiILn7z3kKPdya2/D3wOk3w7s/5W7VhJaC1fG0fAOPgjrsyL1TG
xvbUjU6U+SOWmwr74M9aU7rQ60+yzg/DaebD0hIjV7dXPwwq3EIybQcWXpvrRZ8G7BNVTP7ccMYG
yZ/rJpFFftFxdBamFAb+Ll/ADnv44ZC7QmBYPLK9gl1Tdf7TWseWezIDlUooMrHvMnXSb7Lxw7ro
WoeBh+IGOBvY+Rwd0fIF9RBbp/C5J5ben5+aM7Hljox02/D6zhnWwOd8N37wT8w/DQ04Hw3hXQgG
NIZpAyESMioNykDFnnufvV0mwKGIJZHLPBmdE5cMEd5p/hM3+eCK75XpA/EApSxK6DqMrVTczZRY
egBO4RB6kwrJWotg5iN9BW8w7P8r3VpZYjlgfgmqZTHiWKt6wfNYIxzWDsoHmPV1a/fbcQ9BSgZG
k5saa63bBBeOF+hyqNV/0JBKHbjyerLKOcb8iO5hEV2RxdXii47oa2WGReH8rLYnqBJwXhKJRlFg
2jiVRpp8/3JZrqokQ/ApWzZF681VDyneN3dxAehyrybvqz3CLNRxgjAT9RatRfYDwg4Mt5/D2FgZ
KbLJnbjlJ1lgg/jd412XixRE+ecsA4RHbUb48x57/qI9ZSK7UoAbBTlZk400OF3DIMVYyszLYF9b
RJNaLeOzCUDZAkHrVuc604LbqJUSJBQO/8w8uvq3MRby76MQsQhsioXGPa+U6FPT5Nu8IeRAspSH
Xn1e6SKzEp3GIBnLKp+RXpmMOjqjJBmcH09zEAVVaoGK0xwE2JwnQQtJwyoMh22bN1K4aTX9Kkko
I+DwgmOyDcGKJUPIzrzGYVXmgRR/V0Wh8jGC61kG6D3BDnAKGDo+ypFfrTn4S81pF68qP92PWZ6j
tN/V5sSd+PnTmAjwiOA+DAkhE1faYy7jCC+dWTzCtY2gkd/b7VMaAVEb4sl3po397IodPqcngskJ
3t/Yaa9lKz8vtaUmYLLIe88wzlMAuTD2CdK4DAhAFqScPJKgq2ICzCr31fPSaRYP8PzR6FNVk7OX
V2mWbiZ/WEhSTDxiEHxXTxGSuDpbgvdOHreV6hQ+RyglVo9BJX8kfaMJtIu+2r097hTJ9vzvN5ap
hqqOJ0OVMginIG+wzw4MpNwEZZGWeCtCEpdLWgC2HQqiVFz7492wBP7x7iDDOMxmT3VtsfnFDFQF
rjNqrXJDSPal+8l76Bqs7fwQhiPcbNn5aNYb/8A6WKwbekgt8LW/ME4fOq0NhvYrvwGTOdG+IPUe
JWl3SVBBIMCZEAs9929kOiFJwH0yqxGTuty7H9QsfNvP5ZJcK/vq4n8nEgwGruBMvkbQjiByHOBB
LyB4wHeCSjAIFqtrd7iWSPbsx7a4BAZBH/k9SZmVJGoyRvsTIT8MOYoMr+vheeK0kURYeteGRojl
Mi/QUkWx/zswv8R7wUQlRpefW+SqzR5iEGbfsHmBWVtPykC/hK2gkDWmI9ofaBO/Wms7ZfBfQjg4
ujVKSaBfSCk9y2hUbwvkqaGPlZI3wYv7BUu4Y2uouZaHLR7DsRd1mJlTMubW1KzHw0KuY66ONvDl
LXDHMmzXAEwxSoIbgFBE6m56f/s+M49ybCRnSduBWnTw6dzsv8qpJzTzCLKWjV8e0dJg9m+XzP5x
0wlcuLu1vwk2EMq4d89/ow95izzXMVhb28xxR3Uw+GVHAsTGmaV6PrHYWRq90oNZw//fcvUivUWa
QdQZBzYEVA8jMzAOQDB7oOe734V8G6jER32jhzWaisgaYcVywxFgTae2vXYTX0LoQ5L6KujuUs1O
w69Fv2qIBdsPzsMbgHpdgi+TDueXJJ/KGXNX3m9SrwhYTtuEb1ilgWH2kntzWlPge/ReV3xHSjWL
uXejWFEw/V2MOSiV0gx/x+7tIzA2NUpACcCqdAiXfc6IEQcXXZmd1O6xX6O0VNOKWUreqX+5dQmO
xGD6bPTtwaqrksnN+TjTaZr8WC8DxmBVLBrXebVNXATKU0KC2ocbIJWkybYNjdKkYbq0cutA/Uj5
whzjW8ZUGpoWNNzVBu+3Fy9q5uxNddVRqNxV7Plh7Fd7RcxHIlhZ7q1XuyJ2T2yH61C1QAuEDCJu
CkoGEuSTv5XXoqgfo4uDwV4LGMbMLp1Dh9tG5+IdKvoujpvYcgHU4u0V6+IoUyrv+VVH8tFirK0j
VyrGn/BueRwyDlaFtA0URKnGPotC7aQ/p/clER4MGeb9a+q22tKAmDklVc3ujlg2LuQ6gF24RYpU
90rpsbbrCgNaLfPwzQYx6VxNOkTUfJysriitmSIJi/BiJO33IvuXqXFxzV/tvknTEEEfVAM6oDqL
wCtjJe5IprXNzxxangbJ3EPNqwTSvYeTHqjS/yEpzzri1vu74eSP0krJ7gWKf+ln/qfJX1rShHi8
XZ+Fg2eCrRiFSwlnPOH52+YGthtrgDCgFq2eX+Q+BsYfm7LLsWgsRHwg4kdZdsgUiAJmoo2b8lrs
oQPoUSNGVFnEcjVI2r4Ox3+lqbzCC1yw3iad4D9E/vH0FoC/wvXgsEOy6xLf038X2FjETfWcDrt5
6hUaAqZAEWy6JsH618p5eXZ4o3tPmQo1tTIFnNyhoutVtx4B3Gm7Va3PW99+hbz+i7eMH8KgaDIQ
PAkVRYtsWKVrhM2YNrR2CjNu7TMQChLpeyp1YWne3A2iEppXwWEyM/WMPk3v5+LD1ErKIM512wmn
w1ASU0x4j5CTXvL0cmh+DdFyRsYNEDu1TVM5NUz+MNf5uhuU6NPpAzD953sBkQELqet1+GG1Q29o
/JmHwaV1BSmwWnA4Jaw6UpT8qfekYTtKbBYkbRFMUl+BOy4mn9vua81mTbqyar01eqdGGBWVv4rZ
qyqvqDmJzn1ntEdHJ9pvL0P/+IZgaq6teUutDuOloyzA3B1lu0XOV/PchLuMxEcy7JmKQ9RkggUq
9qtK4vhpoxhtTzU16GkoekP606cdjUGxhFeL5nr0R5xaEWTOVCzINBDYce3pPbeyZgOxFVa3An/m
vtGmvhWi89uy2kR+3lT3HmvmHsfymQy3cOf3Qc04HlmH4UegHu9nIMBLfRkuYb2RCWLqgn4elLqR
9YQX03WjJCw4gwskmet8HRbNpbvC1JEGR9/2L6nMF0NuIlcZHtz4dcI6rtt2B92pe0ODOxDgcbXu
i+i8kPE1Z1XWpi86nQBbjJpx0Y2efVTSz31sBMa1tcQEt4pINmLB9Lg8ONW6biWrBbQiziznVCo7
C8Ew78Y6vdtYao8QtGgbQf8H2InEZ9S285SHFJ/aGDyxw3uejVJ5axUIMHWpIaoFrKItaRpqZnQz
odgD7PM37XidxCDxG20+pL5IzqCi4VuSpC7fOGsCpBzLmvrAFRHdNOAvPXeT9MIt0Wa/Wt4tR8vh
y/Or/85o3hTCmolAYl4U2SvVD9YK4K8/CdxvmdTFbHqcQrdxA1pfQ2/IInHXWZeXhZjmqF+mTF+T
jGpkf69Uc305ytacS6O46bCb/irN4twAbVs/JP619YDk8sL8fYppvhA+PBxTABIy1Uu1Bjs3r6wq
JHI55g+Z5KwN9cIKMvZRLQIjfW1Q2wqng0ceWwLYbkYfTyepVM0u/FdY85y1hNFToKYbJRsbn/A4
sxM5CbIdESAFH+sdM1TKv1TTlwVP0c/PZ1XBvSAAVV8uzPBYgOeOMuv+fSvKfYCuKuiMf/ie0oxO
/oGjaqk53n3PMDDN1LkxybjlJPnEhfVQ/ltltwpYA72jV4IofG23/Yb8482Dv6FCVB13DyXCClvA
Bfw0R0gnmbtwKVcr8yZWDNIQVEn7FJahyI1eYJMbz/lWPWOVWG7B27P4m+8LCVZmd3eQHKAo/snB
5rbouYpzjKbaVeWPELzWaOYVkz84ETT/Yu1RYXoXkr1Ng25tHVEkcYGAmDHQ8FYBVNjIhuVCislr
m5T86nCx2Zr0ADvvhJV4MLi8pwiL4F9p1N72ytsIZ9aecJWVaVbWryXWIxNN2Scusx+s6t9kxHpe
V/+rmyP97uetow9b5f5uENOYqGYpxLE3bkavkxWJM/rsQF2ZnjLVlmWo8JUmgtJmniqjj9G/SEpo
qOiiDsCTwJaDsJFV501wMRSnqxfgpgh6zhBmwDDzoqdFu7DZO4SWUy2qS2Acihak7cfA6+sgzFAZ
vn4Allbbt2UnuO7vEybgcPfSQ4COoFe0oNfLiCIBOsSzOwIQ8OHE+8VhVL+e4VoNDzuPEwAZZLWS
yTW1KbeCbOAL2sbrfYAXl6u334lyMB2z4QKBVEJ7hPkqqD5w441daXJd4LLY4ewtdENzQyD7XTZw
xWGzfjv/cKEIwIoPOr5K/7hed4x+QRfT4NtmgpEDdVWanyKvFUcrt1mHqtav8K6NYAKDzMCQXxg6
nJUxVBelq4s+wtap4RNjR3DmiG5bC36xVBg5txrU4BTIRPs1apfV13jG1JxOS5cJrP7fpeJd5O9B
OFvPRss3iRSEKVkQtlYWczY7BtWqIGm+KDKDVyK0h5HpFfAjuW78Uts0k+UAzmnakFLUaph8q8Ua
SSm9hhxKVcJeFj+9foYz8ijr07agIZpHh9fZ665VT6+uYlIIrd9CB12/qMoTeRTPRvtwPZl3ll6U
uEWP0GeIV65F2/kSAyGkzZQiTeNe1BIJDdvMm9gZSlDwJhFJPt7Hv2RuOPCDY58MqOLmpNVQG/ht
J1NS3ztj/0yQ1Ye0IjYfbbIJqYR6oKuJ2SB2I7i1Zh+xSCesLxDWvXiu0aQVkT+/+VLw0N/OulZZ
5lB83U66zq/e/L0lUhXBPo/QCQmZ+9ceuz5vsHlVERpDxlMb4dii4qJRw6Ke81BRwQ5ai9N5F5XP
el1J756cFuEyFhBH6SgUayJrTcOKNw2BqPpWK7aV6Zv9Q5kZeae40fg5OtDAnd1KbqHUyhhevfXj
WXIw0unYntcUbS4TJGsFkUEaQtLdXWdWe68h/SfByxWMXQJvDXFgPu6dzV/eZlYEwpRrWVhfTTm+
dLlfgi1/h9UrL0ccF+rWWxMffK2fjg0SKfJrm1dhrurOT50cIP+LslWDv47Og1VWw5kdC3M4jJKv
Yg9tnx0QfR90Loi+QcIkQ4rI/WAmEfVj9VFZWYQdDsQFo3NXthKPIn5CQqEeH3sueN0OkMGFqErn
+qyQU/8vB02yIrGKICTXGF2BDOobWwqppzcLf6y7aTvzk7ZPQrwYjwesrVL4BDi3CXW+hv+3OZbu
KD+XCMljIWzXS1rTuT8YT/zetACu1L+5IgohWl57kRqiXr79CdmTAxDWkZyAcptQqCd7IZG+IcHJ
nltyihSFLfA+gm+zqsVLAnWASazI7/caFNo5n0Vmko0t+BZKaphppPz+qGDiFcrU11w5TXAxPM22
kiM519mLjEw1NLup0FI8dsXrIyLvkAMWlnlR4gDPHT0rtIUkmjkO4GbcCzZNtLXMvbnfnENj6tVi
aAZGR9/Y7f3A+X4E0io2zLFB34bbql8WOZRFfBMvHZLEd9torBJp5P+eDdCDcFuupIzkHYGwldA2
0Du/kvdGFskIHtPqhWOjcbjZWJXo/MsDq7uIVj6JBu1nii/Pe9jGyrT/8xrjTezu+pU6YyuVbZPG
HUdkL8FzdjccuqkGQL9+TgVl6sC6GbbdxN31xJqZFzMBxeP7mDJQWawhKUN2XbikmV5PDoDJUF3C
jtMe73uv4LvjijhoQAJhtBauhY0TXB97pA8KxRsyVX46cECnNnUX/zNKl6OEyYKTuk5Kj0Ch3GCv
2CHEvNrJHm/ro5xfA19qN2lt30ceJeEFyRrqXV5tTL3Q9G5g6ZWS4lB85LK3DHOD5Tlui8AnFWwx
g0jhAEzNB98l6uzkRbLq72Jnv/kYiD4iftpLvj1a3sAWnXxfLSe55YBhEojLxP928r4K2IHYLCni
/eN/ceRMkEOg6nQzxkA0lwq6ldm3+ecbYFUgG+M1JpICvom5xKNd2rGL0JP79duRnXzNzWSNuxnM
jQacKZlXgmGvdz0wJcOJonMxGHZBwNfYWsiya3LGGN/D3gteBuAZLEsTvxiBxxZDFjSR4fOJrDgv
NgNuk++By6ihlSB2WLL0SKv7x3PFPnqs7J46YenjXrfZpBnztsHQ+Ihvm6q1NWH8hVCFd2C0nCOS
o3/OtPPvLCptVsPBy5E/oV+urVgPHUckFui3nOfYG0kx16qVCDI4/x7HsqJ1kegoEbGeJxJm1JkN
I6pLFL9I0Iq/yCXbqSRnVdw5QVk6kPfbX9mLzlT2CyWNtX2IZYv+UNwWvlI0W39ED2/J8DriP03N
w/nq73Imi79x9uQnIFsQlZEwUMtiX1xJR00TDtcds82MlEXz3eSJ2UnTCfGQcSBPuERxitTsY9Vl
gVCeaYccTFzlevOTEUE8WdFzsOmbunn0HRr2LtCnoeb5sqUUMgby/p49x00WCkxmSiMpxl6d47nh
FgvNAAnkeq/vsHjIPyV5+62GysXjw5dUxGOCjZFmXG2K7tK5lWx6zw6Z+zgPQNRUg/xekH9aHP65
OFA/pHDyBPeoYau3sf9DZV0tOJAa5CmgHVPv8pfCSUXemzcBsZJvU9Y6CRh8GcEprh+5lUUpa77b
caAyG8yAJlNp373EprKZytsQG6brrAyEl2mm1wrbg91gejRACSBRPY3lq6EQw4g+9+U56d5FvgH3
1Rb8ikOe6+COGgrndFsUdJDFTmSP3aAz0Kp4HsEqMumb48BrsJETxD/WYy2pFODTnaMGW/11CdxL
91NbqYRDeLzrUwbNfrMkC66V7dF1L6gp0SY0BujCFBbs3wq3f9TSxCAvmWJhAVQ+Gsjsh7YxuAhW
xxb1HPyEgjccUOu8uRrzqSIbAI/kxRWgNoLxgcQoIhYcyQnsri/6IDcxjn7gIt3Vg8GlUTK3lJ8r
T5Tv4Sy7+gbvGoLTvfKxvreWHzpgFKM+71bm1ODHHY08t/oaYK8yLk+YHDgCVavvQBeSreu9bxaL
Rs6Cdf6mmr2CR8zjfXP6XnqFwXGyDzeNFN41RDS+lIExLOk4H2CjikbpRkPDp/7RPTFCFxYtP5zd
2vIZPtxMkDH+17TPS+Z1rVzpPHg7GiBhYJRCuecJFfj8mj397W5i5cGY2QumrL8SwNkgH78cQ7Xm
5KkmHrgSAR4Hm7Ci3gmuhrvZE0QW/EH8LzuRbwaW/n0uRAla4KMxN4byPh1Y0PKJEZFT5Y9gvLMh
8PIwWQxjfrKSYLciABejDLOiLriDvgMlzAFL6a9kXW4o0MbopEIaPgQE1JdcJJlv/x1fg6UtmdIX
F5uBZdnIeJYcEIMGbFNarZttJDId3ZVBzt6DVQytdqF+JWHYb3LvZ46B+Yi6jQv/Qkw1blCvhxH9
7SCkKCTiWVQt9xmec5JRcnhVZbAZi0epfCsdb9tmI4VzToxHju+O9ReA7tgDvpM9rwJ2D2j5uitX
J70N/gWF58Sad1WqmE9LT/Un+ynltT9UsLuhlR4n7PlJXF1N1x0F1W+4y68KUs5Pp3/o66KUUAeA
zdyNj3fN/H3noGf4sHDF4ZrfSkye7cMVQPoQKXd6wtiO1fCSzC7/7e+d68QO2FkgXpnhAIVZym54
DMNJUw9sjqf/xxBy9jxTmNLEp548p+00lCrZj1s4I++ClxGofXw0UQr15L/I3WjTgAP1hNIxsxZQ
6wKdQ7WFK4pXFhL9EHb4IhOWX+ufQvGGjVmKybYOIIX3reTJckfoCHX+82w8KM8K3P/QT2VjSYDH
nQFHeY4FRjX7ZqzOLAa/V0FGqIVgH9qWlZyyRRhYNUuLUa0hf7NSwUvF4qif/kktAiV6AZJCpLLJ
j0Wn5HLjMe+EcUYMSqFuOI1Ipkn6GcOmHnG37wVWOfaTKwWirKrrsfNnhiB2n6GEZpD29OFpvFTc
E/tn+z1N5zOiY5G0XyefncQqRQOGdahVvEAGCk3aKi3QAWUdRY8xP48LXy6C9wvHUknhc7QVrTxA
lzinYjiPpogYU9Tsa8yPc+DFUw96OnKmUwqXNphLz20lQbPulSrFN/0WKRA3eHJY/3Hx1HniQff3
aNiC1/1GlU9E44uiXuhlSJWX4Xqo3Urq8YIeYUfAtfp4mtc/CxVsRen6ixcis+KoH+6qQItpICVC
4jWm+ZCp8nBOhgZiVMukyWkKkTcti1YPThgIgXGj9ECGt837+XCHG+Ui+8IFFGa+tU9iK5ZgA8bM
mqyWHSjp5wjQz3ZxEb97JlwXQlLq6tfPvxMVRFZ6VUA662RNEBZq/ou2tsYutdJP5S7ziWgLzHf2
tbVXNWD0z7g13QFCbAQcsnaCG2f6gQuGaDB5AXh2nexAguCCMG/+1XhjZWZ4Ejj35GOR4rcAXfS0
oR0x1FOgwZoB7xjUymp3uwyDWnDP+6zdY4rUCTHLh8vEl65hwHeIASpr7/NArl25KgVyFx0qBbkm
cIjE9Cpdw6N/6n3L32DFUxMSMyJTHWmPBgBJ3shm/mqOMFclmMOWXHci+q2TBbWiVB4MzzDIW5Li
ofV1ogmdkTqGCSEwhtwVId0qRBaQXzWxnVT41bRH1/sWUfLMx1UOULlqikQ/fZUapwUHU+JK03v1
QoPRQbyB3Any9Kdduflyz9VSNG14HyHtFaulVpes2DZdE7SiIKdB6B/TTXRQCioJmplBu1J3kpPk
zrm3kpH+OJRk7NvHjCx95QD6NpUlREY39dpZOUIEXzhUphB/Tmf2Jh/KGbXzSWs4mZddpLAZba4E
iEKUnpMWCxKVCyZTjoKz0Vr+tAuh1bFYIZAFCjfbcNX+akk4D58ONNf6v+oKbaD3J+MaZXaqOXne
n7D3xqFSGLhRTAtm9w+1PVfdhOmqDxLLL7l1sl60iHWZP4M0JQAG7BWHgMKe+G8rwJ3QRwY7E7Bb
bHGPEs/YuA/pHkpyIhr7Q8mF2yGUkot/0TpiHIQH8qUyEA52kC8MRloiaFIjajOPaT1zqBbNLj6H
73XxgGIZeUnL72SReB4M9P4Ni3d6QtQ6Fk2mWPkOduxNU5JK8Ch2bnZMc52/+XxB3u52BXNJkTy5
PJpOFy5XtA7nRc4QkJovkfVEW0HNNewDnI/HAkTeNa/xUAVukckOvqw1XB31p/wj+EvlJ3rsbDwh
Q+kB5JyzyybJV/J4A4+vmXYySupFgsOfhOSz9EvcejQfy7+6UObqtwofIUgh3pcLlMPmSOeIsDdr
YIiibHrX9lX8U+v+ETroBHQZHl/Qga5QIEfPonDrUcXQSXmT30MD8lLBX06leWcRJtVRvmlHWcm2
Exks10mmHHdS5m1ZDvDNQCGWq6mzXbjHQvE5OMMzfz8YhQEabAj3s3b+gJJay7uWdZHP3NaGt9xI
EhL3JPR6AX4jA5LXTR+GG/tNIqDeAkX/Z/0deEYA4J9o9mJ/S6vanc6hDRYlnfG8HmJ5zSmfFcDX
mz7lfUGNAtUvpSwUmaroowFoO4cyW1kIb9/WoCEBiQwSavpRSdc1T+VZg+pCLVzfeI75HDly3wLf
5TEp5GkQXRmbxg44YPjX79NFe1xemb5Gkr5am2lRPgvwKUN3nsZol1CnQiDqa6unBSLTGFaqRNGO
q8D2rRcf5+Z2QPMFHJ/xvpZbjyKq8MW4gCqF9CeJzzec6pzNfio8bMjdqGWxtAeNilSyFrhf37Hd
AbCBJOy4UmqNT3+uLjFiGtcMyTPEsRrIIfCpE/5ZkVmcIIsHGdtzOj3oBUmohY5UWdS58COfyHb1
5VdBNq7/jUV8vWY5fv9+dZR64tg6Pmkp8gKuU4UresG9IBoqplEQ6B7Lo0dHHd9qsg5JZYRZ3Em2
1RTxsuGgzEpUcQh4f2cHY/GTv+2go6tykMmThVLmUNUy14CVfsaEs47VVx4+rAKi54pef1Wjs7Vj
L7D4oB0AuV0Jrz75IMi1mpwOEwRfTYIVZmNK2nVwY4ndVaHU9Z70HMk2emCXpJ59RbEInUufZGPP
uI30u85AujXgAvqIN+2mXdz8CbyYqxqEOSEHOIAVB1HZ4rQLf3MSQak6tv8jxe8fehkxmo6hNPXU
uLkJ/TI1d5wykXypMUh2DioeEIEIG6nFhxd0iro3CtAmu9nGu4hSRcIS6ewI8EOJZoJw6eats8b3
j6snqw+lqSbY5lp/RAcHRzKNtSwQXI755CtPjHN7wvZrfFQvGuht1NY3Jc0r7pm73tD6HxgcyMpQ
YyhZJ2oVaqiCNJCw43vzODSKudLfENYMhuyE7/DfkY0WEKpkRad24ArnI1pqIFF2sFO0xgZqxs6z
upLMNN5+2GgLlnY2Ss2tKw1ZJABwd90sSU7KSTRbEv7FYHR6rx9yt1wT1tCv5/SqlbBq/6MCa8YH
GkNUo2PL8lrnpYzCLO1eBYj/KRvrrHWGQsoCqQivFXICwpR5Y6WtBB/b+4hmdy3+hhKQWackDmJx
oy0Rz5qFQU8gOCaL9DJXMN3LEYjshgVtnbg9K+iS9Ll0pjy7ut3SLaVcee8yvfQIc3VlXtOLrgCD
2uCTb4DG8JW9GiPDn6JD1GUHWc2HKkjj7whkWXwpi/V6pcTaxWsuNqrOusD+6OQ7tMhuWbQU+KQZ
4YWKDGPADf5jSw7u9HUoZ4OuLbXqo1mBT4eA0vpzy8M+sux3AaS+8QjRT9PkbBfGjFH73Q4Dptyz
aR/yfEerK3ORMy7ILNKofsizmhbRQ2rLgYaNXxoQgIN+8gUYn96u2K3l0rkrKRVdyNpWtQ995l67
C+FcPScwKj6fr2lJxN1psXxgpCa9y1Ly5Y+8VgnHTbo8TUPRoKiBykLWcIXe5FD7TfjJnrZYMSWK
O0+0s49ye4BXPZ1eY9YFJbgWhK3XroNHNTR7U+KzFgh/ZDLm/UWbQUZGxsy7m/ZTmbuhddc/gxEJ
2YA8cssH/FHiyeG66kYlSp3P+NaIAlyPBxZtqy0xwAXwx/CQmbOsJLV6ztmmA1K0uZwp6wKwaIRo
ijdW7YSXK3IHjzNvG/AhIW8gUaTkW8ukQQbsLEQT8FHRw33QCzs0rKJMSC7UkBEdBpwSA3eo90g3
sLdDkJXuR25PktTIQS+IgTAX+QKvOflJYniSDCbO4HL4B50QZXbIl2YJ1oTXed6yTfr8CyeBjLsL
L3RCEaMcyxvRGlzXkwZWRqSdRfV0WDisnx+N6w0s/vq/Duinn8ZZ1Y/4LubrNtG8bi7CsKqCqWw4
7J/Lv/H9feRutiG/JMNp1AUEcxPKFbq0vKt5UpuB+YoTbUH+ve32DELg11eqODaAtRTWBy2UWhvV
txnOxX2Ajsps3CfwrFyf1R7FaJQnmL4OXL/QKBW25YPThFZ3wpXpr+kznrkoWisOxzSR7EKfgJIc
C4J4vOex9i5KpMWaaR/luxWHzPbg2twp+rWvQbwWRePdJso/H1nYA3hKDQJR+OuMVL9tW8NVUeCd
g8gIhsoW3fNsmZT8FXJbD3WPLNYGshGd75R77j/t913BdpvnZYjOkCNGhg7Pu3bh2/1uYhw3FX+1
SYnWjc4RXj2znukygC6eqCavPrlmMvwl3GUcOpPSaWyJhWQSlbAsS7D1ZPAsn+IKxKIA0VXDZLlK
BdkW3pD9P1G5dpzEpKPxUqTlIlcuc8bpTcubrN9bimxWHeuFV+o07Py6z2t5IHgrvRavCsiNeXiR
DtfxHsJieA6uMf5ukTdUpJPTOjN4KobOoejP8gTEkbPhq0GLjuEuHz55Sm0gbwmkl2M8jphA0Mam
Q13dnVSdGFGNRDXJw/+n8RpLt/Bmi042y3NQ50LOEP3lk4dUqN9ttpnNxYK277UjvDwjH3zPzVhL
rZjhnaYZsM/maWKKsXzM1SkC91qx7ulD7aMRdYJUbpVUOJ6kVmQ8DPB4liP0yDbBtHvl3VmD7KVv
ezphBVrv5aMXHXQwUbbfLeA1pbQb/fAu7EyBK6cFeVhJrPyDpDs7UohrJV/zhAH4ZliLOWNXdgOv
ZYkYBM7zWfDfeElO1feaCQef3gIhAF6EO6t8Ihjw5oQggXu1g2kK7+HBFWLuGITEVl1TQMBqNROS
EnPC98sTUDUvewNxFdcNOEUD/8foQ8LqBXj8rjsSSWH5ItPGnBwCyu+3MFVCw+oQ4AXC2qyOCnBR
T/n98TV5BANwYpy6x6VleS9QbZUpMV01mHm/CDCCRbj3H9P/ZDmq++EUJYEeA3RaWw4D02alfDww
w9ffe80OhItHh2HTrA/RgSylAMtjg38muG9rzaOQ4K2nSm2UHeWqcSZ28s+1quu2Kz3E2lpdcSB5
+XTZfnF7lgXTRuFDYlQHJOtp1womtyXV6lOgFmdWGvD8GrEFdILlxO3VKMJKi7n6y8bB/+xnDJD0
epIp4dcpo4hOxsLmbcqzf08ElNXusFKxBnONFvd2CAzWgu43LuHY5ebj+7IywWvQldt8jX4EOjq0
8kapfCxAJzY2ul9oyZJ8TvBmK6hkyXitTPJapwg2880CVQO4PTwsGQUqR9IkpQk1poyfnh8aLzJ3
J6uYsKMDVascWDFFLWcVeOSgZZGZ3tHPlmSciYQT7KnkMaXKkfQZD8bR0d7x+1xYFHcF/21/sHAM
KjHLo77QSW+ryjk1KQDEhlPmhCZa6IRP+3Ja99wxUcPthOFCQtkCYdKiOGh8NbOToezlL7HSw1/K
ywrO9PeELUICOnlAko4bFwPiW4TUmT31TDbR4dvAA26pFEAOmkRwCXV5cV1NTAf3XON9HoYtgafU
kYQm/lkV5zloNGUC680Kny+nbxK7dWnUqqYb69woeiGcyv9b3cvXVSvEWMHEpnZGbYYqM6JSjsCh
39YliMLz07Zj7BcNTK8pgV+nVC3ZhJbcMJKhtqxxY0RkMI6gJst1825jnyt/hOEll4RgPSI+acIf
DuKvyWGuQ1/13YvRrSKJlul5+HimgirmHV1APfNej9gFvzzu7pGLSXTsg2ZPoiTmjt8kraVf4Xj0
tOW0ifyGElcGtq/zLVBD70m/Pj1g40P3Rkwi4rBVcspGprWNAb58DbW3PKzjxKAD49RcQZ+niY5P
0UUutdYAp7ZwI5LQSrcK7yxF0KWaPaEBgbLvNYr/NnVfTwS8U64r53CFPts/smc2NTfJJkfzwitG
1dGSEGGHW0+zQGx7i0Fy3is4mjaAXCl/Aj17VaqPfwSJRvFywUvfH9Uux7H82Pw1M0PO73hx2ULL
3LmSMFHp8gnk70Voq0gygZgYySQQMdtSZBRYg23Nd71T0oVwlCjm0K+++qudjMWXIbUoUqNHTMPs
1I+0MlpHYPezGHHoZr7wNQHZzt+xSyIV6PZyPoL9lLXWR7+QBqE6tg7TuQt5sIQbm016X+6XEDTp
KxgW1hSm5KTE67nmehjjjn1OYrKKj0ja9PO5TsO92CXyGCiWgAQo5JxZlN1cMc0fBckxj0Fuy2Vl
wr2M0VykBgXoW/7KKYgJRtqWgg3tqyDJXnfcn0+TObwO4W+aRUyGAHRWsn8wWZRiNBWgAQs+ZfXg
GUkSSVW4UK70hiSyb121WY9UxDbBg89Cx0xDMgZO/kES/ukdkzLVZLAvwtFqOD61ThuuHGgVKRG7
6pjdH9WwgOnJAeYASzpk87kbrgoZLuu1s15/7YZ/OuKH5ZGGs6cdf6nmx6rUf4iIxMQO7Nsc7LQj
7fxsd3I70sT8nRQJegstq5Dq7uLqxKr7DOK6q5j7Z86xRLh0rcL3nNsNuV6RL784tieHWLt3aVVZ
6yB2vwiTS9s9E3gQV89QV9/d3EGaZr3PX9vQlM+naGSH+UOgV2ymTOH8BDh0jadegIvjdH9Vnx5t
OFmBuenvp9OPaoEG8htqVIzlLd3kcSR1Lj1dl1BFxjgWBP0OtcCjmOWSUjVDvSvyMWdAfPiUhrc3
JfZbr3mSJ1hnHx5G3YUw75OBWthhMnXetMb4oo/LI0Bwmhad1PPLwChGHS8TQwyAdMOMbd+S2QlX
Fyq/cFP7BKX4H3OPIbYzvY4FuGdTXXdffUX3leTi9zudGmNf33OjCZyZSADpWcn80rPXoN2v8UCH
UTGKd5P6npcqDLpQU+lLh/wbklvg2nyL19iUjf0gwxRZG+BGlnOd1FEY+2XrGWTC9Ekq/4u95M/w
ob0+b0lqyCzuBT3wmAqYil+VXYMucqVlYvLdGbOHT5kKhmqJGHfQNGHwrMcFllEbOfW0yApbdpmN
94x2oRb8ySDIxl6DOvYvW/t7XK65DMzLsVn+6NUMKP9Vc/BB31J1ZvVeCTMmeKjipxoebGPYcm7N
jtgfajSbp0hLWHdZoCCmS+0EoZxQONG2MFt/U24jqrh5LPAo9AN3CGv4AgGwkVzo5z9DkrGxd9HZ
1pLwlfuP1SnuJ8ystR8vJEKP7Cn+amxmF4oIaMuPIhpJOn8/IK57Rem+QhaeciWFhNDrqrr8Hi8Z
ohdRIk6H85PumVTcPrjrXzJ1BYPLqLfgG4Bv1aDp6ZIjSxC3EzuP5Uy4EaSiyciEWH6V+pb+dVDn
AgHYypg03w2QzsfkIiQgpCKQLZoE3GnLZdf0N9pFsNS3rnlaAN/51JdwNbzIWjY9EzJL7eTdwu1/
UflfHnHEiROWqHf2kh7XejFwWxuumsnZhMfr5yz2Ji/2W8GbqfuWK6nCnRzPBRjWeLcxI32pbg3A
DfB3bwtH6pNy/qU4ctpHE0/cZg50Ag7LjQ3OJpPOT1ZZv3jaCxcnSpvLP7de8PebUtmUWZZik9mE
Qj/UqB7uhFxT07sC3hq+bWXsBWYU1jBi05wX5STHjad02Se4lZYt5iyBdRY1A9hCHxdU111zYgwp
DKsaacHKCf0bzfH7ttITLOlDatjwJnaqiZk0B8L48vkGw7xlg/SEQpl4u9gv5badiiaXcJHaMI3m
uIEIJvrraIN7l6WYLFQho+u5ebEJtabXYSxLldS3OPjaOviaoCSOBmyXSC5bAm9YzSPuWIuIKkhO
/iNCkdLi3XwzLRwU+SHIwkSDwPO+clrHE93MtEUkgorO1WEeoY5jYQDxt1ElNy9npEO7ZkIu3J5G
CBBE8ktFRrhtIkOvlbiSmLoOky/8mNtFwDCrmeBkQt3UBjWhBaS+LznTLVFfinr6KH4Sr4cA7nRV
fdXk8oHgs0LT838OaBETCuTc5ZKu8ZNHHjHeP+t380Ei48oDtEkz+QCKAWWCVLhELt+QabnVw495
X/zL95zqEL3uWfJf79WGm62rKUizTDBizpRVSQ3EFJhfxXVBE4D1LAAu6aSJdTOCC86BGknVXAGN
HCYz1/RZNN88H7oE0VtAw6gcUsmsAg919kRFX9/ldwel7By404gm9+c5DB3LUqeWkW+01UCluWbm
VxTk1xrhrIONvtJZd8S29L6ygHNfo6vESzrrKAPRobvUq9XliW9nG27GVOJMi10msVhZ4EokhPwT
CSpnGBSnKudspfp06VevnU3l0ZMsi8pvvYg1HhBNLqlHfiJPJOQgY3BHr8hPsJSHb8DxP1nSAgF1
c1eDVbbRNX+F3lxnOzz54kqRoUpBprJaVTlucmyrG+fHpJ9SuWOwvcHSmfwWnWiYToDSipztcc48
nUjZ4w7n6JIYRcIGe7HFhAeLHk9JcIWK8whD0782EIIk4KbuOAgESbJ7vB0Uy+vntK3y8j0Liw1D
v2ZotoP4iTtX33kEdpycFhxjkS6SOCtvcBL9FiID/KAxhd0BmcSXlhMmVUG2AKn9yWpGhjLVKUE+
zRrsKJHtgyuKr7E+TqI/ULimnCQGWpKcpQw1oz+4wCIY2e5AL4uXUuKjF9c2/dJBASi/Shzt3DwU
Su07frzw8GGedKW8USEb0t3gKFR8bVOR/Meom6xzo4MLtokadqMCiHhU937EI7GwYx3QlHK1AmB6
4KUUp4Sgm342G6JTd2lXiVtqe3p6XJtJgtH0S9/qZYnM6ytl1HTSfCmZbXkOFEJblPezt3+XJfIk
yOAUeb8lR5IVvqDRSAY4jyRDkGMvHrIb6ks45rf+h4RAuUtGQJq5jqiCZeOrx3p5WzCLnX7Fko3H
DYUuZ4zTRAZVGBg+Etk8ph2Mf7VIeflXl/gc1P4VmWWHxaFGHzrLjGIRLE4GQBj0Am7KJUZPsWxE
r4p2Rwa6iOUoAxUoHLRGPsvgMo/HKaBmWM4lsUW/9R618FR9KueXpCBOtqjptaJFvRlOtyoT9EN6
IedrkJfBf0VbehTwQgr9JEebI0FF3HtBy2eG4JNkycH7ox3YHsBS7/3daHYRGc/soLkZQFvf6tHR
/al9ePUelhcm+rL718mB9T9oXwWw6G/+BbACpaheMNji3IFgI5V1vggeL11KUj40E3i4v+FKs+Ol
gBfLjKkPyJTf3FdKG/0YnyVsPVYFTEKK17riezjZFOKNG/cagIwF7jpcFk5QIl10h+ltZVdtzj7R
fK7PmDjduWIrzCErHWCgjaZlmR342KAE1vE0XYierN+X7JFlLcUESjtaN02PuB8uzzJ74I1NAvQj
nHIWYB+aPwKdHlkxHlY+95o8d8wmOJE809d779p4TAH4/CCQVcMHJEArMuZyyImkQKv3oR3sdpaQ
3VlWUx06od+ZkeRuuHJ8BCnJ3WGW3Xb4JdwgOkK1jcVKQY5QR9PhLIsotqNB5e3eBNAujsc5AIP6
ssXEFZaCNYA+ZYPCYv/djE38nhIT5vRpfm3VAHOvWSn4kGG7dJEcbv7MxTK3TCVS+yie3yKVMyRD
jy8iEAG9hV17TTNeoE7e9jjakIiLYgC2MJrMqrX+g/wnXO2to1Uo2lAWAh0qSwhnWrbC10ooMmIq
oA7Z1G1XLI+1mNV6zHCcJo8T+n3WDkcvz0/v7gneLHBpJPfvW8X9WrrKR37RM49hG6LmjcHwcONW
XS+NDmC2AvSYHlVGpCePOpvnu9XUCMfFVi+Wu3YmxTru8CXYfu8s7BK091Jm0BpoTIgMhJiHYglG
awo5QlrcPOwmL+wPdg4I+iQKp9sT8lnYLwe6BbXIjos0IFIOO9+8jqRxwDI1dePTx4U/bZ8gAZqO
TgsUt6oq64lQ0NWOyEe/UDrTEvqDblHPHAnHGjsk30pPyF+2sA+mfIcqEeF4oznWb1uSBCSVBqHs
bGe08dgXwmv1md9PBXTX7XzMn3I4ceF9rS0rJqkqhQXUel2fj2E27iQVYKBSktKqd6TeWLCTOVly
zFzheIRPZZH5Fa6+yMvYd2NCMjVDEb9Ph7tvLMXN3KJUyZEv4hTnqWmlouMFrEXxvhFzrzsbFAAr
6DwZybrKMk/qArcmJn8V6ObleSjzYJehOm9zmGyKnp3LVh9QMlXmc2dGxOAF3mnlaGHfgrML/0Qy
zjjlXy4u96JEm8eK/QvmR/Ps/A9NQevtnckID0eSrbaPR4uadH1+Q6WbczD5lBZ4yUxdYzE7VlaF
WZ7XWz7FK3Byy1HMa8sOIDCWdmVm47xa1hRV3pzxvwJm05Lcvw/e/Dx0jdDLDZIh+kxd2Jm43dJO
qKJpum+z4nxX3WfZWFd4ZvFq8iP1erIMzRa1FNEmRAtktaPHBNKmpQDct7vDOHxswUUeG3KYFf1Z
2B7g+USIwvvRU6gv+Of39WVH0JQThepAFHztSQoJxz1iAT/i51DaQqxMRA+Fcko5w/UcU2eyoIg0
jbGku0qtHm0Z6pp94tkEPdZpCo6vNa5cA50LtcufB7q1EatDmKi+nixP0b4tKikkMoi9qJYVSz4n
mLv4CWk5lQKw5MonSr7PNfCIMHKdA2wET+4vejikFEy0MkaxcrrjI1Wo6vOjLNrbymz2jxj+EzpY
AR74fKotKcc3qRfmXFmoUVcrvcJB9EAVpIXhwgJ63y0hwUVUFWMmHn1q6TEA06zBhTbaM/gTxdTi
U9WwtYT3DXYZsbK6tWO4s1zyYVcBE/2dJU6odc/1dK1fZ9AgMAftGAe7/SH1mhea4LfzH9mmgcnu
XDMMiSc9EQQLqYuEtE3nmr9l9KdIY/jRc8htDTZuZcjz74UUz33Fw9NfhzaWBomw5FjDyjCO2jnk
zQC2RBqqc82KRCdmKqRcY9dI6ICigBkkeQJeVjmas+IvW3G7G5lXbvHp5gc1oAIilLQHfndtEnzk
57zkDXnSEl5QReSb2JHu8rR00E0NZFK5/Snq885XdQu2m5hAg3EsktlB89s37k3KQya4N4qE5L3l
OzRgUFXJKkMVubRJeKXYxUQgEGGyPtyUyg/JU15A7u63KKbYYyE02mbciM2XsvwpDH7WaoAsP/mV
jIokR+v7k4B1rju4KRWwhifw/zNnAZqXjBVzkXSldrHikK49CYoj9yb+C2qTbepPH5IbJy9DpxrI
2rkNXjEQOCjRMrFqbFbu6voWfrJ/rQ5WxtPSTOVYSx3Y2qDeBnGggdCowTu+SjY7ct+JmSJ+5Sl4
oW5Qu4nh1JH1Wz+TpfskchriASJRPa4gymj6KGSeip5u8SjoUzCnob8twhSy60zN+yDL/Zgo6ZEs
07getAoCQj7YWc7X0U8L5TwmSLkPxdXz/pmn8//pQ4ALQln9KxvB9yykZPRbn9PJSQbA88zfWzhp
fqs0QGkj/7u0VVQeC9UnVbceq+8ZJqIDmV8b+oVDuGy8xAXY+rOh9o3V0Ofk8/QNuBNmnIaHGe/u
EP556VCGAqBjTRTrVAveBABDUzdqW11KAndr0ezlgsvoTM0OtDs+Yt5vxcZk3FaB85o7YKEGZ4Te
CTdcvSH/mQ4MC+vR4dKSu0r4bBblt6JayQQaRe0KgY77ToH4hAxawAAf1Cob/UTLPzm5UE8uK63W
7zqT9ETAznYwSIha347DFqBuutqi5KoypurZqmxY2lMaNaqKcH0Bhp5kTIsVP6UF9kEz/mZGaaIX
fJGGAnpSOF63nCm7xhzn8VOdUIKykOeHlI3222ijGL/n7LgALJFXTSwA0cXMGM58ifB2GLdOnPpu
JD8XGYJQu3MO/Vmi8QSfZ2R5ptkYn8QtfsbUPWv1Z0W7SGArHi+qij2ENa5CCHuMA+F4+xDEwQvY
lKkoD9uUnthWIo0bFwWmyRWJlwm7/cHO40iownQ1KY2D7sXFYq1WHAaMQ8fdfrDRKQ6hp1r9OSCz
2IHe3a5urDw6BVpho6pRJiDp8AMA0FVfeLuFbmOtVzJ8f92BilJXsWjoU4TZDFIt8R7w3YEL8s3Q
zXqbG5C67YOE0S+Ha6JqEg1LmBRFWmQTTTIysHCVq6lPje4+4KkjCqU6uQDF8Qrl8RUN/U7lzCIK
ld2AFcMAPpjErwDt+py6trQY8A1pOVrvq530+cvYZvL4IzA/v66O7KwQi11emEeKtWXiIJAhq6Ft
CjPpsIC7exWxpxV6vbjkfCFxq5tAQRsJhOQZ0ueFSqVwcIQ3ELhFuuRuJ9D0iGy1ZIN09naC1U3F
2cAoOSvVrLlqPnl8Hv/kFt5DZJZfCA4ls7ltdkmoEtLNRy/3rh5zu83Xauqrpp+cu0RlYLHKOWxI
6sqMsrUZ28HeLPqZsx1gFPpHLT9Y4KMpxBBF+5zHw3wjZrsYWP9aGnsnA2KFCqUFsMUOQNrUKC4f
eVtEkd4vmdI38xPEHuVykg1krmHhtJZ3CDJSKviD3RBA7OqArmoUheAxWO1rx49VNt58LHhJ2AGi
Qdd6+cLdUM1q8lrfrTzg9aFw5ebSNpqj7ua330lMFmrfP0K7rK/JietoJmlXRg2lA9+OR6OKJnIa
aT9fEMnWeBUf1X7AWcoZEyYXoDylgjhICAWaJquPy1/BZjSb8dcgjLEFI5dfL30UiVIMosFXXMsd
b4IADJPorayvZUBTbvtQ/QYYByCsjO0CKzuC6UPvjtg54gU6qRiDIP1B+IuMTxrl1b6I1laHbylQ
roq2StO0e/3BOc2qNCh8+9urqcCMR/AmvzWN+642fvIV/ev2wdE+XTDOEEJFtGf3IE+OYiQFLT56
VgCRVDyefOviS+GToL33os//+nA1+oEdQ5SmgKayHSs+Xp3kVwmplFsYldlZPyfyL0jq27p+PQfy
lYg5J7GT+O1meN24mjxFXAwpEWXWcjb4cSJyRywsCOgdnKGDi6A5O62u0TkMDa9Exi52wCBQ0dKO
wek4BySsw6lm98VTwQloldl0xkGcWbxN+ZziccIhMUJsUtVSgKUVv5J0tutZ9pxi01wpXydaLY/J
3ByphQSH8jkD0BGui815+Nn1Igdhqhpz1R51duejQoMBYC9o/bXI+z/U8bHkw68GwWOV1Wb3ielo
X8yPrbEFRMHTtYe7bo9l7AzeiHytdrZPxc+Kvb9YXSgvXN+o++9wPse2/fMR3oR+io/TuOZ/uQjM
cz3xqGW3PRO9T1nMYpKHhBCyYSp99Z+wogUio9CU1L2rp2pTAr8UWWytDq/bznBBsa6UYy7pB474
Lr0679aN6hAtXW4kSDRGDop2qgGHXf4q6yKR6AMxMa7+tELYA9HEDih5u+79P659CQOx8W0n+mhb
w9JP0RPpydJ15BLO7s91TXhz/N0Wax5b/J/HMYBnbb2FMtXOlx701fYjx8nyj/yVJKRNj6Sp/3zO
gjMb4UOkzcH9UXdyxvtI6Kj6cN5KBbQaevV8fhuKpXiXHyXXiOeYxgokWQOCzlQoBjD1YmLzgQFX
ZRUpYppm7cA0c6sykh3eM6XWktb2HTWOrOOBlFxMc47k009rDrFHdZkWRZ87+BIgsG1Y4lmOWyVO
HLmLM+18oQUiT+zgivRVVPzyPkFT6ANc3fDpnnQN4nzhLdk987sY1LplAhHfsqQ3xI9TwFkzLFtu
jK25Oq7CBDFNlKB9eaHNTwG/J2R++4KaTACG+5OXCWhPnkmn+hJAN/pWI2ZfgCnQj1hKqGF8fJWK
9BPbeN5Sexm7yyXp3PHMgWQ9VV9nQbXzbYnFlvJsYrffPxh8fkYTIfvGrSEMYrxZYKCfwYR5lBBH
f01CWh1p+SjlrlFxSEWUDmTAPZ5QA78eUoa9r8B0zUwBpgXV2OxkJesSdBKLvhPD+2dgh/LLq8wv
wTNWAQsKVOFF8qEOaZoNz3bZAH3/bj0ulILG2M0Yr9VXxg7n1NUdIaxBsYmpWBMBfSbhLF8rAU3y
J221ny+lDIlLPSQ9Cim7sX8ABbdZXEnld3Yyo+H/o0SOSUKtBJMA0ih4K4MG3QVcQzoRFzMfgfXU
FhagIsABktKDNGKmCi4swL8yOpPwxqIqxgXjGC96DXUsAzMG3Mxe7zhHtxS7plBAYsRLQSD2oEzR
FLmGoqvUdLClP+nney40Ce0yAkoV2C8GHuhniO69XUEftsEUoKnvC4M2pXR+IDFS56z81sQvDP70
khLpkei1NhCiog2YJBqNt3ovZcJ86qHnMWOn8dzdkN2B2jwkFCp+tbbhvbOfya4oCGO9HqxWUB4P
ZReXdCV+kOrC4acb0EMbbh4zUN0ankaYTOpzTV3YfugRyyFwy7PBt038kTCY4aD+wNcboCJTxhmn
TZUtJJLVEHqGLyzxVUT6mVHkFfEe36xj4BMSSG2FWTUINehEbAOpiaWGJShqDP8vO52M4mBQ9Yah
igi9nVze0rhTVRF8NHpU5gwH11majpKOsCueDF3/IdOOBrCnU+trQvbdmUj9d1/Ym8tav0BQsUE3
E0BO+qeFiGLvDodqJnEICdt4D2l0sqNfwWYup5ksikdDCQXUtkyW52S3ADn4LgRrSOTDwFo+RrFY
PSHmfcjn3URXfAVM9CaQcjuJc9fI1CmrJwT1QblwN+B/sISZuubIigRhwwrTlBnHWfZVaS/kwh3b
siCPhJxvz/mhaAF1dNXmKjtDtLhU+/sVxlG0y/bt9KpikvnSkjpHhQkAGOGJDCsVAQkU7pTEAQ92
rNxH2c80zm8txLkNpTxUHrUg5ptXLpiigbs4FjEzi3pCaSm3zt6EvDp42sqwQMpxNfCRSr2Azi73
KqMon/tsyKLFEf4NRGTMIRgzSerXz4yVUjps66EKqwcXsVaxnBdVo5lhyeGle/dxcYQ90D0d5ike
W1lhquQ+22Y5uDulLomPXrmnyyu3MAI/E7WD3HNjFqCwNAJ3z1puUbX1p14H8UPw5QfxJI/RoJHq
3IYUkvWIhhi29bBnJm/nBlBdMAn+RdqqOm6u25QVLZKhRf35HbILmdRICrDGk4UMZoI7y9qw6kre
iCwhfmvfLmUHuGwgeBw2TTjrfnWY7Ek6IFiMX1Cbtup1muxm5WnUOkufJh16St7eWzBJgradQ8JS
klXWV/tVZa051w/eFCHdKN5qJ4GFsinsZq9pmNqp/ReLLsmNowzLNwAFi35KmIr5e5x9ecL2P0SH
ddSQOXZisMhc3c/GChk+IuhmyzhajviipDnxgiWg7jxCIHlHd2pz6uWDlc5ujyYDTXMv23C2VC5M
AdznT6C5COnmUosGYH9iW7ijVgoz/frP/rET4XDXqtz3sqmK7KNotQ3QICHkd40zE68vu4W6QTPb
duwRO83j1NVbSRjlq9OTwmCvycQXveBqL8nNHkQvJEWKx1C2VijLk1HCplxyRN0BvexGfYEgi7gH
WnHXHsjMvSLVgApmjA/OfHBkJPTd0j1LWp6ZLHL5OffI0pPfCghwp+fdn2N2lofjeUwQpD+6a8y7
4NfNfiYdZghvRAPS/0Ubs2E3EkuER8gNKfe/EjERxM36Foh8lzxr5PaIj9SdJIUFkVAlEnr2Ok0s
sOpGFhpZOEU7RQYrq3g62zUlmRq2LIyxMCHYzDAsEQaRxD1XvAK2qdyKsfAs5X6VRXVMAR4wxnJi
xLgEGpid5judd4grtmq6zPjxHphKSAydAoVn585WSM/bVPJ2XPNikAMEYKTm2h62Wbesfkn6pVI8
IdCnw4F7V5uSSqFTUu8uH0C223Z+MRuuwq0g1W9cEEscVfYeFuXkhMjvrxDrfcSF70Mij1QdR+tj
Oz3BAhMQe6f8eeFPKJHukSpPvS8ut7f1STf730KqFpxqCjFt2Io22PEWs8YTbRHeXdb+B4u8qWOy
3u+dko0/bySaTYHHp1DD0cXxcxc7Dkqw7T8WIPOiRbS+XwG0gBCHX7KBz6N1RI/kCP/Ea00+Vo7J
GEK2FFCdBKeMb67eGkTabEgDtfDTFMCBMPlhO3gKYGvhAE8RuDPs0GHLC94hsx7qYXd53x2UVbfx
Z/KgAxvA467FvkXelCXaGGFTjwGLYJYvy/U40jiXUFv/GGb/ZO43bEogPdhUKkpvfN7WNcxR1LrU
E6i7Y7RctZDd64Yf14pcCxKLQcZN8exbiTT7QyVG5hBDr57qfpP4BNAJ5BSbtLS3oIqP369wDI6s
Yof4T2A25YBr5s1/++dTmBjFlx+b4NAvpvRhzJuDME+UcMXvpfuQp4k3KK577DPYTKg4LoKvyFuS
8RKyYJU6l5iSl9njD37ktJPC+4v3jJTmXItEuODHBRQCUcDwO+0kQSCFaLF8ssO/RvdGFQaiRnNT
g5CPXQ0IK4Q/4OzcDKXCWBT2PfjIcHKNTVDQZcVxgN5tlTUO8QPiw1P++H4idquDXlyfWbyyRW1M
MvIfDm3NtI5ovRL/gNQTvwNjLdCU3++QV+oLy/U2AGasUNtsSQCUZXKWZORQLHPZsAlBwDfbGioT
aXKj5RDwPa+3+dgt7vEelL5uoqRH8MsiEpBk29McENa1Aza4BwN0UB6vP3cxu0YTDYFfGoBXpSKe
sf+PZHoXxB/tDiWlJnB6R/Oz3M0IHtqG/mO7ZY2IqOy6+V3S3Ojj8G/UvOhBj6Y3ogYHDhvxkpLl
8DAJW5fNENsRABzXMTwqUiWxcMPvm6VCF+zy9ashkby1GKuH7TAHnWH+8RKxyqw0ofirHt5dVcWY
8OLrOiRRA/N9Hadm5oAmpV9O5glm4/Ct6eM+sNlaYBAh+2A7kt+1v+3qNs2c0Dc9z7QhdHIOESQJ
gkKLq2L6k9V9FT+GsSJGa4LqjDQn+RP50BCUbZH2iU2syxjzIYlaWaQPf2f7j1v72OU/SM2B/vX7
5pW8vIl4ofXJ4gL9rZtQTFqONb0s0WJuqRsWoZwJE4HFcZTfBrDr9vEAKd7y0dqM3qhOg6L1Ynu5
fqqfcLMf9e1GPjwmw8Cb2iVgv4yt12b6yB5leEM/UMrlNQCdRY3cxA5P9gky9i3x0QvI7vIKFBch
vTxgDGcKV2O/WZGtAiYbdzSFhUBLVXlu/bQaaJ7tCQ7XgUPjWt2Zzp+BmJTZc2sL0NBcFYYQVaSn
zERvhtiPzocvaSpjFr7TFIMMpJ/XEr4xSL2QZBbv0kKrJjS3K1Ok65nrp4ILh72PnJXLrrFiQU07
4L+5x49Xr64J2Bo5vZFnAUeY0fMXIoozL9G7z3khKChTjrZzzLMtQcl4d0aW+i2zQDvgBcXZsvGm
sdiR2cTggijmrp/Mr/lhp8HDxIDeSouJc4w/DNn++MGZi9QWEcRUZJ8Hf1HrPF9cVwcueGaJdcSU
RRfkd0SMV7DjrWJmHwbcU3qCVC3nSeMEPtidbaViOVeG0B6rD5i/Ozyt0FDOS1td80nX3GOyErlo
3t9mcrbdtCvGialK6WrxUIwVXYoqPkPnoS/rU9fcb+BsYv4CCfOxtIy/p1Z5vAcV/Kw74s/24hR3
jIiHtvIjUymu5z/ypGHd63hCtaazZwrEwVQavMj1SIMq9LA35V+NY54EgBP/ILL0aYze2DKSiDO0
f7s4FAYp8g8EfD7ioFY/WApnRlhc0QG0WX6Aht7fOV9ZZpJZMSxQnQSyj/BbdpSTwedztFOP+mJc
kIkJ0T6NsxfacAJk8al46u+g4W78OuBXjpBrDgUyIig5GxAp1IuVFBBY494otwTzyXFtG5vjthew
lBMYM8V9xzndeMEW60cjGgLBN5+Q6HWJ4lKVNffsttbZEsbFZGthLqa7vQxIAkPGFpynKw1YNkQt
XJPx0jRm5smAofJIeMINygBaCLMJlvG1qs44eEDLodXQok+ha6kYGEQy04TkEy17CIR8bLn+7Pdq
Xz4SivA3TXxcEHm/USpQS97eJb6SvulwU7cQef2XJUcreWAdrbMEgs2IjlDjCUIlfP14u0YYInue
WNY1cLdDPPK4KdHW8Zy/cUY+dIf5P9O1GpZf2DMrrnb14ky4qQZ8v+GxpG3hBr4eZIX550FNg9lF
uRneK7aRjkAf8nfxQznXnV3Aj6TWw2Kvoryfe8SNuTBWH59AaYxB55tOyopiKYLZ1r1eCMaVYMlY
Txu6bykyCMKCJyVfzlSwbBukJEEHxO5YHxcYn0fbqZq4wHwdHBgEfa0VUc8lf0yHeoJE8eKVxVGo
LlE/SoGWLLmg3mLfKdAgOxKEcfs+BRv/8gD9zYDAY9GIydQYcsAWy46k6XkCFj2SxdTphU+MuIVy
sQFETtSIQF7glCw9+P5Qk3MxxA8ozO0hXpcrSWhiRX4VV12tN05oGU3G5JMhgBpdz8JMCrFSU+i9
W9DkjVXT1hbriGP4lpsDq5glSLPaxBT4YTbAEGDnSbQWhmZ6ZdGanhd2E+nu6DCskSd4IsKxNcYH
pxBM64SOC7EekVGxj7HtSn8F7pWPm/3wkRUZBwTniKHIOscyUdKTv5FfSVKrotxhjmCQgd9s/ZQl
NTiQE/+I1mP0owFXy6tSkzuoNkZVXSNhz1nY4VC71J04Y0waCzBl3TN9SV7zyaZB34anHeCJshqO
hdlpZ7jMrtBpHa0HywdWSGVchTeef0w6ZN70eV5IPdXZ3pwcop4CeSDiTZcpTLO9XIlOXZckIzyP
xZn+mSlH6EXUyGzoJrTwR3ge/Fh6Nirb9gyS8+9jwahhcBzrXiXacP9R/aWaKBGFRp4mJkKLFNRE
kuASOYm/6hhP/k2VPScalBxILSaoaUp+65oL9NZrRUPLkIXOIrFswlY4SB3wG8G6dF0lhP2AUZBb
UV6FDMK0ZYfSVRLo2JZhhp3lw3fcvr7NPRx2v5eyAFjgu4jFeCEXiLYfW/C2IObHEIm8+fzK1WIS
oqNzIK0DVRPe6Qdn4OQ8Ex0OFsJ2hA8Fw/mOODu40e7IcBpilcLfId3EJurY842JYbGTtFTdLsE6
n15y2wsqsjdphxa1+NpaL1PipygWHIwRzDYJgClKhIHcYqSjq1UN/JqHyizlDf7HMVCI8PVUMfX9
Z/jCipEpIQCnJANVxkW3rMG/kcN9sqfchIc1a8/xGTtOD159fs9ahNVq8OTTeyelq1Wq0yOC4qq1
MNegK0ZYeYJvoMVY5z5ghwmewrruTnARqxUt7ygy93aUfb2GRseQjWE41Z5u7sg5E3oLvX6F1oOh
+SIMaYCW/XcDrDBDc0yWA+qv85d1i1E0aca1SUloEkBdsXprCD856ALfXSef7svMOk40RDNZOpk4
e+XLhqlqn6QSD0RNyxrJpj8iUL3QQTfjNGQoGKMzro1m5lyMFXivVdyg+A2YX9v7PwpVGm/MYJ0T
0USog0j2N48RxJFcwj7GkhjCSIsCvfEVrLUkhVtjTSpL4FAOd6D+YfL63qFcn+UyI8srZhKxZlPJ
emQ9KYUNUmBzoDQjqQ1YueR0NX7bG3Xllof+dnLWmDgCbDNgpa3cuSYodVDtrHlDwwf8D58pXdmn
07+LAIb5mWMUvEShVmmM51dtHj9pwV+8mwRC/KNVgSOTqCGYvbOqZJqOU5qFHcgHgb/rO2zhgO2A
GCmsmITt/C0MPDAVqxFtr2V7+uXAXTpAsJil1ehFhT153B72EVPV6BEiEhDu46do3r6GWa1zwl5X
Gj7lydq3ry5sChivcEv2i4peyyaUEWp7WZ8/RropnAo5RNU0cSsvxHN1MZL0RHf9+WXcwve5aOQy
+fgb/V+r2ytr3cdOeK8lr1tF6DBp+9JSE+LBJQMYlu/WZJhGrC3v2kKsX3WB0R3GF8azD+JNLlML
iv/q45goTd0L7Dj4Q9jnDWvldy/njcvkfKXhFAnJvyIp2/1xXks7VpGvkEUmhGSUDufTSizSTmvv
wJwRc/ip0T04BxJPNHAOWX4CpQwno7m2wO8GrGH/ERPGC4mYaUoY9ohCvd/UQ3U1m+ok+eBfMPoO
GSExmtYPwsmdmkGGmMZmaFNviLDX3KiGII+qDFuzgh5bGgjSRgpoTh/phkYXdOvjTz8FZ5f1HcHA
SVGW8aih6xm9BEiCuQcGwxa9Bvh/iDuOaNQ0PCFs9AdnpJLjgxunfrUoohcdJjybK+GOoH10McKE
RN+N6RX+26BPeNPO8gYcpI0ZkXLpdXOHY+ZXleCe97BzO+XZ6uVZ4Z2c0eY0OZkoVUN8K+jbyf9e
oDsERfZce2SRk5r01VcS3CgQXZhVQPxAOaG6ECzPKiZ1ovXnlNGKUnjjenn3gx6KwIsq9+p7PRg9
YcAr3JHBtHjqccGwKvJGqkGMxrOFHBz6q2eL5fXHv81BvnYwGwBkOkBqZ1a1ctLSv1SIMyXtbOdS
Hd8AGA89UcaZEZwOmgVf8cpntj1VTGvx61ucmRKRDDhykDlTxU0piClDAo0kIH72dNgfiB6M6art
n8Kl/GngwsTFTw8wyb5ZuiulirFzVLzaQxIPQ+ZSwCHYYx1yRUHEHCjm71Qv3+hw08CiZYZdMfKE
cJrQYplNxUIU5WHuhYMKMgPx4M5awz/htc7lcAa2a4/wvh2AllBB6zTjJcoLPjlYxV2PLajaEYaR
laGlhY68robPz4Lar4rOzbL5ZgABUmt84TLBq3FtM/qYK29g/L3PNKOjtrSBXzxemreWau1tbYvA
iYe7It+oLRyTzanayTqvXys6lqRKg+NVmXfuGDnsGYq0W4D87XyvBzzqMUAK6oOIeJfqoG7Atdqr
tJH6x0RBk+7NealL1PKy0cHp2RiJCJUSZH9PmNViqSKN3cDi0lq1cCfFs2nao5dHnsDf43hnzXQb
GykZQTK0ssz6V95XCr8mToNd5MulDEYhBRGhy2x71vIKAwD+DAsZ5zlyLp4nxBmwn7/T/Ecq2y2G
MKZNL22nEbDu6+86d5h3jga0DNGHe8Tuk1itQvwsluH8tKtFlaN4vYRxf9PEGDILz6Ig2ehq3Qjz
1RV0yYuUisCZ9N16qzpGrCrtkbkb1YNCZGAy4nSrNpBDSuRdLlz9hu3PFmT4G553V7BSNOrr4/jF
oke6OQsSSycuuqnG5KAIp2c3nAPt8od5Z4kV3XncnJx9vqz3JIVocGumdAIlGWlHykV9YGEnxG6q
qjWJpVTBLidAA3Ro6nOLaC8YMlAlhalkHiAQC0kDOMvhbqblrSj/lD0piFmwAgTZJ+RRmGQnXOtJ
fQyI5p/xjAdfLpjfxBqeQZoyymzkjZlxOoFShgjgaXLYLiT++z2MCpLVNssodxuaifjitLC+SaPW
pvqEaET9cSCQWYDyfE56RA6v74lzad6dJyIQW56xdZOg0ZxBvlrgdpY4eDd9ojWPmh9DQ3XJnAGY
uPhIr/FeRhcGrr4Ir0dssoF1bL+rG+gWxiYsZYPK5co895dg3KQPHlLy7obzk9t61wTK4BHpw9BP
3pIJPfQDrU1OxhE3o/f0+XtDV+jf1XDrtKvNZH350UT7s6yHLdetURixTm691kRBKDnQ4aHngDQi
hx6ZOoeeRlEk21fb88Y0oqjAzMEQeW9+wCI20886alQaVYru7R6S9YVMyKBaLJc3yryVtxwYM3p/
qWQJcWEolISrWc7xuKwanwBu3MM4y4fbZ8aD5eifvel30eZw8Rs3x2PE3Kly6ME22PF4ARrNxYEw
DXLawI9J4Z8Eg3T35/EWp9AJhIrmisjVkM+1dDqzu2uLrdYZgeyYWQtFW8Yy388wfFmmoP0yhNp+
h0gCFpuY6i1Wux1VDxAfrv0mbF5Im7IrIdinKhYIZF/lmDHLUgwfsAyoseku5LyPrZn+fjvBZPTM
sHfGIrtcUq0fhaQEHf+buAHPq0VSqzG9Vc5t8yie6IJtuK1LTKE3hf4ikXmB6t3FrRISL1P+fSDz
CrOPVAV3UUHiBI+oEVGkiLcx9BpOMPJ2+zH1cMpkD1YOjLt4ihOdJuhBNIpJym0mEfhs/5iJe9ZK
ptVNhl+SMvURnSLlxIV4mtZLdKjsFca8u7JkKEpFgzt5zP9+Y/L4CfR8U8bB/usaUEJ8adM5dvoh
wDSTU9UVvKCPhy/yeCbkWL781Wg0DTMlq2sQY5qodzzKm0iFg4JEYK2m94E4PsWmJ5YQQFD5hQy6
plHJ6WTI85CcR/bN13BikJvGR/M20/n6+ICmkHn/Y6U5uC8hx7WBibKZxtI2l/fCkhZ5z2k6PfN/
vNcErEzPnaQuFuh4XoKmRm3AvcgTRwjmChko1ri3eKyM4B9Vvv6YR7kL7E4d4dTx/97FadCYOH/Z
YXDeKbKpXURY2B388QpTBXI5a+DuYb6WMNcMSsOqEkzgr72IQDj+keLZMoZ1ax2t/T0MhbcIyLAZ
izOLrw0NDqArwQAZ0NJQHTtCUxDxs6S1lgS1xAvww0qtvafTV3AI8/zROPpOuFYfdyQqrgv7HdAJ
VVvvbIvOiK3elBgVP/Pf5X2Bm1ix2rzMoJABl6In6suCuZt3Hx+GaGWU6oufx1PenyZI2Dwax3QM
IIivgc2ECzrU9uXrERkNU0afdl7oW9MVU1hJyCRuTBgq1lOd0UriPS0ag3/v+jYlaqXfM6wofJnd
mSe791l02ahO1xxFR6EA9C1bvRHhH7maGZd9o0c44SCc+FfHIhpCdp4ODigoOSuSCYnrNXVc6zOZ
s43sYOCAdWxYlsJB021aASF/4ZHWrKc85lQ1CNsxz8rugcrqWoQLFkqXPQ2Q/WJBQYembFvs6/m4
cWLBX+BoySwDX6+KRjJ2DFEI0yQ4uguxR9nvduYI1qN4zxKa9kv18owQ8+Lz7IBLaH7uJ/xYxREU
5wHd1JrVZ9mSG9ky5No/pcO8GuZK49GGoQ/gmFEZwWrqoSbo2PvTXtg1DyhJZRMWacsENwg2QA/T
KvGowjG7KR6iCtBPNdhzn7R6d+HqsxdapZL9GIYttCDjCWrSGl6IC55KmL7DFL82pkDjHSJGsrPy
6sqM/tBdO5yn4ppP/OnxPSJmIAug8Y04J4sqt4Jt5HF1PEurvRr8BrsKDBUMifQ2VFIvP9qjsIbg
qdrawFMrHyqudLHL7c2JTWqILDbhDcwqoxcGqOOklolTPe/1ozamB1Aed4xVqMpnvtBK3Xj71t1W
ySdyZlbKrdofG9oRXJTFVcV55QdUuzh1ntgyj9eHBe4vOYg3xQkVNWwp4bFKRq72vCShAV4my/wh
UNNWK2xszZiD1hxXUgTxN5ML9HB8lS9wgHcvDZgRatG9qf5GpHvTDYGo+sEwTyTMdTaJONGa404n
IgA5GqSBPYgoibkwkPH1wNBx/OHD44APQqj5QROo+o+NH/LD/PsgLifqcHUoNgghSM1MmA4riQ5y
Cba8eJCQD3jaCxQF6/vWHMuJadAw3MLSck/uIhUUu0uOZQBW7wWEROw/S7XMZSU9z5iJs7A/+241
Lsy8qmK2RcVEnSVt5/IrnrK/QIgHD1lAkXVfnH8qPKlfLRrxEuCWtsv1RDxLl7Vasn9jdEZCRonc
EAb5+mZorUBjm0OyXNUmy04vjNV0KdpZQuyaKnqTiwIdjsVE12Qgc9J6I21rJKii2qY5K6a5YB4k
1AWtZapI3XamjigmLZvrFAIvilhyToGFY/WMoxiwfdTnU673BaYKtXlSv73VmMlU81/AD+bayCt3
N3x/19n+JlrIPGI3cPIYizUV89MbTYZLg3w4OBs8Osn/CQv/El3SaSxZbpO1K8XHQ0OEjon8kG1s
Q7pYNyNbcnNV8+FVwoDn8JteQiwC3cLwiljvZ/ASrbB/h+EChx2/YeCg8evJ8mXWx7lyaV1zTWU1
mjsmJUHbEyr9BOnjLCSNxd5+YoAkePfT8L+4BO4U7V0EhxTkAAbxnLCAk1DbjH7Lik09tPcvv4Vn
wEAYI3vW5Zgsh2kbhZqAjtPbkECWaq+lTABwxjstENO5JT5xng239miJ9tzjpahi6bmQLDKCr0mj
pfrXQ0PQRil7QBiVlqGGSW2XI8b5UYj1DsRADZXh70k5I+RjjaYSVOJY5892Ja4i6ZP0r3U1UMPH
zExPRRS7r2nwvmcRYMZc8XDdBKeo9JXY3vNUthblPQzvMoqCpBB69uL6nMZawww4qfC69hwRrXL6
8L5FmHHBjG4stzGOA6aHDX/RmGqRC+chxffEwxkpCniJXhn1ysSUXKF0RqKRYvq8eJ/B7jw2ejcY
5q8RN0aPLXyHU72/QYM6fX63C/Nuz7A4RErkDq/26qqjjqrSWteR56XprggReNL04xTKOZHTvXPM
3fPJATS/M2NRFwwsgE+cdETGcjq4u2U5JJrndDIYfP9MfRrVP2VpkYaql1prZgAiDyb+skM8ypdt
Uu0mqfShQZdV5/jVbKLuoMTLmH5pbNNa1MM66rPnhP0JeFf5mPZM94l6Zncbu/kBHkriUntB1Z2H
78cgbzREj4+NzkQmkhqScavXb2BvBK+uD5q+tu/r36Z8I347U4q9T0Hp1lxWekcCaBg0AX8xQb0q
dc689UlXUU6doIFJd5c55BAMAMHliRe3qJjOcAFKAcWU6LLccZxWJC/Z+rA5SGF8XKK7mNgHv4io
kb/2WZsa8bbHu9QC3k4rPuC6wxE/P01BtIfWXs3lgavqqMb9QUyOBYU0w5zarSJsgmF9DF3yTqCZ
6bidhcY4sihemr3v6AP5x/bjO+9qwST1jRfyYOKIqZ/jiXCVzSy8i/qbUL4Hzl5xQ6CDbmPH4Quh
Jhibkj2VItY+jXwhg1WL9Z68ygHKxkBl8+HPXy2+mQ2eSr0x+sseEPKgjfv1bbl49bOoIWgCDkJm
xF9mk6TWoLtGGM7XpZ3ncC6d0hL1eWvL5p3z4mI6QKxZE+f92xzxHA2YFy8kPT/X8vaoNrMj58w0
UpItI9J9S+XkPM0/ogA8j7sYYF1MpZ41ClwroYLW+1hbacCaT0P/TcAW8LZO2pgkUuNMxSodk1Sn
PWbcurDDTmOKA4SRUjjpXrWfTrdNe8oKnl3GMF7luZKCdWar3GKpbY/eMIDoxpecbIXCkfGCuFxR
R0VymlA/1xCd4b71xTyXMbGAqHwwvHeEJOJhqOIUqN5HPLwWx39mTehNTIYt2lp8GYVQ865noi7b
YzxERcf2uAjGAPywnkDoz3+WHkMTpBr8vhl5o/6/5/GHs5RtbWKPvvJdc+bXjrHAn4PnVt5FvlL+
7CcrlTOLKDy0p/LLruUecko/bj51zVbg65Fj00vebrsXtUCtKjAm/3eAa59X08hXivU6aweiI37t
rZFICTe5kDQX2C3bEqGISht1EiCYqcBXI4NrPiX8ME7bL4Akz7GOSsIn/lB5fzkDK5U6et98IFt1
Pf1hT5cbZLuu34P12FMURT0Aq3W9bNcwD4NnrvN5D4Gr+OTLp/jVW5sVGBDEmeKx2ksiVWZaW8k1
AFHQQjr55EyhaM6GcXz5yZ/N5INQj/rZjimvRdHBcilapNHn2+qwONBhxmZgmWbze0QwzQO+LbBZ
1KhPb8JNSIj6uPFl5hv7bR7vT2ZlVsBSr8QvZMLbGnhGE8efZeUWSKWQXAKLxee7oxJJ2ixSZVNk
VtT/Abwx1V+GnkkxFUMfSlJfQVB8+H1AIIFh5oIeSThpbnhS04kj/WFZUi9PLQHBDvcRGkQbtw94
0JMbMw7zQgaFSl9GkWetXqdDWe+XmES5lVHKfthWETKEPrtd9EFHdyWmKqX2mKv+OkjXkYBueEaY
bjsHL6MfrZQRa3Tvz91fENmPtj/SRH8bhZDVmtx793LrXIX+Qd1F1OXkafnWb0h3imNqUhFeufzt
pRrcm/WqA60WSpKgmcNDVC7FL17zpjpW1bG888yrpjQAicNwP8SilXV1Iz60GM1cAwd8uVYsFPRO
LD/gtEyYK+M7TZQcM3lgq6DF5Iya+cM7M6aIt5tpUSDx1kCIua6yAy85+0jTkSPSOAAZqItCT6rr
TITwfjioLzQdny472aPM6mUNoy333bPh4ZOruqql6cvynOsk7eKlSVMbgq83UYEe8IONvGwOReZv
Ep5iAG2lMdAQl1xJmvTxVFxSlaNlgyhjgqd6e3arR3kbu8MlvwMknVRpmBDVnQ7P0Qfb7N3dS5tO
MSZIoqI0oGxGJtvswjUcf5dy5VbWb3tMAuViRc/ROechRncc43s/Fdp9E9fKlLZ9w7ZAW+30nF/9
tbzWT8lZEoM6i1XGBk4+j/YuGCawLGocbNuIL+37w+16pWcJy/KZykFEQN227lX4oSVzBBioT1ey
mfi2QELBdqjbeVpLy8uZu89Ov/kAUNTSw2f4BVqpQ2ctwiOe8fqYGPYYtZ0XfCga9oJMw9KpPWL+
/YzMDmlGeyv+rfJ2D707LSmog4s10VfnS0Kv4QvdvKnrDrwCyiDko37IcqUNxqa2p0xvJmg+hzKo
6a+bv2bX7IibgaQQBdpXpBj6yeMTukRbfwTA/Yx36aJIw2AtUag0piUJDtW/Aa2T+XaPkuLzPuZB
lcL4SWv/ale/K4V3+x9OT9d9Cn+N7R3KOwo1kvudN0KyNnMz3YtB1Ml6gz3lYUI1rFM0keBi1+ob
TnxgMZe9j3bmY2PMUuTYattI7S27kZ8yE3wjC+oUGFvQT2p7vYDOpS0qXB+sZIZn9QVMqkk+jXFL
ZgEqaWy7cgJtvxyJFobPvQXySo2MCTuOuY2krKKJmbSnkz2DlXgjMIXpemgvgegaBdFZqWPAreLN
d/AXsK0Bxm0ZXQqg/2vGjFDJkchzHZBsKmXyqYt4vQSOHyTEFJ1g0RwKPd2xAz7Ob+Vk6uZaZS+u
lsPitAAKL5NLpg1RzTgWWUH4EEwq+ftO2CXKNiNeXDfsBcac3Z+f8v2NlAwisbVuT0+YrOwWwqMo
CEwpkcQT/yNMfgAs7ItvX0tQViPZlpTzPvhPV4rvJu3ID2s7I4KS7Ht1lbCzum5f1GH4vxMqvnhW
qmAcJ9dbGdpOrnA0iWS+Z6bmnuLK/+E9AxRiPnpYbMycYfpfP1hfwNVxG10nTUscmRAqjuXQQOot
efe5Ye1ubMLROXhRMRhMyp/8NwZ1NkCp19dQ/ngo88XHMwoeQ55hDP+NC7DefzdHu1HWG2xZhan2
Kf0EBDJwSyidhB6B9MGTU7N8x/uR3lCGNXzGwGu8ibiJ7hsKXRn7cz4Z05141EANLF6u/XeSTsh7
91HJTlD4IX9B3QB94NQgI6P08FRjckN/0YBCdJ0xXP9edbS4QT2YnzoVs+76t+JhbfbUTAbfAe4s
k1/pNFWwRJnYk/u1R7CgFk28Yq2HqX5EICUBXc7O0adUVz3d1Yuo/yugIVzN5Fq6en4XXXEOco3Z
cT/09wVqU20Gd9dPyJ7neMWIONhuFjf9J3v3l3CyAgPL0g+zbIR76hlKTVcchoEr/3XyFgMWiiHP
9f+0hOFesXCaMGQJ0SoqRsB9mp+rhyGPBSZ+Cq4YXDYWJ1rvLTrSb+B1MjEwAMgQRELTXZocyqF/
0v4d+RVWiiMFOlBwnrYw7lD9L9bYn+MOB9/taei0QqkwM/ZNi72I8A6S7sBO4oPz0FdmxWzjN73L
qhtT3c/TRukmhGCL+2OaGF7WHF4Xf509C0m1Y1YJqSe5JOFi+T+DBf+E80GxfFybVd90KhgLn4wm
CnBeQ2T6rPPskwgJ9ImQGwutZr+acL3cHRsUQpAfF1AnxxxF9+C340gkhOK5yf1Mt+oNMUO3l5zR
By0O2mAi4J4wTU0jGJk8CH2L0DNBIYBou5e7sV/eym+om9x5I7Q5x5NswIsKnnEUXtJL23gpKkhY
uPkXhk7DA49B1M4pyTAEeEsTxksuTkiFycsFArcEH0OLZgRtf8thWWLkHKj12uuT/imIYHOakG5F
sgVOJbtvCZiFL/WmGD4dlRQGG+Cn8lH8nwM/uGIyKrUOGc15SHGwYEwRZV5ybHCyqFDycA6JeNWs
GUfa+T8LjEu5ZH0JB7lIRXr2ml+RkWJfppuisDLiEL/LihraFGSKyO5b39L8MiX7z1fC7Uhlje3L
6D89kdiSKF6Af73x/19hYgVuYeZHFwoslhOJnFM/HSpaayqN9+ZZRK8YnHyY9SWyN604FxZdCchx
xWuFWEiSUyvs/lkdlOXPVs4yfMRPOibXNCRujodPBSMq026sxnfb4hOkQhZGq7UQlUe91H4V7nJk
cF/etLn+zC0cOD1vOBJIPeRgxxa4dKrhcnMSYfp7YoSSUB+KWtIOg0vYXq8zS48LpfZ2LoS0Etv+
eG0WfdYjT3lu21T6IRZxI4AdF7t0azO1pHCMTdpRXMGnO1ZLF4OnTvaRj26YgcL2ozZtDjnX8e+M
3mbazEEn2oDCNRHSf7+LW7Xh973DNO99/dhC8whlrh41wV18WhlztTrfA9S+ETTvMVjz1WV/djCF
WMZQmAFDNBSrFfg6BDB5PwBOVd1uQ5AKZkJuWDJlfVfD3rsge16UxLW3S37KIoTbl37SqU8U6QVU
3yc8oBbvz1XjMML+L2PVeS0XzS1ESIOFCZhUP9g2oWWZnF5crEHBERMdJwJjN2QmloZsc/0P8dDl
cZdNb25G2oL42Itn721cCLkbM36C6VQpYoIuKh7X8WnWQ4mXyy2+ot2I3pUWIQ2bwjhhd1RWVjYA
v6dLYyDIQdL6akGHS1Xf8m0h7iysaXzhxNzPKW/v2WrwGUKuKbnjY3YCwDC4TaC8W6WVx9Ka/mGQ
I6OCCRjkNhOHzpKIeT9cJSaK3y4A9yKJYokc5bpChJQGUGVqpRJjlQS4pVHEcPTO1QPfNiHPGS2n
UU0MDFlCBtESHa29GnIGS+SX9WitmqqkRxNY7RaSCFAFd6t1axURCtNalzOMhH8jO66oGg5ZnMts
qhLhCq2VMQOJtAvFmB99s954k78y3Teu2X6W05EpgGoGzj03MFQp4ZuejOUd7nY1E+Ad1nEvyTWa
ewWNv/74R4I9YtS7ipmiVymFgKOuQI6ZXUryLqvreeZP2aMjwT2movKZCValAEVW1qDTm6/yd3Wa
bDTZuE2tAZz1U3nPb9jlmOMBF7yxzG5Jm4YAhBGlZwBTCsYhtXAZ0cXLj2nZH7/VkRfgY69aj1Pg
4rSJnOBR0bk+6mxIMPGLqEzLzYyCH2kDN9ipry56vjectiW74efp6wy8gyBYA4onO9ux+029o+iC
TgtlCxm2fhxAfzxGwqET3gb2HA4HSLSqCZmohBo7gJaccw5l0wNkI8pI+FRjSLhsmu62gH9F9kNS
WU0dxk+sXeb2O8AYmNwO5sEilrRotO7AVBR/v0gdJB7RBrOecJZ05hX73Dr3FaMZl03bgsp5z24x
pzIpwjhJpHtHnkXy0oW7yuzc6SFlGu9V/dr80wBcqIwvnHHKmFxvhL+9Iy6zOFwbt0pf6c6R82ME
E3Ty1NGMnWtc+IgLHgJ1DRYgmHdcaeEy8lg9Ytrg65qK3CjNrg+xv/AG4HsP5d7VIo9OgwYW+Ha4
teHRzuTJ50wJnYjdlVHwNDNpOqyGzf6as6asshYkfi0LurHJHlFU4hkMfcay/Ye/PEIVu4kevf05
Z7NAFwgIgdBI4Ag8B7gFkmoR+544yru8lf9j7S5wE/vewKZ4uRaddR+nXlEBhB4+8dJyunki+BP9
+ZYU2F2m3do6LwIp/QsNJoapL7gl1BXaO5v2toKVWMhjt6d67uUbzHlFstoFDED4TIvjN7A9hJQ2
cSpfmNVVtI2QtSr4a2E53zT4l9M5COU46/tLLD0gq1zFrxF+zo4ZM7gI+Ys4k5PbU/Ep0mQ/DXUc
FGKmDBLZKxIkxuoS4X00kSUnnkrhINMuYE7qwLGG93PogWdbPzmUvB9dO9TXVu75+EOsgBoiEHwq
jiMKCFs8e+qNQ1btaPWJ3rkrbY/6wWihBgKLa/4vDo3/70qxsXCe4nRGfSUTB7482IQ+b+Q7+mHv
yrBorz1Bu4cfYzn77f9wm7omiXGRly6jq9RgJ0CgBH5HIkmgoMTj3tRnfISYdxsmb59Pr+3QgsV6
z0WsHzEh0SVxadNp74+YmPcQ79uW9NMAnjqgq9Az/hYmGeVhYUNtH+4QelwnZ1YyemARhvzzUR+G
CSgdupoxec1NnvT70rZvFXSR6JGuGdrx+EX4CeNKYikos8yU4XRF2pDX8+RdC4n4B21CrsGzYxyP
jgUHi56sHmS9SPl005nyikMcwFskuxyIvmZttOUig9BSI0jljx/kIrs3MxYZEJ8EgwQ3qGwS7Qnp
LQ8mC+TnvvwfGUUDdqWoSUAEVQUo0hHEl7otAqqdspWkv00orZoRfsRmzbeB7Y2DITI4tjatc+9J
khrc3czL1qomtzNHDupkPm9kBXoRYc/OJ5d9JOnc9HS03wVgNqCBVa4pGmi5yVfn5puR5aejTTor
4IVVG2IeDAnNhLWTOgGG+Q5TQJ3Y+BL4yeuaq9Jam5q3F85bZqUjEiQ99nyQ9ZY6ly2x7l8Q6y1k
ZYYp9/XiE3PviaEfIAMxjq3L+nB6Q9kS5ZqrGgD1faGh2XBQ5l8Ez9pOfp5J+rEdhEBWg31qPd0g
FgjZaGdRKXtwi8HRBYlB6gmEO0XeLZwJlfPl2V4XPOjl/a/bVqSp1DBXiIshNkSs5j8kAMBUW03E
M1dFSOV7Yl1lrupDnTZEWHlTB1X18CpTuUhFYR/ZEuhXaIh9dfsdGmbrs5wp4XMo+ktpwMCmjC5i
Q7aTvRcDWJ2ikYw8JjNJ09KGAXWXCmraG8a7uq9Q8DOi583xPuWctD76WL4cFWrqQyZ2P9YhCE0W
vsPYMVrtZ/Lstz/rVUpMIZkle+PFmYCmYok8AUdhFsapQnzaQ9QzzWoO7BAPMpef5ERRYHpQ4lbS
B/4yo2/uKG1JedcIxHZFgRqzLp7DnmSIkKtuwnK6IFbbX7NA7n7ifJ6XIhEhWcI+pMy1oJTMoSBr
T3j2bR4r/Rc3qGmnVVrbDZS3wpblWNrPF4ZJ94dWxkM4pVyEaS/YRiYp8JjdXX3WgSDp4bPy2vLZ
G1wgbk1lP7hwY9pXiIaM71kDh+jBJqB9hDW7ModP6Qgr3nNd5DtfDoSwpgrjndSJ+btL7XJYvQhf
R/ezoZHtCXis9YE8tiOboziMvk0ZbzaZ8ac+c2j0J+hzTlWV8ySa+FopFbtMVMl/WqunRB6jExRP
9oSN4cr+teyLkF6S9YjpDxq7YeWb4TIrJhuiwefng6aRFyueJU2WaDCdWBgt++WCSs6SaiATAEQP
the4sxUfQ4zVsLlZtRHzvNqF7borD4MGPSC8LQuB2wnJ7pME3QEkjPhrMh3z0igAE5lxuH42DchX
9BOuEzHyCP0+jrzvAFvb5BWodpqAZNZsDw6q/4zcAnW2MckUcQqn3PVODiErF0dFEcbZESsmomzC
7NF8Q/eQLRweolXIK4Lvu89LZH6OLMV4ZIUakCuYf7ffGzhs9BXTQIsyquc6cxnNLEfRDTQ4buC0
UzyDbF9uugig3WNL67aCFmDO4pFQ2cVBhdlbBBd0t+pEjHd2aHA9EU3pYUkBrI0JhB7i2Apeu+06
Y4+125rw5FcMyNCaF+vIltJ+ZC0zCywxHpqeBB2FmldHtOtsl43f2zbg4GBy+7G1o/neb/wL37gX
9/ICAwW139mDUex6Gmgy51xqIiflyHKq3PnS3W0dO9Se0Iu55xTYG3grV67Pulu3Ac6TQNCICuEX
lD+H6Ia+MEWtvsU1BQXi1lo2V41K9IUbARAuCNBABZAaCfj1Kk/gxWEmcZAFJoVDfOJ8HQMZGwlp
DtjBaBcCQZIKoLu5wBwJlXNkDTPd8QqbLfHprHvJAgYoMlVSA+frEhLFmJwLeLa0iVXvjInVNvjk
kXs6CL++e4tFukqc5M5d4SSn6Xtf/sZkYIsgsIPSX4mcji8eVHTWeY8wZMm79JNnRfiad87vtYTL
K3fny/m8BUmbpzQeev4SC1dN9MaQklSu+Etxr/ZmpfyIBIE8Wjix6tXfjowufAvIzoRqGHkD35Rd
ENxTQhCyeTIuHuyBFYQXg1PT0VF9vlABFPF3xNl2zDk+ie9F30XjZ1cJB1qvjEZbF2TC5uCyZixw
KGsf7Q9BW60DQPsPtoOBVYW6CPdA+omMr529FEiQ8pEGqNLVv3vsO2K9hXU7JqPn4gYuVkp/8yPp
hiCv8X7nnGUt+gW489JhKhenAclQWXSGMxFogci4faS+ELTaNBcSH+HHAOk9QZ7q0g6a2uEH2ix3
o2/RBBg0xfDYFBKyG2n9fBtxS50EI3jLxLh7ZujJZT/pWZneSpAx5Cg1gq9Fhzloy8uLojMD80VJ
jgTlG+03DqyC3MAc1B7Ab45AsH6eEUKkIlF6eLvhXI02evxATKXlbbBVEPL3AHR0WDcclQ6GMMsE
TqqVculYCOxBiShTIdcZWDqM0r5nxWdbFEMf6dzYvcpXass2sk6gZweSxfWaSLXB0IMyoH63rOiT
+E66EJfIFtCvmyMu1dLghaMyuv4VNsyJo6qY7S1R0MBNdw8zeOcS7hSV+Sokwp90D+43vatgjG7O
7U3bVqsOVplsuT1lRTiNvVl0563F8eKli6lYOLgLG5BheGrYsg66/CGfJDuRiIOHPKEmszth2gwv
Jdk8pTIWY6UkK0cqdVXjEqyXU3NI52SsV+kbASmsWt0JdT4SHC3O+shlu0St5K5+W0eb9tNXV8CT
5O1l8LswPZhvF48Y8jA00gOyB203b13vN6lRPk5X+f82wwgapsdG8vE+RfqK7m6zjv8tqtx2pBGy
D11ciWVz4B26yZsTA9UKJxBwRKrW2gos1feCmtSOXuYd+iC9O8hZROEHXqjG/xMDToGqX9CbkpIu
vFUz+A+dDo7uHlcELaVa0+OYgLp9gk0fegZx6jQlN58thVv5IVbLf/ZHljeyVRHe+t/gn5PhJUfe
yHnGmk3R4MAmgMlBUxUpcAWn+Scfvbd2OuS5pVXUUP2iqqvrBRayUaaJrchTuKiFAZ3nX1Fy/hPJ
SCde5z7DND4T81XsVrlPSI3XVhh0C42VIyGgrfCm2UANZ4CH7XIlyy3hjhxZdacZa5aCPJVY4bLu
VIebpgfvg3kV77mx6hixq8Htsju6L+TeoZBfMJgWOWoAb63NT6QHI1vXS2/suYVIjkNAXMcpFbAK
FAkPlkuCVOUtFe96iB9+qL6A7DTP+H5JXmzASf0Bn0fUP7ic3MLZuwYUEUZaKxwpFAYT6EEDEjt3
sxIs4TyUwj8Y8mnyBtY1iK8AQeZM67VRJdnXTsBOQ4U2EXPLcfdZ2yGOzuCtch33Ga/R74ltzx/e
GudVDoDebtwEwlezV15dQXfFzWHKvQZ+XeMzPffXn6ykgD8ZhIFv1MHv5g4QRMQe8ftr61hGTZ8Q
4bL44xJAekhkHy0L+OZFqjpZFY+7nBiCGD9Ggi65hPS1c8QiWpigPt4D/uoacEL2R5lH0DbB95Dl
ubZajg9Uz/R/UkB6ogrZPfnwhN7SYcgkB/KeBmE0aML1RTEkP9Zkl05wfzpfFUU1A2a3kJ7gd7xB
sGk5n42UAzCHXV1C6nsTCzbXs0txNTHVFJYKiBopQiSUACZxPlygMs/I95NE8qsUWrJbJRSAs8E/
uANsYfFHgNpbdfb5UNWaH+p9y4SX8bKNpx3tZ2D5+YUs655WdUzYcITgJuK9qtTDzPgrfNkHWmdX
Qa7oxvmx8fWcdtKxte1xoE18HwtVRYRzREE+c77h/Dw4lHr760Gkmk+AqwjFduNwJ2xYjSkUhtWc
vZUhvFTZevJk/u+d3gO1UBgZhPjVQePDLFRA/bQ22qGg6XH6pThxoRSGXiEwjLBA9JN3gpCuQe1G
kV6eTtyyUoOCbxIjmgpWzXgT4A2L+Q4QYgOqP1BRG6sAuWCd/3mwCLVaEFLqWtC83Trqw1s3U9cD
Vv2GteJCG2x0D/xJHjiSCGbKj9dIo865nkYNZ5O+zvwGcj8V8w/QwQVmjYBgHtdGa5fEe2KEvund
WOT7envSKXrs5L2Y/plTmiBfM51JNZ8mvKTv2vSZCvLptoh2KnBXNN1mSwWD3uL4HlNAMkH2PpH3
jXtjbmyG+32mCDjPiZBhYAf3aZFHPbVFpFVjppZeme357f/iPKpJSc5NzGDMWBpCW2jnZ9LQ5IHj
qoPBUbYD4OMs9vCynTRjuD0AERtAvd8CDq0pcjiyG+z3FnPkUTMJtUM2GuYUmRKC9MHXXXRVEh94
bp3/olJ980bEmkDV4LjYKBmBt/2qZXsy2ytNO+4tEW860UXsRHFFN34VDP7eOR57WeRPGINvr7m2
SH022VCw40bVCPZxTIEm1D8EmTFA6OemzoiATtjbbxnXCSUmmoRg/r+kZemnHA0m+3Vgkfoou4Qo
TvJyjzkqA8zvNkugwhEfPBnqEfdclYIFD0Yc34wIkMUgdR6AadcS9d2g/LCRyZ+pQ1gQ2g6fS+8U
8nsF2YursBdq/dpKJIEfeOQ+pk/O3h+Z2YyOuJh7hIEqjhm/3dEnHs+rvF0CXnVbXO7Zr9JsSIv1
D5qyOEf/neg2IyEdk02fM1sv8CS/g1OYeTME+4n88sXjiBQ5MUgP2FRQ7ACPbLLwHIFBtuuF199Z
m2czfA2wO16QAU26ttLnnsuCYAhfXrRvgKU5DDzup7BC9K99ARfoybEjbUi0nryzf8gzFLIUj6GM
5qMlam2f1O3zu1DRdgtVSU/crPZA7h9ydxCFTqu6B0SGv9xf56ecuqXGW7uRykUyN3lVFZjITt6U
z6HHziWrmc/icprTjgeIiwwVYS0McvLfzn+/5lfd57lWuGbGWHy07rH9gJ8dCH24E2HdI4TK/QVE
IOgHW2miJu7UB5i7mO4KemzZ0Y25Y+Wk4A0b4962vXRaWXuo/P7zk5va5feuA+Py2G89qCa/pLH3
zPk/vSjykbuVNDwsk/Gru29B60CK/W85LnRED+WDELIZWRXSJJE1KU2gvKwlAyg5ZLOPzOmymQ54
xbJbXnLN0z/3ljk9Uqe+zd6sK8Bn1X6EieNoGeBPiw3TZo2xBy1tFJFScPUHqk6alqJxBPtSDx++
ADf8HcqGtecIQkE1ecVD/NSiBovgUB5nNaC/9S72ejLmoL5x/H//ODQTyc4u8kCILLY0Oa/mOc5r
F7BCGy4GMQMyrI5AnLBbWx2zkS8eumuFPWqJd2m2uhyvGwiJUikeF/wo9+UsWlwd4SSCXJz9ApAa
VLXycbvODSycKF5VpFuss7mcFi1C1HkjevHry3CE6yVYhxCBlpMo50catJ9MAUMvOHCHu4qlGNpT
C7ER4rmsWEX4hEL5LV+nD9n+hOnZTCyR6fbmelI6ly1rHZ9/yZoFlkuInCr7+APGZFjrqRZOCr6U
brR7VM8Dzoa1nr215gSCTqygW7dQMkjcu7wQezxkuehoKMx7JS0ZZi6MqRdGiCSyVPptP61xi92e
SNwSwlbmXVuvYKEqoA4i4cxSJcxR/W9zkGrbDf/K7G9QJkMDHKIPAN6efN8Eb4Y+wwrIzeG8NrTx
xZd6bmGuRzsRaoV/yNeE+/H8Wqe6a0TPYg9pUiMvz/EOJxNaTkAUJPb6E+emewbmWtxi+40RDtBl
C61wy5xbeR7+YLmBK77+Qn+6iRs/hUZ8uywtBWLmQXMgyv1gMolnfxDr4pBRL0jOBra9xPO+Vunq
mSIfJVpz2c1xkeG1xW/AcSkNbVS8SN+N3QV0OAx/JX9qk4U4wIyCg+YwQSlNQMttM31fXfCgZibh
MBB8G0Z9KSc3pwnU5ZHAShjyv9PbfM7MumjtUPChykJ0w/qpK1FBQ5tqQgaHZYqDHCndoePfBcE/
sHsf9Xlnp2hb+oL1flbch8J5cSeU0L10ry9iNAi764v0xoobSMItVEWg4BkXjFWBGNvwmgvJ9qU5
ouXG0qSssLHwVe9ZzAM1wNpUdbnDErtWtsEu+axEcNSd3LF/cHBUHohFp5rze159qCRDwMu9k4uv
mzq7ImEaLzXvFVww75TuRWZ4lz6t/5f4yULAGiKFTxBgZUHCgO2Fi3twC7nuPh19HOjqeHKClqaE
LAX6NxzJfkSglIpMg9S7oxT0PH2CbigWoMIsE1z3dPaE28Hh48K0k0ypQFDBeI/oTwHGSClWucAD
jTXLQvdq47KJZ5N7IobhZ1ajRuJ5K7wCo4+r/bS2gcMBDnr5csh6WCmfuaxm7ULyGADfYS5l4/Ib
m9MpTLgHFt97xLzWKp5/iQq6rUgGIVc3TkPhg8Cua+RPDsi4+5FUMkVhmcL946CSMPzSOajBDt/Y
f57bipwn9k+ZfpiS2PqmWcQ6Syv9uApvmC2HqWFiaShRo+qOvp8YzF2nWv3Mhy7SR7fzmPNapoEb
lIiwos0HOx39LgBoBl3WZQYS4R0wRw1cNjuA8tHVs18JxY6iL+gG8bvpdKHXs7euYU/MPCY/GoOa
DhKXTb01xfBwy2C7523PSRjzUUjqIr5xgKBBQ0kXKG+3+P6DQ+t5qgT/HSNVtAl0LhK1APNE5j78
WK9UM/qEMUMTQGfFXWl7vvRCQ4TeoE6ejtqMqpQ71F84VxTzXsKx3Gxj5MzpGroCjdGsic2cquBg
UmVTi268Pimfsf9ft5i0l/Mjofyp3/3nrsiS1qaGh9MsZ3a0BawkenDRDPNqGebE83qJUISzlxDV
ucYkQT702WdWVUeIR1QRqKpaGQhfCNRx1WV+tNUK2o99toMjKEHyOkgSkEIDVmdj6SgNQ7TKlPqv
U7Vwx4DhI0Xeh0YR9xbHJnn8xQCyD9+TS25qun1YF8JCEaHrsqbiCZbWC6FQ03pia5gNwuts6bPq
7L8gGG5D0y+APWdMzfaoz1wShosfVOumKsDvBgbIdQmJK24lyrlxeNldyX7rzm6gHwn6uK8Nm4F6
AnDcSg0MzlWKyxW7D7VPqbaLlB9eec2wTXnG8zCMYYuOlupwXZnoWhUPckoNZbF0unxjltoQJX7K
YhdDALcr5d4LO9JB5kn85Rw8h7tv6aSUtM6cUuCFSMJXaHtg2+JwTqUk2HjHdQT7eX++xQNoPlyZ
F6+ucDMvksPFdJyf3DL3njeVuY1IKkerHqqOl0QdgA2seB26Umx9doqxVg+itAT3f98Kb1DfFdaT
+roxFcFjyAkPUGFDPwEG2PdtP7lpJT+WBcBctDF8rpzY+1I51FV9MEjh5+KFAwRSzprp6UKjD5z5
hyF/YTNxeXYcJmn1UWxxclCG6mDd2/oCvXM4QosoM3h9zSg1s5YU+hQX2KbBZoYyPVV6EMeZ5pjn
PYmeUleCnR0JV81X5kUQMO3RMYasi9nfwdu7delK1aqRuIQ1rfz7zdqgA83X7E5jtMFL5Y/0jWUd
BJgnEqN30XFdh3hC73/cbu3QGT2DSbzPnW6+l2ulHs9ExSDvByDlJMXHviI+QOao1Ot7tmy3pKDq
EkxJm5GYQYKzFaSNCRfo22QERFPYfQJd68hpFW+j3E5+rsNOJ+wo9fnFn0284VpEZ03854RkOZeg
CVXsibRsbc12FfZ+/sbNLMW9mh34+0MFY64IV3DGgXxA/VWR0sEzBhnwlPfaewMS26FfAGYJHsHX
JumD9wdStxRrahYhCipMuBvNTuOfTsMykKZ44+Pdfoqh23bSkMLxY01s2qjzQeGKDuU2FmGupxT2
feMmw8CVrjrMIMRCLDV4upbQsMSyoRfFkxOVUSlr+lwvLKd5T4gVsMh4JPj9xDirzJLf7hgSKcZj
wKGtFeYgTHun0EsYso/hTRNGMobA/F4NEdLXs40/LC5RlkWPwbVuQkIWoiXEzaZgIXrG2bL7srUw
aEl+kllz91d13XO+qGhMzv/xkilJpS+yguLLyVHkYAQXzmRHrCMF3hUi7n+xZPstv4xnrNuuqizN
sWFR1k8dyqLwr89VYP00GfELFRie0zqDGuus07TBx0QeHdGo3ZEDP6YQhNEnkdxFO4oCHEClpYvM
LxVesSbrND5vyUhGN2zk6OtDuiPJIUgS/+HieqCETOqZ2tlkP1CDa5W75RjTenKtVv6yrNr/N/6W
hLO9YtFhjEHmfTAjUJfoTJTLuGCMzXVQr1XCHMBj3ozhzkaf/ZeG4Ucimcv+oxmgQThINQ1Rt3+7
tj6gox3EqxyUnaTtD98bSqX4zLyUmxM/Quyd/0YIinmZO9krJeo3S8+JrJcDpTXjLbK7xM8KkZFy
oDSWqgKqDdslStM3fLz6O6V2TE4StkQDwNytBGxaaPUUMdqDTuuWtD+IC3IMzOLQazRgA3uTeXkN
8GMQ377gTJbwd1RBQ10gE9tpRGx3UVlyYJ3hR/MfFvrdyzvkIg3iHkGCB31EhHyGyIwMP9lyiEWd
Ii6oRnl0fiWv5qeJ6Hz8B/4+aXsv6o0kP+Ql4Do8Gx4pS1iyMKZp3ZcJkW5CLJyoqjnmx9/NlLjO
jMthFOaRtDQI7gp2NOh7eoUdVSj9In6u90KV4YOjx+PMOfgxBHibeYI1qkdG1uxxQSLdyehdiHY4
j6hnthZaKnuE54mJYNoKfiOaOTNYCu7m80HD8dv8fb5YtpbIH9ZBzjbLjwcmOCiopO1lVZSYXQB0
fu5Ijc9Tnmi0Retml70vPoMKVmIVx9qKXmCq9Rz2LiqHTpZ9NlEkPTsGLv5KfJ7OTQ0/Z6UbkT3y
TuiMF08cDslFNWzJp+LMqhd8/OPnfCoOPdWy4z56TLa/ZR98lHYTxC79mXSMaTBe7XPv1KVbIE8B
hLf0yzwEa1+GErgN+krRvjdIsRpZrPzDCaDLnwRJ9ocVJrkTkQ96y+cI/+2ZcmPZd0KNLXspZXz+
S/5KiKv92ufS4U7pnBpZ1vLoayVSNxwv0JSZVaVx0Z0MbQj02ohHBt8+mEqbKYaWf2FOCD+FbD2h
OqCmPmd9MN/HK0/OUQMx/WSf/o9VBDujlrLgoEekR2S9X02g9/Oh+RzTJ26dEgF95dj80tZyLBFg
aPVZER+VSywN1Xsc1ZrSvAZLmW6+hbiqepgwtDKONtRx/NIhvD+K73rqAvDAIIorTrwy59fac03C
B9hIH6yCD4di0ecBykGy4Aoo3ttJ567L3GKG7eiKoohjB0Y5CpIO5VldAswjtpyGvIDMAeS/tWBs
zVJr+hgD3Cb4YpWu5jz9+vbj7brAbfSxDKsb9+OL4DYt4toeEb8uF0+B5uldz70A+4ZeFqD+S0Fk
1+ew3t13TUwu1ViPsUwR6iFILsCrL2M26j/AenRDXIKAUmUf2B5PwR8XPFfeskuIIcyAoyFmI0VU
YgrX+znKwJuqvmu6RPWWuqSsSnTXyG/Mme/RuVcnY9PP2NLPOyeQYGZWfnJqgJsOCqzEIZE9/Vff
Z/5n/cQFM8rIyLSHanMZIcR53X9uS5SH+rcVcyK5sRSVcxYAWRZgc184+eyeZuLR+NHMsqgbeXwC
gY34XgtJAN4lJbnSsFdu5PXJbcvxTCrPhQgKPCmiFpA70b/K/iz0e1BFBM6+GD0HbZ6y36++hOWI
NrjtjusihCtIo5gazLGwLlnzQGj8zgNGULnGGGiqMd3aiNCzJB594Ul33/q+P5rQvuTY/SdN5Hzz
GN7WSNU2C70Y1swQWj5vj7COz66ifDkfTg+pBYoN4v1yo6BK51Y2meMVtZXEEqc9r26VM9pJ3QKr
fXyQSgLOcvOMzjUGiHoPCZdXuXvipmZd4DLPEEHx9viWGLpzqFJJa77UTMoekIFD9cW6ozclDm1F
2rFhJIgoTYgpceVdyeWczl+KFXQb508EeZdYsPtEKwgM9ptLo6NR/Sa2pwgPNYs+CINVb5Urit5D
jWjzyni1pVVt2g0TrREKipBD76M4qnTXMy8mwprrWWW7KQ5bntdJl6BbJDXjihFRJb2Cy+7OthVX
yQ14kBLUEpE+EVDLCgCtzT1nz5jp+1hRIfslG5zkAuA/4mgOzyXmJB3aO3DYgGTxxZPcZvmX8OW+
oqiHqgM3Makp23SNY8XQUjQNn95OLKDcKRRH7CZZKiWaICAmGfKd90XPbZHM8bmSu7+w5z0EbVGX
xLHZLMbst+v+7M0TpmdA70HwIdgh7J/D2ooEU6MPg0MGqsFC7h5oz+9QTHlTz5yDLZ7uYHC4V+gE
ueRilgA4vl26KS1nwoAaNWcNtPtZpN/YeqCr9CuoyM7OJt993ec04IWxAkuKWdRN9OxLEp9FXHhz
UEYv/ocEyDKUWrStecFywkG5d9YIBO1Xj9zcssBLXd7dfPeJjn4B+6ow8k3J8HKZ5eyWbqpU5SLk
/47SMSbIPK9w88anpNzlhrr1/UZCEkVaEnwcHFvtyGAWFQMH0dd9FElMyQ9BVtjNX34+zd5yjJA7
mdyyBA0Xe9PX1Cj8zQC4cVYqxg8o8PP/GUHS0kqzvlsywR2SBNMNC4wSBKToGsj+JkB+2ETkymBW
e8nXXblF+1rnbyeszjsqBPdejVsOzS9CMt4Rrg2kPgKMdly43mPdwscRxSt3YF25vHnpjyH33ncL
dGeKjrm2Z6VfJ4iY1tiI2DJSeVoD8TO0Q2g1AqwcDnpjpWwwiTTZV9yoxHpKmTcXkJm7laCaFjrC
zEdFRNSndVzEl8yFXjahn2xWEp0XcEWg1v4cU1/xkJzOQYTDhBX1zSpmAZ9lEgNa+d+/NnJcgcNJ
SzzpeYeD+WPEUqoA/mn0QgchqcUoadnCeP6A0vWXcUZ1EKlyX/UsQsl+aC25HK5DhJjL9Rgh9KhW
mcjKb2IEuj694mqxt0/5U51xHmDl37zBUD729O92dqsVsfX7uBvk+DCifLsOel3LkDIJZkOLIpnP
QBha8gAikt57BjZJE9dQdKMf0yWeG+ttKZqpysWi9DYsMiqRT1zqymKc6vHXpOARr01kbXIL2vhc
fFGK+O6jkkL7a33opQ8mjR8Rm2dNv0HogPCpnTGzspKAWSJ+qsJuSLvcJMJZGUA973Ujzn4of7TX
o3fN5q2hE1GK0ZXl4lYh0Er8d9NSjMNW+ManTpX29qKVV9pzcesDKwksBUj6ojmwsNbLakKkaXMY
PK/TNCU0a3bYhqgsCoCBc3q9rZU2lj/X1jk+PpleAb94XwHi/Q4OV4QC54v/vzXSNF0KYwjkTUbp
tmnDYnYNEmAa8pskEtrJBR5TUIjKZVApFL115y4Zavnpc8jgFCb5nib50bw/deaAWzTczjTSHjhl
+nG7Wn/tlDbuUkbykEGVTYeLz5P6D6ssYs2exD4vcZ4JXnBUZkMrCA9ZlkXQMbSRYVENmsLjbqhA
L3u1MvjvIoLRqZuXEv7WgNZndlNOd+8X5dQCxSqwGHBUHeYQehkb0XcZb2UdKfT0hKQVjFjyYlbl
4mFuU+Y9dklRvIawfzfFvoJAqU/atv6ENZQRkUXK4MuldwfoDB6HPtNgZPOdyNIbqpxl35kBkyJQ
APWKESOz5T3Q8quZxEpar039G2UVP6JuDm0K3+U4tt3EAyuyu9SAAZAoKGflBPJUbPPmA2KfPlA6
NnvnTBdelt2uim5z7gY1LPi4MCbgP0CzPCPUutGqwziPbwFI5mYWztAtG8Yo5xtvITv2uqtmZ6J1
d4Flek8AqqzYrCs2B5LbIArS4+8t2Hb3K+wqFzEtsy87BKt5HBaJIpR6xjqq0QF0oaT0Q05ahSfp
3kbW+4sMlhaB1+I8+/18yjT71AlaxwAtjD2y1DczUBLqqCspkPLjcvfcqC6AdRARqPdbgd+fWdQF
Tj4PlZfJNx4Isj22/6vtVhzbAFYgptBYx2lgRV6EPIphaDjYRyo2l//av8roEHRyZgVjyj08EX6t
I9vFcumWc8xNSymG5htYYf3UWu5a9Y3eQ8JCANSWQ0BlpT28oGJ0lSDQKEhoNYIbPrU+Xq09ToZd
97H06f2J8Y8s5CeatdfcqQOckpmAUf8wNhAJl86Ansa2wiBx+79wJs/c2dQ1A72gWYfBplUrWOet
ja1z89P1iyCwOCxj6u3RXjsLTSUswkJr4jDLgXPweOtGP+73LuLgPqN71R6DMlUzXAndEB+U6mxk
WnnRdqlURuf2GeQ8xKhDHboBqLa1S9ssSvUZbByf8VP9ogOXUykvlfF4KBvoj/N79bkR/rD30Sr2
R88rIxQN/5XyzRCQRkPG8SHY7xrsywvBSBfrxEf4pbeEF6lVytkbRuaOmGnMV5VMDNwXPAUPQqh4
3Sl9+clwGpRVIpmPHucWEiYpRvKqWAIZquguvQFMwvGXgHJQizZVLecczvrF08Zj749OEWkJkwdW
T+Br0EHnM9Ge4eYoOqZHnr0Ig1YwLgpWsav8qnGpBqr74nTQWmiI5GxqCFlD60h2JgXpFWtLUnBu
/GJRnqWrI/kTLYfVIldyJAfZZsd1SAFY9ROmlYicbUYfazGRqDJ+UewT5EWXgM4qHuf4Rk0YYdOi
e3KX0gGZ6gHbW8rwXTnmNqPC7yueVgCPbEYIMhkqRpSNFlWKS7cC0wKv3ZFYe9ByFsxqN/qatiMo
WcEfmQ3NP6JtsD+dZBW9ajjXLcGz5EMHk9/Q+2+gwQ5C+HPuD89VfGJEV3jTcAUTjJoG2BTaUw2G
hXwhW9QJGLTPUaiIu2DP02OC/ySmels8Tw9CR8UGgNZMCRzxpR1TLKOM1H4+drlj+y5efxFUhvnV
e9g4TvtBIK1qPH3X/S4RVm9+5+moBoglbdo0cmC358w/viyIN5Pmp9LDLCP0JSI/9e0iEIrxHE9E
xXaPiKyJgGPnI64zIlfYqJRmv4889u7MdXk4LYqonsuh7NpoVqxbFwGnyb4bSOWXN4e645fcUt9R
YeNtPAy/AbWAUcRQ7XVWjej+uun1WGp6OWI2llFTexCWugVPyMThk5QCq7q1LUWttZ+jGS7eDbOB
B34i2U/FHpp1ZKS5cUFURxirN3GCL2xRi5W4hjy91N51UNZ/q1SS10MH5o6SGOMFT5jpGg60ZlYE
nfXe2N/3VsACbxqW0o9deoFBKjbQzCOuOHDdxMMiEehrPv067hsG7es6SiymztHgkj9rBIFB7N8y
RfuE0n0k4Pwy7vce2/9zdTUun75FFeWH0aTJXUCdwaSQknjti0u7Xo82jE2zgSzklOB0J34rQLtB
RwPLNtaGBPXDvuqx0nu95uzRKBXsop+yE6d+lCyH7rd26ZMgWTPcHtv6J6ndKl7se7zBhC1oOAi4
9esuQ9U52rv7u3tPZSCTqfkKK1+AqqHEp8fqTONBpZVGYfGGmsha2mWzyjG8Qk/a1r2Z2SgDZ1+i
NOoYmJ1+6hLK7ARRdCLRcmZcoFwwbj1GUEu7AIwe/qryJvVuT0t8oG1eUOMthjILGsgpdM/gbggM
wq2Ci2PRNqxONmDjVbuPXBrNNsbH+tIYEbDF/IDVWAWFZPoOIOD6e9jcI2DZSINGleQHxGTGYlU3
0cG3j3swxACe3m+iOLR4oAF7brml/iW5yJCjNoHM9Y5DPDvICcNWgFZuXTQzo3x8qAcMAPlj7Nmd
bHez+VLC5qf1Dbro4DXu49/t0atf4Wp6a64tkerztJkM9kA4CGfPEyLxrL+LFKZ1D2vGgbFKL8h5
RHh/a2OFReVmrNoh29PF4Y2WYmZrbpjlsVvYKBhzeh3YRQ68pw8a02+0WlJeXvh59POKu7ZMwp7y
xfd6v4BJmey4KlV37BwXnB8Dw19mJz1k6bl6b5+bUX1AsQJQFzmVX/LrtPreKD0XcCCAy7w18lqn
/39ofyv4KTxgyEY5OPgzjn3IywPTAVEfXw2TAX96kzAwBieWvG7Uv34Df51aiGwoz0Nj0WLXl9MF
gMyIbEwgZPV7Yl1VrR1zbipVpUJZaUcHefw6vPh61A8YvGrmfR2LwLEvNb8WTTZMlreGF/VPt/aL
5RXiQQCSBgdhjmx4TsqWqQAjCexgBEGx9y/TSWd4ztWSgFsD7QKxEHQo5o6QuesNrgpufYo2Rdn0
7maLiLu5PoPNeKyVQf5Fg9kORKuwx41p+VqZA5fma2u0HZeCeawXfOQkKekdFMCnsR3227uTa3nG
S5QrTKSBWeZrBnDmvVvB9L9tiDkfCQ+veHyInuyzr/Blg3LvAwXQOknbRVmSocgeEbyKmdSmlnGu
rMZYm9BMKzBxrCKEgwN+qhu3flIxbjwLbzaHXxijCaM7ybsg/RynVdrUZIABZHh4YJWNk9MrCfMB
1toH8Dx7weS2yA6zRzGbYgawfnHmMLgbM3U9D6ig0Sceb1xflz0+BXZGUq8xm3/DHiwc9jI/Sctg
5gtYZk+ZiMaA7CtFL5jqaE6kT3FnhIcs9FN4Qy2SjJkxRYH2McX973RpWMjxeGBIT83co6etv4Qd
hF6wHffM0SevnE0MHG3IJyX9Zak1JCUjiLZr28voxrq6qD+Kg61rQBrzrXBPimsoiluaznV40kVM
yQYnSR1nUEQ92ld2XAQjSToglerdOsGghB+lrQaalRALQ9Tlqf2tsmBs03g1FdMGPeZmDQibmgtS
srwHqGFyUdgscd2MkKYedk+UU3MeoCf4Ty7WkdkoQBHvuw3ny+2TvB901dRnFB4GTRY+J5GqJM1n
u/dtfh+EsPlchYNg7UDONJQiJkqYgzWfSA/vq4xezT6sKov5KjwAB86t4fQAoy5scp3KPFIk3gAN
XdORpxSweT0FnN2o0OW9ZpHFoGtgZ8mALhAhay8hhex2Q/R2M0PZ+QNi7xNv6kh0dd4/oXMfA9Is
45zdFyfmIqJONj7MPmPMPgA9TBqy/0o/xxjNLa28czm829HMmROT0KsqUIR129Fb67kDbSturW35
hMhHfGThH7ui6fAmjh4QeJ2YcbSLIR7EX5NPzo3NoKJJyUvSo8uyg5uAf469yLqrR/4yf+AekODs
yulCSbnw4nSEG5NCXvNpsXQJ00hg9/lTOvVvorvawBYKl7nDSpSsBQsh+reLAE0Dk2YHMAIDOsQO
oAio1FDuKkf05dRiFXirvzQzhUToiXq4w67+/kqINtgCzjMYxI8UMILJOP/l9QWvsMKGnpkNiz3L
erT6gwddRM8EocnVDJSR5ngR/G+mkmeBSgS1vK8EL0A9XfhX3QjKJyOmh4LUBOYydHjsLKLZUxQ1
cIkTlOE5QbeXx/2ezCovDn31GE8W254ALWI39l5sIRgqAK+0BRLujZtmNT5QCuZ7GUFCNcG7XJJC
l+l/VIITBkBOyO/C0fQ4aU/K99xpXYvJU5wWHMVGYaQdPZWX3zvTTpqpmaZwRA+/oUEN+EdAAWQJ
RPDaE5+W06KKG7ETBIdvzvXFwIRPr6Oiofr3xGgDSBOcJT1Y7bpintJoY955Ejr6RpSb9nwyelMB
vf0a1KE9mKlwPmw3HtyYOrpRsUITNMmPISCFlBdjbx1y20DPFs6ut8BjkYAKNThtjUf+4bu1ojsV
D54iBdd4kE3V1IfRF0qcVrkQdC3JSLou7nx8JUC23hAhQxjXy9e7i2nUS4PDUE8Es4Ca2fAvzDGF
K3G+Gnac5vNz+PB+fxh91OmrL/k+RU0etgrHpyDxr1WHH1/xkh0JAH8LXaz+e6TDixBZn+QCShGp
Ghf2yIYnm68lDvqKvwEP8S5ZP9IcRL9VPXRTMHXmx7tvuFp712JbSXwUSxi9OKtZWm0L0Zr5Ccer
7Maqq1kGaVdX4bILvn2BZPVZUoEs/db36W/jL0NEr+dVZ2WkZLXi4v+jGaZuqy32hFaW5nN9Wm3W
i2WSx+jEc7CFaRZZobImz04o8Koj/81xuZ8ej/hbg2KkIyHYCJgAL5Cprdd9ytT+7QsMLM8V+6jV
Pzro0ppUevPzpYG1/VrFqPMhWGAtKNJMTMVNrCLCHPaKAsfoNVjeqoqE7fPFGqfB3HTndbuboC73
uyvu/77d5AeMPWBuAxCpVCCiD4hntLO8DNGR8qHGxxqfHgyuS7/tpLKlU3XAUM/nQWQEwBozoPEJ
AUbPKeB6Wj8iDGVZ3awAu10dv03psiQ1voX2DHHSHu9uUw+A4TriIQUuepJPvInaXomh3/ya+v3u
YyZSCN2GlNk3ZxDPUOSNSwIMu4yzXcqYGhV10TeT+NFrPP6+z36qa1I3U1Lk1RegyPprEom/wwFo
SsgbEr8erOePjw8hd5mh286LFKUY+D/M8+IKu2clagFq63FZ+mnhP8KFua1BYRV9N6Zj0Fbynd2S
kHY+Nt7/TdggBP5C/ara5p03WUNic6/WESFwD0SNJ81IJHgJmtsOYuTs6XczyZ+ftNn6KSlm/0Fb
9XpDrhn7k8W9+v4iDmN//H5ze+tw8TOmZ4zQ7A9obl+6vswpU91f86b4vpemUE13aoeDhfVmIREF
sP7lqxvkymIUBT3NBjJJYOM7Hs3w4RMOb2+P7E2sJn+INXGhqWxD2i5QydgNooH7c7irShHuBeTR
VRmIr5/37JvA9BZCeGJS2B5spybMReRczvYe0UW8UCbPs60TU86LbMCOMjHR+kTWSQCNpu1GWz93
4R0W8QvSNyzTBIPAmLFd+gSRXH9PP1j6FhvKj9vY8Ls6Zbwh/dFHYnk+RzriuCARTqdMs5kpWxf7
NlAXT2HgoHP6/Q7cxtkkiCxH0m6gkk3wnSG3WZZ0Xh0Rf6yYGVGNGrn82jc9lo/4RlnpjTXCawDy
OoI/uSW5bbLF2pz+rghIWQP+qfbExZE4Ffm7P4WyOEvBkGqnDoKDkjSSXISJ8AuoT/p8WDVbuqVX
CvQ5TlOjaiK4U/iAyfAgj5evrrxvXRLzkoFegTTN+kmrYIHPETWSTut2PJ6i5ifGSOOikccgw0UE
mk5SbGIEJ0D4V4N1akPNJpqGGADkt4d16sD+nuujSzmN/8DrWMk1SZZXh6+/spUyst8fz6yKKfxd
ABIKFBOw5fI+WuSYP+bqppgVUITdd4cQMV5jFQFP2P70qGehcyWs+MsZC9RXUysupqAXwFn0digK
xAOQWrJO1RVU/OGvoib52Svd+QJtDiw890GCOqC52u59u9Qpo3iJsh7AGG4W2DhUrl46rWHivY0K
xP3RFFuszvfdipBCYje3OpLDdks2h/FMB4IgRAuVVmo47LkhGT2NdlJ1BUaXQYnFdZH/XSyqBseV
TBFaPNTFCpQia6eqvT5omZAl0B0ubFfkNGRDtoJMw0vooIlPssaQi+Pq6YHjLo2fmsgKRZrFMdU3
5IoIQnDEAJQcjkN7wXnZ9Ghs5Wf0/oyFdcgwwIlHE2GuOPCo9uef1Q81L1f8kn56kcjYXNx+jQ2e
MlqpTnmt9utw8Q/1ftC/JwIU9E4ZhGNoR13ZS55Ddw4/HGsfD1ZSsczzUjKZhXuAG+DMVFyPe4nT
Or3hVb7BCZLE07IBw5NosBqyoEsHVO50tJEhWU4IECk2P6lOoIoq8TIzSTlKoBh0MwrVPmzwCaUS
5+n6dhGYP4e94tpWlJ+0ZHjV321SficP2Wwcg2fI+gScosHOeXjSEGO2HZKMk1bREFJP3Unwaol0
CvYQiwRK8m1xuL/hOQ4SYRgP0rbZxZY8zWCQ56/y9iguZ05o7PB+qVR8/TY4TeSvuaFxJqNLAMGx
7d5ZJi1rn6lITvPJHX/6X+KjQgE6anYNX9OMogui6MQzqCiXgQjCY/ghJ+he+LbO5RKW6e3TQgIN
dv52pEGv0UNIsTuX72RfnBIQrHO0gkwClNTOAC2Do/Z4IqTtBqcL9gPlId2/UUkpOQC8Xos+B+D4
ZcKIYSkzAzcIKEbwBIuO2d9KuNNTh+xtEiIqe6IKcIfGQNiebOnANenbT338bUpjYd25gAaztRuR
7lIJOW+vyQgSocxmzOdC7ILWR6ajUejOeR3p3Xpk1L559UYUwx7e4bA60IBdwpIyJ5l4jECLkNJe
TpKViff+3QWYRA1x7Xf9dyYyus56kgKkRzfofbqwdQhuAfvkJmvzt8LiHsekEzFyKJZFWTSeSgRh
Ts/v4nm5I6/w4L9UR12qTL5qoYFyvZ7YIJf3f2xOJ5rueCt8HiMytkTdoEXVPbiu0cFzeEw0ITcz
72esUGX26HOkWh9bxGRETEpXIZoFZDv8Mb9nJm15LiJ079HbjmDJW0o/U8CMefZU1Xu/+mSECL4v
PoqwNa+wTiHyVq22FUTnb6ETH8gyguQv8gSbYVdlm4NcT6Upb5qRsfiul7w4qSlPwuRr1vByQsr4
5MdPVYpejJj6xOKyEZS23J4AHN3LwvkBGWYsihNUEJyu71+4yzmWVZMWxjmNKBm1aNbKuAnxQ9ja
MN/k1vYlztX/iRrxtCpbxU9dYSND4mEzbFBR0R1Tv15SP96Jpq+A2xxjfnrABy827/5tht9I+GAd
wZp2+aJ3JoynXmtVFK31PsVYHuVh0h/r08KXZAEhgNKNa5z6d60E7O8mnU2O9JTumuRD72Zuel9Q
+tmPV4iw3LgxssCPuk02UQ2c/PPgXwFjUFtHfEJxQbWdhOT6ppk0ZtLxpKd5391LBGpal8mIuE8S
SOICC6R7971u2I241T0WO4MmFWU/o45IoErjEBGV0wupkbi+iKUHcJLHT0wni+6pqw7cutm1LhPI
k0S5wk9Wr/A4rLWCo2Pn7M7DQ0hO3sh9gi94e1Dbnzz8iRYgIRajtze73T80xIGZSMl5VfxYrL9r
89X0b5Gmusdv+mlZ9PO3BYPOA7Tm0oYrms+3jhKkVn3nFUrn9fxk1FU8zl+ArVrNJy8hVRqSeNmf
tI8Mp8UPciVhKxPtJY5oHdilTiI++xa51eV4fk5PiB9+ZtJd+N+F2QIMEFT00qP3XUCHej4eQcax
yQMYkDjMPYHYr9y/UGGH5Tt+q+sOl8mP5ZX5usHysNMbNdxOcsqcdVZ6dj+465TCDnHtU3TG22Qk
SVKnXmS/lLgh0HgLjdknsdSOk/at65vc1ddbvhHeH4bhWaPrWDunCZopVgzGI9u8BFeZJ4MTPmPe
WinwaM8cUaSDZ8RRz3cygGxHg+KnVsITnI56msa3y/ooiYgHKJuFAxP421a244pk2HO2yZ5GeU54
RYeR7EgVR5Rgi2Ke1li78kTdGeet3CImd8XRNjfli1/hc6bEOfVy4qvHrxenAaWgwCvplrWgkCX8
uDlxJqjuVNMiy29XOmveQoEtxDDTEKHbC5xe8UHwY5zzm3AE8CTS8C8jUCtULP/7Z0DMRV6VQCii
aUsNh5cpa0amd+W5FCmhGDeB+imsCuTVh+PRHv3ng2gtx/cFVV1FaA04Vp6iBSAk+29gyrDrIbOx
j0Y25/7o4T7ULYuh/9QPWawFCbhMvfLFP7gCBUtNpY8GS2lh9iCcnpbV4Np5wRsJx33g65pJCe2k
4aTIKtzou4zsaiBShB+Bnkz6CqFgwEUcqPZO/+W8D7cj2HjtpqAci2fl/qXDpWUetayxykRtbKfc
7XjXWiWnAGXl1/P/LRx4TOgyJeZ8jZHirV+HryftgE30IRE9fiyj+0vETVL4+b9vCnUQ/tkDAGN+
cfM4ZfC7Hfi3vUcxkR0eBu0ACv+KK5ktV6vs3mmh997RXs841O9rBnHL3b456354Cc2S0dd3rUOv
No4VEGiqXCa9sFlObHOgVIQ0LF98KG8JPaOggnYdUJrYVSphqC4h4QvhH9XbmXfU1f0/NPyGA/dj
5KEH59wBl5n1YQ2L7IfugarjIQemOlEbf+XdZoW7VsP7wXXr/knGTvurK+jFks5V/HK/l6jiIEIw
CqybQy7qlGqYXAQDZ4OkAhNnlGzn/pkccGWcdFSGPk+mGZhfYq5acQQH/2+ipcV69TzkJ8lHK37q
aJVkPdDRK5EW8pYlFOUB0/qn8EBUI6owkd29Qy6rbszaqYwQ6K4PDFtWeH6F/f54tW9TypmB36pQ
X+3ntt8coNPHHM3j7+O1O8Pns9PZn86VZLYqpWkUlH0WcnqA9vwmNm3UPjlgzzd691FWEk402E3F
ULkP8UnKKpf36mgfw/u6LU/RrbNUSK2Vxjzcjk2BhfpmOzdjzlV4oDbo7CA7Jd6hfBwMSZLeQQO1
tPDqPCn0j9Wq3q67WN8FkmeGLcai216mTibhnPqM6vrO1ZGDlvMTPx8i/LnPHYRCrjh0MVRP74Td
76CU588KXzz8OlRED31+LH+Z6ew34RSWTuXGuFJaFJdPe2M6NvjqfLq7zPp7ShjPzU0P3NhBC0oJ
Rk3tervEMAQIeQkyKkDeWSEgR1sDmiWhIoXdskdM5/sHSJ1ip7M4bXWcXBLljNySCdyxcw09iIYI
vSs6qGrONJheuSKDXPfW6vLjHDhmf6kDeuoP0gspJlJpN5NQIdW4YDYxdddcVbV0hRL4sbAGFr8g
kPo0mAJI5FUeZgEau8utSjTrewUSxIOHttpAuNPtsxHxNYIsH9UgZeTmsepoaGQKCUTDi6voG0rE
LwJGc7sC/HObaATpaYsxlKQMrWLXjBVsx2+QyrKzlFtAzJCC33+4EwiIU1HdfuA3BmLTsFFa0CGW
VoJRVoS4Gsum56IwA4fzCLaB//QTwfSw5jgvKxDZ2BQ5+yqXcAkjNNoAqvCv8KUby9RjsMRSEaB7
D50ijgoEPTwpSPbU6O+GoYUd4OyxnJ05TNHdaUBjl07L3XkiXFx9xvR80J9p272iODQpAY7miUtf
fTUQWOb1GfUeTyzLoOUBwWh41IFSlyXaMSdvAl/W0enIEZUP9f+Rr1qlQoodtgnsMYVAp7rAnB0g
X2+cK2Ky2IVKIJ+nByShfntQeWzvE6Y04CjqEwjLFm4YlDSUp5ynmj1spu1VpMUmx1mEv01xOZI2
lfMTSofFHPsBS7Yj0CQ3GpQ9PLFXeiM472UwW4D1h3SNPdQYzDUGNqdR0h3wb9yJVVABXN7gawKf
tU0pSHbYwajw5Wn8zBPS6GsmDagns+eDEuIhGtTi2kCn6J+s7W3SC7WA9xLZiipUy+2buqE8KUjc
wIQEs0grJQ3IC8sRZtlNS8J5p4eS3RI+C48Phn0nA6KP2zN05FsX/Y6sihrmqpb8HzyoGAh/tQmt
uNaApME1hLq8cxVXIcKkLFGJdRmdGeuc5mjx+XU3zyLa5hwGIe0QyI8bjoBe2lwrCChEuDR3Kg08
wdi6+JGp1dMtCGv4I4aFBj74QI+wNwoaat90+xyK6Rj4p1AO9Dd7eDhtEil6217v4RGdDJuSPxiH
wd2Q6Yw9+moE14f9Acd1BrctjTO3Vjs68Hlg6+j6JpjFPrcWb4ziNRQlCun2To8ysQ03/PNfjVsQ
ySCAJD9Xots1LBB8D6ludEcPFRlkER36Da6OtN5kH9gsrVgWuJ/cKN24eLvSA/ssiqOlAcvIy/Em
QhggKLzV5VweW2UJ5hbNmaT54r5R2yq7gHUq7bmo8NF50FWfDm/3CURRty4crPv6X9OtCs1YA3xn
O7MHcev4zj4r/IjHEkMIMpBTunvdZkLz4M363BNJx6UYQ3kSeFkryY3YYzeS0crK+7cbaSgO5CpB
G/FNizGZ9/YJRaeRn6Thkg+3UhTrqRYvlMmEsQZHculSP3u29uZjAx7ekOkgiVwH7wP0FPYqOYXk
KKva7tdQ0EWDxYJmytFV8CRsRwKPNfusslXddpnYIfSe3wTLRTNPvtVrraa6cUVa5f6F8qEW2fbZ
fsqe7HnaC+cjhf11FeaQQk6phCmisynpxXSmhOr4n3efyGn3lGQBL61I6hp0jP5lxkw2NKfVtBTU
33bgHEv0X/6PcUWk1+XUxIe4067uCDAqbRWpWp+WuGVXa13hdu/H+JRSUe5LK9tbKKBwA88js5qN
/qRkWg9sNLa3muguTGa2QRfd+J0VAcTK1AWlTXSYglGO+RXEdFEC3gpx3oiGNfSxw7sIba5QSogI
3XkmpIcMJnQMN7Ia54I3fa5/28SBk++rpHPebQ7OtwiuVC69tc06qeoAipWzReGIwNwAGf7c8K48
KrWAK6bEC2eGa7EZ1xatBnxO4CmjJW600Unk2a2xEZnVcEVzy1xRJJalM9Dk2zy+GyXPcLvsm8rs
PTtT4IPq0UaWlpHDQki+2LUceO/Qjfsnc047Nk77Vb1GsiwjbkR7uFgBUynZpizlRNdN0MuugG62
4Opwii0Et0Xuq6iizX/bmCjw+prdIgY3k33fpRExE4IIBi1IxOpB2gJsqSjtJDjxnjo3rnrY3qqI
tHuagRHB738i9ilibaXqBFLT/QlHiVUpsacGalzM54RtFuV9QCxZv3extFAdBDJfWxMzxrxSwbG2
KNa6S37WgcmgweNHU6vfkEIaTQPzGYGfu7ffCkgH/j56F9H+7oaPYhsMG0mDzzJEcaX7LIJYNFje
DLwfWjR9QKHRqO5EyO9HcoucVD/24VRUL4JE0QxIgO6iGe6MAsA3TrxykWvJ76vK4ytAkIOhfbp+
G64Of6fwdFyrIytQRlWty5q7uY26sysnPyrv1kWGXiq56+KkDwF+JWxnmjmBo9YebN6MqlqqRrSr
350vkdWfwuSCxGm9M3JWMHkAT+JJi79s2R+wVd0Qny+h6Igo/rJfojWy0pFFAsEDDNqEL8tij5fZ
GjYAnV2gTB9FFLBoAgK427gLWSCqovWgQloAbG4G8Oat9UqOshyBNfaqvzV4Rb1peswUfxNYxiJ0
gR8Lou3iXE7ZeUrQZU+cbYtFUg9TlNOY0uPHbEVn23voWQAXK/Gpjt2pz7iKg1OcJh6g5GHP0OXq
cjRc0AlPV8xS/hrNn8HiEhcwvgCzlTzzEE6tx5P1BqCapAtT2uht0UFgc2ls9wQAL1JmMWEAc3a0
70Ls5OJcmeYRScLRNnOeUg3gdXl033XI0tHZVqOl9kbAwWZ/ggzc3EASRcJMD+PEojfg4RZx8COr
4JMpCDFwbro93UkKZVUQ8GyTxcGN2Lle5Tk//rkqBslrPVxNAY8KJ1meTBh67/6Ixu+Xeqsp5C9s
eUMnxyXu2RcRFfS924kOPJvWPpRhVEnT/A5guO4o7ruslQbz59SJ4mBhOF2t6zHi1jtQjoXimwqr
EU1xOSjSYJuPnbfllucqN03+8QeCVLjE+FBvw6FURQqGHfOli4FArv2n38zwVvVA2BeXYYA3+CyW
ZMVUuFkndAYPz6KjU1JoBjOHzrtPq/tQ9o0eMmHrdUi/gds1CWxLdqLpUvZ/teRdBqXh8Y9ZTZSw
0YBwos4cF8l1wc/HG/fuLFg0v4ZX9RssGoYdi5EmTDDsp/GGw+U7zV/7hy/t8S81IAgc5+XJwg4b
Qk/Dq70UYBROilWV1aFCtOF/rB2X3vviK9GCDXyo396ulXr6EiWsl4xG41AqYHoOWfTbuczMP5ml
+xPUjsbRg7dog43KP5mZLHAWZ1vxBa6ygck3oStMw8+V3iZ16l+LYDuvlJ0hRGvrmV3v0nJ9wHLG
0gH5FY1ADM8M68+cCtxb3pWkhA3UzKpHGp7ERqVATsUQtSEd5EJ5Q4vBlfYxtt/xGyVIAoA4KROC
e6sXe4nMaOorM3HlnQykxgqEkBIe4pRc7uhvt0b+K1E4ZUWCNZiWexFQMy0BZl9F3KkrsqYJWV6j
CfYMoQ14dgU2vV3JxqxvKWy6X+KwOwE/anc2DVz9hD+jM0AiN6mYY7gs4LnHiAUUtnRZH+HwieB5
75N3AL3A7rVknSutM4SSUIZw+lOYhSXpcnITxBucmhbB+fBXjbJ/rIccmTw6qBzNV9Oj4m9nsk15
AdVKS/0fZszPqCaI+BfDfKqAVibd6szf7V4yfZW3iV4ztkTqOse9FlY9BFzP4xqyZLvF9Wm/oYtD
Cc1BfcUpZz1wvuXu65jBC24AEa0DevTbE0OQ9HED6ZzWfsdkDyNZpfbxXR1ndbL1ZIKCuXKRLKMO
2LStyOMDCPoX6RjVrN2bkspl2JNeOrKqfltOCohlgKPM7fJtA7/wblyU2rcWEV1AGKOvsqfPU6a+
oX8iEN0olDtbq0TcuGnyYYJKitXB7S9oLo8fu3e7S4LRiFsdDEoz8VLitTQ/sSM+lev0TP0EJenK
u2/3kLktdaxh1zA6NpiLiKty8kaj/rTyd796R6FKZMj8AvyUWrwqGH3HIXrh+m82yvSodJd88KtP
7KPOjzyvuewIxxlud8+Ck4xajzphD8QRozI80NSBkwHy6ctMaldWJy7xEkANV5umR2GqiDcNz6s1
qBF1xFy6nYXwK9/LoE3m12IAHMU7G/A2qjcxxLmjULkdOvqXINhkDyLjV6mc4xgLtqrznh1xMH74
GQw3cJ1A1Oef2QG4aIZX8XKn66YwQcDq11/YL6AikQtxdjEfip302VzXCyqXketAyVolxeq52hD3
ng8XrUhY0Z0lso8YJDolr1QArelFjPPsPinkCjejY93JLEvXAsI+A1wZZnBZx7PDbh8si8H1RQOf
tn3G4KoyKxmKTN5XYfLSqZfCgzVKju8dJnYG4JrGTRwp6TwD9u5CCFJw8yKn3NisrSj5tiZEpDQw
MWd7ienu2jc/4fgqZiiuolUDCx6a409GE42xSttf2U2TAmFyDUKU8IqE6KofSsrRA/q79x9fJ8gS
iHu4uuj3K+txmAUxlhfZMqWQbk/TMzkw7ZjXik2kDk8Hi175QaWCmvWsY+z5eL6k/NDiiXKhNbEv
bVAmbEAZ4lP+2ttTMG4qcypjNAuD9Puh80QX2kkYrh3De9ebOMHaWGIKWIuPVw0Y1lFn7minheda
J7leDzLjpJ0ugAB6ptc0tpB6sKWpUAedL6UgQz+K12aS08/Y5LizpYYDSzxoZccXTgv3+C84DDgF
+rf4bXkhzbGe3XKzxlXAJIMIUcPfs2NhdGI4PZ85tDJI9nbLUUVUrnBbfygyZcDqLLBBjpnRFVw8
1bOp0BaAYANG8eXGRZTXgSS4C1pCp54pTCrdRWiyzVWp+sLjvwh9INCpq6QeT2aqzErQkfWMditm
y3OrknhiiLHS8LZol59IhwRrDXifVTHfwOPipK2Q26xhHqNoQplyUfOfXU44bOtm1eQ8FjdT1GOK
j6E2Vp5BDUAiyFW1QH6vxQ8TpoKHF41CZY9F5Qh2Uv0qOVMsfbvo7aaunWOCy/dtseAGUHCXBpFk
89WmuWizVwnBdpeAuYA46unEKr8UgGw4RzuaRt1pE0iQafqD97Xwv6Ja2+p2Z5l7iOkQHfORU/xG
WXHRbRVUGhNbKZbyuqzjL4yOLxoAxQHXR47wAEjqosMa57m6gsWnOl94oKHUepOtYaZRCibH3T/w
BNbFSVzp7IjdlvTwRBWt1LzAobdnIDXX4WqNUuY9q6R+uV+9IiktaP0QXoq9QSzCxziv1Tz6AtKl
PtHSsQUBCNlOSw/2DVPv0pH75hOSCPYvX8HWcftMOt4PfasdHeORFRZq6x9GmI/eJMW5NA3vcroK
nEF4tx8eAoAjcEK/QlD9COaUetOwHL9kknUYIEQOZ6hKLlAaxvl2MnUPEGE0ivR6t+P0COyKnwqz
5Bix4hglNp5dq3tuMRKKYmn9FNfT6PW7Jc9fkfz5iZHWaJC6Y4vvGT8Qv6gaV++jRR8qh77H1K92
/lsuZk3kNimkl7S+TnqD4JrURaTPFo4OoTfcD0X4IReeVpkGMGWVcmONy6aamK/u1MWfDhsL+cpD
KcCjaJiU0up4k6D75HFRJy7WDqWlK0a61Ct1ZT/MdL2oGZookeDfBuwoeiLX6XDGe0KAAVbAuHUZ
GNXUF0VEgWEybw4iaMvAWqHkzo/zwPnF5oey5fjBqZzNYJgnnNoT7n4/edkYwRtjrlgDz70B/c5v
5zbSG4NrnL3ftr+SSs1nkOFiXQHPt1B/Wn+HXeVPKdg5UN/HwOQGkH90V9Ay4ONHulOqZG5o3o3s
M/zOB3k0J43U8P6w1vgklP5FvVYNbseEkruT3Dl+AoiAeES9+eB3IEbkslLXkNpb6r1XdlpJcAWt
PCV8RMJMzFjMHby2b9LuJgNZBXmzr54ZnStbX1G5KTezFTKHo4yUvjAoUBlPqZyXYOjGaVi8ygCt
CO9hBKJwki6snJZ1HpxP+91Q6I4R5PzGPYJGyHXsLxsLN/0Lpb44SaSABDhCYrtbbcyx9OROh1mz
eh41EX51aMEKZxdDJ1/l5ZxixR8KP0iUDRhOZBDgyiFBidNyf+vzCow7IGkMu4ei2cKr0x36zWDD
JjosBJRf7hj6d4OIOHwFIZVpE6F5VhIJNUa0zfwuPeAaLpBhUlEbuyhYRLabRsE/XWGRkIAnzymr
AKdmvV61k5lOs+CC8PlPA6EL/NoIBx0UIIzdDPukK1iNOJTCNAfHTT0qfvqGn5g3TV6UIsr34FJ4
TFuFE4f1poSS7fCcC9R5GecdGFPHSB05b5hzoHmjSxXB0X/JjS/d6XMEgrdB5GgZzHr5JVsTDX0/
ufDwra+uSSXVesNeyxrXAwe2j3P5aS39cHnImlYJf4r25+IavxhkvhfbjpGxaDqmKwzKz4n4ELeM
YJJzyCndBd+mdYzf3n9iSzhwVsTqpvPaztRPhOO0oKG4Unrh4AVhpVFBAMNJIvUBnZ2g0+35AhP4
idBJKsNVqjio+XClI+UvaJgiWCFm9X8VRZ/6HjtGuyenxd7RD0B1v4NyjxueL1r74ZG7UG/qCfgq
mF2F2QDjasFEtt5aQstAjw3QRpHp9apukUHR1cWHoypYVwT3IJ7NcCpmwIMAMvOGYpz0hXL7elWd
wYncIAzDAmmVPDK39UKm+hEfsHUALZArfCLoxZRBXTCcj4iiwq2mHezC6nCkU9GX3MlpQp+9McEz
l3P3GWFRTZSca9kTqExwOF8Ja9Ct27V5VE3YwdpEzTnX67d04shRtWJJdr38fRCve2reqDgXvsLB
a1qrYKrUTYF6jFhYOSrRopdlP3PorADpHmC43RY4CquHARADbZvaRK33l2gASRrIW4I/q7GAbCQB
8OjkOSbdwy52sL5f4hPK0WWYo2GaS46ta0ATSo//FbA5St4QzDUA9WNHN5ikiuQ1r5dffhE4bdXu
R8t0O2yWk2rG2F/Fw61tZs4a+mYBqDL/8dPV66isNtxFWUM839mq02gCkFpoYGUSWKKDiQZALxvb
faXn0kH1iOSysbCWdY7GN9SmG4pDWWLmxMm4h66gftb5vW9Z3UBbrpMYE6ffX7oapqbGHxwJh7RO
TLVO2pkEkLu21j83fphk0hDjhKwY9wnNkicfJBCH+L7/OTdlSsyo/9mpoXzxHxtM0OOO5jJ3C1lZ
VNIpDnbtpnovrlJgGJNsN0P/V3hA14vTFynw4RwnQm2hxVe7AL5Fxf6W27r+zGodAnfua3xffAN3
gKpXMr4m8ZDTQkHetAKjqTQONrl8CV+o43vul49+8dt2kOy8ebb7zp8F0WLxZ/yXFFz8BujtK4Dg
im3ZLPWXwRLV2Myew87VNYL5CHvsYEj/MqrQ9K1MGULBZO4mLeIdbTOX9fiVaoKQ9yMnW2W43G7L
ieoMiGk8r8fvuCy96JJNyzXKpTwr2jj3TIPAibFYx6DQkhLktLJ4/cpFbmLxzj4KI67eqAaQbqtl
fKZ0rxGoTqVYKG3TAzbKRRfwTywbx/ZmPO9Fo0+Mnhtr1BaQej3a83uejtp+P90BnQkzYz5jzrLg
QnIX9FkALE3Gq13CNnmIgka81sgEWpXn/2/vEaZ74Gwq6jUcvwcbmdoz3NNmqgWiRtEsyfYr8GtC
4PeqHbj3Rn5U2RbLhC9jemv0acjIyjq350wKKb9F6BM5vQXytz6xr651h2zpF/3hk1oLuAtWlCaX
e/pADGwBXIk0bIXFqwG99WhqtVpRKGkEBhJ+oWU06r9YjNX+9sVOdXVUdEwAK0fgDddnlJu/NVGG
kc9XRT9VrWeYTt3rU6ofqZLlrzsOXdgN43JYvTtp7xGsVKakxG65t6iXFyRLLMq37aiN9IyowcTb
tN4roqKxM8vkVxBHlCkR7sD1wlIQ0sIAYoqSAuT3p1Hj+b5/X+i93ya/sb9Xkj3RYVB4lS3JAsnK
rsEUjUykJ7Dksjo0GQi6tMszRfnQ0WHPyroJNVCR6AfUnrZ7wIIU5svXLKBInlkJisdT9JaimwK9
6SMz0jt9IQAnVjH0aS/qH8LajGu8U1PH1Y61vpiB1qrswQsn5WzbSpdkuQah5jpYHvbCvB/Ya3U7
sRDYWflcwZhRT1Pg0H5CQzyrqelAa6pOk9vPiX+eJgo0YGiJERfFoyBt6WGWDT9ZmNym3tVdCk+D
cafYrlFA19DKFP9zuEp1fZP19DDAkBv49LUIJ//WVSl2nZTy7QIolX3bFsiJo70lyBtCVJMUc01k
99lkx/+lpJWc9T3wAs7ixfs7i8oJ278Q9dgPacDC16HQe4mtd1rK9dKPxutjLqNfV18ePONVlFqx
ZXrSNw+R8ktJKSVu/u5kz3Mx9dUoXHa1NNO40sCFnDviQq9JmVCD9PGBfGwc3EyK9MQFJdR+CdvU
LUsxsv5MVN+XFFbmyv3c8mts3umCRjOBt9GytabgSRswzuQYTQuQgzPkx6UnaCv+G15iXpKGEDuc
a2LmuNlPJKXA3U0CpF38EFrY+7Xe1Asx26+333eVhHwPktji+yJGcL/kugB0qdHjSeXeo7qVWqIw
Rxmj68lvrtZEi1BbCahDSYU56IhJ1wkf3oxYaXkxj3K0sfc/tzabi14OdwDQzbkPedqTmtfaVDIh
ozrzcOpwCpLNufQY9HQAo8Soh5gPDRvZXrAowB+SXPjcd94uGxsZAvdI6fC3OOnUtwxde/p0he+U
nYzeRkpqNQZGsFu4v0k7fnZnqDzZb1RkL6jpzBGIfhz2K7dj0hzB1yfntFl7DcmjBwsc61JFIhuF
gtq1D3DLsV7OnXUIw5a9NHk18FPlbR0vGnLNQG11layZy4v7jnxgluFmf8E/LmppgGhm7Rx/KMWY
7QLrxip25Zy5TZfSIzP5g9mfxCEbfe3fjsUS0FTpAEpdeom/7Yw0RJ++HOrKEZtWPShXiSsHtr9G
zgZ8RDiR6RlSe4UdboSx4NSJSGVFRZRc0AmH0SHkI+O+UC7SD2YhPmHHZpaWQaEwCyRKk0Dr0p5T
OttuYFNA+iMG7OAI2KUOrrLQpzWoA6Y2qtBjNjMBwnho+q8zmfgvP3jIgRaPuB0gee6RK/Sgqx/O
heRczb4thQqafgO5Nx4amkoYI+gV2k/5ctTZL6rve4awm3BJg+lTumr9gbUy6yHfnecgankrn727
Raq3IKsueWP1bac20opLehlD3GasgrFXyLfdaGxynh9APcynwARObQdNgI60UwHvMdw/makuvyo4
8bxyu+c7EKvU1jWKU9Kyyl43jQNCkVeLwayHr/QCF0F1qJuya90xbeSY+6b8/RFrauszL6SKo3ld
s4hmjPU+5yzmbN7gYzTlNOBqmjoyuoRyD2wvwSqHPLJh7EPgNFrxWj6EUWns45pBizDgnxEmJy+M
Y4Gc3UR2JRVmS29qpqTsLoCY2nzSFun8cC52eebAY/myd4J/Jk3xFo7sAei/4vIs9syusz0nhoE3
ZiSr8x912TrKihT1N9/2FywWcsqZfkWdLOv4kEDmZMwyfFZofgz2GC3K4vc/j0zBLDT2eTTsUcC2
Sqi85mUUoxW0oDBUBZzAEz+cH727gUKLoOA51D6IPMhKUCLxo5GxhdHqPbcyo8vKoI31M1KXKctU
M/+FTu8tlEWTi1QFjsPlD9gVpDO4UWlqg8ssXcKhWfJJreYEi/9h6j9ewbOCdRQ6pz0YvHJQVTA4
iPeeWRYcQ7vCrAA18fGF6LLNGIgltWM8P+IZpeCSwA2co+/Qm0SY2xev5Wk93NwHq7k1XV7kkn/z
+3M/3kglKTcoo1thQvLcDMsvnB8rI0VVBJv93hevpobhLvETsXv1C8diJvRShilgS2ossgdp4PO0
SKoyMI7WBpB7VYzCxnV39Uq8Tjs4pMg/4cLg4SHDW/93XiVH6i9KySDQxq+6G0gr4i7sOt9CoUyP
rkPcvXVE4pz9J+yM4QFjP2Rht0parPVdg1PNvevqOu6+TRqbpIW67TYUb6WbPP90iel+KmwbwWqd
vj5Op35IzMaU8IST/RDDxLoquitjKHHfIBqLbZzCi8DffQ9yKJ7ab4TONTe50DK7wPwuogPFyyZ9
PQh0f9Pe94JPX/fpzW/dSTfjp2tcxsVrIwmOWeedvnKQqBjjIEBIXLnptm6jVGKdhYE4JnHBJa++
m5QpjzftWbBhriio/lWsf4AbrO1CrpJqztY3v2CyNLcuk8zDFJXBb5bXed28IGGE/ZnRtr5VJOvT
LmT6f6zUzw+b+NT7lFYj6e7zGYaOpfpNFvG50mHOJNAPrr30GQz9U7sQzE+43X5V+bpbYOmBAzsT
qkS5PSzHlpZrW4ESw2NK4cIkZktO67DyNiMfa5HObCZmrJP+8991RWtWvgE2I59O7HMF15E90vQE
d9Ng8kvhHYukjSLDN2aEBvVuUmDmLnI6vd5CDZ8z7qFsehmND+SjHzvKEJtqvFONDUgq71UC+lgn
q63v8/lxfdUkQZ5aR6beLGMbWsHf9Rx02agYvOQs78I7KLKAyq7p8LodJotylfIGfEkgRpN9oZhv
BBWf/6QFJtqdKb8TcAT1LpWWVJD5DyDtqD5ryaqLhKnQIn9v5PG2RYwSAnCx3IQp3vLBxqsTv4jR
nrnFXq/VPSBMNqWxvRM2QB709sXDQ1bpN8heOPz9Oio1nlFn8H1/fNFMfPsW0Hk9XDN8Yc6Pr/7j
GtTErIr9oMJB4orhps3uo/Gk1W6TD2geYY+xr8Ow89Y5PI7UAClmIiSHOt5A72po3484H2sIEd9X
D+qm+8gvh7Rh8NoAarZzs9iT9os0Gek3Y2womOZFg+5kr+E7nFhkaQaQnxQbp+vhWifBJ8zLidds
hSJ+Ck+ZuOAuagyW29Hhu8HVTYgGwBONK7Tao+RPvmxaORVrHxuvjlDRrZMQWkOxEPtp9M+x6sXR
oBwJERIZPuRpZka6VPppYBsxOa7IeUcs5S0iVtWDkyejkX7D/kPmP2lB8eCI9UyONOE/xcY2M2es
BLj9JUPQa/jlD5w3I6U4LJHIYDqtrax8XFF9BzemsrAN6cWsZujjcdiciVavjAyhvif01N0vHzdX
xD3ZNMRinEeXSE9PAycBbty7ERf+bDMrMw0EAo3mw0SApkGHcQEy+bKP54Z14c9vCd6vXk47AHXD
NPauqTvQTcxv1T64X2IzecRgZZTpQuYi4gYL/kpLnuOPSRHurhdHd9yX6DzR3U0THI0xO1yHUYra
mlqO6uubRuPZczKTyEzEzSdb/f783ONFzCmZp6pYqBWznQjRcq8GRzEBvq5hjqHnrcLyyBIQltLK
di2RpHNWTWNFsieo3xTe2Lhh6YvC+k/TUGpVftD8D5X249oZkgC4q3F7c+zQf03oc3eVrK+UQNvq
0R/hcz1Pcg/SJxC+GjGM85WiRMNf3IyXYP5OS3a+SWAKmZSR++nuybAvQRSAQGJddkAD84fhhocj
rcgNxiK33sqAOMFCNc6UqKn3QI49MCsB9IB/zPtQJwaUYJ9KR3PxxnzEbEudIxSzSF6El0RcsEPA
6Z7WCwenWc2bLixVmgGvedtA2AdAQvYqQp4iVPjqzrpWmJPd6xy521sVT9BStQopElMUpLyO85UM
qT+AM4zo3Lnu+buD9OH6x7LpH4ZBvdRH4iEU1ECBENZlmfw0ZJ8eac90MWVUwvgh+fLPPIbndUjM
+peRptioLHn2awxjeGdL5AMdGc4xBcucDXVvZVJJslZWz0AqQWPIObXxeFH0NGLdRk64RIxeZKDM
rYBHyFPKd0pyM7xdPoXgPjtSDcz5J8yUPGJcuIDb3wCJvZ46TkcXnvfMhe4BAv9Eg8tYHWp5jXhQ
cTLiWUjTlqBwSRLdVQVojMqvQDD3si2Y951KHk0FC4O+0R2/qbBQ//V0d3n0r2H+RYMqaAvQb8CP
NX6ElYzxDtpYIalHQqwkFGCwFbBmulrF0APYmBm1T6uvDUsksLtND7OAfskvAhrKcLdsPtCXnE4W
VE1GQ2vRknv4sXWYeqhVYv7QEoeXMzozY+f0fsO06+JkeqWRfMcOOMngMl5CHEUsM2taDKQBdbHg
YqySQoZIOtLvSXKP0/VPf5EkJVtoSfzEOUHqZPHPWP8rHLIGqjpkStwHIYLA5nJDtNc5Q1TQGiPI
+56zmxyhWHUxNOpqysIDD2Jqk8jJv5c3WPgvsPauhQJsND9W0+rSLj0tV9td0SYlbQt3/Qkx1ZLC
91X0L/oovfsIhbG+9P7FAQvcPDvxRl3aDsvh6nDKHf0pVjATcg/+yi+ng/N6wzkzP16vYONqpE2b
axrpB6FRZRQmTdZnhk3wBnLdDgMErCZQ9ylq4hZLQ5FiHBneB6kwi7ZoBnqCaReTf+EQoSomzeEq
g1C1lnI0Z0MAh5p9l+2TeqLuufDnrNIObhnGuZDn8B7XdumDPN2bYaZY4HQv602PeAiL4kvsxAnX
wnikDCPvxqX1AHbJN4RhnWXOUFwiWNL1nci1fpc9dHL1H5h7hMs5aaYqKqhpruLKp7BV46cGIrmf
I4xWSNYgFgg2OHRFfV25pvyixzhyI9QpDwZD/Aids7OTcE918QGPUnQwSymX/RZ+IfkQdggj7PZ2
Kc4Xm25IgGanrxrs9bbZX1u9ixJ3VSP2Jbx0vtsf4mcpL/5jOXOoCt4KtpTu5CIRjinbtHk03iA+
rvJIfPv5AQBB8pOHfMKsJQt30zrCKAD9kG8W9ymFtrBExpNELe9sQGfy0Fw2abqSdrHgEZqgd0nL
6NKBH4jorG4fl6Wi04Bj4gpBRPjEo/pvquomaG7AZYcxaXTR6l8CuOa5kOUW8cH7tU2aSvWPGOT/
ztuKWYTz4zRyp3tpGyKpciJaNRYqcWkM5xJII+SGKnJWSgmHsbCF9w0Rq/UgmjgDt/fytWkYZ3WJ
BEXMqLu41r1Vd2TbeZdYs2u4IXIqmD+mPqOI47mAD5VWVmY+8eBiD9/8R1zR0c5sGaRkp5ge9aK8
xemfY1Bk5i0NSibTeqDrphWkDfAysXDdc/I1NkEmbWchicsCF2PFSRZuwpUNZfVKPPEld1KYS6Mh
HjhNJtNwTLsy63S9FqceS8kUGjsIxZK1AJ2Ho4PHubuHrhvQqUALHF36O2ay9CEEQOlJvg0+WYsU
EPeJTFexRi7xNHo3ERHF0CWCTbWi3DsFYDevDYIueT6RuUZ1S4BYXehhF49W+52U50QDFCDvTG0w
58+cbEIQUuHpQw16q3Zh2tS6u+J7566Q3J+9l5InOb3d7prp7Hh2cNprgS8GKITKs9ZpYpKPSxDJ
0srdqIKSvdYk4qnrXSB4s3fBmTqbr/bOW08IifByLt7bIU5ffvrMA92JR69fsIp4UyMfe8n1ES1w
F3hkIsHIR5q7IFkQaj7dFFVKrj8lKUfVYPcbrdHaRGiYA4Akmz2U51fsAhtzjjc2Ae2unXpiodjs
2+iudkbAqaUiQNAQ0/Tuuv2KBb/A/1jr/Rdh7INMJY/m/iElw+0rOxU5405/nY9AHhXzSoPZ2Mgq
cI68p3TVL3/rRiATsNxYh8Bg3y+Ta0f80HY92dZuprPF0mEDBuxiKYXqEH/dG/LW1psV6w7sI0I1
IIazkAFAXThd/uB/O2OgLnUZz6KowHw8OuylD6MbnKGaLNvvfYGbqhoId4SPs0bhy+G7WCTFx/Ez
xtZlWLkKExS7wBY2JufVCymi0Bu1gMPGe9Dx1HuSBrDQRLvgTlC28SzoPhujF8o2L3gyeNVJJPAw
UAvSxBc2QFlJ2X1gCuxTCdv9m+S+YkX2cLkLwojH06CeUL4VtM1Dib/uUT4Auz2m+ESBvx/Mgrfc
hgHSymiIbI+6jcEJuZkLrzfSy63mbZgyYkcFfGEIFzHl0FRcWJ70P6RKQU7KDZ7fwPyWY++G6CyB
xVNMxCGUEeo4Rf6msAjaUJIKd/379HGA53n5FGyYriNlY1MctsGmlUI+lIKV/DxyRY+s92xDU+ql
esgmt4WIkRaVMx0j3omE2RiKArUDzRsLiU7BEhUU+dZZq0mn7PJnngglf8WP2DUmXFDo5XEKaITM
N5YyQ8rwWMSDRh5uPQE9JJ+B9mx9c2AFc+XwmXc//4RDqFcuAApMvE6kaXjinNjcsNUNI37DLvZU
L/W3yYch+OmTtE6aX4jEYIYdakxuWFEXlYDeE6s03gD734Xb455vSCrvgU5OuIxszCIrdm9Nifna
u7oo5kiDBpqWfm3BI6Hv/DV398/3vegV1pNCAFKS0msopSCsm/x4iN5z8bX877dujI3RAPg8Hv35
IdsI7NJnUEq6E+LekdTVhGZn9MwX9uB8ZufPPhi/2SX2DHQA8l7YundrFwBUMZMxNUsjs/oZzg5F
OvWLzsGvwSIF/GEhDNLkFw5ZNRSuDLLPfPumNjeGpB9ObYJok3qokGTgWWpDaCbZe+dl3yVp+t25
U/KFZdcOXBkpNLYP352HRsIhvPDOGuw2+MHN8Ps8zVHemBz1/rrtdUBEe9LSIj72Qa2pkppwN/kX
Jawt/UpzYDGOt/1XcK49p1ykS8jT8nXAfufFMoVak6PoRdUAaEZjc60Q12+MSmIlEyYSGPF/3eoG
E1fwY3wDO1w7th0tLHmsVCdhZQQ3iBkARK7zIjw1OUWNzrTOnN31oYydp4HXQ4DjNt3nFHjLKjmW
8pPWUCEMLWBfBc+1m9KQ3vlkvwk8wUZP66g6hXLzrrKJqYRgURXIB75natAt6eG0q0WqxIm+OAl8
aoDB4MuFZZ/axGkQSuF0H/u7hPINY6lmYBoZjVJJOQ3tQJ3HsITiV6cn9WZmd0doPI8lgDkHo2fF
g0iWZIi01XmRiAf83WFvmAxjeF1q9923xBE5ALE4ltqW/0/AbbxRcmv2JyVX2naexChR7BrSmtG6
wR/mS8iDwJvKJ3E9aSQNkBrWPp+Z3LNyXrCpHkDVc3n8EJCAleNEB+zsngF3Jd6i/kinBO2ALNPr
hAu/njbGvnPqNZSTOdQCksRsxOroQ1LKFcRzAmorgJMePCoO1j0NuXhSDfn48lqeZ/d2CTjfAHVi
A6ExRzaTu7fqzn91GwLf6TasIy8sAT/MXWJ2IdTor52dCBBo6eUkXlmjU7NDWOnmu9kA7W9PYcd5
jV/PfHMiCQTEANXMG2OZdOCBwnPllP851+EmPeHowd7vHQA4y4TF92Y6Mihvlwvcy6e1UyPbzcC7
hHhUNV2pbGZIlKNIcq5huLkkvek6yGqghNLAVrSTugOUfcSofAZTTedaJouXhr5Rss0CIAsXF/Jz
Y0/SXyggOozOLDLO+uALwrjo59BNhl2WHl7AJIHh8j/XA97quM6IO/KN+IWj33DIpNJ0udQ1YoeN
MiWYe9rdGzCFEcOWSxA5IsuXhCc6/V3L5A5MOFy5LlExSIHjXo8C+twZ7FHNW7F0Yl6jh1Bn0DVg
GBsWZu2H+1eEd4gh+x/sZdlmT442fXJ0QLCdCBmtCsO4Z6LNequknsmZAvEJdJ8xH2qOIDKkUxfz
EQNIJyoawHa/rIwFK5PbXq5EhcxTlbgJJfJL+AiGZqwAyX/2G/cB1F9VJamNNeZi44VXvM1c7NTk
orcyV8oSaUPjkfMAztA+5yXNjhgc1qT07TRbZ4q6/pmr09Sv1agVxTFB7/rr1xghJWuIkaZaUNZb
qggQoEUZXK4cOIOkZD6ToqjNgpJVeLxfmIK8o1GkgKD2IWBxnO7HDOmOTROhPVvI2QNshuurnRnW
Jaz+9IBVVsCqfKlVUxzbWZzguwL+ymL2GGiv0qB5lArhjqvBdFZw51i8SmB90OuJUAXUBpdp4TSD
HYUarE1lzFrjtqv0Ycw0YtQzYyv4fRU7UANvxHG5PNP5OBUmofSjDWXj9NHSj044wvAYW6JHz29/
WNvsQjwaSFdLI4cePygJYUB7T7/GQIBdAydVhxygTX+bUGXOxwruswgTV+ygoCsbh6aCkgkAA82E
Uw6ttsEz/dWsOvOS0l7pSYWA7tmmHBJzPJl7H0Yj7iSrFKuNhf+D6pKBrJ+36Cajkq0d+lo2lDTB
uBE0WvxGziRKNcditvc7gCBtY1VmdT1VdS687BlKq4vNpr4a12d0lCPPZ1QxQtpEtazpGTXwdU/E
EjZFkkgffX2wOJgjOlCBQjnGsMrtrnxnJ8Jwz/1YH9jAPcmYiQB3hoQ8/sEkt/e3ek6V61eq8sJd
BdHi/XuOiubNZa/q9lbGsJ09CcH5yo6CzJuCN5+ypuUHJWjTf989DZU3yGXu2Y9A36h32m7ieJLX
iDaqIlj70+S8nzrcEMGfK3CLgwNl7ubO/qRxt7t+U3e0qEJUt8aeOutSrK3KMXnPNfcEsXqQjYtl
o/xFJy//jp5WMQU7Sg3jXq4q0uPDcG/oHYCqu3hYSbQVQowhf+8mhtWEngfGzuFOQG+rZqUjpk3G
hCDV9TJNwuSEiZuipTgpODiUGQXvuoFnTvMxos4Uyc+ttJCLsROi/UrZRGh3zq2vnNuCch2noK49
KKzg/Lv331CCOaZYK+DJqlLhuLaDwoFOOYsG5XvaB5LfW14ORQQdtypube0OPW12r1T9ybiUS/hX
gy44UE1pZibWxKR7sPv1yrpWBKF2q/l9MNWFAH4bS9T01lnHTledyuqeScZ4wnow3/IjjZ89Yn39
XR6hQJ1c30686lJ8Hc4C1dtcN0un73DyNkJvE4brlXDfVqBmVEOcBd1rOtgJZHAPM0qScrlgJEUx
DuMNwNS9kATHnx5pAgMzDfdOfnYeVipcKSQVgB6kBSQpnDPCP/YodqmASv4X6HfFVFcxX+YgwEjN
Vk+uX8T+vVA3evYrQOYwKKwGHoLVt34WlIj1qSTIq0pZNzKO8gq6jYxUAkHAQtayD4jes6lzqkSV
lfMNxZW4pCox2ArWrxCFlh/Xb+nyn22hoZUJsYd2HYc1/LfAnCGcOPUoZ9jI4m5e5aZCT0Ceuhw8
NmW9beeLdtTSN+L/bPM+YH/wDNkOvPLSTjjuc56VBHyeVaBKaJQr1C/rHhBuWwZPRzTaTRGpqg5t
m/WSqtSVm162dyW83QGmVrdTm1zCx+SKI5TF+KzCPAuhvnq3JTfKJiDobUvW79sxZjtqt4CRlVr+
i90Pql5aP0YNDgRf64AL9LmkkmQzJE325ag7M/QpCwUUo8oXgn9RYs0ACAMwMLgjTBEXzu9F5UF7
N/6W8C2c3xUAF58YCgUR2a+IeBI5wcuvz6US+V7bcQEvz4SuU9JAP+DwSuZm8TP3PGSnufLq8pP0
HatRGCcNJs5pA3wNzMgBKQpr6myI3OPWT53inbzV0flCR6w176P9M7XyaBRtggb3k767iT5Tz7jb
lVMjOKdMzWQ7bwI8OiLxNoVjA0NTaXjnOnGMi7BpfscaKKP9VEO9T0f7hDCkkxUx7XPxZ1P5Hvsp
GGdNd1D3GboGqpWMOMVWiMSgT81b9ultsicUxced5E3LkwvYZamIvMiPuiXTDiTNUDBb+nuZRVsg
Ka2Q1s1iRA/GjNKHfBK/mihIbIR/clZvXSni+cu8e8h2SepTJGJUckhMrsmLVJBr0iRZWqQuQwna
saaWEWmOh9c9PpQhgC3VUxwjBJkys8dEOGqXeiKAQpQx3JQMD3MvR3XPNpYndygLaRIYGQnK2wbs
lZOYjaDD7AuusCo7FcwKtu2n8REZFxS55A9CmTTkTPrFiiotGLa2LUoQ6WM04TvenleR4ix4TFuF
1eNr6Msg1N1u5KoqFDbcd38TwuqC59Sm/dRys8ffhCRSnHK7uC5BzV687u2SZHsWMtbjAJpOhZoI
mA8/mimi2Dqb0Scdi9LJZgboWKerGEHSBAIFePfn/uDcw1Km0YQNYYaPmdROSi2s8cF2yySsBcsg
VNCwQx13MStjyKhYftHCOO8PEUfuUdA9m7MGxz+XTnMZJRL++8DPHMxfb7r6L32EVH6MShHteSTU
61qStbXxcZQD3TLjAnrdnnSZf15snLMBcevxx/UWBrPvunCIPlElsulp1HFE/IOZW3yCH2cmNcuC
fCzLLlT2leFaJ4E4Y6XgvY1I4Dh3KanO2bM1LIExUN+G/D4/xonxpjvCpC2h8Vqv/NtXkFA6ZWfD
P50IZStFk1BrW5skYaLY2rc63+oLTI4q3oO6KAAEc0ZkT6TpT+B5ChvkV7ASBbWCui7iRkmagI5e
v/rir90tdWktdfiCrnY02l9TpEW45jg+X0z5/GCCOyPNH9AaEAVtCDdRsNuZpKBzz6w+5ne0ms60
sfILtfQAn/Vly6Z/8VyUM3A8J3FDwqI8Tm+2E17K7AKoYQuXNGLQF7+GjpkSE0RQgVijpXL/Q1Ba
jruF/wg/ATOVcHSi7rrWgJkFw1LHypOqZLsPT81L8nOhiEMtZczsRLFvhiuy2wUEX8nQrfGGiudX
FVW+yFUV6NtpsiTbRyajr7IMTwOqcPFqkL+FWzoXZezApUg2/WBd4zicdzcYPgFJvLPERkhUeGJX
YLooVqdhp07T8v+VuvyRs7RqMB0oqrgH391jfLqU2UR8W739Zzz2AQxOyDXFFVRhSUgSWZii0DMh
Z5t6NkIwsQLRbfKzAhCGgy8oYLIBRHIE1yTMe+Qjo/mQRNI9KiBSQUGpojyZGiJZ5ZLoOWy/KNFi
+tBL85nnY90xjNl5jKiRIJ9IloMLCee1YiFdD1hnodqw8Ulk52pi0G5p7d6a+FhNLEKNHoSp1OaH
XoCDrwcpLf3Cpgiqzn/TtX5NBKh53GfQgyVwZO+EZhdVIu0Q+Db+6xTyiQGh62ILX0el0xhYn6nQ
KTAH6NFBU5apHfj5dbzZ2ItWBYtBx2DDbgXqS+DUY4DbVdH7fvL3R0tTkWrTPy6i9W4YDyqUs3ph
T3N5Fi21hMITgCk1o/mFkDKL0Rrlmjl6oRQJ/j84WHbTlOf3JJM4ha9wq/8RN1pKUBbLeeiT9iYQ
s2U1h/aXPI5UxeJ+r+/70SHN6ZCqn/Q+ImJQxuq6He0rvYcCTQMy2pqkk8hn2EOIRiafQqhzAY9U
9BPZi3JbjUKAubRDXgoHpfl+ulXsYfpYrqoj2Rn8DzoUadp5fTV7SniQ8SVnDauDvzf2l3584InE
YaHkBIiK4RGPZI4M9xASfU17twiWBUbyVi4mCuttJmnLp3gvh2pbvSYU/hxfKxp5XiDmU7SUBmCp
DgmutJRoC7eGVCc1Ik/KteBYmtOJ7+M08/14p+U5pGiP6GugOyy/WI+yDLz/Pp9g3Sq4eZgrpSmD
1/NnfzAXZufNfL15dmd9btrUm17zTEsdS4faivFP0AteOyIsD05bRaWwx2k3vdhaPT33x1BKQYqg
p+wxSV1meuvlJsfwGSLfOM6gLH7QYocq9fsmrXV6EDgmtYyAMutvINvGYtrcLcHXl38dVsE9l9n0
IEFEyhoJ1tP6hvNW2k/inbuLGRc0PJFTQ6YbEgyNOCbGCZKIMrDSxwM1SXjcHfBHIBNp2kr51GnZ
AzZ3To6o4f3AgOFlCYxk2zgN9SPeVgcGHxuxbLctmOyKXBgznuDmYBI4UwxUhVy64sagsOzx/AN6
DuIo8kAGl02+6OYdQnRrhP1D6qFAhEWLaItLJIQmZxAgRcCktnUh3zGO0OqiFEoLZs+uMk4dMD6E
m0S6wztmYl+GctPMeqdhwaiLsmxoojMnXi0E8huLfZ/QaXfdfiG9ciLy4z/RsCExAQ3B5H1tRyTg
Pthe4Ztky91kU1PEqr1fpjyk7YlupRSeN/kjKQxFNna4F6szVZgbNNiSdOwrdyevC+5AkUkQmBX0
w8iB+g9VNDDzjOanTQHQB4oTNX9PcoZVQbz7qWU7F6jkmhNBbsb/Mlp7KcZ8QnztqQwvyBn4d8dd
yyeUHexOQu5/YmX/J+WOjPuUlyCJirh5XTPysayd/Rpl0urir2gObCTqucYR7uznotdp/chhhyWS
Y/M+r0vzKndwg8aaMS4XPQi30Du5bzbwaJqxSsy6F/p0Vu/QT4ET2i2+AmrW0v6p/k0OHsj4XLtY
Cf5CcqeWA3w0hxai0jrGwF+zg0UpOTjPTfmM3Z4pQiLW3gTP/TyVHe7ks8ac64uP+QKCNQlj5Jbk
JqVWYRzWGK9+WK4mUXjYJqDsyl5ZMb+mfnDy0V5GfnyGknd6vGGXsxGzM617YHyxf1kS9KglOu7W
osE3+6/urtHsuiWLMZqIp+1h9+cgO3BLk01Yx3MkjfJWiOjEk2vcNNgwWBTR3OnlRkvXLEGHEsqk
ihM7vIvt/O73e1SBTvPf5BSJodgBkNtZbmHkJzAT4d9mn2l5w7HjEkKIwaRoFbkjf9WQCL8xxvk1
TlhmCWqJYuuGKBPVpQkXOjjT903DEysoWZDHGG18eDNLblXm4X/88Ezt/od60yngmgmjolK1d88H
kAwXudd7t7k6Lm2ikwQ8jHC8fP4RriOXxaTwai8otbwo+I2B0R8KtwgOLTZ/5a7jGmcp8jPIIo2a
/BhejjZDXNEU7Q1EfBYG9dItrFnD50JybAUWP0hwSOvcavMOx86UxGuxd2tRuHAJep8skD7JFjWS
ck95Pz59Vjdmk4BpCvF7Kg7N42hiiaRrF6LtyKFl5emSYIankj9M3oAwxaw+UC1OVbzrqQD3w81Z
JrHxjmC3uoXbq5ILLjA/YniVNPmaDgzuqJxNOhiMEJIJ4fiOH66KJiQ61pKxfalDhcDOh386W4zw
uNhWFdya+Pa69LkJApNzTQPxnzkRKC1KwEx6KbEDShjNFTLfiXGtm1xDB1mXN4o68+Y0LYZaKfht
DUx2CxD8ynMUzj1avZXecKVgDupWkA3StHswuCS5cJR0KDOTh7mvvvaJQOIMsaBad5cm86xhE4cF
5jcSri49d7JqQ/1gRLk39RylIb55FzNS8lmJ8k8sw/uzfKk28EyjDel550xvjrfLx6Pn7SqMm3ly
EW3VoRdW+bXePNsqrxslR8IiEPZSu3NCPgrH9hOKWxT6Chkitg5aG0HJaT//H2BlvrlhL9A+rCDO
WBokL0dP7mpp1I2OLwhD49NLKImr36R2DL/qjzuMxa1TUd9+n/BFKJbLnCkVaUqd3GVsvv2ILsZl
ORioeVxMG7Jd99zvQLdRuOxT5F0L0ED99c7Q41I6hnMw37MA56wlrDLU1F6Gc6rkniSF1b5kvF3d
HjnZrTVn+ilq1+JyqbRfxG4Is/osoxXimKpCWREfh/Kt6NCKomWh8oDazLjWILLtGuHlG32L+BNq
dUoDrwqLVIDTn8tNKGJqtTnkoIMk5P0dSAGTQ1zlm1y1/NPi1hJ+pNUjaGlFLITRVqOVF0hIHZKt
LOyKCJJVhZDtB8nbVwEvLcRsS2RVoe35ZPjOi04LIQETjb2xkvRDjNEjn4wx6azZtBvsbh/mSPF7
qojQLhiI3AfBDNCmXBGIp5Xfpd+k7n9iQXgOm7YY3+YSEljvylQjOSCz0pB2IeJLoSAW6dfcQ0yu
ox2NC5yqU66fGEPhHEii27u5Wzu2m152LbYGuvg/6lQifiyIB5vcdFxoxrTHYeEFYNjddzx87aqX
7zPwEBfeFI+GmxPVGzqEdf17K3ZOUx5DLms7lmKVoCkYkdWSr940JeY7vuMDipAY0tN+qVA/HRys
6GHffxDx/ZUr/9PzhQTrS+udDNAcT+FBfmdRdPli2FWasvdwaL5pru3RQQXe341JVyp3AgonMYhd
lHt4WPVbvSyC1mqPPiowXN5kF2TBgVs529tqkk8+7dBTSKG4Ev4YrNN9Tp+d8mIySrngm26KAcrE
zI8SB8wq1Ja3hbyWvjGnNuuMq2cOzD1sPVX4yc/QyuoshBlyMBbfyua64bw7FQ84snvz4DakjC2H
Vgb4hc2iMVyElKU0ZNMfvkPKUTTIAaHmQwOmh4H9+cEGHO/QObKJx3a04kRL1SR6ONUe4/ydaeXJ
SP/FElOYLbBm8mgPr9aKvrqBvkoa20ZGp1mKmugeYctVTJxvzTP057AaPJPdxsTlfCOGoD/frWQw
zZhxrIV5OFnOlNeFGzwhV8xHE2E3HLjy5O3jihPEWlUjEbDE69hXeB+MMj6dLAOCgkjlnOLRl/nO
L3bnwDS+t8K7mTXT/pVfKp6EJ8smqPKjY38d2c5tev8kBJiMitPP1IzCAm2P0e71z435nh1E1Kyv
lyR91DCAxnUNguvkIx8f4hH/MSoK5jjc44ceivfHyNYfELSBMLKVU+/hK53jxtTq1M6MHGU+DJx9
MqmTCkn5LjQZpRCt+ZPlNVDM4Lt6U0N1hvgwDuHy+faBCvc3Hc5EMRCZOW70ZktSMorpzip9Tr2F
m5QEjZipXhjbyIa8kfx98udz6SAe31jhO6VtymEmZs3R2gk4FcEJkaE8fgCH0IhwF90lVq033d/d
nliM9fy/B3nOjSTR0FrhX9DEThvhyCod/wqdsfJRdpVDbiPcSX/M6G/ltF+9sxWkcg+QUIKFnsxS
IKpsCNE/r985QTw5SQcnUzg1xGIJ7uc3D6orFEXPrchiVXSllJtsEsoMhR+I/ArMboMKqmmR0Vv0
EQOAGd2gGU1tekr33L0qlqjIX5bZ0aeKos8vxoVAd2EVT7tYPn7F/PEpqiJD+JBN5/MrL5F7htuu
DjY5hkpt3Aadq24GFlzP8htB5DVsbj7s5s0MzjpTwXMb/D1FwlQ/dFCkKh60JfFYYUuFCOj0Wgbf
XeF6+BfYYsOO07rIskv5otcPov66V2UxniMoe2+Ft+T3YdsCBDjSsA9o/3ooTXJj0ki5zUE7M+cc
w+1RL7k0QM/yYwP4/5DsdE3q7yw40fIMzKl3RWLxw+dffppOwFp3uEl71AIYtARLm8NRwujNv42U
+wHpOGQL/73vUsKl7PNWi4EmHKFZEKvGi8u41PKTl7ZOl6x8u8MsMMrBWC01rpo41v5C62QymwnD
aZqN1ZirCCmdfWURexqQiM2yCNZhJE+GoxZ97B8fvSow2wegqLKZyyviTiImx21H3k8vE8I4Z0Z8
N7go7MrEoiouPnub07dMFS9NrbnN2TqRBRGVibf+YirocsZtmp4rPnBx7YhfRxUfa66NbAGomRc1
IBFe4fpPFPOAOywkU0tIlB4PJX5iXooc/j9lOtRn0DCMqe0R+cDwEbKcz91DuBeuE1Yuq/z2yrKj
EC8AGb8CCggTT+HUfogdNgrH+POQcDDJYrbyvUmZNUcgLOfGFxsF3JDQfM5v3m9L25y+Zi17zwYo
+lHcZoltpMYzLjVuHkMD7+HiJkLrNdFVmOw2zuJ7b/kVsQy8w6kC+g8dRrJ8myTHyhVevM8LHetH
K+srFra2VUIyGBxPn6L+2iKeSI9EUZx7rkfunxlyFuAChNc4Q4woO/VIvYH/tTonXoCnh+Zo6X0T
3e+J2zZcVFX0XwMDZUPcv4Od/fOS3fdM/Wn6Ab29BB+5M/0ilGdrzNf4rMPQUfE2LL/vhnoXUJSA
5jLxH3mUt9BLUPgbj7aM1+KAVEJu2+81xPh03qkXGoBh+KSuyy1F3YphupoEeT6gVik1QUqWC+h3
kXBevIkfSzEZ+ttsYfgx6vDMTsJb/FLNdPLB6aCmu9QXawaNJygXRtOZ+CF4Qmy+ITqDM2qeDAf3
9YA3rjrZHY3rj+XZcw/j1MU/HHAEwZjZyJdDzzC1LnEUzEmKnUKWaCZo5aodFJjh7Qs6m6IMeRrz
ZTicMtUwicKOASSHEba5w8RLbGtojjc3yiFCBGWd77VpBbEo5ToTusjmXGMxwjcNgGMwqRu0R0KM
R0XREI6mJAZSb5Q73ZyKCRQcz7jPEOf+N5Qb7x93Yz0cwcuvIRLtje+7A7nXP+UfAS3EWz+Axq8a
JAIwR4AfR9sXSmKlB+TyJONPQLIWEA+vLSLoUAmoRup5jKyGno5ESLd9T44jJg3mHp/5HqAurtve
lo/hioKxQCLcRtr7pOchZaM0XBIFvgGCWa417hTaCkjppFlSSTPjk/J+CHKifSwLAHDO76cG/tWr
+p7xrX49JAUiP1IiDuk/3UEqb3jMiWCAf+gv/zTQ/xbf4AeiXojHLiLU3sRIDC+fT37Pd2Ii1+EE
3gf43h8Wa9LJKox338MSW5aJw2jsQAv8PiAllB4ZARIitmxd4oPPoe6jj9xmFAXONdcx6O/gm2ED
CKptvCssT35CM3FZbN6ivvVDljuEBTyY7/qzgxorNpqavA6cfbbIhwf1futFPyQ3VidD+lpLYXEQ
9q2BTmqwGba5rkariBSeUEXpK+PVO1f4J9oyEgForc8yR7zVb/orcbR9d8nEH7VqxZ8LNDBkeUK6
rMw3uK0WSmi73BSsHwcKekPhaf1UuzGIj48j/9UORHLy+UdJYi6smXB8tCL3Pvc76G2yDl+S9qgj
YxfGmwMt+yCAhAzr5sYEBjrFJ1bYYM8006QthBNdPOfZ2cNYbd/jb8YcZMKpeqoy/hD7tJ1H5lYg
KmJ8TMmb4TCAjI9o83QGKPrEbPg3LepkkKPREmnkspGnfkFCr7kcms5hJLNyUoZ/q/GFcj9QfwkF
RwGMgux5qyt2ySDpDE9fiz7lgdNb80UE6R0eyP2iMQFDiKwzBawzf/KEVax7IIJuS0DycuUfUfBp
piIXGB1TahOLxlbRzY3m+rN4H9swciftAO3iufYgVZQUX1k8a9FD57aOLPpH9OhVGgWnAHTu92U8
h0/fMzoYpl0zMux/3JuvUwqsw976A6z8u86sQpYe5Wxw9w19c6cfgIJ/yVIDZsupWLGEoC0VoTY6
lWOmvyrDzvc2F/wWyCo4updbGMjkfaaN6lmaYCMQtX92TVMrXssNJbnHBf1BzFFQvuLryiNJWNkC
h9bkPdq78QXGBlz5N/sBMDF8L+t0nyEq

`protect end_protected

