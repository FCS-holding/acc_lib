��/  ��Q(���]G%�B�C��G�1�*�$�^�Z��%�������[�Wq�~`�	v�.@s�Yꥱ��+[q�~�����h\x�W�f��O�盁G{b�]���i {����~.q}<�	���`�� �)���(�c�,��e�ط�>�KE��u�ɕR\Q�YL���PB����m�8� ��_�LJ���6R�vݼ�����b<�"�i��7k��n�.[����i�P.Ǚ������-:O?}��԰}DHK8�19v\P�X���xy�g�PZ6�O���$��`kŎ֧X�z	���ܶRm�(44�ŏm��ؽ"Es����UG��B��hz��B���;��??;uئ ~�ʖQ�|������5Db����݀���vs��$b)yUoHH�:`]Y�����u�|Π�fYKH�Y;�O����t������PU�Οt�/�Ԝh�Ī1Xt���Ӱp7 mɜ�̺3����aS�!)}�몈5;J?����ޠܬ��Î���W��MňA5RZ�������]��`����F�#�[�f��:3�P�m�
��(C�ht"�^0^sbх�#��ʇ�C�ԛQm�瘞5���#X$US��~��@���-斕�]�Q�_P��]�l	¼�Pq��5������d׋��"� �L�r�P՝����	�'�.��Br3X����&�g�6�w�gt�Yc�$��ב��9����C:��k��x~W���/*�촯�᪥�u{�Xgq p�� q�<YE1�=-(�9ݦ?ejS��ҋ�u����dO��M�q���ixLF����VޱB �u`}�ВB��/Bgn�%V���~k!�|�'髯�s�{����46��	��J՚)�T9��	ƺ.�_ζ�Dbs_(��h��|6���%�^t�c��=+�����-D%���Nٗ�?���h7+���hз	�Xf��� o;��+[@�
����s7����r!��]�����[�S����Z�Ө���)�ZY9�`����<Vj��h9�y�Q��[g<�s����ҩWz�cEui^h$�u�������'��� hAo�٥P�=�U���Q[��$Y
%*�G��J�nT�� �?�j�%d�� #���/��ˋjw���T����r{�]�;�� ?	y��QX�%Lt�ٴ2�!q�f�t�m�!�H����S��?��[Y ���A��� _T@w���G���\c~0��p,��X�>��ۮ����=M+v�3��G�m����jD���JG��5�D�}�NL�����4�_,eS]��ԫ�nS'SP��ܬ��6�ɼ���;�@�[͑�<ώ`�O3��Y=Rx��Y9��P�I�D�&O#/�r��(�o�۹�)�V������x���In��؍ɺ|����q����Z��)T�5�R��;"�zs�vl�N�����%qI<!7�!U�v���=��VuP81���[p����{��s�Ǵ}���l��yCܔ�R�ot�������+��d�6؅��`,z:Ȭ<�vƎF�4b��7/���P��M���c\���>&p2�����8�?F�D�����5���MڦRU���=�q݀�R�:iـ��*�{@9X4�J�+��%4�Wp�i2#�T�)�y�|�A����!�߹i�_K!�_ĕݩ<��n��L����� iT���&��VAE��0+ԓm�q��X�?Yo�s��3��*��ͣ�B��;t�����|霳5[ܣ�H��IGpsa/p���� �qs1B;F:��I��NN�bs �p� W�F��B�:�4[�}�+F�˛�� ��n">��;e�S�4M�H�ț��VX��3�ǰ�|k+��\(k��9��`�x�GF�����.C�aŵ�V��)͡3��=�2B��~�K�8+&ڒ��;��4�#���P���H�����^P깨�U��'��d�H�E��|Dd�ik�mB�`z�L�ϖ�˾�4�q��L8��T.i>�&O��vi
pTT�J�.�}�	,߿���(s/��FP�yM�gWnҍ��$dg��{˓K n.�+g*Qp��P�4_����m-��7�A�.��?2^5i�`6�|HɄ�o}����rY�:�@[���G�#��,6��U�Y6
��g���Cړ?5�.jA>����L�Y���f+wq�>M8�<?���l����]�|��3��:-�n�}�x#���$��A�]x����wp�y��Yf�]�;�N!��n���T�$K��sK��}��1)�{ǿ� ׿!G�6��T4�y��^x��g�Q�eB�g�d�<���\S�)�Z+����v���$�%��!�=�~�މf����K����B=�i�{���&|�"�[HR-3�*����L3����o���`*����	��T$����h�Nv�im�_g*��Q�{x~>�!����IKH�|��o�Dt7���K�$�T��i�����w�+� ��Y�[��3���0	���k���Wh㵉���+a����}'�-����l���@Sv'(���yM�Vؚ�3h6�9S�F b�h��UZ�쁽��uix���E�<Z���C�Z�z�#۹��c%�K�Y\�n��xҘgc�F�}�0��6��ǒ�������l3o���sqK���NC��At���7�K5�ً�@�8�l��G��4[�����k15�ͦ�n��~�ƫ`�Y�l�G�]z�+���2�⧺G��V�eD�]r����>p����,A`�;;W�{AA�����nU�ݻ�C�[��l�&��.wn'H�����`oE�&�z�@����D�e�B�K��b�25�/��,�9��,�a�l%Հ]F��^�[5Gpc9k���d���l�����s�|)]9VlB�!h��Z�f�����i��7��fU����LnQ�z�X6�Q%x��8��V`R����<m����˷��O:��Q�*hٛG��Z1��a`��0vZ-s2��B�t���v<w�޾s�4�3����}y������7}������{�|BD`��ݞ_��@�/o�>�Z�<�Y����Ĺ��ȹH�ϣݧAK�Y��R>޽��x��v� ��e� i5N+�]�'v�$%����t�4�U�c[j9��@
U��#��.50q�]�,ա��ڎ>����g�NnX�@�t+%��ȫAk��	m���N�d"ke���]��� 8��O�{����wT0' duv��㡍+rT��2�� �x�����"��%ӗe�4��x$Q.T)/{���R=���q�y��SӍC��p`[;���qVX�@��w�!�"�t��Rb��x��@��Q�!�et�Xޞ��&d�=�.��rͩyZh"�jD�_���q3M� ��2�+׆�K[I�Q�9�<֗^��
y�iX��o�u�����pY�cLaн�__r��A1X�CB���!����$7����@R��X��E�m�P��QT�QZxZtV�Ʊ/F!n��pƚ�6g����UV��gA�w)���2x�I��E2}���Ό�V�CHf����ߪP�B�C���x~�����X���3y�O���yW#��VUEU:m��:�~�"�!�!�.
��k�8c�b2���8>�2p���4�њN��'��nx60���G�k5�o��CS��f�zo����O:��B��dT�؜�Bk+���ʨT6�`�_�q�S���o��Ƭw��t�Y	�2��Wip5KUP��}����6�tbvpaÖ�^/O1:��?\^rٔ�5�{T�[�]�s��{va�� \NBF+��1�-�!�4 ��b���T��Y��k�^�&�7b�+	sdUX:&U��2�Ct�y�{T Fa���a��*`����������C��41a~�`f���h��^Dj<9Y���+=��_8򱏓�w��ڤ��E�
��n���
80���5M$��|i�ҁo� ;��ޛ�p��[}M���؇·�����E��,^�"�x�L�cK#��|]~^����-슔2ɫ(G�A9��S2/C����K.�pe�@j�@|aTgc@雿�B1�q�y,�&f�T˫,��3�?����V(�0�~�ꏜ�� %fC��ٸ��EZ�c$;�ݣsw�QE��r��W���'�U���4�DN���RD�^�~A�Bq/8X��eԍ�bx���f�9"��^~�����qu�^C4�yd�v|�Pe��o�(��C_c��k:B�΅͓'��!B���z� �������d���;�\c�(���9�")и�^\l,����}��H���F������b\���~j>%��@�W�]���}���*�6���F�y�(&8�@_t�]"+��\��m�������y�obu1JczypQ��[X��+�/Rؙ-�8ܯ���}���_��ucsЀ��\�"�&Mp}�>c�А�}�|H�����ҽ��D뇊Hz3��ϥ2���CȘ����d���P��h�(ɚh�
y��� �?X����m��[aE:zǃTB�\M���Ze������G�K���fH����2R�k�KlI������`��\[ӡBmml��Ţ\Z-"��w�_z{���m����8|���/rd��V��q/P8��Yz�JZ����w�������L���}j�b��32=��5R3�@�"��{Ef37gB���ـEՐzi"��<�'��ɴ�k�WU�Di�����~F:���������.��
辏���K��[�7y��m�i1����BH�ߊb����F��v�>a�^�r:���S��� .����Ui{k�>�3�0C�f��^/��:`�����4�J>�p�d���>��Ꭸ4�I�o��)]y|�#�H�hZ�&��V�s��Г�rf�������g��n�)sr麲\�HA ha�[�޽˲���eY�ł}n��-I��4g�'#^36Ϯ�R|�FQ�.	Y2�F��G�]�F�07p:÷�ւ��v7�ۮnQr4��_c倞�ȓ:���=��1�W����au}�cZ*��B��>��&����uH�V��?�k�+��� �ߣ�5����g�eF�-d��s�B�_���=��������JX�I~�h� ���E�`�bOQ�.�5��Y���dytl�ulL��f�� �+��>{}�y9]��=�����{�����_k?W����hN��CU��k5�C߁�[���������1�/-����p��1w��Vj�P�{0E��Պ%���fv[�Wb(42�L4�X��
j� w�5>r�V�\i���(�F�� D�F6$�O9�l?���'��迾U�r�~z/�j�J�?�G���9�������}ؘ�h�R�'�Ch�<Y�����g�#�~���@��"��.GGkU|V��v0�>�-�Y�����2�3-(�R���B~��.R��TD�CŹ�bG�?T!'L}2��鎫�.J�9:h*�IfH��F�:-	l�!�T��i؁t��L�Ȅ�~�EZ<��)��k� .O!-Ѥ����fi�DBV��s��C2�;)t���x�mS�ka� ùs���c9��J��J����V��S�g����ۢ�#а���/�Ҭ��+�:X�?���=󟚒��򸸹�ɜ��{0g~+�rD�*�J��r�h�r'Ձ��g�o�^�͢�n�#�{��L�8cs٣��^b��A��|�h���)n�M�\��v�i9��m��qO��vS���:��t�M���qP�G�qd޺5��l�$|Q�b?�Pp���6�����rPO�˝^I�C�&���2T#�/�]f����\�l(��~s���e��t�ENB]���%W�����ۀ8_æ��[V��cG��IŻ�ƋT� �y��0�O2k�I��6X�sM���}d�i��`��K[�ب�`e	Ąpy��8��]d���nπ���i⮏��J4>���4�`	}v��s%�ݒ $6�����:��/�$��h�=��{z�f��+AX�z|��{�~���X��j���왚�m�r=�tq�A����g�C7Hm?��yx��x�n�,\m@ZWw;�;�l̒�s�#,ۑ����0:Y���Z^���5��aF��f�U����h��bN�"�j���8ݜH�"o��ܓ|�<�L�x��-�E�"ܣZkeir�����Oxu{>�薓��RU�s:}��vG8&l*�k�n��a
�H��l��'pd�0x���4sf����S)dr��6T��Gg��.�,���O�ۃ�O��Dlܱi��j�Ok�<H�h�D���9�8��4d��=�x�a��Qq0PI9�m@��c��ʇo�	��׾��������K�< �t�w�`��/��"ί"�f�J^�,Qc�͊B1JAp
t~�f�_��U�TjZ&�VDڟW,�D+[�Ip��DM�ݿ��Ѝ�7#�ॄ�]���P�5A;)�2H��A,�9�������@h
Ό�0��A�K��o�bsR�k�b�	`��M�T�X�mmY9./%T�� ��Df���~)�&��i�>S�G�GǾ����-�q!N�pA�S5~yt	U�����	�l�v�w�n?����Z�Mwv�7�J���P�����a��.b�J�0�D�+�$n�G���\�"	�m5�ʋ~����3�%�G��<��
c4t�pGdr�JM���}���<g�U�&j1w�-�l7*ӱ�H{V"���
�G�9r2[}� ]�	K��wΐi���!�AT`��S��EGe(߱#�R�,��V�wk������XY],@Η���?r�~��j�b�w��G�4�r\
��#�ZS�)���iu��AVO8lm}3��=�� �O?4���jG4��(�C����VꞲ9��~k�RY'���RP��Ia@]�i��{�j���.ns��&�NH��ӛaKF��&�r|?��'sT�f�H��Q���p6���B���_;�p���_�Ƀ�`����2��	jn9��s���������}y)���ʧ���m�`0�)}},�䆜����v���=:B�p�����v�xH;@�Ok����HzX|΂�b/ R9	�ĞG��$�V,b(ry�t���N>�9����7ё/�������N�֓\կ��2(���|'�*=�ߠ��R�7���u�BXt9ϐ4?������-���y�\����J#�haO�N�r���1�{�V��	�O��\��Y�3�q�X�t\��w��:w�6�8��'�
y �KccH7�˸t7�F�@�dX��&�n��+l�̎9hF6fz���U<¿�'���H�`��)��vAcEa&A)+��vA�eg����^2�4��WO3�o�QY&J�C��y�=�����h�a�jE{��2M"��ױ�D"���$�1�ػ����7ɺ�K�b{��|r�C�bGȠ�C��J ԊQD���7�B��*
���_+(s R译a�nv4�R���w��:{z��SOs~�ҥ8��mO���<8�ζ7��oMOu}V�&�+.�8�f��*q�?�.|�:0�<)�)��70V�	P��GSj6|ȧKZ�Ig��{;�W#s���^oZ�'��)����������'`��$�D��_K��I��R�錠J�ˤ��<�dU������rً���X�D$��~�"d��b��3�3A"p�(��'��}��n�u.[\0�LH-��뻋
�ehKK6��F��D��oϽ%"�� ����%���ă�xҾ��AH�M4�T���iR�LB���S��V��^J�
�9��R���A �������A�(|�	�j�����q��l�j(���7!Y��*9�(n��P��k�M�|Dcs��.�(_v���.�!On��H��iS]���?l:��9��=�OIΎ0��Q�?$�ȅR��VZv�?��	v���`uJ��4�� ���RJg���óeb�4�����['S����R{�LE�% �f>c!�����������à�45A�Ȭ$�I�l����]،,�6�׸�ṯ�GĄh�C�B�ݱ��lo���&M~���	;��
�&c�*�nZ��Cĝ=*_�qͰ�����4�co8��'&�Վ)�Dgk4�%��Z �V\p� "n����a��^_JK�@��}�r�����p�go[�+��(�*��ysXcx��p��%?
�Cע��pp���d�4-�gӢ�$|w�T�ai��=�v�<�L1O���눹o�����wi��E�=���)�{:�Z�dS��V�pͰ(�:-G , i-�B���o����>���K�2���</^�SUkMG���bȦ۟�p2J:ݹ����� �d���
�p���|�<��Y�я{Y�U'ouQ��S����o��L���SrJ�J���'�-
�v�@���۷�a�S|��*.F��ډ�l逎���[�*�Y�y�6C��X5�� �j��؍�ih�~�q7���YJ�����G'2�-��Qm�ȕ��g��O��
c����i!;ėw�]B ���qI�%v�q� J�p�A]�.5�I~�ze�7�קh������a��Xe~f}�f�\	��if��I�/Nu �{N��+g
�Аv) �3���!K�rA�� [�K�ۼ_Ԝ�H��B<z,)D�`�~�;�t�R�������'u�$n� n=�sb���Ż�ӝ�s�YvM�A8�����)΁1;A�h��}z	`����	�;����;�R��E���\�fe�v]Ro�$�0��u��[��>VЬ��x�t���&�ɟ�)%l��Y$ڛK��.��^��Y��!~�-���;+~�H�<[���D�z��J��� &	}�:��[ҍ[ȯw0s̴A�Ñ-��^����F���������&�W�m�P�����d���̯�!Zm �Q����M��i�`�~��y���ѢC0�?�,L���M	��cb�1�y��j��e�?ќbU��4�N���K���aW ���J7=�l
�讟��7�j����Pሳ���&��u"�$��K޼D 
��:}N���7���Y����
��$�*TC�t_˿bQ�R3`���ύ�N��
�'x�E��o��ڏ7����o� 2���>q�?��J˟��G���~2��#t�5\(����2B$Һ�z\r��� $��J}S�N%��|<

5�1�!5�Y�5��n��]d�8(̈́\�f�4_���n�����4���s&�@����j��0b}�d*�.!�gx��=�)�Q�q�);_���Btg8�w<�:�qv��<���n��EY��-ß@ǣ�89~1J�:T�g����J6\֍���dE��y��01���(�$	�77¸�%r�gƠ>�y���r�o$<�@�����<Z�\+���I)��6� ��uda�r��D�l����hl%R��Q4��Σ����Lz��Հn�K2�� *�p���G�d��p�w�,ʅ�7�?ټΫL ���i��f��B���Y��0�!�WT�x1or��D�/:v�� ���ڢ�R;l����̀Sb-��ѣ����s� ��Ș%�u��t����}mР&�`�W���u<�p�y��יz��t����7�'> V��`^�kF^3��Z�9Z�r\�+C"��n���&�7�
�탪����@0	������u����<6���D��	F�U�{��Oڼd�C����	�?|ݤ5�\��Ɂ)��-����c1����EJ�j��s�pr���]����;�t ]�@ ���	�6&���>
�/l��8n,�<WfU�Y~���u��g&6ԋ1V� ���{0i�(�}{�z�
� ��g��ʻ������Yi< |#����Y�;}�
,��%����Z`l���7��/퟊�N���&2)� �p;��\\慹L�y�zU!���rv��B�	$�_!��^��<��$6�vAz�O�_�d��Sm�)ҡ�v�������BF���V�q��x��"�ޓ$�Y����O��q�X+�TN}~�Sd�
Y�Œt�\6��@��栥W�����=]\�#%� {M��ی��5G�o�@�n�cׁ��=]!<D�&D<��%��f �C���!A6	l��o�%�AQ��t�ۖh}��E�2�V���֖�R��^_����e;ɒH`�?M�;�Ʌv�V3.��0��81.��*a|�u��K0�5a��k��]�� q6�m�ܬo�Ka�+�+
x�g�a���U�Q�7M�:߶�$�>�s�t�^S�m�.�0��Z��rF9-I��ŧ{�ua���;�f<���X�p��(�gs�?�T�V�����"��]�mbT6�'��7o��E�u4wM<�畦PF��y���r"�fX�q��6��4^��Q�mp��إ���f��Ba���#bj�� ��.,���`�� "�Z��ԩ�'�����d�YQ�+�����"��F�<�֫EE�T�+͘��θ.��$����[� 01�-���SQ�p��_ŹF�q� �hy����^жs�Z�cS��[3�	}a�m����ڤ,o$��U�Q�'��x�[��E�Gx|u ��րF��?D�����.� |�kS����[HӃ�Z��ӃS|�`�겎k��B&���s�48q��6�b�j	�7W�$�S�].RUb"\���h��	�a��[������vJ����'�;ؓ�VՐ/�f��pcND�LQ0�����+�\��"���h���7]U�M�"j>k������`��"d��2(6�rܛ͵|�ҙ�Q��G�۹�M����6�`�ܚ5I��3$�q������ ��]�e�P��gAFA�G��yg�z��>�:��O+V���1�OF��)�{��ԙ�}�����ᴁ���t~�|9��B����;֩S_��!���3�Ò^1G���0��F+U�ߟ�$�nR,�#a��c�R�QR.������f�����|���[���a�,�a�'0�pP9#��q��B� W�RWQ����ķީ�g���7B��{�/	gt��5��a����uؠ���^��p&���I`k'�[�1$zn�m����w&�`�+IqȊk�\�Rxmm _�.u	w�����^-|"���:�$J�,��������Z������鹳� w��g�h��|3��r8���y'A�ۻ��-@_�J�^�o�
�8!�vS��xw�/��`��*K9¢q��=  4����B�{�f����]dI)mʧ_���pi�|�QS�NM�@2��$���Ep����G����9a:4��J��w�,��܉�Y
Wx7\ٴ�)	څ]Qh�E�NII�/�x=�DB�Ӧ�l%����-�O�y�9Ԋ9�[�zq֓<�l�=p���k.~�Ͻ�< �x�s J.O>β�����&0�}iru[F�ŴŘ������D�0ǂFr��O�$;��?o��p7�.����吉�����Tf�nDZ�ҹ�3� �n�RDo��&dy�/�������U�9�A)�a���j�h�9�<�X���7̲�\9L�����p��iv��J'���Pfƶ�	��gf�j�,BL��+P��517�=T� �z�6�И�)��k�P�Ⴖ����yX�gɍi�4�����|A���Vb呟 ��z�e,��7L�n���r���	���qL�-��ĂFl�*��Ŭ��BV�	q�A�[���3���K�d��.N�H*��@ٱ�ț��OM����P���Me:Kj�.��,7{D=�!�z4\ >��T��d@�^��m�=�|s6)��I�\'�Ŭ����}�HRf2��1�4;��MvW;n�r�y$����\R�<O�D�߮��,>@e�9<��$5��L��L�5P�#tW �TXe`;�+pF�J��je�-���캟�ϵ3_��5ζ�']#�d��t1����i�5�$8���s�lb=��\�*vݶFH�h��#�Esp]���U��qR��.E��B��=�H^��S��L��b��@P&W#���H��R�H��G�a+��Uu
g��@�_����	y����Wە�9������'@���UQ���q��q7�"���y��NZ��Cݬ;�� XE��"=KL�5� b(��v�tߺP��݊��͊���0�p�hkWi��e��(ΛD\H��@��'�w�������.H ��0�[륈�����t�֓���fм��vK�� H �+��Q�`���h�����| �
 H%���TM�ԗ�+|z  e����q5<�O��_a7�V��Ѵ�b�c𚫜&��^�-�^t��;��KB�ǋ:�*��\���n�띁�[��9�kF��H��˖[�����Sc��8�^���E�0$�67{���ۿCW��cRD�}\��q�~ �Ocv����m��r��	�͊E�+y�����Q=g�¸1C��78��A���CJ˱��W������ŢW��R
� 9q���\s��S��q��@�r:1mx�K����I5�]�Rd㤱Y����� �\	M�Bɢ.G�v�i��n����bHRm3*H�1x��7�n��D��ܢ�{�6�ʁ.�7^E�GO,6w�K�/���;ҴY?}'��_ ,*뱬Z72�qx�X4��(�*�ϒ����16���Hh�Лi�<��o��(qݚkn�B#ηzX���TA�y���ͥ�>,G��{��m������&�	ׂ��Sښ�M�`�+rO�cR�8�m��,��D�5��u��D0�D޷O������X릭��^Q�"|�4R|_�6�^�`K�B3��$�ͷԕ��/��I�����3�(o��*�4�+�t�	�k���o��1����W�ś�ܷO��Q:L�C��,���}ܟ�j�A+�6�>d#�hI���S�z�e�ren�3���L��n��������%���ߑ�=��������e1po�u��G*��8fs��갸̏�G��-Kى,���#����K��wt�^Ė�b%Θo/{��5����>��h\�q�+��Q��Hг���*[��ǁa�Gy4��YZ�:��tH�@���5�G�\a�\3riu 3�	/9&��Ϗ��`��]��l<����3�#?�^�J��V���J�ͽ`*~߱�l�K1�<��h�끼���?������.r�r�#�F���M"�Ԏ�<����ˎ�=�?�>/��X�Y?�R���e����<��A���(��~λퟗ��AH%i�`�����+��Y�)�li��É��9g�"d&���\���]:y
���&�c��8x��]���E����9���M�tn{�W�YH�!vL���r4uy���qB�p]o���c8$�9S�.p��(�$)3+M*������l��C���M�\��v��Tns
1e ����p'S����^e\��W��N���6�־�}�c��Ԏ��8�O�+���pF!/���r�1Z�K:��v��b������.�����*.wK�LĜ5���� :}���8F02Ŏ��#,��~|"Dq0ӯ�ȴ\f�!�M ��q��h�V/ĳ`�ξ�I|��v�}Eڳ
3u�_h?kW�5��oL����
�ܻ#pP�Vtv_��ne���
~T\/o�ž>�^�Iw\W��d���흄�` ��s/�ĳ��g��CP�d��OZ@��\i�������%7�3����~d��$=�i��&���	��1��P�/7��.�Sh�h��b�=R�t�C;�GaJ�$_.=o�sI��[Rm��79-��V��{��$���?��ո;�Gw�q���N�%\Y�ힲ��R��ߢ������3I���^!��&�8���ׯ�ؒk�-��h�J�ɲ�&n&E�RH�z�GgL���e&�4�S���$��sGmo�21s���Ep�
RR�W(3��&J�� ��dV��@�c����~�x��
(�n�o��G
 �G�3I�ryg��7e��&	]OZ�o��% c޸7 �Ϸ��D-���X�ۼ����S/66�Aw�����c0c��d!����G�V �7�F9���]��)�v:�&)!�zv��̑�ܴg���.ɔ.[�r���(��!M��E<�X���>�V��9M��tH���5��t[��=��
.�2/u��V��`�{���|�7��T���g9���_u�4�� M��c�
��{Xb�J���)�G˵���e[XE��6��[:���k�����y�ҳI�az�\�\ol�K7�g@�j;�s��ρ��**~�W�h���*�����b����"Uz�F� �Z��>";��E��@k
�.��ˊ�Vr ��BD��M%����j.&�t��d���~�����A���:gI�y�!��!Գ�%]���c��IE�痸��9ǽ�?��*�J�Ob~g^��
�f̹�'��i�W�2�kfA��=�b�&k�R��v�N�sl�cx)jT1rRVŢ�['�R��F�W(,I_r�M�r��p�oqG�(>��j���4Q(�Y���wh1�$q�^L���-N��{�r�� �w+��1:`�~ �9������ӱ��yRI��5�մ_H�e O�`�&�2�RX�?���=@�~=6��N+!<w���C��O�A|��x@�ބ�z
G�����[4>0�,F'��q��|J����@\i�p���G��ާuz�-dՇF�M�+� bg��@����k4_���Ca�*W�9���#� l�G�p
�{y&��-e��YО�ر��DFٮ+������>8|�=?���T55�s�{�A������͍�p�(�b�Q�l���s{�:Yl����y>�f)5�-���
[�4`'�L��xE�u��#�DK�~&e+o�>�
hyN��#���՜QY�$�V{�^Q��P��V��syzӽ�)�|�VC�q������;��D	�ܧ:ͪP��CC�%�~�PF�B�� �D�Y�����v�Gяu�����k�������g��d�d��2ϜAY��-8�h�={�C�a�Ӷ~v�c��8(��yQv����n�*�V�fs�k�������z+,��#�����*��^�Ŕۖ.�4�xIxe1���5܉�_���:�o�]n-)cL�{��8��u�L�H�N ��/^ԍ���xY�F�����7Iz$��ᆡ$�2���W��r��l[n�l�9�� )���M��?f÷4<��~������*э��!m-�RŀfB0���d���>x�q/�V.���Տz���@ک�K����a�}y�<�>�g�H*�FD+2[BW�_�8iVcw����r��Ϭ7��/ڶ�F`�WIC֬���>���66v١{��~�+�.�ZY��}�c���x�zW��!�>R9�>\De

伇ѭ9���Fotd��B�i%u�~:h$!�@�۝'�l�O����fm�;�ؔ�eou��<$���d-�G�Vmu�A���Un$n�#�d�{��q�~�L�Iw�������*ZG��M6�X��\�7��o�0�m"ヂ�]c<h��+M�f�����!���+�HT��26����c�<e)������S� �
%V�m��V����:���Yo�p/5g-^��v�ӈ���^��UE;�Ox�~��-~�Z*����ޠn�-�飝�")RJM�1���W��ؿ�A�z�bi���#9���&���v/�~���p�FM����F���4�JM`s�U	�{W�}�Ť�L�]�@KwN埌ձ����\����Iv����|��~=����������R$�
�$o~�9�ԇ*���F0��!�����(��u$z?�	{�jN�߸�B
t�Z�ϵ��d+�y���Ƽ�6bƈ�z&ϑi�h�cڞ
���{|������r��=�O=�9eׄ�8�ə�O�L͹���S�HP�,5�\.ݿ�4�狅C<G�8��I����Wn)#@��A_�����@�?"�2�5K{bmi�� ����`	��S��������x��z?t�AZ��v��)��m��ƾ&v�"OD���΍m��t�u�^w�/m�7�*p䖩��_�1
Y���h�����&�噗,I�p��>8`w���n2�OV <0��Hg#�1� �|R3��Uւ�Y��Y�?� �^�Q����/�W[��2�L8����p����	��}�P���f�� ��
�yn-�<�ARcn��9PY�!�ƄtQ����D�UJ�D��-�|:UL�M�EN]�۰l�yЁ�3C�}(���,N��Y_��<�� V��jԑUd5rqK�g�7�x�c&���j��-14aױ��9��7��a�i�X��CH�N�W|� k��@���|�R���7�5�[g��a鹓�e��M�>����z?^��04W�t��Rv�2�T�:F�@�mZ:�g"��)ד*�xM���>�7��̑�����s��7-H���$Ÿ��գS��9ZD�Y�l��Я>���T�ZS3áu%�# ��8��� o�RP���� D���>O����ڕ�]m��pg�����jg����z~x.X-p��T��O;�Jy�U���g��N<G=7<�eu@��e�܂=��r��6���?:��dho�C�J��r���ar���$��ckJ �Ī�)�Br��	��^[(�d���Ђ��ҙ�b��c����2��ad��F2̴W����?eϓA��@*)-*^�%�]�Y �v����.��&-�Rwl�MK�rTs����A�M�pe��ޭo��r�;3t�� -��p��b(�$����S����NCk��(U :�M�7ޮA�qV��� /~�ǝkԲl���F�9ߊU[�v!��47L�*k������$�7�F^s�a�z;��^eU*pa�O6�"��~����j̨J�-XV���	�7�|T�T�n�2ޠw�&ĐC�s��,{�?�����Q�$��h���Z�xk�o�!���`(c}3��!���+-�~R�9z�6�c��i�,9�ϘZ�a�W�� z�$���3�����@�L�vLΉ�:j�J�_� ��D�`���l���j.5w��h�W
���%O���x/��l=~��8�X�³q�i��	��<��<Ȳ�rV}ڒ =8�y��~�f?G��Ig�n�L�
b��i��%�������V ,��w8�cSl�u���`~~\kZ�0�	�$d?��`1���o"��7�X�%b��.�`��S3���p.CT�:��/A��Oσ�#��s�9��,��I�2��I��	}��}���!�/ܥi�������/su�-�d����&�b#����E�{ۏ_xV���)8�'�1n7��~П�Q���]�-�J�l�k9>_�JI.A~���x��3�>6�̭���[ʟ*i���|a�Q֮�֮K�C��%�Өwa��UM�wđ�z!C.����)5���Ꟙ+k���}_YwA�47�1��1�:J�i瘚����\j7"��2�Z���AKm$��ի�G��E��K��y�<ހ�+�?�7A,�KO!bCί�#��`_�Q���TAV���Z�O�v�����#1�9�*~a�w�g�k��GD#g�,j{2��\]��ؚG3��V4[��A����_-�CqVQ�IҜqŸ{�������K��O' �Ќ=�{,	�h�)u���UJ�н=ya� ���t$A���̭��^Z�j����#^&'�N;D�u�	��`d|��ᖵ���2T����8>�:�1�B�<��Y��ۗ/�]�
�&K[.��9q�T!�edm�����P���Q�@��V�^(�M�Kn<Pd�R�Y.�O��vW��K�!�#��7�%�T��-�6�o��lf�B] ��xx$������=L,|�n�Qd�R�D�[�N��V� �uOc��H��' ܕ�[�n\��Z����"�s�{����\6�Ch�������S�)uD_0׮	��\QjFKz<0���2a���_����"�dj|���>y��glP�{N;�x�t��z��R��� 4޴�9w�"��|�Q��T
�X�H80�mW�ʶ��NW���dv��O�qA#�D<�y������L�`}*uzl�]�WD���A������5B����7���)���p���Bլ3�L[5����j)�6g �_X��ppՙ̿���&1��M݅�vSGi�O8�1�_��E]:����U�EV/B7�ief�(?	��:�ʷȀ��蚺���͂��,�O��q����8�*:�gY��(c�h�,'qB�#CZ�e�Ơ7 Y��?������Y4����D�㞋���/��F��V��mǭ-V5ybt���	!R�At�b����|������%`g�s�vΔyU:�_��ke�O�EQP6��.�����ӡo�5�j�l�,c��y�Lk��v����C�4��l�G���t�NS_���[���mVm�.N$�_C/�����n`�P�W�+�Z��Z�LpK���C�kQ��[�1@�h��u�{V͒=��|/>?9J�ݚF�?|�������J^����.s�64�;������܏ob��O�n�Ho�.�~r��� *a�&�Y�7��+�Da=A8������� 4ݏ��ѧNp,�iqF�8˦�n �L���s��8�Bu�`��[�N���"��
�#�=�5����͏��Wx�l�.�OX�UL`�,m\��j��IC��G157��?h�C]	���B�Z�(�ݶl������f��ԉ����n5��<�`j1ُ���qϨ���	��oɱ!��~qF����>�3V!�̴��жB�)��C4��ƺ�[��$o���w��� �� �\�9�H�o4Ns�\Imי͎�x��_R?6��PΦ�vJq��4V*��U1=`�-����|�ۑ����{���7"Q,T��I���2��_���k��O��}�����ݛJ��6�IE)?[r�%���KÈ��� ���D�E��=�岡��[�?l�e�sL�Q��a�W��j?C�&wB�x���AJ��R��� ?�V0꿂���SI}���*�����.x���M��s��0a�����n���VD�{�B�������EJ j,�|D���U7��K�H�1p��*ol�}��I�w���<	����1ڱ�MN��+�R,SϱYv�	�p�?k�[ͷ��[i���?����u�^�N��J�Zx�k ���VAH��jCV�4LW�HV4�C�BC�n�F)�K{����1(��Fn��F;E�g����ʭ~�9�$
 ��.��ч���sK�x�o�߬4�9�F|.|/�� �I������zͪ�70�����wdJ+�k^����.)Y��?Y�(V�?C��&�E���=�B��-(z�eqE�>⮠�&]EV=[��#��	I�ՠ��d+��j���_{`0�Ү��+�q�Vv���k_iz�暏=yS�R>F�e"�(W�
��<�|p.�m.�I�x/�/4�N�ib��K����t[I�;��9 r� ��G��:�Y��:/%��F�p-�f �*={��݄;؇�dt`=Gn_
��&o���fl�q���do��Q?@�e�7ڠlC��n?�D��=x=\��.
�5K���D���w�7��
���>�J�L�j,�b���� &呕�Sx��F�G�����a��MMwD