------------------------------------------------------------------------
----
---- This file has been generated the 2020/03/16 - 11:19:27.
---- This file can be used with modelsim tools.
---- This file is not synthesizable and does not target any FPGAs.
---- DRM HDK VERSION 4.1.0.0.
---- DRM VERSION 4.1.0.
----
------------------------------------------------------------------------

`protect begin_protected
`protect version=1
`protect encrypt_agent="Synplify encryptP1735.pl"
`protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`protect encoding=(enctype="base64", line_length=76, bytes=128)
`protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`protect key_block
YtCLBBxYQ5noeN31YMjslYg5ZteQCAUN2M3dpR+Ebv4R5wJT/AcMgb5y6ZUKwSRP6XMzCRuPb1tX
I7zPMvpDpT1RFl0dCQAtrYb2lbTmJ0FfPUlbUX3wDVFvd84tLnhPR4odPDZ9m/bYW8aBjHew7/op
iiaS3Kls+SdfDa16jTA=

`protect encoding=(enctype="base64", line_length=76, bytes=864720)
`protect data_method="aes128-cbc"
`protect data_block
I7ZzUt0J1qVIr2pudVAfqX4lkRqDZ06KHaodbY8zR07SOmO0NzP5GsiEMlny9S6ppRoFrlGpiWkz
NLVh2cjqxNaPITx0CRjRNHPMYkPigWdSGbrJXw5hoo4IRUcY9gZo8OIlS0GkwLdVpok+P9F6Xs3B
Upwb8sFg6RkHHuQ80e8Mlh5ntIdrSlcnObHYME9mgr1/F1K9OzOAdN50AkuHnE/hj1OP/jkbKUzm
yF4gMczYLABDsepCUiloVUNY6zG/F++0brT07ZhB9OkKCeehuGVMw8xkQnS3ZANqoPe1cjoqReIJ
doS4ICSIFsJhhdhPL5tSRYAmA2bvUG2P7QsD9NY7Ah621LVxw1KthHGZEAHwBwfSgEHiVfcMSG/p
2Vdb/9AY0Khwjk5e+zAcr2360G5VvHkUSvQmcklpAFUk5b6vKXCNH03QDtBTEMCEYQaaAhLRiShl
Det9mXzfHUv2WNs5QSpEunlDkFOj3V5kIS8y4hx5T+Tfj4ascA/eCG0T3dMG52VI6ILlZu2o09Fh
VVdDjI76zYZE1rNtHT2ZBe8Yqg7UqUddPbLrbFLz1UdqFgwNTL7w++nnm3fYTpG7cuTYTKUkVGu/
yjj0gdwh8HcubdwoPkFHWTl8D+GwewUqz+SS0ValP+uJLL1LZjdMA/2z09f7avtfQZ/gfp7GLiDh
aFrm33QR1kwtuolGjDUq5jeXaoL/EINIhtIRlHAwyCkgcvpRoUTObfLhw6s9T0qtCx/VoB1PVduw
cQ7Ey9YiJiyhdqKBtqfCuYdEsrySRRhsDeSMeBPs4AID8p3w3Xoubmmge7Lq430b4pEDn+NMNSb0
wfZhMQxC2ZAX+QgFH6UH3a5TFCqmkIukBmm+75bZPpuL6dhyTsue4Ksj2bwG/O8nVZHBPEvqLEQD
hVN43I+qVEPueMMjS9P6/KiEQVJbrY+QIeFx+CLXWavLCzsCk3fTDDkvZJs0Jq2oDmmA4RviQhpC
H9W5+1shONM7B7NRlq00sqhvPkjHq95IO4GJVyFqndVSV05mgkmPM5VCmCTk/IcfL6/e9Ujt73ji
vIgaMU6asR5BLFdGjtEOJp3Y3soLOX73SqmD92yPEe0MSpiYnQ9M10zwSOcSGhx8jVs9b475YSwr
n8I9HHAQzZG44FGYTA4nKuJjRMoIFYQWWOEsv/lG2O3J+kzNmXAGJmgJaISlqy0T5QHnyPCSFojI
tinOy/X4w4v9akdueseXV5vm6H9l9LDBzChcDGMfcQCGLcwGgEwuOhrgs/DNs96c78vn8PegzOPi
iVdTfIOtvp5Wl+PuZvefuattwGV014tnhg+64he9hPtYXsP7vHbWwWFUqhB1BxBD5UR22gxez+Fl
fHFVnOJKWhVsuacR6I+E/9r8TCjkaPTEUOH0NJX6Qc6xwiIkmo8rIiB7qjhLZfrPEGFIg1RvOW2R
dy4hOhgnk1RtIW4eyzLwrxtUb1V43zR9mR50JAYnNknxIaX1xgg+zZy+t7QpOIpkxSpGXoXG5oyJ
iH7hGqhLF+8/cOfNmIPCCHHpdq7cyBtObxUOD6WtDFozdOpJJ4MhiauRHireh7TXueNKNr8znbgY
xTIM+dxa5TRUDInjgnWbJPfgmEptiMB50RRtszdeVs6wlGKNxx9OfGjIaJxbTl4XXbpx7gJDnPaP
+pgur0k0/jO3zymx7i+Ny06szcu12nkbyIfHTJhBRVUqQD9j77lVq2iFF3clEPUKpaFzcrkgseur
MuwfhibwJ2T89OWfZn2leLgQztFMmZnDCj9dJytE3s1hvyy8roBNNCG3WwIzvrCO56IM/LT4Ay3f
NEwHce9UThWSMdwBs8Uno6nkDuoW/k+g/XGeYVb79PaIvCoRa+jXZTZx6RyKKsnw7FL398XzwjJ6
xUB5hfVrOV7Y0fLm93ZvQTVFsCiz5MhIFKtFFW5J0lCqQUYJtS1dn4m+mVU1xZB5Qc9oEINYekx3
rE5EGTsYnXGdAZlI2RME90r6pIX+P26NFjbv8j0aSNxO/9Vn34z+++lnaLZq3LH7pcVEMpkcsbQU
x/F7G5pLNoA09g+gX8m0DMQ5mFLEYzcvYZ6Lb71EbPtd8/tFOSOeVOCBHDiBHvP1ttEKm5PZHrVU
e8DWcRT7HmE5bMv7wJZ4uGyibQBrW6WYsMVlnP8GTvlEkLBY4RzCH4vpOUTjyr+7DGeFp4hWGnlr
xSczDvJ0tOeZYn4QcUZunUjJcKiW92kUQp/T+zKsFSjzAFGfnr8mMJDy25hoptFwEd93NgKWmEkp
asdnD93lEcnB4GerJlYdmx4mU1TXZZtBSMCblZoAe+0HpUfSbaSVDTS3h/lOERM4o8lFWp7dJDF8
khNtBPXvLkJtaeXFjbIaXDYMLP8fx2fk5VK3yRp04Aymd20sxjXUXZjnYp1wlSe5SnLyvEXZ20g2
ot7+a5A4qDjduYw/O+KWULB6TDxzrQaB4YgcrxTCVChCYW8Hcc3vnPP/y3ZXINUZZ2DtRKUzb/xq
HV6jPUSvXvRpBFAhXHWobRAxVom5aHnxYK+v64IwwLNOmxLcBTHp7CC5uAzJVR+2srRo/omvO0sZ
5MketIkEjHXMLTRuQyuGzPGtqTta3qxDNgjg/Vf7906QAgmwSd8fWKkKYQFU2NqylxsNnxqN6lTt
spfF1nW5cUNgXxlKO+jcn4LwrZ2BgEmPUj/2WCp8TjciwFwtaD9ZrAY7ndUvPEWuVwb7QxbyRrtm
FcuJ85S2F32pf/+UIGLkxEHFwVXByVcsNGf1l9PFy5jgE6BSvbHZIhTxOI2s+fMGOaOVD5zFn1ht
E7lrS05zIhC2FNrPDdU2QOGmlJTIXNEfJjJiUr9ghK8ucuqf2wtvMdg1X+mQ7edCJNQorWNH7siP
74uK7L+Kcr4pR3PoFgQC8mrqQaoLW/VE1BqmMiQaNxL91UseJtazmdzxSQwULjKR5MqXX1y3Bqrm
2NoMBBhBWyMEAxBvZ4Ut+deEl6fcSqrxmF5Fvj3PN2MOWXL7h9WahZM1ggmzfcgbDBWbeWW/q+/G
s2ITtjh4hu81u4tnzL7+FiGuJrwFpYNr3X2kfY2Io1Hb+QZve/YCelcNygvcPjVVHKH5EFWXQljt
jYRmyCid6EfVfziuubJxJK76rETKoiAocJ/Wt6EdbqPV1OTuwl5xCA8uFhWFWrLykMfsmYVFdh9H
A/CmdTtS2FMAcqNlF4dNn6U1kYZazybJydvdHp9D7PqsWUY+opCme2xexue+moDNc5uU4Kh8b6i6
xdranXitBRUZrAPBTRM9PGl1Sp4gqBO0alkJc+eDD26jrnQLN7rCLn2gqTBle8FvohRSouKgpBrV
M99CJf5qZR+BIlCG3S446GPoW0z24V+XIEzrDlof0qfbxXbKYXxMj/WGDyVj+JQHekeKRQSYMTWk
TtmKvrW1Q567IW9FDomT0Jvi7WEXMnlNwLj4AZaXrUKBeL2L067R8xgdhlp81rB+gqhkj+V3Q9VY
yL/grdhfyoa2ZGTOWh8g1XzVOTzm8kO9O2o/zizCkTjNJn6vhhuGUeK79p3Nc9xx5XjaQYndnmtt
BSSu52NmEudy9lHOzFQI1GrDvRals7zL6Ie/CM7/tE0xw3rMji/ATa1nRuOV1iL3uftlf4KgdXLv
vFZl0Je3RZ7b+5qQUm4eEUXfq0XtBWOi2IvGVj7xMJa1F9yslGzzj02QFOvYpFV3ZsuOAyE8CiSb
gfdb7Wb9wRuvdAEQxVltmVraz7x6I++DZqgofztqtkc86S2nIXLBidgqREHMGkSu5l9nCngYCRZX
YX6JtAkzyhJAoRQwHil7BrWWb7OLDT65HD5IAmtJxrhcZ1wMpOPjQbHapBXJFItNsRZkmZLVs/JI
XdZHp8TsAxwVoMtJu73bPmNdRQIDTU0pBrB8Ww2I+4141gyvWKEzqAj92U5EC6DAGzXbh1/Lh0cc
CGFpfeK1wuZNSTLoWslDkDnGFBwDjRFcL7P0ja6gjvSR/hRFQKstb8ZJNpigrM+2WgNvwuYgj1QF
d7Rtik144lvDgVEM6jyAz3KVXBCZ9o9a51CgV+0FR+oNGGth+xDp0drgGCsfGXznasV9XkCv+Udx
w4Y7y4IJGpbAwjV/wVwONkE/74q83W7V3ahHz8LjC0GEKRYsON+rDyNdG+bsWmcgApna94dU7RD6
ya82konShV8rh1XVoJNaabe1M+wqEqavdTrAKvp0FreiJtpvYP6c8hco/FmVpbB/SZCs2L19QS4G
rjrn69cjVWNJemSaGmK2uVwNecm9qWi15M3y1IFzkFiwjARYU5nZ3m98bcodPMCaslfR07buPZL1
W2Ji4/pg+Sj0VOk0mgkdmWliKA7janHTOGOhxxbam6DyVvxuLhuAXFa8XaDONgQuT9np4wCjyox6
46Us++eAUM0SVNEnHxd1C8pVC8KzVv+DbjpBphveSPk+629UcfPwij69rrqB1iiSMUXYlmkNRSKH
3Z1vR9oi+hjBWnBHHssGUoiRkseSHdihUo5YuytjD7uIHMk+baWVbiYt7H06aIA73QxT1YZCOCm6
jhqdD97GFFn3UwJXMqqdA0WAkXj/piBbYzxpOZSIBPcoVMesptaRcKGtb5C4n1pglC05YdM0iAQX
jWAcW3eu63YkHlP6CpVjVIoTGOJ8wA8JjgZbP4xSdxSOvxgEI5ySnoSQMY/fGGbs72+mATZrAcut
v82I4oHnLEimqPwhGzV66WKQXpMFU5JKoThdDC8LM6oc9mTECVK+qh1+HNkDVFamY4eE2pyKt9yZ
vvdZaoP8Nw0F7p3mICDJcibVWgotjCLHaCtkEtWq6ejdVLNP34IU8zACywkVkZsCBer7+2ujEQMS
VktlMO/zNcPH49zJqZmo3BFnQ+jXm4QM/uuf+Qwb4E4t9F8FpL2PxUrHvHgsgECSGfhLFgz72VJT
Oo48IwcKkshBM9UUIbHsZvJiOtgkl3woZgZMq1aYLe+xwmF/h2jB3x6pqBN8HNV7IeiPMwB38SH6
rYX2bK+kf8M03SVOwytAA91USQ4TXRCbmhOf0b/MQaht0B+qGAZYb1mZhx1Ezzlhk6C3wanXm2BO
YHZHJM65p+tLzLiwBjqwdslFT6g4NsmbvnlDBI7H09CDzsrXJ0cHGSu3tX+vZHtQLWklcYxmtU3M
TpB1J27nzt0qiIdSkskhh/iy9V6FfWtIw4SrZcgqp1pjy+V+634ibuYbvzclKjMq9ffITn9I8L30
TZLT5SgR3/zSc8cd/5u0hFsMIdS3QxAKSDqu3Jua1YfhPpkxp89OOrIP3c5AmpMQ4DVNeHfXpKTP
YT7dEJThPj8zBj3rbhK7McWzsf2+YtcYjqYJklY0awhgOsmiyakWeMaKPJTZFA/2xCPdPGHA7+GM
7aoNmZu8sdorhkBt47sZTQVOBKFDs7EOVmLtkTjlOsopjTKLHMNmCm9GTjegpiPazjX6NnO4eCbE
c+GLP37V74Y6+SUt9tCqu6+n364RXpLr1s2dtYR/h9yxk9gvNckzE5ZEThosXuVYMEuBL9IaaHR4
y+P423gXamACgF16LDd5RYN/zteU02FC0x73XBWdJJ+9xGt5Fn0mPPS76WYtelwfxRJFKJ/rkFru
ogbbZwpXPW7eLSb9SQ5nnj8C1RNKd6nBYZU2bMqKCrobLB7QBqpn9SQjK/lKQUhtz3QtBYoO4FYO
yqQBgeqErHY1xBlkXKe2zmC+vhG0UeJ006nb4HPI+f03D3tzjgVUNVQ7CeMXrVtI4jUpwnEoK+N/
BBKDyulUi2U8bGofHlb6F3ASTBIpU8saD9xYSdLkHmd+velbs2ZgD4Jvt4TmDKt9TCvXIhRCji92
XQaYCFPRDuJKbfR8MB3/A/4A7zo7rI2dOIm6jP0JaLClXRButCjb+DTo5o2qrdu/cjcrVsNqXS03
nuOnS7ye+JGKK9T1mNhIMy7p2yzWHcLJKNAaZ3D784wazTmcCu8Jz3RgkGIRqSPdnQfrovVBZoXg
U3naRzOsf/lITVPtKSHR0XQHyWp5XWqOBlky1A/gGMSsC0Xp2amVBw7IKjmpLS89OJ4HXEPBUR04
Ppsf/J0EpPhIwf2Ek4yUQqCc94dEzy8hfBHVbdv+mqEEjrX4tJPyb7Rp5WgLkFtEG2G7k7I7Rh/q
7DOhhJczTDLahM/IK315k+SgrzNget00BA4f3Uyw0Jv3jsgbdJaq9rrISPjReDOZEJIDS+iQNeeh
FKmKmv67ZwitYeCeNZ3Bo1p0Pq1KwHwTx5gz+LkDn0VhMTsLkU5IAxxJ+pB8pCA+H+T7oGuQJcKw
MsY5pWTvenqCproR3p6tPWXzCcOfsL4xWaHlfQQ00jg78b9O8eOZNPEzHiNu68z+BOSHghBkKxf5
OBWnWGjDpSieq8aMD+DnrEFkHXzi0yOAaL7OaDGCWfQVaxktxFXApZC6bdgdaN6mqiWBlMLIbKG3
BzHPILTSfMtTKAoPe8nmWmMiQUr/AxSCdUPsUE5bkjs1tuENasXg1RuQVf42W2sZA+Zi7SKEOXLU
vjUacKEIaLXLGiz3nphfS7qHDdnKv5MwZdlH61NdDS3tfm/YjAzoipXHeLO2/CRZ5MJn6cLd9Le5
6yrQi33Fd2oK1Y4aLLWSVwAjbCtbFzvaksrMUtlVpQ5EYeolJ5oqLVMlM1uHBE5GYHkOjyY+6CEA
frrl+HOW+N4r66qNYLLsEKjYe8rMdXNe6bHN22ucswopeV2HMxts/6iO64Mhq7583qXOjNefc1gA
RakpS4aNRktzo/w6HaD4K4nSQevAnpOnJaGtgJIPAB/mkEG6tEdZy8ldCDe9eL3LhiAzFiJCms8k
yn7Y8fYznC4XjB20laAQTCNgw525e8k1ZWQJFm1hBwobBqdaaoIFp/ZdMft4mKAVP9DdnENJo3Wr
9SsXmqQylxbbeblpeet91WsXnPEbZzp2QEokdQUSivG8rVU81/8SOK6v6AfaQmVWJkmV5L8vGwBr
PUbO2pPQsmJMaEb2dcT5ABjdZWC27FrqKud0tvhTsC8QqItxWtx6jYBWQwiFcx0rZ3k/SHNKnFyQ
REvnfHdwWPPWzOq9m4O84Y8o961+glrMWdtCA4+pHDuy/pDxcHjrYWHa68EkIwtlb5JfOc4SR42T
U98+IS35uX+9UNByqXP6oQa/uvi7d5vCVKdOXn/ZoO8LKgXZbB/8bKh/C+c+E5975hReHkklLVOA
yChCDkyovBnl3MqdQEGLcVhcVDxtodjX7n4jv4bMNGN9QFw65YMKsFe6My9j3ZkF3BlkYzMf259M
ZMd/mP0t+B3L6xduyelU3yelPbBjEzKCxZUMT2mSdF7qUeLt9DSjPgjQVWWS7lLg7EgYaJZYMjGm
A2sbPAO7GIoD6FueyBHQsi5eoTo6wHxk3A/MblMHYcrh5oOUPDgUAf1zeLa9IIsLafZjRLyCrozE
BSyEfb5L3WorK1irllETqgiOlZoMX102PTcglPHyvCh0E4pamiNEpRZbAIJoTp375NA8oDnFmi3+
b+6ABvuXxkFqC9J3IiHjkiTdZKa8sYqe/qLLjjfhcKujz/wDW6Ia8NbtX8Xnx6w4UeIFjw/tuddX
BcYzKnf8vdkVdnIVNVE+hs/M6+U/bllr2KRWBZbRPZVfAajozaF4xZpuVD0XxNs+bp45/9Cn/p/f
q8crseNrLGxKFbuIqBmtHHsNTQc8VtajieiV7i0GCvA+wwRYV0kv8lfXu/dLDdJnOT083jHI/EiX
JV5gPDBhmU8ez6l6nXI5LeWH97zKaOX4ewJAVhhHR67Ma/EJmwxU7Uvi92g/4o6k5s1+amlZkt04
fR3ak6znKbwo8OP60Zk3lgLG8U9lQHGNitu2miamwKfQ5ZK/viYwSMtankgdtGOgltPukfHPJ9EB
Y00zoflYT8stiZgWVwWKBTy53p86JzAi+uN0eCw1OgzvY3+umOIBSKP00IGRvocXjTys3Edfq2YN
5eckk2G35rL/m/l77qRkbrrIvDUWQORPVjGfnd9seu/Iij/PwOYc3QdEHX4NK5tTKi94feMfn8eN
D6iTy7TsCUzbN1YSCHP2PHr4/GMlZcV0To8djjsvS4aBveIz37EAWzvIuJqzxTMEZBC5izFYLBp5
p+FvRjaIHVAyNmg58yb1TimjB2fkh8tJqcNkFp/cesQIu5h4cOtJpZ3KjKDwr+GnHICpJHUtFjpr
M+3+swoKsjrj4t/IpfHLNmL9XE/Khu29Coh+db94oT9DplpMzw1itg/XIbTJvxQiHEM+fOsiXKmM
tCHiOnuAhvja6C2WhB6ke2MVWMZrMnVCKUuulP8Qy/tKOr034E0H0tNJccwQJxRjASPCt1kkePBy
crphM2UHwn79pyhfSRKe+rVOxjRI+FY01eob3Qc9n7EnEi2yNaDC2H6zWC/vpAKue9r53tE1/GGi
p1pkYM9oYM2jmxEC6qdKUgsiR2E78ae5EdhDkuwUeHnnZfSCRIsMx1Ne/LuqFGVpNJhcBkx9R3rp
8r9+9mok3IqjCsA3MsfE/FjuYLAirjWtJgABCo3YYJYk6lctmV0eUT3Vm10C4nRzZEMSU/mhR+iV
nXIM2+CWhdK/4fF6f/lSNxA546eVAaSV4xLH+7eww3/jgKUH1cLr/em3yGdRVDfx9wJ1tHnWG1GJ
ZSx0rWAblTw8m1OYE/6SbVeJInm/fCzGAxSBTPh9NePj0SVY0QSi6wDpg7H7njGsrWMoLmAJPxkP
3gFQO+6r/3ZzB8q6o+fum9c0vQVBA5m4M2u/4V6XJV1RoeHpWhTknPXRSx3x0sj+zkNuabZiZIFw
PAsgz5Yels8Vq4T6Nc7xSjuSTWzgxROSuZapey/rXK/ldaQGB2nOBYKeTkY+cYN/bXbk0Sy600Od
eMCnnjGQ5Dof2yl4iPD5tenkd7XGe+tKahjhQq97r3QqUGHBgd30WGUT+zE2pSDxNxLISGS1ngz3
qLRU2XINy3pgm3NULr7WV1W2uBrSD8Im7ao7rHNimsN0BIugdRm8BavW0lGNiuJbM1thYCzfjtCH
9dH6RFNG5zfXi1wy4yO6AMOMgiidulOvEuQ76TkXh2beG4ow5XM/EK2pry8ctzz6/2t6BE2sxU3g
mzeaTtZhU8jwa6kzZkhFEVpzp4setdGiO004wMiqlDA4gD/RN21Ij9DvOHt3nZS7qOgbyHnMukbA
hOXxjl9oKQsGomC9vKaV8wAu1kKY9YLp7xXqauKktMhjZhqZP5fnGVJAHCoinX+y1XgRblUn8Dy3
rfG4U+bQ9oyYiNL1TE7E5jfmm4QiVnMHzWzYxMJPdpJiN++v3Y+RnZdMP/k9vHsfaTOGjEpitIfB
WIW447qOLUK7rcwrXU67pX522Oj+dySY+bkK1uSGqDQGCe5aEFSZPXtoAL65l1mwYhWVUXo88JCQ
GfAwx4pjjunL8f+8iGUmhEnIrv0XNAUrFcOgfHHBlU/719jDFQjgD8v6/ArhCYsbWcd1wobia9jt
gpDCk4Nar9U0N2ZSfdxHFMZnPZQKTH+KVBpy4e8dDYmCClW2F57oExKv7N0I0pROYf07fmagfXUh
OODXBhh5tiw9i0OCCCZH70CTd5MfMGSe+X6++GzLvB4XIe/SGL1H1BgHgADahYWAumexB66gvg0r
7otW26L1JcmwozRZH1nhv3EAulk5giWHjpjT/pgdDL2eGRsztqv0c7FHedVXGh53OaeLlrDvYbNt
ZeWy3rxGdCxbiLpeFkNf6Cj4YYkLWKeJGv2myE8dUgsYvhV8185tjulWRfeVhbZyWnKxwrasAfN3
dRLpYq4zwM8Oiw/NFQ9Eka//8RJTlCo3pyD+YXnQ8gPRWu4G0T4C4tF0oXNl92mAomWKuRP+fqDy
Fd/XY2z0MzELlzcBXpMGjvycT66pvjiJxVbo5I/vOgSnWVPXrR2jEbJoU0ipgOxVUn1CnxwttJk4
Av05tOU/vYds/Wr3VOVk/a8v4Gnd7XTMYBIWjfzAIRcCGnfxyccz/G4hq1t3CPG5qSI3zWz/t19z
A4eGawHi3uSpKAxUBXVWkUJV2cO8BJXA6wUs8i/3XCXmFfCuX89C2tWpktqN+3t9V3Zfy2+zgt93
qP3Q4/NSaJqe1pwcaYIA6U4DIHHSaDUUkjOe9ySmoTleF5l8NibBBs8WzCAjyrwhv0BW71BI8010
/Gn3b6OUJbPrswaYppe4DK+UuaejRujQEbBTFnoh4GMalfPzlYuBDkukDk1RjbNOjLfqOVWRoVU6
f5IG8l4CuHaqlsY/oNHw0lkbeCWTojp+EaZWMhjkM6Ez6FikR4+S6mPgcduwK2os2tET3UXreoOV
0hYhExdlPX4s65SLDiUwZAAnzbk0wFar4+60SbJJWeacyAe551keSOCDEO/Mfz8M2nGqr2oxN2Mq
ENFUE/H9PhvVmyxK7/wJEKgf/aUIH4sDFtCd/KqqqwIGQDTCwULKQq20SStgUc1LSm5H9ixRNYDi
8cSCb+3/p5GyJ1zoXhcBa6trueSMZoCxBLTh3ZUaOfVE30iiQRS8Yg+1oejXi/0wcNOPihoKV1X2
p+2vC0GoajYeveuHRLQLfZOGoaYGMY2BZqgluE/G5SXV6v23XG3a4hal8By2/FeyQR6LmCMeNOKJ
uJtL42Rn/0PCvyRq5uD5hmaOtr0Xl8qzgW/XHE0cnkvRHdp3vJaOEXGFtHfvrwCzkuWTitMwKCur
L1gkLH0UyIQxxWveZdQwhYeFTrdZz/DR+YFmoNzaLVYW0N5ApzrDVY/+YVXZxmzAiEhh9gKzdZoU
YAqgumz8CsFX0uG1v+LeVDyHxhyTmwSx/gx/ieTVQqAzgbTna13l35dLntnpko/zpsq36BCyJ0HD
+bevebZ9OhgNoK2AJd9/LRr2Bd3tE7xk/7yvnv4V5ZQWRXHzjQEb15v8smY02U3azB3EHExaDiGV
c+8TkAGEC0KPcrqBHEnRcHQ81hv4GZVzroxDWeAkOW9a72lclOTgVt6DSN+mB5jUgt4qJf7UR3ta
k1X2bpB0RfW71ZXU2pkvCZJK00IBKDkKcfXaiPaA5s1bRCMr6PH9g3jXfovytoYPWWR0LDJtqoVp
Dl7CdPAgXcY9UOoZ++MoQ3YtXe/ixVvpBlonpHcwIHXi71ncmj6+oiZSsvhf9gi44rxJCPWWI1XE
rs/A8t3UW7OegIXru5wH2i5G2VEPl/mZ7dsAVzIK6k2gwdDRTcBWeA9oE+pFR/ZIbz9zc6rbEcVr
1LNBsH/t0fRJMvim2tdhHws3CH+5q6o6cvvATLQVW5dwiV08V3c302ZpB+scVv3JflKwA7UivK8r
CApBLexkMDMbdzmxxMMwTKtI37nx4wyd9RDeDtomhYlUv5Jafnz5/phJTDkNh0185qZiGTsHG2AC
WEGwPZjkPOQVZoGZQD6wjmdGN6fpvrLwgJPs5aXcC5u42riCxEBHcUUOLBZfE+X0iVElRrSzeLO8
xzi0qyCDDhL30SpuMP9OIDEwqL7pZ4Lku/gAJ4hHUx256Hv3+e+aHapw8LVtJNVR9CE45viUf/18
1Zlu3VDTHGgxULXqZCbVQUIOxYjfE8/m9noCPZELZ6JN+eJ90PdBOQYwTUkZM63IKzy/E5iV6Cu0
IBkuT989nCrd1LfZ3cb94CruD3xIur2ng1Qdt5AlWy0PkKl1y+0nANUFDr1hhEypetK0yDaK7qUP
CXzWsm/hJDXFsEq60Ki6HppzsHhkbvCocr2GCQukJ/LPBMS6aXgjqyXp1qElEcdwMU8+b6yYDIBH
dzsj7xiY0AzZl4QvXjwryLJu5SFzJL72PtaB/CfD1GH738vv6KxB4lqkSz8OcGDM5T/8UL7exbBB
EadWiSWkjzEnnNVpUVM6Jfhi08JHPETj+AjF/6cc9N7/ylFDPxy0US/QmSHo9CrE5cYINUBnnTUP
RPXNB5r+hKr+zcwWpojM2TdN5hDeLmBWjr/cTCDmrq7XyB+qzoNnAIcrWX+0TCIdedMbcBfEo/6m
lhlMrBNp5dphTeNx6eEfjitcMVFVtjgt5GV5jMmdzKq7z8DKBa7ys9zdj3LoZEwkQGCAFVjRsLO/
tkCzSCeUmEKH6hhv8MD5sJMOyrnJhACjh7rC6jbTfrGVr3eGJfyZrAkx+7dyrjp+sSUjezA+LgG2
wZGk++prWO0Fdw2BRlSZ9QI921I2r4HoY+RJv2Je3ixalRQ2fXdQR1wDmhQyM1eN6SI3OhFcGS6J
CxirAd5tR/tdzNVX/CmSwaUYZkgFfHZIWMAYi6uc8tJZQJ0m/m2c1ENkoZgfO6yf/p2/xadlBxTi
2e2qi0XsyQJWT2Ir/3sgjUmz3YW6GNuoNodGKddAA0MzMhnMf7YkHrWwQFxYNpr1yfCvesRttXwJ
cLp7iOjQP2Q7Zx2hfwZsHrXtdX3ezzL2bqXGwqNcfy1+wCWrzKwhVM7m/4ljxV4gJq5aAAw2Bhua
+Fc/alPQCnxpzlgMz9nZbXSX4NrJm+9v2eouFF5uSevny8+XaVHin8z0CyPbIYVb0wZ8Ita+l4lj
19OMXnNAfz5bQrEKGMahWpctK9wPw6PgiC2MW/gbrdlI57YiEu1vrDtAn2h49n6PAIAWj1kL9XfE
HDg1z9RGYX20maLk6t4dZbh6c4ta0esGT7/2JzAAw5oyRrPAQ9kl5KXGngBNc+6QRKrbei2sSDTJ
AdJ4zgoBznORu7QOqYxpSyjvVSMTHMXz7Hvh5UX+ZRpnlKMlPktO1nEJLtp3e5iYvj1MJK376RrF
rEpPzbeoBeyK74x94zSFS3d+Ea0ARX3PVYmt45PPIljSNHb+TVwKy2EFcrB5zUqvQoTitkKbb8X3
YukEbmxhnKeDk8KOzFlKJH4RsY6Z3/QM41ESWhqHombMdW/3CI+cL6l3KJLZJPvCCjL7ha1h3/MY
Vw2vGWKm354AMT6GSE/hrxvx9XIZN+tP5rNZ3UCkpCBin4VW097O9Nw1ZCF0MH3dz6YeeYuVE/R7
rMQD8Yt/GAOadN6k+ZggWeq2DFcUWdn1LNNSNUqILULw05L/txtSyPXjDwnxo3Pshw2Sg+bk5aXX
H6WcOfrHEdGxKIGa/MqOyg/n1cmoYGjWsHvfMGKkPxDNOQVItlQCfuhisgovSzYU0AMhzKA11g6o
JPsr9V76m6FhFJ1mt+/Re7IexqgIGPzgffkX6QWeI1aQk09eV6w1BejNAgcDpysB0OmEnmk46mUV
wkDeT0W9hRbQecpW5BGC16GPdj5tqSTPoMEkwoiL9TRH03pKv9dB40QiszURCj/SQrzb1rNErFrn
1UL80iNjVAIXnzehPdWZ0tWUtgJowUxFntcR+sXWFe1PF52ifh4FOh+1EmlEmibtqT1Z578j7V2f
z8gUTw21bSXcfEbk9DDlD9D8P2/uO/jr5FRHNWvMbY/kDBKc2MDPdXiDCV4JhybAok4XTxiGtr5q
XUWATqsiKdSC3T4m0PhhrFeUz2eCbLRxUxgz3G/VQMTuOYdP38L/qESdmP3q0i2h3q31+lA1Uxjw
kCmAvQRoMFgHDm+JoKs9AAIczbtj9Op0cfS9scxRbnphQAYo93wmN8vo7sFykwUpw/c32T8tArsb
jWMNoSGpX7dzWm4avuiJGFV/9zq870I/mXbLQRIHSeN2rcnjpdfcg2RuYRSPWAA9XVCTSgsqNAiW
0z+r6G8N+1qU5YzgyLpSA2aSEmY7KaOG9J5W1CxE+xcKsSJU5+t876cnO87F9v1atTOkMy3/MYKj
e00yFk96Gw0XZ0Ex9lRQ72weOVM0CWyTj12Rr35MO03M6ld+q4XiVh/GEifHWB//QIkR03P8tcIQ
ptXRZN/9RoQ9CFCqQBxmcuPJaMe/My8y2bsWnFJVJcJQTxC2HMNA5rZtET6jj65U/du5UxwT9HAT
A2/J//zHbCgbKYX+neldYBuuQ6lcTrUuL94AGXtPv5SPidpt2Az+jrflIe9wG6knu2JWngnMGcgS
mVNRg3ikSI4bNm417boggncKZCen8tJpxZFbip815f74WOg/DQ+N9eE4PbyS7MiUyqhR72Mw0PL8
kx7I5QESsges8LHlUEcTzRgKT6JyCyzLPOKSaEEJ+PNbr20Tiuj4LcJRV1crm9DWUiNrcNqsWOsQ
DVVFX8s51KCSbrTDhI1hXjFBf4M0AFDZEN6YiIO8+CyPv5jvdUxjmyhgWbRUIn4QNEOyljhTdP/e
BgVSpgu9VB5M/hm5Y4gb7XKI02BUK6YVPmnMLqN4WNAlJnLRfAOvSiUEPDanlFgbt/iVCued1rJh
x2U7UuyayWrVPs6X+OtojO9XouZ10klBeovRas9EVonxrn3JPKMD9hT8y/7+N9inzo6tfX69sUZY
ZbwW9ZbxcbBupTci8vtgiAx8EVrJtIdaSvlz5DxwcRedJQJGndkl+/7NuVnkz+eci+OStDZww0JK
5DTs18sIjyj6mJcarYBbvwJnMiJiu69zUSYu1705h7tWZgXIV3PSdiCDHDBGamwwdHm8RVAHL1Pn
xraiR0EXUoLrSJ3z9Eas1RMh/H2jDmfkC79T1gMbdIG6rya3XzKZvsHOj73a8dTM1fPT2WJfB9RM
3PMt2ncv5FiXZ6MPDYyUujPxqneuQiRa6BKYobVe/DNuXzQ66L51qMqQdVKtLWAEKHKHTERvHpPg
tjWFZ+H236ymzlG+afp5ecxN6NW/fPkzXjS066iqnl8Xj7jhZ8mvkGWscdkVb8Rrfl7m50s2nrHW
Sd5ehNYYab1uMJxzlV52jNx3ifcKWCuSpxpRI1WhIbBd/pNTc2G5d1EQlASpkPQvLf2KocEXEUgr
Zk68x9Fj5VU+DdvNVMJmTyELw2jfsjUCgQrZV84e/R+zm2b/1njgj5uzzHLgaWuzZOFV+B/ukwYy
OVk7LGe1tCUahLeaZcPZLjINfGrR5eweEZ8gnBysTTqESmCTCwcs3kQLcYE3umKZscoDXjR36kW6
iFRH//Kix5U+gtrePSKFPBp7E7upIiLXV6rDb/jBYfhL2U00oyPCV2dsEJWoOkzC+5LT/tOClRWd
XqHKR6cEFQe/85XSfEoBbbxIYB3iyzo3InoLCbR6WaNgyopCHymubMXT8HBZzWcq1TmFF72adOt3
ORH8BIcK06LdalJFw0cXETEfD8A380G0aYcNMGlZ7dfwr6rUJzx5U9TrDfDIaYVTDwo0t5pGmTA9
QaT7b+GwZgFM8pSmxg2C+pzd1TTmmgcGUdiW2Bfh9iXtwMMoclcfXlRyQd7GW6EManGrDusZqMqN
OXBamEezpVxXKg4+7qYw0OmE9KSh8gHyEEuAaL4SvDY/fJwWBB7Orwz2bkmHtITcFqJeE0HX+OSl
okUs2kJPVn6wHb1f/U2+lBOk/e1ACII2SxhUF1LKYM2pAK9gpxwV7gvgMZwWYaujiE+bD4co/mAF
5ZpiBhD556531JN5GgR9QTVvwRmBUoYBzqV/fx9Xd290R/LWfgrJ9GqV8hAjE1mdgIUBxfxqwt6T
vdRvjtNYjTw/UpB7/iVl7GqYDKRnL2lQXYWtcJpvfmaGUL8AYboeqOyrzsWE165Y8KkTT2jVtAEX
4PxPdoM/swoWJAAXE2K4axBmyr1qjii328cdmkWRaUicg4ZAI1pHwTn6oGFyDSDyEY3674LghInf
l1MpXtwFo52k/qbDIiMi1E3I5VwwRKgxVBMTyaWXrN6f3pd8Q+743YomAsQG7tRplArP1ZQ2ly+j
RLAzkuSgDj/X1qRTfyJD7j8WpnaVMvDZMPbgebicJkgJuh68Mz46ySx+rcJxV6xTPT3pr6x6OfqD
f7SRryecD46eu5Z7XHn8GbCmr7uzGbf8tYG7SUH/Lywt+uOj49A0ExDD56dW4wHpsQFD6OYQoAAv
RE5Vg5WdcrhTE0o/jNCPBBfyhveADXooqo12EkqaCBSRCnhrQY7Z8cOPmhH2FQ/plI5OVTsVJiY0
llMo4Oe0UdxDB/VNxO+Zfz1GNHYyApdDwWMpnkEJdZ8dtQbxqpT7qBE7S9PtxKnRfwa+3ki3+4mW
S+dblPCxWyMuRvNnDwijI5S3lhrKXxrc97V9whBGHX9OEq/ewn2T1AVNb72nNf9NsqmggTXMlzb9
YLFuBmRWq9/WDX4C5iC1JN8EU/oSGh11VIPWX4v2Sd4oKQbsS+SmW2agGomadTGDt6TbIXiGiv67
B2FRvaamb7gTbtBivxH9Vh/+p6tvkAmhNkJoaqD+5c0k9KgQg7+7INCnf87oM5L002TDJbgSdilA
eu2fAR6FIbhwlIjr0qBovmTYv4J6j7nYZsL8rb2ogROzVnnkKGw1KJ44U10Z3VzwqL8QI3ra/oPj
b9G2upuK3GnDpE9Kuvs0qVwL61rM4WGEJce2F39unpoXu2F2QOCuzPCnFGYg+z1IwI6HiuKLUOYQ
Tfd9D3kJSTWlqXMP31Ls8/FU9x/Vz2R1Y2C1Cf+GnYdrDC7/lqeCEixDGJu7U1UEOIwqz1znID18
CWf4MAoQPLkt2b7SdqDhseU++P2jq4wvl5rmrDiKj94kRm6Ol4wtdFYrgU3tD4kLskUzPtJK6Nfg
RFAB3q+vgGrI2xmfxc6Xoq0w8GzZyvp7AMpHk1AhmXimcfTEGFW+ZC3cBCSkkQt5nIF/vomABNXn
CXDmVpjd/ZOUwKucDFYo3Xp6SG0dsVq3a+dlt91dDU0WDZl81b0WHBO5GY7XLC1Q6P0o9AuhgAUo
1oCowNcK/L6GkdanOtEpoFWwiomN+nRKQaWT4XQXJiNARzcIFQ0kHhCb/ZAQQbkh/7tMunWgYj2U
eZvUJKhHJHdL6uCK7FP+zfoFmJGfGEIW0Xr6EArYZximbvWRkIj++KOLE6q/p/XUxSUJ/T8Qf7/b
lM/o/8gBxCga66x5ZiJeY1sBCJfvPLstyMPCuUEp27WwgLv9eZwLcZzSHBc+uhkP8XRg4ZRdcQ0F
kOtprryrIkwGx2PIwA2LH+Q0xP7FwqJHs8WpeUSb2gDE8l54GNMLf3XwXEM+6jkVu4YBy7UTcCDu
SddqjeMsr3FXTIgo+y8t6xyoJx5kJeKGxVeFTa7EWiudZDM+PtSpbeG7lJC7HigCK3Oz3TfOXIan
cw+bFJxzNliFun+zKKOES3JacJyDKNyfl+0dNyN2ouf7b41AF9UKD2GsG2Ok7x/pfnAQDyotW04i
OL+fJeVO2L2em9vBbBgy3SWN7qxmyFGBE8tPRKnrPGw9GKCcz+w4ARrkgrefkGlWZYwMYOkkUaRz
5MRbA8T3Xw6cqtCZGbIhs2hLPwFOPX3UX0iccxG2cagxBb1xVY+/UOhRffC62IMT5SDhC8+nJw3e
wGoDJ4b4tWtSmqV+ajLDBLdD1s3G9BzZQJB2A+Ys2E5Eu4gFhTqkixmmCWtRuqZgp6EvpuIy3X10
0V/BQtJOtTLwgj2ywzOAYrqNYpL2YlWaPG4qx1p7RNlScFj95tMKvP+XAr86K3b8JrqMV6HVZv92
G0TBNwRJAd2uWbb+TtTKw3rFHC5g/TvYJw+H7gMcU8Nt/5H2n9bDkF/p75n1QbX8pGXLjJEm/H2V
f5e/vAcDRE/yKFCV0bxyTE9JTlaqXdwP5AYF/4sZcamaRJkqB/Gh3/Suc0ROv1CGbtMC6dzizaVY
AzUII3G3xMZ1zKQQToxitS6UsWrtJKz8EvAXD7tuwb8G0AvWSL0yar5pj+gsrrX2OQOHPu266SWT
92LSH97uhwVzMUaYzgjfDolpfU6G7KEf2lP8Ha6NmHppCSXhh9T7xDh6a4xsiMhajRCCVBECrwFi
a7OwBru9f4XElvIVXomdo4mqNcE6pZVwmx3t2pLJXTiVIRyiAlSkQgp37MXopDSRGPuvaS8LZjIT
tYnMbS+kHL9a51YK5OJdlagK4vZWfQUWulec31qaOkdieVC23/YABE6V7RTtHOYkZDqqh0G1KjsQ
e27frgeGPE9/amhLg0v7yqqBa96sVo/ziTrZQzyYMgPb+Ff5seGHVrn91svMEg4AupmYwY7qRQf0
2BylKSjgMJlFnKieAAVQ//f7POrLNH8Ln74EAi+GXUpVOoW4EA6qdqohHd4jPVvfVSKagHetCGqz
IT87SVChV7bN4l34SSQJBEO4S1IvX3cc3TRmIVsZmwZm99krMw3nuubb1dRCc2kDi2+W09Z8FNOH
NnnoWTTBiiGisjvT8YVCattDR94cF+Z78f/R/IyvnabT6GY8zUoAqtIvEW1GJzDjv1SZBfGSnpwU
PY7uOwluFAhOHjNGWVz6MOvrXAIIZcT4bqx63P/tINC5+3751yKfL8qIv0hJiBvFvuPCVy0LjteK
sSCIy3eexMEsGKqAeE15wNqAErPozIlirWTcAj0gW3EDidODMZ5qUCN76OEjp3Jrz1YxrtzPPPpv
CTo9390haa6+PebS1wnYGdYKBhVqKt+DfQ1eMfgEj9zv7EIF1lmj96P2N8viRVSb8a2Fi106I2ob
FjV9IEcS5TojLTZdf5XUF8dsmErJzf+i5k1upIpbRJ/U9T4LM+AtUa7JHglkRi9ZUKbGqyq0RdoN
mel98fmCdRyiYymkmV/hmJJGag/gF1JIxiwVdUeh6HpeWSF5RBuxGG1dQNR0bc+EqoAFnA2XJEbs
g4+FVu4yVZ7cPqiryp4m7KqYaJZ7aC9fh2yuY8fCGpM8kYk/Ysh/mOz5k82MPY7m/coyoLqz9lQ1
LEo0Dp2S8t88AWGOHMyMm60P1gnjYQPiUoMo0+cyfk9eqR7Wgy9TLZIgOgfYVk8DiC/xw/w/514q
w9nGquqdISXdj95n0ajGN9rTTi8WpR/uYj2poC+PqX9FUgvUjZxolqMj+ScmUbC/IKtSdkeyOMeG
lR+W4ZCFQwlOtM8MxKWoAWa6cgQ98UXQR+C2A345Kpi0T6kF74krlSPSAThk638mCIJl7I3LTZvw
u8pwZ6H3zTjvtdraUoMZ0IkLrTTLp/oXWst/IvyHOCDaewydrTKTAT2msbysiI0+6X9Eo0EEZw5Q
xpOa0NbPsVbafqaVnsToE5EXRLD5F/2lAA8M7mh0pHWv2xPAGOyZ2+BqTyqOARaDr29t0xKqgvli
W/vNJnZhf5jPoeazfA1pgCtjWUibQCxYWEg7OZeFJfICwy4vCSbhrBFAIuXJChu39VuYd/6NrkM4
9AZsLeQGXImmKmxODl3KtRyz3kNrkaRRaMtV0iQAEPyUqMNNXGo2MVub0yN8OEThZmGGacw+6Yme
XMd9Ye7RMCe4H65t9oeUu+3pZmgO31EayJEH0ayIfmoKzhBGh6Zxm5c7Xb+5VPVvHTBAEwdKbao5
/2CZ14ZWaCCpi04XjvMtVdhReGD64RoAXmdDZBdkaUGF0RQqquEGTUnbOkbiKbKR4bcmbUn7UqXE
B4ySJtzmvo07MjVorRQYWwmrv/hVIgQPER+ulPIcL5q3jFqnCYnUvIHbytyUyRb/oGsErPo06Duf
0j7RdMkhPUAKGQU5mgdLglCOyF41MF3h9sO3VFP/Bub7yBa3USjQ9XgkDW0RC2GRZCXttVY/KIPT
zXFZ4d6fk8+2fCXoVS4hDcRiSEpnDc+tkmksxKR8cDYcZCUrRV4S0M6/h+17d3nBIbM4dlnaVo4S
IwtT2IPTelhii0jlHrIiHSAVDiBRktdecag964Qql8NEqpfONUlKFSXjNrfAst2bl0Si54lN3yiF
Vvr3jVJzSoqY4H4IQkg82R36DLCHTjGVYj5LRLVW8XRVEti3M2EvovYQKnPLVvMdKINMzMZsBA69
4+M6iDXaB+NbDvZTC048V7YSGvA92GPlsEG08pRr3ImHUNiWs3p4R2fZYENYUpw2JPtS4Qz95552
45Bh2lVASAEtHIByEV7wwC63sx07yyClkLD1rsxnVygofk8ivIw8vfy1gBZr0i8Kq7PakqNDzKYX
EqBOLX5DUIHeQDDEIN6bcLbWd0nz6Wwj5zxGpFROPeIVNuG/4h1xUj/1sVKjmvMAaWj6imzjyZKX
DQM3OitMb8V8mV8ETYo7w8vpabGl//xWxqKkIY948VQmb16M+0iTXj+2AAwbxUkHFJkmCMc5DQ12
LrA4sGPHq7n6g+Px16PtyFYjzcO9R8yqsVWBJipTR/hM6zN5tRff+VFo6PpQ5OEYjww5NBr+uyOt
qZS69im0Lc1ZqJV0n2Om1XHCuq+rmH5fYw2WUX0lpZXmXMvXZ/xr6y4f6NJJ8RInrW3XKPNt0Dxf
uIqdzlq5Li4ZNSku69W/HUu/Jz2F6ljeWM+EgPvf4uuJKoVpQY14HYMaBdNGyjI2Szs/XsPg3OA/
V22ReWxoBHwozGFrOaTTI/Rbeo7MXUUNZFCPGnsLkHb5S85QymSIBgQmsWiFG3nrNKl7AkNDqf5k
8LjlBfuHIlG0iHkjuXkAq5Ncdhw8XtCC9xKODM11j2FCebBPHNGBTi97+ixBzd2jel5jg8CmMjRE
7kmIkZModntD5LajXFF8DNtFY4DefONVoMX7pswC34S7F8CCZpiXhbojBcb2YYAmH/P87fzy0rBL
Hmfw3VzX0BPFjWuZgh1gARY05fwJxJxf0gY0GHMxz2OTq6rZlK20A9dLqBx4l6TqowSvoXVsZILa
8GDKuYNcFH8Xa6l4oQK2O5IWM7KQ/RJ4B1T0Sp/t+AIwNEQB781XE59MJpyUKmQP5rPjFr8Zhzr1
AqfassHYEjuKgzFmZ2V6Xw18W2ZoX4VFeSV93k2b1sPPqDwJn7qdqYP6laEwy6YxZupF5POpUw4u
v9LokjwQF2yauYNwHAneuzIAR3NL/YOFxvFQW0Mwp9BKtMQUyshKY0lBpWpbGzG+a6L9Fio0Kak6
0IZD5sNGi1nRaqQK+wsFnKdgr7Ioa8t7UW2h1x6k1lG0XzZmSJpbxgsJSTLpZPrExBkfrx2cQycT
In+du9fHkYhLfLUi1UbSdwo7lxahkjCLwwn2PB/Ub30a0nUZQEfyTL43/lSXaXj4pogLraiHE+8f
P8fTQaQDtT/OqyosXg01qDQyrnc6PcDnxYahqAB4WsDS68cUX6lWVNMPy9HoXz8jDDR6a+3yZtuj
ZZCJRDQF6zh0ShFLq+CaiwpP73i/YXMZAhzyF9jtBpOvuy4UVARz4sps0CxmtKUHtleTLgb+scjv
QUUFxu2SVoBGytE4q0Xn/lvTNEQsEOspDDCeEDbSEIPQXucFEQZYtgqEkfdahA1DEAh2Lqsa5cHN
Q47kFSAxbXuKZ/I9CFQYXqOTAmmHJ2tjJd14Z1ahmq7VaS7gydY0wMBriLhpG+fpl56fnfJNETfk
L6mDBjmNqWWew3dOnffMHB1TQl03oyDIcJthbmd3x7XKtn7HVP4nakWP5mtz5szP20TtVZAYDS/e
0SdEwjeQrHmxtqSEGCN1S+zL0TeTuSJ37ZzY0hAybfImovMFDwaw0kC82HtriBUAu7T0OgiEdnUY
RiBbrNabe7ZGawaaOlBkScpV8oRUcMYcznL7wyPqfH4+1iYPex419hCRvDJ4WaWdt673MLdI2xlG
7YsAo1OXlCdni7c9dH6KhyAaKiWwTgp8KhJJG45KsiEK6zL8cfsjz7mjvOp67WDbfwQciIcvymFR
9w6TGgyzoyis4e2YoXg4O+3yGqaaO1GLr0rlkutQdoZ0W1bwKzQMatoLyuCAK/lTH5fXCDaJzd6G
sdJbSpk9tcCl+14pAlcLCuOlVsgvlTbEG5dqimzSaONh/a9LY1vltzZ5vP0xScW06GYCMs8wr5ZY
O4Q65P08WqVAYkM2VxNJDBwiVKNbez1nSHXZNfN3EuPkNq1eniXouUA6ADXrbEy2M7Xxp5okroHc
h8S9KSy9TV+FJ5DP4lYhCzJX350Ec39RbGhWIlI+4O2VGlUmG6oDLtCMoIyi6mwXJ/wBcN7grGcg
ub8ROg4ozK1vC4XYf7qJFcBPhMLpSzpItsqPgaWz5m9bT6XHwJ5xpxiSDUwEYjmHWk755OBGGwB2
N6JzVJkD+GdgUbn5+4BJHvRCyBwCfaY3uaxgU0laNdgjZaRyDjMKsXNBuEYw4hoYs+84JIOHOGge
c5augVZERzuavMdh+VyrjOTXKcpGzMaHg1eOEc1TsvYcD6QBxa0km7xC2Db+0lZifWVSSQ8m/Tjt
64N7nw+FF/yVZ2wcg3Gs8Q5GND2EsjPy6YCMM8Ouw1nqzfBGeRjSyeLFGiMA8/l/bzNSEOF4e6VI
fKpDISqwIm6bk2zBgLtZpj46NSDVQjGeyib6wzzv0deaYFD2Y06kQ8ehs2oBDMqy1Nrd0jzuunx+
Ml92GzErGHmOwwrNha6+VXUl11+Y2ySGYZq2uNktQfUf52Hbacrp0mxx8/2ZxiGsIi3efSFRH+t4
Reinla7fezQP1hvYPaL3+aPyDPye9nmaQFLP/KX2mKJzpS0xQTBb3JGkS0fdnntbqjP+rpHtcnmt
r3EMAD6Nw06tnnWASVeoLtE7BD0ePwbEPAEWM8IxOLwzpv+R7TWLOz+cJ0vHnuAP8PlDuXrPkAOC
5Iv122ffMtp59GL1p1U7S3XrpgnAZAVxDlflYx0MSUf37Wey0kzuJ7O7ooclOKQTMXSpILJEPPEW
geBph+CarJq/lk6FokyB5ereiRt76Mk+dweWUk7fkIcm6L9cDvpfcOqbYeJ0365CLuchER9S/Wle
PpcPS5jRRgnwETuRnyaBP2Rdiym4WVDjKTR8HoisEhu21543/1BlpMS+6bcPCi1DNDrPU30eoo0m
rk2phFHI4/enqGfqNaSdRB/ifaNwsus6ZJi89tP+oOvhdyfR/d7XLJ2IWuPrOfg0iNYcgOL2ZWdw
hVOr/jWPu7iZK+j7j/Rk+5dLXWWu19JZEianlw9Rq3C58bZh4B4QYO3wHzdi/rpcKzviINa6Vfk4
13kuCiyuZNksF1EIByWtuCWsqCzhddF4D2Lfy+qYcby2Zb5gzY2aS+Iu2hrZ9RTRWAB4N4c6qfpC
vuffX40vWMHL5EgYfuWpkjwIMmCEqPWYY0qLIzYHfSc+Q9hJoVPD3QFQA1uFEd0/VyRRmstWYyu2
N9oVL5NgKpRu3EGSDUKV8A+pc0/X/Hzencf3FAKC9Idh/bCpDNyG857APGWNcWAvYMx/s1EQ1u6z
67FappHAtX34mJDwOIMfbw0RK0MpNCTKvxMzpSIkv/G4g5VvwxMe28dJzKkc+JfBS/njWWZFfxtn
hwgG+YAsWYg3xXw5QBhI9doPHV1FW8zq7MyceQ/OQ+LRC5Fh2nWp30Fo/MbhsRhXJ4b0BAcfSYDx
LqwMKqeJogByL4BfjHifhqGFjc7ZXLrkVXj0kwnhVxMOWg5zcvIfSb/ct022Retyf+MOr7maYkbi
S8mJX31Hs1Grdutl8NTjM1gcSxFw43nuSwg8nN9IV3jtJsAUBLxArFGYdRThveo8tVh4/ECD9lYR
67s0VWXirnRsCi8behEzEHLuCk7DPZrgZB8NiU7n6lI9yTOSjj/hbwq1M8hCNFdnVo1PSRYELy8s
l6ePHLOpx4Sm2VRF1KHVHpczq0LiKrOzHp/JaI2O4oZd0WDtTMlGpEbxCHh0QeJIx1rEcChjZfCW
fWbFkyhDyuwYuS4xEWqj3a4Y7kHL0yUShRf6ZdnfmCb3/q+ZpBnRkWoI/3VNdyDiDQFHhm280sz/
vGeTCt9mdoUyC1Ij53JMIbJRkLEubrtZxrEe7oz0QEVE4pp/BuR+xmdfLrqKPDAaTk/NBH4XTvXY
2VvcM/oBfrW5AueaYJj6QJCiW1zXmaR2xs9x2hjgF/vGgLa//sPsPC+gBY9mJiL1T0gnA+ATBLSY
33Trg5595hNH/JnxqfSaHVhk322rCpbcGDKAfIBVHAth+czqU9xx2Z73Tapb7SsU1hq01GRPOGTi
klWikB3x2LcN7mcwO7Wq5QZizw5xv9rqdzNC8lmYzjkz2TdjYBjpl3fO+DOQw3KR2TZyM2G4YWSi
ax3/RakeEeKVt4BsGue5TXMMu73ZQpaKo3bTB3GREGQa3hxE6aow2idZqMEKI9AfZ/sS9sOlEEHA
CSzVhMcQKaJZRY2U/znVAyfBoF4HpLH11VqX+RfcAjx67x8kEqZwiYa52i1Z+2UaAGWgBqObzJJz
TD4XfPoQxcFvq/wuvUJcisqRe9c7pHuGQDJWhWkjrwQJBZ1goZHJjtvZ9gmgrJdBtwpHfjQZsrkV
Uz0mQXDo6TaK/n1+EM/kyzbzU/7slHnOQsmkpkQBGibMbzbITbRwEPBHjZTiUYiBuCPkvvQsco0C
QfCAJuVq08pLpOyfgv04SqJqqScfVBEwHM/PUCZSY4BwHJMZxBCNz7XUdicOqZ29qdOb1Vd70m6A
ARTzynqkXgDBqDlPh5Kt5EblwaaDqqhOJHtP7P5wu8LmhKfjlydsbOeMAigy8dpyJCQ/xCgCstUw
KXh3ubJSerkLeZOsbdO3BHSuJbNtj0dpaAfhyh4N1vGlCcSt5N/rnQMGJcHzaABIQ4vln8n8EMhq
f1iOrb2itEgfmWNE+C0lEU4Gpxk1jJuKxO7UVKPzm3XhfMQD6CZg2XhbaNL+MIAN5t/NCZLLbnPf
S2zNMmGPDz8hvlHFBMtfWR27HZAj5E5frcncK2MazbVVflWtDM++qKGbHK4V1ockG3yVZb/04JA2
Jvqel5AgpskAYS/U1DiTfEmy+kgOgGHT3XGXMKZgdB/z17vLdUryw3UjWxBz+a7oaobtmYkwru1J
6IMT3VgPVEPf9H/Pc24l/wVxl4zPgmPwDaOmz7yEG7/1BuZqR51gvOexk+/HggRdPEwnqkPU9bBn
7b7SxQRE3l8151yjZoQ9IFtUTPJbfZrZCPUspu00Mg60NdS6rRj2wYHVR63zrU/OZPSYdMcphFBQ
RH9Iau5BP4/tuWeqdlkz52xWO1Y6Lx5Dp0KgI7k9v1QUSthXVY1g914eMgjXudJI/ueIglrts03K
iUgtEy1H/IYUlXSxT7DUn29R8qBG299tt2mdtXHP4VszF9/0EbJ/XUsIkdTCZBQLwvENBv/SGFBs
AQs6HssQLZOXE+cazrEzr0KK2IGYTsGyiFzQmZ52fFcjBPX222fnLESPgqdoCrGg3rTppJOrcSSc
4bUrqzsOtY3x3RxodQgta7hFJoZj0um9YpRJo6iTJgnuHjQRV5ivqh1fJKd2/BtH5u6p+veF6rl5
Er6IYpvDDuPnM4mTjRglK9byMnvq+KhMNU6Xj3J9fIrrhdNybNTNuEqHmKmC03GkCiHalpco9nMW
fP9xmj5tNZ6hE0eFz1AC2B9dN5xQJ+5zSU48ZuMWf5/B1H8Eu1abjZQV/+ih5aLbYE07LKKtYFwZ
GquuXgARP/CC3b8/LEGDYFk5bLQl4zXeXG3/kXaUnL8+XTbg1dZqug26lqxR7XWogm9Ji4gFpFIW
Xy2JV72/Q1gb/yNoCWNQqTs/wx5NJuD4+COBzYgpja14cpDAr3slilkahSue/cnzzp7ApiOhd5FI
TBiEW6r4Dv2noveO8clHPYjzmqTzAiJzB3uT0JWGjShC25Z/vMXT1aNF0n6dsmHJwPs4j0g+Fc0a
YdPjHG4qo1FQGsWWexgk8Z+/N10KhvoMJ3I2HbMSGlb9693sLXc5Uj1CfGFHT4AMNamcOWjEXbLA
GcmSV5CqbUqG5R9XmzwcKK6aJsp+pwUPKA390CxoKxgeNHu2B8dmNhN9w3bSfsBlydq2VqQ03mFD
fBPdqy3Cn7Otn9eLuqBKwDl25nF/WJfcrDZSmBIEeu6gfLRB3Kns/+WrWJof8v8IUZ8Ypn8aePtn
GugrkABlHtM/2M1iBoOWHiw5LVSHNFlRGETYkitH1yLEpXjZNwmA/Vc0CI+BWayALy0O+2pUOcVc
TZZFbQzzDRVFJ/xPfJmOfndcuJZ0suNCQIN87RXQyCAkAoH0zdVg+KTZ2vjLnEtF05mbFeAD+E3+
Sb+HeXleOXhk3Mvn+7ncZdLNomUlNEI27DUR80UW7GPWGlJBe3YbBwog7gEnbiXnwDBaCIlkh6TZ
FBQbHTkAxuqzjSPW2SrOKPlJwp4CZZxiiFf6h/9I50Ngsp9lDFDyFQwrtbmgQsH6SbLpzsAv0t3b
p5k0JscuU7MNt9CdDSnBmuloO/B0KF6qJUumi/CXgk95YmHrLw498cEzkRRWuS6qRm4uXpN+EB41
IDYAvo10cKdlf5gTEZixlbDdr9O5T0BlMICzgKbq4upl3ftEGAuMiSDR3EGco5W/0Cwl5pjWmFZG
JkFeTV5l0jHeZJSmkuH88y0k1JH8laX+BGGIUml+vwn8oaitexN22wHIkUQ5Hl5thW5gClEnhcYR
sTDdpezCvLFXw2Gmi4vBBB4KcAZzUUZ+WuZK2s27OzuitNl6EpQiW8HWtmmKO5VUyCAFiG1KVRb0
KLJWZIYRKtbQB1b6HnJi0QNsD601i480CdcKeuOg8dOZrUq4kkJ36MTgyfBevPtDANWyZVbtnNwu
4xVy8oBCBS5iWlC8XWVUw331CG7NE3pEh7DQgM8fx5ixU28fb8i6UjsmbHazn2SBRyre1CizmiYq
pPDoluRtYopT3N8CpsbxOfAgk5HumadJclYCQkON6YvI8S7P7hNJuxvV0e8C2d+cHu5K+4jKIY9Z
TZODc2F+tDHCOyjoBepmvHbf4htp5cNePo0vf7rxQQ5xnSHTjAzKnEZPefP2nm5zzXy2bH2nCYYd
zL8Vw7AwfOESGtuHARhbcxoUZ9N/gA2Vn310yyQolzytDy8mXTCO9FTjNhhzSDB4oLDl9EDo42Fc
5omov9diMmBgunY1RbZizFv3lXHHoHwZ6BXVfdcCWRsDLgbYsOC2hPJjXRHTTNAYdEWONjIK705n
ZAI0NcUTC/dk29TTv1i2BXzy4wlrnWzFxbJASy4vWiAtpj/yVqeSe4vGBGbOPvPpl6TtlfOkB6F9
B3Fnv3NXaqqUaHfi4rp1m+j+QgFIev9pCCnbetSMZlThvJiCeLh4w3vvmuhpjOh7fiCrz102g2dC
gbNor7cUKjtAFIzvMmdKcIdGdLiNtlViuviG/Vqj3Uo58RDRJjbCIC/pRM8dmAWtDhkoZNngfTAP
ScGVZZ7UyGZd3XjFAYGNVJC5Zfv4DQAT8xRCsScxObTtuvSe+RKNVA7CXvqQ+u7GS4W8FTn8lBhu
vNgN0/Ukp/3pkYTaYPTCFKxUPAq1wthd2hwFqhyA0L4wRiZxL7e0iDfOrrznETckYS6v5ALYPqWq
SBodsa6s/LBL7KCwurQMo3Xdh0o0M1/w9jb6Fx9ufdXfThwbKUPb8+vHci1T1mN5qfi5B2umYSQo
fH1LP0p3Iuz9bgjy0M94MkyzItdrTFnAQ9pQ8G6Nl4e3MTXOww6TD5kwQVazeh9r6LZnlJDUEEQA
fZyD3G6i/N8cnLDmyLdtxWxo4BsDxJFFILuMTrBfECMasmWbJW1abyuIipwebEHIy+VUTe7qhl6o
f5hsXSixX/VD0ezD26jBFN12RmZwG4mh/dYUgMwwlNl0wEsBmKcjUlf5nsKL7bqEnyGQHiWZF/BH
dSXLIuTwh+HtMtyZC/L2yLacJRIb4L5gPSW2wA5NBDyLgMCZ0hu/PYfnFLATOLAHja19rz9cTx4m
QZCWUZABdwgx02d6W/SOXRq95o2dalqpvhf2lVzABsJDu6htPt19kWkeYf3E8QT9LbCGdiYj3KfV
e29qwOnjeqt/a69Ds1Kj4U2PwSKRP3xGfFH8HOK3QMUnGOc2Rf9o3400f4c/pEFNkEDOzAa1wWtO
p4RJ0XeaqzFG+cYiFeJGP/ImGmyqO/lRfRNwKXFial8fUoNCGc8QUsP98vMfgSKkKzRrDf1ywYnX
dhmPzrWR8WbgIvZxdcLRLB9A6sazPoztOXHuBXmRQscGdiMuxoqF9na4sSwvUnD5slfnBT28IK7L
ya03nlGErEQ6/NEeTrzTMfOlglLvRV57I7Rqix1q9t0Zvgq6C5qcJmifTODm/5ZqBkSIMSqrflDJ
jnqBei3KOj5x7ArgkaUglFJ50HUSdlNSq0sOuUsJbTAGd0BahcGMCoE8jJrurl6s9KxM5REt3DCK
+yYU14quoevaDHGApJm9pvMzxGXvxS2ZoTWA2jIGJnmcmxoHvxHRQmpkRBmF9aDHoYI5axzZ1m8/
I2d3ZN6LGlZKdTs/0VgHeHIO7CrYQXrOqsCDEI+2iFlPi0RMqvZ79god2NwYcEY75ZlmQ2PBMi+L
1Jkhj1mzvFXxPUu+Jby+QMa1/29f+BAfao6d2uQaX2keG4sXvS8nZ1zbXu4r7TgJq4BvX4GC18t3
ndtCmF9dFmNLd9LYucYCH9zLsMx1FcpfZ50YTN2qtk/EkAq1R8yRBOkjHEDzvrsotQO1LCEXBT7R
d8eZsshNbEnnLB8rrCauLpU1Ff9Q5nLj0vp8azAqM24eJqFqvU3BH1AJ3OsJQvwyot0dqQq6vGca
+B1/PhRZQ8DbpWglKPyswIXM1Ao/j/JbCRwV15QqQS1WHwLsODNgYD/+Obrfw+WiZxOGSEiTXtjd
5L0yu+BzLUs50O6iMEoZ7UeQXUT9MEtKtmjBrj862Cs8GDG7VTdHCdVMBL7MWbT1UtE1qoS0BB3p
Jt1zUKqTedpSr54OQ9W5pzrDywX5C6Q1kGjhnrRjBbWk9PMSx09tC4W/NWzeclAQ4+1iEFv9wzT/
+Twi/GhbwI2pQXQuUZ+I2yJuok1AOcJ/nbiPwH4TO5di7WYhQ/b0Lq3h997633H1wu8H4oVH0LWq
VLuqrbYBwPe37GADinYa4vO0CfO7X1QEtbmx2r6W9jlIKOBK7oP2sN2ySqsncgwfTr8GCV6NMVMR
yZpH+vk73n2VcySSgJ0ozklRWJzpYM3+mJnQ6C9D2Xyo6rd7Arbhdqev3lCsFgcWjjSVS/hvYI9f
KTjo+1kIY7SxkIACmZF1tAORsU9Klf2d9sd7DBCtYA3SwHsYiuwLPshkzzUHo/gJTJaW8dpY1SXH
p7ZlQE/SyYxjpyznjyGZxuO954SygE5cIsw76dTNvdli4XgLahaqnRc9KkJZGUR+L7336ZZ/XyxX
MA1qAWyRuGQNxdFZYtxNusSdMuy40sj5hinXCx1zrCqjN46zMT6yP9QQakiPN+isXT/BTjtfDxhm
YWAfI3tqLzZOHubaNVB7PLMDoa1YHxBfrLARd3Amu2DUdagGMhjxZ5uwQDJSqZowRu1HLbhzKy9i
yEgADaVhVk4WJtcrOpkXIBAoN/6uzQXmwGpE0R2/p2+fhoqrUtBXvG0jZs5k+ZJ8bFZDc+gXcUIp
oLzElgmUvGFFVhJ37NNQhL5J+LMn74e8VZKFwDDz9jwg+lmj9jnp7vMFJU3FOGNkmp85czKvI1Le
PTx9kaJK8+IupALDWBBxGkVyYFcOwAQ7wZXTkGG/h5BPP3yvTiD6CwHLPSdBCxGZfQ/jfyIcBT3g
NDRi0wDvqrXZ1OzJHP1DnTfD/Do0XiI7flBmFY5oPLMHBrls0Vqq6HVmiIrsa81a5rGseyceAnaE
Dz/8dbpvzM1GjLbuBOV0Y6c/VsG27xPg11d80YnopqhYcxHziffJGKdfShQb3LWtZB0kaiDKSIft
GsiZPX3WsJ/WxGstb1p4i2ahp0jLwJ4OGYEIDAFw+qXQBjFB/X4mBFJ8RpKvekjTU0lHEHna63Zq
QAlVnNIL2K+Rgm9rUHsI5CzF/MWChioMFoBanatX0edDkyXHserNv0100ucKZmFM7lACwTKuKoX2
wEKlNtUEMHWC71gCAJAvCoCZqOOHT4DF+beMtevJUIXv9KXqUWNdZsXohXKv1eGS3vUMP4WO/Ey5
pTcQP07SYpdEB6EPAAPcBOftaFFK4NGVfjeT32cNZFH7SSsMdudf1eoD/NyJb6BXRatGkNOQWBba
XaIi8Pk06UHv2faNBvCWKefCBNokXukeL1akKggENlmstIP6GV++4TsQQ/Xq7bdnB4XJMzWqvPS5
xRQfalqIEn2j1gpd+LrYGhkiRDaKc8OYlp1CKt3AAFQmmffM5Dyv01mAcmysO7UYQXS1UvXprNdz
wXv8O8usZNqALF2JZIwkFDMNddBo7FcTdAWIEWFMrcxhqRq2sIbkq/peoLVZ9Dpaj1TY+s0G9AOC
BE+nFNgfOqcGB+OrFc9ENPqhv7Gz4RYYzAY9bh7L29rAo/F01aRbGIxOwYgkCpFDmQS+TOSlxRTp
rkF/DHlHogZT+wqBsmsMFXYv3cYAyky/EYFDt9NKKp7/TJ2+aY1nww5e5ak6vog2QAyPFaLfEvoh
/8OFT99Nc7l2RSXAq0kNTSqStphoSjme6RUBS36CZGyw36gaiG9wJ6Hh7kliO1MybAFqB5zhS0IL
uEq+zKsTppaYCumMFtIqO2BsDDsUo6IEahezOUrCdIsUIFMZQXWBz1R/eVXe/8Yo9/Gx8M/Q1O2+
IWljgp+Y2gNWA+552LbyZY27BFK3zXsqNq8fo/7Xj+NwGp1336LRvBL4S1kMsOzAYDanpbyzBTAp
7oFqXjMKCFioUfLcbaTJGkoDXat4plIt37M8cuGeYSSbITW8aw1mKN34nRwWpJhF6XRbeFKmpLNJ
nJ0hIKNGWr6RkJlT+p8LehC4mfw0OgeoIjee4cii4CMK4WdY415KtEDngPslPNvRdEyuDKXs8Tk+
RH00o2+72iO6j8D6jqpReDhp2orn+eoj/SqFgmQ64i2C1tj6Jz4jFoQlJ6Lb+KM3wWwalhr9ZOHl
uEkzruqKBAPTd9Oa/hQ4umluXmwntLMUz9zJ4lfIgZYo/L6VD6mkWzZD2hxvxSD0yCCDV0ZAOImT
cfjejkc6WoCm9GVEErh+RNzyBC4pvSXfQfxao0emiXBqGRRXxAqtQGXkRS07O3wb02S0y2SpDIbk
Nfb4KFsKn4HfKENcKPEqCTeAN4m2hbm74pKsP1MXv+C5xpxXsumorUoCGfIF21i3KAltrRuoR34C
BUD57kghOAcx7pkpZZvbD2EIuC5y6FBzzwmcoWadTzn8nI9r6AI24qAKhAkRxHy+lPaNBcEhoXam
SXjRLTzSj1jjcmkJbQgqVyhznRRLoXWC6o83v8Z7LyEQwGuv+3R8gmVgMi2FPsF9ZuJpXGl20KYS
Qwbl6haEPRCwaejEWK6RiM3hluSW4z9nSnH4yVBI3VJCuY/pwj7hzxthjwNgi8VJ/FE6Er9JXkfO
6/dipNintdmpZg0LPeDtIFl8YgR+k/i3yiBfQiDpRJaikdP2l6VQcd7yxrv5N86VjGSbX8JpLnJH
reOCePLix8Yl36V2LP5VcFg0rcM7cM1wNt8W5UAwZ5x2D22+Mj2PvyCb3/uGs5b4vR/iHcnZFP/c
UsSrX46PVyepxCAacbP0Fck8oNZOaja6Pi7kaW8RGaM2Scz78hGLGUJI9vmVtBHlsZbC7h9CGAJC
Re3/01NLEjJoseybqcLffYG7MPSx92AgC5TcuHnoyaSINHHH5k6e6AH79FdXbfDXaMu0nr4QIedt
m7BO2QG9ySdAEU9IlTmAzAAtKBI0WT7wbT7dAn2jqWQru8f6ccsCmR7qV9hHm12Yg9Vbh7x4bbip
R7xRBZwKJYv25rdjdhHgr+lt3DreGjFDXuBjU9goIK04yzAkdY+YRiGmjmG5TthCNXhtTProUi8Z
rq2LNPyp/Pxh04rrwn+Abyf67/2FA0uPZq1UydXcU1xNxbeGEzc5RL5kQHO5CXp0LmGbzNpS2/k6
+Y2eMlqqxahojcF9rjUelhIW5thBsHxvPNQlwJ5QG9TpXI/48LO2k98YuXO9FxQMyOVblEL4NrTp
QEp8k6g3wxFfFHY0McfYzLkBUdlJWXnErF2MQoDmZ/z6famEHY+naC5fZ/bzSAvePgarfTL4LyZT
IvtAf+qHg3Sc/nFK73DbM+i8VVnSSObdFd3cZIiQC6OcVdZpbVQRkHBaDTVZAVWih3eBK1C93nTm
hBTopZPBpua8nz4levyQMay4PBN/Oy95NX3WyQiCjCjMjGAFsWlRiW2jCsU2NcAZ/22pr8WlHb04
/zyKi7ZChQ6d4j2jTz5lyOktMKYQzXvV3ek1Ozkju8N/2VTosMwrqWc7XRrb5VKieU4woXbq+nAD
G4EIbVhqMjuGljhRc04Dq7p1XoC+XFGyJvbMGsFADEqgVb/ZRcV7LMWTk35jJ4m/xt7or+7iK89z
/M9690vudC6KijC4KwiiEgKtFWf0bOyKZlBwKW2wQzyz4WwyIJgJ7qeB3EJd2LSqKP4GSpmdk0e/
z93A3lpQcglNOlNXTZab8BQ45iEEMdWKdt63f5tlhJjb8xmyCNJbLCDPLKcuaE4WHNz3JIpmywYj
ZxuBgYf77ppmI3WJKY1aS1CePOrKn9B9zVPWIq49TeocDy1ZrwKedcF/Et9NJK52EbWCx6lfhpxf
rFAGwMh04u/c/dGHLNyjTS4Ick2xysHiL7zPYI0d0Zy4NXL4S5KxXGGIFrEdV2M4Yc2JaIven1Ai
jDEO6JPXERW/WGbN2xjApieem57NgcxPEP8lyy/GVc4toByNCCHvlq2Hbd5sENOC5WJqz+BuOBtR
MjFS9xj1H0z9PuiVzfNH7cXeg+fgS55izb0WfNkWbQTygkLzfNlr9YnKgOTBVfGGO5f+qgVfKghO
ipHgtYoJAauow/2lYHpV86TDxBt16SBqml/PinKKcXLKTyDLiMvgwMZX2M8Dz8eEnH/5hPmBq6wR
y4KBS887PVdLVPXoqeTpSis99F6gvmF6KeGEkZFPdMaRI52ku1qwZCnBhGvmYsyCLM7cHhJJto61
nIU9dRT7TZDHhOWdMf2IZbGyTOfnGBaLSAK1unwDkKeyfxJDWcRBsOk3ByYYAxvwzncdj9hdH+U6
sSmlarUB9cR3jZuAltPlhVHsLgLTT5sY9cwrS9YtDtX0yraHIGI2Oj1d1Q/MZfF16aAiIps0uGVs
FwnaOKsZBEfyOTXRQ5N5yBLdjcl+Scrp5rPYQZn8BVNYu00gfqYgYWhcH3B1Bxu8RF7ln3SXheuW
8tNIPFO0oBDpsjAcQ4js0+0cP+/Vjr0jZz44mWGTIc8HsgCMiuUcpk2Qzn12QWzrDJQbEhi4RQFB
3WHpTS1LX1Z+RmMVUo5hL8JVxSsgLo5Z81EaFewE6gMDT6iZQrghl0T132V8zEQ5yn7FAHa694ki
MvQ5NJqAU+emBTFwqqNDmgN3DKuP/NDrJgBsDtFkGyGLD7XFDwXhcvgJtgoHJzgmOHlxALRA61AI
nxmNE8BmyKrtxWrF/+SR+vwEIb5bz5FPsiHVJ0eIPnQWsWZdo3uY59mdiWmRllBWdbL4d1IvXTbb
Xr15/t63bw+gMbDPDQYjXdhs9YHqcDN7gM8vt1KCdd5llYoV0zDn8ZCNFm4K3ilZar6/f53/UoRA
GYSXK61q+Y2zuzFg8G5tk29YS0u5y1HgnabyilgFwuFJUuwgd75EkLzT24Wn390RXlEPV8+RlLRO
cDU1Vbz73/SfuDc+RsqlAkiss533NLPVHjH3W6+hs6y+BdydRQVLh3+69LacJQAZwT0soX5Jz3Q7
BCihscKSdNvlYk8J5oAXg3et9CC2tLHuRYCuSyvTgkzd40Midy0rx4lCnasjB50zONjxLrQN8Te4
wtWNB6pxqZFU1+rlM9Ucu0SF4BMO9F8UkJAzT+dnMtr+eewCgGmPls8UhvGVipZYIeS4I5Xk+bg/
jY0qZv5mN5VIUc+49v55rcEzwQ5drASmbeE4ZYNow3vYZWmehj3V10Dr03dIs/8x0uaf/m5fAGzJ
ncA4eVIsBEO7mLKOg6S44wU4n3omzFsVz3OFRi7uxzplNHkSaHgFdNM1mgq7o4JxrvP91Luch72m
+NTXapVnH4DMEHfyfNqTqW4cuJIpMdGMa1Wt4mjJEd/FVkhl2m+OENQm8A+dqgdK9XctXTO1OAvH
T0E6NkRrX2mrsj5e9Ry2BiUcw5r12MGRAUrDvTiUxwTYsICSDaaRI0kSsARdRCNWqdXsyOOfFMLg
LU8rqjzm4tmzvGBcCpiAAsj9MjmADvcgB4T2i8MMDGm3E+cI76I77IXZeBn/QgTRKBsClHuvZghq
r9DHdaFkOKCLZ04IInkcAooLgA+8K2s1wSQGgpweA2zeKKmAUxf2Wkpt4jEJKwjJmHzvXia+d2zX
1+7mx+0hEV3YVkjoMsaFrY90clHFvYFPrOvACZpyJf28/karCU8t0k/aLx3V0k/EXzjxfk2CG9sM
vOgWXh6nubUKhgaHqqtYDJfRR7f3YHlyzknnfc5IArpXSlJ3VzLwWbGqOv5xC7t/g1xGIj/w+Vz1
3qOruBfSJjiihCEn4Zms3fKwFHQlDoUPedbmt2ZeA9i5GwW7HJt1DjK3wL4KiVM1+3OWygYinmYo
kMZUfRo15NthDBNdFiShk2yb/iPiyMgDVrNEpLaCLF0TZ4vJxdaIbsINOVpMjoA8b9c8+vSqVQ1j
jS2RnSjTeBYjNOtgjHXFN6F0EKjK9Y3e5sJTlWo1NSZQW+qZ7Yy8Imk2qxgDltZkvODrIhcPs/Lt
7kXjUSDhXdswOMxX8IOPYphUB0R8BXhkRbmjKB1Fn/qGZ8Ui7BnAkVxrIyKutQbTom1ka2qlmD4N
jY1U7ZUnDIlldsRi47evT86aa9HJKeNgce9Xh7KDAu+3GFGIngVoS/nx9NRTuvL96V+gwyPzA0jX
YjvfFcLe2FFjK8BydScYHE35DK5DOcFYPruJR8owVxoPrLqNHG6hXmmko9Mv4FZdPB0APgh3MTuj
jFZ7PMUKexDWJSqxvM7iTefCBJu/rZbNjfOAHk2yBunqvNMWj4sPMbVa+QDsZFkNsUZSaqLumGmE
PuJZjTZGITHe5kA+Ey1gry0pGJut9XcXUS4b3N8bAiVjJKIHmwQi5R95WObT/pgD1+YS3lBaITFW
jClypJoyWvzRsgqHmdYXhDnDdrA2mvJxaguB1Y0qG4ECLYsICxk6QaL6XXM8uaj5uNUN+BQZDwdf
2MNVk6hnbfqfK0uWeTobui3g41iS58hrXPv9KRsu/NiHF3n2xey0c8LfQxxFqQPsan8RVUPX7GXu
oEUgH8b1wlQBOCoaW1WXW2LVB5WkEhe7W2C60uXuLnsKwaeRRMKteu2cCL58rGQh7Cdb0CL1Q4UL
nHYK1hxAHzDQCrTc3MLuy4N+ogSmWDJ2v749zx8+YlSrMLH0LTvdcK81+W6N936Vx19AzSdBDd/R
SLFWzmxMWia650D6Z4xBUGpQEMdZptlg8yy+I+pBQk0hxNQYZu+cN+XfSNJSrhOnHq0W4csuV9nv
Ky8A47ij/2OCaAeHSJV4cX8cZ0cVt3+8B81lMM1ZNGV6zqjISrHlIVpPDw/POn3AQlZl9PHphnU0
VdQ/l3+N3cJ/ZB9hOYNcN6B1lrFibbULCzpOgfaQGM/RtqnDAgpLo80zs4L3BYQl7AYXbztba+WX
4KlV/8I+8ONWahDYUWOETNxJ2B1sbtD2i3ph3a0vC1LDUsOgH1Yw3HPmEAiHMmc6xUZctWnZHAXz
MZ0AgCU5rUMDB7VOoEqgh2j+T7n2IMm4AZY0NdHp1aTYqGaGbVOM78N0nSJejNWu0Z6qi1Z4yRl7
HN9JEEcv8kWjg5egTgIdVrLzzzRSDfu+nN6PRfOthtSJkWfF4otNmF3DQGwTy5IJqYAOaMpoFnQZ
brhZ11HxYCOPHK001NpHb6Z8/NeNkK1lJSoDdSo8Kdl3SMch4oJMEdsdFvBAR+szezgLyPYlhcHE
TL8fRwpDLrbDlKymBGs5V3WK1L0ewmqAwuOHEd2RHBKE79K1uAMdXPHKkejgWQ6wLHs/Iy/M9Lai
ys0rch5hg056Rc0+lgXfoWgcV5r04DmM7opDPlctSXDnr5MS67IW5wFAYQSBAIvS8/1rigomOe55
E5yvg8amjltikEfyHLQqx25srJQH1zGo479MiibFBH531R5qBkh21LFvCyQn58fh8VgiJDYTyrWG
Ns0PUNksd3aklfIIPOLpai7Oe4uzEI3DxXS2gXhnp4uB1UZCrsLC/rWN29sqHP6Fu5WxyFk7yUWe
7E1R/m9C7QEz1Z7IcydYqN8YUwhlFuLEn+QY8H8s8S/swfymeoXme4s88J6ynmo8JP9zCGqBPnqg
Pa2IuZXxNz8IimtJvArIdbhr3pNXag55ta8ZDY/YQVAb5ecC7v/PlJ5D4HqRVyTbtiAViN7ll/wp
TkTbE1/uH/xwnydbDKNvgVYhojSfFluPH83Bo7bk+s9WBtlvNeZ/E0DoTwKeOJe/CZrlYJMJNhj7
aA9cZOe/JN0Ghdg8CZdGTCNSs8ehCbfJprQNCcXe5hosOF0rUY9gI/n3hE47rv60XH6me2+Aw36s
PA7xg/d5lLWduOZtOdPOY/CLiqWp0x8b8vdkidySQzS67KqZkBBWwBGlOuzD+QNq5kdqPGYppRIJ
44y8YFW0lEAOQVBG0LERJr+XS5DBwariuipaShkJNRGKo6KR/kr15UrvRgX00q0Zo2w8vVRJ7uAG
kzPLwKE0wvuYb5RjWO/bCDLi+WikYp9sMA5zblsahEky/1oWd0Ax8eAzl3+obkSvLQefoIrXyoK5
MUHdJWmhv6eTywEDmvFKW18v5g7TvoDQUIhORz8CETFSiIt2dnnuJmMiirbXZuOg4RBs7auvy7KO
BaPpjpxT2hzXVdWh67/M7rlhZSYxMUOO8gn1uCGWuDCCrNfRpBiybzwoWgruMqbPG4gYMQvvxcWX
/S2cG1BtgWHl02ucyOUA17Ptoc/3uecyypxgzcl5oatJ0CNBuZPyGTof7q0QhyKtiOarDTX83xfP
WmEaNuH2tkKpP0rElCqGAEDi8mbdvxhw3ovBWYfIPUtakPmqhxZWDjk5hI5V/ASDpLBnJxDK/8Wr
3kkw8CFlfxCpV0kLIe8nWfr35x5eyDVj9qewEmEMrAsa3fVCaP/B4qoi2lK4XN4SOTHDWf5Tk1Xk
ZCnl/ANFcVm+USC1Uv1zWMqaZNEv7s/D47rIAR/ZxNnCGSP3aNKsnWWPrFwjp8CU6lLfER+Z6pJd
PCPGIqZTtoKZnE/Dp4cSYzErfRP3W80W2oXRrjJ4MP+MmmtiKJmfGK1A+mj3v0MY9KaJi50jP0vq
xWeUBDniNc/B+YtaRgNa8oAlvmlwEFSrUzFy8CMB+b0iQ/8e2gN3Xvd4wy5N36PGXUv/tPBnOnbi
yw9LhVMIo9zSvKP8R3uCRWDkf41vWNR6nG6Ho8SMy/8L23ngghhRQxgZdfv5/LoPKeA8MHvFrH71
/uifysclZXdXVfuChl60iQsme3XValb7fLC/3Xt6+NuCKCiRA8j7QCyqvUXimVuLw3/sdNPFzFyB
Hf+F8Wp75B/FPq27FOjO8PFfwj9YFLocW7YyLF4pWvomjiqiD5Mr3n9StSfPYQ04dvZJWJRCOzff
hu0dvjaeh3S7c15ghWZFZgfnOdMGDNBqkc0imqh+0+k1bVgVz6CVDd5NuAuWEMZTLTIlciu9Y6mT
xSOnLnsP9rba1OtO+2QM3r0LKCkWsS4b5K3K7h0EFi18D3IPZK1Li01t7ztm7XOp3GHrhgchlTOC
KMt5zMaFlOWFbvvbN1ZZjrz4N0l2+tK4lp9S2orI3gnpr0gQgwYvlNjcSDXcHMtbqyVEayHMFxIs
6tdCcp1LCRL53Gm4hAU4yF+vsb26y42O9QljtugWLi1pprv4C0WgMEDBRX2+YyqMQS0A7wAqpfC+
WvnZEiFjuvny90iw5iaZFxko07QCLX9KGYrRGy173Ddu7AAaDvEa1OhKbJADrleM98V4nn+lNevD
ipxMXJro+UTT2oq6Zk9L1vQfG7o7gdbv5SdtieAqQyjVR2d6bhBKFp3wsPG26bzhrd8sZ+JtkYrU
4ADNETxVgPIRSEzPRjufGhyoVSjic+7UMaFwq8HwKJv0iMYY/BDXAUTeQDcrJ2/Djcf7vUvS2D5a
I55Q4xvpXw/R741su5ylFLZq+lcN/0/qtRMnJPuLKvmGWphL2VouDqSt+OgqKTecfcEjr+ncb25l
8n7CABixbvt2rEurP+97P1m8mq+K2KvNnoyBW/8nDjdgxTiaLC1sLl+djVcPoB65bww0KZwDBUyA
2DGIR8CWVgnhW59maH6z1Kd3F3YZ9WT4RXX6hpRoW7EeWE1aLk5im9Nq40P+WXSRmc1G2uAOmbww
lOi/N6+3SfDIWbE5rOUk57dgwbeSV1wvTV7fnzlQ4TjB7CHK8JeTU4iclZQgRa8gGj+kQhnQYDoL
+cGWBhD3GACbFkY8aHIyGkOVTpadyRi6sfZpkpXu0yN1+kOArFzt4Ko2W0kRFoG04Y1vKWqqfvn9
t9wjoNtjMZqcKpvrYDJnPYCLAXFwkRHToc45IwyXExNkOHxMewjvZ9y07odBXwa0UKG1BMD5vSUc
q7fTD8FsfJ1UTZXFlsguqsq48lfKy5vf7XN/Q9nTotG6DNgfKTzb7f437m59vqW3Ne7FY7nNZW3+
ovFc778+gxPa5pIa+1cbNV81sBNzxtCaCNcveg4t5SW+8gWBOjktcB6PgVdWhGqnhQg1qt+pD+z6
bSH36xXox5eGE7JSzzN0L3jz+ZE9n0TDhKc7fEGvrhzQBeSPq6sAYz23/0JdyZcoSaiAzPZIze33
mpdvLfQugfSKcvU7NHcQiRih8mVHMmt0tYyJ7OoBzP7HjE7e5gq79vT1S+hjKgUIu1Rc6iSRsNM4
EFcHLXb+XQqHSBj1Ohoby0P5V0c20QBUwytzAQv8cRjKq2LgSaYdAJcWaHv4Vs8G4sTZ8tKoSb9Z
LJMwYMPgzitUK3N8K+ZGG3h13IB2erD/YwK+nAl0O2j/pWbgWwMyPIb25nvCKWCJFKDAjI7kgDn5
hSH4biK+BvSxQwsJwO5aT2Hsua6+yE4ijGts0Kx+ReVSzRdioPaZ5PQPa7BRf7ury0k66MV1+Yz6
N9z52jmHllrf5x1G2lSDnV/Pl7lYELiSXvywH9eoYWrxP5/LwfaPRRuUAtv1xAnrONTkOcEM0081
YIsW27o6mbKpajM2bNVdeZiyKGTHUJPYQ6r2xxrrUC1ANbicbjop9ff5m282ejItH06id/9k4Adp
EaozCu9CvFC/jXt1XBKDBrR6Axs0/sZBH4OVW0D0656wicM9peFdxpjYaFYLgZ48HnKDjAyTrnO3
jI2KfYch+V2q+RIFqSD9X94ORqp9GUPVdnmxCGS1EbFuHxct8lLdXJAdCnB1t98SKL6xkhmGnZEA
xCzE5jrcv+czwpJxl6Gveguq1FNgysaE6q1VUKwr5ClD28xE3BhnY1VpBTDe9kJtdqYkPk/0KBqE
oRw3+0sFmvk+rCz2hV7Z0tbz8pIgl4F9cM2Fci6IE40BUn9/uRWmletU8T6LI8m4wSvsJfxBBejH
xdmAgN/o/FHhEMqQKS7HI2QBAfzieoINRquU8J3xAqgMShvMvjJE+FziKDYtNraQD2/op/Z0pXOq
TdLuFM+JL1yJeh9h1Wo57/1TOA8fgA9rLy/r70Un/Ac6u5zjungOQ2D376AlW4+gwrTb1y1jp+Hk
ab9nEtnp7gWJD1r5g3QKpugL5xQW/js46QTQv7D+aFMpMGTUejzfKgxVu4M21nal6V/eJSZUbDC9
2ANnaEYyEEUHQ1PCHkLj+37MyFNDYK99xJLrwyE6ERKjhgMhx3o4uM4ncHV4GfCBBwYxSE4J+aaF
12hnvdfrb0V4zIt9o7w95+aPtK4qlWdrIy5pip3wSXQDikLYAuZfCSYhRInX1pQ4o3f00i/ANP55
oJTvSiez8WQlsGvYo7lX57sz4/E44/hv4fiBj0yu5KJHra8UfqZ6ctjQ2B6jfyguy5WY1yz0B886
glyTT2d/GLP4ZpdneX/fNM0xKrNQZY9Jl0FiwiRt7erAlnX0l8JjSgU9KAueRJsXIqvNLmvrBRP7
QVBIyhrQzWgjViqm0QZUJl3kbSxmVGvL+UlkLJLaRGocm51JlBj8cgOnJqzinBaCFrHNHO1jSf9J
kQlWz7xfdV8kELLscQi0u4SkOfFVlyTvMl2XygOsvhqv7kVVnHAyqnusnK2AAnSVnJf99E6Smxx4
CUi0rbM8nK4qfAuN6uZJ8MFw3FR6SqIB0drNJKeebt3+VZ7uBjU0KjhYR9NQKCQs3OMUHTYZzhT3
SuH+WXL0JBHF7UYAZFkTSbMNrGlSGn0P6pquaJY/EdRRA5qo9G5qrDtOJ9T/yNlb7aMpivjsv/6V
46hv0YehICL59CA0qcYk7gU9ajZ0BKLg0Gayf601Fd9Dop77Kz7+dgKTBMx/Rww3ylmabmnikW8v
RdUcG33DEYsYFSvwWycGg46CnwD9R6VEUj2itdU3i92V3iTEpSGYfBe62fzor11VSAjjHnJ/jBUg
w0hRv/S66m/ke78xYM/9uUZlsgQc3y2cj4RVpI9sRP0HGlJTXMjSnwXeQMrRRbX8ZW4YrY8AWI5N
v5RRrO92dddzJh9p+IaNgqIw/RkXJpoU21pFR7drbzSPhqtb6VBD/HVe+IHcWEf8Uo4FWXXnQSFy
XyuCUuB+Bjd1Ededf7/gY3ohLyjmGop3CCzZ75Zf+ftN4H3AaTZ1A++bsGuGoVrZ5bwKR7OsrEFk
hlH1nxMJXgCtATwSMUYEAp3A+zrRMzzlvJGxYoS8tb4OByRC2wCr3B7xNTVjjFS0pdpmAa50ZArW
FztWvqxSYw3YtNkF2lBuVqPMQYHc94rgY2Qe/wQGPZdwZcpWEVr3gy/VSaPZ9DadK3R1kW22LwOv
NeiPNuIunPaKH4ctW7vR3viJfttIgBCW5D/EQfcrcPmjP+i5hmOoOKOa/KGSq6H1WCj9ekuoz7Ta
JdcoILYDvUBONu0OfgpdkWgEq9HS0XCszx+k2l8Amys2JhIS9IxxjDeBy39mrscpMx+gHn6Lsv/F
/AvrMoNMm3mbXA+6dagdMMvemBiaIQNiB741dy0vtTgWGqdXhRK8TbSX1H+oEI6lc7retejqdfuc
hIsEpRzbLRDTRFPBWKD07G/hKeDyeeyPuENKWZFcP/XCKJka5oFxZqRXhT+PxhlQ3IMav2elwOhk
53sq7J4idlYl3AUaDUym5M0J9EHqHdkY94JdpA2E68HOrzekSgtms0s/GYKpoKh/O9hIhPT2Y48s
n8OKjkx0TFYSmJ6BExYplkqHjYQ6YjFYcJ/lRBe0ille0P+/Eli1Mui6wXWt8IhxCfsm1aokl1bt
x9oB6jmF/hCfbG3DKVy1RNgag7CFREX2i/7Ger+dgnauzmUwYnIuDx332QcldOEVV/frm23WUpEK
BFeArQXD+ojw+Ix1p6GY73ar5eozyTmp0xQQWLYUgnZgb5RkGcRpVCyA/5nYSqHOYcdJf1CGs5ca
/ndc5+PcIePB5hq5HdwmahaSJknv/8ZF4QaMI20tlaZi9AIQSmTAz2zCRr0Ihx9UC8PLK/0O/RgV
J9xrH8u7ukkJUgxVyrcqKiG3yJfOLWPo/I7wG7D7cFNPnNP/GaYD3yP38tzNw9y8zeaEcsocfiOr
bxnBOL0KrxhBRWTj+ba4I0/1LSMRB4FT0ZyQ2oyaPjfpUdrGsK7Ns57LtbVf1rwU9oiTpXJojHv1
LkiLS6AZAiM4qXxLcbV8dbQ2yhhp3H4xzyn9IZK5OmabL7J17FdBH/20UenDe+RrJvIikFL87H08
DKjpvEv7O4FDh76tnb+GKGMv5kdPYs6wFTe4iUi3X5I2sEKI9J9uysS9MLnUB03IgdqiLO2DcmZk
VQ9d8CK3KsdFLTe0tIsphNas3U/44yEj6lzGHbeXPU2XLd9TLkaPE6zHcOU2EnTvLGRSduMo7Ntt
HvLf+OalQORePOp3Donzo09A37LXp3jQQhXWLhfh2YQW27ogJ39K/FIuqkjSm2jznK2RFx3BnQdP
VO0U/F7JTI9Xuyv+KscEDKQ5eJz7wO44Y8l573jS7H6DT0PLB6wd+maHe+l8/nfezKRSege6vIg8
Q+sLsylCej70U7vQuR2fQbjG86FliJ7XeMwgx7VJZotmP0WC1s9Dbbkbk0mtHEQyzlGDWt7r0MnM
WYAMVrlhDHDVG84LhA1mYITFoib31eXdf1vQ0sSR7+nXdjdwRPzlCTqshoVz8PVBSXaflyNCH1xQ
L3jrIAPUKZkiHA8TDRSBQQE+fKpv3aVWfIrxLvLZL74zOD5nC9bEgxvDfj7nlUI/eLxCGk7k9x3N
1JBGZ4f+yBnbbnF0aYWGIPPny3DHtG7/ZGTlRXnTEpzZRT5PI9YVFtyYmNhiGHjlO9vlCMiToBQ/
k9T4EHz3hGGEwzOIRg/DGmwBlGj6VpLrH/jEbPeHP6J7eHDd72Ca2QfZivybBM31C2SbP1GZn1t2
RgUmyRlleV7blrMdxPzmwNoDWbCJncejdvQzsK2kMi8PwPFQnVBIL7tJ467q1ASC9GDJJRzkXsE1
9LzEWMPCNMk4eN9+AaJ5jgxhsNvI9MFVqDqgrkQt1Wh49lM63DqFQILO6YSb/UBIG0L6lT/YotkK
vHyKMNDysZbWWXvz1aQ1MkDqNchD10J9j9wt0J1ogbxeUMI+acq/rPJFbx6wYw4bgIkUbTJC/7vT
Ur4EqDCPDZoew2R6HsBEEpdSVfnNfMuO3TjjlROHooPc9fAFyv4SzD5aLZyQHNM7MwwG4F/lU8ZH
UIUIYKH95NL3/SjuZw3XYSuVVG6oaExxSbGmzvuCwG3jPqQT+feOyRvFz8VbTeNb3ZFflaxwNaoW
+uJm0LpbyrHzuknMRLuJXlNaBUPg+qOmUdW8RL2KqblFuHlcLAHDUe1pVY692wG9D5zataPlfL7b
rEAWOo011yhsS+vdp7GIv9dbQFPrgrSjVKfVZ1+6xSUlEEXTGbQWHhfgQrL0koaF29n3R9lmMNnm
8cbl5vHipt34l/KOZcEe9rTTsSAp5GoY7emgC/8/AQPtHBSNf4l0ggBaEYcEwRzXO5Chc8yw30pe
WnNZEaV9oYFcbHuGWscU4UinX6ytDV1CLsrRHD+IR977wsVLSBo+4T804lcaoObGYB0EUvr4Oc39
IOyjgx7Wr0r+0ZR9NJbPlbmqRIz7ImPA8HxDbq8R7LBs/x2pacJGcY1CEMGSuF6ef7VANKHjNfU/
nT74kKTkxXB8p2HZ+8/9WBLTfZxjfNUOROcgGozbO3Kmy+CkJzcT7fcZYBBgZuZVdnWHgs78JczR
l0UwKviE4//Mz7okkgA1xGCRmjRzrRrwMdsctqEPuOcqpAHGkLWfeNneIQEJoI28+j8f8zYEKytj
QM7GBmHuR2Q97AJaZeAH8qYIAWsmFnBDR5++brjJwf4VdMERXxgRISzdCe1wxsB0mam3gKThyoff
NGt/jMOUuODhZIkH5Gkl4U3V8a332eNYBDWIK5oR21EWoFyNeiXjlqmGf2/EbGMc7PtSknahRP3d
upnzlzysXwMmf2VqDpTKmEnTaKaBHU2uFfOZVY1DhgFRRnwunf8xyVo9cUo+JEzx7NIVcgSBgZjQ
VxnjLz0y47UewhWB64gvkCFtEQh7hd464rAzshP2GFNp5WSHuOu8b3rFg47L6GItHXN82dpOc7am
6FxZjGQd6vYEUlfUPZI+bvUIUUYKqFNvBGfnJWMKNDxTSN4f/YGyRkyQIuNH9E7a8h2lulmutb8p
cMlhg475PZn8Ig5cECS0Xf0jW4GDKbI5FNDS1KusmtAs6ZsUfQl/TePlGuc5IT7/vjmFBhnubXD+
RNhVhDkbh2kwK3xAqN9lyf/q2gWX/LuV6KpQlJPCyP/V3WRb2xGEPu4rIIAZghaNWAZFOHIlc1q4
aQ1plNGKkOqAA/ssCYAm3A6XkhZO1Oxv6cAkBLpiW3TYErR/dBK+k4d5cH8xmmgqgn8VxzINJNuX
f10SreynGldlbPyPi4P+vK2u+6sbbHKMV3+2DZ6WlE4bGSvk+RI/+EESW95buwKWPuc2VPLU9oj9
jML9lE/mBlcWWSFZHKWP/CsCj8lle2bXrz2EodlmgN0xi5VfqnSe2QRnC6tmGvxxRqONRP6RirE3
CtPOL6DvLjL2BD/FEbiWQVFZu8FloUzdz53NaB4l2pfLnb6o7GOcDQGL8OGyfOED5NeLeOzKQrq9
OR9MEarSPMJGoL8tU2xMCU9paFregPVyKH2KhU590xzWqtsI/R65inyivjIS51EwDAPVZSVKMZAG
6zceBy+zAF5JF2N1AL+kAoNmnzlyQFLDABXl4Z1CyUno5VORLjsmqAN6JvUcTHD0C2L6F52pEiJ4
1G/TWJJCjcjIyGxUNETteGhIheDScRu+CCkoUrj9Ehgk084IzHRG8sC90IXAMJTT5C6uM94hCeBG
I0bUVUd7pscHK7iB4KwBwEQ5bc1ml8nqnAVYIDA1ftR6sY/WeCWBfQVw0NPWLvnSQXjlbC0SM/0K
Z3IxuZHNxZFAkh/DanTJEiJq/31B++IzQXRtZ86MYLa/+BbPXW43Qk0fJCvMQ8gh4ZVoPoh8CtXG
D4eBYRXvRA7tBq/9ognhb7RGnqJNGmDQll7xBylDQPhwC0qNifOWgmZWW8Cw/KCRTLx2sIepg2d+
Qgxu7cDEtAUxNVVecSVOI4Q0aZQJIYx+BaMkwb7vZ7PLDACOeP2zZhKLNSlTgKEBgmGr8Q7bOVVJ
wWkHRGwAFCDujATKY9UdbTklfNHY0BXkaV3wgQjrLeSd5G2RV7d73NQq2FNGgM8/i1bDmoOKRBRJ
V97RUbvfPglHTkm3Gqcjr4bJoWM1q1zEAV3ixtY3jVCG1rdhV9nwgKsOgfOcZVL0gHBIfnT8RjxX
cbLQxH7EA3sVEHRrs5MUqLczLAd+lZdQmdadzjLLMnmEVoyZg7sBleH42YUp1icDhHr/QiFJiTc6
s5GNYKoCjxaKCtVjW9JKrSVuI3VF5Ga1XJOcDme7Xn3/66wDmqPYJzhBC0R/OnH/L6cpCl1vdIB9
wAKXSD6Ii2mSb9LnrcWoxLghqdTtdDoi5B5ZrZPf2qEsQXXfPAhi2kOJ/dPxxm9qhG7QyRA4N97z
5IYgaMdrYQvmE1XuTeBhcwdYtjOgY2BQzHdTVNFnApnF7LaYexYXvdfd+GeX5mt5ZfJih/1yQP22
tSwuD3406JR+od5OmhSzb7yR5t1uWHLk2qO7ANRh/OUGTve8QlpdvY0SUsBSCEr5SS/7SbmCIGmF
aAEzlhEy2ts1ovYhAvyvonfeYqxFSS8xvFgS97MzyMs0/DDdL6ozxPDao7g8M86hsnI9ltgg/qoY
Bq0SG/fsyUpLHqiB2stLAs8L+UR/Nlpll7PQlQd8lsQw24/H6PNr3CChCXlf2DDYczcGvB/X+83Y
1w2hrXtXFdol3uGMjGL1E9Dk+8J10PjelgigABoMq5Y9ni/pusizL6KdCkA9YNuHWKGR+u5P2BXn
Byzv52piQVqpqt6d3KLWaXBJRkB3sXLgg/NCF18vtOusZRvsI0C/f8Xel5iYDh+SEnVdf0TJkQ6E
uBI+pWThNLFqoW9nd1wLFgn68T4eOMwYhEnY+/NTzwFwqCXfbzDVvYZ6iFuLbgiRywgG5rrcjDNq
BYqHq1yl9LLZpOpnKhuYdYrgTAYjYKmZ2EqRdSoucjetJrLx8k+j4H01dHkjoRpbHdOnVaZsbG82
qr/kVr1GXQ2YDi5jzIkUV/Hv1hXO1BxNPqT1S6VpQDJ9bpOo347Tmp+XOtfcMo88s1f/zna7nSox
NIZ+Jfq1+QXM39VtRqK88omi6CRwDFaNzdfusOdyTrDXU8fl3bDxED01jAuCtkudzrEEKEY74ZhU
nK3X3E3+y0r5V4OQ2P7qXnKNSgPsIQduZb8aGN9iEzODPqKKcxkuX/a3D3HfGHT1tL+qMAgCxpET
6GEodDqmT6Rfj6ED9Mhk5b3R38KmwTg4oobfmCzexL3n3imGa7zsMrZx769Nl4iszjVXvbQDHbKL
ZErvToRtFiXYdNClgqnK7NURmNiS8ITMsCcS4oAyAnQW1MADxVIQOWrCxMFiK9WGfzoCVcl+MNwg
cix5XtXgwRPjIHL3fsojIp8k/igISA6lsffYePRsW4fat6sQ6xEKqZjQSUegdiIOhJVkEOikt0qJ
11TvIHUd/jkqkvef3Aad2VFKZRSsYQ4AxK2N5IAWCRlKl0Dj1tzqloxwC5CU1Qcao9L2e+CUaHYk
I5PtDAmVB46jz/8FSavBCaJMeTeTwzS+25EYJQ+nN82IkLfrVYAT+M9pKjYdsBuv9bnBoQPZCMr5
Ni6eqXbSZU+AbIp2fpQFnTRpx5Bax88x1P1vhJopoEpAWhrO/uNmg5LvJiFOmhQgbanI2I3I4UNU
4tIfGlEW7AQhuvh+UXndKf+t4AOs8k7tLOS2RMLIK/NbxVZIlHyL1h8nzsGtitrkyCo4yRV1Mjtw
b/yZc5rQzMnJUvRSWLTTlfa14gWDojrEZ0PBBLNgtX4qGTATGsvC+4T4p8GYS809VViGqYWGUQjK
761oOpIsTYIawuIWPqXwGpEkVdMiW+VRdj1KQ7ni15WQvw1QYD97k4AZnxU2ywwgi6ZegI2kP0gx
mZZZgQjEy0XwRJNr61trSNs4c8TuDIwKzq5pwtfotYzUBW8ycbzFH567Rt93fWnxI6MAkuX0pEVN
/qGWFCxHsbLQy9seybOxZsQ5TC+Q8Db7myB1rUvQ0nLhP3zWbn0s1mrqxan0d/DvpLOOecjxur1t
lOO8LuzO0qLGiiZzwVlMaCluviDd5D66cGIzdwBhDq7/pXpMTNn1XmJ7W0i06AuJ+X2tdRkrX3UO
2+THZgsBy3gyybR+mxLzEhEcYWuyX2rNFjquQEeaPEa2aYRIPi5eUt35EgirfCCycLawXOxEnzrr
e5bD0Ag6xPqd1JBMoil1oMNd7bazznAOhyNJMA3ouvmy4L/Q6PP3naeHh3ks58XvgBp6ccorknIS
XatOXg3hEl6TPsbXfvSJ4epwJrGlMxEakVxXzvJaTSQLG2MhWwnER6UWcZz8Ioa2aFYuw4kETIbQ
9nM/kP7/NnnSzn32DmttuyGGK5yjDCfIRct6AslMGUzVe+l35DJWceT6ESESUPZoUm8uT7aKXe7w
WYnmvXCyc3YqWNnH9pPt/avFYiHzPAs5Kb2rbkV7mfG4F4HnSuvXUiXdvfPp8JFz2i1Jm2cfhoKh
CgtnHzB8yldc5b7nCBvPQo0WvYwC5nEN6vKNZSkEyFfiSUOeRpRygee+xHmdo7pffWmjnM3dStEX
e6Qe4UcN3U+v0r0XIjM7gVladlkEDKo6yMj14DWvHZms55l34d5wDfYbEeNjS112r1wn9F8EFG6T
4B/ObweVYjiZYhFZHPR2gWZ+anW8DJkR6C9JAI+UCBcdcgR/MNvBtqRkOQZIu1nUsDdykxCizKx1
vGgKLiAbow6Qwf69d+65m+lVjA+zOv+fq5OYHgjmIUHzqPW1gG/e1XvOmP62uL10Ax8DpOM8GHc4
uj/5ij49XIg8XRLnfHm6RIITzFGgZHjp/Y7ArfZ+u762JcLrx1TjEJZUpjzB2Gsc75QdC1f1y1rw
yF9NIKpjyXeuasbTx0bo/lzgxgGPNpoe/3ruasFBctggiQ6ResXRNs7GmM+bvO9l5RKHj0nKsLpp
znJE3AAY1cme0TdePWqsPinlEfmOFNuffd/B1fhvvXMsqn64hzuQXHGstwVEcjoHaU2r1oR08VYx
Fy4647fdiYWTKk1bSq9X8POoKANmA8KZEdKIRLzw1u7U902QJUGpnLbCKYJSSQ/8GPNKQk60Q7rq
Bx2tb6/BpF1yRtgFfKpihd2EAKj5qLRp+/XuiIl4vgTkOhuXASfnRu+SXrPXVYCIkorwR7COjUW0
bF0YDNF91SD1Rmuis+A4Vj00rlt73qMlju+cRhSwY8LTl5WSZ10prxRawo5DSZSles4DperdBuyb
usZ6lnLRy4aJ1iwbiqFrg1m7/4tDfJH0lTmK5zfYP9M7Lcg4FQb70UMb+wA0/JZyNaUkqcNAB0lf
UJD+ynR/tZw7/rvtK1yw2i+l8eJQQ94sccBWVXCEoveL4+dAWxvxoSzDpF7kjlfCENjdAfxO/+Am
Vml2Oeqr2vcUekN2rhijXy+7EKRFAYNVQbLN0aZ7gm/dlS5lThIKStENhsv1KTb4JtcXJoygZYv9
iVIHbfTgjiTHkLUok6ifq14Zw0hibSQRD296AjU+kdUFIAr2678L0Em1trLSQ0Gg3Ltoa9sp4Y6W
dOuPibbDlu2A40rYVgbdufpyK4OORVsBFHfIM6Q9G5cPHYLkU6mHl8nSXCE6brFMkXolSxDaAEhy
xS0TLe3Wg+tYHxrDvAXXMuKzRxYmtXL9BDsqExRrTlSXQUOKFLr2wgnMigvUCG2UBwrL9HP2Issf
nuN3DdSA0jxOddNRtJwNoxv6GpRbYWyMo37b948pDC8N/0pIT74ndCSTp1xCy3OyaTjdI5auLyWv
D4KCzYkOUo8P49amctcFnE1TlxbEibQOQgmVlddpG++f1zx2o90fAe5RhhPKFPYy1T2ojQqybCsY
S+bZISIDHxMKmgRK6cvtGJoHNleVfGhXsF+iaQI9WnJXoRy6gm9G713E8GSjKk+Fokm8187qPaKp
LrvPJvXI6WwZ5x5jD7sC4b6s3dbU/MJ7e+/OaxN/JJOotDlimlFf++DC3lTzYTKkoVeLihytVq7o
lI48FkM91A0TYlCSlcQcXjtiGjxJjTg8a8Zwt2w3DFaXl4WdQVfgTDU4lJopeFaSpG0d/zB1G7np
3sXHNjsbuQx2g5ByaQwLX6t5+MfJuiEfwjaID8R/koG+1toe0qLaIuyLJlxCcsztGFlymoYoULd8
bTUkUjXiSCELyJ7AHom8F9MXABoqRAo3T2ozGHmpOrXTGuV9//RTJzvGbYakU1SGtMAb1MUQvcl1
fR4nyspX7GFKNvYrQRu4KI/GcDxvHVM4g5oEYb7cNDjad8xEPPxY99ILE1n5du/k6BNgYkCNcD0e
OenA0jGF9lac80aD2gAD9gBZzsMiSJG8BU6sk3lven3U2ONn4KS+MBSRSAbKVFDjCX5xmLxSWgNf
zkZbZNqZBCOhDaC/pey8EuCFOg1Gc9nzTgE1+rq2Rv1Ww4mHHm9F0tKbTCulmG2LxeSMQ9ajnKWk
47mK3f0EKsKPw+svjMnK7Qbn3ss8Dzw2XFYJXECBIIqv+OBswWJeaVXuPHB3tig63cV5/vWc57Rz
CE0rEg7Q4Bl/nRcjBvPsBZdfFtB5qOOpQuwcNGDfNAmAufkI43L2/kJfQtOvZ9M1suMpmQNJ7KtL
s+1zmwnv5O2mB77wYC0VUa3PUw2yZVCVoYwYyy50OTUXyQbxEXRiB6NNb5KDSYPXxYZe2VoU69+W
yP4KqDtg33KgVrcyF7K2Pc6WoEPMbNEtlsDKwcyvrb2pLM4d2xSNTxdL74zLmpJt2CRZSgURmVgU
jdvdeEuaRrxWwoJEO0lvO7Q7sR3bYlz3V9nWuDsjq2bZp72Z5IiN3NVRT7EG4bQtnEKVSOP/gBea
Bk2FAvaYj1fyBu8QwbeHE5xYE1rC5lzyl/5xXXJZwRdRSwqKV1DkOTtMkXEiZh2P+MU0/T66gcjE
xwf+s6qpe1hBjdhBuyQwGPonAVsLQqlPJNuLFaYNXv5C6zZb3KbmpH/9KUBDJkH6VOtd9ZFWpar6
eCuVF63kSqDruvMg+s0sFhpqUKo14xn9Iih/0f95E61rZL9xEUHAjYtdT/CDirllKlu0egjHS2O/
MfFAPhU3AA1NPRx+zgdK+WP0Mb0jobsr7iA1yTpBqrHTKknv6am1FP2t/X1/u/yiMM1h5Y/5W/mQ
Huc+l9BPKne22NjkgArp5tYqUf34waKzOlH2+DEmVqR2fRd+L6xKf1xZowuUoA2HZlw7Gj5ql/cF
GlKxTyY5yVG3/ONoJEssQvgctiUryYSNviAApXmREpMGNeSIC2RDmwo0eGAh3cEk3igPD8tHhye7
THq4bRM0SLuW5MC7d4br2bRcxM/5lBLtc9VK20HPS2PqSpKkb9b5sF+YM1869Rfgn+vJM6Te/64s
ThbBjXNazH3+ZKQbHqv/1ZNNmoBkY5mWojZ5c9iEY1By8rA9FubvekneboA0zlJeGXiBpHcN5Wkl
wtUXctfBofbPkVezmVV0/gXdSD3MMLkT1X8f9p8bAM9htHJ0S0ygUgf56kGw4JtpXSoU03HBIf02
tz6sIRx1mJ4tONYpdCBAwx3EsXAEAEkB/Hn0jfUhrY2npvFWPnO1gTNrbv3gudITDjXrX4TKbZ7Z
S/3si7PISQhOCm2uSlmXGLd2eOFwtY9fVtqm2hehB5tLpe18TAlwrw5PMl3q9Qf5D0DXjkADc3Dt
FQlU0yzoMysRb6YW2XzZDSnup3EopenUn8O0zlPj4jFyYPaA1ooV2XaXyNC+Mf7l1jZ4n+55lHaM
TF+xoG25kytf5N2PUqrd8STRw6Xyx5q72vj4gWh1IEfncIhGTyLBdg01haZ5xkBPagrbTL7KKMht
L+k52x5qcqUHlY1vto4cKqhEAGov/456E3HGuXlNvHP1n/1U9qTfG2flcrUey1A9XOpT21H8VPxe
GKMtxTicz1xfLVNq0Z4JEOAs9JdvDmO8X+IOejbzyxlUJXLNpPGykiTFMHVCpEb6XtwbLM/uetIB
bEvsPQGT6KFn0nSMa4Ep2Rj0iQuuO+lZc48INfn8ATjBI64PKMpLQP3y9csJO8Eamw2wBqUy+SCO
x3PiZ/FfnbaYJ20kQhhDwk+5nc7DiDbJGTTH3DdCXYXbmvdyuk3jhTCKM7+24AuhJ5NOCxB1AQh9
wSROhOKMCqKE6ScD3keAc0ID8hXZ0cHpBvriK76phaA8qoms28KnzX2yaJq74xI11FoX8nyv5N4d
JZ4OQkR1fO8pmh0k0EW9eRcQdnXftDcIA2SCgA7MUV4PHyNRSY/5eDO3EAs+JpFBSz27HLLMbFmF
qBprk6alkAYUtcD3VGCzFqhF4cDX1j0xQR9R+A+PIyD3P3UdYyunFxb+frldeJ4TktjX2AvrHqz6
uVXr7omMsUecK5GCrKHJLwLRG3nnAQIs1EHnHQay5YSZdw6qkrjVNgvIj2GPQxJUZAOOy/ITSWAL
Ru515gQ9WR5Yi3l/ZDlfpDhYeqK+Be4DItdb8DCfPUjAjcMDEPhx1o6DccWRI/XKjXrea/q9MS5F
4xf3c5w4dRD4mN1N6F8lvhFscL91Iwa8iXMmGEj06xnJde4fTRuuwzJb+Z6+G5l2TRxCj6AvBrh6
PqG1C64kj5aT+ilypbjxxr2u7plJHUXy7y4p+PkKhunYnx5V06VpDmC8OO2qVvwEoHQq31lkCe11
jykmrwZzLn8B2uvFrOUzIVjp6k6PqhZ5btuU2ctRbZNtauGcEi11HhB/RNgB0o1ShFlASeSN1N+c
mipzdtDHwAegLCUnVCkiLAJFjOr7zSi0x58Mw7oYoCxn0XHvgFzsDj0R6vKm1US32eX/7tKPwZU+
OZ3uigccx2uAzZqwrbAJ/x1YI+gq8JIwefbDU4KfubrJ2hXZpRFtXVmorRce7o7m9phxi6GgKIAw
+M0CiHNyHHlIt+Sy1d3d3jBTXAYMQJT9tPLXD3ensN5z4ofyM5+fR/gtVGEawoKKeVmnuDSzajbG
YFKRXXsQGA1UYIc9i0FcbANPDbUnBehOTly00Oub7wI8np2UyxIeZRsnDXf1s57XuPgLPDhVlND/
lkp2/C7ShqMsVPYx+rzUnLlD3WinpxNx8MsCr9MBxcURfrfpahpLxSoi0YRk23DFN0AbrMtrT7MK
hx0qlhzYlcRSYi4YGCSLjrqzhe7ixUGiiqDrda20IeQGPUK5f2w5fQyTlSdjDZ3zuRnljJ2feprX
dCekrtAtISqH7g5AD3LyLw1sweXjD52JhjxM9+B2I8+TYQDccLFeZe6j7k4IdwczcGaLpkKbP439
nhFk6BgcF66LhVjFZFMDcH10YhigxXD2JgmcZrAF2Jgdfsu3R4kC58W97WW0+Dc5wCwF5Hg/guMv
tvC78xpXUZuTOvHUiB99VakNwdJHldAXEUuRQVx2CczCsVZq1Wo1w+cNBfa8ZtbtBMamV3gR0Z1m
rzs6+82JEPijTrx0daCfAejhx1edkQ7xyKtMOiGtQVkVg3qK07DRu0x2nIYmQboeyL4LM/l8jooD
0qdR/hsN2OvuJSWm271rdrxGQHm35J9GzSUaHooC7OBoonNFDT7NPqhoZsjNDy1a0nN8130ECk1w
UA5aM2gwvPwiSjO5SXooZonZFNA1LpOT4Mh/Rh1UsP07pTj7e0ofPhLIEyGJGTlGfpRnFvPwAVGK
XOOUoWAfdn7posV54EPPJQ564mSYsPAN2BzaSARY3blJXhUxDXkIji6Q8Gxx1wAd1SgpeOQTSBut
MffL8V2zxx78KgFDQ8NdsSa4yScCt23XYfbcGrNMHuZtL+hfUhXMvS5xSHOvd1lcQbLwXdxCFRGQ
+EscmBWTHpabyrHWgBwkXgKuQNz3YoNQG3vPm7ONKkeoYBcGRWyMTznmw/pWaPgdIcAdh7dkX/z7
MAnUvUCYgr4S3/w6wLs0WQtk5wkgy9Vg7Ezq/+8dtpe6yTIdct6RFF/536Q6C0kbPJ6yrhQ1x6Qp
VLzmCj27VWqmXxHtYM+eGZpbvR2x3nqJkufmVhALWNfbTdRDORucYgyf7kdteUf7fnRHWUMjBuIA
V/G+diA64gqUVDXMtjE2Dle1DVmODjcNNv3xQGKTjPOs6oL+V/PmAoNX3BOlIoMAWWQcLAWwsrR2
KiQkaGF12xa4RfCbHmRJ4Gw/xAbQXpNXVj03eRzjDMcFm+BQ6r6PZbvWpfFcH3FcUsq8UyHl1+jG
C3bxbilkdsSbJ7IE6i0oVwRyAlIrlkOrVXZmBPZXlcuVAxhHx+34aO5Ql3JaRM7w8v6SnTXUjkd7
XfpV1gc3yeLna6kHgBzZUP0fi1Az3Wnx+vc8M7ICBHw4bvEbzjhvelgqWvJSVm8QwY0DCV+/2GXy
+mKN7HTMJkyuNfks9b6Y4GMEJptIOUzL4a789v3prnx5LGavfOf9we+T/iWkdwJPy2BzQ4XSS9zb
7hfJfzX7ISUNu7pc/RoYpypiS5Yjg9ZMnPQhcHaao7hEyawz8GBAcUpXkRNa5o+dJ+tz4cVniRVy
jt2dkTmpPUcgHL0IqhBb7oHQz5LdPEqJaj6hQ2ONWOy4M5n6C3rQ/N+oIn3vYZDlSEH8h/kcYmwg
IgMMOOqyXb7SNPNxpkTgL7LQN3UuiPyjixMZV0QfCafgtdMCeDi3TlL8sBHeuDLmjDNLrD9KES4Y
b3urgkNsYIQXRozQXo5t3QwdYDwVTBsqK+GOwQ27YWYpp0KxMQAipM9QgTDDfDpETEuALcN1ww6M
eCw+A8TRoiaXqr2jzPmKfkyi5JCDFlQMJcO1ZrDSXWP2PQsWzxvgW7K3h3eXJfqxBjkMgdW9nW1c
fx4xp/NmmWIx63Go/NpMbsOylIuKB5TiOrHuRRO8tWogOnR2YqyHRUK9g93en5+n7RsU+wDAbrVS
mzgW+hbL8ZMriqFIf6lzP5wELlmkcyBCoLZFupB22TUHsme+kZW76bBNdbSEqe2KztFe2qxWVITv
v7g8u23MZUh/M59SwwUrWzsyCysX24hs5XBMBjjtEQwFVsLkoqCDKvyrHdo/uE4/gmav90M0uRPr
0WT96OoySZoZJzKxYG2cSiy7J75FXF21pa72a2w/B6e7S/pAnfoKUZfoK3mS0MxGQlbqtEFcVmJQ
DAtH58kj8w7LMZ6CUR/x0+Q39A1WsSWtUM7YeQq8adf6ZgXemz7r59YisWkmXSYP6tm7aZkWigty
n9sWVXKoFUOysii38NdRAgO/gE8ub0XwNw1uBMUzZhPZglgEV8LSSQoKXkW8vKEqpBrSN5Xwa8Mp
YAtDHLwY27yiS4gFSdGiYXfDeQbP6isq8bcPqJ1zCTl/un6nBTbM6FPSbZUHJhcaLeCMDbLjHWfF
tk9gDMr+3wUyVoqr+hrY2mOA0/A/QBPybynOTgjjoHIy38NIFLgwm/kBz5ZBEJz4qupoe7Y9K+RC
1ph16BmYUkg0TqFmWgvRIdOGcjchY3e/7JmXZjVI3tt9IsuwNK+w8XgM1fj4P6LAatk7weON8pxC
8nCZzuVFTWrW/gHORpg2stNPr/6zAdgiO9/IdU+bMyai7n+1KfqCDEocWUfaVYLZDSm9GmM67Sjv
eK8pGCd5eUVnHp5zVrtJdL3nInydwFwk59BhtXhgDHmlXlynP2nPfue7DttWqZsnGuoRNrLhPdMv
wHBykZ5RVbtybW3xVMlOVa2ppY+HLreaQu6wNi2tXVUairHkhf8mVbhu/cZY55aZleQx7Bas/+Pu
hAVC9U07cv4CJ5/BwwanTxCHvSTMzEgIaF+V1W9V97d9zBK8KlmaKwebvD9iBxeDleHpMsJ9t46n
ZqITMLUw2MMasD2QFvUFE0l5tjJjKE60HsFycXBU/FuRwQNOpXi9d8zwifkpnhmWYzKlarljyyJw
hsFf26YnEqL/JhR7tuHMUk0bvU1pHtMNMX0wLtJYFyoSEQjhBeUgQIX2ktnLXG3x8GYPVwdqDfRD
Of+JzqyoZqOLL8lwIvIif4f5pdAwTlk7OsvKK0/Sj1kpcRlgP/bX+gjH9t17C32RV8Jd1rkIu7pZ
0eghmIO9GgwC7qvJYMsGFknNK/RpR/l+BKGV34jSV1TB5r653MNAdaku1i0c10NXsz7TECv3+VKk
8YqUcrMsR1PVZtbWJ2tBD765qNjuQuQuseN8jXLrIt/JtlawQPsK1vrk3ALCxCmWaiqJOyIc3sS9
wdhQ13bFK+XEtFqSC9fC8LkBCkyB9Ihxg4PBfAGKVsWGM3bKSAlXVcPkbARwUHbCtexKQe05nSec
WlVGBBKl7mhWVyi6DM3FgULB2V6TQOjZdTbLAjI/ayoKZhAT2wvmfghdIaU0i/2ezHwwzNvEZQXL
UrtSHft01kq9YloOO/5dRvQJfmOzK2h92VkwHNAsANpiGH6Z1A4yQf6JVFljcM1XffCWOQD+qOER
lA6UD/z9SPajaGlsc5oS32PKdG/3NK98vqdzL2rTAuSfCps5Y3zMkfxtO9fzOHkmuU12psociG8n
jPlsb1VxDeMO9LNSorw68C1LDqqkMvk2KMz7Vk9oViudFlS8JtwTkk57BRRO+uknqot0wDYPq5Ff
n3LDucMQBcYtGk1PX9g92ZMLUQ0uFupStC+LO6VmZcmsxxhQXQe5PhGJOagECj1LHWGdOK1VBUck
z8ThpbOr3SnzPBGBBLwpWj67w9LxAh2Eeyfvzq/aMFD97Fp5rykRskAi5wpFO9Y3idOMvMbyE0W2
P8u5VXIzh7Flme0nkW42boNkl1pzHrG6ZhC9MWcZj2VTVSrjhXTSMu22WJaMdZLY3T0TZqjq4aJH
/2zT3jqX+mpri2x6Ahtq1AWduuYVop/SFEs4jWI6IvoFCOSfWpbYhsFyP9Vp2NtPqoj0dMdjTTzP
sjW4rMFY+HSxKunD4a8PQc41BdRTCFex/9FyaYI1lJK0rvM1YD4tMRtvyaI6cqokFJlXE7Vpi/dt
aM5DWI6rpglTVQpV9LVm/XlX69u50sf/oqu/B/LhJ2mPzGrEinV3DpIZuDWPzB1B68JL5TfhwAgV
tXNp080Ovc/FsxrCjBmcpqqyff3s1WXthXnzrpqIdgQY3rbI7L+r9zE4HFug52Zmd3rHLAXpz07G
WMaBzHENjgoZpL9QMBS00PLOUSOTDKf7J1FuMZOlR6zAr05T84FzPsMks+5Y//gjJb0xvAZunF3k
Dg6W4QWJI1vx789IOPlOmobfDrG/OjXrVSW839DfBkOMMnvK/kY07PFXO2fmwSMl4XGMC5wORhgR
xNIJfGoqJ2Gx0NeopVYocR7ykoHEyRnjBTmF8rs4NdfkVBMSS126BMpwMmy53mkU8iuIQD5oUmbe
HabEA6z80RjsQqAsMWUbKJHzrZj7u1dr6v4cQqjwJY2omY2hjkBgI0GnMTZiPkMCswbJsDxrNZ5y
DakaugEkYLTXVA3LE/ZuX8nToqNyDiO/BU1byRi1txeiaOCXd5eU0SZKxfhLQd6P2wKeQv2K7ZOz
TDUdRp/GammEyvA6ONpUrdpv5MxQCeQzm/6Yu59OUHAqYs2zyDhRNtHokt4gNKImqFqXkoxVSV81
EF6SwDJabucSxGYcPmxHS9WP/GoQNhMsihqjL1E+NdunwpKFrwZemrZ8k6TU98Gxw0FwkYtUD1Ig
BJdFeekC7cImQgJJJ2emFlV9GxSxVYIJUT74y0h962sTaQR2BkX8jUiaelqzNhou5HxZOi++jPzg
yJJZmkgD9WbQw1GVgzUoFT8UzprSuv7YgUePOXA2LEJxm5M2VT56Bw77g9nfLlBVu/u7OFIFH9qX
58JsbpA5SiUuURcc1Mpix/BXMepy4IRdFAu2288XWmyn0gundYVJOqV+0K6cog2h77LJYC+XjtYf
lZjsByeJRdnhfrmKRElJOxYd7jqQ9R1fwera5rxfMMyoYFpSau4joam7sKfSUr642MMwxORkUnLO
m9qV6KxicIjTA76uKiyhehbd9dGnm/0HJvmPAXFNciTB8TJ8eLw8Zcvj67bX0s/uML8UYmn4u0Cs
I7qdHfZ3c8Ksak9Rh1oGaRTvvhgKqoOGO6FuI9vz9ppAUA+l8DleSbf0rQznmtHVitRkXxs+BjiU
ejAJtGz1NYSAAXBRsi+Pk9kdVgkb96/0hpA7Rpyhw3X30iIRpoMtSPz31K2x1H5LBRBrpH51WJX1
t49adTHGBP9tItrSJiKiulJSB4ZuBVT/pvJwbmO7kWiiRtZiUQ3b1JZn875UhmNqyfwnOlfFTFXF
e1kW9wcge8MfH60f8/KpKMgS3h34RNCZsyi+hjYzvPDFwUqaqrkntNbt7LlcLjc9+AyKm/XHSt2R
an9YEjTBgFLTRuCde6NQYx8nVTaR42gjSXVuMut9f4RqtGVhHTfS7yNADLrZ0mdkJsGY79Mj2z7D
fuqc1xbkZEGGKhv7CCeGJ0Bs0d81owb+6vqiFqO1mQDioCKwjOrpV8lnmaMmJvtkZrp3kOQVian2
JHlyikWMgMrkBRTT8qMt7n3earwlRdVUDukjTbG3TrToK8B+mfewpX8K1ejFPRBC147r806XEP7s
J5CDDMNE+lK5xwNuroZ2GDve/YkAtaZI8MtQf8Xkl9XsYEyVqDEqkZ3EKX1NNDGxxIFBDJxJmP0A
NuIZ6wEIiKNrgq0eMMUO6kantfXlMqCLrSJm/TfkEU0uLw0F/NkTl4lr/LWE+NUhIvit1vy/7109
qJFIcRCi6R1A/vz66b/iJAljUaTdJl87j/6Raav9ssGo+ey5Q+a8m4rh5A5CwuV2vPH0cyblbHNy
R6kEDHpdKTcjbyABeLEyPHg7sLF1/8R42hX3pwxuTpmh5gvtp3Q+xrHXZpIPJZD+/dwglIobhoNi
aFPKR7lrlOnTiiL3l3k6wr7vQ2T2wGineHPiedNbrPhZ+OK7EX5+d96efQ854B7wu659UYGe1XX9
1wcmRZBjJjSBFrjr76byYMEbPSeM4HpfHwM6PMbRKqT65DNv2SIx7M2iz2rBd4JSFSMl09hv7Nmf
VkFvqj2F2CF4pO9gxX1Qa4pmpfXtxqQRE+SV8XP+f33p4LiiHfxu2P96Tf7+2ii92fkNfP5C0lmm
ig9Ox6UchqgGVc8dhLURz183l36cG7VTXErslnRXw98DZL6j4qSCEZ8r6Khh3xY8kTZG4i8QYALu
bvCSoZaVTreQkPi/pP5o0V7DHjWOghouyJ47faSvyZDRDf/KNtB2jXuNO9GVAuuGnI3fO7vEmJQe
AC/RHfCKdwsnJEQiesSSsIwIDC/MsE3JsKIyYMIDW+AK2tjCUWatEGvyRMDVF6VmDGW8NAgZ+q5s
WXkpGzQNweLO6LI6rP1Ah1PaL6JdaqLhNrIuFosP8ArdbQsmzNcN0Fhu4VXLR41M2BzdP+4/w4wP
V503C67S9iGYZ40djR5lEZAa1e2YruKo7EExsFoEhQkrAOUf3YUgwngMH5aXNnH9AVNyZxOIuXPH
K6SOhCKXF6YtH8krYx5yQGtUzQTWI3ECbBfR75tNwC7xLw6Z0D1I6ZGFClTZWEpfTaB2/+gFVDHF
ckxWiJstOnS1ZhtyeT7LykSA5L9lNlre0PLyeqLmVq+ll6Mr92hjSeqghyrm+tr7rNvvf5sXTo4a
znQ5E7s6NIRZFhQX6D4nXx/kX/Q65rQmJXJes71oZSWYSE9cBM5tbv7SMFUcIxLC3Y8siG205UIt
g80PzgNwyj+H7JVU914P7uH+V3NcX4O4e7PwvBaOqQwW/IsSjuR9OhbT4k/HTVrqbY0P956isrUM
XCPUIqDeKPUdwOb0oBDITHahwixvsGX4nOcZnxWjk4t5kN/+89yocaTlaov2bmrHXvq/4kp3k2D5
MysljW0mS+3pP19PQdWjZeIUq5OO5OGr5MIdXTpf8LKIa4ZjRYOiBmMFCiL75CJcCO/1ENAgodpw
TLQzs3trQNFrNRKohS7JUXDF2oTcEyLSnrixBNsu4cl0HsdAz1cvjb9hh9LTcf4Csb9qDdX8tSPG
KVe8X5pitpLuNADvrVex+ncksrK+JzYxsnxnRkJ5MOEMsPlywFMtmmuj7/Xxk9hu8RjaFvOaMu4P
cd0kIIgjYOk6Au/I3uOO2Gcq1Tw1rAGYjamlB+3mfKbkL+jgE87TApGmBIAkpco54fJaJkCwxLof
9Ib7A2XZtZcWv3df6P89Y5TVP90kkDmjO5wH9sCsNViLcaKEk6tdqyi0a6bgl++Mt+TbEMITxn+p
lnJvNilkwahmSRXLD43+gTH4Hg7j49UUjojMkAwsrSX4BSF9wZIY648TeAJ+nXZyh3HksbH2XscS
onGez/65fTvOAbhDvjYYJHBKZa+eL81HNdqIxfE+3v+pF8Gs4k2qsafA/wcP+3mVqnSc8SULC6Yn
r1/lljhbnwiuBi05XznnCD2OhU5B35SDIKrG4Vuhfqz/hLluwIGW55PxqBoGSg11z9cpDG6cVUkS
HWP/HhNUaLtalfHRHQXTcQto+Mn7EIZIEQzV5ZN0g7TT78dD9Y82H5ZMJaUD5X6l9fSuJ+zH5c3s
vntbzZxuD72n3vbhlKIFwZGvA+dDXs+CyEFDqOIPMULszXwXnrcfKyyYl6zuRcFkd/zE3BhBRULJ
dsKZO37gKIW3rmz5skSxsjbyyRKqJZHlh4nMTqvkfTdRiHzrfLTDe+zjFipnwUziQh906KeYKCSt
joogqDbHGUk/2wE/DcLuSL0E4s0LWW78U49OAIcVLo9GXMPdH4mm5WDdy4rtkPdxTkULzVhAKlK9
vGztvtrRjJRAqzSLYelNXW58GvjHZD24Bd98n8m5ZdeR+y9PPu4nfyZMbl+RVFf5WE9Pd/oA2XXx
YKgf2IhalgDntRpXlI1yjQSudoIGDPkNodYqKu654sEuAG3j1lGg+Z6hzkRxtK9YPrhlrMl8NGST
BaNFf4s4O8iJBXItR/AAVamnSH78UgT2CeHHVMEdJTwfQmR1FLQ1Md3gX+se8+V/orQ3W7zfoS4h
Nvt3hzP4WIu+UvtCJfneawQ/Y7ce01Q17XInB4F8AzyWrifZZ9jN5qTC9UHXJNbQZU1azJ5S94gu
F5ZEajEeRKHJbIjXBfHuuT3RwXrZk2kZ9ozCrT1lOapotIzT0Fss3iLt2kCicDUMg3zMDW5jHnyD
PAGaqn6a40lBO7VdJetIhCdJHYsIwE8Genv7RyQHO6AGKGqftxAv/xpflY2P9L8n8H9Ka2g8jahE
0maFuX7Wq5c0iP7UisfzvCao3U73IvgqQqxjlPGlo2UqcRwdbw8F4t1ZLIVsZOAv7lIp7B3VAuCt
1Y5n81ktZ8xqOWXLatk/Iwn+1LQpkvrb4YGjkcAF0mOcbBbmjlfBZtjynElpWRvB/PJQcfTB4W/V
+pSVdTyMuXe2RnEbJmpnta0zJctz7yrllg0gkUYWj7nU6Q7wO0AN3MSWbSN7ivUkAXWhjZZe4NgX
ISCcMCCR5eGLkWWsnu959tZkseCM/EoNQyznkCECK/f1sHRA00N02n1DaJULSbCR3RoNFGN3zb6O
M7LJ6D+3CYEv97rfFpGM+ecfdiI6oklDBP27rQscaJyZ8xKWAqttonk94rHG1YswAzkfUVHzh97p
MoMC9BXfGrsr/WKD/RkrrMQ8f2JGvAz4or+JiXyjH20Ov8CfRG/mst+twd4Js08is6Rb2lmaDYup
VMOkHSqAiLtHas73xIjCdj5Gr3G/mXLU0eVLIFk9uZphhikVPq4Q75ZxS8jTban+dpoAU13WQ+7q
meXG4159851bh8HKjcPtKAXC1ch/QTNoihNrRKgRaiIchlY2fTLJrU2u/UMeuzg/Hn1x1XDGaL89
3NMEKx4jsLK793WRMjmfl9FlP0EAbPCtmSf2J1nu14Pdx1RX+0BMA2bReUcMqNG12zwWsyAuUfaI
DLhJBGycnPoqxtg4GnVDq5084EInaN53p1/xTmNV2JzOWWtjGiYG/toGo7EmZ7zRE3AQBM1A7Fvy
SEsnoqf1b7lfy/Fbf3ME3tWR1PjcGfmbLKeVW5j9eG34UAmhBeftUH/RuMp89goUehvpeBAvKwPz
y8Fvy7bd629kwB/XlWx2FjPYwnI/Ww2APb9+9vYz0OA17bprTGvE11ggP479/S8Gw39LjyAM9QfJ
dfeWe6EQ9bIVCkKbA/8V0CZFLt9ejPIDqqRa1GMI/qNC+W5Pznr5ruqpfakUA2VGjnchPwbHoq1E
hXzbnQlXPFHE3hZLQi+Y0VzyFJc5kfHVgGnUCYEMi28Wh1vHGXc779WGrAPK+CkWSTgPjeRFjPKO
ZmPvnXKHJFCwmKeTxf+VPoI0HPGH6NV2BB93DGIOqGPrsnGN+IpRabmGXP9+lIEkLYxzOhKWTa5k
Sgs3tVmozyVKOScDCrXnIzSGTM8mT+CgylCWPPNlnHBDPYg1/r2YM0QSxHTlAEhoWBVgxsEr/geq
M1V3sBQ6yD1kwjRBLfWzHl8a2H1jyNqyOQWedKiILMiukYUpo3zP0rbR7Z0gRt9lIL3oLQeJp4wy
g/WlWMzgzA6ZSzGJGc9leEBR/ncxCYlW0kjdXi+Lu6prkeqJm+Q5q/lKtYhV10iblkSCUNVTtsQa
k/zh+SmXSSoNTWvhYWbfcIkmGyYElW9IERCU0TJMRrkyRaXiFK+P2XN9NGnczfK/Cq0jViRgpe03
iTMDZ3Nn9Wx2zXQerbS+JZtcov2OmxHv8iQrN9Us33n6V60jLOIedXnHLYlOE1GiAD9Kp6NZM9Ws
0GKq++tkwqk/3UxrJhjUfnAc3fHhzdrfZkFONBxfO8J67imFlDCBDCrrYxtXRJY9DV9aejtXviy/
C1LBj3LLMmT7MtqrBGt7muxvwTB0/OBjP1LqWF0zp+NDeBLZvKyS1ZICdjfn5pvy9iU4WyQlD/3o
MmqsS26l39XIORU7APE2cKECm+xqfgZ2QMT4IUD0MbblE4Q9f8C8LRdHXUAW0RJBhExOhES36OIh
DZcraBzUWgFg+ttRiGXk6GM4GtS8/MytjzAAgR4K+bHuUao6bKkhfi+cyx8h42ipZUGIUJeM6708
nP1QVejHc4grGmf/+zRgCLNhsAK6eVPXYnj4FPgZcHXwPl0X4jc1OcK9tpeHTajHvkhHoBLAEuL+
RGSPAAH9MulmCG3nRjvJqTcJuKcjqDgbb47qkrh4x+EsV8yQ8IxTtEKdU5THk9cQwHy5XEQxxHqy
uqRVDoulVhXn6Ym03I4VHEQcNooeAuUjAIzcEoPQIpJXivuLAH8iYuO2FV+nOwTha/16NXdofouH
0z/XN0eBc4SAkTBuyrV9Z2YeZQBIqC8RWK9qhxvNkU8wkCll0c+HouagpJe5iyID4YysTHvGxSWA
LgTj/S0cK5vLonDKHvRDxtRXiyFULeL0uWQaDWaR6MDcCaGg4vRqact26qJOKb5FjQ+tJFKDfVNO
3NDXvC3hrOKfUHBtO6bRI3D1d0X1Bc6U3C2KKiVPzm2LBzJxqgNfvbMB1GiI7PRZu2fIyaO005XD
RL5K/Jhamdyc2TQMXHwgMKH8OPnaTNYkuYs+RMUiyCPYtvJm8w7KVIxewV+yFfeAxXRGjRngpb2Z
TDV7Tlpd78qGLVgp5a7ha8xqVMo7IPm2Q1KUcY0gRswOSkGc1NcIkLlid50nEVoGeC8cP/+PBuIG
BDBH/OWgp68MDRnPSnRdfIL6wMGHHETc92uVjgINYRSZYbKjetxagmoTCoHgKNoH/QHCYioyWqGd
78BdqGQ8qWL98yCe9VB4ukLF0ar7g1PXUvJyu1o3b2haszzpppWZpfeJnjLTD1RC9q7xs/RmPLKK
K+JZhFx9GjJknI75kJg0EJPvrY4QLQaBuDRvHsCSofSr/dXs4PslwlOhOUWLCOLv7ctkjzKFxx0+
12vBrBZ70qUWyAaBcNSQcLxNHdCs8Yj0IcjKTHlFFIQ/7QkzOGFZU6ssqk4g9xezxlZY51iYBWws
cYRjG8KdVjhi/krL1rCgsKQ3jwIDDjBkRiOdTTUt0FkkmVkqpCgWbGsgyPmSn2dzH4tcYa/stMc8
tTH47CNenKoxlAFCHOFSXpAGdJERSFOg/hXOc07PA4Tc955uGeKP87vaiuvS2PgK1jpGo0OKxm3Z
hjbC84ntSRyaxaelDKZq41dETg2vNWMKqBClY4g84D3bkhyOSMIxC6w/kOEm/WFKJVSQlCgaNSi7
1RkVYo91LJNeuFL1kmyTO/W3v2wcrl4PVYHLJphnnPCFLEf1fqylErDmoyn8yQ59bx7EDNcIVelo
CyYLaQvhgEJfsn/uMrwIHsZ4H+wefdKNJnDtASZzNiVeWSuW6DJoamp1fp3kN5x3/sPLN/jQHeSR
kJlTYKnfMUMqfSpi4QMFLGQuJj6A0rL0SQzZl9PfDAlBv3Zmyk0fda44WS74a1qX43cLBefTOjHi
VdtnJB55zzqFxXp13qilh2iCO4NI/ZzrdlXwaNRthoDNwev/ncOLghXoXQkMRjXVCpj1bOT4MplD
ukpjNmlG2NuD49JV+3sRYxicvLl/0cVrM7Qvz7XdGbHP079eYzcFbr5gFHGo7OhD6bJluBa5+DyL
E5lIEXKITcJh4oX3SY3euc/oACsqRCQHzjDcuXPVtgZTqP8GVwKBKdUxTk7eXJkhcWQw6bThYMn7
2O1YQsZ670M6zGa9c+kP2Qz9TMIS6hajh7mIHZKg4CGupzkrUQ2t2H05bgep13ScrgBT3wVB7xdK
1QcF6AjPGCGk3cOKLAKn4rOZ5GO43l3Fr+L4JNu1BVaI4uL/ZrRyTmzgF7zi//1t9sV0PBpGT/u3
Fdf0g2sj/JfUrOuBV6f0hTI2a5L0S5c5HxyTV0YB+ad/5qN/2SoHw+VzDB3bvWMUzyUjyG6sf05F
Erue9WMW1gh2gZn4USFRs27fl8fPuobMghTKxA56pyOlSXwYl9sbG5AtXHjMOiqGZ8vFLQxeKZ35
TVDPpiu2ZSYzzX0Awq9aEGuIZ/t/kpq0SKo32Hbo/CStWYal1QUVrzhdK4AOnAS8vjKWYK9O7sO6
ims6kirxLeo/aHyHVGUheb3PO1laGJe5/HXszXGuONxxsadZRqKqXAF/on5iC7lOUHNnToJ0HQOS
xfXVNUxU1sBxoSxiAah7dsitu8sTDTCQStD8fxtn2B387lVKEt89llhIDELSE8si8FDtxAb6nfbJ
er1iTiK3N14aWOWZQOyJonZPP2uyS2XHvDmQv5AMKkWSAKM7CNb5/7Yo7t8Zq9H5JO+VWOJKXHUJ
IB4xELXHnaZ23QvL2c3yxAv6SaDb/v0xc4jzbFNcskftnZxdNDa/dF9EHFu8VkTF/nu65mn0r47j
9jGO/eTQaHvCpRy5APsRFeV46SMcRb9X3YLHJr1d4U1b2EZLdLyCR1qAqjgzD/C2tKhw/6/wyJ1U
l8cgJJUa5tG8Zpb+OMt8C0I+xLmY1KQfLZXiaj1kKHwjjGS42YlqmUiIgrPusG5I2nA/DucTVLX2
Wmx8N2CktIdrQSY/VETpCpigvhjCG+L0dpgjtGexXTjSo8A0pZGdnVSn60G02nrSuj37+gZV57VU
4r40o27gqqgzN9qiIOb4vL9KjlOkdQWIT1rbpIfQtAj2bZcQ2cJ65af24MCpnjlLQz9wrU5KFfWB
ECeDjdh261ERNEw05aZQti4wyAW4XunRX9kWLVTWkC38uNOCGyX6THK7IChWXwSZQna43Hj1inlH
tYDF/7ytLoB+6rLRkE4fM4vSYyS/0z6equkkqK7FR9r+vP2zSztBUG+1rVewjJd7vENDq1RL3aM/
U7l41Z0hrMv/BE+Gq/QgaBeO5Ae6fXu6UaO57183p989LTnBszQ/s7W5LcNrfgGozLNVa/uNDxGW
29cRMWErdE1TuyVsYSAw2Dg43OdUNAd51DyPGjdy2VVAoFp09S1OESiCu0uPELsNYzPJcv0PFIXc
Fkt42QjZcR05nkvgNYaU5wTY2ZMwWqlbvruufODWnQOXCHlkNchMJiQxtB95WpwmtdYOc3u8D7Bt
LJ4/GeqzlznPiz88ZB7F1HMElr18Zu6PnJimwZCWmmlcYRbrapIDzB070NN3zmjN3X5oWyeB1a9J
SWBN2z27bjGD67iqk+6uYthpfELZm9NLyu38ecgmkoet12OE/MBq5+EBXOtdDxnMiHc95RIVCW5E
uk2ru93m0qlVwcSln8pub0TAL88GJ1eHJbnrwcjwYU9go4+wJTCA8o6YTG6pNAL4HSk6dlsINzxy
rU4+fDHbyc43FKi28U4L/+vnfLupGeRau+y3H/HVJ4izzS52Lbi7QigJfgsCsrbjDqz22kR1pTDC
5xrnKDS7rB/GPQzPrSo8oVZKc6yD/D6rcG38VQ/a/YSoJX/WJhBDC4x/+sX98OTz82SyYe4ev7Cp
TalAwsHmn+4VIEfCfBEjMcq8zFDp+Ne6DZxr+1fD09q7pV64md0NcBunZDesNn7l30xfWGPW3fxR
zCwG0jEl09Q/KGa30IPws6F2e1E0q78SB0eGl5RQBGCoFvsSMQhpyYsr+KFhP4QmWS+ElM8Z5tu0
LRmJ/OGRyEWrFfP75NhN4fmSazL/j/RJd+0yetU+Bw7Va+4w/U4CI6qf2OjT+6R2TFEBEGagxmI3
E5dykdyK/Oeve2Q4aPIqAKK/UU8cTNS+jaRTwCLxiRm3DTz4uNzuzIgXwDhoWvK7OShR5NINXava
Z7E8Fl/f4KW7xq12LIUd048wApWNfA/tDBXs35fDbc6OXc5vPu0IYQ7UfF71Ah3F/4UXJs+mSNIE
j3e5TtRqXsSNTueF3xAEqMCNoaRFerf47ZYeow0JhDwbmP9CK8TVg6bVl2SsaHlJB2lvK5osrv6o
u4ztGEqlXUtXkEGiQpeCDWvSYwiRXxkGz7HTkRnO5621mfzzS6k6NNm/tZlcSShz2iU+xAyUeEtz
V9sTQ5BpDesEhIbnZzL4w96Uh/AGusoui6XAMRMgsMOp45nVKg6ukDlT+tdR9sTCBjhmJ1vqEZ1X
Et9S6YTn9eeHck8PcZYDUzf0nnO4s4lO9xPyX9YuZMQkEOVTdkIGc14Bq+cB1l317GJCq+nOZpGM
vdNZR/NABbBt+q8ZekvspoCYBwwyu290ThwsYU+RnVpmW1JjVGoqbPUZWH+w7VBqoErx4d4FNYLa
ViBefQAfTz0mLvF4k/wAuMThaA9JeYwu/xQlINMJZ1vjSpEHjv80Yj9XuK5ghvLzhZl/0N8aBIT8
FryOxk0u7poKQUDJMUINmAM2fGcwNbROJxoUhRsYnJ5RT72tnGr302UImP6tFEVVxNz6hq6r3XMv
aFkdm/w18uIn7eZFDrbkVw+2LQLTT07BFzQBmVBcU7yPrUPzeXOoViXhBKt85Fr5Po5d+OYTObBj
F2B748oFaEvtJNsyuewf+Mwi6KDv4PyApJKoVFUaTU9VSqhc1LH3HN1TB8xMCtPyR130718tF1RI
YKUkNkPGMSV57Ds/v4RFenlbrC9QQQMR+Ak9z4AStOCJuuOU0CHbuHgFAkCNkSoyFGlKhjZhEGGZ
KhV/PZMak96zKZKW+jvqQMp2GFOY9CfzFpShCfkrboisuoogWavi0bcDdK/v+WN1enHSZKxxXL0u
c97paDFxwSSRUBV/8RI5geLJm9lHeY0hEqtXqsn5ksL9otrxQkdFBzBrnYBu+Gmhpmh41Zhv+3ke
dKDkNYQMKVcHcC6BpIN7H6UX7HySeXtdfu7QWLNGUCLWxYXF1yjbiJr2nVmEvvavnbv+k9RqPIyp
14CJay+zlVNEmUAdA+8dDXtaK77a5dwlSed1Mb4kGqZs1lizKIQc1/XHRyDdb84uZ+imWNceFiKW
jyFnH5Yw4kN4CLpGDtTOZQwb5ZiYwEUcdZ/O3dcqYOzJPla9V0RFrM+Rs5VrRJ1altnWar2psaiu
+G2C9G4yxMuBQPywjKO/TIY0hZvWqx44nuKYameKhcdiZDnTMfBENIf46TKC/2lfwxj6JEZwZXPp
p7Xr6AcRuypJd3uLffbc87Khoi6xfDQb7hqJkHsApec+Z9Dyacw9fLuv8ca3Elgek/91kgdby/7q
/WbljUU+q6SLDjZZZouvan712co0FcGZ/GGTxiYZOpZmgvjBj74JVFDS6ox5YDLHH4JzZ1BbF8qs
dRE3X32J62ZbLmOJ4zm0aFGkd5OWcZWuDPxwUm93STN5OCTy0ABlNtCLt8f3t+Yq/tfNyYzkgZep
VreV4CkdtN3FGCipD5XKdGVViy95ajpiRHC8Auftu3LmAQkmIBYITwP1szxZ9mnIULBAuAbyDTMK
bkDxbAGSkhWvql54W/qbQ6suzQbjpYZM/0Qj56go54x5jHXSsnTxQktHDrPMs2oJPEux0d7GPVNz
fM0XTy5egOcp3eq+ZoL16Icme6AExutqKWN7HdE7OjttP9WlAauloGqiZ7SeXBg3/rjrTkoNMO3z
Ogl312iZuujwiSdRnAe6999tlkiYX0rkqHNongE8eleq+sPnBCztYkxkOuQu5SXAoDAdrnNs1nOE
DGToSnB0bCLgKUARQ5a4uZbzBC6u5bkp0ffHm+eQgdALXdVkWvC8OmakDfG6fYYDHsH14fNRjfVy
4VQARHhxHEBRw3OHBG74vTrATGECx+wrMEnR+WbPyfZ959mBGsH9IAmdg3vbiWZTesU4+hDhCt2h
eOD4gt3VrGEOG+OEHJZ18PqKWrVerV0jlzWXDPOb27QFoPVkzbDqnFctAyf7e1VpYy6smUmtoBnH
FSHJOqyl/8keHgXtFdR+H5IBS2pJAQHYdqm4KmJ/+vGA2tZ1E+HFS/bJ9+tGGzbaeuytd9UQgxGW
bp01nOxYtolkEj/kMlt94Vw8UzueA/V3/MQF9GaYgkr5rZ+F8784FXPVV9s8JvWJ0UU6O6hkDwqp
L9rhOa6+fyy/eUCfDyRwTlXb6kQ/lPOabtSZ+8o8wSuVriNmEFbjcnXKqX0KyfpCgdjBJqrYAINS
MeJJ+A/rdIwhsUFnmlotuzFUMS6zE+WJPEc8L/PkXwjfv2KbpVZvwaST2puAsqQGPg9vVMgF7pPY
xVZlsRFOf1SWza34JKRPMYkwT7vl8StCvOsMx9EpvjY8UNVzG/tsI+B9d9PAKsILywCqLtwE/n9O
nN5q9liwnapv99CVRlmRh4j6a/iLMIiAFJe3xUl32fTytBVau/FP5fOgMVOzdzYtcbInfGgSVqpc
4/kMzy8jLf5gUfRZe8URrfHDqg8mAUmAZ2yDOi1syW6G08L/vGH2BYwmRHJjujO11LEz9MyCDlc2
QgZvvPHXgYga0S2/YXC8JgAOvTh1w7/fa/1Qkuq35MBb5Zqpo/TdPueRov1OXjPxpWrRI9cjHP6g
4AqYiR/gBIrJbz+h8kE54S2XG+SwtlWg8KEwgzNBhEBdeIKwQErdLRw68nNdH5y8/pUUaGE2rIE4
muq3YxXyXeNsRms6ztRt12DBAUbW40MPerZqE61Jufr3M5LeY2E2ac2qpjNK8LEjYFiFr+jPHuKE
ojWyO1EQAlHZjj7T+sTQuvOLY5JCw14UEV974D7iOSE7bKwoB3wwBSWYmoFoXzAaNV71VBujtxmL
T3QwAaPlVTQVEHmo6KG8vOssuXCnQgc8qQbV8d1w4NdcWRHQuqGUnh26vkbEPYhz3jDRrl611YMQ
KwF94oJQ2hNyi0VXdvf5gl7UEMFXTghY12rk2V8haAE27wwBIym2tLZC3snWYgTTfLYFMWVksdfm
jsI/735T7EDaHppz6fpvhZbDSUoUsQuQU2pDUX7I1TpXku34vqWAykU5/6QVkarASV5+E5njX+te
NP8Eu0HiiKafDn4sYUZtpiBcFLMOANGvmH3E70QCOyZ+vn3SIpiG864h8hA0Ijd0fvwl+oAgog1v
uwZ1FC3FzXqgHA1bwq2I6/cT+owdF/vF+uSRAzh+fgdFwcEMdOkMA/3RfsKHSRcFoTSM3l5L40vU
xj8Q+wHJCYidVZz2/aCMpX4i2XyBcduvzLWFlOodjDYBzDzv2tPOGJgA1mjP5Cd4jkfvuOvRIDAe
WZDn5maNCFGc4tDRvmnRXkSNGYQPk8SkqU72/hD7/uzOtuld6AKb4Z94mQklOjGDPYtGBS8BDp04
Y26W+S9/wrQWZNgPQlcEwt21sT6GtMmXVWc1+GvSl5xElUrUS0iSaH8DOYzjZZnGjfD5ZB2m1ca4
xbLU+2j7ZlUeLPMOh7M2eBiruVzV7eoUn98RfO/LbwZvHuqhMgWs38KqWp/n8aI3chzQhaMwzQYs
IzlYJXUrGx/o3boljyUZuLEjd8LNUbt0EXcgNH7hV9iK9dssia1igyXMehZ+L4EpuG+oxaDoghIr
FCSlFkTsvclv9EVickQA6lc5FJdToMZhijR9degjk1GBNp3uaFXTg4Ln1J92+3S9iBiYO6PBQ857
EhkrbLlJNRujUaoQHQb2cq/hOIq9zErdPtZSHTg4F7uMn/FntmlvM9q1M7BJdrP3Pm3hwvR8c/FZ
OV4VykoqDSziKq7kgXswdEIcp4xAHyvMvkgKrvm3kwWwb26BMlPAvP6IZCaRngkxVgHl2c2d5UO+
QgQU3p/57CTcW3sFwi8T7NbMAGRg0e6AN3szgrDRSTMMA9vLT5wwHg5izF22xW2SWlVLsPvlzEhN
OInoq4VJaoGcgvDPryVgW3zOm13zJ5nr6wkZA3TSjeKEMMuLeZ6FaUSOVVDEKNrYWA4adzy/eAGJ
eiSJzmqXVHeLPtDOYmO320hn29YvUUxvEumOPdf2rHmcppmNtb0hE/zL469ujK7d98vfzixu7cdh
6OtJMLduUpqmuodasnWPzr6o82Z+kzh6QKnbe84YpwE6LAEiMEKEwFrPTWc3XUbHJe+kwcZemsLk
v8vDSSMbWcdwV4q7KSZPC3hnYmCVJExJubURPAXO73o5rvlsNE3Siai8e2Gp6UjphWrSBJd6UbqZ
4z/bCuLYruKBjA6HdsMecgziqQXHDOl0jnh/cU9pTO6n5L4d83HTW90lBO9pxJWftGwIuBsIuag6
THK6pyFwupRJWGes2GUkZ4UJEvAHxo4SoD/CZfcOPcrkzDvtjqxxHLNexLhe3ZoQZVgm4z3g/lcn
oHLS9psETUwyUzHgvmWQel9NwGtQ/QX7OluGZvzXAD497V1s6K7+vk9Wdu0TKUOAh8GeejKBwXey
UC3Tx3YQwWynm/Tgi/sI+rFP8Xal5w/IqoGD980Dn5pEudr3PTMCTxgtMwJ8Vgt3Vwim5zAEkfNc
27PqYHeM/RSDtBOnWdJUR5+j0e5GW/f8ZyTmLU3FBb4Toxa0j/fHOdcgVxSTwY21J/QHt7hmmZn5
IDSwYDNjvv7+Ae7zAFAcGPseR6YSbDuRuN3hgSh2fifluuBqMvnNcx1NJDjUYo9WUiqglnp6Xgyj
5bnjvZjpXcTyJd6Pq57ikYhpbPpaP97LWtEG7cCmZ7hske6jBijB5CDue+q1oXTjnmfJ8pxVE6cF
TdIUK0Gn3SctD3IXJHy1lOFLHuO9YJgGWqKcAQLUjJ8PHM8rPCB+cPpJpCOlv+biWNAKNW0AEe/B
az8SIGcdBf5VTbDiQJ46I9lBO3yD+jwDR/libDH17o3shuoLlR9cY2i4HcsYv5DA7nw7DXmZXfnE
YXhD6wOLd29bxYVz6uhTjnjU4/n4lTCjf83Nfs3RpG9FylLkm5PlxkjHN1Rlrm/5afIsU7+8md89
MT8hxumEPHvBQKWDmbThuknLa6OH4BANhm5kiUoFpwrOrPF2G9FDwkBHt6H6tXXrH1k8Mfrv4+QJ
MMfjl6dd7xB0CIM+3DZnABn9wA6J0yErRRGNFxMnnIXvNM6HWwf0YNIk1P89rHpSDhTtuz3gCAAr
hho2gNB/f9v7M6AGGYMK6JKqVLwlvF3+fBEeMDSoKuunXQf75AulZo+/4y9id/t1vvAxn+orbaaE
kFlTGSSeqYPu03yf4xhWPRDaHl0sBESV3MNTugsskzASiVFwkOYrcxRmndhDmmHBswRUJEOAk02r
cGmxfa/o6ZOE2Va+ecENcOOt2YQ90eTe1vK/92P5fY5NsN93zzqp/N5Rf2ZMZWJnGVUYrpHUDfNs
wvMhoutPajSXW5N8QvrGGdwajsxSpeI/l8wzA4fDs23XjqM/BWlyiJD7x5MFSm40QnO9eRfOcNs/
EaTuMeeK3UBiZpmgfKj0fFWNoaD0Npb21wD52/Wy57KaHg2VpyskZRcKwBrwSguHr5JHv+9VO2Kr
CG+SH+XqnUbNZmeQU+4ipaHfZcKfOgc/IGpQc35ZgpRk1YXl2Dbwq7TpKKfQ4lGDsXQxbYesKAp0
1FURabM2r5UEl4pDZyaN5ZG98jK6T1IA0g9pefAPR6sJAhytEMFVRPFMTngdeuNEx3srp1kAtF49
iv08Rq3jT14z+Np4qahZXL3T2DcViJBQd5RulsSw4L+aYvDPoIC7SZm+slDNu4+Dw3BiFQDgOR5m
MjR2YSyYQoJTXqIIkPGTJidL9CqeK2PHhaQhN8OFT5riQe8fIEu1rdPR0JTdSYK7uuqFDTDlPRAx
h31GYAfqk9KQP8O7RK7XwFQVLZRtpepbGyd7sKVAsgfwYNNM0I8AU4OQ5JPokAuLbYp3NEsGImHj
olUEYpxTWb6myrOrOMv6DsCRReu1denASBVILiWb6M2VZyQzInwOyAUM8I5DpjJt3hWqguvAjY6H
vIa2YsmmsV0tlwa1g9ND0Ev1hsQAyU/T0vVLjMIVV7bzWTgjVqnU12Ypo0TSL6IOXHGgbSd7cS5O
QNFnwMUM/8yhkJNdT3HRqgpwVFp5mho4FiIXc2v4mQ1OanEAybpVU9II6QDNLZV0VPKCafyWRxiC
h3JY2V9aYtrDCLZjQqkulBrYkk2yTUWRbWaONZzJoAwc1H7VQH0QgA4AMdU3I6WIA8CsmkexEvt9
TCZG3USII2JqsxBkPqgOOs1O64JnXrRppENdjQtyTxqLax5G6rqftd3sOI+4KMlMfoqHibKNc+XN
173rvFOqxkp76a/HbNpJrBNb/ngtE4QFNQ2OC4tizEtQRmXmPutJM902Sl6nERX9ksH9Tq+k6Pp/
D3TjryXLOIh+5kQpVQdt5vr3UPy2ZsmlIirtL42puIRb5mdSTTFKF5MpkAaw7Vmv2LqekQMU1mg8
ymQ2d6s1JTkG8FESnZjoS59Rlxrg6kEazc99JNRzN6runWMamln7BCTjej8P6AHxg0x9M9YbhqQ5
ZkxROSt6TlLDEc91WvgWQKMOyn1kAS0d8/DzYVF8MwJOuNtOULTuZ5S2WRff03B3V7rIolH/ERgo
0ZIXp3OyarzIXevpRy2lnqXOe6jAoaZaK2m1q/JbXa0g95RcV5UDG9DFgp3Z0C4hGGMzn71JpNAf
/5k26TbhQvPBYVrCsyBI9tmi3syQDAkfX+wzjvnEOSUOp3anrbnWKmkepVQQmdlc1Z67Onbb4c2N
ZshjdF1uL68FLYbW6+KgWODx4GM33fBUgVw7KwDtQxBt1xn5Lj8d49irCkYvA29WX9lpuAEl2aG7
ejtaDFU2IU9tN/FtBWnvUlrAHGHtyjmSlgdhwLb/hORY/l2BNzoXhN6CLgEYGo/j6pLL8r5p8s3Z
ogge7SCQhCi6jDixGzV5h2Z6pRQf1ElMTtRzk6zZp7QEl/jKHmAhBz6Oq04x6U1WINQdQYuyDmcb
7bjkUnzlJtZDWH6QSybnzi+gbxf08nJSPO33s02E0Xjxk/9chE98YAlh0BHnUk6L2+OX4SOROLzs
wvR/4gh43OTjDKbwJTDHHfdZpifGYi13ZSZCKL3Ro72k43UnPam5B8kWKD8pqdzhWLvHT9mbcFxf
2TamdBbEn0V7PAWj61kKc8JzbUFb8c0yruDoaLlqiUDvMYcY75Tf9V6SkkjC1bsMsjCn/j5tpZZv
g9owmYwp3wcwwSLHiPaXJo1va65dIjyOr1zLPh+t2pJ8/F6LtsyynDiSk0oR2PdgW7BMF0f6hZEp
xMXRApJIxFmic0gMzRcwlmtCqbhpVK2jmMeaOLF+V3D3YhwVV+flu7Hp0qF7+bAdmeQylvlCKLEc
D6q9pocMJB+sdph4E/Qxb8ebzI0v3q3nk/NuJwleXmqGCwxWB5rROOlSUU5ffaZCXJibd3hXLPf3
mu+BAlLvdOT32+CTIlY0NQlRW79wvHQIgVbTXnUokB9euQWs0DDsnxwlloY4oo5q4Npw2K0P4xy0
YHCt4fyKAClpPjCs7R7eYqAr4Lw4z1dkQFIt+2kzbVUOl5gi5xhC1kdhe/WAYt/x92Ezk4FjZi6m
IVa40AhMXmrvZwC2msT3qYXNbJ7nWpx0Ttp+33vKL2fmt83V4Ie7ITGo+f/9cCqZVpQablVYcOyO
soJ/3egRydPUffqjaFfPmX3DvhjPD4RDplnyVvfqy+DVGhQtdrYxFJBl4SLBtY7emkV6i9Zswi+u
ynDwytHfw6GcX/2VSPgIBoKILYFadt0OsD4O+RHUsitE8r0mOG4u4mUOzzJATTFIUhyhTHj0QYiD
EIzg5LE+zqNFGKiXOiQkIoZS3xMfpqu8ZN2yDt/fBSDJLcA7Z1wKsO6GzNBnsR838UBcT8Dn03cz
WT9o2rY57u4RJJNO5ltu63TnYRzuhRnF1b9Bw2tLbKs7E2nAc8pr96Qe4sMVVGGloqczVOSG1jVI
UrOJS02ULlXPU3mtoU8S/IkBAZv2IVenU0O/5Hljj+N3TOwSkKRh5dQZ09F877JgtZKuQRZMZ0DS
NwLfmjSLaQBYxGrL337yPLC2nplN5BNK2xmR+VcLPXo3jY0vBuVB05O2+KDrVyQ6vIM6d8/JE82E
GnhN+TsddnTyhy8+RRPRBfrS0mec9W4X+10d6hYoMfwptoIvsTbQqNJyfctUvTDJf2V7doraiecX
s9rJwzHiJBP/Rp5BWNzVT5u0xK6f8qJSGcKWhkDD8z2k4TuXaYMhWW984eB4kC5hr9iQ6PUFY+1Y
y9DpFeBVgx2ZUZccPBDXW/DXG95CRW0J8aJKCEqAo6iJSrtSfY7oOuznHh5tQMtDPw/+2230cGQe
evThkNGaOLZp5yTA9XwpEi5cAD3TmiZSZcGT27Sb3UqRkid/S2pQZs9vqgGaqyHJMjfgyQ0xaMyV
TZusSjnGfBz2ThfR6IXKoONi2xJHRnQEq9Xq6q5joNEQZh78QggdtlPk2MIsxGg8cFfoGFT+ETxk
ZpekvJfnUtIJE0NwV0dyvwwfE6CkW6/jNRTf63QrlaRHpoOO+wHjRiHUjzYrI6bilrvLaNpVmkei
Bu2NPaSJ9TwuPeKU1CGc9yulKvauTeqK8DTRZG+6yhrkWwVWiYahvMwQkuW33ARo0U9IufNPrqNk
KnjTgh6WWpesXQqxVFiu83WbRBCSelPq2PrYJXiGaK0XBzBCXCMZJGOgR5bgQi4Ba/qEqRBof+d1
6SCbPXHRyF3apZm8UGBs8FuzbLVqzb4RYQhDi0f5FAZfemKGDfsjGyUTI3s3PZMCUHXU02hdgbW4
YzPikRCE32lpZqfKsQBI2cxkHflHcwM34oXKqFmQ19fJlFDm9C3rL+DfKIZvFvS6FzF2JqgqrdvV
DSSX2BB0Y0O3jEWpLIi36nBFihHb4DEwRPBLhavXHXz+b6Edju1j85x8G/M1X3hPBHMO0p43T1JP
UT3t7145/SX6C0dOhoNQSUUP1ylrn+dlXbXoJb6OZexIvpLjZz1W2mwo9vtEynoOWJCW2MoqN2ut
dQgBZSlqiBgz28leXYfyczc4tO/lNqrafHevOJ4NQ6/s5opzoHy0Cpqxvn1qjL8F9b2ud5N7SxY3
3dDlis8XzMzyr5LfYGNBAxXF6FzVLEJJ43tiU3KBYrX3O44P1b1ggvjqVQVkmA0Q0RH8mZFOdbA3
a0R87mRH8638EfFeekHkwUrfIOmh2AagYz/7qE/ao13TQv0qG1FYrzLkIRIVTJsmq1MTOTED72jB
NMRGpdXS7u65lpnN4DEwp46nSYalfUcn8iNz+0WMWTbX8biWaniapDP8ocacxsztjHnl1idyRVEA
odQ28mohq0NpMk+LMxDViOoio3Wr/XrTmUi7EYjBPBnqZwPF1uQOwjRx1l6tOO/hojb4yWIANISN
mLEbiuYBe0KOiVuDjHXVV/Xvouj6A1nM/9U9Mdt3VvfXE2UvPGTBYGPWs58grv6zShbwxrFoN6tn
AfzeZqiEgiIwk7gVJ5UEnaL+v6H2H64B3rMACl6L0ZECM/h1s2FG5VW4icuoGWj0LdzHnNBpn5rH
TmKOhP12K1isrTVivsfuob7jdvDwfYsRxIdyic/nS6RWKYcG2YbO34XdxSsuXx89hrEV82jXBZMK
B8Y+L7YiVLoT6Fm3TP28M7lo+L3eQ8fXzREaHgt82PhTe+TILtKMZOJVgaLF5X9hQo6rltIuWr6z
VhyVhTV6gN+p7LbJxEvr5Au50mu37KTEXfaXkNjqwONWkZB1QMdxbzYcn5Vy3Uq2wtU29AfbPIZC
HrbgAxEZd/FU9f5QG2KWFoDbti7PwjKFjAm33LAIm9ZAppWmpz0gtu8pkF2oQMRQLIMhrmtHFHGK
OaV8g6gJklMGmm3sfziJTNgY/CFhFdDEOUdKMDlJ06tf/ygmUXu1T3gwMdmSjhaHpfacKvw+krRT
WYjXCiKwIwSQFOymyHO+IBHGb+d7TYqv0kWbj8Rhud0XC/UrNpssI2DeMiYDL4zZ/ozy58NoGfaz
icn1fwTdvxu1oleSD505Af4NF4RCsiC6eSp/msPWT4nNCjY9XxTrY/Rc1fdb9SfBASFG9BxofSMG
KQocPLkPHxIrxYT9qm4xHnnjlcnIEOC5uqr7aqVAPCXTfbr0Y5csKNV7ayaf8RCAF+qELr3cb9Si
Tkeb26c3yAswcRQwV8yeSo3ORZlolrqk/wuAJftDnHY5y2gBXJ5zVz8A5TNvNrlNJ1ECQr6d7rkW
bb9HkRDeR0zrwFfdoswlsfHVLTwhkAg+xsOOg+2uoiboO5+fk6evgfmcXJZsziPIj9X2M+O7QK7V
ibuNJb1iBB8VERGGycVE82GiMv1nRN094nTw18kULz63iK4Mn+Uld19pDw0XVUcnkDJI5qgoXu1K
jN7GPD82n0T4VCi6VeDqyW9CIPEFV/RZFZi6ldUeQWUxKbsFKFwlmYFJfeQQeKTJYS6ZqE/6h0pA
+ttdCXyNiI6qlVMxOT+EQg4xVivXTRQ2egJN/5Z3p3OhIIf7PThSymfuB1KMkwXI0NRNm+TyL4hC
AgV7KwHdAi2xiPa3+ViUc/5NXt+irmAD9tQ6GugvCqgGmgCaOLTlHk/RsH+SwptqwD2u6aOrHFj7
j31uXssKqg/rIjo6PJrMT1q1EuLXWL/E/lJNlSJRg2YfdUiWAmaD5pTh/XABHrGrf8jGXe1Qmgtd
wFUuG6KGXKoTmsrayX0D63sKGixnGtVc2tSq4JwmNmdy4yZEGuG3KzVpW/S7mtcKnhQuIltWGLyw
l5OqL57x6OD39cY9H8XwDXpDoVDGIkn/0HI/+0Lj36zfmKMJxiA2pUMhTrEItotQvCqbLDUKfvbE
KXjXeDy9YSOmSu/BWQWcIlZHhOl2/A9Q+PkiVSvJv3gXnwPbqdWiDgQRDaA0U+VCCme4/LNmuhHr
dijj//OaHNgNabwRasVVH9dL9g0INRmjRIWdbZYpdJZs17jcMhMb9etdLqcxlsTuZwsR/H1JlzRW
tOxsAQXFQDxs3qOF66D+PU8CYAytDcoq7SX7OKvxf24M0V9ErWdsMDxEfDUp/KCyttX0drIbXdaG
7xMT5uuRi0KaVXbYS70UmzGtCCnJMjEWSDRfiNFqirY0bwnnZB4Q8mwwlnJXzJcf3V/swJw9qRC7
9258jXL3XJzTw/eBE/M0bQK/1HyP3ocYrd9Fh68zWLePHUAgVipcurUg0EXRdHanYOXMg4A40h9A
7uXG+yhrNtxsAtmdMXdjq7Ujfc9lc4U+vImEuYltdsX24VHG9fLpyBu1NbAoaZVptup9mq+no1jq
NAtqR68E00Kdqnu0m2lUtJeLl503T34n8EftCKde8z8ZkFDtrWwXm5AO4lN93cdHtw0OyMM7JUlq
roZ4Ox3we6pTVJg48h5VVns0t9j2Zs9cM0w7HpkMkfUlUP2H64mtGzXaEdln1bGRq5BtLUzF764R
2zbJ1dvASlUob8YyD50BeQMaBjCgDJ8pNuUA4DbEb+2gwk52zWDZhVQeudHFn1/dAHkBbKwMAsCW
ZvpNLss3gaSN1w6jDL2qmIEg3F9FccU2qObepBwlYirH1tNi9rusc/wq0s/OrWTHWXsNckHbhK+P
Fmj4XP36FUyxeKKRZUyt/vLQinJ/78UkNYg02pzfDVoQmZJzsbByb/oMgZEsdzpy8/AJw+iQNL3K
dVu7nPaA/zNq8+RH2MbKSn3JLCfjyc+qBC3X2ogShp0CQ19ZjtZ2FujnSY1olnNO3VIOA1P9PF7Y
VuMV+lYpNaz34mXj+SSFOT6PZqH7Mp5zAxeYPB8OFhzPICefQSGZLNzAF8hj5LA0hnUfe/Z743+c
ZiXUcYxVaNVfkEauvSv5vCpQ5wR6Qm1zLbwxVUYc9PvcIyEGVHLQOjEWD4FRl/0ff5JJLxCTYarm
3oFsbwDZ+q5SEDqcLYhv/zb1IHbeFaRh+OGpm4wngRgF0r1zJEHO0BiCY/2NVPTDwobjKZF/tj6s
7g5+aRSlxzvtKkaWrxJUMpZYZIwwJcHAXz6zuohJyVBPXA5niILIj1g/hRz1ouLBh6MYwG1RnJnr
WSgDjF9rKGDl7sXadMUmGX+fZnmtLlA34tbWk7Ckh9iXCmxbIG4gnK8c4aFjh768ygrKu1Uo8hYe
3DMKz2rWFojqLHcNBSL3iIj14ITylqwLUP3Txdo7ofy+ttsNkYEc/Ps2A/3JjTdvMoDDgtdAXT+T
UrTQQdVG7++FzT9TNP/t/oymg9A1jWCCHOPsaRN6RNOSLd94dCLd9r/NiTD67+NNIOM07PxWqnzC
7b20Aa+32fu1PRT9t7EQdErMgur2qkmqSQVLumfvz/Oy1NhC1LvmnPCG8gpUZuyAYPVS+L2nAMu4
cTkO/LTLOJplb5FnSWNArRawJmweMmbCofp6NdrLK+LeFC+D5dIZMHCItZRZL//CSaYNG95bHu/d
yl6aM26u5aunTy2wreanhZc8NsBPDV+JUVSwhlJuCcZsfTvJ+hWOUa3qJnSZxe0LwGbaQXAuAg6W
zUB8U77mPI/tj2QDTN7Nr5TbKWtcCFDqWWLrPuzYYUxfm227lTY7l/6n66b394RGSBLiaWpMjA9U
cIldVnpk78uFcrwU81N87Q6BsG2q+EMsiLvPoKsMXAxr05qM0ifsYckxUq1eOXZAUh8QcRd2RKop
3zq+TrBcVqjUgrr/mjdcNKc3RDXzIaXQeZIkGHEOiThrOsAjskEUE54vNI/0G/BwjSJWjM/hDJ6s
lxXxdkSsakjqD1/PiK7O2g6/jSU3zgclQ5Cm3NeaAyqFA6NQBht4Yfvb20hqBWNHlTQTAPW7P25a
m5l0Y73E2Q2kgOcAYJ9G+Phie6Nd2AXhL1ogYSglRKx0njIou7yiH7T0DBeB9NKBITTE7+yXXyQb
O0Ui+9srkwmcWRnf4AUqGIgV9MsbiG5Xfr8ucvYULLQG8lI6G+71LtxG3zlWJ9ZtLV6CGWesKnTZ
OgU9cetqSeiwkiDahkpnAoixgKcLueXwLtRU79gpjA0HJHazEwpG1Ye7XX8quoDw9oqaQlWFziFK
AIJT0RLhTy0JfCJyv3u9wgAW/VR6Fxk2FL3jJ//tIQpOrmUfMgTY+q79sTvygngGTTWdDyzYM8jk
XtSOyFLae5NyWADB4y+CayErZYlMvm11qu0y2RPQxovQZ/c2JYtX/hCsAiFkrmwgwUVb+SNnlvDw
7/3ajxpfFOtXtSIrgVIhfD3bUwaKA7JLiDwkkPBnElqW9uedqIU83irpJe06vP5coX3SIfGhWolm
5ezRwjB9oRWbTD65Kvp5hpPRIPISuKqCVrHyckTA6I6HGq1UAZoNnqOJ2+rktyOjkBV/57CajfLB
9RX6HVwD4UFCE8vdQx6QJ9DRaM2tr/uxl8d3/q/zVCNrFKiKL0upL9TgDAKWNy8LCVohQlyBLRw+
E22l7wGJl9O6vLs14WWQ1I+9WBq2YHexcvV0CBFvBjU2NsLDIl5N3V2I26KI7dKGtGGati4NXdD/
U/iMwYOjDMxAyjdrbVOxbrd8KZ2QBV2LI/R8aNf1IBj2QkaFB+MTsujjYL2T//Cp+Ktj86Up/Qp/
1g5LeOAzo2hCMo06Ksslnxo9r7PqU0DQKFFxrdaaO8+unv0ep9ij40oE6L0o5lIMnY3hCE2cCtpc
PLbgvwGm3DOGpOhNeHh+J/eWzXZ0drWHy1Y6+Fw2XKyIwV7MhLLwl26BYoaeqFbyKxDAKFoRkuTi
hxGFVFexny9yEfW7mz7FC7LhnhczIMtNEImlnbswIGWWcesG8HdNV+wSbhOgYNlPxqWsr8NeuL5z
VKwD4AXbXc+E6QB1IbgHLtzN8i/IoASkFaB9h+lSpVgstu6R1YbQu2x6ZBNJsMIuwPmSTKGmuF3H
0VFuUJkBmjENnx6wXzQ1BnllOXQ7c3FO3KYw24uF9V6IZzeqPBsq8fSfYSeOT4RnLtr/SYAjp96q
zW40Usd2EccHoxlwWGqjOWZgDn3nU0oVpo+q6KNu87zc8mJKz5dinVNrRTlg3N++XlHosU/RhnJQ
Vk1YrVo8SyML5q9dwHz/xQ8bckY9fchL0irf7sMdB801ktdny8AZzvXKxTsaQ/BCD0/gDcYlLaOH
/jebC70g51TqHmcyEtd3ve1cbIupHrm1kfaDYQhg4B267KmfFyBpXMx9DtrCLR7ZNcj3lZ4GeOSt
XeGKp/LsAW1aGmeeXTu0c7rNoWPvBoJjS7aRM1ffvtCgyDDKEkVdVx3vb3a5WyP1BCr/p6ZIkGOb
F1nXz58hSouvleJmuFmVmNl1hs9QkNr+gsZyVordx2crrnEMyGzkq+tp5YrAsEM3wAhmRYV4diHn
97I/k5usgg4k7VbypFPXvKQR6tw5SiFVAJ08o4yeCLMqpUkrgIWxdh1NBNSAtmVnuqijywNPhscZ
uneaN01K231kD7jH4LleHAjrODD4b84qPqlB9wWaR6DdQ28pTC+x2QAk31uEtTRAhySDYNMheJjZ
vQ2S9mgE3LP5sxj/qxP+LEYM8tNtNbQaJCRwMa5hPAEN01ODavvRLq8hbjTTpoQCav4V5DLFuFV0
mit7oNjf6d/kH/8q6Br4bWqZ2kdPIDaXYqhB2SBr8xXTGIJgxkX15tcpX7SJQ1v3X5RJkoJyDslW
VMx6ayAGCoiD4AzsxwIUByR0i7FXQbJbY8lYSMyv0AbT+8kpbDRpaxd67i9hUkTUkbV3xY9q4+pa
Ws5ZWJyHGE2YEVn/YbFTtgck7LD8pSRKcKmGt5J6p3TZEvYOKcb78OnC3v6SU8Ax8FxRjXZ37rrU
4WNiBbDV2ABWtr7KMMGpFBZKMDpKT2hOXdE8MryI56LFyFcyU4v5JQ2yQe/g4WyNeyBjI2EXsWCv
QVTHgSi8OFoOHvhOs/3rFmfGt4iipgz7Gnv0FNbtEdmU1qX2zNwCQab/Lf8ZzfQ1zUKz1dMaGGjK
PV4WgKkVBVU8Qc8osKm1mhL3bOQiHG+y8xZTv8Oxd1l/EPZ0JY/c+pRDuMwgA9NrtLMOrXp4TWNN
9yMYmIwvzfIoYyMOE2uO78uYjK2fqZHU4bm3gITyM40W5YUaEo9JGmc1qMGYTNUxcjmch9dtnVQe
6iW7PtBHMr0UOhXxeHrhRfdm7MlQvrBkHruYdlElUXG0B0EG715Vn3zPgmuXHQLpO2F+5Qnuojk7
quG85NMJhh1Aefg8Hh7fBzDPy8LpllOxffagWALvB1FlBF6s/9VEKPuZAOEATLBd1EEC8r+uYsU7
8eVgzRCjuT/jnW+ChNGLrvoR+ojlgIRq04KN/GA29nA7AKE9e+u2GY/rYP+nR4PIHEzAJWbIGhuq
TvmJ9tpbBWqPkGA4rePfPb4WQTYFHje2RqfsC9lE0weH+y/Ory76RFf2MsRI4BV9Bse3kBWPhjq0
UnSAmAhJxnwVnRAApdakIwdOkqDVzSsrTVBm7zTasO+ucYlO9/SlnEjUjRdsooZw5kFrLwH4p3EP
XPP9SUQgooBRrPNYTuF+srfNjo0d2AgFyYH82Qt5OtTpL4QznCHyT9vcrUb3GvjzLaP31p9Wa4Sc
PB52lDnYnRdSQex990TN44+Y9oyIos49DjoUz8GZPHyoH6MtloYwAaSDPJbWBdOb2oOBChI4ZqN2
0D8Bb6EIAwaxM5Look2be3aOQ7JKXtjPZD9mkJOpd0V+kckshsB1eIIxpk8kXLMZVYsmoypMk1CR
JuWTmoXsI1WWivGMc5/2AyraxAQOWOkKSdMvHVVxsM7MeRq9KbHRc0g+hmAglMK6uEvr9gt6C4Nm
uOVZrpfc5LASxeeYilorF/C3ns3YCk8Xio+Ui0EvGrRnoJwE2E9olo+M/r29MxmP6A2HWqm1tVFE
3tnrCkNW4puw98QLw0F7I54ZTIT/buOBvyoHW04x/PokEHecbGIXMWtFhFnUAh6cobNmn5ezkmkM
7y32kJNDP8banhptwo3hi+LKh9ApfrJ851Ewqsu6Hs8z5Ibo+m4u6G2qb3Y9N3Z+sKJgsqnwjfAz
lip1sryATKCcpsEZ4etSKKJ2yNgPUke8Svl+PBDUgjKml7OlB1cjmDKsTbqNFibjkwBfhEhmyHug
G0pJPBAAqd6opyvQfHM0w7jboOeAuhnD5uarRPF1bIut7REw/3LDyfkWit+MZsuhuKUM2IhWmrux
HGqcZfjjMln9Ovqe+BmU4384v/7Sj5QgBwSknOI9ogrY0pkTz0yprDhIwm1eXhNLrJRmczlcguAZ
XgWQif/Ck5JbYWF8JUx6dWPenipT4kCrDECMLCk6oxY9Q2Vln3XTh+BL+jQVOHjE3V34AjSxji6y
NUwsjec39IfmpF7pONiipEsAf3bhmzTeCc+mugNcDDW4cXiy4GFlnsdTnqpkSJfqEaKsMhqmycVr
zBHJftFkH+4mosMr7xMwBRCLNnSs3SZw5u/ncVoehLbTAB0XyLyepwEhELV9bJ7ylAYpHDg5/0D1
tauxDHlvA8v7L48UEr+xOXxk1UY8WuGXPl9K0ssNTb0lhlrBWyQS+m5EvqEBatASA0HNGjAscLBb
K35bnMdX83Va5S3ejPVcGoX3OrQSPaP6C/oJ8NybJlwkq1hsGl3lrE3O+4OxmSj1g+7UP5cxCGg8
6Il/YW9uBxqMa6QJiDy2H2IKrIC9x8X5F38y2Xz96/ejUMBshjup2Trrb+psa0Jigj7kLCg5tpXc
EUmu/JRag7x70ICFbjtek14WZKoFZ2nHtVDzawzv0E4GIxVBjm80XFE4fneNxKiBC0TU2PH9g9h3
pzDZn3PRyXJBWuTCiSpqItBxdb/XuedCoAvX6UiompiqYOGlDWeUO4LXi4TY64JIWlgnJ7v9G4oV
56sRS/0IMXrAS+P3jznOk6UVxOm4vA5KX/vBNW16+/WjZ6ZKicVVEAR3gcK5tJGcekrhONcfSw15
exqsgNA3vHTC10a2g5/H3xhQey7C5umZxyn5bY4T4KhFj6Q6w9Ca5uAqpnX7YgOX/LLeZcloM1OV
Q0s3Qp9N/bRFqufH1kDJmrs+dNQf53AkO/c5AH00oliFIfC8HG9bddIvazwV6gxL1J7o2s5AYSut
m1B+49S5C/FE8bpESAOWAWELIHprVARr7mNsNjtF00a4HBtgFJ0ZhPbWWgE+F8V29GMBPM3IXLkd
4AT4oA+m9YXP/b8/0Qr0ysyN2abUFRjIlNIaiPHDZO5oOlheaGDoNpSTj0McrWCQLGIKSpr0BmB/
8iHOmuSY0YzvWvwg0jNE5Yl5cPMH5f6LheYDMiCfjpFUqobGn87pi5IPiOXD/IE2CzWpqMA6RgK3
Y/ZnGMViUqEZLfXNNuzW76t9Y/A17J3h/jo2tbTp2WDbcDAgWgW9bdVOyjZkYMXOlz912fVL1MtS
DkUkxiuz9NsAvpsqSQdMXM6pIOjSAK7UIFeI0u4xMuAkAV1kTjzrokQ0YTOBsX10ixWMVCjFMzkf
UPr7N510aFbINICbIQzS3ZLb9TuS9IQIFOQb3Rw9+aCtOSw325DtTcCWfqqeKMwpadC2rmbxcY4o
daEM3DCWKkBrNh9bc7Uz129sJYvjdFpguGJdxGkkf6hddMabvrMrDwqcI4PERZtoXG+QOOt56gNm
Wpsc6Ylqn33YGi4piUu6shXiWD2GWAPXI4stK+tdHAoD7KG/DOzHlXL/FfyUW3mJ0ku3FyuaqR69
z0Gm64Vrp6/Gm3I5bqPXDEsvR+xfVEvq05Q0bfHyVdqEd54c4NXMqCj5T/l81p+E9lwwI8fXb65B
m1MgWpb5R/0MN7sAUsNSYN2ePRORr4P8GWr0f10AwkohObWnyj4l5iQ6OfzhRvT+p7Q3SUN4Dj/M
yFDRHbF2jWmBVbl2mnxBoj1b7LOYGlGtJ+56nQdTir8XGjnviW++o51wZu5g+bnJ/KBLgthWuP+V
EjCVBZHDKHTbzRJKUUhomrkonUXfhMnHm6qb01L1csJAuTVrivS9NhG+rybLk1VfknE7SAx/wuet
6D/LyRQAB1pNFwo/q4N3lL5/YguSeJamoJaVcWS3A+Qr27/27DTkxuNDcomCdjESbvRwXG3oVkM/
2vC3ZgAdsq580gSJdpLCmZvI+VjYsp4uZa3+M7imnaeErR+NA+EDVcUAVmdnp0QWtw7IMHqn4mB5
7DVHqxH+4WIQrl7H3JKguKcnIt9sB3Hlx1/J7lIgus0jop3X1fAa5gL/Ky7yCAzSHtb5TMxEBCwB
bspmufck2cKWGiMFhdMxtajAVMI6nPpXvOQvGoXYZjog0UGK5SxrkKNewUuaKc/degdZwswP3w+i
nZrmlzO0lekQ16TuiAJ0ZRnNim9b/nYX3IM323VQAeA+IUGvsLKYMKslzjZEeCtAcg4Dof6SSK7J
Ww0YCtlmq6H65sHMxRj+qqFs3Zt8BZf0fKUpOtphINbIRTTfFAzRpqPK/qyBSAj0ktwgZMOxQ9BE
zNZR3dzFAL9Klp1U/kSpeNaeKwxjVbkSbsBk3/N3RmJdxYKuyoAsQzpmdMW3WoxOWo8uBEVCff6f
O9O/lHHllzymkynpjpMq95Zb5/Up/5X0/HfTbSw0ftXELc66HziGExeB5hdPcsu/pH+Tt3kpiy+O
sUDXp5VYDy5onnJYHgRlNrDwoGbNjGyBCdSgAA8iganI39WMfKjrNMCgFM0hmeNKjpUwdZmUSxRN
w906fTn+zBIhgv2vpZF2yAG5FejTKv8honEQMG9pD0MEGWwubO/WxapdR2kf2PoW1d6g50+YNzRa
hKkEIH2o7yG+vVa3I0n9wz4HTgjpw50+C1JCyBspgmbZEr8lOmtWuYSKg7IbcNnLIxjMGrc481FQ
3D2pjvDh2bpozkYe4Huy1jOLcCqSXZtMUhgdAeqF4el8h6etE4/qNTeSqY0qqfjhhPythKI5LizA
MthPWX3KyGHCKBnLTZokCgdRQPm3CT0OYn7FNIoQme3I6opNfrPXuONq7qKTuR6xlWeBhtBKH/8B
EH1hxcwtMH34DhZFmmvV35zjSMIbi2UoYe+z4he5cdT5JqudCQz43Gq7KPqKPyua1SBdva68FCZf
ncDfQ7950ryxQ7BkajsQW+pj/xbDjhAeh7dVpBth5fYx7hdMeWu+epLAmJt8Cup3PEql0TrFZq7K
vxttZ+yqwy+svDm2Py2tm7abInr8DYS4iTKyHotRjg+rwtJqz1Xpy9xXxnwX2SBhQUtRjXqsB36G
GBiZm9l5kgNdSWjlBF9B2ksGCEwi5bwNs7C5jBlUO9E2Ox0EIsW7ryCT/0zO9Cz4Vst38fzQVg3G
E+1G6aMkuiwtxGuNgYghF8POHgsJlSDWyHAEZGgfkoX3t8/q6gvhWuhoVd2PMdaQCD0jho/ShQI5
jtQ6wVdBQrSTJkx2JsKXVEu+geQWDR307cXs88nRAMdkCx/Lw/OiHT9F49pQU5bi/dag6elUoeQv
Wmqsr4dRJRLbdJJCCprb6QmN9Y19MDxYcCZJlO2QRxsmhlr+28yzf6DEBkRlywKkN4qM9ZWumeOI
EiTIcx14k3nirJFJfXjmmP0SDdjeUJIUs7B08ke3qUPfSOs8mKGB1UvoWEKicJC5ZJgTXytodwU8
WEVwX9T9DDZuos2EGV+JDbFRx8e49CiqNd8SZ8B9aI8wTqAOq33K1VNL7jcqToBnM3u7VtFzuwgK
4sZq1CDenjjrZoLpJEhe3vzu8eFEH/aeNlUnxxjgHpBqSIHXFw+9HDpqPQ5/6BrMeSLAfgIgt4s6
RZwUGelqW6L+m2OO70ubC+UETiTp4r/cqWk1cwVfiMy3BIK28CyPkDr1RuaL3/nFJ62VDDZalwUz
5VMdcWlwSc+TiZm/xEYbFnN0/xT31NdEdQ6t1Re3NyKi7P1hubedl8h8jQpYpdtYrAiIs7C1bTEG
l417KEHsmOXuzizESsjxsNdxo1lNpsQRmIr4aKriwfNQibGgBySaYyY9yDbe+zEQlJE2CNnGk8Hp
n+2/oUnJoMx11m+ukJU/Bwj6X8zUIiX7gQCo0Lp0SXMgOWfbe82QKkyaCpM5qzV5j6VvE5A+Hy6p
Kg1AYT96VQxB09GnlVhellT2sqXSFUoIHT6ew26hSZEB+XR5FE8W+88KoyBVIaO9s3FMN7SuYqXw
AH0Sm6CDA7eJ+9fYU61o39xIzuB0mf3oH5oLjUeqIgnmLTqlA2sI7xdjpdKIVXppUbWfnyW0wRRo
RHKOzgpMmUpZ9ZwSEtt0RExs15XfRDSEPLbIMsysCnn7cHFjg0cosoq/KJZo8WhmCkcnYlA5ZEhH
v/TP7WhiRR6AChC4t4wYkne/UyD4Yfigja9XTNnvnpGwGcz6zpsCrrcwe/DyS0my+iWLW4lwh1Ak
0G+eTFZOb8jRakSZO7buzEM9tAIm5aL/b2mGZg5Cf2rhlI652lQsUX+U+y6pPBUHLbot9P4xSV5D
i0UCioVphmBoBXFmWlujhTp5YtRBjF2S5CsxZhPuX2ga6DH+p/6eaOrD1M7T1c5A1pG3gxTyRfXe
ELLzgE8ztBC16PqYD1BRS/A5S09cP9cINLskusC8bPYJCbdEg4bvQPQh/2Uw1f0nOjwS4clwsj46
906AX17bIMIMbXbuw3vkG9yJgCAKVTmnLvAVYbk9sTjVWkMrgQwH7h44RM0KepLSXjdMx46kp5Nh
Q/fyJCTT87LlKyaTcUvFFXUy6kXL35B6olqd8E+dt4AlqiddofzmE5fI3upcKaXNGfFDYaAwOH8J
SYlt1yVI7fdG90+99n57tzkK2qBhWiJpoIJt67eJKJYgp2U5vjJRjho9bxzYQAC60l/xleX677qt
HRR0UKOabPWqdPJue0FvCw60P88i2TYzxmbxs8lwSZDz06eJKgwPwauQdkgr9x4JIPnHneieCrXK
0h7LHwmudQFZAh82KgQHqDOcHC2nM0jIgNtzr4z0+BjocgfT7x0Yar63017DbICJ8w4OoPj9opbr
KT1jCvoZzI3ViwwmJRm3MZWSKrol5GtSiN61zafBYKIDQXbTneOjJXMe2oV0ZglzyEHVAa/fg9hG
+KrhC2Gt7bPsgNlnZ+u+18WlRul8MwhLbueZGcd+FGowsTh6k4ElixB4pA0XTYivoN4YtQa5OIdD
9xzgjJ9Ai9QoSOjIqzelHMWeiNr0XWxHccrjV7kjmUDQkP4+aEn2Tc2LzQyKPxl2nAB5hUUalhyQ
+XFBbF1kCGqq8uYYEFGXGC11Lw51hCABhejiWhBVuyb4/FHpfkVqJR6EU8U9bWrq6TrWMOT53Lo7
SCLPSS8Db29AZqDfwvRSOInLzpbHigLibi0Gn8ikXGhSNwWBluKFxMbwUJzJrDFaf1G1H84pKncW
/Cvgo9cqDrDHmlrNS5wWYW/ZL9JQqZd5HYNxqtkEB05udVmAHz8lWKddUi0DZelf9NEz13wXWoXt
VgZ2mWFFpnbeOK1Quo8E8mwW4hucFfUTcUZLgsE1otMbBIphgspWlmfCAQzCtCXu1uSt90lxMrKR
VCiT4DTVJ3fKC8vNR/EqTQQM/fTIpjhQV6+9chECxTXgr4iIjm7eHC9lMNN8/QB9wiLBCiHK8y5Z
UKUcW9wwRpgxsfB1rdLShseNCzKk7B82Nwgks89Abn/rfuRW9NiymfRXoxi5LofSSWiUWh+eRqOh
r5WIAs9ma8zwJ6B7Tr7TihyPo8sCTebnc57PTqWpXsz9t1m6AVqdmOED03eu+jQBoQ1rneHKgjms
SnB8LPmBJP7A3GHPun8rLYqPC+mQWrGcZJ4Pb9Q2eh8ChrnGnMgjT2e5MpACGkkIC1604eC6StWS
kdTuYumOkCvy1qSZMCeWxb15K6nOgbCnCDFlHRMU3B88fjwsn+wxVjPgtwzDtgfGoTTXwpC7TZrd
yi1GCngtHB2iuHI9faesqNyhn1cqzn7tFgpiPArkGAnp9Hc1RncSE0/nfMBOCyCghoYOxSKIekc5
gWRUDGVxF+b9EXjiU+5OKN5p6ZrdkhvIi9dByPChZGo1kySbwGLiNb8xeeGbFmX1OJbxOtJSTchP
PExoyu1jdZS+XYxQpGKtlOzSuiqpl24zgj0SuK/rZV7F5YbB+8EdoZBJ9ATgzNUQEp5m8q2JWFmt
cnzitIZzgVnN+tfSCQ+RxSCAIgWgxTf3fUAUtVJzytkyM0mosqms/FouID9vNp4F2tMIey9MAyfY
KAcnKHPzUylzaoeUZA4hBd7warMK7j4Msc5U0wA4ulECDhXjdOEAdUYQkhP4G+LsdWx/YF4Qjz9S
7aRhcVdI9FWtzt7iitvVpNqPiNk3LG0hAgN9LBBdgQbGdmSrzcg4ry7nHNiAGk0l2otiuil3VXo1
ElPDNs36rXbPxeKKsZTpf6wFAUyXepBXPmac8Qad7HkLFHP6+BpYW84j4GeMiIZx3ZF365vzJUAM
eNO2KhOepMKc4+QSyOD3bo/JCi5piBdlVGKXxcgMXYzgKAGJWDp8/KVP/9RhRtxmceAGdY8+vclA
qv88OwenxbUtYP2lyhGPznibvfGEVRTKYirL4rjLYv38Lk2Sxp/08gdoKZV0AFseK3wwVSp7pgT+
QK58soJwfiT29ULxWHdJQAU0BGuocKHnl1/xEYi92UXpGj+w9ZN9zz8gOKQKMez74r5K4p6Z9G6o
Xkl53nleexIG2bcQRevUkGE2xaZ4SCONKYGPCpCuRKa05CVGC9uky53G6aCJqSB/hoKDuKr6edtv
k4kn5USbkG5COWzH/uTshMrirNdlP8zEBOapmTCPX5Lb9RlOXi05W8Ez3WkWW9aHOLymvsJ/fOzb
aMuYlYLiVX6QDBXJjwzTbnlFXgMoTEuj4dNQ2oNFt485qAOG5fgjKfWsagipsrT+bCl0FTnXZuQV
Da5BMArHFXJ6WsQ9utYi3DDcKBVBJbnwIa50scua5mfZ8/MK0mqZh1y+d6VN3Y8MY4+9ObSYkbp/
1zxNrsXrpiaqkWWW3jnGJqAR40Ugq+CFMR/vmRInZoXe/9/Mi7nh5Cy6gMFdoDjyCGKybl6+0E80
KZxo84e1VQBOxtnzvzLGaMUd2g/qPrHOHU7oXKtcnn9AHx+5o6Fq+OzXI3yi7b9EJ1qwFxOqiCCH
BzGh4yYK8JfDs17GHIs9WaACRCB5qK01kGUjLs/LwdMjb2RC8Fd1bqB7Bi+dYfpOn+Xksd4RWRer
iwze5i2mQqM4BSzvrVOMfLetJDkz+kwxKIPEGLjLENxacqthI7GKDB1wh6aRvsV1IY8Nws4n4i+7
okrfKZRC9U5NDD+szSwks3s5dzI4eKnNFRlfvsYC6a1tZtswuOrr+TCjracC+syoX1ubwnHMLuso
bwyne3AT3FPNaunuYzchdbdI7zfwMa9hyGxXK6trhUvvUgM2Uyx6xnvF8o6HAQmNCmHU3p2AeQtG
uMxaJbfVEFlfORCY/FbuyFm0p1qadIpjZdb3bFaskZXWBhlstaJ///8/7qht/rlepPAaB2//BBJ7
RC9hFgRoVbkbDnMAAvADkY09yU2qnmhqJPLlKzglpXF+xI6NzAq4Pwp+QsVANUv6lUNqKa33PaFm
oU2Locz2ImaeD6m9uS98p/+SX1vlrWA7dl6IQUvSoZDccblk7NBYkCL6DsvWWnRTCRlB6JZ/7Hp/
4vpueiOfM7HmqD+4UkpGRTcSz4oxeHco/ETXfZmH96SKNuvpY2Y5UQD15ANmeZhNcBoYEa1KLNSK
IdBtXwvI7afXirlJKq2MzNJIN3QxHkcklQWZ2yZAAdEr71TF7vBDjm35dddDwqkXH5gkcDmG6xJ+
kKfzuqVdMPP4DqCNoCMZYK4tg1anRYLTebLGslCrGqemspHGoivc3Q0kRo1dOfs+3WIMcDhqTKeF
4WLUQ/GEsOe03Hutqy7LyRUwvRH3gAWIdZyGGtPmuB7cMVo1iPYgm0mVjdYu+wGhmamke4Ws8Dm5
6NGEzfcgnsbtDCN3nlzLMbdVnNb4nQ+YAH0tE7DlmQdBeidhShOny7z0yCQSqRGzGtpg5knnKafb
SLerhyMY5hWOLRcHby86J9wixxCaUS3PobVgbBinnf3bX+BY0NNQivjjkbzYu63YY/SvNJ2DBkPh
9XeCYJq52imPHfkvbgnF7sc6aVQCFXG1fwStWkPp1z19ZlGGMRFyhGdagFKmDzLCXAjvnZOQD8nB
wG6Azp/Xbc4C+QmdGttb1ySrFDIA42r8djA3oXhlotInXVL+qvzcZo9qXS06sB6hGEB2+gM6IGHE
9JLLmWG7+oxYeogbdd4F8k7hlVhlrNiLXObiVbrgZdQN++2/FAKBHbs8PAg1uPuRyQgur8ttd9Ab
k7mQIDzD3QruJu/6pnr/4AFA+TTLxXflh/HzTLHfS3jcyDvxBXmG+6MLdNClefqzM7w51OqMBbFI
NMy8zzY1SVQbThjKB1YQi3fc/7Rk670Qde1Mw7Mf33AQ1XIJ460w57uyfwkohlyGS84fnpSzqUGj
edDVhIMo508H8XuzA0I5a6/rkPnXYLw3WCl0LM+SzYwBLWcCZVaQxukD9Q3lwQzc8xNyqhs8ohfb
WDblKnMchxckeiihGR3XGqv1VI9aKNIqgxPGEZxR4d7aoqZwmDkV8oj2W7DqeHpxw3IJJTG1GRo7
Z6n0XnElbGhdmAgv6OktBB5F74FXymj/DDUUA88mdMdsL6MucQV9zBxxSNTcSupmEzeNmPczjlWg
rxx90bknJa//pTPmvCxzqVStRMo2VftzFCGTwmhit623XwWj/LtbKdQ1nHIwC+bttrvX7TlJfT9g
ZwbypffMx4LbTmMPaUrudNe6U8WoOLxQ1f6ni0Eu6SGWxMR8OIc0Ili5ciZ2n2564pYsC3iYLHdO
s//UGse3+5j6Ju05jviTR1I8OdVieWbtx3nbz8tN4qwX+3c1JUOjcbAFlKewNCho0HG6a5vMB1hN
TEhEzczXvdQAWxsDpNo69vxTu5S66lcPoLVNtJ+tzxaMvq2cmfYmBpwzrZx1i33I7xoB/P0oYxGd
yox/+I2uUJ4js/fX8e3HCDom7UOJY86P1wHYhPS+ovBLvYuSo1VFhJdMAnMY/EkSYPZcjn9EEjZO
WgXvAnkYLGna+rmmCfgRRidhNfUIOXpu/KmFh26XbyCMblvTljfsuNJX4hOW9/cOoFLz/04Rf4AH
0kRtn0Mu6FOk0Bt5Qk4+rOkfKnsJEyjbaWZWab7aNCmuCLsKC8fh2kQEQ7DIzYkMwaHhxqhNidZq
uo0mz0jDU+Zin61w2dTISrTGhSwXoJh5UZvF68rNi/mtwERHVNV1jH6Fc/hyElFJx59cr4FFXoPd
g6ODpvgRdgF+YLjh/fM+3K11uQdqXgn0E8lOUmp8Miq+wgjW8ZuoXhXn1GVopBRVk4DCdxF0AKcQ
HeQ7tix39jMaD3lk07Amxf1hEcmpaP16WvCodrPNlFlcz74RDjua8+taqFirMUmRHM2R5116u0sr
zUjJ6DNTvOwoy93ymDzv22CaAQHc62z3K0YFWS2jH3q3jHK+yuqaqPr08FQ/DVOmNyEz1pQNNjkO
ebCAhkh/IIeYRHJd2jGXsij7LCwxKA7byj2n0MsPD8Hs+ZaMVzRL2QkiVPLfLOHRGaL9/nSjl/Us
VjNP76UXd8bTAwdXXZV7/Mt+Z43Rxa43vi7On6OaBADmfE8s8e8zjnJJH3gpDZyeTBoGI9bv4TJ1
nkFb+eZPFrnb++SV3OKj7hT11RwlFGZ6E47GUkCAsKrTce7HzpkChjGuufQNkKQE0wh/NiiJpcUq
NEA659tfkGacSCR0GzzAMEowHe+ewfnBDv6UCFyCA5DlaBeM3ycNFTX45ZBf8LCTQkZXyB//Km3c
g4jl3ofMlHb8Lg/aJXHsOUcYQGxH2gGqLed03Gvl1v61cJr569BrGI5p1h7I/rmqEXK1JuiJYlH2
zZVlw4boxeHuyfH7sFhTahVoC5LZFPiftl3V4CStT3ahZiHdsY1mlLkEG260wTIdf+bNK/mh2TQf
rOwVtVKvBlNY51ni15zmdB/3XLzYJOsBmtxd3Y4k2hi5MGv0NX/Sohv0AC+RFPhLQIUbCcVxukqN
0XaqcfYUAvqHJ7VB48xdP7aF+XuV4VIgHQeo4s0GXpNN//wn58is/dufYj3/kiumvZhJs9PbxjL0
ckDAOC0UnHeX7y8QNRTNGMUegDOKUn0cELmiiIZY037cvAE2U9ax+aiB3v3J3yoTHL8YIC996y0o
Gwq165ftWHVYWy+Zaa+5MJ0OFPAIOf+yp+Rhot57027Ex94/Pm5v7dQF7JZwlrh5GA9S6GGZcFYW
j4nK/PamuT29jnM1I8cPa0+wlFNbyoL5tvvcgVo2jIzizTvAJEA4oKCDS06KGxe2uyBLnTrO1EpY
hBTPbORiMQdgDjNKrWJhnEv9/dYChAQTLhG7EYWZf+Uw7IVCWrGcCOZKDUg4e0rHnnjw84CXQ378
3YWNWtSHoAXEeEhsmQRZLat3PFzJlLDA+wY/AYWSrS6X2DJQsCVEmZWJvmQ6/9eauCLKXLr6pgT1
tH2T2zZp8C4Sy7tlQF+Ea6t9VrDFhq1c/F8qySgZTHhGMb+YkA7QJS7l+OSVL5D1cJArrXtigDZ4
Wedy3OMvIARd6bqHfT7yVIdUCG3GIw2MZDOaySpDVt/W6d/5Gv0KPUogD3E6fuBaUdmvkVjD2n/R
8hJzYlgrf3ZGIArBL3PMvAads60eVikiVRFJRr7xrG97ZgZNc5uU9LWytGUOuzB3hPi4wUdXJZY/
JgUhBBXY52qEK8kPomBg1m6EW64Z4UPmcPraE3lHuX6kPHF7cet9IMR/PULbcoV0eFx0AKKr4ClH
M9QOvx/IzUYLmecgmRgGuLd5GOEzAOFtjTsgTsI5fLlluwvMO4KvfHX+fqqphyQotrvrqgDNaOfP
pdE8E5AnLsXdGPAqgeG7U9ucW6KgNrrO0NV+U2kzO5a4yibaMZrHA4V8BQZOl1hcr6IcDuhny41b
t3GVE9Xqp/duTj+pYsOdqQlrnyYRnH61yGScIpHm18Bx24nlJruky8ZLNBTeMBaGMSCA493E6YtF
bdyYejHP9cSd2CUcP+uq9/UhdeGd07Xu7PRD5K5rHeTc84i6p2+UsabtJfFwdZ3W94G0IW8B7RX0
hIJgzqftHIq5q3vuztN0400mL4WkVVpBKeDeYSYF9xwwtyfVIEYWw5UlFgQhrAdiLRvnHViXUeY2
8UQC0WkjCSPMgdczkSebwI+VQ2JxjwK6jzlj2cGcpZ1boPWlxH2Skf59pyx3/Saqidg8UvgvZDyC
BdUTapkNy7y55wuTY+BL0sPnjXFbuTeZrW5WFPm4NufzSApzvcFwa0vPaAaCxHxwr0OQemYRL/gw
ZtuE/WnT088wIq92rzeFXLDemwI/sOTS41QggLBNYp3MemmuI7j4KpU+xkbWtdKyHskpD5TNih/J
7dWdI7363ncznObK1XynA6AQH5lAkwgD93YdBhrUauFYZd94JI1R1hQuusjEXbt5/Q9mpk2jWgZX
DdODlWhJHMvGiGpaVb0sPjuOXCp1RNY88C8ifWpZglp8G3rMSaBX+GsEJDTfn47i5IchMGUDzV61
p5YkWX6JVpnH2md6K/gd3x48MAPycADAehZEfojQUj1HZAnZjc6ARBk0yyuo0mHhS+wIvHbcySXj
clS7JzwJznT4AuTsLYxbN+8sxOQ0YKOhZzvlmdCG4OJvMA3Z7PvJIYYOofm4ZWMI4HnsIrISnXqF
VXR6ytEBk/4vkDnsdEQ31FRgCCHgPKqkv1h9UJEPoUIDGh1wCck5+fsPYQ9BfWAENHwwG64p0/Kp
wEj/NCMOjo+q4yeHisI39g31xfk8fr2IVS2QYMbPki6PKYHWeF1RA2JP4DZR9WBkMHqFVqiMxMro
rjmrNyJ2bzdvAnZzGIzqq/FQDjkzZ6ACduGDbIiyzC+CRKRvE24S1DmW4JV2wH93bI2fHeSNEesF
AAzWNYJRSOjeu+w09G7uAjqmjrVC3zZTaX/kaLD7peOe+JAc2r3R8FXoLKSdbhnBCoHqMtFOh+dB
brP/X2nD4vlKSJAArGHmQLCPkuW2iNN2JqfVgWS9XfZvZ8HJblhDet7tbJdfN6JZuRwCOuvPwF6Y
ljlYIY8dYqEts5AmhbzOuzb0Mq/j4QC7FGNWqZdIGQHek/vIZsCpWrMDWzjv7mxXarbI3kUquEsK
8HGL1jJvMLFr/6vbdlj7ORTq51BpWw3sjpf/wWRmCkQJlKiBLKb/BL2wvTKU9XMyOs72XOnjfFhG
QsgDGMPI7Xixd79vbER3idkXeJFR+v82Jr1NTIeyVJaKXhNnKcQa+0sEQbnVB7O+3xELyDiGu0v9
fzWXeV72GkYagdaoVTfDvLR8C7oVTfqJYh+eDzhuEHn3B4zQNu/Hz5NYMphkGgtu1VgvbqNLMP2j
5E9T2Pt0BuL/65VgBQYjNcX2Y95RCS6bjCUVN3cXyT+vDdLMbBNpOuduheu9dkNNbF4iUPFHCwLP
Whb2DfDWwZfMljW2D19CBoYJZgxx1CKsl8ErFTl6xvOeitHKy7Z39+zXjqav/ODNxL0A0XwXQMBr
90rp7jIShgwaex5dm5LFuH1ElQTDXzvGqeL1SOlN40z5cVqG3I9ipzy5lgwPeLhITq2x1WiQlwwJ
mvSPKKQZnqepy6zTkVC6t+8p9A/NegkiQm31jmemMxrHD0Ew1YgV3y2g6BpScx46ghwmfurAHmDW
+xpt2VcaF4WR6AxLh9lXkBF0s7vhsOTABGsQ8P1AeBdyBQQEuA45jfg5YFdjIYULfJxN9OBBCCE+
9Af1DCs1SFUdEh7OLn8R089RYhr8MEzbZTtmTQbHqhrPGsYdPpz9OKIIL8Bc4Pr4dHjzxPs7FWBG
PfXAWm9glY3L9uuoWc0+JArVNZD7PUqsmbPPhik5iAvVEe0eTPS2wzDHNVWIJj9Uk0pN7ym6cuaQ
xKmuCaXqyBiH3a8kHHXilfmV5WSe1h/+W9tXsc3yAGSC+iF5CtDO4GgEPK6g5UY6cM9qpgAmBkQk
gxsOjl43LoeVXhWmnXgZwYH1bT/iGArnxy82KvmmhjELyUNMTckA9ScyVgB22w+mTOVSvTpjYyiB
cdyF3x1WnskVqADRcm8XW3BwS02YppYZPNyzf6FIqxkRLXz9fHbJlruKaZrfg+ngZlRUtXO7869r
651H3OgH95YXuB34Q2isVCZCZwTVZDh0NSHo9dh9iNKWkDvMsd1tXovFq502n3uqx8vl+26idkcy
eeRuHX5r1cHAeNjJlPbobH+IPUm3BJ9JcdAt6y4YGzQq7JQFSEijPIfIi1wHST1ALb/ZOL9A/8jk
lOYIk4i888B4UqgrJKx3aqL3G8VcenGzMSKvz8i+E4dHa62qYfCVL0IKEB7oglFTjE6vFtUAt19Q
sRNfQDXgNquVON9EEuRHhLO960bytl6IZXdboHCuKvjZ6top0YcQv9UbUsf8/0l53YlWNCh4aUh9
/NM1eY60BcyG6U7OhY16PY6lzKX1BFlZv62qDvQChC/qAuNkDTPYTVKI5TzXLkLmCH6Ip32svQsH
p2BTot6KIfPC55xP68wjvvmwVCPB0nXTXeJ/uho4bKMQkBP0vmV1emh6jMC4dIlI8CTuRWwhSl+5
SfrKMgLgFbeEm5WRSW+Si8Ks90dI81FPy+Tt+dxKLGXVztti5GT/5Fl5voV/MR4yt3sUpi4GwboL
CAyqEvMs3Ila30oByGRwQfhQ656SD/ovSNgZ1Zx7REReRG3kyeEOrZU9CxaXoYucwn7q1Q3tZEHT
GMsTxWmMjxRX/XLcMetuNwxiRH6GPfn3fke6Y9gexCDYuGqAfooCzZopANpj1PcnjBE8hOKCZtbQ
mhe294hONufvylDnzLR83/z8BAYMlGIs3rRpzYDh7aiVX0S8uO1ZFiUpDVG+50Tc/tpI0C7ZvW5R
AMh9UeJXsnaXRgqho7mfRKTYdQTN1UJOnTPU0DC0ys8EMEhbJfBL5iBV9SLvRWvEiXGpZE494g8q
ku6dngs3ctysVEiY688fKlLrH6QOReYbZ4C50/DmSdfRq+eiSkbK9Ifo1beLHYpArG5PsPfBsKqN
qlsRPjG14Z/6FRHN3syIqLlxACurHqtdZricHvsskOe8mQPgj5u41uNFKaDHSB5WNz3NqF5aqiVo
aW957rH1yOjikve21XD1GxjkImuRMxJ/XuRDvxkDXFoJMsT+Fu2dbwXFDuqlRaH5+hK0rSZvBJqg
MYvvzAGy8+n5ZSiFGQ4/4FRSYtnfTEfmVkIEKD4mGijl/UvtYwiRc0//s+klwSTHRnLwf5L4EaAI
CYPuNA/fqLRU78V6pf3jbH383zOUkXw7fVdyZ2lYfQwW6NL127N2RFhpoSc8q6+/zrdc5XgmOQZM
EUF8tRp6J2DsaPEKigwEtiqYY4WX8UlThZWmaCQVpJeFu7ytkusQNdQ1F+JQBdnGeKEG+GqclIJL
UONJy2PbH03EcForK/dvzCEoQuW3TUvRlc3pCr9pLZiouzfgqlCO0wx6yrrl1LktXjIyhXjgEvIk
Ghv7vORqv5RiHWwD9rbGJtBe/ePG6wmAeJuoxFAfKi3Pnwp3xBK4/2t5w+EyiWx0XUPeqw0J70UR
ygWm7e8h91fEje6rmummNBwwlQRa7n1MBJ3UcFFIWS0YcpDzNIovBpYFhreTYSQJ+ZZX+B24ZUO2
il//NuKoI2WyzSU2RzzCO0HOYFljtX6qj9hiNCOouL6KFWNSKHvnyHJIXQK4jrByQAEXpw+FSPZz
CEgUfNSUATdMqqp/rEYYsL/reMoOpnGCjUsulgWIlLyhSfTSgSd71Aszh15xVvdLGJnuNg8goC3p
2IDQpuIZY+ZFV/Axj0G8KZ5MOTZi3LoQAbVhEnC8U+zZKbJfcs8xxAKO1vT79m1zJo0TRYgyC49R
TSuCADQruHmCupPcVItw4g9MNHebrNDIyHdsitX7T9y1f0F83XdDM1lQgf8Fc061/dWj0CWF+TBP
lO1d53bs+FdWHlDONhhr+t+0Mpv3ONi+XYDTcb59HoSyGORPZoYFRTPQ+r2iDwMhHo/gt1t6q/Vp
nZZimeUu/JzPpGBMJAPTZ/WsiVf9UyP4Y7b13KllYwu5pMiwaiSjWlR89KPwkGESYsFZNgyabii0
FLZ/0qlA8V6XJIaWlZW0W5koVCbUxw5TP73+/eDn4DH0EH7C8ulzy7JFgzOCcUjVn7DRUqXPV3dU
nNlpcyRkHexOSNkazecJgdgth7Nt56tEmvxhN9T6H3nXgagCZaClxLphd4CRBI3Wtam3YOAf7hd5
gpPgJb7RBGnzmoVZXlCsuPaZIa3p14P1vq8YjsDLLks76eIvdh4Ua7uiVBTYrU/uQ/di0K3Mm6PF
abXV5jFTuzJv2m2ESOpCniJkcp8di3N5gtNzbYUinGpEf2TQHLoZz5WiuXcG+Ee7gP6w9uFBgLOk
a1C78sfqsnqMY9gXwaJyPSumaVveHFsMjXFgaVU50eipT0nENZRBk2NaJraoSHWkFA/+ykq+UVFG
1e6FdoeFG3qW3QgR8V1vS6OSBYAu4qeNkEqgojzkHo9gwn+2SNC1k6IwFM8BHqw99wQp4ITj/tzB
lYjfVyfgmPm1i4hBtKL6ipREXHnnP+dVvXN29KY7VpmvOYerjlTDO7fHshVzzkvNxIKHIJsNiPG2
VhKykQ9/vMKY7bU3cYc5yqrDUOsbR3CUOVQqTXGBJ5YMEuX8O+C7SIXjUKfwmnLSTHgOzoHnxZ0a
O3IMNlsYJWOTnbgPdBJqATH+QFYAyKH9trngSC6mNY/8+VG5URJyWodvexl23D2rDOfdnRAvJGOG
2J4+mRtmfBwyHQvO0sL9+Jzdv3xics5mQSmuaZ2lZ5XtLkQu5CL+gG4965Zw1ABMrcyvJhT/8hMo
YaYcz8i2EvPKIa9Y6BH6XT/KcHbJVhYPllg1zEy1uER/uiLTpQNPaIYPQdTp7Y+nI+ye9rTD+qHp
AAHzLWSkX1E2hEg0+wzG0jJKodc/+v0pRKcr3By2R8wZ1iNL+XpQ/9Xg/MtSE/95+eXRmslC9yIg
73mZObc6pI0ssZsfoAUiIaAY4F9MvkvYhkqTvFDZdwbLf1nzwvgk4K4hv558rroV3C/0pteKuxlC
gPMcU/LzOtqko7khR1xKmWGlSGlxNknUq8Dd2GYzgQG8ftRpi5qis0lTydZivr1LEVEl6L4+PChd
gD/9uEIUHyLs6fJcbpJ7If02NGcQdqF/FWF/wL0JMs1AKDdCh2vRLGRP0rMAwm5AcPYIgPoIIUB6
/AUyQRqd0V5ku/sbB7hXFX9HGs0oJfswdCt7YhPszIe+aCwXou3Kn29DxriVY0uj+3YXBcGYWyAj
4dQ4GkEwIN8FyPvQr6wLhZtprcQ58B+n92MwTIj/1TQ2VKtTwWrMfTsNGWEgvXDVjnarGhkiBfYv
uADs54eMl83bshtidkPYyr0zjdZ1cYYNu8Vmq399hyKo/UVoX/8PCGG+Yo9WhKNx7HLhLG3lf9kw
k/kMOzLOLJPKYpeEJ7wZjIn7L/1N0FYbz1ccdjSqcJ1T+J87UC9VElsELNXzk9STJABdkBPqGuly
1mxTQL84Lt/g1TJJneusqRx8Pn107f4+mc5HM+cOneknHcHRoE4lTBp8c3fc+wKTOBnoKvYAT9A/
khNNYPfm2zjiT7TsMJy9e3BJDyi/bvV971WFP5Cm0Jcgeom3HMjDXYNRG5ewu7YGuGWZ4BQxxAKL
TGUjG2Xmb/+DQYm/Y2oYV/hE6uJyNLy3cwtW8AkFkgFXcSmmAgq1LiONJcVyakKGoziDmd97wCEA
NeqZx7VcAyMDAhhan5KzdIMUhWqy2UuuABE2L3EJ7pJrZPiuXzSvpnQ4D/fSG65L+hjrXkZJI1m8
5PwNHHxBCtjGf0MAqpxHoohH6dwwLUnA/1cHVNXAVAkAnldqH1jKJHE6q9HZzvl/j8b+gNApJ37o
5kkfDNf4skATSparUAC39LO0LM5kCiTa5LFgWwwRk8rD0enn4gqnRp5hDb9EojGAxam1e6btrsxX
mh0TEwWkosml6RX/C/Zcc75KJP7PDvL3ay0pEg/p5cjgErG1xGipx84mn3JvTiDAomdmSK37hi6R
1lly0WMam8hyvkJubKwh20Dk6veVExdu4qRGwpQPjVlMjeJp8W0ucA+Ih7+4vQy+1tKm4P1DAomp
wdnAXjbf/SEnnJOPI8QfKHQ5kQlyYm0/M64g/V53PmvEIpalDEpVC+OBfyzimb5f05Tf5Gvew83s
tZZ5V8MDSD+jeQBtaAY66kFyhwwqDtGm9gVVlm7eblNYLwKHXpzbABu+nOfoIyQ4lH2e+JO7mdli
bwP7575jjIOhzPuAMEjaJR0qk355M5sq+Hb1Ppaf3mL3LDtB7cwNBuxNqUVpYhFzVpJwKGRfnVsS
GNBx3E9kH/TPpzFt9xO7tRicDkiKLDGqPTgUNh5CAGTe039YrccS0cvUIkq0lVigygIUfhyIKUaD
Kvp2r8s3wxGqbLAkp+jWS8oMxU0LnI7I4y1ZbjSXy+OZCIUeCcRjCMsckMm45AXAtFlmbBGObEU3
+Yx1d8AJIKxla1WJtWagbuDeYGsDo3T2w9IQzVGYBEegVMtCX512+7g0WUaALZo5zS/BOY4sEBA7
R9eZPuXBBdkEq85M6xl7Wr3hZGquw+6dDZpT9nbrT/FiuWd1b1zk/gfkqTXFZKaB3DZkzgZAvS8Y
c+ACrCYmtyMcScxpHmoXLsNMiwz4DpNxdGqwhfhC8c2GYV/dQyj5w2200E3zqFZ4elTf479sfc82
RrfRwi9hgmj+PGfXbmvgDEhZK7lBbMsTrMLYNlOMjIX0+SKoD8l8j1s2kluTmQFEf1RYUdwdbmHx
nxgkvz8dYIRQLNop03SZN5ifQ04+7BhKp1v6iV9YYdckP10teqiYgPViUL01FsfbKaJ0c1kCfJ6P
X1KbX3XNm4uc+A2Y561E9CpK3kRda1TFLTGnAcaAMiNS/f1ouC6DSvTC/H94gMrHvv38OFNNM07+
ga4jH3+FnNNj8+YLU07n3CoCtbkM2anINDDmq88pny33s0DMVGirVucDz6IgBzEdx9C6q4Sl+Yst
+PNkFGUX8eLaPrQdMh5V1xEUG78/Z9nTZFNdv637osFFlm3nASK42BYvSOHaCIcUI7zrFOzxbORU
XEGI27kVzGzqPsjel4PLWqbN/WgYUSBeMLb8NhtmJ1JqPNU7MDq2t3P22oKBhsUOYQmkMg799chy
MmdlhN3tReM0oIrnpUS6u+cqwA8wViyg6oqOLNNXh5OiJcdDeie6/BDEExakyp94Wcon6DxlohMT
nU3C/uXy8IoLtjxSUj/qM5xYqFlo20PY5N71xGB2Rk/OaoZcrQ5YcRmieqioT8y3l6mbRoLBKHe9
inEIecG7LOrnAhEuSKkrgzqFeFCCBv2/eICaLz1F3JnjVEidHgr6sbMN0adRO84C5Vp2y+SiXNHG
2794L4qAu8DeQZiV72FVFsOGcAiYG7QBMrztskw2M/zSeiFHfXc4V0n1LrlTKQxGXlpbNgzh9X4R
89cmcrYSleFhhVccMfLtMDDnzTGcLYTRLhpPN/1xwtyVwCnURZOGf09cxijmwTLn/50Oog7Ws9w4
AqAWikYl14yPbkB4+fqKFmN0T4h1fbwEExhR4yweYSdHkNhRashtnt+hXUA/C7fk8jYszodVGvCu
JmlqTOP3GBOpCgBtd7pNU9XKBb24ndDUbQYnH6wrvOVWr1YfpyiWTr2jV/Y3YLLSukbaJ7Tg1dJ2
lXOXj5uz7zJPGske4lka2xlxLxiJPWncPMUun/cjN6IWbr4Kowx8tl5O1keuXrcOMzzmBWx+FNUV
9DtAaf2RetduGBndhXV0vcLyfX2wMyUP6BDvhrdEx0jDrRe1YDNuL7VM9IzAN7NteQtBBYGMEwD3
b41anG7m8GvalY0PMNYFDbt1W9VoBIuMx+MNiQWKDfAgOzeTkpI3fPsJZqe4CGugx3WGd5YGo7I0
/j4lofYGYLynkU1wwHsgJSefkIf8o1hGjkFoprnN/syTGyCaRNrmsExOUL/4qj9ChP1IFLaajKe8
Zn6qk/mWbzgKnt6tVKBMQp6BVZnlc1VwoItJlI+SIAOOVdZUcClTulJBnp9/bkQZrY27h5mTPOue
QVBPmzZirEypipmPhxqxum3s01UzCafrQsWyqhqMVDJDK315WATKOhrwgB8KHrpbujWnXcaIIrg/
Ne2jtD8prf7y25vlL9Klz2Pyh1rNqziizM1vdm4Z8aX8Caio9Cgm5IhVLyxQCcxch0PtvaaPfUTO
cPTObqZ6nePPT4bE01nreGS365X/fXkiwau+XIZ6p/wTDK7pAT5lcQ0WTJ1oZJBlSKo70D8z/W9I
2it78wS9QO44ffRhMlzvGDlTGDtJl8eu5ns3TXuYv+IJG8GuY6vsSRGxQmywBsk2peRbROQRbRBv
Vxz8vIJCZf3ORtH8tEXaHbAzZ8qjpk2wG4CzYkbMqpvCUMtOsvNS5uLXoR58U/oVQxd9+qwAlOz1
NrASworVrKqHPYwsCgMyuTc3vuTLe3/byR1RPHX/+U0ZZ6byeUvp0VfzV9DF07B09L+RdxRELXAY
2u5FbdSstysBF0bj96gz0ys7m/CWkby5NRMCqDOH0WugsBoqquLAgzWkslh757bDe9AXR/fWn7A2
RisARlM0zh6zu9yiVrTc8crVp5nNql7udsm/ssc/M2PqAdnp5LW2STFh0taxlsVW0HUdjGCY7Mze
LAKB0jgj18HyzZBmKdRpRnHgveuIKINp8YczqTDLHp6VeQjHLUky2EkUjQOksGo7n98mBVa8YLVQ
AVHJLwxtBfxDIQSsUYxwsjEmfrxKbpJzERCFhBxUFQza8E5G0xGEcuXXKOQCqy9VoVa36U0yr28C
Qj3nRgzuDRNqmrUSAyHmPAi/agz/3nuTdcAKPY/Debcb0Bs0Xk1JyHpk0vKnVTXIG/mKtoAXwdRN
PY5m0SG3jio0ORFDMwxO62O8YEZYObaaiI13vxBg/+JLsPpAmiMHuukZBjjo/HyH77ioX9SVzJpx
1bgCFk3B8sycqEtAb0qo5MXPGESvO48bsM6vSbd7mvzpT9yOI1IorSv9cBDrJoyk5A0nkTIRyo91
BZyZVIb2IraL+l57DKlhxWxWgivA8LPCrXEKKqE3Vr4he/ve6Y6JfjvXkdhm1CIbzO/K470TYbwW
rgcHRUlRjppVXepoQQLZN/M4HYXDR5i9Z69nMueumblzk/GYJrhGonx6B9CMLQGdTtChaO9DC8Zr
uBM172v1f/gbfGvBFVOqDT/pH9SgkO00Hm6mGxSMTVZs3Ky7Y3kQa1BvG+ozd9SqedyXqAbZrFvh
AdD2ZWmpsrYPLdi4kaHhLkKg2d+D7q5Yy030AyTHNR79q45gjldGZHdLx9/3SX1pAaeGLEH/hM42
gtDRlEsAsu9N+a6poiT9OE/OXPlH7rUXmwR6dsvpSWAaCSIeRqRM0tl0a+ZLlI7jvhpFyxZi9Ghp
oiTNj+U5YQRxYGXxN6wBzIpIHjcx6SlzTORtlO+bfk0KivOQy4fWOE430EEbWk4rviUK2TsonETq
FkWivhdiDq1ZBleZfhDtK8vX5B7rUiEwpRq/f+Tsr5R4QKa+usCcUYRauAs/g2KsF37NdY2+Vf8E
L7lQw0hMwy6oZ2IPGn+PT8QPyuZzLmoKCxinF2mzSFLdZNdJVz2ZbRafLcTb2HFt3UHW3KJTYPmc
Rky7nSVOwELxHSQlUwnHZbENQ7zBFCMqJkXLfLWGn9VS+/4scX6koAN6iYWxilk4jAig8j7YlDGb
sskV2A8827EkFIcKJfs9KfeZgRz9B1Ryy1e60ul4XElBjUVoDHIP0czGhO3bVKICwjcRdiSMc744
Fg8s9yGa5kvBNErdfa9rtJ+E0bpSKPCeD7fVAa5HOh1SMWv2QtE4zN2wkAPKGzEQDIMW0Xuqq1qb
+wGKRdYHffjNdrqYBJ7BJL5CfKSbOG6UJtIfnPtHNNe7MdkQ0wBojc7RvPL0Y8tG9wEHINY1ZLxT
iAZcGUL4I8teDdI3jxVfyTPo3ZHDRe9hM/DZkMnzIr762sE4TbwcEFjTnrV0zowQ8BIDxW1dswj7
hmQXnncdNt9+r5wFeZsSTtwES2c7OhPgh2SXT6OqQ7sybpC0dvPuwF/v7Wtg4m9tK7CBdD+wJEQ+
NotPvTPL89Otrkr+zyb/d5FDKeARLxtpS2yipZquDGGut7H+BKfLqGNh1weL1B+d3SbmlngVYoWk
3zKh1exQ9LyjOT4yAKLyjm3FhnhAPZsOmrHj7GJc8w3xMgbyzbCNVgFwAKsgzuVRzRu8EDydCpZE
9FQN1pAuU3gP/j0s4+rNprCgsN7kpZh1yCp0vIQ1WSTqIqcS4LByeVNyYOc+Dr0NRstgG6QkwpOE
LdbQ+954fCfapocB64YJbQ/cNq6nor1MjnILtCW3cgqPVVvsO0xIE1iz8GKp2Fx//VBWrpb/fUPX
py98JSCbyAVATDSmNUb0iXZf0/DAF8y+YqcBb6OvXS42n9i20e8N9ZhyNRGUH9S58zyMOQR9ejYF
PoVpRZMbTm1S1Pea8g5zvAs97J7BOVmpcm5jYqBZFKKe7OSwTZj8UTmJM9+SzpM0h4x67xP6Clhn
rAfABRKzEQx5o49nnTtGMgyCKf4lVSzNgopJ/yf2pKaObNvp9nwcuA6uCrzy0dj1/BY2SBVUjem3
EdzR6ZPPiOKG0MKjxUwDVx5WzY6TlWMtvoC+uRw5HV0z0zMxqy4GxqYoQwy8iGvqblLEQhAmo6yr
gsD0gsBxC8JFdl4eTsVL9+yeZ7jzolN7CVSLlokoC6xE9j7jkpQ7lXfmf7OeWMY78e8vC44Y0clo
F+Z1/6lvpsfIg1LtGDiVScKU/xs37QMfEBYV2LEZNwMAjTVioRl5X61B03GR9gkrmi9mbiSvUJWp
qMVLlmee0O9EZXzRoDo1IYTMSEvdlqF6jxRnYlNmSa4gw8IyeUXcuKUxWOWidg0eaiPaeg9LZnt1
6RPtCGoTD9rXEPb+0yFNEvPWhi1caKlk6glKLW1dCzqOF6DRRt62OQLbmRrCQM+e/I1Eb6khN5+b
t5WV0SclErDH0DpF6z3NLOiVQCvB4WHfy4Se3Ntcd1+cAtFrKCodcEpQ7MlV6ljITFpmTmrjBFJl
bxMm8jgDq4WoFo0t4iNqfxK9wJEbnkeqXN1tQx/z1j4TV/jv7M7FnNA/xHyBjNWFqXZkPSVAUaV+
H+HeTptMFiuaL2ik05Q/iKNcJm5mQM32U3F2xYBG9YBd35zk850VbHmJ5EFJMp37AIhMxrBNn+2n
AiShLy1Ze0fHTLgB9cKcxM2Z5HXiZ+b306fsuypjmcAgrZy0ahcO9WxGt9423S7ggyAsJg7MXAFw
LGnV487aC2q/gjiSzQL3GPWXf61QDjzTVhR1iHO6Fyd9q6kvCj/zopb0Y5m552iizrK7Pmcpu15A
OSC+c3G0ncb/o/yeMsrteLUUBFvMXSLbW2DC6zaRhIrUrA4e3z4NNNNdCBZk2B4ozYKZBpj3g7p7
cYIFg9fsHloMQHMSuHicWmMyGBk37DjvpBZPiyEBKn5g1uq3MqWiTR9wOHJJZhnyO0VR4+wVZ7Qx
LjjyhbY3faaJxAOFhFhqVgNlZ6HQ9XCTsTGsQkn8Zre5E0bcYPsK2/XPhwRcxiXo2WCnvNPs94lF
Ftimsf4LQAUn56ipIJ6mfhEBEew5wflmrCYIMHsyL6S3J10mqWl1xzPONNLHe+/mGavu/0NExn99
C0b1UDg2Uoetlc5MGNqWPfVlbqgV6YPHvAtO1vrMs8z/jvfRTZDuM42+7FZwO5Ly6sz2kloWY3R2
hrrZLthMBEpNBo2XORuTm3lu20PVyFqHagH83Gy6g7LDVQXqLRABqQ1dc9q8voMiPIa6gkb3Qaw7
mmfrQpFbgwPdqApw8Hzb3S8kM+dRq2ewCXsM0NCFhbgoQKl/O5aKGdTxrk/O0K4RKfdDqQ+gbX0A
cFU5YmwWz73gjyWcUIOUQriFbuTZAyxITyomQ811BUos610ZIUNAq9tvCfsaaPU75eSu4ZwPwIgy
egpNy6SqRnWO9n1jhRrfa2eG2aqnW0zD51MElGQxI1AINYtuWv46YHGK5ji4kVNYox/SjWGptPWM
M5JhmhY2LmTJkOQ5DNSZlgTaYwiJ3DRIW9QSr/g07SpUvR9gIIBE1Zb2rTLkZQLVLbALtacMfhif
09GS7oKahmVtwWW9briFr6rgL6PGqDpQ2FH6PJilFgN3GH7E3LFwa36g4vCOnCPtXxMK3UsJyiwN
/P8b8ab2BFO8lScYWrgHn3o72mmC0mLwq8U9fvYS+P13LtHkO/syW+1JwDb4+JMDRcI4LdIq0xQg
lOcnntn1LKIgvJHX7v22zV3stnp583T5VqGYwEg8Kj2r6Sspx6M18LGunHkA92d+huGyEzb6m1vz
o0e+nGPfKS+nZ8g0gwACaWr4ZlJFpoes58BpMrKnrQabcA79ioY6fVD4rvq3EAizD5jrBzDR4N3u
7pQopoIqotE2tsLfYPu4HmJgkVRerqkH0ZiTws9RuryKMMNQzVXC7nh+r5toIfvddtD4T33xmffr
bBzCQZHDpFmVonE/AhkQuJzUlxRtgy3HZHWkuNnJuzHEsXdV7yeykV2aS4ljm2D+t70YbOYsbxW8
8OSmP4+6kObQzLUYnCcYnbxGs6WLGccQt69LhykEuY3lfgng6dP6epcloLW4qjKliohikA+eKIzq
UKwuxc4KysHT2iVZ/r+TE0yIV8rX2Y7vqQXbbsDsSeZzy/5wOya0fUhBttltaerC5dy6AyXLU7p+
YU1fUGxuMO5ckLuDUA0c9p3DHKHK9xxFD6burJlxKSpjM19iJaFNfaTx/WhO1mtVCWiJDA7No2Cm
4CUJ79JyGmjoPnqbipMv9UuvdUWHPr9yWFxpA4T37xozz3a6A4NCgq3X504yIbncM/0SMXf0Ljqv
ocpNjUiCrAL98kC/bcaMHnk3aD9RcOWCyrxXCuR6eJd6xsaYXISFX3w+B3ayvf05c6ZL4LY2n8pb
1IyFus2A6dOUwLbHmkcR1zVuRq8MBZhVaH4Df/LBHP4rTe28WVgyRqAJqbhWlIeOB32lkbPAlsMR
vFgFSgVukNtks+uVysFx0lvH1FNBW2dCmHIx7+VOdTjgSozJdVbSNtr4ldoBGAuL6RsO7qUzAFlz
mbtgolrVCoh8MKZKNllSojWMM9tlUlZlHyyQqhtkhwrYWwbIaKHSfj3Z+k9sp86VSf81yGNk6zW+
CJo1IDsmBnSe2ZWlQsjD5dQm3uhCe23lfTLRGXbztW71BoZKINpiUgYbgcMz8XISKyf+TjchaBn9
kEl9qn28DS2if/VCSwfo8uInbW1BDXIp/oSiq5mNyO9lC9yfTICf5fif39UX5MRZylOmWr8RgwVr
g7AEXYMdURCfGQ7Fi5IewRsN20ffhv75GV6mnsYjurVSZMH3LjRbmY5L6cvRk/B6KM9MWFQbqi6J
1UL5iddkggCYM13yIkIuxbGcVWfZz1kq8hYFsPXvp77wGENe4wr3hqXdYES4/lFzAhvDvRHDYHh4
s8kzQ29rTDRF1CFO7gZIFjTVMDcTQ2PWbyFeTkkG1QVoBzEFa4gNm9RrH+c2no/3vlXVJSxgbgbU
XlZifUK/jQUBmeMXrfQPPHAj2NFVJRmfnnK5vk54S1BiN1BnHhhDaSS0k9+2xrthwLUHfToDDFf9
TkrGD+guxIZGnee7FAfbOXSMZhDqKWni0AzLHlBlejfXZJWCK1826g0RiVILgcpVy80ZxHySrdsL
pWjWeU6Jycyv3qR7OxbhFydyOAa9iIQmzlbfBcudEdMlEC6TsZ/yqnGOee25hlJvyrIvC5clCLKu
X8Y3hIGT7TJfeuiMzfr6Asad5eKyvcgyrvU9mNMhJK5FiO3JgeNvLJIsxTCWWRjJ5FTzYyTkcifc
lYXMhqZpCmJLh51JuD9Z0Sj0DmdvLnJ2DZagl2hNJy/vK/MzNyyFdAQ8HhrLK7Un9MGzs4LwcTsn
55hrrZ0tkZAUHur1b45L/9RYueWPJaQodbmYqsSLbANfhHxgx5Fe6QXVZFPEN4WA946FH7j4wxWN
cdKDbr6wgCY/UB0TL6pQuv+L57igO7oPgywmJdUhelwoqtI+oRBMB8wrJImSduYG0A1dt0d3z++1
EJBVnSmTLlbjl/9itWd5ipuxhzwUFusQuZJDAnzFPenC6ncmKw01dFu3NUKYYQx3RreqcD9emitl
LC7LiiCni9yfRIbyKk0MQw5rmWGe+JKnXKiVXSVbAALhBlkxRcr1z1dTunz9hWVQeDhxDFuy66m3
9oUtR5RaVv0xfFDMtN4lNvCVZE3POMqfyVa+XSqw20s7OOT7sWJ3fR00ziC/Y1zWuW4/Dh3jmCXS
pUJvBH35KYgDHVuc7wIUDlrY+cN0keQFV/Ec6lrei2r7JYG6v5AGwBFTewdpYUNUvrDxnFoZRe5+
pnnZq0ArhHw2l8moCJdNDqRwg4nfoNs97t/lGFfSiqYsEIbwoJpft4fcHer7JooR2k7dFgC72+ls
Q1sfnOTuiadkwBc50RhSpXLqoC8IKvYycn3agBymw6i1KvdRyJPX2HaIgb/niuAhpr57X05quGDG
ozbLjzz5lor3nBu4AmUG3TLWdSrHhjjp5p6nvMLyMntKMsBFHq9lyla8eLL94oKJ/XslQrEYgark
HB7n+Ln97y17Aj0K2SQGsFbFlBt4dglgtHu18uuX9GwwS8eLro+RyFNmNViZf+gWee/MevNG7nYU
9Zt3rIqVBpjYW/e2z4sDsqzH6ua59YTC6ohHADIghuhutbQasA8aNB7jYk6m0gxA513m6Jn44zrs
dFFBAYuYZ+W+yoV4D4pnp4f7WBUV8yBt0fpzjhKhcGtAHD1wOO0Erc/UIMnzHfhQHY484/9HkjZ/
Kfa7OnWJcWfbaNAVTWiNm07IW3k/if4iPZcEZeKBJm7n6ZH2xqu907xsWRyGi1kYQSWiW0gGdxC1
TSz6pNpGWf3lfz4vTbgmd5dor6qbhyiLVgpCRj6GDCKFk9U9qr7xpt7IyGY1Pw9cwZ/APxrb73pJ
G0m8NOEKboU/EdboGUVebnws1sF5H7xuZ+rIJKugjewUz+4CLWcpbRIFTrk20952p8uvmujkJB1t
gKZylfETzBl382dClXwsqj46gXn0DgI9Y1hlu6k2mhbWZEEwpPdMejCEQ4nIm9OAv8hXMcHYBOv8
2krymmyFCdZxgaFrDC8MNdq/Z1ccgPHmvBcJHxiqB0OUMgCbEO6qQYN8kbzgACHRUGWtI15T0WQ2
KF2ji0ywolNUNz1gN8eq+HrhubPFZ01bKeJ3FKfHsSNe/sTww9nBWhJvh1+pUtPVSXZaKOGCEaf0
HwbOw6+FPmvoeJt/MunLJjq60n0F7LXBNHs1VlEJeFyH0Bgl4vzfpiJh/b0X0xcFoOFxjHwTCi4W
XT0+1pu1j/Fo6b2Fi6z9etHAiwfBv9ie9bhcBnBVpTwaIzfTWAksvB0u2NlitGPgdf0cNbUzzhEu
9ylQAzH/I+vgaI7AVq5g8OWCNona1C6rI+6ur/TM/607GWbJoVZmsvXHPazyR52a+Q6BuK93hR5E
c5SEsG+B2Sjif0awMrcwPl9O6kGJOg4upQA8Mhor2MIW+mEXZDjhJxNxLc94Eg1ZM1FzLYeCH6gR
EMAw51Ck5meheK30JFZXiC0s2UQ149F4rjWzZeTnML6e9JXXSm3K95qn3ufebqB6KFVYfeOaTnVY
vIfW4WO60mC8CTvTSf2IB8Bwkn3zbBQdTtPPjoWCo8zgCKhqCVwhhMInr0NBpr+DwOk1tiMOTFrL
1d+b2rbugrYP5K2HWYB6z+TxkXE7HHEHvUou6THOpbVkxeuSEqOFcY/ADBqJqrV1hBqgQrTYcTUk
9vEYoTCrKaB2gr88320blk0txmS5lw0os6gmLi/uQfadhBnTcMZ+6tR/yTLdC2hdO2+hHC+Thu5q
Jxv2NaUkoE+1DwMxI2OF70Htyf1VH9TWntVJGYHEyYI39RY0m9AcsuhTLTAKuJQvmplQb8KD5a3O
zYVoHkTur9j8f3GzqEDqZHPautNp+sUBxl/WtxL+Ko7MpZ8CXggsAM8kpm2nChGBAL4kg4DMkU5X
hIzeBeJ1IGn8lCnXs2cmSfLjVa+F4sHCn/0sHceD+3WElVXLUn6Dn/Y1dWG+2SWKYfaI0VyLNwLn
eek7996A+LNYZyF4v5cdxlBhp4lRLDQ7aHzQMVS1HYqtRcoOe2g9PHNbl3i792gN1/AElK4ZJ+SJ
/qSvbtgNhbkOXf1tAijpLHOHwAUTmzUZAAoPP5mXDskUyuRosiAcl8EODg0Qxrhxqm7yNELobfn8
GRvMgERpLNSzx1yH6U3ARGp2ASH9+llcdYpQbVlF1T4EnlsoPCGLVvjsZqjFEb7aaiy/Bf6OhXAY
aQL4flvFojjBCBISGNYQ/KaOHKOvxRqXvWIohCOkYqI0ua3U5CnbWtmNDVlOKXU/U3lqnGd7cS1d
bH0/k+4qII7nwWEerLUgdNFhI6IwSiUYvJNxAwasm7tlYLKiAkfk5yrBS0Tb/1KyAsGKp3aJn3p9
CmYfqs7EYUFUAUJfFwM2V1Fay8dA73lKigZUuLZ0CXppY2EUhw/tTdnt4M+SQ7oiwZ3f9wZqs99Q
eePb/ghPYTZ9HSTFf8b0Yq1SADc6wGfYsGL9b/3IBHlQnptJvSvWWXVDYtrrzhwoceESbPIIpjYz
gbAcmHHtod5pHLcXPI9MrfEuVubHF23/3KbbtsOqOUqM6rn9ewIvagPyw4M8WgmpAcwCGPi6QKIM
3N4W5ivnaIM6WJCZwTSrWpbv773sdh5s574cH6On03pwwoYtje/2iUZkozSRwMHqA7W9LOT3OJpU
0FDI+whYFVv10ZUpOoxsViMj5HWUCtpgJcdV5jNPTbVr5MzUP/yg/QqEoNq0t5BPe1usaQVfkGCB
iZc7zOWwrAW46aPQfIjCK4NNW6JWBO8QmWZwvzhtc+GJSVYMliSddO+WV4JbrLm4tuV/ZxD/X7lN
kjATPiBL4PzXa5tXAZGCHtJLMv/P6oD9DztYlWxthwsOc+/m7EIpqDoyX1wqobNJ9NS9ark/9Qp8
WQDKEPuMaAlCwWsVy/kNR6rwTC6g54JNi5MhEaxD4YglUcAPk0HAYsIugf1w8IohafyWcr2dfmD0
3GmQRz3sc5eQshceY6Uy1ivgeKnZHHKy0Fqu2OVKrc9Q6ysaaF9F8ugJccXrjUc02ofYAcV9GEhz
EWG6JrX5YskFttVbhx2G1d2seCbYR/6QKCvLr3+yWttRZTFHoXDgDYwy46MzDiytSxJ5lhJ8uG5w
eiUH1mVz9zFhEUUx0xIAMXY9trJCLAAoI26joRpCVZmXcOxzt9Q4qn1gsnKxOC67Xg+1XdOwYTYK
wGMWWdOMGR02Wqk5GR/x4hDk7nyY7ux2aQboEm8yyzSsEV70Z4aW8s1FmP+6qKvmAxdsm7S72JNR
Mkl/81DlmukRh23uiBIqbYD1uU3ZM0Z1SIcnBtLDVeepQfXUZIlRKQGGWoHXfjTBt5hX0qR+hm0Y
WaPpE0wqQGR2nxzn5eDJyf3BwqokTDnoPKfUOGQPYZ6aPlC8HsacGFDMaZbJjEXFrWEoM/fNFr42
jiMSfqz265LeOonUUK1oefEmPyjFBfjP4/UJWZPowZ6r4DMnDFcS2xEy0yLPUW/GkjS2Q31ZIKs3
CEPMsJ+XHF4yDf1UXe+Bu66QMhvgLb78D1oeIfARjcdZnZGJBMXvtOl6+e4lW8jJ9BR+oJR4I+1t
S7NERU0vZgipRIERL7/a19tIncw2BZo2M4ouyCXT9nwmKeWZC3BkLdnNm1XSQ9jCEqzFJwSeQImB
TbB6Rm+Rgmw9D6yIRdLEthaQifEJbwg0y6RO+NiRyTBPZsNItS2YM2TjT9rWoI97zGflPYzeVFDL
axK4PnYdS5VapQcmGB1xUoHcTBpzbEGpAx3OmygR3IqPqvsDUeh22UCJQStqCcIJvMKYzGWRAsAn
w/PU5rqZ0hZMXHyTSe2BU32MhmL7p4HgdcKSjRfNTPNGZ4nra3VoxgxFPkobmlaxTAvoe2zWKa37
dcO7HHKsZtsmarSXblOPbxeDCdAHykGinPTYvacezsI26OKlHvOzCt/JhyhmN9H8KZ4GSNvC+krd
pxeW6rt5sXak/ff8lBU9Tp81Ze28d7yzOdn/lGlVx4cANDLUX4GRCd3rpdW7BIY9dPjrgElI0c87
5+mBcnws3M/w0Nf5uKtmCBlRJ7OLI36nAEF1q3KSMkytI9vlWGmqipbWuBzI6tE/tUKQA1HcDZyd
/1VOtZoXL13Df9jqkOAsDO2/29K+fKkmp8MfDM7NoGHsTo1bKri5r8jXGs8dBEVCCmUdDy9YvVDy
PFZQntK7xspL8oRpEabrDDWRAtcmlXtl9R2lQ6GaMJITrnx/ob6ch1x89sNZS64pRJ5w5zqzEmlR
rh/E76FGneHdxsv1VkLfSLXsXvo4x+uQybG8y5BmWc+oWSdi54/EEK9c/70wevnBwh9gm7ClSFsx
m4FuyDcdwIV6WVZ2Va1HghlFDWz7pIgPfquT4etXKH5GUXoej89cSjWn05OkhBo3aL7pzmyMfXQo
9z6mgOmE5I1PiAYX+tS/huI7WzDjho4Pg/7Qd0AkbJfxQJoc6otKEBWb31WCSzDUr1AYS7asrCQZ
I0sUJv5DEyKQ87WO4MhKOo69YekSq7jkmyR3wCHdX5eOcKFlwri1sx9RE3WROKkPkVlczbWMgp05
rdtSGdc1xz8/ZhO9H95WqEqLfOQRCH3Q3PfZ9bo72UDpk6A0IXv2gGtT95+vsbtdSmozHzjDbZSe
F/oUsV6Cd9WsrsHuuTWxHIcl4LHrQ6Jyy8Oc0GH+GfjKBS55p8D3pG7G9BslNBBSbVqN6+qOJ8ix
VanCj57iFzN3q8kimuD+8WGlaLQn/++o6FU9hn2lUAoHcbuDHtv2SlWaJqOqYp3xJ6mP94/8nI8h
BMNlND8hMAYigJizGXnqytt20O27GXk6c4wDItYGuTpvyCMBKs99Oxl/fcE/iPa3TOyDv0zprf57
XTXacglVwtuBOwKA9U7y0fuPuWWRNS1NQ5wIOe+AQe2CmU63BfLNsJhfrPbC7xHKWWtoqllnxJmm
HRbkiGaP6Wpw6j5FLFiw/AMuG/DL9XFbg/rlul1EZcqN5uMNM3Q+o1AbIsjsMeA9r7aJgiW/DSG0
ib+vfF4AW3qOmh9VbKl8oe6pkWD3oIcsTJLzC+7MCDFC/ERJYMmvlJcsNcJoL+ZfXEzJvFN5AnlJ
1uyHRm1y206rgwAVOnOrHLsPJ3FW9JhrkefDNxhFYEb9U1BNyCpn589msWIF46KQvPQQ2Ngq6mMl
NXhrsknXyumbqOS2pAaNUNzqBUFdPZve6Uz+54SxjDLCftjC5ziR246MDX0LBYLsHo6yvXcly0Uq
rySjhS6ZYeE1XAbW1O3LrdT2McjzWoB900BmEeQlVxNrpD3WAVr3SBOkj0XBuQ8yGpIZHVv1u9KO
QGpFOb3Awf8E/ePKC9e1WZnCz2wrEaJ+TnOWKTzaHDmlrRkXSCcvPGwOYQxmyFdWl+NtfDL1NlkQ
P1xqeEUuY+CwXmPuSFl88p73H+i/gGwVuxHf7GYBbVFGr+gUiuGTvB1iL0cXpiCIqG35Dpld21ow
UC+ebOtcKhxzFTbj/9S2hRTqd0ZX+Yy0McJC1QbaH670EmGX7l6rsmsQQZw354et8OdnSVA44uEp
PfqfS95ClNLva/HoP6iokLHzc77EZToBgu1+xPa0h9DOaAxuew5toSuFWeLjynikAyVGpb2uofOc
uqHS35pf+AEg+9SQ1uhRm3lyGuw8DEQfyyf1s6s2iH8fdxVKJJfKQt/dO1s8JJnvyhfRwF8R8Dha
bOGm81V0AjfVyOwh9IK6jwsC6xsPZlcbQ1iuX0EhftUIYl7SmpLoMlP1QL6JFARfbznapPSxQO4h
aWPxIhcil6NBVTyq+9xh423zf5TvIZjNBUswrZBgSSq6+0iUb4D7txtASCzPE0J40fRuHOLSLEmo
ONpYc5iS+uIGLbEi7hddTV6xdhfpouDjssV0IULVXwE9LyzIDpPHPs5gjAhbebgLkzRvm7cDQ4Vt
oHSZsaU/GrNVxEu/b2kMzwZLJh3kynQdW7QWrsosbUbK3D2ziz/nKIVnex3KhBc4x83xwBeYNwcm
RvHegrZB1Ai/KngaCs6GHp7ZbkS4Mvp0QRgkW4RtdpiGxvjmIyEj7lk0AbZZC5VDFVMaVSqhZy8W
ZB5d+HGims08rcDcSlUN6s+n4uM0fgIsyBBsmqSJaa09S+3cLobNypwz+wMWhRny6Yj5U6/ilE2m
4DArSmu1G3jB5fg9UjmC/aAGJSGuxumuTMH2skPNjMKWlBokgW3SqlW0Zm3swQzRfPdwwtXWIvkj
/J59NzjVRggM1/bxr4Ulo6k4E3aLKn3USBbhScZs9io5IlNSFMN1N5cI0n4l49I3Jb8mJqUVY/j3
sxm7AZ8wkguS+ZsDprM/lwLe1+qiMeTOZ2GZyQAqOic6rXJp1iXMjtODslTtDogCXzr3SiWjQyrV
BNv1DtEwD1VvFa5S6xxqzQzcHRDW2NraQdBha1Z3gknqH4VEM7qrth5vstIh8h77qBpVicRIyM9o
MchKaRVBhUZsGE9Migx89iZSgplrM8kNAQg4HS5YM94mYqFeVJMwo/pNN0xQLGKBNsCFY3JVeYMV
MOv6RuQgkI0uDrCAtvq4KI+MPqOtuxtg3vcSBrGQVSZJhbtgX64x2sTiiJaeOq8htx2qYA5msMvy
kDtrhqqxjPAiQWd5KX3cSuQ1N1r7W2HAzW1b3oa5xPyZG8wMrw5JwKAtufpsW2O7MCv2nrtgx4pa
xxizVWUR3QaIHOLaS1HZvL2n/YRnY3+crDqIyThjB0F5ZquTJWaMZChy4ecD3Y62181m/cDJ51Eq
sk8mbhLUsScGoFUWh75VbMXqsRr5Y5qTf1GHCiYWgD+1CLq8fLYxaDgOyPaNzqijw1HEKlDI8yoC
8RrXp0HxynjHNWdTrMraH0HTBbQc8Ibe5GVMIXNrBeCnvb9ncsqvvGW2Q2o7Z2+LfVQK3FJmFIjk
sFHNOlV0WM1feYhrp/1KZi7VwNdKMrIgwioKOzFiAnsjWefrY011zn+M+nwqorryAh71iNaH/Tpg
XNdQNgZ+UWidI2V3celWMhHztBa5PY5Z0PPQQhBHDTPDMBv2XJKnmJGbPSpkWV6JXYVbPw1EIDkJ
O7OJbc7IhgCHvKzwEBsDPTOx+HFoHTSRFUfiSvj8D0rxSUl9h5Qjn94tluOE02jF4NBo+3hXhcis
Aat9m2KFtbJ3xjaWAehcoJ6V8nhyH1RdGkRXBc894p0pi2UnTHOz4NKj1WCjqQ8ZtM2fGFiFqD6Q
8tBGjEt6Nc/LVAMYW2aTCvOutWIGHhvnRgsGCScAJTlWePPi1s5yAMJFfbHIzQK3e0WsFsNgaV+t
qBS+SQ3DHom6hEDwTl1eKQz0FZHX3AA0+m16Hr7flxh+hKfIbc7JFkcxQjFyl1eiRFTAf4A3K53m
cMwNo1IYQKt0IuvQyRyV8dJhM1EdABaWYhLpU4OY1p4+xHikHmjJriIBaj8tZ/OX728tbdyWztw1
Kx/Pe9VSM5z5Sa2G8S6q2Ongcw+1Po37Jty39FOzaDuiNcwSaJUXn9zHCWQ/VtsL9AOS7m/FnICh
wt4y2OGwq4Wu85yMflt2F1bSWFzZ6YDEdxHVifjb/TE7/Ns4ZLln0mf1J8ubROdiW68STCBsUSSS
C3b9avpJ0rj1ReJe0ZUUBlbWrCY3HqfwAbGLvssZC+AyOW7TdeX3mXeLcQopPo4qEYqqz1iAc4cG
jquwKdh/7LanXQ54PvLro5OukcOHt+1LjS7UT5HEqHtJVHxO145v+ditSfw6MM8waWO++aNxyWlC
uOz3NZM2/sBNLZuTkfm4+t+fuSPJXlaqRamnKVpQMycOELne3IuL9heJpENMyiTPP11aSW27+Ph0
sxUlhvAPQPjH78x+xrFmWr5J7sYf0CzKEnZ+qiNtS8sRi4yXVTCgcvF4Lt3RV9WkCFZmkfzTaACe
0HjjxMObJ4sUt99KD0d01hy4pCYC5My/dCyYjGLYKZ2vXS2gM2AYmizcvmodIJ6JTiaDHnSXkSV9
5ceHrfBtJDyQmMVy+k1pNuJMxbH5IgUw3CBpvpM8lYYJ3AadCX0OctkFdZQ4l8CVMjL+hfsswnSf
BZGqzCynHoFAvSNZbmZhaTgjkm1RC2kAiX7YCbK+R0ZFDYNxGM47qT6ag9jUHDYjS8gCxBZEMlH7
UC1xIzygbCAMPLr3GG/R7WnJwS/FqBXZriT+butGQ3zuqF3JruYSZfrgPwetENDzwvLTvcQ+l3sa
Y0tn0nsI0UpZNfjYAklahiJI6xGX37pSozCctxCQVPapZdHnRW5YGTgpAjwkgYvcElXKKrRje/uJ
Wj5Q9ogbB7dL2w3v+3R2Mm/FL0NUDCUeIshngukXX/iLT3CNGxp2QXBPbsCpiivOtKyQRQubKl+8
9UUpTxT1fOlyXTWfgaZJyKung9wfX7tmtt4B75zTB02C4sTx9EpQivMKlpXpLyf6kzO8H3tSks7a
mLKG+RtQrems6+vliA5c0OvW1q+6MQt7IXctO7M8f5Q58FV63UH1dwxSOCpfvN8At4QXFjSh6vFc
dfbymQr1CCO0OvwHBQtIYvBCsbXiKM5+BCDHu0Wx/WCKo/LFPI4j1UJET7eVpeA9JhSeTSCN1Fgb
mkbiufdY9Cr67S2TF2a/KHuht7tOblkrdd40aNWPo2TgRweCYSsU1x8RV21N4sI5sVZsVCsEWqwQ
5VQ+YYUjhxtVPbIYC9W9BRZZOEyuyXKPbsDMPFkuOgFM4VZ6ag9xETreMHUEtg8Kd6OrXMvvfU0S
sVVJSvnnrnXjvzSvYUBgQGHpKzepDO+4ECraPk/fyWk9HSeWE+75MTBstBjAhsaZkiM42N4NH0q1
cWUFPNli816rKBrBYzDOAOJ5AJa9avW4wfSK449utUFwDzJ2TNFbXSSFhFUqDVFkVrCPEpTiQtbN
Lopm3CCtZE/7LbHpUlyZwTfcUMltYjdnNormghak94liAeAS68qKLV9EnW1nJEAixSbPvUsWkoNm
wPPRnCKc4vXvjfZkKvuSwqet+RpJkRyQ5x7CDwmdprw4GolSBwNnbVJtNrNQfXfoVApuwxF8rxTH
vW4W3ghFbmYbJ7Kkr9AS65u9QFLKu5L8KLXQFujbQOCwCJ6fdiz63s0432VGXyNeq86mdJrPpXXi
rU1VfIB/kUQUsph+l/VG05jLr0n6oWhPBOIWLyaEPSyU3x/Z3zSkvIaNdzNAZHvgqmgLx/jo7xyh
meI+bpcvhglfsrjOeVpJ5r1vuaZj/E9DA4qhE+Zk2DjUSArz/kfsse2lWo0hB8A+ZSfQd7Wp39KC
9BOq9GeAuHg6m6ZQMil+hdriwUCcAhDOtr6gFfnFX2IIK19M7VJKP5WiRROYcpJwpehs10SiEzjw
GAQafqUBGkPSKQi+d5cGHvRBh/GZsPJ9O+uIvxY8GQWJa+4dVCVfmFnrsoKF17ELLtU5b45fgrbk
aD1WJRPkFR6TwlzbIPDansMn2AIAVhGWUiwFGjPu9BzBrdyjp0vVi9oFa8u1hsy+WlKLLxF2xJFk
jo8PyBn9I6GHczKM7BVV9A/z6MwYP8o1orxtpMDv/TbPyCs/pQcJZc+brCaMxQt2gFM6w/SyRx3j
18zMfuvDIuwR8b1+hMVXRgxSre1zG8dGapj/R5kkd5ihjqaYisA6YNl6qqgJd7Nkg8MTGdv35J4r
cGV4NvCtYzCc2+7qyci+M9nxiPAFWBNiT0SztkXLvfjr0L1nPji0bjbkTAHRbbt285c07E0NtZwG
YGSJElw65zJ/ZdjiqjJrn0aP6SgDaNlzPlgsmfe4mlxcLyDVtQs7cpYxWU1c17JJrN3Kbi746/8F
zinTjATgz1ZuE6CgobbcTkHJDTo1LV3+5TIwCkIFmJ1Jf40gcPsbUhYcVN0o5HPC7ipqXhYfQcqd
Lr83U/0SGqHVA6VXJdnIqTu+3EssH8/KL1jCYiWwsCeZYC1C8uen1znBC5/ZpvVuRy9I4xDeDg43
IVk9CRZuk2l+aPu8PHOTvOF5qmwOV3BSf555nvBk0YREGTxru5vTorzG64BAbKdvf1lTJMzf8I3Z
Ejwnuz0vWsZSabAr/AZ4W5oQm/vCocDpaE6cRSscdnI75Z51Wlze8UQYXJlouGku/KQ2R7Gavude
An4Nf2OHhXgAxCC5AdO4xwsHwc0Xotvz2pE6V9D5iD0Wt3lYV6Sgqhj42mSgThkwZ5hMqCqUCMTa
G+Po/sTuC0D45br+88cFn+NJ4Oj6LZH+9ndydNvaaBz4RkFpOaRrg0K+q2C07Yo/ycajrhvf6Hmw
D3bk3FxnNm4buCjxN4A21zzWC9DDQ5/IAGOBQBEtlHQayl5hQlcDh5x9HLQwjxcFFS9xMv87H6IA
e+uNHb+rMbrxO3UhTjqBgZelG6VwzEiOV1H11Lx9iP6ITXhDxNt5gQE8r/++DM9VPDl233eCAeHx
AYXhVHr31DM/oAp9/tte63Xbs8SrdST+DkkxvqbuUkGeHgzzF24borlCdXh2O28LfiaGVd6MZjEQ
BZci1BysbXR8WrgCdjhM5WrKn/Ft2a4nivQfP4/RG3MP5EQnaqbsuP1klx0eC4wzrbOtBT8dnu7F
HibB/1gCiKAhdwKN+iP0zGA6gtCLL4DFjq3R6iR1/w5p0Nh2IkEFsRVcEKN1dUUKl03qt+W/9vK+
Fpy/iP3r+4M/WcVY3mBago2rRKGgQkLgACn+JRaXD6IBLgErKskph4WNZahVDEaQEbqvkUO288ld
ZiCjwD6810eAxzG4ZeIL3DVrC6qt7yoLq9kKqCHgIZqOcVxb64N7ZGR8C6QgOGyqsKmW+E9zQt5V
9/ORF01uBKjLD/JcF7hR51nhQpE/57BeoDJS3UJxV00zlRz8LJpGAXIVxk0GU/qxgRoxE5duCKAf
iCuyzo34xGleJp0sMx2me0Iabe4FGYppYbX3GM2gZvF0DRT+APYKp3zCo7PjPU3+fe1+3mJTAGtN
49Wjds8fwD0d3GNNJRdVLMIE7xelxICX/OwtFMMp95kvrqR6olQNnAxZhrrkySZWXFxtIn0k/TaV
R+MdhKjpm6ADVUb+MWc7Z1+NPW/zJO3NA1eg26iAGWiwHdzUOKfnEI9RjcVv4PZQ27be3Xdz+r5i
WUHNvD2z0sRxZw5EQyPMK1dQbo5MzcNEd+5r0Tv70Ga5hEQsqNTsIbV8QVusVpVKmUoRNUEVF/4L
KRRUYh3NxnSb9xyoYBb8yUPTcaRObgNhzD0zsOC6Vwr9zT45AzTfHkeIAnqL+ee2pg8pbOWtcb9J
8kVd8Oj/Fzvwzx1DTFewdSg+l6MnibavBgi7K/RkE4L+VEnTou23YoPS+QmnyHe/6Wzzv8idiL83
eVoTMZl0EHzWsmaSevoTqHLAHrq9kkVqqYuRZY20rih7Vya0A55wqL8a6NR2HEYMToumbK4OO2xS
t9nZR/8ae6ULOXEpE6Y6gFKcGjKCMVrlRwkOyayBNc2rBdz3eiIZiFbsyECigTFY9roPeUJOoUZ3
goo3O0gqdBZiHbYXUm7aPfCGFmeAhwPmlWB0YZ8zLb8RfWprumf9J6b+nE4jGq7QJDuBjMTGlo7J
pLzPK+AIaeWi1QDbvSFJTjTeXkjSF25vZKeIJdaBHavSaD2GpIYFcS3qfiRwzpUdSUZvWEvoH8Y8
cDEyYSpDn+bq2Y9QU+BPVu2KwURgwnW/EtHA+pzakyFWe//ns4xNqD9QQZPI1Drc2EnluXT3JIPF
kILUZhYnb+0FwWnSPniPjd9dNHo9Sf20BXFuuWvwiOXcQu7uwBJuxvoTsmQMKgm4r/E+czuTR+M1
rsaHaPBpkKX9ENpT4cpIjsbP1ZWItaCWXl9KsYDlzBlSc1sFA26FhPFDAqKvaVFlyOa51nSYLK6l
z00cBvrtgO29RCShwSkTKgc/hPwAWnZPWShzhwx6nAtNpy/a3tTUmJAHUUTFTA9lj/FiSg4FPMgC
8l3kk6j/n7CRTIimTrNC8ou4lVnEF4FR71pjCTtpuGcLBDKyss09+DZ2E01PtlFgB6r9q/P+xry0
OaFqbhJLExBCby9mzndTsrZm/jeRlfryAXGg5KoSnEEEJfint6Swr0xw/ioKRjb8AvOgMn4XSO09
q4FK3HywDl83vG423i+IrHT2fboqrt1BiAR4DAVQ2hwr3vBlEIMLPs2wlq9Ea38IfFxBbmvbG7G2
i5Ht3qZEk/6QGVn3zvZZwL0Aqt9UVP1D9y1NCCaOcbLtc5PEBXyFDcHR8ExrEyifSoSN+VXNdfGC
0ksHv2viZ/x6ofHi/inJmBJDHUdvkXhudhXaz273W6cCwvg1d4r2hYZDpYvDEOvA5OP9dwEuC6ny
ARQSro5iQZyds+b34FIctaeskAbvkpSVlLNQ3DYk2knjEEjfOuSvBUMDebU3ZWwRr4e/Ocq1uF/u
IFxqrMAjkMtSRCVV9vxthOH+Od0HimeUPsax5LD7nvDAak7qNBs/k5xY5PQnYpjWKc3g/utgxOqI
Ah+qhboxYT2eTNFhk2dErKnInUZo+4DNblzzj9VN67tl2Ikcm4rPlOpZSxzoHVSO5QbxhLp23kTp
m88N1w/Dxu0e/E+7g3Vqw5vi4AGxms8i9109I4CSI/7rI729OjkK7ITsiknb6bFWcWwEfARQVdoH
ImY3I66T3QX+7TcuAD0dLiVByfgiVUlmPZDkE06dJXzvoQDiz3umAqnzjGlHkXYCmQh+a7mL3MeY
MIHPmoJVAUFmAdVWr7d2Ren7tXtdEvZWOJF6TdjX5QAcEzWx3Neabzet3Gp8LSSzyLIHS+y+bLda
Gy1bKer60W4CxPwT3lEnYFf7GjkudfCFzqMr1d/1JobJVvMLVxN91YGD3qkZvJuV/NIdgQDL8wGn
NqtlLsSKFFnZ50SU+v304WrE2jbmQj1KNAFNmyJFO/zw2DqHoofn+HNehJhM1wHBBeS9QiZL+Zg0
BO1CdJDGfAFJpewkGgQeMeFM1iRXmyrBoX/jmeznjkvA2ULp4aBVE0MBTzq7HquBj9Y1CewHL+qb
4Uaw1uUWiyGboCsHMq8lz9tw6EYFru0oOqHiybOwYwaMrCrAfRyHjCzUAMt5tx7KKTEEE9y1YTZn
7QmVeXWOtry26mw92yFbA1l8uDC3t+MvxrQoBaHrgLWH4Rl1ziNr9XbI1qjWajGKrFJ7hPsY5om4
R2Gu21cRG2XjYUXPb3JYvlbZMsx8nDVpErpHa8qt0LvRHCxhVnrEEOnLv8wMPXrg0avOGgw6xSUB
cOasgAJdNbtgRSdfycWHJmxMZ/QlmDVpemJb/rBfFRVt/VCLDtf5BK/dV7/0Sy/vBZ6zTZXebRWW
QjXKURJxcLlwdD2BgdmZQjZAFnbyxkZvW9/mClyD5WPvNel+MZ4B9rGbgvyPxj5C2ffsXLepL3HI
yXrATEQd6DZNBgZo+PhmH4/J3qZIuq2kEpBXNpC3Y5EeaA6FZdXD0oCmPpUU9jhcNKjpzjlZmOgP
ZxE5n5HkKa799fjFq4+49dwQYVJYLGH029orSa7XxzFh3EDYWYEvm+HwLKTmmaVEQgZURWRKYIn+
/NGm+5pw+elzkNXgAgZvlBjayWDNBn75jJuQP+iEWaK2uF83+dkMOKDznvUs4rx63jg2qDObeGGU
Sc+XNC2t4MkUAejsMWsIM+rMWHxaBSadDMPN9cHn6DoSP4AatMmg/wOEo5J99eMszEWEg8us2ohc
Jccsf/6qvM9pIdIQc02nj5LTN0SPSy9llmOhQ6HkVZ1iseJIApQQsvf+hBwS2MHriUv4dLlpBe0q
Fu6ssCxlclohKDDfm83lGeEPzRBWwP/kvije7DipGgdup75jLOMJ2EtlgAEFfoRDfLN5+AWk4LrO
w2OAA78rYRVN65kleq4zIpRhl8ICt0auVwGQepjbQaT4Ip9daxauJWVbW5IVzUxTvlkSaLyOtXtw
xr0Y7l5OR/+KXvdVvebyBFBcIVBtiRhgpwtlpHZj9ysMsnYEVf5vv/E63XO1Mbc39Afp6DfnMU9b
F3LXjx/MSQ19OSB4Ei5x0RhEJXdijqYsWsT7MCOnJ0zJ6705H2HhxFULKpS6IUqu80VNa/DqFfQn
vKiHVCkVkTQX8bynRgaXm4eIWQsLwXhMNIdhjEEPJanuf/slnSQuf/E581BMqW4CPSiKzdkuEBD4
a7z5v/tboAY/Ufq55fhGjRZVY4lSOKmi/51UN3Z0D6Cu01fHhYpTTsp0S7UwwK/RLfYUWKxlAcj/
5+GhEmK/hWTfmPE5YhfjSYejT6w/fgCZLmi9Mxqb2XX0U3C4XuZSQLCZGpdoKMNOMcNVL6rDUxg1
8wa3itZQY4ymx3dGO98Mg8R/u9hYJNE+ADJlyDaXsckenbsP77alQWdBaaYVFSH+J70RzEu3+J4y
cTdG9u2A52pJhk993ji2mUhDjrNNp4Eolu1xVKAPYyoD6XDq2L2iGmzl5ldk5TGQA52kxmUle9SW
8D+k7l9N9oKfiv1oyYNxgdTkRdCdm5aZJMmT2SsJPQ43Tdt6GwlPFasiDPEHSxw+ZuuHMCZm+iRe
IIEkeQE0iBWtOPAzQN9qqe1fsP+3FdZOT3/YjnLb37ZJLJspMunW4uvBmXDn/Dcf04wXWhjJ23uL
+sc8NSPp8iCr9mp1/gWAf+tj2QSf2h6wCXleoXB4uk6JAyH3dP6dZc2y/SsWx5RmQR9rmoef1/Uu
BxRnp3etrVtqg0e0dgCTUrvjW1DWNkZJBVD1Yue68UQX/GtSmcetkVoy4PGBuNwQvpu0IWVUA/r6
smX9OdjJmRty9XELJk6140gZwcABWeuYGaxySzHZPB7pkqhWUTsBoL97Fq53mzAtBBIWaq/tgr+g
JxYqC7uX1OOQg9DNla3FoAdfog8CUCQLr24dWJscuDo3yKyuVoPJkLdyjvO14naJMFau5OXwfdD+
q3E8Ib9iRakJar+c3OR0CKAL7tTaW+prU8AZWJVUFZw6W880QQ/aS4bMx9BjQ0Wpv694vS0xS1hU
QJOALB4DiCQRI8unj/ItdCan9daKPmeDYppDt1jDzV/2c7bAgoayoN8K2YDFtnFz+8r+N26KSM97
NexfRBzze58fMTNDBz3RTMLFHY+1LkOfZtRbjtUChUqiOkMwG7S0IT+e4XuUAc4xOV2Cyz8fzQP6
zhafVUSuKSPYRgaCnklrV19m+Zf/dhWUvMK3Sce702cTL404Vk3YDpy/Cg0CebyrPZrJubptsg7I
R8lrqylvz3rw5JUG5VCCkV91r09fhjFSczBt0ud6ZZ77EvrEMH6tu4PBqQEC+slM/dzvGusiMg+E
TWoeW51XUujXI1Yp++1gGaJSDz7/tvC8d//d6S3f1HxhJTbA8a2c4CXqc642qfX4bgBLg+qSWWSd
GNjbYKnB1hBiny6PPW3H8lTfhQqBOB7u22leZX4uwRqxtxyPLWj6V5wUbSv40urn6MTLdo+6YR5J
68DT+q57S3ErE+H7FwaD4xnFwkqxOP6Vuoaq57hc1S96yLFEe125g/q4OKOt89vT8Lzbzv3AJten
vO7Ci32SkwsnS5P70avfJ+Uo/RquoOH2xo30R1FpevvxXg9ApXCaI0UevpRGLnLBkIv9cVwU3c+s
EEoRYBNa/rSd66dK6Y9/ISML/7bMyleoZLQETrO7DFCfc8fvip7XkBc0es5duP1PL/qgSLuKKXZ1
Mxx8X+ldC+CJ0CoarIwme6MQtyOUUyW6SJj2vyOYYghNdtEZMbDod30mQA/eVGmd8q0S8ugCEhBa
OGSU3pfWTwbENuycBsk2xzQE2GPsrV88K2kvmc8XPNCfF6XCeDYQ6fb0Z+oX4Sz6zOoZfms6IGqR
FxSognc/ugWJkIWYh0vbJaS9p50O2/yhqQAqCDKlA7VkBHNoMfqouBPbIE1J79ZE1O54+wZJbafR
nd/adbHNNXrmUKAcS66VGpl9+Dc0cuAeaYn14t+xVY1GAH1CPy7pKOL5vcIpiEqqCd5s2IPTLKJ3
tXc+mOeZZ7Dosvsj7+oyV8XDrurjBYYsb6DCFdZb+JPuptriKNKr71SNPpLUYvWdjgIduGvWwVDF
a59HiRvkb7umTjW3DjfR2PwiuJYIhxdqoPyeXu0R2wV8v9B5ZwQQZ0axIGQFDxaGQZgfuy0/Bg0O
T3r+hg1yk+1REeLSth/Jx8YjWyGva+9DA8ph2/w9c3px+AZoSCVJLsr4Y9nEI/eJg4RgxyABx6mG
P4lep7hEIdHfIUpFZfLsZ22eCyYpIXkX6DXOW7UTr8c7tL5+rXUizbmP0EwJ/ibAM4zkiVE8jMTu
oa2FBg+QBZr1i8nwEg1vHxcnermNPsM3NEmO1CRbjKbYVEcZSr/Ja7tcb/ej/LJrMzKZtZEytdqS
0F29Az3zy3jVfLrc3pApfajGSZHe+g/XQYHYkmDnRi8wrN1oA8ug7iNUSaDV4uEkRRYmZ44mIG6q
hUam967t5dGC55lCDoQFevBufXcV0knb3uIymfK9vQ/hHDMkJLsMMkV6SlYI1i3PUsJoBtdLJ05i
1zO6pY6tqr3EeOSicze0Eq6kqGFsukaWjgkhuJfsvYfEtJxVq8MhxhFeGcVrGbFSBmMGq913KqFP
cLAFXrPfuwtC/KElY350IqqG0dgBXt8nkfsc/y5fzRhLKP7gcKnNgE6pr7hGBcJCCMVhZDbJof94
ZZLY6j7/PEMYj9f51EkRSmGCMCC/RtZNjLqHzkqnkmiozhphH9wilvGGmm4GEVl1XR/D3umgkZWp
mXrs0iH1UiGdtk2WaBvJZftCv6TuLb+ViiqoNAaXCeWSQ+hXfBvQ3C5vpP8pln2xmTeXoUEeiIZW
nuBVqSCQ6ADgI2dvGUtItqp17m//7Xx3FYjKK5I2K053kY/7rjJmj3A7jv/xctZ6MWfZziDw/i3E
SmcIGsOVc3vUSaNlx7puA+nljdN6LK5MVqhhT9mSQe6qZNyXQYlluIe6FGxqizVqBQSENPceGjRi
AmNhAU35Cir5+WcSJ627QrI5ocBNh/FhpntaRK/AytKpwhOgv0723PplLpX3K8C/KS8G4EMDxBcX
IAuLclh2MFV/2eR2NzK15/7YOmCTf9GJzHvvc6lLB1ge7xLqcTAemXOWWTBxD9JICjIDcgOTU6Re
qGsf03UIoK1wSKoiYLEqfVC5yT4hQQEx8hhLFytWpGb8TGLIaZJxY9g6sHttBZCG3I02jsZvxANt
yRg3ILScqXlzvngZ7NRjurx82pZtAZhpMTE9M46+Yl5whMS5sxx03hJsnRavckNLHCPxe02JvRj0
yGNpO5mprhn63hbc3ZyApL2bKRZLkfXBwRhTWv1/if5FPAKCBjif36CeNGgtcfegIEUu1FfPrwh+
VLh8hfa1eddAQB76KJpB54EiFRhNKmkgkcRv5Oua2tGd0eTKnwojwK7BIHuL4WtDQvmHrXVA3NrO
44SBsb5lMahNSjEbRQJ+NM3SLVqgaLDOeI5rrI0k1pbZdNZmasj2p/9yjPDbhBsYUDo6sNfrnwNa
trXe/CY8WGNxh/ydw7UOdR8nFomwVzOTX2Mjh55dvZRZFYqobRn/TkB4F/IOs86q96pqsjsBGU0I
680DCe/OOD7W7r3Bd8VHkpJ2KzhjTq1OLAtmsZk4WFSShiYTSjBD0yKq0wMg9BhoR7T8UJBKL4st
ZmzCrjUPGYG2nfTxTk5S/z8KXEuBLr6xeZdpTfd7lrTEKGabkMu38pVrwBoE4oghRyFguNXKIwz8
UlZmbf4zYbF71K2Bux1KAORgB2erCrRsBZavN0ITgoQhy6YCRLx998X3B+xRQS9prXP3KwDpB4YC
817DJZEKIQwDsATrG3Bm0aRbaSCYoDN8pOH+KYtbWxrZI+uQg4zDFJlmsY/+Un6uaSqqS74bxxFU
54UyCWsygSjaWxO51OAmj11dJGPBapbplHTqBHKMlALAHl52X16FglmPaItwf/VrcwlEiGQdFsYG
XV9DN9mEzw4RfCpv3Y+Eb34ivOz8DzyD8uApQV6pPWNiBMkeRY69/sCd6AyoI2F3M7CGsGtKhf3S
W2HGEkgawYAFf+u6rxvDolSUgX8fVDXcuBjR3Xs3/Wd2BclhOagDxoM7KqqJJlUDjohvIrUrn5V6
aZ7tcrLH7somQFL/k8R9ZbCLWZs6LaoGY/CUypPmYv/ReWwjp+Dque9i2j3FWfy1jJ4y6XNQW3oG
moENpBH4YPqx2S0IISO+5yZ+TacpWbZtQeD2bm7yJRfFyY/6Kfm15oZWWnERzOoE+95i7trIws03
1Wbp4EOibfi2sDwMW2l5xoG6sbe4bFeVHG9DscVqhpLDiLbvlAF5tR4tSJjoD2v5wz/zSs+aAZ6k
r/gzc6JH4TuYGZ398OQ21qgsqNEiJ0kccQMjoHsgVgQv4xopynfQitzlENhcAT5R6iKlec8gZmoC
DtBKX5tHSWxJvuKIHWtjI4vHrnsFBr7sSER1np/zS44G1bicsF5sRuunhHZCbvCszmap3KF/Qq8d
GCicwnd6otrRwqTA7Jao8s8inBDAGw3jkCa9JhHTPuRoW50JLlDTZVHshcyIOLrlIKFotmUkvTU+
Ou+4fhpen9ORZwaFEXqOwwuE17vzR7MQSsaLyWmMQ/pN4kQODCqVg96HpZU9KWRDdAu2nTdqrxsI
2HZ4pDE6Uz0ibeYRiFh5Lg1WUboksEPWPq2nNwTifgALpKt+XUCl7gIiTzn8QrHF3ecE5u14EHz+
ejJXU0cR8xZkfeOVLPVtcPkPZr0Z+RVBQX4xgQW1jYrPXo+Hjv4Uwb2fFI1tkRPdKKcBnd+A95ZN
vrC8NrgrGN9AYMQ1iaOXitYYYMt/3iKNWFYIr2UxPC44ZYr9RDEeLDNqs/vpHKAJD/Rb4mSPiwx/
qo0ALsgy1aOJhQ6KkJDSc3XXyF+7+VSeq4TfKPjJf7qx5UYUfYvEZ/BMwhbH5hrBUHEjDVcD3GFt
HqM/BqY/PiJyDULB0I+/ZedLdj5V+o2gVYJ9ir5liuNOIUofezWCJ2hAkiM82fFaaUFOHO1T2W+x
e/5ui8tv/CVZxVpSIfle5+gRifG4CqVqWa6JrDvPu4wQnZd18A8GrJcc3ZdEbTUuixZRJSNOs6c8
x6iIIKDpwZkis5zVAjobA/GfsSdZjHVECug692tLQrXumiAJBcsfpaCYCtL14kSrKMiFYRu161e9
Nutmp7Lmxie0/B7rvPSUnE1nFCAOKyclVIBvW4s+DanCxNf0dNoJQhq6Rfi+nZ0ICl+s8Uwe7rYW
MAk84J6YsCnaSzWd8zVw4KHJqE5JNkULx1LewgexrABfWXVpliCIJx/ni6NjINUgqu6Ql17QHTak
2OCjV9QoyLYj2b50iaSWv0X7xQmbJ7gMVjS1Q9Ks6IHDA9Rb1FWfEIP8vr5shy7P81fwMD20lmUk
4hw07D2W0NIeg/WY6QMYneSWg0RaursWy5gkQPAHFdzNv4m+1179n8efRRrpWkcM37fEWz9B5FMQ
hgbHl5B1deyvkn1gxq5jBSMR0lQSS5jUXhQPXVgzGpBl2IhDduSh0kK/mROhnK1Ds8a1TXjlFzfs
JKQtYFCXxd8tNqCONuNBGRVNQXEZMX+PP8+BkIZfha3Ne0IyafQMLSAZxVmDOIFKd3h0t42QdSJJ
qVA3whEpdsTHmAt8QU/KW6cb1ytB3xKBZt6eBPm2ALL5vdSDXp0sbtFm4D4LaE+EX5Q5Xok7/ahZ
iFUkB+UAXwf4KLMApKuDF/K5PsXHhz2OXf/dLzPwp2bmGKqYsqKBCo5fwBhUgXgK0hRwlp5y7K05
faFF5d4cboOjF41GY3EmaJjy0mtR+Wq4pNUWnoKcgleTZkIFbD8EtsiR+rRD+NN7tI/WpfWGfBsg
xl32/BIKfgh5ceZgMVdq4liM/SYJGbRo2yqWokY3ek78hXzYmKa0IoM05OO151N4i6KGfXs+GnNZ
N05mUaJSgOOICJ4BMwTbvDJ+K4JDvZTT7vviVjiqaO68zryeTpqy1cXO/mWgSD/TnECXn3BQQpa3
hJlqsyOoRLbvxqYsgJYP7vvBAdaaucQ8VBFSmiNvKrE/OJhian35yNPlC1rOTO2yVvd8sCcmfEVK
pvu3IzS7XvQbCts2JIBoTS92QW156IT22rnO+DeUQN2aTVThoYq9d/XF0hFGRvv3mpk6O5rztyXO
SbsS37b5/VyXjcVY1D7L6ACeE7oIo3bE8mvPN3B1XAc2TsybiGHMTK+Qbcmizks2hdoWdHmYbkLt
Om+yby1bLdzM7kdvdY3poG3fVH4mTu+dB/bjMNow4FfJhMI5l7aDbnOEbrGQVKWQQbo37ako9Wpq
w8vNhI1ZTCGZNG6eCJrH9jyrvhS2S/cJdOLWyL9E8ak0u3pDwUnbh4lUL8ydB1WN5erryx5ZOQ4E
fEEqfW9Qq8FK1Jwt+AxAIWyP3lseQd7vMGZv0Rlcc/5O/JJGpSyuwKtlJLmr++l8kVP5SDIEPENN
PMWWyg39ms9zoMMgMI+8cAz0YCafkEZ627kNiitqeqIcwp5v9rzj3YTh0IODG8zkqA2rZCxVgv7K
VVigfp6etNV9hR5KKYy/M5rKZ/cqTT4CxjO5rwIelp5LRm3etZQm6p71OA3CukB1sC+s+YNPZka1
cZTwCfgnOhMApckmwIGnx7r3mviUjSmygJTxtmgm170ag+Xlt8JC3eP+CxqwxYWSsmaeBTAd+Iua
fgDQBRQGDEVyU9shijFTbPvabC/KSJPkK5/Ncbwi6i7hsITE6KbgGrEqm120ZFIosF90C3uqPnqA
RmOLx3Q6A2K2klhEGSWQjVQqTs3srXsGnZaVUO6sgXBIanocBUmkBWeKNmSeRraail88yGpuug8o
oNv+dTLnQnG+2apCMNJKNwSUssdpcSLzkxuhRRkODvxuNIzKih8gqj8b37Z+qCuwZBI7B5sD6Den
3ppRVH+lMdiz+Thdi7XQJ0sL2bi7jyuKbMnqkXr9zjooHq5C3qgms1NmI3ZMBwS53//hFn6rl/Au
wG2h6xoSB3eHVFv+trY6ZHE1TfTRhoG83ju6uHhlCcGIdctQsFqcSK6GQgxdfu3pcg+O1M8mAE2b
m2lsyYNjPlC3ZewKVI71PHlleq4jh8TIzgxelGI/KX4xQ9rvl9ufAnjHrVBeqAdSDwI76eD7P28V
ZBUXGYf7HhdD5jz0D0vsXDdGS+sqEEq+2Jh+3KsP5ZeWMZpb5Foi8wMECF/AcLvEQZlKOuC3Jz9o
tETp+Ib5/c/FYxWn8scOpdlJHOToi4WwsNLVaixpPIJVzIB/yTV7lrpKHbNB9SwBoFwWk+SkCjCR
xVgw9dHrkk9oZBtmXyM6XekCIM8XhUK/F227ZC/qqWyOrw5fk6T1fPFId4aOjii7BgBxHS0b2zIm
aArVSShL/XNIfc+uZ2hPiOMy9TVRbASfG2JP5lG+TbW3AS93KwcUmVWdr3K8Vq9jNuBEqmPUbFIL
ERRl6eiddSdO1KIfyk73gOBTVKKwYDTDRmtoqzUfuQP5rh4rCAmBk4Fvxz7kETJzUGxm1dLFBTjj
RvuEKZfbznRJTlmq3HQVta1vFQWqHyv7ALsCF24eRoKoAc66I+G/37hsOnRnM0wdOMHQq4XR3vON
gDDt0eBLIRuQ+B0Avb80atEDrAbGDLtE212wP9ubUw0o5kwkvN/GbqrdYoj0y2gxLrPZqsRD/Fdr
0q4TA69mvSCc56BurIF5ifcZoCbroNbGOqR7ieA5ANPBEp+RvJg20gFAI0m8mO5usZkN9s6Qz+nl
gtoZOZmL6cTe9uJWt0H3J01iRMU9X561pIE5IC8H2UEholYqk7N/i9UycXVNRmRgzt+QbKRU3XrT
dozJpgKhK5nuDoEZFv8o/pOvcTvQSnVTa46gENo33zaVjXidSKMiHhV8bUeTQRPAa/luIKj30JoF
S0oV6f/XDMmiCJ3H0jND4LREJqjfE6QAYX/EGW7w86fXempaUTar0/3w36033XSnsjsvieN0cdRS
NhzdtEwiyeauWTsha9J5azo3Mtmv+e9W9oy0cJ2fD5gC0mQzAZcOpONHxne/oXrAfrPKf1TQ8aA2
tlkckc7Azn+Eyoa7BUON9QyATNed4GByyhurwRP35kjBi52K2NUWHHjTelKAAhShUknmpsKzveGL
GLtOqBJ2cZJ4klZf18csp70Lz2MAiTAsNDuJ0CWGTXYIX7vQCXwcdQf1RJPt5gmverqblOBVWW09
Eca7ufLv6fNrG6wskIr+kEZDLYLZevViQNsfOcALpB6ilfXxuljhnjtXblsKenAnCIf2HaY7y1UY
LADUni8+Rpi42QhrnWXLLWhoB9D9efRHT4NCGGmsAROxVTsxmawMJEALX/X69wGSmHeYo05s/muF
SdIS1vHrzxvOHm1Uqo9HSR4sDPrJWyOEkCIrrXm9Fn4EnqXNz50kC35P+LD8NUqvmtmHNqAlcRCr
8lRR45FPZglK63f1O1WBBOaEhV4Mxqi3OcrYZAFus9hTONPv2/mm8SexKvtsSmYEeR4h+vwxaSUc
Bp3iwS5wimbD8RhOyLi/kDbRF4Jdzg/wKV63JaeCk2qThVwyk4BhX4cpPqbvuCTtlreeO5zfZGGk
KdxgEoYI6cns/z+DqrgKxIH+E0B/c5OXPNJGZCaHKCoifWsfQAWbAjezPmMDBTqqSLULr/BryfIn
JX45t4E//yPnAI/OQ0ybTuyNX5tVsB9PO26MtEhJU48waNJN17MmNhzFPI7oa7RHGr7z1XmRLfRq
auLyTY+RswgMJcJqON+SHY0HWOY8Sz6OAYskwBjPYThoCVcAkhOK1zSN21i+/xHnG1ypgSe9u+/y
PxDmfDd3gp4FE3b7RfAISMyGx2DtHnecdOvlOpk2PeQVafzNQMX7CjqV16xFNnN7hrN94ztTY3Bm
6FQKVrDU/uCuw7qvRJyz5bdb37EHckl+0cYRuc/hYIul/hUe5xqqve5PmQIzPymOU0sU/MH7Ms6j
5x59x5QjEYjNTqBfbqwzsAbjb1v/V9vTqBeRm0bBUzrW9Marbkx8Wtfyykz0pjOzAZesOf3ak7/q
hsklAGmdxqfZG/Z1SeqNn+QvVjqWW+u3EcnIGCkRMXkcG/R3IDwRKVOq30KGkxLCUccuZxAhFyUy
y+98pyhpYRzuMSNHM9gMm8ssYdnQMHSZGfJK4To392WAB6vE6T7r4Jei/TfPJ9JQSjuWYnRUbgrJ
6mgM50RUuU0JIFwVOXP+pj7YmtND39Gp/HaIKmwgfStmkyM1zil+EVplYjvUu/Z9DCviqglCY9Tb
PgEF0oJZsAq0K/V9fNClncLRnJSulqPLnDNnMAkr/a2o+i9luruVZhF0vRTTHcydHkGpEShebol/
4HFGbOolHUb4bOSiVYBS9+QxSwEAhqmiXgTbsv8DLLi3bL8VLY+InNghNVmsKgii1QlWTHEZm2gb
l+1ofoE8uGmTWcah/lVkV1QLivGJIt/v3Sm2aesioJ3MrTmaNe17j/QwS+ubK1VgslVMjygY/FS5
FdnYOU9YwKNzBkaaP/uJhMS6Z+vswHtS0vPWk50fJui4vmPc4988phUNETrwIdbR+Op7gYtF3q6C
g8KIxxgiXege3/KObSLtNnR31LeDxHhzAvhR/c0diGDHfJMqRghw6fVWUL6WX/9V8fhFmR1V0Yr4
EixvgDNdoBBcaHgSbxbPb+yrxOk3dZhBjV395UMMCcZolstCEPhxTD42/r1T76wfYVSdntTGkrTj
Qek9ofg61iieALBPFnrcbWz2cKNQFMGnpAyWmYBMSOBeypIgMvR2cN4g3VP1LGZyUrDwxCJtu6lR
qwIOQhZjwAtu0MT58CF7RBQXKk4fW9VsG8ffvmANk8AqEZEnsqFkz6EOxJt5RLurkA1Vxn+x8KB4
q2//w8VLUd5lGnx9bYUaqPCPIk11NA8exHvjnhz8x2ikf3oBsWbr2YYfFylfvGgs3T8YN55PfHrJ
455SRRCEwNtku84O9AZS0FElxIH0envwP2ZRw2G7I1mBym/y8mmDnhn33GcQFMR2PUIErtV+7Iuk
l+TKBW/LAtDty2zCYCQq/UMqX38nnYZKRMx5z9Qi7H1FzozK2QfZN/2Uz3e3KGuX+ZBuuwxt9qd7
4/TH2jA4bZQfO/9M+3Ux3nCMNbeAojiY1qebouvP7rAQKmEYhuY7auaWB1y1stm73I9HKsZdiECq
NG/0w1uD0rL38sHzywGBGlgtIBgbB0ge80uQHLkH8+R9R7zYCZsP1UdLDiwLluT6YJVH6VVwJ6bb
IleAyurHCn2GPRNSZ8oKj8b7WA3tF0FrMxz8K3pvIjzJxyEq/pp/6V+Ca3ObHhXUtA9QsV/e2f9W
mS3TDCUkpFOEY2YvebKdztCWTKOVIembhdj2L1DHJEUpe13kcHf1Vdr19tONzW67yxl1866k9kxt
y2cMLwxhqVu1rusx/oqjFYP/V74rWZPjDKMTFlQ5pdmjYLGZgfkyDawefJRk3pSxUX38eszwdJ5E
qhc4vJIrvA+q1rnqRP1bi25UFnVQG/8olCDcpUJwSke8YFWWmtIlWeUSplNxIvDySFYHyKcMXM67
SuoD6ptf1/iEfp0mn78ZRpz4fVt0EEtrKPGQkTHqQ8Z4qQ6QzJDjMYG8M4+0T+w8aCSQ7EsMKYM+
lcnzJiUNfCWoImoIr4Z4VgzY3gOABQX2IromWXy1H8geFZ+FQ4IsBuoI7nAS5OpA+TuCI+Cao9a7
7LU+rFurRWX74YGKoGg9N1sJetIAxk+xX4Hvj5xNP2+trS1w4yr+9oIlzsg2J0suuRMJ01URRh9O
DSP9I5KS5T8WkydHMgHJRiT0z3Qyt28xZQYTl+I3fRr0lgJtJF2FtZMMwIE6XGwNTll2QYfQF2de
o30SqetdEs1PiFPdol5vPPwT1QIWfz5Q1H1LY15UgcPPPjeMbmLKFESAmiAlR/tEFHyFfSc+pwpI
Zyw/oIr/gS1Vz5cpKhmqxQn0wKn/l9lmqA4Qrl0EpkRnOBjK2XM3LxNv73w3djlXYeQ1AKqbvlg/
XTWsUFEl/eFvvDt0TWW+zHPWiP4sNLhq9U0zi2bPK8gWptZpoptOoeKkO6v5Xy2JW7pCEhTvJ6lL
QfTyITAbGnoM7J3l+BpuKwNNxXeQvDagSLgTlrsnSz7U8zqcWyHR8QRJFzrZcIh1FgLnZcJu5PJn
P8FoUQ7dqeWbkyIDrVv2RwqsehlTgGLZOk2fWjm9zvwbUmqgB/poLLxVaBrTWNrnGBfMkj4Tm4Tp
vJvZJBCdjbCKnt8/QktbI04mWH4RM/7upT1V26EqmLecC50pNtet9uXvGTYl1+hNs9tVHi5+fxcO
opNraFjOScRbiSPJs1uUYFqMpDXx9hAfiWezQ0G+gsklTiehv2pdJzrVEz+We5i6Ta2O2Kmi+pKh
uAqUl9ElhghEHTuvOmTpAOY00cQjyzqtTQw3uWFqC+W1UYNf48k5u/IR0BAEod7+nfgdBluFzSI1
FFHE1c7IWwyN1RHnFd/YCVqUWFn+rNHXAvswNADFj1BOi3hAOF677VKWQd6f1xr7hntsNVnGM8vw
eeNc2HAB3UE4SWCOVTdfMurLuf1HqEmE96l8uHT3X6DWQ1nGYYyGwMNJEhsW+vm+C/foOeiruM2i
SI6Ld1hWy2E+hZZKYAf+/ih6ZntOK/vBmRJPVHdSF64fFMlNhAePkRWVq9Qx1DAnEkvEwl/1Ltmw
iLCnjkCMCN8D8vdSH6kB5ljP+9QFZwKgCAXNT+I15Pf3admlYfXtQmmscBKRHY9+e6+BUwnhLGhE
+gDdywKKu/jMTK9cTy3E7lWZCp04ZdkyERGFbVp7ZGWNkfehAEuve2daluKSTEIkpdc3miI3q1oT
Sm1ryc+FtzSH9/FCFe6acLCFKso2hDcqTYIwcsVS6wbMlXnGmF99AinXEEbldCQdMTA4bx4Wk26u
wmZ5+/neTt8g1GNJD1y5pBrl3hk11kYMoSYTt+zVHTLdsEw+wkFDxsZ3K80gIi6JHGxuboNUpttO
o0PwV44RCtDQ/t2oUiNS1sZ5xVXg8KlKuNle9Yqs/NDwyqZJA7kaedX9RKhWUTQ0xRofphZJcpNS
yKBMoi2u5jhx8gZo8yd8Gdd3d+faD3cP87O2LD8SjqwKPMdPa99SbIWDiXRw/2GOdnck6jT+UOL+
/O/zzpdgBYvz2RueEBAt4EKPJmr97nLKEW6sSZOi04rgNBzP9QBdMDgJgOk9UvjtyVGfXMUFwgqN
FccV3tz5QZuQSaBoPLJHLSW+tR1gSeQ8ette/ZLVQI1NyfOBs610PCtaYjU96+OIS26FxNHiOJTE
wC055gOP9zWIpQFVppFn9wJemgy+4PR5nQ6uSZS8lak4F2XgYB0WpU5/qQYPOplkJKbHBtAp93tL
PG5sSdr2RNsJaFcrrrD4Njkp+LwU99RzXQTYw3Zo7CjPHaQxTKIHDJFQ45znAiQV9I59dWUcR//T
lmxjiNXdTgvcjrhcEyNNrOglM6N5336XZ7JWs2vMRfT9/jB4HHv6/6S7CuKt5rVortG1OYCLoCG+
8CAjW0AKlW8Z4/TL9YY+4mYpAGSVx0qaVwUTyJZENa+wT4SWXwl+EGFmdTyKO4zoXBZHga+w9u1Q
VvAXWqpgKMIQhn1lf8d6q4UwZhNKOCcVlIrK7IeDSp9Uf2ZibLfdV9i3dD4ZqKPi/0UXIKqSqRhy
NVYk5ZwvhZ5FNqNkCXj88p+U5Ebi5npE1vIwHYE557Ihx9o8XuriKRce5pKhBUJNJvoIjUPR/QCy
2KLUE3o1o2pmVMagcKG02F99dhbAov2UaOtpkK0DDouo7atNyfBp2K/zF1IYXHDd8NEljRq7nq0T
McamymC/kriVV4dd1EWj9D2HyskCMRtpNRMSBLnN8iuNeQoaL2KGY/diHq8aXAcnWxpytueA8Ltz
hp0ZzgXvw/7w4fmRejh8oBx7rJBciAV5zXRisvw2jRFCTBvXX8zqeSDz5RrhhYepPWZJ4QW5Gjyo
8sgO6fgg9XE+4/Yv9nITqaYaSu2uogYCYumqmyqqi4gFpzp3za1nKNTW9yTmCH6Q8Cw7Qls7dlT3
IGpfQWJWxu/ckav5JhKfuIVa5qLkJsW1yQ6dHD5pqbCWS9eTNUUNbNBuSXunEg3CuxvehaF3+jjJ
20LJctS8GfEbLq3+STyK0HE3IHvhtgc1REkNN8I3/Gdpf7C0Ee4IAe5zc/sgMZEQOjceIybpzXHl
5vB+ILZBuW5dMZqLRhmjqShV7fPdxY+kOdo6u6M0oZzpGAZxkDxRoEAQNQ5COWThT6qvd7XYytf6
n8aSMooJhZoRe4QBmIFdciXWlW2cIAvwxHt7/4Z+0dZ5VDBRF9qLfARPzDk8PZWHQMC9lkKJzzzs
Vg+VrxlHFhSbYLzT/kcbWrM4yf8UzzQ6L5ZN3WNUBgTbns+j4zwX7iTzdNP5xm1Au77G5pzAQzA4
z/232f04K4r+lAVb0mutTph6vX3k+ZGigb6ApGTOE5Dg+2FEUMMcajDXd59i0EE8uIC+SrWRnhiu
76J6PB4k1k00bi3hk5JDG4rVflJHbQh3HptCdLyR5M2Cw+ZsZ8Izj4EGmn6H4jaCjZK2qlozijHh
aF/1GVupMXQo3pFsgcxZBL3CKWr6xPfy8/1IwCRxXf/hYObUU+XmQ3OGBVwA4ZKCyJI/4f36fIjJ
t09DgNIx6hRPZ1hHQO6evDC2hQornPRl99F+5qwKtWS6jm/ozVHbnx0k67oAxPN4voNw5apeLEUJ
+TW6a+gpIkUvoOQtwZ2HDrzqD5PHt5EuYGfGG+XyTUCWquWOhyF8eYdUrMCpBRBft9Gr6PFWyau3
6tWUxoKCAMLx8Pf8eA5pUkZb2g0HnhuafKZmVcci6Y3/rYuKvqgyqZc4pH187+aQFvu/o1etcYja
g6Ejg7LUWR+jeXQTUWOVM9VVq33FZpLE/UkcV5sbSquzGbusyOWUXVyHPe6/R4+1Iar8mtgAm7Xi
IBa8cLvMb9s53DOEuW/EborZeTiH1FA4AMAJtZr50lA2BMHJNcFLpM3PpwaXV9Ft6VTp5ZSRX5Lk
JbO7k6g6IC3eE3niycp0WZoJLdEaVrtM+6jsbPN/sfja21I95Wjf0ye9kqaEdHPBrfqfRuTUzVGR
9OP6ZGIUhkupKWylD7MF57NZkhfMnbDDHoPPnHkQrYOVhI/P/8ahoRJNRAnV9ka9R29g7ZXW/FlC
zecCC+rV8h/sLXvqv9wZEN1jN2MPJqq3TSl3pVW2kxPw0CXsO6RthgSPEH4cQkteVL63oB5sjoZ2
0rpa2h83EI2k8l887XbzJA5fqpDXpeWxbS0mzoCP5ZxLTmkTI1J/3JBf/+2nLUq4623koKsbo1cK
ipkBnK9VhO/xLoGsRBF4TDg0fpBDAk4ybMS4leYlrJ1H0kN1u269b/f8YxMjZgKyCQrqH7khaTXi
3Q+6y9fEFNPLZYDuiSotOp0pOR8GycSWC7GtMH8xTtm4RZhGcL1D4OEzSQa1B8EBkSiI/Z7U4n2y
QrkvQuvuw7HRS6VgUTRab6Kkd5RcH8AmWPjU1oOy1FzIej0lHSxl2ksxsSsn5PcSf3stTUZjqLf7
0MFiS+XCAPKSudreMzZ9hXe2+0k1uxF1nvLwtJMd03wnvNrn5DCJEX1TwJvfJJ9T7kLNDjh9iOo5
W7Qju0UMGSu3DaLVt98tEzDKRhOtDTk0ARvywNv7NWjAeKlv+rGSU9R2DspFofl/4no4HKmOTK+S
RvcueZR0bT5IqGsHs1ZW1rOao5R6iuCPYD2XpdZV460EGbH1Hh/M77jwa/XaZT+cQvmdZzklZAIe
vrMn6z7C+m9d53G6YGCV/hLxQQQSjotqiGvO/4zTWtPGL1SRS/K7mzMeEVDOQgI2NZHiwDrzHpkR
Qp3M/eYYQYtP7/6W2vtcT6TCJJEhJNLbDhlZWMSqsLjHDETR/Y69lozi8bqfYiv9yzhQ2B3Jseh4
C/nzTnA5sqXp67o5+QpdX/+dPNOah1pNR2lLrgyemzuOJcEUWRr0J9qtUJqdVKci5UqP+8XKF4X9
a73sI/1d+/9nwKiqT6dQ2IMCdaHfaswplFI6CsT5JSsTlBDVhH6uMSfCPP/mnR6ZKU8FXKYbEIhQ
XSBmOFgTYfOLl5d9gBCl7+8Ri4/NbbAgIcUR9szFAUYijVIxhN+Ey4QGFm98dmLlE2Ot8T3lSTXC
URXskdqvGC0OuFUYq9pdLvx+FsND8o7ETK4VfsJ96cwrNT0JVVs1cDHJMCScMwOcjohYs3U1bv/S
M+Vy5hDP2VUi+9ECeT5CpNzgsk1UpB6KAKxrhCMFoSACdoQM2+fbHKYo/W2Gtx8kEUiBU1A5UCRq
Oi3x8ujNEAz7evC8IX3ZN2+tcOVXl2dHHpMli7J9AHrA3uCzVXX+gshLTWZxuR72OF2ohzy8GR84
18Bu/AXiF/lqptMzj57mIkH1rwbLlCg9CC+jrEdVQ3KUZ8NzCVoGnm6asRooWsBH33RlkgqwAxLh
6Xq66eXmHnJCPLBpnufoxtxHhD21IgqhsZELaRK5AM4Zs3I9oBdVy2A3GKshSVvRKGCokyV/pl3M
CZKc2HCtOyevRDC/y/Wj5sBxU2gti0U6ks0kdTeBiyTxvvh2dW8FJjBMrgD/B/hM3oJEMaCyhWw6
Hz4iAOjAYIvr2DvP9x71DhhJgl2FupBv00bkJvfvYB9mH8ge56KemlSInMFud43uhq+qrgpCUGBT
bTvO/gLCj/R1l9gbuVokeortiowMviIO6o1zII91K+N6sa+oK7uREfB4USiVbWMSEu1smhVfSZJO
jqUgWeFqNQIcF2GBqoH233TtilhfzN6KHPWxNv92hWbQyA3g8Xv4zGegDBUCQmijsZrW3eWxgZLJ
RXPJtghDCldOrMRVzsxuKDy2FMYlUOeyK7Fv0TLg4EfYcdEUjxZrP/QTbLayMW/hHpAoTsz3wslS
VmplvX25S4Ykxz4ikfMrVP5mtD1+m+XrJwm9hVnj5m1RKO+GxKCMfX+0uQ2RQiGXeG43QJeUvt7k
WF4zYTXXRA2R9J2Rs5P6p9zClulYSJccsbDBXJGVXe7w61UTOjLSKYZwxu6BEk/VX5r7UGbPhJdC
Z6NxEzm+idu1ER3mF/deL9PcCjjonRhyAasF6QtEJg4SlF++DIfA3zMZcwJAig6WjS+1QVk6ooM1
vQM0CmC6ujvbovHYSr9JbYtwYDJG81MlaqbNidDoWtdKpz2rWTa1DJTWwniCBXuRwO3APLNR6zi8
Gz/kFdu5RnzSKsggk5PDL1geimvuivbPo/zgJWF7va0NAnOFHVh8JC9ZJtwc5EISzpKcK565vwOM
Et32gnwF2e5Y+7kwMznB3k4UDjaG53iVW0gcOtA+FnqpxlfSc8T2ou6nHRAoiyIr9Qn4XYVpzqOn
qrprLAbDS37tlCt1UvvJVFDJ6qL1zkYJZGYj02WO+r3b5bwAqjAbaR53jQoF4GllBRPlywi3hNUP
kiYKgSDn2sYRUywazieOuAkOyuTvcQ3EJfpHfnbG1EXJb7w/PSNeKbb7AisteAS53yTOzBgckYTJ
tZhZGxp4KsZ9cV0Tsl8MGsNWcLVEgOnZSopnlKRYBhKvkq3BKRITgkuoV0Vpf8/oPHnRQV1SUZE7
SkU5xSldfnDgH1p9wZqbRPTP0s35iF7BzUOhCPtNEIVkhZqNPunrEnaXmcvRmr7jxUxt/GhkmCmg
wImr5BMPizhyFIOZ1ZTiB53bKx1+lzQwZuE5DPI58hJW6KIkwMtPIqeHUWb9cpKOyPokQlWrpeN+
/+bUn6Q0G/VIHIrWCjiu6T1WBBJVZvE+oxBALyJiZ2LieFyH4zBhP9nQMxhKHZ24fnC7b8Hgg58M
PsFuYykloZASseqzy0b2UHE7O20XGtx08gRMEznOTSu27/O5NV2ALCdSzZF14mVW0zyyU7SSaWzJ
v41+lv5fYFAQkQXI3HKNTEWkhdX7sTX1VBewp9vYuhxC9iMLkFascm4OcsOGuX9crq1nBJan93Ba
uRoiEOj7MZbAOvBBuE1F6cWh+l8qHEFQAlqkljbxE8rzVrb3OWwX1ssJwsBBxDQu5Wxnf/fKKvSq
hdF02qMDQ5HQ/MguCtw+bu3ZZqD6TElue/5eFc629QVzTYsAMIvL60upmiFncjtIHD3GI+yg6O7V
KbBk/3pOZX2Bv0/QzIg34czyvFHpjH2EA/NWFech5cjElLPxExtC30bNEc0AbxDilvIVCtwfcDPp
oZSV7tAKzI3ptD9zY3sBaW3TidwSV+6rjm8Um4aYn9InYPDDBKei11qBrns3Dnalmn1IF4YDDIad
HPtiSAp2Bw0R4P0zvI8G2CxFwH9oOgVOWrMgXXY/5fQKg95RSfbY1VMtDPeTMBVth4/wSj+pXEMM
0E1Z3H0pHgsw6Bcd09YCt/0m6M9N2c1osxno9+Za5h0FiiX/kauAAL3n3qPiYAIPl/nVTOCn6lcb
WS1ikUwiKXgrrHigyzlr6pdNlMIcexvhPpRMgarfROv1MBVMpGlFKkFqWeZJiRhpljXHL+PeduFp
9yIsi6fcun0+0KLgZ5CwpIZjMC2G5061yYV1qH+zqvFEBRss7FJIkS32bAIKiUFfBkhLeKqlRq7x
rhEXa/FAcb+WDSpoKKmnBINFCjc8WNlGVczz0AlFrzbM7JaYH11+LiZFbDWpFcawouRGPubSeljZ
5OGrXpIKRa5/G+ivoT/bXqYVaAYMb8mpdU15/Zx2q/1eGfSP3gtKKe0tepNc5v9XEcDuF7az93+S
8sn3Fs6Hn9MRw+k+6YZJA93RVBKVGg+WXIqmsV3B2RINgMCojy+PJYDK7mKePh0jZEOYj955PV3o
kp4qHYLjw1hOW5LmqklpLeegi3+Czf6z2+UfbQkmOlDKBBK/hFUe+r4ipU8hhOsck3aB1w8Vm4lE
2O5ZwwSvlMG5KK0mO8Fj2/vq1YvZW3MZUCDqWhxZ6MUimZNPp4TJSkGfoHXsUXHWqIAMPMkMYWCW
weOIinyt+WWWBDcN1XL0cuEVJng2bnlWEPRWm3XEHhpQ7D+/ockSTV7AmgfTYXGIYs8tG6jVDzTZ
mKf3CXl39JhTbnIHdhSL+Mv5aqXBK0k9X6HQjnXzZWgxa28369V4jk4DPGUgUhXu6GXBC8J9DjBS
Ai5ZWBhCBoHOIKVxpUXGmtJS+8VC7DBf2UBKCwHs/hopQkzI3uyhravrilUUu3j/f/PTxvSrXc03
wY3fChKWWvMv+d80hkk49ASdkayo5JJlX56ZrW7VhquefEhwjrPBSDWvZurvhhaEp/9IuH6P8QPi
bOQCnFmZiWuj6V3gd5AWwi4Ar0eKCLV1ObnoOaSm35d3g5YFYmFuvE50P+4MOWatUaektyka/MKt
YMMQz2y5LC2sQx8MobrJKKuXbDUBP0DhPrAbX3fJX0OCq6jFl7HtPecmw+4zqa3eiGSqDvcczWwf
utR0+F6UFA1PqUdzHlpySMl3JhqnRNne5Kk07kgtoL9DHbWH9bOTbK+XuN7Er78ifO7oymjQzZLl
vGdjzmGyayP2qllomaA/+kP1ydtdjsdVFl03O8/XjRteUT6tqSjcwz6eqQzKe305/K+qo2PtBc0U
iiOqF64FhZnJyjpJRVGzP0W2TqChQjZsvByn4g4YuicmacX43pFJJg1DHCogNUxsg0UB5wQdrqMy
x9Xe7VFpTiZz2SgsJr5GunzHxBKDQ/4bVZfidYjfEQvvvCJBPqarYP5t4vuqQMaSp5fYoHemvH3W
gTE7YbYoEGbs3gCJTx+VYfk09jjcJeEhIoSy2UA39eHhn1gT3IgwE1kvG6fey5uwQvYzSeMahBRD
c1H4R4fy+/qWij2jeIROPvLA+fsd7xMiQv/4XyxwWM6qfq26paAe/gsVwvnE5VvREIe1VtslX8D7
5VUYT5uAGyMyL2KMVklDUV1iK+eL7is9BYzIGBwlem6VdhLqNmrUznyr3Tut9BD0Ryu/hujj/FGa
xHusEFicvTspRF75E7c3rv7UhgZmeT6/hz3BqqXmoSqswNsypdc4RGhmmztKJJkG6gUJhIntMt1o
zmotcFhzSRoJegBXhHfBVg/G82D1aAEhR2yqs7b00mDFJaUNTBYvVwcO0wqK/hVqVCxD83iHkkka
3W137YadkHHulluSMtbZn60PrwY5KSlVreCFzfQ2Ep2dJ/gnifnBAq4z17zit/KumxN3sgZwY0Ow
+yX18ldOtJBAdAV+lV2lPWVh0Q9TcSwyQr8IibYDrpKFScCI7wwpWhvwXJXSP4Y0bEwMWCKDyGKJ
We5rdBxEx9jFLUOnDHyiMDTTOchaLsV2p8KZJVgUMlni4reSCR+CvplEV1yFkEMiwa05CZISGMwG
4IcaVVsZRuRp+MdbnTiqBb9GFUL2KyqmPYw7Lu+4V6F6EUnHl5dLv5vm8BM6mgGsYYXQWHDlI1wO
v6tp5hXv84ohdTBjfFrc7+gBFHzZ7onMmx8m0MaUOhT+EldClyoIbNlemB/OewyoYJantXbZcHWD
weMlRU4fu1CotIS0jptwZkDnCoRGQBxIt2AizC0ut3y+mmkxzWZTAFBNe86zCGZXBJGIsmg4NAlU
YdOPM4FC8d8ZLIoP3rdkkeZQTZijjPErZHYAxg4TlAL4H1YF1/tFQZJkH91uWuy7XoJo1yZgRhUQ
ZZ1tX9YPoN8aV5H0sx1zTWOKB3qrpepnFc+BNuNmDPlfvtUAFAGf4ESz8fL/JbO4H1fYPxktUrVP
ozDKIpEXQ+CymEtlYX87KhBLUqomH09zP7vcmCAww9SrHfOWSarMNOd+ldOskNgeq67DYt8r7WTN
mMJ1eSyQkoXkThgiLTBDpk8g9RfZ/EMzmeGNTyoGvyKHlCpY6512q8UbhlG0dATEdDMFgJjfO7AL
bujFOWAf1MblCY0X8DkN1lJ2xuDwgnFabDjqZefEb0UXwyiNw/HV9plzZxLJqAfSXw9JMh3VJ01W
ifQ7hVWkSmeUB0oxS4RbodCI75RUFBqmjwSC7IQOz0r16wXKYA/X8C4wBIxImJ8RZuxKXmc/VZiw
BrcnqUmLFs2+RgfmmbvNPd/2aQdjUzE5f+yAVNG5qxkEkbOp6r5RfrNRF20VCFG/8Bb+8v1tssrH
yuVbdEjzqGcnhS9Ur5tDodoeWjYElp13tWz76VptgdFCJu7z1EC2SWl6/tA/QVPvnLJKm3uapnFa
xHU5iDlVVi1b3pDqmbG4qhusMPe+/mEtxb9xOuaWeZnbAvCKtrj01+0y/FL0Pa4xKzFxPahRiLsi
eaOex/OfHIiotIrQpWzj4a2RUkeMkBt60SNdLAen3Vy7CbVPkuOmZq3JJeZ7NQfQ9OH4m0qGKQ7W
+dJLQUmYGRA1vHMb0Q9N/lI379ZtfCRucYVbTAq4b/5vfmylaH2P1KE4com3OnfgJLsLo/KrZJYH
U1Q1FM2rrBT3zmo5Gk8qlJn/HqFiWlkVvwSW2lddU/PWoXhgPmiACBvJ1yKFPMX2Zrr5PimJcMAW
dBkV1xZr7mVeWt183GQAyXUtmMGj+TQclg3aycwGusoQtVrLUKB4gy7dqmBdWi1v+HTpTpzGm1Gs
n9/IyQgKDYqzIowoWGMswKP58aOVJT4oFh1wz7T6/FxcFRYACUV5XtdsbfvcJK03OvoEcYvXoUnQ
uuHduxMe1NsKoBkcpA1ATzajlI5H/2NzM8Xa5cMDhlakNyw2BQlBsC2qHVDim2l5K0fKoG87UZKC
0X2LmyLHZLOYDT4rolA4wqtw1M66VBWQBCqpTRevvlLxAcoogbbY8X3CcMi1J585Wke8SwnqF/iB
thDaiRJQ5exhuiFD5R962Iq+ZG4Pyq2iSBZo4ilP1tIKF9yCP0AIT/eBMLQf68lVwW0+0LPTCss8
IClb0UmDKyyMPgsn0oY8kb+9erO1efxVA4EgyUaahdms+ZehKrW5Ng3meEOAxhWUCrOXP0NZUWR3
s0A98R5/lV/AXduPQPVe/v+Qg0MSHnqNhahSp7JXZXn6Pu1HfV0hjQ7ziQdd71INmT8KRl45dgm/
KHYa7nqUGIjAcJ1cqY4Gwel5SqCmbcWksspzTBxV/WVGN0dssBSMENDKvSNC68aOvSTOytiaznQk
Iq2WzRDWAMq/j/E2bWzSTxnH04v08RDs1d0j8Yj5ij7dyz//KO+vRsVMH/NjGg2G2+AwFmdN7kyg
6bJ4yoSqN+syWKzc6hxiUg376jlifWCO5nZDXSIJkFtH4IUZyBrgW1jWplbDkMjrqROUqzfP4K1d
+sQPnGeek5XdZ+YEv5cH+3+o0VVqwHuV8BG2btKTuApjCrLoxgYg5nrB9WwqonlNZLCzoR5gSzs9
DYu+Fh0Kciqi1ycoo4YN+ObnUIbbBUkPveDQB8bk0WoBybcuH8Abe4E2N53xtCNEAvQFE6H54CjE
7r3xwdUYSe6fNHLHJgbTC9ppbBU6F74wRd94mfkkTPf5tKY4LF2553pMcQhn1dBqGaHcmI9wwFJQ
0yEwCME1XxdF4htEHFVRb2bTxkQFfEeZIfuoCQIhGJVPFdQKCDw/FPwriZ16L+c9fqKmJzhWKYwV
m1BnFGKcUnqAcGQnlHONLXL+RtoZh+A88Cj2Q33L/rD2aw5UoPaZpv2qAORW+FlaBnXzjUcX/vBl
OvQg9GTOywiVQDpwmW38aE+SXYc8ZWBnmoyEkYS3IWf/8X8xSj/zgSUnvDaKqNT5B17GsUX5+kQ9
iUZ3wdo+F0XfCODyJqe2zFqSusWDX5rHqBF+iRmo+s/nCT2K8UjeGr18a5SyX/wxskiHUuuX7919
GJOK7ZA+pl2va7FdVeysQwALu6bHdtfRt/2TM+mHFSzKilaaYBAWj9RF+y0HjaPYgGR4pmRYGC+f
EbqHVJZZi/dMPNVVkrF3WeGxzdB7VzM/ZrwvCjvdZ9jgG/xI/igTWZWo6EsUskaggJI1Ub8/kqqt
Y4cYU2ZMBleS4aU0nLxUUXyiBl8L40fMbQlWtToNBmI7LuMVpOUc2U/olQhXYvNqFUUGauMJcp06
VgigCMJ1Jgb0xpBEvEkrox+lG5QdmdXTyqmk/y9D+YG5ms/PJTwgv8VUDjmqbFBbTTXmeDblwrEa
0Rrgtqe8+UpjNNLcDEapL2AWG5hKQgLvhtYTpg4EINwdOZxPONDJUQ5nwRjrGnZqvuETMdWnXyC/
tvIU94ug9CLS8VGQPsO01yjzecoCLUBvhxDO/01bbLK4c+beRPid27wHo+rLy6wae/wmjJjeG3au
ldQmQljGqL/V9WGqxeZtngYbpvlHhc6b+5nnKJGvNSxvdcuS3AXSx/W48ie4DUntQnXLPu2SkayU
TS7NVmDpMTUAc01WNOpIIYnjOk8IMiZtqjPL8F+dzCFrI3snfL7gagMPhXa8DwS9V03GOaMvlNnU
MKVQYJpKoGQwwFmIicL5IxfUf2ShwM/wIvyvDZq4eJyFsYcWqOkrTj7ib9abcgtDwQvowp4UAtPP
DPERhOC+jlABG/kUHwU8l232i+cs+BBw4ZoJ4QiP1r0aga6NYjCCyKHFo0PXbMFtv8aq2NdxRD98
jwUG6yZMcMW1XHt5TrV1QD5CNYISLkarQ155iPj22WTL1vYYSMvIPvV9W0F3pZtSK3ZNx6HJ0ru6
GMZZU3KFRPeiSValmBiyBpTMPu+9lGwPIiaY9i3nJcxLL9lOWY5W/NE7X6Vz1yG7EOUC6BDEjRue
6UlE/aQEbkBwPkGg/Y+KVWCadD6sP4JKMyZ8nE0+HtZByNSvnGya88gMYi7Lb+VcT14luAAVwVpM
vB1Jp+ivB5z3YgURxeV91tJheXtPDf5fslUoDhv16fVMI2c6hG73dsZbm5q/PSZiN1RXaf0b0Gej
dSszQ3oW9oXym+1OcdhDy8hhCFVELBSqpOCRmidcgPj5N/UwMStbOmxQ+13KHryc1cwgWArkUvCK
pVRKzeDh8e/hH81GrMW5FDAWn7dydV2lzHTlaiuR2SQJ8s8q+FqCYAotkEUpwiNGEteyGZnlEzDC
idVYvb7mBKsPea9qTDqh8sVINcxY2ExVw9ZtIyOC9KG38JEhc/filS65AX3okO+LQm4GE01a1D7k
vGUaNekqZjJF85jHci5ALACZxCjC9nuXPG0VbdOP/qyppxzDKyu8Ueb70aP+OiSspwoxeuwdhFx6
ocmW5s7fERwM8UFSDJwObzdLmyD6HnFSZf6ZZYAg6seakMzi/wsbPVVGTE2DcruPlvmsNLuIuced
qPsvwvVCjY7L3eRPpv3to/J9UEXhARY/wlcu0h6/6K0F69Y5Vi3XLKAONlnYIMv0IO/PzrrRXXds
ry07Yp36q27Fnmnk/ifPi1lXaPgLusZEi7Yi/aZcP9axzeaBmDl4KWQc6ilWEYhqI+Hk3GrDV3l6
5YoyWmu6fjZ+Fm8ilrdMzEiqMUhhkjWU8MWX4RRQgd6cgTDqnb8Zjon5/WV8o45UJ4I37oOMtM5S
Y/AbpV3AHznf6IYIXWVIVbiGK+GFHSuBuBkVYpbBBhG8/oo8fw2mdeKjxAbs4ianwuBcTgjlwJM+
wv3qOIcbhpVh96JV08IWsGIxUGLknbia3+jK7KNKV9zyK+2tzZyWjKtrFrcHf6El3DtUvZL9zlbU
Ve/694xytB5udHnqLsZurmk/O7sixCP8P0kCQQp0B3J2FoB+Pko7OFVrp4fb1tSb0/19tX37Z+D+
bqhvV2YdXS3J6m1Tf7DYmb3P9pRfrQanlzfTHonpL5w1Lq/GILPHxkDGY5PMdrUUX5qRld3GKUS5
RcjZJIlpre8AUHppPFEtQtfb8iI+oWTOYaffBtJKd2Z1d+8Y+MQJdWEKARL8Y5C10gGCm3iuYH/R
vuc/DUecOhO+tMoVhi1ipFqAQDrU6uYcs6yIPalXLIKDvDIq9cfgD4iHHpRPMnTyawAhbiEy3+0C
xnprzBUNdwrLXfsiJcPsi5FSzQy8IVfFYBwYba3lQq0NUW/K7XO6lW4GZEuw0uTyyUtH1EAT+hDe
k7bocuBkUFpr8byZNLL09n9k6+C9DafcfN5k03gkAf0rFF+3PIcBy3S03HIOKuSfcIq+0fWAOUWd
1tImw5aQnA7y9UP1Qr1pYKD47L36GpqL0k2vFon5Uke3AhwJIbIGKnZixwCFxseg+XYmKt+mcQkB
qYmRcw9FrVWm4tHvrQr3mWlt7sFjrBxRueWeVi1sWTmOmVVPF3/z8hNMGTF18W7a/zW0zCZ+kIfs
D23/PoRgtkCT9bLLHWZ8sD1Qp9sGeCF2B4egwZm+YA7ghHQpgooCvrR+OhYhPa7PAXnh7uZvy0gT
h3KxjOjkjszICvLTDHZhHNEPtA+6RMj91u67TBJMZ5YLBxqxIF0vWX1ZXIzFlo/s8i7RflappIBK
bLZrsNsFSYKYirfAvOgpYQq3NsTNTj4mUallFplNOcUXR7JUrIve7Ew6fUOpYgSewuHCH7Qj3r/N
M4/qFFjfWa3A17/wecBcHS87FaLHKDYMGQN3dHVaupiQdUQbfvj0u5nGS0sL6wFtGIWFjIooSn/z
aJSwOwIID/rhsgfjwEWI2WFijhj2GgaH0ecLBAZ+iqcMNzKK5WXTNARkCwoV5OEfHHkvB4+yB9uD
aAQ+NnmKUzuUw4A5i0yYxKsiRgugnRcpuLxowvNV9IShQtrK3TILWdw8lN9JHEP5zyfpvvbf7qDM
nSiw5CuUNHKuuhDgiRU7n7crHwum6VxG2GlC+bOfMUcqme9cfv4pGaPzMSI7N3qamuVci1OZrLQs
snrUPtnqm5CFAAqxIWXMaC4Ah6SrLC3ENxCEwIR1cgZDJxBIXFR1b32WQZgnKRLLtJnRRB8Q5uaJ
4IofjJ2bX/RIbOXOJ0Acw8KYBnWIi+TWAerbIW+ee+ZDjdchcWOMlJY3XBgL60SvWHdYoeolDvf9
ikfyR5NiSCrhdnERr0/S85nafEykp0JK0cPbWtONOnUBKlpJWTn3vAAUGcCptxPmP2lrFkDvbrL5
Ksbm0JraqFl7XkLFJ351K5aqvKJ1pIEgGk2Ym2p9O7Ylo0mo2YPeugoWKXQUPaMdR73ytE7467cG
iDa5mPGcD8Ix6EQEAoVgJhcQ8Kw29pLHKRG/etpKrgH68pO5ME5Crk75c+XndDGbZYwRhhMFa3rv
BWgCpsCKD2UfTY5zyHdE3g9bfPCPhfJ03uL3pDtvu3O7gCW7qAW6AHK/ReaE/akY58kcZHsxLB/w
6G90WbcMLOpgwvMVQVvxWAzpKDaeC2lm2ZRTxuYpUANcgSo/lmdjLZl0t4mC1kn1YKKIGDEOjjlh
gps/PK7TIoSoZVGM+wn24BS4+PerLu4/9hg4E0krVkB9QHU+JCi2WvWpelGE7OF/wCJZMVwdTmgd
AMtOXoIFaE2O5eKXoEu3U6TR++az8Yy4Efd7aLnqTxbBO2vv3AvRVB38SM0O4ZMSExQtAP2r6tFU
SMngWBGyc0Aywvkdw68S3GksYW47eekvIXU5spuppo2o7/UxVNc3147BVme04KkMWqEbV/8+bMHU
6wpgn+L1zSgJcZSk9Eg8+oCEjfrlZAP0EVNQ9qRm98R5dME5HR/eKQLgGC+6b3GleMRFp1onL4zI
tNfhx4ZPnpik4cuqc7hfKMdgZ0sm5sBcxVzeP+RKqoqcQpmVy81oJYtAS8cG0w+VrAVoxJ8q+Rsn
KCU3bJGOPYdTyfbtldVPjsfQleULxk5XxpKSiUXBtE6ch4EHtKq0H7czV5klNCKu5mjTMPjsEJTR
qv1YU9n+cKe5BlRA51zRWDvgzm1L+b/FCUs79xTA5r56LMoGpwZdfX2v4jdNeTKmQxbQB76AlY01
HmeAl0wNAXTftgi3Tv2H/TsCrImiLe8nW+LZ6ECOnrHt1/11VGXn2/+JDlo7jr9TotonJclu6HGv
9gZYe4j3QfK/cg+EUjtsg2usTuhSsbqkyyVBxOiHw63WVAwGKUTEtVuo3bADFAF8kFfQQGmyqqo2
kfHdW4R1Dwbnr7yM2jMQY8nHnatsMGwyjxpcdSMoJidTGMOJB7jFW5xpJUXY5E+JxF7U+uhK+4q9
CGQyx26T1maNtOL47nIMW4rwtXrYyo/Y2pTn2foyXK2j8PsVygWMixPea/W7ZLfApnwfK8zg3mxl
+T6a90R9vV6YhrWEoirMkNZqQpZ5migV+ng82xQ4pQjfei/rbyN8iAwufFAfiaq9nrOZ3edhg3Ld
fQN9mGsoeHpw10Zr8c/xlc/D013wCE1ZKcqKe8k9AeHhr263Swe2xDtry7+nPnRFHiE07U66lss5
PGm2ERE7wiXix8GjEZoX/+4egSBgJY07hrtVM2mDZur2OxHGg2NGQByK0B3AgSyElIe1s1CkYTZe
XMYIlJWPNTblCul7deTZKI/H52mRUtpJO3xrOcT+QnfvyvG6vqBnuERscGJMTeMEgxZIiG5HKufi
4EKiPND9AYH6o8PPY2KT8rN4IwVNYidzWV9yGpzUYZLeEacBtG8geC5/FsmbUB7pqQh+IuMb2HxO
k+Jac4X3hkpAOCoO0+RPTHciAKhbdEm9MwQcYm7yDYzLO1yxYVLopEKxrtqgfAtYYy6m2luJATjj
aGbWWzluPOFp0wUe04qtVni28uNDK5rPLiwM3Suqt6xWLwHfjhaJm9K598rfGdnX/RpkwXTJapSB
jMTihs9AITPIpZl/BfHlLXs21KCpgQ43nH9pl7l7VrTa+TFGecMxLZPc3XBANO/UNPN8Xd4z+ImL
SRsJTYt66nPkL8LBswVm5cx4CyUvvnL3Qvyyskj9fwR45sc4f2CgWciHaIxyJc8xeItPDFyEdr4g
iM/+6au5JpKcO4NiWy8VFME3IpE2//JZrRH9tYoQtycFDebP7xrw4gxphuzWauVBPWgQgZEgDf9A
pnnbu3sInlmFyTtLARzjGJoHu3D7PFlFI9z2Bkbxd/xGnH/Syb/5/z5soUXdxiWFcAMWbwbn678W
DuaRSwehj0xahyTbEDmGyItBMfguMCQ9Iyazsva9/J1aLWA+JLHZg/fIzdjryf286yzf7jUfxUZz
Bldy0JMp0Mwklsg4+kq2CWQfjL+WLt/FEUMaCqDDIIivdRsP5/eZhsgiZ/aCnC8WehUAcyNcT9Rm
gZ/g+CeBIlzcuuB7LeATJKdR4yhW8MZqcvvVr6ZVGAWJwawOu9Q6XXPRbBCEqKna/iHeNNJNc/Nq
/tfp3AlAWWPZ9FmbMsE4NXmtgAoZ65RXAgW4zRXszcELnwcumyZR1H9NeAOrHZ7cIo4N9c/1EUVr
BAXrfV0mSmYhul7vhFJ1cjcLIsO83ezTaYzkJ20JryLfGXZIL6JoLmK6w/1z5VN6hujHXooZobSO
lDOajh6mEyZXBlZcIB1NM4lsjz7gMbZFvxMT6vu2xAxCtBApu+oywKN5Gu7zfBYsdH0n7tBOQ7uI
kUXGB2glBnWDGzIk5zneimRaYbkR6nng5SL4OqIC8QxIhH7LulD6zAMkutMT4IMDMSrZ2nsaggSM
DfhtviIUf5ECtwSQNOkBKHtN+dWPwj/HvNfrj3LkLOfCIU8SnY2m57NhPfdpCryta4B9XErZDhuX
rDjpJ2e241Ae1T3UbQ00z7n1RxEbH6OI2A3zDQxxJajtOtbmFrBxHj/pnsnU8MOrcjuCvGGZR2Fa
ip20XqGQ11Lcjbf1JqhpW4cOuxZS6ntzvhTHuBIHZFK/icPEs/4cI3y+zeu5o2XYOg+2MIsNlJNX
oVf5aZpR/nTSRJhqZkkBxcotLSieuEvDESQXG9oOFzPlUHQ7aioEjTlJjem57SQDGj/c30FVNsla
Sc84cl8ERNFXRrLxlOdlDmQlYhDx/Y+9N/rhn3JP9uAQdiXNWYO5vxBOSGjqEyehpA01rW3K7LpU
PHrBSjpbJQEYyK8zr4blqHRhpE+PDIl/ZTpPW8IyfDS0LcZadqyjY6JByVg3lnZeeSB12cKcU2kq
/Wr6Cj0QR/CkwAR6Y7YLhUleZS/f2rr1lk8IO4suaGT7rZ68PLXMuPbiP8YBj2THnDBdZTeFVg4M
ChqFryA0DIgP04U1/niQI8YpoePe/3W3ITaM33F5ShgPphucBc3YjibfgSYXygGqqRcXxGax3/Gp
OlyNqAPP/TZG1Wy5wv0gy7kbOQgbGYsHrfx0uO5/RQWsT0Xjp7MiFTOpUWOmaI20A13S7xhl0y6U
p5mLjvMXGyIzlAoHzBjpBE4X/tSba1106exoDqilKHz7UQc9MV71imyonowJj2v8EgQ5aj/kdqlK
JpAh8U47JmNDgj0Y56WXfBVud26o3+y+CRXw03iYUtePupmLoXx/JVIUvM0qIOalU0Fe49aSFN4r
u/Ix0cGytE6xV1/hO1YZxgScZnqdPo9iR/kNP0VF8nHw+hlERXS5QDBeYRFoD1mQUlTx4AxsqHhD
wDF3yzXBsqi4QtHbZQlVV8xbtyB0haQ5fJsEUDkU0OubGsCl/8UsdyIFJ6ta2EyRhuWrzMonGcrq
pUvnZ7qy41f1Wbq9grnaMPsNcyAtDuUIPxr9Iox26ojXCN4EWCa/lPKNmgpXLCYPrltEN5tKol+w
Y6oWCTuplV4FBp1xXtm/AlE44X5YBv+hKKl2gOqX/4DGWiAFimTb/pcMRY9jgl4vz1fOwmzphNNR
GwX6gwnuY3ecaqC6mGiD9lXPjBmX5lGY5TfU9d3k94psGFKgmwpSg8ZwfkkaO3mba9bR5RBg41V9
5PG97UwqLTZARGK7WVNl7njHotGjeDszdsqy+Jf6n0q2z1GYXKP7Zw7+TZLj/1BlgbgSuc/W0qq6
p50oTsJqTD8FzoJ8YnnxanEfSu/lfJyKPO+RtNi5h31rEwmuNYsypx9fxbWQL6WmWkhF08HBswVl
BtJxtN7C9oj1UcPbzkqQgif8a2dbXytRAovHgXV5DeIClW+oNXokBR92YqMkVaRzErWU/6eONOoK
htt/yBiFUQR7mLuPE0sDKRhJ5N+Q/j6w+SnQhowX6dSHobV/egN4hwpalozcqoI8dym7NuPY0iuX
TExOjpFPCZSnnq7g27qTmge0xXd7CdSuB+bRhFrNaVNiBgXavD8Zss2n4YNPt+slnT+cfTyKpmXs
wElSR/da+FYXmt61SaQaDGTJtKAMal2Y2ks2rOMOq+03xrJN6b5CSJd0zruq9qN9Y1XxTT0FalUD
EP91Is/sURiekhHN1stIWE/g0W/zR/Ha7Gk4psyTBOuIXJ8JWoJXpuUog6ExFsmVWlfxQnwrLJfS
TO9Sbc3khXxWZmhPovC6OrquJ8lXfmTzAVSxQtGv0ubaBcn4ouZ5kWe3atKgP2N2eb3pV0/Ss0zx
t5KJMMZaP12PuskzUyicAo5gvZPH5FauOcFrgMixdmOzenMzc8/feitq5jrDpLS9HDHyqkQnA9GL
xR9VDbufqg3sf/Cr0VdRtU3YtHJa2mdTTAnMnF2m6mw+ewYDJPsuojpdnCeoc7woteu5+zlOYihM
CkaI0yEwx5YyTwX0VDOuP8TtlgIZ8yYglMoZkFDUW1aLXuj9x33KARNSWn+YCbg8knTXHe83Xqzi
2tyKwS4l/3BgV0PtnVflj5hYTFDxlpEYomlASiom1g0xdckzVyWn/y4G0U+m/fbTo36IYAnaNLUP
7rhzDcIhi7DAybu3s/U25DpK4jEHX5zWhMh0NOrGKSMNCp1x+QO3uNDi/Dw+P4ysBxArBST4ai26
DTmW3zVvzLvmH+qUcVPU/A8ZA8lO9kNt1woFg1vXQnnAljEdWYVeokRUmaDqrktdWqaFpW5h11Tr
xDWABdhLTHBhkCJb2YrLP0pOuJOnuF7tbWMipwGCc3RTu4v7wY6uHd4WLX0xy5sdPvVeZ8E89eak
a91dC5gYmDuxq48A2rpNEDaqeQkoMsKhMRWQQ4B9fAd7vz0JIHCeU/SQ+81EvKOyM5/N4Dh0lV4E
jE0yt+ZvP6X3rHq7j9ZsTOIVQx5yfSSap8R1yVDHKFgw54RU9p9MZvmnlUgDs0hTqhMr9ybg32EL
Hl8q1/53w+AqPXixxSAHGSESdxUrOTlvRJsQlob2+k7H9itGM35togrUOEl4S7rrpnMczTJWMCDJ
Voh6SmhzBh0999qQuFSirhOklsFkXVQaA+QBaGvYa4cvGpkjyqdtbCmZnVhpvr8VGOVqfYpvOzGg
UJFkc/mEkK0vE1WUYKElUwyj3PYbjq0n7fBOqk51eCCjJ8hZimoNA0D3X9pYaLG37qzuUWTZO6zo
zuf7tdhljbjik0sasUew03/2g3Nz+EPg/4modHOfrgKsHemBfNPb71qv8oYKRMtptXSgQqskrjSA
O1t5S7bIruz/ZLctnj1CCKFsNkHFvxFknkxoCE48cn2j8JBEZDdw2SOp4I1G1M95ReEHE8iQzr3L
6s0PtEVLM1iOOVBHlnl4zFMuBaq6l4YejM/HXdRl1TQIVrY6scOYgRTWys0rRNCG+TpsX9w0mn5G
TrLS7qcVQlVDgmzc6OG/bsQmkpYEGCKpPyRY5+g/8NyJ98hDuuCH+xrLB7Y9mk6EOLfGkRyOWTLi
U/zT+WWGkhMsXrkg4y2PTFDGzz2Px5kyqjlSGXU23vb+vF5u9cVv+PBT2gARlxSbR6ryW5myAzsZ
xKyht6jgzW3IT6DwH8Rig78b3qQEg0Z3rctSMC7JvX+LGl4fYYiKgcUBffVUOyGx0Sk902cQU4Up
WjrJ4DMv20ggrn0CZR3b/3s0ZHitJa+htnFHHxIB5/PgFKS2eFMY3VUixHYfrY4V+IfOalKqlBW1
weaz/4Y8YkT9GEI/TISLToAw4eosrCMLW8OscZLIOK4TaLdfRGRqn4vUmMlQFTylFId9HiSnrIvp
IOwCJ3Usj9oagu/jK6m027fN4BEZC0u7GAbfVkkiMQep+FkcV1+byHXO1VAdLKEZcj0dBF7E6rlJ
EHrSKaZgG8F7uox7M32CT6uk9LNWNjT/7FVKlg8B06TQHCCGXT7+b6YD1YjeEywRPCMvrDgUKkl8
yTP9Ob6IQVe71gQDrFYAs/F/OmIhACWG0BisWOG7XjggZxtZTM2RtYbDNtcMIOxOVXeet1z4X1pz
PBDg0h45sYEsfThfbsnAtiNG2bTuQsVecxednrAHT7ojFNsYlKyHUjGyoqsQFIzbfpFBqj/m29sf
QSsga3g38gi1wQAhFBG4vRXYLhoCpCVTItB+tTjewx43Gmspd5MJMeTChNg5ubCyCvCqlyptXaFT
E0YFz9BjhLgZuj1f9tJrFHM0Uk0kVHvvtdlH+jMM8txHeO65q2CzkFR2GkYJ0fFPSV+FvBeC0JmW
X/qyxE3ESfwFQGCkRoqxugZFkrX7qXra2h0+gaSMoSix/kN7Est5JvBD0wJ3nZ04i6AvyeQTVau7
lXExvyfa4ytopJAyGykyy47eZpHCeB7bycYbxop7MtFF5R93E87oHq7dLaOHIDMPTzPUmMadGW2t
hLgIyNfgsgF6ZRIuMXYWfz4nUGA+hoPZDMOW5L4EIEYf8kCVykm92oFYfh5lqpefF0U5zpOPSx/2
pfPdO8Nktk3m54z1QaqhcENVGZYLLnHWz/FGoxx3mNpuO+J8l3nEkHMbWR2EusbMgK1mVtdhjt4+
zFljQL2iasBUXenSkJcW3VoDoJWqHXusY2nslZvaWx2/8aiwmtltkQj2ATrxDts/ebCEhgBRLCdb
rejVJ21Etwk3ZreOOX2RrPVpX0WetcizAWJgIwcWEajBCAh9+Dkau57Qyz54lcYFOWU8AKEYOfu3
QhkSs5SmM2nPbHprf2vcqlgpupxQb3Udg9fFj7BAuLlX6nvucxzbMe9+/pXYtQa6u0prilf+noot
J8QECDhVKhfjXfEDQ2JQMXSvHMCoHD3tdtQpSMWxquJ0hEfzTn0hm3q96QSr003ZBVSjPDT1FQSs
Mmw9RHmQSZSA1dhzRZhrgmD8UrSWPSASqa5133Iyof+sdFVzzoo3ImEms1hIA3ABCau6TLReoKsp
LLCZR9N3Ys4BQ8FcQT8uHvgQLxARUcn3bwSsaCDyiaOIEz3+RYt1NNr5qiLmd8qIvuzDuO8+4Z2D
X6InDzEJg8A+2W/1IUSxHRilttBmsXNYvzkNRNK02Ff0ie0ZMoy5r2CvTFafnl6suZC8lQSTVe50
VdIgqZLdUAW3gZARcnYUS28avt/rRDqzMhx0wOkHTX1Id0teMsqct0WWRh7FsyF5KpnTnHE8mhnX
JIzaMIeN+vLYUyhi8cSURvgpv+N5rggVpxrxlDKe+pkQyjMra/waNbcKZtL6GSh3JGzuApM5VzPW
VT7qfAIenm4m4G4D7VnqDjridhyS9BBym3H14lLK0WHwa1YacIhXuW9Cmdtky2yeR8wRtdrHCqzg
bavSaeWgLaxISQU3gTxB+VxBdYqhuv8m6cpvUUdHzbuaIYGUJjN4o/pNXxV+M2C8ZZWC0yztQg6G
x35LFw+P8sTesm6fbqBYnOdvUjAuHc7HXcy7vW7H/fxmVdVBSpIRqmiUcauv6OC0kmhGiAS/jmj+
HdjRl96cjvVd+WmMHuo/CginE7b7jdAe7BZQSSpuxqvT99gE/QVaNeJ78jD1YBBK5a5K8++cTEzz
hbLeSNzk2rXKxFmitHVSAMFNanuDAmzEhwRANrzYb3aNng15hewgO1EjzjInWE07BI9KE6YICBXs
TUUdi2lCYrxiz69jLbuxAdFovyu1FSroUx1JlQH1zYA+TYnzZgkP6Q7uL+gbu/EVAXa/03EwIWtL
Mzpu7FSrb2B46duIWTpfMgGLt7Lez+Mzj5XdZrg35DSs6B1SjClqNnau7FXJSDCP2joFWIaLC0ZB
KT08mQBwhRReKYma73Z7UF6m9FMDLFNFX3C960BTZPPxLcaBsxCY92SzPk2T6p03QEtUoyHdQ85h
SSBfD4ZZmJ2/rZNuOUIfaJLXRBWoYUZXl6aCjAKvQGw+aiBM1Rqg+Q9f6Ids3FiPbuYo0QgBoEoA
wufBLU2leezsVHK7JCklaMw6tuJ5yPKIzqA5MKdEhTM+Kxvc9FfbL+L2817tkxJsjBueNqtnr+Ss
RHYGe9LA9jzGMh4LtR66TUsFxDtFWLENeSnY7Ex8zMhib9BIrkLkQRKD4Y5UX7135y5hGrPF1gK1
eWcuGblx0i9z0PMAR8msxxcYhvHAC5q8Fdtb6BCtmeqEylQuymxCT1OF30p1q04bQ9cokCKttLRp
9Ag0sSHX440NvaBfBwSXjE3J8fsRirjrMklExZljjYA5hQQ6ETG30LAPfOLTjNTZgtm6SQ5H35ZZ
8me+V6nCsO5s4nwSQUnjxfiqwH/X9OX3ftE+DplVdYhZkoh1djARzRmvolkGp7WLDTpdZhjtLhWv
rWSGZEyDhzrfeh2tVJDx9DqFxeL/6Q7NDo1L/FmPdJf/fEm4rnHWwmY3/1hDedXhT2fc64fot4xj
+w0Gl269iye+3KWfX/G8d+R5ihuAwE+SQ86mflvlK+XP11vWmrK2pi1piT/Jy7LMc7NBxjpJA5qd
G4RKRyw13ljRjTVXB26D4NAEVbeurCfpLcpXgS5JjaTr33h+CToADUpQnN+Zy0ZVZxOYblSPyKhm
sUAHIWFsJPGkE9Ez121CZ5UgqHGx0gcSDO8enlJAl4JkoidTAe1ixu4YarjFex5yWWqN8iQRSA/a
k1SOEnV3hNt5z0cPSm8HFZhEsWbTB/GTc0jfkBYhAUzv8nocQ4mOfjcXixWufJ835fXiqDpUN6ig
xfXTOHtJ+oG7/5B40YVzav20oICoZxchgku9F4uMj8JNBgCY/0mEs1q/bjwxir3wwz9bU+KToOcj
uvlqD70jgUrbPcTA8E/yvx6jZcxnVw2sNb4JRbQJpJJsR80qgJVjEN1Lcxfd04QCAk79reytQ0j4
W7kBzGy9gP/1wNVcK6qbL0/xMd5TmfTFmDDxIfT+ElJeFi+EhsFzdvRYRSfrHEK+SwOTmncTseIb
FlSweswzPS0FFTwxIVnmt/FfiI6OmHEVbsL9fJB2Q9x3yU5Wz/Wtfy6K9DvVbSPq2eJVADL/1AtS
PFeTlZW9DKOS57MlKKzjTe8ZfycbYm5TelKlIFkFJkAxPfmOY3gRI8Fk4dyWE1KeHT4zGxnWtbti
vkXcIdR9Ns/fqUBVZtlFji867T5kdbVsIA2SUkmWHyT364S1q/LIMeVQVH2L+OR4qjIrix3ZTES5
npk6gie13W97ZlwcM+sNrfbdD1Nzx7uH8rGxtAcbcl4Y5+9N9sr/+g/ZhfjrToVQtpZNzZMZGpJm
Cs6OtMCHDsdM0PYcLR8V8QrwNNoyrj126Z6nKJN2jGtn+B3OpJObz/kjHqCC21xp8lGob0jnpTHf
hirFETEcpGuSB4TJkLp4vvpq9ftaxKX2t54Muj3qZm+EoMQmtfik9sJKo2DDooP42hCC8qBINnv0
Ll7gjWJcKCls+mXdeLLVHpWPD8LgH5c+nMiHSQ7C4tamEbuNriTVFegI2MKK458XbfxzhJmnyW+W
4spYgsjXaHaf6/B2KarR5UGKZJ92Qp22uoHDn/U8e0s5fUG6Wd0xYhLQ08I/aRItSS2fgX5DH5Py
BnO3fz0iy9s78GWsJ1jzo+pQnzQpm6jYJVduSeSAnmplKD8/4Gwr8PmnYEK7y9O5WJ0BS7orpizg
XTJovDBPL4Fvp46Yzsc2UXsRYv1S7jqgKIO5P0ngCdhKdfwpirkO1aln+yBfVpNO1ODZnqjzo1h0
VX54xEZsXFtu8KrEi1DB4AdRaYXAXiYVpAwSfvClPtgaHJmKsDwnxj0Li1wIBz1DkcAceGe93s7m
2Ejjs5L/gcQdR27d/QwrPAYfQcpvzyruFKrGchqE4VX3bS2oaCpFt3+bX2MDKOBLDRESt/YBRpxe
F8YDmHt1cXaDL5QluBniFkim5abxh8e6eZ4d9pX2glXIZPTYS+chJFcyFFkHhXA/0QNh0kAtNNdN
NjNlQ8/n8f8iMDA+kdjVYEvP4a3zJVRDZ5yjctVsmvUORoukumoV9FtFaEPX0ssyjqp3xYko54Hk
/tkb2zsWVTTvtFJoj42Hu8bIUNg5QS9QxejZpR3FPlNhJ9xzfNe5K/8ESchaAQbdHGLiQ5N27CH0
W4ChckeGMtpnj2kpy7woJcdxzVhs2ZhdbwOZvM9sjSvHGaSN+4JkF3ZN0HfYZupMPn25XnVP/ekH
XwjDG5miDZAau01ePk580vOR70sujS2cmyP0e4PhVgdTfUrCJFPPYfsp3GluOsQICZ3yfu1LCnDQ
fpgL+6C8UkVPxFRFoYuu6sBb7pjswlT8OQoHNTvbGVE4nJLxvFEKe0XPon7PU8c+cK2yku0xtJvI
RRhg21cGk6hiQa0OeRgQ9IMe+9+et6l6QmZXUPefpHZhBNdvLxsIfXlJB0OOcZGs01Yux74Ww69H
NvozTW+1j8CftMKitKv8vXONk1PlYYC+3PjboM8kiadcwLGwsGmoJGFuRZACWFqbUiGu381by6BM
+cpLAemqDPTssyRaV9a5Zt2kyAkdnJDJfyIwrsczAtmkRuhhK3Qv/oWWcTxrOqFwzzrdKXGys2v4
qv7ZDF9QVzE/9DrZ7G3cE9y13PbArvbjlgIwKOd2Tw8Qabge1nkpPZxkVumQ/VVGa4wp18B8CddC
Gc+V4VBONzK6dFr7kFekBuVuPYzQcgAzMt99V8S8kSEa2elpHoDF2WAuBDjWi3I+V9t1gqV/UGrL
LFtfnhaCUh9XH1p1C2c0y+Isr1QMuq9Gn+WIO8VRQLY858rdXb6z2sw3zVw8TEovrE8/aurp+pjQ
5lJ27+DjNQhpV1Rdg4fuIUQz0H83VeICWUpoh5jFiTjG3COJhdxsbgeM/mu9K1t4TX/Pb/JLsBSe
g+h/8caL8n92mUylG8yAb7KtPoyk76E/KmZvJTBYUA3r5ZQPZZA6DbH7Agqs+IBaj+PIz+/eH69c
XJ50ssggAQMFIhm8oH/T07v/cCh1IKxyo4b1iMknhU27lyu+gYdThtMsXSaG7z8cEBkdA+RzMOWz
50mSvORZQaMWnD5W30JHHZkx1RAhHAELijejNjD/6OTjxGKmbEkaduHil0+zu2JpskdtXrPWJWwT
90SyLQTiuAWnpSXWDJOn3N9wHlBqqEun4ptByNRskeWBJ/grNeX3RxqPpLu6xK05r10LoiQuG8Gs
Qg4tlTHYf9Riw02vcebNctODfzfCS+3ogqXd6jLgxEackBm+NMaA3C0uWrbb+MfWjGjGoh59rt21
lP5lDW5GH5RmesfRZYWzIqvJs7dO1tjorwIfMx128F1NLdk1pFdoPPoJetmbmXoUDQnGiwrJvG2T
vw6J99jatLVs7oEvurjZfYWLcMLd4Ouc+uy0SjxhWmuCkoNm3B1LcEQaZ1CvDX9CTy9sdkMK2J1S
lSjokJrrYXO4zZWiM/bP+n7+E6d3GkYyaMIqKSD3W1CYzv3cGokc6zkCGZPbxk2k2vRPmCEAY7Y3
ELs6e6Kmjv7jPLwAe7+UWRCjVGttXuzlETnvHJSUFBE3IppMckP+jmf2S9PRfZQXOaRf6cfXHu51
eIDGiXV47sOLkqzwBM8QntwDZTWgLdoMD95sNp78FCWBOBtzhi4es41B/mCCbMtdpZuQuhcGBXHw
S7UQobxSGJqk7j7eOFNiF7UNh3ZxiQxutetqdgXN15MmNrJT1JoBdv3ds4QbA4GrJSqI/Omu/aSH
RH/tfwnBQQ8emT5F1CIQKdw1mDWJ3gR9jtTSOF675P1N4ch8zN94xrmA+htM15rCDtNImhlzaZUD
GnPibASnVjzl2jl4t2FUcEDJiVV8HlD7uchwTq7DU4ZNUqosHohxd88qLgnxLBOLfc3aTnTUVeQP
Zr6UfrVVvhv1gZCR7trqsvNaHK5e4C8GB9mtJ0rbWxpg9hNjUWtv6CCHvJunNU2TkNPdacphZ+e8
0VnEHuIpA9EZM9q+1vH5xZib2J6GihR+PTr94nZkf/JoZXFaU9VZ6EmhJMTT9H0CFXkDik0q04de
TkA6TopQViXVWN3MdIH+u134BxraO0hvc718oIslNtagZfhikegHrpI7xKFjCOs/Xgb0otzN7BSw
TNwDD5aHK98HsU+/I9J6uKygA0yznSpNtBOBypjlQ7zuL12FEyVlBEUhq/c8eplGDpRhpfn8s3dW
AnmtK9jK9ofeXR6v+GRkBwLvv4arNrJHLliVnFV9cALq5WnxHPmUEdYXRk9BWSjIHIhWEiU9HtXQ
QEn0v9A+fYJ9w34vyVQEygEooIJzhHtSeCqbpA8++egpX8FLDlrhlIAllt79ayTKEKbA7NrozN0a
+MWUGFU650R5eGs8wsmffFbkIdXfmmWkPV62TasbYxD/d/pNwubihKuvIigoQeMLoa08us0xhNZB
PDvckp1Cn4t4u6pcfzP0jG4wSeVRlIfg1ZzLKgHJF6Z7i418CUdTO8KT2fVHeSkDv9hWl5D4DZn0
we8JbdrgZo/j/HIDQcpWfr9nJ6HIBhkAxeJlgGqs+QxS3vz6poAf7sQRxAJcQw4F787DHP1sRrpc
Rgxh5fjZWQFNHYCxBiNMtOREPT9+kh388R+6dLFDybuOrUMTwf9SftsXOAOeCQ0a+QgENdJAGz7r
4lp3dSJg75QR5mYA/NGiVgTsMQ66gsIuz3AP+Cov4lqjjZlnXDsAaUiqVXHhGBrrAR4cmiqRDtBK
yMardYhl6wQQPhcEfHzZnoy6TLor0tcDy6TcSiE1XXYkWxYxodHSWSVX9wG5gHzIf5Ohw+iySgoM
HxEw3p2L6ZHn60xvfEP1tcLNi7G84+hCEFYqCuwWmtKwKnI5e4HDiMZcqWZi9/smE7FTTck/Cslm
ftPQZSycN90P2FMNtXSx2Maf1dn7RyaNV/rLrsnmudsYjR+25loz46rJRetSOQOg4G9WvfF3EDzv
PvRiBbRAyVxCt8xxZUlVGxhi6N25HFdJ6lPxBU4VMwhT+a5IR1vYtpjP6eCFj+aLo7Vgea9GagI8
c3Mx+kr5eVlv8aUZsrCGi53nbMJbhE6vA3LjAnrqEz/7cGZ3Tto06xttWh4LAoed0/QvTAvtDUjV
bcgybZHkOwMgPXgMno/nGS7sWMC8looeCKHVQaPgytM1Nt/rrtiBAG4Vdfth9FoIfn0F7fs3Voc2
GnuPajQ0Vm+xf5n2VRIyO5+JNPVzcPuPjR5ZTpIKhv06ycJ26jsUGi4Ju8PWXT7i4+Jhh1UjrjsX
loYaZzQqQEhfiQd0SAaPOckB8sDqgNaAc/fPXq8QWa8wl90x9KDwTOxGzmFLMePV27hULT4a7WSR
pY6gmWRV0XN43M9V+7kS9NxUx3ujq88BkLUkXDSM485HzCDBKoZet2g6NFiikaIufD6CkPDbvC2a
lKYk7a5jVi/STD1kpnsPLz3ogUcGlYodPnZbDZ9yb70uOsVmXAIuwsVb7Jtm/Tu6cfqTgszlMYQ4
D4xvJvAC6FIHSFgY5/sbbRGcuqnlnwGAar5CP9rfE4gTGNUMiu6puiG+U+vYEkpsqxaaU/qhmgWU
S3PHOpnF4qJ/XI8nvGcWS/hIsuFEokePMXJwP7XlcjtVECm7wfNMhuSUncn6l3oufEHYGhY+1Ooi
5yqkebji3gGQG03ke2CRxKDf05d9LCe/PqWmB/YPX6BH7Iw3iBaiHns3l3oHSgZdUFeSp+H6trg+
cvKGcTwTe+zrVSCfkQ2w85jc40A0WtcXuukqlBydgc6d3NekvzSMQAux6j4xYo1fuBwPu3kEdbKh
kd49MizZ3LdbLztYXGaZHQUSXG2ojyK5qyfQHQuEbJ+NkhHDF1sPGXY3eQoh804QGWWqhSPTfo8i
mfQETLbS/NPTku4F9jlqlx8R42laCv8nf6G8I7Myh96Tze4mQw6HQLcnRfoQHhj1zq6l0dbC3lDx
IBEPuDBXRSfzkownsW2b4RCQHG4k7ktV7OSiMAw6RCqOXIe/dfiozaknzsBcB1MzOi2G3PHj1Xj7
fkCDSA7iHStB0QVw6M3H8SNoedLdSDykvxQSSW1nZ4L15Begm8EwuzkQCdRsqt/EAmnFNyeWQ05u
DNHmpi5oXy67QdgroMpG6JPcQwNzbktOg7fyzkoDM2hcXQj4N7TaczdmXgcC/Lslme9bW9PDv3Js
ksalv8XUYAOslxNrIHIxnVvjN6iJrdEyI54QEYtbJfxjEBTYmSBmsbemPH4l1d+q48gc7g+6ixhO
iAJbnuVtjX3/QJpIpQm9ESiCa5Lx7wRiJN0Zi8mIAz9tZmjern44V6mtYolkeAMInhXlUgxpxtwL
fm0wsFjb/NmxOim+JOPy7+7wjYHqf4UQ3XKhsfTpl67Kcplm0Qu6Fj4sEFp1hlLj/j+AyhYcTiWK
g2R8Xggn5beNlR/OqZvIiN9kAEadT2w4BCLO+UvLnwhv+giGaQV/W+c8Bsg4o93Z/5CWWQqZ45rv
L7K4VenBAcXjXgYHvT/sf4Ri8HGuufH7GIP7z1aXXDJEo1pvBR7X2uinxOnwN8DDr7HsoPg/7v2k
jH/rfcpKEIcJnVhy+fnw+Zmk7o4ItyP6MyV2c6hPFgJa0RlHA6/J7oqAevBP22MWIQH0FgYuUABq
tWvfd5meuNCMntEO+6DZ0zoN/r7QUCWiz+SLvjrh2PHdqMjLzoFR8eAzkdPqR0w1vEkZHbKdWItm
TJ0oozTYqTdeMWHHVIb7f/m6e+K8+OSA91mxU5IJ/xJwH0jrHruw3R6XmL22xPmwgSmqNlkSVeCZ
0qczAfLV2B6q/tEyqVrPN1lH8s60ALAt+gJlEI3Kz9cMavwvDdA1xSZ5S+z1ZW8vqHlIrzY+SBXm
uADyzxMjgcIK2IzlWgBAlyTmn+oYpBQy2oOHz0gAWn78wRgWypOvRd92FfrqYO9mR2zqU/X5aUMs
4srGEk+013KPAuo1nM1ZOKUtB/XjRZdY825RqqWvFb6watcY0CEYJwFy13sEIHpkoEP/5WSPS06X
hOintrOcQdd9gC0iZvt4j7bnAmTDLnL4LdARMbsg4PwkRd/Qkx02pnlW8GHnLlp2AdxgmNWyBXUh
nP82Fij/Ls2TOxvJjIgC8PbRkCtQQxNu4cBpLZxWKf8XGxG/irVzOBAb6hJYRKUnBT5243klEMnD
r0v0P9hIEg28iZBlUF/Zzfy1PWm3FnWOX+z9l2jZczCAsNI0RdyRUybjfnXZxTxV0WbAMufRENxg
tZtK6tCaZPGgj1A0saD+Ej1p2tL4AWob1H7gW9iQY7AIABS9Bnd2VeB3EZhKALAo1MyAMyfTiG8J
yutVd53AtG+jL9L4Dq93wf1GPDXqsHNHSB77J7INKK+juNC1flgZROtLaY68hdG85z7rwJWFG8R6
d8RyZj2uhupE5jUHPmSVk9S8KwDMuqMYLKqL85dCqe66CNhlg2Ekssnv+Cl/px2K6qqpZnS8bhzZ
56xBqtWXbVvRSNppQpjHC01K5RNzZT/+xN88mxMT85sFFLMcJKTPGceHM+CvcT7cirhT5fO9J/zT
L7coYm8KFpuCU4zJ3Gk3bcQJFhpFAR6OujWeHQhEzYdwPCGwFmbuaXreAnSDsfPC4l2K6cFzTclw
e6DdtkQMIJEGipTRxiElbr0KpdYObhHdGkz20lY+cJib0NtLnW+rIv2Mta86xw51pAhkrN11tAHW
fTx08Z1DcNwJFfZ6PzUb2ULOVI6DkPWCNJQtRDQafPUYta09eM8rF3U7YTAS1RhfhjO8BsLdheSM
9mjlwZ6K+4+slMVp09FKmFtMZjLEn2Wz1nJpSZGwjoxbZvLBaKOpiK3B/WRzXvUBoqYtFzcK2o1B
Gqr5WqaYoNQyY1vVhCe29VjgXeBa00Nyf72seYqtj1LDVAt6ciEg5OWMuwEyj4jGy086kopRjte+
VR5QMuTR0kLzU8da41VZjGCmuXY8Utx9ZMMBM0uT1r6EtzfpqLnvrfIyR9c6hs40TyB/dPAm333W
ctBNjdBsjefK6tSOt5gYabFWfQXO9OUef40ZDrOsr0T+2RSlF1gtO29E/UHpH+/hxMMzgIW5V+Z6
L7k69DrcCs9lB/kxuKeFu611JJinZ/D5ZOKKRwOxze2k05XE4tk9gt8qQKzw6qL2KA3vklM0l6hY
1wgeXGjOq0+ZlZBZ0H+IXpEsCULywQw1IxiAWaZPsGQunL8cNU1zCsJ4zSzZ03SdAY/AwxLUujH/
PWUUuEsz1rnBCiHuBVT8N8RP+MliLXSZnxIlKWNIOM+9tyCghRb/GQJ7AZI11+CJwSShHiOvS1Gg
VF+lb95ugYe1VuZZuCq4yUOchIgtfWPer7Jx6OvWicGyAhofUTeXiVn/fFDH7iMhFdcR6cG2JkKt
rVREORFPiRwpLY6ArdqQ1Qb8jJXn7RRPUSmncVQplfG6nHJcB0kGkhzsGuwHPyqrq7CldFjVuIhc
Bh++NSrkRTrBw5p+KswEzcyt/s9aJIsihR6P9XSyPId+9CJ5fLOPN4m115/z4w7tfRVxTOd49BiY
5VLXCJn3X188+w4DcJRyBT3PM4GMcZsB/F3bKi0yJn6YGgtxbnIGaGZZSEib6o2yDHS046vuVzz6
atp2lIGTKIerXkURHSs4xI8ADbdU49mf8qVZJeZFl27BQTubuigDG2LamHm26DGLWoAJMakdA9h/
t/ZbZI+c5BG3yG94MLFP3xVmiLnI0Dw2TsFLqcwgjIyod4KMmh3wRCyQItEJVMiaGuEnb4WqyBDG
98VbEK84L/jFFHq0xb17V+PahCwyBF2lBTds6IkGYGrC91C5HnuWjv7LgoNT4XcbH1QEHsiWA5Bs
bR29lb59LAedfQjR71ryJNyQurYVzCnr0DjvcoiAcfhtO0SVEqITgOm0uxPz0yYd4MbrjEA94wJb
qdvVHwyyA2JA1Dswoq1Vl/EM4xnmUvMsghiNP9AETwq5IS+vMxcQAHZVw5ZQWlK001F1auxaBBc6
4Vbl3wdhBSCJChpPkRxut4ImTVLI8Hp0TI//arJc2GGBgxOo0tf2rNtmUQR46P0aBX4Pf26r0aA9
jzKnAQh9RZlIpXPJINYvoR7XYF8v6H7Pb9EQZm3SxRroGPuHYOy8RX9Y5QN7PxOFj+APs+3gZAej
cxBUU73all30EvbzVoCui/Rcru4l3Z1wNBq41XwN5attji/1jC9r1TUCjn8JEsSjlfOEBI0cHZa0
nZZt1Cpvt5YVK9pz/7rY1ZpfqTF1NY//HQcRehBA9OrKJ8fQwQrzoqXtKJRELDShsVz3JrcB0gJo
prhrP0J0f4OT4BPfh0xKCkMjKfO5QCHG/3XnvDdj3ZWscymsqbOIPsVAWIskI4KQGMdBJXUFMBbg
8bXBWvJHiCn8D0OkW2MH6Ygz0yAIshxsIBVyfIIazRUUsqyhHG0UAao3Ah0vnzL3wwnE8aotkVMK
5BhGHZz1KCM2Hb4Ob3mieIfMq+ve/U2ty+LviX44T0T1SPN7dO0Bs3dc+Ro6MJMfGrKxEcDYq8ob
iYoq1XnklHzcSsghxf7H6r7GkV2bpphhicQK/BOZu12nBxcT++c+vHvNQCgcghYEN43TrrtavnrX
qfYXNTssRZrTddOQAvDb8ry527nHFZsA2gZvcSEwcPaI5fdnhOXAoKbjlrTnEJGxPbUhzPuAYwB6
oYfpge1b0069m15A60mqdMyI3ou+Vbm6YDrYPim23VGnRusDSFcpe6dbq8z4RimqoIpVwBKi+e+E
zYYB8+7SX81NW4lEb43TFoxwW4+MG6V8UR02PP8QlVntD6SIH5boRP9N6pjY4q5j1DTg5O0en61c
rHWfmUoApywgZYcq8zEvmmUgrL4h8oqzz+paPo0RcPhEjmC2GQhis5numSWpctPEdmgdUxd0++1M
zS+Tr72wFYCvkyW9KimTI6fcYh4eJPZClyO3UM5MuHEe18kz1vC4NVFuREiK3KJyYvDlyS2BQDAa
RdU0t4IVRkByAJgiPHrczRE+1KzNua7qk2lNohax29Fw/kZlOaz44zgUmejo8kbaB0QDW1j/gtEn
BckEwMIZ3U4o+eWJiZeKYsvwookJ7eSsi6w6BwQR+R/uQ0QuiRY4jouV/BMML52ClTXmh9/4MMXS
VoPLUeTw5eywUL3qZrLtjzZ+dUyCIh3S80ak5Un3CiCC51yaxSBbqDB7bFkHiwDxJtmmQ3rckxlo
KEn5e9SMg7oY2CX+kisnYvyn9v566KMIxydAk7Fef3QI7wRggoGUSGL/v7/jLu5vIyYrzYJ5Z9N/
3OyaB2IYe0rjPX00eX+hNnzldftif5XjfPB5rBnFc1xziAbltSzm/yAxZ4Rp45KyorQ3BWfPm1mo
a2pITPNCoY2STuxRklyWMCYl813HLXTtjjivJS1ATAupp+bSbMdMO1Nk4A4cPB7kRENS6M2YBKKh
jtt0BVeu3Andu4WKwoOtI3bYYa1ZAhXxVtBhp4ibpDuJT3AGFP/kWp+ryDSwc5eeBoAwti6ldoTN
Ykz1epvKTr36lutN92WdEkViHcfcNl0pkTE5g/WHUcn0e2djC9oHHOdpB600ZbZ6rhUpy0d9y0dP
/pmQ7e9LzoWVyP4qkh/LQYDlclyG/+6Lh5f4oLZ6CUdsBdGjIWTfBDjFGqcQTWvuaY0MToPA1JTV
pAdA2akwkOitDgjfKfs0sTjo+5iEYrDpE4semkUHr5UuXkVPrKuf9hJ4rwnV3iSlik5itWSVY5+p
4xcknnL2lkQNs8RIRebXZZ3TOZyQFSwxVsRt6L2CZ/QmxwYGNdFVcWYa6TuFR+y0WXTP+49ICUcE
LZ9sJQgaFJv4W/zjyWtH4xE5Mr+qw7kLQoi5qDXLHDGcbOyJp717xCbg4MiB0+FIO8bXCwZ30CwJ
L71FwxQf/gnwRNYs0JmI1EkOOtDKs1RbbbYnNPqhlQSYLveCKE9sOcmIEUamFkoD+nQUY6iELFM/
sF/I4M2t7p0RiAFlrtykuZAKZ1IShlZjOpTeZIG27Sf2wCS/zd9HUf5tp/M3PzVgXVe5VW5tN4X4
3rFoBUPNXBk/XPhS2GzuQLihjlYkgApgWeip/lcTueF5KMD+fhItulZmgN73psiteQjO4skQqB1H
XAffS7t1iGURUl5Zofft+mIFxG2jzQ4G7LwCj7aIdHv9oZ2QTuyZOPLcpFekp6V5CjICaWUqFl+j
mBp1N7fzaFbj2iasoy3x5rwmqOjgVkyjOIVhInX/EukI717AmpjyEQUuDFr21v84HuvcyXttOMYy
+QnVA+6yd8KvTfaJUtjJLLU36yaVZI4fDcrMH8Vd7sCcxJMWwBHFktZUWSsguL1bgxeXcHHM9QDZ
xP5yhrDIuAKASznVZC+zsEiVnuUhrgf1H4Xdve8gSLikz9lsg+slMvNgZuado1AHDXP0U8VqKOn1
oarvyURAlcitXAfCdezYKz2l/5CTGy1LX3DTZl7UEusByqfHQJ425qxm4u0/hkuJcOiAz0rNg2fL
td+J5lF29nYnf0o40e+YYPyvxXALlqXN8+9ug7t5e7nGxF4lc4DJIMuss1UITTTmnPe4UX0oiair
FSBYZQcqljpvrxmZhUrBEDitS/6LPIJrUniytsESSVm9+tzgtuscL90V7FkvcX3ku8fP11hTvtgj
QKTzkgd5hqJURqIWLBL+FXLDaaZFmYRzyPz8rxQ7rgKZqW3Su1wRxGrQ9vwT4wMPzrSV8JT2kniZ
alyxFgQchXsVHZZyynY2FmP70E/sX+xU7OScIS+q4EnHiwdikKJZrEPs0eog4Ch5jOuDJ52NHoZs
inPR5idUmJvgdkd0FwE5IwNX4Pm6xpenlvClubgkDtfDGfvz3Q6h07REfTI2krAa5ZDDC1J5dUb7
1Oww2VYu4U8RwkOfx3zCiqP3JSO5JVOCSrXU6NFP5oZy0pHUT1d93ArbulS63miiYakmCDNfy0oB
TmGjp3+o2gU9DyhSGxW5cYV4vdwk8raNr3qvv0s6sWrKalBbfqyXMwlvHWf4vSC10bfJ08p50wal
eEZZG1kINs7LuzhBhUKN/WzxteyfLjs3yjpb+mH6R7AB9jmNZPd9SDZeQxBy5uMRkgORQYkBEiu3
DWPVSPfmOvJSTMwb6SYn6xalBdD4miJtHMu57hyms/EIO8jqhk3OzH1x/RGSomBNg48lWB3CjwTg
OOFdbngVRQ3FdmvEaE3iC2VNx31wwFgI8nqrOzYaPXoA9zygnb0aoJgr8lYixpQHybayy86eyjgc
ycBRE7ybfIvRRzijzNrjXPjcHGaVts8CjkOhx3rR/xgf1PRq9Eywxc2Q33+Keu5v7uqVOE7m1IYx
/KzXWkUqO634a/Y3aj89AVrqGQVCYg3hxoumSxSWqLh7tr1Q8zLPZ7M0IYUymNew0Zav5SnH/70L
uz6V0w4kFCmihxtcBDOaA72T54BWLRv5bjjEn10PwFsaXYaR3QoN8dkuHrmgJKbDzmmXiiK8xHhr
SqlFZuXelhizGvZJ+KJpLskwczqPLam/d0V+vcpc6Mbfj/Bh5sdYCKe33JM2mcxCk4RO9HeWGJSN
+YIoyzxHD5EwUggQJy83G5aSQKLUQ6ANaPNHMDB/EAHTqbAPy09inMaZsVMpxCDd9lqbYHuInU9Z
oZiJXJvG7XGDXzTTMIZuxlb+hYrY15E+MMuFSuXJS4E3p7qfd5QXCFHwD0aHKtjxIFaL22H1jBqi
x0UzpSnQNh6hvHaixcgCfDMQoUG6ZJ80olcBbG2BTPMITDqNMH8Fh0SyaycFIqiujY0bgsEPnk3b
T7G//tSiLJok2tEgrQQK8HzYk2D0c6WeTZjXHxnfFFjGmT5hj93njK9x/KGGFvDROiit1F4v5cD9
eNIpU/Su9Alp3qf2BFIeXCiEJrj2l+jPQBUTcNczRdFOcCj9TPc7enOLiaO48ZuD04gwrXiRfFmS
02vogKwOj0EBH+MMzzknov9XIXyTkTajj0CzHPN9L7RcF7w8NuGzCJ3DY+KVIQEg17XNta95TdYw
qDTZCxwfQjYE+njJ7HS23lN5KAG9eE/p93BKmKAM/c5Y1ToZlHIJkQpeytXladNfuWBS+32kYqBG
FAuCZ7X4GOvE9GdL7nhpHkLiLmMq8R97jO90kbDLfywgWO8DvXZjYiGBkMrv/dlS2vjcblBykj48
S4FS+S58Ebjmf3ieThjlvlas3f9C3IAB/o/qGs3SWFdQEon4YTA7clb8MeYCcuwgzUWfQdDG2RW1
xp6cDOvgpfmC5qtgYWpAoaEqceQhzsEMBX6xn5oMnMdEzYHQVJdWeaKnfWIZGrPVFUedHNQ623BS
wWDn/ld5lugYlLiuSMao+Q6k30bHVqaXTJroKUTy8+Wn1zxALB3BBm//SJYkBm2eSTVR8RGc07Ed
BhC3VxGGIk5UxixBQO4idRR1pN7jj8JvrqPJrqaivxNPmm5cimiVAoqUPTTGVRgAhwVnwaqhj1ge
76+fBveYH5VNI3DCGaJObIlO+Ayv3qMen79gZrV8v0iMV1+8xZUt2+v/kqTvDd80K70DCqH0gKN6
Syoj5CRuO8877Ati2PS1aF7NlNjp/SGtQAVWxBOCG6mqtHepIfZt8Lm5XCUtCuWLELY6HKKKmYJ+
/Ia70KcJK2jgzJaJ3gJ2Gy7/t0O32bfTqYQo9BpgdqWDB+bHup5oKdgGDfW7Oax8WOfQvaPD1g50
JceiXJz0SfzdQlZnDtC+5cTzAEkPzGnYatQySw329dmGNQdS28g/I9BZnlsZy7XbDEP5eMtiAoXU
xQtv0r/RIYY8tHCNMuQC0oTlFfrtyNFSqL292m2wDi/u5qdDlmjfo57RhNIwyLLvKchXB7moko5H
2qKlxgSoc3SWj7vdABcFq8c1jGu5MV3mxNU/4cGq83p6JxexmHLdiLY1WujQ3zXiUH04WhCEobKa
O9DqwyLWPt6x1FfCwSTp5ummoH5v5xufeDU3z0b+Ifhg+xbiBv9C8edkkLWn1TgXTSndblg7iUfN
iUOVFPmGTRBh6rzIIk4QjRsVq8yVnrlbwBLhlQHueYQxA+XLEoR8nnwsOCoZZD0/lN62HShnkP8x
mRIuWzdPlUJ0DHIFUoQgqZ+XjrXnp4oHrg9YJFUgDH5jVCvXH8xFNIHTjBtlM53RyQivmgYE658n
LCkVsT9CkX5lNf2ZUi5Zjsz/9L/QlMQPZ2Qsg06TjbfSGZuDU5YqTm99tPhbILv7+LqWwWl/+zh8
VIRWNF4znd7JOpA4BJRMkOQ/ITejQqrfH7bHx7PNfGgO105T4swH6Giiv0UhAkR4I5B5zd0d4R6Y
AM1k847i+/ZEEfKy1JDibBgM7YkN6U81C80/VawjMoatwG2AK2C2UEXyE92eAG8J4RlwzjqyX5Lp
VhQ7WpN09eeeveZnivIgY2rQCOHeH+G7xhsxa6fkGSqago8+V2BCcz5FqenxWd+PYNsVDAOf7O+u
QX3PhbVdYsgP091ffwmdT5GT0zjoTjaHCZtS4tVO+dcir1wXRhS3pAztP7RcEXI1XjlNjocbhyXa
mpr+enXlGmj+gX5RYIWp2bOt7WxpgD+AStwrn687S6DGtwGKQm1y6WEk1OBSuFJWNdPAV1C+fZQx
pW9+nS89Cf0aoDVRR8IkIAWHtGnaQXoURVpB+NIeyF1UT9jIw5vsECwwNNf6NalH8sCRyhLq4kLO
S5d9jRtZfSMGGePhFIAKd8FSiiP59PkQnvVvIgTjnYklBTvmSIYQ9KlISvA6PbVGCG0Hi7OLpD7K
8s7h0twDzHe+x44z3q6477MeHPZIDhPi7f+ZQMOUNReIrsfgoDbNrbHDJ3S3JqxziHZxgX0rafvu
UGisR92uHXBNUHXXXs3tvE7NjJ6yUA53fFDpLMEPiCDammUR6qhcpGvi4qQMxj1X6ihP32kSO411
RF26yo5wM2pi5PhyW1f57h/d5M5gjlDsJpTHGMXeCCxbQAX/sk9wwBGAkkHopTauUCmwxBQ3kLrJ
GqnjChKG/xihvi/mBquzXc/iaYu71AqkNGtzVfYuep4ADc0skiTnvFBMG3P36ePqJKJGaT4nKcT3
2rRIMZmYVktPZI4SdturaTs77WfMVDZTDJfj2rOJZIaxlmfDsOZbiLxPE0PxyJW8GYeFGKw74n2E
SAnHyDsMOBAscY0Y6AGuY3dAqu/nebTWcumEIDeA78fdfFR0Yf2BTBhRMXQx0Y3KwrDvZkqt0HZp
HmXIvYShm8DSpMNWhBr/y6fIzmdFHW2eu2JwSGYxdG0V7VKqhoM0vhit683oF/sUpLYvadIjBHMH
2pinrttOBWXhG7JWfJM1E5fB8lAA8e5e+/OC6aL+nPlmhf4i30hgeneIa204NOXnBsKKjKNDFhN6
bSlU6LOTcyTvl6Xe6EGEOoBLV6JheWYtkTcKmTHhStENS0bKX3usw0hk5UxlQqqWp8+Kfvum368o
xArEp6W+wBSj94B1CkAwvbCNbQIh99UCLjMLiILBqUls7tqoH67XS1hXcUZIVCCALfDHumfr0r51
bt6BRnkkH69HjIBlesvj8O+p0gSEVV/onRY3K/IfdPvU3JKy683vN9JzT9cDKqDA22q5io1+TZ46
yc1h79a9kAO78SEHFaKsnEOHVxq0q7zHZL7FsO8f9F/HRgbAwh6vsbG7dBxkSAntVJvW68V6VpCp
rxUoW+9o//+5sva6xK218so5CwsLPsRzTN04Ax/rpgw/uETHVi0HXWY1L7Mb2wj9ZrgrN7auiswp
nALczYTUF2Pc/oShz6FIa6fcdfdJP6XoCxImwJBM7IB2t/j4rseQ8K/QkXUsLjZWaKJYvo9pjuqx
psWLfMMG2zax1EqU3QpmNTsarmgTz67G8q0S4/3rXHYksLhFCj97DHQRC2/kjBIjDjWwE5I0kmCr
EHp+TPaab2QZwo9zPRhi0J9AF4uE5OzZV07vhFzomxoqUqxZbEpxQGV3iaJtbv3HTjpW69EbESE3
oKYxNIdKRkh8+EqvDANGgXIo3w0yfxGOztTK/VlD7xEUZ9hqd6283xDRn/h1L5Mwc6iwEYsieiI1
sBQ8KFxR0QfkM+qSm3/RjPA8LtGAgTkCK8MAjflzGUWdn4MuaJeccc4cf5IBo2DpbWrIIp6gKtn5
ErG7eqStsSE4PRxUWlC4NFzLlemBpKZmW9OWKuzzQK75ZNxizeOZW6cmrm4keKSnidto7EasAneM
QvVT2kLtye4fGIg/gZZdY5bd4ZIGOR5xDdJQKFPWhCnHR+lTWlclL4LNAVquor3rpEgsezG0iDLP
DV87QkjWWV8ch1d8Ctz7Paq92n7QWtKAN3ftnEIHQvcERKMAD9Pz2NZPyiEcD+z3QI4+4uKBwE72
yCd6oV8Z5WsEaJdhotNVcMDoIweLWaz00pPguzp9Vi1Zn4wJbcJXD+LQOEV3A63OjVTK4Pk9WVwJ
oKNLjSr9jpCvmkTXxzWRMYR1Xsvpr5/CalKoEw4XM8NJ4iuVWZPldPgVNstQ2q2aDwTcZ8LKdAn4
isdrPmCraT8Aj6Md9yoVY6A7Not6mdLmvxUw97UP/F3dJioEpdcqSE78HPaOwvoSGD7pX2Wteqks
9aE7TTnlvoJEriZNc87pP5vR7AQDvUE1vTtUlipcP0a+FYKErefB/w4TXzLvfpEdYWjKDfep+03H
kap3l7XKy+T23JiPFRi4bmdN4x6bFKg3zznKeXJEMjnjq8R8Kq42cvqPOVTmyswrhx4oizQoiohp
VJO4SFpqaQ0ckOP5E60GlCXLXuCgdJUZz9KiPlgwvRIE2n2R7m9Ie1+RllHTKMXr/M/hbo6olqN2
GRFBYuMb4bgNaJ/BZAr+qWBX3oSJhEMOjFNKGhG7v/2hqzHLo0UEBANyRJCo/VCXlJBIPWsFuqry
osCt/R6zTleACRShmbwrQ4QtyBN+9/PWkTIKuDXm9Qr4Et36w3I4WIwg8lKZWc2G5PL1aJdAxItC
9tT1Zmsgf/CC+t34YVv7oVP+9rQEqgCKu8mrCncuBd+c9uK8wTpRdusRgRvvq8CYptY7RWzd+7vM
vt0QYQHjQKEfUpd1DEAgEPX6fJdC88TxomG9TRAikO0qiyKy8LyGQ9Hwjjo0VntapEl/+815YCyu
lCdyYWkyLm4KrNzwGjta/3QrxoCaW+5oOtHo17MSmWizJv9J5oGpz3B/hXTmW4rXgJyD4sTG90tU
jtOxg/OlBXX5/aeAkeL3Q1YMZVXYj4XpJhNGYv52In2Gxh3+cQ6y5buG9tSL4eyuVfMzd6kTS9f9
R+xqbyFi4XOEC7fF8y7c+ANxeuKXtRWAJNaJceVWOaObIHF5OeeLCSPT+wGkIGYRzTCM1dlNfnDK
3cdx3pXpxnVpJPZrZ5omb0SjWUFrARfMC9L4HjkfUP5+NqiVSYpekQYTWuicW0TligHXR3PDaTc6
93e9w4CHaAOsj41qRkzSm86yEX/rrBA5lBSrOaHXAGJJdDTpRugYWNX99mEb++YeLEfLVo5ucTvZ
ngAQw3y28itYeaBsBG9GVZOK5eEqyEG0zcIXrroAWDveNoOIW5Lc9sVu5WxHmpZSNpLjMFOviZ4U
7ap5pDsrhWrEgImfnOieNyif5Tx3W3onRn2EZjiIy4m09tKa8aoFDDwDb+GBo47yJBM5CoERKVLH
Vf4bfygqYPjzwWxmgfdjxB5eU6mWopSXAbWX9Mladi5quPlQ+rznHyTaS3KrwopjmYDNxRpYE0HY
wmSyPeb6czSuwL3cyd4yKNGpmE1ZaQnat3nDdIEgGVmtT79KsCp5wXugbuMOSCruinAe0WkZDtmN
V/poq2vcZoIVDAfuy9uooWNyQMBGD4SmXdKxgazYgXr83F3jvoZm+oMK3s5LoxAsomzW3vDvSVbz
t43H0TItBnMOkkACwKf8e9gaTXZ5N3zQ023TqMK5seE8iiezHpgG+G1JopbnpyR/kbzXIgY7FZQL
ZA2NNfpX1taNktw2t16DIzw4mUAqKTV2KaNhq3nUfOsGOyTwI+DoJLmI4dgD+0LRedw3nDJVfY5D
ClXBK6hpTedFeXvu0Nx3aOz8WHzVv7+cLUER43EoUyM5cN7+KDDLSwW+VU2TDyfsPn/F4UHqDYTK
YigepNokP2wR2o7r3M4uGfpI7HqOvytCT72AAPnDRKrWd1ygmqMgo4cI3C27MyqEODN5n4cS3YMN
j+Dd99t48/Fx78xeOr/gHHNykdzvBkUfvq3arpzf8fh/TSAmmrRLgZRHcUTRZ/5XrBfu9k/0zLu/
nCNmyOnn+q6dc6ftWmPKHXVndSPoHbTLpD2Y3Ar7KGeBXtMPh/Bisxzb/S1AUKt1vcX4XBRfO+mu
sf/Sm74gG775rpnBMQ211B2MmJAJxnI939AwSgcV5X3RtYCLLj42PeQFovM31sSO/Ib4Z3ZCbEac
iOQ1wzFIpyOW73VKG8ZfvmeY5oscX3zLhS+UbI4y/SY2w+3iyTI08W7McK52rGIKt74luTdyhktZ
usXHhsglgmOeZMexqy49my0deUx4jIha0gR3PWE22WZ53Zqr6CcusVpvfm1TMrG43hEFDffVGmbU
YxQskku12q58wxYLcGckqfXfGxF5PBIdSPYXuXDpIMf+t6Xfr3PmYnL5kRu9GxzPGPIfVcmug2kK
Jeoxdd8+xcfL/vONEGtdFfz9K6NY3RN1Eor9BSYRQhNG7m2ArxNoyx5EOq6SRnXwgO3PyV5paMFB
LFrGgP1t5G0fC1XF91wvmAOy4i0Vw9l+58F+ir3HOxTxmUn2m01ZEHhdpwPdSg0fBoZg8+Y5cJbB
AmgnjCikOhA+zAbwdgpOmXoZ5739KglyYyp4kNlrshs2T5Xq3Oy4v5hjul8y7wpXyIwn/QWGBTWO
dwP7ra4i4RHQu4fhgMfIJH8cCmQ8DANASc8AaiiXD8fdvLCI1HQ+P4R0IidtqGf0A/rS+GVgB20J
73O9EaNG/EV5h84FWy1d1TlAHYhBfZJzQAFg+Wa31npQGYarJQequ9q7hCpRkf8MVv5xsLf8LOnz
scPv+YTfFJKlmckHJmv03s+kd5p1bYIBQz5HA6O/Z+e6hHp7zvfZDkpPYFXGfdyZHQ+86O8O6Ghw
tZxp6qbX+lCuqCrEP4JVySY60y9+cGavZsBF1naa499wULbfmftVpXeiue4ezApM8tXTo3PMv77n
JsmxKV85s9BWHQarHNZ0QFZKZtCAL4bUzLOQsypFG4Tcdghgu8ac34wescJvvGT4RDmVrmel1L0j
1eCyrBR0T3GjnTEydLoJEO1lSSjTBc8rhHafLlfPJ1icR/FfsYnwPiRGQXAlwH7Xc0VnvBuHCMNW
2QrMjVz8BH+eaf1vAeI9RhBZn6suqMOTDfvE72DKtHV5VmVqxcMY5/FVOrhFDTdH2n+jdAPRZe69
D/XN3y7XWbH0goBUpd4Mq5VzjFTlxu2EB331ipMx/z9jVcy10l8sS24whYV7VpBMYyXoiTC8YRUI
hs0/+nEnL/geG1J1FARiHnWDCDkhoxvWuJOk8FWyKvCTb4UPxANF3+cRTcYoK2FUB+s4X7EW36iC
b7UhFL0bMc6NbRN+t8bYYuIegiBUYWkFvCs+RDjC+GyPz+aNovV1fFyCjzOFSa8F22BY2mr/fcDD
0wRekmYucCqoOeMFiidVaH26FgBtLe4M3Gnqsue2duATj5LLrpOMbmmjckofJmE7mcICpC73++Aj
vX2t/eeKTk/dAGYvnynFSueWiVhwlbJ3mJBb1nxIyoaRLU1iH2qP0h81GzED7kkzabXDwkEy6HvB
QoySSkD7VlU7o8A22zXExXA+9D2DW4rrmzNOMEmn3gAgiJHGGm85LESP83VDGH0MI5KsB5aItxv1
8bheRQ06aKhS1YWpVBlW9VhyuyHpFc+0kLtq8tPdI24NAIdgozqfbXaqeKVn/eu6wjplmOfQXvmp
ienCtbekEQifYv4C/0jlRA1R/L/tlldMfsIODI7h4tfBjulpGlV3/qVIPExv8KZtcZ6PHGce951D
SOevGfl/qioL+WcRp5ZsfNNTYwzp7EDUKm+s5W3xRlcER5d/poQYoW8iATuw12PMRTUwBiPmcB2w
oo7DoxkeP7b1E0ApYJOsIC1kb8rfvNHGz6amElKJPji4u9rnNetPf5QjqHKXjcfIWu/gHd8XgXMs
EKERLE1QH+7pLqADbT99ajEDUr/GYsDfdvXqiAKJoGlJb3HgW3qhYMewyDIevZv0jUaX099aTOvZ
TN2dFwYwJzZIkFGYTEPSThc7kHGp4Vn992cP/+eXzFXMFEZUz2InHtazF9Fd+1pULPcC7b3voSFg
PZI+95Y0vx2L5vMjeZPYYH476E7lTv+h1kKBzWDKHpDEfR6mPz/sDAsK3/L6ZmfLO9so6KEroUWR
mAIaxCWvPLr0RCFTGxxkmsKMEO49u3xuMg5wt+Nvt0pItZF8GVmzNp9uu1RDw6SPikil8BFLR++y
kewOhSpSgIL/1veM8m/zNiSSrjESyHzXaQJESh06tVx4pCFc6e3xWTqm2MCeEENSnL8nnDRdQV2u
UJprO/B2NEbFvTca4DUzhdPohWkDE5Pc4+P2FKpoI+H3sg2ynyhYwBs12jOkJn3BICX8+WRIKKHm
cnjG9vVBU3sTAbPfIPsU/RASkWcp0kof2m5asj0Vf5J2jabJXYsiIGt/fX19Yp8vSZrAa//4BUFO
DMLCWh143mfQ6EQQzb7v3k4apRK5t2lh6NVDbdoQ56yIFZ40YAmO1WGmkryAaCSzJYePrObS5ACL
kNl15igz+GzEWaygAfDf1+T5F3yhzGTEXiHnR9DJ0TKgItnJPsMR1mGuXzOnCRwPAEoaU7E5m2l4
LVnS+MjriNvqOBIepBkwPkkFHf7R4KC1b9f6xOF9wRjmRx8GTEpUMcVFgQTMB77QSu0abkjjh/lN
OhbegQ1echHPY2uB/ID4mavZED0PStTm7yylPqjB/EJpX1667ThV0yM5Vr6uJBP/f+AlbylqZhyP
8EkO9Rw3gycCEEhiINjJOzZzvEA3ugMQU8boSW4XbYC4AO5Z3KMgVU9RtDVZfoTJPr/8GiT9ZNdd
q2ZImg8EJoeI/8q8SCNa2PN7azOHQol7v93Wu8/r3cEdZoVaDMegG+LbUVdNEKCB0i2YJlRr6vvu
p/WlvijXotsKX/pUAdT5SvFxH8WAX61ZpT+Fp1njjPPrsK8D4IXvf58Aj6mbMLCjPPoiKB0E9dIV
W22Z/obCNkgbtBAUABT6tSVtdbG+BCJt2uaviif4j3y2sUtCZp56TTefvMg8bfPrQVPefV2I2Tti
PExqkIPE/ezRT19quM7xmXI8Iiy5Zk+/n4UfRjpYW6ZjDA6O6jq8B+R69WxKmMg5S4seYmv8U94a
7PgQpobm8kMi0Rk/eDZXU63r5EHa0uiZHHpadpwO4dFyUByKFgSqriRbBTTFgkvkChJRSsPNeR+j
/mzP8yxvY7/jEB8HeQK4blKrNYGpmNjXrrcaqnySvMhrkRjn99bNiLyvgMi1t0cVvpSNVQuUtUOU
dWRf8VvLaQIYJv6jUFm0a3Zuf6dSZekLNXU+ZS3qLUqxszjojLYTMLayocvIUqOEL2U1dZNWl5SC
U6kCtEXO82tVygkVXJ9zK+1dH2ZH/9fUMHnQR48ffCvW7d0+JAAs7VitjvbQsRkp8u/3BGSJU9UU
whOImHVBiuM3I+hCWpaPQezg6xd2U1tDGmJXFHTg6gbzzbgoN+H5hQiI2Y+JC9fETuFzjWT4X19o
IJLoKk1yZJAA38Y9v8loWePdf+zeEZ9xZHMaefSKly+5gt2zMydXM9Ez82Ndb+xVmL7xh2IogIIP
nzML/BgviUAvH2SDIweZErVp47e+TRrmlqtLHqvUvhdCNSVpLgFn5orB6382U+itfiqfQnZIUNu/
MBtqi2DLNu6rCOMeKzOdyHOriyAwC+paoFOMU/bpbgjDBaB1SXMKdTzMreQqGhTbvPCSk2OA+Tgz
gg8j2LMcB2rHOsev+RRLLR66UiFY/cymxRLCU7kCA/J8EiIYrYSbuavhyXrlVJrGwocR9x68dcy+
LOknQETzGErV7cVeCR1a5VOox+VOoYDW0rNsXoqMbsU7+aAme+MwZ6rTxKFWXMO3eGVOvWT4inoo
8mLEvsYEvsGjYKukwGxWEUjJD7eQ1YhKzUxqiXTPUqrr96WGgJZDQc6eh2Se3s4u2r9V316b9O2C
QaKAtsK4S0stuXnj79ZNXnZW/hK5PixwJ1ruSdjGK99rFyplITSaMPlqb/W9s0VE5MQfWbhlnHDZ
k8OESbPigjrgNAJSZ/BQFLdDvlLuZigzgnlL6gFQpQLhPBtE6TweNNKp/f6Mr3UUxkFwe+n5YTce
YlMwrYx7Vx7NGYuIgMVkqKrmC9lrT4anUiAlf+/VcqLJnrlwM8S22yJTuH2wcdpR8hQ4hMsdtsn/
0OUNyaxZdc8yshnCqKd2XMnd4PCxKmGLs0VqD2sqD/0DyD54toF3YwnueKlQpxnoM0QIw8YN2ecL
W0ScIg44tmlWe5Eg9R5MDsXRRNRdNVILerg5jLnOKPSP1zYu2ftIhLlaOKbli9NdowM0fTAGKrWW
1X+NmEbqxTmKNyv2K3Vva4ZrdegGX/YY5ARf7d/a4cksZ1DHya59Qg0VD6vQHhsr+EVJUciJmVJj
2RFeBIxzXW01FCrk0F/iUpI0eJoUiVbH1Gqdj1Gz5J81OCF4o16RR4HuoYeYbvilXq1JgAy4+lvg
IQZ6jxPspb/6QQDGcS+PgJlqdwv+KQ0uoIOAxIcFkA+vntnsVwQqdXrqLVBY4kt/9G1M5bEKTGPM
3R38DJyYZrNiryJE+0IuD3o72BUI/kvMR+idFiGmj1FPn/F/C1otg7a17DeDi9V0oiCAzx8ca3cY
iuRzXspYETy5/sjEPsvktwcUH31AfuUM6FY1knvWt7pUl9ekOUm1cJXrqgOc67ce3jDKxpaWHe97
nSmDmfHtdwe6tkXNiBe+Ote4DOnplgZ7SeV18K3Ol8xIVodsyOFuI7T2p7C2jpXas5kbo4IwYZyg
dIvF0pZ3R58ubWY//yZFF/y0XoETnD7g4sSeeYU5HvIz1cRSGhETCpodaG86betkK1RoCsp1eEVe
I/fk+ClwKxfXpmhL1RlKluXNcpTppgA8YMndQjHNIyxcsviJefSgLQEj90pPujyqJo20tTOypsEP
xYW/U0rqmT3DkPG3hI8EXH/DGzOjzx5if1M3yCL6hHjsjLoBgB9kxdptTdEFImr6NiQTaRGOzTMh
IfzCHB/gHz6P8uIcdX7V4k+Uqqd0vmKbOigMDA+n5KuSe8lillhVqE60xKhHDmVwiHQW6JwXnRbT
eaCcKZh/IcszjzcYBNqrC94n2IGMi8O6P79a8KN/ffGJey0gl9ppaplL8RMgzWu6NH/PmlAiowp5
29lb1TsKym6C4+/IbaWfs1OuEA/XSdRYa2gGq9H62u82rLtiDhWx6x2U+23a1bib3enqq8uFSWDt
vvdOIEBvIjmJiu9E1CVUYkw+ENt2G0ndUhatac9F/TkStd4L9Hk78QCT5uUwTK4xV+jrPAxiTEdt
l7vazFvPXBZJUoPOQDp5LHa8cxOnQ/f6BM6Wd2Epj0zP41suwJKC3f+2iXmqeuuTCsHtnveuQYXU
MdamrRPSH0LfO/IAAIO2lQt69c1+2CRk+x9nkipO4k/chkKR8x601bM2R4sbuCngPpBz44ToLj6S
39VKeFNg403NtJ/ltwR5PQ9EZcYO2N+LNvZ8PVoI/4ob7rmRkDql/e6qCM1Ty00OUmsR27Y1AKyn
Y+swHFo9GbfKwMp/VaETAHMwSGLWu9G0AUJ11DlFsQlfOk5+ZjNr1uDlaUHWvYROmATTykCGtS8m
yPxLZs5+1B1kYFkgV/HDs4Im6FFkHr8gVDffp4ZAnmzhh6r7Z/7bM//tqQwJA1ahdRAvmiFuiasu
n6wUYignM4ZJdClKHqJQk/a4dYT47WknIV8A+XvMQKW9rbvHc8yaCNa8BGi508+EUFXLushzRjv3
30NaxFfV99XLKyyID8tMfoqZCX0mRBRzV4h0g3JsBFc/QCIaAOF7Dg3Mx3YM+l6/cT2DScuWNc2N
WE57RScYR5GRGTnwYSvFi97IJFsiz2NhkQSZ1ghz+ddGMMhhXYgo4R4sEE3pYyw7UIePQEgVj6jJ
3ZKAVyX/kASITcrORyXyIOhO5kqakt8rPBwO5Z205edouO/oZxdVTpf2IIvm9WL026Ro+K3nS+Cd
IMIv4waAW/jF2uxN6GPm+arxSMJfpEl4iDQfSIdekrUvjHMPM6bUfYZXIymRfowGtFXU5fxR2pjJ
OFMjhJ/tjmeX+QsRpx7riqAY3GQf3gRXjpIVHvtFcS1MXZD0TK11O41aUUuEM/Nh+Ic+NlRcJqDB
YvvQ42G6a443obeRvKL+zWI6fTLt2KDomkHDn+4lktwxxyvkJ6Cc3D+5AH7BZZOjVHOfAHQdfAl6
IRlaN1ZeHE6mbObRwSjNeYxbWOH80vR1BAPvfHRgFkMsxEMCPeT60xXETKYXvEbUux/ZLDxvLxqy
VOYKohWK0TW0144PLnWgJRoPMN+US7iUtudSCXs8iFABxZlu5zsRUH34Ccdnr+zMDgf+Jtc7kiKF
nUgQQvEwcSYmrYPKnmnpDO2E0oGg1t3+qyZDUggWp428672Kb7TnkKSvfuzBzPaby36ttl6XCzxs
ARacKCrDwPqdE2zvOVe7qBLR5Ybvij4XaW5cFxb4rMqr9fAgeib1DPQN2k0vNJ3Z03ENCJlB9jqW
rL+XR3O2RaeLzk9Jz5jXRLY8GU1LAlBzs4a+LYsLVInKqMWgjC+L6HPUkn59HyaHF4d36Xi14kPi
8b7kY4L1+ZVztgLb4cSzZ0Gqzu+sjgfRdWodrPwGWtm/WObyI880oSAcgLJ8xa20iHlqQU+eLfXs
WJaP7Z9O0A6IKCT+fcNK2CLV9bLeY1uaNOvEIGo4C9D13+cGSjmi8E5OpKDW5ahY8LiDP+BYfkYC
UXViNdJTfmU+hw1vXG12tQt2ppoz5Go4eeSlWt5kWUjYehuL/WRWh3JfqeVRk5DEZFfSgCxCoh2o
ata81z+I1qaw6Iy1yujiyuuIm9AAfmueW8mhPRVFHl8Q6RkZ0wGJXkfyoU/5fkNa45ONNIL+QTSU
T28SIpOpbyyVprkZ0cmiPza+zzC48Vk+QGiiuEnCY6Kqaqp+TeCJJ9mRYj7EvOB/muCrBg7wUa5C
Y9IOZkAmp+5kdh3/QKhkcLVAn7ZdLa9t3U+Z8LjeJHuGD9zATMaXFgNzFDpwL9U9jqdH3q5E6lfo
m8Tp6rIvGAdpbY8LNGvfgcyd33PdJWRRyco2cTbHoA0DOzTxxoX0zgzibPRR8JNdhykjG5dD7GmI
2qMZHZ6O3TQ9gGre8B2dGgsTLsR9CFTpcnhRqpRjOZqbToouRuvtIaSe8tBlHwCI4CIkTqwcIT06
0Sb5TYZZmSKdZZtlkSxsjTroGMi89cQV4pYgTHniXwkmBcq5yC1lpHwnv7DX/Z2Syj0EAh/NGBh1
mF3s6Bx/Bg6At8kEjiCflEX/tHjaatxDXKlsmGx98GigqM/TEhZqj5xOLa/UqeoEL9D/zFZr8vv/
pn09kdsqWowCFEm5oaOnr8dnzhi0JKji9is5wLHb4K31ry2tzwrMLOVGA79njSpkTG2hSvpAP1v9
xYZjzXHKAElHrGNyd7iuD3rVXDScCh9Jo9QcapFo/i85amm76yu/OCCSvMOzYc2uxt/2O/nvI03J
82fjfh4hAU2pwQMJZoB/JTsnSbiE8fW+H4OscV5FyI2P7CyWDfq8f2irAMvcEsM2DTuOeWgEZEPK
hDcQ9Riu+L3tRX8P+LOHXOh+a7ds/5ClHZxhUazuF75GpQKIM8P5cD3NG4k09aQ3Kix6703HsFrJ
X+ObzLGaqJFhaiqwFIbWKZsLHqGh/gYQoF3yBM50zIkIYm67Pp+hFMuVPnVc+NItvJ/dophYEEc9
OzChh1NDytUZXPlqC94FHoGsb1kbOGRik1bfKH7IbLQS9pQ/cd1J+5F9FBB8MJaDNrFEv3LN2Dfa
PfxnCE/76G9KHNaDR1cT31DyeobfjsUFBhQSrI+qSkjBT8jdGgObdAPRcDMjxTnacTPPVmDVYyT6
EJ+2gWnQzbfM/iYD7e6iYrtctDIHXudd72n7DPBHdvJ5NalpepanoilW0CDtjQwkYVHFLy8fiIAG
qkj7SEpgBrt5iXFEUbOntjFCeXCcRkXK7fJxYaJWAdw1Y3alrFAJRohY8db87NHWNzEaDgubU3P7
qxj4ZYYzWOPBZ40fCatS9ELMw6/86iv0O3ePldpwlJ6VI7fk/aTx0dCx/hyWxbDHr7RCAgTQiKrc
1vA4Ree20TmCV9HoduZQ+L+6UKDBTCfHPbUhKp63LtkoV7AB8r4mlSzrBMGcerDI5KGcV70a/h10
t/kYYf+Ywo/I/fowamwxrA297H5cn207UE8KkYYCQOaGq+cjFEAN1Nj2Y10C8OlgOqrdlH+kIC9g
HDp/SSm+c9lDIzQWwv3LRtbPidIwGrFGd6uj9c+ZQz/FMUtF+zHJNpf3KWZMMHL/vu23K/2RA+VQ
1cLwPanXzWPzaGqvBXh7Pc9k86H2nlVycu7FMGLbyECkIlb9dr59Qc9qNMUBSJiSL62HeKCzQ8bJ
IjgZo4BiRsoq3Il7Zhp6Ec/q16NI9A7bkjBn+HbjzcjGy9hBfsuvGA49E8iIin/uKsYeyYjKTdJY
KFtvTNFOhzbT1+hqN4pWaYcvtzEMN3raEk1+N/i3AN2ToCIDtXxo/5rpz+/xB/ucwW8S73a/mz6b
RvpSthv23pf5TYNSoliY53FZae1xchu1CN7+/FLRJTy7AZaYYnQsbvZ4xA3dFw1jfFYo9Vn8ZoLZ
voxgBRD4w7xr24w5M2UctETfon9GJbm6xeHTVOJE8bVd1lJahSOQJynJjgBZq5qykiBuIuaXdh1m
v3ruF6Bp435mxlEb0JgU6RGSq2NDP/TjCsHzcWz+NW2GA8smtlcoPepzlvJrpOmwpo55X6YVfrNK
MCMZRW5LrL34lyucozBiVrEhdGoZswMQHWdMZjwUQDmgZ9S1LdgB4pKr8/OrQGExA/sR7k3noiWG
qdoJ7IyEJi4vh7QxIa8eqAjRkNBu7L1woqA+NcogCqC21M0iP3gss228rEexoq9NSBDCYlcsjB4n
x2kOaaQhglaMJB65Ho6YATvhfePOfwNFhI7EneWD7fCP+9D31pzpZrIK06n3cSP0slOOPXXniw+A
3pIt/WCSnC3RjM/qWEy8Yxl3rtMfEMyNtQa6woGvdZ9D3qR0K5/bnCOoQ/CeXQaKIv5ZmGRZloZT
uWkE7OVeaeqiiMlL0iECHz0oLEzDCZRFN3iTQ8YGPh0U0MGhylrn/CFDQMuLBfUAJvKV2BA+ICXl
k1d6iX5QURYbjxGcT8mmTMHE0HHg8j5gm//VQfvyEo0XK5Iz6BTWJGjgbGQeWWYgZ7u5YHvGb/ub
IOG/k21O8ZhUCC6c475w2TK2QyiTzvf/SnONbOnXivjea5QVAvWF/brqFZhrLYc6bTzXVrGVo5YE
sLPQtWV7H2hEer+xAr6P5hfzSeDEPPAv9mXGSkSVO/q15BP3G6vpzCarAPcRQqT14GbOAc1wtMTA
fpHXGHXVonfkQIVqiS1rBcXSIsXla4yqrztFDvf3v6g/B0vb+6nkwpf9U7YMokrNit80xsOzjHOF
F3zpowOpjj2RhJLFct0GZL6uH/sfSu0PLrlfUuNkkoUTwbdNiNjNBPG43C9m7fHPRe6tkoaGOMye
wzRPoPFp+0pvGvOkBaGw3dxO8TSEWtPT9mv2nNqOqIlURFKyyDcpKyNdMGVgZgKIRbiAYqELfeKH
ZwHLmP2snRQCbAGcWMaXRrlzvO/Db11WC3IXpb25sFO9Ic3puWS/SiYot8EpHlDH6e0Qk1UQXRcz
9x07gdKeVMxxwWOFXHrE+H1B7vA1leLJw2PmmKOOXntzGlU1qAkvq7Mra5p7h4B7EF92ziwzyPcx
pu9d4Z6cxlhdHiUohXkeZjd05bUKMSE1rpGdIKIJntpM7rpEKjfdfjjoC743aZib95BaVlrCBLqI
Gd+kfJHdFN86Ipxx0wp1dQ8j0qLUu0Uhu4fU3c1laT+uAC9pBtT5/iIWdEB6CeYEoQd6Pktz2eV5
7iOHlqme3nx+VJ6suJiOwlPEbudZHagb53jb8wLTzjT2cUNeCFavt9evyr8fauWd9Gzna3J0/vou
xknPwSdCo7jt9jUCcg7b3bX79PXV4MyWwJxrC2oEGgrKx/MggL5ibQeB0bu2i+md721nvHZTn994
DejQ+F/bRdG5Hi9kTB1nw5BTt20xuYK+ZQ+N+WgqOPm6nX/z+56mYYEXpc/s8bZXndR1V5oPJBfI
d8DBLgicvS8TViCC7MUyL6jLU1HwGYD+T/wA/hLKToCyIgT7EbNNRWyCwsbbSwOoHxjeEaW+u4Ya
D/L2NSuxOwysbT32MZbUHVRHQFdt6gS+hRrKGlkhX/a8a8LTygO95h/5V7KWqE8UfqbUyQB+0Xfe
FNOYpmFV0PcXIPaamceVWC7PzYLgzW6GS5Um4a9cjMiMXG5EZ03VgexD/XgBcULw+S/luN2f8YpE
snouc986kR6Kk0pw8oIPhvCI2/HurFqsX1+8J+OpOvMTq7Q6r3lGkg87C2HWItXKC17fNYuzg2aP
1fHkLtKR+6R1xuvcAZaECZVP1llIsVYD/CS4bUHNrRjUjTlZXIw/Apv0AMSHllwCAnaR5zOG48Vy
lkTeMK1Zyls9mLuaY4EX1zmZIE6rP9OIziFUFkKXaH+Se+0SBhJjBDdsiSuZCmU/1kBMsshr6dS5
ylCpOFvCuyQ8fDVskpg55m82Edc29QsWY4K2MdVWx8lxsKv0sBOG+1urr8kF6Co4aMZ3xOdwRwXc
VHQ4p+3yERFh28J5/h7qyfRTkDylx7JzH0EHjVCGUY910i6PzhGGGnhOHsp5R5VFQ+66SSU3oMCO
nTeatYLVEO54qd02cD7jR04GIWhIsJwtTxJr8jcVtSenr7wJ1egJJld8/Id546IZJnydTod8RdJj
uVDjwoHoqJDeWH2oTZ1MaeaHpFoyrGTSoy7ZFi9wUAm+w5LdibTI/2Kw66pahUm5CYypJKCiCxtS
btPxSkyFUJvDVg9YYqX+zgInCTp2iFBlKI5U1vvGhE8Xix4hnepgSzzZnNnGJVcoM/Ym7Uu4iMqq
QKwTwz9buPpC92JWLMumE15u0Ej37XUXfV6Hq2GimH1joCjoZ29mz7crnTJt90zQ0Mbru2DPKdja
LfLYr6+3PTaX2bkIhnXJglNS6XmuIUEu+XF6S8+Wf9gsz0L2KrELmb2FghF/AbI/XfhudiJvBwmx
drzfUSzAX7SVN2fQEaRIPrwW+m4GGz6Riub8uw0ovnH7chSLNTk13gYVh1+irT/dzKYNs6vQTze9
LhE639kXBhlCtzCy4KkWsQJJ8Pzs1PvujOqMAAAegMdkNI9XUTPXSp/kQ0hsHfgQRusJWNGEaBwQ
6u8o7Hv0pLnn05BICSnBfJfM0Nwe7aZSfO6yMQIP1SMpMHqH85GXgwYlIa9vI2pa6plvgoa4AaTs
TDwwCGwEMY/IN+DXpFBUdjxPxXa5a67FRrd6H5vdtvtXapVowTSIFX0+qveWAGFIEMUgu6qI8RdE
hvpl6U3CSY60VkVxVFg9c8whO9OiCr2+dsKoW5nEk++g42QSUvGajGEDNjvz1e0SZwQEEmAER+bK
4Fzq9V/WSAY9/jTTVS5ujMTZGFUmvXTvpNKLP2ZYUDBF7yi9Z+Nle5OAHhRg0VBAAo3y6H3LBKcx
zzHM0Rzp+EudlLB2q7mIEpuqWUzcVbwnOqykf4Y47XKh2EDJEnv/gQnpMhBv9gPxlYKevoXeb4kN
j0V8rYKnyVF2Fs9fq5dRx5qWZcEVMyMrML1DOq7bbMBk34Qqu1kq0ZY80jkyd30jZWdqyPVixyQ0
DeMO7Apren+ieqRx9GL4XwxiSwngzHvONfb/ut0D0/athM5y97cO+ZPEi3ZEwAM94N/vB0TDGULP
mIdRYKvttFYAboeFTjsYgX0JNnyaFfyQwtfOPsIo6JrqG+UaWASFegXvjoH3p4P2SnAPXkU/dVG/
xchwnDvbRPQPnMrZG66KIWkLhqTY1T1MxjzNsdpGID2iqWJSiGdYsFWciZpcxlqw38bgBi0qmV0A
gJh8OfaQUMNfWI+HdTzQAEDC9hgIsIZj8FOENRdzL5XyzegwTLNTgcCX7S7DsngGQbeI5liVnkTR
JNQ3QMysTOOaMgaGV9VLuSwUupmkOkRshQphnLURZ22VAhheRRNqptesosBJc1E0d3YrsKUM3eBd
F7j97VAtPVxDBP28ziZYECymmbfqNOTP0BJmKv2ARSMQ1aXNaIH2cHLpoILtIQD63iF2GvLZSmnv
tSLAwhfUheggY7QYVGPOgYzlGWr+0RZq3129ABlBbg6ZK4cE7a1pu9ZQG8kkfnQ6AzegVTMU585E
B75lD8sco11Xra5OekdjXzYphxx9n+WUQc5MGTXr/aQ284ibgEtonDTzGsg39D96R5ax0Qoxrj2r
v9cJT3/2mQMYtbAAWS9jryX60zy3BIy+qkQuWCm3TLxAm8YaeEc4GFJ/UN+XNctn1KZAp1vTewyN
FZajNZauOLNJihVFTlCFuVcMQKOTjZkjXRgjxld82sXvDU0UZ4eir54nalGfEAJj/4WfCFj8fIDR
TVIfIVZra98gihgNPiCRGEzqTlpsVuqIRkKIAuCDbu6RXDou5NFl1Ym1ygRXAWdRhHbkBmcJpu1R
q5ZZyPArzzWuLPhjwhvKktYT3xap6qt5TtNBCbFzwWTV5AqCN58to287rXzJxPt6iAWDojSmsatN
YoxNK23m49FrDtzd5D2IFD7Avend9OrIoOEmOoGeKmJRRZo7sru46Fv6UIXpZnXzt5fnMkCPEedi
aNBfZtqgV6eD5NDFERu6g+9i5Lbeefe0kB5KEX3ZIcdXwb34wlb7ZiED+g555NTtVHVovstD2uCy
n26mIC3DnR6P/IIx8BI0kXLxz3dxiS91SlNayOpVHSTHOtnHmOn5RWmD3O/FcsnUnNDDpeal5UVa
RldR5Rg/qj0JPp9gtsUh5Uu9deDdBSBMXHCNYNZ4GrqNkKxqCF6wD/vFD4NV8yEsok0uCP7hhji2
1Xq/efQeClbscV797t0tl795M/cwTmL85KqOCK+1kEv1wc1l2yvSpgK4zXvjPKt4MLSrlYRqM/IX
+xfGMDyxyHNIGlRosHx2+1B+WprzMJWQyaq/1mjzA0l+qKmL1W3ET5KD5hCA71/km7FfAtOl63U6
H+lHZ58+MFDj/Aj9fSAHaBGXPEEfqbMaabdwcKJ1rnsoWT0ZpX/ij5GFGAJ92v9Y033n5yZOMYt1
H0MTqsjPNUzkEngg/tevRAED7QwY0KcDvGukP2/Zxgg0riu0Sr1CFepR+yNCxuDo5yynyodKMNxM
gH5smZECElNPR+mCBpnQFJC5d/Gv898x71Xmav9tlrMUQaZD1cSrcFfVLSKAt+IwNYLtWZCSu/Nr
DgLmHrk8QxwCYXyJp6ct6eCJVPJ6Iq6rZT72vzU18aX/bhEe/qfDYlXsZM4AB6M0Dxb9TUFKFmYV
MFIw3D2usDuWmZ7bOwNoCg6SpGqlIEnQxK0ekQTcVa28MVzs43o4e/T+bnamcYrRTx112Hat+sub
u0NEQWn7xpSBdOBsRlY3SWZwYTwdxXC9e/knso/SfW69M8ps7LdOI7SF9dBKhlq+9dcKEaCNh3ah
/GTe2ezRc4MdVUo8ctMtkTulg+n0vCpGLVwpD7uWZk9zOipi7IT2iNWIv5D0Q6gvMoxpXq2ys/JJ
0HTdhiCYxwBZQABGPaVIY5gAD7oHnedqz8Uc/xhzfnxiMt4eEn9h0pBvXWsiLJbQHdtBilbKzGB9
9JF4WRjIsySZ19U97oVMYA+kcWzikRKaScDEv8iRuxVLg/+A79pHfjF0nFBcC+BYVWQ/xx4IUHdx
4MAUy9LM7Uyp6+qV7baQBcHgX5Qam0KsiwM2XX08Xl1PigsYVd1CH9anpYUk293SwihntgrAWD2y
OK9gxylavI/i4FikWhQ3QZZxGv6pvpqw5sC/62Lg7PCJ2gE7cx3iELlwtwKSiHbnzGLT8HuE5RXj
AYmECF+6jfFNMsfcqjl1f0TyumSg2+GRaDqjk1XyDSX/vsiLgXKpC/tr1QWpu9Qk3yC2m9OtLeTY
5sQCKhULvrlUQiQuqVJX8GnwbZlYXx7Fj4GkewYCclhsw/Ygeypu4UZoCsYgcNssK5dy3t9e87Cw
ITTHVWX6NBdnxWS6IeQPKSj8KXPVWJrQrg+SuXPnYL6DFWBk1xnC3TjOQ+ZOWQIVEZORajpJirtZ
sEPFLqu6olC1KTkV24yRiuGousg7ZyhqJcSkfFW8dr58C1o1BEpHPg+AI7wEdlGAHrWgBVV9ikjn
mdg5n/eF2w8Dr/BQpAJ1Uj+I6QhHqkrxq70ob3WMRTLqG5Olp90I+jfzkY2n1lldaTJNmyDdXDpc
9BzGDiUgyGceWDJCNtqaDXzOo7+/j8YlhSVpx+HE2qqwwtv61feqgQfZ1UKocJap8rKVyrGTvwLA
I07I8mikgie3VZfGBiy9CybNMpA3CXvn56xeP+5WlzKT9Jo6B23wiXI4W+aHaZlYyZ1HBIW7HAX7
zp/06BdDIKSzNOd1hiIX61Xxg9rIQMInersEfjkN1uTHdbURAb602DnlXmYRGFj2OgpXkYXNCamA
t/o7z8thM1vNL4F5cIOum7jVHU6f3GvQM48bu5Iimx7HfznSgnHHN1CgVVMaOHSeG3N60QRRFIKA
RZRkb02MiepUJVPDxgMqLrAYfuZMQ9u82X6gykJKVrRzpzHLln72lndCn6RLCe/kAY5ds7VRaVAR
VVji68yWSYtkSzmQMKkXDiouyWmOJDK2mc2SPKUB3e4X6E11f8kFIjp7bJCptbbUMLeQmmDn+B9N
Nrgtnjoxhq5hSJAtl6a76vlJmBVJN97nL4MAT/XkjqktB22UlTbwgZCKZ9f2LnDyCw270B+ymnFQ
pIpzhT0BP9gjjgy9SBMoAqoeYe9rG7rpoFUXI2rVPtob5tvbvK5HB7hoDEy7ZTpCilfHsyq/zqiq
Om1guSA3tyxGm/tLVaViC3WcP0l9nb/UAw4soB/qvedIZYIKG9FpFxV7DT8bKqVWb0rYGHpe9Scn
c0XhrrOOj3SWUnwm1VGAXkegLplj4rMs/xLlgQT5Yg5daR83RIuXu7SRWSXVluujUeL2cPuMqtgj
KTL4Xt8uvjn/N0U+hWoWz61MpuDmiyNC/anOfmMmIge1B3LY9AWCyhrk/tP70+uWb85j4QtIa7zl
bpedXkUJcVLbHya+Ik4cImj3xCC0PqAB5llbwFDXl8wtFl1t/plnwyVPtxUQgDpe6BvNkpIWo7Kh
DKWIgPe2gCLVG4MUc4MtpBHKrkWll3HC94AaK3zek6v3s5eDvOauJu+kg73PvdI3Go/vcP3x9NgH
1hpUnALi4LeNNP/jlwd7DGj7VxvDQUWF26VMf0VDSm1+gPPIJBGR/QSy3yMCBcxSxqmRvlBt0iOL
D5n0D9eylaSmGeDDPsmEPYgoCteilryUMv3fqGpZhHEDtzSVE7EV1EvpFa+yA82grIS86MnzVOpm
49R39POWU+Zz+yQaYcq40FYr6PTGFLL0/N12EtMgOtKEWeuETMFXh+wytw2SXvZGM9iIUji++DUv
j+rHcwv5791SJgMWT258PKOhCAxuSfHRMat+lVsVyIqpOmAYFnSchMTji/0Yw3YlwJpIhkkQfXug
qK9OdcHUJOpsRGoY0q1bNkg/Z27xM758qFGL9qTVCPhbZlTfSvZ+Lkmvnyb47RCsV6KHluQdrhb+
U0JKFFLHHmPaTExScLjdWnzWoYD/zFPUKca6ai/XpEp2P3JFhKMrxuFzsmq16I/QifaR2otml8Uc
xrx2kLPqLoYJdj19wFeCx0CKNh8hhoaAwfRXzsnZQtcx8ThENfok66Bgbwyo50wplw6QT8GgeH5H
TWzhba91MmeUzVPBiBBBe8RdzewEUDqwlido4XpYwDk8WQaneYZTHaI6NpmCh/ca6IM04X0gczm2
2Z0I1SbDGoBNSSE6WBFsb/DDGEDed/buPOmHt29mPVNLD1upQIM5XspS96sSXaMMMH078eS2mnkh
jcv8oMB2l71s4u6gQ6L0uGEurXpUqKtfMPP/qwipn8RK+0mXlwqsSKz0sEKiUBfOgpcxh3PsX8tS
2dAgwqS+N90LL6cONrIEXTCt/HQGcPUZQWiMwXJVHopPi4oqS3pY55C4HFyGcTb+C20LJbVASe9E
9F2gZhKzC3kAvWMLeRXpPql3rdXPQ27KRBgrRNp79uWhLFILKfh+gB3i5ZDy+mi7OcSDzvx1zk4g
IZTJodQYZO9WZicUtBGmDkMEGdXXuzVa6E1k1fbYy7Qpy/KQPSfTG3D02Dnm99z5OORklp7DHxQm
uDGKjWO50YEm/Qyzy/jsZ0zZRCj3d8RFX2vKoB1fWe2najfHY5+zL9nFvRyHKKmXI1+WliabvmFl
xtcMc9CAAb4dBf3QQt5Hve4eBzh9LhFdJ2PTXLEnulkCrXW3OtfTqqwWucjLCoiuuK0kxOPwD1WO
Z5mhyrulEpR0Kd2TDXycIp3ztR72uuAnVss2Y41vwW5DKvUuXE+py6EKhtRcp8v0Bk839vUdKOFA
6YFUErHjKjjtbBjJgrj1fxJak8xatpA+TWWb13EavqLqE0/BKHB3gG/YGUkcrbMbLsqcA5tBVPBr
meT5Lwiq10hXzK795icMBvdE4o+Ej1r1/gAmlmSQa1WZ2vpdgQ9TZUeZzg+5hIZJf/l9KcAAeDnr
EMCnrNa/d8AMlwdv2XBQ39kE6gZN+Arlhu+NR0Jt5W4w/x1B9vU48FJcMC5xJcN637fF2rfoUKrl
jx5x/ziCt2r/GX1lzmseBANfBya4nsrPHxTLafD5Eur3L1lc6aaJzPsRT/xCPeQlvlCuWUjxcyOJ
Gun+AqoNn6eIn80QfyknlrU/f9ZS0Kj6o6jdHdr8nIQlgSBGg27PjnGNmx/zIwEco1fe0JsjzIzi
s2EmLzrYSa0+Kh1l6ARUjra9pDMBgMNb0M9C1qepcWKPR5M2B3cktdQAb4TmaSHN6psP2QD4YYLZ
k0vPGoJwHQ5hxCxb2iBeY15SYNGKhVVw090VDpPoFgU2FeXEJ+NnlMUWhKzXLWzxaVl/Qpiw1m+o
enOfp72twBoKekCl91AZ72zEQ6EvqjZW69AUttDRnESJtQikqqLE/D/t51GsXTV5FMDPb0RC6lfP
Q4Bno+R1IHpjdYtywQTmp3v7iV2XK7zOFArGPye8Izu7X6iuw+B4hwFZm32tFWtZ8ISgYk1NmKvs
MsUkwjYdKxzHZxQcLANmwF5v3byuBLAY5DEHsDZ8n5932ogFOcqala5/8AoBn7mP88DWbZxrrvZF
/HHAj/mQSLQ2p2/2RdQfkZgTQxlpVKYDgU8UH0el7NMKcLurdayuHa75uoVO5F2/+dqjU4HqSFij
/09c3hz4DlVtoW0Jan5Tp6VXNh7cAw7n+A4Fll+mOUxsyKWyYsd33D40ynUXEsKbHzTT5pv1qd//
SEwL3S62pGFOQ+vaaakUtmrvB8PsRVEgmGCV3AqVZ7vbnWI6gzBlD5ScI9Ve6FmGhMjcAPr3e/dg
Q3V17fK55W10xxr241+OGBUCeGBVVTvc5UebArpHY/1ncXJBENYt6VzVTnNYTsK9NGj+TbfU7zy1
2ORGM1fMYKv7FEiXkoANptWD885IuFCBGrFaQi/inm57hKvddUEjNy7ntgA/gD9BPQPT/ns0Lqux
DOH/9eFfXCkLIwWPhEzmbCBmUiD4XULnPQDFes6HFZqVAkOOWcibglQ56p5+boLNCupiuu4HC3Cv
JLq9Kt9GdVG6zdMKSRb1ia/95Z8riE78cZyCmo5Tvi2xCUg0Nx+JulxaMWE3/qU0PJdlvgX6XO8P
2WO2ByqTCu8wSkq3KIKFpKn9qCSJdvTFjp8RbicyY7N+Qpc7/Z1dvoOcgfR3PozHpkuYVH3AwU3X
QhmNfn9s/1psBVdGKIVkHrcsrlJuPcBWzu6P6dZ3ZGGk2wS1ORx5PEJrDoa4XVEwVUcp+5lsfhir
G2Gt7agyjy9mI8NEcurYKFChqx5NMHGn/pGf1q4zisWShYu3M+RsT5tWLWqbSvgP+MyoWuvKBzhm
rUOIpgVqix3Cqj5TiGR0oLoyj+Dt5D7wx83d2pwleNBMNb+9MlM2vCyZb6GPOWgt3qgfHDCCd0Z7
+OVXsCTT0sAQAMpXGJGt6z4kRE8gWU2nILvTHAvoY+uXy2ZK6UTtt0KHysZn3pnua5pF55+Q8aAa
nGzyZHlc+l0GMv33CNAJGiUj/0Aex+UlLsjR0Lvjfe3nrv4txf7HPCJCL3mkmLKYAJZVdh8wbvZ9
pQYqRKTLeemd2CwWx4KNPLr7Nk4cClJdeiyvXruC3bgyB8if3icB4u0s5F882JQKkxjsDZ/p6h1r
w1slVmBtfkAs1URZKxAfzyUgFgxsctMxfYnUPmQyUbcMdRaS+9n9y2gEUiocU9QLMVH+FcJv8vaE
ynTaAmrMfRHMwDIA4XoCGFHAB78ZASoOSLcnDmEsekR6Y/FgmyNMFT5IgXY8ehp5VU1tmGr9Gmvi
+VIKsMXwHtF9md8gzODnpQDcSAv8IGuB2CTTalvvnuIkkwjeqsfIaM2IA0wBM2YfJN2XnkRZd7n6
Sxz9EwIntvLrekZG0vyku/hDC8OZ5fj8H9TZ8XkhRtYj8F3BqqL+/b5y8vfgte5sbYIfmZevgFF9
6QGegiAhy1JMsvVeiXNUh2bwFw4UNzi+5kqvqcLp5qZsfJdKIhqLX+re1xOYd72ZY/n96iMVrHBZ
/8xdYhglc862UyhDRK9dhI4LAKFREWyDiWTQcG0KRZEg3kelQd9eBtRhh0Ft5rjrfEaUVQsEzS+x
vfXuP5G/zw71wc3ah3/w3R65YsazS+UwhIoxA7YlW0ZwEQxNlw8M/puATBu4/YfEwKbe0MPiuZCU
TjUEaB+muk7ho8Pwl1LenurgnRFqomHnz/9JKJX+AqWqh3xMVFIpOgz0xIWzzFSjbHzxl9LjdwVz
OZeLsMVS6z5dl7g8jqC2QLEudrjwip70QMKJpgwjwgM5sB5k/GoRmQSvAFu0hdRbOmbv+byiLa6/
82+ZWDxN9mStyxxRkSU12ifUJyVt2z0f7Q6tHdYfUu5HxNYc5LsGhXSV5nFvbDNMJRUHcNVPMzj7
VXVJRVXRAMWTgToZXnfhFocQur8p7x2yKdMr0+bfG1sFyacQiFsDY5uTtMa1I0FgtN+XNfAXyFjR
AeytnXQMHfRv9KQNTIbaukJzOEoJ+KX2TrmRnb33aPrkFfQOOMdBoHakZwn5bzsaVxW5hmRTyJI6
R9fai5mPpu3AC4Q2/CV8IkyjBwkPKnc05tw2Cj+LXWf9pgdeloBxgpOxEvmlQLD6hTG8OVPRHVnw
NJYeyEl7ZQkRC86bvhgqJSUePvxdKmQeXdKX5o4uBQRIIw0wdtoFwvWRsD0jkSOumaItII3WdDQ7
tla1v6YpA5PxzFeGKj9NpUFJzUHb23IlAy9zuOyOzntvBbkMsZmGCiWS3wLaKcOOwDnCY0oN+mzR
z9DQET9JhGKpN+e+VhuE0WTvQlN0UqXuJhaVAwhrCGMi1iBVSwpEyl5uEDt/IK2H97bDkDRiems0
IVXEOe5E8ruegjdxSauS3vi3x1ngXt9kA1l/7SeCd5NIP8UNbadA/GVm5kZGuIJ+QcSSJfzz++hg
C9LkScZVCZic5VyLLLXfiRl0WdLrZzoXa+8hF0hzJpQdUgHZxKbJ0BfrVQES7LB2iNk7fhsp6feU
Qnhd/7aSo2WHO4LcDtYuaTjBr+BO8qFp9spOZkxlmn7GtXEzWTFgQ2lykOQfJYEcJSW+yMwzsNP8
LC7VblXkaSueY12JuU0zpZLMG5qs/bOoYVT/MNhrOkYE2IpcAwNMewp8HAb4Y7ex1WVU8FDphLS4
+eE/sFMX9YosZLoHS7sY+CIb1ZK0YAH5k7v/lnNzaVyi3qOkcxDMn6+jvxjTQJShj345cS77n555
3cSBZ8FR6+ByI3IzqiNAXNG96bDxU4oJ2n2asOqk6XtOr6q8uzXoEhP77QT5H0kNPkJu2HBSCmwA
HTb6CyJxw4MpPwd+Rl9Qx8YPXSuie1ASsyOmx51MrKyKbH1IopK8QXktbWGlC1Kpgf9pVu8DYjFv
APXieDcxMkCqUap3ZK8e7+cVE0W2srCZE6wCxoMhg+n2JRu0Q/l1Pi/4Bf6Gk0pCZbh85ZSOb/iO
ib9Ep/6FWDa5ueTxYIU8439b+7CuWfEku0NRsiv7v6SJZfrB6Co7pwDb11Oddx+0sUgNU0ASBYOH
QHuZgbd9gMXClgYybzv+SvPpz24My9gboZpGDS+YGMoBsgDQaivDVPYTmwp1Bd3A4GAAB1tHguGU
btSDAszsnbg54I2yr3tSbwG4phUL8MehypZFJsda8fG1hogcOwfXBMXeRHwFy+1FBSHjnR2rtjKE
0Yv2enmDvMZXW8IgarjLaGzjBnevJk4eyTioXo/r1NHmjAHMRTi4ZwN9n6Io7yENzefTvooENjDh
/VQr6IfpM4O7oQGhpIW5h0s0GawarylTn+957M2SkgQZD0D9j8pSm3T1AC3fsil8pz/qw/R/Tj09
qhS0z8DZeMRWR5zWvwl2y4v3bjdGtmeCKia8CBMhT1hNtjUlFgfz5euecbF8CuwFxNHafy5fD16G
U1V4wlCfoljeq7ytXQApiuGRxFgTfHZOfPpa363gZLNnprWgrWlc1j5Y8jGsPu5qwnY5TI0oqRcm
775TmY3nnRlUTj7/cSBkPdIitFT3myFqHsu997jHjYp6TY38YTJBX/opYrCEq+wVhp2HRtJfVkqO
5gV7ttAQOthdQDDJCg9QdmHrWLB4X2vQtv2CX4xGmNTB/xR/pGQKBr+b3TEtQrIXefeE3NVG29Ys
cFklKw4f5OtGOKOMolv1xnf6Ow0tAbe9ZXxBh/lROCk9F/PkwA3iFFsydd2eB3bsSRqi1Lw0gR2N
U6c6lA/nDo1cd5kGNhK48RGIPLfPbb/f3WnV/tLNgMn7UGFFD6TxK6hYS6QXyek0oV3FUDkvMeNm
gOGSJeduEJHgcAVQzxMB6LZEEBiX9+0J3yY36jRfReMe5oKm9Z4A6EKmmXll1eJbwQ+8J7KGSXSC
rr5jSSKrZQ7Bo0hLisAY4hSve1Az/YFABkQMYqOF5yr0/iPzITG9GfbD280GcEDa3Z4HGkZKpIWo
aIqhFYFO6ppb4jTKrj0qSepY89CpPZxJ48zlaV01ZPnZ6qzGpZsLH4ZlKClbJrb5qd8ptluXw7Y8
4fbHrTsIEi2qGmnJQyM6vcaxj4z0/PW6T7boE1MBPcneriNYG6FgXNHQdfljXO3Rwobfk/HIaegl
qfXQjgrS+l2hNUXMt4eC/MEQgiXsxd6FT/CfUY5Y4zrRwFMTs/OjHtAcp9nMuyHB+YVfVXQztykl
NI/g3VZaaUTgHllx67dDMZBk2pcz6bHKAMzeYMZyzGwAOcvJxsfvV6zZ1i//Qp/spoQq/xKzT1Gc
N6RC83BcoMXhFBm8pf0d7PojCWnvb0rgX7u/4VKoPxtqQr+hCt7rMZk7OcZW3uoC/bIc8p3QjmoU
JIcByhBwDYr06SMACyHw2fDZrtyUyaJo75ryu5SSEVwg8y+z3cJ8tetPoQOtHyY92fIxEGKPy73b
QYJPXfGQidmNF0mvUGUbxij7ge1hOqy7KSzPj+H77L5rFcT+h79JsDepkB2E4t8SI1VvXP4/Bf7s
H/5h9qfjdkIf7et/7kuI9ly6mXTCQpPyqdBDx5OZtB7PfR9vAQLPqWeq1zhvN0s+Mj4QYOPv/9b+
25IKs0N6k2jyuxB7EZgiuoxydeMvydtew4wyZzp6x8GWEw+NBucn9+pR919Qq8pUQVJXoZaW9UN6
AHBKyGc75RLMOHP2SK/AEi0k0cVZQtcFHvLglKNvbfbc5dayMMyyiIEEDtkGI6i2JFCryDEMIeCG
YdNdetme9QxrHNKA/JfHXtoctqQbdQ9GXLhSDwbUAia6vsBdWApwARHW/xQTXVg88rTjsYhEUjGu
6L5/rtzSwB7scC7Hw43rmOyQ3m/NKjqj4Z9pMimAneyP01yN9+jOCl9CpuDu6IYn+mTrwWaELa0E
CpPtdws1wxZAjuzYlkKne2PkrcqvTLdPlIeO4Rw2lSMxsyoiSyHQe6J6pVtS64ov05XXg25ES3DY
J8WmJuJLpUwkoFMRKq1/9QCpEQOyWq+93Lw6cHlofW0apXM6LhLhFXN0DLw/BMXQHlqeMP4AqMOy
oWUhrqJrl8uDM5VPhkuXWJFtfkVmetKpAzcOk58Kw9uBr+q/C2SXkpgDOlysVu+XHJp3wgSlYUfz
4Eo5m/2/wK1fKG1DB7orf3vOGU+mAZQEXERsIHWdK0jx6v0mdoMoZ0i6ZixiIWZ5pQRP/ZjcpI4z
ZMv5uL1x4/wAl8MjhRNcVMNxH7SjT4W/b3uIrGb6hIbcg+znnByK0JRsg9KAMr6oVb2L30cxzg0s
4dWobJKNvypVnWMIOsVOaUoPpkNa2XmoesV9/whMhm/r29Og1LbnBSq9v8jBVtKkf81+mSTfkNoA
ZtXM5w/cx8wFldmEh3PG7pokDMa34k/4GZ6t547Yk/otg9diJ1XEgwnS/8cXP9p3HpiP/bq+Vr4S
liJK6EhU2XhU7C5k4idqM92cWilDuxSmV2GtL8B2PpTQNrZ9fIdROEjBEB0xbpfzbBf0M8t1XUjj
XnhWFBk8cFexqL/D3OdaHsp1oqfCHiED23JHDvyb2lGVEaE9EyrVlOIpKrT5Nc7aKUvXr5wwG+wd
6XBO9H6Gc7Yf+BITbQImlQGs7dXOKQt8RhzZF6nStF+ZZNWLU5IoFSOUfK9yRZMhGhyMfJ8O8y82
Mb4ue54keaq9KyqIDcABowk2sh/HMYy9BKjcI1+W4aW7lW7T8FawGH3NOaQxhEoZC8Jj3sv8AQ/F
/2aQzo4SmYwjCAaTWJa6eV/EZraawA5zHZJZxGmOYNYHxPVLWD05M0+ylBbQPPVkMYsnkjLbiJWy
dt4inF7JFq+2neFU/SNqWgmlrUKqcxwQ93gK42gfjacsR9JZq2a6iCjMBcAde9L2+CVebydk5UcE
Ni3/vc8iwa66chY2gGsFBah67pdqm5RoqEpl/xrOgHNXtJCQC3NH0AWTS+E//KuV6wswTz6e4msL
Y4Q+q9mQAWuoCE1SaJLxx2gnTBY1YULBMlcj+yZbmb9G3vwZO9KRYX3Ed2gXQCJIdt/fYeafG2cX
6v2WLIXQpzpZlrcvq9sDy4cyAko2NVN4KhUjfdYW+oMEXHf1rJf2GBmbw1odabVrwyDzIHV3uUul
xOaWQJXwyDpws/wm4rixsb2tBufyE1A8qDDhTHgafGqCl7CwAtSWBgq44kQsi32e3PMuxRDFcEiR
/My3IpB2gDQ2jOfP/AjLG9d1N4TRkNGTivFS2oHopq9KSCgq+rnjMc8t/O/u3oU6sO9/gOwZL8Rm
oTTxhg2+7tCv0tNTXm2+Ckkyd0lIqnvIcEXzlNsysCYttgjOTeKBBTLN4srsc+joZ/pC5XytXjYx
uNoIr94FUwQCJChdyRq99SlGigsmG2w3L3UEtQ+Ia5JS80HobZ7fGWjgRL1Ek3hE8lBSJbbQF0po
wiiKlpRemw6AvFA7Z0JdPmXQNOBB5tm7wf8soYT+woMnYyCFXx6DcxFm7gxUhvZ/WQjNLiBawbnt
QmB/cBucBBY4PIdXA3JqIdJpNx6f9jbRmtnsDKcR8ttZ+rrmzqFTjplfP4BYlLmKHE0YNQ4ajqyA
0PTUyNgQ21h1Lg5La0BPMCW86sInk9kTjtB/5p/f5kCfBJkEh/o2OuN8nhM6l9HLYcDgtvwSc9S/
R1xQKnZYBOSSOzfYU0/3ZsAR8Q3eotuWASbYb1J4DGjmb3yHGCYaKXVd19v1Vu4NZQfdu8WvO3Kj
w3TtYwj/ny1RRJc5pLYr3r/KXQwPXg7Y/9/fpL59uIFrWffQRrAsOruEYAhgDJbYFUUVKGKXmhgX
lIZRe/geplnP7GbR7/2wTXwS+oTHfNevUb65omyMWgjejhQR6q338g9Er+2w7igRqK08h/7HRpJ+
MnTiKNZs/tg2zaYfKqHUdweGA48yODF096Z5sP2RvT2H7OX44TeSZaYfw1VTxQEtnoq2iLKACvI4
XX6X/+5tcjQqD+mxdNjPCqGi94ldCVUdxj4WXjAm6A19er1qogaFPTaavftoHoJoLNYOVzHI/qo4
wXAQS9CKCShPwnspDgIET7UE5FIbmXLYqCcxEsPqMPfdbFYcx5cUDmGD/8ipSCPqAi9YnF450xsY
AhUPGzdaMETNxszuQp1FV494rRXGTz5+97S8BWA/mBZDxUHTZJMV6X9Ft45wNzcHEnrSBjQzUIDX
H3kYMdalAI82Xyq7mzrBuSbG6H/we9kpu3SV0stT0xA8DK5A21aNlnt5hqArOpdiVZ9HI7X+uL6w
m42Wb53PVGSwZLKwJ+q3Pkktd8oYqwkyhWQFq3HvReiS3D/JR69oVUhXrEjVWNAb8PxjQGCMfk3S
Gbi0x6dOcxsrUn4a5cLlK3AsHKaOKfz0SsADzsVgrX3vGnSsvrljKmGvb8M2RN8Kevlar7CsOWC8
MG+6o36aURgabKunyWgoJzplEFtUQL7DAa5NlXZiegmTpSoLUIN7m2czm6nXPzl5H7F16/Q+Jo9L
rSpJrPzYbyLqyJcR/vMRhjBkgoPaQseYrZQW3enPdRAmP2Bzk7p0myBE0n+rdcptIU7/l2jHaku9
dKYOTQF2ahx8KJgjc89pKLZVJtOrDIQr0fHbWB8RhDfYtea3SttlzSzXan9VAra5GBzeTRNYykSC
R6z3567MzS0DOXzFUI5fOsfV864UdV+/5MtKaeWxYtPutWhFQ3Nlpw9720bFlEUmVEsoXAi7U4rj
LztTlgt8vk1nWte4rfJXFvUSwfhDdI8Zy1WaybPEJkjaQIY+6JLzYEBRfgJTs70Y+yLWmye73Hoy
LF0RvKT9QieBTj0e4rQQhvaNWmNICULiGjf6eIIPuTsMBRZNIwb30nk5tsLf9Y4QfjIA8O3xAelF
ReyiaV9bBqC6Th4XzN4jRPwHuZDUpOU60AHxk2WqLBJmtxVnptIOCEDHYkMoAqjtg1NYZs1vf5VC
CuxG4nQ8hw+Xtq0q8LLP1zQSFrZHznMhN75sZD3pHKUIKWmfeFqEFTbbUOAvsYMcI+9pAmNGb1mV
3srsEOdxfW8kgFiENFyhbQfsYGmDRpl6EoFViolm0jU0+qGeDEqKsMUogBj5SqU/PUBxKGa4jV39
dFwW7yZEHoTVwf37DZpLsm22/noMEJYU92SuBrgXfZED+kED3HfaEvGYmxj0J8L7EknatyMeN2z5
cYis3u2/19Wp6SmbzeLGO1dUjDai35NEdq6bO35XiZArT8Nh+FzZdw4vbbOibeYX1ch2s64rcHLB
SK8DbPPb2yetEr+PORR1tOLQ2JV3kl+HUciAn87bF6d1w7QqLrOZUnm8SxXtGR9uLhspLRbTR3WU
x1j2Dk23WX/CRSom4WnQe66uuQDcsG95WNiHxB/eUF596LiNkuU56oMGrJeSlzkDD6cob87bHGUX
r1vjuap+bqp3W2wweTrfTsj19Au6vHRWMnirVCn6AIwX9XEu3x6V7mqWLaJ6kk+p6LbY7BpdVfc4
TH+APGiavA7y60e3eKQuiwsDiDz9JkooBV+WWFReIBw6G8DAtJs9b+6hnj350t5h3MCAn9meICPA
31JzskUKPxIHTRi3kseuqng6CsB9hHATKJRMaJGfTdV3lI/4Iw3LY4Gf55Yp+/MlwHQLVzKfFrzR
zoe6M6LxrI72BLOOavUFiW7aOR2XqlgTedzniZURfDALr8xxA4eF3ZnevWgKW0eGNZ0RYDeqcshh
0R5bwTd9UEDQi9qhh3/5HOxG98hHW7L61SsnU+vyVrHnY1l82qhZNX5JmS+B6Ll4SNhhJd+of7vn
aoJ2FoiSkrz1jEPn5bsV+cvY0RHFF9mRiwL3Hrj/9Rc6Orna4yGQcDYGrPyd+dh1BLkOIpAKdXih
qOWrvCNOOX/Dda1HxjgSDl3LfmPPfs3yc5BpxhtdHClIvuUCNVPjmtWJR7g9CbUduIpAPN25N8LD
BIddKKWMvkYnjCTUhYaew98BUaONYLwkO36lMRRy2thwep2C411VLL27plbr9fO/V7QlsRZe//hl
S6oECFRf9A8cM4j1AvAMoX/QUOdNGSti9X6lSODZhioU1gI/cgvn6KaN8BZhOf+UsamGLBS1mayB
EnbkNDGmvcIf9mKL3YUwQDhoZ98B27uG0MC0mRHh1awBqDjggQK8U9HYnPFYXZikxPmV/bZc/E8w
Ijg4d5SF1e6zeY1fvRACxPyGNQq+TGFoTClB0AyM/ecIzWR35iNFwGoik1yJxCb5YoAY+E6hzZGF
Fp/pMQoLne+kQUL2pYkSXuXeTzQl2lrKBiAV+4RCL/b5USF9bLkWUoxSKfBpYX41pnkURVg+Xn8T
znkN7nPgzJDyZ8t1A5ayRhvtqoz1DKi47FR0OVLBAIlBv6EBpzfZ9v2C9nga3+/ZOEMWoVg+nL7N
7VJB00eoKGyOvJbzhrWjgwy76C8mTSqWyhqLuD0fkitc7oDoz67F/3ARKVSCEJooSyp7iTzscHzz
18J38oAZYhRBzybY0d2CE5ESbZdPBjDaZ3EhgzfSURldEi93quDN5om3HP8PGiExWz1kgMwSANAL
txaYZ8tsIAfpfg42IQ4sKkzQkH0VhpQjog/zqlYT57BcNy10tKPrtbDRPHoZw67FoJANC/mkWye4
YmhcQ/In9XzhFf5OeKjUOjL+Gj/Rl9BmBMJO47l5sWZGo+c+aNEqG7rCw07A6NPxEK+3KbszZqtK
NMlzHA219FnXsDIwUV3xbMso0wmt8VWiM0tXU/iPC/Y0z2IRT5x2H0GJ546e34491Q0jUzBozZvn
RrkZMKEFwOrbLR0ahAwZwvO/7Js2bqUwuF929YbfttnNlKFZAEk634GleAXarImeu30/yXkCccj1
VxoV9WBJVNvxHSVeaI1+mvJ78dpZbhpTxDEzBP1Hs9J1J3/PPS3nn4hRRckcb/WziQ6DhK2Z/nCv
5p6Tn4ErVP1A90v4jItgtwiUopMowai2/dKKcVGJbwp4PTQ27sM0jIHy9LkOsT41pNc0HnEI3LGA
EzMAch3IlN/8zZFBEKgVRSUAOSfnUU/S+Jfpw4fsOa5PByZpITfRxjgAYncS1Y6zC+eg1TI4Ss6b
JbVzWoRoanTveAnWvEcxgM9tyFzFlQyppIz4FwUD2y+ymlN1XAtSTHjT6KBPqyOZY4sjZmhv9oro
EvlVKwhfzFMdmzg0hwbZC2ndoHaZxt28qjW3U3hcpoADR1yJhSYFvlMzfkc4fbL8lNH0ynfLDxhE
/BCnpv4mswzV2kzIp5YjVFXd7khpJSdgba3eIFxejQxiSP1sWT/v5iIMJ830L/TeNFz5aXPlkKWD
rh8DE0QVZ5lWXCPo/CStIT20u3sdsZJhU539dc1mGxBrA60096nXdiA+hOOdLlXYganj2kbKFnTn
FBmIlJiXfYqPN7O0tlC2YDvWT2pCFTdYU5Vg100W1WiqA5hixsQiH+4tYk40Kuo8jn7/+9ZJJf11
4+XuakXfGK5qfMX3gRgc6qg5V+Nrc2j9DFSod5Psfd1v9/gONuY/Qni6OW/DjPZGObhXu/JgbGYi
jxli4uC+ACISaBeDvvpeqButbzQFOMmjBB3gunCWf9xb/myCZpdBCwaDZgjyLkLzk8943yiOh8ca
KL8chvZb1cFGQA6AaeAuGozTHtucyp1nV4IyY/nL9NBlEb4XJP3nA2BEZhTd49RGQeuuZcQYqVgZ
JThd7si63+tRFa/ff6XRIYsQkExulJsp/aquEmq/SUec0n6+Gy2MVsCntGgYwQQ0QpMaiqM6QIJc
t1ZoFmPDNfWn4j0HJuzunFY/IlC6V94HcHqxh/RJHVQuUfpUiFYpV6btJdTip35rOPBVb74MLQAn
om7aM0ju14tg80TGCq3SkIhtcZiDMV0mdrULsQa23eocYn3QE6V4R3QbHaBgy9M5saz6SwNE4wfd
HmOhjhQiKI2hr2pTrKdcp5EjmYZtiRaod/mmCzZd7Vr0G+D5G5aSdxXjNQLcrYivyxe+Atxd9mhp
Fj10OgEYgadQWegNxtc6kb+oXFPcdWSIgOZAH+ZY22hN15w+BicMx5i8NvPbIcz15z+0ee6nciEF
Cowt5YMMBfhuY9Vjjejl5ldcuXgTO93DWMMle29yyy1WEzTqssZOMHJY8oljdsX5KbEE3H8HV9Oc
rZl29vLsef+gguuZ4Pe4wQvowLWPnBJvCn/k9Ugo+J+XS3R8nD2QGnMM8oYZTtiruKFaw0hin2XA
pe/CFgF14uzWVjrmvob8553R5c49t0K//WzbtJ3jqIQ3G/VENNpvt7omzS1ih7LKWssPSxqcA+3z
9yMNunYnjCBRTp24RppBBAkrIZNffERugToh/9PGO5g3dpO69kMdUB/nXFbLMIhQuATDa+qD6joy
IKPijPdEWDIaDcdukBwOSIk12cnhSnWCiEjL4Hy6Ihwc/o2Wrp6NCGYvrKYo8bGjf0yz9g8dd4HA
SfXA/SxkyIR6FF29sz4otLb1Dk97L54rvveqnTmUCFsuFoc+NzqsbdaHuaOgru4VP3XhhYQ80A7V
jD+QA/F5hTMLZMpNAH9vxQp7G+0LfncEwgt9IVAF/x0Pj0ZKKmHjFAcuQcVkIxvdLJbbDyoiW2Nj
Q0L+jIBUfVu4dmEyK6BAasdMmvdTttEL7/ehZSetWvtorwaQaBjEylOrb0fI5gsQs8jh5bXDE+Qc
0ewjSPOo0/LP9C7s4EK7cx9U1kuA2t1u7ZRmEaQ0MdArBKgiLA3UZvvJtA+0UBaths9dhsZPlw0i
1zMCFkdEaDifegz/XbC3RKV42JSepbHadVRiFEYs+Ww89DVTvlP3azs8CWDiuBZ08d2lg7ghSzpH
6+xcPpch81sv9BsvhwuyooXw6yPrIRPmFOdgR/XWWcwtpYjpGXJsP/njsz4cPf9RZBmInm5hrGd8
6uP4ptXEU6JGkU7m8bw9G6tI7FcEIA4WgE6fCHWpTUB5Bd5xS8EXw8kQgrz5tCDO40JD43Bm4G8k
K6xactgR/TlRD8mYQd6QqMCniIbyyJ701Q0e/Fus0++7+CeRIZfZLfTwlpQkLTnQOsHLnjuds/JM
cSVUiTqwUMWplEadqT5nZiTVeebq0WiaPzv7CtKHYEhxlsXzE3Hou8MbksZRkD9UH61RNXiX+OeH
tUs5b01XNPeEqiqvE80duwu/+PAVc/EGdayzgGxxF2UVPz2BBuFRYuHjUEiRxXs4ryEvDF0fxuyR
39sU4gmHm2OkxjREc/FU/D5nAtQtgebrWvxIlJww1PU89f4pufsSOsd9LfUOrB4B8vJQnEmimdKA
ddKnUWoxWvs1WTn8ME6JzOi6qve+gop8wiPldbopyn17dKTI81WL6SzbPnWfNZoBfzidqxQRGHnP
chrbXQ1OmnCSaNxBNqZgJ7756UcEnM4bKVm8Fe5kH8AOtVIiQc7DbKYY7Bdm4sQllhcFjWyPVJca
u9kjjLxxR2lapTeuh5GgqJxGPJeor9/nPU/3BNJDe91YxSw7zlbu9KskyXttglcndVpLPg6q2iDg
1VPfTyY5VMxYB8O6OeCW6iFIJMc/+nQVl64/XKIdEpdrH/0w2az3QJifSv0yRzKlq7gqLIj4XH9G
32+IXz4ENqv5RwG1sR9VNEMPGWSBmWlq2mPp2RXf/F76c7FyP556R3+pzTP3JIeQhgQeI9fRryUd
UJlFPT868p/svNhB4PST0THheCDuRP+Qz0K0Djcy4pAvJ22beg6O3lumZafLsrYdXn+xtjIHFBSQ
4NB1o1oSmMzDB2w7GSFy/GUJ5bBP14ztOaf5JsEVNgg3Phq4oEskl+w546wdMiuxJ71NnaK9lJLk
H+khVlRpy+SIWHyCK+9J5LxGHANlSiR7mvovXnVMoeIGP1iry4OvnQJyWuaKAttJbpr6uQC39Bu4
Dugf8eVu55vmkNqjZQExgFZZ+P0Hxuo1FqT7solnWd3OXIAmKPGHD4bVxVnyAGJJwxNE9/BGp+tG
896VEVtxTD/LDGUuf8f+M6xF5Mo1jfQvVfmb9L2HzekYxz+q+UjxTUhYi9TtCXBw4YUM4OonrwEX
41NDK92SfhMp59ZbS4du0UhnzAJrMKYgwRvjYReJBaPrHX8mE1DI1cNeWxKI7wYai309tXup+GmQ
OXV3nXmhUmpBSZr69INFrNdVh4lQXqjxY/aGZZq6LUxQJkkOTtoE86VNqPMUbtOcO3LWZNeoWlyG
9K6V3yd+r6K7VcuwiTUyNSNP0cNFr4M54X0yVsXkw1UMge9vjlZTbrs+Js4FbUYA3Xfr0pqt6tmO
2GK7IhoqOG59sh0adZgD+aTun671B5OoCCavg0z5g47ykS5pHUi9Pn9ebOWb6eWFX9msHMYUPni5
LX9GXPZtdPfrA8y6lZ113HOMMi1pUuS94nkoR8scdEi8f2C8plDEiEOE+R+g+QkPvp4lIwcrNkhg
IRHYEwI2jRwWi5nerXenpq5nY1ZyUc8yxBvfMIL4j1xfs3TjkTndgyGK05f+K4PMXqsEDTHRfefB
QrWG27B+QoCTUby4VkAPlwemtHmZ27tEFsvW9WTfbiTb1AhCDWwJ3yvmN58eA5ceY+ORtTJfQXQV
vLzPdj4I7R8Dlvt2k3/L2QgG5f5PnwX/s7QeHs+14/4hqrjNJRfTMaQz2nVAYI95JF0Rnv7WOw3U
VgJOMjZYY2q/eQOycNNaygEwIv0nl+c0GzUnVTfg9do1Y/seUEnpU/YlARCEARnHa7vf4R/n9iiD
/iFUfUcr9BppBgsXnkfpd1EGshagwuLD/oFrUBoGF4cvHkyT0n2Sg/YyDPAQGklgZU0BRmJupl2l
kOsNjBgsaDr9yjEJYHMUd8MRfVkSvlK+qmGm3CmR1KKHvGdErWHB0fVMK1fi7O4VxwJv99h1zlOc
qkwkL6mMYIqG5FX3kvZwkm6HpLLNlm1h4s2DgQVbBOmp9bGPVNXnIdErVOeKAXUeRA8JnERtSACV
//dAf56dSyjVtGsw+mGROfP6ca3wSq3Bmv+tQN5LVuQQUADzQrSzsbbZvI7cgTCMBOiwpWn1QHPZ
/F+KZUl7I51gFkF0PEd2YUGkwMJLwCexxvyYpRtLlUTP2P6TTa4zMBW2jPHTyteg67ruixhum0M/
p/T8Dp2fhbEZs483Y0ZgJPK76mgmtr6SDXUiWqVxVFuc2tdwjchHCc3WralerC0s/wsOIzZkOITN
xqb5WnWeCsmWM5Jm0Qg9Qj6V9BSVpBet9ws6cF9blQYGTrGIBhw6oQnqT/6PDr0dzRcU0YLCwF6K
kUZBorJkZ7yFfz+QTGjeGeN04p9oCrBtZH0vsYVGtCJ4W/gylg8dJqepdYE06rKNUdkgpldFpdqx
AjaLH8EmFx/mdw7cKgqQo5nPhVunvPNb7dGtH+v7iLDnH8kfmgzJr3m9CL3D92/lw4Nk7FSxzaM0
UihuzH+LhA3wS5e7TOqb9ezsoKklG8O1RqCcrYzm0CEoeySsAteW7BFDoGeZv9N6sU2rkYZ6d89f
QF3NocWCTU6O/ccyhU7ErbFOi58Pmr03Wx4DlEE/a9cDD7TOTJaAu2IuEy72AjJTebQB2nNqhNb9
045blgAlDwQXLF+N31Do5Rz5Hxtnw5CGMQZvFNGOhuC6o+ZyWDfrE0w+CJ/cM015Ptdy3oZOaV1c
LvGzI3gwQMQebn6UPvTPrQFmSdSdmNPMy9ahbRYIycJpFTfTu/CWq/mbd8CVLmo097Lo8BQ62n3A
Xs2iBsqQ0BQB7yeeVuH+eXjG4PDzP69ely9H1jevUFKr27S0vjv9Mexype4dEvZtYhuWqFWlpsxL
ppZEofHAERoMyLm+2N31uQuw/bspbUlqq0FRaqxmWrKTweY4RIjxDZ7kg9CLqxdKhUvFm9IrPKFc
VLkBbCGw9+qCkS8KIt8wu/jwdjOAF/4m2qi8NdOi6OfzCiHm9FwU3bVANLWoP+wBAwmpy8ofk/MI
RujKJ/QuFgTO2Nf+JAKd5MEG33rZe+3u91NVz88XXQTEDxPjnlkgp1YpZDM5tTXQIsjDn2UZOkFP
uMdci0DZe8fkd0RdYtpAPNFNu07IRylAdGOE7wQbIvx+AaAplAKaH0bp8O2XwJP06ga0A232zx/m
DOLUKzHnaOMXkEzIYjFDX9Un5EpJuuWVM80dn//leXBWoyvnDJfDGLi7j/JJKeYZnXV2Ibm8VZOc
Dzgf4w4kEB6JkRYhACEgBxj281jaF70FnV3v8h2akmqysoynbUXDZfDC9y4MYZpiTuUcWbINYc0p
CaAG7aVfNKDPHwgj3mTN6Tml9ALB10d8vbnWJ4dmZCX0Xay15CrfCIKWo7joq7h5MfUXa0EKM1xA
CNQZ1HElG3IQt2bluEvkn0CXbyTAZsBGAM+PLut24t+hChqEiUQs+RFSwdDKAjGQIGYAwqJG5I8/
NZk1B60GXKbVTmAD5lkGS9D0sFX1tUOzV3l4uKrl7Q84BNTDHe1wjLZAV4Ed79b1aOdnzLoi9C2s
PNS2AKCztCVNjR1rgWHKDItaUPrxwpHVsjwMy79W/I8W1aECA8c1GAjjCQmDTjt/L5ukDk5ZV5ou
mc+4+YBytceAx7t08aKjkzEHUFXrBJP3+OoO6Im/iw77ErBNq4LdhpgXS6K2oAoVGO/G7j95JNlO
MC5jEiJIR9JUxf8lbvaO3rg5Co6VD6adOHf+Mi2N4EJuT8dCkiesrsz4MEHp9W4TdZb5jiCR8ygc
yDPUhlUZxuH2j9jabC73vpehPKPkrjx/0BudNoHRPwDMCSt8EY9C/exRK1TGIvnuaUgEfq+wXfhz
0RDGxIrvsW2KXwmfuETYP202Be4Tedw834qxB/mGqjGtYQcqezzhMJcj9scjz0LHAGZvPfwjZfqd
tFvwxEW8oaPpJNEuB12550zRCPJeFIEouGUxpR7wpk55+hv6XCDY2Y+95vhPeMPQOgO7p3p4uZRq
ZlmBmQ1SV4OXTruaYo8PvmuMrIQuunjklDCbJ3rRX5jRWHERYIqtT26UwrwEplI+FvHKMm0PkDcF
Nr3Vwd2CZWBKNsqLoKMItdWV0cETwPHxrLtYSA8PsfeSLN2UWJrkHnRL/G9YITi8LTnVID3XpRn3
OJhLBzuKI6ckQoK5rwcQknfiqybQVbmuIo5dv3/YMzNPokR/cBX9zZ8nWmM1p9hfJBqHmYbIMUC3
1KhUHQbJTla8K8MypbiqTUC4HUWkW5HhE2Z6lzNq3KlVqT6rkScuvEZUXWTnIgrrN6S+o8fsT5nU
PpF4uI+1enxgS3QEDYPPp/UxnxqVzGF2r7oij8NaLtLGPwjTY6EeqT1PJUJ0ZKbEPHNuU2PfkQHS
f/DQ3zjUVDsF0L8Uh6ZsIZqkMT94Y/1fy0Pb5WxakaC7aM5mRWwMKRprtxcSv1ERv8NhHENMaQLv
w7a7zJCPCmBN7tq4DVN3MesmGLgyexIDKt+8a4gIgJ2zI0dh4Q3DzMdoewWNjPjEMDfzgIuhDpIb
q5BYlfMyZ+CT/Ex8ZlQFTxKPNn/l/6sxx6YWHhqP9fDHAZidJMgzh3zEjeWZPZSaf8MFqN7CzJyi
oOCUtO4Jdi3gCQURkeFA1+Rkgc+04OxAzGHPbq5xVYexrX9g3YiGD1NrMWN/FuuvnaxRFo6Wr2lf
XDtPppnUxn/N+sApD50zCSZe2NGg9gxo/h4JI7rusBrKp4ZfI/CR/36neKvlhB5Koo0OYB8aJPrk
GcIuat4YewS+JIpI4Puzb51+xGSsdrO2GL7DViiRMvTg81rivUZL2EEkLX3TMma5leH+g0JeExVD
2FcAYsyt4He2yNnyn1L3QbgrKiGarxKKi58kX1aWhmLlX2yS6SwiD1Q+469APJL7dB+Ol5J6CJhE
yrLbguiHwr0ASqVv/YSaGr+OQr4yyOdERC6ZAbtTosoQYNQ2IZyHb3i7YjhWERW7WLCkCC7QR1uv
4nF6BJfpvDSEq7nhCWngjYQu3ZizxJoH0R+csPiZC1n3LdA/YQzt56KdhGcGIzUWClTFjocgEKNk
1zQgEPpwN2H3xATW+CUBeSU6UOarPq2xKQY3KaPHCzHXW1Nq7ZwBy90DTIy4wdpm8y73fq1x9fnL
nnpYsF17q7LfVyQK/2z6hULMaH4S1lCABD1+bUWVt23CuXoq8Q9/OwGNvGSU98NsltNAtA8wguiT
I2qaCojFpED9V2YmEtECOQp6qxbW2RB85CCyAFiis7JPm0Gh1nlw7zkgB2WCoJgrAjbvxv4rgHQp
EjGQwdXWmWdqJorldmjDZ2XbgYfz2QL1dGOzOkjRyJnM10FEjnbLzZmgf+RV+/DSBwV53EkYzYmW
CZvmXa5DC7KIvSfPGzytip1CdgTOWfHRfv9ZfH6188CLaj3gU02x1PJ+2OSPrypqIMUzTJrzd+pS
R3OIWrm+cSh8O82Lzafdexe2If9nhmp54EBeFLWfF9IuCH+0OzjcHdJ6c67PSgcQ8zh+s8He88Sh
VPnY0f2HpSMeBly4ukr+Tssu127FBLxl3jQwvLbl55IUKdfNe/6SbUaVALMB4YjT2tAZJ78a7vbJ
9/DiImxm5LYhAtoTlsT7MBKZKNGipmN0bmexRjLVhK5nl/MpD9oSy+yI551q20mLm5CZXrsqnZeP
g+WK9MbRpe+rVGyjr6AOVMfVnGCmBSVXuzQOn5cdPRXQh536A+iIxCu/dpwYU3QKrPVLrKoW804w
GBY2charGPlvA4wTJO7PR0mGap1wVfFeC3Q8OdLP0N+SgyyZTQJhB8DYLBT1v2HrHQUAHUpEsqyt
X1wzgb8ba8pjAzz3M/a/CuD6qT50R8eVDI651mp1l5c+VIY4J/VIL4S/ZjohOtbnIXjSyMQEBOrK
L1oSq6O9ODGT/flwF1twiKKDqhzbVZad6fELHk2g503jO0mRkauDO52bhBTDhYa28FY+gGtifIGX
2CakzOyI/Ryu5LxFm5dExDm5zNUBQ+GyJ23ltmnVdSVocbmJ8/Ud5aTfXGbiHY0MS56tjh9RB864
1IHhk96IcG4QeSzngVrYmHlw/4nfpqmRoLUfhOpN8c8DacW+aGLN6baTsiNmMmel3jq21TIbnMYb
gQfeH7lBEgjAkMesYMc6+sjF8cboMeVd3mC5ZpZlpqhzaHvThsLDAgW/yAcPq+ho5jbawIGEQjw2
MEEJqkmWvir0K9Y/nkKLw7I6v53f18Njz4KoEggYTjNnr8BNJI4fmAzTnQZ1m/A7Bls0OZkFgO3v
2b/SAfJVa15AmqxCxNTI36mac9TDqJ1fk26bax+FGbGPLimcXp3m0oxoK/M9LwVO8jvJuK9PiG1d
SChJaTZ0V6dGey7mekekgx1HCIDPx/tPhkbPA9uRyiyzg0BjdnJp84PWD3AYdQ+V2oFrxnRunQuG
gpq62mQDZNB/69IGFAkwRW/2e7C67hgI+mVNGierpjwnwiHidBu2LoCYY5n1oQ0KuNXlQnFG942F
xy4aww/3gGIvFQW3jewXRZcpJQsbQrpuJb3u81CsQ0t2/u7bMmpxSdzGcRuDBZjPRowkgTlsE4kW
MWMC1UUQVjdjck9BkbsVkydgWZ/SD3thOpAFB8U+n6a490icjypKjrJsxgOBiJG4OuuJL+k9ULmE
B6nur4UA+/WEF+ckCoAToIrMb0G3ZXtuk8m+4mwmdaqgTucHnJGc9mtI047u51IdeXPAih7EYcZp
v5c23g2F5NwDu7IurMe4qsZC8LTWmucdQ89wi2AiRQ2yR+H1IlPuQw7jr03oM/dIF+53VLOD2/fT
YBinZOKEJlADdNQQir3kf0g0CPNj8Q1L8HtJitHJF4pZCBib9hWi62oiqlh9xGKhhSLwJdDy2/al
6n/1XMV35VMl8askm7c0gPqDsm7u3hlPf5P5CYq4IJuipkzz0CR6SEH1r8YQgIxxvEYdAyf4vui6
5ORBU09uChZt4b42v4ZqaEfrSnV7ICC+ugPzK200abELhS7aBbWPxZgkE9s6re6t1jp3pb8pN1l9
9YNeEKd1PJiJKdSRnOI7bBLZZGHjt4+puQKN9FNNVM1aYBBJbIExnblskhUovGy7p7AoMyVgMxX0
QLloEH9Vi+thwwKZz5R308TOpmFj/1kw8AJSooyReOiA6+yLNwD7ExDS6suxvBqU9qCKiHCzxzwC
qAuFx/Qn+GG548eyTzTejUX2TSeZABZjKdLJfFTeTlPbjO8W5O6JXzBOwnmgOhxyGIOrMxs0/HoA
Jb9idCIncfZu2rSXDesATv/tqlZLldTRtO1YkBtkJ9gsdQ+Q4WBKQ5y4a0DXPxYkNtHNA6Yy0YLR
qXaw/tVBLtvXvvL2uEzsZPzHsapIuURD28LyWTZH6PlujTIizcLrHQG918lq2fgov5kkrfY7/irk
RkKu1EY8TEilYYCH6LleKaSK6O/mQPVlm1ixEh+YhzhPI/FbdQbvTnN96Aifqh5R+xIE5jzptmiW
AKDBwll0IvKfa0yBquY7HazUqe0Vu7YcdvSesIwATKVJ+69RDvlgDtV0yszyb20/iky6vPkDk14f
M83/xYBP1dVJJ9NkTAtcYkb5DaF9hAJJx1F+94hSuluFX8z1FjOWr0p2hta+1d0j9DYHLBmvbUs2
5mKJz+qupbNP/QgCH0rdEetwWtjPaOlgElTwTKQVhXuHxgrFI40+juat0nPDOg/wk5nw0BboDfyU
bjg0UErMhQP1Aecf8YBVZCRWH+VY3RDdWt6zPggG25t0VE2xKhE5zloPV/7dDuBue266sA1rQ46f
v28p8EcpXknE+z3M1zp/eqbRl8FuxI2pEYRzHcXYHKW0jY1C+pggqVXxLFxoaNm96hqvBktTiVIU
IDHWT9wp5Fv+PAVyymv0I/VV17gTviWheUSsPXxSgdMbfp4sRFhSb5TYig66knycv/UqW62e1Y6g
U8y33ezTzrgPAcYEJx5UPHSYnA3VXGXkqkMi0UQurh+NET/KXXykmwXBmq/BIDx1oL44LwtKLiO2
xHeXsdAGah8zDd/A+x8TCAkXSWedVyUOSwzvJO+J9Zox4ofkHDOzhmol0bF4TZ/aiEbM7oUTouUn
po6Izf6YSGFy/whpBa0yszj5iF/4tpSdDPDiTIdeYr2XcqsmggV96G4cbtyWIkgbQqJCPNoSWq0z
9t6oB5N+omOIXxUWag9C2etWgbn26yQeL3g6iZQxBqoejEx0SGAWbjR0Ptz6L5WvJz0fPYAVb8PM
o1Vs5d9s7mpb5HjRX3YezSdbXHWOPhUolGrjktcOjl/YkpeC3CuzZeMqg03fS8LOZquA4uM7SPrH
NYhVoX3n0A7Nn3G04aQD2xthG+ieWQepNFkH6RZaeVXzI/KXGO482qbewiwI4kD3GD8VAzg2zllg
caV34qQIO/csADcPNP0OVtJgP5QICN+5cCeODWCLCAY802NhKjfm38wCiv3i3RiHgTjGgBZ4OsJ2
h2VILtmPjMnon43awvNR2A5/ayDQfjqq9D/d6m7rWS7dDqAPZ+4Gl1yy2vK3Ew+tFOqzdA24CtW1
o79F3VLfZeU6q1kO069i6jK+rrB5PaJClr2MXpoVEVy0kNfuCmELhxR93YixTNGr7Xwv75hBEnbZ
wtvI7zG4xZOhqXigShErpKbArtb6xVRIX9OEAtsMs1bSe00IwPNLuX+WpZtIsT9hPqCT2rdSwlHd
kpO6G71ozyRvO/hR1Eib4goh1PzgKMiRq9OZoF6oBre5Anda4U6izJeky6AbSe5HRWoeiiDmJ4sb
NjS35GlYwubxHBA4k1jOv49RakBZLsh0RQkBpbiFdIa6wh8Y80KUGG+00TWdaaXuo83wnvopgNqM
d3YVhphau6lq7gR/Cd33StXepRVrtB9xKwrX5EEgNyHABlAYPhhdTzWAgRrLD4inynHT7/7e7S5x
/qh0r/r/oRduCj6ixYi9SO14XUx18Pyu3IpO1b+HFmWw4jfBtDk1ZGyy74fnNouKk4RyJZO3eznS
c02BWC0FOyZRTrsTJfqUB9L8+1hnmnmsIuoWdQwkZG+SugRyP24t8EDajtW2gU2wP3y2xVhyV8CC
mrzYRG9NXiEZeXc9/fXEQqkurRaGbxhb/H1WiFUE9dyf+QDO5fOk0vqDcDwnPUITo8jDTDRiHwzi
TXQEpYAa0minXAyDd9bUMnaIg1liQZOUuLMxTkcsiikpM93IELiObZBD23KDVomJHDWzabJIJm52
dJb9oNzFfJtyll0W88d9w2J9mJLEB4zlshjjbt0GwiIyNGdFcdWmlOoXr2ir3s7RoF5i7teXUy+t
2cxkNiusZl/Btced3iEM4MzMXpy84+jla+Q1gSzmgDp98lyJ8nOVbggsk7acdulNpdSDThMI7B5+
QyqinqQHrDawqzpYBAUPMDf3AutRQVJL6fHUB+HLxsTRwaiD2Eb5RsQANR/B8Tix24KQKAK3cZn4
WeCEa31xrhJUNsajBEPErAF4krrAVlHHW0Oa+qr7amqf//hUuO97fOsQkGvwbQQ59MGQihghEKFU
gbhChyevLerAhr08onqti7FCZa7p/iK+VJMe/jQvE2Q7CX3hwei2Rx6AEGJDPLII9m19uqQHW+bp
BIJUO1s4akpv7L3L1q6KRXOyX1VASHsqc2oU4/g1S+huWemztNqBTi1NEjg7YMOD9MOarOrSa5GC
KXqo79/hua/5gBh2izD1zUOZxzSRC1WRfraPcFI6HnIXCPKKGdFTP478N2lon4yR2RI2gmkSgBA/
0Y3GTgQSDuTYC0mTugtCT/m/t1tOdi7Vz9AsrVNmi1QckjDv0s4kVJpKm+bhKynWIjpZ3nFW3mMR
nCYIcqm1PJiYKNkCYP5M2qnMB9lyuKb/X6fw8VLrQwjDy5AqFXj7fSrep9XJURXvpvjvN8SWeX+e
7IIb3tp6SNE8QfIaMyWtEnMLGzKs00EmzY911ZNml9875+Jmu9zKsvPeQgFA5F/5q8J1I+lMh/bw
ZtckJO8gmDP7/hS4iyouR4Woq6YjHNhAst2WpCKmz47Ar1U46Tlk3+fdoj9t4n4vOS6hGd19iaAh
oxmEx6SdOfplR6JYmyafdoX28rPg5wXDOxVK77iZlUZoG3B8EYdLFK4De8G0KwpLZ5aR8LTkqPY0
54Y6zu88du99AzIV6uZPsScalHAkYM4PBZ7HywUevSl77RtScYr8a/j+M/PDCJZbBbHN838eIdwJ
AlDk1xZKM7zi4TA2HoTT84e4mMKrrUISqXr7oGuZwRVYpGZTz+YEFgme+TjsuqM1coo23Apx4Pxa
b2X6Szb8c1NZs/pgKwwzHYF24bU0PevlavvFEc7Spc6FZted3QQvQCDmV0ubcxMisIAWcP5sH01H
XGxcU+tCwfCvld9zcpwqTAgGWg+bJMCJY4x/pV+RSRK1PkZPnotkRsYNm99ODIxGU0AnVgQMKB83
xZBMXZXwZgQs7ITiEkfaJrfzRTP8hVpGYz6Curv5Qe3heKnvqSeOLkiFCd3tovApBbufVAzMnELS
Dd83zl24dpRLfWGxkKANxOtj7Q4Cjl11FsU5JbYvRQ5aJPdc5+sniLtQl/FsdMtrQxQSVyBRyiqj
HPzZ3LOw8sJhokYl0TmsKCmbpu4tLI94kpVaC/6FcikZE9Wbh2GqfiGN4+37T59QJZTqi/JhVzEI
8PNkBat7qkFOoNqaocyDvgPfL1hvBLn1uIMtxHgzfVGJf6G0//rVhhucRhZ0CIqy8nZmZ55lH1Mw
XhnbRLH/DsdIEASItNRs+55fgd46ZDHxKKrsP8zua9yZ0R2BbDuFzVv0mZFRcksxipLgAx3rZpcd
YqMUqJPmWeGIlyFe86IRowrLZ5bWUbHDmOksmnn3ZX5GHyvZJ0S2huPy7ezhZB/5pApDcDAk3UjO
tlRvr3mnfvwF8iF8m6/cTKraIP/fQHnkMDMgrD9PB4kUfmp8QK1jcbLzkH6VSbIu51yHtBKr2DAh
BtBRrURd4vAN9zfP5gJh44ABKhyOy/eURGaaqiWxEefSxzZ+46JduduKKuE8S/C7MSeyGxc9Ag0g
O3lHtYSv8O9dzy3dTvgeynCisX6wGPr9DcdcE4Nqa0aP2qahBd0b6KdqKmMGDfQ39sJoxIblGs9t
DgrJ1n6bDdSEPUxicTLQpy190JgUb8CJzvT/gEoygr6i1AWX66tNUmk3qiOAY/ub2278M1WOQKsc
UdNKGXBRcrWpB86reUr6ahGQrL+ENPmoPReuT78SKMfrhFvEvFUZwuQA4L6u1miegZeJXi+SV/k9
gCpziyW88JOgTqK/wu4I6EMs8b8yMaCUueT+piNFuvR6eMpTCXnZ+cdDzKNuugCX1hQiqQAvMCjk
VKb2Fpq0mogjalefdwZOxYf1L2YmcfAs09YclNoWCUk6NJhviT43sm0JlxAeJVNFIz+iVYFMb8CP
wu+pWd8UB6ilzE5fa0jStWNNnUsndzdE82QMlkDud/XW+nFt9VYPATVdiJzilG8nS3qAlSZxkUfP
zH0+f8GyZpl341EYrtJTw12jqh2Mp5y2Uc3fwEq3Z09SGZit0wCEwDQw+cwpzyTJbDCBI2AHTIvV
DIj8/14X5wAmxzP5ZmY/ATQ9ke3fTz/0ma/IIEhuypxH4/CU9M0d0+pPZFx68ZFbFa1INz/XIEcu
unJ5++f6DeXl57+BU0XvPdNWEwp91xrTaoitReWuWiLnTyjQsLbux3VI7G7XcowXq0DXq2GuSjSP
nry2ZibVVF056jBqaPu7/6lO8kX4LY3dGuHWFvYw20B4PvuqaywvRRr9V6Uve+prxO3nY3a88h20
6jwogbn9LO1vJNHAHOmDgFGzma4GIIJimTur+VPjccDA7PFOb6fht8T1yfkckJ2P6d+ehhwms0nG
4OLEnzy0AmXdsun5Tn7XAgG0yGYYGWE/o/s3vRGK1HHx6rkdx++1JpTThSOsjIki+Ysq9D5CTCns
J1XwKCusKg/0y4NvzAkxiy9r0jJmqlNtij+NziVSXVXd3G2EcTVkI9is9J7kL624v0knqc6UJsLw
2rD50tC3wAjS1xeveCcjyIFNeic4+N6p/Bpfz72Eia65MyGdt4fu9cxBmlR3CWiiypmNKRoujq9O
NWAHIc6rIc3fmy59K91inxF4PzjbUeXrlXPv7byMJI1RVu4Ts5FPZr/D5zZreCxSjXRmk0NvyaMO
EfJrD7y/ctNfOQy8HX1aQLw4dPFsBdRa7VUCjsmG1xPy/e2+QOhTrH3eO+u4y55J7+PT22yp3eOX
Z0SkJRJiRJvKtt0G1jRAxof6cT22fbRWsXag79EfN868O2QB5wGGCtt65qZodwCK8DF+9DUlMIVY
kxfdCyceETmpl/NN6dFKhnpMCq6fHDe+dXbWyPFLlt4PEVTiap7ZxIZFLirh2b5n3MBmDhzLr6j5
sZOIJ/eG92xP4jF5yGDapOhsanqdKO2KI5t/D0Z3yHCuKZwHXk7j/WAaIiomvqtJ8nWC9IPNcb+y
G9gBVUuN5o64y4aP8olauh6M2WesznkqvMv3Gtthi6iwkXNCFVcmUODyp9KUe54Igq65G3p+wa6Y
QwUj0xjSRx3w/itSXznJSsA84WuK/6j8kSWTvagDZ+lx0nqe9nXu+4czcxQVb1h+wmUSC0ZfNq31
VIoAW3M+RYETwBgnwM2zsBJdSsmhoRmVgzgYryFU4kVZPkaL3UcFs/qWT2ySWR/znyX9wChAc46B
vWJhlmIXXr16m9Bc0NrFP8iwcZ3/gnc09TSg4hzo4x+uA61uwNdTzyuu1mjwwa/ricg+qVBeszkh
U02jbnGRB8zwSQIdvZxz2Xn3IxpLXXoVti8yQL1M1AR8DNFHv0Qnh/aW0v/xqWjs1vojyaiBQoAO
uGP7ID/27T9+cu5w+0dQW8LX6FvSmkN++GLw0WmcRN97MxCWc5YzMF+V5DY6Vy1N/t9VdtQijK77
Q7y6CUJS/Y3oF0MYskyU8rhoJ6ufN4b3nyPenWV2gaIMPErAiY3FSPVpQd0vkZN2Xalhssp77tut
J95TSQjltNvn3n2OjsENGRt5dNpUOk8GE2ipFtKYzp6iQc7eD08IRfjFgdGnPSIFYQEaYGun7ueX
bdRdJyd2LVszqCpM2xSrcpTCuYqbPWlH/lQAMgTCzYx1G2K6eoB0XY7Cx52hRBSresyXuvp9hOHm
hNzbbvS2qE2qjUZ8O4Rg7vypi8rGcT9OrY1eGqL5y/K1mNI2Wq4HgVgxxO1sb3rcGzHPz+DZcCuU
MizYbBTNMOjy2zwUighykM8epjlQ0miwmLycQ/4ncqYi/42mBKQr2JUbZxkFvtyMh4htou/mWMdZ
z3NfzAX6oYtoa6twFsCbVOGHhOuXklJSAmAsfRUC6P4Vv66RBAQ8V6g4/af2P1g2sgJbq9IG158S
N6lQsNqg+BIjIniGmHxatdygo5SoJzExyRrAq7TGS37eVpebCihz+PD5zSrH79rXzeMDDgjsEUy/
EdrlQ3IBkeXz0IYs4DoqIkiaZRsd7kTnSO+lqWc/We3LGn/VXK/A13lNS+Zg/ZmQaJuSIvhBeyCv
1MUoleSJbhFH5XjxLZH8/lwZNetXHD8QG/VRA2JmdH4R5NeZLUD7xL76MWAcE/dqyZrgTB4IiK7/
g1BApe9SeJXmu0wyOsONZlGpbx7N9joXV4yJWOkn2a9zsSheD78MZOhWbJBuBNSiThbIOXUaq+1X
DBi6GjzxBs5nzzmqOfgpAemgkMKS5AJ3bUXCtUFMo+Y7zkDgkfPceToKSxD9lvbc2p+Y0z5a6HK1
J5xjusHCJo5fLimOBX3v1Dg8DMax0OO7tk2hXGlBHOpys4djVS3ESM2ohrQuMqrr+QMMvNALPswQ
5AEGXC1ZSODzV9qRwhv7XDsUqu4yQnF0Ygju9a3CMw4lMSYQWyFrSRKZUT/wDkvl23PWAbCL4dhW
sXE8cscfRS28Rk0Eo/6h1ighXFNkPzI5gC7QUCTW2yAStrttbyGNmlJdd/FBVGsiZqWoqo9bVm3a
weQx6ymU4e77fge0YvsOEQgm02UqZ3d564yh2wde3vHnrHe1PhkhQAmkF17njIWQ7epFJkep/Ztw
Sl1IUrifHE5LQXPjmOSa9yg1guIPYI9v0yr0PA10PZ3ajYLqoY5R82J8m6/ExMGnqSmRLNOoW9NN
r/cnC65NuTDOu12yxd8Te1G8ghCS75JejI/XNO1dQHCEqhumKcKS8qwhFzZqucCWApbnl5q24wdS
4nyR27TbkVCZK5vPjpolzIfG8ClJHkiSrGdu75+NxvM7/3UywIg64O14qGBAI6Y6t7yDi/WXpORs
g1+CyP6d9+InwYRW2pcawb+SFuWjFDOri2fGAPb8lICoKg5pGTpfyHcMSkGIn+zVEE6deVP8ppYJ
czJReSRHCXfgPbSNml4+f/0ADPu4B5EIwXcLOBhtuM0aZwcGhjlq1zUDyeEGvXcSDfLT4IFy7MJ0
Q/bApUPCwadQCHT30322cK9DmMQ/PWnAoNKAol+o7nwYezr33GcKO0u2gOFAGP1E7YYQTkwTiDvg
tRRiRuXxzI5iYkojXzyLMZR2EvsRCQu7N9ILxDid36K4sXNqx6UDtHAYB1U3vAylc8KUHzfmi2L1
zhI98OTsSYYcfSvP9EYiUL9zvKAfzpuvLAPp60ryAUwGMxXzR5CpRCdj6bJnge957QTXNf6s/ont
Yc1tPhHaHh1XN/EBiGD6Kr5Tsy2iVPwZbKEsjwzEyYfPPaBPvhHGlvI1uykD/iTbvE+Va4V2KM2F
894mduwYMeLcQ7ihIRu8rbFELFkZ+eWWCOt3CoWNTEtho4mJo+m91vNzC+/f9bkafBP1JPOjjVji
bvtMqNSvYozo/o3vYFsy2FUu23eKP1KnU5ZNc/csp6YmfuNFKhBxB56H3ueXC5dBfjkGLPuHOk1O
DMM978VDkb5475TWgOwRBtpNEEvnFUr7mhJFsU6kVpViPWx1NyiWfVLW3MooL8cR7DktrR/yelRz
sv73dJQH7QUq1Od0rn0lJxDmSC3mIUimGFgj9kl214v3h3CU9DFMK6Hqd+Hwl2/+yols/wGKzglD
iIdaKZikv6NX3kFHEBJ3c6n3AHej4bNrlPFViXUUOv5LpM03irRLAkrkYO0zb0nexVySV1VgmobA
EmW+AIQYSYLAR3UHhJy3i2bOBVlWMoVM/Xtirw+Ui/9mlhRNmv/LL7QG4mR5ww33ETQoIBo7hQ43
ue1vMIQqzrSrlQ6yxvEcQf1Uox1CwZzz1BTopwkfOuqw2/A3dXQPm3xLzPzTFZeOOyfgJdiEmMmg
slBiuyl33UyTFsMja1erz2C7DpbdnqCBX6LeJs7w/+pSOMBAOq5MB/VFUxtTeLOz+91EyquSQqXS
A9fNOpD8TZ/Zp9tCwW09mtvVGsOe591vPk9xXRE1Z0rAkGfEefAmnYFWHRkm7ovR5dn/KvH7I2UK
nal/4eNBZclReXNVluRkE5hS/qf4eZKyHJJLA2C+JQHuXnyGwRTZ79CMyey552rUhKyQlbXct2gC
pHXbUXiAisUVfzwQdtV352q2ae617SNy4NkR5AKsg1s0i53iVMaGchglH9PZphyLR/dtyOD13lze
sAplVMCnazZ9IFt4jN3cVj5QvPxJBw7azinXibJcU2GhlTtL2pMBTzP2jKu3gSpiAA0d7VENn9ad
gQtf86KTDc+IW32tCxJgOEl/uW2mVl2Kvb8TqZBJ+jnrH5C6y03otvrcnkATw0jgBm+NZ+mUCJNH
UImBsXykf+il4npunAQ/CFgFNJWtqqOl5q+YsIWaW2iVprfAiZAeM0GDkqFtjPHxtiI00eNjx2Hr
VGPft1Mc1HrrDfZdBGH4rmuKCvycYAuJI5oz52zGX4F7wx6NVdDW+oDpQ7eXf315Hk9Mix2TQc8a
dfG4ONM7y8L80qS95+LKhtISzrYstYMFel89WMCsWBLzwb4eQinr8fwK455Mjp6Qsbpi5g8fZiBQ
tGdSmM+2fUTrdhaiRRqZMzLRBBEIKhIstsluvHJBj1TxeYBIRWjT88PjGzNfqfsUAHDdSTwFqEQH
I3FvtWrrmuA19FvwzM9NkTEDp+96WRZMnZS6ogn2KjXnV+zPHGPn/fxiS8WKDy3VJEnuABU02Wah
oCiRGTMjydPTJS0z/VsnUZoGSPK+cRjHQUfvE2wEhk+zdXGkEJzLp1L+Zy/FWTNMRi9pg789UtIq
CpMhoBlymjbcGah8hKCKzCAj90rQCPBLyNpmMoQEldvA8gHzOdo5fpfPdfFIANl+0A2CjnuHu3bK
K5loQCKrFQX9IA49dp6Lbqj2O2BC9oUlm0XWZVFJKYfcDzXRnF6TmP93HqMshHA2P5eW83/urJMZ
/vIlsbRpfzpLfGU1PfQNRthZORgrqnrH2gQOySCTwhLT7KZjSYzN44u/Bfi2jR0qdZOQlZh8HCns
/dP7pUikB+Y/yDz8KHJCrVVimLfzKC8joI/RD5djfxjhHa5Urd00HingtszrMg0M/qDEVkIyIyFq
fX5BRtA5XzkeADCJTlNwEEVmtKFYswX2AekbF49EfeBEhVTntCbu3sEhEu99qZfvaw4waSdy+dY4
QiKRAeFTDdWe21GWMnr6SaLkOPnmb2ixMKykbltvQ36vQ9xSkdFkOCPvGJD89PoAa4qMGI/cVv11
V3Gs1KhsF1WsE37HjHIRf3A684E2LVMtD/6YJs77HcOHrPMNiys2yHZ8za2RvYfyiJ8gnUmuGVvl
ikf2ZJL0mlh5HuZSOd3yqRb87f7so+oktromXRLNO7zLotOT6ct2Iu1KBpCj6tklFjFUp2nnAz4z
2voKXZN1Dcj4AvJC2TJOsnHq5LLDD5MZEFRMLdvjlxmea2VLza6M3vmQnTz1ioewxg2pSgDC8LfI
+VWF7MegHQ0JOdxSZRseFXvzehIV4ocLfRacAC3x/YA3jEkyINJUKFBn62CfZnVACo+/XPaPad7J
AVyAgbu30ns4BHje1cZgAzG23mQGaxTBItrQKIz4HPX5sh63+x5OXWC3bnj3vuG/MBqHZxvtG4dH
mMVbUZVRhTNb82b4KKyTGeKK+/y1sON0RORFOZi1ZqzsttFUlAuqjXq38QRMFqrUl8rj7MRmFuOZ
1lZqwxiQMfYDVNNrinxlm7cLxsN+jybb+B5peNbisPL9FfypnxCykP68qdSjeb2W97maWJtx4Ikl
xKEAeCoHXX6mssyXQbCzruKU+oNn9ZZyl4NiuOw3UjMd1KdqysOIn3HFD3gMnong4Brb64lw7ZQC
iij8PappwPr0cstQpp1YVBfqTKRRjYxnThZVKtmP7juZyALmsroFFgy+KPgx8G/0+82oXsczPRNK
r+ryPrmFtp1U/GwvCXXJiA3WzV9cTPGve98BsAZAKQq75kbi1cpcdnHUB+iI4duTdoCFclT7yLnh
ZniStehSkMBGwxyIMYcGMRmBofRF3gEH6EeT1AR08cF9CE0D0rIb//VIdBjr3lP5gLdufNh3QeW5
QDK3tH9OOCITOcDxoKRdxiqih0QL0q55WXW5XiAnz9Xvb0jNhCTQvE73an/FI2Pek13/PloOkLLi
+y9QJQD489Rf9LShy9frzpS+gQ9WR08mRksAAuY06WZgPgUFRfrV/hsjspBuXh5ieHp0FAnJ3E3O
QDmoEX3ANabKdZdPvvAXEpSUnZLqLQy9BKDGlh2/G0VFcR4UolgWSUxKDjqp/XGWe0Cs7r3mLU12
Hxax1zuUQW1r/InVeQmbGP8AVT2IABunwTaQ5ehg5fnmxYxasczjb179DaDU+wzV2nhpA17j2qNw
yxWjp9EY/vXtS1aihvzadA+NcB95ZdxOy5d/sM3J7bQEPkB3WG4eEhHKlM5a6bGz6sv3NPKzL03Y
kBmf8O4bQwOCXu236YTV9Cnica+BtFpmPcl5W4kOyKxImH7p+fnVYn2cOlm/OAbkzqHxuMoO/N0E
Es3eRoDd+5GpkuS4x+QLeuAvOSoIqQWsXfK2VGGZjzlUTLGQ+OUEjPpY+bo+60N5aLz6oCQJPE/7
jGmxTgWHsOw/2pDdMA03ZWHTW3S0KZLWOHUdNlmZurrMsrFJ+wcbpOPjwol4IQzxs5+5pqMletq3
kQ7Vlf4aqX4jZ6YQG9IDOyI5mjLT/Z/gXX4ZBBn5vBEAkXUYVr0pKHHyOY6TlNc+uatReE92YDI0
YHQk1cAWhctZVFJq4yvmtY8AQiccIa40bHWfLLI4O9CKkJpHo+fOL+1Tn1RFUs+hQtLCOL+Lk4Vk
cTW0c4iAOCqWqAx5oHwIxlGcrP/Yj/wABLEZxHV6SCWddpv19AfQ72Tpvq9QD/u8ZVKfi5fvjAvg
6ao5ncnBkKD2Ic0bluTmBeWu2lvvUM15T6pYY7XHEkkDeSkz4b0jxe+L2xkeXp9Oz4oHxyklKSpK
Z2zN4Bv/pVDW3Brln5ciKLRKneBWUpCLQcC8TlUJKR9E5wVOS/9Di1z5tq6LVegVqshBa/imns39
elqtu78rSOgTNp9V1KGesyDVuklQhFXmPRONXVK7wTK4k7yeDKpiI/kE8rbQ3Sg4NWqIKYU0G2lw
DvQ0vRF4zqzL+J+/hB5IlygY9GngIXVJbYSi5GTkF6bd7OwObi4/KBB/HzK2GPIdLUKgYo409QVl
PoJd9Qy1c/7LEkFzFdHxqz8ItES0tj6rOjxAzJA5aHsRXqf2jZa6JczmjVCONlxbbnCaBaWhj6EU
wxjimheFgDLCv0ZiN34Qu2WJgsOAkr0AZTBr72BqYxreg9HY4xMaRHLzVgQe2eW1SJVtXmx9OY8U
zkXUTru4L8lIP1v3tlB63rdiRRT8Fq/riRTMiRARu7mevxF2e1LUsZw/AfgSqlKEVALIJHbq1/1Y
v91IkPTwhrVSYXQV0sI5t9qXRhcYkVS8iewzshmoARAweozRsjSkTeU7JEgF5HvCQsfe5ChnCaOj
Jlslxu3a36brwHukFstMo4LVoOCDwRU+CQHeJP2ZtiahvpGp3VPmtaJAmW0aTXUCADDJZSMQNKq2
1rKipJJn7NySIGSEBH+/Y838kaBBucxE8a3yzBkqBd8d0LHcP3E7JyiYrNqpYZPPbgLa/yNq+fb5
rw2b+7/tga/3u8fjpQ7Vb/EYZL9N4U0DgbdGjcjqKCbg6HL92lJ0RhI+Mw+MW575a6TUVhPqMwoS
vWS/wQ0rUd3XRNWDaS/iGBrsHjpo7FiCkBgRhuK7ggBf+FUHoLG5RcSoYSFEq0WDvtOAet/adGO3
QFdQGBrSPkMxUNXZr6IOuP6xD4GmDp7DlA70iY8v4Vgxn1TpDVAr9YJKUikRKNCG68G6lLir533T
/1nlO0j7OMuWetHQ+VGxYsRtsdpK1J+To3wAjMhTcrPi9eCOKSnFqg+TaQiCFExNNP7ZhnsnONsp
iiZjfNOOa4HkAxrTtKv5I1h54ykBQei9KpAmpbxCZvgliQvnYgOMyqC8tyxy7yoa595YirmCdKKd
39SMxFJDiJ636ZQPifd9QSpAIx4kQtr3hbw6YtZhm02Gev2a2lHSiTiP8L+TSxqYrxgUe/pYXcQg
Y11Ll7ZqJInUEhPZYVPfK/s1j8mqw2C5TvTbnY1mNT9oczifFiCrU71/Iy7JSJDSlia461dNsug3
D3gjyUTkTp3MQVDaUdFHC5rBgwj/VDd77Gd8NaEd8IOXlECy1ULpqFqhyX+7tKuP2oHWN17USdWV
yEdat958j2DIWyDDxImV5ID0wzgo/9f7/L4/G3fEYvRVyCfPBXFAUigTeFqd9NCW0IvLGfcvEwqn
B3RX7z0/yTfu2AjKoqtnIjjyIe5ACD/20WZU5pHwfR/Ubx2hEo3QydzCq+B5b4FZAOG5ohtt/c3n
XfywqBO/hNxZs/oXMFkO4OeunfxCNjHDq0yWvsHuS74KBjwPseNRC4ilM+I7EZh25F0L10sa2JQD
IKW2rVAarReZekp45h2xk2OWEs85ExRUfr21ig4cmuNbhnCxxPW78FEWwsTIeICZkjNomi5i5KIN
Leql0YmZ1ZhUeYrR4KO+ijk8F6L9VAOC5fguJJwVh1AKBFDbTmbZ8//UPDEbHzZ+W5Eu8g65b/XM
N/dABjQiqa0mYd4QsNUqtm7Y5Z33bfc2/nhDwTzh8o59zSx4UTdqRBhgGcGgm3jliplNQczozsN4
WiejbjVhNEKIM0T+p6t50c62mXyzCKG6LNp/rhRhFExfhQj90oO3P+S+XOLAGbLCb/v8YtImfckt
qijFSJ3YraMdQzomaQYKoa2xoUgycLgVjawLgahpL1uNue296TZkjSvOPljWQ1V70LHZ29+7WnKi
aGKY9XQ5vWrDCOll2WA2f7RfIn7PN+znRKKFWkDmWEOpNsAtRjcDhF9FRrq0O4HI8Gx8VIqIAEB/
4HKc07w8yc58XqwtuXhy5Zl7Rviw7p/oet78Qa64wbNh5ueaPKRWRZnt+W4Dma8NUes3gTqwjpsX
9pJt0bD8/NTExV397x0p98B0wD4wvOWNrAkV4A8T3uIcZhnZHaLIjUponrFQgg99usfB3xo9vb+s
NSb7Oc6dF9NizB4UM21RsJb/vntx4v4G95Hp4hKY2ZKkwH7/+3pvHX4ryWAcCfPSws2AB8UD9hed
s5RDZ5SFto7eYK74LVt+SA70+NNRrEZCLP1mh7ymYy2L522YANpyuOZ+hx5/2Aakfpe3GLlyh0FA
Gy54YNXKNmA0xJcbjbbRiG0zx1LC409Ueevpp5m0B+sGulWrDh5D4czyc+KnYwoSc9lJf7coDFGb
A6aT3IyA22RsnrWDfXALasItm/QW2xqfoft+BzrJS/NFp5pRaViyTL9o0eY4bgI1nCtSzcKt74R1
B+xrqLoCe0UbvYoTq2zXYjfRlp5EtQurrcpHZBk4BxsnCBiVl1IURVdjD/F+2mtSQj67fE/vUqI3
xw0QtxY+1gyKR/xL9caXFqlhL4G6ILht9FG9/9opDdcBchVbKu0gWFHRjBFeQu3W6k+1wv65VW4V
gJekVN/Jvpr2QUuWiNR5CCZekHiIK3LRTLNy0fUBYvKat3limgxgrf7DLbs7qdf/vVPsiZaRsWQz
OCXPscjFRpdBbNUIj5uGfBMKEBpu0nOPRofL6qqTLuyzvAPe8G0mbNo9K85EzQ8+tIgfg/f1qpwH
OwIySqMRXrLYiD9V4HmfNN5P89hnlwadGX9c0mS2aS6yiB8udNQztJ0q3tF2uF4sH8NZVi/DHUrN
DyGxR3lTiz4Pmj4Xvmq4sSBD1A2I9yd3VG8dNUXnG59EoOtzHbHtGNIban45MMPI0nypsBJitDnd
BbX4TpsQoozo7xK20ydNfYI1OkBXwYieKhyFjjxlwuH/BbjFKw0lh61ngTqcevs3nLvx4i6Q9HH4
kYWSapgDQQlKVtFHB072Rx+JvS6+G1TTcBNH93SHn04WjNo3pvdsiJCTf/0f/zGNMfMYgm8zOVx+
MzOnldjqr9fAa1aX2kNojppewyEj5B5YM/EFr0tbNnkuvk/qVhMNbALvhw50Nh/7DvRKgEn4ByXZ
qaBIMYlz20tmiT4EGvRtXmClRS0NXBxxou6NSKXgW/xL/ZodZtJpPkbeHrD9vJ5hVAhgr1TzVRpH
I6qWKTFfDWPQMetHT6Iy3ps94RBw1G1XpiL9cLNShJ4lEDPig+HKQ4QAuaCP6isy/WBvAliWRJ2g
3vAQpTYfZvba88DTkLWIO9F8gSz4+555lFCS9qLxJjq7wOokhUY5ZK7ClGQidF7Cx2UDB569UU2R
V49pd65J/wJyDLNFhcwrhZ4HgsJLhIXrPh6r4SyYURgorun5Vn87LjTx7G046WAAeRLtEUldLVi+
rv/kwzc42p3QlED+7/nil+8UZ9lERKUtm7P37+qetl2TROZmxGFGOiYVU9cZigAQznX4TL+43xWL
So+e0bNjeEnh8+Ti/v/Omj8G1VkzrXHm/wWi0u163BiSuAa17mteMD5waEB9jWncrD+NSLGmMXnq
ySGlVnfGqKt4/xBofgciuwoopdhQJayoFVv1v/M5+s7bKdTLUPl5+EMOUxoRQpvUvs4zGb67xeMV
ryYPixH6/j3IfSzfilO2JDGoCG3W/F82JBoWh50e3blZVjv76Zpk57NE91wV2jqmbF2NJ1aT3xnA
iXZ3V9W0egJlek1s1UbWvEoOWmnNryGTsIjapan0M5k7RO76XeWOc+xZwZShQXOXigYhbcxcBX+r
son6FlbvsXSacrDcCjlG2al8LgMrH7+OejqeUb1FV5ZeKWKFXxoHFUSaR51MjWOfOMy5iyy751P9
bGvtao8uIiRtBq3B1tBcKMHPDVIkzlz1fD6dllPto28hns4QrBlmkOy9GzYgZIA/69oZBXINzGrs
xuHtXEOKmYvVLBeepP1fjIfYOObyrVvU0WQn+JpCSXygzIX/EjcV/qKZn/bpz1BV7LmyVysmsKVr
vC1GhWu7hJmEajPBH0AplUu7WxpxYpa9MvV6GLYzxravj5H7dFYy4wMcqxsee5paTMVNnrvyrCQr
MlOvUSCHPZf7dPEjO5oyhqPjOYc0bPiuS41sy7B3FBKhuIJ9792Wr9Ak8LgD1RwpswocO7j9ZfSG
0IIbXSJulkGG+oHIKiD9Q9WAN2d0po6vIab0fGotfw5E/9uo0Dbwb15qE1RdBTeT2Oe4VVpglvCe
JUCQQ+OB4Tp0Z95mJ7LsJhSlH7BqwXD1+ig70SQw+7yt/E++lc5cSnmP8AG0744mEhDXYhDdmp7p
ZUgyPUo5xuOA8DHXo3vr3vAHCCqoikGieG+QfRYgTBwb5dJwC0rb7r8igYumk+J0YMTptKw0uspS
5sjPl2kWafik2E1TcYJFlaPR0l0O/6sJeTFpT3aoW5bbrVO/ZiKjfFR814uxajMqUXiaYJxSzUmT
TE5VXlR5mDdEF+wIiqqlDuYyO7KMBOqMRAz/yRR+muLHFLVZX8D0Z0GU/duZgYjuTGb2It17I4wN
Jfx/yxD5U77vH551FNJL/GwYfbUi3Uj0EKq5O6Vsloo1tFgBj3DQD+bAptQs/0U4UHlIrDYzIXL9
Bg0R3fhKs9+pyK/y04fpzWmk9ouwhlvEt/4jZDaKR8XYoiLay2ld+idPesTFF9D+wumO5qhS9P55
aISSIqgn6BghtHjv8w5R+krpfX4kJ7FDvbq/mHYoyCJa30JB+ZIqQqQXNR3l3Kmjx3GGTB/UcYQ1
TtSkmJWPbT5s5UkXizq3Vq79/7lcSGqWBwHWBw+BWKQLFJwhVsT3lnqJIY6kpQmfqRs4+WwDis0r
pt88vFpMquXESmzAtelSC6QCcSYzK6tYa/io6JCa1J1qQ3EK343LF1LEVyJes7yckvAZQBl9ehDb
N7LKFoT8ew8qw6ghdBZeIGmu0/lHCv3FAlwGqngtKPDOQ2atAu+nL3FWBYIxiqPNaPsq3z6T+8ZA
1txi+K1NecZzd3/Gw7IE1sGd2dIAysa3Ky0Am4+gIeeE4+9Ak3YYHZrRZR56zePc2/KeyytnScIa
0AQsvODsTwWZWtFJU24nPjV4EjFAjX8v4YYp2eCoD+5RwN6gjYdVGEB26qQ3OBsgq09+y4n64x7+
Gv7SVCK/AB+BatTE8npUhelsMjq+FcTIRThFSDwpla6DRJzKA8EssWGtxpYR+V6s717fADfBJFAy
jBFSOSVhppMXIJHe77zSJcCvpqI5WJxS0IbIne2hE5Yygjswh7ZZtVdGDGhYYWqfrzZ2RJYlmUf3
G6FGtzyJLsHwp0ik+m88QgN5SMW1j6dvfr04Jrgh4yDaZbG4C7877MZePh+X2mYy72qnokl4Yt/W
GxGFRFFJijLPuINpUAhZMbpncKB/cj2SAbLBnrRbYBQUYDZHib6xsm1viZAfGHH0nKq/dDCnxo6P
JdOHEV0VK8bWm+Sb/QlMBANeeW8SSxaOjEcw0xUIV23GRATYkXraGg5YJlnpzXCdjB7gAjJCXCC6
mVPJ1ZecGdc3FQN72c81qFEhBT/n/ctosYjzVKGjJvaU2/6NSQz9jSBvHu40qLx1nuRYpLkwhMcj
u5Czer0QKf10cdwmy1nuXmF+L+LHfIqPtrJBQd044hed2Y8/+0aufE27xPLw7LkRTO+ASR4bCiHn
0TrGMQthYEd/+TOdkVmkS2xGVL4WoN0wtcPY3DvH0Ue5EAfaiHT+1EldA6MUEEwTpYMRsFexLm+I
ZlC243XZNT5nknzDVQ3M0+XGVg9zgAx2VvZ26HIlVYa0+vq7itWKFQYRPVGLmrG07EilgxQmoOef
BvFmfx7xVtftlFA+VsHU3ljDKShsa6e0Q00mglNLkdX52RSxVdBeE9D6iuldBzED88Zy/PfI0eDm
s7A5vwrO2TWEUNHlElveDss5XvqkPPdSjLxiygenQ6TrtTthxH1nI7zVITUX1CkLYv7fe6bZJbJX
wJcJ1QvBzjp8tXwpnxH04N6LdYJqH2nIYkBEGK2wzuf4BCCNBSksi5qBM/y01JB88vHnur7StgRy
SJh8Ld8LI+aKMl5dJWBKSV7eVCVQwMR3lbn5sik9KKwzFEABwN2nLSDAQ++myQj90O3Ln6j3MM3w
jjIMjrizkLz814s6vjgsJKJ4gUQNFrb8UxYc51Yv7mGPSeExj+Gle32QBW5W1oD6iEkj0wFFkx5p
NLuIiVAa5MeYfHZzLiHs0NgvjZ4D5sMU6ggz9OPK0DZf2hhQCIpyJnFZnsPn9rV1xSClsthK2OQ+
fXFYqY7t1tmK/2ZlAIJV0Hj3sx++wODIHuPUmj009zGoxZK+Z4fF3xmOc+TzlNJhvrUm2HfxDPyM
LKHAuyzfREv7DcJLA/kmVY39YVYNVJMotZJNLWf2riSE3+HE4Wpn3FBl/j9TdPYOrP/xVRKmMQP5
67qGjt6KYDXN2M4T90KUbwVwlXkPFuWbG365YIAJgHQtrc5oJhBHqiNxmra7t3YVPyXivfmU2QvQ
RA7efNxRO+vlRB0bOlNFsuroiRWUGztvhQDEvZT3eoTQMJrp+XE/P2nJvipqi8Z48F8TIQ7KhkB0
30buhh+965iz3O7rY9ovb2QGaKby65IxfgXCkwj/FyVy+ejdTBz9GmLsQ0U82duDDUPAnOw/QYx0
PP0GjcRw32SAt+mVxdz2cky4K5ZOOPPKtZeM+23ZGH74NFcA0Bdo0E9xirau3fVPq73oRa3YRWlR
3Sr4Y873EbQXDJoicRq434uVSDUArODCvFpJUM9Ti6kLQF+GopkPy+TIE/MXSM9aL/73Gfxn8jHi
cP9DOLADKW7nnM2giHmfGHRJ4XeucL0U3QxtKeu6jaL7mfqSzyCjgu+qr08+nOBbjaboHIy1nHgR
bV1hFl0lz6YIlWzqp6ZXCaedVm/vghFQloLB9LJfJMnT6pxomVmyZn+7WQMhePQYTfBtW5SHn9EV
epZ4s6Tbn902OMivodfGaUQIoH8l9CvPzM9tAC17vNzEOSH0V6I7DY4DZr8eBaWQZpvsMhCbilNw
fmTuSm8fg4cKiU1eEaKPuoWfssvrfsv66nyvY0dLBBeX52onW5XOsjNMsqm9xVeGtJJ5wxAsen/e
opteowO9Qsoljeazibgfk16mzbo9L3y/pducvjqEkdc8/HFtY7E4xf4yMI5PVnh8MY3WgOZQRwvQ
Fw7xE4mwwo8qtpvZbay945Np0q5SzOXpTbU0T2XuYcpUnYoQoFLzS4J5YLJlNazn2e9lpkwUYfPn
tf8XiFVtSsG6hj2S5+UY7HldeVMQG535OmBfPlfPfXpd4mGDKl7XEpdNISmXmzz9p0msSn03AhNQ
c/7mgiQQl7Iuv1bmTMCqkXSmPsUR2of/+G3o4EOBXDPKPIiwa2ye/xQ0+prWNfBk6GefIXRpehDs
ARz79jOBsuqN2siYBjbJck28tzxP/dzQVkLM07/hrrf8zLtxSD6Ee8wjMCUQS+yFIoFtAl5EbSqX
xZ62ale/DjDRkcfUVdcm6l5BRqd4LNndE7dQBD6y8fgRwV7/wWjGaETfk46JuHUpzm0xoHU4H6xF
ZE/j2NC+4JMiUFq6NSoqndEbMrFnvLtr+q0FsF6+V7oEb7m46KN21n35uR44e2lJ3vHeAfF0zbsk
/9nOMJmw2GUAy1J+k3pfTV/inIsPCGLnB4o3hSBfe/rHSzYIlyYGneQVBOR1KkGMrUntu957HHrL
fBhG+qZVbEl2Y9VX6gLCz9YWPwzYw0zdFzNA/FkNWnRaujaWrnfkTo1DpQaITmdezNDnHTXKrwM3
9NvkxGIEf9ZkrnDEvK4RC2qIp4itJG8xn3BjYGq6TRrP4FJdcK0Iuy1nD/T0rdB3dD08WMVdXhV5
1P0FsrKApD62eY65re5QJ1RMAWdkuJj+kY5IjvwjVyI40TXwxrnEfSGT5b1Qx03DsxZ1tOsh4sT7
k+hqJheyK+7ZGXQ7WwkP5+bfdDavY40KJnbtT/cWWWPSOF6VTPs34GY4ETslW6pKk+8j6IH89eyN
vMK7FBOKJgpdE+Ioe76+tKTVJUfqyufP7sp9E3nqiN0B3kJsDJ8JQrvV5Uh2Y6Did6cx5IgzD/eP
8Qm1QGdPn18bm3cXmmwoFDAUtrmpu1f+Qe2/H6qBT3fmcn3Tkfole574DWJymSNcnv9qBfop0StV
PlVnZjlBR/nuNr1mlH0ZileoygPtkndizWJjJG0Nr9GHZhIlC5GNglYg4qNdLf6HF+h00wpsESyy
Av0qEoW/TXi/66mlvjC1AaPJ186xcasjIMqgGbpmFwGDfGUFfSA7ozsdr5YaOHUmRuBqFNWAtGWx
Jswpyr/megs+2fCuRt1JPUZLSUZuZn6qQlrYhCI4fGDQ+XGp2NPxxlJJztfoXaJC1dPMFeTN0PuR
rKkXqOsB4Pr19y+R1KlIx6tCVUbTK7yETKzpjOduXd7BF+XzUjTb3sc/0230AsiVSCNkCm+DFm9P
1enNDEV60iKw5fxRLEuS7f2QLpc+G83j/KE44c4auqLwLhOlbH94n5bGmAAlahtNAQi+dMFE+Cag
9cwngsKhmAkimaSzta8Ze6Ucv2nb6WIzh/+P52fbvtNZwMYckXhq8DnS/vqkasUoGrNDw8xp2kEB
Nc2WgYxHtiOqJR/0ptFfWFT7380E9A0jZViuJfVflmRZS1IEb3wxU2pexTsTlGeQQdQ88mEYJ7oI
P5nU47RACRlaFpBsz2ZhC3nzajJK0LMGvHXMNqrkWM9rqLBV3TrvBSyLOKwURptL2kTKRCHASVbP
ns7RpewZzDEoiSmPLT1lsOi97mJMxMSN5dei628+NCOEB1hDG8EDa1v85IdT4+gFR+6dyMPhdJPG
9WZiGludNh2hLh7YHxgVlDJSn3sPMorY6UzPs5FTaSdoLLoUBey5s2iFMmxFg9AUJ4SFwzOGvdPL
HLmxRk2pqYskXxeZ5P1eL7ZJa5X6D0prhgby7w/yM6Ka+zSyRM3tL6+ph+ft4xlb5x4UJtcvmQOa
UrEcLoKzkiOjHgaa1za/mO1TXQQh/Rw4jphoIs77ma7r6huItJIRCILpUNE3PthUA0Z7KaNQ5aYh
fbwdAY/O7xuSIqAe+27RESduYrVSxJu0GJHPoEwwa+gHthpMgBmO29umyjc0cFSrJUdBawJHyhfF
sD0NICCiYjZ2E04JcIlkMmTB6wWWAzqhxlcTCLkGrVwpXRwt8ighoIDwehsGcZizNEwnAo8zlUgr
eww4uS7Nb/S1tfYv6kWE0gz0l4LhVBXJYmOr/dO4j+7Sc/lEWKmwSdi3wLfDzbn0iSEIpl24e2XU
OgjcVEt651eD3KiAVqZDm5KLOxeyJxOMhtiJ8KLtlHohBy27cWgTmtROfSj2eCOdM/cZr5+PusMf
7hT6PHN9l+OqzQnhSb4Nz7cVK37GcnixrZcfLvwFhzMVGPPYIo1rucv6FLh9G1vYKfFmg2fIBm8U
z4N2h+tTeQgwI2ZV2A56oLv9Csl+8zKsCDPv3XZY9RTTDSKPDzfHOxKFRoJwVn1LhSpOsnnw6nyy
E9qzPNB9npOxLhCdq7Sn/vgtTVw4pZbwH6B/sKyBD1/hiFsiombz0sMs4/575eEl4yeCYvmbimfx
+OI2gMzvkBoFhywyXShTkYZlrGlMLEYaKjUyTiaocUtMl5EdCVThdihcS1kK94gBqI6Koe1644sa
PlD5BCsICskG5grjO7YEGb94KZMG1UV91sWixsf4ewbAhbsFG1Ba1BTQ+tD3+WL7vVdZkiuvLuRi
2wl5EWXvZnLjI67QC85fofm+aU1OVZtCSVIqwW73C2aKCcObnrvhIT6JDxbwXCzhLK/kZhMRJRKq
+PJYYZjPiddxXhdA+UgYwN7ApeN6Zf4VSRc4d9v9y9iCayZzqq4YDsxNOCz3qXRX5arOQ6RxpQfh
L4GomT6FXgRiE1tFPjg/vSUb0uzy3DUTGD3qPxcxPiX8bMDgQVDmYaY7YWIliknyNNLYx/6XOBNZ
aDJsZWct1Ix53LyScxKLdHRyRqf78cW4A9KxcTp+fmepXCqqLLYVzPXIhfw5Yd3IE6JKfreJ+gcy
+rIMjn6Z9cuBu4q79WDLJcSZBiJ9QCTi0IGqt5O/tXrtuZsOcIoFgSGGLXGJ9+OxPsy8+r1/HyeY
r7AbtZYe6wIY4xqkin8q/SDHVhYlLc+KtAgVKl66675rW9uDKMbH7KrUE+fTxVkL+bQL3wB+TnUv
rtZleQNd9wvVPHZE/NQJdQP1gC8Xs+LNFMoq16yAQjV8Moq8YRDQJlaCIqJtB+oamCgrzp42NSiT
BGc+sKQ9QgJv8763QZj4EvaKuaX+9GRg8QCLJs0L7JHiY4a38mHXcsrL+SKqMhas3I0fgPaYtjaI
b+CHby2rYDsXpcjgcgEzMxFPlKqUyVmRcmIMtmLo5ql+OMno9ZoSc7EvtV2fBMguSSwT7RtB6Tmq
quyDP9kmNRUrRtwYZV+9uGZz3RHkjaRosBacFXzDm4CoePqPuGSoKOc960SD53vwCMRDRhYqvQkY
NTEza3p6EnOYTFNGnB8MOm0w8y7XKj/J4IIOiwA+MiTIC56C4PU3R64+y7XxFxYym7yyRwKzHIFa
V3nfF9XLsYy78qUTylLOTth9FxcvnaSK6Vz6Nqg8bakt3d7KFI5/1VMSt4G1NNg7yKwDpW+Zf6+K
0rxi/bKd7VP+8G42Ed7fJ2TyzcTy06zBfwIHeoN+4QVHoueH2NbE95JXpWDInrskPySF/Tn1FKC7
GP4sv0mgGtbf3lbEEnuu/mWWntsx0YcTqPZxVZVoE15qEpQKlKGq0fgc1yaiLaMMsFPBENgFXeC8
eHhSIcP5wtYH5RlpCFzANA9rZyJJoS1hqUyXsC/EyGAupZwvAk5tpzD9rQm3Xn/00Bhrf8ehF85K
7k8s/ThYUHXaSXDPk7udSRumdu+4ksnCNl7KBjj7tjBjKZma1KdPZEYPzgqK5mYMcI7rNNBR1LEs
CZ4pBavjQWpkPzHr85+8QF92j50tCi8I2nhfVY9BfRcPtjUsy3mX7eoOVE1Rf4S2L7LHDlLmTIm7
s1j8hlGEoj9onaz3ahoShoklifSWllMxN+9Q0MKfgi9NQoeTpm6SxANP7tkeYbVJ9z14etHWNAFB
FgmWGVcq+WrvvN5cs9XwacXBg8v8O6epfISYvoUlSKgbirgs1DsK3+sm0PVuFADd/xOe3n4YBY1d
xvw+6ZXFkT0IP1qGyUeMP86VunPNZDflHHsZwjwLpPHWP3JFNjEG4D7tlzIyJ1LKCFp1/jVq6ZRS
BeFlRS+9WpZV6EVu4TGw+glw7LrBxAqD3aLATe70XnxlZy6EawD8zCavkayoio/fCvEUHxAYL/oe
7zHbZZVfGDuul1oUzdtFv9aox9ccTxsuRLHyNgXkOBx15yopNDWxlt+zPs1j9bP2cdaQYKwU+x2a
blAswJ+q19KfxYStzEmMud5iTyPk15sJ+r0ykP2VvD92XVXtIv/cMy6ZLe2XpyxAf/cWlytgvIqq
FJUSImmyiib6GPFYcWpOEW4Kj1dLrtIrHUY1zkAnnrF9C28lyhj9M2pSC9e4OedCkUmHYdGZjCsO
6BRdD2XxZB2VjUwVO98w2B+i1MNsWDdrUCak3901f4xVHzdhdwLyWUmqW95qBWYBkQ4jXcaXq8hr
e+rUL2lQccuyFBEBNCHdH8c47+81FVVsase2u/VPrC1fYBzNH1lJFwjk3wNt3FfRmuOtIPZO0EYH
P+J3J2emZrdBATeNA2G7lPNmDgg2IwY2HxyM3gFcX1l5w87vyASfPNb33Y4SRFK2orDFBinpibqK
6mgm8NhC+oEvvxdb/2luCvcO3T1Odjvor7Qscuy+/M/gISQvELgFQ/qDUZeZhTM6bEqnyHuflfGe
eEnIS/a3Ym11g0tOJX/aLgc41GF6dtX+Vci0ArC9kfzksqaZ9+GfkbzbkrUpXi7e8LxkcoaNWAkj
mxmIPn+HnINW5348kn0cIcWspHnIaLVoOemIxPKuxVt8iaeoPAwSpv/3Rtd4xGzHMN/r+KWCz3UU
E65FWWpydHCRFxBA2Z4uwVIG5xEffabsP+3tZGQwKfQNBPPedvyWCCZH9rkfEU+5gW/wGU93VAD2
tDnjtD9bGVeCmMlpmiX6ndGa9xhzaDftxw9mrmKLKE7oWHlzkRy3+5ZyPEwdy1+F7aZK6wY0xPWc
xVUsg3HSLgeN26hEWFMtUpkRvjRkWdWo91nA4cL8IeF8LAOH/USwbeuF1uG4AHp5xduytLPA7VBb
4kkpAVtBc2RrJMambWphlqJ4oriJBtYB8f9LsbWuQnGSyXafxC0HuywUZeXUlREAzqCYR9K4VCAx
l/o5WUcCbdG8lKY+TwaMIg2oXVxDHMMngBtiL2eTQ+NmB2QbEqfQGT8EIlFy/UgeL6AArW0Qr3ab
xmiBDuakKlxNdmsLASEopoU1Q3q3A2xEq1tPlHqd21aClTeleH6yNrA3VyxGw4Ti7PXJAMoUrG10
WmD5+qDtW2Ii7hoKdsjBKeuyBsF3ygSCL1+qftw2xWh7Z3wITcpgZLbPkHfs3TFNj+p7lcx1xjTV
yR2+lNOcXYTQPrW4WaABwO3RiyuBuN0XERDMuV66jXmGtnOzjVlplFTl/i1jjecP7I3PnreyAJ1E
QcWB813SbsooE5pN0DjTDsKwaPyx639OC6yoEYRkgiCr/gAJ+kOuCb14lldOzwIC3u4zZC7QBc5M
IbjRQQXfN1SYm0NxvyPezoZ7k6fzND+g+hFcGjzIRu1DQvlpKVA+BNbfsnxxJ+Gc021dhiK18ed8
KoLgtqSnF0UkZoGOx8Qy+ta0G2kLNYpRJ4MX6RNtJIrXj+vaOjRGmfTinHjpwEzr5vlUsNgTtFc5
+nuLLlsJoaYMZI3ZjIBqCp481stuJ6lvCWVJnyRS881+D2XPxSia9E588sK/Y6m7Z8qbhl5REcnJ
j4hV/q+e3b+PO/eiiYtmvIre0NEtrAveqQdhobv3M0ryp9vBxE3it1aeytb1+5SLtf6Cl/uArnSo
Eg04Q22LshMw2vgK5uwKkwtDwx0/pXd0J3icXcm9mM6K6IWI7x/cG+rQReztA828lomCfMwR50iA
TFWVoIGn5711AYPs7Yzqm9dgsl/9MLThlmCC8s17n1z0BHCjPvs7IwNFvQTDS8OKoP/DlisVa5kF
lDxeK+gXxMT8/ltA0a8qeUerz06yPcpzlvJRlGz6BqWi/xl0uUGr4ruWXjzWusLzj92yhLiqDfdv
SM9fPWaTO/oVqBUT7xHxQY7zLHtgyGtL9yEEBwZMR9V7NJWUEVP3IXIeZe2SydHgshUSKzSztj6e
RYzj4oAbW+Pc8lx9efRFVuqHhw8TEFR6s1X/Icg1EUlU7k0KtfaFbA2c7qEdrwZmWk0gQMzlEmYM
P9JROSOwMifsgvWYeR2Ijs92OuwkwCOB9LYmNg7zxii8HNyndayouHSRPDb4EEDdz+yidWm/ThvG
FOA+pjYJzvtf2KU0Kdw5OrpOAkj6NEpC1lfPPWMGpDxahvF10fbnB2GGemL7gIQuzY5oTRbFhseb
8h1DWqU6ehgSmDxyUBejs/NOsVu4ODDejCjid++bTlhZIBhepHxnMohz0URMsnmB3k6b3pWZPmTK
uuS+VtHm98lQZJK0wPD0waucrrvJA9TWPZGjvSKVVO4Top4rR1s60miXzZiazzvmceMTq8n+yRfg
uJ6eYF7ANpNXoz2HxCi6zLXdfnBD8MLSJNlgCWiN/9x4ahTRBaV+v3JLBJLouV1IuCIr2FWyoXhB
hb9fjUgsA/WtpixX3RTgWe6TfzfW9re1awzTuTAD52MT1hbVZ0sbXEcfK8UHxIOQL3btbAQ3jqge
EwqIoo27GnHNgvBL10mHaLK1f+T8CXmLBbaBeSitJ3Yp5COJbOvskkK3Or/WO0ziPH7duwV94QLc
M97Dc0inMMQruKQvMVc11+eQCIbBAvoGz2OqMSvF+dCa+wuCMhEKrDYjjfSlrppiB84xcM+ZyVPe
sUyhXSsWNYLuYjovON+3QgJ0rGjzm4Z7RRS08Qs4PGJ5LvnZycwha5bFFk3omkrC+PjIYSLaImt5
sgoxEiTiSJQxRhXNfzYRPyl+E3lFj/zfUzIyyja/4WNcFHeFwuvsb3ZJownjgYTqpvSHWICRzJTB
Tz+dWb8jSj6QamKWTfrlwnnZyK/XYFToDlO+Rsr4iPkuutAkrFIVccjffDdj9OnaniHupfJJKa3R
2BFTMG4RllWXsDJsAxBPpRgMTDVZkpO1gFDl2kMOZqztdQ9y6ZFVWrGGnLR4+Bbd1FRc8dHvHOW7
cc+7cDWWMnd0HgNYoOU0gSQb2BoNmzsOtw2GSFGgQOsngVGzMm5zPwXkh+dtNlE5wv1cK2+ho41D
dy8CkxR30upVPbDyRVjANuR/PIN2Q3UUzKhRu+JMrytCB9rsvKj56O6/65tZFNy18vxD7kXzoIj3
egn/nPcv0RS0UJsdzzSauvDVA72rCoVPiwE8JTmaYiY6vFWe05Z8EAEe9T/5X9rXwfnA/+tt0qaa
h266kRyAb+zGf+8yp6CSsbqzPgb5jqfn8FgHq2OH5ciLo4aE1hGt3+3V+6s9zy1MF6LpDt5jJblF
6IjFoccLFwB915h+6vP0xxUt0qu3WYilivOtHkJw8XXr39bfFdK4KorGruTrm+1xIXGDaTl0Qmma
3oYyWn+np0HrtBOh1R6+rWzGw/tWkDremjB1T8FIyaTStPLhKT6pl/s1wfv6VJpfIWmML9DPLW0T
Al0SoywVGp7XsageaNCjNeXOCt9cxNW7rpF7+3T/kSl7n/TsMIPh0awA4xRj0rWNeCknaen63n/B
+bi0ItCSomW1Xi0ks7iXdzcHl6euHMRxtiVQg24sI0GWvA85ElAWvoegGvNZyyAFzhkab/ve4Hs8
VuYmdEIZ9/EuY78vdewIYuqpdDtC+S9kltQyR3onkrNW3DXC2ZlB75NvvWMmrUJZkILWyj5tl5X+
FqffcKJGHvuNUjxxp2yHr1/ggVsuCO70VdsOED8KfZsfflDbsMkgX4PEvgZefYh44PG8/8cnrI0k
1IRa14f0WpazR+bNSe2U7MIn5PWag+4Tp+dXkhNqu4De2eZXU16eW0EeqcAB06e9GIt6lzCNhrfG
L6QkEZnDc+Ec84yCo/ZPh9bnIdkXuSyHF8txkPOj3FdQaqTO8ZClsj8N9yhIffB7Yy9+hxyDtcBr
cq0tR2xIbuOod0+4ylIZ96gQIp4AueMKv7R0/DCgnPE0IIRBXHfONrgD9X8gFh+CZZETQWogpyou
9fmtM4ny+CbNfvqmWmKMfECie1WIBpPsNN6zVP+GCMr2AFKl6awaJqfUYZk9/+xNbOd/m1S8I0EI
9XgT1Drpd+uetVTUD87NdRPKwBoGBAzfKpCcOJBuFo1TxXj/SM3ZQ2CFBHrd1nXwr7C/aj8nAI81
aoZ6s8Rv+gceVyBb8tJhl+/E9JjiPiXkM8wvt8axVb6WxYF23B2ghnIDjqLAAgggrlDck0Q9lKwl
hir79tyqBpIOoP7xM6+GBn1QbyYP660EuRFY0RwXFm9mchsssJW/Nnry97+J5TL6TXBESy5+9xjc
sdxd5rcjNFDdtSOpzqAU/1wXj2tgtiCGdtn/43SDsYM2YcO0Cq845vsxhdksEGAgarj2zOmppL7H
IYxvBeVZsTdHfYd6MchcAaeiD7jH/yyeQdfEo1h4U7/C35SC7igt7EYHmhjVL4v2NZd0+7qQWavV
S5jYhaGRhUsMMT+Bj7OGlY8cSa+v3WuApbqxO/S6Usc23AGEgHE0iyFd58Czmn22PoiOVCmN0fIV
F8KjJBD5E+cLkZ50c4TXhurIgFnyW0o7aKRr7HB/Kt+I17uUkRsywcE8/fBLW3iBSxtoH7iiaiXf
lldws+pJ11rD+9JVz/5NPMHeRqRaEMyQFe1BCyD2U2oSoJFN0AxtKwttFRR4C1sPgUnyZXycQPE2
YUoOBzKBlxGjbNn9Er8ZUBdsAMuyku5sKy8u8JyAJeIwsK996A1k0E1P44JpiG9Nx6y32jclfPlE
SHpFPOqTv9ZPEdRvp5RVgqnONqZU5Bg2PoYtRGfyn+9ZTho6fU8TNVXhcEPQiUGggX53g0CT45Mc
sw+BbArOS2Sbh5ZtOFYDXMLw77KYG92E9/xaODl3Rdk7qooxGMYzoeN5MyS/gKfJ/Dc5QHwjZ5n1
GdyvQmZvB2D0/0nb/RdsGXWjWPZ+cSvwhJRhFL+BahGzY1ja81ZRyiTYRRjN44R5gDFcr2iRV9Jk
qo3LJE8YEIW9/7FI5V5+A4NhoZ497teqFjJIYAhyrXN/DYowrPIFBLLhMiz1N5DzQLTfgxZcNZNn
QSAlExh9jQZOzayPsJoHkXXuW9qrmD91ebWSIOB9SnJyhRDbf4oxSmDQ2m3HNcasqvL086jMhsWk
ZYy989O7pOuo2480ldmSjcRsxt0CHGiYe5B8XMCNve0oUWyNFP19fpPtG3m5q4yFJWjsOat5YPkz
HAU9OHL4VJZaRx6FpPr7CiDaQI40cfuJLk4mT6AhPoEBv9eAIlNG+cyFGX+qyoP5/Hhhaw9N5FqG
QG5udn1pJCf+ih9fXfrr9Faz0lz59S310HA9uDYp48LnI0canjKkENzlZ4M7liN6HTXY9acVaErP
FU2EqQhumcHK2LsKOnlIyS8ZqPtNgwq4P68lmUogeTjCvA1HtD7Ec259pnllmh2q3LhkdikxoDLW
cgS9cGhJr6cuVaCAyo+NUSUlH+2irRtSMJwAG84a29gnXK+J7GDVJRRdD61rw8DIjGNWvyowIoUG
T81jXgM0pXWFwIWCWwlPQoB6EVE8rmr63W7Y4SSTfsqc6J2S9ibEgOox/LgCDyPkvnXMT1TZzkHi
A0SjgTfJviGt/8hDC/MLMVezsQWOA+sRxHD3VRnzVcCdWRNo6lCSI5GMoIRVkDGcok/pbKYWLYFT
tF1VUqItuLQ6LdTDTIrA1aGLLA8eSWQEdsoahKNXXWYcLIwTknDDvKzP7Nt1pKEYTgTrIp6poX6S
j+oMeZ8dQPS8B3ZNhaglL/hK/lhlZ96xPElulTAAYEPBgF9c1pDtKAl2907YVaz87dYHN1yks1jq
xEyZ6rxkWmV/9f8/qmKn7VyvLmBV1540bjgC0KyB+M2GYQYeo3nM0Bz9DiQoODr7dPiUbUVaVQTQ
749vqZFZcZaGRD2KCaBmKwo2g+KcVM1EZvsg49o1ny2qmR+E+aX+8eXyuxYR96Nas+/jgdADw7b2
Gj0o425/3JXk6pRMtWCNHOcyTAVZKji4FUXS4GX2/kVjRYOjFW/vfNUT/sqcKFD6/kkQIkD+gzKS
YujEgiyZQHZSi1c3iR4UeLtxtKsc6CwqKoQekyPdcpR8ww0lq6zKfgAtSRmgva8AQIb53Z9FVJvv
VvpEcgN1ygETS27u+KHH7ulzqFLBcB0vWrdSuRYCUlUgPMins0V1Te8SP5Eu7/pjuP9/x9Eq0rph
HVa3l47W0QFZb8KF5usrQEnKkzT8Wlu+RpR6whIAuMQI9IYTG7Vz8NuIKPzX7farIFURRo3deoqZ
ReehZEU+Z4v9VStyT/JM4h3H02tT67rCKQb6UyJA+pj6v1sxQQRSeXKQ6cbS5/hU2q1p8trqTN7l
wEzEHXEvGSessRGLgCa6otHgU8VsPXmw0EwD8kPIOUPbYWwNy/i66n4lYAp5jHKdx4QIK70dwZOG
jMDJj/q3L5nLIsMYuslzQlRKUx9pJoUWLwGpZdb6CuNdf+GzEdpoEnYt9TS5XDgjVnWc23Mbk8ss
L9RQIKgqWU/SfJPPS6wxt4Xx/mhTAynPMpEAE9lABKXqfpC2FMNMuzF1aAsf+YC37Ci3yqmjNwWw
Jp8f5+3YSc5ivRUXUuSYUoRM1cCNc99+/LHvEd51WsLsoEZGHUJEh85UjVv2kmHsjfRkl/NoSXDT
8cjbo6i7wul+TN9FC41gXFxymUTQny54Jx9lhM50LlxLaHyWHaEUjMTOzN/QJ2/ICCfDEnI0JH4K
GIJ5QJgYEbzkseICEENQ5O7ZdPBMawJOqcI4wrIzQZZITKc/H0uVJeDyQeMarzD0B5lvA41gHPeS
17ZR1LI1Xrz9h01ppCcEHag9gPCV1ciaPB0rwHe5WvLa+cKkkWzJuFxV+9vGp/vJ/bSee0hgedN2
bW8KRtY0cmyNaTQcaxcxpN6SDqUB2v/keQnZbl7EHgi4Wmt8/kexyiSh8tVM74DhlP03BHc/wia6
2AwIxL/dpP+UyUb7JYUi90WoFpIMieAPtA0yDRfF92LHC7nnw0G1O7dqx4k/oRiPSrAGdfkSXaTV
EoS4eir7Mg1kraT2z1IOaAdnEP39tRPj6m3d/7Oylrf7B16NPvTLVc/+b2oyQyoOsKrBwd7DpJoq
v/Qvxb+qOB7tpwNfZl3HM42h5hP16h3V+NsJIn3OuO85Gk/X5FVp/rmlpzgINIwopO18iLQtdXOh
BPFTFES2zvpIi+A6P7unnMDDnJyxHLGfbA5oChjNCE1xeX6OcbuZYQ3tkXKptzFDAOed+2xB99v3
whXIJHnfaCcsRsCkVpXOo7+TbliuQ0/xXQDSOGME6n9gEC06XBCsObRCIdydbN3xrVbamkljkBDb
MNo+hf1q4fIFlt4EMEQSpB4afKcexrTwhXJzbEM1cpfF+Wisd6DPXSQyf4QB8sEDSihQ05YonF6M
OpYVXHEiQ+Qd20RZtf4kEveCQGjcixFaCkcejTGAxftJ3ks4KWlF9sNLWtpxh1B5t4bZSMlOeAHt
5KVrEbmWz9oJpcSu7Lz5NhYc7L+vDFbRYcAOfl7UchJmob3BuOmJF4hbjgmkuN+TB9a6Ug2yXWaX
GYXiQ3ufBG63L0S1hU/hbCefpQKHUI36nUeuh8GJZhk+1uHOWxpTDeYzHgO5mzSNhqLurewEnJtN
lx1LJ3SDLebRXq1vpxFD6Mf4YnxonkPOul0nW4xjtqHotWj7o2VCTE0vUovH1dcfemHShe+knFAw
NGSV3oOsMrvYFfWo8/kuPtILdfVN2ZpAFZ3NxUbdRGjFaG8QWBifo55BSjKNnq4b6YYM7yEPaCe9
aiBtCgirWd9vT0FCBm6Cxo/jfC10qaL1EXr0AlU6R3Di5jbv4J6LWs8fF1rufY6a7RwUNbw0eKJf
gvdhb0visY1TDEnGmiUK09yrPD5sGFqdteuUrnjW66uCiE4mm3c5D0vb1pwhbOJii7YdOpNFLg8+
9VTGjVX6uT6+XrfcFUKvOw5lUNfWuxwcRT8imkUfkK4H8MK4nrkzpmJIqoDefiXyKfszbbtYU/vN
XnrT0C25vnLMwzksYtCQvgBm59Nh0rsow+VMPm7l3sIHUlXNV7J8h9myh2PzTmGoT52WF3qv3uMj
IK0d7k0RL48nEJcuXMbHmiPfEie2LI8Zruj9fA5tNr1RPmNwEnq3JiKsRdDe6GR2dYiSy6KVfb+k
PkowBAeBM/CIBSbWJHvEhhYayd0dCBE/UgykxNFRIMhxUif8NTRrIcsn1zEwj+ULgB/lNrji+C+1
k59h0D0H4hW3yMotpuJg1NhRxMR6+BFhuP8xq13q4cSb4p1UbAl6Lto6J/JnWYKG1RfEi0U9gNyk
c9p7kjkkzYofb8/2PFE1BHrbFdCr34aIx2fW10sfxJB/T9MnrG/92EYDAdvTJSCzStRYHI/LkFqi
SgryZiRDGaManFMw/RnDDsDoKvPOKLRwXDn9pePInAxje/9XnIdmNCRS13lMpm9Zg4g97x1bh0HE
Ht6gwh6WytDYY0RBwpBTLVJ9pKHym/N0zl/WfT9g+1JD/5Fg6t/Gko0PiJDpPQb3IdIsPrrnDdPi
FwdgaNDSvKxQDtFtFcxvyiGtAdPwC36dvvom/HD2akQcnKucNBlyirT31mNcSVC9TfRc5Z/fj2rh
M+oEhkYxymChP5SCkIQpF55cAhsH+5okQyubNL0p/raQx0cv+FBi94CzD8rTu7ELvAU0HEoDStZ9
g81+FMS5hR3g4WwkaBr7NR/9QEUqk2MRZRQbTAH6oB6C83FhTf1GtsoHZc5Q7Xl3CqsSMUKI1xFy
jHMrkT4HddPqYwQIAEqCpePswLaX4R8FUK3r0cTJqkfFRdMYfi37Ou8KFFt8zWsnT7v636934DBd
HKrZkWRGk0CHAcjNK10ZtByahqMleqikZHlvFEolX6ZwRSZVwRWIFkbY89Hoonxd6cMG3xSqJQW1
2DYP2DazF2rNae1BQnQv7yS3WAdGk/U2JqW8pWmkE8wuCG99K9jkvQhyPJ1NNTElajT+DfLzQreP
nfpF5KEqmvbx2AmZguuezAICfmpUYptwwrkX86my8nVg2aekQ2KIY4aleQAcZgvJGGt2SqSS8T9M
6lA79pe10ShgYo/kOi6hSdbCq0wsZBzRdWfIEntLtu++r6J0MsaIg/GgnZstg6t3Nn4dNWeTtpLr
E5Lnp81UY3qLSZDrzoT57wOA0aGrOzPhn9Vpj/8SYciGNLloL80xFhMXtQvu0Zo4SztJdJ5y8ez6
NMAl+7d4VcttIECVfhaoul0c0W5wfVg49vJOBeBkqoj86biUEhucAzhuuXenQsXMO2F4IXGr/2NZ
+VbXVVlmqk9CIdCqkY2Rw1uvy6Yk8K6NuWTITkXskPrJ/Oi+L02RCdhnBG48kAiYy8KWJ+g/0/FC
VZWDUiDnW6ZO/DRPelIUCqEhAWZvs+ISlSiOuoF5+YQxoccTtLWFLSOzSoAWxZHsDlcP3431+L9V
UG/VdDZIXNlUtgFOKMOkMe3UZKNTXKx2HxCPc0WT6bV/NcgiEV2oSOMXjSN/t+Knxt18fJGs1MqY
BHRsuJFpZWdC5ddklZVIBOxqYCe7IIQ7PXyk3faXY+BaTFeKaG4ab+luBj4fhFOhsV7kjziqfjJP
WDGx7oTdVuX4r/sz6J47lqGSiJf9AZTXxG7aVkjSlN8ExygMXHa2FXdpEj6PUnO6T5YMH+oLgllG
RQxhlvf1uJgEgHg3f49I0I7aJCQtIlHofa33d/E2sEw9gJ/1Qw+kAAU5/ZEp4xUIMAnjfIu0fhWI
mq17V7ihS0eD3FFNmCf7NeCIkLsv+9/tZ15OZnebAyjTWe1vHpkMqF/bZek2B8k82wFHQQcpqmrT
eVTalH/WHkDhA5flY4xQAz3pN7m4i1JPfJugdyNECja1z43Qyg/uNZ6HWiacNVEN3Cdo2el3SA8t
lX7ByrbPz6+ab9kNhuqCX/PTMTwUqUqZUo8mzgVUU6CJPC82vNg+G7yt1zD5+nkbyB8SVnciW1cs
HAKFOJ69GN73FcGhYi0/A4m7YWKVsG0NIYf/PIA+NCS+yxN7k4W3Wc7fxCDGScP0rpff53AWiJFT
qJ+cqUc+7L6qkj+QMLcLAmKsPM1x6F1x7Y11necX0msVW4obXvkOdjDVUtr54ObT2V0EsV8En1jj
QjzVBxRLCf6k45MGooTk/jy9xhNNYyKAeCd7FpLg54/Oyh9+GxgM5MZECm6rlSmLBgbNBzjml4c4
FfLlORyqkV9FLUGaUlmMaPsZCAeeMd42XBzagLwA5XqBIWI/Hix7dXGciD4SYcb42jkkAMmyLfLP
Y2DqJKGalX+wRdru1A/QdjkSwigVPmfCLaEMhNzprfHipnuXoTnN61+wfXXjbWd2XSbERPpReVP3
eTWNk71a2BDEirw7nv5jgWp/duWoZqVM0Xd4co13Mm3zPv6rQCHv219oRvGSLR3AK9LYFRMUcmvp
kr886k1drFuMc9A//i5zrkMygpJFKJ+wUSHk38g7nZVIuF9CSugcFY9eOEzWla92GuOSX+V7BDSS
EvRHGstM1qX76K9Vio/CrqL0ZKLUpiFAAN5klaPOWtHxROVzeTfV+Dt6GBk3h9I2YchLsV+5p63B
IulISjmU9QexBOZd4PE+r9/yLqpTVvDGBIPzMpj4J5G3aoKe7ym1YQLXpMRe1eUv6P3WlyeJz3BN
r527ZBdtgy3QHrVT/OyK31S1oBzaAZrHJ0qm4HvgOlSgnAemO1CbHfzynVlXut5W1ER8xYTeVxrc
J/AOHSVIfxubjqDde8037zQOshCS43SnuRbYdNWLk5PtKP4Aq1dGgs4HKhFIlaCofF1D5OYAMg0g
S4IGLaEmXmA8hG5yM3cNRZSkjaw3PcH2VkSSZViS2NiVHukFaL1KvEVJ2BAvj2DcjBocWxyZh5LX
t/B/o7VLZ3aBO3nmcw53BCJtAj8mhoTVnawqvq5cut/gDtxDdn1ba769kvY84yRWIVEE8J7qg8WO
1XKFiccAeQ5DtD02DpS7+jyMpNQMDMsLo498R0mCJtC7J4PbKvFCooWfEbbydd8AlXhNzku/Hm59
I6Fu2dQ4mQEq5Cdnwx2jnoz/0F/kWeJGp4nAhYwNIwRcUGP9paRKPCzonhdtlOgLBTS6UqaqJslb
4DKqjyNuNs1ZbE4B0Zdo3bADauBcLZctH0s6C5+hct22dwYh/aSbA39t+UM7Nm7kVht/Gn4VK/Rg
7kt+DfFZRDkvQ+nJEdPrK15IWg3G8oitzYygOuTNWwBDspSQecgCysOcbqzZgHWyZuON6RzIG40+
yNsPyvSfrQ9ersZPHF6h50m7E07zM8Wfp8pwSJRqS1MfO/ucrj4+v9Atc2c+rxQYnKS1ZuP00t1s
VPwY8bwdq4vvEUEYNft2xhdWt2L1h8h/ow291ZRh7kkhFWAlaVcD40G/ncm5WzWpu/LCvxclgLpd
50XXBYgoUO/cp5b+a2WwZLpryrX286dIx+ITLeavyLS+iVZR5V/UUzZX0NF5/fIm2XIcoqVQ/kXI
De/eeklOicni+yar1ZuW5ybRfboD4nknVik7maR8eD3HayQhrJJ8D/GvJHiMhO0yKQYJslg4vwAs
e1DmcTkAM26SBZg6oEmTMoNBRznB6Nw+GicIpCV3AU2FVUOkVTy7yjm6pKdbayZq6+r+AAtgFhU8
RxNf+DcZ7P+qIyrF91sxZOL+KOtP/Fp0BXu+MBDy1aRQvjJeNdrGiDqO2dR0Zr/jgkJlXP5zX//h
EYzc3TLmcB0bLpfVqCpVV5XynRMdeNEvj9aSFCIp1HdT+8vS/zRoBfankj0hisMKlYymGO2iAdQk
RLgTVMf7wcMppzQp2Bgd8d+e+PspkVcIfov087DlFxPWEnBbgBXYD5G78TQNJhZTmHVWdqS9ogWf
Iok8vODNXyAtrKo1Kx9JzxcFLNU8Zl7SPjKM5o+IwJp8JECOWsaFiJZrYU8iJ1G603cNuu9PGwiv
Ktd/gxZz8gHYaXRGcxqhQrXnWgJn4mwpyrxU+hR5NoN59J0EyyURKMpkH8DqeVJLBI10QD4Ekuzz
zdVLKJqr020HH60UKuJbUE8ChTTj7byNXVgXdCifIJ/S0rmdCnUiASMfQBYSSYUCKJ4msnO909uU
/tBb+FhJt+rH3EZX3gYAaFN2U0tFIhIUFN3TGfo2SdgkD8DNfZbFghTFGTHLsbsC4Xeexy7N2xld
TA7k3SpGrLig32c5hNc3XedZsma+3RV8g+aKvFPAQks21MtoORMg83QgpppjSCLIWauk3ly6ucXk
sCQaUzwtLej/WqXA0stglAHyNXiUU1VDp23m2Gn+Mmo0NmP36tcu+LCKjCY9FWunFWKdJrKAGjRI
Jy21O9ri+lQ1REr6lG/Q8TuGczIbayj/NqaAbVVq8urYIrxoc/pCvDTKvNevXTpcmbPghZc8ct1e
g4uFMaL+MZ0N6W51+psv1aAvBcLk/5XbCycgWWZz/HHrzBNG7EaLiG+jDOaMvXymU4Z6mD9tpzpZ
q7vAQDoTzcBAJcViwu5czPHgBqRSvRPht1SSvppR+Ju8sLMyNf/Rxh9ZxERgfZHGovMvDMfpJXil
xVqpkOHfqBLroMTzOPNHjh7cVtqTAVRc2LXa64V8Pn6Vmzul2Yt8UyTAyyeoy282nESto2PlEaYz
m7WnSNXoRBL9kD/t7g2aqmNN5XX8AGiA4iRE14zW4J8DhL8IM7/QMtF8Ix/KJ0TQYeGAP5nkENtY
3BTnrZjNbnp++uZh2VEf4drNCQg6Nx1k0+BqRNHrSp8LzKHUmNAU1TJPUS4B7gx89XgLZPQ1tSjy
aWYC07Tux9j7XC9emv23taUUA0daic9mXMmI53Jc15D8UCn49jh75ZIpaJvZ2aU4SZKqWC4GdCj6
aymFFHmS31BDOZnCxSsYZwQbA/GULKsXokqKuqdCtMKhBctnSeNFUudOtNkiELfziTnU6RGPIbT1
dFYYNbRSYrR1zPloZoOfSPUZD35q7QS7V4702UuRBh2hyyZG8gZ5P1w9moZFtNBdFL2SVlT+V+tC
ZRNWzZFdEK18R8ctTvC4wKpQ74dhOATdl/vnPW8+4jMU768NZ2q1GHWmzcfeavK9BgwIiauWJBjT
mKeinc+JInNhulIgdMul+Kk4IqbUfJAFRzhV3FK9pacZ8ezGGxujGT3CoeeSbOUBJ2nhQJLtfnop
s4uvkeSkXqDjudIAqSN+0XaJsnl5HOI3t3emSO/EME44oidyUjOQgW363ykq+IEpdsMqacOZUAN9
xkksf1Pq1ZtUhFJ8BYweQTxJnIXzUmsrOnnKfrWv65MJw7C8iCp3zv8zxKxaBlAEVKF2d0ZuEQe1
oRACBlFpzaozZJe9Uc7k5Yq25TPm/jOaQmaY5nMm2VxCs0JYINGPCTe+4Cvq7/IEV75muOuFahBk
3aSBS0Nx6GQFS7+OE8nUzQXNRgmeNBTehyepK/jLB+K83Mkm8GReYKkslRxIT+Ml5/qiuXSeGhCC
uOdGh31sRIAJ9quyvCknKmuoZpfGW6BlwF4IHBfE03NHsY9HbF4NGb6qF2dmIblJNwZpFp244q06
GTIIGphcQ4mSKng23CZTM5KBbkkOHvUkcVbLuGlc+Cq0g0S83I5Fbdmgxwr8MyuUsHwBvORbSpzx
MUUnNEhLsDtQuHa/dyy9F5rk/v9M62F8wVmRcYoX5UTYJZwfA/cYp26GWyE4V6xFxh2YJGEiQ28V
csWMIvBOp3tfA7BgEaLgyeCZWZZYUqTqP43+ZtPJCDXKdcul70g6V/QT1AptsLDdEcg77i+KytM0
oqUoH+o8zcvFaMO2cs2vBAuo6MjmcR+mnSlEACrKxcN/PT23VdnyafmEB/fIw3fQWW3yVprIeJ7K
mf3wmY8mP3TvCScUNCrjrlxtKX27perR3Loj+8XFiMN7pi+67K7JH5XNqA4wKWXvieXkBfpx1zta
FKFDmxmygCNRhK3uS59GtC23A+TPpo7inw6IzezKGytHklNp2EF+cSq5/dAIsaC6axB9yHOnCoJj
tQIEyoqbGKjeTEaAxHl5w2TqAgBU3CMQhkwSIOXp5UO/7eIBRVDAi/9EjZ+kH16fzifjx/taCeYG
Eaigp0rdIOVCF3Ue4HrgmigslgYBYMrB5SK74ZMLEJxTNu0X+ZDr1nsX0X83u25kC2H9x3YxS/HT
Gv6BpknnbuXuNRfYsCcSkn2Ub2/RwDb7SLHydMvjnGfrdV4alhI9tQceOgkAophba/2RgvaSYKWZ
9448xWqMeyTUxZF/wk0FHdFo5L5oO4TB/Khzx1G+pQel4dmAOyma8heTNA+E/EelF+p3gHy0Xq+F
G4cH9FpyzIXdZa3+/Sg0me8o9iKVLxfG25K54DlaBiAd7co7g39Z+hHsXVil8wu6gZb/PQHRQb5t
SXNlFDj1WBppzYkvvWi+B5rtNkFKl0G1oZXHkwEokJF2QdIaDgPaVJb8MGw1d4Fa2cIgaRN/XIa4
R5DNmBnchp5Qr0mM8h+Ya2i6Wt2dI87kMG5MXppcwPlvCWX6yTnR5ECbwZSO+sqdWKclpk7p8x2i
qdgPVnMrbILXxbX8dUn/T76kLeuGUGZTRlzrNw7ixeIJUHJQCZL2xLkRRqpMbsQahLrS4HR3YrJO
01ocOsnldBVolQ1Q+SubIn46KGskOa6XjxkAHBFUIJ9DNvxlyEzZhUKD5Yfmstocwf6CTmC/mDxp
Rq91ZCLANrBTOvJEcn/uBqAKgCiigB9Xt0KlD+KbnmDu8VylSQIe/0pQmoqGaDsVWVYTwNTHt7XF
AvZxIGBwlEuhRoLatZ5JjgPXOKlpRbfDKfP0gm73NbJh4MtrzbmcYJW5XdwOh5PLxGwyJ5qeqYeO
bia/GRr8/i1JpUG65/O+jBN40VXX8NBxqOPD2sGXM7p3OuZReo7QjwjMoo8c3kC8ZzlsHUuzKlmu
1IhzDjYtoKRGISwNOozZIHm5/PKuL9AnZV8J2mpspL3S+TJ0jXJNY57OROW0NcT9sl8kOxdiNcVW
oReqMXNDDLA8IEFz4nAVn1UWMI7gGtv7U4bopG4ITeSO6/wvC2M6M7e9z/w2JX8jmozzg7fEAsc1
1WfRALf/n9NbVeLrAKJWQv0gB/gAzt8oTcqNLZiDOAUaXAnYCMqLyScEXkwmbllnN/h/9trhz10O
7m5C4bdfTcVK7ZHhaBhtXIM18nXqCGwQpR0SdatJIM0MEkqRDvMNKFPyMEfF6bhDKRHbDWxrSy/2
iz2QOR2KZ8/wTeMoIW5JNvBEnaxuDkobg39iY/SxYLXduJ732mvd8Aq07uu4inqAHigDgB7Gl7gk
B2l3Q3/QqPSmjLwe5UUgqHvx8KpbXBzxF52+L8I6/Lwwnuc54cpd4fl7qBtkEMe7NvCaYwRNcuOY
LQvNipOgB+hbZcx8bnF9LNG/0pRM5MmsgRtY2kGvTTFI1VZVvRN65IIpszPwtOWfgOQfy54fe4s9
z/xGhsfmWC02B4vFoR48SKTZOWEwKMWcgusLesEaTlmt/OKKKwafdyEQ3qTpaVWSxzuIQaQv0Sy7
wQLYdH1nq6pc6OcpOs+F840mTm/o3OVprYC2+T6aopI/33N0wMumVOwN66mKOf47+8b3nxqFxTki
4QoWcNFb37hEEUjWbbnc2BzEp1VCIf8cKWmoWa3CKwpZ5LtIuGe1UDQX/d5ILBbZ9E0mhFULcC2f
1gsLAKuoel7FoVm1g+mryL0DHIyxKtiJPjvgqfMYQKQtfmz8bEXlzg/OObPEAQ7m8E+zfyrNBQwv
+Gp1V1nvfZwflPiGDUwGuYsGVgVg95K9SegR4SnBd9pUm358OhMXv5Yp1eUj7NZ6KAvz8GHiYbUH
YXli+SQY7E8dEUCMLxy7lyQysbv02hIKnqXUtq73NZ94KBxjZz22Hy11K88AgfXApulEry9uXU3v
d9feEehUlbdfj29wH26N8VNx19NvooHkSm/qDS4bnGkktKMs7m9M/pZ5teHArywnOvW41B87O6aA
mAsa1oQwCEf40ni7moFMaiyANnMbeRwRyczT2T95wSa11l17r3jntqmwobwvIynej0o1D6i0RAir
8o4iM+tZapkJuWnQU2bHWwrOldJeSxt2t3R08X17y6bP9G1qffaBR4Ow4cyvFHhXbu6tg+3qQKa4
C8LI2/+3Jd0qScAz6HTd7vIlufyJyzyah/8WwjY30uu4v90y4e2i4pIPoTktZhuSUmSgicBMk5nq
okpSqQ9F8bBTUJb7m0e35eQfs9ujprP0Z/GIFfvBznl11c5aSbelecCrkkwrAluDAYcHs05C8R2I
/x89kmkMXe83i2s7SQ1Uzq9s8VDHLYW3Sgp/N/ZBnth1TB31Mz5v6UXHrw8MWOISvhnZS5NLif/7
Xh17K1+7V3C3Ke3s6QO9uU3NPP0QcndI0/gZkMVd9QXPEGCy9AwWsJLbm0UunYWas2jMPR4JsCIb
UOLbBh8UMqxTQl9eq/uLXafmgj4wrq5WtKuD0mgIrVqQbaHX7VmDT1CpvkjNP9bj3Dcyyq+C3KV5
w9DhzY2p9D4haXCDp7iFJwBWzIEVEYoVhabN73Fsfp1tAbsCfqXPxlsfTQhDz+Z4jq7wdTPV0pGq
NiDIClGE7Zbtql4pfrn3lMLPLL1jNm0NnXQcQhlb38zw4bb3UJU+cuFB/qbfP8rHHv1usssrba5c
29N83EC/96xX3Sjp5OIv9CLmO+CXrzSAbdHjFeUn0nkVpsScyO5ZICG0UHnp6cc/qCs4AN0ap2sU
cJotCwXzPHLFvVXAXYVxqIMmtTuo7ppxuCFBFfjGq0L2C8kelDcVtJ0OZZMUSxDAwo6m+00KpjBA
ScsTSZCwI6W0dBukV9wIPinHsGcvPSWDRR3ECbTRn2Jkj6oDjxwxlGfjYm8OGmsEPZOgrPX6bR5i
R6kMwlXqJbz7mtMcPzAzfhIqKG69ybkOZ+njgZIYrk9jek5DV+nwwwejTZ4b00mtMGyIySkGRgMu
EIB49pNUTf/wZDH9J/89sC8phJlibGzv++YcFNQybR1MapRpnPrETP3T7cxudmFbcVanfiCBvO4R
CcazIq/9r1Mz3z4RXwARs6PqfmOREoNOVQwUvIb1yGAwg35Nt+lkaDOF3zBs8Xx0PWmYzwR2Cv1Y
uhEcs07ZUjTbtcXt1+6POfm+OhXyzbtLHa0iG2zAJeP3wosJuMjP7CqPJSJ6hDCccMRBI/b+/ycT
BEScNEo3Mc9RuST3SRfaltULpevEz7KlHQ2o6LhASc1Cq7cfl1DzhGeAfttYuSaGbFur2Pr1uT4G
jqkExCCnq26Z26CCI0On4WffN6gfG9IKc9UNoUAGRZalYTiAb05AoJdrhHiu3pIoDfqiwT7SwEbk
+eJUUceuLfl34Ocgcbeqsek2JOP+H9KTbcHlHygjYDCz3DbpZskQfHo9dngwWmIBPEtHLCVNRqhx
K8jgDkW1I2r2B2OtAU2GpTy7Sa1XFiZTAW9avCpS10Nk09wEKAmcCLt5tK1LKjCaAsI0HKfKWBjU
CsHXBQq1m5bPDybaO+XHiarPF/qtJvxWNzbcXo7HAAkA82UlMhOz+0qfUUPxPObLF0AU1aiBwrBZ
uJES/Ww2fL/urw+FEVVPMJqUJoMPbMfP39axCYUQrr/FA6L2Z6A0yWjDcEqV2SD7PFNv5XMPa08x
wC3+QB4zRTbMXV0LCxGT6v2sDMToHvKXCZscrm2uN5FmS3LPcv4cwt9Ioax0UNCemjXJ+RCjIRa+
CSrveCiMCKFKAWoFzUuEkWizDjst7/m0DRvyuact4E2jOikDC+WL8pN+ph5paG7jGL7n9NdalCev
1wF05ycyayw6LwBenmqtafbIY3RjZQi0FJLDCV8PM897fG042ZWWm4mqfsxglWqekZoLrfFd37wM
rmPx4Y7NjYb+tEwNHYy1DbHKRXleyHkuagxL04hziznqMH5gadl3lw3QXfIVJ2fOxWG/vwejNDmB
gJVackZyJTvfAbMCOFrWdfAxO8qe9Bl0DvkxIHP6lTe0sS36Ti+cD8W9n3KZncArrQKYxtGBfbqa
GQaYtaUg3PiuVP61tp/CVTikHw0e2qq1F5QTSULE5hFy4YLw2fEhllVY/TUuZqEqCUWl2ZZd2eh1
Cz+q77A22hpBTyHgx9iqQn1G/iGpNe5mV/H7GQebu64WqoxDwC1ybNUErXFM5mWopCehEP1WsZZI
iN9omtP5rbtXsoYmA5nn5jqqmkWjJxPHrSfYYeA25II8l5DkOIycaGoav0CSbfWbobV5phQs4AUp
YbsgHY0LyyWb8i2zrbsSRNoVfEAdzeJKEdbe575OYn/q0NRbUcGCdMwDdd7DzeCF4NzxNAXj6iCh
0Z5kg9JLLGhJQYTTf6rt7FHrHpQDlJROV8QaH1u1OO5IxXAcFjJOJQrB/4eImzlI2FvEsJJYbiZL
ohYjEZSzQ81p419dczG1oiuYhFRzKl9FgaTj9tdKIltg3nuiJ5VIN0R+qvfU8VgpS/Y+codDlNn/
78KmuO2yVJJH35g24l/djtZyckj6mkpMRk/pNVi3rHxIwhfZRbJiXzZ0AdSaHatbDFrmBi8KmEjr
tnLRZDREUfpaADwRbaPRzlJjz2RiaUjQjkB4Dp44ibEaeZw/zkKPsDdlAo0kji7+eQOPHMGZkz6j
ntB54rVkcXuzTPHv7I3wlYTsJgg6WFa0bTndxbHevCTW7b1sMFk8kDpEnLvKdmdY95syGglPqed0
ANBXOJTqGA1lK47yTPEtU5kafIp+1NNFJPFk/sefhQfy3Y7xf7uCAfN/KjWHhW/T+VKz/GpwgsQS
k8El9HQ/lVv4Pq2M+AZeDbtP9uw/LICAteZV7e/HJioEbOlN6P0Mhp0ldOos5NXQNYKJjJ9beHTv
GRHKcG91slIfDwXP5NCICVsgucyEX1W0JHcD1n6RUfGRxt4+ORjphKL5ZCHjy75AWYHxKRqR/JHH
+9oezLnC46iKRSPjUxsgwpWm4v4Nfrm2ZagOEnR1u3ownCU1eUqQ299tAHzwz65g+xb5r1fiGlCn
rqyt/08Ws8DJcoV1at3aZv5oZiQeAwK4VAyylbPlh1rdQmcesZhm848KXQqkDNX4wgh/FQsNKnwW
P7ovW92pxxSjRLbvGytyD8N8NcnsFTK8XQvg2uOBeZmFGIFwFG9D3M91k4gO7MJ4mBRtRFCXloBx
VbfQfl8KOvpdZqntstCgfVkhDinYpFDTaag7c+IqbZiLUS50eqhaK8/qUwVSCmnPzDGPKneHWTB4
1ehAjxfQBG7VotkJkm9di4oizG2Vz3e6tXKeHtjY06dADC44w3S7IZTffIFDns164zfvNgCaUiNi
3xMWBAsfYs9vXl0lTJyJ3pmy1A9SCIFLw5/ywUK5mxn8BmWBQI2CEcQXFUpQ9I1OYJH6VMoHSK0v
gPNtaPFn0LodP71nk9YDSglSQ3zPwZgpued7H2FmmEGsvQgwfSZuQGUtPMvfDmIHGte+tBgnHnKQ
nGpwnF32o65N+1Hoxp6rkChw8d5Wp7d9NVXS3VPbWMj5UXEziAeNqYFJL7Up+MNCg66pa1B5Memm
RzTpKCGFAQfL+64Jp61+1IYiGSImBlnTjUuTaEzYmFlUIuuND97SP94XIonhvS/lsWN+R05Q0l9l
JxUZHt/4u8T2f7c6k8TVAj6yBHlmLbXOYpkweY9CwcUuqkaTnogANfpBYIQkLClhgL4G1JWNjaZh
UEaaB2uOOb/Pdmi8OScB0MaUtSwl2LQ1+96VROYPR+OKwK6NRfExF7/jRNSVxxERWKFPeMgor+NC
+e++nMNvH5uJ39PNrHUNz9Fhe+xQrPqDUjPHCl8oWBChKLq0AcbX9QyLGjNqZ0BP+Y2uYAKeyBc9
ihWQMjj93FgT6Ai5cG3g1wN3AHfoTNbZG1lvq33rpz3uGf02TNCjXmvD9xAVT23spuEbaoHiEHXj
vfb245+obAbbqBT5DIAooToJak+ZG+p9+yAnQ3jyNzqqQe9EQZg6Cuqx0u34u9+yAne5Gx3VKtc9
5lnXCopo//ql+wKcvbYxhL8V6HGoOnCd+ojT4LV/I/6tD6EUAHQUx6lOFFGbiBoU8+agkaQUnneS
yq/xKrMi70MEd8CThbAsAG4GIv4WIGPdZ1PsHF2E0ZXptGPAX/NILmGLcqtKes6s2dzeLCfxlTmu
+G3WDBUg2hLqMJRPCNi+1Jw51URVG0suP9fhl9pOHkBZRuHDN5vSv7LfEir+0wvueCp/OPiYqLwz
Je5ELTx6cV+JrQri8Pxs/d/7BBUVT1hCk9CZzkkFRZr5Q6zxK8U2kxtk2XZRBHjy2bMtHDfRv1qJ
Cs5crnMqH1KMKc0EHsA5JsxdGvYUhEVL9j6JGhdnfd9OK73LlXDzNebg/clNRgyMLBOpEmsmSpvB
LP3G8Cx/ZysdTJSVRglEJUGzxCq3VbwYDdJ+7hp4H3Te3NjPtgcSrmXbdOQdwr7P9sljFOJGp34X
JaubebmgF6jH3yKGFYA188bdNY9yk52yl927h4NoUO64duVYrE+qsE4vEwHMnmU+spfUXA44lNvv
svy2vIpFRbi86q/UY+YG+PTeXqv6qhjXLBeUheH3nlOOtCMI123MalVRBjItA8BCsV3MvzL0Ia6T
ZkOXATTx1N1wO0bRZrCJ52RO8Q/8Z1Pmz6XUH0Zs+G3fJTaWtHYMrwKGS1zkBLyrgSLuZekbQ2wg
nw5FEcyeXKB9/WANzztzFjFq5WXmDoJaK2B0d2ABZCYR/JJsaq38Tuf9WWDzPjJ1wJ+2bXTiwTDg
vVsuVZUGhGQvrj4uPNur96lF/KPu7NesxW5sEDco5QMf4oQvrRkUGQOkrxqt+gd5CBV52LAnjvaB
G7YkLU0oslGwsCuS7akFGdXxkVjuggZwMwoKyQjqQ5RPvugc0RFo0hnBjDGVWkNX86ERH/dQiaNj
7JAEOL10eY7EW8dXqesm4K2PugTadt8wLbbF8eq23oTd65qyhv0j4kesYNRUiy0OzM5VMeOGQacx
IfYdC0J17QS/gp49A7eQ24xtxdb5EDolTVWIQV4hKw4VsfUtW/lC+PAJeR30pzadAtPVowjHtDEU
944AmvPoFMZ5eaIX9uDUjsViqDiGi5+4zGq1EXWY2Qoi8aiQZWESUxIYNtD1F2W4WjPDsHP/Ojrx
VGACRZqeF6eq8DVjugDBjxR1SAYKtbKu+z7wm/yLOCt4IIt0m8vMgUjOrkREOx9DK8n+q+dLu9S7
NvFigXoc025iyYnuNBUXtPKyero98dG/XbELC/rgmSw1Ebh1oECQVAHdud4QDPJWlOqb9QKzeFVl
1/dbVV5fZchaBnllGVWXa/u8B+VsAcvyAoOP8nbmWwncS+AOhr8hezhUrZPWHDZeVC0E3SieM/rq
z/ooyAJVy1BYMReIzYVMezNMZKjX3zyYDQS0Ie5ORtexgQnadxKRtxXBH6fTgQwamTanSMNMn5bp
AVnS60n808xQA+KcU9S424EX6BvHFFWS205de5xcinMxlAJFNaRevQL65DNxGQA8NZtRkWWP59bd
gg+7iSPlXmQ7qLwbCGZbbTCZIsda9Et+jvFV9HRVNSiqJxVARwfsZ0sjTweBj8DJ1wU6zK+BpBf4
AveP9D1/Tv0Xu8KAVzXstKSiKZGumTxwi9dPD4o6+ZKMxuj03CqfLejQpWcOVflFZxwRH8zl9P4c
AXiav+g1my+PDlzIm3lcgJ3ZApUuohtvT4N1toCYwSFN9WXPzxpR5DhNCy3GZR8rVz6+qIj9Rxhr
2pIIkF+HGmtNb8IEnW1uTs7ckL1uNVFgn7RMKi5s6dxx8Indx2FUwOGl4bc3N4DCU4n4gLof/vSg
nZJT6dYPlAF2M49sULTejMB/gN+SaSm5U/HXJAm1H5t1pXp0f1l1UWTuZ2D2/Jqj1qYa9xFtArAG
wB+wyLgQJSg2mm57Y8rqoJIwsrrqx4H3GigQcDfKXTNb+7jhtMwZCsF9jmA9G2mIscIwhMqJy0+q
TiM1PbsMCavtULe5rGjgJYp0SeNLKj0pmmto8vtGXPEsrsMvBwz66X9QpKGPiPpNNMQSgVP1vXC+
8RON8WSxocmoD2H4Cx3CR2AR5SqLfmxxDCEICpiANjGZmoeabdH0W3aVE0Vva2KsVS/JD7N6LMRh
xFyLweveeW69ca5pSdRJ5PM63S2M1dcjLhEVZW2VYtNXPMTEX86MdYIt7xD7BU4UG/V6Gw2WTbVb
3PQNtfp9xSmWqZXOYreJ/RIrPYB3HS4reQ2PoFvIrZDuu+YAdLKOoae7Dxu29kBDidYi3lFfiVKG
DpcpKpRugURMwnbJHRt/xJytC+7/8xT0BWXIATlmB6zObKjKttff5zddrgyarUUGnA+B7hajUFIb
Ubil+Zq1+KwsfjyvRgi2n3Tl889UYPNkLXUgmtpArT4k2ce2wg043lug+TTpImDC/73w96tY/jGg
MV6pL8Vc6WIfT5B7hDUoT3+2Zh1fxN0E3p1BzDEuGyfSrhQQFG+05dDJWANKlBI4Dh6IOBYfkWRJ
9Xl3ccAkplwN8xs30ZYSm1B1FsUoP0TG1fLwEcuICaHoZRyNTo31f72MbDZs3glxNWUqnhrUxufX
AZ7EPxyQ9WQlXbpVVnHR9f6t2Xs6wnVBAgVUHMwFvF3OP/ITdi7VAsihVJ1pRVs2FbuHV+HJ3OOV
lVh61C4RU0OI2nIFUZoSHNO0nXGyIANNQQjlFB7JWhptVxoKfRe/vIsViDuE7z3MvFonwuSabhia
Day05Q5s+RtgjoRxd4JXSaDpaThC3DKwv54hq222S3zpQpj8K4RYHciMDJJZpIrYfTAHX7jMIZ1H
J+UHPvFeV4jiRfnHvqsRthZBL836TGHsEYhx3+5kvRiFCnfdmn0zzorKWwRR4uMSZizndDoZHMfp
XSwyUKJOfCBg3dbLasT3Od7jD8m23YcmKiYKHt5RURQ615aPCZU8z9hYh+KxdGNJa7n4ERDkx+rH
/KeCEMLfESRE8+0+OYlLcEB2K4smKgfzOQYnVnTstHApPs5qmYXtyu2Gc9Z3aXN4yH+0v2V5r4Xt
hlP7vDbnoplL0D5KIROkH9ObxI/rUZEX0hiNkX/XBanyUs9w7e53kOLPBTi4Jh0xFdcq1HM7lEoN
0BB2XcvLSbFHSjzZ92RvaaisJBZ+f7KSsQR0XAuNPIDNqsmVlr+ZhplcsIOIHATwBWIcsZx/ZIUP
EuyQ61lucuw9gu8o/8n24wu+e60CsZGy9OU7AQhxgB6gvg+EBVHscvVGHrMNrfWvyX7wPn3V72xY
s8qEFKwu4XmMk1NG+HnaxURfEn+CRJuRXDs52XkAtR4p147sqtcHrSns+IOXwVuYwU76Y3z9FQM7
r3QRLPorflk81dVJVy4WswKEEObPh38wP11wYxsmRrBbIsPqqY63jxICh8yiAMb0ftol3qb5JXge
v8c1PZclNMODm8l4cV5Be+M123hUv4P8jgj49EVAqy+uOyfJDSYzX9rLHOljFN9UNUMyP8ucRZ8+
F/WeCK5BXvm/12b0We+RY9CCqyQXa/aF9z6iPWptOjHdLcd/AejC3uwRo4+3gVt42cqeYsCMAT0A
nZkmeTf76XcbApU4X+IJSwZi3enDGiZuV8b8xXrxzjrIs4otF4esnT9I5aBwRz5DSK1hVLGIRIin
9vmE0NhnpAIKDhxtk6LIDE5CcybGx3ffZbsVmceJaw1MywouJ/fx67RqdJQGAkDq7ovR5rGYWqwZ
1X09eLpgG5M5RCDSYMnFl8wH7oazxYnzR2oXAmYnAgGVPYNANMmB6X3IWy3wp2qDNuZRzrNO1yzG
UyxAbPYHHYfZx9IELuoY5vxEnoUIU/ApWnktPdUjURundglAYGgYiFn5OfRV/ZdVE3+6BsSuZFa/
0WPkRtaEJVz2jqlHsj3obAgVyJCoe4hqeAV3YZBQBwhOor45xgrZTIBB9kmZ465pLXRhY//Hi9RS
0gJeRA4dgrgUgrlOW+sXPWXb4jvFHqljFLTvMpEpNKILJlU4vEOc6TBQ6fd+1lGeKcgVxS1xwL37
e5/uExw+DXVrAB8vjU/tdo3On5vDffDTVXjvn4FRU/En8ax4HuY2dO/uLg932LJgKhhfyotjqILP
wh4ugsNFoU5wlwTtOVmKiHLmi6Bydhqgk0RHe0m9T26MHGub8Meq4gShdQgsCt3hGI1jC10t0Sn6
TTyl/CPd7T4O9UqGU2crB0q1gH0B6OvWdO+e6Wj7dlfUXa0OtkMl1WnLtyymrdfl3PeHXeg5xOyl
uCALzjh149XFYDSATprB0mzEwwB6hTyXVrF7aRQacqfVVfY8d+KwQ9EgNvwCbYC4bq0IkeF5Oe+r
CHAblGHItYnHUix1eL8hyNzyZXYDiHS2qBlPJHXPBqCmcaTuHbQAEy8SpUlG0qHQ4oHynO9Fk9N1
jnYvYsmZJtZRN4OmUlFlAuxUZKP1DK6DG2zCJeL5yLnSsFmy9uEYauQRuk/+1xv3xUed6As/pD9G
V1UTaZCa2r18Q//+yPtSiR8Q8p2FT45FYmFAUwovyVYuXNjHca6ThWVTuvE2T5/ZDU0/8pdlotQW
S5GfkiW+wRKfv0rg2WRj0FfgoNyD9titY/jZEz0h2xi24s7+n/MKJdnFxKbcI9BkyS/SCie7hCFw
8Ue2LvfpBlwqtFt6cqbFeV/FHeT9y62prPt0UzeUHy++K6PZzA9qJqHwzWyf49yIzPEZX85cNG50
wJhEQto/tHi4N5fDdva71jIZPLmqiCeHLNAKynDdnPbEjVbACqA+63B9cHYKuVcb+RhA2fdP2kSm
JnH9pt5WY0gi7tLGgHUTvWPRPlTfpefSmBtVSCYhSskStR1JVB4vrgte7GHAms7s0dV1EkmkpzqP
DbPLWDF9yXk2j7INT/G3mh55oOlrmc1kDYSqaOwLhEbrRHBBHiTmFz8LPuo7NDwM53txa9X7+8h8
ZHgrgz10THbdwl/6QBBWueu4on3oV23KzrKGNM3XJ3cs4DJlVdUDn6Ohax+JFpPGPBU1ipI/GtLt
FS5hjb4PjW+O7aKM96oAbxRsu9/222e8HBafPdKEgzuTBAbN7CkTad57QDHlQ0Sfgd0X1LbbmBen
Cu8vcnDx+JVdWq/jHsCjcj6myueA3SdrfYsU3el6bWX2BbavfEi08ftTjIYCuJ/uygBQD3ILUS56
ZzYlwPD0r5LzDQes4JXfjDzUzLNoyA0U5CFLv5Un0zgf5nPKubIc/5ap6oCs9LDndg1DmwMfnS7/
zLduVRAp7DqMxO05DqTKdKhZKfP6xyT3IbBQKMCPnjSDV9MldNryfC+Nir06Hhdl69brJMy+Munv
epRxLru/B9PZz6NuYGy4loXbYbq0pXCjYyuMH8goNtSN7OjKBBsTVjGj7soKMgnIRfrtMhtqovmm
vjIS3E0drSfcU/VeMFzzVmKizuq2mf0PKbiyTuzEugqKAL5MdX45fY1P5pstzt149d9djrz976Xu
4Z74J8A+HNscpnaxpyN1YqkRPOu/NzEzinsdk1cfTHkdvKwGIOIcuMNhqx/aZ3BiQdxHwCFvhsAa
NUrJtmF68fveZKQRYOZQ+QhuBIChbTxPCUJ5SRpZPPFeamPuMxXh2BFzBwK7ss9/OCIh4XZZWg/4
A55ZPGhowm8hBGUZV8EId4tYK+nQYe16x6i6V4jQfngtqVFHwylfk64bjGzvX10bvgdFPK1OXiAF
VU/KWHIJPhZ8QvAJoRuFzqbpDOqKlcHHVZ8TOQT7vi4aJhZqNO8D691EF3hELWC5tnhAStbJlVE2
llIp5EuoZhoi5nA6Y3xLJJgzdC2MGCaJelD8gfTDBh/ADK056e99JyfDM09vpJNK2GtNgIeTjiUz
ihZSSeHtp6tHz2QpEkrfH+UttZHmhJBki41f1D9SZUbspOPt2zF+jJremTPTWqu/VQWHWJusvV+6
E/wRlBZF9LkkpV7A3a4vqruTLCb/W4mtlLBuCnCrKYuNZhopUWn8htDzEQBy4UUQBrL4abEdRfa1
3KPcyb+/pmH9GcYBZvyDCBnCO4Z6kzIl6Tgms4sBZdzI09E3hO1R8V9U4iqKMk58k1vWygUnX+EH
cx3nbXrvWh10N2eZhmjONzjroR8CSBfX517l4hhft1281N84Fy7QIzwCGi+sPn8C9VRgn9gkum7n
nTcBwmUrdb91kexJdnxdArY7bSnvkqoGjxq8AORoRArBDktWwyaagDF2OFXpe16Xnbzy3l+04OEw
MZyXpLoZUskb1DBmRADlxk+picoadjMcHZVeXoUY9rME948/IxryFZyaz4ycSL5sfbmd5h9h3XI7
8KUQKhujjnXGNyUDi8PbmSGGfMUITXSJt7iU13eyYYFtGvNx2ajboKdBvXZC+CXft/L1X23GovRi
XeHSeyFfDsSH46a7Ec6FOcCbY457gDgy7PMRMKADzaGnBDmSNANLKwgF8xkrQU44QIwzzGz5jt4T
zHkeVgmrfHLfhjgeMgJs7SScU7a4waJXc4/DfGaquTmtxbLLtC3gnjffDDlQW6Cdy6hziEWSA+Gk
eYzcZIQ2Yk4KRi4c6r54+bHeAQGxwbPauycxaJfu9+kT1fC8ZF8RUtip5ftIreiyq0SFJOxqUcj4
htnnYNc6/D4FIEx7uyj8ri44lGWhTHVYDQyIrPl3rlrj4s0+m4FROptpJj2zwNq/XHsKClVynIY0
U9Pom7bCtgq+luIgzwebGLyYOzYWjxp9JKvuK6Kw+LSEFfIam9jil/imOIvyxebeM14i4DUojDrC
8AKKeWvOGn56Hxy3as3ICsJT5IabEyCZXBgb66OYCp6EpdXwF/KF6R3FNDkn2Mc5wOm9mOl9ewaV
lYLgfY/TcgMAP9lBRxruoNQNCdUJhETy8FKCyYEOQotFpjvsZnhxqz4oUWLh5ipHe8a48GbQHQcV
+AmXGvsgNa9bO6QXIMOC2+MJC3KWcQ0EjelL4rITcsKNl8dhtzOipRGkqFdyNr06vN9P4Yp2ff02
WgzfBDzexONAGzWZSLxhXDy8fmAmMxIX0M6fMdHJ/HYJ7cVLO0z3yJ/XpegExx47SXKXp2MYEoCm
nKp+RUrVJ1XXkLYBOA8uwHapYNXsYQeFn/nzMuqx/qV9kEWW2+MpQmb8NgRqGpdjfnMszRpPcOZb
XFqePKS3laTE/rfJd88vjdlM/YW0MPcNDE7MmjukG8hoog1pwLKff5Y0lMac/TQm7ARxvF5Q1BVw
QJ7tCGkMvHyCtW1a+p1Unrn45MJiKQ+MIbPapAqLefeKTDm386feGH5FCmZjlQUx2esjSPt1GRs3
Yg7Pa0hFmRleNwf9bnXkBsJx8yui3/e5YTUtKAhmUYlUYJ7Q434smjgb/W8eiDwfaSMC2hMQa5hZ
poZtmT+TWTIyCcbLHpyrOa2rv6MH6ovQvta0EdcgoHPHxSwLDoldaTPzW+52arc4F29ArnFKL/fg
WTWVmgxCaPfgxIVy0Oi/zrivkrW5wTpehQ1VQeC895YTN7D8tLyTQyn8bE6/48kBc1DOh+UH4OmJ
/iKrWC6B98xLw/ETAiCAUMbxFWRpCP9Xcm/MPPTMfjVlcJ3RFE9vuRfhTkSZzySvhS3PFcuNv66l
C/0ucd6jVZ3r4wIHBXQDSJPsLzDzV86czpH0z05J1d4E7Y3Qzy4dulQtQRSz0fAzU3rlzXSSBFJn
kahNPqiKkh4eX2z22dQj3RBSOpLANPVsMRcKhiMP0y8xxo8o1GjhOlwGAVy+mdSM1ulpIf20elNJ
+JnYwB87jFx+1rh1IOazFOPYdv9RkPrEfTWJk+KmdIjkx1O01sbAg8E7EYEKXTVZ350tjNHiwoIv
lvqgGGARr6hVFNVHUxZeqDttYqy+Wt/ADXLXms656lXXbL5uTHGgYoGmMYdn4XPuzX8ILAS/3az7
A/AtaozO2h8vzsyWDSU9aB6MLOPNk2svPKk2DOEJJ2+vTJykGHWyetaY3QFWhBGBj+AJOWtN+0w2
NPu8eTKfxob7IjvfzVc71WJIXCA7DmfrRm1CCYmnz64/hRq2yfrVlmZ/aQd85ELbv6SOEAuj8/I8
x28tQz+WQ89ueUIxL28pjZUET/6O3S92fHzFhH8prR/b8ust+ShtSf5ZTw1mqHfmJThAQ/0ocVIB
GYG5fZgK8XkWQrG0p4GlyhGZzVRze5de9nmEe/7psDuasmrLAeRmM+Jtgf6QtxksFRbjjrf3rngw
hfwYfU74IacEv6SGqnviT7BN7gVHx1eCUT05/m7FigxtHFJ0sqs8vm9kerSY2qBHri8CwgbY+rv1
sOE2evdXeFXVcVVjBvvN+90J6PYpR9OsEVlRjhKA5Un/hFOWSnfZPirAAqf+Tvyi043k+aocVxkW
G0fWWg+8sJiBO46lwaUIXa+ObjcYc2yTqLVMu1gq1Em4HyPXAAAXad4yLwuPhcgcuJbKsksr4ptb
fv/+pcNsYdH7UHsmteLLsSYfHoqhXR2A4Am2WsOwM9izzWU7k4fgOCJP2c2RtpBqD3NUI+lc5Y+Z
yF5itBLi4MkvrSyTeJjMmcH4z5WKOUB+6pp0nkWnxllPHWt0KWSUFiEZs7BAFseCsZMCmS0ZSkZa
nb70hBgdtZKZ7lY8aoYWIwQyZvRowG3sxU3nZxHsb2jAfsbAIfZIHnj7tKlr/AhlDfaoeLkMPrfg
MjNf7ZML5hT5WwBy9YN2lrL2eN2SMx/U/099weuofzV3iRBhNMigiDX1B/E8wHvV9yB7SuEOVxic
tkgF0epFRJCFQzAat3Ujp32Bdq+xNLMZi23Mt3K381kdB2XK+qSVACNovOKR1nM6a293UYy85EUm
FzSa6CGmON4HOMklfBbqRkq75P20Gomvz+q7kFnauNc+KeIL5MPbCbSVzKPb3I1qW91sO2em1wUA
6ten0iePu7xGfO8pTWechjZ/EAmZqYif2fvpV0IOGl3VDOrG6taSBEKYDW2ZFU/qJfkJz1LHUGxX
AaXtcxYzCztrE5DEUqLorsk/ERH0I+6WcYuWqmKcFIx0h75zv1/7TgKA2mdnbaZBeGb+UZWfTh9v
LjmoiaZ2JgVA4vnT999q6zVkhhUaMp3OUJWvdcbfz/EWB8rl4mO4ZsUEjD/W23oMLvGpOm8eiZ+T
wzdycd1cKPFWzgXy+3BJdCLtrWwUTIrZ56vmVIoRWRYoshbnqRQbtQJ8pFbxX3UW1/vsroB6Zgtg
uZkWCJl3fE/slKvLaSPGvAsQpl8xe3Jf4m0jqoyAr1enn90yw7rt3fGUn+R50/5nbxjbVjRngQG4
XRgel5y8tHsDcJVn7WS6KfjojbbvEv+4kVBejSoH1SWKxJH5HYpGFaUXk3z6ka9YMkOAgwAKDoER
dYu/eb8jUeVhJaChEexwMTM1MPts4x9vgcOz98q2e+EcWZ8MMGoLl+Nj8LfjHGqyy7OJQg3Z+XqS
NfN6Ljw6LL93aFFEohtu3KH/7tKLIj95dYEc9gyJVlUtIlUPAayH4xhxx5hizicfdkPuJYr63ptM
S+lCNvsGeGjLPfqM+t/1gWdKa8hA48k/vY8CrZisfyjdMNpiCMBAftoC9ThzcNpW71AWEZpD4kEA
ADJPx2pxEJcXKrRnfKGxu/yfWcZR77gvjiHojaLVP2ziQv770/kaWg8+BnrGf4xtGVctAHiS3DG0
54L45X7FX6cKrVF8OGb8NDdeJx4sNKVn7iIzFmo67feI8xV0dVY7gBJs+Ig9+vf0rjSUSR7HZVQR
Vkt+i2sIzQAdDinxTvUtOUdnd9KwbiaifBO8ccxVdlPszKdtgP+NPBLcFYFtaud6ptLN4oChZJhX
dOZVAUPn2zFg8IDcuWZZTi7wD/DgINYfgA/e922RFDRxKgjhCX3dnadJw89XP/HjyKmqwrePX8ew
QMA3XIQxgjfvLkGVn9ixl3wwea52y4jOPHv8QCNLNYRE+pQYjzmN+quEQ6S9tgX5sNjH0O7olNVG
k5iTUC+S+S5xUzkRhHWJ75kIsmSWSAE8UCbIAbPF40hXntOE70BFurxLWv866WcG/YXrpZX5AuNT
FmUIpwWejm5xnp6ov1xRfVRYLVo/Zk14CQ+AOY/yVIi+yaBss/t1SNG339xW1+WZrjSTxxlRIJ2U
8RG+BoINgY2JV1e/V1aUFdGBqeSKiCtyFDXMP0cHEsiH7EIXKI6CZV2mjxPfSr/yBw7q1bgeMWWX
BawOuCvxK0zXd3zQj2iH96lMQ3fJ51t0j6VK9/FOrPz/jAFAl8GR4WkCE3T0F1VL2K5TcIEmo/AM
/wynp440sy2gLjy1PLCrQ5dyGaY1nh3qRuchsF6FeayBYV7V4vSIMO3Z9jhKP+u+jjOTQ+7nkPJQ
5vmmkSIek6XeDhFguGbLI+ND5wCtOuQfgjDDVVMmbCY9N/cA7N6tOBiFiSb5Zw7CxBeuNZRokbot
xlTdi0MxvVo8ZacFV+d3AQhu0dHLquiJktRpZnraLYzgZm1Ux6Adl/Qxoj3R9uTZAMwNzG3kn0Ua
YAMyOy6O7ae1JSWTetJJOXpZBoYA+X6xeaV7l9UAMUQC/XDLC/ved3dMCpqyTU58vHa6E1GdlV/J
myVAhcNQHHhNbownh6Cd/femImXpMav+M6/3M/X/Ul/n1KqN41CgGS5SlYB21HGgiURmR6hfYeEy
cpuCAbXzZxso77i1YktArQ76mH3tuDnes9yQGXaKbeyj50mduznPzu9jlDBb4VCOIjtTu6ktLY8D
x20+r/oOyIcanWFG+/DjABg7eTNOnT6AGNt9p79fdTMEwTW5RfpXouJKRrviUKhRpL7jl3Il5r3h
WpIw54Cln7mnyEOO9GupQ+fZIVWgAP/ZkwqxAOWt9iNQ0qGORG6T2KEteU7zt6k5bT3wOjwcGfEJ
4Uy4jWyEq0Ytgw1x6VB7ElCwoYpaYdeXyBdtcbo+VEGYpHisa6iZND0IbvJ+vOvwZo93tXUTdmy9
tU6ACIgBZzB9oFKsy18ah9lhbLKDuK+xebFudegWSHLHxb/Y5Kgp9Xtndia8Frydp8pePVcl8//1
Y7Lio/iicXJoTPggZzQPm+MdwRVJ49J74pcDPJHX3JfLwp5HepToDbKcn/+MOLKEbwrBckaGmhTz
c5TA3yJ4dgIKuQjEaamZ5TgHKA3TH4SwljZi6OvqFZ6O6oM+K+QhhLjaChK+olc9NaiZQ5ITcbo5
m+uOb6o1dFQJK7a9KSm8eRS9vqwtsBDkls4H4xV3iY7V+wFXmowXp8X0xQRe5uQrAZypfoRjVj8U
saUXSPnj0jK9GAd97G3Iv1rGFdAXojSP4wlLyVfRZOddpaCffWx4N6X+T2cQrUKesWp69lKOJVnz
WWxKJbhcWxmqsPb7DkAun26SZIxKv2FSFIXhNt9e/1j7tPa0IVb1rNWySVu4FQ0e37hifMFsSidp
Xc8WmpT6dzTmljjUcvAeBlVRpJfXEdLjXz7YwN94ceK7ONZVJqsKXXce99IiQBZ8AzVmfVS0dFO7
SEBsjE7xEBkpGuGGZO7xESUWwX3/ApjLG99JKVSG3+HSZWatS6undFeIY1vXdNTwSiTH3gD+u971
XtIR/AjPfH2N8GLv7drTC7j/VQRVuPuExfJ1TweiJ5yA+ISpY0GNyazUCDPswD1TxeCxjlvC0Lh7
Zg+bR8q4NsT3l6MQP3/yfaN6nZYVRT8IwOK9622r6d0vbYVFNq2O99az5N+Kta12KhaIY3PxFoLT
Bd+KO+f2LK7d2csRbfELUDI3mGsnzmS/+tOtKYe8HKtb3wpRnfNywSQT9NaMzbUePrxK3S9c/Vid
Kxi2H8UH/h8XPlJGkB24y1hlrMHCb3XaLTOy8HqyK/KA3XZUl3kpaQp7Pp1wsDJtJQoXSM4bbGsx
AsPcCie+nZuE9c1yQpdcIF076dxf01yHWT05xJPiauUbl0mpZHsNoPYfQ79BF/2Zf2DTWpASg0cm
Sf975yzcM+caEBUfWKFtsEK/p4pJ7ohMTeP6m54jpeBE7EN7LOxx7Pi2C87JNfMZarhT0YLLXV/E
XQCphCLAdxlVL+13YxD94IWq+pAYdnPpA5icT+fFvu1hoGMYH0JYUU4fbINcTgcF12FVfCvmp0tJ
xsy/kx4YErjCDdy/UUdfLDeCJZIBspDMlP2UwdfZDkXlA5xSyGEvgSmgGLIppN3Sb6cDWNnCd0SM
X67xFqgNiy0urUZqBAHq1M23UkLUNx0HKc/7lvhsxlmLAYJqQPl7rREWPdbbNm2M+MrSr0lmgAJ5
UEfJQfF3E13FRzeWSuYx1ujPx0sqhS2zqqaoh9jlkbzowZLqYiOqe3D2VApEDM488yl18kVis7ZW
1q6b0kwJTulrVVdAEtWbXEusH43HR5u8cT3K7xEeyx1OGraKR9DzeJsDC1DRrJPjIZmnClmM48lp
/IEIyap8yv1qA5jKIrldQ3VzayUaG4HcdWVn5TrmCq6v86LNhh6ikCxx02ULlhjsB213HFb6HIy1
KHfw84LerS9usUlUixBYTfyASVr0eh6LCwM6WrDVY3yqgdhhb1Apiyiz4mLxacHcHNkFl35evVme
duYAEGfz5Q0o779BSc7W3BtSTRKRcj8wapBgs+7gIeJdXA9FUweROWl1qFb9P6FE8efOG4XcFcIF
U8grM95crOfq7OuKGoGmN7N7ZM6BjkJBFNzP/ITzQzaUsqnaHjU/z9rGOCQX47d8n4/zpgKJCMCh
CzK85dG0VytWl90pG9aZZXbAjfhqfoPMLa2DgJDp8OzEw12WJvTRhA/Ls0lBacK3VlbWB3/CsiG/
bTLD1KHSiVCl1jOIM3EvNp18KVTzTysw+BrM6lhu/jusTZlL36sda+5APB0X2AvpWHJoIsTc/JE2
aKs5s1gB8EdxbAgtRyc5jKcjHLV5TZUo2H/4J2cCNlMSmpuYvrq9uL8Cop9mMwLaeVswats1M/q0
xq+gcM931Db9S2HBZyLECPmaU8xa8ATBI/xR6Cid5yN/w7/ElLzDnjrc0x7X+RXgsPNxg80rNvEE
0F+CIK1i93+2KOe15zXh4I4SDonSh15RYCbQw19hGtsVXbv/fbZ6EEDxTeCAx0WJTSKMu0FpkzEa
aWaE70EsDwQZbHd/ku3Xyg59DerRGoOW6chHVehsj65XDR49dbG1dvdH/RiZXX1HsDjdRn+Nq+Rp
cBSm3dphMdGyre+i2ZtxBVdSaxl6rW/pnEsIHxplGfd/Ox5bBK3E7v8gQkpsg0MnqH+E7CD5eU35
au7kbVjG90VhvahSvhY1ktsb73fNFtz06h311Sq0nRX2ZFOO51LFWj/knkpz6ElsufV39halPGfm
FDwc8I0pjymShZWX2HI/cfIufLo/Gt4aQsDlmmeQMrYy/pK31CutKHSi8AD/Kt993Pt1nzBwUgef
JZYr5rdwY3fJiGFwTUyP1En0KJd4pNux3+y+kLT5FRVrG3UrCdMH1cirEVfFWd4rxPBl3hoHD3cd
dw0uaVn4pnlO7Vgxndxq+4UJabUFTodir3xVDhc8u59zv3rakGEVHcYag93N75+5+bbsimxX05XO
FwU2wEMQY6yyGEgRdd6m0B/njonFxJ/IC2Qa1iPKZk6IDyYZt4dtCIqatrWN06VokMSh6jjmjZas
8DJr/5LEKOpQOoeedadYC4Ru3nuznO73zenTPY6cfEohQgT5DJQDfEb/ZInXbW3Y38clahlfM8Ne
roWY6t+eSpcHjfx+tHxp2uhMXAoRxPDagQr7gRf3OCKTUBWnzrvzc8S2ilsm0bjsKwuVJeA1lbwo
IAXjYY5EeUYByjL8pySn4aTC+m58w7YpxCEfwMGjG972eO1zQ2mWLHujLVWQ6SOnr1aFDEfZel24
nT0Op/GEJO8P6KD9cVTrAdIiQh9emVELp1Wuct2YtvosFlMgdfd/7QL9q95hP1nZfXlqDj5SMPOl
9jpMC4li8CQkjNXr4w+begdJcERBFbGmGQfgW4PxIapxX3xoUAb8LGYBplnEw2o7kICDZBoOjPSv
j/3QPSRZZcwgHoQbUjQA8BLTiXFuxxNrLuQrEMNx1Ooglx8pgt7/R1KRHyecPU5qjMjSM258stHV
3IK4uLu1KgK5YgWFzZmWrdJXVyP6lkl3m+FXdvjOrxR3JHOr85A++1GOrfLEmUfBtRdLcmb+lrG1
jGtEp+OMMj3VkEZBAlGwFhKszPzRob5CUEp/Dt+i6BUyOhwrHBLAnjTFoIEY/Owo7LUB1L2hlkG+
wJr5aiSxpDqA4/Wrl+YUwfX7HesAgRuaQkF5WZtibeAIyOVBnjl6SWEV28Nb06328Lp7TcSA6qnN
RpeKF6UlysyYZWzgCCFylE6N3sDIAT3DP+FCKK7yYPFmwAn80FVViT7mNLh1b6s2UAMruH9rwte+
ZUXIMuZMP8ZHWMWkRICOrD2EbT8mw3KpYm5dnwzMUVLpKzYqb5OdWgCt3yYVx3ur+D5ps4VbSpl9
Bg/YLU2FWAwZXZV9Ykd6gebqEBh/DfkSjMr6YTVKZR+AO3EKu8kH508clnP2uWetgpGJqu3SUK0W
3j/0RsUqpszR8e55q6ijcwJURxVUeSmR3W4MuTjnvP6whurDEMzOo3GDTs0TTGdb/1bDbqftPVqb
pmilYAdEItPxsY+qEHscLaE7818nT5wt9998GrpyZvPdcG9V7PQWQQYmcG1b3qvUVcyUFIkQNMgm
FKJswhFApLEsw2OXVDDeHlU7HQWNMtQuzAs2N93/1xlrpeSdd4HRBQoRcj19genUE6PvOZwkw/PE
HnzL/dUnpY1/y1L4BJroNIeO0XlpqBFXzV0fFMeLgYeQ5fcFa+4YGuoVPxHlGu1f0O4Kti/Wk+OH
j9rXaFcJzXVuzQquGQtNc8EMMfH2BEHVh31CMfEx6Nu99pV8cUbQL8NlL2VVxNpSHOuiQSjwFir4
sr25izpGFBHbV02+FM4pxhEYWHf7gdh8bYR7XPYbt1TbNL/T4/C8gpXYFwFfxAmH+jXmQRhr4G7A
JcDT1fa3m0vyc94kE30EEineUr7XLcSugUGEe9M6iM+nulXmhWDoWi0ns5j4NBdUpQz5D0xd1aIo
HaJ0390DqYvndIQm4ovJwUdz5mRa8cXVFBFr7i1buufL2v1scqz3eU+krFFXmdW+amCmHuxdJATL
HBmt0ADP0qt4wJjtfsQmLeqpGKH0wBevHD2p/rAVAGV1UmDGIn22Nmj3YIlD9tbndksOA4LUYGap
aB6+TJbBpMEaHYSs9NBsyj8ohdgDheASm2Q8qZpu1ZnzdG4Ygh3bbygqFu6xbdIYkjocYqWdrgxY
KjyS/nOtQC+AAKEtiycrN6G0Db4qjD/bd0wDdHzkOHhuD+GsPJ+KZC9COgiQd+LEavaqV1BRj26y
Zqiwwrca0xZScr+5fYHlBND7uRbxtG7aVmHuWvIxItj27U5DGlv+DphBF2tj5rTTv0EcyNX5hXN1
1ystJNcUX5U8maQTYaqsLM96S2DaVKYQWW9Z8WhTEsBg2MTbm27dOBGF9NsQCqbx24YIRRUURqyE
SAgLCei803PKngvlnmX3UqQHLJ/i6cj1vq3sp2ANFeY1CCw4OlDFt8u5EgePBoHU/Yv1XYg4FCUP
jtGtYUzA4ev9+t6lv5CwymNRQwyTQNCjzjojZAKuD16KtbPpF9tSsCb6rpFbEkS3V0suGxPlzxFG
lS9xBym8YDoN05orsuOv9DJitST3qdRP5q/k05E4NfqONAXXskZhkiYeHED8O6uz6MJLQO1Ke6Ao
CR28eIftCdUgDz+/LtWxUI1zaSZh4T3MNnkYsnOJf8Tv1onOxzlIEVzFLdJrim9hUp5RBPOBRHDK
TclnIskdsmU0RmNBQXYWHnH2hhIgZHywo3Ci9rNJyy7IvTAAla+Mt/Q5/JJEAEnF3WjFgxKE2SOu
WWlDyMhcZkQ79GT2OvfxMx6oouWtrtY7h9fS5kEQVw3jlsw16aYEDm7NmhYUq+deN/EmMMdwDILq
es4xEgI22+oy7TEs4gb4iTOfntZG91zTPoe52eC/xWiO+PCSut1iLWP0jiJR5CC3A1GJUDd43vpe
ZgDBBuRB4OJDI3r3CaN+EQyWGk9hchHPqmX8st/jaWJwNwugkaEGPPNmGRPPHoN8/aqq8Ll6nVP0
GLuUN5SBvRae35oU+yTpu79AicF8K+qT0H/egH7BtbURRXge0+Pkk08UFrGNobxoHKPBqtSB2yj2
wKAY+Qc2FAEdblhrJjTHlljDvuKfFaq3Uwu/S0KLdRGYoGlfR2RHMWD7PxWGXhP3UkhXyhSVDkf0
yqU5CWgHqoOKWsaZ9h2nxpEDI9FUmt6LfY3RdwivZ49Aat4r4uyd4fjqjlzHHLbTZK6wUqjGDO6l
YdkE2B/EhbNatS5gXydoeTDqir0TG3flrbWivTJ+f80B1Pbgtj7vcbsSRcG/sAuopM4iSXg3alGY
heMCFpYH9+BjVvg2TI04zBM3NXbnf/G/ysmBOeuUIOpMqXnP42em/c8EczBtYUnb1hhU3OO/HGHA
QRpDMttcMlfVPOec4QYYlz8X6Bfu2gZy0FkRxEk3Kg7Sl4rwbYpsJxxNPeOATKtXJFVTxRuSZub4
HVuaa7afk6ZzHDQ6Md08TDa794meXbfrJtCiIQhZ6QViEcwAmDBAD9XErh2owzrbh7SrN0YmYBD1
SKMOx9YsrDjEs0L9q9Idczi9ry1cbMFv1JeFWwFS5BBcp/w1l1S4VEio1S6CsqmDdNqWTnnxC+7h
WZPMAvvu7Nwseg7H4CzwbHtAcoQQYU/0LKnXns2KaE8mZal54qVQDuQTVDZ5iV54SY+927lICeVm
iAmBHxne/Q5DBHpN0EKgT8T/RoygEUh2AIrecntV5G1NFXN8/EGCyYWILrLtjQLc0+zXycbbPVjE
8oI34QYqp5S6biJjSL+ny9kljMLXSUpLKdet3rEeezVQGQimJsgQWkdUrj8OWBRtTbJ6xTSgXlNR
yV4RVwktwfKlKhAf0dzTAG8QUirUjED87XoPyD23pv5TW34OnVvDDZM3DxaxWE3Z+ShUD1zwecbw
Mkv8WaURLYefpxvloAhO0DaHIxU1E9+rct9h763A1ElU44w7NMFfL16/2v7gMAEf0LDtAIhjO1QQ
cD+Du9N4/z2zJMjJQJYPgpdJY593q+/Q6jErxGWSf1IiMeb5Pldt1S+FHjvxAn8kivQZMvq4x1nW
0DQ0QsBLnU3g3b4FxEAwdMPsOWy7rDwSL6d+Yf+LLHA8dBHnqpNXAeSI0aQqd7Thi0nACra0Z0Km
AgN6IDaukfyxRIfFTS5AJg8CBAefPw4DbQZnA054Lv643nCepX/E/84ax2JzqY7YE9Y6mvH8eacg
Wm/IjwhAZbLNnjPOpvGDs4Uitk+b3tjFAZgPC4GOBYJI4LLuAL2jV4BTYRGylCJkrBUpEuLNaAg2
MtvFSsSSnMY+mlqKFHfaUl5AiinYhW1joGSNAKjY/4vNM7r/3i9Zu5zSK8ADzUph0MWNxalkdLmN
6yToTwp6T7B5Lwkx6RT5gqPpLedUPpgOJXcerBPeQ9TAN0JRu3+mnPxthqlaFg92rMwTvlCmtwhn
6jrz7jpUXNMp+RncCeKpBNYNyeDKZDqfypuzjgPv+NWBE77SDHW/IpX7/MofsU0YVwK5BUPJ068n
yn9ywBQxLiyK2bnnat03jiAvy69yXpWGo54pX4jrh5X5HxrxRVdIu+OJTD2p6l7YjT+3u3ZwhdpM
yodBBvE7qKaMpt3GESjkjvCKHi+7PHfvZhuQjv0G9jbbDAYS5zZ/aLSmqm4VkKrB/PNqZTbFFrIN
Ne85JM9NJlOK09MC9OJnSIy4IEL/Fj6N0bbSF5VfLPvijytPGoZCsdV5v0xOyAhB2fnPkqWpMz/9
vC5m/1dDngKEwpf+8Ew6XRcB7qS2Y3c3R7cKYg6LRA4IqBwPLgBD8lGfwQrrJI59shacQfX9jEgH
xBLDjISHq4Jc8LdObFcI5Q7OEQKGCT9pQfpgDUcDCAwAqz0SS2gNb2oYFsuTwDD4F0OY6RhFn1Gj
JrfoihGz6L8rOUFlrEVDzur3mqPWJ8dw14BN5mDCvxrb3Vi71OEdiOyX3k0ZBezhv4hE8AGGinDf
3M7BNHHkR15Bm6O+t0jElJ3vuhp43u4Gjl+q3xuRNur8GGNthXuNZshL+u3Lqtfs+d0YCXg7XvEr
Q36ipjFLxdKI8drnM0ceqCXnCG0PUv1X/Wq362qfxoKuhu07k6BwSojL9YhL5Oxk/q6h3aueo2kk
lLB9hK6ft+NADR4S7ZkcOHS4EGs2GdQ2h9yPNsi1F9VO+8m5/t3miwUj671q3mbGJ7KhzfKgqm9b
7x+TcVJocfDVWChoOTthedeBUXoOpBA8b42EFAQ4Y05BqMrNVRNFg27OxMwmhmqVF9jz0knqVGAO
ufLSUUyuLG6ee1jawGKwNVdsoXeO6H3wtgLnhSb1dKhzifgRfROn8KF4CGdF9rn7qGVonimf3JJc
rhwIleIL1VB62pJXQLuQWfol/msPrkMA0O6nRMrcmrmJgUbNmFtuAMYLAFDrHemrZqssOSQ2K1hV
xSyeqa5KIagyTMyBLM+iWek8MqAFANYITXM59q8CTVfJA3jB9NM2Moa56DdciGkIOuSSGn9gCIAG
sTFBtafCGk1PmP/S7DM08+9zfhdX3Inqg4WxaGoIZOfleMtTo1KhYcRE7EHqJBkIMMBww6CrcfTB
Y05sfm/YZbWntyGJp7OzztnCM/h4nVLsE2dpkZwfqv8ADIAV0DuuPL1XBV1mK7yR6IEaFBd7y5Bv
k9VVL9ez1nGl5GjrOY69/G49lU6HuZGvNGZDL7Gt7dS3vwOa0lD55ImZgWc+0HRcvJkSnqR/CwNA
1DsC8dcNGbaNCNgfe0mst1Y9QzSs5IdPqWbseudzd1co2vxkRxjy1LoWOez/7GussHy9EAfReoXt
KqsB89XBsa9zQ5vaXLkiWYDbkdWmuOcgxPNykwT+Q0CpHG56R9p3ccttFsNwQoRGFumAJRAMjBaQ
AOev5yFAeYI6/n5YaQl2kNED/3L6H+2NfJWrvBwHiN15TzLI1gpjG0PqO3wSmeleryHO5KfQUrfQ
PENjtfvO5nb6Hx3RWytHlwHumsGuhnbSLvVFiaZ5Fj7pfrL8HU8z3Gh/dYFSVP/LGmMeSVM1Amf0
JPeIUf6XS8ng3m0+YqUXPow4oYK+RvYWYqwk5AQNGJpj0BW/BjjEHcWrQtX0AibzNgwwRf5ZCC3S
lHHZcx1LOrX4anbWeFNVaxpLWi7/rOcHdMwj09QwBY0P3ljfbEPFpLvFvj+JDOFmk6MJ3LYTtvtn
p5xmE+T9vw18PeRk4m1vD5qOHUj7DEoj8a3Df277Al9JLOA8Zhl5zJoHVO1YzuD9DjTglo706dxz
PWbHoh3CJobzb+OhJCHhhCn/it1Y4DMW5XqinX+BJb0dmcRdzqDib8Saxn0LI6EnZsGd3Abivl+P
6cwOBMPwvsbJZ6UsFf0OLh1CuAEOsca3rYKqIlW4J7s8O/zFRBMI6Klkxkw+kBbKeEbCLdVcHeJd
nftJuByNl0aygzNVagQQ/O5ynIbhClkJGyNNQvuX1Ihz5gfszO64GzNPYYUI6UCzjQejLzOHzMUP
iTE603OGsR4iFBPOgOShhyCKjjSkHGXQhdcwCok8saTTmexdH84LkYUzj7vhnqiWVfE1LMjsxhh6
ua28LUs7p76QMEwZfzCH1FXV7GH367dGH/IvupyjLl07MU4t2HdgV1Q1BA+9aanQMoWUkSQiELTr
jqp3jk+eqs0B/hYDlhsehpsUHhGU7kVgqs7/+u6ou9GcED40g01ieVGotdxKPW8IURpsa8S+xY9V
fhLVHIyvH0DyUTLfP9vOElkobVeQZs+Y8aS5lfK6S3jRFOKDr/F0DOz6L2nfwDCDu8eQ3uBNGhae
/3rw+Yue7ocQ5aUxHnhqBZHPQgc4votBHSugF5der5ezZgHTpSR1mLKfA+4eyMOOnHfsLDvd/XKQ
KL4pfaa4jh/LFNtm0JYhZIgYh0e5S/Jcos1m5b+fxp62CMcf+wbnDlNzhEB0+8t6PxIZuJIoW0xc
zQaCCSn3T29UfItHd/GyGsEFBfm0z+4gAe0XX6BNl0bC291+YYFx1eHkFOhu7vy80F+YFPofbnWw
HVpkXtMVfoOXAbnNdAb3K8LmhC9mR93ZWOJhnKVPrqRLtlM+fQ3v0aswjcsG9bdh/ZEiQ7zscSvm
PsyNC9DFCWE1j5H2Q/dvd8Yjg+RLa6JnENnoMMDkIu+3TyLAZTgKTDIM1mUqeOFi32g0XrU/rzA0
GAbTut1Su9GKMEZzn/xCsJ1aewO22yRGtBnPSSjW3Tze7bYga4Ubt+6SXsVEJzSKdPlJktZjrtx8
tZxhIpy6qfg1a3/sVxDEo56cWqSKwaSf9Q//CldQNPBkxYfjpNrnOgzsX4LywGy7eraxYTGBmgXT
9q927Ei9QxdiuJ5UB9g52SS8MdUwkDFUzwJhSCHLhlGRWoPTwIjWc/RwJvQaF6QJONMy4OyXAcyN
cUIHoO8lxi6oe21+EQm/YcqVai6aRsa1z3S+x4gDL+CjoPNCLGBd29IE1FMb7RQ6LnhTJNQeHKgK
dJobaYWIsca81pBBwmA2sUk1lasy9HOyWuIi6UwQhJA+/nT5jKBDqPL5XKwHcno1woQNwyYzdgMA
eIRWE1jDEh6bRzpkCllteWiJTyy9X3SCk9FwJNSZbiBsoI4PcRtiG75MzYF7Jg25fUXVs+nrYCRG
nqlJtL7MjqFqBW8rWiwCtLPMJGn4bqaYeKbQ5BgRQFGwWc8rH4al8RpHAk+rj6vynEkJ1yvGQp0P
j1fIKjY5hWpHmR4554VohANipblGUnRRvoPGxdDkhvuLBbHr7fQtib0evX4nVbbCAbUoZnond+6Z
tyxzR8VSakLRiKExIeCjgeBhaY+RLmGdY5oKeETrJZr3temh803WXIHLRQIMDdbIn7e2SST5/CTW
XE/J8MYG/qsQPm94ZKGjwQdGqcxSPh/IkDtXcz9TAkCmo23BIG/msmJjRfeY+4fFCvUFRUL/HPWL
X6rnfKU+ePb/KiL3vqH3wikzOq8mz61kbCFKXSxr3Il7i/M+JHIRQO4p9ldv5z8q0DbdJitHssj8
Z4fme75B/lTRXC+VNjmKbrQt5qvuRKWNRs5gislZRuqBEJn3Y44AnVJTdpMAX2eEHfIRvLwwUUAI
ijGyvjEtYgJtoFzhyC+taYMF0csLLcFR7nHj+JZXmCF2J3/RCc2AUoT1hlQ6ZUDfV6wtQ6Apw3vY
+53/fjS6GqzWRtw83JPcMyvvdb57Sv++7d2wAI2zQuBBAwX1Kft3Ok0ToNh8VshHv/B3fBrSH6AP
xTvROjc2gwAlGomZKpAh49ME+kHdNAlN6bpz7rONJeBHQOOlmar0HGglEX2U4w40irOxIqcRKn5C
rq6tOF1UgovKOSYLp2yx/OXvyfmTF2hsw/FPZPSO/eL08qNSwXA92+qqizGQmJoWasuJ43kw+q9B
65//4xbaOwEq0VSqTgsXcY03Wo34nY9W+dF7Y7/C/4BhXFooFpRSYs5cSmV0NlZRRZRsF/0+NzXZ
RL1wWYY+0HLr64IGxmxMtIQdCy9kPLSj9NZzX8sIe0/jY31MWSNgcR4MLmlxavz6pY66Dr2sqLCX
Sgc/OwhfPktBoJmcxRYvcbNBiPaEMmAGnJXpJEy0InORtD+PW7SPVFyMcFNJlxxMZpKsBOXPuK1d
kdoAkIODivx+wCpS23F2XORtZW79da5Y6eT47eQ4tXh15vAVPWWUcan56ZvYuOJGmWcdnWYEbbH1
w2sBi87JydcalSFeyx3APPArpITRECeq5/NaSIMWsBb4KakSiJHjJRlur30mqb9gK3ArH04qPO9S
S8HUQUHMc25jPSMGkfUJEL1bEi9LxvAq4KonWXFDPt8tpik1EQICmm7uShImxOi/ZmAACzbucZ1X
uH9cL6e1UtF7XCUOMVMWv0llGUkqWaRoR+eU1MIqKqEPP+PZhqSlGe2wucy20NXuQoD8B01JDanL
HMAsBHZ1oBRhzlZQI5amVqQ+jB0xOlddDwS87AyReG+m150a024CfJEW90GHYWrrHIDaV171XzQS
Lk49PAxXKw53lj99XwMgeKaMF8uAiregJTFDZjx67cJHeStjKa0OSBw8bxUcac31LTXTNZ3JLjvE
Hv9VOc/UtTcALVVr46W21PaepXoQvNqKrlZBmW8EYsigGAAOKkpy5rcMN7t98mLIgnVLAJkc4W0D
wg5WWVIzgvlqojTo484BoZNNzlNCljVU4EPQHMdy99X49et6iXHi/Ql70wTscj/hNgZRFda8y+NU
oFbh7PjyOHMzTuhn+rtQI+VpPSubt6MbdE7Er9pwcx/VGeXXqtNW1Chc+j7YahUTVmGOz7bIp4Ns
AdgcM/uns+1WCnSyv2FRByxNjEX11JT7sLu8qNDuePVBG7F1j+xdrUYE9W85WqLBFsVs3hoP5cZG
yevHbSPcyVy0WFVrrzKRduJywr21Mk//FYV1XTAJ0FocuE7FtdxG1ed+fa3FmCZDG8W5y7rez4MM
bvR1UonBRjFpxXsnIykqkWNqqgVnvLF1pG4j7y3tHvIyqmu8X13GiKOmCkeXFiSacrr9k7ZV49yS
leEDVzhsqFrmL6RZBACQExufHXlA9/Pt2IVi/mr8h4/G78lOXViubc2DYqPiHD/nCOAPRf0cxltE
p26SOnM+jXhE87/qSv2uAECku4IO328DPwUCZtVj5GKHWE/QwUgUR+b2npSb/CY3Q74V8afwTqVv
OA3HHE6PExFSntr1Q71DPIhfnXj93luAyPiNFWWlZhbvnepsh+HQXf91ZHcfU6zSOYQS9X7FiAss
+H99L7KXheeuxRIQaoooumQtERelHKd1tPwMgaCSGJEtvsS7VgEmTzaTeyXZdEHEhgLIngBmLHXQ
BaHkiTKV3d2MiOIGXrygy8WDtr1kOuMUgjp8C6c1Dc2rcXw/8Yjz9MWbDqoJQR28FX4qXKgJVEB8
7PovktInPr6iE8gVC79tmExwuHVtPXuSGRCYEl1nMnD9gjxnM62DQjkKxXXWW1c5F4O2KrmtKjqt
k6TuMYLLenm8TyQNzIYaXxvIwSQHlIEYevVvaDGVoc+ciEXlpzRZe7cv5xDXShnqGUF//hVOyExI
dber3iRDKsWFxD8y7O1gJIkvjQwcN2IXo0JB4ahLtY0o7Z7xeKnae5q3G6xBjBeP2UavJ1XVp0Lo
gntj9RzdPAwx0Xq0s/X0xaiNbnysHaIpa9GuMwL/Nf0qH6qKjDttKoQoIsG+qPcn0t+oYmJImXZp
E/IkaeOmtRlPWIX6Uu4WygLax/+NmleboPC6JFgGWET3JtjutSlXQtyEDkbTfgNdIZrrz3X/Jnfh
plc92FPukefzvhS7ieMFMWUE1fFr3bb3Svb7Xtxy0ttnC1pEA2BlrOWIct5VakF1gqe9YSeZIpBz
bKqZX3Ssde7Sz/zYUzG6ZRLTRe4/8pgpzfL2wTWTzdQAcpV4gXjmKkbmWafVOH7njPk0ImTVx/Yt
JQK3RJDNM4JFK4EpfzoTtPJiipTMYe2PWsVSXfzIk6y5vYnxwCDWkYW24n5gAq3Erm8MP8FCXdZy
c+F6oxPtES+4FnVS+l7+3IWks8ychyjDl7CNb8yWf3GYPNrzZDIq3xHqdOpJX4vQgQR0CUYUfME8
C2itNilVQVLopmRJ/alXPq3/3hAo0+l7nENwkp5p3VViMds/dBlak5tdYy1Gd//tz5/cC++qj9zb
xlHNwnCsdlNUwoJCinEcxpuowVzHDl87RmvAAS8FyPGFrwKlPjnhLMKm2LI7bOFpMBgZjAgXafmN
VgPX8fFlc/szVcMdymfOhYXYtUasMR8QrHGjdhJYTHB/kX81EGBbcrnBY7Q1oAAEerpjAjL7QA2V
xKZN9btn53uvlRrpRPZRo4X5PRXrWTKwvLqS5RGDa1VfF2Un7jX1mJudcYa+6NPyPzugqkJDYJ0M
kAULNEKtwZ39rruEvai6UHEqqbwvoN3OXgIoGYNHUhLfcDjET0qW6SF5bgWGB4JI3jvY5uMWPNh0
BHzZEbfPm10pKRThg3ykgng+Px7rZUMdmU4DudS1INdgMqHh3wKb7z1aPvJeNYgyuI+C0vJ07L71
UZebF5k5jCDWmHkveyyS0GMqL8sjwCMhw/VSvzCnBnHvJUsADCZwX+u5ZjzKofnWSlw1izgdxPn/
D3FKvmSNGiFdfyCdr6O9X2q7OU7XyDJuqSJtsVrl5iaTaVnchOhmn1+0799gHbTCp9ry5fflDWfs
b89Y2fxhZyoVG0nJcomj8ynAUdTZihKPyiIoACie/HNvg0jiWjU88E806r2anbooV8Dn9QtUMT7y
BVYbB9ebmFZj5zDJ+7CUXJQS8eXXpFXK1FY8gZrZubyXl+gNauk/iA/Dgz0KzzFUBF5iwoYVFBZv
BD1hmXVTeV6iXnmodJSEzHKtqdA7r0MetDHcMT/Mlg+mhXazXFyCAfhbYmINx63dHRkF/p65Gb01
vKGOrC/8/UMsV+yU59g9ejVDP5pH6iqHalDpA+FcN2pw3QmUZBhQncFRFQaxL8R0I8QCxrkO2bNx
qMoVz+/d4ZtLbGvXf8EPRCo+llAxlcuBmYAxx2KoR1ljzF7S6WVxvU236JeioZjfc/HuWPEny78b
SGoYGxCaw/UW9jfhBPkePOl1sUrvk3T6clXdzGFN83n9lLiH1ki6EUOQ2Mpga3yZk2kIa5CUuNKB
SxRudj5Gr/ggL+nz3i3ctFMLWw3RGpnk/Vb9M/6O9aHO67Y+gvDjQj3+Ig+awCg9Mck3G14kgyCK
kyVowQTYmQqci9V119XvjAyjOknug6x0qZYQlJpDIrScb5uThc2NVLEmBAPXKnEh9Sy13Wkdpc/Z
Eae5t41wybWRrCURqx87avCUBa9HKUKOBB/mzoyW/2NAuArInJDXV6TDQ8sSIlif8QnWaZPmlOB2
cvz8e4wThIyFBytuo7WSXrAsKlvDXh+RbBbUQG4Kx7M+m3Vtg2FhQR4TFwmBVnN3jFTJc4D00rKW
q8u1Pp2c17slp8PRWd+E/6KYak6fjC/v7/wp0rv2tF77OhwmWFCp5fWdTkknTIAb4MxOdABqT1QV
5bIXHVGn7vzU7mleQMDd6BaCGkBPgmW2YMJ4nGWTiXhwiR8sGyck9t2AfkVLWGxwTA9dY6wiT3qi
iaLtiP2oOx91WoXi7jbN95qiGeDKL0oFe/297G73R1DZGNV+CbU7YnO9pgNw82A/n+KpFGo+R0dK
AhEbrLmbeAArP2J/1PWayBXiQPSQCEpYMpboVc3oBuWYRbMAvA9plFM9JT/zYTPln7S5HSFI5tY8
sMTM6bXG6HqKXwP3ACCq2TZUX66UXNMgY72l7F41tcBASDOI/CHQ7SbPG5pXRdqh7iIljxD3Pf+4
TxCRG8BTBB7xRDy+TVuhosL+AgYIP3Zmd8FgRZhcyeiZzoRSFIqNNkS3FjSv1TKl7exIbVmdAT+h
RH/XK4+kPuja9BTy24qj/GMdf42lh9PgQIpUjv/84ME7gfox6435217ISC37aJVM5cpRUJj7OscG
W2qEcxzgLZDwtCWnilS8ewj4shP1nSxQ01G0oaWaKbnplqcGNqqHXgBxMFMZEH6G1eUp8XipVh8B
CF0+KNrV1zclOHuELbVTQiFjkHJJTiKqLIkN6TgDV+Bp5fZhdLkrax0r3VP0M5njuP9Vw5ICOSrk
igQpR8lPmMbNcjiD6DiefwJQHHP2Rzwc7DSW1T9+lWdTjx1r1VclwgcQiPD7nDIzoWxlxsgCeuLH
opTIMtPl3aaOAtTIiwYwDyX7Khxwtp2qvttO5mnDEbIrEtFaTppIGmfQ2pURVozsqk7SDYedA86M
ESMQXyczu6w9e+OSJZ7F4uAm/Z2n80pMZHQJQvctfB3nBfXYBO1MLHEIYvmxJPjfjLPnQogKRyrz
S7wLWPAaQhvVtNuuxIuDteRH8gEl270FolzAx3eTLPdxzCq2hk8rYS0CH5/ZxdIpgYIyZVfxC3pR
d6QnPi3NPq9E86gwc3IEtjExVg/HXZWYNn+sPGUOmvJTpopV8gHNTiruOzFBTJwPqfQdFSfKEnpB
rJs6k0q9YB1T1D8xzfYlt0qjURp+vyOZUQ9SvE3Ov4wj1rfRdynIn3+pOyub3Ojd+kksLWIxslTH
n3vfT/KMslejaM8z14Q5lqhnn5/sWQfP6a8NPoxSyU+oI9/nfMckxpu+ziZmU3xX9HsBIznEMeJc
8rRxEn/rQ1qNfcPpPn1LL5LesUW/wWB0idiKzr2xeCWwoAELEhLf8LDXC1MKNdxUqe1ALZT9G7nR
zu1loygILIkJbs/J/2tc2Shd+kM3jMjR21b+Q0HtzD6PPanvWkAmVQQxSm4xM4Cawfb610234oee
bST1tnbDNi31eZzsEs9q0fBh2fAZ5EQu3jAepu8y4mFlXK9sUZlTl1plpcyBWEgZm/xT+5DONkws
QZNPc6pClXLKx55oc8gYTXppHZPz2A7/F9NIWgQAUBV/bC98rvGoFoyQeJjJoUz+L21jP6weN30C
Ic6w0Gsh7TaZi3+art/QgpXnScak+dQL4ZV82QE+ififwd7PnyYMgNO62I/GaWnbMGB82pV/B3hL
LZe9lyQ6HEMrYpV/63w434EMg4lICjfC/Sahp6LcLjYWp1JByzRCLorsJTNCn2A1CE51BDjdBVhL
hIU9n7hAQiXVb9dVkACxb3h83cwBQYiYAgMeTESQw+yJOlLvbr0mCkl88qGMuqcOaIKzPqkCTfkk
3edoVanir4hFV5M/XkskFrYaRr3RaqitwfYJksgFGxL0UfJkD9r6EoAZPm4UdyEq7se/MdMmpn6W
etu4UK3OQUMtxo3hyASGy8wwNcz08Yu7QGZPSbX7bwTDLj/ggkkhBTZGZUTbhjwdeMWLFc5vIYMB
uJBJMPWl9LNYX/iXQJDApOMRqgbjhv0rv2XhOTH/0qloI77qinuyqXqrivVItJM5EHDiiXwrIVlE
iEdBqxSnkSGUVo165G7PHaMln1PiGcru9tN+g29pIR6MMY8BX4JqW0Itdui/FpYd/SD1MR6YlkBJ
paYI8XMeOVOMOerGgrH4EuwXoWPnBwJcXwj0oZp7UJ4dd8GhS/aagZ03h87foKD8dlBNdSJkFujO
qePOdkkkvj6hQr6+oYcoDwFKlxaRsdcuk5mc2j+Y76W5NogC2Xl5n+voskOVWyuHJ8WC8qkFIAlw
G88yRCaMEDXzv9s5faGVQUDrEd62KKBshPPikcmrCmUUw5cY7rrIgDocWdyMIfVOkFMEPd5lct7B
lTIZ4kK3z9fzfQCcHUvmEq8tm9wJyLo59rsvNVq5yS52TxwllcO8KVEKB/2PBIusNUt5m6ipA9kD
/Z4CGs+Sm6HbrDZVPqMJ8UvPJZIcJl+HBnI7Cu/8t/QLHPiOwgtidL115/viyUoaye/ACZznuFd3
SZJECjr77xMuCJN/NnroNNd3hHkySiwR72zvY74pwc3nqbsz6Eny7p1s2b4a99H2mhoSROp+ck0j
HmNj9wz0f0Xau02G9pdy8lyvErVnwqZu3udjHJSXMBUW+BhGzwsrYPtJ3BmEWuOYAt3vAgKZlQal
+0u+t9T4o8Lo4RAmW7TGhF+a+4IGRYPhXpZkXyG3VVwC5BmBtOgDxuwRoz6iRszceRIKTMKzIfZ9
woCGTmNsALvzIl6ewpoZDl3hDmBfMgpegutQL0TW9W+odWBWVOmqsQUx/0DXzrJMzTdaULCbJM1V
LZPQY8HOQ7dKOywXQGzFEOKtz33uH6W+7fhJno+grNTi2bupQ+3tG9LFlERVOKs9Rr9kYRUstbgk
fHpfkizGirg4sdun1C8mMHpo/LlsPcYJyKPiZZcAs69FOJ3FR95VPN3td8UtK9UDv85JlMoqswMx
Tw8t6hz57pYET8MIEoXjMmCUw4jXwL1mLSz9PJOiKvH1cDHcdwrsA0evaMfuzFJHUBjixtNc3v6O
sm0LFJpt9XEtIRqC6sU9cchBfX1Ph7dzXsadyTB5UOF4hWZKxZWnH76QeJwKILs4KHX3i4HT2MEI
p+7z0+ZpR6mkKP2zANiC8+ik/yHbMn31aXIRcczrzvpwkTXlvHp9krxI/+17eN0F05ZQM8PYT1qD
6I/i9fP8nciLhv/qToulUjwQHWEFqlUrX4H7aex6054+y18ET0WMFCM2fGAHIdKDbpyXryIpi6PF
BnI4l6/pLLyumrQXBIv/WW0j4KQiDE82vCzBj44vpuRcZdxyz9npje+ZCdfdR0DuegxAsgl0zJ7S
Y6SvtPDH4blIYT2xOGfG6FhQEXZcqZBDana9BZ29CGblFOjqxn9uaUJBIa4lpT0uEd4Qg1Z7V9z4
j6+gWHMnRyBGD5+f0MCmo0RA30LgpXR6sebC0/ZhvBOuakbC3moY5ojUxMouRzfY7LQDKODtEjWj
7Bpr3aRv1zVFdseeNJVJxnWxUtlUB+efKKWfooC3q6TYh+GBCy9dTp7e3bIPhUvLk3a1J8dTaEWv
TYVr0Iih1fJD1VnayKcBesPRPFeU3AjwkO2U8ckhnLlZ8HiuDVw5dTY9lVsrl+8asYPdbaInSqNr
hnh1dPHY2/TH7bU3UKP4YAFYyXzXJlSOy9R5zH6e1/M2j8OCmqkIXpzqx/XxcO6rHoibSnG26XEM
EzL665P50vrqake7QnCGQVND8XOQ0c+94Vn1B7xnKpNI4boy0qu6K83IrOdcSmJQDD4yVVLq5A+j
yjL9RerXTwS6ghrA9PdZT9Pv3GITlQULG8lvVFWHmoDXdzOhxbczuwGCJFlQWz2VYXj1MAS/GCUh
0Ruw3wCKLn9zqGnD2nuSjYK1vLytLaH/VhzvivROTxuJzs9ay55+OwKUpXD9t7qDxxpoJIJyIWT/
Hze1BAxrJLBaKUtqaDos7tddqPxuY79k48p9C0yNnhjmNQdcLk9A57HQJQ/GYN0n81Ah4GJ4+8zl
LefPIzXQjad3rvAcablzizBfPMcHA7q+QjZCk+b5uPtSOJXArnRbfPO70Yi87XnqMhfM+wUYHbxk
Nxhj5ph6RfQ5YfViKJSAoqjkNAiO2sflHaWCML6ryCdjR6doE3TZwCkJriCoSmxvk1B6BLqJ3may
4wess57lse8NQJQKS1cNGYUCw9IoWOdyoWnkXRIKboihWHgMPkxQoIsIsdU1gQfzzsr1tio03s7T
PnmtZIDNdU/ZIONzmBE28R4Om3b8r620Q/87j+oE4cYVHHMBRZoclNtvXRb+5wKpAP8WukxrxVEV
b5GAO9Tnbn+PaAYIsReZFZ8fJ/5hcoh5nnGVwl4dtznE8ura8W6r/JUwOj10HfxKMZVVekuAWE1s
a/b5ipH8mkTR2/AZ05a6EcKIw9mbG+UR/BKOcdUyVCbwI90mOVwBHtFvOWS6ju/0mNHH5irSRzKz
ak1/HuEEZ9iIdiCyJoNhkWCAtWBj1nviaT/+1dn6TPAwV+UelZimopW7SlNZd+dldKdkydT/wsGe
pPUs1v9hjnj0E3RoY1ir5GeYMkGU9Fk/o2DmIS/Smrpb2Yggsj1TNnd3rh/Ke88GrgMj21COG26G
h7HGU/DhvDWcT+5DvQyVjgmDtymTrNyABKisuKD6+hmoJ9JBCvmryDvn5sr9Ll30YLuGBq3T8g2n
+4VOE4WlvQCjWYoD0eHezh1/WAvFO7JNukRhaxd70sn2xRZYcznLLw8VLzksSENtoDL076yhZ/jm
bwRqvFYy/XbN+CKmmKtCQHVG3y9Qj+FtNo50CrXtEEIRPl77w4I6hEr4Qd5oiNR67I7GyNYLASS7
NFjyIrUsXi6XEUAVGtZK6b5EH7rVHvzQOqFyM7KV/UbKhi4lHP/q0/hN8tqA3Uj7YtNFHo7/wHvd
Q7RSNdZAN2i+UBlWeTdJGKHrFRwkg1eoS6mFf/z1+8kKBEGX7vY0cjZ2+joa4r8B1ArO+eOyslew
XXP58eABDVf1KSURMn0YD7gDEcTLIOcl1ylvRyG4Oqj1+D9ibGx82t+cYKeMRNP4g+fznPbHgVAf
N1a5lGNvFPfRj7ABqXR+UQWoLflZu674HoXXpBymdkCp0dwy6153CNkffnsgbpjfC6N+BrKIQW6j
2V569JVUZ/owZxvEOwz+j7LOcz+l4mhMexOigoUZSxGHrKd/e1uQLxZNajGAkca9y4k2SBs2pbb0
4hTdaJiBDGQAOPJayL7e0thdmpikLTDa+b0son26nvR/rNEVyzHr4Ba/OUhj5RFuc0ATiKr6KBhk
eLCrjoF7VARo2HZcKJRS3xJJhhTu08lajflP9VZJ9Clz/kfvk/hoDHzBdAyiUI1fYn0Ai80aL+PX
3UrNdUEjqXxAvdvBezbhxZnQWx0R/SXF8ZRyx4Z23gJ3IHLrJ9HRmE3+3c1hVVY1B1rSOo9Vm/IP
J3ghRcIKRyLpHF/RZzO8SEnYf2f5BinaNAoOuo8mZN/Zz5ijq2UQCk0+1Vu7pzeOQCBuljWSQHCf
1kzwSfPJLp/IA0BhzoEq17C7ZONGhy19GNESfS9C9nSeyiD6j2cMe5XzQYk3i6e0RFGFWCTVYagK
N+9fidAmIyC3skYEg5wA8OUVZS9ZrxlJ5jzuqGRn6nTGCDxXThvOKdOFPdMX4BVqaneUqmjppQRC
EDoW3ABou4R+8G2agY8q3oDogakitCyCn2JI6SxQOLkaddFBW2nkgCtjdzk/w7A1iIb3JsrrKe/y
k6WGD56rd9mYwnmZV+7Dm85YO0A0ObEthDNEove7h++XRvSkL2mtZ7t5PcpJbu0FxUzq09nZgHHJ
EUeU1OQ8UZdP5aarsM4s0MQdev2n73nmIb0l9aJJyO/HQylBFHPeOi73B8RaL6UDVKi10S2hsTWE
ctZm8EzjPgn3GOcp+RVqdzrBqJZOdBSKqd1D2Dj6neqdO3rmHTvMMJWbZQng4imrCtvCXLoXvxU0
UWqxzlLMzLuB/eoPgM42zWyVWnXGEhkN7SV/9/NcMoD4LZL1p4oLHgDjd31Rr0BU2RlF2W0hpeYC
elYo4XdbZDsxHSkL8tFIUOaJgn3gSz0VzFzdoEBrGwPXdIHAk0/TN3gmqOPDeNl9L9uPPpfHS9Tg
wuXjRZGB/EJrYT9kflxm88+GMlWpSHBdh6zpFQ8Lb8bfkOOHJGvPxhRoYlSCajJERKDbO/T3IiPy
ngB9xv7RftmkletzajrfS3/dRCQVMNbS0/Dw+Z8pZ6sGphaMTfodCtPpkxN6+b0xO2/w4NCPYgdb
bGyKW8/73Fl87HzwHCjdMXAcGzi1rDdZKEOwdD3VQDSnpB7XSVFJ8ocaWkZyFxoKiHZey84OfeMr
rHoVFRmT/14OSQouYJpKC+1brPxnXXGy/BGZTlfcY/ycoUH9FRRpdQJrsCeI9gqzUwzV9UMftzF8
rSNn/nkwsuUb2v4DP+tQocJOyl+qmfzl9AX+VCaM7r+dS21bF85yTryY1PT+ThDcy3zwsIQbJgbO
VbBmDI0q3Hll0bOTsN6ecfhI/LBq2HO/vFfgB9xfuUOtUVVb9rntmEqHqAM1U6COuk31YfPdc4Uv
oVrKBL6EAoFqcwbGMeqikbQt60ybT3W2AU+tyN1r5UUXUiM7Y240LsAjK48juoD9a3Dq530+YgTk
PW2MhQxWRqNyESZdLGZfjw6qX1UtBw5ocIVtKnk3uc0l9+BCWqsurF190Zh08fAT9DwarO1nSfEm
psiY9/VosoJRehHpFE79wzbUV53yW5aVKbYBCrCq42Rc+m071Ws7P80qP3Abdz5NnOTq0R6GQj5Z
idKUtLiGu8w/9yld22kYqVXPp1roLtp4OZFOggwahWSbuKDhAzrqZ3QB0rQId0yiWbi9ecRE2/sZ
iEw+0Gt6jsIqLil3g0vbEnOlbZQHV8osnrhwGbj9vf3lmuOZkk12jBr3NPLeGcbpkLP3Gt4NgFQ/
rilxvYNM6CWJmvXHYeoppkY2EvKaQ7Ckkbpxa67jNXRBvXA6pxXsML07BmR8qEKfZl9WCic0INrN
5fnwKgAyAS7gEX2uCk0dogl45519NO8FLC3dXua7N6lVa7HD8Su3zULkWTOgFmBegCr+IKFOuW2A
bwFDlz+0/NU4JvjRv3SYZ5sD5+1F0SfgvezizsbLcSbYeWOnCl4laJyJ3dWPc/wIMu9XfrZ1HVoK
pFY8Kmb7D1E+Pn5UmT67mhi9xwzEfsG8uI5W4O7aYgoV8ddil3VXKEPHLmA7pLiIdo2YhIAiSGDI
Dk1w0S2vY6IDJz2WaJ1jQB9nAXQc1+6c3C8/BdEDwZI3WNr0mGmPupvfCriHwMtF7l1ySdf+6Mvj
zJ2qojSetDi7Fdh5UXJavtQhM+6yFZWYB1SeCe/ajEZzpWbuQQ1wRgrwFz3H4Fn5ugmAWQ+PiAry
0zSQj3nC5Cv5hDUL1OmI2X6LLeBqv0JrvNKIdQ1ln3MF+10E9BCcOAtF3Rr4RV11XeXx4KwAOCbz
gzN4fetdoCERZvdpm+NofQFtYadq+779Wufb/JN+AHVAfmUB6flUVSqdwDWFtXJJb679mW9J5n6r
6lY+RcLnNtNjIMS/PdGoyKRtFuZ1HUxkwn7WlWLebNMR+R46S97lhDMvwcSdLkyo41uMq3XSyP0S
xjME4PK5a2laVU/vMk+tEBCr+6dlwaZEArxXKb92jdBpCz013r2R5088mzN0NYzvbTwoaNhWH2GI
gF4Wbao1AAsP2ra4luARXWQf3YfhahlmZ21zhEfFQ84+lxdRl2Ij87WqjvmZE6L/AHFfpMI6Lgg8
GMu8PY1zqT6VjOqJgKTwk+u+9W5acDQXJnjDIvzG5UgIKlKlLA1dneDGUJlWAFLftdqfMJsu+RD9
b/Kx9B5a9gxmd0RgEq0irA9bKPVmm2TVEJnS/4KEUxV1EiokN4bsRXClidEBP1XP81IAke/wrsAO
x4+dV8+4B3/QYffGha1HLL+E/TrDJ3TS3sbSdghz+jxpsEIU+837j+lmhd3sZhdxeiwFXfYFlNyW
ez4wKNdnFPCz21unBEDNu4f16oQHQoTC9VHjlZmTvBf4/9vQSIUm9kWnAZx2kZd3NtfaDjZ+qi7d
c9iZ91WwNoJ4x66XGfYGwgSGtAYglDqnYaqJxE2+3Ca0EwPElgQvkA2t537f3Swg+dGKKOplo3b8
oF4JXQRNiE41Y6gLoGKYu61JSR3btU6OS0icFm5tcSPdINndWMnCezJzs61KNMydWr42BNz+JuRv
duhTmVhrP53V115T6/rBcEdaUKtYGjb98K9N3TEOt4N84Pm+lWq6wBl++T9+119mgXVPinEPzWYb
WO8FqgMJK9ENBTOHMtBNrqASVAJ+2RXJq93gGfzahDPhnb3zH67xk5r/IG7OOLukRLch/VTxsOJv
sPJToVhaSq8QDFzmXVd5/9zTNif69zYtoxEWBZodccfAs1Iiki9wkjky7NHxP+jPsCsGiM4TOEJ/
xdEOeJRf4XE7v++zvOVxHEIdmjNAqx6bVymwgcDs9giIZmuk1P7fWUHu//eUnxmx4pWlixQFoaTM
rdOaWkGiOQ0VDtPGGDNVr2YUtu6Vmv1eT0JPOtsqaoxcy1zpr8ExbvjgHauR/Qwsrx2+fFPZtxYI
PbAsFdx/EvlnAgIC7zzWuAtGyqghy8ZNdp++f34nWmGspCFa2P8F1Vk9vo3hhzb4YH+T5lSgz0C0
UQXkAsnre9Ak8VrrqXyWYAiaEY85CTYfN1nqnaS5ByXytTGAwhAkYKKpl495p5nT6ikXE0TwZSrD
qFxh3hYBirolzyegF8WqaB+PuSI9x4jF8/MKpKk9JpoorBK/pYBa+tMqA3jThxLgLeMrG1G67VEk
vd8XdZ3PSl/L6tZTbujxSQiwHY5uJD2z4TEVuoL3Q7pS8ispdGiYQMQ9QJ9vKa+tnqLNTQLw6VtT
zrqS3rbpKWOR3MvmcVz4vnioeshHOeW0YjLcRHqbu7a32UcNa6Cgxp8cY/w64M2zNNnus9L5t1z8
OkyFmH/BLvXMbnFrdmmIpsXEbrgwrN20SNBDZjzaMhTBKn7xxxih6VXWgARZAJBDIk4rQOOCxNqP
KqgF2z1/YwEMpH+aNjSzWOdOFwU/C0lqW69fysP8u4DIDH7DaG5pmFQ+zJgnY9Iz108e12iAW/o/
Kgz8oSN1cI+qtc68k89UlMo1SQmqYxx78zfWmOyf8cUHfmQaqr67P1eHJmkALF3Ij0wv4E5YPC9Q
uVTGmR0TCWiT7CVwrsQNz/S93rkXvBj8SxHc4WfKxKqBk1y0w0T016msaUPXkFGhqGQK97kkBjan
4+pcJ9SRFYMSoxbprj1raoS/8GCoxEAr0uB31uQ6G8tQsWCWsskb+soxZMDXiaIlk7p+NHJq/C6C
gunePH3EmIGcIz8xXK11KoG2eMHlT3q5g3bFCZJTe965vRYCwRXXbyQn9rLE4i9JyDHd2nwC8RYx
NLzg2z6y8zf5J28R5/YzghFNADQRrnRmEAAxGpqIoVfm3LebJ6Gw5Sy/I0n4PTICPwFTXisiEtkD
INIdt9he4nj6T96cr+ZaYnresviERDaPEbuw0YwTC/+MHbGdCRltcNKO06rg/WjyvR2RcK+iH/OY
ByQKUH/8oLsjF7657SghMnh4RIdzdKBl93OywI4uoTJVQ8cC4xGBHy4kI8scaCp2kt2bDgxuFzpt
A/pbYPoSrY41RRo5cTaQ1w7g8NIWCmhc94gn628YV8njZ3OQGkSoyAoqW+lxAc7KpxqROP1Ulpli
cYCMgSDWSDrqtG4/z+zMod6BopRfsnKpE4Ty2IimRptZ4mqy1CMG3K0rgrOS/WKR0vSLmL/hgB9m
bhjVHALL5jBHLYWaoxucHTC+a9yOw5VZ6cGdCMVdGT5330Hq+1LBb6P2wlNB2x9vyCDVMFTgZnCp
rVCtMHJWHIAdcqaR3wYJaMlZP7NRTElEKgOcaNVg+ISJjvj/SadZ3HUqYC8Zah04zQ+rIWGwzrMs
/yLqdpPqABrPv4uC0WTbMHUkPAQC4z3kS4Ku7K9qKI8MjhOOR+JH7CiLg2pe97OWJdKI4sqygDaH
JfwYLcT7f/oDQeJ4eaMuWHWh6RhplESNTwS2NvKTnKyYZFNUtXRYHe4UsOSTuBzEelkYdZX6YMiP
VLhFfYjSnMPFRSjxWGfz097zlT99Cd7XyyDW7JAX+CADniqs6Ltg1nHQIre5jzG2xaPahuTb3bO1
G0XeuohC0DT4FypjiynuKpkszS/UqI2aMgodJmNOHDjrKP1sO0OU6je+UDqZpXpC44JBmHP7Ufy9
s+Fk1dgtyXtwggEqQT8RxYJr/FHBlv3RgRCTJ8thWkzmiqk9i6t5p86TAW5QzZNbrfFhNifxAgQ7
HR9A6CFuXGBFdX+2jCCG6QJTGR5edRA4g5HmJ+6XdMzurMUkO8jQkbELd9dF91mF5IeHYJ+tYLjC
61XBmYnMQxEV8M5Ju3/0YOI8k1uNJhQIIFo2rsL+KZhce/5KslcTF3AtfhKh9PsSC+jmgX7lN4Yv
hzDmNTE63qI4c9lWcs1hL0uHYLp/zDVZDgKgz31inwwyqFndY8hlWTT9XSmufPP2qvwvXcWIKe5H
HH6VGuX1lR3+WoqaPg95PEf0xZH4bHuqWu2SLJNvPaSHORiB+2P1CPHUyx65PXY1jUrac6jfJFhr
TNBuAD/0ViRvUhTYWoiLtXJvrLTO0Ja28ar0df52/li0YUxyZ7UPZowuTO5aX7UDIJvatPfOiGq7
OYtwYd9Jog6d4ZWRKGiMAAaWZIYf6l4TQN4nX1qvX7OLXnMOHgNOLWWOgT/XRp+11MnMlwTSIhSI
SLzZAOPCwyY3EzV9uqaN7i64rSHNkb3byemMw1lT3SlYBGBIgVvpk9jSD0JBv3inJzqq9abEFiz0
BmZU/J46zmRw4x8YHlcATnZ3UnUNuMFCZX1zi0W2T/nQk2S/nqbvJzP6HCjz490Y8UDkR0UBvBcg
qzgD3voD460ccPQ8bbo3bpF/YyBlm05NVOd60IX8jYDcYKpWYQdvmy4Qr17OYtTff9TkaXvM2nYZ
Re/D94EdQMVjXJhu6G5NTYhIEZqP7PxsUWXWTM+OLAN7cCtnpBIX4l8dJKnYwNhLkUIv7RiAohZG
DvMtzfpvl+dtW8jZCxn0nfCErFeYlNNCZ1VBhCo8eFfj7zdTiVlGI2zoGAdjcdKj1cvNTFIggNSF
BstSnNgwNH7BsNhejUqU6u+QS86zCK0BJyxWdVnl2vl6MVEOAkCHKdtQTS8nCaS2XRTGdW/+cmR4
ipQmCqwi/DRg1U63gV9i0dpZxaA1iKUsY1StFj9n/yZ1t8vJ4lxJ2Q7NfKLb9hL0cx+Co/6UIJ89
HGvCpNcsdCEl3O3q/32wTlKVm2fxG8qgAURWol8OmEnscB+GS5vz1J1iNR+pwL6gv8QC+RUNPzu3
jO3YQwlJ49mpnGL0IzvN/I7Y+4dvyIB4/uvCrAMm5EAEOokGAekDpTy2Sh1fGc0FNTeQ/DqslPJY
qXf0wWS8ijcUGyL/RqHx/D915dRRrWe0QLCqMnbvvuxIY2GPBvN/iwizeMZFax7BTizYcItwGEBw
vtTCNdXytmNNlf4Wemf/uUbGPfRxpXkA8BWSSUEDlRdD3+1WiUHM7N+snJLqQx0E+0GVmZze5K2E
vDTDFSF2XuZVe0gxOUEs1fngLzM2MwWzbYJMb7CA5MyzAIdfLFT2F2xnt8dt9tjwRhJm7G4DwEps
4pyuDQGopTokejoUXv6LA5Y1a+jdbSPxqpApcdOy9tLudyOcupqRlF9rvMQwM7hNDDqh3i8UYMzt
FX+EJWvPzln9D/yRhlyvNmNU2f5DwsIYOsXWq0sJZGyPIajyzzwmRt+dJZBJdAqBUopwKOLFYJEa
xSkOdaGmOST5RSw/A5b5R75/7STwCCsezft4WzBVD/bdfqr1CxPd0zgbGJJkHe1fkiI9rbWQ5b9O
LnA7zts8mRcMlCd1oeTeCOoA4RFAuaUinWP1+4+LXFxlP5F604YNYB++bGFPNgSxnxs2bvg+/+6A
TaEx1MNB6bDwJbptlXJxFyOUXu5OlgMigLSEjxZc8c0N3HIaHmHptS6OFiHDqAhSXwKcOWUcYos4
10RuBR3JEwDKfPF95bl+Ye6xKshnoxBYmHVJHGczlGEXcs4meNMK3O5YXxZmtnZvjfLGOlZ7ZMzV
I0UPZJD8+MYbmtHATRIQSP5Op0FUFJzoymjvGdb+0D+TuDYEqjsh20Gn1sXOi9zw6lTNq6jr98Vm
fwoP7PTMf0hovLP/DgAmB9vF9Utp1SPjdGDE9N3+cHxIZWioegdBaBe1n8FSfvJFBBQ4L8tbMDHN
CL5UmJ2gfjViPyftNgGJ5bxDQac0jrlxUM2Fxp/zU1ZH7AEbVkxz2kZNUboMO7hL59Yc66OYH8QK
fjR57ifjQslZTN/lbS0Xxmdw8/V+yNfJ0nlUvPOB8y2cKTDc9aBaz0a3lYhoUFv7qjn5nHwSYKM9
bdZfOc+lv22SyYrQenPNnvAt8x1MW8ijEqwFr1nQ+506sWBNa+3V6M34hwRZScFb+Im5tax1JaoJ
PIBnK9NXHbUxfr+On41UygufFpyT62zzLG4TwwfAem7KofBhPVI+u6NzLtsr+VUsiXmG3/Xi0ZyT
OOPsRYY4OvS9rA38VWcJgIZVo+fwID1X7ZZOSnLDX8HyNsr0GtBD5B1eBE7Q2wyAXvAv/B6Muiay
Mk0sry44pJfoUQwmkwDl4Yd+ZNq0VQ8iaIiqwSVWIEljrGOIc7xiL4F0FWyXr/RWzbRgaZJ58Gb0
lTnUDROnCErNCX/0iyAN77ascT1c+Y2E5lTs5dYVMqk18lsTQkQr77p432fp/naZr+MF1Zwqw+sy
7L61DyHEWzS1Q0egZxmVWsYrD8YfNBXVS3mu8LAsojmjZz6KRoyUtx/07NqzjijIbRKgnvpj/W+k
gfdI7ykPvJaXXZg3VEtHewb/4HW3ordQQtUBiWCANbdHa5SfgwOWkV0oNVxKv+0EVoiGBzvujJgz
b+rjIDibQlcff8z9FziBrwALNG9gqyWRCJomEwmsVzlYvzMSxaAxuOLZt6jNOKEchBvOd+FWc1vf
FfFsQkLWtg9FJbm87JZfKUoPvM+eAe32vnZAmTS4kB1vvCqZKqmNB5VT1Lx+E+h+9OYUaZhIcYLS
bKKTFAlOW3MIXqertWKYqjyEokiOInSO6VOYPdHYU1x20QoA8Z9T0X7CMaq8UEHdlWbBiI/q7Pgp
rvvHoR3dE/Z40VBcrUvI9aEaVV/NY8Z/2kt/X5bKjk1iY7YS3E6q1X+ZLZ9LCQgGtn234ONnCgiU
q1s2OP/I8pMjFd3C6YJz68QGsOfc0hz7utn4n4aOl5tllmBeMeyksWAGgDO1ETLrqD7D4zV/i8GS
pY5pm6gG8CErzQE/fQMo5sK+Ohwdcrjy2rx/hURSMcC407YF9miSWLXlntBdDEdPLiHOIXoq25X+
Za4veO9vXd5bY6zBlwjvQ5AegBtWRLS9xyYfrdPP8AbhaNjyPsh+WXfxQHupx1FePKEn3FzuEYUz
ADLmpADUc3WBSuK9Sj80CXEzHnX1SZqsl8t+2h4ZMv3c8XDMnVaPYri4ob5HOVDmMB7Z9E12zFHt
mMTZ0ThvE7gN5Nf01IsTxJcMMvCG+cB7Ig+EHnQj7MnHQAvJ3jd/5p7Bt79MEXl8jNN7nP6tBR3h
ZwCxd1llXukli+BMRZJNoZLWj670juOapF7EjhlBI9eQWSspx8B/UQbZG/n/NEpgBpoYuMYeXKbK
abLKMi/u42KXktuNbsrOrErXYOzyPElRT/uKejF/1kfU35FSbGuJIX6uw6fu0MiVJqik88i8fWZQ
ykjoZU5tKDHnYoolUvQpfYyD/E3bOYok6haLKf1o8WdjhoRE/WoNh1mJmTfw+SmHgNlPfvk1QrFZ
4A4ZnGr+1krW/FmPjn0qKJqYi5k5g3WQacanmq0b+B2HebWrNLFJWLGfRihG9aAalY5m9WpZkjHO
xPKKCGS/1nmMwl8ozEApdGoO7nMsKSCUw6g8MUyvDpm8eXXGHwpAEDuVpokMbm+9J+fLu+e8txYB
kdGny1QZf991Csc2mvJA8VSBY5QqjUgcyM4bmiQVDPTSVumOmH5WbSoofVaMOWU8+uD1IvDVCtAp
0ES/CAAwhJG/q9PsALJpdHN0mK8RTayAAnDFuctB6BW6M3H2cnR7DkLy5jeU10IGG0vNaSpJqkYZ
t4aO7rxdp+8e2WbWZl2JG3y26bHWQM36BO2on3WI+jSWKwQ1IwbBPR+eB9YwgbmVhVfSXTnYi7CI
0hDGEuPS+zJrcDHAlhMpYiB8Y85zEqm65HCnWBMJNpeMf+04lOwXeqy/SsOJDeLTzrp6mjSHhrcC
0Ja5wd+u4Go5qYyZXW2f0YcqOt5H01QhLTvYNFy3xmWLQ8yqh3IgEfe3a0w8Kc59gIPB//hdMbhG
ughJvkPbsfwAjBuSNbsl95Rk1wgEGay7D/94rBW6Y80JOqaJ+KZXiS1c2J/tWV38IMCUL39mqhVO
iiM2gzCMr8OQVrUfKdAeYr3hJR6u4eQCB72tlK93TzPmgd7/cVgyAy1n/8Cn93zKBhH5np1Svr0J
5Q1dABq9TGlu9zNb3kAblLUUCYmph1wfJIa3xKCfqpuuWMBqKXKbhb12DBlT3nDBEnH6SwSnmYfd
ti2KSWfvw3Kh2vkTPYdZOwL6USaK3BZSzu+MnGHMRLTUUBF7FftVS4Mey9577E9OGZAe6xq636ck
Igoyg9uAN6rsCIsPMo74+BNxW1FKLpGAFRiwlEGTykviAK7KMknwWwoy+Z4XzrAS7NFwxfXpQuzk
o8kJ51sUP2OaR4waswW1qjtJ8s2Q97no1koWvQQm/AhyOL5isrQ4GBSltUNy5M7JfsP/UDfqPi27
/iyKv4RXBrDchMCmb7E6mxLnPdl+FWy0bDSnr0UOqrHcY91yEB+SjB+WQHyv33imvRizlsSQUKOz
tWhBHsdrDVD9TvYKSHDdMmiyAM23Vs+s8YU4KsevBuqpzmDP9X5OZQ3J8/L3lv50tbTAFdc41wxc
qRc672E9bm+rlCfBJgIc+6sItdIsXmQuHY4j2dRiZuAI94pby/bZovKPCbw0miVZSEjQBd3AzGMf
qiiAQYMuG3qcgH8YEniyaNPeeNtjxiDdYRUjonFeklgxdMdR3O4uC2JsrAmkBTDW/S4dSPVcHVuP
t6LYsUTuKW9MFNMkU2ra0fzpkxL5luhF9qqZxfRGl9eFRS4yR+AKiYopkctOW0qdzuHgrazYpnwR
jbO+yqXCSTt0RLiSOkIXJHOXn0MMyicOYAfSkggB5Rafb7QFPSEG+Z1hU5sDDDsnahuIViRoZgxw
MR0uKXqSzeBIWGrmX9St9+9J6MFmoaXCVDG2ia5mZe4uv/CPD3ITYq2UhH26zpTMsNevU1RZvtXn
kruft0wd2FCYQXYLy8ZIsbIcZ75yt5PzFwsl7Tplvwr4ySRXJVUUNTM03J8BmuznhcUMVB6crML2
4ZYgNO+BbBy5C6oS+yPFMaGz2lj7DLggryhPImKe9m5QJVsqKCMlWe170s3Q9kyABj2y9Ou5vlJD
5TK6dlXmUmzzmbD3WhF6xlI5r/SEm4IlAX8gXw/louFr83N8Q7DurG11OlXJ6rycYeuGhjPduQRG
84l/Pj8HNyO8C7RS0ifaLWXZeYuBx4RLVuBTPhRpvuiPvxzbCNvMCW2Ab2moG9MXQr1enZ3E0ZUO
CdcicRuV5mZCzbOW/XCedn2/bzBmGmT51EdBFMs5HsQ0IRs6a8X9S/j2jCkjrPDB8w12eI/nIsCv
Iz95qUAIcI9phRTvx0ndVe50UDkkqW+WFpIOAEecv05LbxLMXoYf+w4XZb/SBmqIunXiQ95DerlE
2xs61iX8n2QusFhCALhWWvVMmiJJTpXq67f9+iWXPTEVJwsCSUpI/DLvMWSHe0aoLTwZVF2+KcVi
IKAFlA/5xZobOlYkA3uBvr3yHxjyWIWLpsShZcqeXzl85FWf/+KJybhjMWGNIFJp8MvMkPYaaKXN
JLWR5MmMP6WNnbXuZIppvNJF6wGWmrdlpj0+umdpe1nkkaC13nge2ya4MLoW+fNm3UI0YOZ984su
YuOa+jbuzIv0chANVZU0ypYMHgo9a7Y8K4PJN8f6JhMpgvP172PxbMneIvRwS5XkiokFuciwOB34
m2iFFeUnJSHRDtDgrJ3A2AJCIgHvduY/CkRQL9jcqJf9BoSrNELJSEx6uidp6Ze5u6mSmBu9Me/9
URL4+94pQZ9P49NhKvJO39u9CBk4Mf9gXpXDn0AFfjZiaStD4Pg6bfYHTma4bLJcfDZBh9HlVCDo
ssmvs1Whdo+rYQcPJ75llrk5RRsb5z6rM4GpGL7XMPPVogkAhAvzSuLumlikHZsibLFA8aN4vXhO
07PBQWwVqE4qIFWRcYPwPNCQu9zE3v1FRKTXZluO1dSx8L0i+5odjtATDgyef7aEIzrMkSE8gH1L
EhaWcab4kPDxWsUQ+WgcVDm65yP9e9N0SDtalGVa0FhVe9tyfYClAeoIPdIVPd9Zzb7sLEYQVyGZ
a3121HAayLQesKL73NnvjkYo3sgEy3gme/Au/LIOjs8071s1x894DbwkWEdcVJHfKc6rcJoIN+mD
UB71ezrgVIU3e2sW1shelrf4T7jZHrK49Z/L0pdUFem2x1YF3X2Pw9X96pkMDmxNfD51iy2SWZxP
Bc5K0xDKS6+QV/jXa6nn1XKuEu6a7a2jhENVMurJBjL4dE7R9zPSr/XgN6N2B41sNt88k06ymbrB
9b4wz5kw+IOl5O6k7tlJLEez3DVulq64w3frH6u+qT8bVw2DkxLNjwVxmjC1s/qkqQzLq47NBRMu
K0DT0ogcPj1HX8HcbeAi62T2EsYu2xaOUN9u4kxZNFLSrI/6Ouc94y6CbnvUYXSuHd3Tb3MGMNPw
eWPA5n5zl6U+OXX4lcxzJr8NiONLYTsEuWCwUdLyFAQq6Y3gnO25By2R5Ntm0SgwkMHibWvJRcTL
q3bRmd+3Pz9Cs1FksjNa9k0NnuKQ4BVTKbjlynYZHlgnpikz4GF68SwJxaIiP5team8kDE5kVHJs
IzODsKi/HpsLck177GSHuxfgNwLivGOS876rHgBKnCM5K15NNLIq3VzTGGU4YtmQClrAWjTYg8Wc
NK2fEP5BlcI4AID/24thhNrkCK5Lu81gRnCHDbJPRzGIsCiy8MUExngfdZZUI51Y++cgjUHXhpam
pXwQAWYTXHiY03/Y48tg7ClXFQo8LQodJcya65ot/qKXH0+XmSxTw3uENSCdmRDZeIEEwVvakgKZ
I1nQJxwGlALcCjDYts4UlLI/aM0FVnXdH+L/yrYrL727xPb+aDfoBp1yrs+KYzJYebdli3vftxPt
RBcoRDpOAopDccM6Um3NyH4eBngq12SqN+X8fdicF/8v038Fwhx+DEy0CX/OTaHNnhlhnWEHZekS
88UtujQ7nIeaxQrWZuK3RYxNp7L+bhh+TfKWEnYYrPDjq60SlrSeBqb/LSMvZ4WMv11Cfj8/XJN/
JIs+LX84129I650duYGlOh3hQWKFqYM44Yre3DEkbQNss4EtaimTuabCjJx2sAiIRzye/aqmC91b
L/kA7rLnCJ6FSObQK6UziNrDLy27M5hmYZIeS7ubyS/yOt4sonABx2qKKJJ7AQv4pLW4602jmzGj
21c0TCQOZn/iXiPew748n5dymE9FDSvQgoEOkx/L/LBE49Kr83g9h89Us+3+Gcs4/ygsM413kTPJ
eaF6e8rQcUosfLX2H9NQr9ZRQFA6nU0EP5d8FgqfdVaafPHzyPnMGe4EAw3Nbyc8FahiEP1GtINE
OPdGnT/CeZkCrcMqmlgKpKtPDuBQJxqyAXDWvbrD1rl33WfUqKJbssUDTvOO/l7xmq15wTIyTMcl
yricWzLjrS08qFpsD0oH5Lz4XrXX3TXZYAMZfypr4umM6bzj2IDtPSLZdQyt84jyc9WJWsxVUk2N
WKptuEm/n8SjZ1H0ZP/XdhXHzoucDyFiMRI2aJywMzZzH6xcG/cPo6k65kwp0CWQHbdInIUGCPiX
wQ0fX+bcvbRS72mlNpNfq2hmU2xN+MJbHqL7Tmy6Kdna4sgC3Z38nuvbH9o2IjZtGi5Q3Ke1HRAa
eAKEfkSb8VLpORaGe6fRpx4ERUeTPHwEjxAUBEAYMBaV7vI/SFLb/5pBzzCKf6AKHM7Q2aM4N2Lq
h/rgNE4EzKz1l8XLWuFQrwiouW66Vzck34owQomPA1LaPpmrMMj0A9KbdzCb5+7sDPu4rRzKaEzS
9tg9TwKv8ieqDCy1T5eiIiymWqL8uyBTIHd7Eq1lh9RE31ZMbQ2OxDVc84wULnZrw5guizQRzj+i
Ifd4NE5nU/Hf0oItPWok0+Q2zceieh6anWGvTuZ8sGOOy9F5s5UBiDaOyjQfe7nnkWcGlO+mzjM1
9z2ibY949MDmWS5wTsyPUprPImeMIXzY8DEcHz51AwaQo+EPmW2TmCzXlImRzQXIuctw2MdkLUVL
znSf1jDvFWSS7nIILFUF6tHzqs0topyA/nvyQ0qguNDQBWWZUD4uuJB+/OmgM4Xc6ps+PnoWydsQ
tfnzJXAg/jyx/76knwvgYOzM9En8w6QNkSRQjUGDgLFXQ347ww+0OC/AwdB8aL/5WLSq3PSYpOdE
Jggh7Z/HBTAqJQDPw/V9wuBvRD1b7M+u8+iXe66nsi4SzTlFH4sPhcehviKPa2iiJrq0OYcg9lTj
xnp3DtvFmvdhYvT8RGnROPuAJREX+83C0u6mtuujpFg9Lu3wNLrC22WnAluADzyvNxAFVMuofK44
1CUGC9NkjcVlTVhTmhqIv/B2vj0S6Fk53XjCosENysaj+ZseiRt8zUjGExjFVXzi/29cA+NBIdEI
KlTp+TdXr2bKAx7fuEcUsZabSMHOax8KCWe8Wzy87unNWtXe0pnWgOjzi3MOD5SaXbitIlgkYjxF
sCzYAo3OGoRZ7nvMk2Dfjoiqk/b2sLNPQuDwUl1Yz8TcqJ/PYsZ1JMRvetD6PTmhjSEUzTjANNho
u3SqlKwinQZYFQvHXNry5KXn1koGEGIBX3YrXjE3O1ofipB7LoRBZEDIU9R5uyUmmjyw6gHT4pwC
nT0oj6bmsDy34u/gM71lsO/qXC4zUmuUy2THqpvThEx3UxiWvL6SYAjdTLt7LqVnuAYBkDSovhWO
OGpc+bXHvlX9mcUxTeJVHMTriGJ+M3iN59bSi1UGUzajZuW4ujv/bfNhDENkcL5s5KIBB1sIsAfg
k9Jl00v/PiokcEFz99k/Qa7SDf+gQAC3IqUdaO/LTJaNj5esyAJLGnM4hQ1d1p5EftkxUbVQkHn8
6uSDU4ghd6wIzlEd47+tawHMGolQkA6HT9sg+vBlFX2zIHwFNCAIerw9BMBkQ5ZrQWWwxtysE6wl
G3MlDHXUbVUCE8z2Bt7f7E6EeKs9tODlT1xt+IG30K4fUpTHm9uwTl15dF1FYW8qNB+AViRbU9sd
nrTtyx/8WTjW98RYBIxTmXn9ixN6OZ/rMWNCh6sPSmB72D1r66gQOXzh4dnfxv3vM7n9xeLK5iGm
xt6rygDqd2k17cHHN5y/zDGY/To2o9H+8rrYKecvpaBG5iNhNsp69VIIf6Dmfzw4/NMX1ZbwI8tZ
eUSU1oAIABeneMpkEgUz7EM6YgBrKV8utqnJR8bQMe0D3mnBUujpc892+cajfS43rmzhOaQeFw3E
ZreyWHQD+wvhxENytVpSD95sXJb9e0SP9/lDmplY0ztnVUtZu/U3rnQBNzb6i5dgd/Ak1l49NlR4
jhHpcT0PEzV0xf/TbDPTkaxrKkuKHOIsaCCn4TVgwmYua/zusqq6Lqh81Y4elbzjk9CkoSSCJXlu
W+R8lrC7rliZkk+6ZVp1/6GhDlKjgm6Xxjkh5E7OJyUj3H8GoDlgYIG0rf0Ad/fwiNkVY1kLRvxS
D3r8UFuYOrA/xy5XELQcoEs1dFC5YABZ+MIN5H3CiutEOePPD9MFpm+fw2IZY5fRoBR2MFCVdG40
sPaTcnXlh3VNL1ZoH2JeQHvpnvzPxhGREV6K9ae4/UsGQOdBxLQK00cp6j8BHZkqEvy3/L7XylVz
QkaBrExrbkbbVT4Hvy7PsgJlwJMt1AzWA442eqpj03AD6QtH7+D7/hXFrbZUcxCue/GxjcX/hWfa
TjBgWduF3BblB6Po3xyzbmcZkDW+pmI7xw90dWFhw9x9h2iCpKM9Ln0uFy+a3+UbN2B8VeCzXw1c
KRsSAhcnIZNEm1fq8XT+Dv+pHFiZ3vtS5q7jLikw8girH2IdPocq5Lr8/aI2CqAlhlRrDkEgpH5q
jwWRzXu49apVgl6XvHxqACSA3qP6kTsyqh54WSDvGmG/FKfZznH/W+0ucBX3wSTTWDUI+FQ/WLKh
a20dDIEY4cmNMx6Rq8nUHh5VjvO4ZDnKo8x5mqYjpIPo9+b1bed9lP2NhqdfT3OpA/mWGDBkVnBZ
+LlTppc49Nb0uF6p/ZMvHvahB5g7OfzlVzMhgWH7UP9x6YQkub5E14sv72Zk3hHdHID1RzKsXTyf
9zRGyeg1qx4tYkGqnRwKlb31ztWxlqO5coFCqF6iTRXvKTBy99Z6MBAH9/ZUg6QafvNVZEoNFngK
CrRa1yIWJnaU8uYHvg3wfa5LDOvB7D00Ktahs6YrCPkrNNqAAoz0xvF3ydfptgPSY8pXdoqCy0E2
1E7tcMWCii71BgLOJ2IbWVqaLTg+qWqBImHGuqRYKGEnHS8IznEv2nCK/fK4IQa0rO49pA8TzGIf
MPy1Fhb37KhxaWE3u6u423lJ2Yk42G30xV2kRBD+ywd+lJKXu+XbjZHUf0PL5pfK4EXAepBLDaZb
VGd93SSjxbn39uaKFWcV5eFvta1jiNbuNyEn6NPM/MPmvb5+GmoPeYXD4Avzzhc2/6pkaIIJUY04
DSzmIbdy3FP7LkJ7MP4o4IZVRKfMKMl5+SOmrvZMnwBeL7efbVsGgrVBtlFkdX5AMXZT/wKe2VWJ
4XFLd+Yzw8iYhMqS3Pl5r9PGUyZao42d8IREA16xv9AbHBOaznregVfad8iO6ABDNcRNkRvCB9NG
GxtqG3vhUluWn/q/jAKwPXkzImpc1/yUJMHOyt6mfipOjz9vuzDoYOB0ikMo0JLX8adZXpWRdAg+
wyWdFfPqwnl6a02Zh9+GsYTPKs/MEjvKvccTU1EQZ99OgfYWC8sfYDCYfBToFd+lKOPiqp8kW1HW
oQoc/T7HUeQiwUrRM6VT4nXc4ThSjD243YMhV6O9r+I9AdBRJxkrxnH8J1morCe3drYJ/d8yFnPY
1XWkpd/O4g020N0IFMTmNk0oCcWWH/rulFIJ5w9TIp4z2WYvX+ixIzHONzq1PMH09YMdu2jF4JL8
pnaxC+xBd9vHRy9clRQs707sJ+1+F9lfku1jHPtKC5od7FL9tgLCdRXs3dVfCmPS10UJ7Hxcgh5c
JJsle95w2Tx5cIIGl1MFny7+Le091seCOxWRslbUE6Nub4zUrNOze4HeMIuZHThSjLz5LVlYu8kV
V9vzizt0gnLjaHjV9fCNvMP7d+HAoCmoBs4hR2O7NlqCsaeccz+Uxz+LhfPyAyGLYXWxwrh0vlSz
PCoGItzsWC9sfweWTT+hjbyPgvlw+QOpQ+jgEpK2F0ulPXpSjmHHtc+D1O8tTRHDgnvFaEW/uK9e
P6iMY2sIA0zUCISa3pWq63DeWN+P1P8BHMzDGpTMKCDW4hwo0u/DYR5iHBJNZ/hCaW0YgvzykIhP
oyhMg6PZW23GO6MJdAILHy5dpwS/NuOgkKe5W5EPTcZVk73h4ndHMCyle8XyBH58Ya65JvW1TJdk
Llc6RxC/HayjsSoQCWVY/VLpa5pvtPrai1zWxPzpyj//1HV09GC9nAvnp2W3pPkuM3pUNi6ef45a
n4i5CwQI87JlfOzNN7JOqsKXlXfDtRy6W0xAPbbV3/zazdbox+c7Yc3G/P5GcVXxE0F9jN1vlPo7
NzJGyWBn5O279AtbunKdTT33W6olpsYnmpycJfq7af7H7YPckiKdQa9fTlABMPMjQ2QMnhyUfESN
sqPjcE/52k6z4A2N8aRqKPbVVnnOi93QafbW7glOnKd7Q1S9Reu1n3mYOMUOoPloQFDZVHRrzOeJ
zC+wtE6mC0dRkfMnchi6926/bpgT5tzmfhI4MuVYOxNN7RvZijrytTqn5zRdy/CB/f52j+zxWx5F
DLgMwN1V8qJ2g9qqjPxJRzRZMqRtTiR4qBPVaD9bZPofeqmnKmiA/8oeiXsqUbrwvOO457PTQuzQ
5IrLoTOIWUzIP3SDZLvygGlnOlO0SV5O9e9Zb2OApXbOZyPYarNTZDrksI7NDRPDBr3w1+A6TywG
qHzZiArmblHU8l0MZFfTFJJ2xEVNHzkbiZ5WsE6HoIvzxSrS2wdVFeFYVD6Kt/kUv55DtCaBoMSo
MLUGL8d7FrooxkMbCKD9B3hhqeTtvx+E2p/fWuGJPgfEdtfqof44/ExmH7u6LVGKywBYCySxpWT6
UBKcVVdsBzYBiLCNSzilt+Jf0+RqQ1WsLSZLqssnRepTxGhWvhQIpxRCQrlKbw0hf/dyXW6JZya/
aZdeJjmSBqXZ5IhigFvEi7KdITbgXLOhwa/eX4wEXRhMY/U9iGlwjLXTuB6uEuqhQ3KX5gbG/kKA
H9/B3FHJH5XAv0iVVt22X7wwEluD3yYn6/frAbR1q+1m/emefu3xfBIk/9Enw/x0pP7/3S00ju21
vzqK6Dpz77x18ZsSuhjjGu/De9PCO5W5oYi9Bs+LtvLkvP/9X5t6j+uaC5cUor9/G8t9Hgtrlc4o
JbGzNtG9JQbniI2//e17nis8DPwR82GFHwqBLXLakubBUlsXiatPSykODjIw2OMbjUBUW06cHm8m
4hi21Onav15BrfKJcPhEbJFE5hU6j+PIiMKlQodE5yQJ5pTAPiFZoTGqTqiX2gk21lrPheccpxwt
9612HiyaXe6CGBYV4SssfjPfSa8YjWwSr2FeBPpm5KhlmHLOIKYwVf+p1r5wb7fhCJ6RAPe3aqNm
Kllojx6m7vV7MYCSg5BIZZNghHMT6P8/NIr4EMfttml4yeVl+EXJ2E4IznJtFV071sE+s6usuhVD
DgWTuMuIGne+9NaNuTNngHrXl+RCSD9KYZVfTRrkaCuzINuDY9jxTCqxI2Hu0RY9ZebMvsMP+8Ed
Ue2GF6xGI6q6bEcNvRjU+wHtAHz4zYer0Y5FrQ9PydG7GRk+pm3dmroEZ1slGWefmYGfY4Auk18N
hlt3pBTjJs+5LtVwAhsMFhFCWcWrusybrzN427jMUBcX9oGdQs7VzgWxw24GfmTlT0Ng0yHaLLX2
1JBxeGYU9gVcOc4vcSIpuyhGDYfsZxEvAzO8BqFz5GPQ+TbDflyLy0VGPrt8C5XEnOcZnGNvTAIC
+yzV2z0IbjvmiDMagyC6hR5jBobImRqMtvihV9NGIMx00rF4bQmFDOVQMxlNq3OyG+MoHWRxCMd4
0bqshALk/sswDvaz4B3nVenfMbCXZJzW3lWxOmjJM3l16WCMq8w82SGtOpLzSnqLoWq75h5Qs5Tj
j3ECWG+Fq3Tc8pfhV33gaVNsXehSI5uvSJ1Dtft/muKTFujW9KYr+BY3XH47osupOqLk892IT8bR
RDN7rSdOaPWG5F4dZwX7oeuBFRyHRJI8QFvvnhFxbfdPUsCAoWNI18ZmO/hrrFZAq/L0EtWKqPcG
h9CHMmxAxJoxmXvagm182Qzo/jjQRqUgycypqsEAHo6Y4OatZOgGitoQF6HlEJ6paKS1zSFNOozW
I0L9gF4YDTwxiOsCdjo8AzbLM1q+gZlzscmcw8xCt4MHjSZA/8NHe202nj9esY5a5N4pUcglRLzm
WIZxkbsushYS5bkCDxyOfMm5fid9Ol1PGF+AQe9qUcbKXxe0k7dyFtyttgvBMW3MdqDKWYC1+GBz
/9nyigSiomJJLG+bWkzIr5Yb+x70E7PEDdWkIDjAF01RsckfoyJ9hizJyngdF/ww+A3NFikw0iNZ
fP0X0pLWgik0PVsKFj9ZgcB72c/dGjJN/9Xmyg1CbtBsfwXdbhyAx9ZDZ7Vd4H5Kbhtw9f8MbKN7
LJ+aYoy5B6dXVIvydsv8mZdNgyt8P6grSCz1RTCEhf4bjdKMRVxNUtJza59k2N02qG6OhVyyBRLE
hUhBCvguQyihgKnQWuA0rg4v94I5DDxVtt21E7MSUPUuI5Y+KWX+4Kv2kVxuDYKPmtkVlPPhq2Z1
dvCCh/pswfrT23dKGZ0DsvCbajicsAR817eTT/qqNibzjC4z53ESmEB0vGl2SBnwi9JLRr4s3xZw
UgewcFuKga/H4SrVUxhtLmWxh7A3wz+Eub2iOiNYjPCQAR3hl11/dOefJ4B8p38knEI99jtzjtQX
gCqBtbf+VdtrziwRp8qa3ThRLn7PiiBjDmnrm7nY7TIJJeOSxEGNgd2COH/R3AfATjTFV8bSxR2x
BNhXtU08OSrXPPvV1XRiO5y5tqtaXRPQvjvjo/iOJt2iidmKR3k2wJNn/PPfH6Ye8etiSwv/hCFO
zVqYvNp5MBXbkzbz2CqN+WlhNT91TUwI3xy0MWgLkkOsCzBxY02MviKnGI/B7vrNXD2JLwj6MC17
sadvC6hTo3YheB9sXR37ip0r8zFrOT63jq3S/CE0A2XEw6d2HEBjm4BW+55y3+DNcMV5H6FlSnvB
fSQLQcJV0x2gtzSOWLEIvW2nuKjLHulXsUXLU5WUu61XfMRWw6PCbdvfSR3+eX1S67glEDjVkiHW
HnZMaLozn/3cbamoBzxXHJd4oRrQpkNaAQsWzipnbX38NWFW5F6ndDA7BM7FKyt1mU+06WykCeNX
q3SPfn74VvzXwSPf9yvBKv+czbkV6m5RWjgsAxCKKhOuTlDu1wqt3P6wXpCbsyUGcpjbOB78vN7k
RPkUQhjskVmhQu0CZbUtziLjiakf0lKNvomGOihnW2tRJoxv7weCc/qmLIsHalkgE5pkwq1ghgWV
YLs8e/tWV5OQJ2QJ8hB8oAc69AdP77XkFy68tZlRRmT9Re8pf9nzGO/sR46QsvZMq6pvab9d2aDZ
ZuFGNk8Aw6rWDC4TnMAqcLJPa8OedEP8UPxz53x0SmSnbBf43TiByfwGaCn2RsxhTZ6PBkI+agSA
UjviYiRhCkyjM6ELR1EqJkqoWGlXHdYTltIf60kT5VJSt4jNoCBM8PM1gHGL2G/opTeDuCGxYw4r
0LJDqa7ta3UXd1UvACtn2E1zOYXH1gfJI02IRYWc6BbFfsk4X/bhqk/2hRSM/ihfVKSRka5jJVrp
VAoMd2T0v32STmRFrYovBIRPEtDKNTmElgx+buByV9gImxS9FlerbFbclr5z3si5YwH+wETHtWTQ
hMUGkiTIuuqXj2jSxQGZdmjWUtEeI6lIVv2bv3X437ibyTKJIBhQJHbTTq4Mgp3K8nY+zCB/8EPH
CTkrqAcpv/Ciaz8sTX7mvBuhpmGWnGZLN0yA6EpJq177UuMUw8U+aL5RqBt6lhXhxfvKhFZm9dWI
C1NfVFKMdnQv9HkcjCuJ2We2nlyBW9CG+6Ase+2112uEaKhWiI1Sc2hCCcIcgdjkK0+fwLQDITSE
gh9bGiJxf0anJ3SzmJqsl9ILb7c/CdbkQn9fjelHFe5dSX/5/WxAxB2pwA7J3E/fgGs8JvQ1hWwf
9LD4FsbSnAATNdxXax+TV4369Lwoflodh287bxdXcQKTy6owUg5lNW/CnzA/VZSuP2ST1scJz/G7
4365IZfJp8cB30YnsH2F/wjHaB8gdcg/1AJp0bNze9YjjZR4qw+LKrtWNZY7xHdsv/kcGSwoP7Zc
36zTyHyz9c6ohrLSJTD2ETxYiwVW+VgF7w1xF7M79Kdm4Coa4MZqCSPTjqeH93sSWculDXIwcSGB
AipafkcYgb/ah8gaZcjzyt4U9XzYEX5z2tHEZz4nZyPucn97uRdkLI5Dn6XMmFRuoF5D9Jb/0CTI
DMR2TfyROVyxDFe7Kn1IDQry1a97M4C2Jsiq0797oTQm0BmlNA0R4GUZM6Jqal+onl8hNloNa6P2
072h4d0rRGn/7yoBvZfg5UX3VVjkXiXOyQifYJuiMcchoTR2C1VFTwPGFwLeYfEmbcxR3Qc5s2PW
ta1uVBsoi1BDuLuuiS6TLwr64LNMeiXMYpaoAzYql7WUsPyQt7iahFORRnSVgCwO0UEoQ00ZUiS9
uShChpj2DGcCRX6oQt/fyY0VuKtzYbAgrQbD+y6P54AG5kLlhF6KJvhfTf92eTs9OH7ZCq2yxJQf
bzfvPBY4el1BtZLKE6FWusZYcaLwFzyTDCopvGSEUiBeZfRPTrN4igYQYa+xajqZfXcksT+zkJ6H
8DqAJ7qeFbo4joxD2dYWTTGu8wj1gVyLojBVDOwQTS0rx+uS+5q/tp3oy3W8WxIkzmlCtO73qSqT
R64zx/O8yyl0exW4jzBB9kbtlWHAneaUmbcBPqM+fCbVsC7rNxYJoKaiftJico/KRcljiUIn79Rm
nxdk8nw7A58GAf43/WVChNIt43ENLoK2li0wUsUDUDIAhAyUTecLr8yz562FrytoX3YhzLzvDuNG
OJExPEWxeFCY8VDu9YJKMjLFytemnhTKiOsfKRpvu/R64Qx8ao3/RDOH/ueHQU0DrTD/D3mLI05t
RKD8vXLJetfhJBVZAagGsk9NZWjc7AwmCB8e0Mhf0mbDuo413Pi0yDZl4xyJKX1Dd/2yl6n6aiQt
tP/me+i7Tgzp8xU+QijK+wRS/Y6FcB4DfG2U8NZ37gAnJlxW0LqqoasjiSWW6AmAcXGETA1fklYL
dwCaYuYOLvp6yPz7LuaZ250g9U2Eihyhlttlp45xMzcQ2Iv5PCpeSppTmv5XHQS3Q7ljnVoIOfXm
NBVG9zFtaSvzcE+CfhRbe7JVkiutnZiu4KyoMEcIxleB3xy97fhyWWUYk1aWns26wB/D410Y2OJE
smW++lv5ogFEKFThbNRjn1cmpPn57hsVeuqIR2pkD3gXfBjkSr4BG1WR3OQ05fhg0ygavZnukG/e
5UfrQgV6PSFvDhouRAcD6j3lZ0KOhBQKv2+CrsFpwbP0hXYgi4y88hSyS2YsSP21owWo8TALvlWQ
1eLRGaPPz2vmXA78mPm+JKC0s8ieD4f/xyHYhT09YOn/NSMa7T0UCD2CzDEOPVpLcnbQ1la9lWSi
FHKcaVReQzJL7EcSjt0rUla2xi8DGzvzPcYcE6H51hFsRTqZWkh7jb5keZOqh2HPkBiMpTS5O+hq
AHkHNRPH6zv/Vi9VEllvR6YdjB+HMq7PpD54vu7MAdxMtI87FosVq52FmuBMhDD/6ZQPmh6PmA3Y
QqzvGHOVkq8c77PE9pv3buwtsvh6q++cZOx6q0DUj0dNm8CHoJ8jMCA30X8pgLY86hfx+2TvoBnt
hHGNyknxkvm4WCjxpKlUI5oQTm9HzC1STWddOVmT9otoqqKBMafKEoMVy5BcU5/VO38bEDkoXHWL
jYsDhq/R/Gl5hmcEWYDnQgEohVpvujW6C+XjIutIUvw6VMFqGOQN/hMEmnsrI6zxDk0mXwq6023J
scFS3ofpSaep8a8aitgg6d5jpdJIDUj4fBBFj0b3saER6sGgAsdl4/FYFk6z1Mvw8+fYRb7Md3yc
dIq9xy9uNT9Qq3fIJRh7CHVTAvYpMiukHyj6tCL+cJ4oLplF6OE2IHPfH9sOVf6CzlRv8gsmfQ0D
mYd6rVk4XrhXfecN8+22laqfw2QfYQLV67W1/lZSXThTnnTuhSLtIL4O/p+5z9LueKss59MUdgsr
Av9P13S6RIhbFrNJ6fRhwaTC5pquNssLTeMOCD/4nqccMMGgtLSBHGt64F6brwDzWsn43QvL5yLn
d0yX85yddGDSQBTfD2tGTdmyQN/edOosVsteCRuz3aIsjGklN1hSiePuvK4iJK/Yc6bH8S2j5b+y
VZgW4rFuG/bxEkL0ZVCKfiTeiv0C3t/0hxPFsG/oAqI0oO2GxSpc2Xb6xA80rjs/rs/XazX1acBP
5/IX+rCOxzhI+9kMDTRt3vplh88wA9LSDvJgLR3+Z59Q/b7nQI+UowElYtW9hVhbs5IgumyKm9aR
nZQJeX5Quq5P1ZQm38vEFyla2MjOgASbl6/fFbD9+Aa8CWU3w9kTSC9+5qCT9DvZlOHaqJN5tcfh
n7dW9Y2hZmfVMJ9jK18/Kbog3emE+jG7vOcvqjfRdRUgwRZ48lu91cGmXuAc0CSfrZ2odphC070o
YeiKUZPLGEn5FZK0KcEll8oeU0f0/nHGLVFTciTIs2dVDYOLjwFNSugs/KZ3ewdMPMukplOKrBc+
cXcXoT+pYjQMlIcp9mReN5yef2aEEuHT056IAaXQRWBX8EmDZFi+ID6wRJ7+ZXDtEitw1xLM8BJ4
rW3TXtUraYFGI2li/QGwvjlKdvcVbLBwvLOBJkdC5b65P9AIzq4GqA9wFkI6RWDB3J+yrtWfPFVC
MVik8jnhyVyEwCvf2In+JhMBl/7EzotWnLwOuQ95houpWE0Le0fu5p5Ut2SdOhWtSUSgd88PMqmt
iI7hZGHcN4EH6UM4A//fgNPerJjqLIhGw03d+p/Et23Kn+dAq+fDaw70E8cT4fg5oW3LWeXQ9R+c
O/yDhPDR4n4erVxI/GPrBTSl5p9IjWS+u6lKbv8wWeCz3QvM6OEjWd2WhaduB4NYz3NAJJxtg60t
jTDOmmWL6dSG6Uv6ze/pbEqrlGHGWfSSUxZbiTVZYDHnMef7QLEjuquJsVhgLPAVlbrCloYUx1zY
PcEieHIup+czCFCmm9IpEb484ADNke75vIdb76NZ6OELgTABBhLU8IJAuQPu1lTCL2y1NxWau+qj
rVBVs+oK5K1qHoRaNXtEMuzVK92ZSACD/x/1vtbtaYuaiUdwz1L8hLMCelj5sK2hzycP5lds5oUS
Kc9XUdIlG/Jy4uN3Hcz/29GdbBD1oBzycoVAmeclGxcnfMXTnHjgup4cLyVs2ddOHFtHqUPWprx0
jrqpEKyXKduGWwDW6rpQ/tINwSvXNaleoCOhdkLWfw/5W5LuGU70mlD8iQLmypOPVjzv16JYTbS2
AdZmrNAi1EePtz0zTPuKOxwdcQ0hOGk0SRzOiQBq5nfNHavT+CIiAGO3PFpI5wBwLX7BkU5oNA4w
/c1vVQeuMVkaS/QYZs0tGCEZ1gBjJHmRIEa7uvDSb9YFTeu6VWJsydScYehBHcPkW0dUjgiop/b7
9Olh3ZgDDEXgffrs6qcEGvxK176pcyOlktX0sLcGYkCryZZw3i4wDz9FLLiS9+wGjasbBtotQDeT
+/PUQARSDozTEPZPzHkBtrs8GJJ0dpUCb6LktsQWHXYjBaL3Xd/Mg9tdm5e/Q0kyq5/Nkbet928+
tM0zKEK0vPmkC5Weudr9jdr8rcql8PEDKvIifQ31m6aIbw/x2cY2eUxGnR3adFvShj98ehhEHJSW
p5Mmj8kzxEdTWN/3m4v3DgWyxkFnRcOxa60e65qUYAaaZPx67gJNtByNudb8H40CASJufORoLk85
UK9K4K5rXK98mhuk6bMMOGqn7weHS3qgVuFUnQh0BojHsXBODr8Mrz695kSMp7aos5tuNe6lholX
IKMpmcELNsG5wyafbjyBJgUksI8iBnrjQF9sztUwAGcj976PA/2+vYDlPMxatt5V8ntoHOoqLNRq
WPVA+6xDwo1yidDv+njTGPz96o5ZzyFeRn5xGW3DO71nfQ2F9PM6VsRdMxIJzAK1oNqm92ZRVbZs
XdtrETpCPClNSDFRlfanIqw/I44xvc7HZMEh6FX6leaPh+xtwbhpzD54/ETwi092lTRqKlpSrHGV
zA3JqVgJko+P1xE1ml3Av4+9de6079XL3nRz/mQUsH6IDlhGyPvuqAwBdHwPbK1BfE6x58VB6NwP
zfZ03hvkx3aZI3fPr+47bL0vGTjPSs6FvfzXH/70ahWfZhDM6yPmtqM9/+nL5gaFQyuj/mRyQcEd
XyRFzjsqvAZLjdZA4yBEUvDCSv4lNsWbNimLHYv58ZgamHsZzjwSgXp1L//3tcrPREp15o2KUcVj
y1SyliY7luwYaJ4NOOzPvWIvEeel9HLiIB60xhBg9YlLddNIW3yglxBitmmSxkgACAyM6B7X4yhW
+279sfV4ICnuDO+UGWF5bWff9sI7yDPA2NQ1QnY7qI6OlykYeDzZRR3+Up5jUPcfGfVs8Dr1mFWJ
KgBRT77VliN1Hy876baSpl2rmqv3UgVlHZwyEdAKKulLl0sC/9wCoN6EML6CyN2+zzAugFhC2/gU
5jQ5Vwigtp5IYnYz0xIYNIOSiAhtKEP7B1Hi/zqgdzcQCrO5cVWRIIF+VxTSAAyH+vVdDIG7+DWI
zQ6VzcGtogCWB+2WgPcv3nqZD4I9wYaN1MUo+XU1vSxYsED82ipfCOGcOsAHqNBdOaBIdCd7AwK5
e5f6FjxXznAiloeHeZe7TFsLTKs2Hjp7sGlZWTuoi41IJ8ZSU9YHxC9wxFC3+HSOclPxw8jQgvet
+6zO1ACGq1FE060FuBKaz2LTq1kp6xT+VhQcVYuiOp80QTnDX5xG4dn11TMLQVNivC8LyO15a+5Y
/TeZGbc4y/6yhp5IJKeP6Tj1pOyT6pPJe5QIeuHmQy7Kj1FDfLq6QQoJurUpZ6pC6refh5dHgBo3
MQW9d2QwlQEZeaoOGP+j67Z2IA9BCXpy9J0Z6TcflEs/8uf8WrdU5hE0yflRt8nK/RGJwnEcvaHB
Zi4oZOT+9ELAomdImTtnUg9ml328Yn8Qru8kE99PvZ4vHtLyjqdMbkbsIsxuQ9rfwuOHfQGoy2+d
1EgaH37dtlECEvbhyOIatVFiLfQzEOWjyzv8kIiyno0XSBLqEHdsQ8t99kZdA1ehiGDo4jQ+GZM3
IK34NrdWUJ5QMvM5Eklf51ToIYxqGTMobphgGhVq/mYNn/ssUbwh+xg1tM54mFH2MGyPt5nTFH5k
yUNJhnIZUO/29dVi3lO4FfpTDF4eCj2l11xcJwBIA2rL8iHWLba8m/YCwSb+IlkS3iyIsfmoHZbG
OdK7omFR+7bBk/2bP2Q9bryoaohLrIpzqVnwdcMGLNrlW1IdZcgIwHFYctoK67MvoN82ZD/Amo4i
bz1phUdu6TbjKvx1ZaYduSnAbBqTk7kY3Oan9COqUwTbwfJB5iBfRxjBkpDWx4SCXWOUY7OUE4FE
tve/hcKAc9ve5hIQ/Fs4rZHsxPytQ5pN5016HC7FGfjqvl1Ac1mqYXW/1HCHIbzNBBWJ7SdcNY9N
eouhOAPHw1WE8kEsPHvCGVPuXupRfN8LhGF1j4/XuQQtcMQ2moyzFdgSqwY+I6QR3hl8aB8R+n+6
E7DQVZ5ohoPxpwzRYDGdQJsTAfmEU/+YdADjqyErx1p/DPV4cKR54dNkXu1q3/xH9karnAxR7lK1
IGynx7Dq4ZVZB/ev9BFaTHSuqbEXHQRPYdfNXJDda/ciLm7ftWYLR1qeTXjxLx+EZrYFd5lCphTA
0pp6eSFVG2mkSAvBGqouUbRwu+DyeNxlO6nhy499BHZyE73Kwgf568JLt3+3H0t/GNGUX6xgQpSq
VRoclhwNrTtfhYFkJTDKhdTFzqYTYneMHPrCz5/4qU9Yw+2ZCtM/dh8qiIcYBU/Bggv8sYI5rznU
Oj4dzK8eWnCEBaW7leNTWa2waXMPZ7pRgc+dCsrfZsVN9SamzMAwZ/ysMHvADTMwo6lY+M4xr1pq
fl10v95uu3bFLYbY8le3OH92jxcbPylh2Qss3neVlonP1OJNh/4gCXk6hibkQga7ATTwuD7hr+3P
Z8tt7C5nH4QF8ycqbhQjr9Kh2x1lQMsL++uyKXirRlXrn9aLsFe1JYAPYwDRgEKITabG99r/kA9h
IZ4nAMZcg1/2JJ4w7qL1x9oV5/9HvMKxFd1JwznrQIk/NpgTags2G2XwPdX3tjR9LrllhflVgZq4
1rzD2nInPQLm3b7y3XrPtvsoE35DrVeNe15WhOUjeolp69u8cuBuuumpjAzzxBCOuDvq3CncfNYt
N02rGzxDnsMglCQSrcFu2SfVfYnMdZHk2H9wLZa/d/VxtYYH2vP7sU603HInsMRsESOzg8YDffef
SLQ333NN9LDtpG0K7j3RJLuhBGlb+vcxvqa6dYppPIPVO1HSkW49ggphBTbZuSdjuXRar2rg31x5
v5bdw43xmGPEahv7OPRaDyG91GFHa1ItpU2l0Z19n0B9LsL1RQOZ9tC4VGToZVTEXqfmt3ONPwnW
5NMJvIeTQ6VNcNic2VEaSsx/lhebCfskw20O7Lrgb8+VEl0zAOG1ZioE/y/PahsdeUZ4cFFCsF08
uv1szxOD80gLTbMPcH0rQPTwfQ6S4K1zXlmTNFFIyDnMOh87OH6yExFXOlzFdL3prVqfxekBYH2b
INwyZYMDXCKphW4QMv6AUtoDoEQcRqOsRc5dnTdPUDYlQTOOk2zorm9+lQLYCkfn7v6cwTjIhzMK
b03N68dytI2fODvjAH1ecl1pjMq2zQSHnJ3X09w3y7nrj1IczUCBOgBcs6ePFNn01LYRTk/Sk3Qo
V8BVytzbleObC00l974sL3q0kwJA3B4KsjFrGaIc/OMgjEQ7CDiKWY74ZBJPi3h1ufIN++z+cLSR
q69OsUcS+dDb2vkOvu5K4CKaRwzdmYRfOE54YrnPkUF4E6fAbfbKSm/Jv22Av/k5uebBLWB+YwfM
BvFsrk73RjaehwtY75g/6OzcxVJOazT916dv45LSMV4MZhKo+tXqQilkb7pNgQuoSPg9Bp9j3IX0
zJ9fvofQsJtC8DUCkyl7MFpzeghdse4efH4ICKOB9dKRINtDC/gMWpZNw+JmIK/zEOT41s/o0MYW
I+vT3PKwO77gAkoRjW2k8BLTNqR16HYvLDRLN5oKSmJLSYz/vdqPMsAsbgTanvesF/RSa7pyR90k
4JiPZwrb+zHqf2r/zRJycfSh+yXxFOOPJ3gWwdKN/+6/Ev0V3gZWTUOqaqhGLZtw5KMFiiza17eG
bL6U36UApG1miK/EUM6c1zUW2I4j429avbMRnGGZ9MiCi6HFnN05jw2pf0RH/8w+lvUd5K0C+SdH
fi4Qe59TnQyqQKH8MkquXbyDtGisJgnyqRY4/rOutjmer5855jxQsvH/zJuhXt30uJJgjKQ4mchC
nodm6w3VTn3bcuJ8kDJYJpsz9tNnGlyDNtVMXa6grVhLdbXnmffQOzsZBwg5C95KAeVPYq5Cy70u
QSRvWbbY++3nq8+LPEi+KRf2i1EUD6RtCe19EUrswVONrzSK7u+2ktbBHMNFmvVD9vDu9q1bd/jM
R/22j8+VFjPhaC31uE20zgYB3xUjzL95uCHtvs+vADIzfYWHT0BY/17dOwLgCTomDtLqkoGCSTR3
FE+nAjzL0I7BqrzCONxhON7vG6BjKx2UyX8GjQy8EC1+l2R87vASd8ay3EIHEH4PK9oJpfdJuuV4
1ssAJr6lHDyzwQYH6osBxdHhw+41F+FjMvHYb8Udhb97bCNRT3oOnL+jVWjvvwsdNvX4WpvPLtkV
Kf6HEkHuQXU9gWcJhfYniGh8XGWhmg9tsVfMjPAZgHdH7U+CWZd4dOd41/Ymnl0AKboww5PS5OWM
eZGjTCFbpQZgq3R4SVtkxRjx/KVXSEP0P3op1+GnTgXonb2sDBYkYiEmHtjjSu8tZgeR/uqT5C2R
y0YmG1z0tr4NR8YjLTQdPfbG0wVkVxIbch1k2870il9So5Hvs6DFsqn0bfmmMOXzyLxoeAq2dvZk
bwOC+nefaV9ZNQxkoc4jliMOgtpcG7O4Iwzpb/c3WpjKrvHJwlI8rk7EhYaAnvtYlg/ic5gdHgwQ
qbkMYA8yjzINKhZXXIIMsOTmmGddnfjqmp19DkPtm5IKNiKaeWQOqARNuxTYoDSzG4Nguzq83AyL
nCqIYwIIsc8d6KDHq8BiHGkfGPN+C985cBRxvxeJwdPKoFwwqYuoDRgAwcAoJ/r9Nb/GzAFPeDrq
/ms4ZGOdOxK4MVttccPiNGDYOu+gUbgMnivLO5CASKnEEsmvxE4g4lFy6SywuBC/fGRAlWBzNuBm
HkvdDJAthASPRR584KBmd+4hyoHgJRKtaOeJEXDHGtHFU1UEjZFf/bBna8meb4TFC6BYEz+EUzr8
ffuTyr46xxExh2RWfghKaoD0jkIUq/vlb5fL9Rh6MMPR04q614YqvS63la1GgoAcyy+dERjyTqxZ
bEroBrPp+GNblNcqkde0duknBmAbOVz2TNEJiO+ILZxqbEpWSPXCR1HUo0uk5lkGv9XQPM0L03x+
5Mb7nl+g/NzeyC060nfdCz7SO56tqj/r4bEsLF8aFF+08cXFaBUnjEbsCMb+NuiMZvavFpUzuB3L
i/H30MGI7QJSgMX0fo25M6dEg4dhh/yYwDTB7RkVNmAt+xvemC1qceCzvK/tDJvWMrJstwAYUrid
tzXgFOxOH7bLw4m//pP83U41Y+oCZnLiBf8zrQHmfoYS1e90ItKVe2bVyF9TxrUkw2a/elG3W/9C
D+9IeV899274INfteJWgUR/5t8KvcSqzhENBYlq3epZU5V0T8+SdUbq/KIeFtAXdpHoVUJpRg73K
NxDM5FFcqUMkKCN9qHjnRRm7SkqkwJEXwGN/eae7MM5obnIq4nL3D/Qn4Spb3N9SQ+OdiyXY2k1+
1ncHLDNr4IhFabRRaWuUtZ5MzzPV6N8ro/dxlaWeY75mOtg+xLA9VM2OMONveQkRuLifPWsaCty+
Gu3tjsSsyjo4e2NGun9qJFiQo4hzXYChIMhhcrxj2zXGcUdDx5dT7UZQhZXxQqDE/RqiwKn8KokR
UhXZ/1YShgo9H80eU/Wd4JNRnf1mnTF4rS4OLfoiPcD+HYrAWFHhSlgU7blzyvSm2R1jOjgXw9hR
Vj95Mofnf3rzOrkQdEY12dmNgeWxbFTfNpSXR+EiDEZZCJFHG4LefT+VxzPPX7mRIwpMR53pJtDV
l6+zIK9yuOVmJfiOGJDqZSXn+4hFZf7SflSX5LTMD8be6ux9sR5qYKDroneI/dmnUMZ5IympsRIG
LQWgTrmA7kKBK6IYYbTYvNdjigueKil6hyVR5lnwYbMMIv8V81oXmrx030mNCoVWEOq9dZnOhGEk
D8ZNfwrLSonWWmjwkqe2VihXYPPLiOKJhUH5cd37KKWnAsrlcXhy1l/ffETjpRY9kpnjXe01g5b+
PfJDt1QfzvHFbIiLnZZnRrZelNQ/lLymk8/pclAp7r4zIQSB0CWU13BoGdNWPR7o1ixPQ5BVX/9d
sOi9Y2JGsbVH6zYKCM851bkWU5vu+7pg8zxG/sXtUJoYtuBAiq+kBA9AqmKG35qbRww1uL6otPLJ
Zo+CiL1EyJPahGIxwU1E3VvDvo6D6vV22fW8rnkw0trL4tAKE+HoYI7Nl8/6SxMZfj19lph/FL7m
xsZkFbzyL4tBc4k6ztHJMN4VsgXi9th89H+ilJtEliT1ImZFefRGc5gSp6YorXSYVNNZJw04lCtj
7w/h4znqpBJA5kCGo/cOzVwL0m4XurVGQ7ntx5UxxdnGyqQG5eAQtUmbzMjUkaQwMcqxXpZlOQYq
STHUMClhNQxP+uDz47RHWAo3FEm7ORLbmC5bxDuwkQJuDTYXrunEXJlCzFMJNg2sufi8PacVY1KW
ODMA/5WuLdGKp5071+6KIPVt+8QyP6u4ZKVqykjo8IN4NDE8nbN6J9GzPmXoJ1KhEoxXf0W9YDTH
pRxIPi+SzSwlaTmHgdTJIM2fap9E5FgQ8ofuGJrGWapPZKpEw5lhIGuapl+2zFRq8aVP1orEA7wT
rKWfPdhRQc6fpfMvAejYUKQrWRFKkA1CTDP48cBXrVLmEFzOOgMEIWwjOq/YJhO8h2z5JuRq6dW/
LltSaMVG3oBG9m61ciyBv+14mqZs6Sb9z+6qqsWw7azda64vOctFzq6DRCR1gzpvkwgBseJbv5b6
DCiMYkeKMTvdxFQQFoAlYYx6IVyhLGtpFobe1kPjB4kNlUH++czIOzwEx8Sm31V3sonHKXUlTi7a
x56JQG4oJqGbCfTLTSCpoYSm4lcc52kSunkeGFsqI0IutYxJ9vonzMIAASgFqtyf+mifYRMyi/Gy
sS/J3cM3buqjHshY7fCUQyEKxw3gYbqudeqiZdz0ZamCoxOkVbXXgG8kUXZr6p7NFG4pTYOHWXb6
JUaHL0Jo2b34KbObRf9lNOxfQW47ynvwjh9QwFu0wUo//GVhoJ1+zbmt9TRVZMZ6ozXz8+GOZmhc
rN79n9TowO+HkM4eHNVnPB7nILAnJ+yMX3J5794ZTPjEh/tBzECmH1zMiHKuq6MVMEPpL/6tOqC/
cNG4STh3p+EsVWRQwP2XZYoyE/9iwDv0AJYh5qL5IxgMab1hQ/ohqASgdnueF5TDfSlBXoNal4Ep
VsXNeNE0m/5Gkpu+rzs2w8LqD7Bk422PxWGxbQ1MKwubGaMwQDMacN/g3+USyRjUWvtcsQVV6WIQ
bnaSV3Plm5pcfThn97xOaVnXEBPD4w/oSnZ4Wz+atxnef/1RwN9CPrTmuvIgh8ibeULXB85VdwSS
yBwkwgMbbjSI5ZU0CbWFzPaO1n2eYOdV4WgmpWeAjof7NviXr5Yr43rdVqoE+Td0VLFL0sHIsdBr
diqA1F1JpuL3kLAScubH0v9eHkj9VtTgm8a/PKs5oOqa0gnkh7Tl1Yacj9onBc/KSG5kuJUYVC4L
JKrIDAP4ZjVTb2zXKpAKdEvaKRsebEV8dXZggd4z92AEhHim+Tqx2BkHQsfSaYO64vBoMXDtjvYJ
9YKdFKAB9bWD1AZRYdzKBzC32h2uMLYu9kfImCwIWhbwlS6xywID1vH2cElyF9smvqby7sXDUCTM
5VrwUSyJ9DH5/eRl/2WqQrJSMuTyXzQ41DZZR3BixyT9sERKxdlzP1RZxqzwknFSQ/Fwa+v1geTH
+OlQ/ldJz0VCi/nOhXTd57BlfNQ6UJ39L1upm+Zt7dc7T12RkZx4Q200fQKiKRm9l3SJ/Qvbrt18
Tpk+x8ZpKHNF0U0hLuelbwsD9j1iZOkv5Bouvo95KTBi5yS42n+r2gic6vTvcpsiyBsOVGejOPhV
lpvUNajj7U0xpF63IwYRMuwEUmGpRbDCgERCf7of6AaENf/YwP6CCJM1So0Vh12Bntv4M7RzPME2
psKxsgoUawR6VRQUVjPVee3stVV3+JdAjNq25y0Lpejv4ghNZnoSdIlWfj0E3B26M9CE25XZsalM
wP6snESs5v9k0JrgRswbzqZevHYRLCY8fJ55oYZo0ndOYsJWNdnNl/vB7gnMxEU5gZHXipLIAswQ
WI3ZwBxyjcix4NGCw1GRxjFkXF8GRBX3Jt4J44oWneTnvIrZo9YJ+at/j3/WHamGbGKYEWLhQst6
FoDU3we0x50H0cE7eGFtEYMHk74l5+S+w/jNk6joEuQ9oysaXJiO/UipjciSbwLBe9bz2TbAHCuT
VBjda8gcF0UiOf0pxdpdfxkWGUHLJXpFF32ZT99eyqyxxxSF8DsnRwCxgn31QLkC+syMOAo3okkO
mLPj3uUAzy7d4i2Qj5PArcqSeAvptPEtY8dsITT7kfByU4fUK66B4kgsLNdwvzNctwZ2Te1v2guc
eME32zxUn+gPXu4jKgqWXfYHWp3+9GJwMf1V06SUrLbeqpg2CepUTFgBrwuKF56EE47eSr3DY7qz
/G6KhMtDmh9krW4DYUVjpsBttPGkTt1t16NTlBZIF9Rpqi31fSQqqQw76B53rc7gryjRs6lKKk9g
8CnTKBiIhmYftdXGx5d0jihZutNuX3CKxrIFD+0XxqYVTt+Q7xvBZ7YH9myABfUvDhC+ZXimoHpn
KFYsuBKt6yYLmxRIJJcJsXWfXNQxMuiEmMH/l+YjRJH6UGcovm6NrBYx0I4Smm7SMK8ZJicrOOC6
8taou4yHNkfv1cxaDvU+93rOvwv9ncK3+Rpjrx+COLHvsz3ZE1sAr1/R/MnFpql/iGfOKjMtSYEl
dudWGsdKZHrHpQ+LndfBQNEIDVmAz/AGUHihVhcIS/f1W9Mdeh0EGVI8JCc2cFRrlePMkFMt9atO
38YrRR/Eh507nXHLV8sCa420sOexTpp8raGrb+2/a0CKTOzosreMUHRNo04y4JZNk08zew4DMMQF
priKlJlFiS/pz1KvuP3KC8z2o8xhvPQmBbmjSnw4/8JdAT8gLTDoRMZSKsrjDdHpDVOyezdi4h8d
828yFVcAHfrPSgSyqQLgvN886NPPYuHANVLvz45PfoZ7WYLkGjC/1n9kEZUvcGnNapVYPkwBZ+Jq
/eCJhNFlyTf/21vr/QrJYWBw+OExvIxTKmtrHnaTsc1rOTBamcIrMFpK8LEAIEJZdDse7iozCN83
jKKGobPycWsbTdEyvASyz0dXsXqsgc24C8XrzRuRkhvZM/hRq3hadBvhmj8He35icgiqsolpOTvz
+Rr4b11H+PnJW2tMI1rF1FprFey84OEtnVSJgvFQNK9cd8jm5Gm9+W28uwvICWadlBblegEaP6/N
hIVX7MAkfTDF/1WQCmZWB3P6GXR2xHCYsL8GaaYWLUCwort75Lz92qUgMY5OxLZG0ngOwet5cxuH
baZHL7nNXyNwPbajCavj9OpaasNpffRTFmbIqUK+JsAZ40S8pKDp+nK7NHHUqHr8EnJ1KyL2X4K/
KSfyLSrVPVYIpdPYLUUefgtLi4sxfaXuUY6UL9sfNViqWDQ42OgcnAnTjkZl2F0kmDb8KmnQ62vb
ELeBgjxULcCGX66TVKk3UDppervX6QOqy9tBxKNrjeJ08yAqpUDCulYoQnIDChl0fMzeCTnEZWUK
bDv5otXrfPgzf9M4RqwJFeGL1g1YpF7gSScXb+oe3Pu+iapfnWC9yGwbvTDKN5kmeytpXks1H+bX
BSLbJTLDiutnGj2WbDCprTJD8xqgQ1SFEGVeDGMgSI1guKE5VWjTXFJQqrCU6Svwc/7/So8M6f7Z
uhnWYBQNlNFEkxDu3tIwz3sDHb8w4PXLWJ9oGcko+31ebTmmUSeQ2e6Ji+kGoCR/PyWJ6ngewutr
YDUExO9cgCA3oLiDwFWbgFQ5Q8seyNtdJd6zONtT0PvEj47fod2yJQZO7JhZ1rAD/dEk4xHYG7Nu
0YNyAFCN22sUv3slkxDPDzlIWGzoURz4qUaCKCN4QcdlNgKGch4TvtQ4pWCtPDkj/63/75xIWfZ1
WiA9Z59kOxht3+gXXvgNIILTtfRuqX+L/TzgrwjNZn8UXFr5633X3EGRGgH3eyQDvbNFMJS/q9fS
e/1tHtO7mqdCwSjwoRimU5rT0mY0y/iqt1bM8PUdpaZ1jc93MsLOhR1Q8/ncP1hvBexuEhDORKIc
QYR7RYFtcK2abaA25Iwqa7swnFqKEYUK6cCrfR4AaSppnKEu1r+aedl48W4M7FB2+Aswu/AL0pjQ
amTPgmop3QQw3ixfyo9Q8pWj2e1mJXv//9jNkhNOiwTpH7SVzMhym1avilI6Ca7Xv+Pa86P/lGiw
/V07mEF4/kLN+hbL3kU43Sz7IJBQ4lqPQ5iR3TDD3EH4jijSrt8ntJJXf4y8ttvqtLGT4xHSg5Wd
g2d2FzV/4tetGJ03qaC1O5EsC2CBoBWoSCT66sRYedUKZqPXDsGzLTenYDebPGaI6+yvm36wIuow
AaXSpMTG3ShV+5qdLlTc6OEENm58X6QBdDzERGCMhfMfdo4G+RbieJ/o8F6l/mwAAVl8M6aNBCXV
RjPjRbxaxqxFLJ4LVpKmcZTM8zj26qLX79Br7jd6JJvASPu9GeL/tPGpK0MrGCHSHpHH0KBAJbXQ
OqD4PPTLw61HudKNgPY43rnVFJvujW/b108SUqekLSrTS+BWM2alV6ZaBNitivjWeD7R5NatJkng
//skJL2j48xiQAWwaaKADt12eQrA8/qgCBCVuF5alene8QBIsMb/67AoxTYBbDj/JfKesrJA9rv1
CrX9BGHEplYyr5YL6wH40i9WUvL3lBffIrMZDW27JfxCj8eYyZa2q+sMHVzgXQf7Y9f4c/B4QR8t
FSDNezmz09KTVjNudwN+DDqC8DuDV1110B3JuMKJqo3/h5E9MmngzFxEmQg1d0OCUFKcvrB932ma
mBUQxA5tvOgWV7DZ5VIla/czktr+PZwdTUC08p+FLT77BNSTp1RenEa9kcC6h3yVRNM7ZqIrP8WV
luRvIoddJ+wLsrx/50vl5THvl2V2rT9GR9B/JPyfWCfvXLBFTSxz9GMnqK/O+aA413SxksbTVCaO
gVWZj4dAxiUMETeRkDuAqvoVhg7NeEzdoy2UEv5jNINo2bq5cXRw4nxLlqZCBx3jZv3Br+wRPJqi
dSqLz+5idaK0M+c8otHI3OWy0lxG5sIA5ilfbgH5czFsuTec5eRd8ZO0HWwC4Ma9L0xufgOpYQb/
rD7rXAhzeaz5vgXx/0KC6msVwLYaIsb/t0oylBJ0+JnqqSGhGsEcyzjZEUyPOZU8SjXfv6L0f5+c
MSRFiCqVLIuD/oPb47/cO9RvasLyT7lA1Nn9NbdfEelXSDIhZTdGDp3F2k+gMoT2Au8vaz5Q/nqK
2wurMy95J/jMwwGuRRZBRSFSsbdrh7BpUlJCil67YrxnFnGH/3B+rpXCj8ZzvWcH58/uSEtsVHVQ
5qDQNh1jfw3vyxQj1qGAc68Bputw8YzN54Dufne/ZrxTsaew8z6DzDma3SPI5H7RofZ48FxEndym
d8zNm0VI5G1aCDyYBURt/hiIeQeK9WL8zJ9eVXy8liOAjVX6wfijVKznq5sbUXIeqkGndQ+eIT6C
1tYkEgFfVtOnOEUyTA+hfnje/iOkJlnuK3v4LQmPdoYmNlPCiliKE/Aw9cLhv1QTkh1EVDEeexNe
cE7MN67kGAd5yKGmKyOPxTF3SrtDw1fRzeozawtt5s9P0AQLpNICoO07Snq10yZJlsSJcpUJL6lj
QZzXGSN4ppn4s92f8+qvaC69UVY8dE7monHbytynniNhneKRm3GHOaFEAWMtHTltoNUyzA4IwTuF
upAoVqg3qsX3f9nCXoZNCpa4qUUCValQfMLITTbDgrq7SibuRM2bMoKjiiqBmjznxq5u1AcC1+mc
W6TVO8mGFHdsrvXPFwu6x16RLsZUAPsqDQNSYQSUJ7wZDunWlxbyW2ledqYnOTgBq/duk5yonspZ
w495FEIKdbkHCrhFFf7jWqVWkfs1mMVkLq11rra+J4IK+3yOJZVNyvhVQI+3BaNCiK+wQldZp92N
W1fh+eKCnvbpJFE1gyFGF+6Wzs4fwYIRvkeSQRFwfj7tgPqLrHop3S86bSxbYe5C+BWjwq2lQIK6
pYipi0cay29m89h1mpi2dE8AYtDH/ZCpZaVmclSeqI3aCkaBAaA/NyJo2283SJ/hjY5A1RGrsSoz
3iKu8+CPb++1905A7DE/i+gWyX/MqSsHhHuL4Z5f7VRHXGQ/q0MnC806zjah7/QF/BMucF30DKAx
/OtcA74BjL3O6HBFGn6eLY/LHpGMXomVzTmKewmvdQJNY+fRm6z2qjL97Foh6XgBCV6CNF2yHJG+
XEH6T2eWtrhxbYdSOOs4s/qiQy4vSYYbPar5jE7J2muekJraYTGsCCSz81N/ChJFHOfQpTBtN7Nu
6O2cD6STjh5Y5sV0gwQ5uPj9PS9vFPfUR1UOdCtnaS/bI5hPqSAb61hCwT969aSlevAajtJEH0MM
momKbSlGKtdY4aWykL5KPAXeoPM6YJdkiHeahgTsASg8XMR4iQEcYkhFNwnz1yxzW0fyh7UytoZD
58dpve5Sxe1jKneycSK6zA7dlKot66EbMqKk18noB2apHv1V+VJLDtZCatuHlmA1dOFk3LqevVrd
JcIHhx6zyTxGUSSLHEUnhgQGDJM83/ia+DUy+12Zlb1zH+QhJff8RYRFvcW/Q6pttRJfGtrHeiKL
et1kyshjw8CiDbrxFV6HSilaGiOCJ67/yfYxycTsbPgv2tGojQAfw+QL/kMiRHJTSkulZcSvdyeU
fHvqWTaq+0mtKIQ1lxG4CewlpBqBufVC9euH4NFHSWTRDhUVpPwyIPednDZFt4Wm97IQdjY13Mnj
cMXrcYbZuwY2qBR2JZEtoB1pJWgifa9jy6Ax7zqxsQgTMhdDpzACwiLRecRK/WkLphWI6bio5eBP
lS+oE/qY7Jpwk9PLrmYPtaIKYPT6V1uI59QaY6gMOlKn1eHwtkihReDOqod5TLsPLOGGgpK22S7w
mp9DhHwxOSc5tTkwQZXr9vcNqb32SzERIL8ia9/zqgLvxkOdpk5LxOM3V8jewllqe4nsDMbp3ow7
LZp535W01xcpnNc/HfiHw41Y0ztZJyrigHt78BdCCjJPwDrpK2APj7RiKTOA7hwRvDaXr+h93u1i
tMcad8i0hIYyaK4qzbMNWRy02esHL4q3s7L+xdGdciox5Q9iisYtsRKVGOS6O/5r+lWGnXl+tnNE
CcgMdOi6Jrfoexov05L5NVXokkambGe5qg8rU9qtQHu3fm6EL1BNjofI103M44xyw+ICOrP5Jbdz
P5NF/yNDvhY4tHZykyGC+Dsr7jbQi1iPCp9iMIYKt27xt45JjGcJYbybPpSsG5rYTGa0MraL0Ifb
M4/QhJ2YW4Fpd/82BRW4xLM5/I8BusO61MGNSHYmML7S/Mg2QcR/9f/PIY7HHK99fCXOvrRp5xhP
vNRn4gDtYWnjlI2xFrKe6ALzIkJW3punvC9AeHzgdMRc6MjrI2XNawOgesRlErSCvKTs6fxirNoW
k23oRqmh4CzDrgHP7APkujhI8Nom1ncbXBOp6A8xab1z15fJAvwfM9Nve61eAyJWb4KtzlSFP5sJ
QLfZ2OHTVizGntIXAWXQi4VIJYzChgGDxvXSjraabW+nRiPRe+Xo0dHFqHhbSSnPgHg4M2y6ekZz
S/o+D0w8JU2d8UTAlDE9aaiWUedxwFGHPZMp3brDammw4STkADYi8X7sYKUX0lULE2se0DY5ogJX
lGm3IsahmM0sW/54ZPVrp2awYHzhQkNWy3kjTSdm5ub1P2FedrnhFdwny/DQUUN1/8yVIc5GLp1N
IEesIqDPCzYT6GBz3acck2GEeZ/2ze0Lw5HorRy4L8bEtj1wUlysGBFYZNB3KvxF1xDWmTQQ1PX/
xuync/TzBSEYp3cppb2R6yzKq9Eclii5l4yg34eCnGRLU4vaTSq1HCUisoIxWWuXPGAhu1bJwtav
DDkbHir6AXmH1FU0mlt3hwUCi04FgCOIFbgE7GXDF0IRrvvpgEuoilC6TzI/Zz/usSAQchgmXSK/
TbVgVOloXgE0ojtfM+21KRG4Pc2MhQgK4VItqRt1QAJ3iWkr438LDpBmj8UzDWWEpVOWJXCfPAH0
funj1S8Bn4Lq9pF8/ZPwNRCW0svHhsDXeAxw9UWkQDyl594FpE5IEqLpEI7yUMgWnZUOATWR9jzg
oNzNJuFLgq3sJp49bkNDAiK27YWAwDGniPegsJppJrfDae6RAZ7E4jJxaDBmoQWvYAMalRQyPSqj
w0poWVBYNAD8Rm1QF2aSXV8frA8fL1XpbyUqGtYwHgQewtbmzxtyiYzc/30jFaMkRjUTOGdqW8wK
KLunt1fqRVisY0ArBV6RjDwhsTCmHJMa0mNTgadeMolt87VCVjaYNUaQQP0zxXvtUR2CXQYzI7pO
5vbua1VOam1e63V1qIJGhcIX22Ditp7yqtWqjzb5af6DTCKy5WofgYxRgVUqBhIDF58yiISPExm2
jed02YzxNhNHHymheUne966hF1j71+4+e4ozB8z6cSKAcU3LG6pkcimKFQBWWA36LckJN8ZyaYvL
M1eK9hhpTaE2K65TvSUaLr8QcyH2mkch2zjv4T7iDBCKy8xGT4wpEeln/b+ptbsdBFZbCv2Cz3bh
2uPu3hfiJ+A25oLjXR7XNwTz+SyFg56qq5c2vt+2MaJQzER+Tzwn0Kii89XHEFfMQSlQlbejjWQ7
6rhHnaJDBCtu1VoZ/FGUF14kryzsJI/JnJlVHZ5ERbmqHJwIWM61drC+pPEDpRzvvmYX22/tb5/1
kpsAdZSC72jdIKB2khjoTon26SviAGuVXuRZbSi6GFPvuYWrM1pcavNbu0OSfsMBgJRyCHbTYIp7
cXsEth0e9bGkaYIewWuVXSskQ8rxN0uAHAfFmCxEmvpmJ8JETrv8Vnz/hMiB6nwOTparnjRurO9G
M2i2Tk1R4X7tsu05yphqxLEQDJl1YeSg6ToFw64pnJOfoOYe6LOhf60jzVSqROU3J1WQsloBbQfu
qrcwwezQnmBUmRBlGTGQdEdXCC23EQ0RBA/L9u/YjBZ2jxtGZdm86daSSA+3N4p54+E3JwVYDZtA
h2dCh/EufZYXxJpbNrUi2YqMIyRFop1XIWU8KdwGk2qqy+q77lkvAmZNTi7XqX6D3onFCpV2sLtX
GgKx05dH8KMR74hAo35169d+wN681b+VdV57pFjQ/7E67uYjuI0GTUh34HkNNhriBE8iig024c4Q
mMKfgvfFneqQ2BGCJ40FQKL9LYaPzkyHHP8FGsFdQwressO+KR77ZbWP486+u1xLaQ1btin6OcTL
FvYNkxHg5ZAxG/nZDs34Wb6b8UbbNoi7DKmGRoc2xLVKe4VZYghxPpIKN/LMxetXjRhInY5C80fV
I2kISp6KKWTI/8MjHCrcMmsDWZqNV5mkXhjWslyWiWgf0vmD2BfrjpwMgV6XcJdT8r8NAncosxLz
omDe8asx0rqk//Z7iOFnXOLu9ZWM5I6Od+CfpwnbI9zzDp/6rFSVZHFiRnDUaSIFySly4TX/d+lj
2nLDYDvK3PzMjOnmKrlDsAvXNf0SqWFo6O0fho/mIKwwN6WqKS9lrjbj/TImsz5Dqcz4gI66DdP/
plHzuRxa+vjaapBW5FslGim5AZAAiyFdef+V9GEVM2Nwk1VjqGa1i8Vy2F/e70Rd2JkJ51hmMLt5
NE/eSk7Zg1Z/CjKwL7FKRueblL7pmZ4TabcVsMt799rEN2OzfsnLIQQ1mZ20SIe23D5Bu7B4LTYB
fdYiM+B4nvg83TJJdj7hK20hzWYjpAA+laRewSPkFk3xSLPoryGejCaKXehCLud16Rvbzg35PX22
5FAobL+7VK2v67A3D99Vu9S6OxPIRZNaZ0bEqIEpJsZciVtWafQ93Ns013r3RDbnmGU2dl85nSXT
7bcyg6y44Yr562nBIaZGi1fHfaoqwXCnhjR2rfljGt47gMMH6bStgUNVQOIY7jGuhsWosLfMA3dr
KkASkWnyRSRCVpXaJ3MCmwp7lN5E6GV5lJeHErCJsl18gS+BVMb1LQB7vaIK5XfOmSVd2csoupz6
m31Vnlchjt1oTTa2mzyaPopc9eBWwl/ToLjpha+vJUGnb/75pKYkJyJSk77Hn0nPkfFZrYeRLlJ3
Kcqv0JvFbHGX257G2rOn/zAGRrMIdlCBrptR5I4JwHz1lGcv2qNpw6tCPc7Egt61y1ocpt9pL7Y0
0km3u9RGhtOu16SDZX/fxzjgmybcTKiseVYoiyjUNGN3HfES1+cysm9mRjuyCgE3PCrcA+TnuPXd
EyICHvGh92BAeqw6I7nZ6+gBOiwcNtDK9j5OVtfMFTYYVg118frMDJatjeeC3mw1eCyPGz7CPmZN
51zCKg7bok+HWFA4+TzFD23hlsxN8TjVbekn6fdDHlVOr/Dh9F0Uj4kp/N73lUHKoedY7W9gr8zw
fH4Bc8kvuBp6Rxg1BsE5rLRE910ONqXqVo2wPFT44a1B0qtjbto8PW5goro/UhVXSJmKn+8twih2
RnvgFQGcOJx+vgE/gzxmhCRSues324dh0ai7Za+T6ezbtiVMYiikN5Qh7Vv7hR82xhI9YiQN9E78
0QtUVS9esrItYKvsAjy+LRnwKMWAOvSVKyJaIgICYUyhAzXWzW8Yw+8YPAp23ILozLelHiK8zrDQ
H6ykXVKHB9iAlRgq4anh/luzfG5X9qu50AQVPmm5dzALgRQUTKZGbV4hcAyJomGUMglMpM9YpdzO
KfHP1qApTmxrwXh4wnFitpPhC35dm7KtQcgfyqvNcYr0erZbEl7xgU3MZ6hvJvp1y6l8oZpGmoVV
tQ5xaNhD3/9zRgJgrqpWwz1msMoWl0jCx9PeKvhqPH5Q03lrxqCq4/NNQhYsQf7bzBtC9E0z6yTa
/bzVwfmiygENXgH2mMVUpx3yx5Qeha5hAoWf9qIigfMiWA1hUhWASQn/+c+d3LAmh4pKBCzaaOxN
yY19MS+tJiKvuPz2qmVjLTWtumJU6E+jr42u38Do43GFxqWoJ9hR1r59ON1x54ofq710yVoMn3Eu
f8YzjBj/rjfE4n0XwTYbTDOq1IRPA05cI1mqsqkzScdI/QVcWOrPv8YDYlHtBusbbsPgOa4e+q2A
esnSGXatTu5/HiSXy4SlwngR6sHmGd8GbMp7WvMuwPXW6f35ZRfvKaiSlCB/LC69gOnVEO2+052V
IBEgnO3ty+KU0Tyrv+ZxP9w2JEbW7/+WEeqlKn7wdkuhVYIzbMaucLEbfJdKRKLS3jjHmzqFmjVn
hkAof/VIDVYRG9JyWyMxMUweo07E9Z+6sxUSUSCc9aPN4rvSIu+xNADKe28LH2jykmht+TU9P8AD
g9RJb2jziSm1NonL+oNR5mjCNNVzdWNHrnzsgJYuZIwT4OMJ0seIdDFZvokS0ir2FBy2CNk8ECCl
gxpgSxEvk/I5qC387ckhEMX4IWCsuBRKpHeIx137GFHQ3nq9OIPJDhxtegD9LFUtPaKJepE2Ch/J
H/NUN464K4lFwhPhfRBLBUjZT6V7+HlHddQcWuwGtsnfqgVj3wnT7v5aQDdwYxSevas/SHN02med
sZ02RQzeFjeQSbkLQ+C578yV+FznmcftKae6/m/PxjdHmpCh8XGvCLaYMUHhV4HRnjnf+FgwJSPl
MSTLH9gOmDjEBwYD/Cz0JkbAExLOdkU3vsKwE2VKUbskO9Hbt4hHmf9wiNWoa5FW6fAN8dMYwBYA
tJdjEcOThyrLae48MjxVKIVbmmczEef580ld5VJgeZx/7lluVsZ3nXJztH6kVawHwlteO8/FI0iE
XJW655iX9piVDa68g6dvQL8imdH3T7yNooFbZ3cYlfK3WeP61c1FU9VM6/IBfmA0yw4b9l0eskm4
0LZk4ut3lWysNh5zEMTl3IICHKe6KlW9iL1v6aRVQmKo8mKYG5KbztxQL6TgcEUHEUy8n6i+MDQ+
7f/DMdvGi1A8B7kgdnsWUuqAGDnumLrK/LOy9Fld5EebcWY5baXCy/Q46tNNGw8yFWeo5N3o7bSf
qtWkBqzGGOnu9M4vrZNSNMVvR7ZNWp+1ttPE/7vBEJqD4M5MMgwbbG23DvW8SKf89wLXbvWQkiTo
wpe/dhA+R94/n/AWxDWhrGTlIqIX2KhPmOyEovsvgb8peplJzqPBiuDCClBPeIgBtXcOmOglCzzW
GmwuLg9yiOmte/1MGz1Jv6FZ4nnGQ8yEofx5u0D7azaSNq93OIu00/yxL8JHXMaJ8F4dgwHop+oC
zPTXrwlryV4C0vhANrmnP7QGQh+5xJVcxYjaE5XtKN4Kmb7z/Aeb2vNEVRTxwpGxsTIuZ1UmwSTL
6+LevvZJP2TwqpVRTRNquoKj915ZnTgtj1Rr2BhSbd3hbJ2yBxkz0bPDh5txsn9VFwGGNC9uuGcC
Eu6QUNVOQYto8VqooYdHrtpRWfbrEcNOAX1QlnmW+EXzT383eQMF5mFQcvdeUBhyLXJpQ17Aqf7e
1HLTiRLWpkkzmI1ob3w8Lq147Lse8r16gkKeQt0+JMpYeRiQGIFJ6z/WocZxTUjL/CJBb+/6MFTQ
V+Pqv3lbGzpig+bo3vV5RnSvGksmSsGQy5zK/JfhfXGxRuv8ZVYFPRYJf4qU44++LwGvdPIlL9q0
Mnz/lb0sjaj+zHj19KLxmYf3YCq7o0duzRUorm7nmj3eKd1qD/Xna/KEvb5Gb450Wx63U9uEpACZ
knF91AmtlvTslMNbqNnRlCNYD9LdMiotIYbfKDNhG6Lh/QX953j+5ziAe6wAx8vZzwS5MTHuae4o
fTRzoyEtdTtLpK8Ftc9BY1D17pKTdYMU7/IeV/l88qPRvgwhp7ZZ5JcILeqaRCCFdXPIc7Sf81DU
zFrHtwp/Mp78gfvahOxPFkhl04z60m8xbX177qMSYiVfWje6inXKAHfz337rUh6ezyr+wSspAN6N
k1/XYmDqlu96m+AldYfyKBvoqTQw0a/6TTn2zHDk6vcxcfwnsuEbRFtwIXbJ0hAmICRYdiJ7KNQV
//XtOpp5qkOJ/H+suLkYmyWhSerityGz/9cJpqSGN9pk3e3rJmeWjcKPFu5XCbUEGNN/dd0gwFoS
t0fX9XvNZrsuDIZtTpy0VfzG+lwsGqaKFkkO2DwL7FCxor138IQY9B3gXsgsA9qCyzLpDJr1uMs6
lViY935wuBf9bJF/aMWnpoXPzJkx7SDIa7k+R7LnG0IFEa/pI2zhwkaldL6fOoXhXoyEo871OdTr
m9Sll634IfoNy7JQb/4ZJFTg1bEgweVAdTED1jPEO/WGlT9xEWy0pT9t1d7g+tnl/kYACcURrFyX
Qjaqeb7lk369cCf+L0eFkw0kj0TAx3MpbUwHm4XFvOB8UU90afd9mqfcdCudUo5R1fFcel7KlXaZ
UkMjoQ9f0v/4HP1IxCt5d/4jmmAMXwWbsHyMeKEaVwkd1ZjfZ4F5Fnk+5Nd5qmTwD/14C3AB70jP
fqSZReyn+QJC7zPO+SyW4IvPhmNZmJZBL5IKJObnnijM0uw+cyk3n54W4HpPYw0r7ulZp2W94U0C
Ki8F/Sds6x2/Pw1g0W26e/xNcX6TIdTVDkLezVVDD9krlxl/yqvi3YQW9MoFNUsKIt+j8Wa4EKQQ
Gi+PuwYNZVctKOzR/JYPEGbnxmUJh21LW5G2WUDfFFh2TXucKRJzDIm18Br5fhDtHqaqg6C3zVEU
LJqd3tlVCt8EoXHRUfA3C2w/I+VuGMNd3z/FF81oKPQaE9fHlpzXZ79VrCTda2IEtPHxkkD82MIu
Iv7NlhUObUlBS1+6pxEH1GQIdJGWOTPWnFuPGyzP8k++KkP4tDW8OCutcG9Eq4/4NIT66Kuo5Dfy
uBnPl+lblqtrdsPCNbKPEobfvbcCQhOO/NrHHwigiLJxHvtb3z73UBWtaYc+6OVwlLJwg3zaRUB2
7loJrHfgb8qGgFwCS+dOnPMS8wVNqfG21M8r9e50jOnFbGzSA5kOwgpC76NBjDjbTcCegKXmVLtS
X1NW4Or4GY5TPEaFhzleJ6Y/jIeBK10lsY/cqn/gp7YHZIr52QPImAmYsDJfXS705cuEUa9xTRgf
HBL1GIqt9BkUgdw+ddFuc7h1KcAnzGp4cVyPF0V/vS9oG51h11d81gjEDlfg4dmbP9+i7g1wIVHb
ZxkxhoATaQL1u1/gHgbNix7DOOLqhTcJOnD2S25PJuLXaVWmUg/Xi8OtRqWhN4M4B1KgvIUuk79g
LyVKMasy26o8De6AcMCm0XkUSEK79vXucXvrGCUC4b1eMLpyczzIG9dnOVuNR/ZZV4fPyL0p15vP
zKDYqmoNZ0k7krTEfEQo4dvzg1OBfCA3MZDnUk4kEwLgJhL+hS7xvQKfvLYef9O9S6V6YdBzRKnd
FCmTxmCffe3PxTRJamH0sue0QKbLYhyrKaV7kyJsp1mWpvgs6L+UAfAZGV2Tz2V9LghhwAw0RgkU
wtcUm1RIHNftL3YXFGWfKJl3H8k78GKPbXAw9olXYx7XntR+5ukgERPuZWjIm9pkb/f+EMwjvr4z
3eW8edotNsi+KeZatNMT2CRrfJ0DLL0MqeSM750nRznE3CWc9mpLgNprzEFCnuWtCr+l88uKiOKg
yo3XynF1eJSaiklxT8bhCVuwAg7NhrV3EWk3xtSr3wX/1viGy7EuPH18iQ/2OfZQ+I702qmiRgtn
eQcfTxfBnJsKSx3GAYEU1j4csv+10I0aXH6i+xxNwtn2VRMo1YazkG+S3l3cIt0yjJKUrUIkUaBB
EwgLZhY4tQdbPYxyDs5RlVd3lXtnNS4fN++jfvwYH9aJOkccp/8Ogmu/oO1p4WYqlSskEHVJUvkh
DghnOsmMRBQs9Fu6698Zx3geWd2K9rFP3FbZgL16N3hRtyjD4j8i1VH5OGLsjxgRQV/HhwUV/bto
ome908WMfLfWznTALuvRW8RO0e+yNsSCVFIepRmuiTvYiEQR3Euc5ALC4+LkycntVwaNofq6oPOA
B5T7w11/oHVN2zvWvmWJS2zgO+JUlNIsJ2J8sPRjwml38tCduhbtPOw8/FMuDGQadJO3USFXjwaU
wYzIH3iZnT8KUklb5jHOFRBlB6YPLGNg4lh+HaE1T8klkOUIRKpiPJaMeoq4wObTBrJCPYeUwCk2
ief4NK6uteye0VFBHHi/y60KJU4+iyHE+cJqdjzZfTdqJuHbA9o5D7wBdEtLo6jVuAuQ2G00uOe5
L9iBdqWxtBZKF/tkDYnFX6DmNTnz2QpMhQDc1qfyqPuHnSottLjAVKWZyA7YM3FieCEc5GN2NV/u
rjOsFh61YBGtSeDqQH7PqxDjT06AZYf0CA9MpI9ZnYryl5GK/NvkppXrWorgvq+F7921C/Yfj+at
H/GQZfucxUFom7n+EufIUaNiRHh3wEeN1zF7A2frtVcS+93Zc1/wiE13zuQc+tRo+xetRG1VOy7/
NOqpWHBjoMmWtOBTpAr6WPUuQG60/ZGg5s47Ct4yHXlicIiNlub1Ab+BNqWD7hBa9Upcd3xRjtNV
oRZPq25zI/5ANtN6qwE1BnELhiMJLU2Etv60aNP6+VLKdk5F8QHSLZigRz7G0eySocFvcmbU3KXU
Z2v7BKHuZWf0sfYKPzosecleypJWxTKbe9OMSO3x86Cbh600y2xy7wsQ++22jH72xt3QWMVW+IZ6
NPJPKmzETrbqNyfCmJCvg/DpMMqCKS5XzG9UZ8L10tezfDJyLh4JmBPjo/068bCipPJpJsAcBijl
05PxsKV5rkDlDsn4wRbhAZVoFmQ3x2DsW6C40IShy9cVt9xnZ3XqXwPTA1UY9Zpy+IBar7DT9Yzg
m8zM6yNYKJyooWr6VjG9CKDgjhUoMb5wLkXXdiUibRqbYqqW5VSoBYN0BolfwmQ8ljRMJu+0tACX
F4tvmP4XNCS200MnXaKwwfHKVajaRetK1uMKBYWBOs7kitipAQxvUP9j+pTifed0NWZ3AmEUMstY
X9McnVhShEgrk4+sQgXXntqs4/PGx4jX2dYY/bC7kwxPXGgIvPgRUqJmwOo1/SjDTqWt9sazJ34k
VzEgG7O9k0Wjz95boZvL+ySosVlCr0yNA1LENLqC5ajpN/JU4FADFbhMqc6katqJYJoqLBlwsiYU
H1sscE807hvQ42d81l9PVAIM1B+p1Y15ITXkNVVR14Mt5P6DCT3wkyqLIxFzc+lqkDU83EJq3gUT
p0EeAH10CLOfONmAkAG3BjojWN+mM98IKYXh1t3iCoYtUbPnFdB4oMl2mnYAAZj5Md7E6SNtEBG7
6aibKrKYW07H7wbBhZH72z5xz/60Hz4hjEdfTqRpcF0i2cNXE9+iDDHXZ9m6Ks5nd1M4YpyRVhPS
8x6e6ZZ+ATs06fNoaJT0jPhY3cZWgt87Jgdvuw+p8L2+c7sx3ecfI60VgRemgs6OksUgSa7UNcS8
l8mlvkh1LXHaIhGoEui1ye8Zw3Kq+hob4QTAO8JXOlUlt+PrUxAmgEntwTuwSSMfCqIGMMC44zhV
h321VYzcj6QTQmjfnOiaMyY73Jr7kCZKX9Dhwdhh4oeDZRA9GStSPKaFsTokcekIW098x0cwAHX2
ElF1UnL7nfG2HF1iLZmCkasNWpPSuvRoyudOOTw2DQLo9qwOMrFM8H+ByRFHnd48DdbvdbkT2RRd
rNKO8PY0H01x3pt2IIqQcQVWxAFz+3iwzkoUCg6ZrdBmazMAS6KKoGis5JK2qE6svXTTxDMu1sFY
oTLHNjIXbgPnfTnRU8TqsHQrHN42LO42tZMbNvsoUcHk9tZgqeW2/7pqNdP8Zi4B508fdV2gjNgH
OM+sIB9JKIfjYn7JZN1RL0MbBRb3XIUhxOR+BSAbkypJPSd/OErvT+nQygGxPfM1fSjBtucbRO/i
6PhCqqAGqleNJgznaOvBdEhn9319JIxjn1c7Eue0ZRA91XoBoKacAoIXhQGRGF/AuAB2PeucDplE
udJsb6wHwBUhT+REzUsugdxo80uDXgvIuImdEd+jjvgXXKe3qfbHgY2Ey3kKTpJc/iwh0TCZWqjy
O29OHcunMNyhg34sZ6+Rx2O3iQ7rmmfieIgtjIm5VDp8mlCireT8XD4PzTXNnA8BgrM/x5SM1QpG
lBA75zK+SVmQsjOy4hPHSIn5A3QS0I5WO4dBXawFm3Ela8mz+xgjGfwodQQ+zw+rIAKbBGeUcXsw
joAqNwSEs13Sei14UQypWMOWICQxlTOKknvNw3W4JqV8ajzcbIzvTWtjTEzFMroQTxIjDwvJfc9l
EPka8NZzOQfh7xoMzEgfhwPYGPzsz/MnlAuXKscNpKBdmrW4omXhhZXZaM3NPCRcTfJTCJ1flSF5
rU5/Kgm/vbuPAZokIut/MCvAxT+3CSRXZmPZSmX6jaraM+Iz1Cg89cCcSNEfZoh/YC67GfPW04Br
u/NU60TZm+qnmTv/tMXYAa/QZpi0JrIC50yHszm2uBf16xhtBLCztnyGwZve5Vs19tyNUayx5YyU
hNGlsfyZwCCEEs0MkakJGnV2U6zy83nPhdb8xc3Bnc68Z1Qr2qIqxlANNCmbs5kgXUI3CK6ximyR
2Fm0XWw1Xih0AjEaQ2H9oScTCHmJx1SR7HcZ4G1f/nOkFfIV5FpE3aWzdl2PV1a0agfWjkmld5fq
O4q2FtROzXHuir7fCXS+HASGE3QK5JugTclaC+mYpS+J5ZEtsPe3Yh5ZNg8y1J+zOZQN8mmOQFwE
azNY+eNZ92X8i1GM3GskHY0/sOTDZAs2ybTn+9CezUQzoop7pWRL2vHjtsZ8JbpPsB71pi4gSqpc
TDsqrrNG+ihjSBDKf8E153WKitrJctY8SoxX+AXxXaVEDjKxET3Kxruo1FhOmMulhmM7/Ejb7hDj
yMJvcoGKDjBduTHpT7FbenmPGzZLPGNcb/EJTYuMqBOLqWfKIq/2JyWGUqkVmhZCbCT+FaIjVc5c
mRgdSE6XnNwY3phbBPiybuOEAWxhcbYKnBwRD4k7ZDk4gzlQ+zHRYFOYmylAFLesoYA78zA4JUtN
Q4hfQjMpa8wQIRzfD2SI8ajVNd7acdDSGexQRkOsobt2SZE0cHiiR9yfY6S+hOcdnO9BLlprogai
9y+c5AhcUeLCFsdDLJ2yH7/ZvLK29DTgSJGJhSjnsXKc61KKqI9mltsh0T7dEXNNmDdCggwTe10g
lOhI3+ezm4qKKDI7ADb5zZKEkqDvcuY/XPlui146IMK+hL9BxMKEX6T2lNX5Z1CCGQMvOq6oJGsF
RHoSVbWknR2bOtkRNOYnjhsynLvdCtL862HQcozgCFGvXbAUSMrMd3YaKiMqif7FaQiO1X1uAvmc
yAQ//aoCoq+gYGemBh/jE7vCP1MdXTxMTIQIrykwPDLfRPkbdMiAWpMhcAR9X6qL1QOADoqn+cV9
34VtRdaDxEXvD60z7+jL+PBQmu5j4YsMSMO4EOWR2rqmJrnayXl+SoXvpe81+3FQ5hok87PzSU7i
DMf18lqVher21lKFChvux4cBt0yN6IItMcxuUHNAlZ3qUyLDwrv+54e2lTz0K6ySFmxAdsXsoJQN
avGZD+uVt9xIaxqot0OpoCjjTqa8RRmCRKGx3657g3vjHndw0hRDKdhMMRGgfORzOuNL6l8hssAy
diXBxbzbUEiJZW/l980aFY31MHzS609Ao41gXe46A4OKRpkhsGa66cwNz3acj5JU0OXelfr9Ao4H
TdnasEzD5lohE36pSoU2RiAf15OfafuCi6uGW1o+VS/2AfcdpSlGgjCCwPorfem+u7B018YZ3QFC
B6u8ivawssQnJDOSfZUIVdhGxbTc/Iv+0qu6Quj2FMTDHzmRrsM2lPJjATHfGoylfX4B9C3JpmA6
Hmt4JZCYVA8ByaUyoYIwlkhi1XEs2pzdoRrTL4klwCa87CDmVzvjdUYr0JbPuJHulDuQBedp+qwM
5ExS8I56M8JZsDWc1Zoi7czKcld0RdkBeO6JVYSTS1G6xgiG4+ITCK8ptzxuaSOVcgz/BnUgOVjU
tIzOAqEtoHtWmo5FMrusXhdN/O47tFmTtJFdWa2754EeT2ZoxM0p4KvN285Ixgz4E0I1tHn2hDIa
wckoP4ub/SjCprld7LkSreU0e3SDkv+Vz8n12pC9Adk4YEWIz9JSGXCJmPd58s1nX8ufHh2Fo332
GAH5aCRV8XNMWFtjnk+6BG4qBZ545QlRYnG1PWcJv4xcHeG27yM8xMKajBke85jf3TiN1inO+HY2
CZg8XI+PapLz5nLrpE8UIKD6VKV+WbImoppOJd2k66KQlMXUMYi5o+66anbkXzyrFkm65lznqGJH
98I6HIOlHWoWsHNGB8+UfHTFzJRtYRXkVdstXoo3ulk72h2h5mao8jnSWQIw7DtGm0Bxq9gtRlIC
sQ4whMfj4hfCPw02yWUrm2hRFpaYKVXG6pbo4HLqdyBBUwwBq1l37xbQEo/DYSXDblacVfiQfvcg
0BqjT2q5pZsNV+OFPm77ts6mammhboVvuZipDshfu+jo92A9gG3FosgHZlLr/2FsGgbyhCEWbm7d
HWG7zd1bpMZ2gKWUgx2nExT5BHil1ifSJ/UfkXIBdRaIE2YjX8UO1/ijYlNsYCBA5dczpMFeNpHQ
Rex2Q7E/fkd0LT+U5QhC7xn0cww2pWc7YB2XpbPRUh4Lpu3kmzOR+uEsxzb8M+62sVpy/MbBiwTq
V64KFYqs2xjSeZB3BgLUR4s1sZqAsrExpCJjPB8HMJsjF/IyCqCvSKLb9dTMOu3UXVjoZQUDUg0F
W/10eFVJcZYV5eFl6jc8xektdc9oIrRzWmiu1KsTFWLrLPpZ5ixpm6ZeQ02PjUPk589SlncUsJQK
U3I0hpPKJ2hxD7V5lQpMm9BCj/1L84SiIsgSJPJIw/SShy+K1lSSZLSujVZCcLNDJmyAkJwO6iMe
EB4qE57yH5ICD7oii0Q9oCS4HVQ3MueWU3FrB5v5uYzJeJD+I4duGqCVcgx2icbeebZWMB4Yf48D
yEvfsAfPs5qiA5C0gOIUuL+SnoeRJWsezUSHZfSJ2VjxPj9144Peda+dHDIWqDehZNNtaJoTqsE+
6ZqtqZA/1u1nORGgS/LbPDlFqACR4X8Y3kKe2XffnQv2D2GaRgOjUb6hIOW460cgqykg+JbUPKfz
5wLiR/3OVhMYfLmz/VjGnDaGWAEqiHyIqmvC5pNB71XhzdhzcX6JgnY90M3e7F1ozq+w/gB+HieO
qjbKsRvuuX2JNl47ACDaU5tUwF5DOYUWYC0EKcn6ijMkQqvkdz3vcsXJZ9uPMTpNlzKAVnVysneF
BkkAnV7xhgSnA9xyPdsr4AmH2hwvsSFwUGn+7Hl0h19OIUPdwHuB3juyPFKgxn5dBx2ZhApxCDrH
QiA55EN9gIUB7BHaFKcyB5NmPdzciftX1fd+KXVz78gTFH7VF9RXLnaEAIndpOqLfDcUyHYhptvK
uzSnJX7NZ3RaAurfAu/0tRIopqmQNlmAIfP3tIfzPs2BgIbNydbJfgNdZIEGkH6kBGY0SJ0xnRCh
UPjbXt5wwedQ4BHqAGnIG8ZgqfhMOLEqfxg9pTHpwKFdle9DqMeS8rDv/9hPvpIDEa52KfrE/uPb
CD2bDcjgUI7vYkffr8KHHMB3e8AaFhr/u78wmQYFR1dtTdEIB7a5tY4JoRThpbDuSRo2RkwHW/V/
Zg9jLwzxegX5IZP2m3M5W6ddgG9FLrig9oFGI614SQZEJf8G1w+PJTFA5FCo6+a0nUSMjXsWU+Do
6hr5UdMREDAWF2CNla5SJjzV+j5xtzG3Ht8pV4jt3XNTbdCnNzgEtc22Y6sVvzvuxNq02W+D8aly
ymyKqaN9rWGLW+0bmg8t5PdKhiR9lII2I1UmxAb0zlSoCGknlGxnCam5qy7lkaatAcQ7TX8/jBD4
TQ8c3dEi964hzKeiMFgIMOWltZ4ivlVMmt1bFH2bk3Qnyhqb10dusoCtppAi5ig66VErggyzGkBD
hpEdYhWDsot56/uD8j+HHWeAZhUyeHV7S5f59S+/47s6RWmEn/WSnZAHk7g2LVeJO1sjsCdLjsd+
rE0jfPYveN3JF7kq0OF7TYa1Ews/Q8oBDWX+j5/UjOjeIuwsNFXfbzNf2WDiI3yhsQpsggE7P8kU
nGRsjJRmYdRGfWfblc5fTASbvW+8jF6AKS+WuWQUfIDVg1x7N5w1xdHXUKtm3UGW/GY00vRmAXOR
PPZU8AgHzdIY9AAUkRgMEs7ekUI+oOF92n39c2MY718Boqb9wDl9PtnBZnhExpQyk2l3Hd/u15ly
qZHptWBrzy6PXr+9M1KNDXXGua5IsjstfPwclKN/Jt/0ApVfKBTCpzkoVHniuzAsPQ3wnov8OC1w
9D75gR6pHqyYVJOr5hxvdA9e0dhb8NO1UuUH2QP4aQ4IWgnOEMNPhNlQdkLaNDj57c+9wVQG7YA1
0fR3uevtByZAIPoBubeKUbVNDC+GO7GGNbrjS//xhIFB2sO9LktenXTIoXQtF3YTxmIFneeO+Sc/
ucznjrqGSHf8K44nXs+aN3Xf7snVViLI+cxc4v8d74JAPJlHPN0aVopNliTkRtPIkYVJlc4uZkvA
LxciXKlw3kMl6BxfwFMnVQBujzXA2R4em1RDR3jmmDsuQDRt59jIJBxtFv62rEYOk0TWlHgEeCxI
DLT6GarjIQTuVCQe9xJYdVlkObBSx6EEUn5NVuZheHhlZ9/Qo+gP17MxrNPKS6kSAcKvyja4AJ6l
SqCrrAqn9FKX5oK5DfDu7EJSjp3f7wGSqxvem9CpCtkKkG9twhEE+fZgdI1Jm8saXaII2X0uNULf
kMOniKWRGqN08eGDUYI882VeOJyFLMksGokVm+v8D5MdcKan/pDOqy1HB/zsdsBuLnrxhv/mRb3v
niBfsSy3tznC1COzIj2JqHNaqu0UGmLwLXMp17e3em5ZQUWJLOB6J7DJoPK/OTEMSy/SuRL2OczF
xXspa/5y3XxpaIXjX4J7vBVDZgXwyxbdIklMgB87RDf9Ua/AyVMT3DQfa16y69cYAgvI5eb9KYFv
VwRLY8LZ2ExoBsCKYy0IKfTGy+hfhNjquksY15CjWVEdiQWEEkqkcKZQIrIIYaU56xtOl3d1GFPm
v/EHnn3U+b18fUWTLFx/acV1gE3NLbJC6KM14VIiZXLlKAprESnTI6buNP9MI9N1dl5LeJ4zsD70
ydNm/oubnKIoyDu4egwRp8x6QQlXvLfgmll3kYADLqoWRD4MQOGc8JNjVPY7rGFjM1J3dkyYgYIs
uKzf1WddCRI60xLv9J5PtMpP/+4rPCP6x/pCWTrz9VjNPM7C9Hxlb7pf4epSVzavkTIl+sKgo7J/
gh8HT/WV8ol1FbkxnCz6X3MBaQkuqzorNKDqjYGkojTThaQP1K9X/idLDRLPptX2Yxu3v5fyshc1
O/nkGp8dvThRZpYZ+giFtE9TLNsenAb+E/4kzQK5B9shJiPB7QxQbSOhH063cOl99/2s7B5XTspa
qNeZhnJ6nkLelote/T6S0bw/gWkBjPWgrwbDLUnzborzTBVQ6c0SCeU205zD508pHZQqz4+FQkrG
3NJGloLSWWzHl7pUfbES2bNxnJH1j1+G1QVda3+bM5KMz4/8B0OFKmG1zZFjc/g5pKErZjR+882d
1S2iAhFGrtLLkBKEnp9ARTedbGqxWHaxHh7xRen7rNTwjm4jEOM6CnfdYvQXuOrU6NNbUrGPfBgI
FM4MysKu+a/Iz1+VHKJM7M0AiTrCnz8HrxDNEChaTdzMcpwvxXDsa7Zhwth+kBD7K95BEDI2E26s
R75AMGEJORJemq0FmKmgvMPX0poknl49u/TpbJiO1ZLI5z27kxa1/ELS14ys7sqbPxAzFavJ3PMp
kI+3kqVExYo/9cF7/MhXHPbF4Mdkt1mkbUOhHArDK1tAjpOd2XlDKqOUGmdUA1em+SAwK4xe/d7a
W9j3jiMpRyk0gN1WjeeyPu298DKwTJ6yBu+gIWIlZTHNh5HEQXws23aEE+M/cQ3cvldFdbih+c8v
B7XQQx2RxdRn1rm7LYs+ggfCKH0WGlyPpdCORIANuZgMgnoASd+1ovJ/w7wUwEJtLfD2QxcvmQgF
rb7R6jkUq93zNLksWAdYp5rwn4v4njRpJw7ut+4iE3P6YaOPN45f/ADDLgLCi1qmcOmtbbm2hEMj
mQzn/u/3IfR8Fk9ZDQTKwqUHAxvCEIA0N6cVHgZecyHXOYKhvoUSUWNs0nvZsm7KZxhKdtRnhXdO
pXSLe8Z0v+J0808rgk9sS4bNytvkxM9qQx3dfz8f0hL/IhrMonAo3DfhXsyBu3O1ZtTvRKembGcC
08WkpPdWGMOrTdQ/q2p6pAwXu70pibSr8TmSgxQqKii6PYwZ4mZyFkVykHWZ9LMnzyoQsGEckXr8
0Atr56ffNUe8nVC0X6Z80OYA7aQWyEZ1fCMSNeT/uPZoi4fmQrmXpZrN+RETHZl2XUCU3ZT+MeE1
amDYE4x49nW2LbOv7p6jJ6YO2t6ysJABmQ/iuqd2pEIcwlhUb5yd9mX6R/nBbYoLJC4bG7y6Z4DD
53yGneD9aCIIAO7Ij6SnVnRVqDxGpXADPJkY/+AOxcSMFAEkHvY30Giwvb+z4xr/90TZYgR3xhuG
NSMFR0T1rEaNs8zZBsSQ2+3t8j+lkwcanrWG/TK0iHy+teSYR2AykS/t2SLnIhTDalyq9hp8ZpAD
5SHdHKZMct7g41ErG+g7luCoOqmb65ir8baXRbwIaECAdgEoUjgUstJmxrcsyX4m1VyWsoEcf+nK
N7s3c9oiFDx/s4OswGCaDm8nHNCjpQWOApRSEq/fuuJY3xRUVHfljnPpeUv88dVwhd5/vfs/ZHXw
k9g2eRv8lCnVTctCfIyMv7712hCm5jYqEWO+KLnRn/I0e7tXZL6nYWoPE+4F3bQ7J47PcvdARVxP
PL5SZiG0AZ5GFl6mOAoaPlM8LCDvp/EMdtmJQG9XtTjzEvp+sbJ7zxFE9y2UWC/8bD+2fPlGIAFl
GIrUf4sylYLKP/y4HxpeE2VhmfSXT467IxX7CvEwbZRNJlb4uMuden63WqAZJb+93gGCEXPDaUZl
8lcii4lmJKBBMagtlUK19CpzGBwHU33/ma0EqnzH9Behsld2RQFKSUoGdb46Hqu8LostkI1GHhdz
UTvCTWHq8RunIphfOw3Kd1B/ERY4ET4v7/UfLdsxjTToChuKwyF6Jk9LzCy+GEw7Y/9jiWvsYwL1
HRwig69y1Y+O9cJ8Y8neTqvEvrgiWNyDjgWVUpMTwN2xHa1FXXCfXQSZ+TYVVUU8IyDM418FpCTu
xnt9SMQIVC4iLoaNf3dmyvWNU5h6WUbquoKtNfvZNwASTAJm7ZfXYG0j3TV1nZWF38RJ8IyKaw9O
P+5PUFWUZaxIncLHumFdeNYNOQe2fWwYeU9bCpxqiDMJkTR0VL1rUr0kojU/J5szCGg3s5pKWaJm
aOdXQdTizFk4tMLovVQLB05z17kEtzrryI9pC+rPiFq3uLbjs6Guiz3MzCk1L3edazUlopxMQttL
3tAz8rwARc5zJrBj1Ra8oTDn/X+eRPygQuMV1m8thQav0Ac+OzW/XZ8CKb1b77wlWJNbg8rNbz2w
TGNbx82CZrWQotuv4xOPzS20oYjvxK9f5Ch6tJndNibRK5CiZzHdIp0sWdaqTtOE9wZd1hjRUKGx
n4rLBjEP+DUU0R1PjipqcSZVP8qL/3BvtoifyED3rV/wW96JaMJ9Eb9dUw7vVvquzGJElt4KhH03
sIDa6UH+CuDwJoIDte+93Z5csjq4LGiYPjy0vbGWNs4wsiGXl6CXflYR9wPZ3qbnuJcwZqze/OOD
9X9NOPzxdhzdQUGIJiI0upluSi0SXdZaz4v95KqSXmeWN87A+ce6GycumEPLbyHPalQ8TdKM5dM5
RzRNbADnHg66eu5m7oMeUxBBGcXp09XWj0sB29o+6jmAA7WIRKE7sJLyVFu2De05qP+Fq3aRPGR3
v20br8hNXI96YMGcQ37PC6L4C0VRDl+VOrvFBb3BKP+XEKF9I+Rll5IcgsJbgEMhs7ihGr36m60K
1jz/37LK6mBTwobWsyFCz0TEOhjAyYTttzO+fndIq+t5dpMSEt3yo6oxhNXbGlps/y/FGayliRdF
Darx8lN2BQUAUzfLw270SkITbbmQL8vfvYJyyAdOAZCw1cOShKjDsVH8HtY3owvez0sGObVYx845
uc0fKzEe+8FyXhbArXQf49W4+FXnwDR+wCFXaCihty4Oabhcij8YcGHbSQqIEiLt7k5vRN0efToX
08KU2BDEDJc5jcgQvQz+bbtvD+GKhyeMhHSENZbHL8X7C5ufiqdiiAUh/eIRBVd5FPZOyRBI5uY1
1r+cBTpsIuwuf9A5yz0aandYstGn+y55enPa72j1s63Tz9PmF8Bmrtl9JN900FB1xV7UXgLEQiqu
GNPB5OYf4CiXzECCcgqOB5eE74kxPDF8OBNzYGlpZ5JUkNQz3br2NpUgErc31KMcMH8NYQqyOh3w
XYOIM14Mvzqej2H0Zhgvg+gkW/aqSJuQIBbLop1tvQLdaXZnzMadsJK9c91rgtCnJB/7k2s0xq+X
W92aOU1Uj0TvOZBVi3c2bXtNfJtSZMOqsbEbKUVf4FdzsSh+19oJuKt55jz+k8hCEM3MirvofnSj
Uia+TjARi69ZeVHlKsWAfKmNhAXjm2Z8JsTl7jjyKAebMEwyAcFMepWR6PHHra7pc0mspWX9A3un
IPykpu4+WcpgC6AyCVgqXKAKVZreKX0PtuICztRT9TZAmBdTdlcpelOHEWBsEleMDRqLjA6Z8ga+
YHfCRBA5vVdzLLhQ6CiYhkRhNJvygtzqsI2TmKw2EQlb+bE/siqD8ayJdwvWbaerJqOKwCv/7KD7
z5OiMorkVW4hmG2HIfRCEWUndBPdC5LXtb75k+r6Qv2Llazpz3y+Gz6bMqIgZTm5OA4xotF4hkKq
iK/2J5VcjFnMDRAGnGeT7Q8wrVXJQNrWCSHO2aUuoP4BNlFLuBLHIVypyZQxD+P/MmIXVAGrakdj
CtzxL/81LAvM2ulEPVjIzrmiakP/yEy0zerelhQ3BVYTajf6r9qpCUnH+rbCnM0p4kCmDNgOsv3N
uM4BhEjuZAaonG63KcK+kBJ3nekNiNw8L7virdOhYEvs8bbClTV+qredXvJ5Gf59Pd0BsvvQPrWd
vq1akmFjSV8jqaN6hw3j21J2j7Kn6jC4Yxp6shLbLaImccOR8H95jyMwMk7NlT/9IMhYyRuSZzKY
/pqGzTQnk+CpIbqkdksI8hwkhlRhsXwCeSU4s6b/dZZkhmux3847SpGiFgMzckQ95UPDWY2Hgtw3
lyWxWE2JSXqw/RU1M/foGdg83C5yKUe/SGpJShfZfO9vE4dBmagTUmvwx/CSkrhL87hkc63kCCC5
11eIxLdjF8bnAtZO2ixUzWLcFJG0nV4LUNfKF7SSE/oG2iM4ETlgN+zBxBO9fDek/vWMmI+IH8af
wNsjxH0wRWa6iWLdknb8qCGmW6sRopFenUXSEe+G0YctUzHcOT+Hm4oFheyF4wwKUOzLQPlsc6p6
yyavM+UuzhIJwvMswFSJf4rrb9qazqrVWNFKOdohDCxFkUXQZ5wdMLEFYNN94V8RlcXiI6WGPBBN
hnt2KSVeIVNCjKmuqjhXyxtcWqJi2/YfniOWEbuowaoEVgSSE8hawEBxeRcVxr5qd3hLzHaFwEJu
n6RSyzho70296qoNxat8Dai+FscdeWai+WkinQVBlqCFpIJIIH/6e5nQah5+dASA4nYhv8nR52VW
OGBhv3O9QgUP342xH1QBFQna0TNJsNQ91kvbIJ0pdvclAnUjqm2E472MXT0+L5NDDj3OGuTNE6W+
T5baR8GZa9CfJCMBfOKdxW/5htMvUo7RWDh8cUncxbc6j16PEpjXdd0QFG81Ci56CQKUDAoKEVu8
RIXBXIxhOKZNkbMkN4i81WMVhBdRVzE6ZX7tjrGZHmz8Glb6BN//mnZ8q56WdyYi39luAiUwySNL
egtiGv0PQffZhPf3reE/yOIUCIna5zJmrRsp0wwWplSC7sL1z+4R36Hc8Nf8UybDnUr04gUK8Nco
ErCjvR5vmZlfFDXwRT7w1ZMf1/XpaZ274UWeZdwHVhE5SImDxx6Z2sPC3yqgL1t26928DUlGuyjS
cMUjLCeV97JyqL/zvYYk6aQTSqxN5ZdLzcQAgJ0DJ2zm39T0B/wZ2rfXVnaYTWDi7uv0SJqYdA5H
XudMGw8NPXKcCXR7LG1tsBBuos5T4+NoxkYcQOM7dabDZxBANFiWqr64tHJeHZMhP34ecmrDHaq7
PSwOpz1PHc2DIhv2AQDYjvkkAFS4qo7VQFrRsHnGWgqOuEVikHWakJBK3uet2QNrLePb9pAGO0J4
Z9jh+2nlDAQrRn1xr+rwuJN/K61IjfIf/6ZI+fkKphjLU8yllQffYA7aXFo/7+3GCrGsJgz7S3G5
MRdxlWoGCFNxAvl2vJ89qP2WzP51ueqmMohQ/RZW93xBkwjnGzySTNO9le7Y6X8jlN/I0PJjFW2e
RiGruJvTKmMa6Kr3Y8pwzuC5UgLfQZy1K+5gOKb1ilT3i3Yg5kNuvD3bNLo/wB5EgqVpoyKurryS
HXwKW4zdZ5cgwUMoqhf7sKYm464H6hXTkMvH1atsGi7hMWOmUQuNRPj42AjMqALTpqP2rA6ZG4an
BsSbBCk8/lOrGTRIDzKLrnB6Ze8sSCfNAJT3uKJYAV3kOdKpzMsJO54+Z6nOGxiwDqY/9KPgocJI
Hfr4ULiYANZ4p5Yf7mfZMoruXqjnrf6Hd0v7FqHbQSfq+oH2I8pyxDJzLM9mC1QrqBWSM24LM3gk
VqcM4IpTbrl7OVf03GdgQECjwKsvzc2Iy7K9OWICkQlMUpmT8aTDpVvLNRheCQFI4q5oor71+jlS
MRDmH1khmWb33K7t4N54S/BT5lCsa+P5cVq7ruDVhgEiYI6OcF3Tpkrw+Z5filp/uzm0pNMIgHBd
L72cuMH7P3DU9rQYZVyAv5vA35w05SyK9iE/t9eJ86cWP2ULMlANXka/Izoe7x/xGqv3Jpmu9uXj
MvAJdKyGevvTd/12uPRKnXnFWcWGqjwTRUsgLKnavyXDkMr3zMrc8zNLwVanvNXDIdlo9XdKWAz1
wLnZ58EVYkaSaJMUjZo9zybZ4OJFcZDg2W5Mqm9mBlVDG/VkC32+frS72nyqm9pBK6XRSAX0UF/P
pNVap1SKQDatsXUHGBgOJeJbkmHz10F6iK1cutjbUO6+YMOamzcq0TD2L7u8prigMdjyv666Prn8
6ErKw/MZT8OxXGyE07DRvMzd6aCCpAYgQlWnxRbwOi8B5cDlJL/XxZROPK88V/FDZDU/KVXitOfc
UOzUr+uSE2VZCUf6mpxPDN3d1xiAA61TQMBkftPwvHU3s15oo9nXvkTuzHCSAqhYxDvToOXliTqx
ViBTfzfslkHUlDbN9Y/3qhUcDS0Yo/xtve9uPgSAwxZcAJBcj/wbj+dYfDoXLcfDRdfq1MqnCobg
rvEJi5RbYNUOucZ3JBocvB311y90NkggbZ49W92bEDkTs/1uKo9EjH4sHMkc0mjaC5jVg/z4cIF6
ZObhtvlKbeFtRIlCxtHADygKqL4ZLWIr2H/zSLlm9IH/p2EUBMtuspJjvF41dTwmc6P+Kwmyq6Nr
35w6MGT4tBoIIyiHYWn9g2OKbGN3rnm5inhrNi8BnYJZiQjIazjGQVzO9uBqOR2bt04g/FbUixrm
yeRRB67UXfazPLFHtuzhnARXStRPQY/sleMci/Anh27udbr7v7AU5TWQtgt9ehEszc9Ohbmy58Ss
FTb4Q/x5118HiuFE7KteLlzqwNJ/Hd+yTzXy8z4okMlSx7IJOSFbUVJ/zxTR2ak27ngWxpItoFX8
YOdfvwW1fcetI/MrsBPtZ76iKpZbUPUiJqDg5fHO45BcEFm0ka+PvG1Bu66eyUv1LN0y2WWnM+Oh
D3OFoESNcBbbsPQMY8TXgznqNhsH4fdUx41CM5eFOD1WPWcjaXBLXV3PisGcCwTwum9FgOYZZuBV
lPdQMcUwdWBd5Sm6YTg9+ZZSdJ+DXefNr4g5AGxIKkpv8cqSwULkcGnFLe6tAoDLrkcj05AWC18o
qiyFL0IHSdDhh7hSLdlQoYJlAuMjiaa6ySkCLaDVdOKl0WWKn+D7ElbGGMTYJvZG1fnGXYIzcEVl
Fev64vzg1wT7ODJ/BqsdEtEi7zmZu3XO25sR3lBDZx0+plP2TUFYeMDPDwANiMeKAsNEGOWdk0qn
tlf8LchniX6FLPwl468ZARLbkDyjjcDrVnGoex7UHrgoI+X2vh4g5rI0DUtZgUZR4NLLAZRYWsD4
NkzlQko1G718Ta7OJIsSFkhiNsGmJ8l7Wi0WJ0QG5w+0yvE8mNyRD76DuX6d0cJVQZ/DFt0hYbvR
+rkF5OwyRyVH8In8MXUbX9M7MPNIdHXSewdAUKxfyTi78IcaoK6Sx2mltdiDyGCvoumnacV3wwSQ
qOFVutBz8HwRHRrbwf606VTX1itkrr+Xbyhw97T4RqvbAp7MRQmlOHtU6QphQl5YgKhf6BN+wGwA
f6+fVctTiiPTCN+MHE2C0DG07ewzMI5iW5u1Oxb8GOV6qIgAZNlAnV39I3ayDlv5hwCNBlsRMg/W
rvQfIhobobh+IVVJMiHFCfqXxAVDBWAX+/yDbtXRtYFzw7X4X9sss8/uyj9Zpyiz2Y5B3UCNGK+R
R52Uv1yEixc4UYZTQMbFfz9VIZBzIHX3uBXiyZeORfgJlN5nDAwFzCiBSpeyZfcbzuHZcA8VHMg1
Ak7kOGY88ROO1/lkb546p2TzS4Vf+gxBefhic+8i4xaS8P4X7tvVs4dH9H4/jE1K09/vgwr/LklV
+0RZJe9uOjE47+yBnY17oOGf53xxWF56AIF90//U2PcGXMYICOolhvb6115GSn+0MR218ii/5aci
HWXAYv++02ratyqy7wJkvIyjcIL9BNYLAR4J0TA3jygTQQFb4hrbzjflfALxJfUiLgyt6EX+TCwP
UaicogJB+M/KQp2a8pUWC37IrtnCRcnHL2FoHABuWB/aiPQfqbtuFl0LwN5yx/kxEgp6rVx+fgnz
tYs0rXMhzvwGUVbc3lWo/qUpzUNXONDxjxzrQq2frCT4lvrERcDX5nEk8pam9Ht9cGvv0OKodnLE
1rYyF3NOurcVJnr5VV4X4eXy4LALv20iao7Ew7aFRWcNBfYFaQYdEFdU4VwL19OhiIx3xNiWT/6J
Lc+5VYn+jeNd9oAvauLUj3xG5ik0SdmWDPBJbS0bqkBhE4TZkKKMbkDXXT4IVQrRqT3GixKOTfOt
IPJIk/RjDoXpgIqDdQZQGcXbuACZaJZoIi/F7vAhy3/qvjoJ9+pTorsPShNucetgS1aMtQZshN1n
P6jjNMuCaMHZDmgyx92wTPtnAKuBlCzIAFTdiSpmBySKIlnfS5MGtCXiq1T7sOLUna/nd5EPl/nJ
WDUwLraITeMbU5HkquQN+gKa0HSnVlIg3MgSQIO9i7Epx02s3GsgyiQS0ZUotPJ5sVoxCZiaYVNh
qZoZSRf5OzdqMDREjH65at2bE5veuVS29akKXbfcW6W8NGQQNeWBHis2cp9f82vLhCZmAm9z1LU9
yYEsZtkm8iVjHxydZgo+0cHEhl8Z5SutWyQf77IQ23S/nmGY/mnzHYmMmxKWk013bXJj7fsliVQk
nbMtDiu92cml7nsltDt6N8CIdvvET9t+ISijPwKLuANh7uDFFcUckLslUOTWW/fWsI80Us0GrC2o
1K8Ta6UwS4UWChhgCy6L1Yc8g8/OqpYvtn7Q5/Ptl7Z7jxWA8k+lmUNxXIgbd9vvC222A2dWIvvC
VN/fHNutIbhTdE/OtVjPTpAOURQ0+aoq+nhoLMqHD6KtlYTOycnKpiXHESu25LKs+HSB4JzcAvZ/
HWoWdPjlQioHt9JacsusDRPcaiuc+GA56RxnejPX3v/a+YD/i7XvFDYkBO76F+S42dr6miu5e/Pz
Kc6ip0Ry2XWiEIdSsRNMQ+aDtvrZStvoiMRzA7ybgJi/jcTuJIwe22rlCCwuqBMVYXhuS2NLsirS
9sC6H96z+J3cKcmOys1D4YgwbR7J2odKzn0w2n8jVoHEwTJl5Y733PY1m0Uh6SLtdi/Jmxlj5KHL
MJxj+HxqATfwE6ZC2BqILWCBkVhojuJQzsCY6ZhHviU43Qa18k0N57suxlmgQ07iO4MqfFOvFN8T
NpF2l/yXfiuTIEbQj9VcQpTc/F597jpr2+GXAZ0I1C0RyWHkAp0HlsknKAclkFScD2wqtoAyX6eh
jJI02v4v/wYr4kxyFWpYy3XmyH39F2KDjAlDux0178Vj9VfSvvw6+aHJ8Qmy3H+EUPUkKIFDqplN
b4udlO9kl2LUfnoxFL1DVxM2i/V/+xEf9uraeBP5V3KfkdPwgyTBxXCGWFbj+2lios6Z0LKneSVx
IpEFvfVRGkaatWUY3AH1d4en54UqaaTveXSAcmWxKOZrQIlY63VOhoKEraFjkPWi4Z8F6hQa/JPg
3Q7txwWtBlVFxlCZvlbiUCqf4YsEuZXW/a7pFe3Fp9lNwsBYfwKnh2267a2yhYs1/QhmiNLb8zoD
GbvQ5MAVtKPvsmJMq+H3SxD/SYx+Pr2ZU1TdJpE5zESCtizdvu2+cBn19aD8I2153E6gfm/WWBbW
sh2TEeM0inAJ3QxJyd21XaY0F7DltdEGZ6U3K73zGdd2KImtp42mOUFsqOHoOEBAdSd+NSNuezNK
SIkoNmB5PV+3vtDZ6AZJ6rx14boKahEs5domTDBENcGelkMor65jQarq7TkHNloeL68bHvJNewLX
cUwXuc6KKE34gN4sH2m9gjwGsfNI2TMZBM3uGoamRnOC2NFEx8VE0GSe9AQTFrYdbV5hr2rGI8h/
iSJjfhAy7ZnefNDb+5ZBvlYGQCCJaOZmn+ZgTwNlbOmxoiRRv2ReG4MmIx99/Bo1Q8K8SfCZtQRn
rUvF3bH2TgctekSYwZchJu7mri3lSWtPluKtGVexdtBJQKO7Tl3cE3lFQJFRa2pS+mD4qhYNaIGr
ye2krNn2qXsbw2n0rN3+d8Kohw5qmRn3xgqm4XDRS37HIOYAGuW0fst+x9ISYr4EzHQc5ZYjblHa
3Ud6auamSVtSC8Vj4203xmS5MSeGDEKzRJyU0tkdjc4qXslEQRbcgQ3YDa6PRlPyxrYBYlHIiu3F
VJg++YlvM8aSoa/UzDLLw3esJFlk+HEuFM0WFNvRtwSDDfYvNnA9TSUU4IOeOOLhEN9+bFd8p3bq
/C2NW0Zqxtb2GEiJDvU6D+Lw1VI6yVA+xDzMO0j/zswFkQ67/TJYPz2RBZcdodJ+kQCK1C1WwvTX
LZ1AAo3rpZF51r2BhtcjEE27W2Acw9X3j48KbE+DU7fXVRCYQp6EefFTvl0y1wjsaztydT2584aR
3kyebPY11WmcO/fi/ooqguLAdFULi+oevZ42lmIGvoYCd/KzxotOdDSVT+PbqCkxPwoeZRF9Lg7o
NF0N8qpTfkfvlbxA8Xh4pybRL6E//McvGo/hVDdiuEA4/NMEKsnUg+5DBAj4UmvLyZyXEwnbDo13
xWJHSs4C2Ufz/jspQAUshPi6bvjEoW3kgc5DW6NeeOlF69WrpuP7ZSPF7IYp310kP8wnpF0zUPR7
MxgWrUM6sofTpoDmTr+JzxZ50lz2NuBtBfR5b0PNPRXofGwyiOY3X33i6JfzcIyACocukMh5Zt5S
MZHYNHr0wAjWDYYriOwtHMDQwlZ6W9IVMRHdGVPjiMSLYLYSj44h8+2SPHZYcA1ychct8hvV213q
wYNRr2tKn517wMH6lcAqeVBpbSYfxyWHq5LU56p0qWcu/RAHACPMw6WuzGf4AJlCloXNc0mdSjgo
ZTx1W4xhA1pBRHApZ0+42PNRypG1mhPwP9cX1ZRsDahnRp+2AQl7LlbJOu0ILWqvRoUETZQ70n5p
I7vcKUppvjsiOekqeYsyKiurDlzync4d6QQm1rUdII6MmDtUilBWwKrsrLFG8e/dkK0GusiTuvMJ
DE2L6fw6TtNjZGM0+ZDIL1pTSwQ4tA5i5I6v4sw25zAemypx9gg39e4hHoE54K/2BWnTZU24z4nW
KeF2zQvkG2CRr2m/CdOME7rmPVWwqOSdxAbHlhqc3n79Arv4wExz2u7AZRx1tXn3aMGCU6o2Ieaj
L0TYxCL3MmjOMf8883wo+SMRes/w711IdfjkRNJCJ1lhoNJW3fAI17cpCtaB+n+rY/V8Zixa1z00
fGnCwRsg+RRFEuafHf9H+RGoXFunzjJpWZ61+9IhFu528eMx/Mr9WNQraks7jSo4zKHR8a1uuzBc
GrU7qWa1+t5VHsRM+eEyprJhtYkiv9FQKdS+PndroAGMgIzhaVKq1KD5ZkX1eN64YM5cvQ67Jt8O
2Z+TxEZqIQDahXue6rsAzUqxd06N8gIs1/9ZQ6qsuf+GC//8IGRApz6txhSQx6kasLQZuVFQaFx5
uqalq2t6+NBth8VtGnaQlktFfkI1N6L6S8YO8SEqaczx9AxpFklbCzxKzVowLEDPt6yMPAlrz/DU
lsx8xSX0UFbDF3Wat9uzlWPNlO+gBFq4kaBU+mByyRKtqf5FlUAyHAGBrK0ePERhtjS7dfacGn6S
L04Tf9UV9kxE+9yAnavz6Jz7dta94HoS35LPlR0N8uxR0zcdNt5XEHQs0rG83LtRa6xA8beG3DQo
qceZm3JTyDDNbrHGR9XY4Ws9b68hbvvMJHLRKgMTu7CFbnVqljo2pteDXTxhNnIYayiKYLABA44l
Bk6cEYzdighBCQlsAY441eDMGk1lfIlq19Q1oQjnK7Qw372MAI71F39I6AWNBFKibCD93RGObxfI
MQfimNsUNW33OUPDjIkgSkyHwgublXoe/IJXHG/Aq+HiQIOJwzbJZXEeYBXUQWs2tFP78QpGWTd3
cxr3TI25SE7YGd1uu+nlMfI63NsYqYGS9YkZkGe2Rr+cptl0iW+q+1dzAcoZJkp0mFa3gwERniA8
pqKFUvut2hMA4CUKzLHIm8hm9L0QM936IZY2Z2cOnK9P+uu9Vno1ZVYb2Y6kjszkkAi2A53tFwb4
SoXqfhdz3gA/bnHkVsqDRD1xK8WotE9FjLeV4QA6kQBdg0eiMG8XsTYDsGr88WR++8kImYI2K7Fh
Sw0GiIzgF7KWRZdugX2zAa70VxQjwsFggADYGKrku3kTLp+K19okX+0P0plV8z7CL3zWuA6zuk5y
2lFWdR4qMgv0UNGcCDwVyHVz+wEdwGOViMJSZ10DAXvbz3HFst4SHpqBtVS8FOijRdFJeuO13Ao2
uLraMlPLQqO+aFANXrvsZpl/wOeIQ8l+5hW6neSC7/qQp+FUGoOxfU/V/noGrsQBMqCednnAxpns
YyG44eh7Iyb0LTzORXoAtKYYnJH9kKRVho7LyM/Ps57sPWAnuUqTFcD9xYCM0XyMPNLfT0prhmv7
dWe2G9gYz14VxcHwJK6E0rT+mxmZknJntRh2YS4DAjC2D0/UUMSmwk4j50BVLj+gM+NyUg0LHYAD
SQk/J/Zf2tqOUBIvmuJ0zid/hFnPapogTT3+nQ6YwdHxpZ7i0RHuXcle2qx426rtBwvwwEegr0R2
Fm3RGyr2+PwVkyJuHAfvgZA/dqV0FAaY0nSVBm3NPFybCZ+x3upK0JsEVhxIK8b/SCZAT6c+h+w3
k/oeuUhpWsnNoIIRjNCMKvGGOMcDlXTFZIaC3iN9pWhcmJITZ29PTOtuNDmCIMFMwJu5zT62AtXo
yE9OBt6NeuByi4AuCGh29ZZo38Jg7SQV/v/ZTBAnC//jvKgcXWKTa0Kmjby/VHN+DJWrhlNkFGI4
CI3Mxu8VX0z5YuaKMZbwb0BRqTZD+lIBu8K9Q0eJRprzR2UR+IeZIyraDtoUYxjAoNzhwela6Exf
7QoirFNxUh0olP20CA7febKa7rgvDxcfdAzd01kg7+ZdddK5jE53/13iKAlxT2l2GoH8s5ZimZ2J
b8cKMnowoP1+2PDjF+Hd2uCcPsePiE+DoCDQ0IH4+sf4d4EChpbpnoqS6q/BBdGBGXArdTm03LkG
PbVRwFkX/DHqXYx9uCQuXAkKNyrpKiy5We7vt6MwIqk8ErsJxbx0lyX/aUlfpAK0AssyXa3KkKob
hy44RixIDlk696AKtT34jyLQcU1DvRI8xvkHTnPiBCwxYVWCjnkW27WfL3GEHzMwnKlT77jzvou/
sB7d8x68DNiR/CViOHmEW5b5IWbk4K9W7KvznROHFfdfWmCeDRsT3Jdy+0uF7lw4eF7ozI4K7QJl
aaawpM7FbJDOsD7sEzDL9UOn92H6mZF2ayNM/q1eY5KdQSzd2JjFumY/dXuomo3A3WRIf3a5R8hM
Fl4RpA51GL0qaRTPunnW0/uSN15TX6cZS7McFowQaxvuu5PvlQHf4EgOw1j6eQO7xvD3djIXldlu
SN4bbSQBOHCNVsSmFIHGrmg0es6fJC4h509MydTuI0XMIjc+rm/eUl40nIh//eqRQ37HXvsmplic
M4qKCj7K1UWsSF6uwcOKHFHPR5pRDLv6oNoc53wwuzTv7yyVyoyUrFKur+DKTMJWgtk5R4M8LhFf
dC3skW2FARcGJrrqWpN0GCs2RiJ5HW8A2EAHzxn2Xs8la5jb/fdq2f8khfHMHJ5n4QDbYzITHtiI
OuGFhHJz1kfqGMwAjeQRzYiPX4YyhRc5g0BN9LsKPwfSyBM+JhEQh3FbH6/GabXrfxVuaYvXPhcp
I/s89ZuprpiQtqnnUkOIxqnHWwL7rT7/jpuvfkT6BThaDb0XuKPEw0M+UWl5ANoj7tr0ExLpFbS/
VOy1S3H/ojNFJ5IL+xbHz0ZNbC5opxtYGGLto/bAvmnJyG9esIGfJIXyWYHcxbELgD5dO3TVAo6w
Q+cgkNcXq6JmwSyc6qArzTfFn+iS81DOlHLOVYa8AfdHnpzBptz/YNCRiWikoWiJQNmv6sV3xWyY
HJF53ZGpoB0BvyWkVebkHXM06dpd7sJwhgLd+uR6b8gNXU/uKFie3wcHjj+l34f7TeilMLXkIzcR
HIR9fMrdjVWNTg7kuuVzQmm+16aOtOFOLELN2PL/YL6objTuPzpMxxcVD696NxXDI4jNIta9IegW
MxDSAoGc9vGwDa1WECMIuHteY8RaNiWt7TLmqqN14bA3JJLrqHhMSGfDaYOXINtpsyi/J2sqJvnX
NuH3tDY2cbpC7vZkXLVo5ppzFF4T/b/DcrGZ6W7QrqlI58nd/K0dFttZOcE6mL6uKZ9sQ3422I+L
3O0uRLx2BW+ehZDgtAdi7Byb/RYyNoKkROKsR3/ZmTC7sQ/ejXd6e5jlz8X/jDXwtLbGnLl5ahlw
wZ4kfvLjjtQ+/FIpTWgxci30fRG7QOw11TSDz3JAewxICTyMSYhjdwFa2YXmjUcJZ+qaC7B9Pw99
2yojmi7ccgQbstc5k45N7yRJq2qqyr3dSZCJd9XQhev1S7ui+ERi/LXbwXwUWXvi3Yb+jL2xB9lc
sEo87tO3Xogrh4YdXxAuE4NV9vN5GcT1J8iAVpn/Cj98ZxpjGSZrrGE6QDARykjvmwBdemwAauZh
j2x7EMjVp7wjKUQGmjdVfEmDdKDPMSFR60k0shnXPdfi4hQVx64j9UQPmv/idKLtqliRVwhihGfB
BAr5JHTy7srvIuonu4KCEveNpmVvcmX8AuQG0EwkEhHaEzc+q6hhFN/o+WjvBwzSBiZxXKfIKiBz
mCphnMV9Ilztdpdqs6VnmIvTr1XGDEY3Hdhz9qU7lzYBrafLP5Si8QiR44jM97KPJOnfByI6hF7+
6W66QihxoQ+aGs8su8t2coIXoz3nFuwPa4aRXwmjN5aXKOLKZbOCN8Xts1foFymGCiSBh4uRBkzf
24TbFcU9/RY0LNICEBAr9SV/e3d39Arjw8QIV/TG+6TgruDgh6UVtRLXXwrK77DJ+HcZ2oeWx6s3
9lB1++MpJtkj6kX7ITxHJHRLsRVuHG9WPCvYZtrOg+hZq7TZOubhpl7XpNcqo3OLG8wzFxHSuOHo
CQUkHKXyKGhtnzcM6m7xWES6PRCfkdeHS7lRJLIj65ZGCYHFQzg5GRVGR96Tv698irKh21bgOecG
sbf2qDkJaJ0In2xUENaKAW8FyUxwu/CckBwyXDP+wQlfO0VYdHWLX0YkUHwKn7zW+ipQQ7wOUP1v
xorTnWDTUdVeAlCxc6qJw62GyJCburJ4gpUiLyMuRAYVRYbI5a8wpkAp0g8vLdr832xdpchJ/GZP
w3NiCFiqTGuTxH8ouqdGtdtudyifVawCtD8lz8WD1TMwfoz55izfULzsk9RJf88x5oHj3eQchHW2
lbCELcFEpAjCcWtSWNjpC5TvG6zF8x8gM+0Hv+ZEXMxKii2KTZ895qWZgHvrESUhfUR+YeSIaEl3
q23tG+VCZZJj+vj85So8mqqhHob48F37i58ckiMiccKlPq47XPAjMHnF6DTLG2tjAtnRh9X7tDO/
p5s/mPr4/jF+B283kOv17eKypCNnBne0wnBcipAvzWNKdRs+qhZtoty+3NXaSps+ZuTpeGJlQvZh
RRmP54KigPyCVGGkvsAC9vGIxsh8vMOyu0WaO8LkWopp9y7NzWxHBHIA2f54cBOCRrw0Zwwh9X/F
a8kl7ijxwLIxdV0hIAO3HVvEemPUt85bnk3PYy7Ng7jwFdoBDrxFyDpO7N5zklTHl7z1PFpWOvhF
dIyByz8AJJ60+Fg3LdbPIaeyvSV7l80W+2tJxj04VsMha3jZak5LXtusk1ufjkIet5jXe9yOZ9R5
sWCWhM/D6MuLKQM7FpqtFRhBQGYE6MAnk1HniOnBnKSHQm56UE5IS7DZDiG9hqlaRgsrjH8RBxvk
SGI/QP15VRE3KNiDb/SVJOBJJOTqvdJw4N/F0wyistG9vfSgG9YO//qK7yrKgi4vOFjwZ1jbSzee
b3aW7WJCknxGrYxvB5X1WIw2epodK6byZLlWIX4mnW4sscAyTxE6djiFxaSy5a7GNI5etEk0XUVA
xXDvWlGOoXrEIY0KsKLGUoxzI22VTeHLAv0+JCs0yYQfEG6B5j+tpv04LRNx229JdLGQ4UnFKaTN
NClJ//dR4eTXunTZ/VT8553YUH1iB9Dirr0UFd3iw29L7jYACLRjgZVx6G0M/CJBjwLexoxt/qS2
gJj61NdQZHMv+Qb5TnuNjkqh0oOfpGeXvt88EC6Oc30QkD5CCmnCZJYpLPPLzLbWQYrvl2i/FQLC
QeP+4F9r4tYPopjAzZCLBWavA7t7Tqq8z4W8VQeG7gRqFlNuhCBFLxmRixLQKyr/c8yD8CgSRjFZ
Gx6xv/72ah3cHbR5XRJ4Nlc7iiWgBGW3oJfv8yfXbWkk3CNvpHRvchoAIFB+SxQLbmfl5zvfhose
IMZRkmjAUehxOfBezmI5xo0v2Xhx/UIcD4dhT28+o/SMlBeZpx3AIGDUpXTtPCnYwg/u+MxvXH28
hDt6pMmU+pDFRUoHKNL2cbs/U8O7hk6xeGPdnVSDO6jeRDdAXywHVSqBtX1S6Rnq3d8KuiYME7hW
gtJV0sEil9+sjDzcLap8fE4bKaqoM70P4Q6SCNyQ1Qi9ZWLXM21jInmXZ3otCfs6VIBwcLiL95oU
JkHi6XykEp0Ik4na7Jhlt1rbqhXTijMWNHs6lW/8Iz/sOsTt3Kha08fJrlXHtBFa7Xpalb9+oOr1
xSlmmjH4MkjIfRw6HL6sidHb8P6D65RSoObmn+foDPPCwQ9EJF66D7qXKSJDfWp5256kTMts09Ph
CvgOWt96ogs1UjDOG8l3AMWZrr1Ig4NXhTg3SZti00k5ho4Ett20aO2w6IAJT6lYXqoUxQMubMLQ
4v544jq2/vpaHYUFIJUPnqVfxcYZgMYWs2TJHurXhi/TNdxf/T3oSUE/S+ox1VTN4twEuKYeHrKR
rZVqtUdny8yT3NThcoXipF1gXRnPkJGe/WYjwWHr1+a2QRYCQOnYMeKms5faCrqfWDzqRNBZTAyt
RoJGdsS9mvoCufD7peDUNOYQnoouIMJb+O8rLOTIabgK762oPmiyBK9qEmNauteZbYcLdF9rek7w
VoNBU5+BPn800/4BFxu6HfGOJhbQMxdcBD7GpIZfES8a7/1PVIEiAiDv0PcoitIpvSibSLvy++fC
9Yj0nEMTaLxvNIaayIQhSuM5nzJiJKALCYL10sasWOTXY5bJWBJbyoJHjaDC667VfzdklPntjqZW
TAYLWfAxWzBoRj8JQ5OFJNPdAClxXKVVTlxFP24ix9VE46VGKC8t01l7Fc+/ofY1oLwqVkwgamQY
cbeZjoalotSjvkyAUrfhJoLrSoFCve9JRignaGSu84wlna5G7TGpeeYE4jgUEOtWA4wPImyscjYf
UT7+2nn2RLsj49zI+xYes6tLYIdghiANYqvQR93//TR0oGGPbhF4E+SxauvTTzD40IOx/YWTpAUd
TXE2RQOTKAINfHZ5WR+pfQofQ5+jMlq5qJl17ajictQ0pqDF8PjFBd6WzkD0KDHFWLQPXVODzWtc
DrxUwpgerBxtu5kKZCNXYSWM4RWGQUZF+2+xVDI+XIr0zNIBIU8LvOnkAXsO32HXF7D/Pop5i5SA
dHrkIihh+ZKioECU3qO2pC6DThpN6uF1BS5FSSe+se5o6CN9mul1dkCbAAp3S9fFIqYGGkE1oWwD
HWktWiq4CoUQNf9yOMpMfqPye6iPzqtCMefBTakuEIjU4xpzfq9vnlukIKOPh8uW3f9BW1+Qp+Ug
7ZqKvcDO2lzTkQC75KTiTBXjZZorPfYWejIiTJJcOYehrT40bL8N0t6GntEBUwmAMciq40Ogv6iJ
/hW98yCivQJzcg0tE/a1uEPwV85u3x6q69j2KCkDURXPxivoyN1LSOQ0ufoWLYXHQeLD3TMlvVC7
GdrWILnRluRS0+Dr5kqzZKejym1GyboC+xRc9KvWoOaQ5oUyFIzMP5zidCLOCrclF/xfEb9sX9Oc
URRIgtHL7kPcyIDFp7CzVqOf8SPjcHWxoQ7SopWOQncT8e/gd/9Dcx5ywS0U4XqS9c1P2vIF4evd
qutoaKVUYDrJMqKYZiR+I59L6WcgyduvFecuaaGZ8nnloRrGas2jRLghFSyTxOPApgk08nt3f8cr
5Fd9/JPY6BapSVe9uH0kQffUcAiJ9N9KIN0yCrDfA0ifnHXJpTGkEfYPhN42mJq25psJrN0kQd5z
9EA6di/kxNAq3cmabBtGuXwtoFbgGzHyi9IsOTxd4mTp3tLETFJAhDXwZab6B127t9RMCNmKN+cn
Vf1t4owIpMbzqiF+PDiZCysOZ4/cGvblcRxn/kUaVIQ29R7aRtg6gumoV4mkpMPNi7cuJyGTepiG
kUAtQDIV4DY/TyQWPtj+ecXxrXy/MHEHY/4e7KFfChjIV7ff1bwMqfsdA6+LIEK4SR5khpf62Irw
yFn4cE/E71tPtW0/7inE323Tj251A7ZfWtJX9Khgu4xTLo0TCixOF5DAWyyREtZslE1eK7RO0Ydd
jTs6OFDH6k3HZzcH7CuvSywtuIVHSaMdIPTdvZg5tmSsUGxoxT6WkzCVsi29mrWxpOZzqNzez1xB
Xb1SjEhXKsfcvp2MeXCA0CZPLESIO6AB4rjtmcGXuM5oSCZjCF1gO8XLckQR1fbO+nUDqagAx1f2
VpC8+fEKv4ehLoSmoJ/XBYwVzrKfYDtb0IzfPHr/nfZy1+VmPKuGdBPrxqwA6S2k37j4u4Om4NH5
+hCDgDya1lxqyMZMIzMVf9N56NfBk/TruuLvlAHb4EwICdmDTh1j4OC2X/fX191XjvAqo3zYYbCY
HB3iv4XM87s28KT5gevdWZc848jU9mIKf4p5a8z1a5QS6T1ge7dzICLCabdTBpO5XATItXz5UCZ6
KtfrF0Ki5P1salF1tIAFsdHJusDCHGVIw4zk1DxiZoD+0kHSbluNn4rBounJOwcogbAFHBDi6MgC
q2/8crUdPbYN3teRQU+DFrb7EGMTnD7U/QKCUKdk8bek7k53Y5rSSy6YEnRHYDYUaqKg+DCvPKmL
IeWeKaRzV6Guq1FWnzuScm3ZxJEC0ioztBYiUNkWd2sXhL7tZyyd47POOgTujsxJNgXDzVKDtCxY
9mjL6haYbzaQt88fLZoZwpgzS1nAX0epux+U6c2F5gXD+8ZqOpK52fuPy7XG3JyV24vWcTf9aHeX
pNgUCgj1JDYukWdUkJBIscISUMsQXj7LIdfFRgiX2N1WYtnyZDcjYYFYwrKx+32708xj5hVymx+9
tmM4f6M7CFV54OC15sl0Q0/1s8qXVOsPy3VP6oKvA334WtAG1D3pDWumJlPDXEMZ8mAWjAxipEZ0
cNRe62292Po3pGXUru89e5WwZK72VUiIdUJUcIL8BV6E7of+jJcSR+7gf8pHfOXX4ET7/EAy8U1k
i+u4fAkaYy/ZZtHPvTbgxvxrpRfL5aEbqMd9xfaYChinhCMLXheYhDEVc5hutmrJXcpAWX+3ZysY
VkTHhG0f5nv1Cgq4tHHvyH+US+8RypEM1GogsZ5s/KJf1nkz6UUh25dj5R79knZKVB6m9wZ5fawA
KfHsmITN0BmU3jyUSn/MjbZi6Awsb9HWjJ/3dBEAQlJNsEkxr5T3NN40/osR8ILYE8/uIvC9J72x
LSHUgIjRRO2vEpbzHBo8Th+wgEDzKks4/lMnOPw3Z2O/yWX0a9/8iKquq1A4JAm/fcJDV4pqrqFx
2366klpNCDb86dWJZZOTEOERViPuQYLXVBXkFS0wLj+QlsUO42sIk0Yi7jLMl4hFy/t2vc8hqaOq
rIyctvgdC0srCwPBOUoVRBAwKhg2saeC/BYixQKKI0kDdBwVe43abtJBpt8Pq8vbRB4dY97f1Wk0
3m+F757tdUbBswxO7rj7nQsFN+KkmDjkeA+bFX6quEdZ+URKKdKqkyUsplbKH8veD+oPwxn3vcwI
Jt+xHbV+sRIqD3Aw75R+7CimukcPXaG9gAhDezWERQDMW6pV0duKoUCcsArB1VRG/P+KvOXDsmjG
/DeTm3Un/HoDQdnl4cRDlJTo5jpgt9glM/k44QJcc4xqTzyL/aWQYfQ0uyZiyY4LvAgnAYP2C7Ea
ziuwi2AgzlitXyuW/8M1ef0Tq5ATOJRtTiYJMl39WnfI/gqmSZJZ8eTuojArTAEPgXpJwvRtiCPN
z/hqweRACTOcU0XS8oTYiMh38tbUzvycDjEeRaRLhsRHEIilFStcDoctJaErxwKJ63a0FQvWQRk2
exgFL2Y7yPnU+QOxAX/0lXTq9LWRoeHbCvHb7JW6/hlEEnew3Jba+hCYgNp6XJlk33nnlWAayGoO
+Qo6LsI37Ykaa43o0qWaf9UY/XN1Ehr58LtDTXBu62D56B14lfFCsG+xaucFrr/J1HFXm6iz2vtz
QZFN7JNCY3CO6dTmMc68yosfvjgowdLiDQy3dwHG7coME9ZX4m2aFKiISPDEq/zZgCU0vPOCrFpl
S8L8u2+lJuO93C8j/AYoyzMukwOcLQLVVUYSWEUUHuwr3tADxtVVUShCHX5ClwMgH5+ssC+xHoIg
HT1NzJYP3t7Gj4v2qQweJtASNCUFRL6y+tpqBlC27zdUEWEnEgg3Yq9Aj5p1DBtBRp1zcFGNpntC
EXn+szyoSTRPU/QvmN46UtWkcaFse3LZYoCOHz8vA8y452c8pTRK/fBoKlBTPCHWdwJGKgPfN+qP
1REtnOt3cfGiZe1dMf19CinwhB6oKYjX5Q2D3a2pcLlAsxenUW2XUbtxe/EEbqd9NrN1Yadjd1sK
8AuwFlFw7uqh/KPL8KKB3rC57hHT+1h93UEOIjV1tWIuBIhfjkNL2GarYuL2ymAUbqBPkvPNY29l
ThszoU2lrHtI4gbjddSm9goood2fUrB4NaVFUNKiOe2Z62ZHCHNrWEJa7CBesSMdX6reg8yZfSJV
gjjTsJeH0ZG+8xCaAoVms49FGtpAxQvosOReNt8WzWnRRvrRX2zzH8Z5/NFRkeSF5Vhe2ut0qIbq
V01hlT5h0A9n1Jt6bo5CeVkQ8EYI3JSmTKWad2B6Y34Q0HgGA/G90dI/QbsOilBvddSArpBtCUMl
dzjz6ssKuCdC83XUkHniADsW+HB8cKa5lh0oF5zQmHhzrl4tjnynj+3Ez/0tf0rWDD2ihnBhCJvP
mWfeSpZSnZIUx8mT/5y4L2afP11/294nMHSqK3G5W8dyNMDIRPpdMN8A/N2O1eSqXIoGdzJ1oLaR
H/FANKGDwhJsyMKbG/zvOSiHCLVvRZv0lfiqCG7PVzyDnWAcFUTcxNQcc4L+Cu8Xz9c+tvy4y84A
plyckuF7UhhW4qvp03hxPp5YWu5zn+rzdxWEaPbHaJolfU5cdmn/cLaspxOfcSw661BaibIE7UcS
KUJT2FkmyehQSULH+4go2PH8fVLq/oxAeRjCm3/sdby27dKcEpO8lO7BoadpUIVZ2RhT+gER/Lfk
+j3ihRNt1/hqw8RTLxbQvCY55c6PX51H0v8ez6zYneMZLBUuoE3JxFKsf66+29hYK/JhtFNsS9/j
yIdAox0bvS7vhpeofbSs6wQJYtEiovES9TUZtwCDOpfnwZZ2f8oKnlLTytZg2dV9YpaMUjDfe5bk
ZEte9H3m/qS3dCH259fHMWJJ1/CxxzFOCB3LAx040MVbR17GPls2NAJUpEDF7vUUj6BExABTK77x
vHyoAg6ttG5bxVqhYmZOD6D3NHVGcIVwg67FXRUs9+bH/EBv/fAbwTW23esGt3ynEPXcgi+iAimC
DvtFjlcNBzdt59QW5HngDPu2/sMsf/e458VdOeegQQlafZw3I+UyBlxnDDrUNgDSsdGeOxH3bVhg
lTzrYLnBzlTbrcGjyi5cP8/sO0EtuUzdQR4t6o8V4uxsnnEdAFgwcBbSQqJte7UH9xwGSey7xLuy
QN+WVuGNhP4ZOr2FgvMsDLReBBBtOrfUZ0oJaSkKwLhamtv4+7r01LpyjZXCPIMGstzRD/FL5P0r
I9kUuTmhX914T8KiP6CksZqbiyuQfAq4pTYltFD5DM4xT21LVlgobst/G2JzLfvNw9CWxUf8VXxo
pIRECKQguEpvxKC8wv2m1LoyLRsY6XZTnXTbrzhhEMC5XzR0Ef0RgjLIUZ7zCDeIQ5x6XNMr75xr
Ym5acVFiERRizpuVoCRiKkdllOaEgPVz0keX8WHjSWz428MOneuZQgJiOT5XWpHgeWfaKAScaBdU
iwBsLZDddASaeNHnqGmZH/ltoxxq2DNT9cmU78K+zTHjA86vZUzUjPKZEYQt/Fodpo3YZd1Zwk7i
Gby11KGd4QilWGmOyd2K16EAVe5GjmcYiix33neb/vn/tf1uoY/CNrBdhNT8RGmCj87ALtfSnv7e
hdWsOGMk2+0Pzjzwm8WjnP/UMUTj7Xgv8i0NHLbWhf88z3UZNJAe8zZT5LS9oOFA7cT4dN73aB/G
fCb4nTsuhJc7OTF8azSX/8Tt1bwF9KgWMLS7IVBtNP5a1DngYwH0gt6ZRNfoChR5U8eFF4o8+CwN
E5W3I9hE2V+mBcLxbFiFK3GQqDUphxvHHlq25wLTW2tOji0BABVf58WwIErSW2cs+w/48Oj/MoFb
08+jYb8yDy3SeXRngVOE0srF/GSlNhP6BozVYCL+aC6WuU9jritJoLXcf1zKf9nXsFgiuZGpgZGa
JENU2nXDJDirqkPwOj4Qi3b7mAPfpI09buvx+O0th47nG549Sm6QJTgSSpvN7w7qu0T/uW4iY2EM
QxMux7ybmOViA5TZFSAYDBjcozJ/AEP2K5+qKuwlF/yX793tIUZnSLaQNjw2/BtI4xLabLem3KiI
60LA4oHL9m+1Up67dZ+COhJxmwAPOJ8IPH7p6QeASbOo7D5D5Yo9mWVQQK4T5bSMoXwAIBMyIN16
3O+zZDueKLiT00ADQQVSkEosSJU3m20notr3+hsj7g68CEZE+fkI06+uy/LfJEyQMGdfXDnxQWJd
8akihNuybxSUPPr78sKJIczPVlh4H1ccLGwSbgl0JwvTov3rFPGemKO6akUs2IxL0gPJxnBe1EC7
o2zV3Cm4S0/kq0ivSWuDssgWNgdRsnsj9pXTCm4QH6AFzOpVbhs6vhgZReaig+SrTeAiGSR1Qy6P
cMRUk15yhCSzfmBIcN69+MKCc2A+DYYs2cWULx15zkXtHtsQRlyjCBaYdI5JDJWZ1FZK5pnXoK50
ijzJDNDUdESBXRErAab34jqhJ1HqvMTSha70TQ5euES/6BWAPpifAZz4MCG9pS1Ad0PAgg10oEgw
1KMhb6HU5zMou6v3/Rz7OfFKKTfl8kre1UaH+TjPUNrou6YPWtBUMSDHLxKRMeb6DTPJG9I6KUgx
fUYv+xIQ7nJwwO8JE4mGiUJH8kVosYxiYt2bYS/MVB7OX0Q5Q1oIQIWQQhfcmhwX5QHok7xl3OJR
q/c94rsgTMtwMOO9+OSScKBv3qJR4y28B1WV2ex52DOkJGn9AKih2U/E+cT+g3lvsRq1Fbgi5KQZ
k8ON42o1nVQbWvPtbQE8koCST9rSxBzpvU18MFqaNqLJaejSLHrF1pAz5jZi5tA0nY7vvpAgdxMD
Hh7vJUNe1P4FK/2V296LaNLIfxq/ZXITfkzuYV7qfND4y35DLLt9pEomzhBw8pTz4DdzgCwYMgAL
9nPKCvD7BanZatN9o6xW6uRNefkDdit1dmbm6qlDxqlw8v4XFGJ7CH4w5TSbhKBbQVwedia3vkFl
PX/cXeJWs3FtT+v101NvSokoH8AZplBvnzJ/l3U4mU+x1Nm2ySGErXGJwiLzYhHrYMaJlObYgzy1
YPdHUipjZ8FH5mh92L6EERLgrdcLh4i+YFHnakQp1U/nFJKJBB21hH6vvx2gC0/gIbfkOKekwPLj
Z/t0ibSZbkFsKjqlOc4Pwyo87KETQg70XyuGeLLZfCs18fFPGc7d9sSVXJzxKfkrEaM1jSVdBuxl
Y+bWI/8WN31NiDVeoohwyZBLKqZVI5wCv4u3zH103MDgoAPWJuHRj9NZjv8gVMdvLG/YntRwatzO
j52xtQ/tqgiQlCQ5Q/p8j3FGXTsqhnoZ3ad400Us5RLM3sGxaKvdRcIZhol+oWyP7OUMU5C++FbG
Z3oJWKjlU6gZ0+j6OqCKFphrH0ypOykK2SjI6UjSvaYWdVoeqEiKPQSpEdLLSBUzYCDp2TScOkFv
gSwDt/gMWth2wM/V/xSjxfOuQVCuZ1Dcnj4/xtT+FiVKmprQWd7dkUbdfRszzyTHbtw+PkQZjh3f
BmymjuLn+Xc4lDhyl2EwmO28zsrC/6g9RZ1C3T4yQ4R3CdKAvfv/+MS88nrgdCcITdqB0hGMbVFV
E6yYe/HviEZlT6H8CxN5oA+GE3DYb0OdkVswZg8auGg+Lf8BJ1smeA223/lXjg/3+uU50AkdvFG1
Z4U9hQOwwDgovM3FMDOatdKgvowF2RciNhyCO3H5gjyuRqZL+GyCab01h41GctzfdWPKRcTwObQr
OxeOmAq6X9TvVdylqzvWpCy6olAYcb18ZX/VArdkMZXMNXpl3Dvq9nXUcN/QfmMmPRJ76dXlIwE4
Ke9EPhiQCu1DZ8Fw95/MIf1LFs/SN19eTX25zmEPZ0KVyQ8Pf9ba0apw04iFtN+wW2BfB1EqXoLX
h4eFe51IcfZjDYD55kBAE+vzKp6KCE4qXuZ0Gr/+WvIadxsdmlLzpb/VK+I0BmHCFSgsRVWLYrJW
MuFeln07shYL63/X9MVv1aOyMfTnfxsvQlg3xjzI61d/JVEGg11AAH2inJJJ6Q9QyDwVtI60QLR8
0Mcy6jtOeB6DbI9lwKGlBuf7ZDj/1fBRFszi7PrUMey41isZyX8ajYM1+ZAROZsl/6Q7CsomDpkf
LBNLwua2xMt8kUbcuswE1VagV0j67s15OMpJriA4V80KtRvRcvzb4VPD/i0PMK66HEXeV11gggZr
v5caK/+jgYAgL6OsY5TOcEvY++u5/3yTMxJp7y/1+eZXCu0ItFezVQgZzckkgOdaE8NA6byTv44f
EbSLl5IrRq+yXM+0jbHEnhTpUFd1DRXoWv1BFbtQCst9edtSmAT/CetYymt+6DM+2/1sEFJ4bgb/
jl3Jaa8LkE2t65Tu2xQ8by+7NXT4NravDcIgtdjAQbbBKq3A8fc5d8r9x0Q4eMBHCPni5mRUEEjB
LHrgLPDddxZCxF8b07JdLUcTErRoq3B5K92RUEFM3C6JV2LVdxebkvQszLNz3ce9OWxWf3tC9G50
aye4VvreHpqtNc7p+37j29cs2muma7nHtmTaKvb+9L/k9MxWRLOdBwZSZPAGHgDqaVlUpHCaeMNv
3Ly6XqMavyA9VwZ3TirUNKzYxw4yrE4tZCZhC+0xMFjrpmzJndaRnu7uJ1imKioQFZ/zD989wJFO
lx3CXITfEFNfywWUh0VjEh4hVmfkS6vJUvzb0ApVLnEgQTr9dVsDUT3IbH3Kzt9vlSdCz+JLMzbn
jgHWH8TEy3enVKbjjbS+r1VlgwVQgMVuhqIJJuHDlseCnh3rN1TRsGP7SUcBbvZku6hD6NOhi0jo
c4cGm7IwqWidyPvWYbxAIaMfC0rDj4XXVHarRgFO/nXJrwCD9EXZALN/lg9Hfh3KsG/scWRbWSHL
zKkCTKNCC2AxmVTUjhsK1p5kdc8c6zoVXBBJi/wIvnZVL8luLob84jNPBz06KWBTxPFSfQCvp7Y2
n+eXpM8zSwwfxVErSMA4aVMl4CiFSjEDG3lg2BhAxax9Mlt/adCVTidOkh97VPk7QS1m6G7h0zKi
Y5B3bvlqLniRzP913VUFCr/9KMIdotIA8T2ObOXdw6qaqsdyHtO8RA2t0Dj1jMtz7SMZmngr2AlQ
0HA0Vnji6RX471go1x5r+vuVRctoeCeqScQRWqAv+MOphLpiyveSgn29TicE2l1AA8SZ+hZOeDQk
OsRfDodTB/82NhgQOID9P2u69XneUiyxoBFk8Wdm5ymMWoRPJym5xnwWAtU/sLtTiBjtfW+TGtc/
bHGnj57KlYX5Dj9lPu23HnSxkL+d+GkNDy57PWrOQTn9Jm1b/nt0HCkk5emm/QL8xKBangezrLVq
ilVjYogcvVRQl39GcqKfkOkGMofwqcrtQnmyP+ZwmLdCdCGOA8vLiswT/ShyOgytzQaMqPmScppz
jo3iHANyGAvZ/cClZT6I4qNAv+MzSoPWqSDl7kyOADefQ4m17r6OqRqKpk86RWBuz25syf1RAeqy
pzcaN5bdFSPzl/wrjT0efhAKu67GHIE9pSCoHi625Qae1011y8O1jOgw1i4Dzg60YdyhPcQxd152
UPMcx9oRw/lFMl9sKIHNSQ6XxHQxC5WxYwlP3R/4TORHMz0qMb6fo9/NvaWjKpVBrNJuGFrPS0Tt
Ahr542DklsWVULRkIu9rvAqv8MVHeGWxaazjw9+NH1EgbjXYhIu1ZKSO1BpdveOQon0pWVGTaN/r
3s3w2zt5wpRRqlt1XUkFcmW3zh0zYnthc2Ok9jIvXjSCkUC0QI0BviDEzm3yCRs+cFo7oi3M6x2Y
VUr+DaL8hwCfdyAOQtjNubMfHR8AgdQ8S2lYhzXkzAvCeEmDxrvIja4piWRwyIvkwpDjP8IS/pYm
ltF77GQWRJF0uhh6VVyuIsftyTwfWC5lXP+EZp+oG9TTgxJYDOA7k6Wn7mzMLm0cwy7chKXaw09n
cBvfAhazkicfzSno1S7yZ4eQzVE53wL+tytbfhPOgk2XmAXnmYy/vIuR+Y3SQ2O5BFtRlYQi3fD6
+IvLJiZ+xv8EHA39jXArxIknBqXSTmqWv5/OxANeUDFG4q1WgP8Pm+St/h26iYWnb1XVwOtLu/p0
E34K+PHai5L6lRL8swCWfFcDHhviiKJCBluSkVtHKd4g+L/dTkGFXYreoK2wAmjwJPomsKeYDwze
f8Tfu4GQemDX2yYbhdX5odW5d7BQVPjxIS+haIC8vmaOkCC4QiR2UHMupYOWBEmz6VY41yAjw9qC
akzGcOXbT8v9mkwI13bKKPnxHbvI5tM2alm9bCDJ87/qs+WV7pcJIUBpf4Rgy0/Z8CY4fX8qgmrQ
cRW7uW3/PG6PkbeGFD0O5TqZxDAf01U6jRMSyZ+7pLMNn5wZjN7HzbmTp6jks/oNzDMdv9DaHuT2
vCCP9NGQYFP9qD26hRVcd4Cu90780fa9KiTGtDX0wuff6Q0tGnwwvsfAj11UN/CsoNw3L5Qgpcw6
4BVBW69LeTfv4ue0Lv+FldmQ9ztbqNZHdJmef1Kmof7ugI9XHa9CwmG0uBUak3NuzRIU0yYlxr2p
OqWj1yoOcGhQ95A0Km1fvoKNyxroZ+a/PmL3+lkb/ZSz+L9PMP8GWPu1vb0ULL/Y0oNFDijfH2VO
yw46Xwg0ZueVZf3o6KMwvAya9jR+68oX6xfMDdPkBOlmRpHr1U1qhBFMDrmp9TTc2RUrFAjbQSeM
iFm7fRBggvYY7dBtbcmQRiAaoAvtdkT1L15P95eoTtc3dcEP5AHWRzzuLz9fcESZ/Nc6rgHecw97
a+OM06p6hP10hJkR0hzLic8N7QdkQ56EPGixd42yRsSnBZtVeN4cXIPN2WbhUlIykGgcyYJZVItQ
rZlFRt5S4o/D4p+H9qxDvz1jxIet8LnMzX+EXSfB2GtGR4mzK7DT26l8pnDANgHINhWzTse5Pyf5
v/fIIDtXdt8lchdce5ZQ+xl/Eg46o1Hy+mtFZVRB1SuJrrL9sT6rPEGWNP1AsR4wm+trGRIs2TSO
vehSxYnpDN2s6qZuTPzlxPB10d4Qyk/xjqjf7Wx7TihJ8QvtQU4IuWjNb8d85lwXlxKqrEcDFB92
q1txqGwVPj7mYed9+BmrhKJIY+IK8hP489qTAL3+EGdGj27SPgwRlKp9eZljcpCTRacI/Mb9kP98
mSYJQxE6RNcld9s9QRm7SvnEQOur1iiXN85skWjMMK/zTVqEdpZnrhrM+cw3IabX/oabtl/FeOS5
VfDl3WGXmaJ98jSlk6SPQ8Ih7LqLlN63KjHYUt2XLNFGfC+jF6J9+dEQfF+81ShFlUPqLBWenrjp
tk9e/NVIPNJkMRhnZdkF8dxOsF7NCkkG4MwAKEfTR6suEsYh1wmZW8UHNvcJvqvse0IXz7qWGaj5
C1D56CNarlJ6z3mdVc1ldG6iRA7hnmtzjNWokn2mWnq72J2PPAcfpUuGiSxF/tlzDw7sLgqu6IlU
8Nfu4mATsdmIYpkgOEuK54fKnC4H7rs3HZ8wkdQA8BsWQh8/SUdn1WGlJ1AQXfS8qoVOZ3BspCsS
Lt5zfkm8h45a6f0uHa+DHfIjn6CEHxJrI9T2XQmxZ/HQoynHb4vEU4+0DoVBAHCc8ThhuPur+OJj
THkq4b+zi7i38/UEdnPL6+ph0uRPiDDYyVB2euW7WC/XUYkjgNIswb+/rZVnSgqGCKu4o+ag+fsw
Dsz7p+tG8Lt5S0iLkvecFFz3VjORSkMcv+QkJTHmROIA7iJ0uFlgUvBuAaaebjfJGdSG8fwoY9my
+FQFZ4fuKxHH9eyWU76a19jQllIDnKU+dlSRaVOwvqwTAY1wIPrJMsdBUbGW0C5yKfjgZSAJJHSy
FpOZAm5ZkxXO7FhDcZeYNli2IAL7tKb4iPN7feXi5Ay3a/7AJZ9Gx14V/mL4uHq7OwkBOzW5OzsP
ZAeFM9Pxr+Zed7qj9k0Qe7+OC/DBPLvOZsZs8v3D+8Wl18g++RYDBf6FTbODSC9rC+9c0l+wHt2z
HwfI8NyMgUPywxMwvAt6dsP/Ir8XCCVc1F4xQxxRw+aH0THk3UjrtuSTIu0bJMQJ5vmKaRvdz7HG
Kc/ivV+WVCTExn2EEWTEgNnbZJ4pstfYTsDeQSvzNw3DhSf42aAKGY1krXTUWv107WW4d8snc8S0
pXhGQ2V0IEv2Hyh/0LUVe0zD6O+iDNwOB9u/igrnPXEtEkt5AIMJR4zQyYfzDg1VCTuLh/vtEsfQ
Mma6E36I4cOryWhNr3aAr6/xPeU9cBJk44Br1dLvpfxbMfttz3ywDWyWafTRL+uzI6VZ9Nc+0plF
ZQOabRRLlGI9bixsjaSkLq6IfKvIYkW+HttEcfmr23JduE+6MDsg6XDMObJ67yFOAg7fKSddVGPW
uxcQ12yNQOj6aPk80TI3Q3PrVSRQf1GLFPjDJiFBNkk6xP2e7IP/7Vic4ACAvJT4e4Xfmw5Wcxbd
KS/0tygtaivg+RO1S89vUQ0TVYiqCXrBttgsNUZnzK5GdXzux5ZU7ZDdC5lwAdJMWKO4HKaC18SD
fxrMuPChACOOAFFCPQUSoUaNRuIiD8m+6xJhSzd7mDEWiZ803STjQHoGwCKZ2dGoeRm5Ks09XifE
porWCH9s0FJ8p5kRabH7Ek2M+pYbopGSzmNkrXYr3WnG1b+RIpo3kiF1bIPnehgvgIE7BnUgM/Wl
JO0M6U1rKQoxZmeFgrFPOSfz3wOtiiAlEIzeOSV9zdVXsbddeL+sUabM0C2c1oHQlEhOuuyZ95fM
v0kEqvxtVoLokO072m3huuezrBeU2utvzgLgMG6jaUwusFXqQdovAlljUF5UVyqBAAqqzUPtABW3
A7kAQoceYz0P1MFwC5LXcEMjhc6AhcQJ9aCrPtkG0YXvD+E2845KMgmp0PnUqkwqwTjNyRRG4vkh
MLL0c+166Rnzy4nK6w6EnkQIMylE0mdzNOfz2dK27Zch5o6qhEgcFhbLu1USFOj6kzUiK4U7dLKY
juNqgNPocr0H0MUjaGQUVk+mI04o/OU3uRzemXqMi0bNKoN6HHvGH2DCdWldDlsyBeThljOzO1HN
8WndN+OWKMuIaGHbMs2QeRHpJRPTi/FQrvCH1OMGF+OvT+8wVDkfeEgLJU9rloSk8U7CTc6YeP+8
o/aTZ/i4ulFt6Dq1uVJzP5oAyaqUOiopx+ZScrENUDrVjKpgIq4cRzsyxlCyTeyAT/B0azj4MQ1P
Fe+p6OFtUtSI3wYJcf7pPxdXxyWBE5+GCRnC8GADFbrxgxgmW0UU2CR/23Ky/e9JYuzoYX1TFwjB
rgC6k7cxvx3CD+ySBrs7wdjxe56LyR1JCmKTHGpmwpl0cW6FRGNjhOu4lNctF2Io3Cqk+TFgENZH
KhzI+MTeHFD5wvNT45nM24mxWlyfstK5rVG6cgQHQaRduSqY68Gp6nnZg8YJfESNnPsf2NYgr2s1
1wIV5xuoDgLWJS81ZTL3urSJZahG2sBSwejdnST5Bh+O1h8MusbNZ9Q0jUQ7Zy5MZtJFFePNDUv4
0xETaQJPPyT0NHuGib3j5/Qkslsd8mSFWy/CJQaHr8SyVElhe7Ud7l7mz86PZP9ZY8iIHcUDwTiT
FUwsvmU/ucAoFHV48bEYEjPwMgTbNfblc15MBU52J7L1ProxhSChYtZB0hlqOgIOUzbzdIWJimrf
hx/uFMb/8LRFUKl+Les5GD4YMDnJqr3YJxVRNRZEJiKDwfNqLSohcZN87iy765YG+sF/BJMyUrHq
eaDNbfbVVTXiCxdrKNr0iJiPxYfoyvVus2dmwgWNqlqxkCFzR63VopnWp7bLuOsZTZLQxdvY29oK
IGqTYM0jFQLOZ5EDHzAAIDW3276yiaHykWxdveP/APymVPJ28L1lnOwoqqfgvFHb+5b8arro5lM7
ib6BPCceaMz7/P+eMDqaoWoOOw2rSkAOP4fnuXPvOaTm9iKQoXzMXVNmZYhrzzx/kVsxf5ySig7A
CNAQLvA6g1J7n42NHSXg46EMoXZ4wl6ejJIaRbNmB9BtWBxMq5I3JX5B4EzpuSg3V/E5MQztA2vH
/XMn0uKn6lJMsaWvlgS+OD8tsz/AIPhSbYiK2wVmuM7ODeEBGJGXmTg3Vb8ZQdRxJB2yR9swIWB9
28AhYX1JPZKPRpYe0XCtMS5fJVDsoIfA0vJnavvlnZuf9nMPdccDShrETpS9D/o7Y2z4K/msdNj0
kDnFP+hycU6deQJQ1NX12/9o5UnEEkryfvzzx0idDTIMh5YFo/8/kiUdXgRZmeaE+G9RU3H0vpbU
WEskHefEFYYB3q4IBxjDFInjLLYowT3IubV/8oHIO5BqqZlw1Thqi3zV1FjunVO3kyVvUtBQbua8
ZwXtpnOmvIioWkJ4EoUkAkhDN91TNUjc7Dccp1w29qy2J1X6T694hi82plfI1tNgSKBkOXN53978
aKz7Q1z6BHjbTNkOwRUkXdGcoFK82iU7EKOsoOA36gK7FKkgwAM+BoamgZyfA3RwJ3Vy9igox4b/
FFmuQoQAKCxOwapGfaYy2/9Yr1bPeWKYxM368q51XTMTRcn6B7kNz1Q5WT0tfQqXSLAb+JtBeykf
rQGG3xcotSNddLvfqh/Aw6m10oHeeJrHVQTgFv65giLuaLCdnQkIRW5zFXR6XokztPfzKcLt8z48
djSEv9r3b609qmeI1jNvjl1RMsRuugT7bCBw79yx4NqmIRCsQbAUIkmj9hLM8R6F+QXfj36cXsTr
iTtkCCpWU3fqjy3vkOM7+0Cv/NkSHSEaCrmiBCv1fXh8flaw77KiYZhACo5l04wdbw78CN/MHTbu
JgdKwSq28S2QtPAN+WECLsRbQE5dYpwx6xsGjsC7NomRg6BPlFgoWY1k+Rg+hZvRA5PtAuhlE65r
59UmiwRCMlwHoVFi2I/clBHuNSWrwVRwIUolJ7P8VeXQ5S3W2WiFm3an5wUI+FyKvPvker6cMOmu
Ckr4erNWtNshu6gFHcT+2OndxOJDp3VZG/500z9EdZ6rvo4/IB6X9iZap3mgevjkdyXDuBN3TY++
wajP1ZYY19b1BjmjfW4zJV2iUI8mouJMrr2FirgWR4SDngg0AUpOUz0azJxDGcVjrcDwO9J4KX6x
n9bi7GRQ4SAqpoMJ5AZEcp7sT7Rfm2htc1XatdbZk1E+bH84EJ4+k0yC/xoeG5NOpwMKphK8mfFb
CoJg37/LwWSW6zYvQr4mCFDhAC2kCFFA1P2EnLLU6dzZOVO8fllpAn6XY7cwQ47GCD3qGGLJfmCp
EWRfo8BBRH4OwyDnXpTp7Pd2WaUzTNwfMN5cYSxecucsWTDPTg9e7a5TThZTo4Kc69wKg3EAhTVq
JbRWyVM/6zI6iCE4nOwwr70yHAnI/MoLoL47mqfAK5cX6EmgAnxAENa4RzZP7D9BsMYZ2pM9C+YB
HpGRaF3koLllI/Yf3bhLWSN//ZfU/DJqfSGcnD/a4ta26Y2DJq6K3EnF5pU1CU+b4O044z+02LWR
4ecjDB+0QD3oFhKtLMTHhv6t0uV8vqCsd3mKE2BrZsaVBRzJYgsKkMlhFUOdrH6dCIOt5Sni7ogM
NFk1llXWn61vlIkjtjQzjkblwYl1fXnheMKBS7KrtsyOyITl/N2J+ZeW8qXgftpM7rBhWDfYiw9Z
eAI5HpivhOdKoQNdT7CyZc/T7eBVA0nDsdZ5TgDe1OzOypqhUVAR3Num9oJYlqhiFwMA9B/7H5kA
4Dd+tGp2qIsJp2+DJstqA79jIgdSdm0QjXHEB8Vkn4iup+y1kgSwKMLDNmmmoiMWEX/Vawf5pV23
G+qUs4QZBX7jbPxH0wMCuNexOiNdSzzvkB89AkLjqZc4iMe0dzTVR/eJHUTgPJM14VRPilk/ofAw
q1ApvaEByLWUdyRjXyqyztFcXB9GpuYKid6cnV4rRn7V2HE+bbi5Vs3CPMrW36dCnr3MmBYzhfv0
x2rjXoAUxj77cDwUb5XHKfkiyfcQHH3L1kyfkPZQ6bYWxzPqt9+qgTGWYQmx1mX+gsDc2Gzt1wH7
F02sL3MrIhDLoS3wqo+icFSgxDg5P3eHtVg8ijDsBAtN+ishT3+WuA/G75A3ttHzqzo+Ktd4vTMm
BtFhDGhM3zPrVenTEe0nSFsX4MhI6xmFKpT7ulMODu1t2M8HEyWDshvqv68plnLc9ux/ojcBPn9F
GhZca/HL6MMNpuWhstHI57X7a6rWfEjdAd5Qo3R69N4s10+XLoaEV6lej8FJrD2O4zDQz8HJI4P/
YV8lEmst/aE/SBJua7fHY0fNGPnKAC7DUYvwehtD0Y4MYi098miuNSC0BJVpnTX/JzeTqJ1QDGk8
X5mTujnKWwQmxQ6qrbDIVe13gz7A5I5yjXeS6TeivPT+DXAR39zBwHZntXW16mL90yMzr0q9xJUj
RQxGCi0u6ecsIip6UJXyzytQs0tDfXX7V15N6aSWE4owdpAtFGNRyF4peb579Y2Xv2jEcdCzsfD/
lrqbKK0g/iLR2oVeIhctazi1F362kzSW3TPs//AlFCizt+UvLCuyln17Pp0FaPG3PTVU75ap/gpi
fpml8PLiZsXTlKaH73VILawNW2feNcarzn4zlcvXaE6XuN62y5T1poO24rCrFSu0MMjg7fmDojjo
p5hXTv+QdY0RDPKGxZvhx1suLnF2B71+bj4Knh0OfxtxU2sIMYhXAZ/bFtAqeIRjb1DBRSNOdxzt
aH8kL5UX14iPW1xVQ71W2o6t4tH32g197buJ/lK7P/Z9+YI5n6f6D4N2vwdrlem1sMJe7CO6cl8A
WkDMaOWXXVwGe9DJI+yt7QojQR2nfCZXPTaCMjbNz175VZdQLvpT6ggU862cKeECxHvp1BdC7jsj
hRJ5kdDJvKMfYr1sHhmo6SrMQ0vLRtaGtxvEw9WNI5/+vEDjZLGIpHgJFnJcbIv1bjf8bvJuw5CL
rhGAY2xqMceNBGxGLuUojIX1vZClB/PPKPbKZJxpVduV9t58mN1drueJSK04AF0GeSDqL7lATt0V
uCsBH4b0N0yovkyueXwPkX7SADIZGKwAgGi4FxKRpWFgLgXUVi4YNcEBhnrNfFLMJqgc5JFXcRci
FmUDk6agK1N2o9KB1z+J+gb+HF6rc1f4zMsM3mS5Kq6bWDZEaASOrnLM4PjRTYVeasJ8GTlvRX9x
4aW4gdrmFxwRKcxyQ+9+RU1sTc0OyMHITBmgFJJtd9K1mbM9gEo4RlpwentMgd8J+cdrYUN0qk1b
ZzZKHS+MvvJyUReExTrs0+6ZwyR2u+uEv11MNMiVsmfsEkR1waAr7Jnaxoj1iRKnPa4O778xXCt4
KjVx57ZiB3ULYJMuKdmCWdgSofD+9OPf7aps8LONRN7U+9+dgxHpdnGcGLHZV1nuq0qSAgfhn4Aq
wpO2fLQr+p41Ic4Zt5mz4WPWHM42/H8GnKy/XEc6RnjpQKrpT1hkXd5gp0h1vxvt0OT/SqI7r+lz
gofR4MJaGoKDb2QMf/lW7wdvV7WQETCNLKUnozIMNLukhEqdC4QJbo2gz4cS4FjTDUZe2c2iAbpn
3qPJ+z1Mv4iuMUEwwOc0CRdWTEqYFlBbipB7Fj9FLqbFL8eibYV1hiloUPYwy1/vcQdk63mf8opg
SiEsbreMVnemKLaO58flzvgkJSRVED00wVKCBYf1LJZF1On4VctMawHOClfoWdNwtXaWj7V7qoC+
SmjWbwUqjPbH2erpWVhOKvoZVuCJvleFcp0yGOO2KUm5/oWuoTwcDmPDbJ+nh3LjgJvUbP+jv4qz
GSmDp4mwql+9VkfEGkv3kcSbaN5Y4jaGIIPzNogwXtrT7q9SZim8cGU5jTs2SgD8DICbWxYhHToO
cmICOf7vgW1HICiTiLThVKszDzzMd46F/Vf9p7T2ZFHeRKznvL3YQEK22iEqRa8JpJDmUyq8e1ss
mHR8qv9qJi2CWhQ0N+kHSITKCQ9zS/Fm6VLut43XYlDJJ1UT35EBdO4bF6+0Zs5yZP+ZHTNEwpx6
sBdK5tF2PLtzakLazY+WspJqnwDW/0nYpCpc5eI7TTOM46nAbnFYXLKC9cN8Sg1+UjVFfp97ld7Q
9hGjLHzsfWNGu4K9lCH0wdyurzA67C23anPK89iW7OYKE7GAd+HQ/9iPClOWHx+VjvN+7bRI5flv
YywAik5NxHVz9CxxzUfhCTT/k8d0/BlNc594hIh0yOD9Md4PGIX3ANj/nyBQvfgYYd4Qqb73U5Kw
OAo2vIRlK9ja1z1q7M/CcelpHNW5lKmCGKtSfwj2YkQ4VDdFo4En5v+LZCHDLW0+l36B1z9p3ngQ
UYdmZgQdJ+GWEVtg60cBDLg+u/0f0tKypgacW+A9EZA0TYz2XCI1qwJwbLMq0BApAtXiofwQX5D5
1iKMHvVI0LXyIKPNEAVPj7pMb9jWZNYtEh73b4CxibQb3OoEbaTXLE4h44NhIIeL07A119BxgAcH
1XWSFGEcYvAURKDid4GLJRRBM2JLFh1RFIkgmmwrZYPnCnjEKCIEhLhdsaD3/KOmh2WmOkSXGwDK
Rn9HRlddW5G9JbJeU1W4FRpx9zDBiavnPGJK4D8Q0gcRuUOD0cJ6Gx2zSTAoc7g43wSDn4HlMXiL
fI60BTZygjzdaPdzFvHahSFeu+6GSYU4Q7ng4x6oo0K8Tj6tzjWjOGu4VyCw8ZFTBVRvE9ZuBVVJ
+UF8xOfppfzZEVwr8LeP7JzK0Hf/f9wpDux6hllMdVu0PZK8bgON7/DEcaxTuuaFBDJu4YWfiy4D
cc6G7pOp3mVeEt+JnxujIGzUldjhY1hsIc5rwATENsBqajWnEt777StpX1sAnhAVU9jAMjoEQfmk
MbDwypW8Sz/qEDlRRi1s126IPn90UVRTpD9oagZL06WAWIIXwh/8EiRtrpw8Q0HL2vRLdzIy9EJM
p0zoMcve4+vcdLqMVgjLhz59VnuXiUWKFdBd1hi9i2Tv4shoyTuJ1O02vBAfYf13S0DxwDKaWATe
s23wwSFC96vQApysctWmjcpIgwbs9hPD1PYWpO0qVsoQoI502I2sZElRni0EUWiD6ZPHSNc0Hi3d
JBIcB55jtJ5zLMupBcfbulo7dPnGP6I43/GLorgwRQ1WlN+WF6vf+rWDJzoF2oTV870+JTWeK4af
FIRRfDDqKrtHsNoX0l7n9wn3CUalfsSvcv63rNZPt7/2/FOr6zVx8GH4cRap1wfbuD0CR9MlXaFs
+9J/BkoxFMxgf0JEaE0XpLrrvNzyq9y+uTePiEF0M4qOUSA/BfxdVV+a/1OlkgRSCJDehXGOk2jO
ByPlSgzQoTd8ZyieWm5SJbVn4S0af8ZgEhZg7ClYOV/oQESSL1vWoJllyFB0IYpP/5Xvll1mBE+4
BUsI3olcoi0GTzdsJzt8Wa8S37QMp0aniK31WZrm/BH/UxXysYa2E9BFmDXx4Xdat8eLHE5QlwuV
upwQHLslwliz2WsERr5QTdYeJ4Ua08e2Ag83xeB/ahEDtGVMdU0NSLZ1Lko3BaZcumE8GnkLdJBW
YidbA6OuO3P05IQVaD4zUz9tRp+v0n0sq0VbCqgFt4kHsxL4JFlnD5xvg+JjT52evvcbO62V399K
muwLz1nVZxgvxj7vZIJ5rw2Nx9XZBRcBFv36zKdu4yrynw2TqjKCG38s135GQqhhJTfnlcK65vc9
tnPZsAPlJ+j/82SkeCTQdDTW8kODeFSUop73Ba+LpJh8svd3u6aPITpOiVkcAzWU4RRPTXKSEVad
QuVFhJnuNbYE8czy7o7QxpKfB6pUwpUFtVrCJUCfgl38JsCrdGKRwHyV5oNVBI24huaEvJMkJ5+6
F33qT6REAs53CBiOwAkN5rUNmoIAx6efC5oimgoETn0iweowGpimVx94TlYF+j4us9qmBRIBpZO7
qtDibbgosIsqFXmZVN852tnHaJnzFBLzFQKjNpWxzh062+8jUq8e/yoAhyyXLWXwkKZjvslURRf/
qsG0jIo/5hEQKmQn5UI/OC+hDfaG2N/RKxaRrM/Zq3yJrrGGUbkUhq+mGa1jQOWfFfOXKvkHaoy0
DOnMJc0pDni+P59ogWnxs9bLyATeHY5vf75SnsR45JWFMUufLciOWi6PKLY5B+IlLIxc1OsVYsHg
VG2U7QqtCXGNCwn9SyWYUSScZ4K+LU9FY/Wfx3CIw81F9zMz/IbRVlFmw/Mi4yHjheG0UO+nfJz/
rhzgHROEcJYnwTS2fvy73FAeNHBsJL+SA89PAJinSayuzKZOoT8lxjtzYT1SIl9v7DhENGwb7ec1
loLXwsl0JFmCz+jeIQQyf8EcLmnqWayWdqoZ/rtMV/kFo5scTlumq/A14L+Y07zxLkIWL6PwFNAT
0wKxWe/nm9ZIuOK9uaTQjDxaloztec29lJlGGwF1R7SGne7c8MZFlk3ezSlyYIYd8qxPOtvymiNu
pswH1MHEEZZ8pubjF+JNj8RQMNAFaZPdH9rRGuQCY1Dc2mo1F/aQ+0WB2VH8xXU+dENJy8V535R/
71d1Jnv04a44DAu8dPQXW4gd0E4ITqk58+x+Zo4q05ktElES24ZqqPVfRP5nSZgRZkZuu9Vb2yiL
jsgBNA4w42xe0S/oRunapwkfI4WQisX4pfa2ChhA/yH48oq/H/SuRTFmpcobeDUdpCkwxhi574iA
S7GvQIBtsnn5xCJeXtGQmyrJO4fjyD6mHc3iUGxw/Sa/aR6QSE9UGOza9fMxTaoO9HZD+xkc6OCA
lNO/1obRP7nOwQoTZva6ncchAY7LHBzmeuJcKvpKfGw7d38AaD8yI4QudsMNyz0mb25pNTWxD/1E
y/VElX2hCxeSoOwqWs5P62/I2YLKgk8yqo2TNYrY5OGZPweU6Y+SC9/wWxojASlRY7chrpuIji8n
cZPQCGLNlSQjY+69SoeM7jMc7xS/x/0tpFkg2MfjPAXkPQbg3peV7rGU0zT2Ao2rHtn/tldTCpYT
ugFrtCK78FQ0GgMJAYf6K5z3uOIHGsU2TbN2TvUmt3AraLxeqnZ0M/T66SXCTVqrcNIfGWd+jQPy
Fud59y9WYi0bnM9vOtWAQC0rztJJNGFf0ZK+Sw93srnDWn0HDodBjskTt5+0cvjhQtPAja/2DhZt
hJVscsShFx4lFakjKczTDo5adBkgy2WxkplN7vQG/7SWTAno9bHiT3muBnRjZuUYMyndwkRihlcL
hsPkRWHelq5urBJ2IlLURLAs3aUDluAYOjuIN7BV510fvewKbleHYjarloYld0GoobhZBTe2rNsm
KavRyFrDKaTukYtZSeAGaH3PTzABOKTC8iW/R2G74Qsan5Ac5UVwmEj5BOdsdrDm0SZpDzD/MCIc
khrwCFfQzNDH+1utv+GKz7NDkJOvEO1Y9HzubeKo+qOGTifZMf/kB1Wiz20gsvYgLLdLsFXaZW+y
LaR4xfkx2c0o6zvHXt7yRwGnvCEQlX4ccZP5Cy59UG13F/okF4pe+jqyem7o6stjZbcor3CpBxUP
mFdxWJNeucKQ4I+9a60vsDzZf1XKJli4LFlpJiAmn2ktKkYrw7GE9Usi21fEb2Yx1gwIVIzg4YnA
0h5YPhYGNXxXZvMy/ckoUa3FXsEBN9XkRr9hmD5cpIJz8NW+hRqGrOsVtRBSuMQ4NPDFR/rNFy2z
YJqpx/pmGAfxqvmKmHBzl5vFfw4W1qqCHNjHg+nIB4FSLcubWgcQYPDMMs+QYwXR1lDsmP535zV+
ORQKZXHv/Bo6gXA+DOaFGvlAowjZI9icEYKIXlnNvn+K1iPPB+yQqVBYBF/VxYak0WCXTQ3Y0XNR
Jh+3NJx8NMMoJUq7+4rzN+AISCHImm2oU5TGt7xQrzxv0kPhFrJLLHek7oOEpNbUemw15dLswSKX
kRv9hzldGdjxXgMK53LjzjgQjgdWNhN0agYW9rQy78QTvmCdcF7FiFY5RZvKlcGCOc/KQeHrBqg5
YZjGNPXVvOL4pjoQul1zUmm8vwX0C+71WF8tWTpo7/aU/2Ci/wu3J5PU4U9zrkka0ZtDbo58KJjg
H1ahJZk4Uzx3etthvjlpkFRmuPrnZZFO0/asJy5C7zAnh66u6tJJlThu5wm5PZP9b1o48sahHMkJ
atcP2DdixvuVE9+rL+9IJElXG2nZcCWBHXzdClFVU6dbJTGeNT4XRBCf4Noxse7pU34l/IugWHmg
j5+S35bv8ieiunRoXvx04B2nwQU4LksQNPJ4hixe1qlKhMfHwADrcX9oxbjaZ8BdvhLSJ4yJOYEh
XefQkLLFZ8J+MPIHBNmLBp4M+svTIK1gzGlXWgRX5bD3k8dJ9h8UIZpy3edqGSpmSgAHouaatpSk
1dba87Tc7zSbKj7IG60Jyd9woDYyw6ZGOTD+ybZ8ABCFFc9/PFuXT4Ti7fbdQUhBdUvn4wQNrZmG
Z2DevgZfrkEa5e4L7wpXeIXZl9p7bTELBkHXnNDnL6Js8K9Im+dk06Z0p6p4Rl3Abhn/zdND19Yx
Q+WBGL079l1B3l08MnX4V4myIzD/EcLtMKqFfk9GdSWRITzcvXVc91jIBfo2dbgGnTOxBT0lQLB7
FMuu1Oh9B3PROQuEmA15MDuW5IuDJmt/RzC3Sy+qhp3p4IkCneld9uZPaEdJKCxqhZPUYulxYvtY
BUhEjZpvuT0joGx37hD8Hku94a0aY/Kx2SqhUomzFr5G/xHkCHk6zp5YxLsfDqtmsH4oozsT5pP4
Ee/d/J2g9mUixKMyoblPr0bgkkXiF0lXmhJEVGa0oC8/lo2DUqvujvF/BCGOKTJ/Z3hnL1wuQfCS
b8QVnRq5Yt+iadSqZKEUGqho4fwj2Ckd8ctO0Uk/mM1HJTrShBdS2Ad+wLQermLiCShBSuX7vnJO
0qLRaqwLMd1cMob+HICvMtxp3iU5FMp2tioNKrwAjXuhP3oLZlcqD0HOGi3B0NFhEo45XZaaXd1i
m6+f/awWH2YrkQtjVxsNbMT3tHLA2k1MTzSrcwVgV/OiPfg66kn+XEDszvC+8hyN/jb8Wg9cfx4j
EDNJcUQBBwbgT9epyLszzLp6wHSdVT0lxRpfXqyeUgL2OemO7LUlEW5CTtHnoQCLjIQTZuUCKgSU
7Vilkn+0sMkByGmAzJXmrigqPF9ld6byRE4+BOKZ9O+3skehELHwvC+F+akdG0nRYfF74bYV4/dD
TWJYCLWdwNHHfwmqJVR26vf4dHINjEYxfRYkK5cLpCM0MN1R+D8iax1RJoBgI/KsWB6Vo1tRzKH3
V7rbZvsw0BF4TqYDUENEEPTAbN6pd50nV5WBs6VxxzWmkF6KV4xjG2DzA1AndxTdGKZNJyo7TF51
6Lk53Lwcx8k+fBOsrXE/9iJfU4qmycV0PfFWikFn787HbcuWwpZiGDxVw2T9AN5Ty0eA4I/+z871
wx+q/FVS9o2EVJjm7j7Q48vnzkC7VGMudTdJNpHb9R6Pc488bzO7rf5rfki7Yl9glSy0WiLNbbeY
SPxoSB9ernZRohRVCMnivhTJ48OaDWy6iOGpv8px2cGLyp5D5wH8TqQhJz4kFEO6xeg/xXx8Rs6I
FRYJd8MCHz+ouCros/JEJJHHmxtUzsNOcVZTfnePJGg2XXyVjJ5JY/SmD1Q/mM/1BpT/qY3Kbb+C
c1YnMLKPT4qK2nR73kuZmMhTPUC5Y2uoNEDYoAy/vnBQ1Vbpa+dZvBtqvBz7UQJW9IZ8tnctXccd
3JnwbxLcEVAuHSISnGkSrNL8rUzmcHB92lnU8yrYoQswyPoH3ODOk5E2v7wuCVl/oTS0K2O636vL
ksY/UDgFpibbqt205SafaLg9GPvCPxd/4yCzWewrW8pEVtE7kVc8t0CB88KM+7bAdS3lV/SgdsmG
tOoCMyuZq42LoOVGcrIFcp0PS6j+jzUYdXFUQ2Ktv7xPZq1w/JdxwaRrwlTHkppg+mX1uQEUhjYZ
oOmkxTjNk6YMCextM9GEhc9+GbfPqpem/kPvHjvyMsEAp5avk5DcDVhc38h7PDj9I6amaoS30d0M
UYMttPtpYedPYZdU1G095LMjFHIZhudmMluHdAWRS10bQEYhfXPglfWNoAIUzjizU8nW8dxvHa0I
TTaf3afYtOJoxcTrl44IoeWrjeNiOmTjYVVY41JxrilML+9yUDH1LHQcp8zueb64WZ4EhuDu8bjs
HJmt4wtHAUVxUwMrwqPXQT9YFkYimWZ8juDdLfcaYfxG4FriNUUFzg2lbPcKMPdjvKRa0O2zAW4X
yUFVqa5mXptO17FY98JgJiOBN204LAHSOP0cWuzgj5mfUUb+rWr0Ah45QDXfCq7W4UU9BRFo6yKU
W6Z7VPOcc1EJ3ZJzJRsS0szGBWQwiv5+xpgg48da9ilcUHI7or6XTWLL167o+NL4TCckLtnWnncv
bNJDkmkYUOIFCrwBXYH003d4YI3CxHgjy9Yq6zQMZNabjJ20HEM04CwzXi7sHF+9mufWVllgNX8L
4+hJ8nqWFQb1Z0ZjNvXSOgI7UByM1rMfJc8zglKS6xGVw3vSfDiy/OhRTZEf1C8SZlG/CIJB4VKo
REmtlYJ+n4bUPNlMGwX1vjGDbStXlwt5yh94TNhxBpJBcXXh7vz5ENrZYL9UK93IStzY0CJZ/iWg
m7p0ygqFABchFciLR3Sr0aevNcYPp0I6t1fTwFlkm2NP1Cf++c0DXb1sUdGuyGm1KI2mcmQmfaJd
1KsMgCLFmmgMo1AugEqKXe+1ttJGwMUisrG71MyhvYNQgF7imYktk+zwJROUw8VcDXDIuVZH4tzL
Altsw745mYlb6uB+uFgMQlyPw14ychUUh3oUw+uOQhsaS0WUR+/+9sPHc3D1iGuO8cYDODkf8urh
WJx75FYZEy7RveQgy9eic/vg/xjk95ljFPqErgpCjBoARPY6Q/CF5naCW9/6XLSPC1O7q7973bCY
9Ad+gu14FTnG1++q4BCGeQWxliGktrDaMIzrdMPoez3s94o29aIafYVMSvQYymDxk5ybRtqZGCt4
XKfDL0pJ+TF+t2mIqpcTtSjqPDplGz56M1vDS8H6RIym3zzp5dzLISlYD9LNozMqb+gzdkAD5GIy
UDPFBzV5W2QekflEkR52iYGjADAQdVO8IQuGIXy3wN4Ct3OIEazKz8opxwRtRBGxQQqF4n+gK/U6
NZ4AJhl3OTVgnUj532nvQr75XUiTa7zU+R4xSvTiQHGeJi+FXIxY0TbHF7FMA3ofSkF5T6KHsYMm
1ANuOjWAPGZVTZbXcKotAt7uIffrtRue752RqM0II4wwDRcui3h6W3it5QeEwacSFczzLX6HSLFe
UDFCSzSXsR9ttQPMKnbXJ6dQKOFXmiEy8IFgvPkRF+RDLH5GEuoWFRkUntaL67gY+BEKOdMEg5i1
UROoRG67pRjRJ1GKMSk8VOJiglq+0NrsAgnSHhv51KDuKaj4V3uqv1bxokc12QatYkYDGIjXQ3aq
faNk9fiAZEhU89H25uMbZPTUpCVAgzs9niXW5XENbFtep69/idXYzmqsR7+KR5BUFgadOVQYCwoL
VNpATv/dQJAKaBQxrvQmS4FkvXqTEUavY6jmJcXOg4zdN8F0JJBpNMpYTU6ILJJKEfnLi6KBtPS3
Q2lLXS2FDF25f6UOkp0eGg6EjaL/hc8Vrj5suRtWAiMCkLng+VOOEuqzTHtTgZgjYJoS7mzd5Bt4
N9gfDiVtwDZtVlGYnWoG+S04fGjMS4JnCoukhRlfkgLA/ef8CtJJvdhRxUkk50QtGOuhgtRnjanr
JLrRhNoLEnDuiua3ghM28aruboXDBA89spKk9Pi3jl7W5kO6XyXKDP2yHi8YZOUgdSu3zlxJx9xK
SQfo11mh6K4hRXGoHv7WBW2FIPBPP3bQaNkEyqXLPnntUxF3Xllr5fGqAiha+xIqHJvsCEpSJckq
4qPKPENEIO+gaqhk+yr4WNkT8GIkOl/zWeP55ryYF7I5uatoBZsZ8Hm0wJ0wSRHS6zCikA1jMe0/
VFrxeDExE4NRHWtoKptYY+28NcXm2JRJAfH3DoZ+T6KilnZZLJhLdnr/B1VOy0EFsdzAizp1RPYH
oyjrYXRZRVl6wPatrvbgKdiWhCEXy56lcGOlTTBu1uUUa+bPejl2M/gTjh678G/K2f8tWYUmg3mE
kcWxP7L1ZKmTT7uOwUpmxIIKpSdYm8KvQwMX69ValtBKSN1zuXQ6ZmAFZkHfvy2qwQkYVeZEt6g1
AIOMb9n+WANaPm9//3Pd6h0myWv0BAfJGYrUaAAldhDsBkian11RoqCVFtQ5Y38XdaQvLjorzZKt
S3hkx0LijeDa80ff1BfSNn5u75WAb+TEpAC5+AioGleESZvdrhnforn0EQo9tIKOjQ6ahlBTJ773
a1Yf15lCYTD0fJgGwFbEbiqhkpBYmvR2qZUxFTFt4KqTVhsP99egIX83u7iXbZXiYSv4eFOacs9a
avp/dXr2/pAtWYI9qMZ7vEw/A8zoUfnJF3s/k0aVc1ioBeQZePa+z/JDiDFv1nmGog31Ff9S2g9N
gtr0oDggwGUBx/4Jk2GXanGJiCdPd5hutwt9w8+dQiBNAP9QIZxdRU15xPcKrfM/jWjB7HmS4WPc
SFE/3WoaLPZXv65oB6sumu60EQKxnQRDIG8KKfpEdHhvbx3JKrUv+wZmN33z/nUoQ3vc536o+szz
JdrfSvWkTWXo0R7nQxiUWr2sQXCS6ZgoAIIQ8AfiE1lnzuRRkeqrgNyg5sDMJqsaqbg+7OGy6pcH
nVQXpGTGer5wM2XWE7gUkYE9i69AWGG380zRB+88RgG5UoAcav4+ATMt8qxNg2Bl8X5KixWhdx8r
1g/ha+sizFMp/6M4bKKUBId6n/o8VCkIVxtDmxdTertIwHYFoA7fF24rhiGW97Slg8rA2VYSH67a
0xoJ96VE11G1YwZxg9t0PodtEk4fJGEIiZYGTdve7budEduOdLb2KYn4OSjZOQ7kkCBrrOl/IcU9
Ryt14tuxxXDyfjdedo/cpzEMiVPNk7kZOt0evQ/cgqgVfJWlIYX5Kmo71SAEr0Ps+z/fbniXIAZm
AamKfQyMpkwNGklyX0eWcBOz8GgjB5Cu4mi28Bddku2oa7rWoqMLS6+wBcCyUCdMUwj271fcSWbF
ViGfQaJOD3Uxp1SKtMsG3s2YtWIKHNTdfkxcltYkp6kUf0HOAfeeTJJVSHXxUqXqQa0P273JGxsk
gnprsayYmlzt9lqOHVMI2UygQ5l9KBbgq27b/CxDLseit0iAiNXpH72wTToTr74wfUo+40V/1QG5
PwlFnF39wCagOYm5j4rmTui8XDgEmCzrH4RLv70vwd8gSZKtgLmdt7UJKxE1t1dIh6FwwNIpaWw1
Hh7k3CUQzy4VF+S3Oz7IuMoBgNddbUTlKgQv2NwBnhqyiXzIGRIwkKLvfz4rojwxUXw6QSb5Xldz
GuSX4YYixJDaG7ESUUoJLPM+NoDnqePD//sj599/GoXqIlSPpvlJ/uj+t7Qavv+97FeTGiwbjcBA
c7XWGXT2Jea3NVJRCXFeEqF8YUpYxne0Zq53sGZZK+RdqrHboTRq5j9NnTIcgIXSuAXVNlV3UfE/
tZhbC7v/faJLo1otMUk7Wo4k2/XPPhbYiNHcypTW/a/D4v8iwpsUNWuqTOpIp83+exL8L5g+FFXY
7z9lYWZfU4jz+LGRzjfb+7jpTvtBZ7rexKBuauWWnvP6Ym8zNbD3VxH+5mGvFQ94ym7QvIxhi6gp
nb3gOu23wwihyFqOacWyIHTwbda+QnQz/0zsILO3fVTV1GcipmbtjU7pVcUOjlfitvUJcjy6FzYT
PwErSF74QStlHUiZePKWOnjH4rBuM5xxGGp3nzYYzIZB6dRhxx0vdEaW91QnRrrYXgOtkvFic1zk
kxZUhAo7gH6050rUDMK5rzqGjpEAtZ55AKkOYtkHpLz5DW4NtYOqMWIzeAbLfcWRWz7hKZf2IZB+
WBMf11VS3RUxlM1hiKyPfyPTXkKK8MVE+TKCc0R227l6TvMsW+3ALNPxWJMfluN8aEVGyFpIKN4P
R20ATMRWWa4m26954i64jnExKwzd/rFaqSZGDBhvgVaTNBnfCCAsdF4OyVHb6pJYL6yUoiMVj/JR
szkSEVGB5huJjZvjKovyqc2yX3hKmhfUrNuJ5uLO07WThi92p7smNODlGiyfdJhNypZe9YR4PvdU
vt8Zh3VouhKSIOFCuimnWSzPWN/0x5ui/MnkPFOur+UGqbdW72w/a67FQN9eeuFM7nHLcrB6tE+i
3jkAYETUKeETv1JEg5c3eNCAoCkq5Oa4GSCfPxqjAtX7q60DvSsnFIwecrWBS70PE2qDN7Q0glBu
DrSVU3xD2HDIVd/opJq5DXZiM5u/LUI5i4hL+LQc0lHg1VW44bBdpbINw3Tcr/W+0nLdmPiY4FST
eOPexQ7TMkNO0qCRYoCGzJbWgW5uxW0sJiQ/dHudoqsGlrZf6LtM4Ur62Hhs7SVxW8j1d1DvVBYt
RqDA1tL08l/9FjhAcsVKySXRCCJc7wSV9vgyGS7Pyy58DalOTFUib4hpxofn6b6iDtjMA9qtbujd
zo0WSE+01nmTKHZCh+OLKnbe9mK04JG9DhxhHsfW4wcBS+4WVNFSz9giZh0lgZRH1BJPMmTQEH7j
Yaqch63w1caYzW4AaOtqKSO4E42p2WLOfv4QZObWbo1R/4JYbh4FS1LF0gtBDL5nNkN+1f6qzvrP
YKe1c9m+3gFaeauqfWgBgKQ9QOrGuruxgUJOd8H3S0Zr8tY24oK7uty2sfohnrM1X4W0AiMU5vVG
Yp6AXKrReKsGea3ZYCi53lmjx8CH/6wDESEoaXVI3PCLxIQzaYkF8hJncrWPVffVNL64iwDT1aFt
OVJgb/ngbSJor9LHLXYxbA9AByhDF+ejLFJn6u505KUTHqldNh/Ox5Q3rsfUVdOZhNF8WWOu3bo4
w5yAxy1YMsGij1Xi0DGE2w/luXlyrQZjQaCMrMLkog78jR1xGelo9P/248iG+L6WLpWsPqWymR+Y
y6IbfY7qTEYtCKombz3IaVa6dlyvMsoKgdjWdgQDgxKBCAxUCeup8LyvG2ytwjp2ZqimKve2PJJg
T2C8CvpQrGIoc0J/7bxppKxl3FCP7mByeCF/o+HVEX/4eIvUNvBfVW6aNxx7if+5AvFkU3B/5w9H
eM06Qu7ESmJ9fN5Ikdr0tv8QUCi23uQwNAtZrzgixVcqXFAc+N89ow5I3m1alWMd//HOP7yNWWI/
P6eZIRCMELRHccu8bvQULA1MbJlMRh/GTgVFl0xsbFrbb9XJ8p6ZCsSvnpH3aExQxb0YMMTZUI+x
6Ihi2dJtGAQ/b/VxJNBEw/3aDxeG14gY4IRWDtlO/kfa/+bHZZG5FVNsSDGe15+MuNRo2z8yDnzT
kMm9+He+lDUz2acGSO2AiiXTq6j57XhiPgkGnWD3Cx+jX9CLjX2ksAJdvKDnefhPpn3T5+LM+n6O
C0sm6pd3Wi+c6HimIPNSTohRyinDKGCnAf25UlEbkZRAg3P8cRs7rw1rI71Jhy5+27F9GJbR8IoI
quXQmZ+K/VSmvSyl29Hn+5M1lQVRzW+dfObQhyqPxfDJezNfgiymB50PULZMUawUtIygs5bJ9UjT
+9bxp8rpFhkX+A4d/9tvr6stZcpHBGDnEEIKM9NpOD7SxTe8EyHhF6FGohhj/SkEHjt4WHXnFd5N
cIkI8NzZSwWkDV8B1vTQaqqfLOUWH3fx2gRc3drEiJ7yMasFEMGwiuOlIDqJADKHM4kEj7X+Plf6
8T3084qbmqno2cfrcGbyLy8IR0YKcbZ6LtPre/KwLM/vF1UyD7+QBQuZQREkg2Ye0gbZ0uShyMiL
42+0k1BxAftm6MttfxMDS8leTuCyNj8rx0eJFS0IgdWhROXsuoMGcr0OC1f0F+Kxtp6gTWK43/fk
Z8xdbEWEsTfANwAUb1HomR5A0Q+/j9fnkd7tf7RNB247Vwg23pYkAkk2RUEbPIXPrx9j5xk1exRE
DHiDmFnQiw/ZDZ6n4tV6JRB2blVGPw3qh5wrBGKSqxXnhMek76Zg1r3nOYnySNa+kpqVnYHYYmF/
k0avW2bHV8QId7OsGeuseh3IJjq5iJLSwK2Oudc47ovjUwJ0gnlnrvy43qB/l0xRdZvx+VN2Thgy
o2LBglQn61jZYa1iCU0oYyZLUBxIdYXB0I2wBv1815gNzm5Aq+l3YAkY9whH9fys+dO/hrhB2KTV
DdEfVjRWdKKP9LdPeT/CZqoS5qcZY+tymyOlaleep+vpN0wGqFCcWgmnNFTZxGLwq3Twow7rpI+T
5/dwr8z4iIu7kiXB357WxwL1S1ePkokhlPVDsuMtFSgQyF/ESwpxMWHGtMZMfr03X0LA4OlGnKUB
C0r9aOR17s7o5zPu1iVS8LFbAAg8G18XaIWLs3ITFoR6127CHTbxeCmwqiro6AutixtOeXsjaSGa
hE0sehFiZzHA7XLaxv1LyT3vdNGMCCWg4Veiib6MV8zPP6EIjVl7hD8+3hNXRfSWeoUZFi0iIUI7
uj68+T68/KWErDsLTP9cpu3EzF4NOcHSB41yF6/zIU92nXS3TWiITaKvIZcTok+I0JgIklLAV2Rr
BriAk73ON5bPSA2oioNKVdZtoq8SvXtZhP/I3F1ydPvXX1Kwx3hr/datHuco6P/6dlQx1/5gToBk
c3dRYnHgt4LGmmMcQXUbIWVBQvuDdZ1XFuf+P3+glpYJ/fShtOnWML9E5254epRDJQwN86aZ9+W0
6JKiGTOhr+KX47MOfienrkB12lKeVUOuGO2yyQCksj++EZnoQHcvXOBN51E4xIRREt341j/3f1fQ
TP8zAkOqawvS8RjX5CrJjUZmv228YgBPWib+Ky/N93FphGWHeuYN0jhhvAA5drVndvz5F627mqO/
/pvnuxzJF2g2vrxFyJXDBn/n2gUA+VXHv/g+6gInEkmvYbSojo3iEaLDCdYrzoQme2idif3MH2R0
wUuH/sgOm4bERu9w+EB4YFAt3TNZ0oZ94PPy4CX/92xmJtPs8hS6n9ckNOp/Q09rXc1+KCO91g76
YDVMCTQ9NFFPw92IeO/LKUCdzGI666XZDgWgdYQZtismK1CEUKnpcTx9sZJb/eODpScwKArUxtmz
n59EjYjAQIo97ffK1yoLYiGK3fA6uUi45gDoBlRQeNakh+ceGERJaP80B4F1UEPLUB6GxZXu3fIE
tnqUveQ3PW92GRKGiGLe/VYxMtrdqK+xsXWFaEmmLxmbDJAlY08dwfFhTvpd2gJI1sLrY5hkXPIa
Emg9MWgXT21fdbfdeS1NX+VkMpqTqfkPAcoUm/TNPbAfUTO7ZY4YoaKREUCjO9mVhPw8msR8Xjyn
ugXIPLRv4I0avdFmQv93q26DmArbezzCCnmaueo57JLUVSKJ+0H8GJtpMjp4golvdT04KYlYn+sC
qzmeYYfzFS/r51HvCHgMQdF3gTfUcEQ4vQM2tv3Vqcf+pztfhSfAjYxhiJuWBdD79VqnkpwbcqFF
MI2O7p9uID6qyDbUlctnIOlcZ2RjSqvdu0D28qFSjNvzJLFKqGHbFSxtxJQWnZ8y4WGW6Tt6DP0J
2s5xNfPJXJ6fCxS80Li84x8n4xXLvzq3+qGa9sVKzLuZAUZbGnoWK3IYD3rZKQAaZfVIodmIlG7w
n1mFDM8yjCzplzlPQ7JvQxY1/2UrTcPnxBzx+DgPMelPcFbCfu54GIUVxLJAtwo9CLCYnNwoF1Ln
iT7649DIgISO9b8X3GhJUb7Rf3qIBTj5EEvZNWtp4JFolmGSyNW84+vO8C7o2PD4erCymF/7uM56
QWzSFGVElIZIqVBWeTA5bQb82Wn2Nr29SLLWBIy+afbaSFh+KukHbIlS2qT4XlWbl0dspxs3SK1G
NqxmMO/QWRmL4zNpwxEcm+akrYM8okFpIcOjmAjNPiIsLHO3Te8YgBZ7N5kj7WCsnY/atxc94gJb
Q4BOexc+lC1Fc3hBcUwoYtoy/iyOtJ32Zsp/EpHrFlKZ/Fts7a3sgaCnyP4YKkWqRJaPl3KllXFT
AWDlVrpZ158ZArpPGQSyZW2d2zltTPs89pGkpUuxDTZIK85HxZ8l5unWAnfnlHsIehzkdLBn1jdb
Lurv17QYkGMdfan0OqcyC67M1nIwNXYHorTkiODMwb1QDKmkydexQWS5cEm1M5VDgPnLN4dF+BAB
G8yvf/ffc4bnwQOCvWGZvrQPARS4dfHQLsQol372Les7fcOApdGdn7/RYApWC7UnMzIfCIcivryl
Fw/fI7xNDGcIqZGj+c1ftCUe5MLEPgjBRuIOvwtrowSidKmt/bhN0BJ1OBUMEvDgt7i3SLb6rhnR
we7WBTmLWriaUX3KxF78YV+R4QhJsqVWKQ/X2P/sLjnjtMGGZhiv/RT0TwjlC9UYJUmy13dIW8Xf
47kYO9TLyz14mKzDsZa04mOPHW/97mQD5xmMM3X7/MU8mP16R8l02D1QJAFjuntBmKlfRUVeiUqT
4xFQDsUW+PSu+f8qLJAZalUPYdVfRxDeB6H9HK1FiZLfa/5Ra+0b+mlDAuCietmueHiNCciGt3uD
70bHz6fBDdgG2fX9aN+M0SzZOo26BF+zXYWjAlKQKMsc/rqJF0CuWLfMQ1rTIqa5iLQ1gkbM0zQP
L0bK98vrpdn+eul1U5IXZOlbCnvgOzZ1Mro5vJ1N0ohK3bfmb+ecHiX15r1xKTkvNfa5XcoGLlTi
TfgHeKD9KLHPdIa6ydX5ovZpO56Sjh4YJhoInx4XzEFrEqeXdripUwzs9eJWd2m2reVD1XRHvl8V
iHNcl3bb8ksFZj7fHUkCF78sEyVps/RJL08GdDb+MtpVRPmF+ULRQhpw6F/vVkt4FO7wmpLiDEC5
lh1tDwG8etCYl2oUaifh+Bi8Dy80vUcuK2S3K43yvmS63yoGuYPDRvgsnY0kSIW40OsSuUmgvEUN
pgKuLxZzk4sKj5RNg3skE1ojHiBuQDFJNZUQjb8+z86ueRspOfgiTHQsNmQhUI/lW4z7I/6/ntUl
bMLE6A4iiyFZjPOvtFb+e33TfWP/cS/2oAkmYTXQx7KLojWscjTmJs8clnPlcw6Ol+PgEO9NQSP0
dxbknb1x+tHw829QU+2AfVamXTFAffUpuLUQ3h8wgLhEz4UXYvMPkEf0nI7DspOVoaQpylngS1by
GrlMVlLFM09C6buKd0QFLx36nmX8fYflQBicBCKfBO5YVAWtPiwKWaT0P0SWvQ3mzEcuPYOBw0Xx
Axw78TXqdpl1N0VNw1i782navDRKFQrahnaM5wnJjVd7uULn80FoUVzaGrAugEk0hW8HDqATjLjc
52ZNh7zjr/88NPxnJqWjGBidt/Qu6RmUphbmdfcZctTuTbmxOxRteh1jDBZxpd/6awh4xH5JEsv5
0miDU4wo5B1bd8Pr3YXVWDhVGtox5VFIz6dAPIYVczWtlckw283cBUEHoI78c3yG0ryzHaTOxef3
QoftwnMY4EGpZYTb9Kmdsi01sJfOgnZWdxCkd/Fb3+j7nwNfkt1SVc8BZc0Ia4DMQiS7B+DCZeHV
j0VL+uV28bKYGP98LI5tB99Fy+9WbWzqrnOR9GcGzlKpILYdySt6iJDkxPZsd2nXP0f3C6Xab3i2
QdcrtDd4H7uiQqrVaWn5GNhCLUc6pWY19vA72JQh+eWtZTq8r07Wd7WhFeWGJasjzClyvV3MaXNA
+Cw508kaqkmOZ5dtdZPMAMUOFo20r8kQ/EOi+WGvHwbsdXHmnWzBRVzuHKF6QTZ7xdyqNJ7AQIfP
A50bvng3ZqXlhM+aj6iKzQGdnAq38ZODpz5uBqB62BUydeq+nW7A4TCJ27quCYQhTaygRGmZ4fnE
cdQM1ZC/XEJdHJKd1WQ+RD/U7StE6aAkPliF+LP4WTSQzWJ8pQkT7r5OjUvrpwEhVwwoMvH0JzIy
d9Rm+injaqf1XrMvKkRFzPVeaauuuiL0nbkAQp47MOk7heuRsFz89JNKmTeMwhw5gy4HLCR3EgHF
AWgdDblZZtWXkJ0I6mva2ZJjum2J+hX92MctKGOQushmXMxHe4F1Ftlw0oMZXzS+tJ4PSdtVavQ3
vY4OVTN/yzVr1nxhCT4TA/PuK5KekXW7WZUFeTWkJ9/3eCsh41Usw6EHl9axJ9sB9LquiaSFibwO
YuBwdbXBwfmD/jLrhxujhLk4aHswvKP9PauBBgCe9dp30rMDpr2ycq7JFVSxukCiL2FMqERjhnCR
JUQotjUy/V+MF2ri3u0MEJUVeeKYpYqwgTmkC75zN3juAju8CCjhpahhBxAcxJAaF91zpxpkFAgx
QrEvLVXUuaan6cYnSvAr5LrJIYfkycD4W1DRrAH8LOAePBQ3EIFNqYy3vBRM0Eg7LyEAQ6Uvv6Rr
SA7qjfrT04a68CRwlNg8fhYZqjqxZnrf/fKCENAjxsdvl+uMHUYH/joQW1lZlcO+weuJyv1MlRu3
VJ1aZa64eDObYt8HhrD/l5E+EaQ5YJY+ZIKuBf05LgjIV9NdHVfbLEIxgmTx31mwcS3fffagdp0r
xZQS9CpTEb5Y3jhbSkpIczlsDIIhORPwb5kUWqG1TbZXIVBenMkh0qdPhN9YhIrFf+xLKik3anze
Mvr6IF4b7fi7WU5egov3XO3BHrCeJWuezho7W7alHytIPdc5nQDXPWje9lZYfOktaSquekHnj0PE
SdSVV4h+VK64J0O2N5e5V4olPzQYWy4ndQF9eoSpZUzEf2Ws0q1lSq8iH4VxFGyt537dfKvcjWjh
eLoIJoy9HR9sDsxpdASeoSERZFoaCOrZoRPQIsxPozzIHngmL54dTaP4x2MXVIf3bfZEKoY5dO1o
7eLZFiYiljoOhJwr16RmuI9ZRx0ZvO4854//r+mYKm/Dqw4oZ8KvFOP8iaBHCEQ9gzjaUrJd/Rk2
bf5mrgn7R2yI2sXvJaXT+Kn9nQrMMnB69DcZxcXDI86aCnxf5CMwlR47zZJQyYAyaG58qdLz8dKu
E/j4HhzDbsKFKV3ItqebzfJ5PKnzcwGi6Jrv1md6/+7tBR8XExkQ2uCSvjegjyetcZnfOJGRPFuJ
3uZJctmXGrNup8sdlEqeCScMp/u2yFmvs8jR7aoWAdVdjMJO+wQx7idngDwAMH5yF/h8wVCDkLGe
xMZBYjCVbkdbMWbHfExx3fRSa6g4qsXHOzvxHXhA4CTyjHxaWNlcSm4diOfxzMEf1EnmKOpXMKvN
UKVNVVAlN0vZAZ6L8acNRerkB1/O38HegSoVSBmDotIP9kEYxj3NDOrwYKrMoI1/weN8WGV16/NM
ZId/kOGweTu3sXm4+uvv8qVGr8HIeDJnhaSzGLHvIt8wBN94+qs+zEiU6SPFdizXt39yCSpnVQ0/
9gKjVzQMcZiL86P1AksNk2zlwGCrZ9by2xmKTdM1EALGbZqiMQHVc20ZI9F5+rUtgJCBhED8d92Q
34XqjCLsl2WRq5ydwvvrAiKsXDSogrDOd5zskl7j70sOnnPyU4Fugsn0dh47ztOBiCfMPfgwkxyd
5KSZWBstOszSE5vxHRb78/2v/8StePBxlUYHKT+7YyIz0p4JB19OAHovXErC3wFeJkyO+Sgr0wdT
7py2we5qLTeboK5Ra02CK/mONzKWfoBJjtyAIYbI0SqtTj0nJqvRz9ecf6NbrTzNNrGX1ISozz6h
3zERuugnRa73UcB6+bMS+cw1SQMUqwDvPyBIffBcVm3PHLS8IsJ8GFlivv5CMxppFRtAQMz5L5j5
S16r17uw1cohZc34HowtyvXqYNTUTNPl/txxM4TMHbcPZmxXIORWx/Ki15D5wdcc6bDz4IEAjPw9
aRVAPQ47WdZqo7Wq11tvhuWYaGqAfv+JunAmA6pwGiXen7Dla943xgqZB9aGtUTqySTf82CoNxxN
ctHtgPWR1Jhr03m+ERMqdx1GD6ipyvUXIBIiMjttIP7+1qPYLBQ/0rSOiLvrEWZgR+8OplDpRr6I
otC/aKdE1Tg54m3WkyDVe9OXriqpFWj0USeFrnxIt7SbnsXHBVAE4w7vzg6f33G9hCPkByzJ7xOp
F7XjOf/EFpfX/Lr4jxh6JwmN45jNtd+6y5+O4IxmfTGo/4oGTiMZvxpeuVFr+2YvhYQ4T9lqaRJ9
H9ylCBPBJC6YlcmUP7srmYa2H/ooVJAsWWNGXfPIA8xVYEoFwTl0xbQ49Fc2zBuLK7c+Ts0dIrnq
ggWefW0GR/Fci8ZfNFmtU/+5hjdXKJI5cD3XD3H1epZmOPWwjitW/Glkjp8qN06yFaYFet67SP09
ZPbkw30foOMkKhrOtswykVkhkrlNc2AqNS2zR33hDFo78pt5AYOV0cc84Z7N+b3JGCSkw9wW/znB
Eb/rLnxI52tdfrfD05V+4TGc7u+t0A4UrYexWQZ5UoK3h57Ag0y7SGxRz4fzv/ZTzBCDC/sxm1rJ
1l7Kod1UtQPE//WhEIaV0V5I2nn/6xEheSI6S7/cQ2gXcu2rNFjXtoBVzLMfEoRTetHnjRaRKsL9
rLSeQyvBLFB8eAFP5/hfE4fZRI3KRNs8WgoUAc2NH26GqM/8783qxnOe7CR75aXCqnvUENMJMk9F
Cv5+xA7sH0CnEEJW/imz3ixNpdorARnhkqMz2I/YmjCDYSlV8k+Jeys81PllPX5CTvoMiDqF0bTb
iV+nx2oHq+gG2HdIacQEenszburlly5xRt00iKd6dtDdI0XU1ur24gnl6irPJN6snGOCiuB+NV2K
K0t1Gkjk2+jimcmgrWC8L1CxHOdEEwCztAL05bNloE2Wn/IekzQ/Le0p1mVt3Y3QQZL6AQfp9QRQ
8IcZJysutszrOfgB0U9UkMcCLpzl4OKli36XMmhZHWq/MFWKF5os9EE0CMzA35xCDDL0YXX4qgen
oD33hSp4dSvN1X5d17Xnd97IVyHLwCeUkpPrIPNOQ38A2xCqYxuza7nUquhq7sgEouo2/lv5O5eI
0yiWhiDjUFXmGx9MYw4c9Zi2COsDzqkPi9LXvrl5Z8IoC02hnq3kRfD2GKV12iIwxUgWx1Z9kKn3
swyo7hot9Cy3uJGFjJPTC+aT1OhX+e8gqPZ1KkNyoiKMr0jNsJTq9u9/Pyc/XR5zw4eCRYmFQ6OV
yNKpYSuMWuT4wqQKwHZzlUg5mVXWsbXrk06+TqwYju73GnTBeyule8fVagH1zCqrIBSVdhA0Q18U
VlByoaAFHv3KcRKr90QfiYsHPMH+x4GWegPzwpvxJDJC7ZfwBArZZrGLpL56b39sAIi6xqFURlHb
qQkNUlGieZ7TEqbgqpVKJGVlKuG3X4ijkI8lJGd6dts440egBFbB8MBRihQa9tea3VbcWgc5k0ab
rfg3VYrd0Qs0qLJz/xahFXNRPUwm+borsvcPxNk25VmGzZdmwLjRD9EvLqjA8ua5BrxhDaKxIp2c
xqUrJRqmHmwkX70gxNC46xdiZyKwmgjrfXRWP13cYZ4LZI7/W80NVdXZPzv1kr6WLoBzNv4Ih4so
qpiuKFcd6MFDrcJq79i7izySq3xfq982GzMaKzIlvwvBHSpUceYZLG0YxLYBx9qjmdxFiPP9Lqeg
wEPcLLc3Xv/ojQkiEh3VtPV48kgUqTdJz7MlBxCtQTbWgroLg70iJ00YEhgHRFDfvYJolXNI5m/1
Q+D2C7zq/2WKXOKUwg8vPr+eBFSarYT86zb+lLKLWsVOxHw4Utj8SoY663aeD5cjARxwNQ/eiu+d
sJRTOICNVbRSWJzOLR7b8mul7b6+DLUm7vpJoWa2X+qub7kZXCZ5+fTjRaDRHmLjZVRH4GUpoU3N
gDvL6NPOkFkZcWZVVSs27o/ezN0TU9leWmIshjpa3de1+LEFvr8Q8+IJW2jhg7KQVVzDB7XzYxAy
RSQKRC13TpifdGXzEnVaOvpAr3zlbg1j3TaM9WgtAwwVZkt8VaBTXWMs8heA42I8A7EBa5XEKHP0
GmoBf1/lgg+umOH/kk+tVZLD5PYo3S+9YIy0x6QRXtQOEgTdpKpPNKkUIStvVo5huRJMYMykOcDo
9JNz7Sj97/fvn7OnD8WgHIRsA0h6KlOTyIjpqfgEPa8rxli8ypJ+SvPaRUrG3JgnV+10GV3ii1uD
KznnCit0SauzC/my8XxXkiqevk9sp+pxnU3uF4e+aWndyCS5tlmGJouOKGoF1wPR7Vmc326q0rBi
gIki/0IqxYatM0YZUgZtj+Sm9D3BUEvmYPN+onsLE0E0fhgDHfnJSd+hgJMc5dz6jun0H1k2ZWf/
RilJxx779gmgqxrxQaG63+1Fga6DsRu2pFcPuUE5RqDId1UEj4f8ZrBCI4jFTI4MCnEgewDyI8uA
T1Ehd9EjxCc/OmWN7Me2DqskDn4qr81uEKNq7NGPuUDsY+UbNLQRZXanq7ENopihPPz6Sfa5YWOu
Y83QyvriZidVPA3Te3jGckoNCqiLDlspGmm5gjuWLxbOoC5Gj1wxoeahpuxmFeAor7CnHh1Cb2sl
SD9zGQv2i+dhHEtLWpXsXzp6ctsTTQOprvBl0BhlG7nffca5w/TOaZEoiS9eMKmtqGtRcOZmX6U7
XtpkJ/DpJwwLGRf6rYkELcDAP2lwv0zP0iRLxwUnE0z2gnKKxx00uLJYaTyWr0Ke42f4haFtfzIG
i5qwSrS/lf6VPDKz156OGzA9ph1TD3Tl+zwMM4ylDLMs9Y4Tm9lMXwAQ/lv0Gk7r5FP6MYg5jX2J
8nIGfDfDcozkUq6xh9vYRd2xscMLDNAz51WFDbEtbWTyrUfF1Cz/fgHnTY8z7b5JXSDQXo3IY96l
ZtDB2vZ6dmC9O9Fb71VWWPQry843b6dKzHXVJsXc49IdrLQFrTUmq8IHzjOUFRJzhazYmxfNvDsK
l7/Oj3zz+kkMtHK27D2RPDWKr02Ni+XgDfXJ07tu0ICeStrPyyQCN1dbkI4rBWUFsSzY5qRUKcLG
iHFtG8NACMj1ODbcWQhTMx63azC2Snq5mSfZ12sdzmTdMiEdBQZ/olRErPhSv4XNRVG/ywWBKWJD
qhbABVY8HQX8dsLgSKTf8EDa14Pzrgzmo3VoXWGYAEy+aEjtcoFiPfihHIDz/2taMcxQsgpoqcYe
INobKg9p5Iuua3gE3uwvnLMTeOYmKrfeL1CR0QKrljK4KYIsuNciDcsdvyDUCyfYNsRzAURf5Ttj
uDFYafauq5HOxU5brp3J+/mQ/vos2EDtadThNzY7Lzi9F4BPb6WBhdfccDZEu34LaiLGH7tNhy+Z
qSOd+HNNBYxTa4V2QZESQI+vWPDJuypQMlCwNauFcf6vdNur0DKSFGaoyI/uBuAi0xyd7IZr6dAb
vCAKpxX31rsoKvuSSGg/wlCV/ESHi6dzScoK/iq89NaGxvmOVmvZapwCAfObHbLOu5CpVnlP7Ha4
bDDri/T4/Es2QLLLjT8QtSjtwHdJ/zh7u6eba69Hxb0Z1gj09iCmznMcmTGRpdy+kac8wk2WcSTM
C5uPM8NCuVFanIpRlAhYsVgg05bL7fJo7Xl9jctVGEGFo4BjJjoqZwaqJ+Mvg7RXg7saVkN5X4Lw
TvGYJhP9LqY5msXhGM0BuuwkTOL1Z+oysA7hOTcziYc8LyFLPA0kqEhrQVrBcJEqiMPDZ8JgwtDo
j/7eeH28bDW7ss9ey6VRNZqfhvzzffHk2cKqLAtv6fd3vwDDYkHXmKjAHgAJrnXNv5a6xecfrqIz
XQ+drcQ9oQIPZl60RO8xAAIre1g5yeKymdK31CYzVcG1e4AUpaSvB2rQdd6ZDJrarr4eJIjXwQGI
byoAus+p6JnRUtrvM4v570k3gFxF8XW7enLetUsqNQ2FS0SWsu9+xk54aNhcT9SBvkG1ekFuL0D5
BJPGYlEUTwWqnSKKOS3iSp/2+7d+QIDvaUspeOSiBzR9paNeIUIB6jarGn3C5V7kO3FVPHVeSNmg
VlbjQYYgrqAE/OMhaM0vOEXBUrepTH/h8Mjg4RD/2Zq5fBLGw9vua9CUMSe196+AKMzVWtPQC+bp
lmJF6NNSZaaWas7Xl60MyTqV8JFf3kkw5bQlTY1H2NOpYTtkWzGqxij40N3zA9HJZacuFUjfMjxt
dpnPUDg/d1U0FRB4kS3Y/NWfxqPNs1zoYgm9aM7m8MsNV6p/9Ek/dvj8PmfEFwMSQw7VPbBbWyyy
wpXzHwmjVFAFU22mEJ5MlF7i/H6aKkYWpgk0Jlo6WtR8Vek+jCPmRdEPA4YYdeNG8f91pDtbVk+d
Cb5v7nubiac4FAbp0U/fjZaS5LvV8J4iVitr7lBgSG/jqVsKDmxCPWftQ7lhvRiOMr5TUMmxBUV/
TIpmKg0RFJIIGQCDzDSndrNsZoc3+g1DNWNApSl4VCIJtNoq8HaRSR8rhOeYRWxWkCCcqzMl9mJ+
vPPboLvf77LWeEeTX9w8oMWZPTlAqkYGC2u1zecu/r/2UhdF4r9YU7JA0DTlWY9uJKSAw1hrT86S
7i4K4PqQOJKsFcfFSdZFgeNllRIhl8uXw28ocrYRAk1oVJxQ6z773a6tqs6W0etq0esx+l9UDG16
MpUyVMDXjPB5INYoNQJlJvg4U5KnI9fzFrOdzZETrNjpR4UbBkl3gsdCx6EZt6skI8+/tIFnClJu
gM6iegQBzYdvgcaEoeiGWzCIKt9Mm1ruy7ZDxdr6dZCP86PG3MkgOHoeKqfKDQM4D9HfNGlOocKa
XfrXx268LrU3UDod5Wv/duOcwdLXpUFsY2mv7qKpd1hhxSdGQ1HFHyNp5+f1y5czvK6tzbyMeXev
P9B7Ho0BAUT2uUX9g+A2k3UD7FcDfB4K0h9lK7ads1BkiE0imoFYHtKoAovrn0/QJm7vBOzjg8xb
FlSxet7hBtiv43rhOpUgW0kqFzk5xR+t6eQTSkP9vttOkxtEiUmVy9aQUOGutgI2RuAQSjo+fVwH
VXPoYbzaUjlHliCDdgdGXRVRlfKhGHTqUwONNPJsyrORf530wfCSCdv2z/1AjkgLjDEXWOPuf1T2
+R3XpQ4g+HMHJe0HXJ8kvCtSBQZpgtaRSvajNNnQOTnuQXpd4k72D35DKWkHzapaHfk/5Z5rmQz5
BUcdTIAISvEMlPQZdEVP6xVXa7r0XJaVGPVFrtvlbyy8Geov46WdNhrfqNelENM1N1bZuShmGVK1
hCymg1NfEb4H9WonYugcigC8+7VXuIL3VPZhfF3pE2TG22RyA/buROtM8Ii5eDtJ78aWwi5Kb9Zf
BxU2y1MQX+1JmpszVaS8zDLewihOCxqBPECI1SiraHuu9aXGOJilTuVQI90DmZgONs2ddszGpmWd
vUGajkosaU5HukZlJGORu0+5uRgTAOo3frrIsuGn0qgnEKrHSybCDD65ShR9P3lRFiAWekEYHXT4
kMubP0RqDEi5q9rCuBC4TcAAKq6rerUkL8nfQ/5FsTn/YJZQPTX9Gdv9OJdvzZ714LLEuvQ4xCpA
HSR3nrFw7sTHv1g9dbetllSv6slbbNBP9+PAuTcztwYx0+0QIeWxhZetvDdFF2zzdkmEbhGFGaoK
bewkpJEXR17mFV127MBkO7JQXhOExCtI/uRCfrJ3IM+nODHkO54vPPLPm9H0uIlehdNOYK6nk0pl
8vi9MhyX5jZ3tIkbso7SkQ6BD0X7pwbd3Yiz0hQOK+Mm3DmcbA7E89noobssE2Yiy3HqvpDJyfe3
UWzLcEJSfVf5DfivYcRNrcUo/h6G/z9MyRdSlbndcLc2B5Qw3VS5f8VhGm6fJehQ9T1K45VmYo4b
gXUuIlpupg/pkWU9McHIya6hC8pJmWslP8X6jcJp7+X+RS/6K3ikNIbxJqmKq0C8UvGSx8kP0iS4
1dm5HEAIoK2e0CCaFoW/6ONrkiICCO+gs1t/V7j8Ykz3ZMcNRxfyXu8sMjfKA0iXUdF5RvwH2A/B
5E+V9F0R/xaRGQ6Ueh7cuKh7DYbsUE/GYymnRtB8Hd2AegTzO9gV5kt7+9dmIXakuQoYQMTlTZWZ
qaPEe4nR7CxNPZtJNFvooEAlG0cblV9hkU6dbS1p2+avne6NOsOUK+TDkDOo3Y56QwR1e5QRogWS
YeQBp0ri4E/6oZC0dEYsAdDnA0zggnsxPfujTR8eFOGrA34qyyYzoZbFfz/LEOKbDEZeWEWBJXbf
cPhtFMOchIJsd6NZqrs78g9ZBr7rhbfk35zCl4j37ShIntC+8CHVr0u/9vD3z0Z+hNi5VVltm2s/
Sjz8wfeQAV7M4tw1yBlD10I0TdfrRKHdn6pHLbMFglVhY6OUDb+PYLp2FkxqnjZb13upXBMg9IbT
4LX+0cam37TXK8SvKNdmzaNzqQhOCiYMdwxJ438ZPcRgFlR4lZPm3GKwhARJRhPnEqCvxbl8nJ7O
sMTRTBgv/BB5e3KtFU4i2SUxB69rFBGjWy03zuJoQ4y8rvG/V+O4KJooF5Fy6usqiWiRpZowvqDI
u1+UT44pb+Q5ynEPSUN5XG37c42A6HHZfltSmhrGxIGvcv+EwHOhYdvgLz57idq8jpn1eqZQML9W
+MR1sJTluzXzpCiJyxzUHMgFoa2qFysP1zX+e8+PniWgjwj52R0/DD0jyoMJ5PwJMP9wGns87Dmh
RVUIMl8X6U+4ltC08ZJm8tiBqnql10uamGEBLWm6zheN01eDK7MRFu6DZMo6P2i6oTwwIPls8ljP
1sAvd5tqNsrpzngnhQdD2DXatyZwb3KXM7VVZlZj7MyNUCcK+7hgRbd7NmvhoQnOrGOYtAeUjQ55
mVTfV+iPRlUmi+7qXCh0gG6drLQbPnf1YfVFbUaJC0mIo8grbY1YZtrVWRnsqrKidjfQvQN3ZH8Q
3o7kEmVrzy/yd64mC6gYaAjsxiaS5ik+YSEr7T93xhCVNJYxjaI+x0C4ksZb+soyT1Rf2GenvVHC
E5ml7VVRkE5SuKyBOBFQe/hSQw23uV6CQ5jWmfyWdVcKGNCl16zXHb4SbRy1GTnz6OMig2Uif6gp
To2/B+pQQJBHuDKhxSrexfJ4gfniM2m7fc1mQe5CTlxS7Mn0wQT+6+BxqiDdNRv1Au+ktKgn3IDd
MbqbdYg/SWcJfGvL67svLPxWeR6F4gM5EHLyyLZFFevQMbNqImhnVfPrYkla3sL8/4IL0rubm3g+
BaZyZzm2SbEYBXx25ZVP+LOOKhw8ItZTTLSyTx0zbnD0vGpzujhdQe0C7vEMPI0iz5my1dB/XQQt
WeIr5nst1jXnNbfid2b8ZPFZ1tBhkvgE18DIhEgwhZrwXj8ECZgy7qhEnijq4uOvEfo9AZ3LdbZ/
WHMVu8/cT2dhHSWkLg2jcRqSImaj0iUgIvoaDEMIcAMUrBD7gd9drCX0Ao6BEEu4ct7G50f5D182
qEc60AoIgOnYMEaqIxKNjzUv8nrtPxbfs7XxiygNzyoUyRjjvp2dBdwIK0zjFPnJSJ68IG5M70H3
F+K37Ynd8DYImSZBHiwKL8v/MAz/IoeVLR8tZh8OwoXCf7uYZClmZwd3rS5pS0z/AatpjbSCL+Rp
DBdyMuoo9DYdrEQEebtjRln1TQxwtB8hMudMQWRjxcIXwdkk9t6RUAvfe06qnGLVG8UvH1SAbfcO
/QBzUgBQSMahkoxNakcUsxeG1AydmZZbnuxBva/w8HkPhlhWQXMdFEZPiclgVIxnHrPEZkUjpkPl
dVIkeH1sKGavtjU0MlKGAYvhL2+J58yN5m81ijBfAgT5Coka9vZ0dfPe1o4I5ifQBDGx55zctqbd
+gy+9b+JaQ4rGh54CIOG/+aBAy2qdpkZL1DLzcutmV/0J72oOh6tIaop5qECsKmJ3ZCOTnCkmFU9
OStWHv1KtZ8BxGikwn/efMeFumCsCZTwtK8XIGbaZDHVty/omslBtt4RUKreTekzteIek9S9vEFO
9pkn+cjvETnAYspDw6i1tXl5MgpocXACZMoCRfRA1AJlpXmjod5K5rsOsRSZW1IqwCh/BNNUESFX
KLcGKkENmO4Yq5SEmZYtyzKA8zUcJhVqDLFRu4pz8pedqKWbTD87kwX/HfOuJGy6iylukAylUe+4
5opVVc7F/i29pAIQ79wasDyf6tnrRECdhRP/Bnr8LKOfqfm+uloC7WuW30UmMVMaAC6OsBRE/0Of
aisuv3Dc23gvqjZjyVr4SC41TBV7fDtE/UL+46GUlnvX6NAv6AStoNIYlHTk7T578A5Tud95onWE
Fpu3f56u8bO/Ux3IUErWl8DDuYdNInlI6WA1oop6mInH+ujLDZEal9ezG8pZ9xUzhH1SDmLbwrRb
dLnfPe/VFsQZNa5/I5yFP6fD08AyE/BjbXRxjvvXRPEVK6KUvXxi6er48gln9vqTJI9Xl1u108xB
NwYaZSs6UPGXhTZEBVN8zv4otROXN5p0115tZ1pDrz+fu9R0G+uEa4mBr99WqSxDDhtECKE1pYsy
aWmBMoAl/mBMBG7slyiokjlaLQjz8ARzxyW3BVPjGU95pwLBhWDifSrykEEYkC79t15NOPmfUPTO
54F9srHpscfmo17FC8tZbEsMGQz7uaXvCiVMXrGT604EwijyPROL0X35QQeDLpK0sfssvCkfI0iC
TCA/Ut97eY5Vu69x+UwHCDAMLfdcUv9GbwBzyTFtvxfMtgY493Fw0xWrsSBhJRD/F8c9C5qAkr4a
fMMDIbdIHq6s60a7ffbwxZZG0Nhf2C/mrSdutfI5VMFJpDXOsk5Yds6iEUx1rONKHM8uLYc5r61G
v4U+p6LCp73H5wICNmulsisXRPfmjz5J8hTngcwRdFTbvmQToziXoi4A5PbR71wMSRePf1WIDKrn
fkDKcJ+rn+fnsgh5A1MD2/8b0NlLmRDF2CR7zRwZWEu4W6F1cpKBS0aMrz+L+j2YVnEerGwjTww/
fenA49AsGPgYrpYppWrgu9Akyat9p9ngtPlQs+5slLOk+8utmFJxsRPnhGq6XaX7f54ELJDuny+o
jDqf4Uvdbq1krYYeRb3VTBlZkMBEKkbksHHquNSheUPJ+UIfL4zGyawlgbm3P0bX4+OjmNwJ+xtk
hb1I3luvRb0QgYE/0QTeKV8iJzysMGi+lDN0nfXPZl6mAAqiDxr6yzVsY3oFQsxe1TXF6pzJSfc1
g+e1ilFi18OxEO/UfcdTsLTWAgNK3QQ6Sgf+wgIh84kVqv8J71OxvbYvZ6eru7Ojehc1v2tBWonf
VNFbUqJvxNpg/G8dx2yA4Pncv+WyoYKaCjyR/9VpDJqqMafY7OvYafWlOYnTJiA086oUul7qLsEg
ozikjj79dF37Zg8s/3z5qC0kuFesbKxfiA3iL0gJg/wmoLd/lYzKHwWVgJPtP6b5CsUJvARef0hk
m1CSXq66Deh/6+g9G1wEWxO0ddqFi/KiH9/5yIqac12+tc8KELUmV6SSCuB0B777BEjQPQpQOAfH
5dg9toQ5p157R74b2aof3UudLeGVjNt5Jsnk1QLVuLENN237DiioyVCN+OrzFYF9HNl8k49OGcEU
ro+6r9eoqPKLeA/tWfCwmAYROvjuJJjnQBrgxXFW32V20noxu7V6FPYnQpQ7TY4pizJevesb5Zi8
qn0ZL4nnf2TMvKzgDoCwQ0CChaM90e7tlTL7N1oWDT3peD2+Ea1qYpXu26Tvu9w33LiUHoPUVd3n
6QmH3TzVhrrhVrxodySMdR+p7SHA6IMEObVmH4PTBG8yId5w1yVlIM2mAPpA6wyBd5OU6us5bMRl
X2tHruooS4ILNpySyeeGP49LvOU8HQSMU1m6kFK0W9BV7TLqMQ0CWYa3npJJ2dMYcTj+fL5TVUhq
HIz7boSDAoAl9sG15duSg5o2/3yanQmL1mT7GC0tEZqX+eGs0gPZEDTqOvQZdRtDDoWeAACPQdLQ
lXPOwPkQkmNA/D+oLsfiiSCBVzryURla/1LZjadYG8nzsz2Ls9/dzPXxGUsssLQxB+DkTULVb6b5
nlsVYib8aHswNs78NPIYFcwkdTdae/dKsNmLu52MNhLPbL13Dj4xag3tvYl9nkKz5Q5Ch4eCQgam
AiTrxQX0IcD7lYTWPdC5qKxY+iISaNiCST2w0HbY0hqGBxDMyafSXu3clrpnpy0W1o4W6v/InoZD
87b/OApwduoQDgPS0EG6EnHvx+WaesBrs188fLTRQpbCQJgGg9uMDjDx4TFzHXox0VJAnq1Ecc5i
fRC6LVOD+eJ2Rzx7Bussddfd4Hlb1HI8lUhmKquXMOgEHq+CC+8DkpUCg8+lP0bvrRS7GPe26vE3
pJ6+oQ9oVcaiX6O7Dm/WXJzMdvQwkdRJjz2cUmjFmo3sPqF/hmBENkLdHkpWSN0A00OVoI+8IUhu
7iBU+f5ZzV6dE3fAEuuaxpo6ZZlAlIAmBQyRJ18LF6Veu8cEG4KKToL+4kLl7Ah5F1dGP3V9pNeb
Sla690cDtarBdAoRSlzgM5jhpvuNLOlENJQsTl0/pdEPfX4mEki+FikUUN93ki/TJ5QdgObU8DcQ
TuU6OE2Rh1zwBRWsJgPW3S2JGI+IO6F14Mq6sVt+gD2rzrAAavrp2ikSI5dsIJSlK4VmKzSmVyAT
bgr0y5SBuGzOjR2APvYLlVxBYu8HY8CQY7ZdW4VpwnjhVhuSdhQLSGTn2sT8x/qyBG3eODCsRIn/
9q80qn0WxcG8eNjg/8LCBMnH8sXdhD+pW7RKtopaTb9I5Gw64GGROCZBW34Dt9Dc3xh4LHT3ybex
JGAh7dYfYKN8y8URLkpdDKbOToSADK2FA2++JE7fV2dEq8v0fs2o+XVpLr9Ni5aBvUrt7tpKvyGD
bi7ndl6oqzSJP2tl47slLcahAPGNXYPdoMg3C88lpC200s4afHZlkQceP+1CzvNdS2qKcAu1MLqw
CfYa+PQbPMxC8WTfCa0thkoM2uK22TI1pGXNgSmr0TQsnoJruN+AikzdMgPqwVBIaJ0AtbDZ6LNW
aCLaSOOjx2ivS4Nw6PmyJCHY+WN2Ox+TOfrcWA66FXsjdgFNxkYkS8/Y9Aly28T4EfyZA3m1uEZj
QXxizQkrSS8EmdBa7HAlUbDElX8wF3LQJZKuFLDp/KTCA2ySq6Ghv/6rCfkDhffYBx2LrWd00pcx
kDSdl4q8FiL9JiEDw56ux3HQmMqc0uOALiTkUZSjJp3WUy1KhK/psEVWe9hbkpPpY/JMuO5ioC4I
Ug+6MxGZAJwdWRB7E9pyXo3Gx1Rz1DOJd5282tImCvAn6AkPKR3eFdOrC+4aiF8UbN6oezVcVVhu
7/XFXcO2sEJOv5nWAPVvqt1cUUqKBmIIFzsfvJXHjGMKVrfhOJctZip6v15M1l/7PUMHZbgA75hW
cq5QLwmpGn4fFwSjhTmU7v4uDBnvMzFGYNCZqPkeO4RDSO0HL/gNFydWPn3A4v9rMBlJwDRoGQ/6
GjVItXxk4Q/wSKL2yEqKSFHNkQE+OHNulHMeXNz3XHw3K/TUgn4+8jyC76tGT/QGcjyGEb5k1c4W
BlzNNHGp2iz9lvAbYT0o5MIfTLMd1KdYAPxq96oMhRx2h5G7K6ygGjqsWXdGDAlaSVbchLKH7yxi
HNP4vy4Ude57HGnjldelIjtgFcfhbclnfZOZsiYwUlp1ZDwsP10qmSjQeY9w6ZpouBMXypKQbbSr
FQu6m8pTRIArAkZYxlCE3Mu8Ja/eubt7mF+0vkZ54JfNj3OwJYJoplTa1cWmrxldRFLXEKSsVpKM
hB6hdIA6OZhZz3+O0DOgzFoEfosDgVJkcllkbexub1hc7UGwbSTGnyMB3AAlZmUNlxWdzS61GQT7
QNd3YgfbkIFB7+CXLLbnagjrU5Q3cEoF6K4Mz/GuJCT8dFQZGthE0ob4GTGsUxniMwYFGgchpxDu
LFpm/BZRHxtfxcjOOsb1/xJvwszu8MFEq9s5I6xA6XvMO3pZYPxat68GmW3rKyTvFi6bNEos1gTS
R3WFv+teq8Id2+jJewTdarVbeoOXPB2XGr6fp9Yb2Snt8l/nGcAC2xbelJxZLXqR0tFb3LvWkUmg
yCKuwSsQoTTw3JP9xJ69M673Cm7HwAJbgw7IVIM+TzTZv+BF3xUtMCBOSpckSfYUSWqpwPm8r1Xp
QT8Cew/dIGFxU2bGJMlguW96nTIloPFBBcAapNwNbkjtwEFiy1VdbtOKfDVSsWbDEjp9sa4lLgAj
n3Unaj5JPS8rFKHBIyvS4vbcuOTR/JVlEnOwFcRNLCyWdihis1Hx5F4BBo6K2NaSVV6vQsqY4pUv
WxNGGBYOll/c5qmPVfadQBkdXUi0hP99WfumjPrumlngEWZMVer290WknkjfZYMp9M1gzB0Xa5TZ
YsyOA/2P14iRKGl9EUQ/bV/D4VQ1BT/6RWRLJ74CJnmtlowGHqOZ970Z9gVFzjDSPDDwXgVhLqcr
zjMc79/KSMN547HQRfuvM5QO/0X40EP2Tuc6uf38edzQM0seFcdhEm9sLY+cey0dyOK/BxpMPHfG
8s+UB+dz+Mxl0wCRQ7EPnEhgfWRbC048d6FpiDdjZcvJUP/EMO91ZtjbCFzX7v4RUkPpeA5xuiY8
2akZSMlI43dGHkmdTTMOZcS+qJcG2fbf4r+fLX/dpH8J4OKwieZ+x6zdnI4Sjc4kvOc6TO1YG/ef
48DtRaPqxhJiTaos7S9ff0UgSi1gWjscYWpHw4pOrP1c4rZT79fepqIC8tTVjM4CgPTGbSZOX3ew
Q1dtalJiXYRbvWdxFAMGEHx7o2IqkFxlgIRR8xRrX0wiC0uKbQ5Vn1yVgQUNZPPzBfen9fibZU7K
+pLvFvpTRO1iyWluv+sB/ZHwsdP57meEd5KVx4+MBW/CjuIHq2845Q0RHiibydxnYj1K9dhcTCPa
e0dR5kiwzd56ib/6GqU3Z5WlUfOcQEuyFqLW7YnKanrvEXkx/yMlfWSizOjyJxkL7ig59vb38Img
8HWesJ5XQ7h8E54LkuStyCDac4OAhzvvB5llNbmZCLwsm4zidKU5tRRR0aXyZAHbfDM3Fgm83ZPL
X+iao1E52qR6Y8lnl7J7n8JqnUipHWR41XE2gxMHWOu42h2eVEAzYmR+97S4mbmFiFyEuKDP9nRC
VUOu0Y8a+pwIB0Wji5l7WyaiLb/8vZy+ijI/1cMauo2nV92rtkegO5GW+yuy3rd9HStXgmeQD7iI
FXWRx0BwQll2+CCqpRhfAFGEe6pkRFdKJu4YCc2D+fFWwXZTyVhIO3uvYhNvOuzaD6S1vimpzA5u
rob3DR2hhjkLMMC7E8iZqbO1bq5hroOHU7f/0UJneK+pl4fqBaZBWoJ24bYKThq0Vkltvu4qdYuT
QURfCMJ7jA2vo2VF1fMF3cEYKCIVEJlsCHy8YwaY7wmb3hIwCkIazspMEZND4wFsmaRmkKTqy/ra
VudfOemmV7+fl0qQ5pju5div1HnMHqjMf6iAdFp68q99kQHyFwGy5hhTZkoIZXHb8lUapo3ugEeb
Ji8t2UlhJJouUVVo3D8ed7wpMFrNwglhThUn70fbr+GBCEQujlU1eMdFRL6Y8JsXeiwekMhjhwuV
F1vqt3Op5VFwavxKkEAnnQXWN+aW6sVeGBhEPKJbJSjjm2PkBFGCfde2K/NGLO2gkEbtsB9Ehfsw
VFz8N9TbeisikUem/+RuEJK3plpJcK10mypTc+xzaQZ0WL0h9QFEqTK+ewxvfNyk+Z3w4cqM3BTT
Jp2P49EL3fTdWRl/RJkMR/vXX1IEEI76ZAcyCiYhYYDuCjTws/1yNptVXiVvl55alvw8D2sxBuIj
DcQqqkBza6ERJbf+n89r8cOuIqUBqS+MIqLjVF8g8fIjfMFm9tnX+Oq8p3N0aHf/D7pAo/HddmUk
o7pzfyE5eBR9VUkpV75bl/yFtm/iNZoMlTSy8NgwTXMfra/4A2oIrk6lQsWoE3+OI7TJMB3Qm/od
30FsRRQbh7HknceNCT2Eyf1kDjfxMnXoXnbNxPIh3zlnQqlcfIxPqTK5jqWdSBTUVDw53ZX/O/dU
DOdOkz8ADQGgtnPRyLlV8J4l6UKlZgZar4A+ujLoxnjABosRH4HSVQbu3MkqO90WpCYIeo1T4+Ot
c/ydS9bQ2/DqFW3ukZPrl35uNmJ0SzTQICca6BpW24mH8tw72+hBEaYGBn2tZnlRBA4iSD3tdw76
6614F6DRrarY0pPT/hIk7q+mX4vMKbNgO0Rwnh3FQBl++hqLBpDzKJQxUg9StajuxymvFoOJBiAL
PceoWRXI8G/GVAy8zmq8mvk0K4rVEBzuPEA0NpxcBiXXpqxj06fbDfJuc/CSc2y/nIMaT81V0O5M
lq/ogQ6VwmxPcDkHygXb/4E31yUWKD9E51UIgoj9Yd3UCWtBZiOnvlYFeF7QA1+k/ydEXW1Do0xb
iqzh6rIkbRNmlw4ttsvII5YBssgDmBa6UT0Mln8Py6aNIS5I6at9eICHE1UyPR9JWc02glOYoIK5
jSX+2C59wRqKi/z0QDXI2M5WztKN9s+PEl1bJ5x7KNtYR5wCLtAlefwzmM5qhjNX7RBpYrVPyRli
pxXBKbbWhRzrWfg6LxpeegBye+NMBPfRMIGjA+Mbn4Lgsx14bzgl8WWTFsQb9nAQVYv/SejbJojW
ee/J+Kz1uExPLJPF4r116VI+wt2YF4dq3hLeD8rzRJHqDr5Vo/0xzs81BQ6vggUZE1Alo36PrpCe
PWN6uhFtoOjQvxjeUDWlbc8nkgR747Fc95eWyW3/bDNcDS+X/ALO9q0QDNvhcheEGX+NscnbHLCK
Ri6SIsbALU8vWnSvripKSvLGsgrffOBTfrwigf8Z9Gy3jY1S9XRG3iznUDW8OSyn4HbYDtFuU5/P
QAKJqNpfPBkC9QJ8v+f+fR7iOFjd1xaeDVpcLqexQFv3VhQ1knECr1Np+AXeXsJFISWy0gsclkdG
50tYgDm1zYXlIxW/Xa6ZHLfHeqSxZ+h1dxd9Ob2bQJaoaJx1P12+sg+esOChIZT2utgabUx6PgLD
tiUlp9/VunfOKv55R5I2YR1f5QK6ft0DJcwGC6U7c3DRylmS6FzVGCUgEuH4HduCHPp8N9CvxGUP
oulxfS9RnSTWgs3fSSg1ESV9ClQWjWYs95XoaAolI7Yw/voEAC0iovDeE3BBZea22rInAzLBDM9H
Z2l6ZGui1qmIhXfbEENJKl+hy1Wz9AulRqeIdqdHHRvi8y/NHBfzOwNU0oGaxBnoYn/tS8SfdMPP
gFJUfXvMkzpHSgD+k4VYwyxVNH1eeH7JuJ1JI76kYesajwVsfNFLe3rATvYEpSg0HfCyPcO6MgOm
n3rMokCob8uDgHj8exXDDCTzxWj9lzj0CULqIuIm5HiOXzlsrlgaXxgSgeUt6NSKgTmLmckN1ybO
3TkLVgqpyvh7I3mP5ZHEnoeqrl9fDuGbbnElh5w1p/YE5cEmPii0kXg7lm3O7yAeBrtNd4lBxxIC
1RzLnaEaQGwSKh/ZCwq3JJjXi0aEovYNvzxTsD9vESCoPW1Ezv5I/13DrV+k7x2E/l7GYNFfN4z/
cX+AuP0setlM0FdyP2Yue6wYWUfg4HjS4ru6O+4etk4qcablVXsa4+MZladWtZ/zMw+UJo7s0iOX
IDAoRF4xa/fQSwHOGScWPpuGETnl/Jq+DLob/LwI6e8m4J8lPVTFJEnG623sIKTUIa66rpNsXaln
r6t+627fHvp1HCsDH/TVZyRJaW37dIqIzRFOrQNP6l3zRQ8IZArpm80UEmVATnq6YaIhE+tvcdqt
vR7X4l99J2rGvy3MIjugLYSdRniaoXEVkGZxKHofv4HJkYXrCUr8kRg+h5jf9JyUjZtoyoLs1E8T
pwIY2heAGSAj7+kxOJ+cZBZCVwNgLhVgdbRnOjujMADwOQNz1yawB8/Ge4NPfzrUVbS2OVtnAySF
XH+vXRQhkKve7SiHG9NL6gkxwHXtmNOykYXBjGu/QeMYdxNnSVASnEoO6ncSsQ7U0Ue+usp4HL9V
Lll2HNlgDxP2yJWqXka0/dA5cWanxyhwxxbCaCPnWcyJk5qqCPkLdPI/IzMr0lTCYHmW/wEdKiad
jY0V1htVjsK6fz9ES4tSB73xmMh3H2+YNfmaGuB5KgpGvb90WTrT1UA5Q69+vZmcfIyUUpQAyJkj
YCgXjdii7iHDafvi0ubZFP+jR+L2TFb3GmzzkgN43ZgWRvXF2jLM6JXq+idCdCXxBDKYLtLZRdWL
9aLdXVuQeqNjG7X1+MfEBqpUY0Z4TbWewIuflUebrtlb5BHjG13ABcoLj266hRLOIVJ1hr3Mvgx+
ZcDNAJYhwGyvYJGebp6WU6OcuFEcc+dFK2QWJF3FsoY4P0u+XxHlcS9uzY1/kbVVDOBIjeR6+rmx
uRh7Nxuo8BDk2G4i5ojYKBF65yMHYtlQ/JM/kj7to1mHGNbAz+AxJRMmW4ubGEpElY62XBcu8iX7
0LI6COw0EeXxy23UR37jZ63wtdAxOa4KvPa+4g+qaxYwNXgm5n9KqPf+4opk4uoEHMeU0MdIkG/W
LtafIRiBazksG62c1o6aWuFlpBXLmmghKPWrghlen6F+Wh71EbVmcR+mMt1qLxjhmrdCg0J3u+AO
7OsQMUzEoFyZrQsgoPJ9moC9ehrQU88wPjxX2XWuiPC7y1Mclf9ZeRe7ZrESnfCMDdw1jFujqtoK
NmsLh3XbXcI8QJzrPg2oi5EY8g4J1IK1lgiciRf2+kg2KFJf/oMHSviHTaFXQxDLvVWbBbRHu67X
1a250i5fDM/lQIjGdNBDxiudwaIAKDVGjP9tYZfPnLdlK4EPavQ0vZBacntqtMkTPw8FNlS90/Ps
dbDnHOH1Sc4XvXSjQcIohSIuIaPEaQMv6mCw8PHb0rgu5NjT3iybyWlSHWApiXnfiZ1q+4XfilM6
Oq2tw/XBM4Z5Ml1hU75PwaqvBFwt4zsfvCnNLuRz6XI9Qle2OCMyfGzriTq96Pfph2bfjEd+98/p
2BblGhgyVmQ2Y7HrKT4fQb9k86yIwOeBVwN6XyAcGeVOPsi05W4H8mtJcqTwJ2Whr99bCxZBRN+s
+tND5sFkf1gjg+6qA1YFNFjBAkUQZZ44PKKEm3NDpWlzgGjR27mNUhYMV38LkQ2zZHkwNfLcENTp
SCix23Je+411XKxLtXp9vyrr3LvOarpSN5TU6YAant8WeMt2vAJB6iFJTKSPLOMBYuQqI4FIDcsd
Vd8uhFUZNY480byKwB1RnJaYitfzYYESYb+/tjIQmaqkYODe1q1hKN3S86nB7fFvGxLKgZ+4yxNN
JfTmivOXXEtvTQk5C2QGUJGpXoZJiFZFfhTYzLTG4eecpARo4BKfAMBq8mlqIDDMxhZyALFIHBxV
GiwNSfXrj1s5l5HnLfI+CRSFD+xrO/qSsUKxM8BO0/TQT6Pt0/Zg6yBv+gJFX5oI1IbXhEw0jDIE
GQq1tdOr1EhPwUiAQPjWTsvxQe65cXPj5FC5eF8AuYBDD3xcJhBwuOyrOvFfMQ0SheQDvmoeyttR
qNQI7Al+LpPyKKxbGxZLCnKgkANEBadIQ53paLCion8iQ8p2P5yUOorH2xFH99P/wkL+rlB51xwf
0aXnZSPkUKO9035uCPP0eWkd0pUPS50bmq1KVrcTF9UVfuo75/TI5pC6Q3CkHUv5tLpNR7P/nVNq
dphvl3YOyUG+WzRbaBLkpCxjre6uuIkBE7CjxA30t2kqqRdRKTHZXOsVlB6s8rxgZNLvupvya/Ks
yHlgJzsCG1xvrgd69RCNy3I6GmJb7J4tG3DwkjxKj07viJfIALnDJu2R5MWfyiysiv1rPNUiLLNl
Lu077KvdemhafzVDHMB3BIBZPnGZs7OBdQaMrSY422kCe7eg/85K9tyV1G7GX0jWSG8SFLGu/GlX
e4k7TuNfXBdqngrmruAVHBRW+GFt3+mOz3KSa4Imuh1XS+XjRHQLGLtRGR6bFSwGx6wmHcG4IiEK
r+VBBGxADQ+obiCqF5vXeQt8iYwkJxleFSydyLIkJBUcmU27u9sJSoDDJA+CnCEaUey2Mcq1rwNu
3m77qJ+L0yQFP+DoRdCIb7BflNwvXDG06eROvVHphCbMCv+rtuck4tk9uE6AYFOHB+Ep4igP9d8C
GqDPH+2oJ4g3NHJK6mMu2HCXGlv92adO8exTWI7xhZbcE2ql9NKUTyIx5yfV7ybDo2LzkQKEbU0h
2hGBm9wP/ylUvodP+tg1n4EDEtraRBL/BYGom+UzbHCQaMcoDtnJm+O29IoXGc4nkCjWG34FSIXU
+VBqR5qLc7ZinZQctEAdIuXzlAKzktemDJXY7IINw2xCkPE0420mhCNNvcJMuG+Jjlb72CWeJX1G
jFYgOXy3vq4XHp3e3Yk4r8bX03oKJTX0RQRtW7oiz98qk7t+K/XK8BlKfolVe/gHms5MXHHb284j
mYr8ueb3bKzR0XlejvfeFniSgyWJRqW+7xcBVNLAm35IKEYq2sQyupBdvPd+QbSZhjkqxnmnhb61
lSK58h08E0j8eZpEwB07QYJeNLKEuuTLe5bTMll9GfEs5qumBNuulwKbvojv2YaMDjDl2sB6F6jl
6FDpOuYZOXN3Qk/iGqn9X3KcTdPRIbiD0Tr5YtAuvZjIW1p82ECP0mDYjhzB4hjogFjMKgYLGUuu
HKPYz1OWqCtccwan9Oxax2Dl0RAP5D31PJlOz7p/ujTT6TKl2vtVXbXes7VRuJFc1Byj0vUon6tr
rS7FcnKxI/f2hmsVntsKglshT/iP74XyEA97B5d4ev5jc04ZxnBfja7MrcrP+D+HVUYF3IHfwkKm
6U2aR+iYu05qQ3SKGJPXKROFkgHDr3zbCutJ6T/3DddsU1MIMLZsaPWmLG8RvpTFIbWfBCXliR1z
4NGJn1xKs9OhK067pzNWEPUn5Xt6tgrb5yGKK21WXU5tTgZOmiKa2O+NbVbUvx8LoTzo7H7OvJMu
muxMGF39UZpFV5aNbu2MlEO1098spVpK3OoioMM3rj28Khg0yYqZ1MAwUYsxRsRSlkS++lhayBFB
iTooHGx4j7Lf4XvuKYmHNPmNVmvR6DbjUWj9jIX/6iA86NKzcaiGELCTvgZKC8TpprjeR5jnee/s
h14EzPxKG70fHdUMngw0NYu33gpmi+0PVlzQH+sfAYsDJfgBHybhRDcozmCp3chMYA7hHvtHmsK0
B5j5K3hc8mLgGJGPkkXKNNciKWGO4JGxD4NR1avLnRUNZNAf3sS65oa6imrPMlm4I4NVuk69qWsL
zdIRdxFZ1j2lpzH3ez6xsKvnrI+49ZspGs5OV8wyU7CKLpuuGgQWmQ0kBwG4nDP+ioGuO2BwHNel
bmWYNWUUmusBju0WRzk5ojrGaKE2CV8VYjrVl8BNcmrY8Ihd5Nnymm0ANLQlDbWrguxoStFgXB5X
zCbqiIID3icd2kInc8qVMc3k5osdGA8rgRVYxHWGtpAONJFU+fbv2I2ca2Z3dd9BTi6fVswuJ7wG
HlD2Xl6QvgbQzheTjzwkhFdpRUzhUhN70rT4KHfQhPyb7dS0WNA2jVejOn+lgp3dc5o2ZQefiXVE
dnDzRmrHn3XtLJZi8o+lha/0WmE9s+kiNxmQPfCG+CuUgVAoCrDY1bCtUWhhFgGxIW6/113j5hVy
HrWTLOfyCmeizxFxAj7KS8XNJjH8H6Vs0+26r7Wm1ag9dZ9mdwO4nBi5HC//yKOOqUntkpPr12M+
dNSDnHMvZjBMi7abmxSa2cxrr46nbbB+RdawZx8ufe9K8s/FsouSsOpUu+ZCSCoElXBSpivY1e2g
eBTjxNe/8z/RaLKAC7sIrew1EBwGoeSZ+5CgfUkWCPdO3vvTP6kKrGqfqldnpWFXomz++bVj7VC5
kXQDgPPsB3wvqVYBKaAYPrSbbXPnK5R2g3xwmWNZZ0n4mRV5GXHiiJBwqp5nOgUrFyRUywwVPjqC
K6+71HFcH0eMp+aMPT+/jMT9BHlcVIiXKCzBrAHIhApsS/qV+Gx6Ybztgb9qGJ3VIs+SA43nMQyB
6CGPg+ICKzt3JGP+Su6mmgOF6dj6l5Aw1k+Q31mNp3/7Ph9IMKplZzJO6cJ5PiYcbVvwHxZnlEIP
FUDU52W65BwJkhq63LdtVL4pOVxIY64N3RiFhmqjSUEdZr+oe8whXrQMqbnXAb7pFcU9VFOE/MiT
SHqA+yALPurx8CImRFPEfONO9wb6m7hkJAy9u8RE8Zi/0g91dWeJyuBQIheqlkNA/qhSZlpwD1cx
iDtkm99Q9oSJX7szOIzR23HrZwGKG1uMvWRTh/SZG+/4NvjZihOb1kC+A3UynKKAah3/4sZ8perA
evB9daK5XHATd9RlI1sLs+zvPLwD2rUa2MIpJaGckVViTFWS5Q7cOby1TL2CnOUh6jbXyp4eGTC8
WX40ctzlactBd309+b/Hg4bRaVzRp2T9zWzQG+CD6fbSoSWeZRLUy/hM7l4gxYgfufTAHpJ8VNiV
u9SiXdoKtD0MIJ4aWJn8CEZU60MSwKuqEGMmnlhyAIcXCMu/6qnD8WTuVdOpcRMPlGetNilj2vQ4
BtTISLclszd83UjGx2JHNhZxhlQgPs4LHfhePeGyvQTdPkXztgDo1qNqUnC2fyzc0XudbTWTK4Rf
x4gNTLL8mka9xjkhngMuIXsUCD9vyQrwvxIovHVHHRbOavOFF1/4flk423K5MEq2+f81HaBlHW+Z
y7Vlnubpc8rlNrFv/CvwNYKI929syD5hWnr9DGYGpPRt9Acfhcwmwa8Ic8wPQ53onPEpoWQ5D109
KzYDvgKIjTEP6JCXl3jCVEQ7YxYrq+9S+YfkitLh7wIV2hrR8jdyt4XHKGTG5qiXEv0Dm9TnFjC6
CXlYeUxm/5yFthba9dNAET2V81favs1dytaInLws+f/2xAj4CjQCBQTgabziDEJmoPnVjySqP0Ug
lScql+C5ppOPBqI27YA2+1hNuUlmH1JZ1t15ZxKSrhIvpKEWMku2/t9H8yy6IK75rg479Yaccd/Z
WE/Re7cEX8qYmr6M7rXE3VRMKSDNVq/ysb44yHS/nm/+cSAMZNEeIDvTXWS4H3x1QHRS4QMX8M0N
zjXNxBO75gkkfkHrd/qZIYtoxtbbd+6DtLnGZj9G6UZYZMHbYtUXv8h5ikl7LaKmXZUutuoogd8t
lzpIuQ7xHpxJggNomFPrvrW1+g74m9a0yGIWhpwIeM2lyTlnoi6lc196EJFXJrh/nILvZ3KVjOwf
7z/KhsRhK8CZLedtvhQdQmgtjq4V1RCvreb6aK0bEf+VKHnFi7lSkiIVM5kKDPGlrxkiM6IjhLoh
PbidSeU+qaakrEJaSd95cBbgCoFPlktwBb7zQ5zrBIaFby6BG/2lj9PrPT4HvNkrhROwoP6TIgu+
toVnDmo4EpxVEceqbqRGqEV6anXR12ev5yAO8/in5kBWYfDC/ity2Wbp/qGDSwtgE3HIA7KT0m21
Klw0ARAoXHRWEVIpqKqrLo2C70W8ElkQxnXyD5l0XNz/jypOSrobPNE5HpHygEskNQvsL8PJK8rA
tOOCL0T9fE9b4ZAirZD4dej7LkquZsNjvIf4+1OfEfkjf1L6lMMC7X/nG+LWelZqV0zoaxfXvKsr
scUvTEGUCOGHUuF+cHG13aBzNs0iHC6yOMeZ2+2vjhCDApZtA3D4URU9XYT9U7qOXevta7ugiFZp
jSD02phWZVHi/TNtO9O4BvNl9ElgkRT4CaqUSMKDDKfCVDH7aT9ABjxqF/yoAav43IEpGmHNwqzK
mhBgFXWi6HkILJBvvWRmvhWKkCz+UHBdQmUgr2WDvEQ18iyIekty5mZB4/Vv9w84rOO/ly1q0b5P
o+Sc5WhP9VAVLPdDyuYx8R1JXphXdFWtXhFdR3301EtRpJ4C2GABMLf+pqEANgTeecfCrM7DwpLF
vV/g6GaPJnfx+Mwo8fW3Fa44qyKTEzdAvMrrh2N1+ncChz6BS0j+sjG+UtwaRnVp4alm2qsELH1m
1FFFD3evC0nsnjN2KpNAulyHs4GecqJTmK36+bw/KP8PZZVjqFDKtcPrJjtCm5gUBIVXtoN0CAD/
pge99CDm4+IwACftwz5+K7hGK9i7xkah2EhINh5cObsUtq0Rx2QrXwFXCUC3eCOjNob0Zth+BbIi
paAlTRATMVCN35BP4W+JRODzeCualfkhNFkIN4Bktn1a9Yeo1J9gfXe5lnQcv0RsCEUASxK9PdSD
rm/WJ+n+nncWJuVPfYA1VKAE1Z0hVTACS51hyqPrssqp5VqmR0yHhBw85yI7MbBo3BAwxjrDlvh1
yLLX6FK5jjaZJOk3TZDWoXOBflUJe+5glzvGzEnLsM21zVqI3RQh5DeXkgt23puQEKglNWk1JRbr
rDvG0xUw8PN27QxKOFC6VqAupKDeVuHRWZNyNbfD3HLIvS7lpnVQ6CgEOFLG2Tj9fLCFlyoqUtrU
mGI8SU2S7Z3DP0hwR8bg536oHD2U/1umIRrBGQUxW6/ulhyeboFRducF2rJ8Eaj1JCHt/QYggLJE
FmlutUw+WdZgTF6waTMEcC8p0+5s2i2w01X8TFWDYU7/8qQ3NbZj7B1TLk1MNguC7TMTEYMj+3+q
XLs4V3LUp2H5ykajMm+2ZTd6UdIDTl7DILVQRPTRQ8bGS0efTD98zHci24iWWDlnWLnGuiKChV1t
00CwF03jbEchewXrNtyJhCbuf4O4C064/Uacb7sGzUGtVfI0tWjCjMnlgjAro5FxplEKzdzWM97K
iJG/1UYOEvWCH2cLl999WLPO4wJ60QqAs6M4Eb56VKdlddvj7FmRyyoDCB2yd5+OwwW6mjSg9z1d
NioRwgu6PQFpwC39zPc6xdOwcWQCFfDz0w3+THGAkyY6NuOxNDqmKgxh23E9b9vOrXUGIg4HKmgj
5n/3g5xGQf8EK9+i1E0WlfntK5gb8G0Pv39Bg0Rfn1Cn/5GOUH6CxkKaWIy/flRsJ04/6U1vvBbi
L3s2LsGuK/Dj34uKySe3Twdaj3jqxbcpUmvc76ERKF0kOv3FdLNUi+cgYtioS+K9XVbXDr4rb5lW
IP/pRzFN/TnmfItalk3Oti8jLRNVwFbT2znx0sZWKvH6LFc1wxtKfO/w0+nm2B5KYn9VjIhWqkKj
GT+vFTiO+pNhwIoSpXSm2YQ1qgzP2/X00YTzdQ8LDArSZkIUtnphJ1QqiVGiuV4dnHhfI64TU4YI
bvDgP+RmMFyqgaz7F3SJWgTDB4mg7RHYWDF5rBzAfNmeBcnXJ1qiFdNyWujGxp8+RPLU5zyhae7H
Z9QaPEPhQ4ngpdg1rNfmpKt/qFXjqHWWhOgDPLuI31vnrYpb4Hd58iVRTRejRSyRfrjxIUIdZd+m
WwmQ4avG83db/+fyxPLfFlYCjuDlS3g+ahXAp6xhn1ljJhVXkJj9pbI5t8sy3ngjvpJCrctXLz4X
OThru8ybFzJ3lOmitsJsW+0X5wMMXXwtUrVAuzcO5HX8UM1uCL07SzyVDMMSp1BEvhwJFxsoMLsj
RKEwbDhkXTuTO0tQhhBn+dB1wov8ABGv/d46DRDqkNw+Hp0uleiccTKEUnsb0kL7MowolJtphprT
MSPbfXQNtc1KsIgW9nnI7Hpaxu+a0FM3HKkUEucwz34ROGabMGamPsoM7SJXH4sqf9yIeH2crY+g
eAtQu+hxygNudeb4ZERW6xR0N9KMu8VyJT9HdK8A5kyQhI/NyJ60kE2qRBcvP/c6AFZuk9dcO2W9
04Gax8WLYY1fv6YNtQQjnVrMw2Ohgu9m1iqi/xNf9qWJA0tgqhH+AqlrC3D9SgFeEuPmZVbscBus
pJcBuLI1LCNYj0dJt4zaw4SolnsBaPTURkpQrfkU+XVGS2isNnt9e3XZE9EdnPQbD6b3/pYBAQ4g
4aiJVYBXY+JxW9ASJKpK/iWQbbKBB5aBfXbbvjMQzZsGt16A9+blaseTJkGpXsvtqL+PGTEZVHi5
B8NnO16uWfjf7bS2GyZfwF6rJ/Vjx2Ig25nvG/FdR6ntI9dEcy4lhoimSGlt+rBTfCFTl+ATS5K2
AiOoN7LeUrjTVlQpFXLbu6+acynnOz93i6ZBw9M7ViJ0Xkr5huZcKyvlgZgq4xT7Tgl9S/O3Xk0O
MpetFpLQPVCBJtk4+7Pf6fkJEWIwkQsWW/8rxYdRw11r7GylI8LUegctYmjxAo6O0vF0YSiC7v5M
cXY/XK2OS3Y5voKJcyfrj/mwUcIBNxAkEESzcaD8mKJd4Wy5N7cuhEJUr60hPqfU6LbGtx5FVMPQ
QtwTdFznVmCevQmNAIh62KBnSR2Id3wUUe24ESS99J2R5vRNqB9L0yar5iSubJvZ9KlxjxisQppK
+8YXWTABoax8+AoSsGgJrDd6VGE3LAkBUTnpCffBdz99XsAze+HxjCr7MqFSY42qyYhwQxAU9WuX
D2cgFL1L1F72AxEscwuTHIsLeJALxPHZ+3naCZpMViEIud0SJkSzH8gXF8ZSn0PabguvP5xaBQzV
GkF8NwZGgJ3iwb/eK+G9d6ETAG8OwnLsWfz6YgCcl1WsAcqE5qlcCSuJwIoQdz+nPTbg/7IoPlYG
Rpx5KIs8HpvfYd/S3d+km7wbvxEiM2PgGPXzfIsokv7coSHjzVCNGvaGom6iglCImjQ4RCL7uzGN
8RPhDruSGvGLuxrzG90rCvtuE09Hfe4UoK8oqGVNmlSEa+Lshvj+vsTQj9jU4nTvXbjmasuotr8l
tqFLDVxu++1PRPUuuIEoRGv/LBW1pJULj+Qs9EFMdwmq6c8iRs2i8kjM77pRe+cU/vZvg7Ukd3kq
sLzYGXt4zfs0lvH94ADT/uetmhrTKkvBFuV7RjpcxFlE/r08QPKM3dMAOXNSriVnMseKmuqIIlJr
qpJroavG5wpP5QXBB2wZFtZdO5BLHLpC6KY7gGiZNFFNw4SKrOfYaTe/OwRWUaMdZ5jATIgV4+MA
8za+9PlWHSIAo9vaHZdfekQO/07pxPWxH95hncIFPlXkEw5/ImTU4ueSUhVsH0PowiAHpXsuEBWN
tg6kEP8c+++4brnx+VJ0Y6ZDFu4lFB47hNOgtjzRFF/ZIH/QbBD8O7ewY0UJ2c+LV9jVySCkUps9
ayDI2zjvoGlMOsaMG61vQKijGSXRImaLIXHfmrDXOM8Sntj4fqbUFL8eAmo2XFcHqyIOWLu/Oa3i
h5cztE1ErU/wf149xex4vLFjZ7QPuanKwjyQucUDOIof+D1yTiJcpqzZ2+XMu7wWLM+q9LPNMlCK
0ak8O6V1+q9PzzOXStkIErlko9u6YI18jE3XaFFmnFOOr5eM/t34PnqaKmTekNUxkOjDvmzOEkVN
ucLIMCbu7klGB22bUm/5Q4wNmP1hIk7lersDYFLcnI51S2EaW1Navs/gMlrs+uEs49+soCvyxUg3
tJYHSsGpryHXilaST5Y3ulLvNGi7Ya40cciSYirQWoV+BlvM0ke/u1C01SQ3WDLI2T004vH8H794
mjsMZVgj/S0gGPaQJX0tADr4CZ116AudRIO1U2VuGVTlaiKXiodj4aW4N7vNVHj6U5oVaUfCIRQS
J42W3WtGhs/fixJD2t1kU9X9l951wwYBW+kVrHTASXVbchl7Z2Z0rZ0ZSpyErHYZGQuu6kJ0slxU
JeES7JiM4VWrtga/oT+b3SF+CaQ2kb1n/niiLssm93ulHEDQNNLiHEBvX7Tk55CmvE+LZU6Mlf32
ShBESb78MOg/K7oXdmi/QBsb0K4HCXu07R//B4qGjrbY5b9ZfSCnpFF9AZn0Qc/l4wJvOknjafR6
HbERYJQoADV1m60iTLkdFXVTfPk0JMYplDuGHRCzyYdZlHbU0tfihbeHShuN5ni9ZM55OXgpLq/I
jjXpDOgYREe270Alt8NSAKX19YgubtYCS8gAMZreBY0lJJ0dG1n4w71qwZLevz8FUVLl6OnvKYH1
Mi3RCAcnzzdq06kZFqUzV0RKrHeKOyIEjDtbMiiBg06RNgMsmgcGFpDxhfoMCvvPTP7w1Fgbs5yf
yW43uQ1DAcky4HSbkQUPgNwhx3Rn2KWCJdgmhxAgOLVrX1+a14UphqInLdePzQRe0nn3PFgEz+EP
LXlbZ6XLrOu9/JCzAcIAHf4h0ke9uLwpIqMx92hHLfO/7JeW71DfynRkSZyLdBSGhN8lhn2Hplbw
OID+jOcdp/Ov9qE5c1hXmxOlh4ormovZWHyh3hji55aTrTGcXYLR/8Zh9c+gN0dkyCh/m+423LEF
3lWOuDzRfM5KqR59v2VD9YalRK0gjWTiuEz7b6BuQoXizOUFuhiCIU0uhAWLSQlzq6wMCrFN/ZPN
ybA1U50EsCwdgO3t0dgqftevS8J9lHt6z6v+RPcrlXt6ghSidY4dDcKFryn6rWp2hqLObKkph7ih
P3RsDkpJTw9FFc9B16+uGCA8qxKi0AGAiXEd7JpzKOwvfMw99SRj6cAIrCfOtGitQ03+NYgGiTqA
bmNNFHczW0ghB02jdQ6ipFrKKh4+wZwrjpxIDY/+pzcgCewcRQZ+qg4rGI4aBXj6F3lrAsdXgAQW
CCm8TxGLhWYl9aezO0WpzMZJNvnwyxVcFyjDLUQZfqn3p9fEFfvFNP0ln5tfFRRJ3eCSuWDa9bUj
/3P5bSs6gLtagJUBGqaH7yVTK6iP/nid46n9chho5cGYihvBFI6A+1079m+O7SHGtbDZs2T9j3vi
zneRDGDla42ZN2mZ1IA8TjBIsHV/1TH/h7UQMoex8Y1VM0tzzwzcVDcaK59B88CPWpWMjcgVCg5j
OpP7kQNqHGl7eacVIDwVg213zJGGIonHQ4v2U4pPSHVMGi18LXtSpI5FeT2rHV9Ki3WfoMWDgNb6
2SBxYkzr7XFkjg8XF4Qg0JN2lXzR5haWxWDaMeTynGyGLJ6wUjZ+bgKRwOpCou71aGxdg2Trcw/K
5hSOISvZ0CGz1baxnbnQ524dhYkfCdMetoXNi1cmjWtjPJRFLbQLWAnF+7P48RwiV+GesWw5wwlK
WHt71KJEIZhHaaFfUE0PdJHdWDAkzR4Y2RRYTaqiQnWA88pT+f/o0LQ3MgCM8sfHzfyvobrXF3gA
xBDaffXSNfXGxaz3T237UkYQDEsrdDSTP7ygRaQMXCoDXFxJdirDXshC04Yd8CmcTsL3Lq2cGT3r
H/q7vFVfQrZZl+vFHZGhwS6XK4cidq2ZTyIq7jaNR35m5iJbao4Bmz9/BM4tCkILRFY+OG+AzawY
3Iw2t511qlR7XgroE/2H7ruy81qEoytaB5hn/6GppZ3cDU2qpF5D2v/RgMPeBlbLgXJ1OGGrtnaq
IbrMDk45/j3UCV1RfX/X4Gv0OuM9zVDejmPHhH+cJGiYMWKwVUsrdMLhrRta/ogoHiKXaj/tqEED
3/PwRYeHoucu9+SL5yyEoKZvS+pOYcy2zNUArBGrQ4LNWbP00+YM4Wz/3eTyPUx+/bRWrPr7ypC4
rSZOkgEeXFB9frp28P+fV+sXUiV3aNHdWcHvO5R6AZZheEhR54IC3P1hCs0TLsEPB98YF6U8u+8L
tmcFVRlOFMgo7tsVr4EkGVrkjXe3l6uHj2fKcFKroRtmIGk5scq2SX6Jr8tpApXmZQnMd7XtqBgy
jMZdrjQZZ75nw7APG815NJM3xcCvjYmoVgWQ9BOGf5lpEgL6sVOk5I8GjnlJ1yJ/v5CKmYfzDK6w
lgnsUrWw52Hdk2QWXeqrUez6erQAun8qdIwxkl+DLmoFCTeTQF8eFn57ZwaFN5GXOJtK6O221T2D
tn+FxhCB23EJQ+Nief+c96rIzdJZ2rapU5WLyDGLxHpVMmrjXndT0cRz7fmZOASFPuf8yE+YEALb
ulN4JMi8YvcKRYw9fFYkdH1Mk2F371dkVtnx8bYv/iDhun5q3n4ql/oCF6T3kHB4aRKYwAhg76JG
YG6YZVmDVwJEBEw1w/2QwOnD9I1Rxp6v2uhVPqpAuoIDXzGhuvmethZkA5HEG3xkvpq2HuqriOly
jnLhcDFyaBYNImZ5eXorPFelOlAtVHyBlHXqs9PqPfyKu8yWCvt3fEbfhGCKB37ZeY5eOgaLjNot
WC8+10bMXllfGqaMPC9BNmHd2IuWhzZKAjg/b5aM7mOB19N5GYoVy0o6VrncN2VzWMJ7vahLSYmR
dlc95yri4z2W18vJj39Pxi8fJUyVF+vXJaInGUY4L7R8Em/DFaFWeVVHK4VRyRKdtHuNagaraTxq
+O3Ya3csarFAVp2UAymLneEopEC5h5de86a1oNfGwoQmD2YeRW26xwTQXju5BauNB25pggVTkjeX
QN0Mt/yrpVcecI+WJI+ky44mrBmEV9vwAmPKpzAkZj7oJ5vq2AXhlcJ3yN5MwZKa4McIbI/R2BJe
jUxlwJtpbZX+fAynBiwcO/QJbsweK6tiq2ePx0c92plykFEuoMISw3EvR7fuMgB+/4F3SmSQjv3D
YoQNeOIBASAquMd6s9SzSV1JH7PDBOX/YQCg0xYcmbeuuJ7q7OY0TSpyqtitbIw7QRoYJW9UngEj
jSxaIK/SfPsFtLHsTiESttIKgakQ0TB5sK/m0OU7bzhz70/77EuUyNj94Imb64uktAT9c4dslAG/
fHR7ZCjreDbXwFaN4hJvPo+3OqkAgWXJBSfk6YNKoXy57q3gJQcw7aSfmkIwByFFoxUYoz5DdnTz
p0TykMHVCUjNpciq9BzYqRTB7Ebm3sni7byMn5Ncg4ZqKCGJLNHo8SR48dn5Yv68ijpfrJL6QxgT
gHBnpB1eURFpzBetY0q8kTucxwj2SvzKpVOpBV5yCsXl+BP3Qadl+U8WdkDnNcXG2RLFLZH76TV2
Xt8aFOgBI2QZHV5tg9NUG9fj3mRfIr1o9Iq4sEl56rRaGBVdzlP1EDdTuVQB53BmlFwZsr75A9tB
6gLVpPQ8PBoix0r4wsWbdTfEYQxUNpnqp6abl3xmdJNdmVrsoJjptSyqC7N7cxvj4PYQUAA5TMGi
C4PoLYPo3M0ch5td1VCxCaizByLryH6pPmVs/u/nd4FU9o9CKOgG7EP85hjpE+xVWZ9dgl2L9586
l907svkqg+lBcVBI3IwD1FzYR/CofuEMP34Wwpa1AYgyfjBLTFqwdnGI8lieh5rd6leZBOF+8S0r
t6+/zAxAgn9iaY6KSf1JjAEKbNPTv7ghai7CaeEgZ+zP0I+6AKCMqu/cW3kY5ZCRO1o0ENUgHHXz
81ojaywCQY+oA/kHdajDYznNKYsU+5bwbPzfftNQYRs4L8a14BleZ4nO65DqZEB0U+d+niXnh2Qh
3ZMzMxEUuC/xZduZ0wrIic666aJ9TRE8fMXXXSt4rXvJWXC2BX4XhUXBiuqWtMBCfllYq7Bw7erF
8e1J7V5YybuBT8WuE3aGwtz7MUEHleQKS8JOQAdHt49CLmsmoFm9n/nbigLcIvzfOK9xgka++aPk
UVrJZRozs637yyvtXfadCvEAeCV/EsJn5Q4lammgnnCrV4xhEeHGuWuhRkXycYQA9EzLvB0uBCUG
J8CVdu1cX2Yf0EOrXRBWx32oAcbDq3wTJ09LWY+9uZicsdrOegHs0JHCneSFZ+juQ8rdywDD0i/z
FxFryKaOXQv9U2oDd3cHTsbPWKUji2aTPk1uyt6X6y5nmvYKzmLfdmXIVj/uJ/T4t7uxc+aiI6MA
B4+wp2DnNJGYfMHD811Qk4+2+0k7DRYmWf2p5IibZ+rjI6kuEufKFlV+FAfT8C0GFzLgGuUu8Z7u
Lw7HCEW7f3T9P4vvgZyqoWZKJGeZZSpPDCsWqseb9TzFLde/SZIozBNwZfUIip+J62A5LH/5KVod
UokwAk9Dm+3JSMhgAvhFtl8QAmfYH1R7olsSXmSOxpQfClwszPgigVmQMEM4o28snXFXm5ZtvorU
2VhLOOsEwzuN1iVVFE2camjiQinXq+4ghkXtoHrZ7wCUCzJkFQcQpfpxN6vuHy84v55pkhYnBPru
9h8jmUyrGny4VIPzjWi/dWO6tUa9x4j9jekvA9MgjjOo3VNcxisQD3Gt7VKR/mI48ksWePPVLLkx
Nc44bMRO3gnO1mNHGEJ9pNOcwsYANHRPJkowIKQKp+MG5ssKimCGAKxbfaZmY5je9iHG01MN4IVH
s2EjNVCMYx6XtKwIJA6NxGaMb7rYqcNVmGe/cPLWjGkPDchBzCtSlH5TWYI7x3xLwOBCsctjHELg
cSkpuMIJceoWkiaOlqy2IvazzUqKuMX/09hBbhr+w2MScaFuFMEC7FSg0iBiFpolwaqSSYcwUrkB
t1I9RTNfnSTM/k8LTYi03iqJ4SPxZW0aVNonkg3vBO0Vvd8Go8jsYWiWDkQJh56f0hid40nvDheQ
M1mzYgPKx8z2s1RuwPFeLE8c7oKZ8PTbP/5me9k6+lxVjYjjqdGdS3AWcbvyc0I8i2jPOO08mADP
3RZSjJYxSkq8AjvhbIzqj4JJSI1O6ka7RfahvA+c6+AmJInmo5kIsC+RBWLABmdCToqP9+HKa/wn
Q4mxOmVQqiuYquRYNTofB8a1+WmDCCmKJ19CQ8GMVKnzLfpxcZWbjQnT7TwdQkZUEaWulzkM4O1a
i31Qvvp34MYVQh//I/0a+KEnUrM4lzhiHuGyrxZLp3/+uKglfBxs96hUCWVMAgLvgAsRH+m6NSzk
hDZJRw/QXdLOItzrOrgw6cCNGk4tFPXDmw+vGRp80q5rtNrdy1XgLpvMLTiKmLyk+RrsWEl6LQk2
1lHyEJduDjxsNb0qDwVbK6VlVgxmTQyzZb0CauTI+ORhEA2XV2SjoEQov/9RH0OI/sfCUlEhyz9/
gqOt8o4iBqjDim2IX3RhOdn2t7fzNIgINQSRTrOW0gP+wxoMmYFTEJuJ+/ROmcvxfFWM4MiUYDik
N5mmlnMPltjgkPZrH3+0jVxgOMNhhgfDP+5391N5dffzn51LbZAXryNc4Jq59sd8F2WKI6Xwhxfq
7VW2y/ir8+eUPRY5RexDHVeKaZ+1m/9/V14Mh3/556l7TgVzHQp7mOhG+Nn+V2UGZ59R43d0R81k
MkDoI8WK5/rYbPtZz1fdwV5JYlyAvx1Kzsie20nxJDNPmPVwo6rKqFpkp+sKMXs3gk9kWpcjrixv
XRvMfaNbnyA0GnZIjeBvcqs621an/JM75dQybd28J1HY2bIURdnyAYYVYPGbrP26milUcPHPE9RM
Jr+P133yl962XIPAK/75GBV8cXhMaBxsOuXQZWoLUaKEGDASHQeaS91oYZjdk1ZSsLIraIdW5048
Y4rgI+Rvutcbs1hXSsl4FlNN2a2HruZ2MYU1PIjCi3GVT9VPlaQ/JnHfK2yqaOYCCUIUOLM3VhMJ
fSj6pNFYGckojBq8bYTDqMxg0p7++yKdf2Kz+m2aYBYYh06TBVbYuC7zr2i6wxVH3Ae8OrbVlc+a
2TxmhtFtmf9X587mw1U1q9wVcztyo0rDQ+NwwFAEsChT1FkCUYBL0EEACoYRjYPP0fd96z9kVmnG
qENEUgwCucoZlWb6rXcfUxfc7S/wqFuuGGl4xlSop/BOWpRKKgHVLmxUCMbe8deFG38aFBDgOQN2
6JtXTekZkN9FvXD8ZpuCAafwrzHj5LDk8R6gTLFIzpH0kYCPiNUVAKgvs6wgUWqYnnhekVlU5dnP
3t4rOs6fZiWW6rKUMkZytpaQzaoOg0/OcRjkVdU35OVdVIMdDvac+7kw1Lz2jBVKkzYGk4kyJZ0W
+1qTFrmQpfSQl9KHPnZlMD/5brINHJV9NoxXWrZKjaMh+mZXGocguj5EAhB3/tSiWbYYLYx5Kzw6
WHvEU2EJ05jjtaXqXIyNd/eiqjH1wINnNIPnJBzM2o6XFY1TWOVUv/YRZS3A4+DsgU+PYe9xF5OL
TnLRFhPKzmRxJuYj4RReu0R0rOma3S8kgCvu3dOBtfgdCL2d3tcw1nxqJkFaMboOyCp0iIJtb1lM
21dkX50Flh5tUI0T/ZMqFCaYvi3hn3bXxLbgZ8ZxjyWtTSVQUqV7zwImEw2p8IKAeSXBeFiFyvkR
8bk26aC65/Xk5S+lyTwQnq0xXoXhZLbKujyQjr0mV9iNui6nQnFW/iSpRHCLreJo9+ednNlIIEno
dxeRYIjaCHHm4R8qkGu/jOi/5OHOFvHsSRwAVMd8/c3ReaiCdhEPLBQwOjhRWKoEBtScE0iq4rUz
fDPfH1B61fHL+ljyIPQdicX7JicWZsPhKn2qseKHnd3/RG6W9SGsme0CKP2oWqJ0oDFEbxoejzsR
95gX0lSG8NHxJC2so64irP6A8UwX9iShTosi4Wd4WlQf2rD08R6WUgoLkATVdLk0ezBUjwwWPS9y
QkuJiYwvvIzS/bkgGephyOW1u31shL2yZcxCK2VPSryzcLFabXuDUQpeXPciw1QtE4o6l9KiXyZg
9DSpljCzsee7KfZ/AWrjSIQoKCtliKZ6xz5MhqB69TUBxJR6rlIYvKNEVN/YiiAofRP5YNFIDqe3
ViqXyjKx7cWBiH+vtdWsIpLLy/XFJr3ijt3y4O1+yJjGuSFQLVEXMK9gBT17TSf8RmlRi6mXRLdx
pXHS7HCG8KsRGCc7TdqReAJxC5xkUZ6lrmAM05tnsV2Jy+XEyr/Y317mRU3vqRibdmEA9DYbjybQ
SvTEHWDKfru0m09LsaWz3wWDJfj7cdmdKxDYaiVB4J8vMM+ig1v3ePeIblovn0grgcIgUwbL83/0
LflF1b6KjMQ3O03nVpqk53DkjTjQeARtcOBpm0NNkVufiCB9HkWrn5CfPY1z4SbFjyrzLIIW6tHw
wnzX2ZLGycVA97wBbR8XUCsIje9fe7FKsCpkOp1lK8WKbIBYUQo/eCv4ipfgjJ6gDytNZ4ABwPsH
zyMsAuJ9Dmwree2x6l23u4UGR0OjPk6eP+0UBX0WiDsGUUF81dXJew0Pj+AB4eNZJvO7RlukMvTO
63Ix6B1pIOuPj8KDRPvJ9N0aOWqnbLadL7hqQnuxrPZWxE4hNlei3USwaw/6r73qET5jCQxCgVDx
VRRZIfSQmTXXicBvx+iW65ScOx4Xh7d0jOYfcsqfjd56o902ztqAnNhMfNj/4BCgBNMME2EhSv75
MqG4VEwRkwSJHkmNxgXAZtLe5nIwf0eYY9zT9NYIj8ijn38CsoZewqikty447j9mR4QTHp12vd7o
GETPM49w8L/Rf2v6rtLrsLI8gfVR+SHq0ttpdIFxAOuHsd+js1UQTTR56rv05GQ9m0SwyQuSAhJU
K6YwgnHaqhopva8r9KuJIQsQK+rrV2pVPhlw21QapMEeyWNCD3AiQVp7AnA2pJ4uX64oNUaUkUQY
DmdM3wLMTUC52nvwkgHV1l0INFMgwwpTnqPpZ9fv7Hceg18v4EqiG5DoKNQ1yph5Gv7IJbHeu9to
e80Yrn3ia/f/PcO/zVsfOMSIVBjblt3Ajz7MqHPS39FApgB15prsO8sAbF3XLNLicAmNKsG8DuZ9
sFk7Kxx/1L9V793XDd3oBi398/tsu8qsxqwu4VWsOsxKxtY9bOw1Df3a4eoGbtdZBtDd4ebbzWKw
X3a9ZXAx2HC6g+qLytlLnndL40OhOvu84sg5mV23SNJew9/pfCMFsUd1dImWey+cxUxpDZTpamJh
b+pE+qOy7wKzsZkX+4Yk+Wy2itG62JOaKTY8YG3zimzJNmr05pUYjLNV4Mq8KeaMSmhxB9kpmZ2b
uoCYvsP9Z5RQNTQskjtelnSEa+eJ9Nc/VkjO0IiqkktWf3bp2XpaohKJm6Nw8YRGtHjoLJc4NAYd
6/H52pIlJZWPWDIh1OS14d57sa/MVXnZNRQb65EVBR0U6JBPFiMcZ/9s0Y0OsqpalU8+p32NpH5h
4pqnVbDmbYd/2CesWHE2klhH0d8xVGKykErYKQdBxqPYt534RLUAKxbvzemlImU3wSaqKR9aghL+
xa9BHbiqiD5DSRmUzX8sqA4DeRJaOpxn8Toz8Nwlya1283EpA7u00/CbohPWlNdSezAbuuVLMtSf
wGBxZ4iMoCK0LpHyjWV5KQPiD9XvVrWdlldT3yv0CvFLg6j2H7MYFVb5DrrSmIJKkBJiebi8zBGk
4M5Qn5gfVKcaYNNx/xmw9hq0Ukewi+tzm6x7DdOeuL4+Rj2O3Ds8fd6ykxmlCvQW+zN+tbbrrBer
Mgcqy+2K8GXo6GiOhU13m+M47JNDJMJSYS5GAdJzTrN0EgtDGQHYvlUzc8LXg35ntsCcz2OERZwa
+icEarmvSE7/Qivn1de4KuEKsPUn/FomN399IxQZhPDmoA6vFzbb6k4oIT6/Y+BwZHmTJuyWsdH9
ctxUdJFLegisa22v0yphusLgwqhnH7qfDTNr8I287o3Ym0Rl86xHS9qiaeD1kU3l8jQCTCLve8vk
Dxi/6ytxMRlAqSsCyaStYH26/w9hX7tWyiqC3fwLeoGFa0IceuGUfC0JwADWnZ+Q7Tt4N+Y9Lhay
giLVOlLtpk3749Ogt1smu/qEp4FcyxgULDicMA0guxMosHH62csxPxEL46XMTjjHW6QX9zcveevB
esoxfiJnHWBsEmEjPQPwiNqVYkY6crhdZaxkCfPpKkeRrCif+heOY7nM1g/UMWuZThgV/fkT2DI1
M1e1ZyCgeVc6iqBDpJYHUn8NbqbBsMUGiP4Uo6KSkw10bhkGPDnxb7Se16t37/lBmNlWVn54Nh26
mUqgnYDIBHqnjaoX42RHd/WnfgGcn+UDPhb6xiu7t1WPsmwRTewLLVJ6RO2SduozGSfpF3YtpLru
JauUGJMzL6TD2zoyjyUJMq/19TuxfE+OLq2kcKKMzycbZpglF0qOmS0d/Q+qq4/D/75976gD/sQH
pXuY0pTUMAyZ8ZA9eC1NloHYBcQRA2Jrh8FvPtOhpnO2NUzbOQemLC1EbdftLpfhBOD7qWRL6yxS
xhr3knUAP6CFcZhq8KDbVrhbkKPbfHr4mB1qxBS+0ES4LZ1Ew0mF/lLhxNr2mhS//QDX2wKv92ps
B15r41zO55y1k+tkmeBNnFhuEYARkgu18JscQViG3I5DCKQ8j7IZrFr3nIeTHkNKjdpuHwaS2NCC
iWzukoHIq415RDyODXduXzGE5HPI4bHEZ0Rtd+cIBjUfk1SEBFAzONAMymud/KdD4Tu+YES+w3sY
Kqs5voujji7XMfOq5zsqT5Iqid+0qE8uoi78Bmmacgf4FSXywm4Ne7VxhdT7KAEUAUn4HdbvESij
Pmt85CUXLkf+lA/rTQFfcsuRAJbRzy8L5iXNX1tMH6gl1DYh8m+FJXSrObc7n+zXNaKpfyGYSkiR
+0hofDVP0ri5k1qj3ETwQJvtDb15XZ3HU9y9uq8+e34sxA61TM1cTbB3yqwwioITXlRKi7gG0Qtp
A8wLKUSSs2xzCioQhDjLK5IATtAUpRzRAV9QiEiacZCMGpC5kyIJeaAm0pnwXQ2P6UcQXdzOG/46
e1Hm9B+xyqICdfbToXYAJKB9PYNIlYy4tkqSY4mfXfpIYpcsdO1OryPI4PyFqFWvO5ErvjEv0QBf
P1iT8PJ6o3rBHADmuGu9hWe0TLcaD+Y718K1uFBSr4yr58xXuyyGuwPFcyHYJ9RMY2TWyzRY7XF3
iIOv/bABzhkq55gnkSlkYOH2KF72SWHOqr4s3vAkFIMxeCeuTtzWEe4X+uY7rGhIMlN79uI9aVQ/
k3qe5JVzUGzFfap6bSottwU24wFWsBfthXR6218f4HQjWNXDUM+ljKnXxryjwUHJlNWtOxq2FSps
8eqRUZ9/oL6S4WGQGnB3QVIvim6yc/lSv84OLorqwMlmAhJRosP+luZHP5JR1glRIwRRX6hlHz2o
o2ImhWmB4h6ZhPb4urGkrLMlFNFlWp/fdepmffPaBCljaglP8b5Ht3JfAgrPtWs1aS1vBxTHiS+v
+LTe8ibihXLYecciK1FxtZRl3I3AFbrTkgUPNlMyKSyTsDb/zKjeQALP1RL8xX+O2bFlTnwSioBW
lY1/qzxrIO4wDFn2RGn6+2Cogim1XN2iC0S3LECfJ4Ed5OTIq63/dZjpKImXrfh0U01JiPhekzG2
YVffYM5QpXE3b2yCSDH5Qo8cSak2KoQtp3ymd/dtrTdwE37d9aKOEw+PTppkoWU3Cx3DgwU48XRb
cW6BygucOaDbhhER2pRbNDo3hC47IN9l6lZGKX+JepdtsRUo7BhtEzESsjangZsoSKVvpAW+yGzV
EQEHza509ifV6EyTFeXh4jkTw79AQyJXWurEJ5XTdnZD2uY4oR+v42tGuMGHw5q/JmshpeRDdEAI
HGk5Yg8KJp0h/kIggX+wOaUqv56fzOjLOlfWxkD8/5HMN0rXR0Yp/6z1YZAlnM0z+x58RoePwz92
8VrrXBfX0vqw7r/4Hgtd0no0v+f4qW3hDmtuHqzgx4RMK6L8aAF98XRTD2m6p9vBS2XXeMonxRCO
k+mv9KAfCZuFnd0b7zMt6jj1EEMpQ4DIALma83bwkUpbfiqfayyeX1nigZafniewyqfo24/BiAMi
teKHCHijBpW7Zf0VASDBpFsALE7w+WtE/e8HeN8+FepiXgMlTndLmt0BvIv1zGcmpk9+imTciEs8
q+2R3BabB4QD85W7QmVoJyo2Ynv6S079YA1rraL/uPJ1+9R4R2Xmv4njx36wtEad+b1MfK64Sq+/
MrCfwRD/2AxOhFFk1x8oDOTqAieaM+9+Xl1rHxpo6yNZl4QIWFmcLhlnE5Vh4YWqgztBmcCY6lkT
sYBOGlK9j0WYLlTqKTJFzlDM4rq9xKxy1+uSKp42Yn2dXMbooILxvo+7iXBKAnS7FUMlewivLvDl
sgdA5q+CHrKOyJlDImQ/sQUCNL4PShB4Hao5DNvQ6Hf3v1FdkF55aSExIlAVenp/2U6SRiTcxeKX
wF8dDhGTLAQxDDzZfMgK+Ux2oKhP1A1WMmRpt2qdGkIQ6XJ0y7/p/4lIKXR4/GGrhvnDWCHo5p9y
OFWgcNbnYyou6E9JXzytSiFccCKVKQujNznAGyj2GBEwVqE6uG4Uol6Y+H3+7k2hb/LFSanMPtOM
lOFN8VVuuYnLQxj1eamtQMOwSA9jb1eAAWlpUUL8rMZja7KyhClyT+fEGber+ZoWwaYBSV+JE2LS
+rMxsKP3r1s+hYplJIf3PkxTpWzBvXX566RtDEFH2jZeaEQDNNgYIEBvHA8GmUWsXoStV9+8/6LP
8Jua3JrW1Vjbezq5eHFxnMWRjF3sbi2/UEMdcYJIU/ttbXtB4JUKC3hpbJrFZVsBlIZbfaZ5cJfK
v8wkLLJN1IctSHeFPNOFgWXd3nIeQRRRFoHTBl5CEtUdFfln87gnl9J3Q6h/KiGOyfvb2gzjjqzu
TEf79JAqpK2zWOS5bDlTigilWDcPLYfUvBnWN+h/eWgK3+s0hDqrt7pn67VopolOHrTA3lNKsNmp
K7F7ZOtkYRNWJa2mUC2Lo81OxazVJZGq4GnJpqrQMW0vgHWM3nCpmL+nuvYDci8DCHac3FW69oab
2Pb1i+f0Z3EnO1DLao+YR/Kw2qwL9O8PlWQ2R9aFoFO4YBCU7gV1sqBYMHL3okKPqp/NBcKwApxk
t9HCrlfi01FhDqXacXgP18dcwLIS6sieszSLbjziFHCV+xsmZjXv3AkZ1fDUox/YVn+IQdHMRtrD
M3JcrFIk6En9h8QbszWFXptEv+b0QXMxAWFUb1+lp9fv58aPrNFP0qaFfbG9A8v7a/+QIAB6GJcN
4BI22xVWXd6IVLZZYyO7F7/4W3c2xxUXcb6dOlV1ddTMrhQe7XDk+49OmF8eKeS2bpSDWuAf2au1
vjRg2BiexdxFY5qHfwUqCvo/PYjyzbMbay2Y9WfvbDxbtEiMSANHoNWTdqnwF6Q/GFqfNqWiALbO
NsMeT/ic3BkEHTgLiE6tb/hQJj9MSgdmiTkRnyZPeVEerpLlJOcsBclJ5jeC5VYCG/Jz6KmeXFRu
ECYVxxA8BMSUDnvkw4+UNw90Uwrtd414h8OKGr6AzYIl5UiLybqtsbW7KQB/LCQ2wOCvbm6/bPw8
t/vfk0XGkeIkRI2WXhUMXiqAVTx0h8Z2TPaf4p/GS3w8eKCxG0WPB7HsWLv470TeBJS/tUYi4EKz
X2C5VDpvR0sdhkxuVSos0mEDtd/XrRvfOS2HPAuSAFfvHLyiAjC+PErFr5VoXSl67FIyfpNGfCQN
qgtph6jSMk8ykeOjDxPD1/6NU7j4m+FHqFzsnvwV0v4dWvyS2LYB/HXzJqYD1rxReQ9eyy1iLHEt
rmPJN/UQfLya9tOZXEZUBWOZxYEJKphf229I9o/VzCaJP0WaE53C1ZXIDFyCmnNILRP8yTLFKOfU
mzCws3f6w/t6WZBL+oUoehihh1SgLJggdZhC7o6uWXZZUhhjyKzGOFVYw24BnV25wUKevpKpZaE+
u2tiOYO8lNKqKf+HTatV2B6kXUS6fLJjSwPI92Mqta+DhRb9xUxcN4Xd6N4n1TaO5qTSBW2zbjXZ
lvKHSFV+L4OZ869CDOHjeBYm8UMhj9d7vsyscQcYZriaas3B0BDnS7msGgwCLq0mW9bqznQXPTnm
2ZdM7cq8elY7Y8MlY8+zTMiFxMMHL+hzaNKpM1SrMBwVhDlxRXT8ykjA7dURRhvDCUbbbqY2Awss
Cmjlz/KOuCqeQcOIg+CFfebD8taKTmfqcuQ1mqdCkSl0VFFishyjaR7zcF/wk0H4vq8hOkLykoi1
3dqzNftrt/yDsPlpAdlsN9uxZ1DawhIEU+6yOYLM/WNcKz7DkcAFpd68W3K6LnsfObzoafeEecUO
KzKelrU8j3BPVmmZhNA3Z5XSkYdXaBAKqE7pag7iGjBnIWrFzt1j3YkgY4gkpDlmqHYIdwt0KK2v
FUW03hXS9+pi3EVWAY2W4bIAkEo80f3WcI7ZbstUNvWVzr85rgwLRAeO/aE5w+eGR8oSoYR8zdvT
hc5+NZnOV0YxSCcMZJHZMSZdsn/QTuOZmV45eM3NHhV0dmymwVLACGUOYdrtKCZO0njoBHNc6N5+
73r5gckCz4AeEGx3RNUu4yHO96jgaJk4dOOXEmaI70PhTTxci7O94cScKS59YeeqK1BpKrj+5qLT
Z0+JNsovMt3dnbPDHyVUtS56Q0cZc2KSfkW2R++6ilYb3S1VBUYZzwiIdN1kkGDfXnt29kP3VPSj
gQvVLnAO8QeTfd8dSCdOxkQWGhiY7OBLldm10gFxGsrHAjHfd6bF/XXLjWpV9PBqcFDxQvjPfPGA
A/pob5dBFMwuotRlSoDGQpf6d80FzTUWGdyNmVNAOKwKeQbnrSxzF8yuWie1VnWMddSPlNQIRwmM
Rj6zbju6FYUBYhB69DnKwnNiRrny8UM/Wa0eqPRZfhuNem+MqTzn0+litvJPwMJScqsAUd9V+5qh
RP96fGlza6JdO+KKKCCJo+XeEBcdN1j01n0/g4cNYgZ812ivnIEWHydyM7QRKgqh94t+pb3pJFKp
iTjFHhWAvw+rpm77ofR5OxNjjLl6r/7zuzssvNOdHaOVV1Q8PICyuXgh0ovKS1Og8laMctGbEhUw
gVpuvBlpS5DnTNkrp26cf9yv6ZX1nT5l+zOyhs/X5yOnuiWaAyY/G39jYpS/7FzntzSu29ahAYPA
Bgo3Nh6UYwpyx+LNjc3t1c3I1VqGueoYjFu0HXyo3lxDI+zj6Bi/wjaae372IqxRzVj99A6ZY9Wc
3iJSERRxocXubOQ7rMTaVShwNxQpgD/NchEOE5A2RkPL0+yYIjhDCveyiPgC+6qDOypwQqHDAD7h
1N2OZpMuWVzOlH5qmpjrmMeneHniMRTyGekK4yCcpW9bnelSbJMpQEB7KmUuxsZPmzZM71oDQ5a/
1MWyYZY7ERowHeugKl50MMuFmZUjTKYOxXj8zzUTzprLSL/uOnq9tM8resO0Mf3YHItZELcueeQs
UV7CJ32Vf78UBKUiIe/TQuR1BluqJyufrA3WM21j8H2SAgJBHU3OOiBJ83WdZlh4yWLLZVHz1ccs
vDw2FhzTdXV0wwHfs6qVDbrEBnTHMRr7xPeo3QwpXVfGw6mpfdTytA3u0LkIw9unGlbzSu012dPZ
7T2nJSiCdRbDfAJZVHoTsylGrEXe6s+3pQ8XJvsfJUvx8RkpEKryui8DoMooa3wfRv2FT19zPmWw
zOMk28ZQnFbkZ2nv7nh3ahCKeAw/BrVbTW9xJpo6Tm6u5t5Sk1ROMTJvNl/WS8c/4e1b58AloaYz
PGxIp7Fr5YuHNDtivVsbP3CrhUBZnwlok+wU72Hu0xJSonvT0S862jouxfJx1NG6DbHPi3WXo44n
IxoJkItkVTRgeg78EeuJ/U0kC2MrDpLLubbbBrXiUAYSmbGbqAaHvTHuRCkb84zIMiuJdl7ay7Kc
yaN3G5oXBGCaiXFSotfr9OLFYgfT0TcI5dwEZUrZRJIfLOIYQ6ccx2OXdkazWBoxo+AK1P6T63ja
CxjC7rQbcoFL+Ur7gO7cspnKvW7u54tGPODPJOx1+t4MnpTA8v6ZZmbcNKNrdQJg1T2xTq6+5rXt
2pSRQ+gTDjiAYcVdK+lPHXAf47r3f3e/fsGvUw2P/ZmQRLf2Dbu7ocPHUnkJ68fzuARriWkWxRZm
7tJaULQ1BXxPzRq89zDbAbIDe42bHezb8LUZH6TtcGjns8bjQ0ALPH12vFYyrUy7nx/ApVqOmehq
9qDrdGkdKEq/k0PBRLjmPYwEsyNATJAocCwJOHrpm0MutmDnDmIpJsL9p7rJxtYsgLkmmk4Oa/ti
1h2Fe0c7cHAo2myaeUI6V1tVpDXEnX7cgZNpGi4efGg2GUc9cnpsefK/EHqzGKYeCjHA9nRfKtTF
/MxXt8Ca7AsSePZ5HpJlyaF6qfjM2bbgeNtdXfsar0NtA9ezusDkutLP65+ssAR36QZQjhMTIbKO
jKvhjU4zqkzcbX/jPR3OQrA+Uzqzegn+shBOMCY3h/vWihvdcN1LK4Sxc2F5x2eFwIlRKeSwUbhq
imN4fXeV7irgvqJjl/1lMpS4S1W4CPaElbyEilejUS7f3Qbhb3Qp/q8n8hVwq78u/ENWLYE/5wvk
X9ZLpdEU2u5yjL/w8omq6s7gCo6kyXeAxZnTDdnqSYluS+G+oLHKKLNCfGDHGOTBS/gpGW8ydsZb
9MwgKzCXiCUExJ6JdFPGnv6wmF3/iRbO7mEsg/kc/wtuf6ZwjRDK+Zm8uKNauN458fsFWDBj2ixG
YxoWB+/frhbEgvi4eC7CcaTlosT6yPmG0fctdjLgVrGkYAmu4KAvfBq5D/X+ARXf1mWkEem8j7hK
OWFl0xgmqZCE5vzZEod55/+lP8bw4nl3eScGi9Q9+3iy8NE+V5vPH9kTOGsV8oQAk0FtqcBRrygX
19UrZx+dYdJz8JTY1RYnpUALp2DHGUV8Xx33yiK1bM/TPhRA8XNqbAiED5juUqKgCHVjX9D2mUJK
yXIIShD0Ocmuv5/g6Et775SDtf2vE66Ajg0zSDOeTW3HyBFX22XW3aThWFSNuHCyYluMO0z5LHcn
ldodsFwoelRyln57M3z1M19Q29n2Yj/WuGsLDhtmwO2dBm3HH2KJkJkchmbaQJGYGxvuO22Mkn2I
ZF/UXkW8jbd5jcnnA1JAI5cIhR8Oib+UsyDhzx/oT33quWGkRwT0dIZo5VO6jKMP6WiOkLq4pbQk
X+a0NR2jCo24fQnW/L531pQpyeoQzKw0tMZSrAQZSSU8mpKIOdvfBX/hkoHRw4ttP9kDxgtBemaY
eZY8ojWh2xDVK6IhjY/KRZYtsj59l1mU2sQWXRORE8mwYyT6dIzyFHeRvFnCI1CimotuJXzHgq/p
DvKNtwBaY8uwfMZaNpkt3iD5nTXvtpVEVDYxaJHrsRuIKZ/S98Do9PlZj8/gYuAqINt9IT0LfpTS
T6W9y2hpJa7nI2OihsI86TFZuBzn5GugKLFWBfZpK+qGYkdXwfHw1xkP48eum4/VROp++UPGF4tA
Yq09GD4hUGDC5whtOzUD/pLINX7jJW2uvBUJBbbEK/1m371Y0Ny6o8jLjU/lwQOMnwt64x9VjVdA
CS797jiMyTwVop4Nd2bofUbUjn1gQm0g4DZDhVHPgQwR5/z2MH5hmr0/4/ewvpWWkaEamMgUnz5Q
pKmTQxrS2TRrOXCpn7vCFTrhtwC+2HJRDiCbcycU468czt2f70VLf1yJHHJ7ZIfim0ft8pXhiO1S
02qr2BEd3kJKGEz9kgM9rkFJG2bmkYfTZxfifre9gtydPEyj/nkqVwJboK0Qb7O0b5YoJt4yEpNr
C1GJ7oQEFHoPW+7x3AeAwMmAgk/++oeFi/uZKXGd6JGSqxnTYb9Q/mH67BPeXNgJl/nuo/hqstwE
CtX1sGZNBhs97TdO4mW7px79+nC94YADnVsrO95lYzM35hhjnKp1iUV0inPWpRnrTA1dMwLl26b7
ghdrIJBSG9ahv4zo7PNN9qQLt5w8vbwueYmE1kZBBkTL1H5rwYvVOicSxMvWYZUasz1SOof6lhAn
N7/5UaCLPrLCSwrw9/nZJGMqL9jxyRNtW+2hjj1DKZUCMPf7cauWOyVaCKKzsUyjBP15VbXJK6gQ
nfplXhp+G/n+ZErykSfvJN+qW8t3dM6hyHOn3gYRKpMeLirBQUZuaGUmAVUN+OfTe/IbtLvpYfwL
2qRCs10bqQS9Y0Z2+W0azfHvpgyqjTcZhMJeN/i85bvLFPHkhWdZpdxRIP9qjDMA3CI/cUzk3GjT
W70h/wkgAHlqrTCc0G2O/yWMOna1KhvKdDkqO1dM6xYvC94yxgiskk0awyKxitnp0M3oYhh0zQOG
IPJJKIiHTtudXrjtl7ZDz80qOf570V/dL1Ri0TPRyTBMeG3faz1zFrukJNQagU0Wu79u1AtCpV0I
gxiQ+uO4GNBDq+ZNwYEhmtqzCWruA9aM3jfz6eZ9ALV6/TXaTl280HWPPGacyUrGlZTB7/GrldmO
rcpNAlY2cbsVHcepu5rINBfh0oOwvVR2vMQ0an3C6mJl0wAUMYCr9/DJ1DYTYNRt5qVBaZL+dmbp
8VUuNlQKdHcdqaIc40Dhd+V0dk0N/SI3543crELBGoOSrjYGQcsBZuKMHXNn7qPg0nLy5xI/xkBI
uKMtbv/QOPMr2WLkG7CGAXECTR1otEvQFWcn9Ge10ZMD6rV0iDf8f1jHkHiNvMEP9PhOFivJi0oK
K8UOq54Q82DujdRUjJyhcFksxyRUF4NTLysLbAnpmOU1kvUlTrkfQOSmqoMr+L+eMt15F5rj/SgM
V2Y8yC1019aIlGECgV27zZgOHlSC/O4hYQg28kMAuO9Jg9p3X1+FAhVG1KK7/u2rpazHbzK/6sGh
4TeXg8NKKlCKjRrBafpkV/DZVkA83rrsorhuXM687Q5HvQ/PUWsZgGrc4lFiorIORwppKvjiUgzz
wWmWQtoFUUHgZ+r440MZrM+icACI+0AmVicaYyopK+fjoGxO8Iw92RTretxCVH3xHz69hMx7f/a+
XEufdauRr1LSMf6E1A8K+viW2D5cYP/ewFQEfvBWX6WcYz4uYwMuOsLiBR/ZQVAiTLHRNrpn0eRK
8aRnoaERWesHs7VUvxiJsRg+MxyNWBx9F2BxACP7wMaY4ITMV/jrWmawxxPnVyxl/PKpzCsMjFmz
5XiXPwqYNT5ul610dwEWoRWGKoULIIkUC7W5vmB7IDvHJQd4b2/ZWbaFbPksqy7AFuGZCBfe7s75
7JzHQllAegCpu2N1BnmR0bdDwb3QiUCN042GanvcQSUS1IUY8CdXAj38fXLcRFsa9INSFBU2e5jA
li+lBo0ZRSiciOmjwKPISfkLE+r33WOnhOGhMmWe3ZHP81SlUQIIEDnAucsizj2iOAq6gHSIjg5Y
dzdS2UoUXjCBe72Os9vpLTcfF3FHAeun1/8cBDmmemrZs1+8svZxbYkP37/WtmzoeVOZOkwrA7yW
DrT2pGsKEPWEn+uIdD+1Wmz5ewIftShq7oK5ZD+ySGlEbEzqivBvD2gryqguF6Fy/WEiLN1iwmBz
WBYmIDB7m2N62yQpy45TueuznlYImIhk8ItT8CQOzkqffW80tUj9U2eA6MoiY5THqWpxEw/kqB4C
rulUJYM4Wg+G5IArGGfuQfqrcwLGCkodw8Qrg5vTenKtWRfqs3XLl8Qs+t2nbSOrMNu/wSbYITun
jYoLwWqWEkFHQltpAWyK91LECgrhMPMxkQ/TuSpND4ybnNiaB2HCyrd45kQ8T1sZyATgC6U1JqGu
wxo3WRdPLnUKja26TP7V+HcGD8xYhLIAwCxY/EB/0+uOllkDMJKZz6PkKEkP2eT9kj3/ImHxyL4l
XJx4Z55BmneqQ8qoKlmuwDUn98XoZ5lMJJ2xq5LIVqWp5/0xbsC8BXIiC0usI/hvOA0Pq0YnSrVW
ugk2ebBYlwB2JfSOZxCI/hSitqTwKfb4lROe9N1fL3m9R7cFgHco3osnCxfGVXSKqijnEqN/o4nz
iQeTFCL4GXlzQb+jDLAbx3+qH8idcC7XKCEQ/+NJTUuO5KL2VxR4M4NuobfwxY59/JpzpJKRQwAV
GRb2MRVQ0yDjiOF3CCju1Itm6UWzU4YmydoGXFB+O15VD0p43miTmiluFajvflCgz4g5EXotgAm8
zTdr+FJjFSlEF17gtUWJvv1u5v5kRtBOhdY4ImVID5wdGkLBKiu/Towl4xoqmriLWeJLPGz0o4SM
9S1S0ZJRdn7guZfvlmndcazuB8knN1npw7Wgh1OyB/8gjgfu2KD70GKtaQBd3Yu1l3z/NsnRPmKo
uyx7Pv1XaeCAgmIwgYCobe/X1OazDWX8LTbFv0H8oso5swrG8b17mywOfu/hRC/ncglZmXju//vi
U7yz08JQsfKffZbOborfwMWqBjV/PQ5d03ozpHwsSc9yZAsu7r1kA8qSIVuzPOgjdbEfmR+wAfnY
NJHxub7j0EdxhFIEnmerCWn3eXce9AYhnbjBCKIx0Sc0AquJPlnWC8W6dFlchZxT3029sA3qqXxC
jjbmDo71B1zW+XLPNqKsDM/SZOAWUUq7yDzjMEJ1fl63tm0mf6SxiUK3vqqJFEfH8rJH/95Jqfai
au6p4Bk+DvAjUbMY2gfnc56L7WXSIsCvFJQFHnZ5G7/UcSo5zF6Ae+v1qHGphrUErbh4Nru4K/JD
W5eGFL2YSSCtPFQ+sSWmIgTKnxPMrsjomoHQswzoBszcShKFQnIqXJHguP4W8M5t2dYxNu8m9CtL
cpErTqOjVMG1vbXV2C/wkZ42rTXebfK+NpX9KcERk3OWJ+6hpRGwYNwXf8uliV6nxfgYku5eeUfx
DPEKHFyIRNBG5QgYoscUVEEUcMzOdnUgLQ3r4ArAQcwy/q3BIKf4wLa47WHKXUWJDSi7M1dNjNoZ
m8QRLiwsNqTg8f/T9Sq6e/V/pAlv+/vlRZ1qAXYBFEvU0Jcezi8uJ15mzS0SYyTIOE5JLFggolPO
8PBOd/iCFJlaVpQjkQAJ3IwRCPRZ6Wgmm8uyKnQOQ7glWSaGS3wNkLHgW2eMwq8F9w9xLow4Qdbp
BPCkCj/UiJmQ/i67Q2eVoF033liBCDKXweIjvygqFvGpFZH4lafttl7FFMdr674ZKmkDnaJl6zT3
0Lko6EDo90gVfcx0iq0Rb0m8oti4AaSe2Qa0bRte54/5TajP/yZK5P58LhtgobYwj4LSFEBtDpcA
9Fl18JNpX+2deyGgvgNEcOPe7LRNNUEVU2HSdasngpQhQyLdHBRk3tc2V9XP3X7QxacYCehWMrBH
nid4M/4T/OttuhwVy2WYEx/0ggZk2LwTCp6FIzBpxvMPshNRb7PmfOXFQufrWAFxMn0dC1ZeCpil
PG104fhudb0XpxHozMknTKM2oj4PorJr0V+RjbL+cd3tr8esTN5t+TXMdwZyI/40A07mkZYfX5LP
0X5TW4AG5ISkKfek9oYdQpoLLHRBp1wXMY/Hc1VAJLo0SDc38GFXlIQRh+a9okE7XDPNCM6eSueb
+YU89AQoeiQZwu8U3+sIPSE+Mi0WIU5eeN3Agjy00FbRtGx59Mmy4d3wCNYCNOYRHhjPsOD7jG96
DgeTM8OO6OkpWorHYOEu4KZ81TFtsEA2VOmidJfZVLDBzVPovEtVBhEP6/TlL07FgD5Gix0WSqcj
nViUzAk+YtLW4YU5PQF8pxxC26O21bnQ7To6T3WXmgjgOozJ50OmobkjF9kGPAD4/ovC2HwjtrKF
ZYnWqmuJpr45BIhT5vTJbZ/lVFrERN4TZxLq2Teu2mTNMU4QW/a/etC/pd+l7skMm+ziP2PjWc5j
2Iwg+4V2JlXySMMGwTWmQHcMecZ4I1h3MLm8QiPc1dprUfpHU0xZ0NfxeNlnLh/FaFkPqaz7sriv
Fmh+TzqPcGiTrCgY4jH1k5BsnIQwRNf16uJNMyCa/cl/Q4AQjKvR4ULaF7CUIzEs3fN03mHLOHmU
pV1VMccj3Xh150M7095Lw3ROBdi/jGvqo+xw7mMogeWpbbrK9hDG6RTsW7TmsfiNkpTGJXvVtzFo
7lb3B+FFZZOJRNmWCsmYtgMNZBoSlJjdqJdZLXdKfKsCe3VefbervjWFb8qp6G30oZdfecUqnxhA
T3LKQtK5Qv9JnHuBnFYcsw8MJiEnJHKM8LWaG8EOvjRc5gwtC87mZhK3asVRfF3uy4bH0IF/vTON
J8rNDfAAIHdcHKo/c5QdBqlsKdEW2hqCYLlsptG5AuLti34a/lXLv/TMeLGiU3B97SizQATx2pz3
qGC1otQRd1GoJmmR4qv3h26d+SoVMTPyl4qMVoHfEqc/lZJHjKDuKA6+On6pROHEKNUPi7wBBnRp
TwDHgJvM7Gd+0YIUtfOOaTTX88v/X8ULGYe6cs++3hvCEn9F+Fl9oT00o59PWh40yH0exTjEn9pD
dwct1x1nUU34iXJaDnD9N74g2E0KX+LXAiasxODZr48WOV+Dsgsbn1CqENDUSoj2EFdvryLa0SSS
40Q358146HpFuoBbGfur7NtYwgyvPZ8ea10N9nlQJNG51r0tBZ6cbTNS3F+wTsfG7Rcbb1LsLFxP
72aIdaCIxXgHoan1mVD7yJget3X+P76s91AVMssXt774cdnfAXDB0iqRyUTnFdJ1HCiGmPbMM/07
22NyOObNovbxL0SovtISjY+YvbE+aGQYTUP2U5s7eJCIwaIPtw7M8fxG+Vgpx2wE8HgL3cNjuofR
cSQK6qVdHw7W95Ou0SJ3WMpqqUGZyes8hJ+mcQ7Fpc7bs397O05q8/Hv7hk1PRGRCBg58R2St+4i
Q0ReJxszEqSVmsyYG7sBwy8ga4+7dR37jpg/zyiYg4eVqsKetKgoZMSmERVQSWBHk2jteZnMv9xh
5OS76X6ol6J1BoDFLLmRh8CnSgPogk3eIu6O5w4kEKJqvAx37hmEjolmn7A+Krk9oedTAFLMJETn
dmns2EBu6Nj2sD/zgpYvd1Wkf51OQVuvrhLdDIG2t6GZDC/pB8pIdxf8HJFTwvy1h5nA7SdQZDM6
yPWfd1E8hY/YnkcsI6yxJwiOIULg3zat1zPXVNZeSgu65DXt/aO0dgBMgZsjmwk/KNeawDRNYhzl
gC3HWue8wr4ImDJ2zNmvcjMunqA5OKf98unOZ4HFjixvdM71c4Ok5G7j15yRxC9gOEQ4Fvz20znF
Gu8FMuMoYw9TCZhYofa82grM9PBnY/ysKX4CTnNHqSsMfKOBn9P7WH3CxLyKWbolLNjcIVwe02oc
AXILZVcNdXvtbt4MbdevimnRwQlVNsVskg7T+B5kwv3luHR+Ko0lPyrOv4kp7RpoH+VXY8gV/wlO
KPx721z2d2Fdw6E+fmr+vIpUt9n6Kw2ipVtUZQje4ik+l685OinnEuLiuchLrfnWiKnSTBLYcw8i
KVdKweqTysCx3PePY+PoVOdbCFgORzM7sCu6UpGHWsy3kU70bJFsDFdqV9dHj79fQ/uvRHbOSzEr
yrJlpX5EiXGcYd5HcJ7zP30UAGqV/7ZaWqOQ1YFHsTsoi6Ug8nphRFcToFqUdd/BFrDbriIXd3g4
3UVXQGhXmN+t/mRladgZHL/XE4+w/DHS7aLY9PT2fZ4EeSUlfDUahSHFjI+AafQvxb/fbAeupO91
ZLre6FnddCvx/iQwNOF8G+HC9dnhBmvoHR+R+NPkbCrvRbQf3O2uW9Ejmbraevn7sGxWHc1MHpon
1ZIpHotYV3tJQv1L6REcIxC5KqHUV7awRC0xG7O+oXn2R3c7RI30fcuOiPHCJvgzcKHWCiz/vCyD
aJZeKlXqgF1e//y714IxqDFUQ5QlyI0ABE1DCXpkTcMQf6pp3LQxtaWOJN/95vZV+msdEhoWaMHY
EXEMZ8noHLzm8JjwLXO/EIqwZgnHFWBEzTGPMEl1uEJUjbH8lx8OWMPuxD8VD9KW+cqzIuZsKWOn
dAfrZQhsIOvy9mNfU8uFfXh9hflplSO5tOAgkAJuV5uZYAAo0USMMBVGXCzu8XAY66ExMeDMNlos
nljf/fKYrsb08BdqrDl3ZoLW8BPpD+rfMBUXbKHM1wl+4ioaIRRqOsytFytBvdDvPcVr3CmGA7uP
o7VucN8+14RgUVgcvLLNume4FNXNmytsDxC2JUw9OPW66K053rhwjqA//hMOwP6ZDuaWawmUQKPd
POTutkEsA1TP02XETRN58oP/7yI9JE3Ysp3HzVS9KA9EPl4j0hLL6LWMelIm9+0eVjzbnaZOeQA2
CMh+wv5j9AMJsXX2zFwo4TugpvygfSau8m5hotvbTyj0L4mjjonBAbDk1MV6EPnuMLDnW1v5Gjll
Y+fy8+yiSMm1QmJcLyXzDvSCiG2BSu3DJmccKU5KH3XKuGabtxdQGQQSH3H17E0VFILxLBYe/fjr
iKtvzOkKo5FL5VfZBihMGhUanAY7zvw0/x1F+YgRnUNP23z/A2y8hlFxBehA5rj/sL9+xVZCkTcZ
S2SvvZWY0FKEIXWUcVygHWBEorINSzqfy2iaVJD1DAcox9a8VdWinJqrChOWcjV+WQaMOJVAbygI
ZC/nysRkjf4tJVq4B/Ga1YyjR1R5P9sdEiS/hRlAY+o6t2AtXzFwO/z3vSFCkGyqysdAM/vIt+pP
ACuCnq7X3i0rLbK/SrGp9tdMBQJM1xqbEu2ZgAoTCdC99d4wj4/cZNrhfv350bn1Kij0QLBtHW82
W+Xae+VwGeZ0tcCF1oNBzttEXJga5dvEJRgh6SRLdlfBlx/4iHmtrfn5gK18TT5A3sDrRiMJN7IL
SHjCmZ0Q+jXsn4MtubnH6wbjAbjiG5J7fpWGPhhgEBVFoRPy2W6n2rE6nfdK9SvFIAjj8SLXnhsW
Wg1h0jjU4p/tmtHLIxQrD7zGt/8MuIjpmRezQPQc8rpMLRKizCa3np5K38ewrZG2rJ8p4JZvQ00r
AJpcvfwdfMfxHuv70+kTMMLUdKC2IDpi8VaK2Lk59+pCZ+6VCO0HbIy/JAimDkvnq18VCsOWvR1z
rwgKHlio2O9TIpmlLUIVBSxngaBwXu0+SmWB0V+7A9wXy4Sy5ahImkk0xvTyaa3esbgEO9/RqMDV
kLQvLkwSPAeDBrhjuoAmXX91gqsiR/b8QN4dm8aTqJWQBTKeBlDsr2pC7n52YiVdyd9UWGPJoBSh
7AGoILcWlOMBCQtQxGhCcofYjMrDn2wzSSZORmmjKwGCmmTIqXhmmo4PriVP14VhICQ+1VeOdHy/
OWqxB86GtjOWBXgRdW9JsOfMZF2h+sMbxhmYWG+TCUqBarROi76BMs8BWwH6I3hzj/lAk5JaUoE5
PhIa/pDjyjDne+ot5e9MNVfj4B49CBDkeKNRcIu73egM4nc60w3Zn6VWxRY+30u66btL34WsB0dP
ZSoZ6M0qTdqA+K4WV2bZzPxw9Z4HBNLAHky6z9UdL56h2bjczxCT3po8O0yqvUBN11SkaqEgmaEb
pW5IlkSJyvb1sp0nWv7F+XAeWlKvmTrltgu0ToYjVcINR2tV/N6lqrqytrMPOX2Av1ha0/VulCW1
vwzOhTSNWDcuFaVDsBWMjaq6ZHG4XhOJcqrR3RS5b3A1mzNbDt78vk8sw0RO0hcRydyZcB+SWerC
yOruHLvdsOfXi4kvbl6fJJdio6shBhcmOVcq2PKhYOOC6FNNJn7rwfRlFXBB5Rl7y0QIl7uqZ1Rg
QG72Y3yxQZz0CJ2fyJKnJCcmvrB5X9+62ErI+lWsrSRA55gYji6a2OasoY4OCcQtxpw0lLN++5qS
7FLfApjfRQd9/+Osms61N92RCE2x4fWQHnJDY0C2f3EvWHWL6Y7PjL16k8QZPayH8Ye0hVEN/9ly
ML7ehptmFb04pWvjHbkH6b96oy7eOL5BzFLVQdkRwUWCOvHmvMzixuVmMRsL0SdgmmZ9ZUpWYB/f
xPmYVfi6hg7H7cildQJFuz9mLzzNnwDAdaIBik7NTDUoLn5DU0ISyyALFe5v1yEVm8IifrTtVOul
1Q/mZwP/jjX8PLhYHdQSO4L7ovsAxMrZAz2/36RZBADcNoueLUR9TD2/vrzZiYgHyk08Pq+StG9w
HPFvxo4e+EPYGlsO0hs+V0m7VwmY4apmYDxP7Nwj6ae2tj19J6VzTCrgbzvzY7mPNCkNdBuLly2E
fuUuDtmm8u8/qMNCFdn89HXwiAvHSALjmqjWH8uo5+aKbh/7G3VpX60zRDb1xDGIRUx7XS9/hzJP
oW3Hm7i1PwPohut3uX1LX1qnRL/Q8lZzlKl9AEl1+u86debY0Z7PgpeORNIjVgfbu7GIs20uYiTW
MmflGumx5pYURZ2oMepd7TI+qQhh8CBtquAE2ifU64E1z4D0WYLdVdx8ZJJprNnva/cyJVTDLt/M
b4cRI5GPf326rx77nkY843HULNxYFQzFN0T+yTDr6tX2CBUhHTkJwec5N9xrPWmlqnRD/kYbYAZG
JVsjGaiYtlK2jnKzmO0jPy2jB/Owbz9VAIZSb1DjP/+fv3tXNEbloO6TayTpmx1ULKp8WJvArKzA
ZPlkXSHXe880r4lxBeL6AGlV+XnOVLRraiLgA/jgkOpldzvP/3FoQLjqSrXdu/dW7IyoaA60T4wI
xvFuZa1ZDr7u6hkXKfhZGlzQLbLArZxm7AH7IhAadk4RFWDhuZt2JRXSwVOX1lhJ+JuTdA7y+dwy
rWzboRqNy1aERa/38oV1MzdkXXPrWllIxFIZ0Fy6OOCvokMTlx/+EnzjMZh0a9BojXw9IdprULNv
q+/LBcOWNxDgXm/uLIM37Zmyl1VLP2vrRE7i8FB3HhYfD8iXQLacdgCTjQKk/ex/88bGG5hyyDKF
Zid90n+40V48mpmjlm4+kXf40BYgROf+CrKEk7VmN39harL51dbNUoC5wfovYRkFI3ueAYEWR1Td
97DpOVooapRCRvqb60TiT8GMQh9hXH7hNp1PZuS7PNeCYeYC17mJW4zFPUSz/JQdJqvzlcxkmSgx
Zy0JKpowwEy0lVv/23JrOkGtpvI34ZjOSQnq2J+PzR1+ibMnq8d1OK1atXF0zQP3gRsgD2K5xqPu
TPe9dbe2CytiBuWSDKsMaRDhwCHHzW6JJgJ4KSBABToGWDBO/Y+3KEKjCHEtkjSJX8aYxTFQnuMQ
PxpYvu+8JeTDEPql8A6e/Pz2YllfO35aqlI1+VDKGiax8btu65S/G6rKUIS4QAbfyk4XM7+cZrGg
Wwx2hOR40lNOjjNq2OXh8Sywp0SXwfA7mfBAN2miEMboRFRSga2SLoW+CcA8OvDKYYwAnkYncmrV
U0gJS/CLkqPIxTVwKnbVMXvP48oGgNwRP97kOg9RojlXlrr4EnAtuUF2kYeTfcQBKTOahDzaQofK
+onTX26yFJ9Sg0c9gEL5bFEeG3w4INp7s/9BxXVepHCCvgpKuZLMro/83tA2D3B9QC8hOnpkvj87
CwUm0QhSgJX1DvvSI3S5st8Unj8XM9gsnqFvvuFRTtjFzpmVgJArewNYZjBX78cKvGjYFWqTOCGI
kopDGhC/E+xIPZfvIZmXjy9A7670BY3c1oRAb0LhUsJIGjX66psLkzxJBpYJZGBnof1HQttCaceq
TJJU0prwkXfkXJnGze9ei1m1NHTTI1+8A9/xOiQ4MbexkiKwpemEsFlGzcJCTIVfIMru9VDyuKx5
Sji4JI6Tv04s+15feMdTlby2Z8Wb2W4FhTOJN44iwChlcGj5Sh9ZJkEkXi+81gWbAr4h6f2ukR0K
Az/8BxjZdNsctmOB7ICQDN9xb5tw9qX4q6z/Wof/cPSSYRrAEgNzUL0Tn5UkrZgWP0G8l51PpHEw
rv7WXRmu3A2ERLONDZkhZ6dLTYhDrXdfVwl2xoqFwnehV75UDU2r17n9tvTKv8Y1KdD5rIQGDea2
smhFFtkBOmK6x2hPNgUOGJd15x5nEaHdYq4T0eu2yPF/X3bH5YASQBC1sTf1A/+WBSsWG9Rggq8q
KxjZ4QkDX5NofxKjnytCtoVIKLb1aIW8rdRIQ+kpa65dq7qfBD3u84MPZbRL09qMmzyq4U2QaKZZ
niVdfyRdf5Ak1fwX1GHc+EtdKvv5n448kmWfNLHOc1au9PCOxcdXydTp7TwNbPQnX26Mb/7DdWce
MKskq6rjzE/fyqkyNhi1xD+/uLAyNxAz5iUaOcPZ/0a327xNMeYUr8zFbnUDYUplSpVE02vySbj7
xGdxzCJgOBWY0DB+wyUCv/Juh/ecfKhs0pipY61ONO1gPdw8lNTOxCSgCPRiVLuHE4uKCulJpQ2I
Db/aVlQ0EJr7DfkVFq2h+h6s9TM5R2WUVlWHHg/UW2cahbqmr6J/CIMRB+MTZNekLg5DID94Puts
gIL0oXKuTx+7McgIi2OWxDTTlvHxzNDeufDgugsSrVIIx2TeAVk/e9qe/v9VQvyUawO2Gz5MNKSU
m/bEj2DgTrN3VitpzcXdniGKl4Yzn9ENW3q1NaVXSse+La9Urqg3vC+C/1cSqKuWBW8NbSuY9rzj
Izs5NmaDc+O+mC53pzcawGXmJBPcSmuzVbLJBSzW0umZQ6T286c9bj5QQLuxjF6u87O1GkeCN/cn
haZuV/b/aQXq2CSYAWVjD3Iro9FZOtAd01TDWiGz32XEUb33f+2P1g7Opxx/z2cjYr3rNhphzfk1
MYhp1h0NBVcj1au6toiNUgcLI+9YjC+W/CXxO5naflHS58TU3WvAnCzpZVS6lPhsuT3ipSdyuUCy
rHfffMUAK/9mX6jLMMtzddsDW4ZXvx2ZZtX9PTJh8H+zfSBOZOqEyKZl3js/g2sB9f9F3LoWlFZ4
A+2QceIhcrr/dtSPE3iAiWVkBJAIFQrLxDX2Lfv4N56+cjqLtOrYnbEq8MAxT8UJv0WDO+ZXZyRs
MeoNz14Ed5NIqCQjgWkRkud9OzKIZB+RjWG5NKPL3/Mp2EtRrGzLstjQAHs6ivcZvGewIK+L3r7r
fIcJJ6FjSkoMUT0H0tQY2oB78c0T+jm2sP5ywPeQR/LGp/CEkFi+9qJCoCCpkgoZhcG6kglDCDn9
qbXTVd2tnrPa/biZIwHhXRMKSatE8ImN3wsxS4t7He2ePFALCV8BnbwdavJU9dkx9nS+Dwd7SMBy
WGOFn3SaxkZvIoTjwKnpioOzqY5U98JLvCNi1QOiKPAp2b6n6e/QPTUXjQJ7o1JaQDqWrZ8wsa16
FXeA7K/3PsdQYVc5fJ0uxZtfRFCvvSWbCklt9PJ9aCOxhpUpurLpoPXZ3Qsiqp7Ljb4Vzvb+nNhh
P5uvsJPVygoX7eWBobq9uS5vDmbaOXhYLhpU7mGDPg13pjeAjQD3XZrAM5usrQwEYtOkuoNezPbQ
FpJXQ3WEaeFa9Fxu0Jy3VwCuC/wRNcZxPFmYymQx8r3n1p82+1ls7OruqefNw8cgdCXCuQoj+Z49
OC57fgBwyhJp8KmnMAP7iEmzoi+UDqs4N/fJKeCHVwmsr5nF8ifOEFXAZTwq71AAagMbG6KSUIH3
D4W0P3FjmcF29zG06h2idyCCnvNzg+YEtPAz+Ugl6cAoO8xcmkQ90IFcSHG8cAhJgjPDhAJDqd55
nHLdHvPvQzSzh9fpvJpwAmZv9XFuC4f74JzkWBkwDnvZqkwHF2L6A7N/lvnlL80/uk6w0jJDdkol
yVbbtr2A4XckaNhNS0QWHGTP6mBPcSsn4KH+mJqEOxA6EMi194W0Pgy3d8lHQ1VgdFliuiS1kLOC
tavOOmvbaL4/NnLZW8nSqvJn66w9rzPMm/uurxnbNHrR2sTwHf5n4gKTnvrAIuzLvL2jE5xaqP1s
hbQpui0gIkAmq576ohyMQSBnR9T9z+0puIEYrku0yX1PWTBRDl/yShWSzgx/ktwx5f4ymLaKPC/S
c6ykSDsKGJN/kezfNmQVBW0V0nIO1g7+m8B5mnhqv8IMN7ub6Ay6fls5Tnhdw9c/KfPXxHg6p5ls
sY3COTHhqJbdzdAP8BT0sENSjCWtlWHUJqy30bhxC5+vQDSKzv0C8IilyhOFNnA1820pjloZMVxv
2/FkDsJPJbdSuCBJIp3gzzlhQekrNFPLoHfMRQUgtr78vRqj05rkpm1OKMv294M+XwbbGtasD1/W
n2DpP5FtYmyF0kL087/167AlETDuUP1wGvSKNgCmemijW0g/GFPOUFWOoQlpB0wDhuDzkpuJa1fl
n3hXndCuGi47HUHs4sdrB2ZcJgJ+ES5u2BQZSL16/64CZT70MsE46/ueyLn7rVnDjE4u4DCq9cHM
R5cu3MwdrNwfspS3UP1Cvny6ebuZQxxQ1tCmjPh0PCGfBWcuavUN1QP0V/CCGXKzdTCWWyQoX7xL
8ol934PZvORl6xTgrSg67KIouz6ma1e2nrmhpKiUvFw27BbInGs8nRDwc8DG8KYT1hK48eNDD7VS
KIFe9/fp9L+EdDMGM5lUXzBIAa0ZUS+AbX4caqHXADsLNN+StVE1NAZa5UH1Cf3FJd+XyS0Ro7Lh
g+bK1EEs7e47hBrYJ7e8KOqvNE4yR9hphZCiDP+krSY3vb/8xX1yvngKC1JukK6lFrEZ/q1RFi0b
77xe+/Gdj2YJ8TZaig6S9EJHpwpr/JdawIKAKbC7qTMD43shsDwchYUpgaUojzJagWhbtARzgGuX
4DKahqwtVOtG3b9YDj1c+nZc8PcTXgp/nvnwsZr+9WzDA72130AUz7gkt8ypPRqJIiVQV+3H2mIg
JAyBgwVixo5n53vd6P4PSqaEBs2yTZ7yeQsw83+rEQMNTNqXV6TSlgpwUpuutZQeJJ5yMm4uPrQl
y7pttQgxgcsqGg+Of7T2omeo3uIjSREYgDXKwlPz2Hlb7yEQatqQ6ULfQXTxyXnzwxq1EIhBc2zg
oknOgp9MosJtJe67v0CE/na7EfhIgZ3gcs7EWUJdlevMBSZoczSY36jO5LLWXf7QJSoeEtYiwSLc
jseJydvqkYaQzWqWLHR/QpbXshiqgTFXx1+1XJzlh65vTUxlbXmmskWXk8NOGig1ByP+Zut14xYD
NPwqvaChDSnY+L3eWG8YLIb+9DJfnt3niZilQnXk6B1TnZkBThP4BCzjlkfiDwyNbEr9Ogt0syKp
O2RZ+B0bTDDV2x/iU87ZQxmLJcgFy2vruoTup3LQ4fL0+3nc0Nx7S+5D/OCVtuGLCftKigFji4YO
N3EQRNmfZLsHQM4ur6sObnCjrYmmblkd3cgwL4/vB79uJOhjFnwdZfiy3A5zp9iidPBf/TQRshf1
PXzftWMxgFxpqnJCe5U56tIaeXtSDk9Tj3d8MhJ49TppICclhRbBODEAzXQ1hMJvG9OmK1cxtvsT
typj6KZxI5MBWHW79WV3K2SPbiIwv5UeDWGt2EuyrvX4/WvA5zYxiSluysTO+M9VhdnaVJlAx6WO
ZwlOPoCidXT+l36jUM12pJNhsX23WDQUV7idWZAhtpE3ubzQ8TqA3znbd2Rfzt42lgE3MwAb6iq+
Q1ie8McD836nERd+i18A7+BNehf+a8FHmYNL+okiQz+jHd1kfoKYSHyD6LBPD5g6XVwp7UzXqLmI
EBReGJyyYzVnZNtdMSagvBWmJ74SQmUCchhus62C6GZPIcXQ9MzgM2lR3nEPFElWOLRbuuhh7fFJ
shdf6CJ9a/AEsD+iAd8UX8Jea3gc5rXcAjmq6/Eg5TTpe+PaQgcTS9NSXgIdK5v5+BiKnm3FIPAP
6zFa1ebcV4O8Ec7MMgfiSXFioj0fej94i+A8lGIYdQ0jTS0wuhT2c5fmCrP+4dwoFcC7e07UmtWn
1uZCJBwakwvrIfz1jdGcOfar9/l/cimGFnPR0y+s2QID4q5ntUZLG0OjnmY8OqzNmEpHm8FcXLqv
Ul6fHg1O5GfgUSfh6FPmLY24NXM3SlQWat3Dn4XnO1FqPFk3+ynT3T0eIQrJ/eyFhoFnPCI9VHsq
kIWQ7QbjpNhRiPyICorQUoXX3JVimogOyDtta2xXgfQQF5S+1Z3Gsfv/guxmuNGu9EYObOnDK4/s
Oi2iRUy3K5hD1ISwg0+3TTLlb10apkpDmqvAzifADHn8hVyUEE1So8Qb681BAbAXGLcEcFwI+KJA
ItB9Im3trXDNbB9wgSWwAqUDONBx5JDbo3gHvKqjH6Z/W2Q92yFxgAtBLAkr5NzfF1IFj41sR37j
FF6TwrUV5KhCUW38nmsXw47cS9q73aV+NKMUNHUnu0/WccCf+etZ6seXcBWcxcPhGUA0ziyZeJ8r
NcRuryR+PEGycWmQJbic49phj/K4Iu+r9FthUkoWpWvDVx9l2yM0Zr6bkjUqlAJofG7nG9lGbMqt
zjsUHtAODehHsPda0NaGLxC1yOB26pWge1fc/fhifMw1IBmEBIl4Tp8EDujXrvA9naiZBk6s1yYv
/AckHkiBbJBJlOpe2JHMRpUGhQ26Se42s07KAXNDKpcpRNDpRwTVBEZTJfI3Jv0qOohTP7poCpQd
otRVH5o4g3YUz9tqVWNaaPF2z8NBZ/rpXRvZNsIRGS96Gv3dqR0rp7go3T8KaknFfJOqWit77wpC
gNwijroydBvjvNtl6FX+Bvgtt+wzJUG7xGhX3+3cJmU/RnGurjJnhtpBesZQdF31USFmTPnRycgd
qGNmTLWHbkngWFAQ+cjyyoWagerYenTL3PtyVmwsc/LSgTRS1fmk+fsrW6O03xqYGrAgkzr7+FJC
6zJMVO1N1PK0iwXLKEup9ZkdeAR3oBlr2/fdgtifuwQI0SpwrLORBwCxg3hZ4r3v3msjimjSzhcZ
gUtuU9qlc/mfizvbH65wMq8e9ln+D2mDWQHXO3+83/jOlkjf3BfS0U+cG3QlHXJzp5VJ6c50nP1z
+TT29AMZdDuU47nIjMIJ0pX7tCuPm5aTnO3mRgYf+lop2QnRbQEuqK5PwRVAfpE/u8k1thsPHj1z
7HsAN1Qcb5zfwRSuz1BcNcPhA90HNNPKgckCGfnOG+d6J+K7FfTlfAFdjpePdr4RRa3fe3T33XbD
DKL3//XKCY7nbMIEoJi+OhYfTZKvJm0bEC8Vft/qubcWpIIQ9+eyPgBMh5S00jjfJtEXqGKI25rR
7i+oVvgd5PwE0FPvROSOLXju831gY26R57uiNdvRq665qfxH/yWGOt3cfR2glqKOJknHVIlP55IY
mNET2l1AH4Ns5cKuM9ifdbnKjeugMBktuppLE2bLJZJd5vpKh24x3IN86CS1cedldSYTuvZozVWZ
gGGKSfAStqdgaxPdnGYYJGPMqWn8jfbS+qTfNeEWj3evI2ZKTrAmQvnfBs4HxuX0zVUyXWviWeLj
wyWgvwP4eg1TFbHQ+sBt4h+StNA6JJxrYRBUws0DtBlO5Phg1XKXoEFz43FJQ+LEKzmAljvPj7bv
UmsvYSbz22jOSgDzw5mkNz1mTU17Zttjy4EJQnLlKeZo+GiN/VxMyKe5OUEFWYMUeygXPla/aju9
DxR2cl9M7oG+EF2EFIo0CjuPo9k7l4wq9VRtlNd60KRnqyPxUrR0M8SxZ5Ug6EEkI2LMqAYKyj16
xkD+vYbtzNK7yRTOGpwDc6pJBwTXEGR3XGkrTWVa5ZSjZf+z1ZzD/Q6lyrLsXX0vOcynaF9zzpTI
At2zwxurnfjOqCDbIYBnXGHRugC5fqiAyFTqkVj+y5b5eImlAn200B4nugxkSK7c6TPj1sVgqdQt
uowaykK7yK9Drz7KeGUFv1t0bJRnr9hRRoHQfuFc4+u4lzaG0HJy73r2rLk1Kk51NiojstFZYLUt
fmudSp1Kk8E4CMKfrhjnFPnDoKbhMrDYPDqWjEPTV33lh9FMwsetPoRcD//MbYCI0amCcoW1LcpI
0iXphrwq0TxpIKiStYaYZEMgP+kmGdrb55rfuG/H14YZ+AEPflNHF/Gp74lb/6I283pqaMyQSDPl
Lq/gIAflwwtHci51SXx7wYAv0fuh/S/p1dsUNssUescH9lwOo6SCslKwj/6nlZvs7DM4CR+rcN/C
9Rz268UuhNeMwtyAjun/yYRoncL5FId+0qlcipJBgAhO7b9XDGrY/9zR9ZpW75ik85SWr3WZERH+
shrWbNFYL62hurkAb21fa8DRfVoaKSVKssOSzOE43McmrsmmU9yo5nvk6s88no8L3kd7LtLJEuWH
Atu5m3jgVH5AkKfKdSr8P8y6U5r37RrZ0f99HhG2ChIMIO/2np7NTJW4QOPCJy72jLQZDlwtZU4C
pWxYl47qXjDUxencgQkOleN4XDboTfCVVOA5UeqAm5pJkkRdkgFewxooFnIj11WNrcTlI6gV3hnl
FP7slml//WyvRIwA9Bx9TCx5klRszz7/aJ+5OBZf2Ew32bs/ezuW0AhNB2W++EC+iuJTJSWKjX6M
WrSA7MRt543jQqhH1uxW9k/Fi/PW9TZvcto4Abw/DPm/Ocrgk9gC8ANpcy1+68Ec5RJvcx0dYH/I
RuYRCl1KyjbgtrnQmfK+OxFOG+a7OGo18bc8F9x0CruIjEIzYvd68kHmEesOWI3V75nDkFcknmCN
Qi/149qiL+Hlnh7maNkVbn8QPYX78noj6tBPKI5UvfDphVR7EyNkQ14dxNimVOwb/F2CbfDyMCac
fLmv8KqORqpDNyKY30EGc1ntRi4ikwdKvsYEHqnBwm57uLkZ1i2NNLYIrr9nKr18Yc9Xgj5x1nj+
4D3M426Q/uDVK5rKod8wA4hDD6uF/eFD4NK3Qq9DI/0xp86ke4WlcKzcvR7o4CyKq29jcMGW7r/z
Zl5oF3fmqqLMDh9sL0ly5/Z4c+p1+KbE+y4IcNguGxMqSlaPw5GAIgVubUMMw1gLKHo2lbAWqlWq
+oy3T/+jMw2T199VPDwBzxZoMMTdlIN0JCICeml4JSiRiKiFUfqCQKksMtk03Lijq7v/XfnsiAw6
+Qfs/oTevZEOhrFXsjFk4ZrAmM8Pfcr0K8vqkJbYwkxZYQaw5M1s4Kmd65/9gwh+bXMPOCl7W3NQ
Ap0ie4Se27RJHteVuQeJj8ABKFAH2Znc/XnHT4AFWR2BOdLqfdFLNwIfuJWQLxhgm956VOHMqHyC
Avs6dvyPRufeitTc9t3lCJsytZFVkkK2Sl5V9ApZO9Fk7vBLG0dTN7WOmu86dAWzt4k4J7YeVQBQ
nsfttHPl5LrB+zAg7KJbrUGa22ntcTmYoZqTnNH1OrBw2RuQ1pqzz8F4tsGojC/lYq9tJGLpmtpu
TPehDWaAmavwVALVbnIo4txdEDERj92+sc17HoFwLQElsfhxD8bfwfT16sSSBdG7CKflvFSoXGja
YpX6KD/iIv55AW+mGvcNDibLYx9nZDnCYlamMHRx3rp7utwXjJ6LboCXw6y7daCLmdaCiXBCdd3s
MjSJkER40dP+RYHUqzv6fPrYuISQDfhcA3tHG+QVQsmB7G9Nd04ub3izgIjhAxwWUDAfEQwbNAUq
uNW/dKuVR303by4z3+odYUf5d7+mvCc9Qyj/L1Zjo36shocrh4ouJEHZu4sRjnsW191qTtBCnor2
zWAlIdxE1wAiZ+juHV3pl8sOr5eXAf3ZiPkE/tLoNLOAjzuJbNO4/aOe4qNQ192QYbEEDPeWBqV9
uk59LOEYYQXJ0RE9m9irEJPuk/Pi/TvjhTef7eVHikaKus34b2JkhRjM4Z1vX2MuQTCpVXnI8h5b
44t/JJ6/iWasZYdaNNF0EmmlILKV7pevy/DJ8gJFDMSfpVTnNntT0pzrA5j7O+MxtjL8lRAQ7E0g
d/HzSZiM2Gng22gFU5y8nIa76wnMEHo1WHWWf2e9PDACjvRkwJkRRTTfCP0O5XoKlHaQIHjzPofO
XTJdztcnR0eM93XusnFmrpclIN+VudOYyesm/tMs0meFgL8zIJVr28c/Ul7zLJl03oinfKcYHV4e
C1ngxW/CW/c2d+fFzrYsmC/4maCvjsYi4W668caUM7GYQEJOgDBbpD87p9QaEk/30Z4/XawKE9Sx
KTFA2kbEpD4aBD4r/nRrG2kGlY9lbNk4BbxI4pejZQsqe4kUMIQqjQIQ5+YtIlWiSs0jGWuz+LEE
E5OjrTcMF1Hyxfivpkb4Hvxq9AdlFSueFJycNCcU4Wn/ZiKW3SiRZq83WJ2Cmb5o7utAcBouV209
Ok1gm+JVzcUCQkQoPRAy8UVUegb4Vo7jsTwqNrpkfyiieJYVjbhE3QEUl+LOPhCPdA96RNGSaAyO
wmd62C/bISxuTE2G0kV312rgJkvEdPQRIaMM2DP6iCg7ADHGoGUpMLx1MgO324m+mdQWDLahqnHJ
66UmExdFwxBSsmhIhRdhMerIfks0Dg0fPWJsY2jmAPtDq9kEJx1S8XTdHJfoNeCfkpRNq5HqoCmW
Dre3/o7yIjt05AGgP1yXdBDcLEpFF+KfmFRPfFKlnC1kPiPCo9qeKM8wgA4AEmgiHHpBZtnshjp/
Qw5HdjtVt58Gyt2NNEcYk1MpgnD1y9SSw2DHl/EYkQfxiNSjuCNYByudeG8P0F1/HZGiRH+q+kDU
N9qb6WU5kB0ItvicsR197ulHndTMkqYVE27qfE5EZU1/26x0CtpJHCizxlZWqJTE2F7McySIF94K
ekb7JbO3CPPAoxkLKvmIlmvaJG3LdESjK80psqrDfa4pc0wb+WKCqhD0br0y4rv4+3X4RjCPlpjH
RG5uTBt8yBIwKTHbnUm/Nn4pfXp67UqfkPO/VEVc4JrKtppiYPXmgCcs9aDIqBcYll6YvNiEDEfB
rhgCu4+XR39a+YIq29SK/DX5C5aDs/8JKZk3apHeofPkjmilB297wBGrvp58TqB8IpSgD1TNf5XG
YpGeLgUZSu0JEV4R+UY37om0gknTIzw2rJ5r6lKs0oDDLnGYMLGFv1RnSSZ3vl0UyU8Q6VCAUHzu
0YXfl/lhiZJ9sC+Gw/DvH19E6ZyUdxrJms9bBhBUUfRX58pvGGtzAP30fv+Eqof+Vy1qOwJUNKkk
4pLabAxgEc+958LdehgGUtO0hVBEZGE53Siar+cDq+gn5dO7Wc57miCq8BbqhMlpOgmCJavI+dLB
lc2iqtwwRA8Prje1o2mY/FETRHJHek1hIrJrbUIcAodrN+jECdfs20rpBd97XP263/ZTOTWxiKk4
JRZa0ybVZMOSQ0LvjWohzeDz04U0ZIwgSHlpxvIIXJzavN90OPsClNH7Q14dCW8AYu7GmDYgH87f
R3pDaQ1I1QUJEXpG7C6OEUAamSRQfWSaD+CrDiz3m+UUgZcNNHQTJP4PBidKEOpuyEPTqNwcPNkn
AljPC+ZwaA/zDl8uyGjLEE35MU8nAYxdCUWLDf1S63bvWfpSFR4JuhoEHOKdcWOh3QLW/l/MgFUk
+5n2qWd3IJnTtYbKRJjVelDkgpON1+iqFmtHaj0M7AljZsHpwAoQNgbhVgC654t+secP1qGLSG1y
eG39C8VAie5amrqLDXB8esqmHicZ6GVxy3ZDh0k4W6wxGM6VqvYfyAxSP23hCRSpOOahhUOUquhC
6eT1528IDVq1DP9plc+qiqgcWtS2q6OFl7RZZRHaVqN+iwJ95uHGk/b1oYdOz65PjEx5ZFbA6GRA
Dk/nxH8oVAE23/wCK6/QaAIw8zKg44LJs30hfJW5Q8i1lOYxfm5aT+R+U5ec9Q5JR8qYRDt4ImrW
7weAcr8jXVje80gnMSMCSojGw0FZbcF9nGouQk4tWJEZwAs1KdNYYbKQ6COP4io6fCvMnO/S4hM0
JohdieO0zDKNMDZ6F5Gs6HtvCVIbSFtO6Xdzl6LrRhEcM1Dxr5Q1UQB/m8yFRxioqBIakrIkVzSE
xV25YDqi4lk1PWY1aKh7RNJpNFoUjUdOqPMF2M83h/7D0xmDzXBm03ronAVJpsqsGNAkn8colLSB
tKdL4SxPMOhHNqIl6vXI7YasMiHdniSpPUmmRFQd3WFCPoz0ZBh1a8y2wTPPNRIY92TfRaiyNicF
a/cWGGCFnh7TbR39/DhQrUkX+aIlC3TTzhsT9+I+0J5UAMhrT6NnfCw5q8aHovEzE+5+qAl8TG9N
8rqLu6X9RY5zBoQwhFfMinBWZ2mKJ/EtwYOeYUyiJcb+o2fihgABjw2iVkloX22le2LHUJocDgdx
HqjjlDP9ZXWZ4pcwFJSzQnioH7SKmtANufDJIU++ftg7brOyoG4Tvl+tnHRUw0GhMD/4P6PS/zZm
ZAYK5Jz/dSrj3XynT4YbQnz2ZrmBSkNamM8WUHEhoqjK/mniuKtSFUkKgr8HFf94ez1AhvfFTyt2
+vGCv8Rcg9M7yML+yXft9t+TOliKYH6vmNWw2YCPSWf34YDXLbwhwZ8xw920sWon64+sWGTTgkTF
A00A1YwATEzxkF7TNnKo+7cLKE9JKML0JmcTy9qYM3p16oad+ILwVQCoMvTbqak+vmenRAh69Ssx
iK+HSLBxOkP/l6jJjqSZuVXTHlYrhuUJuezGUmYbdQT+ATF8k60YxPb4G2T7ek96RB5+zdejRb9U
Y2iCgD1n7RbDV5ccmgDTs9zOZIXZTYfcg59xUlbLww07BoQGcQEEouR4dVwwNEsoBpXvIi8yotJM
rGwNU2h878Yr8l4sX+igpV7HbbeBnozWMNxwYKEJZAmDs+BPxO9a8oPMSYSB/3BM5oSp4XdwJESi
eqwZoWftpkOkBK4AS7F95IEBoFvfCa7bd3SB8/iiUsQutxqdnWRQHYBCMkVv1SrqUyWfTs6Xdgff
NbPZ+XQDeLh8Dla+Yggf5XFT+15cDgW7bY33JbCpsFXCM9ll24FRjXSSNVdVoCBYpxJxFLCQ4Cse
71cYnmh5sZSYPUPEGhmURE0du4EwlMvAzc+yoJJxdaDHq+LNovwWQWt6sqSgi/1o460Pj7zKiu+7
EQ1Lkh6SikM2JtCEqzI5OEWIZ29vlgdhHExuR4JfjEiNlvS3jw/EVQDWCoyoOwN+NOGPh5b0thhq
8P8DYChj4NBWzQ09sbowG6aOhUoTY7amk3Rr6VFyGDt9Ygwn642WpFnwrZ9oiSvMEQ6CqsBrpqH6
fNGypbmmJ+hMgMlX44rYkbSZBNxH8D4oUTAGVZnJktTMeehvNLWnJPKLimnn/2KV4dGmjBBgLWYA
adETN33wTr9XFignuJpSBqWGwo4CkrZiURttVmgfMxJN+VD8d+cNpQDBFLTfGGP+PtCrJEEEgEtK
DK568WnHk4XPvkE50w5Ngcq1JR/Z6JT1DY1koRtrGIA7hJ2DpftrQ9HoKk2+Ps6ZLjJvVbPE+Neq
ish03ju2kTYpVU6hkECMEra3TgPTWMx9yrcrb/yfFoZsp2TSIySMTORYMFtv7OXyDkbiqA3kJMrO
c0zNfvCFRbWvXZDGR+RZsnPCmgLWFC1QFsxzQFQ/IFeyCOmAUhNTVLzlfQgxggAbIJa8+QMRJ5Mf
0bWKijrAEv0K6AnWjw3vruw4uhoB1xJr7LdUgUT+fdOBPBUUFPD5pj6988YMA+M4/U39ZGvdweEG
Wx/ISSo56cwGIH+d9+5Pkbre6OspMEQfPBiS9uvemBcb7alZr3svO5obzMWhOPrbfImPz4UkqXWP
y/kCeVlQlgUSJV0lIHi5nKBDWfwGv03CYR301ANYhFpFyr+3wCA0VvkedURRAHGjWJsNqV+wDqAV
PJraifECVMR5InKAiIWE/KI6iS8ROFnBTWT2v5+0NOzdtbpYjTwnzi6HtoPo4YlOFH4PMGGmyQMb
j5qtxkKZdI6FBi17DiBE2hCl7DC2NhwFA6+ScXGnBH6X7fi6F5fa3hDlR1gfjJ/0yN7XLkPokB4Q
WUhTsva/iSgc/6f92HVUBOYnyPgIh8qApfo+dG+rpSBqhd2g5xzHGGRzY6ummb9YPx4zV8MIxyM4
P3B/IWG2CB7NUpW4dWc3coeO02FPnMsHo2Mehit+4aaVMN+w5zXf2gR0kEXel87gaTadTbhXYeMv
FkClHNf0sQkMGfBVJoTSM+kDU1E0x3yL/uXEyetftgVESxWrbfXhJHLkuO+XTnE9+qbQz91lkqMA
u8Z7zya2gB6SmV3DCDZ6KAIpJGLe8QsWwqZhBvapjrq9yjPQQ186OAdLRECt09+2pHTmzfqNpyLQ
DNwPnykUg0dA0KFJlnUkadwLa5AEriOP17SFsSWYTp5NozwPyogAP0NpgcW4GUMlEuOX9RImiIb2
98hH0qci/IaV3ffd01En88LPUjmCYMFuFSzPZWG4n7rBpIS6sbjxMJ/kzeRP0wwPHVYhbPNJ/jP1
7RuXSUvee7j/chjE2XtRwq1y5aA2ECk/fDRQva/QoW/HY54Py0PyoNzmwgRuJe5YLyt0dRWNzik0
WtUtcJOCexSxaN/9TTnjh6G+wxHNomRYeYNYrNDUOvIwjINt/AovCi2uAzoFYgID8btn7jXZuO2w
s97RoOj/ZSPkxA72Es17QJfdzlvBSDCDYPJII82dSenJJx17vhShGqTGkjsZK5fWnPuORQnr/5K6
tVaAUABM8/S4Xv2Twg47nI9NNcyCNIoCuNNZlre7s4U8/eyfHo08HtuoY3tEakOG4uQIQG4JIi42
/nh/KJbUp1Ywk6m3d14Zu25bbhtij+7yo/wiZsK2Xom6ha0GVopL0j6T30gacsLOQeFiBNXUn7bS
D6czxFuMkruoeNrJ9cHLjFT3i5e7PTmSUTppYCfD90Y57NWYCjW8uNeREnVWMb2J4M4dacxqnbj9
Mjyj8xmj1DBB0P1r5r7u5Au24Mx0O8wiS02jQpDVg+h29jyrdbe3cLryk1faW/6HzReW5aPqCbwk
c9M/GQ9fD3YDYkpV7XHiRI0PqOkFC9O+DGNFeUQyt7qro2WxY2AVvtqrrkfjUXu0YcT+mwAggo/+
Y41gBkBEVPpHY7rLHemHY7YY9n++NcB0U1JNBckZTrwH/1ZdKGbtnDNV5aZ/2TZIaQ0M/Z5LRqFc
sE0ULkAHJLW+wugMluqXlnNIUQb7V1/NkS76cfyLaOj1BP3QbA/KxGe7IcuX+kaQIscMH4mjZyZy
8JRLAdxbvBfasqce7doYDpl/e6WTRCvEivnkZjsClhf7dCFhP5iyyy9Nklefy4O6j2chIPnMQQBH
3Y3I8bDsbSU8PUAByb9DyZz7ghUpAD0AoiRXriNhlFpj3mss9QkyX4ly/YNpU+Ms1olk4PXXtIHS
aKs7kINLlFDm/UVffia75q+X+fKaFl15+oJEV+kZFxBjJ5oFTBwD6zHdiRnME9GT+2JvNL7kmczw
CjKO5b07NPmeu5L47EI31ZD4M+IYei+omakFKtHtZEleejVO7gvL63Ds7mtgt0y6CQgkUNiLpHpG
FXcrpC2W64LNqK6Gm/2cRnXMl2AV3pYUnFGFiiBZX1Bv6u3aSTRTgZLHFBznhLHZPi7JC/5tPT2I
UKURWEmArpiqyvRidSSLJf8f3EyNZxfqjAdfx+FCVBBoGIHww7IEme0DvnBxDp9Uit1NhXTbPh6m
29G5887GMXiwAVA6mm7pWEVlKNtvFv2MLyg+CY4qF04bebHrGj+l3QzH5Mw7UER+9eOsWgOjmOes
+SwwWFtO9SWmWWx0FEnKG/KwTh8koJ1ET06OZylIHhs4TMvlZ+H8OdU4s4qeI55059Axh0xH/n7D
28NJhP4YBLPho9eoiYxRVgQIerO1NG7pgZn86gLvO9q5+gTNEKMqj//Rn4djR36clua1KJrGI7k4
GEbp7ndwiA05RnB+mC0Ba20c1Ye1C8Q0QmFDjccYyGxE9WAvh2gELU+IDO4+Eq2q9S02xapxI2rB
A0/2/jOTok6ThmWomDuPzMYknfNJsi14B12VzAbzmG892uKXVl0hk3fmSkeXu9O+2ee6ht3D/3W1
jiQOUZ5BRpU/jJp1ZectpteNccUGGrUFaviFKjE+/5ij5oVoC9NmPY7zkC8a10llc0QGek1Uy7AQ
C3XiAxXT8GsJjOZY+cLLu6pZ02F9ZjqvWPHuPFASq6Sj9uNJFXRQjrJQw4xBQU3b0dsLn3/HARLI
qd/MhhTAGt16kUZgTsu1ZsnnQCFgAITs9gDrn3V3DQn4Vghu7YE1ZU9QIhOo+IVCMXq384mDAwlg
o8sORG1DH6K03OoFVrC8OpRz4Ra827LsxKK/NJ8ViaMmz6mY7YR4ok3HoP/mY95FfC1hD9eWer4a
Xo6/vlvN+S9H58u8k0wIEjHSJHSZQBDvj65lzmbk4stoErOQOyTNC1xxmO8ThwuHJ85c7zceLzpy
QmZoX5EXRfalQ/1jD9fYv151QvwdDznwIB2IdWELCugPhTMcS/GT7jw3BU1x1m6pKGLyMfADxcYi
R2SCn64hLpf61FoJX1+G9HckwKHPGUQngnABfvAULcLbZfkl/RnB0gzj1kGIlkPz3dDHKauTDo/J
xMR+H7LNBvO3YlvIAcOuuD2nhGt/MeP8XIK7ECCU5KKGkgJSXafpJJym/RWflWnlg4ZH7iC86Ab6
pDRipckDnnnkOJ6BbozeeWhlOHZDJLGDFDFu35F/0vJPmpYDuwrGgjQbbqC0efr+Y2dF6QgNSgbQ
/2BRlLm8F0DJWMXXSwxpsf/6PPYtU8YPGYv2VmMawx7DTSrydNDAYUPoVu6jsGlHkumSaFKARnKK
gYrble22T1ZYPYAe4ACuKA1KP/D1dW2218Jb8Ypaz+ttbXPp3PUBqTReqrXCOQ8hpatjN0TkI+ts
Yt2h+LHjhbJl747khzlVRB4HF6hnVcZMErpsC2IXVY+/T59YQRLrFOp1qWCD4D7nePIH7C3DxgWD
C4VVUB82ZnQLPYHDzk4gGxdx0HjTL9vrquDgrAHTv8JOtH0B+TbWczYnj+h+9Wd1mQL2O57fuBdP
rQfIpEMZVOD0jQT8outH9aR8cw/K2SCNvUhZ4TbaN4FuctRc1bps12mNXtxwkt+Yk6Z7ZCiWxHm0
wurP8YVpraLlKTxajgeZrRN6ecEiXG0G/CUWPmwaOLnCR5RXvwu0RTw5iMXG1gZXfNJwovSoCfoz
9B/Rtf3z5Qa8FzlUbGl439MQ9VR3Jc7Dtv0YGcR6l7wzgPh6OJ8TGfdT0dEli+8UiiVm+q3VEAVO
pZmmDLjN09MQIV1DSbZbm5B3fALuSs7kiE61e6xudY0upvnWOXL4tJ2jHo49qheKru2DTjqngSWQ
NPwXjPUIn/gO+pJSwNzYPTW2eu/P4U1dZKHYTlN4QbyZJaxCyetlAoFEI9TZESKXVn5wqaSd7jey
EZShvIZ9hxYnJW1/9mAinbv02ANCYizsbeiAoz9QSTE00i8eV52bW+fXW607C6qW9rprpzngHwIA
tuopJitOilAOsp1gM63SluTbvZD5XfDgtZNaWgTPZ+EoGhH7p0Hf7Rx+Z/7HE7l3FRd6HvMlrIXc
zgPcfrkzsUCZqobMo/PXNRSoG0CRJvJTYUpN8C5tAHsSAUcWiwPV+usk7xi8Lp4zz0iNqgr1SdLS
Qa295Tn127uhV/E5+47j64GieSakDPGbSUGEUB8NmlRMiKHtfjaYSBVOjop61kC4lD0iEhYX4T7I
+jk+UnbhOQlTPUmZhSBUFECV6jIUu5f4IHV1Gymey/e07OtrOMMZHcP7z08HTgsN9CIwgiDEi0QW
MeMFR8aytbCqqpFsFPX/HErI8wWVrRLEKldFmm3nJwTpjviNG6ahZ5iiyfDfemHmbZi9KxpkWUS/
nQTb4ZyRAuJcJH9o18DEWkXnG2bJSME6ibO4vpV1Ir3RUSPJUrv84EnvWqc9o8I8H5zdS2gP0Kku
shkB/Z5PmEEABOAxJb6sE9PxXgJcrIvAsr8iiPN5LHA+JaXkeDenV9vA34E5fLd/3eQO7oBOPUE4
r+elamV2BQhtcrlk7ooW36IbVaxG2W1m6f2qOLCW/iPYkCDbmAgRHW3J5h0A32k9rz6V2scsNeqN
OQM2X9XCurs4jxRs5DKNYukXvpv1PBJ0ggCTsf97mDKjR1BNeAl/BZzIDabNVTRKo43pASmuG4UL
YPgovO6mLtp219dsJBWuitYALU4yRpZANMILiH0Nzj+hnjRke4wWvqMcj84chsQgjEMfY5jYJOhi
hhqUpWfz9z8BLs2GRB4Rol0KPBI9MVCKEFLr9mAYneTd9Hj2WMVCiYr9z7GzSLQ8x8riL9k/cLnd
MWQ7GLZCprUvEc34whHbf1Ax8GTh9TBbvwairx2AKEXskiAitjM1KNUt8aEQVF4C/iabd+bQUboI
Tn6UUajoFjxki6GbeBDQTzUnN5g7ZdbhzOM+l3+rkj57/N2thdbClONYDf971U+4rgddQ81U0eva
fdiR5bjcjpsX4L+MSwKdZ7y0elnFBEGqx/afsZgxr5mylPckjQqE07mxBemT0wgCUsVANnHC7Mf4
l5B0WiMLzBCTYFhjAAo6+rWLf+H1DF5QT2OIvf2bo0LRuLV9X2VJOdtkSV2FFHlWJ7KizUCpHcYc
00ffRtV9wJV79YxuFL9X4lPXYsyBasCoH9/TkIg6TFm5WiT5jAAoFRYxbFjoUfMAod5POfKT2Xs+
MlDaC5zesojL1RsMPZsL5+ILBrE5LTkTHFUyfkusr67pP7UdulCaL4efE8NVThMB9lpeXaQBUGQQ
o0sEuyAlQFFc6HIq+b2dSk5rVPR4pmb5wdMA+fybGF2D+FEEXkEOatX5z4qQ8Lgz2HNUhzsvUzIY
1KirXmuq96un+1MHBm7cY2zyhOf9i5a2fxebMegLrv8ZtIKL72YpNtqxLnvxuT9HKl7UfSCPMfLB
9QSSyG63vBRJCIVWvLIhzAUafZZHsxc9P8THVopVaQJ67+tAFoZyjYH03OGzFM/HucPtReGZ2RcT
gRbmeC9RdRHQDGUV1I93n6PnvJdyxvr1lUSQLiieQDfLKx5lIbPDplsmUz0URy6jfGP2b/i4JJoI
V55vyOR2oWvWxoYc9StI/+11ZpLffypSUHCsIE+WfVsBW9z+e/+tPlC0WZwXELMfc57JC1HerCNc
7/yMnITTT4CyfFh77i1tjEGlljJ6DsRJnneU/XSImwfRDFC8A7Clm0geVf++kXqXwYudbVg+5KD1
/4Ms0GjUigukOiOgSWguZ6d3Ge5O4n3sU4svlJpDhTQTrycK1/dD5DsODB/0om8b8qnZlcQbWaz/
Ouev8zk6UyPcA7BscGhb0ZJUaKAG7Wqq2uZLg5WAIvoqn9to5I1/B1zDkBAHUXGWUADP1WBG9tGY
jSuS6sFwJSyj88SJ6xEZsqjwXvR6+Xa9PEXNTovhc64DztuIGxxc95PGKO0JpNNI35Qg1xr4oAsj
FsPqBkoNZG9+Gz7s82e3hhVfp3F7riq56zOs9BZMRFFvZENpLOKbAexH8dnJujNIk2Hvc1/3PaGI
SIiZavY3KxY+Hw54T7KVqGNfNnltL75TOe2xiHgtKQnhnqNXQmEJSYAlfSNFabsSYobXRuPdDd5W
VHpZiw4Uk/p+ValpMlPUAI2hGaNR4uJl/X08l8800Q/vPO13QCBkWiYQhfFbDT57OMmzhwAxHvBX
8/abmeJ4J/kgUxS+YKPM6aUpjZ68v6Fo3PU4NX3MdbyMXstPsSS/RmogHlL3lPThy5RAJNNOKv4l
DO//2GPlDixhvRsrDBg6vyp9Mh3Pn2/e9JN581g4eqjpCAvBwZJosVoYbAc4rhwRj2jHROB6Nexy
ydevRrQc5MywEP8lOBYooKTpfljOw2dl4BvUlCxjiya9h1oz1fARD9mrCcIlfaIrPGS53mz7sqmN
7gnA7pwtFWvik+KnqHhczzd+DbZYrJfAbO7rCamPGQ9B5ssaFIDld/noz+GFDi219ia+U0vQYXkR
yhHusGAD/qYhXPGizDIY3Y+5SHtpW9AjOTdy+YOz2a4zKDrS1VC/XmG1sgZKu8WLSPjo/sddTs2Q
kCfYoxR+uHQUXug9RcSYtgIKrM68cgQ7tCTuYrWQsVvBmilM8N7wgnmyOvvC33eahlWiNl2/vInL
CdML3MwZMLdbMdJr9jTp3CJPDJCmyxBjGbKQpo0xRmz41rKO2kL9dEff4MD1aOt93M2ta4TKXlKv
OJUKGrXuFq0bzuwisvKhKu96Fm72+diS0nHhnfCfYrpB4uSbPMSspQlzzDFeVK4L/dEdjHQ+4P1V
2waUgfuSafu9WrtQX+lpmO4Nc7ItXdA4u3q9tuefjBCxuQO9XGnKy2WciWXrYVd5XNfrK1O8fI7E
YF3gEA/vL+obauBAA8gbK6xcSuckVw+OEKHZDwEKGu/pwA5X4CwKdVd0sZOBOjBK6oc2/Ct2Ir76
EFi9AXjD02qxHj/kL8eYq+xBnkS0EadL7QLefgCvK3v25nqITYBmxJ3PDLWTTe0jl3IxJoYyz1hM
/DspHzLmM1Mu+PPyHYpOlV13E3/WGvYGsCU5McWY0OqWN7HCc9q+oWczaWTeXx/U4OoHdVPH44e8
YMDvc4lHKE3l3mxZ2moA5DIj9dtwq5yS5ppmCYMBxuTkrb/XCEL9lbLabXkDbKq3Tq6Wt/rN2YuA
nNvnbZwAkcUfpcSswKrBhvYKWjhdQdNDsKLr0bOX3h0EjwNx9HWHaHEk7IaPhCtlM+zvOt9vTDlf
awXCyHd1wrR3GwYN0iFkAkhuF/IA5FQUWQVwPpWHPvwSo9+qCwbA9Kuq3H/KRZwvFG122ihvcmwr
3/JtwYUTEt+DtYSH+K8FK2ZtNOhYR/8yKhemp5N6Mx3oopC34I7ohYbmlwdx/esr+Wv4fKiZENPn
fc1snJAbdmp+p+I+9Skspwclp1uyWRrl7Uq/6sHI9UhzWE5DmEjVQHV//0Kvs4PIe0ODOojoKzVv
PBDy5tVsJB1IX5sQorjsCLJiuhqcyJkNlgUdPTbDeDQPjWRc4bJVNrMmmuY0FoxX3SD3sPvSSH9f
nFPb9xXdVSdM0SSL8jltGNHWO7pYXV7Mr2Vmf2TmECOEDy/H8FLVc8Vp3sReomD57XIBKpfdiewU
XSrFSjxpUgLAEHXK6xVhBEMYP+LENuCbxHu4C4ZDFLL5BfFUDKPPHf7nSj86p+X7cGZ2/C2Yeg+7
7YeXYmlOYsUncuhk7tMeQR/0TOb3OkVXH9+0p7PuGEjuggmKfiJY7N6Spw6wVSn5JQGuDE/qiM4l
jOJGI28JeQK4mAWiFn2iGlJ40zYXwRwe7Kctm01B1P5U2zCVZiwVQ4/ieHO12GhZ+nCPGLgXlmcp
1P8dpR6bv6NgG5eL4Yra/IhX/FVCErcfA7NG3RwD5/uL6bdhFzDEyL5Byiuf7t1uNtdSbOc+y8Me
Trmh/DEZkCa5JraSwdEal4jc1LTVrFYdqJn8LYUvN4KcQYoz7FFWysx81O4fCK+wRop61ReFu9bw
0LPn8tvPWvyJGqpq7k/tCExujzaze3lcpft+CaVawkVNRZVyo+mLYdheHt8J5TNAhDZUnY4zXTd6
pA7LOx1lUfTkGi6vxNq4lPi57ZqR4VKkb8U9vrsbPHK5FWAfr+hxbhfN1g6nbYGV+3j0O1ACG2W/
khbdOcmijg8xtDajx7omCAle+GHpngLtjBNrGRCJCdocFmqUTqo4MjMHdXY3z4OGXxCKo2XVsliq
mIj6JW7DX3fxm2bbPLYfTWN6RyHhad7I6wh0Rg/8Wy2wqPKQURmWWIG+PsBBx3Qu7oPEV0yHWVY1
n8FOtUxhjrWgnYy5NBV/n00vgxDDHnrxSbDcP37z6cUAka74ZiYJdi2nzDaBpeg2Nq7jnylXcHR1
2E8ftAGqxSRXKfAne1DNnyQFjC5i5jxRL4DZdfCEfPTaOgou+I4KXfN5Jaw/Ys1QDpdHh2y33jXu
p2UEjlObYh9rZ7/J10BjyG/vE/osZzKhy8c6KlJZoGCwEyCA4a7Tl+tAVP4RY/oJgDPxkEfms4gP
k5kP389DEEVaru7KJ+BCgDCwUULBX3iIxQpsAuoxi9ynBBIGmk/yjMJohYEJ7VZ1aCusme5jZh6b
ekoE0Tfa1CNp7TRvE1bp4i+UFbdQhrLQjuWJXwu1I2rfsKPfNNmr5o+0GpHXSvwxr6dGumnxN+lW
w6fwzAmIeLJWJj/6yJSUcqfU0RV1fj6CQ8zhbprzoHR6fo5oke2diDW4DOhVC961ekrJpBVHbUiw
u+nRvYVqTXpRi8MGWtp5XI9PgmEKRvnMXja+xBit0Lkx902lwTNsoyjq1Op9Bnd780ySu/j24uOK
rL3ZNriSDvb0JwnIjjjctUt8wIXM2NUw5xF9EfF48XyTgyysu/lb8mZQ9MUDhe92K/cr8prmi264
1HriPs4w0uR3He3SA03s8+Oyc1BQAJQ9HFRN1+4ah9s+4T5YgZph1tLInEvb+j2/nLQCN9ile5S2
Cz73Kw9SbGIaNOzIZih9DYJ0rQ8KzqapHL4t441eosBOt0Z/uOv4J7E2U0FLvbKvHTzSl0GSe0fE
p4bwKtiehFx4fVZgz7ZFMpQRw8qkAYrvgZny65rSV97O4eBcX1l/ib6rMg8U2DWostWgmw86T2/2
H5regEVYfKcirG76KfUGzlpww1jR+VYsZHiS9PNtOXS3c/r9b1c0UZl25UemsaW217p8qwCzo3Ig
U0lEbjVxCvTNP4fQdOgcqEM0UirfLwTsp4c/d0uZO3QeUtFcOXnPpx5+2C3K1fL4e7XNOJ/KdBNl
Q8sjvwBOqMYIozEGYqorBM+Q3qYXhQXkayeW3Ge9P58hZBd+0cZpOKXlppCNL81XrESKG9JGt9Z6
HiicCATz4nJH5f140wowNV5fn2C/TeDtecf/EcVrzZ6boX8y09nKunYrBAGjJARrnshN+9wDtouV
AWU+GJ0kQ20cRzk1oXCLehkGn+UQw529+LVw80WM/HYRZBkpVEwMe9IYT4egDPt3YBTJfP2Ph7BF
AjYinLZWGlxRc6cmD0K/JUJCplmGSjZEO4exmBZKCX1KplU+W6O1c8+f8oYyg5NfJFBA6+Qj7zu3
EKWdGKNQUqV8iCRFTcHXSTiGkB3OnguRClN/XePr2b5robmqHAQ5wlslCMoy93YvkASWocgy7OaM
EZLPf1DW6pIbkSN0uMoYgW3w1/dfOOQTP+dFArBCTfGNIUrmH1j5Meet/UW/QgzNoYHHhZh6aFF4
cfq7+AA47bNXVHqRdAxVCQwSEW+OL/Y26eBPu6UIf+4gyTn5hUVCufw0wyYJhzB4YcGsZx1PZBXx
feP31dStSJA7vZIgJu8rwvsx80wRrCkxqhGuSiQf70ztkX712tA9Om3vquL3c9++Dtg1SsFA+fkz
MfuJk/y+CTWoy3mdEqWkMXS7uRB8XM9Si/zNbHurfccHaxhDL3aZwFFX0Eg9vqSDEGdnsFes/IwA
Ram/eOFIQ/3iOYLgsW1RTuhqOT9x6uCe0lE/PO3TzCwgWhA7n/DH2T98LLBZ7doqEPgr8hYQoDS9
eDELySSf9i5gviwwubq+p5n1JyYiGuAuGm5HC02M4OlN874oeTUVohX8zfxgrYE5p8JuUk0/qaR5
xH04DV7PiNKi6hQ6fJMscDrHdSOjCKjgt4WQVjjFAgoAAUABVC5xnbPrf7P1ydglhJXCbpTwKkUJ
T8JBQbuell4sdHeZN397qvod35H7KnZzGk/1yhHGSp7iG7xkjWb9N44IeLKcLsz1d6vhYfy04X3d
+v9xVpn1NzG6TLjaK/e19TGosSiNwA4g9k+ZZzL1mUp0P1L3CUFGhecW95Or6q5GNWw+42xHLSjN
b2k8T50i8gGPEfW/hkqEr6s2nK0exWwRj4fKtVd775SqbDwqykx5zQ7aeGa4bjxLUiozWT2Wiig0
J0/5yKUm0NZrPWGE4Yg/1f971mvWbXwoXFSo21aheu84TcBBBgtLg16kyUibvqs6RD/sGhHbJW8L
HY+ID9BZDAbDdxVHf05yiCnrJlLTz9skjiQ9idkZnbDOSdZ3IZMGs86mzrlyUfowG+yloASv5hn9
l1MdfpuTGTIpkiCjlDHgwhkc9vf+PlkgQ7j97+DWO32Kk0shwGAqhGVJqAnIwZpmHqMb3or7Cztr
Rlta9EJsXotwZUTXf7tIj18/1OI5MJM7cO4yQ42c5UEr6ByzqoXsuR1W+7AeVQwGxS3h/c9W6x3v
i/rLPE5vt5UNxhFCVE7AJmhoHC5wV6FZyQlDBqgF0etV/5vtTh4weDVg1NY9ltiOPD7CNBGfbh6s
jyCdsaYNSPP3vctDg2sxYvnSMDvgjurzx0ihbMuuAhyf/dlLUj9UR6EcFfqD01LxO4pQJyDcqufx
bHma9HPCKfZefyZi8fpEhXOHfoGVifESGdFK3043NVFj6HgbQ01jTtzoWrpT2U1MYAezf3ilM4vq
qPPYAcVWsNkNl6Ho61JZyAxYjK1eiymGcmjMsl/DJcopiR070ss92tzRReHvSHr0USdIKFWJEQts
hkzI4TrBolcnWZqptqAlmLTbDh7i31bD/6FAF9x9FtpY8uGDyXLxLBjhcNRKeQmvZDGzK2zlIKPS
I8iF9CI4QmJs8SVSlDrxOQ6be7fYybqGmHjhisbpA3sl8HTwIj9PuJCHGfCmgmtgkMB6AVUQXiTT
UEOpMO2Xgw6tKY1bN1l0ukbmtTXEJ0f66L8OGD77jWLw7fYf4ZbfmmwYhNTvdq01sIeYL6pYwtu0
80P3UcGUqWPoqSzgsRbr1cY7sivaShV+TKGQwQyWL9gf+ZawcblZ+iwd6JU2Mad3S1jjSg4fmIgd
e4Xgc/Av365rMoW5cpMzKf/xFwpgO/EZHUs+1IsuLWqeTz+jUhJg3mzzdCwncbP5b0u8igiiCQWB
t8J+6/HevGaB1t/n+t1hTUr1YAYaJEYUnO/ATryJeX/hXnjaYkSzv+qmCqVgwT5wQOqu030zSq2w
Qht2eznh9SNYy0MvfQXiOR23eQ1u6R9q50+Pxwql1/st91CZQEjNDNEKSVyM3z3xYazUQZnPxKTa
sp0mxww/LyY1OsCc5Q61mcBW5PLz7NalNZHPFfcZEYIE9Qq2haS9zYeukquJjqStoQyijqf9bWp6
YYkVdAlrXA1a0wj6Ne1xEyIyAMLKNhhxiXsd6klm9lxwZUP3NHF3htx68cxgy1znY2C0A/3zwSag
vk19/82z+cLSwzmMIJ9efbOneoDEWUzlaiIlwOOl3uTwPK0NYpKSuOWucOfeMtQVeGMJoUgz2/AG
mBZESrYQ7xDVY0kkY7K01MuemrqectisFKx0CMPUAo4OouCXUssdh544Acm4lRddzATL54RwCfpA
CajSYuTxBACrXj/9lcq5ySdu3uy2anuH40DGzLlqkVAS6KlxJSTwIR0B+zJOxu5mNG0Qorr5/DCQ
SezSj2/OsvU/6T5+o5xQsAmpfs8TeywxMe8rCoDNpCkEK8a5NSaqSO0eS1dAC4twV75VhGNQrGZO
2goCsHleL9nHwZIYyXVQnQcprSkyg2r/ZRcDQdDb3y94c+x6QT499fj+FLtPfG492p3Y3cqP6HLx
m6+0W+LaFhVQM1jCiVta1DQ/2mklfzv4NFUuZOEF6/S3i1Xjy9tKdW29pGFn1mGcOFBMztzfi99B
v6Sx1/V8W99wCsBubmJyy52N3dAC0D9XEaR5Zzf9NhabdTJWHvft/bZ5IoH8p7W8CCH+BoLJ1khU
IGh8cDMc8jP4rommBPqI0q6B/yKkbbyE0QFADSRI0L0GaJq8dPBb9RHY7z49EtHdFNAeiDD9EzAT
Wi8ddl4Fs19NqVD57qApoSfEUa/c90cDIRvFOf1NywuxCqNyK8i758F86JP1DAFLcfPR4lVSR7yM
hucp9Rz7pBhA86hreQ7VfUA4qMQWNoSdtahmKkOp4sL8CtdwqtOramEbgg794Y+xF4GL24Z1uIUz
UnZJ4MP1EG51WKh9OzjFb87YkPd3VseLp3hTA9qRm6LusYL0F5QDgYRP6PhGfdhoVhLYV/ewI9BG
Sj3MDhP0ogbttBNxfUXT2b0Nh5XaRC2SJMcvU/xru/mxyu7xxXbTtIzFNB+pEjlfky3Q233YWyuV
gp35TCayRjF5IcDG/xUFHhMpc6iqJFe3UjSxEJJ9/VKIaEHNsxCbExkinAQV5rUlRpXAzd7z7HZx
UU0SMzma9HRKz2/Lf5hkJ9sIllshyjjbtVxp04L9NRNVeXtvV6slBlfut/QVlBUt/RicpTxgPMF0
QS1Zh64TbEIZzS1RqVMa1CEAz2pt9Pxq9FhJqKENt6cz5Pw0w9ggo2YTLrYHDkWdLpz9LPPNLz/n
orwoqdb/In/2WjxQ/rx5hJPtykOR6GcnXGhQsZ94elc6onq7Wo1juMrifAQkCQDpBNaN06AD9Bjq
Mdk0iO4/m1FIr++EuSW177dtR2kwtMzZdJn8kIKa4nqyVKeyKRFic9NuxjuQu7Bg5qOh/Ye82BLj
8tkcBPTb/iuA8xSVBYZkOh4zo4jpI+g3K/FrYBTdtb96LGB0k3oDWDCvXRZeVC5eFQClhwzeMM64
w3yRMGbZivoWEmXUj8zsvH9PWFF1Z8vB0Q4gd0RODO/ksmqax156jlLaCwzRZooRp1nkfVBsQHGk
J8ZMr2UupwzrXwjD3oyvvvHHDR4tP6+3vW5PsLZb2FU/ulrN6W1ORl5oio+HxKa7y5xNogcMpEo1
rHE5yypo24/DtlG5b3NbXGssGmWrItLIk+cGoTQ8CMamJYzcazTD1wBmDeebVUmLqihLa0FD4KG8
Bwr+QyXXvLaOhLhHhgHVyQ4NOnGJyVzjiCBlBkaE4s2qQiJt6Yd8NEmCCfcScTFr7uta4NoL/S4Q
9+FP9Q7aiQQoaAOm8xPfnvQyGfapajljNyQ5Qxe6YPFCUPjT5Xkvx/dz+S/vJeH2u4RIvkgsFAlU
AZzXG2wcv0kFo11kFJHiJQM5jI6gdc4djH/pntnBzY9XovgyZRk/TAXvKVGLTX8FimLtYC1wzosO
bvAbtiHy7gbVD/EKTou3wxmEI9bfONwVmcmrBQIT0ChjrcV9xaFWPhvywNq2q7Zm4SEllfDQd5Sh
Yob3F6EqhckzUHCs0YUV6gnUjanO7nx2ZTLJF1OhyPfV2pK7mpXOOVw+aNq14IwqbYsh44hEa1bZ
Bbb8nYAWmvvaLwx7rrP6aeXS56sVpG659NmhrxotDGL8oAaqwQfKTP26yfHnOV8MeRke41oRsVTW
FQTQe/pikINzsv8oFHZZHSP7pGTWNsy8fAhAiEEK1w7vFW+1Um5TL1TJC/eRwaKE18PGCPfRsQyx
kkyT818pqE88t28KTItDdN07XvgwXP+aZS/E/J0TkxJrbfVcMAG9Icen7NModJ3ge+EbxMadsCrz
3P4w5nQTS2kpxJCa0dFFgavnw26gt4AKGrPBPVrbIpwv+eh7Dt0r7+PJAypocyStvTkhP/dZ16kN
RrxYcPCoa9I+8ANqJjHuAHMJkjI09908r0zV3a0RvTkKzlvm5KzLGue0Znk1I6GCoU12DTbpBz2Y
cHZykDJxA4wYcvDyIYFPw5CU3oqtxIBTC7Hlnu/sTmWJY1vEKmWxAGQ8hwZyqLWv6Td2EwbYSjLf
F4Q+lhsXNvQdMZMbNJ+S5QHaF6i7/OJo/FgagsKjNBdiYVmXPnOqTPYAwjeEVa9+UmjPD9lM/Eyl
4bjlGGcz2cSfgdHi1X9nASsOj1wPp7uL35IH/84JTuXCTtLLQxVTTee4ZnCXIl9A026F9YC4lG7M
lAimj5psKx7qq2aC9x18oSoFtmyjETlVP7Z2M6ZXRZ8jtplEEnfkI236FdnfIjcMxZs6uHJ94YWQ
Voh7SvHqNvcfpuY26BmdKdEf9p+qTv2UrcYNQS1mlRDB2oEkLt+VY1UH/6adZFh/GthvTXuHlQt3
EpJEzZfDqr/r4nxhuyQP/rYHuzGiT4YNJrr/mmO7Krqd2DEdBJqm/coRl+8qhmEiy0TBmpRGBMlI
GCssvPuNsUlNkfpT+yzN/lbzK/EIhAsKsgDrdbVdRZGkR6SqNsC+KMQMWGNW1qsxG5D0DPd3rb4p
RLvPUFLBHjMep9oTC4dtdCYZdDpMQGSUib6MZhpnHqAzUJclFgkJvDz1Xx62oGt05mJfL8GsTLjf
RzkcSVxv7jN5YtFtz0Z3J4/iJoI1dlANdQRR+yG1iY0CknQSUZL4GJi678EFblgfy6KtoCchQM7x
24I1JnVq7VwHonfQ/vJIMHQW/7cxWSFc9h/uGqP4ywRJldqSkd1wgpsODIK6LL4pSib8llWAaTo7
0Xuo9RVbmeiL2q6+mpgSrGDEbMgg6uu9e8AiJLk3hjEmYm9J+7fISQabQwbWMD5g0BUdV8OYfX/P
j2u50J0zuNv7FF3yXlApGqmRH2hBnk0AwBpWEFFueFsTStrExxYovPvt2OxN6ND5pwMR9NKYTtLc
Ey+LJOqBswBCb/Xk+unNawYn1H3NVLFQh2SqhycihOCr9SEEKaWVPcVSX7lh6tNxx3fkwQkMnYEQ
81FajRWYXN/i6+fHvmEKB6OxH2lBweUzDyWkUAlJsykG+IaASf7QYzE/IFJGm9QnBSl3o+RFLXf2
mgKx31nCfXI5w5RcpttFRZjRwfCQc7mi6M/dxZ7yMtwKt4QI3XWsC75ciQIOAi/+FQe7bLNTU0Ue
BuwDaTNtiSM3tjAfFgyl3FMbMpGOWaoQIJ4oosnZovLFdpoSYNcetWSC/4HrUXWNlPuqp7SHVUZH
qt5ZzVqOL7iYgU3bPg6bfwl2iirPKrdegSf0urNwKMeGEj0VjxGnQoSiAJ8iKFqtkiTUjkrkaOFg
kgdfJZhD6Dn/H5edLUu7Gfh6eTzY3Ost6EOqKYXTN0lHRT+JUQ/KwoIk7LW1bLcmo0zUhOepQ9Cf
sAfMBxxjLl8nFiKZBFBNZRrm+L2vJ5K1i+GtjoVnZEh95GkXpFnwTY3cliyyVdtEplKNhJUiQTge
VkyObHir0g/KnX3vIV83xU12cy217bECB/6kca6XFEJT+7btu9MQMX3VEEu8qRmSzERnr3pfty/D
Q2eX7/+boNKKZ1k/MWBT4BppwnrMxsRKOK7rLuRre/hdQPaXiJDcsrc235THozupIOxzv2NH80ug
eJJw8FpbYQ0tOY/3RDVej1EEFeoX8BsxsxmHtgDn/4K0xhAkkbHezJ2G0qsZiQDkC7TRydgge6vq
pJpoqnLDLf6SIphq/TFsq4Kh1KZ5bjKq9rhBE0GUbFrFE+b++CEC9fICDC1dZTEN93bDkmVIGq78
/t1wVEJaUGUZ/SX+e1HmAJgRD23zF+2K3PvApMtYLNAZPRiIG22c5JWe3hCGkcDULFse+jJjhqk0
luqdwaglGnPXGHEQkkWR+hcE8hiSstRoAVO3MZbYaw4uh/RlIN7Sk4kkPcnH40THP3kJ+X30a9wT
uFAe6VM7TZ3UP2+OuI6CO1K5WxNbCYfnaIcxkVHiJOsK1K5KOTsvUgX9SrJCDcrYEB16i7M7I/Jx
ylzPrLOOhRQyog/b35vwVLc13D2oOcA2YOluYVjsTQawP505BOSXT6y/dgbhRP4j2kpWYyAdnvP0
5LcYs3Drg+rt/glqZuVwHgcUHlGFeo29XCB7Giz2VZAlHafTj/DmGvVM7vKbJwTWExbPSzK1VJAx
g9A7tb4M5I73NXmZ3lR1cJkgQFzE+QgRC+shs9yo25SoNc9rJiP4QO7E40676KARaxMRDbFXILqP
3fw5o03yB2R/weYC4SXcJYSzYjTsqPBVT0mt6vAkDHZuMELLs+7mPxcFYGAYJPLeDtwD32WmCXI5
Bu2RGVV6Xfef6ASkeu2kapZCXIMHhCqai00hPmZxRYuUHCyRlpAAcosfZmLFpDoUeeht8hQVFT/R
BWa2QrG0lSzNB6rLyM9nQyjWFT6fg3u+H8NF7HXtcGjrr0QU3QzzvgOWxAu3Kz4ep7SanvXiOWNY
7m1ZskTGfZvfytsvCh35ZbDN2bpGLynMUCfqP97NfZgU9Jt9OJj3bf70Iu0ZEOxJsxxjYBXrs0IY
aZgqep2vaarOq5m83kOW00x9SOJNEnnzDJ4VtNJa2GiBlUPMaOkEp7P8yuVDIM9995g3RSE+sWpI
ZV0NKVozX0GPcM1WbYiVHFGOQqiMOfnZOwrGLYMwdsJY5EvAbzw8+QFEBZR7zK/vtApJSzrklXdH
S2CQTVISZyTdeZyWiWAo2Nzb51/K6fzelrAYRieCz0qWJwYQStgEUYlNDhnBtipPOkSqyR1uw0be
sIAe4W1VbPolVZx+ji7DAyGPnm4AUiecnQZSKT0RegnsNdRtCgCa33iifdlpuckaD8zcmDBUAabn
IZQhMhRxG7wDGQS5rIvyI+5i2lEC7qRwhi0dM5ZEFvNFhEaOwjUFWuNqVU1u+d1sYRqM40LuvVS/
119HVK/GmU0RY75mI+61/SSUC9FScph8lUwPoFHgcc6VowiuSSNMtLDLh+NllPI/hFTyYoAl2PGm
QnKySeqk1BZXPUUFt1ebEgFFA/Jm/y1HwBNDcpobFRziKx6S26WHLX7KCej8657p7dqjyG/0J0OB
UVpbeCuhwoYcIUIUnglZeb3vNIn1jRxdYWhVLhP8oPEqKVp9WlEg75vb2zOC4UMzZ+z+9plm57BD
9Tb41G/EclTOGEEd9HMa4aQPCdqf0+UMfA2/BmhqzKD2eVh+XnvIU40VQYaWH+gP2NI+5Oy0KvHj
Rbj9suYyfZwQURjf39oWLjG17OWlkUyGsnXKJqLnWcVvsYVHPya6B3Cyi0n1IHwk0MsvLh38G+Rb
HrjxG9SOGqZKiMzEkGnKfb1eE9QnFzQj/R5Ivlp4V+BF2oB6rE8719wa5ROvn63OM3kxwBiNUOig
J6cOdWTFOfWMji3UOzuJLWWCWOYCGrCXsdh+tkkPJrJnHPR7zirYCiKte9/KN6tdlTwNfGOtb/IY
JgQ3GH0m9WXO1jn/UGLQRbzVaM94PwX2YjTnagelNJMCnIumBa22R4lSg1LNGL6ZeVdFk3eRl3Zn
8zrH2qfeuqQTp4zNjVoGmiSze5Irf4vpynZqYUAhSqYWcTFGUk76vBTXN5EYWhpGkETMrhtTmgfr
Bm6UgP1GgvbfooCQRVi5e8nZcKNFXHecGo52KDgKikgRRfIu+ha8xT/8g4Bw5hhYMHIfyXshWZiH
Aieho9HG0UzyVylwn3a6QOs0q0XGyW0F6/wXs3NslnEXdAsdBHEcJiEZfvvFh+I9/pT6lSzP3ulE
NaX6Ok+5xc9ukr6J0oA0fFshvBfNX/htl2fkZwREgWa7qXAsXKlFd/mNGz/+qkpwRObyv+mu1tBh
L5zPsS6Vr1Bp/WNd3QiWnFiZNcWLXuNVghhU2m+MZPY5amyNUdkU69NOKCxak9XQrp9VWAD7j9ZK
0C8AF29qixPrAiGzaXRFSYJhCcoIVkA34IgL9+ObWPp9SMHPcM4nnlhe1BABA+Q+frZogKvGbPQM
0M5RNtFqJVmXxIsTn9mFJ1XWUCY5KWX3gNaV/zdkaXoZWYm5Kwb9s989p1t5FU1qhZ6LpUeaVcnu
HX9homBnHd2OazlvOyopxj5q77BkHoPh4MrVK4ecip3/DUTZdRi09nc9dvpQJeqECSQmL+ylwIv2
aIyrhqzBo8Qtb6ulawq/u/K3n8+aGazAQ0TDwyiElauGYreYlSkoS8IJZJmMnZQkaqTL2ojW+Clr
FnmLky0Dbam+B8ixxxu3g6DkACUrYRQaJ5LdO/aA+dL1sj+QVk07YJPnw8wi/bqRaewOHZBZSfel
OCjvxTYj3iJbKMHHVRniJc0SDxQn0/H8J28U7aSo6FyqfzBTVFf5D1GJu1FPr2vYHjipTpkF2/sv
yQCDM9xSXw5eRGOInT4NtYU9jt9xaLSs7OUk6Viz+c+HU4LDGvdyamwqMj06Audfh9TByEw2ph6z
nm/qlYRaYf8iZWV/htv4dObE1QVQkbLNLtxdOY7ebJ9K1XkMFt5zTk9WtSI8i88l+0IRj5HdsbtF
oAeocH6aTNCzXkC3zzNIrzDMmw6gMwENllOAiQiHHYHnnlS3YwaEAc16Z3d2xtNFux7aevBshYB4
4RCubHmGrtBdun7w0BaU4djLgtADI2Z3KgtfN4uETpSPuv3gpYKRby9PzbHgW5yNeP5Mpc6hqLu8
kcWEIbwDhhH4V+i7uRk2RxmTHNZ4GiQirGrI6OaJzS6x4PutP9JUk1ngvL3yWygF883TN02Ym6yQ
zEpu0XBlg7ehEGkfQfwQHyDukzzpaWxy7EM6WtasLbekYIQBDnXlk4FjcqtyX/epVaO5GulRmH8F
Lamir8PZ0dUT7jTSVI4hmVyAoTKNhm605mTTO7NSEviK8lKFY659UXUXp2K6IEYxiV8Mrc4H+muL
b0RhIoVfsBZi2reJFCage5iSnl21QQSjVBXzzF/aGyTHmEY1jBJqGeKLJjaadW/V12GsobVxYNhY
wtq/HKmhDGhsDJvOtuOWtTusRlBomlhQeknQ2bIjN32BQDZ45eB25NdFNGyp09gt0sYikPN36wHS
Br6YC0KAM5uqmY3t5eLCYMh5Utl8jvD3OQ9bUsAsvhSfuXLDj1LITRVfnWGm9d3xU2rso29eTqlx
oLKnBp6PoOcnEqptwtzBPCD3+A95cF57ojNywI/P6IpxftQmVh+Jbqxyu9aL5kNEP6exvgx9/ZBO
Ut+XBcrtHcXLGD9v/jQZ5nc8yynEPjyS4ek6fsVcup4fDDAGs9FWhqgWt8BITcDCM3eZR6arXQMR
5TsRM4E2jSLkoP68YzfnPReRlc5YrPQvC6ESMqi6pBYdAQMSobbTebRXdVxikppT9DQtSfQevRTB
G6SgOkSjqRoKJdlimLh1dP/8kwhyoQRvS8QfY3TetwGQUzHVAsjiu+rfORWvm7Rrv+JYbtuZaa5S
QZ+JMM7IS3ltUlzoo8TM7chhhnMlmaKYQ5kc12RvSOy3YQrOvCs8x/NqQUysKuYR1dC9pp54lB+M
ucr0HgB7IwYDC2NUCaPDiLKGZ8Vn85QgG+3Kwg8JUz9QXtRyUHB5ru85GRcEtKYlvGHzJ8901J8q
a4keU/FoHWLVxlxypS01hpzRMS3s75xmk6TJa8a2gvBMdZjdKga02O1pWYjavVw4LxodCYmQnvL7
TVFL88q1ho1/FrMFOKH0NTqTZ7BCNak9SK6RL1Xi0+gVeWnzTYaE9QD2LD4xNAajj4D/5yGtj3TY
AMnRDFks7eyW+rhIFtnHqpundnCxgnkdxjW2xGB0BfTl148d1odb0McGz7vpbv+Tp8Q2JzSFItKz
lQ7vud6Kk1aoUeYjeDYyoqArAlmbA6wsB56pXA8nC9orPA+ag1vxaQCDgxFn0NYOGpOd3z32iPc1
9xP2ZKM5rudg4TA3l0YqTu6F3iu2/WPulcPwiauee4UWF62QdkjjOvTXRWeTz/lYzLIhNi9K80Jq
lI1Ep2yJcRQ/OylCybPner0fv4ale2enH8jCpEdyqVabrNv0SDgHeQSh9hWeRQHe47k17do6AMln
o3FRCv1rqUZ1v/z8Qk3NTLGExj+pq5lT0aQe+IFz4yDM+wEwO2vs3Owor/bo6w4h68f/fpHVqjgi
u2yw2R0NsF02Ge9g9z6zwH3tmE7I/YQIP1+YhPOpkbx/uKf0RuskdJAF7oqYZPwBL7XYywUyvFyP
xLbNPHJLrx98qOv6XlDX7xcLPBjmY1Uy/CvBSx+jPzRRxXPVkdA/PRCdzStorEqBaTPzE18fMoJR
oy9C4f682qCY/iJp8NPiN9nQ6vKgZsAa983LoyAzjbqkEOY5LkNnxLNAL6ysTnV5w4WXRt09UKhB
q0y8DQkSms9RXZ3vBV+6i3z9JS6KMsGKRFOYKQjalprdBDB5m9W0MYnQBj3PtdT+s7+bRQ3B4LOZ
UTreCzFjT6+y4WeorPJRmpoiqBzRZbZ4pzNFv62bisjNzLq5+BTzZ1TEUitZYZ1Xjyaytm1ITvf5
/jv8SEe9PwqUsVMDdS6ZdtdIJFNroh9DuMgXJqhhf/wQFgayWZSv3ykJW38T1NCodlxhi5YODXeI
rEzYi0zSnL58X6Ucq832AWhr2VMIwxrMR3M+vyzJPjc+2J8dFX+MLtW8XFQy+Pj6p/0gyGDMZvVD
E5Ba/obB4yZzkdq0w9ReAF9zAYIGTOf4zoiMdjp17f1nkiiVGO9IMrp4eJO24Cjydms0n00c3gYp
Q8RIjDF2DNgdNhRv/sQo4aFYTOQhz9G3t9exWv1OZD7xu2YZd3ZZ6g7I4guHwwN/nvdhVolDYQ+g
7+5iCNYjqaleuso27oKxcbItQftWsCUb+IfplDr4OJJ2oumY/TaKcLeU7S3XRnAqBOCxTTLISfc5
fED6RtUI5tq/1/n4+DFd5sLSYSZTPKBp5wxoFp8FWNnxuXInHAirc4fb8yhgC/NUoaxT2a98eDEw
L+vCpfv+ResmfP7iNrzQi+kFTZO/Wbye8dOz0EazF7oIpw/w7FCqEQ9YE7nlFqViX6s0lYnTT5BV
OY0e1Q17nmUHf5//kDMzAuSII6fmoV5BzwkddFMsUWtOAVSS5/tJTWDOoY59H00VaDaTQ+fcThPW
KNItfb4r8OsjV+AxoWSHj+FXLHTwquK/NXLuWpRhg95iJr3b4NKrepng2D9ItXbZ4OvuPcdFTzY7
PQBsXMJD3Q/qtGpHamkZ5Oopc2OJA6FmqmvYgdllPF0QRKPf0TwmE9AT+lXKn3hTG0r7Vcl0uTR1
0nm0eB+HtN8+LzTi0t3pMWtnmrmhSv7mWei+UlcvyO8LwyizJQm/G6cuf+afA55xZNndo+jXfq4b
X+49/+i0dajLy7jOi1lfOmfm/yu3BmAGD010JqFAZKMIycm8IaS6cCSirVLTfZpKft9b/W6ZwLS9
cxllFkf1AtOcfGD7qP+jE+VZwVOIK63FXbM4UrOhL37I3RdzgnWQaaeX8x4dEuLoWnex/4ik+amc
DkkjHu57WvYssfJolLrMzIw7A8FFwdyAzEoDa7JdJyE7jalID4SdpmcfWOjL1t9jArAmFInyzGfa
O7e9T1ZvnNkWB6SIW0Gf9zRPuV9s7zJ7UAerxABomaw9rf3wteXG2UbwqyPcjfM6GbOKDxVmP2yW
at9tg0MMBRd04RZaG0pxHMgKqrAZT9p+BHe40O2EObZGrXTIuBRJLxQliqPO/J0oWzeGowYNW8X+
Ih6Hok0BW457hZlQj5w6lxJMQtkAaqBYQqNarOujyLkP/2gngENHOUY0hJRCrhrzAyeXMwD+R/gE
HrQUrlmUK5BvXyMLvvJQ2YTrTOOSAg+JR5ifCIC7za6PGg4uR8NNMKFNWGvckQCubHbRHqbJ0gxa
F+g/ZfKmMP9SQpb8T0PA3z67GWARcAavr02dMbGAkgs9Z9MXc8VzgQxzzfYgSCApJ3bq5nNUazQt
HB6hZRon6o0Q3lsvYXljzzYSChKgjVyKO+3cX+zH0pLYjk+dNyn6FJTcDJRpQ3+z1ER8CFC/Maxi
qZH5S9Q2OETEXs9AEDKCA90yl5ffvcJRnFeFER7KxGNwwWkRI88oht2rKsbYZ6tKNRTMJBkXCkEF
rIlpqhQv05+0EkCIXR38hY5IQo8YqMUWTmWTTVQt2B4FBa52HA9nqaBBSEPnI0063rtnwzLuPvym
+QDBZDSmD7yrp3vPfdAQaWS4qVV8EhyWn3OW0DttrD9Amhn9sFPMLdygtmZO13ukWHgTnUoZqYp3
p1U7AOyvwmnSGZ2kuG2PzG1b/RfZrgyFtkc+84tyeK6AQc0AurD9d1CVRyYCflHMCSTovcqf6RwV
2AffghfhAOPdw1lipFNcLL3MjAzpUljXu8SKAuiTsk29M53CRnOnwc094M0HjTJ3iRw2vqFGUmMj
Zykt4npx/TAxJlUgm1bxyC6/G95AWLEksRFnvUHIBQkTPG2jaUL7r7cg6xMVYH5adT14Jpd5eDXA
EvNy0Lm9J2tTGrt15q+pMhTlv6IDelq6ZlhNtvjBRg6A3SvlSIQOMbPovobcl8+rGE2LzlAEIit1
rz00QPSfvg8Ny5zhH7bT+OzraPTQJyU3CLSeIJvg7/+0I1l+yj+RGXQ7PAP/l05tYNzBuwTf7DCJ
Rfjb0Zpgg92KlY9LSpVt/FtOZgLu8GRZKdIQEg3RXv2VTnqJu7hWr/SeUldtXi4XkzZGDQ+Dqen1
foxrRWy9nRf3/4L3eZeDoNnFZQfPFjjopv9KCbBZyuMIGdYDXSKnbiLPnB5wPu2qumIircf7V7HN
CTTtEH08R/z6aJsCh+U7azLZ5aw3V145o6T2o6qQWWsstyIivHTKbTIJeCMQUbSZtGQ1iimDfjuW
PY9jU/pn6SA3pGes0TAz8MF7SWk2VIeA5uXo9Q8JgOOc1SbSkq49QFpyDyk8Txg+bUZtHMXUpXVH
FeSFdhfSmF74Dok6aLPD++lepKSkg9PGqgwVhyeF7mBeaPKukWRntQxbyb0logVV8Pi1LX5yS+RO
Ogcmx7Y7hp3FevQ0ilmMxvyRmv78FeLUCZ0Vfb8E3meB0p1ScGaKb9IdWd1HsE71xXjnXPk8LCai
7lj8xCquqc1KYOGehiMZMSbwtIus/v55cPwVMRpcYvdU0/y2Bn4y4qAcKZLkc/HzJOVZ9bf6Wsj/
jvKCAJt9VjdPsd7Ga7nOV53hbvJkP0ZJhaPc3KDbgsLu8uQAKu0gsNPp1X6dPfz8B+LoZUVVcNdB
cN95CTMwNJC6kCMGxRC+/HDg2JCz3vTPATvMG0vXL2A/joJRcN0xHjx2H9CCqg44Ni/6MNnPhkTc
T4swzdtO1EZuQn+rMRXVG2G3Hbstw2+Gm6TgTmznsGaMq14LloC6+v5BsJZDeRazz7it3ryviskE
rOG3WEATdSRAxMoGC46BVU80BzUYd08BkWTIWGpXfIDyqNP+7xCpGz+b9zVmz2DPulAldX7bHpO7
0eJoOADI2kzwsFyqfmCgusCoDyLsZhhPXulPkAKLmJxYfttvJVMJiqovgexdRTzENGRsEFR6scEH
D9nzTfJQDPv6M2tnEZC8zDX4y2cyitsbxDJu0bRIWVQKmQabGaf0Xkh8a9S60pHd5flv7NBeU8DT
L8u/ZEx2lW8NHqdxPids0Z53M/HZKp6S/1Cf5gcgcvaOxOCkp0bOVWN383dMYNBcDSYW8hGMU35z
TJS1u34gz3YUrrPGQnQdACFYZ5CLdgr+a72CQKwmHMxSqp2osLCXxQ7YaHRvkqTzkVcJD4i69PYt
7Yut5vnq16UFS28/rHP4oCPhJlocauiVxOBQi9v+HiWk7KQifM9ED/T3et4ruGh9clTxnuEtHwg9
qlbcyAj+eMO2USwWLo62kzVuM8FCapYXsy4NKiDtCrcbKLgprPQsrc9Yy9SxOmeciSGMP5prZWst
TP/vH+Lf4x7HE9spcZB+Bsld+ApiGK810z0/t7KgCXE5EcKzxP0YF+V97h9rESJm/qUjCenPGcWj
zK8KfnSK6pUJ/UR/Q0M0EfA9ow1N9HnL0OVCPduZ/U0YaomOV8godeDx0iHwErTrM8HH1T5VDSTS
wIDB7JKLcHb39uFUiWBzxqrKQhaMoiQeJ3r7v8SSOSM/w1SFs5+aRVzsE6+7o5lanhyeZERufM4N
cE/8kgm7duhpQ6afSWDs69egqIYFDySHu2Oq/7QsuswLKYFZYHnkPpN2zBiSpM8xWqSOTm9ayBPe
+gUDurvOcSKb40H8EpVU69MkdaBi5TbfK1dUtTn0ZlIeil9BOCTIuMWGwXJRzAa4KQL2Ktj8/hTy
iC4hWJlD0HDrWrXaIE76GhfT+kOLIUedK47ME/jpoLBcyO+LVHC/r6quPSlKca+xdQmT2DyItaX4
lESgslUYMpHe9H8HPEbVzx62B8F4yvDNDncrcQWfwLeOnX1xcANKFCoZtE3COYsYcpObAlcQoj19
MOtjGfcIF0PEXg+7Tor6DWVnEiutOdYmpJvaqXgLZ5nACXYAjPt78eyVaSfNBdoqXIM6G1fpMD0C
nTKyIxf/KkD5rA4aLWdFYnNb7VsZrYjJ9oMKAWQ1gRJePyqZI1s/QM6HnvVvNyFd1Z+jAFi86NwL
Yg3M7tCHD9PU0OLeSuGHzM04fERcq5IPkNeJf3HsBe1MchhIlcBllogrqKejlTm3O9g9HF9bLh1g
hBDJUCi/ImNVJIxVl9t2rw0GOlrFezBP3gnXXxVZl3rVJKvmoe0B8A0K18naulK2STXXVGxXxXE8
31cuIJAdK8KnQTp9y1aETvz6lDw2cFZI5K+93GHiPIVl0RLWUaBhEYFSfgApIZ6FxW+Ce0JqlliD
OonWyaTKop+ZsUDbjqV56fLG/a1aWBnsk0PUi67gvJ9dpxDZyppPZcJtqMq138owpAWvVo64/dK0
jYHDJXuf14Z3D/qWenvEJ4392oADdF+MYnWWTvN5CWYAtXfPkWf7NscE9iWTPs5ySvtPkpj9NBvQ
U0Vydx97S6lbW97z32xws7F5+9+n1PEbuVHiUEEps15RDjnWW1ZGxxSF3psPy7t+wyWhg0Bc3spV
KaZa1jon9Hs9yIPDQ8/gNcnPZw1FGQzvMEv48W74RkvjJ7AKtNPLZSB5/w4TqGFe4LYrPIUCz8s0
lSj/t2+1dYRbJiEQVsYcLiWSG9aQ1hj7UcTSUF6ksZ4L+ve5U1FRg8nScndbPMAyT82XQGVA9zqY
igyGLD0xClthQcm58T/RnJazNmq0JCEHJBzV9mU6EyY1dYaBWpxQT5akOdXNG0Pvn5GAthwqVL2e
d8XneUQx8T7RDE3p+296YtdkGEEEuJj5m8pOjBcLXsz0s69ST7Yzg+DUyR9tBVpbOebiCYx1H12L
9TLeUrnVAI1iHTvw5L95llPAkLEHLZRYZJr4bsSl/ybbiy3YUvyT63tZk0VI+PT5UNKYPYJ2uV+R
w0WRi3sZQ+sSXitH4FJgdF7f5fpiCMUd6dcDRwvE7/VY0UJLgLgfrLXOPXb1d/6XtSQ9zlm0sqv7
4y9/HsV5veolZOa9MdwN12227QFYixKoI9Y8TIQ9lkXz6b/2ue96xKG2blbhJN97EjDMYX12IxRK
502g/p108Z3xU+eHIc44RhGaROg+Iv6S0fLg4Mni4Og9GEMmJe502Itfcycu/PQAuq9sOoFv0sb6
E61jCZx6vIUpKOXGxjPj0zLqlAL8JgMPM7L4BukNdHundejAXlxzUvrTCafQk/cKZ+e21nRPQqfs
j+XQK4KN6AwVvkpaxhQgm6Yc7Cp1wIq7E0r7tN9GmGTgSbaBrzc6VNVChDZr2w1yEGArR/rh+wpS
AY0GJyMcOJTDQ0tvEaZiJ3gnSKuZygFUEaxoSkT70YcutBSuEHL2d+ZxbsoBGjomPQB2wfPi1z47
KxpG3qY2HIzACmn4zyaqXxuykRPUfTPWaTP1d0+MCzX6mQDGtwvkBndHTAKTCjKVziIZUXgPScFA
oyJg70uzyPF4RLt1zqtrwXbjWUUiuzyerdI1fmkNZKifRPK63GtH+Z2f+IhCP7Rx1UfWSp0P/o6a
1RVpuAxK6pUyXWgLW8e99+e9fNIYkk5o1wShPv7RGoRJM5lcHVHPbiSlS0OIpz99ZVIdkGHd+t7r
YdaBBxBSjG8/0GdKuXNvnuJhv6bsHUMHN27UwasA0aJeSTWPDg73tbq8zlzFip29KqhF/K8G4/+O
AeioF88j4DnSJRk15M9m6Ha8rV9SW1v2QHU6J7+FDmUnKVoUg/VJ7ohM3gv8cPwVQGVYvhKa9oSk
Jv05mx/3Prj5N/Fs1ltt5AA09moJ+CxOk7R6azhvFv/nCYm3iliYE1/FyUN5Dfnuy0WTxFYdKKB3
5YtWRBTZVnDFef4r9GxYbwerFCepsS5AsaVhAb0fskxWaintbVEXwJyXNOf9eKrHZDdKJxkcFFn+
YNocPwt3pIrEVjrvV6MQOMoe8dejUcL3bspGZmFFQDlGjZhcLHHeoPzXhgijyGSDYjjLG5xYxHKN
Ca+573cb1AK9sXtmYudcCHARAKwxw0FBl/LP+l4UjmlxIKHeAfv7HWoxU8vKEyzRBGnBZXcij8bQ
apLqMJkfg9cxqRXW0iSFyhyJ7fS7Z+kNveOgQDUMNF4kEIW24fH1miDzbvxJr3wbrKNdm5fwkKj3
/g9cJ9Ty5eIcBvtI4n9Jg8ATb2mhb62ljTZ7+PED2AIL8V+9F+gDnpsDIiwORxNhiS3bqJh2pxus
EgW77Fe1dchE/va2oTFC45/HcndkFPoXu6DyvBlT3QlIxFxCXNy2VDdb5pQFOlO2ye8G6HVS8e0O
bQtto5cWT+sS635EZFI+7I8xosITHhQscspChEO5ouRyQVsuwM0bM+dv4e6SiNtMQexBnMkI9S+s
5w7KC223YhedubwC4Hweq5xWtKzGTSuxw/Wv5K8lMBAshWyVoYvlFuZvhlrJuoRdbSqa/fyKmjIr
WMIgavOJmVlovjLZiq4dZjihtvg/Se6EypNYgLhm8p9aoAscA15+SGkGY3sOI+/mT72hmiyx17Ai
muL63/7EVwRiEnQKiui8yp2LsJeaRtTu7ww3VXMnCa9zE6lWs4QIxNra6Q3KXVr41h8pzA478twX
Kb3Lro/zjaVOSPu5SXz9iQA+IXRLcq4ABPeM0Hk4INV2x6IBChxjK0t0tRP8sxWGByW3hq7w4hR7
vO/EGWy0MnLMlPizYiY/TEWM8hEQxmTWwMdv6RVj2vO3o6YhDQMeAx3L0LpOmm0gGu3dQLNazhww
8AZ6MyEUhOHNSUKORjb1xIxwb4Ti4adcj+6usCBU/tYkCqy86zIeug5aMRCzQSANJcF7dfA+LwPN
HHvDQ9g5GQxfbV6cGonBzolHZElRu9t2qbfdtco7gi75aYz4escQCEPftsqBr7NuP46XsD28ccrF
XbzZL2+PXUw8lhMue6pWy1idOHR4wBIyTyBMhVS7jJ9NvFOFiMqN4j+xWUC7xzVNTLj2oKLxAEBY
Yz+c1NU9cbrFF0+OQTKw1/ZdxgA5/QzfB/FlX340DST5PLRXNBowNoUMbX2d8K7voo1linoECeik
O+9EHz7ZoxlVk4WVPESMnguciQwTDopd/dem3n5qW48ACBSmQVGSv4TEdukSm8haEChxRqLuBMP1
IcegkMbB1ZZFIgHrYUfxyQIAH4y7DTfwoJlR4GJVPEq3RTvW+QLMikvlPz7ZJqei69faLI5lL5cO
VT29f25D+uroE+++ig/IZy+XOOXbQxjyeytWkdTLvbEa0I/Fd1HUKIdnpX3MQzBWZwk0CCJ1Wss8
aC1ZjNqzE/UzioyHgM7HjH2eQWJ8jmT86SVcuk2Bh0SLfwhwdjoK3+ICmhxV4AFPvQgYIUqPRq54
pW+pRa/+VYIue1wIDRrKzPXyLfjRYggpyjV0vBLMxXjpWubGpOIe215lyj1EZGPxBzaa6tXkQYdr
3R2GoD8x7i876BQ6rYRdKEy8X36BJfeABSzPPzDABSMS4g0v+bxOMNkWM0Lqm6XPeVVglJIUX+ma
Xp3blPCvyxMUuq6KOyjrRpWPGcWKGs91RYZvW7RB7U4PThuKwkt66MJNqvRhP/AOb1BSYRgBK7tP
fXUNo5k147lRskN+TMi1FS6BpqfCo5R10P3TSBJZToUEgkjM1ONtQsJgTVyYXpRcT6KTv9AHXcxA
Z1XPw0njz7m46IfR4G1B+UWN25wa4qlsd5L5D71dGyMOezwHWvRPxLKylNw1f9H7FW4CiBAUQFkA
0/1PURmyZxvGZ6gQAYmH4Bj16L61VVqOMVhYkXo/je8tVdSIbrl/Yam0jpneYU5yKaEmzALAOZwJ
im94oq9FihLVJgVUxQFuKRN+CL8sE90pf0XcoBlIwhc4Ou3LORa4Y1BrXFxK85i6EHcKPMzosUTo
nOASf1JmtQx/d1oYHRHnb2pirkHtKcndYLLEkiGtQvNPprTtoS3LFhbyWEWh+7bSHs2Ydo1Xb0V3
VNUFsNG9Ujb19a17aR8Ql8WdzuXAk6jYjlE0qtAUGpNgAsCFjT4v6mW/dgsceJlI9uMwHkAEFua9
q47qsu1jYbB9/tMF2RPabsmsQhiY2diMiV3GLTqQtqV2pk8f0Sku1Jo6/Vnp/ujTQKKBCVMI4Mbd
m25k4EV5Yws6KIynzJVGuUT45j9kjvVBAUSGMfUwv8OZDPz+3jas7CC/I1izYJ3ACfsD6f9Ae1UX
lmGNXXvSWjRQIGzwTPolnY4GhCuQH9Sb0cU8j87HmWBZSS35F8TK+P5z6ThM/01BbqRytFmAU2N8
vbUgomAsu+KuNlTSqVsOYTVEoO6J0KMQ6w07aAlcoqyzI1UJUjCEAA2eDe2G3D9Jk+hIfiTZuHCL
9RZyrkUbmmYuIkZ9FnMSOtm0h2rs+ICdR/4W11CBUfs17OMOOcL5ERIXc/L07TtV8eZQdRNbYxYx
o6nJvKT0Hr07dEybhVGoEwlv/XQVzFGw1IwYdJ5ZZ5ywpW+bQ3gy6N7YCuPydcifm/SvN/apz5EB
w8c8NKCBMdDu5JiCnrJrj6Ca4SQf7Un8EtEQ2h51auUUcuE6/WHNQ3DVs8rNUF4IgDnhlCSRq1VB
ashpqYylRLw2H/DWlsXhf7fwIkJUyyIafF1jA0/RoqXlMryGeF3aA6VeCt85eW7ecFrcmUX7liV3
XLq5DMcR2F2NAsUrc2ASL4flNDmPpQo2mhbBCp4Ej1sQqbBgF8WPCyVESsipj0PdT0ph/rx63z2Y
EHifC/plX+LjXmapB/YkqsS7PPfUVBESWR1OBqi1J9PqdElAfmFdYHgrk/DprKDzpEOF2qo8AonO
zd3oLHE8Pd0lBsQajetyOfIYtN9EzM/O85ZDUkkS8BJOz2BMpxoh95YjxwmZ/D7rJRcUeBDmRLOX
b+5vLMt6e62OeWGfd6siUK9PhKRIK8uDopEOv/f+ysz8GXRRJCjbjtGBatI8D2k1zzmggZ6BgPhA
jIGIi33TobtpXP9gRxhyvonmIfo85bap5b4zCXif8VWsmRNLW+LwHmcRFfFjB/lYKENijtBIz+Ig
4usUstKK/ozFuM1Oi302AQaHPZemd93C5qztrMnvt27GbiqLLCW0fjOeq4ceaOK+GTfohbIpXsDZ
heRpKa08ea1Nt7W9PUcWq1LIU8RpZ5vaJeMcJsRTQlTH2EpwkafaVV4v+05izgVEXNyDtjrZWZ2Z
7T12TUh6Atd+3TCNB6LuTqcww2Pm/BSaFRcvDAHNCSFQ7Egs67EPP5FrP4CgB9WToq4xEkl4ShWK
SEqzqsSIn7GQxqghbW/sWL2wx4HrAVvs8hq9eETFUYEwG6L/8kVyqsRyV3000Mjl3VVC5R8MGRNS
eLE9o9+u1ifPE7BOoCTaUQWVs8abLbYAANG5QfuXnk/iA2yPDihjO9rpPfC7NaSFnOBnAvt91YIQ
mQxzfCl6pAZhjZQiSZjjWgXFTaZw3urZXfjR7WWrIbkrh5/nvLJ4ATP6h6DsftbdfD8+SfrG5+7z
DNYXE/PuQ4+7jnt4n+jRUG0iWO5pCAgzvSm3veR00/F2nGqn9T+L7SwgMVEmqHbThZvBvvmqQkC1
8hLT/0Ze8VoMo7KrtwH82t44GrwrEv6ukW2PgpAHwrWH5bYMMiPVI3CZ/DCYkr1VYetLMt1C+z12
bCCFzRO+MKxUNfK6WoCbth8UDHx+50b7uXiXx925PoGGWL69hJSoyam8dVtmhkgWduftlpKna58/
lwdYYsvC5DfZEs/k8NvyNET8eZv+dOFZri5whRCpWzJJESeWvegR6RaQKlxvCoxD/tophQodZm8i
3ozXY43LuMSZ7MqDZ8P+JONziwddQBocPaFt21deqq8Kojafrz6x92RK/gmwnILPgquTuU1k1yAt
QVCLs3XaQoY5N7fZ7DPcKbZfLNb3pPBc1PZMBO4uAjHxhkv2XL59rIUKNnivum7ewto7ZQ+SIhxC
CxdEdDT5kAcn0LOF/yS80oJ95hkAyAglwxP6j4W7L3ffg4kDolB09xRVSOLeo11YWTqR+hABGbVU
x3Ys7gwgG3W4DCufWnR3tXdHm/n/Zphv7P+1m0IxOjZr7WEIX8DkF0NsSls7bLh3jG7kwGLD6dJ0
hYkU6EB7ULuCw0n6qBsDyjeiHwKgBL+T7oaj/IKtFcnmJ1IIDtTyYfGMFTNA5yg92WbrecW5VGhq
4ZeNvdkr0Lsoht9kmLJG9vJ5CwKJfD5BxTOGNfZfBWLTcUo6YnYnfvN9d8pLA/oNyZUBJ9XCeZPy
Yg2UBuNALZ96lICH8+tZPIGfhlnnFe3kzJ1iysvO0iBFD3+6MwdznJrwzdeCR9oWzDwm5qY6A790
2MYmzcAx6j85v+MYzkxHW9/nR+5upZnp0ieeA8nwdgmrEUM9XWXmBNi2wcjiVryC5ZJ+WuBIL/zD
6+0nQGD+JxqEPLVFqxj5vlcv+XrywR9HT4T8X7XzBwzIcxvz5FKGU5VtwI/VG46ONkVt83bE3mTt
oK3qB+U07q8hyVJ+dI2DcP4uAbSFHrIUacf7uk+f6lzeGN8ZIjfQuIln8jGL62V2galx3rWJ0JmM
DExTLaXbgVwOEfG/lsBBgJYQVW1NRaBkvtYifQSIQOn3Yf9EL1GJP1dH5EBWqT7Gh1BdBo8GSerA
q74UHQjb+tzdKqRQrunDeUvSi7i83XiWk5pqKbndB2SUHJDhUv5i9edB9A7RlhgmrodWv0GchmCh
OV+oxoHZGHvmZ40aeklhLWa2YOJ0vhFsfsh0bVo96YtKLHROSV5PTlOR6gcI35wV8QoxSWR8ZxAt
W6gF5yODoSp35dCyEfzpPo8UYgBAkEvu3R5ff88beysIJZ0rA7S3ad0P9XXVDIASNWmDwsZhQqVs
no35Qj/9ZyPktT5IrgNmGZ8W1SGscw3D1SEc2IQb3gdgvo5cwdF+1kqzqrlBHtX+PSdNq1OJn5PC
QY0RZORxcHbYv3IYizlO/Dgk1jKnzMPOmhNya6FckfN1PF8xz9WWS4+tFGIC+k4ssNIoYK27hZu8
fPQNPk1NYZLxqGEsL2ca59yGIv2YfAsWvAu11hFLGUVEv+KO9Rvjue8Y97uQmxCd1srUtz45QbVq
5lOKATAe4dMiW5ACPrntVTmu6TPdkDbzVPE1cYfUrYczKrWWxn+lrsl9sdjiJdfPKr+hKg0cLZgV
sb9jIAzEXUBrgDdJleZanXk1Qn8ZO8Wh3AmbmKkr8aXIczizmx/vjuf++fdyQXN6vRqcYGItbT2V
lhSzRMcc3eIFupqQg1bkzt4voOKHEVD4NNswJi2GaryAMPPfs4DzAMreBMKCGr/PWPokPhZNEH5C
+PzISb3NpkaeRs+oWBMvUVqgdc6GhcZqApwAZvAosjhYQG64v9J+mxCm8mja1fU+EUsnYDiUlHoH
0SKRUckJnYPMckSxN/CqEBin5BOUOWuGyQzLbLVqn9XQeTJnlj41hkAshrACrkY+mHS2XisuG3dU
fU0EPO+3DWh1/Ra254Ob1pbh4gWDeGPtLE5kthstRknqlXmAqpsS3K3M2Lv2DlOoBG/ows+SEihn
z71Gj9V043QNR6RLTDA+1l2aeoaHjYKo3w+rhrubaNa0Pw9MUQCkl0AKyIyQ0SpcQ0SzT73oFYz2
Vm3QRkbhjPZUPsa5ZKBojWkHGw2C61rnzNmBYKhi5/5rNpkwCfzeF/M7OJua/rJswCq+FNmhXBMA
2Myq0u/b2oj0+2WCmO9wHAani0YgwiM0OgzgF24REKgYEqc02a/aec8Y4NDakcQJy+96ORPH2TZi
/B8c20cgPIdUxJMYTibE+ArvVsDjg8My7b0TBhRt0SgDg4ms7aCVlFupaDi5hLm+/YaScoDyQ0ec
kKTcImm3qAix5YXvCh3vA2D+Q9k86pLreWsQb74S9KpxgFmhWc/XzvzXUh9dhfGPFcmsARg6KFY1
Ex7Id0x5LnEMhrFf+iXbW8j3rKTWeD2ZPmUcU/ccvZZvwj4KEx2cevx+lxt4FH2+JUd6EsvsAKhx
JKbiL8rMZ57IxysmHkn+BtBZne2cZ5q7UG9xBQTJhNwVap2uvXtcFhhWU4OvdH8i4Xm/1TcQ0BD1
VFLO6hF9CP4qz8JvTLBzgnjo3iR26Fb6KZLL5GG5gyqd0MxYdy76Y5V57rJk96bAieOFzKJbxlGI
uxHXT/ULLhHVXbHuwEt8DAjTwGzWDnRb6KLQp9QGQOuGKBXXqbAjPHa99yrmrufMqryVt7zHc+wy
7moUydsisyEcsBSngxGJe9tusgVVL4PvNDw+rnGP4M+o690Jg7+nNmRR4wRqQH9fbzoXl2dqImhf
UVWCdzOlM2QqplZ1i6wJjmLVi+BcIqHvWjGxfcgwE4AZ8RCU8Tg7e5bwk8w3scaMvbgD/l7276fh
EYu42DqIGcqaNopSpmVcNMVuAyXdh90cEItJSbnzsyaYxlHL5Es9Jiuc/afqcl8RRq8TZfgHWT0D
EJ1dQwDPNOhzkg0laZz2TDU+0MoES/EHhCuCFoyChDWhV4eFir/FIr9I9ro/qi3XJOTd6lGhjf1E
qCtsfjv7pFceF2ul86+/NEIRD0NH0nrWODT1laRCMLQ9oyniqxfaZ3f/5QtuvJyvbix+o5WPD9C7
qz6FtL93aqHe/1ZXiNpMsmi/2FHQzb+Ksuj3i7rqleQ/AAGl9cE+9vTb8rblB3NQZua3Ut+t0YWW
Ll+cMAi02wnA8Q2IerXnl/MLYGcFifXFek7vNJk3H5odsRr1PZoKOD6raD0G0k5+MWCa+DjvVwxs
eXxgJZRLqWOXPwDWHwjEj9G5aDEj5iCGhZ5h2tDsbLI/mohs8hA5WIwKbkRe8uy5GRfKLitVvdr5
Y4DHgUNh924/honlfF3RTTgu+0WrZ8xgtSYLQhTP3i7er34FurWv5QOebPXJxwXv+FTENoLAmifG
fN2qKpj/0ZkjjYXobQpUWGYEH6LiMNdMWXPfys80c+Lt2PDhBaMREwB5St0wgPVNUu1iYoTjP5Fr
AP6jv8NDBKlpA5KbRC5jdRb5fNm2WP7vJ6+NDPH9JXgLWLTE0+c5kMk8/N35b08UCIW/C7a5sWlv
k7nwQuLiDePjei+RRufItEokxwSjeK6tCH1ClhKs3paEDbbieLiCg5/M/e37qp9eRE1SxXdbw0+8
1qxLXw4emOKod7K9xEdNCARLgG2Ztf0WO7i+DkDQeR2h5BXRpcsodrsinKF2TzQ0llWtxoYqh18U
TAsh+pXggVB4fwSnzD9HX76I9dpLnK8dBgxmhwxHb+ZjytBq/sz8fk6CHqVdp81+8ZtSa7PW3YJB
R6kMpF6lO65LTW+gQsh6N8igsrZCQvWcLxA6jPEK1uNKtP4N9dmSFzoCyBNN7N7B7+HdWOUIYfq2
Fwj6LDpF91Suvp7FJgyMOO71Zhc8VpD/5wTIv2EeEVb/7oGXDZbXVblwdaW5worRMRNtafifJs5m
RUu6AC2hxYf+g24vZx5PA3w0hxoKTqbGcPGVvWOmxZ33F1f12YNG6R8KuAU3U8eU7tY5u9fQg4Lo
TbnXrZj0222+2AwVvwOYrO2e9XnjU3S4HRfA/sLbCU2XF20XTKWd9nKIOtYKrFzj0KrEzaRaH+He
EeHMKk+NsWpZcQwJlzqe3MnIziNKOHWB9NgM63F1mS1ldmoC8gJa3M0IwEG7mR6A+dtzjI+IsY5r
V+YppRjM33Nv+P9RmU0i8Jno/rayA+wIOMOacSezw3dSNgXUGBn9YiwdJ1wd/OXZB34YXe2ygrFc
412vSGg6AIwxVKFn7ljndTBe+LSZ5ppYXiflHnUQgsvs7a5ozariebp117X1r5Evpd0n/hNT7h8H
nsZ0PLdDn5s9fUDu9gc+y5qlB/ERQEEnD/FloXtoRdrkD6NKBi+m0ZTnm4rSGmkVGAcb8Nnzlhk+
Hp6XFWWdSUosTO6VVmRz0s9MTJuNfqfybFZmrphEoQTXi6s7vxjQD4KYKVBXiSBNk4Eo1YN0Ws2s
sUNSreZFlG6bIQqEdUnWJYTy4L8GG06YPpY0U7kEoriCKD98Xc7RCOufPaNq0mEcNDZfSVlUhnqt
3zTepqOnP8Y19loakY/z9tGdS7m0ZyG/lvwILjTVouOxfr4Uzgsx1BJmsKOQoHWEKsc3Y7Ovnymb
4USeOeuUrOr7X8TLNuc0t55WnDSrGlyhI+LjZk6He3JC8MeWDzE84QJz5ES4gwebNWx0IO+t4uAb
14Xh3WsJOl7dYXBsVvRQNB82ltBkDlmnISDdtvHyren+adbcRkXisVTH/i+kgZqO+udIS0oMgD1h
5BR8hXspfjdZwVblifOtZww3jfG4A4ejDbGCXoAspziOwuGaGY05RBTMh4O2/WJYL3G2EiYG+Z/u
4YzDNfuwvl7bVsaMuO6ORWwu6SZ6rhzvwbVQiB8sFnATkOTF5QxhV+aBIWOF/mK/RU01GZkQsh58
90+TX4/EiYawPf8/Esg8RqL8TO4Z0nBenbpFQpXpOuTBYPNtVHmKNYY8kELR3+5WgdUoXpf8aQ+h
hHRJamEM0Xj3BvcJwRWX372UfViJWqLvFvBk4Ag08OAY30qIi3ZR8ohown4sIqaEgEeCEGBg74Rt
Yg0OyCun9eDy3T9yT8Yxv5Z/H40uTgDhcKnyWBIoIyANQ9NzREkRGz2cbGMyVkyDu/QSTgtI0dXj
soFFxkz7/VvlGelIXZjRN0n29LQ/EM8r5kF5bR2aR3w1PqK5MJ55VJ9k+fhEqbzLIJe0ddHQl/lf
R/D+0Fu1FujciGwkQaGzxUo1S3dzebB6PmQx5Kk2lfa6nO3EnPJPJBjbFmcmIHySMZ+Ui9Ds6rzV
j7v3bt2jl8r0ZtwYGCiPxVV4uxcBMG99LHmaGTU//Hb+6Z66b6aPriZ3r61FPYmPccGPfhdw1a2I
Yidw1bJRzm/BgmX63wlh0sKYCU7BYVXBu8GvHfAGb4z9fUbx+xubjpnAVefSVPvx6hipdwXLIbo5
C7ESG5LUSLRjNpO8L/tVQgqdfv5QzfwKdJP1JRhdaiUyB1q1id0Lzp1NuXjW0ECQT4NCOdrVCg+R
U6+v59DTbBzGSICFjn0/RkAwfxMlNRfF1enAGy2rQPHmi3RRqK1HyaLTP68x+38oYMlSzu1NG9+C
CAt1vF/Jk768/2SgZ4jcLOATJFYzWuh8czslPG1bzxJXUpU3Vbk8gDsGpGkLkyRQPUBp6EGpPnWx
Zyxk5JgRr2EP+LVpeRDAEs6505Lg2w91Ffdcbha6S/sTWZyFIfXOcDMjsQ8Kmn7YyZJ+4pvx6+Fr
7VWZgh8F2YgdzdaXVsSIVv/6Qm1/Le3BmwSPLYrE2BT5B2SaMY7We6QGA1mpXo1VrkyCLepnot1y
/mHJCxXP5nfuebaew9RBOGdWz/4ygZnaxBRHc6zYqXPLXApSAH8oBzzV1L18X7G+I6tkNrejftFG
J9erj1OH37vnaSq7s2oPT5IsBZwUFn/geek3/FKdmTkdvN6Y8bkkomLdLeXDjtgwAypZxIYCb3T0
Ut6lVKuPWdXJGbIHMD2tBf2RgTrRWyTB3QfpPN3bhfMgQmX2QiqCisB2nH/ryvRKCcpbgfNnsFSu
PYWIzg5EooZSkkRYX//QACywX8YQZD94UJDke+NXlLD7qEj/eNIOlgco/ZMmxG7+bW9ZaOhGtRRm
Sg/GEk/F1ozGfBp1HCKbqtpIJSuPEAOSj8H24jZ5RTqxfLUyYE4jKvhM5e4eUaxzjdEr97SHv5Ru
eyYLfLqhSfmyjCPxSPLOu/vHxiVSa5A9XBaSuYuqcrGL0aDYg68LKosYcgy7vr8ipnDo+zqH9DGS
Xt9osXChI8SrxOsEUW3zOs8pK9exzuugsJN93EzZ6ecwKUYciicPwLlDdAwKtWWSfu0fQ1mWPybE
+iCKS8BHAD1EWOKV7WQug4oCCK/IJehWifyT10llWlAFLkL4JceWyyPVmwB0PdA4xO+ZcEujY6m4
5wdm15OBOB/FYw5PCBUoCVIOyGil3IAuUEWxB47472uupJaA04e4zyZG9L2CJZy/ELXqXPOUVOX5
7xoUis/eh4/kZ/1SknijSTrb/H3CqtbTGNOQ0xAXCuFgbrGfaKg3YvM5SzBlfyhDAHvQMFqrocZW
zgX7eyfK9eKEo6iqxPcD9TVUok9+EPvxNj8eaUmr/WeJwun+NlEIgLwh3oO7Ni+f/gdrN35ihW7O
QfL/8QB5sQTPEOt3bUJbS93+Hy9X/PDCS/Wz+9eQ6+nAyxakMDL8yU4KCL2ex4JPqe/HQpJ8agJQ
CMrEb6xoCFC6h0KPWQ1XE7w9QxBTjuG/T11IIBzCyGSOleLoTmKcOfMeYjay5gQr25NIoEXyvJJX
t9q3n+vZvg8QL1/WAY0qSSRUjthIWB/oeJmhpY7qCtSqfkCw6A21BPI0mfCtji1p7eLyw+DaHf5p
UqC8c7+4qhmvAf+WhxqDQ3COjDM0qXFeUqETMTT0zFQ6B3Dk6/WzZtoNpRHA/39GWGFnmbI+e2Nd
LCDJIbbiVn5eLY1IDPtkSqk00UNZTGqyXOaG2FZfH6qAOpIAjGiZT2cMp22QcbDId6AJx4hmiTat
mhd/0YsNDjO49OickamKbofECQm5+7CdvOAWLGyHShNbQpmOtUdzzVk3xrn0j/z/fY1r0Sc++rr8
VOGmUNvhKbGeEbkrdVlSzaEw1DkYjuOJ2Wk4pkYX4RBrqnOilMkPlRAdLsd+/w1Nar5wmHBNwMtS
CH/V3MsJNExtCFUW/Lg6CLXRL7mRT+RTtYd7hmXYHKKsZlcZeRiytlsZIi5V9JMBpUBIEkL0DZLl
As+F89IVDhbPyPEK8aZotQzxzNW0SZqOEvqGXJb5qv1Wtnv1n8+2+cjcA9ndLi5sPNx0FHe9/Dp7
WH8ehxmQd6W8VfImBNTcqhICN73H49wmmqjjCyIpvmuNLAezyJhrN6uWvZ3TGQ7phvRUp8O/TIWE
cKil1lU4zp0rFwLudZpWocNIjx2HM0l5CqMZ5T83MsoVrSb/MMQX1bpoM7oJCFt8DpuM7IIezdgN
fjMCO9EwE+Z6WK7U8pn9aZQ7Mi5hKTal55YWIiW+4u/N+Z6S8NRZlktJMUtGBVztjK3mNrnDYJ1i
+jWOXH79TFyzYdjj+/gvmrMXRUXAkIqCvA4k2TJAeyQNmx4BzjTEg0p36KsYDF3VdKW0Ixu7YQV2
8zPA9/MZb2EXENbbQWyHPP946qO7UlYaNDcgnY91yQMiBJJhrThBDy0o6JArQ9dYIDCIzXYBSyid
PtbeqPgmukshOSBVUDKuDgTdxzSk4hTI49JM9RT8VxQf27QNj+cuyxLk8IisOJeZsezBJJF63ECn
fM8gnF7PoxvXVTh1wqDYg6q/HXq+POV+7kksS1CKNpvXoEVny5oR+grNsWX92khYYxRMFFYkZRZF
crnshZY0op+112iN+GCy1FLuSSKyQplmrKlJjdxrcv6gMwXeIDpf5ZGDWYjIQxplfT80Giruplwc
uPdwZjSe3raiUeJgj+JUuvp1oMN++W8D41SIfNEPkHA8Pdltnmk1+2p39JvAGTs4QTWZi4bPf+W8
fWxpv/1FwcbxiLr8YDznKzUUVm3oxZnTyk6ir4us/Q8eQCLzW6Erf5jBzl4WlDYZb9xTol+KRlig
gHCfZbHi/5bmUO30EvFM4FDPB5ZjCXpjug1RExeLgjgSChTpQx2+HGQJxuZ/EAQS9wceIYMw1jdR
q6XN7USmmVcxSm2rWNLi/pjyWruZ+efXkLUBkmlRNjOVWbqUcaVkR2vqILLGropsHyMv/SZCI6M9
FSzwiwU9FWgAEdbXpS5PDsdrQ0bpnu1NxnRJ+bvpRvXCTTq4cLlOBbYbTCjp2gUt6LqJJoRxF3b2
dSUboFGwXx3dJv181ZxeYEytNG/dUNhfObvb1BTDe0MOysnbQsw0Cq5KSCKS4IAzSleCkia/xoEm
C8EysxfXZxYF6l/XfIUtSJd/33RRsVT/rz87Hwp9KW3tuTzWJMuv/TvNzWnW2xFzLUASGyjYuRkt
ivHErKbtNHq5aQXQ/eaLjWVrUTH1PuMWyA+GmIhA0NJ9z9ayqZTyaH6F4jUjBZoGbsR1swESC2wo
zNCsmTn9bht3QH3I+lQQkvJsKt8P6Mb8tx39WDLDaLSPM9alkREcZQVS3JMckUaw0iutrmI047dZ
hEsqde38NTruhx5oLZ1ty0r4Co+iqJml0gmTMDlW32VT6C5ngQDKKjB7Rk0VAtQqn/Liuzswzc6r
Rd4lQKEkDsuUP4qQNSKfCSav/uOYvQ6s1BCzD8OZ8AL+35rLjOmgfyYttvCKoNyMpgPIWMEjJnDq
UPgLf5zJSfEQHGmt+jVC52CIiqPB63G6UiiZ/lCXvbu3pb3fyd1W1zVCMbL+QLJpWA7+LDc4aaBd
Oi5TpOSYjUpSfk7TV+ZyrsUPC30VdDzcbjc7w2SRbidNb6eO8GaZmzbGAQfiKU/kgcVVxvMGc+SQ
AUNEaX6Q6f7sJ/v699sIwdUWI/gDO5EdKxJNCX8RJWdS2rVbdnj78c6VFAUN0Cf7VuJ4W53AwXj/
Hpn0T3VBTpWdAak4nXkMS5wWfeeR/pjTEJ00vLSMqzTmuhJKGE34Jzj0nA212w8WoQgPocmKWWTI
j53MxHud3HdNxUUA87TtV8A0cX8sQI8UHGNGnaLtDzTMkEnoj2FGP/UsYOFoFTTUQ4kFnqt1CGk3
M3N3U/A5LSiO+5TGwgB0d1jBCS4VxtnmDD695UZQbAMYXkrdkc7FTiinfnaQ2yFQx3RIPU5Ilby/
aFOq/iFz7HDO35HuYRkbmUIFESjPrgwtBMwiFpVrqgJRd+sJeiMaVZ7JnxjX5wHKM30lH2k94ZmJ
SWifRp6r7lZX4Edmr1VG4haNZW4ifE+9kDMU1wp/ppDxAaVY+KTYZv3B45Gkm0tNaVbxtBjAXX51
Jww75xvuOfiPyeU2mOeqrrgi4zlwWkTTumwiSFX3i8G2FkCinCRROT5N+KW1PGysvsIHw5lluk8i
brsdEsFWixa5A/2y9skj0VdwPmsBxZM18wXxWG1FBlElOjS3xXIpXiuqowp5uEDzHSDupEjqg/sb
bVQOuQvjus5yMQ/ZDz9PP4HwIUyTotdgMPrVQ+cfKAh9LByYUHiV6mrW5Q/dmmNbbUrQvO4VvzBZ
0vxnX03uqw+5vzTWRHl5DRcBu/0Uv3vUO9ufdwRgMbcYL+5qEM1ZirlZHBKWqBqVNnJ0kjDku2Ep
pdSHTnE0C2JVcbvwnY4jO1WjHx/5uvXhd/jWxxvgndm6vmqV5gNGopZgRBNo/kr4XKryr4BwB0/Y
NuSzhB64OAmgmLEJktMf+jFz+cQXl139Xtfxh8wQb3xcj/R3shACdnRToz6uHBkmnEf+yptI7nm8
XVuonRSl/ur4jLf/DZqIeCBK36PFAS/C3UMXNgnoiJBLl6+DmARxP4pmd36kdcuIPQkVjdfsSHEQ
Qk/2d91aZSXJ9t43FvcNQEWjGtnxg5Vn37lWDlcvddgZ4dgnhC/VtrLFho1+OWWkq1SEBfg8Bgic
mkuT0bnkVxxDq+cRWVjZLgCxKcOPOyUlVz2oDJo2CI8kJGJbDPljMlo00XuVcXgW1jKoPRnOiFzk
6mZG04z0DbdorZIQ+eYKncq3HwcouQsQ7uiS0nK5bOrhBvxkd27do7Q7uCFCjFIFWlQIjQvgzgYC
+eOIGPwcd3AdwrTPknGQfTQm5vkCfDP6tltxho93iKW+NbgPJoj01zKFBdKqgyCqs/hTQivvNRBZ
BYkzb5LP6hj7ebXmzNaCq9bdfS/vvowLSj1akecbZcuoYumD8ckYLV9rm25kcwPEQ1zlem/wE4Ub
i/dzS2ZhGnWci9Q57m/PtcJjZc0r3KkOFcGM5NQpzl5Q7ilKY39wCMIu94G8Wxa6pJc0o6R6n/cR
XncUseZ0ICMsdVbYSQYl889tyx+wA52R7W6jau294/M4LmrQk1IQaSdT/bInZ9k9AUP94ou6JRo5
P/9TTk8n2DrZuHKxK+5Gaa3pOHsp295XkhZqQBZtO5mAeJRZDG+U0K+5nNqHH50LS/QWfelUdd3y
CGT+V5MMmAwEothZvc24jnTpn+OW480Z8oqR2vmMEEkQpa0SLThuI6ZYx+ag3JFBHFjLnojhFSTk
p1AJxGMXUlQf3/JJjM5dYd/mt3Y+YWJ4QgT/6lj8O5qKd8fxti+07TKsSiMiF60LAdpJaGbuJXNy
UypXFosrYy3gWDSvzXse70miziE6cCLH3p4lTkK4id1o3SkiibVQGzjHb0lITZd3L0Ed/hGOdgHu
20A5znwnhKUA5xFlFcFhJ2cg+A5s3NPx3ykF5Wh7bclxJh6LItAYeTfNzMo3QGifLaxc3UWhUhnc
UNEGRiaLdKWxYQTg6er0NphtXEr4TT1xCsjU1JQMWBslhVTayBaWwkvib5pUyaxCK3z1fbqalunN
4I+xSb7Vs7kguC5p5S2Q0jl8C2PzCP7tRkanIboBVMQI+bed4ndveuSiQfk65gvwdTbYIbTl3b4z
hN4yvyosyOghDtPk42wSazLCMWTewQT0Bwp0/ChAQOAdO3uCJValOS738l5Y7rWjX+Sm+QqQrVZc
zFD27OtPwB4GRVlYv1EJF5hFG5tWmaiEpihX1FMXDoDeE+oZ4gq1vG9CIWK49XM0Va+kQqjZ+WrS
qLiY1rBCINlAyYOGfX60zJMA8yui5kDVlUMfOocu6bUf1jMTd3s0MgF/RMi+tCDpDUhcjiILRBVw
9idq6yVfHnVE3OXS9viN3KZVIwa7Z4Wajk4cgu+ORZ21qIMifsMTOwHIgFnxzG7q08k12Np6iFDa
OzUe5mmhVUCddn1setuzoskVCwEZJCZITG3GZizOzihBGJBd1oD0Wh1yty2b9Z7Wt4/QqJ0q49L9
CTulMBsUXy+/CvoW55oBm4GktsLag/8BWe6vaWtX/tFauUbkuKvWljc3wy6nAMVEGljDdQ9eTpxA
SfiKYKHtfwqibWSlwfsTrb+sXfKQap0wC1doKmB3/BPbFdgIx1Otcc1ToEGe+l2UnSgrV062c3Df
aBx8vQWLPoCZlyhy22E8gvPkLmz8L64gYWxW2NloBc1jQqBW/xukGMoqjVA6pSa6afKzc2pEcMD2
mr4rlSZCrx+HNZA5aTe4YL8zSaaujGLk0QDvYfj1iEF1l8mKUuR2dpVOuR5PMfMPct9BB0npCoYR
uywVnvzJjTtTGxDDXVNrGeTzRWKCrLypdmPPxA1oDpU+kPoY5NlsjCHyFya0+vgRMamgtKdKMtCT
Kv2RaLM8uDFuqOjUr6wbLfJMViYpCuUD1yNzKXuDZ3Xq2dSpt1J0PrLd9QaJELzhOO/AcTpU9zJ6
xtsNqCltyAZXP/wIIzvrM3dpsa6SyoxInG9BbZXZKVthMNvqmAOXKpaNNuxHiESvfwx22Jb3cvLj
HurLL5AwVnJFbTrPmBrX3vk4dB1EJVihc29YWnyoFXbxreufA+kS3uhP9BUbJjkGC2/03GfM7TG+
67e79UlVLRlzzF5/6MzAsC4n0eCqJpMzEQQ6j7ou7znEagtUxJQRz2knuzxWfbZ8Jibw4J8Aoizq
0Z3TcGs8sqewEiBuGYP+H6v2EIyr9pzlehVARuV8/GLyveZIgU4dOrmiOG41lC2Qnk+5kZMw05TV
mt8nw+ZsfF5vry5s5bRd7ExvgjkjxSs8JpiYqhEa1urRWfJFX0l00jrXUG5pJbSVgIIaZw3Mg+RB
OOLSnO2xAWOMvOx39dz6jFXlaLzkYhuHMq0NB2rZbDP2g6HxwhfrFQGC0DgaZcjSlV5B96p6jlGG
Km/E58wGIEkQU1rEak327qyYx9CU2QZnWSFoO0WrfNtHkLXCvWMmZiPN0Q2746MHZ7JfhCxNYFTX
9vsWQmkK/L8Vzgf2p4UqD/FV/oNHsu9dbyTk8ciik6GU+OEv7xJu42w7LH2VskxDOT6nhPmEec3F
8PX0M7x5Gz+YT1gVvjpbel66P1+BGu98s+pd6NNEFwIZephCYnN5tiXO7NPMe0/bIEpSHUsrcAoI
jklApJ1jeLqiBRHBDqTiSA7lwh8KsDQGFSmF+81d6LSo32osyhhfP5aj84TnoHh1GmT5rZl1I/RL
hrgALJ90W/jT0E1hAIx3I2EbpvwIR7rWrIG4O7IP1vwnTRPc/3AQTnYmUCtIInQa2XRhpDVQeocF
PhEIyksgrAU5/09bTP0qkR53GLAx/pdl5MU94kK9rM506RuYTicGxlbJ7KgObjltWxbtOjO9KqTw
AhLbj7SnALiCjxITyGWVxbcuxFeJ77mVNexVodaqAF/rkTVqIEvmDxbunwkzta1+ictWAToK87wl
aK56McLCJryxEg3OOJ+1o9y3DeGYctMTtnYyDErIjdDHtW8Ye3GZctH1m7nVFVbCffoHXIJdbFQa
moEvjsw7zTHwsOGqKiJk35q2Unz3HudqDSJ5+gl0tTuD6TLkAU7Gmg7vEtHGkXFl3iJ0x8MIXvwh
JEdA7UqUEOppMsDBtbb72zNU+Vf1rJvLZj4Ktrn/pXgK9wOsrlofTuFiJN2n0kV3KaSu+IHcvGWn
ehAroB3zqz3nb+WCKlxZn1cEceDXgiqOwhivLwBLR+RDX89FPvOtezVVEUs+xz1LtyuQEvfN8Yzx
GewaAWRAb2FZzBoV1Je7JZVlEoZZ+Vf/pUh07TehDpWxkfCiFScmE0ixcYrGGGMZEJIYXoUPVaYn
YhRka0f6ujcICmnn68F05J7opEoh5rNBAFcxMqKncPqkPqFf/PKCJn7huZYdScWzJ0nVgbvroVMW
89xRbf6R5P2uIllvkRAfZHtebtJhmk9r8FmUFiFhs7UUAgt+LyWrkCKrI35uPCgl59V9QL5E70fg
ly3LYgycsndwIfWabFxETDFawIpWm1NgHEkQ5JyZLXnWXU3EqiTsLvOf/mVQEd8MysLJ0ajpGbTG
8bfiqtJCa8wpsTHsQjgBnt04n9fAKXkGRAbCJPNeyJ/zJcf0bN8V2VRL2y73JYrfC2z8DH0M1+pp
iUWdQDrtDcCwLrNjBex6WHZs+eX5TCIqwFWtmYrhkWeQaBp9zhvlabSrXn7U2qq+KpuM5iY5nH+h
kaTxVye6QqEzb1hQtiN/eULU5YF6bUUQj4/SYG0LMVGr3V3+ChewJGqe2ITQCRIYRzjpcaS+7hvM
8rgQ8BwiUaK8G3KZVerGlCd1aR5HSgbY1aWzX5Ip9cestr13ak3x8NNoX7yW/qrTKueO3Ud8EhJO
ccnfsH6NTin67VqNr2tGkYQSeC7MZ8ueV67z2SsUrbj9amHGHwAcakxePok7AxFnOPU18KrQlJEb
Y4o/k+ElbraaLzCWAhceeXL1nuEWjHks2igbJsbT8VFb1sxUFOepX2HtUXVH6CBveuDQjlhZQiiG
0HOyG06efcdmPahhASRSRd6xFihJfJRXauSGATEpNSAkkO36rFBMQsMErzF8Bs9iD6fsKlCX5LC0
LIMubVQ/8C3nTHqrM+c96Y9gDllCX/Yj1U4IWCsLBzNYEXOVLX4TI4yGU1E6h0sYV/3DPvVTyXG2
fWd3Thr0m/vqyKlPreZm0ep7hSMwM7DlgGt0FqTH5Xk7kjGCKw3a8K/IKW67JZ+4xUVR9xpyBgrL
yRCZ/UYerPiK51lX7yri7IQwWuVg8KWpcdXDk/KaJQLe64/7V00yZuhOKwjgtQbpcSqxCmkS2f6B
rHUziId0KNL2uly7b7ArwwZT84p+dJVOe4qPwqay0Nx213geZR8dLxwZfK7SLcNiWqEx2rIRap5o
7+SmRPZLaGptvqGDM726xr1HE9WZD/FNaMTQTiDNBugcrhBW+4/xu8wCFuBCWabhkzGBXAd7MarF
+z/3xeDWZKhm5NQjGTN07J8sjefk4/gARSrqUtRx7Hy81uXIrWs7hSBy6boqgQRiS4f2SBqXH8SS
u3B+cR9oKlkmt7SwnwP0/ifJ4NwbYXC9JC8u2sjqXi53eyanpM0JamHeGKzgXOizk59tCNvSONK3
TUz1xpxcbfGg+JPQvC8UWIny1yoFsyAdWlctOM3lzEmscvlC1ngmoxT8gUkSQriL7+nwJHb1T0O8
FpYESH3cWLNGn9YrhfPmkMK3YSXhhPg2iBMAqVRyPpHxcj8KIktX6uDH38eb8vLoVuWqcaH8IUa1
i6OYKXJbRrU5bq7q6um0RJELVl5AtHieGKcL4BmLqe4faI9HWsguJmdk9IuYHcXqQ7V/unE+p5M9
hDln67XMNHswfwKRthVWFdrSiWjWcinkJfICyyWQ4ZmfAmxDG67UbwQwS8YMIymWF/4C5yFpjSzH
L9B4kaKQnwvJG06CUxjVVttfSS4zk1sbae6PJSzAwxa6fQfKB/QZmDEjKKEURMbVJGl4i/IKY9ac
ZoVGQsL7uV4wj041/FsRYJ0EqQ+eph+wX/jiEpD+iUPmvUdO4ht4D5EtQ5vhBwOtIhHA9wuLjQbZ
pij+dEHysUkJC7revdBQKzH5zaH1R7ynLkvoGVMcAbjLoKR47yoO7cZ1fn75m1tMg3vfJb2bM9j1
FvND/FJUBVxezkwGRaGpO0+0yvcpYj+541h6QT322yF672Qc4UKfFuZpCxXMZbHlXziBya1eaxct
4xVVpvk0SHEpFxQ/s6AVRswm3LpQOSVTxG2cInm545LyHueCf2OLmA8AVPpdJnPntUfzPT2+g9/G
Ft27Hivb8JhkgrJ+Q9MNjq5cqF+JhuXhwex78sLLS9P2xO5qmlYebTNxYiboEAxxG8yKDn0Lhky+
pUf4U021NDoZC3brPH2OVqR0SHcvkEzrGO4ti+/UyE2d4GX/E6b3fHJcS5mZpEW2k+sTwPyHH42q
nHkAB1K6m3SCSRdU+AO6kJPqv90OEoZI3M7kXkRNGN8dJJbBn57Y4fU7GZ6uDaeJZ+yALJtG/tjw
q7S3pCPGl/0id+JApW96KMwYEgyOP2RZqKXnaJGjqr2ESb/dxLsV9IzHA5FVicw+WDfpBW6HE6Dp
O5KD9lHw9ehObR+8Oaj+2R/U2P2HGxwne9D6+avkMtpsLjcOW213VXEBUmFec3kjuPrFb9Wvy+Ih
SREXJWnGFM1X2vVb1CANWZh5bsysF3q+OhC0S744ACTlR/CKJTfHJWXQR5B9eTkn8uj7h38A5AEt
eBFkD3ZklTR5f0JP0Ya5BuUgl5JLyP5Or6/R8pmwlVyObv7mWgF1+uR38kLtaUtDknhpA6xNmrtE
CvJHwvFCgmP1EhgiRHXhpTfWTS2G4MYrq2+S5I+oFroYy8+2jorK8IHUdhPWcy2VNsfGVt/v3izH
EBPMruxnA42uCKBaZArzyhXTis6hs8yTLGiXUJF7NaOaFHiIE7+HexRn6/+WRTX6da9gOy4NITWI
pZkkAWTxmZPeWgXFlJHX+vrwlnlnZkxk8Q3wTEPEMKIeiugUCBQ7AgvY1TjW3wD83Tf6Y4FI7a7+
DWUeU4oXjyBiuixiLV+i9+gwWlKNzDkTV1AfKCzkYqvdg2TyZTW7mZtAqbCwdaX6yyzTNrbXIw3B
F/LKAzzKokeMqsBpzEnze1wI9L9JGlmM9YAtY1Qsmq/daCQkvvAxwV+n4+y/JOJyJayTS7lqczxb
V+EV37DbrGZc1dd3hdchRUGdIrcREyUhIfeqsV1kQxZ3pvLe5Ci4okYb67HYmz/J11rdBagtExa7
qHfGD78S0PNVScGC3PWe1MzdIOXRxFPOpEcpLqOnsGIz4HGwhdG9BPM6X0iDump5HNjHIoWuMXri
a8Tp1sil9cftiZl6RiJu9fL2g08GidD3kQNUSSyIPksH/1yWdaEsfal381Ek2qIikw7SPFoqMSvw
e7m8Kd0/BLVTs+4y/tYLOKK160SmiokMl/t3zlzRcsSns/4mseRFFTvwK2RL2FWfp6HU4m+NP5vO
KgG/pjgvEiLnRirWUuqSDGKxk82M7w3D2VrybP1lW3Q9MNvKTwKvIJA0HmTdq87IrmD7Qox2wixD
Wpco5Hq1eFy/2mHjqc4TGuwTHe73+9UFEF+p6vkq/ybSPaGpRDZhS8K8fBxdIVPwcyhoHGq1uJxy
T0yEDQjmR+PBVgpJ5obE8kVoSQnUlV/xOwth70oBlpaFj9zquMqlLNXeZlJdlK2/ZMdTL7KUS4Tg
c3Bit898wB0LCI1MgSbBBp7E7x1DoJ6MWhcb3JfNIo+P3klTbDT6gkLF91TsZT767PB9CpY8WoHd
SERdtB3RLe8ljU2lw5lRaMjDofR/86rIpl6B0Aps1BwnNTYLsAeUEIBhbvzjDlYnr2Jt3317zA3F
c73Cih3KEbFMrCcKzhahI6LLTNQF6IDCx7B5kXCTVHF/sAUgujN8m4MI9dCokShRpGl0x0z0W+VG
CsKDoLqyPC14CMe2HxtCHQL5xWg3hntz/oCc49MebB5NLg97dlaOoDg8g8mOihUoj6wQgRdAkTBq
MaNQ7VIO9KbJGZY8ZBYuzgA/uWAGJMbEUWheuKE9k6BBpM9fxF2deT33ARAJmwngiBYy6BPGz9i0
fWTLncxD4U5sEBu2dYonUuqOgHBsG81ISIOULtysLRKKT8/pOUYXb78ssIojARrscBrpCRPcj+oN
EW3Yr3kdeZ9j3m2vWJH7MK8buNMnw5q3TjGt4pLsU0Te7IFiaVlSNFStItoiyIYLENvjpPwkTVsb
QnyTyfrj2xdVStUWhnci/kawTnLabQfw9Id3DU1y9ThAPV9hxETSPzGVa6vlTMKu20bQC/gTPaMF
vaECFagDEXiKLrlSOsRrJiWBTgwPBjnU5la1Agm/HWmzkwfupyCELuS3orfNZhC7Rd34+PZ+lBei
YUUGZdLg0GXMnPJAIym1n2oFz1PlWVgPwTFbd5589xlFj2qDTm72zu7j0do6UpFYuAjnyHeyhALS
m2wCdAPdy9rIBJXVjuPxASkNomR8BMMIZPuTIju/SuPmvQR+YdLuDvAQbY1Je8jFX02/HMLLi73f
7kXRoG8P53MkYaWpgldhVrQvULNxHALuqB6cscMTOWe1T/2epGx8ujsWAyMWMb/ERp2yTnRoQ1TH
750iWe0b0OaeCn/yqQEozx67eaw9ZAM+zj0tr3a2IsmYxVV8fG7g1x8pj3IUtcE11OSDDfz1Tiwo
t1Wxl5bweKcDmVDoNfciajWmv/40isCAy8gduCVwhJ+VDbuonW7Szv4+9CeRX/hW0z/FxsxQkyPM
/ve7EeDQTh1qiBjBBrG1vBbr5sipK/q2ZQc69FPC/h8Z/WBPbEDrQVuJSLYnSPhvkwcD09Mvlu3k
ASwlnNVQkABYiWG6l0gkeEIij14jfYztEKKwEPUpAR1EUWImp8ceb7OAiv+Y0RT52888M3STfTIC
wJWAawoznT6AZYrH3tH7FHHGOBUp4+8pQ2GjM7sS6HDeptytZYKms4M81GUSikzVBstkIYtFeaLs
SXd0dVvJpj+dgbtnV5PGZrZ8ZZPymGWz962s2a+RVJ8Ze/6RRVrRLkidS7zy5hWDnWUHKe1Tmbj7
5I7ftcZ2dLz1wrVY/Ydx1fYD5M+Q0NEmTBY3peCDrkp5MlCN8sIgm34jK3fU9h/Ok/B8ZOJOj5c0
rNte2t16nm7Dgjc0El1Jh5XJEzdpwKV5n4JLgcz06MdZ47PWCUSW0YqNHXo3/ouqSk1fr4M1Vzal
bPJgcRrZgboaGGAfvjdo/f/M/MjG1LT/VPhHHhVFAp3yRHPITbZoeXeS3hZOm9WRyBLWPJkxWxZA
C0CAo9Umv4reTSQGWTW27hseo5wiQ9RXcLDRgLz4+LQosv8JKVcBs2V7pY1FAS1hN/VJ/nWXs/E9
WEJ2C4AYKVen/QSnAAWNoCSR3w3iBVvEfjxKrJyywtgE35iqyw03UDiZEHyK+uVyd1n7vg0EhRBB
BizOuBL9TWXtfMa1d51VzLqoXS34nmqV/y+l3OArjYYcv3j5W1Qd0vsFPAVMd5feSZ9MFlQ2z2Yz
eww62PTpkMZRy0YOe32aj+eOq03kbsqqHgXcI+CPx3co3r4FivlpibofQSxfLOq2nbbtu6uHM2y9
IDB38ahT8hCQJK/mLpkL9trvgm7mp9g8C/WLMhodVGrEAsnoeFrwCG0Nb+3VbacrEeMWxN3p0Uk7
Dir7hWw23Y1tMPqQ5xp+rQmEdTRkf13kdEY7D0LNEpP4UlJp9hsUTk3iSSMWNAzA6JzkUZw1l/rC
6/eWNM43XXK3Ao/uSSvvVLQGGqC/uP56wm9FbRS5yCAGC7jFYTK/pHdFmnRrJFI9PgOE/c3MRATm
aaGhozUs6Jzk2HfQxttaeFX6hUq1u7tVzu1l1KOT1uZ2veHMm4EXDaSFMw1FWhU2tUuw+U+vQLa9
gVpCpqwDiT44MgGPkSTle323vsnH3ZhYHgXNAZGHvly7ODA+fbRKsI1Y36mluOCRqJ3b0Ef2EA1H
/ZDqWxV71hJ0zZ3cYml/wCfa+JnqxJqtfWChkps+2R5Z1dJgbJoanOzdxh10xqQJ+nRvuV4VSJvH
2PnFeeiXWE9yFyBqzi46aARtu+qNMqTpznbCYQNe0Pb449Xn8xFh7UG1IA0n35r6p0GAlF5y+L4r
4Nqe1TpPLiC4W48ZhArqXF8BtxDnXDx/r86NT+7Mn4uHPNxSH/p316RmamdqhvHL3YU4nwT97ZrC
vxbrkAk3Vz3kX+rpvT0t+zooS/D2mjUkkUN17znEMz47rZOG5kcn2/7UdAcTNNMo+vHxiGw7EGGP
0IFdtKsgxhtCSkWXJhKESqv/5vZRvh8LyijYfW5Kz2DjcnectQL91Ha5XAcROMKd7mw2t3Qxyrd8
6mjP/Hi+IEF7O8y69rmzVt6eq5/HBv8EHu1G0PyezUrcqUXK3cqezvqeSRsa6MhmPNfb1XUpS3eM
zbndRGiCIykgJtQXQv/2Jr4QfClURyzCvIHNgpqpjdkDbPfU+i1gBKwKs4uxi224MioBgM9ja47q
XLnf+pm3biSnH9HPi7We+IJYpq+M+3rPIkUsCZbEIW7UVZL/xSuFZEm45R0r16cY+obfd+rqRENR
ibQhfldwHUhXrhhHGbYMYNfTfcieWlnvMcSf63SGEGskud+S1zydrBJpSWayRLNE0rvcMqKfbAGg
WTd2FqwF6ffrp1CzRqRFZ9vlPIzsohsXM3z1POot5EqLDj3GE1UGSmHCMzhUmQ2QS+oIbFDAQT0n
LaQ03sHAW5MUBTlciDuz9348EEQLs0L6ejtWZiXDSBzEw6uTMgfk7jEpqTobIlaRxg3DuOUSKSOr
CleRNWOFdsG7+S24uWV3DfWZrPkhvcweLR+FmPx/NzTVK4igaDqxU0e1KVdX3LuCYtW0NRh6NrvB
fks7zeeU9/vwnhNJuTfuKQ9fNz00qTaXC0iYbglDKc9fYeMGX5AKXNPnnfWoFvavqjJ4lIUfAYV/
iOI1EQOIGZOBGidSZ5I7eQQGhB/XxWkn5Pi/a2E3ktmdePk91xax3rXDm1oxFuvm8mOujqK0EdJh
VdfCn4UrxGVQ7UrLq0Ijd2SJJ4nafGoChbfmKw06b51A4cZuNAOPBrCYGqunWtIMlkSJirFxeIAx
+vRQb/Fsu8hTNRZDRyA/p1blgk4dOPygvIrY8XsOHrV5UZOj+bOgaKjeqm79LAnL714arTE8q6pY
eNsgLJ+QfR/vXhrhIlV4z2Uq8XVqRAV8daAAqCNUmlBePh4wQ9sHJhCeQanWHT3DVeBlECBIxskY
nF93jzjhEQmclfk6DjIlPFth0AiVD1MCnB7wTxSeGPBIYS44tTHZ9YloqBgUuvd+ovaAj9DBnCOd
P5FzT2xvRK3t3ClzKLJLu6uiPbPtkIETYoxNWbW1RM2j+EOQpjD9QdQuTmbiON6tTC5KvJs4D8WH
1tur/3LTzOxP6uDID9MtMp+y18928+wUDojHyf4vGJKFnXvKpUu7chDefS6t6QvFWbm9WIlXQnEq
oaht9tcUR+3RxuTnGKuKhQ7Zkc06gIQ8zZsu5xLiG86gOe+ZobtsArPu0A/4pAJ1yGsc2Wf5Gxq7
9AIkAWmOvzX4I5JdBL65Hqjyfk/vJevj/8v728z0oVjPtlGHIAE8Wskziq1Q5OVklM4CY+F8FEHN
90pYP0T+6L0soJPWlrbcGCB6/Xn6AgPtmLW/NRI/mw9JM4QnqD9tRE0x9vXgsgtv0IS4GFtA8128
Z8FnyNIyWEAGWwt0YMVV812uZGpNbwZFUad3/MGqNFXy/oLObzbLa6t9I/C8/r7FilkzlAcTGCz7
/TbKQheOIN3Q7e4C3Cp4MXIY/trdoGqwJq67OWxWpaVcZjS80aKZKi1rIK6cizePx/ZG9ijZLx+Z
XiCdYIB65fOJ4SuzZPqt4dHqttdNoiKz3eX3z93vDiUS4raPenpmYCHgfzgNjyi/G28A0GnwGVnW
zPyqQ3ywz1EF/TB38HchGqrHfK4WXoN5+NYpSAXiIwGLFRGWyuH7TNK+iP9wIxMnySSbHeWp8vCU
SIHMKLR8XQ4nE3bKJHWS6jPk7S2GIZPGckbuFb+5uxkQGC7cE5deta4B1O5TwuokB58trFsUfjdc
C9zRwZWS+Ak9BRILVnp/OodqdjHJ4WhEjyCwtXzbrvsZR7vxRWAj9s0BWbg3FY5RaFHZYDjA/1qC
/rnfCPZWYt3tMhUEL73CoCwSEut2pI7Weez9Hb5zVYR4/6JaDOEqzJqdvj41IaPs3LsoyStNrbY+
7eMjoSqz70ih8zepENgbHcWP3ldfco16T3g66xSazgicNYZXIA6erRFgcX9Io9mEKo6B+oxIGupq
72Kl2efd0UfTv5YBPwZjKAQZTO78joXpHXQ6w0DLo8BJuUv8kdc22o7JVuF9HxZFNn9qsStQCfnZ
V465EbO/S/C60goPGPXwH6U7o20yxN0FQbbSxy057lChZmsF2VhLimX66B7KZQtRwemYOOTa3vgc
x7iPLn4xS+kMPP3hoA2TP7kB9uNoANjKcONX7HbtH5MWPQ1pFAQ3i3pql2PoFyZ/TVozhsWg2jgT
0SUNfqvzhx+AVGBELz8kK0FVKiAfSs5/TkJxUxCeM2n/DgVEewtrNlhvZPcgfG6Pug3KFWYizlU2
nfUsEc7h/UrOWO70RFxsx1H9VRcwghwJr7p0lH+EIO7e2lMwo3jcy3wMpuBKc/5vtiwvfAhyymE1
PaKV7fx2f8DDaORQ8B1lYnvbNW+56NOEY2s0Q64BmEFHJwMGMkZp/IZg3Y5Sizc9X2Liw4es7oOG
ciM0zUC29aJDqo3XnL1F5A8KDSwzfp4jyM6kA2R2Icv3S52OOaO+cWomoiy0HJCYwS+5TEUOpKf9
9o/dE8p+HFW2Jx0UHjjnn0LDHOi+Uw857fiTviw/rCT3VgcK/RtrVY+R0RzPNGjKMLQVRr8tOuS7
Omm5tqq/He2xfrb/RD9BzFP/CdDm5KNfpneNVtRdSf1T/JSVSfQifvWXLpCauP6W450kXnzMLu4X
2VK4xriwdqX7UE4tBf1TWHLFAb6LbSW+piENpyg9QqV3MZ6WZQe/hksJIGqguFQpvq7bxhj3uzAW
ory3H2JkUXXIjWPE5uRMnHEZ9HfOpZU79Iw8OvYqkju9TRx5L2UjP5ybetWBk8YHLUYo8sAoc8LP
PjORCOlK2JNzJ+fanNEHSzkcTw/+NuRtshIj3RoPDC7Grfe2lJ1LhWe8O9PGMO5nUYdcy4tAi0q4
F2c54zn1tLiiCxbl9QVrvyaAhazPqN6No1/rzIRi5meeXFqoL+vLcmZSh/JwylxHqXz9ufAERRb9
zERdmtde7vVS+kh68lnvsjY891sW6dUxjUUuAubyO49Fr+5iYnB2QGyI3D6d52Lwk7jW/B4VblaE
g7apsAbgvWJgNoWW/RuJac3BUJlK3cQ5H/6uugxF/hUxz4Olzd6S4RR70wznhUkUAasF34MY1jyZ
TcoRuFfGIzmKfx4MjlFs0HXvvS2hVaTk/E3MwrKKXPw3e4TSnJGUuKANZEubf3va6x9O6CqykUsS
SBtAM1xmj/ULpPRrmLcVQ+f6mPsylzb7IOp4E73J7+/lis/WAgR8Y6kx9A2dtSet1L9r1JaGvFoM
aeeyW6iM4fvGcStV8/5IcdhRoaw/crMgeqtpYrg6WuwzSH13XlnYpO1I13Zeh0q+cf8wBVoBcEAw
FW8uJq1guCqVGwDMhOpFI17p75FHlhv+ZTA1FLl0kR4M+Ixc7cFA/urSRj+pj/mfLLRzfVy1h47S
0i6y3lhfHN7vJ0bn0vkdQuGKzDjedMA9vcN2Y6+QpcovFZ1i4rXSiyN7et11lJG2mWTun/FltI93
Xbpn9PVA+UtqhlogridUmgElKvIc/Dj3hwrT0MIqCtDztXPfOocp9bvE2Pc4TMom8+df5ur/dbPy
Iikr5+PLQlSquExVclMo0o8RLZCLbMyQn/qDa2Xkfl7LNW42oj3sjkFTiwOnNZbhjhcJFsYEGTad
0e4Zn2ALnuxpJjJhcTjMmCMnMKxSR2jb+NGWQAXwwrXkZfjvcVYzHGfnUKWf4Kaja+mV1fdTUoZZ
V45cG8tLlaYSKnCP03aOzZTsnJbgnjZKdMwTYbxxdaBd1ONFADAlzpkUJ1ZTrr6R4R/Rg9STaDQ4
bjBCSXh+49FHl+Lyn4UykGbx9fWQ7EpbxXbtfHyfVLTUe3OOfvUOUjvFW3CBX86Psn0CbpOoTyh0
Jh7T80hkca/s1I9eb3cQ3XdMxZ214yihu7COoZVxgj4z1rMK3tq3VDCRKzvv/KLlfenQsZF0dX5e
aR8bi2cR/FYZAQ12zD/hI+4MIUh3U2rvZKmsDG4j5c7LizBH/UOhzfrJisL+Rn8Y7D9KxeQrDzo3
hCDnUhmTA4OUXJZk+t88kYLWNq3CrW0dY27QrvX7+ouTwK86y+AUOjIxX70zr8YqTD6FKRrvpgQy
Z4jlf85VK3+6sNhw84O3aM/uZ7Tlvr6UdbkaF9f7t4B6ga3MAN9OZ2MezhdgZzlt5FDVQGAjOmz5
npOglSVApFZZHOq6bxIXbGlFUCz/qj/W76xhFfle7zS2w4OZCLju/3g4R7Bo8f7XokIvOmX8WON1
9stR0p+eb8IDuzkPoK8BgKmrV7UV/ihg1RhuYA1iwzTWTQK/skQM6HLYsvsCuxiVv4jFAMqpeKQx
Ab642C9UlG+x8aXII7SJ2dKawTRPKXajrtRinPZ6q3QS+ZaLL/vrny8J3uaaGD/mv2u607/kJi2n
ZfCTQ59DDc176lb8K613tQ9UgN8VVJMhpsMVCU0zo9Kxx1xp9Q1uTCCwrAHAW79QfbLBKAcop34R
XNolGXUqTPyY+1EdYFmNSdltxBkOd+/I2FkE0jll/OllXdcz5ETMY6W8v8irLM+UuReEzn+8xByc
Pw3tzTxAlitDXuR/jMwclZr806+FAK4eYFdFU2tXZCQkZS75hZtEQUFJBE/TCcpOKnlrBWdWsckM
f2swDnJGY+MznQpUlO6y1H1aM7h+rGgl3mbamc5NDPOQYud10yVk3THQDRkQ1n6xRnmmhEN0fwzS
NnbAM0jC4sy/Tux5C/ab1GyNLkcQLC/H64tKRHJL0FIJ1ERyZa6RofyIugyw02qPC5cCct8+LnHG
JHEt4vGXDYq18p5PBsIT0A0AwkAFlOXnhqddhECrG9yRVX4yy5NBwJotC73i5hWrkjCdkdaQlGlr
YHrY2v2+y15J46vyb6nZHFnfjOo1dHV3Z/THeIaxaIHuo4P4+TttMOC4uE+qlC7voUqU75XTkQJA
U7Tvmp80l8g7HMHatQb6HykMwr3yGzbBhYBLCGCWKYytRsPyvJh4dfdpgbGudj8seERfmuKKHhw1
DEkmTdrGV9AHgGo5pXUMXFFFZMnKP3dBlsfbksGcpIlz7uSdB9iQZZQzAWTzItY5rzF6GJ05or/K
BhTN49Mri1zuABK7iRUMiDxgYPswTdwqinBzyshNNgMpFEtN+GbpqMFlzqwp3NKGU/J+eokT3oYR
FYR1yLEk9c2/OOYrBtjhEfcW6cALVZYmCVNjz8REN1tUJg53IIXfsunhixHiq57hz3PItCIDNUxY
xemWU1w+IhkhEce305ogNBMaXMhbZ8joyhsOcKjZCjpsHFqZk/Ah4upfZh0lglZ/92GrUd2j7ubQ
7Q24pVnKnJkR2d4igiv6ksOI/JsWTAz/tE4ZmiXPal5Ibgxku3jcEjXE3FaHpyt+zdh2+jytrIwG
R4AZJo0Qc5dM4RDNITi3TkbJd5rtlK2znKSwvUlBI78S+VY4lDh/2cY2T1VkTz1K8Stx6N0qOiOE
e7Esa1Uxab+96hwcDGU7diL1ggJyiyhVaKMJHJ4IyAalU1i0zVSZVmKj05iccWuVUJz39096jihM
5zmGRnVaBZ9p63UBAU6SqwvWC8niQFX3+PSdcvx+vjtXLLBq68wPLKt1clA+Gh/VvmtOXy+FPmn5
HtIizhRN6nAiB+R3OQ1uQvxJsLSInS3mNy11KoMRAfTVWGzC2Aho2v4DmLgbiePjFJWye2xA9V1/
tyKR6pbettMA34+sHp8TZK4x1qb5wYc046mWP6w3fVmknyh9jrHISkPKOgwoJAhQ8crQLZIQhGW3
Hp9Bij3M38CNLtD7oRs1E+k5cVgagkTyWSk5EKPaDJS8JV2cR87YzFgV3H6TB4lCrAE20evpk4B5
8H6qyOwTv8ipwQKH34wDaYdwv2gFXmevG1m1hDCl+oTb32apjGsLFwS1fvgqHtebXiBXOlM39N8R
M2rPtDzhzOAFsb7/Egnju2hvgErXTcs+9JzYPlJarUF1llA+1692Mht1gJgdHff0aWEe/5W5VE0C
q1jLfG2zguv9ut846owgHSXr4Kp2CbP1yjUeEXA8BjkK4hHDF9GMWp8eDnUWXGOoljsXCMxtxH76
eZNEUkhBzdTZqfUVGWG9V3ZGFMgbOOIPeMup3WYUHW2iYvfHsWfaalRydzlAzcYw6y03/QEsOg8I
mAMYlpUvLrnPtxfAyfConxzkWL2e2LsTsFi1rtD/UBop3BaLwgmgx2gBybnVJM4ID/tyrcsisMUZ
RqIzUMV4anlPonEyC87E4nXfMofrm22J46tbJ0xPo/TS2/5cGQVcTmZ5dUwXeb6Pw5ZmZdoCBjMv
SeQN8mb1ETcnbx84R5hByvhQsQAWf4ZnSH9lmACnjyf672NkVuOV7FEYlaZs9p8KnzcCmeQF/FYx
3tFJIwcgQikDGm3Bro4XR4+8H+InJMPJpBfpQsd5qrqTEwLfAkIcJXCp5qNhZYPtLUsP846MGOtV
2igt4BBsoK78NrIXg42al185caXOQVafZGTNjPz+LBjWpL1AzKA2vidl3zw/fLxAciwi1WPo4SFl
+/5hZedwhGLcT8LTjBkhf6hi99//7cereDXxGsb7j/Wd6n9vvCRf2utlchXzk0SROrRWjKGoRn45
B88H7kVQdi/amZyj0jC5SGfwtVad5eLEAfOsMZt/3ZEic7ZpurvbO6onYwsKan5PoLi8n1jAjlAN
lJ2ibe2wNKLo1ecCMuCjLEofMTFTA9OUtGosvSQmbZWE4C5KW50VpqtVyGpNlZqUql6CPkWuM3yJ
bMkHi+74vn2akH+Ki23ZeP8SGT2AmBJK+prupp3dzEIvta4Yhp5uOJCKvUfAOi5oQ0AEf+8VkMDB
5PMsuTHP6IS4IYOjOQrcGW4YNFcH6wHLjCrBDhakijJJLelcou0vi2gKfOz6/x7u1g6SwPF3gPv3
EONNUQhMgvo+SXS0UYrtDMnaB4JPsxLY79XS/Cae8wyxS7S4xi86du5xB6oUFEg+HNPC6/0mwA3E
j8D364tUboPerNONz9rZXltc0xeSWImEiEAS0qcX1T+0Z9vqOJA3LtpRWMyax8DENvB5L2WpSQnH
bjo5Ovm/4FgDNltzWLfAqdCjfHO7cdeDGzvC9AYCe7tRuj6Ra7ES5AvuVsazqltVcHWau6b+o1bP
urhC/GvYN/8pl1WsdqH/u80SpiJekrUomln9hBg0HPVGR30O7KOodrpzpTJuVvHX5XdmZSlfgyfX
5CeaqnGczkGXpiNF4K07ku+tCTn68nWLV0ysQqgiB3rcxt076+TErFvOp4C0gOlLlYuEOzlyMMF4
RHXixRYgrBIO0CxdzjNqrhMVBkphFuKiXnvNPTMIcWBtoZZV7Q7b3X8itXMokG4SwmbgSCLa7V1Z
heqxH755+WJBIax8N8pDOC4m0RYt+3GWyl45rR4juEFzKl3gmU0x+qZyJAUa6eYOP9eQw9ktQklO
x1xtj4Xqx9zjDy7IKy7ejM8/OTfWPHMXAdS9zJu+BdthyUYPccIspv7GNZfui9wsmoaKv4PnYBq8
aygj7ZHCM/CxD1aG0p6PshH0x0Ih55aJLuD5O1BgskkchlES6YntNySmFfJiFA1k55JLApE7cUvH
ZP+/Gw7xP6OYpOp/abXiAv0ZYX/WiWjCy0XWmfENijZmhJNHhnjgtfjg5TUGN11gPtYTkLWJ2lTa
ASV8a5QyKozMwGvAJxY4ew9bhphEh1CM9lIa+XcbAkDGF8kBCoyVYXOf1P6nlPOlsWaIGgpcnzh7
3OZv7tetgSL8JtG5csNo3ufBgbtNBZk9wGl2JOFm1slSWG10ZmCe3BHoLXx1Vmh7qmhMoNRevEl/
IehMrc9daUryf7dfkI63Dfx1uIHRCTMDBW1jB8GIOXoQ4ogrLY2a3sFx7q3WGLGMRWRBjmjVGzTj
K5ptKVK7TJbSV06dWytP+WS0835/BqaMWGs68bkQYDBP+xTx4QDnUWzEDq7QvyqB7sOUbP5p9ZMi
dqndt0DB9qdSBDqU+VOo5YzvNswBFXGlPOSe/k3+fgrTUw9+octhbwseiXRXaeUasS8fC3cHX62h
5Jy7uNty7oK5gkYJL1ekUnuEW6U/v6isEmejzEsSpQXUllwkcAFJLqcaR/nmb3HL/prl5s8sybjR
GfYtQhHeOQlrw7KOQNmPGE0F2Zeeeix/2VGwPpg3cp+94xCRUE0wVs7T/jShSxwPNQTlNsULoWeA
GyaykCDedVTqf9a7pAJRZ+OqrFMbWRGJyVLTzWWaWdO3v5JKE67vOYI8Il7WGGS0nxUyqGWDflKl
jEBQUDtR4FREVGvqQNJMUuueuvHZF1eFlkVRiyrfZ7IJiNqbNdy+T70N29V4oFwoI8weuBcmitdj
fzFJFqa54JoQh+scmc/GurHsFsQpkmIDEMH1/ZrgO1NgjGFDguWesHmdb1mCyJ78esKzD9m2uxEr
0oDOE3EKFd5As+uGqJZzsfAb4bUX8iCLrNnCOWmur779GFAZDp2HE3L1ihudzUFwq7nTyLqdIGRF
rciwXiz4IObvyTbMY2NLkX51VKYf9aQPV4jTD6SshW3g/tUFeIwbaugUpMf0F+7iUrOcO/fhowmf
065GbmM8ce1/ZrBwa3xi36MvRW4Rrd23Crf0KiL1sm4lhyDaPgTV1XJ//5p7nQ3AqI9/X/TKIRTo
0fZEWkykN+2rf5S3JRomRBSv5l9+KJB2oqXzog1nfqLCeEycWTj460a1vB4fHpd9K/1hT7U0fFbk
Rqj22WqBw92G3mr2T53+2xqfo9fFs2zcK+uosh8rlGR1LYIzK8xOuQFexPAj0zHWjGL+URPlEC5e
qp+87VUJ9zcgiT9BVDf/gFGWi52LAJBCAU1h6IW5TI+qun06zd+s1pwIKADDG8EkXD4RYzCVqG9z
rgxPKiECE54J0gDl6qdqjNnZUaov+DMLKKwXq4MOpkDZn0A6aX65koCksAqZakNc4S/5Lhy7mLx8
L3z1i6BKJYSVlPEneKMMYgJZwEbU+tmnOTWFwZtqanNXuq5nZTYLv9KjyuLpDuR7ahyDCMpcxmHk
FhH55TAezTjJV8NwWcwiLyn3nDlliHpGaJ3YMowsGOOWv4ZUGvpwsaD3fgKfxWi4O3oUiREiH9ZB
PJAkDQCfExhGj1LMJp2+W9aB/Ws67tUlkprCGzX+q/R2Ng7Zmnq3tC0kO253AiTFC7AwrJAdWnJe
1ySIPjynFqTM2ce02YPKKySCYR1WcADpaqlbr/p4oa+4bRLbqn2yCYFl8LtQS/RG08QaT+REbLea
XqlE5ihnvHBHT11YbNe1k8q2ESniTdPi5DVuOFbAi3XS9z45EaQ8ZgBF3nEu9V/TvPhXxOzIsFG7
X697/7X2jQD1Ja/E1mn0ZwfriZM7yCgE7yNhwrgjRv6CyOwRt92uyKAFQBwPWX5BrDiNbBglXBhG
WtnRIwUo2qCoCpdmPW9plku1cXexmmsMI4i+GhcWUKJwN48EDoDHXj5Vkq7LetPetA4uSDBBUg94
3Qv97VMfOqOHcTGRRSzabU+2GGEpcotiQPY4ACxZ5pVBhg7hEO60e1ExRg6YMX5kuShU77nmyYHV
PNMJct1LsJ9r3DM3jh8X8fNiiH5KOFpUoFq8tgEVw7twuam21w3tpogrEojVg9hH52LMSzlTa96b
YZ4GTfP/Pgag7pShlC2GEIj++v8nAt97nmBES+vnoSL8v44g/e7IP79sAdsTOk4vR/gZlSnH/IRR
A0i+3pWzia0ltIKI+WGFurFerA9Du8r6JOmTykkFSN0b/hMh6zJ7ZY7TiDpZbvR4+ZpWwAfle/HF
zayBRc5tuCKBYdu18IEgSxBWz9rcfnsZ9VOAbek7R7Wu1B3VNnDWYXNvMRmwxjwmJvkrJ4qoUKkk
h1xyQBfSpfZw0JNF4FXd21DCCdOLIGgjk+GkmIP53pqV1zcxzLovXtIpZ2Dpsx24DD0AhUVNY2BO
u44OSwhPEoNGOSK64AXHROz1vidrVffNlx4cjOEx1/gHeRtZtWFXiJ3SuOOm+bUt5mOru96i3+hd
2iuSP+kRc1dRNFW7bz4AqC34MlIasYZztqcNg6DP0QOCVDmVlb9l8w1+yBGPArlWlpjMQlaVzlcB
Rz4oZ0uK705QABuarozZbwVDANNuWD6n2rw2nN4R5GCN1VJZ2aiRM8hYsbTyjHyKqQFYnN0gS/4A
/Z7+rneD1U57OuxfyXFsD2dXyWjsMAoMNTYaZKnvr/8175w8x/GFOftxnHI8u0aAZFBgciOMLhsS
Fdi75u8HGmvHJCvyY84IGDzzP5uYQiEZFYh0BsuneVpORKD4kC6yHC+jal8HqNESTm4Pnaac20Q1
asM+NmMtWik5I7vtcu54HUiALfyDsdPQsNmwJc60Ao9MepferyEGwSF3qWenjMQzgIGf7/nia062
lTRjuJuIIdsrLSuMWHwk+VKGUvE1UCV+uDlfb8yOyFWbn8xQiRUnV8c397CTAzFZ/2wmM56xxcu2
DU/SUSO8YoPYG5aaqf+8VLv0UENlM1VYN2crSv7BGRKBrPwwLytpRWwmOTA198ndmFM+HMclkhof
AVqIxpVs05i3qDAmW4QcAnL3xA7dC3lGYw/qswxKMl2oyDi3nMLPzmT53Szra/D5pBcxxm+V98iH
oipoqFEQGctXhhaNE2ogUiB6XpR6qNzModSpwrGSmocbopMzRMPeXgm5ao7HBK2k4Z9pdEfrzw7b
kRTnjg+oqBOR4Er5ek8uYQKMArk5d6Su7/zgzdW4PqjtFkc1WYId8PUIUIxxrZJiMMPI4kMo3ldO
KcwSpkYvVlNypX7UzC5nQ4lh2C8RIDXsdV6bXoGOzbqwYIUzhLbXH/s5OE7ZIbQPIN4snteaVuQv
pWTBMoPA85TzMtf4XHm33pQoDztOPLaAOGRXZGMHtoiEfbsAGugueVq3q4w8kjOpw/NAUosmWK/c
njS4eGXoNy/FYq8suYOOU8CXlM6YpBbNriZgZ4XZZIyynaURVQNMDPf/Rv6+LkUz8jmugq+aA+Ha
eOhCzh+GEUKTp05oUFQZbJUVk62sgCANn7dpBOK5eNYg1fbk8taP4UtsuUs4iVdhCofwAZfPoqgG
co1H0aEzfobS7qz22bn3WgzpMTk1lAGzOY2UPxAwrzaJgOTw9XMIwe1hinMg1GwxMPWHpB0CyJQp
F9KSC6YJz2Kj+pNEUxTEHgSm9ZPaSA30XNHdDdRlUYSStTVizJDanah9dvDDlY36fX4te5QJUZmU
9KkHhVPHM97fFz2PX6H1h4FmdFPecEPRNouPRFW2FWa+WwY9OAE8lTfSQ6whrZOJuxLBtkNXYKHe
sPzxFE/PWcHnbQRMRtVYqQi11uKBO6tOgNeZVFq/XLKmM5pMsOuHCO+dCIdxSWzZGYKKSsTyLp93
IUMAi9FTEh9bsvy8DNifzMf4RQasnGDG1mvjx1xQyP3rk7fOt/pvGDBIcUJHw+/irJ47ysm6DgbJ
4tIP3U11sYpqoXSNLSumHUfh9UkUfZ2wHue4ZZiyzoWHTauRFELpr0v2dDZFbFgH7Oy/Nb8GZQgv
c7hVTqdJI8AW8ANd2oRsMswOB8/LzG33vP9oqil5zHtUFFRowtzrG/Fz5QwVUo1rdRRqK6VnWf71
xbf8X1Bvc5xhp4+fS6ati1QaYUVd88P6kslE6LergycV1YccdPPYB64Akz+PlwXBD//Qysj48lTz
s3nya3BKnvVCJD78ZJfPhFbEM0vkR3tm6r3/V0SHcQtoa8IW0t7UnutnCjAsd44lBbEU6lGNVwvv
TDmtO/SqpC3AujyWRUQBReLHDNZUBsCqVPgEaYTAcYY24JHU6ZwxWNNdnOA+oJK23HPTh2MDlHt/
duD3GvvGnPRWDnE9EnoepS4Z87T9rSbAz9MjbUg9PJrGl/iSedld/gri5s24tlPcHCO5ROOQJj6m
uexXLB4fkHDq20qUeO85eUT0evf67+DYikbPYxstueTp0fsxDxL0iB3w/qo/0lDnbbFe/OBaljNV
0wAL16zN+pfUzEBha97BR4bTaHYiTYZTg6FnRregCELljYi8IZZpU7vvPP/e7d0PEJzah0aVtxTe
Ha8dbt0AbIQmPugzEqmREZRDn44/zzWfoz/ea5aoZ7G8wDQZ/TcMLkXcZQYsYw8CeBInAU74T5zW
+STm7kbW3aDyUYZMyw3yY4+TXWWM0nrZ5UB8ZSfu43Zu/24T6D27DqwhdZ8tES5Z78aGZXJ+uSOC
l6Ap387hRmyGWogsbaC2wbcv887UDMMGHkcaELqxCZqXlUV7N4q35DiTa43ZegVeoE0nH5+n5UvY
3tcmaNfQdeUkDMVlXC6wl4OpdshU2gIZexxNT7BPJrD4+Bu8hGs2NQsMwrv6FYsZjduKO+Wt2WC2
u8Pt0u8asj31ynKbTEZvJQil8GCou+gDUFfxUSMO8fzYGwXGJzhBPM5tEa2Yg18+4MFzff59fGTd
2WBZzV3Dc3UIKCwnf7JUBVKrSNyOcGnwILl4E9rHNOUmUNbszllNfZOy5jwz7h25vuk6JpvpxJt4
PBII7Nglrt1jcvKSJBFiuBpb4Qj3iYVdi6PXTLe0oP8cMcklWICsLhiuzgzXd2hW1EZedS1taMU+
3kuM42+I/QtzzLHoCUUO5FwkW643WQJnnNdZalR6LP2Hq21qElWMRlkLGFxLdcjM9ix9rHMz+0d9
rE+yZ+DRUpziT9wYt3L0Eghq1kn0hfTC5xVdC8AvdDB611JZ29Bg1KEvaW0EFvNlITY5ZH0yToy4
AZlHlAcyU/54GnZi5vuR5IGkKUQH36BK3CoVuPjEVpyscLIHEMdyLE60wcXriTNrpCGsEuzGVk76
72DDZLWg74zXPq1+D2c8lqnjHJTZIanvsb+Wyy04g+BtLr3WiRxCp9EEWeJQKP0tgcdzmwzKBjtd
UMToJkPxwjXfXuqjueYS+dFKQoizP/TbgTSSsj4XPECscr935lSkQKHrhiufixzpfiIUuIHrHi/x
bB0H7tMfO0KoUnej9GvxLcyCl+CUPch1qOe2fgLllpxqXloeao3YE/aE/t9DNuMsohAUBWsjDbQB
4EcQ6I0QrI0thiEh+zC+tnKh19PTEJeZqdfiblbZ7+pnF3WglCKYNnK6kLapl5u7Hfi+YL4jGmox
2zZkLx4CCaGL0IPczlDH/VU8olG99m7XWXQHtEDQpdyXIowoenCBOqbmsOsbaj4K5wDi8WfnVmwD
qdYSP1FZ9Via/h9vuhaoDva0igr/SASBwNfSvdZ7k9wTYz5BwAwjhoOFUTsZIXgRWzwAEHxJYG/Y
Mg5zP3/JO2/yHY2tmDtt942Jos3fOWBISOidWwcThyZZfhLyiJ9aEgrJABN+Ppo1c5OPvmSEo2Q8
nGhcbY8zMKIp/LDrBj0IdFGOAA4jT7CINSSMzj54xCyvHgKtIxMDp2YFtKU/UN+P6UzBaARF7/rI
hgORYlQDVM+G1edopwAruI8MhrWXIbqOULZ/5Edgk3csv3RHrTSWtKLBj/6LF0IA0Qa4As82MgeO
mHP67i8fBcuYRbe82mZ9YRUnRkR/z22o8paAHcFbzHCiyxWiO4SwFWJet80xEDPPiDtS2ifJMxbx
ZnF62T7zs+m0BZ64ngk8KU0edlabW6pWBWda4pzSZOhfN/I1H2nxFDkt3QsGF9ZkUyPn6SLJ9DKH
RTaXJwJSvlyZUqUtmseZMgFcQluiNSinazbKfQMGoHrbE6h5zH3phbRUQi4bjVRLc+n70A8qA3gB
jbTeTF8lRx5S1K6oRzZfTMFslXwhp8+SYKkNoL02uBYC+RQTOnlgntX4m1K3HgWiBxAQJbchlOYZ
5FRStVIKmzdxoZj0FU+1GlTCvrr6DJYS2F9nU5J8Ro9/pLXZjdBiLB4wNrIIm5EweMJ7ZOCbGCVG
n7aItvsLKsg0EemQEoLpM+RJJp+5qnwQuU1h2tl0rgcuL+Zw1lkNXwQaedwKmKRjlTckqSTV6GyL
BA7/RSo+gsv2xCjRz8SuAumX4aSy6McIhtjCvEfw/kREFbAs+PwZ7Cei1YBYItilOsrbA2wDqeHM
YAeJ/NMpxC/zaEQiB3a1k09jG8FfPwZmVj/5+r5Or9Z9GOVIby0Bb3AIZLz/AUQcZVvSsISyfL6y
nLABojZE4I2GJ9Ww363MHh2i6YjIEVxDDL7yoexBo31IfI08+oadNqqMxkjhWTJAkVDkzsjN5pVy
e9Vl5RSsbqtG3OOYEMa76kWafGM8nasPeBdu0XZ2wRX9dBzI1EDKgDUXeeYFcGQcfRLkD5f/WRqT
ZvApo8tKBgixBX2CNaooTZxN6SJMMwwkqi9M0p+z/9pNnikmAJOvL+pFvvAc7RdYlQA7HlDCQ1SC
iooBWOh/77jtT995XW/6Ps1KMXl1GtKbayeFIhduDXUJuvHUoaZX7VLh2CehzTgaruZ+BN4t//bq
eiyo1bM63sYu4X4vIU1hxnsF+VNLeOverVR++n4chMHfHuS0O6papUvJl1H2AEOHJq+dfbW7Atpq
hYemzxTolwo1Wmh02giwu35jVtT7qGg+wxyjbr+8Gki5L8SLuZQ14+xYJTcxVfQfp6Q5yji9w8ui
5HLR0W8l8lpeG2Gt+LToiu51YCajPH6JkJ7mbqzbti3xCkY5FmU53xShdTEpfkhhWcM7PHu3neDl
TQZ1AIWUCTZzINzs5c0DktWtM4oKJm9d1r7Nf9BevG6ksbozPTKYVwnq3M4Fi8LUSjvc6UrvUwxm
x6So2ggVAPYjlnSQuVgeQl6ADQI5NhWYrkMX0R5bECYwv7aZEoOhrQo0A5MzeWcmkZkiE1xEPVmc
VwRtEm/k6KgDeaae9qLEk62NGCf96M84L+ieZ1l9PsGGnh6k/TlHtc+huJd+c0bh6GLp7UMYiTAU
sAClKgozgrEc3yxNOohDlOlrw3IbHsyqRatoxRXwwhYN+cVyGjuKs8FXbhUXAxoy3M+n/522Atdd
HVxVC2x6VjEcHeCLAR/m7vZm4g6cMabJVj/iXWrs0a5FFXJbAPaGlJEJ0M2jnx3bw6nLhhD+KTkN
2/9df8GB1qCtR3nRu3efW6imR2/FKdbUYrlu/Ex8Ny2zj1e4/65Mx84VFzVEZoASP856orZkh5aD
e3Ix4Xd8Q1nlsA/43SNy51zroC2mKHUGStY4n4TTuF898zOUpIkvm40AgMp96vQmxmZ+/jfRBUbb
b3PYsHkemvfh5KejTBjwqCjAUgfcq1zdWfz8VS3UdnL9bLo1cf3NGh3eFb/G2yWdpeJoR1SssYjW
KpE4GEgIksc8vHpOEndD+XgOlsQO19tB5Xwq1lwszML9UPERgfsrQjR20wzEdQxxXZm1GgYr7nFH
5ZX6/6wOmnVUeF5qt7NUDwgp8iKuGYkauUHWcRqw6AabymxkOEZonMDhOmUoeTKJtqHC8apxfSgV
DwHUxrbuIvLYZ4tXBsiPaNjm37qI7nHMrHPR31fi/RSGzd0MO48nxQLG3JUq7/opCIJMl8gPSkDF
JaPjHaVjDusXAe5z1v81IpYpu5wMibU/qEvKzkBgpMDmrDWHfWQ2p2Bovj+80srfZKdsIk8CD0MM
ViSlV33bmKvH1QBt+HEoWrj8FmfczM+9A1b9K6FWhZ4Z4tUjOj3bCZ+RNBA0uz0ERdnsC73eQEuu
S0rLNSv9hpZ8QwYTKTqtSnMprv05a/8H52WAiGgeqkD74jXERErGWfEisbeFJcxI45dEjKlB0OZt
EaqrNEgd7hw2WfqWTCQak08rD+rXTqxXCson0+J6Bnhx6isjuGx9ZpebDk7fYD+G2MXHZO7A+HE1
iR/DW2rZp3L4kGAvSorhtquP5Eb3fw23Y+UUvWIXWjT5rMJF3c6LFZLRQNglmAMwI+TinSDgRXJc
fYXtwi+UV7SynOLhfQbnM5iB8F++96Zzsv/unuDzadyuvs3O7JTjLK5rGB8iZDnpU6tUDcn2VSFe
oYo7MeQ3maN9OXCdfkLt+AFkS/XLQ9zPyS/EkUzi7EJCq52L0Gv6VoGFI6664yf5rLxARGRDXm/c
lh9xQbnZuCCeOfBEtvIf4vhF/DrcpeQB/Qg5wrepZgDOQ2wiC/dZnb215c/TZxKwtSQPqZ15Wp+6
x0Z0roSJNcUq06ns2tOvt4sii6gRwaj2Hh+qPqmLdOc4/n9KIGBf99cpVnfrPX5SQToAOKXuIBd6
BtSCMqQO6PWfgXCJP46Najs7zQLciMpspmE38XKbObcjUUm9CEIVlrhZTja1vlWa1aVz8yio+0e1
keOm4Nz6nB2IsoN29C++bk7CQW1kUZ/hxdxi9l9jVabu1Ipv9sK7dH09UVe5tNaiC/yF+dkFETXN
bCar+mM8lCP+/vx6fTzIOo9PpiYfkqCvs4C2n5k1WL3wajahmA23aMXefHrghhSEgmJjXHAH9kG5
lB1b+1BcCw9odo++gzKCyd+moin0xcw/ihIIOzwaqJaOLdE/fwnrLy8S4zLp3zZWX5bIVIp/fUnP
1m0NzAJozkJv9d0GkeWwOv1c3z24md30hVaoqt4n0Z/sh+hUmT5TmGjz9BaWs9kvZyoRUiCQLUfB
ixsboEtlLiOxoeSOsPwivI0tWXadoNwbVVbr6HZQZV+A43PNhuDgMDmVLHkW/KUSs3fsr8MuUwk5
QL4ryWY3Vt72Oz33pU1IvohvPU5djb66MJn9ej54nJn/tgm1RbKLe0cxQMbv6Q8MGGBkUSD+Uz2T
uPRay9hYHZ/k+HzZqKkm3mbN6o8KAiKJPqtQ05Ld421K58jwJB5V25NthndcepT2gCCnPfQRV7iw
E5grioDVzIqaAlAAkL3G0sNowttNToCb1ti2P04sdqJQ5hY+EJmdy9iu7H9iVUOmTmWJeZC4YgCT
gp93xzEABsFV3GrC4iji1hUuTIhkMmMc1rFtowwQXQe4sIbk2SIb+6AaF4BzlIjJN8y9gf4NnpMZ
s89rylpxLmPszCOQhEX/AxJH5mb7wbpU5qhS22RZYyJU+d4LNNoSXMyizwI2SnfmcRhuegBczSJa
5l5lwu26D8u9l+yapwjs505KhSyaOl9qLxJzoCsT6bUnsNCyA0KD1tFjeQcoSWwy7aaviZsDGlQK
P0bK1WJM1N1A4cbZAv5YEnZCudYmiaKB89wbNLu9Rwv3BYqCFeAYtzvaV2OUDKWsWd42zxsLUdM/
MnNYpoU0r7D+F1Ha/MkiuTul5hH+pMS3s4yRvDYvItR96pP5X60Ft66GuL/hOdzrD/Lqp2vlP3lC
R6/twXe2xYlvvy+I6ETOitCtFYcTqaJzCnpN1IZ5lvKvMJZp2m1BiubfgCCDh9mRfHfEMil8FTNF
bu3sl4NyVe6cqSffsHGCvI6gpq/EC/R4dnAiN34RhGZRW0ZPdtOyAeqhfTgQnZ3JEJ8VbSsP+bL4
ecKDu0U7N1x7DXR/5e2NuvJw9kEsbTl5PXdaV88pwAnc8L02lPiawk9EnlQvoRcFCAVZ80yjFGbf
urj/e37Dv5jSL6M/MZiFCURN/cAZ/KPkpzknZBze0wx5PWFgUZ2xNZUgnoKCH5mvl0aOFYnKaUca
cEf5pUeSkJYKJDKJLBlayIZdXuzX7gh0HBg7t1rX95bykw0tvvDJZog3hRzasZ3Lj7402wRcv3za
FLYLGNCPHAVFVIHyKVeN+S+tPWVFYX0p9focyelUg/GGNFwjxr0+199izcGx+T0KV2rd/RnOyh6h
tVYvQk9SUsp2lOTuuQM3w8RGShcdkb+2fRCeeJdmm82gsuIPJy/6XkgvHfuIaX8GHlD9zdDCncKP
miArdY95QpU/aEO1txXsgNGc5eaO1eyvVlAHGi6X+WybsK07sdAUVr99iTqDm61wN0oK5NnPIGjO
Vq4pTuEw6VKr1WWlK2y3v1NfSHzrVTp78YMuGI8Sp3DTUNnmvKTNlis4OLmdvCRkAzHFYEvS8964
6Ut+RWAwXV1YyrFxcQw430M635KcdsNfaHLZ96wXCaMAJNcb0MdonWqCawSzJcLLeArR1GWEyscx
cWTvO7p1yRmGZBHdSEwCgU8AHfaprKrmqKWA9tqrRIdm+BilfrPsBjzznU1T+WErS5HW6XQRyPH5
uqJRoVuUG2hRDqRlzGNyGblD6br6xGJ5ziBGjxe5qYdYGPgI5Am/iPfd5WwQL3tJZ+YjNVF94xVj
5hOGbiVGZvnwFDnPsNdb5acNhATNguz+fxohoC+GlZhWIBIBplEfKvHp/hKL3nI20X6uNQiXAPQW
VFAdhz3jq2ewwv3R2s18ebB3Ntxq3Br4rr2eg6nqgfN29QA+iv/DI4HyUBYOYd7l3byz/AOy6l6U
N3eqHWsIj1xNw2mapMEbG3DIzQVDHSq0cg2vEQ/SYTM3z95Oki8NMwL3cKCeBFL1UvDB5rb0oGnh
/QyJUyBosnprGzf8QExGZXb2NwwQA631Sco9rN/aNULTK/ifphUH00mcD5Serg4l6bXK4ay+LCqc
l6OuSG9VK6Xc37yTPhRPS5KGp/nNiwFzL1zDYMP3J8Bc8VEp2Am0htAm8DF3NXfiGdK7qC2pDRoN
aeG3wolNs9NE7Sv8Yuf2oH1H7YaO8JB8n/hr7U0HEWqGvGRz5obWXKl9R/JEkEPkbA9NlZ34bPmn
sx12zAJgqKEKu0OsPnal4lF5MMEQpkbvrXhAqgJNQAzXGFIXre02HlAqVnaQakniDa4XlDgoG3sH
eHiZKjyVAGsETzOludEuy39R7LD40aVdEJJeE+0lpF3S9vJeAiquWqgMrX6Sdh1fw+0aHJrwkP/w
Nsw+5kxOoTNVWykOdkQ3osMwZ9AWlTwHVhEfr+srOX5lFMa5/8dwcODtxDSmKIUzZ3COpWWW1J9Z
f+0PKFkozvYUfk4khzi3clWvKK9X/XZObLDMaL4AAswD8xPTG8JeYZEqz8CvtGdk7kznFA2hqDzg
sMv8AcOHNAzLpBQFN+Zb4juzi0p51Ky3BFOf9h+i7i3d70ZwZ3x+FJL0tvp04HBexjXhrKUdEmmg
dIWmpAfBY+EaNlM3fH8HFF5k1YvvvW2EAhCppa5vV64+YF521klIzMgJ7rCEUGhArOKzwSIe/NOb
zi1QKEEjtX3aBditTinktIPH2+JnLWUdjMnJ5LFaDVrXpkgAlYlNLiMSdfM2m9HgWSotd9rHnaa7
r4akDFN2mPP6dtDGYfU9RxlWkHwVXogcW5EOjPTcIS2vPrb9gZA/uepxu3xkjRjtX/Cii67OrYwY
CQ4oKiXmI50MCoeZ2y0oCrgf/2jbayJOmz3ge4AHBnW7X8XpvYRvd5H90qp3jnPOd8EkpPz0nRlG
ir1aGSIwwboQtKUfQiJq5hvv5ap4/ILfamfZyn/T0l/ajOaUc+KnHvLlBaI3zwnPLssc5h+hBIRb
oIyGEqmzdlr0Gay21TN8R+iemXl6ulrTdWXE8dMui/ALZ4UIkgW6zc+0Gx7VQga1zPkJv/SEZMjj
qa+BuniWJfkDt5NW1zlRKYHJYVDARiOB1Wvd3Hsllo+o4vAG1m/sfcbzlactrGa9+a17zF3sNShz
AWh5p6glltHSJHC7MHoTArr3z+caGPO5foKpqKOwX2jXktnk6Nwbqx8t9/vU/c2mWwrbW2yeb17b
1KhQOMeiSuDx7GdUTMcgBIQqhhdzwAAuA109J6hRUqXHogkyUdMHGRYJnXaGegjgvE2awvjbqLqD
MbT1hefjFhtQDxHNlH8uWTlpkYy43hYQA/QEO0ip5FSCaMsyLFZvz6PzPUn3B6/+OslsDHaL6aFn
i+m27mewb2IKPOeQhUVo4w35CPvz79qKdMm8nTXyHPsjvV0b1gL+3tHiOr8YqU6Le/yFOMlV9MRp
9344Z0XeboJ9QPuDKOobBSWLaN/vUZHFLvZNajtn+Z2UM1UzhQb92+mTv1gU+3cRuZxhZUI/yz08
xZIqxbZRZWq2LIhyS/zvGqTWKB6YB5MZlKvoDt1LF9HUZKloWCh+iBWDQaz8Ph+WZQqkAaFknLib
N9q8mIa8Vk4ZS2BZgj1f/GVy1jeZ2V2kwFaZ50zuivzXEol7ViIkobRbtfGGX08T9dI6ZuHo35ni
Lx5/PpWn3avuY3bv8HcDwYsD6aLKSdKQX5viyDs1UXBIUpn6Wbhac/20D9Rw97M8CBiDXfApsqJn
iyElU3SENpPgJ6ThBqtJUgkTMhLXj3eoXCy38B/HHHt7Rhs54t3dcuu5DVNwMpq3CiAO9ULFrTkU
1VLN4O5jj/v1z244EFLaCUtl+1SOgdu8OCj3mgK6ta/xcVFqCcVaAAEWBRUG+knITONXQAIyDr3Y
V4p/iFtxdsK0afm3jUMxXD+XVkKFdsJLKV5o1WrHL/zF11XtEIHHHxLQm5mzL+GhIFKlFZzCo/DT
6rG9AiJ5x4eMvRPZXsTatr7DLCOKZN4jRh97kXuu6pG49Mfw3BFPhi/JjxeNlRgAAiAv2R7gnbuh
CF+EaQSK4+c+NJZOZ+C2n5zzwCvhPOpvcORKpGqUExYMxcrMiKpPZ7YtRYxx6y3Hin0yMoKv95Pi
GJYRkR6A8ZZYTR1Uj555NDFYO6BGdB0owGozugbF76dKgyzhx3P48R/rcr8RTgeUWTa4kwUUO+wE
Ev91btJjCMo+6TiF32FnYkFERejotQ9+WKbg1yUY0qwXtkfYi2gJqhwsccOhM1iHUkoi8ys64Dg9
mpz6CgikU+XjUJQPMti+vX/+piiNjgFH+0s+cZNILUgJVccxQGp5Y0xG5onC4wF+8fC15icdbnE2
OEjJdnuSCLFqV4kVxfw4SV6zBpMQMlmilz16GxTQkqW0wF147gWBnlsMhO4sJnSiib7HbHDcdgqt
Xi5O/O+YmmMKuu40y/skCsQvEJdrI9nWGneVFF9UiwVzPBkNIakLbhbbuYpFy+YArNxXgdQFGdH5
xRpRahlfhyIjxsfpsf+R5Ho+3FQ+VTrlb2Vs3CkDSK2HW+YDxUPW3XmPmKQ31AtFpskdXgRV8tMo
UPrNR2nc3rwS+TuHdYWg2ccbDdomRLz0jwZLiEFuIrBUG6/QIuJpV0nHn7Rwn48GePJ73ZstRoer
S6dL99bbpWY7ljGGnngVeV32qRb4IrZ0LDsRxRcE9EGN59IFwWAYXVS8+tUGcVn+Q+02OvqvkNCQ
FF/wlm2Zp4lGIM+vhVI77NhOj9iTGi7lnE8ECgHbQWf5lyp96F7BeDeDThXQNfKw0LI1HzGuUIZX
Rtc6NheHvWBJsDVHCFmoRwh8J/4193e1jJV6TSf2Gx8VyoJDP8Ga6iZLkK78gSLnNSI4czYkY45j
lZ9y0ZV0i9wjlQOEl1j574wPzR4OHrJFEbhb+SWJeeX8qaPKlTA5+BMhwqh1/EyLytQf9ZJlI4rj
j41glnjpf9yWEyNYBLHc0KAjdnH4SZ4mHJ2uuZrD0Hchs+9JpQaxYRhSu6KyXaNNrmiAdl6x4hPV
0JXca1OByue1ZIfKcqdByiD6gfqiGN0z7oDwzc4ejkptZfK4Mo5ZBnixYb4rlWLiFvb5JS4xnae6
InHI8OjjM38z4Af3O6C/i4/V0nraNPFBimEj+9X2QF92Y2UWe6lmXOKSccAeadiAtb+LgTop6JT3
jWg01h5npfqQvCe8C0zcaoCgv096WVCwxNX0PK6ONHllRDt63eiGtiI4OgKx1XpzJCcVVfQT7h2t
/v5/2Y24x+0JbceiCMdXiLudTGvxbFsCuRZdW4b27Fg5T92thr7wK6NiQDZJWglss+uDgFKdut0E
KU6iD9SVQugAAdjeaZuecxbrrbUfJehyYTZkNjIb5rYaoBvMXvfMxzBw/Jx8GSQ+7wI2USL27SaA
RN6nIZBFRawgd4IOwSoWKQ9jqJp6rmM46rAeqhon0hprSxKpFkvRRqDm6s2x6U4ypuveF50jS9Dr
Yi5hRQGR+N88bN6/lCcg0Vfq4nisiry1Og2kBIteI6KxbDg3cDkBYut0zzKBoNGw/THvPxVKhhin
+7B8C37/EqvEPgWlRGVyUbPzPGcB2r9yxP7tFipH0oiST71pGVXyFdQW8xwdl0ybB60hQ/q1+BuW
frSV1LkONtIE9oDMqff939ZhzfxGYtJzR4D4UoyX4OgO96gp+wKKRkJs+u1IiXK0eZH30Q9vdIwH
zEfApFB0gXfUi48OwJQZn3lOiFgNUGh2RzQO001mAtVClaAnBxb0FQMxR++kPDQoATt+OBpqZodp
d54WtXmezc2LSOAwNoblZhHTRq8Csj31PepMA+NCA/qLTBTCgWVQ+qG76wfB0TDqnUYsDmZyBoCL
7BVLhovE5rLGntSRSNfXyO6zygZ7CFGGDaHdm3ZH1ZBaHZicue/+fxD3OQJmomkalvkBImI5hiys
3EnSr+XrPXKqMVxZDe6Y37CVazUeMeIZd+GeajzVCFbZRnuLJB9afbfv+Zc0NBr73YyetNwH+aRX
0YbeKmdY57kLoTPdeIs3UEdp5ZoazErFnn1d0KpDB1EuMLHl126M3uHxpNo6QgKZWViCAotAeGYk
rj43H8z2QQNuJ7VSAz/NpUAqbiCSZEdrxlqcANx6mt/LsEPQv4Sae+Sh6dG8xwbB0Qrg2Vdcj4fv
09ZT5xaeJAhmbVxppaS7LIfRhe6S+fW40bKnql0D7QNxwcL1c77tZkkTE9Vv/diIj3bjYk0smYDQ
+S2ESRTRbcynjyXUgoISwaAXvcaOAG1cQslj2TLwTtw+RJlaEbZbt6LSZsBAR/MM4tXEwpZeOwpt
XVnynaGe/eVg1cVoJk6WcRG0aI98kihJbNHSIURfFNdGpZokPmGMPxxipaV3i3ExZUgompcil0Kl
p4Lc+JQZfBfD15lxPm/DK1h7HCmwIHyMXcOB7if72dgCNqHZxoltf08Z64tz9byWs0y7Yrv+O/G9
DDdfpIch3hza75H+wRx2cgOzdMtp+cywqGmphoFguK6FNEuOoTuxqQwPNyXxVqE6t5fyjIqjjqiR
mc4io5rgPra7pkCy/PSuG9t/3CSJFuyg6f3CUwCJndNZG2nHe83Uhv1sFvsz9QNky27YGQSR7p8s
wPaEL4aseZPsxogdGXFV/9ll7n+dII+tCWcadzlxHp4GfgcC0ASZA4/1Hd20JdyKeCDwb67DDbq0
4B85ySTadfm2brsbFN1cBinkWdTOxB8PDi41CtzeEO/0fFRUQ3YyAKNNIKchfs3/C6bjVwOAOaRf
X6B1nNnJ3wOTngxfQQKiBb9o087eFrJjrac71R9c9alcOUKUeT26XtPsTsGvA9Eq94G7lNX3cCKX
U9K+mW6siSMUQRvOruemNHeQtXietd9Pq5ltq7LPElNDrK8b/Cbsw3f7ZUa+XD6uqenuR5MxTj/7
FmIXaOYUq18qUNQlA4i7gMjxIFkFj1HG2ZEiFfQYJc4ru3MWbLo7vRYdmJa4OKW74PHtp/zs2PDg
OxWAVh+tHWrcspx+FBGwBjp9uiaAUL5VxaaSPjfsjpc4hlD9FmrEpImUSiEBmPPNyOHE/m2o/AVs
1eJzrCPk6nz3mmdouJEdlr7XNKJJAy5ITSKmAqVisKXH3XJp28JgVttRDRKLcSRF7DEN5jsTbREd
mxQbXfTNDnDwnAJXl+hE+uLzFphg9mtoVs9KbFsv4Mk8YYBFd/eVg6DInDwMKiZWAeRSutUyShil
Ieh3wk9AiFAFpnjcyXzMCo64KJT+iEfbP982XKPfEtysHi1MRz2CPeLvqC+hppR8NZTgs7TjAhxe
J3NnIosHzs5Wxz8kZT/Jpx7Z/zLe27ukI0mLxiujpyGFv0UBLQATg83bbARSCMTulnglUgqGrtcO
x0/2/uQaNuRQKAuA40x1wjAKw6LYa8eMVgVWjZsT52tLGR5fx2DPrVX13pGGxtmMEGeP8O8nyo8I
y6SZFNp18w+G0Ws/absbphhQYGnpoHNKRsQ1yF/pPWvG8LbrV8+5qqkm9CUNpoI53JztQQSImnVS
NtHMQYJRmcy8uknuD8EL4rKbwdTWg+ATrq+HNPkm7SxHosSJgIgrudTSdj068twcH3BuOocrYMMP
07tVe09u6nKcD++Ak1HtgMJRlyWid2WWvhq9pFgYGBNYC3tHN93k4JVxOaglpKRRuNy35QVxUHjb
qJv+DT9PHIPiAHMa8gEs9okMpMrdSyJPnzeoseCBvOspznJnj3XZtIOg8lpriwDt4K+xiWOAmu8K
GJSQvxldQ+Ch68oohSKexwSEgvrvgR609iICmI8JzUS1ow8HVNqUg2aX9LApaucAl2pCffddO4oD
D3uL6pRawcuM4SR47dr4sozmmaBCezT81pPTtXFggh0g5PaBpdO+wp/TAAO7gF7KsgXkgspo82ei
iL5+Qc1dz0aXWY+jqA7GkSiy2tlb5kCPsNMZgFxKbBuZmRpERxjptilOkNjQpKMGyznzj7LmPTrl
9sCd3l1Icr6Lhng3DfQAGwzCYfJFZNTYPDLNfZ2JKQhjtr/LPbAZfUZHfZI/DYuGkK0l8ZZ1CfP8
NbStxnLH8L8JfWEMG3UFIM7s69lyDxt/Bn98FZBE1V9N5TlF7+qe07C70M4aGSui78NPsKyrYyRq
HBrH7NAamiCu9gW58RPBRvTGtKSJDICdsTI+/zbzOw3pKSfFI+jLs4MBPjCu3tps7opZzdApEnjK
TrNZgljHEZb6s/EuzcPYKkGztJ4803ZGsEolesJSDwrCcZZ9I3WOUMgp7dlBS3jOPg+SMiiByNCt
5mCvgsjpEp8KEdEPkwjZBj4XUt/yuTb+IC06AZ+dRLo4xyGbz5wwc+87jgUOIALhpvhTKK0ESDIz
WnNBZ5FPliyeAOR/yeXDq/aG4CjELaxWYFSr25EpIjLDxcdW2ozpWrV0Zumv/JIjQRZ5IKEdV7Hf
uLbatjU+CwbYwPqT2yq3LRyaQ+yxQf+hZUj4qqMn5TU66lv08/w30PCqh4EqVCPJ8p++TiuFP+HQ
WzCSJfzK61TcTHBbb/CK8t2bi8bAZMA9UGQrQvecLDlTvUM+L91wu2piaUPVZle5sI8D2urHrEEY
OqmS5L/ZGKsPHdJ3wdoKtjmJxCxiTT+n+DcbyGp/qOuhDOSiWFjlt3P26bpvGi/iMe24Z81Gmkd6
HGDjtDB9zv5JyXIeKIIipKfSoSpsy9t+LV6HrTu2+0zUiYWObRtRK/OHD8tG+o+At2/KfTXAG6rR
NsMYSRxpziRXsG2zvLBlOkUYGi7VC+NcKcLtOyLPn0rzpDGlQ4flZ/ygdEZRsX3xxb18vXubvtUq
Ut+caM8b8ET3l+5Xf2OM+FdzUEgaxMoENTB+He6ubSw0aMZqpYTRTaztQGQOc+zthD8HuI7y6TJY
aOot7tKJQ0H2RSQ3kLRQyynwe1LHZCtoHFr9Z5esiD3iinifwazW9PFnCexbp0OXQJPpCL/v+0qx
QD+Jv8j/6tDpVpPynxs7aOicgpQEFnt65mHVcAuRx4/tLYjJlBZFplATGM/18Zig58Qmkwpok6pd
A2DKbnlKM0esf91k6TkSPiRgqDKSqq+zVc1sLJwLlMIQxJcGNU6jDeXPtjFoi8aDQFiXKcrfH/M0
SewNPqS8vZYTNsCIo+NDUBEV6OTENdU5AjAAvZ0oh1AILuIGQIRNOBCLYK/boG1kfRn2znVYBMgP
xh0m0pcHaveOsa28l2tEcFKi0ulq98QYZlIxtZBIxFAYo5yylS1vn4FTLemdocjB00X0X94gHPlW
DU3B9IjwQpuDSy0VpKXBxp0I8TcAyd+xms0kg1ljD6S+JRDOKRcAhG6TwEcQf4AHuSL3lx+7DicL
DUSzB30Qcf93CeESTzHBfIilSyIT4yjOEciQfgyR/EgmLG4XocDMERiwba3HICV0uEPpnfAXyd6p
gROgaxrVGQPJ0vqFIG6QiZQ9KogDLfJUcLrGwOYQHfnp0peof6EEHYKcOnY7qVm56pf6IprbtbEE
OK3Hv+8XtvkWmRSmO3MjZVFNy3Fb20WN6jVKgJJXDDlRL2qXmabKyjfxF5YJa6U2WMVaYrAfKL9d
vhWM6jwYDydeHcOXXxeTkzYwqyQ8uXBORq0LMrTL0IDWhxulpvaNPnhOXaq3WXajCzWOTyHaKfSA
3GMhwgEGfIuf994oJ/99wxmxNZDHPndJgHCQV3/YPJXvnyRPztDGnJtVECCHg47e/vwVcBkA2JQv
EjeubpgyrZiNPZSOjBsOynU9zIvU6dDQgMlJ7H0VDi9hZzXSpjEvdOyPe/ew18QfDRbZDv2PGuzw
sK0nC3mVf1cx6B7HYSkd2sEn3nZzFc/4K9IAE9lBbne4Tl/IqgNM9qfM4QLTnbYMuraQhtBVIOIH
Vnxo+F7XYcY4fQ9lL+UJxwgoAa2VS5GKQ1YB0y6nd8VIr98OV7FEBxiYHbsjURlepnlq+44kYHjY
rbRICQrACRMc7flfuoHCD2/UajuusrInsQLzxBdSYM9U1OonRrvXX/YvYyoZX7S0z9Ze+CzvPK64
iW9FxtoKfu6fuhsJuPtSFEoto1SFw0j7Nyji4Gbu0zAvyIL4/i+Rq4y6iZM8sPcWqL8XWEJTo6MF
IDzLkieYkqhVQ0xWp5Qo9isPsuR8EmSpK0op1qZNUVhAcrOpVk94Gtq4cbgkMkaWGiggDd75sbi8
9vrNSmjN699E+xGFt91fuE4aFpxom1PklB67YRNHBr/DseCCBXTpJ7SSjdYcI400t82pfLj37ccq
QpntMS3tMC043L3BZGdWswN01rXKnycnTQcb/r224T96o0Kemrku0D0J7j0tuRzAbqWGa7BzO8Za
WwG0zIvkDrGCF8Ixi+SJpAoEP0yyl9nIqzzQpkK+eozUjGKu1jVzYH9zezmZb8nk79teruWJmUrS
AdLRSp97UfItiQg5auBMPw5AOU8JUI3UObscv7PlB9i1qIsgto/zot6SSEW5vHh4MWpNudGC3h20
PZVA+jbfX3Tr31MzUJKL53DDSn/k6/XlHLBrR21neBIvaYobEt/kxhbRp7e2fIJpsROxsIX5NMSB
u60UdWfr10aMmru4Gc9MEoe82CBNVH2CWxOlAYhsHpr6h5+uyY6TtulCb8UvjvxScAw8h9zFgqGI
zuovVkdLVx7HP8QtVIy6zMmSACtzNQbZ/0oA/Lm31JTeRE98k0WwYjfPYrjlqgXDb/6VeTvRNpG2
CdX6EwMXaU81Cbj7xJcbqCe5X1HwyQM7Li/MUtCaWD0hTl1x9m2TJeQMnSieLzumv6SydUBeAr30
9++4ycyXREPlTQqfJKVuyWV4e6jYtOcbU1czWBK3N331B8030fsbIYZaXh0xOvnau7+jb/jVQPw5
Q2AuqNGGzfiL/XYt1reH0tHZpIjIwytxvqhraf+btMmK5EQcgAYIwLC3ht1mkspK+CAKvW8ozzOH
mfIGnS5TqRKN8L8vyCXZiJ+uidE0cvoZyJJRi+5Fg4fo/5nDRgaJq4RSpsgy9Mk66Z6tchsylvXL
tlbKoioFK/P14+z92IrdpyBrqb7hyerAsE6yNtWQjPg1CBpQyaDViVxZMXEKaU7ZAs5u1cPFESYf
Fr67CkoTBBnRZ1FuXH05yLteivA4sujkKNNIuvYXzOoIZETnCA8e+H1z89LBq8wavarV+YwNzc4D
t/0cut7CUjUUoQVk9FRjQzyPuaQTFtJ9Hehu78smfNguxgz9U5nQN1UtKeeVoDrMVHn0PRQkm9z2
CjIisSnoQ16L8IwRlULUd6u2ZGs0Dx/aA57MJG2KMhozjJfGDRFxBmJ9pWBpbPbZoZ+Yes+K9rsT
31DSLzSNK9+3vo3Wes5zmwubjIM8ka3RfdfAws244gFTKEFajXeY/6oVqUrDVG7aFTSMojGMma8g
YXQFQqGqkjSvb47W32VoUT0jW0bVk9B2EIcalWMNkmXo4+k8kPc1PZrq59p/q/BVwHx5Y9oNuz8L
CvVAq9+WFkuCUn/RrEK7dU+vKOIX5gylZFFXgV0H74f+n1YkqPjNa26cFD0TPE9TiMLjcDMuR7UZ
3MJnUwnv9NAw7pz4FhhyWYxGACzHpTAMXjjVzo5lEsanZFDwpwDMf37+NGB050Jie5IsArBKV+OH
8QBpUCAkQ2XLL5grMmXu6mnBndMAmuvM20eZ2Rh5z6rTR11kaGJm5mb0jc8s2z1QuCfkJhpP/iUy
mZXA9AzP2R91m4oRPJj59kBv3kuFXfGqK+hi3BQIzlG1rpywmA/eqfhpKhpNTjNPBKt+6maj6aMb
B2fztbeTAlk95XRtwZH0TovezTUKy19FjHNEgb3tGIILR40ufQ8YZwl0AiB5F3QItsOWImYocMam
wdBKLXYvC34WaLjijDq4SlajvOGsifsGaDo+nUz9KU+E+qdzXoBfzgoi6oqIwT/iE+zInM+FpzIl
r436BM22NB1htPryOz23QCR5uurKURbJW/cEAm3sSxkABlcYdaq2OTFYcRyhU3k+tU2f15KMN7y2
QGMF/KuA38KAiwD1tQiOTw37T8Fa48eqt+vtwLiQ3p7c8z6FxNt6s9Hp4MXaCYg+tKu6+aps1vZo
Lzir3nLA2quMay0LT2EJLqu75aKRUMocDYTagFynKdCQaO8BHL5xVEAN/xqany3y8x2KgGP+lOiJ
DEmw1amiZAYt+kW5VUXuyET9V7DkV/+jTchhFYcN9hkegyOEhVCL6VfnQcTkgyUqDZydg808hJJw
cKWcK2zJknC93QbwQ5wAEcv/bC/MM1dm6cFr6WsTaTy7ufeuUFRr7bGuy61ujmLKdXOFLbsFANfR
Z/aQD6GCznHcQqgpmCyiAq/RVoc616fEUwSA+HfPlfQpjHvmnBDl2ijnwT08ujICMxLqzTaf9Fel
BM3nQP3zXYGa8z8wK2A8UYOYUyFGDeMoEPLS6MtE88P5tX9B/VsnjMoCh9ErY0IB07XBRjKqR9BV
U7CqwLqi4m/9vvzuBiQb2dAMsJU4L/66wSb+qX1YCyUCoftnK9ntHV8cnV6Z4BYgcuWlghdFnige
hA+NF1lT9meEQk1aZzhJjYo+YqLoY1ToOY0iQ5d3giJItUC7L5GocLpoKk7QFZ+OCjFq+dQSHAkN
Fv7TTO7upfpyj6MJJoak8HK38/ZJN4Rij7zpY8OYnYgTGSGqT3eGLbIBr8j6X2+FYOK7FxCiaoaf
Fra3xoWIst0HF8EKGRKBQv1cCvvizyJyOsbf6I94OEQ25FArKfGMw9lHay570zURskWCSeptt354
erevhW5nE0Im7rsIJmnQHyMJ2qf8xYdSlGTgQeS3Jb+2XjX4UF3ow8+d+4RPTjrUWDvR2ZJB3ypq
J3va4kwdwbX2rT35PVjqFy8nDhBwfnMV/KPxafazLSHcx8vqYwEGMBBbFFvBiBGgiVWVTPaP+ngw
CfW0aSTtH8fOKa8BQVrbFJyqO8xTiUh40yE3HuvPoqCJwnmW8I6qRZFEmbpi3LSGSwqz11LnbR++
8qIzNBDtcFnsySUTFRKg/SXhgksqtZLQML5KAlY3Mgx89Rji/SB7cjO53ne3HlEvILOnnjzstF8V
qTvPmRPdkOGVNFxEtJ/acMkh12vNhGVY3Us0dRbeuZmcszQuDrWSNHuyXn+1OwGX6ZKQfhvg3Bu6
U06R+mmVBTl6zyUhP5m9HH6omsXVDl/IcvIywEMgxlIXN15HvzoRtrezJuxwEg1dUnszziZoOGb9
OQebibqAWCPWQAllUyjpMB5ot4yeotLui0JWjA/5nvbFt8/QzDwxSzTq1xFul23CP7oLuTE+PwhF
H3nDF21koQSqdfscuyiu8Dc+tdW9NbvS5JW8pLDC4d2oMUf63G9Va3X0M13NMSgwjwOZeFzICnFt
OYZch3r5iqYmbusaSpurTrZJPWuAgQyS4g9+EaOQ6lD66NaXR3U37HFb+1/Y4Hezkdvgpb6lmbnt
WcjgH8UUcmcKUGPwG/apVDxQxfb8yXLM/2zF2irU0td1zBX/5c/2ZB89JgBBUgOADqQEE97hRKyl
tg4sG0EovL7mxRu7ecGempd0ipKuGCfxIENDv55RTE+R/8ltSWFVpaMP779uI7EOmubYqEVV/1C3
lOtq9eOFhAVmAkC499Mw/QCzUPFEwj9DMmkWPMAfGEUdG8LgMAL3g5ql1gvS4ichNYeM9AcU5aXU
AXV4pLMou0xxOpttoIlCB6Ym4JL/ridzxIeRp4PgmXKBDRBTLH0Uk/99zegD/JcDpAt9LCsUy0x1
UDQuDZ+jmyPuByQ07Eany1LBzd90Of4p2Y20i7+v/sTXeGa7iy5hrrs5fPRkn0XdgXZHKFOLCSqq
87uarsmZzKdCIyqXs9yqJvkjoOG7RhVcMlENXTUb0uzANezrsziWboIh1CklrFQN2OBJPmgjj/+d
7z5HvVBUSe3hPdzK+B94uOO4E6Yi2nUJpsVARYbJpP4y/jn4x8w8G7s5NcXoEt9QOaXlTAQMopqg
drYhC8SYKt4JjlEBLMgesh5ow5aAytQQQo3JQ9wEkkg1oYiVGCCSbjTK25XsYsan833ReCdjyi3X
7nMs1PjJluLs1qao0s0o85sq6T5s8DmgFp66CgHhFiAw0Q+jSiHl1JFMmaYqmXJV2TxtQ7CVRtYR
gxKcyUKhoD8cnRPstIF6kZ2VxrkWX8gno8OX++zVNsD4MEmyyvP7EsJXTehA0iCGB37wC2WTCkvS
Uce4ZGvVnM2C+sq9O/qR32Cfscpg76hV+7nPdk+o3QxHlxdtyW/05DAoLw6/m19GZgpafH7FdV4G
Kw0pWzvYKcaUBq4pwyK+ZUnQhfIjZZTd+iTA6IMFs4c2jBEWkcclHiOukBZT9UBLlXmG5O3I5lZg
1qq9U+OBzq0jvV6UkZ0T2OmGGqOuBTVpzYhJ/Byag8xElc7etnY6sTJ5ajP1OtE5r99OHRiqB0JB
dxff0gLQUU2T9uJ/+AtiKjx5TPQhQwuG08vEeO9wj61FmCdJkkROYkJWeKiyMcWLcTO0smJ5udUs
O7TjhP1JvDL3NPo+eoe4rcGVhb5DJLFUtFbYWS8/Mzk1DSlwP066uKV8BDl82+g6EuJrzeGErmRT
16hHtqybGm4M3zJaHOyQpndxF/GUO0HUbfJcltXS4jKL1bLytWlOlTga7L99KY+9GMLKKE1y0lEp
6cMgU/4obgrM7aGq6/rLYtqDpRNQ4hHZR8YFyzdvTqoLuunAlvzum1de5t+R5qgoUEDRJxC+INSc
kkKpX0m/81irStMLiyWDmBwupGLAth8cVkC4ngctVE46SQQauSmp4uPZcsv7LpdGprIvtKarJPcZ
NKMtNZOoTJYLzPooMdi41sypHDvJTMpBVDT+/JixVj7UVRc941YdZifb0ufPirdEILcVZwHwD13e
YnpWQC6GFyMFjMAt0BPqfqnRWJ0evXVa3pkyCarkOTX57a9BOB3jeyifrkSHq4u7MCUWVKuWW40R
7+zCaSNtAecsJzjTXRqdaPBZRWeJpikHGxA4aV7UqRsst2KpS4BtUWSBVq1J8e0/WZxbrtccN9mH
Bjb8luwAMbGw8HeXOtqsUOSaLCQySQIZI2AyIOCullBf/pmCTRbUt/nr7u//3OVhL4OXJ1oWyNWG
TJOIcRwZtqQUQ+S5/oR8+9lIZlOjq0IixFtVUg4S72F1TiVOuiZUJn4T3jw1oDaSZ8bkjJbrCBZr
lzcEkgUbvzZ4CStXCnW8nKbHgqMO0I4CHnXRnxN5SCZiS+LwvfFZbj9iWS9b6lh4XRBrKG9dLvzA
pCYQOF4LzI3UoSySbYNZZ22keESXSUMR6u2nRrYXqOENSTutPFbb+GBjSz1C/ausIpvbTqI8LrU3
rr60xHlqsHmNgVfFyJzRMJs+jhUq+LSrSwqGK0/xtdbhbbqJ4Ow0kX2V9ovvMOQEok1gEd9yVfMU
HDPluN3BuKyozR/Fh07DKF2JAaKCgKpFih0C+ibIxo3/Sjlaj3WO3pxY9KiENWVftbi5/hfb3TDK
GANjMygPlIXzAizfQjtITW3c3KeVo1U4Y9SdaG66FApDIhg0JI5p0XOr4L5NVbQDRrkjIzNzOhk8
nxg12NLzlMM2KmxV4YHYi7XfCp/amw0qP+uk1sdU8MmHTX+DYGhM0+pRg3LbXCMyHNnfvqhk2Z/J
pMVsYdNFW1qPkQUzsO5+imBUAAd75MdnJE4V0L/UZHJZV4aBXjz9BLjtm2/Zp5oqMIXb3yjRFKeG
nbeuDRo3oS+O72vVOtHgADr47gpVmtpEoZySlf6Ykcb+h3iKpVb9b0k5JGs08o4y/90EvKdKuyFd
8/gvmMSA3drXf/TdaCFdFwGuH4/ZG0gl3i9HiKEykDVfcup90Swuw697F+c6ehQZAVTWeC7kJGGK
dJ7NqUGiJZlcumPKg3C2v3IN8wsQP+UgVXs/VVn3IwQd/uOMNiYLVzzi96u5NR0EVa70j7Fu3Mj5
6JfWQzPlCOIQqNFdbbDqZfQXkxoEERAKI9YsiSnNvZDMcsmK1zFKJLAqPoztjMzOrpXasejnj+wT
QD+GClV2CNuCcst14wLkeCGltJ2OpmlX8ztX1nF5fV6kwnhQ8uXiv7BtRiJwcLCaX++oIoITEwWT
Ud9zAoLUkSqkd+Qm3gGTr6j3QNGyFB7QED7a2vqmF3jL/ERQ4YBMXisTIc1ZHQsdw0CcNwuuDdbM
/M30LR/EokcW+1VclCKYuh+LuI7AaBClDqw97kbCALtzJ9Uk5bUMSsAgicRsk3emSQmr5pwV/fCa
GzES2Hf9dmJTQBz0lwVr86f1ahE38SvJiIPFNK+z3+HCzWB+tyME7Y4zlQVIyG1UW2hK6wYFPNOy
KhETuAeP0h9XBKQpcw0oRVAS40Dos6IELJidaC20EgVeqWptwvWJc1r+TJCJepUZB+JS1ViYSn4l
xRljvbtIcYnkIVB9xhjCFMQjYTNgG0dlJVoMOgWK3BtZxwO1xtJpC+BMyGCnKD1zcGQPn8PwOMYE
uSAYIjss/q8iSBT8nHvnfZ89lof3AAtY0ApN83ENyKMPJlTHXPC9N/FOhjX93Y8jcIu0R4JIz64C
qXcXPFpK7e67FqeINaVYRC1VzhVQrBqDt+riwnmyavrFMkpN5TJU5TgBV7ZWSkLRJI+HLDLLdZ1v
FZrk6VbppkwXhzX/Sm+U4zfKwP3CVi1Wly7NjunRNLldarPGOIzRyx1j8xz7sOk1Jnv/aAHe3/Fm
do566CJ09DUqL3YB+qh+I/04wYW00hhtkbRVBPSY6SYQx40ekv4H4fp+Ok2mT9yZljcAyyxZED92
EyfFJIKXE+kQVA1Y/p3H37HO5Hipya+60NxNZMaGawdX+ElS660UCvMyd/zotAAacUABcYRXY6HW
9OSat0BjlRJds42TOhZUD/fxgTGSvFl0OL2sMOv/ZPXnnhNgxDARyCK2Vs92o+5Ko6deQos5Nixc
uIp3I/2MVStKPMewktNSlkANdkLUu/MepKPGiymAtSZyDzM3YdSzKnN9v9bSdU6L0apzSQL9Opnw
5qeNQIolDmSVMPH4mH8DIk59OhTjU6CvktqhHrY6ducDPujRqq84KRN1MRj9e6PwXL8MsJjSq9q+
/fhirS41ZqXF/EYqfWh2YT10Mgw/6ixurcNeFmgx0VEgaymcC3ojPBwnlNZwu5YplB9VxhA+azpr
px2hilIJrjJbtcMAT2LECmLtP9azJTJMvn1QLJQ+tOCMqxBXWqAU32qlCX4jW6j0PHHDto07kQlU
tqG+QpxdYCiP5GtTF/gly4hVGgDDoU8xSN9R/K5pIXXyVj/kk/tUKQYpe1nQZxCeZvpR7lvToFfl
vGt7C0kGDBwl4Isc+aL1Kfo1T/NT0JM94Y+CbNlH1zOHDMFBaqgBCja8FMgjPdR/uxEOluC/TBAK
F8e8EQSx5Vj6QKwvPW+1bJDqhWNjt/lz2l3YgN//tW08QszQw3Napa9yS8NPlnXP6tP51Wkusfxi
mF3gGjE1rLQzdZqFPkjczX47qtPE1iPo6jXoPKrSZauAWjUVNgBRlgZWS5WjsOCeMCrsBF1tOWXe
gMkI13RENyVVBE+Ca1DxJuRS6zBD8odQ2MOM0V92YHN27GvGYnoJFYsSc19KbjhWFBe2BKvmyawm
Iew8GUdQEL1+qOWLv98wVt00v3118KSF+2cxGYRsAOOTjRi9xYC4Lqqw/s5J6c1XzJwPZ7bN7YsY
l68Q8HRZIWzLMQPHSaK1K3uxy33YhDUyNz7o502IlkCgJ7L5mxlkQYVv/Yn9AGJ4jgzrvAjG/zSb
BeNg8v4ntZ86uMRWKvIZka4Zo+POEPvCrxQARK49wsRl5ulMGo9qJYYUiQ3TTzSYz2rWaDHX/pJT
zpSDgunNRnlH92m1dUjaxMnBVcLjLl5BNZny3ZkYUjRdUENGfoF1l+jFleoomq52beUpeXnCo3uh
RFHTHoVrLUzs0i/pHV+zzLiEh8RzvtKnMiz3SKgmlwxQ7EG76T1kZNwyig81DRS1XUVYtrFftsQ4
TWQhdnDx6uMyZGAHDlHC5LPq08G53Yd4HFHqC/UrhQRK7SNdvHZRbyY2QWFJPcWEfmibEPm2oh4y
EOY4YLnsmwZUIqWdaHk64YUaSQ/1yLrEi3BxPQuKEMGDblLegkuwWdp/7wWBRaDdh05bIsOloLOi
gpG0HWUMxydC1t5p/e4egOnConmzRB1tGGj59VQq1PiUoEKbzGQmg9G9sI0Xi71jgJmjAPOU2k3p
LWQDJI/+20//yYezZ34mZalN49AOJ9PwsWXGSi4WpubDNI7bDBlOiD8yCJYr0r66rDkZP6knfgSc
aNC7S+47eacC3A9IDmhzG70Ptg5ZcrstfudkjbaN27B/SPykwvF024IgvwUEPYZO3TvrzkJz0hsM
/taS9SPIWwcS1j3joBJnxobKH6d3relLRJ1RXnm5voS+eEZflVngWwzMm8eSsupmI+OzZazXjIZJ
Eb0AymSEB9vS+JW+QaCGMMW/VWHqw6nrtRfZXChL11Ey/E8GrBLcm0J1apqdOLq6oOfcOXaXia4b
QE8+hqNcHj5W15F7WbWLOETK9zanGR6SEkGg8LMhH5fAIDdRoZntsaOH5q01eRqethJ7BcUMvetM
JECPIYHVKmRCLEVdHnUVq/GO5f6iu4F0Hdp3+it/JTunIboL6UpIsmltyiS83jl3akHYXVW0zF94
pnDH2R9yg5SfKYGmg0CGVldFsDb1zCf7OrfuOas9W2+V7b9ySULwS0wI6C9SXKcZr2P7WwH50TKW
f7XfQA2OkiVRSOQiw9/2uvI2kdT0qXqj5jeZg988kP+17yXYYIQnxIpkVst7HhlPuB7tgIldLtWq
ZqVmLY3spF/Yshzx5/eMsoYAZx70Jh9k3PQFIXxD8UsKZUIN/VxRyS83BLCIzIEi5KEbC+bIIeyj
kFSiBmNdFEZfd42Cf/Iktnwdi8Afo4YXFJoP9iqEXRwIkAS4T4riUZGC51R9LMnzzC3NwlLcfmmE
hSLvm2DZCvIoJHAvZrdFNafdx1o4V8dobJuoE+Hito0rqtCBlojuA7Ljgbu0A5V7dCFYC2dpBg/N
ZhA8oa6URTgIApLnBigwK7UORTOyEaOfMcOro95AThqFMHgJ0D+mraSIQYpf2HYID+oim0DU/w9B
RJROJV0nl4HcHbQv9qgip+RjwC4hkMLrfWD+evAqc0+VyIm3pCoxzeKavIq1/fxLrrA73c/UiXPR
+2VDDOG7qOKw38bk/Vqv4AdU5lRvGnb9SlES8CehBm0gI7is+d5joeFc5KejBFDK4rWNHKRgyw9q
edgOO4U+A+c89tF0U/3Fj27pM17qj9qB96issPtrSMZD8ncM2ZSSkT6kbsXeQp5yrE+Cz8gXvUlS
CZbF7Lbkho/AAeKKDbkA8WsoJU2pYTFOD61NzdMVeiXPWT8Kyt8Uc5uPImcFKSw+NpPxFJTvDpLW
iYGclv9NTILIg3XpePO/JUYInmOAwtq+6SDx+sQuOd1bKNOQBnuAPC/kYsQIK//yum7l3CCAAAC6
jEVjrqzYR8rIkei3Idj38isGmzdsGqLFfTbDrCiG+FufZVD0iBPFa2WbegCYxgqCMCN4VfX8cEL9
bQ7G5YGJi4ESJokeDUi5cvjZOi8+4+/31jFeExTzijo/Yn+VwFKI+LfK4Q+EI6o3Q7tGha+cmEWo
2RC4Ewx3yAlvLGK8BpIOsa7LQBX/eUjzGPO8acJlnveCjK1HoN8D8Y29oC3ml8KcFEACN7TGNRQB
8pTxqKCOKsMlMPACUs9VeyGCGouGOCTxuRi8ydbTl+NVAF3TrORLspdJ3kxBKDLEtK+QORSHayPE
LG9SDaYGE/aSzY34tdLom7GMtK5NBTkU5zwGdZXiBNZ91NJQ1vWVtadZsOkDD9b/CZNPzpGE9VT3
hGXQwN0dZF0OTgBmHisulReicVBYsvL1MiuFsWx8xtSXDbteQUPPsyWR9o6elycicL8lHH+5csWT
ViAXCHa622dlBVCOGBXn9xHZLVUmdIswPRVAxVAejDFjn6Xc9hlPaqXgnLazRA2hjfrQNiTrrpgf
BnXutLzlzpYtuv4xFNuC780emP7P4eqcwzO5e1aRF0ceqOtBeBguoCTuI9LVUFo4+faGxQT1Fhxn
07PR12AG6/bgNGjjr9OOyr/MEmNRonuw/V5l7RE+R77GeQ580UXT6TxDwLF30q9eQ/7XFyyRFSwh
iOjj8Oq0SgLSuSu/RWEpA5KGyx2czudAdXzrxMUMf05JSVzqty4H1SpftYuwrMbyJqa6tBA+v14u
ZNnhLgmLTmYNvCG449xddQePL4Vy2b9nlmvptPi1rWXYQmHxLbAfjswTb6f47egftgDBFejQIU44
Y/gA5A1xcLLofmNxSldUR/zjItZeDB9VINmeVhH5HmkedvX9wn/RrXyc/Qp3p/xgC3UB8KWU3A4J
7cQK5F0xxjxLuxSzYhc1gkfxG4TE2GCAEB/EwNrqjcf9plbOmp4bdyLSEJLd2IdSfU+7euA4jiCg
dbxkeU39wWAoz25vFDl9fmNJNgtsm4siiVsMqSxsAuH4HvrCenA0adIiqsxXL9xCTi97/fMaBsVi
IwEP8EkF95xwcFEqR33zKCYtgiM3baHd0vPgrRSgg8HBUCiLoizAREG38+nYvhegM0YKdVqQtPoD
g8reoj9n5WSOHkSpKCosFCQ2ydH7ujoBdOMZv6MUx21wd3pMVdKV3Kxv2k5qXH4rOCWQwQQN76aX
GATEYo8qoylZYXRQ3UD5XzlpUAQKhsnSabEzJVpv9nGhjThCjvmjsslLWqTbVCx1FfQCVmHmOyQn
q3b5nALlUDFGF2ujgH5J6/v4oFQ5OSfjFOV+NYZk9ZDbTmm5HIj/rdXvnq4+IBqwMnSsNJTZIHHN
Gey3PRmWmMBrzKUaY7/TGMYhH9J5NHrRuBFCKwibCl67hk5Hgu1UlcX2tHgdU5DhIv5N29aivwY5
oaZ+j3rQVyp18GUpBoCsmn+qBpSclIRWp3MkrCJkXwcyKgB6eu9TXm3wewgKBhm+14UiAuHCIcsW
WRzrwywuop7wW2COOB5Ji8EHvNGnL0R+EA6CRrx7iCTPCo8gT4nGnCWZWLrdt2f2o9b2MlNGnk3R
mcORa7rhzkPsaej6Zd4USwJHzBNJBOY6rYrnf47O5riXhhdFTlWJ1CbH6tWULgJxVTBVuox+T4BH
2atE72dN65esjyu3A1s2Z0OX8/uITxe+j0OvxEsGk39tLbfRd+5h1ntFRB9T1XUwKR+pvBCMPlPn
FinzSsyYX9ii2IoD3SwHtaeDTHdAvML5bpUMITm4vkzJHkXlkjQP3tYTEjWvDvUDvTE4blcBE52p
8rS2VjhRAPkb6tTFNuYXSxlg0NMbsI+59xN/Ol1CALgq/+LnL3T+zpegGoViHohwvTL8eRfL4ZHT
tdee0dqZQE1S6lTvHZoD2wLTjV1qYTTpHYMPh6hruTc45W5gju+kvGyy34Lv3LgsdRu/FBu4DlSY
xO4Ye3nIsBXUyOHgu9GNMDPj/edGYIt1/LJWLO0BrcCox1YThX9nFKKMCHxiCQhkfzbtyMix6wgO
/alBxFMKTvLs2HgHyVTduJSfCT9UfgYnBXItOCH240AjoiXPSvY9ZtKtPcs808lH/jykWrxzHoTx
DQPMfGIdtKDlJZ5gIgzcOFZJxeUgwRRF0scir3oD2af6FS9HZI2q/LSai/uy1C7Z0Us4U2fVbDaz
UZWcJDtN4QFISN1d+B4I6IqG9GW/qb7KXyEvioPlmHL9s67oOKMntOHswsFlEGgcPk6+1qARn4fD
XxJIb4VqaCDgN4hhITrZztd91DP/wVJq4hin+78Us1a1gLjxV9mdfoKpZ6gqc/sCGxfSqKG0xeRA
0eeaOpqU5X5J/JSH3zKmI7dpIFj5lZ0eOe6oqSK+UegulEJWJwRVH/PfVGfqJbZkQfppsZKsGTih
7g07y+3ZYjC6VM2wblDa0enF3wCk8QoUgFgtx8gHd41ycJJPNUiS77YBFt+DTIZW43HqGwtdVeIE
BZmYdTxyZ5wzG4NDcnGj3zUE3Bm4LfjPa8Oyx4OJtD9wf8sXG87GN5qZoGjteGaE/u5bt2a+MdQV
eQUSqsmbVsmLOkMvt+uuzceS85k89x1Tk+Yle1m3TODN18+jev0tM0XBAqcVmpDzveUuErsNzdB8
G+u0raybJ4MGbp9pqVIs7E/eCQVjnjnCuF104RgNSP3S7ePLV53fQpHFqnQqebOvZcCAYC3bPKb3
8/5cG3370mG/jBIzAndDVtJmfA+1qZRgm1ZSmo4rq5emUB4aqh3AmDiuaVkZmyf8ZaxKj+gr4z5d
2Qqvp//DuuLAW7Bm/XdiZ36e4CnYZN+XAy7PRDQ+Kqo9PFCHRpQgI4cc6dAP3zrb1UK+2I2R4xHc
waRpZg1jDroth94Ibk4kHWbCmcRBKUAyGPRdoBaKc0y57/3ZzI6W2bx7JlA6ncX9miVbG1vCAICj
20ueOyjGgzVLMQ/29tM0OJsn5ZFp645OaNa7MxU8IEMjAWGPDFUKhGw13omtuL7ORKyZY7GkStD2
FA+NaJOWV5Ek2UoM/aC36pHyD9VhvpnWEF7NYDWDvwQvkMUUX97x0AixqCyCGShxXoHto/G4MPvE
Wzz10RSN47dH0tbFAZukGQ1wa3r1eLeYtLykqBpKgvXrAYC8jNBQHXvgRqGHCXzoHj4U/kn4yf5Y
mOcbk6m7cnqfSuS4NGkS1glMAF0wZ0knyoFJPFf0+kN5CuV6p4uMkupn8ZHw9+jVUes+2mVmn6yb
dPhd1zpl4p0dVI2oo9VewvHcyXnvLe+V6IUSRUcDSEckmFQNzAM5oAuln3LDDz3QPp8luEsoGAsJ
EFlGrksgjuH4Y4vYTZgz1jBXH4pqLWSlucK6BGEnrz2bIyQHpRNiUYTX1eJEROooPKii6JJNIEJT
WsEQfvcfUCXb2tdkXhZ/2dL7fzqq63NBux7OB1faXd61nPXyt8Q8AWh0sxQKJc46C5UI/RKuhrJA
Xo8e1yt/f2lkK1qD/KMEFxfZlAL345C79McvU0J5dy5TDnNowEEoq2rQ2e9jzakGubacNdoWF4tG
9NXpynkh+cHhIiYfShpZA9cGoRvrHRYaLYHzfMQ7pTSRTjzBmAbyDpCkHNdLe8baYwGNokfMMv/D
H5jKnd3NK21FvaafjjX0mtxfBjA7wwX5X3984Bfi/bSLNErvI309cn7Q0byq+D7l8hPoajmkb3qd
b+rkbHgxeIsEqPFG8yq0WyPgnMJxFbFbn3DgWe+FbjFoIPkM0sorFU5rbwqqQowsPbQ9pr4LSwHX
wfsQCzXWX5WSTNdnuuRBSS5vlXt3eIbwaX9pUKWyFEcFJDc6qqSRlohAAJIsnAqFYaxwHQ7bK48Y
m1K2qzCpFuuC75bTYda+mTwPqpstJYu2L7OzUXrqh3RSwhFEjK9r+A0DzoG6LqgC+XsqOCysBWI4
SotGLYNWZBVcS7oUVMOFpzB9Z2AH250Z/fHuNs9m9VUeDurhUXKqW9GyhqQVULl/c6GKhf5WWmMz
1JH9XE9Unf+HxMv0Q1tQSGQztV7WGvVRz7a9F9bXU2XGP3WjMB17rp7UpYWL1qHCOjkVObf4DIWM
urNVQuGeo55P8tdYiiU2qxQJICvHJELB7xe56LOmaDjz//1W6/xgHMXUClYMD6AzjVPBTiPIX44C
gGywpx49S3jlbKkG9kWoE1oJwFsvA5vpbLiJkhksTsBmlLjxeeeqzeVYZNkKry9SMAK07M7MRH0r
nG1A4hu6YjyzAjA6z2Pcam6uMaXLjc29lChCkR6iYIx8FPau8UzzEatSb3+0cVeukUE8LmjGA+Jx
KKIlSwA6ga0YaxAMMDpp26DmLFoKcVshylDp1wJ835/8JPeORs7wMLlU8MZZRnlAR++H/wOdNNFj
R4QkQVWbQvpqTfM1/F38b6ShqwJr4zPjWl5IC8opOy4FXDdfqHIWlzPjZhjZpfOtgmUNN8ZwP3rx
VHBBI5LX51zDMCEkktnQuLzgy4W+5ZCtozdQiSiWdUor341vDEOfMlDMKmdYRWRV4fEpWtaLj+H0
KbzjfrSiAilnAiJFubONx41iPAbdxdkkz63MaG3mYedrbS/pVc4+6MdjXXOjlcwnkaJ6imXWti8v
dXZfqKxCb/EyiHadtYqFQgg4xwL1rAMlgJJE5jZDC71D+cL6V/zSrvH7sPIRc0W7/kHTmdVUCS0d
KLFsFdO6qcRs6eHvMSdT2Tz9rsIm4eSpOdgE8/HWyXT8i/DSGFp+uCnLV1Waed5/SCOZrwNuMePH
Dc4a1Jo0XUdOx+B1s2GHtzD95vfSxzdayd54lVqgAcq2ulIoCl64M9iiDWF2IHGpXiZ1rWVR/Grr
2iiLCLmi8CQAHUl2DeZgDMKo4xsAKLIYHb3NbgSnNiFnV+IRii/Ha5iZsUyBnqylCPVE1caLc5il
Qyct9jXA+rnoRxQ9Wg3nnldiy4S7Qwu51kNS1jJ3L255RdRefnfL86yQ3p5ZzDqyAY60iFE9Fj++
QJMAnSX2ZIkb8GxlHwRT7ee/VMzEWu8kjDm/bd+zyd3wh/Z0+0XonMwTtJN+0/QczKV1Tbvwv2fR
uZ0YHcuTDHP4mIX5VSGmY3vdyNlmqab5TdW3wx9ER1qTDYu0RjXEwjuiq/pXGvib2Tkn1jnkH+fU
lyO/lUE+Z782e3xsT7f93NXL6cXGBIuRlFwbC6yy9xJSVcnwWzKcMpBySn63TV423CYrrUz5kFv8
FyqXuyNYwB+uxYdo/fOFBZoMtHHsxAB9xL4cbBELgMr0vTasQjt5ThGcIuENDZWb1INqwQqduTFO
n+OpmBXOKbkq70Ift/RnzqKFJ/sCGrLtJuefuKZ6YhY8ZKGcf5O6BcrZUvRzTmouhA+NHg5rfpxt
pKvN9figl3m7sbzpLJME5aunVCUBPn+PJE0LHA1ZYeRZLXqxVmgr4ICi0pps6z+QQiVRb9NiJcL3
J1j0VgL2mmZsSGPRZpI9PCN5kBBnumkxo3nt15fo9s+QXwmhF5gUrfAzsyJbVtrGxBTNfaJwlCNE
SEKYlXjfy52h2s6bC/V2zT5Rp68ZqR5DrV6F6upQW9gWzjGWs4WFSTqotsBdRLb9gO1jH0Hy3tWT
dqjXTyyjTyHlsZ/1KSrshEdTaTbh5wjI77Qqfs5HbQqTGC+2GC/s40hMrfx+735p7P8/XNgwy6hq
WzH7gTIZUMyyaIYyfMuv8wttDa4BONmFhOlzgHJjpOi1Z3KhZO/A34v4h2jlf5CD7QybUo3WCuEm
ufw//81i0NfbRya1Q15c5BJpsm+R3W5M1OntyzpGI+fSFO/2X2cbUit1mdgTvnbYPBiyujbXz2H3
5JiT0ArfEJvLGWtcg3P+X3W4CtNNLyH/U6J3OmTF5iLF9zoRr04wvBfSvmkhLM5BCKu/v2YgkRem
pJjuMEIFhhmzONk8saaLUyMM7YSgpSUZFt623yaqErqRRdcWuBH9pi9d5AXA1DNYm84b+FWph6xY
4PAsP7U4LUMGYYQtOBzXBHkKo30ABSGAxUFbgCOcMb5hG+Bmh4QQIYlRp5QWypfJ4i2rJq9O38Km
l6CGw7ffHAkO3huNS82I8+E7e+QH4qpitGNSLUGIEMECTQNVgaLCZ23YziiiaSP856zi/FdB8Ooo
M4fDN2xmzGHDVD5MdjjJPGtpFkVVjjPillsT7KW1FSZJgP8oma8xA3ARzvb6FdU7mp/eruOFK7Wf
jDMZ4yKM+eQH16Ft5dcmoFtbjzY7y2TtzCnjVh6GCBfsbx3NFt3xND/jK22nWUyTOrgbv+d9qDZG
eYkUuyXFnTIIhMIWYxg9EcCbA1sxsk0Zu1o5s+JQkgkG2lKVWiAPHIJwvzgVuDT6ilkp74PBoGw2
MdqxTdwiY4XKxxMxI9qaF1IECcIgiR9UseWPTqRKNYstbeH9NkAzL76XpHqP/mMwk2se9IgKVw05
SEOWvqmRvAQtDGu3F50JPP0U6qHJUv2uQt2OX4OBVO+J+OTD2E5e+pUQNFCYivfvU0lXzz0mZBLG
1NUazx8DmelG346rjWBphfTtJEfbEx803Z9y/G4w6rXmQF6Gw1WJb73U/RSnp9dEG0XwdG1ad+em
15B7pWet3sK4mZLFuA21cHxpL/0ZVDst9vsOTpgt31CS8Mo0FuAx0d7xDPiZRb6Vn2/UYauopJhK
dAeUKBu17xyYPGxeW3o//Xf7UTQLWMSGBVMr8PvhRiRkxnIb0yISBDCdewA4kKvTNg8waRxRRbpF
fNOo/Xy4B3RnL7YDh2MQZH8Ps2qAtarREGTV56c6G4XH+7lwYaDeGNtzAZ2lC/MGs0iYB2X1p4Xz
FwIKLEpqaqRjoLoisgU3EQDhotNBU1p3lZRtfrIrzXCAzHcKs4aToVC8juiwP+qk96vu6Jyjtsq9
lJ62Ejps5xgOffib4vGV9B8oqfAW4edbJAcR0cJ5GBMO9QNjE1ZSj/luO4r8Du9xPtmqXH4LMrW0
sf+PnLHlR5gL6RUOIJOBmf3FWS7PwRfzxY3z/bppZA3FiCc55voJVI+W3EJ/qnl3aaK83IqCn/E4
3kBLH0aqufj6tJyYY822Sm1dIKQHdfquN++evHPLztGVYBiFCNBOzoBWha+vc+wcGfYLJYoJhZvt
CiM9YLZSGfvb3MyUkRglqHMariHcmbu78zS4XuDs2fpeEXQl7tiBUouVrIB09IGKOz+dGqK4O1AG
U9i64oXXSjgUy/P3GC8MT+XVuNbUz27sXD9AZEUvPbfeX8n6ngQ71jEOIgS1u9j4KBkxzXOf5Sex
PJgd5G10cy6yOcJEZv26SJrVE67gg56WnlUr90EU+DusEXY2soUNpuVJGAXFBnKWY8OE7mPcrs7W
BHsN1G1b5XA5BziQo8gjsQI51ZVGF8Wyq0xD6zdWNrnBVKeNmwv5Db5rqSkqkNnh5Qf228yjU94K
D+NX9+2EsLTPxItGZibm3W7V2yJHxMF4RFAkJdLSVD/oBXbg3u4Qi5YgfnqfVofVO625L2eZhRiE
0JyFf3pLD4wUHweJAjT4ri+k3UvatcHC0squ5rVQXL839A4RSJq11Pzx1tqdbJywfNwQZaIuF61I
RgAVOgskigTH9CfTJrklPw7QNHv5VQg4U5nLn033iUf8KvUB3KUCHJisTVLrYqbEBn5A6KuROKj5
clNgKmhqMzZGTNaxHqBYb3V1p7V1AgegY2z3HGKqk7t6dDUyhvPJW0UB/cniiByr+9ivMa7cS6mP
+uqXZn4o5JeMhj0nYMNaBDTIkiEOdKk6NSPH3hLMelxhI+a96V+9ZMW1raH+jwPR1H0Xf4WO1qyt
5A7bsHgMx9TF4T897Ch7o0lmE6Ufimk6qZp4miC6WZh0VSHSmxP+PhjghEE6V+ESHdHS0gYQSX9I
/L3euNdXeEMYB1F3i91fznsBFcHZPOZnekRMrto7QbLISWvgl44yQTLXWkgbg7ygVN18iXFMJLTt
NCn3RCtWsYTnraFVls0TzJHHkvzKfqEL6/BZfMr7B7zDOtAzEINaI08nShY13ZyysRebSTmnRL6J
+BhubSQt0k0AEKEzPoijtus08vS4rdc4QfekH7EL+74CnzB/T3wxDTUr0UXZUuls35dvnd6pbtpu
1VipC8koCwe4KWVHTD+hD0GZ/w0fAupy4fHdPt9ggWGX6t8Ygb601JoXy32vyJ9dBBX2i5Mn699f
c6sSsLHXqynsB9jh3GFnmxEPfhEwgOw6JzSXgNQg4RjwPvbEpWnUGA4eEnKCHVS4GSLmByHklbx6
M304PVCIDJalnA5UHuosEKUa+O/eGG65XyT3YCDU6Wz7RyG7jq2M9Ep3hKuSmlZvY1CLrjcM+0CK
eDpJ+we81dm9tRvOQJQueMKiYSwupbZFht/251OwvT/1Z3A9D2BNElgepYYEFgRUdJXy8dsEy3DE
+VexqnglNNOGEi3sXjRisRWOzHNaqzYGsUExXJEO7A7DoUACICx6/a64cKA50qXiEYENv8uxRzT7
bBl1my1WQL6/uCagUW+yy/mZwchg2zpnCAL+BSI1FnMjf2ee+RWwSJjAR2xxa/gdC/OVhu8q7ucy
rH2IZOk8NxFszOttcx3X0K7mLMbUl8tKf9E9KvLOlQL7wczjGLmlYBbsVGW6qUTQ0wsx7UD3yk2g
ORycM77s6k2e7yd296yflk2K0+fI71GMC0ePfb+nHBTcPsj2NOTVdVJX3GzIfT2dyp7oa5j2PwbP
4bpf9LaxghpmGu4bDZc/fGnxQ58gAWichKQWRATs7lD/L2aKS24uCBNj5kXN9V/xY74mjNJKY7mJ
dNCza9S8RaFcGoZtzswDJqlJMb/86v0tc4/vT62Qqjwxf+PNNYaUAfvRCUx7wgnV/1VfOEdWcGzz
qMV0EM6GzHioNy8Gqkopu4cT1Ss3A2AjRE3fMckL+4A9uvWzO6Wx53gmqQHXdaLOVGRsbXYJIiCN
8IE4Z+UNNhNAKwXGtitD/B4Dfirs0aV4fbuiKelnVmAUFUGKzXMmdTFI/exsW10NqSAgg4226cjO
JyP1Q8JU5X3HbobYh1HKjUMzabyq7aAKRvj73+Yyz+kYaSqS6Gtgh0IGg63oueLw6zyuLxAGTrhh
PRGPsVPIKZ9zY/pPj+XexVe3HajFqDR/WQ6pkHtPxKavIjRhmvxLMUA9qCgxx7+MUYlTzrOW9FuE
+L81Dd7Ot4Ajwr9yFv3AdC5wmmqRaPUs13vU0MagoqxM12KR3cKT54ez/tA30BdCn9dAjPTzRXtC
MSD9YHvOUxJATtYjCZD6Kdl6Ur3+wtbZ+iF/qeII423vDmPJoBhp0Skfl0sfZQR2mvOzq8UAvyus
PGP0B1LlmwgUqqWjv1sql+iY3fyP9pXjQjUcVYbKLdPc9aWHhwGYz2nTjcsYaECZcqldxR+mVWpO
DH4JALnYVz9kNHfOTeIM+uuusw3TLeaItYK4UZU25DJYjC4TUwAScsVhaap7OP1GQc7RMTNkeMCG
dAlC7MyvhVp8d4z53q4cfnMjYN2KZ5jpSRv5uRZLz6yyOOnNmS/2UDyInwJiBn/0WeiBfJCUnygM
Wu8++3t4NAsB/JbM19Qt5hand4jrB4hJHYdDCXKuKECdOcMXG+bMYIo8Pg5uQitCK8kOQMn+p7lX
EjkR+7N2LK0EyTwgcWdeMRySELXd8U3bJbKvjr6Af3cdIK9sGSA2vUQy+K3epZeHDbJOfyy2+Uhe
Wed2uVy7ZzCwGyuJtP0cfKV0cZ7TRRKXRbE7XP/ErnnLZXLhR3IR64hbQUx4Ifa3U/J76MYw3Jg9
uEmhIM/CRu941bhYliTW7ciR3wgoEe+IhuMkLxWWkbc62ce7phvArtqZK/aZKdOuBsSREPeNnd1f
kOwXm2ifO0yE7dezA8hn4bWJObB39dactO3Hmk9kruzhMp1M0QcfjaDey4DxTKCmbpLvZtoP0iaY
H52fukSnmBzd/PKdnxlCMm3mEt1cJRA9aRnkkr0d2iFkOvCKmcWQ6nYMHY0R755OXlhS6KWPmw/T
BI4vzztnAPGF/DRp64uvP4yNEKpGhUiz+b4yfB5lEw2D7X6YbsAZki8800HQwmrmB9rEzDZqGNPO
TlemSpWfop7VrfZY67uWfIklwGRK70SAGBzrEs8EG5TND3P9s0lmf/5PUOeiDJSjO8hBN0j1rK9V
3tU6CXJXhhp+C3jd3RjzsksNmIej7YAtVjCRz0GEHfI7a5EVJystY6XYGJyNEWGt4zs9fdTV3z1P
H96Jbk7mxaK4eISSh6PBXIko4IqKT0G/fqd6GKILNUm+1yEguzUh2DLm39LkM6A7Q9PGU1Vqlh32
9DhyWeSrzHqaHlg5vsaPxqxgPI31xJzFPM8cLelF7k7me8E7oNz/V7WLVCJB7RJiHN3vXKosm8Vb
PeCzy9bKzJ7pWVvWMIfDqG/hIF7waxeart/L1X4WOLb0OpaRlqcmOxKNVuGHgrjcqqfNCpS8LDbM
910mtMQ8oQVod0DNa3lBoDLo9RITJibam+NRchgEBn/hBvB0rnEJH2rPNRRC4gOqFLglpk3iGCM8
EESnlgVDDvBGttogKFja3vw/SdEQa+oMlWn2XAKRNOXMCbUo6XEpZ3Aco6pI9JsLSaxk611hFIRn
BorPOj1P5mIQWwQRZm5qWlotxHERm3b3VHMHu6ZNY/vJHv88ySE4nSMxcnQOPvw5rOwrpeeGKqqG
qMUdEmU9AfJszWdau6EtSpbKfUUlFww4KIfWTr4A/eesDH2gV/jwkaV+n+QkyWJSTyIzU7xp9Y9l
GjmZiuAHjH1CZheivNQaAMW2DmTXp1umfb6kTN6OxM/WiO3EcFMA3a7rF/PGzySrKWtCK3/7Y7If
qxWQG8Qy+pdMpgIKhHUXvLEC+L2cfcslGQvBC/qfEwpHsyA+U2PZFGDqH28TO4ALflQPljief8em
4zetFd/A+GBTDDnJu8AYrrheJTjxT4mwZn4/q/2mrTRUOC70HSHR3KDRUoeqShvp+nRlBKO2flTo
e49jddZaqS8xKcLp6vxeuqjuBxbxNEn6bmfsdfdwEHFf4x29cNAKttjtP+nqvd4tGLDJ7o5hhOJd
A/E8/j3vF4gLO/2X4DyWb1tVnE6UH6JrCyrSLgc9OOeZi0oVAuR2F6GhWVxl2cvY23u9RfjMdRkS
Rza2flqYhRG7EEmVE1hu1nLYrGZYoEqtT3JmkS++C0K9O9F4mC6gnRZcqZSFW/d6E0LXf3mr6qhC
eE8AHbWqOROyTkTkRb0V79w4bQaTPmzRTxIX4fKlGRyrvQQNgchBTpt7q3scbc9zwzwzYjQGVXBb
MUgOoReU1pCaxLcYeOwqRaxVNTAQxCeZOnhHl3rm3tQ2g05uH8E/bMxc5sXs1LW8+r6aY+25wzj1
vDY7U33OxOOZPHQNGdlJTmnISrcfIx3ezl3RJ73nMyD9m690LjlMXtzZcy8bljriC64ddJ3WIWmr
gPn0VmrFB+ooJyjeHTET09j382UCKIBHvg/xsykUvGAw8jYOwsf5Z9n2XuiSD4V8uXFJ+I7dEbJQ
NIDa9m69paIhzEktH1FHo8pKZ7X+jKo8UqK5syqbPQQDW2o8TJNp/AiwBAF1IlmsBh05qD3ilD33
d6a1UUZd5cogBhCrsVDlfKi+dmFeznqVqWuiKrWooqu2XjRcNQ1PiaRei0vo3MquRqp+jr0wQOdy
m4ixorzSh6QSB1o922AjNaxLAU3IGST++zs9kBgzRHh0nPxM9zKPYCh5nJ99McnTS5HrJ0M5k9S4
6koCpSUXb6nl0l6UcOTKi+1rDdF7RlpJTjjbXyoHAzHTL9fPYHXEe5emFK69xhqk4OiBYZ5hcWCo
y8NKvCdvV6YGrBGbhE5T4vXXu/Vz9K6Y2BQdb6LwswRHqsgL3koypTEHZwHcZsmZRAvgbh0Nz33p
orxQPTTwNimn0lFZPue/nmPQ6IMZZd1+inQ7FGS455vY7CtkF7dPvkvbVcNPajnrVo3QrHmEq5Oi
Z5CRgxxjpek9RKCZ2vwwF8agldGAeJrp2Gy9GWyLMuU+3Nh+sU/59doYmgyo8PTYy+/Zkr4itim7
ZDRQkPizhrUSTNN/+48oEivURTz0QB4Ng+wMlIqrujMTiXPBH1l2AoBsgmZ7N7T8VEZ+dUvYgDYd
Fw77p+fzLVHO0+nYMhsHpuL48M0ktHCPvzHnx0TWD4BjG6PbbpRZQ8bCf6xAqiYXKpVL3ek27QTp
dhDGntfuaq+If6ze2MTQpo30lLJ6IWSb9e/KiQT2uZSXo8CCuAbETcIzWPjliyFM7YzNGLpJ7U0n
xXQkqtsapz1XdOJsX/JnohdQy9mkWzAF6jkbvaUV2OpCClwP376yRyAAanIE/hCVuUN7FITyxgNp
Y03LBuYpJjB4jMM4oysgSaz6bgWciggnq9KZLeA9bznn/o4LiPkT0SD2KdRfsbi/3/jH8coXaSsJ
EsljGfGx8kvYe4EAXd0Rm3GoIqfNxSRXJqqwftbGgkD/TxaZiC55BxwWCx+yO4nqH9m7yvuAluwB
wPilkk0x5rN6F6/VpnDoSCqzGJwVIibUrN2l1dvPNEn1wPLU5ouAJvF3XLiuGmSprtXoUcfsafVo
QBfUYajVZKCKm8kcBpw3nY3AUBnRQjdpHQ+8Ne2yERpMpFdGG+FnlyCBn8lgLxUg/EQbYVWcMqm1
FE/BH0nJ/Vg0+9AasbHOY2sExbGBdPiLuU1cpe+pyt/YV7sz6FWH+wwJqVXOA1Sjo0ddbwTgSPJy
fEobcuaSUaDPanTrL2bpzbYqxqwJWcZnuxyREW4Cmq/a6wnJgNSRyHWU0D0SsBZKVnuZSMpiP5Wk
shOBiKNmedkydZH+egrmCE5RHQMkIag+pe5hERowGQKeUZOdCbPBMaXyq/lhE//zqXwFKtYGybkZ
kVXyw+/gZ2ugCVFfNQqWtJRUhoFJsoI96mT63yNRrnnDa+AU0wIxWu296kBfzg5ZwlrcjS6XiCoq
iTpT6h2H+yVh7Qkma39depEZeQzwYgIxFz+F27AdhNgXAM9ZDbEl4FVtiFFOflaKOLxWCOCWzkka
bpwCBLC0olcZvtgoRmuw5ooGu1Cc5f/6xw1qjCvwD7OuZwkRh5DGZnSyExIruISbSi6fFMjSKNzm
8vBg9aIUJRDZ/7yyRpXwoHHNdCACFElgAJ0uyu1pAiKr7CYKwvsoV09kYQeyDgzJHDdmXdPFcIz/
Nhc4wTqe29CQdbOrZJe2ggAlSNHvZU6ygcq240lUKpeEL++1ZCQmPGPO31bFselh+TaF0jzp6DZ9
zSnvCniztniL+0hLqme5ttnpZXDNHVQ7VRjvpjJQbRzXoRGxCLcuySw9nCV1uOeVziQtnDlEBqvu
brSKPKs8yUqkOvl4Xsx13Ueaw6KPY1Yr/HJebKA20N3b1OotRloENGESC1TEO5JkJWGu0B9Tf8gq
w0wMHQZnN0MWQMiDm3mEj2SOuR9GRjZg80hhT0EhunSqMTshZZR6E9ZMUtPy7c6J/ngnUY2sGu8e
p3uZkifVzc1TTl3gdIiW0zDzHQGlJ1w1CHRd0SvkjTcjZW6YALiGoWqAgmNRERk7OvyCqz+sLW3d
x/Q7iZBncVsAYEa9a8GeeWvMz6AIpv/OzOAcev2cpE0QAJa+bf2YwChgha737VMRLQQC3JY6OdeE
rGQfLMCjSjcWD26Qr8l0mDW1oNkDNw1bIsyVwvaXsBlhv3ep0h/w8rWSueDKdwYT05elHsysdvxV
APAgaVDHNljYbrkq1CiAQBP3bdI1D63Rgxc2tHDTp4q266KisKRXimQd+XHzx9oVYsb4mJZhp4jO
Zdam7EmLqYO5OOoKJAuFw9gi05KqheRYFWdCR6NBoMLYTA5ifO6TDlWXbvdPg+B1w1AXVIMP3hxh
eNX696Hb3hgD3xl41AHRWooZkkXCiyRaoZc16A0gSNcY6duIH7/GhYtkm8u3yTAne3eK1gLWmTcl
ie6zqsbO+C71U3BUBvxi6pj2NoaV91Wnhu9GMFqTSo7au/2VlouqSjBAx1Dn6xxjAT5WyRltv+uW
t2NcN9z8LcjqrLcqPZm9AwH751WtbFxB0e8GCy6azh7vjTyJloAV47phx6pRT2ZkM0GGHGFsgo3M
1X9BTU3y/3pnWWtecqda6WC+YQo1x6oceo6CpK+fLy9QiaypfhrlgOAEcs40S2yv8EVyTjgUjYTr
PHgNMUyhuGIhGQq/VPEI8wusY5OURbvu2/mu/WMA9SulW6dUuSREsJkFW/LGhVrQ/GQ/gCDme8qv
OoefiOVKMsfzkpVpTIpUbju8rLOPZ2INCDoXUm4Wh1HhrUktbNAwPC0Zl0ttoJ9e7JpM+sjCa8gd
5ZImAQ4G85xk1rFQnU6O7LfqD0j6ZA16qOF009Z0eHnVMFACSrtjrAzvIq83P6ow/pIbil20Kqck
TGxAO3cDTT/vqLcfQhlzyvuOWIp1gIxIdwOcNZRVjeQ3qmjTrF6xGzVvsTWWkmhuuHv8KNTb3LrO
mPfxH9IhvnePnoPzu0AwM/tUB4uPiJlSOsvSzKmKglIYMdjs4lTLZ/axCM4FTWfTnSxTULxX5EkJ
8zCg9jl/Lim5kXFM+TorbwcuO1ZYcFgFyp/6VVjcMQqSeVq4YMDNnJb/0u2BSAwv5w0sfxFVAZdb
xa7B5t0DGBPHs75e+W8hWCOA0opa0HgG5RXKFfjBlWvIS6Bmo9Dj25jfFoWhZG1kHuRZAkVvPSDu
qQ6tH6zyPOj+GxGLfL5NMFLUzfN3Vox50/uJxS8FMFnIv4un07UXkMsQXb4ubCQ+QtXgbgne3H8f
m/kuXevNMS63AoDTKYXnLURCuer2YBZvETsI5yh4T9XLYr7giFHzzi1Y/Ro78ZZOOtoEnkE8bxVx
hsqt2na1WXc/ufSXrhIPx6qXOBtSfzQYmIYVH9R0ZgMyNEdAmkQDt0HSU80DZ0D20/8IKN1+etFR
5VGRvXY4kcCEf91v5zuc6oj/xCx8KNIQ5Y6KSFi3aYDKksN6n/KUtAED3uZnSY0CdlOvHxNurdFG
CarPQ++oQibMY9EzzoAGAt8wDxsJGEx4lkfZ/hZucpcYPJQmezxbajXtY8vxGeSJqHjgYJpEOAIu
QqWJ03EZB66gwo69KoLgWToz95S+TiJLfidPqHB1HFmN5tsk6Rjitj9KOmHkYUq26/4bSBOSoGfz
YtPqjoZMVipgF2Pi3bTrsZLXA23grwFe6rCNZnwqNMf7YJb6W/D6xWK1kpeZKmdNe+Y9ZWWyo4dp
kiCNq0BnkgncfuOlSGRcv+NfHEUFGBmipay8BK73Gx6I/Xx3LwFNhKD6LTIGjyhvO3quqMK44FYG
eA2dwxa7HxbM4aom0fa7vQY+Gcg74oldsCmwp3tY0XbXQMMfT3v9Jh+HdAs9WysT8lAKSN+ZN+GF
droQHofHqOt2JjKpbWZMTIFHjMW4P5Rh1FoBzmwjQ8NN40rJfxz4fXkyUBRe0QFdPhjq4DH9VlGD
K2miTyDuEE/zCKn5TFBp36xZgd7NkeqjMOHY+vpf1RAmtUKKoiVwDS43bdNXB0aStI+d8TCxrLpR
eOj1CPTwlramXuoJ1StodBrDA0ZKDUcsiJQIrX9BS4UuNnoki6q/xmaESvH9TMT1kWC8rC4LY5iw
LNUjl06hOviVUnNMUZgNm1DBmLIvAvZ9uISvdwgoOKd2ue/9SI+WIh49Xy/ja5pMp12RyvqSCX4O
iJSUmaVWz31vpw4MSYbj8WWqmLkReTcgOfmb2cG5MMkbmwr5Z5NZyl87C5IIEHXX0VkVxBvC2Adj
e1kJhhNaoSHIUbhqsOiHQjWLlJdGtRB/Oy9riaaa9rnLexjBC7uOm0kg7hMmRCCLGZ53poQ1T3I0
ISzDgcC6bw7G/4otIltqG5haRPWwYv2LTmLl84wz/Tq4l479NOow0bqiHviIUUZgJ9wylL7LeYSq
9letOiaJVqtaFcZI1XgB8GAtN/Bmvn8RqA1YHXDRVkUSp33gsvO9HQjth5ldumTgM9ELpUGVTyEI
ptPqgcQPBAPLr0lpptcD3NHY4zrKiAciaZ1MiPaHwfm+ngARzvgHICpzR8LFFxdXCXp4w3vavfAG
zIBLaWFbw2xKF2MUlDZ2ELtH9BjSV+LimqnAz56RboZaubCJqkCHbt6QVN4FWvj3/KkFTtzbEslW
FKqXyQcDGMLHWcir9casdKamhX/NVgj6P2iWkWykrFNKutSjrlGS5/58aCavO6IbGCtqp19LKKPL
f6fjvexZAT2AxNKr0+wlYD+dC8AmnBe23QEEdSD4Z+jQAnsduaRbhZQW8KNfXGMAL3k2aY9iXzwQ
E9ujbYjAuLjrFuU0p1sNxicipUq3mZYimHNHxH+0SZUvec2yGH6T2UB8PVZI5CDLdDkzQdD+mqpw
egaox65Dv05c8ZGOOiQqevtVmVAfXFtvdnFonQdK6GrEzpgsFj+VNJ78cPz4/HcgYBjuI2Z5AP1V
fGHzHFsfW2F0Oz/34QF//tKjsPI6f/UcKmIDu1t6n7TdOsNvuIHNpgG266d6RTQh5HdgJghUbalq
s2bc+d8JdxZAUYNHKyq5jNLvukR/cN7125DGe3ZJF6lpUEDIhBzBJvhYK8FCmfBQdiKg6nEjt66k
di/5O8kSpHUbJzLQ+WsTFxB0oRofILXOjsmvrTHSsuAVhGB3nqyOABtrPM5simFQNrmYRtWANZws
UE2TfVg+lBSMCYF1dUFSz8dl0qO05ipx6UbBw5gFKsyUGbgOu/FlxzSeL6wQTtAEUldC9tydI2/Q
6kx56E7zEGfriRnQEjTgbKDEbcSYPiEZXQ3mmRPMhdMOGoL0iejJBC33rIQBRfhIZj5JrwQAtwF8
0/sqoKqg+1VGzsfKA82k2LA7GfJE8UNvPxn4NV2lwQrNcvcwZSiz+/iHTg4g08ytkhMSoqVrlb9o
jvIxVP9tbGudrmm8ve7oECpTUoypbHMJ/byvADXMhxhn+wyrAfPob34ZUCBAh/1sxcQUzmtdQpPM
UT5JD1Va01Wuj/sag0jFfzm8XZ3yN3ubOGb18E226XllqZvqOlplYAbIkYjOXW9qOUHUpeYX5GQy
9FoHkk0sX9041qJjjeph0dY11mStEkjBM1qEMCYYMFGaeMemBXvOtPQi+7M0VpgWi+AN1WSayMWb
rSMIIoN1TOBLztQS/TH/pxx0MXabaXXuJJ1f6/wrIKYK3RMtfaLwfFFUEakWU1374nqClY+ISdZ3
qkHNOx8uhyF19OwrfvrEj4xqYF+F53qy/zWveIqSnSdE+gqZjqRuo9gryEz6VshOj5WCx9Ji6odY
gDekt6HjAsnwsyB+IV0yJebKm8CPiEEfVqg62d+vHMHrmJ3h5Pqztn5nhlNGJlutpfTy9dJuZakc
W6b4EbeArvnVCuPBcBVb2TzHA4ss4nljW1C2Yofs8/NOWqY6waJrY27L8mrZGd9QRJvSuyXQKVbe
/peSSOz57GbtboPEHTkGybRw81ZNSqOeXvnWK9bs33rAuXZZm4udx0PV6Y1kJ0QQL0sK3CTubmYa
2kPWLnoCvPPoWt2Rua/kDR+X1iJnL/xy4+DnGiYNE1lFrhsz1LKK0no0uNca5+8nB2t2nUMNZQ47
2y2M2Uqd7h7gWxNUgeqBVZifaSOJJ51FoXuFai/NSmwG0Mj1bQNgoGN254TUpJSRQWeToKOeqk4f
d+j4N0MeESikF/inbqtLxOyRKjEWQh6pr6E9zxJhcs8uA08GKm/zV5IvTLGA/JCJEVv8fDcgaHrf
mfQf4A9OMaJD3TN6oZ4ITgR7WdKdOJL5XVy1NjB/Y3fe1ushSAeh8+KQddDK/8J4kLq/csNtpIFD
FV7JHiX3MjXNp3yqvXBjz7+pP144LR/auNbhApgjOPBo4FBHj5qa66hT3ZIy3LL5PEK9L4ENI9d+
h/r8lcRgq4HeMzj6fCGq5Wp7iluKx46XXlxqDF03yBPy+Mg+1cMep1pBS38olfX892WzDuTgkEvc
N4dlpAOGmppdxoBehFmwurpAh/nx3l/hNCLS+n7BUQa+yv6olWoiuY41Ksj7X96blnAMnJXL1urr
GBBI94oMG1VCLyQzj0vqSfVn2F9x3lo8/EiaPf0qu7/W279H9Q7h3dl3YrEOsogSOEadXzRQOVEC
zEXy2WD2UndnHP4py5mVdO4LTLcYfnuhUBOhObhidlPf4yOc+vwWQk20kbs1uf43sUDW6419+Dij
Do6Bzl1Cpt8W17sDtfGqW2vmhHndFpNa8+ZoDGa+rjYtRiqlSgcdc+izCXfKZ9vPoAo3ueKITmGD
EtToUT5ZmfCILHsMlGpEx7l96As+VoZPowPXqk6rbHUjLAhoJmCKl1rMYf2QGGZUd2oWzQpQ0pRN
4n/dpaetQWAQVn0JuVjFmXSi7Y6InlJK9SWHuy7UBNt4RH1XX72361meRLxW8HM074z8hDCa7v/z
LRMDmuoxTsMcuJBOmaZQzOSZOjLZP3yvBIuyctjdsBFODqeHIkqkU56HF8iljupKho5mYWfRviZ+
mjfq1PPMSnddgnBnIfo2NWsUEcdonZ6FNm+lBVHyMFzIGjPW+kyrLp/EvYvCgIRSpi9gq6JtVu1K
65kuhgXV6Vn0PzPUaQIleEyLDsOlGpoK6YIU2Ogiq94/LifiWRGr7XJ8F/n0tmzMwyCyxMIEIPoV
WiyAxFP2Mj4ceePqPjmo+puo/gZMWINfKZq0nnSAA5iXcnop9dWz+JYLy1y33XdPP6rsxLnZ0iyz
5OTygReMRH85wHH7KkHbtEPHJCPzFzuIDfCuyaofGiu/pJT1dsCxagI1yH12FVBUl2bZAgwbu+c0
FFpEz2E9ph27Mwrejzt4AjxkmiOdksBTCiyKTQPiyIWUZG/8H2YFo0FxtRAjpatQjqIJvyqJ9Xub
qZvNqMfCZyJg6wfRo+v+EoLnXDPrOdezxS/nXZ1W+vHoX3i9YRUXAAng5KzNoiflipTMJ0cs73+N
pgbX4SZY+kVzXsfRULNC9EjBFYgrIu7FSlLOz/Nxx9IFn3X1xrs9Nqd71OUsq2MikEkZF/Kuu63w
oJMndRwPgzVNyLx3AuJgfdIGlSCUwOMGTFWq+JTB1k3dDC76oyhv1Grj2H0hQQDHq+zbxZqjbPtb
qpbdpbhhpCovGcpU2c9fja/bICqaKB8s/R9yc+MIbeGxJeXdItKjSx3R8QzzRy5zODBccnOTwg44
Ss1a+LmFVpkYqEAEjfxtVqn/i86LKqtSswYfpHqEsBfZJlNUH5WuQZ8WdwHqChvF8I1dLIgIMYKj
qYHGcjmy3qUqGmW4ec0Fmw2tqHH8Le7+P1iWWwLIIi3eT1LsdLlOMPr+yFV05QDhxdPVnqHx3STr
n5HAvXub1HeR7fgW7b3t3nx6IOYKAaMYOGWrl28WlkyUF3YnyRnFMrGb4oUBvnSHH0hqUqH4jeIW
01AVzLMHO6EHf2TfLgjp0cexxJi+TVQXf8eTSCj7kSBcGPPy+vU6Ox3msoUsB4etR2Ez0SYlu1qa
zGbK4vVCbToqORjQ5x5O5kkfE48q4OxmWNCFWkF8Lso6Oezz+0fqjpvG9HvkQUE2m4mI5q+JjWoK
70xgGSdqmGxM9CE+K6os1ZjJtCGocvmZbTAo7vv6hPzOjFwLJC9uRPvUbUTsMquskcYs/LaEVtrh
nbUCaz5ZJUlsPU5bL7frY6jbm9c8PLdcSdrVkmWqqEb5n//DbV49JM13WSMcm36W0IF9sGFwE+WK
LXeiggsAS2AtyYlyaH0pAVfcRBJyrjpV4F5U74GRisfa8u/aqBgRLddiCrznDwkfru40zMhfPod+
bkirXHo29Dk3fPwyAleYNUF8zAyeZERwhSl3HTGB9WukelCqB7GmaosyttSSXn1IN+9qkPT0Kf8Z
h96hXpf9ypXAQRbcuQegFDg3D7wM9/bHm2DNi+fDfOYF+yiiaefzP/jIPM++uZYGGHybI/ubo0ul
rHYt5VxbPPurh0lR8k292GEAvKEjsWf7pPeaKw/I2spjEr+Abehi8PWc4XUnUIYvJiZnSrJ1vzuj
Jdm0KDZrlRcfilDAK0eoTcuRAjLYy6sJ9n2DBU5Dcu4EYnRi4t5Gusx12kjES0gZq2VZ9jnaESqD
oPgGWHeIIswMcJd1PYCpZGr0Y777IpOk7J818MONKFOKO0eotOvfTsuy6DZC/ZzTFTk225Azx/os
TB7onkUxlgZ/mWjKdWoprwsgkB6KWVWMhFn8VQH4YjsrhbAVJqfrBovCN8VwoQCoTHwn/DyjU+kb
7xhNUfeXX9BxUFeF0+gKtn/F74hcxjXI7PERKr4O3dflRy+1xWb5WaTtYC6Esv+/IRVtjWl2qmJT
yNf9FlyROo5fKeRVWC6xMqVJ8bn8UEWcuI9pmwOIEHaWUE0EX4WJ1keSR3bmXGVY/YajX2FAj/7w
WGVc17txpafOTzDPXdocyLeN+5dKQXGXcF0xufEGmDBTyjQfJCWzBygNSLeX8n4D4aUNn9xnc0ju
20eY00wm0jw4ZEQF+yR+uKrlt+4amqDrKMZbgpUfMgMOG5YeOUETewCF5laPrOO0jS8bHI6wYwR6
NFp4kkEqZ6+vOH10Uk50YGaTrwyZMtQ8CftPXpJOcTNCmDX59hZBnMICgeiLjhjU/MqO2vz8gPna
DhZYzjWyuAso5OS/oaq7itwiygRj1nBT9q0waCvHyXkhlpNhwXrbWgHn+77Yib8tzZ6ExATYnY2T
RY9QvOXLVFCwADWhZiGHfAA/ZOs4JuatrMHxlpJuYTzymTZG4XdIaStOmJGnUu/5SEhNL4NWVtQC
/Ad2TKok61LJvYcJPEVy6ZL2aC/ZT8Xf2U9xJbVyy63le1VJ46+ri2PDx3i8V7gDbjzEwpcSga4i
os3NJy5lhDBZNOszQbrLpgPMwCK0ii6MR5HtQ0gRQVDc5uV63ZJFK9bctfYHbdlelr1ioo+hZ3dj
V93DtOSJYWvQrR8K3ruhuWu400M4uWcOZXjCCfGZjJ3g7Agm0XrA+5FwD8K84oCKUv43eK4AG9QQ
xCtWFxuThIvtksFjVICTMIm4M+TMR2tUmEwZKIGdZvkePOS/+/ep9Hg5rH5wUBiw2msS7sJJX3EO
zIzyx7x0/fsylwJTgijNsmi4w7rJNvcdhs88I0WsHvkuw0IomqnVmcvEqkd4dIdB5r0Q3kuj2xAZ
+e34wYeKEyJ3to/bjEMDRdZJuzk6owuXBuRUe6GxY2GxWFeSQN8CoKJCpj2NiXU3CIBN75RKbSYL
qW90ruV1TspWbPqfhm8VcvzbomfcXe0s8sNOh0URFkqi5a6K7QUIfh1LbJbaRrtLZINH5NLyQFrg
z74GNFeJKl6dRvjVxY5GVyeQWEekxGjdt8kaEI63sBfb459LTCDiT1WDGwn8+N6RWk7seiUrkwJn
Zll/q/VtH7IzhbbsBJeSvsQyME5wn7QZyhIUqL4SF8hE490Fm4AxQIDLWF2+4xiWJ7QS81UCh5Wa
9KkakHnuihowtQyM/YmfbIFRbz5sLB/XEjT0TLVCQ0d6lDlj2qAUjSx/OoQTFNROAmwRGn/R5ukb
GC2eZvon8FQdu+IM+QUigWJ0/a1CYueGLbEeMbxT17Kj6IAde9rLugiYpN9EapGrzIhG3EeLyUpp
IPeMIQ+20vVxr4Jw59hZbL9aftJs01WyUvIO9H7U1+eHN9nsz1u+fzclcZk62t6EX+EAfK9Uf2p2
pO2eSnnzj4fPZf8Z2iFyqkxWJFC0Y6LL9B8QjU6pJqw6SJRfRndt/eviJixsGkNohcKxL7J7GRIu
0I2coshaT4CSUTr74jsq3UF9+wI+Ia61r8rMIzHmtQl8i1sBObdK3pSgL1VP9GkGoTWopSCtwYk7
2HfA5kmDoMx2s8ji/iCrezJfbccG5vhqbEkjPLFjMV/4DD+6olzdbAwg9Ch6gKIkEw3iO+PRf3w9
71tup/hKJ6lrSe72habg6VGLVNh9oA5rnB7pyAdLWbfP4bxtK5jsBDzI/JCfs12mCMKkIG4w0BuQ
6NTzSpvXKYZIiZF/TOfd2HPAxDiCfx2nMZlLAC8elze3VGD5jYsNxU4Azqdt9Rns0puAw2cq0Z4j
bmd9czmqzUl0f7Xj8pi0s8DLS9FnlAK/N4yEIMFXLfXHmnG3v4wa0QcVvIsaQN6UsulWaDv4QICD
bRjqiO30eMz4t81Or9cmd2eynAP5hzEbPGmJVj9Y/ZI1wsdG5bSvXvalhv9OBnRNA2IbVjGN/T+l
ihJ9SBEX0Gy7dS1SaliqQkd5u8nnjDoiZpeK1LaGWKo9w16Qj2IwBIIgrRPlps3uy9qVb9K72hgl
lGuSKjRS89ltoVCfQ8WjlcTm/g91KehWzL2Hs6hsrO+QWrR50W2HJHdHcWxJplH6+mPTD7AqVGMm
NyibiCcCjBlDRFPuiQLPbCpq9URtYAUJP8W7NVM1I2LTH7jZSDYJYLsp7/xMhuvihRdLeq19uIEI
xonVbejRQy03b740FV1F1DY9WOUCCRZ0zjH12+shqLU69eywNHxyJDz0kge99m3MwR9SfUIze+e+
YJyUG8XRzqhgo/Tk7iBG8qMV58SjY6hcjIQz4i09EzxpHchH/LCsETPSrd1nrdaqLYlm9/Bm6Azw
mgVXPV/mvaHzhoKqBp5+6wPKvHbo8434pwL3m8V06/vCaorTCfTGVcrtTwY1OMtAxUHCdQ4NANpD
g4Bc7y/EaHzkwzzmVrEn1wNhDQpCjcHj+92iEDG8CmCmKzQnEUkuidd6vCPmcIs5GHYC89SwtS7x
9ee/lC2dIfTCatzEzTXg+d2Ipze+SHfXJDeDPbiM2gW3VXISrnx/+yM6uDEPqUHOJht87R+XTqyy
WdOxjsuVyERIzj828jEOdf72Ol9xzw7Hs+TT+Uzn/V7CxwKi7Es7PUrMoRlgaYsP8t+dGaUou3zL
xWGpUP+s+r0s67z96eLEoyfyGrxeo5DzeoeRNRGl6Q0zbQtFpln2jHlEcIFg1iwWR8Hsqnjitl02
VX6l0GcxaFk30BaqadFDekiLBSCI70xcs4RWkBRjmHnyUbpYKl7FDdZahF2NmGsiuuyK0HbAfReo
urZfQFMUGo2xQbuw/MWKoioMG4fXWJCW5DKIMBvFAxa0nv4d6gPYRaTobi89yoreTvi6/+mCb0Ce
irBdt5ojzY6hjYjvkQWf54khsV5cmB5zlEFBLJ/p9CvbG+ErLBf7N4QGaNfcJk1a756pHuTzDFEo
mdkZyUPT3pbBbt5P2xFaBscpPP3M/3K/l/v9sBEsLVqPkj4qDZ/71uWF94kbUci/pHeemXGUULM9
ZyROVxX94/YhGA0my0tqSjQGO5ac5NhbDr45RRiyJ5lTK2XKl7RzQi7IGpHU238/E2aTGtQaazO2
fr/vuerf93w8Mw4nHyXnvCdWdQMMVVL4Q34ymV0IrQ2Rt/hung0NJTcIjobVAzLqR5rOS39lk1Ol
zn/L7laKoguOHQPKZyPTuU0u1NHcwfe9ethk8ls+72cgBXL+AxOU53P8oywtBhegJnT5B2jjdE6m
FSu8TSGZ/OQeu6JNa5o/iU5J6nVvHBtIbu8eWTftu9f/o/DjNCDibhspWhq5d94CrcOzgnBNRcR3
lzTVxCg6vnB6/4uUn7SlfL67CGhUEs+dGS7VgsRejeUeo6NegvnF6Ae06nWn7r+33cloqNmeZZJB
4wJGywuTZZ2fQiie1sD9rBUoi8S1eLZRvMJdCzaW1Do2ka73w/Sjcn23PrIPJ7f6PESrKvcW1RY9
rTsJzDSvc1bIP57gx5euE0N0gw/HFYbi0ixH28q/a1kL5dflm50AwwqSm4wa9hODf/6dJAcT4e6w
IJRXFj3WDnKcIIyv++8JcZ9WRM24JbQkGyfACgw27cQDRxESogAtw1wFX7euQxX9FMxDmQdhMelq
tqUCMvCeaEOzaMU9RYSRGMv8BsNNtcdju6OeTyJhOEd/9PsUPbgyYhijOi5dicOqjTTTcq71eIGZ
SQ/pEAUGh6hV0fk+ZpVzsjmqup4GJgGBNihxAFIhoQWk3pxW39BSq1QOGyjQjWb0EhHZpaa9PHgF
5tlDaF3oxNfnHjqEDfI2cNRcpaxDbc8OWBHCEpCUceJhcpeRuQKDtf48ifmPdDjT93E7zHcprX5X
dBAe1pt4vLnCnpYt8PCLeNRvayr4j21RQ7fVEtbJPuwSLVP8vymQbXgY3M7WMI20pXX5dDtiNuT1
G45gCGKA4DPLJv1QWcQKJywDmNY9dXT1gHVFlXjjR2HM1VLq1R8ntC0QdQBQJFhwm8wpaJrEqB3b
xgqoWBjOWlBgShLLIkdjC1lzGiGdhsbBd/qh+iy+38k2EDjojXBKp5aTNlG9eUG8woHacfeRrw1N
xerLM/7lvw/JUAIGXlFp2HnwLBptMximg46tfopWDmVPvLUjxkCXEsQbRlKXkP0cYAzAgZtRUl/o
EaxHmUTi5lF63ILFF33BZI+7eSlQ8GIxDL0cgDb7Cn/26vViMZah2XzfNRctSwYkGNRNTFgy7eY+
ebRrUUn5g5HMlt9O4Fn88FDbIsiUhVhV4SyCnytdvMLWI0n66TMNoDloQbFIWc9EJ7svc57Cx7J7
h1swjHOsz2x539pTubIDw+6Bgf9w5HTQpfVpNGUuqssMkFqwkwng+TauMiL6RwQWM/0fiQ9xuXBy
TbX2wFAVCLstnopz70D0+Quj8SShv7PrerespiOM2kG+SbU6Per95FKqTCDSZNBuSuyH2252HOWM
IW7Iu485Ul5Lht+hCYpf7g4QmXrze2cXjgqj55PTbuhN9BEQFS3FSHVuwnfxBSdd2n0iTQrutM9q
W+bmI7qndIFSz6wI9NOc5/s2fFbLRf5N+OgRW7Fg0utSJHKC5nrtJtoB5bz2E+G+rWTjfV0xKXdd
VkYJ3so37fbkiRbXRdTXadCj4dqRyBShnnqUhNfHjlYONRz/rHjeciKeMzc0MMYXNN4lWSP0rYqh
GwIcDwA6q2xxDZt+qqKxFfhfiij2Uth0Y1CRQKWupdQGjffvgjtVCH1fdk0n3+DHt5gBW6frWGTI
xVGmM7asfRopHP3fikUtSeMwkCJ2s92xKwEwDBzjfw+pbrbQjYT0tuT0wq8dle7hN+1zYTaNi5cu
B09ibKQpXhwHqFBc+9UPQ2YpxHie15qCSNcMgJuPxBNLcaH5JcNstQ7vVwk3mgJaQaLnPlyYrHGx
HqVjZOUAmZEemSsyPtk4iQjhUHBFOdr6/zLh7F+EK94DD5TlZq71vEduQ/8veuJGJYrAZ0VpNkx5
1HYR7Jgs+qdOlsXraktYoSgdXHGu3NPdlymIvyjpiAw13qucpZaE035NOktbaFyVzFvIyE35Mmxm
YgW/xCltDVXY4ifjKy6XZCnDvgLVTZaKnfzg69+OfMHBaeTQCn72lt+WJcJuSq5cVvZuS7KK0yBw
k27+DzSyfeW7ergrLSvHyxfFTrjPFmQPNSdmxQqygd5NX8XfEYV4FA5jljiUgIjii0n/kfGim/yW
xLDDxakAcN/Cw7qS0aJ0qA2tgaiYqjCu4kE3uagFUlFbJKWOhxQ+n/ih8yUheSebVzK1PcOyXXVL
UZ/d+JKOLTfWNaQLbUoj7ll/YbYzP9gXv4ISNRAP/Ir3wAgJxsNEChLOB68ufiuJWuHzSMjM/ufT
hhNUnvW1OO25yYjf8uc0j7X2ckoEIK1s2CICXqH/oamIa2ZHgjgtXrQgUTC0dWZkDhaMflblQxYM
QKmDKu9Sb5kfJA3vULRF3fZFqBHGPd1UalTahgcyq3B1fvp6w/Sb6F6J0DEY3qiGVP7yBrxZk8oy
QvtkkUpRwL2oE53p2tvdU3tEpvZw2syVwyrnFXlJijEOaFkApuXo2Hpl5ISvctWAqZPTx27IfbXc
Ie0kt8R8krEbTYwoBOmVKcYP+l21wW52Po2bBt1mYD/hXgbdVFkS7NUsQS/Z8DDYqgTKq7gvOZq+
PScqnQRYHSgkNhHQ4po2zRN+UX0xHAWP7l/RKegLKuf2eR/wYm3B/JYqsAY7oRyy1Z7fZJ3RnOhZ
MiEXUFba0N6SUe4oCI+7w3tbq63GNmoEY8laFgF+lyNeLi2HS7TnsRAtKkes+Yq5uekv/pO80HWI
mhbJJfVosUSY3XsYkxZ3xQ+W+VBGbSdkn99i/SiZnKGHDfMJy/BMHEo121/NHuS8z+PyQdYQhcY+
oYO5NXEZX4agzWjSGVUS5S5WHJAAzk49LuB9oifB3BNILZaj3Kkd7iZiWSAUDDSaYzXAuS0fpLhZ
v1DNrOloou158qS4mlCldKs9L/9daeaQfHgyCo7olHtKa0Wjmv1sPK868Ol//jCIBFIK02FnA8uu
iofns4yTFodMnfW9hDkIyX4IJNd5HoYUb7QtzdrpnHE218BRTbtmai0PyZDPAdi0Ji0c+2u5o+cU
TLsaKKGKOVPHOTJEZeHptvKH4uomKI9daW3aj8B/t/lTcznGV8mH8G4UFn+fVPCx4JFPaR9Av+GX
Iryeew4Ge+Nphu5ENPt5FsHIF1fbCP1f6cA3JzTr5weRkUdRC8AvxWjxXnRYktdmGbBxt3MWts6n
9fyINKa5xT1JFDbG1cco+ldk00k0BretwxZab/j8WfAeclZWow8GDSV4pwTXHbUB7nej34TOF3cf
25a7VXLBPBgXNhpzKGw9ccLJQioYj+c3aVFVt79Zq+vcVE5tl7OU0p+I6ictsk8uaBWyDBZwPhs9
5u1UMPDDfWijduItOzD6C8t4/4S/cCmbI+MYaUwOMFPOeiA6wtb1+jS3QEtNg0R+NZ3Qb5jIxAix
o+HZ8cGBB10H0WpPUdvIFUtLmhW8941KGGFGoQwn6JFnLKrbq1klEZa6xwhOz6LwjmSfMnrQozob
ge4JxGZziqE2dOJhHKRcLAw5NMjkIkNJHuZbT7SjcsrBUnPS3VwymBMCuJFyCWsZwVhPHGKpuNxA
sahImXH8g8mFNNb9y9gXCgJRhgJpI4YCk9RCslMbnMSEBV+yo5reg90fVLYEx045u/hJ7zCc/3fe
te6mib4n8rf9mCRrufx2307Yf44tD5txX6R+rc4CZ9kxbBGKJtSk9shXrnhck1k9MtLSNlNNnyUz
aRil1Gp0FuTKnExsRN8F66AliD+CcNg4Sc4H2CuB6Is8DzmV8t6hyZfjT/bmg3iNFcr05Q1e4Qos
3LHHddqPP5hKCbHAGmXrEeXbOvWr/ZMKObwsZepjigCuFfE1tUBVsdVOWsdasBk8sD4R3eLzTYOI
oLqGUCYdlc/zkh+zlIGChjThCjFHAklcnaCBW4DyyYetMZdad5vMRfbTGf15jqzdLOz3Qq1Jbpt2
yE3xUmyZPeTjLIGD2tLl5U23t0xNP+G9ujuvbOez03TahXWM+253Quo8nHRR9PKn89f4IlS31MJm
sxca7nCOFS3G/bW4IheQjYtQrhmo+W8xnWLYdU/+gXCsuo1pQOBnFY4jZDCsSG5XQyEbUYXuiDd3
9/A5L4KNBtRuCmdcezTGdL/mtrbbWupZiFLwyMQB4dBsgjmKQEbzOCaUEEwrSk4bUCpPcUaBw50x
bUEfagdYX0owBLcqFsi25GmHjyNl4gbItq9efu5QA1gdksLC/sEFk1Oxub8YfIJ+vDeFYb7plBRG
y3qWowCsNwjHKtpylg1kzw1sSu/G6Xi/8G2kQ/Z3p2WdH5km1YRdfqdAdUSRfCpGosOatbyFdNfZ
KYBWUyf4TxlQiK7ZUlzCY+XOdpxr7APh7YFmPpii9LrZlVwhu4xxuUcQX0gbiH2/5EN88DyHzRa5
pN1IuOZ5hcOQopRjNNqtBa0dIXLnL+NHj4kuXrWZXfGPJOC+XC+CuAk4GhdEHo14Zka4FWTPKLfS
2LtEiSrrN/z7IQoVDJeYZzSbGkOBMKjHRjIS5JpinbX/e6zU967eO2o5XXIj7JHeyaGrLgnKQI4D
WqC3XwIqyrzFO/H3dSOFxk1JqJrPs5cJPBkrH0yBSbmIHfZAWt4lXdKy3gBDUbhNc/dI40sgsWLm
dMf6GEK3fY6VRw36O73L5n3FWCX5+5KEZGahHFBMXQ6ZIObKZZm3PL7njmUV0nIFFHSHh7Wy47XZ
IEVasKEuO4E44IwbPXwoqcMhdUIdHtKP/gXJwjZl9oh61DkgRr/zNOX89t0H02JCOwklMvi1d9cb
LEFnyRMe3R1d/CHZKENkx1WmkxbBeeIA/62cLHtMTCTAtJ9SBJfzfRD0/cIIkDIRuZGafqs7fzej
Loi5BoxfX7BdtLgylk26dZ9cyT4spGMqF7AwDzR889P3XFo2df5LSJ9zQ4UWAKCllUZxnJwEPr1t
IQ6aXh1e9QaPKFgTcCxlJI0Jaa7ratnOVvX7IDFOanXfCWyipwKCd3C3r9PygL0VV8+WurSUymxb
QLfjJa7eBHQcOjYk4+0VChg9j0YypZ99KdmdV7+QtTCPijkJGprDTugTETG7P7tnsK64Gp5jm8C5
bXclsF8KYTgvztSz3rLDcjbBV58yEL+hBMguG8Huax7ZegrsoF4ccUKHtgA31RyNwkEAgK/n/cpl
BBmyTTgBAGSVDkfey7eMzhs4JymDJ0fgiq1bNKOXP56WJY12ev2CZEDCY3socwf/bxsoDbfStboR
TEb7CXkT5jd7qBw3KfBYLg9ML4Ab/4tbR8AcqsPVwM/4ELYNY2yU+uIf3N6TE3T1WUqp1FNNJ6NA
sNlZ5w9R3pr6Q21gCiV9JU8NUZKoxs4iMwGM++NhLgk0nC0TmMP5lAC6SdZ1NvFMmtiMMSb6ezmR
OlbXPtG5iu9FHH+exRmJ+RAETM6XWgdezOB28+Yvcly1h2yv2FdPklNh4Qhwn8p1W93zx2jGXq4K
7fZh4bqcrmGyGbxQEesR3bWExlMJcXw2VsdGoL3c+RaaKH/PKkvgNPzPDGMKPSpxETf1Pp30Jo7i
p3WIiGj5vFgF41VMU6x4yRuec9n1wBb066qbnNIJGKAmYtIz7vbuDFkftTJH9RTvZqOd/Tn7CmJt
3+x35kfSaYEMnWP9cJ6f/nyciPtkFJfW/X9MLYS6ZIC8nhbnPQrTW0U0BeFdZZyBL6++gfcFXgKA
cELQzeuGQ2Gh5UF4WuNPxUaZWqOP71c8PPs0UBjH5gCF9Yw8bKXYT0culKxQ0W/dDeK0NbWfjR6F
59jfL+WnrD+K3Gzcu2cjjdF9GgxQtLjbpTDlIegM1kvdR/l4wlXElXY+47/sNculmOVlQQS9E/WK
4zjQXi1NywLyXecCblvmlgyeas37z8pVfDDSa6nyeOzPIUVcup/uQYTZZA3CWMhUL7v6uKdBLS8u
CnxgkgjfdRAtkKNskgGcKeP9OrOS86+O4P+f0l5HFtM4PsctkvLgNfz1Wk7AErpI0nwJK3avlx2y
fBtcIwxpoL6ZcGM0X1fePZdl3KGj4UxKfjGgT3Qt7xqRNTrkidVNzqY7Auvx1YuFJ2Ey0k3EculG
NimD3v2yHOqUZ14ivPYSufBkw86xgySkcpZp7P3/SVybZ+K2rRu8FBPhO+LCPD/YLB9HhdfHwlQi
0QQB5rO+2WZIg9sRkX71yQb9nJg6jk+oqAxIdUiZCRVMTGEmfXFx0ifXzR3Vbxo3Nn5KHFQXIVTZ
Aw483WpouyHkF7CdkbksE4IQwpgK7BVuKj6VqOgvwwxHdw8bUB21VHgHpbq1T9P7BqBdr3qmI/4E
IwuMl6tAN7WxKrZ4BvuCV476uBHTEwdwaENgH0IYcxn+MVnHVCvKC49wEM7NT9B7wlwplQanzaqp
knb831E0W+RBeVA9edw7CDoGn0fIBVaYNTiORjuPzy9fbjaqXJv1jDjKu6lqYNiYAPD/54XLY45I
LXysJtNGWda+Ex6yb9PKX8zui0BYsE/fZA80+eWhemGQcHdoPYGnBp7s08iB9f8d6XdqIAdEt6BB
2IKB1NQoBsoh0gcW1nq+6ppxdYyb9d41aNyWwg6KTX/hxdLp4WusNJJfM/zeAV1Xuhz+E2LOTZjq
LJNo92uhw9/ecsGt1fyfmvyd2UnFToSKODGMAj8Kl1EZm9MRREDXQ8WWHQGpzd9u3MzQcE243iB6
hKKwYqCk6X7MhmlHleXUS0vPCWJMjRCtj0HtTaLMUpXus7edN89sTNTChZGADekZwp6zGefTvo5G
sWvBCztOztb18zWn6cpEHJ0h71jkfbh1g4RRKpd/Ig/LIACA2fFAO+nxnzAczNLyGsV7ryKBAIpC
XsUjq0nGGyd2TqtOckNPGMq7MOvxS+F6rREXZvAUsz3iDiWLfxsNXeiBDErkkBJUo44MKbul4A+T
7h0BvKeYPibJK9rdreGg451ttX/9Q8slJPvMvGTVgSvMVFeQIcyXQqXUO4l5Ldintn8pvH92Jc3y
ExV8N3sEs/kuN1F6DaSzBm9ypbCUiCE/7igQaTM54hI5mN+8MokCQCMpYpZQTCiQsymJaf6xlGec
AoSFGeoX1JZAhfgiolFxTmvQ9/2/eERFsEHNIRr+NLIvbJsA1xum1+b02un2w7E4y8SG49JWhg0e
1GEq+2AbgPCcUWX1AtmlOi6Gr8ofVSdU6m4NGuaiZ9AJWHVEQKT7/IkyMqQTHqk1cL6/o0G32/rr
/sPE0pirYU1ayrzn9uv7qExjXM635s6rTgskbdJqWrtAhSVlg2iBWaPaBzwG1IztEu9g0szAvmlI
NE8wFPapEiDOhjmNScHE7Gx1H4hKVrFcU2i4k2UV4y6o21QqBvN0ZLiuBgD4Gj1mXg80vLFt3web
n6aZQ8ddM+y2m+7JvzXDI/wG0bGqfn2DNMTvNcUUX6NdoIUwAN7WAmcXlOitzlkR2wh0yBH1fv+9
+bTO4yhwlqcLVKgkqqIS3zxm3IPe9Vg5RxtMtHh+PIHg6wFFb0p5WFVgGv+E7SeniWAYcWZDo4cJ
mCFWd1+zr9efLrQvlidWjmzkPXY6QXIujfNLKA3RrtEA8xGs/Sz7TR8advd4OYcRCYpcW/krNi1w
x9hGPJefsXb8JjQ6c6O5iLhGwerTBogBbEAI9eEZZXwjKFzyYSWFIzyyVR8R4quo4vI5L1dA0Unc
Jh6KuFPK4fP/PJ9OGvNHe/4XI9UQodfSm+Qqiipb3bsR0uKM+jtDK+hZJ7iGEtsYIkrwIesIx/Ch
nHRS80vOavhVDITUclHArxeVP0v6qVLNh7icwU8zJd7OZrICkY1iQRFZTq3M9XmuQ8QbG8l8W4LU
atVNqv3XuookXZPQ3BnEDcKLKhO01okZFBRQd5uhM7SjzZYjBs3lfMXhkbu162eYYISc2zpn9pkT
CA25PXgT54CEJadcbw3ylRS7AtYjzQULpKW8+ZsmQWjSKxcLRG7KIuzxGUMMC5ppu+2iZY2bTP0C
imqMTphvynCUH4at8lq2WModmIDlYQZeBgbNHHzOj3apK4EYVEFdVFW3zTumKrzHAA/FYBsTFFCB
b1xmAyRKZMe0cb7mgirc1nyZ4vl++m0jypP1fLiQd0YpFvGMjecKhLNLTLnLZHpyphOEg1xkOmxe
3Rj9uZgFjLaYqjUKevqglnXRJNFzhoBRxhvbWuZTrJC2Yl5ESaTLcrmWlu3FC0P7N7Bzp3JZB4/X
mIpLI7ayl0tE9qLwB4pCxhTIvtWJkGcv2QvGQonZCDiiCqnYUw1lBCeOnbkgVmw0YAuSK33p0Fit
YrlylC+ViAJw2H/1Ib7u5uPcl3Ug/WWfksqtjE0fF81qOd9GPy4LJxA/Hyn5lrhx5rVAT15E0X3R
s3abhjPpoGCuequXU3jpJU2lQBftKE8TF1ej6JoN8zAsMM7N/X0v/DtdbcBLt/h9R6swxMOdON7w
SpSD024Ysx/9C5w6JPQ1c5MBXbvF78na63EDYQNWMuGghvXfw9RcHPbrSqsXomCX7RImCEZqVnB+
5eWdK/1W1taVqWbNLmTzBTo0l+IyEmCPazQYUwYbR/7vIEgdnzLujfH75LIn9wpLnt3DjIoEcuJT
KwWN79MJJ1Lh4lyv1IeWfqiTECVUtAqHLLfbaZuoOCyd/5pdtF7DAMYs+RIQbz1yKBi4wlpirHaE
ytqFZ2xkZoXsTRfMhZDV8O/idwta41CFY+k+UmKC0jMOwp1QzqPXUU1DDCijDcreFsrrwz/mY93/
AT7dNsklKBngBl2O5dU20gsGGeJDCqRSSrYah6NrDkyelGqXa6/QInhy/AjhqrBLSswMchNlQJpD
O/B1InaQywOP0JCZdgt7boUakvlf58Y5sTSc587/VmwyMq7hZVvRIOqnn00VrIHanK5+BC/TE3Sj
YAaE3TSYVldRoKcvTO0CP84YAGL3jzLV0XF8Nwi7ae1qYmr28MXu265F92rV3+eDeiU2iA5dckOt
B+l5HhKQGsCa8WqqpqeR6eS28aJ4hXV8391lx4hrpeg23AhjKzsdoa6+vcenQ++hVHvC14SDg0ia
C9BHRnS7UHI20u70n7wMv4IrRvfr3HWf4GKr0pGvvfqNgKJzVbBB48JBFF5zFo21dmchAHXmuCCp
P2dYCCENaoPcdyYNmJrKVlqutpN5RoJOpSAH/lkzS29BsWcELzPVH2LgfoKcZ/k5XDMNHrkbfDFw
rofWQIOT/Fx35d6lhbYsc8WhztVt3O5KqNUoGtsatd1Nxvj4ZkNQxbmG2Qwl0byIsxtQ9yc4JMva
+39jvzNopBy1kCDOX+FxN/K1gIdL1yi/TjQPjr8Z3FYSOgvDM55iGf+lT3PAOxB/YkqE7APP88Tr
lTzC3Yy4WmJqULCttBoNwOCDoKVl4o0Ape7lR+3dxnpHa8MLWkk3WA/+vmiNaQ4DWpUDr2d9Psjp
gYankA7AjX2ZBbcu05kkNC5d3upFQohcnl7H5+nzgo1rtyd07emUSWaVa5iwKEBKgk7TB2U4uWsD
3hBMh2NICAK6djiNPPsEIDEeZfpF1BiYGEjeOHF+yg4Jwd2bpeYd2vSdVsFC0BNbUXI5qaGI4oI7
f6Wqnf6NcSIbnp3nKohOeOo6wBko8aTQckvQDhnm7qntrP1h6vradx9s+GR7/m6PdiTPkueTi+VT
zIJHh2hlXv5mR5GuzphthZTVF6QmfEyOjX314jbQGPRf7vJ3QNqkDFh7nwzrIkazNhr46v9CFtyd
37LocTlgsA5LtqOeEIrPJ1WXcLwq0lkjpRcooGHAILkn7ghO8J9kqWJ0/WxD7eMQ+XfbMOuZi8f5
4YfJqA1DXSuDKwPu/gXx3Fh0d6/a30rCD3H4FBnhjGB0Um4y/jMW9GXbcwfSs74Hn+k75FVolfAQ
J5CRtBZwVJ0BxTHyhHkSOeqQCCk0ScKs2UVV60b+B6PTlvpsdzbKPtD652XwDomuA8HqzZUwh4LB
5f+Vw+DbbC3wnbcF+/fyTlYeVoTy2eyOzPgX1txItzKlMNIvqycs8hIMmLn/l67MjBUozjsQrzIS
28T4qaXqGsi6HmiNmDQc3af0Fe68z32JFTE7byEQn6jzaD/Ujxo9VOjChDuUof2bW9sSbqMCde2M
75D3GAUlYoHbhJWEzxZy7yD1XResthaKxXQClVNv4txiuYJ3LQ9AF87d25nD0+E6rERzA6Heq3x5
JdF6LQaKjSX1JSoFqpoUFtRbJlyH90zgmEHRHxa/tToYKmNu+q86CYKD6+AGs1CFV4aIfrHk+ZVj
qX0PPfQzBNRnQ9U3XviH4rC16yhCKAGEg2CO1jEfPsAdrWxKsJt/6aAEYXThGBaOwAoD6Mw2vWJa
0BcME4Saz1IjMbyxc7NOQnQ17cjaYAFfW8/vgyZNEbsDr6Kl22dIvigZIRqAhQpEEu3m+aBG8Unn
4OhpykDEQyQy/i35KN47rJHPtivUNhZvMzmiiyI1OGOqdH9iom1l8AHhV+TxQDINSH2AJ05nmFY2
UfcATvHvSYGyOE0wF9mP8XNmZ+1pCNC2/KOLJVyZVgeW6AR5p1W7gk+lk4rts5UOZ5T0RZtKIj5A
auiIUMMN2ssmB1wzropefUylCV9kl9P4qyG6kqBUUKlzBWizsm4cV6um6ohK8XM0h5n0sfBW8Xdh
VC6ZQReM9J9EYSgnGUa00oB1bT9OqWP40xvXJyvH6AbGKrMaNLN042cy6YtLizMZelJfYV3NT2VU
hEImcTitdYoKBTFvlSKWURBfFmjh4ArXypkJ7HyEfqaB5HP4eF6tAtwQORxmppXut4cjsLJmGPjx
YbuPt5KGXcUUDZpdkRCpeh4+m0hAX8X3zRuI51T0FOn6eXO/+6/SjZ2H5x7oppQTewabVlXEcnsa
5G47/1TwFn45UpTOgElRDG4z8voMdK09dGJusWM6KBjKCZzVu+N/X6nLrJIJtKnnFdzD6QyOopMa
tK/htCGu+yE/yV4Dow9Ea8kokOZk0s1LsQYlqCVtc4pA3XqonKNJVCu3NfikOHep1dXHcbo3f9ub
XKSvvURO9f3cc5YsIJuQSnD1S89MKg3ID3ICBwIXHOWZuEHlJniFkub0QTtbtuifv+tTXIcyR72J
VCEzoOF0EHt+NI6kwgjIfS1HYOEyC9Wvsgr78eYN4B7IObMu/HPKnAtha0mTfDZOx2qME1G0LdRG
rfpwA9wTcrGlaF7KHcvDIfY48XacQzIaSSS0V0xQQrpFutpNe1UY8vnLxThoF41CUH2tAw4GP1ig
Ya+YERmJ1xnjmI/ahsUGzqzY+P6d9CwUrgiJbP8l3hZTy0kdaYcu2xDzaSSm7oanTofhWmC2jdF7
CiFDTf3iE2F6xtLYy6Xjb9zvT1pqWhSPjClguPhK5zGjH2+G8rtrGLx2smZqHO5Sj0A4aLh9vGt0
nEmsbTEV5yVxrw/Ck7K23UGW1gBnTsQPhanuYjrqDUw9tWlwHRlLtBDAbpu5gbi0Oop5tblp1Qg2
luLHelnWn8fFFwKV7ec/mcK6f4gNL+f4u6sHynWb1OmhtzQgZVrMlrNU4eU+cALvVJ+tRO8Ijp+h
hZCbt0zjMMYAUQoSj8cDitWcvm26mGw/JK5PoaueIpH2HKi5VrxAfhWcLBu2XtVv/xO3kiFFZ2bH
XHtU4zyfj+hsO0k2DxTneRQzcM4wkAL6W9N/oAjm068D7jmXOelOdyDyzlQRaBAQL+dO10Xgg0od
bTswp3W+mLPGNUHRHxwtKfIrHWBJhPKZL7WFjEPXqqLxMUiUZchvdILKVovCzRjp5kVgEyMAcWf0
8YQc2vKrIM2qrI8m2ooaSbVo3Zhor7nAXOCcNxcMh6jq2YLF1nmsFO/4Pp45VGrjWHGdyur/nfzm
v8cpcN32qFp6GWXSvkOy/YaI1vM4CGd41SzJKoYUchdDt7V5mOTrB8fa05vO3kcwxafH3Z9h8piS
2SMhPa/dME/YXoseqR7ZLll6p4Mu4l4WkFD/KCI8Hl9yk/9v+QuLCFTrxZ3RnPgRh/MZVceId0/T
VMWVS0a0rmFHxOaw0d9zRJCSQoWHbNRgFJuWVW0+Vx3NkzqMmMw/gfRcr+CI5+iKCm5qFwAqvpi/
+gy3JfzWvU0I7GWQkw/+eEyx4RaB12JFScfywCumJcpfXjnw18u0fWv4/2G66Hvh1Ei+fRyjpBEB
vcLM6Hqc4zEWPDYiqkllBZ4jjDh1jI0TCfnmOFSHETJHh8mzix06apaOvq+eJl9OSI8V2es5Vztz
3bbCtcIZ/olZuvkBIxO/L3yAOJ+S+kiwUgQZRpBH3fCMSOdGVt7nk6ru1E3wULehAiYZa9H9zg5w
3ESzL5/iYkkccuDGCPqM7w+hpcTle/3rYCa01bsteI5o7hI2II5USW8xc9hGjS6kdEqDgy4yrNAm
NxuGeCq5ffzVR2iX59+sVNa5iT5MKVzSvqfGj4qUmkl4/13XAB0qEYI4NPx/ncJrDIlqT4SIkPU7
Zhe6/FzlAVtTMVOhX5APEvfBGuPjHHySmfYC4O99eNE2v99JIUHqlVUsZoYF+yUaCIXdXO6fuLtK
FGr5FcptV0rMYap+CJ1hO7lrAP2gbPEISROH9FcYCCdt4rJktOFd2yTKE5n7MwTXTV0OmzT4Qf0u
GdDgL7hutpD0PXviOTAeAW1W3TzFs21ItI5LJ1QnYUnSU9Rm13neuEOs/KqDLTLM0dXEVmcEenZH
BRdqoGS2MPA0j/ddC6kaCRQzWfWGPlcLYH1Wk4+HVgmd8xC23Ss4R+usjW5JL6tcHIbHjq6VaG7J
HJVohXOxct6oEej/ECvB4bcBVg2HQun/jLNpiJtr5+aB2J+tOA9/z/2BXpSGMAfVnpD/GflY0KNf
0b+NHd4vQRdpRYXRnUgV6Y8Ai44O6B1pnAnq+A6uJI7rWltjfuZyIsRboi9JSIdmjbyjTjT7x4kM
ydQVozDFQ5djEOHfZOuzI4taKiso+IiGm9YDqQ9seZ2lC0JUrPLDRgtZL+w1IIxGdTAYmpB8GYRx
vwqZnx0rz4KjATaJQt0zR93Erd9OSCz6Dl+B2Dq+TKV+7rNITRnL2zHdOBq9oACaAGa6f29IwNpe
9RfFgxIbspsToTnMXph2itiFhrNFTaYa3tF7RWGyRzM8nBBdGLenvtoi/dp8TH10iK0IhN3ikN/p
A1BAtNIOyxDvjUbRKMNwVmm7bm9Zf1C8LfpEe/g7e78l7Ybzh7B5k1uBdJNYgEON9HrkDWU9KK5U
eFEG67mF7G1C7EUX2xBwJelqMN1LIXRo2fbxT4HYk9/8xakBKMmGC4EFAy0W0RV5VuiSr2Nerpoa
1tSMH9EtXLrXfeq/WSTTOCV154erLBwmd4WRn1W3jJx6eF74yFfCrcP5w3wONAbkUJRJf3SG43X+
n1KFxrCCPTG5Asp+dtJb9smxoFRfHSl+91ZTdbATZX60YkShCuFsv4M8Yl+6nQ5Z9/tHg/EhZWpa
iYM+yzfuAKrZis5Qh8xUpl7DU6US/pzZXXx32KTBfkCg/aM6+m05lSUSgt19CloynzlJ9HVzZM4s
00vzgrTpDhrS3P0sYZ6RExmdpMMhzs++xtUowEumftveh95EFKf/zjyIMMttzlY0So3y/LUZgRcR
mNIwCffCuaEeX1IABHxeulN+wAuZLU3hlUzWlubOHQBDeEy2cWy0tO+ejdrWjKn9qI1VF4k8NG9i
HGIMI/rztt+7Su+lampimTE6OPYUq8BP+v4tjtc+p//y5ZfAUQFw5GaF0syLk6sShFE7DArPdUOQ
51fKah3oqCtq8vVQ7LCV9YG2x25KyFQYbzUBwJQ/GDkiLNZZfVSyKJlysG6vb9ZvgIpbm0L1RXs3
sDvUMxTzuKIIn7iYFQUe950D6YmKqTPsdKnztNvtuz0GEq36sGCUP/FU2Y++TR/KHGiuVj86V3yt
2zF1WfZv4D6E15DzzPoFXqsou+g/hX43vtdpBc9p4U5x/EMnFuNE1FzYoyQgp4q2Z9Ozb27C1uWg
H6uBSQokzqpbLZJmsqLuPE9F+TrprRL3y8jJjAMPI+p+Ce1hioiAIsVLg0Zd9UeBk30DyU/6uNBr
WmNoqlnRMWAvXlQCk38kNKMZP92K3js9TQ9DcIV63y2H9FpU6qZ1bObmeqbqpuanxvsPeQr5bklR
y3fsAdlBGwx6wjgHVjKpr9L2PT+p40QHkA9jgdD8NZ+SYwD4kIjm+dmNhjESh1laxW6QV+9lDAgQ
SUgt6WcMOHpYssyTqvMRVCvKQWkAKEjv/h12oAAELnRmIGGrw1qDA02ar63UVOJEokOFYW5MjQNX
rrI4qnkrWO07iOSNagUo0A1tO9blUCmvrcf8UtOB0YtKq76tiSlCvS/xl2k93MpSWB9XSCU97i9n
pgFDtz94J2D8XDuvoppeM4Xcxs8tMqM5X57YILn6iDVmA7AvRLsOYmgSWGfkzx385wLXk/6K/++9
3NMazQwLkrA26Ts6DlQAZZD/XWk3eeZkRlvUA9iF2tX6l/UjYjBItAjfbJmO1laS8I3Feor0suyC
frtUXwMW3Co8q1oKHHu7NjjyB/dLdoWQy+jPNTKWHnG8KTXnO0xQxinPoqQR9CjwjzCmO2czUSSr
hBmtLLHGVCm+nAd3kAMUTGDZJz58g76pmbp509EV+h+aBxcqS879pdklpRDrfXy3jVVPQ0Fsf2FD
VQ3Tqhty6n38RZas/QamEcPhD+p/3lpC3K6kw8hyMzPAgNFXjwCUqy5xOeX3eSJnwJRE7zNTigje
hDzzwKX7hnUDP7MmtBRQWxCheVifkfzpyZ4V7qDDjQnYYuznDAWgCM09SfWokSXIlSGaLW4PkM3r
J+tIlggdIT+gDatL+GTvtWcWhlC4dJ8Ukn7VDu0Z5RpMoCO6xOv4y+k8F+VM5zjXFl9iIi/LzHhR
aUbMPtvndyOrfC/wZ5wue/tWat/RgjcLJSVLc/D13Wlgb2Hb+c6EkgbK83EBQ8mWGUnZCWKNiobw
8K+nkYgg7m6zLnzVmkJRxBPgVVd82jD+D89b4r4oCfSrdRqq/cMdTGiUsUATkOrtstBM/EKasW8K
NkFeLwQuA7bamWebCD68n2/xLtZHADlWztvXs37zkR/oEp83oILPvZwyvtknJ15FfOH5fzbh0l2S
yx7nQv95PksU2U05HIEwJW7/Cbe/+HVuRdwvzmpmepPSPGW+EgEJJUwswhzOwazRMmfbLr9Z16Ga
b6iuavA8G0PT9Yrhv1O4MsUoS4PAEZ8uCAaZwH4X/GE2D1wBzxjP6CEEk2k1YAcDlIMG8eMn8mPY
DsH7pXkj/VEz/8Af84sB2YXZ4a8M+NqDEuDrqbH16+b78/phZLrS+5DotyTZ/ViuAUt4srvEyvAM
0rAXv7E1zfIlVxKaIKyKTJwM9GBh0u+rVqrvL+dzzHR1f3kDRPG5pQ/sOceC0HBX+LPzuk4584Pz
8MqQf2vguqYvMZeyIQtuq+V14RgLjNghCCFK0JHbQaknrUA9ZFsGKVnJ8RNZ3SXw5BSEaKaiwDPJ
kKi+Zy6kfZ+5RJlDA9bMHd8fxvMnx1m4ADyhdiw95Vr/a3jsji4ONSkMk14U69FvWgSYZe9NRU7l
bQAbkf99pWi9kOu0Cpaa7pDKXIhvKapeQ0h91wfwPCWh8Pci3I5EgQIBPFw24gKhloUKGtw8Ily4
OJpaRBZlbyWd++XiV5OmrDEScQ92egsRCRVJq45N9OPney4WNGb32PxEYV3j0wqferN4ocKS7rzh
JWYCE6cSkmEOV0IGBRJ7x1q+3eqNtKX3/dRZip+bhEQc+dg6Siet1JpDFyRNud+rZ2DEvctML7kC
5qhGZBq+ht7wcuEL+fot4monn80V1bWj7A2BndeL9IdGdviXfS+5zhDne9hz9/0dUmlUlS+Ov5Mg
XUmbG0RYfGI+uTwc8ib+MBmxKHO4ObbiLC45Hg79Cd9fDXaLoyIwi8L+O1DYaATE1FdrZVJNg7+E
BzATeA2XcJkFKMkjd7/CLR+jyGb0yQ613+OTQM3N9XHVQbOXvjcXrfPMu1qeuPr1pCAxVs39+3PB
zGCpMiILDqQQqD5EFtcQjGM6Z+Z2B+MHIO/mVehW9KyrpNj8xNm7nnpDxHivI3MBfvy5Bn7uxeQG
HBbddVTEJpKB/iL8qqRDcTHc73Nvbo9uItGFJoXKkOnH08q7npjPE9iEUvHCahNnvkLI3KwWeZFi
Gu2hGNuyEK6U8N9G7XlrgWHZkLYroGACyPLr+EEGwZhTNb5vdgaR5U6pwT34B+OLxY8ANe0JA6BN
4EXXzqcjvJ5vaDMwvTRmIM++VXNmdkGb7iA2IU3t0rudAzYgEZDwwrSxBIGBnNjFyhhcjJmFM7RB
eFIOAtNzkENkTcbUtasQm5xJIP+9nLTdxTm3vPb1rSrADxyB4ooIAhHhWmzxlym/cWbevRWje92R
bZf0UzRO2OjGPWLfaEJ4X3XeEAQQc+thBLDtToKvVz58aH4g/VD4cHXpZeuXlIr0sdJj03c9zpKt
+qqFKuOn4WZJJnhF09Sq9xeVkVpME12QnsQWF3Q+ZIsRUyGzJdfa81UAq7Z6fz2uYToTgJcrVtvU
phu7EKiLzxVjYum3XLfDC/aQiF8ueLtU7oH2xLr415qiA7HkVsM6UVLC58yxkO6SvAzmyzJwSd/D
yp7hSdPit2XLYXhj0fVgptRVa94T9YfphUAdac4AGas0FvUA8h1mgar+t72kb4bsLVp8/daYJK4P
xt9b6rZTRwOYJUtphIm2LdWCaKuSHxuhB0jPAwU28A91MYjVDa8fDOQNeiCsHwVDUdYrCt3KKNJB
olNCmC4xUMbmbbCOtP8iV3xIOWCdlX7yH4zXWsfQ1lgsC6WseKETGTBV8rfzjrjhr3LelzNG4o8t
BSEVFLFKMEx5/bmV/qq8LltE17Ts+cGtwy+/EcWDRqvKKYnZss0MQk0pYjwo+N+gGejHwoIEXVWf
6ytC/jirFt7U9CioCYGg2lCQ70gecKQWx+WpvngPc/HEeD0vaVhRPACt0hbTfVYyq8+eqkmDkG4B
p8iTu0wYOm+vaxwp4TISzZLPL9mGCTusvwoYhSBkYsFmC6S69pEI8mxzMzD6ozkYnlIwUInyC9wl
A20kwFhU52ENiu4VnW2KviPg7Pe5tJ/5vJJEfsJotX9gNx+l4g/8AwtwQOgRt2AVw+8qD5YRPfW6
vS4cvbXhvs7JHM1ssWHPqJd+NUy8FYLpSyOJBjAM9OtawD4vr39QYFWnzwACia2kFjVRDdNlHId3
wcUjgPpw4hWchztZWcHi0QoCefbPS1tXLsK9CsqbQ+Robj5uWYCm5loM62ursHPiuwlpGdFEAfOJ
BVCjhAkc/SJTcFLPEB7uHF/CJYlRD3Ma5ymuGNZ0YbsvB4hUuWhbH5/OLHNOmLLzXdJj3e8wiV1x
mWl8EMDM7sNl6KsuCkIDK7v7QaUNWiz3lt62lpjCsol8B8WIpzQH0NZ9RRSE5T2Hq7/nY4UJukYT
QU6BKRfb+e2sfl3OWUVMiTcuwSI2P3+Ss05XL8dYe1DUCnj6fG1FBbSQzJtemBOikjrLOQvAOGaY
0latZxwe86qZmoWvFt6Xa8cyT+0skLmzizu5Zefat5vITNErDVpV1Dz6Mtrlw42TIN0/Y29S4sg5
uascyNNHpYaHhRcIhslm0Ld8oB2DjDPGDCsuEilSkVnMtFHjbxzdsQe9cP7E2HK2SqAABfN+rGBU
0MQyODiqf7OFshfenB3jjgOp3ORPNgeou+fIv9yTU244LkpBKkfgIUbeP1oO5Dgl7X3mmQNRMVZV
GXmR3XD65fTdeREeQWRmm+JQOpOOY9TAv1CRP2CqpAAJ8v5zWZiHWjBRBQTbnJGCWp/BL9ASmVzY
4RVcj83y19vR/3NVR+fde5iW02IaeB1Iws45tublFStFXOBYmhnmNTMNLF/B4uY1PpAQFhuGwTMC
d+fTrpBwEDx08z0f33v6vDLfwJddftvIsX7VL8SoRgrQ9w8SoNS5nN07JRyuIB3+hMEO/rfORH5h
hLJcWSOrFHWVVmTVhQzPdyW6vOpR/hMI/86IlUjozcZI+JbBw4mc8gd8qF5Bz+ZG1i8PBql9Y+kG
P//3h+/0ASmK4H5vAJv7gR0haboovURtJ0ab6OhfVMdPcHy2wMHnpfwb4nht/L1YG9Rh5ahGhWoB
rdASjmRDuAC5C5Dt+OoY18C/p8vwF8WUJa/OmkpiQzbg+NZXQayEHJ07DnzLIWv467CEv4rTAZ1N
qt3pCH8QBd5+ryih/WDNvFEcRPeNXtTLE5WQuANObEzfzorbLmr2hoShtVYjheqH6KLe+Dzivo4Q
/alPqAFdZdhQkxstFaT6GG+6mPgL8ecEllhj3so6qrVa++yOf8ebgiD6AvWgfQ+0PIM8eNiDL/na
bK9A1x3Mw7toRDkhQ078r9+/Z5MQii47FRn4USzV6zxhxm1WU/Qpjt4N6FWacPP8jLIRgH8O7hoU
U3SnscK/B80EBvHsiuKSOlIS1LP4KFlexq6cNVX+Eh/eultAfexJ5AovvkTjghweWtfBmIsiqUZm
cSd+aJ/rWcxZhxERfGJ0SpI0/IaG7EgeVKGzmkI9nx24QoXQzrcxRXyQT18tVQYMSWv6lv+J8erT
E79gwZSVVYticUPx99PwZxRr1EK8VxowhmNzY7nBI/41BzmDlyJ+/GM5UhdU2BS7fw80tpkDi/dP
JCSa/lnKj2Ag/okBxuW845pVPkxDq1AxlakEZmXulhctRYSsO7CWV5mTYk2GVp5PNBm8NMplp5pc
gnY6P/6CUx/QPo5JEharvoMpjsqIIpYS4wGo0wk7D5ZybQLneQ/DbvlOj84VT4WZnqKXwsr9zm+r
rqRbLWxASbkFcM2UaN0RB2yqnxzQU/3hGHplkyMlLvB3G2xH7x0Cvd/248qMSEwROUmZ59ah+/7x
ZSrsTXKQoKJAbJJWiXFs0Ucv8uwAN4MWtqQiiCzp9mjr0PnI4Hn6NFenlbKA1oC2226xRBRlo/0F
Nbscx1/7GuuO74RY7BI3tvPjGh7OgT0nQWdrl3IqcKuY+yn2MmfMXNTakrrCPtGuRGkcZhqZybIL
fxNtF8QX862adoxy+I9PbCi7PQeyOKwhdWw5T3wSegdkiidsVu1MmiQIMA+Gxcs0CfMEOJJ3gL4W
uMRnSDIS3WEkvXgb46Ok8xMYG7kVqJjxWWJlClQxbjpKQQKWQkbnJmcnDx8KZaStApoXSR+9r3lk
BdFkjNYm3pd16ySCx4e/d9DYsFzCJUhNW6GIfh+UyDso1MOgiFzKJxME+1+awIcbo9+8QGVMEhEO
JHTS80Q88y6LtwkeUOKPCcMbtUe1Ocr6g4xcOv+A3hYSsiSUHhogPp6SXb9wFghELmXYMdQUgMnP
xlwuNdvrSIxoIHYzbGvvIfPOsLWIwqs9EEEBfJfBD3OL2MNwKqx04xUCQMQuY90oxf19ljL/u+Fm
CZ9Gxw7yB768/xYzKv8wDcvUVOMmE+hg9035766Dz12n5mFR6vFwoyxVj4tk4j+Pca2998uMjvud
1ElBXbaHOCTHyl9lv34q0rXYTobJtPCK9Y/STzhBx1JUpPzeRXgR4+jej7stiDUsGuQYStvvA6ty
+xVMkUlByQUORvV6Q0pSwCmSnd5ezErvtf/ZB/opG8cOXSfpmXUCrLgDNzSfhrf2Au4/tdEl0En3
JVSlYuVwecNkA/BFVQ5v0yifzSdPQlN8/mA6rR2hXj2E6MzShRShHvLg9LZuRJ4HirCvUHavCg8p
nxZbjTRS4iPAyARyLR+77DKKAk8LNbuEQV6RLiMUeHlbEhjwJA5H5D1Y5dewTvkf4TZT5ugeIvcJ
2/2dcUEFwpcc2p+Yux5spnubPzzvrX8X1AUQ6FFXuGfdcbLaCIGPmpnl6Wzv1vyvC7pFOCH4Y5go
66Kn4iDywlUjNvyPr1+tJ2SoWzFNO3yD3nGHXnkyaoxuJL3ZmiLhrdi/Skkk4sD6ffmGtXlYsr1Y
rQGoYuUbVPHsDqTa+CnpAiKkyzlM9oM7TdPMUiQnEKJpkCDGNOsYZcbCmJP2YwSijh+TllcZx2e7
2Cf8CrC8cCb2loeKWusjv+/YjRisBtBJ0G12pLelCz2Ll8bfCfd9rnQHPDiUDZ+LbKYfO+KdlPmC
pZJZ10F2V5WvEDfRK5kAv3A15tamX5ssyEFknBDr281xJNsTUXPtL9CbPDcFPburb4RLn2KwlA+I
cxCUMR4iFfFgbcFIHq4ZbEK4xc4mkzx9uqSU/AtgHvCrXLGqrnybrOewss89FXjfPQOmrJqKX9oU
7Z44qp5/kLpakhdkIBsRjzWUwYymnC6mG6EIdZ0zM9G63CMV4oW5ToIyJzvfOT510ArHqRLnpZqt
/HT8lHkF6zUKbglZyNNa/GVO9esqijXuQ6QzZzjjtWLP+bvrU/XeACbFnBLC8pLqyisTP7H8TQo1
6R3+i9izU2RbURjTDU5FAO9oCfMLBCIjMQqNSP0v7A2SYDxsifjVP9rnP/4AqEXpH4dJAcLJiZnl
C6sunaiHn6xzA4XZfaHN0Lq16eXLOTTGtbt271YP8umsueOm9t3k7MiMRGpw9+b3vZs174xU3sYt
8smt4Gl9AxVbg0zm2IIl33QNAHqjGcxz4xUaJ+a/rQl1fzaQZqj3wrAYVv7LhHFL0EwyYFHbOSTK
EkmM2+xLVN/iIJdwJiK4Rd8lFReT8mb6UNXDiwkZw3whWCPLB1CX+s7wlxFaxsGApUjqAKvZTQNf
e5+/u+rlOIFhXnDnV+waalmeG8qkUTyIKGrwhoBeyesryCb6HbfC1zVXTUc0bJqPTDBvji/6LRDy
LUm9qZWUTDmmFPaXtAcdQPAZ9CN2j/tdNx8DCzqkw7PDtfpMfTqD8imxqD6uOotd0YklLSF7VRTS
xIkMeQAjYcu8UQAvJWc1UKioKAy4HO9jPQa+okG9WV/WYbdWHPgeBZNHW1xfn7A/jokbTQ7YUCZp
eG5hjEMWxov6Vnxj/+fWxWCaxsU4h7+RLQ/jnof/EPi798nIMDp8IVoIKhwz9e9alYS0xSugDQ6M
0hMvG4RWTwPmAorWgk7dd+YohksrjgoTEwyNONPXqW+99o1xmWWPCM/BXcHg7ooZ0zHmFVzUwAbp
QwBQ9dyueA/iG2kMWEUV4lx3BSdQgpa8NLjgppJGW24LVDPEcL/g72n7w5h4pGLYlOP99KUt9sBK
oIYgoBlOIIOTx1KrduOi+VLXC8zpSAx20DmR4ZMmmzsWOe6u7x7oec5aT+SyAToR1oETX/RYbFj7
61nBK8L1BCKjaiDlZzN4nH5sCrz2TG1OKc6b6Dq8LXX098+vckt2mDIm77ExQn7iLp+r9kl67AvS
pwQ00ulkjA0f3N5Mdc0D8xNaxEncxu+uV6uHBquc6UdeMq+b4CFH9jKu4cnabx3eVyGctv3nS5bK
WoyzrNltj/ldTRMhuAY6SDYNbAC2oaayJ9y1nkcUsw88rNoAZhp0Wsp4Z58oAqvQCVdG3V5fSqRN
Il1S9EOPY9cSQjp3rDtHhRW5p3c5c55OuIBKH/de8p+mrnyztt/6HtpXM3pMx7mh0D0p+5/5oku5
SoRztdfikRRxfDt5OWkBbLmVKYM3um2W9qLrDioNUC+bwUCssn9uxQyB+vE/UAH80pId1ODYR9Ra
WfDLrxnr97ta+RqSCHQF9ahiiW7Uj2GQ63ONTUfmlk1oRe3Zy4RHPtzNdQT2z+yFbTAKHE9p9NYL
PxR0nGto0OPBJblI6nMgiT8Sm1E6+1jJTtW/jVedK283TVM44WGdhFQQ7np4seblw9Yexw1Ft7PJ
KGu9/+VxYHeLcpuNknk1cv5mt4rJQFELMvhnzYyANO0uJSQpKpUXcpgVQ3QsWZaVMO37RZ+F76rf
bWF+2XmC3KWEtbFx+Q9pfzEm47qJENNX9+pQ6IzjmFpf40hs7z4ThBJK+WEbYSzdTV9jb01H+psY
PaFpcZWWd0VGf2KxEHDd6fL5jN57RKGFu/V8znJzlUV1Bp3cwG0TdVYF/cxq6dbCrm9Izr3V+1ux
nblocz3UurQrVuz8mAV4wAhDBFgstrjb0J3ThWWVSDrvW4/L6XxUucOjYL0ESQW7udGp5brP04R+
/W3aNptRF1JmIZ7r9NtT7tg60+f9rrtl7MpT2DSgARsI8yEi56IhATlLbCr2ogh3sd6X+I0uhi1l
kytLorp75PVw2gqjfZeY4itAfPilqKcg/3Q/hw42yjmXPf23mNxt+AXyOBXzaaIrUwEYhat4y81q
6AlfNh+juIFeDzAnXAo2WekoQ+D58SOOhVR6Elh+d0SSo+acI0EIg62wurk9C4esWjPR9leIPk3m
aiLDDlbnIkoqBFlHMZ4FX3khtLdMC9Grt9KD0bzm40XiHex1I91EoYTtOFrlq5t4/Oj/fIM/s/0M
Vzx7YLz5RF0a/eG9Yski0g5Lw3n7H82GXSiAqRa8wOP+dQEt0Um6PhEGKJ2v2T0MwM1qCBagyiKF
JCoTGb4OvZr7X5+K3l7ETFH24V6JN6tqYWnzda6x+3gBVqQp9bXEB1IBavFVSbh2VlEUtAsrHby6
N89chm7mmWiPSaBLF7kzfGMonFBRkD8o3lBrs/kJ3+acMgT+6kJDIhOo5+lPG20Btav4rj3sL0Gt
5iHO898jiL3ai7EPh4UGCdhn9XcCJYzynMX3Gq05Y1GNlo8eciZ7A2cfJyYZeItiQ4hY99kbC9q8
OAw+FQmchx4dJwnR9xyzIK5ACzmqRt5j+m8dpyq4q92b/zJE50Ht1tM3NdH6XQKlUYgnUKOnZVLy
U0WaxjBee+EzeoiliGP2PQr3kTa7nhmQnnHRihbIruK1Ch3l4rG1Kok3bPQEwMNMlVrE/Ym5ggWY
RnOCPr8UU9+MENL2wFiqzopVMPwnQQjTweS4KRBl283n6atunVUqbtZKd8DRKFLJBipPZJaMWvmn
Us1Hgvbx8LBTYmXhJLegr5hOf08hc5lk9oWpxVeywnNa2G6Wl4W5+zr1DZL47lOVEfYc+G13Ilke
j5TJCAK6352Wl/4uldbsN20Bf5egcUWWkmx5VNib8nnY0ovHgTvT4rDZTdKMiCOiyUCLjngUGqA4
WlFIUhH0Q21Q3lzMCuY5rk/2qMu+NoSaHK314n0uR+4iMVd/ghVwPTxn7WbNdhOF13k119CrjGll
gcwHO06HEIP/OyvK5CQju6ekmMVu8oVlov7i/Ri8OlP5lATxji83b40OQiOeh3s1owMAZdB+ilNO
KnJlfk6NYMbhCmi1RqRcSbTh+Z3NAvf2BZn7DfTW6FPuAzh1t6uxix99PXKxPec8NoEhOjt/d1cE
AZdR5qYkrlaPQVhmA3xSPhoswy3kZ16e/4NZZPOh8vMxGlJwfoWpPVP9QYhkmXIfXAuUMCImN780
PTjWF7lYx5r3XYQ12XuuM5wF7+7CWGns/DDRWic1Ik4Ht4NhNhlm90OHchxdumNsEiKFPg7S/g98
TZr1setzZwrdwdj1Jfe+oV+kop1G3miH6hWBMIb+t6utV5y/VQhofMXn3Qh2Ar+/49uJ337a/cyC
y4Nim17IReZDl8YotZ99oHn3Gg8OEgAQ9/wSo73G2Nxhmi+Y3tIYm4yrA0AFaHrOmQoPWBUAUnNs
I0GdCGacoDthkS7953rPw9iVj/ETym16zFj+vMUvhfDuqqmqUskjEjt0nxkGKiYH0L/IeDqDr49x
aPclvNhSdRsjK494re2f5JMFuZ6AxVYb3Aal0ikbVDxZdxhjARW4t7LkJnPm9yiu3nKM3t3DQEu+
ra5farjj9SpooyTas0G9zHm9QoIHX0oPPz3F3jf4aNzXrL/y9gSbfV++Qd6Z78KB8VBZmN/GzDb6
XkcjQkUJqbhty2gr1izHNXI20sOxKsuNO5/CgyHAmVzloD3bxoABC0Oe9lAsDXFyMBjlL152Zh+8
36o/HPFVPcx40VhgIATSy/Sk8sogQxaL69puX0xHLcOcA6rfszYEe8CETypxyjYo4oJuYcGkoB+y
1OXZGFaJL/QghqT+8d8rQclQ5eeYejVxTqmElU2vgyURjFOnmjkE3AA2yX8v5cXFbhY9MlvV72tn
J7D7SA6lMz816krnFhX8UQcU0hzpL7D9LA9+oc6usfy30KkjCMyD12qZ1ZocR9l+1URP3mqa8vfU
lM+hpnq9UoYAf8u49bSt/KYlFS34v0soWuJrCs9k6oUnWaHxrMBU3CMC7dqiiOc7+DDodusFyvnm
ytgK946AGTDYq+IHda3vwy5QLgoNmCn+36d8XUBZO1xPF6bdgwq+A9p1ySkHmKmTg7tYl61SKXZh
XtDeEWYqWh+Wc/2kHQtlcrjy1WNhTyTQo1DBuxy6xHxBqZH7YJnxfIekQwpDG2yzumvFbVfCno9U
y60d+vSiJL5+A/b358JA0eUohhEpelnfUtiwGEJ+chuY2zkE409L3+GJSEdfiMPBI0SLrwNc6F8Z
PJvDanyAQkAZPHeC8UaMUGeCVEsbnNTRDaRxie7uwxWUvEOab1KRyiXU841sEZOyVKzoYik1yjZU
MH74OoqdAXfKRDT60C0Zi9vfNojaNzM0wk8cQuaXgEzEfvkVqhPDZ0Thnhg8jxdg/Nkuri0XCROj
ckvRLZcwiErnX6GO9D1NbJu02q2gW3EeAUGY3OfKsBaRSInCaVoz5l3vNPx5Hv+tqGDtNUMdU1xK
lypViO1cQ4sJ8bgauXx4l/SK2iggqr1S5JBfh3NPeCnR3Wz/Omru2kfk2ongUUAOjLTGoUzwVOvi
ZrMRkPsSucArCvpoIx+jTMU93Ph6s14P9PlJOEShIleClGYHADMkYHAM/Im7rir16Bu8B0ftkGdF
1LmlQ/+rDAm+iHBwGgXzDURHdhGMIPXF+7Nm6ChNP9hp3Gt/IK/MhqKq68vaMCiSk4CFSRc1QNYi
cf1DbsrEqjYmu6DMSQTxkSLEXLguqLzKiHwxqqSqfPak1AYXdHO5jHyKFk53013MX/b9fP3Vhmd1
r0h3u7peF0ptcMCha3QUY/oSd+SEy4TNDDnTwqyB8E+Swzmqd3TukIW1i/FvDCuh7YMkhYdBjwHA
hs/qaxTN7y3ZIgrYYABMk2p1GWUgJrXHd8CuoA9XDXABD8YlZStLiVqwSrvfwSn1roIZh6eDnpJP
pOHbb5rJc1bsOWyS6OtuwutziNndHTuzjxsiHalLLDLrLuntOoPTMH/RG85dpR8Rd0QtTl0ZkbCN
foSIJM2l9CmqQdv1DMp+HN+V4oPUxlpVBj30bEZNL+OhLw4BY0kwlnJU1O2yomgi+66lK4o/pSXb
YU3zgkVAGI2CU64FFdRZgyL4UrixeZSBmrlpiRPPJJH1hh9fdwUOspvYlaR5W3PtJT9RxRb0HI0i
ptb8gyjftwo6l7l6Uv1fgfbtcidNhHGfr0sOX50O7pKgdGSjgrmTokrySnMmEPPv+QwLRihbns21
M6gE/uoS0FtC9kKt+BObg1BfAAJ/YOua+qTmahd3NVLJW27jxqPr73pkSTwhQw2MPYdTL1YeaAg+
0grMNiwP8Sqa4LgtSSN64nejJwE+AgY8Bc/ktZYzJsZ0BsTNu1TSonM3wT9OQ7Gn1mppLoDzTwJm
+0d3iFXOWWq4QLDd9BLXXvMVv4OKdAMvbweyc5VKdRODXld9r5bfmVRJxwmpMI5UndyisswCB4t1
Gmvu1YY6htxTkV3hTZIpoNysvfG8aTEe2RMkGzbB3ydgp/d+o1Hq4x6HclLypIqr29A+8llBFNkJ
MasHDBmvZu3kMHuGLRrVGFbkKOLO+n+cJG0oNl6mIbk28aXHpRTSrwBFJgO7PIdKzfnwbwZ69yjg
Ib8+t8iDwjKfBBPuOxT8k35Ipiwk30EYQDqwmzauzzWTd2xT2ZQiY1ZUOvsbCypL7UOqRAtZW4QQ
BrE6Y+E4T17Hstw5syNLZbHlrTn0aCjoAxYwxL0iB3CmXm7+MMpmNCeeUkAP4wvGaVCJq1asXdkH
T61tlVNgdRgUdMOMh8wVn90LqAyKuGUN+2+s2u2RGvsYyf9rQeDf71cfwIaP2SGznMlwRIegPXaI
KxCJ+AYKIgXB9aJdmXYQe9ke/lmb5dOn7qqumal7vU9msSSUTtws4h5pk+2GHlto+Aj7vzX1hr67
CAlBjRzqleznRlmkdnyLLdjCer0VdZm1WsX1wJhwhKdMWE5uijaKBnlAjirgSqEJ9kfiJVO4TuH6
T9Zf3micyjRtduQJnn/x3stddwZ3VoyYsDVavUGUgRLSEKTDR/K5O9OkH6z5QosC0gibfnwn16M9
CoP/EgwSpa4exchSxQ2ENxjgkXoNSm3PRAmA3z8qoaKIWeHbig4ChDdAsQxMCUbx5cjePPXHRZDZ
2l92x1v5OFCJJWenIRe9F5g5PgZb+QdAWBrzM3/9eGK5d4hEavOtapP78KnEUFj4AEdUBIsPWBAB
6KWNjccqlfbhjnXA3jGFAPjbaG/GkaNTlRe/UDM3BWJNGcfycdiqG1dpIByTjHqVUBVq5hs4td+6
ua7ECd9NKzAavvfBVReuxzxnHxnaJKz2YQb4SA45b0aDgde178Ab+Y57KuBXXW6IaMldfC7BjD3I
IXyDS2l46WYd6hF9hSNbVc6XO6EjrO/VAJxYIDU398cIq4dsA0b+8k+Dby3h1st28I6lElDGWCbe
+c65siQDXNXzzisbEoEixiWX1CRLShSQxcCXaeeT2GiNiiCoeXZ4/vP1RJlsEGVN4AQnLzaCZs+h
dGecrRvu1f3pEmesuACK5At/ElOHO51hUfqkiLHokZKzSdoPMQsVEeAmiaR2frZHwGm8S1KXrqRq
RQV+QdKl2fYzHwShRKLhb+3ez2UHkDdWeL6rLBfZDqYaj8yvnSIevXqqn37yVDXa1gkWJwJGMK5z
gtOm4v+BPTzFq6uSPwYXfwjy4BJ21sTxYR4joW/9VddH2AFCBkjjtSPCYmzpEGlsIVXgugDxhfX2
qJK0tRFRznM7zIGeilySF2FZQNnJU6Lz7vzn3RRqjipn/Shi64zkFT9+VYWJKsU6zrnf5Pg5Lo0c
Q/dlDj6TyLbnRbD646IO7b1VI8vVJQXgJaN0PsJJwRaEZw37eppHZvc9LuAHtiV9y2+fJr9Qf6WH
sWJEHk2DOTAAK/KPo3mpNx3Lhg1qvXdma4SclZWWC8fYDLs6UsRer5hsQSpH66DG4LJI9hJCC4jW
IpAuZyo5HhXasZ8NBl/sZvYL0mc+I7qYsyH0hkxzTDVPLXavVjaoa2HFx+Gkclf1WiS4ieVBtZHW
b4IVZynFEOIIlYpRdMXaCruXQRsEtB5eABUIkNpOKakdhNiYAokknBjzHem/YTOnXatyeEU7n4Au
T4kXeLUho3xRVhXYgipM8WMoh1XAs1eIA8obz1mmwH9RCY4cqhPmt9A2btBL7gHQsxsw0xYrHS6+
q6teQkmAKvyFVhskbxyyADvyep9wdLJwyl3pR0IbB9xiwcv+Gy7CJ6O4f6iJHBuW6dRoKJrvw7vV
COjldLbmQ0X9IKMiJnS5DFGPei3USvnXlPElGdyBZv0staiQbasvctwnceQycFtQfUD3m8GoJZIG
XfMuutbniTAQFI/7gTItrURN63+2jXkUhc52hRPR/x+5jWa1UJ6HXICa/l5PHkz1Rk6r+rGCM8e/
o/5EQnTpeqQt22wcp2yMEXoSyBZzv3ly2VFEKS1PJxrA8wCxEWmEYtkYEid19nnJxmXUPChOG3Td
93qWcBRv73Xjsa2+h8gYbphzdNwZUnshVOu36tnQXCn8mfNlLAm+5+MbH/UkLJDp1XwDFl1E1k8h
dp8/32V3zDYgaWkix3kYSX1eOihOe+ECtuAkfHZUGmZkkuwZX6ukgO32wybKxr6aDWlutZhWpvtt
A+OgODerRjUaKo83UgarfLT+og9nd2jbTwOF31AhrYvA8oFMX5XT5IwXCzzTFcHVZoxShRoDyhwK
jaImWfHSQNJRAiYfIsu2KOy5/3P1RQaQtWgTST4GQLK2LAITY/nseDC6XBZtf4la/p9t8Y/ymsV+
qnsVe4TEykTy70Bq6baBT7LGx8r9EgvEfWOYabE71Pk8UkQTHDBFJZR3cneg5uqmdL2vhCTP8C80
Hkamw59ia1k2TS+fewSuFYMgWpqmUIV3K/943qkWjWu0670c+VXXLaYkYlTkNesCxeHspbcgMWUH
LnnF9+B+g3cJpY/ecg9c+wMfY2jm56UfUm8zFy95GlJ1cLwDB83TiPdJ18XrmbonlLfwL+JBXKH9
SpiJC7TdI3O7B6MzSecwzVIXyg4iTjwIjvk5HnqukdPu0aXPyyTopk4X3TXWD0ekLsyzBNa7DqPZ
LhnVm2OthmYAJokSWdvqmg0Eouk13WVWjJJjSTJj5WOe5/afpy3ABlM55GPNlQK2Q+4OzBlA/F2V
3379FWI0/Z9MRsN9Lt1PHQS3DgbrTNyW5ryfpcNs5ZqWHXXVdi74A3cYddrj/dJDUNEo4iJ1KXTy
b2l3doWEckTyGoNOdXe5wIhDRlaS13x7mHC2wp5xQ73yoYJi7AwbjWe4PTC96+pf3zGAUf93Yxlr
J+Ou02uXaX75qsDYHBWSHSTmmvy/oq4wq1UMiOdRxgbN0TB/dApnBK0QtFA8L8V6K3a+3itSyEiT
hBvcozoW46lv955Pr8TwHs2ywroNV2RlwoDxo7YmFDX4rd88OeZaOJL5A4sP3og9bD7DDsjoDfUt
hh1qFnSCxcVUfGdRJwFgnr/eq/P1QOhaBEyTV14CGEUuEGLaoJ5BSS9Qfi2pmqC5rMiBJQVMxNFi
E2GvKcUtReFM4dGULa85TN61v6YJOGw1btM01QKBx9tXypUPIVLvFQX+Xty5fM+U5LNgDJIHJX8c
sFYyQyzCybrBbthkiyUhLMxyvCOmq5IcBbvTzwzqlL5qWygZ/Ns+ZlvPBtbRrITz3QXoghVLO56J
dWgA2GRrjgLDEMAPX6/oPzB2iWyUNd1evSNJiq9m43C/FPr2Rkvlzb2N98m2kIrQw9hpZhMAA6TG
bPpqBPhbyxZHccLNJ+NBNpcAB+UtjeBdjVXp3rxTLe8IJBORiYiiSLC5XPGswwTtk5kNoiZII0ci
r5I3fVvQYWfVXFBucCCLLcGNSvD/Qo5W9k9wGvAAfR1p9HnB5dgVddEP7Re+7brE4Qsi3G13KpjX
zJ0/oJQ+ZbAO4aPhSzQkIOnVhluS9DRztjfDk8wOJO5z4KfYyhPe8Wgk9mxIpbsrJf6Okkd7mQ5P
hYqULxSwA6aO6WH7H9DTVAe6LLxyhtjzpIyoFEmZvkccNYo5sCQPqVUVen4n9VA81QVqkp44dlgK
SbBHsWIq6v8x5zddZTX/aNfkhGKbIqmHurD6YgO9ZvgZkD+W7/6t9qVuUez1bWBL0UD+9MyTzziZ
dFYJ2fK6CuMhzuAUJBDhjvRNENM6YZl8Qx2NGoq7ajMEADZ8ArDkk9RvDOjW2qicyg7i1lyaK7Wc
ZfB3zr387mh2euuJeGFH27mWz0TuojjlwARK32bp+ir5VUF7HOZT5DliIJKNsHgI6escMqzkS/xU
5dfnk6fhnM1viaD8/R+8y6Iw7q89utYMSGmK2DuAfPNLQ10JQxav0HPdP0XNmHa9REGQLRBGcpfI
fKWLWmIyfx6YkSqIYS350EGcA7fe+Q7wvcZAfHr8zxcnYUo0xjJMpNb36e3sDwYlvq7clcN1OyTb
h4moIPKNFb73XHsjyBWh6m8nNq84YjiIIFjNHeUKVbyCDOlNGWFqIhEqYh6qJbp90HSEVveJyYXW
CVdE2b8j67UGQ2+vsKkWZER065mYX0sKeb/q985SjR0YA9NwuPW5v4ZitJh4fXBh23rf/wTKU8zI
7yOdkDzmIeo1Jw5RB4tEqu5bO9upFeF6H+jLTSa1CypSHZpI4B6MyfdWrzIB5HHYSxfEvS6qlXf8
nACqvkyy9dRApv+dw2obqpk2jFUUb4jWfM8RBYg4ZA/NmRFRnRQOuGFTOQ8VheqYqm6tBjU9/PcF
+sC5QAQbtTkSm5+pYg18ccjZPE8bhAkAi4A94fjMPYXsZvf/vYNZezvhgzgoQIx8UvDDxiB335Xy
7plQR4Wd7lVX6mOtJqB3h6ZDgHAXZVCOFvC2vEcJu1RaOCs1ZB7y8JPGjRRBV3ULsTThBNhG+viW
1+31Q5GBXx5nD3gbGf8jW9rAzF98+b1iwW5op1+3MffDW+rAZnBzBqkNj7yk45jSB7uwGdP/lCIh
/6lWbh9r1g5ewjZljqC6eAF2QhsFL9NKXqb0eAmUI81K75Jov+48eDezz1B590NFKA+f9DypX0R+
UjRNWO1vaOh91GQjqi0IN5IxU8aIy64iW2PuwesVNy2BV6wILf5MsCyGbzTNACCP0Tli354JlqSq
sYwEMkqKxBgGNMhqp8hlLygzQHDed/Bb0Tg9f+VAP+eQQ0F4C6lfhXQim2+M3zQ/HWNvrnVm/k8x
PLVjp19s+sSArGklMAfY5RTorpRyaIvuyQzgoty9Wrb9W7qfqxTuv3rzF6RxToOOPaLFjEzGNQPN
NvSPUS+cKgtNWSnpiahIAM+9ecnwwYZgyYOlIg8IAhkVCjcBUYsr9zZKYbGqJy1xAqYLQU5hwnqH
mrXO03i+Ij/JKE62T7kgJyjK4U5uf2Gato5yxPe42snULgIZE6eG0LPIh8ZNc2LDHaKnfMgfrrqT
5CtjGGLgDcLfPcNQelswW3ewPZwydVl96D6e26F4yHqbh4g/71dk/psrlQ1Xcl2dOWEoayt7DK4X
MER0sJ2sXK1PG1dNPA0bDas/tRAQebMIc++VpNckx8sCv2ptixfsipBJW5vjix8i1hX2e11kKoes
IZKK5STFOxviiT8/aL9ZOwmsvt2wZhRkcVWwFMyIRIB2V3ttAeZ3T4kDF9wEYgglGtFA842oxkAn
DOi44tAMtBoM/YorEclfy9NE5anwNDPd3IyWHiKMyrE+GYNytlguIMwZYbhFNjU5FIUSBe7tyzry
EVNoM3MiExDGspqpnAB2mSKQYy04xOUoXnWAnvcYf8OxwMkjODEjEZySO8rJ+5XoS+ZSgtmBAX6I
wl+Ea/880F2ftxMwsiMGpdmNB7Y0Mdq43Y0ERh6TQ5Lq/yhcLu1Rc9g2i/WRIfjhXvclNAg0gQBu
n8Ur1Fle1zO6HXhU4E3eO8bUjM9GMb5riOjWIlTPqNWIdCpNwjztbT2HS9LKsOWKrwNRMtZVMv/2
iFuLZk7Nwu+73euQy3PM2r9niSpGUZjBSd2FC5fDiBWV7QrIjV/hPZs7LpPQqjYdlCVoCBHJxIE0
AvnRCDG3EAsKZL6gwwdg2Nu0V2naRYrrHe8ZhMXO4Ldx+eNJ7KVE5WHt/8Zhe4sRQhEh/Y9Odlx6
yylBg+owLf1VLyC49DsegWUCrdrw9KD0HhFsABnZ9IU4wAymuAwh49g/3lnjWClqZra99wMsVIEE
4xI3tEfExxyNjRZwuW9bwp4VopSD63SIjNfLBbLgj7kp9BifPfLBe2saiWuLTF/CthF+h0Hmqufx
3tq3UDWqs2q3IsGzAvdNJWofMtbFW2nfpFxPDiQT77OzKxVWbKWgxmCxBcSDy5yWyZRngXKyWIo6
GpWWXZRuxWoDkkMNlm0OjzGwxIidn4jtj/3cseEM5eitM7uPDVP0wxarLC/IUDsoUiFIfRmM5AS8
ZOR/zZfb8j56W6X9Vwz/N6XrrGR/9WBIqfCPBCBoCTynQAgx53UsYqMrHhgWEdYj7noKi9WBaDJI
GAEo4URRnA9jpllddSyMzMXfE70PBS9BtAJ7aTh8LPRs641RF3ieiF1rfDZDcjLk+6NiPJbbEZXK
6iedeC37DkVOmOBH6TVN0t8/RxJRcNh0f6BuYKBEXv3XbCDCi8YOOGc7l4HOmYjc/ULD4nwz8V/b
8kkOxn3HtYOR3hL719LH0ryN9yyIsI8p5lJFZPaqzzWua/AQx5kxFw98SkbUUEXRfJU5g39N31kw
nElsg5WIUHpwPXjf+/fVfenWdd6bse4DmDzj7Pb6O7Zzjpxe5wVgOm873JEBK2xU4GsMIzA6avO+
XtHMhCJQz3GUTszjM+0fKsrYzDq6gGZvKWfDtIaIzLTZmxhYD6yn/hBOrBo+ADuChZUmRto3hLtV
LfIvIjvQbHVQIXEMTXHXloGFulHPRZCcXoafElOhzAzA7GzqHeYxk6U4orJVJOyOqv3up+TeN4S2
yNMzSHCzH3xCtUkg5mIaM+005jDHySNDiC91+dz9lqZ4frVd9Cn4Jh9+Ulhf6zzDlCrz6MRGcqsA
lmAGMM7Tg03NWUAIAvk47aSGdm1H2dpAh/v6L9tZM54IJqtQuFMbIU13YZHBkn7/0vckaUU4mJft
NDJVuvpDWxxOdQwBhnaipZoTAfCxSbC3u77LE54FwDFeh/Nrup5/FRXQVw8CqfiAH8xTnLKYDGRQ
bWUum8Jv3YXZgF105qbr8X9oRJQlB+OZJoh2PqBvbZ464ac/rQxxnz3xAQzF8to6ALFyuRWvP1Ia
ykwMaY4Krfz/C2F0Yp1pGNbTB3rphasIxdQLtoSTs5Cp/Aaj0+5YVLc/bclvuI623Qy4OrpmhNRM
JF8Fiixb2UbiJpLJuqb8juB4uH/y8t4oU09OHR/MhtQNFH5lRM1rZsIXEHJZzCrS+XvSH12F3XcW
/Bu80hRnHXJ9F+3HI2LhH5xUe15pR1zxo0x1Mwkeb97cnwdVMIN9jPKL51S6GqxxUCMNfSBRHgaC
ZkRWKVT/n7V1B2g9pA4VdGXs75cmREjC9016h9boQ4ZTm0OicWDoSUGIPJbOyui1kk7ZOwARJ2yM
wMj07oNTKnLUvhr/JJj/MK4fX37hTw5Bav3xfdSNvrMtncBQLqvuaXxZhQsJ9ttqs38+dMbQ8IXu
ClFIZ7oTV9horPkrtlg0xN26FIfpz6m+l9DfUBbdFVdVK1DpjAjgZ91C5i9JZMj5m7wZGiakZWD2
ZE51Aln3Pb/xyh9k/M5M5ImPmeBP434+egQ0RwqtH358AiX0i+0RnEZSut8VdMwzr7Nxd7/etShC
Lyorqr542K7cE/mXKZ16WKl/UZQHJSCO1HaXfAT37qfRpHRbJ/Jo5LlguQEprVNhvYVGsKzkGbHG
+0kPQOMz9Zgbx7M8nKmljC8rJ6S0RBX4U72ilpM+TpiAAGMfIMks4aghv2FDgSOsQLAks4DE6hLj
AWicGqw6q+xxyBeetUGyDxxMFd476phRybjoOAAx1/BCsQ1nRhaRWEfYdKUex6DVFz6/gpsfI6PT
NOr03rPd14xQzVCdxOC838weFyo+vyN6r/BTuoLamxrdqlrRTzm/ejHv4rbAbnP9s2592Vi/eOkI
7VbzH0rV+sNINE4YdujT0Aj87uWNvVmE8Ik30M8Ag3n2yLiD8UEOAtTNdQhTJ7GwFP4JjR2jsZUl
6NReX87Z75PlNLxU488MlatCXhFXbldzQkEtJ1OMrj7cyb+z6EQWoUaBNpdENebiTYeFepr0Bvj8
5abuQX5cP89SLrdo+FYXzjns1u7TJuVozWwzbVC9aCazeiIKqs0ZuqBYc7ncVM2McNoGt4j+WEGY
cw2x0lfuJmqpqZjlMdZDD9d7iHkoMYYZ2QJBlkX4I/xobLuIT8quRoVKAn9+hNF3uaMlFIwRMtc4
IA+9PIYXZxFv9DBTAcB9DKM6nZQwZpmjdsbcQ5dpYtD7pdu2j89L7d75YuRrAERObXLRGFdgPmRj
37N4YU58r/afpHGOjbbzGyLPauVGbTaXdNl5uwP78TkvJ+iFDIbZV+K1sVmMRFxQqXNQboqqNjTb
XRj5KNfTeJZaa4taBaxwbqYqOe8hlwUCWW/c0ap+KNKrMjjstqQtMTvONMchNuxB0c9s73MleIst
chnmEylYdFTdOilj0ycCryQGV/5xHRucHGhjRi/WJeWBvS8daAUookBgr7qndz1HaDYyzUzjQkEX
oAyhIUiygloKu9zfNOnYyMxt2/F9Cu1WRlgA66MlfhNGGMnZV3p8I3HIvMcjtNXi/+QWt8EtCQq/
H0XbRzFfkdBoTerKB9j5/muNVR6SYKUd3wC6iQgp2kF98JoySXIcgZOJ4agC0KqIYdp1vKi1/hOT
I87N0ozzS+wLrKgXU85rJUE8EGVGjRbl6/HBqfVy8ieQP8fIezqbRQs3W1bC9CG1DJ+VU5c9yPGg
QDLfnzPE0q44soNhhOwDZRzH3rn1VtuiJPlOhltnzVQiKUIKPId7j28s5oUZMkfWKj0ykbIDkoJx
cdkt5mvwYUUAul+uCS/TBUMxsGQcEyqQqxi7lmBM/7jlqIPPk3kGHODb5GNb1OwvCjyDUht0oDvx
ueAoV8LKnFFc3/4Q5I+A0WwShjdLt5nrZtWCtRcNXdX6X/hWguuyUBdvk/4QFvlMjvSQxcnG0qIj
96fDOh2yYAv4JW2Wwi84P6sR/nrbiUXX4uFfZ45uAr3p7Blh49imqH+pAG/tw7EkZSdOmlHxtsZx
443fCefXCfyXSE2PWWOnhIhI1zZzmEEqe02oBdUStpYdnB6+TylTtu9EFyOpbqarfAiCcaJz540d
PO9YSyu2+h5PsQ3rTFd7eEbKd9kJb9OyKt2nL+3mE1N83nb5nnmEWVA/eTJCL0IeUPLC3VEsm9rz
flDARNkS2npcgbiz8ledFfLSZx3v8aISuyNnr5F6l/+sm7wH43iOexF6uYT3JuZt5gi7mlgtv174
hQaqDEK5D+8osME9EgTmjgrJxDh9tKSXb51jzPBW4JM5HRmJr9SMgbZn4uNDFm1vB73Y3rTH3h0V
H+7P1UX6ZEI3I/PtzCD83yDsnTw2t40Y9P0KS8T+oJe7VQMP2OK2KFKXm74Tu9Idav8c5fWiJy4o
i+oJ5HMHM2/tGp5azQzvjcsmNumXscqiAY+z50G2MWkR/ySlbWPojONXMZ4myT9dF3y8kdGw2QYw
rGO/ZeGi8nxSKGR5cPBDEVMflD4YZl7MQLEfOIyPoW/Jr+LfsSQzbLo30eDNqC28z02nptrdCx8p
5k0BUvuBhi3yeuOKgmLiBCQgx6M7KKMQ2VkhcH/LiK5yX4tz4v/KdPe5f208nJnRbFDUp6zOaMY9
PbBC9NX2i0pYfNCtoI/NtR7L7A395tUKURpiqPf/SRLLwLXKHFA4JUzMSOdl/LF8ORtmQ7zavePw
VMhKylo+1WQgjtabez92iKkOCOvm/5q2y91O/NMg1qD6gNijL6rfUFSZulHlBYKCo/BLXNzY3EeE
yUCQKne9sywFiJdvnSEoTRb3VLoROOyhB6SCmClqDuiTEXTZLGy09Qo9r5f7ioUWN27KKMmUPzLx
H77wAy7oh1qjU7WWQsep8QgKVQF7phGbBpnoIb3UqSYRMoFecMDmgpiNuZUMkLokMobullT32qVq
TRLHQS/YthNvxPK0WH6eQhP5dPCYkAIIzamyHql07WPmvtZFdeG3ahXk2PtKSK4rSFW2TAXXVOiY
uA0CZFWVayyfUjeZ2lDUw60I7DaAZ90RS8pauS7QXg6VooxhgbuORrxMF8BToAMtpI6codhERLJh
GUDXFk3cM8+aHV755/mgbc1UwE3Top2suqpfr7kR9C40CY6Qv+Ln4gy/XqXna+MXhEGBXHppZQtY
r7jHBsIFTBDR0N9KJCcvx96lvVmvRhCux/4+bb8ox+6zfbi7yjGlCfOgFIDtqgY/OYT0RPkVtHVO
OkOlEU3AVox/k5BKk3S3X2hux0RPb6Elc5OApsbMSKWDjNt4rWJT9Q95WPLVMdYK2hWAcH7jl2dE
eqbPFrnrCuMYO0ZD58N5KEo2fZ2kwuPZBK9MU0bNR8Dlb9sfyzQnjML/hVtae/tZvALgnMWBDAVz
i4q9i+ZXrkI0KCX6rQK/M2klI2v1gCOS+JtKmwk3zRVeaW/rdvDvUlL8eE7DlsOLul6s2beatJZ/
GmduG62FJTKnBI0viMt/G6gkHuq3NyII5NSeDpORAZyEhXAydWLuxsMNn2KRV8VhhuAdoHNoIPzJ
ZhVj2+hf6Erxfha3ndmbkmEZMaEIxqq9O+ljeQ8DQgsd5zk5vmCOLunROV+fI3BEMETfYzcsci3i
pLJZKVDoOPYC4aUT5ex2SDsWIcVnPDCXvhztbFUpeBXWLlZWQBEIFVoD4Tg2ABHVAJmpXP3TpRaE
KCRmsqdsqKDSJAIGdREq8BQYFEle/jGXI3YRZ98EAj2VuDJRhx4aYOvfAaVtuQuPwfjQX6MqKb3j
rFBaklbqWxnR5fCBwG4/XIDueXK1gjUp3LvSafh1MAkkxWdXv5k7wLwDV3DKDgPvjNQBoAYk3B+n
4Vkk7+EJJ/tGbN3Fu0K/3jTTJra4Xg61fETPMdlGPlOoBBBz/kDkvDvePI9Kt/FJaIMga6QZlGvq
jBTgbM0jZXeWlRRsF99xk+n2/6xc4r4p3xr8LnUtXjjTlZCvC4mx+ZywwR3+UPgTvSC9gSlxKwTr
JDzrCn1UB1fIKBwH04721cYfBnuJ64jrev9yHdR0i5Ok2LKiO0dYvfQFNX121P5NRqLvZi3UH0Zd
89PtqcLDo/iHcef80gZ0OdM8K2FYsNsqNbNmX40MobAQB1J+pEkNPbGfRYE79uOi0x3XYolEQJ8i
IRPAjbpFNMW7CoJnq8qW3pOa1PRWYcgGEdLbgHk8GE7mP+JJzE19jddzFxiVesRsQMS3ERK35Ee1
7VWqKiisozLvM4G/toYBszJq/KNgxn8CU9Fv3KQlaEM5LW9S7ct3cu0cAN0+/6CgXr+TOcd2losO
wc+bwjt1dFAY8QK6QTlBs7krqM1f7D6u6PfnoiIqJzcbwFATKRSVoH47JjLhRwjITlpswSdZI63w
K9hGwHouHeXNpPUuSA16LgQ7NQwrI/8rF/SGYJtROSJ2P3UTdUS3z23kUmTCsdpQHlEa8EmBwjD2
cLkhk6Mn/N4psU+FHgHRAVmeimAAxjjEEc7Y/+T+lxmYJQUtrjFmDrT4ArqvP4/dZc4lmhTt0r/0
sBObVALXq/pV5iKOTrfHadMhBDRIFu10g1H33Lo2qWEZKlb8wrMIZahPfQeh+TSQs79cuV+Sz+sx
E/N5sbnI0iZ82stuSzobqQBVFsXKnVwuRn89sgoh8Ishn0+sCubj9h0B+KrK46G0JPfoKmZj7Oeo
dIxRywx8dOGRABzO3zvI6IysLkaqvgOIaoi79pCy3VIoMqcr9Vle4KlazPVekIlVi+73fCOx+pva
M6KEjVuacJfTZ1SzRhU5bvbOr0Z0gZZwpAcB3gSplmQxSjVL5fhQvz1F/d59p6xW5wlM9oXq8dkh
Y1femjO9xMUZkk1Ni9Tsq026+Qf1Ul//bXaVyS2z7nuz7usjFnosfsCZy1b42NVaYTyJMpPTFTsZ
Bf4huJ7zhc4Rf5V3RH7zG15ASLrz68pX+kYlmMlPkf3OYChfmComIEICkyNLE4dB1X1ND3lCDzfg
Wj3BqzBIuk9GYwsM/qRMic5wU03pvmq+ICmPHaGBai4APZfWMsUI4lHKZnzMOYO/m17koE2Ua2Z8
0qwfCXHDCqz8iGfsRlqSD3QdccDOpI2Fb3eYPpQoKddlc9WhMCPgXt8bD4G6FDGFBAU2Q6x6cXgK
LtWEixL06IyEAElcriqe6C7rSJWP34oYm01ENUTtvjAjNiTqUcH6OC9Vdam5qshwwpP9DHop8eaF
kbZ5jaqFQw45O68hwiQbSkeQsOitI3AnwyPCPHmAumhfaNhL5XQVmV3DFwL1r09oC02BM9OyFtGw
1TQhom5x93b1sPjXfRmVTtxLYl1P/gCQ8wbFm/uRVaixrgRPvN88NB4l2SKV2kaubrUcCWr3k/9d
0NngJUgQN95Oltvzagm8UIt0hAVri5jKrDgKGtGTALpzFBRlWW0lNnsg8evG9ZtXtaeIIKmISffL
uFq3Z4KKJeLcMWRzWqnOWEhJ8MtB6nSe5xWNg/ByeAiHNw8Z5H7tPVdZOMdRRLchMWdrhsui4iKu
FgiYvOWbKTzLq90U2GeA7Zt2YrYX8ggyB+y53LWGf5vr+Z5iaVy0xSWoGdT169eeR6llzZ5i9w66
uzT4odyb7I79FpM0+kaf2aaWdbO/rRaGhOFMby6zS4tMK3r/yGkxJOZASL9Fpt+ISXjhOvkNRQyt
xCgNV65leXD6iDkX5IdF89Lv9NluwdNRD3fKISA34kB5X5fz8EeicTQqiHTJp+m0FHUHsU+jXw+O
VF/u7FZMjKGptmKkm8Tnp+ZQUccAFMtGyJjiMCo/o1l/ulcL/2DCznk+2DJDxzaNcw6HawAl0RNK
Rc05VCHd5WOnJwPJr8rFg4jH/5XszsYK6qleFFm9z6F9z41zhpcKw6N3yfeDjO0B7PXgF1vbgd5L
TOZ8eL1qlPx0HVl3UaC5jZ4+DZ7m1xS+3GoL+8y8nBH8euiRbaTEfoaKWx2P6OuHYgvfAnsIvFGu
dMw5yrhWrx/I2ahelgJ1Ne2wWP2PmDC/qiGaFgca9H44FI8DAfFZyzReHCqZayZweq0veQ0wo4uo
f2iPaziRziRJQSJYgy4cvGwvLEeQ26pLb38GmoezpT2w0pcIeIt1Rvx/nGDJLiM1T6dSEoYB/s46
x7sTB5dGMvvV3EjgfSFKiaJU0Qd9CfEuBS46IIhWYFAEF7Lz9wC95sAtR8Vr4///G7UEF3tP0W/i
aoWtISQ21G1nyXkgBfuMaLmqKMb2sfLwTFpZ/z0yKcu8QB/94XTX8QfMuYJuBu9JMRZBJfhKfzVq
GUA2Ef5jO0ZLffF+kwqLaW71BgNIFeZVzkmcVsJMoznSRACtZTFNBdrp01Mnn/6o25GKZosppl0G
DTH5wBNhcggB3OdqNzD/BLMYCQc/4YV3pmwDBAd1pWM+12kzXRMsanAJy3y5OOUKAdHXAaO6/Vb8
u4Db11GeXDINrqiVVN3slgyggYkYoY6BO6HAVeVq1CVZSRRiUjv6ojcbxzF+I6qce0yY8+/4FzmQ
5U3KI5Lo1BS57ALmJEXZFVaNqGN5ErmdEC+92DqSSvivAI6Ah3kpSuyew0Kon+x18K1FGVCZjbwQ
mtESwn3xU8UpqC3NtVhXZ2xrzNvpm+tzCmOrfimgRuGpaWCrZmMm9EvecRpcefaKkRwB8IuFnZ1D
G4iN8HzCgSVtBK5UnocNejmIeZxauUKEBUUtYaCpuBsP2NVwDkr8amcNhkFHHN5x3l9izfAE1lD2
DWTqZxFoDeCmXvvXXwEYQpZeURWAivWO5x3EZcdbhUBtirpRn5kxk2qWdfzP6zywuQHGCcS8ceh1
aemqF//oZoM4utYPdkCyb5fToSOZrUrfSZkxtpuGA587RlNl+Eoc5V+7vuA1n5fIJrioOG3NlX3d
KaOGjNROG8ryiU7ojXkYqpT7WDvBqJpB1uwq92x87oUk5POH6jfhf49n+hAoS+mWf9MGPp1pBw5p
XdHkruOg8C36La8ZXN+zlFCdhhAiesALKSj48e0CzXTlVsCYa1bbfhGLyqQwy3unhR0Uqeusa8dp
5v3WWkrzsLdnCu01C5lzCkmEoUXU8imIvRBtzCJUS9UiCO1PsdsueriZ4hMOfsYne3WrcBbLKr3a
B4MnLeSEXk7AX6xr/iWC+Ubh3hqawySPZwpJcGyQig2MJ24Ir3VfbZK6qNlrjPxm/bAFOFbufMnj
sFn+W/Wg0kfg6h3nOMpYmNJmmp1EVLllC1xfBDSRgxnRtEZmuorJyHllg7agDDc2P3j+WJPk16h7
v2gt/4OmYZrHZHAaXlkxB23VN1jbDOhcOZrtSamVBy4soXdkIpdgCG0ZsBHU51zEobAQFK6eT0GM
kZsaZv1rLdigYAObAHB9NceEyAQfy16OqsLNjYU/cLPQ3GH1aHb7U2hi2wiofdA0jMpA8FnnuxE6
/tBgTeRjtrp8ZxZD7afh1g9VAqd7K2E8Vbn99N3a8yActLanCMS744VGeKMDxfMQ3kT0olxD6S2Z
uVcftK9SbXmzxPK7fE3Tb0YOoiJRRMTcmDrQTjuLsPv8IEzMYuKp4yi4clPIxf9Z9oDq8snsD/iV
bA7kRCk0lyOZ+K3HjR0iex7WcYsfOKKWh+R55sUJWPRJxfieeU+aL1oixJcKYwQZBTgLXpwn88An
ilU78qIeYZCTJQZc1eoCeQvC8D2UlDXx6gZdFQcdlb7kwG/ahXE0HipRrSkpJgw9e83Fyk8+UtTQ
ZO/l8KKEAdUel+KGI82vRWTqlRFScClGm8of4wHxw8qVDQTBADGeHuo+ZbjVtFWiwLeAv2syIMSB
9SZQKwRKRqiKT8I13K3klBW9n+IZmnV2fFGWYdD45ebazBl2NJLA4JBkkaCsUJiGW6FzHutoNbxo
TH+kfcmNSPHgnhw4QCyvs56wYSPg7dW2ifJGy65/r6LQAxATMnD8R9iIZLuKjipmE8VQ6vwiCT2q
8ypWf0KMdqstegHpRiZOttgrNtEovtYfnX+YTNhN458NDPBKun/1Ok03p/lqcFU5d5qXT+0WxDkH
zYkALjjXH0djklYv5yAbjlW8YXRthW/wWTfaLK9xJg5CtLE0mD/XB7vHD9tDPV/98ZN3y8K7U7xY
tFYfU+51rVmZD3YE46mS4gLwc7mhch5QE88utpRw4aovkMV6Kkdt5CVlyabS56NKnk/WNEq8FF6U
CIqERO+x1Ju9xqr0Iv93QUjgmyyGtwZke94wpyXNDOYaRl8ehseZZCJYy7+XYg3aTDuEjD0Yq06q
j0ci1lYgAl0U+1MlFPZE8Dkd0YCsdsLV5Lc8FV4jiOf/bedUqP2PAKm4ayCZuHPCnM3sbhGG5dWe
Bnz9BSID/YVn2vgWF0Czd1alEA5LwkrYJ1IXxf+LjEwphiYEamDWAzPVkfQPkxXh/SxjxS1zCDIq
CwHH3wVR761aSPOqIHrH5CDbwWJpGy94Mot5WgekvKqm6uM5XmgYulj7DJLmWxFEmWHE/KLdJzgG
KQLLcVNLWK8EBFatKeJUJU7MTJKFhWK2mDVLdAgYWHRhR/e8JK6dPhGS0Z3L4S6aGQ8+pqJLQPIu
6zvdmISR6ANb8jEE1qr6KwPz0K+4Yv7b0u7UwlR/W8mxf10maf6L1SdBOKX7+p4Fhd8NvRsOYgE5
GqOoWipyKxfMCZ+nQEe0Bcw0mvjy0FV+vu0quTdCH+mhperKWGhhahbmjBCOOSkjPTfgLZE/XzYT
BnZg7Uy+DLWabhx08YxYNWTO23+tBJFYplhA1556EdqSaizDb5roqX4ZVzpkpT7k7zG+TgA7Un5D
JPKVGfg1Y009jhvoPcBxWwLffRKmJX41GteNaJUTqg+zNIr1O7+5jRU8tlPqOUiRcCKXJVQj/adI
FRwwrNjLcI7uK5owppDcfh5+AomiTpGnv7/TFy22jSWHhHQTkBgqwq4q6X6JGK6181wEmd87n2Jm
8MH7HQSE1iPiZqNe2vYtMnSmCMr0g2kplR60E/fFrpfXGuzp8XVshn44rHhpN5cA8PsX+P4Sb5qf
LUsXPTuugHYZsTTCywR3Zm78w7NA65/nuDBiMWubPJEWj766U0/MDeSSkYGC8BkFBc4XAcOVgBad
TT2zE7YHEZ/S8PwYghvONUPMqJuJmDqRphHUMuiX2LxGErXchOUo8MEtMKHUlhGpw+CosT86nOBU
xoPTjGl5ShULni3dAxseFaOVjqHLSODvgjVWSGfRbv14YNfsV+B9gd96xot9cKlORh7EU8owhm+b
30tGIthTLGbAn8E+7IHGnYs7rofMQ7MFz2gEVr+4btPe+N+FkaAygZ7B0xC8L6x3ydGkydWxXO5+
Drv6XDmwZMhuV9CpWLlZ8ESaevZk7uXEPwfwTebTR2ru8mlB1oSAsl4Dq1gaYhj8whdV/Up123NL
fcBdy+DpTv4ezDFN/rDT6SMcaShV7vh7z0zr80lCLLzxaRDCdFhBeACj2l5dawhRoYNUuefCDD50
vRp0snMluflg58hnBNy36u556C5Zl6fnDX0WtwProdtsMa4YUjLMgK3sbbXg1/6gUbmtJsV+zC2+
g+W9UMVooC6juA9dKI8QLkNNTZgO8s7huoKNhIK3T00NGzLWmobYXq8/X5DDxfkfmAybrMEUrQdo
tCEnMpQPiU6mEAST4cYAjT1LF2yiXchdK00+1stgZzxpRZudHUiXEx1vJ6oRAzS1KEhwivb/1SXy
zUciv/Mg+I9g9mrzpT2Ias+AGE2XyeBWIwaQyyyyiaOzEYQStK6E9fpoi7BEq+r/AySgkWc64zeM
PGW5GCJvtvsSBaU4ZxEugYAruFTamc23yW/wv915Y3OW19mn8w4LRrCrHVEnKht/hRW8BLdBJUvK
OHEnxAgK/fxEoG+GBKquCOFyaKq4/5hH51n1+sn3NBe5WTiMCKmvPJ5JZS1HNVuzzc6Vinu7HbCp
RkzouZUPowspaKSDCk1xkEDhNt61i4aKxWqrYtatDWAXfoudv947nwU2asXKd2W4YWJZRyjwRYF6
mEzM6JalddB8/Wc9UPwAZ1/w52VJD/vJtTa1ZvrF+N3kxcxIh8eJam/uOZq0tK49Fh4HvB6QDLGH
JvmO0moub1T+D348YhCOk9lhmga0DRkQT+RdRIXdIK3m3b/7hAcyAhfia6F6hgQRDaDBskZiYuKQ
mOziIIZ12dIUSZt98OH4wy60v19xFfKi9EDZMZL003z5w74Aym3ZSNFC0Xd9ct3EAh9c/V8bU9zn
ih+aMyM/Ol1rsS1EroYf2O2JlJLtg4FKm8Imc3F/WSDmqVo4rProHomks9ZvQOKy1BfaA5U2L3fz
KN8PbUvI8CHp+XWWWyziwE9MlGqhTi6abrhvtlb3wKEX1CAv1UwHhAUxBpoH1IFiHIIlmU+/OuTT
aK2+MaYlz9f0GU5HPMslFWCOZBD7mnPlRe4YBoIQVUG2/1ZA+obZ16IKxws0x6y+h3u5lFk77blJ
HQrJEGhXlZIW5lV4z8sACHuNh1iiKhRK0fbq62oFuKw0PvGDhZ1Cc8pIYkAnIG8+zOKcPsp5977U
Wtcj2xsBsl1gCxK1UqaE/u5RjH+iBJ7akMcAw+hEH1tbU01IcT8OQCXJEBFtQ3qyeC4jC2+MUjd3
/Hyoz52YJ8hEnSsehSOVMoG6pC759nK7rCzZc58nwNuyLrw/XvRKyvcNcJt9NeyYYoreIsZY73cq
StwWp0UXiJoeOu9gT8Kt1A102uw5hAZ7vfzkcRx+xW+ulDtFP7slylJBJ/KxyF5yGWPHp8zkFdrt
+NXdJGbDWmKdY/USNeMkcWy8kpv63k5aPYLaNpVjyCxszepTVYEVRB72d55y/AKPWzHRGqoRt8ya
VQOI2VKBdwV4TpOD2bQz5Lqik4WtwaEo1sFJhoNTT+8sG9a+3nzQpkGgNIhp0DHTHRZYurCpOIIv
x+ZrWnaX9ypX4i6Swm04K7rzUtF3xoIxCAQvrgn3/fYvboy5/JUZ2FcM3JW5PMLnaYhTruBYTsov
wV5U+UtJGsTK6GMQUrczVvOkzVVGXnlmG7YzIPAzBcknbICzZIkKrqpwBH1HjYaRVbgpYZ6Pxvl2
ufXb3VhSZ2NzIBunm4TpVfb7IAO0+LjrAjVjARtxiLjamT3A71pt++l9r3dpURyE69ZxctXjIsfI
vNYnBsHb0qSgMX7TxRQ0bGjx64ejtOJ6dvOXladImEipDue0PmY7x5hi+juI+xHACcK8Mn/6w1Nd
LqCwnLja4iZjO88V5U4oBHTubP9hQlAcUdTymMUNSAiQJAs6pgPpIwr+zzs4vLInV0rYu2oeISuW
V1G/w56z/wXuuzBFbkxsnFRyWexkrt/l20WcJe+n0QAnO7p9ltogGANfBnkrk8UHkDjewTpQP9yE
b/RIZ6i17RnnNZFkRBRLEUOQy6vUn/84EpkULlSue7AQZ5DPm1C4a0pq6FoW+0aQTJnsrCUNzEM7
twneYng50afhDfzDAUwwstDXiVeymWostedfMOmyLXdskFYoK4VMG0UyWStC3b8YLHICoVvPOAsB
MnT4R5QkVtJiLyUOeCAOE6OSVSYjInsiDGjGXwFNikJT69wZUmM0oN5IO6CVklwSbUVaAVXS7sAx
AL1eVO9uFWUMMdp3tuh/lmAyLt7aKhfl8+cDVDCFUQ7oiRYr7aJxd7g6A8naNp96/a7FMQuziWYA
gZtr1pIxhkLCJk7dTFEozwkkvwrXi3VA9Ibdwjag0BnJwAs99co2/xmOcoL46VVXsFecnbVN2AWQ
rsk6hEi23ZuECuGrGl++MH+0eJKkhQ/OUWjLQqcYhLaHnO8aFFvSTT+uNI8Iw4R2+B6zc+V/B4MJ
q9VJ/0lIyPKgxABuZ15WX2BX9fqZWNGTr2jbdOZlhJAzdHOebSAv0yvRYSFC0YYZ76DEG0U/HW3m
dZ+XV6IY+VD1AJ4j0ZW4t/hhx66u0HShf5eehyJB7wbFulS1w2uj/NTmOgMdyf7IGbiEXGgXd1u6
Zl8vgpg6TEVxKcfWtmVZqXAjF4SfbWHrvWrV0vdNdXXKBinQNYRhmN16XVRrIOWLzqbgeLIYQ6l0
d1Q5MJQv8kZ5qQaWX4ra8udr9ZF++HFCqNsbRP/olT+8m1nxhTl8kZDNmiwcL873BYmFQt2plME/
tZlC82NDm33/P0KNoYPWWAA9PoIsxmUZTTRn2ObbXuzXeKLTw16QM/goD1aGfSi9zkOXgokDvgNh
OXwlpUWK+U9Uo38AohcxHAyZajlJ1tpXiGB+9NVE0tKimDTVCpY0JLU0u4Y9Eia8fcWA7w7tki69
V+aBSHXY5VXOIOXRDkP5jgBe7dB3BXfpE2skb/dn6trEzEN6NhbhqnYoNy2YqM7vc5+CrsJJaX4c
uKDgT4Eu22HfHQf6td7pBM2qSzXD+ppNT5Vrm4xeS1L0Aupu/xp3TBJjdOLyEC0RZ24dEfz0V18m
4aEHIZja2cNMj+oHBeyMVx8ZaEmwsss7wnib53Aj7ZuB3/8IXnc7+9B8qvxzrFJltJHhMghx4/QT
66awTQZxPNwsFULDZdlmx6Z0O7RuNOTvc33D9ZDJ2OJ9fpSvc3AGkm6BF0xQq3PfBOvsrWF/FMp/
ooLeejBi1TaKioYwvXH3l5LWKBWipXhDcigUsBMyD1X6xfdYg8Ymv3fUYb7qI7GHu9gdSWKHQBZb
3EerDVF1LHS59BMT0pUgLDLe3VqbqqVejuHH3cj3q5pHEvcyNK91SRi3AlWnnjOltbo0mzEbx5mT
cJezKEQt157gXYW0IEGRHYkaYM5F5Xo/Q4sB+qJFp79XOLqB3gYR770l5IVGxN/iWpN9IDcXIUjs
iS7iZNvS9vKxtuiZBI1P3cotJv/xJ3Wb5Ailh0XWacL6syYiGOPAzl06FVXx83UoH84UidJqsumn
8XfbAv8VlpmcU3ahEo5GZynCviWa9n4Mnimi4r+3/oiPP2aVS3QTyJUz+jxNtMCSBMaPH/OsQL0h
sUsG/zfuMFpUIMm20k1dUsGeWM5q9KNX/I+BvdWwQdUv9Mt2k3HU6dkiHRjAtggDTBiskTruWBXT
3Y+t8FuEmTmLgsezh8OgcJ+3WJfOVBPsqlr5AdM6Y++aPEl/yqbF1W+Q7OdmBjNtJt2rm4UH1LUg
sZy8CHo9Ezh5FCDnGasjXW2SxHnLUCbxx0GYY5TbEZadRQly8AzNATKEMWjZjt4rxSGVYUCeOHaY
XvBauJfysjzlvmPkIXkkzftQS8c5xiVr1aHQsy4wDuU6kmo07lErbxvwSqbk8+2ZECU0kL77tU52
cKipQ5y2JwN9pui13uBpusLmgJaQzWHIrO5hHjTiopsU3qCWrmFF3kZtO1qA4K8VMPR0Tp8hx6C7
AXa+rzvFPiwYRnsfKwwSxnfeEQjCkl4AAoY2lw2MIem0a5qwPLw+YY4t26+eX8ft9ZGzKvS13Htl
k6C5+xNpbNh08IQUpdThjYz2mtHcSOx6mPsfZ980nkE+IzuNdB327Grw9HN+rK3dDzU20xUbdN7d
satXUA+VCigL0CbZARXKilNx2p+mgxnOeHsiEmm03fsHSli5LIfk7lAXd83vVDEAUaf0IJlNtg8P
/WdvCybqu8Ay4T0xVtTRl0Xnfbv8udIMpYzoK0WuX3XxqIBzKwDhboM9/SwduJgoK1mgO7m1xy5s
JZukYuz6TE0357LzNW/Xg7t0qbyrjZjgrrX5ClIWKhKbsbaNNS/81nguwQfED7xcxKyEFy6XaWoE
b37+0BHM8QH+hAJdYCQ0OfclmNjuS7d7d0isUFGtMjE+uUNAchx0CJa4XhYVvc/PxzxUHdDYVAkE
Xgwfn26KsAaL4mgBvvPp+hhbEUOn5/M6yEpGKkiwOygC4+k0PrmxJB6n5lgqIuMlUqkmuwvMBIdS
PDX+n0BSNJlVN3ZqWNFDQE5K8qqCUXqmAZiaFVWNlnpDAQrsC6VXdgjrx43e2lU+qRKtE3XZi2ne
8vDV/nVpOfBZJolVkQsEbrTXFKeFx8EJiANlGwCjVRNOBfBq6KkaZXMpUvC+Y/8H7ZZJRQmWyVLq
nZE6PgZGJGpaHVmIiamb7JeMXNOGPlyZ0Qphf/dL+E6vJZN8O6YVB8Jontx+mPTg+MimGUVc7/Hn
YGtthfTkXaPMhgkt9kSZ444JOa4tzzMAvo7wwJqv8zw1GH24RCmubaofZxyGc3C3PQWT20MxFqMm
Q+CDCX++C77ESpYVpy+wCcyJaIl06R8w62Zhj79z5fYf/URsyyw3/QFWjIZxUaPkefRpbJNsokN0
UcnUdoDHms1dh3vbaRnq+Cs5YXLDvkLPmZt5FDZ/JvRb8vKwSBWLzbYLNImsREX99Ne1o3tBvFWK
fOYcgKRMyKCM/2gD40c1QSEbSJs/uxX3ZrpMchhyLLCmQQahN2JFhngI6qrNbUToLfWWvrNEEgcs
mGKs1wPz5Qyw1Nv39L4qZ+WIwO49JD2ywaVnw7N6isVJnegtFnPaoagTvgAQmiYp8lMFn/1DeXck
WrMjaCqEqqoAMtOB1CX2y8h162f3d+fxwRz+WKj6vC1QWXjnoyBNKT/dvx8tjv0wUR1QjzMzdmQ9
m57g+UeCGS/u3huAEPj3bOCssH+FwwFzuefkX/me6RaEw4xO5DUPjipuBhwtgDve59ocKKKOAIts
U9PXEjNOXBZDYhy++4y2YjDmR5YMf7wDIOiQvGsBQmbWRQI5ZY47tnuTSKZnCIg8knoOJ9WNsMjn
rXe7C1kIpUsWec6+NZiJW3pbP/d/wjUF9gKtE0UgtKk/AKipiKL+4hQLKCqPpZx2Uh4dx4dxKlJu
mpDLuC5hXOua11hIRfcf7HpKYKFZ1kYQ3vsjNZmEcMmp2O8/ikkYBDW8pRdbyWrd8R+8Xh9sp9iO
VruzkX/FJQvCsBpL+qgxwFMG0Mo3isvd2OhJVFetXCYwXUWr1M4FxwfKvJd3+J1OxdILsVe1iT3c
dF/DtyVQFBeOzuLlcNl4t47CRTVY/ckLNCa3Z3AdSOOPYvKbsLqDLUF/dTuIzEe3tFH6O/d+OenR
xTzEaGvs1bAfamxpi5qV7QhvGeKynJLmlDNG5nW1yyEiS7ZSuwoDU0XDUCChsR5Qy5FquZgj26T0
VSv+u7I5PHag0j1zXNjRog63rJ41kZXYE7n0c9oM3cCqjPEbEMq5cgt0RTO3m79CH+u4YKo2Xd9k
J9qeu226R9TrVmQIDWlBVDqCD+Xq+sdgUJcpLFssKiBc3uDV4FV56JDWKoIa/1xLkwm7bBGItzod
LpKcvgnM0eoknqC/t5EnDqRfkVrfgsQWTK90ICGayVYpYLm4Ln5OviPX/IymHRoiu3zkKyOBo12d
Yp6JFVJWcb/OKcRO+QLwUNPrhhKNOGIIYSg2nwZuz7slB6OlplMpXKFjRfWt7XiOUIcF1IGzs6Hc
BqoY9AA+XFkZX7sysopb8GUHa04uIH7YEag32z8yTUWELSH9i34umJLNXRFX324yXgHjVjSzbEV/
Pno3oZmTStPmesFIFjduoLZ7nt9YSUaM7YQhNj1WofNOWs+Z+lAnk8RYKmiSQyNe0ucYtwOVZAJp
bMEuDb3JQXWFa/3mpfjL4t/ZWUJwMYbuBnvxuPejMXMe8Bci91iFPjG4Ik0Wfh8jNW4mCTwpQ71g
UZHTfKUYG5ozuv3NRZo+Wqr+DXtBlIZtwKeiw6q8Rvn+q/HSvN29efRaaV6Hauilhh42epOE8yPD
rHA6aPUF26+BOeXjGrSNZ9aGf1dgPRpa2itOyEhh+163yYW4KFBtJDS2XBQANIz8umu0noHQK59J
u7/0wtBNb/Xeym6N0gpc06pdt5aMb0Yrt1w0jmfW57DLtDwNPHI/3slqyFHVnrQWzc5Qa/0cU42M
MSzwdHQg7n90gcwOLVR3gfHiq+7SZ3wm4FiKydHhVDUnoHYXtIeYN/tjolFCMUk4xEZsm4uY0wyg
B3ETJ3zYSgnEWeiI0fjx2Iqc8hxwT8Tzqe+wS7KMDVTVxKYWHpcV+W8dkWvM4WDb2d9IP9aeYqau
+AnGuVD6PuEqchytUlU4dyAPgy01NXqZK1JPtSmgbivmIdu0texVQVUAHS2ozqkMGrxuDJWokkNR
dVc26gl6S8a3SSvbMMjxNMneuOf3H+2692NSMHnOVhhbj7e5X/r81Owfy+EJsZ8/iB6tFdo+XCJB
oL5dxLSC4PDC7OydpWlQ1Lx1tINpTOASQHARxEm8lSBPsAIiOCx7CcO99mIqck/sdyTeJThYhzEf
mkt7I6niXKr0ZgUmyGNaQjff7n4bxXSp41jyGoMhQHwNBDAZJ7clTpjiN1P/WVL07+itKnI4YlYd
SI4PZECuiCm4pDwwsyOJiAkTvf7S7q0SmKQSr/vflIe6Gb/qjLuHesvr1SIvvwoTeGOq+IFbdLDW
zNd/Y+lhM8LqoUk9sakBdprq4QwjalnZPhuQVIz0AP1GxGopPBBwd6k6s4A6h+pBSayTqwaqgqrg
OxVtnXA7E2HjjhWZDw7qI6xXPqis1b/bSJm5FTcyJM3i4nH5Z3SlEqmimsnQKHVS9ynEPbm2Fb3P
h63IkqxO3wX4OatEYpVKyukv3Ki6C9j6HHXNhxYIo5SWfQpNILx8Pyx1e0TlDIVH8yUqpKgz9AXk
xwmgYDpZn19qoz8oe+Ngf0MBiHRLfsAVSG79f/HPAAUumINHIicq1e9HsifAsRMF2J5qAj6sbatS
68VmITTfZ8G9YnUCbyFVtlst1MMmukRbDyHYw6fPROIbVNQ0ypNLvPXGR8ZoITBaLwJCE804lqpy
MjRxrUyxR/w+UlXGYwvsl+vxRO6LikcHhwF9acP77+F7i3bSzQOJ+y78ebADvTLBi25Rb6MYTrbM
Zqxop+Z3JJG2i0kJ27TYA3x0DGg/i+IF3bUn8lxJ/LtjtO+fexOJHEoOokKsibVgfqdnNP4cluMZ
9dhWihmB2WN3fcKUVfFRkQK7yvxF+r4AeKlUzTEKZkuvgyL62hmwhC/dcE14imEevTelmh6no9aw
ruW+81Scaf1qMhCd4EJNfmA9Rw27/LJATcDqunLk+46FfqwklJ7bZzKNgHxa0oHMX+qcTRL0GNPF
QLCsy4pq/FRjNfWz7KXHJoHZ9Q1YXjHMtOhMGF3ab5FdDOeiNQPyfELUIMx1DkZ2j6OtnHwnpyeE
RtoJtJjZRwRlwTfmkWbU8XkmsoWJECivabQpdU5eywC8Km4CS8x6C5hzP6DstmzAnqz1KwuqbFFm
RvNe4XvjojZai8LX8RRaZZZJGKfebDV5WbSlriQ+g6BVNFx9uj4KxZRksrmAhtjE1a/ZVOvrmQVA
2AzsXZaRto1ecPgW1GgHTCirc20wGzOXhz7rqLCr1jMyR1KXPJaKDuGdVjOkraErOKP2HN1siFan
/4WmWno0lPOMSvOPilCa1sZeET/OZsAWlhSwzm2BhzQ2FYQJLVO4+D4QH0Nc306qlkYhzAxW3lvl
o9slQ4TWVauDF+rWnC+QowUcgHwlqyIs5VzRUE8/UeiDmXdW0SX8WR+J4ErBxfAp4OgYRkj8Mdp1
tsgGXQSrBlmj1PfE/+R65kfStvD4ptOXaj6Ldn13V2DO8OaLa9kKFPggOnfn1pmPBBFpJuMexu5S
R0Ah3JBXM8/C4czWQfIWvJvp7cyh9VtbCLml4Xnubp8cY22lAURP4xKbYgs3j62MufZKfpBan7Hr
+bh0VdsHvtdKhQHvtLG54OVimiVENRQZh2SOSw1JIjDfMMuOhIpcPRhIhNixybik0Erl28Xkja8R
F8vkun4K2sK+UGj/CfL9H/oVSPZd+8xyA8LgxMKYwHzyobkNOiQ4VeV3APFpiNxEcuDPdFDaoRaR
9V6IazBQjWJDcc7WJFEcfkUX9mwIINlVjTh5DhEcnoTClUHAHN3AhGNpEzm/Zqnd18CIUh6e6eWO
roqRteYhEhI0RSQOljH7nbkNkSsfrevG04E674bj+JB1oNcXEeYIQXBEyZBgWrcAzE2bFe1+82Sv
Rgoq7roXloHdMgz7pwkr5lLFYwBJ932HIsr2xRgfW+iFVWiZMtUJnpezjxqvw8nUgksKsxl0AsSx
iBFL6xc3v26hO4uHbBAmjgKyA8Ejso3wK8UGvcNhyh1HJtpGarYd8tJ3nwTXEWqA+LIXnkyez/6g
sIAz1nWdA31XZ/DJybTZr6ld33hWnDTfZcmY/4vMF57VqeTS6VO26kDaeBkGDiyidxPL3I4xbSIq
OXszU+R7eqrQJBpARiQdYglrYV1lg/LTIhjnV63iAjORrJCtLk12elynUpJn4n5p7qt8kN9/2kzt
osrhN/PkEpGT0CHFUoq3XUNrt2aVLKfxpm7JIdmimy6ivfnGDPt6eN24dt6MSrjtCL5HmsSd+puK
6m0DWW04gCah+fEnU4unaKF58LnXHp1V1YbG/9voKQEXxw9X6GYXSaEcc/9FKHKIdDlyAIJ1DKA/
jtmsHrN8v0SxI8XiKh2LhnHfd+dk+OzYDXQTxB+dGsOgd0771m5g7ml6KjAPFXxO6qRh+fZ1N4z7
AYKaVbs/o96yonFl8rq780etckj5KxjkeW3BjTFqPPhVwCOeKM/Qc1Y4zSPpuZwlhIjkbTzSHAwN
qUZ40XO3EhgGYp6Sxhm3or14e0xrs7dcDiQRYacCJePSTUyBe5Tc9skBpJFJ6Y79Jf3CPkuBS1GK
iuQXHyPuLfPMOTcNxQWEXRoLk1sYSus9mi+i8gA0SlaLuK/7ZR7eB0UKZ/vszFgp+rgXaInUvkDF
4W3IUO1n/lfRyFEingBQ2RowVqUcqtEtPuA76FPdLMCXPuX9ZGgizWA5rcCd9CGXZMasszKvNRoy
9a4r0Kk0R9wouXouXMuqcBhlcMoHctAL4ewEOJ9u+Fh2A5buBIP3kVpYbmFe72ecLWJE/sBuk6rr
6R3XaZF7qZcGcDySgJeCTG0i5Z7P99RVY76N9ogDLlJMcUP0egQJNoiZ7pe3kR5V+B6BKpV77qGx
/BiHWpyTP+zZ6+cFd9b3npjuCwAwG8qd/bRKE3F+2Y/pEZkPUfo/xzfLlHTdKTfCSQBYy0WPhXDU
Xs00XiC79R7Y7KUb7kjqThQ0KByy3mZqhoZQQzbV5T696i0sBGjw7KfjQ5sSXHBazusFMDtlgcTi
YX434a4Ky1o3KNZOb29gBZXEyHFT8mAR7edb4RKQ1+w7Aa5NKgtOH9uaCjMQgy+v3V63zD0yUCTr
WM4S53iM0+uf8463fNn5m6CEhMxAr3dMCkADVW0EOFDYKhuJz1dz54IJsC9Iq7A/1akzVFMu+XkV
CFACqHY45+em1lFcoZLmT1Lrylt0at3I7+Gn9WpQV6sKvod/JkwyiYLuLLGMpK7x4HOfgMqOIE+H
/lf5krz9EDh42YDj6vfBBy5HowbYfBhdghBd5u8xC8zW9DBA4IOCm9aVISUcX96bso9zoILyT3vE
9FlBqyRPw9TK9sQqr6our2FoNM5hy1kWcyLeFTM2l0/7qAJuOCvF7sLQtRYszrLcs9q3kJzyBESs
lfm2l6itkUn/huGBdke3IHC9Q8p8g3KcjWZIChiqMYdtgWq9BZg4k00eDd3YT3gxFSDYS8J0yjFb
lLRUYejrxO8pgYPZDwHdfgI218SxO+jQF6lzxB9LV3if+Ayh/E/e9bDkX+JmOidGQ5y9kGlOCK96
qDSxgY56sZnMZKzSX4UMtEOWA/dljPDcuoPz9YQbkgPozB4KEfjhuA4RYGPYN2Bb8WCZPWDYJePW
HMCsM7Ys7KlN8pa2KmhWWSpREAM6c/jDXZ4eSAHaTUEl4aXoNpJRz4Z1AQhdleSIkKmCwpo49R49
3z3r7Q9Ha4T0bfigEFUjBCbgDNJWG2y/+JI4mYINOzNTe/RPpgpclBVQLBVzlBrLV6aRTlYI1scF
5MeX7Dj+3PLxYeAy1L05iGwpaxfn92qpIKcZfbLN13nZpO5lSWLhLkLcBrg+ojirKyo0dF9XZIah
ajdC2su4bVimLh7nYGH1MC4yHRKvaPjB1WInu/AbCm8pUmVo5CxN/cTTP3FP2929oJ6Lvmvg0kF3
EDcNR0MwUgFbsgZREH+I/rixg8/WO7T87yg4a5kpVX/IWct0mtNsQsOj3FmQ7qbGJJH+gsbi8MCy
+91hUcTkSc541t5O8HJaxu8U5oIaEQOyTjElgWYzuVW2O1Um4yc2bSxHtVzrtEKTXD9apV5F0G+L
nCPYFI10vkSu5q9WERqcExUa+WgZ8dtnmZLI/Bw/uNRXq7iSKDSfN1kz+0yWgMQ1/gp3eVKxEcfF
bc/HHTVb9Smi2sAwkVEWqnfZpzvQerEpKgCK+w7b3sCnnY3PWuDux4LUVcRegJxFsgyfSyh3XPdz
3mIUjl2Pd90JzbHt9UO31DEiT0fal7mqbMXxNPIKo/+Lwv29VFt1gRWff0G6LKN8WmUorzofN0Id
BclmOw7CVplMN+17fSGmvxzRvO9fWrzxLg0kfA42x4ddlAue2nnTU7RdSquKGR5aftr5iUHvD/ou
i8WF81AmWNrtHkZX2k9IIqyPfeMi4aaLGTxpWc8ez7dNDVbHS4rIdhOwtxb1hP/FiXhiXWPFUaGF
/IqR3THdRccKmkfY+epQ8NbUbtbB/rL53UvEjmhpgcWDxdRxWUlk8kim28uRQdGUqIsyhs+V8jke
yYwa7SMzmVBbaYCCc3T+YtNsz2b/EnyeQmje2h+JOiH/2P70FD3gKsFc6cCxOQlnH1Y3flG+xpQV
TC+LS/uiGccJ09Wo1HjBbyxqdOv74lhEPyBqtIAzx4YG9zBG40PZ73cU1XWJhXM0kYqwrXIhDQVE
0xydUhg/dHkXd12CrN253B2AtNo/x9vammXA1PufyaNFrDSkB0NwRwuT0KTmkFqYgchUSVjUqUko
wYAS42c3vuS5g9O0N+QITpOYi/czkWUGU60gZp5ukCA1neqe+iHRAP1X6LYXahUJF0GhOln8TG59
d6nsNvVryfw9NzaiJzI0XadTGYDRrmjxFNGep20QLYlMEQlpCGbTIEWsEHLPouaXf2+azdLNJBvn
Pmje93A215rSgls67iH3WIqxmuIS3Rs6bXb3aLRaJDDYRSl4Ihrs4DRvLpZSUZvXXCh+/IvWSBts
LJdYTLu9bmNnMFn0B4lzKckYaM5HdQwSFhYE8Fl/dua2VrGVhqA+czwzUHoZBVmlUDdhu6uae5wx
Kwg3Qc4J1i5GJVfZJpldaagukPLmVLwfGSUWGvSpmBX0daWhaEYMgcWBR3ablj4gUMXdwhGwbQuB
Bz8FiIKZENeDly501a56QXbTu4JJVNWVPV0N/wXPyuBiFaN8aP2hT6EHNtKCffet1vvkfsjMOX7W
vyMgQzabdg7HHPJEHI9PAFicCdJbAkUxWEns6F6fcye3xN03j3faK0caz9J3xOxBZiCvMZMe+JGd
pxAbfpVf0he55yHjwUrUomagRNr7orUCzZhhaWACm82y7XLiQTLZUQgSNqDTWMnz1Pq9YpqkuQnE
6hE5Fomn3Vbb6CvAlUirrReqbHZrvQw6KDIvvT7YMWFhKMQurBnrHLBqP16qFhDpJipQQYJ1Nin/
5iZruhTuSBo2MkdS7T3R2Z2lG4HqofsTaTVg3xFFTvjNDmreczynR7F3STsyyCchi+24vI6n070u
bvCxc/G3XXp4sFZQfkssXK1i4GbPJKUj3+JRtACWOkgLRhx/JKkQnLej86bcjzMfnAaZOK9ZzWg/
+a9Hj/b4KIcbA1EctKlcsV4PptthtCz2T+riGYVaVbfw5FIoB6pmK7MF9Qbr870Bud+eaeD4RK8S
lGGGe/o61aHTL6SsLExRYdhhPU83wA9xv13vCtiu8OTo5GGbGD5o7Xikc05j5o7k16uzIziEVxtK
lUEkgfNnk32YLNjBs8HSV1N7ukwCJDhADVAnePD7SOrpoK2TZIN1tR8Q5TOsNlhrIHJ2zrZKEhht
FKu0GD9wJnDX5R/uOsLp29ZKO5aKOS88GPEWJH/+NXcRlsn46G5PVowfujpqb+2igWb2COzoEGIV
EHh7/a3l2Gkkd66La+QwyHwalxKo014q84BZ3OzU48KSZ31admzqJ+mDlVqSDQUJPie6SsuIamUo
G09gccxN7qlynS1WMerG7hphOvS/AKwRJLIVxPnQ+0Eo8GCYE4zgoURENj7kqrpFmsRdh3wUFLrp
4wxmNT+4VoHmhg8AAMfNI64SPYa0icGACTf5GnT9YEBl3LcM8ZuXPGJNCj68fcW6dwzUqzavFIx6
tcs7aEegtr2skpYak8gxR2/dR3i4kZQ2TTpsxJldQNQFaGP7Dj/jqQePCPvk3lX95ksTJql/g7MB
RFjwYvNma2i0Y5ajnJp5BpicRRvQmYiFX0Kt4B1v2zppL/jXID6xEXGxCPZSS5WXADezvNBmiDhq
ChGTzHRQN+dq0Z9lvLPxE6u8doH4WFyhpw9fbRHCCF6bzl+H4isWKHK5JccMx7ZtwWDCyDZZUhk/
ailpRqaadtotTJRT/41JETTqXfrrTyw26Eo/pCAnKZfH9fzwkHmTwPdTuQdKObKMlWuy6OIu9EEA
Ut8CC/8Bz0xBvxu0opHLuk4JkAaVbLxjqe/oQoCu8LLSyrQ7PR3I4+iQNvd1Lve2UdgrwnBH71UH
30l9xcch9sjxrFcN4Wqi0h9hg4CFPZ7GnWT9JNLYe2Kz0KUS4/qhuNkdnEkI15MUHX++cjQx8XZE
JXYfd9ldAqYPNPZb/aKaFWU59nyu+H2In1JRu8EswR5HskcVfz6Mjw7L/0zxs46HrhTK2bMGOjCp
4z+cEW/Mg34tGJcu2RWGqe64ROCku8pbre7zFPHs432EoGGv2O8WXRsW1i7yofu5UDrmTpxxkbGr
JkhHuPNVjqLNKnxb2vE+CrnUfLCch0sPwfb/o6JYRl5C1128INvpaMrMwdAfBOgzq5XrcNJ/qlli
M7WCDfcGQng25yaIhDmGdPtHiqh5Mm/crkWW8NZFIC1UUiJ1j84G+x4uefhi0xbrHdJf6/2Za3Ly
YTWUIQOmYSzS3IFgSnmhfscrKOOlQt/H7UOtGmwmUHYDpLnjiJCslQxJa7pksMKSLEbTYg+srcib
uGHsDMtQIyVp8oh8R79yo79L5O2pMIpiEKG76B59PiWOyR83RC3lbZ6I4S9JnvF4nj9TCsBa2BQL
Jc6osZaVjlmf6eF1Qi/r6fkOQb0ih7Lrs+8y0bhwISqpMeBXA4V340itkzsxbjnqx8HN8w59yTe9
BKdgkk7FCJEXsenQ08QQAkKze0568BdYldKi0bS8blPR/HniNCuOrlCUw3DDZan5SgcD3sTlFCRX
HQnrdiNDu5UXpBd8dCgPiIIK8irjlCJMIfBCmsD2EZjn981K5FGZE1qn3ujDGG82wSmBuRqPD2OI
vH9Zguq41zZXZICQmbT8HOSzRrQslzNduw6jmTizS5lPjACF34u7VuZuZTNgpUTm3OBgOJmGW7PE
5Ic0if9N152tQ+ceXBB9ykAD66cPZFXPcJlU1ovBOPXvGgr8qczZwH1jYx6eCtH+cuJRtOzvijuK
nK2cYo1t21RQuJfw+51Iz81hiyRbXujGz5apOQ0sJQJaM8B1S35Oil7Guz0Q4k5b9u/rkQw7RcPx
AUcS04KU8kHvUO7qNT78NPt1lX+zZ+zbZiB7tDEUCALxYiiOJ3KytCaqBXS9oWGrEdBGPQAfaeSu
T1IRMPoCAeqsHHyNwwSIm74GWPcXscydHYn+4vHbm2L4ELakDkRdIrrCZfgbiNj57OnTWpZzOMmj
6PD2/HtSHWpO8O87AwPu072exTd5bIceJqb8+nIpo+dywmc4T0LAv3Si6BcuuqYkLHI69K0De9dJ
I0ZPhYYLs3eIjt3EjraCZjnzLMpaJH1ZCTCdSpvkDcuJDneSD36TMJiqR/EtW5vQ8q+BM4y0jnki
dRqB2eSnCw8sJdw7HkRgIXu+pFz3ozxXfjrY6odh89HwVnStL0Bs+Y6EMs3/Q7pBy2uUHnp16mO6
tCOYSwjiwP+hUzYecMD3GV1L5WzndGGQ8n/wBaUUW7Z4VFv5a5YX4x8UrEsljbQ27sWLT5A04lIU
gWqxM4dresp6yRBxUGNSEywxn++Ef7B6FHC+3pPAg27+kCtiykDDkxq9kuomJxMUhEr7g/934ooL
4zzIw5z49DC848e7ZbdzzjHoLwReRpvhHJVsE765asp/B+tcc9FdzXWygNohNQeKufGowliUbT79
jG0YG3pKLRNajTrMXmxTSSmQH/mU0PKZWGXBob+HOn3d0bOwmdAedP9y4b4hefSfPVwIG962Dgwz
jmtDdSbKMRSHQlbTLQxAiC3R+HiHmbbSk3wual8avMkhdgjR/vfkWnE5LBBw5fjR57qS1FruJhbq
Ta40iqgTHz9aS1rAIZdVlhnye7lNwWdc3DLjG/NsZhD3tB2TMlklhNag8kIripwJoFnIysaJ8tog
5yz5CLtmFGFdKwH3jIlooQk1yoviE2e4IobcRuw/3gJCs8CynmlqPs5V9IZsRffrYa3r0x3Gz8o1
pbs2X7vFbyhhmD7iM3DHbMNnodt3nJ5j4IOdMIHieLjs1GUthZvKrnZf8W7qw7ubjkMAZ3Z3ojpa
/H8mRtNGndcyzCmR1PoRFXocjQImYwiUhg2Jmq+9aLkJAovN7TvHqwlFrOeWQGcLJ0xnC0n1f2Ye
pg8SO68+J/cG0rh9ViLeUOiD3bN69bVMeBXjVDuCaAld9F6fkJitLC3F8vXxG+azw2oesRXQNL1Z
NJ3eIGsvZJO2kQiwCpbpW9G54LKOqhMr/WZHTjVTPvE7xdlKq87CdRty28FIyyBrCBQmbH3juYJH
bk27Avew4jXu7uJUOKHAdIhznGjiLRXaKzM93g46THtbJ18bZJvV+YFhGL5ji3+xgZozlV2HF6hq
RN4wbpI6v0nOyNJw5UAnYzdI1o8jl3xGJGyqp7fqxztYPt6croAIPDsR7DD7Rf+SiwFX9k8htc+m
JNJOksN4XAfLe7kFpNl88INqsTMi3MNYf69fCYBqY5dtSiQj0wr2UbZb801qqc0OlxzFSvq1M6Kt
qcmsOFv35H38IgH27+iwoYpuquhmwz/PEV2HsX0BiEnphxUTS8kGBnrQ7WAE1Lh7iX0w9jJq7Spm
02kbSiNSy/DJUdLDWqVzJ+/g1b0RpDXpQ+q3gx7D+4n10BxgYgs9dEYGf3cAIx5EEY2EoX4WmePm
4kHbltmJj/c+bh7o+iuolbsjKpdfyAo+0SFZWEe86jgIpmxYaocsk7bSWagl1iGeezVQeszZ4oPD
zIjrd1FpiojWUG+3qAOUAa7bwDExNPUysgaFFIkbifA/QowF02cv7z/SLy6paxIHdrkxtlXrRptj
WoTkPtldiafmmUASdOGHvP+eScJFHnv862r/gSgHBBr9aeVQNlpSnicdKL0q2B0v6NJkTf/P5v30
JQRH0ucLK3jRfWSv5vLsVVPXeOpa/1byqSBkT7z2WiQELqEpHCy2luMPWD0jtDzoEsSAq/Tnycav
K3+mnQV3nUB83Z8OheG4ksFyfsEdWk1WZDLjun6nkd1WPAWT2qKNNRHvX8JxFO/NLPHn2GfdKKj2
XMjmexG2LTPsHxap7xCl0yetVow784IR0ivXyk01PPwPXdiiEvGFmuCmkcIXsQJ1Fz08hORHNuOM
cIYDdIEEHVfI+LtxO3fWNlY3Tt0jYh+V/3DgE1eOMS3nu+Je5RDu9hSSv7Fr8oUnv+GG3gtGcVn+
JYgRSJXkj5Le3wj8ghNegCnS1/u0mTGE9tF5UV1k8cwpupQcFq89yggq/SdHALvn99zoonWo8ja9
huUoBpADpdzCKkGZ9TljgCa9r1RZxQ7p/HXDlXau5gDu6FRRspCKkUu3IcFXAN4X64trGdUUbBSG
1HSXoBae6gSMUTD4Y2u99knzSej8yDZhq+wvw81oEXuKEMwTaUUhGm/h5ina933gsaRl/juJ/WVy
m5aUrNqJJV+m6Dp+8tda/pP353mSEb3ndsjgad3ZLWo3G7+FfgYjPRrINAK2g1iVyyBa6DIE+7re
ijK53nbip3QznJycUF6WXvz3YjnE5sM59rfMe3p9DoAwqQ+2JYCzBhUm+VRItlu0dUk2V+FW+k2C
6M2o+s1H2Axe34+ePQVlln4cdpcbaU2+lW2cnWthm75UOzWNq3lS7LupZthi/kRoN9bINQd25KLQ
B9KQTYdVCwEGY0m34jLnU2nDvLkyfamXs6ElhnT5SGa8f0aabxH6NVeUqma90nZ2sfllIZNUuBwI
UPRQ0tC9yNiIJnU6unUjzLGdFDF68VMH1+PiabJ/y2JoDwwV9wXiiuAmSQDluCEREkFmIXjva7a9
AjET3em6leijavyEzArMOUAU1WGxM+uQZCUJ0rdJg0wguMA8Fp/AI/5pe4xmiiOy5j5TseLuelPc
VwdZSAsoNEkAygR4otSw2NWh85IK54PUPgieUKDhs6fvAxfdZVWQA5RuoT7eztHffahF52UCiaDN
IscXSX9sXT2CkzUq5sDkikZZ5kYEDdAL6aJ+sp9ZxaiggxXQ3MAqIEahrMJb8K6yVvFjLSee05hV
hs2vvoNm6rcHyAzIwj+wSSltIJEOMvtvZduH5jpjzAAav2aT0uUIrAZ/plYWdzhE5hSlsxmvL/tU
swEkA+dpLWST9dl4ujWYsKJstn8FJE4FgjYkSrtGHQjazSEqR8D7leYDy3Z5WRtNDZyLMC2Y1wRz
Dg3E00TomUq8P0oOgA4ceghh0rtmDEBCCkoOwBk1gmT2XA/EwJmzo18pTJYeJ45E3JlLxutwn8Tt
vzp1xdjlW/c7/gJOfecWKJQO4zsaABC7KmZu0o+OTQE9JaUBHI9rEdOFJNOpLPI+9kDonbMix0Mc
wHYt04JVv4zQFj+JRTdYJ/PGI+ga12kfssMVRfjgAWmISakcnLfwYCQo4sV0yHPoveOWQKCRdSrG
elFgLQ9wXfgogjM37LiG6f1r9PoVddP9/TMvwx5Zw7XgWHtaMxqPshCWlCNXF+ck9gHyoNoCGu5p
LdhdXna1dzHvEJPI8iomiTE6LyQkavEKobJTbgYYjn1QXHRytBjgEizYa0cpkaTWUeGTcbBRGd+Z
CanqEUUSZ4ES24BI12HcKZl1XOfqGkNgPV2TDeJEycEMdcKtNds4MMQiBP4aXLtSkycPjqfqcaUQ
Z5fqyHvyo29bMOokUTqbe8NH8IAWpAZg24q5oOkL1KDPCGjC8ZRvX4Ua48i9DncbgXL59H9HqfQL
i2tkhLnAF/Cc1858Ybl2DAAcdmjw6qhr/oAyvbOEBwftEQPF4nqAJ0XWM1IrqVXjolQRZGcXMRJC
Ax5Y5sVjlquiIduhZvPsEpLJWWFgIcskWm1geD/DxNgkMrkh1X6cSRvRmsMYT7iD89/aMaWIRw6g
4Z2yolAfJFuCvtquQlKGQYdqTyzy7KmpHI4hgxdTRbgDfUDFML4X5UPq4yGEazPV6ZEZ+e/jwJMx
lBGPu0OtbfVfsZnrLPvtvEPfRL3xqSGl6EBxTQfEbzf46Rtv24R2xQz6yvShFrMZ5f+MUZXGvI0k
TvrkTa3rvMDy6zkoYx8C7cNt20bOS9gWGmx6WlcOqvfI00v6S3OLKp36KsmMvQt+wktZq/o6rJYA
DPJtMJx2NXjjtsCP4EanA4vFNiJ8dxI2ma+SUrUWTeoXgE8r3TyKL9uu6+7YYimAAwoI1v9q8Aow
2eFOQGrmm2r1XAJhcFI9G0FO7OGvoVv40sNAC7OyD3w3CYYZNFQJgC0wdKvw0V41Q3PaU1WCZrXG
KZdNzfBXtN9uf0TS8J7xOBT1COzLG2DjfaRRS2b01VD+2x+0S6mh+t8UC6Qw2WLU4UfHm0gbudD6
3qsIPo//TXC7wV1xLPG0VyLOxi+tpVtZUaYZBRTd1egg9jTNVzi9yrtO/NmXOBY5gp5eGsENJA09
xZKG72btgtW/SWloVBH1Xotu2bdxaTLGmAGK7qW81rYLINysY2TWU0y1hLc0y74AcgLYeMzeo1xC
mCqaw4yJtjEhJkqwmX3osUav4a9bSyDNBWWYZibVlGm/d3QmoO+A0h78fjlUygNr+lR29giIfiA4
IiSNVktILpNr5VxCo4r+LyGffyiyZZXQwDN2eQp+WEvtT6CAbpRyFdiOMYXfLQVqUppgEnJ4gvvd
WNhm5EjjJ5onFiBZBSEtfwZLegnHtxBec/aV0zrXR4jbSwPB3/Vy3kiMQIEU+lrgbHip6ADuHkm+
Y3d8F5OBT0RHwNaPWysG3Jm/HrFyGDVdK7ie85OYTUSeF4c01yNlCAyzXhLcQXfATdLaiylcr3QQ
u7+ZZavgSeni+TDD0d5Hcu83yPiIhle6qZrGodIap0bXzh2236+YRSu1J2s0U4iRvY9TsD8QdQtG
8z8FmMzY5zOyek1VJ1rz1tTF/4G6Rgc0FdmM1vcYGHt99k+CtjaRCxUWREnNZebxBdKDBBWPqOR1
fuh9NhR+qmv+Yzrv1RPadhBs9G/o1K5UW+Pp2OEozyb+JpktrjlPEk9E+UZWZ0gcJfxry4pGWRFz
/C2TKmR0WWJyT4b5EiVIdav2TrZNw/S8kcgv+ao9YIBF2Cj1YB6nXp/6FMM4OabA028ukG3cvuZ2
VpVXJ6v/nXASX3KtgHdEoaLNxt+HM3H5mhgKuk+N2KbcYyFFzW8+8QrrWIbQf2qqbVS+Bc+MxqnJ
vdnkhRBCPxSLap92LLpwVqkGIeTQa4ahZiKNH7b0hKtcHKhgJlxOklUthVb0U4lR4EkBU1fbKu0t
q+4qJMi/334jXSGs2FCBz8TQjnF4AZWOuMPU3vcwp8TQnHQRrXv4JIfkCwgdjqV4bAOEdAIL2vh2
f9UABQZ9kSUti+BZiEYcB/e0DaRySFVML9DVATVEV/Ryrb0fUZyeTpbSVZgL+9T7aBGDrSjx7Lgh
PLCah9qhsdc5lDvFe4CGK+sFSNf6HzoswBEppUoOIt1GYh8UPfXgxR73xln7tVEnl6iCDHTbE286
sfA/NLayIfNrBNNLHd+uGBWKQ9ClnegI9tXSqAWH5NPDA6r/3+bhjJ8zwEtoZIgdVPpGCAouTHYx
pxOOCNeFad2E2sTtJ1wdE2cQCy5RWBUtuJ9POTpP7Q3HEsZ9Sw+pmbo2SULApnh37TYd4J988gAe
onaz28dFIgkX6EEEA3n+7SOl0BfyFRDrjpqYEtsG17e0N33H35qEzDrGzFJHnP63v72hsOvQXp+7
OchhUFnmSM2x+h+vbNurQUlKh5ucbdSsOg86RsIV0l5VK4G9ciZUkANX9S3jsBTvT1yBt+VzlYyU
fBv4Htr/G07k3eMGf5pFOBDP2KaZq2zTSGm3ZgzVJtl83DnIpOGC7byG3jtl8sAW6n2mlHp07ysE
9iMHbZdojWEWylmaF7gtozis+JZZHKSwuNq4SHkRExdPpBp4t9CDYgqFWYZAD/7pMLVSfIAevEzF
gmKBJTKAkfbDpKbkbqkj/+EVK6+eV1kCPH4+0jcwcZePZdRUqSuNrjYGk4SSaxObkIcuLUAuqPsO
gblExtMMfqdHvpdusuDdUrkqu3ZdTpfDBVHa2+y+m7GNnPcHEVS7RP9ikxK+1/Oxbz4peX8g7I0U
0N6a7jomEiUtHB8axfzZSQMldA1eklBfsRlMK2fleGvj7vnsQHchIBsr1cJOo3LmwxbZxydCN90F
qcHa44XZ2mAp5wqJBAt6Y31zB6HBMVVf470POc6HcaK7/p1nrzrWNvMaexphoabEUU5+fuT/Dthu
OQQOE18kziwK76JuRc6XHt7RkqJDQQw1902hlJkNp574v1RTRppFeT3O1TMNcihr5GV5o+RZDx0d
McSf26c5Bxw9kauuLfUieTKc0SI6+dBUEUHxtfOj0im1+cGJT61b7i33QyQcRlqTs9bc+wWdmQz2
uu1qr4JSXrSodx72c0LJE7o96LaaobiJKPd/ayXbpkLmnZPqjDHFjSFvaoKXXFSWduZoxZXRqQ/B
5JZsP9oi1mZFnVUTzsdi1eWxIFmHNyy18mvVTF1gT+qwExTdDHAUACMXrzKxZwVmDJQ8i3cBpvmz
/2Z8E+Gj7a7drsC8+m0SR1c03j6Q3gsgSSRVHHltDGF/YeFZVrR5PWYMwRViqaRYQH/0nwJ2nKZm
ep+7ZLVC6RxWTx33svp2CfEL0JasRATOgHyalwS6MRAbyb2QPYwpvxLEBZLUfM1cRCFdRyzueJtn
ePqIbZ+pAnWFQyi7lT3Y/0jjx17ALPUcyykO0LCyE3v2wUeAQc1CWigIl/CIluqwUf0Na54vyhnK
xKaaLmxYz5oqA8JV6QOQj/5sDfAS/yeYWxC3vYPyWuA1S8KtFtdhpqHPvmq7NjXOxPKC3sKa1hAK
Y3AzrDqZQC+Z2JIkBZX+1Am/Eyijxx+rIrmKNOEsAHaOiyVNdQ4FRQ9f2nuQC57TUGESuXEmleFm
7jIt2s2iK3GLVh7TNq5TwrEloqZlZIqxxsn3QmSeNzcwDUfffRI3KKomn/Uk43f8xkBEEPO5FzTQ
amrjfDXaTCK14+o7lQCnuBPNLe4TCQY5m/jcevv/+584B16RgBk3xeuEparXNtWRW4H/vu3G/kEf
DtYxPcS+ad6gDGg/OTniyJVntNP66oZCKWgbE2WBamsDE79OqwHe11jAF+sHuGMWIGhjyyUSOyZv
uu/EZrhUZ2EIMM9+bxQqPEtvqzxw8sioVaWb+BSFbtbOOa6P2JO+x8rkmWT+3I3ZkhJw29rHvBqx
Wgu9n1DiCr+ihvOhQgqWK1VRVfy1DBZfx9kyD2P3gu6/Ge4CC1bf6AAcViFJI0MFMUebbvCUQzMC
8EfJWFnbr12qRQP6c/XcU2zBXVZAsrnSepvzvRz+lx2MP95h/v7xG6FI+pL7f7AM70GwmrzlpQvH
RTWgJ+JsQxxvVt2YX9E/i+J3RO9mOVRqD7r9SXCz92nI9TXC68FtanMq0ACT/XE+tsZBHahiSwwW
NWP56qCFqDfxQ3R4ZfeE8czVgli1x/cnf0+01Hcz0ErKdpG8Imds92FsD/SO4YkWGPMyM48vnMsz
yudhXHeP2D55nIIDr0tIe1mug6bBTr5GWggW89NZH+EnGrq94pyCGvqyxBbkCw+gAO0zvmUp+RM2
Tvrv2J+0OKClNGMf0myUwsX/UcZD2UCgsVCN6kATHy0xw2QMnukytSeyrDxSBflLBdsz1td2mVcF
pj83T5glFsRyyycTF7XoNJdWtC1E6eBzvaE71ng94RMDEcq633IWk3kWJUdJjhM8LUHhYmTLMo/h
VttN8Sfq2HHGB9uWUDI2BPf7m8mZEpm7Le/QJhFD0sNsStcQO7y42zcmXzV+3w6dFDH2YIu1SFDv
7+TMn+sPubQ0LtopO9aJHrQBgpY8c0DjGRepYCSUuPd0BCX7R7CRuOrUWQD8xwU7RvDFrbTWZNTQ
1C3hlpTmRFf5kJaDpq1qzyNJfmLQKbT7OnFXIubBxf/xVsnywFtn7gADJFOHpdq56/C//zS71mAy
NoskPexG53UxnjGy5oRTNqwe9yaFk39NqkjRLuiZZ+7CHkb4HtrEYKrPBMnHp73sah1F4MaG7znx
8Aysdz769WGjiAla6PISOKaoiF0K00qLsT9gksgxaOfdGVBD0eyAu6orF365+iiPECte2+je624W
jn4YB4TUWVWjuZ7/uOyFrWN75+737JHszilapVuIkY5T7QvID3c5/MaLtFzgt1LzXvm3QAmbE3A6
9bWbN7dG4A7pSOUzuYDgXsCA9SPiyZkKll+e61/So/OR/ki5HBCwdHgEtT2gDftfJLjkLT/TMR/+
rMuM9xfCM+cG809uIzqduYIUJPzRzzoXq5lHc4kInCD32tXNxLWNnyy39BHFYrgzyvu+evSaM8yW
nQh63mv3PWfTSZ39aMMZ14IIQM1MK2n/kIO9BrHin8JPiarp4g347a0XduHUEMjKReE92lcOoqdK
+4Z1nX+9JQDaCdbT5Dzgx8JVRUlC30fdpWFfOZlBZuGoynBcNdlV2KxSetOp/NjWjwSSA9xbhBR8
g5DPpxBC3vPN/zM8j8zkEjAXUX/gv91zE/26Id0njZhBlm80jBudE0HYdSXNC0/bALqDJlHc1WNw
LkordEpErTIetoXNHEho5c7iqo8MSMzJBsHLW9zzxp/JSc5Ojh/Jlx9LpWBgBF56pzr/yNvtKak5
AiGeA0Zc+JF45w8Mw/psW8+SUQx3W83GkdWNcV0Mx5cpxrDEJ3drx7bR+DFPxrB+P5Q+YR/2fKsC
t8QRYbxGPRaW3q2wDdtXn/k1hA+3wd7rBvMRcaanVbg0kOkHy1lCVV5Kp6YYMoAlTah+ok2Wha5Q
TKM5AWZrjMm9BNei4IB5laGY9ZbPjZHxtiKM5xe8gbruppGYDCdK9C4GXQEMY6/e+bYGFnryn/NT
83fUykRy+ciBBVl+3bY/pXttPOAk7rx1sL0Lix7m+hoqi/0fTqacoRhU8YARZ6RW0GQOJCoHyA7K
nHYMYH1cvFJ/EMGx60XdRAJEF5X26UTxi1Rdr2CYs7x/qEtWCiNGNsagJhgkCcbhuMxJnr4Bl/q4
e4nSlZJhnHB7i80HZntaMnCsy1BzDg8m45cPDXo7pLaELaQNfKJazCnLq4wkDW/oWr9nkalEjx4K
uG7NCoMiQefoAbM5PO+koaEEV/II6tY6L9RC4+phc/D0bRi3e1uLUsR1aeK/WutOl/MryNTuND9U
OX6khHljpu1vHX0DY2I0DI9lCbgG1mQ4tK+Kortu3grdcSZWDxFiqJgngul/jbiFRqj3gomQ1NuA
YcAkGh1aiyjkNXW5WVd8pd0XfY1Guz98HHIU/nnQNGlYdfIeKrormMoHrsCvceFDPTQQm8PMokk/
4XCIwQw7r0P0CxljK7ZfUIWdSeE6c4Z8OK9Dht2PckRyQTgQtyKm6zNs8knLwTNR2pPGyRh26b/w
mAgMs5nL9KISQ/TqQITACJLvrrrMHNY+eHjzzM4Rv1nf+nlyKrcG934oF1ZmLELBWhJeJ6aIrn9m
wW0RHVySe5W8r27fiN/x4FyFM+EYzb6orGGN2t8HCtiAyXT1x+1wJ2evvNljGXGYL0YJ7XWG1nMh
1KUN3RBpvfrwU5XNKnEwnl0kvNWkkGB5B0iuxpFYJ+o8sbhsrQJdtfrOjORuveDADX803qBFD355
FMZP75ZFj/mGv4TkBUm1uR13BIr9GRf6Mc0h6zC6d7GQMLAd2qpc/K2kSW3Ulxxj6VjAcs5/rPeX
7UIFz0LseATIStxRTh1Y2+7c4ybDFKKecnzgwe8+q9BodziHKwfpAUUIEax4iXtCZrL1/LgSHs9X
hdAiFe3ye1z06CcN47ZePZOevP4to60y6GcENdVPRUY7+WRzi30CmvtZktyeIigx2zK2lmhAeZqi
SefXZZnMcqN92KXhULGSKc99AxBwjVEPWkNJydHi5CdgA75BmmKipQXrI8qMcL7OsdK7GwR8Hwji
dTZfBjn+s/j6BpRFHuXP4mqxEXAP7ZK5n4w+zNenmXf7DJZc1+zAruWfgjnCy8Wd3UIqRLvugSN6
sJhQ7XjTKQbKtd9Iari1js18sQq/WPSfN7tnzBY0j1NlUgZMHB8yZSZSbrXasztchrFF2MYF43iW
cQCv03vmcetCDrUlz8jNIgB2niK/lu/B5ILsY4DAM175L+MbSgEeGR6NFUwe/5QZUI2TWNfzuQ6w
ZQS6PMMWhApI2Hv8wiDlc6QU8GjKGxOE/0KEatR5kY4fJmpIhmeKmgaFiUQxddAFEaYo7iLMQy47
FzV1DIZQG+UPAVOOVwJQ+/WxXo8nokBwdZsFhODFpnDle7unlgod+bwl3tdel5hDgHLW8MGEivtP
CPwkEQFfANLlRN0xZ1XSDVMlYKCcieW7kuC6Og4b+YrqXhHZKtIGythjkcB7vh6y3Ur4TlpIVAer
qdBY45y9sIHiMYGGpOu1b3pq1m0+fhUiFfxU4qpM2I2x4C4d7GWkoENG+AgnBZiNxaDQjWRAZyj7
VoG8ViUG37/peeoTEYCRzLZ0J+CyzJEZ1ISaYHJuF7jkhAjNbWE2wIEAlytFOGkKqqfyq+Pp3qpM
Ir5Fs9+ex1JtsVjFxxbqbDr56Eo2McdxmZbBhoTHmDlQFvWhHC4ZzRpasRs7O+s2WCjAaYus/5fc
8dUbJgeBwA1zNQ7Bbd85rqJtIYBYwmHLUG5oBBbxK0yXb7w3/e3VSTUxH0yMGJQz1lA+1I8P4+UV
WsFxZOm50MVciE/9dSj+7tHWGyhfgPYMFzgytAvz89t9c4E0qh2MZMefL10oBIMq//keh81a0RGi
l8TwoF5ycXFzrhfbDhUe3cEcETOiq5Uyq2xuHN7cIq3KG8urJ2amfRVOgfhfTvkhalHXiQAPGNek
BAIZlCYwRAR3lLaZtrwoxhdaZhd7Nqh2lDQO8OzYwA3PVmOC0yzuoaYPerKJL30RxKd0O5RfdnQm
sELEjEGDAojwzcznvbJQ2utdfSDBMNjOxGNwSOj8P+sFu3xGYxwWZO98A9NJ+wl8PEfTccbo2mSJ
qX/AUcslWVA4Ezkycg/nWoof3ELglD4eg2zfYciNVI3/7q1aEj3A94Lsr0b/ePgoHyNCC6DUGsY8
IXCequ3PSSVQOwiw67LEu1e64Q9N+krm9NMUYkOBOUtYXV3Q2OvkKqEE/d8A+UaUXz5tUFG4ECTJ
MSvgFAzEjfX92QyqimVhMa0+sdawLz86+7FW/IiWdeVeO7dYHwJHj3v8eNqXQWPtQtvubBi2zlYU
Ou7YAiWaklh5CqJjPEN/jm3yly4a1AlYBgSmg1F3GXDYUIbVJ00lxhUTEmtK1G0FFfBK7JJUhVc3
cXmG6NdkANZMM8P324QJav3CbrVmWl6HEiyzRtgvw90STpCldj3l83H8HKrhFzKSWJCsr9ASRKuh
G9uuCK3u4CT+vwVA9IAnaZ8QtJvYU0r3sn0BP8tqBLMxfiOZPZU3FCmwRyLYAL88Emjpgn9VhVbC
BlOSdQjpvexLJ2F/75DkC6vlxpX9HbTbCJyPn7rdYSptqIo9qdyDeuGYyRtLbii1UxB5VkboS7KN
2k8DRsyS3HHU2gE+TdLHDc97zG+xn3lOuKcUO2CJjLhG2bvnO5+1/lGc1XA8IA77FjWkIhIEV3dJ
GuopVfUmWb5UQYMwW24hAUNKWaKnEQZ+VpXB3M7VJn47x0evThjv1DEpmqArmOEKMFis00fFPAx6
EjJ9n/dDFdZTpDYDNlIasrspqLZLIxKXXZ7uojV251h6NBFRK0b1Xq9KkjvYaxVZbXGZ92/Snba8
Xo09Zui+sI78vXgYg7cELEUTv/CVDPB5LwiiOmc013CM/OtEb0mg5SliWigN9enNVa8RnzLwczl+
JVlEcJC4EwYNCPwgIrEADtvMRDqydaoMDLuJBoAMca94zGL64nMNhVp79g7bt6sRfRnyCJCN/JpK
nyrJxLxc3ZAij+do3MmampL+fNVSBLSW7uT3Pz3zb+r3ulGWJ8/5T3i4hs7qUBh0Ey+zSJIvRxR9
A55u5MbdeQjmuVa9db4zx6J6pIO0YyxgJ+Ykai9SWIruekl0A9r0EPkO1tjivm9YQ2FcikAo0ULj
4TRmLkjDlL0uEWFiJgB7FNp9TUQ9BOQ7sPfFO/TJlXKpLSEMUOy/cv5oTnSjG6UU0QTvFS9Fezoy
Ojyrm7DphK1Nxl9/6FcoDggIh6mfu6hULpeypsQczec8YTI8x0iWJhkucjdjz76R7BAByHuH12yN
/xzGW1xktGyT8cBrLvxtvy0NeeFaL6iQVC95yeEqjy3lnb0Xb4Q9hf5HD2dkB/s1vLC9x4gK+W9e
xej6wGg4jZ7y7mYQTJtbTzfePEQWVTcquZfBc0R/rUAtAQJSB5wwYN5z49vJB7FrJ5CfHSdiZuua
af2CP3orIFgHqII2mt87olEVJJxjYvizoAbK8E4HQSsWPlrWjrj65Khu+ZkpVq7NHVK6CnbkPZqU
dOqiVqaHFr/xNAminHd9wxTKUYeIEFNJErq5mEofuqlz6LxGvT9J6It2NHGuFTXUBvizsTwztFoc
5+eDiE6QSL93A3tdSUASwyk/nUBFwVYBXERMjCvMQ0DVXhwaewubzhRQXNDamhg0Q8X/9aAlotOQ
Ii3gjkdILED+7YYb8A0zqVyDgWEk7A0tw+ILeACWZnvKtlTPiHTVUtz1grPYZTSOGh9J2WyOpqwf
JOMtg4tl2Oq6NajT3S0NYCmhS50QeKlcKs80fH5NzGqwv7SgUi9/3PKAYLhpa6E2ANO0X6x6rhp9
lqMmNqTzqm34PAwSA0PEWVTUZbAnXQJZDDMiutb9Q/e/ipswSLcQlt8KB4LOKDGTaIa6kezoyTaO
kXdIlHpBaGSCCqi+bo1LECyLEEI9v2w8X5XJNl950AT0Yx9WqyoryAQ41va8XWAWcCu4imPgV+5W
VsnD8KFNkVUrhQieYzo2VvPk/cBRX1mAdz6dmf7z6IfLCd6pZIt4YpVfvxz+BkEiRuHfLZ7bo4yw
BRCrNNZHW+jkGYfphXsU3O+IoJMt1D+QEYIPxdEHEuIv/843/+tSX66dM5urI/ejhoKPTFGbg4VE
6t9D6IugGTFI9wusuddru4bAjHMNGlLFotaA4za8oAMI5OMeMbqmXPwXk6yc+jFeGfeTEKzveTEZ
HNGIVm6bBaBRaN6qSj3ZcgNKz6AriWNTn2Ci+tZlApjXXXb5+HX1vvivJ3+n17poaE1sQ6D7E2iU
vs/ScXVAITMHgUJ97yLijypX14vHBvYVWoAxvwQA9ec+T1mhv+YpwzinMYUAaUdOs4OiZVm7vXdS
JoDvPC6buYU9UATaucV4xYEsYUe9eOIL+4OQuZUh0CHueb2baTHHhx+mhacrtc2D89sWDvPL5+wK
W0GJdTZSRy93pT1WlFdmqo4sIdPMdqRRbZ+TQ7xzhJU2FkFuiZ5YFLZX4AQ1I+qzx0safRHEKZJY
i7CNNpDR6WHlvvFTPPJvpuv8t7Fc5kzES+G9D3TGdNKa6J/G1VFOH8HNuNZGmbgRPbxhh+X9bQGy
MXB9w1nBG4ZHFDmJhvziRjjsLAfJ1ezVOn62U9jtC39OhVL7ChLgI6pIk1qP5t3CK/ZCE1RqOl3e
4LUzjGFDmddGIhALou+a6Mih1nzHKe2SSeaYVqkrP977hzj23nsnzgW/D8RvvFPNxVMCgAHN94P2
uR8MRAkVnXF/wRRurzYX+KhMyiujxY2MRKMRTv0IDF/5IHLANxbwal/KwbdIfY0Qfnmz7p6hLHKW
dNsyztklKpa0hfI08jshNBq/Io0041gtJ7ApZHcyMZpLdJJT5CnCanIr2jcAFTL9O9NYdhvtW8XD
CgrkIf5GRsqWcZQWJpFnTY3wd/s3RVb7kM5s2i/8aDTHd4SgAdNKK22DOi0eXhWXJ7z7afEXe0Lk
0dcMx1FwGABYBiIPNTybqSRgFKuOYft6BKyVQMrGQneXoy/vgshgWWdfzPATwOn+Ylx77nRG8pt6
yPyFEQKMVMCU7TOGi7kAjEksDz/GTCa8jhnoA/14EXRpku/nb9oiGE0EABXIx7vmaMF2SI3Mt2Zq
G5nCC2r16zXIQ4wwSY1Z+JCiu+PjGpGFBPeLKLh/Tf57qAW6mcc5AM4SVKl2glz1Le9I3IzlAEK3
WyKOio0ZI3sJIuI0BY82vUC9SwIQhot3ExKnwXyxpdWl1yoz0g0VGWpPMehk8qPjERALnoEa5YY4
06o7VGiUpTA+uC3C2lkkmonBZapg0JEcyNQjy/cFerhw2ZAgcumDNVH9PgxLildspfoAQzrFjLYY
P0zTR3r7EjjDv5ioBzWKK0LA6kxRXspiBmhMqezuSrMYILlMRwg4ApSKIagyCVJXond24ypOgbrL
XwQ3Ecacdii7ep4BdVgnWv4udtltukb9SXsMiXeKu5kDBE0puPPqfCxrYR7qnOXAk5fK9XbtQn88
oTOaP1VhDHrB1Qo6XlKwuOkT5qfx+HCiXnt5ezNFuFGNSyt8xxpT89+7ac+bETyDlwxvqm/H5TFq
t4E89UJoUAS2pllS6UCwfAdUPWgDoF58h/+EAwdldDVFMrJQ75yitbpPzRBITQaG5ZQ5l8FYoiZh
lEaLUg7/jIR09gmmLVPT0jLs4HVlq6oTiwFy3yB9qMHmj54OzbV2CHNFJ6BoM3AI1rF8TXNYgKeO
nuiAkIQOvDzR43kPVtvztvbt4qHW/0fTwTraukOO2DZeHvlm5M6zodKHhlqU44QHcW3UYT+HQH9G
UXAJjgPflzfocBQlOdWagIJPWK5+C0OAnCgFJRdrS0OdEJmjhpwrRAJM40VtGAtrdbJwQfiJGcdj
UrAT01hRD6+yvi+DgTxpTuoNEi0Jxv5Qk6aeU1njkg6+gTNbPvcMnQdxsoUZNC3f+RbMRYzU+fag
G+iCHNthsEYXLu0emtBwe1maDGVFaXD4MCiJ2xeBb6brJ95SyLLtLMTSvtcf4Vpw8a1y+BymwGNe
cLISBGB4Phaojk5zlrOq7yzPdJcyPIgjam5auicxX13ae/iLFIrm1IA9DrsK/JXEsRCjGj09rBeh
QdaV7kmyW/IrAQWHRrmS9S1d64lw0PiCSCd9CRzOIvzxCK3eNByhcNwVbbyils5OFu4vyq632Noq
IOp0sFN0TOKP9tzGbXSCzDxg14bV9ryjSWWDnIR4a+4Nf99ZRr+mpuwjabgtdUTb0FzgpVAqV6DL
Kd5OvEtSlmWzrKVN7dOAs2XVhl3YFUkLIPnBV+eoQ2TkEpnQUY6yHm/86joQc+TbxxVbn88in3fP
hOHS2VL9wJbASPcvp7vO+iqvdNkE2l+zXiY9bkJXASiNQ18Ex1UQsavnO+VqEI7IJ73v1jfXSeJk
aymq0Flroi63EAIGQig4DDrpiaF9wbC60H+pwLxjU/YamtcL6Q3XwbD62hPDnHahnoWE8X2ud6e/
aRFjnkuBWQtJS34WzoTz0LgZA3rIiw5fuAz999AcR4nw9LlL1HJ6xmxVnt5BOP3Fn8K0Q/Ah76fv
XUlYHtn69JDr33LDi9l1BJfJgswwYHi/U3cH9I2lgqQOYEEX0tBxuXM8UOrDI55iq1W22rC09Ys4
RFUuO44j47n1iTBGBpr0+cujhsgAFsAOXu5lO/SSjXPbdfAfdJaeicsyun4buzAqrRBQC9uwFeZC
5T1P7JcfXke0jhqD5xp2pGpiXmsDsjFsCZLouEmgIveeMZWPDxLEQIi9D7OQ1ShBU59ksixkZ2lZ
4gUz4TsauFNsfMCFv/9kuOoQJrdMYvHT78xRmdweZCiUfWVB86CJFmd23B/7VpRbONTPmxryHRuD
8JMjwAQifXro+PMTFxBRAmrW3FpcmPuYHjba6tfsqbvnvhn+BOaaIk91dabKbdcyNkSisNB17UG1
Z6qcNcQpOj725hDxLlP7HpGjUKFfkG9Rv4CzmVIXZEQrdNHNPMW7WhPxuoESygdoRWpr4sOw/rOX
1PnRcNRNcaF/TR0pb7pDoBteTvfCuahJbTHzFVI71bpk5jnGvc1J7QeeCukZFbFoY6k8crZlNm8u
wJDVQCfIteSDvOI/MMEIJHwpDidlcg0vsq+ggyUxo1Btjsyls5BVo9AZ/dpfF3o+PEMR1bJruKDH
MLRBxswZlIbizGsi15PRfzsDFalvhlISl8zkI7/oBPF1IHY9l+qUjDjj+rSn1hKONZvi/TQwNh0r
xgrcYIaDbBpfjcJktEMmsz+UidShVkml8Olvb6sjLUqK+A1hkcX8o4OdpYBISAFvTjOdHThWQ1aq
iunNt42H96jrzU++oOpSga94HMpAfj8URkjFSi4sOskC0auav2clszwiFnStRe2s6ykKJ2czpWAr
UX5w7oNJ2M6xrN951B0Q4kk/tjApz1mTi9NsrkhvjaW7uhZfPAhpuPCOZcLEWkLxKuFXnQhl0WXY
6P1q//k5mz9R20aURBDp7LywzPs15cL4L5Kgj7EWlAc/r3Q+4GYodPFDXKbPFw1/QneYtoUq6Y+Q
EoiP1dIJHQxj2B245FdYA4hpJKESOiItpynJjpLd4/A9/iawT/4snU5wkhi5NASxcjnJ+0y7qHup
b1gfZPnA5mQ1RgKh2aVC8LEnZHIPWXkrZGEC60eEFTVapYjQZS8Jf4FmzLaNS2mhaDzmqkc/f4gx
UMt4cIa8eiHcfyplF7auLJ52oxphSNCrH4aG/oDbE6MB2rNWLoyCh9S4TpItDIggn5gMild35BVv
yT0i0A+UILb7Z3aM4v2+6GZPt+vPjvyrz2YW6aHL6UdLv2kFxJvFbdoh++6Qcho7E1AjAmTmqaoR
XlulSpNTn7kaHsSv5AuyloTYmEisl3V6c5+tRf5ANXUJFmZchPzJZcqaY0z6bkMRanMkx206jnTb
UBb3Dp6Dn+zOaHBxb7iZe7iZ29zaid6tQYyqCwmjQvw7tUjwZwh0PSII16j4yKvXckDfizmfwYJZ
kk4D1uH5+sm88G4fsrvTay4cxCyYh8sjMcKwlL+tA90eVgPymz6BWrHA17fOQiuQ7/aLlxfpWHIo
kKwVNV6p0HhaLARuMKpRfvhFvEkUCNM3RfqgMOHeCyyRG3SGYFwWPWZw8+9ZxfY0v4QrFtArK8+b
ZP10+zM7fLniWXIRF19A/QBk0s/1XUe9Sc5HEc4v3/qEnAUHp+hi0luRpHHgGWiDZzJ3v9KA1uB4
NMLQHTvuRNWta5eG/bc4clJMDSL/jUU5fUh6b/evSgLyzoPJZ/qBXi5BRsPGqNsd2cp+oGkFZ0y/
Uy3x9MceU8zLNHGClQH5PCM8jkOS0KwBCGi4RSXKVXaWnOOFIB/e5pqIwjEp3RRZTLD1qAJu9aL1
qsUs2nnaFlJTknJRcqo+tsSxO/3JaHReMpVoNU51i8pm0lhDLm9v+TM19XCGiSvEVUkNEmMaxi2J
6u+VgF4rlGltOjdtyu9VAWzAkZTD1lV5Boyd1ajQXGnTFQ7VciYx3ISCAI+QRSRtzgh3W/c+5Yob
QB50Vax6D1MSXRQ6araIdBjeEDNJ3OMzdheM1fMbW/krtKErH+2eoHK2GEhmGFEgwEikiSuvainV
5d1h6VpClUpXsiBXtWISPMjNiSpVqBXBwyhuKyDkVxk3BwiT2m4xO2Z4h2ASQcag2dkeosd87fVc
qLNtkULDqnm+NIwxQHV+0rReEBs3RTXn6n7Y5HiHDyZ+QgexkHMAXjiY7q1j76Bj6uLSdVcNnb1M
srCiRUvg+YnFQg4PYH0pHE6iyb0557fkHfZEPQ1EM9OFcWXhccZtzQ4X9OkwWo5zgFdhMvTz6D82
HCVhHI0A0wrU03Gg4XZc8j5JZxx2hE0sDQCZ6dgdq/jl0gXZcIzJe3dLgm/flaYrcXE5IuWbAxp/
sYX423uTaXvBpVIDGgBdoccSpqUudTpt6+i+yweMFSRj9mfv+Rkh8QEeI1OUzKA+s0Ed/FHMhqrL
Dcb2TJ6443jC3RrTcXppn82BP6qGjFh8fbTo8hzqZTQBo38qcEVb7mygCNOYKwvLRvZWS4kGKpls
4T8+v6U69RCN3MgwmO7vPiNBAmUyedtRRHjbOGriVfuSEuNF/xYFlbZcj64/int3UmrO4UidksMX
PbzZoCymqCFaB0nCIUIf/YmADLthLXAiXTrnFW5OuWWIBgIKjinxTc12Nb79bLbW7yC07FxXxmk5
Ts6xRAr7X0sUzi1IbQF9qXSitxT44V+ZHlHv44CTb515imZoynNes8Vuv/6QQ1Q1KRy0cUflTKO7
SUVkQRuBIPy5NZj46RnEZLIE+l9XWu3s87s+86A35NhT1THd178ebZ+Sg+3UszwuS+s+l4InCz4P
0l7J2ktk/fSFIqnbOwJZbrZ4oNDJmUn1R2ldPkxGnDnoAAz9UYG2Vutle6HVwWW2e1VvZJYIvAP2
VBT1IFg/wvFghZPShl7NIQt/63LRoARJIbdiauIt2Hxxp0sj9lcQW3QcDKRAHv7I1rkwPun+veSX
dC3hgxoD1F4tC0/DL1NHkW3rHXJawBAVxrUgKrLifyY6xg33uGykGLbS9hcZYmbYYwzjZBXi2yqz
AWLaP5uPXBrb0B6rt2U8f4whWQRpvoxK15Q4+vCtINaBBRKVtOyxOuSTEid0HTCZP0QK/SZeYONw
PGDxeJNnWT9O8Ddb5NX8QlotBi8yEruraZ+ODAskEA2paqk71+kimJShSDQ6Kb9mymPuat84u98K
r2S2gSGex4yWJr3CxCssd9dBKD4RscLHw8xu7LaAPF/DbOPg/2L2rb+t1HvZ43/eb5B9J0yfDvpe
PywsX+sjUYeFzWQSWB+t1+/MvX5iiUuI1ezerBY3O8K5Fx7+Y6q88Bv8xYa/uoPxAJK261NODApe
IgAtLr1lc3HgRIvP8UKVCkr2lU4/3IVuCcmolkrMn9Nkad3+0ogcIxcRjJD531wq9s6gmOzIM2Ue
IFhT/NaaGfCOucCB9CrsziPMaonkm5qyMZVwtnPOwIicqJyD9Ez6my79qajPfdNkOc69hkyt09Gl
UgWnWAPqUP242RDqtve4m5jMM4fdXc5vRJ02EmnfXEacF7cT1G6IVZ4BLAjDhThMzCccJfRM9CZ8
oGcxU6Iwa3H/3zw2rfgke0gwlF/IU8aQZ/trlxCDEXuAxjzldL2sBLUUaQdYn93l3HrhU92/irNN
s5OVfiQ3AmSQ2/ssdyt2ix77Pcgr01gDTtYHlr0x9aPglY10Aq0lY0fUt597qLa1/sJnwHprWwZM
m57L+OXFmjfTfWWhKUWtOnubMb6kisV4T9y2ZP/EuF/TgDBbNHw+0XhW7BMXORiwF5XBO6FOTtRL
4cQOY9cCkocE7QXyn7H+VToUe3mPbSBWh/v3bo0eGacMVkT/BDoKtxCNdOWHQ9s25XY/k4YHmIXw
VN7KqdBg+scESfzrVMcBu1sye+9hz/bMuj+2DKBNXza4aZkMM15tKGg0kLp3PKMkELKFrJ5RBugQ
03CPUr754XShj06QPKwv2yGs348EVFDPwTky3h1QNf4Ur34Lp00UjXx6WacK1sRBur/RQ80u3O0L
1pl/eqKFzIoJl3HT1A99bFbf8rOcJKmK2jQXK+3u2SQpykyEunBkoF2o9RM9i3FCcZGyahtm2TMV
96/uKo2+4KIDlxWpKI6HbI8hwGq5EoHny7jI0zPDSuzGxpKD6Q7uhBRoCZ8Br2E6fEImAunf7RS+
CuLP1aqPHKlorSeR/HxO4hsFbOnWBjZE30b2c1GuhTOu19dP0/Lfv2ot/kcsNrSDxy23Ak6jyqnH
WiwYGXKGE39XQqB/pu6qstY7keqPytREV+1k9D3fgcSCHJBaO4EFt7IzCQszUiz6/isKXmWnqfy9
mQQ1cimEFSKAqbE5gAXwA6Ms6GGe8tCy86WqDAj9E3zvGvJh3NYeOqhxamM8MKs63U/JYRokDzAT
am4RCDehvH+RN+CuetPonHgmbuLDVtFyDgFGMc8Zm/1lMLmKXLciPnmlQtDkEYGQfr9gLeSFL1hL
nT8I56iDDZHG08p/9bts7M8x0HAzV7LMkGLcjRYjmI8XIqQoUDlDCMNk8J47/UL5s+GiPbQlgBWw
ALUlkJkcUVqr932ZCoNexmCI56+TeCsfxTaPCO8nTHS9ajIfqPFq1RIgAMIzT/PSJ4pWQbHrF0LV
fLbXzps31JCqhxGZnEprwIIVqlaFedQHpOyItBjex6jJTwL9FJU3BJMp6fjLLaqZQ7eMGLfhX3Nn
yzKWLwWqfDTEZveOJClYHwTsamDthziLtqziWF+/3UwBa15W5IUTfhM16GN5+O2p0adVb9B4zq9K
iJjclrFEuTq52BDsDdX0JCxGrSQPz4Fyk4i4LrIquq3ADeZ7XWWdnB/+8BccidyIRAXyNd+HLQy+
Gd2lvbsWQ2hRC2Sibsm7nqSz7oAZ+NhSycDgJF2k9+/xHQeHA4opFZ0S6K19oZ4VuTdOCjuJ8Ouv
WON0yI1t9pZLhN6BYav/TfkMYAiyjZqE6s2Run551Cz+QsjFtEAyWEE5oom9XSlq64wqZege9VBb
u/AjJX78tKmfwqs5Aup7RTf2C/Qq4yY+s+9oUC3TY0iDyDJh80oB+c5w2n0FJa7OO8LRcbgtILjl
K8lxxM/3jx4BaPu57nSnrE3PKS3xt1h/KExaKchY/SPLjYEO+k4lMANqwp015te5BeEDfXIyxarW
YIs+0fo7twsHQGJ4r1qtgqNuFp+Qrjc5bN+MMdy4sI6pFDTIb0bB8/vNPlFvNLkMr9iXLIqV9ZMm
e5Dp2qYH4yjQmgqe+A7WyWMgBs/tCUUTrmOqWdKEjr6fkZgO8HQqGJZqsNTrFkJ9kszgN6FUwPOn
phpEHqqt3q2iYGoTvRowotFQDW7ziQ2Kp31MuwhiOYW+FpeuD5n6qzxZwKaAKkfnaAHQ9/DCxQFW
1xX1Fqk9D5bUYGmSq8h1kzVhYoEjmgIHez68aNk65/YttMSPsMoqC8qlvJ3mhlT/Nt6jDkMGyWEd
C9YMv5r0H5Hn7pIey7nAo59FlER2qWezIQVqH1O/+e12YMv42HyWDdrDUVoK/qR6KO881EdZx7MU
stHSQqoQSD+70SaqYKfKqqv8LS8L+jVSnwZtuJmmQUnUJj62mNsehiH8j8t+DCbnHto5tNr7M/B/
ovXpzredzM4s8UlWQpGJsjAv2EctDeb0uED8561mxQzM6KC0hGA1rQcqgQx4ptPM6gFbDuuTfXvQ
Jmxq2h82AJ5/ZGZITtueRjt8KmkQwwERkGERDX73v0ZpuQmnjI/aoq48mW2YyzZAEBnsL6mpJcAt
XnjS+SY37Vqr3LlI9Rn5oV2faTqNxqG6QDqAYxiWaxcodmfIsRNjYd3kxJ/PjWWeXfrlV/2QO1n/
PBCZoZYc1d7Xt9DSLY3TtIFt+8zPNeUE+1EkbSIrq60mTpsSGk03Rs9dn6VTuSbrdV0TcQnlMEZP
74DyVoKljHWEokrBi1s2PhCKdfoW6aWHqz5QFWey5QjYVo2vzsi2taVoiVAIpFPuZG5gA1sOfcwO
9o1JgXc3yrdy1E/j+jItKmPlxOe6Lb9+5aXvYxrtm0XX8vEt5FcTzgScYWT1wqRwRDye6yKqLCiC
ZMGLJL+1l2CdrnWaWW1TBsp9pHHxTz2thLJOb19HA35Lp+HVJ5IsZE0zqxFANu1peu7EYkBra1sC
ktJEum+ykqQA/nbLA7k4C1LuWq+1/LRBQrPxQdQgkRzvfgoKxT/7Rei5eiUIxrjOkgpc9ituDbgW
WTvi1Y8kU6ID+9cy2/bIeikyHKz0pUDnpCHfLK9puTci8ph29iW82LhLOXKjCBihYyHjIk1rkxat
lNgk/mmIQiK76JG6UQkIEgcUyMYrSZrBW4FJXcDFcPxeJn7bBZyyhEORACxuyfwd5VDghU0onZ6h
33z9JkVrDwmac9gPgSHeS1pt001dOZpDCZowI/t/le9qaxhBMNSrxyx2cgCAC8u5Jf6+q+3dcNS9
FdhOwVDN5RaIQGIi2ZKcbRU0pkF18Wl7/WdEzLNeumq0aUt4krD5c6kn9PDEz5gf4Ze8Bzj4yaNB
gKBDKl8ZwvXeQ2mV0JI1JGUtgaQhppOEGO16hG3Mi4fndAYd32qLjgcVkWa1vrCXESwTWzNsxSHz
70Q4U6wuo3IWLjArwLdXcYqVY2vPCEw9tuoVBEgvWlJDd/7OTASa+5ZB9hmAYvHCUb6hyaBHdzk5
UNAaXqatIpebGl0X9h35ppps0+C9EzutURoXWndmj9gEBKqX52okSIfc7Df9SQDuc0OupYygvejG
Az0NypkSsPJmrM5Nm31DxgDJIkvvhfqYk/tNOSjvataOhGs+w3F9rg0bVi17o6gQXkQ6wg6tG3gj
sHz3J0t887gkfriDhaTdjndzFEubK3AJmCGrLfY2ajaUXH50lGBIReZjFT9e/8LKgnSMjQlH+/Sh
u9tZv/3/NqHgUIuzJPWWOTLWdE0Rtdd+OO3xT+KtGJkr3DPVQtUXnbpQPnkQA+eWYrbqSPIQ9a6J
rHdzN9CYgsrDo45EHKkPc+IkBa1t9lEj2hH0jRLuRiEHYYBhQ3weEPtbaf8H29B+RJb3K6GmNmBR
YBnbxVtyhdt+WdsKAj0qN8tBz2Ru3d5uHVTuruUNBa38vU7DzreSPg5A0rnqYeDFhMBoil5fVZBD
QmzbcoEaXxM4PTzvKIE3VEKHqyUCzXAcmdDlQrRspZt83w/ZvUIBiEympQ98XOo1I0Bcys7ctU4I
nYRq30wUUiWiaMe1Kqj+R9L2A80WgEm+PntLElhFb2MyHrxiErT8EaMr5xJ2UZI2TL4qU4g/AneV
hbhepViHUzplILjdtORBTYUZuhxX+HtYwIo4qO2gccQuF2zlsNe3jBLR5S8c9g3n4J5gNrSxFQpd
AKv0TKfLbhDYGnHZaJHzIHgpJoFU8BKR2utEuilcuI/rXkheKZeKi10UnLAG6bJNSYG8HrmhfGY6
oP+JSK8Qw/8wQ+Dr15ELjL1NOtFlPJPYej1IKyxi5qTy4PlUn5nhgAqkP9bvyKc1scfSqIFzUzul
NjdWxXDuTgnpoZH5t0Q8e0qX+pM2ah8Fdc+dNlzYKJ3aZPEKqvcbCwyurFfhLKFQByTajj1UZw8N
KyFMsuVn2/y8+Lonnw9gIb0FraVdnKJbVYLHRjxEi7YqBtzSQHx9k0fjouQ06I9uYl2YZsaCeCcr
MWbpbM2wn4rI3iMlHHAyJkWgtRpBLuSrvBc338OUS3hHPkgk8AwMqi6EUR19JKS+hZfO71OzZ5J8
UYS6veEcbZhg6muuZcTsTLh4wB2htQeJpphEKjXKMY9gdi38vrylqmd41XXqXXA60nT0hQ3mwPOz
5J5KO8GwIU/JiXUm9vcvYY3vx+oGMBCjlBtFi/XQR5Xa6cnxNNnFABOEkNLb+sBAIybaFQTvi0FM
CJkD0tuUpJkqINhvBWSH+aPSXV6JdNXVJ6xWcAj0AqLKkBQK7qbkdRZokb93bwtvUkXbQDURtxFl
7faG9ajB/UoL4UGhRjz3nWlkA1yWbN3z4bPfdkYyJvdt9rQm2E26EaV/Sdg3EMn9SnYXONgJXEQ0
1LMWr5/pu4oukGFK++gXePH1yYPqXC0Iz56MPkDBuvVvPOBJ/j/wFJReyh+E+HJGihjyGt2xutnf
777dAARVoRB7UiDRUJ3VURNR5VoMGDI2ZZNe4jW+KfTS3DX5eTvroQnJCWXTZ25P7QgBhITpMOof
UeFUml3n92ABGJiNRM7FL9/Ru7XWe5IdaZ9lE7yqC+k8w38YOQyY2yF3R6g2H4ub9YGQDmqDPxDj
S0M9yEtRci8D0VxRqY5id2Q2I4Zyfael+J1t+VWRsOPeVA1WCQMw/n6O0AgNDJCBAMy1XIYp8hBl
6JTjwqJz1XSmED+8iVjlztbo9B8Eq7y45TkUwnX3ocpv9Qn77xsvgRfHfoHsK5W8vXD4W9nOkrrJ
L/41b3FwLXi7RjLwoFWogSKD33N03m3jzje0UfuTDvfteqyjX5dvzPMlvJZJCgrzGYGTV0KJ7UU5
ueTvn2oKUOH4RzygyzZH1CV5ooF0F6odA86zH2ERiOzd8a3SFB4QHF+5ljj0mUllWuIW/wQ2MyOZ
LvkQdhDB0c633OG3SnBqJtRestN/+TePbyuGQxbteq839ZybILnM/7Fe52Zo3EcKk512cdzHWUQ6
BhuE1nZ+bgBMRMf+LKtkGHlxdzqHzP5+YlcFA9L0ypqdr5t5nU1yU/XKRzZfbXH9in7L/FUyo04Z
n8YraPlHzglQlz3bY4u3mmr89MTKN4c7AaNfDhuTOH74Oit248yeSONbzDR6m5HoEp/iBTY30a5H
/RAjfmJcGusN9k+sD0Lsatn9d0xGVGPnrBcjl/Z7msY5QODEb8J+DciNzZVVU3UsXCBgjQjtJ69g
lW/NUYsfHDLgrVHPrEz6h4LriFS6unC7srDo/avSp/x1V1xaVJu3e8GNxvYh9pjeLMbvAx3Mg/fb
muvolJ+JsFwSS6KSaN0DVE3QfXKLXa68BxG7J3dkuncxGVVbn7BLKLEygafvAtEhmIEJxd0aHqDl
IvugtZX/qll7HKuxM92floyxifFOmZRalClzo1Eok2jYajybUXVnvTzZCxvZY4kDL14ZB7zTXPv4
42BrWDufpMRF9PUUD8sDhZ90terVMu71nemKawHiEuQFSLX+GTjU37p1o1/IeGPVzCq4lYjMhdql
3Y+/sZeZg0SCKf7siYl/Y1RSr6BfhGbxoS8z5H6tqrBheYOzm9zgwSevWsQwwqEpLYM6bo+FVP3C
jwPBZm093EDTUOdUZohBCZYt1xqIkLEsJXG6HVs01BkAEXD7cuu7SZuHHq27T7dH9hQYllNvzZus
JvWXIfDm2ghTHdhBajkTe0ZJMxOHYDPQzGviB2tdD42Gl68sPghVrvHU4o0xdd+Hc1HPSupkes3Y
bI4YdpbtrLJqVxpUY2uMeJIEH6KI5pfISkxKlNmxvzTOqKxvHrC4Vpa7WjOzYGHxJsWA/RMKq+Zj
588Bt5PHgevFJTi8llEzdOy6rm6QmUGw6MIxoo7nARPT+MdjRhs8rlUi9ZJsL/ftbCQAOLJXF1F/
NAHEf5iR5cZ5Yx6MHCL4NQviI8E87gwvFc1WQAdu1AQJTS7iKWteth8ujcdsWAQ4tt63kqfMLBIE
Pn7ekCZNV7IJv9xJ6MzTnkXJ5fE4pGwt0elnZ7By/U9Jre0BXBjQBTHV08agI+CMBF7Fru6JJ4kj
c1wuu0F0DDfzhTw+h0nRur8DGsAAKPrpDsdc5Go1Q/5p1yuLpLQDzO+9X1O0GM51+r1PyXFAsQhJ
uGDrdkdke45KABcYv/20E76ocXDkgl7RNQMe9vnQxxNWS44NSf5qYzzgQ4Xn2cgXPtfbqpEMoVvu
aT63No83wgeh73idrM8QhdSBAsTYYptEG7ROlOOo8ESjSurSvHJhN7Y77p4yDe6BRA5yREJp5Uo+
34R3vIJ6TfJ/g7mTlpevWUbq6L+CQuZS1A12h0AHsWeHRigE8zXWC5LhcvD8vvkPvBUaIaSrmNxb
E+JEK6XV1EyQ6LNPl8+a1hC09ua+CpyddGXJBGLQszpgXYm2r5CVSkipXLwAMsClkdTggnlXOOUI
JlYzjnmSEpu37BLWMKRxtCYX4MSqMcvGYiTofx1j7bjfYYUPUA1GvEIti3ag0GLDh+AvHcz46/tW
vPs5bBCK8YjHQ6whZyOap5mCEv1pS9N+MznT8KghQp7FjSHae0U3TW7OfNkOXyYhQtF55qi5wG/V
/TjKV9dH4DvZansi87Y9PnZacY7K51MQrVD5pka1XeNyiVFXAeBaU/b77W7JwdChvBQ8vW8+XtML
nD9D/Rlr9TQ2aPwO573F9ZDIiVB7clxqXkpCZHQe6uBqrkWzt73u2geQpJnk0h3Nqj6nlCeNb1SA
hrIdzVY6zSbv8qbrTCGOiP3YnBd2BLVqzPc1EUxAnmPi1ZF+KTx55Df9oCHWmMYcfwTbL/9D56Dv
t1PyFvm9+qVma0RUEEMrjcYvUZi6x5zfMQEt4LK6KFO9ZN2aO5vrGFQTriM842hpAWo/N0qFuqYZ
1tAUz9Gm8bdoCn41QdQ8xvetZhsqOjrjTO+WXhf3oHJKUR5adWJvYTQVwTCL6O6KRj4TU2GB5NRB
GC0LqZl+7B0ewrnEKjlAoxFiat8hH7+/chZfzx+eQSP7fZEtA3HvUt8EbGAMowEvcvM2BHcDqSP8
JhocjT0aml9WKBIyqgsbXUD/B/7zTWNAPYhPQJecH62iQ8FyUyYqaFseD3a/iLVTxKUSs+ONGmsY
jnhmfip9gah7Jod2OIKFt9RZHWCcyPacglVCgu8JgOaf2N1y1gihp4oB51Z6WuFzkGEiSxjKndw1
YWw01STfF+31p/zeIJUrxu2HvTJpLzR+71yZUODo/Ix8dt+L/0U0EhWP6Px4Kn08gQz51UePlofW
GC4Ea2MkkLjkRD9YBePVl81EgTC/cqJP8MzI7n23lmtT0zGK0pIkHTVhpzqmlI6dUMTi9/HES6dg
UitAy/5AramLkHWoaUNmk75MuIuk9wS2tSNLUnbJWIhKZDbLcdeTnOThLzh8y+WThwCxzlLDUpCX
DfLC7+CzmtXWwI5OV/7UXMPj3v6IGyvBdFhoPAk5UyqE1CBL1qIHfxHClnXzPQYsOmJpUfQiptzO
jWFz2B61HfTxwRNleN8b9tPj676gfVsGr7TVCFVVK7BKazHuBuOpRtPudaPl9raQU6Hqg1ohEfvt
LsNvtSl0T6H+J0JdgFD99d8jtJLiU5nvuq6qFe0Zx1gjEBo9fqzMYCDqnA4jl5YtF3wM9wj2u3n8
KFjqbk3uiII9oup+JFerDKNEl87Y3bJSDOwYQbaqn418G6zpBigBfcbOqMGHqwEX6H8vY+muEv8z
fT+BoPc/wyNcN9R6Xs9jvls20F1FabW4hqpqhoVGRH5ggEM61odQZ5fG9ZxFZ9m4pC+3b8aLX74i
zjIchmxLEgPLrBr4cANGi7crqlANFR2MLzwGnDWzZ97VnwdrWcPsi+4T92V+NCH7oNGo1CvVBL1h
SMzxYIZ4buTL8OhY1FYyXffFWH46QQhB4AjTtLDgo5GLZm8Mmfa2t/EjVo9czZaZXLmlrMp3JWnF
hChsubqlWfVOy1zsrD2ZqGUnLv4R66ZwqvXbloid5gC1FFdABRXF+znKtEoyL2eK1oqYWw1tb/T/
tBX6l+H689YfhkMRcMpg2kSSoIBFYdhQ2L0F16kuUCxxGpkld0f58jCqF765F6LgwCzoSX/YSxEQ
rG75uLOMtvkhgLNvOBR4Xd7kqVIgNx601TObKHjbtXzzAu3jfHn09ZhGyHNuozVShuwfD+SMYHC4
PuGFqFvFsIRSBwo5mZWp5NYg4bJe6pRzqPn9WuZW3Qf5FTlbOUY1Ev3O2HjwMfCHXklOxYMT6wY9
NSZPfMhGa5NjHyb7eSPBKHTXgHNoH/RX1PpkqIVdAlwGDkcduFlhXJh1L/oCLjSldzQZi9IRTZi9
POZF0ktTW0aGVvDzBC4GznjyAMFaccSc0NwQPB98rRwonXdrX8hg3Um7IzNDjkLjMKgtiGqaVQsm
I7BYk6EO9qHoZBoiYvbrvUI6u6Tbeynv9dNxSyx06HYKz2lK8J/ix3yRBGwpuPViHNOWr/dLCpKh
QMv+56YcHYnY3HV7wu1d22MI6MwcKTPEJZiy6sJlD52MaG/VFp1uETlBLFiycaB6SwlYrItrX/Bq
QMFpQS0//ondCUOzy02DawuakzAkiUMmqhpS73+NmSscSRHJisKASVDGb+2aS7ebiuDBSL8ks0KA
Cx2c4yjedjZQUfR/b263RNL703l7x5LOGvWVbQlv8MBOJqAFJ5ED9LYhl/jk/mI+k9MFz4rhcHnd
7wcclqIYEpa+SBxvun+GeR7Z4WiCWJVukBucoUey1FDqhhm+ER86tPAqF3HXZfcKljg3gQT5VKc6
7/et6iBw2iEEPoRTaYiRo287F9qz3ynGZp0A82rvGQ4fKZXz9xO4dB9NVJQ6K6OU6vEKQVnsd1tR
hkBFHCi6EdFO2rUvHB4VSn7HGTgdGUw6jV3/aXa3smZ8m9K2LVQW7WcLBSGfQjvJymYmBuGf4u86
OQrSgnJc+4GB7KrK6yTVTwci1jF7V2HkPFZS2r1krd8qYj0qN0KWWETR86aBjMa5wYMCdkPdF+Cu
CI6c8jxO0ycUvKx/LFfwLQXPyFCTwF+8T2RU5bXrlgZ9ZJe4F0JPQoaPV2CMvtUPxhW8OFL05TTK
71erZXdIQjdIqyoJuf2yXzfxZhA1eLv5O8SsbfNsEcG3kx+c2DGcy1cuin6EdwsM/ymAzTAVOZkr
nLLTKN6+Qw89jaYtjl55fg/L6ZlyqRMKKXwzR+eTju99iCqzLQ65fqB2nw+AaoShEFsuZlw20GkL
wGIkAB+xzg9B6hey4ryxghNbcJmhfHchTQOijY1hYbUP9Y2SJ47RZTQ6a3x2Xcc3jbvmRCRtfZF5
Dfpt4YRgZL4mHbKoPmT/3Lm5BMs4sJuUOKxC9KTx5dQBlcfSp6uedN4F817OtEkkic0LoeBIdcDP
zcVG4Ju0YEXNBEbujAqhYNEWcEc4Q98puLHBZzAaCqNrCKwdXk060EQ+afPfqbrUp5zI83u+w1zE
34MYQb+wKP3H5Vcg/Z6EYhHOzJsk9N5BDUPmrbeUz9SYVr6suMxi+ydV6CmBBuW42lK4MjcDguKe
6LFOOGY11NWskxxZUb9twcO8g8Zxq1Gw0OwNu5bjpCg2E803GlM2VwQ/PgmamP3EkGCM6jDaUtFe
zXQQn8jWaGRJrtbdkRtXioUDDgQ8P4rkS6+Su4SbTyNVLbHzqt0ATSs85Pujmc+xpxCvgpG+xTCf
8GGUcFeBa7Ymnh2uKI/SS7ywM7nVuOmzQWFTd5HCoqTim1HhK13oclS26yHb42PekJSLWnlfzMmA
NjyEpoQrq4qNuM6gxuZzZlHz+V9dRcG83xeeXl94/jQB1TPp4jQL7QGlHbxOh6oN0Yr2cdsbeFub
LbAqhhzXXiafKA2XoLRDuKIoJWngdIXWF2PYlN4xjJE2263Es922g+7iLpfSsRqFB57v0y5wXN1U
usQQa3P+Q+DJIDxa9OsgjWEFi4g3lRairBMo/9ISHYkGoueVYxrA0WGJOl9JlnaJhiJ4PSZkrpR3
VI1AmErcZ9cRHnltiGGO6qTfF1pKF5KCdBwIpTfeyWzaM9tgJnlpYY1MnqfpGUFMd2xcuhBsvURJ
lXsTFhX6SG+dET4Kjh0sCfCw2Pm/d+kYmTWfCrkTA3CoWhS6nnNL2pYdSJfPRo79d/iklo+GqN73
67pYdsb+jqAaF9TlutxM8pEx+n0/xnNTd+uOJwdPA9+EikTMWkzXi63g9b1lEboy9H/Uqkv9gUSI
vp6EmjEHCh6aTMk9NP92Dv2vTRzACUaH8OoMWkYU450a2vVAXPcHReqMQZTyj6/8q8q1i5rc44Uc
BSmWf8Q+AhrJM0l0Gne9cRxxMLy/FZqozdsaoVY4kSnoEVpXLJ6nne4X6LNuPF22n+uBhCj7JxnG
qWo1F9AVxTL3DLM2ffWwqDdCBsaBAVQIUGtZwP/SxS7E2FbLWgKtVi+eg/vuoTgPgZp1CC5e9rMO
luB5caBIOyVjmvYxSFqiTuNl8gw5OGpC5g4AEL2mR/KWvAeYuw2BqCmaztpaeNLdyO9HrZv6Imt/
lkptPqqF2uSBlVEbkMUSLIZiGxerViroMM++794yEgy/ZVHBJ+BfX3EHQO3OkWuo2+RMe8PZe5ya
8J97YXxqES21xLcvZQll/wdAmF1UuOY0ocQrRcTeDWJ4q8W1yullofv8LvBfQaCmHk4g0KjUBsBw
6LAJG2JZ7NgY9Y56Cz/bfHZRFD1sMoL3+9ZQGSuqE6hU0C6+4mb/o4tsGH5mVYgtOj7ti5/2T4ls
qcGvoHNIY5pkUWXkX9jTnb61UZnk6pAIcWmwrSB2IgMDqCmlaAqxGdN7ffaoJmWl/GmxFYtew0Ys
CLiYNRQaBoU5gZuX6q2XTSP6rSjdqylZvqmYbtCJXuw3HjHiXKdUAi9EWGdxVpjaRD4nkHUBGkks
ZQqdNIod7dohF4NKljL+HMVaeRjJ8NHnEAwwEHDjKE7Xg7zTUHIKg5eUKMYnLPkgnbPSZQBJ17QV
3WopgbeNCUU4tgIx0n7eMJo+1xs9S1zjCqNLGc/lEb+3eZsxCj+2E4j9xFQeco55pn9Yj1b+2WLN
rewbYCZSQyX9aao7mDROR18oapDG6psTV2929sqmQ6FJb4VC0WsYOdCy6Pk1dJ87yoDUKcZqLsHN
qNGQ2cvFdl3KcPBg8jyTKu/GA2B+x9RfCh6rRTv5poeO3XsNec15CJIoYb7kyjF316oP5S1FSwJX
1i+kr0p7ZusbE7pS3LXuJfKRLj+51FtpC84oLLaCY/CJPwpMlO8ZpewYIA87DvvdJ1czojFRgEcr
VfCmstqqB3rbjqJ7P0X6yaXXI5V0isZ3aOERfWCesc2Wjo+wBcx5TyEvbS53FX9kx1K5EgetpYNF
GnJ+2d6kVoTLQOETFedjhR2TkzRex17EKR3gVPqU04aTUJRa8WJO2bD8zylSmlT8Jif8YAge4Lzg
7tvaUydeJIF1ar6hC4ACumIZl0zG6CgtnBQMpT+MKJrH4pRkCEmwqC69wSY/inytkiZv+tWCxc4Q
5Y/3L1qpd4b4a6zX74wKFs3C0w+ANSsbRvC+jti4e4ON1cY5WFDmCHDeZEqzsfG7qO+jbnUXx4A3
Hq11wVTNmbIYP9eFHkIU+IlxD2qeWrBra8rNSyPCReXKObzH2qJPLeiyuLG2z8ps8AtzeyHadDB1
PrWq3IrbnvaVeFkzjKu1c1yvQ/CW3gwN/ZsD/AiSS7E+9IoFTeKra03HLaC6S2RT/4Ky+a0+nheM
vD8sY0T7jy229oaNUhbQVXb6RFA/05ErUJCPyGehZT1jbCsaAzrwY+mjWzd0QFbi8dwaOkSqI5SS
TAVcA+JpErXsVvE+DeuDhCNqmku7lNb557Xa+6g8UiB9HbTBYwg6jsLpT1+blCqgnzU/jZ/LCaAY
D3V5ftb4yZs0yFycQmkqa6+kQTMamO+TSC2u74vqsqfhGBilyCKcAw0ZYE+Fd2VPskBEkQJyUmhv
Koz4uZJq50HdrTW+WYVpvEAKcLBIIK9SxsZ9Doqso4NEZWxZiZpjBZXjoVAJ6n5Tb4EHEDiVlVor
4ztxXNvy5MnnmsyRhnswdPWeVxzlfbvY6XHSgmD2Mr1uNbnXZklWORIZclRheukUilbVdgolBQCO
1f8/JstHnWSncwXUyMOmJfsFaGpDYcHsRHhO1J/5ZvVxdlwef8/ImgvYeQ/UJ/ZogfOuN9uI4lwS
2ZL9uydGoQVIDjwYEoXIo9aOIRPiHax+bUtBAV1jw5Md2s79/DHbvgvSK0x7L3OcQ8wmdGH+GNcM
6FPDGR+mJ7KfmHXdWNQmAe/jwCCidxC/BeBuQaiRKfHJM7vcfQVMJBGK8EdN9a0zhZNX3fNlSZO0
AGPe295dRmQuOgTszkwtoy78KsQ7/gE2SBA0rouaYPiUpDrdcqKDn7Pd1RrzDlQMjym4wau1jTfb
DYD6NU1sv6XFxikbfMvZ3p8J3X8ds/y1qFkSlsVq1PzTz4lmsKz+ojWb0qgLsmme/pLsbcjMjfEl
4m1bZdcybWyGpCYgG+7/++CWNMJ/3vV4hlIifAagbwmxe5fVZAfIvzFOPffFy9TKmV1ZwbSPisCt
DR828Z0p0cGdqvtGAJ0AlrE9UMlb2axsxT3lKEa/dYcBINDKDVniaFw+D7LXSq16Eiz5uSyk34r8
086Nh6hUvIHNReSaI0wNZ9wnTmr/qqA9KIK6W1q2Gmm0SJKPJlq2/OLBJDAgIRaahgt14ocI8KbM
KZ1SAiZCy3/60IcLT5I44eaBfNegOsT6ZBBAypZJX0uWLapse6YDdqvXw8kN4Glbp3uvVLsxxwK5
m9GSZqYmCfE1h+xJLzZOe0Hj6Kh8TTDJln/ZIQsWx4BNit6aQWz6ERFV4hys3aw9lJ6OF0WB++Te
ocHhfmy63CQIa/xM8O6Yrg9HCBbPeUpl6mbOjVjnnuCLQXNtOUC7srry5hBkbE0IU3s+w37gSjTl
76BAQ3snPpcfp6IqACCK9oWBei/Q4KLMN8xZD1ccdgP00c1Y22U/n12gSi6LxCOjpjr7LWs6Nqq/
Csacfq2QHD/hbXhZPrAm6kzlXm970oidV2GESEnOmME6B+XbCW29hOQK31v8E4UqTDJMda1Vjjlk
uMhfIRF8nlVWEEgwtXatde/5cpU/JoVWBojPAwJhxmgUok4I7Ob0vFufPWJxoQ1+Pj/OPaOxFIkZ
A/ibBkOjYFoc9q/5sGZBZANo/4sZ3B+FyMsV7xMQbP+SpG76l0ns0aqMvgely37e3iPDruEoL41L
IHPtGYgSkTxRcwWR45N0zKmXVAG5oNAe+sCCHe07zIkw2Lk92w8IUob/yuMIk/PzGe7U/dfWnpy0
N7xvD4Vkx/1+g6FjAsDwLFoulRjAsDCAXxlu+cVLEELHEzP3t/ra2a4vzPSCewv/M0T+hCeLU3H6
URsQphout+C1agPwXKRex/oDudk95ELGuTJbVzB3XqG81KptrsvdFgK58MYUfsaPV8fPVd/twM2g
wnCOHQoOAzu1y0SV0te0YypRdGP/YQIfKVjETuYkCFF/r/Kg4UYTJ9dxMnW4C4G+B0WSmkyi+N44
BEcOrIJt2pIdr7Jngho2IjVhcnWQO3+YcQ+N4aTMhCbAjaoOs+8I/UJseKhwOejndQxUTaFCpMBU
3iZ7UPTBtuiNnAc+irfGCLpZzzyMudYbSJT7f61B3E1FiQfnGdU8s/1xubwcpo8F+rN4uiZrwct7
gAa8ZgoMRspsW9pt8MKA2uOA9WmaVoOmnVNZy+GObSecYaHwXnHOQeSGc0ohJEDKWsJRwS2IBlVG
XvMWWbLh/Ghm4X1BmsGZdhfWAYHrlrq4kcmc+BTJnMs/kIoLnFrjZWsKIlJXMsb3YwwsTamA7TAd
Rqka3JLDHLzZFR4Z7XRWAkFeFPuHILBlE8uEGWORz2NqYlqb5K269jDPSKTiYE5Q+uzLYbqm3qtB
acr3BZn9zrdytFeK1Z9/gbXuYbChuoSmWsvWpyo2NPRsckF9E0WnGBTGFEVYS6F3RgxSCxBeUgQl
s/4REn/gR48M4Az5ybvWYc52yQ9vI8XfpJsIgl7rMGX2tgszIhlaAdlQNnPquA5KY4Zgx/zBAcoq
hPBux0S0pncD5xlvdeEZntn3iAUKUp09N2BkCDNASWH+Yzk3nPxhQosH5lxj8cssve54zllu8FrH
NmW2OetPMzECtd/JD02N21eiScjv0MkMfs1qG5vQtRkZIaq6p+17Med2/VucpLp0zq6EYoyv/VPB
aU2CwjhKfPHEkVDU8wNGmecebSiyBKb8M8OZ49zj50pBcxIBbMeElq4yTCStCS9NT7tDLJzUEsVm
qzMrPSBAa1m2teYM6X/UWkCouxRADJtJWlCaoSMZXgUC71T47No0LwDzbVr+Qh3TkcGj7vvv8lxQ
gJB0ugzG1/UhzjLbOS7eUatwJ9371vrD0ILG9yXENeX/FiQ9nBh5tidWmxgwXSJ7QhvwwCLrdIY+
cVMXCxZsQGWEuSBj2LyYYMGoYrXtMYdJZW4zh+rcnDlwUVVABoGHO3DWm8DjoEIp8Ie9iga5+5zO
PngWldRRCOQLAS5mdoTkndoMG5EQwY2RfKgNumlSIJZGzq4OLXbg+JbJepk7e2ElOV/6z+yLjSQM
Dkh0vy2pwKr0Iu3/X6tCNz46PKKzRpudhg+RPNye1ADuWAe9vUqwZ6GB/yVQ02ZfFSCQxToS2e69
RIc6h577A9JPm0Pn47eQ8os2SSP+u+fLBTWAOFai6ePiXCWWCvxuIAc2d/gf+zj7ZDeoyYvxhhuq
WwKODIp9IN5znoy3NNhpN+SfWfvgoL5dMqkiQMkoU584quxAtH/DwU4cxwuCkbs1RnL/mAPGX7Mq
I1KNRt4pG37qUJMC+NZ6SNl1ahpduTQwM7EHujqBNYoRROJQ1xGDK+sqpMSRcaMghncQyXttmxil
gwBbW/S5s7cK7xqTTk4g9dzJujCF0ZsAnwimydziOkVtN+CfA5LxPNXHr+CiRel/Deid/CyXLSX2
zx9q8nUjB92Ouejx0NFz63XBDZIlGPMSI2OMnfR4S+RCVStgzySeXEudr4FGhlRsTUKVKtZCGow8
XCA2BzFH0mqhk5vzXNS7vJTIj2Ri2wQDcQwMCFVcODPajv2gESiPL5mEvjDMAMCvwUbSNBVYHZJY
TP7lsimLoF+OzKTwclLG99DFj4JxPatqF+KfYfO5oGt0WSBO8ORgTSDYKJhPt16txPQ6W/+cVZWq
+7r1ZpOmKwF/IsnAdAjRTf8gk2A0clmMlG3ccO76TnhKYo1g/8VmCR++isU7mS6PXu8WcNJ8WsWh
3VJXQLhIVU8OaMQhDQX8jMkAUvrvdZRcLIvU8tTHm1rTz+neZFFbA0MyKnRi7In7NlcV52SI9wfg
OJjZNpvkFJLC6V86iNyGn80xr70ur3+HvEBKtJuj0PThjH6ScIGG/b+/42J9a6/dO03+h9t0M3iF
OW44r9Apr4f0fOviN92Gm4MgBKTf2RNYq7v11ZjQQlndycryhNWw5Cy8WOe5rGmUIDB7eb0tkvPC
e4slJAiL2qo03bP16r6HWMCBAOnO0xxXb6NSKCLNp3R6cmT2OPhtj2LIY6h3ASvHUB4wcAxuF/Ud
E2441d/syV3/Ma84kRVUI4eUaKD43uLE+NCHzLjaA7zK/raHmdNy9yfliXZs/2fLQSxZ/pp2ZJyd
RXG8FlAZ6Gu98eRek45pdPKsQKisjBWYC9ci6+b1WWcatIpCKeUCNl+4mM/O81BdvNIEpEPy7Cu9
AHuucH5Doxo59lOAJmWpOy1+DlmwAAARhAWTiYNneC53UU95hkrJiLLj5CexdbJSeKr0llTNNum2
IyG5svrQPJTO3dW69FOxSWdGWH3brnQAOV68YZQAHTIv8ZIBbQMQ+QTNN2QklopxozAQ0BUgNLur
7QMbRwDzA7CGdUAAcrDEIxJcCrCiTlRXzUPQ6nOXzgO3V/fWI8GKk0OKaj8TDzF2FfB3r4CifiFJ
NVM2BFJu+kg9P/vlK8IBGcIt4bXGIUglD3xwXk/DRiV5wqLDOeAnHG0gPcTTy6AKDPeUp5IrpGjw
uJnkbpw9m1ppayhhd5Go4yvslZIzzxxAUqLrQlmyz1XIcLfVvh2sXl/aG5EOf39C69CXPfomvjnD
tToGzRMHmwG3AU4Mt9ZuZrrhENr2jGLo3Kv1MAeNJpFijBXyWFwQcUl3Ep8HklF9UExlo/DRL0b5
HDjZCF06JHlq1pa2zhFRTSEDCRqdBB/lUK5OzhedCNH9eRYg9+9AOjMAKB85c90wiYOw1YnbIdmG
rfOtCA9Eo+QBT/pDOBr9a0TaJDegY1NjtHactAhHz6bfGdlTj1B/p6MzJUgbVCBHUITb8IDSPrAB
+iZeIvKC+wvRGqBxIO6gfG+35uVqbfjSBcm+L9lZwtlRCxy81Q1r0ZgTF2vuVqnMY8/hy61aPjSb
CCzye27Syi5v30nxjQTQ2s2QAjUVKdvD11KaTM38X7mGAEnfqKGab/QWLWGTXMn3ZLHICLlypV5w
BmjUn0gjjo7LcCUIp9ySWHfE6iR4tkW9aiOY/k6oVBmiC4Tqt3CVEIMSEoa6CcpoJp0smkJxa+gC
95H1o59Iyd840Y9nvyJN7CStb0tMmSQGhfgQ04cpisZ93ytTbllssHjLViL7+dkKNfDZdPHxeAvf
+th3a+PorXie++j6G4yTnnJ7MFrm4uN1qt229+nLbscg/UYKcIPnvPX4qx4ytmxn5GImdZziVfin
BalC5BRp9rErwoSz5N7wgQi73wv7H/OR68vfrwD8ZucJHC4BCkZS6IxVklZyTXS9kGLM+xcrnHzc
dSlhKr4MpzYtG6kqKUQtu27kA1my/tgqLwsaX5JHCyVmQtIgIRvY0ATo7fWRfOCzZO8i+FKQhHXI
wwbNEjdVGJ5R5Yj0dwqEZ55qLziY+cqUKRqLeSS77wv4SC5XPJiv4N7KDNSPwTHkCi6PaE5IjAeD
FB3Os5tZuRX3Ixx92f+PvDNAyZqoSHWf4I3h/2XERCKanGUTw68DCW1noX2Z4P+I13+WWyFd4xal
6r0OURcZjNf3Ih6NvXsqpoMQSez++4N8Bn3s5E+7OV9ZIyVznbBka4zwB9/bm1olx8fCVw0DVoXl
QzcDC/SS3DK9yGN9wRqKk9oU14FzTf5K9IyPqoWuQJOtdT+EXS55p+k1CL3arLHlt9p5Ywe10ROU
ucPhxvYw6EfN7IoFOv1nLtuBFLtahivzFbGbxbRIbFbR/gcH+QxQyTcDISA3+vFKATxE04QAxKQD
AqJhKySCOPLcvO70RhAOjtf+XZ10g2aI6LFcHs1EwXPNJesOiE9hU/QV/PE+ucY9cYtGGzAf+tEm
bBgR2SggeuYPXvMiwOBSkrPJO3QqKgN3/bMe1z68wVUif26L6yeXoKmoEDNrk0ZUTV6U00aMnueL
THQVFZ180rJWIH7S4OwObhNLuPSlMfTbvye2gQ9PAhoDtDnyB5HhKxBCPtM6nZVMjxuuQNraSjg5
vgJb55FVdUgRUXquI/d+FOBeDh0gYr0iX77QfFWk1qefgolQ4em+bKNmckqd9Twh3v5PtQQEjaF8
0ma5J5uv2Q4kF2CGxNdh7T/Pkyv4JIF9bduT7Pk/HrGykiWuiJ+I8aY5C5ZrXXCDieg1bVFO/2Zx
21s49UjDWrH2RMPwiQ0knHWpLzrWV9K53anPUps3wbZr0wOUBSkxNLc5pgtIe9sKvmwx81VTd2Fo
+tQFDn7l4JtEYUQPVbfakjxXhgGEegeuevcMW5cvDPYRIfGsSw+lX2CIpgprSvFiFIuqXj+L+x09
cAw9bY9NGiHcqFnt6GX9laDsp/UJgOszNyc6Iu26TVMM3iiTQ1hQpXhXPJ/DiI30DINVyNh1LNEQ
7x3o54Ek1JAro7ANgKK0/GAN9ft3coRDBEm2oFOA8nrmQMaBYHBp3hOgw9n05Kms6th1QuUS+wEG
r8hkQ2AZeWvoPEyiAHTXxtwXquOxpsqE1JruA/JFBf6UoVXo29+XgayYhUSZiTjhhdjF5uTZVpsx
RZ9gIHDKlHqVlmt0tBDcLrUL3KTIWqCu7hr3jzrQ/wwABqhQ22QkIHWOMYJnxwVfCKskDfZO0bC9
H0x99xc6DnIO+iLdwe3fRuZDltF5pt3DCYrLHlxoYl7w/8Fveh1oIZnruyMG4aF44yH++nhzIs3D
/v2y5Wx7hBW1vHIMcOibBF+VRzGxBT3B5uSP+I8pELGDCGWXWooTr2PjCCJLNBk568JVzG2LrOL0
DmbSyAwbZSEJa0Gn9FmrUzXTSj9pxo7ecx1fFVI1VR46Vos2GLEe0Pw2seShv/5LL0hxKCr9ynfi
4s//Mdd9voQHT3ON9EB7u1yMT4uVtFatUIutonzj73OeHqHSke08Ug9FhO/1gqtuemy01/VW/3u3
uTfI/SuNu5ky7ZzI8HURB+lQGrBguX1mlfuIJ4kvqV9gcs8O0AyZEciWqITuXyTUY/ihf8UcNJao
z5wHF2pahbQtna7m0CxqZ0GRZ4rl9M1Q/68sA2+svhsZlLW0k6jbcCMlWZJPV1C2eEO1PzKnA4Nu
JfoIOyL+aXkeCrvkIPTacfWThGJrA3FqNcFtvHXiRniJ9ucsPxnyMQPKzwECinBPgZJxVqCdEitK
dN03SgY+T3MXwD7FB5cVv6o09x4jP2x8KkB8C+iz3vWZY1AA2k717HmVouExcR73pIY3yxTncefn
L0n32HoBSoXOMoCS5Zm/U6Cuk+aVb+b20zC12RlBdJXk4kcMxtTJ2oZnEZ174W75We1KmX8W9UKR
G0gI2qPtiuhhWY14WcYbPvGryZjxJKn6ug4Bh4qo/no6Y1riEDl2ObQDvlbo0a5jgwfXa+wq9GtO
PrTEEI25rR/WmnC+6fD1j+qBMxcd9BYYZjhyQiZjFdPGwKIoF4GBBbobv8S2W7o+PjEtBBaypb6a
8Ge+v3qc4YbDIIy0Q6mnGmTI9Q6Ia8TS2sz4xhhjKUvepzFch87rX6i31ikvpyT8p4uecSw3Nw2o
/uPGAPacnQ8Pvh0eHIvmQ+INq4G4mXPD4yo8/LkMi3Y4pPE+elOShp6XT7PPS2zymi9nV0OpLg0O
kCZmhJfG/cVOxjG0jmyxS2/0+wAjpKw5EYByvyDPIzB0QAP6UWCXx5I/ElGxEfKwP92N3JtrMXZb
EnT+8ENWI4BdS0HO4RR3/GDSTW2NV0vMaIUZonvNAKyTrs8o11NFPZ+BpmX+Z+q9/HVIWvoJX6//
YqljQVaavXodNqGlWmmYhcigk3QP4d8F9tMlskYq3+Tb26P17cH/L6Nn5llNIatGKDzcwGil8GJq
If41De4XcswHf6kxMuEfBJ/b+xOH63qwCmYfAWkn9WD7Y4EAsfb7BVabPoSnIF0mi8/H/4Cw8V93
Mfb1DXO6dv2MsKk0v82VsgVY53aWYwkEwgChYmY5AtzD9cWHjUgfyeUQr8B8QWJmm1SOooc3irAz
8hz78+Hx+c+uhHGCPbqpkgQjC9USSjoIYUoHcuIZnrJzDsG1imS+sF5kgGQ9Gamlt8oB7c1PFN7K
XwA0+nuCZ3LzwsvbhL2a/CqI6ftYQ+RHzhS923fwusQpMmJxk+R6eTwvXDQNTuf0JcW3TZRK+84D
4ChKXfbKaMxthu6BzzFHVdWzrlxla42NgraRKUpHd/XP5oc/KiQfo7wvChbCl8OpZjIbGjojv1gj
wYVWiVG92WK4KRyVaRY+cx+lTW+HNR4u/uTHHaqOlxbHlsNrLjHiN5Ti8ErY8xlA2r0B7XxyUwG6
yyqIurxSvFokNpezuQ0mLBJXr2kQTXmsGZn+RqFlbSkWp2xz0usBrNa86oYTeG5+I2YrDiQcZEii
3aHE9uOz4hubFrZ6bbhzUPUu/Tw69IA+djSX1NrxYy5YbRgvJDMT5TxkAnKYOn+zeSQ18sojPHv/
KE5fWZzOb2Y5LJkT/iRxzuz9MhoOWj7K8UwS41G1b+cDzTAxeWLmrOR4VOiQvmoGqOTSgjhj5s6I
BS/wImSOaq3uvcSVrZtGQNr6RPxcfTs/8YDRWuimZnoybLrd/5ecH8ree8xgzR7Px9+Bzs5D9FKz
gXC+ZYlAsBBuWXlfI/TVLNUfoW/jNn2cbkTfoFU8WLRWqSZbpR18kY7gaebVlqcsopLef/jizB1V
eq6PlVxcbynXQu0QhVphnUJzESEhRzYEMtXy8xCxNXrvPDm4wHNzVc1IKyQMb9MgylLU1yvX4Sbn
Ut8+7qe+5kEBIeN3pRfO5FbjaChMZbq5ZgBvCAIkhJHkpD7SRtNwAtQNThpRM7zWkAt6pyNmvayx
fvO/E6Mr85D9WjRfUBl8xojT0/0cV6Q4hIwV3b3sb/iqSGnCMOvxT/pNtpiv9dJanMYIY2yW5b/s
ZH3FKtVtakpEXtGpoIjHGOjxdNd1Jyw8zmCRrt+5htcD14Iw7G/LyGrltFIdR4WM+ZkZPJyOh56h
ejagtHdt/ju+PQd/S54quYQb9ZhoI2Q1TbBXLJnUIdaSjyAuZHipLafc1zjLTi7EMQT2riRPd3Tm
PT2ArWP5CP/fejLXbWSqxMNGghVvBDprVIuxidP7w18n4yJLJ8OqLqYVM4/++u9mz6/Q05lw+P0W
KoOOLMlqeeGA+tJpF0aRxwXpUkAfqy5PN9JdfJtHEuljS0ouvB56IcP/YmKE8B5MbV8YGxMy1C9C
fJkMNmzWspx4gbaBOw1X/INyMqh2O0ahFV06yajVO6G5IokSIosChn+YG3Ph8ScnPmDcn7BwH/2K
lGsAKwWEXaZbkk0y0kqQQx1qUUrSXKWh90eVOgRZ8B/vno/0latoIHE6sQ9xbYr0k9GdfO/9xyb4
cX0SUfwB3a77gg/wKO++2iPZTUBnHOUyiPHUlm1xl0+CrFsAiOFeWqwybdZ30sTu+YPDhXwMRU5D
89DaOMoOSSVcxJOsebrM9XKg08w4jXd/Cwo5pzxGg+YNEznqt4+3RMBJUT4PCeqlsqnyGUL7R/CP
VK2TSzQ+zfSK9RAbLmq5e9lLDrSIMFjASATT5jq2CBkjZN6VEXpYm0JV6u8vxGbm/ptDvwGJXZNa
K1z7uDQCt9xxTo5xIiK6u/00AC0tSTNkKa/bV0taZZyYQmb85iiicR/Sp5D9JmsogDgVX82DRK5T
dqXxpwBg4/tq78tcZK51RuIbtr28CRK8E+t6oyLsHubMhzu1OC2RK4o90M3vVgUULgbzFDgNzKm9
ULATkmRxlKHuXEr6OHaaSS7K5SDa6q7aOzM2qw7LaWswkoEgza7p9ik2KIne2+NnPhPJN4uZmuxS
nouXjfj7PUBCkvj52EHX5leGJxvXJZ4RJzoxeRwrSRGN1bjEFdlbam4CbDW5BKavnb/zSJhKSlGu
JUDJbSpgGxzS2I7QTIsQREjQQGFq/0Z5Jpmf+Sd9PFNDhqRMBZadU3XoXIF5NdCNtS1DDmyeet1t
ft3zU4YCKLKk/AZe0FB679AAeqSSpxGBbqj+xylBZrHG2ddKFtNUHgpFcj0C0z3PF0VsWxNfDTh8
wi8cnVxhrN8tMRhh3hxICeVGIDbT89bo+k41KQqVKJ5M5VdTm5EClDrN9NktAA9X1UZPxkEPe0Xu
fYgO9Vus70SQaGGMU/IMExfNbGBVcp5wI1gte9aYc3OtWyYQl0dZBVu61yqEDdgtrXWpygkHBObq
5xoEpjzEhUhInkxrSCJlHxeX2qVccEaeCc6RjXANB4v+9hJGE2MP2pgDwWRCNFWeIaIXWtTJyK4N
q9RcFf1qqyfJckSr+13w4pR5PIEdec6gI+mMb894fpstX/FgPLtHcwxPRbg/JpDma6JijK4SJOYX
dGl7ApHc6L/dYK059FOKDS+oZJo3z1iyuvmvnx47kR0XsKOAOUkjpP/P4jdNAp9FHvyLCbBqlVPi
RSCNDwm1vToqFdiZJvKF9CJr8yyrBd5SFW5HVw2AdjFFLAFX8wx1h8ViTTAgI6OESzJ5pL5vvkof
BsMr0SZXocJEgbPGqdGN0gYOUwB/PzDKECmBx0HRrIQJipaqiNqYJwDimotx4fq5b84EzQpDQIcu
QQNQQT2HI/+FHPtUeFX0KsnEDNbbLk3JJu4AwDzHDFYXERRyjuaWlDP7G7quHdyrJOhRy1chhfBk
GWc33glJLFRaACqsrGumryA1HyyTEdUTcBm9sZBvPo7b7RTxEru4xdSdDQBLNm6LAwZMQOLKyeUb
ieDjPZ3NvFRcBCcyt1EgfMDUdZHnQsXRqrb8Cv4kOwesG7Zj54T9UsFqiexui5nX/qOrQVzlzWUD
nRT3ahoyx0qAFf6gAcAL+sTetpoOLVCL+MqCI+HvERlboU/cYEqNlV8h6MRoFDiGjJRj0GA86kpv
t8bwsV0M2PUE1B9XqR1jXZP2Enc5Cp+doi73IxGkmJxiGjiPNHz69NfdR4B4s5WpkaP/edEVcIrQ
azSvXD79UJroj7juxF/I7zh0udORE+dO8FGLv0kT/bvKj5vb10QP8Odguf2f1cbJUUWo9Bw3SLjb
nJPoxA63BHIXfEXCpsPgVDXcqZPcPJlwy/ghdqJMeygWeKPvRUzEpcpEMSGhKyS3l15fBG2r6dMh
bKE8g1rX9NkvFkNh+Wq5chmlEClBrWdOQTWgxxhL8vX37NOYjzzdzy3eCrJMaZ3Q63Yy0f1Dx9Rs
BUcn9OTuIqFJAgNHQ2CPU6dghlqrUAfeRF8Z0YdyKYW4eJgKFPtA3RxtAWny7RxpZ53mNYtrT2r0
T4fcR0pI/rr/iV19gLvUK7tujS6giZaeJDlztGRiRXfW58N84Q9/QM5y4QsPZL/hc6tMNfarADp8
4InV6D7iNwvlT8yC0gKAyPW/0DrIkZNp5gdSbwXzDmHZ4q/tpj+jb84We1k6z/OopoRwZlHji7A3
cM6BgLfkEGDzFvsirUI0uE3BJu0xkbJloCcR0k4XZ+tb9GS3W178VuJI5gK4pa5NEPnq6S++PuYc
9QHWEZWUwMcmDumnJJ1IaT88aYBcCaglL4M3VG++77xuqPrLdx3m8OYXDeD3yCJOZ0NC2LoDo1P1
LCYeg9GE3Q2GSsjvIwuIWQM+LkfcXkcz+WApf3bnS/joO2IcON7iRKB0pbMGIzy2lRKCtdQa1KWA
Rhr85yVj5ZeCTCVvNdnjF3auUNyo/3gSQUguKnMCYhT76VB0fklgFMJlnG9oZjJHjykBKpCNxvQE
DZ09Cuo6+eukVW5fHthIWHiXs6TY0tacBkFprmWtG6PnpfRFboU94auZIOfNd3JIpY6EBSHwWIZO
Ui5v5/rbUC6zMfJrwU+uZzBvG5z25wN7ZGvKQmlOmTXM6SdQr1gmSlXYE/4MM/shXbeai2b91ETn
lCpeMo5p+qeQInOitBNYOoKKBZVAGwyAKo1NQKslqdy1siqPAA69Ab4T7SNGRYKR2p9nsW8SwNwc
NvwJqDRlaRpE09FEBMZd0Au7oAZESxOxtOpZfZQliz5Ks+WJl+KLfSsk1yNKgyjyJytzT2g5Y+7a
DE8mloobnZztzQRNGuZFB7cVeNeiSP/dSVe4paLEtp5pfw/XsoLipUPVc/72ATd7xxQeBGYNp8AZ
+mSn+8e+/2+HMYNER2moHove9Hy3iWQ97yjxeA6m/jWQG8X75SQis3Llh++DRhT70sSUpARu4j+1
q+tuNfz6nLt0DZx/zDoMHc4HUpYXO1E4uNbO5LdprDKXDQVkoLcZHTm7w/NqGOvoSzTOY2aamdLT
jy/A0ESsU/fcUBoa8wbadbzAIJs5CmtAsIzSUTPQSYEPFBhiZR/AXY5Tijg8Xd87q+/xWXrrujl0
QrZ0Cb9aZo/+BatX0hJT667TdPb0gAjzMna57kAtkr+EjTuAfTW+uydONYA289h8AM7mZ8ZC3+Vf
v4+mmt/NAvtt2rnC1t9jflvtg6m0q27uoN+n/UEu2nfX6AqtgLq6WZycBvUYTcZyGElHnzRyUGPC
jqInH/IFWhuG5q0EVz77eZmOG7scqp2bIw8G/dYyRE9MhIk5dLROrkBFWsQ/LCkw1WQMnH78P6pw
7GsDZjB6R5siix9oD9BmgeYAZFSrtZyA0rCUqIXhrN5IYZE7HAk+U6ibPQBQOKxQI/TVD/RYTo9b
lH/+w2uE+UEYaDESqBpOmMa0FAIgKp+1p8DgzWagK4kWQpN0ty4FrnDBlLI7dynnYBG5BwXyfKG4
00RzBWrwc2M615kKBeWJ7BRWTU/y8RKWrnKAeCSGByJbQUWoWjoreN5XrJDo6gW6kHwZ8JpFpKDV
RO9ku9YNdiwE4EuJ+CsnrsOZh7m5S6uL8Zno3GKN22AnCFqsO6dOlGsC3Ngbg888n8lGBJJuD59i
3mqWlw24AKGrTdcwZ6OicAxRhShjYTAK6R+im+dByRT7DLO48r1l+G9aBjE9ReE/GE/0dhew8uHS
xrPFiHvUD6/Ce6se0Or/QgwYlqYYRsQLSUW/NqBnA4tDhBd2I4ewLcknFZtnnWt8LBTq/+0k+PY2
eVPHVifwQncRTTxFflENncqGQ7kgRwPZ76+owTc/ZMX9VEUEn+QUOc6gCR72cSaln7In3x91TRz4
BhzzTarWDuN0E5XAYWGN11TBpbn98Uerx7rgrlO6pFFivfht7xtOt00f9rfMJN15TSOPEEHywnkg
anq9XiRT3aDpuRniKH3Ls5H/cWwK/RSN6kww+Tm0mChY6Djx98lT5aUnx3AeaYVOwDQXehFFlgzI
b0oKQGuoKGPQdqvwlZJJ3rwTLEAwKN3CvJAQGNFSk93AcGf97XlMyrQyP6+BAgpedPivzo1nlqTv
5blKGtfzs+u/Rdj9ULHIw6xw76A4G0vshVSaQYQkSvkE8crombw8VWHQgxIvsrWWjcEOFy3kalgM
DCBdprAzcP7iMuQCHLWRjsXDPOIAE1zqc6Vt/ScPbEDdQe5Px/HC8mZ/CH4nTs06wEvDt0HvhtBd
qv0M65XFaBgru7Pb9ETSk2c6lEoUwAIf5Yhwq+cC6SoNt5sIrO829+wQ+6AE3zHbG8CqztewxXSR
ZEM8KcpoLu7FI+WrTXf+otM9RPugS0JmESjg31TrPD9ywnRn30ji2w0XdkWvC2hCLfJ81w5tgBvv
nhilzZLpF6ZKv9ntNRfQSOuomyyByvZXie0z+4yQFm78w3+a/d7h3h6aMv9htkUG7PWmaGkl5Udl
qRF2Q3bmFzCzNvBkyEI6x4iu3uArRt/+E2I+XcRU0pLgLh7ml5QYKKO7pxpTNtFtlshXWZxmEsE9
hWEvC94HfTbLemAMdfjeqrXhqadp8w2rw9ERhVjKzfg5jAiiz6FRAKf24NxJzUd6gi/IVlkGyRyX
08wRypWhCs27oK2mrLccjugzQJPGk86oy7dYDtYUwP/U1fsYTlE1MQ4So+lqi9Cun1KTUPzVu87e
ASKQfcyivzBPD57m6am3rbapBLFBtxLEVUPfSwjXimMKqThPPem5X0lVzOTP0MB8czEVXRsjfIL2
WIoVvlxpDqUYzEZMmHcLqixzOa6KnySwvbhVPizyEQe5eYByi3vIZ2/UiAoYizeD1if9uj8Az84Y
wLcA88VDKKuI0NQUGks8cnpDh9xkuj8k4aHBbfBOzMEOSMaZgHPVfSJ2GVpD8Vlp4E9ahyEA/HPo
D+Hj+KrZEI3lvvJ68jk1ueM4tXvAJ0n2rDKodRaYcJmvLfMtnP9IAA8LKKm3m5GVY7iQ/1UITCxZ
WxszgGx35bAkI5TAmqRDBz1VUZnayLiLj9vmplem1QW716QL9YLqb2zNbKHws0MNjGbmB3tuZeKA
HJNWrIb35lyGksUZqt3x2qC3QG/+2lZrCL1wQTS5Qg2kxu0IYbPvXK6mKGBZiySXZegqSfgSLCLz
JNiiDsuxXCs7c/X756tZOkWxSF2aXsMcxS21toTZnetg1lOJojHUAQU3nyYMFOfbThYVg4Zg19F7
KiJJ+aB8tsS94u5GM2GAi15Bls+3L3zEv0VVEAg+HN7JK4KGelLmduwcHlb8FCmsUAMcVZbTXPS/
96z4Qc5b7etTzMMhKdQLmMu5PlP8q6W60JEt4fHdDjyMyukpgmhZ3WC1pI/GoKcnL9rcxwuoQOSH
Z6maIlKXuL/dPdtxpD0uWOkSyM4sI6g2lTYxJl2X0WWl+S3W6IipLhS/SMk6XDruI97IAOmGslMv
H52uezVtzd1ZIeE7XEYTzTtsUcK2d/ynWh4b/HwR6P5WNWJN+fhP+aWC3GODJmPJaeIzXv0FA9xS
aEBOX9OvVwCcjALL4oZrB53ZZJ455ukZxbpCAlzRBFhTeV+OGDMyGyRozYOmyuJX98kB9Is78H6R
ypBe26FyEEILKJ9OXlZxaK/DDr+t0BBX0AwjR2DV2hAzb9lzTFs6Z5PrPG9HMwlKxzlUtHP8N7EJ
J/lZnfSkbkfRgkVIw4wt3kTZ5Rl6Ff4TtSan746IkVp6aobMBr2PR6XMmRPprcXTEMHaYDwCehfU
K8SJYa2uLMAcz55P+Dh7dbsyWC2YGpaEjuzIFvxiwgY94E+5AAREB5g5TzT+EO95BTojpEYM7Pbb
Uwg5fQbmNpTfdCuORhnn/Cpgu7ebCF4glRsGg6maM249i6SImF3cydNaCkb7ODv1DQmQp1UB5DdS
ztaoNAIPW3Hli5Se/uy+jigzoho5+MtFFG0sUnd2/zjraovsQ5LvVL7C3JLkWaga/13nA29FMGbb
IqtE09jfsG103Fpqu5avdVuoLCx4/IBIjEVYRvGP/IaaKv0lwZb97gh2UUe3KOJAO4HfT+cFz5tu
BNKUy539EXCxsDkpnUbbrpKSlEEUzVehyteqYZ8lNEa+ODhLeejGL4/nniQjAWF3ZtXyWpVMyQNt
tQmsiXNKEnf7GQXX7OucyBBrRgLVpbp3Y5YN5eSELCPnrGP8OwuGTWtaMjnhDq0KAqa/ih02zGa7
yM5wDEow0bmWiKduC8BQHhA0M8T5J8zC2UgYcwV5JkQeIkLqqUalcBtZUoEmDjVdXpQVFllqKXBN
gHecYqoKTHsNsGMqonsXL/fq2HIh6vybbmI5fNCOrgFrZHIhUrUKWy305XNv48YUBJvD0HWEZ+0C
IMzWvky3Ci0dOUDO5rsQ4oh//fxP5iaz9+OqHJkez42TVwaSnNK62iNTJ5YcJtMB1nyee5hkEe74
Wiiaqrd11mHwQUotrT2XkS/29Ol8eQltuFcq8FAqqFKCO0Kdm9lVYwojM1Ya2JiLQS6+C5cvR8qb
xVwyqO1e4dqvup4lQFu/VYmPhq2ggojvLy45Ctx6qf4QMSqrNRW/UPyrONEtXEjYccD/0u9D4NiD
W3lK1JYTzN2PeX2Q1XTcJcv6eYFYh1dzV2spGz0PO0UkrXyVy2zI+a6V3Vu5UW2aV8cPLSubvGFs
9Bxn3srPUZ7GA+Z+79/Qg3WhgK+Km19nnM6nw8rhvM/Phh0/mPAwN9/58qhycnD7AWJsD666+moR
s5tk3Bjkt+VPVij1z7Pd74iTqXuVetBfqD8vOkw6VrIRPze3/YwMpI00XPSS1ZcrZTBkhGgSCGlH
ZzzgF56zjvIf9fAZIeus9S+WNYxV9Ja8+dEs+1vfAovS++XEuykmnU5X+BuZ76gN1WXWNuA3l6sl
KurCRlYgnBsyln5smrXTYzE6Ir8gaMPEUWgEUv3VO8K4CNv5BjCoP85H/bwT3e6j89s9HszepPhJ
XfQPns1kYSR9zakYrZeaIHPKZ+ptq+lE3rzvDtLmTbHy73fqG0FCu14Ep3CxE4L/C6LUFxtj01Cg
0wBS4PKz1+SvcD6X2qOrr0vEOVI/kyP8VeyaxSeq99ZY6LJ+kWW6F57CXymaxr282vo+3qQHGlQz
rp0KL4jutqhXVi8dMWBqchrgX7UncIaMB2uEoLpySEe9KFSNGUh4mdwHiz4Yz8LCUkkLpVYfbeSC
b0ol7ZGMkoAB0+qvHN0Sqef/enx5wR68vwqRGrINJxg1nsjYRjD3pfGRVGnNpDqmGgMEq2guWN5G
GxWe3W7m1In/Y8N3LCsauaG5lYz2Yk2YEJMIJZdsNdgG7Sbm00L223bctS3qzMnQwiHIKMUKNNkD
CC+XM5/7j0SZj/s+QDvILjfT53ppblrTCHd6EEybjfwUj0cnFQyHhYraHiZuYvrhffH4CDvQ3/sn
SyKzbrtShHBzRDTVqOiNTKo8yFuW0iGVAFSm8tcQXRXVZzgfAqA6H6moGPclN1BervYWviUd0XfE
3W3qoZJsQtkRwp5QyGytAT/QIzRhgMpEMalz7fbgyzwNf9GSxJO1swYX/cJFphloTIZ8SAaN8B0o
rRaC1yfUGzuHF88upM8CU5gc+AOEbBezCtiDhoo7XWUVSSLN9wH68dH5n9vYHJKDLtb77JjwJ5+U
5ABSSFqi2nFwQHKtJVOpp8AwJ4DN2DdN9SehHoSSE+wcfDZiXWOt03m87cJsYqepZTNjiwqwufVa
C2uFzHiaC+iHT26ipil3cHPQdxMiFRLL8Ohg/mlHzDJKdGYxyX7OBGJhesvaMFNEjfio4wIOrnSU
depMIgg3khENheREgmcBcTbrBgYeQmUgdD/rTSjfS1LDEfp1hmyVgLCTO5ibZnoae4y5+AbPgXu5
mgIJKDbdKVI+GMGoBpvu5zHN9B29asAvwMrpir0VV+j4mo45X5/jre9hU71Izm9lHcy/6K2zp54x
ix09cQaAqFvB/cQscNpcd00AZFYR52UAJ8YS8kDYaWrwuaXAekwuvH7E15VSgeaQuDxmf6/krTd+
WsSs9VkR9LmxZe+gWqSE9d9Uw6ZBG5mbpl3ueMxL1V1nj+aG35aowWlLmffmhreIxUlJNrzjUn0U
rYRAKQMvUr1sUjj20Plapyl+mmR6L0R6vlylPPg2TH45HyPRC+uRj2CRJBGpPQTHgfeTgaMXeRn6
6rXZtU2g799ePD/ch/ukcSBEn49BSXEPRtNaJfFChY0EheToS/nOjfvuOjD3yp+tLtM9hWfymakg
xclvmnSU/swpyPRS0dOIWLbyhljA84n0tkTdPptKK0dl9bevma2qFAGYLXTzAhthPmFPux9VPoGE
+mp2PQjdxkoaTJjVE3sW8/HbUXG7aBJ2LrLodgqlUTyqdOpL0KTejKIy5oamdNOzqX3A7rbnGpMY
X0SrMOz1fLpl66wMVDaY3BsphSo4nbHds/l3BDKBE2bebgh+xu3iCqpH+XIPM7yP8Wb/Xe23EcbE
yJKu82TrdLyC/AjpGcYLbbi8yM3Ek6d2cwfOPaf5pZMRf1iH7pOdVNnqbJBMSar6Ws4hk6tjtDvd
xcn927sqr+5szRyhQm0nBnyuOuiHcTfO18XZp9T20CYW4cIi676KLeklp2TqLZ/BKl0S+mVMSKjD
odQu8TgarU0cDVS2R1G5HjrA53CM+z0T7/tN1/5358nqNT7nwfqFZFBRgZGYL68AYpzHyBfzqiDW
N9aKYV2Ed0TYt+OiNHwJlxRiHe7SdRb39qzxjcd+ztbdJoqtKLX38eC/PTZolXjHet7TYQcqJ2+G
X0I5SmjkRTwgC4ElK1ooNRrIQgy6az/DuttCHxG5TT4Z1JUopV4mRwHPpiLT5OJ1tfoS/5Gm9fZH
Sk4eul6N3E7sHbwZHfqw1vSyfcfg7J12qvamJzBSqefsUgv3Qnk4pBuGaUWHsFL/Q/b8d0OUqHzw
pZ5SQGg89F2v97v0RLoasC5JEpucKCvGXXurY63MO59awffoA28RQUjg/fxiMB0627KoZJ4pKzH4
HVzBRtLQ3Z5OD/CaFFA4gH8mopHaMujKyE1kzF4ZF8uLtYj/cTaj7UwY0mzN0bafSku7tdlOAU9h
07Ufylo3JorycfGF6O6KIy67fDJAcO4AgeoNn0ORtEKBSBEp/EDShryN1AZwHQxgXcBY8yNVp6fu
mxNIb6ncba4BbNbIYS4e6bdz4eNmRuj0w2dKdxndZgrP61ADCpPCVAht8euK884YrWrjiiFST8lX
YJm156s9Tpnd6uAz8EXlkar5gz+drqS3JQfZBZIUwZo9ydozE1z+zriYQUeX9cm+a53Z/jKxJHZ2
pz4pQjWV/xTPSltcneTUibo5KAoL4tFzpiRp/BX0HI6JRg+AzKG2di+l5kaOVVUbrzkUolNcCA3P
IRBP7wXYBbMT8XHKoOdKajGSfbJyRcJs2+uHWWDNKSilTBZNQmwLdd2ad5ulPOdfNfaJdWbXveBd
Puwt5hXFYTIGt09NEjDxTo8oCc59n4V5cgrWOXSZ2Txl3aAKXXdMB7PZw7fzBXBj5dsGRDkXC5T6
KBdmp9oMHQGhe9TZwy1vqvzE1X5wmgA5qXJ4KSx4biNwKAcSg1GbhzYwqzKZJM4m7WMf0dd01rUw
Slz9FVBk8dlTn37Bq9IvA629jQL0d044UD8qwOgNq2fxww5OUpVq5g8VEj36MiNr9eBqrf8AmQlS
M4qkEB5EPUuPwk45z71iyKA2QBG6E8Ch3fu0RAjxzQ36SXMr7rOy+vvEZ1eNeya2PKMxEUrXFxSQ
KjFpHvRTAX1SJ2xgvFiUWkR1gQ2DeL/uNsyb/4DaVSlYAkjjjnrCdUaw+cKJ4qSJ/uIllcrZOnDr
7HA5N7AJYN+C6embvpzrKYaJ3gkd6tT5swmAqCiBf9tXQtqRC00tiq6h/BWq7gIpXZsrpf2p/l1t
7LvJjhqIxQyI+kQMEjMd6U0Qj6kW/AU1dCKyUN9+Voh97t+p9jvZyBJFAVwFdWkm/OV1HhIPtHvq
99mGMxVWPFK3jTcrrzJZ0F7Cs736WAtjM0mPKBeI4fpBzf+1iMg3kk9CGVBYVuGLEI+GWBuf8MDL
StrieAC24JY1z1nKEbo2X3J0TuIc+7JvriEGSYP1fUlUMuPGybXEVjrdHIJ0T8lDvUc8MxHaffgV
cFIlINSoBd22Wyx5H7phrvzEOpeNqsMRsmHHU4CJtSdJvC8odyqnV6ounc2AUAZqN+65MDqNpmjs
Hkmuvx3FBH781srjz1g7Aqn5qrmjbXlhYzivhf69Y8HEeMRcK5G2Tvx4SjpxvkMcOE0WlKXT9Lkk
UG+bDmmk0H4gJOY03iDOx6syN7jpb0UGTpki33MO5zm8tYWBtssZsHeSsrVa+3xFyY07PDZ/Sc/n
9boNV6V3KXTqND6IUeWXpjgoBEomEX4+ifo/HPJKIHWoiJYj5FTFcemK9qi/ubTvlqPHa4EAJmDo
vpPw5EjH82CIAzwSKU29xLHi6XjIN0gB8su6vrIs9Y3WBNXfFlwC76SOc/Gs9rCPVnCD0xvN36ax
5YBWtqDkC+8KqWmD3RD3Mcfg0lRc1Dz9WQppZfU99Js6mcqojNUUfpXLBaovmAIdtywey8cdTF8j
IdQzUdvRzVRtJN/2xMGOO4hYyJLV3I5QuOC92ZKpxkZUJj0lqmb+Le0HU49TGrWhZeEHKgfZDUHd
e9erhaR4aFBLu4AMBjP3YDnBXrHce8y78r0ovACI1aklE7mRjbKsEVXIZESoyoRyTTMUq1i3eNa1
qG7kvATP7U2UdTOlqgxL3Ydbg4V/LWZP7k/vz1ink6c0G8sPRbZ0TsT2OYLX9/HgTEdO9Y+6l/Rs
XVHLVppnHM4gKphAJC1Pf2L6sj9528kvFxU3t5MVJpdUb8meG4Fk5N0MJ4MTaSg6JoufA1qUbELr
S0KKeRJohR5ChQLC+JnKJgQpw3owFl0HeRTgGoKxBaJ4hwd98hUgkgaB5hpuN7RxdXIfdL/3lQUN
z0HprolMSKXw8Red6fdXZYeLo7vCcB1YP40dtxKeai/9nhJWXBJ0m0Ay9yKb32EtDW2AeG4w1R+J
aUQ45w1VJQWeGQkX3dsjFWIOn1GdtH62tJ+MJL0KRBJsTgeST8iuXnl6vICSiYflYifG1tpxJ0Sr
yGSmsXDvIF3B/Ab2uc/3NpkHeu1UAR2lrXMyM+im++XXPU/qOqBu4ehAEf8TxoivkjRSdSCJn14e
6AH7dsq9b1ZL5sfiX1TBldKDcQ8IHjUI/EDAAV6PBIHPK2f6bfy6k2H/vBRxUs7vmMo3gtGNYOHw
Iv4LsZPg42EXyYeU7Vjz0RqXUu7MkQ+OSMG8LQZhzbJZAEs2hXO65JKIUm9cK8wV8/J1mnCYg3ak
EHHaquSCyfzDc//b7P98EZXlD44cCMYwrhI72Znvx8bqdsE6AGo001bvHKp/9Dq1+wkp9YQJmhL9
bFLrkuCT+G+WEvBf5eisfL3OZWYGFDSpQt+VHRneYpOIXnM1VE7aNSKuLIkdDk2BaGqpiF2dtzXH
rCU2143gOKzDeUwFaFrf395HZPcFZeNp5W2D1tIOI4n4Q//6StQzUN52lbd9UgbFC0ygAkAGINOo
UCYjx41XS4ASW9MDGPnlQzJIaCzuUwK9qoEqwEmRVG6KWl8EhR+gVw1iOcS3wn7M3qmpFqq1Fq8q
Llk0SswyTO09sYYiWp3q3Qab2YpFoj0Bmsf7XTS+018GOTHzlGapWn8HcpUD/6dklBEF27uCxgF7
JCTjAR+VEL3p4LMj3bTD/nDuZl48+QoW0S7otvtAsSrw0mTrq73MnTpehui1X2GGk/xlTorz+usz
KlJAwrC0qU6DfGbRJCTAo7f0yI0bG5TSZR3W4gPY7zbbxOF/o6fbDSbuV1USHYwE1AnmOqRUuIrk
91W7cpMvRmu0EdPVmWr79xYOGkX9Z/ln3fMHCdZ2NpADts17o4DotE5SALBGpYMI3uuQ886DA8A/
63ZWi86AiKomohgKRlE/DafqQSAHl1slbPBj8AjItzUEar1La9k1gNXC6IBTxKqYUU8NdToE7HAQ
QWt0gni/Jx/FTbXRY8qPp3oKa6d5W8htl85IUqZGcGX37D2f7wyNbn/QPleREq7/SRsNmoJThHKd
SLGREIqJyPJ09i4Wlmf3pRkJOn9SOTUO6ILrpuH96b0WGJ7MYSWHjONMjdIIStM9kdSt95ZQ8X4H
svmXaq0PmH8kHioHiVD7JPbNWayNdHTUnT5cAuBe49q3MFP4oPUzwvLahlOqkF9HaRDx1LCow69A
YvRFoYtd2VC3mJ1WkcjVf9wUrw4MIJKXxpu8tBlU302eIv3TULgCr4m0wa0H2n8Izuf5dhBbzAva
umpFkJfYOECTFppwfM/5OVRNe7efLixOpvDeD3K1Xv3AfW16iikQRGFyRrf95Q7HFYynQgc4eV7V
7seOhzB9WeUQea80/jyyT1+R5+AI9oB7ZYr5Ar9Xs763ZKUmfWkoH3cyCgsXJoAl6ygbfGIMvJws
MrDL0AFTKxWA33BANLEClT1WylFDoLpMSBJD/QlCoD5O0aF+x8VPSM9kDZwH2y/wXq3kb1O+tkXO
MxRE12GkKikNC8yUVvet0ldNWz1Dswhnd3LCHj19jx12OdHWwsuCku7Tx2EMRe/n2ZNsGobepdLI
wmwJKkSwKG8s7mqBu/EDcz+ZOISHPlAHgqQyyjYKF2OW7hAsSJD3+av9BvfINmiae3sWHQCTHL/B
dx2pSr7NgpDxd1Pztm4dpKelrbd5bKTPqk1LNGEpEubMpQvMg4h4/to9QCU0mrdPwbDJbzs0K9Ll
KNRz1IMGtdIgvb96rd4ItFhvvfkIOS+9dGdGMAc55Pl6cIwmzEFXZy7WGIAtjP5FD/fzV/KxvAe5
oKKCKDQT6CtyxTQH1QaFS5VhUh3tirUDVA8/vB9cG4tCDTbbk0SV0oxbVdt/lQ2gBO6Z1X9MGdn2
Jy33BHea50cuG/zmIdue1KhF6pB23e7WB9dfkhQoUbPeEuuIv3paCazVCauGznoalkgmXB97z5D7
REDDv8aBXjcnMGjoKfulMS9NH4KmD+eLWk971Ib+lPEWf1gQeoVv9JBvePImVOkFetA/C/Eg0Csk
3sdwxFhDOeUzdU3JL7VQj2iduNkd+8aCR8jysY31aebszqHmLPUu//4/1y0JxE6tKl/zbxFqBzGh
vIikuvOoqOizRIK7sG7vadUd9eWpGA8FsEhrIHAS+/6QDqBjo881H7CorCXMXCtyidCgmbmSTT23
q/zD5yR+2yRWl67iLqjyQ6MwOB2KsW1sJN/GvZBHNADSm9p+ng1Pjz8gim6a/MP8JWQv54kqO6ty
V3UgTSQw2OWBS9V0bgsCucpMoXwuFWIErFQYALKcZLGVj0oqHAEGZMSGWnUBl3hB3fCzEoVDvz64
zO4sz1/xpzLfoc1kHhtwDgczYkC6JOCGkIrYUsifwRbnwEo38zUl6Plc7W1nswdtldTGO5b4ViVl
uSxFUJR98ONN3bqS0OkKT2dHded+//mrloRAkbcvqkBXdG5NjwbPm+9Z4ipo/lhCUgxgAr6Ipn5V
/Xs2IK/JUn3E5LMK44+mPZiHw9+Yskay90MYPAG1x5M+Pw5kzlBErm36DS29008j8V7n6921w37s
fSkOxxAmskR9s6kFvp0QbjCgbCybEz00kio/05q8hroAouAduTqv4cetU2xqD4KJ79nZED5iiw+X
IOD2Cj97vxbLYTxeRyEHZvuVOF8hduKrstm7F9nl2oVx9EubCfQpJKnSOKH//Ofq4dT1jJYPzl8U
4xh2TRVMs9UHNXvQi5OPoyPaO/qYjJJxI23EypAIwz9CYqAl9DNzloB/ko5s5W7kUyyUWxe4Y4GZ
Z82PkdJ0N8fKm8JTzOP8a560fvChWd/ZDHZ1KuJMdAPGlqpFRMY1oIWqKAFYB8Y3GDc0MNrKEUu9
YHe7dgpPmYFeJHsTUPeB7hFVkjuQV3Siwrg4R0Xg94rdIhlXyTqM6QllJNgcAtYJdM16jGLL6kpk
sNKVQQ4f+lwFw96pLB+r3y8W6wsE9SQcekS+fXxQ24A9RZKcsHdpjD1zlvMvXdbAEaTbxqs4nFCQ
sAgA2cWBgcaYt44GsAqS5/QNhCxTZ5/Hca3LrL8cv79B8QnV9LxuIG7qUPlFZSvBGS9Bvm3IDhgu
L812U+2NocIWqW/il9porv1BmmFvtyi41E7LEK3NX0FHZxeymf7TDSvwEGY9B8gLdD2VYqgOju1G
B46wJYlRkZCoLuNDBJmqdL00HpMWneIhmyFtdpdjnMz46k84fv6jyY5OjxDTtxpkbAbzFX6mhDA/
M5zOxpqMOdcgaaPC5s1yOw5W1fBPfSA7YIyRWh7p1qxW7+vS8ZgPMBmgwY7qBygEQMHNgxXzxXLS
ytXx4BVIWBPuIZaHmyVs4O8ite+J6IhJogj9CFrbyycpYlLk90UMMqouW1FrC8fVjuBLbToZ+/7A
U3j7pXZYvraI3RCFmVxFw0Af6fD2U1Ln9bAGO6mUo/2/6A+PXTXvxePDXJsjK9EA9uDDJPq72QfK
Jc6oNlwbdR10SoMRCHcyOcXwf0Xn8N3Zt8HzMmn3YMgR65KIG29CayN0RkGkWdP6uBvLJe0OSyO+
+LGmGYPc8yG0R1pKpgd6ev0gnzDFCk14Os1Ll1heooqUrZKJFudAhOYwrRVTPJ6FVo6tZnRa8Uqt
KSluQcFDuP/wOz48JzEobzDrT7GfJKx6V76GxeyFS1xH358lra1H4yrvqVsBiW+jKFe8dnQ27zKJ
bEbUmVTg4ILWCtkfx/cR0CpJxGwTcuVrtYt74oIxTP2n1v7HEjyYGvcjN76EcNbc4Z/gx8pE4hWL
758buG2l92ktGM8rkOWOjhPO4BGl/OgckhfgZzUqUYTZh8JzCh0/UPT/7d4B88EO9zXEOWEso6/4
so1tn88VWynYO7SLJ94rwiExH0nBKAcKmy8yXKRJMIiqka3ZX/YQ5YVcIjCx67dkpHWCSdgbWCKK
TFH3w4poI3PUzWCx0LVJjsa5zWHtX1G1cyYWrspKLS3KTEf3hagQQ0QmRsglVobvhVDvjGkw8o9X
zk3NA8VCnkeNqGuIjYp/Mi8/vWxpvCYXAnyMEOa5K8ySwSis+RE+KfrswTJtmlzKxm0zhhsTn6Q4
gP0D8iAJ+cd75bwGPOBbY6ckYFsArU1CJFBNXX20DFLfl9igPOv67lbLSgR/UIl8U+DoWFz9ly1U
nChzkIiyyWxA9lPXQjmecZXWWTsJ6gE4iXF+NyCYBM3pnb5CNwlT/1CZEoZ1didSXpLIlu/nvreh
riZkYjYnHZcrCgzj++S8erPolaUru8Bl0NT3BybKONnAA+tMJpj0cJg+4h3ve7GKre+z7mk8qpZl
A4kp6gn3q45PCou1wLvM86QRbICPPQDb+fXpnZudmRfnVMlpQGjL7u9O582Fa9vBp2J2iGZBoTpx
XVBqsv8r0sIujXSiYy9yKoKAl+YTooWkNk1j7QwmuWn282OMNBleCD0sGe9EQhUM2D8M0wuUDlX6
tCmq7wVttx37nIZRGxRPm5ATKt5X6nXWFToJGFmyuYLWJH45+K2YKP2kHCljyEVRKV6ydIXxd5KB
vCHLbhYfaqT/81z48UtKkQmw+1R0yQkEVrLGkT0RH3206j5WNOch9gPTVguWq0YEiIG/iqftxfnp
TV5EXAuxA7ZKiplmHZtx5qsKbGEFZJaIsXP7kT0OgGb59iAswAQF5vpnDflSg61cK6mvbmsw96fx
pPTndlV/NyahrmNyQi5aWR1uR37cQ0nt0TG71k7wv/yOMPVKBnh9psxwpWopjLewrCyz95ZVeYaf
YeWfVEwaV0RMJqhXiFD7F+nbgLOL4W1S1yb2f8Clhz3nS1rqcLHOSv8sbacHFzo5yBEkGwq7+K4J
tun9afpgDk+7L56SddGBEIy6h7dUAr+PbPyNjFy3X+MP61UhDl267UjdZUSh3Bbj5QaegUWjpg6X
6oyR33SFJvHY/qVSFFlSsZl615/9/OLHsOoOPhv0gPTtEK11RXQpTJ1kYwl0HmNMv39Q7jNEP72J
rghi9ijvtoxifX3D++wng8onAorpz7xMLK8y22mlZkn1rcDaANj0T2N5Em5q1uZJOg0upTNOJ7+s
KH9W9VGCvH2nZ3uXwz5sugUTJDC5YJsjZdqfIGPWrvF3qfdHGuEpHp6106Nqlm89P7i6KZMpPyn5
K/uTfgBrjsS2pmU40E/teUuTKYkKyyU3O9xUFR18DnWU+EUBWfgfHo04xQPrxGyknEhYFDoABRzY
40zjK5XA8eZ5BvyHFals6nTQRnAlpRo3T1DDJ680t7cEtfBo2YC/VuGsgDqXzrDyX7ZGc8DwbsDV
U4Qm8OJBP1cNPPs7q7Ld5Rkq5bNUft8HkkcnwCNdOZzINzwPZwf9YoKEccncTxB/mtGcMIUIh2ln
YcMSlv32e5v/z/O64NyyTi1kQsKK0StNhoSgij+bhpzTet6gmA8FxkBqx+qCAqsYWSOyGBbzIbAF
9x1d8UbRuPaUK3Wobh9LauE4p6x6bzT+R2TAST7I8j3UcjiWw06wV7PoH2hX6Z5rCECWuQtANwJ2
B28kxCg9DYFKM48/lQTJf5eyOIZgVqXsKx6z67eVaCob5L2EDH9sYrU37/Ae5QvvtUtAkPmftjff
UwLhN6MphqjQyL691u6/65VZRyjjaa0diRd3e+ys5D14zFsAm7zqcw4l1NUiJ/UlDH5PrRjz4pSZ
RP5AeYHom2Kl6tka78EFdR4SFiymobbMFFaJpHXUcmqHMJKiiuco7II2+TaOA8gHLM3Q6MeggZjq
8Td4VynSdyNq1DnIbdI8x//doWzY6FcGRD8uKpTETl9zBNVBfu/8oC4qLQaF0RGEukhXnL5EzDlL
umCJ+yQKL2Xq3WNpoT+pnPHslE3ydqOG5sZ10UKiQeGPEulARBc+ARz9ZGgfl31oXTECBr1j9vQ7
nEquIUBBDY+rDE5QjrFYmUvIISQZeOn66z7px5UyiaHuQ0b97CCTa1ByxI1Jek9K0qT/xC9eU6sx
kOzkm0CA1rNmX2Ud3HIlFIzBUPcL37MxcXbxVCmW3/qjyw1Bo6ymvoTGjoYaqdNGA6g9+kRlb7YP
Ozuk4xF1J5YbMDq9FlyCNQf1pwPYStjVMaxbzYu/22xExvfQwJLQsokHGZxlVpgUs6FeLxJxB1ez
3/AUoUgtvhLkKDv9j5/zaPyA3+Q8BOWdqI1jjJUv+N0Xsb7XV3Pq1KQqAKTrgeY4jSq/6NmGWyxh
4sV7O4O04CRe6pdp1FmX5nMhYzeePgxScULadBypaKzvlhp49JgRTBN0e5EGP7xcJuxtEbbLYYsT
6uyO5pUj+h5rZY8cuMFoSaZLsUbYLUyVykpVVTVLPd6997YMMS7K+ZzQkITR5wLKzHYhXyU03eAw
ATysHEFNNJ4C5I6s8zqPY1ZgSBSMry9nY9PhHPuOKa275QSyuVE7H/lbP50kupOK4l3OVaADSQL9
+GDIUdneIMICwT37skDyLRTJ0y9ZwOhCGo4nmaT8hNMNVxv3OkFANtOxsELCrbRSpic/gE8PIK5d
O8jQ55vXqQuv/EH/VutxbXE5NqCM1KhFRpxEZZpF/Sx4bIMMjkO9k0CigZhKP8eS7zlpfrrzq8ke
x/F+74JPb4ZzqFIO03yt3XcR0aYTQM5F91z5At8ylDG6Gd4Hox68/l9S/F9uxNxgSM+HPJoc1jnZ
Dm7SalyUj23vZjkf2YyKU6j7BfWlamRGDIHS7ZIsEXPnxzAhgPBez9HX+8m7s2LXPbIxgD9y5A+3
4g/1eDAqlvahNoXU0C6tixwoqG7sdqqhDeri44ZW78zZKLIpy0aVApdc2Oc7SWRYno3hPz06d9do
fMkU5adnCsfbCXBNbJft8EBC8IkDRyYOkz0vJxjk34DBGWfgCBaevdqUUnGYrE9qlk4hoOoxpn9e
ot1pkO4hM2EK6I1qc4p7R8MF9PLRASuu0cJhYgFojFDsCag/WnOAbBGi+utDn40AOqQUaP7K2tTI
R0o6XpYJKhYB0na1RSTkC5+fBg9WqQ/2Wh0F9ng2ur6BnWh8p9z+m68mBkYi8bY708kUQ3rnayOO
pb4tjXQZfaV1ucrh9nwNoAps5E30JWNJmCAfUUTIdGk2keo/CqfycxsS41ZqajaR5O0qrfJvV9H4
2qTJqBlUC5xJnpBel2EoKGElk1h7naFdWWo9otDx6SGZh/DtC2/Vb+X+DLRLPDzZ6ZZw+scMweWi
venyAYJAPyI4d0cvgvWlLrBGJeFsxUTsYYDv5ND0SFN/TOw4FKNanRcNC+Z/N6og4eYbauW5Q4l8
zvUQvimo74JksNmzuF4+4XjZGjNcnvmrRLD9HzVEHRGiiziBpZP7sN1dpjv8CDfDHjGF+1FejVJe
+fKt/buTHTh0u+Gmi7YnohNtlmtZ/1GtS5ZjOF85dLGzqpEqMk/n7V56JrsTwy7qAc6Dfi0DaqF+
OadSnZ4TTrmX3gugYZ/PNr4S+kn+J1LGTpJkCc6jCyArhvj6/dJG8KObAzHewaINSSxtxIhSldZm
QKZKHTizUPG8ixMTLQHabpwCa6BGckvHddFj7DAkS6Es0nLdpkZrwF9wNJ4Y4Z2vvVbHaQ4Qigmm
B3NDjKbAB13BtKWjePgUgktob0AbUrtoX6LcSFsz1bd00JFDalSpwKOiKygPXfHXnc808b/SvJAa
JPyK8uZGuGXKe9TFi7UFTn+Belt5ZltZeknnozV0OlV5hYJJDaamQ6PyXkV5XuqZPy7l+beaGQao
ecZ0g3i74zYzv++WEBAdkyqE/4iPUmL44KtwbbyFkz8/MFrnfePbF9wCC1etFUQnd5fVVemBQSoe
C/YM75BVAAEK/VSAYUpEtKAElFTJEIib4SgqKRLrtepJ7iZW3iE1MWsY3r7DuX04/c0CsLo4rk7f
Cz8dz8zjh1xAb4Ss1jAIiWtvH8XWqfMAkZbn4+sDw4K+/GCIAmCoUZBE42FrNnH421GbQdqUG7MT
L4mYObJmboiR3qksKAOhoF5uxVXxvd9OSFpLGvp8ZfoWwZbrx2jl6t89UE50TO6r6e/i9z/1R9Yq
b0H1ckiyh7wbFS/kJo4NxqZjzYI5nyfbAkpOJPCGEZAmVnm8TCibi8tP8BZ+iJnEDOQ3ZKLoj+xk
bARMmOOnSpkMnpWklEfUhL8p3qdQilonTnI9MBIHIB8JKw/gHuR5DdZWCOwixGkw3ZB9u44jwfDP
q96veeVcgF3wmoo+9LuqM/Hz7H+5CjAEfwpYehIL4O6iYrBLlvKZp7/fi9wtKBunSPDgbnHTg9W9
ggYgJz6XrZ/gWcuL2+wWF+J4vm2f6K7aiZxg0/LYXzcFVgKiUkaWmVzTify/CHCi6VNr/mmUy0eh
Q+Qz10GT2qGysqx+2kQYPVeG07ROZrRPXAbdsXZGZSoqRq0mUOe7EB193m9BPGCCIL/kN47+9SV9
2/P5CMYg/afBXKot5JoSYD5CDKZEkgLWewRDAq1s/RH1IB666x9vZ5Jo+0R1alpoggEPr/ZP0Gds
XSHcx5seu6cXWWzNjgWf1o7paEp1H1o5WCQ+fAwhYfkDFiEQEEs1w4pC0fIKwnCur8UNzZROm7rW
vvJMTcXdQs3rCCrZHIg0hmp48eB8g+bta8nFSRVRgmclUEnIZDtZiT51AOJbixd1MVJhg3KcdSg4
O3KcsRVM4O0GTufVRQ2526/R2Q/CkfeG8U8b1zUQYv5ZyBI842GRjFjGgeur7DVo6NlcF0RspVrL
LxZyaAWXqLMkJEuh0fBS27O0YcsxnrEVktGrIPAOBYEQ+6rocHPU8BwPuLnS05nwWx4qLnJP+ZYW
aIeXEo9y4Z4x9R657wT8pn6RPxkeHfaG1ewww4XeUs4do64/tAe3u2g+rFd/diDFk9hek9Eo7lBB
qVl3O3NUwdXNh81flhyM0O30Tv+9phAbGNL3jTJy5JdkPmhQNOBGApv1luBLXV/h0TSolGS/v/xJ
z7LiAngnJN5GOmZrkf6FRmS4WSIlGcPy5MAm6H6ajPZU8LtJubt7NPQSCg4hAA8oPsQh8vXP2jng
6TrwXKZwfUVJQ8yYVJeLdk2PO6JqHsLpzU7IuaEh4L0G23LYUJNCfxNerTpvY7phfNvv15hRX3yV
GbYQXjXMJSRubYxukxvXFHLwQQippFuULcVDEd6NK5TEiqFieQhcHp1ffkKDJYmw2lVc1gXqXTzX
APl1ILzW4AKoxY8aekvigdqL3F+4D8mjxlU35WgwsipfEjy1BAgSM2N1ZIDD955+rUGEZoevyuPz
d/3CVi3TPRA3GgVBlO41ObJANSAz5Sj58/xZHjjTENZkd4sGGttJ6OmX+l/dVYWhuVJ5Lt1uJ/Mf
114kwjfYlQNlB60886AU1hrs3mm5qxay6D5frLQP99+9hFdYNIvH/SQju2Ecwv0ilGV3Xe+xk89M
G3Xwe0wOLXvQ5l/zlJh2G7Eau4LNJQ5MrpXQUwkTPcStlJWjyNFgqv6slux0FwSU+5DIUsK5s2Zz
HQPONq8xhun9RjxgIxge1/6EcDzKxlrPdAY9LUUGk3jl5cLlYVeLxMCTQYuR5TEB9gFZqB3d6Yo2
5a4j69HRRTRtJD7JmwwztHH6AZeyL2lrR2CQRhIfQ/QtyQ7cU1lSeE9lNHUOAFRLXPKfF2TjoSCf
P6R79pxWARVHMDUw2j7bZZkWInatW178Zv4gWxkosdHrMVK5ur2UsXu4YFFxF+iVM9oikuXsTtLT
WMiaDTdobI765z3Q4sl7eoVt3tvVYbpiL3geWCPR5IsIXVnZzuY5WoyrfAzH1yHCUiTfCjqfge2i
GrdXzudRnBlXNdTNgQ1CP5v4QwgSXq68RtNVVMbu5ATaKD8q9Fo18jmANnPZNnBpJ0i/dzllfJBF
UloLKq0JW+Qu7RAFaqnOFZrSwwLeeewrzmpp6rxwVb2Hb5o6ai/aSAbnkMC5k9iIWi4GOY1wxOkP
GTpfqmaZMf1ONTqvIwHPKbNlPc8adiEAbzGUsdd8jVlxgHPkqc9PVC2MGh6R1/zdSK0cobwH5qUe
7r9eGk3bXMHy57iS8BKHZGvB5PGdiOWH2BHqPd7f6ic3feVLOTRL+pNm4Tb5x6mysZfdWdH13kWq
iXqzjX/jkt4FKz55jsNaPA/j/C8XMk5zQHtl7ARjIRApxvHtfSCeGZVHexAe6O7f8jP/ewYt2CZk
4MX9aYTGgYxOmb/8t3F3SE70U0R3nlGPmY4sRn6Hq2wu+pB7o4WNAKzreVs7+vBkp5nXlYcEZ9mF
4EWsn451S5HtRfuoxwUXZZdYa5qcnFcsdIHi1GHw/cY+C9rCkOlR+Z/ogCg83HImb4CopHPcPFfo
z5d8rJJ1h8W+B7rqG8+YCuRGX+vQK0VhomKw5Zxoxv1pHyW//+73Bgt8oebKDm4BBw9l1lVcMReb
Lu0baC4zDfkj94F7/065QS1Q1lbxXQ3XQXpecyN7ZBezWCk+4LK8smRCgsyzqBlJx29wuX52RDbV
Sy3sXhZj9VTbGUOG0SdQfYH8xIbN6oZeEohBmnNnVUaamFnaA9XXjAvRV3zRmKSSzyPAefo+lFFi
/SamD7aUUj0z12NiA3RkvWSZmzmbvgcOknYoQLEBtHjz1PvHKoqGUkjJrTk6Njt+nkHHenDwC5DJ
yUuGW2GZMWvj2f8Vj8phgKHQQmHqnE0hwLWVzgu8G4LS7bImFRT/2uGUqq5t1VoXERhT9+gEUvmg
pLAFxpzxr93CRv2yCcdFUDfGCfgggJmcnlPCddQNXHeQU7WDS4Z8CFT9+6REs+LypdceHCgC4Bds
q95Jy7zP3g6KiG5OHaOBZYoUVcUo4GaCnjsTZgTQMxLGl8kQANPHobWSk2zN4wnorNIUiXr7SzEE
0MxiZafLVtRr7syVYFtUoR77aM4MmUhaaxvxKKaPyWCKUblziFRgEDxnze9trx8DzLh/oIpek2kE
QeFJd3c9u5gbWeabFyBd23cPD0qO5MC/Vigzq9AKgTQ29hushzf5tPFpez6bWfT1i7QXScbqOeC4
QS//gEfDxc2tuUeCkT6owJfU1xQDufR81H6MnjDrG/YHI2/Pp7NV2/JfEitSWXRUzp8bges4DmqV
YQLmfYInf70URff9C9YF+hrLfwUPlLanO+scDS3hEqIXN38pZhU4ghDPKHSpgXJErNN94bayeWhh
vw/PtEVpUii40DoXie1/Mq8zrG3pJzKs6ZmlQoRHnsNno5sxkXwXeGB4IOTOdxpR/wi4BcDEtG7N
tsngBzQhoZwPwoLA7rd/dpwqF3+/06/nIo4qoX+DJU9LWAdHgJ5hk0NaYJtJiW41KDZqzyCoD7Qh
rJ1D1JBuSGeCA4zF47ddxP7e14Vt4BhACEqUf92t2TIdlmtY42pStJbn1DsFxWCX+AeU3vTCFQh6
orf5+W8jz8O8kGhLHWvvUDGKCaeZ/ecWVRGrjsfLxitVD8H24u5Ee7w4fqWlOXvmTJxSXFJ55kFi
73gIsRsVGHfV5/PJGtxpNqlbPIkgGjIKEqTaY20H+rSqJja0ClBxGYDf5nO8P7EXcvbMz3hxynJp
z1FRwdBpvZQsbIeZnkWx5eMfkszjxeXjaJKAZ7jd+SYnUbmUml58iR8U3tY2CHOVt7t9XhdZQJzJ
Pcgt72vB7PHQiCHX8lbiOjAL7e8l/6QxfeJkjW/dKZeBKCkq9W1zYTjx0zS1EV3tq+u+00xMnFpK
zo0viMU2DbRxP9mBS58VpqoFkBbCaQahc1Qf60kQLqlF404GmYQ6cGnnszBSyoJBvUPnHaxF92bY
PZ2s9CAQ7QYUbnKiExANjFkcEXVzvhycDJyFuxXBJNml5Cd8tPmYoIqfCiz5HSVUoPz7okpMdfXy
p+o3BOzN8QhXke/YJIyr732uei2VWyozucXpxH3tYOOlMCYfJh/Pm+FTgoqeXhGjwlbDpGMDUTDd
1o7rW67YAV/K5elytIagG+ZxgRdinViQhuSYYOndTQK3cf8Nyr6ppkYFweb53k3PfIz5nYCtSf2H
QSYRbSSMXEdLX632v1SB0iy+aNU1yI0KBL75jWJnJhNGgdkGpQ54QgB7gjeUyFMCPsXMMHt7D553
sVSUVn1OaVtEjb6C0SMbbl+j8SX+0KLmWAzzPl6397yvpuO6XP+XPuu4BpRfsf4Tksri0VIO7kFd
s8s84OhIRCTmiTsfplC+g6kJsG667GsEDzTm2sHGmTM0u9MSG6ahnZoQXSsmVjVBF3/uam4zzHB9
1e4lkebJ0jjLGVu0MAaEQVBGTiieyOF9p6GY5GIjzYyoc9VydvRsRj/ABb0087MNBCEVIAu1IMzD
dr2SrsEG20R6JgvDnsohWZOl+ZiHZ8OIdN4F+zaeVGw0qJfBqSEodO9t84Zb8xmL/Zuv5b0liFak
iGBuALTrGoqDyDTBEWeNKfZ/KsiohngW6ZSCZc6HJgNAiqQzsFWERFOnq6g68v/qiuBoob5sHd43
/ipqsmc4vQ5gA2mhBgl8FJ5JsXjoZtxDBaDJx2FZD6NnuHtZe43B4/iWA+d4Gg90AYNwp6INy4u2
kpgaI2/8j4+XTWj2YsIgj8Tk4YCbx3qoNUGX4NAIiGZBigXNOw6aJD7YcSJFqlo1+zZ0zQRgegeR
Xc7fwkhqJgNCYDPq6s5dwRJDg/E8ivpMSPk/QE2MDyWrNZQ4CvfONYwaM/6nrrpgfxSX08rUJhji
wY688zHouKpqdQ5WLhczlXUY+ellxDn/1Wg+fRohzX2Ngqz3g6G6dTovS7TYiT5lkWhHyT++lget
Y/EPBUmOMrHvMyzP0ipX33Sw4i4DhvDw/WoDoMoTEAgsCjNm2RIA4tqWePVLq1Q7gZPnV16g+u7G
4TXH684aikLvbIg2JShJ1cur6H3PwRJPaHi8hBvkqn3+bA70bZIV+poEj8M+1ca2yS+W8luhJvRH
75o9Me9zUtpu1EhWpB2REyUgd50z0NpGUlO+GmTOQ0qOVXX3zS6ke80ydc1XObkYHH8idkSWVDux
n0umu1i0rf9hZhd7AkM+Z79emd/q/omSLMy4xbwwpllr0HspFgPrcHRb8stuN9eQwOyvj4zYpVQ2
RQbFARntJoXWOq0p5iGJMuZrXGq3QzXz4UsqJ9cWri/ta/eZrM5vBUQSvHDucSdzsH2Iw09iHAeh
S257e3oLEAXAGxBx3usk0mQjOpeV4iMnQEPvWHfbx9+uNLauIjxb7e/oHhMWC99OXf+drr8Rj5+e
WY/uQ6Wh74GbZHUBoqoKEDeJV/ZvLHU2boURadt/+ThXJ9cU5NaSHCthf9n6fa7TwcRpm8d/IUoc
R5ddIg4jeDXvG2ZhkJxdgHG7vyjL3jLJjprroy7cE0EyYezZ3KQg+qyccuclF4HWyr92EUu1ASS1
UNg2w2z/pTKnZ61ifiugSew/RlMdHAGB6ZLTtkp96Y/J1s7VTBj3jgxnVQaiGxX0vMpxa1jU3fHj
AysYq1vuJF5RAuOM2uqZZD09SI9tSV3s4flM7oRef+O5zlGpr3y2/5VRUCe4rE1TjlN7DHN3tC4Z
Z0jyVeQBAZb3oixpJ/iP2tKIII0cbGulVx7G2nPBjhQc/l61zYLo2SS2gMMSR/MsKsQHRFLblID5
+wuYgIT2zvBv24bNkRrrYQhl0vXM2NiatIohh6Np77EeTRr9pg7JxvHtvUlQuO5Jg6coP4D82Qr7
e/d+KNtR/1TvMavi1KRL9VlIYmi9JLHjPlt2KkFMk91MCWMyvQV+2NKSmVSQYSnn13jkRialBoJL
tpXV13sCcrQoaN0IEDXKh0/PtWp6dJRK0lhPs3OgDjnj8qRx5Isx3IA9v86183cR6a74yxDzbUK4
nsxrBWa00q1YuJw7Ew8YwEJ/8szYmbeyJfCCmOTtGWVvNVQk6FUFOWwtgI2pKVuyXpME4qPhAafe
YBy4h7cGPD8XKO6Kreh3hWRMn8cyV8mz8uwb8gdcRqwLCegAUPcDjcPmhaQnEsx5kDA4QlESncPf
GG6eLKTMmWh/QYbXzpEsey/ppaYF//n/bKCLDNmU7LsvMGezyg5Bf5/aF6Spgx6VERAct1euzHCI
70KtwafaSymKza1JJ+/Ku8qg7KtgfAb8bcKLZnH+sx9EhQw5l9dBMMSbHLJHFn6cFXW8oN2Xajt0
IRS/LrmmYKynun5I4IzEUvAHQcmqpmGq3PDQIv3Qz9iMgMvJUyHc2hqIM0UacEh7sPqliFdq/kov
GGGgA3a1ZDusVgn5AA3usX27Z7V5oRGr/fZnT1KBphYe9IOAXUlagnc/rDjsIPHwUkOGP0qWGucy
jRaXQNP+phO4iDx6vmI6Gj8E2gSiFiNIMxSU0zfYcbTstUYMAsdApjzKW0WC47ojTSaHFeIGCil2
ks+tsBE+QreMhely8l61GeHVYGG8VPWV1z2gi0JqshnH4oNF9NGLby/nBnVY2QC3Su4rIzqNDvQv
B3jfQ5fg89VfImrZjriffa8jiEUX+tNe8VjgiELmIVgj3kE6/90Igbpc0KQ/QjZQlW6h8VA2WShm
gEFF33a/hFBgGYjUYIaNDBn/UvQnulsxysN+KBNHlezhhVO2CCC+CrF94Uc9wF2trImXScgG6063
l+WCcuccLeITt7Xdeu2cfoRe4rejlDyWSWTh8fMT0pwx9epL18lNkyoCFt9v8sBLpiyY/psol3j1
mob5ldFmXBiv5GRJyDmkrXrpW5zfB0fK0Cwbc0rO+m9Ou1fRtDSPIiCSva07aWbcHxzA82Q8OHAB
15dAli2vErq/ZTK8fceJ0O1a7Gx3c5baSRM/0z2RubxYVIEDBYhqoVsck/8zbfQKvV42q/YOAo/h
348D61Mal//BsA0RuWIsTLeCTl9jsTzDKujKX4NIztUGphS0busvZ1BSjsK8HBpDa09BkvP6zH9H
hIr9yM0+23VPLrhODMc3Cb+a/FYWKjcgzqUnRh8PQ0aoE7JxFTyS+jb2AV4Mot+3XqpWIyPCRWfI
/5YIHLlO2Pig8inR9f8SJJL39pSaFIf7VAJTWsMu1hXCvNVCjuXEnNuqcthIryLXMx/WuGZ3Kz5p
iUddtKBGKmVce4FL0gfcFEeB1XGrcEQpeZhrBufe7+cTd951Xo1Gkdojs9FY85LilDv1C3WEt1EY
gw6S9JihV9+4CozA7Bv91YtBx4IKrlhAr+5Y3AT8XeoYpgz9ZiUUSWPKD1le+cIZ3anz78t7oFVF
WanpTHaw/IwtCYR/m4BPs1inzf6m9kuvON2waJ6OscYxiYA4hyIUAP89Qv82Je0E6/yD5zF9hjXc
ftKIRBfg2XF9jEticR6/KrjNVhQ/F12zsBliaxoRMLB6l953FRGvhCWav5krsszi6BN2eG7IB5ju
3HMxbXjrYTKw6bgryLLN/1ofQ4c9LwIP6S7F18L6YBvKuFSgPPB85wY+G4MkHV+GQfxUXePjeJQM
c8Oi1grt/Qx/bfK5ULNY+Qpem5Vslpjy7hvTwlU+jb+gUNJKU9xZ6PrLIL8yDokg6o/JDWsL5NT5
Q8SgDzQprGw+R10ue4gkyKj+NgDr6WFOiGfTnWmXGMQKZ/+99snLNAiMqqdvSGUDgdyc6g9ZuXIA
qJ6DQMrhWxuYtGl4lsc4Yas819phiFWZNcL85jXe6J93szZ/jzj0jjJkbJ7mMqPiwpTAHgZ0trYk
WReHRkEuOdUoMdKSsa28LNn1nIdd/OBoLByIJzpCcln7SdvY0q9IjMhPeAEuv+jevTZBd8CPvl1E
vul4yFhTT5aAFKq1ebgRK9u55iJxslrdbDFZ23yBoXBwoQgJaMNfQiGNcY5QSaAFOcx9A7m6kgPW
Gux7e1TDsS1T64CTIKcEFevk1Ye894iX+DTzyF8qQTJKYeGocC0gs+Mws5lVKNnz6/IrOd+GcitE
Q6LNTNZvobUxWev/78Gc2bl/xrfNVniFeWuFj+EN6+aythfgmAd2hjiocIHKEbR0rbCF1C9ANgBj
LV3vp9BxeZks40K8JyfuR+w7SAsLwn8xsHpfVjIG12+6MNaB17hdcSpRPq5ZsVKO29FjsZ0FDGEf
oKbN94/bnY7fwxy2r2oZrAQQ4H4s6R0668RfqEgDNVfvG04Oeo+xPVl8KdYgoAE6dG/BrzoAtEkh
er9Q8slwnV7tD49/K8ZW1U4+JLCzPpcrCvJVtdPz3uD7+mM4wYTUGepyzDqySgRNFU8JR/odvpRU
DSICQSU1UOr23OQGbn9zQuQ+Popglkv28GycH9K4arff4YM+UMWXZbC/+yPESGmlAAwrQkWI+QnP
scprBM/6XTKvDDR7xzc4lb5lmZdTwVlOoJwmaZk7l1091As8TlrZ8B2KrVvvcSls4elpiohKC9nF
PlYf5S6B/nULf/hlh4aDGPmE4tXKhrRqv9bWzPITr/GYdrpn+k+IjwEGj0V1/sdKLitwGUCPP9UQ
Th6Ixgd1zZ3xTl2iarA4cL0yl7XhGqbeOveQ9Vh5T/FI5nfqYe7vY7tAvMUDzZ7YwWOECmXvSiZI
GdVSgsJnz2wSA7r3svjN2neORzJHG0ZE72agFM4WnhpbolM6sakvlB0EjomqqHcdRtXFbA2EAcdi
/f1Y0+fT68qZj5NlVP11NAXY3J0cmrelN3xrJJC3TyEKpkz70CTDqR1nexzNeqvp40DZfamYpvkN
NSJBWZ4b7vfg5kARncNHwuFZwGTpTnTd+bUMcjfBlAlOTyu+aArcvkLiEvtybG1r3BJS3Dl5o+Vj
b/rhROOk/7Qha3Uiqu4lDTotfCC2xfful99tbcFWaJl/CKLe4usgQVcpmeB6LhOiZM0U3DQicMNv
eLxekIu+2ZHqxAaeYFJ6rYjYCDCdO4ENDePyz0yKEPoII46b3JdVn9w1ozMfqHWuu5tPsAjjtzjv
wp65cF3s1YuInURH8xgWErg2JnibJBYuaRkTC6X12yPuGCTiR7P1UHM729E5GzUQeTXIvwVoGYQ/
GYz/GjtFgak3oa90AzHKYuueXP6lWLUsZ/c3g0GEDPDOorTNlFOB6nW+gI+aPtfYvqWvwTIpoXo+
ww8p8nBKDk3ZEjQp4VOZA9uiV/Np+ltIpGVR1EGbaWcyYbOYByLQGGUU2qEqQ3ibGIxMuwkuloj2
Jj3kJG91GfXb4XeN1lFU9BK0iizqvS4qJZ5UwI3hCs/DwQrmKNCIVybiUIU5LI4brlgHk7Jyx89Z
1KY764JAgJcmoyJ52hCyt8VPwu9+wgF3yE8oIU6OvOTAK+UhUIULCnOa+k/KOg/b4BLsLChJPYsI
mvPWz3D9+lrcUQcgMKYgEbBZQSYzy/j52DghQoui0hcRetM6GQApPhJEorA8D13y+76CAV2eFW39
qH3oNOT4MNt3nNLkjdmTzyetOEk/LvAXlxsA6MD4P+SSFUlacGGZs5i86kk67gXs0dY6QwiRBmx4
T31QvlDEG2qVFh0wNuiHtUBFek9njJC1+5rHVNxkpVL9f/G/5ZyDv26+/K/7KqSKYfa67DILxcyj
93tDJ23AxAnmF1SUyc3CvfqOmzI4bUETrp2UaFQEjVI31YAXz5DUHQTbxFTutVAR7WsQ2Zvy1AsH
8REfPVHMQqsI6BD2KItTyTGoPiZF1iyi6yU9D5wjCuxeEwxbT8NDFV5lC+QwMMOiEpRckVKKqlef
ETGEESDmMgk9SPeYVwzR6Sa0cbMDdoxthSf26maHp+CKAqINuQXJ4VsrDxjRu1zebib4gCdreQHf
1JppQ3AA0D+w8D1v0V2H58Pg2nE9DB62J2mSXCdcbN44eDFW085WHjyLZVCkXbjFznapGEKnF4UX
rkiuKSaE6MHsOlzo5yELNiuq+hiFDIQZJI3AY6lhNyzcBPT4s6fHhtx+HJbhDXmtQY+ab54FWudi
tcXnnsSfYMAz4M5KzzNHO7nlCpSNhtb81fmODyx96L94nXkO7I7SlEqQJPC5W2WHmq25LLEUO88t
ycwhqswtxC9NzoIusWElFhw17TNTdHupcRaiJKjvPsGu/GJRGCcan3eLWeOFcp1q6xLZCubZYf9w
3+LmR08PicoYlVIYeGe9LfYOB5mKTEavd10L4JsEKouZm5E0WWwX113mGLFU9RmMywsx4+BNw5d6
qFOm9Hn+jnWPQqSGV+4f1YCQxLPcW45Sxhu+SJzF3hclg4mp3g7o7JQLjS9SUm+TTphC/fXntd9D
/boz7VJKx27f4FI/2Kx2/H5IMWGQ8q/+BvaWXytQH3D+V/VzyxYJyyFXDsra9D31/wN2K+o2kKN0
pQ6OUBVKuM84/TJ5hkV8VkhO/E31YdpkEufi9SPy2xhP8EB5AAir1Zv88w7Pkh+vqjphpVxsRD/t
7Bp2PSzc/6OcY1tzSl3kq93b3Akfx/jutY1A0v2ToY65HmHKwButeTaMfZKVcjUj7TjoCB3CW6W3
fwVqfl7sEIvkJNzwHdLgIljSJUPN9Aryqxhf7fgO71o1266YYAFxPoi+001itThuxcCtHQ+74kCi
gO015f7yUOIiJPLWW3D7R3kTyGUOSurzHRpkLCHvwMf916CP85QoM58WTzS4a/TJKduvLmVgZmuf
VkTlePQzhyMgIlJnLwQh8CaUwmpoNtW6rEOxumgdhglZvtVZzTPsqlsdeUZUMBNzH3o1fFWM97Uj
yfLnOBv4uksw0BlBYFLJFW2z4jh7Q/yaeaDJkktsrIj6/l75HQQv1ytK1Zf5R74Nr+qUMI+O4l7S
3gASyPnauXK5X27ONPmTV6Dz50cSa6J/3oJP392YffAYBFvUPouslMmUd/8EXVhK64GAFru21dwU
ICt5ZeTQCwWPwCs9QM3jVhDV5oqLKmAgdOc98j4p6vL/U0v9yoo1gatJmHaXtjxPthKEhJ6Kw0C3
F1WCafnZoYqLRaswYPD9HOVr7P1yI99HMV/zW4T0xrjfatasT7MgbUt9qCGnoehlpSCl4LBGOivf
UvOBvQqWgD/nupbsQ81xg1qhbLbkA3h877ASlTM2Sm8r5H+5WbQKM82y5Q8ig25k3vXt2kjWaFwM
+EvAs9uP1UTkC+HZ8ildVXzS3ynmf7Gr+IhmesEy6PYM3os+2NDHtq6T1NQtWP29Li1fBG/76H9Q
tPGt4J/gnUvBYo2Ze/OXRjPeX+1WZHA3z+J8NwJGT7oUFlXJaMyRnTXYfKqY6xMTr6CbrFIDICca
LCMa0+UpOVp5w33mbnZO6fdfUdc+Wdl9MoYi8/JWSTutxiOaQR03vRgzLgcVanztH2XolzYd+r9k
Yqb68NOHT79uujF2Ffd66TVw+KNe3ysX4cSuxl11sfdKZ1v8NbqzxRGzrg/I30Z+PmHApw42S0e8
UVj4DYYFMFq2TBTtXnj0K3tHJsc2IxI0+Y+8wY7wlr+F9vXRJ1j39+007RykLsM39wisYD8fI/kp
Y/N8KOFrEOmn/JA6/+225GMiGvcfVEOXfy5bTXC93qQp4Zp1G0RP7vmV9eAGdAV/K+pFz2MhSZFm
+3ufCU+noNg37a1uu4g8RCw7Rp/g1qBOK7ifW6xZZSCfUKWXctCgpctDbroNI1W7DoS93Py+MNSS
pFWTmZEJu3sqNkxSoFQm6eQojWfoIgA/3U8Oc0uwFBFEirPEHmKRaPWRFREuUFIxrKwFf5ujOlly
a4HUAsJVCol/OPtawbC4RYBicaVXO+xGUlxN8kno6MCSCJpP3JWHMbdiHCsAs4N6ZiwBv0YW25Lm
kyaR3h8j9BZwlY0+Wjnp5OH9ytLEaHoaV3VJDT7UYsjdvb/ytC0+jY0GKEWNFd+OQJHev1ZYT/Kg
I1lFZf2JjAn00FEMukmh0Z2T8JSs8S2BjG3de3zbAH8xW3wLfBpVO8dZy6pF952Ln52MaZnPrHKn
m/xit/7KBvrDZtV8D8ntBd5gN9kLfxxCUVsRAC58o5co5S1wdsanlPQGnnJt+U8nIwFuEfv44Zy7
4jSnA7P9+D1CpReJBa4drb3B6n8iHnyGgL99BaX+8fXozXwNymXkYmPlWZ0s7Fc9jepJ4xKlrMQ3
kPXD8rvgGdNb3rXbg6KDXb16TIL2Roi3l56DrpIwDQD/2JrnmyDm+QJ1ix3oydAzBOjRF6oD/oK9
foNQXsOjcXP2ZyiJaP1aXWg+fkwEWJLC1C06YEQtVXYPc+90UaMl6+JUAUgvOSPbynITFckdk06Q
lZUuCuym7LICsGPMXlk3ix8KlozzzNOmYmiN08fwIqNAsJvhI4ytuyiC07i+lkHFEmSe2tOloFQE
ML2Xi2z+8Cyy7kXGDcHDWZL4MAPqRHXhEmCTMQO+1XHNr6Mz6DjRry72iVqdeFK/zJod1Vo2dVfg
2zxX1zD+/UOzRP8kY/bhyXRc7xum7dp0Vllq41JvexO1tP9nEbEnf3vm5wYAc4leogHCrbJVRJMY
pSqBFAudiT8qM7Dg5BA2Ukk6qMvYTg3iZBGYlJkZVx1xRrK9p7DFdO7BPmNIY8Qq42YN/j4WIoqG
Mc9F4OAUCYWvJ+Zmi2zeEchieEqDdwUqb5HvLIWcMbAdDUfJ+Z2ZeBX+54xfWclIbTS/paOhKuLo
Hw7icHnc1aaBkMU+IvTwO7MwywWJPQZwz50nSeVI12Q2+sKF9wFSNRXzfuVFXqCFKloDEfIFehAu
w9J6fm84n1vvUdEWlz96bmCxOGLed5HYV6X5vqDelfdCq80fgsA/q/cocYNVVFYFUGAfSon9IWZu
uELCkVYeVOpoka6a21JYdUWOADkLgyy6YjLudJ3jrGygngjija5teJAxqUU8VllNhNp1S/3+6R27
DJMrbmS+zLDzmobATvzJZJ+0iU37QbqqWnGYkpNn87ELmaTsd6ZgAdiRkVw/KI4zFwZhQDWWPSsy
ewHqj99JbHtSOOWz6rTzKrw8Qy3IiGwmTmlRLnXFo/9l0itDscrTBbf3fWnN3TGG+42+VFTvxOFo
WhNm7BEC3BhMnG+pfhGi37nra3URfNm8Z3rnPUBepz2nZkPqlqtMTk0h8JOWiY1Bg5nV7DVLPjHX
LqeoYEhqgC1FtiQ8ax6NtVD48CQyqaJSSEVDHq0lFYhgU4bnhhcKgo7PWH6LZnBQlHbRNGkSjX5b
wj3nmc/MQaR2JU/mj3yMXJDoNUz4HGv+JEgWPrd9TN7KUQjul0uddsGbUaxNtVH53fvY98Ha+YQ6
HaD6lOAKb5xXfmMywzT09TDgqxAdYDlThiUcO8JiKnq5cw64sj0HRcGj6a7k3InzDtKNciUchf/7
p8q8rndumohsYPmP88Nl85qahmB737BQgqDbw08Zprsav5EIvXPvsmomk58LVkXse0QheOPlyhVe
kAuAJE9ZcMb1Tp6rKMUjJa1Y8w85cZ5E88d8nPWN/kjB9nC25AmqQw37XevMa594k0kefJDWmSwp
gexOWJoMgw+YoZaltDRwwYfFIqdqZefQekYzGi1fqnCaHZ+BH+KgvX3KyCVu8U25E8lJwwK0nOX0
69nMEHK+poEE084p7h3C6TFaQ0bv4zt+o5F8gt9jic9z7ToNnjWFHIP+bjcdrMvi+LIUyv836Qhn
DgSc8GItmUZbT+pT8ukPaDn40E1Zoe5OwrOjRy32scccYqmACbNOZRoAwIertLVijxX3x/M3R0nR
P9iANNTNRLFcsZYaeq05SOPFiXSPPTrLMGs6dWct5x/l5LYULe+Obtge5CxtjpmWV0QexyXDRsAA
rciEXqTpmrYL35hm/xbkPylRbrFQ0Hwm7HS3y1V9WfO1/WBEQPhTh/yowm99eWDZHIqVR7lSLVyk
f6dIyk5kjN2ATKcyVy2sUdxSYPV6dLGoxwxkXiPVZkzFhPiD07wBDna6AEtj2Jg+hUo+Nu0O2bsJ
0ErltghNT8/0kCzsNaQH+wS35q38gj6HQv/W4K156xqxJGIwQd/zy83yw05NtMhsU0xbbwcZyuAC
J68oEYD/IOxHEIj4d/4l6ygXy7RMSUg1zGZTMr5p5KqZU6DWBaV2oIndhLaiemQScfigbTiCkma3
YV2bEPT0UtF89KtyE5ObV5Man6ApGAK24tgV7QGhiTVLSVWH1r4ls5/1KRNNGDHRlCVx6M55FAoC
lb890caJO5pgfY+nW9e+MELAbgnhGSPrZs9Z5MpjJW54lSFvABHhz75HW6Cn3lWu8pceWsjVJ/tp
HmDKLBREkEKGHb3+cjgdDQzfI9IOQliI2Jv+Jo2vNmHLntkXPBjopFuaXKbCNuSMYASrfil7Hxyz
iQm8HJeYEPtTLHpFxHk30e03n8/+mumePUC4TP8lJmJYCm2U0v5eAb9xplOAmn9rHwRxeDOaucen
rqc3iIR36Gtlv1usYGmU663nNQU+J3YG1X+Lp42vAeFhLb+FXq+6oWioW9LeYnvFlZnw/D0Oqvuo
AdYVAfYDjcLutFpmdRuPp2NrPf0MkfYHH36vdNW+84MUka+WkeuDafkw90C/BYJgrzeBZNeS0Npu
T+QxI3N6EZLhEbWoks25D1xl6eXewmaCZi61dZ6U5S0t31b8Ebfh8jOWK+PvF7DzbtRRlczsFcbO
PfJTBThpf2dtVt3MMc6TgUall9ApPWu2DMjzgx7R3VlEIT5nppPeYB1fGHzmjURE9q7fqm/hMzx+
TbGJIGehszGbHiTDW38hExdC9gqmJitqqdXPAXyA60ykvzFa1KayqZ16ukwENyIoJB14/AmSzu/M
HC7mqeg6K2jR4L1i3TwA9gtcuX94MwCaInOLTAtInGCrpGhbzcVAPDBYMLkJuyeQdzeEqglHsqYm
4jDeTnB+En3TRn7JyA4sT+G14s+j6Kb6T1yteZHu6Cpnsd+gpBgvRDuXhqcqjtK9uL7SGP8uXsDT
rF042iB4tXLk6/lb3c5laMu7iOyhfK72IxgLf6b1IlPtkk+ieSvXVpEG+G2NOq7WGJu/7/8YH7sB
PArsZce0a6g/RtxQ2M/S2JZsrmJo5F4Wn0vYPL3nYPsFNT+NxIfKK7rkKcgLWbh0mP34w82BPZw2
jp/5lZLmvMza/RgFXHwNH8bH/MNUkvVGRjSVMLQKhg6mgl7CLzA/28eOuYKdvCLKze8pUlrOrKxm
WAGpejMOe5Boqsc1rYnsSTP7CYfDabMwT4mskNyhnhUbQ/EgK/XX6++aZH2UjH//rdmcRpcOXHdB
tT1Xy8yrN0YZ6bmaZ3B8eIrIj1pSiZQ7jmANGWnRKxQckKyctpR6k69o9JoaddOq/4kz9NVgw0dP
bmgtEH5JFvAVeZZxNWgdQR2ogwb0hBbhgkq5xfvmxMKWQf58Ug7mpawPeMSeK26jDltCazlJRS5x
ObzPD3CtkR2+MBjA0t6fIC3jYidD7yHhOOSsid0wKvPXmSZcb52k9ctsVaWYoyIqZVqoXCqyin6E
siz4ubaV5QQko8KRlPjspA7jqFbGvRnJOKjA00E/9KztHMHoCVKWLcUezcaXL8W688U1feX8mBdO
JECaomwDiXRGXJFw06bLufHGMfHz0M7loS0EeBiVTJw/sMb5avlzUMzzrmsppFHclfzTz5AnZk7E
/tj72cuKt7PVzxQVrpdKRmeMtblNge12plC3sr8EoA9jM2utSZYA0YycdC6evCLoB62/zbHhmBVY
GWkOw4cAzaECNvFZZvS05JlFP2moPgbQIBG5R7rOckY/vtkLHJXYr9Cg1RVrkl1bPE6Ud4p31vRF
grjz+i/E/hzvsd74C9N+oS+HF6+VDrmYtqeB8hgu/L3fbVYvdsOZ4n3udwKiUQ/QJ2H9Lm8WpLaS
A6Ws6Td4eMH2RVDKBadpZubESxQDhTheeuJiU7qN4usVVagIjR3ejp0mu1iIFAQvv/lby/EeyV0F
ZmHk9TVYCCgL+qVb9F4BN7hJNi3sq8XjKH/TvQwF415HNEHMYwg9KmBJmuR418Kao4Xcg14hV8Qs
NVpXpTO8pUe5y1cM2H+icJintELQ/kTmBL0UG3myXmIO8QU4X0libNM1QZAAL+t2cXZBuRgcKCS/
+vw6vQMMhq+cqecF1mUp3hHcFd3BYf/5Bifww7jNfq2G4aBPAwwIrj0uCmvAqyWbccJBCalewksQ
ErRRrFL+cC1NEpLSOSS65+cZFBgaFPhJtqEiR+7JAhT+wZ2+QB9JvUXjvJSw6Fp1hjHTjtKkMuhE
t8ulgfezRN0P71ixgbojShKxDeHTotk3+E73h7deB4xHA9QWJ4rxPqBRGCVAgxINi1mD7ggCS8hi
jbTGjXrD1XPeTrFDAoK4RISKjgldln6B3n6JwBZkc6X16UEoDHn6JLpKl1h5wP3rdzsir8ttqJ7s
Wbsg7r/odjAMz/aiYsD5JnfAqt4SitV8q0gwhW5LbV/+f4bxJQnzntJUlVW9p5yE5ahRFsHgekKA
zRuTPfCxcRBoi6r7V0e5kxj6Y4Bdt1vqaBoRr5BJL96H+KV5aoacNrafs1T4bIk8dEAiep7D7Y3U
ZB3aKL7sJaiS86jPPM+F5BvPqkzEEAzqbxtFG4GfF+6+PwrM/b5hZnZCUCie1tabGshxS5uNFPbN
wdjO9dZg+cNt+tIfOskmN3acaQJuAiwEFqZP3DJC/7TqLJYVqGLYvyQ61KPPMUw1x329xC0CX63Z
KCNeoZpFQKsXgZ+wcOyDEzKqwaldCMR0zpKMt/AlgCV5panprPhb2X7Kp9at3cUekBATVVBHCQfe
SimbhJY18WbEY4RdOf4tPWXuyzf1FwI4aXRzLGBKmHEDkdf53vRVisccHddXrIrt6X9M3oyEfWuK
H8NBEwiC+HdJHXJkOofzghdZEu8lk1MZBf4Qc/sUjh69oPoeU++wSdHARLXhd+oI8GQjX0A32XGv
5m8CroOi4wsuVVvyOkxRvfxbRo4HgJrArJ8C7x63DaJjIqmn77/M7WIJJRwM1yz/lnbohsii1O25
HKPANFJ3FPcyAn0Oys0LnBnwVFFKoPVF2ofroCKOP0YInyb+hxYgPJbvFmpJ1brs970nwylCr6Uq
NbTPQiSfrlLh6tqr6GStrbg8X2Y9y/UFVnn54mEMyKzTljnLMixZnyoxbnKlyQlBrkdBhbnUGeXX
gtkXBQgDdK7eE1ChE65vm+DRrdL9tmCGFBIKCGz46GW/YnMKitJq0asZriM5E5N2RAd2LwntFKuz
L7aaa4u5bvm9QoWyOwpvxQCt4yyw2mBttvLG7b976X7ul0fiNxKQ3ADulMeIbls+FPe9zeRTPrX5
t3eSaMiwqkvcRGAfd/sTzoZL6npsA1AXvN/FMKg5MinmzsJy25iDttKQ0fNwUrKZyW8Mdmc/SQmz
s6rBKWnmQiyGBMMYOrqa5ORTV9tuIQQBmcQ4rCxD28WZ9JWzZcZbD/7Qda01h7Cncf4xI8bcZAWh
wx8gBmFAdUwQ1DlZ1QiYCqZl+I1CtzmpFqpk4rlXYtPrOMFROSets6biDPzS9Xnhq8kbVVpy+Iyk
L7Z1tegT6exB0djXDPFb4xIGwxOHPEkdSU5w/6clCqX32hlBlwz4ZDiZ6fTqbWSUJI1OzWMazMgc
3fO6uTfw3OaeLjGvanbNDo9XLZCQrF1BLUoAIWcW6j8zPRxEaIY8FAqpKeM41J+CMXL2PfXFn1HT
xj3/NtpiwpjPrvRA9DG1XBHN5RdZSK6sJ5+be2fjctYWJnn/QZXpwh25YUAEnanh2jTKVkNqQAgJ
6g7IvdQeXyAw3gXjF4eAgiRU0i+qVj+1ZRDhQEHkRbDxjX4iy+TCAGYeKNh398w/f2ZUDE5ASmLc
bz6wVfQFiOh2IwkSRPtqaJFCwaaOiVuM3GrlPQ3QXrYIG0G7tt8EssorzCa8RYfFW0BKKwXim+kn
zuWeE9O3eFE0tWPfuohwzwQE54wEglZuTy1AHHaRudTM9uBDMAyyF117LXdRsVe1nwS0rHWYcrGB
KvFjwthx7p6Pr3R6qcHkeKSETc7xLDkTKqav3Lrm4E/oorcaLC+U9obi1iB1wNFnQHppP6Vf88lj
lKgya54xNw0DvLt+V6SEXs72XpQ5FopWpCsg4WeK1DQNvxONqH3paAX5OKcxJyWVsN07DBHC9cCB
+/1S5ZvgXbcMLAgiudT69I5MWfUb85VljA11JQiYjzlni+od9HsI/mpLui/GHvVXdnLYWCMrJncU
Zlan/7U/nODe1PVG5OboosmqI+ETCIdo/WnqsZC11iK8RkZHVDNOrk0sodJ6y9roPF+O3Skpg0ko
swewlWiygrXZ6FFBpgXrmwe6VCcihpGWEH1UJYwazDHTXkXuTbfxkF9BWRfXe/8K/2juK7dvWjMF
TtNCCqhUJHQ29d/NHB6eDyC51x0criQH0NRK/rfEM0zfKMYVMKyN4IYJuAm4gdqqsCD/Ov4HWe8o
0Z+atV8PptvICBoRBOXCOrCDkEZPdiDFnlhtJvw9YCOYXcL5BGwFucxpTG4fJtUlOuPY/u7bLaiB
ialqzrTp4imAfhHdZSq6JaPfS/SK5WcRaCxoOfYX5jbkMwoBXkCHrsr0ZOCUmQmNoZxeZ733lZEp
TMYV6dhP/z84QUtgZcoIeu6AMCidKGeQkQFezsPDP2HAVhgLekqBRDNFHB3rd5Lecd1md4w7DDYD
MKhbm5N1EBf1Qp4L0mWQxhy1sGvyjalluxrMi/duoPUpVs2/TcEFVAl3+ykTkEo6N1UcCVoYucux
E+UJ0adYL9Cgu0pDG467txOcGzCYGmiM27PuxBWwt99QdFEVTJAQNqcBfEELlEkac9BM8T6LBulZ
OW8GbF8yFDOy9SNzs4VHncMflUWsYqzErgLbW69VqGVfbT7/5Mxl4xvXp63AoW09leGHMsQSVYtN
O4wRCc8GKs1kPEEEh3VoKVmd1dr4kdOTO3RiooJblLN+IqpSdGzG2dWOXdNGZyODX3Ykc8WSlVaS
TLV61dU93jFA8m3He/O4l+jLjJLA2GLuel4ZpcfAfhmqdBsjQwcdHX2yi+hUtw18Lw4jy7R4rNBn
RqrJ+3hOSmi0m2Z/OHyISO0TiOsVYcPfc3xLDO1H2zwtBY00PnT9kXheknwxrRrFnB0AVGfxaJ8c
HVoUHlE26PgBzkH24Kr7Udoy30d1fpEl7BijDGa+KdIxaSV0RQZcbW/K5InKRQgqSsUwKHW6MB63
p58grjaD72omv8TIHHcTH4JDaLSR83EfYMdvFzSQoZCRc9agQWZ6PHYVl5tKUxAFbRzax2Gp4Qxg
7yVlpo9oT+aux9fQRzrr+NgAtWTEftbTwNA3dV1cFleaPUCu6L8HQA8mwalJD/t4ps8QkiVPh5wt
T3vSYOQGvfPtPysHyyH42pzdnb5sO6PB8o7LpWPfJj6joY8ERnd5qdd+AJ3vfxyNqRo0j1ORQcOj
oVEXF/bVkhKJmWxgSP7Q13OIGRLMIURMrmO1hnnhTmNs96ibJIE4452UTALhH3sc2a6IY3MJ85va
bDhcxjFnJ7OG/7bOszkRiZWrePaF4Cbz8dUE37guJOeAgj7Dw5hCm8ceo/3eWiZwY42e3CZWR1l3
D3z6Pkjt8UJQQHcqlpsNDSBLBaOr/Zo7y+hYo2MJY1M2l/riDF9Q1xSl5DaILNV+5vhRkl2HK5T5
cvRtOWeQbAvyVk5Ma/1Wdqeyism8eZTjii2eXeJwjvhoJbLj0I/OO0FO5qtL20QBS1ouXNI0pXbT
MLMMCt6+XNHKS4tAkz/GmGua3tbju7LyWfgX8yb3T7i4kJBe5UC6R+KX+5J58uJPQAFGl6KBKn5e
FGM3mJ6uN9qG1M/ShoqLe0ZLd97RVoBbe8wbwGjxK7RRNW3IAC9BswmRd67XNAmvMgR7Q3vk1Zq9
GHf4F8F1sRPxPvaRlaVUvzdjQ13CaYFKqA3AkByLGSA04ga6oBWfhEGtGB2Aud+LdyNj4jyMiFSL
3RCX+fWGahnhDC6eDDx32y+5Pos4LrIeI3kYDTOa9iMwX/9FVzff14CMKWYn5UFnjSMNxA4mKAZy
VGQik0W972pcFRPj3vip1D1UigqTq7reAZEClRCLQnAFsA0NggTP8n3GBZqBKBBchvK4+6cVV5RX
fMnVHON0cQQ2pKVBMO22MjNHhO2OsG0L7dHXDIGAAXz0Snd664ddJPXD1KAf6UJPIS5t8P2G2xK8
Ch+x7NRZEQGnv+ogmoyLSD4k12Q+lBy+rEFrJIZMBKt2RifzjQD4WpcWCaPUzEWrzbouo8txPrgZ
xjyCWfIJpvkK9Q2oxFT1ahbPXPpENlSUvkDxa1Tk9UM76qlv1Tk7kYRgW6a/J7HwOzLoNp937kC+
8geHS7TSz8NNvdFrSpWn7z+PUjAjIkkZgdIdFXeM6wN0Ecrx4IU7rPLntn4bhp9HAsu8FoZcAoE5
bVtQNBox4Dgi33M/OosOiggkX8rOgo5HQ4jzl3WN7pw4l4uVhYuTQG70Tf9PiC8K6e0y/GUN52J+
bJxk98USPmg8vMwtd2F1YZTrznRZUAgwS9bZ30b7VbjHkH2p80d7uIWh+YP9B2fbDFRMKsoN9I3C
Aia1niobYT1fJV21olk5lL7e0XnsEtuMTbqsiGEoAVZADbkNmTcW6FOyzoFSrcFdk9P1pwBouOp3
GlRpFIRQWIqSqbECdQrkZdnFQueKzTikmnrm4e4fYlL+sryq1FfCwwMRn4u2HY6OxS0+1Z0oGWDe
E8rwVyJ+ia+ySbAEPv7NZft30JKS8LTEy2pdJfynhEY1blAqe/Q7dXD30j1pl5+kGCHbIbjak01k
XePWRA8B6VlYRgMDFdyNxwPS6cFXXyBie9v+Pknlen/B5oHd3m47S68gBfex27aMRQwwWAGyzoB+
JseQ5KzDA6WCciFjVYHVvCLp9Uox70yDW9TdSJ/m6XJpzSCi1DFssmfvmacPlfSHYo8QoU6PT/gj
5IAC5GnEm4ExXpGec2bM9WV3uDtWUG6/EDdxM8FfD8XPbivDkcD1sGd+rz6Fg8+LdqKVI9vBdvBf
3ICn7pLQKLIfmNB2SWeuAfFwojScU35Sr+4JObNUtoB3dAYijS+7+YlxC2n0Q56QTeeXSwQVC4eV
ovshSJO/EwZskP4P7UmLFHni5MY4S82zEEPsKF8eYKIev62MkPNzZNWECt2pkjuKLoHzzKKWVOgD
toqZEhOrk9h6U6bKzuW/m/ITAaZlUunOTgQtYvJXGT9NTtM06W4Mq13v8Yy0Kg/uZ4wIc3mXC7R+
Ga73FrUpcdzYLYMiMf6z6PxRGNMUTLjNuqZ2ewdaUbxyDg4XT4+0GD2ZKKppDZSSWeJb8A1HWLNA
iHBTX2zIRU6n6mykffSMmqll8hCkj3+2Ukqdz9hA5xpifSzsLaaJzDBvDv5DJMU+/uJhzyHR++Yz
Vgp1weBndaOTva+R87YpujEQ5HWCtiIywkCLGTjYrF9cR7dL1zJjWO1FfMkt9xUBinuaL2Cl4t26
cqBq6NcrN+jBWsntKRNloeHJ3D3kAWFfBcDKt8LhGLKdIFm4sY8Eg3xhxDk725Ihf/p3sXpZXAwi
rOB8g6s7c8pQY1ECCayYa8xkdGeXwsV1bg6knDNRUe/lpQWoBQdYno6SWgXlVelvBJWy6egHFT2z
dEqtVjVsCbWxI+ZMVkl33Lbb77z6HgwqFy+6I1fq0usgZMEl92qXMM+m75Eu5R4bd6eG5W+ffuhX
5lBkQgnPoBZw67H9E7R3ObTElVJHnos498UHpbqFLekG+9/57ZcoUOUXSuTO87E4qZGE9GUAzpkD
WcIz765hXH/x6QAAyW2GjLKjgtTyTjofNvryV8cA2YsjKVMXC+trEwwbmjTpOogeD3bE+s2K44H+
50ENrVjyMRrH6lYhEO5RIuJzEuP2kSL43nIdUCMLmkwXtLoDHnW3Evnz+gEpesbnE1rhkxcyvuoa
1hav9fIF6jupmX67Xr1UZnDYWvENerRdVpyfamL/NGcylKVaffHxNoDn5XSIABDnXVFCd5b3WvFU
hc7wYw+6CR8AD7dJWuTJGybxW/1Q3Pjd+nHxOqpL8vLA2USkC5gFtKKIYHsMD7NrSW+UWdYQErRk
aB07Lj8jhCSJSlaORpd+83rTNPIVFxrXoHGT3IhahOMvvOr98NMrW/0E6MkZp/zCwH3BJ726poQl
hhFHDWkvku1kGuzqxgZoBPPs/YOT4ocenXahvuu1uzRJqwclx4weRwPcNmOm/qcT3CT9gUX8T9ox
PzkSXJtZuT9tHB1f3IGM/AjiMo534Ok+CR6Du23z9VjzeTCr+/hr+P+LXstXWN71fyFRnx8gRCB0
hKadsdsEk8GSyk0F7zolLzH+jZOBRnZjl6DwO2IwhcFcYty0mLnSPtPywypokMXnXUVpcaxwb8MO
kFoRAjwY0E74RrgY2Hc3oPP1deEsfSIUj712URdRj3Vbzb7n2chuzEW5SgUpnB1zwoQklcmRG19z
7PDlx1LqgO5cP66exRQhnB0BxPHqyNI+2BaOvajeAE4UgrTJF6DKQIx1pCBVBhp8XYxCz80JYR1l
wrmnOuTLJlTFVX9f+9LCdbNUuQsqDVoZNzifXUphaJC9+Z+5YGyhKNhnWFLNoEOEYI//pm7QzzGP
2jFryF0ho1VUeVlpbs8CHNoUGjWPwsdHGYCnhSbnx+65fMPalLMxdEbI7WAMD35K6kNIvy1INH1n
Ey22cMr93Ev3ZyBiJUFaW8Q0KJx15rOJfWWWepGSKAQYTPnPDBCDIPTPvX8oA6en8yfFT0NO0lU0
S5t5TJO+QOcUWsiYKpF+thycPitU9QU84coux7TAGAeVxl6cObbTMtsnN7o0MgrRkWf5jXJxM+Yj
6jWDxyVB29C9VeTnNlo1rbjzT0VW48GbD4knItbDl0ZqsXCkNrPIcizqpc6P4A4QrOoVenyB8qn3
lod8X83WwGGN3V4gsuFUSEBudncZsX2B7rx6g1XBtUazt+q3DBdy41QmM+k/KXtHyJ/uXTJ8bmi5
wyWEyDcnwqrma2gtHAxeB+A4sA6C0K9gf5L7khS6mb7uJBQvDSK0/3eiNq1Xd3j/H5DV3XVpuCXf
YjKNwrHRch9pxkIqRkpXM3rMZBQS3g/XTe0bxqHY/CX0xqPgbQjeKlCyrH2ymPhJtqm/+26/ycru
21CMpuuEs12muC7+xDRIX7mkC6MOD+QmkPq4gPxjDzhUboOsF3WklsKr8fi2EwEC8BAEMcCbS5tD
C0hNCWzFp77XoxPDAxTfij7EdQIe6eYAbjydD+olvfpKcPI0L3H/CbRR2nkeP7rIKRVeqveWrbxH
1o4gaMmaeOOue9hCCzActabf3i0dvTWLdeQHAK6l2HVKHMEPgDMQkTVeyU+KaxckFAy3K1YKD2qk
0VXlGPfm2BO0wdDG3adHNSEPC48/EDjajwvk5McBiAwiH8obNJlu79utUPNIMrMXY8fop/Ave4ml
9OoULK0rdC39QYYjV+GNQa/ATl1MwaQCpcQydfy/XjcqIodAgsANhLErcud2okklzL2wz2I6+XpR
cBW412dp7qLQx3lLC1JAcmoLlr2RYGLPms785S3GHgFVindD3jKF3FE80FuF0RuFU7GHEz1Grc+F
TJ7htfn5YZd5zGFjInjnuSKyoMW8wrYDjUHO3tN2MyGDj9adZGrKS8b+cVBXIiju3pHz0/4qQIU/
4tpNwQrVLmSSrmuglpoGSPOaABqH41HOLsHGaqAzRUWqA0jm9KYzy1EvqQ6RSWKE0St1MkLa540r
WNcp0yOMJhAQ1Ui1qmERx1nlqc+pRzxPbEp8LLhxC+13eBmRKIaHQqmXE1SrNLmx7EsEt15+sLlK
sFZMZp1za6LmP1HjlkxIaIcJu6/4+QRObg2mKT25vMQ4DHlXZ6hoO3+2m/8EjYMu1udaCSO5Qn+F
mH5KeI5E9P1WhqmlsHZnXpqXwiFgmoj5EW/OkZrcFAOH1zgkGNr0c/O/scuN3CVzKQeim95c/4bu
ottTJdGVxRq44vRxfC32PeJyXdsxS4SYqbiuta+y6DPVwSgxP19/suu53jRBJ4Dsyv31q6B4nhYR
rPKfIteDfanr/gxPpBjbFFsjbWiCKAILR8cBHjSiZVxixArBSM5UwLaHmTcNe/mGZuuqY4OotYVc
Zqowa+kdhjy2nviYiKQBSw/NwCurMKTAx6NMDFb1zzeVVt1Ewvh9DREUrbCXg7EoaVhnHAgUZwm9
4HCOBoLOQWDC6BROgvKp+8XJQefaXBnfJGeemnuV40SARwU2PaQWysi7+w1FZvtUMvEv9QfGVtML
1FmbuH1WoIpK8iy58Ucyc/r622RE7QIjPp78n1eCy7KClOyRtgxKJN6qW9c9KSwWIgqsxqfoesXI
sSY39aB8HV+WnHSRCel0FR2+SapGLZox0buaF7O8rZUqcrVoe3Maw35QsNHRbpFtloOYbr/ROi30
Xfij9z8QjAN4INquMPlu6UqK6fEjaOb5em9z3KtXVSnyRtnYgGKjqHTRKlLAzMWhWxNBF0mMQ8lX
CjAp1qu8fX/X9wWHF5t1mz3sUZ3jzCIaFofuFVBAYo3qPOCaHChHFnwppHld4rWJPc27MzoiMgw6
hd7ptgeziN3LL1xUrTBqS2aWY2kAI2Nd/gJGI7zLBDoQmOm8rtmRUEsu9en5KmQEIVNpRhFVeKoy
f9xbaWykrDoMoF91izy7vftYRb1Qkllnw5ls/eiqaLdbhJ62e2lFsG6TQUHnLB/cXhkPX4FziqEo
vQwE1e0sAyx/tCtGeuF/1mnhTFiN6gt1DEthAU3rSQcVMzpwHxqP68kvDmJfHPqocDjVD6/X3vey
6m9niX/bFe9vm6o1ZM59If8gurEAKI+/JRvKzrfl/Hz5gVmf/Enz1uXb4jbaFtZHflshPNq2yKNc
Z66DocuiOBnYRWu7CcHKHi5jOMokAdQcs1cjKxMJX9P1oq56cOfdu5DU8/1Sl7jw1ujLWnrQ06Eu
vM8pnrHQgd3jn8h88jBoYRooOg1YGWFhCPhm6Gl1wexNlcfNU4mi+2/XvMbIqaVYMWzvZgeqWlx6
qunvHdftKFYaOE6DWi3E0dkpYWXBOkdGHHAvONYc3beN2IQMX2WyoFS7uSB3JNUWQmrLRo5xXqAy
TcsewFkdOpzqTn+i+Cx8Scj4FZ8vuNRXxySz+wDIqaPH8Zxk6uS5bynoezl8tD5xI5m829nK/OxB
3dfR/H9Bs4NYN45TU5zWLiar0K9CMDvVNmzVXSplb+THeNBojnjMPHZbLwIHIpt/UDExkIezTdeL
xbLPtB9ft0IhFo5/IxcVoc/zEu3c/gP16fVwS6/dS3G3/5RCvQKrbPNh0d2SVLNVq4eOOMmnNtnz
nw8THAhEOICzRxThOOPQJtkTODobf9sRZZgnd+diThpJc+pF6+z54bIEyN5L/4wjGGDXSfnUX8Jj
a/KCtQyqMpg6OsfNLrg4Ew5RAyh/eUQL4EQeoNvqrAAoO0ZaEfFKgYY2G0neERXLDNj6Vv48dPkr
5r8KfzhXjl3/OCbJjxl7JTyii/DGkeGSC4E32Abkq9d1l3rWPphaF69A1natHW+t95p9HlQbQR7W
Qcfdu/6Lw0jVk9Ovu1h5kbM2CvYI/t3rhfxWBwoXtBd0422/c7FBRbtg1OCDSf+hrKvH21xdGLWk
EBrGmLzIvPsWHBcXLmfERjxVi6hhCqT9UBPZz3NAafG0WQoVr/7M3K3RsKGJMITwyY6c5KBdy6q7
wGueMwvYrN2MaTvIO8C9es6oT5ff/z/YBvbeVEjvQMjneARQAcFxL+8Vn6leTKcNPqFmA4PL05/u
GYAEcXHSS8IWwPkvkVsXlVm7rfszsk+I+io5dGnXEQiZQn64Z4FNY6voZdctqs3ZBYcuqzfs0K7f
2+CxPilWOvluvIX4FWa0phBzddhLq6mvrsWeFdmi2hN9x+D/NBVsMgHglNB6yIHpWgPVb7tmWOny
ZcIx+GVl+42jap4iQBvKA2FERAvyH+GKxqxGmlpb1UzkU5/gHDm7KHFDF99Pj4FxZtNU9cLcygAU
FW7nb9w0ZfmiXaXaZkPAb2BDQ45HAIqIBcoL9x/iXLMjiUiwWYGkdeXT1lmkoRVzIWJqc6iIhUM0
RIwHdXFG0twvevxW+VUNOOmCc+qw3VWemNONazeel7mLhnz9g+FL4AmTRWcC0eg4HmOIA2C1CCc7
nF/W21hcEubV/iOsIUB58b6Tri0Gadb+II13KmN6BMNHuF8emLGuDk3fZEOAMWu8h4AWtSkHI8w0
BBBjio90DWYXDfz7ERb6uNtTtcN0H6h42oj5i6nBpDWvhrIqh6tB0a7can5TZ8hFrOT27uA5jIix
B3nnow+HAngIh9HuURP8WUbCc1DYyX6DZLEDHKPGi9ZTISXqpgl3TiFh5pJfsUmYIgttO407N9tE
qWqVRmIAg8qhdlp3P9Tb+6h8zqbev/xnV1tJHaQlCeQy2c04Z3NU+wgvPrtXQ5lFPrqeYNyRk18z
KUYOkY4WEROpiq3kauHv8tQ7RiLLiFkKUbxgCtN4FPbPRAFgZiT3vwy75QIkcnJj/Gq3+WGVpgbZ
nJSJR/VQynMhEeGdjMl/BsGnj6DCbe1l2/rP352evg8OmOBduiVIUhC4Ly37Fa/dvyTzSqcOyANp
q2CCtrEE2x0ttfZeVEAwPycObruupNZmbtkRFzekU0FySEMih883pGLLhKZSUrzGpt6idM+HJXNb
d/PaSKVUW3RQM33kkEQZsgmtQVOXJwwsESs+zl27vMhItpM3vXi7cGCT4TGuGNCbsCenWyayWnLT
GH2Vio8/4jXJm/BveNAC3ONzFtEVJ0FvgMgK/+TmDp6rfArNtH85HzGB/WSDrs9Y0LAENkPzSY0w
A1OeSR6xs2/uaT7jJbK2eGZGTYvmJ+sCiuBgbBX0k7ucenLHZnyFlyScopXipCqPHYXlHndTFj6R
lzxGX3v9SWLJUMccc35P84yiQ27dmSpEvjznPkUvy0yheeMdYCb2ldWY8U0jT0vWeUlpX67H4YO9
za01OIxKH0LJlzsYUssMPYH2/sLiugS7WYGz8U4zSHRpkwsi/9L4A9CiL+wGcz1umsbgSvK+c2wt
RtCfDaqFJUH/sg5wgmFusoxu1Ac8kpNcDKaPzZJ7q/Qi/JVlCBOSNNwEwRbMwjgQNZz5W/jjM78Y
WXem4gIb2EhRhNimy99ovyV7HWi0DR7W8OoFWJkAqq02ZEU14RKafwh14Tp8JWdsN12rWiD0/O8R
dbF5QBKh4aIsgcAnbCNBoGbuf9Q3rwYDvRED0cYU+wYXeVmCJfOH6S5GZBaSULPYwB/RYR25k08m
iR1xR4fWu/4ZcnmPt+tPMmq1/3EUl5SzvksXdDRBwtdakhkJ1voRIPvnbB9bjXebgzSinnZtXJzs
+8tdOZkE1js77D8iCN44DJD4YmXUaCQpgH7wdDMcTlYoyUTs/08jAaiQaoE2ah9pMYy4shvsdtqa
Kc/FrlRMAlQr4EN7AI26j2jods6BulhqgDKxwJUxlgQDnbOazVAp9fRvpP17aZnTW2lJDAnTBIEk
ZJ2ccOqnNNl2J3eDsboblnuSgQApFc/anVQxUb1q/32AfWbk3ah5C0zZw6pnNzGYCYXtB38gw0xn
p/jWe26R+ZttOkVsr8sz+WGioHBCafQQMuGVTUV/KemOGfdUtf9qRNTzzJFh2OkvxjvYWBy3/CR9
+ZZMuxiHRBuEY8FaCCPqbGaauigKRQTvKVsNZo4dkneCm9llsnWcOrcuhjLnOgMVaq3Pyo4blVeH
gCt/uDSzqj51v4o/S/obnC60Ic/l0jLTU12gJYjuX+wwdIt1P9oeao75hVom/LrXuZZTsVEmN/k+
tPaIhvz+0n6nuCXMoqqU52WHvVbylyfy2NC8OJv7NGKdhP3hJlNUgO2lpxaPqyu1iEV1D9K29SdG
YQKz8EAePQDHVgckxl4AZEphQsRPKaA2qUFltP0ICptwHmEOmonZvMj+4Ds1F8LcboCONOihxQme
zcqG1v5rCqJ0e3hJvcOVOHMlNTkarj6Xigr5lYo+6SlT3/2Dsn0wcrPH22nDge5YCMBttF2moBGX
HlB966pzaAaTb30aWwRN1kCkyJzrs2JNVNqvP4/JaXyIQRuJV8QIZQ9iz0nRG2svoTQ9HfrhD6wl
E0EATCPZJyIjlBj0jEoJkOUIvNw22l9qn38MVSVEhrBOVtu6kz91RyhanBo+wj405YM1ntlNisHV
GVeuceR8whKsTZH4eUw75nK4RG9MRrAh6iRWLcjWJf5Qflhd5TlLE67h09eHqk0XPMGaT4/MO2y3
gOA4fmJoI01F1m9b0To0wd4vWTiQVIWgCeEW4QaK0QoPiVQFbLQCsBe+bSWkE++DJRs9sOg3wQLQ
Mm4qQwPjXB3ubzl06DHO32UC54JtvP7yNbw/fWZPIFv3x/hmXeN6vg39CaAMBD7vzIwtSl8OERR5
GhMHleckgv+r/SVxGdlD0TM3abwajGLrnxt7oj04wJbN4rWzl5AtO4TxlYSWZFWQB+9Bc2hQSrWn
+NcwsUyWUbkmlw3UatLR0P4k0WDMYEwUqc6BzvTDYBd8anu9aPSkEUOuXfYCgsXkqx4YekzBbpjz
Olgdg94JnsW/RS5q9ig7YWmt0fNUk3xoHeV06EeHs7Stas6gQY8P1cxnaGJgndjVd8TMuyA71Awl
CpdYJvI+GiIosoYd4bB5dyYVhTeGFPiqoh7K6O0TNn7ikVhckr1/s79A1Y9EQZ0IRp2h0w1Jpxyk
G0JV+EFMaShiYrRFtuBXjOdzq3IzjibfFcEUW6vSI4PfTgvyTbe6qOWEgqF12VVTZjnT6sbzoIsQ
75qIysfji0FqQ/+hbDbbwJwSXjL9IXRNvmOUBFT7itfsncphrmcvG02U4D0ru56H+iHy+rrFJLac
WIDDxVK7BD9ByUUKSCfCYpR1CbtoAzUtzjfiZ9o/vwz8GPOoLqfJ7FP4AxjjMnf84RvYGZnAnWlS
DIp77o2fYQ1qweghKsoVye7wD+pl9FrK6IFGqYNzJTnlUNFDaiWPhpI3cRyLNGIBWkUOfidQ0aSL
4LdGzHVRu9fiIJFvOdRuAr8g9Sy8MTntA8re1L2CC/70QlOH1ni7KiyZm0RK2Cdu95w5DhykezF/
7Rf+2zgGcg03HF3pXXatXUE434jT82bRBQjNitbsJhIa3PiB4TPZEk6RHOmPkNn/f9z42Pbs2Bc2
Cl+cQR9aRKQXygKUF4iw0qIZsKyYl8ur6E+LeKh1CWx3YVwKIVnfqBbBuOtQs+nxpraasGHtwJ/a
YYlF5j+10UaP5tVIKiKxjX1FzRMczSB3qvCsZx9FQESP7dPXDs2dzjtMXq6BMFV43S64YCIxxCe2
QECziuZGHZbNcn8eAIOL2oM+2wpzYh+exIw7PMg5SM+lyh5wfNmt5r+zmcpQtRta2Zlvx8FtNyWr
eEcKDl01FdKyWQ71danfuoE22Gu+huiP6qEahEGjPPXJ1sKMogDR1w74Ntcy1RjilTvhAfgh0gej
LNLT2LuvQyxRca+EqMyuXIpCltdK+dtdx0V1iBvx6p2Nhvf+Gwtxand2btx7M1mtmrcMu4HrSgcv
TXsiUAWjKx/O1cRLB+2Hv7CG/gV+AUgNLGhhbiziUIT+aTy251gZT/a8XKwcjZSboM8WNrWekxm6
pgylWyza7erWpqHNJ/GF+oZrcjAonpUBx7IxfZKVyEp2zvW/RhRJeflLwzizA1iUGPYK6VvhK9Eq
BhVxcEfelLB9x4Z6JVa2OCr93jhB3yYG4pj3zRhs3WmzeULWrxZxuCLJ9AiZ6ke12dXe+GWQvlk+
bhnxvBcu2/zQIWyOwdmgyVN9xDvkrGEclKJudoF8tQoKulh61Azl+7oZ+SW+k9xDNG6aLzWsGNSl
fx3QX1tvAdBdhU+htt9H44/+HEo+LSooU14cb9jZWYpFAPUnRns9ThEhAhxVLoeQYjbQTTvd8Etr
b1IIGVfc4hF9gKwE91JXd9tCnhFpDlVYjPJCbWt6kJKCShuFQt2hIeeHVXxRyS3fljkotY50/eAG
Dfe3hZaZkJVZJGZhZ50r8UQ1TKPquIFVQk+x3wfjkPUUPxsOxBfuKUJW+Mc1iE00jrnmgd8HkgZp
KjY0i8QqDkmGcjyEvxpzDgNbU1INT+Ji0Z02JPv1+AJ4u54TT8VPlNMAtN5BMZhnoiHyaeQdZNQA
2TS9eE6HpSQuCAhIP43GmiPvp1Z2gnUgeJUdAdgyaAyRHOktitdgfj0olhA5vQiWWzTfp9KeoZON
CBe5LzJjWcaQtgVKB47+ZT6uUbu9YG0bcVxQzGArbBiehrOzfTvnQVpjDyYoBLcC9yJewR5Nznjg
7cdEMpaFq1SfPtH/v1iFG2Bn41Y3idbvOSAP9GKndw1CR8E2J/wIIF0vr+AciQWrzIhd16e+Ptf5
ED8yZ+fL1lOXM6uSI1dlZAPmECUeGgG1Cu+/jK0lGXSmZBObkC0QpA7IB2CxOwMaqU+PINRc3INU
De7XE5q8roKDSjB2UL3yOWWxfEW7BfXQFGlS2z4wW9w42B6MWUpPuzDpch2JLyomgWVEM7lfW0nd
vSHbKw+96UmcKxjVChiH/LqsuQgX4fTft2HJVsJmaqriDTasDXKiRNuKSNXoTIneYrcn0jrWlgM/
6w3lLmORyIAixxbCukNhY35Ig4Ea6YDOSM9JV8mjzMgBezHVEho7UstEQqVr8331mhIwo4PvAWVH
0TwwK9+SqCZXoPlkkysdVe/G+nIO+yFSvt6Js6X9Y2y4bhWYOjh9Mr4J8WQv2tMB6CS/4q9/4ggY
Gax6OqcDzZufaWVy6tweU4fOU1D4J/hKuL/Ue3iojE3c9auQzTsRUhLEOOu9JIWOrooFmgODW4ax
R4iOWrHl+fRzh2SCGd4GJk9lQBNMnO38PaWqX+g/h6cEZs9veRVCM6J7tJGgP7z7+KZnw3Z1S9HJ
PK5Zi0gPHLrX71QsmQvXt8Qd4EA5WBdy+i9n48Zjw/R9PqZd53lmSytqQ4iec0yc4cqmQ6YYliNb
gO64iQYDBmn57uFSuhTO//1J+iSZC6ydTbM8KCfjM2OHxgRrVO0xKK8rTvegYV3uTDZfMXNFMjzv
cuiB6mEPiNouMypjwn51kUELAaSNNYsURDkt6nSUXyrgnATcBe8NDwaRXtWuKJSY1UriHzx8jjx2
Z7bH1ZwaLHuph22VdYKCu8uncGTEygyziMK2b9fsS/GpsoNxWRMEokPIND+aTmDJQIlKKoslMOqn
J8iU2z/b2b4Jr+/lspD+ONS4CfQ6dUeC+1yce9uAqUDr+B6w/8OKRVoAED0Pv+DVcsX1UDh2dfq4
9L+WxOU51259yqBMKzFtoWDzspsZA69oMXklhaZUyf7aPGOMUHqiP5txjmMoiZINK0vyRIMUpnrh
N2l7GcAjIgW47sTVkRAN26qGqz0iVfCVu4aVUk3jy7G+bTjeC4f4X2qHw6tcf1+LFqJCGtnilTqs
wlJQI5IZF4xVH63r2t1bxzimvAwcwldObriE0eLM8qNOz0fcsP0B1w0+5/le9P3yg+gKvBhERXLh
ccM4+O7pzoHCg9J6upZFWwC7rrNjhjweDxjXCg5fnbMEIA8gdiizRi58WItMt25DKsPZyD4K2PKG
9GtSdnWOUv7jao/5JShgVr0GJZb6JTPFjuCgoTkkwSV5UFbVT+llAeY2Tv4UK0CCSHAFqjzzMsRs
nOR1mY6cmmTdqFoguT/JJSkO5VMDvigXfh66euBDALGNesvRWR7hekJXL0hq8Ya20fbQlwYZC3sr
W8LpQVldBzosRcLXjmQntWpvV4l0ar9CdH/mxja5mTznyKW2kHXGq/jrTktqtabpClgftdqjrFmP
J0yBapOUL1BhBZXqG2KjKs9c+M9KOqP8bQ2BXp6qW0BPkWBfoj2rqTNU5zzX8xENiKu2rTmciDFj
t7L6YITms+rm7Oass8NDCWNwUC9A00ABNsQx5zAGJuE1+GAGGCERJKn3R/izC2lp4NdGGNbCL83u
/+4+3HrlTIUhPHbXHaersPJ/b3jD5g81AQ7SDMTpMhRcwSrFmysE9VhPQ3tnP6Z8Gg7BwMjYeHrC
+sCRONrbP71u/L9Mx4KL5riJ1Y6gM1Q8vYQKIBvV+a3BLe6hxobfHbTnuCy7oE3qlb75QvCcgqyM
Q1C8bwZV/IIKj/mrxPvKsuXNZ/QC1fj6Yp5LdywVnKy3JV4QJx2P+goKZGYFW2i5Jsk4klcUA+WB
acAnMmAz2ENTSROMvZ7YvN36WaikThSExR/rDZtPlPH+rQPg97XMIbUa3w3D6gKZrMQ7yJW07jhW
yPxx6bSKuqR9jAJKo4LP9QTjkcATkavqCrIKBHxQOEMxPLWmVWqY/FK1eATaor5kuARsoNyftXRF
lz8eoqxD9YVVvyPue5gsf/NCOPWfNIMQR145ss9+IApi1CeL5R3cnYuOtaIDZbdYMAcoHAs4k9n6
xqvDzs4IyKvgftG5F1Hcc0Bfuf7NkAIi9o9gFXHDQjEPefmoScZcMl3zAV5X48oemmF/ar+3UDVb
oAvOtVchAfbo2eBWcvnPnAnLvrx7Pi37I5j/JmaGb2HaRLmvwvSrBJSH2h4Mc9gJmWjeljKXOZlX
LZXl8/AAzKOZjM4ygTkbBxZJ2Nfwq4lb8hfbDybZTV8DpsoeS77dBtboqCCsCChGZKOuCMTTQEEx
zAX6oRyTD4C1XjisXtoypwUIu3qmKuwqBdGW8gBXT9Z5vkEyzMECWNPsj3eGR/zNa4ZLD87uELh8
Fe+U7wKlDekFj34GN5zUpRX69kjFlMMX5VKctwXYvl1fo6JRaV6Jhxq8v67lBEGWBfHgHKIAI4wO
XkXRFPm0SIdlRlkDCMZ6TyVzGozMcdZ2kNDyKAXQB84a9YIFD1PTyKSHPJ84z90Q4K5iWkPgjoRS
HLvJMm5jq9oOkZfqIEV/VF6kYreJd0CyjwtB2ZVTwmdAYCPN7CF2i/9fKlbvA/Zw7RlvjGwMA/pt
Jm85Z6wVWn+w6VLO4NqtQUznY6IgRDwLeVwRrdOYX00ntjjDEpdRDLUmfYbj8zMHPMgOA9dnPRNE
eAqB0B8cg4A4GRIWEkRx3kyJGdo0HW4OswvTX/N+E8ivsyA8jf7bZRzRihx73p9MVIdRXznWpH8Y
7Nzm0GFC4RbPLZOuO7UGwfaPiqEuORQMIkrojIAtJmXykLVHm2LShPgqwHo9IHKIF9smFx9jCo3Y
D80ogvsjM/LV+SVNWy4EpoEOaJJih/qKWsCiMqOpSGO2cDeE+qNkb7GG96oIECkaOjbMGMJR+A+G
+s9ElXIWOD/6LeoHVP7LePhJ/u7BNI29HwL8m0BrFHZKRSuCNac4p6f8sofX0TpPkt+D86ULy018
OFAlSUroBy3PiwkPiEy27pDYmRgwNg5wkPv3zvgY1+L4K/A/ezXVh1eEr1SKZcXPADJ0CDL9dAzy
dcBKZXh/b/hCRdNkVg6irJChiJ0b4Vo1pjlcP1FQQ2FY6D1irdju3P91zYsnso2hWwm2aJjmOJws
c5bdcojfLzKX8oyJKVuq6VT9MfVq/oRduWNApCriZ1ibHkYoBtgN954hQam6rdCcyAfkaZnXzVcO
R8MFAshasHsoZAbh340VnBeDS0NlI5y8qak3mOn+wGr/0rtN23yCfoqwa0Q+9U2knOa8n/EN9VsD
ppkEfruVftRH5/HbTXNCA+5pUtsU3hpX7BfnuIh+J4tXUia1yhA47JSpwJytzFZ6bL7HLOib+iAy
GfpogSzOG+3hMi2OIzLpBtX55+kjEMCrMz9TMspKDQp4HXhxwuVUBaEEpcBFkem4kxvoE2mizGuq
gseQ35imtglwEcqBYlD5rUl2CR1Ir1iS90YX0bbF2t1M0T5SNJ1kXZT1VDt1iZb+1GU4PMB3SpYv
ysaWxOhUm7T3i77gLfqR3e6p9K4nR5r2REiPYM1zyiAMUzG+ktej5AGfXC/mk7x2V5gUC3asF+0K
8HFBHjezxaUXHk5JFa3JljrmX2H6wEl+DmwNhyltY7BDb5fpReFM5tkt/f/59n3a7At5bNSuUz+k
GBctJO7oWwV5sIOXR+1Dryl0L5m9tx7NkPrGkzlCQ65NhYJpxHAGZEnPtGBDw2UScWPXaTdll66f
WTzrifBu29tqExyUtrw+ZWK9JPWcHfDu7wIk7j1OhYz5FHwUFX9ShbjzzRrmYxdMM7YH6d7Te4gd
vjAAqHxL+hf+2R6ZWsfGIKmIEpTmj8Ngo83JadrdIkoL/Pt41/hh2jqxh4M/WrsH3WQYnhjaNkql
uQbKeLbgJKHB7N/UIiqT/UTnIbhe8TfZIHsc/5U6lQHkXmkWqGUy82P+hGwtfQ2C6752rEF5rPrt
TJZUwo9PDXMkCCb/6gkdIP++mjGMqJqw2ZZfjVXjlauqasebf+BQo6Ytn40QBK0yHyNcDTr0jcxu
yzlLraXh0aUDo+U3jF8VuY8sQoZxOx5UTxUJi1TyzLjqdegHn9fS6sUyA1dA0g9fO8K6Z2qX3cYi
irukWOrwFtL5zDvWzGKCYJxLEVVzsSI4tkcjGj5KoKrdq6Unff5YbsDpIh1z1bUC/UXEvApCY3J+
/j9kGvGHOJ6/4kijHt3tHUjXqhuM5EoOWO16j6AEXiTwZ51pUj1PnILaGWNZg4BKlWvGpwVhHDjj
Nq8uM+ukCr8Df5HxKk50C3Lm/7GFXoK2Mp7kFdVybenzDELaYuGYmLNm1NHvSCP7LLJY9nRfWegc
LSoPrDQowQGUmMpxSC0WcgkdWTDtG+SDQJz3KKbbaUjbZP023VjOq4fuW8O7+qv69eN0MGM4xlqA
reX+pYgn5s1DrKGobhdbuJ4ifyID8fjXhlGMwyAXARLVjC1WhUaP+zGgzjfs5Zy5Dc3kByW6Q+aq
vZGjCWHf3z8qJpATPQ8ej7TikKBZccjg+VHr5jPFraR0ugQVu/jhK9nWCLcsd8I0k5IS/YmrQcWC
zmLT7HhXnomQJLlXP+tF5087oJp01Y6FQKvLAfZbJSsudsWH+C3cJzlKSjehNJsBY73G9Oka5pPO
avflDbjfneVxrFhDZ1IzC7jvLOI1yM1o7xovGNZcA1Q788TKZJk/Sr84RNHRKZBkWnTDmdn8DwLY
WdnqJTJhFwr8D3mVDcRtVdlUiWK/loHkcrneYONdidKR2GG3U1jByyU+8pbBNIh338q5MLG8g7Fv
AO4umGMBeInW7PhR07VRD6HCn7Hef0uFrwm4jmlV+UMDRIZC9yorl0eQNydo7lP+2WZoH35C7GEw
Nqa7mYa4QH/oE+qPGzIvo1veXCtm5lYDRbbGVyZVNqLj/1RZIoYUxKKzt7dpJbn11Nbq0qLUktcq
0QYstRpThQVPvG+/qs/EkevpeBnedr/wU0D0baEXrroN8CIrclVQyE7EjbBptbYCrQt2JhAYyw0F
0nMxYmHhmOG2llUDLGQOTwe/7RAweoy1vrcKgPpx2FLBMZmBmqwM/e6pbToHTlphwL4dzDi/hMA2
EREgbFB+aH6rLmOlNDROBN3IHF0ZjJg5oLcDAZ8PcLGJ59lVBpbEp9fR4OgmPgPWaaSrNqfOV5Cs
Cok5jEaHWD+mVtHc+h1ECn3lzzKIbQ2CsoFC1Juji0d+72fhrC1Y6vdH17IrkT2QNAgCckatwWWM
cCPq+npztxhzSaYGhqBRW8KZm+uZLrbIe7mXC783rqmBA0iHOhnLEkHKIVecj5lq4qlW1QBJxi+y
ataOhHlLxfkAjV889970k8qqYLuaEguKxtKHy4c8V5kFYLFZ7pG+6e2hKHuKPxh2k0RP8kZ4Sqia
U0Ud47EDD3eimyYi4GMfH0JpgwZr/RZ/22Knvbvn1W/Y2hKCUwGkoZGfOb9rXBmzpY95HrilS92q
W7F0/MzF+XnIGufWFdbBSU1oqzN9py5HYL0A1MIzK5v8PWVAFh7A9P5D4htLge/nZke9BG0JKEhv
UaILtD9W99BTTjkin37q5d8VFRAwMjh2K4OlCP91XwJAXoYuSwWpuLuZ7YrBClRK08/NjM+FL8DF
gXgUAnq/hE3bn68fykKwV77mPh7u6iIPKS0yaJQy2FSfpWWoq6pXxR4GtrAhmoYNrQQDyn9jbkwl
NkhxWHIFbTbhGJeYORJIa7nadBc6J0uNNNtTIh8cpFUsib1d5MGGWR8HroWWg9d1b/ISQtk/4O1P
k5IIgpUluQ5HMYePIvyiIjgRs9t9pNxMuIPutvzI9Yd+FO/0wTk6gY4tioEdjcIplp2rqoeSJt+D
1bc+OAg44Jp8shIbFMw8VFnAAYevZDEsTfuDpJ+ZrjUeg4IlmDfGxb0JawPqwSE7/bE5nnXwxQcx
2P6dReuU2pSxexRe+cRjHMNxmB/sF0583Wg7Zr2rYVZf6T3Q+z0lMTD9P3ycE1BfkR8pJw6hl7EZ
dVdCIV7eZsao/c2huGXVeJdLVT/y+QEErSxFX4y77EHz1Qi68Z4wrfbYfwneoYPhM4kBQuOZFjNs
gG79uDskpJzAnQ1Hqh9OZolOFWWB+BsTpl1A2vcCwz+2v75+lMiMHgDu8uIMu56JX4n9GS6N5TDh
jkRQxoJ3pzHL5s2S438EmxJDbxWZOG7buee+PKEioJ6DXoJwDksZWPu4wBfmxtI5MB6HI3aklVlx
VZtnk2BRYMZiXAJGZONOH3hqOswUbsyPrwtKD9IdU9o7FFHfU/Z7QgC7MGSkjXuLr7jR8Q7DF2ik
tvw7AL0D7zROzxjpLgC6JgBZ6hPCjAaiu0XnnMa39iI70UN/hxWzheuwBaFx+CssbfBKWNuIa4DH
RsSWS7fGgOXEgM3jzEj+g/SErbNw2SvnvVDwZofKC3vsdMl/sgAeCnLvWvck0iMt6pn3XzHQwS1M
HLsWca9q2J4Bu8CbZfbtJyfcmJPNML67+IqpOBmScF7MwYWyY0SCYvxW7yxGkZ3j3p/6NbNyLyYR
+W0t5+nc+gDDgi4Z7DskXwqPKO/N0XTn+v9DIqbyIzXXTbfrFZtMvEqBMPfdZd/fVD4qDlJgYDNJ
FX593u5VNjdJQrxeQJllBlm788eAHFKf8XweHgDtgoSFDVPVm61Vmo47KxmpO1YONoAKGGrIel37
uZfa5mN1MxWgfho48rrI7jRPIZq6l/opK/uzVW5rXWPvBnbbX8h60ZZel6XCj1/BPCpKvnkhAwz+
wqVZME/qikPo4tIibBA2u7Zr7XBvhaJ48IZKpVv9UVafYNgikPqgyYENhrXJSIhNZNwW/d7kF3JJ
yKX++QplxZZ3+B3DVxlEIcYs0L+tBF3FmF9sgJrg3vfExjIBxXZdw94T4eQz1y+ylyhkwin76MI0
V0ud3ItPbmJ+0cFDQD0FnwXZj4OgWBwAtn85bvdAIdqwguQbrvnhTZlpbzBn08Hne47ZMm7XWU6V
NOxB45Px01ufohLvPqoxtzWu6qUm7iTPOqIF6axWFgv0w39ET3JalGpAOECkj6SNpM+bb2+IkANR
SOhLeGsGVwGayISjINKmXfoPd8hRU45joIU1mZJjH/OnQf/5IHFdkUpeKz8k8+2l5f0knYfowpt6
jxUhPI099hFGrArgousOSRZ0Km1KadvSG+WGAOttZECgM7nXB44EsPdzGsLau++BKtPxasb6Dm7e
7wzxokF9/Z7XuedGbDENj8iFejFUnUpL5rRx6swudpmkOlV97RRwWuFu8snAH+h3bwMBTNbFi2QJ
pNA1EkIn0E3x6IOuz8AunMrQehgjpWc6IIbEFCWers/HGm02er17u3vvGLSJIVYn2JubT2+YPRtx
XSHMkdH5QFTRp+DkQMvg9JTmkDQjtNEbb9Vd/lA5TPFLQbp0Xp1k9OU5rohTouqabI3Xt7d9vgir
dpLyyeDrBA/tStG7jV/84d/oHokaaJOlLU4iAebyCl1Pu0wrrAsUf2hszwDRzYx0Ve+N1CEYfFMA
4dzJ634hsqS1oct0b6UpdTH5/mYMvK4F+QkLdxqHbiInrZNjCUT6Mege3eKDvZBa1miS7Y32Cdu9
O8vWstlbF5W5uoRJdcwBqPC7AT+C3kCLj1xJ8m4ufsPm1r5WUfq3opogxrBtsq8FdB5zC1JuAQTq
AzSVwSC/3wXaNa0WOmbRwNmF6q+fma10UcOYuswwhJijNXR5Qu6hR44TJ/aph+Eet8uODou3S8m5
i7OZ7HyCbgkjP5Z6X5F7PYe+iiBDZJ96kRdRygMSEUEbhwGXs6uTFHzfl4fBBnXLwOjY/Ug8K6so
sZmcEkFdCmrHhS4Eu0u2U4+Tq6bt7sEN11w/7hVWb+hwgtf8NIqztEKbFOrjKNmW+3+jfS0sbDXd
S47pllmIXxNIaCWlJTWs6FsZabtLIGGIRbaApgw/P5wBtGqYW4TN08lrRnxl4odku02wfDiCz8D8
UrdwLT5Sc4rx7fLrAr+NlytmrY6NBGiQWQsKKOG12KoczfJmcgp0JPtSkPxm63pDRdug6Mn3z3JK
F8PGsipWgBzAjLZ4uXIYCaxlzGYEonmMulNIoNCcpOnM2/GuC/gZ8RFoMusebfNBYewJJP1KlYR9
7p4xaAi6yx9dImSf4xPJj2FmcVjNP430P6npSZVnWX5KlRsIatbWnu+ykbafk44AQSYT3EUjNQe8
XqxQ+IBJ0e8unVL+OSP0mn4heHBFZmMo8YEHSAT1L2oAxs214/Oy12TYjQsm4w+zEk1ipq7SkSUi
04ou605dHH1GEexdM+vNqj7YK+XJVjTMtkkSN8SorZytsYz7uWmmhB9KO9uePi7Q2jpmpmKcwEW0
PuuqVQ6MqMebBvSpUJt3AJLMJBXFGUt5vTmcaV6G/o4oA0xppOUqsR5q+rOlCLh6l7D93ivU7A/l
QalMOmm96ztWWsFc1G6ijLsVpqWizIfKklW3z3bTprIOOpzoY5qqMbg7ISUg98Voj5Z9yErPSJ6P
ZYebJ+QKAgC9Whsl7fpZcOmcxX+e6AUmJKAAYK1uQULvy/M+AtHEvva5Rz+pYzbr8ZjVkL+yj68e
o0D+HJd5lcUK+axvtjipR5H6kulvZIXBVjccXsdC9357yOOrcQbs4XdM1M1/+srYXXnZS6XlDK1g
8T7L9wCipFzL0tDVNaFxHZ3/hqO5b4XvU3qLAnE+mCnuGz4IhdW1cEUkUihypkbsK4rW2ucJlmPR
SKaRKdzY0iMda6J+0nYBA9NDKauottvxyb9NPQ7MUOQhA1BEnFPulYnuD8c2gVwdEjIFUF5+htbg
/NELLIhiC2cBrJkROaiFi+JvTFPlJVCKpuVvCxbyr34Tjp0Ko4+PIwIxDstuUUfmQ4vTOPs2e2cB
c7LijeNlAtRY2eGzDX9YS7gcqjcRgiZ4eWaA75L5au0Rgq4OJA3dttZKySDQnq9Y9DL2OUB1CQIw
8nw2ZVtSbEsoVBIbjPKcMyoKlC5RcNDmMaczM+cdy8q5E6eSYx1vasLrMfCpTkLFWdyAR04+X1Ka
BQIuaFcsNuVZOyFrROdmKThA0eKqH0oRXSa9f6n0BEYSrgtUIsqllodDTabHJIElAYhFBX6pWCvY
Ac7MJV34i4+jn5ldnTZq+Pq/fftQ5iXQcDcz469zviqpgcV3BbrRVfvC51arxJaQCeJ9FoEFBtRd
iotz1kvMzgWWX3oUteIHffz4Tg8aoaIOWzhXtWxcFX6cdg6iVUufWp6QsDcbmfWzBAzR7gtaXReB
R2LoyPdxPP9bezJkq0CjX/pkx65AQqJrY5eStA7QJC2fz/i/NxqGvYIUB8NqwulwTM86O4lMVo9G
Q9OkShGQmMYYHraE8VX0B1SEI40Qp5TYlgTRF9pCnV+xx6dCMUuDrnoMAKkTihCvML8OhzQTzURU
Ka5mjB00kspLjSoKZ1pWx1thz4PNEV3MhJFHR1dKn583g6tRLOBNubdFAc+jV9qZ+a8SF8lOhlE/
3VARFflSfbH0zTjQ2BsKDpYk+Cjkbr+rK1aMKQ+tRxnzESA1aENyURSDgIu2p+Voc3LmOhFy4+OZ
B93kfXrRQ5M72jkfd4PjQsGzKMFRZb/3q+Qg25ZK4RKweAylK3yJRkEHtuzyukdu6UI6d1ZLGuXc
//CBCQRYtZin1oE6JJoKykRqRV5QeDkrK7pTXhBTcQcu6a3y5OSBZd+uxAEi3O2C9WgQ1Uhe2FpN
KIm/jCtvqRQQz9efGcpyC2cdXuIZu+t2NP5Z6Gwa/lA+Lfyg6YYx0SI+nArzX39z3LhWQpTMTCLv
qyLHYCEEIT7iQ+1wiW5CGmbStu2/BhFKodas9x8Sk4GqiZvl6lGmPr/uGeDV7uo4uWnQVTq0jr3h
IlxohOab63n5P8bk4iSke8Bw7uY5CELEVNf4dltgOO7wClqJlNFADqssBpq+VJRljONmZ1031S6t
uCzgMyhy+2yIg6C4QyxoxpGg0yVPj7Tq9wwqIbOqL9vQ9Nha6sTM/RLg4fIY8GLeev9qANRUlsm5
vm1xF8H79NrW0tINMmmP4Poj8nA1dTMm+Ydk9i4qWCpVVCltBbA6HsxsGPNYYLmq1XzqEFKOH1mG
yYLK2KJTonEYqZpbZynWsFjVktA/095zIOhKj2MfsfkKH+6RIBJa0PLsScdYHVVL7r6iEiD2WNcB
5P1kFw/WeCgjluXZaqtBVPZ016t+AmsmgY6HElGdmhEq01V0eKQlC4doJJy+qRHmuOSZFlPj/vCC
j9vdWoMGf8J1gOJiq3bLqYkY8WI2kQzrw3HbG9VhHtr/o0M/xHkUg3PF31kZ4fBmqd7HeSbVKlPm
IbTJjnSqTwlvoVyTYp56OZkjhVhz09d1KXhtWpYjSD/zsCLGjBptXo3t+W7PNK74Hk6gilTgyvpX
RAI0QZTeuIydWp7lllkQttTuIyJnVTypqGSRsqQZ1q0gHQ23OVf5oUQ6eqfE/ZVe7z+yScH13WiS
qPjJ5FvUifDF2FPVryo3uZb6xZ2h+iNXoDja/F5kmzBeaEKPiizk9i1FjLTDrx8XM7zuhN6WvQQl
Xp/CJ3DCHYl51UpGPWurqjovoupq7aLKyThHI+oqWd87jaQwXbfuyeNDq+U8tEWDNK+CBSzf7iSF
Ppb+PV9oTq60nvtsFkQ2wHcuCIK3l+osQpbCUftm3rnKIRgqoK7rH7pJZU0i/mywTZ7dBJ0P0Ln5
ZPOYymE+Pg+boLCtR9OLcENemRUwz1dx9VLH1sIfy4PFQcc/DP+WbPpLKfy7eiVuxGjZL2rGHi9Y
uBYgaEbKUuW3zKIRrBw6fsT9M8cWWwJhvMDhjqvWm+QsVKIvDFqXUdNBTJ566TKE1kAwFZa9PeAQ
+BjhYvlL30cRrK8zUbx5GfaVHR+oDyKqVmEKhbd47ogdtqSP5Bxc2SsVZM2Un7PYuYWr4Pi845yE
9ehjG1+rXv3EPVVU7qnZ6JED9QLgcqRsRPWXr4enn1s0/6g06oRJCNAeKyEzmn+FhaeyYlG/j81Z
ssgXSYMENWjdUoxdqFnD2t00Y1RUcUzCsMSuE0hMbTG+velrwqjrZoWNxCUPDTBxZ1tuBtzQoIGP
YGhONkGikyhbPhk9L7CWCCCevRvI/ItHBt06LxBZ39XWrjCR+pARkL9N5w04TYKzeLl+1E8LbFFz
TwD87uiIU31jAerQMg4lboEZXx5m5tNy2EQ9Z+5J3eP5SvpMZUkp6+mH3IBUTCnxwmoPVOos00IW
eNyx2f0RsQmV2YXhFpbidm+adFzC+MIKGw5lejMDV02ZXBVTB9iTfgYC8fRSJykmnPWjyb9LZYPz
krfJMPc5OoyEZJgQHlMFKhnRVNMC9tCY2mZknhXP2LzPCEYynfofHIh3HVPXoOYJYfXWZfhS0+AV
F22nP5q1NxasM79WoTViACHuPJmggBIcRDZs69MBxy6NvbTsVnpxwfJvCJ1SGwGJjKMAv9E6034K
ekSpEhnzfidVL/67TZMdA2Cvnoi9KWcvvpQZCJpGGbai/sgcOpImtlurBIXuNnS/9jZjLHXY/D7m
SW+M8/2unPtj43A9Gna3jSI+CR2t5Kypd7DsQukTTGvDqt+sBrxpzI4EUQ7R9xPKDikkFMsRmjmb
6uH4SfShrs859YbL3Qr/F/SA99ktNUvJZBiYlFNziLSZ55hc37UDtkIpWUG/9RF7OZrOsQxVNNtY
RrNhysY9qK+yK/2/H5bQ41eDiURYvlz4LQgdN5pJJiScvzL7sicde1CYuIh7FEmmvuedDe/qizM7
Z8vMFoRKYrv+DEIU1NaNHn2XT1iErVqi3OnlZJLmOFA2qz6HGeIUZHXJ1EJsYYiE0L58ur6IDjE9
nBFmaVt8SNu9MwMABGHX4Amo0phDaBToxRp/4AMoYBUPVRZuVEYbRwj7FVNB6YfUcHy5IYJ16Odi
zsqNmSqodij7K9WKbODlgY3HFQGKBIFB0YLssbWr6FhG3IEVPAGDookDAiO/fWx/+uLqTaUsFrk8
Twzw3HY78bf7aKGyBijwsW0zxqIsYBzMVrQ/zB9lrFQu+WljuRLXT3v4uomq51UlNPMZUIgG8uGR
sKPuojwRVcyetDlNxvFufmQCp2L7IwsTZisWxmOU4o5eHDzBEMOHmxX5US30EH5YemgAJqO+eBOF
pKKi0jZ54vsG41mIgwxgWtbskp/ga/saPlEcXwsGjZ/Fno+hk8sTiXYNONpVel8s94spQ0HqFu5v
MKSwm64I22TxFgw92UtSHYN1OViXiZVYOyhu7H4hY7kWvL1pHKb43YqwI67lfTpXRVA/t2Jb3T6K
rddZDaSav2WYe41mltmglcHByniCYCZzCuJ/BPG1dBrhSddNxh294YPxG6eTAB6zBVkPbIaxE9eE
/3jaJ0zs3PI11hTUU0dbjssRQRFGDZr+cyrxnJBn57yHA6FmmqrqqyVNvDtp+79lYUg9rZXaLTl5
hl5VN/lmOTKKRV81ZovmVvuSxjoyGs6FlPk55EwetQCAmacbza+YzKbzdbpQCShA+gKOhzk7J7Na
zthwTQ5P/1nbdKTrS2HLz9vyOBiLsVAXqzEWVugwbrQZRjLmoalWnoCSYF51Yxb1rhXl5CbxWOar
Qu4mG7h/sIxKlxyowvpUD4e6ipVJUZ7waRpgHUUjWgPNQlepvDK8vq+KkbNrFTxxsXQEX3X5DGYq
HCmqC/xi7n7qCW3RgZdi/KLOCIpIV5iHKR+7kg3vOy+xwRXuuKy4u7nxVwqVR7zqW+mc2THYwLnS
ypHnByrO1BKXPGKNV64NXOUnl5hzQXVqgy2RoHIgDWk91zmkaChWlGnFHZe6lMMSqWD0yQxn6Ks6
hDqFTRBSFchXbPtB+g/RIsybXN9YJTOukOeSWlDEfI1NHznqeWN1sybIsOHs3Sa61txPVckrGcxX
ptzolmpNZFYmkF/zPoOeiKTqFk977xb35Jyj5dbsZe+2EiqbEJJzrVs0mOtwqhaPHK8/VAAIwjXW
gQJsl/p+x1CWP+QDxxzcD4HphqnQKPrr0S5TBBUSQ1kDOplT7WeIuX0+m9Gu7KBW75SwT0TO0kD5
Khm2Ggvq4asVDaUYcTILbfVDW8R6naJZ9j0P9ZW3njs/O6W7H5Vxwsd6R6GbQaX8vsK5ujQRkLBY
snlXqYw3i+BY1hDJFv1cDutuqcMvGGq3zOLoLGnCI2vScs+JGQiyoRk6lJHLYarJy14NK4PLpDpb
tOreHNKHNggjxPJpp4z23cfVYQmgU1WKOqZKlHmq1oTya+klyJftyRJF/LP3VV8A4ifQF1DWc0EI
qQbtznVl3InftC2wA6i4w/KZZFk/XduzlY5qU38mn3Qsm8UUg48RL/ZM6gTyv+xq+BCGMWC3GenE
aKrr1JrTO8+8gC+bjgLixvYppXbhi9vf4w1bzwQ8DaeglSIozSfWrB9e80cnMGafRaMTygQwjqpT
uVl1YRF8cGN6WF0lXe8xX0HOFHB85liYBYceoywBL8hs6p8kTC1LXWRRlosFBvrjnp9JrC//Oqny
1mRSjKV8Jzgq/XcnHGUV8d0ej2Ztt308/CcxAzbz7Bt2ruWZVisviMXrMpyyaVHGprZtv+TQ1RY2
ZEZ122TDCnAec20fP+NQGxsXykaGp7TWcyhgeNG+ArJsmgIMbFJ7nHonCydjVCYPVPU56az/gYsk
J5RXEmnz5q5wNLgcmWx+2jRwREaAAaNARznOuMGXGIBSyv3KNMfw6GLJHeHNF5wY5PsbU06faSfr
Je6RBQBmjQZQgWJHzliVZM9qj8IFl6tJb2VP3eUUIFk62vmviyrLTSE4lpRhQ+qzNXKDfW+z5ILg
Fb54uZbOg7//DhIK9sR6WVjwoq9iHdZemglzdmlLVDy99YUGVvphYiJ6+vmHH9WI7PB2TSKToPGI
pNdSodtusHzqjIUtYde8CNl1W8FO34v3+3FD7PDXT/AUENStchEgOHYAXZrY4skspAWw2AIvqOk/
2TjwANjx6pzBT2dhDW36tTUwKod/LK+GTL5A7rCJfvvG93X3Hop/GXacV3o9QWwDJLTmsqUDM6iM
64exFIVBq4IqjCjWU+KW/BGRufWfyt5isMYATh6j+320zn33LBXV3JdHmVbSxGZKP7aVApEM8bzr
fc14ECJ2FuEuHRcwGiYdqkaFhagcbVDH5InKRVt1rbA7dqR1fAeW7Dkfb/v/JCsEmZH8B/ewFu2l
Tav/0LkUKseg5gaqtXwbzgW9NX0feQPHjvbjeS8a0KmALqkTrNrtfnCCAqf6jkU/jr5QhU5O38KK
L+HQOY0gc5twM3HxBOkVtXTkMmQDCqSztcQXJt2f92G8kDbEwgZmVVAABo+3u4IkX/49nNt+wtHR
6DNh4pRuHkM8a/Lv0/V+1O5/RTOWD28ckNZXTCsaLf/hDEuzZome8IUOy6aWHD+Y64WwLMcaLjNP
4bEyNek5wY5DMpq35hjaOq01htsS1OXjuOpinYF+Io01KRodNAjUCcX+Muy+klyL/CG519Qn8qhW
o5DkmVZeoPopqoVaCluwlEJ6zw9SHtah2PhaSNBOOVd5k7oqsId//i89+huVWaPAWxqpjVWs6sBH
VKcLzxF9F8KW9kKfzpXKhjPxmQAnKRdQHHapjVEgsbTSxGx6+w/gHaquzM2SdYciMkWkeib1T/Vq
dLdCiZEkruB5CpPYmHi6KyCETN0Q9c/GBxvPZgLraGVFOq9VbGPxBAN25xEqjtGWoxldFavc1u6P
SUw1rL7nY57CGq7D3M1/um+oRdxs/witYIZ7WBZhsOi3i+TlcFGWJIidCkuj3aBE6ofK8RZa1Xn+
cPat7uXyABIJVUN7iqWPaYI2usoyvHIz35XZ1qmxKEl0un0Yuk0BXeJ/ZsJjk2I4pFv++WP/5Elt
11Ee8iCVRSXDRPqXKFJxKYkN2m9fNmUshvwWeJ0Bzu+JkkFJ2XGK19U4z42NJ5P1FHeQdFfgwoNZ
Kt8XcTLsfL6jft5gsknADc/C2uMykw+BaCtt4L8Sm+5HReCMAYr/ZZDtFH3zWfzewQCwU2CfaKHa
uxui1OqFk2vVaBbxOyqXlM7dcMVS1POCRk7halVmaWel6H6+vAZenHqLC9VVS78HIkYV2E3auD5m
k69GFf2GjlVH0iGxaKIte0vFBouSeXV3GxPGIBRBMKv1lSlYhkeJTRMt+96bptY8JAhnudIr0XIe
2WpZwz5jvEaCKOVr4xtqiOG1YtHN1O5zHYiZUiE3r1vlOWxpEZ3kU/XnQyPahiP0JcYs1DpA3P5l
ttp0xvkvXbSMBOKvXj8Uk4oAxoBezW/UXvtKpdQ4o096ratfRzup1S/acxjRDkKTpHqAbAl+y8BO
p1VWwNWUu1mQ4pqrjBQo66tlKd3l3CWt2Nap4RvWGzDOeMaIUmUujYIrUix4MYrBRawohgZbOGV2
RvGUBVeMilvCmmqv0oHCw2sUyi9Yrq6JBMJlQpwIdE/UYOzSVA6Oj2nh7o5FI3uRbEfnPSBmOg8B
l6sP8Jrpfq0Cpu0sauIoQaLIvZu41/lpr92Fj/g6RfemZjFHR0DXIprG/3opnN9bb1iwoHz2tGhn
rbHVHmQx2RBPq9SuVSN8OCbEzx98GYIMVh5UK4tTvdQXqG/GZwhAnvrj43HcBFvSp9RdVzhiHpHf
yOJVaBw8zP9yd/WszfTixmFGJOzorVGUZlGRpvMbf6lh8klAa07lxYSRIrXvlH7WkY49oaQzBSi7
6hHu+fh8FfXJoDUrKo2CPufjVCsznfwFYHvegAb0jFUzoHs1Xg8XujB6XxlRkELWpBMwUnux1bdE
KBffgLksvAuurILWb1MYO2nH/uWTyZVkZXMNfP3peA4nInF2NzblodlI6gxqAtYgLoAE4H7b4L4a
QMzzEukt5EOOwmlcIoB+TamPesndxnn7OvuyTN+99i2r+ZFMTQ0AUkZ7SM24N8AvRAQv0Aqd1efi
lmr6BSO5Iw65XHrdV232rzAejYyb116r/0bXlpZtew7BTGqURdjttIxSxigDicNmiBoiNVvrdiHE
ufZcmOJcgmeo9ANFHnjzE8DD7YoHDEKnTptC7kqkduPhzDwar7ZkQbvSY5tChVqd8Q8sQPGtPL0Y
meAsimWpumiSUQBJkwsMYoMfSaazFORlhQTPMBOm6xnIQtMIskpl8IJype5B8gunBlhix4dgjrKf
5dFJDoavMQ6q6o69cJYaCY7PsRVHOvp4pPwetbnHngsvaQ1NDODVrTFRCrEHcosdWbOHeGVudgHl
AAHBrzDGtrHmMZW4HlrUe+5lP8P7uPT0RsMXroomJFyj3edG0DjNo60R/dslmHEeUO0+AEJWINP8
xZzcz6XRWq3Bxt3L/ppnPZ4+r8/wN3meqFqfu/J1AqO/d4O42ym8mhpDNTAuBwYgq/CFbY/h7iBe
qv3wvcpSmK1oj1XQiZchqVK81IVYM87TI2YBQMcJ0qvy8b4CVB2tE9Oq1bhEyPqigjtFGSVoJ8ip
MXyT3+NGRJqgdWB5vSIr5OrEY0FZbdlwDQOQeq09aix9gXpwfbnzg5j9CR2xtADXEFwlUchb2dVs
0p3hVCYzBwiohUCpvybXvc6CisYV05XQgWSbQXDNvfXOBSLLYynrRnCzF9zBrFbMGPMA5cFx6VVB
OVPLAY9WCjz/bwAtBksGWSOZBTEj1Y53ijR/WSuw8zKiBMMl8I+J7fLvAnLMwl9GrM8KMpBcBZ67
UpNg94mdzba9u3x8k865mV6yT2HmsCPr70CiROUpxHunYk+KHfOCSnCbQIj+88iPPazXEHCLVnIW
LGw89epa1+hYayrGq9vy9GQJQJaYgwlyTdze+K6mi7fLFs817jWV1lg2qRO8to8xOihlMF/IkH27
bYA6LHjtgHaScEIFNOMClGmiyB0BDdh1bDDJqdP7Tc/fGYTGx9EhAhXbYm6xLdncG1ruzmTNWV7M
IWcrHZK/oCbSIpZqgS325v7PIFKnP6z6/FenxCAhQ12pAjHp6Mo9SbNNLW/P9YVaAxOWtLxTFFBM
kMarM53hHLGpigOEYXTj7FnyP0R8FrO70d9MXIUyMXEV6YvIAmhyM8hOhqOefB+gfXgjb5ACE02W
XQmqkDIvAPkruuoI4ZVBt/bLVxwsFBFsJ5QlxG63hTkI3Ds6Jpiag2cWPiAxNMMqhZHBhlhLcxKh
MWcADjUlehaq27YM7CHaVTF04WpI4uVRLmmMccSbsEKI7C1CiBaEfgx8KvN5YSUk6oUGEeimHPhQ
Isz7WOg3OBdoIX7XvQyK8TqjyQfPk30LKAbXl8manfqdTQ0h+XeSLQf9DxZ07cVBa5cwptd2Mknn
atH8bm4DeCjHV7XKIkeU3mQ8mJwq1Kxq7TIOxOaEXLbAbCzvGI2WiJKbOA9USFRTvmOG/Pfw1Cvm
zo/zNHK3WP+GRj4rMJ0ysQn0LuhfCFGwXG132K094Uy7kwK1Fh+Vozgmg6YjvmIl+i7p/TMXYPhL
6Ka98jg2c4iAAtXVM4IXqN3oIoIur/8+hIVABBvAUwvx4hReuanq9+FNdOkNsOwmapRUKjht9W7f
Y/XtSitDaCS02FLPsIpovC8+J/w8UOqK+zj1iSubvA6DzSwRbwSc1IIC4+rlTZKVF+/HvfgksNWv
w14bcBq+o3N3LAiNII/4g7LE4O2u42twUfnRU6QflNcyukCFhisLKXZPbYHvL/4bDU6HmaAV45Kt
M8u5ErA44Uc/tiD0mO3ktGv5yKXmB1AwyYEou0zsgS66+4lsbA6zT77oc4Nzlu4JWY8q3DOWSOmn
p/kNq/wenAJzJCtiBhrqDhODKpm1eF9nb6WnsmTxpNT+g4XQs5S/EZbxAfUESym6U8Jmz/vc7Dny
aH6C3sjE2EMDfQxRAgngWGYAHVqydWaNFJeXSKIq4lNkYCFofa5rB1jAObS2vpSOpstGW4f81rkr
kVZgkTkAWsPXHGdAfm5qBz0CwdkNOrbAel6ePAwBuOHa1m3VU9eVXuLzmZiDGO1xr3PFpk5pcv5B
qRGqSJ096WOKSK1+t2zTG6x8/uBWDmF9Ucd+j282vhuIt85yKHR8nytfvtBreSeos2O19ykkRjq8
KG63fV981u3A8NeLKexMFgYORaAeOndU4KaqxOqn9gSSJ7khVwBKDfFVjehiN0UgyP8fWeOi5VeC
i2Qy8zzPBfgFcIC2yDGwth8SuAwqpuptS0n4tASOaHLq+xCAa7+CENShhJ/K/AGsSKB2Tcj/jeK7
FhVDBunzw+GYy+3/pYP1F6zDDmIsX2/o47N/G76gBTgOWrrCCd5dS1jpGS9M9XNeSiD9MHOxATHl
XYwLPkffkI/FdtgDvb5yEjyi+XInT/DRK5w6tIlnqB70DMomBsCO3zvtIgZ5Bg7sOAf/NRBMY5VK
+fwO7NbbG4Emo6/74S2NSOcQpuN+IpohVa6UpWj9dKsjrT4XAzjHWR4JiyAtfoHoj0KJCeSYNRhS
qxyPzvCTpNR02Bha0TX+bTYwisSrMOgWVCLSmW/4HwdNJK3O5ZKItRnm2p1BNHFR0m/cFTin6/HZ
z3XnkQlB4rmHeWcbF9BtnUC0tQ2za/0SwAVX8bAci/+6c+ReRLAiWJicp0Y/ounGRF2IU5/nKfJ1
WsGgMejuYaKz6lqaOuskll3EfxVPePXtX3iCYW+YBQN0o/Yw90odK0hSURaSBjkuInJOfGetF4y0
OUyYPNaA+grszC4ZItyISG5SuNSDrGFStDDxiYP/OADVHpe3Pat4KVGf0w0PgSTfRtUeD5BZcHLm
if+jCClvqtwzf1/kRGhEiZWAlMqTgdr7Yqg1HxfzsJOmz4VbjRCk9XU1A+EoACJj2k/rN3r0MOIp
Az5CoxjkEwxmbzZx0Prin4ovBQb8OuhAoVKMMm6hUIbXZPq4RFlh2ayqmgQ4r/+yiBiQoCSPfn6d
qlqYbN4Lapw0M5Nm4UnbI0kkJqM7OK1XFX6irwLBxlo2cqpNxTeK+teHb3JvpLdJRlGkUK2KvNL9
IPckzZO5GgHobd+8i7CM4yZupTGz0jkh4n3pd2P24Adwt+Gud5DZhwsJHhVq1jPFH6mtzWOr1x0t
3/V3HpproO5fpEPD3Ab2FM8pqW/irKAOakmEDtvXezXKiFhFfqhqW5LFRUVVD2iWyzsiyhLkP2PG
NcJWj/wPWeswIKNc9lC/ET8u/+t+9W78rBrBZhMzGLJFdKSd55ua18SL3bQ8Xifvod+he3hN0Hsy
Nas2AePP9dENJ4ZUa7UNnHiE/dlP1u0tCDHmz+gu8WaRc35jNWu4fxBGufFxKd6YnIVn8xeyQC2E
lVyhVx661QRPx5/JOWaUKvNHr3P92ySAiuL1bJnoHrtokHfsHIst6j90ppxfzgYs1TDayOOpsyxH
boaFZAua3G/X7ogcsIjtljvVmPPePxg/p6aS8k7UI7KXFiMn1JNe3hT0c+ZbpBxwraGrKjq1z/cE
efTy7TCOo0GHDen950its5PUV0OdmFKc9PB/U0obJAOtsCjCs19PxcLK/xpwM4uDgnDbYYtbVkRz
AWnExmhfJBZ4/uF8hH+iHn/tcJxPar6uwbuxCfxm5R/2gR10iXh4oLty7hZ6XZIx0c+OjzzNHLR/
NjBdtMExdgIwpai3TMHkHxLFw2d6vIURDeEbzlK4aJe3eLd1q5qNsudh02DCUdYjzAgUw+YPiqFt
3wwg0c7l4HZCjoClyVcrADp0Zr21zSNLSMCDAnz5n9//+udeJaeat9BxyfzEJdAdDTkWdC5AYV1i
hSSlytpRpsusleFhf9CQlauMRIkpopzyInR8r0iz42+S0Kw3DLnNoC28Kj+VIpKdP83KZAkDtyfB
dJsQ4S7E4/cPXq8aHGys3uCEYgomYJY1mMLSnu5CxVbszdZQMaPlzID40tUnCotlYnduXSwRLe3I
i3Xuc3vXEWOUtXQul3b1poTudIeCrBDdXYaC//lWjOoO11X9K4ZF5vVAcj02bpatfyAAQRCNntrg
Q6HmNT6RQLfvTIJH+niU8zt5VXcLR/MHD5ZF0yh/sGGa0KFWiQQBvOfohN0CoawL91fNbI+Kzlxe
EyLKDhzevbr5RCXWbC3ppmWEakYQtduENAFd1Fs768EIGWyYM5x/Iqv+Ef+iKEuER7X1Nztj4dBd
agt34aWb+wIWvxDr15VPYW58MqpMAO/tWymceadQUSVVnf4YvPKpRn7DHSOLuppf5zod+c+5pllQ
cWyJKv3zIGIbboqP3ANNINOP3m9OHbRF5ghSNu8MxK/xrEjeDKY8IFrt0n3jXUlRVONquqxkL5EV
VgABSQ1Pu1UPF23HijCBLey61tBYSYR80vlJcdBzo9Wajteqw+LyTrjh5ehVBLtiTGxGRo77JI3b
RtuC4faJFiOVRdxmLWlax1ymwK9UUIJnaMvygLW8qZ3sVlyV6YrsWRXq6v6r+Z5WBYvcLDk8+kup
RmgnrNIIpHhraU6j6Xaa+SXIy5TLARV2eIt5ZZ4gE7/Xix5kP7JDvdYtkfzlpj3AI/+Qm9RW8aJc
TBqISADyg/ThjUcr97BRTVAiQUDO0kQnDs2O6U+Kg3ULPwd5I7d3MTiVo+cmHQGk7lkKuRf4wBYF
2ZVjhZUIrtsQQfmNbITCaFLP9rs/R3qF38N8BsdeuiTUDA23Jl7TvCmRIIOtwS/5Fi4RFWNY2Tlk
9mYKqUiHtqH39DalO/HTXHGickW99JbR6qzJ+ecHM34xM5XHI0kGeL0ZyosGCHb9U4hcy1TLHzEH
bfRCQjFhPoeLQ9b2tAsQLKU5oc4RF25K0I+iceak/uyc8S6l0lzX4edWlXKNOrmRuYvBXmltVkiU
cv07OrGprqdlzW02BJ1hqhazHzheED4AyLhqjr0mHM+T5gvfwjlWtgiVQzJm+NdzcsLVENT8xXXb
evSDSlcTkuR+y7LRvevEucuEVRbKH7OGHr+X+tkHRzoDF14g6gond5LM0g56SU/gymCwYCY15aza
jvwoAMhOL0uypppWTxRy/Z2bVP8/eTvQYno4BUB3Xw2cmcBQT7TJnIj5uUzguKlvG6PlxtiAN6Wu
nvwLJep1fPx40MahB8E7tTpoLjOsaCBXIOJu/pY5sAwKc933Rpi2qyxueeOlggfy+NRe1Fm9UQ6L
5jIJGz94btYYc+Wl+JjyulNv2bw9W24ahMnOml5a41xY6VG3Yg8OPHcY8bo1t4DS6lZojgcGaz7e
tBFf+39lsGdMaQKqxA2Ou6SFrgjeK1ST/Dey1KbApC7VsndQhGEnsLHfwtrxNltmR8fo3Sb9SS3h
C9sjXfQLeRii/UGJJJcyefLyaISGXf5Y/1hpK/4SSwM9qFPpS6lBVqxSLcs6JGF6HRWoWNr8g4D0
2kOiGXFeT7sWOQvcYvd9DxX/RFPRdVRNN5bJ7fjjdbapnQZ2t/LF5OYfK/QkOrQrTxd89e8H190U
IUTWWhxHXPw6M+VotEwdkC8fAFkFw2i71HPcTKmx1qINW+6/uLwFpgdEOhjilniUcemd7yxtGHF4
RuQT+UPFlpywg7gkklGQpAuCHq9cv/RHNjBXfNW+0aVAW4w+H46hMfWM+PQEeBIlIqCsdTyk39h4
dTHekYuVDosusRhw6pxw0GJ2gkW5zwAS3Oer+fr8VdSesfiBdFq2qxsSN0JnaAI8ITCBLCSbgRk6
aUaTyniOSTq6lJ6mS2Q2FhvBHOItqfo9UONB9VSEmYFdmO+Ya8wHZoaeMk+aoBbFtfaeGFq55l3L
ZAo2+aIdSGoYKWUFl6yG+L3HLxHtHYzMPzimZXj9I08f+kFbYpmH6o0aoIf2y0sajKsiGQ8JRYwD
zelAryk46l3DxAgRumsyXAyBGQ82itsWZAzgRANkNi3LQtqtIVDwzEmV5SLpR/F185HfNy7irJYd
tIwAEp/SJKKImlNSlGvU9vdo/G1LMLXiVyXwvW4XC6dYG9++la6MnKqZDi39oQrAAUTK1rYHmuuI
dM0uEOVigFVtwlbZMWwcxCZ5PM0cBkUpbvBwFVLGUWJ0zZALIGFOtpUdmaFdDtLI5igQGVl++27s
jtch+EkaBqPomNSz3O/iDlvdpYVEicNC6vhRvOXvmXb5oir8VJzvXiBN8H2IXsIsyh1Wq6qEiBiV
7aedpAqWTamWfxMX9htjApPNx2F3VwA6qnIjeY4ZuizraNmRDTgcmqoQyNmmQ1mZfMcd75B9oYFU
RjlrFVu5ZKhEuAtCirkVNBoB9rP+kcGDV319qYqTdONnGWGXEFnvoyFPgvU50npMSZrKsCta2Ctd
wZSApXiyb9jPib35KWatjX3wNXTaSTwWm3LGjTKR7hOYE6uRzEngHnMFX44JOI6+QTw+ZHTl/VEp
fZFoZJf+y572mHlYgIiIguyDlr6bXKG43S17BvFkjYFZUbEzY6QeZ2K4jpl6RSQXnwHrU51afCmv
xEDDqN2UoU2uBt3bN2HSk3an8nPoQ/H+e5xDEII5t/JCDLNDgDEJxDnvhYUU5ugFKxB2dttjHBZv
JZU0c38NuQY1yyeeSQWk93MpKpFx4+k7KpKMQuQJt7jRUwSEa8aekSzb+72eGSFZkLhZkjum48OF
I7LoVH3WgTiAAfDfT0nkKY42FhnJJg3evHnQlzuTA7MfiqeKxzM/gCXFYsx0yA80xfIUuZy4gxAe
e6DzCWWUvQvzoE0gV5DqPpiwYsh2OwxvVpdjPYiNYOLHZO2ROBL+jf3AeSikQbnayTl8h3L/mHm+
kVq0tK7licMeRdLDHDjQx+Rkqa4EjJ2wyEfh1FbGONkFiYSwhCFQ3SbT+q5QXfYOZGV0Kvrjwn+S
g3NfDJvQgytytk6xmkSxeWJRLes78UOtvrZTHDiRBBJPXQLFGxSIV9xGPTdlr/c8OyDnkP1+GlWp
BMezNUAPqjM3h155oMgsV/Pn026ueXxLsrTshZ68BQqRq3wvdDIIYYReWOz9VV4ovmsJBhEiBiLj
XO2KwBg0QYocVYuUjy7MkiZB7umc0zBcmk5BPGo+3VUMQUw+xYJjB0kgQ3Ws7/kMFDbcLvX6bwYv
DhYiyljZGTMXkzzgRnkS/td6SkRWxJjfN/Y3vWqlKKxTvgMt20JWlBfMzUzISOH3KLnEjJC1Buud
731n6jxnmXoQuASti2GyRB6OkxudIjp2P8V4quyXMMh4d7QNZx2vW0NdSk/rXg94QrImugGQwTL6
z4thKXhghVcKyH0ZZbW+pvfdHAcwoTduqaJyZJUMsY4hG2/kdYm/J2OCsvwExE4oMSjoQVGL081c
qrgda3NrPo9QIonmIoVwjy/vaHfbM1oqg+KA0iE+MOOQyAd+RUrxz2BB/gYjDPhsngmXV8C25Kwn
rqazNnULjeF2IYOvFgzTBQB/fg1i9XyJpa5s8Ry9wZUtywamoLkSR1K7PCLexet5bubiWH4sqTi8
i0/63hNHHW5MP916jtw+w7EFYweeX59Fs9HUvPNWZNYodOtlkWDukCdwsIH9jqCjxwkpj1Ps/UoD
utOeyqz0JnLV+no71/jNi9tsodZrfAOujAXSLd71WPJigKmLeszMOJfN3/dj3QIlZq4j82fIOEnN
jC5GnthaIg9d/bGWGTihOppj6jgUkFXHazji7dfPO5O5k3Wcmby+fPDvuxTyeL0IRAQQGGsgpm2z
SjqdAIk0zyI/Uuip47ekMzqCWIjhMUE8Kk75GewJ8JB3FdMf8BLTfNJ82IDiQgzEQElCo5R9LmRM
6/+GakMMvZGj/QOGXfucYSG+1sNfuPMhM+dPQklkHKBjjbLefF/dwnNmIdzmGcrN7S+VwILG7Ezm
shnJXj6uvSVj02vL8zplnCxMUUSTTmFh1J9n9nALB4jw8jzC25Mog4xARtBb0ewlGQxqhW6T0leq
9/1qX1etxEWmvH+iZQCU1QG+X6l0z2gYz0/DdNGtXzZWuGJ7qa4NpSq3BcOC2awNbR9IRUsW+HTy
pEFsSkiUcHNRwq+fKrb+Rxnko82GtILf9qLnkTOCid37obPZuscCtNIz0P/Dfv6AYC/oJRudC0zL
yDT05y9IljiEQPtvT3ZacGWD3P1XiblgV336q5zprMLrS43skUWbh0ictNQXZIWqo+i80NYg6hNb
tguKF3sK6JwsYX7QAo/H+BE6ki8nbK2YhuVqhWbM+6ImRQ0Vws5pCvNn+g/jSsF60hXSxOQrAmUc
WoxkH0HmvkMOKgCfmLmk7RqsNQt3G4l09dpXGa0+xZyDn0BDBc4IhtZXH2ga9hhwuhxnPtQ7lGaf
elfHdZ+214Jzm3HdeT+jw1EkB+ZzUqzv2qLN286Df6TShnxkTK4zi0Vgy8ia1+jen7i9RcCnpQN2
3kik3Ahgiy1Tbp5+8a4DO/kwgbIoMPpO/2JEiHtexrKf6UByH1IE7Ic7h8IcrgPLonnQEVIqZVrn
NSNafltcFD1iSEyrPTYHWBINXqhJNSwEhLKXeHP0x+qnVKEzFgCcCy7v9GmvkatgA92IRYjD/yTk
60JTdS8XmGOj4JJTbBPe+CBkpovCQO9XryzJzdiSKsERRCDNzlocr4DdBVn5aVTgwXo+dzBIrXeT
YUFVt/f9xaE87l3Cp1EZ8Wb7sV7/WRSsj6HjxC4ZLpUqglJVUrJDmMxLAnJvPKB6/yQsj0gUVa4H
QQPgq4rzFsmRbbHR4LVKEsiLqNiGbeV7b3jdSdH62RgaW/wxvflU/lf6SOleaFUQh1vi7aaT4Q10
rkos3bEQ503LpjRzojCG2BKxDGhpaG549PoVkadKHBbUUCezd55MjR+iVlsk8fH/i/Cx4VIMstvd
CiSD/z5G+ZgUxXhFMF4uOGpk4ypMgQrfHKun03ncxsoTBr3NcHZ4PhLPRqOufmOJge/jMspemBOM
7EMUwxAroqYZzVZWNJdt2n6qrelYIqtZIylSPjBn8KLsVAakW7fFvqBTGSIEtUmz+MBRo2tSJT4h
Q/PN9VxjOg9aJEXwPMW3l1gv/AmNGAHfbWYMl3TVF8PFBZ9o4clcvKQu3s/6soRqSGOgr5yJd9m0
2hnsbNcHxbXU0ZyPyNYLdkY/rbkuu8cshNK6dD1cgVVEhxfpdjwZ4AD1nmnBekeNNQCBbWqmB5Gn
X4MNMzlyV6tF5Zx1NhnbrbBWITDPgMgHCjDQWNytgWddI4KANCPQ9+V7HYeF8xDsbH7yPfSUKfoH
+EuapaxmZ0jQtyWeHzfFfEJWnuyssJu2tINrAOX3xgNdakD0dFV4qmkhjA2fxmw51i6D03gR1zei
9cnbVLuRFxjR/plsQ7rb1sFqPhaW0rArGQ3VjSmD4lyUY5IiKrQY/3dJAoocd4Uok6jtYF5MztpW
TAjGI7pvvK1/doolUEolGxoNja+lFC3iKBP71I5gfHuVt0dGG3m8u0c+KOWS3Xi2Umh7zjobVaS4
tgLSsbmT35uHshxNQxDBfgG5/uhXh72kHiS3hUYHPZBowRKEZbbTuxltlrdUNfB6jEG9brDdI8fp
92soHcPRG0EeIjrNqDRIGV2kCDncu6s4EGsD8ruBxfT2FhLv8LOskFQ8EAxTwrL3hapxRY9WtCdD
io+qyJ2BFT7lk2gxmJffayTyI4cqTcQ3DSQHKYlycjuntxkAoHmGDNKLJcE5+Ik45prcRY3BbDVB
D/jGH763zL51FJhq3zAmUAtSA1v1yRr6b4QIeKpU50nIGTJtqI6xBNBegYIn0GYUT379H3VNVjM/
OU0yTP4eidUxchYhSr5lhxd1A91lo3fMM3uDLDF3ZR6VNfqFIKGdixPV7j18pxVihptP7kXbk6B7
htidDA6xRH+5gSjFWUxM9IGj1MiMZPFmajtCPXTaN8K8d+tCW7LsxJOJkXQGWvHavKCHmnAdxs0h
GUAZTcHVczuTp3F5pgDDdFfv4mZ/wjIXp+tCwHbVahC5Al43u3JGaAGFNEMg7Bb3n+S4DnM6nLOp
KUC25HFPELuycrLbYQ99TgA3bgNgYYC5mEvZr7eLlNCoB5fdf9uBYlfD8FF/YaezAxh+saCHtFcb
PtR+Wk1i81uIMJGWW1fzJGt+5YOfKHe+xcUMYp+1BfCaJWjrN8NaI5gQHHkMAUbUNXZ5upyu+D6M
nhIbQG5fMrAOGh9qe7eTehX4aJmjdvM3U89/Hc8pHx2UXwDzAsdRT+rHqcm5x64lTOWZJcmzgo/V
zcf13hARKjw9bjpcY+p8m2VvYQA1EarmQldZ6JJQwx97kpkwaAfpU+VeCXoxWgDgdm+w6fX0PnGw
tP+lAFazOVfyCiiNJr+592uyvzswdVWFK8llgbTcokdVnTQFoFy3hHO7hB94SWXFqiLgh19c/h8X
j6AzLV3fBKnePXOYPSOWgJL5E+6Fw5lOHJFfb9EUvgfg1dKHbrZrPbY+TevUnzB6To8rAszuPZPc
66LuvGliOvmA2JCyRwsYWPPIsq1RDH+mu2QtoHYu3KW+FFJ4KY7K6Q44jYY3KP6IzNdqpaghd7CM
KdqjluBd1w6JrJoNv5o974HHNfKtG7zdewD0GLpOGaaZmX9IdaB45YVEJEDZ9Wrh6k9a+IBTO2L3
6YQ/Jb34QenaPrWhu8I7rW0gZDlWwNmiD+tZdWXPfFvm3zlHFBM3Xp5CspkN1n1kw79hO5IuPP5a
TlEon1mxoBRyPmhm9GcxmntNO8r60EV9qGPxIL+C7GMUvrJdSVsMKtXDU9g7rfhnROmt1+DVfA8I
Z021B6U97QqT/qnw3i9r8Ww5ZG3prHshB7+JMcHNkXyVJDN9/Co9gjy0l2RpIvhqj1Sk/kHa2Qq2
UgAXu42e/dQwdU/TBeA0/9bZr9Ej2SLPoY47OAk6zvqExLoMaluBfCw7sMhSl9lZ9uWn3r9a498C
4cy8aUiQvkEceEtVLR7CM6J5CDYF4nM0LF+bhcgHyHo8zgdwsMUsIKroQPpMo5gENFIw1DmwO5Fe
pLe8sInsOP74klz6cwtM0KzTirk12rCUDkWQxwTljv6sTfkEFJnPPrul0xk9VbhGsl0/lG7nkhfy
Jt9Wh3lKZ3DpVkrzDtECZ1sEuemUUHTg3cqujoAbdAR7N2OvZf9BWswghrNZeJi+A8jY1XyFGBcE
GY8SfP9eNUWWHWkCVFiP8ySsttNKQUqUh+tj4qsQGFWpuUFif1w2MTXxlyPzPUJ2IIAFkovV0zxk
Of3ocri6LecdgC3qNcmSnkdFsgfQAgR+UEvuOCSypeASwl6cAOgS4D2KOjsYgOoS4E+Wwp5Mm4Zq
LrmsrJ+qiCZdqZupoysxU9LZz2radDLWZsITAyYFyWQaf80ETopW5hHRo2xUQ1tQk0FcRPJLViqj
MHkyAzTWTZ9S9GppZlsQ9ORxBJ70qQ8/yPqJNxkLMzMN/iGGTak5CneJMqHXOCESUyyxaD6ZBIF6
a47V3Qwvp3cwKDnUITySNjez5/nkZTbtLN958h7Hs/g4OKkPwXUIuou09TtXVk0pn8PynZ1lNMbU
b5jAijo3h4cwdAdrNQdUmlzDSQ2M/SY+MH7Ilem/W7i0MqkkOwDy4OZK45Nk6KVQDpyzgz3K1qgp
nmaCjHID0Px1x2kjtM/dirZ0HvqLNG2DtQ2LbQjlnusN/UVlG3QM21wQFj5ldpFUD3b6LQUvzGOF
Ti9rU5BGJfKxl2qYJaxG0tyYv7hrb9ggKZ06EMRIAkltClikFELu6C9Dh2PeW+60cJmP/D4vqcI7
zsNvkbRxch/MEEmLZ/YnsHVH1K+mGxuM+zoZrW7UoL5A1/m2HQHSu9IvSOpZC5hmSj+Ic6PXMUVt
ZMsO09d0SlFEqiwL5BeqmIalp0wlH/jwGU6vMFAt17SHODgSan0U6gGLRyhuUW/Nb7f79yDndMoa
VcnfZ/aPArC1pcJV8FjUNWgs/u2fwHcnw8gw2NJr/NPsB7Ci0uUVp2+smQQn3dmsxcXNKWoaoblU
720g+axyZPyfj5e4euirBRM+xFyAedxMj3UU7y+PuqR/RcAGdRM6YM7RjMpXOu7MVvWcklyATdkI
iSpeZDzr/w2ml8XIfgnrHpWCNg4L7DEDBAveN0lvWxmkgbGyD2NkLuVYQmAeMj6tmWFabwG8MZjG
/n8wqOVBML4etCHcysIVqG7HHRJMpQXPSepuEHwzFgQCWDT2U65H7ZlYkCyPaZIZ/2K3Xb9T39N9
d6qQLrjVmmToglYFm3NCbeof8oblsQFu30LoMcmRqnlvRayi2ThuLtM8Go6XLJYeoGrzCbZ/U5fZ
qbc1GgdsZBhMWHkj2mPG4Q7kEq5KN2BSHS6mwM8gd/04UV7dVOmnYbbhWWQxoJxseOBXx1ZXKsVl
pwmSnFvCVlnuw5xAWUov4Bui4DiaF1RqGVAdK3CI3/lqBoeKt4JEwYVwLAf4Iys6f/ibl4LVjGAQ
496sX43OvcwFl/Re7vt1e2reknVQknFjOTxStruJohykUtcJgO1tgTu2m5nFQb6NaNL0gWEYVcRg
DC9fAf9IKYGrmgwFFx66vmCkdyA8QqSB2PV3J/PJDtYpsjbfJYeDrooBVMd2nSi1CrGwiqCfox9G
t0nuioEemYkxGrARjBIYTnhFZgXRXbthxNfiP1Vwba8sa514gVz3PqRd56IofIpugBMYkVbE6gtn
x6ZH3fpUeKWq8ZFa+LlBRqhp+/lLfDApnDwurL4GeKph4XZIu8yRnEa0lga1zhjN/dhVpsQ5mGBu
/wk00UnnfkMxc3jf/bvdlHWBO/jMV+njJpOyP6U3OvEaw21X/9rCVyV1mhRUETfc3ZmrhQNC/wPV
E/uBt97reb+yyhFns6TWJpywQo+8OaPKwVJKcTBfUStkcPFhKRxsKJ9lWAyq5IOpnuPnQNf1ZBgB
Crm8HIC8CAF2f9yNk/wpEkf6ohOokCp6yUFiHqy/GB6ANw2k5O9BksduKM324dygYQEkqPjvWGAB
l+GpD7QiLCD8LKS+c8cXOljnX5fr/4VSMac2t24a6ZCaS9/j2esn90KwIx2iszr11VoF0swEktKR
ZcxgW94OO4F/HKQDw72waqindpzDvgsSLy8oJ0M5jycaH/arBwLidN2M346jgPp/9XvfVwG+2oI9
ruzymhQDMIM1SHOTapZ4yhLGVxp5sw/rxUA1wvmzjaExfa83rt2kSvF+jiIVJVGuFg3CJ29lWptx
bnYFqMMYmOd6tQlzwwHM/89EEvEmxrXDVWqc+1aGXzi2nnNH8L0jZJcRG7EApicSYyr3xI1OeiO3
W7YwTcWL9laMnUOx7VUekaqDbLKzZtEwgYRsw/mGBRFsEAjweV4vLUdQtwqnW0MDidz32VydX496
0UWkRoWlWrSgKLidPwszt9EY7QVN9AoU36Z5nLgJX7io43B7n6bz0AWRvUNHX8Kw3Su4PpLCQmfR
xfa2DH0YXP9GVPtCmdy6zBXYi+7d+Gty6fc7G3F5FTd5U/ehDFFu09ZaoF0oJ63TXr1UVpI0P+p8
OesykM37tuZ0/KcFhC5DNPskAFCuanhgmu3ZsP/3sZibjAdcalZWwvr6l67UBSXNyJBC2J7mMyFe
H8i+t1d7ViNR9XD5LqHuMb8OpFZPOSm1bQvFS8UgN0HsqpCU2YX/rImojiyzNhgg0adfKRNqI4Gp
ePA+9bpkGK6JDi775ocf8GTlxg7O/P6d+y2PMVK42X0VEuM8pGZtnalNd1hzIM73y+SDBFqc92o3
oEc+16Yr2axu/STywFcMqL9MwCLE/bUPQFFfd84OvhmuEDYpmU0Y39b8fBv7tHNe7E85Jm82noFK
fPjasp/gByEwJmg229Cq3sEVj+GB6k72K0MeqUjq8T5ky5C+LYC5DaFh3cD7Wx3SqCSg7YsyNGwj
Qvkj9F+EACvhKN2lk1HCl+NH2XEa1bZlRZrDun8sY1mUbnmZFX+9GHWBhlUPSk9H8fCzyEbU3g6q
yV33xwo0Prb6iVL5F/p6Ofh1MQ6igBO1raj6aPJU8Neu/uYyIKVoLTzuvg2C4WQqu+QN2wcblQVZ
Z2AXzRP8TqHCZvmG0dskGGBkMSTKGqC+auIFHF3oOtZJCEJbTjUdiSuzGWG1GU4gVpcMZP8AQtji
Eg1D96FWKMDDoNE6gwHLGVUGzkczp+99Wq3+ktypkInFe9HSQHMXTZQczyir7eZvtoP0zkIfw2Dl
IZEJkQ8lXJaPiWd5U5Sisoo+vOFsxQUtyjeMF4EfD8lzySwnlE70zlqZx3HvOoK85KIf7I2E5SJF
tTQDl0K1r+gk7UWXxqIdiZ0JWSGrzqOKw4npZJDY6yCmmoyAb4pkSzNcawO2jqg/eEsv2KitB7qH
Nlw2KQeJK+31tY69MmkRdn9pURIczv1hV1xxzNTzJLzge5aHPKiUXtXv/S9czJHzXJQDdCC5qhkB
Mbuzn2bMKomymM7BYJPjKh/JbfQSZCvphp2iPcSvlfuChknrTlHiylJh7Hcl6IEGAmQ8UJlPOL7b
5CHWPmOiD8bAVvoe4ZEV6sFLjd/5UMy+s7ahkpiXaeKoqBT0OZKVKpfSimyGxo7wu9gW5tK/KNMJ
kZGUnFs0RoCv+bDJnirFAObcBw5B03PNXmidSe+WjK6YUV7fH56qydRd9x9157hn0aeZ+mjsX10Y
f6+/4dQ7+aBLHQf4Q3mk4F0Su9KhUpmfhv0RHdiwi4+OPbYd1WT5Aj2X3PNaJqgxtV/1/c5cs0Oy
BVrS97Fyvf0rXWNBZXKoRF0fSf9GSJcBc6oHtR3+l2bwqwI+0MkO0pAA0CGVkbqnuSrS4OjyzR6Z
n1Y/4UUF/dFGS957vL0Xf6iR+YDuV7R0bXGFXnSfqkorSI6dkG0iJYuaB3Jbedo+pD5CSxEiOna8
MrODzrYe/BpImdwJDhLi/cyIvA0yOTVoh3kccTPhh8BHFfU7bzHYXwsnRgBNGpg2qvZZNEkRDU/Z
0wJMqPTGXYgVPOaqpkfP4HabieuBJ0OWBoNa8FY5Z7dghDhPJZW78N9dVzoHHIR507sXgJ0xypDi
gXf3FsAWwOvHKcKrsRN4KngNclbXwEbSr/LnDZYzWOpWiYRrr9uvIbu49yQHndubtblbtkRyNjfz
WHnBscR0Yc+JUOqCaBz/rzrj66Y4m+X8UL6/8J2BtzJaKHAHz/5BqyII2C8JxgIjoyW4sTBuM6aw
c/sbiypgOF+Ome4/zSe4mxbZQZXcjKgZqKrNntS+OY21DURHd3RIdnSDx1mSh5t0NUhO8xgoHCsq
44Xh1JVG40JGGG+gI6oHQ4BMwUfJluXX9pY17QTu8lTQtNJpBtfLtTFgEl/fwhC+B2ZdhhkHh8NX
3BXDy+LRZpg5Bu+GlhDTI+roIrucLMFVkJSDN01/DtyY3fhTO8iy0k0FpZPW8PwhXVRL4hB9BpLG
g3oMWEPtZTjQl+TWu9y3Vdw9aFb4z11WCx7jQtTr+vDOQlxYjor+ywfpkx565UX/600FLPzFpwZe
UiOxC8HWUOLWo2NtRRZnz+vbiuvdZz9kOatXpkVvyWe+qcO17YOy0ES91SFd0d5gtp8kO0+l0M7k
Az3e7ioYzsqspxVfrjslQfD35ifhG1zXW6AxonF2gGtbyMq+YOL5fU2VwyxUItaj/6N2xA42cAFe
Kmz4B4aPQHmEf2nvcP9ktZ9Ly7xeKuO/M5QxxkKiOCO+aqQXmz+5eDlL2zmZGulRJYoJ3PxwTHae
HC0Zk03G3UeQbLpi81ts/WdponhOiVnIUl98oFZwQx/wrZRoRe1FSyQVDTQejmqgNxEG+3QeYdLn
cRkSBu6DEDqjRQd2wjssBlepvqSf5HNt4aEASSA8ElkBMSz5SA2zr35md6GzZ6lWftSgXtMbUbbR
Knm7XMGeRXUdwLkUUijkyyJOPaYL0LBn+6Xh3yihzVs3Tn/LbUW1Ac81XiSKbrbgyT88qRfqiLJn
nw41Jpkpxju/9UUF3jpb8ecZSsdswI+UEYN+c0ctHU6Tlo8pleX7bJg5lbTlrUax1ccVI4HrIm8C
7w/kN+ifU9GPFxlUVKO28z0g6Zzko+T0FMgKv8dTKKKKgrC3VvAQjtgIr8IM4yRSbXFw3I8z5Afq
BmY8ReGCo9jeevyuCuSftMwu+skvmXNq7uUP7WixLPKISalDJnxckLilQsG5h/jJuHVTQPwBO/5Y
KuD0ABtgrH9n7Y1OOhgVbxRTu0479YXCOmhJlvV+fffHGxNir6HduJUJL/6+YktOis4jytZbXlNK
FTVB7RXhfcbUkvtqih0+j6edl3gXNrLFXa8GADBraz5YynhJyHr+KBFqGUQtGGbIX/sMexAZ9RpN
mxC+1963ilqOah0sJSLfvSMCt23x7iENhXkxCJhi362oYxWSlxrgiMLiD25q96kTXnBL3MOl5ZsK
7gL158cWHi83PN+JbpX3fwgbP8YShUO7E+CmQXLoykc6SYUOhCWS4DGqZagouR8uILETaOPUvMdS
jwcwGk2rMPSWjBuMhhjml1gvcfY7qfoNcrD/Y+Zs/zly000Nx3Hf4JpmkXp1fORd81qWkwQVDtW2
xY31yhXVy6+SKIFvnyckr31aoDOuLeTq353XnLk93TjIHMX/7Y77ZjfMfkKmyYf/lcL8A9JqGi4+
wAbw3Qs/Qv6F1rdtODJshj1u67xdi7llqBSW5Yc1jK7KK5Kc6ZmKYhjThhBAaZyb2I5aB/wsbMAa
IwDLuTCHRYkQUkCQOo/8IEyJRF92Q9eSCfbhzHRYhXI01V7ldKHFuPZGfUuQCTUi1G+0o6T3F86a
f+6EymL54h9oTMt97XDyREl7UwkVVeqXLxfDNtB5r4BA29xWeeKYRInFiN9Vzmw/FbPxWGAFUUiM
i513+y9ylrGgx/J73AYYlxvWLJD2tyqWNqkAtZB+L1EqAm8NQsX84h6eZYb3iF5VWcy/vDLwtIxt
TaK+m2++kB48XXrHqrl/LBjNrSlRORqThh445pnh6cMmeLj4kMP4v7pSXXMAiXz7QO3NT9ns21cz
P/93rlyTp33UkPAosRI2m1Wghfu1Xo4+Ayi+TtCBQVwDBq6+Y8aSCKCk3N9TDAVLhknxOuaqRDIK
19EAk1Cg8c77/Js6qvIQfKVTjw/quo4043xMTx+ly+N/RXY2Q45kljq195HwHj7jze4XMwXNzbic
p5IAzpaUC1rlVthdvPNhnkL/Yb7pHHPt7T897UqlEwEifrjxLHue0z7vmqbmCHssvAwTXtAtiYca
fqkzLbW3CyO4zGqQhNoLGPHQSU6rfbyUdst05icky926XyX0tH6HeHBUH83dTd5R7k/TwyViHwhr
AuF/U5MNyosSgRm6IvQ45Hlx6Rz+I2TqLf+WWHRU5AbyBlKnN9J/SQQVuZE4My4AvypDtKPDJ1vZ
ww03qQ/Vba1SF9U+zleef0XGk/3s6ZUQmx3I05af7mT+dwQD4Y9fQkluYSeMiQK89UkAcCMZ+EfP
ClTwV8lpNJtKE6OHg2aYdtbAf9Z08L5KpMZy8U5w58HB7eGL4V46Qd8ZsqhltC5qUlNuYkX65TWg
JHKhjoZBe8m4pgVjXN7wPIQEKbeS1NLVe1C8+hICzd8Un0GpX6lYQQiy3i8VqHj8cYtaQm2edJ2h
xl1tBjAnu+0M6VwJaLo4vZk/uKoL4pJJO8ZXagN9j4O95m3P4nD6QcfEJlTiv7QCsYFJ624Nj28M
LSI/MVdOpaRhDQawJX+oTFYrToLp549wKne7Ilae6ym+NWb/6orrzvNPNLe2S2peGUB1tDF+vnO1
eOj04BrOB8PYD74Tez/XCEh+z07QXzFS9xH/kVeiUOikwIjfbfvzYB9pluawX3ztU14kflNA+3Re
vtd3Qmzb9y4EfXrFBfb8FRv2Chf1SiPWB9VCAkgP3UPnnlg8JqFO6PoT8cFC1nlfIYoe5I8b8Mwh
3+eYvminXN15wPSkS2ZdJf/9uSldYNjpjwdhN5Oyjml+i8y/n2SniVG2f1V/oc3FTow+UnzMts+6
4Zc1TxP5tH2gQWKw5qtm96yr+yqdBnEHeKkH219Cj7sfJP6Ne66wmJjeepNxX/pEooQBPGL/m3W8
MyNZudNdH+nDrWQn6JPNqCcHSqVCWLw8UzV+O2yYEnqok8aDZpz0aX/Yoxr5VTs1xSk3MH+uVSUQ
tT20wF0wvClHhVB4cwpw7BQx+l650eq62JM/wEtjM0CHPGIss0hFt6cB3zht9S8eC6wL9FOZtT++
RLQyoE3d+GE0tN2BT81molByRdbwVHIOa2SpTdcPc0vEbjweMmaU72rcLiNnPGoasrkL8ex+nk45
klgrXaz8/bB4l9vwdxntVOD8UiJCmCVsC7HUhzH2L067D627Ao7MtpywwqHFmWPCsV7nbG7oxFbc
hSN0P6E+QuE6tJnHrwbmfiLuqOSNxc3bbagMIcsx0qEop4WwQ0c2B0FGDXGRsQ/2Ml6Kd5zvJlGC
BWeVVmkrN22oLpEsR/NGWYEpHeYRtr/G78dH2Jbo0NyCLHWP56XdPVh/ug+VAR6x0j1nTwJmc4+B
a8/XIObHbnLz4ob0g991p6d/Q/qxuUe742OaNEb0JX530Sks4p/vYz6QnmZDWjUB/nkE6Pko6cYH
lW/cl5LD0CJaQssH88lIRFaNZOSo1ieqIhAuHGi4A+ZoekbuWrAmyot+h/M14MHLll5KQfOsoL5x
MsXDAtCvwVbxhSNkzf5c/j71f/Z6oHiH/lhM7nyd/nlh3VWTW643zLp0+vnjLOlKFX2mWBHGVBSj
grATMOnTcXJIN7WviOjbxq+tR8gfmpKZNp71sZtrnJNhmSC4N12F5a19VSdxrzUyep9WdtQ1cbjS
4q/oxfDJ7qEu55G8hyIeFr/UWaH1ZOgh+JrI/ocKkI8J0TOd3cP4bTE8dkspsHwmVsH9Co1N0C2g
djtdo6vMfCcxWWfNKrzpFasTPtC4NRN/WtzQt+mBstDbhJvdWKqoXpPpSZAf7OjNrNmIJzl1r0zu
yAH3AVvJQ7alQHg2pI6FZkjVbR7QirOQIrIMG5ztOIfqevgRykkQBAqKnXxB4M8zfqskblh8Cco5
knBtu37PGVY9Jj8Am0nvXfmOedPR8MJLgIWvfdlq+G95fqgVWCPKL5BcxaMG0IEuxmo9DQEzuJFk
ep8WwltWd2OMSvMs4R+0UkH3evJ4IaI2sjKt8dM5CsBpZ/MosV/h0JWX4bcc8G1+Z4v70qpGGgzp
L3BniE9o0u0YAYtJORQpikZMxR1ebAKXuWKfKD1fH36TAy/XCytQdasvMMwR12bSZjyW5O1vTLnW
xwjdvZgADb6R58OIcqwl+JT9uxgvmmAyC7SVyIJiMg2bT/ap+DtBNOHrR8ME8jK9GZZfOqxKR07L
jJJ/r1fQ7Us1UEU3t77mxMxV4Td7rZjB/GSpW+5ghIZj8PxgNJMVfYbGfJHhnxAukpTl2f5/A1fx
93QwAumAbIZ7ZQxpoWnAMCpa3KJV+F6NzvB6jWVLoFm9tQCFuJ5Lw904dBXSnTgk1PQL6iZiUSJf
qPBaJt3QLtE878csYBkJ/DxTsVUGCTelkO/F6y4RlHYas0ihlI1TeAzpzbvV1puiR9Vj75VgrdKp
GMynmZVcyLBLx+dP3eZLyJYrAe2QAzfaYI4iWWOrN7ffwTvuGzXXvWc3B1N7dhG9pnDMHDRdJvWo
hKKWpvc/KRhXEatdQOZfhzLdzl9pZkY4TEn/74cC9+Ok8/zGC/5XhtzUz2rMDBqsd3MH1ymgQwD0
sKlWph2q51FtSh0ZEJA+6D7fg3OqStzic1wLOyiVMZACakX0VMrunjbwwBFye4V0+lkAxK7LvLKK
VZYkyvqd2oesx3Wd1VUL7kkwTUle2qmednZD2GVhupwqOCA/6/QYgpSRs4wjqnBrN3CxT4JfxfEG
BGbd0atyC+IBuyRyNcM1oaxeyRHgr/1WXNodgE+14fg+iklCTknE7Z2klCjqiX1038qBom78Yv8S
zHCJXzlZeMKzc4ES1kP3vycSWNMcdVr0gQfxSiygp8qMVjQOFmSHEo1eZVyokKaeJCYMBpDCP4+i
PYjqffWhwyki2ZgOVDGq6eLpGDOaOqL8vkX9JxfaHzVdMA9ck9kruWuoOFqquOy9X0GvSohLLISx
okw9x/oDhiBeyFGNSdb9Yn3gZa2KKnmOYhvvFw6MHEXChfpWNxR4INxiEC9GnEWXthtygjiwQWJH
1gjcd8DdZck0rtjkGpui+mUDPrMcYWHXfaAJp7sMsAeX73Oz+6ZGeJ17i9owVnPXYkRfwdBT43K0
AuGGaESAboH5awqwVMK/8c/r9zFJaHhz3iEI/IPWPniHfFsuOfhcNn1B5yJjcSVMFsR69eSJHmXy
F4G3+07N4lg2n5cwoFYWzO7Sc2Lg1HcZW35bTbPeVDuiYijeqBVFb0gIeALxrwyEzSYL8LH0KRIp
u6njnzm1ezAzfgpTRw+EU58dE8wZpYwPBjYNxiPnpLx7qaCSnDAZrzhlg+RCY7VUN2hN//NAnU6f
U9Dq1q9A8agv3U1lm5S7f3ou/HkCIRpND82pRbp3VOYq85RLxeWoC13aiui2On0wRcjGc7qYN/0K
BIDsIjSi3rGzvMZJDZjsmx79KIcupsMbyE9lcR7BCgJZEhFq3GdE4W8+eNgOjJ3Angwl29KJW/pE
MsiY30oBVdtUeXw+GiNLm6QruRg9KzSGrjKLirxF3XB+9g3nCAtSKXPmjyie3WjcVnJDHjSWgBPj
xB986JVZCe811+SbPO0DA8Q7SD76RIF8m7EliZyXbcAdqBpElCzMVC9XPefaq7gwVRyVlc3VbxcU
qxeOX49me9ZLlWp2RKtAaha/PsNAKSoEE7552ag7vsLQO/W/KikHtE3kaQoF6us395ltwulScVNc
ufnoY+Dz6yTxP/uW1fMEeUQ+a203oIsLg2ottijwDx7vUzpVjHN0vZvwGHsOTTVq3HXwGfJNLSMa
Fv+MKKYdnADzlnJHGDR/SHQCaQPzSV7mRNzIMQBJm2U6CcPbvWqUVM7FCk4RHi+k9JL1kUrWiwyO
ckBHnHk2BPrO4Ocyj65aRHvAteRFVQQW2Ze5u2MUyJ7VoavjHAPDpfKly0XEiO1rRFHc0FBQubZ/
Rba8e8bgXas5LuNbsCXuJ/8j3kHq8g5n7bWBjSZ2zwd0jAPH1Gytry+YzHZBMjBkn27WR8/U8/mq
vp2b5GmbUZrebqLNLdBtJ4CkCM4bwLBSrjb9DW/AR7l/8xPpH/Nswio7qkB3Up56+uxo0KyoYzU4
Q0Hwn1HlfzKVwcj7Ra+r7V8WDm/d97kg0DBK1qMrdrUJWcdthL+7Z/LSmXQVX4gjJcRC48Y/3xUV
GQV0XWE0tTbxOw5MV77rAG8kAor2muHQlB4S3+kGVHi5NkopMPyH1Z3W/0T6Y5Us1TqTk+VSSdMN
67WGqaw37y+riFuJqIuurfawwBks6znH7d3EIprLXQ2jjHkCNGt97YbdFwSoXuMJSab1vlvaFMh8
/VIalhqAqYCZ6rUUpCGcLVS2DTxtUnaAKJIlOVmPvD05RnjR+soUirU15tjYjD2CozjI5hr5mZGX
MLdTfss2M8NkySEj7mge9YviUV+cZ48gjGM8fQOHEr3oGABxmJP8KAFcpSECgkbDhTDbkcDwKhdY
L0Jv9Q5X3RT3tS+KpJqlg/APzjX1Et0Eqd9GdIxsStNlsrFmvuMO4i3MCuFO+5UDiT19OoofXxSO
0JBtklB1MnwfeMuMaBO+F2wwoa1YDK4W4R7Qyo+I6R9hbNqT/mfsX2u+d1ZB8EXjDFnr9Pi7llZC
iziPtqe0/N800PQKZ32ILibHyn/oBWNdcD+LMM2452h6NXD4U1UMLZn+8GVV8Qrci2ykzcbNRsau
8a8DW+NgtFy2cSXnt40RWuEwIDrBKhWu3duuweIr9BYVl8bB+CYKIqjLfEVZxhQXMZj7V0YPSdsK
xqPRjR3DTDP7RfHmRQa3Y2kAF9zB4OSHLTkJuPlKcofai9X1mAJQybyPyisL7rxJ1hfYFyUsN0Ag
k/m+vfNNibugqhHfkr/Gxd3BtxQ5AkUUCNe9/mOeHGod9vayXM37EvpEXFgdsLm1sIzGzrEFtn+v
4HC6mEFnt/GLZfQ75pWgWhzZKBzAXXyNCN1tMd5tv5/tzSzlg1g9t8u2gIDr4C+PhvZGoIS+LZIm
Da5K2Xsq4Y8Nsq2UriYMZMXeAmCTYufq+angJNJaRquvP0zYnlh52LaVGxRlJUicHt/LshZOkHDI
b0j2rBHdcPsCs68Ni65i0Y/NU6WB/TqhoHkOdMyDEGvSmzdajmh0PirCxNqEYkNkbkKPLs33rwRp
mAX9GhZP8uPg4YirwjN2hPHRJ+IpwvR8WSBVMGWPiGG1fEiuSdf1zh6MEcR4FYXngfcK7yPXzo3H
E6daTnvzre8HcGsySD3vwlWgXPGQShy3ArHPUR6ndX2B2BmMozMpe7FDog+/ZhQq7fmvRh/OUPhP
mcS5fGav08Tpg6Y/m1m256HuCpkWxHAFSL2z2srvsTO2HNVn9X8yAgO7Bu7n3hAFt+D351VpAG+Z
HMYv8daq4BtOElLylH7rmy0ld38qZ4zGe3k+RiCDjKl5+pwqmY7paUX/jmuPOYtCy4CeDnN3WqtV
bk/49WTdQp63l94ALP3Nwx18bsfjZ/hOYh/5N0gDY7yh9xKy8mIScmxe6lLrmnNtacWCZlFX0qE0
+KA/M2bBV5/li6uu54zZJmfr1IfWhnwbfF1uSVLmNQ9scui4Z1gzHTj9Jv21V8YfQZGMu3Fh40Tg
ITRwbvEFsAG+Pet2wompL96xLfh5chJUkTtjdfsiohlcd0dw2uYGiTv96n4Z20EhAm1Rd6tHxHYf
PY82kPN4nU+3ci8IbfZi8yUulJ/jd/TfCq46iRu8lq6UC6H/1+qVSXzhO4Dbv8wuVcsqvtKl7TNm
8EcXSdKnDoVChHU+Du0q6VGXKOLrfICGAyZF940SAE2eCeDlrOo318Mxtw+aa+TzMaRF8JgSibkd
gPfjdua4lqUuZM2XH/EVB27/gKnJ4QdiaBFtfK6sjZ3WRFLCr6D8bkxjlndcTRBWJLNaDt4byv0q
ci4gqvl97Xmmtp4/pVwP4WaXCLtcYQF+DA9I0f888Yfqss5dMxnKXSRhU/b9wsHNpAIV45Hfmh4E
aSdCvrwfi5W6+E7v0hhAztxxn1VVRKldRRa2wEfktjWveDyLB837CGaWT/3tKLhHYrQYUPrIj+TP
zEeYVwnjdGGEzCIsAk/KxqMm7ax4uxwkcU8+AjdL1iEeeRXqzBwMHMhdQIlgrZORoJcTPPCgoZXp
dBOdtjvM1P10Kjca40A73+K7PjOOF6Y6eFEHHcw/Hx3Z9Xb4MSQNpf0C9mp1qZrT2I/A2dFjpcLN
bSlBVpk8JcveOScTYfsThVRgxZV+POzbP3H/8SwtM/QTI584RNlWMRwwHaxsaecdhdK2xfrqEjCK
6yFUzHObx9/N3jMzQsOQBh6EyTpJT4fHOMlo3Hgt0G7W9FqEvzYC+j1MCAf1/Ue45HUmE3+3gM5Y
TAP1Tbkia0/hrTfNphlNvebnuCHy10CqSaFgxJJicnGWTCNR0TDnDeqfaeipfs8C82m9FxHNVEdZ
DcyyhGvM0ziAYkTlxehTZmQS/1Vq8645YOhF5HguZORlFylrbnmbUP0lwngK612eQ6ecGZ6p6L7Z
naw+m8XeX0SPbwbIk3eb6EXBtCZXwATRLX2HShfI3muoVxNpym07Caf0oup0uuAJfyu4uXhysuL3
pk/+T/GXNFNSBgJgtPLJqdxRE4i6mIEs/8+8EF1ikBAYm6pwB9B5u0TAmwbWcNUpEp8Kp1xnVssG
Ya6G+bZb3cgTh4MUnMZ9yYfBLnSyuWCb51qsvn6J7hh4zVe1blEMLY8ouubJlmZTNJBNWuunyD8t
uJMMIbHkFgbqAiVxxXfTmbMt1cXN4nGo3CRRfzuvA9QE/dX6d69mAGjFLWhp2pm7+Z8C+mdcC9WS
0OJt/pNwiLrFI2faSrAbtWFHZHotPkrItGL4xt1WPVUjPz0OhpT0qteSdnlKefYI+ae5U22QkbQi
VGfb2jHWlJnj4mdmaLodJVty3gaILU3zedRnfTYZkWoFm3axFX6XFZWyY1cqeIdSpahNj5CsWr+t
rUDLmP8yfOrF0TxVpYr3m2Ny90DRoNDeX9Z0jxsPrKtaVG1TDO0pGDd4mWARG8IEGdSDaXI1XbLI
v97BsZxy7HAkbDys0kYizmfFnJe3Z1n5uJZEKqOuRXqiIKA+ANKttLOI/F25jBMH/u62VVcv9rK8
ijRAc4GoZqoU+ven9WnmGGA87OC576fenbXJrz03gj/FUR2QQHhgsQPM4wN5oCJi8PDTlVMOWsv1
qnLZke37mdRVK9M9AYagnQ2UKBdmRzyk6zu6AQh5uar9XpRyGXuCgT7jagmi6aG5yy68cAqBHUDs
daYnThMjv0Gez31Lrp0wBV+rdr6sHQDUJ3TunfZJN3lp4dYAzNihrXQ+HiIzs6IYHpX81tTT8h5P
/fl8VnsaP24IVc80YEVTaTqGxVnOtFClHt/8yJdSLwIgktZtXw8axKzR1IgkJ/RJ2Z6XKv+BVutl
5HQZavi3BR7WBVP4OMloMmem56lopzWsl3NgOllJ7GCEgeYpV2zy7scjj0nYIpBX4rZQja5wFpxA
j5TKsTC1tpSrF7jDu7LTQJaMIXui9pxk+gcXOx/6StGpQ0+4NeYsgFTeG5PB5CElD/23kxS4MLJw
d1lnn2RkFzuF+wkV3HzLZlySJPjPPT2LwPiJ8eJIM29EaGu5SWSc+NkuEaoS57qZkGOV4to5aAm8
CUQ2DtyDxL8jNKk++fjq6GILL8uxAZvltj7odrgg/RJrfaSD3QbW/A/OzIWWAEUSpIR1Vr9wrq0G
tBsgQfPIJ0PRT0FcRakzWgiSCYVmvcW1O+pq/Q/oYzbQEp9g51doKFywvnFuFIP7ZaxG9li+fT8A
JrP1tsD6sCvRWHpn/nZiMzk4vQral/m0PNVggXAUjKiRMUcoSAdAHK1LDxL7ui5JlxQ7D+gUyVtV
zMk9rqUMC/XjRmNVXH2pQzrBR/iO/oUinlcsEZLnNqqZSM8gY0bu7OgqIuwdAa54vC88Rw5Q4ui7
AVwyFRuOPKUJ7iSa2FvBnUdzhNVcr39iMnC4Y4dorAucaiG1WRqr+kRomXWtfF1SAvzc3vTNKc1C
8DY5NSTKW7l3C01selnX8MSxim476abhWYU41VFv9/eSq5ZfswXewFOEk3pFiMtKE6Rol3njCRXs
X9xXQ5U1fYvLYWSGE1++cBNXQqFB8zbb4tUEzFPrw6P5RQjavo9TTNz/NEKb1OYfv68Nfun/Y6A/
s1T05q8bmueRPyndzoTVfTKZJmH2Ac25Q9XFosRmt5wuJ9+Z4hIHY0p9R+svlhkpSPyVH+X72cjC
rRPqu6Y6OmBhwUeeNokjV1dhIvUrP1uOyerwi3xmsppAqu/yKG449iNp+Omwrt9+NlsAaFBNT5uO
nj6aIpbuGBYFLQ9MTmh0H2Dsc0qlsCDIibVGsG0FTbc+6PRqqUCcwul/waz1ZGoOl8VpNDtKt2H8
URrDCb3Z4y0NNGiPZbOPUnG/I1aPx0it1WjciJQxuCjhUETbkTPHo6GMrkxNtddj7Bx3/qY4eoVw
x0KjYv9l5X84c8akKb9sTU5S+vVG02gJUv77Jf4eTGiU61TtFjesEGpk5JDGxJJezGvkSiJPZO4Y
7F3evBTcPnbF5sOOVm5anmdEt5ztxhZp0OUa2VYdVL+40DiaVsrUSCh6TxtAfzdwnonBElDSQJSy
PZ6VZOgIEWbwC/Mt2DWHIRf8keT2HLJ0Og//F/uHUbdaNssMqcQw5NX3j/M1mNaJK8BxO8fLs7To
zPCCo+GXPa5mtpOmKcnvofrxQazc+RbpBRmLDsiAw+U6LG62jrKnY+3EPmN0CqjR72wX5WqkTQtQ
RQFFXfrcxHfpirB7vH5pk1wR5jhxUE6PMsNjA6+pd9BJ1jzk85ljnmSrBs1Azox2gauSh16uZFFP
NtzxrkxyrMlTlyYNDfAtzMbMZDOYOhktbLV4e9Rn8CJptFpdMJj8YMxGzWfbMdXx0pp9sIcvHnvO
O6gD934zw5Wzei0DS8GAWqmSrFqzs8gGSFTNNtnWfxV/i8SF8edMAOLULSFBggv6p2HZaNUZkvRb
Xjpjsda3l6Mg1og8jVecfH4ZNLCz2El6xR8DfJuVn5geceIaxidDhg4YRtUF91Dfy0//4oONoqoP
l1W+j8l+jQW5yX5m2zs7B5JVWN1US8/GslzBq+QrdSZReTkYRkvc84FWJzStkQfmx5rfonqY4ksO
IK9LKmwOLxWqo+76pbzHdwTu9mIUp5gw/qnIUGGtQsPrD29bIYzJf2tkxrrtbj1y398n72NOVOB9
nX0MNGSdbnlMa3qSKCjsiFR8iXlsWiDD48oVN0FeX6NO+/awJRdg7jmCogQumJ7qvol5BedU6TIy
Y84kSP0+81wJpYbpi4RcuHSseAy5dUclOXtR1pXM/SvU2jfejkovq7unfFZK2TZNb1iyil9CHb34
RFF/gAnRpO+OdZHQQjgLOQNOBUZTiIpn8l5ECGGS8TMP4lZu6HdHJ0e5h9t0siGJJUb0jUzAMPqP
aacxGhPSrxZvRrX/OfHbYNZQuqDTpFYVjpDbSLqALKCJHejssLlB583/tjdGojFS1FDiJC+A9mLh
3vNsjK88rV3b+wbKzhqR2SMbKCWzz0uvmutiNQfrW/NpJX6lpEFKkct0ZNvDePQJKP5U5ZOz11Nm
Esmokln67JZbVQXSWBun6dgvM2J5Ncv3X6XQZ/+9CTCmZZzz/z8P1PkYYXrUb7j7pAxiiPBMeYtE
RTB0fCI4SyHQrKt2XdGxhkgVgkcnN1dMefyYO3mkwVwd4Uu6FlEjOCqiCVPplWDReGRQ6utQBU9t
RXsvr8a+aPa83Tz6T9Qp/TDNiiM/esiEuYgiiM1DkjznrQQCeN21S6kkDL/qx5ffkpU6q9cGHYUj
mULIdB5q7eIejwB684hl0bAbNF4Hi59/TeS0wbZdHFgFUzjXJyk/RfFHAFDDvpHUa0Dj49tV8F1L
uoqMqnRVSgEtJeWHAt+ZKsDmjWMfBIVH6LwRzjYaUV8Wjv3W/JzTLwqEBJ9yRpDRdI8vD73/bwtg
/BhywEj0rAtXoCe+ouxgEB0h9HU6HMVpHIVYXOdRiWCgKlIw3tBTz+eJZB/d7jdCOdu2DbbJEJbc
ZiG+U0HZJKwv/A03pozFLYlgX5bylBXGiKX8THyUMOr+vKmTH8xREYZI/PA9Alrkqw1uMF6GtW5u
mcvf8xt+NOTmkrWu5bahCntgMAka/xU9+74NZqrlP/ovTgk2PCrul6psbDoXVT72PtOFukBQjvkM
KYdNUYbIMSPsZfrQJTG3J1CqT50g4gF/dossP0cV1yZpxY4Fei5ZLPouGQs6OerZyxS/wJYeeWTd
6BwkrDbtKRnBA+iS3Wazyqhs9N8POD/oj13M/fSSW4svEzj7w+heIPkKIm0/NPRgxtrf46smrnKK
yUJFPiIVB1rSmnxFVnDLmgtEC6UDcQhJuC+VfzbOY3vk3cUeAT8IBiZoSO3vzSoyz8i+kOKTfL0S
0msA2C5bJdrYchs6vfGAPKfok3se4e9X9gLV8QG5+x8X9Kf4D2WC7jp2/IB0MVZwGVNnLYJwjbQT
Y4OWm6aNX2tjId+BB8hUl3sHDU8AiDA7j0Kv2GTJIvnDQRdDm+/XvOqNn4gcU3IEX13dZdl48Stl
PKiTUAHoQsCIonghPbOlO/n3RZXKYvhZwRnmEL60PEcoWFXLhItj1fjrrfA0kbbMx+TRQ13s4abN
0qfJB4xlECS2xT9C/rnspbK5OraERpKGXXMzsHeyPg0N1Lb7iQvzOGekX63Or90oTxI9R9zKQ7y7
TEjtXK6k/CXGTtAvwZs0R0C6sUAyO21uAhBmecaHBzBy+1Q+w87z6/3L+eEpvHMpOy0wviwkVbIt
Nj2OZUXdYCutSfVsIZ8tws4QjY+5044h8jWrUi+DH1PDHAsafPhQuGnAIQyU/VcWjD+tvDLedXvm
pbObqMS9EKtcWTwFU/B1fAkBJvR+r+oEurcjaXqBbxpsbUfqGQgVHt/jZvcdbuatQw+gJ+6UtTLR
3+JlLGjMjWn+nV5E4MPbD0Vx3HFiJ0ivo/NCcDUqYsp9xCLc/9s8eJfAjuNzIyNedRd/mrFJuHkr
PUj0Ie6GSGqN0SABI7rhOj1fJHXW6sSQB10beroYhQWm/Y+XOnyy2QHLeRfkIbC9gxT65txFfRxB
5nTq6yS9zUwWlwcyYds+HCz5vrkAD3mefLDJiGXZ8ORMzc/M87Ux9gSd4IHuQiRk7RA8tIzCaB9O
60Jxcfz2ZINf8bNyNYmjeoAw7KKHqlprgnFdfmol3khLXtT6ZQW5x5/zsrGu6XzaD7rQCt709cWs
KGoDFNtxZxKqSfFgw2VVqaDjjl3pJj2T5zblS+c7Hf94Si+RkJfnMCHv2BZOC4awlsLHFAtcxgl0
HQLU5bU5u2J/OoT3PqIMoz8e+1FTh+yOih4WBgKRBb1WssOKg6onXRzvUNelZKIgxNs4WZbSbuW0
mkd4nLIupZNd1LU95N15XWNfW9bR4n654kBVGo8lnzALDRHPqCXWuk+5Ogq/gDGfYUSGVgUfaS3u
r27XUMTqyRwSl9M0jWYcCKEIliSfTWfsD1G0KJkFhF10mKCDHHA8jd5aomuCPYMWbK1uG7/O7hBh
ElZjaGdfj12liZ332bw3MfeoJVPXioHBKdOVjt6k0YaUi8/R0rVKl4VF25owEBCgDVb9FA8/VwLv
pie58B5cVv4+IDfOdTJXXBIBC7eTVdxeeQVkyh5LSn8FkbXp5YbAiKq0/8cFLOwgzk0ae/gC0IJX
d4os7zsYLgi+Ial+x+z6KsO/77W+NDJCiL4bhU2NquPIq/kKl3uTOjGLfy6vap3oqhRr7b7/AvS+
LkAAJBClgKRUGzCYuIrxK092pwFCN7TeX8yE64qG7hK83jYda1LAHE4kJl7b65xmSH3IrQ1ax1IY
yxFdK3OdGwnmXUiCKCzkIyFb+C037zb2Yvwp5j/3oU76WFe+6bJc82vjabUhB2DFJMYfTAqY5ON7
YulNaVLWpyBy7bHjmdq2axNpYUJdvSnHPlsBuSqoYNOphC8hTGnv258LXY3Ow29GGVMMa5u0C1do
qbYISqWT00LcYkI1IAvquW22IjQNJMM+govH+xffZz3r+d663YJPWo1oWAjrq2PtEHUsBmMErak0
7VN+TUCYVbr3nJiF8gz9m7VjPbMNMEefrI1vnCX10QhEgJdalSSmKB++s8ptWSLMjmDPNVXy5ELQ
oG2mP2wKGGQ07kBPYekhr2spV34d4qTsHMXTKljsyDHd3rs4ANdA96YZhNftBOBBPOQ+W4XPTMQg
GBC3uedpPWI0xDlt40tVxB+c4H4puVBayf5Pq8Tm3qqWcpxvILS5ZzvRFJfAdDeDfF/3dDKCBGht
QSuIwFOYaxFl4ftdJ3hd2LlVv6DYLUZARXTNC9GINkPyr/4KN6ZVWSNWwjhgT9XAqF/h/9pzWQzK
MeMwSzPIPHMOOFhcA3UR53IJfPPxIsqPvyP0Z6JpBxHbtWLKMNvipbRZR4usMNaMcmu0iAFRNM/v
e2nsrOlTawwPL7QW/+SGKQ7w5cAuuz7VHsvO/2//+M71PReg5HskpKApyRk+6FJcueaH/j6OPyaI
yh+JLmjNQNl/IOeOWZoEiAVTuSy12VKcFK3nSTaiOmMX4YC9DEb/3Hy8oNckZ79SBMN4yPl0ayCP
NEHfny+6Dhapa+QaaW9+IpWVy4DssJxeUiR/2WTAwAmC80+urk+jB2Bx1uY25pb/UE0v6Fhp7K3E
24teifaE5nOM/XoivVi0hmxdlmYncGIUINXsRgRwdb/Dy6rAqWCiDzSJ4tNjPCKKbNzI0bSFTe5w
Wrj7Z/v/O2iIuUVdkPc46zXYYDjmvs4fTzlwJy5l2RlnpPHn1yaRRNsa5o0YQXPExUU07O8VDHJ1
z6o3mkGkWeaz+Qt8I7Fu8XayW7WIufZUKbIW8/Y750jFOT6nQbzlgF3nwv5VsDx2+2gC7EIcN6a/
ViukyUFKuhXkpIlVbSWcMeZ5Headi/DHLk/JTfbbllb24RZjT4hPOK1dTkDgJfBEu6tNUEoil6AA
EyNuTjE/xsIx71h1/JJFsnvI1060rfnsMNd6wASQED/MhTQ6htFyTV14SM/gi2vQOYK4tEdjecMF
XWfaje4dyHtodC5XVgLpwOtU47GFhWIKR8T9pRK7F3JYaG6GPLK5r/xfYjO/ck0hyXiKb53vv7sx
7iRtADQ/Z8LwmkRBmik5ldBIxawp1esG1QHJjSEiNMOgoSB4agZNypcLGng8/kw+mP0FpFTXKpvy
al5AujPtY7nLqO0KQixMINKkA1PcoHufbjMzYcaR2OzLhAVab2bhIWZlbhH/9jB4+oXX0fQqiAvd
flrxsWtZDrROlPmh2DDb2cMCVADdHnwQ0573r9GwKNrFl/KIw/U+3GWWXyTEXclyzxoPGmIGjTFY
QcdzMdRpzxAs9ZVFhTRsj62W11TS0pT4VaCQ0TjOBmizFZemk57/zC0xnKCCDvXMLWUkj4vNxhhT
CGJlRh7fGO74hVnY/05uaLVlSgqY5rFMx7Pt/6yu2oBPwkIf+DBkLUABMoaTiI3Hs/9Qn5AGHj0T
bI+u7maoEbC9DvS/1PE95hgDbDPR5SfiVICdkTuzQhs8DwgkqbJyvKhZH9zbGmuRq6oxjYOmIoWF
5paJY3bb4XY+Jgw1QruJ4/8yOevMOsni3QGQPvDlmQLUI75RKcll7iQ9AwXbMLfEstqJneBiVDFR
kd1oWHZGlC6bOPe/J70h/gSQd5Duo4X14mYfFBmlqoAOuMDn/N16xQepPKFp+PWg784cVZhQaG6t
odEcwbNcWM26mEiA2EllGKHJBTFW41etzPGB8HuWn6MO1VahmScXSibnbKejrKbTfENOFhPxkug2
Nrhhwlsz/+JgywrSengUKTLiAAZhF/hNIRYyp4dvspbSb6xuCPGSV5IFm7+OdUmAPkwjeLOuV0oD
Dsoyy+n43jlpifNQpEPMdGC7jYJVwLZzas6mt7K0ZSs1s7rFh3dEHIxd05/YoGlJ49/zuk5hzJsA
X6u3sFKcYUoEp+8BLMfbBR9fojcdRTvIpoZd1BIoAMsC0GeqzwIMS2fxdQBMP26iWGH61fZada2W
qwLfFVehe2lT0RUDi6efT29c3UKa3i5Apm8/lry3FFXeYXtg2LBQ+0hTxSY1DiTUx883nXBcsXw1
twmVr30ovAKXCq1j7mWS38O9ehrXsNMPkeFORY8FSHDApV1dPktDFYfu6uPQK61a7luz8twRq61W
KEirXZdce5anCDJXZrCYxEb6GdPSGX8jxUvh3CBMli0+0CgDX8knI/fTVyxopvqYth4YgencJnxe
OuHYzHSW1yUBWNMALqmZ3UtG5G/2+J4mSpDSf/E2H0LNMPPLLccmfoYH8Rpg12Pm95LcgeUpzavn
4wvbBpofXcRPwlRe/mV/IR3ewuZiB5sWeuCFxtcg4Hri+Ns/Xwtv5AHdH4fVrl5hML7gYUamh9oL
IR+nOUGbC7UR352Q2lJyua2+cdZ5Cou2PCjJJpBKQ1F41Nlro2Zdl+njmTiQ5RPsuDv8MCAmBNGu
N7jaUod/kq01R+FWVb9DNtH6DOfaRY9EbAJSEjwxbHH+gs+ZoYPkNMI3rtasiEZyWvqq4WHxUXfi
YMcy+efCxo0u6/pWzImYycWdegZYu5skKbD4POpvtOZqdRKRRPD65+X1w1VzJu8TKZv4P8xmZz4g
J9Kpzw1MfZs2FcIxw+/jHH2jUAL8wsZFI1VmRI7FYl/9wDcnNJN7iDSJryK5z7h3OyGXHKxnGrog
n9L1M8mPQylYytswRLW4fW/ZXC1v89exD4h/PCL3VWOnTOrBjxOEWedLc2f4CMdZNupB0gt6Iv1v
6teHf66B1Us1BhzZKNR1hnLGJJgoPBMlxnU9h+IV8RskwzCCT/Dg18W6XxoK/Y7nm2rfwziMF+G1
AIY/TgSLnIkvk7Id6vJSxooLAwUycZiQhCZiHt6j1Jf3bootQ/FaNcLBi0EWc+zWhrL3qOxJ7lpR
Ql0W0o0bEtgOfqlafDX+K9Hq+rzvoToQYuYEqkbjxuqahV7ZWR0bMB7FYyur5PGPlnrc6I9MUZPl
3NR2Zu5D1fuvU5e4f/nHeEXYDNyn0vzTVRyqyIRyhaGOITIjIv6l6opHaWXCfWUsBBGRMaE9gOLv
oXgTpcDcBT8zTYd6GIoe6YhNURv5glfaD+dyGTTpFQT0SO5oBjiyFD72Yo/wjdHmo1mOc9YH7Mtd
TZfObPi04fZhW2xPK5YTX9G00A8KubHZ3UlIO+VIUNPvEU33+wYsF/q5j8zJlRQ4MhhXs5LdxX4u
pIzjFnQc/C6PbreDFMVpNVjyPIHxumtVZqRJg1PQqJOCrYHB0CkahYcrHx3wiqdzPt7ld2o4kWF8
ZtiYO1PEmILMaYqUVeJ9RWQf6l4Sykw2joN7N+mdzr/xTs1B65jS3qqPtP3XntyitBSn0VFWW6HK
mfnQef+yfoBePS0JBwvrXTQZZ1KK+Lof6FgthEsO1T/zlxUbnNeeVp/noBOmBQ74dEbRsHOFOrLp
UTEkYWVgEhaC44Y1XTicp0CzbMGGy7p2HgjAnLwyhPYLQdGqgPjCFXPiYwiWT4SLz5IHlerba9oJ
3StoWqScz0YwqrbrCGhHphp3AHPX3gotxs11yiwcun3tfCwi3QyvvYOQscGgOn0wV4SMbI443Bum
7+s7uZ5iMqPppnNhaYnW5id58dCXoBYozHDp6Solmhvi6blvbgspPxAcjVnG/CMnTbVYiOQoiS+3
syHJuVHg99nv4XoAd3cpEShY0Sj2W6MzgrBsw9xYMUZnu3VVHCiyiWRu85n6Pp9W1tvGytuOTn+c
2Ptbv5R26TSS6uA0PdGo9BoMzozngCzmrJkWTfMv0JdmZWDwyktOt9wW8A+K6y0zqf0M/1p4m6P0
ffq2v0WaVB2vTejC88V10t7kBCZ6/yXHeOyEGi0nz70RJY517uj8qiANhJaZeFFyoGCxzMGpcmvC
IItuKH6qenRb3l0CK3Y7PS7sfZTXEd2yLOQGHjgZ9WyrXEBydjP7F2+vpO0kFp1tFYUl4RxuXMrT
jEe4YBKdAv1ybVC3t189SaT8usK2lexNwDecBIduJH62FnXeOjQSFVNSjzWIWgmbsfqYPaeTI2tc
KQ71SwtDkSZ47bi0+dWo2n8hOUfG3pHVzzSaoFH3DV32SMFNPVb9DM50UHujp8Mjh6e5H7suiZ+Z
2ARkVvS0Qaik9ykjr6k9mnbI8vvtWNMAPtwQ+n6GHlHohjlToaloKKvQVkQcZ+nItqLjyCC8yMxE
uWMRpbMgpe4qIS0FgpEjX5n/nK6hRaWQOXcL5G+ctI4ijpSQ/Z/VuK4tZWlqqyMcr2KON8QVY8e0
t6xx4O+b0NAtdJ47i2GtZMkOul9Hj1ILuIcObumCRJAB7x3BFLnxfpWiY5sWPnq+gW4amKY5yPBG
mf56U3QSpucEnKEtHWTtpBfY88YfeErqjX+zGgmw+5TttfIreuLREQdLkafyncuTcSmsOfhdLgRN
EW+uogbYM9xU6oSp3mnvzMmft8eCwHEA1yg9yJatVGWedPC/KAva/jEDvQTwRuzFmSbORWSO3H/m
yRHNmZl7p2VZsxo9WeFuo4aFX6xsnKQWJI2TWtvS7/sgYRHo6bEOsOV6xqSAszsUUkGwtRIynEwL
heao0R+1HzrbChM70XHN0ct/1HBAV0nKIy7xSv+7xnLzjMBdh78O5b8udiul5INT921TFTJpTwm9
lNth8vNgKjiQU7odBUyJsfPZBi8JuZmDV4CYYFy9oWEwID1g5T3lFLJ2rFeajCRWNjEP/sCllMA0
woKpx/hZaCNvlZ2X3WSmpafd0My0Q0dCqcro4n/Utv0E4BasLEnt7LL0EmEK06ESqUSdrbi+Hbj5
+OuktHPFwf/DDou3Adwg6hOq+JdUCBvC92L2lguW84zFvWDKBwuzDQbFG83nD5uat1rvKGrVc+nS
V3oj5Fba6AK8UKH+3mfC5T6oe9Lll26eya/PJCvE8Ky/qUfVoqh3Bjh0Y/BLSyt3J+esnI0AttrV
1F7Dv8mDzMG37YHgudIFh84IYcv0iT3C5De5lbNSTx0CLUZHvFaNRpcHuzlVr4t5aRIKLYbzTPMG
8AzW6Rh0Ihy87nIZDYIHaePdb8at3WYUuAndzvgM69V47UqzTCa/pfIdj0Stmjf94tf7RTXuAFD0
MrtZZy0FvaQAOperZKmD7uvkfRHQ/w0ggoUxTenblAgpDTwdZJRRLr1LqmwC/jch0AMfc9EgJSpA
Xb1XziDNSfrIaMazNc1bIiF+VD7KiTrzW1Nsr2jRKdxluUuK6PZCh2txgF0eFLM8/i7zFFcyj6Fa
DYclgHwptn9wufnXr4060i1bP5luH9jzQapSDXZTaxQKENyT68e3Kv1h7SJvO/Y5OLfG/vh2oty6
uWLNQyPS5Qmw9E+U6hJRes5VnmtsH8tSVqQ23VUGcbbCi+d6Sp+Snp3fa9zYLG5kXJgYHushOuLr
rjRhRCb6jbDfw30nGQqMhPnU+mUhs21cliR4oblswrPjYHCJ85E3+ojHGD02haRtBrRpOGc/vdU2
7cP3WKEuYDiBr7riVPo4PDCowK5cu/24NnK1r35V/9KJ3UIaq0f8cCjWacD+zjFSGFcesbiZRqr8
feEjasdl/7nBRjBenOsZCdpVqaB8B2BmqNy8uZAun3BQCRKArpm9BzQwugmvM3/BwKqNjV/BZtw/
eLuLTrZX6AEgVEX8Xw1aNL8S+xc44WDLztUKw/IOAwFmqp84qTkF5CftA0H2Tvg5RP7U7V/6vAUv
GidaDiAAoQCq4CXz9gcFsVyt9sMRzLrD4dyoEk8pwEGg72a17Jg0+MjwQSmP+eCGY20eqZDrwkY6
DqZ4XW+GU8RjyzGKlmu5tYx3HGnSdh5tL08Olm12XNbvUyLPq9/0ZYjfb5h4wELYc1jLSz6r/Agc
Gw0tbaSLY5GzF1v7sjXtU0w94JnVfZlVkbvEf1KaL83HksF59DhYw8WlJkrgqolVNZ2qK8QavFvX
JxD5YVFHSrQkeXLVB4AG0ubpZ+MQ93BBWLuKhopy9ZDV4dti2Y+QxsYKbPlAzgvdYfIB7LOycfJc
uCYmgNdh3b7d+Yg8oed7QiI83nR4jA4MYH3vUOmyX072OenDbyYnsj9iN637nR2FZW4VBiS1GbLk
3YjK28TdHiKIsk4mzO2Jgj5QqG+Do24EMj4uLTChh5W/1yAvYypjZQtfoi4a4ems8zhAxZ0Y7gOI
TFaXnU2uCGY/QVSceNLxE0pp2DHJptjdekBviobdFWT4X9dx1hc20MtPNEbQw/VJLdGbMU6iw0P6
7AaoRRqPrZNCzBcw4J0ShTe8xO6haXgaA2tnW9P6nXOKXw3Xiz8T0KIMcCbntqlA2O56hnPHgQGG
KxUIuDtP8QZNQUVJ8lu77xi/kQ1hwQ8PnEPiqoZ1zA2fKGHPiaOElVQF32peMoGrx9GUmGa6iMU2
ygJFtejwGj6217rdUyDZgRvxJT2BBDEzD65gr3Ws6bilweyhIGGRdnYRtAHgOxmJwqzwVK6LbiXJ
k9/KU5O4dS8uj7uhZvBgFwCWaQvCS7xB20iIPIoBFplVdpqtIt1w78bo/Vi4MFjArCIIJd5Q771W
q/LcmQt9PT7VEEX0Pwirz/RrQhfYBeVzfs3CyPy7iRbGV9RjDsxHHizGEHUJ90Nu3E+GNeqADIOw
I75PGAxdZFPhD0jY4xDXhLPVeDykVSCoQZMof35HBBoqTR9RnXrWS90GH6p0/f5kgLNTHhUjmBjD
fRzDLOG+sty4X0iqUJGgSRyKEjCy3LeH266WG5rUYmSVXNxsNAiGDUAdwWdQnNMQ+zkbQ04At8Oh
Tn3hpEyAw3xHBM6kpnCMAo4vv19VYsHHcC4e90e9+U0ci3dtKIUSj+IJG7oKh9os4qEXoPU4hNQ+
YcTjnsGpOPWchvPGZuEyeqa4t5vpvJVcZsWQTjCzQwjmvEd2ni52Bj8MBhhrSkDZB3tSLiPtlTxL
j6TUNDnYlhTv3Ts6n74tA4M15nIH+RcvHp/dXtJxBY9desNO7LliO7b7szDnaYL7bfYI69XwCV+1
usq4G1DLGFF9RVBz4fQdvRodMtNCgnsoSIeCzZq2f2EvraV1QQ6jREQSXsDzMlUsQgmjxwmc9ZNd
Awc98p5AbVOOXQcKXCU9tTEXLAUd02aa0C5KHO3GeJ6WoafSt2sjLuferd540nrbnxIPP607HKru
b3e81wMDY1XnGgDi1hCtMtN38DMBBMhMtBgZ/XY+GEOdnOWA3fr0sgFDRK/c0Vu0SKqdm6ZnRQZq
ATOcBKiB+Lp9pYxZQ/i4Q3zEBrhbw7P7OBtuSfqnbmZt+kfHaMMIMdD9FLX38jj7nqwPM6uFUXzd
d3dZhNFjwen9BEt/lD1lzpcyfKm+V9QTvfNEikHvvQxQ+tttTQoauwGdpKEzOreiGt/p8ixSg9u1
DPAGI+D9vfBwqf/lcCP5H2GGBTwS1lSNYbjpruliMhynHKDN4RryY1Y7sPZ0oBPFvlW7GwuG+oAX
4LSYK1sK8QnuZ2fm7pjpvbe27v47S8engwcobGcUUtRb7+i6QE5w15q6t5Uqi33TMgvfuhnCyKAR
wUWUyxWMAbkBPp3QbYJ7IC8J+9u53RvmAlMoKvnbDtWYjmNYmB/VriprmZy8jrB7K28RPR1tI3Ww
RE5a6K5I2WNZlIykAOzzwDpSMoN+Hg0Fr1W//15f12Bv8XJwwVseRhL2I3pc30bLFhVGap9XP1YD
E7hbSbtmdeuhLnkhCobotd71lWqs0qZfNMn+Wfjjq++gEPUxmYh93MK7tDtWB1XuHYXfSvsshvHG
RXoxXjbf0zpBEeuJvjy6FYiyadTh7R9exQGwuSsgnuq+YLxPhEJPwR8xwn9lgSX8+ztTF1QjpLQT
/vWKklk8tEH4uQ/4TQI0pRVIXF8PF+LehsAM8+eZ7My6WYl+zC6c74uFlSvREHnK+m6AfS6dz2eo
eDGWzaXmL8qjM6IGxCsrjnft3yplJISww+iEjan4Z2UXQEcRHcERuHmNPqel6bj19LPBszYH2fkT
xPQ75nHiPh4QPzweE9snmUqaF1kUvLDvzodV0XqtGe9qk0Gbr+tSdjOgqPcaoI3Z5G7pEgfgmvJK
/2ktrGFlNek2N0A0ZLPjMd5KINbbKDOLznGKIqVX1C4qNRiM6sMDtagYYjuHxi3YETIqjOtThirq
lMF89ln44r/Hbm/n7xmkvcVSNFbJmj0KfeH42ythsou+DmoZD2fIbbv1i0N8WJlfRbWxrQVVRhpV
KOmiTEyT3LP3v3MuiBNJ/ZevHPH3IgLwlBj/AEYIr9w3aGDGkcpnCYKaCGKZ4QqZqwIxvT7ghX9t
8NjIg6r7QA31/MTWjf0JHZqymu8je73r3AO7RimL3q3s6+EOQveO9iWVJ4r39B5uXO9QknG/8W8r
yEHZeBBXhIWspuf2ByV7Bx/m/7isV29oFoWB8qb2HCpLaS18vI1eIvA+8zYFYRHDAyp31oTSgXCZ
J8CgcRFbjTIFrYZHBhTw67nQv0cUbIordxEckK9zKMEpY98zRsirun4Jh8RJ/FLz024OuMaWbueV
yyCa2vv4/YRosgnw7llnNL2sxZdnVS+RjtIgrcVNzcH7CFoJR4AF02xvhpaXj89YFQ8tWO1yg/nP
+7hpjV+ri4iRgCtj3Wwily4+Nz+J2TpiD9zPti+PRN2kb3I2IcvNpimnzGRiPKrOGPCZwaueFxT5
puIaDpodGjq0AHf9o6FLB9euX4q9eTP8j3VaQuwff/FbzeOXeW5Iw/Vx4M6d4Xr2laQ5jo33BFza
cWV6Wu7YmAkvkB4uBmZCYl1iOm8xNbEWR+abblq6746Ke/DGHgoWv9gi4Psji3srYnTPOEBaU9Dc
x6ZbM9uNJ3qK2HPzKV+QseJEuH9tztUFSIkz/slllrckJraVVOBsohdTP+BJxgVE/197Zqc5UvWO
zh7yAJXF9e+DS9HYTM1szHUiyJPns1Af+HMH5qyp6kux+UvTZO85w8XybpkIDvp3/ALDLF7im7hJ
Yk8Q+bdeAZj1WysItqO3d4SZXMqA7WrXZZ6FWLN0ZEywbeIhHFT322x8p/GXEf2BwxHZtIbss4uI
QAT5/HlNQQkHkK3nYdRYOg9KD3jz0FfQzCaxB2CRcJByJi27EcL/9VOTGfRmgfQEP+4eXht7CNG0
tXglXPl9KH+WEhUoxhP4ZoSDT5vavgSn/Wen1We9g+DKz3N6z9VJjtaEQine2vLm96u096Wspvir
zcgj04iBzkwWNIMUl7YxrGujZJ0GVPQ1GzkpfBK8CFSYHWQi5mJ6SeiFYbf4qrYUOLCvxTUpJjrx
2QvqmxrQp7TzQQcaxnvK7GJ0n4/RveUd9ICkDTcaWB3+jY+PViv4gFD+rwsiLa6RA65HgQTD+x9p
vmI7BL1xy2VAzpxSPw4x2hrWQLoW2Kyuw0thtb1yi/KECXmfc1T+O2LUKZF3E2/jvz33HNgFfYMG
SmK1rrULQHTbz89DGJT0hcmPLgrOaBbETxNjegkCu9eF0Nm35PPYggG/rYl2X0Tiykfb84mMQ/WU
awLymnptxrHBpLcuX3dYHeWLxrqth7x4de3MuWcH2JdRTcy1Lo07VJXB7IYwvxibj7eeSfcfyMTL
dcoYdFQOTBdE7X84VYu6o3YJC62jAIi5YOkb7AbwZ4cvWCSIxwSDeycYUWWZXobmb3CZ2JTk46BU
DluMeuHKaTyoAGvQKC6AcIHmwFRUgkPcwKiCRmBWL+n/YEPnmoI6uFm4i2EsmW4up+RM59lBvCHf
WM1410M2NEQoqJGyVD870A2ErQ3VefSwlsxsOGL0Uy3NLikEKFflgCKBoytU4sKRoBMsi2EzXmcd
Qwqqb4m1iMiUx7qN6Shy+P8v5vZ+xqRcr+QGa7SxyxXgfVr66tKjHWK9okyvIQb8Pej9qB4yTyxJ
oCzgDqczYtb7O4v2BbdYgVwruKJkNwNLwpAlggs9dEppU0lvGk9V94wbJxXW7pVXZtRICP9BC8SS
4stKYqe7GjkNbwazZlRVZzhdOLOUu1uuM8mcmsmajsrXu9Ioglc4uGLgwFyGSDSyV6U8vjmucup/
eERT8wxQCPhH2g1GTOpLZntWTlcmadKbg/h3IVeii0VVJzC/EvxLX9XwZXt0YrTfoHZmIONDowOx
iLkfS1h3E/b1W6O9vsi5zeSLGsPSq1CxUKyVCC/n8iVB/T+mecc5IBX1vk1HlzO2lWh9Bdv0mmuV
f1JljAzMU8n6/JzZHa7OCiyZM/vmq6LQoAdwpN7xXP/yZ7uairDZxdZvdELce4E7rp2OdDDOyBaS
nZN1OgofmCWSbPXxit7/3m1wKgmF0Inu/zmWZW/OPv9JoCrAOxQtRU3yzm6OUNb/B6FNW9KMwo/p
ITxJPo9YcDLfWYYzpI0sMdm/YESuswu8kjEm0RKJaXmvcGV976/26WHpsu+P6qbHcmDamAW+HV4d
Npog+CKZL410UoPk4G86xramWpZBI0xBHWMnQMg8mBCExve/FPeRa6srDU0CWaBHp9D5xwihCQZd
LaSFmLPldiG3wXt4od4rQ4RECXlh9nDJs5UhDdVMqorM3IHMTaHy+PqY3HSPW9IMA/2qUk3UUdrI
3u8ZySnggZJLtH2xeF+8/+3isHvNXGgBA7u4jhvzJ67vjEMdP5wYeJ1GyCb+EqYZGystTUkDN5hI
NYTQ7l9PWVg/cb88MVn864nMjWUzl8f3B2Q3kZzE4S+Tw+3ld+FxVMcz1qKfZed2uepuxl7wmdlp
x/5a3sVTnIfaZFInKsnW3jYS8971cLK2nS8QeqrzyP0GushFjcHqy8CDAIxfYM312J6Zmc2Pf+Dm
T7V/iZ4tQODIUDXm0Mlpmw3AS87t/61CtHVfp1tTqfp+TH7BbJA4IvqXKkPtnABdsQEH0KGpaEQu
s3+tVF/M3SUgG21vwyGtY17GxNRAb4DtU+bewHoSlwawriFquYjksYMIcYLVCVz3EdFZMWkyEdYa
pquZJAZFJajK9KLiSQhFceorNAkY8xi9iYoInZqN3DoWcoxi3qQZlYBzUMSLpsLExnbBq9dI+Kwe
bdBhFUSqSIsJsp3RUQCTVDxL8T/uXYV7++RDXOx1Xu9LsL9qPDEVzaEA8Zz59ndIcpXuUIYl76pZ
xUxLQsDBRBJjHn2VYE+2wjxwCHSpSmWCmVuI6vS4NS616aV9UEKKQhApqNjdMCT8JpS23Dq/Gkq7
v8jeNeQZsUP64uVUbLwYrMTGKe7jOMAXtEadFd3GtNOJsW2AmW92IoxxrE31Oys8qcCVDOQwKSDk
vJFB7VfVCInW1Y8oDwXvPOjsdwvw3zObrP5Nl1oEazleCVMbKjNKBBRxnS8ytFN3M7S0uqq+nb9N
UrfPrAcwvS5dLwXmZhlVbl8xPFxuCvAvxfE6IfkoHqfdXU2yMG/4zO6lD4E9T3/hYA6UKZyT18gE
mr44OMC57QbooDC4kwszLP454qUKZ2TsBcrkJaYhqaWdMzJXRihYh04wf8NasB2IS1cMcD5HkWSQ
79ZW8FBSbo+emD5cd+U+GnPCggSIfqfCHOhQk7FHfCoZGo9nOPbTsdrlFzL2tgZ1cVg4OBZiLzvQ
61Cv5Z6LRTjDEJnsndqbSUWt+eQNI9np7gRJIQG/HGXkMYvLsI+0YV351RttFCye3YG5+ogU/dWr
RLzLN/6aYqc4bGPgbbuRAqRgsWunu3L9j7KrWE+uz1VZOoz3eWol2QSwjEhJR1OkIWwkvHgva7wH
wMdYVGszanVoytcrIKmSJIWh3QPo9vqqLc4Ae5iYkumRaQB4GcXcAOlx2mhIp5Zt+UNU1RfCWfve
aVH5pEZXl1RxYWhFlujPxw9p2JVcjCBAotBOxvGjp/ECGvisoXenrjp6tq0MBhIZEPh4ZozH853q
jSSQjEUnaLoCWAjBUhWH5wGhiAcf1zH9WY+KTcM/1aDiupx/IBczjotZmu1AhWaAJA0e+Cz2fQd5
b+YojouXYOxKivYvidRnf6rr5J8+6GO903SCfUbo+4bZgzOQhZ+H6f0FuatXmD4Y4dns6GmEiqnP
LnhWCeymDaigLbglbupiqMWJkxipHnXKIAcrvjaZhsYxEZqg+PzH5ZoeIvkblNOqblfhsrC0Vt/t
zPsAhiV7aruSzPer8SRz9D3GUvIe/5/GavBbRLchUAbA0jIUJwBO2ax77ywgfJPAUExo+2RyJSyS
RPLZsEIahHyuKaRoibErUtYUugaGZUegk32ZlPONZW5Mnn83yhUNBIWRfiOgsHumbbeMd1u1MWe/
ZfhnNrrSfhEJVbEUSeRi7c4550XZogjeSHIRNUTbs+Hl7DqNL4VJkvh0+lN8REZM37Muh3tWeo9A
Yje8v08zqaxNhrajscTCN5uQvM8wgAfGwzXnh2X93fuDNA2s7W52fYv3vVYr5Fud6XeyD/ZigZtw
wM48FnOQKdxmiL4VTYJ2mNh0kIl+RahG+iGXrdpM64yVw3cILiJ65l2g8/FQRaoMhaOfN0rpcRZF
aSY37FSyJxHh4asFUGvL15NYyk5/Vp/oVJPQvhV6NfA6SwPVMdF5dfuIhX7IbcAm2CfVGUI+m+jY
Z5h3ncunQ8F9J/Gun1shEy5Wxvab3Wd+N1e8n1maUbpkkojC8oK65ujlafbVIwcn54Ecxz8L+pZw
4Iho9O9d4EQNrZ8umAC3R82nNJ79G2QwcmbNj4h/BBBlR0YxmIoaJlhbxWr5QRE/JH1D0ZpQvTAN
wF1ib3TCNEzZEE8VmJjjzQX1T68XBLZZawgQIvVyjkzQC9LiX6ufxiKpuAkrxbliFyflmyQoOnW1
Fy7JKEEFmUjfgIbbUorJFE24AZjcdboZoccaatG1NLRK0iaXgXG9yAskGnFY2OwWRQCiOBEcKvOh
Z+ZGP7EY28dXmlSI/3Xc3jpCrUFLHcKKjZZTdQOVlO92p6M1ZUdaKFDmtHLb1C5o3wMgaHY1iyOu
byoonUrhL1q+aB4pgMypopqVekvzUbw5Ddq7h9i/p9Z1gvJqyvfn9mHjMdv8jc9sKKrB6KQoIdw7
KAWwyRQUUn+ETqyeRkxSP1rxkaCNEu7hR+EAvyZErzVsbGr9UNPkr95cVEM0V3Gt6f0Un0G0am0d
nS3i0GlLeOoGVmO2I1nWMIwkVYREJE637DMh64hd/Vufs6b/LLrj3x8ihgHlPXnTXprl4L+CQfan
JTYPMJT3i7tzziPA/tyNs3w+BqlMnMhV0qy7JPPTNEcGGJykVvmVi3ZGLzcz+EooGDy0bauCOMsg
zaPYqQEnMt3jt/tKlxkNtoL9225tXeoqHND/yrBniO/Z3Aa8jq70zc6NAS4MaWC33DE1Fgs2/Nzh
EeGvTTy/827orN3lfTDR3jjyCzcTlWy/P2PyGfmciKZ8GgNMfcC8bpsZcgF4ZI+qizdPQPbdh5xL
2ljr0n/Wnc1xcRKVKq4HR4ss/I3OMOiCiBjArUqiRoL6Xz7rtROrg365u8NPnjXbonpe+2NGsGbv
8reTETS1N8V7qBgUC/hOIg/nIoCfeU6vYOTn36fNHdY+uX79vZgw8JD8czT9lMhOYnlwqmPC9Km0
qKYEqQg8Izt81XMF2duFx5OF4Up5iPdENiWzLnZiYnzm1XJBce/87cI5sbrXwZFUDl9Q3kVopkI3
tcCsxGJVayA0T/R5tYVqOOGWs1L2zVD0TAbvV8DBRBU98nQW6WzW0hTEZ+q+8lsIfBevu9lD0RwH
jV8wir6w3XmpGhfNaP+dTGfAEKtBqto7edMefIG62ZASzWKiyrg7x24q8wLZYYDF3+BGXLG67nmb
lojYBC4Uiwv5HNSvSGb49PgO3enDoWYGR/Lr/QbFxd1kvP9xBSeejOoeZb6cCmcRCgb1GVuorpph
F+mvM1siZy0OYEA7DC2fxcw6ZJTOnpOJuBaFCevk56gLT3eHhqAYpckIga9AUuOKEMPc6/8PjBwE
HtVH+muNJvuruOOPO1T1MWGFHyVB8tZYHm1dQbKLZOSo1xNp5mfHi4eV4PbUuQrisD6GRB39+tVc
odnpoMtd3PuD08rLSNnEiKiOSRpPtPzB8NwiV8Pb8x85BDiK6CMs7ibgkM2KRQLkSqEnl4jgmhBr
tnCbzgGxen07axBTtWS9HeB/fkM4Z/l6qBB2WQ6RvihFjwGjlhsaMr1RNQql+k0xDzfxGo/RWl1j
YLX452ij8G+K8zmu4VMBSBa5X4Pved+2V3GgeQj26QeZOm98ALSDzNfFrYioarmYijxlkk0W6WsK
Dx1of6szvLFTLZOQnvuLqoGEA0Q2SeiUuF7j7Yl4hlnVMmy0hUo1u6q1ZHhLSANWlNXC+JW0AgmS
KFXjtbsRVexTa7TVqKtZGv17EGOsbicTGEznCtBTZ4OALW4rgFWP8OEVAPSMWyg7r7jy8NbldvKr
msYreaZJT/BgttwafKbeuqK0h5zAKhhPrZcjAz2p+mQ8WE/SuOblKvoarltj9SOIy21a/N7VZegj
cv5wHW3f6c5HCpZt6tryYVCR7zfBCvE5MZHEkK7RgP1Yu9eV7p5yt2uL/K71MYodGsjeqRLWpduK
e/CsfHiNoP+ET9pdm4nxz9UBlnTq9W3Pyqbbjq7oGWDtcCqlcBwrzgkefEyly+b7vPSJqlN8KSy3
5lv2VCU2EHKfX4FUVrFnNyGLO5RFYa38FPRBe9CaiBRhJjyjaGsDMCSoigrKsbaK4dbyp/mmOwA5
emrJGVFeVG5/GZzHzTPWwZiAt45E26gqICHJi47LL0TfXUyQO5LurbcNnc2ZS3BN4u1Hy7d0VF6J
TbxHTFDeZjYhKu2khke4mYyJSL0eWZuThBnQ5TNzX6BylAQhSoUnBbVg1q1/rfY6A6ACSga9tzZN
ylz0xfYsRx/e6QlNbNStE8qvOcWF7NXGnus9L/VEG1ONd4FFylSeuxKlUT/aqQACMkh/3Pug97ei
wFvhAkhAjN7NX6WvL5lFeLSdpn2WBmoIdlipCLBrxfrtLkFwrgjJMxZGjWyEvM5h/cIKSSZvXyLF
8yYPGuwoZuO0EBFNFpJJd+S1TzXIMyUX0Yy//GBy13RI+pvhTJ55ykeKKSS9YJ2cedrP/30oCa7I
JdhyWTXBG1plYbNOJvya68yfBlcH1qDNozsDxyd+tlbu3YOW7cOKPpF5VW8rIIS4MVCvsi1Li3hW
OiODK3aygobM9ANtC8hCg0jTqxFxDl4x+8P6rlS/zy3mypxO3uk208lCFow9neKbcNfB07cb+I/P
da4wVpoHWlVfSSyVvvaEVO1L+WXcks2ele8IB4v7RK0i5vlGUORtAg8sdtq/51n4oOsZxCPiVISF
zI+NsDrUSXq3SGDanj3lAOYHk9Kpyla1SLkfv/bE8SwM7cA6IYdsIbTza9PyeKeGowEzY6l1iymx
JGELGtafRxgyrFnOO8cpyGDBdDDzFaODqX+rXzjUIB6BvbC80WWGFSVS0s20brhjPIim+9YQhkfm
gI1My1+ES+4ZufKbhxJIeLtsxm2Pmc+Op2KsC5HNxK2R1UJqjA9FqlodpMlxpXMQUjd0r9x9zUZR
ui0DKSCtpg0XAH22Xhgr95WhVTKpXDdouOHNhkIL0Puz98Ol8ZE/youMJiz5jHPM5+p8qQXbtsWy
WnJDsD/QVGiulek/jZ999MWjHRM58rkhWp3kNNWQ/IGXabtmQ0POBy5598cnyX1QiC6zJ3uiL/EO
wEGszVRo5zDkZFs49tyQC8vmST60SfpRlsGSqpqCgKP2pDlx+VdiwYFh+xScsluUq40DS/7I0+z3
2eUTSU2gBqbG0Nl1LWh3/KxtSUZaeEOeP71C9MKF1YgKnEPr1TpgbcE2b6jMgcn2u9tLzSyk90sH
IJjm3rIgsYv/rLltaYdB/WqEPZVvWd2bwbleUwDNBJTyz+pJbuPf9ei7eeBiOFC4tLtl7palDTeE
q0ULqyjsAlfRGMqsvNsMTw+5fjTFFB3uh93JLK9Vc+T5tsE3igC0WWvIfyKrNi8LSDsOfHMiAcDm
bFrGsYCkM5+KFFu2AxslBnDXrn4T6gKZdAvvzksRicGGfc7FA78qk8ja8Do4PQGZobV+H4lpb5LA
lAC5oAQJZLBfjD5uiHsZq/cX9JtErIcgx8x0fP0lzAkuWpVjdzixT7NAm+JcdKgE5zEjzURejBZE
Lawqo6Zrx6T58kugOtnPdQ7n3ng/7G2q4UZwjUrycPOACMTUO7RyGq+9zuxQLu2xoIzuEma3PM1B
6MGEswTJo0ZBl0l1W4EHt9AVMKaDC9xNBRym5e+5LTwupXVGQQ6XGkWD1neeR4jbC/8cWekMHtjA
BZlRa5nlGhHgZc9os+s4GXstc2Pm+ZHRKjrVCo7UNDeRVheJkPbE8i6m+yNZsRe8H9UXyN/9GJ5X
6OPmPK8yB406vPirr3xB5FVNSWi2tbTjuL+4ll5/hBMCQjLHF99E5RMDZpJQYq7M+zCVBtHb9wne
JWP+IiNbwJ21vhAEh1Zt3XH0it7wEN9IIvDMpnE3LSLJVNkOhhhzmtJ8KbSLSZw1VGf3fGfZRNFA
+a3Zgfhd2/gsF/rM+Q8yMeL9RNwvpPWdY4J36ZylDly/8CE03tH/tq9bp1YnUGXaC+Ai9qQ2KGrw
UZHJY2TOD9TmC8L/gItvo2e7IxcXF2aAtIL5RjM68n6OQ0TicDrUhafmIBwAK0hBPLKYJdREkdzd
YT60Wti0Z+AhenY1pQWudCbEhFRczI6pjRyPEEufOo/fAkS6uCL76FOCMXc+8WzvUaY403XsMpcM
JtuAgOGHmYAduIpp9pCn0sOLCOdmkmP9pux+Pd3qcwA918uYXmgcgek2sbxv6ZUjq22WpFdzAM8Q
JiI87IvFveco1RSow8KtWfK49x6fFZQHhTCZRzDzOZ8qjrTWW3bN5mbVoVIxmWzxwsb+Oi1UeFvh
MCwKIpQghXouYjrA+PGEUTKocciQ6M1GpT72EMDfTGS0CQ78v0/B9IbdXHYQP8wbx9vlKtJeXTC3
XFk7DvKHSYg8J42OBmn38pXQjq2vG2M2MIjxdt2v7EGsENs5oAs4SctkbEol/7/ineadWEB+l3vN
6pU50IJCbGdrx0zTPk996jHSDTxK4KZzb8YFxodyfqFrdLABnUk9t6aR3Fq36NucyTQpmpN2wwit
Vf19YjvKHyV3L5AmlJEj2uL5yhRllRFMkg+CSiTn09Qp7KiBwhkEj6mvoqAGzf/zoQnF+5JXpcMn
GU+jgiVO8PWSkY6JdkmFpwQxUvm1hZffQpoyf5H+TfYgQ4S7KrsbFVCWnwi0JNU2DaW4ZxX+KHtH
5FT+2SCSlNIK5p4ZMpefw04FASMeTTJbnmLJI1BC0KQFUx+AqWy4hlA912x8WoAOuKYhPo3oLU1z
UUs8pFZQ2vt3vrxXsNQjPwMwkh7H81vyxVcobWCxlZmSbLOuUkfSuioZjBnWUqk+07yswYExfxGg
kHjd+uQBHKf76Ma7Bsx+XLShDOUsjwstmvSKE2UI9V/G6cMAyif0+4b8pBzDUPYiWqynn7H/YlIy
JIhtW3uCrApcsAIr5y4T0sZnwxnuXGLuzAtBu6OJ7f/U12nA1E1EkPB5SnlbuXkr26wei8wMB6sJ
NJ4QHSeaQtTcrsssmMcFZrTexsG/3czh9RGB6xWGdVnlEB64tYEQ1IrhaAsD5bcQxObO2KGq01bD
pSLLkxEFkw34+QWr33vXviqeDhzlHPgQx5i53/QzMNoKbVzrfiaBCF2pDw7TkG1gGv6DVrsdTBRI
mjh10FgBHtJceahPkjo0FhVjMkCWxudCVdfp3HG+5EZqo7sseWDaxWIyvhTMvNbfqeeFCYDe98sD
y1XIFYAf3L9yz87noTQbntiPnyfvayhJOJ9GsbepgK3eBgAO7ef/vxa2Hnb4pOczuOvwbrpomlqO
w2LgLj30at4v8g23/5mqeKr1Xo/Sz/gQh89j01GoUe5DCImJcfh1UukEpg9AQNvNyWc+HKAmkV1R
S5MFZTk58Bt+EW7qeLH8Kwovpx0AXa8LtE7BZv+n9rvin1H1Ut8tpfwPB28PgHFbOBIQMh92gG0g
8K74syICfAVy0inx3PAZ3F5bZImR3xAKhUYisBOnUQiNZiARpOaZvTeRHeZ/1TQeJdCgHwMOm8BS
SRIOv0XNyB4Hdtj0+aC1Gw7VoAvVeK2tZzeFX3xQ5Ik6Xmdf6N6gOsI/VuU7gESM5a2FPx4sdZln
BNU3Q4nxybjZYLgQOezJy7OorKI1EQMY/8EZ3SkW+9Qxu96PDv4cC+wDe8CA54G09ec5jTOdYeKq
FGSBPF/GBSr+Ak6lXALp3L/6ciBHs8P6VwXHEaOGY6Li/h7wJngJuC8MwsU75GVo9FCDqmKZU6r4
PZSupyEX1KFbBbdBe8hZF8AUwyVr+nHg8K9GsC8dHOgUiB2oChWgc0gbBcMLZdyQXWQ6psdabwyK
awf+E2DAmy+fLsXIDM+y6eiMdwF8UgzUsCYj7pppoEn5NZhT23pXpCfl9987ip3gocM4cR9MoqQ4
aRAI3Nq3aGToHZa0XuNeXC2uAloCxuAW50LkQFgqaU06qKMSxJLkwE0vjFJ/sF/Qnjtbw5oQPvZg
HpYqr7rOlAPfeM+nLeyDjr0c4n7GfFhfFuq8nC957pUC/FV6Ut59S6SXGmZAq1phG+yW6+jLH1R1
QQ1awR6L9zQA+HjAJVWhZQ+fgf8pTWOrzFa8n0RTdz9MI5m3sLWsOY0LOnKUK/YDNUDtAuAZLAc0
i+GUmF5L0vKOJ3SXNVuwif/As5eXkanuldEOEIzFzrOTrCiY+9HR8dAnsixSZnfC8Qt2wwCqr/Di
Hj7A69OUEZpTLIt+8RYMWUfHMjR2QQAazfEQ2DRM0jRJ8+exewc5J6ghq5G9urFFcqEr0E2ByPI9
jsUTbqS7rjaWdEUMicINBaQBj4P6Zf3sO838XSfP8htijACw4+IkeLAAOrMNoyiVnwTl0VJEhZZ4
6QLSdMWabOBjcHhdXBYOefpKmSGB0zG4Gr9QaWx8yLXxWairPmuCIwEhQhdEJbigxC6TCISr8y5B
RqOV/QoOKSB/+j7ekyc81uRrCI5CdT9r/px9esAFaX/UNznnHwh1PLMAqiXruvp6PK7av2Kq/Nbr
/IFwOg1BhTXdIsBYzfl+zPvQMvN9BRWENgHF+S58oXB2Xnizhr85y+Whnywmgpv52/rn1wkIKzMG
3O3W7LHAdcFCtZPtopva51s/FM3p6RO+0ZB2EZXJfmqKvR1wVPxPn44aCbz90PGA2+sHLmKhAfZP
pT+kf856W00WHh6shWwV6wc4e5lXFh8zUqNzgAWlHaiEw5O8uUEZGOYH1DCA+szz6MlJZZOiX7Ep
0zZ7MVlt4Cj2/zJljsY1ihMORsuU7Y5hol2TqIVmCr9/xntGTXxW/V6JRfJFnp7la+34eCQbHnQ/
BkfzNALQn4Yj/C1UMu6a9xNnDa3K83d426mi9GBmcpZBYiL/Jib6BG+yJtieIsrtDp7wk2/gdNHL
dqdQmPNjzDxnKT/ffgRXcxazJ373yIQfNXqUZbXj9sGdpeuAZw0942S6misLLD9WCW8HNRXP++1f
Xsbf1AFxc4LyZLFDxiYrH5yEsPQC6n/BspilGPEe1fY6XNsPNUQyeZ7VLlMjtAwBgfVE6czp6U+F
FM2WKopk5TTyjrO6YshUPn9Ddf2ZYiaj613i20Di5IHGP1ANzqr384piEfmlE94OlCAlf1Yih3Vk
9CpDwWfsFZn+BAAQj1v4IxrlpHa7e91C9K5nrDIO5QkCBXKxDpxqaVa58s2cp4o93NtUY2F8cAJX
mc9NpkFozSYgkGho1UVDWcxq5OOX6Rd4uHT8oEUVnNn+FniW4cB7BW++qEgJkKSB3hD9Js5/86Ey
M5mVzIXGbyGc6wYNGac4xJHORYP2YCzQPFEW2uPno/eoFBOa4AZ2ds8oOHzJHHOdcL97qGiabeL2
Qgrnk4i0YR4RYgl/VGe20tE9bj57Vmrjayr1XrJ0TETCLHsgdXabwgSjZ/ur3kbcTrTsUcrCu8r3
XAgVxU9ahSGRZzMzIQ51lo0CCTRP2Xxgg7usREg84meAeb8kbwx4lp3mb+uAQqJo7VUjKcGKp0I4
Im4r/lPCHlxU+LnLH/PubcRQVylLwmhdeKW8EU/Z5ehJ8I/mLp/lRCcsKuVIYaU1OVq5PAxoWzJa
Ql0hupOc/451KCj5CXg6Z1+Gtjf4gaQIWcT7mrXOnksj3fnNacxVCMY4bfYaoICpjI4XUllJ65j5
OHroeVxmVXraiQCxB0+7u42BQta5uvGTWJ8AbZQ2aquvo+LjGwtzBR7DVkrmrhrp0wfkwmTsZuOc
AhJEJKp6Q9p+0ekuOm8EvYr4LJfPMtdWoSdslMwyg6epxyzRm0sdRB/jUP0Vg096TcLcyqw1n8DH
KVWv2peaWkfiLvzQvhWpi9AfvO7x3UEORVDAqTHQig7DiUVxqs+Lg/V8M08cspUwGXeD74S/YqOl
lNIE6/xexh8lb4MrV3paSzwlhVwwZM/zT0qqvclyZJkMzm3ZaAEefZRKlWiiC49i7vICm3h1Dm5m
/HgqCVr5CXHiARtD7VR/0AczQYO2FpnJaJcr3DqSYv+eD0U2j/5RBwlR1AepaV3YTXfP1wX0X+TT
1QGo79vp1I4jODLTFdvzPsYm6BLfBowWGiUADx10c8KjBeCLM3LPew7cXi8SNezwxhhLbRFx3GsH
g6XCK7WCrM4wW/8mOhvC6EIPh/hG0FqUKThlo4u05TT9BSD3hkz4QgNrazP5vZDOASS/2Gn3vi5n
T7ujSGZjoJr9nNb6OJlVph8cZGoVEir8HgmB7EBVsc7XEIZ8XMCnGgfjaCKMF4hNshvYApRndmLs
sU42IzB4gV3Sj767j2BDZK1qVw8JrqdM9bYb335ZZPDij3uYu1SzmxoDqW/bDRvi4eDlHMTdNQ1s
k+dRkGlavkieC8Cvx8mkhTeYXhzyv5DbzMUhJhb4f9cSD6tOcgkeToo4dDdfEe01fZNIaMiGRvNw
Aoxi3jn8ebmc1FDEeHH4PZ1BYb5n2Kbtmo8gejvLqAVDzD/NKpIv30IDb6ps/MuKHVk6hLfUhEWR
6Rf/pOj50FUUEhvlYFg5uAC37JNo/eaaJOiIFOvD0gh3+CzdXxY/90wf/EF+zDDZEUyu0srIHkSK
L/BjCbTJzudQT1lEvUyk//moK4Z7fweIf/P8rVEMWMftH2+IS+NFHOW5btrxyY8v/CN4iwS9JX+q
JfqS71ScregokLKP38BjSMXI7fYrKJt98AA8jSD7YcjxqA+5F/knRNdQFDHmm7y6Hq07KkSzRzdk
dWnEJzIZmqd/ueAyPSBIsE23N6zJfZp7a6x3SZ+2FTFMCOEzAayN0DuGXkC27BU6kFLkgLnk8czK
jt0F+s1nVlj+nprsf8Q54i/IZS4IPKBUUTYWo2PLdwJYDQOpIjDR30zrLOtIdbFFkGVMG6cwYSrq
jWUlHUp9aoC2AcPK5TCRgRtBRnRMIu4sqDj4zpaXCqF16zPvYSrZuIjelLuG059cVQNBBl3oHHSy
KorQ+ZwoOjiR82ariAn2/1DvhOZ0dcZCN4QY8PXKJWv8PAklgzz5bKp0ZC7eck7V++Mx2z7WRQa1
fvMF084Uc7egzbVla1OjDbtB3zDiwvLYTNimxI9MG1CjF7W4wXkxYpzBnYe1OvtSbScU9bKdkvjS
J7+FWQ3vSeHnSBF2PIO9P+ydUK2jTvHZQ4gye1ZV+ArRDbRg2AAg2YrlhGYMY1mTUgbkeEks4Im4
OslUBhl4ljngwCM9HFJ3T2fCjqWI6n23RJ2+MWB593TEXIa3AI3Q+JLZoCe0aGx/E7/FH5lVB/UK
KdEC3z1HDQmmJHcjelpFmNUIcBAJ06xIqIU9ZK7SSbdebufl/dgHYZWit+uJ2XaZW+EtY2aTgGGO
q/QMxGFU59wSzx0JdIOPpYjiH3wloBv9UBwR3HeKXUW/HypZyBCmc3TM1OcyHATU4Jr/QLboMlSv
IbDhTMrlMup17o0TJZoJGE8cscxvFPKOPNYD5l729jkAZHF7BqDPsut8/fmgJuo93pxlc9n4mCzH
tZGG2GI6b+XwZg107ykgivpp0ebrQabUoNC1AGgWwLq8lRPqU10vhdRKKHzKvrUuN9k26grQQ1ud
piX9+NmG8Piw+wT/D0mYgqZAaP8SG40Ka+AzDHDuWcorjiY6FgS7FjoqMBWQkjAMaojeC3U44dMR
+WNtSZ/UuMzdjIusIVaaWBAMPzHmUXgwWBzz+1UUEhr5m/c47ToaJ4vizM/EoevXOVPcFqcJ5y8d
R2TVB+ZCIOp3ycyE0m6AbPywukxglsWBAjE4TKPevdVkqAZu4UcKmdr3cP4J0m9/8/FDi8O7m4Wp
GSMsll1bw3vbh3g57Y6aJUs5H9/arr1fqeRzRZiMcIbDLynM7ZaVKoSiAyGQgx4PonwzXdJyDZvG
HL6ShFxGRFbS3O/HSUEORxkfwlU7n25uM0hjhAOlA5AMNkN5hMEKAwZNlAP9KizgfTg5SWRULjlw
6iSrJ1+WsObaalgA67qTsEc3sWgcHhDJkwjh+7YAr7fYlR138NlupPYbHuQoiciwQTz736kMi4cV
PHykO6gKP87YaSEOKKpp3SnvrlP2aaAYns/ACWPEl7cj2aah/IA0Etmql2jjrFyGD8XzIq+asfq0
9LpOLIGwCJLWFehhF0PydFfx/E+MDZJ3TOkP9YXSXsfx1UVVOCo+vwodRf+BPOgx8u6FYsDiJLFJ
fefsWwNYxZ+wFM0JGT9Ghdatt083FkfnVGczNyZA16Ex5r/LzJNfxXk+CUiWzMhZZHsQyk42UbCI
WHfxcRcsZYNl8s3jgVUM52ewZLTub3VrcK9ibGuk8TovBjImaBszriGU7fyqliqlaDgZtJ/24oHp
Efb6ofIh8n4bwv81fwOzlZgIOoOPxFezjvsMIlHgK0oxYvYmuk7RAd++ES+o4Z2hVyDJ3gR6s+RR
rABunaiX3Viz7KyqTt9nWfqzFyaAloq7KyfCAulUMVjjo1vc/5UcOn3nKdZrw1tTAQjyO3Yd1Lnx
7TOw+jjMBJ3OcI8+mAMve5W7vHUg2PUUahPgURI0vm2RS9T5ZIVKsw01vwDezdLS+KFE3zcn9UX1
oOdXPHtHFdqqGF8dtGdKOflf4T3AAxcq4Cz0ZNCXCwdzv4QEdT7msAhjC8OBKvtP+ChDovfemFNE
KKtUppEexaXjn92gayrsqhgVlxJeXj/2OsTNE+Xatl0xRf9dksv3wEM0FucnAGZnf5KdrHVR4wcl
VlJCK9LXF68Z8eK7U3lDV/aF7/Mi34XaeOY0PoE2K1eK5G66WdrvozHqJYQncJ3dIncYScf4vBFS
IyZBhGMt+v9liNhKlRov/jOfQnXWKByQYuivLmEVzVnXwYrnerUg+VMaZISf2G6QPlCbRFm9bYaX
WLblGhNLGf9lDgAeI1gEiTO3Q0FjIN51sBu0zRLX7/3E/8eJAWugoSRgBn+quIj9WSz5AlFfj6xF
OO6SKAnkDZzV2v2RqJ0BJOngW+5KcdMzlIAEYATECY4E8PwzuORhfuAXNfiqKKNWxQC/PLHmLCLq
4xtqVPqjNuotOwIKk6qRW04tbAvKvkDGWcC9uDaJGK9IItgnPK8oMZfg2zSJINVb5UtseZ7/3zOy
YZ3qYbxGabM5Nhx47SzzdhgED3G2yHEkwZHlIgvjrHzWoMuQY3F2abo5Ov37WhwY1ZujGANfH79r
HCeYmISyIXyHOWjMX4f9yTE0bqa/r6K3f7ln5TFLXyJ1gaDn77QF5eJArd7OFWuuNHumvMqglOnE
KF+wRNTmUhKQcuhJ9i0OjqEBkvNXZyt8T0S+laIRY0N030vjit23xWA/KXQY+bvvwDaK0VKv58R7
/Mxl1pwrmz3lM6cXMMgiYOK4oH4gbaYbJz+7vLWh5uBONNvHjqVMw790WIgjp92mrEm5D8YNeKKy
2COzfdiX8NkO4bixfokYi70Nt/pZ7zBbSIoMbnasNfc7JHcYA7+tWSCXoC8CwPKWasEAVxks4rFy
PRtnVEiHGISMUwnuFiZ7XVjbIMPOlUSQPhlauQrtu6/nssWjGnPYjRkp3z5TZ9GMKwgnR9gS3yci
RuTi5tIpgDvu5xU29NPzPkJRUQTijrqG9hMBO/ehJL0+xmt7qIKvb6Rxq4wi8lPsaegaXAl7yBTL
t4GvujsKPk67jnfVRCMzMu387YhvV8kqJQ9EeA7nb8wSJ4PsAzkSvglX4GK0SpmaY4d3wrFIiDgk
bwma7QN19Gctc49doHCpBkYO8wqwZeSPz/NS6PAnIqW0A0x3GtOX+VUrdYeuzK+X4ZbXczY3IE/c
u1EeonfiGHhSz6GRGPE/61FmkXCfrvz5jgTKrgftle+vPsHK++4UDVuryJ20wr/3FrWEB1cdP0ec
GeT1ULS9FEqtkfoKXM3OZNTnMiEur1zja1fftsdDUCWBYCTi5+oBw/jR5xUK2x6Td8fmOoGidC4B
JrvS9V5vYpfWeUfYwvcho6z3Os3RCMbu8EE23DORN+K0rj5Mw9cH0DXEm+GpLuxvrI9bU6gQZ84D
jtVlZjQL0LXG4Thjy+a8/g1Ibr48C7cvwTxg2U1ew99o1as6lzARoB1BDfJ2QuA5ebCZAjhtDbvA
8Ac0jyy4v0KOFXw7+9cjH1Tu6mMRnTBAr+xiOC8594gIqj740GVteU68m8Axk/0tMnc8nIvhFQMw
cZ9Io/FSzuCtYiTJ7nRyOK7ubMnVWdPphn3mwJtepFebZvNlFfO6gPVm0NSShUultFL0GH/dEQXL
bBDLxGy43GkvNhBhO9jqOJjAXSi+BdHxuO0Ykn99O/DuCReDK7PvDTrWKz+Fx6iBcMbLUZgTuL6n
HcSY20Atu5hRmjq4e5wRsJxmf3CRWf4+FAdxTY0slW67NYG59r8iGQOnmuj6UioZJZihstlEMhaY
sI6HN6ettMwRVkpBZAJ1VKGKZACoo/p4Kf6WxVGhIGUoStqxZ2RVakDXzGaNt+D4xux+m0KeRaAy
FxeZHU4sFRPZYuaf2kCIRyIpt8fbr74cAdDf9p6Csh66sAPRYO0GLbhoeSJJJbvd2GvMq/FTvIQd
XKpw7JlHJCuLj3SNp7zG7O7URhr4rXtdHfrgUsYkC0E+IaoAjUl98VL4EgDSAyX3xPVl5hpjvtkN
M8ckq+JiGcs3WryRS1rD/84fMvQEARRCL7OmVwQaut9YGtmw7OPlnQ6sNRyLAEulQjuzSKa1n2rx
25dc/br5oRzJhhN3kGRSJYf95tNMk+sLE/eduGoMymtnlA5zzKM3E7YbbPZn2yTK2bl9w3c/EKHd
LVwVUZv9deWxr8n0WXL5XpAjNWAWL0lMHxvfEzLadZmZFXK2yF/jEbu+KSlK1NVLiGxN7/5oBUC/
riRv315j3SiISVzx1DdLZHc/kZl+g/cgm/CXiJI5RBa23qyAejcD/W615NvIJgta8WjnCZnzS1El
BsDp77AToQUTZH4LKH54P7W70SeCELnkw4qDNkrjoApJWIoFlF9m5iOm1afluFIRwSk5fwVTXF/4
C/4IZsy14GnAlkaLB9aRX+TgGoxJP9jgwChjfPdupqgQ0ddLvPGs8qigMfeo0y/yydcyHT6tGHRa
/JJpqtb0k5oeVkkUF7bhgKB+PgWTljo6NUpsl/kqG67jjV5Hpnn+Qi/8rZYy2KQbCXTP60S1zllK
dX2gb1U9JXr5tqvTbLc3hEQzDYm676apoaJgMqlng7kbbG8n5lCAnYfT73BhaPqAh6D1oNWqpoU8
8v1+CPfoa2GJOhAB0WEPVSUzjUe/72oF9BM+GUYIuCWAzuvFR0BgQ3KvKLMCH8Ff6JPAsRKGDNUj
F5emj4ns+/syBI41KFIWPqro8VctGSDqVmzZvHPcLRUNoDwoF54tAMt1axVQWevV7iurG/scIGaZ
Lk7m98H0FP614LGsf6q3dBhH9KPlbacXzU8Sk/t67W/Q+woEIrvweFrerikAFdm+FIlTFt9TMU6t
ICTFUrhG0l3O7mLY2mh4ElcO+FaQNkZ4hTasXb7j8qc1hpubxMTJhF3NMS2DWdXwv93mAk2axOYU
x6XwN+OzWYzaGxS1RI21oiGy7my+UUkuWoLzVOyimAo+A6D2YeSm4AgWOxhhO0QQRs05eekmThkd
q5gyd2gi726LA6Bk31xfwflZv+ziKwX7i9wOmXb9Te2uXsECsNsPXpyLkfhIjHQ7PrM5lefIWU0K
j93S+5K2MrSr1phRwAJ0O0tyVR/U7coNEI6Udu5DVspVtaOoodounrDoyJVtjYrvM5HAF0dxpzaA
52jm2HkIAe5AyUoeEZTqoEYUd6o2r/FDFbGHEEO00sO9bhudL+E1YpcbGk9ZBLqPdPD/+dLmQLWe
kuKPP8jNoWN7QGMUrZ5umAUv3fL6G2yjMB6hVJ3aHoGJkfTa8FIzYr8qAXe2UYZ7aSZ5GKYurXR9
9iAYjZMKWd3Y8BCH87u22+b/tOwa3Wi41SJD0JFYINx9PjlZ0l4yrGG1e22fBQIVPEtwOO/4n7Os
PqSCFfTEhkZjZgKKI8xaoZ72I8i1tdAxszSjgc/fz6ONbFi4YjxDNL0GQdJgFR6qtIRag6U3xtfk
oJ8JM1XT0y6KTjYBkLkApvth512pMYDTXQdCr+5rWUbDt6F8yCb4YfAQCvcLy+7b1zWlBW+ALzkY
m8wIWrv/U5VqyvR077FNTy25eKAPAktOSrxif3OM5oj/yILScM1KnOoCUZa41MKlidO1iFXBBSGo
Y04+XIGqJheQdWeeGdhcQ5XYJexwJRaBmGzlNDdfnlHuIr/0qf2j9v5Bd3RpKnkEJF/i8Yrrr66p
xgJi1h9tngv6fkUp+gh/deLYohThkIhv5YUxR+Zvjd4E6QI1K2yIfB0gUj0xU3HcKbQbAy9KPamb
luAKI18Nza8+I9O31V5q1woEheqzRaB+lYQICRvNZKqVmImARhIjishgGi5fd1oVKSybWLJGv5WN
tD/mA7iy/WTbGIUiTB5iLLHaaqZr900eGRmgx4SmWH8TB+RDqbv1wXn1xMb0dHbYBpznhtkqsneQ
M+GhddZpEjT/nLgnDriud1KuPACXHgWAC1Jt+t2lNWoMvx4QmjUyMKJ/T6etVLmJhYKdeuGl4m69
ZOkZ6C3J7OjzcqUvcs0lnhFebGvb+KBVwsp8MUuyXeBdPT6NQ3MyG8e6lyYXRdj2fSWiv5Ey7aXE
uABM0PhigdGqXsyGR8zfBmSJ5ZolZUYIKlaRiybfuiLpfP+dJyPRypac5EfNyFz6Ba1F/nrFHkS6
ETsnkubaUlpjWZ2mzVRQDolDqqD+RTzOrO97M+qwQpsXPznFuY+WxU0jseC3svxQf1Ep4EYbOKwC
X4C1Etsrif4Jz0ENBa5sYJOjXndNzh4nr+AkUO8xS4LwYVJvdrSn7gY0e5y5elB/q5iRUB2dZf5v
ctxfSM3CaNjIJvhBrFqIq/0/ZNs9kB2Dfo/GyX7Jz3r7GFiu3338MR/ABhSkvMjws7imuPjkMzIk
YJj/XzvmTgx8oXlzrJltyJp1R4wzHCCcBDdOc7liwl8NH8ct4ISoVz0tty0Fgkt5lYlRnL2p5TvG
H85yDQsshrEsuWGAAzIXnomdcAoj/virk/j/eaFdtA8jSxoCNx9KC/wfR70QQzLvQpviiq+ErlsN
y0LjmFC2G6xtYGDVOPEyXAUnbG6ngMyX5cS7496Sxel6aaluopkD2Y1fW2uuzPkVPjy1rAx4qq8+
hkjrgUiIQGAw69L7pkY2dq1C7xJPu1o7tDlXKewiGQ2usYEiJMboaIrZST6CEGFB+MB/oG+a8UVa
FWs+d3BRv5YYbdiEr5Am0kvFIRDKFbETxA2aheFHM6UqvmqfpdwOFscKu/Mo4ZkH1QN8ja4srrNi
oLNwBDrAcICWpnCzPLFCZt2188wQpEfbMlQ2Ma0Pepr3b45BgssdB0XZdX3f3SFJOCAQw0MsBjol
0KdCrya17PfKNdbgYbxxLFBoi0wv7mHFPd415cYCP1AydKWsAf+qO1bAaKjhvpYhkivKH4wutGm0
shbOmwXUczN/Iwj3sz6EbnkLxJl78/Dj0SbUBlIljpyVYlIZ7mveEgNouiwH/Cqi+sJYaPH5cKqc
TBpTaARP5boZ2CbTstjbEbNxdlaS/ydV1gdFi+ufTkgnIzDJRcOiqjes0oMejHmBpDsjQkqT+qRe
LvX3s/4iXCJ0T6Ltgj9HBnEg1mE5QKjmJSmgXK+2piTviwbvL2a4KdxOSc3k4zM01SfvvMpVCGRR
NCQN1IOWU0zVLWbW91917k+9lzpiqMA33jiAGL66Wm/nF4Xg1yoY36IREhXfotXBWg+bJ1sEjLx8
eUwLG491TWR+zdKLZYEC8ds1aDQ7A86PZGJc+I6GoWv2mtnGQ0S1qFX5u7kCZLfA48JvR9VYXMZ4
WBmRw0oqdDbFiBfzCL0qZ9apmWBFnidn9NXB59naY/u2PeY8T3fmN7pfx56LThEm00BJEsy1aJk3
wbBl3iG9uTXgic+aSrDU/YzqpjNNiecPz2HflesRdagEQmTr82d3Hwmh+iGkQ4tVnA6+IOAtta2A
L23KPNCB+8MearSz/SNRB25UQSYhnRoKO310vlYWbUErPwGNrvmQpVwgzSl1swX3K2lgFLm/czih
WE8aPO1cRFDFS+lSXaxSl62I/NE9fg4kkQz9dQ1t7cNP4lf9Q01LLeniO3vnfLdWYLve2pguaHPp
yo6hTtZ/nguhUWiuNiavwHIEP+v9DluDRCVxpNQ8CCfAycpuCEppeWwt7dLDw015hGKW602u1e8o
JqOkE/Rj+IG2FwMY0Mevi6mMBba/HzZhfvSImurcPkDWPtDwx6yCJJke4LjBszlzhdx9xURNRl0X
xI7D/ZO1ASLsr8Gluyqa662KQOpq7KN/MINc9Nuqm5i0cAOn9Zuwrx0MaE6OjPMVIjtlEm3n46ak
jUCAYS1fG+TK3MuB0wrTPNuL0NhPK1OJyVbXq7zUrsn28vwo73XynmU1JQgqDTJXUKpoVPZC2+li
NZnpws6cuLVTsxlYYEHphuFhDAhKzOoJ+r/Y8nbNXuVi/4wjV4zevRHTdSlFofgJEdb+HYChF2Fu
ZcjeJTNfp0lfQ2ESDbbdf/t5OBPP4qZO6idaX1B7uxdSD0mumMntpRzKT06L0yxu9qi+ttAXjUCC
PlMh+QzqsrJcvPuzY/TUT8yMW58XPjeXB+2HQ8HkX52bwfpjk8OqcgiGLd7mmaTbyQgIBp527Yn3
yCxaj6E0n/w4D3zlYFUch2kFue8IoLOoWmZZ/283O2mE7UINGWl6LyH7DAC5eNg42EahSCZwrgCj
r1gcriKXZbMoQNxvEELMOUEmone+2Y8p7EWLdLEREygCU3VZhg53HW0aMW1jdXFPptCMDcROF8PN
80MNvdpNzZg37CU77NhFwoXI7T5o8t2zENgFlJj2NiRCHNGiTDfjbpyMuiSBS5wqx9FwcCWg1PQv
ajOQCei7QtfLRCWZDMuqVwLaKQZniqOb5b+RNlhwreoBXOwYE82DHMURo/JTKGl6h7qpYvurncUX
q6z8W/UMqK/lee/UYIcrPDZa3UoFQZcB5UJg+65ShCMWvTpH5YVzK3DXv6pXY4HcYP3sWElT3XAf
wJmkh8m8Q8D21OsiGlPYxuT7c3CqLDInzSCrmcAmfJ/MjzzOiOIWhZNfvdUQxAAQgqwbYEr6qFVe
D5gYi9STrjAz4UcVEfeIVFjFA9nkhAwQMhpf/BVsE2ykMJMsoS0UmK4QQAFPsv+WxR8KsoAQM61u
mCzYvaVSFB+RMCxFVxMg8si3zNBV1lV9gmP3MAFNh6fDZDT9xw2T4vs3R7iTiRKXlaqH+5o/05ZV
JrsUhYQY9clKK+dhwDlejApREz97f1E3Phszs8u6i+uB4NG6cNDgSBgS8bHiAFeQTQfjqsxGIuzm
C6Xx0nNi75MPXbKa2J6FF1GpxyOccBsabudLJHgLP3CkGgWZfsQDZt+0YzwET51h6n0Ge5uXZrz1
thWAZQC6dBCKIctlfRno4ixeizTcOSC8Rc4zOimAKgNw+0W9rPU9NqMHPcJPJMJq+RFj5qmqVqzB
IJnCicmq9uvisE0TwnH5fXdjeaFw4jmow3pH/FD++LuxZp0uynfz9OVRkEo5fF/AjEAUBfmY3my0
tPIq1T1U7KBQ0y1J/DKv6N+aSuW3TjL1JVPv6vX7EovfUsWKSyOgC/8TnnwYyNFMDZcMDYyCqGAx
EsUr5Lj7tpsWGzbtg8MPskSwvtz7ZGU7vhEJTsysceCV+QewdNkqpzO+MgYWcTNCYvtBu5M6EFJN
iSKxCQd7q1nXSwtQYHn2BS5+k0Q0DvislE6IayQgr3mpChfzq1byKdUOMVRQrhfwIabLpZHk2elU
xEWWPYVZJgd0gE73FZ89JjQqbqGTx6ME3vqQJo2H82H1LKMOC9nDyNiHwS8UEWS4aR83w/xP71f4
/3rBLU/vLAFhaxk4prV6WMvjwtyPBwQLDv9znXb85zBHh/r2+TEE+F2mSEEQ2vqghQYpivMSvrc/
LshACxWaTGpATbY4XWlxMSZeRdj7fEvCfkY2LXjBUYCgq3GNjMqoU4KmTRBRRgR93VhxjBvIfb0z
MoEbyEZxVoGuV7pzWCaSLYLun8MFfSAd/jY9AWmFmtlpRPgVXxUo6ai5PbfkTqd05ViYemlUZ0gs
tC9p4h4OJIa/HJbyNGcmrfc5wt7R4n4GV5W+xXfHMcEN4n6X1AjHBbjpvCPBVN0DkrMvPtUtSugu
9O9uD2kMqPfuSVxTtIp2OT50K9DiGAHrpviCqXtXgZh+EmNAbrskceSLKZNYAoK3edufTl4Ok/ac
e63QqTZodb5Nhb2ju3ze7cWPgaqRG+xQU3UbuiBWayu4gC2YC+ZzkTszA6g1H/SyvCLTWyFMznJD
WPwdPZbo8sA6F03pyQ/Mw8pncetn7E5xzIcedP9gRauUK2Kf6jeDEl02e+GbHUAE0or8XDngyZRd
m05Vaa3GcqHSKoNdVMUiALWiNG4PC5cp9dtZA+oYye9iPUYpVqlbSFYUJ8iQTJluzJ6RpSe+kOQf
aD4DxsBBp42Ve7o6yvL8x8IsgJ82O3adoPxJMze1GuCdQKqCrej2B4UleJ03v+OdLIuFTztztnju
XMSTIOztYBbzGJMh8sqTnhQLqH5gnEVPvEDA6awxC4iNIJU+S2ANDt4Y71ITxC1bJAkCJg8jgKsx
oxUx/uFf4VA3vRnopk7PQW/1A8+0ZIq6jr/LPQYWe9e18ecfx0/UKoeaTxFaqD8YiCLiN9jDNOCE
77cFE5dxkMEhAtP+NewXXwvaqDlH8uMQnO0tHQKTTYY/VtLCJkrmMjNGKaHupxiXmsZe9sHt3THA
xzXTmLYJrED1EaaThd1bRB7nHPFy3sbDgfDwrN7HxQngrdc8iDLDdrNoXprdb286sgdp+YXXIsQ6
CUOSBcypB+DN+h/mvL01RjkS/dhr7vT5dNEDprpsvgZXS3BEsu2m571N4LXr0X9ctJbQJjdGonVL
EH2U29FCPcWS9EiYNBDhEykxkbEVdm6os/PW3YTDKclvy3fvSQGZB/wAP9pHKB3JB5LJqsKt+14F
UrdyCLYWX8sCmw0uw2UOt22cVfHk1ub1csZ4ORavbNDu+DL3kjzDBNQooZ7QvPpSeh/mkJugcc70
JeCONCuQPa26b2qPC0OZmunMHICF8nRJgsutFpeOeAhZaqNhHcvOLPo1hnKpf4+dV+MglBOwiTpw
+6VhybXPTEUQc/CWCCP0q9IyGqNmC9G13l2rJIlQJHSVtRkAuRu4Vmkip94+fPFUb+WxAIxiV/jq
8fDQK6n8q+mSV5dmJQSoxpMLPeJLIRFMkspK9rUSbuBhvKY07mzenCU5W+F3pRIlDtSemLfHJzJZ
NJEuingytzspPr0qxOBgvPayMI2PNvVS/sMGz92Hv42tq9J/kL4LgamktQXHRqe35l2A0iSVN/Jy
21HISK1TFmFx9MVGaLxR2mNBdqH4MiU2YJ05poghRCHj4/UqDhI3UZAK4q9lIMdYysvUDV/b9D8i
wEuBHV1YYtFLZWWXW0QA+4LYtRrf9OL/BO99ye8CQVWBFV1/52rfSuM6m7a2MGVpK/mt+TP6rqHO
OEKvwEJ1lFhJHJsqYwETK1mrrHXq8VoqyoPsZ5/mO4zTHI8vGZC4OA3uA/u1G+j2f6oOrbxMPlBY
a0X+S0of1+DH4bCqG3zusakYwOWY4FWr2gLdAtPv7nlv7Vdy4IbVdtjvQx8kdVu2pZibfCCLKdrj
GLINuJgX7BarbevMMXb04kkC4g5wWiFzpQW27z72nYZOyMPUX7FZEUE5fDQPSWBczzin7r4IfG/f
HDoMm64NRfRMaafZZv6GBYKqmNAR46GgsAKDQSgx7w7kAAMZT9QGQo0J/vORYVe3SDnhPnbk0+5B
JF4TX+LNiNptJ1ZdGW9Un2piqi3So7EU5J04eT4RJCC2F9Z4YaozCpxLK654ryXI9M2ufyFDYoP6
s/1oNmYSNdZ0+cDrr8cG8Td+glnYTwGEX4i/aOhZ+CxiNezriU1c7ZaAo0wkIRbo6UdlCBChMhM9
+oAzRl484ekOk3VzdukgXL7V5MU7RPahwlEhoLd6kyAGFDMMNcwOg5XgvK3lGgn6OPGUyDzYh7nU
i+XO+MF08bTGYVX0uLtXgCN1krGTLqDi1M34JiXnvQfJ/h9CS4EboRLy7hNyYM6TubnFltcOGpMA
vskwOQGhwDMRWMJa1SYTOns6lsW35E9TxzVqtx1zSBdBCQ09BVlzuYB8LekhA8LpleZnhQG5rp1q
B4MwSz/Bdz5YTRNku5Sjc+JfOrE0iwGELp7PcQk7uj1Cwbi1XaxDgvPRXuHh0BVak/nbcfmJeg0d
T0mDPHbeKnFv3H8HysfE0fMpQcGvxL1pDZ9eZPED0Aui3Xg7Q6Aget00cpmeR+oy+kZcNW2hhU5P
cfYQUHWzmYVbvZyWu5+Eeqe9NzK1NJe1odoJejLuKE3JGPc9VY1tjYEoCTCRYElL/yzzGxktKQbt
WOSyzNEHPaP3sDkuxA3Qwvx6675RAEv3K0GB8oMjG118mib9bp/CzDNQp6h5UrjTehSAvByDHvYq
hpHsSdi53lKETXSrKpyjwh3wevibMANe8y4KC35/FodbL0i269/rA646GLM2GCfSCRwP+A96j+AT
4SXCX3qQ8yF0xwkPfrQ4SCsob3+QX2PvfZwe3KHNw4staOdlVRzsaJz16lgk2uIt7gqPMcQxtQrG
U2IxbCwh4GTENKjOnWzuEAVtSZT4y7mxZz5E1wskrpTYMatukHp35FzkRydHC/t2BvZacO76rdxE
UBvFfcBoRJKDwkRZD6A/EsK+aCPrsrr3gpwfFKsc0WbaWczJQYFNUfJKaAiHfKB4OXZuLfgwPTpj
uOw1cvgUL3/Yhpujz3RUB6kaVZ5FZJqMCiL6pcVtR4SnfCjvBxohhoYyKxknTjih653ncHZjSJaK
Loj/sAw1G/fHfHY33aSE7V84xFJjgbFeiPnQwg7RaBFcQAam0WIEkMWrJVzyvNC/1p4JT10kr1pm
Velw1OqG14RjqTaxxwrzBTsReL2inwYyK769vCjnK/+8q7JsdEtoPuKQaICIi19cZwlWhsmYGUF8
jVm+oA7lJSpZFwKghPVE2T9VYPGkYlPNBgryJ/eJv4UzBKYE23PovXkE7r1EtN9g6sBdpWz4Yzy2
hS8DkhzIRh6Licw49QQZZG1B1W3RupIlwKRfySOrOY2BZoZbp3fWPcYu4/FC5TA57/5fJJ+AizGO
16ReE8fxKDA9oeBHcG1FkEVVESq6EH4pUPmGr2zSBpkdjEZDbpUE2qwNcpa9Dm/SB4Rlqvyh3Sqo
VMC2I7oEOJrobccLXmibGcJaVmcZinERZIZlh4p2VPIQtUMzM/s8FBWQZtJAkeyXG1CD+1a8Pof3
FhAh6uIWJ7LbkcUSTpEkMWbzOpfCIU4UmOA11/ZHW/1KKuZTLym9FaRSSKVBDsyU55lpzxl9iJFa
L5ojotDWWl4WwhOBpNBidZ5Ksl1EZoOdn6oyaw8bS4/BwcRAIKOJUUhQz85TDs5mUeP3uFILzAvl
RJVvJwUg5uV8UyIKaSCx04Wrp+mlLq4owEdKCGrKwkdNdE6tQ80QkeMEqQJdtXoOT9CaQUT98a9V
q11jXhD0ixRw00pKcsGQNBG8NdCGGLfqzOvTwaSHuI8wxVmyxBdOJDrrbdvFLmU7ALXsuXl2/xeB
EKrMOg8K/krN5BHnb0lNSX4SyQzERQLrrYLemj/PwKhRhZ8zMIc4GNKXQcEjf+DLdG1ZhMPqkh2P
3YQAOBum0Mw1L+3eYZnGnn4+ev8pTOn7LHAziUVEEAS8PD5boYfWZf+mkPRxQ1OdJAygAo3Z+Suz
vKfU8mnc22cPKRtEyS2HxNK1l2KpJieoaKet5/eO9bx3XalyrOObeVyRqqJ6WtzfhtzlC72kAfTJ
tuQtQ4tipzZ/sgMvwCRXd6oKJOleANaIzcf7HzTFteVQ/OOq+rdikDWXHCVDO6sE2pxqiwlvb6aE
CD3owjG6WEmYUfCf0Ply5O5rVpj6xivIKY7WzQyx+f75Ejy0puMRvZEwmBbE4wZn89zqa8/HHneb
g34Yx5SiJ+EhTVoLqhuQ/ntVo7pNc5340faPoICksdpQ0zY0nX/Pr7fOcD00h5MwIFvGtGTd5l7u
frqDXM6E2DHRrHCut/K4YVT80dyLSiSHUeR5N6eQrqHD6fHutIfAE/AzKMFYbQ2MmNOuMik4pTAk
uJ5gebIpl7o30ykAWggYDWwQ7MvUbx/V0X8oMXHllu7rBrdd1YkBI9OmVrRqQ5xGblwE4YC5TOrM
qOfUjPby0OCaw0IcYvkZb7b++RfDH4yZ+5x8ef3EmkSj4A/xAvPJH7LFPwH6ye161pm3C2z4JXVc
RbkZpDVWDVO1BgXzS0j+HzxLXAjAbT0voMl+CFN7Sv8vNw2aIpZWnelh1b9HSkAVH1yhAiUX8RZ1
/9Eqs+E7ppJEpS8uunXYxzbJl6LXoTmuhs1FuACXedRa+VctFaBWmveEDKuT2h909fjczPKoLsnb
py7XpPovhigr5sMDc4ogh4ZQxfJBdiHTB5S2AGJEgbO9mOFAyQC2ca2fbOFv4Cbqpp/sExIbJS4E
8cYGPARelGf9cThVd4hBmc5hAW+TY6QZDWcwrlzRoC5EkfJY2LVfEyNwA/9WEd120wQ5KdDJu+N/
JBpnwq5aZBQX1kn7gG7+ec3QuPzjKq8DrsZp/afh2Auftqxdc/QvrHiDUBhIsyrh9djM13m9UrrV
eO+/a7jhfIdnCyf6dpzNDfcwDxxI/KBPHDYF7mprA35OoppbjbPi2kTR8zmtFpKJgGrSMBaRXhuS
2HKIhQLwzhdeDRrqJdL1PcaX/NpH8UyJg45n/xqQA/IPqCiERHlKmOebda31KovNoe5p8mEiEqLT
5SSI3wJ6eJfkGV9IrOq5SCcDe1UDqEJv596rmyZ2MiCw3m8OTZnUDzaNHZaViUx+94iMFHeSReGk
WbrMb9WCdLDP/ItilRqVDymxOzP/ZCVZrsNO77eeuQk+zosBbIli0ZO5wM8ndPCr4hVIuIiDx79m
YH3RQH+dvfa/gF2YuQKWhPsvpq4BIFTS0l+uEaT58mo/JVj6V02bczpkJr69KC97wMHFg/png6lF
P/HnG8t4YYLfVatKy/jiN+NgqCSlXJOgSWjBqsEsL+MQoaz1V4cn7ebZDls/wWS5Sp+8vJo0YXDh
zldMbawb4xQxEmXLSbLhXGH7Y4lybBX8fh4kRe3fIgmAh2HyI6SZE+okoc4bgYpWQduIhY2MytCw
0zDok1ZpE95bV0ZiQnn/a60rfsXXSci577VeQzU/d+mdIAW/8yxxxri/CK+uJ3aQp+0R2EAxXmW0
YppRUFAZW4tAUDw6zjEwCc4vEmSqGQVzdNodOqSJN50LuUuV90za37HAOQqObwqWDoNYwxFwr3N1
rtZfPnxR3WEU8MMCG//hgnn2Lk2rNKf58WYALUS0wIeLMAgch1N0iTcSshK12XxbPX19TWi0b2vs
iZwPmw8PzdA00TPIjdqbm/TwFn0OE8jzwgk2Q/9DBuQWhr3ki/WLsPLr2RnbsnAw84mtF4SwDVio
eMZr6JrVX/4Yp1PNZqR1dLatwREvREsEgoY1EA1PDIsJq4dsJgyhTPOTKFHQEos4wrP9k1ktG3OG
SekO+h7aH9RYi8RrTxzGuAWA4G8VKWSr7mp8G1BH7Uj07TlBkxrX69dwDPQzSFEfNWoD8QlN2Yue
LV3bsIkfchHa+jkRBVmujd1Xjp9YD16Uh3UOMzPAUagD2jKx9tgXwT79P3MKQm2GeTr45tD1DnWC
/2Gq5Ryvgd5XU5IrPLqaE82LNNh3ctCMKYUj7HLMGZZWPp/3jrBo874wIR/TkhK+DxPoU5G97wAp
dh30mvbN3FNjZcILknuY9bNEj1xGIxxzPklE4fGbfChTn/Yg4krLwNzrsuri+UzOYsGjUw6uAgVq
N/giECrAd8PSQaS//hbOX0A5ov5tXr4r6hk3qp1lgecwoSKkF5j+G+WEPoMA+uTLFmn0JtD3+Ygr
9in1nUx/l+pO+V0WDYgDuaaCBq4tMRxciWw7EjWFDyUEuRJoy9NNdzZQOAxUDabeLVOytJ7fHNR8
y173WFjsTkjYAFCNwU8NETAHMPegvccbYAVAGiweBrrLjC90ZQrtg4XyJWBr8Mem/9i8+6r+HDaw
C/uk2yXHbZzVH7mVkKzcLUaDt+Ho7+kihGWDszQfHImnb3jpdCnb+gRpSqavaY1pxcf5eX5sxkJs
b/0rp0p87HaYp4g59io7g8bQuDs55OdSbJqOmvCevvE6Qf8PpuEtB8S1mwyoxV9eBr5kaG3ltpBS
K/Q94id/+bEkeqjNIpiHWLPScsNTXI0oO0GvMphcoJjYq8nCEoiANePV2yFV0NOMMD2BfYSLde/X
D4nm5HMAn0I2ssc6qHljv+Ijl5CgxZ5eOJBHGUuLJyT9udTTC9Jb0/PEyrYPZO8Czi2luW8HNFRt
YF+O4lPulYr8xyZh1H89UKrge6SzpFJcL5UcoJhVzra9hDB37vboBSR14z4TQImoIBiCnwjMjTfd
f4L6coIVbc8mSxsHp3k88rkePa94SaiCYfeOgZqjXaoMTZj8KLv99rzBa1pORbanZ9SZYBbgRwNo
RMzDbdyd/XVzmAYt6mQJqe2Ci5v8hw/BTuo4ydg//x7uXF1SnXsWxiAjJ59iCTHUMsqTVtlpFFLu
VgqF6B/oewjZOSngYj2fqLmGqSmq+6ioNo22UdNv4Y18P3ke//HU/LHBl6MKGwKVm9Njbtf7/B2r
5b3M5YWfXXaurx2Vf6es+EeuSKzkFk3/KTr4/ey4sgx7PmnjDP8WNX+gWO/rVy2VFcR0bFvmVFub
eNWNbN5bDKzSJb0NN43EQbO1dNHYcAtjG9tGwCRHGFJSuQVz38n/nwuaLD5SS7PgewyG94W+oVky
UWGAVABIHL+lS6IACjR1x2G4JJ+KukpfZF9J5/WqF03OvSFc7pdOSPZnYoDv/lv32RGd3I9L4DJN
tE/5QAU+RLGB4hjJgfEKtrK/DbMGQewA0iUnSrI6cUXViFLybsFQyYjDldQcY9ixHHpyXFWikyp0
LkUm3Ke6ErdeFlIltOHzGZoj0pSrjgfVsnZRz4LqmYYgmaCdXF+5gEX5z9hvy0/BytMJIeyRII/P
Da63EO8GCUDoXSTl2Evujm/IQeJaSLifN3v3oyygIE2WbvjV8QnTWDz7u6AHwNDfxg++U8b/usU6
V/tmVygQMgVacbUo3Az4pDzo2952mWO9UD0Zgu659GiW+lrYM34mpEX//FX5wJgjb+AQszDmP7IH
R9AEE/i+seVzSGjWrI98MXJa0EGsWkVZp9OVKPkoWyR1ngy0qTLi2Hp7IS67y4iIKwmCcO7VzOYb
ZbDuLfvcktIUOBJuQR26nWj7T7aC5WwyLum1pZgL/zERrM2MvoiSXTJAZ6Q7ZAt9DuLcNFg0vnen
GGCFlNhlOSwQAaFlXnXHz0Yi+rIuNJXfi5TpzBNSDhAakF1VJ2a7WZ2sYF2vaPB9CrpSsy1RxAqn
a5XQ5zh4iw84Yf0X9dV0I0ynXvKhqMGJTPVNwqtM9/ibX1Dt+SB4A+v6Tm/kic9J88scV6kK1cZc
lHm328ringdu6rZiPu+dwVzvDWUgsReas/rWBTRNngdY1XvMvwOpPdbOIb0gsLXY7zRTNYZ4KFiB
G/vgWDJCf96l6WINN3ILqXfYw1oRSEBUUwXLfnzGqCWdXRwddyo6Z9rledgutOdZ/Hq8NMhiM0K+
iuBvzifuxsZssAvgoPfURWD9ob65VJ1NRO1+QUi5gxCtxPDCQlSiBsXjqG9KtrvaL0QzRUwn8tcN
o2M0o5UQFfPYnvU6XR9AzoLnW4p9APIXT8A3zqnLA8mM4RLpq6ddfKSBAgmALrUJuWqjdwvRQyLh
NZX5TOp5tXwK+5mnUVml0yX8Z9oFRzNoW/RNi8oEt66a77fSM0shDL690AtEyKNwolNodIZxaWCI
xCD92cptYBCrxWpV3vVeD/ckcKUaxbbzEE4XFsgNFBwmRdTM3oz8yyCcQArBL72OkpIWFbnyTW6u
DptZA17CIcRYzPKcw/dvIsNPPzk3PCjSycf1vqtid2r5iUMGd8y+6v8Gk3J1H6FguKq40dCxLH2p
qJN1y00maZ8Xn1HXBt74d8c6n1/iNt8VT37tuyM7wZ7AL8SRXAUW+vYQNgP38nsHOWtTjFc0ja8Y
SetKLJlOIs7hYSvEyiVAUGSFAuny9zbCoscjxbBSTIuQEMJlCv7zNHLZomyobjWxb/1Ja1iBsHeN
LNQvd1ZRbi4d9EjcdycOYZXiO4C0JIf6H6jINbwp8YGvaP3XYy2NtQzqKdpwopDaBZg+A45I50jU
BFwHVdyjtlKqgEzgn6IwDszqC8/u5Y6mwcOY+s00BYJL3jg2zg5ZxJq0XY7S2Ss7pXtQE+bkKT5F
MffTMc9KIhyTFmZLRzk9NVdMCPNqXUDIhv7RQNpPOAQRjukIjVPwBBC8NWrTQTtFanqqieL/w+EV
S7gxexHXBztXSH/IbzbktDnCVm/K1UIQ8QJzwJ29YmvDa5Lhla5XkBx8RDPbHjD8wydMLuwRTq3M
XFE1sPb1FU1sGbJcp0oA+rxx1qkgkJvzKoVbK6msPPyodpb4IHcu7uEcH8H2qRUlPi28LQFBkzMe
eg2H+Nr/P+hhRy0mEYnXb6n0Sbv0lS4jAY533OFc4LQ7Lq/VT7VrYQXuTmAih1WdrHttcBmHz4RY
MLFpdk3LKnKTspnBFnENS7UHf5cpILRpXd8WFvQmB30Km06iJBISnKuFh6mSpyWVcqTk9VoAiCDv
J8WP2Zw7guwswCoxeLSoCxyr/dqCjdKOo6FIF6O0ECOXdo2w5wmWWnKTkthHWaI2eVRQF9nXhz39
4s8q+5K8o1uoQJfdb2H14visfHy2Z2hgo0hL7bnYPqGNxQeoc5Z8iNO5MuXugoNeoXSOetan5oRZ
wLhUXi2+OGym4Bh96Y3mKPbMnTGCYM3yOWY4cvaG1hm0eAl0vk0gYOoXHKCW/WN8CWlRqAWQF8qv
Q7Lh6/fxxMRHL3oR3AGmaDwP9WxoYMMFDguRH/O+G9jg4Hq1gZ96LxlfDEbqPckHcfrjQ35D+smL
W2tCXA453o6w0sZmfhj4A03LHOJopLLfv6wTGMumq4jjUdDzjZrG660rQzRLBQG/BFqiQZ9jDq5j
XmOdKtvwg9wnb+M2hNaM6APsE1mWw3YVGFfmPhr0/9Kk249Hu2/+5GOaMqE7GtIXjcvUHr4+gu5c
1EQsXmB4rTmny4/AFVJYSSemkZrbsBw0g6V0PsJnTJw7A+1daH5v1BHHTgIOszkun04FqU0zNysN
QiQH4TrbrjBAilIfdayf4aHL2rpRZvDWK4nZnO2xBYa6VWXKDNedAJOjDCO6bSplUpdHjM7ztzAh
2OfdCOTSEcUGjTJhCt/LSpQyQSR2gsUYZYPqW8fXLOKcoMr3u4MtjIM+6cJdxhfgFQlObqI1ap3w
Bh6oQDnMO9Sbtv75yq+LpQsz/2WJONV3mm/LUblNQyy3JHUC41ktkTP7pw/TR2DtzxNHmmZQEMEo
+o7tfKctDDSfiVKmEiDdAf+Xa5yOR0WNkV5PEGHn4uEZ8nD3M47aK042cYmAr/q4stSmgLyXoSel
KzMr0kX/qh4sAdc3a4EBnq1Acndv1IsR2SqwDyz6xHeGouNTbpkbXlJ+/5CxM9EKs2XuZ03UfsyJ
i2eTFhYby3XcEF/0l/t+SYoOsJGwhSHJOtX+KkNeDFswpygqSKwAV3S+VrD3be+OOMYKU31HHQn9
nSFXicj63LeQAxK3MtmM5EzBpMibEFusIjt3ZvHmnLiVH5EQ8W9YmIaDKRoBwKzQkCL9Ci5l4T0R
kt0aj8ISNdInUfXFs90AjJ5CrCoHPu+Drsu8BqxTAOIsQPHOFinyFY8kbfEU1lmSaMYaV1+YlIRy
oS5l/wk2hRAwL1l4nVp2E9RWO8RG04770wlhKU1pGFluReU2vLnthYG8er26qCnGd3E89jARqO8m
PQbos07Uk/61JdkA9sIA7uNaB+rgNprArtROvVGcDrSpmiYhEuKlSSNV3/ukWxp/87gL/vKLZNaz
N2/D5/0dI62RI5Xq2b7dUawFtF22fiZj9+fIZhN/nD5thCAnUfRX8+pKrFSEtllMs7IoRLSISvyE
7ByNCxcgS5phkSryfa/Tbv5rABhpwbO2BOXr6nleRFSFgDIHg8uOxenf/FihsLWktLUjCMGswqba
AzHVQw9JocoT/e38N0/ozEBJG7CSc3Qi3ebHXd/QUc2IaHrp53T32lo6Hg3GXc4GbWX2dG1R4PKW
DHCPnuBIhqJUMHnsBKh1SoMHi4gkeGZwhY++bbelVGJl1avs9NuveMxZWHu9vPSMyALrbz19J3qf
fD8mUdpEnpjhfNxKS05lar4nm4w5yxknU6pLWSFM2+yqDfjo1wkA31BrBkY3e9fcvfC337646+Xy
QkLo+G9MSCL6rvTm9YXxxRm4RY2v9MKNeSiOj1Gg9TOrcssGJutcqnlz7HTUop7Q+OL8afWyrD9L
+Ir5Dke2edZnw0P8Ykh/BLgZXOENNIhT1kIH1PggCHJTML1uABHPGhsbE0/r2xDegZ+3g/9KEw6F
Spgi/X399CYIRcuKYI/g47tUnV3Qs543x0AzOq/8r/Jj64Oqp5Cq9WRH8+Idr7146u500t1GWY15
5x+3nn2L9NrPSTUO49Y+5bV04KhVK1EXYbj3NzVamaofehdeBajkdIWPctLbNpc7VqTGtjAHUEyu
A4ZwW6GG7QfW6uS6JwVOGPe/vGMQRjFeT9Vp6o/3FDdia8o4DDRdvCIZnl895O/54xk1ho9/CVS+
AcqTK4GcMKCsqiPoc3kcg1LcPzFpPnGZp0YXbC00GK2+EvkNqqUok3kjOlZ/+CZLa4yU3HO33ueh
UsyXDKWk7yg4AFaiemHPMtAuD8RsWxtGreg6QdrCRcmv008RqxZACggI/jRaG92q8NM3aXMtKB8f
cxPfUayej7NW3jRxVKMF6u8MfmVsVGjDSzkagpA1kkL2YOEHSrd5SYuaxuN2RSImB5ZjXjDee3g0
UzZxUhAml0IFWRxaHl9+BKIjlhi8dug9O1st/dKmlCDzQBDQVgtfD+6T1CK1ReIKFBehniztaYO4
+Sn9+b8XfMnAYII2nUzp23napImxYnPxcsVMIdbGJftD322ObnVBTTqvGQIuyv6agR45PZJLNLfc
UwBllaNSSS+DO/H6j9UJr/FSI1yN1xsPkiscDyZI9n7qhcqfkV1XOBMdYGcG+0Vz7cXJvMomru/Q
YVIiIm1grr45BBnfbpDDg35k4xdDS6zJwnssTsddPVBfE+Pmk4Zyt1U4+4d1G+6/4KCJEQArvKYL
saHhmNNBK+nOmJ/2WcFtNf60PpqLfg6hLd8yjQU6SqbbCH0GNcqpojNywS5fjKLAw8IZY1HaBSUv
gIQFyOpaLczO5XZ+oa4dNdDiwYrW7ZTBSLVR2fif0BkFep63s9RoX3ChQI1mSu7oCMqflLBcZwnQ
pN6KezI3SpyiIELc/B9y9829gYWD7CBy9E68wVcmfmZck9Su3PcyJ+qph+IsFgwa3w36mOEZ3xYm
ItxkzgDsQ0kZzOowD3zDhZnAxreRpgilRQGgX+RJ4njA6QKZLRLLRM7ME6wV8M8TthgnmVg660gJ
qZQCShKc2j/28jlhdacZsCXvNkGXD2jPDQy6+wmRo9jzxuCwq/6z4Q+E/9+DTgBE8fJT3nkYn99I
Tl5cMNQlwivRtGBk/pq23F+CcSHZ7+6vbHsak7yWN+SCCv4cZHWAmJDxv6JRO7OPS8qUmcbwo0Lo
IpCyrc2v31qTXwoHyqmEtX31yTe2q6KcLmxlyyFiK523ICSMyQF2FNP1In/NcCa9lZMvR4dcBEo9
7szaFWmMKR7MKNIWQgYMPv60YY2AccFBKtXcsUrH5hgtbI80tXm6v/aohiZduk4auukyz05ySMgi
UpqRMgrB19LXI3QowDscsgz19sdY48bIAm+rjPeGjrQKNXTW1Srp2FHcX9pbLFJbn5mjjxrMGWM3
2dQGRHtPmYzxRuSVFqSgdfHgha+LPLfFlfQa/CO4mD/yheBnHPEAx2MVzQAPHtn24ilDL2lIjoYd
1A/GS/VfmWvQQhTIF5AOqxv4zdGWzvXk0q54q7BhS7r/ZZUoLn+SQ+lsID+ThWW6tAq6Ij9zk8Fw
izd6VpERg/OCgPJCtQDSiRVZDgwezdvEIsiwNgo4uW6rJ2xXgk52Ip3oIMXEDCacLVPMj13ZGfh2
YDZvYykl0SMBz3zaSnHQdVsjBpBPA0IPBYPsyf0G5GP3x6P6B7Iis6Gwab6DRHTiPaQRVKu4Heya
vlhDkp2NVhBYwiseIBCN/4KpTmaVn3+2+9xobjFd0gEso10RCIE0Gag9MJ8hCQX6irITtnx/Ia+p
J7Xcmf0JruFpRS97/4e3J1ttC5uaAvJuJ3Khu9dYJPn3segfZke777e45KEmS2kRuH2EJtZSGXWE
WzqaAf/GzKzKk2NcXCORJuaR8xFT2r51U+Ua7SqR3YasJgX7UVTOY6hATryskEtz5O9RdQyWnJZT
7sD2QOcx7XCp2Ju5REI/jC0xyslOzQ6XZk7Te7R+/0XMHYTyAxU/JsWQRAlGN3bMYvEQVGWmuuM3
JKeV67eSKp77q5ZnI0RCuT5B3h1/Q5gnLJ6ZBSicto/lW51Fe21pNaQUi+S5dQcBmQzmHzCRlXoS
Hdg1wVuDvakQ3/hN6xc1fGeotRYvsc9QadAJQt7t0aEpVHNyfNXHru9tpOfBVbeelbIWxoHzjcYv
7hlZ0sXVXtCaf7SR5G58bcN5ygo3bs46j9YCnIArCcEpydZNq6XkGZLBVj4tiw/TbNNG1mZTCxPV
xd3tkfqFtGI+7w8xplSKPX5qCPuMG2nZ84o8HCjy18SARX28AgpFzsRnVwOHTvrLUZQbliMIccqx
kBwpHqUG0Tw9ZYV4puYgxP6aszSWq/JsUO85SvAtC/3IuQz1snenR9gZ2SF+/sg2goLx7UZgAdFV
fUGbT3Y3Ab7XfFaBXtYR8m/yXrV+iCDzmLAuB0dEcheTa6DsXtEJz/XjvOU0etAZutmKeISvioXQ
gUDCDOsp1g1NEHkB60B7esf1uuJOND5lgCwZSviptpKI3Zy4aoqfeNYNCTwgDsbLfi4NPbJVM5se
nMWTXVjyX00Qz6NXGVW5p9rYyK1dhapm9RqKtYPmoyo68shD4zY6omuiVzhIurh213cZbxFT52Sq
Z02+/RUrybXAJLzxgjW28wSJsDB04ZPtAVpZmS9WKWUTJ1FElO98RQS6zdNzQTu5xaWzIQOsoIfe
ImLZTuZ7Y7Ke8g54bkgZn9CcZVjSTjDeC5fbqE3git6Y3RQhS97lgsQ8Z/t2xv3ofjC+jJTlJYjq
5xKeFuRdMSHm6YpHGZrJ6preNt4NTQXs9p9KUomkHmGzCniRxwK/SPPORQfEbw70+eNZm/yF5EKa
vKtOpBAojAqE6xlgIMVZu0DQk4PvDoeLKOAMK3NfQwmsQkkoUaegjKJKWVmkLsTmV6B2YrJqJ2FF
BVlr3LRwVlrL5/CMMHYAmy6++qT6iemeiB0SdYGMkNH8mH64i1xS6xe4/l4Q5AuHBkwlAiZ91puk
FzrGUjFCfJMu+XtfjfSermQnUSQYWzAUb9OtSpWT7GgBTtKPhPVGJPkYzir73981mRJT0220Yuyf
eTm1oW5Fxsi4yPFobyzb1KCBGuWAYp8k9iOwss8er+GqclFHhXXNbBVbPKF01ap7Mx1gBa99XX4t
JBVAmKXtU34PRibb6kPPUMW90iYEmQwP3Kg3J2BRrSLqggqRma16EcthpTD1kWYq2GUEq8LN0ZF1
jsmXgQJ8wps4BnLijKredp+zVd22ymBPurNuUqDRtexO08Yilvmz/VYbGBY/AxkiI56KyZUAZZvT
5+jAsbB4nIbgPDXZGPJ9r/Wesxcgbz8yV3ITbt4oEoLR84CLiB1pdn0OJwkdOW5Rxlm0jRAUsYNB
Y/dQ4+ZU5Xc8N6KG8NLTBSrUznUWkQFJKrSxi2u9xhnePdieGWm7ck/LDS8qvhROynevmmt2Bk44
qSmXJOdxWFobiqQLKgeQ7GO1CQSBSYYMiEtJLQmwHnYWXgwVx/SgH/g9PNaxditNXcGkjVJo61K/
ljPLH3jpViG0+WKciRX+p+r2yvJzjQ4hnexOAPwYWNvnJM9/+CXVBSPiPujjTWnisPLFFgeKdTRm
Q9i2DI9n28GqPcDCXP1gIZXrI4GmiFRMI2uu/GtLlhC4TmGRJu2SVP3hvCZ4mok4Bwvhzhf9oFAS
oxhtVz29TgdxEnOlCUoaT0KmtcQn5neSc2A0TKvfL2TAoS64ZhZBi8UvijtNut1ZdBt07le2fFRB
H2UxbgVeOmM1nLyjXnTTRpEpOkEVWw+44LhNBNTpRzJtnUPYr5rTNKTEWQrMCkXFRSqspDQuz3oL
E4JX3yjgY9VAqOSZUHCh1l0GfID2W6H0JmmL0rthF0nChAoUriPEJ2XFYrzAguZhHj3rQUY+Zwaz
kvDx5Q40htAVc1KW9qsXUOIR86d7PvC0rpxbq5SaAzmCeIDOJvAgMCL48p4jBFpIqTtBvNkFoChr
YKNpUjaA+ZAK/Ii5+qShYadz5zZUXu/TjhBu9ciNBb1giW0OO6GTCKg73GIAmUx/9IgwOKMT4FWd
OIIpFMTX6QRvTRz7b1VCIHnKfd6mTGn6/p5uZ+1zbujByxgWB5+I2B8ukMblWQYPT6P8z50rpuJR
K4yqzCVkmq+KP7QR3BtMK4asWaPiEbxyaS1NnUh941kdT/pHt59Y0dkYWyrCY7iZG/1b/qfd4iRZ
CMCElwRaVHZBVFlGV8D7WKqgAea+VxldVgHs2rVmM0HJJFa+P554UhjPTTFMf060F3Ik7ih7tfDD
lz3ImxCdHjYaatgflJ0HTGTtVO83FkFFzbKez/6k9anDTiW0nSwF6sVj4/Kh9QP17WV1t7IZUuhy
0RJdRc3G3ow4san4cDRPux91rUOw2RwPKj7MuAJX69576Rx9Xs6WG+aLEkBHEE5/fFG88UOesRB5
P66opatydCFygmGA54hqW4WfdEqmgIh2Th7C3anAILUMdUd/7Ep1MWDfHOqBkV4f4Pd75vtW5mvp
JS4OZ5+fiizqDTKB1+qejROpRCNqx8VT1NK68pDOJKbQCBgK14H8do6YO5iw42cFhJfcZllh089h
s3MSilh8/0h55zMsNxFmU3rRzHr/rdefKjOoAhM/GYhngJzG1A6DXJ4r8hULI4GoUyCayqDrWMhF
MPjxRVYWJu4aiPlJ+a6Plf5CLe28VniD3FuJl1iWJG0U0Hw++FpjosLBQpyT1Rys+HiU0qRgmZOX
VCUuffZgAHMixRgTEyHy8EGsyjcUgXlrOJuv3v0X3BwvCfkDX4KYYWWLRkiHJ9F7Auqmk7t3ajAJ
kn3mOdSrM6faO5KSgt3gtSidG2AfUCN6LGQsMRXxuYQONFmTZqOBWNATwXU5/cbD1UGa+641WY4y
GRdns7vqvnKdy+sSbkkYzrVQUUeK+aojlOiOV71y79OBJIeTEm70OdrlkHZaOhZB9PgNzbjcZJx4
NFrlA509Av8JikEO+KNGaSvLR+ajJhHGLxp4fazfh7QwzndY1okui93S2BIKaImdTc+Wvss8zKT+
oiJYChAB2TEu+1NlOpA+cr0kYNwnnS8ffbMK9ElnPlCSqbeLtfgb7do89CKHYGeG//OOCGNqc+Cq
d60aeCLtRUf3hIBaoFLGG9YneDYqHidXXPZdyZmlQ5zObtNt+aCDd5GNuCx2ladNmSPjUl6yTVdj
Etcd26tseQAflLQ1B4T9Sn3qRiwg9mfkAvFHq59AS+CvWI/YiUxyvW+T+u/GwgLvOgQYCDw7NWAA
0kE1zatWoEfMy/BTvyIOXaMBlevbwmxmmp3XXXWkSyeUVYVmSSWvPgnQMNkCNG0sRV90c9q4XVGx
pHFLAEae9DdHDqtBFPD0/P/6kPDR1ds2ctRq0gRV+QxpSmGQAyEPRZKUUkw251phitgYBJCLXk/4
5JJ7ExRmT3Fgz6CcO/pAZU7/2eL23ZFDs/hkRNXGb+i/HMHBu6R9ESDjXdqhLe4YsMneCuAh0BQQ
QRkVGqEDPmGyxSy9WWkL9/fbXsSn2cUtxMufjy47ZK04O8yhiCMvnS/pLc58BTX5YdTQ6EOCfa5+
LKXPQDNMKio5Qm2QyZA7AHvFhrkK9MYrKyMp2xPFT5vpaeVsuTf7FRFGnqzBJ1cj1qniah41z+CW
BZyEaFD4T0ZOoGKwJPC71swaTd0g21KoPyLWkfFDxUDO4kDMfcZG9vzNLIRkcQFGju38BlOb+2GQ
VgrLiGTcAwKGZZAFLneh7AaKPsWoaCTztGQvBjW9lm2EnXetq4/RHe7ZNy2u1WN8ilANrEGP9VhH
DQ9Lfapi0UPAkYtc9ZICV3DSy4Bz4/WU4sohDmV66CL1GKvVsdBKPbXHFJh0pMf/WpMsjZw2PtJa
WlAWVKMGm8zOytH6avbc+XLXvaQ6AFuhwQXsm+QRcxEp2fYkg77HrOuDWT7Rfk4ST7mfgNsNfdN2
u7NHqDBrr1Xv0SiFs9DH0DxpnQg41yzLPDZt16BHtvt++fNfuZ7h1734aN1vy4rqttyqtIFXB29u
Qu2IMQdOqnukoRYQ6tg18IZoEEm3KPbkzHQPIGBBHcyDmCqk96i5ICFQ9DiF3uEj2hK1u7vpc8ig
NDerQKBWlVDpx6J+goQDgScfcsEPZwPWrdMRqDdSyYlxY3Bst0Nee4ZanWfspr2nRmJP7oUAq0QH
tBzG516OAlWS5mkczOu0O0jrfrxnsGUxbwIzcIjojf0rC32ovnFOP2LJwVRclTYoIlAab+eRyHd+
ecEG3Ror8MSfqmz+/BFcnOxIA6iapuw2MM8fmx5DcN9RsykYET0/ZVSF7qKZ2NK7VNP5RHPXmhkA
/V+/9GRAPpPmiROm4gLJkPTw9JVQEd+KVujSsjZcKZiNP5boUfsf0OdzIz6Eq5kyJpohFXBe8YkL
481L60E4JC0z0/uJyS9rdPJWgELaqNTGszajTFd1npW4rfdyN9IQ+n3Vc3fzo8P2oLLPDJMBeHLG
K0Hi6tiDPTtUzpxsZJoyxzXbTGFQM0xizVvyIQdqvCFOjn8ueY5IKEoqdggxs1kNN3ryVcTNZd58
uMwOR2fN90L0L0JE2fLMG7IIZp4vrv96t796IRzL1Vde0t/yNc/3ND5zKderhK4o/t3rJU5XOUWq
fdp1uw9bzqUksgyAQ+ATSWQEIASQaphbV+G4z+rIsQSM9oKWzDOZWQIsMzkHx63oEveSzBBIAOkD
bnEj530YEbRRpmEN2hi57L8uT0NePb14Tihu5foGaSumQmPIqW7I7oKyZoGewdT7f3ZxQHD4218X
rTcobjkdG9w1ZFeDMblccIyuAbKjoZmixG70/VukGzsdupxEBOFJ7rNon4a8fcR/6gRglPU8k378
IIGsQrOiB7MCZsGJx7fUlxOxCEcFqqAsT2d8MozABIcdkbSuQgcvtyL55N0B3rgJaAb9O5flheo9
bpNi0I3cEdDKIWQiRqECrW3kF3chOUfEwhogBaTs8kvrWsaMz+qLatmkiN6zsQtF8nSxEC2ODs2X
pcMS9HFyGaYcdmuFuW27pXphuzrevXSGgszJjTNLbbYCkqbhtFWXpZe0gSmo+WeuHEL+Z+EhsFjl
WwUH3MNeRBm2tX4AcrxfoZOdV2MkVy750C95lVIHZHhatGRpFtbG6sUTwbJrwi91ermsLlxU1S1u
0qHh6DJXHo9NsUpWLj8YJE/1TkIPSDVdAmtn3hDpXrJK7bPNQQoufQBsyhC5xkqoxURPxubnflfc
Sj43L91DVT9VomnGRMIsmRuM/efesAVj64TZsfqkrYBHA7b2jqt0lxunLaPfsqqDcZ+AmFAeUxEr
A4dug4AnlkLpp75YAU/A+vvZomzI9fUMA+qU2/gegwbpVVamntm7Nm6vdmsLHA1xdoSsIwqDQihw
6cYMY3JqFznydz78fuDLY71OkvJy9zmqCRZYLQZBjFefjhgQRLHQimQEjZ4CnWc4Bw7wdGWUuuE8
+BPOfUhWXMsgQoN4puzbUBmKrVSP9dZn4w43eIq7H0g0GmirtE67NogNkl5Htx1YQwCuf6j63Sw+
IA7dZtjSux8tNu0hsB1HkAyhYA8x7DnxT4oh1Nfy5Y1EY2CAlqqwABt31DRpF1g0gr341gYnB1gM
JCmxDnUzcE0OCiLyihadTCpBszbAmxg3B/6zlpV4zb4EThSiZQNTPtLCXUrjspFnsb94moVaL206
GBkjPtFStUVxSCs0dq/l98IzWU7Q7Jkg/VvU6SGgJvxhZ0jkEoPUhHNiiU+X44Y47TkgkvRitBfi
JaSQMezHBAxp1WdBUrY3aUBjBo4ffwCBEJs8OeFKPILQbVDiU+achLmnRxNHuFS37uPtsJReBxHZ
cGRbrlRLN0dmeG6AX6QeJRHsVY7i1mvy0x5EnaHpQDmM1ljo+3E+D2GKDP1zJYzN0AAXehoS8fps
PcXFQlic38FjxsKuWHVJ1H9NXHh/089zap1FGP9gViVLDOZwOeKPvFueS6Ya7uauuPyYB9B8LqjX
I7LneBFy61mM7shyRrzynlCafN0kEF3fgNhNxGuK4emTYKh+1+a9h2ZtpYJbhiqsElZ/IiV1bPAe
9ljhahfhq3VsrNsuUxVxyJpm8ZTyO3UQtYjjOtBQroc54gSylpFPxJG6I5qSMISz1LTA7H17w5or
Awf3+cxa5n+SKj8OezrwInEkJdDYrPn/74H0rYmoJa1DXrGJwZGVF/13vpmeE8ZeupJZkKE+J7vJ
GlYdWohMC1gf3l5AXEaYDYs1GxyT9Sg18dFvW4SS5d8XhwIuGrkMeK+NS7sSdWWcQjTJiVTDhFCe
KVF7svb1yfJY4ipq53H8StxubomyNHSpoOHreGivmM9g1RtcbGgT2jMsVCBZNrHwQTSSpf7K7Vxp
k2DyU9KxvPh0c9VbDqZiL4s8A4b1bclUkd9JsBRxc5ah2BEom7SFyPUPFpc7gtZfHBmJfqjvgI6s
EdnUbmAgsZx0iIRndmx8Jjst9+Qj4ds6KxmMrUNB8scq4H+EG09Bs26t/vfkmTeTmUIqy6xhRTGG
knOVcsOCG/uhm2bWqr2tT8/rapvkr1qpvR4mYUOmJo9J8K54h9zafSLD3gj3xnY/quSR7J7T7ASe
30KIOrdYGk0KEYEY0TKTsZNpYICyw8GRWGpjznal5AgqtxINXr4XghTgI7ohnWH2vCxTCzcnic2p
CC9qyvv3JD64gZASg9RsppgSlxNoDZ7fE73nVb+vQqV1cc7kpmzEMjS0n+q/EdyhIf3T74Vk6STf
AIKBW8o5EsyecyfNQBuBVLhgGPwYeBhDI1qNkFm6K4ji1UUHmMDZ38ogdOoBoVkyf2xZybra+Jes
2bKUM9//AjJAM1Z+kTz0U61ELal3ZJNjkPQqaxWNR82DMPR16Ltuiy5z6E8H+0o4fRF9QEmCYo1f
i+gPzc3y4hv4gkJLkiCXbVbsveko3VaHQrXnUgwlPPDm5kaM3lOdcBcR/OTu+Y9uFxSJpo3UQ3z+
uUZbWrlHIlJ/r61wDbm5SdaArTkz1gbgsGBGfF9hjfyzFmujhfjJXWpJTIDBo9dGRrKeVI02jEjv
cKmVhZIbZsGfi9EOP6DSYYvMaSeKkdD6kthoIgPrNXPnted20McXSLlumEma6ceHlWP7DT/4fr88
5wMcU1KQakhkmqYJ+ZmjBK60d2GbljJIcPvcgQhRo0olKSQFPJW/JStTn/Ykw6pH+7rtKI4m5Tdh
n7VedDUhZCQxB6q7wVoS1+A96D4yvBlpZ/ZK/jVKnhxnA7GCRP2ml5ZK62mgLIKIkrL4KwTUn8Tq
UZi6TU/JqEUS7of6V3O0QSzKoVWwlZ3j9J2q9PbLjzadIFCZVCScMx/GJO5zbGh2v9Nm5+soPUO7
nexrXrpRkhZJPijXIjoml7Xj9I6zDkbFNO49Nnh8Z5xzPFe6G4kgUaPNmYD2L0+mccIjaN2fMWTN
LfJl8V20VDqgdA5PmPFpY2WIPmWQxfuLRjV8xbQ0Eyth7nhPOP5oSFIB04KEIXsgx/cOj9tNuA5t
qBDeqOb6A48R3/S7i2AGQXd2dJBWDSOuSKZ5SzZE/iAb+TLaMEjJuYpuiuuX/BhRN8rTsgVDRfWY
seCThgRdb5W41MBPwhPDdATsQvvnes10Yw/HuwsaoBH4HNNLJKIx1YY2iwDsf/h7/wwKgmoZZGCs
bTd/fMgf6fn0b1waUmgRpo0Z5SfBEkbBSVEZZXvb8qIXa7RJAIlb7OJJOKHtLBtkN4GAL9Ixz8Lm
2nW1OeCaayd45pNd3NNSr7CqW88yq+Y/5UG0Kym/4CJBiolI2Uh9pB/dPkQsVDloV168oUvc0TZ/
8dIMDMfU/RhHqwI1d46NvYAm4slela09JiwpR9iqYsyfp5uUTZMYjY/tiMzx1Ozjpw0ZM3lmAnZE
xy+JUCwirUY21f1dx8/LlCkm9Ee3vNKw3ycOKlAH6ovWoA7HDwJB5ePt70MdYeCX2kVK/i0HvOhS
msWILesu/LIPM1VpivBztdWjETc7SC6Lmaf2TEyxS6wLz17xomTcdFtvgdX8NmP6PoBjIwKX5/DV
ciVQtBlghgDYNWnn2/9nfmwOWYbOTw/djW/QxoLNg2gxxtqH2hNkcYFBtVXtvCoM2GZkGQXQ0rz7
JKUeEtPfsmX4fA9lwVCCU0H5BvrScIN7hMg1LXu61HL+85CxHKar35B/Nvm5KYtDCvVI22i1DPyh
299p2p3gd8PZtoSugN3lSDaEIV3OlRydZY4SCqMcBZYh4PUbIf0IUhU/oMlJGI1GQyH0YfOGCQZV
1I7PQYblCeji7afaeFYkgohZufJzbmj6qtYyP6F2YvTWP/FkHKAXNqCwmjEqI6mIHAi5a2lLRX48
7Qhh4XtEqVOQ//PfFTN2prW4fWPgEL4X/p7Et9wLMulwQ7lU8k9JWGxv9vnziac4dRiCx6c7SxeI
wex2m6KIFrcyJhPijgP5Pw1L0Xh3bGyWjmioalEY4uID6T39BhN63DzsLZaIa5pUKNz+iJz3ezYM
rTQBlyjuODbIM+UYQckULwCifSbMd2DKMTMwPeeUZp9qSxCwT8QrcbGBgANhjyTj9nq9DHgnKPdh
e5KXNQbTArRdrM15gmnua6bsWiJElMvhGEUfHpdZC4zYFr9aVAsadreXWvjr+kHeAnc5oTK/BKGp
P6/3W2Mv7xOZu0iqyPR6XnBYNbJD+Dqw2RBexjvAafUTZBM1hAh+tCXVSK3UTUBLKyG0gPbUyLhW
mlGEThsXrnrY8BfsTAXmTaMk4OWwziasHh9QVX+81jd/OvIbrf10Y6qWheQVhoFKHIX8RWDP52aY
hVPPq4WIfQLlkbosse38S2JTY0uI0FRwUbA3fMk5QfdBLtSxxhqvWFPue5rOKsiGrwY08kjQOQgh
YifOtJPZdXbNQEhfmSSnQ7+6G4OHAyanohPLm+Kn2cxjZyAlGyUyqx/bQLFT6auBCEvq/sB5Ova1
2O+00lZ5QfznswcMOHJbvlwpAC4i8QbmM0hTAmpQ6UND5llWzSh9Tjb4c4/sy/vILRlggMu2WgkJ
ONOeBl6KJDvrGeFEJenlML86RaFtOQFaMADpKaOzTm0M64FN0M6pN70mBW6BSD4AFWrleTPYsUgV
tWJYUY/SXExag4x09U5xvzMiGKJI2pj1b33ozs4M2VBVfEaE6WPwMr63ndJLWtfQuoSq0f2KfeDI
uZNlPnZTnRtpVNoI9e7bQribEWzDqgBuTf1wQ7brrYmnUxLmhasxoqZAJcZfVZACZb8/cOQHa+fW
vSOEyDj7xrW4cOz10NtRi2L+Qk9HqWui4L7WYCDLzF5A4BEpgraj0J3Ljn++IVJHfKvRI9o91xbI
NndIVR/Xw3KWUzf8Fk7ItCLVhdyyGMveypeQmGPDcQ/tHTpW/Kyj4vmO5Q0F5qrH/ZMyLPWIneDf
GrQlO7M4+1J63Gj8z/SAq6lpU2Mv1YNDtUvU2TmURXTPjkhxCicAGqy18TKaf4WKhhkFGxVBfiM1
l8WTLzhVQDKY4QmugNC2Szy8PlOogvwgSoAHfGAxAE9YWSNBQdyb1o4giSnUiZkO611Ok/FwOZlW
x23Nn1Er3G2nGoqMMsA7Dk6R2iNPfr07TBqgxD47hUEPAnhcFecrVWtZpmfI34ZxLSbJi5BTQmXt
CT8CUUFI13ty/jo9w2hrsMq356MOgq4a0nZp+gX0/xcY3z2nHaAicnUbe0FWwfcHdTGR2f9CBB95
ENbJJTfrjCQZuq05O6IanvN6Po6raDowFgWQX+elH5VmLqgbiJjMDWeyGohO5ta+yvlDWx2MLSRO
pVEKf9OA8/5NhFVxIGgAVvAPadHe+XO/SJFIEdq5sUmMqR/wf30fhDT9TvXanQvjNjQtrStMyx1N
mt3ZA3XdnBh840f/ya5RINwsMWnauQPTLFHo/3DPTbnLxrqVnxyLrjTXNrucJj8bwMACgZp5IFxP
o7zXUm+JRbST5MoAwxgILDfL2V1P5EAp64BaNH1d+otcPyopnLTu+seLByWfFll4amaRMhbkl9bg
euwmNfVjXC2mE8Rh+vWQ1NKiYRAdzURF1s6UYZIJEgeRyDjCJxQvbVjV6g8NA75egpMK5bdcRd26
ieDPFcB6bKTmp8lW/Jwgka0KmBk/6UTQOMmlaDxmDRtvCIBKFXnwCurHvR0ujZiayhwAnGn080/1
PGBISDaMhMwIhbytk7A7Raaw3Db+Z647KHxDiqxy03iSZRiIv+YItTvEQ6Lfg8roFrgGYjiG9pfW
HQHl8ukcbW7D8M7WN0xyT2AkpPkFB8duTMUVCj8BC2DhyTExfuDcY96MO4HocrOtWnjPz+jA0Ac4
dEDXmdS7tw2lGTmqJ0Fs39rY6jdFedMyj1Ay/CLQjZqyfdjqYAUnsYYr6Qakma/WNhBRDNFIPuXA
tuFFRjxwgyO6X4GnyrETjyqy4m66bwOqP20OWfIw3kIwhmCKCj8ofohXGj5FQwx3Xsrfz+1Ot/zp
Z/3RIxB2K86oe09X58mKtoLQ1aj4sbj34Wmu/02UhsHrCHJMQiSlGTGqdt7L45FjIuDF0IYIg6XS
d96fVVks9kKa5O8hrrHxSMGza1CCbdKAQxtZb0gpbMTFEhDdUZevbEqiSgzbl7XV6NucO4P6eLIF
ReFSByoeVwlCt/FvyN+ngTs1tsHcyvpnR7gFYvrlbeTtud0TIeXEYB0mYcpw4/YKqaqvJm4WePuW
o5kG6SwNUkkhD3hGP2XpOCNwP/IyQIkcXv9R/SZlTvmXMb9lBM7LeFG6UGLInSFzKQZrblLa9I6g
E0lPKQxWk0wYI13IjazyYvFlexU9wiWVOEpAG8cWhz+19Wog7ciMvma51BLTdP6TriC9ux07f336
wKWKLlzl3hRhcgfhLQDvDMbxsxmoMfy9dRA/Y+e6YKNkXrqiwgfjHbcbauhEp7qUrR2ZcjjCbwAA
56gU2Vres1L+DyuaNG7eq0jEBfbtL30D3lJVGyqdgwcmEZir5Ymdfg+YyocQe2qydec+GsGF9pJe
/3Z096VAH5ETh7IeaOe2/ef2rdZdPUdU0t1wGtEwBgqQmrq8nUW2ykj9NG8YLpTOJdupv2A6akOa
pp2ycCbybAp0oFoRLe007K5UVP9ZER1A9fOEgAX2gdIefueU69kX3WTpQiZN/binjGZvY9bk2TZ2
nciIg4nRi1ggLFFgNdLGDHTae2V4b5avdOh9zLNGvbfXBrSKddK9G/GqYQLlLPjVLJvYfdX+61J5
nQCbVjZ9/c4pFc8xtQ/vc8E5Ar9k0htXP1EzyhfAo1tipjyGl2lLKyA4wqzMkBCh1Zmd+zubWgHA
gKUOm6RaU1Y1u+wqgJhIvaUd/7cz9qeiLpfUeQjFgTt8jX3Nv406Hk/aVmIw4paSkT4WOsbfHjMj
6A6XOMvW73nt3nurmj/nWo/N2zUXnoC9S40cJTIIFjpgrScnKWqxWpMwrL3A5ZgbZVqh+AGv2QnJ
l2316vysQoyqHUzrbWPNwf9GWAq8S/btQxUO2fTt3Vi2TaKlIG+5GC96uI+ncoY2kybQs6e8N0eV
Gq+R11tEnb5GKZPV7CuNLBDnLD3UHHVTjzI3Qyk+BVzY+2W2qxRdbv61jM18BQLyPSnx0al39wRV
Hgx7PTJet8jNppO9BdlrwK3hCt4zJ4PyfFYn95iMEnRaUxI6QDO0z+x4ZJ9Ov1ru6vKv17WotkkE
4s2KMHuW7wbyP3n4Slulf3etfiwFWeZKrS0yy3T5oXKJqLylkiH3e/l9q+8TeAgVEO2YMgHc8Slj
M2iwRIARBeDYBmFXmXZ6TkZXuePX1MyGiFksiTieBoZxPP42EotFzfUIm7W1WLIO4Bn99ZsecEdR
IMgQ16VkqWqqd3JtVwavnO+uF+dPNcUAA/t0M1vBJwUZssnAdpzpPX+XC/OSbyaOleXl2o1RjN9T
2MdCI/1KwlRhlD+oTCAkAEqp2FMuLyvMnXQKK8l7B3EhXYSYDHFCNRMXejYJsud2HPb3cZgEaYOn
ISWWWjvqLpbxbBLzF2Oe4SHOEOpYkeHSiZq+dy6hA0Vgz93hGBcEC/SgDzkyK7JcQJ0sx+ANqD8q
P83yP1N8XetkZzJ6qtg8PotDo97eTYdjLX4RK76RTknrmZKLg2RUycChP+NuCOvwUGs3/wyYIZnt
9c/FaOZSYk52TE/QEFZCECfb94Hc03r5mSR2Ybrds3nRTzTMXhEmZWlrRS0TEezxjbhCl813Cr6+
oYaLi0Mw0eMOGjCPoPyvgqHLwF25rwpAtH6Pyzj0e2QvlitHeQgEozjx21rbVMRks5Hf78lwgP6d
/OFUeBA18Zc2opaKxEbYIjU4MUAyevFqyRad+zlvki/ixF2+/tJGspcGXFpLBCrxW8DcOQERqtJ4
RDsjs7WzVAuxwxlVX3Ln3eSc//ANX/jrg3X5jnQtZK1jNRZ9rt1c6J60lsNZ5TMu92Eg0NLdYz+g
A4msixleb74jYXI9DvbMSd7bGpmfrPEVuSr+RFx7FAZVmULiOct/wd4BnyOvj5yBcxDScd2xVoEl
UNDv/ic33QO0VURlTiujLqQYPlHY9P0dUEcMGDatEb2JgIyMVQfzdfVD8LCwwN1C/7DUS7yOr5NC
lNhu4YTq2Iq0otkBH82VgnI/KRAUolkpFiVah3eMMgMxQK5Jg7UaJqGLgkuEVLzaFFzSeFyHvutR
TSYn7CnH/QQndRbcX6ARN+YtNEdfE+S7ollWMs/BLUV+xS/SCdwW7eUMEZyr+Z8XmIUgvGwBlLa/
YVNKReJdl63sAPBxJG9hQ4m5BnypKktkXxuAgaOtC2Zmlz4uAFoZSxn0SGFk3wfR/OVQBHtt0hq6
Vf8Vhm6xAWvHawlYDVED0pPLsMMVwGQ+AxyYWmAPjT7czs+HhyGyNVO5EmDvhF+Sbf77ERxUB5s+
uOlgI8cY9kG+9GBGztg9LoMK/rLK4u6e6NvrYeUDr8ji+boOZMnPbrtexJ4fIuQu6ez787DzyxEI
+e2z7nakRWWqdHwMsfs2e+OHYtMOxVbinlKoOVDas0nHDBrvwIuqBkuesMx8znUoBSX41X647Q/E
+t8ZsGs6411ZZaco3hZqO/pwopvoU98cVCbBzXW+m/qN0C0ktN4eiEanluyTaGUm7MuJJRznMi/G
KC/Sy+DlyapgSUNIG3VX24gVl3LIBefKBn+ur8JS3dUlBzQieNoa0B+VAGEJatTGm8EUUyXUlpLw
F28IYecjzoNpA+L984Bt3/dQnNOP9BvWdwUJ5MbyDBPnpa+97OpGIHpBHz3fPXuCK4zKconP186y
nOHz3N4CBc2+CkhDog7W7ZZjahVWJ2MuXmb1+1Zqd8Xl82yzg3/sBTqWnhDbnjUrmVVOUjT5o63/
JEqYgRJ9dUfKRL30z6v6J07B37rdllqpDaoOZzSeYyR7ZWrzsQCXo+zxsM12sZdORkyVsuPMImao
8pK2vg2bEPu19ni0+q0rntQG1pGf09JAf7nue/WWrtAuN/vVipm0AHhUlw/aW+BYtJA3yMS/NRD1
03JckZ65RgTfZBhVJwUbr81dFvrkQQGcaEBT029iy1u1Wo7zUifPrN+uAfFr5LZW/+8GMqXquP0l
EoIrBfaLmEyDG2S4gbE1osPNGdkEULxuS97DINxL8LCCtR+sPOHRzmdSIDtZhdxMSIvkUP69BNeY
+2V83ZC8wS3vNqWB6Lk5MbBLK0AS3xzS6Pvu/mj8dWS2b6Adu8MpilmhzcZ8UF6t0Jf+gU4JRBqx
2tooNMYxULNAN8cSr+/xUy2IHo4XnRLmgh8JF/UnscbsQCKqLis+P039FtR2/KwVYbQj36JR5iKa
/dF7wBWsaPtTPx8Xb0TZlH/m4t0J/pe+eJfwKIVNt1hh80CPMbcb6C4NlnuqNKBqZrXBTOkrIIOW
gomldm95TjxULzb7Pot2yuT7wqCFoiBFqXPqEpt5uIK9/XZIomUnT/Ti9MX4e4uTWNuhD5abpzSH
ZfECa+dXnHZclBWyo/poLb8w1Oh6EhsVlbqrLWrd5ZpIS9Xt6FapqldwYlw65MtAvLngnd+x4SLt
U+sEGc8GCns957ANyHOgZ20hREjrZReF/cxyWkS3SDu521Rweze1Pq8rfgeQTT2JC/g1FJD02/Vb
s01QS9uQPawxcDMMwl4ykrSGWH6aVLJL2NxzLWRigbCzu4vjjy3A1irLMmJYv76DJJyqHWn7voNH
s4nlCqbDo9HKhuGH9Ars73wXysHYGJ250iwz36f6bDJzXEmcwjRTGNc4JR/hzrVA8QJVXKKDbw5R
B2Wa0ps3aJQZy9ElaRJc5MqwCKXZ2niyIh/cGUC4l8uMK6oV8SXxRhtEhJC5kEc0xw5/iB8tvE8D
HvmnIVmrMeiWYKGtFrNtQT0xezrKVi+0SEFUxgWwW4S/89mDjk45qSJDGgBGUsgmQFmLVxW0u8/y
kUZr9pJiiZyYrrgwGi/hMT5T3KO/s5mGp5sxl2niGRjMsMKW+nS57dxmH3AQwY5Jaai0mU6sXWWc
ng7Vtu4GeX3Lsys6w2Nmu6vpjS6pqL6RjYXshWCU60R/vlYZJ3WmTe1HBShf4iZdLkqTETCQulDJ
xAyIghBba6FmflJ6jLZv2Sw0bsI1wjhGy77z0t3s2maSjYPt3LKwhlT+j6c8Zmr52hG3Tp7wyj8Z
/pyvoFnB0DlpZIkj2rbQU9FLwC78r0tLNCK5Lz87r4kgc24jfTHTPtFxsNJFuZ1l3i1zuPXFJSrA
diQpvxUyd7w4FLM66H/GwCR/A1NhAFmPoy+h1bT0ctv5O/XG/8wIy5bOmjkS9MNVq7HnVrmf+XZg
v7ZWi0Io2Uryz/WB17vbF+04Te3f1UvdD7s3xZmXOdycJNtJebk28fWRO4sV5PM75QAncNfLFfQK
/IDBFFGyB+CP97VB4uwXX37MjWtTK7oaZlW//+MFBO+1wlD4R9sHUaHgLEBIc6J2MoFQJXNTqtPb
RZ/aPr6c9Ir4cdOGeay1N09Z9mI7QWop0Ws5d2Kgxfj+yVLAzW0/4sG5nH8c3L6Gj582En/tgWGe
l3Z1zXFV0QGQf+N7YgCGzQlh8GYT/9ywwPVFbHv4JshadeljIhHm3U0Dq6Rfy3ZmG99qPpyR+NmI
esDiM4KeAOiS5Xh5cwDYKk5P6j2epEG3+bcY2ao514lT7E0aVTYCGq/JPS1NoU7tOntWLm6PGAGK
Ghp4h/PSt/gjggxwoXIlR6XtxQrIb1FOHUFuGRzuJOiYskNEk246zHyT2JaHw3CGJE2fsW8B3ebE
eqMb6dw+8xbpnl8W6/R/W1snhW5xwx6s9OPRSH7+7ZLJXRm6SrWyboAmcwXuVgUsOX9fsYvjTohr
eW+MgtMLpV+j4OlHh/8TAXoJZcfPPRLz69DGgFIk1IkdHGxu50wOBGzM5BoFy/MmsJTS3tZYcvTM
t4Xdfs+Vl/xedB7IdOkCi5WMeAH87lJngeFKluW12wb9k2AK+ha+Du1sYuW0vH3sVPZadqu5iMNc
pw2RD9ZtsXSnkB0p2Nk24Sf7lczkKVxVyveThAvhsDMstmDVOxXhTZ1uy6T+GASJxmqBjpZm+UUJ
KOs5L9tY9njtAPb3xGqjS4xBcgNZfkHdGnB94Gs0S+D8aJk0we+xeeT8P8E3C4nuTnBYdozDuIsa
ypziHO+n8z0/Zg2IOJ3rhdM2rUebFGJPuq9lY2NTx6CaDRWOXwj1MK4Dn+v9Q8waOLtSQRdURx7u
ovllg4bgxjZMdosrIbef1eIkSutAeeah3VN9fx8jaf0JMEnFi4C27k8cOqjul3ELiYc/kPllhDKO
eWSveV8R2CYqGcRJT6m23q7dKXFoC+jm+zDsbbNJTwM92DYPHv0PYd9uvZO9a0EXNfX0Oa0dyE/j
clEzSLscF5D6IBOgXRU2+UcrSis6LeA3gp0b5K3ITlX3zj6oqkUGrzdeSjzTFtnerjWurlKaOcHD
U7q3ehdDWZFinEWVpF2UTB+R5qYaosvHHQQ3PUNVHMuKhbmRLScQjOntwG/XXXdEDZ67A01DOPne
CIerJXYIzmqsyUpC++f56yAiiJ59XKLODyhR963LC3L1Hx+5jbXFQmN+ZZ8zAYpfi9wccNd8cJx+
2wpcjWRw2wMnCaX1WR4OTcyly9HYCtKuGrJBUA9y01C3Vra/mbyL+D2YwhR3+Ce04Gz0DnqTDTSw
1/slRg8oDYGG2hr1kPDagbsxh8lwwVz374sMOCgnu+5wljbRNKNjNMifwxMrj3qpDDjALsBvE+88
iIghxLOl4hd2bshz60v/7BDBgkdo9AB4XnXZDh9nn3af+dMUV5DTdkUXT8JDZzP8i3ZjlIPJfsR7
x7hDlLcGlyAnQoEWYkBse94UXBdgELGds6P9kQO6RwU9qm17G5/0zrxGLy/TIOB8u9dOYLjG7Q7i
wnGr3ptKOk7xCyVcp+HdmIiaPiRR992bfVzXQulXXU0XE3Ff1+r/D85rJaf30IWyDarIe8NwSjNs
lJXpiKv6BrdiwgJpfjlSQrK57yJ1UfPJKrveBIVHEeZeAC5LseF26hsZX35fk5T0yvKxwysRpLQs
FW5VT2HQiF2kjdFwuKeQbWvDG3QKblF6hKBPqH3Al7suvL7kR2wLOo3yQml7AxDqUvX/eBRyHaVD
FyxqNHTIyC1XkLx2EYM0BzkDLx5OTH4CevZc8HzgXN0Qc47qj6AQ06kyqhdb6J4ULU63JU/0Lp1W
aIBFy+yBsbEeE/8j08TVH1QfvEV1+A9OYea3wjYeYdCOFZICAs5p4FSOW14YgWh2wNfqAB67I+S5
+UsrMUbJGWrT1wsU0Ngv0QJ/IkRg9cKI2hyxIpcFtaZUQSIwV/cL8DPuwjjVNjaIu19A/MKdS/8j
kS0w6D6LYuOOY1oHHhH4G0bV8y8R5fV5JKJ1zIcFrmc2fln4r5kFQ+cBIv1lxCTsK1K201ZUZQnZ
l0ipSB8ee+V0k5psAghjxmemhvALyiO4DI4ltNgH72vVoT2BB+yEZK8MxGlI1t9iidHXUo0rhw8u
oBoPwcd0lBCgN5ln8yaHRTSGmPqM7Gfs0ojpJ2S92mhcv1+06Xen02FdbJKtzLCvfPeK2IoCidQY
nci8cmacbTcQTZsOwPYdcM4/HDDgK2BxwRVpiXspPWPlPUitg4Em2SYgntCefChhzSonnREY4cV/
KOQdktj9z9D8Oajd9TQ9HiNOmoLpbFe8HhtwtOTmtTkTzPAFyU8WzMXb3GeVvKHk2CLoE64ewlRl
leAf1p+uas2crhWa6dt2RhP9PphX0q5khbuf+ydw0H9UGt9nhjYkwB+nsKM7weysN8Dg82YuDIvm
sd5wWYUzYCDjZ2hG89akUGh43TdsUlVWvXFuBWr3jMt7DcG+filYPwiZ6t8L3ZZNxjWBZ5OTV29f
23+Rt2gDskYA63mHZC5ZBdZpd/AUSP6xCzBgrnRwPoIvOx410UhASOD1cElQDKTBtS12SRPK/IGA
chIhOEplJdU0VJlIGH4T1/TVN4BHjQX4Q/lSzRRMxsl8vM2ify+D2qt0i8DoXbDbXDQm0M0pzKMT
/OX6achiDGt/ujaZ1OfJwMH67zD7YjSF/HA4FLdDlxA7y9FgREkM8scevDyBoHLefOGi8o11pEAz
8clDq1w4LHzy6V6tXAl/8Otwbbu/U494GMzSR8PYHxtdbNF6W7CzrX4rt+4cK6dPHiat/uasyEQj
+I37gAp2KUGMLIA0+4Eth8jpHq0LpKmkKycdGOFb3bA7lAZiYyTFLHeKZZjEVpZDxxdNsXjGiy/N
Wag6Ghq0OXCRMx4of6IFoNKoe4pngJMNy1ZxwJQEbm+OqEJ/CHY2nb1JugG5Udk88/hRuZwUQce+
SCB2eU1h70sa2lhJihncLFxyfmib/lNpAPuDv2LAglazHTpCYuGHdmqp7xw+b1FG00PcQigPEEcF
+aRZJoDwb5jCwmKKaYhw6/MAaFLSPm0Wqnlx+Qs6Yovy+adNXahPgGfZusUBHYctdSb/Z1vrZdim
aBaHyv6DuAilvQKSVMccIMeM3TcGTRrDi/BAChCscgsMARp6r0lqzzMG+AwG9QdMo+fS/VpXz1Fx
3bxg3aodz2uBb5w96wlsQoMDj2sgtSc+/Rmo7DtHJJ92Szf0/GGaTfX1iTPnR5GJhQRwkXg81EfW
3BtVOmVGNvyYXEu+huVWfjDzJgv5Ib1gQCmnYbN0oLH9Kw1VmcUXSDvylRHi6S/TQgIVTRcY26zK
IMIbZna8Ef2E614R0vFc+6DiOKcjhvKMksCX5rAPZXkARnhRo8YXzcv+AhHtEp+kvWKqp22F3zUr
V/4KJzaMdBfpk53ZgG2B0bleRIfZajrdoJPqabSOcM/3T5uIA1HyEyCKiFM4/LXtu4wksZOBT89Q
kwhWtPS+Lber951eV9Vfy0SO+KJ5/Jx+FkkDq+yogaSIoHeWqlceS+Jv8BwTmmIu7vF3cE4WdWIr
ltbUHcuaYrgDGtfQdtakhag2F0x6FPY+Nj0zzo9da4GR9hxhRGG9HhAFaIE9DRQqPzXsbo2la6rR
eiCgsdMWo6UdChH0/a47crlPT1yrmlArzAKRlRmw1mxobMJAOrQOhYTz9cXuSDoTDUKwAe104Ers
3Uoj6IUwU12TXpM0yuK4d9wTUyljifyNnJwl9DS8FQtEvNuC87Mr80Qxv7JdlaQsFKbCL0y+6sU7
i5cWYJDfedbEv1Wu2QXNH798VUKf5TdJx5/gxn1R5yHR5dD1b1sh7IfGrmYfTDl7UhncqDxS628O
dv6pvDn3TqxGkzhRmIgPiebq/VVUXp5z6uW3RJLeOh0tkv5hgKWoWglx6KYHbHsgkpjz1yPmmzqR
RHuLSnXr4MgQoKS9fLMDnisf5Cq8lH7K3jWVef2NEdiBWHhxkB6XcHoP8jDGVfvD0DNSXNWLLgB4
6YugbmUEPAsRDi2v+muus5EpSQ947UqMkhzjfeGkDdQ+DQ1oiPM73s+St3FNmfLPe88caDrPSZ/d
gC/epmr0CYtmlSXC+C2MyLE8ElvwBlXGspPSluSfpKhxRRvnQlIUyfzJ89EEZ50ANnnh+v7JNKeB
ZwbHY3XIk2GC3twARNX+5TVbKFFqU5BP+15z1n4RCQSfy0ARHt1ayHgcveRwzPStLrBIjP3FE8T3
XiSxFmvkhO1L5BATOcsOvIUpoGLv9uWVRCrbaTpnFoqNH4eJcJYx0DKhBjFa1iM0XtUo1LrpYA+/
R9daFX1bWGEnImVeRFBCOu9/1XuWkExh8a22flzuqyTG2sV6IrV6GY3KrLX385r7njNnxTTIclDb
t4kYgireCUaCFI3UwlpJkLb5QYWPLJuMzBKD5yzA2WchsV8sQRXwfSxc3yvMeoKrJUEpyDskHmOS
hxTBaMNcNAn31KRvqONy2DZtELXSbOm/6XP8UFgN8szgUPiDGu+PlCtOrTL/f2g9fk2c3wkJxBdV
BfPg6W20JFPJS821MKnysanSPwhlE2P6ehIpVIuGR6Htp5M1TDGKe/Gx/8DK+wjmokf017AwZ3ux
9Z8YbsztkZUmG4N7Vg3uZD3Cxr6Eemdg5IiKyj65It+77jNfzAJl43ZVBXrUmdb50aALDCIGNsaw
wB+M4jTIhZcE2K2wVCnCq4ayuzr8gRuWDGn+Jmngx23OMenNzLIgxpC94LFwsleDbymTBmmpajMw
QHQNn+5xj5qSvqGX3oypUAiZJmBJjD2ww+plSxibDkTgYF8W6VotkVDNVk4WVnG6PQVz95eSaAwu
FeANTxuUO9USIxiMK9OdKMKtP9iKMtDih3Ute/ca4dHKyj/NoKasR4/Nmr81nJXfaQ6vbVSPzq4i
Y7vm9R5rFfWFTrnDH6rxjqfphpJaZ+bz82eLbLUs1hs86+UStLr8aRpr8ufgaueRBojEMtJD9owi
6RpUO2ghT48QGNOlhqHl0mBCvBBOHdx0kIo5mTXskrMwHO3KBGS43B0zWBp57lcvUfi6H+Bmq1Bi
LOEzEVSdWj8ArMdmtiEd7jErgnHB2hJbBkyLEBaTPJLr6oCPy832Byafto2OamrRy6MK1G9o196a
ycgQNTwm/Af2biWmLkM9j3s3LVraiQpPaGC8i1Ge72FXNSQ7LfReBsrdA5SwxwbOytIExwFwB0de
B0hYxmMDVPh12fAGCtJyP4bVtUxledO6H6reFEpnunPiEh/x67+yNvg3AItkM5tqKLYAHM43Aw3u
Inm7iieUwWpjTGwRwE6nBJYFtdi1oe/SfHl6vd1SRwOuP0IgoEYW3E5MPNn8OCVgJ3NMv3+Hxbgr
QSCbko/nHplCNQ3Rz3PtnrB2wg8FslHecQgQHnEbdHOI8/6bCdsPG7tvu8aB1jBBJ03tSbCzk2CA
gm+29iMpx+ij8UtZkM5B2qxZTsjvhtCVH+rPErbegXXIIuDYBxWRotfdUNsIq/HXVH2kTl44dHnU
lhOHtZLteCEAfoO5OYCwkpfNZbKQJTlvo9XVh4EoACegz3BOKt34PSLPdHjKHEXiNtF2KY0VevCI
+c8UF/4u6ZeuXiwp9MAzqFE2t+pedgbl0IHSto1ZjnoPCQZXweuYCDO+2PD7p1q9EO4l3R7OrQ6O
pfJ+8vbOoJc2KIQ2OSDeqxQyeoFLb2oYEe4L6pJb3zgBOoRcoJqgfm1kTIm1emfTU0YT4RiA+uuq
YSgEofhs2b9ADFsACXc3R5AHwwThV4lCtsY5N2DD6/no5HC4Lel0WaOxvhBNtqF7ze/4gOoLCCZr
d88/BLpZnxynBHZ9T7E4195EBYDM7lPue17YXgWI9XeLeZHZSCQvpWBSxPBaGwOnRZFqcU3c1z3w
A3kg3nUXpNYhHuCVSceC6IJqX9QNz8d+rJTcNo4/TeNmCav+wD+mgSff5+57WikrNS029ea5Is4D
/jV9BGkP4IHx9+nQwaKuU3eogRV31lDC0Vz8ArM5KP17AUg4q92SCZ+8O2zbyi2Bq3YlWRNbQmCf
jT6SkEGP0LP6MzNkiifG8aPy5/zI/Vua78kQltRdNzJv88PVvSE8PFXieoxnrxGUSVI7eFOk2XID
z2ZOxYSTMgesH/eiSLt0ZTo7emfIpz9+p5ONqL6feRwFBkv6hQeho1kmUiyf+kaRhQuF8Mj7Nnr/
pH2EXI2WA+YRPVaMXs/yRENDarG1rhpA2ngPRU1Nij1nh+ylvYs6eqS252YiTYDcK6EL5h3atUe1
y8GiRsbQ8QIcqGHyNivImByh7Oy8PUV+d3Tqlwfk1sqgPCZYoK00vXJGcwlazaZHifXxBntQ7ngd
fm11RyIV5UhMObaLEbKqC4c9LkXvmVVCOuGHUlAnpI0o+Hs3/Q8qxo5cgvwNmdVhFOknjWhNDjOS
V+JfHXY1Ydl3m8FC1uMsFIKmIfZ2xfbdo5K9Sk5UxD1CrxTm1l/ayaHHvipe3n6ycKaeulYTJ8bD
J/yzKA/z+2GND8CZykvQw9TRZ1666qZukykKUCn/jC/nLbQ12AWaBtV7Y9/4CV3QFdCdZ/T4LQor
7Hy7EfsVpl0y2XvYJP4gpJbP8BtIn3zCiNfQ1D4VC/zfpEjrek12gX57ByJ4I65+Q5FA7USKpjK9
okUMWXpG5DLINeLROYIpi5TCnUq/RDghS1fppBX0yxN2I/GpM2AXSfuzzbRV+/doAg87pSGwDGut
dOLh/Z+f366FaA7cw62F8J2OPNQIGmQuy/C+5krZailVOPGcVmRDNcy/VIINfDihQTgd/xmtLVvY
YEiRJuVJSQ2l72NCEPULAqs/Ey6zIBtdA40fgmyC4trS0LDuucSB3SNN00urIDkJFMxYKtWXO879
+BdOmwDlyVZ6VjKqMjtrlrAwNuOiodEnrqhZn/lvHsguenAt5FKKuZgKt9o4RHVYwZB/1/hmySi3
Fpc8JxZGjkeWZ2lK+6ewo+9lXTyezNYlqnorK/vNxg9bMiW3FGsVSUw8JEnxxig6WrbrnC7461Zt
fYp0oBbMdWVNrwRZ8Nt99aY0aiJ22OjNlPEWTtYc/I+1auibIPxvcYmLSLdpZmvtF+SESwWcPBGB
VbKoJdQ9APlvsq/5XuHnmKEu4a/aFy149eASQ3tUi7cLnVKz2w3nnGPzfgprw2Yld6kVsQt0rxPc
GI7d0Uj8cwDo14V4Ipno2Wm3TMNujDBSCaFuDg5PZV5WmzSPG3VX4cVD+jCjexUTnHR73FnscupT
yFoo/yGuUCyq9it15BTdYhZDiCQhi1BZkspNMf7TsvuK2yI4fW2QiTHgcnu3IVEj35Yfin70mrFf
jt6RWQRsuI1aI3IT5/XCKoyKs8CHwcD2PpXUSruTcqKupv8cPmuFnXuqHdUDlA07iS1nWCE0Mx79
PFszmD2de2qf4E8dlFC8Oa3sWSpygtzGPEw6lEYH2Cq3e4RsYAODC01wRna8dqXFrkXVUzWPaIvL
TUXf6mYQF8X0eGub4yBr3CypPBIgTsDRM/PeWSFzMCr0Jt4+dTKBKk5niIcOIQVNSlpFNwnBfftq
dXQBdY8tECTkvfMdh8AGHMyaces3O54PZ91cTa3LGwb9MJUo3YOuIMf1JMHU57BOMrLTPe5iHEOK
h9QnROB1FA+BrrWrE+mUq4cWITVr+XiTiOLnmevyvo/Af7ywaFWJRI5FLbGc9YUtQzoq9uulpY8Y
KQiOPqsEka98Jn0nPpTKmyIq8CDP+/mCK3k795+BeV9Q1ZzJx+Js1ESYv3YPUasZejlQAmd8aPkQ
zU44tS1jlYUDfAOEwXMKPirzhDceKLWp0iLISP8hvd/RO2XS7mERq0pDvEAG0Elwj/wuPSIXzDry
9iL2T+JqyaVTbXy/zJh58ZD+oeRlt1/IGzQt6nlTnNw0K/iyRb8iizNwG0jiM8+u81zrUHb5kGQx
3il+wPAkO7Om29xMEOyaM7fHU09btv3BF+BaRV9ebnYGivFBtwkQgI+yuNeM2IaprNd6tFInMs4Z
LLavXXG0Adl5n19RLhxF9/HDLQZpgQlNFzTw0qzt7X/fymeeypr/gsU7kZcbKeMYkntSFjJlnuqj
QXKUmQfOcyHLf+3g/ZuIPDWaNfCZlPNF3vwebR/ffzh2ldKfizBHScd1a9K2XYyuOp1uhA75kj1Z
zQLI81w7Vv+efRbxbtmOXTDxemuTbV4MhESriHr6aasZB+w5xVNA6F2/9QmV0HTy+OILIATOxLwN
EHhrXS5cWNrKBmZSPFYAomauq6LcCPDoKlpNflzBdRVGgtOC86z58SCFOy5FLs591mYekCYENlmf
n9z+9uTw0TLzljyZ45qxQTElMcF9BViEZAY6Cf2Hd7nTQ1/mlgxladoP6+gu26Zi2ihukNDwAYzJ
gHRf4q4wdqnwp+fH41f+L/o4Y5eO1rsXzPlAFWj3sWZKGyQS6WJA/ukU/NzOwPXmFGukDoJfHatL
zfDyTH296Bw5+SuUf2PXF7aed+WkujwSmngzZx4FFkenhQ8SsWMsaP3ppK36UbOw8cowIeShjPaO
z5mU/aFsl3SNWx5jsE55qvjpbDSAWy/H1l2ioWQeocLhmKR1t86REr8iho6YEG4TXNxfousRgbEY
J0zq/OITwExSu7TnVEFq5B1UZ1yW9BKDFSakYRHFbc9SqhTPIORFhOJh8iYsJp1niECNC4rwA2HM
Kv8Tcs/52D0jQc8PbDPlQrWtG+3T/5CyE78aKy17xxZu7wxZvtXDtGes+GGmRYdA724BIbVv97Od
XMvsR8+ebmMFCnkCsbvm+8JLn/vyWHIVbBTc06763us3XZyTvEI/ogBTwIBB9nuXq1tYvPK/Jnnn
554cm6uwPIsjt/kbhp9+VrbwofzWb+bpH0xpkC5+QikymQZYDDUFNGe+9DZNbRlt7bsLbU364OK6
7VXO/1RZOf2prcHj6EgqKEH3ZErlqG0mKQYXGdfRAN5j4ORRipReEHq2hrB5LYIF8PyWmTVBBS49
ECd3+bNqn5AFr5YwGZO+Qh1r82Sujk2fgkQNqgGx8BClMbOgJhufvq3n1rq6xKt222B+SG18wgy9
ri/2OSMyZrC1DkcMkhChuWTWAV0ZQd8Xe4qXxXEp+SA0yhWgpPI13/3goFi5UptB9qwXjzJw7bZ9
k3YxyfQiPLDSHHPeRCi+a8yGHjblOJ88RZ5Iw9VCKKhdf4pq3WTmwAYSuk3N0/ii9dhKZQEF388E
keVE0NMns2I5EW8Kex5DKZZ/J0FPFgELwZYGMMiY0I7ovwfIfpeGpNPTTIQIQsffWUF+22XymlkV
ttzwqquOaYR21jpfk3/9a+Lbqx6Cx99sbPy7kJCQ5tPVVsVdz7854+kRQ7I2tK0lgF8487e6A0y+
4zpyrTECVNlkP8PG5CQfDo8mN7BNzI16VwIo5+6MNllRcMj40UpV1QoR/VMDHp1TfVXEpfTebFqU
0Qa+hyhHwBGRVyqmx/iVlJ81A6SEjNfidk73UA2JBVBUZ6Bm0PzqOO4Nhdb4wlRthz2DOSjM+QeS
6ZKTPrcIMIdqawlBgEUVaXyqtAP65eSLsG3YQFi743FPMndJ9eSXr5vSaGSbg8AdmysxhlV6Q+PA
8+I/C/W6jxgAa/1TmlfTxIR9bZnHR8M492I73+4PBuoDg5IliRuLNUJUfrovHuUJ3HnLmeIf1KPs
GZriabmW0Fmxd1fIG3n5Neq2djlBYTFrHrTvaC/rC/GDLzhcmKMQSXPhRVqQUCNdf5HAeJJeeTp1
m5KeD5d0AgWShkbylGNL9UPLhC4kBk2rUFgt8HBQUty4YV6jw+Kw6DALBDBV7Nd1U0wlGwtdRXyf
t00/9lz5rqS/glWBVHDX8hFkCwkUIyND/k3IKrvPGgrSvqgDjbFvMGby6fKyyPndo21Jo2YEAmH9
V8pRKjHIULtwn5p4hcsQLsarKe4VX31uUTC3Oe9iO2pk+SphT/US6nN1YVpqr2uZ0s4V3gK3NzPD
uxWrPiZUAPTvXS0urG6dqR3Hcv7ldo+5tdKG5IL+0rEU9eSy/q0nFp4f0U+T02HWFAl8+FZEy7he
lTQQLckYsU3I/LplgkDB1E7ZPOxxOvzup2S2D+naSWQWdb4rZdQalV046+5wMmLRTwPkvCXz4m/B
3sGMcq24IMjFN3LDSI2MisD8XAZFKfAxLYYQ1/14J4lFvTEX6LGMP8HmEJ8PzWKdGiS5DT7nLpEW
Ho+y+znTS4Fi+ztDE3oYC907BbSyvbQQWIe59gxiD7ClpBJ/e6Djx4YP41GpicTSfCv8ydRtjPka
als+tx3gqLhfasP97eMlDntBlozSJJOo/4Ox73FmS3Pz2ic+/SFb+wbyYYG9J86mJKTUzCScgMHf
w/4kv5g8bF6xBE/Z7f/bnKfMpL/hcURbBRpP9YBjvaE/pMEzclOThAQ9pJjLpqgCvEvAJhqsK0HK
1+zG+43lEOZh4QIobpBJyuVxTZQa+GAMZIpcvrYENe4dI8AFfU3E5lm1BhcQjIMjQSXS5BMmU0xB
7htn8QG+JquV/IgtcOWJgcGzDJGXxQmEWClqntYNp99rpUSG2GSzzbYlkGmzIVVEuvQzQNJPiQcy
bb/ECJab7z6+IUhzexve1dhbOiodXhvbNFbuqGXs4ZXxZ/cicX6huPXypQAdRKJ+WbbI1REv+GrI
LccqWC4Qeexyz9DSJdHL2qbzcRMgnDCLkwlUQgEkZC5XdpuHeIEySyIquXiJ6VCGnS2E5JRg8Zdp
u9oo4DVIOIuPdfqNR3tEsgHzywXBRch6jPTr4a+AFRm1203jFOpzrkioUcS2rVw9glP6R3U1MJNk
VyJ4XXNmXMMQLrncs85MCReqvP4Tmt2WEpUd2QKvEw+Gtx8DYpghO6yTrncmluS5Mc6iPWDCG5Ui
XQYWIz5KPyyZfJXLsDemBqYx3gHAlc3V6iD2Rca5P8R4ef1MylNhySmTSYVdwFUV1ZO60hmLKkw5
C95cjD9RpLCne55x32fBdchDhjfOKAx6KLzCngvc8DZI/rIaNuH+mlUJIYhHNRzfwZ8CLKG7vWDu
+ZvpooL9cUeObSVI8qxNpYlzmkqcGzpE8+EtF6nUhz4ViwAJBCmSDdwgXH9ljy5TbV26VPBaYSyh
Mq6+fC2cDRJ8HjQBZ4TqKkLkgO9Vi81phbmzSN1XeFdSrVp66z/BQa1ODMV6M/HcWhJ+6cK95zV9
hHfjHlJsLOx89yDI2X9zMCjdBbjICocTdzaW+ul/bCjXYMnYIUO2YSomPvdB8pYzwO/iBWK8cmTv
C4zfkSRdKn8SQ4cQ47ZEFcSzrRfDGVc6k4FCAXm14lmSNVv4c1vfVXK9AdPxG3EgSeCLYWak7Rt8
koa6kqnp1Cm9PJdUTM2YgoBYnTOx/JkHfQHQpDNgFEZlI5ohvAOhgmEL1Yt412kJuyJWSr9VE75N
8i/rR6gemb8mK4FUGhn3j2+xOzYVMXRaPtzi0yDiOQ4Jd0sr2sR0HqIixJrIZ55dld+/+B+z+Ipz
Z+kNhboTRAha8h7pGymX+H0YtV0+PQ26EorpoEyutxnwKUOea67F1t/o52YKw9zp6zch3nZgrGFV
Ry0PXuumcD3OfMboOwLcCbM7wNrQmhrklVEGb04g0Xxqo/wnSLv7ihmfYdbdQbPcxXIWx7q8SoFf
wABaEwxGsKuysFyQPgUV3hxGEPwKaOyJtabGj6ae7z9TV4/p+SgeoJ6GA4IPnfBpP4AfU1zUf7Jv
t17G7hJbKc4o6ohBnPMJz84oIpWXKGWsc336x3CfpTURCKSyelKRrsazbYw4u5xGOsS7RB28/Xc+
NjK/4LArR3M3wWgQqfcHWf4BDkTXYPVBV+FHa1o3CtK13aCi20H56DEpPbC7yIEGGtsX7sGu5RQi
QcdOTmcuXhA138HydIPQQxof5JKVnexyxc6To73QAq5tvoFlVQcvq/JEWsXXCalS5nHbybxjQBY8
l99ZL7x0D7L3UPfDa9kuxzxqcq6y65e5f7Uc5mYq18RCw4R3OnOX81iqFVjEzhsOiqAvrcInwcnX
MROOFEbA4hIivEB0fE3FEPTIqlZRTKSVKkGUGrkL9QIt7z5lb8AwZtAAChxNI3YxGnC35/6SZTik
YM56mf2D2fdMni2ViQkVc9Ukmi76tVGG/dujBLJprqk/BjH24BZr1eOr53IqdL57jbmJEYHJ0gkY
7iPSYF8N5NpvlW/jfpdFkBfkTd50BxTA324Ygy2wY3USTA9nodV5RJnK1d3FZ85AZIXyEH6WWqwF
qOOWegeKgjGoVnPIWkGmRPqyiPc8A4qgpUiJmlh9XUVMjAYtKZNUT7dneKwuSnRwgbAWytKii6mR
JvS2Tt3aOOF+nq2ul86LWwUaVMWy71278vzU/thi03VSIaW/3sIacI071/YDvusHDg7W/RSTCoJE
T0x7ARG/Ob65lFfUoaGTSYpzHy414KgHFsKcYYt0C8Md0q4fJRgPyzv7cT+3LL15DvyxRME+y4SA
G8Gu/rgKPHk6k+xrnuDplbmudybHM8W9rwOhfbrVikGgw9sU9XSTKi2rZpflExXIR476d1gSBH8C
swwhoKh5aSZaN6qsPVMxEhBx930+/aSKTBtemqOONMirJnmvDbs5tXF+UtDscAlmtM9ZGlkqoCUe
grWNRemnYkJuHntQsE6UsMqjNKJEPvxNAp1RKdEoXkVHZCN18SzSoBzshStwt3AVrLc7YtxJ/5wp
Fm42hp3ImoF1OVGxWClzN8JKMuJS/zJ+dnAqF3S/HzP0fF07DDIVbe5ctMJvt4O5fg61eim2RLcU
8zFnC8lC4MYJ7WgGvWXxKhD/dWHg95s6Vuy0EUvcVGGfmknmujK+D3YEYAE3hXC+AEVKMVKNgaX2
k5T4mNgtbWZh1NtkmvkLKYY3yuGmg1QE+YvlqHZRoq88bY/rnn3tsofbw6Comm1A+jjWiP6vNNJZ
pX2ozDXmT+5ZgtjufNe7BbG/obxiyCtBekw7gfoabev9atcJW6APPbbZF1MUsLterpkk2lx+zjcc
THSFHBypVO2oG/9D2BWWHMh548s2GF3kK9yo9mO2tGBtin4gDeabYy4v3LNGuzeap/Hc+w9PtJSa
BgNlMBOlPri7qtbDiZWqfMyFCyaXgZJ5FI8r1wUry8gqCC0ReKvmDp0GRwoSPQLq4c0CnGRfy55Z
OYlsm5MeDeooQQ6qXmHMOfaLqo4jVaA76LsRDOoEyVpivay5gpdGTwEKYxnKRuOXjvsG6cxbChYK
8lJjK4a740FgPUCg+ITd/9VQSqSZhlMhUWBvxExTSbCVYf8NUXlFyDGPN4QOBBguyTm2YIKPl+7d
9yhjieCUqgVwe5G/xNN1NS++hmfCUXSyqslFU7H9cBrTgrxCelYnkNhlHry2aubyg7G1bVKSZ+wI
cr/lXiKRlLmQmvrwKsx0mf+u/qyWfy73jT7P2bkEVFzNsKtHBzG248Rv4gjjLO1QGzdyZ/1vs8Wy
UWLyb95cr6p2pCVtoMA82mMZWw96J5tGRURMd9K50NlXQv+4OL1SXisr2iD8bpeVprDHeP6Nmr2h
BlLJzaaP/b2YdtINrqfA5MuY/rQ/HwrKgezELv9dg0qlv7klJrNgO6/IT6RJ9DsAxS6dNQLnGMvd
coGLY1Zt1t3tUgJlAsJvpykMMhGFID4I2iW/WDjDEFddssZIpOSuhrSTlU94s8iuUFlIlso6lKvv
lCNzbRcYoAogOk6ZVpdfJRYyNVCODAK+cNYqkXO8vGRoef2OnUJ6wfrTXTtOoTj9f8TgbqaBiFlS
PecdzI5BO+7+MTGO0WKrOZ46GkIIAm70USlPEo0seq3F+WGHRKLq8Lv5ItoQN0bxKduXOvFB5/1G
dmTCUuJ6ShTETyQCTlxeAuGs8DCNSb0Tu/EtuYjouTVlOtFASQgYr+uhYOjekKOJemyuA24WHe0c
KjoCLChfOh1OJUPG8v+rVDHLGxR3BjpbIvaY5dkdCZmq1FNKXNssx5EdE6imSz1rxfWjNgUk48ym
B5m3Z3K5vaPBCR+Iwwl4kCGdsFMVM9oH22ba74gqceFcOWM0Pr8AXMcl15lq14U3eY60lwShalQH
2FFBokYUnvyiT6X1CLTaJpyLXnHsfwmvrwN0ppcMhARdAc++ny3Yoo6RkwF4X6XZQ5y3KzX4Ubgp
EhwPYzR6iNiTdlDQ5n5QwhKq27sWCkSrYKT6RHuS+qd2Glfe4gPFYD8LNpOl2HSpNvuPC0Cfq4QJ
UTZfQaCW/87nZ4vZxrUUCfTTMZyHjhhzTDcAekZbUvIynKCeM1QWtuYyybrHTkpqsmeZouizID9F
w5psg+su7DKRMGMi1Tzow1J6pHvUWGvhQ3J8t1WCRXHTTgOljb6ThbJjmfXgz7T5cJ0mFt27ttL/
4bxeya0t8DDzZ3wNOXqieNVZDduDqRFttsOGi6lfpyMRl0ORL+MQgptDWZFSH547faFn2U48FSoo
0CfukdJDLDHq8ItHSlyo3n+mqOz4RH9as0jl19ijhaFt1VcUE3TCBxBNIFWB25Mknw/YWL0G1DxT
VIN1YdDQESbi+zCwXQMXsJXna8ML1rPaQpomNkQbgJxh4+G7MbSaQMh0jw0a8dRvcNWRCGaKsotE
O9Hv9EnE8WL4Y7yJCcZlZXtZe0/szmAJ5MwWYEmEUfLOUgxBck339drUARnPP4T5OZJiaKvtqp7W
vOSt/GGA9nnt/SWHklxKzZfFArDtb8XSXgH6NA9HmlhSUzmOpRAoilFUv9RN0SZE9FNNWunN0cCN
ykxnj4Mb36GcXHyTTB6N3mK9yRTfeo2XU/Yi3hQFqblBAy28ulO5urWfuO36YSJpYwoQef2SY9Fa
NoCnA03pToJgJKluB/2UF+23fdahD5bm4mSJZleKv5s7b0MVqXwGYv50CcwTjwx96vkm0cDgnkKb
FofDWIr4SqJivcSCbSa2GdRDZP4c/C/SphlrkkqCXN/m71XOlOmf2/h5DTq/ny3mO8bzX9m1+xUo
qBMNPci6UjnAAY9wNYMEBOQrHd40B+81vRZ1hQGaqQWVrx+haFMZ1sL1/AmPy6Q4nC4J06JsixQg
tC5nZ4IbL8Rg8XJxyS761IOfujmdMAwgsBpjrCycpg/tbYOEsfEW/Km3Xfdy3gMHYwn4jZ+IwJWA
rWET/mh4R/Oxi9NRjMuVGM+jWucGP9cpQoN+hJsjss4SmsYIvr52K35PWdmSl6u86UbjCMREhX/Q
iC0JYMhLH/jVnIiZ9oxNfZgT37cgkUYOD4Eqzj22EiOVGKi3bZzFPS2lz0uK4PQyDUqnHiwCf6Xy
/23+6lcs8nuaDhveCFu4bOt2vcrvrNDGuLIpb9U1hF+68ACnmoDyJj8DVPjZwtjugEkawU2a54a/
DysYzeDBiowerILHre6sbkltZCJg9x6YxAkIIMaSBVqFevb9boCs5Nvt0R4c13HyFRIiCUSZHcYV
b167yzZa5zMWyoKb6/86cCKBnMdLJPaeVwf13rFkcZsKF8SIXN4TAU2coM9g01GZaBzco9GZQrVX
ul8ZjjozqZ2dLlMp8ukZKGv6NR5Rul8XF0455V+28ebJUK0pmr2pvBrUG99E4ocXvvwYt+KS0KZs
BwEF9MjrAEfg/UiWxTiwrFmDkXOyKNGf8e6Jroj/Mk+zFxKDVbovkzwhR6XWblL5IGsUJqvJPHiN
fNOUFJURVByxoSbYe9HAgGlGbh1CcSk7/0vHKP2Z3r2ow9p10Pa/mm6OZJ1C5ch8Y/FqFmirVw7f
ZKoNOwgi9wxWkeaqB8CvmCS2LZqFIFzyN7GlPKx/r0RFaAMqF1MjUtwDTFpR45dXMRpch4uTXw51
t2dIoEg00B+oRaQEhZctoVYmQSTamRbgsgRzdyJtIyaeQch8ah0gK5V0wtj58+1uouf27ZfI6+BH
fTUXbnX8A4Ft7y21mwas8ODB0PyZvfX7E03zzYEMbMZVMRyFLPj99FGVI8ybTXao0N7fZ1NGQN1p
b1kmZho87c2Y4Q6Q7JYf8EXol3FUWy3IoDfbNttWKBdxCh39LNbAfSrIZK7Iha1DcIUaDbbMyaQ8
CX/B7nkO6+AydUFWgnFg36WDpQttBOLdsJy4oaqy40lXGRRNGtLzlvZQPW6cbOOY1mYw7rh3sngp
ehfrgtSi53mTeQnuk5hdhTGoQP0Y/QduDlNHxAaYITh1+opC0fDooZZOnJtIIaOdrBgOVDQs2CE1
tcsmYobn8Swa5s41s+9qCE3vUpWOy0QFMuzfSmsynuMxbg6wkGur3iAY7GWe+HOFzwBAdo4v1ZIb
tCpd9xca6o+2m0a24xMenDAkVAiwOKoXoKr3f40JaQZNNdreuJds0n7MDxP0cER0jADPL2W0miCJ
miKUik30RoacS3F9pNryZWlSxrnrTzefd0xWyiJn4oZ5BK3q/0s8HHvI9g+A5ewF+IwFrNUQ/KzG
aeM6CxEPU8VqvMsHjMKvhnw0NHaZi5+Ckm/JOhlk28Hvf53FJ0fMjTC1f6pQmfx7q88FzMdvvVz9
MPcVLhTp5OmZ/GeHhjYls+KfAvvvwbV54nnI9GNIjfK9p7P9BKux9SPagx67hRdKOBe/NamveDn6
66ONI9vbQOxqDQ7L6JpADI6ECzMbpM/9JKAmVOVU0l6MDBHoH57ydj1HZY7QHPaoCIkA9nL2JTxn
6cihVoUQedzPu+wnEOYCK+l2WSdcC6Wzb3lV9HqeKFuqtV9uBBwGpCGqX3UkXIkpZrX7qFBWjup2
Ou89hjZTk33+bargU8wOi0GdS+xA21z9u2Lym/hidFe2njZ2m5HGU6KP6uQQ2EYPE+G/ed9ZifQ7
WBYFtAaqF8xCDZiXmYRy9oXSf4+uLxxBX+V7P/gHtUVbFswrWbgdYiP+UDsGLBUbP9U2kE6ATBVD
/QUvkjsK/SJgSKzQ9nxQPTgKb7XGcIg/DmMkVDI1E7G/mWwp6+nch7baBjuLQk6mFs+5e8gTN/Q1
MzRND2Y12YuNXXowM5HgYlki9aelGqE0TLmcif5abrWrFtdS6ELndVwLQtz1KaEmsa7B4ruUzah5
mnDmvWNNtP5F5jiuBgGgo3h32l5rVyccP/b9/YUD0msdhV6U9vUBxnS9bnAqUBgj409dgNX0M+io
gkscQgUWL9S6xyaemD0Pap1W+tVXA23kcUsXrodaNBbIbWQHXIuVNrWme1HsMMoNAkTsCQqJEkW7
19w4W6c+Mjsah49J2kPnL6u1x2GbauLcLDb/1Y7tXf6ElNRY0nN/maHtBZxpIHSBD8uHX7D4j2ve
bc6ymZ0E/SQmvdIwJVCjBUFz7mOFc2NzzdQxWOxkggwK2+hcgc7cGdFmFbPxDqg7rB0LAKLj0zXC
HH1oHfqne2n3PLQFAY3N9IpDrDcj9RYpZPBt6VOhIo8f4M3wX5NKBwu1xotI3tybXdRYEHohmwGU
reDihzmWRPlHF+/kTTQkd9K81GU+zftECqY02+kNiLaARUGOoc+5Om70ZXWwWjNPraWw/ycBCIi1
N9wJXbcEduqUb8VpFiGSJCnIZyEazuwQKk/sYZnLo8IJSmIg4vdpJSmM4oUCvivoPtPO5dzURDlu
trckpGp+UyjdRq1BxZhEnn6r2GQt8YtLOjjUzO60jysnQCjXbNcpjUQcIDvn9/EVF/CP/CstUCo0
hQmAkJOElL46k0fYmAc0Cqex66/UfYTrMAKS0DioUYFdn8VNxsRMy9i57URAHcXHa3r2RchMtJzm
2DlRWYzbzP3bzR/1f3VzVIueGA+c+eLfFlcJScxXYCgOtep2VlxXIAxN64PNj8uFTI5p7NEo+ZZU
/kCxFqSV7w533T50Pr+Q569L5t9TKq5THnMxqiPuFfwMNPUHTKfffFKmB6/ILmB/7agNKgPpHsHh
uiigOZ5SaB43xyXt/0zi0Nptrwqc/RNYumj/LFM4kIdqRHhCSgdoJMR1b6iC4FTF2P/ZhOnf3kWC
CpS/rub04kyQCxwr1lE5m8Gc2y50InsKA9NprjXeh/nwSVCRK0q0LjilaIcj0brcbVLNFV2QAmrY
2AO/jDVVW1CWpguKGnBNbVkHiHj7urMu+dKymtCPJmD3FghL4uxt+yKPUXn671KtOuMo3u0KM8G/
WqR02pSeab2ko6EveNCtwlcVxTNXm/1q92ABzAmub5Rfb3toOXeEyJKpWCuwY/7v5NcF9qxJP+4D
z59RY1Am1k7YSphHJtdRJXI8UKMu1rIFH+a1H3T3yS/dricX3ianB8aKHBV1aKmFUSpD94Q9C1yw
zT91O40CVXpfUEwgQbWuJlLlsDl9HQnI6ZjnxJpV10lyEf+HAH/ho2/Q2z8BVTeI4qo8PZCoh+vL
BAjrK7PJBi1zG5aRMqzqD2gs/dIP2oYTqzH6UOJ+HHOdG9kWiF8oj1xUxyiwKaLmtFl4ZjsQTCyr
vjtFA2vBBw7rrX0vr2DDuNNvhDWwywZWap5Dlta2gSOTQxPyvzks5vE3LXxNT0eZiTqbohJ5C7zk
ZrxQbTVGtm1cFBWM1lKe81r+uyXvxSGQHMEeCwVqP1h9Gjr2WwiAIypHA0/IOLH/Tdapu5otHeFA
Wk/LKEMZnE32dEthwQcx7Q8Lw+EY8G40nf2WSByD/puagfj0KOnrfMXb4KetfHbwJO0o1bEu1C95
dF7AwapBKeljBOYb9mUrfUmdjGagbA+lqW0p+pv1ryGszXYHZgVsPGJq6P448XBU4I84RSD+NOoT
0yj1bgtBVKqyA8K2meCDgicYQQ1BSQVilhgsgu8XRa/K8o6AMenEXNdrdnD7oXJYsUs3aD9fbH/A
P2R7aA8yfhvkJV9c9IgvaVw0Iw9E5eiY8zjyCoodVinI2pjg4v/GOM1qSOryGYpbQ2lz5AmGLu0z
LPEKUo71cwbpMdqlFlLIsn5c70Vu9UK1RFHbP8H+HALhYkvoXTR3hsT6kVBbZWWuhgc8vD4Ue4U+
wl9ByuODl0II8ePaq6mWqiiNQ+sPCB0cpTnb5fY6hKF5uKPR9fSrUAxR0EpQIhanHNCMADLm+hkW
yiv+q2mE/gS1cNiyc9Gra6HDLecQIM1s1Fr0afVP4//iP1M3Sj8VJ8TpcNOWk2LpqMcMtS5EhyBE
dELN2iDU4t9L7TncCSuF3jQuSgO5+frJ7XkD/rc859DJmjx24rrSEAgFkrELxMkCXphyTdsRX5+R
iAO5+AqXSeT3PPL2mGmYvfDXcMmJFsz45YgAuoyRMFUvF7LjZdGTsT7p7sLLJxqUtk0obSiRvmlg
x94NqGIZL0EkF83fG6fpiXbIRjgq3THMUvRmgk5Uh5m0uc6vIDBhkMhcHdUnVbiJ+0Sn10e6+WrR
S0D3i0uZUScUGnljk6iOrNRmUvJ0165YHQ1O7e6tZDCSXvNZig109+aciINnwx8WFYZBUsTp7utH
3Z20ZVI9nhkM80DXomDw521LQ/1nHaKJKJtMgRS+XqKXGB/Qyc4BXNeTnYId0l70c6BHFG0smyW7
wt0YDXgPKiogVSd7krrwzF1ccg8griA+CNJ/U2brghCVWQ+/dSAtGwn7m6O263/xpbgUprHST8Qz
+Ra5jp5Ezgz+YAd71dXBznHxfTJH0oFdNr1TclHyXksXunSbeJT/Q83V0frSjdPpV3GRBqmpPN6B
alYbYz3L6tT/yCLA+mdHLnckHr/dSjd5ZOu0r9BPUn8i+EmZHTs5Aw9Kk2L+A/I7IuZCcbZVvoVd
Gpq1POyniHt4CZQvyUFOyJOJ+dBrPrk2aSrjqRMVBBmA2TRibltsv+c9VS3iLG9V9ZwFwDaCTOUm
67/NvBwKV+A8VKyn7VejQApePzxvQBZ8Jc3MC1gr/TSyDIsqXURJCon4xarTAg5dp5xNX9AlNy8F
ePwyzVVIr43zWn9+Eax/AH0q7wi1mc9RbPybFYN2nrxdT1s+x+8cTS9V3kKslCmYRdj3forNvI9Q
Kzc9Zvu+Qx2GP26XfsDAV3VI0J7lq6ceT87qCzWsZVroBcAzkg4DPpv4+L/d2Qq0+G7fctGtz/rR
yyJX+nhx0GKibbDD0gPSsjzbN7g+grK6abbSq985TdIalsnq24R2zSuJarjdbj+1Bf+GIXAci7my
glRVSjBbJkdfJXfIj0G/4Mz5cUB0lAGzWe/3hiokKkp02g7Rk2gZITDNI4e1JY58uSAes6bb/Ryj
QgvH0OCOI0mloa6H9YZ7nQiwj79SR9KHXc5XM8apBJ1VW/rFd4Ij+hQjCPH75QtN69Dn95iC5DWh
gcFW5kRRmkOoSZZFgj7/Tkn2y/+8NV3DVotwdLeKfVanH4sfvVLQryk51dA5lUkoesWoFkvtqIPV
IawkdxQkxPOoJeB4aBf7WmYVcGXL37RfGhJNMplssqbnV9whEZ8Yk7xKtkDlQmivo72JpcRFECl/
aEuwyJGvaB2a9lrpg9FldKbHx25bhQtMZMTa/rVTUYWZHdZR0ikdBBUWt5wexBaPc/e38GM616uJ
b+VLkCzyQx1qj5dkraMNIQu42F2p9yI3suOIHzQN7ksjalfbGwqCi+nKdXKbbCjGfwQrkcHT7/p3
ie7Xey7/AZKZ6gD95VU7Ef8FJ0Mym5Vw14XcJqvxgBcWRRGs20KImpYzgM5Umz/hXExJmMsmCJ1p
vvfUoXADGic/JRHrlYpCzCo2SwFZ4+J/Fq6GVpXBV1lq1ZzNxe/Y20b26KfEGKFFrUuccU5e/Dmj
+MRBol7D0TWfRfk9KJMl0pAjCJZhjGMvd50AJC50JSiQI9h2uqlU9UzUueSoHt9uPJCHwGJkVrUO
nIBwM37fTflWa8inJH17r5hM9ng0Kl/Yo+PKAWZLw63XaVXYkhz+ucIq7+txFvkr8KQRsaB+AMHR
zhp6/RpEHKzxdYKl4RQGGx/G+OthZUh/PmBBoImG0SjgjYHmGuFNgTE5mULHrVszPHwXS0aoyGrt
KsqMt2iEYT2Ed/jO2uL48E+epEUA8n3lSDV9B3BuHtgnICMmkuwOeyqQmURnR1e2r2l1PPJCrbzj
cb7Jhhdwdk80OBaPcp8ue9RZmSCVdFliRN+cMMdR3IC6bAbKsXx5fXvSUz8433lYFeTdo0YXkwkc
eBn7e8p7+ZYAdsjoLvznTq8QGO7eGff8yb1eFlpTQ1hce8NTXKRhyMDiqgcr0cUPgpA0IqknWpWD
CGgyE3jQeYiM4t8/dKtk6DljJcHHOkKQcbhavy82Du8lkG+0GHFWMtkrsYKmKET/aC3Xg3x7VAZz
qX/Nm8CXKzQx+x6NnxmecZqvbddy8DrRz6bCtU8knvhQxqGySX9c9mwHwLeWgBcpMEsBRzj6Uu7j
3AH1Wk2sr76afNQLFs0tbWoIJmbZaMb8o1wD1DgoQ18hxiPSKdBCIFVnXUnqXoQXsAj+koV3k0sv
bsYIn50H8Did5MbhhBN33Q5en6GdNNhI+GcI/rHw/fdTuWOCgNyOXBR6zQe9s9+0gyOFipL14dec
QEyRCjJW6epi5dROG1Vo0HRBU0HDEU4FU9a9gTw+MyNEt2wZyJ2M8pmimKFAvg/1OkyTRdShbCBZ
DP5GEgUXX1DJChMbD+tl2V4IYUf3Kr+B+tsToE0nQI9yTVKWmRZhTG7UElkoXmoJlDzVVU+pR+jZ
NmBEMB7BMU3g7fXX653K4iBJohCtHjv4wlyioneZymxdl2Yd+YploaOXOvzQeIMSBnBX+V46KPVe
sIIsREWWOzRsI2/lHBH+fWBUYTlg/IlD5Qpcd1PF8qFpTMdHP0YGO636RvbJR2SzHkmXgKAwLXCX
p1X08WMsO520dxz2astIDYupdoaM73qrUvCmgBsXc9/JvkSSKosKV2QpkXipQOr/TOjNmXOAnu9y
GNZ14mjjjAiLwErGDk4AzraWEn+cSAuux33Io1iVsFSqNJ+OsWCpf9I4I9JjhvvTpQlXr4IKcYUi
oXHmXAmXUa62v1aW+vYL2L0xkitVOGXcNBFUTX0NcanFGPWznrX9Zb6w7NzTViBO43OTCvBOb5+w
TdVgv5oYAr+tHUMd7N1HvEXbXUoB3gt0YZgp9OKkIE00uBMCtDanP/WLX68w/72h+1+lNaGEPxOp
LelQRkrPNPMqytWpJb0IzR5ZlD/Dg4FHnGdcpK9dprd1D0X5sR+woNiR9E6bfckWenoPAjLIK3fn
DR7amoWAHXLiwoHz/AvQKrnEHXMDcXePwfxp+DDj0PlmKdrk0/QeHxtUDi280hrRaP6jUAptYWO8
Fg98KBtaW9HF/NAsetphnMVOgF9YIw0Hn8bbXLxEul8MPN4OBd9D4FLQZaUMUJXn+1JUN+E1fXUp
Or9I4i4AeFIcLrPkIxWvAOO6EVgdeSKIW/TytcB0oq1K8KGVLovj1I21jNvrAg4k/SJ7SiDi/Ht6
H9pOoVouxqqfRAz4YflV7sopq7KnWllCNVu6Y2Up66B7+oKyVyi/pZYy6ySnw3EYngYbY5J3Ch7R
83LlnsIA0uWYvj6DGpoDTJ9lTUQclDTYXwc+p1r8+EU4af9CKmwVUl67/5DeVlc4cEWuVZ8vJzY3
Db6T96RmXRNE0clVO4gDIbMaqkJAGE3qsSQ6TLCVrw4paUfSbC06MBMtqGaySf9JRd8k3a0LiW/+
cKLlQD7FYKLQsIgFrPIqqmGJ82qgDk+3TD0Jq+++rckdOQueeMuY6fBc8lC0RSpV8G1HUdVvIiYa
bzWgneqKXzNlypZJozW+OYzNsx71LXhQjSY7VwImuCOh83bhtpLDm+cqKmzFDtzDpHPMvXz/LQDR
02o6mkF/oxTUQDGDApy6mOoYAzgmefONfTaPX1am99bi3eoSQeUSP8mxK+VWEjgaQNYVyDYcy60B
OzAKTDOTsTOUqNNwkHC5nOpA7PgJEsAyV50DAkKgRFRYDMIf3X3Xa7Wr2YUM6tUwYfG/dbY/X14M
RU1qmUPxIMjwUuI23jQJ7/k+zuUi8EgtUjqYw4OiPZNtgsMxHeoD+4+qVwBrYzfDUt4+qV2pZ12X
6sGbn7YlAmY4srElo3mx8cEz0EwsvINiBJBPXl36SXhnoOIIBTQH37veRCTY3ByepPvhtvgKRHf+
i8YMR+r7U60b7sDBFqArx01U9FpSazsMbK3n912PrGrg0RnIjjhcH+J9FPCCbhnCrn4KXOveesHm
GocUSTYMzSq4xp523Q0jnnDMJJpiBu/DaZgiN7oXNTEqyip6AZCg64XmvYo0A0GlqLz2kPpiaDCH
FJT2i1Ziz3WDOEoEGEN/NpGDz3Vfe3J6ijONKXR+lwSCKgXzC2LtD2An1cheJsvyzLdn/Ft46Ttd
qLikPZQgu5PuPfWnHxCpd2zXTGuNBQL00yIemaBE6yUzZdTt0JVRCDHQtluhce+UwWXHSGxpwVbh
qpBwQdydA6k/9EZ2YZicGvzYNPaO+luuQXBHfIQ8nNu7mwejEUPPQVpPaEduF+bKvaONCY9aaZvm
qAOdjqcoegnEy9Ul3mAPO9qXy08nstI/deuTOgeYUpqLMYgSTfQwKG0ISeB+y2mO3AOPL3y4sPtx
k+4qSOi3QSaT7nlQvJc6AhAaTs8keVwPCAXTeUIOsHWtVD4tkb+BKf8m7De59+xkZTiV82ypGkVy
3kWcQySpuaLYm2SPzHLPip1wJVjdTsb/N5wD2drVHK0aWhg1q8obqelDJbQLii8TuSp2IpzT1PEA
t644OX9FhNnR2JHZEQo3EqSztKx3+s6LsFPDtRWNXQF+lbDupuR+MD8SfRP1baCQG5o4KRIQi7lx
Lv2MN7xfuAT/Xq4K7kF8Bw7dPov6iCOj6pHj64VPKw5bW+go/HC51/reOeQH2HGdBg0tT25F+FDv
B9tAui2fyXXnYJCGjBmxv0MZM5Zu5m4oUXL9YoX1KlrtwAQV50lWpSNDmST8fCSj41z07K/Rt1o6
PMy/zDbpgM8cP6q6K+1RAuPbBRkXLzpDXIT8mr/gzta266dun/K5vkfbkEkOKgQqSr6iPkiY5oHG
PaX/W5NvgJx/Jdr5xHT5jLp3gnyWvu8OAoI1phIwi6/QmUX+vk20+BcSuWEr+CyzGScJdOD2HnMU
J7ArVX6M1Dw2cbRd7i7H/SYrjK6xppFSW6kK42oxJeUsFrOV27vg3/BntKSdoDO5F4WnvKolAFNh
IlE80+Eo59EFElV2gEIBwLuMh6dA/6ZcqMzY/sbOsnDGC6hEsxWWj3SxHj2hxBpwUWBaMceyI8KW
ovf2EtM150nlzchGFKwhtHnNgOLg0kGiAShWImKa+hHPPK8eIRqrrLH3XpPhvaxHcMgJUNvOfios
T077MJese2Nwb5IVsp/Y1a9Tnfz0G1yQ+/OIuPwtQcJpjEPo6MEgkFHRlmos3/vMyavZEx1pUAu8
fM/j+I7F/XBa9N/A5ywZ4a3DkQA4TtOKKRDo8dIuyEviIpKAYM++xn42HzMbrSBVj6le/xfdsIbu
AJnkBmExmTxhmbQwsOd6k8rxUWxPoJRFFK6W2geDa28Qa7mjmkndPyljo60mOZrgyXM80AQ5dmR+
GfZw0ajkNsyEqdDBtzIbh3ntBWF7cOJBEXpBkvWnVkhT0rnNazDFAmnLROzTw5qikDTs+7ZF9Isx
8HQ3Qp/E4oXiK3HCCEL0j8o1Jok6gWqTfo6HOS/lxBbdPc5X/GrWu1QUURp2n/UODEXCKv6J5HLy
hEifpUnDRjnMS1aya8zdVxpOPXV1K+G5oeNn+KggfBLUorslaTHCLJkDU68xhDxrZhKFRlsOHYxw
l0BQp/hYfc2JIeD8kZ/fDY3Lm1rQCVb8apPpfRZYuFwTaZyvf8JPWqrH4Vr4vE91vZjKJ3VpBKBo
M3h1hy9Kvulu2lAa1akjeobPzApSD+vpHM9pz+qWHm0hds91yDW2fE8gXdz5LpzKsGyh5JRpziM2
nuyxcyRg22j5NmvI1fAuxA90WxAOoWO3RaAjAXtCJdj/h7p6lBK5oXBhQHZo2Kisqrc26HdbA7wp
ag6HASF5vaqZH/KRoAmmLa2S6pk2x0w8FA4khPkSErrby5ZndwkSb0RUgoAqosDnUwqUwg6ROgtA
Nq2rosG8ja+y9bz4VIwvvRlYllmVD0dtyns7KTc4cV1qOBdQTuSBsEk+UkbGuNg+D6lXbG+Hv1Lo
xw10755X5SL8FdBTgD5TNg84E5v1nK3qD2bxk+1STdcloafDz7o4dgCGJkF8u+jPH5QLBY/KdNSZ
EXn3cq4NMWOjjgF/leb0oViP9bUf/y+wRhhGK+mLq3EUAUOia/7VytIVTHlcTSwSVmmfCvxuNwLH
SxnPnDW2RquzC63jepYoFlXVLOA5rq9EA5pyXbv3z00XPwv5n+k7af0WjpMHVuhqgErAMa4CattX
OF1Y13ss0hI6QBXSqRHBTYqq5eRQ6WjXYL632/LKrGXx/4XlZwaS0Hy9efiuuSG5CmAqjkA6tygt
BOWCna4dT3KwNqo2lZrhYWr+68FjwCfdWV2znFxr2lcZNhwsJdQp56EB3Bhno+6OQYSanlspaa5+
Rn9boMHd5its4shHQAURsjMM97/bO13WtQWACbTik2LVRFYCg1CcKtrSNr7kA58Ag5g25JqFNHii
ZYpHmTYpUFFRWKtuMZkDqaUZTLeBp3u5Gc5h7HnqBlCz98/3/rRsOUlHwyccDtqYFTjrbwUf9LJB
9BUISZAUoB9g5Wk6uAETOy1gcn2f5m++8Of5EzU6G5VEIwU64x1JD/YWmdrXs95N/jIhXtKZ+ilT
1dxLXYKZF7Wj9eWd7QahObV/MGZ+rQs+Y1o1r1RzEJWNbLS0HMYgDE5L45X+rEq2yeOQWusIXSCz
7SGRM6vOpnjr/tsEPfm10BdsP5eeT9zO1gNgNKLN0b/w/GMUibz0wtTsybzXviiqylWsZVez2uO5
Ff+MwCUSwg7PNZwN+CqDG9xHcVA5giUGsx3kZ0H/dYaVx9i/gI6ZoXNoFzkWOmIlnXK7Z4d+Sk3o
Y1Qr4lavnU5GuZyIZMwN2Tp+tyfK7EBe9YdwmlB4eeWODRapuN90PiaU+0k1VW7mrq+zdOxsDFDT
QaNBjjfB/L+PGqTzXuX+Xy5ZJjD0lM6GnceoLDsgp02Pm4s0s2qQhqAdnT6j1TxI/1TP9Nfejmje
+bnw3hs/uN692fIMTd75zZwzRwOSiED7jEQHlSjWWc86GseDJoenBAM6GOxqIOQXo54nFch+rFgK
zDEouPTDq3QYDnZfcdCNdhPTOupFNlra+IRhi5RtbE74O1uscoTXJ7YBv7KBD0NqAzsFPHedmcgO
tqQaK+938cVHja62uTkv12fcWyfZFzfbK58eLLVQJu8yu6VHNOgFpbb3+SyaMRmo3ZzOct7eHAbd
xuUs1wT9Yud76uFrp3kUI9S2VZUo/T04UyJQ+MYg1dR5I9l2Eosi6ej13lltuvhvbVvPNe2d8Lnw
z8YUIR6zNjqqEr55VXw7DTjOuCwyWRH4rjUv2brBf26ItjurnhPKi+G7tBgyJ0o2O+AzFh3GtbgZ
DipLT8bafhnOxMc4fqEYE0qf+ztBmr1f3B58bV6IYDckAvrDQQBGb8tRX+Kjd1sEzH7DSSfS/5mp
Ra07bkNgXXJ2hK6MndJR2q9ML3G+BS7rRdwLEA8N8rpXLhZQwznSYxISC+avCNR5wlGE0x3YB+Ea
dYt+QQ3tsbpW7cJwmILhY5Yxv6njZCAdD+TFwy/W//dbqUbzwwxPK+5iP7e7FfYH+fYuWz0Y/vNl
KTwzTD88QaozyDGNE+Of0X7cwzsdBTuVT7jS0F38OIWS624mDadzw4Q8datgytQIiiFb4LPviHGJ
YhimHdPEC5Aj0pTHUo6neRgPNkpROI3vr1s8sY++QXFSE8Gi/s8VIdGSxPsYVoehvMTl8FpQfCJf
940lRxZrM3W5G2g4EeeszY4TtrMhIXyGfkUQkc2Kr4aVe7smXlukpUtSlZA6ojWf0oxzWjbeIsxk
8+J/He3paMxovU9+HMWXOHnfIf9PypjeXjei554bPunGPcK8uOvhkmfA0K8NqlWQdesCU6/JbXfi
k9nqe2u01SuTdsu9b2lRXlhZdUb0c5XQHDUWqlq4cna4QVjG5TPmR17B5gIbpPjuYVn++mCDImBS
tJrUV8sp6GQ3Tt8vWcBe59GllKfE9ki3aDVw5VAobdPFlibu2BO9NJqwnIVkRcqgxWJSUf4rvIeM
jJnfmHK4meIgpCrb3J1rV+sXaGSzij5UzQGUnWsChxVHPgdutYXypkp9kHHtxs/LSCe8ki4hp3vN
nF/PcQYzVXS9+7fuXkjY/cQjIbaoEiUx2iGRVXXr/XSXxxq6m1PBVy4TTwAESMfMFa+FETgMN/YJ
rK4QzZFmoMnb5+iJLnyXAvW6ap7zaNbPzy7zqkjvCgXkkYBc2+5EXspaw9Ka+hhCQxqPRcnkqilc
myAU+K2G0Cigb6Pv3T9N1epZEN/o9D229R4U9s8L+8ck1x3IxNA790uDpeuO7eeMXosCNjdiavSY
niEHIGJvbkcDu+xRTay6YIBtn5/X26mSPRkweFSjLnbtScFfSQKx/dthE1rks2wkQ9WcGj1D+rjF
AEpxZjlISvlShQXtWVg6wYFN2dWyZwqqddXz9EUln+OZp3KmzVT8o2VGWXgcnz4DWIIK4W+y8LoO
v0WrM2jolZMvt7PN/Yw7nQTDJCOiBnBGHr5Kuv7aTJL1F+pqo+0AZ9yvq6U7QegZtzBrD3X2XwUE
/QSSiGUSJILISERu37x5Sdoi7FjsN3tXNIrcvlzYS6bYRsB0AoLLXhILuu89g1eUt5jO5yXfu5cw
QpAXKEgj9GwLYrHaHNOkL6HTyczP3RF+HIg+mvSDAgZ3CdOPZHRF/MiMcyv6qYY7OAySt6FMNwea
NpLj79aF1r07j/v/TXPUcg80ntm1piX+XbxDTvrBPsTf/Hlff6Pz46Dvdou2NVNjvNqr7GeI8eSI
2S6JKTTGbqVPlGm30oYs0TWKY4IAShjmqJJA0Y6MLpqJ5x4H9a7REVgnmq0/BDSLzsyWbu51CCzF
17jteG48BwSOK9ab/UCvfah/a97eLnCvwh10RwwykKZyZcwI84r+CXZdlpIseeomukFKky6uEn2K
Xa3RlZ0G04RLp1xqCJ1uxHzqgIdjis/P88tw0XU4qHWCTwFuBmVK4/GqcaA7RdcrCHnQWAdoOXmA
Wi5bVaDdIiJEzIzlLKFtu3C2aASVD219RRhIsCdiHDwM7+IHUQkYxcN6UCuUENVATv8XMXl2reDg
kux3qUzjB38Iu1GsOSqKM14edClpkQdGPh1gXZHMo7aK5SkMRpm6myX7BL0o5uAX8Q33VdtYCXl6
hgvRniNuo3eiGSlyySuM1YjqGmhluWIhXDRRPbJ4YbF61ShtJnbjz0xuqaiqUnszagi+9Boe7Lwd
8zZG9/atMAwRZjyTwobkXhvXlqAWhW7d09WocMc/i2WbYCA0aqf95k20BumZMQTjHemxYx88jig+
7/NBqU/hmnL8aD8iJ5cLsriSVhggAfOX4NQx7sZCUy8LBx5jid0/qHG3JNkR2LhBon8FEhyI5F2x
/WhHlSKWN5mzmgAJNnaL+J9pwLE+58r42W/6iIPr9gmfstTZ7G5qD+n7Yci1WLhK5ZRpL8XE/7kW
taVrRL28PA5JTWU9NImc8ZKsE465Uv98GVuDcOP1QaUisqZ9BWDQ9+HJkLBk5ToV2NYstM2g9GlG
C//7I5//aYV90KEEwi3DrtIBaeduGy/vSbjK0g3FPRmg5MUd6Jq2cHkZMDIenmCsAn+Hx4ty/zZb
xnwdsa3KX9T2UZHhIUKvcZmvYXqDY1tm940fQ87cC5Sav5vGG2aj1nViMTSwBk1l8lICT8xPZyxA
Am9VcwwJ2SPgWPuHgicX2mcvqbQMxE9IOyyDJkHvb2g7kWxKzxWmK2hmOOUhaV1WmKBtdjBEJGbp
bs/AjTXJn3TCxO4Fi0DQzbQJ691qKZM28pvOA/6S9ATZ3hWs9+EQMKy46Y2LvkUIczcL/c8fLeoq
VVkhCqIfaD6RKACN8d6PabVEKn6Cz/QPiZrqNrhzYBWJG5RO4SBjbrSEmsXTMK9+vpvFKwIi7pJq
+Y4yHFZvzctWlkP5S4Q6a3btDbQkkzlBWbUDsBnDIcoG16+JkFfVjkpf5Y/gQ5LG5TL/05C3poii
gtnWCM1NHFzikn3pK2anupBoxEUIiyEr5i0JJLUajPkgGuEjXENXXI2o/2pTT5N5pfM4ySC5CO3Z
MK5mgjYS2/TxKbl2iA2QXB86hkTIResz37LLZPvKISPrrevLu0XWme3IehEUXc9yUg6PJ57pkepK
YDtCcp3IQRNc+CkC7aI0PkkDvazMCmCFv1HeqTUJfVEBK8kcKUBrrkVQT0R1//Zh9OxRPItywLA0
tNhn99Ej6GvCVuSODaQ6+gwBvirYTA0gLsIxOoaCzSH/fZ37ORxhSaZnLZdHVrWUsPXHx2i9uM+D
VX5hm0AhUnJoIeXwsW+BNY/TGMNpLW14OFRU5iQ5Xf6cCinsZMS6ydtM+kidAl9mKG22oe2qI2k9
vG2tTKR6m7vq+hw9K711TfKS0nATjokHMNQsaCw3NQCh2KMvpcZ19znQ+Ljb7Kv693CayBiiaRlF
kqyEnV4aUtvVLQzxKFFEj/4T5IZgs52QC9xezqaddsi+oedBoHMi8S7BUA38D2O8/pcfL/j1CEsY
8UlK3LsE6NxlYE6/KfziQXeMWJ5ou+mWgrGpRxIKuk15zfMb9p7uKwAegMszOxouN+UFXQ+cRgBE
71u46BtAtEKriwY8yn6NzUplG3QVfWvAOqpnDxLcgbuZ1CvmT1czaxSic4r6LfqH0GKv1WYQJfYe
+zfraFHBjgRNMqq9N3PDm463XrRm3hs+uXPeJRG1JmdgIdupSJHdkFJL1oTyYpvNDaWvkBElOF3k
XXF3hHgjx80Ab44eopaiaRAixrQgheWbOQ6K8RFCEhCBw5yDcVTfNwdtntCSEmpSFwoW9NTG74WJ
K4qP565rfo2yBZu1J4R+7m7nAJyQxM41vpEoibuAHKCD3WiGWfPEAHvLZCUJ+CIlZEHpGgCuAdjC
pCqrZ5icsyIkCGIxbaKMyFdJka/KHRCP6v5xJx6ZAFSKin6VajhYhtLbzS+Ba8SfzG/EKIVXO9cM
6l3iKbNMTE544gImp04NHxyCjkY9/iB33somOhciBofUKXeMQCFPDqTAJqUjqvAcL0l+oIRr6VAG
WggdOOEGrfTq+bhZLqhTtoI+A8BOc0B2AmDDe++Znrhdb85NoF70u2sB8OfJzDBx5c1Y68xD8bBa
ukFle5Od2vFEbsXm6jU5Q9APTVrtd6c8pVEZeUiB3eB/QbK3+MsJ7SLRxE1oL/zF1FuyAnUZj4o6
8WX7jTt+tq+b2P+24Tibp4b1oWlracSId6/V10ZtvTQaq1F44X/Uo8+g8vtCDzJz0ZDcLxgRix9X
PX35khwoV3fIWBHBq6IhReYK6BIwwJd+HzoEtEObS52+HQDnT1dlhXwokTXn0kjTJmUjI0WPuE8R
a+kFQz0CwJDjXSDD1dNMdvksjXLWQotqOmZ3nGpjWGcPqCjKDIFUTwjLTpws5wmxYMlLyB5RDA2F
lQHBFWgXSi11WglXtm10aJ3ULL0Ld9nAEvLl2LRt96NoVBd2uNfSmDWu7DjKpUP2NBBi9nKX+3Yw
uAB4Mk0Et0H8JfcSevJTGioppDaHhuALlABZHhZKRAIgutLM5gIuAjTqU3wwsR8TbWryiImrRxoe
xTByqVRGkF4GJQRZNkVIcTp1409tI4gQmWG0ls+I7PWRR8ILyb+ffKldZHyT2dVbAO4F9ZorS2dc
RdiiClhvuIebFUmkV7vKcKPS6lVgPbSB2lSgRzL6ztV+KKY/aiKPx4VFEQ1jFBGmC6TsYihd8eHh
Ki3dFaFUPsnG2Rc6Ug/JpW2L+7Frumh4z2E3kPb+wt9mjquDW0OcGNQROhaR7/iUBv5Z0BhhkGM7
Ap2iZUltvq5v2krAIxtEPeMmCS52d9+ZmEYum24isjbdkXMs6pz2oNhWM6LQ+sIi/Tl944UlAoeh
dHRv5EhsquZFDjaaVkZsHBoTzVO3LQGFVW3RqzBAscCer2gMW+mS6Rg0w3zJzx9e5qKuLa1Pi6J2
EHvhxpAOov8Saf3GAIdz1opbNHGoRZWGe3DUTzooo7dBIe/sJZg4PrIN8ZHxQ/4yuuS/RvdMbc2F
vFQ1CxSULFNxocQNTY6QjFGuCfZv1DE1sEc8em8aQcu9JGA7Yhd6/lO14BzM3njfjSMBPBa/kK+W
voJ7Wgs5850juAZOG+a4/24uOWUpNJExxCPD/Ai0tr5QxT/J4yz7Phz5W83Pnk1TrLyUFuj/kIdK
dKAZm58LslE/hAwXxTxlNMrcUwdZQHx5h52+hC/3tFHtR7WDoVo/ycY1IjBqUYndHfk68D7coktn
R14W9xhWYWdJLRsLJzrKxCtt7mZ4pZH4UC6iP8MuA+nv4FPHlScVKkOfj+iZt7ZacUJBnhjEwJ5/
y78IL1vfxw75lLDUN0fRSdUx8cAV9FzA6MdFWmDaJjLw6CU4yxYPBfJkDGLw2iu8Q64PFaUExqjv
ubU/ZM3PKE0nHRjJfNSRCWQmtvH/q6KjO1MjrF8R60nX31qgiAcgCBAZdKJaTBnmEcyNkXKt2h+/
gpSAnta7xNKnrraO1lcv0ASOn26UdJa64CiPS7zgsK498Sm9d8CJyiyxZwCHD1txn3zHy4JcPSmw
DI8RptzYoAgEmcnLsHhfnSC3sukVdJ0MHX0Q4dP3s294cOhbipMjyEHocfu2utl4nkSnewMTW5Be
+OqZ2MaJcpy93kQQ7U72uRQtGRuaQ+sTiHI468eNydPheo5L4IntaloDNAHdFMfDMRzoFG1pKq/J
QOwzGPLYu3mmHN0PFGZSHiKje6YR1Pv6P7PGmLa1MmDvKPUlvxVEQzMPLvM1aTMeZrffnx5HiwH+
xw5/OkIcH6raq4bnJX0sDbf+B9Ig+AKlt7o8nxLJPhkGwfyu/zwsg9I/7FGGdl4rJvSHVwATYcXu
EO6KXcj+prZEP8e4IDQ19pY/xO8vUkviJtxumBq5hK2WlORee0nrXDmje6yZ3k2VMioB7g+URbPh
dJsFmKuDfAyOGHTv32wXFSWFfJr4d8YBVK+iW7HHAYsOUM7MKyk3KYBIE4y8d65HRnM+53tRr3aO
kHPs+GgoTvo/xQt0L32kxN/u5mQGgD4TQpBQMzA7713nj8dX09Jzqo5f1HHmaC7OkLPyD2pKCygi
wozfXi3IFLRO3ppM5IOEDPTnfSV3nJUQ81huBLNsUWbhodQ6mECehKARsf4Bf4ObK2asBSs9yLOX
1VXBcAPufbVQzSDIucfGrnDaQhAuF8IcI8VwtU6rk5LXHLKd2IoTIHAEozEOzPahZD1REbos6R6k
F6IUVbMjFlprmGcSCzExoZvzjGlz+sdS3Nul/hNThDFj41/MdLXE5nZ38rIU81R4RxYF3T4Wa4KS
Pefn1HAhwLQYS6HHLzeSAJUtg5B+MSJwTFefv/xHdt5+JYZcw/KvsFJjEApr+rRfzfkNq1bo2NJU
rlrKuvvBEw7KKCuT/CC3+hi7spyy+iQ9RKob7zwSsynTqc15BBZ4jPIDaYmQbeTaddqbui7PfttL
U7nWIBYIMJIM+cr+HvZdR3SG3BigAv6K2oVmRe83beqeyVGURFlscGsu9xpv7YjyAYVFlE6BRaJj
FdjOhJHtja0K9iTNzdkOTRjCWuSMHjswzS1xTzU9kpsnIsbf5Go20I0YQ7GKyEeFweBq4wXwY5TC
SSSXM51Vw2llgqPmAOROfNOYKFM7cF3dyyt+AZa5bP0Ysb3kequyoXvZhFP5LrOZ97u0QmD04PXV
ID0vNUTxwjKBPTkNaYtnFGqlCcg94LYkw5UIcV0BcEiB+76yHw1+qzSGJgDcfYcN+plOrAHt1j6T
XrDrlQa/aDXJduOCE6e49eNPTNi37knQvTN9GRuHvhpTYuD9aFbon8DJ1u6BEG1AqUsQ1rERwhcD
IohrE0jnFKvMrQhw+Jt2AYiVCEDw00QoR+34w7FCQCqVsKpj//wASFhwobtpP+KLw965vUqZ8iTB
8vKbx/Zs3TCK1t2JhMV+hybSEyiqaVRDs3TO8oqeIhIggHEk6wSdz/mOnvVkrYTTdDH+FHPqNWUo
SXG1e+lWTyihPY1W4mH8teR0gflpo5ujt/vJbA5zDaFB0dpr/V0mFh+vGqJWZcZUvOvuMLHKHNp4
QZlqA5LhdkOVJEraptBur5kAZRFWG7pLaRJ2p0seKjRwvYjIfI19ZjpodL7DV7n7q/UAg2ZUqRHd
deSaBpsyubGydaaHm3OtE9PfgsDHL5Am5DLdWCu//5US6bu+uXtnwamWMZjltl7T06FiJLNmmK+4
GSJZqO0f3s8byGhGqyc1X/Rpu7qx1oNNQLFLNtdZF9elYmCE/rTxU+cg6Z7CVXMbtmcyf/gGIyur
Zu86I0sE6tMb91Q4jrN21FiZXHf+kzPbC2UEaAZlPYi/LqKO8++DJ3I1VqaG0KMggD/wJxIl4/Jo
xV01rTyt1IMzz5lkCWAlF3aPFh71niNHpXVYTJcmoxAvU8AD3V1SjploEI3M//koi2vKm+w94kPX
Wv9KlXpyTVAbxdRIjdks7nv6O0NoV1BpyOqaaDCdNaLgZNA0SP869bX+/pB/ZNhex1WjuCxahkqr
QT6yPL3zo3tBwef8cUR/Ktx4tSg8/PH8x/OklBtNUw3LSycg+tKfd0kW8zsx7okxhHTjK1iOC1OC
vVjWMKy1q8d7mcxL3tcY1NV9qOwUiUzceLin9VKTknivkl2WPbWQjd//8C3WNZt2JVcyhHnvqTqY
KPbowavek/xwvnZudmVkF6bT0f7qr2NtbPQrDb0mxZMQM2N87s4YmdGqkVqE88vMQLUCN3i2dZIS
z2fgJe2SzCaOLHMyKDldNDGxHa7463GIr1VFtBLh6+Lm0ChfvQySQndbybAgTlZkkJk/+k+hsoMO
ZUDVJT3b4s8TxLji1rx7T9k70liUgm5xy/6AeEnbOoI3yOF6GMnyDmVl7790B1Hy4zB9AbG3hIwD
klRpnxnf43SCI8mmgY/nSdUGzzPPfV/lXGORyW3DuYPpC7bHYwIfRWW8IGSnGcqu38tySO2hB40g
nU5+vfL7z2Rsa5p9VxXLSz0JOJDyOZnrQ0oZ3j9upJ0lI4uX6CIIpDIt29hY5dHl+ER53f+vylDX
KxQ6SqDW2PRbx/dgotSnAXsdJk4xazRVihp6YgpKYXOQp5pdD+dBbJrdc6y/34fKI2RP+lEB1Lhr
dQP4vcioRUc5tnyEY6H4KP5x/zMnSFTgFlA7MtQxx66qrrH3XcRcCYoQHOH9pCjpSvkoV71F3oRe
E/82NezPUVbtdbKuDfRC6EY0DBrvwzFAn4gabDdbe7Cuq2Nmg1sw1Cn6BlXm5kDOvJrGZd0BgOxN
6ySDc3EdBU43QWSDRbI1rycU7b1WkVF/yGQuZh850ELAuuZB5YDhYZeceybJVpaxLy663FvfYrXy
2k4Z0gRq1whcYC9LGqrsugyzsSe+d4CFrOK7F/O8VtZ/ZTdNdbHh5N54gHwscAJfh3Pl3gltbZMj
11bkxNRNf14cQ5YIZEryQY2jVn8he9yym31ydcA8RH7vXR8imanygFDYZCkTcZqPqzhxP5hLqlDT
6epp3sOfNOyOGd2FAzKgG8Bw+qdoDtZqmwclnag4OewYq4OBmkGGQQOg2iaQGMc2ktO7Ntkxf8TA
AuXbsTc2D0L+ll2pKyaMy+BBjGSRzoPbIlJS3P0ak9r2dTIw0PxXgKCNI8KX2yeuuqWxpQOqrXZU
eTbsVdxNtCUl7hsDJjtVG3ZsqiQrm1xWxB9z4zY6eiLEJMSyO8/9Vez/lQWTec9D/+Vgiupd6JLj
AL4RSUzzlp8nksP25tFghFlTAOryhz3EfVu9TcwizrrtaqB1pNpMQAWRN0AymwRT5Ck5rN0Zvf6l
H7UYRr3V23ROnkiUqke1zYISqTofj8bRvZKhBrHB/6ElSq95rYGDjim4PfFWVBobFv9jGdyQQJ4u
RJfz3iNwNHtOJRaoNhrIJn9Wi7hirZ9LC7ST/qBQmWPcJgUsUGFAXq3vgZDsl+wk/S45hRpJ70sV
u71CilrfsnCnfwi04pMea+uZ+Qzc9WjEMqjS1/slBQWLcH4GtHrcJ8g53vunZ47P8rgYB1QumxXg
agMnoqBQNsBu4jh1LMcu5hC9dky6QEU4lrRCtESUHzHjlzrOppj5AofeNRuDTskJg5DxFTvcqy6c
nKGfkCgY8n0bFARhjg/ScYm8VYrA0Mw9YUaGaXLsR8otjw41gzfbmQvDdXcSGh+swz8WSqQGgVOn
KZioYvVlx6XxnRzpBl8TAuLJuKwDHSnJ4cPByJ86RGxO/1hk7MRG26p9cpp1m3jGfDqAYgpyPlxh
WkwNatHuw53TlPu6LYMEmREOdyqSSBq8kQPvakNiPGTjSgCzOr8E9gHpf6D3UR8uvnnuYSH52d8R
tVr55UP758FL8RcFMMfZku1WYHMpT9hmbIwoWnGBQa3Yg9PZrFrWrscZmBJ4TS+EyRIvHKCMzajx
VwLmvCXHK4C8kYT/COhScjsh1wYpPKvPtwDWUVXXDyiZLDCE/6BRQYMZZ5xRibEN9dGDuZWnt+Kl
3xI/1CwUHObC8R063zWxUAUEFb8fc4+ZuuDLO2todulCh/UkwsFLlXYEFgOXB2pWw492rOHNSONh
dAyyDPfcdP4o0MYRCjqqTn1JekhW3CpAwDXnIIhOOOhrqZ918lu1/rEwpYd5pHkCsdwCjIcXVMa5
6ocVo8i6U3w/ZGfvBVqIce1BxHbpzr5ftRvJzC4OMuavny9x0QmuUuUc/FEk8/2chPczpcJogmSk
3TpwznixiHbKjqR+zbjjtGuu4jeJYsosrIMSHhNvQ2ZmsMbVS3eeiEz1vBYrijifni7/DpHPSjPO
PAU16fdneTbA1OyFhItFwF0Z99eAvbUCzLJRxvHGpZCfslTmSOB7E4adHmAW5AEJpBiTe7cxiW6N
AM6chsbe3muQqmGTJgDnUBrYBHgEf+ftVzdKsXAdDfhOvIy5FONMqApYeI6eR5x44OoBKCkXvb3z
CFzt91syfCIdo3KLhvTSMyskXMXGS4kLJrBcNpSM6c12ZyxG8zQr4xt7H09BqdPRxnPZ+hnr38LC
X5nSRTw/XWPXW1CeAHMkeftL+u/f4ShK4+Stb78T/eVcha3BkH/kXQOy67APPkGgau8UuE9qwVRO
fx5+tO1t9aJdGcYfifnNH5mTP1ProusJwrRDYiPtrIWSTCe3dOur6gswemcs9A4Vseqh0vUe7BwC
/moHtpC9UM143MqiHz4jgIrp7GqmnUV76V5pPSrplaG69dk71ABBPU8skuoLdMxc/59LZb5yojQg
TEKJ7MINwG9o147qP7Z1HE/pFBgDcLPGjqOboU7KFKvzujkjWwBlMPsqW04i+SOp29t+va+jBSM1
dPybfhm3FTRb2lh16Kjp9YXmQqxBVGWftxZByw/u5JB6LQC+wj3HMbPq5ig7t652IRzWmsK6MnNm
a/LD6CHGeWGD6i8vb/hwpmc1IysT3VQUtFn/M/Vr2SAuYI5h0iz5UCf6glNXXoyBiTctGpvn2tPx
B/bgGKfYLFSVeGLCEx2/1gLbOc1ulJaEYaaa+1cdFpa2EgfrVg5MKiq+/T+uNAD8r00e1C3WLipv
CZ1K/21ueQUAXMcoFlNtK8G3IajEGr/ZaHEc/3QdYk9Dx5A1N/jaoJczc63ZpabVDLQv5kX3Hv3p
Dcxt48mO+SVcGpS/GCSpCUa+ZQWvBCZCR1voSBlgdOZ5W7wj1UB0SIKHafdg+disrZlGSqg/wjNW
xfcX30wQ5ywZSaLGifq03kLKtvS7fJjx38i26LDk1/GutdzW/C3kLPodEkkiubaSkbck2t6b4z+z
vWwmDkvHSqy2J7Hs3oOZ0uEs7kPFzjt6FP5qj9KxmzcYJi7UAwAmMrpoesd5AjUBcrDzgWbPqjnN
AQld5VfRyZUGlNzs0qL6gylG5Y7OOjnJdoH+N8/wxbU3t7RzWFF+bWUvLGMihZLlU5Z4pLdfaD2Q
L/ph7pyhqFBSc0+ny6T6b8ItrhV2lOv3qTLjHG4Lvln53b45iKJYl+FD6I2y0ZzC/rpERNAbxt1U
s+zEtQLQ3lPBBQbkb2sNa5PdgwF7ZxRXYG2cYH/Wb70Q+qvIO45zjbya9uvojAVdv1cGDbHR5nW0
OqjHxFnrKa6nI4JiIt97Bodp4OfjGcOIumfytMDOlAu1MO+VX72VexclCrFmUENyoQkeNeSbGaKc
Xq4WMvhLyz3kfvdb/9hhJRPM8dWULTGQ65FtkkrKJnbPjKkBwbxA7hUfZEH75wFsQdSlyt5PvNiH
O54arzDz5Nr9jHau2ot9A8dK7PYRrVruPeJM61q7/sM1XWBEA3OiE2IuNZRA4Vi75bevWELqshwa
SZu99JIZ3Bfrv1ymRu2SjMIp1Ur1OwSbXpixc8hu6KPJRx0tL74ONPxAswjoFq8zSI7TdA4188b/
IfYu3IVY5xPAWYaiIBwlPxD6mmNLd3D+24BKIlRW9Vo3DoaWO/DgcTYzprMkWuUszyXaeW+htUUI
fCWYUNxoIwKnxKGmUBgX8EfvvEx9QT/ZUpWBzfSy1/c1Wco849H0iOZ7EOzCLyuOk9pScFlo4zku
Sq0teNhkTnxYrw1XXu6FOR/+yxTU+X7pQpav6Yk4B1k6UBp+/gSpgiRPUcDtItUzA8o9ScAwoJeM
KQMR2ZvtnWR8f/NDXVbkvPyIODnrKkFYeakxO3N92Xg9VU2cf6Xnz5D1RVupS2159WPv3qS/3x2t
l0O9uJs/AElKk4aYNUSbCEV1XqF5jy93dqYiaK7mX8KmvTaIUScxcTfYOr/L8VJVDaKlQXAS1X0S
mm13tT6foc0AOf7NL1j7465IxWtvdvGpZbWiOn+uNw2bG0LQfN1r2p+D57J1/2q8ViYf5995SUqH
BinIBgzVBvC0gmjcg5DNOIedJC1PNcc8koQFb5/dsHt/24b+QwNdgSrTvsp/nWnBRDnSEpWAQ7Bo
TwJwxP/YsNEM1FXVxaI8vkhcTwcKZzmkYKXNxMRz4xQBDacfG5Kl/fnyE/f2P0Q4ntZBZ3IfF2rO
xfcIW12/4sNa2rkkexuERVGhA4hW3jdeFczGTNcG4hJdouBjELlHkr/MwKb0Od39kBIiQPbjMA3f
8epzuPZmU/pKfBrzx5Q3Md0RvVKSg/m3IToUttZo5IuKMHZnO/UlWOpE0OdyrlSK546vVJtPWV/j
yXkL8TImFZdUDMwNFr59pBHKSQDqR2FiVcs3EkgZxM2V/EY65oNTKLzZe0geqmj3/Ck25cS4fZZN
tlGLeKUtGnRMduebIJxbQBYo/qmlBxrLQrbDCjdaT9oUCyhejjsFrS4Z8jY+9eTNmDd87Ed1We2c
zFnovXsGZgnadd4SCGdPQ6XqC9Xoa9Y4D1VKs703yXIxakiipd2D86uHpbJZ0tWiYBtClUNrPkJ9
4eXBTfjUan0+FfdE4KXuHjYbK90BcWM6xQq5ypv60rWZYihw54OY75PG7FoCM6jGCYjYneEcma7l
PYOmWGlaAm8vNPXbatwkK0k5b4dksJic5N+AzVOsZTFA0PQAM53+m2kd0bBnRO7dBjjBnuW6FEXx
8EDUBxwQNVWEzPSAdvGSnIZC25SS2t5ctyygRibVM7zFw9JrZuM3Q0eaDEnd5XQJUmTky7J/zafF
IfhbX6hUDPInSs7tSGCGqTfrCMgb+kCJ4CadNHIgNqXiFzAR/aClKQnSEsejb7S6jaGYrEEMD0jj
pdS14y+hB2qr9cNldlZ5F8JaRTJrItiOv1QOGr3IUW+3vOgWqSg2XtN0RIc4H9MKx7Mqo4laLovh
jAYqC15KSjknurAJjNJtWTg83O+2Fbm/M+MCLnxoSAaeJFBkGCquISe08sfo6FR4Nyge9A/+VcOG
A9TkBDwIeKtF7/3+c/l4OsdkLxh7GIez5VHBi88RvKqHeqXVSDbTAscPPx/ozNXNa3vFAjc/dhSy
zY4/Yx4J8U6xd0v3RtdfVtPUHXow5DzjKH1R/JLpBN0bI8SJMIIYtdt3oEl/Ya5Yi9MofbrWS+IL
Y6ECGiB/YOJVsOLluRuDC49cK9weINvGTrxdjrlHVKw5B56CiW0jroNYeXKhIXYjR822KERt7hhy
jOEUjEQCr2r2Ia+WtOw+xgKHgzjC7hPwT3mIKTfgMcNiON0B2R11D6+cNfue+hQ51x3iplDEcJZS
4ptJRXUcxxEg3qZcXXeksZiJjiU/7MvUr1eeSL2J+YKoZZw9YU+KgVRZZMemmq4rbdQz2hCwg9AC
qNU+GC9/+BCKUDFW0XnSDQpGNv0C8TWjs88aVxHk/aud0C9eU8DzCgq0JcoDuArDVSCGvUtqxZIn
15v+VDvD0yAdn0WZmuHQfBhFe/ZHFa5z2kfSpDV4znGIyvN7alLMVnHnezSDxMoxjgQjTF8NWo8U
Zb/vu0nYmboh+J84FcxnxLApk8d4POCLpK22CoKHYP5QNT9hUkB28cS8FwDOw87viQG/4bERS30p
EFMXsWuK71B0vWxz9ro1R5pWRf28WOSw71CR7+NnYZo/ZgaFK3pXwOroZm4/cMsEc/0IsdL9HYPh
qa/CPukrKnE/UF0BeOGjMaMJpxj1F4K4ySOVykGbQxFke4mc4p8EU0r/EuIrPs4iy29nGtOVaiL5
MBSYpGIByKEQo3fWB+snuXpUQtb49gsrEl1u2O8pb+I9EznA4vcpTHtuZ7OCXv3dKMbWL6VC232O
0nOy1+KbqI7fg4zRxOAQs2pd2vQ78YtK7EfxAMMYOm8U4uCi3xnwz4Yr2v53iPnzTUtKthPqb+pO
2iESN44VnQuOpr2f9a/ujr47w/N1ZAmjAEu5eSr60obemxyP0s594EFBexFERMYmyXWB4CrwKP69
yZH3k6RWWYcy6ty22ut+xoKShtJHv7ZsF5JoAAmPCpi0orNrHdetmSqpz4aKGRbduI8lmrccTrzj
TvIYGyF+XWDi7HmCg5n0I7OP17BLP1bygXe6D9QVEwPWx2e1D4bIq+w3fB+ZBoXUTG4gHSy/ThQL
wHDtAlt7urqV7qngumsxCrjV65/5JqJfxqZ/33IaBNc4jmirRwY8dYoD/aMD0RztkynfDP0RQsEX
C8HvMT8qyVeDtGz8Tz3apI3pyqcerRy6Y3/1quUuIHI6GTkv/6QPZCd3VsObFViLXi5+ICzjPl3n
c7316MVQKWF+v5E/Afk21vQptf/u3PeKKYgp4aFfK41v7EEr4NmVkW0H0419E72wOf80HX5x7Je1
AFMpYZffo9rW5p8gB/1LwvcfE30LxAvAZdcODRD5RzX+fL4n6FiNn3qSLMhj5uYnboOgLzWl5cSO
4diaUlZ4aIfcg/jWmLVqItQZVRzUPkP4eXYkVL7y5ZlaLk1bGAyzsIQWLITZKGKamKRDsO/2iPL3
mn1PmJYhA9PjiYPGUsLXvRvcbbin8tjmgnxQ/8m0YL8/P89LyFwmVMJRetFlQLCs0VtVM5Vm5lUO
1o2TlxfjwFZWi5BHvH6PYU0LDb8M4J3L0hHFimHqFY8TDse+BtYH4pO3TLcbR9/UHygqHlNpiC7U
a22gFhy7rQUvdDwtxQPwqyKv/Jz3s9JvoR1GMCqIwfXHxsnJGaoGUzwT16WHhuP5anyQ6kpQ/Ixp
pqL5YrZeV0mvKh9oyGckDEiRZhexiMhjgX022adf3xnvcnoD8xmY7l2OiKh22dsfkYQmSF3qiCfg
KSD5KoFiLxfxu0wmozSS9oI7cmsnjg+RINWnYNL0afVgxtxsBiNOsxJCqjpgiiQDODa7HLnjwqeQ
JlrF6nr+iUocKLhMARkL3tCWfyPUcmDViV/OhYS1b8svDxUWAJQs/6FgUat8njrTyv1u9boXfpG8
GxKANnnkZ5oSgRE2+SzgeSwmn2kM/7sUD1FpZvdejU5GB9nVsATxqs2PL3sa1orGwFTp9jJkR52H
mkIMzcvwR/CpgAQgSJaUJrwmm7ZkorbX7iU5jZwO3lYTCU1A/mD6l9DZDfi4Glo0qzc+Cw9im1Pu
Xk++ENkXgoYFTVfl9DduTYcJhAqiKabuxWgGrI84aihtWpd+lXxqvZMkCba9D8i7YVILaXkUW4V7
ox8w6ZSG/vx9TFOHCxPFhsOc5B0FsmCv80Iit3eJllHHHXJ09UBc/FynahLUSPUfCgf3HmYT0xl0
ZSZqvBfDPUHihZScwznWHsP6GY9w01A6s+ocYr6mjjUZxywgfGU/A8q5TmkmTvumVnlIUQT+ydTX
U4/KNfDeAY/l/ugPICzPuWixoUIsqk0xgwBUKnao2Jm2T7jt4vDr3lsIT/g2vejJW/VDPRF4sKft
vAGvCbsly7HBhZVhNp/rh9YSss93KlHnJhniODCwn1KlnWEjpA8u49VSP1SRV6Q7o9DEcVHBdwWq
WsjnvadiJpno157JnlcvYS0ebUnMN1tO4gYJwQg5wZvCD3Kbm1d5DdKztT8Ge6ZDKzckKTindMIs
vqtClnmqiOI+gX5Wnf7H8Ge7N3m3mY0/+VANK4Cb4qNcBtrzWSh0lLizpHHCT5fCdWHkD+46MwEp
1y5NC44kwtkIdxkozj8oxk8ixfaF05cgQA53ipNqaSyyF+SZeJG8Wy+yp4ox3bCKSKQdbNAyGokR
unNoTF3CGjYeFcQgAuqcqA+3MLBI+cUMZRXDDktivlLMLoQaPUNYFJVLtIIXzNCGvmTcitovYTNZ
UpL0oKGB/3dhmdG9a6G+/kQvHkjmKF7RloSrNVXSFgsKhNNDQOHXOoFR2skYXZ9SRHpnXLFvQJi5
xZ3PT8SJbovTly+hfM91Fd22TUC8eLnzA24LuUKoJA7Lw+OaWbkU1GuY1ErZVV/DDGm2KM9u7e2j
FmrBmtwsCK3kftCkKGsv285nRmVogrf+J9HaOuPk4psU4WwTJsEWwsSUCWPpqaR0DM6JhUE5WueC
lOdv7v6J89dQB/opFpUrehqgqKy1khzNmZSpCnYPgz1gp23SbCEWynjqvO8CgudcFG9eqS8e+ufi
uOTqVAiMxyYSHsLRhban1paGVAUuqHtnra+qQUxV09wX+FLQpa7rXVfqLoI4JnvSaenLn2/HstyU
ybj7CGK+YXQrkmFi5ypUJ+YmERUsRuWK+OgIus42/aX7CL/ctU+WweGyQHcYk6JHA/fUHl4btKNS
V0ilF4HEjzfH+CcMeeuoNwOofZ7a8wGg8NV2ejY1WeOLQ+zWzgEF+b32l4SBRGtKRCHvOSiZXd64
29xOegpvfmRG4s+90wxepca//K3oDxYdFWTBFnXuULrajuEPSOjJLeYrubSEQqUcWTNDqAmFEu9X
awVS1A62QEj86+394/FASPTkMy1nNGq/usi8GzWTSIFKgv1cYqGFdRe9v4hYickJoHBiwx2DSB4E
+TiP5s4s1vUP8Oh8fULOTw2nQvdQGQKc3aCt2D+1vz4XNQ38TmD57PRK01tHgPEbfs2JGFfjFJgO
+TY3TxtkbZtBh87lqIdQ7G3zf/7A/p3DhKYedX0/rYI4HoycC622pW+b6gFdvzG53djaEb7zzohL
SpJgZrSs0fOWIPkkrcb4kAcBR92+1JOsmAW+KHQ0ZmX27brjuN0GW2GPzGDfZO5HpIKn8/q/DOxJ
vW6I0rZ/CtJuSC72x9CCycP/MEV5pD6pviPpLa41t3Vj60+IEI5hk6q11Zy+PpaS3s2pcqGu5uR/
XmvNUtc8isefIMSZogdpdkeTQHBnz05GqZCVFOZD2vAlrLcp/QUgF8TGvag5RJk7U3caUgoCTThz
07Cl8PXpI4XfEeVnufgg4niRYXgCxpaU+mrvxOPSbkKt2k+RBguDlAsFIygoc/vkjhbmrKm8X8cS
QlysJ+UOj92n1G2UuxQIdF2+kmJJ6nQRpBvbtKj1mRwaMwnj18Pd05YsFhhvxijJNUipERfpuZBG
8FcZ/uAQeQl02gWWbOud782e+QYviE39MQtFD0BfJwE/1lA4QHe5LuMbOj3u9aa/sfnREDDv9Efc
5Jx8gR0jFYf7IjEGXI7utEImmiUZcMGLUiqNytz8PGfCUB6diDTbFkU6EuLVThTZhiJu/RiKUuct
zwx0uGax/ToUkwXaEAFZIiQ0JAwxGn7/w3pYKkEBbX+Kw/WKcHBiuHA1/wQeuS3kR3qhp7vTCUos
mSfJfjdAe5dTj2OxlM78tgbgmItpEfLATYnqAI6+NQf3HZNgStt/U92gYNUafqqT5rzDQxkYL9li
dyURXMUyv+kPwXK4MHmKWoHjgGBxchQskJ79ytG2HQ0yz00lJ41X9BbHfTUqfNfPlSu2F+BXyIgL
73EFwRX9hgt/NHCunoGktx5iTHPZULx+/oXRdisi70Iwoe2j7Le4M83Yuo+W6sfgjYZTuE2ncs+m
81qiDSxhI4FAPh5PVWGkXGejx81t8c4x19SOKDiTZ1dnhFprpfH43dpC+yAayYHz6BRgv40maYoq
pwTyLs0h5ACdFUnOwD1JbOCcnO6UpUjrO/Lv+hoKkW0yJIrntdwrZHadPgc2v5hrr9lUjk/YHtrP
zJ6BdUhVwo/+yMuQoTbiGKO02BiN133q0GQs1DJA/n1AuMBD7SdiPpLKuSB9uedJvKWT4+m/Sq7x
TZ08qkZixcL7UvRyaIvALpGCYx8qN3OVllJdVIVhRTT37jEk53J9QrJ50NH9QWGLuSq/4KmGsPkC
jOStQbJGD9YAChABl/VZBN9wpuQezYhEqouMEhp+q9npPYDFbv7UWvE8gp3mBPcnnUeDEogD9X5C
vTk6ZWq0MJJXQzgSGfCSobBVKZwxuT1Dn9ncTg5ihM6WBMDAqu6KIIPq51Iyq+dy6O5YYZZWJTT+
F4N3ozMEFyFW1VO2GBtVUeFhVVSJatHmi1bbmE0qskrp9fGNtk2dBsx3liXkqKBH9AQG3lXA/Ljd
tPrSdz3UsEsRfXuZO6nDw6rZHIsz2vcPGmV2+g/pwQtRCsG1q+m5jefBblXWV3bD7m/flpve9VvR
CLJ1/gpBWWsx81PnWilSf/snM+RmviD9VqV4xAh536WcGy/KOiysrFUaOq2j4keIoqeW9bowJNq4
Mqfyt6Qco9cd74j3yikz+ThKHWOFSG2didAghdeC88uS0phFGTgYaOeF8dQp/kyVKufmD0WNhv+w
e20j0wdUS48TzxHSTcmxKcsCQLYcP+fckErLdUPFpDjEvGce3f7OaO9p1QuiUlg0giRKLFwBGL4u
xyZ6N1glmh/924BI+Ovl3z7Epi9+/jSQsGgDjCpB4sZc7fNTMIp7qmq1Tbp8WIu2riD2ZDGH36gE
YQfruMwMLbQhP7NeIOZQ6Iol4LcN2NspNiLlW/Qfq+39qIi++fxVkLY9TVe5KcsIaSaFrnaew/BN
x3GR34gQEANVtwdKZmu+rokcNWDqpMa8vXrGmml+PQNqtLUyj/AfOHnDjvJ6Ic2kMnsa1u1f+bzy
kTmaA/9V2R+6FQzwh0aYndSdMl3z+WlQxSFTcpuR2oRWXkZOC641gn0XpQ4rIqsY/zrATVHriWwq
vbSSFh9S1mp6D2GIfLTeSWqUNI3TsXK2oKhtL0ZY1kNcE9y35UiYwAwkXo50gyXL1al1nHllxJlh
n8kp/r3ALcWAaa1AakTQnhaC2nPH6rt/u0178AQwSW31CZwW4m3PiLSQGPgj+ybw5KZ5sXF/E7aM
zviuqEuWT88LIHmaCPcq0Cg8ENqraAoMXWOYT51cg/sd1e0ygRXjtR6aEZMkFGlE50dCjRoqD7Cz
98A4nwLqmEj9nmeM2Xu5RC7iCZ8r0BYEM2FhY+Zn6+741IJrOg2vk4Pi01iYNwjVcGh7INQpBaVx
+4sFLNrZ7/xXc1v7GO+ZLn6PwHjoirbzxWtaZvKee/DJWQXCm94q4v5geTHi8jEbyN/+mmCwBAL3
c1t0mlhCtjFuaxsfHAugAH+ix67sWB+1sVSWT7E+I93HptM5i+p8W2et/IjDWoQzxgnSrMmJ0bpY
qKfukbOrUcGGdy+DzuhTC379+Rh8IXVWk1gGGaCCpBdeSl5nF2AwuaqLxaM8p5wlxsf9nf86WKJU
IK7hHPu802ZShxecuXW5p7MH0bGAoTaNKtE9IYIqAItpVAw0I/v8IoPnQIM4TP/DD3xq0QfedlsE
bqekb7GtUxcXfneIL60G7LVAyEcVSygUMv1OTAgSOLSi+tkYienIYJ3hOcIcVnANEnxiRZHCtlbZ
8V0zzUi5aDZd4gfZ0hwVABRqOIWGSv3VsT6PO7VQOwFE8DdrZIRr4mBhKQdRMcShDOZtAUMSxiNi
2eJ2dUVW6HiyQoasIYjUlL3Nb0qOCkBNJIwHiDvyFGJWefLtiBhIk3ULPGlj+6Woyn5s4DNNMRmw
TpjQdsdwmmLeSObpI5QkddcbhA2oPgVEWTLZrnp0Iy3YPyARv62kOQJjTVXvY0UbyRfcimoaNmSA
KtfqoB19V6RFC5rrjoxJqkG+lhxFvEewHLubpJiAFcSAOBQNZufY5SjY7kArNOQExhwjqUQ8s1FX
Tk7SuhWFFT6OZ4oXb2rKdvgOznUoCVJJeydTGsdcySiO1/SrAiZr1WGTAPCULqF3w2qKxNLXSL+6
HbfQg09r+3FawPWwduoGwIh8rxd110ZzAhfR0G1L7nFgjUYqzwf6YGx35gsdZpdRIoA/NFd6kvTI
8umj7W3ZYyF8QC2DCA4DJvlWj2voMxuRxy5gyjQSVayORVh52ggZCbrISIVL0mKkWgfXEDPBsaOu
H8i7oWpRhk81kQ8Zx6t8nLxPv4gmVAQRjiVw8+95PTNqSiYhDYqAo4AYgqauDFWUVLt0n7VMA/oG
wCEnPUVbqVF9u5OTvnefnRvt2wY2B8oRzkaSPydh9Z+ipZCjcZbJNHaTvAnM/PqNozXc70GZkK0q
tVeW9tAMTvSsbArX3lIerVwOLJ4z4RPjsy6KhaGnA66Poi95kSSxAppSAY3Lkqx/eJqd6KvKhQ4d
7NDK4CsZViZeLpo9Uzs4NeJvQ5kmAF2L/4QuRjj8nGivlrdM8XhuiYSeQ9dxh94MS5xavQzPmnkB
EBegt7xFWmdpWgglZJruLn8GuKf6UkjOlJTRSvbQH3r6QH1g45s8rpEWm2HvAQqXwa4YtVBKrrnM
l/n2ATC0D/67i/dC71XB0U8LrGqtkZqw4TbJH+hAK+K0D9yXuW8BesLRg1EhbMThZfeHJ55TqXmv
QkWaCE4IqHi2C1mqeDJoM79yS8CvbtmCpcFtZjLBi/w35DCIgEGklyNGaLb0BAlIg3qjELxUbL1k
gU5DRiu7vdw2W7Y3dA7R8ooowoihQmjyjizvWXa4phHXwyLjuHEJL8OlcLdVSEPvYCSoFg5zuTly
DrLwhaEiI3/T7MyEV+Y/WHHg8HYLlauc3GHNoLoktYaRAzGMNaYY/rvJtPfF7xK6bZ1iGV+++J0N
lCQkXQNF6Neo4PlkY7k10ParxSayAXCLJKaWcoctNuWsNouMCx1HmjYSGtTRC9DEcjezy3S3GL8c
Yz+FH+fskDM6ErLYTL4uQYrksPJ/KYgplA1nMQykxAOm465Ospu0qHBX5vwMcgkjtF8i5dF4mZ/O
nhcPH9TJNo1WlODhot5fQauZDXMMKElJhCDP5YiIasitzxrGvxBlutraOzXCu1y/1RmHHRHSFQXr
aM9ZC5GvlGJxJPkExdyzw7CgKny3jALbDKNrnGRF/ORxXrpvWDaOQJNjddRCHSxzhd2n0NYOULSp
xvYNuNOxhqh1x5r1OhUoGXgxRmwcvsfRKqD/IIodCYnkPqOr3QcXpAyacSAvfweUqu43l3CvIFRq
hHF4TvxUc/ZpdOQHnsUITKW2FDNZYtKqFROPIwDI4OqeA3xNE9UKItVKImPvbZGv/vnc7pceyVnd
SbaJL8M5iUsb+LCd4rf1399bWqnSHmBhTRXBB8yM9FMgbvQDiTK5hNP58YC2PavQTuvjZBJtx50K
PEt2PXbs8Kd0EmRktUkv/xk2uCLLki+RiTiI9qy+FfdW5BXO95CbNv9bftjOl4aZGcdIokzo06lw
4HwdZD8U3NDgSsmiXAIHaLelK7HsLfulzaCduH/5b6bLkwBcArKtImn6EbyXft+3B/8op1TqKj2M
TagPdCVnw6KxD8oC4cesk+Rd3T+3t3ESBSjREndLig76RhdCxEeAR+jalp5tj/I6bEhpNS8tjGRX
pgvEIxTieZSXPiEB6tlXoQGrmRKuTCKv/gFAW62AeThE+DYl86tajP343pRhNhv/uwOYmH3Uckz/
YP6deZa1wb/YGyObqZ/45cy3Yhc8PDvFTQlPeVBeNWWeUhhyyoBO8m7wtKfqxNefYckl4VqUIO87
jqaPZej7L4uKs88XU4S0bUvIiGb25LtLKqPYHCr/vSYZAb/zbEExq2yZKPTFiLtoVj9D/0C//019
/ZBgeb2EtDKAS4MReEGIevV5xEB37uTxD/kqKjfqlMAxUqISYtfw0JTo3tA0WVWINI7rv/9bRFTJ
9Tn56MhY5iFu1TdZdYRR2AGus7yggFNPhhxDPhuUTf3YTG7HVsMKH1qTuxgyQ3HuyYJSgVqb3kPu
3SdI29r94Yj/+2ioWVwR5ilINcL+eFmnyHxnKCNwGgWqeT+qX0fNsd+abt/xgssFqhWu+XhqHcKP
ufL8vfjGq96+6ztN2digQheiRdPOv9cpEJYbEvkXwJSktyLhYQbApGhnDwYQElMbjyxYQnkGgUGL
Y2CJewS7uRoFfl4KZUWds0qJnRDKFepQh4SSAZHVMuC+8T7yoc8m0enOL/4Gx9iONSx/mc7/FreZ
bp7i5eY2oTauW+L0APU/iIZ5sfgaKMTBmGpojnaPjI+YZq0RjSDBP2aqpJHeZmqkguun4CeSpX03
a/ieKYX1mGbTlfD+iVAfXL0HLuCcAK+LquK/yKQyIgv8lGHFZp/2zCJxnQgHcPblIPKBGVWBCKNc
gvAxcydqHBlpFQs1xyAGT9d26vh9vfce9gAVVxHzZp7TiiW+yFBaWKoegFyhcIx8FQ5bqRPdhHAH
ggJIY0KcrocSevynwMkH/JBpprYTY1zhzf47cye8hXzy+sHz6IVBmrhBcYQJETp308yp8eMTVabf
rPpgtHXYg9KBIqq8SxctUr1EBnCcX/UtqpS9HodeQlkrp133EWmMCxtBb/7kn+S89LtpuhUpln1s
jroeJFKpejxAz/ElEzo+SUiJdXXK/V5I5hxLHuL7SXF3gCxdcQAPMJMJ4YGU8sQMp1YP+excx0MS
rYFq3TSEINDck/5jxJxTFREhTEILFSE0U3OZb4dX1C7XVOGa7Eg40QhSP8RqydI4uWIjpyG9c7xH
/VMUj3QBQCKTp1m+0uyfDrEFEp3xOi1Y/Uc4BF+R61ogsJhNBFJ1JmbfzIp0HQLbl6eu56P+4YJM
xwbFSLISi0Dw0uVfzjYDxyMsgMMtfUvn0vh2kUqotTngbJe4rEIQ5+rprNg2tIxDeCw7KbwGZxFR
Nd2xFnYXCpMvxAGI8gR9Pu+TyfpsJZbJ+oDHEg2jHXOr/vgb9TTDHkDuqq7VBukFgGMz7a9bgPdM
iKptOoADYIFIKJYrGZPptuvRgntIP/e1gsmqJy4sIb0b0TbD9chIy1sLAucRTFyll+vOy4pSAy7g
7cnhtwoytR6wfSA08DmxjElXH72+YIRumGK/FcoWPHd+2CNVpoj27E1WfTx+nzKwaPulY2AM6D9+
ta3I0FC6tLrH1SH3obrclmSda8g913GkDADEbDFsyb7O83+25HbCoImxafGQCSshEiiTq8ldwnfQ
NlyejpoymHgaiWwKBQLpS405MNPsFVBradY8FaPIGMNYJ8Zoo8de8jEn9LPnApmj+/DeJWbej8Bl
fHT9ce05BZ7ZYObwPq1g0MqEMJNbdfCIF2r2GxwCHWbG3rFyKx3S3o742sarTChvTVtu+9nZuPrZ
vHNPUC3l+Z/HvVdEJBSgWLrw9VTXp0ELycNaO/g+qicDTcOomj5EN7klLC75PoRMQDtyRzYrvn/D
5qFsvMXFjFJ/tfdLA2ddFTmX6zJfLvW7DDI1f9jXJ1xNOg1/agULrKAM1KgtX4ofsVSKyQpLDly9
0m4k9meVZDkejJFYkBcRfdWx5R7IKyKFLDCGHTUiGAqqMirUkfrj5AQvLn9qYTTnz4Fje49rog5e
E88HNTxpyKQSHm0i7uUPKfaCxQ/52GlXRyydKB1PE2IEcxJtXo3OK/DPPC3+fdHyb/g+QYodn8fg
kjrBoEO1ITFDBSadQh6PJ0M+JlgtSRfoEkuowF6+CTpcpBn7kGpwj5nf7nbmT3d//RUhTfAGua4s
ZVPH6CVqftexpEUdaj+ciEKJFtl9vh1D7BSwg+t34p4Z42HM4uIpLGLtrfspP3nTT+XzbJ292TKX
3jIMhff/TmC6sXzt+S+3bEQo5uMkAkUDfhPLIz4pLGrBI4rjpv+yOFAEj7MQrbKrLqCgVqJw0u33
FjOSw2AE8azxsyKfus13SFFh1LKtyUcmwaUKn2yEVHFi672rQYHfaLvZBnCHxGabG/+Rr73alQIT
Rs7waFSH4G9IU19CEZarlg2Dd9Cv/0eG2tuG/vlTwS2fcfdzElAehGZ0K/lUViRDaGhN24VW0jwp
+aAq/pTQZ2FYx37fRDeUgFsu3lNSQXxCxOxtQgh2vFM5x3nrUBMRy2ITv13xb0kRe5dlcJuEFx14
le8F0lXxyfJeQAtmXte9jkK72+HqhE4wX7QmO5X/CUDqqNIOk5Jo3THwHIQnGRI352CFr5eiQaux
l9/vDC2wksR/FmclOQsF1Q303VutupLiav4EyG3LR6Ib0mRGEZWk7dAfVvHKJCWq848lwqDFgVGj
u+se6HffM2DTqYdbvcCWcQK840yEc4klb0apXfET6JVeYqP/P28LzBgQ+xCWL9Edrc3eFbXyEJwn
alZ8i1j44E3uRzqcUvsvupuAjenHSdmKItyVeHFVXp2IRJecygieClRsjVe6ddzS3YRrSqhjfMwh
8qojbtqv7yFmgZkrtvOl2/MakRihiOSI7m8Gz072m6eOK65q5R2/USMscj3yZtyIMB94RqIuhy0e
mwr+eSzEaWX/CYpXjo6+W4KbFhMyOnuDekpy2V6X2DFyjCFLcc0AS0GlX7jeyHeJCrqH2glWtcXZ
GEcagbgajztSKjKwKUt85Dhv9cOfLuOoQNzu3DJvGOBD4miH0Nxy8Be2x2lph/GZSHC5j9Ebcxc0
rwHX1G21MqgHPa0elp/XjsQ3UNKEx6RZXOpgMyLMCIv1AsajXlhqn4eUbQwC5bgYOG68KmX4r5dT
3mAARtMFX2DwYnQYFejLdc1wWvkHM7Aw8bnCcZl1RerTO3JnXoDoF4GPSgEhVGgy9dleX9AvhQ1Y
PRj40+CFkDkOvSRpNHfwXS1inZB8siXSwx4Vjjybcp3TYsxlM+vlYuJUSFblgL8NFKU9nC6ic7lO
evWSI85yfTGT6FoN0i7ms4a01CN/iOQSnrSRLIWPJQO7NIuk51ph2KZez8RZYp558pTygxYnf//x
s4d+d8f36NIL0JiQXVNSb/NbfHbncaDHrz7JxN+RaOFjkalOMd7UiYcOqMft6RRNUeAay2K4JDU6
x761BFmTtJ87+6WQwfD7Pbpe0SWkyj7kWoWgjEIdSaF16miZXDxveUfAFkiKYD88avoz/LwywFP3
6llPEeWuvTa692pphAq8OszjVPqjlnNuvrYqsWPEULywCrBL4I5+iiDL+keooB6mwi5l/vg5qYI9
uhcsE7606tRT60TLmsVrNKhuk3w7HvzNxdGGjd8mQX8ofQuCpaKR4jDRtnFinwt8etiZ47fk3PKJ
CumbM5wcg8ITh7VbbU7FAUPWyAmQrO+gO2senFBur/8bQhNX27jVTEiq8/EZFKUHLVJ1fB/eUKzy
PFabzcv5G+BdmRFZnUzmwM5Pz0vEUp4+RS6wYSA3/3WJZkIRTSpQpCazFaUHHXhOsFn2qMBcBmDI
KKJKW+D6PyWsiJQCntF1skcEZZjHm29+puFSgAALbtpSkFL5fGD7ce4dpisbweASApCVuEqYKw0N
kDZ2BcK4HAPTORX0cTesOSNxw+X54ZMdZk4JV2tOeXKJcrwOvAuBAcQaLTKMZBGS0Lq5ajONcT3O
xpmA/kKFWyLsOdVYcCyUX8eP3EJSL/1zP6/qSy4WmW+ppoyCE3qxaXvus/JM2KXk6jCLUtnDFt6U
SH4Tybn2uJRszpVlNqvEC23qcdEpusBpSfKWMrxHztsi5doZqYkxIoK+3JnOHJMQcV1kTkRZpi/Q
1OmlL7NQMX6DfXOUJbtqfumHosqvz3FQhMwgLw/QzhrzMm1T6Mhg7gLwaUFghzXnhla8PgKmtomj
70C4YsnQP5+lNL9O9vbx4svMGL0W/4IkPSGH0/HnTHrZ55GN7JOjtViNwxkcMGVkAQ4OEKi8uRtS
hjZmGnD1mGHENhzf0P7+OMZPkXa35Yu0vBKQyriYiY7flELTvqGLCrj3QliWIE/u1XQR4YO9Uaeb
ZsNet2JLMAmFoOMK39mgCciqd9tl/qhkl7GOFeh+guE1fRY/KRPNpCsZFsC3Fo+6zKlttThiey+6
lHOyCbqlrEFsLkiYFY8a3MeAPl/HrIFAqynDE8FgQUmzcnGAd/FjfCUks0zwL66mSiv5ngmtFFda
roxJmyvGgS+xpNQOhOSp4WEk9QkK7DgWQwYVNBI3EZdRzyU4+dgIbsjsxR/w9SCK521YYYVyhxbh
dauH+96kkM1eG3ZjP/aWZIczhUeCtVcSW1SnT4iPnRGHZbxUzgBhot2HHJUDgDQaBZ1Ljyx1RV3H
vzJZxmuqnWn01LeVX1A4kutHZdebsiMICUKZDIOKm++FkRsIQHl8DpTtqikgN4LVeeg4cbF24hIt
8k30kkaMzxozJWC5lAXpaxaIEP8hznaGkT9IcAKCvoHVu8qbD9/TDv8mbdhDoj1CaK8WJ1e9FdE9
kmsSaaNs+qL/IKX/90SyaUxfTXy10juyHCwOdghBlB8PUJ3cDv49EHz0mTolvQ68Otmj5HZCjGfL
Kn1VaG/dfddiSqw73sJbHLEFph8+c9pYNe/HinnsDdqm0ceaKUVdT4yjLUiAq+HvpGOFWMke2boO
VNjMNBkuIC1SouIOBdegUlU3sBPIaEZODTz1QgwdPgGxxKOw2qhf2+OnsNQ210gHnY6fKrf7rsU9
0J5bEMNGpMO3zJlEfI5awSRT455KmJY1J5NtRTGij5bf5JRApspnmhUvLrQ1bkH6XvANoUpvFZC4
xGoEJfLQN1auQgQFanCtTxGeLTO0KjqdKfVtyA/wyjBMGeczY5peDaWbFJcW7A7Xus12rESrH1Pm
q817Q57tTtbrz6C0RzgPgQ7I2/5BZbDXJkAgPmrRDO47fcK/6ydyNlrrZNl8TZalJA4T515QIWU3
vQaa/ytYEPUuSiqXnEc2121la390JMSE2336Hb4sbMy94jevrPiLwIxQaHjagH9eGfenGvjlgEhp
zTYAxZ2pb/dn0v/8/ZrLcfbeVTVvpg83bVXe3oMqFFzeewflvu/wigOwgjEsD7qX9+cAhYDSTOJm
ZNDr6B5M2BUaH3DRv0ynP9dD1VK5M2Gku7b9FOzX0mgkPpKANos3fZvwBiwCttx6s/TFt1FTspkD
YMgmDM6enkTMTCkGY0HKZxoaOf/1oHRVQwcghImz1cFMrgtyken8RglkoY+bYp3snodq8bWYvXDG
3gyACON3pdexkMUG8+/w3bsZsGjCo80tfWaWC98X75yZlfujDY2lfSN4TK50y6dqKwxUdHPLae2Z
XlP3EL3c65KG8exg6PEKHnwBsSAKhsu1PsZkBWZ2yJ7utDOin4pxVsHApznCxln+bMl3HuGpIMzh
SI/nY5z3kZD3sUxMeF/uN254km0nNngPoGbB0PtxRJzm0z0nzV0YIGpcOmWPaUDi0UQ+KG/MiC/K
8t2rYRd+Va3z3vzm1MZifSizo03KsCHV1e3W6K0QQL9pyWR4PTe6OYonq5Dj+YtXUMOzT/eQHPkw
HRL4oOliMAEZ8yiZ4ONRTB8+bQJ+jWxKKHLd1CnUkG9GuXwvpsBYiPiawPtZM52g0zP+I8J7bTUh
jUH+nBqZbuwD5TKjZdu109OMd0jLMay6ogWztknGntJKjtJsGZhvp6Z/Wpg0Vlv13G8wyjfYfiSB
lRFm3GEfaahvBWY6GD7UiJqIIn9PokWnIdbPvzD8BkYeUxSYMwcrw/xdPUmHhKpFTq0W235i5Sbx
FTGAdswD6iKZ5jTUqJ4zBqlG+JBGW48H/GZ7H1I4N+DOttO8nzMMzlY7zdXCgrjIyrDGIn1WAuak
UFCBUs9pd8zwViAl82FzsUtZfTTIAz63RH4rnFVSHAIFdxmD0DxNwEEl0LjWTbJrPSp48qDk+HlH
f+zNvwvhUFRBQHRVDtzOII/2GulzcZb3w+iotDWyEknNOwC29VDBignb0Ivs4YmwXDKu6uAyHuCQ
ZCKNIuInNy2p1ZFgWQPI8HRXI2XM/M+yALxlI/GYlXhzxNBMTJ3KWzZ+OOp4t/Nfz0BTrB0sLOBI
L2+1XG7iuERDAnwLgo46WDX90sPyOzu7WyHVoztzR4iezpfcxFYntqcFN167ZIFpmoni/7CgjDYY
FaGimSb/pPdfplchYe1BoALXyqq3gt5aqUeueGhNxjqH+Txw0RzDXx61MvLTJ0ydrko8oF/Cmqld
6vLDPLTE6x1H3RNHJOv52F0D9rL6Wg2ulRRF/BvHySqOgfKw3uV/rwSSFShcDEwqRfM9WGLmBijB
k8JtSuOsh/YM4s41NAYFhzO5WASDm2/YlDPNR2E5T9ETjVxweEkIAjkVegcU82HtAsEqb6omkWtU
8PBBOfP96y1yfak4v3ADaLnfaPotdrAaRDwCYBbPis46Gj+3q+l7ZwkBqTkGNursRNoZlZ27c5Ir
D3Ur9nqhDUt/K33anSBZIWxjcEAPaXyGp3xcxw41M/6PGhvwpXoMbtX5RuRCin1SBHrV5F3k8ikG
ijnik8700knCnLjTZxYPENOgTntTbM5eQF7XFOi4gO1h7kS86ZTUBu/25tAKEpRi0ZgAsPxz57py
O/IKp/AuVcvqPSCG+7nBPMBJxQAPy3o2AiCjwnD2tm3EIoDCAALZpKgpHHOPdYBBSfvhLegt4rIG
Wl+v1a5C0tb6fMumeXkxG7sbu/NT6d0oLLmuDmLf/abjLajKkASaLfrF0l5064K7UKHQEfK2dTpQ
0sTA5fDQHpukVQjBYi4Bwp8T4V4wy3kUejFod7EkFrgW2jo2xoYwMW5J81r8NFE1wfbHkPU4vOWl
Ot9RAm3MyswH/0Hxipr0omrYEzS1CjcXinq7+SDrsZNVzGIBAItiZiVCQYjXBRodppwzR1dS5iKE
JZ6cot/ufpL7Uqme6b2xtWNrkF2u49S4qQLRiG94tJgvpBBSiDdZ8+aiZOjgFEYyk85nqeMnFQNC
hhSCm1V0QN0HXtdSG5xS0Ys9VzU4azWq/3CU57mm9kdfLhs0MxZPU2AC5EC5sja+efO/wp65GTDj
hKb2iA9op37BLAByRdb0JXyV1+CXXgsdzq4pRIdAO3fPnScpK90K1izvq/B1ugSH9WAuWsO4jKZ2
V8NSwR2QsJ7xSJ4eGhSCkNumiH/YXSXA0OiCeJy/E5ROJ4kH2S5KdStcn85O8zne2cqmUDf+qAKG
s1rO0n1gGsyYD44O4IFolID6HHerOUDP8sg1D4bbjCeCTXobAGmTFwJAsqF5MC2JModisZFtzHhT
k/Xn17wljAz1FKVouf1cVzC4e6tYQZtP1vTQo2O5Hgq2Vvf0m0IOboxXsSDSjnsKXE6sHpdGY7HR
TACE260rYbf16By/96jKulhx+sClZumsXHzGrMlgupacMQNYXXHdIFbN7yOOzvCuOMmvWIteYKv3
NoNvT4hwGVw/ycMN+g2zm9GHgZxJuKEuCRI9gyOYG5KtNTHFeinBqHFOBJnHgP1JRo4dSumR/f10
wRRFodMay55OATsv1qhLTEtcKcCS+MkhsajUDL3cnd2RhISeB++GIh9aqGiJ5cznpkfNX0YkzEKc
S6f2Kr1uhmMPHSSt6Ohad2e98B47o6QjqIulGCW2ZivJsWXZK6Gj7zf+9A4rI86AZCjmb+ex5Nr0
XTMMFEFD1NlCQ5ZicdjqkdCxFYU+pHG2JEkrGzf9tZJRzjGuhePhFYvxDjjzOd2HoENZFscWJ3TQ
X7cjxeOIqnZcCdChCElMWvWg9exz2dVIRzTxgpo24xoRHqkd3Feu81IvN87I7qzW6nzDQ5zc9X1q
ndaPIx0MgoUme7aGZyoCogmGNm1NeFYaJNub4rQa25TACmoK/HPyLQUbg1CpLuxGse4/ro/KOvsl
MaM9nmZ3hXYB87QfeFR7q2oM4Vi/XUwbPvSEDV3/XOmLS4vSGrL5UTKeV7uKnJJTbJyF6ZH+e8qz
bpg0cuySVeqD/Trz768mZAEEJGGZxp/sOA/VW5ulEC1A6WxQrrWuo555OG34SFugKECfQymisq9y
RNqXzEliWVK0dizuXpCAtPeZ+/QoC8dtc/cPvZTfaRbp8J6//mWG4+MlyFYwdZyKkK6eDnbOrQ8J
b90yc9EDqUVA8ceFXPWJiSyX3JJ+cX9DSglpaocom5gPe4VEqwNE2OT9LVWo2SxpqysDj2ytpE81
ut1bz5bM5DiAaG6i4xUPpGheBs+wtqpoTG5rBSptZVOZGeC3p/ts6std5eJNz2T2FK3hcwmPAGsT
hHdaTqIE6Ps6N154178qM/Y/vo7iRgxcK7vcKHf0juQPlIcEwLPVOZI/gEdW7amVAAjUGs3IBww7
WojWR/M2AcpPHiH3oRZDzRiox/s09wWvGFnCXfBt5o6C9v8xFA373bAQPuRJWAVgV8hbn9C4jAal
s+ZpAP4oEN4oCDgojreDPBJcC2qnTo/yAQA/32BB8VSCB78GAGuwM3hc9/rPcV/HI6kTtvtU4Mgz
U32nrnGsd5uAoOmItipJe431edgTjHnSKsrBtDowAA0tZ5NnQKLOYA9SqKMSn7YCFyxzrIizaBpE
afZlYXmwWmMniGsKVGe3QLrsw81URjVGp6YN1pVmdFkywsKEB/Uzl+qo5JFUD7hF4+SXAmMx85SG
xr3FIseodFc99X5Q8IVHmzfjWcZan7JTSPuaY8w+D/rXEzqhrWJbmHbmgVGjKBW8NyWCSssKaU7l
+x0WJK4NRldZ/Pap9gcfBq5orsIltFWaQNYkbcjzA9oXZsVKg141Fy43r5wJV0WfVF2fMbEDbrA8
xTWxkCMscF8Z8NkSvf1iUqWMQO7o0HtuMjCO4LyABzyMhLgOraFkpriN2vloe49iygVAwNxTL+Yt
V+zsqe2pw8yjTubDhvIzk3TbR6BdaX9QaSuOKZMH7/LoK3kNx42RiQx3tfw0CN2zshUeJLXFyWKd
4Rwn+k0D+YLT8GnvEPvamjCI1ef+YGRjJ9mfODf1yqzRSMYScpfprOK5nHzqrnlqzvg3t5LxC54S
DqaPgJ7DoHlGvPvrVv8Ov/ohtboHeCqf/nfIdUHZhd7PfCnuKBTS83aGmvNrhnR4wyFzOegmwLzv
7wwkw6dKNcpZcYoF7+IyDZoSfGcWGsEAJRW33Pyj1VEDTdMjHkCOc9rMr/zbio02UYvUXk357iu0
K8IgXzrnkJ+25lVomnmlcAoh9YdX6BVyHbkGT+Nqqix6w7CxF0Mh4VIpJRGqZNk+BassokHpDP0n
s2KJvO9hmoMFtrJLxv0qWTUvLbTTR7p0/edM6XsBI+EIx/vTMRYLOHR3ZUZhsC3PSxE9OGFuCeeE
cM1PHgqc+ZBTcec45tnPQQAwis63HKyUGcYclx2JWB+p0HwpbKwgCWOCJmakkfjixaWx9OemFait
1gkz9UtEWA/WohnrZRhI5jt0pJd8lx5uMK9d2tLx4Je/UTuyg48fbAW/u35TYKioltht96veYTy8
2Bhe5xjLYtm5tD5L05Kq5ZzSC5yS3ldqxrpgUChZt6Xs89j2bze6hHFSWxjQ2D7L893ELhkpzv+b
T+L27oiHBlqgKrNxkybAv/Zpcrl45e7nRJA5Kv3R7BhVb01KQ8KAAuHS9NWMnpt/Yl40xvnJzKd1
bzKpLVtffWXY7ktVw2/DgwUNroUIDYMGUUF33jp/CJR+uVBxoj3LPlG2cbsJ47rN9XZ5qIfFYlJa
JOcgRBGF2HLZcKVStagyqxNAK9z2iF+rMVU0Fhz+7Tvo2dl/OCJszbw/KgriPSe4l9VUehxddZfV
8xqrLghE2eKKZGvgfyAfGx6HBbayOwZIqJFJPPo3cypMJlxmfu1k9GFcW+d/JZ454BhHQT1UfR6i
uRUxkjxvQ/Ie3uqUcPC0y0HfKkp0dDajC2lJhe/2GUHbAS8iB7m8JOaiUhD+ZAkyVxY8iEAkJ1wH
entTja3HbewzNyI2g7A3nHIHR+1gcEUWCUpiRhihajdlOeFHDhfSYrOHCM/VLtmxPpxsne5YFv9D
pFqoVGFMdFcZggNjSoglDpbHQjFPJRVuXXRfkSSKcLgZu1Mocp/ZabsSYH4NCQjnitqjMbnRmJE+
69BARSWv44Chxwphkec8cbk+ucSmndyABdNibkUgJzAco/v8yTVolL4jts1+bHvVcIEzJrAjkObB
kinmgzOiZjckNGeJ5PD9+W7uOc3dYABJkp1mZVXco+hLNJyP6Hwakz7D38n+uNHkZP+x8jDxZCRZ
R33rEfLZ/tWWDURnZxv9JuPLsUl3YOZqQMa4WPSaTFqRUKNYo2KvGC6g/FEFpJ+bQ70OkF0d3nZx
cFhVRDziYuvMaAe13LN6H+smvfrmyYGfhpvAAJcxy2Lzre87ez/u4FcLQDbNUuWUl48/4cnqercx
8wc+V3Rh/x1DWgRksa9CYnEvLolCHspitpPIquESaCTuWd3Tz3thJTY0qX8krLARV0E12BScXKEa
womJXmEhCJBYGvL8fq1O+4O5eZARbmWi9YFFw46jfUu6EXV3fkP8945z32o7QsQCnTWSNe7/0+35
F9jAXBphAPfKyMiceuW2YoQCkyQ9Ndo/Ajd9b3FoIXqjdAAhMOFOwrTyP1DbgqJR+IkHGZO1CxgM
M2QUk750VqTHQ/3DZWApvKqi6TLfNDrjgqrJtTESwgWmFAyqLu6k95k/S5tGMZ+eZO3dKj93MNkV
rT4rPt3RJBV6TZfpBwy4wJuNxrowYc3lvl2LsVUpfgfaLC+P2haGHp9yVGEVezJmEv/iS+pJcKuc
tq/1Hxsnk8kAY4OZ99YhmmPXmgxjf09yPEsv4pSIIHcgBgOtuILAw7+Pxd9rbwzig8plk4gnqLaJ
eTZjOeixTFGdPRKPb4SwkkBNjeB8ykfxqfF16flUm9no3v28MT8qgIcyuarZ7lHBBMcFn5b0G8gs
ZksAkJWRXsXyLV2lH3/towl7l+p8bIqcdTnCo5+B/5u0fmn7G4Gz14xm+SsBWqnDB7468eJekpu7
7PlZAwG2fin1ULonTl7b8N82z7MGw+UjVyFQE8+eavT0MiD6sEU56otno6LBw0g4OK5XylT080z3
4PinOVAUTES0AKMO4p0QafRLQXUpk4lLQ5N4f6wqH/o9H5HMflQoeXDlj79wtf5e9VJ68Y6cvKx0
3WU+67se1zDmTOjHvzC39Iq2V4FZ4nC8v4/p5uDCGAea/s3uTBz1a4g0TtQYqqhFBO5N8YCTRgNA
aFf/K8+nWluCw1iMy8oz1eNUiN+CwF3ZRo2vxKy3gYORcf9AkkkOutGZ4gWXzcWviINXuVvOahnw
MislnZoD1wr05ouGMwoGXXsGQvB2tEkl8zKR18xys4GdKznL8GCpCFsqGHCTC+ylwMGx0X3wMJAh
JxzqFPs0ZS8JrVFPy2RthCS/RS3t5mKL5eCmHXuHxq2hUIOEeXzpQLw+336UHW6LfKk+/Je2BOq5
B5LGIQuHoN6SvnvVtzcFOApQjFBLptcVjGLWJHBzPXsK2WnJ88DpB2tKKKz7JJnJVPCHSVhn21aV
2+K2DslTGxhiR9na9joaClMarFh07IUkXL2UOg48x8/NpA0YHzg25GbIb//zI12IYgfS+CoBvKNt
5WvQQANidGQYOKo0JB31AMzn8cgAbe2rF8bDpYrNQZL5fCLsb8+nRmBP7encOHlmqRzL8LKlIVWm
zxIJi6EbraiFwTb+vJQE3DeOuHF3M3pr/hCDJAN3zFqMfUzvLlSDYGioPFG5tBHUSMI3rYxFfDPJ
2DI3r31q0K65ba9IzYqGe/yO5OIZlxRgetNSyNl8gW1F0pwYHZbWgrDIhWobxlLVZ2HBplqlCvlY
LGyNWv5U3RSx3AJRGtbtiuKSNeQXmdmEipEo3yaeyT9OTAcGOZoCp48SQMxi7B80Om8toVX9lela
M0Wlw78iwqzFRY9oRYeB/HeZmaQPixBNdsxF7JENgPf9hLxfNyKjGRAzXI9vPjiyx5edFDBTsyK1
Q6C0Bvg2vyMhaLo+A7pYqk/0Wxl61Ag3ZcF9IOfEWuYeRE5kMPVmRStgb2Xy+vTxdt3hdsp3plZ+
gOcOwe4SNp0JIfn2cdG96C47z3ehSKv/kLvQfB4sNmeVoAmCXyPm9daYdMhNtFjtDChhFRw1ZKEt
RUik50nqpAjsu9pGGGy0SVogTvyoXKzYJeGvV+Hf3R/8yQHlJLY9Sw4DYY5Y4N4kE3nczTQFDOh7
wT0R3CfqkQy5Msat4Q7xVuFfuEnvTEzvbWD8YodPYxwMCcceVhfJKbJhKP9gaeHY+Xf5MrybMNZz
pyaZohO9vVQ9VM75ijcPTXmDwP20n+nIKDTDYHwFkcoM6mhWBzb80qRt3+zM/thfM40THYCWlP1j
4hnGTNCyXcu4tOFAD5m2xOwCaKUw1WBhL5K3w3C9xGwSHmoybqky3VxXZcfcZ1qf0OHqMOxLXtIy
B+JN+0PuuprTpDdTUWuZId31CAaVbJgXgFZsCuKRV7u7O2BGL8XToUKgfcK8dmSjaCazAN1AeOKr
sZvnItzU6XwnsP51+OD8eVaHU5NeeRFW3A0nxOw3oyj6WSDzjHi2XVRoYS95ZQoV1NuW29P6H8R3
ElWAuwhM6ASGngcnblrpYkqc3ijTw2BSCDjLxJg5El3ye1mmD6PVMG9mcMapsMVmowfq7U3TjKKA
TykS/jr3ZtfSERyPwj8mBPwY1hh0TbSscQ0KkeMsXat1XYj1LSoEfBnXhMK3uE2p7KjMx5xIY0dN
lbU3/MmzvBTTeQOEs/kxTPZ5OETqPqDWzNyMsp849EEXb6rnC0TVQAbWrDD4bN3BuJp3MG9IhkQv
90GYfXqVkMW1vvgVy0GVW69Ku8MrOK2/1CvRqGGDZnE+sBEBOyMwKMHhJJkxQ5vC7aRoP0kwu9BW
Nik/aMDvDW0mVSkg9JLWvddA9Qikwn2JBO7frrHV9lM8hTgdVKv0l+IQxWgaxaTvM37o7FKGotGf
p/hto7KgDLRUbINsSZNQy5oCqC5WHnsxwlubh49C5tW1ZIQwNYoTRD8f2DqUCdGxHFw+IdwI6D9W
7eAe30YGec0gdONGShpBTco+aXzR94+gon8/6whZYZJo4SFaAADw+OWhKOO3rLkVSNPmJOFimsVV
qxaYk/HtniBh1Zw+lnwUMIUcMWzAOYCPHj8RMEhV1pqnxjS6Q33wJaYpzbDy5u879gxzqbYeLit9
8HuAHjGQ6zHWojG1Mo0R29FiACVX/TL8YNDqW7Qr8cWqQbyw7bdNNvf0oUQq6e6f7rBdxdXwk9Gw
lpiWN0NQFe181CVNA8UqK2ck3ycx+hja8rNbOlXJdJNSzMWCK/EhhuwKF9Vx00Wgtmc4BSB6mqi6
HqdbbZNn/X9SGuRta54vxcZ895xssjDNJAsLdh/vsKUVmbvqzrJg4lvY/qCpjHnmbDPmznNt+CT5
CLuOhHRhyW5bx8ov3oU3dLu4yearYdnJ0qHbL/ZFt27r6D1o4/IHM9eKX7+GMXeF812QS2ZH55Bx
DizgFwe2mPGNg7/Bc7TXwxtV6uP99MH85NA8rG4zwB/e4GvzGEu4VhtGsXQhVDu7LiMyEht7CVjC
N8v0TAVi3VxC49qs7wnM3YiQIt0bV7U1G1D+ps1pjHnOnVpQFHpdRHC6bfMhNdRDJIhbD7BJA3CT
HAQcODjzL4t9nxQtdzCddpNobXMQY1CP4KLlzW/e3vmGiGCkmrmZK/7p8LjWDFOHCuIKLtBCsSxB
fTjJnOi67IuzJV9ybJjFu6erm27qddOTjAo0X3U4yCaTypawUKC19IaTLywNEeEGWUhNt8dDtZaC
Ngs8MAtkw6KSip9NaPcDO0UM2fPWHqC2b3XJ00yBq4UNWdT7THbU/rpin9DjruqS7THoBQeD5jEx
dqZPDiqo1icdg6WIjyjtGO285aNKeb0KPBGtfPtsGj7XG0WOL/gtcuBZPtP5p1HFI47CkKk+K4zA
JoVk6JRlg2/Q0iMwzHurCG6TXwxsYku7qMsNwiZTFf5sobYAAauMQqa6sd5e5JzxjofG45BLEULd
Wo/a4vc9UoBOSu+Ohi0Dye75bIZOB7skL8ChGCL5gKHY+syPu+frsNmGZAM6aqzWtVDuaLTJtVOd
RxFJYJuAsH/Zs1af+eTZ3s9aJWVtEItnlzOEh9KYaFJr/wNMPq1uM+7nq3t8SXiE5w6ABEFaTJHZ
9+Yj5W1NIL9X5xuTK2/sghrM902ZBHHFj2V8qPlfMwyhDZwC9XiXlzPOWDeFWliF3ZRp1gisKd7F
nueNSskUJV31KoCBOp5NvZVPLZ2+zVwAJ0Y+NVN3P4wJd6OWNvKFVlESZykVQEzEgG7YNPzlk5nZ
mIsklFTboaS5kMrmmmbF6zmVh4767OWFxjLvXP44bD+4VDhFfGJ2gEGRMDLteRBjdQBTfBAWiBmk
Jd444x32Xz607iEaBRuLOFq8aK9Tiwf5UrU6/DXM1rke7A/D32Ut5/GDeVxuSAuEYZwVcziCCB3l
jRWvUjLWeX2c57EjoC11sUfLrCV8/0LMEOwzMH7NDI9EozUrdv0QSCbEJd2bFlF6IXS4at3bReiP
jUHsujc8KoEhOHQOAMNaz9/VvijmNN3nx+vvNmjOH2sWZvQ+gMLa1j6rrwhdFV13MgFjyxywRsOu
O7CdNjUalefoLbdsvvS1LkmYqg4j3AmfAeRBIAPAO8c/4uinS5h3ilsfvZBqQalnvTKRnFfjxbVl
haPkagwlp1ywiDyZwQckmITZ36u+O4SGWsYh244PN+hNokcBdt+1SpESjvpTbwbrnTZ1etkLjQG7
vC5qYbcBG5E1HXiqlPaZuvg3ZyHI0FhTq4SPs6wREA2bZf7yNwwMehOCsyYml6z6+XdFzrLl7qVb
wQSY1jaB8ZfGBvyOQKhD4rfJW86SIk7lExCOXr0XbfY92dSDKzkmERv0Jok4NkFDXPKW+2aQ0e05
jOzWVaTGOEmi2xf2jgBfRf6LSnUN4ARzd8bbaCHryF7YSQQRtx8XXU9rj4R6I5a/YG15WA/gW1w7
GCjEzoFQtdkzNKTmkKc4gOgMztG+dmu++aPbufpFVVhLbEHvgVBP3TDH7Xokw4fG6SW5EBymJDNY
8iN+0uKzZALzPaZk20b4s69DtIYTPVXl2iYxqzIlsC4AetMBc4ycW1flBRoqIMjhU1oRQUv82XGK
eFyOK/QIENYmuFakxS+qytAHMm1FIUgjgJRYVWy5a5m3vmX+ZUUmNdmNnvu5W4GJPc8XVF1yzHIM
l9c0yiT8kcMWgvndniGYTXKfI+IwtEJ+XNklG2FOFmDXrGVS3VZYZ3xjLL8QPVntOXGT9M5d3qwb
gzBt2bSF9FNCS9XRP7MfJo3bFOCHBbDvtCH/+pgId3mU4fQi/LZRJS9mHvMdKQb78v1b+MJQkQLU
uY1YUjPJtq4xcumdiZYDCFYb4rBol+kseScSusX7yb48a2DMXWPksyOCSnhsoKYBHWAlREPZUe6H
q/7KZjVNB86BvQSGQBquMXoZLC6Qxsfx5pYS7RpuqHVC2h7GUFWX77ip6ja7PTvujY4pwosHqCAd
X4iB/udkRYlhUFyytGkBejdSp5sx/blrrOyYTo8bgZPpTLkcMwZulPbrd8fTA/imt8kt2ACoe2uD
Zc7GfLs4Ri3q3EpTXBBr3GEOKMTxkp2COdUsOiAB3HDHMNB+PYkCc1Uv0pHO709GCvokfiZM+RXQ
dMxWdDZf/0T7hGvbtZsoll5IOqJBtb8JVRsFydTOiLK4Kb4pcGelpr2kU+AQFGuMJTJY5D3NolsN
fgnz1w8tNL3ENQiU938BF2fCyI+vOJecmT8xpzXA9FZSZQtvnvwYE8uhjMMnEp0UdE+atZeUi1Ce
OGP7t0vjlwRZ1CRgg+/OiS4N8Id05kEWEgQvl6TGJTMh/1MPLoW10Hnjv5YDbhQK4TUc9WJhHjj9
aq9zbqenboRmCS1KA0utzl1pslVqAQEGOzFD+y+dbHQV4K+wsy6B8+jRYpL0+FJlsOhl6cS3pqZf
vQ7+Kduhlvt1VjY6IvzkOgxbLGhG0n5DdLH7zfAF53jNxWM6SebrAcG8yTT8MLvSElOfZVkwcZI/
PW/tl585PbyUkgXCUJGL1ZiNQKx/ZIwQDFbXxFe09EgrDCEPqlzVkR9pyZpiRyUU6O4CCrFKQisj
1TnhoarfzevPe4IJdaM9dSJ0KKpYjhRniakvx0/RuKqu/utnQKjGS/n2CYoE0jqi+CntiZAsgG4l
XDoOaAFZmWRuJuhZPbt28x3lmAmtbfZOq+pQrkShvA/cU7Qutle8XWbC2BG75D5v/L85tMFxCzpE
GXMycMDWMvHOUDIFV2rBPRQsidP0j/FUt8OMLMtlSLq2Q2QdmquVIJkH9Cycrb603q05tA6aqI2d
GjTMlYe005x82Kx+2+915OOyiF9zD6rwN0qch+nvzxGE92NA24Ltk6uPaIcmF+Xu7zWsuGjm/pzv
ny4JUMigslEzN0P+/JaqgGdP3rnTcnRNBxYhfL/ChHsvkSx4zO1tyYTgnQ6nVk/7L+YvW1MFLrbZ
cgWU5vgmWfbuWmVFA1pIXkY2ZW9dXK15vyZyhB195ZCUbC620zkkRJJlRFmDwucE6l/FTol0CzI6
QVCTfV2rng1z1ne2VW/ovpCGpRNdjQvTMz8EUSgjsyj2r7nKufUUO0oU2m079IKZ1JipGe7zuQP1
B1M5AYzBxxM97dSOhEWXFecd7MD26B/ZNdMVQ0ivhIyR6iVPLExgGvjTzGJ6qxn/0Q1Eg5t27zZD
uN8nHUoXHJCMhaxaKwBZUfGjcAUZWLaTAo9jLBbcfNn7Dku/mCNvW1WSINFSrP/DMa+4AzXwBzDU
T2aaXUdJIUU76ugFUoSSPWVg5t9QEw+EpTmvL+G1sIbISbHjfdEPhqu9nBO/5YiA1NYKTxx+HR9/
tvEg1aipkHRdmpEy1Hb3wDrA/zITVlPC2sG4gxxYUmot5muexIMT/xc4ob/Kv+3gxTTel94u6TWS
45I69IVsxsODry48fe4fnp4o87ntOhqxqAmlQ5sqlZwDg7a8XSHqxjksge8jkcQLl5zoyXk1hFvZ
8aijy6AGWSlKqYJPNokL4rKFdXWuDvsgY7u3SFXj859D+KsT0/GTzZdIIugwr8MFNJEK8WLPlJZf
qOCNnrd2VyvyCZLSAUEuJjWcY6N1Edc8xU/77p2KtAuhAIkIKpKcIJm5e8LSdFTaYqs8zH5YDYNA
yOLEvSooJSjCPm079u6e48zt+Y0mzxtNOyKV9JR17O879oobx3mPJbK8c4VaUjAEm8J3bRzdqo+S
Yz7CUXiX5NOuXcePGKRdUh3jxjUzXjewTyqx4E7Ju52s0OOhJWgi0aCIOzHFy8ZQ95rLfkgKJlMg
7R6Wohqejclx6OAjhGlSroS5mqAAqaRE3RlFm6DDtMBPhGhpRbimJbNmaxYvwEIm9rC+hPAp/8bX
7rc9wtRkHjcN586eN6x9A7KJs7VYQXHJyrgvVWwuWe7Ga+LbiRBaUTH+lFtS9J0Z4aW8x2YWw8h7
mZGYhiLb5mfZtjvZP2d9SnFWt7sbTXVh/y3Eu6w8dvbSrs8RqYPONoVBuQ9LZ2eBLHs9bNARFtjU
Gjf3YxjlaXj2ozJfpMgUE1QVGswSQHymMTls+nz4Yfcso43dgMw3o7OgiJnlv0hQxXcovkq0b7Fu
YeImDmHYj2QBFX1oJechN91gZO+uqh5c2cRMK0GJNpQYRDIUmC8M18ZKbfEj7fzhoY5nRucFAP/3
tTB7kSqnbsbnV36zKDF5ViLrULbye7m7ho5i20cxAwNwT6ZUN4nRBaUMqQJxqvHIAIgbZlZwRxmq
eV4J0mOeEF3znaQOIUNiGG6MH8VapS+TRie+UNBToew1gz/ILdVXuB89M+y4yZ5D98dGOCJfzo9j
cL5v+avtVhRTDu9E2bSFCrbSM/hk/WyjEv6f3zOdZpbzQubtAyGvSMLmBXm5qSepGL59dZzxubNf
wO67cs32vEXwOsgF6HzpaLwQH9EbWPef9HE8ZvyeXRpc0sg6TX0J7Y9fNBAQLVOa0qh8YpTvXI6l
2NFbzOwfauMSF6PWC7TCF8eOdy2nJ4R3QMNrr78MuVJuzRZCs3UefeQe28dytkRMIVya0aMbxFfc
aoupwWSn5GvX8mYHX4alWnq0v4zQ1PdywHpKVr0xLmUiq21EMmUXHwkh3oL5W7ahTa6XpOKTnHCP
S3ZHcWv2dUcjWV952uUCnutbmCIwdW7JGof3eEX5kRAndkyixe+j59AVaLL7P8NJppU3bNFpK++k
1jsFOuGpt2WKeCa8hiyZVacP0fLCjRQJ974c+ltj5UGj0DVqoBt4AcXtQO0jl1n/vcIDa6xBgEIo
vsbr18Jwxb3xJ42HGUyu6XEkAGWcL2uMgxEZVKyybLpDFeFTOI1Zkn+Zf0Iz+CHdpVWN9Cj/oTYr
01XRIeSnbgluu8fE273UnEWenO1Jc0QIkiBaFAJDN6cDlI436UHl5D7PvympVwgZLoJ488l5f1Ep
vKDrVfjtfSE8qhXfD5r5NrIR4XV3gBbY91PRlI8KO3VtL95LI8IK29iZEL3tAWFKP4jcrI4xsOyj
HFTtye1h3ArxITntz9lsf5SNSyNxUNY+dvawOf2ql/yy3Wvm4pI71G2rHCHx4zEfBHetXG6+FXBq
R+KXf5DrrKAC7v3CebbJHQBbhlirg+MrGA9XI9tGKC/EpFrssdZt06AJidWpn1FV0O2i/V6iaeKj
91L4i+yprj4iVEWv2sVZU0lRurQHMV9QHDTjwaC3/yyK9BVNAYUfUJOfUZP5G9PdGvnWaepEPwTN
P/3MByAX+z2oXqWRmRu5pxppVepy7yoa2R/0LjNxjQsfC5tg/lioi0nboYzA5c++wdiXJLPg471C
pG3nFiqP7iYosuZpZ0Vg29iMuTZXnw5+h8cIYN/WKD8ay1uAXU++6YaTARxrtuovLXj08OVG3fYz
cSb//tk4DRbIJzraPXXJiajJA4zjCbZUiFZGll1g+GATXpTlY1VE/bEvgLbeGnKB5quaLZwnW1df
Nag2nnGnzWU8vhu4G61RleanBWbZVh8kGbDlJ2CYyZeO11p5mAETqDhcnW66QU2NmkHGUy6F1bCm
7lOMGVl0LSZQ7mj2072FQgCADZEp+G8gSs/i7xcJDNt1Fpbx2NsKQRhhGhmbYHZEyXgO3MdgvzcD
q61lC1yC6F5LYGhq+FyCFrPpu3vaDnqkNQZGXsmICdlj/OV+jK76tGvHCiZdI4KX9TXgRBaGh4YG
6k8p1wjZrQJeBmW8qp+or43xw/A5MKzbgWS39qa/IKMxZHIGzLFq5SGssiSMMBdDVccI1voof8Eb
t/hDzr8/eb8466Hk+RI3iQMweEFZ5UjYe/py+zrGGUB+3JUBKBumBsEVd47lEYbbOTVzs9LsDbV4
ILhW/0yzr/LhKmCH0OP/nIeL/dL2zVIz600QRfxwfigtCP3SEkQ0JQ4R9ufRaJ1kKBb8uHttOMCJ
iTJ5X9WHGHtVkbkbSkmiaGS2AJGzg4AtTZK0dfDSFYKwGpept4wqBznj6cRkwoyQHuQID0897t/0
3qSDjSmA7W2I50gHSBOeHqTEXq7xYymBJFP/WZQbJQoC/G0AvGRBUAsthQMupZiqsyWxCan+J8ly
PFJQWbwbvXEbSdHawkh0jxtbrk8sK0aqotghGk6NQXuF6y7TExzc8TlD/6pCbZ7DHjo2uGdWVrtU
f5KETi3yeoxv6noDPwWft0l3oDHp5qrP8yC8pqU4J8XM19Kz+n3ZKCWCL8WlXBtfH6CX0lhf5++7
vTH1NK9MtWJQpI2H+5CUpVijk+IAhKpOnCxQ2lQisdze3WzqUMUCfqKM+agaUi0LJdZIjJx1qGHQ
XU8U53mkmF3bhjb515c8kK7GdwMzBtgDuCzpDehN53QFS9Eli0wB+caIKYL6fm3PDOzbUznPA8VR
MscVJPcqqdjmxuQYua9QWQP3HDDwqybAU/XXpU9+0VbMWm1xoIM1fJx3LAVZFERqcLSp07aVgkyE
Uxdt0+AtNRROBI4ozPD2qjuFLQeUb9nTXuD8+YjAj/HktdC31qrKDjVV3LGH3+bGcpporJzqdors
i8ZaPWu00eE+OxQdO+jA1/nASmHfuMUPLKbZ5LIAD3wigFTeL6Pn9wHiOW7XFCORSxEtKUuYjoz+
coTz5NNqGrZuRldemhcZ1tJJibNLlKP9uzbLlgcK3aNiiXfOZSE6wc1mYZbbMyCFJHCfWUW+2mve
UKa6wmttvaCLC8eGRzfbfWW2pzqwNkjuOsLPwSVAFbPJHsbWHYBfjLYJys0k4nFvuev52lnZ/Gao
L6pXBoT7pu/pRB5Kfv4J4CoeVHsWm/qvd721dKIPOuhFVhfquDZ/in92Z1TTJAJEquzYXJYvnqO+
yd3BY53EhXBFs2dfb8Ld2h0xnVjXD9FJAJf2ysBMSfh4uUlJjGBJ9W9uZDXQkcLyKSv4UAk02lgn
AGUHHewRvfimj1Wj5umhbyU78p9+ELymcZ5PgI3ucgIula55u+eILIbeKFKabRw9tFPjpxR3je6Q
H9mq6uh6eO2NMxd9crF3WwajLd9NPR0stvmaxYO3YTj4gSnssa6FCZaAEr0Du7SmsHK8ztA/JOFR
aQClX/DxupFOVkQsJ1dZF9qo1ZhiS4e9O/GImskxNt8JRo0xZebDO148PQuChmNJEVCRcYnqwc2k
oA5NsvxO1+rVY4nHDwODsXwbF/1ObVxUoR9cBtaANC6HrI6feq3r6Q9+a6UYCjXwPf8tw9uszB+q
U+zgEYCsFEBq2SPWHAr1Kc3SnlrhsbfDGZTqe+N9wBT02TkVbUcgwcjsZhOxWoa+Ax1SWpIW382a
VHr45U3WUN1Iixrho9lJniC453jHSHdg1JjKFPZOuRKPtQc5ngVrwJHsFQmv7tH7pJbe3qmoOnFo
rMHUEVsc8O4DN3N/y4z1dajG2kErl9S10zOIB9QJ2y2EfHW3J1yvk6PVB2b0wTPrITLO3mvvynu5
9IyDKDi3iACjQ7JMB0lVUJ7zdLUtMxOJJuLed31SdP7EXgmSIN/QCeH0kg8UrNbwryTHEqYdIEoY
jbtMGNcydzTTSb5PRR5B59zl4T4Z6aShFhXXRrRJOb2DSdR8lP6i7m61fzlua7cxYgFoOBpzo1eo
aAtGNIW42NqZb/CNXDr4RkbrSjy0btAFjMFLSx/tA1Kak/0iAsSv4ILEtH2HADdZBCNt1aQ/2IQn
4QMtgebb1MYAkt7cex69d/lGSP5sEzv70G/vO4+QhwcPXnbm828E+oz3nD+CovxrGGYtIPSMQt2F
JdIExpeotjYB7LWWJ+ridqaXaK3YUHy8UhYSXW8de6TqniD3fu7oNugqkODPiredOzC3eKVLdISa
/pEQIOwSYwA8NruHpvE25696/9S+TlRGuD1yqmAs1Qv+gPCvFiciYYIcvj06I50p8t6cVbS1t5wr
gDPjLM98eWlwfyT5jRQDhFy7oNjOnfeaC1MLYMu9/esF4ttVOYCswKbEHfKW/1UzNu/m32a+2SXJ
I0DgsVcSbn1j04mHoer9U5UjJX+tco9s4cG9sipiTHhcbb9LursoZWy4YWLrAcBfNpjsGJGIU4DP
ZcifJl9IKuAJGg2vxJxx2fPFM3PZWYVHc1FvBNaQgwu8zXtqoLJv0rj6QMHMTfHgvsfNeoVL27AU
eghkwP8x1kZaeXLWuBoRvleG1uzGrng48t2BdIsATto8fA30j8n+f7qlVwEgur3WKOlQuXK6oA6u
2IlSbgbw6BgRo9l5dCzGPx3HnHk45UhtZLSydpBQmiaLgjCJRqdYVriJjmJjf1zKShGRgD4j/CKE
eeBU+bdQfxJTrAoQHg/tKjQag8fQEVXG+v8gUe8QEXVGSzrUeYvQrWYjjJg3vkwcLzN7vj2GGrGK
cCHtoKsNrl0O4NRaa2+yPK2Oh57dDGgyJ6uICbhCIqT7xyyFFpGgUqZTulZgKNevcwdl1nrvSzsj
43b6c7+F0ygqGANNTXUvKFyOJcMZ/AkBMtoZ3JV/tb/CWjl4L1KaoIEzI+pktmD1tdUyrjSghd3q
7Spkbr/BPxnDQIuPb8IDiNlUO0OwYVhQGT8RZCtkYjU8WqmVV4QgIOH7DuNEHp2UxhHzPJh/6YXu
m8kUvf8WsxUtzW30fDfFEIfGIumBYe5gHFfy7m8QaVGeFrudn0IhMZhd6gdLQeOM32AEC12zJSs0
PYfQz4U6o88XtQVCey6ePLP7euJDCydFyiUMoxZ0/tNHoiTGXKvq9yjlG26iYU8Ayob++/NzgYxV
CxnGUylWE5/ynYmvDsxzjrNhjnkcg3RdPs1EjhQU3xfl+Y4gOfq/WJanLebGnLaU7sOp/G3m+74U
dxSxiIl/dFcZNMjukp7rnj8QbiuTMAd/Qercqzv/kSxNdZAdBGolBBwC6BzUdaE/o0wpnEdlUKIH
87JAF+vl3jrcYWLRrGeO8RXhwy0dkiqM96Z22HB4Q5ZF8rKpJO9xffLR79Sg8sP+yRMJC9sDTo+k
UJbHlrJNx5yMX76nvArOejeNNp44ItOL9vGfxS64nPOSoFW4pn93uRPV5zEUnwG4wqDkhXpYhYDV
22jt9Edl/dVz4H6j3w5izizyQPDbEy0L+iqWbSVgc4uCWzZJtdRiILz62zp1mK3bDzWw5FqWBXk7
+HtfsG6Gtm+kMPX91a6YiAlDINMtT0D2MBtJ2Mx0gLNb2FmMx3IUrhj+fzAtLchpX915YD/umAwI
aP1DTFvz2dDN236l8wh5PhMzP3Df7oP49XG/h1D8a0fngz747DXJIkLxqVwPrm1HDRKUyyr0bqL5
xWNOEJ7f7ZCLO0WdzbKkLuMLzfzW8aKtkgEku6QlErssVT+ntAVy0lCeNipaJtcAHBzJAzbCx7Li
nzGZjR1J2MEz0R1jcNMYHSZ2yaTqo7SBh6DVUgBU3zZRqjADdt4R/vMm7CTfuFlcvc4Dja1diEhX
IfqMTCB+6TChb8czQvVZqOH3sVzhMvA7G/OKnh69tIYeQ4NUnGFtbLbemsRxgw9JdnwR2JmGx5nG
4pSCJjepahcG+lkMEnAXdyuNdeaamqC2dxThEPnwps01EZW/dH7/vIjIISUUrmfhDDAnkG3vqW53
T7C1dCVbMRv0vsrrsxbLmUMK0trrAClRSuFsAISW6a97pKBNEEN1hDG5DZSFJW7YEMqfVQa69eMY
7DBJ9/smj/qD0F5EU+Si9tknQbYOEj3eO87ovDHFqC5GB1RjAAN8ru6L6IUjPEB5kxZ6pc1iQDXh
BgjIJwHKPc6dKNWx6FHT3FdL0UE0AkXhbziT0iRKPbIpo4k6n2iv29ELpD6PzKKPz5b5BCkard3o
81qgoPaovpvhz6Tnc8i/i/rhy8Ht19YJQ8NN0cGlZ2PDstfW0n2o1daXRPi4Jxvo/e6+uI4lJ+0S
3Q7SRs7lzUKib2E40Y7SfEJghdqTI7qoGVS3W1uP2reR7+jDYW7Ggi74Bl8+RvzyLoSeNpTwrD0A
x2JBPC2LOjFksVqpDHjUGjga1LmTG6WqmZZz+3q0DbZ1+Saxre7NDl1bb5jWofZv3iDlm8bEh2Dp
qY/MYC9m2V1Gf/PHpTioWEyX9X8p80hEWo0Vdns2qEAMEGl8/i40uRfTNH5LDl8IMy2MjMm1acS9
U8KuMZkWo2ah3tdKaWgECmpVLDR09mOjUWmv1CMi32B2TON+2pPC9rl4b+ZthUP22UmkMXUBMD1m
hOELU6g5lrdZx5vhPogwI3w8TY/FhvZoOacJXYrOxhYMLYlbtPblLN7AqgBxSZCK4K21aku1JC2g
oUFvLikI5RlJvW7z41Fq4z8x6X1pB6n0wHPvhmY/TmLAQQuyGVrr4Y+9nxOtVXXQfgk6VCWsjeeA
rpOKzsx1aEku79ZbLT0o47rPJ8/76/d3sa0AOOnE9Bd4Kjlvo3lESMVikuH/AjcqPMuMqZmeGeim
G13/lf5ZNAv0KH0//o9feWBO4VxHHPkP27ePE3FAqi1tfgL3GQ4/cdqPdwMmCYDsYhCXSDTUR3en
VpYzR5cxvgfTc3rlD1lE11P8mGSHZ7fWDcbS4plpOjG1bx2S7J4KmNN1/xFqlqEczldq8tVih23I
Vs/7z0yyah5PkhpX71BmF4b6n5IBNcxn5ROEkwkwLQCjvvnjn4URjY8ySE3PNLVbvJ6TKR1bF/AF
642SiDptqCmHmswHpS206ksWwAlX30dmPAj2NderAj1ATHunQB4Csmo+F9SeentpfNs9rpHzAFol
mahCoBQDRCashqUTeWbvX++5iIxcWGRrZ9XUSvN2krYqqD9Abg72J+42QLCooP775VbeSVKhmqUG
lJZnDrW2EqAPFv5cHFCt19snriNwFhB+yXRpbKTqsZ5AwLkyE0CEy8lwJC6y4yPiXVndEcdPD9iS
vk9Jm6UOLwMk5CRLMbLcoT300h1gJh5d4c6yUPy6fQXHj2dt93914Gt6AlxVhH0dzVCsrx0qCF5u
mlDCwssvLMwltcE4edFiuv3iRB+q0mx1MjCWBEGHxH0qjRXmsD/R6ivssi7+Tk9XgIji/mN1i+3t
aCH2iQHZLS+GVxZSSlA1QeTsBdBS4CcsrHAGXb4T8omvyH+xYhMneNQ26h6qHRPGlsgy31Tn3kBI
lpl8vIVF73BVLvA4Eu3gnquSRaEBhM5VBL8kMY2Rjex3YpRKaX26gsXTPjBO0fPa1Yk/uMVzZKDs
catLlV2npEojKo2H8Ljg4unzrXcFJ52k8AJGg6/M+1EJBgUAcFVbMZseYN9jqIyniY6Ta5tbFNSj
Za8+RFGXmOmOcCjxSejvLj2QdN5dcsi4EteUpC17ucMT5ZA+a41869A+kWZQ5AHpP6gk+Lemunmb
6IjWZ5bouAOMJgXzx5aDtDdKXbKq/BB4C/Xd7Oe354Hs13ppNYsTOkhQqjZ3uKFgE55qluUhISBx
gHykaDIZBFT//Hn0G7tg2Uz3BD8trTso+7HOecX1GGnGGzz0jVJuf1uVvUWez0mb7Yl1zm6f6Nl/
BU1tNldDGBRLzY0wWwijZQ4kWnSVagFMggl7mAmfKkV+eL3JMuF3hIUiBwbXWLusDte0JlaAP+rM
V0wX+BPhP6sxgfZuk8x5lql0zO/BxORz4x3jQUQm6T2reOljKOfT5lCpG9Exqed742cbD42Jd/KG
nhxCS3ygOwYYyqCauKv45mf7jezfni4K657HC/qyyB0yFGxJaTAuiCU14yXwCZ6dCGBa3rY/tIGy
hVFLFy3FJ6iVTCtNTquxZBoLfms7VjIJgVxS/MK4Wq3bAnIcE3n62e+tDPMMfEbqNZsc/BMrjYkT
ljmvbm9Nu0yevblmegDah8us6O4xOh16GwnpAWWCXp51Vdw+Psu+U+AZ6UNoAw4zLWM5AuGBe9w0
AymerN4FiKLEE0PzFskUHAXb2eQaDn6+42gR6qBF2eOKNXswIbMwBeMahWiqnBdFcxuJEIWuuSJq
iB1N9GLzdOHaJcY7Rfy7XBk+FKS0fkPtz7bLZk18IB2a7qC8kdJhHWAj1/arYk0tDQ9Fg2p69MEf
c4CjsBspqjKPEyVo1JJwMVd2nzE9kqaRY0I+LjTBlefp15/5/YuY5GP5oCLFJkEXR0CQXlmK/0f9
QmpyYJnDSBIR57nM4ZL8CRR5kxSMoTqlMN6csOk0WpCAS0qBVoa67cnLekdNjVm/QvpPIVDja1tB
CTuxnUo2nCzhR8AdVuFTU2E4vXXA0qfx5oHgnc10Sdwa39nU7tq/AEIR6M+87dB11z7oTUwvRVin
PJkEE3ScMEtimn7B2TDjU9RqsYkj8EZMMJXnXg2/JyNACi/1cx+enf0qj68rkmIxWYe+vef8Sq2b
V+nBvrXPCX5O6fGdrM4SYaIAMAyfve6rAmyxizFQlkW7ltgNMRDN7xRcqYk5PY6WgqESztngjqWE
aBym+w+wGjIpungtjFbXe5oqjCwfzwcLXdRKJ5qHby3vNs/ytG5ZkQJOu2ISNNPk1coidIUYG4s1
1XKaRxI81NIQGZJCGdMRrmBzO4frfmbqSvY5T0cEBiLo0CUj3srLlKutok/F1dFoz7aAxzUtC4D2
seVRZNbHTIx1Rfp6axsq9wbTczIEsd70mcXVzJo4QeaMnLbC/wKnqiskCsfMShy9MC3qJxoyl18J
5s5VEBQoBCDconJ4C5GBw/X4FaKiWnH6HwPG8F5BQ3nWI7YQ/WAgAb+7iRZjwbpnzHGf915qkTOH
ILM2cFK8BalODH6XZCAUba24mEEd9qn2CL0yB7RgvhBcrUKNI1GJ8uXZdsWTWSvujd4BysMeJS/6
6d28ze6HqGYLu4PK+bXcM+Y0kgvnHt6RHkc7ZI7obB9hZO1TzBsyX8kWjEpp5DtN51ScBxWxED+f
4JRv53IE18QdW+oDtaS/aBSgS/kRnrxMJ1+dgJwM7+VS2AChX8Bbi6ZUGjgVNJkCf/dlWZ3pnPcJ
tL++YSut7R6MLjddz3Z2gg9IIXl+iylAJHacVxe9Sp7lBFgHvRIo3qZMnoAKN9d7fke9V4jemFIy
sM3QRD84RCIHsjg3/CJbSq28W9MqoP/stsDWD9kBpQLPMIfEIwj2Hft0ibvCWZ7nSIArUbPQfU0V
GiMoiwkca8dkfeMBYrTCRYvZU1lYdAxBF5a1gkme84DJkAFN45JlAWeI/ddn5UGW6FOk37lQlu0A
/wwQ4Vbf6PlYgibR2RTJlRw39E0eTtmnz0Qfoiu1Lj6ODUsuN3jxMjsXUUzw4D7qnCPQnQgqJN5H
Cb8lwYLMhhfoOHgbqMcRlEc4GlzLwHazFzToPQRUTF6fBxJERV3iu170aN1IR4KuTREo20jcNKlc
MXe8Dhl98OPNPBFIk80Sto+SugRZoMPu+NI1W5ne9IzgDGSR2b2/5cEjjnQjmggoXAd5xlfTJoax
Fht4odfX3gqU5PWOQO45KX9eUno6WLy9prWQI4M1RbtOhWNWdsYOsk0DTh/vpPJu4mZ7+ibbLybq
kWGC0PGf73YieOUaWXIkBWiajUkncFOkhb5VwauLpYf041zTGL/pcYXoeEB+XS4FPiiQUg0bF5mv
KgdkTkZ/lSmuZVdHJSLR42imrYrB1KDv1WBKVdu/LJU6fqs5npSsdJ+2PJCdz6EhoHftX8fcmsxt
zib20+6FboRhzFH2cVWRWDL2owxrRBcQqVrctNHKrtZ/LJ23qyYpTDhe3KRN6s3nRdddoLTayCFf
nCVgrWAuMiv1GcKUC7bJ3qxlKZ5dq9wvv8CFMpX/EIoG7m/u4OLGVEROqb8KSFBOvq/75IjltdLK
5kX6YQZyh8Tsd5DzIg2vpDkf3m2JwobJcjTI1MAGnCi13KSXvhdj8Rev+L6zExqiKV3Af7Yefk5I
siRNzlgHtZUiisKJS4HdFFCnBmBGIT91HHS605K8iRuW2Ed1y6qok+sDj1eyVRY/vO2wa4Ki/k/t
c+UyTOiD/I8SVZ6NyFFRpGNmu24b/AaJxXAAemu+0sWtrUVzD/cjUx5avhv26684/fIvTWD5qJw7
N0hGwhx3U8/9Y/otZ65Svy75qTWRm6vjmwDqiMOReicltcRh6FQ2WY3zUj2yrUXtYRP1zEPxr8d7
/cm35Y8YrlB2zqc3b7/y4yDU9K0IMS1kmQXyy4W7Lrs23BIzsNQqr1xkQ9pRqB2hvp+IfbDB6Q66
wKqgpl2ECGFVxGN9GjJofb0xi9Oir65gO+S5PzEKFKXUphiQwt8Wsqd2ZnmfuGWqMtQhFf86jBzX
nx0n6RnuogjkavzvqR0WFgSQqN8b02heBE0X75bbJgHyUolYwSt2poL6mmTFzR05C4szLbWCulOx
Xpjw9DZuHj1qZqSEMh2DIQdZaJbO07f8i7F6kZQJzjbbgtFstoYBNLndboi+1WRJkyAm4HnlO/gw
dZ2p4q+Rq6jNWuAYXOMpIMD7y+VprrUMi+m1JwTNUZXwYV1WEiOtDfCpgcybmzbq7BWQU9N4bEpF
PtZb8s/O4k+/k2bUlAmvfpFSxMWPzIyZY4Yi5q8Qy7xFxAidAZa+pLqP7zfP7xWWnQl1uDFvq848
kaSai6zoFMG5uCjJ1aMc7CicKQM5r92JQHnGPJFVM9BBYn0/G57HhlerXWjZ5MywzbrCQ07kdd6P
3XN+bZzntX/Al8X3nA83gFm4PFdBESzyXbct684pS7RZXGhGUA+P4znjLhN/9+/7wBZov2oEEKvf
9iA3k52UddwUOHd34iYR7r7o15/deTFqTBd9RCQfZbIlInwywhQ6ojUgNgUH0+aJZBdhsShlK7Kp
X5kVtZ22cgDPFgrlfNsAj4hyP3P6ZDGAWG3woD3X1C6qwAs4AJAeNPosXRKuS+8K8t2J+/teKtzC
LgJel8pQg56IcIkhP6zOcoerGvSdOIhAZyDj0yr4x2YJDOyy/MOybWYUZvtUXnvm5wgOQ+d8GwTh
r9K8vdBKcpfJvBQd0nDDX8wxqkPHOI6OpJJCE4dRN/JS6gKhl3amwMahEwT+7q9Tg9Jb5+ELwHUn
/wM6KcXAXqdbLecAmCAS/B2E0gEXr5+Wj/l+6ndHmV8KABF8LpsW6/i67aqoUTQFZgMzbFt346Kl
E1ELi2TvkRtbvezwbt9aVfQvGDDukZw3wMEpn467IA14P1EmRDr6W4VLEiQ2YakBu0sL9HoI+pFa
RJ7jMw0nnVc2RWZEdWK3RC3WnqrJNCyythRnrkfH6hE+W6Af1D48Hy9PQHMzn1Kt4WS489c8IVOM
X9Hm9xuHoUupQE5hnDpiWnkx06XVSbof2OpgMMMPD4Gk6fFlTdMirZbdki658N0cKW9r4V482+yT
qmWLILs1273eAbSeYpFxJIkkkE+yIz9o6ytMr1+ovaw1DFceoYm3Z++r2e9CQVQxJJzEr4DdgD5w
4uDsuFD90s9FXUTVF6myKdxV9oFg3R7RKn1TYtAGMqwFg9nqADJIvBF+197qFdA6HYr5RRvWrmXx
0nJMfGf+BH2OInFeVaN97HM1Eip7D4dhTD+BSYOPxUpc9vlVnIXJdrTej1FSf9aRs4FpwSsDwyPZ
PZwzZiBDjUxfgrZfvily73AUwnvWDpCNVgJt954EYpI6TT//3jIXi9Sw+xzUPU9Wz3qvLAvPfQri
kEM4YuBk98ROYVB2P1bWt52yz8nDvg8VVjCEcAtg/k+My60mRsfNM1DVZaZOM3eBuDzx/8d6JDTu
hgiS+Jld1t3M01TsPA0K76ieYOnaTRbsDZZO8XcRWchqob+LMsGFBWf/OGa8Z+R+l0xcOX5s41IT
5D0SdpBr9afCJ47DnSkfbpMYp5MhnVXfq06PqoyWhk0hgGCYNmEasb75TAoDI8ovk0fqSwC64F2e
8Gadx0kk/ykOxKllpZ1OxHce6CHlSs06C9IMm3OPhkRxyE+P9q9POV06XmOfGTgad2L40Cfygflf
g7GgoPoU+SXXssxc1iN71fNEXquL8WHC4vfURnctd17dBlBSMiP63ffEPvRovgcoS/eaVt2xmygg
gpOR6ZAOFb8IabAZ+qGYqDGP/VjJlytnpfebRXbFtb70Lt2Qlx9SRtwdUdbPZ9c91pnRPdzzAW4B
pUGQLBYLPvDVP5dt5gV00UcLXfn5qAI9GbdvhzOfKA5WDEVY/RIaJpn4VYBbdyhgREFmoWmxFkx+
VZonLPaaQUmpZWpHtEGkd1oYyeq1geGXYQ6E6+Y01M7W+OLJNb0pKfDehacOUxDciI9E1qkjpUz+
eLIH4KiyzQelbFrFVzWpOITFcKXZCjKdOs9Wc/RlUTVyoQUyTJ714uOGwEn1V1qmEQSsBL/eQibj
hQrHTCWQIX42PNZQA5FRoEeDkjyyL7ZPl1ZAAmN363TDV5nPs6LQfSHj9biq9z7IC0/VsYH1vghS
myqFx7ZGMLUHFFt7IbgfQaLhIocAGKmea20zV4WU3zIjCqVaZC1mWSNfdRXfSnmYfsgxMBdssCIE
CDZGmm8GM36b312Zpy5Psp82YiPOZdxk5MMMlXMh+IlmuM8LVvaTzmI7DL6PyBVh/dOMdz8bWqXe
cBE4DXfYLUR15tOOElurbOPWXf62HXmc5bj0JSYQzULJlaY47uhx7B0g8pqqSTd894+LVw5Twv0u
n9d+o0uCUo336geqEPo+37+CoJmjGCj0SIdT7CkqQxdkAmbbvp6ORKaieGzT01dhgyR2NsZx+4vm
ZD7Vx3hC+jTOK96aaYhnwHyRrZqVgEXrzsZq3jk4gbcgN+giK9MHuciluyWmF6AmoPewvzNrfJ9g
zjFSdE8YBQRj+iwR5GYH316Q/Q0THeHMGEgkeOwDT7SmA8ctSu11FTwfq9sm8wEsifgAkkXKa8XO
m5+AKckApyq4o6XjS4DpiVPko8y2c62rj5EJE54czdTga1l+dWiv78DPUuCH2+eBD6Y63Kszsodp
HlkkkxGeOgEuQmqbxyFE3GbuZucZ1C5H5AtlM+neeWA0+okFYIoWgbFlbnzehju+uEWlqEG0Lb9p
OC81IVwM482UMZmU2lgVOyWiviOeYShRZsMA04M/U+mQLkkGs403ThbUNwOB9t/mZ5Pn98wSEXE9
cK/W+arKPdyj98KruC+HNiMC2gyBM+I9TaFKIoXlvN+5uFEAfX865GydDyqzxFwSVCR8KCbKqFre
FxZocUyuBLj9O0pAGufh3VY4dYkXtTTXNmN+1KiSiO5q2wzFCejPg4+w7TDuKEAx3KRkTTGVq/81
EEqdDyXJp2mrhJAukw0yhRf/HC9PEwUI3YhO+PiR9a0HfYci7WjUnYTUdjP9zT7zPxfLrAFwAYG5
cG3qk1+NC/8guf90kIsXmxvmxV6XYwPEMWx7ZJzDND+nCXI5BhE4l0dIkUr3n79tBcfXyEwc3jiF
KqDMyjPD7cxhXXgX0AwQ5REeRHbs2qP+EWUJLYqIJgwDfgClM67bvuhxXkpJi1K0Kr3pB7IOpbsq
csX+hCGintSZ+tj+sM4XhT4BULH7mw9hbzITNQmMQrt4k9qWueQHQmS5h/FvTNGlC/1TC6++5J5B
QaPXl6Ejs117pKKxXI21mOk6gF2KZbd7pVdciT6BVK0Cn5tWwELA0KFHndu+XvzvISuBHo/M4+77
yc1jvYzd2CoeRj9BC8NLg1nLtsF15kOElyjT2In+j8QSaEUePyd03QPZLMaapKL9ZSX0CEUBgK4K
GdNO4UttgWuPzw8lUycovobEmFZ6KNKQe5Qe3jHKpqWJljo5WWs+S2LsSsRf6DTCAFKb/k4xRImU
3DR/2yn0sZt83JJwWgxje99j8s13gcG++eL2J5vsc8YJijif8DF94zy3lL3xZ0s7O5ChxU7fo6We
+My0LX4yrq3bDQsCpNp0ScuutoL9sBETJlOheP5L2fufjgm1CdbFGY8YVJ9Dqstf81p+37RvS9Sz
xFuiF2kWV2WkLDvvJHwxLdvxCDuf9Q9KBLQpRw682joA6AoNC2JU3JgEOY8hA9KTFr7tPoQuavI1
+p69MfBzStnwgLN7ZGxP2aIwccg4Z40wdb08vRAOc8czucLymOJkTOMmlgT937kpy/V6lCO3jQEB
XdFmVUMl3BdXSwZcany1F50fClcHRZUs/iwnXQPoARnQMJ+5U5l5CbfO+2bDCFDpIkihbN82UA9C
Pv/QCPK5EhdvvNYIpjlpkv03DRd4HyZmB91OqHWdznzrEm48iRuI44pzNhZYqFhzA54t306OYRlD
jzSJzP9TKMRcMBStF9rhldkPi8bgam/NWsxxr2byviU2m0wbarfkbMJ2V0SYrvVHii1PubGKd4wH
ypnZcis7TQ+eTW78qPvN2SSMxXZ7S8cZ0MV8w4cqAqhKWnY7SXKUTngV2bczIBpLap+S+Ux5qwj1
z98Lk7gBWQ/EKiXL/CAi6dt2qgtlZ3JMbgXM6yzpexF3f49gKvJRET5fdIbdpoRu+Ea0vym0JUwp
9icVQonn0qzuKtLTe6sMaVyJ+fDl0gMjAAPIy2NEfsdgc3JRaum7wWJk40xkWHC4DE/s7rKSXzby
vAjbFbj93GzKxw3z6KZgJJJKGz7vNR42PcYf+Q++e2aZ4IZhDsCLhcvE4zCMSpz2+/40ybpLxW+2
L3uXIE75kE9b2/3RE/uDoVrQPtf8MJqbkYLzZrqnZKahhMBW+oM+0kgwOwzYKY6/j2Uv+WP0gV1W
DD4nW7XTYyToXkdyzjJzNwWu7rjbEd2O0hMHlLgcTihkKnGVb6WEHs+bewmq1j/DV7lpJN2/NQNv
EeygsEpCwZns5w8Ur99rSZSxyrJpSlyx2gO0VxVuqU2Jky/9quWCNCmzqiFhMzO616Q0qK7AF2pL
QB+x4O0CdzPY1WUmtEMnFp8qaBdtINKrzc1RXgmOH3dWQPUZXylFxRbD+9Qy5NHWOBIBff8FIwJN
L2h0o9dwmwnaGIV+KYKpULrZqhIzlO9QJkbYfs592uNLXqk6yqQTpGryFWTDtt7Z0PlxnKqADaHH
Y4tjwjBhmKAWqHd/6+8ivSFKzUIDkoswbe7gLTTvmzWHwAlPoTZgX77lL5Bv35usHbFloFsfpFmE
BRU9HvLe+w8GSd8aSMU6sbS4rKKbnmrdu2Or7Qe3UqzM1QrGcwITOQwxlAECeO8PHNipluUi5NBO
PujyyqWTQ5zpbN8SRJeHkuGd1PZ0vXQ+5rQzlRcFQG21fQkSqwSJxPnuOM/oOOm4PTMN32T6JrSC
zUJ2LviDMQmJ3tkeS0C56eCJUW7SlBlI4G73/8sywbJrvDbzbFM/D69mCTP/GeEqZPtzq/a8mrZ2
zd4VemjWumCKsXZriqBZ75va4NaglbvCwFmgY7UvH10awJLFCMNFrNBW7XF5BBsUwJ3ngujz8CqQ
4enokmhz1iz1gXakfXWgiD9Bp2xo9pRs2/d8T1VWKM0wH5lejnsGLaaaURN4TXB5BegUdJe2IkTD
3hoTgqxyykqdouZF/0NFsdqV5I1A6C5v3alNAss5e1BPbkwVtOJDYV87PTUvKEBWS69dMntJqmVJ
pEgLHKrZVWy5iRNNhmIMmcSJwusBi8I/Y87SPPjZR34FjcvdBlfXOdyU+QOZrqAB/A2PY9KIFnVm
KPFDpzohyQ9a3/IGFSxH7hBI6gkrIouze37daJSgk3XjNH068lFNluA5SQ3XsSsfZxLwK/y+ZKRD
mO0V2dM8bJ1NG+xtq5z/3rJ6km1y9XHKOJFoulnPq78sDACFAR1WbmSPP/QrH0aXDPLknmeyuC27
cjWZv23BU+TDMPijjNsacRDGDAWjesmhUHaV3QN+TUtFcOeaYvileyX75PILRxqEr1S7HdRoThao
9rRauDjU6EG6svX3T2qtCnpDo2RE96At9tyguZmIRFEnURZCeSdSiv+9JYQnbHdF9z5XCqPr2q5w
H0H5Y2JueSZPNYZeJkKzTAlt81DmVonjbryfD9lUgGj0YOtCDTtCcA+rqwSQ7FmTzla6HNRr5rAs
HIKdp470XL5+IxYGiJBP9I11Dp2rE03OBLXApXs52gH/cOjLkMxrMkuTDWXVeyGoQOq8KoUd6e5c
M2Xumodal39fAeANiEevK0CdMMAppgflk9aVjLet+sDCJ50xaqMZMGb910rvwDiGOXRHCOK3C+IQ
hrGFNdC1CEVtQZ5mEBbm6oA3f50FiCTyncAGuKycuKT2iqE/PkdZ7HvUYGkxV9WFiPAXv1g3Aw8B
0jK2AhGKDpVsuUb/Pe/vh9rDYv6jFbl08PzAtsdrvvfvkwjftGF7ZYd2IwqAekNTP0NhbaH9hpHH
u9JQ+dMjlknqedZSKQ/w/Dv9dsQqxF7/PqU8Ft64Qiov+vKWP9Zdq++Y57ozHBs400aRKLdxdlFX
Lz2FLzpH+JycF89lOoHO95UTFTnn1DsH4dAl0x1VMAF1KZGdGyBrXahqBbxKHhFjubjpLOPco5WN
0N860I6Wx799DCtDMZFg6AEvGhC+vBRHR/5zmsOfVTwNy1JLh84/o11o1X1Z0+rlZCSKln/clHuT
QGNQH5oDSJ4/z69IpL8V6Pq06NhO/+eevSP7olD29C1bdToPyp89qzp0i/nA3jLKdcTpgHrKJOJM
lIPQ87+mIInRGJucyLvSTR6GfiUX2x6EwJumVjSsIk/vjUzed9MoMzdQoUidqL+SN1h5vxmQWDsG
rLZvn0bniJqvmAmrMY1SGCfKN/DqgQo35ujrjSjdd0q3N7DdPxN9mSrWJPj3IlMrWqd+sXoDHcDm
m2S24WRr9ipCUfzmv8XpJhnmcB+PVGOUzANpf/+Xr/hIlCJggL3pRSdN+cbQcCBRRiXCwb5Ifyq0
dr81yo+7jvSNMB6aYO0CmNSAmUwmLKof9Yh6xSOzj/dtsNExWPY9IErxYGN+p0vYGjBtW3rwu32g
6ERvSQP9AxLjAO10x2O/pqfCmksXxDcuXcik8sJYuEDWPxbhOMlsvhC+uTxbym31n6fYN47cOQ4z
pF78IZI1PrkZ8oB/Puo0tyyae7X+7QQHx8f0mqtaPzxYIS4dBYNWKWUqxLxhoS76Onng07fZdTha
Fhqaz1SW/pVytJc0LN/jc32wwJx6CbfDFhoTYsktdcgIB7HK269XGlQuKqiKgkVlEC6+KhbnBzGd
mIYax24uG+OEJBYXmi25ZLl/ayPm9m/g25KTMP8vV9f9NR5+KxPe6iZyLz/73+hZYxlrZ73YtKnT
AMN9PpvfnytSSaIKITtZwPwjDqzLdrd9v1RL3mwD7KCFG/bw79N3KXYldqkvtViNluqN+z9OE4d/
CXa2eexavHhrREaFfssA1AqauOFYKZhLc29kfysa4UGgX2koZwoyyfulMM01MjzAYiRfsHHomNzd
qG0WZTmGP0r2ciACN6icdcOiz/kz+zTXwjUvGZx6i6GT68wjHHw4YW1P5yCm/Qlw6n1ti0OyvtGn
w+oaP7cFh4YbhEQsSwaRiJIKFrZBPcbjKV+mNxVYEtP1toV+XDA0vJW7xtmryqm3ej1yXd3L7fwq
6iAlAeeBR52ZZkOM/SImPX013pNTjqe+mLIGHtVndamJ8Hvn62ZImufexPDz+ZS9+EISxOHeXYuq
ILZeXkKyD/eexDCIslv7B4LRX3YRMkmke61XhZWO0YSuOwo8kGAV4px43Lk7wDe1zkn3XVPq4rjS
exV/TSHoZ6E/l53eW8KfFIXxSc2HdqeorVOdQvTQ0npFJhA2VoNEUk0OokgO6iPM0vE1zeDZqE+O
LqhkuOVn5Wl0QSPJC2hw/Df53TvVhECR8cd2PTcaUbF7CWWRjIcf19hdKYdfMS+NU1IeksGApoot
YdXx2HAGau73oO6iZLBfI801TUDoGNPjNduXEtlFQnwrWbFITsSfLPgaOKQcB/IeRqeSqcEH2QiX
fPMGvLKWDwWmlkW6n16XTM08TFcKDbsmvsn0ZxukhQRuuldQsMXc9K4mwxwJV4wpTxair9LOxE+J
zI832VlX9lKD36y6ueuOEvl1kSOUeINKjJ8uNjz3ae3e7TKy9XH/x0TDoarLbKW4sZ3vlSNZZnR7
iOqPw8uhyxo3MhTI3hqaFMrfWRqaixyH9kB3MTys++s//FhJHWHEcaWaH/9cF1aA8oR0BNhxrCGW
LOdw0CJaAbm2FMck67IoWaq2n55FOaLLHI+oEKfKXNhkVdgpXcO7Of+RP9zS80HnYC+5bhbhqw16
8ItHenbbgA60Dmp9ZaxEiwkvgOYWvY/GOx4LGjDhV/R0oSnETAgQagbSBy/mcqImcvplRsp+1LLC
o9z2KV0h9FOi3lZOfKnvmZFKGeMjrYTj4WueSZrcIIgdZXesPJps6Da6c6uxhB3Oz3lHr4wKiGhO
h7g1rezAkT1UKy///7uh/9fBfPGXgHIDdYFVHSED4obVmitB1UM3t8kljEE7w8Cej582Qjq2fpLw
rMceP4le5fAnCSYW5G55NrLYWhm+5VuUryGHmj+ANACOruUlOXsKH4EuYAlRgDCjIce3MklQtI5E
atHGVRUaL7DC5iGaYSUgiIr2xAifxLEeMTaXEOQ5SyEZNUkJoKCDctY3emtZ3Y172t8tVmFJG0WN
g2BKPPkUwrJ3Vfep6+UncFKnh4GROMmy03eWhYehwCrv4HnkgK7sgbRcd2pc1wnRZf8adVlbkXKi
06I38lQMw4lo27yG2R5Fy2lwkeicvphpM1enKk17tlXPqPX6JtSGVPKTvPdXPiguluB/+5N392j9
/jNzatzWMNgUHPuj0VatuvBcxjoKcX+HfwNbh9rP91hGXH4NwCk0RuQl0MnqprHDwIdMYn8ql3cw
lZ63vsSvGB9H3f77iWyG87jvBNQU+TynQxBGhPUZLb7UWfiFY4sACrT1kq2Cw6qQJgoqnFTz/lPd
efIho4TPGZn3ZrGThKhRh3MYftWCc43aznzbdvfwVXTsoKfzp+dEqQR6LssiUcEhrkwqK1R8LIX6
FxhKBmfHf+5oFqluHG9p+viPTgnAU18B7YuRMvH0SfcKVrKWmtlZLOTzf6K+xN/EnJ7FVUOaShB9
bQz2LL7Z/c/7jaDoGXcmRWRWfjkyISGSV//Ni3QCNIPF2aQ3Nw9EzVBTrfxYd0Rs7KagdmZyjycn
qJMCALetKCWBlh44Od81l2JDqVGzT/qOVlx70KwX/Bsv/oIsD8/5Z7Xvgu/hxYTLTcKLHe4QuWvl
itV5qIwMhOdritVeOtzVHqVKBbPVFAkbWl9f7sVE2lOkmhEJvH6Kg3uh/qXo2mW0wQTmsJle59Oy
zLb2ef8Ixw1vno97PaFozCrF0ctSZlEsCzC+SKDwKv1sfIF0ZdyFgu3f+KYkgh0tBjEoONJfr8Vo
WdAaIWNKIWLVyEaQPbWyt2XLwvZ3Hf2jqLLHUDIPXMYe3ddXj3E13y+HPOtiwTg1ymjXdGxqpkJu
VCYvn93Hu9HovoeBPCedQT9YfBwANnKsAp42Kj0+zoWI5q9qwuZfSQxjMYpuvkaBgaOY2U8dwA2N
CUYG8EVDegBDKo05uHEDA4t/y/P4yyy6pk4toEOiIjUPgVKpgHTn+S1wM6LlDysvo5UHTCG+gYMo
S9ZGaqrD7ORN2nIDsth0CjAer0fr1t0ob1U0yLNHM6U98y38+CPkiB55pYGk3leaUulGe/ofipYY
HBJpXh6vuUofzZK4e1kjw1rOaazaNmLc+c0lNOz/zm54ztjfDiDq7dV762VfmROm9vg0n/m3XxfK
QmcZDb6EeME/D/+M6rQDW+jirHYIE6dApK0XXaeDtnw7AA2O6FO/4hwwh8jfu660hvRvjjheZFMs
vC62e0K+kT6UIPqMRpYOSDgne6VM1PHUrZi0AVjOqCUAY0IU4wikqZN/US+JOIIzUg30GrQ5mtuV
RfRRMm3bGQJIwAUPod7WtGY6lgWkBgN3J6kuX2VNq0jG8zjLUbTBIojXrlQ3eqVdErrvXCI5yvut
L1mDgoTAvD8ntH0T+yZvUyEDlXzFYJLQsI4kQlB68a+VGYDE2KgpdpwR7mKAyT5hMMPbi8zGbI8n
ctvIwTG2BoBFV3JTBYKFhCYvFk8uz7QqNu6inI03Fe4xQ2KpEIRaLg5YpkZTgDA6KUITQ2mlh8ay
uudjUZoQ4GcVR0SorKZ7SfABPHOaDVl4evhh5tuk/dOF4iUg95bAZtorhuqKnhGXDvAddzjkopCt
kyLgfWugTY8eBn8xgQiXcNaMR+5bpIRveMWj52KBAZRnJfljzVTtQLxnWB+NTEVJ5ZGKUKVLuLsa
FuE9FHpu2XvkTs6dPKnfDdWJmm86l5RaLEZS0Cg+06+c75OWvf8aQOp5QLs4AgzBDCNPWxH1bjd1
L1zqmnqxth22uAWPmgl/oB+8T/akQn3OwdAe7aFw6V7sTz9u86jOlD3LB5urA3Ev6fmQnOYPI8VC
Fhw7hqnTKspSkN/zlWjX5bkmC+rGSr9Bd744IxsWD/0ebN2Agh5HIGaeBr58V60FjxPigWX/K3e2
WETAN3dGRpf9VPVgKDJriyP/nS1GRVRhHZC7Zp1bDtDhV4eM4Dg/kUCcpnB2HzeWvhf68DDULVmA
haWRbLXoSVpLwVujB6Nh8qK6vUA0Zboc5Q2/ZAPqWyIjv/BIzZWRbew2y3vRqd/zLhMg6BfJSVPl
BkjiUsJTrRoUAFbMU0W9/FEU+BiKUgQtk9kKmYHk2gjiwXAVp1JXBEa5l2R1TxST6R4bx64SyDrm
UPuL+aMsV44RHlobH3BW0Q/ROn0EwnqCniZ0suPhxdE2cAC1gSnZzaVQE8pC9ZuMj6ndnRjryjsS
vKFYhQ4RbRM4WcE8w79ZZJGv6kYDFiUJq8GhJ8yv1PiW11Cryuw0XA4PsD3Kdwh91k2HC0hySkNs
TzNxNRsajP5DXpKqZrMER9OWDOphPQQ4H9OxSsFo+8VuDVFnfDaREEnvB9K6/4t8OW1ZMXgE42ze
agdaC7AK++iHLCQKjP5OTEPav8y+fphLmUF2MDrP0heky0R7ig2TjYMtMwKzQGxo+lhvDQJnbO7r
QF4cgTTJDTzwzdWt53NhMX7yPQBW4MtADv4aAJO1hBEKQcWZfMpYBu8rMu64Ef0nu19Hve/KrdHm
NpIr6begO/2DEfWGxE4MT39SwNBSv+9CHK9ZzOWvjZTrfijU+K0YmooMTTcVy8nA8E5/utCjv6R8
GUrwvC+L+dgAY0z8HEHgyBUd+wQuK/fbt04KABpUgXLohSd9C2lpmTQV0F0uz61IaT/yMaVZb4Hv
Qw2sBoXF3OQ/lbNXgbrTgxBZDWN8irYQDK10pLbo9wK3mdAnjk4MV5ox4JsRr+6yEtpKBqRf9ble
S/hIYxU/eieWylTQrCsTGJCK/mYCgPJNKlQ/gpz58ypmQd5jKCjbMa1m9MXrBaUnvM5WhIJZ0NF1
S/lYy8KOsXfKR1i9Ef20CzCWpla6s9JxEY3EivFUh/GyfV0Jv+Py+Kto0qbsoxEP+LQJ4n66YQYp
isb76TXBaJppmLw2Xy1OCeZbSPpSUZ/+6qi/8nbcKrN8HBEpAGWgOliY7OoaHH/BcDnLp3Kji9o4
EIEesFQDnE8+bp90ivd4XKUaAdFv9fdc8NgU86G5MrLhYTjES6R+ltRlKDEghKTB5IyR9m2FXQdz
zerq5n2/HD+XEigkZr20pK9NWcarIJJYzZAp/FGlfi3LX2rT6CC6VIaxAmP498Pja+E4P6qMVYgz
LKNgq+3ljRUWSN6O0/quO45rBtON+KPSb8p3YZqiAipQEV+zlH1HlPPksdYBlvwFluU6Tlg8Z5tH
L75y/p5Xy6SnQRqopluNfDSBsjlZk3wCWU+wfGEXnnFOy5erw0py3ygC/5KItjvp7pnaVimEUe7J
EbcNV7L7MEUmsbCtI3IHoRLaj4i2JMHHM5jD+sZ7MXUMOCDA769Wxn5JBdoHM77ido0uL8fCivMM
Fhdgi3jNsOuRDqmA4Dmjo6zSEX2dQxgez41AYrsPlBzkCaTPAXJ6XNn1/N8ewaRuTi1KuEJf28+s
8DrduxNWGtFf4NnOu19qzPQVGQL8EmEcENMzNWrs2z1A19N9OX2kO2ADN5LeQusOFZqTucgoK5V0
NNNaqIgNMV23vdbxkjpIWRJ8Rp1k3lIhTIn6f6yj9gOxvH5NPEZLmYeoQ0b8f2iejn2q3rCSECil
S7gbdwPAm6Q6AtsbMtB2wmzpAw5ZYgWKmmn2XnH9znJ2cuVmruEAD8O4r9CCxf+Ojt2ivNB6BIw1
YPki88+bsNF0cXX8+FIBFJzwT5CnwhVS8zZ5GJbGx2yXnqFn4T3OIGYimG+8BykvZbSUg0BWgg2L
Hu7NtL5tXKpqxX3KbteELyLrSYUD/OfOKlcvPPuIciWEKWpTGpcHNWyP7tPZcQPA+Qp4FkcJaj48
GYT9X88TDmW4zXdHO6iMFXxFRGXFaxM+08hDqCZOeDwJeDciDo3WUYp5D8QNS2BEha2xvzN28hj0
ZuRJpmijK3gbBsu+QdWtrOej6KqddoTRQpNEbaZb++Qw+MmaTGAC4n1gIoMlvSl2SXMejFesgMqZ
tf0nlMtj6IfqbUeX36mW/0uCllSY0oCFHbvnJtnVHdIAO/DsFNO3hDZabCPJzfQEjGKIZapgk+hm
8qg/ToEfP9AGObt2p+OmJam5lPN68wrVTDxefF85rvcskdTHZuwH2DbymJW35bg18qhUeHsQMOc/
thhvFh7Zgx3AgYxF4Hv4AA0ElYa6ZLsK/0rJMd+r0BRwO5idfxe3j2mMLP5U5XbjemPtOa1rJ0/O
xDvDte0sgVhf1LyaC3bo0OuM0SFkIGugNYd1hmxFX/3knDWH1NpOOtU084lhf7Ksh6VOB+Umj3Yw
2qC2luvpSbhK+7DgLy8vScZ6LoR91oUlGJK2oAFG5UZzCUxOChTfSFfeuowzk4E5B513bNaNx9yL
KAN0RUo8+jVSmf483UgcYGKlsNLc71xSl+2ZqNlY01TWWWUYyKqXHwwfDMKdx6a1Xu2v9pOmnsRg
qxZ7GlFI9191EuuMYePpiwZDGrP7A6qNIJ6Iu+Y/ZDDNFXyNr7z1OWZe7xdDWufgF/fSAh/1b/Jv
3ZoPzGKDVcX+rEQPPl+/BPs/KNmHsLUR3MfmmuHim0erFEFtMdFz5AGqwrDWe3aTQVDd4lxA3lCd
iIiXcaDC561+P1MbT4PhB2w3z+9VTi9ACW/apuQnbLgqOy+vmPXSlxdqApBDjSS4LrLl4O3sgLsr
bVOGeh2tfuKti/Hua18+UZqAF4A4hjak1RaBYLbPNtO4dmSiy9FYfOPGbFR59W1XDJQGbt/7e40x
3VMznSt7W2VPqJYjs/qaF94L+ZVysHTVilAdOgwqVvzVi2EtyNn5QES4pb9aI9eYFA15z9uHKWY2
ZVyPqECs/gavAPMXBtu/zZtGjxAS2lIzmvPi/9FxwOE2jdaHToqosu4uAERgY0/flEaOtIQv6829
5zenv45Zk3mePCUdBXKqiY5LlvLqaMi4WRLHrInWJWrTtaPtr+CCJmVrShG9HXSaWeMmoBCdzgvS
8k6IEilhCrx0FR2ufiPsT8X4YWW8ubEQhVdbwms/k3JN7AVIuh9DuLH4QaCeUJidaNVVUJnFCr7p
4E1iJTEz/+sDnJX90F9B/PpnLJJYDjnop9hF69CckEePyrU6P+oCfxekiqbGnVVICRJcjbzQA/mp
XJXtS8aO4v8YwI/4+xrPryWCtFvpt34Vg0MEHE9jLShht/OjPNUN+BPDjgDT+gOqztWaAv2RFiyU
2htrPU8Naat463D+UXYcM+AttlWgk/AibR6Sr0tX06x9oi5alQYDs0wus0HeQ16DhXiUqgFeThg2
YyrRaI78Ta+fJbRulIqfYYLW8Q6JAMAL4XstPFG44lOfHwyUQZxBlNW73rjtsr2F8PdZXK4n5IwN
BLX76mhYUg9hW0x4gXgFDBfSzI6ACACHtcNJ+AkLtTfy4I/kz9F6D2oo9JaIoo6h2n8+Ae+wmYhg
Tn2v4Dq7jeruPvY0IWm1w/HiPt72XCprNvzlztJo/6Bdlcw8vPtV1JAPyG8dHSU+mgVHPV4IVDsW
ZYuSyEsQP6sE1kyBkl2rj6qcHw1ISwiurSqga0eLevLs6RNwdzV5V/xJSI6bSpjF55FOHJLs9O5Z
thuwSP3Lwgujt5YfsjR68PebSUG1CrpDjoKPXdNmqFpgVE372ciopmx3fRbUyQNJmK6ySL8UPGJM
VE0l9D5vhUwsVLMFx3k7xTZImDXZV16zgkFeYZOJdUNMu/wNECifcr0hsBfKMWmwK9xzClLfVF31
sP0GARFJgrGblTfe2QTIb5BmFlSeE5ReqykyvUoXoF80YUf7Q57O1yyOLinVAsAFQLLeRyIps4Ph
QP/BC7Z+nsFCnMztzaiO4CL6nifRoq3ebHFEZHKgNnokBzNDCb823v8rO3HBxegb/G83jGk8SrZ+
UM84dOZ7UCSWlyhObs4acTMjlLJbgSVcpoG5c/PtgEgYxc4ljHKP/E1HuJ9qAuyEWC3Gf+PVkx4N
4MLH8GvrwGzfGvgTv1ZKQIXD+vBjmHMqf57zEaJ2uTw6DPL2UJzqkjO3CsnmhtfYa6Rt2mCaKqHB
H1LqniEyCweJsJBXOaID/M7oDO6U/gvAEN3WYu4u67YdUmzFHuKo927ts3lJIp+ItP0dlofX9yJl
rHzSsa7nR0viF1JsovGFPK9vZO+jpjWyz2co9q8dJy4QgB8TNo8myMpnDizgWK6z2fjoqNu5Ku/e
5bMqv2X5HxADLgq7sU5ZWZ+K4cl993mEzCRRrBdjzEUfDpraoplokYcy5Vt2ssgBxCHs/m+4WPeT
wiwbGDuAdRKcFy6h09V74wQ/S7w8etNqT9Z/0dE5VVHiOdTCxVt+GySgvtoY2vCuZ6+MG5EPLByR
a8CD2j+JcnI1Ua5PfZqQhHfV49V/ECi7Kt5ufmX0NKLu53NZhlP2lCKqNw8e0I087wtoXYQX/gzI
C65uquboJpL8P7refHp02QPL46DI/DhpwjUGuPAYfxPHh9CLJFg3aiXjeU0p24cIh9o0zbcpMguu
KnAK5jwScVQht4kdvemoUJGc26Pbo+ph+DBJ9zRrJ9tpTjwlTJAFGwqnx/Eyz25EZZfGwAd/W0t/
0kZkRpXJPp+kKDn35uhFZZg5iUkOtdVSN4GFKdnsvgRZrMgx7aEIkpOhOchGzq3wRevMpkhc8ZJc
4x7c2EmD6Bzvo5S2AKrXIqs7KPphP7KK+AQjBgX/WvzvGlQiC8E1Y4+8vJPHy0pKVFL9HrjaTs1w
sVRZ5sdV6Ztd5UFBkf13btcLvcbJVK4S9YqX/7c5plBiDukHPFlNml2CgJQwNuNkmYYPUm2h7HHn
Ax7vpdLCiLj3RpDEyanfaRA2W+/JS16PDquWqab5CPtIK9gMsllfJ+l+RVu+4yRrJNGvdvtcgKxj
v6eOUaI3hbStDS4b5ERB0zudyyRd5Is430lVfuYGx0x+MOP53VtlTnvyzD4pjAIHdQp5KYUks1L7
jP32VVlT4oWeRpba+lPmMTFOufgHYjjKK67qtbxbjbIEURITYoypDwSedRo/ELHKESu5PW+qworq
RuKO5A9ZW1ZyhoBrYZIwg9LOSdTQurY9sCC9/rg/5RGtDEOo44odXv8P7omDTjaMqmB1T5bZAHop
fjIpPR4o2a5hodth/kumbHvTCzHUNhAS3+NYkm+/fZXdYS7+a03n9+aL4/JIeGBZjKd+iHfEIlrm
yaZ33d3vAMEz3sHxDaXjgJqk6kx/93Nb+wKoXcWpvYBIOb7XKWerKb2OnS2o+2uZ5p0AJJHQq7zc
/qTVSxiN+mgyBgKAKZz4O7gPd+pIM3lDBoshxO5rM7XeDRwX/NwQGNGoMh8wmplPU/o5wO2iVcik
AK7miJuDYeZisIludvVKKHo3nc2qAdVfV+5Er4uNDGpvDQmG98WhUz+2m3/0Gko7uCdfMzAx6Uw8
5DOsSqfEKlSZGEXO7z++ZIv+yp/SGlRrgnRSHHUzhgEHJtQwDqZkNWkWiRRqetipbNLBXkjWqwFP
D8U9yJOVcmHm/jmk2jvD/SBBgWkuxDlzkgifhYKs+fZ2IQyvDNK2dEybgBiveYK+FV3Yjt2ZY3yV
2TjH6k+zIo+c0MBopcxHir4a0uZV7ssFYwRoxwnbFAe6763qPiEOvu1oKQz2oWW4aHoj4CMh9ACJ
FSm9ii4qhxJp6Xdl1122FaNSazqRu9Xko7FwealH6uKHfq47hkTVvBt+tDqa+hnDGMxD5QmFRlPr
AZLq1pRN9sCNIgEsuycxeor4k+tdMhdPA9hrozE4xOZAelYDOR6ylNRnNuCYChOIBuDmD4P6Y77T
Hrb6M7XDpv3x+yhuv/2+B+6xora1FPOLQqOol3tbAQcrDS1tTw2zUcyta0fqA/gF85+6WjeXVzOe
qosDQxQLNgEqyp4DZF6m+atRDKcrIVPtUGlWMAjrCkb2a22fwCi1Sz6GHGdBEMm7/5h5fNTjoSwr
R1SShiKGKbgOZo9DKZAkMQJA1fi/RHkF6Um8jelMlgcMVs2ZjFCcLtClMIDntlAEjMoLUFg/75hm
fd9qmP0LuWjaGBTyHFoTPvD/iECSTK9pXgpj0MNWTgd32YRW+LrzYGhL1kYmEPOLpaVGrhH1UJbk
o0KypgyxpR0s+u6MDogMPifRFS9s4P3lpVusttGLPRn0ACx3m0Kd4eldGcXdJYq9uT07usm4cFet
kwcj2Tv55LWrc1SnIacp+aF6ZQanCnIkcfRadrSCI8/Qw5PwFfSllj7Xctgb5+bZYOejIERFkkgd
c5ERSW7mhHbX0TSR0AF21dtuibt+8Mmjxcn7Lzsxczpgn3qLOfDCpFZ3PMdFiHhV8bwznlj650KR
9ldTZVvIvZ2C9Y2qc8soi+adw+1OiNz6ZiiWZ0GEsJpOO5Gg2jv9gTcnJi1lM2lT510bsxNHWynB
t/MWAo1EbT/M2msaMZvChFnEbPx7lPGRFxPTqAt6F3QHkRuU4OFgdmNq61VVwueTtI9zZ+QFQM41
hc1Ah5+c6OWeyho2+zNDltaK+qkIBTuLXqh/wfMdvGnSO6knYqiJRUAv2quriBW3NLUBbMytJqr5
3dijSm+5xQpi3r2LhJIgX+MtrbAkOJVvVGZPdvibh/RG3WDV5apNOtRPHuhjILO3JEAKGiyvCOhJ
xkI4K7KyLz9Vn0f6jj+Yf3iNDNwt9HhG36RliQCqabC+CqtrvvLHkwpM3wExYYNcdM09If/Mq1fG
pBuDIK4hOtqFlJa2felr9AdEwM05+fRfc0d8UsjQvQ63jO/fG0b79sBuItb4Ko+D4rBN/mFC97UO
5JSn2QPuHqsuNnSW6reax5SRAUjvLWpRAdYu3U5++dQsosIDIZmXUhS0ML5DGFMq2wtWW6W27f2y
yjBKUS8aMmXLoCqM6o1edv3X5jylvZ+cFH79B6t9bArXHfQOum6WtLyrG62ScRXzalJ6gyVnnKN+
9P4wb8BOD0dwMaQm4DX8gh0okj2RoBD9sM3XUS5l606VJXrxeGjXbBrTi/JJYvupCaGt/fd0hAvn
wUnmczi97tqHvovfZFW6opfP7NUS3QYE0jWDoS3HUviSHTiuy93qzMCgiP3u9zeEQv5iBohR+2/c
4G+948Q3KCjqZLVWkA9DZoddmcdPKQ6dEh/Qf+DvIODY9nCFqzdDIybVi9xAGDOl44yIZN94VWYw
puG3JDbJR+qpCxcsp6U+PWR2B5vwC6+sO2+QsSYu4PXKZ9WG3SD4xky7U6huBZV5NZ9dRQJG946k
2fjHQ6vXvd04qgn2f4PUvIDpIZ6V0POh2bst6eb0RI2gPNF2rIbtxrjSKSRKL0z+CbDYczBUrFGz
GIuEHdrvcVu+jtrDtBg8yGrpeYlI9UBKJOx8GA/WNZEnQRKVQiwz5LkamlbwJTL6rTblNZEAdhcD
XtowBM5acOHO+lTnVBUcTjurRZLcXTHVqdTjm8mDKmYeCtzw60UBbg942+lksa0uBnc1/t1qhJlC
uf00Fpkyum9EBM96zBEz+zue8eXDlwsYjjCz1NvjZsLc/FIRT91eErhHgp9rb3YrUfv9x461QMOK
mFGH8ds4/e2K6F06GZIOmMA/T8LpgyePMA6gULvZr0nPPqiWvZegHeQlHIqVP+WsgmTfZV3U/wpX
oOqHs7RdD2BLGWEvssFSHLxaxuLip34v/ZUnQYku4K2hbn3IZubzMnAhDoCWnV6fWaoMyLr8aZqP
OKzN/Hnfpm0WRx2anOCGsGBR2weKozW5wgtJe3A8M82s/2WqMbKPb6MsX8MKUy2lz8QJSdXFeTvx
076W5m/tD+f+3W28P15KUxcvHVcdAkodOGUpFOxV6IV0be+ZEBeK9Ma2HZXky/q4BMWR4o8ZjN5N
2bbts0zYiUy8B2whXxIxH4TGKcnG4vQvOLo6urdGd60E0N2ikYjNzGxFsVLYr9Q0R4qFV390LVGO
ZnEYe83uTAqBmKuREydWqpgJ3oRZBCqaJkF7++3NcixgaWZR+aB/QWqr12OKdcm6Dhs2zkUG7P40
MxsbCPPj44OwUXynJvpZ2WWDWCi8asWcUUa5GSnvbqShAuDwtRQVpTLAtXoy0x/1rQI8JCRN5fhL
N2jukS+OB2MhSVLu8LzUo02Z0THbZME9KFgIgNOfJxj2GXprtvC7noT7Sb2VVNJy9D8/6g66reXw
CkDfFO9vt0xBWy8MJ+X2cPYGz7lDIhVS9OFVAekBl+E2EvL4nYMjXFqUQNiZ2sqx8Yb/C4ANBZIh
FTAKS7k086JfCpGgKLRenDwLZnh38iqsFQiZtfpFcEZOPjE5mdTtSJLEajhSk/yqM7t6fX+BS5m1
QoqF5XRAMhi7w4KzW/o2WMYEwc6c19lcD8ry5lFjPq1iz6y2Q1uhNMbpZxcS5nCLaIfpLMlKsgyt
VzrCYFLp7JXOr9MKn/1sUo3YZ9mwTozEwXN0ddf9Nw//r7AKzrZWB8+dDWkePbIBgOm2TNRIOxpF
7M5OTIi3b0nN1NvDFmM3LBYa/5yEN+/V0+A+tsCukoGIeZ/bm7pVIepG/JDvrFdCVmWtIrXqIgC6
KRJ2QjyJ+LpzdfupvvqHXQSA7xIraqcFHIT4sSVqTFtv1LgfrlTDvZ++/zclrr5w0zBmqgw8W7cO
pN4nPtvXUKKzoaPAtTckVsOeOUumieeGU38WVkcbjseuZZSkGeC+j6wmwtg+ROJBDGkmZslGeko2
p98nJBiNFb8kGhqf8Il6U3DBB7rcG8vYWHZlZPflG/iA8++dYmX6b0Y07pmpFM+OqBTFEEvEQRdE
PvelePDYhWf6sQbseMMuEwfmlEVvrVYSuBas3FJYAh/39zZxI9j2kzUivV78a07WS0jdXi8HgTSj
Dfr+uYgP0uRyP31Rk59rEOBuOvXJLt/aruMmHBd+ZpWhW7OgBDdYN0ewUZdAiCVm1AczDRYZJgpw
FLNOYeRou8A37fzbirwS4DT3+ouQnvSOV4wBOMVnamFrWOj8LIUiW1BKoI32ZZocLrJ4+DSax80C
kGMerJpTFsqheLLZ1Wuf33duukUlLfthx3t+WA+AH+cY5SPJRLdCJw0HgLjrfV1wYomQ8PurY7zD
xYdqqUhnNWIMlXP/UIwmIE1k5yxg9LULSv2fxXEpNToN5jGe3kEkZyZx3RAfZNy9xFs0nyU8ovAy
wBRmcBc4PnHGrq49agHmUE9me+iPxpVXuSHcSZYB9iwOv5HLzSWNJziGcvv6OwFV1c0Fi+k95weD
wu5IRHAgbheERoeXobBTrdvsJTsG3zB6TA8IDS3eQjbcKmH3/M10ayIW49KSKdW9ddKoQ8szi2NS
FZZJiFghAAnjt4ryC9BFY8DTX4OoenER23iLTIyCAPt2TrY9gVR6zCKDgQ0areXrDysV3vn7N0g6
MWx99sgb7BDjoWDsILIeRWtbBdgpuFP4QPAoxNv34Rw5/tajUx/Zud1WLT98Mbuwqx9iVv1M7h32
feUMdxqcvdkgtAH7UIIR8ouSwpohzMiZj0j2Mgyp+0hKfL0PfOzpdQqVMf5+nmW1spC1WHP1nOIW
sgjgh2vfjvkWZ9JXs0h8C3DBOqYZET4fP6cIwKXeLgd9lxJ0wsZYeQCe6oumxfISG11YKTMl04WK
lpZy+QBN8PBmedylznPvg2F6Q6Vxf9zw3H2NqCLiasI3b7e4A2CXxmgh3K4KO5R1SexaSNHwsqhj
TXHv30geV/dYaM8kG+qha8dw6PlcsY9p5xaUA51om59/zEFScUokFdH+2Kj1TwbRSEEoBvyFWHer
bl8tZnpb0g+IBYbrR26Pi//drtXJqwrI/+y1xthCjHqPkLzoiFMY7WSConuPTeq7Fxon0ljkRL/6
O5goyZwEMM9De8cypiywa5irtfGIF6M0r8nBvAQ9LrhZPeqLd0hLpnC5DVBXPu2W8C6Cp5jE4Gdm
2N4xvRFTXxjr7hiRJTpkWjSEiyEkjXfk5PXvWenkgJtjzgovBU7xvEWKzk3VbDb5430vWfLTI/KE
fMKne4ax6YGPvpv98bcoCPQOX4ar4Nwlf3fXPlPYOej7A7aNsw06K4jmeORtFXsFw6+SD3dSorkU
N8EEdPg4shN4d3MxvYrfRR7mCFfYUTXWtg1T3K3RfQPi93x9OP+1ePP+R7xeLIHEgl8wlSz8SBZi
iOSAlR0+uYiH0rf8LfKvathnv8Ik7TEznGOPEgiiDYp9Yzyns/7+0iVO5PbN9EpekCDuFZ/8vGp6
VOxW6VSEUzTl0+woB4Q8CVA3AR83RylM3DxIKldkBRVHO/Fox79aCbK7Fuh9046gRG1qECRqbRNE
H/678Dfc39hkjGxJjr0WVefLYgazqa6x24cSOJlz1oMFftgSKtjtdcPsHNHTVbaS1Wd41wHwXIhL
9LaK7M32hVXblVOkSlfYP2tOcwHyA1+v7O3a0o/ddKB0XIgsKF83UNgFe0ypJbA15z16S9prGkuG
1MixDfHu8Yj3FLVHCASH8Q9gSqF2j4E1h7M0X3A1mvlFj4n+5QvO2/pbirQAmoLaGfizWFKlEiBY
AquYVBcVSTmas0llx/qiM0z/5sWt5q4XKS5GiFNV4lo6KOsVpiFqX+qN9torNdcxy0nBjNxg1ulB
emfZFeokGVIVKjb3JngqwYVQd93/FAYII3J/gMw/F8ElHJdGaMPsDFLrPRWMZ0ylWJ1rfTVMFFh0
Y4Oq3Ku8ZPmNPkBHa9eC7QtYGRj8ZAKJxXwgUyaTIzZ2sApxROrHLP7yOlE7elZxkG3/he0zMJPT
WLc6iaj8KTJACGRAg1pkVmMwdyDlJkHWkLtJM4j0fvepT3SGlBoDETt6Rq9F9m7DYY0vUp22i2Ay
YQob/GfnFM/Ku+pagNhSaNAwT2EqzOlHtEmEj/kTAnMOOdVWh7E9cA/A2neT1xM4EMcUjpqaYxL9
jAxo1pTh2DfzUrW6lsXQFzdXkvluqeVbbs2MpHiBadOXTsGsFTuQAc6a8KDFcdyLwTC6Cku7mN9G
xo5wMrChnhCFsEwb9Zt7QOj88AevdLRV84fi6r4VIsBcyqqCHQw2TU6nDff0a4h1VIxRq4ebz5JJ
/ULaTo3weewFg/oJLldqm5GRqvjxh7ob5d2zJmA9KmX0IACYNawVyTDrQ7Fj8tVbj7HS9dfS/ZB0
SWYCFoqPcrkj1EsP9+q4CPruJIknSlp5jiq18B8f0xtjzjmwqxhsJN/FJDIj4puuXtPqToKX523R
sxA9Us8j5YmactVfzRf25H11S7rjfATNyg4Z0CawHhHA3dj0iRO/cUum9XW4Vx3LRtAfk9vEjdiZ
HYcQ+WiPsPP8U9HHDoFfIvp45jqNSGhJjMhPqYtSzcqVgPTioLhweN0nqVN0+juvxR5J6uDR1WD0
xJPGdPiy5Yr03nGziYSwzQFlUjeX+mOjiMtDvsGgvNMFWhnIRCP+oTkQopxirUmKJqKCRVNLdpy1
A1Gvq9mnTxS2JnZ4sRzbX9m4ZvkfThhTZoaRXJbPpUAPOIWaCze/jVb1PB22gmV72igYxEK1bWc/
60DQdx83lJNFbufjJmmDNJ7VKnVVRBXY+lG/Od88QUFo9swPsSuTeohAOIlg7kiobWBreD7+2WSr
XN8Iah6U++d9O//PIW2rerEpnxW1wWgu4K44sDX7pThASSvhB9VXqhABTPenrYtLiTWqbb/pwh80
g+UQftQ9ciGu1ga3f58tHu5OxW4zS+UffvWttbJQM3V6LwPxv50coCLOYYU6cPMQSlOOvkBjaNIP
8y66iAlT7/9Q9MNFwcT5WANdEDwpD+tqZph36EGCYgLoHfaALeNn7uSemRHzVbMgIn4EAY3TR6fP
GvnM9LezvNXzgEUXR3bJpMfcpD4026b4LFiomeYbD2Rxx3S9+hceO1eSaPYQQ49iRE6H0fC8a62K
XWbTRQHjT0KrMr7pR8aAIifTl6DtA3U0QMd+r2goGATNS6xaxWix5/5Q3LGgDflu+RmFaTyfBhvL
ENGwn6oJZt0t2uO41C6OnNVqS9c0P5lIASVSPcK4ng/kTNfwa6I6UA27JFvscf/ZpszotO1raMFC
IbFv5qfCgFe8wrGLOKdawGohaFw0/VJkbCXb0YCERHzyR8aDr7MX0+4v48q1/zTK+4rSA/wrLaWa
x2s2oGntoDy1w2s05zc1KDi+yP41aGVW56fdx1ctd21dZQ7fts55GKI/8YS0nupTHUvVrizijbVQ
LXCpUV0PBbexGFhs2o46guQE0+F0JQGnTDn/RsUsFppSxUf/RjQi00bSt5azUhZIM0lztEhDFYCf
sJtaLQsnrKpxDjzKfPaBejA9dnVeDeC2n2YyvqCaOhdtcJdJcvH8bVgqDSpHCxGoQQzjgWyGfomV
gj6ikRa5jttcJyqbkU8/xuCOIil5nhmjroOsBb6rbOvNdbfsQ1Vxj5Zu6g3sfNs5r6isVt4XmCT6
ZK20gVxRxkpvJuqIqRBiEd5bQonZ4FTadAlfpVgUhFAamGIoMBx7XfnpVhDArspbGAu/Ok+IoyRA
j+P+PNuprbEtP0HOQqhw0Jhyo+SVqNw2RaJ8/TL9ZoKZTUGgadwRtvRMwv/HOlguLUAKeILYOxA7
wXYwOFHcNjCUXJQC6o22S5uN2WbwT6EGNAg+0kNj9Ne/BWoPe5Z+Yc0bxR0o+Rrtez2CsNxgGefa
xIwsYzlervLdNP94nl8HenG+p/CiBXX3nsRzoQTFrn50+hMAlMvaGjRZxd7tzfj9Ai5Qf3t1glPA
xvWFhW/urhVVithjbjWswtOHjz60/Y1NGvVBRJ/v6ARurpsn95khxYVETUYz0UCHUiq8jqlcNY3H
k3hV8WGiP5HXi5i4TD/s+vQjebEKzLOaHmWvovoAwKVBx88vB6JqoX/iWDLoGUpaZ8OLbttctyRF
Z8A/4q4qgOrUzuz9NYaBLeQX8uEiuhc9aph9MUwDFm1kjDZvronUImKbaYTkeRTgOEOKbbGWCp3z
SVW6zWBdQQpr8ML5OKm1WjXzHO257rt3/SJN9shQiB0LLZdPIvRp0y/mrCcfKijyYVZOOGnhyIom
WjHTh91dEYlUPtCXmDFwoof6rssm2n5JwwkW8KvFQXJ49tC1qkpBLuf1dscPxj+P3dHF1h45/R2L
Df/hinjCCrADsPi/lj8OzPjGrEsyPuRThNnCEW4x/1i3s31ha3xDFHsj9q4LEHBf4vCL50I38BmG
yN1UyNLunp7Vy9E8h3JuUeoAQa54ZRwTYdsQ50qfZ0Dh6k01ujtheaveSbkVeIvIG6R6rrMqZ3o+
+pqbGo4/Kp9HHV6ujNf9+BE6PM34o6OuNAn5JPVoASovcMO7+sOQeGEf+KBsUc5jBObM2742CvP9
sHepYwLWEgVTYXaTVuJeBm/0M/jKMscokWtH3R8C/tfLkb8Wm/taXSSXlqpCZCYJZGPRcxLWAYNc
EJt86mRFRpv59x0defhnQDCfGkixR+G67QbADRGg1Lao3ExurfFdO9KPUjHM1oZMmOT5Rc3RlvbC
b1E5xfkPUFqUwjVsWExEFXDdZ34ow7rJYF0P8Nwrihlewin7BCSJrOrDCwNAqNnUk3r4GJXeQb0e
rewA7dMmt1I7z6lpXR+a0f7/VjG+9w6gZGgLxYkXSc0mvW7OegpYGbqT/JuryP8TlmHcTwj0uT2Y
WKafKc1SoIWj2VkFffd3qQz11lv63CukjY6apztZwVOhzagvVkM9gfdtuHvV6C9uA9TX9NRVr8VV
cNK0DBsXUYLzvKUjTFeo04N0ueZSOTpfyE29GNG4QdSCCNYBN7A5F3DF7iN6Pid1LmYBmhsLNxto
/+2KVcsjlH/u74jAtmkPSkvZTGchOkVd0xZhIYJDXJoTRxcmKKERxSssHutYcYA0WP5EE2F8yqtL
rZu0R/Y5pNw7kGkHugVxgvL+GUoagswG++zIg2I4Sy8i/crBCumt8ki5i6npuU/u7Xg4ZfNd/ncA
ir3eKnCYgakl1eyI0G1SY7bjY9uMP4CahyhlgmYrmtkIjMX458EeaJ9Wh71fYevDnnq+7BwDKfzX
A7/Jm9kH1XAOfpn/ErTGUurATlEjUCBGPVvFZiQb8zUBtqqE12u80grupKPXtvJ9VFeHVKiRex+b
YZwXjHyerubiig2u1tp3uzhoUWXz0QPj46AuBw2pL0y4HBkuIfon2n2wcwkJCh1kqUIPqjkz9lBR
rmr+yGOetLLw2uRne0+7/sJF+DOuFr4kv/F9t0CJKdK8QeZ1AN+EMlQ3NHLvfH3QREA+ng1fyYjq
Zfrizopb34bZfDz8fuAvgG8SqyuA7VStkLKxWMOdeba/9Me0LDPtvX6tci/M93Q9vfrA3qL4fbC/
gUdx9zNuA2SbELH0JglPejnP6tJCoxzjC+xPHFp+1G9AKMNr70iU6TxhlYbQ7gJOkE+crh5p6bAo
kaTLc2LLEoYHp/LtAubFXpprRDPs6ASaVN2JeolG5Wfp/9ooQIA+oXIkuqpY3MdQWB1RVtL+0ZLL
bm/0WKkZrk3FhJt6OroFqVDAEn9hafPAQvhx8AWjctCUzw+cgfQWgTkuagH2ppYqj9J4G9M1fegC
ZpIlC0Yt//KXAqwC4m5BH+3rWinHDcO5pazVefHr2jpY1tAt4U5G8CO20YwQVuLrUquOgYr4ZuHU
Ep/WeuVI64vgLo9lkTZNZRBua6GIi8T56XxSCUFW9kWjFTPPHPJP3E1npH7oJdEynLoGyJvV2H7T
/Zpf/06fn+eVytIBxpRmNOwZ5/6zLgzgvHtUyYMeNwbteIuutYyqG5YSoA6jJxCODen3u0rCP43T
fuivtfsGn8HA1htZhBcf5OftpNyR0wDjlHEjz6I4m/afOAL3tUOGgoK9ib5CBceWV7WNcFC/BZiV
5SnImQar8Ozm39tvMHwFvgthqK7A8jjyFt4+ryDMRcHYC7b7u3nLm+jWMVjaelDYomvE0eekseka
c89KUZWd/QQaWaR6T/5t6sjb/iB5L1izBaS2zGUdBaGaCJWyKRSoFyNJZAgkhosCNavgV3TMrzou
zmdunyff7320CxTqsPgYT/jlpi+S7WDz3Uye/5opdI09CG9GPmjTj/D2PPT5qU08rRlmXgBUFiXc
XpRuYWKqW2hY5laJia0yfzi01jPDp83t288DVyb+gG8lUvXzVjaaomItUhuIymwYEMD6t4ypJ+62
CnncqzBdlzVxWQZxEgD+jrpbkOVL+ce7sFC9C5waudmoo8ZSlSVDU/tq05zTqJip83eWkV/+X0XL
nnomuLFeSkEyU22CetCJD7iBi3CpFpJ4JK5rIUTsbjsoJlTweTn5tbBATn8wZAwv6Oa4J6RUAQbN
Fy39oL4lLemvs8McVbRiPiZe+uffNLnmxFkqzpys3N+yym0CdO2eRpPz4yR0K5AH8a3/Gi/2r93b
y55Ehv3m6QWCm/+KwtvAO1t+EXE9K1TDZXPrZBeoHZjDL6NBSmwj7ir/xA2ZEQRU7kDiphx3X4+m
wjOZQk3YpcjpYJP9R/VtiQ1kgFGKEwatM8ky09HYZGHnVGzQZGJhD6rR8dgI5ShoxxUECjKG9Zdn
CPoBvsEA6J14RWSBXt40vWrt3XictkeUMwJEqdfnEHiu9YJWC5Z8oKBG/wO9ILnc7MAWvW+uWDnq
DhtTg73uXJhj4+9m0P1rD/Fr5ykZcV+kVQa06Iwh+1quG31NKO6L5wxBIyTtweDviNFrvzk++ERA
JKsvpajYj0u8Hqa8VBAF4za0Uvc0Zoc0RjJVlwWa50rbiZB655ucppabpOZkD+W6gP2fMgXC/m/p
DbeRe6r0lA9rPIqsTyzqRdvwe5w0MpU+ZoGimxjYQuXwT2QFuAfHswZBanmUrLzbHKboAmJs2mIJ
PHHJ1V/Bob4cVQiNt9P1cUCE5f+50nZwzglwR+ZQ52YFdl5quJ2LBoKfe7rHKDoPlVAGZfQSAnSL
Re4Z8eDfcZLbpdzlKk4BB1W8Ni6JgRARf/FnjAI3NHQHWXaxVXCwkJm6lb8LdxxAWMIEi/QXAlhU
pjItrWSO3UUDTN4ESaFlyFh/sh74G+o/FPUAEI+Gk4yFsfrCC+Iwg3kfRoC3AoX6zW9irDqtiPr1
OcMDFPR5ThChrRjJqvBIM4WzWJgE2QoJkJhK9FklY3vjEotQXyvgMNOzHqYe3cITAX6spNBmNkBB
jDAMQ87dws0cS3dVKQuBXcQFqXm4sQK/fMODRlEgbBCct/VDDtkrxedsG3y7nH8QDjdxYwhuX3nw
bEIyt8ecCCguvSgx4OjzIWLI4tGRRCYJI9GApNnOH9YYtiIbpDAYe3UVRqkQtxnfWLvihsk37b5X
N5kstczE+TEEkxO1YLWKH93lvJCsnlmBopbMSxMmpZ6UlIwicZ5deHF1aGiGK5vp74mY/WZE6E9A
XmIn3H4ywMhlrNg9boU7XiXZ1fHQr9p3rSrjKGTbw922AQsHHb4m8ajbRAhTUBigidXpLc7AeW5M
QmYli86hdVUH5ivPjYCvT2lK9J4XiDp4jdpu6px1znJ7k1GMl8ksESJvutXsuZXwm6GlYIgK0n22
pbVn9K6UNgPCH/iJMrpvfgLw83DWT2zoDFH99gWcc2Hr1bvrjbxMcaP3uFvWNmjt1HbPkVE0dIxb
DGfoPgm6tVokZ0zWgaeVyeEYSL3Yf9KuExtPZ10pJgIqKk3NFcVk48KrKELLBBTn/CHYZuC4gXYZ
cBn37QJFiaJ4vxBxk5QSjMgqJYb/qbUepdRDBJkDhNOY4eVwj2bmAAGHxIs3A7XhACsOmGOFJnFD
z0y8xAk0x6Rbb+H7OBGgaKexPenPJk4IirGoBAEJ2xblhCGDS6LLeGSdtQFmZCTj0SHvsz3iPK+T
lBOM+RpeFBKglye79AQ+cnykhYIwiy3f+Og3prxF+ukItXTjB4vHGKxvHkNcZHHRCn7d7GF1Lrlw
1aew2j89PIl3bfz8Rz6RChncjS/zImJNlIly2//bnlS1YWAXBfhWuhXJeqdrP4eh8W75F6OH/okc
g8/BQ2Ew8XgD4MUdeaqfXb44X0exnm1rAf1WL+6ybiKNffYrygWcu9XFfBfToa4aNz8mEtomMSUQ
rG+Toi/ycB+zOU1FW9qDycCLJVcs/FYissT9u1+lvvL0DqV3dlgc1XK2VRb4JUil02bBf50qzYHO
xrRCYUaGwr95MniNfvcAppo1r+J3M/7nCjebvRA3PxYE/yCQZ7bNqkpGtd2jHr6rVuNeklWjPMaU
jSwRwn+qIF6YOn2sAIW7joJ15EJVegy+5TIRHO9a9hYQpPjCndfudxtKYVlMCvVWRcK5j4vUjMs1
0fj24LnvAvdyFF2BU21OTX8SFWh3BPlDSdfs1E904y7eTmQ2Bijy7JJHwHZNKhLfWu118+Ijwz1+
Z8vMyNc0mKsX5C+W5MLf8j1ojQ3Za8VVROJJEMbTh0RU9hsYO77NM1R2oFy2v1E+K+UcZSXmekCj
jzMF7sqq4nly7ALodW3PPuK+p1bH7Re+l6xR5stCcR5LkyAe9O6+pxl73WDWKXNXSlyZwysNh2QO
jUXQLgmpaGAYX+0SFDGXjTMVI52xY3bw7dM1BczvKTlpDfOQ/M7/tRVQFmTuCUJTBiMW69Y+lbXL
4q+oCnd/pRYSBJ4m0cLd0iNdjJNFUmGJeMYz59sEPXUk4RBkMkxBofM4BCBYfX7Yh9bZ590TNsc6
mwpZVN8lLzA6wdz4Wp4N4o/oMLQ2KG5BnEz5Wm77yVHNwTLLADTnLHh7Yg50CqLd36FZlTCTskEL
Ve0CcXNNYxhxTjP6rpnxSS4IZaYr0cE0vwWfOaKqdqCO0DVwxHENbSuXtv3IzKWUzxs8ivYRZC8u
t5MsTNuNUKI23kCvvjqEo88B0FCxEjw33EfRWqp5B8/ULI3hVzOyfOF+/vVNO25MnzEdiCsy94tA
4R+iI3V7VRF64xtLMHm93f+H7vChgfzYxaYj9GxMsFFXD1Tjp/7zTdDEz9kHeeVMo3WiKsw4Do17
EobP6cnYDZtmxliz/sICTGy4bSBs+3sm0j1mPZJp2wjtPCeYa4a09CxbvRC7R6KY3QbhlFlL2pZU
Mf204Oe3+NNc+OlwPoov41enxDzqGUDDzjv8S/xXwreEoBQIXIxnaYLtZOVC9DRzP5peraTFu8ob
f3Y/wIy5Sj+FhJtqzHPx39cTd4hN4EraTicBKDfTb09lo5XKMtnaWvGxMx0KAyCLuIUGXhUD5lvA
tjKQDly43G9JT+8gMc6FjoQNE2S/f2xNLiK3Ko8FICUEqMqRwKjBzZd+61hAjUaFX5ezsCTDuUJf
9d5OUvKb7AgJWO/TcktVYSFPvU4bCWldMY+cJ/+M64hLriVvv7+RvnwwvWx1SBGQgBHH2HlcGt6d
6vyPHxIMFneQ4S/1ddIvwHUAgwOCmj2fHMTEvGSZa94LhLOvZZsvIdUForOCQF3uD7EvdVKgFOk7
SuSkORihOndn8pPB5MAHsnTm4nhJoLCVj6RAfmS6MRsgCOVIgVoTHYkuTYDEBYrxQ0z5uLvKkRMy
qCQQZxLSLEsdI6Q/jKGVBK1ZrU4MZ0BHk4qmXks+9cVxi1LqBZVhQ8Vo26mXTDrSz4JyhHZ1CSaM
egJ0N5CxOwQlvoQO0OsV0dC5l1ESP+8Zv7yYv3oIomKFLcsvCQz4L9aJ3JguyeoY7pO9+UDA2Fwy
uPuWojMWxjoDv+6YjOI3cP6fuLCCWIIx0fo10ApGC4gsZ1t2U0Ptlj0VQl9ASIgjxdxU96T7n8OV
S81W6Ny9K7y4QSRpN8yH/jpBAAf8kbReOP5Dffmcfw9Jjrw8pFG6WXcTxjjLEPDc451BHBol7wJT
r/UQKXfX9zXTVVGia3zjJh3u1UjGvCSbhOwPUGuoUaJ8SX/CcjKf0h7vBSdKesO6FJScjJd1/n3E
CDeDGI782yTKHLw3/e4R3niQ8GlAYzQSK9j/kwhDQr/FVhm9jb66ZWQmV2xyHH+2hhelNwEEjvWG
ietIMbYCgJ71v9P5clE1FuQh6o/ZXwCu51tJ3k6MyLd1F11DFU0G8AQfPbUaWMdupS55PRO1N2jg
wpkv3guzLFcr49vsOcUpq9aVHYyO/oEsFfzu/CRKH0fU5u/vyhJhdRmlyvlDW72oe2vIdZ9WdjuJ
wPIYv18UK8WjbM3OXHIbU5nWrDTzX2S8nImu84i28k2F4xSqa7muuXRJK1FwVRSJ2nmQ4qiLmuev
sSvT4/dJVUj9oKahNqBiLR6tBWHZwNWXuCIk0p6plW/X3jXtynsn3MQxYlqFFmqg1jM4dxeHOtWo
h6H3wXnGT103VLna8ZnycUDBEDQ2JeXT7wveZf1i9HiYrEbQ+gzVXHkhjth9Nw7mVrMImfBlcKjP
1s82SW9Ir1HoY+KBh7uICxYvQcGYXcxXC8P0Jo0IAaEw774FswmadUp4C5blEqKR3sPZkkk2Zs9z
bV5XPgFkAPuD4SFCrqlwRFCPzWtwdUcSxet2NNf3YgqHnQlUpwemWIyNg6++DEfFnSI2j4eoexLm
PC9oGsQGOk0IuKGu5PK9dEeOPdyn35P9ccYltivj4Agkw4AKv/+2HJvikL/fPYoFuKn+oHIiji9P
UHoy1mTBQ2vTdegcwXOtqi+YRLNQ6gmmrSA9rpS8WBrmCvrADju4tUjG1baP11vt9103RWvKm2XZ
VKyH6eXx3aJQdtTuGee5oK6zWzd1tXLRRii0sg4ybAlcFB+/O22e75rxj+oQh//Xkm+WJcsnNXpV
ph7Rwail6ZyfU4RatRu9YceLQRSVZ+LiPB3WiJtwtejf/BeohGtwxYCfW+V4teS90zId7Ql7UE3/
1jYkZAdXrHnto9QrhvO3qPIuFvaU0VD2WDunUBpbecWGeRoGRP65c6PuAHq1jep4S7ezhciZj5No
6O6Z29NARaOkiISeSjdvEgXeo3eFTZsAWbVH1A2zkD/VyJe2T5Cdizr9AXwQBegVOJKMukuzKojG
W3dykwFZAiMoz9AhdM2gFrb7BmQmklXcC0ie613N3y5YRO1hP7qOmKB5xZn5R2Z7iklfw+WdRjl3
+m7hbl8YpVL7qTDPHhDvk1aJmPA3l2Y9IEIkBMPhHpltWcxozpbOJX+85kv+FRhh76v6UXp1QLse
0W3wNmzGulb9OVvNWsUtd3cFAQANxBUHlszeEc5L+X08Uqp3oho0giR0iXRgaUubX52vrkiZ/6dZ
TsbDdh+y1aXEbLyWHB6myjg3po46V4gu+BvqqtGCYvlSX7Sd/gDUh6NCt6E+duYemxMASO94U7m0
vagz+H6VlanFwcqzvZB1wCFyWjBDXsgXxWmuWzEMkM2YYtp5PNIcYFtK3uMO3TqFJ9JZBTyqXh5I
TXbBOKqD9OiCKaUVUT7JKn9titrHfBMQQJWA0AVsyuQpZoVzw9dJdc1nfJShOOd1Cs4lWAPRWKOJ
WgmafnJhjslMaDnRYNhK4JzJe8yvB6OUERBL+v9/eswj2MjMGgh7x6g50VUFLLwxAtbfmarylMGs
GHdij4XPgsWadtJjxKNytL+nWkVXXXZVK1u35ynOJ3qn8qCVus9lpPnx3lBRb37RyfRQCoNvN3cH
NOWHT3+vOAd2lUvlA1OwuEbvjF8M3KVSz139y2d48bmn06JlDa8IHPdwWeXxjOEkpPCUmejxo6OZ
/noYJLPafBPO6c0JbYG+zy22cM6rndl3uGGsgvDkQDZoDyPjRpHKRwU71ubmONtySSwFG1+nUqBy
3KsHNgtuRRJbL2gdD239ZHr8b2Z6Ta+WFOkCBV3+Z7Nc7MQrVPN9tsTopKEv/HzdKzmUYGdF6++P
iyDpi8XI86AzMXCmwn51I/euUCvp8gYozQnyE0I80yAOJ2B3iBEYGTmbXhqFMIazUwYlaAEeq/QC
oUmt2OSN1b0TKq24qNqB3RhcdDtp0s7AZ8xrh0PtxhK9s3K6ELMvC98UVZANEqDT8PqdnQWWx9cw
rs6v7E8BSDv0d6yc18/8XadEi0Nxe07Em0ZmkM3knAeTapxUqZrJ2V1CI4gBaw9ifv/mP9DLQy6N
UoT7dMew3YUbevEHiKIxodOkzfo/zeCfv8MZtPGKbe8RTaGEtxK/MuCCjgpyK6NWSUKDyKi0EOfY
OpATZTmZtz2Ti5TFlKOxHvgrXsxPze57cCGLUlPc6WMjhGKvjCWdP4BJxxWXUe/gJcjnqmSr3gVR
28hiJ4KJ52+c7tfrGTMLFv8I4E9VtQj9Aub/a8VJzI6+Ge544NT/Oka+CJtRrKEA0cdlyNNZ/eI2
kQ402PZYvw9pK/Xc2yzg63AvVpzC/eZU34rVd0pJA3SLmXqyWrKqnPTgw0J1/2KA2XXV+2IZyBmG
xvnibbHp3Z0YXnnrkGi6DibVLg7UCCP48PHGHsv7h6nBkBHoe4Wkga+vGw6dYktQxkUB6nFQFsA9
6ZNewJv5WRI+H7zNMrCjWh4D1q6O57r+kLEXou9qCw4Dv1/h/beXM/ArtqMlQEw9LcWDSnc9Jg5f
1MEJdJ580be1Xkut7XGFpbPESvrRiCloSNBEXOePkUOIblKjz/y/jr+Qc2ZIwny+iDqNeS5m3Bpv
c+Goueq/1moLQCke2mnl7G0QfB3pNWDzyUZlMEeHG2Fcm28eqhrj0WZ48xzm2E48JTdr7DFnRrZS
Fo2kb+O3NznMIZB7GFtBe7Of+PaLVr6XCTqLKJfEdYtyuVr2eodL+3Y1oI1Rkx//js9hJFQ1URa6
gzyTtbTdeESzHAMf2TjkLBfbv41SKdZNA+nSCskx92uuvYkSYlYFPARALzvw9LD2eS1pyYzazGOU
NLQCIahQAFRfQVZ/uc8awgzWfXKy4r9i19zTHkp/zyWh0pa8Q3YHq1sJ2ym7v27F71cargYhr98/
3ebuvKnxfswKcyu2pYDHRikQPgpeS3Tn4iFK19fSc2my9i9iUB16GgYjrYe9f1mcIZfpd8MqrNf3
xfkWlacmFNfY65U6dRvTI6hw8AxONK0crfYO+O8DMexmfNeAFKqlykfEdL6zPPm50S3snDZ/QFf6
SsoVcSmWxRPxi2LwYUZ5YSoRZhhPi9Q8ilnwB1zBRcyQDVtTUmIvUCYrGsXum6p5oe5SEpuvgLuO
EiAWx/sTwks5fIsJBeMv22TZSfQA/fqncUfxG5k0DuNBUVdoS2M36VgWc21YWcQO9dDpIcqWz87I
dLGl/H1UImfYZ/GHx5vqMK6fbO0qp8oTSfIX+eR8vEYxtNL8VGzw0vI5YwBfP0fiVRbhHgFGqUh8
sU/BqZ3Y3Ec9ysxomizU/v+sMW0JC5LGCRalFZEhjyLqU+Nt25LxDqFan939TxLque0kmMP2XYyQ
dJwcpuZ/cS14uRNwV3TbdEYKenCY3J3n1ILF9IIvF/Xb7wSI9HHk0YqQ0D1nYTHOqTZm3yulOzAq
5WeFqrSlTcuhD/JguUhQx/ZRhm+9OKW3xqkkExJlevGDshlT0ZwHRcCvEChsIDEE5EVoSKMaXdZP
aZwOr2nc3ewVuzh7YhvEqzwh7KuLS7ELwiX8+q5adDc+Aij66VQKe88m05Gs/hDgG5mr85jFtTIi
S3voYOMp5LTwLgFm1ovoA0SMAZv7mNCHOpm4hJhdqTTFEQyZWjVvA21lXGWMVCoKHbkytf3g5Bdi
naIGH21tYcI6YVAUHt9BPSyvaPh1NArw/ZddzKRUML4HdhxbpiYUif0JqNn6ZcqXMKLzBj9R6O9j
fSIxHhj81CXgvBauRjmB2FYrJv/YwPowYiUoNW7bFJxhMinoqS0KASlO0svU3hbBbZldd6RYYsD3
/GubIXaRrrKOyVEDTGDMJmzlXKQzkHMrkr2+hv8NqkWMHF0q5Ts9h1Y4D6fWLv/Sef7Nxrni1P6t
UNAEzXcPWUM8RwDF8+KNVwmdB03Q6ab8RERQI1ZNx8sVUPyJK0Q9vZk9SJdCx5ka8PsN5Ysuhgjp
UsVstsTtDuVvijK/eir4pnzV8iO7xPUM3Oxy9gSNajRIbLdE+6XHTXaj0856jIOZX2ICt10tQMkM
xNDNSaJZzCE3eLglHJsGgAB+pwgAb1cG00P/TeT+Squa1v0OP9eBZ7auhf9rRlHfmpLT8KuyGIPr
aIfGoWPNqPV3zj6ODSow2syUW9TcNcd+N3VeVyA8gOrUWlspK4WSu4hUHuKl/x3mddP4PCcQJ7Mc
JZts+acCBC2apTGT6tW8G48pKQN/E43NInv4ubhd95xT48YkulVahrv5UpKSGfWZxxKZ8b1vHUb7
ccFjgBRi0ynUKe+e4ZPJNRVNVHp85ZeeVYx2FBVZufxKPnQertitKYBYQAgHjWmpfR3qKFEpbDO0
U7ZxJwJiEmJ+hHAiQRebtwnTlHGhLHvH+SU40b48dhOsOsFLp/mLLsnQhr0ub9ZNdD9tS/hZuC9W
Ec9B7jY9oPADfpcf4BYN3g+m0uhJcpG6p+yBaVotTJBauk3aGYbpSVRxH0QYmjGDPip9MRYmJrLT
8NNvsBu+WRIEAPRexV8hKGqKIfgfuimUE/0AmjKLFeXM2BzchVv51//PQyQZXZPhSbyPZw8pWC8z
dxJCn96ven9BPZPnj2H7NJvQGv/Lby84MmsmaSjD/+4fkU75HgqVHaRZ8DuTJ0vbAu9fEPa0CgdC
FZYY8NZGlClq9a2Yw8I1mUme4lFNFlgO6e1F3MsSpsd1B5vYLhK0ryPSe8Fe1/CnQD0qDRssFxg/
kYLXteFs+a2TS4PH+l5oodWW0TEArGpqxVaARIsMP6jA8qvGHKt2U8KMTosTmkde0Al87fXZEMxs
zRTdUcooTe1GDdI4ZVtD3Y5OyaAZftr5uR625jGMBNjQdKk7UQyZaXlikS2bHksgb+u/TglCZYOm
yyHK2MEX3hoFiPUzpyrcyHWTJ/uRg2of477aWg37U9D2omSOc0Ed46gJXB+0bqcVj4YHXFx52wUi
fBKXqS4lr0tjQdWy9jr4Bq5Q7oDCM5S1tfO8PgIQvWr3attLP8JwyVYY9pvpn1evyCgnQlgjbd/I
txkUJax7p3DBHqZh2VqgRkj94EZifK7+RcmvjnVYB6ZRnaEKVeYg9+xO8cOlvZGTk1w7yxN6tFDg
P5/Qx+9HlBPbk7xR/vdhWKPe59PZ7Gyb6txduHN4VsSEtGf77utdFqriWvPMkPhgxQP+iKqClI7f
IoBQJWVj2x9xlOp8jEi1yyNyh5a4brURDfDkbR3O2ql9u7QOKLQxsY8e/0qVwjoeHsbqfKK0htha
AL+hGYnZFU790Q5ZZXalcJWcdD13Qv5URyPsPHHLOi/qFjOKcA9nYMDWy8awsKJ8UfkGWkOkPHFu
DSMwHdZB/pGOp8HwUvcMbPtf6n3sUTvEXivOqrruZXRBmcY0Skr3KIbaFnihQt2TsjbXkrp0vGgm
fVkOAkpZKKZ/W6FMm8sU+2WSsIxf1VQ/25p+61fauUmEx1/CTEqRaq3TAD673CamEWKG7jlYXO+d
VctVnR9GEMJ9iOoZzmkgvLNKFWhKw6Rdrg87ZP8miZwCSc4azeq9Mj1REQXNWiVupgcausHeA0JR
FYgYpJHb5d7Z9WI3HE8bBpEXL5DlUt/5RRax+dOyBrTau05fnDzVjtnKE1Id4IGPoJH3pI5uVR1q
BISQ07X948QO8hRKFT0fW+Plb0kTSA/aJ3GKmTVh8KmaSSoAVyTLILN5kJujJFDD/DMC79Xy4CD6
InZGqj/hfa/pKcovkZULOlZAyyTKIJ1Ng5U1LsYsY3yMnUZtniKH8nIJHfSYT19c7epMwHFCLJWe
XwFZStWWI3Y3xM1AXSWJtAdzYpC+BhBtrh+ESQ6xtR5qjR/N5DVWoJcdUUdzVNxpn9gUxr6qPUMT
4yKI9HEmyGRNy19oqEDle1r/6BBvjIhPmQSXshlcbwiMIr+amfmUvvZJ+ISkVjAIYh8emS5JARlK
8MT/gUIg1ZEnQ5nOMNdOcJq0YLtIp/9Kb+CLwOQyNP9BM+NbBATfbuRRCiQm95qBBAcVQ/x07L2x
5INrBmXeXVRY0BMWBrZKltslnMiulnh6c3EyMrQI21yHyLzTtY+evdA+UROt4FSWN05mbiWW5Z1q
6wdKqxU5tF+5mvWXnIfAGwx8mHqj6/Kt3BBQZSEHmkmRyE9Gi7pL02jExTSYMAUltfIeK0kEn4Tj
YwpuAzJlEovnsxxXwJJ2mSq2edLMtkC2R5vOaS1rxElGpnkaL6I63XuVcmStiMnaTI9ViK+UO712
D8pP5Xv20jbsE1EOIFobetbZwA6F0ozWHN0G7lRhJ03CPCF164GQdhcENTeIXfxKwQ68ueSZNVbm
4aLTMDb9RSge6rfQ/CGAvu9pqOBbZvrG+qN7iFFU0EDbwfCx2R4+kgAu4qjyNbGEaRC31tZMQviy
XXeBb7XB5Pgq0Nkhsbt5pwBoE4JlgEy2e3fOiJohP85RbG99EwsZofCmC+/aQ8IzQ7OhpliX6pyT
y9qsV7L1wVrsg54qz9ijm5FZFJU3lZKXtZCRtceIZmsjg69fM6vpiXR8IcgK9T3o4FXsesvfiew1
j4uD+Q1iRSmyU9CYK58E2xT7JApSKpvXQQLDPkYwx/kVY2rwgb95Htn53CuFcVTE5d20rajcjjUp
650J3XJZm3Sf4YEhhtbzM1D8YWiE3Eo0qi8TQpC2J1BUvrSyft1U9sBc7exx7bz5lBD4MEtiEP9h
KFgpnJJBtZKPMuhxceeAx4jifIfVId+SI8uk5pCrGXZIncP/tlfAyKTPXLs/upim/hy9Adoi7wcn
QSS/DVpdqDYTroUjWpv0UeSSDRTgvbBvHDhgDKtmt4zr63zokoD1vwlvMEqB3vXIpxJbjoGD6v4/
339kKdLsUEIl6z0XLfAJVViW5MtggObJQXEzWd9N7m20G4fPO/l6CuGpnjM5gfdjmlrs3p6JuBq8
JHM6JmXp0yckx/FNJE2X+sv/yOspPovWG5QYY1ooMuPoSYUqbo4pEJOhxVLQyiq42a2Pad9fhr8s
7VHRUw+FOhKODLu4Wv3yNNHzbnwa76xgaCSoCm736fbjdXaYWs46xhgHaawG/AdfNwq0UyeQqjSG
xYvaJMNxTzUlfqBHuK2JT034pbJKm8xX+51eBRpBDv4Vy9Uvqu/WYwEcr5jr3BHTSYuJRYeqNvZ0
Ot51OIf2nWHrcAwXmhmtZTl75WAh2nHgi296JbIBHJXtIak21I3xo+PMZAH5chGElCxVyEcWMY7k
hx/utgyHcLZ55DF26yCaoQWmMFS/x8PlFjfHfh75ttOX9jfGvH/l/j/4eBtHtXrsEKyvu6xAEKj8
DVKI3Q9aWUNRIm/4wtTOMSEFFDUunrbDP904dIoHU7Wky2hXh54Wj4Uo9rRrfYAJOyL2kzsIa2K0
CRP/SEu7L10aXqJNaJrEbQ7pkvqE6HezVbD+rnFBbuBaKrfzKSx5daD0m5ONBSuaJW7jCUKKg7sQ
sr9CmjmASVTXMz76k6lkfuL7Mp2y3XkqNya6PG23sF5hZRx+j29XBjvoKIlvkELGSpJRaWHmqu2l
LlT4TeSFEHRyWUhZBh3knG2eLg3IhD0LMv1RYIhfB+/tRCAAZcQspvkxGceVC/ttAwQcbLzRPpNf
iH7lbIr82QAZTJoMhAVr1X8EXhVNlKVcpppEtvcb2xwpwBbVJtHueR4qFTMXaTvgOAwPqdEcUN9I
mUDu1d+uOFBDRoQ69yJSWjuLu/IeXcA4Z1RCKsyhkds+aqpMyDMY2CF5MS7OFXwa1b62jXfbdrZN
h3yX/l59ZE1IqH/V9m9P4geous1ePlVZkWyggQwgefPuewWmnH4EmXeZ3kPhH28cZtilhvKQuFoP
mengX3Q0UveDQGD73VTa9eMtf8nOHoPdPe7I8emHCk5LNqIsFFBOXhXkHVgyT/z45HHNJEGUrp4E
rpr2wzo3f8H3a+DkoTcanxoQQmTVtMUq12LVmpUrdhrMQ8rfwYElBbUe9ktutuONsKmSsLkbcgiq
27VrXu5ZKns1FztcXJ1WqBL64G1TnDk5aHNN9Q88lX0js5dBGRkbI8Q91lANFXkUdnDOXUC0Wz5W
yrJ2CbY/sWVqyt3CaWfgmGhJq/PUU+bzTyYMWMFNCaefAxzOasWordAocKNHOeNUyKhGLiivax7a
znzV56ykG/7oiU9/nXdpNDBRnyTxtMU2lxgcEAO13hZwUVQ1N3ZBnBv/m/aLB8KjaTfWDpbRNqkK
agylQzi1nHyqsXPuCVTZgAJOFPywRRd6N0CPydcgdLwhqqWDl1GXc7hRo77fOYZpdAdEYmNKS59v
PCBKvEPRuyyXPAnjxOhkqg+SOA6WzbSKOSGqOCgtS9WS3HF5wPIdfYcaMTy4c3DsPRhcYhiB4bXP
oBG5n4e92KlqFvxI175NoAb8ois4wdzkUjzhgIi6F4BGeaPpGukok4gZGoFMhWX3ATkvYB25yEm8
LxZrXChZZNM6VoGFyEusZi3AsYYWjUFHBNVO3uZygzNiiKj96f2EhklM60o6WuzJsbwKi4Dci7O/
vcgnSZyYl+Y7nTnQA2zdvLL2JLJuFfdE7LG5bt2A3LogOGhWEMCgGTPCkm47j93x/7pQdVxsr+um
i9MS7z2s+RH9Xp7E2u6aokJemM4xB9ET3eLkUMfRWyqgkAY2+ZkQQN2tAzYnABjK2UQnlthooM0o
UcZOptnN5ym2fOlRye454jcgcl70NkdKVzgdDb74t9ykhIMFZShrNL6OvzymmDoGltJmPNAwau2p
aUkvn4ufxKh1T8Bygr5/mGgo096fYqYOd6mSw6tGbUQ4F95WF4dvelOEbsgLrnWZ3c2xZbhjdi0s
oxvdRYYshS3FYmHZx0A9jhe2D8d9ERgpB3q6Z4UKfwxecY4ENiqnUqxgVopiAfGBSq0Vb2iiSmOo
b1mDwlSxVpdr4+nTBeTCb6KZrEr7mhgmDir1/kvdZzloXn9Ceu6bRymLpafekpiW4tyWJygRsHb2
bcraTEVVDLgSR2iZ3z8/Lhy7Fe5KE4aWGfs4dGORufyawB5zJ2nzR0e3wiMq+cEBZvj8dNxAcTyY
VaZpT9pxtHa2vYgBoOafBBC9ViAW22ZC4DyA9BRnxWsTzeBcqI9oAGy4VxXLe/mm9txqwhPjeYiw
D8P7y+YMK8ZyJ5R9rgrsGU3UbebG6IvLbxfdNftfLCWtReQ/s+LT28YWgrlM/RR16XQDeoccXBuy
ebHTfPKm6jWxDYDXytwi13s6iTfDKGrN2a8/YPxuIvmDTUUaKxWcMdmOX3P4DTlWYHhtrdH/F7Xr
4V3AurDMv6DzVIZBZrNHa5DL2oH9uh8xAqz2pPRIWjHWEY8vvpHO7drwH4XBvmMsndUogLP+ebjS
b0owo8ilDjp49Xw0KYUojgIN5qvkMN1SfJG7/RFeyGamrap7whmTg9WDOzEs+gTqp1b1zP80F7Al
Y9pNl5hmj4TuqVQlTXKYugYLvbE2bvzm/Tlgp+ZiJCOBMv/McLBLVNRC2s5Cid7Pby7uS1d17vcK
VseQxr5ankXoaF6M5Spgfcs6t0md7HL8SrzZAyYAFNdt0cH+IbNmKbRli71p7mq7hpgE6g8A4Yu5
LXz3Ut2fkt05x60W/eO5AkESuL79cVGRO4nQbw4s7GAmMAuuS2MYxUQRUTuH2b8gv2x2H7kDor/K
kMoG5I5C80m5Hzyd+ssU5MfWN/hYjCyiwel8bx+QJu0mZj/XlqJUaXE8U45luTKVB/DMl4QGIwvD
a807UNVYm5XysJ7hxtFemtzpJLAmjMfnfYTpJEHUjZkGMv3/1/CaXWaZVHVdxNH+RSmK0FPXEpGl
/zF8hVUibAUBy1l9yIbc7hoeXcbWRJkigsSKKUiS/J43UKJ55dS4qfVgTkQQ1wzNbQbeiM1e8soI
934eZ1QYJmy65DF+y3NzL7jdY0CfaPO3JoxP2QpR8D8dL6bHBX3MeS/4tgdG+xhJtCWkI6Df+wQ+
7noPlUvXa+mC05MA8KvR9QGua4c8QNZw6dhw59GwSOOTN/vocfehcZudccobZ+vvP/JDn/lzlZ5T
rfwZNOiLw5vazJaXspOX31rVVAcJWOYiGag/eMcihtnST4EBaaSAgsZWlzvXBc7E+NXXahiEOrz3
b1DOPnzgL3Du3ryOFAMIWskPMmOmW5+no2S7nZSZc70n32sS9RN6KWjzHEwbKodhr3Y/PK6H452U
SiBDqyDeY607OUK7tpGvkjK11TMdMOciqbYmzHFpDwod0Xagv+3ZbZLC8piHZ3+AIMQuBAk9WTi1
U6dA/fCu0z9bCw/AylqP789IUsEdxa4t+UfIOFL48zSlXCBlDO0uLZCxeJrtIiHIHiVMmGAl6kKl
n3stu5Gd7A9iI+8m6a+e55i1xiF83P+6tryV+J6JODRuvDBUHt3b3fkRBT5FM+PAkJxu10m3GaH6
97ti8rqvN3bIukrmRmFBU174+ygVz8qEw6LiGvybYnqruSCFLwRHuA7gqEjZVO2FwMJJayEFSxeY
23AkAd6ThUNoCzxBfhw8oC/9klLRuTVwCWdc1yy5M3/I9aoAkrNR3eYz7tEdFeqM/NCCJtZjWpw/
yd/RxTsJ+cetWjrcig9nw1xABaTdxGcJi08jJuEIS07uLiupHiD124YUD9Fs81265/LcSvnHSiOP
g9XJI9itUWtA2VaeshfA9Xm6pf2D1hcmp79MOoIhk0ZSXt2f9askJUG8gHQX/zmQpziSGzjdhliT
/TgZ3VKuTTWPDUgqAmifWhXI0onu+KxgRLzIIBbT19sSCWQdzZ7NTw/htD9alv38kmpiR1rHYrDs
+RMvVyEo11aYm/Kbr0ozYOhZ009/EWazV5HkSq7gPXDA/zglCSR1cg0KeldY9lU0vW3LRSzXil6/
78zuOBBrq4lA6w1uS789YWGFBbsp/IoVJgL2DAgu3X1ydLZOltgDpvCv/SpyuGkw75pkqtnQXG81
7KyUVLvZ7RoKnajiwRi7XAjEn/ycSLmeasoN0hTz9JESYK7SxI7itJ1rRuM3rJV/FRCD0giMYAOf
OXUkDHLlsKDXGuEIvoCAGrr39mdR1Uj/K450xPyT3nifSLUKjpxaspqKYwvac1PKlTeEjlI47xZh
P1ktPa5oQiQLQ71jqqrTDdPPoLV5IXxhC9+TYrBFDxDpu0ah2rDGkWFh/Udg5qlSV2PlYjqI2Ybi
NdT8zmWMv7EvvO3XeFT8j975WG1S65obHFdU9lLAw7fqeKWh1EJndYMkqQrKmXvwsTfQLfNQftGg
E+p+KvT3NWrtaLHPN7IvM8ol+rdvJVI4cOKfthFOQeY/l895kbieI01vVC0JuDUk/yyszkejPjtn
9kwiu/yi8bFvvKGxMVbkSGY9IjyirtvdaNRjnnFVyJaX/YQc+utHm3RUypPfs/ddfAgFJCA0e6fD
CbAXE+H43UN+OOyH4tVqzPD3GbudeskjUUIBqv+WNSw1xX+DLSkNWVYG7OXDmAHBwoSqQjoHfPt0
KW7FUkLKk4RTgIWw3G1pJMfzSfO8WVCw0uXyqjx4TZCNZOEhrq76NJC/QjcTNVX+9HRCRZn2mzi8
fcUwQYD8LoowHsIxIcCDqsYuMCYyHKHRirrPLlGesUnFv7siS/gETehl1pykZFa7oINfzcCBX9d0
3EJCMyweNOYDSWhAmd9yVonbKUnm0ToplpxKRukkReTFyiCWyt6pCCcu4xzTDQZVB1ED9Rg0/3pv
nsEJdaPDxoM9/xn6UsO20ZmlTqv9NalLQnKZz8y9XgI/7TumLN7fZcBIkdXdPqHWpx1GEDNjaQIw
a/3IbWea4lNtALkUVLFrbfnsnYBiktOFmL9yZuYpjo6qnOZZ0cn4krZtIUGoU9+oAPq1n3dPFXlr
PY0+6odBpt8TY3CU8PAuhmn6C6bZhmfIxtooonnfMoPHB7h5M+IABrtoySqPK1470KXDR/NWJD6d
DBqdzvXrYT+XnMgyBKTXKeqXqu2Gf/YwZVYfA0OIjU5YpMEOUzqqV1s7vzvKZVEhtohmh9ffSGRH
9JpcZA399lsQu0Py0piCyB4zIGtya/bOlZfT89y2+/jyKrfhoXD2JZecwapoYgaWlYUpLFPiRqmT
39exc8qMl0v4Af2J2DoPQMXY+DZyJqMLbYExCdCc0ZLpYS8W1WPmfOTUbtOI/dM0qyqAIsqsxbLc
wAJ42Rk7CmCYPbtutU4qSikjl6O2dhRMP+qY+jnD+25NuW5s7jYkknVUFGUIk0MFHHT4wDQV83YD
bY5fxuXjqK/sq98NaPfFj9a3O1hRDQwKGxsRw9CNJPpnuT0L5lL4H7YTNqeveHCtGpoBSRMgaeGg
I7C4sdWgm9tZfC9BOomYXmkRtjxF6DEaANKrWg+a5caGfNZ1fk/oWLkD++T0qgA72DNl3KRnLZE3
6qmkyLs4RxxpJOcYR3aybQtoDRy3t+3SkpMuI1gENzjp9W/9m2rTvu1Kf/Y2k3o5IAfnwqYAMJsY
cmJVjKIihwUczIeF79vCfMqfpcFP6EYqNZ7y1MpudJfU2QM4k6/C4C1VviYK8vt89WJTldPqdXy9
jxcqm1XORGmvCp1Ps8MYU6ybsgZk8UJ6t/BSAt9Ow8WVcNVtIHpnPCfw+YG8U89tS+vdiD5gyam9
Mb1StkntC+V51nG84IPaplxUojE4VEHpJcC0tObOgTsXgNJALBOQYG7bNpvXa1m6m9B8sHIxbMj3
P84wiseiMKRBvUG4UbJlarQu4X+QqdYe5k0zaoc73Nm/erh0LW2dNGowW6UA0WOEzoQzn3q3j7c8
4qdhLHG3moYT5xhblsxY+qEyJWkN2ScHjRG+iCUEFmn38WyEK35B+ZnRQXzDTYWU4+mpUenAyo83
Tcz+JRuLsH1M2HP36DZIrDQsKmwZjlD8p6h5b7LmCXRrSWTX7S3MSeCLyH/Z5bFXMWuyDF0KZi1W
gxUP/IJ0WvfIwgJyIwY1EfPuj6boV0O214/Stc7/NmkbwceSISfOjWgG5XRE6pFy9sIjxmw6JDBx
Ue7u8qXOhXSHwIwtc4CTGqcqH0qFBGUSS5Y87CrACto0GQerEhtwX6q53Oy2Pt4SEkFZj1eAvV5V
PTfbOEKJxeakmvDKSFuc8TQTyyaVYnO/7as/D4srh3uvhdYKYwVe4ALeC9MCF42g2lXjkdnnmlNA
FlziiUF9hl/HhEXVu6Ytn/B4j3MnsY7n8K/SG4FcVqjHmoFmN/W6Ogajg5WCED6cobL0/fp6wE5F
sDpSKLjSHtvPk0poTlXoYap+oZmnCPHZeo3eadTsTCaYrp546Eu2w5YKDSGlGd7Am7KwxV3X9GEY
pWfZF3TwfHHq0w2u1QfNb/+1EpfYJkodfXkaL1+MCo6haiRfFaNkWfVa0ct89Bdw21Xj6AhIVirp
aHcRl3KPCaFN0wYLwd1czyarYESHIGgymR+iRANCC1PzO304CDkFMFrCAIkyeCebqHdDYb/4ZwP7
PByOB5dBGE/WGGxog7osLS4HODZOaegF2BoF6bpYiJdO9ulIcN6hrlHp/dcDL1EmwZ58lfA3Emg+
8EsJ9AFoBQFHmyhiCK3p5miouW3g8AbRMsJejiTEdQVG2AUweAlP+6MpkGjUmjUJ/7v0ZFceEJdk
J03GZ8rMcWTlyhUaVIUDuUrzyL3ykgX/oQYfKph7DB8yv4xF65Q1yAJPWXJmNTGA+zvUmQ7nrrV2
V3R4Uaad/hilGR9KnC2S8W+GAFe9ZjVgA765CXgSZEASzQYGAKzgKPFaBSoTOK4b9wwFPV1XIJ3Z
1GYarAvBkbXQ5aq67emHCbwfPf5SUwiN0eeycx5gb7BJb9DLHbsJoQqYR7O5l9/depkBpR8mrmDC
IfgiWcZyGda7Q+KOKl8hMyRnpKTshMUjDcKNfl59IGKHN4uqpPXR2EdbXGmxOTn+ddw5B/4ilgzp
WLaw3yCR9wUkwwVd0WpTMmmgsVx5Yz1XJ8S0r4W0RIdkT0PAO2Mw8Naln+2cTHjnlUi7ztX+6lu2
HUVJohLCAhTBhPwwtMiYiRrzIlaT6SdYC676IboVxZKjQz/1qTnVfh0iuU76xZjlAvDLsQ3Mz1rV
KTKqchyWRdwVZuEiPzmZl+gWjkponmA1cNz0UOMNh+br2A9IUF8rPg6/P32W0EUV9jj5In5YdydX
dHINrsEVKU80SdqnmTG6X7ZCqVIqH8nbMmRa8cp2lYCKsRA2iMKOGQ1Q8H9+V/p/ugVEsj4LBudC
seljsTkCas8IxIjGYiUut1jnTnTHXPFOW5SrMtsFjhHMeZeNtE344PPrKfVozknV0iWk2HkekTQ6
c+/mlgCYha7ogZatE0t7yPR5pUZeZ2D19W2LVnSd9Rqo6cQYpJi8f35ripSq9o7gmIVUCf7Ow2/T
A/k7EXjh5nbwHCEExFeDRaZjew+yd7LBOsTLWP6ozGfRd8wLD5o6mYwRzFZNcBcHT0RXF7lt0Frd
Aeb78sdw3y6bPSV9XMacBmQEXad2EW7KqWhUstIaJMFKF7DzsClQ3gABXVXcmM63F/haBHlCQk6T
f/3v3ZnIWk7wsm9iJgzQhHvItVBVYtF8cfOItjUoDPpYFV//XTlyFGkFCJTCTMr1ad+T+TPrvUzi
2oKXEAzfAB7cOuczoDNa6K5661J1AzmiY2QnMeyhyUbJUEtVvkwIIhTXwFt25BGKc9pqqX/bsaHh
ErFe/DARWStWxwgORLF3a+UUwJ7h/PQbyGDI0KWl1R53ip9guAAGQpQfe+3pqenTS5cXYLMQhDlj
9VYDSDLEfD6dllGGBd8z3MCiKX/OypleurdAHQ6AStIME7NvB1I+SrCeIJMYZ17fCS7jPSQPQWVo
YCSIFKLzl2cKe16fCPZSSxvMrsh4R2SEHmr5yL6hzWo5JNXQu8jorJfZ01zq2gOQEe/oX1zgBh7a
F+R2dWwvNtT8XaOuX34EJwsKpJ4zLU473MxATl3KZ7P7c2CQ2BQHKtzZTq4x8W4zYobIdKIffrxd
TMQOCFanTryMcYV/w3Uo1ozp2e5Eb9XU4QbNRjZPzmpcjyVQX1GIBldgaF8W8sJJfAVCxlgp3psX
Ssbhb0kAlkgvjcqC0weUr0bJj7fdSYl6Jm99jEdNhQ9tRCrypsLNYaqByBrEOmDVsfHMuRF86aUY
vtKPyAkV/Mfcy5Ec4a8O9nS1O/wv8wwnmDZIQv1qW7IaHguTi1/e9GZvc3EdG7u/VO/PXELhErwP
o1C0EI2io8/ECYsyAL+gkP9j0+aY/s6r1PbHvRQxwltLZeyrrlWPFzD/Sw4nzwjW0hHsNV4svCJk
EiLFAhvGNcEmQGU2IKC6rIivbxvoPUVMRV30IcTlPJAET54NLTeVZK2/MXOpFIwJf/UwiLLBZyPn
+1Olp/QU7me7rWun88hoaz0AqnnPN/tSxrC6vzybZsieTWVRwbF/ZaM9Ce691gsM32IUofe/9E3M
yBGtyi4yO6jSAHVny+SyRzBoXRjF11wQ+V7XcJua9NDHqjzpYRTbC/if9x10DI89SZFhJN5K008M
QIP7NzQBbZ3AhyUEzfImSDY3jNHz8J1DX3+C0y3HMSZQxvAFrkdHnWt8gZoTPs5QA7tXwOOKgVy/
YXpfwAeUEvJjtCg9iyxKYJO/Fwrl4DE3t6zsh5XoJ+EiizMSYcBoFOFyDldGjGfV5cG17wraiLpx
KSIxQsNtAUtU+Atld9sqzz/MjCPTwDSEuleW5GYGoU/NTJy5z3yBh2vFFSVY1ZzsoiSiK9bQa33o
IcKvGLBenQyCNnP2cTigsxuv22hFdv37eW2mkKrFd59s6NAYokSucHaJHWIk0nhrypW/ko/sD9Bt
po2GJLIXxzSx/Y6ysCEKzjM/N3YUBFxOrCxHiwPhQsx8xfEy20NgwooZrjmZ/1hULT4g35I0y6hC
zUU2j/4Q/lc5RPw7ACc2vjHmgE574+1RaFX0w8FOXycvbdqCOrGWiH6lLcyNnavwRxk5loRq0xyA
N3RNUCkiVEvzuxPGwYxmGpKqceo+Up+YxGK5WUtN1r9QtGOFKe5Bg0J8bGPh1n/2Urg+c3/qUQaf
JJQBk/DkeYiIjau57DVxyaj5slCLzCF9sqIB3Tj0jNM3AADG6Scay07E2jZCVLMReVTssg1WapLE
Gqi1rJR96mN33/M/rxdjBzo0zeYLm0EYD7KrdXjS0ttBJQ7WeS0bVosEFuwqKaznx969uBbvP+H3
/QqC/4Cl+rkmLNf1MNcW/aUB6uIdkxcb/lno9HMjG2KhE0S5km0+hQjLXIg7A7AFx0LuGgAgd+co
g1o3hZ/ZEDz+o5Eb43Y56wiPeKp1EudcVCxzUtOxBu5UZNSuqukkGvUWHG2fKZofDKvfRdhodLmE
marariz8LrOiSbPOAJNOn8E5WkI0b/Gy8ChF7cCQrYvBgoAjtgAL1C4KVo4vtTSdahibrCP7J11i
7KzFvPhooqP+40hIIqhkIWA7OBuks66fRGmCyvTn/D0NKEU5jp6mC8OyoIJLSs3sHZUjYOFZTRbZ
nLOl0fl2yDij4dTwnymddtBdwTnGSVcdVL8RvnP4s7Bvo+nzbcomUsxcZ6/KPm6aFYogpc3afxXs
C+C9UgUsOWo4mMVQYO7fEcKC47kEaC1Hn47P/LwmDS9MwaVW2JmHdQvMKbsVueGqBDL0ZMSrHTPZ
ya5XJJEIVYB9gCotpK8ddr5rmqf/jrfIxaxivwS0C42NXhNt2j9iB7gbRvC4iTdTNiEOFxN7eEN7
OUQ4uorKDUMcdgwP2bROTxlqDGvMpaj+KcHye1GMCtFAjkr2pHREuEiHYgTCWLI4BGmdgP2sHjdE
akdkXbDsBFF1z0hay8C2fx0U8mnAjMT4+T6HnqsqRulZgVjAmRML0Xg2CtJrvtzKuRNIEI8k+wZY
Z8Napj4gy+z5miguFIQJ5jAbU01xJLEazmIYRI4vkXqzP2sG1a0wNtIY1oqkwZd5QJX9QUvt4/kh
RM/xpdMnuYBIqG/os+5DP9liNeXCOJ6mWWYnSF8EI0H9E44DlSzxl0vNjwUSnC+UvuPpOq7YOgTw
Tg99ZniAMcba16QgqZgtq0xLaoSaKM6+Cz50Bqy5bnHrJywU1A3dx8ZNro5kPOmsGFhXs59fz5mp
TRMqzP01GF/Ig0F+ONSEG72PKm8+v83dl8vIGBxWKuupvGha7w9Mx4T0P5AuybCwyOlk+mEXTtOb
RNX7jmKodHf3/Qp34Rn5pFzcqG8u1B1QQqVFwNtql0KPVGsBV/IokRnxM5aBsMCFqJh41BpeFY5p
46sjvHaNXbN8OBVl2kwzXE8AfTmx89MbT/VdSw0YelHFsukc3ovX/W+I9KWO4qoAI/g0yfn5IlRP
LIJ8PFTtPRFypGpRStlBR51d4AkiRE3j5/kWh3EajJks7JtG274tDKcYfrrAsOBdJKk+hxGCOLhx
ZCFrun4W+sRyA3+B9m03vUD9WTRuwVH+X+xqInbLUk7aatJvYiH7GENJSt+i0sv1sJ8BtOJ3t1Sn
YI9evmyI5naeblaiT3I7RkpjqJckMGq8LmfhYBVQJ9qYbb6fsLGlfC4S4AWLHaVLxQwjXCn/kiVC
lKYE7q7j3JXY63A+B1v/xDtYzz68Q/55ttg4sV1e9t1QhYYee5xAK/IkmL55qvaoim0ycGFVe8Ki
btsXGpKnX7Si3n68va9lv+ljuH0TLJDTJZmvolUcx7HAcUmk7vBOmh2OznnJ962562BeKe2OC9Be
76WvhAnMq0c5670ClkEnW25rBFiLpPQj6jvQHdKSbqGDyZqPtRQlZ7EQVY9kD8Qos9JLNXhBa0NR
C3UrVhr5+r8YNwqlVZazAETpMl6VQcAv1cOhHHw7u/+N9qYn6FAiN+PBcOLJUgjHo6s1ZFlEVSJf
B1cSpsZltUJgwNKjR0LX6UDXRSjML24EjazcZpBkLj1eVnQd3GrC3ZWpXe3Um9mtnJNKB3R86rC+
QyuAFII3yCGVrn3xbgooEAZA1lUnzeAWNiYxxxw2+sW5IhCTCk1tFbHK8F/id/zV+fcZVWl4CtTM
KR6zgsniAiZCq165H746MXvKtf9gltQkt126PVuwd+Y8VioIljbaX8nK2dCyj/vOAQmLFZOzt35w
g0qTfpi12DQ1AP6xoaFgiL936GPjJShvOw0SdndD1tWn6iFl9dertKas8AMW74IU78L0tGBLw5nu
bWrCBKeQCHDlvE10FM+D99r1DmHIvFGTxdxbbENkRQSZjeXa0DX5f4oMem20Z/rjIwGPzzaR4ifi
oPPqQUuJn6lS89iB/dGaGzCm65pzSUy2dtLo91vJvV6SAQ9emM/GWmFmGrPhghhTklTRpKC8bAnB
RR7l95R+kWB6rlPSCHJAkreyakXggXGTU2WJ7xwQ8eTOjO2iyxjI1ET4s32NQ4F4dWcgkm7ku5Z/
In4zpf9KbECjN1+HmpIW0QjK50Uz4gXp2/Q/ujDqlUNioPebNzPpT41ejZHVz2ghLyHfKCffF3pZ
qxC++lyzDTEmDuODTgQFd0qB27JcyrLrQvt9fYLYDJwF+TVL7ax6/HtbCiNgaB6UVCN0Dnpgy3J/
K1AXORHFwZAUqc+FBmFbzD6m47Mdxmdsfd64eOlEGtWYtSNXShKaZVGtGZbLo8tUIwReXwvVnxJ0
LjQKz5Uq+mp5DuksNsjmPQZBAOPs8iR3qllT+4LqLU+2hBn611Pn5N/qN82Ft4eQJ6sWH/TRqhZp
lMQyfZGsHDw6a0hXjrW+ilNJgKUx3H1VdOAGntsivAs5ZLfVDxB7BjTP+45MqJM2Y4F5B4lhcW9Z
So94QRPBL6demGdsiF2HFVtoIblfY42SEu5CSz00wGq6+VkKDjqhK64wBTvWoWaiKpLbfTazeW2n
ehkCliHKEuOyCOc7GretYiEnuPpI5rXGBoHxEEeIZCz2SPSciE3WHFnFHLfr8mLBl/N9OeXhAte+
cDIUV+9WHJK+OkD+06kmmES0p6HxjkaveX1533IP42XzUdC5kBhZuYYd7PFbN62h/KYnhv/Uqc/M
Mgz6mIlpGfIh8YGiuk4/uGEPJ7XZszDAhTRSTf8RdS5LpJo4sTiLo0oIn9F2sFbvwfLQ+WSwtk+n
iD31XdR9jHXqAMMfurEQ9VK5xoc74bLJaBre9m8uqGVkM8IEKCjadzgiNm+ZlAVNRg0VnHlNGWxj
VVj+kaMdsfuCu4l+fqdPF72LGOYT9rwmVz2KtC8KHAmsd/QigZUjgTsFn72+mSTtAIeuzah8xJEy
WhOEndQkWeIoq7BJyfeWqfOj94ZoeZsF41FJw4q4LIblfryQWdGN2mAcuRFNCPvA1kbHg9ujk1rk
zwCtaELLiQNcXZIBPIf1yrSiNInlCU9MfrCXVMYeq+6oAqfPi2N5+wtPrFvHAWa7+0MgNJ64inBf
5FKq8r17idb2pLM/SMm/nbZeiaQtYNFbrJPqwbiKvXOaBcl+cR+Q3kbGMTThVa1aZUtRbG7Lc6/r
pXF2owUlvRs/w7SsMlFyjGYF84BJQTQhMcrahVR8YwFnCqF5VYOGWLwjSgA8hgtUvQFM9rr1fxQE
CZJogb74YwrVQpWqeusj1MCb0Vfjlvi4ZxtWELhC9xR1k4cWMlNcar6TQPHVxXz1Z1gcUxfVyGZB
d+7Al17/R/wfsa/EfIJZFvzfilB0T/DhUf58YtyQQlZLJr1P5pNb6KH9pantHDBGQDBViOb606QD
L9xSDAlCzrn+9PH/a4we6jME2Bc9dzc7FvqFQl267WnvAhjchbPggwLg31eM+ZUyOwbJGI/IQMjo
/KaHZUTLwNkp00fZFkgeAstkTEOzl8M+SIGFxlJSu0Km3cf41ZAPX+U3+fIdTzLxOG2VUfGGpBTJ
XUMXwxWAeq/83TQbQi2ZnvDwsy5AmoqYwBLad+QbfzU5+rwlMx0Kr58whEPGYo/NCczzpU6uSCz3
vAbRzUVADbL8NPVG/PmlBq/2rvnhAjAlGDtIh68T/yjROBVZ3kSOZXoD5GPoFd6KWMUkJrOkoUOf
5giUjq3ZvWW8eOy35EZu+TrjoBDS00TG12agkSK/CDbpGNeM18duBUuZ/tXcbNSDOFd5reI01pC+
wwJasfIk85ki93tniujbCyQCcxEu6zp+62MLsxvV0wBqp/mcpq63dxjRwbHyxYJuCJQA7xxNHyLh
7ViUsFynyr1Vu/XxZY156ibB8wNdtggGi8nefXM88PfCs8Y1RMDZMPdJ7aAEoVsrXRhcM1iDxd5A
FFFQ+A8y4fAWnIGX91sUbZynArmKOyvyljfyycGEvCMyy9QhA7qQ5x+H8luw1QGqBWXLpKYotLb3
bCHKcPCBTT5YV/I9iWQ2CcmeYcDf0tL7L7YZnwYBza+rl725R1UmrdVQanvkqQXm3pGtIT2pWA0d
xXP1OV+JA5ODA1pnDlC8fbcp0y/9vkkJJTYk/IXXWvr27jXVvAAb+DGbIqgFywPvdsfsHV6WhDBx
4L8IoOs9ruiJegJPzsk4fHCav88yjVYK8KtCPkizwvDmCAZmmT3jkTvjqpfQQTl8qhR46lMi0aZn
r0olLMuMmjMnyTqBVmY/kJ9XO3gjSn14tGBaispXRDGmkL7D1ERXF8YI//1JpxCA91Ur1+9omdeN
7coA7XSbB678wJZky0PXYg6tlOxXpGwcI33mGay4B1jVcpZMuPXA7qIopARuqRx9n559iZj1NC7B
9IRmiNMrr7RBrTfBSazMjtj3txmoGvyI7P05H+aqM+18oJSTf/xfpX4LRndduAAqDAx3eXLTtJCk
PpXgq8ZhaEUd1BD4O2dAz+BRNAftIowfK6VJNe9neL7IPWR6/Rn8dfWVFqGGSA3tYmR2m6Mouxwr
AjbBjV3icav9RMxx1irhgyF08gAeMeRDFhmFCrix6Hbfkphu3IyM1fK+Dq2n9vacGu4l/n0v9U6V
8LnbZTaLsR2tKI8HJMKXqP1/Hv5EI4VfYO0YWd2JF+y3lJu1Lu8/WQTeg/tv19G4n+47/4c+bAZO
NCDtsKLHxut1NeG5WtvAH6c8WriPHlLYePwXWy4OtMRRCZevMVfPzqCVpojoMkKt8YKXB56u9lri
GWbJKPR/u0O2mnSkF5zfG9gzooZas6GcGfVHitYmJe4IrexflU0e82o6CTZ+nfqUBZ0KBjQPgaq8
GIkq0MPFvnju8O1YyYMHQbLPNPi5Wlz3mPHuFgD+VlnRTApj8w+OECb/r/smtPC8hjlkA6FV3YPV
IdpOqXEzsnXeJFj+1EyzWIUJSeEGv1k25hhJrEn388FRTiGHwW6xljaMev/KzrpTPD/MRHnF2NKx
8uLpsIStkZ4SUTFVQ0n4w2aV/8TQLRNdQoudshzM3tj+Qg+bj/C/EwFGjcb//qHYcJHiSMV47DtP
a+dyizHNOonfCHNDr1yXmubzgpaxfkvFyVtRhMlRjhk0gzhlOnjAhKcaDqX7xPC4D3fMbEqYNz8e
++D6tvm5zZi4BbEc8tGUvGkw81+KDKzL57SuhbV6ubn1o4byLe001oSgvfolhS6ny4zSFzbypFbZ
wgSG7SeI/6rSgBXGEt4kj++bPpEVMtnDxxDsy9Mf/a1oywfyYSfw+kUyeX/FKdnPDg8r7+s/xLMl
iTtNgpaLGoviiqwTbJRqDFzlsRgpBffFqJhGBAw7HKxvusH34BheXaV2YBFE9fhurH1MouSrjwHM
79SgX0ch7hBbQPy2c/mxzNI3DRK98x9C19gSmUdci1BASXAiA+tJl8S5DSdkRkHQGcKc4EbwBNHM
9QfxOt+MCk4tpf2c5hZOnC02feWLWacAQYHK/YLHb5nKphQ+9URUpPaouFAr2Karnhn//LuUKCDK
Mk2BfJOdYBjZt4+Q1JRUn7bL6Gh/Fi5wi+LrTfExkRoBO81NHNJW5NuvtfFvpqf4wxx24bhGdKT5
Hf4ZIAg08DKPNbtCcLzcV3fWXvSlRQwkz9q+xPlXuxkRghObdV3IUZCnhTN5zCE4gndLhwBNU/QV
CPF4qifDa3As4JrCoOeBdMcInTg54/mixFmV4Umj09Utpik3jDlJ4x85T6AexsntnwCv+oZNK40F
KhcOneSZVezO7zniSRFaTFXGdOtgaQ+9eSs7yBdP7rRVTt4oezemRbn/MJhp6t2L91m4cmbRjp7i
USDrpYc0myFI47McldoGt1xDv61Tdu3jVbUg007XMZKsMEm8wwScJaJPoFW64PTDdikE6NALsPv2
l4sXu8RB7AduW+G2oQV8Qq0Yd/wPivr/hlf/kBcq5vLBuVgN0Fo5tz0UI18iUmkDkNl2fxOhV0gT
C/LpW135vo0SefH0oe/9mgo+cRDjoeu/cZG+yLP0FEMklFkuIVesp8SVG3mJndt3OyVhvpWr5NRx
QpnB0oxlkaKVwYm6orp75dQ4s1aQikV1hl0/mjEWuDY8r+KqmDScuVil0FUvrG4OzaIBsohm6Afr
oafj+Gj1pPzmmcMNxcFUh6fyx9eag+cRah8qLnPCQAqhQEBPo/XNDmN+gnJw8riN/cFtnZwogiVF
p/buJUO+Kaw5TyJiy8j2D1fP6Sopp2MHckLru4UHpEtCSuVDjoGojwDqG+JfTiFbnPY+1yigmneC
G1MO3CCKDa8s8ym6QErCEETk8PAsuW1ogxvtFtPF2hHEFcuU8zct/FJx/o8OhAAFwfv923zUUJq3
40hGjc7g2LzmELZqkosYIn2+F51unr3RAydU2bW5PR0l/sxkxrj3fgm7RV7EVufR5qzEw0xKodZU
bfHfdqodfAuwXLAD4IiCHWrhPjYkT8PtV1aUjH/tu7RLafs6/wiWxma8cdnbBrquqji+Jq9fzwn5
IfmGFHMb4gjubS9MwoSumXS5Tz7K4bTsDFmXjX3zbVA6TdSq9IaoEnJcT/a/tuJGOilt3hNWsgfn
QswFCe53qKpAxkJaO22hmqpdCIKieWXuyypq0CoMsEYPL9ovnxA6ULkrSzRvqtcX4DGS/0/t7dHK
8f59fvaWU1gOm/83N7Ylew0gqp8Fx6mPqYuWzgJLQXmsXT7aqwyVswdJoMysxgopnaTw9xIDvelQ
dRMcWG2RP0ssShj6PqHYQoJAcNIo6s3Hn5wn4Le6igNK6lu/6M6gaXe5zNXXVpFbzcrnyjapxcHa
iwaz1U6u5B7RzjgBTskCbw3Xp1vFS57VJOgjS8gziCBipkdOwHmnK15qoAouIy1zvnhadG6M4ocH
DDE4v1QBuziM9AXLYR/b2MxpAH401WSI8wZdN54UvKB10n0vu+fIrBDC3EkWKTIM6PIvCEV6KGH3
XDu+jlBlusYmPcHLkFEHypbwXV+QRJdaz5k8+N9xxRpWS8PtEzwJrIGRFMY62YIwr+Ya6PIqPSa5
Avvitmz9zHhyZ+QM8oW+X6NDukV5No6CJLtOZWq6TaX+RT/r1ENJVzl14u3YwVNeIYMVsI4Xy6fp
zklf8jZOX6P0Kz2AO4J1MOqvRTKMnAEsoyetyOpj+wd3rl2lL32vYEOFnElrBYqZXrsrrA0N5jrC
Dvkb/jrG4GvZyMxmgkkNAhUGW05+UH1lPunf6imVTXiDnqYENV/Ys73xwM1MPfPHFE3KmYmwnlVu
0zg375mcV4n30G8VP713IiIKz5HAAvE/L0F10ICEW1tF0eWim/Oq6VzK89WNAqCoZU4l1MkvFlJz
DZCRoMcs+hOX2X8srhdfzqLR0CMI/8dREw/Hui+WsJix81jTpUozNw9kar2awVO1N8G/tLC0eibo
IagpfVkvVoTid3/mqcZpDfngCimU+PIpzCKrUlM6Oko0e8QGvF5koh+FxgpkOyhTGsfqeGIYGRCO
ezdF92skMlE6GzWtbFssklRz0kpTDs6NOV4IjbSBqBekt/lzQxQs3t5ZY6RCs6GlneHbtw69tE0W
dvSQPwOM5E6LFtIUBjGQEdUBYkmipCc7Yd6a6IKTUFPzq7bH4ZtwzOdl/v5+zOUBireAX0oeHe6g
QBhXQBJvGDVC08P/CGqPKlRi43uWe77ekPOpBVumY+otmyVXvgCHLa+qfjc6X8J+sjbFkTMbdFaE
StyceaOksx61gbeMaG9E94B7S8hQGgLACyzGJuOsCzisvw12N3SS6WEDtP1yU7YP+HmH4AOASNEy
RZDX0RNS2lWbMccbSRZsGd31E/xuUPe/HFUAkRFt/EUu57dQ8KxfNOob/BKBM1OiXbOmwHKIYids
IGmvrnJb0cXEA+EKllq9v6LUOklGNQ0CrjrJypqMS2y7bq0BO5R84ZkgJCZKNDFJ548dzjlgS+4S
EtvoJ/2Wy/yFgOUlKvkWojRIol/8zURBG0Pxcl3I6r+yzyHCKPn59mE2RMwmYzOmeP8S0hC/xHyC
8pQ7kEDGYQVFhX83s98KeEToimY54V5Vm7DtheA3+amvNfCKCStcJZWXJ9/fG+YCnln48WVi6QdB
RMHwph9F0GjO+aknjpN3uoFnGU+7r7JtjnmUOylDULlWeNuwpyjTCZH2HBmuM9UbZLZBr2kA4L4c
6gZnFWk3jdBXZHpLOMpLfsAClc6YcdQPKwVv5XAoHzTSTCJhshhllFTnH9u7O5nrP8ESmypZW608
6ID+jQ66kRNYVqmsgqQngyv+m5c7+LRBXSpnKMIVysCxU8XrMcf2VzQmxewXNgOAw+nL4BOBifRn
GI3LufuvQ3bmSFWeFq3A2KMQZQMAb0CMHpEAtwNV+AvfJZ38QG4IbFRxHrh2IGoMQXNWYFz9lfhy
SLKTGYcRpiAHujkPJt9i1TfV+EUWZN7bhumGkpFbD/D7bAxUCOlgHVkxQxXWZHFHCoU35h8AtEeK
U8jnsoOFhkhhVJC92GidQqR3nOp0JuI2pYJMq2v6M3ZsZtT/h326nb/ZrT/8IwiSMdZ28cW3PO3a
FMhTwgstWsvIeGBcq91QJ9CqMBbAcWGy7LwNKKIDAtwZh8shI0RKx51f05CpTiTTmvKvPcwEL3VU
3Z7lryINt4ildEmEmqZpLT6nFqpUc56yxl7wbO4vliSlwuZ2sMQxgJxh5X0vQjixDlfqvv9+RRQA
eqObte1JHWZHrfugW6zMNpsHbtKIfsb75w6O8CPJEqiQV8TcEAi9GWyowTE3mEcz8LWXJHPBuIHs
Db2q+iwFWHYdfUtC7lTnDSfP/MhiVqjzg8SUI+rBlxV4bvCZeMEJNhgQYAnn3+g46ISrnq05aOuT
xyy0Y46i+FnPQW49/6XoGPJLYwCnrkaD9e9wAWiqR2VItXzAEEFRST08h/4jk+z3ggLm95P4SCMV
v84dOHhHMbaPOXxmG1sjxKmcqgs4Bcm0jRVxAse6GB+G0u4ZWiKUsd30q0+RAIJ6G/Gd4vuc1CVO
yNhZNQIkqbnHJb+CQ45TL9vEytYiI1kqMRlphX6R6R+MQIRYziIveEU+L7Zjt9PdvD0LL2hB46pE
oIiA08NG8xj21xY8qkExE2hu4cnfo796t7w2walbtr6+s27DkcBHW9TbBsu3tWp0g/ZNaBWi9cHf
GdcsyPKUvIvf7gJNRS7rfJwO766AmCDnw0n0p8Kbnw/dCg7QvqmDFHQMxeX9MroGdJfvsH3HyZxv
Vghjm/5edBQEpPSHECZi4DMaVGtAH0WpTLQF5lxxP/J1hCJiFpWvwGidRoqbfozQWLIHQCb3g/rQ
p+4/JAl7YvwYaJFlgDl3WL+3fpbnjpd0kcnmH+MF9x0ShS4jWzXISxQ/Cr+zX46AagbAeYkTHJxa
AdwXTNISw0TRkDKjMQD0i1/+B002Pw6PTO0t+Pu6zcCkbISiJ/RVn0i0B5Kxoj4vVIrtFvC2pz8Y
iK2T2ioDpNIQOIiDFA00b1idbvTTPAhriyOKHXBBrNJBXweh04RPqiZeYPWBDpw5dLSAzUrA43GW
++libQYpRtVAyCNFOko/Jy1PvE0KcNTC/zRkSWLKlFWLFl47y1PBq2ZZXCTuTEfW7LDRI8yhe5Oc
KD22Bz8vvd3BaM84yKwK6iXaD8Fu711BsVM68tedo3qqnD0Do2MenotxtNz69PG8Dm215/fISPCg
90cSpcXH8q9KMCXWORS2wc3PRDVozKb3ja7j+VvnA8kl23N+VN1Yv5uiA8upSW/0AivK772du0zy
ktOckzrhM2Ri0IiZHOAqHb3f4/uFFM7uKt+loCuN6TrzwtRlbQAzlWlNI6nHSK2v8opcpJw8Ba/R
z9U2JVjHkWrVoysyck8ntqCXb0SzgwIfAGr9wdEWTlNZV1M3sRPNntJ/qkThuIZPAtKR796/1HDB
C5cCP8TPmU3/XTMddNhb/2PbFcGyxzFpENtPFxz+d9rQDdWKB3A3pBta16kMxzeTLOwgxgdXe/em
D/vfHmyk9eZHanIOvEa2S6m1lVQNfUxQ4Pk/FPKYvM+u/AVm57w4nCppBY85niC6zpGuwByNICVh
2QZSEit2vKmLeUh4ij5AjPyR70P3pKEI6ad1EyJj8rT5EkUmLpAVXNxhU/RRwrbpwp7ZProBWWxK
jpcB3iCJmsqox4L1ueJv0LzNgGRIPuV+vqZBwzYQpGAcepjePZyEDDAWvpzxOaeWi6gGTpYx/Oi/
JW/dbKZpWf9QZLJ6I51uHiiR7EBfkHEtcFc5HgFNuQ/AIAFAV4RF6qCsj3M4l6pE20TiR0qB2C+V
nbAQ82NBNTVGpMTW9uvyuOZdiPzeUD80U9an4s6YqHxew5wf75pxbzbZpOhxPgeUQNI/GWEaUWrO
Pq0EsWE3z/RuEaoFyL0r+Wda42kny4P3jpGCXaY0iDsrQHi7AhZfe1o7mdF/u4jwjpmXqOGjPmPW
ZruOZPdWhJCYIo9W0dI1/snATKxDPsllRmIGJDeRSdukw7zPszUvDlcmRV/3iV4NGjXkYiaxZ6b1
+oReGDMEO4W+TJfN9SaZloL4Eprdl2q5lNqkK7oCl4Kb+O6VaoOw2kHRIiIf9PUo9JurpTvmHQ19
vLfqQ2A/d4+O2KzNYN7ZnFIOfPbKOG0wu3f0GaiqV40i5hEVKtMV3cNkKX7G3glgz8Fc8fQyWzXr
ekncJnWoE4zDmze52HyTTb21YXgd8ForB7QPHkVahLgr8VXJfE856KuIGZliT8yT+srEl1XMihZ3
L+briVqNzLtJ2lnEHONZLRJoTm0zsP8fCKrscdLV3KLDqi8Q1iudyrovXNqwyDKjbtIgTA6P9Mrp
SLfd5P1xtipS2X6M8e/DpimIyfdrL89j5RrVBz/YRp0xeyuziXZegPV+Y3fYALNm2Nd6UmJDMZQv
8oc6Tel9n9L3YyMGMtwOFh3lgyHQyxxSopykPgn2BDyklnavlLw7okybtJpypE5t8ESY7BQvvTGj
1Wz3Ckim6YInpmQDwcsQsFkPiKupb8Y4yP5k4d8fCOOF6eKYt8XjURouF45P4L20kbMXPGav0vGg
3J/p6zDbT33cU/K2ZTAe7w5/k5NgIYWlD4CYUzYY/L5KsKQQ5R+zjHXAIGusrK/10sSTKCaAPUxm
nZwxIpGsjQ3+rzS6r52e4pSQWhuseplj6rR7PThRIuizx5fl5Jo/AQCDaFHZllpzvZ2Qr9M4pDem
5ZrDRIy6xlYRniCDo+oHQnVeVi+p+nf1H/psCBekxULnlV6Jodh4karFKn/J7YCpvtnh+kBkIgG2
HVla2Krpl1JvKPEt8h1kYKrXV17k3CrMCTGseHB5CnHtHShK7rC5BthzWsZTPgp6lghuR3L8GabF
OnO7l2kvxdgpTRVsINxqOtpEveNXShkBB7+34PHtnqCzhM9HKZe2YlEwg2oHlw40VYt0F52SbnpQ
2/nFjg3wLdfFokjK2g3XDj54DyrA8ZFjf+OgZvM/T1amk0YY3d5oek7qzgroBy8UTxZyhuJsaiVb
AWuJoNAM0Liar5VStXJWFLId8PnQXJcP/hSOg8rPa50pQpybDutdFHDPCq6/K80nyKIGFve16ehh
pCuDxkMO+/oAacsNYGSGibTMR9NZnPynB+mjEtqjgaBsR0ih62f3imR08u1dsYkeKQVtm1z3vKl4
s2h1ZeqXnk1DFxDw8/IBAo7VxMyNrm+V0RoXMu8EKtwgf+J9JcOmS5mralD9WTfEiyUL5TcNbPko
DM2ma8zSLE+Sc3lxYijIMQ/5XySX/CBBP4cZrW9dbD+VrXUyHAT+72AK2/X6nhFdhx64XGyqJPh/
roExRkcTX7D9Uq76TxWs3gI3hDYjjFicoUT+PTH9c/jZfut+dtIk0Bx21xCmqTHuKwtLaFEQYf2L
KfFTkRrSHjJl57dM/x4SjuFGzWPTCmm14n2nDo9BQqNKpETxUG86a+5+KvS1ONgDtyEoCtJtFITT
nmKmhYueK0/VmjS3mxOFLo+EM4PpClZHEFr32OBe3Xi1AxFY7v8datOXRmPM525rizj931UBXhHg
Rl4puAg/wHFK8hol6aZdmjghqTtlCEWJ1D4zBKetk7G2AW7xmEfFqmSqQFNsMkHz+7n1FjV6gxMi
tJ8wVUNR7CmeiRK+khJTyeOpxyYvbkgzGyBt4HxmXbTX5srDNr3UtXWB4141DoMRiwyvi27mm1IA
TdYEIiQDE1ICRjmLrsYbLcE4ZlFs0X5uaCOWBM+41zw1olAAWPMQZPhM8c87tfMWgoILmEcozswp
UMgfuefWEyCZgyqVO91RYCIm60JE+5j5IziKDRqBqSlQNLJM6HOTcZC/XZ7pgKVfosS+IkFHob+U
0I+MgXQIEigB8CMwGe18Dfs9EEQY9/tdSL25K+kR77ChrVvGj/DG6OkaFEaVw9Mu2m3Lm1ZDGody
C/X0TiLRfibwrAsoTDophVBdmTWZcBE7NyK0XMkdg+NTI4S0lRk4kRcPzm3mYHooeN04nozd+Ui0
G/7nnX90htRqu4//PuhXgbPyhjRMjuCuNeYwLrVqDr8a1YcKbwCerdPeB3A5HQ5VfbHEWjmXKJtY
RTzyuMX3xjhs6ItcbtTZ0d0kYHfLVuKeTzjVlZxJkpaawGDT1WsHomy1OMdVcA3A94UM1PBjvKo2
gaSHeIKo0EGMax+7Pz/xBfVgiw8TpIMoPnInLolQkytPS3IML0bDpnITsDhyzaHygPX2SsM/Xb3/
qRymO8rU7j4v1e6jjo9Fd1Mu/r8EqLGg7ighz8ksbgm0nhvSXc8uXdcbd712hMPESxnS+M3fD44w
XLgP8fxMPm2HFncXh5lj/M9ElPFo77U0OCy3QZvd8BB46E+8OdqrX7/HYOnMIVt4zzpLvTOKkRoZ
N+tWOxjWOEIvMJLefPOWchHYDG2t3NM13KzbOk6aQxxwpEI6dXqz88mdt4DwzhhpPB0T8Njhnuo1
6gFtuI7S7lUCUvgaEJTunakpav8knp12xycHcvbcHXkKN7jLCJ2oJ9kBA0+PE0v85bjuJSuXS0kY
HOHHhptun8doNo+zEbYci8xaB+JBo6ZX/3llZVT8zUYMcpuvGRWwNb572G6K1e1MlB0/fzrADBw9
BQXLo7T38xQkpaa965ecfqoCqf0kFEaWWfBNSMcjydvJzhH8dR6HPVCt4qgvbf0zTufd5+6ZRsxj
GtSEzNpShTTY8HWLHQPhFvZFhDDcz2teUh2eFKxo0jL9hMnxVkB2SActC/ljpqw3IEE7kqNicyjt
B/gaUYY8lJYCLaQAmQ66hsw8thStG9I/se7nXJr3J8MvO8hUu2i5kPue/CL+JD2WplSSSKljY6/n
x/19Q2fAhGaleTVfw+yvuIDpUDey+HmSkLxv0XsceLiZVICTDSYFTGfIVd6FmOBIqbL4O2IKfPW6
FsdPdVxV8Omei6DYTQzBdESxUzLqRh5wp69hDMha+p9Fq1E7n/0BRPArsOLqJLT53goAf3Usr8kZ
yh09viizoEZa1Tng2dphHh9K/qLfXFPl+YJiUmyg+nbE1HZVpT3Ce5LTk5otiR+RENQjeVo7Yvmk
ltRxSJhBE+vv+JKjAZ1e+M3oyCzDa8AYlR4CFliSRu9oAG6ZcMdoANRw8wjYSeU9IOP6R320Zy/g
2P+6mxBRmAN92443GCWryGbFs5gOXUki7UVxKZ2YAV/6EipbMymcQzgIyIIt0F6ve4ihQ9HW+6wr
2bS/T08OkohHmcMDCGKuhugz6F3tiadHsq9RvNvzVp3YxZ599/ADdk7zuLSylKzZo4CrUzcSi3De
rwO86eObewLgH4CJufQID3bW9r060M1yJSpLMUT4x/ZfOmn4oHTBlos4nvvSRB+4hJb7Jooq0OOb
uwJ5Da1tfDDSrVWCtwYbiBN+ItSzRne8a0lwWkBPMz3TumXCkLUhQLncvTV9FnExIKIbnaujEe92
UBuM9C64AgjdsgMxgclEbgafNCZzONuCzAFrAU2lAvPczlQjm1nM+G4sA6yT/c8xZiXEZ/rftjn5
Q33QO0afxNWAK460i/ZsCdIERWmTURnjhIFRzsZII+9PY1X61zibtJJVzNeM7Aa1cKbkiV06bgh7
UaTd0hBqnw5CNegP6WJFta7/FPEUmD6BbWsQIMl87GQUcl8j0Gi9vBwuzS+z6u9elgu1x4HS8gEa
imEQAIfbRfe7Iwvp4lhuZqTBxN0y1EiuEl7FCSRg0HR4PS6AJnfU9xlKzcjmvyQFJCeD5SXtzDkm
3JcdzRMHESo4pLlgfvV97AmNctn9rM4wwWb+roxcwYpQ5IgWCqK5hFVcuRV/Q/8zL36lPfAlwNlr
qPVCii+L+tTLtT2Pg9D9BJlEboZH6My+SUF/3lwpo66CgamRbV4nEqpE1oftwdP5Rp9W/7uxLbiK
CfFzWJvybIn8MKlx4kU9ijzPngzCpVYLm50vD28kr2DiT36B2+A4Q+2gg4KW3Sl4VgaRKDApJh0M
srhBmDaCpPUdBY8XWTN5uhos8FpnkZGdOrj2RhT0yRaqXiZodEKdz8cGIKOp9RxPnF0mD8eyyb0m
PluptdQJGt4lgA7/48Uq6TOIXnGWhKmxF+lHJGEJ1OIS92ptdGuLaQi/jKRLF5FUDoH9/5Z0/8f6
VUPMNoLhukZrZj0VWg4+Rm8zsBOiCvMsrFKPPa3l9POJeDM25O63+7s9nBSCAWKZ5Q1xwRgiL78B
ui8742TOHQYd15dUeMFQKD2mrthmbfIXWnyv1sbnif6Gr6HjGzRFvSuUBH+aLqjWIJFMK3cR31zx
O1kYwvYhCaQe16tCROvB8wzqZpNWjs8VmJ0E/hSgZCi+uWw0OCQQHZsRabrTX7UzPipJJNmObDvH
kum1OLxsKEMR3OyCOVbUVxffF1vZ5LKBV8ioJ06a26SDtgTT0GIkdZzZiApV0cEJEXc0F4odonLc
lHsXfiv/0ICJETuOjilscP1x4LsyU/4UERNRjh5T7i0IBQ2S0i7plIjVYEDASWxzM2Biakn/+JoV
r+JGCKmiXtRxt4YNgdhborWynELg21akk2Ta0kpWscyCiIhfbEHFwXrGRhWazpKu4NPgd9eoPZq4
Em9s/5MJrlPKxGQio6ZREdMzBScuEr8Y39Y4uconlq4W8ri28snaX1wy71LQLr9hI2deqGVk9dxw
oeBprG5XUpxlbdqQQKOds0MGTSnEvtDOYVTs2XxnTPrE+odOkouk5ZJuhNtIgH76W/rSXBg5nc3S
UT7XMYYtEUK6OT1IOQ03PZW/+xRAd3NpsBpOe/4LW9DCObUTOPJCZdSBWIwECnlq7xTMJQx0Id+N
JOyi6rEuMeiRLv1rI+XnjGrrJoICWgZPkvLNGcQYlS3y2tp+y4TEOU6NNsTl0CebcFZfB6KZ0Lae
/k2evIAQRHAOnT0eYDhnwpFlNAMBy5C6/oiSInnUwOhfrKr1VJNbKuFtIM+BNXxic3+PXxRP0EGp
87W1Ec7noK2o6ylsEa2TLoQ/F/jpGhUyq94tSxM6SqjC1ARXR8oFQ2NDJKndq8i7v2r1WH4j6Zoh
K8s18cp0mIwQNZQxrsNRZ95F7Ci4GzNomcdSfedNQjo8Vz1UOwL80ndRJXHHg01/I7p1Cxh/rjVk
6VX0yS2+RdnmbXNbQnxDm48JiObdVjgbhx8EyT5eUFAqX3Wo6UVdqAOo3cHpOV0KuebotOHIdwKh
/xppJxC6YcFhkZH3oZV6Qa+RZasCzhLcCO/OqWj1tGXlMWYt6mufo6GNcyvPCZbTSlDZCH1l2TlM
x7sHIKwmscG7Yi2x6By2xWZuNbntklI5cX8dnq2yT4GLwQzWLAmHElbpeC7xlPUnmKQmdbr/umKp
HA5Qp5x5DTEtuNnvC5LBKXMCiqUGBNW6l7UykD0XbNs3+M98y2B4ki7MQkCSsGehMwmWj+QKECt9
F1uIhfD6d8+k1t+U13d0ybUXpySskPunlrSAwGAUNirGRaavCuqyX2ZrEwenU9hT/WvWWYaoaW2D
vboXQxfVSZ8oER047KUs/eRZKRmtN/AcFHcmAzcvD8D19zv34nmlfwUKeu0nJcGOA0IWnCEmkiyS
EtONhWJt8005Ur2fTlk2aDthDthYNOjkPp7jGMVRaGOa3sOBmd1XB21rA8D3sbzpq4B0D+imYs1r
wrBvmuzGi7aqkiBYvgzox+GGmKdbpisAWoBPts2Muq5fnHZqMAMqYKkm5kXdcvpON69QHh0Ked3+
eAkYpHhbI7jCJXVXfzvJ93s2Ti3UMwXtlWXIEilx8EVM2uUjRC/VIyoQLt4ZzdricjBR0UbAXEBO
hgEzJDmYeSRzEDJnnbagGu3tjOpG1DCT1j89K0r04e76QaLuTgeGJ8dLkr0V6O7dR7K1ZeDODUCX
iD8jCVA/g83abHpFJ+KHKpgu0fUWoSAxFo93z8WvZlz1hQH3T/aWuncflu8YkXfdz7GhGUxKQvHL
QR1Q1ZDeDOeKieJvdVmNFePwXfdSQOujMqdN/hhVxWLiQ810vph3F1VkGwVzufCtNnKyBGN62wkX
HCVndxxjf9oSACQRsSL8+Oap2k6uvfzQTu01s3eM3D7fBleN2Na8M1Qn/TU3Mgps/31sTXdCRxgM
qXPuh9Ls+LIS+ywk2MmQhqZjHfTWcIv2erGvRdTHA8j1Q847WtmQAfwjN4vhkcZJ2V1tL8zSvw5T
xz5umzabM7QyTHfDrWRzgpqQsSJ/5mGD3+8mSsfXaFpiFux8mMVevfw7L/sb+DtBXxAjvzmpJO2O
SPtXJw+Tyx5L7OMLYQ1HtENSdOzIN+vK/81Vn2AXYr82y378YhTS/SbhUb576D5x4S0Ky6mU6ikv
mgVWyPFWOpSrdf6uNs/V+0sMfLPO+XngRT+iupLJSoCab1OCGUn6XeeECzvjNgQyzqUIn0m6g6Ib
8ixEMa3IZ9JJiqrSdwl2UU6r8TapQw2w6FCHpMqQRaz0O5kPY+pbwvlU1YLomtgOWo11StKl3AZB
P6dw1raPmGD+441uv9FlGewZ/O03A+pRJaQx3bKuhoCAfztQaoi0Jcqq5jMPF7101y+5G3NN9DGi
prN3E1jfSJw1dApI5zPvunWJRuF1OCB4k5Rtx+8ef+tjSrICS3YYBGfyH98TJVffU+51KAMTOpZI
i7da3s/gyE6EYHTRJ2q+PTgCyKwz0Kbqm7u/Tz0Kh/vZ7C4SJCPQ8LoC2iOC6m0EAk2zCigtxQDy
W3hEvN2iBeASGluGdtZWvcdSnMMzkBGidq840981gjysstemyQXe8FD7GjOPxZFVPXwlKKwVg4Lj
dYiJPhufjFO2QKx1fxVFKt2QndrjzsoYwlOiziQclc/srXu0Jvgu2s6YXqMgVidvnt4j4GW3WMb4
m6io46ko/v1Z+w+SwjaOYuiP0hyBOMImcL+9QZhbXGBu8++P8SgOrkVLxIROJgzn3RrJwd+AYwxZ
pO5eJS9VVJpW5u5P5jBRIkjDRLlau5zLApffRo/BG46lBUt0eNu4EIU4OtyqlDcUFZovYI1N/GqK
/S5eSfZtj3UxazCgNsmAa6E7aJmWI6/Wth+qy3ecU504fqthxKhA2rm9IKk8LxbcS0O4u4H8eCpF
4eXl8d6bRdH+WzMxu9X4zhS8pRj8sRCZhi2xgMOuUPnSPsiyEd7pHgn/yhr4I87rpDSLBPAek5kQ
cQCSuO2byiBumiOP4bCTYPww16EqjJol0LmPqyoggBAsssNqTFyhKpZ1sBSC5mde28DTdpeoPtBf
WL9SM2GTJYyZEnmp9Znj9O6mpmXH4ZyUPVXLgbtlRhocIzwq3Gm5QLU6pz7AkfIlxBnkI3OQ9fh1
he01OJOKMLr6Jbq2TVByDXW80Nl1Un+twItX3L2oYMfoMinVrTijHxZPNhwhs9CUbmn1Kq4TlhvD
QclH0CjTZbXHAATUPdShAMse86yHPTapM4EJBek1zwGLOH6nif72/9VFwNIZVtWXr3lS3cxBjiY8
+e78FZDJWUdZzgEiAohtYan8vwax44SkVoQz5kFVhb89MwzoOAOdKWNdQY7B6fAifH8onditqidU
k4DApnObLm6pfTwt0nGFbjtUZdPH87m4gRXar1OB3NbYKRk0hKxjg3+DFs2oxp/E0pF1YdsXbSak
GUqH8bdfeAeIJEECokR9RYjgvp6w53UntYX/JcvR9XASmOJ1ZUyRO1auxCjbVYv/mO0p37m17odQ
YGZvm71+4noWeq6pVRK74MH3K7HsdZ6d3M/0Ef0LPC5+Z/6aJiRWu6hXhv3lXYXUrwEhZBEK1sqh
I7GEyJ+X6Vc/UfkmNmYM3tE0E9dIzS9eMGy4yLiz09SzlZQbPg84I1nSShT9I/ILhUC+GvOntDaZ
OL+C39O4tHf+r4w0vhvFxMPqPKYlnGUMBlwbVkDxgK9pvC2HIaz1vLBPkFYWLOQhee/bUOCS7A77
quW9bSqWWee+syM42E6xwaK4/i0rm10NBYPGxoqKb1GTKWlog771tOA9nJ+CIkji89Itg6tEdn01
ZDWIRvmZit5BE9Dhdk+R6AJKXAcH779n9yx6TlaO4lWldX2wTByENTbIW5fK1evhq2Y+5syWNgl/
wpXZ8AoYzLn1/Iz57PQ0dzgOhgsCA5pMINv+/JZXZDWlPg80W2HIUNFe0mnglcOXHlMMzif7UJLn
ekHaeaBc3uVWrpelZOrDoJ5DP6WKsc1fi8M50/SC0bAnIixIm9RH714Ju++Nx/AiemfANL/o4qNU
aJkai0+KlGSaVlIA7v5MnChhJxRoHb2/dlEux9+vO7IgaHlkP1ceCAeItL8BA4zrP1TgVAjickkX
JMlpsNwzuq9zUSg4uhdxZwglOl9n1itwuYqoUqAAlLTVnp85o4bTuuKKP33FO/NxBBRKX8O26JKL
AkvwpayE30M1kGI0CPU5SXkXXMXuNsFUWise2F4mVP2kTFmDKTkef+czwo1yIC1iZ2AA1OGrMxRS
mt7F9/fPpUs6p/Dw022JzAkzyYpza5RUF3waAGycLXJPtSumQToZsl2PbRYxOJq5Tnl09+TI/dEx
23yXvDuerioEfI8+qVfn+TW+bwT4x74gFORqhn+Wum79ysPv96P0LVeN6UmEXqdMwm1LM7qxQ22P
U1LfYWf3nJj2KpRkf34S7Lob1R89+Z6UNlblbgDyRUt1N5C/aBtOaxLEcimE1Vep1Im+g1bnC936
IvpcD6J8UIcMxs1/UQTOMLJ3QCiy/qrLmTPZfuVPbfS4l457pY+fOjttzl5DDnvlgJG2g8fSfKgJ
Ttbl4st7mWIGCc6AKmSMjzg8A8mz5eiCkr1pLtuWoFOMoIyVm0P9ZMtiaZkLeytYxHfNZEZRlSYm
gwb6CqQgWCFzFhYvqh1rF6aZ74W9syltEbcEB2iEpTO6PbDk74MmUnoUDSgC2Ww/GaocMXLWMbMX
SAAxMCgBM1m9ycwNe+XpO3UxLLcU24WZFYgO2adtFG2q4Yk6si4WtoVOCmYsiXTqhtKWjnuSTl16
1Yut/wiysjnVQtRqJmtDT7qn2Ax95/UMRh/+xZu7DOHb2mQkTZrCYSNFPuP51sENx9pD8hcvtKcv
Ni20Wt0alyGDZckJ3NikXiU1SiP9JeA5tVTF1C6j01kFnihF08UGQHxb2n2MpkfRZb64Zwk8oqzo
85/tiO1ot+IwHzC/KYFBJzSRFwzpoUBtZAGSfa6EctwIrIXtMJs4PFW9/8/S9ZTFDwpPln3Lh05T
X4wNJGuUKS8GBrtAHYRCUiKGDOartd1XY+uEYHLTBn7ckI/QRYjE78dS76mPLzq+52Wrg3P3W9yY
ymsxGBRcy65pNrmDI125NGI6WfalNEtM8/hBZjgVmOwvptyoD9YszBYFkWm0UJuca4+YWbnV+5vy
Hra/ResvM1T5YiKNcy00WiSgNJPz9Pn/sKT3VKHn1CuRLGC9JrrWUHnr3fVZhWmJgMlUs4CiypQk
MuV03Looizn/lloLMWHLhJVwVZ+yHJxfOe18fWC1cJ56xqhfHVMSOuY52iEnzMgw0e/kwGv/8UN5
s/w3aWxpHm4cJaJuOMJLzvXt0rk4bP4UPKqUv7yioH5h2KaqwJacB4SvL75WpJZZ9gNQNLew9Kfi
/BpW8WqfAlRFIQ+Sd+WuH5Gy7ssdpCL5dJGvRutW4ZxY7NI6Lj8XhS81gaQq9iho9ficerJdb2mu
IUyh8q18+fz8zSu9c9tr50X+goOM6i9YvOP+DKLt1GEerOfI/qO00JVCuiGs2mQt9ysmislrrSAM
r15byXrUEpaIvfDmE7jUE92bByYK+ocRznlge23xWDChV/szmKSO2JwzWgHtqRXrA4K0KRPOMNKZ
mXTwMlPZ1LzpDA8W5fKGUTeDLmx3k8wV74FE24W8B/W3YqfKoUilvjl6tH6ZN1BQNWC7nIgR7WKw
uAavWmHMeKQQYXsfHSAkVdNcjUSQcS4HQ5pzL87WUBQc1cWiGFe1HiO4ZeRVQpv3oDSYjyRPJZI9
X77K7g4RGzyD57tpfe+9Jp9jLPGH+IO9QwHRV3RoXIC/IC3fWp0L6C5QckIS3PF3V/Iyi1K66dZ0
EQ7jbCTo75H6ARw4QWDBZHMYB9aFTlatgxoig6UJUn24u8flQvPGRjMWbJCk9uK6d4xoz9fGIBaH
6mDEvncMbGy2Jy5J99U69nZRhXTeoLrpLwpJJ5YSG5rn1s5W2s1kT+RoGvG2DcKJ+1J5MBoq9GvB
FiFCsQgtZiIqR09NGPn7lbz8eG+P4BReovNsQBL4OHfWJaYvT1jB4ScvACzIdyaf0QkWP6moIvCA
8vYs0NbP3OUfv707FAm8OfqSTmYXe4RiyoSvI4BlbU8DFxLGe6ctZl6T6BnnvdDgKuzcxsLXRWoM
S+FLtIfZszu7A/DbCtXbSm5Ss9RTneNHVMBieKAsCT7E0tkqISTVFYIFnLvv3j4Uy1YHfpLgBp4c
cdnJT99Pb26vkOn03tYVwd6Nzzb/PLx+EcGzugVY9WcYbfW62+QSA8nlEH+yc8ovKnsKprqCkEmr
BRzx9745KOqFmvbN2m1EOCqTQs17S/mbdBTcwWxWDFsFE/7b+mSz7fRhkc1+PY78bI+pNpnH+fct
hJWLCXBtGE5R03lzjgZ8kiEAkRH5ljrHoOjfyFEtHIr9kAxVdnTXn/XsawatfsJQeSg84AgPxD9f
D03dG4sxqJdgkwEyiXFz9cAdCgDwg1mASV8FGtwe6m5ntnD8F4yDl9oMDE11cYGVoKlkhG8W2P9b
cK8ABg/NA6MljL1SLiD24/pEe4uKFVQCy2SNNE8FYw4R4UKe5zISFDD2HZm+b4nyzezBheoVDGGQ
Vj2+9zfu8YIGftIKsiAxex3piKLM85Kl/X7+ZLUOlBLq5tT4BqIXF68Smc9ljZ2jhrTEJsdJMIW4
6Y7Mkyg05SOHhR99F3LMPfZpxtr+IpaBZGZveWEPjb77D9oErSC6BYtA8fboWqYXGb1QWQuLHT6C
goiJ1XmEyhw0dBFvcL7LwUiurbUCPs9uFPZVsF8gcZ50t/niZX+QEMetmtZiTcJQxToj5wzsPohX
Scrksoh/0im6TJLo2T31+7cGw9ZV0MtigdOKcvBXeTrYBm0i2+CGwaIe2kN0907W11tTkIK+wWmQ
wDhv5sUVqZHjob8M5wXlizFUWxKmiOIWBNJGlWqKb2o+Tj2IJLO4xpDfo2TvNHXnZ7wfK8BVrm0v
gPFSVQVqlcRp+hc0kfeTHlsRj/YcJcyRsmp3CTGGPtmfonMEzAF6iLtrhYAIVEPEkX1CTxjtPErI
yzubajPld2QJ5YXGNv6YYJObPti62VY03BrQc3HYg74C3/kYMggVBTO4qIWYAe4a2kjixrMwK6wu
PCdWU6maCAByjBCLmzGo+IhPum/Nw2hCT77GnHq7YXFXksNJY0WhxJgOKehbfZ68Vm6J67ifFjEt
xzP/qCjDdM9Ztl1W3h3Gd0aY3F4mEqTsFcATbRzS5W4a54TAFtKyVHEZbbC3qUt5vqqLShx0fn0G
C54caPpm2NMEps+oroqQx9Z7e0VJTPesqBFsyCd92TvSiUfrUuCyUmvPALeXX624c8KiPHFO3UuZ
+ZvNleYn0fl3Cj2clttgWHg8cLgZ9yyDYX2OT7Vu4VJuZDEAR+MnFO/F0xsYrZj9YMqPRQgMmm+l
RQsQ0tb2G3NTe1jWSAd8rBtDeu1Tc5IpktNOnRfygIYlE/gsvGfAriQzxB2IQcHjyCOgHh1caMDz
WMbEkVwSUGXLee6lywO4+XlI0iyBVhWx3m8AcKFR+9eAbdSs5zjFBAv/5BNOmOWy8NZaLNHvxubC
RkUpHP5j5Ka79C9AhBOkFY1pa1l2CsrxyK6o9TGbZJ/Uyn8o9FKhgL54BuSTpq8xiHQ/kjfYDz62
elvJuma8S3Mq/hVEmXKhCEC/sPa06F3trq6z31iETTukAspz3ithIlZAMBVLVokf6uM2wEpypKzh
OzaRUCmNUZsUKzGKspWxj5iFY2RrbGvS/Sgdm7owh2U6qPS2KlHuGqRzsbS3ofq0v5gBisRvoaKs
JN5L7KQbLGxzG8RFR6GLQVnTDyc5aGZriFd6DiaV5S9zEdhMhkuD6ZQZH9kDFi6YIrOmEZVR7PwR
UYKCstrq5FMRGeGcnrXx1+GOVPXv0n3vjMok1rJdD+W1RzIpaIG3casVqZOaPOuRB1LI7kSmoVhO
jk1PUV0GaPhn50Jy3v6yrBKNfN/BP3XVMvNVwUQJ6vAJYtx2qNEwFoARbfCFFznj9xJMLqlJ6nhe
RKLd5CMULwjqM72aHcyeYWVORB38YHV+WK+dktTG5UwfPVIWOZcqf+jo5s/5uaVXOqmIWo1qE/bE
dVvhHQMQtn9MQi86ntc8UPamMS7/g9sX/qyV8i+ahspB8aWU/v5RE+91p8rgwXyMPyfMTq4V5Wji
dGhXdJOzbNjsGmsHBBrQNjw2PWEljH1zVX7nQtnRXLopKVprEPut6ykBzyfpEq5VkAZ5Gnj8J2EX
ib3228UWcULAid9hGjn42RSobJlOTfKVm84qTNCa2K2eg2gFEI3p2focEeHdFVbzDeeEm4YsC0Tj
3zMNoyzyiQSmyCxFR8baqaDU2bxNnvcxrdGlIYnGGhnide6ZNCGuQSCnRlv6qfHLT5JJr350oBQC
36a83dKRol2MMfRlw7MPstrrpu/w7vsup7gFvzrDym/3jbzCE9G/h8kCRH5GXSHbx5bmGZLFyVQO
CyfuWT/tEa9FHGOGguNYlhIYsPVYIPgdxyI7WmHt9LenUObjAue0n9LnIm0Fx5A/eMG7KMyDA0hL
n1rPPB5dK1DwaEz574lxkh9v1PaD0EKXOjMVt7XO9DNZogA4VRGWe3n456evADeoNK8/IDYeKUOc
dRvxD+xCrN8qKp61MMXRZaYg3Bew1Q2PikBTUI07t8TaHCI7kwaK9GGpaHDXMIHNmWpDlGpRSPgg
qIrtO7Kn68n4Z6oDMQ3TnkFh/mInI2EolWeP4xDxIz9AppCJ5Hqzv2twFV0ZnZ6PFzBrvqq7GrOX
CV87mahTk5u/wNem9lN+dTEH/YBnll6us16jFzvA3kpjHnQ423uSLSm1WPlakLLt+Z56FaoNUADY
JaHLwxRNRzfM0GAoIclDNuRisN0cVUT7v7YW50zRwYdSf2QGvv/fDuTpjzd70yIMe2tu3EOuEMUC
LpGEh8zs2ZsSAXQbIF4QtAQKHlI0k9r6vPdH8OJZwLBlSPNdfmjKRl+CU+t3T5O792FjvT/m4h88
ZzJQk3tr4ah0Els2cqUti+lHNobxCoi1O93LyWbh74+8wsJCwFEaWzfMcKPkqM2I3BjVKRHnd2UD
BsOUiiC3HMdmt6kF7auw2H93ZzwCoMngv94noqcPoJfBQrNNbZ+1/06kMiwzjM1sgWZZLnG8o23m
cqWd1qGYIaO3VwzChm+LnFA+fbvnUINg92uesG9QhPePTxBFS5sfe78F5DsUygLJwaTmsls3YEfr
JpVFzAdg+2KBCXqJcdouMSdTrE0QBXgUzomSfyeQRwxLDsvaW4kJmQWra3bHGGljgbr/rBRsWaWP
3WDoYooDRXkmyisTQ4nJQb9OpgecnZ74dWjs/CWt9cOYswxyWvq1k1p5MioBzI7R0yCyqlgHGPeW
2d3HnFqe3BdABXUShRhAtF6RKj1XX9exHtAz+yRIqX22s6cige6sfMiKR3XfYwXjfPyMF83jRVq8
8BC8AVUCZVQiBL4a5emLhKzbiugwpgd5s75uNGfEgE9EzDNSEdRHUyoESragg3053xnY+6j/PS68
fUhz5FKUKgy7W3KzKMHpPcrEkCpWV/SF9PSU97PWxZu83r60E5n11I0kLhuTzccGFgGUwh/Fo3Rx
5wMVVvuBDJv6WZJ/vSlgPmPHv4s9kOfcOAnaiLr0+QJ9nzVLOrb8YV6URIFzooIe3/NFto2mfEsp
HLLNUcdZ9Kl+QqHsR+zMr/Br+A2Fqiej5LN1ub+qFGXwUCXZsDS0q3vFIJPTu0sEMwgRKOITh2yG
4IQgJ6C8x0NWpdvb6IRxM6o1XlyD8RsQYFHd8KfMcq4PprEdRJNb7RoPrJOv65Gxavp+nS3ApShv
wEAFZSroRT4D242UDkJwcYuu/vqF8D65OiJGz/TTjUPZQDiVpdB+t760N1Qg+J1EPMyTg+N4a7Xp
ja3NLQ1jTjNxYkBnALf/MzodEZJ6OY/abrQT/JQbfrs9U0L6z104z41jB4ihjtXs00FtLUPhDggj
AY8YMBMMWj+R2GaMyWBvgjHf3PTOHycKTPmaF3N440pS7DSZZmLVAS7eWOoWIlMLJUOuu5iAvh6O
3D/+NMMQyxpfZcWrTbEd5b2M+5l4GKANS/qTpwrj4s6nA3BYQOqSHrHqnYmlRc8Gexc2OUTmpRj3
UcEyUMV3R6J7ZYmofoJoYZlO48n9a1fnBfegS1rqnqJT9Tb5F33b/dbxJq/PsIApo7NBsJrDofJd
DuIHRvuKR+hbnv8hxaGeSqa2zM/W17EWl51sNHQ5mOpDmYqDexQiWaS2dBw2D1ZvGj1rSLA2+jKD
ctBEtrUPACwL8qRyn/+z85DV+7yz79ORsAuPKnfEpGcjb20Fm0ezCmxGsp9qth8lufWqxB5yxjAA
JAFzS14Asf4z0OziqXUZKc2m7QVsJIyPH0w4v4ZnU4ymtJpzSE6MUm2AzpK86VQ5GXvyacbTeNSZ
aLQG5KmgF+RagOdlDCC5cpKJ95KvLZ3MGW4WU1WtTsfpB/7T1zk2HJ9Kaauh0kFVhkMVtK2NdEAL
XW8RB/A8+hc3Fm1P168PjJKsMAHuFwa7Ri8lbwCwHz5QYqgDhuX8/47ybji3YfOdQ812tP26FFC1
4/wmidwDv+13LDX0oL3TShuhSCV58k5xNIWxVn26UrRzJ6H+HPDRcsxQz5oUM37QH4QaR6ctWU/2
FmtuihrjPyjG2w1dAyqm498grs4Ahq1mpLMtyynp31loqjhGl7rWC63cEXprw3eKt9YNl5OiUFLA
6yEGJebxdSAf+sdShUnwcUCyf1j6OBcM+EP5m6wk51M02hGMuExBKxOqYJyYzxqVn8zxms8DiEet
6FVk93vX5repjEtq4HsFkj60yXN9WqvsxzQrEtTHIsC6JBLHh+apZJgLzHhGe7FC2QBIQA8z4diA
RRSRfA2jflo90WwzofKMvmzkgu7JBXyya1yyy2SHZDaPLkasgaQjbkT3vC2TJNieOc8k5MF031g+
XCgXwDydtrxzFR2M0RJnHnWyZQfRuq7/dWiaomCQmwyJdAIRpFgqQ/sC6k8V8vGa/1fXgXQCOZpJ
xmukU6UDm6/Y1mOLhcPQ/pyym4+cUT6Sxue+7FT3f84W2Ri5LnwX2cBW/VywDKvJCjlWKNiQhfOb
ssCEzrnWi3EKBgDz/Eh9SCTffZGLgmWjzqFqGJoqhCrVEjPwNQyud6zSNGweSvLgun1RPsZFR4mK
29r1asVh52Y81euioGEFqNBISGsNm3nrZVhPTIcIIpk44uyaixaL0Tv3z9Tjdlq+cC8bCCystTGX
mZ7hPm79z3y4fmT4MMK5B6+EDe7EHEkBzrE97MvkuL8SpuJPdXZwwMTdAreWTKpkFCM3deqvE/4z
33q3NC58vqL1xnpC5DZ9bLxWQd8r3dGh7mmp7WqYhY0LJvnAg/TqIp6ESozl/RgerYUDFkk8WBi0
iqlGu7BfFZTDNRxrFaUBEpXwHq0Nn09a8ye9V4Hoj1y50pGNhKKJrg9s6jvDAdj8dLJoBLEAV4G/
9Z63DAqBhjBDzdVsRTyeY/gDu+2VCwTx44s07XR5ZORXLmQr18D2RvUs6M0D1Gpj7wmqavV9pajx
LOLsjRwKPmL368HUN5GSeCIZhZoOWDYJ+BJ98nPUlEmAB2igbAVbyDHyRyg4NB24IEqcjY++CaJ+
nmgeOpNwByMfflYvBFsLxmQCEZ14Hw3Zg425WJ+x2E8f3ZlWDb+Tc+6Ks9PH4jjwhliwa2+YkW+U
F+1sG3cxr9l/yCbqRhY6WfvGRYqZmyRegVuygE13eQNw1Rm5Eg4LKjPHUdJSgAwUIpDKsIDJjvJp
XwPBp/FCtHuJPcAiN70QeAMEa9SX1KtIDsUNWNpuw26hv9udSRtWTdGsO3DJj2tZUUNkhcsA0/jq
k3L833YhalFsHDKnwPH2el257KSJB8x14tk/6nPajwKZCJzHkKXpshvxpkf4MGyU6QbRtP4gSqL0
1AJqldKdnZ7KUwpZAOw1yJQFHCCehOq9F5ziOH1kL0oa7DZuuY2hWYjYs0m5+uXOSIn7NrqncUSa
aziV3GVlDBnHLw3Qp7NHwn7k2XT49GR80AMbwwBNeHNh8FA/dx1u0cnPyTOID7DUCe1CRZzh57yf
50SUTRTwBHaqs8FhG1ocw5t1Y/VkslgQfrhu0qCcAJALeX6PqFc3hYC3tznlwYsc6dL7P6oMqff7
qDeb/3rEYqJ6mVwaUDOPbU4M6c/9EAHnQwkgoq9l5/EHfQ3KC4GprbFGOPqT3BWSvYjAjVW6BMPq
dlErru8SNfOZJeWFKxodD8eCVtzZFtUDRDsp9lcOf/OlokdLVZC4YFBxAQjZusYnpM61ft9Qpe98
FY/kmvqxFQcKFlbhS+bA559UOg5BmMIGpf60AT1wKSt/Psd1PXJzwLAtKOKyb7XEHT0socgqIysC
vVgUcs9Gu++pw1piWyhlWhCPOa6mPRMCQD7pcDhdvk7t0/8/IbFP4N3oowylOaljek0EvmT6rw5G
KFg0b1weVd7hMx68Mxqc8eCF+EbNwQYiZs+vvFFznUe/gVeceFOTTlU1zeAiYZ07gDii6tNL5CTP
SBdCYsar+v6ZzqvxntQLatYwNPNXI4EJiGxcXouJSTjpX1BCUND8Vr8Pv9Ct2hV3NwM9oExFtJHa
i2azQ98L7ODN1T6zRcsYaAd9m4oPcdJQKywpsyRz67BbQF+DT1sZx6Ll1Gip3P183YwM7g1puiBS
58c38OTHllqIS4JMnVmsyWm5j1J70s9aqUQP5WNyN/atHH/X5zSvLNE4pz61P8uU/qWzDaIJn5gl
vsdU2sBbHDoCqsV7YdbyLjb1zTtJsDvU0I4cklT6WBQIJOq6sBwkCGsDVKLxU6u2WPdEpP3Wexb0
6HhWICH6YZMI47R5eVNCIhA85B78i+z3wjD+w+Jp6nRR3j5Xbj8TzGCg4lHzThU/bSA3heYndY6C
CbjfeoCdOYBv0ObOznNhpUg9RYrCkPqd2vQKRC53VbfszbZGqYuuaEBWiaU63f2yr8CkU5CNtXdf
gt2hOtQ7J9pFNF58DZKUo3hLQdQRLGIYXhPL46E53zsJDMloGTVOIxKw5cvgmKazJwlipICfCWtb
tT74ieSSoR17XCNhEMvnvTsQCBDCjuZHLmPMROL3w4OBoYlCo/6BqnAyEql23wiIzLEvY6KnpkND
WII79CpXUc533+F3ucAlrdc5NOmjlNCfDMKzblCeKb2cJxyKLp23bq6iZ4rC2ywH4r4RsJJMSQM3
xA7Q+NVXl0D5BPBFvbiKh20/IJGV3DxA24jbLGCClTJhiv4BBXu2H1jMi9KIrmugE6548v5RNIlW
bb9FwWz9d0nvh8CNsqhUt5X85ZDy/6Y11nRZOwtC1j9/Lx2V/KO71S2FJEG4UcDTJvpaxjMnOKRk
ZH/z6jjqFk98smeR4Exz9y2t0GRCgjXPuDTOfmZRTBdcUOc7QzHAvTzLQ2kOyNf9MORoSZ7olepm
3itokHj2xcXfRfY49d/5gcTaBFldI+MngtRrFWJO+qL4PRdx9ySVdWD/rwEjbbR5q3Q0OpYdczL5
hMdgMC36rF4Sc8UT7wODtkXAWtLKvzNf/9e6oy008z2dKvUnOUkOwdk6XuhQ0j99jGqRCn4Krjf7
Ax+A0LrY3zDYu6+0INrtPUUy3KX28o9nI9GMeZ/YbIcUAylwtPAqjU33b7FMEaHD3HzLXazCKx7G
RVEtK1DGIcvk5P/bE84Wp53vp14pZ28oZXV3YPATHxtiWHbQr7Us5fQXR0xexip0Q5rj1ZqPbrPu
RtZAza8jEbUHE9kzAkgvtZD6jY7HkhHGIXSAph42RTm4LfkxG34wzeW29tdFwVHKl9ROcP16DZF7
f+hcQGRyuR13o3T/FfL3pCLKBTYTHO+p7nksOB5IxdAHXPZ9o1zWHjgwQ9aTaQPYIzm07s5YbrkR
X1twFzoa4EW36aOOtFqZoZ2OGVu76aNCddnvqvEZixmjtBeFgoOE9QzsA11skPi4u9LTynRgWtkn
DqBgM6OlKpfU6zBnvqV1Y1++06rgYMsq2nLiGUi2lJwfIIFtg4D8MiZ8e57aCh1f6KuF8mfJiTG8
mPDptTJg6a/Us0OGTBGPQhYx+eSW/ZGtJe+Wpl8H/ZZT8Heh0vUAjnvsxwvHPFMGCWdn2tLFrPTG
3j5Y/jcs7OI/PYz9W6bHPO0Mm0jBHVEzi8s7lh1OOz32Wit7C2OD5RTUsyCKP3lbI6luJZ85Pqvm
hsmxA5zmxI4TngxL8h8CIjt/MSro4Tbh6uB2Af6KNhjaHTAbNxtgRTWFzdq4rNLjx2c2aLYaQskE
IPXjJjTm8ZRAJ/Modj0E6akfmsqiB0vvkQ3l4PVRKUWVZsaTMU3Rj6YV8QsLWqnL/Xzzzc3GumcR
rJy/qc6OHLkxX4v+W+utR9mG6nMe8thkalJityhptSQ5k/oS9xv8blJx7JnhEznf0UO/sttB4RQe
c3Ol9/iAFm/L4auejZLw+9anBkTQkKhfOy9lswrFq9XOiFktENC3eH24E+ePJmacdKU21kKvuKPa
sjFRENUEwz/RWblT/quIhcbkioUfdvdsJ31d6PZ5hEiftJe+TfGvmWMrWCnRBMK8cmKi2R+CGGLv
uZTl6YUaXLQlGWxmwjN6uYngv5eni1QE7GfRQ7KyLE2Y2m9jWgKuppxAAliA4SXvKj1+pqXf+WCH
3y47qmnnl0dGzt7ix+cFt4eWgevLqjN3uaf+Jp3d5QQovXG49qxD6xuzgzpgzmvNX+qOG3qAU/6W
qQI7F67/g8UkLEVSb02inaDFBVA+vfd/wrcrUKXkCaWe7WQbPlCoYoYcfU2o6pAw/FVf4V0Cf6Pv
bcQknlpFgGp3f30ByfVcCkwM/mUGRuiioNMQv2elBrktMg2gfLwOGGkvPzNZAqgVk4Jik7MEPYvX
qyHnUgh5gC1Lgdj3SSYawymxQXHkcixDDvyx1e0MDMMOt+HJo5ueakgYMhqQf29VMmm/ANoCZoT1
1zWkJhJNZk9qjw+8QQNL4v1Y5bRl1KpLVdNHhq/m0zTVYmp7KXo/UqjaWtVcfcdBlH1dox1ljMzP
F/BwzJgcnyIfcbEMmW5l7Y/gtDOePUpELw7fYJBNJDrREjBc6sRT9IcPLs5ZpGG5RFQtikzw4jlX
ka2hTgfFWSFPK2saKJj7Sh2fV3tWNyDu6UOzZ3S9mjIVXjtFxJsC6sAm7xIAC2djZJPLR9ztwhmz
8clCB3P2GY+ov1R47Khj549v1sOxYK3AM5sMSdsBY50RKYb3m0mTH7cNmg4zZkkSYS9yvhcbJhFZ
QAh0kI2n2ksIX6vI/98SggzwT97HNviva0oNHGkCyopbfppa+9KcITvDkUC65bbOAFw3Z/3j3pwL
tFxsMMIGyHc3Y5mUIeitLMe+2rCUaWcAvQJox5ftGKhIJuaW0IxSo2FuX3Pwxtn315m5bZVo+RFz
2rm5mQok1AqV3kRlFLQVAnEmLxbePIYVxN+HzUVsH/Q1mz/Miqy+jh6+T2SZB3DmaNhHe6GLX3G7
XE7dznAEs17fV5r4OQWOP36mxSpFUIq6vWbUrEKo3BjamoNIipn/+wcy6k+vRzKpCSkNUcegu1sX
LbhLCZAJk9OQqVt+xbGOBlhl/vIRZkWoF2UPenEeMiqGpQaCGfxxH9wpT/kdlQ/4LksO+x4zZtox
T4NW2H2ALGygFDUGLwmStBQ5iB4n1Gq+i4Ygow9QJvi8BmTsopRqjMUxZyRa9vWMN+igBnIArR1J
kijXBdyT5yWUsyxxgS1RiecuRIJqvRgSKpFS/AaAMrA7JGwPvXo7xm8Sx+e5tRPGoPsipvdxORwu
1BNb4ilQLXsuPrNB09BdsBDycLUwvnzJT8pTdSxwZZvbrZ7s5w8R+ntxjFL/3XBIhoizuam8Hlh7
kT+/4jOrYcQVHVviXp3F0DOGgx5/VLcbN/b8kNuWn937KiC5jzyS70oMTgLzh3LVRggbAMxKxG7W
GjR0SFX8u5LRVmPhCg1N4JDsM8BwtGrUXTNK5WEhOupebBkVaaLU1+QU35KHjfkbxEuj42p95Uif
pE0CN3/T4nIkQWAZACDSu4v7y8wi2/eXg8ebnUGDuvT6yhYJwKW1G3my1owanSx8hwyJhVxl/4zr
zWpueNd11NyuQkfVOKSx4qh+vqUdLTBpJTcuRvqi9BTInwr+Wt/FoKkutmLSeoOy3hYE32WPE+dP
8llnKrYjvM0PlVIPbLTwBv6XKyhZz4oCh7wd30yG/OlKJEuzGQgMC1lG4HOQqgnkAJ946g0SWc+e
DF/G0vs17BGvbXlnqRPC/t63kVefvOD68xK97cZ8cs4lNezkEi5px5dP3f4zCfFtaFIsQbR71+lL
y4VxldzIdjA3upq4mI/QZDlKfABox2rbvA4g/ZppSzYCYBdSnrawmPqh2KgjPzW4peNPMg5lPNB0
FM/pWXhfkA/FhNqYUfas9TjvVTeof5wThaffyG6/w0FEYJ4p1F+ebndKlrOviCnl7HjrSh9sWUmv
S0T0CFp2pSSO+BWc1dNEPg2ot/jNrFwVI8kHWw+27uecxYqPB3rnEUvlryeiJrUgwRshLZyqW4w9
4U85YisU9mldIxmD2K+e4vjGncBnLNxDs/Qjzze9z2/gM3L3EP7PjF3WLPwJ1pseFHf5JWz3kGrY
G2DSPN7Qd6ulD9AplC1mznNGTjNZbTk7yNHuSg7WRuOUIBW4CuUjzxxbJU4f+ytKX0TrSvp+ahgD
I/kwmNv5ygjB7lreyXso1U9BK2D3N/T3TbpxZvwX61MY1tQiWk8jlN+OtTu3dHPGPIMETWP2U4Jc
fXfirKz+1nZlqVhlB5Yhv0cQnzh4jEM7QYM22Rvp5OsRkCQHAGQTJBg7R/R9Pwr6kBwNMB/aWpg6
Bz2xBbTSVlcfg7Cu9B2o7HYGB0yzHF0RQ5PghS1pKSkDPuLjoFTcTbCjzlmGoSxT2yspjxWrxFb1
KYLpmV/uuJpKygaBefPnDRt0Sc+Da7rzhneKR+riRcpSvPSnUKAmcAKUup2sc0oEfPcUtpXx4QoK
+8/HdB0zoMO0z9Y6trDYBlk/rXKyoGQFjKtKgZ7RckeZE+XmzgELj+hZ5mODpCnfyHfQZ3DTVXCe
RCn1sgv0zuRZ5r4pv9Q+RhJ3y7tzlbBUsB61zXHQruJrWPWoUmgr+rUrsSZKf3uOynssPlkEeshk
8re5OzTcUftSwfz9x7nT/HKyLnFGz7LlOU6m7tcNp1Uw37x26frfrsqDeI7zcNU0aOsKBGz4XHK1
zaSzebHup1UVKwlN6cFoK12iIvjiRqDuLlAvBvEVmZ1Q9IiYwXrhKMFKp/pypZXO/yFX9Z1nZtYC
Yd2MRIUBWhKaXwlwhy1UgGJ2CHyjodGGD/H1R6qV/bNAsLMYnMnVt6mDLOc46IXsstJBhT1Myt4G
yEKwkmf551oOt0ejiTrvsk6fLAE0epidw2cZVHg+fPp7yqmaSc5r7NVxOytbP9sIrJd2kvkKCoV1
NruKcPOhijhEq+EQS1Igpn93AVpKyKD+k+qlbUpaxDKwjRk6S4QA6eXua3Kdgt5gF0xEbHtDCQ4E
aH/8MT7xwoGkJQl3arC2CH7fk1dBq80nWcziu30FUgP29MTrYPW5gKF9eWu/nvQyQGjkpfbz8dKV
lfmbmlv6fas5sbx1Kc+3iIfkFW/ghWrxfgU0ste7L96hPJlbesvc+4Wh9QTSWsF4GrU/HHXtZ933
5nWOt/Vgr3yVp2hkbU97Zqhv3/xK6btLs95RpxwYg7z/LjKkXpbsR6R23ZwviHgD1uc+vi47edqy
MHoi3YKRTj0CnwYVpX0SAU4wjX7BG+znCOA4ZLJ3qQzd1SN5+7GI/Iz9p4woJqepNNtUGDQSD+48
fQh7mORl6DxlbjGxIj81fAP0xSkA5uEdMZCRpUjoXUM/zNX2ggAR6i33+m5icOqE+gE3JmSTVzhY
tqGQLizPzVbZWy5SZY/LGuX9v/nyxYlipTGEPxdVTDFSg7HBRMUs0vKK7JIel2klDBojFdhbu2x0
3xh7bcwMO5rNTHauSM2ywc5e8v1fxtFywFou+EcbOqncoQzARxeNbdfOeRBdhYdwHdOADur8EQj1
k65DrSb6A/dyoJW9/B2BLwky3o/Z4kC95dcRtsE+YGLY1NH52j2ukvCWedHgyWNz5kEfoRspL+7U
6eJwOpYMVvAQUJGJ94krSLidjJIbikcuGFtYCh3i2T/AP3gG1li6Q4/IKiQbv+Wk1C6JqtxwTeJX
7pwN7Hfbyayl10p8vePZmMuvoeMJF38G2JQYDmtI4RiSgR4UIh4TEzUWE6IiM6qBZT1VpxTAcDsK
QjzEniLfQX8FHziHqvAO9u9slr5o1BTkDiabBHcHxM2zMFWAHaqbn6xbc7vWg9Z7MJiCinvKFhDN
kdWuGHxuRYYW/6zq5JKreBbgQaVJCKc5Kpjjf05mAHvjyimB+RgWw836toVQ3YBFfX4URtIhC2Ft
PAHpd6RIAA7sNa4eUe3Q/TVVgGOXkJV9iAzTLmTyOf0fFq1wJxn2Fwk+907EPkvNSi+4W1uD8oe6
+ywkwG7RQVOWXKxASvnKBPv1G4cGKOJRVJ6xVpEANhtq3mAjdBJ05aZfdDpoPE+NA6XwmxQCze4T
YBLFkXFtZtvRVHADrHjf2+zP/0uRkUpkTRdAFKxrKi1cPTNDaJsGFLMbf2mTl1Kc+pvA/0w7cLNh
NXdWi/LU8U7sKmV3pchjLP48k77WAmsPJj+pHAVyXYtnqGyvPUH+v0wm7/B6SH75Bh7I5tzaHwPX
IM/c87mCRpG/0ushsLa0Bt/FqY0YdggQZt9qNkfsq0P8d3xOQER6c8XuWPwYlXPmnshX4oQzJsTl
AWuKXJFZnlHLi+I1oBEE7ZTsKngMdO0OeUQXMD5tH2unE44av/R0G7pNeKQNARx7coz5gYSAh7FE
x5OatKQmNfYunUavt0nkJDfP6qT/w8G3fhyJuFU1TG3iwEwr1Xc7MJer58yW4+y9q7DlBtlQM/Kl
GJ8tqLxGGEUbZ4l8GyVJsPmhiZjaXM9EBRgqpxfuC1gcuZrvdfjtpV0ZIpSW94335CGBJMrWrWlK
9/7uzXu4nc37Gn0CPfVzEr1Rx5uiIrUHfqbiKhn4W91TOsrv7ZyCt/XxRbHVSMpqldhZwYYlom7P
iNRQ02rpY1mmA4WawX0sHvmUWxbHXas0KioYWs+GPFMOpcJeDOI+aiSDvDTpzPjmsVpIjtKAiC1w
urCswfBrfBV6gyvwfNcGyDbvk/Lx/6xveA8NPSOMUhllxAr/1tDH7hO+faKeb8zPuKAfNbWJhelD
DROMr811mcIF5OL/h0NhaUvhKPye+YM8zodS64xzMRIaAB34fQm9DoPdqy0HK33FM6RPiUMDN7zF
fYMeLTc7HbQ9JVp09fD/Oe0mHc1y8saJe+L28NRZzZWWzfV2/CHNyxL4nSqNarUdbqKqJgNbmXSU
2GlopVNVu+howwWGe5RhDvVZ4H3Me73XpQ+dkUZD+N5dT0AopRO47RfxPiTwQ7vwGImsvDawaRtn
SVB4ea1vMeRcQUVay3QL11UP7H4vZehwPtwfDQYQkCJQ0Z0LTg1IqW/M9VgQT/d645hBEVqTm75G
yU49je26U8hA5Ei3kmEa+zbnO+RIIqP4u2oPzCMcn3UQWXEyh0JlOVaL8BZm4/mY129m320tO//D
PoLc095BTfLbP9ReKWxn9I27jk7H7u6Q6RsVKoBYE2Bmp9h8Q2NSWKXppxRKJ5bWeeIJ4EitJZ4m
as8reut1foxwpF6Y3KKFvMFYfUSlokFi/62CVfh7L6ed2A3dC2h1loDRHZfZra4c/sCvZYqea5MG
Napl8tXi/JI6EsEiA47kTc5ajgQGxs5r0Ju9JXvOEcsBcDo3ZSRrNB+fWKEydab/okBncdjBfdzx
V8QvvfUqupFipZvUVSDLjO+B2Cck6L3LHtRZYpqlJl8xGTQ6yYDQx6IrFHFHsfFCOt3c4hoUd8GN
zDZLpDmQaLXapb4FQfo3A2b5bioETX+O7Gt7O2NxJvXOYzCbzuJjYC1y44MwVL3dpqU2HyCHiapg
H3bIPfW6ZhvDzyZTTNhM+wuDanAkzzt1lpUPAW/eY89s2pvtPqVZBNg1fA//VcVyh3zGs+vnvWWT
WVPIsltdzxYIf9HYzGUfv8+RvvWAFvhg6U0jVq9pbapC9/38a1uokOnegWaNUSaEDi+/V3sSk91v
ADNlji1DEAxODPjDIkhiF0gpR36BzKabqWaicNNcTNHuWqlFc2TCdPKALCLI6oev5SOL2xPK9nA0
2nr/EwYFj1VUz7aXNgYMvsTI1nR1FHgDugZ3E33p089JFM/jGCH8m7jjLhI49coKjBcvEXYTqKlM
P2QLlQcio9ACuLXY7XWH52iydjLq/cvFdxUmikuGn921IFWmFBn/NqHNhjiFtrpKc/BmF4LPNW1M
8eG+nFphf4vWMwMmq3VU8+rdJqnmecZHgD4kOBC1NG8anIX4qL5hUTyVbGr7qYPpCEriqTulghOn
9XDUS+7M4KCL5nhEBC8/QpqWgkbfSzafqSrRNhYNOYH59RBH+H6kOGx2gZsJMcOR4S1gRt15VM0n
TvbVursfw5bhFljiHAEbXWAC/7ll/9+pHaBuq+4av1NHrsXjRj4cgT0j+0sq+NLn+cJHzBaupIi8
Sm5WruLHm5obGoW5Ekzu97og74jk7s9Oql3l3UCnuk38byrf7rmx2r72xzxGP7+O4YVuDKpmlE4r
Jpt9V1ZPNLpgCScJ3GbWtGbgtrpuG4joqpuicr1y41lk/hOjIEX9jwdxjs4dFaSab7cLe06m3mPh
lluM3/HAb6qFKwSkoMazu9yUioTgI0o5kykVKnCxROpjJXo2YiYYG28u7a2uZeAvLAVzUViyngp/
C7MQVPx3SxIi0M7CfLNVbSRkL43Gdnk5VEAwxj1ZlqbTl2x4MnM40w3CanPam2OUZV/Pz1J34npz
rNIYu1z4IGlVKNvDAlCIXQ4KzabO7CpIKqYtAj9ZpG4UThfKFON17Q7QD4ouRGycxvKXu26CN8E8
yZXcOADFnZUeyAjqE0mELYvMILMAoSqNKCuObLDERZXOHCfo/YF9lgqrlcZeLhP7CIa9RR6wCq/P
V7TUm9HPxVezjgiLK+Dn91jLfVDYVvCRZPfCisCKtbne7h1KJC0r0F8uqjYzhmq1MJ+eB9LfS60b
PovR1ZSjPBP6zTXYh1OF0QFmFEzbFdqPlNCZsKwfu1VNwxc5SwO042mJ0JkhY8eSp5r4Bv4UQJuY
G5C7+XMJcY4lVTzTnCOXColr0VzJURllzTtT/+g1HLIZLss+5QyqA+07Ob0Ww7OpK/WBCMaHRtFi
zD0z169nXKz6gCnrXTfWvk2CR+wHKiM0urz2s7q0GOP0KtU9IR0V94vs6Db+o+ER8v5GZ+YP78RV
trhoLdXYkI13t7wxguZuswsoQ4zwnBF95ao52EbRBbJukpRkz5GPwyXh5xxxNIBgf6UYsl7rC37I
JdWxtj+uKtQsKJd574sO742U3xkm8UEFzRl0Nyt8bg44U3FmaCZpOi9U4D6uLzR/ICAkCeyz2GnQ
09OgQ5lDo0/1QbEwSthhmo5J4BeYiKQZUMaa7BsoyuMadupolJg4lFOafJqPLlwMHpi1Meo7ndRw
gndc77T7W5RhbM0bS/llBRW3NvnnuQK91+1Tvi6+dbCbbEdjystcWN7Z91Elwh8IOPx5MAkI56D3
6AWTDBLANI7I34dmHF5vTUOd8+L0itGFoaQ9+kipB/SN7jkTG0TRKZIK/5PGpmng+ofe67NYz8Ig
VfbHNJvaBf/7xnjKPTJ8DKKnjVxZvwb/k9BRF5rCjfhIYG2bCAlg3z/rf6PN3xXfXBm8xmgl02z7
/b0NoGYtV4SIpUr8PZn3vrA51as7e+F0LAntytT5PL9PDZuy0EImseAeZXGgetdqhB1hsIU9eK/s
0D2lojrWzbzG+rOTTZAuw7cRxCsZJhOGFtCwJg/r4k0toBPj30BJkviLv2Il9dbYeogLELYFkqxC
E+yTxHRPMzzP72SeXBtoqvkgSZBaCRAop4ZFz0XvB7UhFfMdYEOs50KtcezlurWnFZ04aqrLDkqu
l2cZUh9ew0Okfy7cngRE396BGsEO0MHQG0PiJyb4Bun/uxPaREJMjYjGGsG9GTrd7RdvBlcDA8Aj
4dJy76TOBIBTqr5APC0WcmWFAOK8JDLHaGxBWUm0sg6pp3FLryp+e5NF75xhvVRETzn9cXGsVmMr
tn+osstgQZmf/7i5WjD3f5i0lzNveZboaX5o7L+0JCwNhJbAfIgBU40tG6aM/LPjhe/Oi6L8QuYK
ZrmZX0jAtj8GD9B9ZG23lkiBmQQP66m96ovZYIXe5kDjD0wjjaHCUtylnXhb6pUodl/a6gP1bxv5
TVvQvbQcyumio9xy20osihwyGy/T6tgtrYw/5Lp6m63uerb3n0rlVPy7iKEHcShv9B9WzxpHt2nQ
VFQX+h/X6pwalvoCd/gN2dFiVG+2zQFO3fZz/UDLPWQDQJjfUY4zJ7u+Z0kn2uueyrocHQmJd1Kb
Ye6y4AkNuaa2FTBt0JaOT3qPOJWtgZpoMNzjNCQYhyAmhrCB1Ajiqavxot650VHR/DkdinsTEXb7
Xsp/SCDGHTsExWkPKP4d70dWGnkLJusctqgqNkkWy7phFrQ7faFbA+CaJeGZAtZ45MPrmqcQuR0G
vd8oMs1lz/9LmLhPrUEN+WY3mAJ46IovUoJauefT4myjBdZS4rFazHocEaSjvlkkBrLXyrpWnesh
VoLIwPae7XR1HRsAfX+ZdyYU3j8WW9NXdHn+Q88YrcekBHOOB0yN8866IsXkjbxzban4KhbWCgdp
pcNzXuezyS3PdVln9EfHxaHPDGnNdARiOWB58uAwH7AJUWXHGmLFxYnaMb9oQOnZNKeSGuV5sWmp
aNCEC9c9RAoYQJS9UhzgKnmat0egozn3IBUZxc/EzBeTXffFuGWMCYQxUGpRDK/Q8DX75a5kIPMJ
T2FkqjMRhXC4u8ceoaYnshrj4IdYDwSQ1TxJzNHTzOjMOrgsk/LKBv33XOD2H/8nwa0c+sylu3f6
Q1nzeVEnTZWt5bF/Mj/P1/a+y/WgHYmE/sBK/OhR3wo4VZOPsaBzk8V7a8LkrRQWfk5fEIDvsIEr
hIQKtMMsI+R5NXgAg7JHsYFAFcen/lJW/ZCEAHwdp3q9K3tK6eAVq4a7auv4fOiO6EUG/3Pohfjz
BQSkaE+N0GRGL6A9MbUqWsFFQ8/k3fvQNH1EoTYM3ZE8h+ZeDxp3/pnPd0yN/HEG9P8t+SDun6DB
OTUPBmRtH1z2BA9ggT1XtYvV3gDNG2xD6apAD4VVuRGVxvNJronvaUpWjhLaH8z2xQzYyBSI0Xit
i4OpAgKkirhJGYButYwNIZJ342g2Jbbxp/Fatk0sdUuhBZPNZCKVJAQzmoOOxpQb0zKAblke88IY
KVjJAdWWYLuOs1+8jW42gmOtY7P2jVndRKDc1S7ycQg6XrEC8PY7v9SCmVo5O/z/FTteCRaNt6J3
Xc9mwppYgZOd+Dp57duy4pqwOUgao8P1UuOCOm/NB2l2F4XrrrWkfD+IiMLHRH03ehO+vjzaMrfs
UnM2sADuKUyDaz0OsSxnq8Sfsx663EVDIRzS7Br0oG7ZNAuAjk5fsy9uSE2BijrkjC1Z3lno5NPV
uS8/A+J/OXx9u85lsgSpTW78BHLd/66jcp+Zk0zVyy/RmHsPWxXnaAnd2YBn0CZc931FrISFiBrS
Kd+wOcK4no53vy9p4NNNDzTXbGuUulZk3LJC/jU/NQ430ZMv047YSVfbKimFzPQOdgjsiFV92i1q
HNtzirhtHPBf5+UmwyrHeER8KTC23x/UxBqwDDpK3sJJ7UXqTLDP5uHzPOH5C2Uk7srrNA64RU5x
8liIz4xiSSdpGuauVt6uHeLMPwWuWi7FpLXLjccOsaZQnubVsXHFbMwkHblEpeTiATUycTJqIc8O
SX7dCdTl0jZqWkzEoogxqgzHIOn6nJuBnC6R2/IxV4kw0qufnMLUfTy2H/UTIBmiubs1s73HOfzq
iZBu71KGgwJYn4rNnO5GAs6K0xINPIfYM/KT4+h8T3OiTJbTyQdpukZjy4lXqddL1xj7aYfYRK6R
ZOjEtrTSWOLcQtKoZaSpwxEfNfeJ/0+EL7k13bnOO1JE+uhz3r3rztVtbT5DLM9JHmeUWLl6tFD4
hyl82qewoNj6dL6dMDs8Dg4ugI/wWSFmy4Ll0jSlt8J1JwesLwqdnR/aSNBWjFiZ80oxpPQFPihw
pD7PaoUzC7Ns6wuR3qYx/7EQVuhccxmEFqZknk6fgUTIfCzAePHXaWBOC9IDcWgRVMJ/VON5s/uK
dWiML2iQmDc5QftsyYmpSHGButpLAwgsUS0PnO0AUbjQ592bNJ107nEgvj6qs4iKk8/wtnWheZpu
ppmAJP7Ao+qaA7fPzGqxQP8yEiGMl0insC73klBY5uCK1l20TMxZY2ppady5atwOQR1c32L30OYz
TkfC5FOc0Jsu/rFbKOIMvK6NYfV2nnes6pwubycRW1xn6uT2szdstE5OUKQc5EzLMhBXwgpFCvxu
1v1tAymeQpQJHgBEDlcIiKaL6lh1i1vIOg2oqnvNeGJv8JMPCm7zFR5FnfR7MAmd2K1zzxA8O6sT
Cgx7p0A2t5BJjOjmi5tpFeSWPD4NM4skZEtZmi03hM+8gBs6IYaO5A/Z1+0GrOuNir89//eHPK38
QQ8hVsuip2V3yZmbRxtWMAufi0+BqsKyf/VjwpNlJMVLmnoOpo5c0fkZeFjKnjY9u5kkoq+DLQEv
jqxUhPryro8dQInPdK4JfkVVyogcbEpYVptznpYcjUJvdUkiQ+SP1iqzbhYturXiueBdxqNTvNE4
yWDUhWrKA4iA2n/wEvPmo02reKCoF99c1BV1uWT+bBKxTNH00XvbAG0sSsU/7PI7ev515re+Ddhj
Ubk8ykPWZD+Uydg+RfVgQQwzhwRsDQ/NT/49NyP//P8mVU0VpkbCQ3RYJWFN3A34t/c2bGK3d9eX
3y4XMXltLBSGfmGc02KnbFlAeJvQqBlzO5mI4g0GZbtePjrQy+IjiJh2DH46X/qMlrMSmz63+Dpq
bHkjT1cJteCV+JKm62B85fj3doGQMmeY4pTkcoV8k92vWR5gQimzCdu3V5Fk+AJrXxb4zEkPZTwl
k/Gtvk5ynRJ3RzIY7Ack5nscQ2ThQvdGIMRuR6Dop0bPH2yo9AfvlCrg1/zsi3oh7X0R5hp5JsSM
zBqxIVS+Gh0E2juGpgU3St1uKZhWzqTtCtf6pUcTHBXnXjtouyXz1sc3RXxUg5hxqzeop05521TE
HntjvSv+dwiYvGFlIOrropKH8REB4MHTSxQYWK1jvAOSY9HB8xihNikj7h4LHSQXeC4e/GzN1tkv
RHqVzIkU0/WsabZ0U97YodY+J13Gyod7N47rwYhDZHOnCpdzuO/AhiLQDdskuhix1exSm1I3A6PN
qPZuhetYDzt4mOnaNAU1NoXgmHhsdWxu16y3NX6EweORHCVLOa7baZ0xcG2hW16TgGGfB661F5XM
KaqT+hwUQsMywC0rIUE+n1gakEawDGmd30Z2wrK8OjlVntWiWw8WGP9l5aOICK02dHod+lPRpL/k
ayFkyyRpfuFeIOKBwX3SFvA4yhV4RpP0/mFUbjYwVHWmLZ7BRNMdl4APkUAnjAwDtkb4efjDbuOh
A8oq1lEUtpyBo4gsdJn4wLHlDVr8iFU4uFB5OkJJsSZ72URwpBPd15DNVRZby0STX3zScwCRctSS
ua+ffhwKnE0HxCaFrqxhZoF1k8HcmCrOWOWvCVhPO+90VIfjzdvfEuKczK5aML51qpfCGu52xatl
oioPYaTyU7+Q8kgmr1A6Epx6VjxcohzFAr5uSDzPz/HP6/r+yeIGjoDWhuJVNg+DCNyWm6qD6n4z
19JNRqjXnWGPrgKq/dTug9Tnb8u+4tF6oug1MNPzTDjR/hkzJARhhZ4ov7E+dozrLD8nSHHMqnw4
7laO0lOVqKCyHZGaQHmEBFerFeqPNCKjO7TjUuwnOktkezycHYOO16nAIHhJ2zOAiplzz28zQgN5
CIgeiB+28RFN7lFdy/plWKbh6/KWqcHZSViX1UQmhqK0WSjvP0mFwztq3rmv7cgk/7R5ZqtgMZ7/
AhRnO0oPf8pf5PUQ3yHDl7iDiiSU/mqFivozTiXj8d9UM1obrjW5HO4CHk4EJfevOFnx3fLAhjrG
nry+Dcq/uMpZ2gOtzwzWl/szfKNp9T/Q2d1FyLV0KG02arrNGrIW7DH8+3DBqEeBFdXZot1exVbQ
1Ws+AFz9hSUz6+aWDIElSUfombgbpwBjjyMR9yEWJYH/VHX9dcTMtbO002dPgUorNLLGwzyFg7xy
CeNDx5XbT54mSzBCsq1k8LeQz6aTVnj0g5t9/iEPeYYA/SF6r8gO+rkJHu3K3LyWpFNAiN87UK9M
IDYZRB9U+zSev/KjgMyHwlTgvsNvh2wHL4puQRgpQlSMq5cb8MMlzB6WUX5pMgAbBpSyy2TWek5j
UILHhv/gxtgk4wATw0Z7XWCHDGqskRn0tsV3UTQJ/9yTzVpx6uJWlFTO/LRUVfWXh7/SHAHt/jM5
7u2Qy6H86ebPAxj1hYHYjoZPnmSEzXY1z8RDjNv4Uo8utdMVNoohOaR1SjVstOPR0gjRS6EKs5jc
IMRdSJ3NIv4AjfSYpguDGnMomDqLLZmxGsEno38aWjSBgbeYnlMw/DfstTTo8P030H53F6/DMxk4
XQ+qRC/GwyqjSW3/tawqYY1O2sqQpSsednSRYlfOlPz4zZxVU4iHl5zojR6M3Wc0aP32wLvj15nz
n7sE2NHl8vDI+jDFTJqWkgSpA6j2wWH4VORphIRuvn8t07E6+LaWY2x4EJ6hcZsCMoOhgdl8oeQb
XhE3boMOxDOYiG5qOxWPx99JuagR6LHw8msiSC07kTN3NcJ4r8j5Fg/MfFPkIes6E5kASJR7mANM
KFiiwI3DoO0S2BzLbDtiIxX/x0oRUGQy7PS6mvAKOd2tiDIanvFyU6ZpXUh1k91j5s6NiLp6KVED
9bpzkLQuuPnN1L1d2ZCq1m38AzILy5add1AgdC0H9jHFhSdprSj9BSnc5Cu50SJkUiAHgPOuXg6U
+TvK1XQHRfM5XLTEQNbk0hpV8rI5wOjXoWDRYYs8/bVNvGqbTqgA1RNkxzr0IoTY4dwgMKZVrDDG
1kO4O6dqMjT6x9xSuz8seHxAU7QR9cpwZjmtfL4MmruEs/DAUQrxZi0jGvCAr1HG/ZAUWwxGo8pE
2veYl0QDWhGl//EDcbxgUjii8jUSqh6lhUdZGWXlwRt65uZ4hb4UWdFdaCusuu8orP7Bcv7DmMSD
+7kKN4WPtalrjI7iBzakwsdf6o7mnqXjCa1SCYx9ltsfBxiF+a+4B9cXs6E52zvMdPay3oxHKhKM
HPtHK3l6PYRjnM0xHDJISxFMudS2T+A7E1Z19s1yH+pgfbQ/Ndf67ppfwyJ2y6xwNZT8poqHUrlr
DShNKslJeFlR/gZe5/27/lX/m5OFGaQxyoiV03QLGQJGQj9Em96v7ceLk+aXJ/RsrvRs4pIONaAD
Q7X9dS08JB4X9Oyuxm60kLWcuw9KLj+fA30roPlk3orjIDQefgKxDfpY3BTOPVxQGKWZqUs716AA
gYWf2OWqPvZoFKhV/kZsomMMKdHCpXfhuTHdhuVpKw3QQc1+ZWj3m99anNu/eODlxGYNn8lMvyn2
99dRRR0xZjlH0uvug7FOeZwXvLQPUUrQvZWwSWqpm0TABH3oZNf5JbK36Rk2qtH28DMcKprAEV7G
NBxhP9QlR76+uAgSRC9pb4SfJubXo2CKCkoMRJuZlA25yjM4fDxw/d9mcNNPye0RlvoMpWBzz5qi
e63d7d1rgOlvEDIczMP+68S6u3nepPk8jP+UrWjVvNr/CvDuj2sZy23sXoIBUoSFkfoPMQ6v7Sd9
ZDV7hxXstSbZmKh86SGpoF07bNQTQ+k/49na/HK8HRpnte8CHfLYedUS5vkBLvUyIzjgNCJNTmdP
wZlHP+wxMRQrh5wyCC0yew89G0eS5MyHrdw3iQxnlEGL9PFpfj1HSmkDQt1FJ8JagE7Ck2mxNfS0
GTLQPUMQRmXPW4uoVwCXlu8RwkkU3x3CS8PBA6d4RGYTfEy8wbT70auL6BZ6oMY/LR7HPwA3JCPp
cXCdkdUYEFouG04sqWQW6cJ2ungc8I9YaddzPA1F5TJx6R31NAJTLcE/oSyTjXoTFblfORkHhZZa
q3/kEK1i5lehxBBl9fe5GojiQW5LLl+kOkbuJtB3DfwyZ2TYdgTxFAWB1zPfHlCKg+/XgM5MUdGf
RwA05GlJc7j4IQlfyQaRCUfE1BTxaanawidKEkRX02F7mh5wfsFZ0ihQr2u59FZSj4nPouLM9ttE
Fx0ovXeRiJPRx0RzCjcQta0PX1305dBKmvsG8xDPvjH3oR3CWLzKI2zCwgeNcuQdIYTfGglTUSqY
cLDRQW9XiLGtF7Eu026rv8/nnbKPbqzQRRfYfYiZSoBdK9RBzdWNZflJ3aOMvPA9bFiUBEcPbiiG
COICIIJ8MDGbIJ9A1yDWMzsTW4ke1Ywd49jgO+e/JqzHoI1ffB8eRzUY0VZ2qLRUXBqAx8emZBso
ZiluI2cptOyBiCbFPPwMTdtqt32hmZRxoz2T5AOsLYQ0d6NVxeCGYaVW6L1U37rtsfpksruscg6G
SDb44u6+e5SRe5ryJ6AQpV/QMzhTrbugX2002hJYG0DiELvQ6TIQvTRXrAoev58Jo7YETU/f7Nt0
WRu+TjoN9K67WlhIrmb8f5o1FV+PJ5+zMDgtYvNguWCx578F944rb52atz/xpkLbJNoDQasfT2K+
8vdo3v5WNShTbS+ZojH4U1qKwRZIT11vXQRn8FClEt6EMeOx9UY/C2HIfREqaEoE5ngDDF8wp4uY
dLoNZC396mYZZIDt4JabM7KGaaLtvCbYGP68hpeEDq03VSKSMttZjM6MGNjC7tyHNvm3GCJtYtWH
RdK71KlHCBU6f1dX8Kqhr7eK+5FK1GGf2fOivCrdLlH9CaRgM2NVfT7ISN3cBjwQaZMkYqRsyvft
j9qs3mG0A8FD2Fwp6SQn2n0s0whE8lgrJpyWbKSfvcs49GmoZfZHBtXNNDHn5k3nFadfrJpLP7PT
HRdzbrp36043TuujwdHX0XCbRWS2o4TEMquTSeOSMPYdtu+Vvn6QcE5MhjbSTTApDv+Msa/S0QTc
Go6D2k0sk1iatLAwaLGGCST+lJDPxXmIX0odEEkPJP7Mn66yOWwiSpoh0oZEb5VXCqjQPbfes0Zv
OPmdl/DmSgRtnXV33tt7LBlYHYO2238SD5RWOpdDiJVuycyCAc1x6zit5IWHP88IetAiUBtqcojO
nZ5qTg9Y05cKkIehB1IQZ7WuQVSEg0OgONVBNl9uLjnVrz8wEhKG21KFroNOb5CJkboZBsG1FHnU
x5+K3vx++4IuEMAhxhophzT4YEx9z22s3wCdyDhHRRv+7hCU1eQjW38VWDFcQ+0IKT63HwKgte/6
UPN2rQwncEJ56TI8BGkhrhSc65/pAzHeUygGFGJ+Xn3gMzD7z1PBkVqz0iSjfIcRx0zZdYEaZ7sf
QS8kA2x+XqyYWDgG5aB1hIkzf518ze2GdzpBFjSNsTQOMDnfkABlT1G7HOTWgL7OHSsDgIb6xTu0
Us+ha0Jq4P9tJJLUYphrsFf9WUyQrgv73kCP6oWKlc+vxN9ZF4J2tj518Uwz2CCL748B/EHpydbg
WtBS/aIOYWTU2pvZZKmQjCCv7+MgUduUyXWzyU2SR1L9iWNepRDLJ48fGiNF0/Kj6jXvWcjT6M4h
x6wf+Q5Q5ekJOp83MG8cwTQoDsrjgu7TkhK9uaLHvCKd70BGwOD/2YStS49NN++0rBekyIPF0wBh
pCO4BTGMKK4amxYZ/YXbNddOZdcnwVNjMyFk2Z7icYsjZz+fCuXfpN/X6fsLEPP6O3cxDd0gEfTF
j8+8SA+7NFYayEJ7YhmNxk01Zj9HbeqJ5Buq9VQYAEGYoK5E7Nb1gkipOlpAuw3UFPIi1cKiozyn
VKCPVaBHOfeqL1LaN4YO+mEzPDpkMwNNC92yfINK9Y8g5twUM4lNqhqgTKaoUcaeye6riXS3+Ibi
8pb22ML5oX4vcLJnHpV89zoQsOfWzX+kn3l+s676TDz5uh3AC0ploaNhltMRgB8YWXT6V+cTP+mJ
WPU5qedgCG/BHMuRlvs5uI51hjouHp7yvyKCVhxe+UdtyZXvRkUUcqp0D8WpYPNY11YfoSgeyraJ
tucw2EA57SMh0RX24xdHGwfIMB9pFyzD51xFiuLzapj+PlStvnu6KoPK67P+RxjcbeKALW06XO/g
an4NyBfu5rBQnstIAwSrWrOjN+FGUNvPG3uKAaWzecrIxRK+Ukzp/kRDh56B7KWLeLFQIKWaYXdl
r/wkd5M0qBy6pa6A/GVOz5NbiZdb+6e9HCw9KuPBZEC8fILGNusJIhKXQf6tAZ1t6Z0MH6AkjMj8
+9Rxbewb/iPZCx9GYmd6yryzDJqgpdWx2AOM8EnMcNhUnrPtr0aUUHgpj2z4+IYFR+/pOvPpO1FH
zbNXZMmIiyXixnUI8Pydo9mcS9FBlsfMEm84G4klFxGq575zAr7fvHduw5ZACEHm60Md4Os7WK2R
WowRkWhWRVNRMrNNj5RNtC6CflHzMvBgVmfdHtUqftlUNUBDQdGKw7ubopNanLaq9/PqO7S3obud
jNXZI4z8jSAwUJL8Dd5zFNEN9BuaX40bpdOmg67u7bjNkH1UqrbEw0Ups2O+PHfypmNsmPem7on9
ZyGQCRmI/5e8lAkblJA0SEXrFqVAxqEJ3FYrxjj9Pya4Ol7am+B9mcCz0oKCQiqoYqvjQwRwWZAe
Zkmhhn5axYgtkkiBFm87DZDIEv0v2u2vnGTpJde1OuIHrjXP8Ozx7nklhrLpxMnoEnivMW2x4e/K
0quTdAEDtRQ+pWrL+37fqQ2OLr1CiVUcnXAmCtV1TmKqqLkdP3s1jMBbTpLPxfgYESzc1Ea3BLEG
bnXAafiM4l/T0/plvHc2oId4FW5vX/D12/KpcUAAMbFCeDfQf7SMGO9zHd0B/sILbqsQIK7vxOaK
ggNItQWQ2bEMhDJ9oeGqIQe/wLn05ThOLDKwJp0Q/tAMKiMjz9TITIUbbA5143jYiRUx8Vt+dKmG
1+NPvuXhQL1LFF2lZYJp7BO3fM1Lb2t0czRCnH+hMpbjbbDg0Ve6/TAfB7yQEuWz8v1ID6Wgtdnd
aDM/QKg4euYIKYRG8aP5D47nUJiSRcikHEaUx4Kt8OXccgveFtd47ECNRgqkg3nIRtIC+SZROXBs
V6UduXWIeWkMTxSub+PNR/2APEYWRthRzmtCHCizgyiipNG2jUzcW/P3NPRA+jBqe1hBkpHVSFNk
gyl2/ds/LQ+50/E88BdkHEo6lWbqCSYczVk5R3huPcGJhQfZgLAb075AOxMZxGuVAE5S4IDcoyh1
VBx+2i1XDG/XbBzSy+C6jth9iLxKFb8i0ZsUkJbpLbgduM/xe8HhfJ/lS19hhw+zidvdTxJDCawc
wTv9tANTFazYVKwG+VSzB3ahHGlRzEXSGjfBJougTe7ycyYKqZjdfEv3iIDKzMV59fQNgFlQiXch
VB19aeRxPOWJXA3d/VTjLtphzapTNuW3en98N80j4eTFEW83bolerwGEnuv2Ioaxm9R+5dRDdE3g
jVmx81pWVJ1siBIQO4yxrNt4yeCfIpb4LXmTnIYZ+3/mx94a2BYlilXdpwRZHB3TZnDVRC/bvkQ4
OlD7uzqqxzQv5CyVgTZiSTNNzPerymeN5rSWPU6PkUebo1DzkqRhWQntv0dT9BdkYRVlxVYy5yox
Guk2bfMoyovAT869HMI9P+1OiJ29kTtmyBuLGwKjACneoaxERnB9q7mYfcFyD8maRwpiHQxg/cYj
9XSAwxEAuzjTO/gJhf74gpVZRWnf+eZNRDu27pX71KIP6/ZMFUjiNKnVVp90H81oq7jAsHm35aBy
2CWNcGesBJOaQzGkPRggl0qCgNQ8S6bXJSQnOm57/nCV96xXEfDg6uyTzXgi7lS4SbV5eVBppoAU
6yX1WEMd8JalU9yrdrEEHv0zUDDHgbub4wK6BQHA35d8x7iPNOWlZZGDLABUb7jVPC72WGV49nrw
o27HnNkeJceRhaZmsH1gHvuJuHCJsGECbwq7uxuBupQxcCHBoVuP7syKdO5DLAnTqmWeGwsinh+l
YN/riUsXWfNNiYJTnI7nXhCVWVL+Q4FHSW74Rnttmmy+7ae5DiDAYgJn00b2fyxF6/6iao4+vxz/
2iIZWIi4sGXFZgfqgfxQP5azbyq7VvZydldn0hC/C/A8JvdDdZbeTj/dOJEtXKSaRA7jBNV3nFnQ
rfd1HywpQZ4Iw5l+miADiv3cTThS2y8PbzMRiq95Ytk4IkIlPn2j+AMeAduI/nMWI3HrrUe0Xg5A
3V9kKbLulhKurFMYIlQ1Y9oxj9MpXvgbNO3RrVOh58vkhWSr3ojCRg5Js+ZydaNUorUJaoGP811/
EzXMtMzgh+bcQyPrK8icyb/bucpSazGihhPvXbo92rbpyOdDUw7LS3CDpgdGUZnquIvNXrdO8hoK
ZN5O//hkd9GQpdLQc7iGcmqkJRBi3ZudCjWEUjWNo9pQS58eryjvstWnLQkImcEyYts2bmHzHJKx
twr2ZWCWgy4nfjA+j8/9U2ahaKq3F1+TZuWlaFAArB9SIwNCaKqtxhpHh8dtMJp0iyNsnadEd0Pz
i04FWIh6K8qH2ILgIYgfl5Kehl+hxEKS6eHLYbEM2MWlCOnNPoGol0jeYpTxMkyws73VDtOeK6ei
Uaj6Drm9IrTbzdM7NGk3OWYDJcPrzxnSbbttiw2fXl89Aa6CZ4lymh+snl0egMrRYWKWgP2lYL4E
PZAkZrVNoEqznhfl2jksYefpfH1KvovWTi60sJvqshkiP/pEFsVGogjDpHM2+wNkJrg7Eyr1FuhP
2YwA4UKVIYA5q8DcjaXwmG33o14/05ycjEtJgwmoiPfmthmPq0OxIe5sAzVUzZgJkplQy6659kbb
t/SlgPNt3aYBANkOQhAE0EmvNFl0KY0M75YFLDQRARVoSa/h4mnjPFLOydD9doJ7VzGqi/o7Pxkm
8iUltbAR+PD8twJ8GX1QNsRZUgEj4mcki8mGFi7WuSK3eksgzibIkjc7Sr7QRr6t480jHN/50/U0
+dcCJ33I4IRYIcpo+IhqwJSE318tu3AWn3AJeHUwzLg6Rd/HEg4tX7MTkyDUcyagODSyAg8vk58Y
+qh1NXOgh9cur9lqLoEZwx0+qDNacG4LZ5o1ha3hXPqSVFBUNa5iC8XJ6+wg+7CFH+6ljcqQczyD
KO51sXEeYByhKlebWnTfdOD4OtJtVu0kMwvEcYL6EMukDpl3utHzfuW3exMGZHVDmjFf66kw9biP
BJBWcu8/DZmaiTChyNcusKyU9QwgqCLpcmh56n9XglG0ydpZt+6D+gaoKBfHbm3pNbp2oASC0dNl
lQIBjFpzoYzQvHVUG+54x1sxLjW6ITAoyS5RAKRVQKMnRVQwrjzLs/dC7rWigvFEnD6MVzKRnmoq
9qvlkff8BGOVGCNlyKT4v+ISw+Cp1EdILd9erPtZ4VeKGHAmbKRHHaJCCYunqiA6+PZksWHzcTdO
95naEzOWi+IKNAFnGxUFIfK/U7x11t0v0zBH3n6bjEY1n6Znbfmpa/ORU3wGj7TXbr6t+YHXS5wK
RnTAIVZSrqQvVciHdKNzCgMfIqXePrUUx0maywDqu+kXMKH4bwOs+r9vj1V11G2kopmhnPZr1jrM
JqDF14b/EKU4TBtyE5tCv+HhDAAn8ImAV5Q5WyBTAbyZzsuSQLVSzTpCxgeWEHgXwmuzS5duRsQO
EyZoald47q4echfTwVT3rzej9fcmmaQpv+Kk4dMDAqunQzsuEfq4c9GG7Vkmxwq0Nt9SGhY4jfh6
BibTUgSxsIfqJKb3UPd2HYCZxRUtaVocT9VvDIKDkCGt0dPRhJ8EUQdkKTFuqDkUO3SVBAthLKA2
EvgPk2kMjeVtNdV90fhKE37aejp8sx/Xr3ErpBSrn44tkTjU1j97QGEBHHS/2ikU/W+gbg7I9RsH
g5pwsCWO2PJ+6YyZ/ceQWyUp50M1tKQxRoDcSyioZ/PISypJWCit2/xnCYAwr2AiWvfFGboum5EZ
nObIHvO840c92pq31LljG0ze6rdS4S3xeI7QX83lQrYoZo6UFP2UslQbUNjoALMBQ7Bu/0RyZmVi
6V0cFxNozQOlkIF+6dOO52E0ivNE7Pdeb+NfPQfu5ijRmdRIwvFnxP9jLwHsDv0VexRNkCifBtEh
qr/gTqX4uOdPGNcTMvmnL0VNGNHK7mpQ+c9OXWCUcF2nHhrobtmYFFqsFHOVMRlocarWF/eLCfCh
NPUmF878ozIKxHK3sf2mztMpZ259E6OzJuh5GtRQXKgxcrlPbV4Fjnc5Iq6ESI5/62riZmd5cj5R
2Btvver/Inm9doaU6FmsU9npjRnzuft+iDv6zDvvvFe0N8wK9aXDIRzxDts2DNKMggJ3LL6HpodY
/lDHc0x8gr+mxLY/Ij9oAzZiKLijZj8TcyvrB2J7OjHLp2q0utS4VK3ymWibjosou9+HQ/2hZz21
82ysyHvsOKePSsw35zGt4bSG2AcEOZIR3LEkexg0PtZMi49tZMjHT0+pGH4u/3H09JnQ8qNxM758
Baku7+vu+nyUPa4eY/DSv+P66Wa4JkLccgNJhWp+8oDfPnTd/PgBF1dwiN31leJbuh8kg/gZDoyQ
U1nzf+CxggtK/Kj+0MWOm6N11eZFm5O4FLvuxwGjBGS/wP6BI/vjdiBMV4iEw6DnloPqYUMEF6FC
Bh5iGV+Ka/XxwlkPDkNHtFNb5nRlYf9/ulJFEgVxIKtBwz8oQsQPyRcHG9Wbdq7gpYKnlp4QbN7D
TQZQ5M8iePmHvH7olhnI33Q1Lg/iGEH+GO0iVtFlcI7sNfYT4Szp0VQFTRWFqB7yI2M1hxnVDajh
RzoTS36lzNKbsg5IX2HBlfUQvn5IEVVaCcEkzJ4BCu4tmf0UGdGlyLGEO178Nxgg5oQsdizKh2zR
UhP74GumENh3jSgwg5MnEJKJGxees/cZN0mUpX7qPYUvqO5YwRzFQauqoUq/Bn7JoM0f8HZLq/rq
R04KYMporeCyse6BAsa2qwNaUrshXcQbuYRwRRGPaqAhtJX7GM4wxNYIdVGHpMZHXkCFcbZrW+V4
xxBDT+HhKPUlbFv/c3o+hvXHZ7569P+5JiPxS7H33NGllvgzfXivaruVzZzyzW06LFS6hMWR0hKY
pRZ+8EAhWBP1M4IFQI+GqPaVdJ2uiug3tVQ+oUbgCeugEXZKNo6+K+rh63AX7thUOXgjfIPY7KOm
yZXzqONkA130gk2vXusBPUeFnl5QKWTxOclU/TKLWo9iBf2r5JT3PH12mqZZof8yAZvnnEQdhFYy
3pUNaH6Fo647zS5TlkUea8QiECacVEAMjSszX3B0gFmywZQMdjugwRpc7Lm3hllIe1hvZmAZutW1
0MC9H1nJyN5kp9olbZ8aXso97c2kKvwKISbFLpiJJuGwVZdiNywxsS2FpfvQpJ+Uc6rkeJ9oho6H
1ldlDnb4dcAUtuWFxFc5vobGJxLc+KlbK2Q4Ve/Lwq6l73Cl3oaQ7UtZyBlMj5CKQ/YYntBHlvuC
qbHwH0AY2Fg2JHJBqG2Y/CFkyBlEIIwvcgQDyYp/aEuSQTs3NtPaCVWyoHs1sNnZvp6qoluh5205
uqjozkJo9QlWQPEJKLMK1Gzt8pKUrO9azIgV6HHzrq0dV4tKzV7jhT8/1NT5SK78yQXTs5Nx8y70
ugH/1Ssk9B+GRn+f6D4XK7dMkqDwSdW1lh38+ZHyOjLwX2ydKNXKW4mjEyvPELqXg+4IWjQAnjik
WPErJEf1JjIAYreseONdRYdAJbH5TQR58Tw7yQNf1/pdDZiaZREebsbj+WqL2ZpzURo4P96SGwDt
DU3zTm5fkGtDmZj+FGShYmRqfOwm6QfNfk7ePveNOXGWiCXCUW5dX61ESVf0+DHlIe3u5LA1Umqa
EfSSqKydDmLS9l0AS/iLHMGoVRsaUEBxjivPiAUF14s4ONMpFJlUjH1fwJx+5DgEgi4EXH25Lzr7
Td1FzB7/S8J6TXwS/pO9ACLZhxvo/kQZRVimRdqtaNBGoHGWmosIG4xJi0lojWK7VawppSFE4ZHh
xzkaJldclGqgOOQ3yL9vJBne9D57731SrVuErIVJY0tJGKsWi3ZAW5SWP+o+vfKwX5mortLakPmg
BAgGL97JUmGGRrkKLfqAnZQmWwAr2OJJZ8/q0NTSgpTgNxJI9GzElgCGa9HjIxMc1pcwKYdKvoVt
JG65q/tjFwCLBGJpB2KbrxXXhIJxHw1jWds/QkYg1PpgILUunj3ywqFtvlROXB8fsMEbn7XoLU6M
Qp8rfX28I7R3WNgVdkk/rovMYUPke26Pvi6thzzIZsfLu6BTTByY9fLA6M7md+CumWmvU0G3z3bX
zgDPG8VNmhRSPTkkfqOU984EnARgFrcOCuJ3aSp3dKH1JSdhG1uqYDJ0MRTL/kyXB2xfxtOsJsJd
1NtCdREorp5NIFQbYsqi8Q8NYwvrhrKbkl5wYJjtEOCnskN4QA6kaw1xpYJ1tq/kCFeodsefdM8v
g8/8u/5SI+Soyju3pLM6EreS/5ZuTCW9FG4G9dLo7nQMQW5hIZs8QG1n6azn2Vx6/Hb0V05pQ7FC
TN44GtDUpavZ8Rpg6DY7g/RHr8LL+RUFyfx1oyElP6Hdc47TvpZLiZ/36wWEgbpwoPUkcvX0Un37
MlysPPpxnIa7+0Q2YD/VNG4fZNWH793E5xkGWQraC4YxXwBULAIvywkHGfcGp8bKR6im/mUbrU0y
WmuNs8MWmfw2ORfHLYi8qCcojnV2f5wCTFyKanQ8OBXA89r9pWrPT1bNBtPw9elzhsf9bOQ53k64
SEZb+uJ1Ui40qQ3mNL8xM2arZiNIc6BZYZwF+5FiX2PF+XImZucAFp67uKoZli8PU7fm4wKwtKAS
MfCeDLv2ucRdwm6kYv+/G7YI0asv8r4eIvYE5ui3tguF96JDjkFXFV3zIS5j+wPpTgO5yhX9LtfP
4oBhNkqvy48M5JbMAaJM1hC6s2pK4MhufVu8AIWtXvpK2W61EZU1far39ZEAN6L8yijVn7x+wGiW
sVThyv1p+oVJl1T8f2UZJlv3OENykqJvBF98K32NekCYbsAeTuz9bId+yofQZ9vB6af8lRmA2m8T
Mck2Eg4iADvbZUE7sWGutQT7QX7W6X2zH0A321JMGmqEWLkI2XQ+9I/grAl0IT7bNu4ufq2ak8xj
rhgJDvmVfVzh/cPSyUCT8Q2VJOp6rLy7yqtCIHWoYjQTAl0O6GpmUS2QHTruRRgojNG+t6QQGRSR
2/M34g60bBAJLpZcH9liyc+Pp9mBGlKJP/drSPQ56avcvJ7/jSwqLCjPzCoNCSFVX7x5EkpAIEbM
BiVGo0FUO7YBqQfh+KivLAGxIO0WGwzRGMlFAyQgKBJtOpdSNJCWPa7wa6eMafFBmF5wRARUt9ZL
NCL9daxRxHyFbU16fWnzhQHNQazMkQGdic+K9u2rFEVvVAaJrnoETE0kUTmIa3Nja51VwnMLAqkm
xSLwGqCbp9e9pVXWHEIg5UF9GGSJSoAMArIIhQot2OfcIn5Pk9PTz87jCCFfJm4lMpgZ/q1BC+DV
DKNd+QGymyekUCXS7Pdc8R4AcngHw5UVrCjXMyOKvtQM74lJBskSfrgnTrmi3LxOvLbGEDE3xqUE
eENV0h7ZJYbsO5NSJy0gkEzolwbU9hzuQ4boLwtyc8AWBV6tQtbSd8eIGRlmwSW397CoJj2r34Cx
Ix0a3UaaeSAQwtVwFkLLKEx5eLovQtLOAn7HdfSWA76LjEcltTiy94nbuhUVMGKI1jtiNpwmz79V
17U6aFyp0YZSV9RQqp6dg0s56cHATLMRBFgtdrSGuNDjsSzPd/wHhUk9G++TpwFdOXMXWdTH20VC
qvGn0KYT/3RVGDyHepyUViswPhE80pCO6w2lCFpJjQyqn3GQITrwvMvLz77zyTjC4AXOuBroRuJi
UJFy2VQDqF78u+Om9f+5fT1R2KYjDcyNwpYU0JRj1EFrwGBlOBcTnmoMn75AbynfEuDCwDes/vIu
gjVeZUCAQyEV+GAqnfa3KqbEYLhWnMHE5z3rViHqpyk6haMDtiCCsew7vIgG5g4jlOsdV0j+j5VK
nu1dsBG3XbtgV5qKqsYy/5DxMF9+cFomAeR/e3ecQUzYm39WCzHJwofoXOeDDk1/G6hWelkacLRP
7tndg/XiAR7HNOS6JwVNnMieQcxKu7iGRgR9JfMS2XNksghXZ/tCO03deTWBFA0n7H1UOaSnCCGh
c3wK0Ndqp8ny+VzwF/O+CZ4ER6S90zLFgQr7d/FdJuaiuI69nnsQKyKrSWYjp9yY2NECaiaitI59
PJk7+482TGA43yuZE3bLICDIieVfKEpV4vz+/JuxrZzZ72MNK+LX4uALjViey7z7rE98WH4nZl4w
HEWF3nqk8MNghQpgmnGhZGfHVsOIdntMEkpQggsPtd4BSSgWr/qwgKM1p4L0XBctozV73qOLDcku
XsXVnGu0P4NZrop5Q2nviWeFPqK4Aq6Knc9BORaCPXw6RvAT4KK4VFCwj9w7hRT3OKjGJF8BNmGZ
vgnM0gTSaQkW+oTdQio12WwTpZGoMbgojtUXnoxd4N7H0MJVl8/Gf5LqdNKXOxUSLUlpXox88pLS
LWjDxb+hwPVs7uI7jKdvndbV5enOe/SU7nNgWw4pPLmOkZKaha4VCazBFG8AGWfaUEEDPTZ6Qw9m
9Qm3T5sTXlrE0SY7p6iEifoedbSQEQ4XcVAvaAztAcFrmlZ+59VYXoxFufBEn1TRDa/ABJPN7Vyw
b543pUlf3MVyfJf2G0Xyu4ld7oOucjsNjZGWS2ups46uasBViLZplxKYEcp9DYyWHNrYaK41229e
MzXrbhcTd6/8VmLJy2/pdGC+M5X/pSzCshuYzPmfBZtS6Has8cPLmpL9npPtVuYhlml7cmeitcLE
Rqvg0yPlv72b4DP9aKKuFvoNpSYFHkVgtVlieqQsoSCnV93RQGv8DBEyghJ+qLjA7wFIEWPqyyOx
iPj4cjSe2KDUAXTeppZtsXpoSfVDKgnRdGGGcHH54DVu3ogn6QiHRTePOIk+/0EJuWZ5+4SR203u
XiBXxPzBn8BL9Wihwf4JKDEnFRW3O8go7+ynEt+aJN/A0Ii+fTMAQP/9Aq+ZBCfHu8bgPO0QMWKw
XeYOqd4yhlGe0ab1mECwLfq1ndX9GRiXYHhm7p7v1QZaE12Gmu2tgKjeKTW4g+8nF2xwxAQkp8oI
6qHettNh/WaXug3dK5kGUfPybVCyKSSXmF4NEwis0tp0NB3y5w09euD31hbJogzjgzumNzNST6Y0
gAtxISGWB7M1iDfpgm4d+1poUJkNrhOJ1TB9EUy39O1zm4ePe8zmKBB7YYFq7JgdoLpw8Zt74ioR
uBcMJqqJbbtVWDYF0ckkQio1rP9/L6QC9SKVbzhNKDLvPZRsASe1cf5oHcCRHMs6qA4YWyU5PRNA
bLm2qo53Sf9P8adjP2UU94glUChQ1nlYxuoCemeWupmKtoUbtHQ+gykiKjzz46CNqKZQ03DZwHRT
Iw6PIcD6CMEE/gH8J6CI+3zX8Z2igC0dazrdMF/QikrHSe0UEBvS6aoZCrX0+CgHWDaUZsS6RXsy
4BwRplmQ/yWy5Sr0rWnV8ItD5g6asPMqLlC2b4dQVm/YDtLwdYPgHlfjE5ohdDb/3qslHv3hBv+a
juTz99+SL64JbNnPYNW2BrD7Tfz1ZeCKYoRHSx0ktmcjlHySNx/GUvk6QpavXT5TVND7e3PAll60
ZOlvLKiprA4NEUSyMZ7Dz7uHLY6xtDl20b+dSvUgaroy/k+TgZlsSUWbLKvkSIa8/bNjAoj9k5pS
CfV6a90o2096p61I42XaaWzsbrjI8Qw8DlX/Rkr3+1GFhXOG5LW9npsVkrATalFir8zc9nEuM3W8
f6GJL9EVOco/lV4jF/LAEPKvhXzT6WLBy+HQXh3W3CGOeQ87riI6UcMh6LdK0b/7f4WTCM6QfJXu
Yuwmzit3CljqNHFRicQhHq1tDK3dN5zf8y4ZWrNiCwuUW7/E7/mTGwhQ7utWtYI+2iLsCTIKuRh7
RPuS1KxslCI2E/r2h69oY+yC/8pLFpjvAv0KGE2oZWt33JZkiQNRhEj+6MODLb7+0fVhCxSZI1n5
Kuhgn8NKmN25lYR5HlD/lyj9ZbpyPGAAn8qF3PsNxe5K5d3pOkJnSoZOLjE3s5MfPTMp+CuUlQAX
fUrqmmcqFPdvdsEU20Krp88ooXHJDucWfjjm+pligKtNtPxZr4aqq408PGNr7idOQWBbHz2OQ2/d
sTkzCEpq/k8ViZYlpQONPP0l+l+VCj09FPmMWuReV/5BSzQ+VE3Tx1GSzD+/EmlaO6Rc6Y8jz/6N
iOnPvCB6yW1wWqVutCasZYA9c3M0JrkAOfdTi6ZiMRfRyN7SCzR6izKs7XR4GxxYmSQSvvwRjEf1
BAJpUjECGNTI1NPJ+dlXp/vpd4jk3Jc1ArMfTE+VWd6+zYYpKyANsJUzFBGiFJDIPczHSVuH3sc0
VyKwM/hOjTp+xGnjR/3MG07UhCWvZww75H0tovoEbiCZKhdKo54jrql3GaAv41SH2wKt8CkSvOzy
cUJrJBz/XmIlAD49JLnaFsBhpVzdFdAntaJ805mrybShOkleFKCVtN4rqAl87dTFRpJqNwiHRIjx
mVmu28Ddc/rRRS6ScYZrnmcR/4vCNp9Xw4LH7k3e7a2UmueSvbY+xRjXIeTxxc95qnpaIOsHjHp2
OjBG+rU9OSDecAeEjkBg7vOXID81ELWk0pzG1gaTxVi7GRjXrjVYCLgimUG4jQrbdGKpmHXBFN0M
Lp8dK9D11cuJMn1S6xoYahq/LVSvwANY2b3xyJdCCyq7SdCjC4mOzcbnxnj7CYpJlBI0pZ4LhbUW
o2KutPYA9r4Ben7eFiOhy1PI+RJZen6IiBnD0lfZ3j0uW5XfBR/s2T7+3qS4phvb8Uw5zj6S9zIN
BEAkxmCCyocVP11WCXWCYd2hY/oZfgSYKwWR44sdtq1dL0SFZ9EQeyewqRc5Gl3YcW1y1B52wW0p
y1Nhtgw0+KYgN+T3O4SINmCVWZOM094RPvd72AUk0f/RVcL/6AVYpk4PS1VAZyft7PefjsGMDBut
9gdUZYrqeFbEGbOiUpb0IZoA26dQNrLsAx9L2lK+E/oeT3rkCPwPETsb7sadAdIs1BHzcyGqIlul
SkaHo4eppmA4spl/4L2E1ajh1B7V85z+6DbhRyzDRj2TFo8B3OEKmcENaB8db67jNHmaa7hZJSvc
UQ0K1Y/LlbC5odXKSgD7mI9a8LboKEY02Bm2jTuNmaYmfP8W0wqqQPHo+MxcwAMUPQC12ClQ2V5y
EteSR+UPs8dPax4S8fwU1GhdmEFfQCdIih1VyXykboeLpaoJ2L2hJzKiA6MmRMBiQiTfxN0l0bb4
OMiOGAJU7wcDKrIVGzQgq/LuNx9qj7VtfNq/Uu9wJq1fSXdlOKodWCobOwO25A2tER5yJfrqQMmm
N8uB5CV0b1F41pm8Fg0IkkwhzbJGgeW8+ZG//KMCbnv/l/78U+4oJtzyZf27CkSNcwzWGxQfiQti
lSxdCcCjhgLQcL4mYq77bICh8L/cPBE0Gl7k4hIIdAvXNPNp/5MubSCYyOwiO8VkaBWObq0hZtXP
6S+ObhusjRs3VNrDVrvoFFE8kibXtH4+KubmHH73XQ8UEXVOlJqUgCIQHsEWKlcCrZKQtVeOt99e
shrvAIOOl+KZv7LeJ4UJdrlKjGPe1AUVlSkkwO6MsUxIwG+h/HeUz0EKFIc3obdFh4FkTWFzP2lN
P+NVWSRzbfojvnDiFZFyUymTTno/4P0TDNu8ARVrBrESZOz0gum8L2zDn4LMHlMAGu69sDCqlJxn
2oo/aroF3uAL5uYBs36R5A8orqNUizIN3OFocckd1Gzb51zeKevzOl1SsSX55bfiC5QAawmk9rre
exgfB3HCyb4GigsA5Pr4L/c7IBhR3m579Ckr9RUBI6p9cH9uZDlZB12fV1j1eQ/AyV1IMtYjZDdN
3A2fvW/+6mD0XlJsm1mjY6EtWmg5HTrZt+lciUZT6doMV2kseApE/aqEtKX4PyXHSiiBkjZf0jxd
6K6Mt2TQ85+AG52fPmlgQ7ZG4j4NQ6FIK2s9bHmahSzBVoAzyvQW/6+f3y0ItTV/KvjFoFyflMsW
2ugGhmsm2ggooJZPD9L2fAxAOxZ877/l750ljBvw65y5nvCVlwPUVZk5Se01yFqB57eQque6hw67
5eZ17WmPMb5mVFA+s7JfY2w01hXdRATqV/q2R566so7Z68RA0ArjiAH5zWA0NxARYr3vKrOrv53k
IsxKpCBmVfHu6RVMH7ssPRzv/q1jRhN6zEDXVqviyvtSDjXaxjlmjGU6CkdWgpSft7GKiIFlOfuC
qkGzHIkktlD+u2c6b9nE7GuKFU7Gxo3WbjY3buaiu0ORyKteMBGNwjJ8CWtaKo/ZHkVkILko9NSz
x99Wxo5+xKkqTzsrORiZAosi+LOQzIjIqYI+L2UfjAc/T3xATaLDQXia0jjg2lfFSwCqt9NEQaJt
1gkMJZw5EdtQFLbTG2WYrWGRunEX7of27Tunz8qtwPuyRH2z8OkevBuQM18oRKifx35ZzLWNop4U
MPlok97EppiXatmSCzLibOv0KamBsmW100Fp07Xq6aA7iRqkHJXXpdSj9YlHiblEAdTHCyzENduB
aBKiwJiEVFsdyjBNQyy+Zxun+NqPhWx+bNvXc+H/N2ABmG7ZBV7J+75aq5BiqhXGhOsXm3yIYO6O
1dsFTjw2MCkbZAJXFUbXdEhuRZ6DLp9V8FlwQQlmNk4P64E0qRq1XoZCO7dcNfKZ+s9MW2RQkSId
DlO/MRxRaEO7yxRFQXQkPPdXiqp77lGQMX7EWGfWCb+Dr0CgT+2MXdzZEwvvj3Oxkjc2MGFHO9AP
qZiR93jZfiHhlgLvN67DotgvJfBUN9mBj+2NjWwHwOgi7KudDeWwipcv/Vv2/yourHz1dAtDvMDi
EuMthdgk7uSLJVLMAYemx02kCNStjbk+OYoEvKB3tLz6rcKfj3k+IKZ8Ck3GqmGPQz73Tq0+Uh/9
wrhbHfjTUpmmJsjmAs0TPTrbjuFdTOilxGHYkOfXDKQtnvILJWANt8k6FoK167tB9z0Ut3/SU8JP
aQrioBmQY9G7nXzD3YGekCtFEQ0l1bpifnVqlj0Tkp9vPOviprzJTWEs6WzE/RqzuYC5H3Gkzi2P
HsmfC8xqcWfDma7vpXTr4WtTXGk8weki/qA7rntSsowPWG0cki+E8z4EsWUndlmJtDOw6Bb/Qc2g
3wuIgm6BfKFKpWyMl8zDeFp28rJIKEQHVskKHm73B3CR3diRe6O5NXOJK9auZ+SX23FVOlEaba0e
si7wMGjoQZWWgKQE9VMLR3o7DB84Tou25kk5wOw1DD+cG5lGj+YnHveOdpF7nhwQOyJ///aFTAJ7
/LJ5YQc0Gv0omftGdHA3vkre/tA3lpN0Lh6BPGITpRuAXPpFFaIi7K/emoI0Hom1naCksxWepgEe
7gT6LsQSCXjG3wpLsunzZOCcGdVwiHSlEDW5j7ONqmLE2bXLqKKSljADllLbrxyGLyzilMS+t4nP
lDT3XIMKM6J8bd5d+o5M+t9moQzZM6235tNFXphJdx2vOZJgqP0XTWbLoU+aiJ67h/fWU9xJPlPk
drXTg9f1lOvUakIgFBCN36D8alHBYlmEwijq7a+9ucR4r8guC9PMfOzVgD1KT2X+CECalCblwvuk
07ZKHOvuhLuViTUYR6stJq7vQcMQFDTHzTlVNK2rZFdmb0yyVeX5xCdMjhZFn4M8l9e6kFbiGOlf
AsnZkeu00bYnH4IscziQA6YySSO7jlEgw2OD/5HSAo5T4ROKA+WLfIqIRph77nepN11iPK//ytlu
1bIC/GW41Dd3I4dPzMii3qK/+O4+b8E/bURfQldL/GSw2vP5+uVZtKUfr3eKM3TYY0mGdY9zoPyj
MRi5uIIq3t++UZmwTCIjx2b1d1MEOgIV+fIGoipF4u9uffMCwrHNFLLyd0lOvfwcqfIOhtNZLO00
nkZD2lPae0SB2EGJah3X5GQtVq/vBJS7HWhkOPwf0Bn83RRweqnt5wl1FsS+jeFB4/1rODCVBiPV
2S86sWdu+nb3FDMsV0hY8pw9SQBnGJzA+8+Y4Iiu8hcZ8EdyBfrctvTz2e/xE5GQj1EYY6rTCFt0
Zd+UzwkxCHvnzqdSS9tirdHNGkKPzq0UtYRRtS3gwTSnpDmOynWyfCcT6mg6D3QpCEYb/rTPiSPb
gkh5vUWlABOLMqchNdQlwIz5ZdSeQoRe6sQoHGHGGrzmgV6nN43/De9KfuSgdEJPN35dpXO54BqX
vuRyI29m3MoTBOkT4jzONS7gQ8QSC45ApUm1YFSs2j9+OjSKVtnr5QsIjhCyhmuySdYlFE8vT8I9
KVqN59PHy/fjArYIXcADijTJunpGqZQN8FBzYn2LFcuCEB5SVWIeXuIITiJ4qtKDkoJPQdf9Uu+X
IAwuFCeMAXe7AUxeyWjjwJ31le+HH6vP68rCdRXKECywvPTqqYBMOXOAW6u/TB/Qy92adEjKwMJ4
NUT4+Me/7BbMqCkV/JunZst2cgiAzKFAk3E5nqbQ/WnBaK5D/08QJLJHfr93cYjhM4VtlWOHgX43
aO/R9FauT/kt1UxFjJX6SN+XtOvKeH9exm6yk5Htu6ft35SyL3Dgv6FybPOBMzg1mTfOBjDiwY1x
0/smq5Dc5NekUa78VgSM+9UBnyhKu8uPjZ0dSZVlCazSJxXQOeWgMTitaGoWYxerV0yptLHjXf6G
fSmNSmJ94FNVQvlOGcTc66pRhTASXs8D2iGMYY3wlHsORUXVp5hUtGW9cw58ssJucauwjptAN9PH
DQ6mtiQVzjomB5w1y15T/8Fh1Vvq9GO8ndQfGFUxCgjY1g/2OGAu/N7q4EYE3J8Ma0LVejLFn9c/
To88V6GOu+ublZlm8L2lUUZHsywG9rV1v3h3FLPOOwnmu4h+8JLJWEOLqXytVSiI92PXAyaOxABN
M8z6V47pv11IgUh34p2Jc88ZVsIH/n03ASHyjZYXG8LzbepAeNIRxid17bZhbRoLrqboOsGcNA55
uB7wBUZo913nqCcGbvmVOgF/hIunKZbZeJEdn5qLM0RMOm9aM+mLNSms0TXlI1207ONsO/QdrqgO
m5IuXzBQmFOO0iOHVAnxTngxmcckKI4awJdZ9mniJX9d6qocgVQT/+0YOEFoZAAnAubBlZoPrula
uaSQd/bSnFc1DB5hMDJpNwplPHBf2OGKCe4PaWbMEmepYqF1l7FJrRNWUklCt2VfDeYgtjCQ3maL
WBUrRoRD8I4lzj8mZAISHFRCbotyq7lLUCAQC0agJWzvW4h0dzWWWavjkG739sIeZUozCO+djogq
7KzIMIoSj5rlTTPUJYouAocFRqMOsOVaJ8cQbI+/RxFbluuGCDj5UyBAWhfiqeunXwu2FBduebwg
/dyB7ETee/ozox5pwwVsgWbDz9DNDRoX2R4NwLuBzi8wk0SBk5BQesrs8XH88ftMZl63nqYk5zSj
kDW4hGSkBjL8zmMQuhrN6+YDWgy33s+C6S9m0IFyidCd1MamBRJloCU+C1vBRgDJEG1PTnivODMR
P+WpwNxn+xjWey01sQ6/ssI4CdC7OOIsO9IsWYyDEZgjY6i6WnLdlwwh3A2H8X8dHBNRdLmTTC4b
WU1EDlAU4DA6uZOHcL+Pzvh9oSnBfaEwyfKBwcXTyCVef0l90QuOr5E6FxKMpjo/eJxihwzpHd8C
OEQ87aet59BmOUsf+M61mCRkmfILkSqmvf2nQqFh0dp9fFGTO50Tqc9duYBreoXT89/DVq08wZIu
ruCA3IEul2v2wgBseaaZrR6g2klpHgscOdzoNtHLd3OA8VbRaza4maRyqI63GUPSh7AGpKG/AOIb
sXfGX+mgVJGOIkt5DKao6qj9hV+LcyZ6S8WgANtwMq2mDGvdmOzx2Z6OtR2NeRvXZ38Y6oL9FZKo
3iPC3eAhIwx/41hj8BK490nT4kBjxv11iN00H2JSSVs8HjWb6xidHqXcMr/8yYHuRwb+MEpAQyPt
ypGT8aECWtbCuwLnwNoMkAL/DN8j2dAIxFDQfbEU52hy1U0Ln0SzHVf7eoZWUJAPyyuA5x7qYnku
VacS17pn4Y7DTd3zqYQXiz5kKTqNI7/FyyJNnizY1kWArVdIne6etiaIC+t1KHY37S6On5c8mium
/2nHJHttcpLVMeLpyLTgTRcV50VOOHd8FVKxu1si6wrpJTA7YC0aDQTHOJE6VoyGh6d2uN3zVvFo
QXVm1MHrOBLgJYNGDNw8SKB9jTUYerjzafCU9RYVoOh09yX/H3jR/StEAQ0kQDs6zeqA8kFc85mS
6w5SdVfcE4HdhtxvZe7dEPYodHm5+PT6llHnvgEKVXDKfccFqz9BMzBkIjbLb66bvb4Ebqc86HBl
utgc6G6wap357ublnpa3U9REHuuFYMWR5zsaUbwz8SJ7kEb1niB7yLbOLgqxXtWj+jkJcRDW9gJo
QW8mR/emrgDkgFG/02XN9lUosWPAtPlv4KWYJ62gvxKh0NPxxCGEUaqHhyL2L6m8VLNNyqYQrhJX
nHoRTwW74I7EXo4h187GJkl4hnty9Xy6FOJZIfsKhXuWYcG4DxEXK09xC9WeWx424WEq+bdLfZ2L
i+fHD0oOC9hsKZLRb7pLUPxv/O9L11qyEd6yP0nzZiN0wtJ/3tw2T5lRaJGNsGlFyQu1b0pgukaa
e5UZuevHOBBk3S0yTAoleYBgpMaDaygZbADEiV4PtM3SRvoioSClJzU2uZJUz05Zlus7QHCTMRdI
W6LOBvsJC9AyFOUmHNYpdffAOQfGvfWnZcep4STUG4NXlw6mfD9oCHbsF+OiL7rkBSVrFiIfnc/J
lMV4NriDXG1yPsgKbLeNDb8Hto8mdIP8BzQkBy8sxmNVxPn8jVeskGSEQVe6LtPjQL/NOg2YNKBL
/ztl8uO9bMSyjAyUDML+rFnxjoPoUPctSod4f2YamIMeCy06faUiSvJXMECVAYlqDe3vp6xqcHu7
t/ZvhF4H2k3fQoGVgM4PUqCJfohAofueeIgm9nwFxHO7kWDROe830T9S0c5ogf2mIcfb2YHpdYUW
Ynx9dux14emSfRU5lR1hHHTj7t8XHdEAdDqbuI3F9OPx9PPVVvo8k76Seran95VkbUu7lrb+Gzoj
y9UMAgrQf89NWuxyPnUzRMKWNe+XYzlzC4bjFIqniw027fwCB3XAFKMhaHS0Cv/ckazYV2+59JTP
aUL145zKNZvzo2Jy0eB/v4Aj+Afgs38dD2B7XAay7NbQzex5GM9P2a3BU1gB/oxydEp5Tw+YyF2r
7Dk/fFNO31S9ApAr4nT9CvMJrRgEn8RbGREdVkwDE6aGjsuoZd1g4XRlMzisJQsiJLZR4iIuZelv
dm31Xx5bHzYhXignVHjWZzXltn4utkcnnsLfXSIuX8+BKZIWzibpOnrVdHR7cjgnhnxtYfSWMQEn
4tePM519v0giqW9x4AUt0CvlemciIuiHXAn9FTjyL7M5U0mxV/rGEUCRL4j6CEe0+7DY6UN7T0x3
8OKg65n8+OKveWfIyzAeKE4hEqb6mYRHyJaLNXT2Gh33646ATtAtzOguwjIFJtl+oAd1gnSAfhPg
cWcb1tyWYDJ07s8SFv/fNr3XxQiYmuxd+SCkZxwLLKJL8y/XURdYn6dT/VPgLGP4bPziM9ApzrAy
IcqIMFeI+Ku6934nFqfyGFIM2nXegYrKWcTw4Nco9uELHofnZEeL8GgCadPobZiDfrrgNndkvA9i
vqVZLPui5lnn8TpPiP7PmPRkwDDG5FtXYfHV6IasCuAiqTbONZir5AEggkNRr6i0pmfwCFg3FdF9
cnP0poXBXzldWSekq9dHE7RkWmTX4TFSwCnKbD6dXi9ZvO5LKkABDZVgxPxhklexxsZmpKwOnXrq
XtkzYY0/ADR6nvyyS8DbE3lE0BTj86zLTOTLOk3BY8gVsBQkDjZoDhTSG9bZNdAJS/p0RKEtg3kz
LrzfiGbvPVr49kPq+/yczMpx0T0tPXjZR0SsOXNIbpVRnV5W1VOarF1V2x5sad6dY4B+drh6wfPE
epr/aVr5IXcTBs+uqgIWAqCxtaQGp97PgJnJGdQTQMnupXKmini8dEDD/Ob1+lsx+RHRCWkCObuk
Ijqe7LE7ThjNlQeOJJX7r5kM9tlO6W1ZvT3xFkkgjMU2ZUqqyjHKHEKb/0UnsbywvivGHX9gqCjQ
4OM4t+ubzs0UOkE8vpc72rIGtup6y2iuFblgH/MjcA4maqzTp0z1XVHw6+ZuwjLUOtz4CsjOhyd4
l/ShEcq/2cwC6qc2DZEL4Dks01UdMVyJpgqv8iM9dZ3vr6Y3sbijmIpChZmWTxRY11+/NnvJnymU
zX62amng1vhlX1+bGeVGzc5Qdb2JTukEKEFe90Ii4jD7+KBLvHa+TPe2tKzgHcA1TXMSJtYomh6J
QkBR0k+h2S26Xsyw9JFGxxZFLiPkaCv6LhWSw48e+ByzURJJIsRxf7SBmFDCJWfS+mk2pBIjguW0
lwx9zBeh4VkbCaz//6yRSRuiXVRIcrdb6eLrLKTH7hcR9WyK0Rr09O4JEGaJcZ310NYEXfoMa/Qh
HXqssbBrZ6+mGqokSdgNRKoQ55WVIs8UZqmNHLnDl5GMUqpjagEOBEExmEk/6l+sOyNZy44GPWty
bFhkN19HRcph/3lxT88R6w24tsHpldq5/TKZpELW6dbZVHsZshb+8d1SvsPU+2WVOBSfJIqZf5id
tzz+vmi7mhsXDMvIH0iOTgMq9841z1hp8jsnidDhoHNUqDxP+qTys57O5AleGtruulKaDKy45bmb
J0SPXr6ivWU51OkmPVE8pArGz9jxru05+PGny55D62cF2I9qUruRityDPHN7tpT8BdrrOh4E0qTJ
jkFTrLvTwg4kcsWITFE9IUyupEU4ORXO9UxIVOiOzECSDNjV3T5X7SePCdZBsDANRCbEX1Eflj9F
KiaFpqkUTTcVJPgsAo6x0H+dqV9N6pW6PXF1162qCT5vqPPlhG0fyuDnNf9egoMx5i+vG164Ozba
udGu//2jnFmbB5rPDu3xA3rlnZ/Mf7zSjmqanWXSG+W2ANIRRvgrHs5w4uNLevVC0bpG5zS1smZl
HckAhuz3qIcLveiMzvgfb3p50VIowjDGFiMDs2KpGfl+MKaADZpKOmiqMuFmwljIhPjZWzyKLxhZ
QIcvuvMJYVwbbqPKSf62YRYecYFau+900mtI6UA1IbKI25WcbWsBjY4d8BenKCIitVbA2RkQRXKC
ggJEV8e4TeE4y9oqqQxjNgbnQS40RVYK5psVGk6xvUsGCZp4hEw6HEcQlxENSMx5xoYHjhZzzvLP
6YlOLzTkB6liiM7GzVWp9d/U07EMWZ9stvxiIbvX9+UbhSGbmpA1qeQm+ubRlkMTGaEkM//t55xK
EXARhlMcKOnJv09qep39ghhlcK3zuhLsvzizX0paWA4BCuroK+MRNuLPoCil0E0SBzJ1lwXWVhbC
lU4VfXDrI1eosMql0kc1ssS6XmUJuj3pUGMBdS6N02q7IbfMyrVPvMDlXspmVnYpUXeo4JrxaBLb
AAnsusQyslzv1J7l628LvkwoAJ3cb9ikkxD8AmUN3CKaBrgHjU6H5ixpUjjPvpaP/9adbC/GSE0J
hqPFaOZT5Xketym6yqgoHsmryU9dYtKOoTZsebiQvc5vHgAx3eLyyI17mkDltS7+YSJ1jktIt3MF
4RepA7zCoq2w87RNtoDeBTVi4PYu+ccjmmeqD8eATR2csmM/jUc+1epWIrFBwTLz85ypXDHL8W2l
cX9t2gPGAc/tYlF3kApHAg9YVZFj79Prj4XR+gbPKenn5iWIEyeMpEcD5blmhm0io2pHdsTowkiF
MFODzx8ryVxich4IMWIBf/ESrnNBFy9z9NzxeBd0E8ehzUpJtGEWNkg1mTv7mRpoXM8p4ua3DmHN
SxAHGNvQkBgWHipJlAQNAIzqWz/WZxawEWqOMldFsBETq4/rUOEs5tXrK/Sy4kxMrX59/w0aNJ2m
meu8LOtvUGpLR4hTFsjJ40ivoRS05vaAnjKH9PzQqOKmPBgvzFG2tlzZ+Yq/MfyY82dfA2KF/lMt
75O3Vl73FsUsdYFDnKuipe0JQyeXuIZrlgwCWmBXSkvZuxPNpZyEbnPaUvOY1Tu0dCaGtj882agq
LulX584VJqrMS3DBJn7tUAc1ux2kVlSvZCfA0ctDDymim764OH7v+sVsjtGLMFtLEBIJ5iZ6EJr2
L89HAfBBzU7PWK2I8+LlHKAaLXoAmbaMHkEwYqFiZn1deKWY8cuVg6vi2q6F1P7k0oCtzNXbsErO
XZ25XEIcNLE1tbKZAgAwXpMsmOsNSyR80CbutkQu0e9I8WUiUwT1v2nI43CN/MUp7o2AZ+zRUsYq
8vKTHPBs1xKeBbqTGyClChD/uUFbSQxHIYxewgyN/JfgsmzxLV3L3m9GlxNMT7UI2GZ0BXp+21xB
oBqsaBfq231TTQUmLfW0ZfYzMxb/RjzyM7qGSOXPsbVGo/Onx25dJ0E6uUfLFUB6Wlx+nHcnwqON
b49dSa2FmqacmmIvUJdMsHpEPyzWT21r3Vwi4cbuaHJ2fLCbzDMbngG5M+EreRbwzQfagyjPECY1
svDsKnJNB73dizQTFqRbuvqeR8FL8bcZOtFuO3ATCM//tlFgG6T7uNCUTSWj/zOqqNjBKqcdgPSV
fPSSdviSAQfuYDC5MDwHQR6JpUSY6NbPEiHvA4ZZWGiIhPPuUu7uxkRDjm+WUzTmT6vB9eZfBojJ
CpjNa93QIqvkQMZiTVN2fCb72aMtFbfEICwPavlh/LdXWaQMWWSznskwbi+ylValWQaMe5q3jGZf
eaO5/XT4Kne+Bcq4BjJGWesjEXnimzICSkASynAeatDtfYbEMNd/RKYlaXugQNerTQnNV1TTr8Qu
HuxGE7G/3hzvQAzAnxPXblHPRJcoyNgAActc76Ur38zu0R0YEBcNKc9xjI9zRzBap7zMNAOfHioo
9tt4UBnz+4DidqtjKq4LSZjFxkRxqYhJkhFaCJLhqMl/d+ye5QVTcZgAmQCGqSEWo2wlC0xU8c9u
D9vp0r5QeBrOX9C5Atc9RHW/I1TSxZzCpjfcVjgvU6wpHCmr+0Ky/3ID2DiNu++vfUcpprRAPsrs
XFswPi3O8yk3Z9CBSuXHFA1vQciEsJHQlrsIct5/U5RYQTid8owouAXoI9TtmcIjIm9TR6JntDeX
vK37k/zBj0nAqMiYbA0IxrA2maVXoHk+ZoVb4g0KKlkP1l1H71npYKAskifeRZ9EUi72E6EOGjmV
es+IEBAqnn61FYsFlRiUQNSTfJwMI39XC6KTlB0JPdTiR2xJvO9yT+RvoRwsjrhA8qqcBUF70kWL
FU5GGNGZHK0o8vyEjhcrMUOvDcK//W8PTLO0YRvNrMLaqgkeLmfe+sw5CWiAKIXpxXKsBMJf5lp8
vnu4fA7VSLns44gcbldRKvIXh3Ci8s7e3SG2TLBqf77UuF0cyBbn1uuzD032fcPt5vkG1aRe5/zM
0/zgpizVmdGXhUX9F4RnMAVtDbxfSIfO2K/okc197TZn+oajV7k5D5d5uG0Sn0kRh8PB1aCSHI8F
5oHAF1JfhC//W3v9mXQoBkVMkjGNBp4bmySJiS2MslZhR0s/0z++MEja5QY8IfJdlaLOiyWiQFyh
BIG23WN9673uCrb1xDQpHySfG27IZ6c16q29ImI97jipd2O5/eOw2D1y/bSw8LPd4RuFEKu7bl8u
Aah/5Zj6DxvjUXXklEaCOSuvHeZjpAx4Yx+hbXMSLWQ35qDZ4hPQMGmNJLTieBHn8WgbCnTlG7CY
bNryNPKYmeV05h5Ayn7npv+nhajk2zVpuZekHZdYmyG6U/2+h2J1FJMFluCBYNNydc+nBQyHXcmx
r288qc9wMU9bGol9p7FClXZ6hRtFNEWcT+o9iqcAtWnW/f59KiFiev03Dx6WeuqQ5AaeKSZVLYf6
oZ4pnj1BAuDustesJgAAFNblFIqSH9Y3KMepFExM7gwnJ1GGIVtU2leVveueuNGbn5c74zkmjhcu
WwQ3TXmEhrnNgLWvzaHxy2omj/st2wg2rD4E3J+jDtWnw1jQeP6MypFQaAbXpRZZK9qbSgQvgbaS
frfG5tdqP8QNbCQyBX27/Q71P9MpAUrb+E6M0ksf5/0I60WConyNA/CUWHdIXwzpy5gAoAk+wn98
WpGgcnMJP2lDf/mvqF66XhjyB09HN0sc6ySf/IPbXDdAA22KDJGX5AEWDaGxdNRTUp+/rYobLNrS
4s5ZELMqgAXZ3mn1LuVhYQV276LZQOssfejj9c86/QQeYN1tLs+eUxMDRy2FsDcnWtC6ZdkXbBfI
EZasHrOmhKaJc58Qd9idE6qX3HPzTedfs52xky48SDF9lM7Z2xVtArgZg25SNNP1gIf6wLYtNCP9
r57AqW2YS6le0dPQnSbDy8sG9omakALFQPhjEPd5JVU72vrOVTjt3X1zbZ8h78QxQn9q5G8e9xix
oJwQpnQFz0mF/Cwd6xB0ian1oPAfN44FqJqjvaAKV0Ci3+q5dTjCBoGaGm5w7lqF60ntBET4tIYY
CF5Kz3D8HnYmP56DG2E9R+JBLWUQ/CBCCSMJ6S5q4gRtfLCnYxuZzKbpuvxrGXcAHCErio0PWBUs
TXB/a0OzYQDhjZvU6gXe3Gu6zD7rM2gEsD3ZAl2p7QpQ2OTZiPiDVH9dvVas5xw0F2pm/+S4jbhC
hOk4vS9Wcy5FArCRCSSAielq4CkP28TZ85j49x/Enxl7am3ajbDj+6LDZBDz8GOr8mpJOukyHPzT
dAIJHV1IzOSNodks0eSPvXDie1UdoNYdMWVFO/tDgqWZqSTFs9dnehq7wg0KFnprQAJuPutIKXkm
uozGIfbw0ZeRUZf0YJJtbqHaZyaoMNcxRk2l9OeMLe2bJAxIrgdGctfSpRxjIuZDbBqnKMUGlzfO
+/mn15vYOaoeoJZqzGuk5eiTQ9wkDOgabIs3rSGM7D3GvlIxo9DFF6V1w5U9ZhY7qokx4SrfnQTv
wZGClg5W44+ltTraBYqIMScJi6uUWBhYMfBL0eCUR6UlSDKG57IQqSJhAxAOj6xyFcgOPjaTJQgG
xU0uPWwrpUeGQc0n9dZJWzMxT5Q/hNCcuun5d2I668z8nnaJsHt/cyif/6hfr1Mpa2Ha3u9tbOwj
+O9XiVoiWcn85d2Ez3yeZDQoNrcEdqbeQiyChrVxjIHdpE+UmeG1+wbRNodCb/6RFxdjS9EuuUc/
mKyE9loguwD7yo1hq/Nz6DAdl7E14Y18aVdlUg3MJpwt0Xj1C2B0KVFKySf5KCmyk7MzpQ0i8QI2
QYVmiy8NQ/ais21HxKkI62M7ItWdOCJvHoNEzbGbTtZlZUsk3fujTTHyowgm/1Qaj+1mhdE9766p
2Rp512HCeTtry2TEGeIlN7hCcgGCBKmTqkhUz0JY5x1NCO7E/3YcB9TDQ495N/WIQmpK7sEaGrHN
HWCb+KriXeuru2JJufVaC3AmS+kz2DMxhHXtDcpc48yYB1W9KVmD12N3M2QNwTYxRl1c9WOO7WXB
OMkOfLC/KnlVHHptNYkBztdYZa7DETOV7cZGuNx6fEaCnN6OQf2RF01MbjvGhSpWLL65A1HM+du1
3QSdQYG18kFz8c/iNFQ+F3HaahbLbf4aStfbSOH6au9Yza9+sL3IIuICz8/8K/yn2jDE1Wb+B/gV
WmhElt+clZKdywd6Wa4h3/Ez1xM4RWSF9+t68UnrgucQ4kQ7Xd1bUn0TFUvkh8513XE9GB98bEBm
Zezv9NZPBk1kMNe1l6tgaOK77CH+CYB9449rSuDf2RB5O2GxpoIH/T2bhIwkpODO6Bol22O9/LRT
24Am+xjaPeU93YRk3YJFxojjpN/rDyuCjtqKudOQk5sjQfr/9D3AOpV/pXx9LweyYDI8Wj8pheGg
ZaIga5aVM7df22Yv40GtltYWKvGDPc+TQQWLWoXiitcvQ2X8RCX7qaq11oOqDmk+/KKim4voHhAe
ptlC/DILViyeSCwvXMVxaivnk1l2qsGzG7m7ZWcWtAmtm/JiuqmdKNiBcxe62fbKPU22ov4JBjWe
wWCl572U6WJESTgZ9y64kQuNrDD++PG9Lomm22y8glLpcqzsSfY4PVbQFFuu+9NKskKsmG4ClGAE
6mUUGB7SS3n3/yRBg7b492u5kFu1twlyinD1ZDe/py+0+puhnJHMM6OJvRUov121vSiUgJ36QujP
mHmQyuXmehcs4Chr85a3K5EwxOWlRbbeSFCffalILwT71C2s4qrB26Pi4oQHuhcIHy/0VjM+OtgV
62xFVi1JqPjsz0rajZFR2O/qp/op2glnN3++cRsDgPgpV3lUfvI7O4mq+Efi17wYd6uShjqKFMVk
qHSYYhKg9Cs/r8ciYFYggzx9veu3S7L5sbTJSj5RoFEsiTxvQpnMxcc4VxXJuxf25iwsJRaP/yOX
8ZZDsHNcHIKQroNa9FVh+hm2RhWhlTjjCwfNfTtDuhKEvGG2Yfk1zOxFiazRFrsUIPosaqTPVOQp
e52IQKdb6hUF1Hsbxfo0Gu4PSAdeRBNB3nV+OhNxKachg7fxfcgFWGeBtubOzUvmhDtOcweqOF0f
6elGumRopsj3sRWLir92ciAgNkhA6d6+CxQrR2BAbWDFGih/OneQhUcDtq9VSv57bJwx74S5yxJW
Qx2F3EpBVzJuFOBqHKMzN5L770tgGyHiXHrsbBlV3I+ou8Qj/UmvB+wu74GuuDw/xUi/VIw8kSqd
8WBZByN2k5Z5MGw2Usrr2UVl7MnnwJ6l8m1uOsdGKnbvTYvCaBgoThf6Uwa8iEVbjeuEaLCWS/78
i9qKtFjOubQthrCDW72Y/5lqxT3HO4+eewFfHe+UZTyt5Mj89dEr1Qk5YHdBXXfuuJ5SdzN/gWqD
kPOp8tSCPwPQHbpr5x+vZbsghz4lfa68rJ/AG0A7MQcUcEKZ76Fdb9qXRkelAdnHyk39g1Bc+ZaB
sVSglZlfexsT6xK6u/l2oiu8N9acodHzelus9piXH9vQlzSfDqDysQCTVEOvTSkD/2ILK+xNXSv0
a0Nytc4zO0UQAOAbv+M0Nb8IYP5MsYVa7Ylf5H5W0UoPbSXkpGFDzpGpTr0DsppbhWNCnctb6DQA
ON0NsSnEcJhiOxnlAKB2+c/6H9Uz2mmycJES+eX4+cvMy2mbEwHjPjlls2HDZB0uZ3B6l83aCEaG
gvU+uWRtHKc3YtgIbqCrx4poHor60ujYwaSiAUlB4wG9QBi+hi9Im/5aNIBecjzSKYX+6nU29PsM
Ix68SC5g30piUgrJ6fRYFYYSJ1ZTYTDoLHHdhnpWHTVOyY/FrfT9hoqhHLNbAmxgQ2rzZxRwEWd8
KpgyiK/gpIrvJ9XIxtQ5NfjOE0w5Xmz1fwDwkEixp0BhqjDOdAxkzwB0VAlPqauMqlOs93Ng3yVd
y38RgJaRFprl6mL7Y8RUhB+diEu0iplGiCzodLhPrdu/njl3iWNH6bhuIUyiWTKf+bI/+RTONpb3
YeeJGA0+ALHzY6CTNZAxNelo1wuskqzgQGR7mOqY5lG4CH+SKTwtmpmrmKyHZSbsM/juKRina+P/
lAWNfi9RRcxfd22ixIV62rNpbhyPryC8D8GLsL3Ic70F6Yr09Fk3PBpjDSVyUvUHtZyJSu1LtaAG
a38H/Zacn6FKpaX9+WJgqz+x3R0acgJG/y0lo0s1SZezUtzYwE3ca6rlY25+i6v3BqpTbbM3lwZJ
zD0ydnss5EC28V1PHd98NpU4FkbOR/NTcbHDyZR5M9Yz1sMMnsLKY7DAlKLRi0ymZdMpCOmnS+bJ
OMq8TMWZCZbSF+8noUVnQJ/LxenzRNOOp+iGKlKGV0QDUHBgRL5TDo6YlX1hKEYOrsd40bH+hd9B
UUyqijq5XrcSUcz1zG2I7sUsvpC+flRY6qt3Fkfnhas4a+2wIBdcvEvxXXuttEJwMOG8DeNMOTnS
wBTGlpBplYSnYdBTP/EsnvOTZiEAYoKAquJhqrSXAiFXriTOZ60M8B0ylU4qrssSRTPSYqTKJIVA
d8CZNUcs3s1sIJuIvlKUZlyYwVx/FOK/POe4jclXRg7FWj3eE7SMk0PdwHb4uNkTmw3keWcEC8zv
kauJtPAXWmKFRE96mN/XywlTUGekjDxcdI6RBqfC5PzHfWBtFVGVeyxutGojgVpxKrlihhwTFOSL
3NPWfRcKMdrnSHRQIkn01AWaa/f5+AVs2ARQz8k2E08Np6nzvuc0z6v5VZMauxrg6NCTBMpcLHRP
bQGtdMn8fAXC3ayzNsyRvXueTUlcX8zLzcPspcb0BMOjCETquCzTcMEQLHkZEvBhvDS+noG80CgV
bwmD0kk9sv65Xp2yYveMa5Fa4O+QiEikbzNip4ozDo68d3KdqYrb3pGFkNStvRAFxgaBQVyYWHXv
D7t7BYGeqp8/0/FFiRobN2sM5zEvfhlXzW/1kOemazPjXuBbSeq+WSznsqRYbsgh9X2QXPTmkY9L
d3KgnBZIM3T5or8/+5wGsfDpeNMINKhi0jYNp+hao9SOLeJDkdHCB4CU4tUccN7G42xXCki0HuuT
YV+x+4usrYO1te/hJEKDkvCgnxKctGCsFahLDsdMLYpKTC9TyAdVEWtULCeKDPafrmOY54Krd0WM
cA3uKelkgRQpAqdK67fDIg4LEIyou2tXM+6t9uQ1Tz1JElexo0xuJXUvxH3YC0P9ABZ/9+ix6YvM
N/v74Y83UIW0VnHyJENLpy91Mt2eH9BXDxziljyQmWo6nKDxGlEhyFOffqx84F0lPi1Fx7VR5yYG
wEAnsstRrF71XpJAfrXFBak/FWu9wiMPOsmkIB4CcJ2WkmDs6amNiBO1bmn3gHko3t5s+4cEq7Yr
vTdUvryeBXtdpYhEAXB6E1cuCuBpaF0r87G+QqFhstOgG4hN9Xbj3m8fCYRYEBMnJlMUdQz0ovfX
uJ0YFh2PbqzXq5CoKzdTTrpuKDzWGAyqB134Ebj8J4afUq09mfts2b07lvBt/osozQAARGbiLz4O
Adz722sznEUahWSCsiCg6YoBGMM/7jTdAB+5oVBDRDTyiEq6OnqItlRjmEr5o+7501JYi/oy63Lt
K0/FT312FKH0ebUMt7XEQxQGLxOzNA7Af6O+HPPi+SZtPexQRUSqs6NXnhtheAVJ7yKzToq6gtuj
hsgK9SGeZyaPILQzO8u7BTOHzwBsVCOfy274s1w2o5dz9E9WIRH62Pehmcuidj5cVeRv6a7JINFg
wEsEtQxIij0/oqCgkU9bnGLE4+vp3sBOj5FMuHgyCKS/0oifbaplA5FQY7n0ENDSAXb0VXCYX6H1
sD0TGJaT2k5JpwFh3Xh/pl2no0kCDP15TxAaFTePhBdti+l50bNRfjTvvyY2d6Hj04y5PqdrMucR
cuiOAjtnyCkKNM1IihmGpcxeEue4XKSJ3T+8HwHP0ESKF8BdBI6oH9K/hWVy64bsvtPw76Hujdz3
3ok85uGklV5gOQyjRJwjb0QQGmwrHNaP4LyOHvtSMRLwvg6cHeEfk2ERxygEtMB1f3tO7TCU7vk2
oz2zPCNKQYKZEXN0PcJGIkFTO6r76EZHBiWOByc+JLdd9WbO6LOm1DBV3FZzApkQMmCrIXxC0Hn6
sS6qrEvL/yKNFIhGpY5ykAhHfEb97oPqev1ujMR7lfpygkh0qK2TI/41J6yMDj+X56NApr0n1MyV
W0AbGIt5QwrohAls5UrR6pvQWDUlI+efiRaLP1b1Em+KrXmtBTEyVDsHQJzH26CWcZmUUYLZNypE
o2oDHZZjPyj84AuIVxZgaO9rpgy0xo+m3dhxiHwfsrZzu+0bSz1SNQxsy7NyZU6X/RboCQUHWeWg
X2BtjlRT4bmRNndyPsfBFWIpvpxiLY8AACV85DduSoW9ysGTTBR+1GdXoi6+uqsC5BNrvaQQgkL2
Ze+kwgv6hicQKQ4DpkAQ8MEy6/nWFY41/mdgVg/MVR9Tgbe47BYlTi/AvwZzf9w0VT60OwrrZZsw
JTAKHZDDEGroPS0HzLJlhULLbO7jYTliZ6ila4v/LBdeiBll1UV1VhXFpwuEKXpD66MCXHqELRrN
ogkoBhXGIZZvFtXnFtEsgFQZ5ncf3d1GmU8X6jR4trcwCVzSRMsjjujMe561ZRsrhwQPb0aD1fne
cBblxmU3inQTNhxhjOIGBRKqs7nh06FNKlGQj8dk1nHKB47OiUkyefozzPF5Z1oZ5LkMkES1+uWQ
fTWiOpdy6EZ3jLxPyH/k2HVKwRPVGIFwUHnuT0zMfqrLd9h/KryovYb3BEfXq/TLq8SDfeYeCCbK
tBTh3Vv9a5QHX2QBm7Bz4Qzj8IsqkFVIVsmieVhvitJoAVShrFuhZSbapbasX47wD+ESBD3fw80n
a1DL7WXGMa81KTPHw5FY8YenSKr5TScKIzjiaa9oOntaaZ98Tu1j+4tGtEQW8wVufnw6WYjXej96
Ou6QaglFm87y2Ddqp8gtnlk8bYkrbI4QGT9uPMbU8GRsAv09id2xU8aK/tVBqa+CWNsaRqX8528h
sB4EBKXgwaVLIwCClvkXLLvQdqVQi6lcyrKEnwPl9TaCJzsoRBbmC0X8bqfF4DmIfdFwh4taPTzG
NJpCAd/IFa78g9RG4V7pj7vtMMDRYi8GvmpHfLl0T6b5mOiF2rqaQU3BFk/yAUYJ6MoFNWj5CoTi
IB5tcc4t+5YugSPMa6feuLFDCgi7x47Rec9ddrc7U0OaJ326/i+q5ZmG5y8rJ3zuLvy9ZWdOPNyk
AwVZCDmcLhMYeUIIUimcQL10jrjm+FUyOAEnht5VRjx+hv4RbfpnOt2Mb62CMtDzumLb6+fU8aQX
rhw48TFy5jDaxs5lbH6wJYAy55zc/BQRm+Ah3WeRK0Pqeq8x2jXehC3tFSlZMTmEWK2jPSjKTXME
x2kF5GLWwWLprO3SHHzb+UTyOh7a0hbOzvG1i8DEsUhjsBld/5C8UhUUXVbHxIT4d2eLAI5uwFyA
auBZVeUrR31vOMNrKjZAL0MEzep8K2OslLK9T0+zQIUMBxqOs6IL2I0e5OdCM88aFTfGCxTdsh82
ghYgxjdqFplFdHLY1ky2/WHewfcNxombl0c5UT4cqg/0vSGxv5WmAYr4Uy9u2Ag70CvlVAnVAYBv
Z/P8kYtiMVYVw4+IF9myj5Y8eNKBcXeAG6n2fZh3Jt5ijZ2vgsva/Bz76X5uqE/hf8LJcWjwoYIq
BdBsIC9MSLY4GAcHmwNsHbY7RZBQYyXFm1pEuK7gDxJIniqVGP0kjYsoKHFaZw4gAXypzxHevj1O
l3kSbrksXYfqVovh2K5ycJ56bBJ1X+HwPMUYZ23UPcADzc4KJ9L5xIl3BVZZTFEGO2xjgZkSM5CU
NoafGCGYqm+uegPNWrw2FUgYqhH1JQHn86zLknm89c/BFVA3u9GpEm2j4eZDF67CRFBnxQ6CVDrF
9JNI4eKfE4q0awBWYrmTPVGXZHiadBuWhAwLXjJ8c1XXUqd03SuOrnhBx6UP2wLOhOePLqMT3M95
vE82zuYkVBOz4xGgxZVp2RpK3SxdUsx6wK5rIPxUP+PXEB+0lKZLxTvDPs96itgXBbgEqO3zPcYr
6XPDfJ4M/1oh8quj6Ha4okVxGtdx+NbBTEJy8a3Qgo0/2DeEROVNm0p7uRDSl+eTzXCDNSR0U92X
XkQJK+cOwrafIvKaH94P8lwwzvoRb6WK08FEXwKQ+JPr7WYVIXQ9ETxnPde5D4ade493aM6625gv
XlTpqHfLgUC3uqo9avFfXzIvN9IE1mk+jLrLCVx3hR+gjt9Xn8P4754navwqiynmAn/CGX6zIZ4b
FwQjKkwqHYfpGaUvy2jlZZQYuYJhK+EdaWBYvGVSRBlUoNbgYXL/0bqqWopl6sYCvXtNzgRDNhdx
aBIj4Cnp9PnqaxcyM9Ohatrh597Mocg5KXVHMM/u30Nv/sNwX+8a759h47hw4zqMUdJ9153fwaFU
mSW+LOPEURVQdtcFPAqyfx6NNHnH1BuSeRxunMjZgOviZSDDPetz5KAI4QtFELtzxyo4V9tmIE5m
+Xv325SE1lHzKoc2WuzOV/zRPx05LT0tIU/G0/cD4GI/3rPtqpswD4ctL4JWX5Lnsx2CLr0+i0zW
zEXhSKhQZyHTjaRLpOzrDckn5wLXn/BX1cpFcIRck1empVs1tMzGk/D6n3zUJtiUI/ah95eUa2qW
lGhjVbuhsz6dfZ/3YYKtH1t7RU9XxwIT1BhI/9OEriWmIDE3eTExfHfMOVUHJGtPgyP+YDJ7/1j4
J8l6Bt8YT4bspUsAXDyv9zXmOldgXr5mS+nf11AYh/wDNF6eAG6dcjk3PjkRU6ZN3dOPm1JySV91
OtGRLHulw5e23ELlSehZEDcb/Zs9tfokkN2NqvecgojJEcaghvLHU3yJLHQeWZjvlswHnHPZf3OB
wpqEPEzUWhAkInLvft1iIa7w5Z8TD5x2ta5RLM6aBXF1SJQrzGNixhmXSTadsvTOYaoWL7bLQ5QS
rrAxuBqymGVrgyH4dA5g76ri6+ngDOW9XgbGNfkpFevlQ3wkYcucAV1Nv9q4KXzLvKux7TQuAEur
howiitFevYQFPWySmGku7z/XranzhK1vXow5zRoWrIHMzWw53mPywzj+tTblsbRNiTGUOvtevs/V
nLaPpxqx2wK+NVKf9+ghlB/HtwB9LMf8Q1jv2zv6S3tsZUGxMtt1RQ8FKnqoUjD9SQwgaESIKvZS
7rFuu/kTT8XeCOP2IfxH8Li/sRZp/LasBZQSP3++MwD7cy6VsXKpDccSqbJwDlzu03BM3h6hk1g2
AcNsnBvB8rKIF5HoRWCUJ4fizem+WuxF6//qFGn5gBU8SiFegwpO3cKe0UYtsIR+5O9YFhVKaxhX
zeofCmCm5QXfKkBTXAYhFX7s3o5JDEJbYyGcydr29+wgYTHGClUCAfVt/SZC+qIXfrE3t2/oDH7y
8BBouSSFv5GjJZWYarclyaqkNBicAgVFu20x911fL+gXI0ra7Go7P7q+UEpaloTFsr7sbzPOlqf3
cOtsioqdPWIv2YBQxKx7/Hrros4yOVoyyBeBaFyZ7fTeR7WH53X+9DzaTB4QOEzpH6fAnLZCqNsp
CUg7kTcaJQc7JsqpeuQz9fWxwGh6559vJd2x5pOb9/ffHke7Iqj97RxJgttW/d/U350702TV2836
xMJOjvjI5QcjoNtQyB4AHNtMtMuYCjo09FKlkk4oNdd3ZGPXjPWzkiGsvzHLmREFOZJYh/Cl6qen
RAfOnnSRyNImIUchDkWuQAmbOqXp1bY4RUspr/I3cbI7b2JnP3GJser29DX5BK7x12DApplQxblf
QZmcDEgJoVr2ILDFhgDZwlZoDi53iv5m5i8lj+9Fq8JftUhDN6xr1tQEf1XrDJyDow6J/iOYNNOp
gse6qLFkDaYTOnCxcN1dNaLyrGypNqk8f67fQ+iM2ctmjlmtJAFP9OOk9KWjRb198g+bB6s9DzoW
+4Q1zaH7XAqj8e4wP23OqH4DO0AGiT+tILRUK2N8ZFoUacurxeLFAGMa7+/ukXrk/Ja3vx+hG+9q
X9ztyfm/M2xHfXALBt7V8V2x5Nf7rSFRdPz+4DzeKYudxzp+xWfPxNCTp4F7RZlDNtFVSQL3ciof
e13Z9d958Auy6cHXaGpOdyR2tb+/PUF9iFoHZTYOCNoElKSqw3u6wxfMO8V8U420+MkU6npZ+EsJ
pPYxjAWN/IEZzeEtAUh0+01qeSS6+gd3t8Ey1KkSeGTlI7fmPAl+GgEI6JpK8frUWPZK4ZRp935o
6wGDHal4d/o1d3cU+hNa6Q+7OuHk3vIkCAF8xrTjMTysgP+F+94/Y+I/oQUk5mN/An5NP3eO1efd
PtG9RrWIj3BdlTt+dLVLKQ+QuMj+SUWaC1IcMMXG2z3n45fR/ShpG4dBolWQR+M0E04oOOVMZVwF
wwSrPA3TP7zMO7NgngctZ7Ta1sTNalu8qLtUQ2xiav61fHPrnKp57pTmoj855CLfXjmPO7mFteoI
+1eRb9IgyBNtGyKjvcqhp7Iu65pq59uyVdHZwZTeFBG9tYFRFgA9zgpqvkLoZXlKRhj/9J7nn14h
2QEbrxbHda6n7UDPm5g9JzNaNh5lQNQrVlIVS0jx2FkBJGsxvDiRw35JbsJkbxuCbh4fMsXu4yxZ
pNYw1B8zLY3BamkGBcccSHWopKyP96hJVxG2l7snbK1McaQxxZKOcr8bZOnbAad8MVjS5osBb72+
gTRlViAVhrHnbW0GffvOzIErIaS2jztMpJGjireX1bQ6ZGGD7nCIES369R6xFWW2pV9QXN/qsI8e
FE5N4s5A9Vw76MyXW34/MhzRjE0d4x9qR7eL0zVFXQWQpTiKGXFSJ0a7TIw/ajkVUrduqRvfFpHd
UYEdMUYalrbBL2w1UHYiTwRjQYk2Y1p6MH6Dqo9bhUWbqTmRV7LrdaDEBuJWoCxNtaD/71yLGiD6
VrWmJdx0pWHIPtaV6aI/2RnzLBCScxxcipE1T613eiu9KTzyOnA2LYIbUL67FkD07da+ReU3QyEu
XiRfjPx8XuT9d1OY8hHBJPk6rsIoimmNiK0RAETrjteWQOGiM/BGTtngeZ2q8GoiabU8nSbcfoy5
ZoTAl5rrBNu8tuwboT26L7AUvMGY7lAhg0F664IfX23lSeXPdyBJXP/40HOIu+hcaHCyxPC56FPt
rLD6JCd+m1qOEMd0cjNhTnRUp1CFx0LhENmzmWm4IlBYo+54+6jJBtJruNg2g7eELO4U6JhoT3rP
fqA8kdfT8QDNkoFCzAmd5/gcwJCkBnf9+a8voWkz8LDHG+EBG7cDyC9OATlAcoHlioM7NRS/N+oS
Lw+m31Lid3v0YO9xVNRu5PYqbf3DMbp8N34v1VapmwvYZ+ZPmQDRYBUFcdZ56S0yMHalXVpw5/N0
f3zWhZmAexzuaCtPHQhhNfZWHbounzfiaLVWhoI7MC4jc12V54ClJB9/2RDxisL2P4WR+uTkq+DR
ZWwbL20wvHCYz/erdaWHahV/68BjSBWnsVtWpXMWlVYHEIPQk9aa1NWPpy6bPQcEdQ83/Nrw7YcP
Piof3kAgDNyxf8yTAmVE+vFYJQRZuXGJ3T6ktS3Rc2LyBs9THx33217WaoLsZgzPUEWJTPtVKQQE
h5/USmXTcLyPjsYyXMOueUZ3+9aGIupua0r39HP9HWE2f0Vc7KKEWraMECJ4IqJonF+ghVnNCoE0
P6M5Wv/fjX8jcLEFph419NuoyIDkzjsRecb2wDilTKh9nTNjJhvZ53HA/+XbFMF2eqE9Ip0oG4p4
UmtbelYNKmReo8+u9IVr764xr8or/Rv0P+aQ775B5FByZ0vyWFRhYqdAqWutK11GUKYaPvx7lliW
LlB3QMKuziK1rToe7P+3jdb5t8vqbnKRQRFEZ7zK4X6jYMTsn7Wu70czivTM9VMhiR+2iWF0OADP
vQyqRERCMcYm+rzLu57VMsk4JE84Uk1s69AMOKTxvFl5D86RcsNdfaFMKklj/H1LbUD+uyTxLPYm
CD+F3/O526higAX6KGVp6ErPxnSjHPEjZ0IMXVY/gY5FVITZTi2+N4hLaixEd7gEThVz6wH24Gmc
XkuLw3IzNXJjK7bmYHKrn96aDtKZ8DYhwE4mQzaN5WX8pjnQ/wn6DPEDf3ZxwSeoTPc7uLIsEIQV
mId7s6B5cAookLFo19yo08e1K+3xx/qmApvRVeqqm5/2pvsfFUTMURk6vhoGTbUTXXlGw8D8/sRL
rArUh/dk6QdLCVkMR4c7bdvAz7Pq2pXEu4h1djt5BUlz/Y9DlI1dnutZy7n2Zn8Gv77AKule6UQi
GNXgunxQayeTuSJNK+FhAvJPGLytmGjtByIwlSS59Ot1B0i3mL6m3epZZnO+vBAY2/i3hv5KIpgE
eOz+4ple85gLU6lUJDZ/yg8YWbABG80vFf5eMhpVUfpcecAMRh4dzxqffCg8UBZG1IbXCzp48Q89
Oe7bXb4Q0REYR5JIdLpAs7g2IrnS382DQ0OOq35RY08V1a9oYzA3n5dukncUrCADhQjUFjeY7OGk
n8LsJmYrNn0FNTmvsa8+Gx6fdclM+VRcb4CZvpf/B1sm0ZZXOkvqzt+KW39fJcSFJ+eubL4kD/IG
eW8OXFlonGBhNdLiWvcP2Z2gX/e4PVMqsA+SzYu7axzCqeOEn2qyVgjikc+5Oj3DW/lTyvp6EcSa
Sv1yGyiuTblaRiK4uYuf8CI2Zj3GyRgOFbKlwRX8g05188cM8gQg/EztmgWZi7F//0BYOsw7TtkT
6NF0DwZJC3WTGtLejHgiCfIpZ1MdIfWMKqsBDMGJf7NU3B8QcRKbVHOQEogPYhKJvggDKKky4FUS
zHoKXfWBV1UYVqJoxHjr+QQXIhsqbKHWbQwFn/AU1cE+N++QQ4y/kmxedZBPt9Buth4CcuUpE6AU
9+bomJbn+yxqh5uQ3dqqyWNEmO/FMV7ox00DBrWrSZBm/5cBCYR8rvYBV7grIXTQcwRfMWtnvHwm
YKEGCLKekJr2ZhBg7zofSeGCAZj5KyIJdkupKSnFB37XxYnpmTqQnLKRWhvo6sHI5zHGJxjfqC8n
fzighzMAWlqmqSTnMMKbTdNTYw+4gw5W0mcOI+dEJmH+lU3SrNVQue0buEMS2AOM6DxxCdzEsHdi
B+ONeRCYnpG/ZDVj02P29zLgaFxl1i84yqrH0srfcKzjrNbi1yX1K3Wwgh0qAc+4onch68b6PAnH
yXcz8CUm6t3saj+KpBr6lMzLCLbK5N0XUMONMnstLmJuwB2m7tiew7nMtmCOQIq2vH2fiQQiXsIA
vvg0D0EM/D6J2LGau9oJ2pSl7tG6EasoETTm6b2mzbc8OyX6TVqojzWJZKRM2linFdhJ3txoMpao
muvHw/dcD/XF/0HRThWhichzA5TwgH0YSw7IJYO1rrXEXn7VnjZ4d/Ev3ZMqOAjVdNEc5qh8McLz
iUELjN74YXUuLdJrx8TZkApQW829znNxGEfkr1cGdiEDn13mU6u9OeCilymr7Z80tJt12YFPjMUI
Ar8ZkOrXI6VAY7IYa5Qwa5n1rakFLcPUATy7xm6yxStT9ybyO+J1/uZfg5BEU1XOlQKHg4KNVRXr
1988KprqK7CZwhV4M+DH+U/FVY5nH+JddS59vhGItquz3cuYGXzB9BNcoQnEkCDbeCCmo8TTZiyV
wRYOaYcW22BO6dKbvmR0iQwNFsaCrQVh0n6leidBReFUk6wrwoqvaiCZlFIdKo/VXgYDsnxrtCHM
O4GP3Vr0/en0qlUsobIZSgfi31GCfqMTtnLGs6fhIj9Rx71WEsrCM63wvp3JIJ/UW8TfMn7/YlQK
/QFHx9kJa4yWDIthemwMADpzh94UUCUS2PFm/LlYBfD5Y1IN3QTMoDbPOQQl+r7ZpGN0H8m3gNg8
ur0f1vipYN1zYg92h7r+iJNXHYduZi7LYUxN+xb3SQVNYEdMBhpVPZjgPDngPYwoDgN22Gzv0fnF
SkcjeQcysVwjb6tm9bngAs8JWbm0cU92V3TPxQ7eKjoHYC1R1Dg+NbJeY2JhdDuYNWKyAW0UIIBk
KZKk5sXMlHz68Z2GQO8WOO+Jp/fSqTyn0kFMi2lycDgghGXjVGnuJIG7zTrHD8LxJ0xqve11U1/9
qzJzwLs9D4nYEKBA7SyaDHwXq9Do3M2yZoNbCTeBS0jObLSUO7VLFseF3CO3sQO7r9rLtF89zLpW
pb7GUFw413q59m4eIT2eHmf+PYlD5J1mqnSjONxShf3wrUvk3N01Ay2XnL3uj/rgBxH8PBy734uL
ljljRHOLIG8BGibbwwn01rz7CQWwjxiG4sWcHVBcYeZWmtJczNtu+T06V20RaGvrL/aoNc9qfIt8
L4QOjgA8mXQGsrCax3DpKdOY7J7DmrXTl5ir1BPu5e1r2dNXeitUC/jWHrxcvm5YnpFvxPn+lvFr
0QuUqqyZPjRWsBH7RwaW4gVhkcK98SS36x7XKP9TnP60MlJWhG4aAJW91sfULEFeYVotojKbdHl0
/uglORG+eFUV6DQahJ4z8kIWDqcoAVpEptbuzGYx5vsRifCzAIwB4xpem0Vw6hKSjVL6Kohzr2hv
1+AcEBE3xjFB3CjGwszrwQ6wI6uyY6IwArdFc5Jxu9BLZG3cSgL6e1J5ogPouIzd3B6nrxYkF29m
0CRIBvfyPy7si1oVbJXaz4LYewKZE+5YKAAYTbzrbwb4f8kL6bzy6/hZ9npsrTiByCnHDQzXVF4b
HnwTmlWcZG3LW+YDqV9FzJRZvsZKoCHPsuuHYmsVphmIIvIHK20gv8Ek1hxcPbCXoy/QjKztgzOA
l6GiF1jA0ilH27dX0ao49ZByZHgov4kYPp6uHKK5tZ0aakvj/FXbStKF2C4wxHMiWjla2yxSQThH
HlwylOQqZaMDdpLYtZE4imrYNnMKJxArcFKWXdXyT87hpgAETPbgbglUuBs5AycKDluTcCGsWOue
whXJ0+ggeXpBkcbGGjgE1iHPdA4lYIGSAseb2tUSB03IMLJoxwD8CPh3uCA0r6sQ86JSloakuAY0
RBvo/ht+YE/fzVza/ETMJi5Ul+Kz0NguCieEbA2mtF/WdVXc4iHbzSFoPLZ6T9KAfNl4LcX5UCRr
79JxEvfaolk9vw7iaWz/yvVT9xFlTVK+1AWvNmiiMbYsA0qXmkQfgG/kcLFp1ZSd+P1qntagQhzL
orb0v3xQzpSDc+qYkWe+MYI8PZRbdToc++xZmhzkH5xc0+/QmYYIXxwZtcH62VWdgkRpH+8PckJs
bZfcmDJR2MHtfUc7q0XKK1gu9ItunRUftPOOqQflRwsJa2ziZkAk6/yD0DRtfc8J1mBS9XlFc1qF
u2fxpgjovfSC2fKY8QYFSgHsgcaVcg8cDGA/j1cmTm9CHiXwU/u8AEnyEs7YWCcYDzWgEuocu27L
S39+vjvFqH1irY9QKZqiz+b9lYzOIA2N+s2U+VsmXdyGNwaT86BbdjIGhsy1gOn19XWR6osoZhMj
RKc8voAebiaKlF07qnztxuh37Ib+gAexDlMKHVgxJdC3bG9YtOsM5eDIRF1OsWkm5rv/lpLKtGTr
zYYLOsDv4cK1OirQ6eS5wioAU3CA1bLQ5Btlc7RxePnMX82EFZaT9jdhcwR6HzTkksLl09wGMPYt
ywHB3Jn572eMYhGyK1Bo0FpWnXrDW7d7Qhem5hnTsNRZ5s2dzAR3QI/ynIhE2pRtXds8y9a7RSZb
M/8xuL6HwlUl9b7coSxKn7Oi54x4xl2koqNX4dQyV+Q8ad54J08GOjHKz8SIDK7vhPVvDqnYHMhG
ijJm81Zyb7bJNlDop13adcirovhgSs9wSO1ZH/UxI50Rx3yU5/f4EKWyTOzNpDYMf6dR1xinCWUF
n472m0k/kNGFiiMOrFr1U0vzYATOeCVFVMb0E5L3cI9fepB5N9ifLxhsS1D5lIGNF3OwciAVRd7O
DNd8b7yA3IgwwhYMR9PSXlH37yEsFh1TXIxManyPxnzndDJ0QtWP8KvmIptYKePZA+A/ocTLtcZy
wpEORr2ROfmETJoVUG1DQVlkjytrDCMrSobluZW8Dfmqvxpf3xEv1eQ5hqxCO97uMNjabzQDqmbH
H1v4QB0TGRBjojC2Bs63bWEYIyOFK3OGyXiZh6pFrqigq/1IXNpo60YloNnZDUQdbOJ/einNW/9g
ACihsm2xqBucTqzhwyuPZLrCJs7hrPn0ynWt828Ej/k5kIyX+4M9gyJQJA3uZVW1XYiF8KxaJAbs
l/f+1aez50Dk4Qxdgum07XzDGVAgJhBoMAqpdJztYmobKrs9xYbgq0os+/coWFj7twxSd72bReaX
VQ9d43CeXv8dyHDA4KGo1swZ5qBAkQGSwjnmF+N5wTwtww1iPdGj8DE0KldRwoL5cnl98fnS0X3L
Ye2q7sfvHGztdUKvaStwgOXQcm4+hm4no5gzjCLr2CGbkzDRo03V1VBUMy0+TMJvez1YEhlwknYl
iLhuIbI1sepsXfxAx8FRowHLQPe/JK7Oh4D8i6pIt78syVbMS1feDblTwchc+JGThukU6GStp7/w
VaA0xKxsjvbg/UGCIjVr4JByFhNCbcGtIrDyPbhoHNrnEMxMUgZkt9uIGN/CDl46EvRCJrANPwSG
5TEZJk2ZIdltShNlBxTSa9gZY8tJSOebJ99DAjg8Y3auFbnwlqu0l2y5h/joH6RGSWovwIYMu7sb
Tjzw+yPRISzN+FxbPv6/+9tBjAZkpl6gZsHA1db71W4pdMGQ6MPSBUQ/KJvVMvUHnLsQDbH4T0UV
l4yww7Oe040TP28ecsG/6URh8iZ+0CmuGjoQ4jlhmXbKyKVq9dlftCH54y1blTzVUzQiWfgw7aVe
PYK2hwK7G3CrCLpMt+WXr/ilMl1K1qAOQq97iRWTAeX8leL7ZjDcUppEugSAE4G3CkRihm1lM4/K
Et8H+vA1/Wk7xowah4c74QF3us/yzNIh+X6BpUSurWJJjyPO67r45X2Zx+P0YsgPO/R6IvlLvO2J
GUWnTKB+r9IAmLbe7ILxKQIWWue8Nu/FovU204iMXrjjdbMk0PwNzutT8U6eA0L1RQpl89BUj7Ys
NWrn/L5AEwKvUlTLiyu6y1y6OcXBmsUCGyBxifwI/LquFb922nhEGvlXZwOW0ZfCMM93lW2hNJ3K
6Lw8fFJrxv8Lj11g6hV9PBcbPOkzndGgMHxoBgbRqQ0PNetf0wa4FlYY3Cfww9KimWh4bYS5yKyP
H/aPaFI0sL6ucPNokq8WEhjL4n/cn4voxwGxeMq28+521W98VGHfuzPj6BsrDeR3teH1L+Tf+g/w
q8dJyBxHMIraJlqG7gHe5V+sDUJ8gPIrBqo7nbFq1d1VDzi59WZt66Y+V2mR0ctm523uyUcrcTm3
iQHhWlMV2IOKV6UTTaAogtDE7BU4uEuhB7cFPLIQqHx3lw5nNzyiBRCwN8lrTf792jAhD64wXm/0
Fb5zKuzeCxle+abDhJn1L7DeV1XNxMP1vJegTUE5HuJAacG5NOE8GfdJsDaFaWvsxQgk+Xa/RG53
kCjrYgvpdEkBqyJyK/XTZu51BG3Mb39XajOXnc9Up8ZEkRIzGpUlYX8/6cZYvfGE4gU5lVDkHY/B
wqHomOEcq9o21p4i1R2zCMrI/m11R6APk/9igEbuU5V+FVssczfeBPiorFT0ODr3dsAnUShaj1UB
lx4INB0pmxdGdLC9o87CjtOs2RE4mMJ3MtApymQuZSRgHDsC3X4i49G3AtaIlO0OQkSNMTXviosq
eMC+VysYdsXh7CgxZ094uPJIhDjwVk2KCe61WGzyiYwFCfDSfcauq2+O8ackFn9hIThbrizoieGt
EHHhqi7UYhEaN5ALvXFh8bx0Ps8RqLASGZuEiNil9rA1XgonsS63X9AlP9vfTJt2bpeAGTLCbmqY
E74/TjR4q37qv6pObfEBoNRRv94Picc0r5hj+gkq3A03xL2qIcx2L8qi+RM8O0cUIHKbDhDzEEcw
Gf6D79EhIClp3IrihCXu5kxqXGV13GLWh4wln92iDYGZsCCgY5f3B+m+ffg7S7OheTE3Sa6aD3jq
qONtAa8BRyNQpKMcvDRhzJxGQifPWcOcSFvOG4SttfrfAnfxjMl/OYMhIab/YtKQ4krxFdMW0Zr7
Nk2BRQnPtOYwXVF/8lPUK/sl4zfw1cK4eOPSNZ8s4VDUp+OAjd7eMMRFz45jWJ+ctaSBiEZ0efEv
aurrotmvaOhH37y1/g2LaH1jBiNPPMl0koMtAC/XghIqrfBkfFRrcvWqymo640pxroYphQYz4yvm
Qtaw9zZaiY8m1UJf7J0Y0anW7q9IQHH8HSS2bvyhCmZai/lkCXFR8QTT0De/V+7ByaB4PcUvTSO2
bwKNsccDGbxOFmuBylvKGSDNicVgMYpR2AHVY+OfHpxlbmVaKOeqrlU7meuGGBQRDPaICwWCbqmK
echVWFOMK/nAT/Ih8JCbh8x6zPjnS7mwwifeJFEO5HGNN2n5Mwl8/UPWQdXNj117f0oPiwgypXaO
dEEetUs4R2rGpysDM2e8PoGW/gYE9B6ueHRvX1MFfHdS8ySCuBPiyFchj190uH3ocV1g27QMMTGT
RcHjmwCbQTQgFWAUaIethwnN0QbSOg/t/eayNwfzipTqwlYuLpiuk9Gcp6dg2NrfZ55aN3hrvslh
zr5HGGAYYe7uHwFIyk6dM3MbaS2m6w6MYtmvtizgzvs7xLizBeuB34ka8pQPlNumXHeftT9Bjk6z
tQxH/CoKBz3aBwc3k9UXa/P1+T+KZ7Lm/g6/LkxlH9ats3jzjGy0M/oTBSIf0mDpKAL8Op/RijYg
8N8edkaZGIwwaDDbkVML32PxEiqzoFOrC4D3+ghn+9l1Y+h/eRNCw4WsKxP575G3SFoBkECB5MQv
HHand0xMyix0Y49gS+vLFVFefBBvimp+q2J79GgVHy4k2mboAyPOmeCwm8dKxR7QpgthAu9IMvs4
bdEkiEyHaZagIBR+Pfwtd4DdKXwRw3FEl+4KHNL1AeXxJfdBuouoxKmzHoewcq4w/zkXShWStbj3
K2mzWIcD8ekMpZtxA+8if71dW5ZC2mohV3pu9ipuC3KcJWCc3lBy+bY15wcJQA1g5YH7eIpk0Qbh
hjDI4ByyUXXgNoYYZT3YFssyvo09iL5hnUSVLMQBId3+TVY3ZuGFmUj0D2nqQ1ELZNGviLQeqQpi
dgsjom40exfJyXqQFxaB5ti1RjlVfatqj0LF2+I3XGhEsplP2cHj/0vyk42yUMGasBjrOrdJ9IZn
mwo3OUfnAtKUoxO6NZ0LVoAPRAm1rmm9BbPsYGjO73h2CONK1GDWm2mQXJnEcr5wKuBG8BGRbpal
9e/YiChCFzljA5TRPxL5h49c/k1ZZSTEAPMHQ45I7M62mVVSUg3CToviFPh4e/5PLD5PWxUOjrxj
EyDNSN1naELnOAvQjcP0FwMfbPZIKfiid/XxHEQXdWBwo19hJ62ahpsTQV3zIZ0Fr00zgC9xqBE4
A2HXoOuJoXU8N2ah2c4pQmEYHZ1Y47bpp02G/y29pdEKhewe/haZW2K6CRidchbW6ykaGaUjWNz4
xzRSxmtjwKikRZuOX7btWh8wS59Q6E5chV8T1Tj57Qa89jYKN2ZYUI+NpltKdJWBiRstnql1dNJF
DTRBar0bjrzQS9Go+07T7JSuZmSH/DEwK6+qi0BEnUezUaQMskBdfZJfsM+12eyf0o4koJtFsRAC
lkIaTDay88w9Et7wlpRxCLiLbuydYNM3zzSxj8OoLtDd+UgXWlSnr24pKLAZN+mlHu5BxKTkFhTw
wcbUDaE5hnwtgPMOHcCmk50MiHhTT1ideWM0RCttguwpCn6OFeI7QP1LITQxnGeWBK6lIOcTeQxK
PYKIL5qPX6Qll2ZUUjHiZbvl/v8ElmBYufRvDvQF3Tj1y859w335hlDxcQHk/8fUZReDKAFUsIqJ
1pxcFsg5HyPTQPxps8NpImOpiBk+cx+xS5cT0TTYuRveBhK16/sfl8GX3nCzyeUVIoK5fSjuJpf+
hdXepNQfWUyWFEky/PYRgGCJVcW/f6l0O35qzqnWc8KL0cKQMNg0oMldxtPij7jKgBQSPxwPb2P0
n4YJ8J6BqRKI0Svqllmxx9tIjs+OM8vzHqu2obUJz2XsBmIKJcw+FVcO2fRgmkQ57ZCsfOyd571x
Gih99iGzHGjQIn/VzpGYf3zT0Fwczx+kHGTztpbW9Fp/52PLpzz37+2IUVkuAtQOb204iXT+r4q2
Qq7q6ea9xye7mC5W1vcnFYD+b0Do+sTGPh2BCJbtrYgI7TZIrVQGKZmZ4qExk9iG8PQE5vOvH1Ty
AcKHxfaIyzm7ElIBNdhAO9EJw46slnGNfRUpkRTEa+hz4F0mAkem/jbfyyYNXd4SPLJamrLLV7DJ
LMjufv+c6vVpknZy6Ujana+bP9Hb7dlo0wcF5zSDpHdb4YaVQSihHpkLvqb+5xqZ0QNJ8nWECGfQ
eXeCicRv1hlrGSVYNaJURbZ7bLJOfU1Syz43D6vli5w3pQKuz6vB7imuQzzwM3xK3NXGx9MS1Sub
79b4S7ss3m12ngJ2Oq+5ARRvjsT6tuAZXqNfSdT5UsVyBpdC8fcMi3hmmwQBXUi1SJAqtPdSi3BS
IMZXmcBrFghrRRDpz8JXPapy0pCdPVcKfO9gQwmFNfINOD6fcHtl11ogbhevDlb8QmWC68i3xEt3
qUKNk2PGkld2Tc8GoEJc3oK0V86jnVbg4P0xbqpn/NyotKiRFKraT7Za/vFstlUVIOxtW2hA8pcR
stRG1cq8hzJjfkuFsvByN/Vi9JqLgckZpLihBwaoL3KMprOy3JCadeSP6SkjeV0tNtH4SKfs5ddq
6F37XhahzBH0eRAEm67T8c3kPrWgbW0kYM6bxcQfc0YAccJhuXrGlPtkcPnUIdiTP+oTuTxRyH6s
rn3Hf2UU7ckEnf/B/zvEOKBBhroi8iMkicKtPt1kTOlGqOg4sdGEuRmFMzGgnvfPNHOo4UwMEkGp
2/lbjFbxzQQRHqf1pvOQsTksnGE9mvOsUrxxM7lDR+DHy1jiPCtxJ7A6McRbk7UtRdkLQ+tH1qjr
civcxIqLNVNlK301jBx/cM0s6UmYcSuERvbxBWVi5iSPVHMiJ+vnzNRe7UE4IojrSVe0y1KbAxg4
K4TS33f7YzEi1tX0XhFO7uO7V5/wktPDPPTlfLnzyfXytfAY/FVJ0oBzVd/GxygchKyp+z9awYUL
0ptzZvKQIzQiJa3PzEVRFmDnv7Rpvyq9mTDHMlac7hv8pe6jjSWYiYlTIwL1V0jmIa1CE2ELXy9T
C630o+eSTM1cDaUU6QueGXypHNxaXzoqVvBDRTbJY/PHDQYgwTtqEzlQcu3Os0XiplzFDpggZOtv
r9Qb9J7+hFbZ3WU3Qq3akBQsh5Ktc3l15bWp2h23zbwT7WHINDHWfiECoQV4IFQQyiZiT33x7rLS
q2v2ACwZUYGnociMvAsU4mLLkYOH7FSBCSKAJlzZbkla6Gv4g5XVLw2CeG8YjfMFFDWG0EV2WA0H
m/f9BSk5zpBrSSNmsU/vyekBrNfqPw4uiNb+Q2zuYPrhrv7/BgnArz+LrJIQTdY0+LWeerUAA9u2
iKu5QyoTLHggel8wpRvfBv367mb3QMdQUvY9iVKE17QxTvIMA8KYFcSZwID7qTyrYouORtcrsk+i
BK7XBQdshZ82SnDuf0Fi4FByYp3KpkYHBJ67xR31rplMBJQYH/z2zkOqjumXPP5E5zvwGg67Xyug
wyRZUaUkfH4wE5NFugHyoQZBmRAuePULqL/FykYh72wLlTg30r0cjDZnPPKt5zTAVr9qKZ2BaxSS
8pj7t08impk3RZhuIv5qBxG2/d6kzIhDEL0PsuDOC7H2bYTLiyqh2UavOlce8SyisdhaKiUuV8Oa
6ueelWYqGXRP1YtOZ95tGCF/Ez0qdoOp7HfIRrzp8diTJAekM/mkI/vEmvONG4ZojmG6OLSj/bqy
jBacwNmbOkpZfry384yVy5G4Z2EftTtilZeBT2FeLwKSdcJEIJZ0H9sIaPGVoLszvEtbf5VT3vaw
rWtEUOD36SDrr5uKYNrdp5NQt3OrGFrcGG4ouMhT4sOSHGhQIyI2QuyPYmCRjqbz1ezeMk8qaliW
ZbosW4wNxzDG7HF0fLUvblkhRJAri/mrnwWr/JrkFoivhocp2w+sD40EfoYnphQK0fmAcaW6qPEu
aRpM2xEznmf6wW7XHxWscF6NuOch4AENbC0IjeWeTEc/Mt6w+ngSS6Rg1cjaK1ia/hJKjENeO8/w
2QC9U3mX1Q+iHeC0zFzVn5kZxuiLqU3hWrg9d/7tw6ga8TA5F1viBx4TesplXiYDWb3Kpeti2KKW
0Z+aYW5nZEy8juEdR9XXRocP7oqEYuRtvkufSeU1QPkGzhrZG5CsfS5HAY1JMtdzeH9FIDBF8go8
FicCLva/ev9FTHTx0qRmMGthhJxsv+7yx5+FUwgiC9EIEGzeg22fq98JoC4En7qUiF9J/99f/vpn
hd+dGdZf8zWbwzJGe9p9zrKR1zb0e4FGBEnhRUEbI0E7R4tAJPINjY6ZGTqFaG/vKKwSMHGHPPT0
lOB/XdXl71Qf+VbylR03wI9uApPwQUCNaKu1Kp7wQra6VeA71uaa8mniUmzNNb9nF3uonbk86Fpx
K6qYd2WNWwr18AZ7PgNyjjWmIZl6AQNbpR7t2OajENRb8XTWOLcwT0Z5Uyo5AsMc/pRyvWx1fmVj
1gGi0A4N/TMDsZaDUrza8d0uTL9ZG5oVR/A2Il8C7w6zcVjUFfdjzqlKXhG2kALoVdEKYH50xnIn
9uRxcxTTK75hAFxXTS7ohr0laDFuzppAJpnow7/6l8Fq8qnjeDet2IyYQFLVzjimjRRsZbW4LJXx
8oa9Sn8DAU31WUPsSfC6fgT5T0/Ir37M3PQjpHZ5Hg4FQFKA5BlJ2YTUDIqEDUBrdENLpE/j6RmM
7nY/15C1PdFtOPn0or5vcj4JOKfMfPF7y3DRVUG3CBIaBTmEOxZPv3IIEFHhEUFWZ6MdEqYVeuG0
UaYzE9VtHA/3+Qctsf5jSeTiMeRVnTle12DUm1faWtUQjI13fcTDHiE6gwosF1rRBvMJqIClEvex
mZAyNwlhK5KRxlYH/gdjykEafn0jproK+EbJjXv2ZNl8i659/MecSd4e4qguyZ870jUm+FZmCVat
ccwHBsWptoArnaYl/GcEEDJ15zAdPZcOIqcYdLA74HLrA2ID7KoPqmLELPD2QVduexF4gDZG6iCq
bzW54bUTG6PxnW+9xwhaqn41Xfe/maadOVAZliBMclYRO+HF9RaT+hNX23B1HNTHHxavIu/osg/G
UNNecR+L8jBT2K1LGMc8BtNzABn/GjTwpZAY9NmPSLbpN4U7/Kf3poohTPVqeYU5DojlforJ9sBB
uFtdKrjwMpSskfiMTeW3kedf5cE2J/prsOmuo9N4Uvj2eWmd5Y/zG1MZllnF8vWHJxt+zclM00Z4
p/USlbaC47vbtojN7KOP8GDwwCyVC9WgspwazvuuRDc6vWGX9UjcRyNBo1Izc5/I//Sct6P9TV6G
EuZMpyntrvpElD+se2DnuLUI9gQUeXKF6de9/AKDwQV1oeWfb72RgHTJer4lMFCZHqlIMEd5cf0X
creLcsVqC/f/u8Jn3jVz6p4coUHaVXkow37FOV6ep9iz+ZvcEFUjK2whX/QuxAUxGrRiUyKGxKE0
wttGhmwe3udlCsD6/KS3AYVnKBBTgTJneVpL+oK/8hTnLhyi6+kmIzgDu0ZYirDRpkblzQHy0Lyd
Pn3J8TVVuJo+VA0bLU0PJGWFcmWHjHNpk+q62BpYT36+W7TuEyIsl80G8a52nlEX3d298jHhx9r6
HLYt8FeCU+WXruynTSP0NslcDDpQsjMYkBRQTp3OOkjrdHYyHUU+K7hR5zFm1Fvcu1B/yVGqpbHE
abJURPqzbR9pIOL3wZ9vWrz/R0+Czy/Ycvy4FiolROosr9L01KK2NkX74wGFohGWdjoRbDUJwjYi
qkKbf643RgkR626OVqRxwyn3MxeHhQS2MK7oW7I8KusDEOKK5KIuqBAFr1fiDqbUkTfMmP2LJw+t
+AYvQfm/+MuYvzZtDCq4gFDChqcyyNoFJeXnID3dSzCa09ujgf6fLuVHRUogbCG+ylGSXJZsv75W
KxyzdZxG0PrE5sHR90+IgtedA0F+cX6dMNCl5NBsvxLmXwZCajEj7kGBliIkNvivXEI9M2Mkv6jw
jLK2ldlzPcZ0xAywLhJXldLXh7FQ28a0jWVu62ccBCFAOaoU0GrV6qyeWka73DlgtgvTpYPbS4bn
uRXjIXBHDVB+tL3QvsP8WjQ8anZfpJo4ab7eBneZQq7dCPdU3VOiKbh5p9AFhe85rrthgRfCy9+R
KQuznQld9raLu6PSmV6ImjhmjT+c70h9Wtu5t2tQORKp3g4imkJThJtwbwuIQZdzgKCZJYqXacaX
Pni4v0ZGGJTkIckRTOJFgzgt64t4J+E+Aqvx43ynmGw0bJPWF3Ffyf1r8i0bYt6940sL4cmuU/TI
omcToRxBSxjYXb5g7iZpNtqBFn+rbSwsYe90TEgP5ORlMC6vhk25o88STnCOuczu4T5UvlIGU8+D
ZFhAr10jpDbakSnZc4otNyzV8sDBiUduiSQQzXZ3kfnujBfgATvrOKdiWzDo19h/vBx+bFkfdiRM
3nma12nJ8o9khJmlywiF7zydYj3/TqUyFIDImfH4lePnUpYxtKwUrcok0ynG+5FyXHCsCa1+KSKU
Hmir7oZVij1YXgYwIr9ysKSFPJ+mEnN+bJd2L4eZk2cjRL027owaEgjdCp5+q4k4AoLyA8iqj9tT
g6kxlIWYXN/h26Ao/fZ8fwbS83aZ7Doa6QC8HZBmYPIZUfPHSgJvcRKphXU0kw5Q/GqDekQMvQIZ
ZWAPQQ657o3CpPnLvAD1EmMQF1OD1N0PSzvhgYMYCi0+vnLslvcnmrQYtKXoDxZxkbfsZr3xmfR0
E0t2mXCspMnDgsSTI30yNYbJHMAjwvaKUUw1yUM4LS2wstTAtYfARpX7TzWYkEDgzU+b7B5os3HM
oPaoVm4KmxWpxssHuzxg5jX9LYkNZ9RPllsumjOZWduWQT5fVLKRSw8tl470m0Q02Vyz1sYMXVuh
0TS0KOTzhFoctzENyk/MS/2IKE9m9q/asiWuS5u0Y2aJzkFr0n0/boF9G/zZIFARFraGlf6QTQ0/
HLdqD+2uLKIAs0MRi81eaxmXK9TnJFeNuJRBFx1xSMfhiKCVrPDi0yaOFBO79qyNPXpgcrAhCZph
kuuVWQWp4ziV0boQAY/cC5/09czIcvNfw+EVoCzVVzlUjaDnefuFikPf3/MXLu1djdQGjhf6KULm
56Njguu9QucgAeSqAtNbSISKqP7MqtWyeeI9eM19fpBTMyXxvNJiTmIhHRdq3xlKQlky/zbvvo3j
CcH9P25H+oozPqCvKK11k3DMKZs+6YhWUyaVjNXgh6vG8T8W/BUHo2vZ4toxosv4Ozm7bX/jV3aO
8HZqwNlFdUgloLiq47RoF2t5SYyIITvcSYDx6I2bLDE2B4uU1gsjlk7fn+r1/S2TgGHuGo17EaQX
XVZB8A1HsjlM8eUyF+Pw7pa4v/FRqVZc2UZLcljzy4GzCR2ThCpcKZuJZLGC0clIHynQbl8q2MOw
jKg134Rm+e5BxN4UqD+kBLDGEGDqK+Xiyd+PB37MvhVeOvaejMOKKsYlCwwSeeZh8n8hMaO+lPql
ngi+aGdW4DzoLcTOkG7EuOoH7roODoR9e2Ww6LR/vE0C7EpI2wS+c42KU5fTT/Ulg0UOn1a6wnH5
aooreBEKhHVzU7pDQ4wHpBomeBDycagR5MX4T+JkJ3XYCkUDnRlMawFrxJOJ3bW99dNxFnI40p1B
C0SJOaIvRzHukoS0kgzRdm5R8BNmQB6hHT57lOAv0aW+El2S9nUGkZRlyVCqOrNAgZti0vopIOhu
6TICjSuN05CTytj9OSK1c+M6usjBX6xtPXtXkklqfX8pzi/W5IOtPUQD9jWhZrEBPmLlNtm15zzQ
WuJvqVt7Z8EcYbVcoToi2IIgX2iXxyAyzrbx8PekMi2xLDQK2sfKLbOCqoSch+I4Z9ozwx0uktt7
bx8PWVCyPeKwwya3rFu+NXSL0fSNbuY3wxV9/59oM1914s9+6IrX7zDB2B2RzX1zmE6z6IK4QeIS
zG2QpV5cU6pwboaHwXgT9G/gnN2wAqaKnFMQsq5LXQ1zAXrZleVyJZ0AT5XGTgePcFAYebJp1vHP
9wNzbunerkp+RBt7OikXJKaq4qYlxSJlKpb7OHWuwNmD6/6bNxUVi1gPhPDdrQKCzymCng4RD9c+
LvWN6wwEeesAmfZmUnQA4/IqozCTsCN5m6uMjspmVIskHn7XRKvgh+X9XPnaAdVk1Fd/mayBahSl
CuwStafeAthrYESbAY/sQV339cqAVwSvyb+F+mJVCm2LQ/JQEQB33SbBSAU3JMO6eh5YCFvvvdya
Yn2g2/GXBZTelnfVFw7uI3WYHR5c/F46kdumTFN1NvNgUk+2KcAxhtgHPQw0DwBP8nCGXGvAykCT
irblrkdPPv1SQ8Ecd8Qh3xmJkPEjuThlVF1e2aV6NX5U83k6r8UFeoVUJROdsjVGX20ybA33qrkA
/tmjpt1hcPlgTQvl4yqZv3Hbq0GRGFZ7ElfP2rLvxBzVK6A0jMUMjEW6XpRY1eOkc1EnEgd8gM1y
PlVK5rAVRfR39kBv67T3DSJCqXo/tD93FGCe/1W7YQzL5NmvjI1Qfuq9s/RFbW+azvdCpJgdhVx8
T3oVX6geXsPMqo/bj2OP05Kyj2/RsKpDnht3wUIFH4fOGMKIkQ8J6VVdE5O3F50uSCwF0Og3FZ+y
85vhWKZZytIaZE9LqgNV0PS2nh5SQ/hJa2H+tpP54QNnitRfL2OFY2ClbksOeEkM4OlPC6lDw1X1
AjbOG5zkyMWRrF4dhkJda1O1wic5LBk9kLo4vtaFUPf1JjLVRaHJvhyOdsFRvkdB98YlwBsKCnIv
qnIPItfsUBUk3Y8EmYKj7ivGcZiUMEiP18F083V/nfN9Lj9kVtvzEAte0LkM5cQGE+Jm/4akN/Av
HsZc2JLpKWyKvxqjy0cJNm+lZSIRvVbG7rzMRAaP3EQNCU4SZMYht6Y1mU0eXSb2/iKEgsA5N96H
1UufyAO3cPvvd1yHJZcM22GPEM4PTV2gQVk58CawJZ3sOiLQUVVsQT94r5eUqTgS7uWxebvR0DMk
NWOLJksJa3FtkqOAevUtCMUoIn7b1PEJu2iY2iZZrW5Kvzvu3AaqQpnGDY3hShIJF/P3n0M+avdD
4zXMya8ZGxy6ws1y23eYJXV2FMEl86dVeGiUUnFhdcgloFVzunnGon6Scb1yCcLAyj3vKp2hZGe+
XcLW21uDj+0sKORIpBSl/wBuUcVLxrDUAOK9ykFa1/bFpl6vFTkrJfS7Gue65MeBF2zN4FexncQh
f86LOFRqmdY+6iJlvtg8T+0+T472aeg5s3nPIqkC+q1xnE6tmYQ4tTQ2EoPGiPGG2mLdg8Io5MFj
KS3Y7KCp/U9m/NhgfLKHHa/W3HzX56IvWL60MhOUC0YEZqTQfVVblQ0bFOG46B/PgwaKccTHp0aZ
bKEfl7hVgiV83j1EuJHRyOPwKXgqRkJIJMfDGzlTQiu94erUZgeKVt9batLgytRd3bbqA5G/+Ohp
5lAXzD1iZYMBi7m4zDK6PamSyIatEQQwspG5czi6cCky4MN7xEzdZxZlCdezsWbKyG86KhReO0r1
u+ZpO+pXrHMOz2Kf3BWJZVYrN7hhLJs1gYz9tKB9syfTE9L/5KzfOVr66kxMZtWKRhzDJ9U7xLHo
+oxHUv90I9rscRnzJ3tiF4cI0ebPqnEeMlZZf0xjLQsJxgiQb5yfytO73Fa8KNzhKIKjri687Bhx
TbSrQ9l51owMkLnB3KFHt7ADEsJSlDHw551JrkJRHZt1G+s/nICWWwJVGQc57wIBUhTAi5sHmWy0
rzuhY5IQ7Nr+V1g1od/QLODZ29wL5JbNyk5C3rIxuseINd1wKAjKhth/o43/9OVGBSnl7pYJSAaP
KvUHMYtC7RVNpLX2RiX0n9Wkd6K16FodCLj7BPSd/hXVMkWkS3oPXtMEjhv0vxl7RxdD0jwqSUAO
JUI/Nn+xe/vfr5Tzomag0bECgH+svFy5E1SycjIPkiB9rtzdovPO9nL5xMht291I6gSxMG9qucBm
O1Uepz4K4f5PcbcbOdnat4gIxJkacrsWV/2IETW6fxgoKLjBX7Wt9w8qAs6YzfBM43SlnVjGq3cy
N64hcYOtsvZTAcZBoSGInD6UfElT71Feefr0l92TuIWA/CXdntYbS/jJFVaEoUh/CkJY5jCpFIg+
iK/iJ4oZJ1QfgcHoEWT37qLRx5RlTdtGZejMjdYT+rpvaMH/TTDp8ZuuWXzOfssnz1JJ24Dz/unQ
kyU+vXudwh7OLyl6FA8swnqcJ1PDjf0BCLvXfBEeF09hUWqPblouBD0QEl2IvZcrLGgsAwQv5x8u
89zKx2LyEND8savtodV5NXYiHg+DO+1hGOkKOyQwMmwjWxuHK1p9+GQohlRBefAWZDz4pi6bH6h1
HG99sn5gW4snU//T7bcYQz8fn4MlUCWu9XevPm4OfYqobGnxJisVyJMooce0OOqlpBOJtynqpmuN
Y5NFz5EE4kcNQMsit215U12/NL8PbdOlUghb3rOnTwdKsjKzJ4Sd8iennVLgnZ00yzWzv2bm8PEO
rPIaGoS7DuvvpjNtrYNJScL6f2/sNkOjdCM5xLYE5atqoIiy+BW0pvmQJxCwtAT/MaKjZ6EYeUSz
aYNW+6Fe2C+PpVIdZmR9wExD5y/7uO0SSELOLB3s08yW2zrGz0GmXkIecXWPIEc4VdXVW08eUEuf
j+/80+ky2M0cT/yanWaEK8Ziyp4xlBiy4U3V623R1xTIrpozp99ridicuOgQnXFNRfpx54f+ISn8
NE1ror7232+HsqeM+KalAoxajq6XOArOTIye8E2SOLp5Yz7Qo+ykY154DO0zcOzOvXFbiTUnyuun
LiKezEIXCMkf5QaiBq5N5v2CFSkog2dJA9O3jRZfkYh85sa1EDuwayWeKenxTH9Q1OJxDFVSnBtK
EnptZCkZlEOlieWtuFKnbd8IUEVqZXk6Ht+jGzVvkthvoQkeXBzVuV1HYS+K0qL0pOZNIO64TtFi
3rhM+0D0ic2+bEPd7R5OtfkkFL35HHgvY6koqGykdjxAyz8yK3h7AswUJe3To7GujwzXXNQaqnF0
RoTuqhXU5ZsOg3kgY5me5SYhoWGoD8W+YvLM8swGdMJe/vxG+9dSomUS26J0RZAm6UpT1PiwzAg/
s69WJQ6ZG/kmF6i9EWV+FgvDpyS49/88jpzzLiO9biIGAoHnSFRGOl7yL34AHhCzNfHCBla03HAs
f2a44MiVD+l6Y70efXhDDAFZ/dfCyiQGiAxzNyYr5dZUe5Q1n3lv6U0Duvz0leLDmrSe/dxXLIEj
RFLCjxOcHFjEDkEmVkRdyqnncbEVKY5OyURS7+mFeV8qyqXeyAMkyCHAPnl46zW5N9AYx5h5XbvW
Y9tpDTaqbUz1igD/dY7X+7y32he58iYMSuaE9llWSX0Y8IR4iRe5v5W/O6bgklwu71xdoA0Cd9oc
wiBuetq9/PaH5+kR77v1y/ic+6jdJojPuCFz/FeL45Hn3cBJe5fdVC4VqZe8EjujayQQayosL+4d
fwqkOv5ZoE107Kux6+Rs3QmIbtjDqsYds9aITnsyl9/zhrp+IQuh7mynlIetzBGAD37Ll7IbIh8H
9oQK93ZSWCnJVlRvbK/NzypW1U4FXMmBBAgfbJzZhD0AHk6JHPQkabtTdXOqpQ6E9F3gCOtAZzto
M4/7AT6Jd4jLYAnLiijwpnm7SkkAdzweVcTaGfR0bRgpmRet/is0ans/5UCbktlHnDDdHKK74bM5
YmzJOYOb9aeBVOBTUI3xAbzo85ma+KS7/fZ6NkLTIGsh2HHwrO777K5nuyJwln5eWblK8eq8KXNB
tkpnGKcc0j+L2lvblGkfa3c0wDwlGgGy9vPdM7MuNSIC4TfTrWKYXAPYrQifbHUlnraFunhXjRqD
tytAHns2bR4sdGs/ptbiNUlX6KX4Y9gYkA3HglCIxWk0ZoQ9RNbaVd/GRmtvsZBFkL+igvs7UsWp
v0e69l3xhYLFs0hsBW0lq4+7HEXLWlT/jtArjSS0KxM2QXWv1tEXehsGIElQxbsAaHLyynsh0VEp
ZwNGbRRtaOlc/xM3MaIP3ETrpZfDYe9XrqtInp9Mc/D4gkP4D9raxniFf+arK294jVLBe4IGs09u
mqKMd2FCbjrkflF0cxHfYpjyytFcEz75CPAwJcn4d6eJ+Pn9WZpyMWT2uj9nQUnSvE/OAKY+ehUi
HnQumRP6HH7irD1xC8AIMrBorr89g8P99eirYxSEQjCxot7Mkootn7S1WbbZvMxwAchA7F5RWDbc
6wu2Vzr8+T5BDmXiPg5lX8vCsVRjjPtX+uyqrSbligb8hSi052lNe1vA2SprPPWQDjZFHo8Pd4DO
RWzvdnK0sXzwr2ugf17qTB/G3YYP7McGhU0x7B+ULIGEuzroPfRb1gOBeX6WP4KYmRMYZnivFQp6
UIq5bQjyip7EbGmut2fwqMema/jfpfZ5ONfDXEjgxPtolm28lgGuQK5JavNCabgTS5GxQKIwfegH
WDBpgwW16TU3rSCGhyRBaC3m2yQzdrqjsqRSbADvjO6SiTVqYRp0v02IWaEkqp15nQv6H1SA72ze
GgjOnvb86VJSvFgh1QNUHl8HHTP09/eqjWLxV66+mqvER2NL7dQXLEq5qWU8XDhImpdxc0DRViXf
UawlFq3GgnY9mDKSw0b1Y6aDAPjzWaImb3iBMOU/6F05jHsao+e84twwTSaKtVqdVblVUEqI/F9d
quR3nkTpRQOS1SKZ60ULj7kJeLZbmy3fC4eog8JFHOSNuUINsxBvpdPgVNwqHhreipPiMZMvUFCD
l+wTCmpd+wUeaDNbUfZdZ3/jcbscfstEwkD+e0ciPtoQqwNA0w+U3p3JfAEiW4kU6pBstm9wuY1S
uB5o5uoy8BUxErlIKBwNOS0ycefxy5O377gzaj7yUUQm9GpU7/qCJYNuh9T5B3StDLvqj+R8w1cd
xyTN9yjFkPi6hgPjK4wjSgIXmqNl/QuMHGvo98gnMNZoHeuoBFEG9HBapUB1AFZtuvIfn1ANDmIi
f9x5O+jJUWKFOOFel9MIUUYw6dmGNwh5waUn/peOKyWI9ScK4YNZ9cXEODBoiQ7nhz6BXVVBxXjr
915k5v6DXjDLSlDSOyWBlzcifL+/K0qcM9t77vqwnQVKo+KfhTN2B8JVOPG9sk20Y/y0fD8sH0lX
sZUaj3FcIy9uPNL5f/heMcyfni38F2zMbcJdZPogEVQFUPpw3A0BB4dtKNsxTeMmxt0kA4WOvGGg
YjG+lreNzdA411vNlMGsCUSEqGcIBS71T/APGca8rMZST5GauZoyPalC3bxGS/qMlnfmNNzYy35T
KNHKGifg5qs95EW0X1X03hbejW2OrlB3lVnujFaYVkBURcv3GXtK81gK23mJRyuAuhnNftfzb2gs
pjESAWXxUEMsu9GfwQQ/+t9Wq52dGLV2Z/pJWTlOvCp+qpfqm6XphLchJrCrMaOEuje8JMeSOH+Y
/2RQRqFHBzo8NOZOD3QRiWB4DK6cTuC6eXDZ4gEDSt1C7Nstv5cC6tD6lpqiQkKpcENDDntNEPum
GwjltpjCicULBTjKlJxa8q17pAm8Z1XlP2rDN4Qp+pm6Fi84LNqqsyJflbKXK1rsL/YW7+EHYlq+
VvTa1wtLhaFe791N2hgM0Qkx7RfRJqc2TS96z+JhKJ84TQE319+/IvAk55FKDLeD0f0gyNq+qeXo
gX4xWAe8nptTUoJn9P1xaX316KhbFyrwJ3892PJb6pWYqzH6AXr01usHeGVM0yEaySPAWiFPuQ4p
KpKwrZWHQdg1D8lFuTd1dyVf4RdrYvrPb/NmUAf4am0cPw6tm0VSuu98iUhDIflrKvgM3b9IJIcv
niOdArMq2xXzBjKcunGXaldXsR0+RT5ciLoH2WF3KK/92M+GGonZIKAvm1aoP+RF/otPrM/zE9sf
EUhZ/gSfmRecg08LERTXWlZuRrtqjx2vBrtsrBE1SgMSv5qaQzsC5hjT/XrjYxjFJ9vVWgq/c9eJ
oxTI/9p3Xky+UJ/vsYKCr/3d+HXGsQj7JjQzZ3cxDZrC/3hXAFAM5prpv1gkdajtMzDEULle/YSu
jtDvIcGAaqg8QXrxOD6zkNxTbhuGGUgyRph3Ut9N0nN0PT131Pkb0NMFAyQO/tIBfNOVRIN2nL5l
aMRyNPV+AYQ+zdv6SZJe000qmkMA6wb+/MyFJF2Fusx0zBD4TfSnk35ZrgtjPvQzrNcpyYLRR9gO
io0EsSGBl1m6HxH7yNecKcQ+ofRbZDJIfOf3TkocD/Y1RjB3udCzTgQFE99jo4vJo99Qe3kNkDhf
UVMM3A38+uf3F4yYYZCL+Ppm3gMVa2UzNV9mgdbejafG8+31mU5Dc29ySl7JZplrqRBDtJk2rvwm
adPTEEEe6DaopJUEX3IvH/zH1jzXfxkREAKUW0oZy5FhSTL0y0LY3XwL6gD5f6VC3seQV7zhUqiZ
3EhoZd+g6BT3Ll6FtM1nGkDBP+YhNO5fH2PnDWq6oa9JDYI+PtzkP8ZKr7CUEv9dVd3vIiLNZWOP
fYn3MM5+cs5dy2Us3e/31r1B83wNh3+Vp9pch/Mj9rqoj4rsYea9OCtkQAWDhhr0T315NY8C3zuJ
+1Sk5EGuQ/hgDWPK3TmeY000paMJc9t372klux3soxpi+JRJJXveZEEATx4IRrcbPjP4ahrY02RJ
L+Jpx2CEsS8aqrxkJSb3oT+co5/VsN8VoTanWt/LL0by1A80U+z+V6n0ip23AUZATUXXkJtKWDhO
T68C8jixWpsP40d2N+TKiaBrGjqPmZki+pd1FamyHOgU1DxV2qwiOrH94oP14m5BP5w2Gk0cSdq1
wl1uWw9DVS1PDmlEk9vcLkSK5YiyJB/+dI0m5TLruZjZ6ZwoD71FU791b0H0l3DFirYwCoqE7tGi
2HG/MKSaM6XtltewvdteUwcsnLN8ALcMUlMnNRLkqyS18nIQPSL0+AQZcvDAOYR5CIKTVTgOgT1n
LzCE5psoIQRwSqFOtAfdYaHY7+8Hzi9/ky+CIYCeu+IaE9uLg0IRK/nLZiQcIgLittNy7BrRv/qJ
+sKoNT6gSFXJJEyEov/z3XcoEWEyydcC5Q6aJor2mes7irliZxr5ufzj87yHe4MiUs4UMf/KVfZX
TmNEogk/q4Ufv4bS+pZtH55IWrqjeFrGCk1sOr4Ix9HIosyyYU5PoyYd9CggaBs+eKizNKE+s202
ROwP+xECJUOrFvXTDaNrychwsS/dMRste9QrJdPbJSv+nsi9gBi8P/U/HF2cGkEq1Y3JZoPINBS8
p8HSQtTvrZLjUqNLKLBou/K4lFk6eBqsj8+L16+W+wqIvEFpZWvpuH5ZFsiI37eIaKD1f7mbCC7e
fVxx3ll4TsASLL2jxFOpSLK1nrJ/3Hp8Yzc8bH5B6tl92+Q6asQZIvq4teM0KDV+uyoPKhsZviwS
S+d+s/K2hiFod/CcS1+WbnaKF5Ra7S5uXpdxAq7Sf/R5oHt2D/LWq3QJU4ndjb88ddWT0KtJQwIN
yPCCmGQbXeaRZfqm+DWz272PeD+MmXjOAT1WAGs1xJRZ9YBLgeeatvsAZUqMDjSGGsMj0d9z0QrQ
nDYtZxlxrUFJO/whpv0NCWGeTm87Fud84/s0s9jxeu8rIkh8XN5nHACS56WdwtAtIQqhyvrNasuF
knuog1OdvOkiwbzJI+oUllw2xiYNZcATiKja7lpaRfb5DrTrJgAMoImspbdPrb+9QewVKag0CTSI
Ubtoq0bIHX9i2rQfGDrCdgehJrtkH5GERnfsigQR0QnCHqw44/Ge9LsD+FxUbRc/lDD1ACXR4oQ1
Z55JllJ77lwaiqWgsMFkC6eoho48SCjfRuR3S51LKmw02naUjL43BEylOflO957kbL4UNG7F/Hoc
K97yyTrmBDsoKwm4idwTiRJ0i6xPDUJaFgDm0rPQ99l+GdOj3hez3E5QtIgSOijE4iVPxtrN/7W4
dypqP0Tspv00wsg9jADKJ7akHbKZKJkTN/Fq1ZynhGrGmx1ZdKV2cIJajmwokqAXum40RE03dWEy
Ruxww5Ufv2EffO/1ZIOK/Wk8AXyRSoD6ka9eR6ANBh3oQBSRDNO1+s7Ac/LATAWqunUrYzKMIPFc
aFyB9Qgw0FjjfCh4QPTNsDQT0vxDbna8ldy3o7pHK1vavrapPYv6JGkb0wP4KOH54txq3L+TieDr
WRTcwExYRuXmVR4N2wf44j3hGflS6o/MVu7L/avvFDkLVU7Ynbw4U5Uh5RSMzbp0rJwDXXMuaLxU
JEriM0IV8ddf9OMYjLxKkVUB6J4ulHh7ZUPpqWYEe9EfleDGCqyQOplIvG343aJ1seF1wuye73/T
0VpW1q4kohXSfNqZFfhuR+u5CsfI8kibcnpwE2f/oRNujGxGXV56E6miKG3myxN7a2bDw4neXLg+
7gxGAGL9sVfZTeTTzA8mw6U5DeJjDtjSyaHbG4Smjv7ujBTJhF2Mw7hPNy/wZl94/Raxi8jIym+j
9TQRH2w4oGko3/4WEGmkhO3zLztctmV07ayScJ8grKuOXa5idlyPsRBewbC72pHx1YdSOSzh/HUh
uZx9BRgiQx5xDXtdobYEqcfpuw5h1+BgK3L+0iMc963McJRfj8GxiPODXrGSZeziTC6iwnHdZONb
VTgx/UypkU1KDvf2w3ejV2k7900Eo560SvY0tWJdyECqo58vz89lNTHjMVejLekc3Sm81gNEcg2S
Ysd8nRtxR7vvYJwdFpPmWw9c/BhHFzH5HQZCpe0OG5ZTdyB2gIvkcCv3iQIlJwCiAa+l8csWj/uZ
Eb9h9pl4ql2thc2nDFTbL/+z7vZIUdVb6tOm7k7HUDYwNBg3vAcDMpF4rYmPdIrPzC7EEzs/H4jN
i68bMKGAia1y7bHoPmbtkkBjuimryplLjdy7CuCc9n58MzMciCQNHr73NM3H33FKuMSKWiw5J1Ha
ZVNrvRwFm4BpdUmkkBPuOIv0mno5EPNC0DMk3cAqZMgjzqTac2a6VEqEP9QW5/H9R3EMsSPdHe+X
+F60EZ9Yhazr/gmH/+D4A6vABgU+X7g5CgDmoU3A6BLyfxOvsvYh33RuHHpI/toer4d/cJnnT5jk
DHxuJcNpoceR0mIHMMLDi1dCtKISUE7K82fFqn1tm1eMiNuQdGj2GL/U8DDIwZ0OiuPvPnINrcn0
N2QXifp4pciRFSaN/ZZi5JBVG5hKhvaAZVkf8beLTa7SngDFFI/3Qk7O6i/deakcPb2foT/MuUB8
Cev4D0xKnb/S5NWODuXqgxV4s6NwZwuDcalPJevRJwOrgiPT69kjyj5joEIXnYFduC58biteYdtU
UuWuGXohUbBnw7hsjkmgZ5I8lgqU5G9XBRx1EgqVuRJaov7Y0mxD+1LRfsY7IkkS8e8/8swbCyYk
X8ihxmxvKebjVr6GQu9uoPvwgGSCNn/OsmYdcopm/LOjWH/BNBFo/2RHwQUegOiVQhLUWvnibRFd
wN337kgN+yTPjUQbSYg+OFoWl1I9nuwMkR9kMq2q4ZDKlKKo+/NAepjqDGNwajDyXUmHu9dtMvMe
PcJacc3UR5KxSteI5BB5AL17MKBtQLGOpGihDvYGnfmIEm5hrHn6qsllZFTeqVISqsKsf9imjz87
WulkFtwMzmqBnUXA7fyw5vxhpXJ5JzFzzZytGdQjO9FreAfFvEXFDUisgoS0fqAg+XkClShnGJQ7
guzkZ4aBgGFHh+0GOuSLvbdHY8ZPJmxE/Ed+EORQeb5kq7RHT3uc5kAufhQtb2BgBXBCKR7ugw+h
U/5snwDFvgb7EdLqi4QKp3lxBHrFP1EUEgE2EAxcJTQxf+rq3wcfDsaRZTX2M95JkjX38D2XT4jC
49zMHB9/1Hr4r3bzWejje9oSUuzY0IQbQT1HlNZQjePeJgTs7lJP5J4a1jZj5kJFCXxptQlXWa/w
8kAvQC5+M924PXQRVDJlPQzxBLzzR2fjo61cTF7DJ0WqLxCLfaFwhl2ku4iOmb86//vGKDTBPQ8/
8tPA71bJi14n72/1gtKUaGei7fH7ieobhPKwAyBS9y9aFB7TzUoPGdxi5JN7g8v44h74bg0foFXO
22KGKtOf71L8fsN+0A8G4Ma9AZmlZrPSsVbkwYRf9qI80pJ6QcDTfUqx/dNChbKnCZRpAdpXOwBb
vYsST+/9ueUe8SJQayCm3IuFv4B1H56Lt2UA5i0nlYqpCiSnRcwASHrQwQs+qUIVS2ZY0+bl3Wcb
FsE9Vw0xcHZdl1QavUhHh7rj1KLI9fGX3D8t/R8K+FcjwYCSSDbJZoFGam33zEthwKhtjLPHBroz
vhzCAWgmffi1RjSTMCcgWGzmAn5Xuy4COTpdC/ug0nWb7JQc9rY5CQrnbZFFRWreiC0EuvXhRgWy
b/jVRvSbnfppHM+25g/FHDgugsEtfM6AuTtBarWGrvvl8ZuIiRxak98wBBd5cj3w05ePst8mYC8k
odJ6mcfWOH0HNPtzRcSZkJv43BaHsVO/eJRwWaxLXcujrDAIQjafeWbLbVYCjuMThhByu9kL1ef0
hXBK3QwYm85n3nTixZjjhxFXzri+nf0/JnLUQPUODuYY8ELc2ZEkq1++Y+Fc690wsV2l9Eyfuff9
Dh5L7nEWNgmAXHx5ydJWRk+l9ZSXFCDR7RL3I7lWYTC9+VoFGxWSE/hikzOACIv7vGiOwoFtSeiR
YxPSWIiAReheWZgKLYR6mr6Oqfy/4LFEDR6r2yrap1yTTPL3SMgFSaLO7qkHdPwE/moKSV7SDGxR
u9SJmcYJNws3RALWuIqo6ZO7jKqFMFtbjYes1RxnAsyz2FR/mQdqWWk3zjZPbavfYZhNVBFHwdK6
OFWoC+zAxxIMiOxBgl0ykWBTVFPAOp7YkUXfj0icteyziDI5oTIoiCbKUR3w5ShU5z1LP9tFWLHY
1WR6BEUc3iMas7X0Dk7N9QyDI9iXD6rxU7pzqPsrmvYe/NyGpzHCjiUMuJQRiotdcX3jNq4/K4Fd
ZWmiIAzsvEykmrWV0x7z3PoPHtKFKymJffETUHIqFrgUp184RQ9Xxl5Bqq7o624ynl+gQrGqL8dx
SOWAeyQVFqBPZ1VAj+Sx2JQ9CgG3bD8Irm0IL44cGwnEdc2QeX1YftQ43ENcft7W40GEjTKYsSFT
Vna/3wFcn2IThGXnVZVddXX+wIGfCsVbtJ75lWCGCH0UfezfX4/hpuwPM0ZLt3nA/HXmv47Zvj/2
1eIaMPtI3XpU0VKwJ7sANTwHkYOaFsYgYH+7q6DyPjM6RJyiRbmkIUp6fI/RWMR1hkmcaC9wBUqt
hBWu2LsiwCnBksF8Cxle3ewD6/ZLCK8Dyvmn/cXlQLMYMai32a4MWUbItiyInjcrCTyxjCgxHOHi
mhPRr6c4L6Ow696pcxqciKHEmRYCpax4CZorITSL3pvNI4poio1OP+0BuRiA7JzfekQ1hb39/P5O
gojVNHJ6zJRObw0VL+aA0X4YTrptUF/KiLf6L//pRScxfkm/w8ND2Oojxc5Eg8U3qXr8sNihNhdm
4P7bEZhbQk/+LSsIYXESH0+wNqXsxrB2UtbR67oNcMfMxwl+dkrxBYQDyogrskCaRNR3uDKt78up
4vR9FLc68J/sw4Np6eLnq5ebmUscmizojNtO2Z6hgZ3mF7vwy+PFf8yF0nzpn8CAKccZAagL3VrD
s66uMz474GVV1CbbO7yrNd2AGCTGbdP3FJI/0S3GUgfdrLenkFm4c2lHQpHkzIlj73sVS1sW0e+m
eoBENZLcNlH4FsaZvp6U2ZR0z+fBe1ZgZMlKMTgllPpnareCNcTP1/18dL52l+BPkI5Es45pN1sI
1XiFAQXAkMfXnllYv9mRP7cxTzf5Y0/efBem2eBeRHBHXwMEWS3W+poufDnnJnY5IM1Mh0XjeRHF
MryXx10VtXN1/kti5kgUeLw8QFk4th20scI1ILnG4a6qU8EdU+ggsPOwLCPxvw6G7Gf9SBBeTgZS
NDODmoHIfkJFBjCsvhKKfae+VUNnAp6jyV/Gs0Mg+8GmrFyevWg44b6SygYvUvBYApPdBK3XwMh1
Av57/6Bqsdf/kTuRBCbAN4ZiCk+hrQgR+4LZivAOhE3VNvSpJvH3fXBizKi8b3H/Dim7BLd0u4Jg
ZBbbsAtLePxUTs5/noPmOktnWilLwlAwyNRPu5vv7JhgtqpZE+M4cbjtZ0LA4ro2kQD211hABne+
DrteTnl1rv8/VRR7WCnP5h+oj15e7JDFtkgnz4x5cRsoU1LdLlArNycc7Y3PYpz0TOv6tNPMm4z3
XqteO+riJIaLDH4lBSe6m609wq2du5YRA03rLqH2qOoeVHjsh4b29+Ffi/Y2Xvb13h7UCATruOyV
HGrt7+eovU2tl4WiRqTRikcCrP8w2bnVpwo1KiuYMaEBL3qlCM5pLBrfB3cGSN3BNJ3TDM/+VqtE
MHelEBmIgNh5Ii1S1YapSSkWzSbBp5nEAj6rasBqyXU8pTarUpUqeWLzvyOi+CMJiE4oFlECewYG
VUHEFZZFUlnZ1P5LP43F+0up8sKnda8rCvSfK63cVLtxeXngxsZayREyi2A/oGxhK2ekczt3JhMx
mT/84ZD05k4XUEH/z9ule8+nv7ObGQDYjck2Hpjtfo3Ks5rfn5NiGM9jEnnCZGRnt9sZQxw/5hhT
FcKKKrXiVUXIsrGlwbOQKkhOk6E4ompcz3IPWL8HB3ELGJdye2LOURhw+6j68JshwY/UH9rJOZkF
uE5hzkkDOv0lgKIulrFGyDIlDyt9Xwv9oQ0jytHPVAs7Q4fOxD1vhMtAAr1FJ3QXSkiOBQlG5MmG
yoKOhSXvJLr/36LIgCCOD2SpX6lsh+vZ6vH5RkqYfCLPYdHpCQXNu64a+ogDDgyhGdQ/sLZkHozx
/vewBynQmSgOul+SKP3VQ/82jqkc5OK7Ej5LtUGqLvdz+KqzQACE9+/k9Gd05NEOTyGyUGgHYEMV
pqvzXOOQ0hjZSnV8mDfbudVQ7RYZwsh3HAjk00PxxUuQ3ds7qDMv/S3Lm+zC5Y+bNj97j69kHrhp
FbMEQtqE2aIPi0RYxgurwuH/x2qQteePZu6Vo8AV8IKpXn+mVvuGo4eLvIp0GubACqU8kH15FYjb
evmdqPDyrbZAaVpxHxbWyKZUPwa+o0kazBlYpDjVZ13z441p6a4Ih1Vmc/IZTq52R5PL9FQJQ1KE
hn+Lezck74rEnKrbUKh1qChgP0nY0ZHKi9Jv//ZOHKcfbNAhDfpAY4tgdQMo28+OxCVFWRYs4ePT
uAz7iuEWuiUFvJzkYG4FWnXPmhCKlWBO/XV4UYf+ZOIxCnwU4i5E5cOj/LCKdplUMRg5wYRRQ2qa
ZxQzQ5K5JloVBJ1zYpYXeZHLMWcuaSxj0pLMJuIxRuBKYWTVt42Z4YVLfG9J8ma+yICgkE+496Oi
RcuZMA33KkLdPROuUY7X9F5LQb7skO3XpiCcYfz40PL3iA/ixofsY9kQniFQF+CdHeUTGS+grjhB
F+KRBYv3cDK7fB6BsF9IE4eBEhr/oj6h4KMUledY0przEId1kNH1Ocgy+R/ma2xeN9oIjs33OPxe
a66k4eeuyePZ3W07VaC3/az8g3s0/pXCk+4A0bc6mg+q7vj2wuKonDQ9u+w8qJD8s7TvfkmzwVYM
afLaFMEeTbPvyZ5Ll6d/l9jx7FwgEwf3GV37bmxxRnT1WC+loMFtaR51WR78ld21AKqad5wAOo0V
x6l63VXfnZdb0aGJZ+/hJeP48a/AgAAYYWuWlmZ4vTC0RN9U0Kf+1ixw29zTYygqXqnReEkxYAXm
1/TioeqqYRF/79l28QU2QwGX4A6rSrqLawof07TbXVfXdAdvuSosry6r4mZ5fkuvS6Yl3XHVV8pC
uUbNwtOcBgAJN9FuMuQUd/MjsHrR8GWzfa4MY/VRjDWTWgxmRjZDpMIn+/W+U9o7RGqjwGtRGgFI
KmZZ1c/tO6R5wx7gARQsPvltI0jSbLsUHWEA2f9H9sm8CIDL6pcHS4ma9bTBNPH/yHA79X2hsy4a
loPVO/wkZmph/yKlaAiZEA0aIan4Cn8SghRnjgN6XGVYURFm7zv/pJfdXG25fz/uCmNDIXCi2v4e
EuURJojdnXE3GnOxKiWITwG6H4vlhol/bxQO70DI+tPiXn2igc0LrkkCuIj1V1tj98u/fV82IFuf
p6bBQ7VAHh4aWBkXroPyoyv7ufBYqMOHEil0Oth2a/tanRjWAqDOYTuRV5lqMP4NlCRaIq6TJMei
KFkM09WlraXc29PlxgI+R1edG9ageUzFCJT0/BCR6lsLBdK+qUkqN0a+KRJmMarlmrDqs7iiJMTU
fGF8LKqkPYRKuuIgglhr2OJqynzZT0uoJ+sXDSJhzcmU9aS2G9SPg5x2kFsMB8TP/wSPfjoDq84d
nirg5Lgp8rmm6UQOmL9rNJb3Se+x7yuWdwAMhQKORgfavKAlfpJv1e9PooZcHpR5aU6D5lqEFgMP
/p7FpijpXhbIpV1aEcCjU3vIRPrrjMs55fsDgMMfbFL8ek1h0j3PPXeHRUxUQseAL+c3LRIC2gEc
fahhR/IlKsyihOb4myEcXO/MySXolSVX0KHG6QjMQZa5kxUGeqQmogfxnkYqTk/evVxfC4BqCuzx
TpF/LUrRxwVJyVnri//DcYfpMls5cryWAJfHhOHSRIGOiSMAw7uWm1dB9taQwXPZc+O+xSAeEWFh
8DPmX/F96eIiEGla6BHRXlgKpdJ+7NHBQHJuP9imHNDJqNpQbIJDjGdNS3/SqvWXEkP/jNocq1D2
uqLJyHn+GdMY+nZLzgO6zD1dh+RQwQiaQk16lFykrPcqaJmiX4ZPR6IVOi2tFWg1L6Le6BGLfVEp
USQ1RPhg5faCgUpMmZRlj4MNaqycxJQ1VHdK3yJtUcKuOjUant5pGIxIG+B7hVoNB35hZwo3ALhr
SK1RcldLozu+b6X5f7FwDIVqJ8/piKcSci2rNR4DMTA/e7CDlNBSMXpfEmAui67APK9P+TCWcwmn
1qui2bdLWC2VTrYSteV+4HRP1K3Jw68HSHw9YdQiunc9ZXLrfUaZy3OK23X/AshbUyo92IUfHclW
rkhpQMe7QTLhB5Vroz5sBP/lFTsOGcemzL9kaOUW4/5DCPBGMgAMG/isOBdzDjp8EL78cs1wACQd
+6b61/YLfp/8MBIADzR9js7WDfjAOCvnwDltKgTsUT/Awsw7CpnAjTJUDaKj3/+GS450S34LNf4v
5MSoeADvKpOfABoBE/g/BNKwP48L71JuPi/o1JTn+Y7VDLUYNt7UCiveCncOpsUbwn/LympUlame
b0OoerkT/J3G+BXkm29E4O0vjZHYQbgthz3zLgUx4rR6TI47WG1ZKcgwIi3OILYNKWzcGcnIeReW
L1IafjkpYLvbYdPiivyJb9Gmrvi7VE2py/qaSHfMlzEB/igsXKn2KJ3J/Is/A1mclRj8sUonTjuQ
knU/V/TJvbQl8BsbbQTzNYJZ4AQBKfVUeEsKKhTHkOz071p1k09A7yq5V6NfcoOSTkmvVwj1zXjP
KuCIoB6lRN/muPf5+l0vdlvi34xOYee0OfGigyIAoJBs9KZR2vnSu4ZzVNRMvYrhe45kZQkZg5jJ
CRXabSoXNrMBZ58fuxNONgg6aFOPPcX/slIkx0V1dAGuQxOtBw+MbCEAEKczPcWkt8hwLrxoASOw
6fpWnoa1TeJ3lbox3Iw9wDPQpCJfyjjy9/CjSAiYGOzGk199rFaFcVYmGwraVQq5lfHYxsigf/up
G3dToElxrl5+f3XRnUG1MxunJ9bN7WEna1lZLW4lrkKntL86ASGKVksvUf8Uhi1YzIX5WppNaVrc
DanPn5dszWE9pbJUiW0zB5goXC8+RM4X/MqaZqFT6U7r3a86G+hjLqBqhc78iDJsfYjqTjWUHX10
QDJZgMDJ8ktady+HWb2i84TUHC1iPMyhNQlXxGbrUAtfeJn4EgEhV9Cn3Wy7w0AMStRYLzrpot1E
xVXA0BsBbR3P5TaCKEX0fX+Q8YexIpktZJDRlP6z2aJN0yueT1y+h1+t13xd9JaIdWuQZKedAnsN
sHtFByLLNgNRvnqueTMyi+qMV9LikeShuYmKIUeIpIw33+miywTTBoGhV9BLFP5JWJZoDYiFQrXW
DckJ+yu1w/hsNHQquIvt/F9lbmF6713nMzAQew/O/fa/xlZZRodY55mtE3x4DMfr/eAXx8nfhSfw
BICG33DhN7v2oXxfvukky2koL5hYS7Ss9yLHVJ0hyM6q/OfvxMaQ7rrTiGlmNIPeezrwpg7JOUhL
Dv76d57O/FozMqUybFw9qlzmJ82cmATfEJJlu+wV4F/8A/9T3od/Aiq/RbALjGx1MlXST3MOSXgq
zWiVIiShB/w9P8DBydCTZwCFIXzOfvf+LPv78flGpsf5Q9jDl2K2jd2pSoDzECTjAB+GgBQ4KgoL
sgHbstXYrKeNB/m1Ji/Yg/k15AwqlVli4vWe/20/9rBxnUVnEyFUVZfgrUxO84RTLI3/ifb+kxew
ZpXw0UQS0rSYMKc4lEVhyG67S0iOKzbIX17gmSYMS0HmPprjgK4sGq7muhFvkSCSAmJttBifyHgu
DtEHaD85D++ZYfzD26eCYATu2GnCn29ehIYQ2ShexnvwNuv7idQ/lbuZZgt6VFJreoy/dhb+ONU6
gdE4dcnySfqI0JUw/waee9HKAqKtXu0A/3SjohxaQ2srA7moQF1Cen0swqQWADVphSY+QL68+DiN
C9xP16PxJsOHNOlMC8SvJW9twWtMhy/+bY58Xs/3/33V4u2ughbolHJqUF6sV30LSVIVewmLhNoW
5SwFWCL+eG+2lQKqsXJpHxAUTFeJpcey8dAluNR7EJQp4iZSOqgx+N2wtX8v5YOT+IkPv78obcOo
xw0J+kNjlOVbtlIyL+OA4Lcprb1GxgvUyfjxQkLHAWFCHtZ1U3DrB+ALQ2pPzUrsCp2nJzWSQesj
x7elT4V3ZrN/R977Wm3IQiHuRy2KrHKuz9yBv77UZmVNnIrDcglWc9rZxNMOJP2/WN9dlWUtF0ty
FhD0NxygS2ZF4HHazZ4I3nBqQaf/HwJvugN5USl830K2Y/IQUhkeVwR9+6rHtRvHE/0DiENlHv33
x4kKTbswdLzh9Oj6FrS2AcqRZLhJpVqAvx59c0JiFv3HMwa0R+x98EWgSYoBZOk7GBtmd4rlpy/N
Ep8zSTccr2jxnmds9q40iVBkR7Kw/7s5nsFnp0Awa2ZoRraRD6Xwk++sW0Owrv3U5FbeGroP6qkL
ZBre06Bvrc1JRvaOTthcfBRFj5EJIawLDFPAJj8j5eX2kUCNvGZX05YhsbPXRGOdIdUrKqzNkciI
LdkwYaMhN+Uezw/ap6+89Uv4mSSXtL0V8r3Mzt3WgIPOakopUW8sJFltFvnBR0lIFbmutjyjxazO
kqW2X1kv6+c694BWutqK6VkUSZniQf7gQeqGtl3uypUqtlzSwMNTJVTHIRDXmVDkyzwiE4bvb2ba
sBxx8WCQ3iTBMAWXOEwnbk7ptOtpRO5VqZK3a48KzAOUqXiaC5QhHH7cWYAiqDmJ6D6DG5imlUCN
/32v9F5Z9tydQ8ivTdVKmoCfwDcXg2oVVh4eJj3HqwnxJWCgMCYSrv75gt++agg6tswHZo6l+DUp
noouLighhpz/Vcq/6u9QtN+P+eSkZBI6jVsVjrHebACyOXS8hJP48GVRq10s/l17iIqqOanzpRmp
A9TLQX2GNqp7U9RC1SpzYGmHPTAh70v6qTgxaEtd36NVWwZRd0J5snL5NdCEYmVTJycNlyrmdS0N
OtBynikL8etc7Hic+52WchMkMwSyZMjUmTtaOyDhlqjqdB89nGBiOu3sOxfpyUQ7puiMjB5UkwbB
fdEawtVC/enQr2dOYzeeiYRKoBWAdnS/EIWai3zDNZVB+fInDOjK7Y4ZbBbHE3DhiJOQ9IvYgfqL
UsgrYRBwnyXYpDYtFhiePj9/eAmeO3M0sFmvywhXgTPEXSmgjvPvlmQLm8jY39f0sjbXpsGAVdC3
S7kx/TVZ2oT2ja1iFCuxiSmDsfM9V+hBd0Su5UI8pGaBhSb1zi7XHPZAJZ8kRThGlw3ay68seTCo
JL4bosjCl2kYeVJJpvePWcQ2tNrSftJBfDsich3TjiEpVxExl9X82nAHMQSeykYzBFiox6mavS8U
gbnSYYurkJ8MybgQOLf26L3GHqPbCwUwfWE98CD4v4yjrg6fnIx1tkivrhEsgL7Gp0D2kSiOfnmh
wclXJTLk+zQXCKIDsKblQ9W4qXehLFAFXJU431P04FVgBFhbDW8DYPIYkv7z1TzrPdtvwqWt4AFm
7X5tMB1/78p+f2hnBNBJ15UNK1NA4VwHHnbye4rWCQrYBo5WgkwRu3AKYz6D1l7KMS4ojqP5NzE/
B0ZoCz3OQ0dKGun0X+TVsmroBzDhM93PLXxGX5TBXYQaN563qjpv0r75/pAZPFheNRBwkDX4Vz5m
PF6u4IWc/9fFXC8R379zjdV4sErgPuI057HcWKaWJ2DCj2ckBD3TwkvVrdOxH78kw9rjl+f6leub
YxmXEOFQBMWLp4t78HR3iq1UsA0j8A0bfjBtKYlTxEQX+EcVKeNawGQU37thGcTzcIkngG5sFjdK
Qc5Y8LzW5pDiQEybX6GAgecYGg0Zde85FM3bGfGVUxEReKuFi0RKsR6I/4zZwFh5jIdMSPmBtBQg
I+1Aocl4Cttn4M3GgMeLJnkGQ9kxZJzDG+sY0FGYzxsVHN9sK5sRfXlNPkYQn73weYA/ZPeUEfTI
lK7TPCEIM0I9lr/h2N/i+UA3le7/XLmXS1HGWGM74MJCtiV5kTr8dmEUbzIgjhicT7BvrHXFSj44
47tvodKv6KDD3flqC2+GKGrBP+oX30VA7TFTMJdJqeqzlB8DWauLCZeItYotsoQrez1aqM0yzzas
Y/Dox3HafMjP0Z3paXKzjT1P28LzYa1qv3asZhTjMDR5xjQaNeXp8OQaj+K+OAsxVIL8DS0yiw2y
ftrVKjAf/JKw8KQMw7t/edsxmGyLTOzisrGQUKy28uQJby+d7NffUNzhJ/X4D66FGypUAgE39VP9
nb+OXgvJAp8Zlns5CFF3Cv5OvvK8EFNtgLecMsaw31r0Hbv96+4/DOH+N8R3XaAClil58RPYSFlx
BlhsiTqddYZM6GTu8yP61hZ1SAlWwkwt9M/EyopazSTzpqhJYkKPk/4aLIiugmCOtILojm5qXhAA
aG5uCqGuP+HKAPmKhah1sU6aVOQL1vdWG+WT8nX0YFX89hif793fGE28fAOW9xWcdV5NE9W8oWZ3
/anOfAWph1sydXYsj1O8+Qv3B7nZjDrsSCCzlkwbv1I5fXuAsEB1VZPAc9xBf5sBPL1ZiWZxJj/I
XuGIysHr3XFe0EgYUQ0rbdAsV0tEj3yEoYMSsWfTIpLGfoOvfAIYrBwEQRJIcbmckrYROnt4fwKD
CnatEbIfZrOaZ9oE5lXZD4Va36gNPljnlw0RZiy7qYjaQKqrBGc9ylV+4mbIAAFFCYf+gTSVGeYJ
PRNrEk1qFSL9AsTRlM1KUCiBWebThZ0zqKaJ38xOrhEFrMsS9t5d8URP12zvEaI+p5M4NcRvFD6f
ftiz/SHiqzPDnu2tz3BOhzcAngc5gKPA3ww8DqnPMcNkXuRjJ+JLOigQe04Q5kyuYXO4A+tS4Dbs
qUGBk7Tpp3j+IM9yqlyeWXE/hI0QYMi6ymBHdna0TlmiQR4vs/uIZh112TZvMOVj0iZbfjx6bmRw
dEYjysXyO0LqHk0s0ozjj1tldRpW29wtC8EP1/7eavgQLYMiueLxcxA2OE+2ZcPQxDnXiyyVm3fr
IOeJrXcGpz9NrN+udCuIB/dHmGcrkR5KEZlPP2D6XkBt0qobKkKcMMtg+TWSohHbeCnGuhKhebUF
wspO/eqZHiPm6L3g6cOodB7pQksyaz13iZvze/Poq6CAmvzRgTx/013jfdge14dswog1B8HPANCd
0Jw+r1GcABC36B0/rlFJhWG7ItdObRltqTwl2E5mhh1XGFn2xxJg4sOBeD/hYw1NFfIdVY/uOfJB
x6dJ7J6yfbHyFkKwvtSpbcsDxmsdq+5qTEeL/I6qJFAN2yz/K5k0yoW8oitB3pSrYLYaeoiiDzny
99/nWDyn5UoMRM7CeRobG6FlwKNSxK+LVAA6bbAkkEQTzab/eI4ou99pXM5UDnWQm7IjLMqZnDoz
f6k0kH04a6WeLpMZ3vURmyy2/V+oiDuUc60OR4KqXPSPyw0S7lckfKvyXliGT+d4Tk65VhEb2kvz
XS6U/APClXKGVCXu5VCIRFBLUfMnPilxSkDcnG/tqX1wTA/xVXFwM5SWJGfMTm2c2nWqzSjuzTjq
UgkqUaWVjceBbV1Z/cD193TvNXOLCK6r8x7YSb4jlwZpX0W5ULBZlArwaoHWDLRMEFGVRhWhANW9
UwBjK8Vjkn3fRmWf37tBsIi4dGnmwOBWsN33cqFBDlrIyQvjhQ5Q2dczlfmslFOJf4nF9KXkMwu6
TmG2sldzLtMUrfycwp6w2HDZnejXM1HslMlPm1gHjVpUqRG5KvzM38s29ZxW0NCfzaRqyo2sNTvi
lAJNGAMeciDn+JImyjheTu9GACa31TD23B3G/ggdjmP10hFl3toEUfotmUjXhGg7kxssnsjwF/3h
VIx8G5/To1ZMjYubpat6v2LsCkMeXyiOpRRAhRSCgIs1vMOk5x21s5aYLmuutYQ9hwyDnt63t1SQ
OHnqeXjNcfDPYpmwG58RFD4yrWy7mIPiDH1JqPYvrO+Gj+iVq0hzURoF/zV/5PZgbe/c6Oe6ARWe
ysBi0OSC1FmZcYkZLZ17y1tDZnJ99zG66lG97cDg0OAlY2CG13HT1uUlKsCDFTHSkNUkihNevh0/
HjaxK3Wy6TQ28vOgghYjedBuvivQywveaLNDLhuKpI0p1tw2aJY1xg2fil1bXePwaf6S5vnbIMnp
YRSovHCLjB7ERSEg34H/3Y4dgGJSod5g3xPRHI6eOfwNuunykh5nUE805l7RNHWRcQRDjL/Hl+nQ
hFuGo12jr0Fxw3B4wUlQlosu5mY6viUt2ywGjrZltX6idEA+p4TtWSjzbqdOWEifrEmUUccMi/Q2
FvzU+TdlYcKS/LGYMMXD+uTw5Pv54jIQI0jmnmJfmBXvwbJXvtk8+GtcHEE5KHVmrhypjXgej4Wn
00DM5otDj8i8E20U1x43c6Z+oRpR0vWfRyshYfEQ1sZ6pExkj5QD7ZwkiO3bXS3w2ktmmaOIzeM8
3BHdZRNKFmuuQq+qO/hMpwNBkfSLSDaKGy/LiLFQzRa4zLx9QG1b3dv9hPv4WX8fSKG8eDtPGgPu
0UFD3DTVS2nNxMYV0Le+XX5i5sVHcVskBl5ObBqlFchKodVHOahzMwFvUVqOf+9rNLA99C6TDaIz
iGOoWI9Xy+JvrBho+bXQxBc1pIrNiZzOwdaZdQWqYOUpKq6xqbH8eGOBBKg0PWuDRmv8g6k7RM3n
FyoJ2dTzkt+AqNh5yl67jfxtT7PfhQ81bdXXhycAgaXxx492Mw4TT111uChR5X75roOTs5Fk9sGv
8RY+jf6SHnvAFga5Sz9jRiWxZINtmGOaFDqxVnG3Aa5F01S9iGlvDwNo8Jvq1ldEM0C8bD3YIGFX
X9S+MBkH14zR7bLgy1OWOCpkAsulnA1l9ZJT23ByMbOUTqdcNxXUZibqkpkj3n8rnK50Jhq8YUgh
QvZEipCyysdruogg6ALUsWI/8oI958eqV4DGDCmUd57FtRBSEOQZFRddmuO1gVQR5VkATS+/59QQ
N8C54qIPKaGYbps9FVMZLCTPqWQRbhv6Y5lcykSMHkO/9kJ410ZsfKn8LzWv+ZFyHk9XC6g0OMDf
EzDnKQAEGYOAV6F+TiSur5FSLJsGeW/FPbsUYP7SEeNEaIrKAOUeApGGjnwTrHNWjx/sSeX+a4NZ
htUJu5O5swyENM3z5X2E7/8fS6Ml+pUmFbq9IJDb6iCKaIeF4IR+QXQaTbMeKzSdfUVpyfCHZp9t
ELL924G3rZ6yq8cj/o4VzuMssKvqqH5fF0Dvi9R6Ev/xik3RI0FOi7tUad1Bee72AAgqP4IwaITW
KBuR1bWogUqr30NQc73rGvDceEDCTu6TU4Rb02+qdK2prbGOlBpkbc3iTh9RANkXXkvd3h5IuJUA
adybk9QRvf+tnFg1yu6wYrD7UbdTNa+JpR7zpDN5maRWzlnb2+9MJnFzaFeUAFBM4J1aaptOs4Gu
s3MVwINRJ/XRgzGSqyzyStQwRntMHvwHP8pBEZ1iAIE0POzUY+ji0uEGANJkU9k8dhso7+PGy72i
kP+0rrRsDOD+cKTG/DfadXMPPVKAkP3A4RRZZZBDk6DWOLoh6iTF+n4Nor2KdEIDzS7148z3gg9I
AA0bxoGE2bcUqYsYFKw0Yr2cE7TyeJS6vAKEkgGpQpSgU2m3y+YujV4xcPGDfJOFn0p3orik+7ec
GTggdm4eIO0n5r6uJRwCC5EsoEdAI4tzENgc6bomm3cebhp5dvZdUpp8DavCdMLxnnd2aH01VfyM
/V13JoZXpcq2KanPNSZ0drpVz4QviKMX7eV6vP13c+aaMb+5E9Hzf7jm2Z2bS4QVqdKrImoxmjzZ
rU7wKsrc2L4v4stv0TuYBaDB5yIAczvBzCwITYMtsD+9Pbv95cNX+24+AhQkKarYGkXPxNO7tpDh
PehiXQQ7kRe6yfa9MPLVpay7z2Ey46m9OzqiEfsWnb1fj4djjOq119E4QzJt4Z+DNMQ3VMLEtV2U
96tNfPLfu+uRAR60jh1IDRh9tQTbAV1EXJqVZzH5DaNf2yoPWFft8/BwiJJ+X1pSevUkiAq+olsY
e9b2VaWJPgplEvzQ6UHrIeSCYU5GEK5UzeAm7zef06bkxWRzWtoxbVubMGOSPBuskmPtDdbR0TS9
KZijnBtppiI4hsKaizkErC8gy+L6bVuY+DOEMcs5ynp/mPWkVW3D4ZhXGWpDFmst6NeUVdSYcxcu
/YuwnsTReb/4Np/siMWSIxGxF7qoEKZyLCIgypgKuRNmx5Ne3U5W4k91o8naKs0ac3ncggJ4GyBC
4itsw2OHhdXsqHfIs0QkA14DAlSP6CsoHsTpLu7xur7q+fBVNMRkSri4fB7rnfAcCQ4gNG8/Lc9+
jCqcGnhVG8w6DtNVn+VPtvy8tzHLhqS4sTn2VxnIxKffKEY0+hvUOXcn015SEsVkw4iK/OhyBDrk
SlbRu+h20hOAt5bV0ddrfByV/bYiL6i6Og9mkQc+PzUONrbNy8BBroKMuEZxbw4hHRJzyYHyxtvc
9afxbe5rZTuCaloF0Qqrc4UpCTJ9aJ1C7WbGF8DRoYST+hDD3UP07MfC0nJn49KZgwKDdipzZtii
2p+/ff6izvQu2au8EaVWucbVadwWJaozSNYv7Oqv25PXm2mLd6riNYobDkLhC5B+5O4JDIzJVWdY
i5KNwHuaSpKRKNDE5vewaKkBauryMEhvyr86Hl4LGn9TkJYICEAX0lwoZnkVTOE9FC/FqMAKzZV7
VPKfRLWrAI2zsW3CJo64zmR/tpz4/9Bb/HnP7fc14Xchk631Y1TLxar5JBaX/vXeRBQ8w3fWiGtB
r42zRhHRzUO41+ttCd6+bzAhf5E7B3+Z6ege35AM9XxPoHv5IUof4noy1dy4NHKpFjpqAqyOGjd1
bbEblI4tBq0NDHfqNvxapndI91GXA0Myln87K+3I6LeAOz2ZQlLp9ETtT62cFtvFJYANCgaUyYU3
VMF94dzPFuRWcuZ38Not89zjJr0pXlm+7VMNw5P7VhSkB4/lZwLmbgXdCtiTdsg2lfDDEEUK2tSr
ZNGBQE1oCDwAKCkHoveUMtZAJ84KrlcLFAfxBEKn03DuIaA1aF1z6uRUfhMFQjhHiYSuK/rxqtzY
XI9dr4MS61fpfeFf5gADpgjQr1j1/2yd9COzx0bUzJy8Y0gFDgLjqcjcOuSk1QgE29OsuFC+KLLL
CE9/A46rtzKkDpEXYc3XW0OVuo1XMK+u2D8kngJhKBJkySWc9JAuizl+v9mjhouo8rnuEWfv3dbg
tmcFjoa/FQPJd9dEHt6E3ie/rsGjNjYAJTdyFy+mMOXWffNFlHBghQCzrIVo7AMywtlcouUGdMqY
sv2JujKLyMlsvAbp/A5XtofreLd3g/cka9C31yzJ1bdM+i2KUzaM4TX9kGlsxfFTUe/Yz6WBPpC/
3qa+CvfksxctTHAmvjb9K/ywgj2XCTVmzxJn9VPAxq1rA2F/evCxoAprqUYSU/NqnoHMrSgKJyLF
y0Ar5Vabu/Ga1u+P18Cv2ew+1oYi9MoZpl0ydgpY4ePPnYuTAxVteHuBLPJgUibJW+7NGZ8a/fe0
6usGPuLfbgYWPLXRC8mrq3av4hcRjwVZPUlgAeDdkSoPRxcjye2b6a8kT8PN1Hqq+rJreEVGcen0
VCAiSQN3XPrq5O2fvSFz4oFvaTSEzVVDr7xJjqhnXGQES0I8mQBiLBbTrcfRVemisq8IAO+q5all
1n/rgEKgH6goPK+MlM3KS/K4oWAhqxE7tWx+9xDCKWgTwEcrnqgg/paZBD9lmBCe+/7j6HLxqxjd
6K7mjhRWZFZQ0fc98zQZvko1cI6qYhw6vn29RViRYaWjs1z+c+PfsCMaTuGKIxcjg/mnxB5uhy+K
PR2Dk4uy7gtFmhFmaAJRT2yvurCscZqKoi1Dc2aR0DsQ7xcHGDkWbIhOc1m8O25yi0JQyy9sGEbL
COjlk+RxAhvsctVNBd4DOcAwmH0Bstc7Kg+pt/xSj/2dkZWi/44o25TnHBC94CP+gDajHo9psSvL
KQR46d43nC0k2uU4PB1NAv3M2FglhBR4lop5kxhWQ4mc7JkRbODRZZHlIGsWaf37OaifC8/Nzadu
qxMnQUgKxC4kTnC9KlreipVT76a9kK+VVxR6SCRgosldnp/2SjXB4tTauug2Y6L77QvxHiiChDsY
uigY6iHH9Gk5ssehky5JkmTn9kGWsWW43YA78qbD/RnnQPReMw4jpGBTFhSkRPPyORH9JEuDVvyR
+priOj9wwFWpfOhWmDV11BbB0R+5wZdWUjWjZBxFKR6OYntXeUzHPRVfuYjg9OF9VHJsKAC4e3Sh
/7QIeAhF/eVKwDjLad6zxazt/O6k41nKzJzlEAAFA8KOuxFrWSJ4Q7WPGb+dfL7Eg2mB7LQ60tY9
5XRMZVvyi2Ow8t4z7DfDx51xjWed7OmJPVLvKMcfcyzdpRr6onBFQoxghuD7L2kD7GFy8ln4aG0k
QzvlxDU6le51Nie4PLbC/MdWpJcwTiUfazxBBvz6LrPZKGBB80JuIKaH/7pqHcMoVitk4hwG/BOB
xkpylmoGOe0VdBgd+Cgy+rQQ6JSXygE0UPBVHMbpCPvATpNmEWQ0Ko3wz4a8hQvL7hlcPGi5/AwL
j8QjrT0+oKdtkh8+Scar+fU5p1ZH0DnFifyuG5OFnSmZuhdjtKLslsjszY5wtujQIHh0XYd4jACZ
gY9zoCTc0FuhzmIt1I2AFq0LJye6Z13ZpgWC54ouY+I/11KrV1Vu8NW//USkzyJu3uyhL2uzVogQ
zhh3jDRC9prFldvCPKHUms8KNLm//DtGEOupIWClHqsqSPh2IROWk+YBXQQQXNGlHvWwdlUCQR+P
wKhuNyQUCeNT2oZB8nDvFYtFInMqptlL7ZbQi6k99L8iCirqv8KaWUMZQ7ghzRkPRFctrC5VrdtS
RkwGYoAcLjcBynvUlJjnB+L/QHXXiY0E2iCJMOC6ky0/WqdZJOeQpyQ7aElEtuaJLwWghN/gVpSB
cuPyZ8Sxp0a0L8q1sMOqmJmRUl+95rv4/UoVPT2tS6hIJvIhciwcBtE0C5Vys4k4DF9qGK8q0/vP
Otn30IPiOB6pn0TIT8yHUM9P2VnjbT/vgHMZzbuGn8UwJSgX3lWZkE0kYyWZbPE0xF458nUWx/hS
Zk3dtb/5j3Gbvl1FWBv34wch8RGWydF087VttN9QW6QdjqXyxZBXQyTtdmbOTYvJO5qdrG7t3/x6
jqS0HpTqppM27zcz22RqnzaJmEPztOKFAj+iRvJAlg0/dhAXYwEGohcxEY4FesbACgpjxnOp1fKb
GmbFWXpcEsehFivM4qZeickDfwytS2o3tHPW8q/fWkSMtG/zBDFhMl+KAvAtmbide3L/rTWNxWqa
OFOW75wUImukC68C7DZ7jst1dG1zcyhEjCd7jObWOTl0wrLoX7i2TcyDID429d1Zvlme+WFMcHCc
P+30ERFX98GhSNHKQ2634axSBNW9KzPgXy61lemx7LCGWVwW8CjNTQihKfDK0SMcQTzDPSbIxaTd
FUTcz5sEVTa8unvxdIjL1jNekFZXu2h2OmJADgNnpEHqlhEvKCtLVqWgKF9uTz2QDKrlqVeXIM9O
txbFmi3INsCen81rYoJ8Xp5qGXUPXUArQsgAxK5CLFnMtQsfQRll+UWYoFFQYMwmVz2POtSbqN7A
6a2GFhv2dcUp7tZ1ISA55n7PAh1ZMrfFNjKfu+PkH0A+Fw1fO7Nf9jwlE3fuXloSR+QF0ga89Rca
+O4zPBOOzqQe8D1SYQ7fSeQX27KiCqMuURlafUOnhE0QstjHpaLXIHmd48LAI9QZ/TnEef06Hu2Y
wDyTLwaZeRkFMrqbId5IpChNCOwGTh53AiP4NKoP5BqqJlRQqZXhNO1uTWyffjfqjxt2yf+tnFfM
xRULMwWqG8SbtgUqIW3a5q/3N6AK7o+gfx5PD8ovgjiov64qqSJRZolq2gOujmKsdFGzbXE95/Ll
Uce3jaOMhvVytDw+e16CYB9zTnxDD72PeGJg6vCgW9STp81r+LyUUOXviDKQpZ+WgsSYThCE3siQ
7mRbShvk6kVaGhp8HsY4638BO2DzXDmL+ApOsxSCo4TBAcXJyBywM3siw6yN81yLvKlisSyLwYcM
AeiTjQ79LXiAi4ZNW2WnrkWa+QAI1CmTfijpbZcxCHTfgeWQ0eyUCHd0iXG4orfZMZeUgSzDPp5J
1z1ZaR0D+e4hFaCxCzLU5x2hXr1+9FXZeANkTelLtshZyDJt0RSmwoo5RzUIEoCcjNimpWXZaC0/
bCrH0ewRW+H3izgxVH1nv87G/m8O49A/VDcnuKmDrce5EIFyg6fzlKCXVDsgyb+aaHdPfZ0MtlhK
LHEIifUySto07eZPm7oZACXhkvLlj07ZmOQf8rG5LpurBIMBlLCwhXumUURaK38ikAlQOQn3AxeJ
ODUoO1oMM1aVhw1BnPS+6KS9vDqvFaa9GSoPdOekDXD01zAdleCdsSwrM58jgN7oXqmRRy49foTc
wgodCcfScHDAGwcqIIB/EeK8wWTJEomjdk2SMAz6Vvbbjh+vh9tiLzekjLVLhNrX6w/wgDJvM9j7
HkOACbWok0nyDhJT/RRm/Gm6exRkitJHI5GtPr/g0DINTdBJvs3Yv14tarHX7aoJMNrODeqow4bo
rddLz7/ngZpf6+YyreFhtOY7+MMmz7PT+mehrsTkRgh5VN3UNOTJJkBH2NrBRq/6uG/y7Mgs+Cpu
18Om03mcfnW8n/qQdu63pVHtj8BwcasaxB6+6z5RANWElAellj+GsVCIDxXIPoeNSWp1oYHpZFp4
+QyERNS0YFiVeyalDFowSU4kcmbiDvIQ6fSHSI/1KRgScRIRzdtrotpw0CVWwGP8K+ehbA2rfQ5k
IciXBw99Z5hXnaEdOJMiZ0eZu0TIJbpLPocf5YLfbUmKme8aHPhDBhgQ2JkBWAMKCnm/w3o2fwnp
0OFQAyqDDBYA6gMWTDLUGoEES//sr0a9vppzh+ZtxKvP1DDFb7WVRHjp1d40BmDXIABxSatxeh47
f+V8se7cWaEVVr9BwcJQtMzWuVlWt28oWxeaMRufnCbFWhWYiPoWdccrCSwFY7VOK1OUqKuzYN3o
pkiN8X5jYOjBCbLnV/9kigXHxBGKB3h8SdNN0x8dBX8dzJha/QUx4QBax0StISf6WcS2HKiVk+EP
DZTHjh32sp8nOlWx1eqcRO9WYyvrBHXLsXYnqZG1LdMvfzohPJGJB9fARPKwphfXffobwu1LR/lo
Hdp7RvUpzPD7hrRaWcvhSdFCcw0aS/P8s+V5Nbk3V0IILy3WSkpZD4IcLnGfm+Lzavc49jCqmjLM
sgb1cb13BRE84rkPzwUQP66bADhvSzNg5wyHSSaMVjjedx08lVcV/BZYGw6na/MABm9BwKsjkGy5
7rE0yNbNpXYXF/sgXjM95kPBjvaRydL5xuk2p5ZobCSL81yc5FPvI5y6jIY9AbkymaLO4rG/XM30
1vqkzpHuzbPeJdLNU33yG8PAAA7f+e06VrfJLCsPDdD5ttwC1nyBkKGxuqR6IjMxCXq9s31qZgzK
YuDXcIy9J346dy2/DGo7ZBhrBD2HVmq429031fnMJwkghAZfMr9Yv65rWViuOIH03fZ0AYPKagk2
CrLtES4TW2V3Zt1zR0AKntFKvP0xMhzjYE5yoP5HUjqv8fq2b39JtTgwEMVQusCqhG1N3J4Yq1Mb
YNREm+BuDXVMJdMhhxJ7eg8upC6uJBI2fM/tfocOvsM/O0Xg0WkdIG02isekPu2CHO3MaqIxWlML
Aft5shnkCBmAF8fd8RwkBkvyMNHhRPutEIq47xO+tiHI6WFtuw9tTpDSlUplWey7ZzHuw8bBVbit
WIyNwXpbAxmLVxUHHcPLwUrIvL5C1ZOTDyh4+Skr1mXjBz9+A4lG/pxgkwbwTyGxrgjBebboCCZf
4ax2y+RfVAzBncqlH7uCRvUHh3XDTDeNZGaD6YnrBiX9DqGsZyhSenn/+S8GzwIFk0Ujipb9xj7K
bkGAz6K26t12QseD0BK5pao+vWlbQtKW+HHGdDLTi3/N8ADYap1fCa/1D8ubch8KaA10dJqsZ7AP
LtUIaS2vgFnH/E5y05gEbnoEMuXdZuRohaSLy03buZq7VGoiGIwY1VBfTHe0hUT5Hjh8ZTGCU8sG
BlemxKoDIOHYBZTGi7JprqOsrVHGsyAh2PEKX9e+6wFHeKRDsKjlcU28Yfel+K1FctnjwxohxKS4
y0CiuQHq8abDUrw+1y8XIBX6ERoDEpZFxr1zv3+aO7RIOo9IL6NIQW4m8qL4eTmBkbxQrVnIEchb
vr9GToS2y0akKGBAVV1BBhUgBjFBGUh09XoU69RUkp+1dn6QZYULguicHEI43umWQiVNK84y9grG
M7GuZBeXSVrkYWe0Vvthmjf7t8fyg6SEHfibUCl2BpAODJ9lZRbEl3V7TQdXYWkr3YDX2bswBIke
3SOXPDIj4RiPsHoVa+pgmVXOs07cu0qmyhVQJcN2XSgCZ6D/7370gUt7234X/7K5T536pu6A86oa
F7qA0Z965HzkGbSD9srxj5WbfqGkjFZya3KYzOcua42mQ3MGDuYKen4oQsQSGjIC0Wo2M8/2Q+qq
M9Nk3lxCB6LSt7/N5atG8P3al/T4Kk3S75b/gjn/7CfdCYeXGXBCG6aGzIbShIZMgCvEwcm/zDkU
e+ZgRhWAjC+zmmNSBT8k2XAlv8/syUNAlM1WTls4tCIBfiuEJSU17I0tK7nxdOZOhVkWas1X+hlT
WVKYdahQrKAsxY35xifQFeOZusv+u5zrbMCWiedNfUkmmpeivmSmmiZsdAt9f11/JbNNBEGQaz20
GbejaFO1CBP3/cH1A9kDZxZGgAIzR+A1mFUjJIveQchkHfIVqLCKMoiTHqKIGjWEeYU6nvT8MazP
WJ38CI1s2g8SlMsPWyB5ivzvcs1VqL3dNZUTChhSEzGzVbIUnoPlAYFRAAhb79rvBgA8M787HTEd
aeLIhD5aOEZrcsdzdjhXWJnWN3mBNFSS10du9opmNJTN6RMizomDywyCRX/ywz7hzKMaxCaciapZ
ZDdZI/YmUiYPhvD/qU0unxhEG6lWdfg5KKURof2kRPVFL9TxWuApmJhf8Vco86gGzqwUZTeeCIlS
OX+iWPhghXwz9T6bdJEgDAajxQqA3EqAOPfQ7VRIUC0kMxMH5wiUj2FqRvqydnLCqM7zDPtMmmHx
ev0wR6qVo4Pf6Yrjca7IAAEngqd1hUhqsPcQkRHTPss2B9Io8XPn5EhToDxEZM/OEZqwlImw58pS
ZjXT6p5b60GDkQEs1gjusFnk/FvPCuC3tGbffZSWPuNPggxaeOtfen+0VJtWWSf6xmBw9JWQ6E7D
B01kiUC5fIWEUidHAEekC8YAyZwBeHHw0T09sDSZsyxm7b9NBs+4fi/NS6T7360ScUN/vifGpQno
1Ko29eIyk7oS0rKSfiGyFWTtCYrN9sI3N0DZI0jdVvIASWwikg7NI2o/Sy189s1XKjZwQChmpoKH
revi38XRiwwoguUK7IGJM72q0dvFfyKH3PQ6I5AxlH7smI0lYYcLxqm4Zc1+rAO3FlmVJfagDIgI
mKm2vB6on/eK+wUzwJYO09QSI19w1RaDWi4b2nZwIUokzZQBbh46TFJOnrQ8W+k1L0r8duejeOIL
gDabF5e9eisLJ8g9RSsLhzZBsYW66qKy9vgScgbIdpzoGW2faq8sxQdg9lWn58wrcMjNinuNjFSD
b8Qk/N8om+90H7HlcT7k7xTp9X7VpTUr7OvTj2BjxZLzgNDCY4HEaRuV+3f28q1FByhSe28SxZW6
oTe2UICEUVQ4OTsRQw+O57wObPdc/OshPbHELokOPB2AHB388T+Lk5tUiP+8OZhSg1kypG3uMCB1
pJfQuhY7lwYbZT6Bly3YLiyWyXnhdy5cypLnhXvyyLgl/emERXbmdhtp2PKTjI4/4GqB+L3YHxI9
h2Gzewjqsp2L1epp2AJ2s7oxA5nDb9sm5Yo7zEv4LBaY8FdergA1Bfd4DF8sfPZWWjgdt5vWenKc
tCDUoF2Oxng0XKPZVZuvyNyGS+PelpeXiIo4hmlUht7LmF1P/YC0stNBGsiumYKaju7ua6oBSNsz
HV/PMOSs+tlP8hcj4G5/QzF3n2BA83mRkSClDSLucVAdNWMDCQZM9H4TrGRFvbX+NkAu3/2/aC3n
t4ACVNcwgmvlwbdy5aeKmTnf2qT0oVWZoGxVZXFS1hOu3VQCdORz+3UqfVds+Y2y4Qf5s+EApJoX
dAj9mjsUs5bnZVIhw4HMNsxcudPg+nZAGeNfvDvFnb/jmR2Irta5g+nIcMbz09j6bn4Mb+H0TYQh
ZZdvQ2icAy7x1ji7M6StBYwe4zS7sZnxJbO7grVZzePiiHDXf0qOLSFcgEX4NoQ7F9CzQkyptl/K
5c176TXuNk9VtHUsG2m/7Js/GKtk9C3U8IkMJcGB64x5Rcap13AwNd26JATvD0fvojsWuqEVlddX
aS69dUKxq/7ypACjBIaOnHgHhfAN/yWdvGC/5g3CpspKy/bPlhWsdfqcW+dwIDxcODIPIjsvonBs
ea7OMgoAI+2EkYtzjntu6ROaTuHb5xI01cea2S/HMvp8Vq9XDuR3T7Y4ElUSyP5gl7UJkW610RCa
KPbTpbl61P6n8gD6BLmlHiTaj1USbyG+BRaRyyPeA3S8i/ZsTb+OUg4+u5U4J97ljDKgfKXwUl7O
Wq5YVhlUVfh+FbYaK1aA9GeyDGeGWfi1yMfdmFl0hAaY/DYzC04Vcx6mLRZEYC74qjR8agf5tjvO
0Nw2WpxyJ5xsn27PYReN2WZZjoLDApa1GudyHX/eDzA3so4Mm6sUL89JR94VfJT8/Bfg8pW3+Lbt
T6iFd2yvG0n6OX6f9JLDFrU/kcvW16/xGskOJLEkl/qu2g2NZKfj9qTJEKo3TgvcIuL6JsRq57B+
9W/BoXa1vpQ9ISgLKbfauCSKNV2M7wF8z4oyZyKBpZdraCsu7N0UCR0l04vY5JEt39TUx+1E5iPO
FzBhu//tel0ujWgiHZdbC6SJ0MI7jdyLALz22Q56r85c4vo/9I75yU/Ipg6Sf8s/KeU8dn+SqAfw
6WwM+b1Oka14MUEcGKp51RXulevC774NvJ6cuYbJhJcNWLiBph7GGiTlj906eduIhZdIrJeHIoGj
yQgpbmrmXsbGTHwv+qNLTMgy5rLIL6F65SfiNIvgufOMGQfgknemr4fbPMAPS7eV8JtvsygnhjW7
ybzTRTSRUho2ClxBeSCFasndIfXQgt6IvoaA8w5srW+nVAAp19rmPI61XyJCgUVhgefROVvt7vJ6
gtaMbf2bFBRtjKz9OnM68TieNfegDILOZ+XAu19lVzUupD/o475yh7nYx5KB4FTiL+Klu9DBoy8J
RH8tYPd3y1UNeQ7Ux+CD/GN80Yrbe797LgkHu2HtIYjq3t53IbUQ0q0QkMyFFF5NyWt/2fFnz/il
67by+id9fqgUbp13kVN/ZdiHT1+Pre9+LWuCPmzS9xY1x3DnRv4yF3sbWvlP/3inLvwu9rCyg4CN
mdyG2V5511GN440t+n5mtBx4nSUvJOPIM95i7oA48J7FIr1/WHHsNerbmnxhP01nEDxg/mLmoTCL
uweERYSyoTWOaXL302c5V9L3fJm7w0N5On9ykKIzYjPQepEguLpKsyHrsrbPr0AmW/22DOZ9NWGR
MBq1IM1Tzp/kPBIRcyMxmPNyrk81k5Z9JKp45RA08d8ySgLgpN8Y0qymQa4uFgjMqOKjlW7vpxnG
wGRHzhQ8PlZrXj8Nw04dw+hCZlUcdieLUGBThjLUnhIbbZWX5SNYGwqZTZPcXYbsGda/KEDHy3uR
N4zyufiqLkLO9LbYYSTYxlQsx21KJQW4v1dyXlaYy3T8fpSLyoJ55ddTfOFfC7BeTOX8EvDIr2S2
WX7PcNmwzIaFg766C9j/0WDHuGz/tWaZoNJ0pq9jOQOZRi4SHx/SbeGsHnf2RSPIu4dsA/7ro2W5
t52J5qtYsirrL4VcEOLjMLU1/CX2eAMo0YbMs1m9yfCvfbm2CU/fOFG9o9iQthmvUSMm4jXjJdBa
KnDOKrI07hQyptvhyn00Q6xBhCODNr6whyZuaLlaI9JzEnVbjK5tVdI/DcwxCFGue203skQWdPrF
RsaC/aApF9FPfXdeGvqeBMF9WucVxRfvy0jTNeFQ+AJ1Asge0nMQwekOqK+6EFeYG7HGXcpqz3aN
g9ZYNd1fcJM5+0dD/ILxV7ey1SdR5bxblZ3K9mTdep6kKNtx/I2tyC8lyKxZlLmTNBM4w2p/d5hX
g9CmZAteHMiJs+voc+4kNezjwepEyAX4YoTOG4t+uIz0rBHUyi8mcSnr8bSgc4ks8f+HP4YN1odR
+RwpM4fSPPzE6QFGvdPcbbM1C9WX9+lr0AE69JEjjTUaOc2dlia8fyv7hEhScTycSOY1yBvXFJjZ
wKc+Q1G30vGs7/g0Q4EOD2RjpZ9CQbbkcX7yJ9Y/vWQ00g+U+MxTVTG/0JYAnKN376aTGxY5hHkT
XOjcnG8qPkA/E2e46P8uLPl2Swb3xy5XuXEwXXJzajU/gnYefwj5COIWaMZteHX5fH/KPOSM1k9B
aJ4aaYXFufT1p4oSpBKXH8DV/BibOYMy8jrzAdLYHo/qfDqbQoGMeQ/DamFDLK18T/tZu8k8e1gq
7GSSUd9rlgBoohP6UzfMOd3pHvpBj+a2gDEn2aNsJHLsx1AqdHXMZqwsLTbwSaOGFQ9OItquvYd5
Fw7EbcT22JahPnpmWcbz2SbBP1CYQde6I5ltEQ57spF9z4JXkc7mMlkA1DFwizMyPoWKrwhifKbF
sbfILN1gWYtJzbO24dX4+OkeuijMPEDa+koGkLHlRct3lhtInr1lic/kwxF8CfH1WegXyFItNswO
MoA0AO4mhWt+UqF4JB7PVDptA5VHZOsx2K1N6ikuF98Uy1Rmb7oFWHIXaVPJ8mRp6FSjhqWPLS5l
No2qqIuDW6TgujmpaklOm9/pzEdS+fEHm3dYYBxF//fNjRtpswq7lr3iaYnXY16F0ppzzeh80Nwy
6mGN/woOg/eA38/9Ra9rXPiKBcW1Or7btDGC54ENvTtfHvR4yeAvoc8k3UNk5PLvjkSi3c9qVzcO
SxA3BRHoHWyTASZvNJn7WrWipAo98ySJJF8DaP8mQI+qYm9USQt98fHxZRvL4/bzEI5tlLo1M2Ga
1qxkwD8iLfdkQD7GezSMFzUGfFlmW3/JauAlrvZRSTmXe//O3LpGTC6k+Nusd7jgGVTAT6ZsMyKC
y+t6Brto9anixeRTYbEGbtOaWtlazk78lIsVUllRERHfOAxdcKJ/DoHs4BTCiW9Bf6uOLbjhkIHM
gGq9psfDlRkq7Fk8i36opnWwkOUEwY5svNZ3xthl2O02mywMA4ahYmmvXFBbMNpRiVTQvB+Sk9eJ
AqlReOhSdWnvKMcdq1JwT+kYD9EP1mmbhX7MBmWcjIj78hzLUV0+tXyqvq9vBtpt2V03mbm4Zs3s
zd7Ryz8yMK4w3ToZ9w/7lRdjct2IjH7ebQyZswF0Dau62Sw2kaJEatfvXiQgUxATti7Row6eV0ar
pRJ3+YSMs/Ekxl47C2rw7gXlGU6gBdZU4BJNdanm/ONNmyQS3SgaFwI0aQykrq6APo+oPmY+/oTY
DN0szk8hkd3QmC2KEvmpSc0hv+jLV4sCa0m0ZsxcEfvhtWUTdygLCKhg3dIdjExq89nUjHwRBZ/9
Ivqhk59zhHLUZ+hNqbkn+aeYbI0lza9JUXclw7+Rh/q0WEkTPltpuchynxto6JKm0UE7F8JLKpvc
DD4loERzuypqxWTksFz4dd2ilmv9JtdtG1/TGuQJIXDeg3n4Ru6Lg4Ah6aat8ZdSDDNuTUN2Fzlk
6wDXXVxwxr/SrKGztcLBXvwbbQsE8EkVVN/AlzixgEllAn9pm3Ecn98XwMvbdVdrMl81O8XXGjeK
C5kuEl1e0NnTfL6WbqhdcFZLjldOGT1JQ53w1BYKEzkDdWnQ/U+Wby/xr4XS0AZzulMNS1R2RmW/
GvyM7j39wD6GL+RGSsNm2/rqE3tEBuy4LjB8Wm3KYpYr7wJZwYQ0/Og4sxXTIECaogQUn53GWVxd
vHlvYIWLmHe7RFVmK3h1UE8xyh7MvIfd9VJ8MUyFo2z6ztifXZv47vMuelXBMKzef3tKq14joEpN
DjIJdk3zpPWn9H+OZeqmPn75ZSAlL5O+AuQrFG3dymXW4+/6nlze9yLIhoKus3+tb9eOE3CGsg0d
kBosCixGraGFW04fo2GwuL/Z4XmrD25wK3nS9j+F10zDtbTQ3NbAaeeVnU0DbJwCRBuHHjDclXz2
oFf938SpRgUPcUY78UMJQ6+jb8jAH+lxdAn+/ZH3lE0qxxr1HAXet0gH9XPhQRWTQfP+gO5Ni/ht
TIpjl2j+M6laOaVvMHygLqxwFBUxEV9SARlGdcIvRo1B5mSyXntXYy+avhKff5N+SkqSvG4CmEeF
nn3IO8WU0OIyR8SnBIMErZXB3oRybZ3qI++Yodn18It80pCE2exFjOgOqfLQHPaJir+cyTaCLaXT
y2XMFgcHiOCDbPJajSx8l+KvAL3Fh9jB4cqSf2zOnM23VKZnW9tvlx5f0CjkgJJkuKT0zGtzUfC2
81CAtlBCrMvmTCKN0lxwiYxjcHezODVJclUajioEuskZ5r4K1txX/ZSASitnohnn5JV0OvbZPg9i
AyEy1EzHpN3mF5UMJ8hE+Sk7i620FBkVWgiQ6BD964eTJW3HEymwqSoG6Qd/gbBTZixjxH3ARb6o
dX8YF2Kri+U7Kg0NUv7md9iKsYgZx9i0b26Nx0xWBv5AJQry1PL1ibWOssLJXiZ5vWNjjIrrZxz9
gLie/08/SjQ/fWqog1/vMR953itJ5T5nQEdth0ohvO4M4bQRNc8rXzNbPl9lyp4w7+AMMhz6h7VO
SNcyLrsNXxsOQxGBh//pTbGnwyfQP9SFIZAm9citw3HAgh3b97gZsH6/Y+qKU6q6y8t2AbpYqhGt
2AiNLNwnUtD3tVIWNuHKLxjTwenGjGZtJNlgAhaRVN5QlXTUIgOYlN2IDRzlXKjJMaYECnafiAva
lF78u3EwdNJSTf686xnlc0VUDXPHq1wFZwdSpaiHvZRrjwbvHwcc0IrD1iAVLzf2TiPz6Bz2N8ty
0vJWyg3jlObxQ9/ptPbaoWs5NfBiaeXcQbg7xEd0ZEa+rf8EtibHifmFIcub/bCdLGkLOJVFORud
UUoR84lftcsEQ4pc3wSvWsysI1xO4zPV31ECdD0wfAopblanwC/VRKgsETHgSR6llACg8T7fpyTn
0zLic7qU4VQId5YWAqHYqRKBGG9+UFWJMq3ig3Xdz34+PmWeQwJHMy7QgpLD9TJZE3/Jtp7N/6gG
hKHNeerP7sh0qevjM2o6ytZYDnD4YrVXWe6bxwUnse1Eto5D1BrjK4BpwuBpuiGHBtvbvkPe+1Mj
Rv1O8PrcXD/lLOi2LUFZQ/kIEh2x7yneNACWRue5Z9rCKotwodUQaUpFeHFqvlUlJDxumyf9Dgsl
tOP8C82fLrjaMh7b9EL09trgYydtWbiSU4PskGvO8hQ07H1fVpL7xLmjQldug10zVyZe3FJ8LRMX
bDGUkjUsu0WP3hdgxRKQqOFS4Nqi9eReCMes5GZSb79oRDXs6mvGrU8AZ6E0/70m7Nts7LPeRjTv
q5fWiG4rhZcFbiLamqz/OkrFAp7fS64rpU/mIefcFBXtaYS64i7bWbvKaumlMQI9rFmdhfPjWIhQ
9z/mhI9XqFgR6zK+El2abHy3COxCK8QgKr89CmR0nkt8e+tL1kVOrVkslr6Fzodi/b8pkUqOFqEx
QuOui2cigwWQIEB3DXhCdqDSKB/0Ole3d8rRoU0Ak40IES4w/ULbXbG4Ap57eaw4hi6jG4J+RFAJ
EZ8cKgQmAUqZea3MGSF2k+aAiFYScVXrH6245e25NacGXHS1LZY/2y4MXEzRdfwhfhFCrXpJv8t/
WtuC0dBemi6RjC1/55G7uJ9mMZarII+hT4SbLKZukNR/Jigl3GtsamVDeN7DyUsMDfxLCZ6UD/xy
7VRYNPtDPi3WRXu3D7mC7L3VoTjaEXzf8gdWdw+5ltlwk2WjxHTYmtwKFs65TRBpq9pOVisrQwGJ
jczINg3FkpvY4A6yI7LFCo5IxKX/Inz+6i/kpTfxCOOP6xgVfnvuS77dJ6weBz5Q9OqgPVQ6dSkV
Abt5OZJDVqBAXmi/8Rcf13aMXzUXglECzcR4kW+QTq0ZMc2NQsHzpUiQLn98eLvBiWJNgZ+/EfxA
rRLwhqC7593VwcKZDjSEbwm3vMJHkbqjLrRs5QhVU2y/EtUP4yZUXhkdEHTVM24AgmPD7Hg3Wo5G
8PijFzKR+vbXGqbmEtbfmTd2vzEWrK7T3dS1rRXPTUmoySERmpkFsBd/+Ik0iN3cwnTjGNGBOIG9
xnz5bgkJX5kXFMjpXzKLW6FLpbnlQO7QVtKYydqIHoL1auEjuQEI7ADiDvfQZTTrDE01IQ3YeWqh
fUag+kwVEBi4dawSCtL/TF8lpxog4inEunZ3PK3IlSo6VYkK3WD2nqzorb5tiHqHJ6M9P1b9hFy2
5accO3RIceug7nHp74uQMmkA+QT8ErLnjIAsAkdNCzSDxjb0ksCTtSsCuROx06hue6/lBgXoh/Dz
TaRZLScUoKq2gaEkZmEXEzqKyskepUhKpLxpk+7v5/QKDIFRjdDmQ5NAsPDB82GJi+BXfwOvs6GV
sofKQ4mkgtJDXcGP3nqAyFlAdgiqLrTfshYXRC6jqxH4WmdYWP+SgB5KDqH6IKmgmwnGWMQRmbk2
MZk16bynnhiw9Sabv/h3xJBB2KcNf1pjS+kppgg5R7ODHGAlVL3/uiy1B6EQtNBnrWIH8ubvHnRv
8cflerCYiattFAmWFJ6i4himD4jV600dBnR47r/Nw0T4wl2Hw+xH/bEohKBYklZHi9Xjn0nefXIy
NPxXITYu5lm+0kkyzpztp1AdXdKPB6Ue8T+JsKwhlg/7ZqIJ44h0YN/E4WICwJN94gtbLa1vhpz6
oQa/1RS4aOOE/08xfgi8lAieUlqsgBDafnCK1j+eDl6NbOmrmp6U0g4BuDmu1pu075VNOH5VSkBu
fHO54woyR/WUqvSxNkr3I2R1EYH5fW3TYMoNWsy92H8da6MRK/yIEk5AF/KUOEvWttCmiG0c+TqY
kxCfuUtoKErTg0tIm9+y1lytRqYGEWJrbqWnHyYCul1RIIv64q23Ae0ES9Dxj+EwP0miKWZN29AZ
7HBNaSlcaWS71eHxn1DNZLKENFSOCssz0LdIkRGjZnTvbq2t5kNZf9uRtHVSGN8ky2MXAWpjpjqf
W6j81+LBYPJTm3R0T/Xr9xeDuaJGUbC/tPNGdS+hMGHN7cGWeWQG23Up2/pdn4hxaqT6yQeckas9
RsWPE8qehN3xb9cmkZdqQgtmEd7Hm3i6pbtvchhJizEor591hub1Hf7+FAu79Xri7ucdPfvU4gCX
QvInjQYEdgrropjQF12pKADK0Yp7ca6z1tAFJCBGoNeknmx7iJrxrl2cDzjVotWCXAfU0dKlOBk9
5HL4xqtJ0iScWUBhD7/i+W0BEm9ZvoA82s7gsFVXriPsQ9+rSTEYPfLEpCuK71Q48fHdMQVNV3eP
60is7DJtnLAgWbWTLvjCEMgwuI9G4VYv2NytTmS8G+8j5//OHPjOfRaSWl2tyT10N8qNs2bd9/nG
EPBZabbpqIYjggGdDIYVYQVkXj/UFub6IwtNAej/FEwgKswpJ7L0gH5mvAK1kf3e5oiJ8XkpAONH
keOBnN7K35wnzN/FaaKfhyM9+b7uMPy+cPE6Up+2YOxn549zJg7Jn+gBNJIuMYHRrIrz4bK5+Ii5
SFypss4CHaMo48F0ZTc4Ht0RUWcOP11O2vT5jLwfiViTXW2Xjnbzxk4RPG/+d1Ps2bRxDGJPiqMa
ZDTthf4alIAfSRtSQ4JPAtMVNAfvF2F14EBnY2WvtrD9NSa0LOHsxqYBdVpNzkQnylQzxmfhIfjo
5XhbTpq7i6bgFdybNTrX9GTJoRihR19SqmPz4IMducss+8Sd6jU3pdNNIGQ+fS010o7YobMM5wEH
jFo6whbqf1yUXTgypWldy356SL1xYyWcxvVNGyUEINBMH7F8fMLNlCJDVqhxbm/7xuvbVCDHvaj9
iNxdNg+RjOv2wpSjWNd4PyVnkCQrVa8zKcwCs+b3rAE2B04sLBSqvUSBqc3hDWwtO8bGR+xa/aVi
E4e9Pd1dek8czFS91SITCBYQZSfpUtGE9SE2O+O1IYcE3V/fF4eYwG6GChfzNPvYIDutWIbPaXzH
8O9jO6t32QehiTYUmLhO8I4hgQco9lJxXiEb+Q+JglsQoNxSSDqqk2L+pqV1c1VLlWyO5e700Ev0
QaQjlRGOU443WTVQDCmNZgxzc6F3zzo2QLPb1XK6wmeitRhjS/i5sMdUWcRklF4NIPl8OzGmxJgm
qoKNy1mqSJGkZyNirVzV7oG8trZP9f1Qp+brJLuAsKG+3IT6S89aRvXezX71OHb8bRGy9wde3Tnq
pA6O4qpbgY6TiAynbB1hwGu97qwFv/SZ6o5Fg5esQWZruXHr3z1LoScRQmkhJk/UQmSruL3mwrsX
PfYi7aPQYcaHe+PG1QYWmQXT1mm8HsQYWpj68jY9Gmdnu318X6r23wNRni6J63/xkBaOx9qgpwLe
e4p9dzXBC3pcD5rgjLEsCbdFKKwn5ZJQrlftgKns++arfGijKC5OyCOzty3CAC6HZcSCDQZypoay
3lzrAerxsE/WNXfTvbHY9jXL9lVoSnbgx/3Qgyv8yIpXKOCnEG6cPDZQNCoKwZN3uriefYhFQc04
43Gh6dLhGYfs7LHhG6fwIjhdlzhGXOPN5UmQa+R2mavPf+3yV0LpbLudQofX37Mlt6sWcCjxIuLW
5wdMI4YZDI09VBVjTfmR7XYi1Lqz2aAk+8+qSeFZ7pxgj/vUADDtEUoWHRk5rdK7hmQnh2KzqTQs
iPaZ6VrBS1/Iqy2fMJ489JfrUhWl10qf8MpqqAVjI2J8fx7fR8bc4jdY+rtLH/nP3s9w45SCYqWJ
3YJjp26hdud12Xf1hqtGalZZqCuUVqtUe29ThApXwQ/g1645ZsgNFusFudgmRVpRKE1xzk01QR7o
FF0vYumEuP/Ntqp14KAeUX7Ow3uRS3TTkvL4h4Ye4GZBJ12Vgny09NBlbTbAFZ4Iq6FdsazC5FdO
K9zmbxPkZ2S2T7wrFnQHe0DbhWre4ZbKHwmlF2RUDSBrTOBvTEqVA/G8mXAnrVV37hv6cn4HC3Fv
ZlU5bx6sYQjzbNqRY+NDebhFx1vb9shXG2Spa3YcFwaJT0kPPqwsl9Gc+8fkAhuhzOssNqaLIoQM
K/St60t39lWLkFh71H97ltp9Ht70lw1B4mpQyLhVaxBvkRJcxnD9OXSKNBTE6/A8V3bZqa14zLC9
wGwqlUK/umNKzYwVEyFNMdgTZdx+pU+Cj26v4Zalc0KGsZvOjiws7yA4NawKpovCOcyV3xKmDtzL
CO4m0qXu+takxWx+WaHq9mSLFlsBu3YewX0OImOalLveDeoniWHEw0Fz++R8N/kxmooL/pgCdOg/
sUCi6st/Rys9J9hjSIweI9oOlKpAOBd6eub8/08G3JBNPfGVzyF4oNzznUv92RTL3E3Xn62zdWfn
m8htFl93+qfdNGpXEJ2WQ6t6ecp6uoOgDlikaP08yQc6ke6nW6ENuCqUsztiUB5FGGPC3YLxVVwQ
Gf5GF2/Ic8jHvxeHOQDw+Ak/AemD0bsu7kCVunHga95akyMyLZJNEO5vm3P/cavGkDuu59AHprfA
mJMf8G90vidJjQWoNgC05GqTIRUaWmQpgEL8gv+QN9VcnRzD0cBgAKYDmtsr52OBdlJ8vZ5bQG6v
UHQVHETOni3/EBqs5nntOz1Z60GyPRmwseLWqHa0fFcYEXeWAYbseH9r+5oTBEPTB5czuKYupTSZ
Eo7sn2vitO4bY5I9x06t+BDyFTh+Kx4Is4ry2f/R50CJT65UYqdJKadO2AsE0xw1yL7MZvcd27+K
sllqxF363WdgKKIWcawb/K2s5pftTXbKCpQP0K4gAvO5MobOpl4qtrGp/G9unt6t26quzSB0CQV1
MPLZ9Up7qnQ6M+qrYXj3AvZF3xHzogP/pYB/OvPGP/kAneJo2DEtOoAH40XGibycNpXhzR3vAdD8
TSEV2YYAfWW5svfqIelxAUyG4Kp/cPDJsWMSnBRamkuXf3bs+28JuTKrRDBbbayglWyPrkmG7hHc
l88wzMgJKUO3RUSIWrKNBVL6pogZGQt0Ew2Oxu1yE2UX5GNtvIuEL0fxHhHmrgw+xy3qWgxY/qDk
PqP7DRNkzbFphNMLK3XjYaeAVQTn+9LHs1gryakzZoElO7dUPqX19dLc4DOYeyEl5HRYEvi8l6xk
0km4WKW82vJ4YqzhRTIz+KPXXrMMA6M33VChAwipIY8llDyKcbjU6AVdaeDFbac3ShswGinir/z0
SByILSv7gRtydjn0edZkTQ3Zno78k7UPRdYMgn5I/cnqhlPNT+mTiU1mnEHTxMsLENg/SRGcOeOQ
dtdxmuYmmx6nGcr0+pNITiguWoumI5LgKwI7kSQbVtJJZMj1IoiMavSCwuClEKfXloXlqRg7wM6w
MCnvSgkkOescoGUhZeVFeERRrMgiN7ozZQSO6F+VPzQRDCLafl3VeCSqsodFjiLj+FHB9I+doEvr
WCLX8QE7+jc697JPvrkaonaCj9Zjit29oegANU1c+E4TzJnoGBOH8ytzCKPQ3ENkjQJ0eVSoLcoL
K56z/zG/qO+yuq2vy89jQJMqAIFXt4HBkhA1K8RVA5wQnOOp3zJER88ebKBsnoyJVLhLErSpmcLl
IYtJZggW4boHNoF8t9RffyaZ/kvvrCFY/fNpkWvQAfmuJ1KTVLBQ/TKLzXfxpa7tInxddXw099PU
FUPIAiw7BlNopbNxQBA42mLgRg+b02MKxSJzwosbULTLRZzzSF31wQph+DExg4I/9C/b6HjzvtlT
B97ZBI2XRNIELfRqEVvtu7GkvD3PAk7CrYxGUyo3DK6aOH2GV9R512INiaaXzEVRj1NB8aPwkZSx
MUszBg2SqHfrvb3JaXwUcdj8qluiC6f5GwnRrJFJ+k7plpuROHUbk5ZCA2yK3xv6bCk5tplytkCd
T4txj8gcwTNI5/k9mm3IXf+BZQeaP7VD0Fkk+uWlporfIEiGvx6gLihLjAZSBhaX2dA3InqN1f/+
XI7WKZrY1WTaV2A5kT9c8rJXgDJ68zd4He1q9JwG7c2mFYRS9/M5/b6RUG+7jkuYHQKCK+vq1L5N
/rO8On3Ok3HZnU35k7m35ON78acaEK6QS52aeKiyfULTwZhsf6dMSjzD+UFeTMTYvu/1crYRyJLU
RNDjaEEREQbizAtmsFaeOa2HNvVl5C6fgd69uq4mankQdj8Tw7feE2Baoo/jEA+mqdt7GxTnwPPr
FpyA7hx+Np7xlNEPzG955hhx0CiIkn8Pe6/If0Ec57cqHbSndtJC/vr86WdS0ARBY2xnuie0sdMi
Us53IAjz+PPJKRYZ6viQ3Qs1CaU3mFzE9Odrb4AKvHgQPz5piedTlzhVcGnBFJ68mI+7ibeoI7iU
PDmyv94zdqXDVgxlRV2UQX7u88CrDxxLCnUHSqytEkvp96+a2FJ9duSIM/v8p0JWr/CcVfemE/Fc
/XMM3gk9m7l5d0OpqpCi4NtUHgCQ3ubrhBh87oO/FSeM4oLadQ3+8hzAGEMlRT9XQSQ+hO0MpDYN
Ri0h1l+z6tn2EfiNaFoKQyJNj36jqQjJOVzqXbdl+mnYdGdKsibp/yzSk7FoSeZZb2vhKXEv5ZYD
DS98GvFgJ/RuPhiY291wPyYmYIPBrzMYxTppJrkpin9K1MdGozFv7CROtTmos+ZfP5avl17Tkrav
W1Qbu6nJPcwhv1OpS1RXrLdCy5zEVn4UdD/bcmgVIo4XemFS7+uOyrjoWbDeFHBHTAEtUT9bpF5A
qd664eOW69QtmK5+eSnbywYcmzv/zn+yH24jOS165N/O4s4KPnYNHo86jneyPiypHxeyTYDlAZbR
3gDAT9XlzKH+yQT1b1F6NRaPoeEGf6UakXVfwZeRhTuXEnkTwKfTeIPZq6BdZFVemNbPbkSx9rH5
O0hVfamGtnm+KT23XmKu5xesYgvGEZkmP4bUSWCQ9bXYnudqa7cM9SmxhNQ4/u4Wbyg/Lkp5zl77
y5RFPqYUa3bv3067Xb2fL8Osjd0tflbuQKwOnoOo8hZu8xfYjzpRB07eDK+VSl16H9xV2rWYH1MK
6CUc0JnvWgtg53/mPpLgWmw84bvLlKAcnJsacq+zVDFN+JiJE905whv1BXNpeCUQqf3/vqNHBP8J
zsJh2vX+PP3dC3BlXtO5OSrgwo5kFtqv/rwBim4GyxSWsXjtN7JtXV08fP5S7fzftvFnU32ldEW7
eUi0yZXCnBJw3Wa1rbY9riRjOJvyqpzoMo0lL7nGgMYr85NHM9KaBnmQdVpUq70wuHbIDSNLxHcz
4I7hxEgo2v8YubZjrIeYo6E0tq6VT8ZtUPg1H2fQJ450Mj+x9cpBrk682MaRxiV7l5uSTRPIYiy6
kqE3/kzG/cG4VPNHQ8Iy1z2UISNgR65La81OQqWcocHVAwsbJ7UrKNhjTNsENAylyq7Z2tC6Etml
eKqIelrQ3lieEgkadcL3fJDwNUdcyeNahFSPvjMzzY3vle7stpsBickZjvtDMm5bc1mN3hH7yyZS
E6eIzBzoW5kC/gIPZWtl9o2JLec6bVO6O7oOMr/aJ6nzCAdVSCJRaVJlFbkRha4U4ONOBByHU65q
L1EKiiez7m5n1LjJI6VVvW5EY3zd4ZIGymo43Mo0cHzMnMiZ2lsyQmo0Q58c3QfWbI2xKkf8kKIO
FBbupMt6lDTxX58aVEzPQeAgTNcnxRuUkCBhuL9dzzaS13A9+mXIFvgfb/Pgy+5DZ7Uw2w3OSr7i
RiVx+6m7E0nQ/laqt4ZP1xTLyLiYcJNZHJ1b8mzYAK8juZ3n2lreF6fDdMZexKz2iftPeRD7vJbq
opp1bv+fnNax4lieX5/2KDT2+se50i5WdgSTPO7/aogaL4Pe7Rrc0TuIcEbt5pmWaI5bO7pfNAxS
OOiCF3Z1OVCEh8e7mffvWBG6WoiozFj3yteQinOlu/6mDhtV/ZxdZ1YLIHxq/Lpl1lJxZ/h2fCC0
furX1pCXZIFX6DsXkRW10VXtYR8fMDXDGaIvkL9UyAjQVCKPbq6cFeiuIDtJH29Xs5ojizgOGObL
VcIBTa6CR19FkjSq6uHw5F38xW4kyG+B0QmPnYwEQC1L/Sk8ZC9mEFw59DWyDHvw9IC8RIvJbzX3
m5Az/2ReyW+xcBJql4SwFNHPChMP08ghwKMU/iBRRe55fQgMyUnZcWJHygqZSrokJ5NT9BpJPSda
5W3GKfQCpxgCZOyoTtJrO+t4rK7lxRUySUisSljqioPRSvqlHzfQTTO6tjTa2l2W0rWDAq/sBvSu
QmGtPB7DNsHdErKg6q9FgBwX9IJW228UZ+n2sUEF6sl53I5MHgJ3L6vRi4T9SKZJOFioZQ0n77NU
+efRKRvFy8Ib9qp9zK8jGL0OPBATivrHKgHjdF8dcv9SwtIMGM+9jlZCIeA9Bhe1CbdmVK81p0T2
fWLQzJHzi9AV0JFxqO1DTPzbtunAwFF/GPT10oc8niMnGong/CUWmcYTadPMNVo6Z+2nljx/P7Ih
0FSaRZBAO3BRGaUvgswn+fzg45HcEGTtc7POtbzaTbC384/GJsmtZ0O+uXHYBgVWAN2pj3hkBiYs
WGr9zWwFrZvd3EzV9GYUNdxGbgeTipcJdBtXq4ApNw87sO0tOAQubTHTZk3p70vVgE/Nm8elCBsb
B7CA92+VQALiOhfTIFC8ca3szUuZV5TnW6Mnm47sFXGlT5oxhl9SXlNi8dbY6J4tEv8K8xR4PPPb
h4Wr5hFHmiP4ECcSFmFG4srCgNPVhduUpyYTWq1S4qpx4OO0SlhpjwCzJqTq2R44GtN0tKSIwAkY
MCE+2Gaag8P/cSEoUQE23Eb4EIqfeHp5fifT5Rt1rqxMOVBHx2iqyhbNEWEtVgo2zREONaoYivMG
D1C/2rCxWsI1kj5XNDbJVc0qWvNSd1zCd48pD+MhJ61FBAEsXV83H32DgBaoo8AjWWy2eBh3g9Iq
9i6gNkTvvqPTU6bUNXGNAiN5xKjBYXV1IEBRF1dFtTdKZi+A8jVkfMm/hssoGJt+i3CC/RzKdCpu
5XgUw3bmtZLUwHMYnVwytbMWE6hC0ea+6eE+LGWP2Eo530JRP78HnTDq5kHfyEXO0v4I5aRDhrHw
wqAtRcRMv3ACp3UZWvBNMd5QP/KDgSM8BW83i852xgcrzenCQS64DJylYYApwz45xqjm6RgIK7lo
LK/q5yqnkeFshep4A+fYrKGXMSyHTFGZjr3jL5qGqDizZETNOtybIOkxB8ks0aGNUCyoaDLAywXj
T4luFOAROo+5Xcup1q0Nb/TJjOBTlaEeKOypML5rkDyURKLgoF7ZBwnMkDsKjuHwq3Id2RHOBDuD
lJ6DaWMTrNJ+SVFxsF0Q9XfUBzUrYBC7plNBQUpETCBYEJk/nN7AfXBq6RiMpPNPO8sgLrLsmjju
LK6s/vRq5KEKPIKZaF/SPLAu4RZCP7p1sMTWH+ThAGPlLCeqF3ciiHL+Dd3+9LPbcY4i1DbnNyR/
naIsU4kmsWBwjkBNAWuP1c5qDzST3FtZo7CWAIdXb2k7nmWyVsSPVvzuLMrgmOvP+kqs1NUmOmnZ
QRwV2NfD+3t6D3WLk2CAxT+5iW6eVkN6fwnT+qvUqfNzoReKilhx6Cf+5mnyArV/fQlc4fILHZz3
mngOtO1GVQ6TMIZN2T87o+9rls5qDWcBt0HlBKJoQDiDtphlHAwY91/uC2BaZNtaIuZ4Z+KyH0gV
Je9K9UBAWsWB2xRYUpuu1xB3Y4lJxgJVLEzKz+x+lg4ityTLR4pI2sdaSZ6F+MeyR1UIG4CJSB/N
gEYw7xcez5GzdtKsm6pBDivWZ4JXywZSDQ6TBpa29oKZ1Kw3uvP0rTf15iYabW9tP7WstMKGq/G+
tbrd70tBpI5gEK5IA3sAtWUdXoGsmFg+dJBWPE6FoL4rGlSUJAN5OVzCxYHZh8SEdUG2DrFUZChE
SM7btbTfy026uImkl5e/om/p2+Qpqi1wwZYyKp1XC5m45BoLs1Y41V4HeQfiCDZ7pVv0b8rVQdgl
w0p92VYaTFla09VcvWP9UtqClHsje2BZbw/xYgPHCYiHNgYyANSWhk9kAa0aKktFHJOO9XfkvcHD
mECIYOGFqRVthFt2VDXRIB42qF3mDrAg7X7r93wCFdfhra7ctKoFLkw8eLNS5+tShT84pLnM2Q/2
GG/zz+PKbP9h5FN4JqiTbhsnBaUTOBS0Aipa084jNqaIh6hHaGEYnsUJRnQFZEUo7o1qa6ptaPKX
q53lxtudqUumJTd/LfL9RESPR9QLXilX+taMOfVWGOzxauPRLSLo4EYWEwKpe6MlkTebCL6N8skB
cB9LF14qLqzeQfGJtragWe8PIKZmNtClIbQAkzpu0aIzOPJXxnhlKmGOpCBLQ6/GHgdxHMzf/GBz
ppIC72i9pBeRDX9roI8TJCyS/AiGkqDXVluaztZlrYiw+orG8Kew8LZXBj+51BuvysPFwpOGynZJ
c3y6wrOy5QW+YyCxhQMOjHSm4U3XxgFiV7dXXRCXifiFjzF919gs+oYbm9ARPTXhrz8bmsmw00ot
Op6W6uPwm493SqaHQqKraDsen8/qdaPGKdw9wsDRMCSYMtrBlHil/wsjdQOItOXDAu1NWffosRwa
zNkphGhmFgb7MW6IqNkXEnVJaM70U+/MqcV68X+2GqiT6l+woZPuN4iXraIQfVq3ERN1dkeKqaIf
kRFiMcD0cXZ6TQ4VG1hC4LUhek28OL4mtULLV/gcTuYWcwd0V9VO/5R05qmYgaKCKuGUWlDH1cnQ
Z9Xw9XyISHrf8/Hrfo/A6SIy4G7MU6CIc5Cl93WENiKN12570dw+3aCSsy+ROhvnZg6nrBIhKFS/
rJ9Wnbh1L5r2e9ZM8y4VmUAZ4yJX8ZUOOmuYP+Sv78Jp43h1pMJ58lR7QwoTMZDX1ZGRsavFOYCP
RUTAsmx3AL23lFyKgMgaDddOq4OqBP9OQWLYTTUUb4XmXwXzafsBGRC6myNKbuudM0t8N/RXtFIo
cf5D2t2Nh3Jp1iGswjfU/yGHdxJRXbW8zrzOjfHO7bN8KceySeip8Tw0ipzo4aHvn7Jv41ve5qDy
pbcNVy12K5VRPeU2miguGnWVBQ/uSQjiT7BBIxaKme22CcsvcotlMEfM7ZnXSLvgJfkzzdfAtgQY
UHU69JbwpI00wwFKbT7MmEls3H1MTKiUIzEQ23HcDceYkbV3ZNRJPcFikbtUGEhF8VWwVQkdaO7k
6IpFPAeS9mVJNy+vF+vbcjt7pWpCPuRm+jm3reeb2Me50mTyyszg0SE6qtRPUkKutV53GOL5Gg2U
3PlkJh6QLk98AD/Lg8lm7k2bEb3hlnrT7KCNjtwgXL089uintgIV2NCOjiHEahwbzA1HkWD8AVFN
JfHki+MGzgtMsUJrejNBZgfoSQjK2K9fvBOL/294pQbSYpmVdS3GS2h3nHMwyJnqR1HxOzv6vF4E
ZnnhJosgp+S0pbxK8Yu9di5tgQV5urhVYRIDZD+ypnrkS9k7/8h0/VT5CUJHyciWhvGJ3pH+QP8C
AZ5UORZxWu5WQ03USlOL7OdFetx9eXO0MUqk3pa3znH21OI1rwAYqZNLO7fxvjM9yqZyUXrM/2Or
8OGnF0CHv3b+f67Dep91GNkxMBByVLHCBQYVzBBI781SnXgPgjsaffSEra3D/Nsbfe8T8XUN7dlC
3nBA69t9pTlyX7Ifrtpwxhc5mzpP8qGBIgfgHJSFgaMJxC4iNd3j3DzijjmU24zKqfa2+6jzQaRo
woG5YYwlvTc4xU+MDIyaV9OT1ifCyCLEE38s1JVzyIMXWhjXP3hahFmwZlOkpysaM8RL66lqkEe9
8l31BfLUGnUNQ2m3YU83Jq9DOrJsytcOs7fDksVkVdklNUoUorv42DKzooEE4QR+N/jCunNGlftA
ZZCg/iRdMf9PrZGWvL3fFWxEe21d/xpzfBJD2oF9fPg7czKLcblaf5oefPfGXDEo/0LfMXkctafm
Lu2NV2erB6Sx7vSKFpTDsgKZpdXnq2JYc4XcFsHROCHPR356KOEejZhO744dIIkvpKYOF89DdQ/L
BZnCcFs8xi3LUsdetEh4icHD6gpKciFUshR1gdgExeQ4lES8ELcFmr91WzhdWJd/AH1MHHvQFcMH
yDuzZrOo78VrfFEwYtloA1B9YKcfhaYRRTV7+h3sw5rpwFaphpY3ThyCHWWQkmHC8UoY4ftWzXXk
1LMyfq0MIon35uI1imGG3TNeIw7dLhKlq42KAQc1v4M+MA+cx4a3AWGSFaB2HgJJ0bUK95CtPJPR
r3tvKR3ayjrJywmTiQ5wgFUFRKYgISL+47TIFt/r1DtK2GUvew01IIuhdbdw+3IuMYYolR9UqLpT
Tt6kLlIxhV73D7s8eFf1TKRosTbeIkAcqdNUb9pj5lH+9K9jdOXfCB6dQXXiABmwOf0NhrrvPn+Y
A2+TDhdnJ1ilKBECmhkPmjt13uGsapRoR1fxOmlAhweykl0Ap/RC8BMiwdi+OJtaiMWc53CpLE7V
Ps2EPnP3H3brRwPw6V2G/W7bcUgA5iP+0aoCEbSNllzS222h5auyyLPpU5bwW4mJgHuW4ifzMB2j
Gpo4GfEKGsReLbu3iMGD4Ml1N1iYSWecEXKNA7DDC4aIiPpoadReJT88PeipH6qapjImnbbnHKRi
GPyDY6LF6Wj+XhEhB4QHfVtmxaLImmi6eM27aJLK/vd738LXRIEShIdVx6GPebIZzOkjIrokviZc
/9KiG8RJeMdEIo1pthsqWSevH4OjOwrFxxWq2EQfe5b3HHIZtRBHTo/jQh2Q1Pw4ZodEQt3KDm1r
fvQ6qOCIQRthLd7pkfiQ4YZAY5YJ1LjnxhQRQSAvRxr2M5tGIK1IjA7xzHZh3UtQ67scm37s0h6Z
bAac6ktfEMD5q+8HQ3b1NV6ibBTWqwldpbsH97BWd6WK5lgn6CKHUXidbI9zRXLyZHsis4rzFSwO
KWD8SbJbSG8xewxgrue8fKmLzlTI0WNzsYsSiVw5KaSmO3g3z16LgXgbAdb3Ehk7Dw89NzejkHdf
KWVIfObmWf6HGk8yghPlAmALmdXoxJa8Aq+W+plluR46gbLjAWOYaJFmwyoJphQBmu/vDBnMm5Dr
mt+ZmXA1okkPCulUXZgb17XfZxhQsUnsKLo7jbQ2PM+xWuWLTbFTVUeyyGOydZn6dV/Lor7xxBDl
i6sHatirdGUK85Avje2n7Wgme3T/P2fKoMiBEyLqhQeLxvn2xnj4sRqGr25rLn7CBmIM/DW2yIC7
7u7IksyFxSJ3GbFoxh0tYtMgsmtIPeDAZiv6OOnC0TFXXnr6+hZox3d2bsVCNMu2ohL0fPeT27UB
lVpKgsBQEH0vPNxsXTfpbd+8xM9dpV1B77tzrDSOn9SNOw6UbfWuM0kDj9Yq/Tjj0jwE5fpHEXxE
qJPHdkB9tyPbC0BLdcxUuocHE9rXdCc4pVvG3rCxyf0j55+VLzzLjWnCtNI958WVdpXw3ZTeKTIX
ogPo2Z4Ei83TuGvrreEhZAvFvQr2AtC0o98qaKl/Xwijkiw9sMPQZSoyafBsn/Cemj/JmsW+NY/G
HoJBIo9F7/FNeJ3BZD+Xk878Ung394DEd9FgkgHmEAu+1++9Y7h5fOSUGhYG+cIyGAaVrW4i50AX
EiUt5OWRTZzKKlAgVVKyctWxA7Aa9tjBYj28icv+7MVqGihUlpkQkt96vzua6foI/ufi34cZ6P2W
Gh2/bxfBOo4IHQYSxfKry4Hwhl3c43R8DDYAdt0UyM/CWt3m4Hl5NZliu6NuPjZPJ2KmOTTk4S8s
n0Y2oCEoF67ie7gclDmKq9KVhDfDfmsxUgpAXMHk1rXpM+I/n9ww3VgvSSaeySKd4R+BV/UT4bVy
wUxP/8s600nQXQigkmEPtqGAHDIp9SPC6kDiK9Szdb5f9KjtMYH4hJjJgS4hSB+GwwMsNxYu49sg
8eJzfMbZxcuTY6mUqr330v0CwNy5ui2eEBgvUdgxdhuUfhP62exmubqUCZW0GDvK5q6x8pAgkt3A
fuDpVjdvtRFjMY8TCUY1xBAw5VRGNbJuFtSmnwtJXHl6GcrhIys0k+6iyghYMwqgjUDUFYcEC7tg
xFIrHNRZVsNseaq9M6xVItaBd9FtpnNvvKjC/w1LS0keA9c7x52Z+mhssnVDUjsljhXJ356D43fq
wXNn7QKNUuF071RX1kEjYdyyr7CyrQ9jAn8HoSBGtky9t4t+h57YKnCDXzAf9ySSWTltEac4YEpm
BVqjZCZWSpPyTPAsVqY9hIKYa4D4TTsFOj2s96Zae6ylfZtMWtocuD4MvVOMU9bwztfru8S2Zyml
mFig8QeojlQ72schXsHqBD1koLkjvnwpIe4cU7Vs2S3s0pzJ99UV+KwB6fgzZNg1JT0BIPquFgJ6
r7mNF6+OnhCUjiC5WkJD9lmRR+7rUQZTpi3x4ZNAVB1CRR5x2l3JkhHgyjJ/39O0AVW/k6yDYVQi
0ISgroOMSKIOnH2YeoFGl3Y8/3mC2hbgRTyhYJ5YrYqT1uKYpOwABwsDT4YSgmIbPns++lf83i/A
FAguVTuacwxugVpleEBO0FO8nuyJauzrhWCfuTgl3kd5Z2EWAb+u8GpBNR+6WGnhekcoGXVPpsqo
5DH0W1n3H0v4j0voWXHf5X2Dfrs19WqLPbckhtxZAIftWpUsy0eFXaAo46B39V+TmDyJ4GHO87AJ
tf789WkixFdJAHxQ6tLYV+yc2SGHTFYzolGWeCSoxlpNsFLGSuihKBM7BHJz1BflGuLE5R+I4Q3C
zsb5rZpQ137o1yYLmGHgsf/JshdOSpaOWesDuw4xCnfgO7SqOpFuI+JImyYC2fUAlaAXGQWGfz02
evXf45QQp8oYChIv8Ci9zsqk6tN2FqsyxNoppKxP5+DU5AXa7TLUqo/thSXr9ZHHr4y7l/OhL112
7SwYB+j4ZzuWAGlrKHEvu6ZizN6wy4GCv346aO9vvzNeOXMfwhADYB/DCmuT2Eu/WmULMk07g7oq
aEwVDbgGA2oQP8MFkWgPnmxaYJLfTRc/UYLt5MI/bqBaSa5D76np+SZCatEzRVGLPgjCKjPhnTBK
tsX65iMFUvRrrv6ZnpX6DxbuFTMJCMDmvVt4O3RM3gWAREsppLM8vOOq0bbxqlQO6g/b2HNhABSS
o4zmLM9qktEeKdRJH/CQH618AwNvl2azlycEMf8CQtgngoFz1zmAHMCdCzlPdGmXphhDy705zxeX
lcprmKJ5i4ws89B3x+3KpQ8rligVTdhN3b1sxqcZyUeBsDXKYSDwIZ/FgyLo8SRxgJkVQRhEHZdr
KvbVYD9JUvVdxYDzLuXtXuDbee/ZMeZ0TPHjnaJTsL7JIflX/jKJyQpNzL1ldfpXoyDNcj7qIDml
GLkUXwVkXBstvssf9QrnMFU542QZ1sdPi3f+xqtne8m+ty3CdFyqwkB+z1FJGFRDT3FTonhaycZk
wXUIcGmfLih5vHQg9wqAD4K4gajin8uF7GoAEgRTvuULCxXYrsRIH30SqTrb59E1qZlQ64D6SLsP
7Hp8jkk1cGjGbGdtYpUf3GBNKFPA5sEG84XgzTl8Or/J0qSTtmL14cYqDxrHbCjxdFc+w9Qprr8z
8uFGpCdpgtp8hRl1SEOgeEL5Lv+pOcDNWqYzcsWL1RHE5miQTum15GDznTUIZ9BuQwTJPTh1/pdI
uUMyUmJHV2ehnX+6T5bUR9UjWw2sxh8XSi5OhW3Og0dn83r7TqJH0N5tQ1AjTLphW6FDuUP5Co/X
TjNtrbStVRD2IBABEaCm04vZmXqpdxquylfga/UOAscc7/xVt2/8AN/PKU8OQJXeeOoaIzA0zbuH
e5xuV/618FXxxjBQv3Jg6m2KAWfwCYzfAp4x/NS2js7joYDOuZSXu7IxlXomOEK92AEROeAyOKR5
AVZNkxciqkS7wzygKgFf/VFigu7jI6JdZi6o/s1JBNE5CsrIMgmTOSIqy6SvhqI1oPHuTlJDkbch
cuCBmFvcqQYFq8p06XJeaj7wPh1KsrM3Z31/CNugpvH7ea36dbntdPM3KwanSHqH7vJS/Geh2ozW
VmDSo3Vx/1eEVOnZGXpa/Ni4u7GAyEdp5PqBZD9SJFyxSacFP8RvrBDGh+PzhazkNtNFNmEOLLaG
qMv/7j+vyQICRRYnuvvxAzzVgpNqMUIKvemEAa2R1GrsCS8xB7Jzn0hCZPmm7nKek5KhpIyfDJYm
GfvbEyFjXDRDpWJcxKGMmXBbAiCCRMGEZk9M8WBri156uNeR6Uol/HVMcFMk36bdXFRcL8yYsQ1n
Bj/3RZC9wDv1mjPKoqDodC9RxiCzWjOz+bFfgoQzAkI64Sbz/3bGVOVgHlb0lq+nRlx2VjH3TkUC
0LH+K+cjfxsf5DDEz6WXDoIF70TRSMtyWc+bPC+/OGCVQRU2XiL0GMdGSKOHcKIqPgHGFPNo9V5A
aMThO3EhHRX7fppLj1PkaqToBJb6V7PtszKLa+Evi4yUwtOLxmdmOfPSJuMMEslqabzgbvdwxXyl
czw0DON3E1VNo5tmIYkV7gXIbRapwFMSFR0SIqQ4Agj1jjGwAd/iu5vyVWyl6qj0vcLpULcdlfsi
n3G5mf0HsyCRF/mmrTjQvXsJS72L+ZEtk62c448GeyFDKKkge8hVfKQ579VYN1B7/yp6yNkf79mM
a4UR5W/jwyLXRgaPNFVNtof/KYMU0R/p9b3I05aCFCcfqWuH3ditQMC9BJHHsJhSvOvPc/g4HAOQ
cFCrjo+2GbdXChohVVaxUzrjCcHkI+QH/gzUKqZAPIjMd0Fhs9XZueMCxPNqCDMlrQdIr6TP/jF7
ZXEOM2ggpD465zVuUfvkWqntq7nkHC0UVXOMctOs7adnGRPpkDPL5QeDSP1mXdt3Cu3Yw04sp/iQ
0Io8X7SWqAQaj+yXc91ht1tIiXX6nlvaq9opQixS/ugs3KtpXvSk6ZREU962GRFo+cayGJ3w98tD
3PFubmvr38dvaHGP6aNDvwy0xNCfyQzZAm+uHwg8mMP5erP+UoyIbYzsktu5mvYNFIorQkT+hpD9
kAvkoI7mJPHItSZkIWRQUbS7TGGGali69u+RpW4dwc6URVpFUBsQZ5w6Rxnv//ihlvNRPyisz+Vj
dp5ACw1tKQplyirAKkv9BqEQ2a8LwWEpVrGbHzoDzj9jKEQgiBQbH3zAdhpa/Ebvz6Anco+jD6RS
4Eyp+66sIsNTT08o6heiDGXk0dwaajEqAQbGMqSzRQlhVl6p/+Bgrtgc8kUbzXWAatVHzSuuN3IB
uJcankrLo/b+YVIrf+lf31dBdGWkCButvbAfL2nwH986bhy5OJHj9SNAwVCb0dTxiQY4CQwEbLP+
qRjTcxFPJ+0ZcZZrOGiV50ZOzlJbo48t/r4nfB0UYntXa1JxgjArlE0gkyrbzDOz0yONySmPmvM+
498zNlAT0d1Vc4ebeVQKhdBg4jRNEsLzyLwLRQ9Z/Zaw/8N238BzV+uonaCnoZCkLn3pzUS1UrkG
R0YB85j3pBmdxO7kIYKBK74fgGUxjOoDz5OAf2zWyGefxQwXF/UEhuJuoBXOpF1a+PkbbaKmJZfv
nIGHqESTqvQRkix8HFo+Xv7ccScUOqHld9NmFg87dEDEOqqhNWNWmjI2S/2g238svrNKxuKCHSaz
zLxUPxEWIDY5jAyBpp6JdW95CaeEA0Fx5lZZjYjuvJNGbZtVIgzlp7jdq5eJZbR5rvyddfEu96/7
IU0gZ5NR85T11g+vKFxR+0+6Tfi1e0Fce00g5rMbL6UgDnU5TI/TNFiw83VtG5+3oaNUlHDiEgVT
WHBN88WsFJ/ePbDJ59nW3LluFwKkUCv6FcOdZse+7he+ih7HaH5Tlltly3LkQCSetltE6HHOrFQi
1Bd3kE95sF3kHgI/3c/TNXdg2c6KWooJjYwTotyMuqMejB0C+qU3LNBsepp25C9gsZV+nV4bPRsV
G5c0T7Dd9FOlrRn/MqaszXvC7/BCbRoL5uXw78/vOX1LnQvN3ZlsRnJ4I8vUkJwOE50/Yj0wT0Nk
TWiLcH2K+fCogccWkvmW27EX/3w6vD+JPmP6qoL/0BTKMHQ6G1DYlexPo2myqFtlbmXSRpFk8SOO
jjbmG7LQboFD1WpLaZM2tAJ8PZvgob2BkWGj484YdVvMTOBptX/4KZllZYJCj1AogCiilDCIrNzb
mgD3xEdhYrp+M9caW6gyfMu2E6uwJJ6+cHq3XsgcD4ihHL9TbxfwqN4zc9SI6mGiVD93XaITbaUD
iWdE529PwpfuwE7guyWEEMmrCm1o4LkmMzye/yOTJiG+lUKPt4uh0MQmpr1v47ab00DEUFCQip+V
p+OKrKNYbERv//IEaaBuBSGtW6lO5LiA5dnNACx3P3zk6UAotgjWweP+EcC3XuY5lVpXZsfm/Ioz
DPPGeZ1cYBwFGIFkbm+r3ePMXtFkOBHDtg1o3YLE+yqT/bBGa7Qd7re30HMh/hDQGvpAUjEwbEpp
Bq4yB4d0JjEkZwVdZqrcMpZDkjztsKxWYwJx3GkutROvmSmW8rcJ6wVuOYCHuAySvJy5mXr1RA+r
6cPsz5oNhCi1rHNxTLeBYJjYDwSeGmc7TUJcm3R7UJAd+P8wZWw31232tu46tWwSSMU16FyLLR6+
8eUfYmG9B+PLyQGB/oFDBEIEVKVA7L0rB2GMcScUU23CocM65ppXbt7NubW1wvn1CXfMZDm28KSd
FFCq0bhy89+cUOwsm8T9qtdDFdpGu/fQZlkXWX3WT2zvvSwLhLndMDle0xjOxkBCNSpFVmQ2O47k
h2elkqYGbxvU7Xa02cK+HtXxYR6enAiofEp3sRna/VtxALlCx+eTSGZELFLVz55ARIBTojne2dTs
k9b79x5Pb9EhbpOjgWiWu6JROoZhMoTP+VfXQpStgPXaXLYCIetITtt9RcF8KXpRkETskgv+pOBi
3WIHVzgpT/SRiAw3UHJ9T8t+vmkft79mnT9HGMII8ySTdP+i8C1cBWxZisJJOhqykwkb5xChsihC
jEKq7tX1Ujl2d/Czf3AQXdrJ57yaZpxrDX4rXK5k8BR/EYY2nLzDiOfuZSKhkNhsWq7z2fYF/xVN
+1z6aRPyypqOrhXgT1XHopQniJe+dsBurf1iSrvstrjrVxwGo+MTtryfnDrVrmMprV08Ny7Wwc/P
dE4+dhjqgr4whJKrcPLDS4AceOS8ZQKeozeEkPo5fdMAFnjS6Y/Gf0/M2Jq43w3dRcHYVuAgHkoC
K9Mo17XQnnu97fz5eIQ6qHZXR+UG4+0uyXOa4+AgbJeZSqEsbteK3/0qLL4qz2QBPOIGZ/LkZ8RZ
iSwrctrFQ+K284J//ogjWqmhTOvZsISiIH9dCQ7MKgBoJQV0NU0ugtQI/7BEVhmwdiXoGB/NXwa7
AI3kWe0tTcCzMirasQzmCYgc3Wp4uTDEY7q483QKLLz6H/7k9rt4lIigJEEBOtz8kDAQNpjUkiwo
0VuT3ppNKH7Y3tTlQAfgvnUTDxMOufL7+RQSPaMoC9Z/7wR5/OWfBjW6M8y0dmp45oNRO2RY6M6p
og1BXgNX7loFvQcry8OynPYO6B9ZThM6CBi0iuQT1Yilz9AF+3gY9ypWj4DsQ4+cl/SotEFTbtn/
ljmaYJpNjltz+fgrSyoaY5DQr39vernQflzbo1RD20874tSQ/Otp3CV/polT+K1qYO4Um+qbxN2X
9ovsx5BNkro7s65dDpfNyxa5jL9D/spn9qI7yxcG6W4c6pshHa6dM21Tw6EiK+4/ARmynltkn6WM
7BA+Xc0+rS8ZRhM5y7nYckKgvUR/qsx2Amp5JXst+37PqZdirNXmUBMqX2/iUtnBdzaakxuaSjUS
95ZKxgQfqwEWlCN4ezqg/5HBgFqWLyX6wY06ew66G37a677qFRHdPCkyDPaygV/ZAn1wHdLbVKhI
Fc895tJYbR8sW8JmD4XGywyzzCa99ZLYgeMK9Sq+fzBYw4pNnLnuvCTCvBAb2YfJGgoPEgJUKhjo
oxZQERR0bS6c9l/KsGl5B+1dXb/1oaGmkkZNAHuSEZU0dbSwWKnsp6IxbeSGtTfdT0y7ixj6/uhR
BmzTOcZS/JQJWqzfFdyTnC1CeBx3k9o5n72M3fPBrLgljVtVI5j7B7jIGQu1f6YkRLJi+i8y0+zK
rFfLHqhf6A5MzfQlBmHD7Zzf0uQ66kjo7iNWKizjpCZwz92LCh46xhW4CfF3kKQmcGw4d4/3k0EV
z2V25CZJE6D9MuRtRUtZHim4VeMRnS41ThlMRuA6jheV23/e4xiJY/rnRo19tX+bQyTlKtpxqkEP
fl68tgFdXOxdUBeDFW9HmasHPZAU6kusB+qz/IkFRH/LfufTEhpfu/jwU/MFIL8w/Gb9cKSu6rUR
wrGp3DmSBGiZczyOdQ8OjVGpAVXqBkDlWj2iUaqyE3uD0GuwlTVUTDCF0Jqzodv51SKtC0uP+I4w
463nL6vgCE0Y6OJuZZdEQ11HOG8bVaWQ5qiBFzfm+EC+zIKQV0Gx5g82MpMcCTF4lEHyk4y/cmRN
fQ/K8k573K/GIt60BZgUjydi/YvlhWvp627Ff9ZmlptabdX76Xu3d8kdNL3B56x+I6buLpXGuN8R
iyOriCoZ68uJ7+Kp2sFo5i0SEjWXhIq23pNCUe8EDG3QxsL5rVWZdjeH2bI6d+8Zup5skx7zGZJu
lAVs/hK9Hxkj149oo8qo6pfKzt/UgTSloxJwC6wrLA05aVH+KjgftYikV49YqDIgRM8o4RxfXKr4
njOOS/m+QTXuoE1SQhDA9Tr8UAPn1zhkaFvzSxDMWa7+iLa2ns2aaNVoZHdw8V/r+sYqkBu5RKE7
LOGr22VOSWuBE0+SMRU2J8z5IsxIr3PeWaOCcGTiABfbGN/M7egUjeiL+etCEP0/6K4M5cljkfMk
vq4za/eW7g+QC6WbpR0uFTtE2ybmm++2QsQ6bu4Xcc+ZayNrXx6WPrq87wP4QemTNc6VSrmiO/3a
u7d3KA9b8oChVqu/mFxsk0/P2YghWN3j7AnKhPtgnoGJn1R/qsjOQ+9/Hx3lLBah9cnGKj3tdwQh
Pj1mDzYJ52S3mZELKh89A6jvrbOFwVFwCe17w5AkzHOYtnGJlhZJzUHFc77r30YA3IEp4N8iUyJf
Fo/sUVD4namyC1ZFnQtQF4ieZ6qd4TzkJf3OiUAGkMmHnn5cHBhbIgf0wuNAdy8ktBvGd/jzQ6Rm
GFB4BtJ2LyKScJaHOxXz618z3dayqvFQ/f+01PNpch/NjSCfrqtYdlUJ8M/L9ck1Ajokr+2bnEr9
Zjtecmfe8snm+UxGYqft7n4OOFWofd+YfgBZYp/5F5BZsNRjrzbFkdrPKR5zQ3sDRQ+Ah8c6ntwj
JqzPwmdvVNwgNsLmOKkpa2EeqzD4Ce+kMUOow9tgEqWtOAGZoGkBsg28i8R9N6RQRlG5uhoEKt1S
Toq65vHN6yAgJUn43ppjGlID/9LwOb2sxhcOmfH18jTErJN/08IhUpW3lHpyyiUw0KzpgFxNNeDn
wGHzR7MkoAvE7vmTEI7N0ZlAsRDvrYlykfHU5h4t/fLOA7vnmCB5XiUzSNfH/8rY+kmLyqiHOo8+
oT8EjSobgfheo8M45tBf9gnhd5IDewF1EqdDc4vOIm7XdXENSnWU+eEou2J1gMGjG5vEvqc664WH
8w8vW0X751DLRFKTPO+zQnQX+251qbc36pSEKipioWnu3ZNlPnZgwD61FQfoCKy2GqKF0HjU9oNZ
0oLkSxLd9P0DU6Il6d24BPg/RCkQp58/TJ6REqPU416QW47LXR1xFRsHkK04DKf4YbviLX+1HzTb
x74OHY/VWm5aFiVkZrTWvTLreBUBLc2zUxb8AQ3mjQKZReSAscpLE0tG4m4LLCBuLSlAM2OybFDp
M5bU0SLMtHUdWq3llJq+IEursJeK4cS7j40eX1XWoxEOJjWJSUMvALVW985UWabsuSek4jre19+/
m3S+L9PepVAvf7op4oHAwB+iLkhoNlhl7oH2YYhaDl+Y/W+MnEomKVvsHsNtf+ul0QqVuezZ1oBP
v9e9g3jAtgxRZRf8cRQDxcLY7UPK/PBUN7SVyISFFM46WeDTnUtpIgPvv8LsJ2R+icFdiMXkmDJv
rbAEXVwwQ/SPwv0zZEH+3phPOIeWI0Gs/WlRWNS8HVN04xY303jM5oaMIEwuWS4VgdZAPSYhnql+
bHzoVOChIOplb7gfEQAoydl5MpnuY69+OO+mZQcRBlDCOXwZb+gR9vV4uBVgFWNida9awKDbBX9G
VjQWP+PSR/TWN5Sy+GnziJsv1Ztw1PO59BlX/+G2C6Vzzm+/0JdwehQ1umAs+ApO0XjruzN/4DkW
TucUJB0GrGCEu3CVc0YCIRKS51DGmz2OypA5cBvcWx7NQk8fyrerEEMeEaxQ7kGof+ssgDfHO4ag
BXfwKWvGYigukN0JLffBGfYGJ6YZ7zRal8L6sPiahx9pY7Mz4Zhhn2OL4E+sMssAQsZQIWHTnLF2
LLdL1j2Q54+n34IiKvmm7T+WWDhqgyRXuSA0WOaM1KjaEdPDo6grCivujMO+uGyU8DviExV0zeef
3zaG7f/B7zUQj3w2cbZInmJktLPdRgHlkiq6IQn71oX6kdxohSXbNRGTsQhTM3bFiMaSzJyWukgj
E8S8QnZULh0S7Dk4TW5dvJAGmR297sAaWvqwO7aVkZAtzxNW78avLouwfa75ctnJPV3kBHWbjw7N
scR6Z1NwJhpYUm0n3e3StMXUwmDONVRoC/z/AtRIhaw129RueYUhn/omX+jhKM8PN8Xtlc+jVuBm
WxuPZUiHYH5CyoUWzbkEV+320j+nQTz4qDm9bl9Li38vk9uK8M9kh4C8HR4AkKnWYanFHQvxjwpt
t2I+vRtZHodoyKlTHHEfEla6D16XA2ddYZVwUYJyu5rj3bxuRM785l8QhdsSBdZ3MLhHRoBlNvMt
ceKz9tnPGMvC/3z8mccHOVog7UcNNQZWmrHzyXhisicRdNyM2R5vsdCqjpRNJo/IjKqp2xSze26n
f8KcOjWjUoi0ls4qc7ki+C1bX+aTZHO2s8QyLMA0aX8r/UaePRFgWN38nRIUskT7oO/Oqdps6qCV
0TMpdxTYPU2q3rr1OfhVkMa7ePGBaY+hKFSVQBkOWVDNawNz6wRRqyeGQV7BMXiMEAFgRMcbocyk
dmz1Y6i7URKk6Fwx0aWVRSZn+Lqqg0Tf+rruHaDallaQREis7txXAZvH15rHAh95rqD9trn3pfDj
03t0J6L22FpuObSVjUIXIrj2KR2XbmfHuRUNb3IEoFH8KH1WNHiBhGYMYxQtlG4lgArrCQBEfeAR
4LFjRxNeM4ke9fdENuYrCtbGv9gTlma97onDM40mp1sLL8D1sajuuMhqm+3MmC17MjhZFECBXRp4
sPP5ifLUdQi354l2XX84opAx/VWKpRS/5M1gGpU1Y8iF8RahMO2wSIpmFtUP7Lr1nI1afCQgNUto
Merq9lLD7wTYFoY5dn6Tog9rDzUPVHfb4RQqVZdcggQBiRfV+eoNIF5fgFLALJR0elb51d30PRI6
nYZGRIHMfpI8paD0m2hK22aYmf+2kl5w8SJU3fsD9qGg2wRPEBEf1bCmRKOjcJs6ZbHVxKiOgtrk
qpJ4ZqZOJbHDJBkNOR2b7nBE8By9dxprsDPbSUymovjsle418GS5SkM990HX/sDzmAXroJL6uZj3
NKYErKKgA1e6qkVB/2/XCr3o5Xpvy7WMlzv8OmeyOCb4pdLKfOXqVu/sdBuqcRDVWCAjWSgekBMw
lTId5nDLt9j1lpM0it3l6Cc1CSwUOvNcY+4Bis3fz0k+kpUKvcWXdult9vFTFTLRPCqg5hIeNOA6
AMky+jSr0OZAsi5zCxDj/VFMJso6s8nFvwACPCaQhLhmQBXrpflYLGJLhAgMSyU8TnDHUwl/nz4k
G3mDEv7qCD0Iyyt9YNsRNh/K+R6u7JHpqWWZ+TDw3sHzJZ+oNqiUU0JL+s5lqb/Hvrq6RDrbB8Ub
AOHDExB9F7txcz47BAmHaMSYoqq5nZf1X/aAefpazxGUmtCF7yPtxvP9z8rq7Jm2bt+EeZdvyiGg
UTqyRdBMwHqYfTP5/EIPqZoLWtGHorg7MZBpBH/AnM3mCQFkqNpctNUqoVaD7DSZmC9l60zLqeDq
xkK6hzIzTqX4CWS0uofMw98dIDtc91ZI0J4j6qtjS6gNUniGXyVnbYtVP+1rrSPMR76xOzZufnXt
lJWhH3kcdVdqYKSfZ6/nJxZr2wIRNneS9/KiaE2AIeMmSuSB8w3AB/PSq26/dM2FYe7QHSwReB6E
l+xsQgKbrfLtB+qB0estsrZ85fVfIVPArE4mvye0env+S5qGA08qUS6EnutRmKt+C5R9XJmePlAd
oOEDFJpI+gnAYZJH+itLjkCM3xs7UcaoAOz1Jf5YMW1B70Qym/ifoKLBXr7AMxKiqWKUNBgrTAmi
0i4WlMM2GCfqpgP1m3xW97tMx7hDsDTwfTgomeYQ6I0WA+ye9Kac1jANUPOogA1gVlAz4IyC8xYr
+25CNFWHjPRTAwWGs4c7jkUKyjrnhBMY3SmLgoUcwKgveKfj+Fznzum70BWIbzvi/6lvAz3dmPXk
TGiAfKyF43PhbTm5LIUXMbbq693I3st5UDY5xVgDWNn1RLkMxhhDcYoshPzCX8Dls8VKW9i+ctgm
X++i04qY0n0okeDlpq8pvTeLHHDLSstbnkfL0hrdCoy6sMs2fM5sd6vHPFWUMvxCIG4Eo/5A0fS6
1s99IbjSsGRadjT0SPyx3fnruP7iM8Zoa+6HQUsUcm3g5r++chCLIzK/K8czrZWLE8lzB4aGqZM/
W7G1YCou739axSrE3PCX+qNP+HUzCItL6+ZbtbT7rxN53kicf1lK/6mNjFByg+ZVNNAsNIetVpBP
0an67QJOe186INf1yncEVxChBAouhTx/+kaoFaoOfYTlexXAN854eG67xPo7/h0H+nBzLNkVnLgd
/XRLsAhJqR/WY9oYcu67wFMrrdQ8aCX+zYOLzmKV5ASiNnxlnhSmD27Tol0Xw5d0LygvF0Aa9Qb1
oFNLfoGuG+zncZ0Tr88CsHNnvNAmmGYeGj7ozjxIx54aue7vRr3Mk5dNYOfcfu5uqM65ksMAiXMh
8agY4FbydRI5vFW+R+LY9zdrRzUz65p8feA2m0//0NAJlkXb0WcdjPa8wj2Zys9K8Aoi5TY+di5o
slF+v7hwbgD3OA4x0onbpb8W7jveP1wmMAZ5qMgPY7Afkm84ukeDsfkcpiYt/QcBmGUNXoF71/q3
IhNrDyfW9bZGhnWoGV5yeJ54eN6GlIjxM+3fHl5LUcz69CCLr927xqIJmHVrCnUu1CZ+YdHftD6t
uU16oLAPVgU3lAXVI3rGTYfzWpKpYeH9q70J8kRv0vWyKyBBGP3DPF5oqB+DTSlueyExXOboMFlz
nLd0PkI4uCg5RPU1xXkhjmANQvVvSAcIlOreLv4KXCqWp/KkA33h0w6CE6AlQuzn41RoeWQe0Yfh
jh40iJOmsh3GpDloLe6qNmZ1yCB808lwIxPTxLoH0nPhUH5s858FeiyO+m/jXj7vLhu+6YsYDMH4
GjRdzWvfWJCl1ffIjTMmnWoQZ1JCsoiBuK46FcPiN2Z8oJV9DQ3EtblF2H4bmurwTtTRQ2P1HhDb
U4U6oVyn2rVY93+TMnYSUQc0DnHpqbojjLXdE11PxOxnhjmjekcGVTDOVtCkFADvRf3Ykxyn08S2
v5pUIeM1pYGlm56NE0nsiRYCHvTsc3Gjy6P3nitSDU458NcmOozWzgdWugJcx5JBkfNDH64a92gi
cXTrnnMLkPuVchFGX94Wxjg5MTqeCgmdZ62vIOZ7AGJ+P3Umz0wUa6B7/ICxKdyssWKDAI7yhaUR
uLcOUn3m48VteQVZj+4xywJb9ydQvZEPRK16xguTS3ALpvW3k5nqfSyL1QE9++Gk2JUquXv/ho9y
ibw0h/E7fe7qCRfw9szE3PD0miTPu5verSW9rJRfpRgOtHGLcIt7IvbdydcsE4XLcF0ReT6PqCrc
nDvcxBnNmzGJTPD1KAWFlZXJIOALKNqNLiUh2ljuLJstL7BNCTkTF5215Hme+FeQaHV2IKy9fjof
/q07wdm5+W6GIwTspkfSb5Oc9HmuYUI4xyVE7gd9bcPdRBbo1jCzjdaHkYJB2piltV29AWroWSoK
b4FVhxmB90vToS9D3Rc1/SDyQMU/+/OHJiwIXt+vIBDMCm6YFNCa3J9pO9PhoRXRRTjV46EO8u2n
o6ne8WLMgI/aSUsUtpKrv3bXXwrmd1+ZqRnGElvD5cINNWXEAj/lhY1+cEtrhMEclHiN1m1yqnmY
3Sx+7x6yzr3TZE6dHRXEI7i3O1i1kjpzYWQaduT/t7GQc9Rq/iOEweuCcZpGI7wh1CLIhmY6qyDd
nHTSdajM9xidX+/Q3Z8okRevrolZJhpmvF93QlN4A5dGgNcJzNOm3G8MSXaLhSA5x6uYkR+ozMen
by6CI9eomhqXClan89NRfSCZwERsNFwbza0UlvmjPqYpWep6OMt4ZrpNP15pzanYaBpD68ZUV+v8
UIBNMRGKppjkp5YT5U1I6zTE4Lvol+Ig2fInIChQTtRk0jNSJNYaqHqt+F26YDwnZ5VfvDENqBA1
/JD6aUcT6mNQ4JqRwq717Er3AWmf0nDlZAEAVicEMd+beJQlP0tvaOs6+sOUkGSN19oou8CF0cgP
CbJRCpBOEIhCUTEuvWYLWdFXmgphX/8QeWHmU72G4PYAD3NQcwWv5pNCVHtGM0ph4RNlzJgwtKGY
U0PD4rm08Keyz8RCH8x4rq6E+MJXhqQWTG33rZMNKkBH4Q1Ra+IRDpKEVFsci09tgI3EKCDuNxRE
H4BOSS8Q/vHBbJgXfP0A/S+5mCwManOA0RrdgVYtLnXkcyVWnJygIGUl+8ivk0E6VE+98n1jsJBj
DY2ClXXXUuq/gtkLGdCHgdA8Wx31J33+HqnIcFukq3ye2O5n0XAlOdqFEsnUEOGmcWCGNp6LMy6b
T1KobbynHwLoXCJjNQlla+1WrQNPMvBx9/bfKmZ2Kaor82Q/Q8+KK1GG4UDndR68mZA1ibMgSwEb
aNtPMELTVElE1z90SioiFnJQNeXRNtBnW0LQBGceGSPS2cYGWm2F10uMfBknAr/Fyt9WwF/wa2BE
ABbyybuUKkVRjHpyQEouJziuZ762utEuHAOLw/kZAAcW5dLvSrPmb3Ak0g6OWG+onmgOsWnfSXhu
kaVtjCv9X3H4U2BJXsSJzNbq9aSn75f6JsZkKlq0FGeM7ogjeq9GwzXednHqreFNplyJNTnw/yNm
YbeZAC00DSP7N27nVWhfy2q4S6Gd9Bfge7ZuU2XiCZndJQDDvVcU4gBs5jSzAPNkpF4MwoSksSOG
79sFEkiHmhYE3N9999hHOxUpgYlH/CN3ocvSWH8YjgEM05wDudVjaqyy1ZSX5+4/bI/7ei6SrquI
OLa8oaX1u26xNh0g0oEx6fPLF0EZtwtLZBWB3nBH+Pcn87W3pqufmfA7hD1gnegHeFs9R0c1R4Q3
R3dnyJNi/qK5uIYu4x5LZoobQ2bTgqcTsXa5TcCN0oTclHDow/X8176rwud9cG9LAhrpWx5YqnPW
otoM7JILq5OWsq6mu0d8cquTjOVE7ziAhJbZnK7WeNqs4s7CHigGa52XoeVRto4GA8ZO/xnykMcV
dFTnSwer4NM5tf5woCoTCZFEmLlDYOCE2iwhb6EizkpenUxppKsI/wjzhuVD4VtMFBbLKbbVlEm5
N1zZLnsm955qjLyKxfd85XjyfV6jhBfJTHE1Z7GSc4vSEHcS23o7r+UDW2KPlOiiusk8vZMuVYxB
y+F4EU1isB3g72Xa/PT+eV4w6LVyCdzF/BwLBgLZaPmN7BM4kQgEf2Y1o43YsGq9kX/eO2JnJSe0
Sb2uR3jpL5U5rrnQ60Qz0hON4UI7zbew4RxZic8gSKXfKn1k8pz2BYM3E+4PfGXK4yAIX8pg0ssJ
maMoZ42SiQ0/dOqWtEwWcrvjKC652Wk3kn11NKfUmis37Qg+2NDY2qPH/GCuR6hWPUNEOw84GJZH
iz/5hSJ56wa/TlEKfBQH8Asnnefe6Jigkn7HFPgU1Dw5PpoP1NhGVrRCUm0/lJSS2xh+YgzYPSTn
BIBiB4cBnp3SXaQgA7r66HNEE+Xb+EOD77AM2nengopL5D27KaLv+gQanxnW9I/J8+BqTdxp3KDW
R7yvND8G5be9bDbA25BuSRBRSnlxnpPCwt55VlbeXFd7SJQZu6LUrisCO/d+5uXSHhMb3Gj/03Nk
bVqjIuYM00Abs0xTx4K7ZDx1Eg5NQGyD34dgS1FhZYfxEZ5SUyfCLCVQc6gHEuA+MtaUkQNL9OdQ
WySIkZRaXt/R628L6j4TAxT2/mMRxTRDca3YYURNzd9TR93H9JHRDwgZSbcLnKIq8ui9zYE/jDnw
riOaN+kBzMuK9Xr86dE3RpPns25IWAxEe3J2/iiOyTJNktjrVLPwi3X0gJaIwa3rEvPoaBfa8G67
i20xQ2OhmxTX2k5r6Y8GwFwgCDzTJqvguVrHvwWdZskASPpVEgd+ggC5WlJlQNxRwO13iQ0wGcfx
6hsRWbU++DiVEeqUDGKXw34XWTkvU62wYh9Ot5eXYpVCYnYXxh+8z0PZZJJcOoAx2PUWktb3v444
PNJzh6G+fjsMpuyDyhXmlJbfvZzqPAQSyV0vCG6c2hM8z9mlt+IoL9+4OPTrP2KIJzUa/q5HX9yS
kh2hyCHRhu+tEkGtCBigwUvVZF3DGUrYNkbg3/PEfKgoOVQ7vFmZdNClNBsUBPBjuhKOu0WhJnVX
4nr9lzPcrTmE7/91IhVr41CJAMX6LtTPT+1RViGxCqTyED7LtqG2nZYU49N2PYCp6h/J7LkFWB3W
InYONnPRxXYtXB7f6LUx3NgfNi7J5CqscGYXWpmndZYZpCWHsiHXhhMlaw4/4fthACGac/VobMel
8ZJHElR7mYkw/LG4Hc0QmIhWuG0IJ/OTs2dVJm2azXidvCaPEMJk13phCE9N2YpnkJgXvuq4rN21
LHcuAWSHuJxMe89pY1H/U1jr0nn1KWlT33L5q7i2/Jp9RJt/w/dDxTbwI7Rm9KepRV7/2VWd6sx2
dzBwRq3fyL5EXyBnQO0K8S16nt7i2KTDje1/hG11t52iWQEfWc+J8ayEct0m7L69hDGMwWJdRO5v
KJx2/mMD80pwaKjD90QQgxY7iTW5kaiHvBTOgteFC3la3wnMEfJ/Uf0exCxDk3siDIrNbFHdy+gd
Uf/dr4MY53D1zcV5nGW24zMCiUgeCM7aBDQz5B35A4jiPo7cwXaxo8Jug9E95MXdzhDrCl5h652I
vLuVc1piUfgIpzpN3xexpMPQtKUAuGcPGkoEiC6U/icIQr1EB4FoDfgMs9wFY3onelfkTJnp2N4A
HvGTOoDC1d101IoUS1jv+BfUMaBCXrtSLariKJj8pv4/mmw6xemRcWtc3disKRPBmvckImRDO1Aa
RWldV1dM+vSKs2IIQUPpTBnDgb/zlxYG7JE1hxIRb9oCEcDMbduo4IogZn8HH/0CexSwNbm7mEAZ
4QRc9U3Uf3rQKVkumZFy21dW3ArFXgHfnsZ3sqAwYlRLVJGSafiGJnJIrqSUbIy1ZGCI8IMfbf1F
6Ys1qEbvpGtefpnw2R2D2fjGKHqfxt7+AlO3EApGqPhzYTf1AzPDH49j8BCipiPM1xGn5M9mnSN8
XUs5oUF+9M0e5IXh3jmT55L7t4GB2IYt20OMJb6n1j2KK4RTpZXiVZBVT1/MimpFYppgmmZPY+3r
4u5tqfs3Wpv9lJKPh+NnkHeeeDqPiAGG6sawVvAQ3YioyWQobs6LpeXzgH8dwTUGNCKhA0vpf/vY
eD+vEMiweYYx1TWe4oCAT/v+BjW2SL+BZ1aoEwEuHxDcqPJdz164gWuOzZPzMjP13Ea72+hSM4mr
GKwy8kkVLHdKr1xpZbIRUKFdVZBAzaIo5LVQA/UPZpiYbGQE5u+tTtH97JBIexaGG1wIRVK2hzub
czcOikJFRfymRuNcdXUO50QSTearPCBlPHx7FlaoVyhJ/NqrlbvCXosikRdyHgtvKCvwzS8z9wp1
NmT9GiX1+47Qc6Hdsz5myY11pA1e4wl6rrpDCl77lyQrSCWNgEHfqQqnNElrAh214Pxgw9A1dVQ9
Bck0Br0JGiVfzhJ5GAI2K1vrBSu+Qw4snOGp2xAxE5RrrugXxFIfw3f6DaxxcJXsENkiRkDOMPD1
CKBgAaTPLqv3EzUSNo7BKqnlHCWMd5DIvNDHujql5ZiI4qtN+RauevId2pTkhAZEpo5NeWsux/L0
oce1nLt0BehRkshRvemRGtqHUYOkMC2QSKBjPeT3hsOi+kYuGom8StifxEhWxchOElBwBMkHrvlX
KH1kHW4uxrzxi6UsGcKOVaAHo2RYcSpWNLR5QhOZOynXDKPdOV0TqAJqlcUKOgJuftDf83sT4YOu
7TatyME+IrNDVbeTy6rQWgRHZA0ira96+Wj4DXsMYiTf7oe9GSjf/Tc+gBPMZsKQtZuqIxXs3zUg
dZ4JJDm1GekictK+AQ5Fh9TDwXAe9fHfiOh3wZq2W60NdVWRSmDcF4uw5TSJiE5NEV70QxyG+VGX
9aF7HrdT6PE/IBGTHT/UMFTUye5sYt0y/rkP5FW/+hQws18rRItv5n7J87v+Nco7raypnORHyL0i
pntGMLCIJ0LeIwHXeyr3Knr3UGyVkarSiE91k86eGd85GPYIA1G9cB7E0l+AJ5WmJ3IQKsA8UU9t
0w8LrPmH9S6CvOlrrqYoWZZ6viGcO6qe9nr8rY599PIOCk24ftrlfxtUDqBXxpxVRsOjBzn+2veT
CAJO2oFWs5qiB5Qdnzrlf1sKTVCLRtx+qCCP9JqHOyozFAyvSOIDq3tSdiTc2EReHFOUaynYmgA5
UTgEh7uflTBHGh6zvIR5vhB2mG9Xf+iySy1ZjmjWA1wAI6pvKNw8b9G664sskl6WdhqpxZvFWzhc
iWfoewjUayU105xAW1mvrofzgMLINIkWwywBW34PsFX35lQgOojzqOIVnIuC+L5g38nWL/nRcS1z
GtRJAjCX5wyOdakKjDcgASPb61dO3+3jqjthvlZrdfQXL1LHRDHi4FuyMiOR+WVnV2qI92bHg7Lp
s8HtOsJrLVTkOJWqbgEO4ZJDah698Env81MEuA9MnJ34tNYeyCtjE/DxW2TovZfYhnFmZ1JxPpfr
90tsU6WlA3nt2QluKZD+EQYZoLlqGU4b7MUlHAKB/fJEwfXQTc4nU/bZLNewbajYfZscO/SMICm7
L5GMEjXWUHN1a3N10kP3qtjASNf4jZjMV1R2vaa0ua4u/3+bzbpEd8mjE5AaqXPam6OSuXzcfdD5
GTNKhXZ7Dq6b1hLebiOr3pBbxXgLZDKSubd01uTSxmrLencphTCs6j9YFjfLzBMampaXas3/cFqB
3ORMVGfCmLERbv7vfVnUXv5dlpj7buaGUg5jro1y2UGN1u8VuUEKyKgBvrrs/wQhn7PGfSxaUQfn
5X9vuD+q2/tgthWqAECeH4E2N2dj1cP6wBvCu1xD90vRIonhX+6uQE/PmwLaC/+rsLGH8Zao/fgE
5GQ2H7d0Qag95gAuB7aLqMxOx4xhn8RHC8yTaCuHKUjqJCkprfszwwMYXIadnyBVfx91Vv34Tq47
daq3N14yLKFzMdh8wtK8ZoTqqppoJIvuavEz7wvzS2+svGZaJ4bV1RA8x3ua5IS9EkJWcAeDD+Nl
TsAyEnINcHlG7O7mHPlAzshsQ3QnlC0bKP90zlCfAZeUQHTavC6oMwML8GHbz4cLg4361k2trpBA
Rq+cEdUejOw7bRi5bXZfuWWL+k7+N1PhbC2a+NJVruhKPRRmvoQrbvdzxUOUDt2Q2mpr70U2+3SW
E0ZGsHebcf5VRkOIkkehW/DajWspSSYN9V+FOFJZ9fbbiYbFq38x7TMJjrwREqKac4kotQY+3YOJ
ij12iPKGvZ1OTtgQ2I/Vn5TKkpi8Qd8RuzMYD29KH7dlK5qeSzmXdIvHNPSeWOlwllmxyGTaZs/g
mk0ed6m4e7/z0w4PHMLFx3klxHdu4fik+uzPmaOnGR4XPqJilRAANzYKi1/r2TDAoyELkAMNB9vH
jdgukSOgjWYIqGlvEVB0fvC0u+oG0ghg1lRjiKzwzyVIsx4wHNc0wsCA3NNuYbLZFw4ejsBTDdLc
y6SpR/Nt7m7zHSeA0n/Yi1zYGNZL0pnZcB4F5LkfBZxd7eOwmeXJKliqNixFHJrFDCs8vulzovTJ
z1uJNNP8m7pdAwLtclHODuk8P11JRSyhirA/j40BUeUwc38N1KBm40vAPjzOF54bkJwEn2EoNukb
ohgU8DTeaFkJAACuqYisWIzyLCHhVabL1RSPx8mRPA/FbgplVXrEj+DtIj55RRPO3o8qUStB++Sn
X7C++4ZdzddCr+V3krG67Kg2/i5ouY19FQLVZJGPyjGbystO0mfsqGaYtb4++XorM6XAQ675hCle
1NPxTVx6COyjLuDlhtzL3eCrj3p3CNFnE9khMgAy6LkuXgljEQqIvPw8fDgX4SQhXrtlSSWvdOAM
keBkS11fEU57uqgiuSiRXeRyQXHSMPTnvm4o7048lTQgajgQK/k2fNl9pOEdTJp6D7+puaFVhoAW
gMjp38804mpevUug0IiUdJXWwVhEbMNjEfKr4Wp9+KEfo6jus9Cuq/8icJBpT6vg3vezTqsxp1jM
CNSBJ9QUfiit02IktyX/uifYa0IA/k87/uiQyGrv27AxpWNxVT1wAE36xceGjxWfHgpnKi+3ZP6q
qT/UVgtKiE5aA9R4DJnT6FzawFVoKWu4BnrDIqwsBMK6KwqP7ASwbzJzfpb8MZ3Ypny68j85nxP8
WwGcCdD8fL+18kzTp77MCoj2/6zWqSaPFNLWQ1CNaJtc9PlHhBFrGKL7tbDU6wr4si6/om/2funT
czhO639FxCbQR9VGwwQ/kNKG3sCaqyLT5Pd0qO482JXra/EMenUpS+y+I7rSOPuIsNMe5rXkSThz
KQ2YIrudDi7OHXcnuADYYRyWUCywuI691Ud4kBEq3RUvmf2t1MgrwvICbwP98bzvyh/MptwBAZCF
Dv2dw1irL7bmDzJJOZLd4F/fOQFVQ9H0/oBBpXhlGawdy8txJkPJaF7lCTNISg7GxRWjeJsw5Qhc
EPtCk3I7ZAedHhJLHokrCvgAg5h6CS4Pc/bAJGnxhv5V6XRUZ3v0sgkbgdSouGR0hYkmInHVb112
OOZ/Aqq+MyaSgMAcVlOU9X3up7Y5g/KfwTl0mhrp95L0t6O9jXbAY84Dxk2OjSBd+iqngJkrg4sN
65lyOCBd5lKklNo0mykoV38rpEbtE+zH2wafkYN0qReeRFQ3hepXWITX8ueLG6U9VA4Ac5M2g2Ou
Mu8rQSQgAYXwU8cRWtkQIKwwhwsjYeNNYVru5nPBKXaZOcZv/Ge3qs2nfUh0hC7hmR+pxijVFHco
oPZrnfSo5uKLYWyZlSnBXSxISQivs4b6FGW3a52mnbST5U0DfVGu9qkBWjWynxIMbr4leG1MH2UD
OJrwfuE25HJK6Uj0UNSkRl0fYpn6/aBWgNmHxhJrE62+CmeYeS/bEEj/uh0e9eDYD07WAyhDI9eF
Fb54YG+gbjfGbMHLE+ZLEyUmVppmweIpjjY4ZAz9uzspJZ3oQydwliXLJOQ2UJuoQfErnHYkWz9Q
E6XKxg/RdBCgGZQScl/arzSima+i5eA7n7zquPALyZCdpFaOkLLaigcy/uUbP1SBi+eK/Hol8FiF
6sbRHwWyUsBpn78UxctxZQRXFeFc1dTX9I3k83kpW/XWlMgZqDY4BdkPhDjASo3zzjMlqu6+4e7X
yrRwVr43mq0tv2FRESght5Nf13QvQOSocVIIZ8NMPzCsjA3GTgeFKcLUydQk8o3oQyw1uCTFFp2M
+fuZV85dhFSiUgtQmFmPJvNqA2zc99YudQYAIWqjfw0p7jbf25zaIgR0papXC7rtPTVBeSeXUISB
2IF3e5T8Bq7uZ/65gC0RVCoCjBIOade+hD7k7ZqxQV2DtIGgmaFAW2mc7cR5lalxPUcEYdIyzjGn
cIOxkcmMTYolAX4vKx/9KSNiRcaID6A8AagFhojyZqSkD8dPy+Uxv1qljjSFxXeohTZjMp8tlSxC
AE30mBPuxkB8gNpPdU3fap3ahjiLiIpjBKEWB2yfoqRgdChYIOR85hyKUWY69GlEFCSWxChiAaN8
plcFLgksniVwLJ7FPj0K5QXaHWoeljgkWE3vZgMA29vpk0N//h0EQV2E9EZMCLQm5Ftbs4TafGhb
phVyL0fXMfmygmDya3U5Gi4xMRfpGjk1kvrBs/lq2rUZd9Ep8fqQJk4ailE21MIDq6pqmellF0+T
ezI+cMukSqPoqb45D0iIIAiAbM4Cfx/PHVVgaXEAnGNCB0YZlnr/J+J9WIbAyvheYjSXmC0Y3gh4
6y3dCmJM2yJfIbeWxqXn1cbPTLF1Y/kfcdZMSNLuYyTtAtfBXS3y/J0qE+9o38xDWu39sUkdmTZ7
gDHaA3IAANqo1dpMSHmp/0fhI7aUCXrd+3x+P7QjV90qcRGyokO91dQOr6mrZKdXppafDhd6JWR9
W9ONEfxr1gpTi+y9miE7PvmgwEfdfN7gQKXn9MUg2yN6RGpwIs/AlzivnC5oQ2N79xdOu7RZFAeh
QM78oGNoSezrZh/rut4V0Gyu/3Fmz1rJ3JZIYq0lv1xMfpDzHySWsAi/Ap1zdoBoMBEV4wJFVYL2
Ux1GapKvysJ/an08ThNnkNqC0Ykxcs3/8md2rGngqTUsHCSkWA+tEIJjfKDKEor9PkThQ13pVJqR
624fgYb1j3LYG87s+2FT9bN2WQxawyUH2J9gfEb8QH9gm6BZh8kjVS735VlnTD8+l38D8BmHanXJ
It8PZbO21PUlbBfMWu436FPaGo5YqSNCZSy79VqjqTIlJGAQ5syvmUgoIjHXU8/tAj4iNHKkDrJ3
L/D7XoMwrgT89FUXgyisiVDjRsQ5LrmA/ECP2zQ6q27nMLrqFjwUFEtQD1m3bmaX73BwwVziwkdt
dscrbSlFUZPVmO/LQ6y7eMjLTLILqHWdbxPtIsYpLRxbY9ZO1jGkV0VueMkEia2b55JWJz+E+J58
unwlQfh8MMTOR1qFs0LBfDQXpzEOeosaNf0s2UsCmVhOzTPpDUqyEE7bpINvMnaVdl17PLh0+o3o
zRFa/mfP2T2BCYAIqn8R2qDeeJsOb4S5+sJRSB9gc+1xKH6PMMLdifPFloQdLNNOu3cBecWoa5vq
erEpfhbff2lAENtqf0g9wo7Hz6oYZ9Q0FUyYlNOqsAvhX2HSlEz2JIhcw4ISqWjPJrcWmBr15Jeg
RMGkWGPHW4rlQJ6Qxysvm4ype3EzV6rmBKEA5V5lkXmgMIZT3esztlHWz8aYLTGaZqI/GvU7jOiz
8NRYwZ4jpYs40p3UiVJc2w+gF7h6V1KKGWqqMLH0zkpilGgaPyu798lwbupaBBTMrK4O1T+bRDgZ
Z0VmXNSxEmbmU/A9gmI1aMGp3mNxtiagDGMZ3lNXLSiXIPRVOE+qD46JLOJx8P7NSYtF7JSDIdKA
zlG2r3A5h7etqZDX3Zac1mySDOxstVXUWIbQxkyB7gb3d3MDl3KLK+Z26hl9GTVuVoUPr7Q9m79a
DORA0qNA4/BiDMvl7j4X0AyzeL/IE/ld1Nk5a0XBKvDheWnQ0GXkg12WNg7S854C6kT1agoVqGya
ZroebO4VcEd91U8jL0WTAIKPFcMSWxGoVvAoXp5GV3qNoELBZ4+uFkb/92FjWOJRpxwRcpEKiGWn
5q7QiOqhQVzvB+A9jTDm1MAgWOfJXvOseq0gQeWXgXA32phVUt6JumITIzeDvk2NceYHf4K7iU65
p6e5j38MZd0Vx4qEcjZBrV2ryQM4+ZIL6/4BFQHmkjKq7lYiJlOBe1pkVQMK5iTAgt4ThP0mMRrS
EbXMUSse9QGWB79F/MclyG84qYa6YF/jLk4mvrVrbQhckIoyGm5UFjSHogRvyA5JfYs5/F55N+tX
xuk6qZYj78JYUOl1p7cbWtRrKTOxfHFTmdwAA1WqG4Zr1Xged5K33qjvjtvyAG22oCCNPIDTNMTp
XkwaNIM07oPx0QUYMjwHbgMncAGF//6WZ83zDnbGeXSwuVjQwv24giGC6WfSA9BpAd9Fmo8uWnOr
QkcoWw9AhJFSAOhvh4bQwqR7SfVmHIFzqYCUJ1PGu1pUMrS2KOxhJNNev1V1kwBCndmLCxgMG+Xg
rYmM2/GBh717iXWj3Nd37AvcTXCS3SeaEOagoqBsf6PO7W5iAJjxg0xxy8BdFEvLm5raEBLEZR6m
aP7MEg43xqpaPUki0k6RN1rq2bCFfDDcluuP49Wlhc+cG+g/aJayV6JamYHqnSxivQY29A6zJFqE
a35rVD+EldDGziHLFVwEGJ7/Bez1EeSZjhou39gOJMr4ShUUCD/79pTsmW/MZRnEyipUpAjZLUQr
f08LlgB9JCDw9mO/cQLWO8tl0KeEu7ME4vJLCoGN3wAAKFqQFUwhegzFk+38yYrrU/P//ZtDOiHP
jT7kSzWRd2hstkLx/hVAKEWOaF5C4cdnyvses7RLJBPskXA5aNxQaZ6p2htfbiehKqqzqzSsAIAX
zIHYz5aO8dTXAxcy3f8y3o7qBkDEGKpDRY3sXrkPw6PvSdphX8HXoupG+pOzhiY/1gEIB3wr6/XL
rBoES2kTiAtOnfd9IBmXyQFNe/DwNAeoisPaRNd9p6REVXFYecVZJRVbC8cF9df51CO5jD1PurOa
Nv1VWoJW1GPHmtmL2X4Wf8x7Kx9KCcGIoIxiwsWkSi85k7CGsDjK/NnuFbRcDukOi9A/ldTdqTxC
r6UhEUo0hiAnrBbqpJtEnHNXiDW6mF7r/8X2Sni2jNedA1dUCYImBY6fqJX28jxsRJdN2B7FCzZl
uOYfzlHd/bMGc8FvyrOjqWBsPrxSaod5V71yu5821Dc6omK1H7anUlt5OJ36WdxXm2bDe7a73cY5
a2aq7nAXus1KC/VTXgXeUTzSTXh/RKHyMVjwLqwvQTv0FhBs1Le+QshAdjOSQs/ofranXzZ4Sg7b
YoooftKJb9W5PPnAGtE8O8tFq7K5ORLiG0oqPDf8uB2jlYlaoOsgWinnL1qCEPSa8GmWzWclkxpm
u8rsJTkznH/2938F02Ayuo9vFA2lmoggYMDrOix7F23Crd6ck4w5SphyNBEdpR4YjhkgsZfB7zGa
ePLb7pzNBvLDAPk8SHy7y8FrpZ/YlSF3aD1Q31ViqYEt4HTrj/DxHiy3Qfej0fxjSS3HYihB+rKS
affN6CSt4vLaQpnB5nslStUkUXWjCaYBoU/YQOTHqQuRfZr0Ix4tETepZjYZNpMXy5Te5pi928qZ
Wy+M1NNTbYtfzgR4BzEoTKQ/MnUmvNt6OVfJ0xok0sE4DnFqE8h2SoLNcxPwpsTu44o/r1k8aSSD
Xv6iezCXIVxoEiJmz2+S1pBnBHOVoIFXSxAWr89n2O12L1pm/IlvALEkqa9U+bQv1gqFlRD97Euy
kN0+wi5xhDVelJEOvRgqx13MbVnc6N5N3m3jezrJk26TCQTp0lHtwT6gW1Bq31FLKD/LQ4Py8Del
nvagfylGI9gOilT9s+Rlgr58iQk8F/iUKwz9ang+mau7GaeR58GbWaG0PsdptaZsYQliSbGiEOWx
IW0b6I7XWdZDTFOgYAGE1H42DiYJBWTb5sumr8qp2edwX4NHng29KkvYJwztUNfUMUfUgbZX3aDL
HLW81cvFy62MAXYnghzJVtaSpGdFDKfFuKZ9EKPiTeRjiOcmNAI2ENwULeMjdmT34aLr2sd8XaVS
kj5F6CUA0AAtbJaoAJR5D/9I9ZgR4a34gg+T0ikqcvkGhShd7XamB0SAuRxBBujk21BLCFibxrCG
OExtndVSvU0Brt4Vo775dJwu7zTwkASVACGVh2XTpMXoCW8Va2tk5cd7BbFIAuJclAAi/7cygZKo
K/0mmfQpXwzKmGLs8X8XdEWRk9eY0FTcd/WKbgFbgpSJduPK6oMFzVf9ig7BTAavjDzZXvkOqYer
l4TYY5WlNhxlguKu0nQ28zHUwoepeYhl+axj9ckMExLsAHFwMxTJfBVbVLK7B/YYRfu3Ko/4Zl57
DNoChNYL0w0UKQaMm40WOmFh5vvbaObczP1+ZZlAE1Xm7hLlv6jT/yt3w4/hU4JEbJqo8iWaJ9KH
uRek8DQElR9sUurGlGjUzElthE8/ewqh7piLFgCKFY8M8Shc1YrI/jCa6kGk0W39BtXmgcO0MpnN
ApGo0CSeIOJkTsWX/ls2uQov9CpB/R9jy9OJKrtaatcfzQgnNvKGRvsb5FW1MkHu29EAtlYZbPod
z14e2VPsyTmvvM2vBJzf8Jan1q9C5/P/4PJFVfInelHtUi9KrTkE4YVuiNLcm+Ex+EGyclS3K/sg
GyTfEKDPDl/rpwQCmSPx+GDSTw1vTZd4lkCiA4IoensA4Zbt+yodjJp1Jy/3TdHnKY03Vd9OWG9w
N53VnMl1XS2nXWgKIa3Jj3MXkM1vB49yBm/NqfRIK7aVX9WKsxg39TESqx2MZkcOTd66EHvPkTeK
6vDGYCw2szs+AN8vMRtFQDu8KJTjR6GhOEQk4BleyF7nx8v/J+ORBMcDhC0HzqaQb7ZQsS1B5/BA
LvX93Rt5qtbtzN3NNVLfWm1SJNfWbsFXYdBhl0fEKUJxiGHKRpCZqe//I/HJqsPB3+6C2m2furW5
Z5xuBRgAMR24tOHk8gwDDe7XnUo3K4tZ3csudgvq3SHcy7gUUw/ttQjzmylr372DnPjUvzgVpcGU
z3+l8LzCP9cvmxh3sCOTQeE1+j6Ub8hhC4FdwxgyAJ4mkGMMBMeUWdP1OUsDKrZad5hmo2wQOHjY
rF3hOTOqm0504KvVFGZzvToAozgX2s47fhR/p6xht1GrgRddMkZo4CJVuKrlhhh8CoAvZrQ2W0uT
8Rcm3ImQhL+Hl/Hi4JDF75X9c+VkNP3CGSz8XYs7alY/nrssyl2KsIij3X324Jl6I3tACnZ6pefB
LJHIcelHGPo0Xjq0veEIM4pz8wJPTikh9FN2X5KlaDSKxw+qNGs5545GTrqbrq2cgzFtJpHPOpPW
dVdS+WIA5RYHosGz3Cbt6rCVWrLSkK5MGj1RdIAYDpjCqSk3spf7txKpum7M21xkZDnZ03cHyZQJ
vnd6Rr0moZfAO885yPyYkloEFOzSk3pP8swyMcGxQsJILB8goydb9iG0kUmZcmRee4tio4O6gx0R
rSv3ug3hy/jraoRonvEE0ARtmZ2GqMWbqTuNM+FavbVy0oLVBhF7J2BOq2415rCManHnDCv9Daqg
GVg4jovSbrvIlKomxsFQJ7No2hfyri/rshIvM14gcLWLkqANKADiyCRKj/vAApYjvossQGlPYt0Z
WkZ7oqMShqFVMiyThcEy6wn9v/hHgEFdE602+eBQzHlz9lKlzdkdA1FZAK5d8jwd113168Qy89G3
TNVM05GXLBINgXQYzsqrzIjQZN/OpobPShTVOpQQZyZVSX/AEhiuZga2K1ma6KO2qdC+d6JvI7Sp
G2bpSQdvTacNy6VClp3o0Y+P9GCe7yiIbY7ViqTlPNChprDUs5n7ZC6VYBB25R8wRjsZ5cdjJcU0
kcLsTtQLxN1U9cSHy6eG0WmBwZFCZqXwZpCrLT6cLX45DdWN0l7lKfZlt2dZuQUd52D8lp9c3/IZ
OI5+Rd6vkmsix5DhpJDPQq1cgi2rxYlbL/OscGDGsJOf1ZbV1GHwJwt7UKFMtRW++vCkTJgxmpjx
y1ZDQipSueweqfEH1kz8sqGa3C6PrAuX1zedsnqESOrUUG9xN+dMS/wWxmK9hNqTCK58mkLr+9dN
WPF4Dl1Y1AOTlLM6X+5lsP2m03T81Q8oJCMepYi0GYwbb2va8razsp1jgvjxz2cppKM59W75vTOS
w4OobpzrUoPaRLNLKgT0b54WCXHauFcjDvKCvIFQCBKYyrKUj9sNdl5mYhx64hSOi4Qf9WxsCGKg
CNpAkyj8wnVSMJ4v8PJV/1IKzijGhLxNnZVe0cAl/kzbHAHBvP9qZlmvl9vWV7Z1MDLg5yVvLMlB
V6rQRXxcB0buezGRks3zujoi06v3NxogTq8NXi3xL1RAkZLKEZEPTbB6V6HvSXCCTHKVUJ4GBvGS
M2syMmfiaJ+LGPQ3wNey4hZ8oALppcL9ZE9666ni9z3dhEYX2C3NBLW9VS1MDFYWB1x6xe1mLqZL
u3RRdzNK9qztonfqp6gL/PQK32LxyltQfvNClWh33HGte1WXA0v0Y+Ry1CBmP//oqs5Nvn13McSW
SpW7peOUd+Gk4vEojaNMDFNd6mSocJwbLBQW4QyrJj7Q1IbaUzEmG56+TW94f5aFLB/ukfZHwqE8
L/IKrXLB/uywGNjp8gGMyQ6YR5Jco8LHE4L1PAjNELP3ZD+1a3zukTVj8S6o0kqOhKyrox8qHLcB
UdJ4n+6Ryd1csf8qebWjRqRXMrLYBJebFjmQZiSvdu/B1c6KHWDaNcHh8l6r3viwhLNPpS/vrOC5
0ozjojZfaKeGbLxvJp+8ih5XMTZCsU15REVUbZb43nArE7Cvt3jqGhbVutOHBKZxtpPmOEojI494
4JMgBCTLUcJEnhhL61tA4lmoI3t4t1Bt7NoO/fE2FjgCI5J2ki0IiRqiaUWNqgxzw1sZ7oS0uSS0
z0NRDexLYtJ6HTADjLzUFyGmFWBsRJBy3uo1Ai2atcX96Tj1yqOhPB/W+Yk96+DbyCaKsDYox33e
oDL0GU/uqXx/hTi19TEXIHsiedDKKNWxBE+SBrDKWKdT26XCxQ3dTRMlbcZqFE8RjVp8R+91UxnE
RSfqZkp6Cft7f+4Kb13wEXRt/7Mau4S8hlA9HJKMbUx8p0R+LISBMYx7K6P1vnNNppLerU5U2lbn
BIxgVDQX0BigqzbTob2k/wMFp1kLVeEKYCymsHJgUPrHSzBjdUvNpu2BJut7Cjss90PCXO+KUe5I
h5Giz7wFLv/FGNKbFvEnVl9dTqK2a2p3HLT4MRHSDoiPq0G3GVS2+g3pvZlYScy5QwAwEjsmOddy
CNQ6g6x0zJABRKYQJfnj7u9ttx06bsvYwiC/SU02QVbW3m6HAcJHGqcW5F+azpglyjCBlarEnvgI
rDKyyXIrBBAdD2KO7dZet178vkEH4IiyG3VEvVm614E7r8jMHnHNwsSjBG/58qAQV1J9XDI6X4Fs
mv88Cgc6jVbA1eWYH3Px838wDCT3ilQnyuDPY6/C8+V/GrpX8fzdjFhLpZtJe7kwtJ8ZSuFIiFqk
ERsopUBu4aNpIMl0fj1TVSQlxlgLExlTbSmpQJCowGo1pytf9lG+ALveh3KDlStLcjpujITZm1uW
War2Sh4PXkzSBK6WtgRE//hCnTx7zZE3rzjg/jncZWVOum2F9ARXuDnMlAb1HSzWOKfl9SHQ+62x
oNwAAESTbaU01mt0p4+arnkX4BlKqpEIaMXb679rS7zhwAqCdnsmp+k4QO9mgumMZlp8WV3YBOm9
wl93MqmaF3w0jorhyRIF7/WM6CR2KUotvyIUM2SPX214umG8fpSsYgbIea+WZyaKoFYT3ZtJ7QRJ
aQ75x3aTYQSJqpPH5LhHd5aY1uB792NGKMOfRJWfqDdUr/ERQXpXjLCwlznBzAPUh2ko/V7WV1ba
wcOXiMziKS14uFOUD1Icx7Aqb1CDDkzSFF7EAeJ4qiQoUlVEN3xYAXUFnlvdr7OFMwLiICk8bcGF
sTBojwmK01riA3T+B4J8koocTat7saHeeuYbqRQu6MLGWpxCrAujgIUtijn5GuJVmmGamkhbgids
nTXRz3rFykKx/d00INTRrHkqp9vIoUqu1JuiT9VMBFPn0XsekG+XkzuoGwEgz/qnemqa3A5gUP0A
1raljm4bU7EgvgZn9BZNDV2FyjHv1WyUnl+twV0BU22nuKtotyvNzaimbdj8LtNsOtyDb3wLmJat
EBaU1Z7JYPY8AuwkaLfk05ibI/MojsQem1PNS4VAM+KdItMR0oDrJPd/QAAIglgmJmMQB/lpWQyc
72EKRa2mSAbIhhoSevDL1qBRAPzCooMrgjXRU9nte86ZaOzNj6godQI8YQDAf3fZ3IhWdozZxh3h
n+HvMFD0arfFb/HSU5AW4BU8/MEeQA3lk1VZsiBQgOoDaz6PsJT1DLOUH5vKLakOokDJsx9GfLXr
DKjO61T5BbAgo8WCfQ4JyKtIuFkF6T89Lh91k55wv6p6uQ53f5PrrIGiQP/JXDnbYHNDjqEu2P5o
FbwvfYXA21E2OzZJ/65UeAjB4La0YifI34s5g3VtVfln9TLQ8FjVI5lZms6AbqfzwrabhJzPKIUw
DDcLCnvG++dsEy+e3D6bVpvO83eaJ2TavFvli62aueNxbzZALI/tZNbsrvOtT5KPIv+GPvTD0qSO
FkbV2EHavRH6vPbh81VZ2O9Coi5LqZbkgl3KHqTrbBA09hkxWNjwzCl1mqa3e/XMM/JSLAG0ZKIF
vOuDABh+R4IE8PQwWi70g8ULjCLW6/QZqiNyzxYCVSIBXuzJKW7niSZexrs+gar51pfpBgPEVZ4K
C16jXUUhVNISn9pVyqo6IQ/6hAQnaLoacGzorf4iG1OFw/e+WusEjEiYo8dwmoHfyyzJ8nzT+5pU
uvFEkD1DKY6sIZgzZtFp8CoZTRbaYzAbX4kuSHkgL7aJb29nM5xAuF/y+xT266/u4S/wyCAtY8S1
7s2pw6o0X3kuQRenQb9Bgx8MDL0QbxEI/LfUT+yZA2iDYws0gV1tpBL97Sw6lIU3/akiAc1vVFbt
KihCspgO2SMQSDrgWrN+7t5BBF0MWG2KHn7LCvj6pFcFHXrM08UpxpajIGV4rZ9H69rXgWKRL4Ad
vFtTCefMpa+IJz855M9rb1Dw8X1ciCDM7nj7pQnwYlusRz55zrdFtIyuLE3XwnXROPlDksP8Xwwr
cZu8KPNjX34OVB4/i3SZscPFXO4ZzbqdEiy0pnk7s6FDkcQ3RGLZP4R/KvMKOIqfEU9N9x66AFO8
7KGG4zmvreX9zqYr2bRMDYeIZ82QfPaJ5IaGnQEiVJqQ4bR89MzhiOGjLfCLLHlDq6EYAnGh51QQ
H0I4gy/oNie6qJet7sLpKgkCwnlAsUJxXlcVjb4YLDLxwDAF26oocpSywpxWP3KPOfHpay8IhrOL
NiCvWaLY6jpe6IzmjyHODbqhvgA7vBCb5CgsKp+Jufby4XMwx+yWGnobJgEiCqJeH560OAqTU7f5
n9J92b/Py1IeFRls4fLm6v1O53ESOp9/70xZV80CkieyWsPxVmTwkUEDyaVnseZBCfC13oKJoKM8
seFvj5v5D7tsbc66TEI+n6v2hvfv8E1zpqQpTGl1pWHKNhEvls0Cxtr1FNcBsJJf/iSYp6RzAVgp
Nhh2YwvZtixCO/J+leSpqq8+9xdaiL9sj4TB6OfAMeGdA35+WMoUqRxpguxaouKMfDuAhYG+plvo
lZsiC1dGaB7PhrGeeY2skV0sBVK5z+/s7f3jMjFTGQdPy5OX/VMalZyIuFYgZ0fq7rZc2/mF2WpC
ip94U/VqVo1OPayOiK0OyVNpMyY+Qs6NXdN36CJ5JXwyYVnCno4JhMfHLj/vgam1Ijovp34/bORy
6fAd0sgQN/01WbK6BGefMbZNnI6RwWEtFmhMKZ7PxauCvWMNx/L0naw4tJgmCgrzAtHMnCOYR4ty
5tyFuCtF36vw50jjhbgPmgQYPqAnURtBu5AVWmG2RMSvKkNG4QQaY3lx3eWjwt8152BYOzdM6GTp
HijFz9AMa7YTlz3DI+1Na3XLHWwCDDDcdpuwO7ECGWLWMyezeBMu2vwcWgdlkP94L6DNpjA5j+gE
TeV8qk0e1IJrMsqP3AIwIloepRNOy+oJXPTF4Va8+YqkIr8G2rFYA/ilT1re3oiMwW7F4jOlMjku
6lgp5S0TdWt9imF7Xs9vdvvBAMDP0AX1l2epAKQckYokupl6QRr5LnUXc+IxVZeiCeVII/YI3ThZ
9JqUhEjIUkN6rw52IiVCx1qnLRJhhUgCPlaFKBiCtjotHDtIqGP4bZ752tFh0EAEdXKA7ihi3wa8
/L0UzfDZeTFYilSrUe9k1BXOKrE2YDRNpAWTqh4xT6GV5uBF1GIzZFv5539vjMbcgl7LGDp8JkNE
5AFTEVWBvDCfNv6rjAlzxsGT/gEp+axj4WZdhKNHU/Hg+jz8D+xQnVZJeSdeR/UwwXzlGopp5CiP
1FThRqzhsMuw6OiQUCVa4me7jRIXqgafpZiVmX7Skv4eDGCxaB+15J5ydWXpQeHxdgB5rR+fhCPj
6RQjm1+lU3hYziDx3HX4aA/ESjHOxeOMpbkSihMT4YTRf0izfBOEWCIN4awVHHsQZXa7GisiCPc/
/CW8oqtKcRmSqxAZ8UIFSUnFnAChS7RG2wp9j7lpLqPiFphqwXBUAiymixLCcizw+SYRqev9KXUs
dVRZvlXUI6deKebyYMgcWMEQ30ecRFnVRge/Zuq5cuyroQVi4MIUMnTjMSt9/6DdHSc2gaqjmnlS
vxLabv0OFuBcjBlMsjHlSDcEWpY3Jk5asw/BbDdNXXvifuNK9Jo2/7qqMSnnByczROv+1m66dxWH
rnbLgb7Q1Ip1jKYQgtu73VeLQMm74W0I3x+VquQFNXXUQRFmlf6PkYtw9GSIIOwBLmFKt5hEt0Pc
ZmRvvgVLTeBeqz6zRQmLCfNnWOtc6I3KxSCS0k+QuVmyRNN2MN0uwYHQOmLvXRJke75nGKiwOIpd
S2lpzi5ejZUtXGwyx2wV83FzqzDDv1PgWlZXRWqUwhwGvDwSiqfpZlVMYyuuuvAtUtthJNIgoNL5
ZDV26BwOVxDjUBEnDTsMavdediX9v4G58ylL0YIKfAtjjWVj6PJAPk/ojWZsX6yqZ6iCLXCGFrcg
WNAbU7XyNZNsWWeh9dVVUZdHcZTPvkDd83nuJEjdLIB+IuHdflvA9KlJLfzfRctwIzwqX4jL/7+a
MwB9XjzgtVQksxWLUCq6PHdBv358y7H7PWJlPsOVSiniiE1B3m8DVT+OU5mBpz20JbUc7jSFE+dl
bsSyqv29IozqC/ygxF/YFV4ZH4VXP9R6cSFT7JTe2hGAjrfeRZzPa3yxUG8zysleUDSlEFDOYaNT
wmdqe9NJaVPAEvZKUUevxyIm/XSRP6gQq5pEkfpViyS1ANF+mJF7MN3or7sbJALBD3COKp6RCgAc
guNi/2nm3IT77JfjmVunSbOJhp+K4y2v+pjRHyiIsSPKmmbc8wQcxAj4WtVi734MS1dDKuwT8Z4Z
97GuCpZ23IvVmsdtdfRjya5AX9RtpDF+7CC/l9lsV3r4k84alv3h4WF1/htu+qIGrhXPTIqqX9n4
+ZqURJtrzT1M5me2AL9UF1R1MCgXVhmmkWPdz+ATb1sBKoGV04lIWGnNt3hx7ZGqiF0kpa3TvGpI
Lo5jkdgX1FFwWs9+NIoORm1fuj2VvfGiDyFZsHdsjC0SXqUMf+F3YMoi7jn/BsYN/H4Fc48rdeSc
I7ictAm/jU+2nVcwCwWi/JdXV1RVcVLjy44kQX/962ytY9iVBq/9wN6zVp/B2dtGj3cIWEr66TF3
YXB68/NRaYwx05rCxMkxwkQhmzfW7NXtgZwgBb7+QHHUcHJ5N/HI0WcQmNpPOk960gr9DeKZ+/+r
e2EVyTSwhOY+HUMwVnZxm48LPWzmGYmuAAaldX065ccn/sj5yAr4Gj6e4txWv7IfMASRNxjFmpPr
PxhzXiXnTXRyH1hgpFVcO78lPCGFsNUu7udE31cBHNBMs88y/bgecee3X8oB7vvty4yKcG0fy++c
ZZDYa2hHxdTi+oE8MJIIgVSxJReIE1yypVkMV1QYBqBVXNfHijd6CNk425Nu9e/BIecDDwq1vkwr
8H4kgUSOWrzl52WOKKCXxt93UI+IiDCyx4cclt+z6ERpAFL/RC0t7CWYrTXCSzLiM/6OTfFsjncO
fyulqd9IOZZv/j3V/UeEAY7w5jtaEH6oFjWPpmNvnB8bJgvM2nEDtmis9YzYyz6hNNBYj5XWzgeU
l1HnEjexBxEYvcEcb/AYgCyzSEqvUxgX8+hZ0Si9f7aHl5AQnQigah9BEEe/Xps5TGAcfAlwmLcI
3Wn+KTL4rolynDP7kk++mkEK4WKMgSEE743bP3sxwaZJiz/lWzrKBUosxZ3yQMjdq4K6rEYdWupo
ncACvt8t7zveQhdogUWf+V7oWp0ydvtKuPC5GSUzfLfSgdNbcO1LV/nPUuzt/t4ASnlJ8H57xKQ4
3Y6h15OighttMPXtac9zMCb1wQEDUjheHp637oa73DUvhc+YnTdxP4PxPhifWrskwYIjcoPg9+Od
JD+X1q4k+2zsfE55nMaJDDeL1AufHkNFsoDXnTKrGEqziyhdVsOroGCwgInbR0vTXBV/oUWdgRuW
e6sUZN/Zz5RUCkx0RrhUNSoqHwf1FNKgi7zCsVFEimU1o+THSopd3OEYXxTvxzp+hUuNtx/VXwOz
UziYyto+Pn8ue3LnwEGByRaTse2Posk5aPaXopL1nbAT5ru6L3Nv/7t3olcZLWmlL52veygvqCdm
DQpEs72OCg3OyCn6XeFTqMD6s0eBav/SaOdcm1IOccunBEK+WGxmyZDJKwLq4PEOrz0IAKZlz5i2
m1uMvJXZzezG3FffIQLXVnLJuyaO1RFFCKV1dO/piMb8NgZwh1rWXFE2LefMUINm2bgTx7ZO5DAw
0Z6/UTLbbwyLb49r3XPMANXcrjU5QKs2KzCKsFymXbEnM9imFx8ggKV0an9ntWnACo/dQKaixLxa
hABlFwxbcL+7CnhmZjdcSKzqeEzzS3rYEboR1E5o/cmw3hF7vUKOGjmqu1JSMHSa0KNdrE/FJkdi
aCaVWHve77B2sYAYOvUqRgJb2ApHWm136ncJ3z5uDFY1+aLLGNm0OgwZkjDp/XG/yYzFnwa2dIS7
/j2LcAoH8SK6O5J5fHg3xHxG3cBuxcxy17UcrQdF9j87GwxQWk4M0i1V2csKZef7FWc2pR/akXeZ
7YjrbalSqSrULfLMjI6sLzWp0H571s1hpVYAfaX0hY1t3ZCbSI7LEYfKCJnWkWk1ss1KeYzhxraZ
ZxnwrJgcC5vZ1U7G6gq7taQePJTe5W6u9X2VQBRIaOZLsNzqX1t/J28sfb8SnnLsaVcP/wQBW4Lw
OG2LT06xtlgksHQF9gI/N5AQClENQt5kVG9/egWoecYtsdGrEeEKPmkibVi/kAELvFK5T0cWPWNt
uVl6VMFmjODhMZSF6XlFWtXPK3iegVTx9kPgwSxQIW7h19J5yuULKHkxHJrsiUiCOsJLxCnjWQna
JoCp6nutaNnu1138sYSe1AUyPDV7JN++ErJu81IYsdp8bBrkCdOBSP7nW7bEd1iQo3/qar611XVX
K8Pc52h/eqE7Wk6dgdhKhGZT06RafXfvh3qYChoGiWlacXVGsJvM86Q9QI5lhc46N8pA7m6wB2CC
1LZ5u41DIgBF/HCqIEdaWvyFQqfUn3STUwKndfgh278KncD6RWWSVIn6hXSXWbG2t2kL3/xpGYzd
X280qOgG4VH6dtTPq38zhiOvZ7JLRH3Fu2GnF2/WGnxFBeRN4GLQ7y1oc2MsZUb2U4uw3zjt/+Gi
TZCq3YtjCwdSGDLymQuyPqFzWQpdPw1p9PMKdcn3intYtYJ7fC9+bpdQx7vGPebHSgJzdggBzFGp
Oym4tM1HbGgeuk/RQSg33xN+4SiHgJKaaWXlhD0BHw4x1aUHkkKmJ+R5N24uUfMFQqt0GFVqn2+Q
L4xeyspgW4XtwbIHt685I+U/0PRJNobP5pN5bYLUsri1KQu4W3BBrLKQHXN23wHbcH6BhawSvvyR
JhSR32gwyL94L/abLSE49POTIaKluMEmr8TZKORoFp5MS+/PKcF31rDhvi5kh/c4rTt08rvIggZu
7Yta32T9hMuML2oLSeWsRY6wUc2mMFrq9f9IQXk22Ac+bOyw/ac3a7SMGhy8wMAOAfgo1o2dKWHT
fFvg73S3jciaSmpU7tf7FiDjeYf88Mp87gCrQZK7+jFybLR1NBvhcazgQIr+HhcgCbZMkeGnvp12
lFccsJI0FeDaLquw+H8bWH54FC75/qOqhDloXmP841j/Q/2fotQaTJQY2+XS7JLdrGVajZo0HDiZ
F6vc71IgEk93OguGWiNbQpOeaOIvdRyIxmIPL1OONv/qT3H0zV27Fl2GKNG+bF6WV7nSjKCV7fV7
cyntC9YqwNazpSeC6UAH8HE/WcR8IY8vx6Q8BdvHavqaZYC2SPd4DibWiJ6O8ilpAbXW23zCAcai
PIKu27OWTEy0jESSHDqoi4PiuxwvDAvVtrzes3WEol+zLJ91rYpzUL8ti+l1KMIx71RU78POqFJZ
9OpgIT86fP8n91qOx38JEEnuBb/+p4gU6XRcDLFeP2h4Zo51g7s796ZnHdV+uKhEbev5cH3dKq4O
VkcwtAa6NGFEju7SWd9oHbQXBooQC7oteh03TUv0OgqSNGpuGIU10rXoLCuJtxpK5v3Jb6FRn1Fw
Ae90Q5oOOrN7F5jTNOrpE6odniMo3tak8/4CTqawEJC1LhuKB8rvNuF8CwjdjzVyYpjjTK3BL1yQ
OxOjdOyQOwdAmuYC1F1EyO2n4+KDvjmlJtKYf6Brp1ZLSPSj1MkDxPwZIim6NZBA5odEItOqVG6M
AS3rxGKrBLXiknbjGYqRr3Zbg2lIXr9ZjuSHk1Cl8pW8eiR0wb8CphbVuBDCtNxiNGuH664NPNjB
7uM0iv5e5Awu/f/mMGjoxTWMMFyUyT4KyAKawxNzvk8wfYj3VpFkad89Xf+0riD8b5s2s81P5oRw
7QHdWyp+z1hzR8dmrfxd0DUIFTt3x2+a7IPwal5uUDJqxJDscuCGiAikCjeMt3uYoQT+KkUABxy/
LpWFW8S1V8SM+DnB0iA+5DBcrWkPKRxrZiG9ratrul12Ya2gFt+uA6/dwYQsZ/UoGQ9jEyUcbCvs
x+R9UEeH0M875LpP+JOIGNWwDwkL/O0Pmn1wWMaBbxxcGRPCbjpZ6mbB27iyrhKChy9hC1pgXYXQ
UVHhMHI84FnSv85Z8To9r+F4sSlZCvMn9JPadsReCeYcDOR4KVx6D2KdQvbsokijy9urp+DWErDh
ghygYMf9Q/IzLSDt76WezzpLDZxGjjBtt1pdvR172RVxTsqhc0Sbs1j60X6wIVOO0HM1VvJMo0hE
1ibAkffnQqDpvUo7U4JFrgy3k88JtGF3/qOqjpS/iYYjPFIeOCW+ywdad1FRVUHsUCoicm0QUZeB
6/t/HNEB5C/0mA2c88KEpVXG8ERB1dyvtUIiWJ9F7UB1HBG6VjZxMuEORZAlGzvWrHvqKa8hC09U
9fuyUGiGb/c4Q3G4ZiMusSXcShcy9x2gHxCswgCDr76TZK1a7UqeyJUvzL3NhiPJGoweAD/ATuFs
slwpXVfNzTcBFaUjEUPMTAYwSQ8/TuBh/VNrJWBiaqN1mmDUKuVOY9mPgsoGXnvXNnlfmEkJYvDX
nD1hpSXWl3v9cIGNAuK+yd9pjYhRC1D5L94e3n4g8/4UqHfCJMLgj6LQhQdt4Yopj79Ked3rdX4O
hBCaEW8iHejNO9CIf0h/txNqgT/kbXJ1XBp8fBgLsWGLZwWdclg1hLxWy/69e+NCGOEWFsIQFU/l
XJ2b4jp5mpyqi8O05L2OETnEbg+T5yrNs9mswViXfq0j+kpswzjnb18U9hVD4MdYBSN3KEdXh+Sp
NODBbxrbJZJwU/bYsG20vxk1/1iQKNJws288u+eUe1GnxKtYyf32rngu38FvcYQk1lw+URsjIdl1
fGbXEr91V0gzzdO0RribYA2Kl3cXco0PPxMDD42E0MZIZArhtgSlex+6SGpzzK0Y9vG4NbuyyEG0
hQvXN0YP7jGhE/fuWzo4L0yET4mGovEExZWT9//8Snq3Y8VQTdrCUb5xYPbFQ7ttR0Umg3L12pOl
vWgSB+9EH/uR2JLgNRhBK8Tw+kiJLtbECnq5m5Scf3FeTFBECUPKjMaCW/Ujc6cdmJGj2hyr8hB9
5uOwu0/8juNfPecEhDNpr3DvQ0xO46iS9M+gCuvCtqfaW2kF64HLDBf8zNucpoD6lEgAl8MhqZPr
BVyjOLjWkndwhzz5bJrkz9CbdvO6ZqZGUHqhjlpkKlgaTgf8JTmsdL1txlJmfNq45lW+PO6CGbvP
tb1eFGkAVMcWRphVoIlX4kaJGcv5GKP2vPUQzM7aFH4s52FQb91N5MShGmjMXgdzEin7GnrtDgqF
Tk0i4DjVf4ngg+Torp6EAry5NU8Mfi4LAgyeLPoqfPhHKpBpgUuz7aIS2SCwcV47wnqSdiy/L2Qu
aBOa1z2hlYbaBeXQ/1QsH+OiukL+d3TFmZGe1ALFiih/t1vZk8TTaFOkr/LzGoFsUbKRHt899iOT
B1dm7uE+82v1YmsDviyPp50zbWIrxrcpBaFBwOq2+8tKEkfvbEIYhJ9QJpslnFYkmAu2GmJF/JVr
O6BR22aU474rMXf53sBOiCw7F6lHaK1Ib6SZ4osoJmPmK+6vEOLrympp1YSPLHOkkVZU9+oUvBi5
CH1Sb7+b4SEw88QrB798jlOZWMFGjPRuNYOHr2vNxNsA1Buv5o5mNk0of++hshR+vcei+0wLEL/S
owNdikhGe3917eDTj7o+N/Ll/mDzYFyhNjmgEghdB2/skoVnUUjegKbOqkAeNY2C1gPuiVEEAKdx
Ql1r/G02tRHVyfGO+qqmlFSG6cJs0XsKlUNSJ8XyU0MKFU/QESlQ3ffkhitygcgYXa1qrMwpwn+d
xvzrc77PoeTE2U88j5OSgCFSjwoPg6ZRH1aOWfTUpDI75NdXYyH4y6bVMMCqsCzy8fYkBcC3fN/h
8YzmwP/xvqOcywjqZFpr6hNW9O/8lH+zuOWLOGBEZZqkUURi7MapDEOASxjhXTO1SlI16epUEoJz
m6Ouidt7MLuiDZmwB0LYNv2Z8BVmb1En6YbjntxVrnOIWRcY1r24n9ox9CNrV6xtxLvJOShzpYk8
5Cl84VBePAxKsj+wADA0vwsFvCvZ0bGKBUkqV4RQEsRk0JRofahfQajJl3irz3falk4dSW9WyRaD
XjdMdN5GFRZX/8lUIE2ZQbSRNYPKzSizl69hQRZzIvJhI2f+gNx+89lwnIuAQ1j5P4pP+IRNNNI7
F7Mhqd3WX+sH6RRB+zYvJ73ByqPRxgMat41vnrwOSdQ95CM2QWUlDzINhr1xlMHhcTt411nOB/5q
FarmKljTk3IWmAsGEdvMfgrAEDwHO3e/nPacK4g7KDmVL0buC/ctTzhzjLlfhvHdSSKsr3DlXcI+
L4dlYM7TF8w6tjpAVq5Mm3drZvX5bb9RP9Qi/bA4t/pvlEbAzbXAF7RRup1al099bClX/jBuNJwo
R76t6BaLAh6Z/jEQDyqn1CmlYCwIJPumdKA92ZJRKNhhnVqWvsHMDh181g8SJwHBqN8iW+zXz1Ba
6tGaQpVr3LUzoEPhPzz3JeoVh8HNhUNZ2SknyXLpXNQxpw/a+H5Klq/Nh9RK15aay35Kl179Mz3M
GvRLktpl33kye3Q3X0H9NPLXbb37ssm0lok9EyF+G6Rgm0N80AAB1CTBa/Z41eW8SF+6VplnVH+q
RHiObWng5n3bEEM82KUZwLwUBLjqAU36BvrO4xI2i4MXEoxNWEOs8D9Pn/BIRYd5Mn+4pfxx6ZjW
EwicSenjAVXK0PdjehUhHPGt0tuNY8wD4AsV0+rKvTW5c3wuqqD4iC9rxR28IUwhI8LO1FCnHcj5
TpSH819UQM01xGSJ26bO0ZPsipIDI2RzyBlaZ4i9Y9X71N4sQ3s8gbw9iq8EskViBSBziRIU5vPA
QRlLEs5JcEvIcJivRl+BVuMT4M2F9Em+05UcwRQkTZtl7GByDmjDdiWMVavvoWdKgIYNluiFK+d1
Z25ihxAMpu6PAgvGD0CORrYTQie3p3zah+B/F1i6t3WmwNYcz6MpIK2/2x3s5laCorakvakccPzf
M90I1xeLAgwRDwkIOaCMw7m+0fGAORmKy/mpt0vWmWRxpnQFnaIogo4UkYlDc6jkQ5BYZiD5gteb
mhpeFjSfsCsCYv45elk5OgOMRLv4HYpVVMCrlhC9S3SQvo7Lfs0U8YH7RAioFoLDJENcZoYLutep
XGZ9l21/mWtvxgNhpnger+mzc/9+WrVDXFP1kuKylGTgJq4/awJvTtQs1bjQ/oQVhWvYSp5pUMNW
QY7dITjtJQaSp7uNuTgPxL+CMqS4YwZTE9p5ZDKSN0eJlFF/Ilm6+TP+d4vUjg/FEcumI0L7Repu
egPKN4Soh9SZd0hQo9I64UAJIzshDIIFKXH4ZCmvIWb80b2f/iuRaTLXUJLjZYg3onv4mR+BY7tj
jfgWbO1BZaORuquNzq9b9HYgq0Tsz0eTTLYRhDYakJnBsppW9anJNJcsbUfCJ2uJPZIzcQ34dqtr
tcDBywMgv3cWlR56mePKVy+N6kwrJqHh10NAevf1GmVtOCkIHbDVFkSECYKSjWrsmy945dNnEzN7
7wFgVdLcqXsf6uBTkIvuuB/+n4bdPkA9KIWSlF0KxBWAnk7ald3uavUNg92inrUexvaVl+1TEueG
k/HlG5vpdQSTUaZVombvXz3xFDZW9CdUIkbtfVrLU4luNelWugdWHrgC3nmfA6SU+Azq9Nt1LlfL
jbL2wSSFEt1/2ID0+3HeAARdSrJpaiAJRbJ2OBElMzFdvL/z8cLokBYl7HOgICBwSk9pcnsQ4iPk
wvVgQxYxFcVzmKyW2RY7u0IHbcbb23Dhy9qTp2l1Wp9MK2m/ZXZ3Pi4NT/rQ7tB6fGp1+d5WtNX9
c7d8EBi4ShJxh7vT8+ccZdH+ycNOSzfuNllsZqaDkiwT9IShR0pPBgv2ECdHleJPKTmjaYcBAFOP
dfqaJEqIc50PFs56njl9xHu1WriTS/nGZFGYpi07Kv3rb9PNdS5I6+S0T+CHhqc4H5heYRnLcJCy
aZi1Xt+CmcavuHbao+85q+YbjtCJEkEKUEhkQbw1p+IbOC64iHS5xTTqNuBJ++lEpw5xyinFFh7o
mwNx9J5Goeem5+NGL4X3MgxPZS7CxhoHkumz4zRqcwVtOlQD+7DRJpVjydU+8AX4TjkolxX264Bp
vHiN7h068hn0YpciVxsoEdmpHP327mEDZJ4hdq7ZJUQLdQNlt5a3H8OKIHwkBhf95jdpBVWNbxih
2GzYJ5z+Vc8hTHPEXT3q+dvAB384ByzaJmrW2j8iz1KVTB+LBxbBR8JLNATahi4WcI1omui6FbD7
ZUn4vZJb0dn1/jz8ZnxtjjFy9ds9rJtEUIgX3Q6e08EA0eMBn73XwuiRa9UI8KXgDDyZKnlJ33vC
DvqLH038uopFgTrWaR5aGUF3JC2Ld2NCiNDFME5Ln4xY3vFenP128e0dmQYLZhQD13VeLboZlnAZ
3WqDp3gbQZDsfNr7nXBA8h1iJGcv2eDZbPQqWPwpSvo4J98+lVYuQRr4yIHWp3g79RCE//WCOtVt
3P3i95uxdT4iCp33gdXu1NNS+MCOqe//9dM5yjGhZ1iQA/zrKKTgWgzq8YJ+KON4YurT7FwE5Txd
aVyCWng4MtmAW0DIg1lDZEr6vBVhWhY+/NX4t2Is1sn6mfRLb7+RFpyqUWqFgUhRbqR895eeCNn1
y9rRG3UT7EltfkgjAPi0IMWX7sCL2H8p/29kn/B8Y2exLR2adCnEL5k8GSi1gy3vMvg3eVhZl1K7
hzO57v7hfHAzgdmOo2EbfM010HxNEH87yludO1nXWooSMPZJBslu2+dktd1enDFjeRZwcwNpVhbD
fhysJCyTLRcdPJWdLQcjvOtGuSyNVuY6nzofbMdimSNXcsqIQd/X3RU314bj8iAi0RnmZuI66UYT
pHh5vepAn7TIku7kV5OK2JXHV0MYFrC7m+qe+qvjXr6PTzs4FiLJ6HCKNC0u31/ELgGKeGCGGJ82
WjZm9uwul9pAyP3BzAwAIoqndvVRa1pPZjPnDTiJiZtZeIRNQKWqZx5y4W+w2W24A+L1qDYG9rmJ
RuUdhGyBbCIuHa92kjlxCZtWpndDg7hL7cKeb99D1NAAOaPpYIsacV+1tzOCMOUvGJ7w0CPKfGWk
nlrGLlmH0RRBwAydUwfmaCcmC1sRbZzUvg3LGBhed/6wtLiTreqTnlNfXJM5oOUa6l+Dmbvk84Aa
uO/JYlBOhwrq2xDZqfhCGghueHyw653leBbe2P7OQVpMkbUMsySty03dPgjfbB7iQu3STuzgmpX4
MEv0bQnVVnkS6yU2lXqRiFt0i/0pD2Eq1Yk5Fnaw8Cs8aALMIqy+RUh+GxMRl5Vn1S5K/GrWiHAd
3XcWHcy1SpuaEehIF8OvRB4NUKWcBdeekXtCoG8Lv8dGAOICDX00cQ0bjXvtzH9lav+x7gIKkxnF
5axFJgA1qeBoqgeUn+dfEsB7Y9kdgFUC+TeZI02FKqMrUZPpW6sBkI6QIJW3JrU+9vxPqMwK7a4y
KaxvXbroe+6V84rkbkuWYZSZkVM30PGKuKECs+hlfyq/rvSrYB1RwnRp7AXfEl6XOAv1Qu7EJ6JO
9KGxFvvon05d4howiyCW0BKj1inpR+epa+FC5X9BEq/9trKz2BdpU2W3UZn2Gc0PMfXb74gd4ld6
SGWJlskRwVsuzLJ+iBJok/0RNOJ0R0+FqrltP1PaNCZLfUcdA7gE61nOBjr4QtcPEnm7Kvwe7FBO
WS16pF7khNlVaVAyULxPfjh1wlFP3plPz6127O+ASlwLokFLR6tRprmc0Twt2uMHUxJ2Pq4q1Vcl
YCO9EXomiaIjljwuKCNKRzFTjUWDwcpRe6klo5hcU+78N+HkfOi/MT//Q62/xgpgAMYeK/VlEgGJ
0KR0qXfu1TMw+kigR/bUweizPU7OzIo4iO2EVvZSy8o/f8u1hFvHomUY+i8BO2JLSDkQsd+Ajxrl
kuoM1+MKOHXyskDHHi1PGr4cKq5khU5oflqrs9uRwI2DF+daqaWafvdE29bOSbpmBMxMGu7xwJ9V
yGZtH+eBmZOcjckuNDbkRx175XF+8s59jurSgcuCEAeiakl9y+s7ysEIkDfX1VMNDyEd6gGAdjsK
xV5/ef2H+yOKiqBAx2QOD96SdBnhoQpdJTjPvce422w4FCPU5+cBvYs9v5LSdTCk0oxb7UK/2VN3
5zgDaKqYN5DkOqaH7ExNcsomOxkCjePBleVwP9Ogzey0O7PkoW/Cew/OacSx2gfunQ9zxKGMqbca
r6PK+D3a+L84Z9I/3rFSTDCBUdY9INQEy+7o+IwSP3XtnE9+yHJEZjF37Rlwfhyb5bkZVaj+spPJ
jgJGmRmNU6MRQoIs5WqCeS0eIXTUNoGC66pdBdTd6Bn7Zhqjgdrwh9vUKD062VrX8O5PPv9qFLrI
lJvoJeKqTT+rh4oxcbbHcBBbGX+OTzbotK7zDP3iT+TELM9ILeMQG6So7OPZQUepdR1nlwJVGbjC
uatnedFlb32nszlk0xFZJ0UxuPxME9h/LaBvthzDXdjuxSO8g5WayT+1jCdCDE2A5ICMyAE+bR/C
HzkJLxhTAImyMv5fRfcCiM+t32UJg8GBHO4bf0wzisZsCjDZazE4GvbphX7JfMIlIc9iEQjpygCm
Rnmi0CxFfdhfT4GwZUY8xyNkdRN8IWcAlAJE5MXF8grht/EJigkQzDATwJKVGra5El+gdXoGJqJT
NPOCc7OTcA0xl3RufBzbEUHYVvb9TPI2E3mWQnNI3rSrdnbgfDpd6iHaooaPsZI3mo1TICpEUH9h
rOYd0nf6XxMzr1PnpXGS/hSFUtxJ7fSaQJPhjgDDY/9Bblt3PmwJUCFRXLKDpChkB5LW8PMAzsWx
7tb0IO8fmleVVRg1IQyXMprywFbv5VK8hbRBV97aPKaiBZIqI/fCmaVd/fslIzfsnlZRET7bH6fY
hSmvGTJ13KW6svsLInwRx3Mpx62eur9gcVDZa06+LPyue8mb6PNecCeZ0N/XyBsWjrNIsnT4XSAP
gE9L+75t+yS1IdOMEvASXXyie+72KQwkrgH2b6H3mtvUs0JLUYCebs3pnJoH7/7IXnjkc1mw5Mz/
H5At3/cFrhfPzvx6b4EL+46pNeVgZwxdkIY177fq528a5czoU+JNA9k++JjQMmGIm6FpSwUxwXGL
jMBglzVwba2n65ypJ/EELoFNGGcdnN4GqO5uW7WhrLuhXwfjYFaevkuPQifIfjBSxF15jXrXtWZT
SPmblJCJT8JLgVraw9H97jUZLBfNrTJAHLL5eWIGXzOhy6jHqBobbZwAvN9ZAQzeXrnFU0pkdaWH
FTt8KcuTtiq/VpefSUj2h3S5XlyZraKI0Pu6RzRscTj/dmKZfHCLKj+R/2V00tTdJCl8Fpm/KK5h
fkTM6OW08IGKTvyky6I45Vb2uCZ7OLxIiCbKzKHjnaGj85wzoTd6ot+7PMAEvUoQgMmVg4zv03I/
tsPOJa1ZhxB0EC+7sX5/89SLKALAVZdTkZpDKUeuUlnlNYLa55Zcve22BATUVe1L1WAQ35+pSRx+
pniiv2sUUEVNjcZxFQoMWCjw7Z91mTHlHLJ0D5TBe+C6SVxngC1hS8sGFIKaGBIZiWHwDTt8OdEp
MLG7EUcCjYXMLQ2nF2UUTJnGvsVydy7WRz7EG+sq3f5nTECaxkY1CLHYxt+MbZGKpVWWA7SKO/RA
M8tIXmmwiK2DvLzXxY322jvJRhEVbiYBnWqoCfczkycolenQvBBNREf5hBD0t6nEtrGyocBAlIUK
9Sdbalm9GIUdGam4vwfB63Q6u0TfzfFmOORYvrFGShGbvZVj6KeIMIS1UK0+pvubW4XmTIKraesY
CZAELYKIcKlr7JB56M/3vINeJoD+nOG8qSuucGF+nAjSYob9olROsiasH01vds0rbgTt7e/chhSI
zO/2PNC31iK3kCdj8bFHVb9OVBADSAnFjjM/73KjJNbrYnH/JcDVC5eVKJaGpTUQhJBIBF1qAR8G
FhOX05/qhO4Pbj9FamKYZCIp3PLYuV3LdF3ON/4p0acmecM8o+ECWp2WNwqJUewYqTgVdXXTk3Pt
Nc9WdsJUJP72AGfNknowFqprc64Cii5BEiy7QIFv8wflaNjk68yPJWhRR9nu9LveNoUWl/U02ugV
jMC22Oi9sQickieExvXcImUXxBqt0LlLqpaD39LvBLBNW9umGvUoF/Mh3VHhjjlJ2efsHnCHVwA5
PAUgEWjQt6UTBfoYD87vIB0WjBJ8V0N7ML59qM/s9caDzEaoP4naAzSurFwhkat0RIiZnzF/sKQx
XE7CYBxYP9bAF4x3r01D/yczbOGBs+IK5DK35tA+nKt21XI3vJbPFTymAT6RgP7Dca09ZygR+zO6
JM9Zn2igvHi+yeQUTP1JVZEi5en4PqDa0FvyQuBluKrPCpPoUXANCL8Wvo9SiT7zvU9/ItZdbHMC
/jr8RKiaVcU09hqWdvaVGrhOzpObXYgS7Ara/mp9Ma5I01L95oKnrTkMzyU+F12hkC/R1NskTlEc
xrge/jASuUbmVx1TPCRTO33f/wQ/111COqzLJMXZ6QZtLx+SfPbFalr7p/ctmJJeZLpX98gmiyon
QVti5/Xk7ZUi3urhfaZTBCG2i4oamOoxgbZlmrppZbyl7DgRuBcRUe5lStMnbuix0ddwls14Y0au
+4hCgYG44L0+cNp4OxzeOGS27By6EDnmzsvIky/0GvIlubijmLT3o3deZymZ3P+5M5awDF/ORr2d
XxcmEZCc8dWX8uw1KdDLlfOIzcex140JESfS5VfKsDtu1MfGTvESm8C2W0hiP//RKRxKtSD1F30f
zVt9866D8Snd2I3riHqYAJ662Hm2z1IFqm7jkPI/MgHbM0/XWWTH4zH55EZtBl6Z5u3yKov59f0Y
TXZyeTOGVvo8ATFVLNrB8yzeOAGWmx2IZsfKIX6gFHODXWHJYiD2b9Yz8dIYFj8PTJBwVtwPHbGd
v+Ge7BwGQe0C0qTFvy2RKJOm3B6+xFw7SEhH9prJ5pSS6xfdL4/5cj6qIXrP2ldeMgqTV45vOB1I
AxQCvoGGEE2ub19tyvIgLLtUztagLFGqowVIjsyPt2QJwfTEjb7c92QUmbqFdv3Spr7Tfytyorf1
2YBYDVy9CmWzHGVblluLs09SKg0wguLwUvNshSEnAo/skau36adniqVazj6NQ1LcGKsXLHjHtGdb
WBb0/RF2e4lfHfzi8oeP/u8nT9uLQBwyKJTneNXZasM7kx2ovy3hDQdSfc6lnVqo8wKFckIG6j0w
u5jGbN8DI6Q+dZOSywSOizBAOlZo6QnJzwpFrpv8khs7UTj+u4q3p1oMNDqV9D9qKsDo6B/LGWC8
zs5v5vb5e1Jqwo6Az7pKtT7WkwYpoMbyeTMsvU1oOXMK6uSlWyxIEZcObCkSLjomoXYMXcHcZqCk
fNP8qdqQYSDKuYqUL9zhwYsIa4FOLQinJLJvj/1RdErqV5CLW9e8hnfEuSNL8SqyDzkhagGIcA4B
iVyOiOXwxHsGO0s331uaaXYtxlngN8e+JudlDMXUQFJMwq22p490fWdFY+IxdsQvfoDWg6MthX6f
8M+CFyesCTv0PhwJcjK/vT6QnVGz2SCE3//GAi4KdvuQD+5NOR5ZPUFLnsSWzIE5ev4hGZRuwE1F
yPB4RPVWiyUJiRufZNs0DfZnWLbHOSBmFKMgVr1zg3vNuZXssDkO0BAQoAWOTv7soDSRy/WP5Av1
lh9NOiWShXuQjLwlTVley6cezb/AK3OaLZR/4qH1bkko9nBAqBvWvERV/3L7xz/6qysXZ1PM7BU1
z8FwKrJ0JBm4+VToWuy4OetaS6aWevoZRY2OTSUfjS1MRuB2dQ95kgnzag8VvkrSr/Wgu/BQtu+C
tWdMUwUobtnKm55s5elkxlsoNGsGD4qYPOdeoCragggczctsaHewvkcu02xmjkQMO+lvajT1cyri
+cQNHVSsig6stL3fIcc1/UUnciNEotjoOUJfL96ZGFOW5FuRbkKMoVkYlppIfW70lCG086f5Xgit
fQKitKtHS6jX4IqBPnjom/f9F0iWnI953G4o93yJVy+PhOdZs3IvIT/tb1bwtf+z6jr0HTLiSFix
jUMO1YD1+C+EbI3PqqiD4J8BOHqhEoubkCrWi4J2TFix5Mx4uKGESkZrI3s68/DGismIPbujZHhz
csDv+BflPUvlzGgK47fv1NjIL4la9TZdKeL45Xy3rYPllAAxLp++wHB7W2ev18v+fF7jug4vTlUm
+P8a3vnQyTp6UsCYfuXqAuDVCDwMEsM97q7uuK7HMyunuXejJW6RaHfc2NT/sJOEiaO6oQ2CRJQi
nzQjmOwoPurJCqe5iUkBHAK9DmGObGz7jObJo/IIt8quUrETqpmS95reYoeKIBmzcaKU2BTokPVQ
R/AiGhLy/gwUvVWwKtvqNBlgqQ0qdHl9FLVjdi+40bE1ynnJSKFCpXQ/TOWVoTEdKR/NgirRSLfC
yh5xAmLsFaBue+USQqK8+lnz5LQNG1bsbTNO5Dep8TyeRGRzsUGrk/ms7emdCmgdZXPCJsPCf29U
cd1VV04EyvzjoWW8ngFveQe4uXPa2W3mDoeIbhxC5uok7gDBNLjtqLrbX/WOnxQ9aXxe/+t1qVwg
UxWDypRa0urIX8fGHZEnhJNBHpm12br6ocOH8B46lrbm3LTcSZq3Cpax95GaqCFbOY6Y3s0wx6OD
DcY0v/xXJ6s+dFuYqEFO9lqG/M66kjwB75JpoSX/jMCZiC8k9OjloaDT946QrdUG3SOuSqDsXf5j
p3ez6KAbFbBNeRU7+sip/XSEmt79VDCUQBhHsOg8YHdr+McJxAcoFGi1f1rZTqt5rrSY9iGLUJe6
IzSyi+R2eV7CwbPV4mVlp3EtFHbojYJ2yDP1C76oSsumD/FAdy0l++88aNZpM/gcVDPj4F9h22aA
2d/pPBfJyAcQnRlFUXrZ+ANfxSAfoVVGbfiRvbEXZ9aLAzgUUnds0FLGb+oMFc7pTQzIHAeItNCk
WsBujzIxczw9MbQ2dGiQuXlJupYpyGUHwLzT4s5j35eqrPv822NxJW+HvASdxisax/QboeRugAsk
XxjUV0DFluQTWln7Ui/bWwLRk6R9IWmu6/XXaU3/Numgr+pwPMVjSqctg7Alogj/Go7VbigioeB0
sXE80UcwhAFfSFfqyF0QoK07vwaCfppg0XhB1fsM+gQz1mdJiws+5obPGYSK6pVU/R7tr6x4cdo/
5tl8St1NYiELSU/eg2b+msDGom2vOCv7uutRrHlU+6Orsmpc5n8TQw/WmpzrsAElBOwacPfsS8Wj
E0trFXUyHdaXrd5dRq9y8SrP1/GNbjPYQBLau9fCp+eyz0/yfMlF0/9rLFkwQTrdrVOb4WPSs1JX
ZLALdW0WMk+DUE6vGAX1IomUrfXFhpRJyaALq6qOVCH+kNMgOZeBgm1BR4U2nynAtoMLEzhVxpDO
1GXkFgIjfZ3aj0/pVr6VF1pR7FBnXUu0kvdHwr7QrpGa9VwUYRUbnpnMJN6hKBQdEI2af+5U3env
Jfgce1bEscKM0ErSOgRfL+7uyIrT2IvUpYJ9EG74mewprvCYJPYvir00hw3oIgj9CAl3Y1fK/rEs
NkbLtph5wgnwK7m3VkVDzb57IGycp5dO63m7HC0Ua/4/SwgF0MSRBHEKJkfPPnQakkSpwoVZIMQM
ywTfuxGwfUb28Na6CR/LBKN2fylkwYoX2/9Z2AIRD6VjdOKrF4q4k4n1bi7DPl1bAYLl1iain5Zx
2fa3M5P7nZw33s9iRtM0BXk2aMaTtvjW8r3MOIgQeqRPve6xwIEbulkSC346vWTFeqv4oarDm/ED
qPG+OhGYLYyRb6o0hSlAOooxy3kW4dhySEKExkWNqvVQsgYQaKxoziQZuk7h0jeYRq14s002wf4s
GLXGaA0PhpFyHmsE8dx1C6B6+Cmq/hZbuQNaJri0E5TftAcOACY5AquiXgFPNA5+n6APBDBmelCk
/dpitimgz8LY4b+7BVZaiMgtUzZwxUtkWtHpxcfZLVbZe8RadLnTWywOsbKf8p763DqtlQOFrrHE
F80XyGCTejjvJSTiQ39/RCTFnn2Pv/+SX1rtEmoJyBBfc3akO1kztT8OLtT/0EV22tPnLiRggmbs
KC+htX6K8tdhItS7Swf2bOLx8xx6q9X7XVFMUdjdoftA3lrxP/6eQiRTSgJPnpluQLAgLWxhNv44
l5TXLV8Gacr65eZx2jps/xCYh8LRd9d6RqmdhYLZa7XxiDdWS9io3xhDpygsTKnFeRop/bO0Mgmu
hv5fFSaX1PPvB0Q7JADl/OS9JcCxHLW/Ww7u+ShuGN/tFW4DRACoV35TyH7T5aJYNcfqMDdbbpjI
I6rLlx9VHaUl2afsOUcaIN2sl0/nJnHz5MxC0bDMDF6EjBBc16RjssyyVNfrF8nQVge5s6ti8ajY
61MP/P3byZfaJn5OWiNSKwtzS6FrS67h6iNrM1RPALJblWG1FWtfD3FKRvzcHtRgRXk+9proy50F
YCZPVFdnc3hZxfdlL+FWhi8F9lpUSrsRkdEmrsNy+1MN1h0JhqjftR1zv36ePY4OJTusY9p6VDQM
NX6eI2Uo0uGCvZMzRUr1mfQ0CPSL+DE1y+PUO6myEdlkQVpdxpxar+c1VAV5I7L35h+IFeJmSI0D
R4ovygMnLEHOR0MeX8/t41WZG7ObgdSrrcwssIC0RfNVYjAVVzt0/Ak0Ql07nvVpPHkFJchKKfoD
pHS/dKS53pLIaZS06PTe/m38MrGvi1b60m78rEdh+lFZ08BqFgAatEerTQf85INeEmSh0aVVYUl8
kx0HFJy+dZGsR+nG3nkoo2Yn47UI8JYBVj8quxuNxRddTJpqwnmQWsT9ZhAhtZ7inSN1fWSLle64
tE+OuKhDwwQYRPZ3AfX0bxc7Mz8f/IUJgsKouzpMXEse/2qvr6zdrODI9E3uaUEP3RxDozcI6dK+
rQE/s+P92jxAIxGTo38tEMDgjQD2Dt4tbADpGbyyHYc+Y8stAQ0XfwAztIqk8So47kq0oTs2eDmq
6s+KIAlC6G5l5lqB1RRqdQHpG/w4Y3EWT800QfRh8AqqGzJcQqOONkntZLbQSAApT9YkAtPOASEH
kooQNsXKkXNRLvkX/4K7uM8kv8C/QKwI/WH5U5DXjtenvPCfCN3KZKYV1gb4PgGLTecSu9ImXMiA
IFJ/qC442xX9WO6cU82j0PhauBYtqyapglEMAC9hMc4mTYgTMGXgINivfHJ0qyUhCbuMX6bB/6k9
k5KtC0Z1unSnH1HoDEhyGdeCLDUrqJi2GNsVl6gc/9OabtqS5g0WaBC8sanSyQYDZdMrRK6se9Oq
n3Zu9wt+bzIQdMWd2RbeVQIM6LjxzcRPoiG/nDCgTU5Wb5nvNCB2ZKse2kEivDDXQtVWRQ3N74Sw
L0T5njR+H4wG7xYhMPX36cCAP5vmawMzTAOkxMoIty1iEqULeuxpNd78awXBA4oHUG0g/DNY4THG
LvyYOHwlEwL7+IARTFZgs74poS/tBdPzrXuwcWEyAHrTGQARkwjp8/FCwRnNpUmJcu8v01JwicYO
yO5b6w2us64EWsedOebgqr7AmJtqrt4Z/M+ENirDzuBUY///XaaA3HRO8rpDRn8mVsS42f5O6/cd
HUPltBtLOwXgAYYg18NKRNWe1sQtZNaxhdEyW7ATxxKARNWpiy6n3Y2wJEJwSN3KOcHyp4uus60V
l4TdHyOIs2GT15EcJ6M+S2lYCECbXyshhy021YcCyUI11aFzNL/nvcD2uLI2dbm7ixsnHdYuc+c6
VjKRDizDaBBLDjJ+DwurGWDfkHVs65VNluRdk1RxmtxT5yhHQL8LdMwrE7uAARV2vumeamVwt0f+
1ud17r0GUOW/hAA3zZfLC6qUtOpacnheOZbqCAkRKmvBbHtsMnCMgrCgCja11mSMLpVvLS2U8X/a
Vn5YtUzzgNT3XTBtd1Vi4/0CZgNnmSPfJhNTHMUlhNt15UQDtqBMmsryggmzcz1riwfo6WpAziub
zsS9dZZ2L0Dmq6sxztivIUDfdootv64EBSSNTTzr4GFTrRo1vshEgP8Of9frAmrpv2xD+/3eIYFC
CE5RK9eZ1FwJOcjjXUL1WBpcCJ7AMRheWzkKpHQQUSfUh6vMiUv12IElBWRqzFsHMfvOJABPxbU2
/8WJDarmPFuKu6qZfmiV/RWX6crjSBsbx9XUG9mPKwMwwbcxL1Li5QNNu3w83JDd+Oij3uVMA9lb
uDNOQWZUBrND0F+JLof9Q6Z/sPZrcaVrhuzL69hxi/ikMKOi0zg3TeSpCCjZrfiyG4vdd1Un2AT4
xRITDN8Ic943jqjBH63XuXYzS0yqzcS5MJ80PHQLgJcRHpWml2Hn7SBbUgMq+sgGjJ0KAQBCsL1Q
Y9fx6vCyim8uKnMW1/7jmva+OjzFPXDhRme94JTGp9cN4iADvTfPBtYMxVbTy1pbu3zzs2uto75V
k2RN+AYQH7+oaGillKAKN4K2CGjQi6tvlznEqOv/Bc6voxREgnMrHBMMYb1+YICnD0uGJXZ2TrYF
sFmtNmeMdCyhyP6ru5lRF7UpymitlaQC+V2ZWQfiDolhzJxmZt23s4YqM/j8uJB+3BZpxQ4ctfTb
5j1PHZoWV2nM9/46oQ1yCqVzhukEKJbzb/iSbbx3nMdZAC0t1Cnvk948IdlFmAhoN/kdr4ddt6hx
5m3lIrpzEGCvxIpaoHnT+iQc1nNjcJOaJ5tV8XS2k8W9RmYmme4EH6HirW+TcmjA4feLJjajWxJ6
RPfS0oTCjFEJh0zau9RX+7RSqtp+SBCeE3KD+THbb1mnC/06piRDwhmo2+lX1CqYKoWqsu/6ESLs
kOOGHidycRI6acRP5htBzBFvTUS+HKSMTwWxtcxU6X1vuuYmkHjDOZUnpqYB4q4uuc1DNM3zOt/i
Wnamr1SuDMMutCUkH9mQSI+qmUB6h8HcizymGd+ZmxoLOXKJlIqsouae53d8qC6H2XyzLYAmxH3m
eaRwkgM/Jy00BZkDLT0np/XIhWdSOJcKciDUSo7Ev/v/CSYjtp8pzkjE6Xixrkg8JCS4VELvaffo
zUxG7yk+/p0oiIOkRzL4mViOfG4mdFQycFfbhIa0Zzr9vWMHT9/lCUIMG+k37qlZWPxycLImiO15
LuSixLIauVeFewd/XyboHs+YF59nD0M/D2hTO+M1uMqG5bOq6B62qZ/bdUAXuAs53keUo28lOV7u
lqGLHoyVWcySE2N70rrSxCWlT1YzQCeGZoLGXw8ZJwk8BOUoVz2Xi3H5l5deD0yXzjlYDedMPEjC
ktwIiRpQfU/ohDF9ZJ42KfDGekUPbH1/B+kggvm20Ja8M87stogp+eslkKIkUoZ9h17uWHEWG+sK
ogKIX43mrULsrb6h0oVJjd/VdKCRHuC5bIH0rF/HsUJ5YL+gyEhqPDtfqyFUtPFPDckIedeiEomT
i248nnQXsf0vtlpA6PlE2VDY3/LI2zpG4NWeYM73M1fQwAWh/BxrQThttYR8KlqAy97BG9Wqplp/
oYOjRqUapU99TAtxuM6OnKKHwf4HRaXWxxiEY8p9MbpU2z++z/pmZOmZhlsrd4xH8/xJAdS9XcWS
rBonmdiDvE9lgfi+4nmPYhBhsiXSshKHgm9qC/aiwONjtnCJfLdnH79mh/ESlGXv1ejRLmeUCM5C
ksvElz3GmSosaTtrjEbHboOWBCfU8X6m3bLxLCC61tisuCaNIMLI8+unAiObLH3wK13vAN1VqGN6
aRS3wUaDe315jE4UpoZ/jPd++Uzmheep9DWo4m/bbxwRiWGgUhQeTfFbVpRjK77fYJBX3Kqagy97
BsNWxIF9UDQGutF+HMWqYQQHCE3h0iw8RWL0lxJgjw/IHx5LautnXYIGJMGHXglgjv2s00A9e9rm
Lw2i+Zrx5l9DGlT/kZJi+NR3CQKn1bZWMVZTO8JoCpb/5RjVLDxn0qxctDn/ITRlvK+R1z9NY51p
9O/ziPk8Phn0ruHpUqojrYi5wGzNLpBwpYQ8G9vxxa1e4Tg1tBMuDWu/6muoq66t7wLHqKvtBREK
yf9sp3RqJSXsV7B5PR0Pov8LhQf6RPIAGClXykX8WNaxNiA7F0aj/6TVEC363LLNEiDEMR/KhHor
mGn2DbymFHAwY9ydl1hhjwusbUF8Q6dRCrqpihGozLzFBN12T0xCtqap7HCNVLX6JkiVMx4diTyY
9QJoNwvu7fc+a99xayGZaPSja4DqhY6A+p0B79FkwnI8Un/xKA0zMkuc6qUU4xhBxj5Mn4cxvl6r
hIhsciEJ7bT1Ya7hYzQ2lOt359grusrR/DamuLzn65SPZKjI6jl8ZMmxe4EBdr+FwoAFnecPQD2y
bH+H2E8avoB9wMd1yv5ORKN3e3/ZEJ5kqx/pvo42mUwRSncVoKmoIfieMW2NdU6SqYJ27gla7+BQ
Odb4odDlAszPJCjDPpwoAHLy/nmBGL89m5L1YQGuhf3SVmcwdUWgYK2p92O7lKpTN08JJpT1BHkS
Kd00iJ90d1czQrkzl9ikFbjdOWgJKTosWy3hkKfo2bAZv0wAfVrgAratXS8uT3Tsly0q3Rr4xkvB
M1vUhkCh88GbhdCVWtDUhyZpc4v6GZ1sxK+aPUqvdWYTEB4TcxD3f5u5uU3uR11FlenShtIAJuxv
jDfz1jfwbHY3X6/NZKQjTUrQgQDr9nZXtpCpWs68ka6baYAtUTd2RjIaNJx2cyQ59lKBFUmzvuva
rwteiIGeydF9oa+yDTUWPqLnTZKSRcKQs0esrUX3Rf7YLfg3ePStphoEYKyTVd59bzJE5JBnLqQq
qmviR9Yv3BlfmOqRgDSc0dQmW2L3OjeWEJx6X6XAOd6LMxliSXTsaCLdqn57lwn657Or+pAu5EN0
UcMNJTbLCV/cSOuB98FFGvmeJAITKl6m67ueoSHMCmsdZlONbHVfBA5AGZZCuyZMDLu0E3hHIby1
uSEA+TU/x2av5hhA0supqRhHDSRdeBhuUpEpxZxo990Rgq7yxT7Px4x8dOrW3Aggxinv5KE5vZxH
0Tjm9yxnVnHcYd22DpdpHcueciiuvsOJTG3GduB7slJQeoubFN/smbEtBdwCns5E7aBvr0ym42TA
r4b+PTIl+ysq9l+E2zlBw56RC8raO6wTypTAlvtr2SzgIi7J3cBQmBVivOtwWKNdcZseerRSwjMj
lTFuGyaJZZUQE8HXAs2iu3r2Nt4PSPv8ZIyt3iLhg+z/oa9ZUgRBWTUd1BZx/jHk2RcNM2l2wZuH
ZHIRrBWy8VCyKsHtwZTGpNydodZ3rng+rQUm3th1M6FUjOys5/G93tsQCWI0eEWJlf8PUqb30XbM
SpObHxXvatTX3Jmyhke2YsO0inqIW2GMxL+ba5flVcyd/TS/L6pDKOFbxDytUH14JKQAPi/iAKqE
c8cmK+8uqtjAqgoQqLgOqzYOz2kPRYr6EoFLl8JZnehwfoT06snZ/Vk3siW3asLlg57G4F//SvBL
3OVyubWGYbgrndwZC6+Scp/mzipKGn7Gk+Z7/zY3hxRV86LwvLiyeciGzNwtT3g7bMeFBJxfTGZ9
RCUM9Ao+hTmCSUYmjkQn5Bzg6Y7oaFmJbdVaG6gompwTmC5D6cjPyP+sH8D10wtO0Jarn/TA0ZyO
dxc7vBxWxBz65R1WSwjxNAYDz3/e6sJ1OK6CDT9aAXrKiV0+GNZwMBvdZu6UA04E+VybT2nBKVgc
yktz5hhVdBU8LT1VgA1AnJuws4wbsKgSvjkjEKQHkSMcBaSabnQMrUuUyBrs1qFqutl2a7pifmvm
VqfHS0EKnsC4UhD1m8wntGXD2764qwDSKLGcmvaiB10CLFIoJ8JjldRBW1ljr0ZZkVhxPQORPY9p
gfslwP/en/c7hzPvQLM8aPlCos6hjDCAuZwb2bLrLgRiCurBPgxy1ZzXrdKrhD/fwGfsmBEQPyb2
ZqXWVgeeHMOa6Uwu3gMAMs4gcRDyilC7+8DuJdTAoXW58DOLoB9tEcBtSwstHE8tFHMLpBLLAab2
4F6G5ahMSr+q/zaJriDAWxAto0iFGqWtcsba10giVhwQyxIWcNHeo7hvFXFOD+xRS1yOa870TSF5
3c2jpRWTTvfqKIglLEVDvzpR75CqV2zKOMNWmBdmhAHo40IHy7B2nGfPYmvOcnJxHADfJXhGYebr
LGQlT3loXyrDvcNHYl7wW31QXFMA7+cBy837sl4iEr1bZbVTOTBsLKfL3qoGfeHD5b3MYpRTwLEv
ImHPjVKZJ7+FQU5D0PH0LrU8FToIlfdemMVE7GHBGbB92viimLeNSDopMgklyP3zWNzwIIHHhLTu
W5KN3ON+/Rc6rjGkS1oqK1/Um5UCkjyDNLGKJ4Gnxi9aLg5rJjW3MoI3bL14QBn11Dv6RRyPFpEd
w/gKE+cXur3XpTD34049ZMHScp9Mdt47FnqmHMS7dOqcEexzlp5LhaMkn4721bnVyqoEl7Br9Chv
4llr4ULjfo+0a8IWqr1Q8HVLQw0FbpXVbpYd6LncRsiRuyz1yw2ry27P8QTTdqvp3XMTipol1tlc
TaG+N/ZenX8OQPaJLy1IhikqvHD0g36YHphx5qOp5XdlJz9TZ1/FA/c1KjeQsPtQ7dSa+rkvT8Pp
nvPfmuQtKhFnNxTinTzMCb77FM1o6AqSmbez70BWGkGvGc6UVA9m4pk5uiOUOFrVGAflz3YDF+NL
6khgz4Lt0lFB4KWOkx1PgTvNDwK2IM72loFyEpivNNO2djbxY0audcxxNd1fdVpE7sFakZElGW1b
XqHyQb3ISmRTuDFdbtiQOQKgn9FTbRvuoRnerSnrAxq3u+OEu/TIKq1v/0gOjrLNiZi2Z0BzfVN5
y9tj6fjwvIYPyvBNMSQ2NDiIAd8CcLOWxY9gNi14+nnvC4fMYyO0dwqUYPk66lev8z1XtclEDytq
GJK4XEb47HlWg/hECSMHmd7ciD740T3oPxL5MXECZimX0+STIb1nwZRCrXi8Ne1r36ta/cC3J/FG
Z59iX3j4BrD0UyvxBINv9vAoOHCsEovS8rk/Nzj+iKMdizBoDYLlaOex1IKEMgNUtaQlB39xhAHm
kczQZONIwlqcuj5CiHHec/zLCpV3x+IfkhWagZXI0D748HG8CziOyAubVfqYm6YiE+yZ802Ze65+
hygMBZFBNVsuHUhGxi7ARbT89q6tuNikizxZJbxh2TMCB6aKTSMxeEbhsNmx7KJl97Ghnxbne0NE
6urEPjPX3PgYrzNOeZAygXzVaKJUN8atGhnOYKNZyc5t0E1ljrXsWoeBPkV1j2m5KrOuu4fMBSy5
tFeV1ycXtsLOp5xINCGt4MerDvX6o82Mj7eB9OvcuvYQGbWArl1oTo6QJoQHc2Yo4hFPpzU76qw7
xMz58NrIP4sLaNJfT6jMob02cufRtj3ic6DjbOqxjHMiuhA5Mb6m1t8qGKCEh3auy7XDOqP0EYHe
/ftq5cqigOtSCbnetwaLfnTYB2GvxKgtHrTS9btJstuFDGfDxRoT1B0n7aMdQbt1sFsFc8VgIk+J
pqELHMnZSt3bKFrEO9S3F2iYxMsKzB0xzf+Zt4XXVwth7J77DsPAqIM7WvkVLj4cOBJy2+51F8+q
WUVbjokCMG7gWuXoHyLgaPSAM1KxnDPhnMyTyWPiLhe1Ecc0ygzWSzS/brt3MOkzLmU5hjQXx1PX
dYTBijSBzAxaTyhnoC7TVG/VJfyU0E5JuZm9svqkn29ELJtgn+TjaxNmmiAeOPwvMqgfd2KetCwv
TvXrfo+koOvfcqWNNK/p4B7qe+rAp5UpJGzpKAehwaTXMkJanJMkHpiWCNCn4DprE45+rwDQ748G
EUjjwEIgd3dy9nGf+ci3VFxgszekGiYvXguS9vdGFbDEcqn9L3M7HdEeXjBmc54u1cGjk6cwC/Pr
mdcMm9PYKm95HRo1BYA/o5nhGJkadBeIUffdS9LiMvUf/Z6iR94ku2x6atj4DX/MyfXwDWFAskpW
y7Jy37LgLMtR/zn7d98GW0m03LCHmOc+y/aPaG7qAByYqfULOwaFshj07nCNHDw78zb5cwavscyg
xB/AlniyCEr+8VkwaCQJeFOKYue9XSjMm2OA7TNCPDWukoaEBovpjEwl5sJNVTJhr16Vk+xsS+D5
dpWcnVOKN6T6LiDxiJb+jOyRN/DIa9BJrG1el9ji/EIfmYyaUlwXcTtpmzyynRhAY/XtIvAgjl04
Thgcrc3tW7tqjQ2HSXPqoCtkWYW60uv9kFmoAsJ1qHHNrlfDHgVlwAwc95TBAam3epwCmyWtItEX
44LAC2sh8FYPiphFaqPVTs8jj6u6U+ISPlH3R2/bL19qULM5dhoBh0Kkl1ygMet8rLtbsd354vtA
vmqjW7iCbaU900Cy9T/AbFBgY39uSPPFLhsmOtXzkXbVB+JUmixdSH3pSLCRsdeeSxIpXmrpgVkE
XV/or5B2mkEXScOwbKSEcXeIW9/nNoWbPktYno5UxLnjCia8SOjfbcQA/OXB4vF7JzXHZ06XLNdA
d5HogvzJO91ure9dfirHbrPJ+sDuetgU2mPF0rc/xouz0U1snvEwADc9GUhXUWMLm9u18F8wwbze
bqHBGq3/8U8G2+YpvxyvJbrmhHzcngTeKLe8gWpV14nrp9AaIV5nhO+zKnHpRCLS+pejCXlaw3xy
BUtKyXwCUqt8+l+8EZVtPhfDO3kGplek1GMWMIVjkfpdWX4k+tQtT3jSKshojbUAd/KUa+i6GYjs
nDCaR9x5MGHVyWDBQVf36cBqvlMRw6/KLi3gL+0pfMrzOr8KeACgteYbbc3QqoNpKU7yfBfkE46l
VZI+7T7qg6EOBL9V8X3ik4fBBZfP6fy6OtiVdUAMgiSX4Q48laLUJFT2E6hVI0k1gF4DkW8gBAi5
caxZ9g/GhOkKmx8jFtDjLAL5g+CLEFOUwZV9jM8cSfRHOFJF1FFDtFDnMWBi1L24gHomOgjOm092
H6wzV66uFZ8AOB9f7u4s68gKyu80RMLTNBcRdpvmGm6bUzIIla1UqbZ5oCMpEfIWqvRsYmU7bCdl
T7LsUFxt+IsWwI5cJXUWSeA0EuWNAw+XnQMi1CEwTNRxIKvNsfkgkqzGEOXdyPYlaDwM420kYFv/
Y3T3fa7zUgKpBjMSTtjOdI0e10IxCVD1J9smI7+FAAU+pRGlkQG1ae3HUVKBx0ypFutKZhJ0tdmG
OaM3qX2DWEfd3zLyOMEKpxZGvFX/Tj8wNCFX88gr2wUyapXqh+116P8AygKsX12NWivU5JrRnT+Y
5uY88KWKZfbk61PC1URFEZLqaHhPCTUuIw3RRlGicpSrx5JuVZl1yxFErOnqbeH0sitblC3Vqyhh
iCPvocps8bRGRfOffqamZpQNl8o0FYuFuGlOFQ63KriHJGNWrSKGXuKMe/hjHsz0gBQh14I2yWyY
GjvLvNIHH+LGun8PR/oT2yZFVl7jiHNLc5M1mxVXkGUzUmLZuXWg/vBAS+nLMRyXq8rYg1MWCVj/
dHpTDywPz99IZb+aPsndlPRPbi+UmhTGDUa1DuGzFw/LHGbW+RxVIFJV0OtmeD7vq3nydWBp74bX
Y5tQm/LXgP6VoOubfBJVazeHXG5Rzfzpq81BU+1bcE6GY1x6F3rwJgJA/InhsnwL39JKEKn8pr2j
CuSk24Ri9fVfDNihYofaMbGQDW0/EJbd+vfzUM74iU0VmfQngPhkQmI9RPA9GE5XnM7HviNZPC1G
B/ECMtloIk6WvPb5NvbJNRsKFFZN6s/0NGH7Kld2ukyulRVeMgL7G1zaM2V/MIhO3CAZg2+7jI8X
679hBuNzvJ9wqytwTbOtHDub2i6RXpOP67C7H/Pj8vhPMZzk3SzdF79fjgXEmIuN7Id2Dw3NVc9s
qFpF9apcdJRZgF46FP3gSGbaeuP1KmItdKiitNzQrrvyRlXe+nrgUOTVB+IEyN24Uq4A2bOchHrQ
DlQtipO/VJCmi7Su63alhmkeDjN16EgB4JTvhYuLBEHsFeM4Z94Bp/o1wYtRHWnklSJTCb0pD75Y
AhqP37URCmVyD0nWCDSLBTyNjyGMYgmgezHbuN910HJXlhLH9bt2hH84MV/MMJK9GiZeKGetzf3I
SJvndi7hqbnDSXpx09G6zpZ9Ows6QjTWusCd0kmcET46fY8vLGPR7ZYUKwpB1CPKwr6NeXyHoRZk
WS91BC7a8o2NiLeH85PXc79Ix0Y2o9FoHfDt4VfahiJOj7xq75dlzvq9cyMTBeeLKeXSG32xQfuR
8YCc94YowJ+e3WRp7ym3VlWAkM29OpHydc+qc2PxEJ23yXhcCpkItVFTEWKUyg7unDe9bvNkxHtT
cqAo4jjpdKcjELFXJIrt/reAhwnF47lpUA6kaDduc7lKG9Hn3Tc7cwneNGdFRqoo5WXWCTvdJQ4+
OoF8WyxgQmPbAUleygAxhEp9C+ejXVqz6KefTzbjgWWcfZwZ5QqL6gxvRGb8OczzMdS0lGP09nmA
Wi4khiGuKP/jJseEoA22tmIdm/w+Skm3jUCAG0aGEH7gocwWx+0Pb0EHT2XK9REJhJVpC8IckO3P
YV8Oqkp9jY86fF8t365RWwcPW4BDAcCZpcykzm+YkvjMwGsh/3YKs6iIyJJo/YbAemtANIJIzJV3
grZUoEkh+U++GPIXb9PqACDxTP3ylkbZopcYfDhfSuFtF0FUbj0ZT8eZ56MRgRelmjac582BBP+R
W2dmyn/CTNo7Xi0SHUcRj3l+PZzprFqXMstKPFMVyuhnPGFOvChXWA4yEMfb0NmlmvpOz4HPJYRE
DY6xGZChlDXtA/BzX+CZjzsp3yqbIYAo8IyCE5o71KRsYs75J9mus7NRHzh/HOPX14LYMYMl9K3G
jjENfFuNxjNz0e8bP2+LjpmsMLsOdSoyDj/f0k8+E9LBf3DogcP2tx+7i1OO99gfC3WYqf7fNxtb
4MVdYSjSWVp2KbOFj1/6givCbkr8r0edZtza7wnCSJevgTuQMY2PYTrL1bPHO76qyIXliXvOsm/G
yHokqOXYDUpleantOGPpFQZ9P0yFJaKYck+mwaezOYbtMq1fb5BNDO/2g/9GEpxANKJtOaDsdoBo
4iH6EsnbpHB0FFVZISJXFXrOiN95ZOEoollukM20fDUSLOWD/wPMQX5cLEOdCjSmj5RxyJgx9NDy
8SEX5jE2COKi0+TgtQbyZJ3Sz2KHxGV1c19qxqiS9AwzWIDRT+Akp45MSiacKIVpqHl1tYLosvYh
5+Zu5db5PDaMXTLlaeUt64hF8UjPa8MMx4zQevjAMai+1Y7HV9VZaUelOUtTiPGW+QpUL7v57O1w
2CGdYX8zI1q/8H99HF39pxoOZeotN5GtUW621AtmOq0BPVbmp1vMf/R5W/MtDeVzT7p5C+RVcHNH
sZucXCfx0KiyFrPOhD/i72U3iyMyEHUWCnmE8yryTZ5nOkMcY9Wo8nW359BekTLi5ilWa+ytGvC1
zSdykW9LPnRvY3/+lnBLy8wpkVEcS7WDDE7Cum8wmIPKb9n7Dh0cCyL+zEVhVQkiOayHBOHX2j0M
zupWJkMa28QEymBacVuRXZ7gSOMDDa2o+IrT1ftQW8K25KxvHebcfrcaYP17KaVNmVQoMele5Fkn
1jCRs1HUqYiJzhhXmkvOfgI6vMCm45nBkYhi4L2x+AjB99APjYDCRqwV6zRndyG3Dj/VK0ZRYtf/
DdG+VQ++VKtTqBgQjjzIQhsRds3LJ95SsZW4HK3feLqhd3fZjWKyFEP6EAED1opqgU0MRO7SKxye
h2RXb/toKAJsVukwXYD0dE6GK1xwKnUnaYgx/6WU1sqTeeRhXCBvdiCOqsC1QZM/MLq3wVUD6m33
/Opvx8KYlEdn40yNuRGusWahwYVagpjKvrUpdE59WMWmkUq6420OGKMQeIbUUOVMZdIVsSNE8X9V
UbYZn1zOVatRCUtncjtPNFKBBG/kXa3h2BS4wb4qLV5IBpel2dzd9QR8PdGqmLHSwz5fVsA6fUSG
9y6rl2sVZjUxqxXLPUShpq8ak9/E3juclXm7sioju1qNgGDsa4Lwo4kC4lmFmm7WzHWWE6LE7HL5
2FfhNXeE0C9u7H9rmpYbJYlGswi7iL+7p7cNBNojRMwbRKJC/QLpPhUGP01KMNjidP4+dLH9Rf0v
V4+9HttymFA34YdFeOjFNcAzjMt8Z5lQovU8/wI67pUcMrLKO77IIamlYCqs4gSsP60t64972F9M
yphw4hXeCXTEUgaB5JQi20Qxvy/0mELyKE4ggqcwVlOrvNETz6zVVZ0Yw05KT6ieryukvsVjlbg9
9DrvmSS6WYQopnDwrh04cTSSqtZnKARrs3GmuTizo+gnP2OG5uSNr0QQgWI0P5UifwsBj33KRy+L
Q2TEK8qs8o10fxKLjFdzIQoYKKBHyGREo9mNGauPqjcZbVeQWRwFQdLOpC6yAubh2AR1Rqg4gXzK
8nzqQRVc8fSl/9WIcZySTCprUWz9p9hoxqU1vuedybTMVtakQsbzZcZ03KvuIEXqgVVNUTg0Uq8H
U8QdGX6ZaaXBGrT2gpNHNhHBkJwl14VxAoo9oDTZlhflkFeJLXpmQJY7t910uaBFELcuusFUkcMw
sQ/JZaS9AZTdn6UvSEf/H2IQhcjovir6OFfQ9xX1w9TmUXHZN9GNaKlLRieerjOExYTV7RkvrjJs
I+jmEGZ+eGLis+ryHPeN/OK5xSEIlxDRTcuPvcL6jukht/CkDlPvBX1v9ohIXAHOID431jGgl8Y+
KJv1ch0EMcpy+QaXhIIkyt4C+sd9nQ9bYybSAujKy5V93TOMTWKfb+M01GnBQa0uQbNQe/G1RSOf
VWK/ifoQkrAmIPGUBck3BzVsktsZwH5/G0Jl0r4Amk8JmMpnyQ+sCDgVDuqKxFcIlZ59kY+HGOgt
n2q5zmrHX2p9Fk9kCb+0qz/yZdbBHW4oZnh/arHzJ9fLvjZ4M0gGQPl6mtLa/ZHnaKsPYNvLftH/
d2HgvMfNN08DpUtkQFmKansT2HK0cNCAG6cBpYTqKJjpzUmz4KoV7yVxBScSwBNJ4YVW8KrAlBKy
8fTzxiSFfr/X5iUZXN5XPatSyMk6fPwNkpyT4GWH9F8hn2x2XgPLWFIoLdqF/OkymKUw+8dMHsDG
mq4jqMvsjARqs12O1bI5j7UZELANremCNP8mj2lxI1/MJsTTP5tX213PKP/DBNi5daezTk9JzUVy
qGRLvDvD8xWllpQLfKImNpYqThQ787HZVDX6W3Pwdi0s5DvxNBWJ5fZCAGdVOf6SoMOrgOjj/POs
jPfIqMRpuqeexRCkTlqnL75rl2M/ZxrTB2D7NKIAMHhrRno4NlASWNbykhoxsErOkFiUWuk8vbrs
s3/XXk5ms1IncqkXbSaN9cs728Ak0qeTT/8fVezU9G3/+wj78GNBwJABZJEQDYtg89RJIX/5x5yR
X4l/eBz4g1CgntgoTIOAtEMMBGWXR12UPfIL+BIiR1czQz4WS52a3Bh4KaQp1JVvnNMXKub8lDYG
wbmYDcGRuUDk2KknZQ4/qZ47YqY33k2nBwMlmx83zsPPn8qoaHTzmOCgBf3/Dc8S4caOLCPjNevz
vbb77pKaZXhsjUMpMTe0mSpNRRFtamUnOyZIfkkE4cVKSlheAlVTD9fS4+bsVCyas1/GjfFAmY+1
X97xqj5AuXOIGR+BAACnfcZ271Kum4tuuLsMhJ0qT1YgZZMvGAchEl9aHnKknI2Gn4xyPYtxnx7K
dOzB5/Gj7TJeSkCYUzSgGb4SNnaUm80uUxcPZkE5fRDWQk7/o8MqMwUgt/KBrlF3RupKq5+zVghH
o04I8tBzWAuvPQxc4ubjoJHtpca8uQteeBxNfDCKCq9UJqt6X6NPfxo84cwO/5ssqcpOpy8bfJqz
P02dNQnDnns3GXJEpEx9WEPce9CctrzJAhsT5b9KkJmeYcNckgTuOPQKz7EPLWqjuRn0/MRdRKGq
CWx6fZZcrHfpPhisQNJFGUrzNue7HcKUjZK1nrtqZxbLP7efYRf47isltddF26sbxXXwLMY15fE/
LKFs5+uRItUds28cqxhjvhyDfUtI2Lm0v5zMPBdI+8827Z/5pJVPbCIGorLh8JvhkK8/FUmC6890
VWO9QF+nLU4YI4KteegyEp3TL0Sgfw5/JQPexDWkBM8oGivi62U5IW/xa4wdV/rIyk4XXk/CKmBd
2KpYGM03vZYfOHS1B8rEwNScSsBh4GXD7rEVnhycZFUu2LsrdKHERanMXZPSJlFMejt7tjtSza/x
LgG5E0+WcB0SCUHQv6jAaEB6bpVqrbmtQG7fBBZl/QfZ5O+7jzSAm5TrajzL9rIXZquUe9kgwPRo
6S6iQwUPJSzTNx1TfvVOM2jn9yfU9HEIqlJW4f2uzrEqquQEETNZIHiQOc59H/FB3ZivZ/r85Ut3
Yo7EmVF6pd00gsvjRfO2TtBqEb4YFxlA3EVMhgefozIKhfo/E/RRig8wDJ5ZBsMx/7ccWi0C57gk
N3fmHl50E9vIVu5CwoaQsVYyVBq1FZbURP3ubim0z+ykhzSQDPePfPBru6wfjseq9fbJ38MQU8Pw
ywtkQ18DHMNarXmAepQo3oiD1HmembBOjMHG/aT5CBKQSShwFB4ZYsoXVfd/cJXpGTKjgXDZRafG
b27/0kEd6juxz4L4UnIzM0WH0j836aLPgdE9yC+CH0zR40pgXSDrhSaN/nsXubIkNH+rGWmjA8eD
ApPplcad+EQ9WpjHzPWh+2dG0BNU25uBTjHiYijeGuMpf3mBX3WUf6QT3WdoHkE3cZ0rOYB1PYHt
J9Al2JbiGF7vRVVGl4mRfo+/yynSWO7CXWMWs1giMW6fFfOgnNaEwNpTLFoX72bP7YJE+v8WMAI3
wL+k+sfVBetahBRG/8Vw4WmP9x18JJ/SsugVYvirz6tzXW+kovmTLdMx8kUfaUbGI6Tbr/z8PrWg
36s2Zr+UyOG5NgD+3wIgyw7ccUSVn3E8SnynBNbI4Kd5Jl6Nlrahpca3AKVEQ2H6o2fDc8EA479U
iqREWcaoE9kLzq8VcEIHIY6Nekn2AH1Y12I6oe55A0LdMGGUSrN39RNet6VripJcpGME937yZT83
FBqj84TqNzr91P8fyY8/7WLkE6LZUJ0BkAm9Y18ehJZxSU/HzW22fBHJ42PtDBG2b/i0jHXkUI1+
Lkq3ucEVb6+bXn8sGP29CwkXHS9IEZhK2PLHDJpd//wNxp6iybIK5Dz92JfG+abWdPNXOunMBfGa
Ln/xUIkdLNmW4NogIxgsxtwkX6karUrjHU2TE356QfASqW8/M0GKIT7D+qyO+mcU3COU/q8eGu3J
apHRxcvz8ju3ijK4nUpq1M9zv3lMXTjK8bBI4CdaWLnBSklqRfjbEQ+xl28gTWcHaMoAYAWPW2WL
kz+iCJlVcWk3YAX0XEN72gwDOFrPWbVNnzif9aZFV8+opAiq6uBJgx8dwMg5wsfMvA+FD9fZOXUo
d2aD5cBgm5VsZVq/eDMjWTa1xIJmdgXdOdsxbQV6Ua1/eU9rQH7CrY2z2FrthqFXsUF868sPAZ1u
czKa746pekfXqrFTAp9RSpo1LBO+KVEinWjgL7CHM9V3MiUop2ephBq4jIEg4yZF00vVr4o59SGG
jZq1tucx9Zy3AQRWW4xVV3ojukAlFcqI7k6Oc+9cN9jza1+AwBLspOG/n/T7Ry+urMrY8GmADpQH
EyYB9wFddNFevPU4MXDzTTFJSfRhOzdbWNW1QPzN5PugobhInMWkzpy6tnxNPimc7C77/dPdPVUv
0wrZ0WLtkn+PdYnhLACKSjO2INhiEPVzRQqqF9aedsNUrfiJmx/7tJfAMuCsOBpJyNWJiwmmULNV
bz0EN4Rhbh2vrNPoJI1C5fweGjyFO8Xew4A/2eCkhXicStXxs1DH/K9eFQxdo/0CcnqfRnL7V6wm
GyYBMevklofAScwePTE7UhfNJmZAaIf1NUClDWFQBRzORBYNvvR1cSP+7BvgKK3jZVIkbKO76AQG
xyS/68R+2by8Cs73gSk8XTbZaeiEwwfnxo1CMUQDdBw2kk+DVcHzyBdRWj4B04xlwc13fEK5wDIP
txjM+VuBg2msew5l0dCdOG1SIu+iB32RXRzmhLoZHTS7WuBMw2nWJuP9nI7z5qi2h2COTr4b9DOK
UG17198sXkKmy5VAiwiUEsish7Lv40voh1boHDqemFEHhUNMYX5EWA/kGd9H4K93PDbxqi6Fgvqb
ar0ccWQ0VLvRc0FaXJJGEObkU5KC23sf4vU47RiL7SvsR8GaPIR5U1RJz+lmnm5UjgqgCuBGdCQE
8XTLereQZXp6GrQqxrdSS/s/f5CRuNNyAsCzIRdbRWnB9kmqW2B6HZqolAQ1Q6H23iCN3Hr7jZ5r
y9+Z8rGdxWLWR8J1YLBKjZKz11H4SB9HDTtmtC4To1IkM/VHs64YmCGSnfrF5vp4iqrKQt/FiO1n
tadI29Yu3tgJ0vqqzwGMOjXd7+BbvVG6GTMBe4uVMP8eXV7FcHZf9mdy8hGwSfYujyFtZ+yS8fz3
XB6VMvHt8VLc0yMBPq6bDux9/0YaiWDFuBvXlQQfP9TJPG1wyEtzIhF2nXtHGSCtMKKcEvnABFwx
QJeIis43NlzqKd6kwttdZQia3g7ckP3fDHD36htAw87XN7h5DnukYU/PABi+kKQBaxGWmYsoL/Io
WldPdCj6TVO9lssotNxFCyGoh8LqeDDoGusOCWFjHSoxyB85iECsimpG5wMnMKjq9gwcLzz1hQPg
ybOtEK8Vrh7eeInqJKg9mTtofNvym7nxPIv2l47q0NPo36/K0Snmr/FbSOhq6rh/296XT5ks5HG7
kkIr5fyItP4yrnwNLmfAPIHFcLntIZmizbmJeh3O1UYIMlxMYwxBrgDoLCymI0XBwxCQh9mN5DF5
q+JhPK1WJCBiofBpFFlqf083wr4fRCIIsh8MzEOd3YbrU1LieCwPkgU4hmFpvOWbAyenJgkw8uM3
hfCK7a9ORRkZEjH0uP/YH+rD3d18bvewAusxVvgOa3Rra8i3E5rdhUzmtA5a/phn/JNnW+CXNPPp
h8hEtVFBwtKUdDRGYchgQg3cBFCUwX1e1tDbqP+jVK11faWAXgSocEeAvduh3kLV3B6z+O8SgQTj
ECsfwuNUq+eytZy81jDjmG4cx7BtzFKWv4c9lfD7zNwDJgQys81vC/59pF26r6XtyidwGkC54Izf
S9iWhi8dJmJTwo7KMQuYKOsu4kndPC+Y9mJnzyWA4Xk+aZzkqQcUuAlY67Lb17Rs9lGl4O3CNpnk
ItxIAF04RJSvz6dcHUMtPfMEYc3Z6evSOiYVcwHEeKxrTpEZaGAyDycVscxC2oxhfT17kWp5pBV/
823XAJW7a59Oh+hNxi1Dm4zz265Qh/ddEiJQqEGh1npL/ZD2dl7h9xiakJJyXlw/+2BhYHoASyaf
xRfHWvm/Be3fuptWKQ/aU8HHJJPpn/lhIr4GNSSR4MM7NRjfhzgnwRlyp+mUiLOgqAxskkntuX52
lYAnSzOf2ehjrP43F6Zow1tpwF2ii3V8v9ZcVuvjHAD+6pNJOYHFXC7cFHJbtKrTDMfPwmnDOmW+
ZcsSIAevX3il0TUKsFv2GSAi/UarfuRHgnkrk8ouOV+VMBw2XkkxdErYToMm9LNAcm2eOZcDc3/F
I3j6+Dcu2Ebszl3QoNhGBmxOYNTs3B4MF4M9AgMg9jlXJVRIjrwwlvzUk7v3mVG/vNdHFTHVClz7
+qlo2Ew3Gt0q/fSb/LfhQ6F868Aux4vS61TuzaerWfa/hnz0+YnPy2MS2k6Pr12udq7oBGSW+jBw
jDYHRZWmXCxlSYpL69i8IqdqHQ2+SAbqAsIB7ehhafEGjWEPr9VRnTqmviqrHY8eM2Zm7HT6ggIq
AO7aD7fmXE1W1hWqbWXCx17nhj6Y7WJX4I2FRSqOK9Kg05UcpK+Qu0eoZpdW5CZMxxC7eiVFCQs2
lW9RxFK86GrtOCg+DUgF98snJAXve7Hz9GWv5b3xAcI/89KD/fPZeXvmFGzFRbp6WnfmzCP+ht6H
DLmiPJ2bzL2mk8qibWoyQjuewD2oTmdajMf80M4x0wxGSBat1IkZX3NaMTIhl1RGjZt+ktx/slZt
7jGdGNNghWzwxvgdwwBVyOZNe7w7VquMKA8UUw7WhFVRq+4Kq+M+jqThnRNmj+eq4YrLcDUiGVp4
GyL+cZqrtN4ANhOK5W9u12MKOzbcpSp4p+ZqNV+iI/roI6BNOtNYTr3dLYnwv89dDo+6ZZyy3n/j
6gwWiWbYlMW5SjUoI1Bb1MtEzNKwFazJPC+c3zPyIiIJRoJV6DPlLNOzgQz9eYM37Gc6lU18A2uh
2RT1ii3ELGBTiimEi7W9XjNHoujtSWzvMFv19TBBt8oYpjuel2UxUT8Kv804ZTFfw9RDSVRKYW20
QWPhjlP9FAgbbE+wU7mNnKQbDKG1HZjkfT4l94WFr/R/ML/cEyQDrfcm7aatu748pjboJvPqGm33
0AZ7YuzvfFdjsstE5MGppTgRI/m0rNn6b3AvUlcazAA2dEGWsJALIsV3zq4vqWtvqscGpzSVlzcQ
nfoEuklkZjTG488/hPuFJN+bDw02DADmKv8EfBqrfF3+WkwPOaubV3DO8hf7MKwWwhlSjWr7/ED8
jEGrxX+dHE4ovd7m0wbnGOqKkDu55HAseGZPZ+auMrL7HZgEWV8YYqjKPTtTmvRXyLbhcKm2QAHI
VqPJUb96hXepl1XI8VaMzYz3eKRZs6SkPRObGhN3fqfyb/38HkkhmCcZd2Jm0YVD1dbGFvPxpZ2k
8StVbUXrrnDCGCKCdRJpR1U5hV0F7i98Qy0+YwK6Z+bIcPOJpAu0k+UXn7hritRWi7BopTBPUwxh
43hDXdvCGPfiJiDfGrmR5eGZEPwLfAVr2ndPsP6ivM55DrxEN4VH+JbX3SYGbMojhXG16QWRYUtv
aROW3I0HXZ1anhRHBQ2YYmGoYJHkzzyFQIWCLCshXeKEpEbt/rp/4VC+CdpEtqtY9dV8SGokxhWs
2Aa06KDGlq8mNQSvwzybfBxGTf9mUps50qM2PvJ4TV73nlpxXVilfkl6sT2xAi0yqFw4m+aUR0cR
aE9fH7qGZqjlAp6S/ecoq6ohCy74Ufl0UWFKEpw4m3d2ZEEAgYbdU9Zj9lS2FKX6XdcmK7q3GDuw
H7nOm1Ho6oF5m7c3nNyztU+3VOKBQwXPqePTN9dEXNzLr8pKGkmqHG9JFK6fiApsI8J7pjSQePMA
jrRatyikKOoePddQCbOI+eySNo2iQJ541F5RoVexmKs6yr7W++mxqChpixTWhMNRuRmSnzOzH4Pl
Lrr3Mj9lxH6KTpfNm04zxmJAIaTzetaYnW+IXVtTeMyYByTr741wecKm41qEziEUuF7eVNAdgF4Z
2sXKZmjhqvKk8cM0d8EqKld6wqdb9VKjwJ7pTPWqytEEWNmDHdX4//VDrfzT2bBrF7DOJ4YpxpyA
gLiKwrTn3lXtkRRtAJzyTZx74LM3r6R7gTx8CZGvdXg66XITNO2Esk3KnyIdNolez5CJFojOl3SC
Wk/34Nkfc33G5q36wSzDbO7Qaz5YrWJ1gZcq0+LOGgBnc7n3Zp5F0+pmEdYcQagiL7/1p7uOiZ/h
AnEPb0eqPLIu1xHmuveHS//eU9tP1Vu4WiiXMCMqH/Y10y5aZVtMajCauOpNrj6YZfknWKOQrsEA
iEUO9++E8CapB1qbnx+fAQQvSItRrY1Ee85OnatfmlvpkW9uqyFXEpQMNDVmBfUoreo2/6fFFhZo
UyfyU4RlBtGd2rbz4xvDJ5rsJhk6ltmY0e8Gk/gHOSgKA9BYQj0Z3eJovTH7CoN0LXQ/IO5hMVXn
FkMz6yv1/4YCL5YXkB94cfH+aNkSebEECs9Z04QL0C+ynqRqU+/QnmKZS+Z4EeMgb3j7j5AEqn2W
kLK4ffOHfJAtVp8sxk20m3eXLnyW2tA30mkAYFyazyQnR0tBRHtAqk7sLlpDL3IKZMx599VOJJlI
U3zRjVYlqIOMWm3bH/3FgDExiUCLwAu0VdsS0JOPr+5c2tlWiGadkxiytz3BwzppBabAQTaZE86V
giq5vhHQWTrLOlcCwDJYpTt2GXNKDNMjSAWoamsvuFuQfEBOGiZrwoT8frDTFTeXlLYFDwfXfFrj
opTd20hnuHU7ihp+q4VvNkz5Pz+DcQFq6BVXc71mQuQpthYZ2T/z0XBpy04vV6FJluZeXTzVsnZV
6euDVG2JP6Suemouwsp7U+rnOXuXNto0zFqnd2fCbDVqa823iY7CWkZKFNeqZTzpapunL4Me6UZN
Jaa1kl1EgtdDcZUp5LnJLBcY4q9rFIjHjV8NPpudrBmdc2Kb/fS1HRLz48uynK6XVA9ODxRQJPSv
1SyzIsBPlw6axjdVxcJmglwO6vDuV8tzIAaAwFH+PrN0hcnFx0nWRAVG6yQbFNY3Ta0agsKjPxc+
Ih1SSzFAOcH8HW80DtpgHBNSpIwhbKE9bRJEqn5yaUcAA51m/2n4cp5hJAevCS8/0YuHG4HOOuJf
mdmtT2EAYfqv8UEpt8CEMJk2PL4jLcLx+FarFfV1e+wUJxHWyV7S7Y9PYJ3oCJbY3Z1Ymb07+EAF
Xae3pJKITfd9zpI5POFt4YuQTGLMyOVforVDMleOPCipQQLEV1CHhGV0sH95b+oxgcPxaSjc0KHx
6Pr/k8leBTmDFaDSILl8kOL9H7MEpFQAorvHKO97E6EFNGV7rc3zylQYdIvsZznASrlP4QzmeM5Z
bSlSeinjOq3uxv88dp9Gb+tR8XSNGIaG9NbTwJAadhkH8aXVkt7SNGB/izX0T+j7bZVaNzALf25t
Ypmz6XYt90rwvebtTBQpyX4KVtTTxw9Ec4l1fjIIpWrcV6XRH7WzhjVFTrpZBAiyYTUjIDsAtA95
fE1YtltmbEaq6yee82/gPGAL0bSTK3BDIKDdnl7TEyHto3aCyxKXRn8wZTbRFDpjoqQ0v9AMMJ5I
wu2GKhRs5weT0Hu94faneTSWW+llSBdFLbwA3yAtL3fHkyuUcxuW6P+s6q0loIPJ7ULBgi6JSao1
aZUIxGD+4T+wfrVzizz15PC4HOpCNOh528yLG0B8MPd+tUr6LXdVERFvw8X/ABa7kbozVjVbYa9a
PNi2kHHKg/RALjrONkh0Lh/7N58VM/gib8rUAhdzuNhB/59B2gPriv0DxTsuHO0a+ai8o/NOArBu
AVIQ/SpnF1WbQzBl8Kas1qUOtmv0vqmo9gbDJWPCfJYNOxU6EOxAlFB+0/m/3nxZfOqlRSbUxK58
lgt+M5vHD3EBF+KaZqM2nSam1rorx9WUalMxdVMfh6aGkrGlX+2B5tMWJVsy+7LHURSLOw0SBQd7
+HpZ8iD6ZtAElImjMW6FYEhMBOjbZ7N2uXxXG0Ht8PKsTkTIbyHgGZiSieIv2wv8Fbm5xG+uR9eS
UDjZwsXUm8Zg+fj4y2IIJxRS+mIPPsW4ObnOfmALt5PM0oLwPXFxe9z02l39fzwoUIRZxKnV641k
yaSn3X/lx/j4eDgY5+rUiuRa37dOh1wT6Oc1TqmiE9/O4AQCQs2l1btxM+Fo+BAt5fwSlnpYp9/g
Ep50KEan9M9bO0eJUeCQzFJVvAkqvU0jbC+Yb+MXjN+v7ZE9oo9FcbLlxE45n7JaRTrqe4+jQ6Ej
mugXaEDBc7rtpWgwRVcRSQ2mvVE1O1sPEabXmztRz5Bn957BxBe6+6BF3XTWl4T8cPceP7F+Q38l
sE+cv2ya1zZL0YxGKtJwWuUC9g1z312rOyfn2YuPcY4UnDWCTTAa9L8X4TD5+qOeH5CTeCHXo6Vw
n4VrTQeGBWIwkVqYvE1Dm+tUl/zIUP1uGmasxXzRvcsqTLQTTTejxRscCxK1C6BF5D+qrzYpzHek
QCwiO+ZjU9q8EbH7zLXYHv/tVg5q9L/RTievF3u1gdAxCE/C4M8Pi29TiObTw0KCxVU7eDMebcgy
PZi7B4aMf/okumA8rW6/MLRzYgDSUxfaTHKwtwcYuw1tcBYjNspwy4I3j8CXrFNp4DKfv8HU++S7
vI7IUPbvxXRDoVFXvkNWvIvnW+rwd0ke9MCDRqywA466/T+B4xtV/8M8ooYniiWf1PbG62RkEca1
CbUq1U+SZ5lldBZLco34v1YQ0f2dGjN2ZmA3Js2e0tcqndcBY2j5rbT2Pry71a/fbWXL7AFj4bfv
uScX9cdU/C2ZOnOFXmU21yjU/pvONJmPmGpr3l7+En8pxm1ECpLtil1e5Q94Tvx47vZHYMw9wPQ6
KDlGCVdZPXBKtIl+i7CDTdcSZknMFiwxLpB7Q4UvrZ5yjTUH0+EZzsTbeUD+zFouOnfbtIf6yO7N
ogTnyU+Z8sRN223d7EhL1Xkqgn1i0CY1sBsQjMnmBYkwdkMgIBSb3XHacy4f/NJAphMGoFDoUC/b
176ZU5blmOcM1pRQHiSh2s+1FgMYD1hE/H7BUjeCc0hA4x+In3qpjBlla2Q7dSlIFZWZXmAYjdJ3
FYK22FEQA08I8uP+ZjUJwOc1k0oUZ8M/FCnWFfQHcpEHDOsOQGCKI1R43wPeGBZWrum/dl+wIVRz
RuC23K41HwLqkisGPDulZSKPV7yT48i7rnJf2RJ6KsSg2DThfbD0eLe3k3ykJtPEBmhpAOt8m3dJ
UU15PpzbmCDriv91qCriao4UmJTIZWk+f4CttSRVw1DUsI0tMEWDKnoaUdGH5zju6HF0qua7cPeL
bNMMKLztGGLYRT8pcweZOfRJvWziFDoIzmg73fyogE88Ayi4QpabwP01R4nBjLxPRZDByKm+WEK6
vYd2f9CiceXhX3Hj1QNZCc/ICzaydbHkaR4jrd22t3+wDztsMeyUezyDyzSUArDKKsjAnypO0MK3
i9kq2kjOIGjoMgcRC6vjY9UZFr1Vk9R9A6krND+dWw6WsXa+9ExjazfNTBebRCDRO9LAZ7GAcKqU
TJms98gPfvtWp6CmYWEtE09K3vsS0JuZ1TbJH1uOQl7z5RqMyup59HGyhDABN4CkYhpc0oFpM1DG
uel6rVarfI/gDXHFK/ShF6z15HVjVm5kFm5RWPqzkPQlaP+o/iLZnKizFnFZagNjdb7+6U46oG1q
xkb4NXgvDRjrhGYwXpyyA4es0z+UdrwsoatyagPdHRq79Jj6JzMQXeUHbAeNM/2lWwNLr9e0ydZh
In/RvavFM7extAe42OX87YuOiI/JpJfWSIvXboYgN9oKy8+R9LkHoNkT/uEcGavCUC4ZvFbU+VEY
bJWRmuYYkTtQNppflamGnTNykcc2Lz3RASZXd1eLysyqIHjysq5qqYY80GskGTL7Y+In2W5XNxQ7
1tSwjZjY9ntM1LMPc+IgNuILAnSz6WG3PKWLWZund8O9bgLdunHTvUtQ9PnhHv/Eh4/IYyCUkDxb
0fg4HN03kJfSJq4T1Wrdh02/ohv7NJOad320mfBAEeWyvPzGKsd0kETbTVHMitIt0tWypTI7Ecgh
i3MEOnBn+Kh5IQEV/nzeNbQvWLoCOqx6hnhOxCbIgIh7LWs7rGUhlUiZWERwoKYrnECVKzrNzdnZ
dNasVSIuJae7vtf0qDutks2QEbcrijOG0Cbjk1qfxuQSMtptWrN5lsG6+Y8C+/zYUtcjnG6uEiOI
kljYxyXSv8i8LDtZvb6SRyJtdowYzHuw4Cdbb/EbIGfQjAm5iotPlHWBN49gdCj6DuYcLdE0CM0X
jVDJq43YKQQncEMjFxWeXsD72M0lQFK46Fshlz55XUC7W6ryAvD2vtmCh52A2rHQToVWMySTMgkR
a/rXOT8+PFBP9bZDBACTpfHIOj6KuYFOL2ig+Q4mUx4T/QtDOZ2KcJylmJdnOkC22ryeApyIgHTy
lsBGRNodhszBMa4kPtyboAPfi8mwAb2K3fnLYJg4TqBGrha9SGH4G+zUx31Ei9ksJKoSn50r0M1a
NAt/qr87DDPB3pUsuRf2Y/ap5LrTn+IqSNEkLzxYJ88lmtvqoinXvc3jZiAjFsxSKMdbwdcxJOkk
VyrcIKcxlk42EgMwF4ACjGzp5ku76w1g3FrJ7bp2JF17kxnHQiunAvlEgCD6ANTx+r/xf7GV8QkK
H3GO52wBsykMWSNJqbxmBiuG/HzKr34KvxK1N9ieOCQ3hDnuVL3ioRer1ujy5l//gQbQFBoIm+i1
Hz/4AzdP5PIzIQuwYKvMtPzzPSkt7VDfMivTd+IF3SmiDudDLT+qL5Qkp7Oxthn5ksxfjbJP3JFp
a/0yroFPGN3I06SQnQ3y8BiPsjCo9mFk6zYaFT5Hb5obIz1fgds7jbgNs98JrdEJqUaMOFBKwxkH
JaTV5Zn8Z0fC8TahgRllHUR++6/9qYQYugC5nebysKc8YGg7ofR48GuvcR59VVbv0BPUd5zhO536
pQvnoRV+FvquWg+t5YWg2kq5sK+d+0eDya/G9/WQ4Myh3ufbNLuLoKzaAmSJ3CwNowvBPKoyoysM
WjoV7j3egoxCX5XNyqo0PoMAZtfY4GV5QRvt8kTG/VLRCss63s/sbLCW9sNbLhOHjfHddAJwRbQj
6JymKvAqaHffl8LWO8t5ExXZT8b7E15SGI6TCzr1kSEBIxmZ+y5hcC4bYoGLkAZUmFIsFREj8PUS
u5xhEvCz7rOSv2QYe7AMYQwRhuUH7xYPRu4Q3WJ9jus9Nxv+aCzIQ23ic3K6VtGLOYFPHf4TnNHf
bFMoyEjJ/v7rFVUS+E9IG3yah6sz7J2gBSBTHno68tBzgXIp6lIDLW8YGHVof7jWqQsfaOZDiJ3J
ubnbHh0btJwH2PxtSw26M01MjJt/icrEFCVHA3BjfRY3RLAB8/+GK7sbKBakmt/yahmPcNqimY3d
LMku88Gvp4hoC7Ugx2ozskYRAzhH1FMYwBso7FS1vHs01vSh0rtT7RtBnFq+B3/pKrn4xNkuZ3jy
r4/H1z9Pp5CK+7hauDI0IS4ycOYR2JBXD+GmT7KwWCErpUGKEMYWSWOSyq0qN3A/sxqjBYeYgdG5
v9zfW2G+yz8jgkxsSSW5nr2BPR9PHrQ2wiCow9dbrFsg2hDdCw2kB7GQwoSfbeOycwWrQgHXmI7S
gFpa5WADUW/6vJywPVtpic/y1SyawfZ6gRHoAUiLe/dJ8NYCS17gGqd2D7/hzrqGdBa/8YmzTesT
SWg7h1ksoy7VVBqP8k1F09+njr3nPU/dj/0s4wiscpSy6sg3ZW7uJ8rS45C5WxpS+KOIOJsMy+Bd
BB7GB6/gl8PwrRvkFphrWHa/D+KnanpC0ZnYaI0CQ+tCTrnEb3UaD+ZO7rJsbMje4C85EQWEzk+e
W+n85xB+i6JJ26sgN6IVcsiEAQvZ5dR6B1HFvx2al6lITTXlJr2JHGdxq6XGLp0WujkzVrlNB0hI
yccLATXM8NBbL7o2KX04h+Yj883MD/KrEC2Jh1xVnzQHDCXuvTU1SAF5AZT7jLQrhQHXETcKEenz
ejLwKWkgEr3cgVqvE5tCQ8JR/yyzZ6Xljhuq4/jKrGK0mpJcqRXt/mAZJ4jp2jqIpBaKyb8PqLe4
qR8cb4V2RNA+i6QHT2cp6Wj2r/Qiw6uR2mV5w2XUx98J1P7AKo75aXcrNOCXEGctkd4rCadYdVPq
KyYV0n7cgKzyklmBWMB4WNE/og2UHsRWuMXF+EhLpgJCeYPeiXo5Qqzdzbjsjvriaqz8tFuY6Uji
2jjIoRU/yEs2gCzo6zV5ig/BfIhxbevgXNQxGeM/0s+YL2FezdeDSxxMe9AR0MDU2MmhRG3HroUS
9wKEBPxzVtrcFmkNi0afc5gtyp3eojDWnqWa6WdEjlu47+6xxY1oxJNFZ7AcaCKUg+q3ysucum01
Rw7tz0tqvDf0k5tHoTO/vPsW8M/USZr1X/b8aEVpTcswUwj1NQ2IMOMMBNVBvun4nGBQZZEzb1do
IiiITHVjC0GF50x9RuMQZYXyEtwXMlQQKYyEba1sNy4G6Wq3BoRWuYBlbQE4fqvdNUiRQzq79/ce
Qc4pf16NGyD65GQyxIH4TFd4lfRRV7S4aiF6Z7VRoq6I8kMk+SzVC94HbasJTcTvz5e5CZ6+CHOS
uVPmz6sv+41Te7S4LRW+Cssd7A7yXFyJryFiLvJPFsM/PNPr3Sgj16oQCiYlJcurkpi6sn7ZgZAU
7MLue7MhPCYZ92P+nJu/UHkvve1YNa8v+G61VaTRiaYdmdADeDZp2MxiOwVkdx0um9WdMdSl8u7s
fp8U2E8pJjnIAyNpqEprVf/V83FM8IIPfnieEgn17ugt2FNSf6TA/PIVvmAlMWAIZe5iBeUyT3B4
OSQRDlgXyDfHu0PaPjfO0IbY07H4tYyH8W2LoY+752S4wtWf4334sD2aI484iwbYzn3EqDWkyQkx
6iH4aJfZTLD5x/vpPMqlZLKX1PR6JMeU/OTvNKmUsXwKh0xeZCYKlKSh25e9rhLtLdOqdltoi9an
AkJSETUGoQobjU9SMjW7SGfaN52jhRVmFuIpGknQk35VTjaleWHnDG3zVlCS6XLd1olVYQ5yvdPa
L+w8Qw8TIVCujdUH7QVz4Y43mWZf+FambhHMOP2FSHajljp6J0MJsL9kQNu8iJkKjgOGBbct3oqD
L14gWXPMmbMVDVfBdE2zVFk59HIFOCpKzW4CTo7bTAxFhum6T4t5wQk4fe8omaP1r+57VgjgJoqB
OME8mCKe14PUugvNuPJx5NUzh/pplFg/TV7iEuT4J5Cf0ry7kqVpPjoG4ClTJMj+WuF36i/xsjcb
6SIadVIZeWhE2InYsSaW3Ue/dcwxzglH5nyxJpUH/DaAE/VXbtFpv6bPjRJDkmtK/Rqndl74Ab0R
COIsSzlmTKyeUk/eU54UTk8tPQygNc/Gp/VnIVdaPYcDWvKety/gLJlg1DKCRXZrEOeC21B9HYCi
nIbiNdCPqMSArNoLPgMzYCyUPl3IqNMfNN2LBIQFqkZyPuxG6L6ONRIZbpgxPZzHB2PgZTHWuy85
nvaG5IzNDdO0tNfK+mk+/87HJ42wxMWMkZ5po+8DhxCTQynxE24Ne24+d4CI83hNPs3qmppUBKT+
77QL6erk1YN/sfeV6UGedvIHqIZ/+RZkXDoADIEiYbRUSDqF+buh1n8s6t3hlSn58xCqTkZMsSbd
+qUQOD/wCR5tZOZ3P6jXnJjrEg/StjCcl/VT7mAp9+kO+3BoqKBZ+zIQFdAVJYP/CY9vmg0BjW7Q
hQi0GUYeuG7qOsNKC+vgnEtlXTypNabIv/zqXi9Wod1J91PJTR+IFx1vhFgrcM6Wgwtl+tTQLN6H
Hxeg3Lzc7VZfF1y/hw7ehayoOe4m7dhzNzuucLNCcosBrrEhY4jHZWIl30QM9zpljh2wQA3n6JQ0
ISXX1CPlSVhZqjOttZe4rV77Ac+AMhix6sk8A4hvo1dxhTGxibLt0yZywZX/kU1XaQxY3nYb7aGf
a+En7aZA9bi9YxZ8POlG538YvxM6wQhq/gzkbNdBUQSuQfgTskRXxubK2MHPfcVFlHqiUqLeVE9a
kWea+XSQddK3ne2cs3ryLEMBbm2s2QsFO5wFdmHJmMOlW4myZfQjuLbbkESvKnSJzofBSHL4MLUQ
zVj0Ykr0+QongJF1YT4rMCAXZU6Y/emGo9CVb9moEWJ2IjaiEMr9E/CDWXQF7+3lHG3o82N2HZz0
IdAO9MORllguO42vc1GU8tMbT9p2nXHzVTBN3lqjeoaLX82UxaJkeKQn+7j2Nsqz3lhT813GaGfl
lDG+NSDwxfWjDWUOjyqyX99o3WP2rIrZCzasdkDzIM2e5MN0k7JlifEOla7QPf885/ed2oSOOMq2
P0ewBaC8x9+XF40likYEY7fPgjNHkQZMOzgDs/5Bbo8Qp4MH7XHN6zijUnKFprfLh0qASmpBPPnl
Mb30TYv3NHYCq6NcPFqxERDz/NP2f0380m015AxVacoAMDho/3b+Oyx0wTu8x0/YrwxPm2Zje6LR
UeH1dPfx3/uAlhYzvvx+q4grlPo0j0mMRCKMIDd8TaZCte1D4gcDqW7aiEAhX9taAhhBGT6MvpTC
JrIG1wJjzaL2FXNpKGbcK3/VSgmecLOq2fscA5YTEMZZAQ0FVLa1jl7YFM4jwGZgGDEVgOLr/6dO
c7vQ7g0dGIe6eGEr6Py/VX4Ap7St5ZbYu9BPmu8ElJAoGJum9IIgh6R9mDKQg+sE2mW2W9J3eWH/
FF43gSigUodcMg+Abt4RufRX7tyzXVOlN7opT8Xphug9cYcP5HCzmI/ZghnuSKqZfSD0KHO77etI
Fz5u2oT8gD8HtDsh0eB1KQJM1/Rjn2DpUNjWRE4vzGJ0iJcZIyTe/1EFwZVyuU74KAwTRXDPhnNq
2oocGLkFunr3kV+swSsevVFjYSKdMoKcVmt7S2JUsLyeodpTgosw/4iffdMpm2gXYjzQ3mlkDTPv
Z4pDswGlJKOEjWav2FKM/lURx8IwmXPv4ZM4yn/8hmGge14Hae9dkFqCF6uPnC5lbWKr1sNCSgf4
xr/a0tlngJle29wIGfknwo3H1VrIQUGF0gDg9qfSfGF/QbKoEPty13HBEwE7iQGiSHXZy/moda7o
nwC7ndNQnfROG8DusheRMC/YRHwUFJFJ2bRmD2rBewhvGdrCgwGRMkLxROoz39G/bujIB15Y27dQ
WJSDrKn5Ymz/wlUFs+Kzeug/7xpSJasVpeJnvXFs65RipEOv15THFivcFKWv5jJrjrtmMk7bnUjT
2YKEU6kbxuDphw+WfEN9uCdhtFVibNqkjqxKlOoD/EnJIftwIZv8BcsiD5lMM8NEEFWuGaFLQfh3
sBwOfwEv19/nv5FMPV0JAXQY+Xn6KxvYgw/b8yF8sNWrTVdvxGoYxvV7e+mwWQAeMpuU4ohsIZyE
fh9gvKoAXT80/GG9IBDoGfuT1zgIzcQ6q7hwMvAwVJFubaUcxqW2sSVcJx4pF/ZKA8Ts0zjJ2fLt
JeAuy5UG+uDm96//5/02xsb4IiEBVt4p9w1RunY3zr7zvIxiepBrmAnFeu/Farfl02DdHutkGxRB
E4UovA3imY98V9EJKMhguJs/dJJRQsZsp298OcpqsNrAyXCiDhTNJl/Xi/6gBWtElG1mtLrOsnCE
sx8Xdq4uk0MwBAp9S9JtfASjelf01gq6kh1wfBhh58w1dqbdiuZw8QiNyhk4LRTO2AP23wUpTZBJ
h00Pg/UAnifcQL4a+2qy14QI6iPhU39PWeEe0zEQEGIGqySaPFt6QbdipS6BC424zHV+72RWeoU3
PULeFNRiWgpd+X9m268NkufwwsxyrjJrHBPr7Pp8PCkpuISNqaXg0DvpUDt/mdhtxRG7JJXgHRGX
7amzwAZVNZfMdZv/kmJPjYlp+Tl8HQ9/xLHzAZB5HSl742bjnesNt9yTEj5LZ7WN2rhEmQZZ5ixm
/egbn8/e/BbGhwCg30sjS12E2micG559O3wvV7yP+45XoIutLtpSMs4HLk4+T5O2vl9BI501q5Pq
69jBMvEmOFEF6XN7vPleP2h+lYV5lH5MLmHiCktJzgnPU5dgp3vQ0TNGKKDaqtDAD1FtDL9pmEJZ
JBvA4ogQ3E+ESpI+s58wDOS4L9upYkgqvjaJ8JTrzdaJ7vAzKzV3giy5GN6VmZ2Nw2aTHZ9nyf3Q
kqj8sGCZYy7j+Qo6CFmEn98+gaD/MZlYY9Qrd3WH72Q6hG9uDmSKp5fzJfYwOHZdO9UuEtzQQNYF
J5AzCBStJR5a9pTW4yQXM9qYnlQ/Ztkucmusu3cMFDvxq4fMaYlNBlPcSEp/2p90zJnFWBIDi+A/
5nl9hIB9KRosRhN0Ip1MRCJrb52qWT5lCGRsz0O9vlFAqPZnnis+tQkFCo2ksZqKXsH1N2UUOSH/
WpOgrZqu7qm1R6Vl3SV6m8GB3YJxzE4ZLO1CGmHqMk4AzJTarZtiAXPceTvYAbGNqG5K9ieN0teS
Anyml6qFbeZceBPnFeS2wawBhvCibUHEZL1AxsHbcaIxuLbcJdt9MtPkf37yLw7QFgeA6Dy3h5/P
Ju+GRMzS4IW3Tk2Jz8jsp+TO0ewH1BWHlxoRse3JJvPh5HHUcMpqfWzg1ZpgcLTpBrQ68xetbQuS
h83VdQ6hTY3co2FX8o8ivf/HhcMHUEYapg6DGermGsvh/iCRZdBRldnQFLrY1POEki5ZT8uu34YA
lWxsfvt2p/bJDM4dEpItMIQE4GLkaR+q7Ago0mGd75/7RllwQ2+9s98fWuHCXSG9BBY0EePNUzMJ
+fTMlkMsMY5b1beDyNGrc0oWtkHK9TQgWUEZdRYZce1HGuNzDsDDNw38No/ktXt79mdjunhEoldn
Jms7Fj+m1r2WX2hr8IYOkEM1SzxcyBtu9sHkXeyVwVGe6jzZK6VL9EVP9VoPzYxVHfhw2wvIHgXf
oH3gVFyo3SFMNdkDuDL3AhiS6KiD/DtTHaTabNmafzXqAgLzmoVdt2+RfVHcsElZ/y3lUVyzTyXH
gYKbmMK1tj6rGBugHGwRxyF2+udUnZUmpn6cBF80tJJsSr1z9TtmclLAxqSKdt4Oe/AFa5FNNDX+
hi0Ow/bSvwORJhUXdqA9W7tm+VVLoCkfp8ngqJ0ecJanLcvkSKVdp2D4G/oNBjZiYyZ0C/zTRPEZ
UljETfUlWM/ExdTYQzXmItxtDbMMV9zFJLU3Y3R3V015wYyTsd96zQ88eEQdUPvnZDpSw2gXOV+3
aBWU2nNehZlcD7269zW6HUfepk5YKUsBLaL92jlcIGCCtOU4KiifzEK28zP8vIvrxczkORjmf7Jg
7bk0MAjx3Y1qeKPCNbEHgdS663cZR9MgJWIjZA8ULFJLCnCGxG6k4L03WeSFfpMSitC0yfgf3DL8
oFGHJFSi8bYUhNOrPAfwV+t39S7m34odrIZ5KIZfCT628upA2mwZakfyp3xuzEY4JbhLUqeeJ4O/
gsC4WtA9Fd20CuXFBfkOplpw/phMcX6HR/n6W11SjqabSyT45OGl1Y8XU3SA9m+Jyj7fw06WS8x+
buTun+KGn3DG5lQt/67zJYM3Vd7Nv/gjgZpvngafcQCtHp2hkHWVnslAVQ3mYchrxw5AZZnVWv3K
9V6ag2jIlr6+jjv/AJdZae2LlPvxWRs6GFz7yrDbNkaM0NFPVDUvLI32A8R16I1u9eLLongQ/hVF
jOQi9NyDnQ5K2aJ4OeRxR46zOY/Hl3wkBdhce2FiLQ3TAsbj3Mivs2ef3q5kuGL78CgqZJ8git+p
W2HlTaJwNUbrXaHKsz9eGIIJgi08szI5no+dVBiB8SoKbQa/71rCnEhmKJ3pCmzLYI96jK3Zxc10
aIPrTr7W+Xs6sJHVHcIE6nu5lE6tMMHPaA/gB96qCcoQuGJtY0O/GbBxUO0p4j1RHg/2wJR7Ktkv
ZXfAh4W5wDWowo2DKJW78mGDvgoGRW8naypNuq3/yp2JrJtMeahEp3TKwp54ovjPm0Fz0vxfcM70
C78CaSe5WahE1SRrlSBBDWShHnwx+M3IDHNzgpXwVURqyUgBts9ybAgvJ4CDjTk139OujwVbGXEJ
hEeXJ2Pmmi/B5Mo6BJ9TEufLbhVfKxFjeB+hvFD/wvkM0ncNSztg61I5sHVL9PqYUC1/D+mt2+uR
uD2r0a9aHzib5FR605CXD5XmdJ97y95lGTKeSt7btyMk6RIAibaziD9nW0b+WKEOrTT+D49btnx5
EThJ6mDUC9oq40rJF8Mxnz1PRbTkCL/jPyjm6HFQbls+JVTREjixqgLTGKKTEv9tjgJX9fZQvCl1
EUXWynrJLmlEdkyKCJtxO8bJ+MXZIAzIA+Wa8W1fmw8lKsUQfGdKO4cYuwZigMxiDN7Svarnv1Gb
4cJeeQj6/xMn670iReSp4PHOzZtpguyJx/q7FBHK60rlX59mPx8iWLVU5pt/vWKL69Avl2YZaHRf
dfAjbCfOqyzQfa2iSo1jfkaqsG6APZRqbJ0OBjWU6uxF1d6Sa59GagV0OnKApMToxVpqbA1ek2Zq
O6OMGC66kjL1DerTNOKCuWQQEZzE9hCMRVNLGnSxSJRsUpoA4KnEBdyQzFLp/OR38H/xAY+L90wy
wfBTLEUV1e+kMVTkSglj9LeP8R/ZVzkVhUyuGOEIYxfUzM7fGC6PvBNgXN8wqzXIVj0i1j3HM0Ma
60vA+hcLWunJTU7MK44QqnGAIWybgDpptendCcwAK5/LFiHDoqYumHXnbfiejyKdlBBYMtNmEeH6
80O8d4QQ9yyg7IVBcFwiY3MMnSR5LaXiNe9/62vOsAXbL87dNQY7mPjayyKGXlsGhWk7RZ+cYh9s
OSIi1X9T4deBSdL8N8CmcIdIQre1P9UonCkNNZ4XNNP9VoH9KAZpcVsLhgQHL0WGWJGKEntaJjbu
NWoVT/iVGsx75nqELyiGhwKtss/EPgAP+HFUZ49sn4JeutygAaX60BBypUBxslwgWVDZ0g+D8tdb
boWzqUFTSkpLIen0IpXdPKWrRVCErMxpsHfJO+e5Qfxq2Jk/37t/M5nVzVnSLsuzwLXdao2UWvNG
A0yB+J/AFWJDZIL7vAYGHkwF49iJP6CPFyCu5iFurZBK1Z6jge4XGH7RfZquOTi9hrF3afpy4Mfj
3AC/7eKnP5IJe9Nxtcarc3HRSPMQiGud+TNMNYFyXW6O6tp7HN4lD/bzFx6YukNtXui+mZQS+f1O
liM9gw2EgxZJq20MvZClm9vQPebNgIraPjzztB11oP0yWAvyLNqRMLvIIfCZxC9GzAfjxTyznVXj
z/L55rDEoP0NY/ErRPgl9BwNHF5fq0itwwIEmdKvCtRW4FUvY8jUmSYtqu9SogwDTIzL2iLAkowK
Xof3+wkrD8y6c9CdXUSr8jsf48lT2VE2chLh8AmQCa/gwbAwa26LqNGsBpomUA/Rxhf/H4Du3wgm
R3TJ5+HEYcZ76A/yqQyo1shcS2Kry4wmqmd7TpRWFWFBFqtG51DQmowap4Sg2EMVL89si4YoVfgB
3Q8QlOPTGM62eff6W+9lDzCjhqQKdXEEFZxqLj3CouGlplc/yiCyMPrcKtoJ7H831piaeZa8DbNH
39aAwHKwkEuN5+XufraooRbSxC+GCcTrHegPKMwHZLCtg5mm5xa9+uZpAHpN0SnkUYO5lbCgLCAu
RQPnCt0WUqLExF9q61d6UW4Z2ReO6m1nnl2lLYiDbpavnegRZw1RPjgOcJi4D5PpyqVSlwGHHHXH
9uVuTWA1hVH70hBf2Cc1HJNBNjPcqGLjIJLG11BDxuazw/gaWLiXG5mvxLmgsg6sApCvVIZ3t5D1
/1zFwDw0N1I0wFVJ6+HzfVas/BBLib6HGpDw9WZ+

`protect end_protected

